H   E���}H@                        m��b�@                        �%�J6;@H      �      �         �  v���)��Ɠ��h����2w���*�!C������U�U������7�ʾ�@���ܣ��J���量>õ�v�ҾO1�w�'�Jaf��X��'���::������/��w<�����������R����f�3�$����V,�p��1HF��ŉ��Q����������hr���\���"���9��~�[��P�lpƿ�ن���?������������죡��!����������e྇�^9�܅���Ľ����e9S�?e�������X��?���qV������I��1x��m�M����>|�	o�����h^����������@�� r��M���������JƉ��WB�0K�ǽ���jo��T-�+��V�־a?���&���s������K7�� KǾ��ﾻ���
N�nl��5+ٿQ#�*�m�wܡ�W�������<����G��Y4������ڈ����7����Y��CS��1��x�D���K����N����(������P���z2w�}�*��B�a���I�U�p������'�ʾ\>��}ڣ�tH��u����z�Ҿl0���'��`f��X�����::������/��|<�����������4���щf�ٕ$�,���+����GF�Qŉ��Q��\���`���>r���\���"���9��D�[��P�pƿ�ن��?�A�~����󖫾���"��$�������Z���^9�C���Ž�Ƶ��9S�he�������X��q����V���������ix����M�k��}��o������^����������@��)r��P���������LƉ��WB�HK����~ko��U-�&��{�־�A���(��Wv������9��CMǾ������N��l���+ٿOQ#�y�m��ܡ�����"���y����G���4�����+�����7�e������S�1�x�YD���K��E���  �  >�����ѱ��,���G�l��l$���ܿ8G��J$U���w���о�=�������뤾x���NϺ�T�׾�s�z�(��e��9���h��3��~�,�������r���l����X��%ƽ��9���=]����u�����翱�
�X�>����rʬ��e��џ���������J̹��Ñ��S��/�}����L���2@������K�žB|���N���ȥ��׮���¾z徽���9��8��#k��K�	�L�J��(����������	��Y���Ш��)������E��H�, ����b��2U�Y����������6������p`������r�����:�|f��d<��'�m��R.�A���ܾR�������������,��=r̾&����w���M��N���Xӿ�n�D9d�����n���b���Z����/���_���ݣ�z�v���0�F>�5������H`*���m�>W����������������������l��l$�,�ܿ�F��x#U���%u���о�;��E���S餾6���"ͺ�N�׾s���(�0e�M9���h��3��~�3�������w���j����X��ƽ��9��T=]�A���������I�
��>����Bʬ�\e��������������&̹��Ñ�IS��/�+���CL��62@����<��žA|���N��;ɥ�wخ���¾o �R���9�e9���k����	���J��(������į���	����������)��*���i�E�bI��ǒ���(3U�{�����������?������p`������u�����:��f���<���m��S.�?���ܾ[T������������.���t̾Y���y���M�|O��aYӿ�n��9d�����������������+0��<`��ޣ��v���0��>�l������`*�w�m�zW��ף�� ���  �  >D��e`��nu���5����Q�$��A�̿��U��W%����2ᾙ^ƾ	���ȅ���깾U7˾�龞��3f.�{�c����8޿�m �.a�Q��4ѳ���������K����ަ�\E���C�y����޿��ӿו��yX)�B�h�����w(���y��D5���׾���K����;�{��&۵�O���TC�-B�2����־�1�����{���j��n�ӾcV�����=���{�q宿XG��B�4�"�x�Lk���Q���k��t���m���ӛ�O�p���/����tտ�ۿ�Y	���<�J��F���8��tY���6��W̶������h��&��|�o���Ãk�OB3����UF�X�;qF�����ᚶ�0)ľD�ݾ6���!��kO�8΋��Ŀ��10J��?��e���`���!���������w0����Y����#����ѿG��R��1R�f;��1���n���D��C`��Ru���5����Q������̿���U��V%����0�V\ƾ����h���,蹾5˾�龧��_e.���c����n8޿�m �1a�V��:ѳ���������@����ަ�?E����C�#���޿��ӿ���X)���h�����J(��~y��5���׾�����J��ř;�L���ڵ��N��9TC��A��1����־�1��2��|��ik��/�ӾVW�������=���{��宿�G����4�r�x�xk���Q���k����������ӛ���p�.�/��Vuտ�ۿAZ	�>�<�%J��4F���8��}Y���6��X̶������h��&�}翿�����k�=C3�����H��;�H������T����+ľ��ݾR��	 !��lO��΋���Ŀ��~0J��?�����a���!����������0��)�Y����Y���ѿj ���2R��;��e��������  �  &#���
��Y���+d���-��t��E�������x_�Ҟ5����������"ӾZ$ξ��վЂ�
���q�ͷ=��j�����g�ȿ����9��Vp�����ġ�Gԥ�T��ة���bV��� ��\�%����:����Կ7.���=�9�u����U��bI���ٙ������Q�JV��
��M��o�����O�U�*�q�����	�ݾ<оeTϾ�k۾J)����b'��K��7~�q	���4޿(	��K�����ؗ�'���Y��"�����{�-�C�Y�O�ڿ)����ۼ��K��8��P�F˃�'!���i��0���x��9Xv���?�)��pzϿ�5��'!q���A�� �&�s���׾4_ξ��Ѿ"B�Q=��߿���1��Z�Y�����������R(��	^��q���s����������Ŏ�	<i�ʚ1��!���ʿ�ѵ���ƿG�����+�,�b�L)��ZS���"���
��=��\+d���-�)t��袻����w_�ޝ5�ۋ����h��n Ӿ�!ξ,�վ]�����yp�޶=�@�j�H���4�ȿx���9��Vp�����ġ�Cԥ�I��ĩ��abV�z� �Q\�r���:���Կ�-�3�=�ݡu�譓�+��;I��mٙ����d�Q�V�+
濩M��0���N�O��*��p�a���
�ݾlо�TϾ=l۾
*������'��K��8~��	��5޿o	�_�K�����ؗ�W������U����{���C���$�ڿ����Zܼ�GL�09�4P�^˃�7!���i��6���x��CXv���?�B���zϿ(6��	"q���A�� �?'�����׾�aξ8�Ѿ�D⾬?������1��Z���� ������;S(�K
^��q��.t��9������,Ǝ��<i�^�1�W"���ʿ�ҵ���ƿP���.�+���b��)���S���  �  {�v��+m�$:S��K0����t;߿"�������}���X��89�^��_�Y���۰��E��#�Ok$��?�B`��`��S����p��(��Z}��a8�$Z��p�Hv��ug���H�n!����EF��+���8��˩���Nۿ����7�)S[���q�A�u�Df�k%H��.$��[��-Ͽ,ʨ��S���zp���M���/�����p��U���W��{��y���,��J��Ml�y����J��\7ʿ�����0 ��HD�NKc�U�t�Zs��^��;�!G�l��|������O ���c���%�*�(jD��d��ku��nr��L]�3d<��U������ˬ��8ą�2d�uC�u-'��(�ng�f��������	�Ô��6�P�T�y�����m1��l�ٿ�]	��>,���O�R�j���v��nn�8T���.������ο�˥����ۢ�^�ȿ2���Q*��rP��Sl�/�v�V+m��9S��K0�W��;߿���&����}���X��79�.�=^�����&����C��"�j$���?��@`�~`��􉛿�p�����M}��a8�!Z��p�<v�|ug�d�H��m!������E������������/NۿC����7��R[�H�q���u��
f�,%H�k.$��[��-Ͽ�ɨ��S���zp�h�M�y�/�����p��U��XX�����qy��,�&J�UNl�ۼ��K���7ʿ%����0 �;ID��Kc���t�cZs�Q�^���;��G�<��H��������;d��&�g�XjD�6�d�lu��nr��L]�Dd<�
V�'����8����ą�;3d��C��.'��)��h�%��V����	�����6�`�T�y�z����1���ٿ�]	��>,��O���j�j�v�!on��8T�"�.�����ο�̥����ܢ�Y�ȿ���XR*�sP�Tl��  �  �M,��Z(���-`	�����;ֿD\¿�����V���b���Ds�E�N�^A1�>��T��[�!�p�6�'8V�>�{�M����O���=��X\ƿ�|ۿn���Wd���'/*�l�+�	!�ŭ�N翶����9����|�xu�燿2����5ѿn��0��U(��A,��$��Z�9t��$�� Ͽ���������4���ˆ��yf���C���)�F�������'��]@��Ob����`�����>ú�̾̿��:��c�S#�v�+�^)�� ���~�ֿ����m���Xv�I.z�����򲿓�ῌ
��.���*�a�*�m; ��f�����@޿FnȿA���B���ߓ��.��,Z�%�9���#�(�����k�.�W�J�$�n��1���P������k����ӿI��a��.�B'��o,���%��F��E��Σƿ�ŝ��u����s�������&���������-\$��M,�wZ(�x��_	����;ֿ�[¿����aV��b���Cs��N�@1����۟���!���6��6V���{�����1O��l=���[ƿ?|ۿ?���Gd���/*�Z�+��!�����M�:���9����|�+u�g懿����<5ѿ������T(��A,���$�\Z�t�-$習 ϿV�������n4���ˆ��yf���C���)�_����Й'�K^@�(Pb�S������<���ú�D�̿]係���c�YS#���+�t^)�\!�P��F�ֿ����Yn��)Zv��/z�@���	�ῼ
�/��*�x�*��; ��f�I����@޿�nȿ���BC��R����/���-Z���9�)�#������ .���J�K�n�`2��vQ������k���ӿƑ��a�/�`B'�p,�O�%�5G��F��Фƿ�Ɲ��v����s����������Z��&���\$��  �  �=�L�?��4�S�H��=L󿄹�߿~�ƿ�����L��%rg��J��A���N��p��x��${�� �̿��� ���+�+����t����)�V��ܿ�������q܆��3a��/G��XB�$S���w��C������pYѿ������\��GN���aH�O���-���>ؿ ��@�����8z[���D���C�n�W�����+��������տ^^�=m�{s�߫��c��8��2�%��Y.Կ���������}��IV��&C���E��R]�k ��,������ɋٿ�����"��Q��L����S�����Ͽ�㲿Q���-ju���Q�h	B��H��8c��Q���=����ÿ�Fݿ���:�iN�[�����q2�;�+�����g˿�ĭ�g揿�/n���M�4�A��/K�,�i�:Ќ��Y��kPȿ���=￟K�إ�\4�`S�����K���.�߿�ƿ����K���pg�ZJ�h�A���N�@�p��w��az��J�̿���s��u+�������@��~��)�%���ܿV��������ۆ��2a�w.G�jWB��"S�F�w��B������Xѿ��>������M￪��
H��i������>ؿ����,�����<z[���D�֨C���W�;���+��򨹿M�տ�^鿥m��s�_��6�����؛�2�֋�/ԿI���[���U}�KV��'C�דE�T]�� ���,������ٿ��M��`����쿶�￙��S��忽�Ͽq䲿 ����ku���Q��
B�H�	:c�7R��2>���ÿGݿ|��Z;��N�ʚ�` ��2�;�Y,���⿪h˿�ŭ�T珿�1n�o�M��A��1K��i�ь��Z��Qȿ)���  �  �|��4XÿP�׿O��`
������(�F.,�!�#�ώ�?��g��FI������s��~������1?ɿl��Uz�f�&��r,�I�&��=�]d�����ҿ>v���ʮ�qL��R����l�}	I��]-�
�I�J�$���;��/\�I��n񔿩:�������|ɿ�߿�h��`g�`	!�*8+�=�*�]6����޿[���<����y�&w�&ŋ�k(���_ٿ���:/���)�S�+�`�"��e��� �]��{�˿ֹ�%�����v|���?`�ֶ>�-�&�����v�*�f|E�Гh��凿�=���쬿ܐ���(п��7m�
S�"h%�^[,��'�6��,^ �Q�ο���T����t��*~�gܔ����꿠���!���+���)�����b�R%��#ڿ�WſnR��!S�������y�JCT�~r5�y!�U����m�2�EmP�]nu�2y���V��/|���Wÿ�׿���i`
�W��p�(�.,�ߓ#������￮��}H�������s��}�����N>ɿ����y��&�zr,��&�z=�/d����چҿv��\ʮ�+L�������l��I��\-���%��$���;��.\�wH����&:��V���p|ɿ��߿[h��8g�=	!�8+�$�*�I6��� �޿S���>���y�L&w�Hŋ��(���_ٿ���b/���)���+���"� f�7� ����˿�ֹ��%��K��*}��fA`�@�>���&�j�����*�q}E���h�1懿6>��@�'����(пq��km�IS�lh%��[,�s�'�����^ �4�οﭣ�4�����t�g,~�%ݔ���������B�!��+��)����b��%���#ڿXſS���S��ǥ��<�y��DT�:t5�7!�������2��nP��ou��y��VW���  �  ���>#������rR2�$�T��.n��v�%1k���N��(�ʚ�N0ƿ���!<���d����ѿ��	�W�0��V��fo��lv�y�i���M�9*�����ֿ4J���[����v�US��|4�GY�7���;���E��g�35�-�(���D�v2f�N���'I��� ÿv<���G�b>���^�)s�A�t�FCc�ORB�b����b���%��ͭ��Ʃ��n�q�>��8`�>�s� Mt�%�a��TB�N5�����o�ǿc����w���>j�4EH��t+�
\�sN�����^����2�����h1�!]O�$�r�����k���&�ѿ��r0&�OJ��Yg���u��(q��Y��c5�%���ؿiҪ�����f�������i���#�ЍJ�s�h��Qv�%p��hX��]6�������L�����/4��O^�`>�E#�M(��� �o������F��h ���:��xZ�2�����"�������IR2���T��.n�Țv��0k�f�N�^(�g��x/ƿ8���0;���c����ѿ��	���0�_V�Pfo��lv�)�i���M��8*����t�ֿ�I���[��G�v�� S��{4�hX�B���9��\C��K�4��(�x�D�q1f������H��A ÿ<���G��a>�i�^�s�)�t�3Cc�ARB�Y����d���%��孙�該�Ln忛q�0>�9`�j�s�QMt�\�a��TB��5�5����ǿ����Xx��%@j��FH�>v+�d]��O�n�������4���yi1��]O���r�����������ѿ���0&��J�Zg�E�u�-)q���Y�5d5�����ؿ[Ӫ�g���?������~j��6�#��J���h��Qv�Op�iX��]6�%�����~L��B���4��`P^��>��#��)�L� �����!����G�8j ��:�'zZ�>���  �  �"���þ�5����0�%:g��a��ȟ�I ��ʍ���ъ���_�)�(�����1�Ŀ�����HͿSQ���4�|[l��
��Gh��s��㚜�����Z�D�%�uc򿄬���$��{nW���/�d��L����jѾ<�ξv�ؾ|)�(P	�Z#"�3D��Lt�R����ӿtY�U�B��Qy������e��W#��#��aU����L������r���ǃ��*�ݿ�}�u�F�B�~�����u��qG��&̖��3��H�p�+hڿ`~��K�z���H��f%�ñ�s�siھϾ�tо�޾K�������J,�iUR�qh�����~�\	 ���T�6S��=͚�M���c����~��s�r�1�:��	�3<ҿ�����C����4V#�m�Y�����������%�����FPm�'�6�E��y:ſ`i��$h��;�=������n3վξ�Ӿ�3�:������7�}Bb�0"��/þ�����0��9g��a��ȟ�, �������ъ�t�_���(�����>�Ŀ�����GͿ�P�	�4��Zl�z
��h��@���������_�Z��%�c�3���:$���mW���/�Ec�?K����hѾ,�ξZ�ؾ_'�O	�X""�2D��Kt�攝�1ӿGY�,�B��Qy�囔��e��L#��	#��ZU����L���������ރ��L�ݿ�}���F�b�~�����u���G��A̖�+4�B�H�Ip��hڿ�~����z�ٺH��g%����u�lھ�	Ͼwо&�޾R������XK,�0VR��h������꿕	 ���T�]S��j͚����������~����r���:���	�4=ҿ���D��S�V#���Y����
������!%�����hPm�L�6�q���:ſ�i��Bh�'�;����<��
�s6վξ��Ӿz6澌��P��і7�xCb��  �  ����ѿ^��|U��.��V��N��I@��/���q���>��D�N��t��r�O�ѿ���k �/o]�~(�������S�������O��8a��fC���|F�6�z���GW�� JL����t�4�۾uþ�-��Hܳ�b���@Ͼxﾠf���5��po����G쿎F*���l�?͙�"<������9������ q��^�|�dr9�'�Adٿ(�ֿ�����2�P�t����_��,'���������x����t��1��+��������w�@ ;�X��1��e!Ҿϓ���<��~e��K!���eؾ{����'�>F�����lw��2��1?��H��ݤ��
��$���M���4��� ��de��M&����$�ҿ���d��NG�ZC������������Q��zF������(]�%>���ٿ "���P`��,�D
�����ɾ�E���v�������Ǿ�㾺���'�NY�����Bѿ7�c|U�o.��C���M��,@�����G���>��؅N�Mt��q�B�ѿj��k ��n]�8(������KS�������O��a��EC���|F��5�!����V��PIL���s���۾�þ�+��Jڳ�Z���>Ͼvﾨe��5��oo�)���F�cF*�{�l�.͙�<������.������q��V�|�`r9�'�Ndٿ?�ֿ�����2�l�t�����/_��A'������!�������$�t�'1�o,��O���3�w�};��������#ҾO���G?���g��w#���gؾX����(��>F�����w��h��U1?��H��/ݤ��
��Z�������u���d���e�qN&����$�ҿ���de�<OG��C��ڡ��֭��"��b���F������(]�K>���ٿ�"���Q`��,��
�w羥�ɾfH��fy�����F�Ǿb�����'��NY��  �  �b��X��3(�bnq��̡�&������O�����{�������i��J'�k���x����:4���z�����0��o"���������e�������_�7��ο�q���@J��D�����ʾ�4���P��x9��â������4޾َ��1�;7r�Q⭿�
�Ƚ>�	F��*�����H@������8�����&b���CQ�+��ا��^�I��
�I��׊�(R���9������ƀ���,���{���ۊ�c�F�����x��[�{���6��.���8f�����4���ƛ��XZ���pǾ���S��uC�������ſ~g�SVW���?ڻ�b���jF��9���H���?���i݁���:������濲j��5\!�Wa�-���%ɿ���������c	��y4���O���az��\/����ڟ�"�`��b&�����վs�������ݤ�����P��]�ѾBr��tn!��X�;b����(�@nq��̡�������2�����Q���Q����i�J'�e���b��@��4�C�z����D0��2"������y���<��z�����_����ο�q��J@J�:D����R�ʾ3���N���7��Ǡ������2޾���1�a6r��᭿T
���>��E���)�����;@��|���8�����"b���CQ�,����_�Z�� �I��׊�8R���9������݀���,���{��܊���F�#��]y����{�
�6��/���⾹h��(���������\���rǾb��2��vC� �G�ſ�g��VW�9��iڻ������F��v������������݁��:�S����濦k���\!�yWa�W���Hɿ�̞������s	���4���O���az��\/�3�J۟��`��c&�N����վ*����"��rा���hS����Ѿ�t��xo!��X��  �  S����~迓~.��{�V��	���YD������K����I��(��%�s���-����%��	��S;�҂��X������F��W������8���u���hi�0��OԿki���\J�������ž�C��F���]���ѧ�͏��Pپ�h�%90�h t�4���oL��{F��+����@w��v���!������ۖ��������Y�'$��h��K��1��9�Q��Ր��$�����4�������+������������N�r������
�}�<6�&
�}�ݾ�J��P8���꠾�q�� M¾���p-�zIC�:�����ʿ����g`������H��^���:���4������Y��ep����B�&��M�O���	�'� �j� ��\,��m���V��9N���V��H���4���yA6��W�hˢ�
b��%�,��-�о����o\��=��S���O��2�̾&������-�Y������~�n~.���{�F������BD��ޚ��'����I�������s�6�-�����$�y�	�/S;��т�vX��[���F���V��ƀ����au���hi�����NԿi��C\J���B�֔ž�A��e���l���ϧ�Ս��aپh�@80��t�Ж��AL��{F��+����1w��i���������Ֆ��������Y�)$��h��c��B��O�Q��Ր��$��'���I�������D�����������Q�N����K���7�}�T=6�c 
���ݾMM���:�� �=�,s��O¾}��Q.�OJC������ʿ���g`������H������q���q����������p���B����$N�E���x�'���j�? ��,��/m��W��IN��W��T���A����A6�X��ˢ��
b�%������о����,_���?���U��ER����̾a�������Y��  �  �b��X��3(�bnq��̡�&������O�����{�������i��J'�k���x����:4���z�����0��o"���������e�������_�7��ο�q���@J��D�����ʾ�4���P��x9��â������4޾َ��1�;7r�Q⭿�
�Ƚ>�	F��*�����H@������8�����&b���CQ�+��ا��^�I��
�I��׊�(R���9������ƀ���,���{���ۊ�c�F�����x��[�{���6��.���8f�����4���ƛ��XZ���pǾ���S��uC�������ſ~g�SVW���?ڻ�b���jF��9���H���?���i݁���:������濲j��5\!�Wa�-���%ɿ���������c	��y4���O���az��\/����ڟ�"�`��b&�����վs�������ݤ�����P��]�ѾBr��tn!��X�;b����(�@nq��̡�������2�����Q���Q����i�J'�e���b��@��4�C�z����D0��2"������y���<��z�����_����ο�q��J@J�:D����R�ʾ3���N���7��Ǡ������2޾���1�a6r��᭿T
���>��E���)�����;@��|���8�����"b���CQ�,����_�Z�� �I��׊�8R���9������݀���,���{��܊���F�#��]y����{�
�6��/���⾹h��(���������\���rǾb��2��vC� �G�ſ�g��VW�9��iڻ������F��v������������݁��:�S����濦k���\!�yWa�W���Hɿ�̞������s	���4���O���az��\/�3�J۟��`��c&�N����վ*����"��rा���hS����Ѿ�t��xo!��X��  �  ����ѿ^��|U��.��V��N��I@��/���q���>��D�N��t��r�O�ѿ���k �/o]�~(�������S�������O��8a��fC���|F�6�z���GW�� JL����t�4�۾uþ�-��Hܳ�b���@Ͼxﾠf���5��po����G쿎F*���l�?͙�"<������9������ q��^�|�dr9�'�Adٿ(�ֿ�����2�P�t����_��,'���������x����t��1��+��������w�@ ;�X��1��e!Ҿϓ���<��~e��K!���eؾ{����'�>F�����lw��2��1?��H��ݤ��
��$���M���4��� ��de��M&����$�ҿ���d��NG�ZC������������Q��zF������(]�%>���ٿ "���P`��,�D
�����ɾ�E���v�������Ǿ�㾺���'�NY�����Bѿ7�c|U�o.��C���M��,@�����G���>��؅N�Mt��q�B�ѿj��k ��n]�8(������KS�������O��a��EC���|F��5�!����V��PIL���s���۾�þ�+��Jڳ�Z���>Ͼvﾨe��5��oo�)���F�cF*�{�l�.͙�<������.������q��V�|�`r9�'�Ndٿ?�ֿ�����2�l�t�����/_��A'������!�������$�t�'1�o,��O���3�w�};��������#ҾO���G?���g��w#���gؾX����(��>F�����w��h��U1?��H��/ݤ��
��Z�������u���d���e�qN&����$�ҿ���de�<OG��C��ڡ��֭��"��b���F������(]�K>���ٿ�"���Q`��,��
�w羥�ɾfH��fy�����F�Ǿb�����'��NY��  �  �"���þ�5����0�%:g��a��ȟ�I ��ʍ���ъ���_�)�(�����1�Ŀ�����HͿSQ���4�|[l��
��Gh��s��㚜�����Z�D�%�uc򿄬���$��{nW���/�d��L����jѾ<�ξv�ؾ|)�(P	�Z#"�3D��Lt�R����ӿtY�U�B��Qy������e��W#��#��aU����L������r���ǃ��*�ݿ�}�u�F�B�~�����u��qG��&̖��3��H�p�+hڿ`~��K�z���H��f%�ñ�s�siھϾ�tо�޾K�������J,�iUR�qh�����~�\	 ���T�6S��=͚�M���c����~��s�r�1�:��	�3<ҿ�����C����4V#�m�Y�����������%�����FPm�'�6�E��y:ſ`i��$h��;�=������n3վξ�Ӿ�3�:������7�}Bb�0"��/þ�����0��9g��a��ȟ�, �������ъ�t�_���(�����>�Ŀ�����GͿ�P�	�4��Zl�z
��h��@���������_�Z��%�c�3���:$���mW���/�Ec�?K����hѾ,�ξZ�ؾ_'�O	�X""�2D��Kt�攝�1ӿGY�,�B��Qy�囔��e��L#��	#��ZU����L���������ރ��L�ݿ�}���F�b�~�����u���G��A̖�+4�B�H�Ip��hڿ�~����z�ٺH��g%����u�lھ�	Ͼwо&�޾R������XK,�0VR��h������꿕	 ���T�]S��j͚����������~����r���:���	�4=ҿ���D��S�V#���Y����
������!%�����hPm�L�6�q���:ſ�i��Bh�'�;����<��
�s6վξ��Ӿz6澌��P��і7�xCb��  �  ���>#������rR2�$�T��.n��v�%1k���N��(�ʚ�N0ƿ���!<���d����ѿ��	�W�0��V��fo��lv�y�i���M�9*�����ֿ4J���[����v�US��|4�GY�7���;���E��g�35�-�(���D�v2f�N���'I��� ÿv<���G�b>���^�)s�A�t�FCc�ORB�b����b���%��ͭ��Ʃ��n�q�>��8`�>�s� Mt�%�a��TB�N5�����o�ǿc����w���>j�4EH��t+�
\�sN�����^����2�����h1�!]O�$�r�����k���&�ѿ��r0&�OJ��Yg���u��(q��Y��c5�%���ؿiҪ�����f�������i���#�ЍJ�s�h��Qv�%p��hX��]6�������L�����/4��O^�`>�E#�M(��� �o������F��h ���:��xZ�2�����"�������IR2���T��.n�Țv��0k�f�N�^(�g��x/ƿ8���0;���c����ѿ��	���0�_V�Pfo��lv�)�i���M��8*����t�ֿ�I���[��G�v�� S��{4�hX�B���9��\C��K�4��(�x�D�q1f������H��A ÿ<���G��a>�i�^�s�)�t�3Cc�ARB�Y����d���%��孙�該�Ln忛q�0>�9`�j�s�QMt�\�a��TB��5�5����ǿ����Xx��%@j��FH�>v+�d]��O�n�������4���yi1��]O���r�����������ѿ���0&��J�Zg�E�u�-)q���Y�5d5�����ؿ[Ӫ�g���?������~j��6�#��J���h��Qv�Op�iX��]6�%�����~L��B���4��`P^��>��#��)�L� �����!����G�8j ��:�'zZ�>���  �  �|��4XÿP�׿O��`
������(�F.,�!�#�ώ�?��g��FI������s��~������1?ɿl��Uz�f�&��r,�I�&��=�]d�����ҿ>v���ʮ�qL��R����l�}	I��]-�
�I�J�$���;��/\�I��n񔿩:�������|ɿ�߿�h��`g�`	!�*8+�=�*�]6����޿[���<����y�&w�&ŋ�k(���_ٿ���:/���)�S�+�`�"��e��� �]��{�˿ֹ�%�����v|���?`�ֶ>�-�&�����v�*�f|E�Гh��凿�=���쬿ܐ���(п��7m�
S�"h%�^[,��'�6��,^ �Q�ο���T����t��*~�gܔ����꿠���!���+���)�����b�R%��#ڿ�WſnR��!S�������y�JCT�~r5�y!�U����m�2�EmP�]nu�2y���V��/|���Wÿ�׿���i`
�W��p�(�.,�ߓ#������￮��}H�������s��}�����N>ɿ����y��&�zr,��&�z=�/d����چҿv��\ʮ�+L�������l��I��\-���%��$���;��.\�wH����&:��V���p|ɿ��߿[h��8g�=	!�8+�$�*�I6��� �޿S���>���y�L&w�Hŋ��(���_ٿ���b/���)���+���"� f�7� ����˿�ֹ��%��K��*}��fA`�@�>���&�j�����*�q}E���h�1懿6>��@�'����(пq��km�IS�lh%��[,�s�'�����^ �4�οﭣ�4�����t�g,~�%ݔ���������B�!��+��)����b��%���#ڿXſS���S��ǥ��<�y��DT�:t5�7!�������2��nP��ou��y��VW���  �  �=�L�?��4�S�H��=L󿄹�߿~�ƿ�����L��%rg��J��A���N��p��x��${�� �̿��� ���+�+����t����)�V��ܿ�������q܆��3a��/G��XB�$S���w��C������pYѿ������\��GN���aH�O���-���>ؿ ��@�����8z[���D���C�n�W�����+��������տ^^�=m�{s�߫��c��8��2�%��Y.Կ���������}��IV��&C���E��R]�k ��,������ɋٿ�����"��Q��L����S�����Ͽ�㲿Q���-ju���Q�h	B��H��8c��Q���=����ÿ�Fݿ���:�iN�[�����q2�;�+�����g˿�ĭ�g揿�/n���M�4�A��/K�,�i�:Ќ��Y��kPȿ���=￟K�إ�\4�`S�����K���.�߿�ƿ����K���pg�ZJ�h�A���N�@�p��w��az��J�̿���s��u+�������@��~��)�%���ܿV��������ۆ��2a�w.G�jWB��"S�F�w��B������Xѿ��>������M￪��
H��i������>ؿ����,�����<z[���D�֨C���W�;���+��򨹿M�տ�^鿥m��s�_��6�����؛�2�֋�/ԿI���[���U}�KV��'C�דE�T]�� ���,������ٿ��M��`����쿶�￙��S��忽�Ͽq䲿 ����ku���Q��
B�H�	:c�7R��2>���ÿGݿ|��Z;��N�ʚ�` ��2�;�Y,���⿪h˿�ŭ�T珿�1n�o�M��A��1K��i�ь��Z��Qȿ)���  �  �M,��Z(���-`	�����;ֿD\¿�����V���b���Ds�E�N�^A1�>��T��[�!�p�6�'8V�>�{�M����O���=��X\ƿ�|ۿn���Wd���'/*�l�+�	!�ŭ�N翶����9����|�xu�燿2����5ѿn��0��U(��A,��$��Z�9t��$�� Ͽ���������4���ˆ��yf���C���)�F�������'��]@��Ob����`�����>ú�̾̿��:��c�S#�v�+�^)�� ���~�ֿ����m���Xv�I.z�����򲿓�ῌ
��.���*�a�*�m; ��f�����@޿FnȿA���B���ߓ��.��,Z�%�9���#�(�����k�.�W�J�$�n��1���P������k����ӿI��a��.�B'��o,���%��F��E��Σƿ�ŝ��u����s�������&���������-\$��M,�wZ(�x��_	����;ֿ�[¿����aV��b���Cs��N�@1����۟���!���6��6V���{�����1O��l=���[ƿ?|ۿ?���Gd���/*�Z�+��!�����M�:���9����|�+u�g懿����<5ѿ������T(��A,���$�\Z�t�-$習 ϿV�������n4���ˆ��yf���C���)�_����Й'�K^@�(Pb�S������<���ú�D�̿]係���c�YS#���+�t^)�\!�P��F�ֿ����Yn��)Zv��/z�@���	�ῼ
�/��*�x�*��; ��f�I����@޿�nȿ���BC��R����/���-Z���9�)�#������ .���J�K�n�`2��vQ������k���ӿƑ��a�/�`B'�p,�O�%�5G��F��Фƿ�Ɲ��v����s����������Z��&���\$��  �  {�v��+m�$:S��K0����t;߿"�������}���X��89�^��_�Y���۰��E��#�Ok$��?�B`��`��S����p��(��Z}��a8�$Z��p�Hv��ug���H�n!����EF��+���8��˩���Nۿ����7�)S[���q�A�u�Df�k%H��.$��[��-Ͽ,ʨ��S���zp���M���/�����p��U���W��{��y���,��J��Ml�y����J��\7ʿ�����0 ��HD�NKc�U�t�Zs��^��;�!G�l��|������O ���c���%�*�(jD��d��ku��nr��L]�3d<��U������ˬ��8ą�2d�uC�u-'��(�ng�f��������	�Ô��6�P�T�y�����m1��l�ٿ�]	��>,���O�R�j���v��nn�8T���.������ο�˥����ۢ�^�ȿ2���Q*��rP��Sl�/�v�V+m��9S��K0�W��;߿���&����}���X��79�.�=^�����&����C��"�j$���?��@`�~`��􉛿�p�����M}��a8�!Z��p�<v�|ug�d�H��m!������E������������/NۿC����7��R[�H�q���u��
f�,%H�k.$��[��-Ͽ�ɨ��S���zp�h�M�y�/�����p��U��XX�����qy��,�&J�UNl�ۼ��K���7ʿ%����0 �;ID��Kc���t�cZs�Q�^���;��G�<��H��������;d��&�g�XjD�6�d�lu��nr��L]�Dd<�
V�'����8����ą�;3d��C��.'��)��h�%��V����	�����6�`�T�y�z����1���ٿ�]	��>,��O���j�j�v�!on��8T�"�.�����ο�̥����ܢ�Y�ȿ���XR*�sP�Tl��  �  &#���
��Y���+d���-��t��E�������x_�Ҟ5����������"ӾZ$ξ��վЂ�
���q�ͷ=��j�����g�ȿ����9��Vp�����ġ�Gԥ�T��ة���bV��� ��\�%����:����Կ7.���=�9�u����U��bI���ٙ������Q�JV��
��M��o�����O�U�*�q�����	�ݾ<оeTϾ�k۾J)����b'��K��7~�q	���4޿(	��K�����ؗ�'���Y��"�����{�-�C�Y�O�ڿ)����ۼ��K��8��P�F˃�'!���i��0���x��9Xv���?�)��pzϿ�5��'!q���A�� �&�s���׾4_ξ��Ѿ"B�Q=��߿���1��Z�Y�����������R(��	^��q���s����������Ŏ�	<i�ʚ1��!���ʿ�ѵ���ƿG�����+�,�b�L)��ZS���"���
��=��\+d���-�)t��袻����w_�ޝ5�ۋ����h��n Ӿ�!ξ,�վ]�����yp�޶=�@�j�H���4�ȿx���9��Vp�����ġ�Cԥ�I��ĩ��abV�z� �Q\�r���:���Կ�-�3�=�ݡu�譓�+��;I��mٙ����d�Q�V�+
濩M��0���N�O��*��p�a���
�ݾlо�TϾ=l۾
*������'��K��8~��	��5޿o	�_�K�����ؗ�W������U����{���C���$�ڿ����Zܼ�GL�09�4P�^˃�7!���i��6���x��CXv���?�B���zϿ(6��	"q���A�� �?'�����׾�aξ8�Ѿ�D⾬?������1��Z���� ������;S(�K
^��q��.t��9������,Ǝ��<i�^�1�W"���ʿ�ҵ���ƿP���.�+���b��)���S���  �  >D��e`��nu���5����Q�$��A�̿��U��W%����2ᾙ^ƾ	���ȅ���깾U7˾�龞��3f.�{�c����8޿�m �.a�Q��4ѳ���������K����ަ�\E���C�y����޿��ӿו��yX)�B�h�����w(���y��D5���׾���K����;�{��&۵�O���TC�-B�2����־�1�����{���j��n�ӾcV�����=���{�q宿XG��B�4�"�x�Lk���Q���k��t���m���ӛ�O�p���/����tտ�ۿ�Y	���<�J��F���8��tY���6��W̶������h��&��|�o���Ãk�OB3����UF�X�;qF�����ᚶ�0)ľD�ݾ6���!��kO�8΋��Ŀ��10J��?��e���`���!���������w0����Y����#����ѿG��R��1R�f;��1���n���D��C`��Ru���5����Q������̿���U��V%����0�V\ƾ����h���,蹾5˾�龧��_e.���c����n8޿�m �1a�V��:ѳ���������@����ަ�?E����C�#���޿��ӿ���X)���h�����J(��~y��5���׾�����J��ř;�L���ڵ��N��9TC��A��1����־�1��2��|��ik��/�ӾVW�������=���{��宿�G����4�r�x�xk���Q���k����������ӛ���p�.�/��Vuտ�ۿAZ	�>�<�%J��4F���8��}Y���6��X̶������h��&�}翿�����k�=C3�����H��;�H������T����+ľ��ݾR��	 !��lO��΋���Ŀ��~0J��?�����a���!����������0��)�Y����Y���ѿj ���2R��;��e��������  �  >�����ѱ��,���G�l��l$���ܿ8G��J$U���w���о�=�������뤾x���NϺ�T�׾�s�z�(��e��9���h��3��~�,�������r���l����X��%ƽ��9���=]����u�����翱�
�X�>����rʬ��e��џ���������J̹��Ñ��S��/�}����L���2@������K�žB|���N���ȥ��׮���¾z徽���9��8��#k��K�	�L�J��(����������	��Y���Ш��)������E��H�, ����b��2U�Y����������6������p`������r�����:�|f��d<��'�m��R.�A���ܾR�������������,��=r̾&����w���M��N���Xӿ�n�D9d�����n���b���Z����/���_���ݣ�z�v���0�F>�5������H`*���m�>W����������������������l��l$�,�ܿ�F��x#U���%u���о�;��E���S餾6���"ͺ�N�׾s���(�0e�M9���h��3��~�3�������w���j����X��ƽ��9��T=]�A���������I�
��>����Bʬ�\e��������������&̹��Ñ�IS��/�+���CL��62@����<��žA|���N��;ɥ�wخ���¾o �R���9�e9���k����	���J��(������į���	����������)��*���i�E�bI��ǒ���(3U�{�����������?������p`������u�����:��f���<���m��S.�?���ܾ[T������������.���t̾Y���y���M�|O��aYӿ�n��9d�����������������+0��<`��ޣ��v���0��>�l������`*�w�m�zW��ף�� ���  �  � ����������6�� �m��W$���ۿW��VtP�F����)Ǿ`,��G��L���� ��ߒ��/�ξ�/��L	$���`�Tk���g�,3����.������$���~~��C���X��͝��q�]�=�����������
��>��g��H��5���v��]���4z�������=���rS����"�� 1��i^;���P��3F�������]o��4��<X����۾�%	��5�"|��׷��	��K����pT�����"���G����Z��\�������)F�(b����6���<�ƚU�,���7���`��/���!z��l>��ѣ��U]����:�j���р��A<i��h)�����ҾQ���gP���ŝ�+B���/����þ+�W���
I�RO��
ҿ�H�߰d��������e�����������A��Q�� w�>	1��I��������]�*�rn�Wş��@�����f ������������Ոm�VW$�>�ۿ�V���sP�c����'Ǿ6*��������������5�ξ.���$��`�#k���g�,3����.������*���}~��9���X������$�]���������u�
���>��g���G�����v��4���z�������=���rS�����"���0��^;�X��� F��������o������X����۾O&	��5��"|�Wط�_�	�	K�:����T�����S���{����Z��������N*F��b������5=��U�N��8���`��6���#z��k>��ϣ��V]����:���������<i��i)����*�Ҿ����R���ǝ��D��2��?�þ<-�f���I��O���
ҿ�H�-�d������������ ����������ZQ���w��	1�9J����%����*��rn��ş��@��@����  �  ����=��!���ED��x�c��Z�/�տ+	��V�O�|��o����/̾|
�������"���ʧ�#����Ӿ�� �F4%��P_�It���8��e,�@�t�9���������%l������\��KZ����T�����1�[���8�{j7��}�����C��ƛ��/���Y�������
����J���&���¸��"�;�D���徢G¾�l���}�������ҫ��U��P��,�ݞ5�Ƭy��������C����������N��a���,���%f���<���A��b>��a
����)鿘���M�K����i���%��^��������>��r2���}���3�f��W,��ãg��d*���w�׾����XL��'ڤ�5��,�Ⱦ���&���H��M��*�̿���][�-���UF��l������`O������t����l��M*�J����޿ƚ��0$���d��������T�������=�����-D��L�c��Z�֟տ�����O����~���-̾M��{���� ��rȧ��|����Ӿ�� ��3%�9P_�t���8��e,�J�t�A���������$l������\��.Z����T�t���0��࿉8�j7���}����eC���������2�������
����J���ԏ��������;�������pG¾�l���}��I���8ӫ�VV��D������5���y�3������C�����쀮�(O������`���Zf���<���A���b>�Gb
���������M�m��� j���%��f��������>��q2���}���3����,��{�g��e*�����׾7���~���N���ܤ����p�Ⱦ���'��H�AN����̿f��?^[�X����F����������O��9���5u��%�l�BN*�����L�޿����0$��d��������T���  �  i7��٭��୦����ΨI�6��]qƿ������P�b�!����O�ܾ��¾�Y���c��O���Z~Ǿv��u���*� V^�=�����ֿ���%XX��?��Xˬ�����U��� ��dS��D5~�!a<�H	�?�׿TͿ�c��'#��_�	��>��������3���e������X�v��4�����dc����}�e�>����;����Ҿ~���I䱾�S����ƳϾӀ�r��[9�Yu�2���f��i�-��n�.��^���]r�����B�������Xkg�Z!)�xt��bϿE]Կj����5���v�wޜ�\����T���S��K���`��F�_��� ���߿yZ��Ơe��;/�������1ʾ��Б��ve�������YپQ- �ۤ�{~J��������p	��{B�����r��»�����������މ���KQ������ɐ˿е���8*J������������B7������ĭ��鹆���I���qƿ|�����P�x�!����,�ܾ��¾3W��Qa������|ǾV�侀��:�*�wU^� �����ֿ���)XX��?��_ˬ�����T��� ��PS��5~��`<��	���׿=SͿ�b�'#���_�O	�����k����3���e�������v�Ԉ4�B���c�� �}� �>���.;��k�Ҿ~���y䱾�S�������ϾŁ�,s�L\9��Yu��������-�b�n�I.�������r��?���v���ƶ���kg��!)�Uu��8Ͽ^Կƫ���5���v��ޜ�k����T���S��K���b��N�_��� ��߿�Z����e��</�����辔ʾ���H����g�����)\پk. ����J�I��4����	��{B�����r��J»����ĵ����)����LQ�C������˿��࿛���*J�ֽ����������  �  8���1Ә�����d[�;�'�������tU��fZ���1�0Y�9��Mxྑ6Ͼ	Yʾk�Ѿ���`-���8j9��Be�����r¿KF�
�2��g�s��q��~T��,���a��� N�r�����'��%��Nο`H�sf6��l�F�������<ў��֓�Ӓ}��I�����޿�v����~�� K�B�&��v����Yپ\3̾9�˾�G׾*]�P
��p#�YF���w��h���׿�����C��x�	���6��ޞ��\��N�q�X><����#�ӿHe��k����߿,��
 H��A}����k�����������l��d8����tɿF���0k��=����^���辫�ӾM�ʾ6ξ:�ݾ�$������-��T�|��H���x��,"��U����fL�������p���)��/+`�`�*�eR��U�Ŀ4���)���@O���n%��*Z�&���������Ә����d[��'��������U���Z��1�'X�����u�4Ͼ�Vʾ��Ѿh��8,���Ki9��Ae�M����q¿>F��2��g�s��q��{T��!���a��� N�-����u��h��SMο�G�f6�fl��������ў�z֓���}���I����H�޿@v��c�~�B K���&�|v���� Zپ�3̾��˾�H׾�]��
�.q#��YF�Y�w�Si��e׿�����C�x�6���6����������q��><������ӿf���k��C�߿x��I H�(B}����t��
���������l��d8�����ɿ�����0k��=����_���A�Ӿ�ʾ�ξ��ݾ9'�� ���-��T��|���H��@y�+-"�n�U�����L��ֆ��7q��>*���+`���*��S��~�ĿV���@���IP��Vo%�+Z�Y�������  �  �m�Ld��3K���)�c-�wLؿ	��`���0w��`S�x�4�����|�S������[���$�� �SN;� �Z����!e�����vx��Q��1���Q�ؒg���l�Ww^���@��}�@0�ل��J���!��r����5Կ��
���0���R�9�h�Pl��1]�0�@��H����(�ȿ'������Z�j�ղH�#�+�����\d���m���K��I�	)�JBE�s}f��+���ɠ��5Ŀ�����y���<�|�Z�DNk���i��V�T�4����ɓڿ�s�������̗��۳�e�lE�w�<��[�<�k�
i�&�T� c5����(W�R?���j��<]��$�^���>��v#������"#�������e/���1���O�O�r��玿gD��	�ҿ¶���%�Q�G�r�a�!�l�]'e�B	L�Z9(���Fȿ�'�����	Y����¿�����#�NmH�U"c�Wm�d��3K�Y�)�6-�Lؿ�������1/w��_S�a�4�v���{�����[��.Y��#��� �#M;��Z�T���d�����Ix��Q��1���Q�Ԓg�w�l�@w^���@��}��/�A�������o�������4Կ)�
���0���R��h�l�p1]��@��H�K����ȿ�&��¬����j���H���+� �����d��Bn���K�@J�~	)��BE�~f�,���ɠ�G6ĿA���2z�5�<�ӐZ��Nk���i�_V���4�����ڿPt��w���͗�6ܳ��迨E���<�%�[�S�k�-
i�4�T�0c5����hW鿧?���j���]��G�^��>�Jx#�p������%�v���J���0���1���O�N�r�u莿�D����ҿ���%���G���a���l��'e��	L��9(����&Gȿ)��� ��Z����¿o��3�#��mH��"c��  �  -�%�u:"����E��3^���Ͽ����^����כ�������l���I��:-����#b��h���2��P��bu�Z����������������Կ5
���.����#�??%��!�i����߿����/���bv�Io�RV���栿>sʿ���ed�4"�5�%����5,�0L��2�H�ȿ�3�����S땿*0��s�`�r?��&�X�����#���;�c�\�B���擿�F��f��z�ƿ�ݿס���M��s�̠%��#��{�����k�Ͽj�������j@p���s�j/������0ڿ�!�@\�8�$�ѥ$����T�
���g�׿I�¿�Ա������Ώ���y�u�T�c�5�G �՟��J�O�*��E���h�n���㙿`����ݺ��wͿ�)濦����0!��&���������]Z���H������m�	~|�L���6v��\W꿼���P���%�8:"�i�����]鿕�Ͽ<������yכ������l�g�I��9-�4���`�g�+�2���P�jau��������\��<�����Կ
���"��z�#�-?%��!�C��.�߿]�� /���av��o��U��"栿�rʿl���d��"���%�Q���+��K������ȿh3��r��'땿	0��H�`�^?��&�+X�7��6�#�'�;�ם\�����擿�F���f���ƿYݿh���*N�t�$�%��#��{�����2�Ͽ1������Ap� �s�
0������Z1ڿ�!�e\�T�$��$����m�
��󿻉׿��¿sձ�s���.Ϗ��y���T��5�� �L���K���*�W�E���h�o��"䙿ն���ݺ�(xͿ*����_��r0!�V&���+�����^[���I������m��|�8���w��'X���Q��  �  vc翛l�W���忶�忰C�Sj�1��<Tؿ9y��/����y��j�a�d^E�
8=�.�I�}cj��f��.��fƿ3vܿ���2U�p迳��Vd���%B�1���Կ�ܻ�^����6��>�[�3�B��=��N��|q�������ţʿf;߿���E����t�[��d��꿺3�Aѿ�"���噿@~��V��U@��*?�K�R�7y����
ﳿ�ο��R�꿂��`<�+j��l���pG�[���ZͿ�Q�� ���sv�QQ���>�A���W�Tw����������t�ҿ���+	�X8�ʴ濤~�1�I.��k鿧V޿�>ɿBr��]s���o���L���=��nC���]�眄�]��Oi���ֿ����T�u��)?����դ�@a�K��xۿ��Ŀ����c䋿Kh�[�H�,=��kF�(�c��툿YC��j����gٿ�b�'l��鿝��_��VC��i���濿Sؿ�x������y����a��\E�o6=���I��aj��e��J-��^eƿ�uܿ4�迿T��o�o��$d�����A��0忟�Կ]ܻ�����6��1�[��B���=�SN�H{q�G���y��0�ʿ�:߿v������bt��濻c���꿆3��@ѿ�"���噿�?~��V��U@�#+?���R��y�?���Oﳿe�οL�Ώ������<翶j心m翲��H��࿜[Ϳ�R��� ��uv��Q��>�`A���W��w��e������Āҿ��g	뿔8����~忙��.�bl�PW޿c?ɿs��+t���o�#�L�B�=�9pC��]������]���i��bֿ��aU�ݩ鿖?�o��_���a뿸K迒yۿ��Ŀ؊��O勿-h�=�H�=��mF��c��D�����jhٿ�  �  nd��ɰ���ѿ� �#�� o���"�N�%�&��a�ˣ���9����z���m����� ����¿t���^ ��&�� �����������M̿��ѩ�蘿�_��m�f�6D�Wx)����[��� ��#7��V�(�{��֐�����ٸ���ÿ�ؿ�A��Ow�@G�8�$��W$��n������׿�U�����r��q�G��G���>ҿ�;�~�u�#��n%�����\�����j�ۿ�ſ�����Z��Ⓙ?�� �Z��<:�^�"��L�����!'���@���b�)@��w떿������bʿ��� �l�&n��&�5�!�.O�����s�ǿ� 2����n���w������Y��=�J��@���y%�ʒ#������V�:�ӿ����*��p��������Ds�mO�=H1�����P��+�U�.�"YK��o�_���2Ϝ��c��]���^ѿ� �����n���"��%����`�$��f��p��F�z��m�������¿7s�J�w^ �Q&��� �������[�俎M̿���Щ��瘿�_����f�+5D�Xw)����7���� ��"7�ĲV��{�=֐����_���}�ÿ��ؿDA��&w�G��$��W$�un������׿�U�����r��q�i��u��(?ҿ�;�-~���#�o%�Ŀ��\�C�����ۿz�ſV���o[���Ⓙ���k�Z�_>:���"�:N�)���"'���@�w�b��@���떿:��5���ʿև�7 ���pn�&���!��O�����U�ǿg 3��m�n���w�^���MZ���=⿎��{���y%���#��H��%W�ӿ�����+�� ���~���uFs�O��I1�>��eR�--��.��ZK�.o������Ϝ��  �  T��>���5ۿ��	�i�+��L��d�,m��b���F�=�!��A���������>������<(˿6���W*���M�qf��l���`�0F��$�^�kпgp�������p�0�M��_0�Y�����><��dc�L` �����$��7@���`�'��������l���X�h���I7�iRV���i��uk��qZ��:�Q,�0�俙������������p����ݿ����6�܇W��vj���j�l0Y�%;�4���~�i����&�����~d�z�C�~�'�K5������������o�t��gc-�TpJ���l�K􊿊᥿�e˿�W���2 �[nB��q^��gl�q�g��1Q���.����ѿg�������츚�U����������B���_���l�~�f�4(P�b�/�$��ۚ࿂����땿^�}�j�X�h�9�Yx��0�Q��B��Ni���\	�.���6�x5U��_y���������ۿ��	�A�+���L���d��m�Yb�f�F���!�A���������=������A'˿���:W*���M�f���l�S�`��F��$�3��jп!p������0�p���M��^0�z�����0:��<a�1_ �����$��6@���`�����S���Rl��MX�=���I7�HRV���i��uk��qZ��:�H,�(�俜�������ʔ���p����ݿ����6��W��vj�&�j��0Y�a;�t��V�����1'��M�F�d�ҐC�ڞ'��6���f������p�y��Rd-�$qJ�a�l����᥿,f˿�W��3 ��nB��q^�\hl���g�2Q�6�.�~���ѿY���x���Ź�����^��6����B���_�%�l���f�[(P���/�O��A������앿��}���X��9��y�(2�PT��u��ll��^	����V�6��6U��`y��  �  �R�����1,��#V*�:R^�Cއ�ш��=����S���^���(W���"��v����0㰿
ǿR� � �-��(c��a��6��zi���{��ʂ�i�R����rd�O|��7���EUR�},��M��A����ܾ!�;'�ʾ*wԾ�꾦�����2�?��?n��@��:u̿�J��B;�ʧo�YΎ�y������u���tz�#E�e���ܿ?��(<��&�ֿI@��1?���t�!��q���ٝ�>���Ku��	A��%��}ӿ����(�t�;D��!�������wL־�5˾�̾YpھH���+��_�(��eM����t���t⿇C��L�#������t���5��伌��i���3�[���˿����=���꿇\��"Q�ں������w���ך�pG���&d���/���d?��p��bb�Md7�B����.��O9Ѿ+Gʾi�Ͼ ��� �,���v3���\�\R������+���U*�R^�/އ����� ���kS��w^��_(W�H�"��u����/ⰿǿ˽ �z�-�N(c��a�����Hi���{���ɂ�,�R�]��d��{��韄��TR��,�M�=@�� �ܾ(�;�ʾuԾ�}꾜����;�?��>n��@���t̿�J��B;���o�IΎ�k������l���tz��"E�a���ܿ?��?<��H�ֿ_@��1?��t�4�����ڝ�Y���Ku��	A�5&��~ӿ����b�t��D�l�!����C��O־O8˾a�̾�rھN�����5�(�EfM�������Vu⿿C�I�L�7#���������6��"���ui�E�3�����˿����"������\�#Q�����"����w���ך��G���&d���/���?���p��'cb��e7����2�&��R<Ѿ+JʾW�Ͼ���L	 �d��x3���\��  �  ����oʿ8���JM������@��K���r3�����bT���Մ�9�F�o2�gI޿;�˿ ��6����T��m��`���W��5��������ˡ������>�QR�Y��󭅿:wG���9���Q�׾�����������֬���m˾����g���1�ji��T���h��#��c�ȓ�����������Ջ�����L�r�H�2����B�ҿ]/п�5���4,��/k������	���-�����Ӳ���e���'k��y*�*��|����Dq��6�̹�s7ﾆ;ξJ2��>���7��!���WԾݬ��F����A�&��س�u� ���7��fz��i����������������~-���=\�XA ��P�̿8�ٿ0`���?�������������w7���O���a��ТT���.�ҿ�ڔ���Z��>(�
0�Γ�?ƾT����T���۴�|�þ��޾zI���#�T�����.oʿ���JM�{����@��3���U3�����8T���Մ�ͧF��1�hH޿-�˿�迨���T�qm�����������Z���dˡ����Y�>�!R��������vG�I��������׾ǘ���������Ϊ���k˾����f���1�@ii��T��kh���#�ɕc��Ǔ��
����������̋�����D�r�D�2����O�ҿt/п6���4,�0k������	���-��1������e��!(k��y*��������Eq�%�6��� :�>ξ�4������9��K���
YԾ����"����A�����س��� ���7��fz�$j��"�����������Ǐ���-��>\��A �&�Q�̿'�ٿ�`���?��������������7���O���a���T�����ҿ_۔���Z��?(�M1�����Aƾ0���W���޴�)�þ��޾�J���#�T��  �  ���cZڿ�!�)h�Ns��ƿ��A��X����B��~�����@�`�?!�y�����޿ğ ��y-�%-q�����~B��'8���������a��"����7W�m�yȿ�����iE���6�Ǿ����y���n��,���=��I�پ���&-���k���$��P�7����BM�������6���o��|����f��zȉ��PI��B��5���z��V�A��l��P��Y���9{��j��C����t��wi��*(?�Z,����t���2��G	��k޾!콾7���â��ȣ��E��,�þ��Q����>�	C��裿��rO��@������	e�����,���B������V�y��4��D���߿m�����X�f���L��?���P���.!���E���ɟ���p���(�&�79���O[��"��r����Ѿ�P���7��@��#.�������;�f�����H�S�"��Zڿ��!�h�>s��
ƿ��A��<����B��T�����Ѯ`��>!�r�����޿4� �8y-��,q�U���;B���7���������^a�� ����7W��l�ȿ.���5iE��o4�WǾ����w���l��0���;��U�پ���?-��k������#��%�7����1M�������6���o��s����f��vȉ��PI�C��5��俋��l�A��l��P��k���N{��&j��]����t���i��j(?��,�Uﯿ��t��2�1I	�en޾�����Ţ�$ˣ��G��-�þj�/��r�>�oC��P���G��O�A��ҁ��8e��3��i�����������y�Z4�4E���߿b��}��Q�X�����*L��Z���d���>!���E���ɟ���p���(�e&俟9���P[�7�"��t����Ѿ�S��Q:�����0��F��^ ξ�h�����,�S��  �  �z��@��$�'�(r��c���c��[��o��������R��}���/j�'�����Q��3�H`4�"z{���q���;���W����s������k1���R`�'��1eͿ�j��}E��R�mq辋¾�A��'䟾9睾����|G��UվƩ��5,���m�i0��"� ���>�]����ׯ�����P1���r��m������v����Q����ߢ�0V�,���I��.���׳����Pp��q��f��T0��I����F�-��۳��6w�2��D��{پ.񸾊U��9���7���z��;�X/㾸�w�>��ۅ��qĿz)�ĲW�~���՛��
���E5��;���`]��G���*��NF;��������o���!�i�a����]^���a��Q����������W���{��`/�>
����+W\�s!����E�̾h����������ƍ���4����Ⱦ��|��NT�(z���� �'�r��c���c��D��S��������R���|��/j��~'�����9�忡��_4��y{�z���-������� ���{s��Ԩ��I1��_R`�����dͿ�j��P|E��Q��o�����@��G⟾I坾�����E��eվ֨��4,���m�0���� �c�>�J����ׯ�����C1���r��d������r����Q������GV�<��1�I��.���׳�&���ep���q�����p0��2I��'�F�q���۳��7w�;2��E�H~پ���W���;��:���|��Ͼ�61㾘�J�>�2܅�rĿ�)��W���������:���{5��y����]�����++���F;�#������p����!���a�����^���a��f����������b���{��`/��
�6��X\�3t!�h�����̾�j����������s���v7��M�ȾE��}��OT��  �  ���cZڿ�!�)h�Ns��ƿ��A��X����B��~�����@�`�?!�y�����޿ğ ��y-�%-q�����~B��'8���������a��"����7W�m�yȿ�����iE���6�Ǿ����y���n��,���=��I�پ���&-���k���$��P�7����BM�������6���o��|����f��zȉ��PI��B��5���z��V�A��l��P��Y���9{��j��C����t��wi��*(?�Z,����t���2��G	��k޾!콾7���â��ȣ��E��,�þ��Q����>�	C��裿��rO��@������	e�����,���B������V�y��4��D���߿m�����X�f���L��?���P���.!���E���ɟ���p���(�&�79���O[��"��r����Ѿ�P���7��@��#.�������;�f�����H�S�"��Zڿ��!�h�>s��
ƿ��A��<����B��T�����Ѯ`��>!�r�����޿4� �8y-��,q�U���;B���7���������^a�� ����7W��l�ȿ.���5iE��o4�WǾ����w���l��0���;��U�پ���?-��k������#��%�7����1M�������6���o��s����f��vȉ��PI�C��5��俋��l�A��l��P��k���N{��&j��]����t���i��j(?��,�Uﯿ��t��2�1I	�en޾�����Ţ�$ˣ��G��-�þj�/��r�>�oC��P���G��O�A��ҁ��8e��3��i�����������y�Z4�4E���߿b��}��Q�X�����*L��Z���d���>!���E���ɟ���p���(�e&俟9���P[�7�"��t����Ѿ�S��Q:�����0��F��^ ξ�h�����,�S��  �  ����oʿ8���JM������@��K���r3�����bT���Մ�9�F�o2�gI޿;�˿ ��6����T��m��`���W��5��������ˡ������>�QR�Y��󭅿:wG���9���Q�׾�����������֬���m˾����g���1�ji��T���h��#��c�ȓ�����������Ջ�����L�r�H�2����B�ҿ]/п�5���4,��/k������	���-�����Ӳ���e���'k��y*�*��|����Dq��6�̹�s7ﾆ;ξJ2��>���7��!���WԾݬ��F����A�&��س�u� ���7��fz��i����������������~-���=\�XA ��P�̿8�ٿ0`���?�������������w7���O���a��ТT���.�ҿ�ڔ���Z��>(�
0�Γ�?ƾT����T���۴�|�þ��޾zI���#�T�����.oʿ���JM�{����@��3���U3�����8T���Մ�ͧF��1�hH޿-�˿�迨���T�qm�����������Z���dˡ����Y�>�!R��������vG�I��������׾ǘ���������Ϊ���k˾����f���1�@ii��T��kh���#�ɕc��Ǔ��
����������̋�����D�r�D�2����O�ҿt/п6���4,�0k������	���-��1������e��!(k��y*��������Eq�%�6��� :�>ξ�4������9��K���
YԾ����"����A�����س��� ���7��fz�$j��"�����������Ǐ���-��>\��A �&�Q�̿'�ٿ�`���?��������������7���O���a���T�����ҿ_۔���Z��?(�M1�����Aƾ0���W���޴�)�þ��޾�J���#�T��  �  �R�����1,��#V*�:R^�Cއ�ш��=����S���^���(W���"��v����0㰿
ǿR� � �-��(c��a��6��zi���{��ʂ�i�R����rd�O|��7���EUR�},��M��A����ܾ!�;'�ʾ*wԾ�꾦�����2�?��?n��@��:u̿�J��B;�ʧo�YΎ�y������u���tz�#E�e���ܿ?��(<��&�ֿI@��1?���t�!��q���ٝ�>���Ku��	A��%��}ӿ����(�t�;D��!�������wL־�5˾�̾YpھH���+��_�(��eM����t���t⿇C��L�#������t���5��伌��i���3�[���˿����=���꿇\��"Q�ں������w���ך�pG���&d���/���d?��p��bb�Md7�B����.��O9Ѿ+Gʾi�Ͼ ��� �,���v3���\�\R������+���U*�R^�/އ����� ���kS��w^��_(W�H�"��u����/ⰿǿ˽ �z�-�N(c��a�����Hi���{���ɂ�,�R�]��d��{��韄��TR��,�M�=@�� �ܾ(�;�ʾuԾ�}꾜����;�?��>n��@���t̿�J��B;���o�IΎ�k������l���tz��"E�a���ܿ?��?<��H�ֿ_@��1?��t�4�����ڝ�Y���Ku��	A�5&��~ӿ����b�t��D�l�!����C��O־O8˾a�̾�rھN�����5�(�EfM�������Vu⿿C�I�L�7#���������6��"���ui�E�3�����˿����"������\�#Q�����"����w���ך��G���&d���/���?���p��'cb��e7����2�&��R<Ѿ+JʾW�Ͼ���L	 �d��x3���\��  �  T��>���5ۿ��	�i�+��L��d�,m��b���F�=�!��A���������>������<(˿6���W*���M�qf��l���`�0F��$�^�kпgp�������p�0�M��_0�Y�����><��dc�L` �����$��7@���`�'��������l���X�h���I7�iRV���i��uk��qZ��:�Q,�0�俙������������p����ݿ����6�܇W��vj���j�l0Y�%;�4���~�i����&�����~d�z�C�~�'�K5������������o�t��gc-�TpJ���l�K􊿊᥿�e˿�W���2 �[nB��q^��gl�q�g��1Q���.����ѿg�������츚�U����������B���_���l�~�f�4(P�b�/�$��ۚ࿂����땿^�}�j�X�h�9�Yx��0�Q��B��Ni���\	�.���6�x5U��_y���������ۿ��	�A�+���L���d��m�Yb�f�F���!�A���������=������A'˿���:W*���M�f���l�S�`��F��$�3��jп!p������0�p���M��^0�z�����0:��<a�1_ �����$��6@���`�����S���Rl��MX�=���I7�HRV���i��uk��qZ��:�H,�(�俜�������ʔ���p����ݿ����6��W��vj�&�j��0Y�a;�t��V�����1'��M�F�d�ҐC�ڞ'��6���f������p�y��Rd-�$qJ�a�l����᥿,f˿�W��3 ��nB��q^�\hl���g�2Q�6�.�~���ѿY���x���Ź�����^��6����B���_�%�l���f�[(P���/�O��A������앿��}���X��9��y�(2�PT��u��ll��^	����V�6��6U��`y��  �  nd��ɰ���ѿ� �#�� o���"�N�%�&��a�ˣ���9����z���m����� ����¿t���^ ��&�� �����������M̿��ѩ�蘿�_��m�f�6D�Wx)����[��� ��#7��V�(�{��֐�����ٸ���ÿ�ؿ�A��Ow�@G�8�$��W$��n������׿�U�����r��q�G��G���>ҿ�;�~�u�#��n%�����\�����j�ۿ�ſ�����Z��Ⓙ?�� �Z��<:�^�"��L�����!'���@���b�)@��w떿������bʿ��� �l�&n��&�5�!�.O�����s�ǿ� 2����n���w������Y��=�J��@���y%�ʒ#������V�:�ӿ����*��p��������Ds�mO�=H1�����P��+�U�.�"YK��o�_���2Ϝ��c��]���^ѿ� �����n���"��%����`�$��f��p��F�z��m�������¿7s�J�w^ �Q&��� �������[�俎M̿���Щ��瘿�_����f�+5D�Xw)����7���� ��"7�ĲV��{�=֐����_���}�ÿ��ؿDA��&w�G��$��W$�un������׿�U�����r��q�i��u��(?ҿ�;�-~���#�o%�Ŀ��\�C�����ۿz�ſV���o[���Ⓙ���k�Z�_>:���"�:N�)���"'���@�w�b��@���떿:��5���ʿև�7 ���pn�&���!��O�����U�ǿg 3��m�n���w�^���MZ���=⿎��{���y%���#��H��%W�ӿ�����+�� ���~���uFs�O��I1�>��eR�--��.��ZK�.o������Ϝ��  �  vc翛l�W���忶�忰C�Sj�1��<Tؿ9y��/����y��j�a�d^E�
8=�.�I�}cj��f��.��fƿ3vܿ���2U�p迳��Vd���%B�1���Կ�ܻ�^����6��>�[�3�B��=��N��|q�������ţʿf;߿���E����t�[��d��꿺3�Aѿ�"���噿@~��V��U@��*?�K�R�7y����
ﳿ�ο��R�꿂��`<�+j��l���pG�[���ZͿ�Q�� ���sv�QQ���>�A���W�Tw����������t�ҿ���+	�X8�ʴ濤~�1�I.��k鿧V޿�>ɿBr��]s���o���L���=��nC���]�眄�]��Oi���ֿ����T�u��)?����դ�@a�K��xۿ��Ŀ����c䋿Kh�[�H�,=��kF�(�c��툿YC��j����gٿ�b�'l��鿝��_��VC��i���濿Sؿ�x������y����a��\E�o6=���I��aj��e��J-��^eƿ�uܿ4�迿T��o�o��$d�����A��0忟�Կ]ܻ�����6��1�[��B���=�SN�H{q�G���y��0�ʿ�:߿v������bt��濻c���꿆3��@ѿ�"���噿�?~��V��U@�#+?���R��y�?���Oﳿe�οL�Ώ������<翶j心m翲��H��࿜[Ϳ�R��� ��uv��Q��>�`A���W��w��e������Āҿ��g	뿔8����~忙��.�bl�PW޿c?ɿs��+t���o�#�L�B�=�9pC��]������]���i��bֿ��aU�ݩ鿖?�o��_���a뿸K迒yۿ��Ŀ؊��O勿-h�=�H�=��mF��c��D�����jhٿ�  �  -�%�u:"����E��3^���Ͽ����^����כ�������l���I��:-����#b��h���2��P��bu�Z����������������Կ5
���.����#�??%��!�i����߿����/���bv�Io�RV���栿>sʿ���ed�4"�5�%����5,�0L��2�H�ȿ�3�����S땿*0��s�`�r?��&�X�����#���;�c�\�B���擿�F��f��z�ƿ�ݿס���M��s�̠%��#��{�����k�Ͽj�������j@p���s�j/������0ڿ�!�@\�8�$�ѥ$����T�
���g�׿I�¿�Ա������Ώ���y�u�T�c�5�G �՟��J�O�*��E���h�n���㙿`����ݺ��wͿ�)濦����0!��&���������]Z���H������m�	~|�L���6v��\W꿼���P���%�8:"�i�����]鿕�Ͽ<������yכ������l�g�I��9-�4���`�g�+�2���P�jau��������\��<�����Կ
���"��z�#�-?%��!�C��.�߿]�� /���av��o��U��"栿�rʿl���d��"���%�Q���+��K������ȿh3��r��'땿	0��H�`�^?��&�+X�7��6�#�'�;�ם\�����擿�F���f���ƿYݿh���*N�t�$�%��#��{�����2�Ͽ1������Ap� �s�
0������Z1ڿ�!�e\�T�$��$����m�
��󿻉׿��¿sձ�s���.Ϗ��y���T��5�� �L���K���*�W�E���h�o��"䙿ն���ݺ�(xͿ*����_��r0!�V&���+�����^[���I������m��|�8���w��'X���Q��  �  �m�Ld��3K���)�c-�wLؿ	��`���0w��`S�x�4�����|�S������[���$�� �SN;� �Z����!e�����vx��Q��1���Q�ؒg���l�Ww^���@��}�@0�ل��J���!��r����5Կ��
���0���R�9�h�Pl��1]�0�@��H����(�ȿ'������Z�j�ղH�#�+�����\d���m���K��I�	)�JBE�s}f��+���ɠ��5Ŀ�����y���<�|�Z�DNk���i��V�T�4����ɓڿ�s�������̗��۳�e�lE�w�<��[�<�k�
i�&�T� c5����(W�R?���j��<]��$�^���>��v#������"#�������e/���1���O�O�r��玿gD��	�ҿ¶���%�Q�G�r�a�!�l�]'e�B	L�Z9(���Fȿ�'�����	Y����¿�����#�NmH�U"c�Wm�d��3K�Y�)�6-�Lؿ�������1/w��_S�a�4�v���{�����[��.Y��#��� �#M;��Z�T���d�����Ix��Q��1���Q�Ԓg�w�l�@w^���@��}��/�A�������o�������4Կ)�
���0���R��h�l�p1]��@��H�K����ȿ�&��¬����j���H���+� �����d��Bn���K�@J�~	)��BE�~f�,���ɠ�G6ĿA���2z�5�<�ӐZ��Nk���i�_V���4�����ڿPt��w���͗�6ܳ��迨E���<�%�[�S�k�-
i�4�T�0c5����hW鿧?���j���]��G�^��>�Jx#�p������%�v���J���0���1���O�N�r�u莿�D����ҿ���%���G���a���l��'e��	L��9(����&Gȿ)��� ��Z����¿o��3�#��mH��"c��  �  8���1Ә�����d[�;�'�������tU��fZ���1�0Y�9��Mxྑ6Ͼ	Yʾk�Ѿ���`-���8j9��Be�����r¿KF�
�2��g�s��q��~T��,���a��� N�r�����'��%��Nο`H�sf6��l�F�������<ў��֓�Ӓ}��I�����޿�v����~�� K�B�&��v����Yپ\3̾9�˾�G׾*]�P
��p#�YF���w��h���׿�����C��x�	���6��ޞ��\��N�q�X><����#�ӿHe��k����߿,��
 H��A}����k�����������l��d8����tɿF���0k��=����^���辫�ӾM�ʾ6ξ:�ݾ�$������-��T�|��H���x��,"��U����fL�������p���)��/+`�`�*�eR��U�Ŀ4���)���@O���n%��*Z�&���������Ә����d[��'��������U���Z��1�'X�����u�4Ͼ�Vʾ��Ѿh��8,���Ki9��Ae�M����q¿>F��2��g�s��q��{T��!���a��� N�-����u��h��SMο�G�f6�fl��������ў�z֓���}���I����H�޿@v��c�~�B K���&�|v���� Zپ�3̾��˾�H׾�]��
�.q#��YF�Y�w�Si��e׿�����C�x�6���6����������q��><������ӿf���k��C�߿x��I H�(B}����t��
���������l��d8�����ɿ�����0k��=����_���A�Ӿ�ʾ�ξ��ݾ9'�� ���-��T��|���H��@y�+-"�n�U�����L��ֆ��7q��>*���+`���*��S��~�ĿV���@���IP��Vo%�+Z�Y�������  �  i7��٭��୦����ΨI�6��]qƿ������P�b�!����O�ܾ��¾�Y���c��O���Z~Ǿv��u���*� V^�=�����ֿ���%XX��?��Xˬ�����U��� ��dS��D5~�!a<�H	�?�׿TͿ�c��'#��_�	��>��������3���e������X�v��4�����dc����}�e�>����;����Ҿ~���I䱾�S����ƳϾӀ�r��[9�Yu�2���f��i�-��n�.��^���]r�����B�������Xkg�Z!)�xt��bϿE]Կj����5���v�wޜ�\����T���S��K���`��F�_��� ���߿yZ��Ơe��;/�������1ʾ��Б��ve�������YپQ- �ۤ�{~J��������p	��{B�����r��»�����������މ���KQ������ɐ˿е���8*J������������B7������ĭ��鹆���I���qƿ|�����P�x�!����,�ܾ��¾3W��Qa������|ǾV�侀��:�*�wU^� �����ֿ���)XX��?��_ˬ�����T��� ��PS��5~��`<��	���׿=SͿ�b�'#���_�O	�����k����3���e�������v�Ԉ4�B���c�� �}� �>���.;��k�Ҿ~���y䱾�S�������ϾŁ�,s�L\9��Yu��������-�b�n�I.�������r��?���v���ƶ���kg��!)�Uu��8Ͽ^Կƫ���5���v��ޜ�k����T���S��K���b��N�_��� ��߿�Z����e��</�����辔ʾ���H����g�����)\پk. ����J�I��4����	��{B�����r��J»����ĵ����)����LQ�C������˿��࿛���*J�ֽ����������  �  ����=��!���ED��x�c��Z�/�տ+	��V�O�|��o����/̾|
�������"���ʧ�#����Ӿ�� �F4%��P_�It���8��e,�@�t�9���������%l������\��KZ����T�����1�[���8�{j7��}�����C��ƛ��/���Y�������
����J���&���¸��"�;�D���徢G¾�l���}�������ҫ��U��P��,�ݞ5�Ƭy��������C����������N��a���,���%f���<���A��b>��a
����)鿘���M�K����i���%��^��������>��r2���}���3�f��W,��ãg��d*���w�׾����XL��'ڤ�5��,�Ⱦ���&���H��M��*�̿���][�-���UF��l������`O������t����l��M*�J����޿ƚ��0$���d��������T�������=�����-D��L�c��Z�֟տ�����O����~���-̾M��{���� ��rȧ��|����Ӿ�� ��3%�9P_�t���8��e,�J�t�A���������$l������\��.Z����T�t���0��࿉8�j7���}����eC���������2�������
����J���ԏ��������;�������pG¾�l���}��I���8ӫ�VV��D������5���y�3������C�����쀮�(O������`���Zf���<���A���b>�Gb
���������M�m��� j���%��f��������>��q2���}���3����,��{�g��e*�����׾7���~���N���ܤ����p�Ⱦ���'��H�AN����̿f��?^[�X����F����������O��9���5u��%�l�BN*�����L�޿����0$��d��������T���  �  $b���}��A�� ���R���+�ƿ�0��S�A�UW�N��pt��dF�����uە������\���zþ7Mc��P����p�ؿ���@�b��������8���4����0���������]AE�Iz���޿�Dӿ����Z*�mk�и��܄���^���_�������r��/���#<�-�羮���q�;�.��j��Ծ�J���"����k���c�������W�Ͼ�� ���(���h�ty��=5����4��!{�;���\G�����������n��+���Ds���0��D��&տ^�ڿ��	�)2>�ԓ���6��G����_��a��T���������j���&���"�����W��F�Tl���IǾ����_��� ���R��lm���7��V�ݾ�'�.�:��؂�]h��{��K��މ�j���{v��E���L���>��?đ�~�[�P]�9��Laѿ�	����J�S��������Ju���a��t}��'��
����R������ƿ�0����A�vV�h��gr��?D��Y��:ٕ������Z���xþ~K��b�;P�ؿ��\�ؿ���N�b��������@���6����0�����o���AE��y�0�޿Dӿ(����Y*�k����������^���_������ur������<�������D�q�Ӑ.�Hj�nԾwJ���"��K��ʟ��򬞾����J�Ͼn� �^�(�o�h��y���5���4�"{�g����G���������$o��b����s���0�GE�j'տ/�ڿ-�	�{2>������6��V����_��a��P���������j���&���c���Y�W��G�<n���KǾٞ�����B��=U���o��7:���ݾ�(�3�:�ق��h�����RK��މ������v��YE��M��=?���đ� �[��]�}��bѿ�
�t����S�׼�����xu���  �  �n�����!�����EXJ���������7��,:A�>���E���̩�\i��b��zW����Ⱦ�f����O�Y4��նҿs��QjY�֘��t���l3��3���߻��ġ�T���m=�Pi	�h�׿=Ϳ���#�,za�kE��^���ء��)s��)����V���hx�p�4�'���Ъ��ko���.�)��ؾ*﷾P���AV���ܚ�
�� 4��1Ծ����m)��f��룿`��-�ޘp�4�y��>�������v������fi�$�)������ο�-Կ���϶6�vix�B������|������Ϩ���`��za��V ��ۿ�!��/�V��:��e����˾?4��x���9��䚜�Z짾iཾR�b���:�>!��p��������B�b���:��_���Q������㭫�٪��%�R��z�v濭A˿���s.��fK�"ч��|������n�����������XJ�Բ�����:7��`9A�]���C�����ɩ�g����?U���쭾�Ⱦ&e�6��?O�)4����ҿt��]jY�����~���t3��4���߻��ġ�8��6m=��h	���׿q
Ϳ��0�#��ya�:E��0��������r������V��Chx�8�4������Ϫ�]ko���.��(��ؾ�O���pV���ܚ�����4��$Ծ��sn)��f�:죿�`�7�-�/�p�`����o��������v��! ���i���)������ο�.Կ��!�6��ix��B��#����|������̨���`��{a�W �8�ۿ"���V��;��g����˾�6��oz��6<��B�����⽾|�m��	�:��!��󥹿�����B�����:������Q��Ҵ��-���&���šR�9{����B˿γ�/�0gK�^ч�}������  �  *ۯ�GI��2ٓ��o�c�3�r/ �����큿k?B��z�V��3�о�c�����V��� ���ļ� �׾�� ��� zN�y_���
ÿz�
�j@��e|��G��;5��P��������*����a�.(�{.����Ŀ�㻿��ۿ9'�@G�����i����������H������d�Z�,!�P��<����j��1��������2Ǿ�β�L����4��/3��_ľ����x	��-�6)c�0^��&<ۿ@=��@T��߇�ԋ��8K����[���Ą���M�cU�e��Of������C��gL"���Z�u�����_���i���ӛ��x����F���.�ʿ$s���
U�2�#�]��z۾�'��c[��Ѐ��� ���d���M;�U񾀻���<�K{�8ԭ�����J-��fh�����M�������r���Җ��u�ZK:�o��!ѿw_����̿G���4��o�	��ۄ��ۯ�'I��ٓ��o�8�3�H/ �����=큿�>B��y�T���о�a��k���S��a��[¼��׾�� �"�}yN�@_���
ÿw�
�j@��e|��G��A5��P�������*��d�a��(��-����Ŀ㻿��ۿ�&��G�Ȅ��<��|���{���!�������&�Z��!�����;���j���1�j��*���2Ǿ�β�|���65���3���_ľ��㾆y	�{-� *c��^���<ۿ�=�3AT��߇����iK���������*ń�j�M��U�C��%g��K�����￶L"� �Z�������f���i���ӛ��x����F���c�ʿos���U��#�
^��|۾*���]��C���d#���f���O;�W񾌼���<�I{��ԭ�����;K-�gh�������������'Ӗ���u��K:��o�#ѿ�`��ǒ̿���p4�o�A	��	����  �  푍����o��3C�)���8߿J�������J�&�5�U'ﾯ�ӾZ�þ4k���{ƾ��ؾR���My��0-��U��4���{�����#��kM���w�����K�����+�e��h7��
�=ѿ���q��������󿆷"�КQ�D�{������܌�-+���4a�*�3�X+�Jʿ����7�k��:=��#��������I;�!��"}��4`˾������h�8�p�e�������ÿ���I�.��_\�x���T���ċ��}��V�4�'�ǝ��!����ʤ�hF��W:˿0?��*2���`�5K��Q��E׊���{��wR���$�����D��� ���jZ���0��=�7���^�۾��Ǿ���K�¾1�Ѿ)�뾢����"��3F�`�x�Ⅱ�P�׿VI�U>���j��9��g{������@Ls��0G������F鳿cx���j����ݿ���S�A���n�����Ǒ�����o��3C�����8߿񝦿L���J�&�	4�%�V�Ӿ��þ�h��(yƾK�ؾ���Dx�0-�U�l4��Y{�����"��kM���w�����K������e�Lh7�ٯ
��ѿm�������
�����&�"�s�Q��{������܌�	+��u4a���3�#+��ʿq�����k�):=��#�_������I;""���}���`˾B��^�����8�6�e�%���;�ÿ����.�I`\�2x���T���ċ�~���V���'���������{ˤ�*G��;˿|?��*2��`�EK��Y��I׊� �{��wR� $����RD��� ��kZ���0��>������۾,�Ǿ������¾��Ѿ}�뾼����"��4F�X�x�^�����׿�I��>�݊j��9���{��9���Ls�N1G����'��o곿�y���k����ݿZ����A��n�+����  �  �R��J��5������Gſ}۠�U����Fe��D���(�����= ��뾱��ф���v�ү.��qK��`m��ċ��맿|�ο@�3��%�:�l�M�$R�/�E���+��2�Wؿ��������È��}���Z}����5};���N���Q�n�D���+����;�9����.����~�x�Y��:��� ��<�=���$7�'U澳$��G5	�\��5�7�!V��Gz�.��ˈ����޿x�
�2�(��B�Q��O�,D>��:!��J ��+ƿY1���q��3����ѿ���7P(��`C�P�Q�O�o�=�� "��H�K�ӿq����z����q���N���1�~���`�>���%�8��aa��t�� &�<ZA�"[a�!!�������|��r��;���2���H���R���K���5�`F����E���5��q�������8t����俫��L_2�J�I�ƖR��J��5��������ſ"۠�񘆿�Ee�#�D���(�y���< ������2��vu���.��pK��_m��ċ�I맿T�ο6�1��%�:�j�M�R��E���+��2��ؿb���Q���j�4ģ���|������|;�j�N�`�Q�)�D�q�+�p��;�䲷��.��v�~��Y���:�i� ��<�A���T7羅U�@%���5	������7��V�MHz��.��G���D�޿��
���(�v�B�^Q�|�O��D>�a;!�YK ��,ƿ&2������*	��ڄ����ѿ���eP(��`C�e�Q�+O�{�=�� "��H���ӿ¦��{���q���N���1����Vb����(�ߐ��c�����&�H[A�\a��!�����}����ￄ��2���H�+�R�'�K�:�5��F���G��7����Ñ�4u��~�����_2���I��  �  %|��e����5D�LwԿ	)����Ed��gN��;�}��Q[�8a;��!�g����b��&��B���b�����ƒ�\�������¿Z?ڿ����q	�e�����!�
�N���7ʿj~��
烿�}d�0�]�:�t�?y��"ѷ�^��*�����dw����Ï濵X̿�����-��N����,r�P4P�h�1��F����r9��Z��/�Z�L�Xn�?#���֗�v�������ɿWf��Q �Q�dE�H�����Y�ZU��'��g�x��_�Qb�8B�������ſ�q��a	�W��s���
����&=ݿ��Ŀ?\��Q:��{���r��?�f��E�$f)�����T����6���&8��W���y�����Ĝ��g�������ѿ ���ւ�k�����%E �cVؿ ���Ȍ��"m���\���i�{������ܟӿ�o��|���{��e�x���C��vԿ�(������c���M��3�}��P[��_;���!������(a���&��B���b�����2ƒ�흡�Ǒ��͗¿2?ڿ{���q	�[������
���7ʿ�}��}惿�|d���]��t��x��wз�����)�n�Ł�#w����Z��XX̿�������~��!���o,r�&4P�T�1��F�����9��Z�/�ΕL��Xn��#��Tח��v��<��(�ɿ�f�/R �bQ��E�������Y�!V�������x�<_�wRb��B��-�����ſr�b	�W��s���
����a=ݿF�Ŀ�\���:���{��Ns����f���E��g)�Q��TV������(8�*�W���y�����3Ŝ�fh������ѿ� �<�,��˝�$���E �YWؿ���Ɍ��$m���\���i�f���뺪���ӿlp��̹��  �  �ѿ+�տnԿQ�ѿ�ѿ`>Կ��տ�Kѿ�?Ŀ?)������y�3BQ�I�7�ˬ0�<�Y�q��N���c����ǿ��ҿ`�տ�ӿKdѿ"ҿ��Կ6vտ��Ͽe9�����Be��Rr���K�~x5��I1�s�?��e_�~ ���џ�J"��Peʿ��ӿ+�տ{!ӿ�Dѿ�cҿ�տ1տ��Ϳ����즿{����j���F�"x3�1l2��C�<f�$K����4���`�̿<�Կ/Nտ��ҿ"<ѿ �ҿ�fտ�uԿ��˿Z��������䈿��c�|B���1�t4�o�H�Z$m�����R������ο�7տ��Կ�AҿvLѿ�Iӿv�տ��ӿ �ɿ�涿a��9����=]���>� 1��>6���M�͂t�wԒ��u���A¿�Jп�տb�Կ��ѿxsѿ��ӿK�տk�ҿǿU��v������!W���:���0���8��"S�],|�.(���|���4ſ��ѿ��տԿ��ѿ��ѿ
>ԿK�տ)Kѿ�?Ŀ�(��i�����y��@Q���7�3�0�n<��Y�����~��c���ǿ�ҿ�տ��ӿdѿ�ҿ�ԿvտX�Ͽ*9������d��hr�~�K�Yw5��H1�2�?��d_����!џ��!���dʿG�ӿ��տ!ӿBDѿzcҿKտ�տU�Ϳ�����즿g����j���F�;x3�`l2�c�C��f�]K��J��������̿��Կ�Nտy�ҿ�<ѿ��ҿegտUvԿ��˿���T����刿�c���B��1��4���H�i%m�����RS����Q�ο�7տ��Կ�Aҿ�LѿJӿ�տ��ӿ��ɿ�綿�a���S?]�[�>��1�k@6�)�M��t�Ւ�Bv��B¿lKпq�տƋԿ �ѿ�sѿ�ӿ�տ�ҿ�ǿ'��V��淀��W�i�:�]�0�h�8��$S��-|��(���}��E5ſ�  �  23��=���>����տ����L���Y_�o�W��AEѿf���+��kh��]��n��g��-����ڿ�E�Ї������@H�$a�,Rп���\�������Y�����w�\�U�V�6��f��)��� ��m�*��AG�L�h��`��T��	���E���ƿ�޿6���et� ��
�ߑ�{2�	:ÿx���. ��u^a�ļ_��6{�ܘ�T���ȥ远��+X��Ŷ�l�����A�ȿZ ��:���Y��m8��Wml�U�J�5�-�Ip����iF��H�Kz3��R�1t�`܊��Q��G꨿����ǦͿ;(迭��o�s��c���7�aa߿��������Ħr���]���e�H��L�����̿��ū���ъ����"1��S�ؿu������Ϡ��鑿����`��[@�bx%�i���E[�H�"�/=��2]����-���2���󭿴=��2�տ���L����#_�/�{V���Dѿ����H*��fih�]�:�n��f��9,��ӰڿiE�v��W��v�H��`��Qпg��'����������2�w���U�t�6��e��(���Ӷ�>�*�t@G�*�h�D`���S�����@E��gƿ��޿����Bt����	�ˑ�^2��9ÿo���0 ���^a��_��6{�9ܘ����������XX�8�������.��Ћȿ� ��ܦ����9���nl���J���-��q����G��I�S{3��R��t��܊�R���꨿�����Ϳ�(�����Ŕ����K8�9b߿����������r���]�O�e��H��������̿��� ����������|1����ؿ�u������3Р��ꑿŤ����`�P]@�z%�$�����\���"��=��3]�M��S.���  �  �܇�!���9~ǿ���������6�/�K�ъR���H�&�0�ѻ�B��4$������������Ǹ�q￦�}7��eL�	kR�&�G���0���X�쿪;���㛿�삿�n_���?���$��k��������`德��O�()��+3�)�P�x�s��ޏ�v�����ֿ@����#���>���O�=&Q��(B��&����ο�����Q��S��ힿ�ɿ\��#�-�?�DP��P�MA��'�5#	���ۿ��������x�DT�396�/��H8����徏��P��<G�`�!���<���[�Ϗ��A����ֹ��翚��wx-�d�E�f
R���M��:������������9f���s��Ȗ��?����6ۿ
�*q-���F��IR��"M��l9�Y!����|\̿����q��8Pk���I��6-�	B��������뾒
�����Q*�|TF�tCg�܇������}ǿ����u��^�6� �K���R���H���0�y��}��]#��0����
��%����Ƹ�z�/�7�3eL��jR���G�r�0�����c;���㛿\삿n_���?��$��j�(�������^征��wN�(��*3�$�P���s�9ޏ����%�ֿ����#���>�߯O�%&Q��(B��&����ο�����Q��j��.ힿ�ɿx�#�S�?�DDP�K�P�CMA��'�u#	��ۿ����Q���,x�gET��:6�����9�%��9����羌��@H�H�!�w�<�Z�[�#��������ֹ�G�Ҽ��x-���E��
R��M�Z:�����������*g���t���������W7ۿd
�nq-��F��IR�#M�m9�!����\̿	��0r��mQk��I�8-��C�x��G������������R*��UF�yDg��  �  ��?��u�⿾b�"�E�i4q��3������k����l��M?�����zڿ�Ѯ�����Xϵ��V�y;���I��ru�>���#b�������@h��~;���^Կ&��={u�@�C�� ��|��龏kо6^¾�˿�K�Ⱦ�ݾ��������2��.]�p'���?������l '���T��r}�1D��ϲ���r���C^��/����vȿ�B��Ԅ���7ÿ����o`*�CY����������V���+�Y�*,�@���e���V����b���6����Q� ���wʾO7��ހ���Jξ�i�~�t��/h?�Jo��H��-tͿ�h
�n\6��c�����}��}���6�y�~O��2 �7��!㹿52��/諿bԿO��H	:�^�g�����k��w[��uu�%�J��9���꿨���WN��tR��W+�U����b�׾�žxZ���~ľuվ���]|�k�'�hM�����B?��&�⿚b���E�B4q�q3������I��8�l�UM?�-���yڿ�Ю�����Oε�zU��:�+�I�{ru�����a��r����@h��~;�����]Կ����zu���C�d� ��{�`�龸iо?\¾zɿ�1�Ⱦ�ݾ��������2��-]�'��I?��.���C '�p�T��r}�$D��Ĳ���r���C^��/����vȿ�B��넥�8ÿ����`*�3CY��������%��q���e�Y�F*,����f��gW����b�+�6�C���� ���Szʾ�9��5���Mξ�k�g�G���h?� o�DI���tͿ�h
��\6�[�c�������������y��O�V3 �>��"乿+3��髿5Կ����	:���g�3����k���[��2uu�D�J�:��������N��*uR��X+�������T�׾�žr]��܁ľ?վ`�}���'��hM��  �  74���������6�sr��>��9��@ׯ�4������� �k��1����{ʿ���=�ӿ;�
��t=��!y��-��3���ƞ�� ���I����
e��3*���� �����v�w�9�z��x��ù˾�t�����z���i���i��-tݾ���!&��rX���T�οֲ��DJ����E��c��sî�Y��S����W��|���뿌����X��\忪 ���P�G`��M�����,��{j��5K����P��Z���ֿ剘�b�_��*�Q�� �ᾁþ�p������������>�Ⱦ�@��m���4�S�n��E�����d$�GQ^�`�������f:�����^̚�����C������ؿ�Q��Ѯƿ)��� +��e�����P��@���O���t����y��*=����M��i숿>NK��k��?����վ�������H���|��\l���LҾ����Ji�d1E��3��-��޳�f�6��rr��>��#��$ׯ����W�����k��1�l���zʿ����%�ӿ��
�at=�g!y�r-����������Ӫ��#����
e��3*�%�񿬑��T�v���9��������˾�r��,���~���c���g��,rݾ���4&��qX������ο����DJ�y��5��U��hî�P��L����W�|���뿙���Y��~�� ���P�W`��_���2��D���j��RK��0�P��Z�p�ֿx�����_�>�*�������
þs��9����
��E���=�ȾhB꾴n���4��n�/F���违$��Q^����������:������̚�H����C�H����ؿ�R����ƿ�)��� +�Me�᪏�k��U���^��������y��*=�(��"N���숿>OK��l�tB��b�վc��������J��t��o��OҾ���Qj�K2E��  �  ܈���ſ����N��׉�T�������h������=٦����y�G����=޿�{˿P���:�kLV�p����:��(����.��~��T���&���V?�h��͵��^}�-�7�.����߾�U�����&A��*Z��X���g��:�;������!��oZ��5������#�x�d�`?��P��{-��G$���Z��,y��ʍt�o3�z��A�ҿ��Ͽ���\-��l��ט��̵�2K���=���µ�n����l��K*�=W�"���4�b���&�4� ���Ѿ�䳾c��⨚�T����]���Z��&�ھS��/�1�K�s��b������+8�*Q|����g����������y:���b����]��� �uB�%_̿y�ٿr����@����|�����o3��Fq��@<��<���f�U�}���Jο�Y��+zK��:��ﾭIƾ ֬�kΞ����mם��Ī���¾�������D��ۈ�W�ſ����N�{׉�C�������h������٦�m��
�G�j���<޿�z˿/��8:��KV�(����:�����w.��O��-������V?�8�b͵�^}�~�7�v���߾T��,
��F?��9X��^���e��F�;����ˮ!��nZ��5��C���#�R�d�O?��A��n-��<$���Z��&y��t�o3�|��N�ҿ��Ͽ?���r-�4�l��ט��̵�GK���=��
õ������l�L*��W꿳���a�b���&�r� �@�Ѿ6糾�e��A��������_���\����ھ-����1��s�Zc��0���+8�nQ|�������N��������:���b��M�]�W� ��C�.`̿p�ٿ���@�B���|��(����3��Tq��L<��G����U�����JοZ��{K��;�d��=Lƾ�ج�)ў�?	��ڝ�yǪ�i�¾�龿��ώD��  �  )����0˿g���V�����ű�mn���Z���v���1��ﶋ�%4P���q�֞ѿ��WC!��a_��œ�	޴�r%��c!��
a��V���҇�JG�ս	�[Y��BG��ʷ7��%
�y5۾έ��d���P���n ��y���Rͬ�WGɾ����	� ���[��<������*���n�2�����B�����v����X�����:����")ٿ�TֿsG��4�Tw�k���ս������2���˟��	w�1�I��g����bd��&��9���f;�E������m��qZ���蠾����[־F�h�1�ɫv��������к?�����bI��:��S���Z���� ��׿���+g�3A'�\k���ҿ5��8��~�H�Ĩ��歪�T��m!���)��������3�^�=�c9Կ徐�<NL����X�ڣ��
G���y���Ε����
<��� ��I������E������0˿E���V������ı�Xn���Z���v���1�������3P�s�p忼�ѿ����B!��`_�Pœ��ݴ�4%��-!���`��.���҇��IG���	�Y���F���7��$
��3۾$�������s����������Zˬ�gEɾ���#� ��[�#<����翫*���n�!�����5�����m����X�����:����/)ٿ�Tֿ�G��4�ow�{���!ս������K���˟�,
w�P1��������dd�5&�H<��xi;AH��;���qo���\���꠾����]־ZG�7�1���v�񄲿���?������I��i����������,�����],g��A'�ul���ҿ.�࿩����H�����3T���!���)�������J�^�\��9ԿH���(OL��	�[�a����I��Q|���ѕ������>��K#��|����}E��  �  ܈���ſ����N��׉�T�������h������=٦����y�G����=޿�{˿P���:�kLV�p����:��(����.��~��T���&���V?�h��͵��^}�-�7�.����߾�U�����&A��*Z��X���g��:�;������!��oZ��5������#�x�d�`?��P��{-��G$���Z��,y��ʍt�o3�z��A�ҿ��Ͽ���\-��l��ט��̵�2K���=���µ�n����l��K*�=W�"���4�b���&�4� ���Ѿ�䳾c��⨚�T����]���Z��&�ھS��/�1�K�s��b������+8�*Q|����g����������y:���b����]��� �uB�%_̿y�ٿr����@����|�����o3��Fq��@<��<���f�U�}���Jο�Y��+zK��:��ﾭIƾ ֬�kΞ����mם��Ī���¾�������D��ۈ�W�ſ����N�{׉�C�������h������٦�m��
�G�j���<޿�z˿/��8:��KV�(����:�����w.��O��-������V?�8�b͵�^}�~�7�v���߾T��,
��F?��9X��^���e��F�;����ˮ!��nZ��5��C���#�R�d�O?��A��n-��<$���Z��&y��t�o3�|��N�ҿ��Ͽ?���r-�4�l��ט��̵�GK���=��
õ������l�L*��W꿳���a�b���&�r� �@�Ѿ6糾�e��A��������_���\����ھ-����1��s�Zc��0���+8�nQ|�������N��������:���b��M�]�W� ��C�.`̿p�ٿ���@�B���|��(����3��Tq��L<��G����U�����JοZ��{K��;�d��=Lƾ�ج�)ў�?	��ڝ�yǪ�i�¾�龿��ώD��  �  74���������6�sr��>��9��@ׯ�4������� �k��1����{ʿ���=�ӿ;�
��t=��!y��-��3���ƞ�� ���I����
e��3*���� �����v�w�9�z��x��ù˾�t�����z���i���i��-tݾ���!&��rX���T�οֲ��DJ����E��c��sî�Y��S����W��|���뿌����X��\忪 ���P�G`��M�����,��{j��5K����P��Z���ֿ剘�b�_��*�Q�� �ᾁþ�p������������>�Ⱦ�@��m���4�S�n��E�����d$�GQ^�`�������f:�����^̚�����C������ؿ�Q��Ѯƿ)��� +��e�����P��@���O���t����y��*=����M��i숿>NK��k��?����վ�������H���|��\l���LҾ����Ji�d1E��3��-��޳�f�6��rr��>��#��$ׯ����W�����k��1�l���zʿ����%�ӿ��
�at=�g!y�r-����������Ӫ��#����
e��3*�%�񿬑��T�v���9��������˾�r��,���~���c���g��,rݾ���4&��qX������ο����DJ�y��5��U��hî�P��L����W�|���뿙���Y��~�� ���P�W`��_���2��D���j��RK��0�P��Z�p�ֿx�����_�>�*�������
þs��9����
��E���=�ȾhB꾴n���4��n�/F���违$��Q^����������:������̚�H����C�H����ؿ�R����ƿ�)��� +�Me�᪏�k��U���^��������y��*=�(��"N���숿>OK��l�tB��b�վc��������J��t��o��OҾ���Qj�K2E��  �  ��?��u�⿾b�"�E�i4q��3������k����l��M?�����zڿ�Ѯ�����Xϵ��V�y;���I��ru�>���#b�������@h��~;���^Կ&��={u�@�C�� ��|��龏kо6^¾�˿�K�Ⱦ�ݾ��������2��.]�p'���?������l '���T��r}�1D��ϲ���r���C^��/����vȿ�B��Ԅ���7ÿ����o`*�CY����������V���+�Y�*,�@���e���V����b���6����Q� ���wʾO7��ހ���Jξ�i�~�t��/h?�Jo��H��-tͿ�h
�n\6��c�����}��}���6�y�~O��2 �7��!㹿52��/諿bԿO��H	:�^�g�����k��w[��uu�%�J��9���꿨���WN��tR��W+�U����b�׾�žxZ���~ľuվ���]|�k�'�hM�����B?��&�⿚b���E�B4q�q3������I��8�l�UM?�-���yڿ�Ю�����Oε�zU��:�+�I�{ru�����a��r����@h��~;�����]Կ����zu���C�d� ��{�`�龸iо?\¾zɿ�1�Ⱦ�ݾ��������2��-]�'��I?��.���C '�p�T��r}�$D��Ĳ���r���C^��/����vȿ�B��넥�8ÿ����`*�3CY��������%��q���e�Y�F*,����f��gW����b�+�6�C���� ���Szʾ�9��5���Mξ�k�g�G���h?� o�DI���tͿ�h
��\6�[�c�������������y��O�V3 �>��"乿+3��髿5Կ����	:���g�3����k���[��2uu�D�J�:��������N��*uR��X+�������T�׾�žr]��܁ľ?վ`�}���'��hM��  �  �܇�!���9~ǿ���������6�/�K�ъR���H�&�0�ѻ�B��4$������������Ǹ�q￦�}7��eL�	kR�&�G���0���X�쿪;���㛿�삿�n_���?���$��k��������`德��O�()��+3�)�P�x�s��ޏ�v�����ֿ@����#���>���O�=&Q��(B��&����ο�����Q��S��ힿ�ɿ\��#�-�?�DP��P�MA��'�5#	���ۿ��������x�DT�396�/��H8����徏��P��<G�`�!���<���[�Ϗ��A����ֹ��翚��wx-�d�E�f
R���M��:������������9f���s��Ȗ��?����6ۿ
�*q-���F��IR��"M��l9�Y!����|\̿����q��8Pk���I��6-�	B��������뾒
�����Q*�|TF�tCg�܇������}ǿ����u��^�6� �K���R���H���0�y��}��]#��0����
��%����Ƹ�z�/�7�3eL��jR���G�r�0�����c;���㛿\삿n_���?��$��j�(�������^征��wN�(��*3�$�P���s�9ޏ����%�ֿ����#���>�߯O�%&Q��(B��&����ο�����Q��j��.ힿ�ɿx�#�S�?�DDP�K�P�CMA��'�u#	��ۿ����Q���,x�gET��:6�����9�%��9����羌��@H�H�!�w�<�Z�[�#��������ֹ�G�Ҽ��x-���E��
R��M�Z:�����������*g���t���������W7ۿd
�nq-��F��IR�#M�m9�!����\̿	��0r��mQk��I�8-��C�x��G������������R*��UF�yDg��  �  23��=���>����տ����L���Y_�o�W��AEѿf���+��kh��]��n��g��-����ڿ�E�Ї������@H�$a�,Rп���\�������Y�����w�\�U�V�6��f��)��� ��m�*��AG�L�h��`��T��	���E���ƿ�޿6���et� ��
�ߑ�{2�	:ÿx���. ��u^a�ļ_��6{�ܘ�T���ȥ远��+X��Ŷ�l�����A�ȿZ ��:���Y��m8��Wml�U�J�5�-�Ip����iF��H�Kz3��R�1t�`܊��Q��G꨿����ǦͿ;(迭��o�s��c���7�aa߿��������Ħr���]���e�H��L�����̿��ū���ъ����"1��S�ؿu������Ϡ��鑿����`��[@�bx%�i���E[�H�"�/=��2]����-���2���󭿴=��2�տ���L����#_�/�{V���Dѿ����H*��fih�]�:�n��f��9,��ӰڿiE�v��W��v�H��`��Qпg��'����������2�w���U�t�6��e��(���Ӷ�>�*�t@G�*�h�D`���S�����@E��gƿ��޿����Bt����	�ˑ�^2��9ÿo���0 ���^a��_��6{�9ܘ����������XX�8�������.��Ћȿ� ��ܦ����9���nl���J���-��q����G��I�S{3��R��t��܊�R���꨿�����Ϳ�(�����Ŕ����K8�9b߿����������r���]�O�e��H��������̿��� ����������|1����ؿ�u������3Р��ꑿŤ����`�P]@�z%�$�����\���"��=��3]�M��S.���  �  �ѿ+�տnԿQ�ѿ�ѿ`>Կ��տ�Kѿ�?Ŀ?)������y�3BQ�I�7�ˬ0�<�Y�q��N���c����ǿ��ҿ`�տ�ӿKdѿ"ҿ��Կ6vտ��Ͽe9�����Be��Rr���K�~x5��I1�s�?��e_�~ ���џ�J"��Peʿ��ӿ+�տ{!ӿ�Dѿ�cҿ�տ1տ��Ϳ����즿{����j���F�"x3�1l2��C�<f�$K����4���`�̿<�Կ/Nտ��ҿ"<ѿ �ҿ�fտ�uԿ��˿Z��������䈿��c�|B���1�t4�o�H�Z$m�����R������ο�7տ��Կ�AҿvLѿ�Iӿv�տ��ӿ �ɿ�涿a��9����=]���>� 1��>6���M�͂t�wԒ��u���A¿�Jп�տb�Կ��ѿxsѿ��ӿK�տk�ҿǿU��v������!W���:���0���8��"S�],|�.(���|���4ſ��ѿ��տԿ��ѿ��ѿ
>ԿK�տ)Kѿ�?Ŀ�(��i�����y��@Q���7�3�0�n<��Y�����~��c���ǿ�ҿ�տ��ӿdѿ�ҿ�ԿvտX�Ͽ*9������d��hr�~�K�Yw5��H1�2�?��d_����!џ��!���dʿG�ӿ��տ!ӿBDѿzcҿKտ�տU�Ϳ�����즿g����j���F�;x3�`l2�c�C��f�]K��J��������̿��Կ�Nտy�ҿ�<ѿ��ҿegտUvԿ��˿���T����刿�c���B��1��4���H�i%m�����RS����Q�ο�7տ��Կ�Aҿ�LѿJӿ�տ��ӿ��ɿ�綿�a���S?]�[�>��1�k@6�)�M��t�Ւ�Bv��B¿lKпq�տƋԿ �ѿ�sѿ�ӿ�տ�ҿ�ǿ'��V��淀��W�i�:�]�0�h�8��$S��-|��(���}��E5ſ�  �  %|��e����5D�LwԿ	)����Ed��gN��;�}��Q[�8a;��!�g����b��&��B���b�����ƒ�\�������¿Z?ڿ����q	�e�����!�
�N���7ʿj~��
烿�}d�0�]�:�t�?y��"ѷ�^��*�����dw����Ï濵X̿�����-��N����,r�P4P�h�1��F����r9��Z��/�Z�L�Xn�?#���֗�v�������ɿWf��Q �Q�dE�H�����Y�ZU��'��g�x��_�Qb�8B�������ſ�q��a	�W��s���
����&=ݿ��Ŀ?\��Q:��{���r��?�f��E�$f)�����T����6���&8��W���y�����Ĝ��g�������ѿ ���ւ�k�����%E �cVؿ ���Ȍ��"m���\���i�{������ܟӿ�o��|���{��e�x���C��vԿ�(������c���M��3�}��P[��_;���!������(a���&��B���b�����2ƒ�흡�Ǒ��͗¿2?ڿ{���q	�[������
���7ʿ�}��}惿�|d���]��t��x��wз�����)�n�Ł�#w����Z��XX̿�������~��!���o,r�&4P�T�1��F�����9��Z�/�ΕL��Xn��#��Tח��v��<��(�ɿ�f�/R �bQ��E�������Y�!V�������x�<_�wRb��B��-�����ſr�b	�W��s���
����a=ݿF�Ŀ�\���:���{��Ns����f���E��g)�Q��TV������(8�*�W���y�����3Ŝ�fh������ѿ� �<�,��˝�$���E �YWؿ���Ɍ��$m���\���i�f���뺪���ӿlp��̹��  �  �R��J��5������Gſ}۠�U����Fe��D���(�����= ��뾱��ф���v�ү.��qK��`m��ċ��맿|�ο@�3��%�:�l�M�$R�/�E���+��2�Wؿ��������È��}���Z}����5};���N���Q�n�D���+����;�9����.����~�x�Y��:��� ��<�=���$7�'U澳$��G5	�\��5�7�!V��Gz�.��ˈ����޿x�
�2�(��B�Q��O�,D>��:!��J ��+ƿY1���q��3����ѿ���7P(��`C�P�Q�O�o�=�� "��H�K�ӿq����z����q���N���1�~���`�>���%�8��aa��t�� &�<ZA�"[a�!!�������|��r��;���2���H���R���K���5�`F����E���5��q�������8t����俫��L_2�J�I�ƖR��J��5��������ſ"۠�񘆿�Ee�#�D���(�y���< ������2��vu���.��pK��_m��ċ�I맿T�ο6�1��%�:�j�M�R��E���+��2��ؿb���Q���j�4ģ���|������|;�j�N�`�Q�)�D�q�+�p��;�䲷��.��v�~��Y���:�i� ��<�A���T7羅U�@%���5	������7��V�MHz��.��G���D�޿��
���(�v�B�^Q�|�O��D>�a;!�YK ��,ƿ&2������*	��ڄ����ѿ���eP(��`C�e�Q�+O�{�=�� "��H���ӿ¦��{���q���N���1����Vb����(�ߐ��c�����&�H[A�\a��!�����}����ￄ��2���H�+�R�'�K�:�5��F���G��7����Ñ�4u��~�����_2���I��  �  푍����o��3C�)���8߿J�������J�&�5�U'ﾯ�ӾZ�þ4k���{ƾ��ؾR���My��0-��U��4���{�����#��kM���w�����K�����+�e��h7��
�=ѿ���q��������󿆷"�КQ�D�{������܌�-+���4a�*�3�X+�Jʿ����7�k��:=��#��������I;�!��"}��4`˾������h�8�p�e�������ÿ���I�.��_\�x���T���ċ��}��V�4�'�ǝ��!����ʤ�hF��W:˿0?��*2���`�5K��Q��E׊���{��wR���$�����D��� ���jZ���0��=�7���^�۾��Ǿ���K�¾1�Ѿ)�뾢����"��3F�`�x�Ⅱ�P�׿VI�U>���j��9��g{������@Ls��0G������F鳿cx���j����ݿ���S�A���n�����Ǒ�����o��3C�����8߿񝦿L���J�&�	4�%�V�Ӿ��þ�h��(yƾK�ؾ���Dx�0-�U�l4��Y{�����"��kM���w�����K������e�Lh7�ٯ
��ѿm�������
�����&�"�s�Q��{������܌�	+��u4a���3�#+��ʿq�����k�):=��#�_������I;""���}���`˾B��^�����8�6�e�%���;�ÿ����.�I`\�2x���T���ċ�~���V���'���������{ˤ�*G��;˿|?��*2��`�EK��Y��I׊� �{��wR� $����RD��� ��kZ���0��>������۾,�Ǿ������¾��Ѿ}�뾼����"��4F�X�x�^�����׿�I��>�݊j��9���{��9���Ls�N1G����'��o곿�y���k����ݿZ����A��n�+����  �  *ۯ�GI��2ٓ��o�c�3�r/ �����큿k?B��z�V��3�о�c�����V��� ���ļ� �׾�� ��� zN�y_���
ÿz�
�j@��e|��G��;5��P��������*����a�.(�{.����Ŀ�㻿��ۿ9'�@G�����i����������H������d�Z�,!�P��<����j��1��������2Ǿ�β�L����4��/3��_ľ����x	��-�6)c�0^��&<ۿ@=��@T��߇�ԋ��8K����[���Ą���M�cU�e��Of������C��gL"���Z�u�����_���i���ӛ��x����F���.�ʿ$s���
U�2�#�]��z۾�'��c[��Ѐ��� ���d���M;�U񾀻���<�K{�8ԭ�����J-��fh�����M�������r���Җ��u�ZK:�o��!ѿw_����̿G���4��o�	��ۄ��ۯ�'I��ٓ��o�8�3�H/ �����=큿�>B��y�T���о�a��k���S��a��[¼��׾�� �"�}yN�@_���
ÿw�
�j@��e|��G��A5��P�������*��d�a��(��-����Ŀ㻿��ۿ�&��G�Ȅ��<��|���{���!�������&�Z��!�����;���j���1�j��*���2Ǿ�β�|���65���3���_ľ��㾆y	�{-� *c��^���<ۿ�=�3AT��߇����iK���������*ń�j�M��U�C��%g��K�����￶L"� �Z�������f���i���ӛ��x����F���c�ʿos���U��#�
^��|۾*���]��C���d#���f���O;�W񾌼���<�I{��ԭ�����;K-�gh�������������'Ӗ���u��K:��o�#ѿ�`��ǒ̿���p4�o�A	��	����  �  �n�����!�����EXJ���������7��,:A�>���E���̩�\i��b��zW����Ⱦ�f����O�Y4��նҿs��QjY�֘��t���l3��3���߻��ġ�T���m=�Pi	�h�׿=Ϳ���#�,za�kE��^���ء��)s��)����V���hx�p�4�'���Ъ��ko���.�)��ؾ*﷾P���AV���ܚ�
�� 4��1Ծ����m)��f��룿`��-�ޘp�4�y��>�������v������fi�$�)������ο�-Կ���϶6�vix�B������|������Ϩ���`��za��V ��ۿ�!��/�V��:��e����˾?4��x���9��䚜�Z짾iཾR�b���:�>!��p��������B�b���:��_���Q������㭫�٪��%�R��z�v濭A˿���s.��fK�"ч��|������n�����������XJ�Բ�����:7��`9A�]���C�����ɩ�g����?U���쭾�Ⱦ&e�6��?O�)4����ҿt��]jY�����~���t3��4���߻��ġ�8��6m=��h	���׿q
Ϳ��0�#��ya�:E��0��������r������V��Chx�8�4������Ϫ�]ko���.��(��ؾ�O���pV���ܚ�����4��$Ծ��sn)��f�:죿�`�7�-�/�p�`����o��������v��! ���i���)������ο�.Կ��!�6��ix��B��#����|������̨���`��{a�W �8�ۿ"���V��;��g����˾�6��oz��6<��B�����⽾|�m��	�:��!��󥹿�����B�����:������Q��Ҵ��-���&���šR�9{����B˿γ�/�0gK�^ч�}������  �  mv��'&������bh���-�m��.���_m�*�+������;-������B���\ˉ�j`��W���*��A�׾n	��7�,��g�������::�2�u�wo��v���	��E����:���[�7�"�ؖ�W㾿'��Hտ���6A���{�-ݗ��*����ۯ���\���zT��=�+�ؿ����,T�������+���T壾���㊾z��[����~��XǼ���D����L��:��пgh���M��K��.���P����*��{A����o�G����i�ڿۉ����7�e�׍T��:�����7����+��j����{�k�@��/
�����)E���n>����;�ܾ��������[���쉾T���nܕ�p ���0ɾ@���&�r�d�6����S��L'���a��D��{���^��䤥�᷒���n�}�4�GC�s�ʿ�����?ƿ�����.�;9h������!��Fv��&�����|bh���-����~���^m�e�+�̥���;-����}�����(ɉ�@^��F���(����׾Om	���7��+��X�������::�I�u��o��������?����:��b[���"�+�ￖ⾿Y��tտ���H6A�Z�{��ܗ��*��¡�������\��TzT�L=���ؿ���O,T�#����ɴ��#壾��䊾_z��餑�z��Hȼ�����W�L��:���п�h�,�M��K��]��������*���A��>���G�	��N�ڿ�������7�ee��T�
;�����:����+��e����{�i�@��/
����eE��.o>�i�� ݾȅ������]���� ���ޕ��"���2ɾK���&�m�d�����NT�M'�=�a�E��M{���^��'���*���N�n��4��C���ʿʛ���@ƿ/����.��9h������!���  �  >��d��w����^�'�&����k��Lj��y+����#�Ѿ��|�������\����<���)��GC���K۾^v
�]+7�)]|�?���/ ���2�ik�� ��aϟ��£��Ǚ��d���R�j��a}�RT������xMοf��$s9��*q��i������L���ٗ�����D�K�j��<ҿ����@R�������Ͱľ����3▾v���!A��&���N���0�����뾭=���J�[r��F�ɿ����eE��I}�kӕ�����
��s����:w�]�?��K���ӿ�\�������࿭i���K�ˇ��y��DS��?���e��qAq�6�8�wF��l��4���t=�Ѓ�k��З���+���<��S���-Ώ��ؙ�n=���;V����	&���a�$������ �!QX�_4��[{��X��������]�d��-�"���Ŀ����N��������'�T�^����w ����E��^��ɝ^� �&���쿹j��YKj��x+����B�Ѿ��Y����!����:���'��VA��)J۾�u
��*7��\|�-���/ ���2�k���jϟ��£��Ǚ��d��VR�"���|翓S�������Lο����r9�/*q�|i�������L���ٗ������K��i�|<ҿu��J@R������l�ľe���3▾����A��������� �����Z>���J��r����ɿ��fE�@J}��ӕ�����>������V;w�τ?�cL���ӿ�]��ˊ������i�	�K�⇁����IS��=���e��jAq�6�8��F��l��s��2u=����P��癹��-��6?�������Џ��ڙ��?���;a����
&���a������� �qQX��4���{�����Y��������d���-�S#�� �Ŀꕯ�DO������{�'�͗^���� ���  �  �����]r��MD�&����׿�@����c���,�x���޾Ҽ��,g������T��{t���C����þ�,辤���7��Ys��㦿�1�N���O���z�� ��]���-�����h��y9����]ѿ`���zݢ��㻿w���QH$�PT�,e��9���1���,��`�c��4����;��{�����N�����u��RIҾ\u��y�����������������tξ���*��uH�!ˆ��?���\��.���^�ui��&������������Y��~)����������������Gg˿��U4��c�T���A������FMT�?#$�����h�{�;�<�Z���%�LLǾ�^��l���:z��/͛�����Pպ�wھ
����'�4p\��˕�}пʱ��>��rm��W��sԏ��"��q�v�}�I�Q�a��(���a����wm޿=,�9BD��Pr���������*r��MD������׿n@���c�2�,�����޾�����d��Ɠ��]R��0r���A����þ�*����7�(Ys��㦿�1�W���O���z�� ��_���&�����h��y9����j\ѿ�����ܢ��⻿�����G$��OT��d�p9���1���,���c�N4�g�;��-����N����6u���HҾ-u��y��ܐ����5��?����uξ:���֌��uH��ˆ�|@��]�\�.��^��i��W���%��-����Y��~)�����i������S����g˿���4�G�c�T���A������CMT�B#$�&�������{��<�9���'�}NǾ�`��Ҍ���|���ϛ������׺�Ayھ����'�*q\�6̕��п��c�>��rm��W���ԏ�2#����v��I������^�������B����n޿�,��BD�!Qr�����  �  ��g�37^�#VD��J!�z���8����x���a��q4�������yؾ����,���ᜮ��Ҵ�ž�(߾#��|��|=��Hm��I���4ʿ��>o)�,K���a��dg�U�Y�b�<�A����迯���6I��g���<!����Ϳ�@�ք,�$AN�O�c���f�hW�A9�����N�����9aP�/�(�H�K��cϾ�̺�����������N�̾*꾷t	�%��AK��р��ܧ���ݿp���b5��]T�T�e���d��`Q�ݜ0��G��?Կ�Х�����1p��������~�T�8�dW�z�f�#|c��cN�+w-��	�לпL�����s���A��&��b����lǾq ��ˮ�?���`���Pվ�f��}��7`0��?[��Q���&��dd��3�m�@��	\�`�g�FH`��G��5$�.���z7¿d���,Ӎ�t嘿����0��� �:�C�,M^�F�g��6^��UD��J!�(��������x���a��p4�&�������vؾQ�����k���wд� ž�&߾!������=�_Hm��I���4ʿ��Go)�',K���a��dg�D�Y�?�<���������H������y ���Ϳ]@�x�,��@N���c�o�f�W��@9���j���������`P�ϯ(���cϾ�̺�������s��
�̾�*�Fu	��%��BK�hҀ�ݧ�/�ݿ���c5��]T���e���d�KaQ�H�0�H�[@Կtѥ������p��d��G��I~���8��W���f�)|c��cN�/w-�	���п������s�ΚA��'��c���⾕nǾ�"���ͮ�����ʆ��hRվ�h�����0a0��@[��Q��'���d�64�½@�V
\�Ϲg��H`�j�G�6$�R����8¿����Nԍ��昿¼��1��Y ���C��M^��  �  em-��G'��.������п�Щ��U����l���J�2�.�������p��3�ԾE�Ͼ��׾mK�������4�`�Q�9�u�'$��ʞ��t[ڿ��������)���,�c#�*O��������͑��cx�Hsp���"���jҿ������!*�5�,�
�"�2��-��U�¿�����Q��	�`���@�oi&�-��������߾�Ѿ��о#�ݾ���av�.�#�I�=�(�\�с�Ý���5�����^��� �JH,��+�P����n�׿=d��㯈��q���u��������M(����&!��,��*����(4�:_߿>����1���z��ZU�q�7��m��	�\d�r�پ��Ͼ%�Ӿ6���� ��p�G�+��{G�+�h�����4����˿�Q�������%��c-���'���o���ǿd���w���o��~��嘿���y�������L&�m-��G'�p.�������п�Щ�6U����l���J�=�.��������}羛�Ծ��Ͼ:�׾�H�s��l���4���Q���u��#������e[ڿ��������)���,�N#�O�?�近���_͑�Tbx��qp�I��i����ҿ��A��=!*���,�Ŕ"��������¿e����Q����`�c�@�+i&� ��Յ����߾L�Ѿ>�о��ݾt���v���#���=���\�{с�=����6�����I_��� ��H,��+���2��?�׿e��������q��u�W��������(�0���&!�1�,���*����34�^_߿t����1���z��[U���7�o�	�g�(�پ5�ϾƢӾ����� ��q�N�+��|G��h�󒉿���P�˿;R����R�%�!d-��'�0�v���! ǿz����x���o�&�~��昿����N�������L&��  �  ~9��<����ס̿���Ť�F���.�� Uz��d^�/oA� m&����h��1��+K�����,���G���d�����ƌ��z��td���V��;�ѿ���|���.!�����[�Ϳz<���U��#g�jJ�v�D�ydW��/��~������ݿ��e���D￮�ۿA	ſDE�������L��_ׅ�Bq�]�T�]8��q�\)�H� � �;�	������4�q~Q�W,n��m���萿����7����¿Jbٿ����R�����f�¿n��!����Z�&�E��OH���b��%��U����ɿK1�I���������^QԿ�����G��h����&��쐁�T�g��K�C�.��+����X���%����z�#�)E>�_-[��Uw�A���H��������Kʿ���_g�Gy���&�x�׿�����h��u��5Q�(�C���N��op�f��������VԿ�*��8�����㿁�̿�����Ĥ�틖����<Tz��c^�nA��k&�/�� ��.���I�J��k,�F�G�z�d�+��qƌ�4z��<d��~V��&�ѿ���j���!��\���Ϳ<��mU��
g�4J�+�D�"cW�;/��`}��u��9�ݿ���{d��TD�9�ۿ�ſ�D��g����L��(ׅ��Aq��T�38��q�^)�`� �; ���	�)��W�4��~Q��,n��m��+鐿^��8���¿�bٿ���R��
��n��+�¿5�����@�Z���E��PH��b�L&�����+�ɿ�1�;I��������鿇QԿس���G������'��u�����g�I
K�� /�e-���>����������#�LF>�h.[��Vw��������{������ʿH��h�z���'�[�׿�����i��ńu��7Q�$�C�o�N��qp�A���{³�6WԿq+��  �  v;������L�������ô��d��\�ղ�觿Ԝ���́���Z�`$9��$����[|'�ϥ?��Hc�=���`㚿{��K��M��� ��͐���������-��������i���I����|�xYT��4���!�rk��*���D���i�r���󝿣 ���+��
��b����{���8���߶�L<����������᏿�}u��TN�Ȏ0�H? ��^��.�wJ���p������࠿�ۮ�pݵ������g���u��)���q��֦���B���ꟿ�h���n�m�H���,�P �O� �9�1�{NP���w�A��E���V����d���ζ��"��􀴿�̵�]��洿YV�����䈿Լg��C��{)��1���"�`6��gV���~��g��C������=ö�s����崿������g������F7���ՙ��Y���a�`�=�{�&�=����$���:��\�J���{�������:������PL��6���>ô��d��Aղ��秿K���X́�k�Z��"9�s$�J���z'�7�?�CGc������⚿��cK������ ���������������������si��tI���|��XT��4�x�!�<j���*���D�T�i����^� ��T+���������e{���8��S߶�<��p���񾢿�᏿�}u��TN�̎0�a? ��^�<.�fwJ���p����ᠿ#ܮ��ݵ�����h��v��������~���_C���럿�i��|�n��H�D�,����� �i�1��OP���w�������������d���ζ��"��<���S͵�����洿�V��L򜿍刿d�g��C�f})�=3��"��6�iV��~�h���C��e����ö�Ӓ���崿+�������������8���֙�eZ��la�:�=�W�&�����$�E�:���\����"��������  �  񵊿�E�� ����᷿��Ϳ�5俲`��_��n�-�ҿ1౿fH����m�xUM���C�˧R�H%x��(���g���7ٿ��]�������߿��ȿ�s���.��h������I�u��Y�c�<��Z"�W��$�������G��U��z0�¦L�f�i��I��׎�����>��i澿��տf��;���������,ȿ����I���_�`�ׇG��/F���\�ӌ��z�M�ĿZ,����&���Z��U ؿHS��56���K���7��l�����l�"�O��w3����������3� �����R�9��WV���r��������.���Q���Iƿ�ݿZ�H|��]��Sܿ�%��X�����}���U��bD��K��Ji�����X��v>Ͽe���y���~��p濴yп-,��]w��$���.��~�~��-c��6F�/�*�<��ٮ����r������'��C�G�_���{�|���.E��ɧ��M᷿=�ͿT5�X`������쿝�ҿ�߱��G��@�m��SM�6�C��R��#x��'���f���6ٿ��Ȇ��"�񿉈߿n�ȿas��\.���g��{�����u�w�Y���<��Y"�\���������F�uT��y0���L�Pi�AI���֎�����@>��澿f�տ ���:��������俴,ȿ����@���d�`���G��/F��\� ����򢿐�Ŀ�,�u�������ɒ�� ؿ�S���6��`L��&8������l���O�"y3�y����9���q� �����6�9�aXV�n�r�K�������q���]Q���Iƿ�ݿ���|����TTܿj&��4���?�}�u�U�HdD��K�vLi���������>Ͽ���Lz����jp�
zп�,���w�����������~�:/c�8F�ԥ*�������_�������3�'�C�}�_���{��  �  y�n�⿍�򸫿/�ҿ� ��V���'��a-���%��I�Y��5��<���,}�PJo�U���μ���ɿiq���Q��c(�]O-��%�������~ɿEF��K:����f�b�E�I�*��?�> ����Ӿ о�ھV�&
����+9�.W��l|����ȷ��ῧ������.+�%;,�#- ��/
�SE��O��j���t�ՙr����V�����ڿ=_��!�V�+���+����J�3�
��*���^�����Z��><��]"��W� N��x�ܾՀо9	Ҿ��MR������'�I�B���b�����������Ŀ�l�&��q#��-���)�Ʊ�8���LϿtܢ�>ք�b�o�}�y�!�������������#��*-�l,)�ח��C���׿��������Os�XP�,3��������7׾�yϾ]�վ���y����B@0�C�L���n�����������ҿǟ ��V�\�'��a-�n�%��I�����4��f��+}�qHo�_���ػ���ɿ�p��DQ�Hc(�O-�i%�˛������}ɿF��:��#�f���E���*��>�e ����Ӿ��Ͼ؞ھ��%
����*9� -W��k|�(�}ȷ���῁��u���.+�;,�- ��/
�AE��O��l��6�t��r�������-�ڿ^_��!���+���+�������翕
����������8�Z��?<�_"��X��P���ܾ^�о�Ҿ�OT�������'���B�6�b����	���#�Ŀ-m��&��q#��-��)�3������MϿgݢ�-ׄ�0�o�2�y�ꀓ�������=����#��*-��,)�����C�9�׿񟯿���#Ps��P�Z-3�[��w��%��b׾�|Ͼo�վv�������cA0�A�L��  �  ��c�~���B���ǡ���U#��F�:_�+�g�q;]��'B����Hu�"�������񍿏+���ſ�U�zL&��FI�k1a���g���Z�~�>�)�<���P��<N���sX�/g.��J��G����Ӿ���� 5����7ֶ�9�Ⱦ݃����"����C��'w�^��7�ӿ��
�w/�W�O��+d�"if�K�U���6��l��"޿�꫿����?��cƧ��{׿Q��2�G�R��te��^e���R�Hm3�h����ڿ�P��f~�6�H�vF#��'��=辇C˾�R��P��
r��\���a�о �|���*�S�Oe���ɯ����n��(;��hX��g��b�v�L��s*��B���ʿ�e���f��R����&"쿱���j>�l�Z���g��a�ՂI�h'�&��ǿ���Pj���:��I��� ��mݾ��þ�3��Ս�����"���0ھ� ��"/�ׇ6��c�'�����������pU#�kF��9_���g�/;]��'B����yt�5!�����������*���ſUU��K&�/FI��0a�F�g���Z�;�>��(��ￆP���M��'sX��f.��I�+F���Ӿˊ��3���﮾Զ��Ⱦȁ����+����C��&w��]����ӿ��
��v/�7�O��+d�if�9�U���6��l��"޿뫿����?���Ƨ��{׿*Q�>�2�m�R��te�$_e���R��m3�����ڿeQ���~�o�H��G#��(�o@�F˾1U���R��\t������]�о�!�|}�K�*��S��e��'ʯ�
�迨��(;�#iX�g���b��L�Rt*�<C���ʿ�f���g��S������"����j>���Z�Йg��a��I�/h'�&&�ǿ���8 j�	�:��J�	� ��pݾ��þ�6��Ȑ��v������ھ���10�Ĉ6��  �  G�g����y�ۿ
5�x�F��ct�c��g��_4����o�.�A�P���ۿ�P���ӡ��x��:7�����SL�oy�z�����������k�W6<�X=�p6̿N(��2�X��|%�%:��[ؾ�q���ϥ��u�������"��wz���ɾ��� ��5s?�z��3G��L-����&���V�⏀�Z�������u��tIa��o1������ȿ����Kˤ��3ÿ� �� ,��(\�#����h��
R��&}���\�7,��%���۶�R{��KbE����W���̾<ı��a��百՚�D8��ӿ��CԾ�1 �[� ��R����-�Ŀ�g���6�q0f�*��'i�������T}�`�Q���!��𿆥���j��ZU�� |ԿA���*<�L7k�������甋��x��YL��R����㣿Oo��Y4��'�N�徙W¾�>����G��� ��^P���:�� ᾢ�	�+/���g����4�ۿ�4�Z�F��ct��b��L��=4��k�o�ΏA����ۿ�O���ҡ��w�� 6�T��RSL��y�A�������ۘ���k�6<�'=�6̿�'����X�=|%�u9�PZؾIp��)Υ��s������ ��px���ɾ��3��Ur?����F���,����&���V�ҏ��M�������u��gIa��o1������ȿ����bˤ��3ÿ5� �� ,��(\�6����h��"R��@}���\�t,�(&���ܶ��{��|cE����
����̾�Ʊ�d��p陾Xך�f:�������DԾ�2 �� �:R�[����Ŀ�g�
�6��0f�U��Zi������U}��Q���!��𿓦���k��KV���|Կ���A+<��7k�Կ���������x��YL��R����h㣿�Oo��Z4�)����9Z¾[A�����J������R��8=��`ᾤ�	��+/��  �  �n�2���1���)��a��6��5ҝ� ���X�������w[�%�d��wc��e¯�-�ƿ���@�0���g��č��;�����٠��PӅ�|)U�����;߿�雿Q�]�Ll#��w��)�ʾ�᫾����~��E͍��ɓ�~;��KU���;㾠��b�@������1����p<��Lt�����:o���
��������`�H�E���-ݿ�R��<����ֿ����B��:z�B˔��W��O���Ô��Qz�%CB�[/�3�ſ����$yG�7�����N�n��z����뎾�����@��x�ƾ6����^�tV��앿�|ֿ%9���N�����Ϙ�D����o���9��.n�r6�T4�_�˿Ts��!庿�&�Ds�.6U�1̅�5�������/��#č�; h�̺/��f��J���`�w��"4�����ؾ5����1���������琾�]��ڐ����Ӿo��.J.�e�n�亨�����)�b�a��6��!ҝ����X������Ow[�� %�o��ob��O����ƿ/����0�7�g�sč��;���������+Ӆ�?)U�`��6;߿]雿��]��k#��v����ʾ�߫�>���|��Vˍ��Ǔ��9��WS���9㾸����@�&���g1�����I<��Lt�����-o���
��������X�H�B���-ݿ�R��<���ֿ2����B��:z�T˔�X��O���Ô�Rz�aCB��/���ſ����QzG�n��2���ﾾ�p����o���펾�����B��G�ƾ�����_�3V�8핿$}ֿ]9���N�����Ϙ�y����o���9���n��r6��4�u�˿^t��溿s'뿧s��6U�S̅�O�������/��.č�O h��/��f������%�w�{#4���,�ؾ����D4���ő�_���1ꐾ`��;����Ӿi��K.��  �  ��q�5���0����0�9�k��w��F���p��xP��1����d���+������9Ŀ�ʴ��Ϳ����7��r�J���V��-A��□��ҋ�uq^�?=$��濊x���O`�_N#����D�ƾ�ħ����o�������叾G)��D��w�߾"��Y�A��釿��ÿN��d�C�:)�&%��簨��U��v���/���dKQ�3�� �����7u���޿�T���J�p���g����황�Nv��
�����J�ǋ���˿�c����H��O����.㺾(X��^���L��� ������E%��˾¾^��D��X��(��.Uݿ�4�b�W�}ވ�Ѱ���������Ҟ��V~x�>��B�#>ҿi���A���xs���%�a^�U���u���GA��Y���#��?r�7��-��8���l{�	�4�Ch��վ���g(���荾忉����\Y���t���%о����.��q����������0��k��w��2��qp��VP�������d�3�+�ň���8Ŀ�ɴ��Ϳ���(�7�nr����V���@�������ҋ�7q^�
=$����5x��<O`��M#�������ƾ=ç������������㏾R'��B����߾<����A�W釿&�ÿ$��=�C�)�%��ڰ���U��n���(���\KQ�0��#��)���Nu���޿�T���J������g��������gv��%���׌J���D�˿Rd��*�H��P� �復庾�Z���	��UO���"������;'����¾����X�))���Uݿ15���W��ވ��������ݙ������~x��>�uC�<?ҿv���;���\t�P�%�ta^�w�������ZA��Y���#��?r�.7�.�9��jm{��4�Li�'վ����+��z덾��i���[���v���'оޅ�[�.��  �  �n�2���1���)��a��6��5ҝ� ���X�������w[�%�d��wc��e¯�-�ƿ���@�0���g��č��;�����٠��PӅ�|)U�����;߿�雿Q�]�Ll#��w��)�ʾ�᫾����~��E͍��ɓ�~;��KU���;㾠��b�@������1����p<��Lt�����:o���
��������`�H�E���-ݿ�R��<����ֿ����B��:z�B˔��W��O���Ô��Qz�%CB�[/�3�ſ����$yG�7�����N�n��z����뎾�����@��x�ƾ6����^�tV��앿�|ֿ%9���N�����Ϙ�D����o���9��.n�r6�T4�_�˿Ts��!庿�&�Ds�.6U�1̅�5�������/��#č�; h�̺/��f��J���`�w��"4�����ؾ5����1���������琾�]��ڐ����Ӿo��.J.�e�n�亨�����)�b�a��6��!ҝ����X������Ow[�� %�o��ob��O����ƿ/����0�7�g�sč��;���������+Ӆ�?)U�`��6;߿]雿��]��k#��v����ʾ�߫�>���|��Vˍ��Ǔ��9��WS���9㾸����@�&���g1�����I<��Lt�����-o���
��������X�H�B���-ݿ�R��<���ֿ2����B��:z�T˔�X��O���Ô�Rz�aCB��/���ſ����QzG�n��2���ﾾ�p����o���펾�����B��G�ƾ�����_�3V�8핿$}ֿ]9���N�����Ϙ�y����o���9���n��r6��4�u�˿^t��溿s'뿧s��6U�S̅�O�������/��.č�O h��/��f������%�w�{#4���,�ؾ����D4���ő�_���1ꐾ`��;����Ӿi��K.��  �  G�g����y�ۿ
5�x�F��ct�c��g��_4����o�.�A�P���ۿ�P���ӡ��x��:7�����SL�oy�z�����������k�W6<�X=�p6̿N(��2�X��|%�%:��[ؾ�q���ϥ��u�������"��wz���ɾ��� ��5s?�z��3G��L-����&���V�⏀�Z�������u��tIa��o1������ȿ����Kˤ��3ÿ� �� ,��(\�#����h��
R��&}���\�7,��%���۶�R{��KbE����W���̾<ı��a��百՚�D8��ӿ��CԾ�1 �[� ��R����-�Ŀ�g���6�q0f�*��'i�������T}�`�Q���!��𿆥���j��ZU�� |ԿA���*<�L7k�������甋��x��YL��R����㣿Oo��Y4��'�N�徙W¾�>����G��� ��^P���:�� ᾢ�	�+/���g����4�ۿ�4�Z�F��ct��b��L��=4��k�o�ΏA����ۿ�O���ҡ��w�� 6�T��RSL��y�A�������ۘ���k�6<�'=�6̿�'����X�=|%�u9�PZؾIp��)Υ��s������ ��px���ɾ��3��Ur?����F���,����&���V�ҏ��M�������u��gIa��o1������ȿ����bˤ��3ÿ5� �� ,��(\�6����h��"R��@}���\�t,�(&���ܶ��{��|cE����
����̾�Ʊ�d��p陾Xך�f:�������DԾ�2 �� �:R�[����Ŀ�g�
�6��0f�U��Zi������U}��Q���!��𿓦���k��KV���|Կ���A+<��7k�Կ���������x��YL��R����h㣿�Oo��Z4�)����9Z¾[A�����J������R��8=��`ᾤ�	��+/��  �  ��c�~���B���ǡ���U#��F�:_�+�g�q;]��'B����Hu�"�������񍿏+���ſ�U�zL&��FI�k1a���g���Z�~�>�)�<���P��<N���sX�/g.��J��G����Ӿ���� 5����7ֶ�9�Ⱦ݃����"����C��'w�^��7�ӿ��
�w/�W�O��+d�"if�K�U���6��l��"޿�꫿����?��cƧ��{׿Q��2�G�R��te��^e���R�Hm3�h����ڿ�P��f~�6�H�vF#��'��=辇C˾�R��P��
r��\���a�о �|���*�S�Oe���ɯ����n��(;��hX��g��b�v�L��s*��B���ʿ�e���f��R����&"쿱���j>�l�Z���g��a�ՂI�h'�&��ǿ���Pj���:��I��� ��mݾ��þ�3��Ս�����"���0ھ� ��"/�ׇ6��c�'�����������pU#�kF��9_���g�/;]��'B����yt�5!�����������*���ſUU��K&�/FI��0a�F�g���Z�;�>��(��ￆP���M��'sX��f.��I�+F���Ӿˊ��3���﮾Զ��Ⱦȁ����+����C��&w��]����ӿ��
��v/�7�O��+d�if�9�U���6��l��"޿뫿����?���Ƨ��{׿*Q�>�2�m�R��te�$_e���R��m3�����ڿeQ���~�o�H��G#��(�o@�F˾1U���R��\t������]�о�!�|}�K�*��S��e��'ʯ�
�迨��(;�#iX�g���b��L�Rt*�<C���ʿ�f���g��S������"����j>���Z�Йg��a��I�/h'�&&�ǿ���8 j�	�:��J�	� ��pݾ��þ�6��Ȑ��v������ھ���10�Ĉ6��  �  y�n�⿍�򸫿/�ҿ� ��V���'��a-���%��I�Y��5��<���,}�PJo�U���μ���ɿiq���Q��c(�]O-��%�������~ɿEF��K:����f�b�E�I�*��?�> ����Ӿ о�ھV�&
����+9�.W��l|����ȷ��ῧ������.+�%;,�#- ��/
�SE��O��j���t�ՙr����V�����ڿ=_��!�V�+���+����J�3�
��*���^�����Z��><��]"��W� N��x�ܾՀо9	Ҿ��MR������'�I�B���b�����������Ŀ�l�&��q#��-���)�Ʊ�8���LϿtܢ�>ք�b�o�}�y�!�������������#��*-�l,)�ח��C���׿��������Os�XP�,3��������7׾�yϾ]�վ���y����B@0�C�L���n�����������ҿǟ ��V�\�'��a-�n�%��I�����4��f��+}�qHo�_���ػ���ɿ�p��DQ�Hc(�O-�i%�˛������}ɿF��:��#�f���E���*��>�e ����Ӿ��Ͼ؞ھ��%
����*9� -W��k|�(�}ȷ���῁��u���.+�;,�- ��/
�AE��O��l��6�t��r�������-�ڿ^_��!���+���+�������翕
����������8�Z��?<�_"��X��P���ܾ^�о�Ҿ�OT�������'���B�6�b����	���#�Ŀ-m��&��q#��-��)�3������MϿgݢ�-ׄ�0�o�2�y�ꀓ�������=����#��*-��,)�����C�9�׿񟯿���#Ps��P�Z-3�[��w��%��b׾�|Ͼo�վv�������cA0�A�L��  �  񵊿�E�� ����᷿��Ϳ�5俲`��_��n�-�ҿ1౿fH����m�xUM���C�˧R�H%x��(���g���7ٿ��]�������߿��ȿ�s���.��h������I�u��Y�c�<��Z"�W��$�������G��U��z0�¦L�f�i��I��׎�����>��i澿��տf��;���������,ȿ����I���_�`�ׇG��/F���\�ӌ��z�M�ĿZ,����&���Z��U ؿHS��56���K���7��l�����l�"�O��w3����������3� �����R�9��WV���r��������.���Q���Iƿ�ݿZ�H|��]��Sܿ�%��X�����}���U��bD��K��Ji�����X��v>Ͽe���y���~��p濴yп-,��]w��$���.��~�~��-c��6F�/�*�<��ٮ����r������'��C�G�_���{�|���.E��ɧ��M᷿=�ͿT5�X`������쿝�ҿ�߱��G��@�m��SM�6�C��R��#x��'���f���6ٿ��Ȇ��"�񿉈߿n�ȿas��\.���g��{�����u�w�Y���<��Y"�\���������F�uT��y0���L�Pi�AI���֎�����@>��澿f�տ ���:��������俴,ȿ����@���d�`���G��/F��\� ����򢿐�Ŀ�,�u�������ɒ�� ؿ�S���6��`L��&8������l���O�"y3�y����9���q� �����6�9�aXV�n�r�K�������q���]Q���Iƿ�ݿ���|����TTܿj&��4���?�}�u�U�HdD��K�vLi���������>Ͽ���Lz����jp�
zп�,���w�����������~�:/c�8F�ԥ*�������_�������3�'�C�}�_���{��  �  v;������L�������ô��d��\�ղ�觿Ԝ���́���Z�`$9��$����[|'�ϥ?��Hc�=���`㚿{��K��M��� ��͐���������-��������i���I����|�xYT��4���!�rk��*���D���i�r���󝿣 ���+��
��b����{���8���߶�L<����������᏿�}u��TN�Ȏ0�H? ��^��.�wJ���p������࠿�ۮ�pݵ������g���u��)���q��֦���B���ꟿ�h���n�m�H���,�P �O� �9�1�{NP���w�A��E���V����d���ζ��"��􀴿�̵�]��洿YV�����䈿Լg��C��{)��1���"�`6��gV���~��g��C������=ö�s����崿������g������F7���ՙ��Y���a�`�=�{�&�=����$���:��\�J���{�������:������PL��6���>ô��d��Aղ��秿K���X́�k�Z��"9�s$�J���z'�7�?�CGc������⚿��cK������ ���������������������si��tI���|��XT��4�x�!�<j���*���D�T�i����^� ��T+���������e{���8��S߶�<��p���񾢿�᏿�}u��TN�̎0�a? ��^�<.�fwJ���p����ᠿ#ܮ��ݵ�����h��v��������~���_C���럿�i��|�n��H�D�,����� �i�1��OP���w�������������d���ζ��"��<���S͵�����洿�V��L򜿍刿d�g��C�f})�=3��"��6�iV��~�h���C��e����ö�Ӓ���崿+�������������8���֙�eZ��la�:�=�W�&�����$�E�:���\����"��������  �  ~9��<����ס̿���Ť�F���.�� Uz��d^�/oA� m&����h��1��+K�����,���G���d�����ƌ��z��td���V��;�ѿ���|���.!�����[�Ϳz<���U��#g�jJ�v�D�ydW��/��~������ݿ��e���D￮�ۿA	ſDE�������L��_ׅ�Bq�]�T�]8��q�\)�H� � �;�	������4�q~Q�W,n��m���萿����7����¿Jbٿ����R�����f�¿n��!����Z�&�E��OH���b��%��U����ɿK1�I���������^QԿ�����G��h����&��쐁�T�g��K�C�.��+����X���%����z�#�)E>�_-[��Uw�A���H��������Kʿ���_g�Gy���&�x�׿�����h��u��5Q�(�C���N��op�f��������VԿ�*��8�����㿁�̿�����Ĥ�틖����<Tz��c^�nA��k&�/�� ��.���I�J��k,�F�G�z�d�+��qƌ�4z��<d��~V��&�ѿ���j���!��\���Ϳ<��mU��
g�4J�+�D�"cW�;/��`}��u��9�ݿ���{d��TD�9�ۿ�ſ�D��g����L��(ׅ��Aq��T�38��q�^)�`� �; ���	�)��W�4��~Q��,n��m��+鐿^��8���¿�bٿ���R��
��n��+�¿5�����@�Z���E��PH��b�L&�����+�ɿ�1�;I��������鿇QԿس���G������'��u�����g�I
K�� /�e-���>����������#�LF>�h.[��Vw��������{������ʿH��h�z���'�[�׿�����i��ńu��7Q�$�C�o�N��qp�A���{³�6WԿq+��  �  em-��G'��.������п�Щ��U����l���J�2�.�������p��3�ԾE�Ͼ��׾mK�������4�`�Q�9�u�'$��ʞ��t[ڿ��������)���,�c#�*O��������͑��cx�Hsp���"���jҿ������!*�5�,�
�"�2��-��U�¿�����Q��	�`���@�oi&�-��������߾�Ѿ��о#�ݾ���av�.�#�I�=�(�\�с�Ý���5�����^��� �JH,��+�P����n�׿=d��㯈��q���u��������M(����&!��,��*����(4�:_߿>����1���z��ZU�q�7��m��	�\d�r�پ��Ͼ%�Ӿ6���� ��p�G�+��{G�+�h�����4����˿�Q�������%��c-���'���o���ǿd���w���o��~��嘿���y�������L&�m-��G'�p.�������п�Щ�6U����l���J�=�.��������}羛�Ծ��Ͼ:�׾�H�s��l���4���Q���u��#������e[ڿ��������)���,�N#�O�?�近���_͑�Tbx��qp�I��i����ҿ��A��=!*���,�Ŕ"��������¿e����Q����`�c�@�+i&� ��Յ����߾L�Ѿ>�о��ݾt���v���#���=���\�{с�=����6�����I_��� ��H,��+���2��?�׿e��������q��u�W��������(�0���&!�1�,���*����34�^_߿t����1���z��[U���7�o�	�g�(�پ5�ϾƢӾ����� ��q�N�+��|G��h�󒉿���P�˿;R����R�%�!d-��'�0�v���! ǿz����x���o�&�~��昿����N�������L&��  �  ��g�37^�#VD��J!�z���8����x���a��q4�������yؾ����,���ᜮ��Ҵ�ž�(߾#��|��|=��Hm��I���4ʿ��>o)�,K���a��dg�U�Y�b�<�A����迯���6I��g���<!����Ϳ�@�ք,�$AN�O�c���f�hW�A9�����N�����9aP�/�(�H�K��cϾ�̺�����������N�̾*꾷t	�%��AK��р��ܧ���ݿp���b5��]T�T�e���d��`Q�ݜ0��G��?Կ�Х�����1p��������~�T�8�dW�z�f�#|c��cN�+w-��	�לпL�����s���A��&��b����lǾq ��ˮ�?���`���Pվ�f��}��7`0��?[��Q���&��dd��3�m�@��	\�`�g�FH`��G��5$�.���z7¿d���,Ӎ�t嘿����0��� �:�C�,M^�F�g��6^��UD��J!�(��������x���a��p4�&�������vؾQ�����k���wд� ž�&߾!������=�_Hm��I���4ʿ��Go)�',K���a��dg�D�Y�?�<���������H������y ���Ϳ]@�x�,��@N���c�o�f�W��@9���j���������`P�ϯ(���cϾ�̺�������s��
�̾�*�Fu	��%��BK�hҀ�ݧ�/�ݿ���c5��]T���e���d�KaQ�H�0�H�[@Կtѥ������p��d��G��I~���8��W���f�)|c��cN�/w-�	���п������s�ΚA��'��c���⾕nǾ�"���ͮ�����ʆ��hRվ�h�����0a0��@[��Q��'���d�64�½@�V
\�Ϲg��H`�j�G�6$�R����8¿����Nԍ��昿¼��1��Y ���C��M^��  �  �����]r��MD�&����׿�@����c���,�x���޾Ҽ��,g������T��{t���C����þ�,辤���7��Ys��㦿�1�N���O���z�� ��]���-�����h��y9����]ѿ`���zݢ��㻿w���QH$�PT�,e��9���1���,��`�c��4����;��{�����N�����u��RIҾ\u��y�����������������tξ���*��uH�!ˆ��?���\��.���^�ui��&������������Y��~)����������������Gg˿��U4��c�T���A������FMT�?#$�����h�{�;�<�Z���%�LLǾ�^��l���:z��/͛�����Pպ�wھ
����'�4p\��˕�}пʱ��>��rm��W��sԏ��"��q�v�}�I�Q�a��(���a����wm޿=,�9BD��Pr���������*r��MD������׿n@���c�2�,�����޾�����d��Ɠ��]R��0r���A����þ�*����7�(Ys��㦿�1�W���O���z�� ��_���&�����h��y9����j\ѿ�����ܢ��⻿�����G$��OT��d�p9���1���,���c�N4�g�;��-����N����6u���HҾ-u��y��ܐ����5��?����uξ:���֌��uH��ˆ�|@��]�\�.��^��i��W���%��-����Y��~)�����i������S����g˿���4�G�c�T���A������CMT�B#$�&�������{��<�9���'�}NǾ�`��Ҍ���|���ϛ������׺�Ayھ����'�*q\�6̕��п��c�>��rm��W���ԏ�2#����v��I������^�������B����n޿�,��BD�!Qr�����  �  >��d��w����^�'�&����k��Lj��y+����#�Ѿ��|�������\����<���)��GC���K۾^v
�]+7�)]|�?���/ ���2�ik�� ��aϟ��£��Ǚ��d���R�j��a}�RT������xMοf��$s9��*q��i������L���ٗ�����D�K�j��<ҿ����@R�������Ͱľ����3▾v���!A��&���N���0�����뾭=���J�[r��F�ɿ����eE��I}�kӕ�����
��s����:w�]�?��K���ӿ�\�������࿭i���K�ˇ��y��DS��?���e��qAq�6�8�wF��l��4���t=�Ѓ�k��З���+���<��S���-Ώ��ؙ�n=���;V����	&���a�$������ �!QX�_4��[{��X��������]�d��-�"���Ŀ����N��������'�T�^����w ����E��^��ɝ^� �&���쿹j��YKj��x+����B�Ѿ��Y����!����:���'��VA��)J۾�u
��*7��\|�-���/ ���2�k���jϟ��£��Ǚ��d��VR�"���|翓S�������Lο����r9�/*q�|i�������L���ٗ������K��i�|<ҿu��J@R������l�ľe���3▾����A��������� �����Z>���J��r����ɿ��fE�@J}��ӕ�����>������V;w�τ?�cL���ӿ�]��ˊ������i�	�K�⇁����IS��=���e��jAq�6�8��F��l��s��2u=����P��癹��-��6?�������Џ��ڙ��?���;a����
&���a������� �qQX��4���{�����Y��������d���-�S#�� �Ŀꕯ�DO������{�'�͗^���� ���  �  �m��.�w�J�Y�Nd0�g������N��ʂE����߾Ż��`z��d5��'z��u���|��D��׫����_��O��A"T���q�Ͽ����:��a�[|�{&��^�r��Q��&��a����������a��U����ݿ�����>� ie�t�}�)̀���o�*�L�j�!��M�@���u���1�����ξ�֨�a���X���v�@Hv��=��M���C����ɾ*� ��+�v�l�ڥ�-�� ��.H��ll��P��e�v�h��tC���3快���n������s>���T��H"��L�ݑo��̀���}�ze�/�>��\�`�׿����[�8� �Y�Z���y����m�~��Vu���x��ф����꯾��پYY���>�A��	���C� �O�+�φU��Ou��[���z���]��<5���
�1Tп�!��S��N����ʿX���o0��Y��w��m����w��Y�%d0��f�V����N���E�J��n�߾󹳾jx��Q3���z�iu���|��B�������﻾��ғ��!T�
��~�Ͽ���:�%�a�o|�~&��R�r��Q���&�!a��g������`������1�ݿa��&�>��he��}��̀���o��L�+�!�9M�?��E�u��1�����ξ�֨�1���X��d�v��Hv�7>�����0���4�ɾ�� ���+�Y�l��ڥ����O��f.H�[ml�Q���e���h�(uC����忎����n��_���,?���U���"�A�L���o��̀���}�ze�%�>��\�l�׿��@�[��� ��Z�\���{�����~�G[u�Q�x� Ԅ����,쯾��پNZ��>��A�������� ���+�'�U�cPu��[��Kz���]�5=5�!�
�qUп#��OT��|����ʿݚ�p0�J�Y�a�w��  �  ��w�a6m�V�P��@)�� �a
���^��NC���c⾻�c����&K����{����(������J���]&��CQ������)ɿ*D	��l2��$X�Pq�?w��@h��eH��7 �BB�b���<w��@u��	����Eֿ�T�J�6��[��s�"�v��^e��+D��g����R���q�O�0��W��Ѿ:2��D#��_���r}���|�����N���ҡ̾��p�*��h��t��:�߿?��;�?��Vb��u��|t��'_��m;����ݿI����t���u��܉��������(D��ke���v�� s�o�[���6�C����пe����X�=$ �f���`Vþ�颾Ib�����'�{� ]�O2������.��/Qܾ�w���<�v���GO�������$��L�z�j��w�po��lT�A�-�<���sɿ�{���s��Zy���ÿ���W)���P�)Em�Q�w�%6m�%�P�~@)�� �
���^��dMC�U�����ﶾg�ꗉ��H����{�轁�����������\�:&��CQ�z����)ɿ9D	� m2�%X�.Pq�?w��@h�beH�s7 ��A󿻉���v��wt��9����Dֿ T���6���[�ts�Ύv�t^e�h+D��g�B��􄧿sq�Њ0��W���Ѿ�1��#��_���lr}�f�|�l���	�����̾���5�*���h�au����߿�����?�Wb�P�u�}t��'_�&n;����ݿ+���}u��iv������/��B���(D��ke���v�� s�g�[���6�A����п����c�X��$ �����5Xþ�뢾xd��M�����{��a��4��F����0��,Sܾ�x���<���O��b�����$�v�L���j�[�w��po�rmT���-����7uɿ}��u���z���ÿr��qX)�I�P��Em��  �  (�Y��XP��7����'��*~���>�6����*¾�g���z�����Bć����"���֟��D�ɾ����k���J��Ї��䷿k�������1>���S��Y��)L�߸0��:� kڿ�(����������U���џ��;�����!��aA�yU��rX���I�P-�Y[
���ѿO]��gf�O.�����p۾ ���u��S���Έ�Hj��� ��]���e��g�־%{�nG)��_��4��,˿v��_)���F�M�W���V��QD��%�d���yǿ. ��h������Aޣ��ӿ�W
��-���I���X��[U��CA���!�����%���o��XQ�C��?��_�;�i��������ㇾډ�5��������k���k�P7��9��u�A9���߿�1�g;4�4FN��bY�p[R�[;�E���+￡�������>���3��R���s�6�q�7�*}P�߂Y�mXP�ܪ7����'�4�)~�J�>�r�߼�G¾�e���x��Ё�������������ם����ɾ^��k�8�J��Ї��䷿��������1>���S��Y��)L���0�z:�xjڿ!(��չ��؊���������q���_�!�oaA��xU�prX�W�I�-�[
�)�ѿ�\��wff��N.����mp۾Ø���t��S��ψ��j��2!���]���f����־�{�1H)�h_�u5���,˿Tv�$`)�!�F���W�!�V�-RD�Y�%�Ԭ��zǿ
!���h��S ���ޣ��ӿ�W
�$-���I��X��[U��CA���!�����%��#p���XQ�������M�;�k�����i���凾u܉�� ��4����m���m�D8��9��u��9����߿2��;4��FN�cY��[R��;�����,�է������k���U��e���r迪�׻7��}P��  �  �0��)�+?�����o�ſ������n��X=�W�������3پn���k������<���$랾�u��%@¾���$���� �w�F�<N|�v����	ѿ���6���+���/��%�R��F�T@���9���u�%�m����y
��՞ӿl���?��,��H/�s�#�x5�-�{�������\�t(0��6����Y�ξ���ꣾ������������ʲ�Hg˾�0�u?��,�C�V�j������<�h�*�!�;�.���-�b�����
mٿs���ч�ko�� s��ߍ��1��iE��;�#��G/���,������ӴֿD;������L�xX$�ٝ�����/žOv������ޙ��<�������.�վ���bt���8��h��;��N���	��٢��~'���/�w*��Y�j���Kȿ΃��^���Kl�w�|����Q�¿�\������)��0��)��>�m���"�ſ\����n��W=���������1پJ���"���&��ѵ���螾@s���=¾���N��R� ���F��M|�i����	ѿ&���6���+���/��%��Q�NF��?��:9����u���m����	���ӿ���?���,�JH/�*�#�65�����A���\��'0�@6������ξ����ꣾ���ၚ�����=˲�0h˾2�@��,��V���� ��U=�gh���!���.�`�-�Ɉ�����mٿL����ч�
o�3"s�����Y2���E�H�X�#��G/���,�������ֿe;��殁��L�=Y$�Ğ���02ž�x��G��ᙾJ?��u��<��Q�վ���Su���8��h�_<��̌�����)���~'�F�/�xw*�nZ�k���Lȿ򄜿<_��9Nl���|����D�¿�]����=)��  �  ���0����K%ɿ�⧿GK��i�i��'G���+���(V����jɾ?����U���?����;��辯m�ڶ�-h1�-N�|�r����������п�c�v���)�Φ���ݿ������np�m	P��J�o�^�Ap��x���JͿ����	���#����߿�ǽ�ޱ��$���*]�d=���#��������ؾ~�¾��c��F�����վC���O.!�J:��;Y�����o�����S�ۿY��]��������!tѿ���������b�$K��N�ǖk�����䳿|�ٿ3������ۤ�-n�}|Կ���&���Vw�I�Q�EM4��(���s�.aоe������������ƾ��޾���Κ��)���C�`e�Y���k��pXſ����) ��}��F����!�Ŀ�y���U�� �W��I�mU���z���������8��: �����/�����$ɿ�⧿�J��Īi��&G���+���U�����ɾ����S��I=��j�;!�辖l���bg1��N��r�������¹п�c�u���)�������ݿ9�����lp�&P�aJ��^��o��Nw��<JͿ�ￇ	���������߿*ǽ�}����#���)]��c=�r�#�������Ѳؾ��¾J��{c������V�վ�C����.!��J:��<Y�����p��>����ۿ�����\��� ��tѿ؏��a���_�b��	K�d
N��k�����e峿֜ٿq��������>n�|Կ9���K&��Ww� �Q�'N4��)�-�����cо���-�������,�ƾ�޾1���Л��)���C��`e����#l���Xſ/��.* ��}�G����!�Ŀ�z���V��$�W��I�wU�q�z�}��������8�-; ��  �  ��ÿ����j���~��4�����ݽy��e���P�5e:��E#�Q��ш��i��G$ܾ�"澦N���7�;_(��?��U��j�j~�Jӊ�����)��트�3�¿^�¿�������D`���g�\A�Z +�L�&��\5�Q�T�mc���J��&
���m��tĿG��X����/ǐ�r��V�r���^��I�I�2�����J�7��%�޾Ѫݾ���G��T�/0�kG�%�\�J�p��؂��<���:���������Q�ÿB����1���������Y��8�Щ'�ѽ)��>�7b�\����a���5��?¿gÿP������5���(C��Mf��4:l���W�B�^�*���ht�'7�&pܾ�ᾠ`���~�1� ��7��bN��Mc�	rw�3�����������ĳ�S��KĿ�ܼ��r������[+v�`eL���0�CE&�ۍ.�އH�q�9������4b��6�ÿ0��@j��`~��蘕����4�y�Q�e��P�9d:��D#���0������n!ܾ ��K���6��](�q~?�'�U�� j��i~�ӊ�����)��ኸ�#�¿B�¿��������_���g��ZA�(+��&�S[5���T��b���I���	��Gm���Ŀ�ｿpX������Ɛ�#����r�z�^�I�
�2�����J�<��V�޾-�ݾ���%H�VU��0�G�ށ\��p�(ق�!=��9;��W���������ÿ�����2��a�����IY�:8�C�'�,�)�>�*8b�Ϙ��%b��66��8?¿�ÿq�����e���jC���f��;l���W�/B���*�F���u�
:�sܾ��Ac��2��Q� �
�7�tcN��Nc��rw�������������_ų�����Ŀ�ݼ�qs������H-v�ZgL���0�9G&���.���H��q���������b���  �  ������&���P���X��J%��	픿=D��&�����v�îV�"�6����
C��o�p���!�K�=���]��/}�/����{���0��K����=��6u���>��w���[0��������q��:Q��2��Y���
�m���g�9&���B��dc�M�y����;��|J��)Ԕ��2��o���tN��'2��:�������FNl�G�K�'o-�?�0H	�(���!��j*��:H���h�2��o���ٓ��Q�����"/��w����P��K���2����t����f��rF��(�w/��L���	��)�P�.�ܛM��n��U���c��%Y���J��݊��G5�������C���������+����a�W-A��$�Î����O�r|�'�3�>
S�y=s��Y����������6���j��	C�����?#��3���k����{��#\��<� � �e>�_����X�g�8��X�Jx��<�������������P���X���$���씿�C������z�v���V���6�k���A�)n����x�!�ʸ=�o�]�s.}�����{���0������=��u���>��X���30��g����q��9Q��2��X���
�;��Df��&�c�B��cc���홌�;��J���Ӕ� 2�����)N���1�����u���
Nl� �K�o-�B�IH	�V��9"�9k*��:H�w�h�h2�����$ړ��Q�������/��
���UQ��񨓿ᘍ��u���f�7tF���(��0��M�د	�+�Z�.���M��n��U���c��XY���J������5������CD������@��h,�� �a��.A���$�U��(�����}�o�3�fS��>s�6Z��{�������O7��3k��qC�����#���3���l��N�{�|%\�\<�Ѥ �:@��`�o�����8��X�YKx��=���  �  �f��z�ٺ��)n��mi��N8��_r����ÿA���)̧�J���+yn�>�F�x�-�|]&��1�gN�c�x��$��P���{��� Ŀ;���"2����&�����_Ov��.b��,M���6�m�?m
����U�t�ܾ�V龲c�����9,� IC��Y�iWm���r��������㫿񶺿�Yÿ6���S?����O6��P�_��z<��#)��(�;z9��C[��u���`��4=��O�����ÿ���{����V���z���9��K�o��Z[�c�E�V�.����K�P�뾷GݾK߾e���Q��D�3���J�J�_�+t����k���pl7��ڃ���Ŀ(־�?쮿D闿~���R��4�	�&�C�+��C�yi��Č�+F��@�-ÿ�3¿qȷ��>�������';}���h�]T��8>�'���.���X&�Xܾ�X�6(����v�$�̫;��Q�)�f�C�z������m��'i��8��	r���ÿȘ���˧������wn���F�Ԝ-��[&�I�1�ZeN���x��#������֍��sĿȘ������}&��m��Ov�N.b�n,M���6��~�dl
� ��|S�5�ܾ�T龅b�h���8,��GC��Y�uVm�� ����������㫿�����Yÿ���,?�����<6��@�_��z<��#)��(�~z9�CD[�v��a���=������X�ÿi��󰭿W��g{��`:����o�>\[���E���.� �GM���VJݾ�߾����R����3�%�J���_��t�D���������7��U���GĿ�־��쮿ꗿ�~�v�R�M4���&���+�fC�azi�DŌ��F����-ÿ�3¿�ȷ��>����y��<}���h�S^T�U:>��'��������)徱ܾ�[�P+�����Ɋ$���;�"�Q��  �  ��H�%�k�����A���q˿��뿗���v�V���Y�N{��R����;x���S��'I�Y�WЁ�s����ƿ�꿊���p��;�����7sÿ����m!���Gc��.B�ȷ'�5u�����6ݾ4�ž�;��h����x��ȴѾ������f���5���S��y�J����v���Zֿ����`����~���*�׿�˱�8Ŏ��Hi��)M�a�K���d��X��������ӿ���������i����ڿ�)���՘��~�DOW���8�A���
�m�jԾ;��Z��Bb��|�þ�,ھ]���/�%���>�d,_�{s���Y�����N�����>����,�1˿*q��y܄�X]�¦I�'Q��r�y�j;��{�߿����5K�ƈ�;����ο2������SYp�>RL���/�)���b���� �̾���E��=P��>5ʾ��W����*-��H�s�k�M�������.˿=��l���v��U��0Y㿡z������2:x��S��%I�ߖY�eρ�r����ƿK��,��`p�\;��V���rÿ����1!��6Gc�.B�?�'��t�{���*5ݾY�ž�9��I���~v����Ѿ`�����e���5���S��y�강�[v��QZֿ����D�����Y����׿�˱�0Ŏ��Hi��)M���K��d�Y��Ѡ���ӿ��������Թ��Kڿ*��^֘��~�wPW�9�8����k�
��o��lԾ���� ���d����þ�.ھ����/��%�G�>��,_��s���Y��h����Nῒ���+?������1˿r��h݄�1]���I��(Q���r�.�	<���߿���cK�������οh2��T���(Zp�:SL� �/�o��.d�����̾/���2H��CS��!8ʾ���QX����+-��  �  ��?�c+r����P�ȿõ�������)�70��8(�xm��V�����|�����z��yl��y�������˿8 �����"+���/��&�N�A��^㽿N"��:ye��6����x����Ӿ�Ǹ�>7��+䛾���"���e����ƾZ�����?:&���N�i~��_����ٿQ���rk-���.���"���I⿃����G��
�q���o�q@���뫿 ]ܿ(	��� �pH.��J.��� ��	�BU߿h���j5���T�E*�i��A
���ɾ�����ס��M���@������M���[о�󾘻�GA2��u_�H��O���O뿯��X�$���/��Y,�G�S9�P�п�բ�؃�6'm��bw������պ�J���Ј&�g�/�x-+�t��K��;ο�<��R�x�|�D�������0�޾����{���e��9���mt��
���.���۾���n�ů?��*r������ȿ����e��W�)�0��8(�*m�
V�����������z�xl��x��ے���˿�7 �2��k"+�z�/���&��M����㽿"���xe�e�6�����w��%�ӾƸ�s5��>⛾������M���βƾU�����V9&�±N�~�������ٿ,�ˮ�Wk-���.���"���I�|����G��$�q��o��@���뫿6]ܿ,(	�¡ ��H.�K.�)� �N�	��U߿삮��5���T�|*������q�ɾO����ڡ�=P���B��1���}O���]о���M���A2��v_��������������$���/�MZ,����9�L�п�֢�ك�)m��dw�����aֺ��J�6���&���/��-+���
L��;ο =���x�\�D��������޾�����}���h�� ���Cw���������(۾���o��  �  ��A�4���ڮ�>��T�HX9�
OQ�'}Y�{O��6�-�Y����?܎�ʅ��
���M�������/�<�t7S��<Y�N+M�Jz2��;�Ibܿ�p��Z�q��B6�VU�Y��_���΢�L���������������n���ݯ�sо|8��t!"�m�T�GЎ��V��7� ��#��B��V��$X�oH�:+�i�:�пPԡ��>����:����~ʿ.��Ay'�^�E��=W��&W��E��'�5����ǿq���,�[���&���hzԾٲ��Z��^���g?��w��-���n���C?��]�ݾ��	��0��*j�����aտ�O���.�K�J�a�X���T��?����(���Ⱦ�V���7��z���Ug����ݿ.�ɂ2��PM��DY�DS���<�!��H8�մ�z���оG�F��$��Ǿ�C���ޖ�����+����݊��>��ڧ����þ�z��ȫA��3��Wڮ���7�'X9��NQ��|Y��zO��6������(��Aێ�
Ʌ��	��tL�����3����<�7S��<Y��*M�z2�];��aܿ�p����q�GB6��T���証�j̢�PJ���������������l���ۯ��о�6��� "���T��ώ�VV��� ���#���B�jV��$X��nH�:+�i�3�пSԡ��>����[����~ʿH��ay'���E� >W��&W��E��'�r��o�ǿ����N�[��&�=���|Ծ�۲�:]��ґ���A���
��G���^���A����ݾI�	���0��+j����bտ�O���.���J���X�=�T���?���3���ɾ�`���8��j���2h����ݿZ.��2�QM�EY�cS��<�9��|8��մ�͑����G�G��&� �Ǿ0F���ᖾm�����~���uA��D����þ�|����  �  [�F��؈�}��n��<�+��~R�YSn���w��l�^�N��'��'�����~��&���p����̿��p/0��PV�Aop�1vw�ʈi��{J��S"�L�����|~�Ԝ9��^��پ�`���g������(�~���{�����G��_��Εž�`����"���\��Ƙ�LRԿ&���39�]p]��s�)v�W�c��B��l�@�翝)��˕��S��F����࿻����=� �`�u�_u�g�`�Y�=�u��2ܿ�����d��(�op���8ʾ�`���!��^
��k|���}�IG��]1���୾q3Ծ�M��3�&uu�X�����|���LF�(�f���v��=r�y�Y���4�5(�1�ҿ{���@�������(��/*��t~"��yJ��i��yw�_`p�mLV��$0�����ſt�>�M�i���,�.꼾	Ş�#ߋ�&X��lu{������S���.���Ḿ������F�H؈��|��R�� �+��~R�1Sn���w��l��N�2'��&������w�����T����̿z���.0�KPV��np��uw�v�i�|{J�WS"��K��o��s{~�:�9��]���پ8_��:f��͈��}�~��{�����E��]���ž�^����"�3�\�BƘ��QԿ����39�>p]���s��(v�F�c��B��l�:�翠)��ؕ��j��g��������ף=�$�`�9u��u���`���=�����ܿ������d� (��r��q;ʾ
c��$������o|�*�}�^I��J3���⭾5Ծ�N�H�3��uu�����쿸��MF�}�f��v�$>r���Y�(�4��(�H�ҿ����H��험�{)���*���~"�zJ�8�i��yw�{`p��LV��$0���Ռſ����M�M���.�y켾�Ǟ��ዾ�Z���z{�[���1V���0���㸾�徯��  �  �I��鋿�Ŀ�����2��[���x�9i����v���W��.�Uu�Sǿ����u��Zڥ�f�ӿ/3��7�6�_��"{�kE����s��_S�
)��Y���I���΁��^;�I+��׾���r,��ZZx�r�u�����֋���>�¾j���~x#��_�m�����ۿ��[1A��Hg�#�~���o n��^J�]��Jh�齶�3������w����������E���j�b�������j���E�܈�5��ར�oQh��	)��/���cǾ%�������1���&�u��dw��삾ȹ��k���ҜѾ�����4��z�0�������^8$�l�N�Aq������}���c�-e<�ݵ��Vڿy�������O᜿
E���? �i:)�AES���s��E��k#{���_�,�7��N�?�˿I��UZP���F?�uι��O���t���"|��
u�O�z�톾+���䳵����6��
I��鋿�Ŀl����2���[���x�i��Y�v�K�W�K.��t�\ǿ����t��;٥�D�ӿ�2�{�7���_�m"{�9E��:�s�N_S��)��Y��NI��΁�B^;��*�w׾G���퓾M*���Vx���u�����ԋ��_�¾�����w#�T�_����T�ۿ۽�91A��Hg�	�~�哀�^ n��^J�U��Ch�콶�@���������:�������E��j�w�������j� �E������g����Rh��
)�2��QfǾ����-���������u�iw������0���r�ѾP��m�4�� z����������8$���N��q����6	}�u�c��e<�i��Xڿ��������I✿�E��@ ��:)��ES���s��E���#{���_�?�7��N�x�˿TI��[P�{�LA龷й� R��Qw���'|��u�y�z��{��������⾒7��  �  [�F��؈�}��n��<�+��~R�YSn���w��l�^�N��'��'�����~��&���p����̿��p/0��PV�Aop�1vw�ʈi��{J��S"�L�����|~�Ԝ9��^��پ�`���g������(�~���{�����G��_��Εž�`����"���\��Ƙ�LRԿ&���39�]p]��s�)v�W�c��B��l�@�翝)��˕��S��F����࿻����=� �`�u�_u�g�`�Y�=�u��2ܿ�����d��(�op���8ʾ�`���!��^
��k|���}�IG��]1���୾q3Ծ�M��3�&uu�X�����|���LF�(�f���v��=r�y�Y���4�5(�1�ҿ{���@�������(��/*��t~"��yJ��i��yw�_`p�mLV��$0�����ſt�>�M�i���,�.꼾	Ş�#ߋ�&X��lu{������S���.���Ḿ������F�H؈��|��R�� �+��~R�1Sn���w��l��N�2'��&������w�����T����̿z���.0�KPV��np��uw�v�i�|{J�WS"��K��o��s{~�:�9��]���پ8_��:f��͈��}�~��{�����E��]���ž�^����"�3�\�BƘ��QԿ����39�>p]���s��(v�F�c��B��l�:�翠)��ؕ��j��g��������ף=�$�`�9u��u���`���=�����ܿ������d� (��r��q;ʾ
c��$������o|�*�}�^I��J3���⭾5Ծ�N�H�3��uu�����쿸��MF�}�f��v�$>r���Y�(�4��(�H�ҿ����H��험�{)���*���~"�zJ�8�i��yw�{`p��LV��$0���Ռſ����M�M���.�y켾�Ǟ��ዾ�Z���z{�[���1V���0���㸾�徯��  �  ��A�4���ڮ�>��T�HX9�
OQ�'}Y�{O��6�-�Y����?܎�ʅ��
���M�������/�<�t7S��<Y�N+M�Jz2��;�Ibܿ�p��Z�q��B6�VU�Y��_���΢�L���������������n���ݯ�sо|8��t!"�m�T�GЎ��V��7� ��#��B��V��$X�oH�:+�i�:�пPԡ��>����:����~ʿ.��Ay'�^�E��=W��&W��E��'�5����ǿq���,�[���&���hzԾٲ��Z��^���g?��w��-���n���C?��]�ݾ��	��0��*j�����aտ�O���.�K�J�a�X���T��?����(���Ⱦ�V���7��z���Ug����ݿ.�ɂ2��PM��DY�DS���<�!��H8�մ�z���оG�F��$��Ǿ�C���ޖ�����+����݊��>��ڧ����þ�z��ȫA��3��Wڮ���7�'X9��NQ��|Y��zO��6������(��Aێ�
Ʌ��	��tL�����3����<�7S��<Y��*M�z2�];��aܿ�p����q�GB6��T���証�j̢�PJ���������������l���ۯ��о�6��� "���T��ώ�VV��� ���#���B�jV��$X��nH�:+�i�3�пSԡ��>����[����~ʿH��ay'���E� >W��&W��E��'�r��o�ǿ����N�[��&�=���|Ծ�۲�:]��ґ���A���
��G���^���A����ݾI�	���0��+j����bտ�O���.���J���X�=�T���?���3���ɾ�`���8��j���2h����ݿZ.��2�QM�EY�cS��<�9��|8��մ�͑����G�G��&� �Ǿ0F���ᖾm�����~���uA��D����þ�|����  �  ��?�c+r����P�ȿõ�������)�70��8(�xm��V�����|�����z��yl��y�������˿8 �����"+���/��&�N�A��^㽿N"��:ye��6����x����Ӿ�Ǹ�>7��+䛾���"���e����ƾZ�����?:&���N�i~��_����ٿQ���rk-���.���"���I⿃����G��
�q���o�q@���뫿 ]ܿ(	��� �pH.��J.��� ��	�BU߿h���j5���T�E*�i��A
���ɾ�����ס��M���@������M���[о�󾘻�GA2��u_�H��O���O뿯��X�$���/��Y,�G�S9�P�п�բ�؃�6'm��bw������պ�J���Ј&�g�/�x-+�t��K��;ο�<��R�x�|�D�������0�޾����{���e��9���mt��
���.���۾���n�ů?��*r������ȿ����e��W�)�0��8(�*m�
V�����������z�xl��x��ے���˿�7 �2��k"+�z�/���&��M����㽿"���xe�e�6�����w��%�ӾƸ�s5��>⛾������M���βƾU�����V9&�±N�~�������ٿ,�ˮ�Wk-���.���"���I�|����G��$�q��o��@���뫿6]ܿ,(	�¡ ��H.�K.�)� �N�	��U߿삮��5���T�|*������q�ɾO����ڡ�=P���B��1���}O���]о���M���A2��v_��������������$���/�MZ,����9�L�п�֢�ك�)m��dw�����aֺ��J�6���&���/��-+���
L��;ο =���x�\�D��������޾�����}���h�� ���Cw���������(۾���o��  �  ��H�%�k�����A���q˿��뿗���v�V���Y�N{��R����;x���S��'I�Y�WЁ�s����ƿ�꿊���p��;�����7sÿ����m!���Gc��.B�ȷ'�5u�����6ݾ4�ž�;��h����x��ȴѾ������f���5���S��y�J����v���Zֿ����`����~���*�׿�˱�8Ŏ��Hi��)M�a�K���d��X��������ӿ���������i����ڿ�)���՘��~�DOW���8�A���
�m�jԾ;��Z��Bb��|�þ�,ھ]���/�%���>�d,_�{s���Y�����N�����>����,�1˿*q��y܄�X]�¦I�'Q��r�y�j;��{�߿����5K�ƈ�;����ο2������SYp�>RL���/�)���b���� �̾���E��=P��>5ʾ��W����*-��H�s�k�M�������.˿=��l���v��U��0Y㿡z������2:x��S��%I�ߖY�eρ�r����ƿK��,��`p�\;��V���rÿ����1!��6Gc�.B�?�'��t�{���*5ݾY�ž�9��I���~v����Ѿ`�����e���5���S��y�강�[v��QZֿ����D�����Y����׿�˱�0Ŏ��Hi��)M���K��d�Y��Ѡ���ӿ��������Թ��Kڿ*��^֘��~�wPW�9�8����k�
��o��lԾ���� ���d����þ�.ھ����/��%�G�>��,_��s���Y��h����Nῒ���+?������1˿r��h݄�1]���I��(Q���r�.�	<���߿���cK�������οh2��T���(Zp�:SL� �/�o��.d�����̾/���2H��CS��!8ʾ���QX����+-��  �  �f��z�ٺ��)n��mi��N8��_r����ÿA���)̧�J���+yn�>�F�x�-�|]&��1�gN�c�x��$��P���{��� Ŀ;���"2����&�����_Ov��.b��,M���6�m�?m
����U�t�ܾ�V龲c�����9,� IC��Y�iWm���r��������㫿񶺿�Yÿ6���S?����O6��P�_��z<��#)��(�;z9��C[��u���`��4=��O�����ÿ���{����V���z���9��K�o��Z[�c�E�V�.����K�P�뾷GݾK߾e���Q��D�3���J�J�_�+t����k���pl7��ڃ���Ŀ(־�?쮿D闿~���R��4�	�&�C�+��C�yi��Č�+F��@�-ÿ�3¿qȷ��>�������';}���h�]T��8>�'���.���X&�Xܾ�X�6(����v�$�̫;��Q�)�f�C�z������m��'i��8��	r���ÿȘ���˧������wn���F�Ԝ-��[&�I�1�ZeN���x��#������֍��sĿȘ������}&��m��Ov�N.b�n,M���6��~�dl
� ��|S�5�ܾ�T龅b�h���8,��GC��Y�uVm�� ����������㫿�����Yÿ���,?�����<6��@�_��z<��#)��(�~z9�CD[�v��a���=������X�ÿi��󰭿W��g{��`:����o�>\[���E���.� �GM���VJݾ�߾����R����3�%�J���_��t�D���������7��U���GĿ�־��쮿ꗿ�~�v�R�M4���&���+�fC�azi�DŌ��F����-ÿ�3¿�ȷ��>����y��<}���h�S^T�U:>��'��������)徱ܾ�[�P+�����Ɋ$���;�"�Q��  �  ������&���P���X��J%��	픿=D��&�����v�îV�"�6����
C��o�p���!�K�=���]��/}�/����{���0��K����=��6u���>��w���[0��������q��:Q��2��Y���
�m���g�9&���B��dc�M�y����;��|J��)Ԕ��2��o���tN��'2��:�������FNl�G�K�'o-�?�0H	�(���!��j*��:H���h�2��o���ٓ��Q�����"/��w����P��K���2����t����f��rF��(�w/��L���	��)�P�.�ܛM��n��U���c��%Y���J��݊��G5�������C���������+����a�W-A��$�Î����O�r|�'�3�>
S�y=s��Y����������6���j��	C�����?#��3���k����{��#\��<� � �e>�_����X�g�8��X�Jx��<�������������P���X���$���씿�C������z�v���V���6�k���A�)n����x�!�ʸ=�o�]�s.}�����{���0������=��u���>��X���30��g����q��9Q��2��X���
�;��Df��&�c�B��cc���홌�;��J���Ӕ� 2�����)N���1�����u���
Nl� �K�o-�B�IH	�V��9"�9k*��:H�w�h�h2�����$ړ��Q�������/��
���UQ��񨓿ᘍ��u���f�7tF���(��0��M�د	�+�Z�.���M��n��U���c��XY���J������5������CD������@��h,�� �a��.A���$�U��(�����}�o�3�fS��>s�6Z��{�������O7��3k��qC�����#���3���l��N�{�|%\�\<�Ѥ �:@��`�o�����8��X�YKx��=���  �  ��ÿ����j���~��4�����ݽy��e���P�5e:��E#�Q��ш��i��G$ܾ�"澦N���7�;_(��?��U��j�j~�Jӊ�����)��트�3�¿^�¿�������D`���g�\A�Z +�L�&��\5�Q�T�mc���J��&
���m��tĿG��X����/ǐ�r��V�r���^��I�I�2�����J�7��%�޾Ѫݾ���G��T�/0�kG�%�\�J�p��؂��<���:���������Q�ÿB����1���������Y��8�Щ'�ѽ)��>�7b�\����a���5��?¿gÿP������5���(C��Mf��4:l���W�B�^�*���ht�'7�&pܾ�ᾠ`���~�1� ��7��bN��Mc�	rw�3�����������ĳ�S��KĿ�ܼ��r������[+v�`eL���0�CE&�ۍ.�އH�q�9������4b��6�ÿ0��@j��`~��蘕����4�y�Q�e��P�9d:��D#���0������n!ܾ ��K���6��](�q~?�'�U�� j��i~�ӊ�����)��ኸ�#�¿B�¿��������_���g��ZA�(+��&�S[5���T��b���I���	��Gm���Ŀ�ｿpX������Ɛ�#����r�z�^�I�
�2�����J�<��V�޾-�ݾ���%H�VU��0�G�ށ\��p�(ق�!=��9;��W���������ÿ�����2��a�����IY�:8�C�'�,�)�>�*8b�Ϙ��%b��66��8?¿�ÿq�����e���jC���f��;l���W�/B���*�F���u�
:�sܾ��Ac��2��Q� �
�7�tcN��Nc��rw�������������_ų�����Ŀ�ݼ�qs������H-v�ZgL���0�9G&���.���H��q���������b���  �  ���0����K%ɿ�⧿GK��i�i��'G���+���(V����jɾ?����U���?����;��辯m�ڶ�-h1�-N�|�r����������п�c�v���)�Φ���ݿ������np�m	P��J�o�^�Ap��x���JͿ����	���#����߿�ǽ�ޱ��$���*]�d=���#��������ؾ~�¾��c��F�����վC���O.!�J:��;Y�����o�����S�ۿY��]��������!tѿ���������b�$K��N�ǖk�����䳿|�ٿ3������ۤ�-n�}|Կ���&���Vw�I�Q�EM4��(���s�.aоe������������ƾ��޾���Κ��)���C�`e�Y���k��pXſ����) ��}��F����!�Ŀ�y���U�� �W��I�mU���z���������8��: �����/�����$ɿ�⧿�J��Īi��&G���+���U�����ɾ����S��I=��j�;!�辖l���bg1��N��r�������¹п�c�u���)�������ݿ9�����lp�&P�aJ��^��o��Nw��<JͿ�ￇ	���������߿*ǽ�}����#���)]��c=�r�#�������Ѳؾ��¾J��{c������V�վ�C����.!��J:��<Y�����p��>����ۿ�����\��� ��tѿ؏��a���_�b��	K�d
N��k�����e峿֜ٿq��������>n�|Կ9���K&��Ww� �Q�'N4��)�-�����cо���-�������,�ƾ�޾1���Л��)���C��`e����#l���Xſ/��.* ��}�G����!�Ŀ�z���V��$�W��I�wU�q�z�}��������8�-; ��  �  �0��)�+?�����o�ſ������n��X=�W�������3پn���k������<���$랾�u��%@¾���$���� �w�F�<N|�v����	ѿ���6���+���/��%�R��F�T@���9���u�%�m����y
��՞ӿl���?��,��H/�s�#�x5�-�{�������\�t(0��6����Y�ξ���ꣾ������������ʲ�Hg˾�0�u?��,�C�V�j������<�h�*�!�;�.���-�b�����
mٿs���ч�ko�� s��ߍ��1��iE��;�#��G/���,������ӴֿD;������L�xX$�ٝ�����/žOv������ޙ��<�������.�վ���bt���8��h��;��N���	��٢��~'���/�w*��Y�j���Kȿ΃��^���Kl�w�|����Q�¿�\������)��0��)��>�m���"�ſ\����n��W=���������1پJ���"���&��ѵ���螾@s���=¾���N��R� ���F��M|�i����	ѿ&���6���+���/��%��Q�NF��?��:9����u���m����	���ӿ���?���,�JH/�*�#�65�����A���\��'0�@6������ξ����ꣾ���ၚ�����=˲�0h˾2�@��,��V���� ��U=�gh���!���.�`�-�Ɉ�����mٿL����ч�
o�3"s�����Y2���E�H�X�#��G/���,�������ֿe;��殁��L�=Y$�Ğ���02ž�x��G��ᙾJ?��u��<��Q�վ���Su���8��h�_<��̌�����)���~'�F�/�xw*�nZ�k���Lȿ򄜿<_��9Nl���|����D�¿�]����=)��  �  (�Y��XP��7����'��*~���>�6����*¾�g���z�����Bć����"���֟��D�ɾ����k���J��Ї��䷿k�������1>���S��Y��)L�߸0��:� kڿ�(����������U���џ��;�����!��aA�yU��rX���I�P-�Y[
���ѿO]��gf�O.�����p۾ ���u��S���Έ�Hj��� ��]���e��g�־%{�nG)��_��4��,˿v��_)���F�M�W���V��QD��%�d���yǿ. ��h������Aޣ��ӿ�W
��-���I���X��[U��CA���!�����%���o��XQ�C��?��_�;�i��������ㇾډ�5��������k���k�P7��9��u�A9���߿�1�g;4�4FN��bY�p[R�[;�E���+￡�������>���3��R���s�6�q�7�*}P�߂Y�mXP�ܪ7����'�4�)~�J�>�r�߼�G¾�e���x��Ё�������������ם����ɾ^��k�8�J��Ї��䷿��������1>���S��Y��)L���0�z:�xjڿ!(��չ��؊���������q���_�!�oaA��xU�prX�W�I�-�[
�)�ѿ�\��wff��N.����mp۾Ø���t��S��ψ��j��2!���]���f����־�{�1H)�h_�u5���,˿Tv�$`)�!�F���W�!�V�-RD�Y�%�Ԭ��zǿ
!���h��S ���ޣ��ӿ�W
�$-���I��X��[U��CA���!�����%��#p���XQ�������M�;�k�����i���凾u܉�� ��4����m���m�D8��9��u��9����߿2��;4��FN�cY��[R��;�����,�է������k���U��e���r迪�׻7��}P��  �  ��w�a6m�V�P��@)�� �a
���^��NC���c⾻�c����&K����{����(������J���]&��CQ������)ɿ*D	��l2��$X�Pq�?w��@h��eH��7 �BB�b���<w��@u��	����Eֿ�T�J�6��[��s�"�v��^e��+D��g����R���q�O�0��W��Ѿ:2��D#��_���r}���|�����N���ҡ̾��p�*��h��t��:�߿?��;�?��Vb��u��|t��'_��m;����ݿI����t���u��܉��������(D��ke���v�� s�o�[���6�C����пe����X�=$ �f���`Vþ�颾Ib�����'�{� ]�O2������.��/Qܾ�w���<�v���GO�������$��L�z�j��w�po��lT�A�-�<���sɿ�{���s��Zy���ÿ���W)���P�)Em�Q�w�%6m�%�P�~@)�� �
���^��dMC�U�����ﶾg�ꗉ��H����{�轁�����������\�:&��CQ�z����)ɿ9D	� m2�%X�.Pq�?w��@h�beH�s7 ��A󿻉���v��wt��9����Dֿ T���6���[�ts�Ύv�t^e�h+D��g�B��􄧿sq�Њ0��W���Ѿ�1��#��_���lr}�f�|�l���	�����̾���5�*���h�au����߿�����?�Wb�P�u�}t��'_�&n;����ݿ+���}u��iv������/��B���(D��ke���v�� s�g�[���6�A����п����c�X��$ �����5Xþ�뢾xd��M�����{��a��4��F����0��,Sܾ�x���<���O��b�����$�v�L���j�[�w��po�rmT���-����7uɿ}��u���z���ÿr��qX)�I�P��Em��  �  25�`�-��`����!�¿���GjU����o�y+�� o��]݀�P�e�q�V�}�R�JY�J�j�:��D��	ľ�%��ʐ(�b�d�1����ο?�y����0��4�*�V���Pￚڹ�j	��ԉs��k��d��(����ֿz��=!�¸1�o;4�>(���dK�-�������@�-P�7�ھ��l�G�v���_�qT���S���]��s�2#������Ծ�
��R:��?}��Z��`��8����%�ϒ3�l�2�A�#���
�x�ܿ���6���ll��p�7���m�����8��t(��<4���1�C@!�Lk��,տLr��}l�LA.��~�Pɾ;o���F��r�m�*�Z�bS���U�ʝc���}�ce��썵�c�����AN��C������2�������+�s�4�{'/�.�+�Ƨʿ�՜���~��i�d�z�⯘���ĿO���&]�*�-��5�%�-�k`�§��إ¿G���iU�j��2n��)��Zm��rۀ�A�e�?�V�C�R�[FY�[�j�m���𝾞ľ�$����(�L�d�1����ο?������0��4�*�6��+P�ڹ����d�s�M k��c��X���I�ֿ�y�+=!�h�1�;4��(�Ү��J�� ��7���@��O�t�ھ<����v���_�wqT�F�S���]�[�s�$���K�Ծ��
��S:�z@}�E[����ῌ���%�0�3�ӽ2���#��
�[�ܿ�����6��Dnl�x�p�뉍����Y�d���(��<4���1�;@!�Dk��,տWr��M}l��A.�1��Qɾ�p���H����m���Z��S�x�U�-�c��}�jg��ۏ��>������BN�UD������x3����5�+���4��'/����+���ʿ�֜�F�~�}�i���z�������Ŀ:����]���-��  �  ��-�0x&�C?��>�;���=��ksQ��^�����������0���ebk�E\��(X���^��bp�FӇ��n���ž����ۡ&�g�_��і���ǿXi���T�;)�j:-�x!#����*�濶���挿�im�lCe��؀�������ο�H�����e*���,�M2!���
��߿聫�l��e�=�tq�uv۾x���x���d|��	e���Y�tY�p8c��y�����"0��͟վ\*
���7��^w��&��i�ٿ�')��#,�G]+�m��<� �Կ�"��}����f�k�j����Y���������:!���,��^*�����6���Ϳ-Λ�+mg��,�"��ʾ�ڣ�����s�	`��VX�aE[��i�W����	��8������;��_�J�6���.���D �;���$��|-��'�������C�ÿJ"���<x���c�.t�e/���>��J���D���&���-��w&�?��>�:��W=���rQ�@^�.��]���"��@���I^k��@\��$X�ğ^��^p�qч�m����ž������&�K�_��і���ǿi���T�);)�m:-�k!#�|��ƅ�0���o匿8hm��Ae��׀�������ο+H�L���e*�3�,�2!���
���߿~������͵=��p��u۾����x��Od|��	e��Y�+ Y��9c�< y��Ꮎ:1���վ+
�r�7��_w�'���ٿZ��)�%$,��]+���j=���Կ�#��[�����f���j�Ő��򴮿�����:!���,��^*�����6���Ϳ;Λ�omg�,��"���ʾFܣ�����!s�}`�![X��I[�<i�x������'������!��E�J���������� 쿍��e�$�`}-���'�,��)���r�ÿ#��e?x�D�c�`0t�z0���?��2��)E��&��  �  �?��&�`��-ٿ:<���6���G�Wp���`þ��G����|�I�l��kh�|ho����������˾k���o"��T�Xe��<���i�
����R���O��*����ο���:w���Q\�3U���m�׆��Fk���\�6"	�\��������t���ɿ����o�Ս6�+�
�߾x��.����L��}<v��j�:wi��Mt�`�������T��ӓھ~b	��=1��Wh��u�� YĿ?�������[��[l��`���l��$�r��aV���Y��$}�:���.~ɿHX����B��]}�		����|#��񥏿�Z�h0'��@���о�_���H�������p���h���k�x�z��늾 ���྾e �00���A�q�~��h��\�ӿx �&���*�rr����޿𼰿�1���e�D T�r9b�Ǉ����4�ؿB���2��?�O&�1���ٿ�;��~6��{�G��o�,�þ
�Gތ���|���l��gh�do� ��	�������˾U����n"�rT�Ye��P���i�����S���O��*���ο.���v���P\��1U�@�m�����j���[��!	������i��tt����ɿ����o�A�6�+�M�߾���Ӝ���L���<v��j��wi��Nt��������U���ھ=c	��>1�}Xh��v���YĿ�����G�3\�~�4m�a���m��׬r��cV�Q�Y�&}�Ь���~ɿ�X�� ��O��`}�	���迀#�����q�Z��0'�8A�Y�о�a���J��F���i�p�m�h���k���z��튾.��~⾾="�1���A�Y�~�qi����ӿmx ����C+��r�v��2޿����2��q�e��T��;b�'ȇ�����ؿ��� 3��  �  L`��:�,pٿ�����d���n���=��	�L���=�Ӿ�?��혞�Ͳ��3Z������`ۆ�骑�����G��Ϝ۾�L��? ��DG��~z��؜�����f�߿%�������Ul�=-ѿ ѭ�o����sb�H�C��=��Q�d�}��������aL����[���i���ο%;������t\�	10�]�.�-�Ⱦu笾����x؊������U��R���r���>M���žp�辥��� ,�Y�V��-���V���&˿x�� ����_���R忹�ſ���Ӂ�|U���>��A���]�'S��5ө�:pͿ��꿤F���D����ÿ����|���TL��	$���!�߾�n���\���C��]����ӂ�;����S��o���^����Ͼ���w���8���g�ξ������տ�#��D��U����ۿ�ٹ�����q��'K�j�<�$QH�%{l��Ғ��ֵ�T_ؿ����_���9��oٿq���od��� n���=�	�������Ӿ�=��Ԗ�������W��[���ن�����o���E��6�۾.L�J? �IDG�z~z��؜�����z�߿0�������2l��,ѿ�Э�𺋿�rb���C���=�t�Q��~}���������K�h��[���h�o�ο�:�������s\�y00����-��Ⱦ笾c���{؊�˶��)V��ڹ��'���"N���ž���a���,�J�V�t.���W��l'˿%��ڍ���`���S忋�ſb񡿗ԁ��}U�Z�>�d�A���]��S���ө��pͿ.���F���D���%�ÿˤ��*|��UL�8
$�a���߾�p��)_�� F��̻��Cւ������U�������`����Ͼ����V����8�m�g�E������S ֿr$�E��6����ۿ�ڹ�׀��H�q��)K���<�CSH�(}l��Ӓ�o׵�`ؿ���  �  ÿO���y���T��������3[�۬:�g� �F�����%rվ�ۻ�Z���N��;՘��E�����>����۾Ć��c(��&��FA�sc��b������籿�࿿��¿����B��A<���4e��H>��L'��#���1�'9R�d��w���ò��j���x�¿�E��]Ҧ��a��u��O�Oe1��^����U龢P̾#����o��k(��神�2���$Z��fɾ���(�����t.�\�K��~p��ڍ�Om������,¿���h۲�YY��^���ֻV��4�*�#�R�%��:��<`�[^��gա��ض��¿����
峿P����ڈ�Եg�>�D� �(��c�9V��߾�þ��Og�������y��i����[��UҾ�m𾥲	��F��7��7W�"O~��s���s��9L��ÿ�K������ړ���t���I���,��G"�K�*��E��o����F���^㻿�ÿ⟽�������R���O3[�;�:��� �x�����pվ�ٻ��W��CL���Ҙ�jC�������z�۾�����'�Q&�FA��rc��b������籿�࿿��¿�����~���;��4e��G>��K'�P #���1��7R����ȋ�����ˬ���¿TE���Ѧ�%a��Cu�N�O��d1�M^����U�MP̾�����o���(��J��������Z��gɾ���Ȕ����{u.�G�K��p�Hۍ��m��Ǖ���-¿У��,ܲ�#Z��+���o�V���4���#���%�L�:��=`��^���ա��ض�¿����峿d���ۈ�/�g���D���(��d�2X��F!߾��þ����i��" ��E|��ܞ���]��9WҾ�o𾎳	��G���7�a8W�P~�t��.t���L���ÿ�L������ۓ���t���I���,��I"�J�*��E�Ȇo����������㻿�  �  ڲ���C���؊��O����j��nW�ͶF��57�~9'���K{��辺y;i���L���f[����ҾC��[������*��:�rBJ��|[���o�Ă��ߌ�8/������S���z��cX�R�6��p��A��8���Pa)���H�P�k�v���@���_��T�����l9y�5	d���Q��A��1��!�\2����mW޾��ƾ�����׸�o�ľED۾����;����
<0�h�?��O���a���v��\��������1D��b@���o�v�L���,�b��v��r>
��
��3�fyT��&w���\���ޅ���э�������q��]�2L��[<��,�����N
����jվ����"巾2i���˾���5����2_%��z5���D�uU��h��&~�Sŉ�f����哿f���^���"d��ZA��l#�
A����-���� ���=��9`��〿ڦ��]���}C��/؊�8O��=�j�@nW�*�F��47��8'���5z�I�%w;���������X��ȦҾ����Z������*�1�:��AJ�2|[�V�o�Ă��ߌ�(/�����~S����z��bX�k�6��o��@�r7�����_)���H��k�����������T�������8y��d��Q���A���1�à!�2�����GW޾��ƾ(����׸���ľ�D۾g����;�J���<0�5�?� �O���a��v�z]��4������D��A��k�o���L�+�,������?
����3�IzT��'w�J����������э������q���]��L��\<��,����P
�0��Rmվ�����緾�k��X˾O��P����`%�Y{5�g�D��uU�ڈh��'~��ŉ������擿&���2����#d��\A��n#��B����
��p� �7�=�;`��䀿m����  �  ?�b�d�h���i��hi�oi�|�i���h�Ncb��UU��A��y*��,�����/�澔�߾���`��0%�d�/���F��X��Qd�.0i��i��Yi�Մi���i���g���`�{R�|>��z&����W���M��*��y�)�������3��
J��B[�ыe�%�i�x�i�8Pi��i�`�i�K1g�h�^�fsO�tF:��"��������R⾴I�1��4�	�v��Ӱ7�@VM�x]���f�ݶi�άi��Li�ٴi��i��Af���\��@L��b6�E������"������e���=���#�͍;��zP�;{_�Swg���i���i�sRi�T�i��hi��'e��yZ���H�Pr2�w�����\5��߾��%�����b�'��U?��rS�Ja�.h�'�i��|i�Y]i�9�i��i�x�c���W��jE��w.�L�����u���u߾õ�� �e���+�C��=V�V�b���h�(�i�5hi��ni���i��h��bb��TU��A��x*�r+�ː��;�澇�߾p��ܓ��#�
�/�i�F���X�Qd��/i���i�9Yi���i���i���g���`��zR��>�z&�9���U���K�r(�}w��������3��	J��A[�ϊe�7�i���i�xOi�b�i���i��0g��^�sO�8F:���"�������S�Jᾶ���	����V�7��VM��x]�e�f���i�íi��Mi���i�G�i�FCf���\��AL�Dd6����$��m%�S��_�⾶���>���#���;�7{P��{_��wg�F�i�&�i��Ri���i��ii��(e�{Z�:�H��s2�����o8��߾���
�������'��V?��sS��Ja��.h���i�K}i�!^i��i��i���c�;X�GlE�*y.��������ky߾7�羏� ��f��+��C��>V��  �  D8��G��nX���k�2퀿P^��7�������d�����eE^���;�	J���������$��8C�f��c���-��/���x`��9����|�~eg�c|T��D�2�4��q$��$�9��� �D�ɾ=庾���P����־c\��VJ�����-�a7=�9�L�4�^�� s�"����E��	����>��{_���Ou���R��n1�����	�p	�l��".�R�N��q����㝑��ޓ�H#��ƅ�Ҍu�Z�`�K�N���>�3Y/�d��?������پ�þ����󹾁�Ǿ��߾�n���-�
�"���2��]B���R�w%e�tz�R��ȱ��'�����������i�P�F��'�2��l�V��1���N8�YXZ���|�����7�������a��V'��tXn��tZ��\I�\�9�8�)�4 �Ua��>�=OѾ����񘷾�5��Q�ξ���q����#(�j8�S�G�.nX���k��쀿^��䅒��������P��'D^�4�;��H�N� ����`�$�37C��f�c���,������`���8���|�eg�|T�sD�М4�Hq$�$������^�ɾ(㺾��������־Z��7I�����-�o6=�Z�L�j�^�, s�Ҕ��{E��Ψ���>��T_��^Ou�\�R��n1����	��	����g".���N�g�q�`���9���ߓ��#���ƅ�ԍu�p�`�t�N���>�}Z/����s@�� ����پ͢þ����"�����Ǿ��߾ep��T.���"�|�2�^B�6�R��%e��tz����;������D������c�i���F���'�����������P8��YZ��|�}���8�����b���'��"Yn��uZ��]I�m�9�o�)����b��A�~RѾٛ��:����8��\�ξ���Nr����$(��  �  "�K<��:]�:���]A��xî�x=��bÿ%"���^��������l��C���)��`"��.���K���w�J���C��󽿾ÿʖ��8Q��*/�� �{�{CU� �5�����[��]�о�%���ɥ�������6��� ���(ž��
� �w���0*��sF���i��� Ġ��ڴ��1�������䵿<{��;���]��=9��>%��+$��"6�<Y�������
泿�������Ⲷ�+7������	Dn�EJ��-����U��5(�d�Ǿ@���M���r��}q��1���õ�1�;�뾙�����e�2��kQ��Pw��������������¿#��r����!��V}�YP�ؐ0��"��(�D@�L�g������ͥ�󃹿��¿�]���ిǛ�N)���Ya�)�?�f�$�o������5ھ.����������ǘ�w����=�����I׾�������J"�kJ<�-:]�����A��2î�%=���ÿ�!��3^���L�l���C��)��^"�.���K��w�:I��+C��p�(ÿN����P���.����{�CU���5�����$����о5$��ȥ������������y&ž���� �����/*�sF�!�i�����à�Yڴ�}1��y����䵿!{��)���]��=9�?%�,$�;#6��Y����C���U泿��N���L����7��r���En�dJ��-��������*�
�Ǿ�B��_P��u���s��53���ŵ���;>�@������2�lQ�LQw�ޥ��5 ��5���¿�#��8����"��	}�(P���0�м"�;(��@���g�$���8Υ�b���8�¿�]���ిIǛ��)���Za���?�Y�$�������8ھ����������ʘ�o��@��%"���׾����n���  �  ���'�?��q��<���鹿�ۿ#2�W�����/�ֿBճ�1����i�zG�P=�y�L�}�t��^���ڻ��{ݿi����!��8��>Կ���"�le�|�6�q���`����;����~}�������p��P3�����j���x�����ȉ�<�%���N��!��4����ſċ�G���������d�˿Dק�Q����[���@��e?�xW�|i���壿W�ǿ��濬�������h�Hɿwg��ez��U6T���)��z
�>R��[þ����ѕ��0��b,���탾�n��⃙�"<��mNʾ��խ��U2��G_��c��b.��u�п������Z��й�ֿ�i&���z���O�Nz=�ƣD�d�d�x��ѯ��ӿX�����/���Fc޿�ͽ������Ow�w�D��e����A�پ���T᡾x␾`p��֪��ϯ��xf��!���Z�����վ���������?�Dq��<��H鹿�ۿ�1�V���𿖜ֿ�Գ�g���i��G�a�<��L���t��]��ڻ�{ݿ���� !����i>ԿE�����e���6����h_����;(����{�������n��삾B1�����[���w����߈�c�%���N�4!��㍢��ſ����������m��J�˿3ק�J����[��@�f?�]xW��i���壿��ǿ�� �����Di�wHɿ�g���z��k7T��)��{
��T�h^þw
��Yԕ�3���.��<����p��΅���=���OʾR��u��{V2�RH_�d���.���п��쿶����[������ֿ�]'����z���O�-|=���D��d��x���ѯ�rӿǝ�?��u����c޿�ͽ�5����Pw�,�D��f������پ���� 䡾C吾:s����������!i������������վV����  �  ˟���J��7��+�����ۿ������;��������Zֿ|���)#���`��(T�<�g�S���� ��ɭ࿿���!���#����Jѿ���S�z�V�>�� �-<�tܼ�Ϧ�������ky��Rk��h�(�q��C���q����oӾ)��{�)��]�+Б�����<��
�u��S�M������ �ƿ	����cz���X�!W�'u�o�����*����׷���������)8����d�\�.���1ؾ�����Җ��΄��bs��1i�Gvj�!@w��+���훾]3�����G9��5s�TU���̿V���
x�*��9�u���忠�������%�k��T�B�]�����8���0ѿ2���{��=����.��Ɯ��O��>�P�J ����O�ɾ�������Ne��^�n�0Yh�Vlm�:,~�-����n��>1žs,�����J��7��򬭿x�ۿ�����V;�A��[���Yֿ����@"����`��&T�%�g�G������Ϭ�L�T���������rJѿ�����z���>�% �;�,ۼ�b���i���Jhy�=Ok�5�h�3�q��A���o��'���ӾI����)�A�]��ϑ�@������
�Z���R�;��o����ƿ����cz��X�3!W�P'u�Bo��H���h���� ����;��}�����8����d�{�.�F���ؾo���lՖ�ф��gs�S6i��zj�CDw�l-��<�︾���l�dH9�A6s��U��&̿����Vx����������忢�������,�k��T��]������8��q1ѿ������?�]����_������WO����P� �݄��i�ɾV���f����g��Ʒn��^h��qm�I1~��⍾ q��)3ž.���  �  6��h�T���������L�����8'���-�c�%�c��W��Z���8J���Sr��d��qz��/��	|ƿ������(�O`-���#��4�5�}���h���OG�2�_�侞W��P����Ӏ�ch��Z��X���`�g�t�c9��r����W;����.�lPk�]X��S�пk����E�*��~,�7: �ٙ	�B�ݿ&@�����8�i�yxg�?���4w����׿6��o ���+��+���e����ֿ�����Hs��4���{�Ҿ�I��쟍�ۋw��[b��X�dZ�Z�e�B~�)В�6$��\y޾�����@�U��&:���⿹j��)"��-���)�e���� ��̿�l���(��d���n�����N��.�鿓:�>$� b-���(�]�)b����Ŀ�_��D&\���#�s��-þ�Ğ�����+o��]�>X���\�D�l���������|N���������T��������OL��e���7'�X�-�!�%�����￀���HI���Qr��d�coz��.���zƿ���R���(��_-�o�#�V4���$����g���NG�v1�-��QV��☕�Ҁ��h�u�Z��{X��`���t�v7������V;�� �.��Ok�X���пI�� ��+�*�z~,�%: �̙	�2�ݿ@�����R�i��xg�_���^w����׿U��� ��+�1�+�������ֿ
����Is��4�����ҾFL��]�����w��`b���X��Z�qf�	~��ђ��%���z޾<����@�����:������j�	*"��-��)�ܐ�Y� ��̿�m���*��d�j�n������O��ن��:�u$�Ib-���(�t�Tb���Ŀ7`���&\���#�0��/þ�ƞ�h���Bo�Q�]�yX���\�+�l�䫄�����WP��d���  �  �q �Y�摓���ſ�������g.�95�*�,����`����¿X���b�x��i�-��������Ϳ���ok���/���4�+�4����ʳ��^牿��J��Z��6�zU����P|�a�b���U��@S� e[���n��s���?���̾:��z/1�ؒp�����Sؿ���Kw"�?2�|�3�l'��.�3�忹���;ߋ�rso�IQm������򬿑�߿�!�%�$��.3�>-3���$�7���޿������x�Y77�y��N�ѾE���^ߊ���q�_�\�S�S�V�T���`�yx����b��O�ݾA��pD��H���߳���뿸-��)�x}4��$1�6����i�ӿ�q�����Zwj�!u��ݒ�����]y��+���4���/�vn����˿�����`�0�%��W���z��~@��������i�K�X�3�R��xW�Ng�jہ�%�������)���p ��Y�����a�ſ��������f.�5���,�q�������¿f���Z�x���i��������ϓͿv���j�?�/�1�4��+�����o���牿�J�4Z�|5�+T��p1|��b���U��<S�Ja[� �n��q���=���	̾a���.1��p�e���Sؿ���-w"�?2�g�3�['��.�#�忳���>ߋ��so�vQm�������Ů߿�!�I�$�/3�k-3��$�n��޿w�����x�s87������Ѿ�����ኾi�q��\��S���T���`��|x�O�������ݾ��D�$I��೿���-��)��}4�D%1�������w�ӿ�r�����eyj�	#u��ޒ�ď��	z�`�J+��4���/��n�3��I�˿ĝ��}�`���%��Y���|���B��󃾞�i�t�X�_�R��}W�'g��݁�6��̍������  �  6��h�T���������L�����8'���-�c�%�c��W��Z���8J���Sr��d��qz��/��	|ƿ������(�O`-���#��4�5�}���h���OG�2�_�侞W��P����Ӏ�ch��Z��X���`�g�t�c9��r����W;����.�lPk�]X��S�пk����E�*��~,�7: �ٙ	�B�ݿ&@�����8�i�yxg�?���4w����׿6��o ���+��+���e����ֿ�����Hs��4���{�Ҿ�I��쟍�ۋw��[b��X�dZ�Z�e�B~�)В�6$��\y޾�����@�U��&:���⿹j��)"��-���)�e���� ��̿�l���(��d���n�����N��.�鿓:�>$� b-���(�]�)b����Ŀ�_��D&\���#�s��-þ�Ğ�����+o��]�>X���\�D�l���������|N���������T��������OL��e���7'�X�-�!�%�����￀���HI���Qr��d�coz��.���zƿ���R���(��_-�o�#�V4���$����g���NG�v1�-��QV��☕�Ҁ��h�u�Z��{X��`���t�v7������V;�� �.��Ok�X���пI�� ��+�*�z~,�%: �̙	�2�ݿ@�����R�i��xg�_���^w����׿U��� ��+�1�+�������ֿ
����Is��4�����ҾFL��]�����w��`b���X��Z�qf�	~��ђ��%���z޾<����@�����:������j�	*"��-��)�ܐ�Y� ��̿�m���*��d�j�n������O��ن��:�u$�Ib-���(�t�Tb���Ŀ7`���&\���#�0��/þ�ƞ�h���Bo�Q�]�yX���\�+�l�䫄�����WP��d���  �  ˟���J��7��+�����ۿ������;��������Zֿ|���)#���`��(T�<�g�S���� ��ɭ࿿���!���#����Jѿ���S�z�V�>�� �-<�tܼ�Ϧ�������ky��Rk��h�(�q��C���q����oӾ)��{�)��]�+Б�����<��
�u��S�M������ �ƿ	����cz���X�!W�'u�o�����*����׷���������)8����d�\�.���1ؾ�����Җ��΄��bs��1i�Gvj�!@w��+���훾]3�����G9��5s�TU���̿V���
x�*��9�u���忠�������%�k��T�B�]�����8���0ѿ2���{��=����.��Ɯ��O��>�P�J ����O�ɾ�������Ne��^�n�0Yh�Vlm�:,~�-����n��>1žs,�����J��7��򬭿x�ۿ�����V;�A��[���Yֿ����@"����`��&T�%�g�G������Ϭ�L�T���������rJѿ�����z���>�% �;�,ۼ�b���i���Jhy�=Ok�5�h�3�q��A���o��'���ӾI����)�A�]��ϑ�@������
�Z���R�;��o����ƿ����cz��X�3!W�P'u�Bo��H���h���� ����;��}�����8����d�{�.�F���ؾo���lՖ�ф��gs�S6i��zj�CDw�l-��<�︾���l�dH9�A6s��U��&̿����Vx����������忢�������,�k��T��]������8��q1ѿ������?�]����_������WO����P� �݄��i�ɾV���f����g��Ʒn��^h��qm�I1~��⍾ q��)3ž.���  �  ���'�?��q��<���鹿�ۿ#2�W�����/�ֿBճ�1����i�zG�P=�y�L�}�t��^���ڻ��{ݿi����!��8��>Կ���"�le�|�6�q���`����;����~}�������p��P3�����j���x�����ȉ�<�%���N��!��4����ſċ�G���������d�˿Dק�Q����[���@��e?�xW�|i���壿W�ǿ��濬�������h�Hɿwg��ez��U6T���)��z
�>R��[þ����ѕ��0��b,���탾�n��⃙�"<��mNʾ��խ��U2��G_��c��b.��u�п������Z��й�ֿ�i&���z���O�Nz=�ƣD�d�d�x��ѯ��ӿX�����/���Fc޿�ͽ������Ow�w�D��e����A�پ���T᡾x␾`p��֪��ϯ��xf��!���Z�����վ���������?�Dq��<��H鹿�ۿ�1�V���𿖜ֿ�Գ�g���i��G�a�<��L���t��]��ڻ�{ݿ���� !����i>ԿE�����e���6����h_����;(����{�������n��삾B1�����[���w����߈�c�%���N�4!��㍢��ſ����������m��J�˿3ק�J����[��@�f?�]xW��i���壿��ǿ�� �����Di�wHɿ�g���z��k7T��)��{
��T�h^þw
��Yԕ�3���.��<����p��΅���=���OʾR��u��{V2�RH_�d���.���п��쿶����[������ֿ�]'����z���O�-|=���D��d��x���ѯ�rӿǝ�?��u����c޿�ͽ�5����Pw�,�D��f������پ���� 䡾C吾:s����������!i������������վV����  �  "�K<��:]�:���]A��xî�x=��bÿ%"���^��������l��C���)��`"��.���K���w�J���C��󽿾ÿʖ��8Q��*/�� �{�{CU� �5�����[��]�о�%���ɥ�������6��� ���(ž��
� �w���0*��sF���i��� Ġ��ڴ��1�������䵿<{��;���]��=9��>%��+$��"6�<Y�������
泿�������Ⲷ�+7������	Dn�EJ��-����U��5(�d�Ǿ@���M���r��}q��1���õ�1�;�뾙�����e�2��kQ��Pw��������������¿#��r����!��V}�YP�ؐ0��"��(�D@�L�g������ͥ�󃹿��¿�]���ిǛ�N)���Ya�)�?�f�$�o������5ھ.����������ǘ�w����=�����I׾�������J"�kJ<�-:]�����A��2î�%=���ÿ�!��3^���L�l���C��)��^"�.���K��w�:I��+C��p�(ÿN����P���.����{�CU���5�����$����о5$��ȥ������������y&ž���� �����/*�sF�!�i�����à�Yڴ�}1��y����䵿!{��)���]��=9�?%�,$�;#6��Y����C���U泿��N���L����7��r���En�dJ��-��������*�
�Ǿ�B��_P��u���s��53���ŵ���;>�@������2�lQ�LQw�ޥ��5 ��5���¿�#��8����"��	}�(P���0�м"�;(��@���g�$���8Υ�b���8�¿�]���ిIǛ��)���Za���?�Y�$�������8ھ����������ʘ�o��@��%"���׾����n���  �  D8��G��nX���k�2퀿P^��7�������d�����eE^���;�	J���������$��8C�f��c���-��/���x`��9����|�~eg�c|T��D�2�4��q$��$�9��� �D�ɾ=庾���P����־c\��VJ�����-�a7=�9�L�4�^�� s�"����E��	����>��{_���Ou���R��n1�����	�p	�l��".�R�N��q����㝑��ޓ�H#��ƅ�Ҍu�Z�`�K�N���>�3Y/�d��?������پ�þ����󹾁�Ǿ��߾�n���-�
�"���2��]B���R�w%e�tz�R��ȱ��'�����������i�P�F��'�2��l�V��1���N8�YXZ���|�����7�������a��V'��tXn��tZ��\I�\�9�8�)�4 �Ua��>�=OѾ����񘷾�5��Q�ξ���q����#(�j8�S�G�.nX���k��쀿^��䅒��������P��'D^�4�;��H�N� ����`�$�37C��f�c���,������`���8���|�eg�|T�sD�М4�Hq$�$������^�ɾ(㺾��������־Z��7I�����-�o6=�Z�L�j�^�, s�Ҕ��{E��Ψ���>��T_��^Ou�\�R��n1����	��	����g".���N�g�q�`���9���ߓ��#���ƅ�ԍu�p�`�t�N���>�}Z/����s@�� ����پ͢þ����"�����Ǿ��߾ep��T.���"�|�2�^B�6�R��%e��tz����;������D������c�i���F���'�����������P8��YZ��|�}���8�����b���'��"Yn��uZ��]I�m�9�o�)����b��A�~RѾٛ��:����8��\�ξ���Nr����$(��  �  ?�b�d�h���i��hi�oi�|�i���h�Ncb��UU��A��y*��,�����/�澔�߾���`��0%�d�/���F��X��Qd�.0i��i��Yi�Մi���i���g���`�{R�|>��z&����W���M��*��y�)�������3��
J��B[�ыe�%�i�x�i�8Pi��i�`�i�K1g�h�^�fsO�tF:��"��������R⾴I�1��4�	�v��Ӱ7�@VM�x]���f�ݶi�άi��Li�ٴi��i��Af���\��@L��b6�E������"������e���=���#�͍;��zP�;{_�Swg���i���i�sRi�T�i��hi��'e��yZ���H�Pr2�w�����\5��߾��%�����b�'��U?��rS�Ja�.h�'�i��|i�Y]i�9�i��i�x�c���W��jE��w.�L�����u���u߾õ�� �e���+�C��=V�V�b���h�(�i�5hi��ni���i��h��bb��TU��A��x*�r+�ː��;�澇�߾p��ܓ��#�
�/�i�F���X�Qd��/i���i�9Yi���i���i���g���`��zR��>�z&�9���U���K�r(�}w��������3��	J��A[�ϊe�7�i���i�xOi�b�i���i��0g��^�sO�8F:���"�������S�Jᾶ���	����V�7��VM��x]�e�f���i�íi��Mi���i�G�i�FCf���\��AL�Dd6����$��m%�S��_�⾶���>���#���;�7{P��{_��wg�F�i�&�i��Ri���i��ii��(e�{Z�:�H��s2�����o8��߾���
�������'��V?��sS��Ja��.h���i�K}i�!^i��i��i���c�;X�GlE�*y.��������ky߾7�羏� ��f��+��C��>V��  �  ڲ���C���؊��O����j��nW�ͶF��57�~9'���K{��辺y;i���L���f[����ҾC��[������*��:�rBJ��|[���o�Ă��ߌ�8/������S���z��cX�R�6��p��A��8���Pa)���H�P�k�v���@���_��T�����l9y�5	d���Q��A��1��!�\2����mW޾��ƾ�����׸�o�ľED۾����;����
<0�h�?��O���a���v��\��������1D��b@���o�v�L���,�b��v��r>
��
��3�fyT��&w���\���ޅ���э�������q��]�2L��[<��,�����N
����jվ����"巾2i���˾���5����2_%��z5���D�uU��h��&~�Sŉ�f����哿f���^���"d��ZA��l#�
A����-���� ���=��9`��〿ڦ��]���}C��/؊�8O��=�j�@nW�*�F��47��8'���5z�I�%w;���������X��ȦҾ����Z������*�1�:��AJ�2|[�V�o�Ă��ߌ�(/�����~S����z��bX�k�6��o��@�r7�����_)���H��k�����������T�������8y��d��Q���A���1�à!�2�����GW޾��ƾ(����׸���ľ�D۾g����;�J���<0�5�?� �O���a��v�z]��4������D��A��k�o���L�+�,������?
����3�IzT��'w�J����������э������q���]��L��\<��,����P
�0��Rmվ�����緾�k��X˾O��P����`%�Y{5�g�D��uU�ڈh��'~��ŉ������擿&���2����#d��\A��n#��B����
��p� �7�=�;`��䀿m����  �  ÿO���y���T��������3[�۬:�g� �F�����%rվ�ۻ�Z���N��;՘��E�����>����۾Ć��c(��&��FA�sc��b������籿�࿿��¿����B��A<���4e��H>��L'��#���1�'9R�d��w���ò��j���x�¿�E��]Ҧ��a��u��O�Oe1��^����U龢P̾#����o��k(��神�2���$Z��fɾ���(�����t.�\�K��~p��ڍ�Om������,¿���h۲�YY��^���ֻV��4�*�#�R�%��:��<`�[^��gա��ض��¿����
峿P����ڈ�Եg�>�D� �(��c�9V��߾�þ��Og�������y��i����[��UҾ�m𾥲	��F��7��7W�"O~��s���s��9L��ÿ�K������ړ���t���I���,��G"�K�*��E��o����F���^㻿�ÿ⟽�������R���O3[�;�:��� �x�����pվ�ٻ��W��CL���Ҙ�jC�������z�۾�����'�Q&�FA��rc��b������籿�࿿��¿�����~���;��4e��G>��K'�P #���1��7R����ȋ�����ˬ���¿TE���Ѧ�%a��Cu�N�O��d1�M^����U�MP̾�����o���(��J��������Z��gɾ���Ȕ����{u.�G�K��p�Hۍ��m��Ǖ���-¿У��,ܲ�#Z��+���o�V���4���#���%�L�:��=`��^���ա��ض�¿����峿d���ۈ�/�g���D���(��d�2X��F!߾��þ����i��" ��E|��ܞ���]��9WҾ�o𾎳	��G���7�a8W�P~�t��.t���L���ÿ�L������ۓ���t���I���,��I"�J�*��E�Ȇo����������㻿�  �  L`��:�,pٿ�����d���n���=��	�L���=�Ӿ�?��혞�Ͳ��3Z������`ۆ�骑�����G��Ϝ۾�L��? ��DG��~z��؜�����f�߿%�������Ul�=-ѿ ѭ�o����sb�H�C��=��Q�d�}��������aL����[���i���ο%;������t\�	10�]�.�-�Ⱦu笾����x؊������U��R���r���>M���žp�辥��� ,�Y�V��-���V���&˿x�� ����_���R忹�ſ���Ӂ�|U���>��A���]�'S��5ө�:pͿ��꿤F���D����ÿ����|���TL��	$���!�߾�n���\���C��]����ӂ�;����S��o���^����Ͼ���w���8���g�ξ������տ�#��D��U����ۿ�ٹ�����q��'K�j�<�$QH�%{l��Ғ��ֵ�T_ؿ����_���9��oٿq���od��� n���=�	�������Ӿ�=��Ԗ�������W��[���ن�����o���E��6�۾.L�J? �IDG�z~z��؜�����z�߿0�������2l��,ѿ�Э�𺋿�rb���C���=�t�Q��~}���������K�h��[���h�o�ο�:�������s\�y00����-��Ⱦ笾c���{؊�˶��)V��ڹ��'���"N���ž���a���,�J�V�t.���W��l'˿%��ڍ���`���S忋�ſb񡿗ԁ��}U�Z�>�d�A���]��S���ө��pͿ.���F���D���%�ÿˤ��*|��UL�8
$�a���߾�p��)_�� F��̻��Cւ������U�������`����Ͼ����V����8�m�g�E������S ֿr$�E��6����ۿ�ڹ�׀��H�q��)K���<�CSH�(}l��Ӓ�o׵�`ؿ���  �  �?��&�`��-ٿ:<���6���G�Wp���`þ��G����|�I�l��kh�|ho����������˾k���o"��T�Xe��<���i�
����R���O��*����ο���:w���Q\�3U���m�׆��Fk���\�6"	�\��������t���ɿ����o�Ս6�+�
�߾x��.����L��}<v��j�:wi��Mt�`�������T��ӓھ~b	��=1��Wh��u�� YĿ?�������[��[l��`���l��$�r��aV���Y��$}�:���.~ɿHX����B��]}�		����|#��񥏿�Z�h0'��@���о�_���H�������p���h���k�x�z��늾 ���྾e �00���A�q�~��h��\�ӿx �&���*�rr����޿𼰿�1���e�D T�r9b�Ǉ����4�ؿB���2��?�O&�1���ٿ�;��~6��{�G��o�,�þ
�Gތ���|���l��gh�do� ��	�������˾U����n"�rT�Ye��P���i�����S���O��*���ο.���v���P\��1U�@�m�����j���[��!	������i��tt����ɿ����o�A�6�+�M�߾���Ӝ���L���<v��j��wi��Nt��������U���ھ=c	��>1�}Xh��v���YĿ�����G�3\�~�4m�a���m��׬r��cV�Q�Y�&}�Ь���~ɿ�X�� ��O��`}�	���迀#�����q�Z��0'�8A�Y�о�a���J��F���i�p�m�h���k���z��튾.��~⾾="�1���A�Y�~�qi����ӿmx ����C+��r�v��2޿����2��q�e��T��;b�'ȇ�����ؿ��� 3��  �  ��-�0x&�C?��>�;���=��ksQ��^�����������0���ebk�E\��(X���^��bp�FӇ��n���ž����ۡ&�g�_��і���ǿXi���T�;)�j:-�x!#����*�濶���挿�im�lCe��؀�������ο�H�����e*���,�M2!���
��߿聫�l��e�=�tq�uv۾x���x���d|��	e���Y�tY�p8c��y�����"0��͟վ\*
���7��^w��&��i�ٿ�')��#,�G]+�m��<� �Կ�"��}����f�k�j����Y���������:!���,��^*�����6���Ϳ-Λ�+mg��,�"��ʾ�ڣ�����s�	`��VX�aE[��i�W����	��8������;��_�J�6���.���D �;���$��|-��'�������C�ÿJ"���<x���c�.t�e/���>��J���D���&���-��w&�?��>�:��W=���rQ�@^�.��]���"��@���I^k��@\��$X�ğ^��^p�qч�m����ž������&�K�_��і���ǿi���T�);)�m:-�k!#�|��ƅ�0���o匿8hm��Ae��׀�������ο+H�L���e*�3�,�2!���
���߿~������͵=��p��u۾����x��Od|��	e��Y�+ Y��9c�< y��Ꮎ:1���վ+
�r�7��_w�'���ٿZ��)�%$,��]+���j=���Կ�#��[�����f���j�Ő��򴮿�����:!���,��^*�����6���Ϳ;Λ�omg�,��"���ʾFܣ�����!s�}`�![X��I[�<i�x������'������!��E�J���������� 쿍��e�$�`}-���'�,��)���r�ÿ#��e?x�D�c�`0t�z0���?��2��)E��&��  �  A��]�濞οw��$?��$[S�{L ������7m���gv��S��P>���2�R�/���4�v*B�'FZ�'���˜�˾ƾ-O�]�*�Dm`�搿uN��3�Կ>꿉6�}O�+ǿc1��Hf��&�U���7��L2�'�E���o����j��z�׿�����߿9tÿ�����H|��@���l�޾􈭾�~��,i�7jK� n9��0��I0�G8�[�H��)e�sv��E��huؾ���;�u�ޡ������c@ݿ���}�쿑�ڿ�/���ř�i�u��&I�d83�^�5��9Q����[����ÿB�߿�����׿-��|Ȕ�2/g��/�,K�nk̾ѷ���˂���]�DD�:�5�c�/���1���<�J�P��q�E���I���[�j��M�&}��������ʿW�����!z��aѿ����Ď���d�x+?�F]1�7m<�v[_��:��笿�ο?�濳����@ο�v���>���ZS��K ����a
���k��(dv�S�S��L>���2�2�/��4��&B��BZ�%���ʜ��ƾ�N�B�*�Sm`�#搿�N��U�ԿT꿉6�_O��*ǿ 1���e���U�R�7�OK2���E�L�o���Ji����׿��t���߿�sÿ2���H|�V�@�]�|�޾8���M~��Z+i��iK�n9�C�0��J0�T	8���H�a+e��w������vؾ���;�+u�s���o¿�Aݿz��E��c�ڿ_0���ƙ�%�u��(I�:3���5��:Q�y���[����ÿy�߿�����׿
-��|Ȕ�N/g�R�/��K��l̾@���{͂���]�7HD���5�Ŵ/�,�1��<�p�P��q�(�����e]��j��M��}��K���2�ʿ�俒��{��bѿð�CŎ�
�d��-?��_1�to<��]_��;���笿�ο���  �  �����ݿ��ƿ����kJ��{N�S��)���L���ᖾ�tz��>X�1�B�E�6�L�3�u�8�F�}�^���u��Ȟƾ� �%�'�t�Z�����q2����̿�H�a!�}�ٿ����ş�	����&P�y�3��A.��@�ti�nX�����غϿ8����/�׿����y���tu�/�<�c.�P�ݾ�F��"3��gm��O��=���4��c4�}B<�SDM��oi�Y<��9�����׾���[Q7��n�����'���տ�����㿪}ҿG����䔿��n��(D��#/���1���K�F�z�1��������׿��>��٭Ͽ�ޱ��A��_a�c�,�L��b̾'ۡ������b�$�H��9��3�6�b�@��DU���u�����n����꾥�LwH�����9���Zÿ|�ۿVr�Q�߿��ɿ
Ȫ�Mf��%j^���:��[-�s�7�)jY�m�����ʪƿ��ݿ�濁�ݿ@�ƿ<���#J���zN������`K��_���0qz��:X�-�B��6��3�]�8��|F��^����1��֝ƾ@ ��'��Z�Đ���2����̿�H�_!�^�ٿh��^ş������%P��3�E@.���@��i��W��;���Ͽ���R�応�׿����x��tu���<��-�a�ݾ�E���2��cfm���O��=��4�Pd4��C<��EM�Qqi�j=��|���k�׾���LR7��n��������Gտf�俶��{~ҿ����唿D�n��*D�G%/��1�E�K�o�z����宼���׿;��E��խϿ�ޱ��A��3_a���,�����̾�ܡ�����tb�K�H�d�9�{�3�r6���@�(IU���u�񄓾Pp����꾂�0xH���������Zÿ0�ۿ%s�9�߿��ɿɪ�ng��vl^��:�9^-���7�ClY�f�������ƿA�ݿ�  �  ��ͿS�ƿ,����k��
�u��A�E{��0����_��a��bnf��6P�+�C�DS@�B�E�=DT���l�0ň������Ǿ?����  ���L���}ȝ��㷿�eɿƇͿ,ÿoج��Ȋk���@�Ԗ'���"�,3���V�m������K��L�ʿ�Ϳ������ƍ�Sbc�Ǎ2�B����ܾⱾP���w{���]��K���A�!A�_�I��A[���w�:�����+!׾���6�-���]�)�����������h̿[�˿8���Aأ�������[�$76�2�#��&��=�:f�vō�l穿�
��Ϳ��ʿ^���렿 ,���R��s$��� ���̾ׄ���?��'Bp��uV���F��x@�!�B��YN��kc�^����:���1��b辏g�x�<��eo�6���د��Ŀ�Ϳ�ȿc3���u����|��HM���-�Y"��w+���H���v��I��r���+�ƿH�Ϳ�ƿϞ���k��z�u���A��z��/���s]�����yjf��2P�߽C��N@���E�+@T���l��È������Ǿ�����  ���L�#���ȝ��㷿�eɿ��Ϳÿ.ج�~ˉk���@�~�'�=�"��*3��V�Yl��W���'K����ʿͿv��p��2ƍ��ac��2����ܾ͗f᱾�O��w{�;�]��K���A��!A�k�I�C[�P�w�J�������"׾���$�-��]�����{�������i̿�˿���٣�w�����[��86�ȭ#�F&�=�^f��ō��穿�
��(Ϳ��ʿ^���렿),���R�	t$�� �%�̾d���hA��,Fp�DzV�"�F�\}@���B�a^N�-pc�b⁾�<��h3���ih�W�<��fo��6��ٯ���Ŀ��Ϳ�ȿ[4���v����|��JM���-��"��y+���H���v�{J��3���Їƿ�  �  �g��<ꦿ|̗�\���CZ��I2��.�>���
Ǿ�慨����趀�>i���Z���V�"]�j�m����e���򮾒�ξ����D���:�q�c��퇿�͛�6�����_ţ��V��Ԋx�D#M�]�*���7�����O<���d��̈�뜿ù��ѫ��Ƣ�+I��	iw�XJL�n&����++ྥ����������5x�9c��VX�X�W��a� bu������������۾���֧"�L�G��|r�� ��-��mU��N���Ȟ�>����i�0P@�`�!���������'���H�P�s����Q7��糫���������sR���h�S�>��d��T���Ӿ���혾�߅��p��s^�w�V��Y��g��7~�}ŏ����PFþ���W��*>.�/�U�����߯������Y������阿҃���Z�Q�4������:��,1�	AV�UO��oʖ�:���Zg���馿 ̗���CZ�I2�G.���N	Ǿ�����۴���i���Z�*�V�x]��m����������\�ξ��������:�w�c��͛�;�����9ţ��V���x�O"M�:�*���T6�N��&N<�6�d��ˈ�iꜿ ���qЫ�nƢ��H��+hw��IL�em&���G*�����������I5x�9c�
WX��W��a�ccu�գ����T�����۾�����"�Q�G��}r�����-��!V������Ȟ��>��S�i��Q@���!�R��b����'�ܽH�9�s�����7�������������~R���h���>�.e��U��b	Ӿ����	ⅾ�p��x^�BW���Y��g�T<~��Ǐ����HþO��,��?.��U�/���o�������bZ����꘿|Ӄ���Z�u�4�"!���-<��.1��BV�'P��(˖�ه���  �  ?ɉ������y��N^��6A��r&����Wi���t۾��������������~�>�x��|��Z⊾+���/���}ƾ�����u��,���G�\�d�@�~�v�<n�����jl�K�K�x+�7_���e��������	=��^^�h�{�􈇿撉��g	q�8�T���7�j�&0	�̀�s-Ҿ.ݸ����J���^����z�Z	z��H�������頾FD��X.Ͼ� ��a��;�4�LQ��n��悿�M���&��%�~�P�a���@�d�!���
�'��� � ���a)(�7H��i��恿���m}��������g�o�J���.���� �N5�dVɾ05��i����a���U���y��|�����Mܔ������-��dNؾ����1���#��>�[�`�v��ǅ��ω�q���v�W�:�5������С���*�`��M2�DOS���r�l���ȉ�����H�y�EN^�L6A�Lr&����g��s۾����!�軖�x�� ~�E�x�ez���ߊ��)���_{ƾ5�ᾈ�iu��,�j�G�X�d�@�~�o�'n�����ljl���K�.w+�"^����ɞ�����H���=�i]^� �{�Z���V���Dyq�e�T�"�7�si��/	����,Ҿ�ܸ����lJ���^��J�z�
z�)I��d���l꠾PE���/Ͼ2���E��9�4�+MQ��	n�H炿�N���'����~���a���@���!�x�
����~� ��t*(�H��i�灿����}��ɢ���g���J���.�������6�HXɾT7������ud��vX���y���|�VĆ��ޔ�ٟ��}/��.Pؾ,��������#��>�[�l�v�Aȅ��Љ�8���v��W�-�5������ҥ���,��a��O2��PS��r����  �  ҴW���V���M�5@�r�1��v$��u�	��4�55��yϾ0w��i񣾤���*ߓ��������������#վ���D��˔��
��N'�x�4��]C�6P�a�W�;�V�F-L�d�9��_"��N��$�%�ھ�U־�徿:�����/���D�I-S��VX�V@T�1iI� e;�7-��U �����+	�d)��ڗ�i%ǾQ���垾B�������g��&��rmľ��ݾ�^�����__����ٴ+��9���G�PS��NX�C:T���F�s2�r��d����o	׾�)پ��������7�tJ�&�U���W�u7Q���D��6�_�(�X�w���;�ھ���׾����ũ����F	��Q���
)�������̾�U����~���-�u#��F0�N�>�8L�^�U�{X�n�P��r@��N*�����7��*�6�վJ޾�X���0���'�;4>�LNO��W��V��M�y4@���1�Qv$�5u�Q��3�R3��wϾ�t����}��tܓ�牙����z����!վ���k����
�WN'�B�4��]C�P�<�W���V��,L�ل9�*_"��M�v"�ܒھ�S־]��s9�k��̄/�p�D�&,S��UX�^?T�QhI�8d;�a6-��T �}���+	��(��`��%Ǿ�P���垾3B�����dh�����Knľ��ݾ `��{��&`����е+��9���G�VQS�'PX��;T���F��2��s�`f���:׾P,پc����j��Y7��tJ���U���W��7Q�C�D�_�6���(��X�9���<����]�׾%��Eȩ�ۻ���������+�����۬̾|W澪���M���.�3#�eG0�'�>�9L�x�U��	X�ܶP�Rt@�7P*�̵�];���-��վ�޾\��X2��'��5>�iOO��  �  b�*�.�/��1��1�� 1��0��a/��m*�� ��9��|��Ⱦ�'������5��^Sξ��r��{�Wq#���+���/�Y1�1�2#1�F�0���.�W,)�i���}�.���a߾�+žU_��ie��ꬼ���ҾG��Y<	�_��_.%�I�,��N0�S 1�1�h$1��0�[/.�#�'����L���'��>rھĸ��X򳾏3��0���"D׾q�����<=��&�d�-��0�##1��1�>"1��|0�l-�0C&��x���f���Ĵվ����Ⲿ
`���¾�ܾ$��j��:w�9C(��i.���0�+$1�u1��1�l30���,���$����M���\1Ѿ�û��2���굾`ƾ�ᾟ� �D^������)��/���0��!1�.1��1�$�/�ӌ+�D�"�,��(�����@�̾�G��iⱾѷ�
5ʾ�5�8��D����!��*�n�/��1��1��1�t�0�Fa/��l*�>� �����y�K�Ⱦ%����;��sPξ!���p��z�Zp#���+��/��1��1��"1��0���.�,)����<}�����Y_߾�)ž-]��c�������Ҿ���,;	�>��N-%�K�,��M0��1�U1��#1�Q�0��..���'�C����Q'��rھ˸�����3�������D׾�q��}���=���&�'�-���0�$1��1�X#1�~0�Hm-��D&�z�^�>�����վՖ��2岾�b��L�¾�ܾ���!���w��C(�:j.���0��$1��1�T1�$40���,� �$�!�;O���M4Ѿ�ƻ��5�����bƾN��� �E_����K�)�o/���0�~"1��1��1�#�/���+���"��������龯�̾2K���屾tԷ�>8ʾ�8澓��x��˒!��  �  n��.�+%���2�� A�K4N���V��~W��N��=�IZ&�����|��� ݾ��վ2N��:��'���+���A��_Q�v(X�~U�a�K���=���/�`a"������%O�����=H˾�ҳ��P��cA��-���\���Ҫ�Sm���kپ�)�����z�g ��|)��`7�G�E���Q�PX�{�U��I���5�5f�;��7쾾�ؾ�|׾�-�8������Y3�G�G���T��@X�6�R�2G�T�8���*��Q�?���5�~���Gܾ�þW���`���΃��a�������w����Ⱦ8������	�'F��!�X�-��2<�� J�O�T�NX��R���C��9.����*�~���־]۾S�򾧁�x�#�a�:�3�L���V�|VW�OtO���B��04�N�&��c�]���:�|��Ӿ9����������Г����ڤ�����,�оS��F�����z�s*%�i�2� A��3N���V�~W�7�N�s=�Y&�f���y���ݾx�վ�Jᾘ7�������+�9�A�s^Q��'X�U}U�ǈK�M�=�R�/�a"�6��C�7N������F˾ѳ�$O��Z?���*���Z���Ъ�k���iپ�'�����y�����{)��_7���E�N�Q��X��U�ӍI���5�f�+���7��ؾ�|׾).龍��H��Z3�ۯG�5�T��AX�
�R� 3G�P�8���*�S�t���6�����Iܾ�þ
������X���Đ��ʮ���x��D�Ⱦ��P���g�	��F�l!���-�b3<��!J�%�T�OX��R��C�R;.�x��=,����־`۾3�������#�h�:� M���V�'WW��tO�3�B��14��&��d�c���;��~��Ӿ<���Ħ�R���ԓ�<���ݤ�c�����о���?���  �  pK�������'��B���_���z�"������u���^q��sQ�Œ0��l��G���f��v�w�7��X�_�w��m���ʉ��Y��gu�rY�փ<�_"�Jp�`�����־�ּ��y�����#���8|��;y�!́�#+��Ժ��bv��c�ʾf�������j0�~mL�Hni��9������ 爿�K��zFg��@F�2�&����sX ��8�����_#�*�B�q�c����^m���"���[��X�l���O�%_3�����
�
G��;`���7՟�9Î��Â�(�y�<6{���(��6���,��ȰӾlF�@B
���m9�0V�7�r��l��Q����/��H�z�Q�\�-6;�R�X��?���J�9���%-�w�M�Gn�����>�������ً}��c���E���*��E�� ��Cྛžk���ͥ���$�����a�x�%�~�����ΰ��u ���G¾N
ݾ�I��P���'���B��_�K�z��􆿨��������\q�RrQ�R�0����������Pd��t�ś7�i�X��w��l��ʉ�Y��Nfu�xqY�_�<��^"��o�������־|ռ�cx��H�/"���4|��7y�ˁ��(������Nt��d�ʾ���� ���j0��lL��mi��9��X����房�K��DFg��@F�$�&�����X �&9����e_#���B���c����m��P#��Z\��:�l���O�-`3������xI꾇�;�����ן��Ŏ�5Ƃ��y��:{�򄾳*���7��Z.���Ӿ�G��B
�����m9��0V� �r�Km��᫉��0����z��\��7;��S��eC��-L�����&-���M�Tn�������������f�}�* c�/�E�M�*��F�| ��E��ž
��������'�����R�x��~�i���b����"���I¾ݾ�  �  �����W4���\��K���Ә�t����`���⥿f������+�S��w/�,]�����&���6�MZ]�����򙿗F���E������(���C�~��5S�B,�>b�F4�0q������������|��f��rY�1&W��._��cq�̆�-(������$վ� ��,�A��#k���������M[���u���e��1؎�� q��F�q&��8�fB��O#��_B�Sl�@t�� ����ު��
���V���؍�Xp�ɅE��� �E`�fqپi����������St���`�߃W�~�X�vd�<�y�����衾ؽ��y�FK	�KY(�=�N���y�h��$���� ��F���򛿾����+b��Z:��V�Y�����7(,��_O��{��y��	����6��ܔ���Ԛ����]oa�R�8�/��D��\�̾�f��b[���7���ul��}\��V��W[�0j���������e����Ⱦv�\���V4� �\��K���Ә�!���o`��O⥿г�������S��u/�`[�ץ��$���6�xX]����(��E��*E�����������~�5S��A,��a�O3�p������0�����|�*f�	oY�F"W��*_�z_q�ʆ�2&�����G"վ� �2,�WA�F#k�G�������[���u���e��؎�� q���F�v&��8��B��O#��_B��l�}t��H����ު�F��QW��iٍ�G	p�ʆE�� �fa��sپ����.�������Nt�{�`���W��X��"d��y����� ꡾Xٽ�{��K	��Y(���N���y�rh������(���F��r󛿚����-b��\:�lX�*������),�6aO�A{�z��y���=7��%����Ԛ�X����oa��8��/�;F��L�̾ i���]��n:�� {l�(�\���V�O][�A5j�b�������g��Z�Ⱦ�  �  nN񾰐�mD�q�x�4������Pǿ��Ϳ��ſ�������?t�e�F��h*��4"�v/���O����2�������ȿӰͿ/�ÿ n��㚒�B]l��:��j��)���q���pЀ�j�a��|M���B���@���G��W�
r�D���-T��PMϾے�/�&���T�)Å�xy������˿��̿����i��U2���ec�<;��W%��*$�2�7��+^�=��>a���Ͻ��̿�̿�ܽ�M����􈿕�Z�u[+�H�xԾ	��@(��ڬu�� Z���H���@���A�~�K�#0_��x}�����泾Lf߾X��e5�fZf�ob��̈��'¿�PͿ�ʿ���m/���傿�<T��1���"��u(���B��Sn������I���ÿ�Ϳ(�ȿ ����3����~���I��������%}ž�K��T���u+k�A0S�*-E��C@��0D��)Q���g�7��%�������M����lD���x����l����Oǿ��Ϳ|�ſB�������t���F��f*��2"�u
/���O����G
������\�ȿ-�Ϳ��ÿ�m�������\l��:�!j��(����3���π�U�a�ByM��B���@��|G��W�/r�\���XR���KϾ��o�&���T���2y��Ə���˿��̿�����h��E2���ec�<;��W%��*$�r�7��+^�p��{a��,н��̿̿"ݽ�����D�����Z��\+�b�fzԾn���*����u��Z���H�p�@�G�A���K��3_�&|}����`賾�g߾���5�[f��b��D����¿IQͿ�ʿ���W0��z悿�>T�ټ1�s�"�iw(�B�B�Un�2���@J����ÿu�Ϳl�ȿY����3��l�~��I��������~ž�M������]0k�i5S�q2E��H@��5D��.Q�0�g�'9�����,����  �  �1���" ���Q���m����0ȿ��޿���ݿ�ſJG��b^��2W�X�6��z-��<�
a����{����U˿>���O�y�ڿO���H������E����w���p㑾L�s���S��@�~�5���3��[:��I�4�c����'ӣ���ξD��SA/�g�d��������>ѿnG�:=��]ֿ��M����w���I�)1���/��E�
�q�����n��;�ӿ�`�hZ��ӿJ���ו��Dk�a�4�P�	��Ծ�ާ��̈�S�g�:L�O�;�14�5�Ek>�PQ��ro�湎��~����ྺY�ù?���x�fZ��M��@�ؿ1�忺�=Kο�@��ƕ���Yf�c?���-��4��^R����n���������ڿ�Q�t���F˿�X��9���t�W�_%�Xo��,�þ�1�� Ԁ��\��wE�,8���3��?7�b�C���Y���|�����\̾�{0��m" ��Q����4���W0ȿV�޿���Lݿ6ſ�F���]��aW�f�6��x-�t<�� a���������T˿u��=O���ڿְ�����a���E�{���v����.⑾��s���S��@���5���3��W:�C�I�d�c����]ѣ���ξy���@/���d����I���ѿ:G�=忱]ֿ���L����w���I�B1�ܲ/�M�E�]�q�J���%o����ӿ�`��Z�f�ӿzJ��ؕ��Ek�j�4�f�	�c�Ծ�৾ψ��g��L���;��54�f5�Ho>�Q�8vo�n������.��]Z�k�?�r�x��Z���M��Եؿ��忂�Lο�A��Ö���[f�g?���-�̐4�h`R����������A�ڿ�Q濶��G˿�X��l�����W��%��p����þ�3��Pր���\��|E�(18���3��D7�.�C�L�Y���|�Y����;��  �  �/��R�"�+�V��$��qo��Q�Ͽb����s��fd̿����~����\��,;�F}1�C�@��Lg�
���?���?�ҿ1V鿢h�"n�
�ȿL���֡��w�I���r�辸����L����o��xO�s�;���1�m�/�n(6�PbE���_��+��C���PXϾ�V���2�z�j�n�������ٿ8��E��޿�����r��-�/O��05�}�3��K���x�������ۿJ]�^Y�,�ۿ]⽿W���h�q��68�:���[վn릾�����9c���G��^7�a0�&�0��):��L�	>k���0ԯ�� �2b���C����k���UEſ��?����꿑ֿ=���14����l�(�C��1��8���W�������F�ȿ�t�hi��O���ҿQ[��)����]���'�ۻ����þ2㚾y�}���X�\#A��4��/�3��6?�WcU���x�4������L.����"���V�r$��8o���Ͽ�翧�����c̿���:}����\��*;�9{1�+�@��Jg����G���Z�ҿeU��gￍm㿏�ȿ燦�������I�c�Y�辐����K���o��uO�&�;�<�1���/��$6��^E�ʁ_��)��}����VϾ/V�֞2�Мj�!���W��Yٿ�7쿧E���޿�����r�� �5O��05���3��K��x�!������]�ۿ�]�Y��ۿ�⽿˩��`�q��78�O���]վ����t>c�>�G�,c7��0�j1��-:���L�iAk�����կ��!��b�U�C�w��֑���EſD�����sֿ2���25����l�2�C��1���8�E X�M��F����ȿu㿾i�P��ҿ[��[���r]�P�'�D�����þ!嚾Ⱦ}�P�X�E(A��4��/�3�W;?��gU���x��5������  �  �1���" ���Q���m����0ȿ��޿���ݿ�ſJG��b^��2W�X�6��z-��<�
a����{����U˿>���O�y�ڿO���H������E����w���p㑾L�s���S��@�~�5���3��[:��I�4�c����'ӣ���ξD��SA/�g�d��������>ѿnG�:=��]ֿ��M����w���I�)1���/��E�
�q�����n��;�ӿ�`�hZ��ӿJ���ו��Dk�a�4�P�	��Ծ�ާ��̈�S�g�:L�O�;�14�5�Ek>�PQ��ro�湎��~����ྺY�ù?���x�fZ��M��@�ؿ1�忺�=Kο�@��ƕ���Yf�c?���-��4��^R����n���������ڿ�Q�t���F˿�X��9���t�W�_%�Xo��,�þ�1�� Ԁ��\��wE�,8���3��?7�b�C���Y���|�����\̾�{0��m" ��Q����4���W0ȿV�޿���Lݿ6ſ�F���]��aW�f�6��x-�t<�� a���������T˿u��=O���ڿְ�����a���E�{���v����.⑾��s���S��@���5���3��W:�C�I�d�c����]ѣ���ξy���@/���d����I���ѿ:G�=忱]ֿ���L����w���I�B1�ܲ/�M�E�]�q�J���%o����ӿ�`��Z�f�ӿzJ��ؕ��Ek�j�4�f�	�c�Ծ�৾ψ��g��L���;��54�f5�Ho>�Q�8vo�n������.��]Z�k�?�r�x��Z���M��Եؿ��忂�Lο�A��Ö���[f�g?���-�̐4�h`R����������A�ڿ�Q濶��G˿�X��l�����W��%��p����þ�3��Pր���\��|E�(18���3��D7�.�C�L�Y���|�Y����;��  �  nN񾰐�mD�q�x�4������Pǿ��Ϳ��ſ�������?t�e�F��h*��4"�v/���O����2�������ȿӰͿ/�ÿ n��㚒�B]l��:��j��)���q���pЀ�j�a��|M���B���@���G��W�
r�D���-T��PMϾے�/�&���T�)Å�xy������˿��̿����i��U2���ec�<;��W%��*$�2�7��+^�=��>a���Ͻ��̿�̿�ܽ�M����􈿕�Z�u[+�H�xԾ	��@(��ڬu�� Z���H���@���A�~�K�#0_��x}�����泾Lf߾X��e5�fZf�ob��̈��'¿�PͿ�ʿ���m/���傿�<T��1���"��u(���B��Sn������I���ÿ�Ϳ(�ȿ ����3����~���I��������%}ž�K��T���u+k�A0S�*-E��C@��0D��)Q���g�7��%�������M����lD���x����l����Oǿ��Ϳ|�ſB�������t���F��f*��2"�u
/���O����G
������\�ȿ-�Ϳ��ÿ�m�������\l��:�!j��(����3���π�U�a�ByM��B���@��|G��W�/r�\���XR���KϾ��o�&���T���2y��Ə���˿��̿�����h��E2���ec�<;��W%��*$�r�7��+^�p��{a��,н��̿̿"ݽ�����D�����Z��\+�b�fzԾn���*����u��Z���H�p�@�G�A���K��3_�&|}����`賾�g߾���5�[f��b��D����¿IQͿ�ʿ���W0��z悿�>T�ټ1�s�"�iw(�B�B�Un�2���@J����ÿu�Ϳl�ȿY����3��l�~��I��������~ž�M������]0k�i5S�q2E��H@��5D��.Q�0�g�'9�����,����  �  �����W4���\��K���Ә�t����`���⥿f������+�S��w/�,]�����&���6�MZ]�����򙿗F���E������(���C�~��5S�B,�>b�F4�0q������������|��f��rY�1&W��._��cq�̆�-(������$վ� ��,�A��#k���������M[���u���e��1؎�� q��F�q&��8�fB��O#��_B�Sl�@t�� ����ު��
���V���؍�Xp�ɅE��� �E`�fqپi����������St���`�߃W�~�X�vd�<�y�����衾ؽ��y�FK	�KY(�=�N���y�h��$���� ��F���򛿾����+b��Z:��V�Y�����7(,��_O��{��y��	����6��ܔ���Ԛ����]oa�R�8�/��D��\�̾�f��b[���7���ul��}\��V��W[�0j���������e����Ⱦv�\���V4� �\��K���Ә�!���o`��O⥿г�������S��u/�`[�ץ��$���6�xX]����(��E��*E�����������~�5S��A,��a�O3�p������0�����|�*f�	oY�F"W��*_�z_q�ʆ�2&�����G"վ� �2,�WA�F#k�G�������[���u���e��؎�� q���F�v&��8��B��O#��_B��l�}t��H����ު�F��QW��iٍ�G	p�ʆE�� �fa��sپ����.�������Nt�{�`���W��X��"d��y����� ꡾Xٽ�{��K	��Y(���N���y�rh������(���F��r󛿚����-b��\:�lX�*������),�6aO�A{�z��y���=7��%����Ԛ�X����oa��8��/�;F��L�̾ i���]��n:�� {l�(�\���V�O][�A5j�b�������g��Z�Ⱦ�  �  pK�������'��B���_���z�"������u���^q��sQ�Œ0��l��G���f��v�w�7��X�_�w��m���ʉ��Y��gu�rY�փ<�_"�Jp�`�����־�ּ��y�����#���8|��;y�!́�#+��Ժ��bv��c�ʾf�������j0�~mL�Hni��9������ 爿�K��zFg��@F�2�&����sX ��8�����_#�*�B�q�c����^m���"���[��X�l���O�%_3�����
�
G��;`���7՟�9Î��Â�(�y�<6{���(��6���,��ȰӾlF�@B
���m9�0V�7�r��l��Q����/��H�z�Q�\�-6;�R�X��?���J�9���%-�w�M�Gn�����>�������ً}��c���E���*��E�� ��Cྛžk���ͥ���$�����a�x�%�~�����ΰ��u ���G¾N
ݾ�I��P���'���B��_�K�z��􆿨��������\q�RrQ�R�0����������Pd��t�ś7�i�X��w��l��ʉ�Y��Nfu�xqY�_�<��^"��o�������־|ռ�cx��H�/"���4|��7y�ˁ��(������Nt��d�ʾ���� ���j0��lL��mi��9��X����房�K��DFg��@F�$�&�����X �&9����e_#���B���c����m��P#��Z\��:�l���O�-`3������xI꾇�;�����ן��Ŏ�5Ƃ��y��:{�򄾳*���7��Z.���Ӿ�G��B
�����m9��0V� �r�Km��᫉��0����z��\��7;��S��eC��-L�����&-���M�Tn�������������f�}�* c�/�E�M�*��F�| ��E��ž
��������'�����R�x��~�i���b����"���I¾ݾ�  �  n��.�+%���2�� A�K4N���V��~W��N��=�IZ&�����|��� ݾ��վ2N��:��'���+���A��_Q�v(X�~U�a�K���=���/�`a"������%O�����=H˾�ҳ��P��cA��-���\���Ҫ�Sm���kپ�)�����z�g ��|)��`7�G�E���Q�PX�{�U��I���5�5f�;��7쾾�ؾ�|׾�-�8������Y3�G�G���T��@X�6�R�2G�T�8���*��Q�?���5�~���Gܾ�þW���`���΃��a�������w����Ⱦ8������	�'F��!�X�-��2<�� J�O�T�NX��R���C��9.����*�~���־]۾S�򾧁�x�#�a�:�3�L���V�|VW�OtO���B��04�N�&��c�]���:�|��Ӿ9����������Г����ڤ�����,�оS��F�����z�s*%�i�2� A��3N���V�~W�7�N�s=�Y&�f���y���ݾx�վ�Jᾘ7�������+�9�A�s^Q��'X�U}U�ǈK�M�=�R�/�a"�6��C�7N������F˾ѳ�$O��Z?���*���Z���Ъ�k���iپ�'�����y�����{)��_7���E�N�Q��X��U�ӍI���5�f�+���7��ؾ�|׾).龍��H��Z3�ۯG�5�T��AX�
�R� 3G�P�8���*�S�t���6�����Iܾ�þ
������X���Đ��ʮ���x��D�Ⱦ��P���g�	��F�l!���-�b3<��!J�%�T�OX��R��C�R;.�x��=,����־`۾3�������#�h�:� M���V�'WW��tO�3�B��14��&��d�c���;��~��Ӿ<���Ħ�R���ԓ�<���ݤ�c�����о���?���  �  b�*�.�/��1��1�� 1��0��a/��m*�� ��9��|��Ⱦ�'������5��^Sξ��r��{�Wq#���+���/�Y1�1�2#1�F�0���.�W,)�i���}�.���a߾�+žU_��ie��ꬼ���ҾG��Y<	�_��_.%�I�,��N0�S 1�1�h$1��0�[/.�#�'����L���'��>rھĸ��X򳾏3��0���"D׾q�����<=��&�d�-��0�##1��1�>"1��|0�l-�0C&��x���f���Ĵվ����Ⲿ
`���¾�ܾ$��j��:w�9C(��i.���0�+$1�u1��1�l30���,���$����M���\1Ѿ�û��2���굾`ƾ�ᾟ� �D^������)��/���0��!1�.1��1�$�/�ӌ+�D�"�,��(�����@�̾�G��iⱾѷ�
5ʾ�5�8��D����!��*�n�/��1��1��1�t�0�Fa/��l*�>� �����y�K�Ⱦ%����;��sPξ!���p��z�Zp#���+��/��1��1��"1��0���.�,)����<}�����Y_߾�)ž-]��c�������Ҿ���,;	�>��N-%�K�,��M0��1�U1��#1�Q�0��..���'�C����Q'��rھ˸�����3�������D׾�q��}���=���&�'�-���0�$1��1�X#1�~0�Hm-��D&�z�^�>�����վՖ��2岾�b��L�¾�ܾ���!���w��C(�:j.���0��$1��1�T1�$40���,� �$�!�;O���M4Ѿ�ƻ��5�����bƾN��� �E_����K�)�o/���0�~"1��1��1�#�/���+���"��������龯�̾2K���屾tԷ�>8ʾ�8澓��x��˒!��  �  ҴW���V���M�5@�r�1��v$��u�	��4�55��yϾ0w��i񣾤���*ߓ��������������#վ���D��˔��
��N'�x�4��]C�6P�a�W�;�V�F-L�d�9��_"��N��$�%�ھ�U־�徿:�����/���D�I-S��VX�V@T�1iI� e;�7-��U �����+	�d)��ڗ�i%ǾQ���垾B�������g��&��rmľ��ݾ�^�����__����ٴ+��9���G�PS��NX�C:T���F�s2�r��d����o	׾�)پ��������7�tJ�&�U���W�u7Q���D��6�_�(�X�w���;�ھ���׾����ũ����F	��Q���
)�������̾�U����~���-�u#��F0�N�>�8L�^�U�{X�n�P��r@��N*�����7��*�6�վJ޾�X���0���'�;4>�LNO��W��V��M�y4@���1�Qv$�5u�Q��3�R3��wϾ�t����}��tܓ�牙����z����!վ���k����
�WN'�B�4��]C�P�<�W���V��,L�ل9�*_"��M�v"�ܒھ�S־]��s9�k��̄/�p�D�&,S��UX�^?T�QhI�8d;�a6-��T �}���+	��(��`��%Ǿ�P���垾3B�����dh�����Knľ��ݾ `��{��&`����е+��9���G�VQS�'PX��;T���F��2��s�`f���:׾P,پc����j��Y7��tJ���U���W��7Q�C�D�_�6���(��X�9���<����]�׾%��Eȩ�ۻ���������+�����۬̾|W澪���M���.�3#�eG0�'�>�9L�x�U��	X�ܶP�Rt@�7P*�̵�];���-��վ�޾\��X2��'��5>�iOO��  �  ?ɉ������y��N^��6A��r&����Wi���t۾��������������~�>�x��|��Z⊾+���/���}ƾ�����u��,���G�\�d�@�~�v�<n�����jl�K�K�x+�7_���e��������	=��^^�h�{�􈇿撉��g	q�8�T���7�j�&0	�̀�s-Ҿ.ݸ����J���^����z�Z	z��H�������頾FD��X.Ͼ� ��a��;�4�LQ��n��悿�M���&��%�~�P�a���@�d�!���
�'��� � ���a)(�7H��i��恿���m}��������g�o�J���.���� �N5�dVɾ05��i����a���U���y��|�����Mܔ������-��dNؾ����1���#��>�[�`�v��ǅ��ω�q���v�W�:�5������С���*�`��M2�DOS���r�l���ȉ�����H�y�EN^�L6A�Lr&����g��s۾����!�軖�x�� ~�E�x�ez���ߊ��)���_{ƾ5�ᾈ�iu��,�j�G�X�d�@�~�o�'n�����ljl���K�.w+�"^����ɞ�����H���=�i]^� �{�Z���V���Dyq�e�T�"�7�si��/	����,Ҿ�ܸ����lJ���^��J�z�
z�)I��d���l꠾PE���/Ͼ2���E��9�4�+MQ��	n�H炿�N���'����~���a���@���!�x�
����~� ��t*(�H��i�灿����}��ɢ���g���J���.�������6�HXɾT7������ud��vX���y���|�VĆ��ޔ�ٟ��}/��.Pؾ,��������#��>�[�l�v�Aȅ��Љ�8���v��W�-�5������ҥ���,��a��O2��PS��r����  �  �g��<ꦿ|̗�\���CZ��I2��.�>���
Ǿ�慨����趀�>i���Z���V�"]�j�m����e���򮾒�ξ����D���:�q�c��퇿�͛�6�����_ţ��V��Ԋx�D#M�]�*���7�����O<���d��̈�뜿ù��ѫ��Ƣ�+I��	iw�XJL�n&����++ྥ����������5x�9c��VX�X�W��a� bu������������۾���֧"�L�G��|r�� ��-��mU��N���Ȟ�>����i�0P@�`�!���������'���H�P�s����Q7��糫���������sR���h�S�>��d��T���Ӿ���혾�߅��p��s^�w�V��Y��g��7~�}ŏ����PFþ���W��*>.�/�U�����߯������Y������阿҃���Z�Q�4������:��,1�	AV�UO��oʖ�:���Zg���馿 ̗���CZ�I2�G.���N	Ǿ�����۴���i���Z�*�V�x]��m����������\�ξ��������:�w�c��͛�;�����9ţ��V���x�O"M�:�*���T6�N��&N<�6�d��ˈ�iꜿ ���qЫ�nƢ��H��+hw��IL�em&���G*�����������I5x�9c�
WX��W��a�ccu�գ����T�����۾�����"�Q�G��}r�����-��!V������Ȟ��>��S�i��Q@���!�R��b����'�ܽH�9�s�����7�������������~R���h���>�.e��U��b	Ӿ����	ⅾ�p��x^�BW���Y��g�T<~��Ǐ����HþO��,��?.��U�/���o�������bZ����꘿|Ӄ���Z�u�4�"!���-<��.1��BV�'P��(˖�ه���  �  ��ͿS�ƿ,����k��
�u��A�E{��0����_��a��bnf��6P�+�C�DS@�B�E�=DT���l�0ň������Ǿ?����  ���L���}ȝ��㷿�eɿƇͿ,ÿoج��Ȋk���@�Ԗ'���"�,3���V�m������K��L�ʿ�Ϳ������ƍ�Sbc�Ǎ2�B����ܾⱾP���w{���]��K���A�!A�_�I��A[���w�:�����+!׾���6�-���]�)�����������h̿[�˿8���Aأ�������[�$76�2�#��&��=�:f�vō�l穿�
��Ϳ��ʿ^���렿 ,���R��s$��� ���̾ׄ���?��'Bp��uV���F��x@�!�B��YN��kc�^����:���1��b辏g�x�<��eo�6���د��Ŀ�Ϳ�ȿc3���u����|��HM���-�Y"��w+���H���v��I��r���+�ƿH�Ϳ�ƿϞ���k��z�u���A��z��/���s]�����yjf��2P�߽C��N@���E�+@T���l��È������Ǿ�����  ���L�#���ȝ��㷿�eɿ��Ϳÿ.ج�~ˉk���@�~�'�=�"��*3��V�Yl��W���'K����ʿͿv��p��2ƍ��ac��2����ܾ͗f᱾�O��w{�;�]��K���A��!A�k�I�C[�P�w�J�������"׾���$�-��]�����{�������i̿�˿���٣�w�����[��86�ȭ#�F&�=�^f��ō��穿�
��(Ϳ��ʿ^���렿),���R�	t$�� �%�̾d���hA��,Fp�DzV�"�F�\}@���B�a^N�-pc�b⁾�<��h3���ih�W�<��fo��6��ٯ���Ŀ��Ϳ�ȿ[4���v����|��JM���-��"��y+���H���v�{J��3���Їƿ�  �  �����ݿ��ƿ����kJ��{N�S��)���L���ᖾ�tz��>X�1�B�E�6�L�3�u�8�F�}�^���u��Ȟƾ� �%�'�t�Z�����q2����̿�H�a!�}�ٿ����ş�	����&P�y�3��A.��@�ti�nX�����غϿ8����/�׿����y���tu�/�<�c.�P�ݾ�F��"3��gm��O��=���4��c4�}B<�SDM��oi�Y<��9�����׾���[Q7��n�����'���տ�����㿪}ҿG����䔿��n��(D��#/���1���K�F�z�1��������׿��>��٭Ͽ�ޱ��A��_a�c�,�L��b̾'ۡ������b�$�H��9��3�6�b�@��DU���u�����n����꾥�LwH�����9���Zÿ|�ۿVr�Q�߿��ɿ
Ȫ�Mf��%j^���:��[-�s�7�)jY�m�����ʪƿ��ݿ�濁�ݿ@�ƿ<���#J���zN������`K��_���0qz��:X�-�B��6��3�]�8��|F��^����1��֝ƾ@ ��'��Z�Đ���2����̿�H�_!�^�ٿh��^ş������%P��3�E@.���@��i��W��;���Ͽ���R�応�׿����x��tu���<��-�a�ݾ�E���2��cfm���O��=��4�Pd4��C<��EM�Qqi�j=��|���k�׾���LR7��n��������Gտf�俶��{~ҿ����唿D�n��*D�G%/��1�E�K�o�z����宼���׿;��E��խϿ�ޱ��A��3_a���,�����̾�ܡ�����tb�K�H�d�9�{�3�r6���@�(IU���u�񄓾Pp����꾂�0xH���������Zÿ0�ۿ%s�9�߿��ɿɪ�ng��vl^��:�9^-���7�ClY�f�������ƿA�ݿ�  �  ����:y���h��*�g�Lw=����龖� g��R�g�ϦA��@(�K;����;�q����+�,�Y�H�JUr��얾y<��~R���]�L�F���p��%���z���`�����ȉ��ԕ_�7�8�J6�����`)�ZK)��M��v�m����S���������M���Y�5�/�s<
�\�־)���M ��n^Y��7�[�!�-��]���#�� ��5���T����F����о�t�RV+�G�T�}P~�C%�������������
fz�fR���,�#j���&d�r�;�4�[�(x��c�����kN��u挿#{u�<{K���"��W��ۤž�䚾��w�ͺL���/����/���S�t��x���
&��B>�ۺb�V׋�����U��
���8�nc��n��OL��̐��b���Nf��Fm���D�)l"�4*��w�q	�N3�{�@��h�������������x��)h����g��v=�w����T쵾�e��7�g�g�A�%=(�j7����7�������,�e�H��Rr��떾�;��8R���]�j�F���p��%���z���`����������_�=�8�5����G��'��I)�l�M�Hv�����4S���
������YM��	�Y�o�/��;
�A�־B������d]Y�U�7��!�1�������)��u �w5���T����:H��q�о�u�VW+�f�T��Q~��%��W���F��|����gz�R�[�,��k�����e�cs�^�4�[��x������B��{N��{挿){u�L{K��"�oX����ž暾��w��L�l�/����_��#X�������&��F>���b�ً����XW�����8�wc�Co���L������?���Bg��S!m���D�an"�q,��y�2s	�V5�^�@�Ġh�ۂ��`����  �  �v������V'���a��8���s��Hٴ�6���)�i���D���+�u�O��8F��
��[��D0�f�K��Lt�����¾�������A���i���u��8��+>��l�~��Y�m�3������pM �@���%�{�G���n��n��D��"甿t䌿�z�5�S���+������Ծn(��s�8�[�%$;��F%����+������e#��98�n�W�����W䢾��ξj"��g'�O�S�v��y���w��C}����r��0L�#�(���� ��������/�g�T���z�팿s锿5?���b�� *n�[F����Q����þ�Κ���y�k�O�F�2�������_���U ��V)�L]A��e�#C��O ��q྾8��R4���\�gE��n���e��ϔ��Y���f�V�?�s�h�dv��1p��Z�܌;���a�%9��Ӓ��Sv��>����&��Ra�[�8�^�I��ش�ͳ���i�O�D� �+�1q�C��'B����W�3A0�b�K�iJt�	���s���3����2�A���i�����u��8��>����~�%Y�t�3�V��9��L ����@%���G�-�n�n��fC���政�㌿�z�T�S���+����Ծ�'������/�[�x#;��F%� ��b+�~����{f#�~;8���W����墾��ξS#��h'�0O���v�mz��mx��F��&�r�=2L�ʈ(�S��� �������/�T�T�P�z�S팿�锿G?���b��	*n�oF����R����þК���y�ĚO��2����9��gc�<��$��Z)�2aA��e��D��"���rྛ9��S4���\��E���n���f������J���f�x�?�:u����z��Qr��\���;�S�a��9��w����  �  _��'��3o���N��,��>���޾uﲾ%����1r���N�#6�r�%�O���������(���:�c�U���{�3��M���`F�1)�T�3���V��Xu�̄��&��7���Kh��.G��#&��x��������1�|8�G	Z��x�Lr��]冿K ��W'e�T[C�� ��Z�P�ξ��������Ve���E�6�/�/�!����Y��� ���-�B�B��`�P���颾��ɾa��Z���q?���a��}�ʅ�����D�z���]�Q�;��G����n���j	���"�D`C���d����ᆿay��r:x��VZ��7���+��T��¦���j���RY��Q=�}:*������Ʈ�n1$�j�3���K�P�m�#��e����tپ���1(��"K���k� 0��FQ�������r�W�R�_�0��U������������-���N���n�����^���&��]2o�B�N�,�7>�\�޾+����R.r�L�N�P6�f�%��J�������ŕ(���:�1�U���{�2�������E�")�a�3�͚V��Xu�̄��&����Kh�.G� #&��w��������{0�	8��Z�;x��q���䆿���_&e�xZC�S� ��Y�;�ξ��������Qe�ގE��/�4�!�q��oZ��� ���-���B�� a�����iꢾ-�ɾ�b��Z���r?�+�a�^�}�|���U����z�M�]���;�'I�t��{�h���	��"�.aC�F�d����&↿wy���:x��VZ��7�P���+��U������+l��nVY�vU=��>*�I����5���5$���3���K�
�m�倎����Tvپ����2(��#K���k��0��R��a����r�O�R�q�0�X� �����7������� -�,�N���n�{���  �  �g���a�k�O��6��c�Ѯ�5Z׾-ѳ�L헾�A���c���I���7�Qz-���*��(/�7L;��N���i�e���ԉ����Zf྇�xm!�g�<�sqT��d��lg��|]��H�[�-�����`����޾��پ�&���
`!� 
=�tMU���d�2g��\���G�B�-������%�ʾ�������^x��Y�cC�H�3���+��9+��\2�	�@�=�V�7�t�����������ƾ�����6�*��&E���Z�M�f���e�W�W�z@�<m$�'�
��W���ھ?Fݾw�������*���E�ݡ[���f�$e��V��?��w$���	���6���ru���ވ�[?m��fQ��=�0�'�*���,�h6��wG���_�2+��3;��\����Ҿ����e���3�c*M��	`���g�3b�H�P�X�6�PY�T/� z�cپ��� ��f�Y�3���M�X�`��g��a���O�{�6�0c�@��Y׾�ϳ��뗾R@���c���I���7��u-�6�*�)$/��G;��N�L�i�Ꙇ�����C���e�d�qm!�o�<�{qT��d��lg��|]���H���-����^��T�޾��پ�#�h��^!��=�'LU�O�d��0g��\���G�m�-�������ʾ����_���]x�_�Y�C�O�3��+��:+��]2�c�@���V�B�t�ě�����L�ƾ~����K�*��'E���Z���f���e�׈W�@��n$���
��Z���ھIݾ�y�������*�A�E�_�[�N�f�\e��V��?��w$���	���K����v������ Cm��jQ��=��#0�ӭ*�\�,��l6�#|G���_�-���<���]��k�Ҿ0���f�u�3�w+M��
`�f�g��4b��P�8�6�J[�_1�?~�x!پ�� � ��h���3�%�M���`��  �  }�>���:�2/�Uj��������s_־k~���u��\��|Ƃ�w�i�,{T��hG���C���I�?�X��eo��>��b��7������`�ܾg�����f"�~\2���<��>���5���%� f�`B��uA׾��¾�Ͼ��3̾4�������/���;�]>���7�1�)�)M�n���7꾓@;_Ŵ�̟�>���ߠ{���a�{"O��E�щD��M��\_��tx�Ŭ�����H��FRʾM�澙��~=��%(��6�>� b<��c1��c�kH
���G�ξhs���d��M7Ծ��� ���#�I�4��=��$=���3�5Z$���& ��ྀ�ľ2p��#o������Tr�+�Z�W�J��C��F���R�?�f����+c���2��r޹�EӾP��	�vc�k�-�-�9�S�>���9�n�+��{�FO�@Sᾃ�Ǿ�%����ž��ݾ�
�"��*���8���>��:�k1/��i�i������:^־}��Lt��ZZ���Ă�6�i��vT��cG��C���I���X�9ao��<��p`�����v�����ܾ�f��y�wf"�q\2�ۂ<��>�_�5��%�Ge��@��]?׾[�¾L;��0̾������z�ɬ/�~�;��[>���7�L�)�\L����P6꾐?;�Ĵ�]˟�Ì��?�{���a��"O�E���D��M�:^_�Pvx�ȭ��0���cI���Sʾ	�澏���>��&(�S�6�j>�cc<�2e1�e��I
���=�ξ>v��-g���9Ծ9������#�ю4�q�=�%=���3�lZ$�# �� �����ľ�q���p����LYr��Z�E�J��C���F�F�R��g���e���4��๾�FӾ�Q�v�	�[d�m�-�S�9���>��9�,��}�"Q�W�f�Ǿ�)��[�ž-�ݾf��#�S*���8��  �  ���;�_������� �:p�*ҾC��P`���.��
7����|��*k�f�Mn�z���ȏ�|/��{k��0ž]�վ��S�����'���z����%��z�������(!ξ{���ԥ�Z󢾺⬾�¾�޾��������d������t���������r�ݾ��̾3e���G��K���(����u��g�`;g�P�s�Đ���_���>���i��z�ʾ47۾~�����������*f���_��)��� �c3⾂�ľ'���cl���ݤ��в�p�ʾ�*����(���L�����*������������羐�׾�Ǿ"l���1��i���������o��;f���i�Hz��z���1��W���P��zSо�ྌ6�jz�C�
��*������Ⱦ�X
����s�׾`��ƛ��[t���1���湾�ԾP��Q�����$���:������������n⾞(Ҿ�A��w^���,���4���|��%k���e�n����hƏ�N-���i���ž�վ�澥���؎�����z�[�������c����oξ}���ҥ���AାE¾��޾w���o���c������s�=��j����q�ݾء̾�d��1G��2K���(����u�h�g�<g�Q�s�o���^`���?���j����ʾ�8۾0�뾿��������[g�@����*�� �H6�e�ľ����o��JाӲ�{�ʾL,龬�����CM����=+�Ԯ�o��n������׾EǾ*n���3������ �����o��@f���i�Mz�}��4��Y��VR��Uо���8�,{��
��+�����%���
������׾􂼾e����w��_5��깾��Ծ!�󾑘�����  �  ����i ����t3��1�C��vG ����Ț�/�ؾ5¾
������u���ֈ��~���~��͇���SǾ�=ݾ<�z,��X� �8���6��+��������3��0���
վ�\��6��9-���7��W$��xK���}���;���"˾��ي񾀙������R8��"�v|�O���>8��g���`Ѿ%���wӤ�^ʓ��8��س��0Q��G�������]�ξ������J����V���7�a��A�jt����l��'�;l���y��������z��������量qͻ�
�Ҿp��������H��$&��7�7��� �4#������v߾��ɾ����w��ۨ��z ��)������r[��Ǣ��"=־I��������������-�F5�0��� �`����@�ܾ�	ƾ�L��ʄ��&Ȉ��ꌾ٦���㬾�zþ��پ��X���Ai �S���2�b1�����F �j����9�ؾ�2¾��������s���ӈ��{���{��'���@QǾ`;ݾ]��*���� ����6��+�k������53��S���	վ}[��n4��S+���5��"��&I���{���9��? ˾��ƈ񾑗�����
��7�/"��{�`���y7�����z`Ѿۇ��VӤ�fʓ�9��/����Q��𤢾U���X�ξ���6������]W���8�t��B��v��+����;/���9���:����}�����������'ϻ�y�Ҿ��������������&�J8���u� ��$�����9y߾�ɾf����y������V��񚋾n���]�����!?־�龐���L���I��P.�6���� �����C��ܾ�ƾ�O�����u�}ˈ��팾򩙾�款N}þO�پ���  �  �Ӿ7X������(<�D^��d��^��S���v��$�ҾJ�������^���qb���ٽ�8�پ����@�
�L0����������7
��� �/E�C�߾^iϾ$X���T���7������y��di��of�9�p��F��D����5���m����Ǿ��ؾC�辦���:�\(��~���u�+�0 �~l羓nɾL����s������鲯��eƾ����{�����m����b��"��������Oھ�ɾ8j��
:��k��kȄ�͇r���f�eh�=�v�v����B��TK��#a���;0�ݾlb���#2	�����1�����*,�W?���	ݾ���m��Q¢��[���8����Ͼ�g�PN��J�E������B9��
�&���'�3�ԾD%ľg���+��"ގ�5e���Dm�#�e�Q�k��~�K��[+���a��9¾6Ӿ�V㾏��I��;��]�Od�^�S������Ҿr�������D���R_���ֽ�J�پ4����
�;/����0��j���7
�x� ��D𾙹߾�hϾ5W���S���6�����}y��`i�tkf�ڡp�sD������3���k����Ǿ��ؾ��� ������'�~�+������8l�tnɾT����s��N���h����fƾ���r|�g��`n�����D��#�����@��VRھ��ɾ�l���<���m��˄��r���f��ih���v�c���nD���L��^b����;�ݾQc�{����2	�����2�����l-�B���ݾ������dŢ��^���;��K�Ͼ4j�UO�cK� �������9�A�����)�2�Ծ�'ľ�i��b.��ᎾCh���Jm�V�e�\�k��~�����-���c���:¾�  �  Gҽ���׾�������k�0�m\;�cr>�g�7��)�������}ܾ�žt>��{�Ⱦ�'㾎v������,�f6:�{�>�\w9�ǧ,��_�}��Q�ﾅ�Ѿ���3��l��B��k�e�W�Q�F���C�/nK�0�[��s�}툾�z��i����
ƾ����S'��P%�
�4��j=��W=���3���"����Q��?�Ҿ[����ܿ�� о���4w�l� ��72���<�"�=�k�5�l6'��5�?��&微�ȾU��В��龊���v��(^�}�L� ND��aE�z�O�gc��;}����]⠾R��2�ξ��뾬���S���*�J^8�Kv>�?*;�G�.����F����/˾�����fþ>�ؾ#m�������&�x�6�l2>�'<���1�hi!��
�.���P ۾����;穾�[��A[����m��yW���H���C�K�G��pU��k�3����X��+����н�`�׾������k��0��[;��q>�y�7��)����I���pܾ{ ž;���ȾZ$��t�<��w�,�45:�w�>��v9��,�_�
����ﾹ�Ѿ$���3���j���@��L�e�ݭQ�DF���C�jK���[���s�t눾�x������<	ƾz��6��&�'P%���4�fj=�PW=���3�x�"����4��H�Ҿ����ݿ� оE�w�� �+82�T�<���=�4�5�I7'��6�A �L���Ⱦ���D���k�����v��-^�l�L��RD�FfE���O�*c�#?}������㠾s��<�ξ���8��;T�E�*�/_8�Zw>�y+;���.�&�����S�澇˾֑��jþ5�ؾ�o��.����&�]�6�,3>��'<���1��i!�#������!۾���L驾�]���]��H�m�{W���H�\�C���G�8vU��k�~����Z�������  �  (�����پ��v��+8��P��3b���g��`��L��[2���� ���K��<پ1��_]����i�8� �Q�s�b�7�g� @_�O�K��)2�t���s����о�����듾�O~��X^��WF�R�5��u,���*���0��	>���R��
o����]������[v�"Q�O�%�j�@�e�W���e��f���Z�6_D��)�ވ�_��S�ܾ�O۾z
������%�zA�i�X���e��Nf�p�Y��C�	)��(��K�W�ľ����Hd��¬r��~U���?���1�+�m�+�UG4�FD��K[��Pz��V���[��֣̾SL�����,!/��=I�ڏ]��gg��d��#T�.�;�������Z��v�پ3�߾dg��0�ZA/�1�I�{\^��g��uc��IS�� ;�������޾"+��m��}��=h���M��h:�ڮ.�|{*���-���8�K�ʴd�vP��@K��������پ
�����*8�u�P�F3b���g��`�ĤL�/Z2�t��Ģ����ᾍ8پ��澕[�-���8���Q�$�b��g�0?_���K�A)2����	s����о�����꓾�M~�V^��TF���5�:r,���*��0��>�ĽR�o������l����t�pP���%���@��W�7�e���f�r�Z�_D�y)�ш�j�󾃎ܾ�O۾�
�@��#�%��zA���X�l�e��Of�5�Y���C��	)��)��M쾌�ľ� ���f����r�w�U���?��1��+���+�bK4��!D��N[��Sz��W���\����̾vM������!/�b>I�Ր]��hg�4d�"%T�͉;����i�����پ��߾�j�����B/�C�I�`]^���g�"vc�dJS�!;���� ��K޾�,��S��3���h���M��m:�E�.��*��-��8��	K��d�dR���L���  �  ��G��t����-���P��p�^���T[�����hNm�8�L��Z+��C������%�]B ����A�2��sT���s��b��A��򬁿Jj�13I��L&��9�U�־������Mrk�3J���2�b�#�1l�S��]��+��>�z2[�����l��e�¾>+�:���9��.\���y�Kƅ�D�����~��c��zA��!�5���&�����]������=��_��|��G���L��VH|���_��}=�) �PE���|Ǿ(���`���_��MA���,�7 �	1����ZK"�Ҵ0��G��$g����i���؊Ѿ�����"�^NE���f�0���@
�����-�v��-X��66���������" �������'�I�l�i�p����>���k����s�y�T�S�1�Ph��`�z�����WNy���S���9�E�'�\�����8I&��27��P��t��8���������.�-�!�P�y�p�
����Z������8Mm���L�#Y+�B����2"�v@ ����n�2��qT�)�s��a���@��q���2Ij��2I�/L&�9�Z�־��������ok�}J���2��#��h�������+��>��.[�O���k��˭¾�)��s�9�R.\�/�y�ƅ����I�~�vc��zA��!�:���&��ߦ���C��t�=���_�"|��G���L��I|���_��~=�!�]G��Ǿh��@c���_�ORA���,�� ��5����SO"�y�0��
G��'g�H������
�Ѿ ����"�OE���f������
��7����v��/X��86���������#��B��"�'�_I���i�✁�X?��	l��6�s��T���1��h��a羊{��̃��\Ry���S�Õ9�J�'�-a�+��(��N&�e77��P���t�C:���  �  &D�����j�B�:��Dc����t��	s�����L��-�_��9����)��֞������ �ޯA�u5h��腿&���R���Վ�gO���\Z��$2��S�hݾ�ԭ�p���y�b�_�?�tK(�������#x��H��� ��4�,�Q��|�ǜ�
�ƾپ���"!��YH��Kp�r0������N���|;��b�x�֟R���-����p��6��A�rQ*�:TN���t��Ɗ��8��5��I����t�*�L��L%��[��̾�Р��/��ْU��6�g|"��2����"\��P��?&�:�<��-^��V���W��s׾˖	��-��U�B�|����U���Ⓙ�����ul�{�E��X#���
�� ��I����H�5��C[�Wf���܎�ZS������م�;�g��a?����J�07������q���I�/����ߥ�.:�G���!�Ī,�iF��wl�?x���B���������:�`Dc�������r������K��ė_�z�9���M���������� ���A��3h�$腿k��R��CՎ��N���[Z��#2�$S��fݾ�ӭ�S����b���?�xH(����1���t��D�+� �/4���Q�z�|��Ŝ�x�ƾe���*"!�YH�pKp�70��y���$���Z;��1�x���R���-������7��A��Q*��TN��t��Ɗ�9��q5������Ղt��L��M%��\��̾�Ҡ�22����U���6��"�W7�(��U`��T�[C&���<��0^�X���X��[t׾m�	���-���U�-�|���������㒿u���^wl�X�E��Z#���
�� �TK�0��ƙ5�<E[��f��Yݎ��S��#���م���g�-b?����2L�8��>��Ȥq���I��/����ڪ�-?�-��3&�(�,�mF�P{l��y���  �  "q��� �V�b�?��j��^���������$P����^f�Χ>���A��������$��#G��^o��R������|��R���ul����`���6���'+�~���l��fS`��<���$��O�}��dl��$�d����0�r�N���z��jȾ�� ��$���M��w�����`���qؙ�)�k���X�q�2�� ����w�ܜ��.�UT���|�Cl���T���P��L^���"|���R�J")�ؙ��ξ,��Ji����R���3�o4�����iK�� ���"��y9�	�[��������"�پ�'�A
2�� \�:[��JV���8���헿1����s��zK�{�'�N����l4�����:���a����^���H}��V��?=���n��pD�tC����=���u���J�o�M�F�,�+�tU�����/�Q������`)�:bC��Hj��9���o��p�����?�/j�x^��T����������<]f�3�>�*��`��������$��!G�]o��Q������{��ȫ��l���`��6�\�*�o���M���P`�L�<���$��L����h�,!��|��0�зN�z�z�=xhȾ� �u�$�d�M�_�w�l���-���Gؙ���j����X�e�2�� ��������Y�.�kUT�(�|��l��U���P���^���#|���R�=#)�ښ��ξb!���k��I�R�U�3�9���&���O��$�5�"��|9��[������c�پz(��
2�]\��[���V���9�������s�e|K�k�'�>����:6�Z����:���a�����ѵ���}�����{=��^�n�8qD��C��󾩘������o��G���+�AZ�y���4�)��z���d)�2fC��Lj�B;���  �  &D�����j�B�:��Dc����t��	s�����L��-�_��9����)��֞������ �ޯA�u5h��腿&���R���Վ�gO���\Z��$2��S�hݾ�ԭ�p���y�b�_�?�tK(�������#x��H��� ��4�,�Q��|�ǜ�
�ƾپ���"!��YH��Kp�r0������N���|;��b�x�֟R���-����p��6��A�rQ*�:TN���t��Ɗ��8��5��I����t�*�L��L%��[��̾�Р��/��ْU��6�g|"��2����"\��P��?&�:�<��-^��V���W��s׾˖	��-��U�B�|����U���Ⓙ�����ul�{�E��X#���
�� ��I����H�5��C[�Wf���܎�ZS������م�;�g��a?����J�07������q���I�/����ߥ�.:�G���!�Ī,�iF��wl�?x���B���������:�`Dc�������r������K��ė_�z�9���M���������� ���A��3h�$腿k��R��CՎ��N���[Z��#2�$S��fݾ�ӭ�S����b���?�xH(����1���t��D�+� �/4���Q�z�|��Ŝ�x�ƾe���*"!�YH�pKp�70��y���$���Z;��1�x���R���-������7��A��Q*��TN��t��Ɗ�9��q5������Ղt��L��M%��\��̾�Ҡ�22����U���6��"�W7�(��U`��T�[C&���<��0^�X���X��[t׾m�	���-���U�-�|���������㒿u���^wl�X�E��Z#���
�� �TK�0��ƙ5�<E[��f��Yݎ��S��#���م���g�-b?����2L�8��>��Ȥq���I��/����ڪ�-?�-��3&�(�,�mF�P{l��y���  �  ��G��t����-���P��p�^���T[�����hNm�8�L��Z+��C������%�]B ����A�2��sT���s��b��A��򬁿Jj�13I��L&��9�U�־������Mrk�3J���2�b�#�1l�S��]��+��>�z2[�����l��e�¾>+�:���9��.\���y�Kƅ�D�����~��c��zA��!�5���&�����]������=��_��|��G���L��VH|���_��}=�) �PE���|Ǿ(���`���_��MA���,�7 �	1����ZK"�Ҵ0��G��$g����i���؊Ѿ�����"�^NE���f�0���@
�����-�v��-X��66���������" �������'�I�l�i�p����>���k����s�y�T�S�1�Ph��`�z�����WNy���S���9�E�'�\�����8I&��27��P��t��8���������.�-�!�P�y�p�
����Z������8Mm���L�#Y+�B����2"�v@ ����n�2��qT�)�s��a���@��q���2Ij��2I�/L&�9�Z�־��������ok�}J���2��#��h�������+��>��.[�O���k��˭¾�)��s�9�R.\�/�y�ƅ����I�~�vc��zA��!�:���&��ߦ���C��t�=���_�"|��G���L��I|���_��~=�!�]G��Ǿh��@c���_�ORA���,�� ��5����SO"�y�0��
G��'g�H������
�Ѿ ����"�OE���f������
��7����v��/X��86���������#��B��"�'�_I���i�✁�X?��	l��6�s��T���1��h��a羊{��̃��\Ry���S�Õ9�J�'�-a�+��(��N&�e77��P���t�C:���  �  (�����پ��v��+8��P��3b���g��`��L��[2���� ���K��<پ1��_]����i�8� �Q�s�b�7�g� @_�O�K��)2�t���s����о�����듾�O~��X^��WF�R�5��u,���*���0��	>���R��
o����]������[v�"Q�O�%�j�@�e�W���e��f���Z�6_D��)�ވ�_��S�ܾ�O۾z
������%�zA�i�X���e��Nf�p�Y��C�	)��(��K�W�ľ����Hd��¬r��~U���?���1�+�m�+�UG4�FD��K[��Pz��V���[��֣̾SL�����,!/��=I�ڏ]��gg��d��#T�.�;�������Z��v�پ3�߾dg��0�ZA/�1�I�{\^��g��uc��IS�� ;�������޾"+��m��}��=h���M��h:�ڮ.�|{*���-���8�K�ʴd�vP��@K��������پ
�����*8�u�P�F3b���g��`�ĤL�/Z2�t��Ģ����ᾍ8پ��澕[�-���8���Q�$�b��g�0?_���K�A)2����	s����о�����꓾�M~�V^��TF���5�:r,���*��0��>�ĽR�o������l����t�pP���%���@��W�7�e���f�r�Z�_D�y)�ш�j�󾃎ܾ�O۾�
�@��#�%��zA���X�l�e��Of�5�Y���C��	)��)��M쾌�ľ� ���f����r�w�U���?��1��+���+�bK4��!D��N[��Sz��W���\����̾vM������!/�b>I�Ր]��hg�4d�"%T�͉;����i�����پ��߾�j�����B/�C�I�`]^���g�"vc�dJS�!;���� ��K޾�,��S��3���h���M��m:�E�.��*��-��8��	K��d�dR���L���  �  Gҽ���׾�������k�0�m\;�cr>�g�7��)�������}ܾ�žt>��{�Ⱦ�'㾎v������,�f6:�{�>�\w9�ǧ,��_�}��Q�ﾅ�Ѿ���3��l��B��k�e�W�Q�F���C�/nK�0�[��s�}툾�z��i����
ƾ����S'��P%�
�4��j=��W=���3���"����Q��?�Ҿ[����ܿ�� о���4w�l� ��72���<�"�=�k�5�l6'��5�?��&微�ȾU��В��龊���v��(^�}�L� ND��aE�z�O�gc��;}����]⠾R��2�ξ��뾬���S���*�J^8�Kv>�?*;�G�.����F����/˾�����fþ>�ؾ#m�������&�x�6�l2>�'<���1�hi!��
�.���P ۾����;穾�[��A[����m��yW���H���C�K�G��pU��k�3����X��+����н�`�׾������k��0��[;��q>�y�7��)����I���pܾ{ ž;���ȾZ$��t�<��w�,�45:�w�>��v9��,�_�
����ﾹ�Ѿ$���3���j���@��L�e�ݭQ�DF���C�jK���[���s�t눾�x������<	ƾz��6��&�'P%���4�fj=�PW=���3�x�"����4��H�Ҿ����ݿ� оE�w�� �+82�T�<���=�4�5�I7'��6�A �L���Ⱦ���D���k�����v��-^�l�L��RD�FfE���O�*c�#?}������㠾s��<�ξ���8��;T�E�*�/_8�Zw>�y+;���.�&�����S�澇˾֑��jþ5�ؾ�o��.����&�]�6�,3>��'<���1��i!�#������!۾���L驾�]���]��H�m�{W���H�\�C���G�8vU��k�~����Z�������  �  �Ӿ7X������(<�D^��d��^��S���v��$�ҾJ�������^���qb���ٽ�8�پ����@�
�L0����������7
��� �/E�C�߾^iϾ$X���T���7������y��di��of�9�p��F��D����5���m����Ǿ��ؾC�辦���:�\(��~���u�+�0 �~l羓nɾL����s������鲯��eƾ����{�����m����b��"��������Oھ�ɾ8j��
:��k��kȄ�͇r���f�eh�=�v�v����B��TK��#a���;0�ݾlb���#2	�����1�����*,�W?���	ݾ���m��Q¢��[���8����Ͼ�g�PN��J�E������B9��
�&���'�3�ԾD%ľg���+��"ގ�5e���Dm�#�e�Q�k��~�K��[+���a��9¾6Ӿ�V㾏��I��;��]�Od�^�S������Ҿr�������D���R_���ֽ�J�پ4����
�;/����0��j���7
�x� ��D𾙹߾�hϾ5W���S���6�����}y��`i�tkf�ڡp�sD������3���k����Ǿ��ؾ��� ������'�~�+������8l�tnɾT����s��N���h����fƾ���r|�g��`n�����D��#�����@��VRھ��ɾ�l���<���m��˄��r���f��ih���v�c���nD���L��^b����;�ݾQc�{����2	�����2�����l-�B���ݾ������dŢ��^���;��K�Ͼ4j�UO�cK� �������9�A�����)�2�Ծ�'ľ�i��b.��ᎾCh���Jm�V�e�\�k��~�����-���c���:¾�  �  ����i ����t3��1�C��vG ����Ț�/�ؾ5¾
������u���ֈ��~���~��͇���SǾ�=ݾ<�z,��X� �8���6��+��������3��0���
վ�\��6��9-���7��W$��xK���}���;���"˾��ي񾀙������R8��"�v|�O���>8��g���`Ѿ%���wӤ�^ʓ��8��س��0Q��G�������]�ξ������J����V���7�a��A�jt����l��'�;l���y��������z��������量qͻ�
�Ҿp��������H��$&��7�7��� �4#������v߾��ɾ����w��ۨ��z ��)������r[��Ǣ��"=־I��������������-�F5�0��� �`����@�ܾ�	ƾ�L��ʄ��&Ȉ��ꌾ٦���㬾�zþ��پ��X���Ai �S���2�b1�����F �j����9�ؾ�2¾��������s���ӈ��{���{��'���@QǾ`;ݾ]��*���� ����6��+�k������53��S���	վ}[��n4��S+���5��"��&I���{���9��? ˾��ƈ񾑗�����
��7�/"��{�`���y7�����z`Ѿۇ��VӤ�fʓ�9��/����Q��𤢾U���X�ξ���6������]W���8�t��B��v��+����;/���9���:����}�����������'ϻ�y�Ҿ��������������&�J8���u� ��$�����9y߾�ɾf����y������V��񚋾n���]�����!?־�龐���L���I��P.�6���� �����C��ܾ�ƾ�O�����u�}ˈ��팾򩙾�款N}þO�پ���  �  ���;�_������� �:p�*ҾC��P`���.��
7����|��*k�f�Mn�z���ȏ�|/��{k��0ž]�վ��S�����'���z����%��z�������(!ξ{���ԥ�Z󢾺⬾�¾�޾��������d������t���������r�ݾ��̾3e���G��K���(����u��g�`;g�P�s�Đ���_���>���i��z�ʾ47۾~�����������*f���_��)��� �c3⾂�ľ'���cl���ݤ��в�p�ʾ�*����(���L�����*������������羐�׾�Ǿ"l���1��i���������o��;f���i�Hz��z���1��W���P��zSо�ྌ6�jz�C�
��*������Ⱦ�X
����s�׾`��ƛ��[t���1���湾�ԾP��Q�����$���:������������n⾞(Ҿ�A��w^���,���4���|��%k���e�n����hƏ�N-���i���ž�վ�澥���؎�����z�[�������c����oξ}���ҥ���AାE¾��޾w���o���c������s�=��j����q�ݾء̾�d��1G��2K���(����u�h�g�<g�Q�s�o���^`���?���j����ʾ�8۾0�뾿��������[g�@����*�� �H6�e�ľ����o��JाӲ�{�ʾL,龬�����CM����=+�Ԯ�o��n������׾EǾ*n���3������ �����o��@f���i�Mz�}��4��Y��VR��Uо���8�,{��
��+�����%���
������׾􂼾e����w��_5��깾��Ծ!�󾑘�����  �  }�>���:�2/�Uj��������s_־k~���u��\��|Ƃ�w�i�,{T��hG���C���I�?�X��eo��>��b��7������`�ܾg�����f"�~\2���<��>���5���%� f�`B��uA׾��¾�Ͼ��3̾4�������/���;�]>���7�1�)�)M�n���7꾓@;_Ŵ�̟�>���ߠ{���a�{"O��E�щD��M��\_��tx�Ŭ�����H��FRʾM�澙��~=��%(��6�>� b<��c1��c�kH
���G�ξhs���d��M7Ծ��� ���#�I�4��=��$=���3�5Z$���& ��ྀ�ľ2p��#o������Tr�+�Z�W�J��C��F���R�?�f����+c���2��r޹�EӾP��	�vc�k�-�-�9�S�>���9�n�+��{�FO�@Sᾃ�Ǿ�%����ž��ݾ�
�"��*���8���>��:�k1/��i�i������:^־}��Lt��ZZ���Ă�6�i��vT��cG��C���I���X�9ao��<��p`�����v�����ܾ�f��y�wf"�q\2�ۂ<��>�_�5��%�Ge��@��]?׾[�¾L;��0̾������z�ɬ/�~�;��[>���7�L�)�\L����P6꾐?;�Ĵ�]˟�Ì��?�{���a��"O�E���D��M�:^_�Pvx�ȭ��0���cI���Sʾ	�澏���>��&(�S�6�j>�cc<�2e1�e��I
���=�ξ>v��-g���9Ծ9������#�ю4�q�=�%=���3�lZ$�# �� �����ľ�q���p����LYr��Z�E�J��C���F�F�R��g���e���4��๾�FӾ�Q�v�	�[d�m�-�S�9���>��9�,��}�"Q�W�f�Ǿ�)��[�ž-�ݾf��#�S*���8��  �  �g���a�k�O��6��c�Ѯ�5Z׾-ѳ�L헾�A���c���I���7�Qz-���*��(/�7L;��N���i�e���ԉ����Zf྇�xm!�g�<�sqT��d��lg��|]��H�[�-�����`����޾��پ�&���
`!� 
=�tMU���d�2g��\���G�B�-������%�ʾ�������^x��Y�cC�H�3���+��9+��\2�	�@�=�V�7�t�����������ƾ�����6�*��&E���Z�M�f���e�W�W�z@�<m$�'�
��W���ھ?Fݾw�������*���E�ݡ[���f�$e��V��?��w$���	���6���ru���ވ�[?m��fQ��=�0�'�*���,�h6��wG���_�2+��3;��\����Ҿ����e���3�c*M��	`���g�3b�H�P�X�6�PY�T/� z�cپ��� ��f�Y�3���M�X�`��g��a���O�{�6�0c�@��Y׾�ϳ��뗾R@���c���I���7��u-�6�*�)$/��G;��N�L�i�Ꙇ�����C���e�d�qm!�o�<�{qT��d��lg��|]���H���-����^��T�޾��پ�#�h��^!��=�'LU�O�d��0g��\���G�m�-�������ʾ����_���]x�_�Y�C�O�3��+��:+��]2�c�@���V�B�t�ě�����L�ƾ~����K�*��'E���Z���f���e�׈W�@��n$���
��Z���ھIݾ�y�������*�A�E�_�[�N�f�\e��V��?��w$���	���K����v������ Cm��jQ��=��#0�ӭ*�\�,��l6�#|G���_�-���<���]��k�Ҿ0���f�u�3�w+M��
`�f�g��4b��P�8�6�J[�_1�?~�x!پ�� � ��h���3�%�M���`��  �  _��'��3o���N��,��>���޾uﲾ%����1r���N�#6�r�%�O���������(���:�c�U���{�3��M���`F�1)�T�3���V��Xu�̄��&��7���Kh��.G��#&��x��������1�|8�G	Z��x�Lr��]冿K ��W'e�T[C�� ��Z�P�ξ��������Ve���E�6�/�/�!����Y��� ���-�B�B��`�P���颾��ɾa��Z���q?���a��}�ʅ�����D�z���]�Q�;��G����n���j	���"�D`C���d����ᆿay��r:x��VZ��7���+��T��¦���j���RY��Q=�}:*������Ʈ�n1$�j�3���K�P�m�#��e����tپ���1(��"K���k� 0��FQ�������r�W�R�_�0��U������������-���N���n�����^���&��]2o�B�N�,�7>�\�޾+����R.r�L�N�P6�f�%��J�������ŕ(���:�1�U���{�2�������E�")�a�3�͚V��Xu�̄��&����Kh�.G� #&��w��������{0�	8��Z�;x��q���䆿���_&e�xZC�S� ��Y�;�ξ��������Qe�ގE��/�4�!�q��oZ��� ���-���B�� a�����iꢾ-�ɾ�b��Z���r?�+�a�^�}�|���U����z�M�]���;�'I�t��{�h���	��"�.aC�F�d����&↿wy���:x��VZ��7�P���+��U������+l��nVY�vU=��>*�I����5���5$���3���K�
�m�倎����Tvپ����2(��#K���k��0��R��a����r�O�R�q�0�X� �����7������� -�,�N���n�{���  �  �v������V'���a��8���s��Hٴ�6���)�i���D���+�u�O��8F��
��[��D0�f�K��Lt�����¾�������A���i���u��8��+>��l�~��Y�m�3������pM �@���%�{�G���n��n��D��"甿t䌿�z�5�S���+������Ծn(��s�8�[�%$;��F%����+������e#��98�n�W�����W䢾��ξj"��g'�O�S�v��y���w��C}����r��0L�#�(���� ��������/�g�T���z�팿s锿5?���b�� *n�[F����Q����þ�Κ���y�k�O�F�2�������_���U ��V)�L]A��e�#C��O ��q྾8��R4���\�gE��n���e��ϔ��Y���f�V�?�s�h�dv��1p��Z�܌;���a�%9��Ӓ��Sv��>����&��Ra�[�8�^�I��ش�ͳ���i�O�D� �+�1q�C��'B����W�3A0�b�K�iJt�	���s���3����2�A���i�����u��8��>����~�%Y�t�3�V��9��L ����@%���G�-�n�n��fC���政�㌿�z�T�S���+����Ծ�'������/�[�x#;��F%� ��b+�~����{f#�~;8���W����墾��ξS#��h'�0O���v�mz��mx��F��&�r�=2L�ʈ(�S��� �������/�T�T�P�z�S팿�锿G?���b��	*n�oF����R����þК���y�ĚO��2����9��gc�<��$��Z)�2aA��e��D��"���rྛ9��S4���\��E���n���f������J���f�x�?�:u����z��Qr��\���;�S�a��9��w����  �  XpF���@�J�0������ ��Mо,���$у�?�S���-�I���� �����޽�2۽�u���H�2����4���]����Ư��Z�ھ�,�ED��4�X�B��&F���=�D@,�yY�WR���^־p��z���
ʾ#�龣�
��m"�7�l�C���E��C<�֌)��~��M��U��k���A�t��qE���#��N�����彁oܽ��۽p0�.��{�	�uw �AA��n�k���c������k��'���:�PAE�b�D��8���$��g��V�k�̾�ӻ�������ҾQ���ѱ���)��Z<�g�E���C���6���!�z	�� ྋ3��7C���7c�7�8�8�����@񽣐�S۽��ݽ��:�����*�N�N���������8˾�k��6�Q.��H?��[F�*�A�"�2�mA�������žd`����¾@�ݾ��!��x�0�h�@�IoF���@���0����$� ��Lо���σ�t�S�{�-����>� �p��/޽�*۽�m���E�L��c�4��]�{���i���<�ھ�,�WD�-�4�R�B��&F�W�=��?,��X�uP���\־�m������ʾJ��9�
�7l"��7�.�C���E��B<��)��}�2L�T��]�����t�0pE���#�j��������1pܽ5�۽p2佴0��&�	�wy ��A�֔n�����#������~��8'��:��BE�ңD���8�-�$�~i�Z�̾�ֻ�� ��W�Ҿ�������p�)�w[<���E�%�C��6���!��	�R�-4��D���9c���8�s����UH�Ϙ�h[۽�ݽ��1������*�ƮN�ŉ�������:˾�m��6�$R.�J?�]F���A���2�YC����J���!ž�d���þ�ݾO������0���@��  �  ��@��;�O�+�,���d��y�̾|��M8���%T��;/���?F������Y�߽�佃�󽝣�C ��h6��^�Rԉ��n��(�־|��#���/�77=�TW@��q8��}'��y�XL���Ѿ�����o����ž��bP�b�0�1�#>��?�|�6�t�$����VZ��S��7���	t�PxF�ys%�e[����>=�>�ཝR���b���J��o"��8B��Dn�w��l���B�b?��"�!E5��|?���>���3�:z ���	���!Ⱦ����5��
sξ������4%���6���?�\>�^�1�������X�۾@İ��F��>Mc��2:����m�����潜�߽��v�������A�+��jO����� ���Ǿ����M��)���9�?�@��:<��-�R�vU��ܾ���_���=��E�ؾn���Ď��+��;��@��;���+�����c��T�̾L��7���"T�m8/�\��B���!��o�߽Y��,��A��O��f6��^��Ӊ��n���־���#���/�/7=�*W@��q8��|'��x�xJ��ҵѾ~���*m����ž2���N����1��!>���?�p�6���$����X뾉R��r6�� t��vF�|r%��Z�p���H=�����S���	����K��q"��:B��Gn��x��*���3�s@�,�"�dF5��}?�!�>�4�3��{ �3�	�C��8�Ⱦ�"���8���uξ)�����5%��6���?��>���1������ʻ۾�İ��G���Oc�t5:�N���q�`�����߽]"�����������+�nO�j�������Ǿ_���N�:�)���9���@�i<<���-�9�wW�$�ܾ�������B���ؾ����a����+��;��  �  �0���+��b��W�0��0þVf���=��,W�[-5�8b�l�
������� ����z.�c*�M5!���;��1`��#���̦���˾Q��������!���-�U0�GP)��C�����i�z�ľ��������I�վ�-�����q#�L].�x0�$(��~��V��޾����씾��s�>�J���+�����B�L���!~�f��a���������l")���F�S�n�����
����~پ%���h�E�&��/��/�j
%�I�����1WپrU��ß��������CH��a�:<�<�'�"0��m.�p�#����p��iо/���t5���d�_?��#�q��FW�����D�)��C���3	�n�Z�1�:�R�[�~��ћ�达�v羐	��{���*�T�0���,�*��q�E�Uξ)����]���Գ��ʾ���1�$�Z�+�ە0��+�9b�W��.쾞/þ#e���<��4)W�.*5��^���
�������a����*��&�02!��;��/`�#��v̦�r�˾D��������!���-��T0��O)�WC�˨��g�P�ľ����g�������վ�*������o#�\.�Y0��"(�	~�V�,޾͏��{딾��s��J���+�@��aB�X����~��_�����d��l$)�O�F��n����ā����پ4��j���&�a�/�	/��%�������HZپ{X����������\���lJ��b��<���'��0�0n.���#���#q���iо꟪�n6����d�b?�~�#�>��Z[�4��jM���ｻ���7	�P�2���R���~�Cӛ��龾gx羈	��|��*���0�,�,�����r�fI�Yξ;����a���س�9�ʾ��G3�w%���+��  �  ���h����n����%ؾ��������N2���3`�B�<�*�}����u��ȗ�^���w�SF�!P/�J&H���g���8�ڒ��=�߾�y �5��`��.��n���R�)�̾O��ʛ�� t���V�����t�޾�Z �����/��"���E�a����̾����~���x��SU�#�9��$����	�T`����"��{��"�A�6�h�Q��Pt� ʏ��L���Tɾ��H���x�&^�����D�K%�����¾�Y����������׮�hTɾJF꾄����@|��v���Q:��n��¾���<���l�k�XMK���1�����ҋ��� *���
�(�5Y(��%?�Ex\��؀�V��3���gԾ~���j
�~������S��X��
�׾gv��f���+霾�2��x�����Ӿ���F�
�������g����*����$ؾ����S����0���0`��B���*������+��s�����s��B��L/�g#H�B�g�7���젾~����߾�y �)��E�������eR�����̾M��t���}q��CT��e�����޾oY ��������$���D�ɰ�\�̾L����}��J�x��RU�/�9�\$����	��`���#��|�~"�<�6���Q��St��ˏ�;N��iVɾ3��i���y�s_����cF��&�����¾�\��j�������ڮ��VɾH�;������|��v�0��:� o㾐¾����T���!�k��PK�:�1�� �j��K��s���.���Z�,](��)?��{\��ڀ�����4��9iԾY���k
������b����F\��Ɖ׾Bz��Nä�
휾�6�������Ӿ �����
�����  �  �n���������ܾ�{ž����ٚ��P��m?t���Y���B�A/�h4 �v�|~�����
#���2��\G��J_�R�z���������ܳ�U�ʾdh� ����\ �������7侟�ʾ�l�������z��U��������������,>پIG����e��3�������Ծ�ѽ������������j���Q���;��)��z�}{����b���'��U9���N�	�g�K��R���Y���9J��^Ҿ�k�h����<�� �od�ܾP���7v���7���`������{ǘ�����՜Ǿ[��FQ���� �� �_�����9;�P���G��$�����}��$b���I�s5���$�n����Px�3��9-�r!@��V��q�����ZĘ�,���[�¾� ھ�����&}�����˶�+tӾ�߸��.���Đ�3�������I)��k�о�K�
J���m�Z������Ȁܾ�zž`��Gؚ�wO��Y<t�4�Y��}B�/� 0 ����y���7#���2��XG�kG_���z�����4��vܳ���ʾ(h�ƿ��b\ �O�����6�2�ʾ�j������Xx�������S��������;پ�D�I���d�2��֧�?�Ծfн�����������j���Q��;�ҁ)��z��{�7��c�?�'�oW9���N�Th��L��м�����L��`Ҿ&n�ƾ���=�'
 �6g��ܾ6���y���:��Bc��B����ɘ�������Ǿɐ�eR��d� �8� ������㾶9;�Q���H��bᎾ��}�}(b���I��5�=�$��r�ƞ�}�����"-��%@���V�q�T����Ř�������¾�ھv������g~�a����뾀wӾM㸾,2��uȐ�ދ�������S��N�оTN�GL���  �  ؆վ�վ�Ͼɫž 	���V��I	���˗�	��9��u�f�TFO�^_<�N0��,�^K2��@�+T��l�b���Î��Q��}����簾���cȾ�sѾ.G־�{ԾC7˾�t���㧾 ���ns�E�o���|��<���螾���:�ľ�FѾDc־GLԾ�̾A������퇪��N��)������@/w�qx^��XH�*z7�Q.�b�-��6��)F���[��bt�Ұ��⫒����WD���ȴ�����=�˾M�Ӿx{־5ҾM�ƾ�-��	!������)�F;p�#%r�G��?��/���Yg���ɾ��Ӿ�n־,AҾKɾI���P1���Ħ�/���������n� �V��B��l3���,�ds/��:�:�L��c��|�G�J����ɡ�5��<���djľf�ξ<Pվ@�վ�Ͼ>I�������~��e����kx��n��v�?톾�U��6a��Be��1�;�վ_�վ��Ͼ��ž���qU����Qʗ�m�����i�f��AO��Z<�"I0��,�_F2�@��&T��l���������TP�������氾�����ȾHsѾ�F־;{Ծl6˾�s��t⧾f������is���o���|�:��W枾�����ľgDѾKa־xJԾI�̾����e��φ���M��b���,��[.w��w^�vXH�6z7��.��-��6�+F�f�[��dt�����.���j���E��pʴ�����a�˾��Ӿ�}־�7Ҿ��ƾz0���#��Z!��D/��@p�*r�\I��>��碥��h���ɾ��Ӿ�o־�AҾ�Kɾ���?2���Ŧ����������[�n�گV��B��q3���,�nx/�ɧ:���L�S�c���|�
Ċ�膖�pˡ��������lľ7�ξJRվ��վ�ϾL��ܟ��D���Σ��qrx���n�ϓv�q����X���c���g��O�;�  �  �V����������ڹ��չ����8l��y𰾹���������M!z���`��AP�w]K� S���e��G��my���������v���4��I��<幾�Ĺ�\�������M���[إ��������uu�wS]��N�L�K��kU�7�i��������R���ƫ�K|��г��:u���깾o����a��e����L���أ��,������p��Z�p;M���L��#X��n��@������_v�� R��g�� ��>���깾��������X��Ь��������vh��g�l��/W��9L���M��%[�jr��ʇ����������Į��<��g�� ����蹾g�������&��#;��V���7)���遾Xmh�ǏT���K�
O�lo^�~�v�sX���j���{��������1θ��ɹ��๾u6��M����� ����S��͜��9�~�k{d��<R�%HK�i�P��a�H�{�茾�ț�1Y���T��=������pٹ��Թ������j��ﰾ	���� ������z���`�W<P�XK���R�S�e�+E��w�����'���u���3��(H���乾�ù�Ե���������uץ�����s~���qu��O]�	�N� �K�xgU���i�o���� ���P���ī�mz������s�� 鹾4����`��}����K��Tأ�*,������p��Z��;M�;�L�}$X��n��A��x���|w��gS���h���!�����칾����������~Ҭ�Lá����� k����l�5W��>L�Q�M�*[��mr�<̇�k���Ά���Ů�_=��4���ӵ���鹾#h������(��=�������+��.쁾�rh�L�T��K�hO��t^�G w��Z���l���}�����v����ϸ�6˹�y⹾ 8��/���������V������S�~���d�CR��NK���P�b�ܷ{��ꌾ˛�0[���  �  �m��p���G���V���Jƾh$оk�վMվiC;�o���D���F�����1�u�Wo�
ty������廯�48¾F�Ͼ+־�վ�8ξ,�þn���m��2,���㕾^���a{��|b���K���9�/��-��4�wC�!�W��7p�{���~����1��e��?ײ�������ɾH�Ҿ�z־!tӾ��Ⱦ]��q����������L�q�R�p�:�����FA���@��_eǾ��Ҿ��־�WӾ�˾�쿾�!��i���o��T��� ����r���Z��E��U5��b-��f.�2:8�tI���_���x�I���Z����퟾P)�����7�¾0;��Ծ"L־��о�ľ\��ʝ�N��
�{��Yo�t�ۃ��7(��z���t����˾I�Ծ�)־EѾZ�Ǿ� ��sA���夾宙����y݁��j���R�W?�B�1�s�,���0�!>=�~uP� �g�qy��Č�l�����	���3����Hƾ:#о�վ�Kվ�A;�m��aB��ND�����r�u�oo�ny����ꖛ�U����5¾C�Ͼy־sվg7ξH�þ���=m��+���╾k��a_{�zb���K��9�./��-��	4�/C���W��3p�z�������%0��uc���ղ�[�����ɾA�Ҿ�y־hsӾ%�Ⱦ]��-���u��������q���p��:��K��B���A��xfǾ��Ҿf�־2YӾ�˾��#������Iq�����2��� s���Z��E��Z5��g-�3k.�`>8�FxI���_���x�����m����=*�����N�¾P1;?�Ծ�M־��оFľ�ﱾm͝��P����{��_o��$t������*������v����˾��Ծb+־�Ѿ��Ǿ2���B��?社ٰ�����߁�i�j�n�R�8?�?�1�l�,�w�0��C=��zP���g��{���Ō��  �  �9���曾�:����ƾ �ݾ(���d���_����M�
Ͼd����ڝ�����K���Pr��[���U����Ծ��쾳Y��#�%.�����ؾ8����|������򡆾y�o�#�U��>�4,�C��4�۵�H��AX%� 6��K��c�Ԑ��ԏ��a������@�ξC�侜[���� �K� ��a���5�T ƾ�^���ٗ�dF��I�����'���t&þ�uݾHk��A �s"�"���I�3ѾH	��ߙ������Mr����f��M��<8�4�&�m��s��H����6b*��<���R�s�l�Z���8��� )�����5־~�������q�����S+���׾�=��к��ے�2̊�����l˱�^̾�徚����3�m' �`��i1��Xɾ���������y���]�F���1�2I"��*�q�Fm�'� ��/���C��[���u��7��W图�9��i�ƾ�ݾ���oc��_�F���)辛
Ͼ�����ם��������o���W���R����Ծ��wW��/~��,�����ھؾS���|��'������y�o�ϒU�k�>�r1,��?�1����F��1T%��6��K��c�8��ӏ�5`�������ξ!�侟Z��$� �� �%a��^5� ƾ�^��ڗ��F������~������<'þ{vݾ\l�`B �$#������J�Ѿ=���������t��j�f��M��A8��&�8����������e*�R�<���R��l�~ᄾF���
*��%���6־��뾖����r�F����-ﾛ�׾�@������Jޒ�Wϊ���⿛�α��̾��h���t4�( ����2�Zɾp����������y��]�"F��1��N"�g0��v��r�`� �� 0�$�C��[�c�u��  �  �c���o���U���ھ����������� �ZT�|�	����Ҿ3@������������򺾽`پ7�����h�=��\���	�kE��o�Ҿi���/����g�g�Z���=�GC'��I�J~
�������l��;h��L3���L��n��ۋ�������þQP�\��������N��"����a��Ǿ��������N���l��QľH����c��"���-����[�����Ǿ�����u�� .r��3P�/�5�P!����Ŵ�$�����}	�Ե�%�+�:�wW�L�z�9ޓ��0����ξ��h�P��������>�X���}ݾ/����_��b>���/��T���܆ξ���%�^X�������,��+��a�ݾ�ϼ�i���І� �e���F�,.��Z���Ȇ�]��]��;��ј�^�+�#�C�+b�kb���n��{T���ھ������������eS�^�	�+���Ҿ=���|������������]پ4��[��0�1��|�B�	�7D��j�Ҿ}���I����e�Q�Z�T�=��@'� G�{
�
��ۿ����Xd�6��3���L�i n�9ڋ������þO���=��9���N��"�����a�̣Ǿū�����N��'m���Qľ��k	�������8.�a��.�����Ǿ´���w���2r�)8P��5�!�P��h�����/����	�t��S%��:�W���z�Zߓ��1��*�ξF��2�=���ܽ�@�a����ݾ����Kc���A���2��T�����ξ3��#&�FY����������,����ݾѼ�pj��s҆���e�ʙF��.��_�?��	��������*��p����+��C��b��  �  ����	8���Zž/��M}�TO�H,�2�0�U+�$3��
���뾬Oɾ�����u��Q����о�}�����{� �.$-��u0�3*�[�����徍̼�i���|���P�*v0�=���s�a$������l����������%��.A�kVg��ƌ�9���өҾ�����2�br$���.�}�/�I'��3��>�	C߾�H���������Z���^J۾� �Y�%�%��R/�_/�z�%��Y��� �-4׾������9El�y�D�Q�'�4���7�i$��'��}���U��H�����>r-���L�ףv����������p�0�����b�(�70�7�-�}�"�O�����X�Ӿw˸��¬��p��>!ƾ�羭��8A���)��p0�9-��!�~���L󾃺ɾ=ꤾ�����]�":����NG��� �\F���e9�_����S��~�6��\Y�����6���Yž'���|��N�mG,�a�0�Z+��1��
����tLɾ|���Jr������nоZz����� ��"-��t0�A*����r���徍˼�r���|���P��s0�����p�����{ｏe������^��>%�V+A�Sg�EŌ�Ď���ҾV���2��q$�o�.�(�/��H'��3��>��B߾�H���������Ԝ���J۾g� �����%�qS/��_/�8�%��Z�x� �6׾����'����Il���D���'����m<�v-�������]�����/��0u-�N�L�O�v���������@r���x��^�(�@80���-���"����|���ִӾ�θ�>Ƭ� t��Z$ƾ������NB���)�hq0��9-�!����M󾭻ɾ�뤾����"�]�	&:����K��� �`P���;C����V��b��#�6��_Y��  �  ք���� %Ͼ���B���,�\�;���@��y:��*��K��d��r�־����Ӷ��3¾�޾����V�Z�.���<��t@��9��n(�
��VU�Siž2��e}�2!M�;3*�١�� ���콱���߽{��9&��U_	��(��'<���e�
�� ���QL޾	/����3�2���>���?�x(6��$�����n��̾���ې���ɾ����3�!��4�7?�Z1?��l4�c!���	��x㾹o��⠒�Atk�<'@��� ��H�{���2��Y�z�k����k�2�&�-�H���v� ��'�������K��%&�Ц7��+@�´=�e�0�6���[��k�ľ�)���^��AhӾ,�������(��%9��u@�;�<�E�.��������Ծ:L���"��]�[��4����h����Y併v߽+]�V~���KQ�T�0�g�V��Ԅ�T���#Ͼ��B�3�,���;���@��x:���*�cJ��a��#�־D��0ж�0¾I�޾:��<U���.�'�<��s@� 9��m(�Z��)T�Ehž0��Y}�M��0*�2��"� ��������߽5������[	�%��$<�Z�e��������K޾r.�b����2�/�>���?�5(6�t$����gn��̾7���1���{�ɾ� �p���!��4��7?�2?��m4��c!���	��z㾲q�������xk��+@�k� ��M�������#ཬ����Tn�''��H�Y�v�X!��e���7L�s&&�է7��,@��=���0��������	�ľH-��Kb��pkӾ���N��ӛ(��&9��v@�۸<���.�%��S��� ԾM��9$����[�Ð4�$��������Xc�s�߽�f㽀���>U���0���V��  �  �~�����g�Ҿ����6���1�;A��kF��@���/�9R����۾�¾�{��EGƾ���P��ڐ�64��jB�9EF��>��'-�K��ɡ��ʸȾ{�����}�0OL��f(�6`��,��)�e]ݽ�w۽23�t���W���:���e����~��T�� m
��8#�s�7��9D�A�E�H�;�4�(�_��1��^ѾJ^��>I���Gξ������4&�[�9�X�D���D���9�9�%��A�p�'��yӓ��k�k�>����5�������y��۽�ܽ�u�h?���"� %�r�G��w�џ����þ�����\�*�=���E�ggC�#6��$!��{	����Y�Ⱦ�Ժ�N;��'ؾ������>i-�]�>��FF��\B�*�3��������ؾGv���눾�,[�23�\���d�R����߽r۽��޽������ ��T/�]
V�J}�����Y�Ҿ��o6�c�1�^:A�"kF��@���/��P������۾�¾	x���Cƾ�㾊��.��� 4�KiB�DF��>��&-����������Ⱦv�����}��LL��d(��]��&���"轰Vݽ�p۽�+��l�-���!�:�x�e�����}���⾊l
�K8#���7�d9D��E��;��(��^��1��^Ѿ{^���I��6HξB��[���4&���9���D�W�D�S�9��%�zB�J�)���Փ�5�k���>�c������������}�۽8�ܽ[}�~F���%�#%�)�G�u�w�����þ���>�*�=���E��hC��	6�^&!��}	�A����Ⱦtغ��>��\"ؾ�������Xj-�H�>�^GF�4]B���3���A��ؾ�w��G툾	0[��3����Vi�����߽)۽7�޽���)��p$�1X/�vV��  �  ք���� %Ͼ���B���,�\�;���@��y:��*��K��d��r�־����Ӷ��3¾�޾����V�Z�.���<��t@��9��n(�
��VU�Siž2��e}�2!M�;3*�١�� ���콱���߽{��9&��U_	��(��'<���e�
�� ���QL޾	/����3�2���>���?�x(6��$�����n��̾���ې���ɾ����3�!��4�7?�Z1?��l4�c!���	��x㾹o��⠒�Atk�<'@��� ��H�{���2��Y�z�k����k�2�&�-�H���v� ��'�������K��%&�Ц7��+@�´=�e�0�6���[��k�ľ�)���^��AhӾ,�������(��%9��u@�;�<�E�.��������Ծ:L���"��]�[��4����h����Y併v߽+]�V~���KQ�T�0�g�V��Ԅ�T���#Ͼ��B�3�,���;���@��x:���*�cJ��a��#�־D��0ж�0¾I�޾:��<U���.�'�<��s@� 9��m(�Z��)T�Ehž0��Y}�M��0*�2��"� ��������߽5������[	�%��$<�Z�e��������K޾r.�b����2�/�>���?�5(6�t$����gn��̾7���1���{�ɾ� �p���!��4��7?�2?��m4��c!���	��z㾲q�������xk��+@�k� ��M�������#ཬ����Tn�''��H�Y�v�X!��e���7L�s&&�է7��,@��=���0��������	�ľH-��Kb��pkӾ���N��ӛ(��&9��v@�۸<���.�%��S��� ԾM��9$����[�Ð4�$��������Xc�s�߽�f㽀���>U���0���V��  �  ����	8���Zž/��M}�TO�H,�2�0�U+�$3��
���뾬Oɾ�����u��Q����о�}�����{� �.$-��u0�3*�[�����徍̼�i���|���P�*v0�=���s�a$������l����������%��.A�kVg��ƌ�9���өҾ�����2�br$���.�}�/�I'��3��>�	C߾�H���������Z���^J۾� �Y�%�%��R/�_/�z�%��Y��� �-4׾������9El�y�D�Q�'�4���7�i$��'��}���U��H�����>r-���L�ףv����������p�0�����b�(�70�7�-�}�"�O�����X�Ӿw˸��¬��p��>!ƾ�羭��8A���)��p0�9-��!�~���L󾃺ɾ=ꤾ�����]�":����NG��� �\F���e9�_����S��~�6��\Y�����6���Yž'���|��N�mG,�a�0�Z+��1��
����tLɾ|���Jr������nоZz����� ��"-��t0�A*����r���徍˼�r���|���P��s0�����p�����{ｏe������^��>%�V+A�Sg�EŌ�Ď���ҾV���2��q$�o�.�(�/��H'��3��>��B߾�H���������Ԝ���J۾g� �����%�qS/��_/�8�%��Z�x� �6׾����'����Il���D���'����m<�v-�������]�����/��0u-�N�L�O�v���������@r���x��^�(�@80���-���"����|���ִӾ�θ�>Ƭ� t��Z$ƾ������NB���)�hq0��9-�!����M󾭻ɾ�뤾����"�]�	&:����K��� �`P���;C����V��b��#�6��_Y��  �  �c���o���U���ھ����������� �ZT�|�	����Ҿ3@������������򺾽`پ7�����h�=��\���	�kE��o�Ҿi���/����g�g�Z���=�GC'��I�J~
�������l��;h��L3���L��n��ۋ�������þQP�\��������N��"����a��Ǿ��������N���l��QľH����c��"���-����[�����Ǿ�����u�� .r��3P�/�5�P!����Ŵ�$�����}	�Ե�%�+�:�wW�L�z�9ޓ��0����ξ��h�P��������>�X���}ݾ/����_��b>���/��T���܆ξ���%�^X�������,��+��a�ݾ�ϼ�i���І� �e���F�,.��Z���Ȇ�]��]��;��ј�^�+�#�C�+b�kb���n��{T���ھ������������eS�^�	�+���Ҿ=���|������������]پ4��[��0�1��|�B�	�7D��j�Ҿ}���I����e�Q�Z�T�=��@'� G�{
�
��ۿ����Xd�6��3���L�i n�9ڋ������þO���=��9���N��"�����a�̣Ǿū�����N��'m���Qľ��k	�������8.�a��.�����Ǿ´���w���2r�)8P��5�!�P��h�����/����	�t��S%��:�W���z�Zߓ��1��*�ξF��2�=���ܽ�@�a����ݾ����Kc���A���2��T�����ξ3��#&�FY����������,����ݾѼ�pj��s҆���e�ʙF��.��_�?��	��������*��p����+��C��b��  �  �9���曾�:����ƾ �ݾ(���d���_����M�
Ͼd����ڝ�����K���Pr��[���U����Ծ��쾳Y��#�%.�����ؾ8����|������򡆾y�o�#�U��>�4,�C��4�۵�H��AX%� 6��K��c�Ԑ��ԏ��a������@�ξC�侜[���� �K� ��a���5�T ƾ�^���ٗ�dF��I�����'���t&þ�uݾHk��A �s"�"���I�3ѾH	��ߙ������Mr����f��M��<8�4�&�m��s��H����6b*��<���R�s�l�Z���8��� )�����5־~�������q�����S+���׾�=��к��ے�2̊�����l˱�^̾�徚����3�m' �`��i1��Xɾ���������y���]�F���1�2I"��*�q�Fm�'� ��/���C��[���u��7��W图�9��i�ƾ�ݾ���oc��_�F���)辛
Ͼ�����ם��������o���W���R����Ծ��wW��/~��,�����ھؾS���|��'������y�o�ϒU�k�>�r1,��?�1����F��1T%��6��K��c�8��ӏ�5`�������ξ!�侟Z��$� �� �%a��^5� ƾ�^��ڗ��F������~������<'þ{vݾ\l�`B �$#������J�Ѿ=���������t��j�f��M��A8��&�8����������e*�R�<���R��l�~ᄾF���
*��%���6־��뾖����r�F����-ﾛ�׾�@������Jޒ�Wϊ���⿛�α��̾��h���t4�( ����2�Zɾp����������y��]�"F��1��N"�g0��v��r�`� �� 0�$�C��[�c�u��  �  �m��p���G���V���Jƾh$оk�վMվiC;�o���D���F�����1�u�Wo�
ty������廯�48¾F�Ͼ+־�վ�8ξ,�þn���m��2,���㕾^���a{��|b���K���9�/��-��4�wC�!�W��7p�{���~����1��e��?ײ�������ɾH�Ҿ�z־!tӾ��Ⱦ]��q����������L�q�R�p�:�����FA���@��_eǾ��Ҿ��־�WӾ�˾�쿾�!��i���o��T��� ����r���Z��E��U5��b-��f.�2:8�tI���_���x�I���Z����퟾P)�����7�¾0;��Ծ"L־��о�ľ\��ʝ�N��
�{��Yo�t�ۃ��7(��z���t����˾I�Ծ�)־EѾZ�Ǿ� ��sA���夾宙����y݁��j���R�W?�B�1�s�,���0�!>=�~uP� �g�qy��Č�l�����	���3����Hƾ:#о�վ�Kվ�A;�m��aB��ND�����r�u�oo�ny����ꖛ�U����5¾C�Ͼy־sվg7ξH�þ���=m��+���╾k��a_{�zb���K��9�./��-��	4�/C���W��3p�z�������%0��uc���ղ�[�����ɾA�Ҿ�y־hsӾ%�Ⱦ]��-���u��������q���p��:��K��B���A��xfǾ��Ҿf�־2YӾ�˾��#������Iq�����2��� s���Z��E��Z5��g-�3k.�`>8�FxI���_���x�����m����=*�����N�¾P1;?�Ծ�M־��оFľ�ﱾm͝��P����{��_o��$t������*������v����˾��Ծb+־�Ѿ��Ǿ2���B��?社ٰ�����߁�i�j�n�R�8?�?�1�l�,�w�0��C=��zP���g��{���Ō��  �  �V����������ڹ��չ����8l��y𰾹���������M!z���`��AP�w]K� S���e��G��my���������v���4��I��<幾�Ĺ�\�������M���[إ��������uu�wS]��N�L�K��kU�7�i��������R���ƫ�K|��г��:u���깾o����a��e����L���أ��,������p��Z�p;M���L��#X��n��@������_v�� R��g�� ��>���깾��������X��Ь��������vh��g�l��/W��9L���M��%[�jr��ʇ����������Į��<��g�� ����蹾g�������&��#;��V���7)���遾Xmh�ǏT���K�
O�lo^�~�v�sX���j���{��������1θ��ɹ��๾u6��M����� ����S��͜��9�~�k{d��<R�%HK�i�P��a�H�{�茾�ț�1Y���T��=������pٹ��Թ������j��ﰾ	���� ������z���`�W<P�XK���R�S�e�+E��w�����'���u���3��(H���乾�ù�Ե���������uץ�����s~���qu��O]�	�N� �K�xgU���i�o���� ���P���ī�mz������s�� 鹾4����`��}����K��Tأ�*,������p��Z��;M�;�L�}$X��n��A��x���|w��gS���h���!�����칾����������~Ҭ�Lá����� k����l�5W��>L�Q�M�*[��mr�<̇�k���Ά���Ů�_=��4���ӵ���鹾#h������(��=�������+��.쁾�rh�L�T��K�hO��t^�G w��Z���l���}�����v����ϸ�6˹�y⹾ 8��/���������V������S�~���d�CR��NK���P�b�ܷ{��ꌾ˛�0[���  �  ؆վ�վ�Ͼɫž 	���V��I	���˗�	��9��u�f�TFO�^_<�N0��,�^K2��@�+T��l�b���Î��Q��}����簾���cȾ�sѾ.G־�{ԾC7˾�t���㧾 ���ns�E�o���|��<���螾���:�ľ�FѾDc־GLԾ�̾A������퇪��N��)������@/w�qx^��XH�*z7�Q.�b�-��6��)F���[��bt�Ұ��⫒����WD���ȴ�����=�˾M�Ӿx{־5ҾM�ƾ�-��	!������)�F;p�#%r�G��?��/���Yg���ɾ��Ӿ�n־,AҾKɾI���P1���Ħ�/���������n� �V��B��l3���,�ds/��:�:�L��c��|�G�J����ɡ�5��<���djľf�ξ<Pվ@�վ�Ͼ>I�������~��e����kx��n��v�?톾�U��6a��Be��1�;�վ_�վ��Ͼ��ž���qU����Qʗ�m�����i�f��AO��Z<�"I0��,�_F2�@��&T��l���������TP�������氾�����ȾHsѾ�F־;{Ծl6˾�s��t⧾f������is���o���|�:��W枾�����ľgDѾKa־xJԾI�̾����e��φ���M��b���,��[.w��w^�vXH�6z7��.��-��6�+F�f�[��dt�����.���j���E��pʴ�����a�˾��Ӿ�}־�7Ҿ��ƾz0���#��Z!��D/��@p�*r�\I��>��碥��h���ɾ��Ӿ�o־�AҾ�Kɾ���?2���Ŧ����������[�n�گV��B��q3���,�nx/�ɧ:���L�S�c���|�
Ċ�膖�pˡ��������lľ7�ξJRվ��վ�ϾL��ܟ��D���Σ��qrx���n�ϓv�q����X���c���g��O�;�  �  �n���������ܾ�{ž����ٚ��P��m?t���Y���B�A/�h4 �v�|~�����
#���2��\G��J_�R�z���������ܳ�U�ʾdh� ����\ �������7侟�ʾ�l�������z��U��������������,>پIG����e��3�������Ծ�ѽ������������j���Q���;��)��z�}{����b���'��U9���N�	�g�K��R���Y���9J��^Ҿ�k�h����<�� �od�ܾP���7v���7���`������{ǘ�����՜Ǿ[��FQ���� �� �_�����9;�P���G��$�����}��$b���I�s5���$�n����Px�3��9-�r!@��V��q�����ZĘ�,���[�¾� ھ�����&}�����˶�+tӾ�߸��.���Đ�3�������I)��k�о�K�
J���m�Z������Ȁܾ�zž`��Gؚ�wO��Y<t�4�Y��}B�/� 0 ����y���7#���2��XG�kG_���z�����4��vܳ���ʾ(h�ƿ��b\ �O�����6�2�ʾ�j������Xx�������S��������;پ�D�I���d�2��֧�?�Ծfн�����������j���Q��;�ҁ)��z��{�7��c�?�'�oW9���N�Th��L��м�����L��`Ҿ&n�ƾ���=�'
 �6g��ܾ6���y���:��Bc��B����ɘ�������Ǿɐ�eR��d� �8� ������㾶9;�Q���H��bᎾ��}�}(b���I��5�=�$��r�ƞ�}�����"-��%@���V�q�T����Ř�������¾�ھv������g~�a����뾀wӾM㸾,2��uȐ�ދ�������S��N�оTN�GL���  �  ���h����n����%ؾ��������N2���3`�B�<�*�}����u��ȗ�^���w�SF�!P/�J&H���g���8�ڒ��=�߾�y �5��`��.��n���R�)�̾O��ʛ�� t���V�����t�޾�Z �����/��"���E�a����̾����~���x��SU�#�9��$����	�T`����"��{��"�A�6�h�Q��Pt� ʏ��L���Tɾ��H���x�&^�����D�K%�����¾�Y����������׮�hTɾJF꾄����@|��v���Q:��n��¾���<���l�k�XMK���1�����ҋ��� *���
�(�5Y(��%?�Ex\��؀�V��3���gԾ~���j
�~������S��X��
�׾gv��f���+霾�2��x�����Ӿ���F�
�������g����*����$ؾ����S����0���0`��B���*������+��s�����s��B��L/�g#H�B�g�7���젾~����߾�y �)��E�������eR�����̾M��t���}q��CT��e�����޾oY ��������$���D�ɰ�\�̾L����}��J�x��RU�/�9�\$����	��`���#��|�~"�<�6���Q��St��ˏ�;N��iVɾ3��i���y�s_����cF��&�����¾�\��j�������ڮ��VɾH�;������|��v�0��:� o㾐¾����T���!�k��PK�:�1�� �j��K��s���.���Z�,](��)?��{\��ڀ�����4��9iԾY���k
������b����F\��Ɖ׾Bz��Nä�
휾�6�������Ӿ �����
�����  �  �0���+��b��W�0��0þVf���=��,W�[-5�8b�l�
������� ����z.�c*�M5!���;��1`��#���̦���˾Q��������!���-�U0�GP)��C�����i�z�ľ��������I�վ�-�����q#�L].�x0�$(��~��V��޾����씾��s�>�J���+�����B�L���!~�f��a���������l")���F�S�n�����
����~پ%���h�E�&��/��/�j
%�I�����1WپrU��ß��������CH��a�:<�<�'�"0��m.�p�#����p��iо/���t5���d�_?��#�q��FW�����D�)��C���3	�n�Z�1�:�R�[�~��ћ�达�v羐	��{���*�T�0���,�*��q�E�Uξ)����]���Գ��ʾ���1�$�Z�+�ە0��+�9b�W��.쾞/þ#e���<��4)W�.*5��^���
�������a����*��&�02!��;��/`�#��v̦�r�˾D��������!���-��T0��O)�WC�˨��g�P�ľ����g�������վ�*������o#�\.�Y0��"(�	~�V�,޾͏��{딾��s��J���+�@��aB�X����~��_�����d��l$)�O�F��n����ā����پ4��j���&�a�/�	/��%�������HZپ{X����������\���lJ��b��<���'��0�0n.���#���#q���iо꟪�n6����d�b?�~�#�>��Z[�4��jM���ｻ���7	�P�2���R���~�Cӛ��龾gx羈	��|��*���0�,�,�����r�fI�Yξ;����a���س�9�ʾ��G3�w%���+��  �  ��@��;�O�+�,���d��y�̾|��M8���%T��;/���?F������Y�߽�佃�󽝣�C ��h6��^�Rԉ��n��(�־|��#���/�77=�TW@��q8��}'��y�XL���Ѿ�����o����ž��bP�b�0�1�#>��?�|�6�t�$����VZ��S��7���	t�PxF�ys%�e[����>=�>�ཝR���b���J��o"��8B��Dn�w��l���B�b?��"�!E5��|?���>���3�:z ���	���!Ⱦ����5��
sξ������4%���6���?�\>�^�1�������X�۾@İ��F��>Mc��2:����m�����潜�߽��v�������A�+��jO����� ���Ǿ����M��)���9�?�@��:<��-�R�vU��ܾ���_���=��E�ؾn���Ď��+��;��@��;���+�����c��T�̾L��7���"T�m8/�\��B���!��o�߽Y��,��A��O��f6��^��Ӊ��n���־���#���/�/7=�*W@��q8��|'��x�xJ��ҵѾ~���*m����ž2���N����1��!>���?�p�6���$����X뾉R��r6�� t��vF�|r%��Z�p���H=�����S���	����K��q"��:B��Gn��x��*���3�s@�,�"�dF5��}?�!�>�4�3��{ �3�	�C��8�Ⱦ�"���8���uξ)�����5%��6���?��>���1������ʻ۾�İ��G���Oc�t5:�N���q�`�����߽]"�����������+�nO�j�������Ǿ_���N�:�)���9���@�i<<���-�9�wW�$�ܾ�������B���ؾ����a����+��;��  �  ���������^�n�ɾ[:��MD��W"e�,9�L��_���V�ֽ�J8�������j�����
��v�½:yݽC�o��7�A��Ap�$��� ���о�Y�˂���F�����zu߾�ľ�+���O���R��T���/ϊ�'���5��GԾd�뾔����������%ܾ��������烾�SU�)�,��O�(��2ͽɷ����yC��hP���7�$WʽJ��Dc
���(�bJP�=���B���*K���8پ�ﾀ;��Ê�����־IM���Ƞ��}��p���n���?���M��J����ܾu�����l���߫�,-Ӿ~~��������u�O�F��!�8���!��Ž菲�r˧��~���!���鬽x���Gӽ}���~t�Ҷ4�g�_����rΧ� Xƾd���_��Z���{`���8�D�;Q������ˇ�6��!�������� �ʾQ�侟���������?]��ɾ 9��C���e��9�{��<�����ֽ�罽�0�����b����������½�sݽ�@������A��@p�ී�����оkY龏���	F��;��]t߾g�ľ�)���M��LP��Ш���̊�\$��3���Ծ���?���]������#ܾ$�������惾�QU��,�fN�C�1ͽyȷ����'D����@�����]Zʽ+�轋e
�8�(�]MP��ှ���6M�� ;پ|��>��|���{��־EP���ˠ�ŀ��C��Rq��OB���O�����^�ܾ���������R�뾒-Ӿ�~��T ���u�0�F��!� ��G(��Ž����jӧ������)����Iɻ��Nӽ�����w�(�4���_�I��;Ч��Yƾ���cb������c���;���;��x ���χ��9�������������7�ʾ��	���  �  '�����G�޾0ž3ܧ�>��j�b�p]8�L2�����t�ٽ�&��4c��8è�k������;����ŽOf�S���W�@���m��H���n���5˾�~�<󾯝��c���پ���^s���Z��ԁ���~����%͚�r�����ξt��9���1�����k�־p~���������S��I,�l��ｿSн@�������H��󦽌���@(���~ͽ)���<�Y|(���N��\~�Tњ�y>���Ծ���Þ��������� �Ѿ���PX�����8]�����K\��������m5׾����7�����t��	6ξp���Wo���s��yE��>!�U����㽡5Ƚõ��᪽����+��8�����`Wֽ�d��~��64���]�j
��"���d���+ܾ�	� ���{��\�=�ȾG���핾�/����}�%M����!��Eƾ"�޾f�����@��ĵ޾�
ž�ڧ�����b��Z8�w/�����Ìٽ����[������ec��[��s4��	�Ž~`ཡP�����@���m��H���n���5˾�~���5��������پ?���q���X���с���~�0��ʚ�������ξ������x/����뾤�־�|��g������S�@H,�$���ｄRн� �������I��_���|����*��Ɓͽ��?��~(���N�`~�.Ӛ��@���Ծ&��S�����������Ѿ
���I[������b�<����^��*���T���6׾��뾿8��r	����s6ξ䷱��o��]s��{E�A!�(��U��<Ƚ�ʵ��骽ᇦ��3��U������^ֽ�k����$:4�D�]���蔤�R���7-ܾB�������`��ɾ��w��3��\�}���祓��$��V	ƾ��޾˗��  �  gk�J�޾�+Ͼ!���	̞�hc���Q]�:o7��u����t�㽝w˽�\���F��ï�`���P��н&�H'�mw�j)?���f��݊�ʘ��0����aӾ�ι�B�۾�>ʾ&�������R����|u���p�\l��+X��n���O���վ������ھ�6Ⱦ��+%���z���O��,������Ĉڽ�@Ž����8����U��ox���^ý��׽����|��%)�zK���u��H��@���ž��ؾ�M��⾌�־z�¾Rʪ�¤��偾�q���s�/��lw���<����Ǿ _ھ&�㾷��Xվ����4~��्�	�k��*C���"���	�y��քҽ�㿽c����ٯ�A��������Fɽpi�{ ���9�3���X�α���图�µ���̾Ήݾ�X�%�߾��о]���������{��p��Jy�N܊�7��u^��.�ξ��޾`i侎�޾Q*Ͼ͉���ʞ�5b��vO]��l7��r�������Gp˽KU��?��$��������H��1н�꽮$�Pu��'?���f�E݊���������aӾ��<�x�۾�=ʾ��������D���*xu���p��i���U�����M��
վH�������ھ5Ⱦ����#����z� �O�s�,���������ڽ/@Ž����粰�KW��^z��Kaý��׽�����~�P()��|K�H�u��J��B��C�ž��ؾP㾭��V�־Z�¾?ͪ������灾j�q��s�q1���y���>���ǾC`ھ��\�ᾕXվ�����~��������k��,C�|�"���	�2��?�ҽ뿽����⯽����4���Nɽq཰~ �c����3�ڷX�v���i盾ĵ��̾)�ݾ�[��߾��о���Y���b�7�{�np�,Ry��ߊ����ua����ξ�޾�  �  �ɾ��žo���e��uҒ�O�|�:X�o9����q������޽�Rͽ&ý�D����Ľ�н/d㽀a��}���$��?���_��ۂ��u��绫�`Ǽ�:�Ǿ�ɾS�¾����~ݟ�:����#u��I`�~S\���i��^��節��&��۰���Ǿ�ɾ�~¾{峾۪���勾�p��3M�
0��o���n�Y	ؽhɽ�X�������ǽNֽ�6뽙����%-��I�	�k�����`��	챾00��R?ɾ�EȾ�F��O����R��twl�T�\�j�^��r�j��^���%���85��Oɾ�4Ⱦ�U��(ح�gƙ������c���B�ɕ'����Z �I��Eҽ��Ž�_��|n½��˽�Kܽ���t	��:��6��xT�A�x�M���o,�������ľ��ɾZ�žW>���������1?�{we�#�[��c��{��㏾Mo��.i����ľ�ɾ�ž�m��Ld��<ђ���|��7X��9����n�s���^�޽�Jͽ�ý�<����Ľ7�н�\��Z�������$�1�?�1�_�qۂ��u������Ǽ�݃Ǿ��ɾ��¾����ܟ�����u�UE`��N\���i�&\��q���;$��������Ǿښɾ�|¾�㳾X����䋾cp�2M��0��n�*��?��ؽzɽ1Y�����
�ǽ�ֽ�9뽂��2!��'-��I�M�k�˜��b��1�2���AɾHHȾ[I���Q�������T��}l���\�x�^�Fr�!l��!�������`6��Pɾ`5Ⱦ=V���ح� Ǚ������c��B�~�'����] ���iMҽj�Ž{h��@w½M�˽Tܽ���jx	�N>�6��{T�~�x�����B.������H�ľP�ɾ,�žnA��ص��"��qF��~e�p�[�"�c�ھ{��揾3r���k����ľ�  �  +����w��<���ܕ�*���Q�r���X��wA��$-�_:�6��a�����mhܽ��ؽek޽�콽���+��p1�w[F�1^���x�V֊��٘����'����-���楾���։��s���W���F���C���N���e�qt���撾���l9��0���Q���t���6���̂���i�d�P�\d:��&�
������H��?�㽗0ڽӭٽY4�3��T������$�c8���M���f�33���������s��}���Ԫ�Rb������NH��Wi���P��PD���E��PU�v�o�����}���̤�ѫ��ы���M���p���|��a���H�[�3�o� �{���n�����߽��ؽއ۽i��$'��`�	��[�+�w?�b�U�*�o�� ��rS��M��Lѩ�-���캨�TG���Q����}���_�+K�u=C�֚I��]��	z������ʜ�6ݧ�F���1v���:��eە�򜇾��r� �X��tA��!-��6�x��P���b�轖_ܽ��ؽ�b޽j���	�|���
n1�WYF�z/^�s�x��Պ��٘��������-���奾�����ԉ�5s���W���F�$�C���N�)�e�r��X䒾S��O7��8���3O��)s��5���˂�[�i���P��b:���&�&��/��6H��U��I1ڽ!�ٽD6⽼��EV����4�$��8���M���f��4������]u��偬�lת��d��i���K���i�D�P�VD���E�UUU�w�o�?������Τ�ҫ�_﫾|���,N���q���|��a�T�H�U�3��� �U��s����.�߽�ٽ�۽X�潫/��d�	��_��
+��?���U�N�o�}��/U��7��pө���������AJ��U��e�}���_�2K�fDC���I�$]��z�u���͜�eߧ��  �  ���F{��>�����D����ir��wc�?eT�q�D�#(4��r#���Ie�������� �
�	�'3�I'���7�W?H���W���f�R�u��g������������P���M���J����g�u�N��9���,�c5*��2�_tD��P\��u�EF���3��ӫ��赐�V?��J����u|�~im��z^��=O�u=?�k�.����V� %�����A1��*/����TK�5�,�kg=��M�E�\�v�k��z��ل����	[��nÑ�BΎ�TW����x�
#_���F��44�*�*���+��7���K���d�X�}�]���ޏ�iϑ�ꋏ��7��?:���mw�oh��uY�� J��9���(����!�Xt�GG�������<�=[�j�!�hF2�B�B�/�R�>�a�2�p�-���;��.x���C��aK��4̌�s���+Ip�*�V���?��/�5�)�I�.���=���S�Psm��ɂ�`�� ���y���	��� �����wgr�-uc�_bT�;�D��$4��n#�����`����x��� �m�	��.�P'�z�7�V<H��W���f���u�2g��U����� ���/P���L��~I���g�3�N�N�9���,�1*�m�2��oD�L\���u�#D��1��񩑾-����=��㧅�Vs|�Ygm��x^�K<O�I<?���.���V�%������2��0�����L��,��i=��M��\���k���z��ۄ�"���<]���ő��Ў��Y��3�x�Z(_���F�:4�+�*�L�+�f�7���K���d�=�}�P^���ߏ�CБ�����L8��;���ow�sqh��xY��J���9��(����%�By�*Q��{����A��_���!�=J2���B�s�R�U�a�8�p�B��Z=���y���E���M���Ό�1���Op�i�V�>�?���/���)���.���=�|�S��xm��˂�t���  �  ��t��i|�6������8������	|�vtt�d#h��fW�C�C��Q0����h���� ��T#�ă4�VH��q[�zJk��v�A}��<���ƀ����Q��� {�»r�*�e�kFT�"�@�BE-����/�����`���%�׻7�N�K�"\^��~m�v�w���}��a���ˀ�*�����Rz�M�p�q�b��Q��4=�>Q*�p�
�˔�T%�fi(�K�:���N�q*a��o�%;y��~�F��-ˀ�ju��k~�o�x�8�n�,;`��M�W�9��x'�����a��K���G+��N>�%R���c�ށq��hz��4�ș���ɀ��U���}��}w���l��b]�	�J�o�6�(�$��������=��?��B.���A��OU�
wf��Os�!u{��������l��,����|��v��j��mZ��4G��n3�51"��K���g��� ��U1���D��hX���h�j�t��f|����T��������_|�|qt� h�cW��C�aM0���P��������M	#�4��QH��m[�Gk���v��>}��;���ŀ�`������{�:�r�K�e�#DT�i�@�B-�d��P����x\�8�%���7��K�X^�{m���w���}�s`��9ʀ��������z���p�N�b�Q�4=�Q*�"p�\
�r��G&��j(�� ;���N��,a���o��=y���~�����̀�iw��Vo~���x���n�@`��M�r�9��}'����Sf�iP�@��K+�R>��'R� �c���q�jjz�M6������ʀ��V����}�ʀw���l�g]���J�W�6�M�$�9��7��
C��D�gG.��A��SU��zf��Rs�#x{����4����À��.����|��v���j�sZ�:G�yt3�A7"�R�4��
m�W� �;[1���D�;mX���h��  �  ?U�(Ld��?s��(���b���P��g����ߐ�A����.��~l�ϓR�$�<��#.���)�4�0���@��X���q�씄�K-���j��\&��.��nن���~�i�o�6�`�w�Q���A�NZ1�E� �V������*���z��F��o��"��_�)��:���J�>NZ�Di��Dx�J��������Ï��ё�����������|��pc��J�5�6�R|+���*��
5�SH���`�S�y��݇�L���ˑ�)+��p@��Kr���y�x�j�x�[�4�L��z<���+��j�_,�U�������=��ӣ������y/�	&@�mP�AO_��=n�L}����󏌾Oݐ�x���)ލ������~t���Z��@C�z�1�	*�8-�x�:���O��*i�N쀾J���̂����Ԏ�� ������^�t���e���V�	XG���6�|-&��Z��0	�DU ������X��{�� ���W$��5�P�E��;U�IId�5=s��'���a���O�����$ސ������,��l���R��<�-.�.�)���0��@��X�ǲq�����d+��i��%���,���؆���~���o���`���Q���A�X1��� �G��"��&#���r��9��S����^�)��:��J��JZ��@i��Ax�����������'ё�����H���֨|�]pc�עJ�F�6��|+�<�*�}5��H���`�'�y��އ����2͑��,��B��t����y���j���[�ʣL��<���+��o�D1�!��;����F������a��v|/��(@��P�GQ_��?n�N}����:����ސ�7���*���𸅾��t���Z�uFC��1��*�� -���:���O�j/i�R���h���e���"֎�4"�����u�t�"�e���V�U\G�_�6��2&��_�l6	�[ �	���c�����,��z\$�5��E��  �  .�B�/Z��St�Cl��k���4Ң��ª�+����h��Q	��(���;Jx�!�[���H�gUC��	L�qga�mr��;��-���$�������y��@f��#����4��=n��T�l�=�y�)�4t�+'	��������-۽�$ٽm3�F���'��]���!���4�&J�ub���}��=��G�� ��$��њ���9���2��y�� �m�I%T�PvE�H�D�4�Q�q�j��5��G���Q������c�����j���Ԏ��g��{Ue���L�z�6��#�������}�Zsٽ�xڽmr�Mv��������9�'��;���Q�c<k�:���������U���n����੾eg��w������bd��M�4�C�Z�G��Y�H�t�F���mv���j��R���H��'���X��Jhw���\��E�:W0���S���Y ����	�ݽ��ؽ��ܽX������U��&�b1.��B�q�Y�}Qt�k��A����Т�{��������f��:��Ж��Ex���[�#�H�kOC��L��aa��l�/9��� ��}"��˾��Bx���d������3��i;n�=�T���=�r�)��q��$	�����k��&۽7ٽ�+�q��$�Z�2�!��4��J�rb�ԧ}��<��-��
��R��#���9��S2��:����m�\%T��vE��D�$�Q���j��6��.���^������d��� ���k���֎��i���Ye�ʪL���6���#���Κ�M��D��J|ٽ9�ڽUz佊}�����q����'�7�;���Q��>k�W���M ���������V����⩾�i��!��ӊ���gd��M�+�C�%�G�HY�b�t���x���l���S��XJ��y���h�����%kw���\�}E�6[0�B����^ �>����ݽi�ؽ+�ܽv��R���Y��*��4.��  �  ��:�I Z���6���~~��EL���Gƾ��ɾ�Tľ;z��gN��H̎�	z�/�b���[�/�f�ǋ�� B��է��$���\ƾ��ɾ�Dľ������Z��vv�¢R��4�����d�8۽
 ˽�&½����>ƽ�2ӽ�5�F7�����(�c�D���e��6���ᮾ���_�Ⱦ@ɾ���-}���g��Z`���p�kc^�Ye]�_�m�KT�����b�������Ⱦ�ɾ
����밾n:���w����i���G�F�+���������+
ս�Lǽ���c���Ǿɽ�ٽWp���S��y�1���N��7r�F��͡��ڴ��þ�ɾ�4Ǿ�ڻ�3�������f����h�l\�`a�
�v�a�����������&þs�ɾ_ Ǿ����Ҩ��L�������]��=�D�#�\~��������Ͻ�NĽ\2���|ý ν�߽9���p��� �ǯ:��Z�����X}��K��FFƾ$�ɾ�Rľx���K���Ɏ�Hz��b�9�[�Ѓf����� ?��Fҧ�]"��xZƾ��ɾ�Bľ����o���X��Ctv��R��~4����}��^��2۽�˽�½�y���7ƽz+ӽ|.罝3������(�=�D���e�O5���욾�ா�����Ⱦ�ɾ�����|���g��A`��#�p��c^��e]�N�m��T��f��c�����ƔȾ	ɾ���P�(<���y����i���G���+�4 �Z��L��Rս�Uǽ���������ɽ�ٽ�v�ך�����1�0 O��9r�z��YΡ�jܴ��þ �ɾ7Ǿ*ݻ�	�������i����h��\�ra�ǻv����#��Ί��s(þ
�ɾ�!Ǿ�������AM��h���v�]�h�=���#�{��v���])�u�Ͻ�XĽ�<��Ɔý�ν��߽�����s�0!��  �  OT9�n�_�ھ��?���깾Bо�m߾�e�8޾R�;y��О�cމ�}Ex�:)p�%�|���;���b���
Ҿ�eྡྷE�d�ܾl�˾�]���u���^��XsV���1��/�������޽�AȽ�_���f�����e��W�����ӽ*h�&�
��4$�W6E��*n����𨾽���GI־�Q���㾉�پ>�ƾ�ா>���S��hBs�cr�䮂��Ԕ��'���"ľ��׾�⾪� ؾv{ľ�Ы�cݑ�]+s�a[I��w'��4��
�`cֽ�s½;�',��x䰽!��7ƽj�۽�����p��R.�[�Q��w}�����e���kɾBa۾��㾛_��Ծ� ��*����4��m���p��Tv�Lꇾ�:���P��Ii˾ �ܾ}=�#��,\Ҿš���$��{��#ed��.=�&������l�^�ν쁽��J��#���S������K�̽!�չ�@��sQ9��_������=���鹾�@оjl߾ d�H޾�;���J͞�Yۉ�?x��"p�|�|�������_���ҾmcྌC侞�ܾ��˾U\��{t���]��iqV���1��-�������޽<ȽWY��`���2������o�ӽaｺ�
��1$�H3E��'n�M�������]H־�P�X���پߟƾ�ா>���S���Bs�	r�[���UՔ�N(���#ľ��׾3���㾑ؾ	}ľ]ҫ�5ߑ�;/s�t_I�;|'�P9���^lֽ�|½����4���창�(��!>ƽ��۽����:s�U.���Q��y}�򔗾Ί���lɾ!c۾���bᾇԾy��O����7���s�
�p�/[v�C퇾�=��]S��pk˾��ܾ?侁��d]Ҿ좼��%��F|���gd��1=����~��.u�x�νp����T��廯�囲������̽ )�t��z���  �  �z:�y{e�P�������/�ƾ�߾�0�i������c�ݾ��ľ峩�`����]����}�3ᅾ ��h����zʾ��⾘��t���%C���ھdO���񢾵���J[��22�b���1��~�Խ�����z����7����T��˘����ɽ���.�#��G���u�m���Z����Ͼf��g}������Z��N�վ���TS��j��c����������f����z��Ӿ���S���H��7��іҾ靶��5��~{��iL�ʠ&�=�	�ڰ齷̽�B��W6��̦��w��`J���󻽿�ѽ�������9.�zV�񏃾����\��#0ؾ=��i����z���b;�z�����1Q��B.~��K���`��]ئ�X����+۾GY�׿��io�"V�K�ɾJɬ�ɷ��f�j�O�>�������޽��Ľ;t��Ƕ���Z���	��$��n;½b3۽gO��.���w:��xe�-�������ƾ��߾]/��������ݾ	�ľ���C���LZ����}��݅����*����wʾ3����J���LA�T�ھN���𢾪���J[��02�6��4-��H�Խ�񽽐t��	맽Z����M�������zɽ��彴*��#��G�!�u�'��xY���Ͼ�澡|��P��������վ���<S��"j������g��j��� ����{���Ӿ���HT���I�����`�Ҿ�����7��܁{��mL���&���	���齕&̽^K���>��jԦ�����Q������'�ѽb�񽧊�+<.��V�-���O�������1ؾ,��Ak��v��I���e;.~��d����T���4~��N���c��%ۦ�։��.۾$[�l����p�SW�h�ɾiʬ������j�T�>������޽��Ľy}��=���od��������C½,;۽vV��U���  �  35;�*�g�}ݎ�C�A˾���۝��͔��I���r��Zɾ���c����酾'H��&���~Y������g�Ͼr辁���g�����I]��ľ���)���]��2�k�� ��y�ѽ徺��T���褽�����<��kd���Rƽ���7�"�"���H�^�x�����3���ԾA���������o�!J۾����社ZE��5��c��Gd��p$���ݼ�,lؾ�ﾋ���������̼׾@��������~�Z�M���&������潓�ȽW�����2ɣ�,q���'��'���t�ν+@�����.���W�Uo��^����Z���ݾ��a��|#�����$�Ҿ�����ٜ������}��T΄�_��$���1<ƾs��Ǳ���i������\$�vξ�[������lm��?������ �Ө۽gT���D�������Z��s����ۮ�1��3ؽ1��@Z�o2;���g�\܎�,מּ�?˾}��n������G���p�>Xɾ)���?���7慾�D�����V��_���S~Ͼ:o�� ��Qe������[ྸ�ľ������]�	�2�=��a��D�ѽ6����N��V⤽Ē���5��S]���Kƽ��|4���"���H���x�S����1��ܵԾ[����������I۾�����椾eE��d��fc���d��%���޼�mؾ� ﾴ�������y��[�׾�������~�\�M�Ω&�#��M��e�Ƚ���#���ѣ�y��V/��¸�ٯνF�����.�a�W��p������P\����ݾ����
&�����9�Ҿ���Cݜ�5������ф�b��🪾�>ƾ��ྦ����k��7����%�5wξ�\�����Rom��?�3���� ���۽%]��N�����d������䮽����:ؽ0��`]��  �  �z:�y{e�P�������/�ƾ�߾�0�i������c�ݾ��ľ峩�`����]����}�3ᅾ ��h����zʾ��⾘��t���%C���ھdO���񢾵���J[��22�b���1��~�Խ�����z����7����T��˘����ɽ���.�#��G���u�m���Z����Ͼf��g}������Z��N�վ���TS��j��c����������f����z��Ӿ���S���H��7��іҾ靶��5��~{��iL�ʠ&�=�	�ڰ齷̽�B��W6��̦��w��`J���󻽿�ѽ�������9.�zV�񏃾����\��#0ؾ=��i����z���b;�z�����1Q��B.~��K���`��]ئ�X����+۾GY�׿��io�"V�K�ɾJɬ�ɷ��f�j�O�>�������޽��Ľ;t��Ƕ���Z���	��$��n;½b3۽gO��.���w:��xe�-�������ƾ��߾]/��������ݾ	�ľ���C���LZ����}��݅����*����wʾ3����J���LA�T�ھN���𢾪���J[��02�6��4-��H�Խ�񽽐t��	맽Z����M�������zɽ��彴*��#��G�!�u�'��xY���Ͼ�澡|��P��������վ���<S��"j������g��j��� ����{���Ӿ���HT���I�����`�Ҿ�����7��܁{��mL���&���	���齕&̽^K���>��jԦ�����Q������'�ѽb�񽧊�+<.��V�-���O�������1ؾ,��Ak��v��I���e;.~��d����T���4~��N���c��%ۦ�։��.۾$[�l����p�SW�h�ɾiʬ������j�T�>������޽��Ľy}��=���od��������C½,;۽vV��U���  �  OT9�n�_�ھ��?���깾Bо�m߾�e�8޾R�;y��О�cމ�}Ex�:)p�%�|���;���b���
Ҿ�eྡྷE�d�ܾl�˾�]���u���^��XsV���1��/�������޽�AȽ�_���f�����e��W�����ӽ*h�&�
��4$�W6E��*n����𨾽���GI־�Q���㾉�پ>�ƾ�ா>���S��hBs�cr�䮂��Ԕ��'���"ľ��׾�⾪� ؾv{ľ�Ы�cݑ�]+s�a[I��w'��4��
�`cֽ�s½;�',��x䰽!��7ƽj�۽�����p��R.�[�Q��w}�����e���kɾBa۾��㾛_��Ծ� ��*����4��m���p��Tv�Lꇾ�:���P��Ii˾ �ܾ}=�#��,\Ҿš���$��{��#ed��.=�&������l�^�ν쁽��J��#���S������K�̽!�չ�@��sQ9��_������=���鹾�@оjl߾ d�H޾�;���J͞�Yۉ�?x��"p�|�|�������_���ҾmcྌC侞�ܾ��˾U\��{t���]��iqV���1��-�������޽<ȽWY��`���2������o�ӽaｺ�
��1$�H3E��'n�M�������]H־�P�X���پߟƾ�ா>���S���Bs�	r�[���UՔ�N(���#ľ��׾3���㾑ؾ	}ľ]ҫ�5ߑ�;/s�t_I�;|'�P9���^lֽ�|½����4���창�(��!>ƽ��۽����:s�U.���Q��y}�򔗾Ί���lɾ!c۾���bᾇԾy��O����7���s�
�p�/[v�C퇾�=��]S��pk˾��ܾ?侁��d]Ҿ좼��%��F|���gd��1=����~��.u�x�νp����T��廯�囲������̽ )�t��z���  �  ��:�I Z���6���~~��EL���Gƾ��ɾ�Tľ;z��gN��H̎�	z�/�b���[�/�f�ǋ�� B��է��$���\ƾ��ɾ�Dľ������Z��vv�¢R��4�����d�8۽
 ˽�&½����>ƽ�2ӽ�5�F7�����(�c�D���e��6���ᮾ���_�Ⱦ@ɾ���-}���g��Z`���p�kc^�Ye]�_�m�KT�����b�������Ⱦ�ɾ
����밾n:���w����i���G�F�+���������+
ս�Lǽ���c���Ǿɽ�ٽWp���S��y�1���N��7r�F��͡��ڴ��þ�ɾ�4Ǿ�ڻ�3�������f����h�l\�`a�
�v�a�����������&þs�ɾ_ Ǿ����Ҩ��L�������]��=�D�#�\~��������Ͻ�NĽ\2���|ý ν�߽9���p��� �ǯ:��Z�����X}��K��FFƾ$�ɾ�Rľx���K���Ɏ�Hz��b�9�[�Ѓf����� ?��Fҧ�]"��xZƾ��ɾ�Bľ����o���X��Ctv��R��~4����}��^��2۽�˽�½�y���7ƽz+ӽ|.罝3������(�=�D���e�O5���욾�ா�����Ⱦ�ɾ�����|���g��A`��#�p��c^��e]�N�m��T��f��c�����ƔȾ	ɾ���P�(<���y����i���G���+�4 �Z��L��Rս�Uǽ���������ɽ�ٽ�v�ך�����1�0 O��9r�z��YΡ�jܴ��þ �ɾ7Ǿ*ݻ�	�������i����h��\�ra�ǻv����#��Ί��s(þ
�ɾ�!Ǿ�������AM��h���v�]�h�=���#�{��v���])�u�Ͻ�XĽ�<��Ɔý�ν��߽�����s�0!��  �  .�B�/Z��St�Cl��k���4Ң��ª�+����h��Q	��(���;Jx�!�[���H�gUC��	L�qga�mr��;��-���$�������y��@f��#����4��=n��T�l�=�y�)�4t�+'	��������-۽�$ٽm3�F���'��]���!���4�&J�ub���}��=��G�� ��$��њ���9���2��y�� �m�I%T�PvE�H�D�4�Q�q�j��5��G���Q������c�����j���Ԏ��g��{Ue���L�z�6��#�������}�Zsٽ�xڽmr�Mv��������9�'��;���Q�c<k�:���������U���n����੾eg��w������bd��M�4�C�Z�G��Y�H�t�F���mv���j��R���H��'���X��Jhw���\��E�:W0���S���Y ����	�ݽ��ؽ��ܽX������U��&�b1.��B�q�Y�}Qt�k��A����Т�{��������f��:��Ж��Ex���[�#�H�kOC��L��aa��l�/9��� ��}"��˾��Bx���d������3��i;n�=�T���=�r�)��q��$	�����k��&۽7ٽ�+�q��$�Z�2�!��4��J�rb�ԧ}��<��-��
��R��#���9��S2��:����m�\%T��vE��D�$�Q���j��6��.���^������d��� ���k���֎��i���Ye�ʪL���6���#���Κ�M��D��J|ٽ9�ڽUz佊}�����q����'�7�;���Q��>k�W���M ���������V����⩾�i��!��ӊ���gd��M�+�C�%�G�HY�b�t���x���l���S��XJ��y���h�����%kw���\�}E�6[0�B����^ �>����ݽi�ؽ+�ܽv��R���Y��*��4.��  �  ?U�(Ld��?s��(���b���P��g����ߐ�A����.��~l�ϓR�$�<��#.���)�4�0���@��X���q�씄�K-���j��\&��.��nن���~�i�o�6�`�w�Q���A�NZ1�E� �V������*���z��F��o��"��_�)��:���J�>NZ�Di��Dx�J��������Ï��ё�����������|��pc��J�5�6�R|+���*��
5�SH���`�S�y��݇�L���ˑ�)+��p@��Kr���y�x�j�x�[�4�L��z<���+��j�_,�U�������=��ӣ������y/�	&@�mP�AO_��=n�L}����󏌾Oݐ�x���)ލ������~t���Z��@C�z�1�	*�8-�x�:���O��*i�N쀾J���̂����Ԏ�� ������^�t���e���V�	XG���6�|-&��Z��0	�DU ������X��{�� ���W$��5�P�E��;U�IId�5=s��'���a���O�����$ސ������,��l���R��<�-.�.�)���0��@��X�ǲq�����d+��i��%���,���؆���~���o���`���Q���A�X1��� �G��"��&#���r��9��S����^�)��:��J��JZ��@i��Ax�����������'ё�����H���֨|�]pc�עJ�F�6��|+�<�*�}5��H���`�'�y��އ����2͑��,��B��t����y���j���[�ʣL��<���+��o�D1�!��;����F������a��v|/��(@��P�GQ_��?n�N}����:����ސ�7���*���𸅾��t���Z�uFC��1��*�� -���:���O�j/i�R���h���e���"֎�4"�����u�t�"�e���V�U\G�_�6��2&��_�l6	�[ �	���c�����,��z\$�5��E��  �  ��t��i|�6������8������	|�vtt�d#h��fW�C�C��Q0����h���� ��T#�ă4�VH��q[�zJk��v�A}��<���ƀ����Q��� {�»r�*�e�kFT�"�@�BE-����/�����`���%�׻7�N�K�"\^��~m�v�w���}��a���ˀ�*�����Rz�M�p�q�b��Q��4=�>Q*�p�
�˔�T%�fi(�K�:���N�q*a��o�%;y��~�F��-ˀ�ju��k~�o�x�8�n�,;`��M�W�9��x'�����a��K���G+��N>�%R���c�ށq��hz��4�ș���ɀ��U���}��}w���l��b]�	�J�o�6�(�$��������=��?��B.���A��OU�
wf��Os�!u{��������l��,����|��v��j��mZ��4G��n3�51"��K���g��� ��U1���D��hX���h�j�t��f|����T��������_|�|qt� h�cW��C�aM0���P��������M	#�4��QH��m[�Gk���v��>}��;���ŀ�`������{�:�r�K�e�#DT�i�@�B-�d��P����x\�8�%���7��K�X^�{m���w���}�s`��9ʀ��������z���p�N�b�Q�4=�Q*�"p�\
�r��G&��j(�� ;���N��,a���o��=y���~�����̀�iw��Vo~���x���n�@`��M�r�9��}'����Sf�iP�@��K+�R>��'R� �c���q�jjz�M6������ʀ��V����}�ʀw���l�g]���J�W�6�M�$�9��7��
C��D�gG.��A��SU��zf��Rs�#x{����4����À��.����|��v���j�sZ�:G�yt3�A7"�R�4��
m�W� �;[1���D�;mX���h��  �  ���F{��>�����D����ir��wc�?eT�q�D�#(4��r#���Ie�������� �
�	�'3�I'���7�W?H���W���f�R�u��g������������P���M���J����g�u�N��9���,�c5*��2�_tD��P\��u�EF���3��ӫ��赐�V?��J����u|�~im��z^��=O�u=?�k�.����V� %�����A1��*/����TK�5�,�kg=��M�E�\�v�k��z��ل����	[��nÑ�BΎ�TW����x�
#_���F��44�*�*���+��7���K���d�X�}�]���ޏ�iϑ�ꋏ��7��?:���mw�oh��uY�� J��9���(����!�Xt�GG�������<�=[�j�!�hF2�B�B�/�R�>�a�2�p�-���;��.x���C��aK��4̌�s���+Ip�*�V���?��/�5�)�I�.���=���S�Psm��ɂ�`�� ���y���	��� �����wgr�-uc�_bT�;�D��$4��n#�����`����x��� �m�	��.�P'�z�7�V<H��W���f���u�2g��U����� ���/P���L��~I���g�3�N�N�9���,�1*�m�2��oD�L\���u�#D��1��񩑾-����=��㧅�Vs|�Ygm��x^�K<O�I<?���.���V�%������2��0�����L��,��i=��M��\���k���z��ۄ�"���<]���ő��Ў��Y��3�x�Z(_���F�:4�+�*�L�+�f�7���K���d�=�}�P^���ߏ�CБ�����L8��;���ow�sqh��xY��J���9��(����%�By�*Q��{����A��_���!�=J2���B�s�R�U�a�8�p�B��Z=���y���E���M���Ό�1���Op�i�V�>�?���/���)���.���=�|�S��xm��˂�t���  �  +����w��<���ܕ�*���Q�r���X��wA��$-�_:�6��a�����mhܽ��ؽek޽�콽���+��p1�w[F�1^���x�V֊��٘����'����-���楾���։��s���W���F���C���N���e�qt���撾���l9��0���Q���t���6���̂���i�d�P�\d:��&�
������H��?�㽗0ڽӭٽY4�3��T������$�c8���M���f�33���������s��}���Ԫ�Rb������NH��Wi���P��PD���E��PU�v�o�����}���̤�ѫ��ы���M���p���|��a���H�[�3�o� �{���n�����߽��ؽއ۽i��$'��`�	��[�+�w?�b�U�*�o�� ��rS��M��Lѩ�-���캨�TG���Q����}���_�+K�u=C�֚I��]��	z������ʜ�6ݧ�F���1v���:��eە�򜇾��r� �X��tA��!-��6�x��P���b�轖_ܽ��ؽ�b޽j���	�|���
n1�WYF�z/^�s�x��Պ��٘��������-���奾�����ԉ�5s���W���F�$�C���N�)�e�r��X䒾S��O7��8���3O��)s��5���˂�[�i���P��b:���&�&��/��6H��U��I1ڽ!�ٽD6⽼��EV����4�$��8���M���f��4������]u��偬�lת��d��i���K���i�D�P�VD���E�UUU�w�o�?������Τ�ҫ�_﫾|���,N���q���|��a�T�H�U�3��� �U��s����.�߽�ٽ�۽X�潫/��d�	��_��
+��?���U�N�o�}��/U��7��pө���������AJ��U��e�}���_�2K�fDC���I�$]��z�u���͜�eߧ��  �  �ɾ��žo���e��uҒ�O�|�:X�o9����q������޽�Rͽ&ý�D����Ľ�н/d㽀a��}���$��?���_��ۂ��u��绫�`Ǽ�:�Ǿ�ɾS�¾����~ݟ�:����#u��I`�~S\���i��^��節��&��۰���Ǿ�ɾ�~¾{峾۪���勾�p��3M�
0��o���n�Y	ؽhɽ�X�������ǽNֽ�6뽙����%-��I�	�k�����`��	챾00��R?ɾ�EȾ�F��O����R��twl�T�\�j�^��r�j��^���%���85��Oɾ�4Ⱦ�U��(ح�gƙ������c���B�ɕ'����Z �I��Eҽ��Ž�_��|n½��˽�Kܽ���t	��:��6��xT�A�x�M���o,�������ľ��ɾZ�žW>���������1?�{we�#�[��c��{��㏾Mo��.i����ľ�ɾ�ž�m��Ld��<ђ���|��7X��9����n�s���^�޽�Jͽ�ý�<����Ľ7�н�\��Z�������$�1�?�1�_�qۂ��u������Ǽ�݃Ǿ��ɾ��¾����ܟ�����u�UE`��N\���i�&\��q���;$��������Ǿښɾ�|¾�㳾X����䋾cp�2M��0��n�*��?��ؽzɽ1Y�����
�ǽ�ֽ�9뽂��2!��'-��I�M�k�˜��b��1�2���AɾHHȾ[I���Q�������T��}l���\�x�^�Fr�!l��!�������`6��Pɾ`5Ⱦ=V���ح� Ǚ������c��B�~�'����] ���iMҽj�Ž{h��@w½M�˽Tܽ���jx	�N>�6��{T�~�x�����B.������H�ľP�ɾ,�žnA��ص��"��qF��~e�p�[�"�c�ھ{��揾3r���k����ľ�  �  gk�J�޾�+Ͼ!���	̞�hc���Q]�:o7��u����t�㽝w˽�\���F��ï�`���P��н&�H'�mw�j)?���f��݊�ʘ��0����aӾ�ι�B�۾�>ʾ&�������R����|u���p�\l��+X��n���O���վ������ھ�6Ⱦ��+%���z���O��,������Ĉڽ�@Ž����8����U��ox���^ý��׽����|��%)�zK���u��H��@���ž��ؾ�M��⾌�־z�¾Rʪ�¤��偾�q���s�/��lw���<����Ǿ _ھ&�㾷��Xվ����4~��्�	�k��*C���"���	�y��քҽ�㿽c����ٯ�A��������Fɽpi�{ ���9�3���X�α���图�µ���̾Ήݾ�X�%�߾��о]���������{��p��Jy�N܊�7��u^��.�ξ��޾`i侎�޾Q*Ͼ͉���ʞ�5b��vO]��l7��r�������Gp˽KU��?��$��������H��1н�꽮$�Pu��'?���f�E݊���������aӾ��<�x�۾�=ʾ��������D���*xu���p��i���U�����M��
վH�������ھ5Ⱦ����#����z� �O�s�,���������ڽ/@Ž����粰�KW��^z��Kaý��׽�����~�P()��|K�H�u��J��B��C�ž��ؾP㾭��V�־Z�¾?ͪ������灾j�q��s�q1���y���>���ǾC`ھ��\�ᾕXվ�����~��������k��,C�|�"���	�2��?�ҽ뿽����⯽����4���Nɽq཰~ �c����3�ڷX�v���i盾ĵ��̾)�ݾ�[��߾��о���Y���b�7�{�np�,Ry��ߊ����ua����ξ�޾�  �  '�����G�޾0ž3ܧ�>��j�b�p]8�L2�����t�ٽ�&��4c��8è�k������;����ŽOf�S���W�@���m��H���n���5˾�~�<󾯝��c���پ���^s���Z��ԁ���~����%͚�r�����ξt��9���1�����k�־p~���������S��I,�l��ｿSн@�������H��󦽌���@(���~ͽ)���<�Y|(���N��\~�Tњ�y>���Ծ���Þ��������� �Ѿ���PX�����8]�����K\��������m5׾����7�����t��	6ξp���Wo���s��yE��>!�U����㽡5Ƚõ��᪽����+��8�����`Wֽ�d��~��64���]�j
��"���d���+ܾ�	� ���{��\�=�ȾG���핾�/����}�%M����!��Eƾ"�޾f�����@��ĵ޾�
ž�ڧ�����b��Z8�w/�����Ìٽ����[������ec��[��s4��	�Ž~`ཡP�����@���m��H���n���5˾�~���5��������پ?���q���X���с���~�0��ʚ�������ξ������x/����뾤�־�|��g������S�@H,�$���ｄRн� �������I��_���|����*��Ɓͽ��?��~(���N�`~�.Ӛ��@���Ծ&��S�����������Ѿ
���I[������b�<����^��*���T���6׾��뾿8��r	����s6ξ䷱��o��]s��{E�A!�(��U��<Ƚ�ʵ��骽ᇦ��3��U������^ֽ�k����$:4�D�]���蔤�R���7-ܾB�������`��ɾ��w��3��\�}���祓��$��V	ƾ��޾˗��  �  Up��)���鳑�{ၾK6_�!�:��8����}uν�w���Ε�>���8�v��nk�D]h�63m�/]z�˪���[����
?׽���V5 ��|B��g��������f���@��EϚ��쎾�U~�;�]��)B�M41���-��9�'lP���o��6��N2����������N���܌�t�w� �R���.�4?���
K½!���h���ח��N�q��{i�Gi�J�p�)b���č��⡽W~��%t���#+�w�N�|�s�*!��z�������@��.s����5s���S��;�f~.�0�R�?�0Z���z��M��8ę����9�������������k��F���#����l�۽rQ��e����E��|V|�c-n�@sh���j���t�B1��邏�c���?ʽ���W��f�6��[�����#������Y`���l��u������9h��ZJ��k5��g-�k�3�+G�J�d��Ԃ��������Kn��c���[�������3_���:�L6�����oν�q��	ȕ�G�����v��_k�rNh��$m�mOz�r���?V��鳽;׽R��.4 �|B��~g�˲��w������U@��jΚ�c뎾�R~�Û]��%B��/1��-��9�3gP�̆o�#4�� 0��U�������s���bڌ�x�w�a�R�U�.�M=��~꽘H½U���=���K���o�q�B}i��i��p��d���Ǎ�_桽����+y����&+� �N�]�s�F#��R|�����$C���u����k;s�R�S�B#;���.�
"0��?�/4Z� �z�O��jř��������6���J�����k�N�F���#����<�۽W���ǜ��L��`e|��<n�-�h���j�L�t��8��X���%j���Fʽk
�����Ŝ6�#[�����%�����b���o��7x��p���Ah�bJ�&s5�5o-���3���G���d��ׂ����k����  �  �����Ә��d��nV~�R-[� �7��������&ϽH���ŗ�巇���z��}o��bl�Gq�\�~������C���V��f�׽�c�f����?��%c��ׂ��4���H��/d�����5�����x�<Y��q>�h.���*���5��AL��gj��������#��"������f�r�:O��,�:�ON�AUýe[���������	
v�-�m�%m�<�t��y��eЏ���������Jk彿&�\)��AK���n�R���锾K͛��k��rߓ�6ˆ�f�m�OO���7�c+���,��<�|�U��"u�u��=��)��eᚾT���z����g�_lC��"�0=��ܽ���꟞�|W���A���Cr�yl�J�n��y��H��c���+��K˽gt��<��j4�-W�J�z��㌾����c���R���y��^����Pc��`F�2�?U*�X�0��C���_����P���!䘾����6Ҙ�Gc���S~��*[���7��������� Ͻ ��+���߰��E�z��no��Sl�a8q�oz~�2����=���Q��N�׽�a�3��ˊ?�;%c��ׂ�F4��4H���c��������۷x��Y��m>��-��*� �5��<L�cj����æ���뚾�!��J���m�r�g7O�ƴ,�-8�6K��Rý�Y��笑�2���+
v���m��m���t�S|��~ӏ�N������Np彖)��)�EK���n�l��씾�ϛ�[n��⓾�͆���m��TO��7�Vh+���,�q
<���U�&u����p���)��'⚾��������g��mC�1"�=?�g!ܽ����R����^��)I��USr��l�e�n�q y�[P��ԩ��M	��&˽{������4��0W��z��匾F�������)�����������Wc�hF�j 2�\*�i�0�֢C�L�_�����s显�  �  gő������C��N�o�TYP��
1���������Mҽ����UX���}��M����
|���x�H�}�#ㅽ腑�����Rv���ڽ e������7��jW�jv�����7ɏ�4���2ǌ�U����h�	L���3�C�$��"�2�+�zu@���[���x�s���V>��'i��J���!���`e��E��'�[����꽑rǽAZ��d���i��}y����y�yy��R.������f˩��Ľ����;	���#��9B�i�a�O�#
�����P���Ӊ���{� _�3<C�<�-���"���#�=�1��I�{�e�	耾^܋��_��wO��ꈾ?5y�m�Z�YG;�ۚ�i��a޽�����������膽��~�3�x��0{����{��C��׳��Ɏν ��j��;�-���L�]-l�H���򹑾8��Q��"�r��qU�1;���(�i�!�A'��8�$GR��ao� 	���b��hÑ��~��+B����o��VP�%1���#���HҽI����Q��pv���3�{�>�x�*�}��ۅ�7������q��[ڽFc�;����7�-jW��
v�?����ȏ�����Rƌ��S����h��L���3���$�"�p�+��p@��[���x�3���6<��-g��z�� ���]e�W�E��'�}�����(pǽ|X���b��ui���y�� �y��{y��À��0������ϩ�FĽ����>	���#�s=B�>�a�BS�a��' ��ճ���Չ�F�{��%_��AC���-�.�"�z�#�ò1��I���e��逾�݋��`��?P���ꈾ}6y���Z��H;�������|#޽ސ��i���7$����
���x�kA{����V���J��
�����ν�&�������-�"�L�1l��������v������#T����r��xU�;";���(���!��G'���8�XMR�fgo�����d���  �  �,��c�	�p��'[�B���(�í�������ڽ�2��)��� ��L͏�����0��,/��C쑽�G��{d��=�Ž�|������M.�O�G�td`�\�t�-��������c{�1ki���Q�h�8�X$�pL�!��~A�B�.��uF��K_�fet�ȹ������a�{�3j�N�R�h�9��� ��
����F;ѽ9����B��Җ�R���函�����8������i��)-���2ν�%��e��(���6��2P���g��z������ ���Iv�l�a��9I��J1����?�tx��:"�hL6���N���f�F�y�����&���v���b��J�?1�u�g���佒bȽF����韽�	��LȊ��?��V����ˎ�i�����p���5|׽}����I�+&��4?��uX���n�L~��*��e�}Ap��Y�c�@��P*�D{��l��I�,'(��3>�+W�@n�U.~��*���{��p�E%[��B�D�(�)��W�����ڽ#,��"�����vŏ�����(��9'���䑽�@��^����Ž;x�0��p���L.�h�G��c`���t��������b{��hi�)�Q��8��$�DH�����<���.��pF�G_�at���������ؐ{��/j�q�R��9��� ��
�����8ѽ|����A���і�g��x懽ʠ���:��f����l���0���6ν�*콜h��+��6��6P���g�Hz�Á� #���Nv���a�?I��O1����-D�B}�?"�bP6�	�N���f���y������&��s�v���b�X�J��1�i��
�7���hȽE���|񟽫���Њ�uH��ۥ��Ԏ�y����#������"�׽!����L�n&��7?�UyX���n�uP~�	-��wj�PGp�C�Y���@��W*�'��rs�FP��-(��9>��0W�<n��2~��  �  ;a�c�^�[U��.F���4���"��B�X��7�G�Խ�)�����,ۡ�?����`������^��uu��,xĽd�ٽ���V�������&���8�d�I���W�-`��`�o�X���I��t6�^J"�ta�G��/����A(��V-�g�A���R�0^��Wa�EU\��P�.�@���.��+���F�����ͽ@��������B��J뗽+���N���X	��W/˽@e������e�zJ��,���>���N�N[�&(a���^���T��C�u�/�m��
�wL��J����_+ ��)4��G���W��*`�v�`�fY�ؑK�k�:�*�(���'����08ܽ��ƽ6@�����l͛��t���$������U@��I��DҽCp�"��6���� �ެ2��ND��S��^��[a��W\���O��4=�M�(�j���	�š�������R�&��:�8�M��G[�B7a��^�kU�1,F�j�4�q�"�Y@�GU�b1콂�Խ�"��9��ҡ�����(X��g���V���m��6qĽ=�ٽs��*�������&���8�i�I���W�`�v�`���X�h�I��q6�G"��]�@���������#�fR-��A���R�,^� Ta��Q\�֑P�g~@�B�.��)�,�W|��b�U�ͽ( ��$��&����B���엽�������d���2˽�iὢ���xh��M�z�,�D�>���N�`R[��,a���^���T��C���/�����hQ�OO�+��D/ �c-4�n�G�1�W��,`�8�`��Y�a�K��:��(�-����	����>ܽq�ƽQH������J֛��}���-��7����H��0���KҽAw�r��i��� �#�2��QD�ʪS�^�,`a��\\���O��:=���(��p�D�	�P�����߭��&�[�:��M��K[��  �  ��?��@�Ҵ<�ru5��y,���"��E��l�W�}����߽�˽̺��g���[����������@Ͻ��㽛����u�`��m�%�q�.�tE7�g�=�<�@�h�>��7���*�G���&�7�����뽢���@����M����#�2�U<�Ҙ@��?�/�:��2�+P)�e�����
����%j�gؽ�Ž/���ƀ������R���3ýI�ս���9] ���
����q���=(��1�e�9��_?���@��<�RX3�4�%����N��,��E(�[������}	��-���(���5�U'>�3�@�Jt>��"8���/��&��}���L��M���l,��aѽ=�������w������H����Ƚ�ܽ{?�q���J�,.��!��j+�5�4�<��`@�@��6:��%/��U ��B��������s=�3� �������-�:9�%�?�Ҙ@���<��r5�rw,�%�"��B��i��h����	߽|˽Aú��^��XR��w���ｽ88ϽI��҄���r���k�u%��.�@D7�9�=���@�ݻ>��7�o�*�����#������n��T8�q������#���1���;�@�@���?�2�:�V�2��M)�X����a	�r��h�Xؽ`ŽK���v�������T��6ýO�ս* �T_ ���
�D��v���@(���1�O�9��c?��@���<�,]3�0�%����(S�v6���1�f��L���_�	�1���(��5�y)>��@�v>��$8�W�/��!&�U������������}4潧jѽd���\��7���j����Q��ɽ9�ܽG����GN�S1�'�!�n+���4��	<��d@�r@��;:�+/�a[ ��H�"�����),轐I�� �������-�>9��  �  ^�#�k�(�}�+�t�,���,�ns+���(���#�Du���~H�����ڽ��̽�Ƚ(Ͻ��޽����,�BL������$��~)�%�+�6�,�t,�Y +�(�5a"�S��3��'�j���׽�i˽)ɽ�ѽg�2��9	��)�p����%�*��,��,��Q,�ܿ*��D'�/'!�("���� ��罧�Խ�Jʽ(�ɽSӽ���c<���L�q��I ���&�5v*�	4,���,��$,��O*�Ho&���U[�D�
�f����P�~�ҽ�sɽ�ʽC�ս�.� � ��[���T�!�B�'���*�d],�2�,�A�+��)�!�%��u�@�����e�������Yн��ȽS�˽ˌؽ�����k`�	_�5�"�F>(��:+��z,��,��+�*K)�&�$�U�����9d����-�ݽ0lν^�ȽvIͽ\۽����`Z������#�Z�(���+�ߑ,��,��p+�Ư(���#��q�b��jD�͗ｮ~ڽ��̽*�Ƚ\
Ͻu�޽������H��}���$�K|)�6�+���,��r,��+��(��_"�_����P$�E���׽�b˽Sɽ�ѽ.����5	��%����;�%���)�,�R�,�xO,��*�C'��%!�!�A��D ������Խ�Kʽm�ɽ�Tӽ��b?��aN����lK �;�&�,y*�K7,�E�,��(,��S*��s&����`��
�"����Z�	�ҽ�|ɽϥʽe�սU6�P� ��^������!�D�'���*�N_,�B�,���+���)�9�%�;y�8��܆�����h���cн��Ƚ<�˽Z�ؽ��L��Pd��b���"�^A(��=+��},�5�,�C�+��N)�<�$������}i��󽱟ݽ�wν�Ƚ�TͽT�۽X��T���^�����  �  \������u#���,���5��=���@�]{?� �8�8�,�?�����������6<��𽬛��(�	=!�B�/���:��9@��B@���;��
4���*��Q!�?��ͽ��Y�5��۽YȽ����PZ��Z���g�������Հҽ<e�*'���0	��J�2�v�&�0�Ǐ8�ϴ>�P�@���=��F5��(��H����f��VD�=��9���k{�^g&��4��%=�~�@��)?��`9�31�J�'����^�R
�Є��$��M�ԽGE½+����ݭ�����5��ƽ�:ٽ��*(�=��2��> ��)��3���:��?�8{@���;�XO1���"����
��K�s�hI�C!��������Q+�ٟ7�f�>���@���=�Q�6��.���$�e��T����M�����o%ν��������G��F°�i���G̽�6��������������r#��,�$�5�=�0�@�Ax?���8�R�,���]��ͱ��_��1�~�𽋖�$��8!�'�/��:��6@�L@@�h�;�	4�C�*�P!����	���W��
񽚉۽_�ǽd���6S��ܓ�������}��yҽ�]����9-	��G�+���&��0���8��>���@�m�=��E5�!(�H�����f��
E꽁���;��A��|�"i&��4�'(=��@��,?�d9��1��'���c�xV
����q�齳�Խ�N½`����歽yƮ��=��Hƽ,Aٽ٣*����S��@ �5�)��3�f�:� �?��~@�l�;��S1�<�"���G�eV�2~��S�M+�����=���U+�y�7��?���@�}�=�.�6��	.�ч$����$�K���V������/νu'�������R��
Ͱ���̽�?��������  �  � ��$���#�_�5��G���U�`1_��a�J�Z�c�L���9��%�h��l'�����
�UX�`�)�hV>��uP�O�\�ha��]���R�`C���1�� ���V����ѽ!
���u��d ��_똽����^=��Bg���3����ǽ��ݽU"�����L��޺)��;��nL���Y�Ѻ`���_���V��F�3��#���+����������0���D�7YU��H_�_
a���Z�N�%�=���+��\�(�
�)��e�8ʽ,���̧�'��^×��p�����֪������ν�a����j����&�/�EvA�!^Q���\�aa���]��'R���@�1,�n/�:0����Q�b(�-X#�#�7���J�ҁY���`���_�(W�1�H���7�!�%�������c�jؽ:Xý|�����������O��� ���l��yǯ�Y1����ս�����!��#��5�G��U��._�Sa���Z�Q�L�%�9�%�%�'���!�"��
��R�"�)��Q>�qP�\�\��da�-�]�i�R��]C��1�6 ����x���Mѽ����o�����䘽�����5���_��I,��T�ǽ�}ݽ������c��5�)���;��lL���Y�;�`�}�_���V�J�F��3��#�������������6�0�c�D�?[U��J_��a���Z�2!N���=���+�v`�=�
����6�;ʽE���է����˗�y��0���ݪ�\��ӵν=g���������o�/��xA��`Q��\��da���]�,R���@�l6,��4��5�N���V��-�]#���7���J�}�Y���`���_��*W���H���7��%�W��/��tk�:sؽ}aýI���ĸ��v����Y���
���v���Я��9����ս����  �  ����x���,*��}C��{\���q�����%��؊}���l�)�U���<�!'�)��^���&�mt+��PB��I[�,Xq�l��O&����}�?�m��W���=�[�$���������սR��F%���阽�Z���o��X���$��h���}ɠ�����ɽ����R�"z2�G L�l.d��w�~S��柁�b�x�1�e��oM�W5��V!���2����W�2�9�J��0c��6w��O������	9y�P�f�(�N��E5�|��	I��N꽞�̽L��������ٔ��Ӌ��~��%��}p��}���1���͹�G�ҽ�����j"���:�~^T�cXk�%L|�
��>}��Lcs���]��E�H�-����� ���%�i2:��S��j� |�s	��(���2�s��_�dTF���,��P��� ���߽S2Ľ�G���o�� V���ډ��!��P���F���ܛ�	*���~���bܽx������Z**�d{C�y\��q�'��"$���}���l�s�U���<��'�d��tz�� ��n+�&KB�QD[�kSq�.��u$����}���m�ZW���=�s�$������F�սdM�� ��?䘽�T��i��Q�����/���M �t���4�ɽ�����O��w2���K�Y,d��w��R��C���`�x�t�e�CoM�&5��V!�B �ԃ�����2���J��2c��8w��P������;y�d�f�|�N�EI5�F��M��V�7�̽������b┽�܋�&���&��x������7��kӹ���ҽ�������"�9�:�(aT�b[k��O|���q��,hs�$�]�kE� �-���Ӵ����N%��7:��S�=�j��#|���������s�m_�	WF�^�,� T��� �j�߽r:ĽXP��y���_���䉽c+���Y���O��_国62��"���Niܽ�  �  �U����x�2�-R��-q��腾'ڎ�����t���b��6�m���P��c7�X�&���!��l)�Bn<�|W��.t���nh�������W��A��ـj�/K�~	,��3����P�̽�Y��WI���b��,�����z���x���`y��k���s(���$���2�n@�Y)��=�G�\�w�z��x��"����<��a���.��Cd���G��0��#��"�w�.���D��`�ug}�s\��Y吾J�s�����}��+`�|z@��K"�����d� \½����o���ϓ���h���?y��2z��ց�G
���R������d.ɽ7�^�Y�(���G��g��؁��x��d���B����#��'Kw�+CZ��?�i+���!�q%�l5�w�M�܉j�L���3��`���B}��w&���mt��U�h6���H  �ؽs븽苡�'����Y��Z}���x��g|�sc�� 1��\_��!����.Խ�O���� �2��R�U+q�3煾�؎�4������i`��Z�m�<�P��]7�Z�&�y�!�jf)�2h<��W�:)t�}���2f�������U���?��^~j��K�z,��1�����̽'U��.D���\�������z�i�x�;��[r��o𓽚!�����f,�y=��&� =��\�p�z��w��`����;���`��p.���d���G��0�J�#���"�_�.�"�D�t�`�/i}�r]��z搾��؉����}�*/`� ~@�mO"�����l�od½�������p���!q��OPy�rBz�Sށ�+��DY�������3ɽ<�a���(�!�G��g�Xځ�cz��o������� &���Pw�IZ��?��+���!��v%�5���M���j�l���5������~���'��pt���U�!6���|# �ؽ6�I������c��m}���x�yz|�ll���9��>g��W���5Խ�  �  "x���}���9��+]�j�����X9��菜��|���፾>~��"^�
KB���/� m*�B�2���G�e�z����������fv������Z ����x��1U�#@2�����2ɽh���e���\����Ox�Hgn�f�l���r�π�"3���ݟ��\��?f޽)��{�#��_E��i�����$��^%����z����A���Xs�9T�3�:���,�Ϲ+��8���P���o�b����v��o���]���CW��>9���m�'II��I'���	����Խ�1\��{玽�⁽�t�`�l��m�u�v��M��`��������6Žk��3����.�
5Q�d�t���������C������"���C���h�\�J�{�4��*�{�.��?�B�Z�C�z�\a��o���Rw���򙾫����g&a�Л=������ �cwս���	���퉽:~}���p��Gl���o�(�{��j��'՘�Ո���4ѽbr��]{�#�9��)]�4��r���7��7����z���ߍ�I~�i^�3EB�u�/��f*���2���G�e�����ﱐ�@��at��󁗾���#�x��/U�>2�������ɽ����B���Ǜ���Cx��Zn��l�&�r�Ȁ�F,��2ן�[V��`޽@��ǿ#�d]E�pi����0#���$��b������*A��jXs�T�J�:��,�q�+��8��P�+�o�=����w�����������X���:���m��LI�;M'�c�	���9ݽ��d��	���*끽�t���l���m��v�ZT����������:<Ž��콪��m�.��7Q�E�t����������E��򥚾����F���h���J�Ƕ4�W�*���.�ò?���Z��z��c��Q����x��������
����(a�f�=�`���� �B~ս����.������C�}��p�=Zl�"�o���{��r���ܘ�⏰�:;ѽ�  �  Q�������<� Ia�ق�u��{����m���7��3B���큾��b�#F��#3�a�-��L6���K��j������,�� ̝��R���-���X���}�K�X�S�4�h(��Y�:Ƚz쨽��������,t�s[j��h��n�Rp}��"��Q��d��]2޽�n�O�%�%�H���m�w�������󞾴ܟ��7���z����x�\�X�+|>�:�/���.��5<��4U�
u�̊�b��{���n���ᗾ�@��`�q�&�L��F)�X}
�������r���ڌ�x��v�o�/�h��i�e�r��5������7��W:Ľ^�����0��T���y�����(������q��釕�8S���m�C�N�w8�v�-� �1��oC�#W_����(���-K���T������꓾�����ke��y@��m���<�ԽQ>��(��Tه�=Ty�6�l��Bh��k�hzw��T���ᖽI��^�н`K����R~<��Fa��ׂ��s���l��6���?��T끾z�b�:F��3�z-�eF6�T�K��
j�����f*���ɝ��P��,��@W��y�}���X�6�4�^&��U�.6Ƚ�稽����&���� t��Nj��h��n��b}�����������5,޽�k���%���H�c�m�v������#�ܟ�d7���z����x�.�X�B|>���/���.��6<��5U�|u��̊�`��0|���o��0㗾B����q���L�~J)�6�
���c���畠��⌽l���o�X�h���i��r�u<��M���
���?Ľx����c�0���T���y�H����)������s������V���m���N��8���-�8�1�kuC�}\_�i��O���M��LV��h���\듾1�ine�2|@�`p��� ս�E��00���ᇽfy�z�l��Th�
�k�ŋw��\��/閽H
����н�  �  "x���}���9��+]�j�����X9��菜��|���፾>~��"^�
KB���/� m*�B�2���G�e�z����������fv������Z ����x��1U�#@2�����2ɽh���e���\����Ox�Hgn�f�l���r�π�"3���ݟ��\��?f޽)��{�#��_E��i�����$��^%����z����A���Xs�9T�3�:���,�Ϲ+��8���P���o�b����v��o���]���CW��>9���m�'II��I'���	����Խ�1\��{玽�⁽�t�`�l��m�u�v��M��`��������6Žk��3����.�
5Q�d�t���������C������"���C���h�\�J�{�4��*�{�.��?�B�Z�C�z�\a��o���Rw���򙾫����g&a�Л=������ �cwս���	���퉽:~}���p��Gl���o�(�{��j��'՘�Ո���4ѽbr��]{�#�9��)]�4��r���7��7����z���ߍ�I~�i^�3EB�u�/��f*���2���G�e�����ﱐ�@��at��󁗾���#�x��/U�>2�������ɽ����B���Ǜ���Cx��Zn��l�&�r�Ȁ�F,��2ן�[V��`޽@��ǿ#�d]E�pi����0#���$��b������*A��jXs�T�J�:��,�q�+��8��P�+�o�=����w�����������X���:���m��LI�;M'�c�	���9ݽ��d��	���*끽�t���l���m��v�ZT����������:<Ž��콪��m�.��7Q�E�t����������E��򥚾����F���h���J�Ƕ4�W�*���.�ò?���Z��z��c��Q����x��������
����(a�f�=�`���� �B~ս����.������C�}��p�=Zl�"�o���{��r���ܘ�⏰�:;ѽ�  �  �U����x�2�-R��-q��腾'ڎ�����t���b��6�m���P��c7�X�&���!��l)�Bn<�|W��.t���nh�������W��A��ـj�/K�~	,��3����P�̽�Y��WI���b��,�����z���x���`y��k���s(���$���2�n@�Y)��=�G�\�w�z��x��"����<��a���.��Cd���G��0��#��"�w�.���D��`�ug}�s\��Y吾J�s�����}��+`�|z@��K"�����d� \½����o���ϓ���h���?y��2z��ց�G
���R������d.ɽ7�^�Y�(���G��g��؁��x��d���B����#��'Kw�+CZ��?�i+���!�q%�l5�w�M�܉j�L���3��`���B}��w&���mt��U�h6���H  �ؽs븽苡�'����Y��Z}���x��g|�sc�� 1��\_��!����.Խ�O���� �2��R�U+q�3煾�؎�4������i`��Z�m�<�P��]7�Z�&�y�!�jf)�2h<��W�:)t�}���2f�������U���?��^~j��K�z,��1�����̽'U��.D���\�������z�i�x�;��[r��o𓽚!�����f,�y=��&� =��\�p�z��w��`����;���`��p.���d���G��0�J�#���"�_�.�"�D�t�`�/i}�r]��z搾��؉����}�*/`� ~@�mO"�����l�od½�������p���!q��OPy�rBz�Sށ�+��DY�������3ɽ<�a���(�!�G��g�Xځ�cz��o������� &���Pw�IZ��?��+���!��v%�5���M���j�l���5������~���'��pt���U�!6���|# �ؽ6�I������c��m}���x�yz|�ll���9��>g��W���5Խ�  �  ����x���,*��}C��{\���q�����%��؊}���l�)�U���<�!'�)��^���&�mt+��PB��I[�,Xq�l��O&����}�?�m��W���=�[�$���������սR��F%���阽�Z���o��X���$��h���}ɠ�����ɽ����R�"z2�G L�l.d��w�~S��柁�b�x�1�e��oM�W5��V!���2����W�2�9�J��0c��6w��O������	9y�P�f�(�N��E5�|��	I��N꽞�̽L��������ٔ��Ӌ��~��%��}p��}���1���͹�G�ҽ�����j"���:�~^T�cXk�%L|�
��>}��Lcs���]��E�H�-����� ���%�i2:��S��j� |�s	��(���2�s��_�dTF���,��P��� ���߽S2Ľ�G���o�� V���ډ��!��P���F���ܛ�	*���~���bܽx������Z**�d{C�y\��q�'��"$���}���l�s�U���<��'�d��tz�� ��n+�&KB�QD[�kSq�.��u$����}���m�ZW���=�s�$������F�սdM�� ��?䘽�T��i��Q�����/���M �t���4�ɽ�����O��w2���K�Y,d��w��R��C���`�x�t�e�CoM�&5��V!�B �ԃ�����2���J��2c��8w��P������;y�d�f�|�N�EI5�F��M��V�7�̽������b┽�܋�&���&��x������7��kӹ���ҽ�������"�9�:�(aT�b[k��O|���q��,hs�$�]�kE� �-���Ӵ����N%��7:��S�=�j��#|���������s�m_�	WF�^�,� T��� �j�߽r:ĽXP��y���_���䉽c+���Y���O��_国62��"���Niܽ�  �  � ��$���#�_�5��G���U�`1_��a�J�Z�c�L���9��%�h��l'�����
�UX�`�)�hV>��uP�O�\�ha��]���R�`C���1�� ���V����ѽ!
���u��d ��_똽����^=��Bg���3����ǽ��ݽU"�����L��޺)��;��nL���Y�Ѻ`���_���V��F�3��#���+����������0���D�7YU��H_�_
a���Z�N�%�=���+��\�(�
�)��e�8ʽ,���̧�'��^×��p�����֪������ν�a����j����&�/�EvA�!^Q���\�aa���]��'R���@�1,�n/�:0����Q�b(�-X#�#�7���J�ҁY���`���_�(W�1�H���7�!�%�������c�jؽ:Xý|�����������O��� ���l��yǯ�Y1����ս�����!��#��5�G��U��._�Sa���Z�Q�L�%�9�%�%�'���!�"��
��R�"�)��Q>�qP�\�\��da�-�]�i�R��]C��1�6 ����x���Mѽ����o�����䘽�����5���_��I,��T�ǽ�}ݽ������c��5�)���;��lL���Y�;�`�}�_���V�J�F��3��#�������������6�0�c�D�?[U��J_��a���Z�2!N���=���+�v`�=�
����6�;ʽE���է����˗�y��0���ݪ�\��ӵν=g���������o�/��xA��`Q��\��da���]�,R���@�l6,��4��5�N���V��-�]#���7���J�}�Y���`���_��*W���H���7��%�W��/��tk�:sؽ}aýI���ĸ��v����Y���
���v���Я��9����ս����  �  \������u#���,���5��=���@�]{?� �8�8�,�?�����������6<��𽬛��(�	=!�B�/���:��9@��B@���;��
4���*��Q!�?��ͽ��Y�5��۽YȽ����PZ��Z���g�������Հҽ<e�*'���0	��J�2�v�&�0�Ǐ8�ϴ>�P�@���=��F5��(��H����f��VD�=��9���k{�^g&��4��%=�~�@��)?��`9�31�J�'����^�R
�Є��$��M�ԽGE½+����ݭ�����5��ƽ�:ٽ��*(�=��2��> ��)��3���:��?�8{@���;�XO1���"����
��K�s�hI�C!��������Q+�ٟ7�f�>���@���=�Q�6��.���$�e��T����M�����o%ν��������G��F°�i���G̽�6��������������r#��,�$�5�=�0�@�Ax?���8�R�,���]��ͱ��_��1�~�𽋖�$��8!�'�/��:��6@�L@@�h�;�	4�C�*�P!����	���W��
񽚉۽_�ǽd���6S��ܓ�������}��yҽ�]����9-	��G�+���&��0���8��>���@�m�=��E5�!(�H�����f��
E꽁���;��A��|�"i&��4�'(=��@��,?�d9��1��'���c�xV
����q�齳�Խ�N½`����歽yƮ��=��Hƽ,Aٽ٣*����S��@ �5�)��3�f�:� �?��~@�l�;��S1�<�"���G�eV�2~��S�M+�����=���U+�y�7��?���@�}�=�.�6��	.�ч$����$�K���V������/νu'�������R��
Ͱ���̽�?��������  �  ^�#�k�(�}�+�t�,���,�ns+���(���#�Du���~H�����ڽ��̽�Ƚ(Ͻ��޽����,�BL������$��~)�%�+�6�,�t,�Y +�(�5a"�S��3��'�j���׽�i˽)ɽ�ѽg�2��9	��)�p����%�*��,��,��Q,�ܿ*��D'�/'!�("���� ��罧�Խ�Jʽ(�ɽSӽ���c<���L�q��I ���&�5v*�	4,���,��$,��O*�Ho&���U[�D�
�f����P�~�ҽ�sɽ�ʽC�ս�.� � ��[���T�!�B�'���*�d],�2�,�A�+��)�!�%��u�@�����e�������Yн��ȽS�˽ˌؽ�����k`�	_�5�"�F>(��:+��z,��,��+�*K)�&�$�U�����9d����-�ݽ0lν^�ȽvIͽ\۽����`Z������#�Z�(���+�ߑ,��,��p+�Ư(���#��q�b��jD�͗ｮ~ڽ��̽*�Ƚ\
Ͻu�޽������H��}���$�K|)�6�+���,��r,��+��(��_"�_����P$�E���׽�b˽Sɽ�ѽ.����5	��%����;�%���)�,�R�,�xO,��*�C'��%!�!�A��D ������Խ�Kʽm�ɽ�Tӽ��b?��aN����lK �;�&�,y*�K7,�E�,��(,��S*��s&����`��
�"����Z�	�ҽ�|ɽϥʽe�սU6�P� ��^������!�D�'���*�N_,�B�,���+���)�9�%�;y�8��܆�����h���cн��Ƚ<�˽Z�ؽ��L��Pd��b���"�^A(��=+��},�5�,�C�+��N)�<�$������}i��󽱟ݽ�wν�Ƚ�TͽT�۽X��T���^�����  �  ��?��@�Ҵ<�ru5��y,���"��E��l�W�}����߽�˽̺��g���[����������@Ͻ��㽛����u�`��m�%�q�.�tE7�g�=�<�@�h�>��7���*�G���&�7�����뽢���@����M����#�2�U<�Ҙ@��?�/�:��2�+P)�e�����
����%j�gؽ�Ž/���ƀ������R���3ýI�ս���9] ���
����q���=(��1�e�9��_?���@��<�RX3�4�%����N��,��E(�[������}	��-���(���5�U'>�3�@�Jt>��"8���/��&��}���L��M���l,��aѽ=�������w������H����Ƚ�ܽ{?�q���J�,.��!��j+�5�4�<��`@�@��6:��%/��U ��B��������s=�3� �������-�:9�%�?�Ҙ@���<��r5�rw,�%�"��B��i��h����	߽|˽Aú��^��XR��w���ｽ88ϽI��҄���r���k�u%��.�@D7�9�=���@�ݻ>��7�o�*�����#������n��T8�q������#���1���;�@�@���?�2�:�V�2��M)�X����a	�r��h�Xؽ`ŽK���v�������T��6ýO�ս* �T_ ���
�D��v���@(���1�O�9��c?��@���<�,]3�0�%����(S�v6���1�f��L���_�	�1���(��5�y)>��@�v>��$8�W�/��!&�U������������}4潧jѽd���\��7���j����Q��ɽ9�ܽG����GN�S1�'�!�n+���4��	<��d@�r@��;:�+/�a[ ��H�"�����),轐I�� �������-�>9��  �  ;a�c�^�[U��.F���4���"��B�X��7�G�Խ�)�����,ۡ�?����`������^��uu��,xĽd�ٽ���V�������&���8�d�I���W�-`��`�o�X���I��t6�^J"�ta�G��/����A(��V-�g�A���R�0^��Wa�EU\��P�.�@���.��+���F�����ͽ@��������B��J뗽+���N���X	��W/˽@e������e�zJ��,���>���N�N[�&(a���^���T��C�u�/�m��
�wL��J����_+ ��)4��G���W��*`�v�`�fY�ؑK�k�:�*�(���'����08ܽ��ƽ6@�����l͛��t���$������U@��I��DҽCp�"��6���� �ެ2��ND��S��^��[a��W\���O��4=�M�(�j���	�š�������R�&��:�8�M��G[�B7a��^�kU�1,F�j�4�q�"�Y@�GU�b1콂�Խ�"��9��ҡ�����(X��g���V���m��6qĽ=�ٽs��*�������&���8�i�I���W�`�v�`���X�h�I��q6�G"��]�@���������#�fR-��A���R�,^� Ta��Q\�֑P�g~@�B�.��)�,�W|��b�U�ͽ( ��$��&����B���엽�������d���2˽�iὢ���xh��M�z�,�D�>���N�`R[��,a���^���T��C���/�����hQ�OO�+��D/ �c-4�n�G�1�W��,`�8�`��Y�a�K��:��(�-����	����>ܽq�ƽQH������J֛��}���-��7����H��0���KҽAw�r��i��� �#�2��QD�ʪS�^�,`a��\\���O��:=���(��p�D�	�P�����߭��&�[�:��M��K[��  �  �,��c�	�p��'[�B���(�í�������ڽ�2��)��� ��L͏�����0��,/��C쑽�G��{d��=�Ž�|������M.�O�G�td`�\�t�-��������c{�1ki���Q�h�8�X$�pL�!��~A�B�.��uF��K_�fet�ȹ������a�{�3j�N�R�h�9��� ��
����F;ѽ9����B��Җ�R���函�����8������i��)-���2ν�%��e��(���6��2P���g��z������ ���Iv�l�a��9I��J1����?�tx��:"�hL6���N���f�F�y�����&���v���b��J�?1�u�g���佒bȽF����韽�	��LȊ��?��V����ˎ�i�����p���5|׽}����I�+&��4?��uX���n�L~��*��e�}Ap��Y�c�@��P*�D{��l��I�,'(��3>�+W�@n�U.~��*���{��p�E%[��B�D�(�)��W�����ڽ#,��"�����vŏ�����(��9'���䑽�@��^����Ž;x�0��p���L.�h�G��c`���t��������b{��hi�)�Q��8��$�DH�����<���.��pF�G_�at���������ؐ{��/j�q�R��9��� ��
�����8ѽ|����A���і�g��x懽ʠ���:��f����l���0���6ν�*콜h��+��6��6P���g�Hz�Á� #���Nv���a�?I��O1����-D�B}�?"�bP6�	�N���f���y������&��s�v���b�X�J��1�i��
�7���hȽE���|񟽫���Њ�uH��ۥ��Ԏ�y����#������"�׽!����L�n&��7?�UyX���n�uP~�	-��wj�PGp�C�Y���@��W*�'��rs�FP��-(��9>��0W�<n��2~��  �  gő������C��N�o�TYP��
1���������Mҽ����UX���}��M����
|���x�H�}�#ㅽ腑�����Rv���ڽ e������7��jW�jv�����7ɏ�4���2ǌ�U����h�	L���3�C�$��"�2�+�zu@���[���x�s���V>��'i��J���!���`e��E��'�[����꽑rǽAZ��d���i��}y����y�yy��R.������f˩��Ľ����;	���#��9B�i�a�O�#
�����P���Ӊ���{� _�3<C�<�-���"���#�=�1��I�{�e�	耾^܋��_��wO��ꈾ?5y�m�Z�YG;�ۚ�i��a޽�����������膽��~�3�x��0{����{��C��׳��Ɏν ��j��;�-���L�]-l�H���򹑾8��Q��"�r��qU�1;���(�i�!�A'��8�$GR��ao� 	���b��hÑ��~��+B����o��VP�%1���#���HҽI����Q��pv���3�{�>�x�*�}��ۅ�7������q��[ڽFc�;����7�-jW��
v�?����ȏ�����Rƌ��S����h��L���3���$�"�p�+��p@��[���x�3���6<��-g��z�� ���]e�W�E��'�}�����(pǽ|X���b��ui���y�� �y��{y��À��0������ϩ�FĽ����>	���#�s=B�>�a�BS�a��' ��ճ���Չ�F�{��%_��AC���-�.�"�z�#�ò1��I���e��逾�݋��`��?P���ꈾ}6y���Z��H;�������|#޽ސ��i���7$����
���x�kA{����V���J��
�����ν�&�������-�"�L�1l��������v������#T����r��xU�;";���(���!��G'���8�XMR�fgo�����d���  �  �����Ә��d��nV~�R-[� �7��������&ϽH���ŗ�巇���z��}o��bl�Gq�\�~������C���V��f�׽�c�f����?��%c��ׂ��4���H��/d�����5�����x�<Y��q>�h.���*���5��AL��gj��������#��"������f�r�:O��,�:�ON�AUýe[���������	
v�-�m�%m�<�t��y��eЏ���������Jk彿&�\)��AK���n�R���锾K͛��k��rߓ�6ˆ�f�m�OO���7�c+���,��<�|�U��"u�u��=��)��eᚾT���z����g�_lC��"�0=��ܽ���꟞�|W���A���Cr�yl�J�n��y��H��c���+��K˽gt��<��j4�-W�J�z��㌾����c���R���y��^����Pc��`F�2�?U*�X�0��C���_����P���!䘾����6Ҙ�Gc���S~��*[���7��������� Ͻ ��+���߰��E�z��no��Sl�a8q�oz~�2����=���Q��N�׽�a�3��ˊ?�;%c��ׂ�F4��4H���c��������۷x��Y��m>��-��*� �5��<L�cj����æ���뚾�!��J���m�r�g7O�ƴ,�-8�6K��Rý�Y��笑�2���+
v���m��m���t�S|��~ӏ�N������Np彖)��)�EK���n�l��씾�ϛ�[n��⓾�͆���m��TO��7�Vh+���,�q
<���U�&u����p���)��'⚾��������g��mC�1"�=?�g!ܽ����R����^��)I��USr��l�e�n�q y�[P��ԩ��M	��&˽{������4��0W��z��匾F�������)�����������Wc�hF�j 2�\*�i�0�֢C�L�_�����s显�  �  �fG�4�B��6��-#�S6������Ľ�+��셆�OWc��rE��(1�fS$�T�ei�nn���&���4�*/K��k���I���ͽٌ���6���'��v9���D��0G���@���2��= �Q��k����X�=|�g������o���*��r;��oE���F�O]?�DB0�x����y�߽���&����}��"X��=��,�d[!�2������ ��*��R;��T���x�H������U�ڽ~-�f��h2.��>��pF�]F���<�-����]���.�<ὸ�'���j�
���n�0�ʟ?�D�F��PE�;���)���Lu���ѽ�������o��0N�*�6�
�'���q�����8#�X/�h�B�l_��ۃ����������,�
�� ��%4�3�A��QG�>�C�:8�V�&�C��4��_���߽/|�~���2����$���6��B��bG���B���5��*#��3�q���Ľ&�� ����Jc�meE�1�.E$��E��Z�S`�3�&��4��#K�{k��
���E��R�ͽ�����5�ٻ'��u9���D�/G��@���2��: ��������P但s�^��@��2k���*�Jn;��kE���F��Y?�!?0��
����:�߽釸�#��
�}�9X���=��,��[!�����+� �՝*��X;�.�T��x��������e�ڽ�0���c6.�>�NuF�)
F���<�6-�3������8�6"�+����^�
�
�l�0�N�?�\�F��RE��;�g�)�����x����ѽ!������o��=N���6���'�P�1��O��yH#�<g/��B�?z_�y⃽H��������
齲�
��� �*4���A��VG���C��?8���&����;�*m�e�߽t��8��1��K�$���6���B��  �  ��B�!v>�r2������
�@��T7ý춡������Pe���G�T�3���&����:��H� ��@)�ɖ7���M��Mm��S��ؕ����˽������\$��s5��,@�]�B�<�+�.�"����	����$Uཙ�ܽ�y齚H��R�F'�{A7��@�-\B�0$;�̓,�������ܽoN��x����~�;WZ��E@�%�.�"�#�����Y�r#�_<-�M�=���V��Mz�;����z���xؽ#����̖*� �9���A�]�A�o�8�u>)��n���n���,ݽ�߽�������b-�O;��cB���@�X�6��}&�8�����Z�Ͻ�!��[��+xq���P��9��w*�f�!����KZ�h�%���1�|<E��za�_���a��-&����!`�*���S0��o=���B��t?�}!4��*#�_�e����5��۽�`�1������!�x2��>���B��r>�K2����
���2ýj����GDe���G��3�|�&�^�����	� �3)�"�7���M��Cm�uO��T���Ƀ˽������[$��r5��+@��B�.}<���.�L����	����L��ܽ�p�D��M��A'�==7��@�oXB�� ;���,�*����w�ܽ�J�������~��SZ�_C@�$�.�L�#�K��\�#�*A-�E�=��V�&Vz����f����~ؽt&�=��Ě*�D�9��A�%�A�k�8��C)�*t�������6ݽ4߽�"���;��`-��Q;��eB���@�� 7�&���G����Ͻ�%��e"����q�q�P�ܟ9�K�*���!�A�j���%�2�4KE��a��e��sh���,��K
潤c����W0�ft=���B��y?�I'4��0#���Ə��NC彊�۽�m㽻=����/!�
}2���>��  �  �(6��O2�dV'��,��V�&t�5L��mC��s���.Ul�kHP��U<��$/�!�'���%���(�6�1��$@��U���s��㍽Kr����ƽ���
��V��M*�y�3���5��=0���#�#Q�v�~��=�Խ�vѽ5Aݽ���V�����lq+��W4�(�5�Q]/��f"�������T?ֽ����S������J�a�l�H��47�i,��j&�S&� +���5��rF�t�^�	��Ż���7���Aҽ�x��\��P� ��2.��b5�	�4�6�,����p��[���d߽4 ҽ3�ӽ�9佲0 ��Z��("�-'/��5�!q4�֭+�F����
���R�ʽ���+m��d�w��X�XB���2���)��%�0/'���-��:��M���h�F����A��>���R޽M-�z'���%��f1�U6���2�h�(�������｡Yٽ��н��׽6������+�V'�`#2�%6�'L2�ES'��)��S��n��F���=�������Hl��:P�qG<�/�(�'���%���(�.1��@� �U�U�s�ߍ��n��~�ƽ$����b��L*�I�3�P�5�<0�m�#�RN�0�!��4�Խ nѽ_8ݽ����}����>m+��S4�x�5��Y/��c"������&;ֽ���m��������a�D�H��37��,�Ol&��!&��#+�Ŭ5��xF���^�Z������`=���Gҽu�����?� �37.�pg5���4�#�,����*u�f��#o߽
ҽ�ӽ�B佚4 �2^��+"��)/�+�5��r4�r�+����,�
�u�@�ʽ����er��9�w�5�X��-B���2�7�)��%�>?'�{.��:�˱M���h�(���EH��ٯ���X޽�0�++���%�Bk1�%6���2��(���W�����fٽ�нv�׽���ҿ��0�D'��'2��  �  i�#�>� ���M�+���.�ؽ�	���%���g��k%{�$�`��FL�L>�Ԣ5��C3���6���@��@P� �e����������R��q½xu߽����0�n���!�c#��A�i|��,�>n콜<ӽ0�ý�����ʽiRཎ���Sg�1�*�!��j#��x����p6�x�νeE��1Û��\���}q�EY���F��:��4���3��9��)E�k�V��nn�uo���d��Lo��݆˽��齟f����R��)#�#^"�z1�R��� ��1��̽N0��+�½��н|D��y�G�M�� #�Ut"�������� ����5ŽJ����ٔ�����)�h�KR��B�۵7��P3�h5�M�<�4WJ�8�]���w��R��F������Wս�%��\f	����U �У#�צ �Ŕ��'
��!��M�ڽ��ǽJ1��	ƽ�ؽQ��K��1C������#��� ��	�y�Ο���ؽ-��$ ���a��p{�Iw`�-8L��=�?�5�L43�;�6�۟@��2P���e����������N��½�r߽=����.��l�>�!��a#��?�z��)��g�h5ӽX�ý9���f�ʽ�I�����c��O�!�2g#�@u���^��1�]�ν�A��W����Z���zq�'Y���F�P�:�C!4���3���9��.E�U�V��un��s��@i���t��Ќ˽&��4j����{��~-#��b"�P6�J��� ��;�	�̽�9��I�½h�н.L�X}�?��O��"#�5v"�V��F��z����89Ž ���ߔ�!ǂ��h�\ZR��B�)�7�Wa3��5���<�gJ�e�]��w��Y������y���]սS,���i	����� �y�#�� �E��^-
��-���ڽu�ǽ>���"ƽ�(ؽ��򽎆��G�����  �  ̛��D�b{����_����ѽ,���I��G|������&{��he���T�y�J�!�G�XLL��X�*�i��K�������KK�����l�ֽ��2� ��	�����9��|	��f �)齵|н3Ȼ��������(�߇ƽ�ݽ�������������%��l%���h�=�ʽ\���Bt��DK�����.[s�8_��P���H�UH�siO�gK]�3�p�Ň��0���s����t��edȽ��ݽ���J��t)�x���+�
���G��Ļ���Ƚ�t�������1��+⹽��ͽaQ潋Y���������>�J�	������ٽ��ý�P��!ڞ�
R�������l���Y��3M�m�G�f�I��QS�;c��sx����絗�>L���㺽1sϽ�J彊���4�����S��	������U��vؽi���-���)��\����ǿ���ս�����K�
���-A�]x�������|�ѽ����C��
v��ō��P{��Ye���T��J���G�<L�"�W�o�i�E���������F��/���N�ֽa���� �z	�R��38��z	�ld ���kvн0���K ��v����괽pƽ��ݽ��������������8��. ��-d�;�ʽ����xq��I����Ys��7_��P�Q�H�~WH�mO�#P]��p�H���G��� ���3z��CjȽ��ݽ������-�˜��0����`Q����ཫ�Ƚ�~������:��r깽-�ͽ X�u_��H�����|@��	����n	��ٽ3�ýV������X��ʱ��T$l���Y��DM���G���I��bS�hKc��x�
��缗��R��G꺽�yϽxQ彂�������˴������ a񽓂ؽ����f9��6��g	��uӿ���ս����w�
��  �  ������T��S�[޽,:ҽ��Ž�k���L��f���������/t��\g�p�c���i��x�m(�� ������ E��sB�� �Ƚ�Խ����6뽣��L���j�5��kڽ�Jǽj���ad���\���u������ݫ�io��^3ҽ������3���H*���"�ʑ�V4ڽa*ν����4��ɧ����\������&#o���d�,dd���m�x��G��g���FC�����nn���̽&�ؽ�W��.�Ȳ���	�����>�'FԽk���1���w1����������;䡽Ū���Žegؽ�a�ߪ�J��Ѩ�=�.���:ֽʽ����6���Q<��ጕ��|��.�z���j���c�bf�C�r��1������"��dǪ�x���M�Ľ��н��ܽE��U������"������/�ͽ�
��a<���ӛ����-嚽����e巽��˽�<޽B��h������o����޽�4ҽ9�Ž�e��AF��d�������y��Pnt�'Kg��rc��ui�rx�� ��������Y?��|=��˸Ƚ��Խ{��4��	��I��Vg�<��[fڽ.EǽH����]��sU���m�������ի�Zg��}+ҽ�㽩��w���$���ｶ���/ڽ{&ν����{���Ƨ�-��[�������c#o�=�d��fd�K�m�-��J��╘�RG�������s����̽�ؽ�^�[6���c������G当OԽ���������:���Ǘ�����L졽)����ŽHmؽg�m��N�����RA�0��_?ֽ�ʽa�������pC������L�����z���j��c�tf�ޠr�:�����*��yΪ�*�����Ľ��н^�ܽ��罀������!��W������ͽ����G���ߛ�d&���𚽏����﷽@�˽�E޽G���  �  үҽ�Cٽ��ܽ�c޽�Y޽Z�ܽ��ؽK8ҽ(�ǽ⍺�n�����%T�������+���"��-�R䞽����Ž�E�ʽԽ�ڽQDݽy{޽d3޽Kܽqؽ��н�Ž����p�����O����Ԅ��`��d������r��#<��3��_̽�>ս��ڽ"�ݽe�޽��ݽ��۽h׽v.Ͻ��ý#����ɥ�S���>Ԋ�������0ˉ�]6������γ�_T½_ν�[ֽ�\۽��ݽN�޽��ݽd'۽S�սsͽƒ���%��{s��XI������sQ��[��р��E���4^����ĽI�Ͻ=k׽=�۽�޽ρ޽kxݽ�ڽ��ԽC�˽2N��/W��=����J��T쇽�A�����r��♽9L���฽՚ƽ�:ѽ�^ؽ�nܽ$<޽Ro޽�ݽX�ٽ��ӽP�ɽ�񼽇������W:��浆�z��K����뎽�U����8V����Ƚ�ҽ�=ٽ(�ܽ�^޽hT޽��ܽ�ؽ*2ҽv�ǽ����������7K��c����"�����-落�۞� ���U����ʽ��ӽ(	ڽI@ݽ�w޽30޽Hܽ8ؽ�н�Ž����k������|���̈́� Y��_\������+k���4�����.X̽8սۺڽ��ݽ|�޽��ݽ"�۽1׽�+Ͻ��ý����ɥ�輖�`Ԋ�������̉��8���
��Hҳ�`X½�ν�`ֽsb۽ �ݽ�޽��ݽ*/۽�ֽ�ͽ��������N.���|��mR��`����Y���b�����Ү��d���Ľ��Ͻ�o׽X�۽�޽.�޽;}ݽx�ڽ��Խ)�˽�U���_��%����S������/K��#������꙽~T��M踽�ƽ�Aѽ�dؽ�tܽUB޽�u޽�&ݽ��ٽ�ӽ�ɽ����������LE������$��/
��v����_�������^��U�Ƚ�  �  -"��֮ƽ]�ҽ��޽-�齤� (��C^��d��#TݽG�ʽ߶�i���8���&0���_���'��p*��U�ν��[��V��׳��xr��V��,ܽ 4н��ý0E��-��Me��t䎽+����q�0f�[�c�.nk�G�{�o3��S��E���w��)\��w�ʽ��ֽ�⽋��;��D���E򽂢��e׽q�ýJ����3��,p�������ٟ���������Tս5��e�"��ev�����u��{3ؽ3̽?���n岽�~��*͗�������}���l��!d��<e���o��T���k��eښ�-����е�6�½��ν��ڽ�'�b�ｺX��n���Po�W���ѽhO��)ꪽi���N��u���� �����S_Ƚ�_۽��꽓��@��ɲ���꽗�58Խ�Ƚ����I���W򠽟K���r��fw�t�h��dc�W�g�adu�����Α��k��U�����ʨƽ��ҽX�޽��8��9"���W��t�뽁Lݽ��ʽ�ֶ�����px��6&���U�����C!����ν��/T��P�������m��R�m)ܽ�0н\�ýwA��	���`��4ߎ�X���_�q���e��c�w_k�d�{�,���K��H���q���U����ʽl�ֽD��T�콏���@��'C�y�罁d׽��ý䬰��3���p��%����۟��������VXս*�Zj�'���{��ٻ��㽛:ؽ�"̽A¿���i���֗�������}�"�l��2d�Me���o��[��Ar��<���s����յ���½��νn�ڽ�,潛�ｗ^������vｉ���$ѽ�X�����;s��Y��m���Y*��=ƴ��gȽ�g۽ʎ�I��eF��и��꽷	཭>Խ�ȽG�������B���$U���|���zw���h��yc���g�Gxu�V)��fב�t������  �  �G��k6���ӽ���"��x���w�\����
�!*��F�tԽ�Ǿ��|���B���ܲ�.ý��ٽ6��`����������*�����6��Hν�ҹ�yX���ݖ��E���2w�W?b�t�R��I���G���M���Z�Lm�{d��a&��Yȟ��Z��H�Ľ0Nڽz9�DF�/
��[�����<�������&�̽� ���ۭ�@�� J��� ʽ�$⽪���NV��c�A����
�XH�$�򽪷ܽT;ǽg��Ϛ�����ʃ���o��U\�l�N�� H�>�H�_CQ��.`���t�����"��g��b����˽��὜M��9<�4����<t��e�]����ܽmTŽ80���k���r�����$�ѽ{�� � �	�}U�
��;���& �d��qսk��"B��c ��L茽�%�D�h��"W���K��G��J�Q�U��lf��m|��T���W��TA���0��P	ӽU���������t�!��$�
�(&�>�?kԽ½���r��8��Ҳ��ý��ٽ���[�,��\����r(�6���P�EνϹ��T���ٖ��@���(w��3b��R�ۋI�'�G���M�d�Z��=m��]����������T����ĽIڽ�4�8D�<-
�;Z�����;�z�����ş̽
��cܭ�SA���K���"ʽ\'����CX��e������
�ZK���򽤾ܽ�Bǽ�n������^ˑ��Ӄ�d�o�Gg\��N�31H�
I�NRQ�i<`�Z�t��Ć�(��l�������˽B�ὮR��?�Y�;��0x�Fj��f����ܽ�^Ž�:���v��W}��ü���ѽ�� ���	��X�&��,���) ��i��wսr��MI��/(�������7�7�h�\6W���K��G��K�>�U��~f��~|�i\���^���  �  -l��0���Eaڽ�a������� !���#���ϙ�g���@��ֽRwŽ�M���\ȽM"ܽ2���]�
��=��!���#�!�������_n�}�ӽ ���tf��lU���:v���\��zI�c2<�+�4�s3��-8�d�B�AiS�&j�\������*T����ƽ���S��%w�6��"��"����
E�����罿�ϽoB½y���<�ͽp��A� �������"�#��T�����t��|�ɽG
��G:���|��u�l�.�U�VD��9���3�L4��;�9�G�29Z��s��T����q���gн������7��M#�e�!�ou�D���"����޽��ɽ���]4ĽhcԽ���] �N0�1���x#���!�����f�����~�ݽ����v����������Hqd�l*O���?��6��*3�J�5���>��-M���a��|� m���e�������[ڽZ\��}��ѧ�!�6�#�m�������7��ֽ�lŽ�B���QȽ�ܽ������
�:9��� �u�#�����l��/j򽏰ӽ@���rb��!Q��y1v�L�\�ZoI�X&<�e�4��e3��8���B��[S��j�ڥ������VN����ƽ�����&u�w���"���"����TD���������Ͻ"C½������ͽ��佪� ���������"��#���K��1��P���ɽ���BB������E�l�&�U�gD�R9���3��[4�\;��G��EZ�js�Z������B����kн���X�������
�#���!�z�:��6-����޽�ʽ���2?Ľ�mԽy���m4���T|#���!�����i�?���]�ݽ����G��핑�� ��l�d�z<O�J�?�"�6��=3�
�5���>��>M���a���|��s���  �  bȢ�!���佇i��*��(�]�2�j$6���1�mL&��:�C����0�ֽ
�н�Mڽ�/񽸜�z�TW)��Z3�&6���0���$��&���Mܽ�湽М�Yz���g�jlL��9�:�-�'���%�]�)�%�3�V5C��"Z��y�n����B��\n̽q�G����?W,���4�r�5���.��L!�b�,������(=ӽ!aҽ_��6���l����`-�Q5�S05�f�-�Q�����V���Jн;����^��<�}�� ]�&OE�M�4�E�*���%���&��w,���7�|�I�(�c��5���뙽_��x>ؽ����I�A#�t�/�$�5��4���*������
��Y���0ܽ6ѽu~ս�:����_F��$���0�s6��x3�7�)�J���*�轇�Ľ�٥�����#�q��LT��?�\�0���(��%���'�?�/�F1=�ƎQ��n��(��]¢��������f�(�(�[�2�!6���1�8H&��5�;�����ֽ��н:Bڽj$�Y��o��R)��V3�u6���0���$�U$����Iܽ~⹽�˜� v����f�9bL�ޤ9�gw-���&���%��)��z3��'C��Z�S�y�a���=��i̽�������U,�/�4�;�5���.�L!��a�ӛ�����=ӽ[bҽ!�����m�ʊ�zb-��5��25��-�?��9��]���QнĐ���f��k�}�;1]��_E���4���*��	&�П&�f�,�=	8�
�I�ǣc�;����d��kCؽ����*D#���/�	�5�K
4�e�*�����
�$e��1<ܽ}Aѽ��սfE�����J��$�B�0��6��{3��)� �ǎ�ӱ轒�Ľ�ॽƣ����q�s]T�*?�c�0��(�T�%�(���/��A=�Z�Q�<)n�/���  �  �f��>DŽ��콧�!��2���>���B�r>�f�1�� �|��~�����7ܽ�?潵D��C'�g9$�"�4�^�?��B���<�m/�}���-���h-���ǜ�!$���_���C�01�_^%��0����!��++���:��%R���s���������ѽU��m4���'���7�*0A�`7B��:��),�����������޽j�ݽf�����;*��^9�4�A�J�A�0(9���)�������\Dֽ�����t��ex��FU�&�<��},��"��5�D��Y^$�?�/��uA��\�ͭ��픙��;���0߽���"B�҈-���;���B��@�E~6��?&�d>��]�|P��Oܽj��hz��b�
�����/�Q
=���B�`�?�V�4�hE#�5i�X���fɽ�Ц�BV3k��L��6�ޔ(�
� �_��n �l'�M�4�9CI��4g�?���`���>Ž[��  �z!�A�2���>�"�B��>� �1�� �[��������⽎�۽�3�?9���!�;4$�`�4��?�D�B�1�<�'j/����+�ֺ�L)���Ü������_�o�C�+%1��R%��$�	���!�>+�W�:��R�A�s��������ѽ���B2���'��7��.A�-6B�)�:�),���q��ڼ｡�޽��ݽ'�B�w��X=*��`9�a�A���A��*9���)�>��C���xKֽ����z|��gx��VU���<��,�B�"��E�U���l$���/��A�/\�:�������@���5߽,���D���-�K�;���B�]�@�&�6��D&��C��c�3\�t[ܽ�	�A���v�
�f��T�/�=���B�k�?�%�4�H#��k�ߩ�lɽ�֦�4���]Bk��'L�ܜ6�y�(��� �[��#" �&}'���4�|RI��Bg��E���  �  �ꣽiǽ�>�w�uU$�y�6�+KC�.dG��~B�'�5�_�#����jb��)�潩�߽q���x+�-�'�9�5VD�CG��3A��63�x��&s	���'���$��-����]��rA�L�.���"�̦�����h��(��	8�]�O�~r��l���׮��+Խ��������+���;�L�E� �F���>�I0����ƭ	�=8���|���b�1�����.�j�=��IF�4F��N=��'-��b����Y�ؽ����k��w�v��R��*:��)�. �I��;���!���,���>���Y�������*���?��3���@�x@1���?��G�EE�p�:�}�)�3S����Q�콎4�i��"������R!���3��hA�FG�m,D���8��&���F��Q˽�s��~����]i���I��3���%���R�����$�H2�|�F��Fe��ه��䣽� ǽ�9�t��R$���6�!HC��`G��zB�ۡ5���#����kW�������߽Re� ��%���'�N9��QD�1?G�<0A��33����p	�ɤ�������ɒ����]��hA�d�.�.�"����܁��[��|(���7���O��q�g��$Ү�Z&Խ������+���;�ڢE�κF��>��0�w����	�l8��X}���#��U�����.�U�=�'LF�y6F�4Q=��*-��e�J��o�ؽ~����s��i�v�V
S�N;:�Z�)�B' ��� J���!�$�,�!�>�Y�Y���Gƙ�1���R������C��C1�F@��G��E�[�:���)��X������H@����-�����xW!�(�3�LlA��IG�w/D�x�8���&��������V˽z��`����li���I���3�H&��"��d������$�u2���F��Te�<����  �  �f��>DŽ��콧�!��2���>���B�r>�f�1�� �|��~�����7ܽ�?潵D��C'�g9$�"�4�^�?��B���<�m/�}���-���h-���ǜ�!$���_���C�01�_^%��0����!��++���:��%R���s���������ѽU��m4���'���7�*0A�`7B��:��),�����������޽j�ݽf�����;*��^9�4�A�J�A�0(9���)�������\Dֽ�����t��ex��FU�&�<��},��"��5�D��Y^$�?�/��uA��\�ͭ��픙��;���0߽���"B�҈-���;���B��@�E~6��?&�d>��]�|P��Oܽj��hz��b�
�����/�Q
=���B�`�?�V�4�hE#�5i�X���fɽ�Ц�BV3k��L��6�ޔ(�
� �_��n �l'�M�4�9CI��4g�?���`���>Ž[��  �z!�A�2���>�"�B��>� �1�� �[��������⽎�۽�3�?9���!�;4$�`�4��?�D�B�1�<�'j/����+�ֺ�L)���Ü������_�o�C�+%1��R%��$�	���!�>+�W�:��R�A�s��������ѽ���B2���'��7��.A�-6B�)�:�),���q��ڼ｡�޽��ݽ'�B�w��X=*��`9�a�A���A��*9���)�>��C���xKֽ����z|��gx��VU���<��,�B�"��E�U���l$���/��A�/\�:�������@���5߽,���D���-�K�;���B�]�@�&�6��D&��C��c�3\�t[ܽ�	�A���v�
�f��T�/�=���B�k�?�%�4�H#��k�ߩ�lɽ�֦�4���]Bk��'L�ܜ6�y�(��� �[��#" �&}'���4�|RI��Bg��E���  �  bȢ�!���佇i��*��(�]�2�j$6���1�mL&��:�C����0�ֽ
�н�Mڽ�/񽸜�z�TW)��Z3�&6���0���$��&���Mܽ�湽М�Yz���g�jlL��9�:�-�'���%�]�)�%�3�V5C��"Z��y�n����B��\n̽q�G����?W,���4�r�5���.��L!�b�,������(=ӽ!aҽ_��6���l����`-�Q5�S05�f�-�Q�����V���Jн;����^��<�}�� ]�&OE�M�4�E�*���%���&��w,���7�|�I�(�c��5���뙽_��x>ؽ����I�A#�t�/�$�5��4���*������
��Y���0ܽ6ѽu~ս�:����_F��$���0�s6��x3�7�)�J���*�轇�Ľ�٥�����#�q��LT��?�\�0���(��%���'�?�/�F1=�ƎQ��n��(��]¢��������f�(�(�[�2�!6���1�8H&��5�;�����ֽ��н:Bڽj$�Y��o��R)��V3�u6���0���$�U$����Iܽ~⹽�˜� v����f�9bL�ޤ9�gw-���&���%��)��z3��'C��Z�S�y�a���=��i̽�������U,�/�4�;�5���.�L!��a�ӛ�����=ӽ[bҽ!�����m�ʊ�zb-��5��25��-�?��9��]���QнĐ���f��k�}�;1]��_E���4���*��	&�П&�f�,�=	8�
�I�ǣc�;����d��kCؽ����*D#���/�	�5�K
4�e�*�����
�$e��1<ܽ}Aѽ��սfE�����J��$�B�0��6��{3��)� �ǎ�ӱ轒�Ľ�ॽƣ����q�s]T�*?�c�0��(�T�%�(���/��A=�Z�Q�<)n�/���  �  -l��0���Eaڽ�a������� !���#���ϙ�g���@��ֽRwŽ�M���\ȽM"ܽ2���]�
��=��!���#�!�������_n�}�ӽ ���tf��lU���:v���\��zI�c2<�+�4�s3��-8�d�B�AiS�&j�\������*T����ƽ���S��%w�6��"��"����
E�����罿�ϽoB½y���<�ͽp��A� �������"�#��T�����t��|�ɽG
��G:���|��u�l�.�U�VD��9���3�L4��;�9�G�29Z��s��T����q���gн������7��M#�e�!�ou�D���"����޽��ɽ���]4ĽhcԽ���] �N0�1���x#���!�����f�����~�ݽ����v����������Hqd�l*O���?��6��*3�J�5���>��-M���a��|� m���e�������[ڽZ\��}��ѧ�!�6�#�m�������7��ֽ�lŽ�B���QȽ�ܽ������
�:9��� �u�#�����l��/j򽏰ӽ@���rb��!Q��y1v�L�\�ZoI�X&<�e�4��e3��8���B��[S��j�ڥ������VN����ƽ�����&u�w���"���"����TD���������Ͻ"C½������ͽ��佪� ���������"��#���K��1��P���ɽ���BB������E�l�&�U�gD�R9���3��[4�\;��G��EZ�js�Z������B����kн���X�������
�#���!�z�:��6-����޽�ʽ���2?Ľ�mԽy���m4���T|#���!�����i�?���]�ݽ����G��핑�� ��l�d�z<O�J�?�"�6��=3�
�5���>��>M���a���|��s���  �  �G��k6���ӽ���"��x���w�\����
�!*��F�tԽ�Ǿ��|���B���ܲ�.ý��ٽ6��`����������*�����6��Hν�ҹ�yX���ݖ��E���2w�W?b�t�R��I���G���M���Z�Lm�{d��a&��Yȟ��Z��H�Ľ0Nڽz9�DF�/
��[�����<�������&�̽� ���ۭ�@�� J��� ʽ�$⽪���NV��c�A����
�XH�$�򽪷ܽT;ǽg��Ϛ�����ʃ���o��U\�l�N�� H�>�H�_CQ��.`���t�����"��g��b����˽��὜M��9<�4����<t��e�]����ܽmTŽ80���k���r�����$�ѽ{�� � �	�}U�
��;���& �d��qսk��"B��c ��L茽�%�D�h��"W���K��G��J�Q�U��lf��m|��T���W��TA���0��P	ӽU���������t�!��$�
�(&�>�?kԽ½���r��8��Ҳ��ý��ٽ���[�,��\����r(�6���P�EνϹ��T���ٖ��@���(w��3b��R�ۋI�'�G���M�d�Z��=m��]����������T����ĽIڽ�4�8D�<-
�;Z�����;�z�����ş̽
��cܭ�SA���K���"ʽ\'����CX��e������
�ZK���򽤾ܽ�Bǽ�n������^ˑ��Ӄ�d�o�Gg\��N�31H�
I�NRQ�i<`�Z�t��Ć�(��l�������˽B�ὮR��?�Y�;��0x�Fj��f����ܽ�^Ž�:���v��W}��ü���ѽ�� ���	��X�&��,���) ��i��wսr��MI��/(�������7�7�h�\6W���K��G��K�>�U��~f��~|�i\���^���  �  -"��֮ƽ]�ҽ��޽-�齤� (��C^��d��#TݽG�ʽ߶�i���8���&0���_���'��p*��U�ν��[��V��׳��xr��V��,ܽ 4н��ý0E��-��Me��t䎽+����q�0f�[�c�.nk�G�{�o3��S��E���w��)\��w�ʽ��ֽ�⽋��;��D���E򽂢��e׽q�ýJ����3��,p�������ٟ���������Tս5��e�"��ev�����u��{3ؽ3̽?���n岽�~��*͗�������}���l��!d��<e���o��T���k��eښ�-����е�6�½��ν��ڽ�'�b�ｺX��n���Po�W���ѽhO��)ꪽi���N��u���� �����S_Ƚ�_۽��꽓��@��ɲ���꽗�58Խ�Ƚ����I���W򠽟K���r��fw�t�h��dc�W�g�adu�����Α��k��U�����ʨƽ��ҽX�޽��8��9"���W��t�뽁Lݽ��ʽ�ֶ�����px��6&���U�����C!����ν��/T��P�������m��R�m)ܽ�0н\�ýwA��	���`��4ߎ�X���_�q���e��c�w_k�d�{�,���K��H���q���U����ʽl�ֽD��T�콏���@��'C�y�罁d׽��ý䬰��3���p��%����۟��������VXս*�Zj�'���{��ٻ��㽛:ؽ�"̽A¿���i���֗�������}�"�l��2d�Me���o��[��Ar��<���s����յ���½��νn�ڽ�,潛�ｗ^������vｉ���$ѽ�X�����;s��Y��m���Y*��=ƴ��gȽ�g۽ʎ�I��eF��и��꽷	཭>Խ�ȽG�������B���$U���|���zw���h��yc���g�Gxu�V)��fב�t������  �  үҽ�Cٽ��ܽ�c޽�Y޽Z�ܽ��ؽK8ҽ(�ǽ⍺�n�����%T�������+���"��-�R䞽����Ž�E�ʽԽ�ڽQDݽy{޽d3޽Kܽqؽ��н�Ž����p�����O����Ԅ��`��d������r��#<��3��_̽�>ս��ڽ"�ݽe�޽��ݽ��۽h׽v.Ͻ��ý#����ɥ�S���>Ԋ�������0ˉ�]6������γ�_T½_ν�[ֽ�\۽��ݽN�޽��ݽd'۽S�սsͽƒ���%��{s��XI������sQ��[��р��E���4^����ĽI�Ͻ=k׽=�۽�޽ρ޽kxݽ�ڽ��ԽC�˽2N��/W��=����J��T쇽�A�����r��♽9L���฽՚ƽ�:ѽ�^ؽ�nܽ$<޽Ro޽�ݽX�ٽ��ӽP�ɽ�񼽇������W:��浆�z��K����뎽�U����8V����Ƚ�ҽ�=ٽ(�ܽ�^޽hT޽��ܽ�ؽ*2ҽv�ǽ����������7K��c����"�����-落�۞� ���U����ʽ��ӽ(	ڽI@ݽ�w޽30޽Hܽ8ؽ�н�Ž����k������|���̈́� Y��_\������+k���4�����.X̽8սۺڽ��ݽ|�޽��ݽ"�۽1׽�+Ͻ��ý����ɥ�輖�`Ԋ�������̉��8���
��Hҳ�`X½�ν�`ֽsb۽ �ݽ�޽��ݽ*/۽�ֽ�ͽ��������N.���|��mR��`����Y���b�����Ү��d���Ľ��Ͻ�o׽X�۽�޽.�޽;}ݽx�ڽ��Խ)�˽�U���_��%����S������/K��#������꙽~T��M踽�ƽ�Aѽ�dؽ�tܽUB޽�u޽�&ݽ��ٽ�ӽ�ɽ����������LE������$��/
��v����_�������^��U�Ƚ�  �  ������T��S�[޽,:ҽ��Ž�k���L��f���������/t��\g�p�c���i��x�m(�� ������ E��sB�� �Ƚ�Խ����6뽣��L���j�5��kڽ�Jǽj���ad���\���u������ݫ�io��^3ҽ������3���H*���"�ʑ�V4ڽa*ν����4��ɧ����\������&#o���d�,dd���m�x��G��g���FC�����nn���̽&�ؽ�W��.�Ȳ���	�����>�'FԽk���1���w1����������;䡽Ū���Žegؽ�a�ߪ�J��Ѩ�=�.���:ֽʽ����6���Q<��ጕ��|��.�z���j���c�bf�C�r��1������"��dǪ�x���M�Ľ��н��ܽE��U������"������/�ͽ�
��a<���ӛ����-嚽����e巽��˽�<޽B��h������o����޽�4ҽ9�Ž�e��AF��d�������y��Pnt�'Kg��rc��ui�rx�� ��������Y?��|=��˸Ƚ��Խ{��4��	��I��Vg�<��[fڽ.EǽH����]��sU���m�������ի�Zg��}+ҽ�㽩��w���$���ｶ���/ڽ{&ν����{���Ƨ�-��[�������c#o�=�d��fd�K�m�-��J��╘�RG�������s����̽�ؽ�^�[6���c������G当OԽ���������:���Ǘ�����L졽)����ŽHmؽg�m��N�����RA�0��_?ֽ�ʽa�������pC������L�����z���j��c�tf�ޠr�:�����*��yΪ�*�����Ľ��н^�ܽ��罀������!��W������ͽ����G���ߛ�d&���𚽏����﷽@�˽�E޽G���  �  ̛��D�b{����_����ѽ,���I��G|������&{��he���T�y�J�!�G�XLL��X�*�i��K�������KK�����l�ֽ��2� ��	�����9��|	��f �)齵|н3Ȼ��������(�߇ƽ�ݽ�������������%��l%���h�=�ʽ\���Bt��DK�����.[s�8_��P���H�UH�siO�gK]�3�p�Ň��0���s����t��edȽ��ݽ���J��t)�x���+�
���G��Ļ���Ƚ�t�������1��+⹽��ͽaQ潋Y���������>�J�	������ٽ��ý�P��!ڞ�
R�������l���Y��3M�m�G�f�I��QS�;c��sx����絗�>L���㺽1sϽ�J彊���4�����S��	������U��vؽi���-���)��\����ǿ���ս�����K�
���-A�]x�������|�ѽ����C��
v��ō��P{��Ye���T��J���G�<L�"�W�o�i�E���������F��/���N�ֽa���� �z	�R��38��z	�ld ���kvн0���K ��v����괽pƽ��ݽ��������������8��. ��-d�;�ʽ����xq��I����Ys��7_��P�Q�H�~WH�mO�#P]��p�H���G��� ���3z��CjȽ��ݽ������-�˜��0����`Q����ཫ�Ƚ�~������:��r깽-�ͽ X�u_��H�����|@��	����n	��ٽ3�ýV������X��ʱ��T$l���Y��DM���G���I��bS�hKc��x�
��缗��R��G꺽�yϽxQ彂�������˴������ a񽓂ؽ����f9��6��g	��uӿ���ս����w�
��  �  i�#�>� ���M�+���.�ؽ�	���%���g��k%{�$�`��FL�L>�Ԣ5��C3���6���@��@P� �e����������R��q½xu߽����0�n���!�c#��A�i|��,�>n콜<ӽ0�ý�����ʽiRཎ���Sg�1�*�!��j#��x����p6�x�νeE��1Û��\���}q�EY���F��:��4���3��9��)E�k�V��nn�uo���d��Lo��݆˽��齟f����R��)#�#^"�z1�R��� ��1��̽N0��+�½��н|D��y�G�M�� #�Ut"�������� ����5ŽJ����ٔ�����)�h�KR��B�۵7��P3�h5�M�<�4WJ�8�]���w��R��F������Wս�%��\f	����U �У#�צ �Ŕ��'
��!��M�ڽ��ǽJ1��	ƽ�ؽQ��K��1C������#��� ��	�y�Ο���ؽ-��$ ���a��p{�Iw`�-8L��=�?�5�L43�;�6�۟@��2P���e����������N��½�r߽=����.��l�>�!��a#��?�z��)��g�h5ӽX�ý9���f�ʽ�I�����c��O�!�2g#�@u���^��1�]�ν�A��W����Z���zq�'Y���F�P�:�C!4���3���9��.E�U�V��un��s��@i���t��Ќ˽&��4j����{��~-#��b"�P6�J��� ��;�	�̽�9��I�½h�н.L�X}�?��O��"#�5v"�V��F��z����89Ž ���ߔ�!ǂ��h�\ZR��B�)�7�Wa3��5���<�gJ�e�]��w��Y������y���]սS,���i	����� �y�#�� �E��^-
��-���ڽu�ǽ>���"ƽ�(ؽ��򽎆��G�����  �  �(6��O2�dV'��,��V�&t�5L��mC��s���.Ul�kHP��U<��$/�!�'���%���(�6�1��$@��U���s��㍽Kr����ƽ���
��V��M*�y�3���5��=0���#�#Q�v�~��=�Խ�vѽ5Aݽ���V�����lq+��W4�(�5�Q]/��f"�������T?ֽ����S������J�a�l�H��47�i,��j&�S&� +���5��rF�t�^�	��Ż���7���Aҽ�x��\��P� ��2.��b5�	�4�6�,����p��[���d߽4 ҽ3�ӽ�9佲0 ��Z��("�-'/��5�!q4�֭+�F����
���R�ʽ���+m��d�w��X�XB���2���)��%�0/'���-��:��M���h�F����A��>���R޽M-�z'���%��f1�U6���2�h�(�������｡Yٽ��н��׽6������+�V'�`#2�%6�'L2�ES'��)��S��n��F���=�������Hl��:P�qG<�/�(�'���%���(�.1��@� �U�U�s�ߍ��n��~�ƽ$����b��L*�I�3�P�5�<0�m�#�RN�0�!��4�Խ nѽ_8ݽ����}����>m+��S4�x�5��Y/��c"������&;ֽ���m��������a�D�H��37��,�Ol&��!&��#+�Ŭ5��xF���^�Z������`=���Gҽu�����?� �37.�pg5���4�#�,����*u�f��#o߽
ҽ�ӽ�B佚4 �2^��+"��)/�+�5��r4�r�+����,�
�u�@�ʽ����er��9�w�5�X��-B���2�7�)��%�>?'�{.��:�˱M���h�(���EH��ٯ���X޽�0�++���%�Bk1�%6���2��(���W�����fٽ�нv�׽���ҿ��0�D'��'2��  �  ��B�!v>�r2������
�@��T7ý춡������Pe���G�T�3���&����:��H� ��@)�ɖ7���M��Mm��S��ؕ����˽������\$��s5��,@�]�B�<�+�.�"����	����$Uཙ�ܽ�y齚H��R�F'�{A7��@�-\B�0$;�̓,�������ܽoN��x����~�;WZ��E@�%�.�"�#�����Y�r#�_<-�M�=���V��Mz�;����z���xؽ#����̖*� �9���A�]�A�o�8�u>)��n���n���,ݽ�߽�������b-�O;��cB���@�X�6��}&�8�����Z�Ͻ�!��[��+xq���P��9��w*�f�!����KZ�h�%���1�|<E��za�_���a��-&����!`�*���S0��o=���B��t?�}!4��*#�_�e����5��۽�`�1������!�x2��>���B��r>�K2����
���2ýj����GDe���G��3�|�&�^�����	� �3)�"�7���M��Cm�uO��T���Ƀ˽������[$��r5��+@��B�.}<���.�L����	����L��ܽ�p�D��M��A'�==7��@�oXB�� ;���,�*����w�ܽ�J�������~��SZ�_C@�$�.�L�#�K��\�#�*A-�E�=��V�&Vz����f����~ؽt&�=��Ě*�D�9��A�%�A�k�8��C)�*t�������6ݽ4߽�"���;��`-��Q;��eB���@�� 7�&���G����Ͻ�%��e"����q�q�P�ܟ9�K�*���!�A�j���%�2�4KE��a��e��sh���,��K
潤c����W0�ft=���B��y?�I'4��0#���Ə��NC彊�۽�m㽻=����/!�
}2���>��  �  ht��꽧�۽�iŽ,���Z���o���D���"�	���N�ּG�Ǽ|
��Fｼ�D����ʼ�qۼM���	x�y�)�pM�/�y�N7���(����ʽ�߽��6����`ؽV½C)��ꓗ�wz��-����+����㷽�Ͻ�p�7*�_������Խ�鼽o#������`��u8����9��\��g�м�ļ����V����ü5ϼ���ơ �R���4�44[�B&������#�ҽ�F彯Hｱ���$�2jѽ	v��������������P����ƕ�Ⲩ�o����ֽ�V罃��a����vͽ����*����~��Q�W.-��z}����ݼb�˼5���뽼k��]�Ƽ��Լ4��`����O@���i��o��$��1�½��ٽV���V�bY�1�޽8ʽ8����g���v������zV��v]��$!��yǽR�ܽ�E뽅l� ��8�۽�cŽ~&��mU���o�d�D��"�_v	����5�ּc�Ǽ5ӽ�\)��-�ʼ	Yۼ�����m���)��hM�ُy��4��l&����ʽ��߽��2���5\ؽzP½�"��،���r���$���������z۷�~�ν�h��"�f��d��C�Խw伽�������`�>p8�@|���C�弎�мv�ļ�����Z����üM>ϼ
�⼢� �Q��<�4��>[��~#�������ҽ�N�7Qｪ��+.��sѽ���l��'������9����Ε�����D����"ֽ7\���Z��J��tyͽ�"��X.����~�+�Q��8-�~�������ݼ
̼�����	��������Ƽ��Լ;��v,�s����@�j��v��+����½ �ٽ��?`�c�(�޽�ʽ`���t��s���3͈��b��]i��h,����ǽ��ܽ}N��  �  �$�彌;׽�����V���{���m�4D��r#���
�Y/�G2ڼa	˼��¼>���"/ļ��ͼ&�޼�������j*�ӜL��;w�G"�����O�ƽv/۽h����꽏��:�ӽ�K���ʧ���l��������u��*����'��E�ʽ�uݽ�轴}�b���н�q��֠��N/��J�^�^T8�$R�����S/Լ��Ǽ:{��+����ƼscҼO.����u���4�9�Y��v��"�������UEν^�z��4��X߽��̽x���UР��؏�����7����Hf��۽���}ѽ58�k��5��wݽ\gɽ����`���tb|���P��h-�D�=x��m�!ϼC�ļ����EH¼%�ɼ! ؼ���7h��C �Q@�&h����1j��x��ս;�佫 �罔�ٽ[�ŽN���l���勽W��F͊�.q��
���JHý��׽�
�C���!5׽����Q��v���m��(D��f#���
�/� ڼI�ʼD�¼գ��Zļ�ͼ:�޼����W����)�:�L�E5w��������ƽ -۽��罂�꽓��x�ӽfF��}ħ�ջ������ȸ���m������I���ʽ nݽ����v����M�н�l��@���V+����^��N8��M������}-Լa�Ǽ�}���/����Ƽ�lҼ�9漼��}�ė4���Y��|��v��������Lνf���&�齥&߽#�̽0���ڠ��⏽>!��z@��i
���m���Ļ��ѽq=����4��ݽ�jɽ{�������j|���P�Xs-��#��������=ϼA�ļG���g¼��ɼؼ��Vv��Q ��'@�w3h�ӱ��8q�������ս��
�G!�z�ٽ��Žc$��y��K򋽢c���ي�}��?����RýI�׽���  �  �ܽ�׽ȃʽGA��⭠�6���=nh��C���%��K[���y�%�ԼR̼*�ɼWeͼ"�׼p	�3w�ю���+��:K�\|q�Ʀ��:ԥ��컽�	ν�Tٽ��۽�սtƽ�ٲ�j8������2遽A�����ԕ������#���iϽ��ٽ.�۽�
Խ��Ľ_�D蘽a1���d[�D�8����K���S�fN޼B Ѽyʼ�!ʼ'�ϼrܼM�������z5� /W�ׄ�uM��yj����½��ҽ�)۽{�ڽJ�н�A���׫�З�8��Y(��{1��z ��������foĽ��ӽҁ۽�ڽ)�Ͻ|-��J`��#0��ev�)O���.�'��W'�Q]��
ټ�μJ�ɼ�W˼,OӼ�;⼂$��!����"���?���c�(�����QԴ�ÚȽ8sֽ�ܽTHؽ�̽�����ꤽ�����
�~�⒃�Z��餢��j��8;ʽP׽5ܽ�׽j}ʽa;��G�������-ch���C���%�m���@��^�t�Լ,�˼�ɼ�Hͼ�{׼���nk�F��u�+��2K��uq�ݣ���ѥ�껽ν�Qٽ��۽�սRoƽQԲ�!2�������ၽb���醽}̕�q������#bϽ?�ٽT�۽mԽĝĽ:믽�㘽s-��H^[���8�d}�$���O�L޼� Ѽ�{ʼ�&ʼ(�ϼ7{ܼ���l����܃5�@9W�A���S��Uq���½�ҽ�1۽W�ڽ�нK��"᫽�ٗ��A���1��C:���(��c��߈��euĽ��ӽf�۽�ڽޭϽ1���c��4���v��'O��/���Z4�Ly�S(ټx3μ��ɼ9w˼/nӼ�Y��A��]���#��?��d�������۴���Ƚ�{ֽ�ܽQRؽf̽����m������������������*��揤�t���Dʽ�X׽�  �  ?(ƽX�½ya��iѨ�����Ã�o|d���E��r,�����������m�{�ܼ^�ټ�޼��鼧W��z0�m&���1�(AL�5�k�)���G�������7��.2Ľ��Ž�����ಽ-ա��鏽������n���j�Nw�Z���������x����ĽW�Ž������`䢽n6��l{�=�Y���<�k%�+��t����#?���ڼ�]ڼ���
��Q�K�"�b�9�e5V�ow�����נ��뱽�羽�Ž��ĽK��Mz��ٽ���V��.�y�:sk�hBm�\�~� ���˟����f���.�Ž��Ľ񄼽oj��.Ü��q�o�
O�Q4�B��������A8��޼'�ټq�ۼ��伳+��o_����)�0�B���`������f���٦�#ֶ�����#ƽ��½Ǽ���§�����;��-s�y<j�=jq���������p˥�c+������� ƽu�½/[���˨�|���l���Aqd�
�E��f,����)���o���O�Inܼ'�ټ�޼ ���<��$�M��1��8L���k�݇�w���ޕ��c4��2/Ľ��Ž�����۲��ϡ��㏽����>vn�N�j�>w�@���ﺙ����謺��Ľ��Ž����睳�Sߢ��1��Xd{���Y���<�/%�d(��r����?�h�ڼdbڼ�%��n��X�3�"�k�9��?V�]zw�����ޠ�󱽡ﾽa�Žc�Ľ[������KǛ�`��֗y�V�k��Sm���~�u��Sҟ��#������чŽ��Ľǈ��(n���Ɯ���l�o��O�C\4�kN�f�������V뼼߼W�ټ��ۼ{�伳J��kn�v���)���B���`�/���~m���ঽ�ݶ�=���,ƽ��½1Ƿ��ͧ��ŕ�hG��Es�xTj�q�װ���˓�xե��4������  �  P��m�������ᙽ����j���e�o�N��:�/�'��$���
��� ������[�=�����l��4r���+�l>���S�pdk�B�������w���ی���]��c���z⦽����#�����}�͡d���T��Q��B\�ѻq�C���畽Ȕ���ɪ�n6�������`��н������?�v�:�]��{G��3�3]"�e��.��������6�h���!���� ���1�"E��1[���s�����L���/�������NR��b����n��̰��ݑt� ^��kR���S��Ib��z�~���z��L⥽6A��$���:l���ĝ��p�����3&n�EV��@�7�-������������ e������ ��	�{��%���7�%4L��#c�r|�
����P���	���=-��li��,����䵃�ul���X��iQ�/^W�9~i����w������n���������蚤�(ܙ� ���_�K�e���N�Z:���'�`��
�� ����6<�������1��e��+��a>���S�~\k�ͣ�����������Z��ؙ��cަ�/񛽺���_�}�t�d���T���Q�3\��q�t���ߕ�o����ª��/������?[��ḕ�b�����v���]��vG��3�(Z"�c�.� ���7���
o�������g� ���1� +E��;[��s���pS���6���������Z��B����w�����X�t�;(^�F}R���S��Yb���z�!��π���祽�E��h���:p��sȝ�	u��#���/n��!V��@�R�-��$������������3���� ���	�m���&��7��AL��0c�3|�����������5���r��3������ ���Y5l�*�X�ӀQ��tW��i���,���Þ������  �  ;���c������F���[�������p�y]a��FQ��@�k0�� ��5�pH���	�	������#���3�gdD���T���d��Tt�Դ���爽GB��瓽�ƕ�����&��Ȅ�.br��Z��F�#G:���7�8
@��Q���g����`]��_���Pw���"��˖��Jދ�����{���k��	\���K�2;�Ұ*���f��F�
�{
����d��|�(�m-9��I��:Z�\ j�]Vy�� ��������vڔ�s���}q���V��S���@j��JS��xA��>8��n9��D�X�o�o�L���N@��
��������@��Tݏ�æ��W���s�u���f��V�Q2F��|5���%����E��
�]�� �v��5.���>�fO��_��*o��b~�D����B����������* ������.5���Sz�$Kb�ݖL�!P=��r7�s(<��J��_���w���������ӡ���������wU��'��/�p�XQa�	:Q��@��0�O� �b%��7�+�	���������#�l�3��WD�+�T���d��Kt����L䈽?���㓽�Õ�o����"��SÄ��Wr�=�Z��F�;9:���7�3�?���P���g���EV���ّ��p�����u���~ً�����l{���k�n\���K�8
;��*��������
�w}
�����(�49���I��CZ�L
j�bay��&��%���
��┽m����y���_��4���Rj��\S���A��O8�S9���D��*X���o�6����E��Շ��3ƕ�(E��}ᏽ��������v��f�ĶV�=@F���5��%����+W�c
�ļ�	���UE.�{�>�HtO���_��7o��o~�Б��zI��ޝ��_���x�������>���gz�d`b�¬L�Uf=�
�7�0><��J��_�H�w�����ʏ��  �  G(��?��䓆�e���[���q|��e��Z��x6s�3�b���O���<���,��8"��\�#�� 0�]A��?T��f��\v�{���侄��ӆ�H����s��G/�������}�Ŷp���_���L���9�l�*�R"!�VW�\�%�ی2��)D�oW�W�i�<�x�F���0���������!P��mօ�%߂���{��n��\�xsI�b7�(�S? ����%9'��45��LG���Z��Jl�c�z�.j��A���/0��+���� ���o���-���y��\k��{Y�x5F��C4�/�&�N���z �")� 8�րJ���]�4�n���|���:��Z��,�����F���x����w�F�h��SV��C��1�|�$�A,�}i!��<+�@�:���M��`�؂q��~�����D��#x��$���R���!���󮀽o�u�D�e��S�%�?�/�$m#�@��n�"���-���=�\�P���c��s�T!���8����������ш���v�������)s���b�(�O�`�<�{�,�"'"�O���#���/�'�@��0T�P�f�%Pv�������Qφ�����qp���+��|��Z�}�_�p�Y�_�(�L��9�Ѕ*��!�AI��t%�<~2�D��`W���i�5�x�*���q*�����S����K���҅�܂���{��n�&�\��qI��7�J(��@ �A���<'�95�\RG�4�Z��Rl�$�z�o������!6�������'���v��v5��c�y�ymk��Y��FF�NU4�m�&���� �>1)�*8�čJ���]�� o�[�|��������A_��ʬ����������~��"�w��h��cV��!C�Ҳ1���$��>��{!��N+�J�:���M�X�`�7�q�y�~�����K���~������7���~���඀��u���e�I.S�a@��./�K�#�_�-�"���-���=�?Q�|�c�:t��  �  �>b�d�q�7w��-���?K���K��k���鏔�Uf������Tjv��x^���I��;�Ɣ7��>��M�ׯc���{�ʈ��䐽	)���r���^�����+��d�}�Zn��^��N���=�g]-��W����y��'
����#���h&�nr6�D(G�Q�W�Mtg�t�v��킽I��j+��m�������E���̌�$�jSn���V���C�P9�!�8�}KB�l�T���k�����<׋����⥕�ӷ��绐�����<����|x�? i��QY�~�H�z:8�V(�j�����P
���
��l������+���;�~�L���\�(�l���{�Z���7��ؑ�<<���[��f���JӉ��B~��Cf���O�-F?�X�7���:�F�G���[���s� Z�����})��/���(����뎽���{E���ns���c�R�S�gfC�`�2��#�9���(���	�M��ɹ�%j!���0��A��!R�1b���q�iq�������E��F��{�������n_��9���<Zv��g^���I�e�;��7���=���M���c�]�{���7ސ�#���m��2Z���댽H'���}��Rn��^��~N���=�S-��L��x��l��
�ɫ����Z&��d6�G���W�~hg���v��肽���e'���i������}C���ʌ������Qn�"�V�;�C��9���8��NB��T�+�k�ݳ��ۋ�f�������-�������Ǌ�����x�y/i��aY��I�LK8�Y(�i��ɔ��`
�b
�k{�S��l�+�s<�<�L���\���l�'�{�(_���<��aݑ�B��ab������'ۉ��S~��Uf���O�QY?���7���:���G�I�[�>�s��a��e���N0���ĕ�g���,�f���L���|s� d��T��wC���2�#��"=���	������`|!���0���A��0R��  �  ��O�*Bg�Nq���ʍ�׌��� ���«�j���f>������>��.N��Mh���V��Q�u�Y�F�m�M���}��������ϩ�G=��̶�����Kח��ӊ�F{���a�GK���6��%����?	�<M�����
��s}���f�p�����H�.���A��aW���o�ބ�x+���d���ا� Ϭ����_��_����9���y��8a���S�<�R�Q_�Cv�2����7��dI�������������엟�M���7T���Wr�n�Y�+�C�8�0�������m�s���0��F��[�������#�@#�ڻ4���H��%_��x��R��Ho��K����8��*u��e���B��2���@p��M[���Q��xU���e�YU���������fT�����)�����؛�I>���䁽,�i��PR��C=��*�ċ�����M����,����KZ�Z��4����(��;���O�6g��k��Gō�X���B��߼������K7�����`6��@E��@:h�"�V�A|Q���Y�*{m�(����{������_ȩ��6��2����	���җ�xϊ�� {���a�;K��6�y%������\5���}�����b��Y���f����.�[�A�VW���o�%ل�'���`���է�6̬����^������9��y��8a��S���R��!_��v�񍉽);��)M�����v���������������Z��fr�U�Y��D�E�0���a-�F~����������U���*���0��K#���4��H�c/_�j$x�iW��vt��������m?���|������.���;���Tp��a[��Q�S�U���e��g�)��������[���ì��/�����ޛ�eD��끽�j�M_R�vS=�m�*�J��1���`��?��fS�C���l�њ�����(��#;��  �  8uG�rTf��Ʉ�8����Ʃ�h���.ý�ƽ�<��Me��#פ��В�e낽�p��fj��6t�����Ö�Oƨ�A�����½W#ƽ������5䥽�_�������	_�GGA���(�	����+��n@伣�ۼ(ڼT�߼3�Q �6��;b�8�5��,Q�V�q�J���̝�+Q���&����Ľ�SŽ�����<���˞����)L}�g�l���k���z��@���Ĝ�\j��)���}�ĽahŽ�V������ӟ�����xu��}T�>r8�Ə!�pg�?V�F��p�B'ڼ��ڼ�⼂��'��c>&��A>�As[�f}�>A���⣽�s�������Ž��ý����੪�;�������Z)v�A�j�Z o�hd��7א�"Ϣ����y4��l�Ž�ý.���u���գ���҆��j���J�H0��	�fN
�����_�輼�ݼ7�ټL�ܼ缔���9��{��*�-��hG��Hf�)Ą�ǌ��S������v(ýQƽa5��V]��~Τ�Mǒ��Ⴝ��p�]Rj�v"t����8���M���򀸽&�½�ƽ }������ߥ�@[��}����_�	?A���(���������)�zۼ��ټ)g߼��6 �_���U�e�5��!Q���q������ǝ�WM���#����Ľ�QŽ��*;��˞�2���L}���l��k�>�z��B���ǜ��m��綼���ĽmŽ\��z���ٟ�;����u�%�T�|�8��!�~w�vf������^Fڼ�ۼ���L�34�""�?I&��K>�*}[��o}�UF��%製�y��e���� ƽy�ý���1���Ę��ć�)>v��j��4o�Dn�������ע�5����;��J�Ž{�ý<���[���©���؆��j�[�J��V0���0_
������輛�ݼ�ټ��ܼR2�6�����?�Һ-��  �  x�E���j�Y܊�h���yp��#m˽6ؽGܽ��ֽ1Wɽ(P��	���KH��f'���� ,���풽��L׺�o�̽��ؽ�۽D�ս��ǽ裳�+̜������a�x.>���!�-�������K���Ҽ�.˼��ɼ3�μ��ټ)�켼�|"���0� Q��qx��x�������J���sнqaڽQ۽�ӽFlýS[������b���耽Ad���툽�ܘ����	U��l�ѽU�ڽ��ڽe�ѽNt��?)����� }��U���3�ߑ����K)���ۼ%gϼ��ɼ��ʼ��Ѽ�8߼B�����	������:��]�.g��1���*���Ž�Խ��۽�ٽu�ν����^���ϔ��J���]�#C�������J�������gǽ9�սX�۽�ؽ+ͽW���Æ��]��'o�NAI��O*�
X�� �j��Ŷּ��̼V�ɼ�5̼sHռ�t弳�����qO'�vE�s�j��֊��k��ig˽ؽ�
ܽF�ֽOɽLG������C>�� �����!��7㒽+���ͺ���̽�ؽ	�۽�ս�ǽ����ǜ��ۅ�z�a�&>���!����z���]6�ȱҼ\˼üɼ�μ6�ټ���0�[�m�0�9Q�sgx��s��n����F��spн�^ڽ�N۽�ӽ�jý~Z��b���0b���逽se��b�ޘ����BX��$�ѽ��ڽQ�ڽ��ѽ�y��Q/��c
���-}��,U���3�Z��c��-I�Σۼ��ϼ�ʼ�ʼ�ѼS߼���,�	�����:��]�<l��S6��^0����Ž��Խw�۽+�ٽk�νJ���h��|ڔ��U��&s��M������-T������oǽ��ս:�۽x�ؽ1ͽ!Ǻ�����c���3o��NI��]*�\g�K� �l����ּ�ͼ�ɼ"Y̼�jռw�弁���	#��\'��  �  �DF���o�:㏽1ɩ�z�½MAؽ�l��뽎��X�ֽ>½Jn��i����W��)o��䈌��}���c��{ǽ��ڽ���p���佱Խ��������N��	�e�d(>�����V��s��׼�4ɼ|#¼����LżQ�ϼ�S�"c��n�//��)S� �j���e����ʽ��ݽ��TV�~��bн�{���?���2��臽�X�����������νS�߽���8��ڑ߽ͽ�6���D��g ����W���2����D�伉~Ѽ�	Ƽ^��������ȼ�ռ�d�-$�����9:���`�"�������Һ��ѽ��o��tr�ҍܽ�eɽ�ܲ������������`�����I�������b�Խ�@�.���j�X6ڽ��Žk��������t��mJ�I(��I�]��hݼ��̼{�ü�����ü��˼�(ۼE����q %��8F�T�o��ݏ��é��½�;ؽaf���z��ֽ?
½�d��3|��,M��_d��~��]s��|Y����ƽ��ڽ���?��}�Խ����E����I����e��>�ƾ��M��_�W׼ɼ�¼����2ż��ϼJ:�gJ��!b��#/�(S���~��e��pa����ʽl�ݽ	�T�H|ὓaн{��X?���2��/釽�Y��̟��������.ν�߽�������߽�ͽ�<��NK��8'���W���2�l�)�����Ѽ�(Ƽ���3����ȼ;,ռ_}��/����,D:��`�C������:غ�F�ѽ������z���ܽ`oɽ�沽x���̍�����Ik��O�������������ԽnH���6q�H<ڽR�Ž���w���d�t��zJ�$W(��X�&9��a�ݼͼw�üû��j7ü0�˼�Hۼ������%��  �  ��F�5�q��ϑ�`���8�ƽ�ܽ�뽴q�[��E�۽i:ƽ$讽�k��j݌�و�J��v������Q˽u�߽\��,H�齘{ؽ�6��⨦����4{g�|>������F��Ӽ�+Ƽ�G��c��'Z¼��̼߼p���j��/�G8T�NӀ����������νS���W�i��^��%�Խ�h������8��\��ɉ�Q��G'��Uɻ���ҽ���	'�Xｵr佇Eѽ����+��������X���2���~7���ἻRμrü�*��wž��ļ��Ѽ�0�������k:��{b��'���dW���$ֽ���[������ὧ�ͽ��������_��C����ߋ��w���]��w�ýPsٽ�n齗L𽛘���޽|ɽ���.�����v��-K���'�^$��	��#)ڼ��ɼ����3Ƚ��1���yȼ�׼�𼟩
���$���F�ئq�rʑ������ƽY�ܽ؉��j�Ѱ���۽^1ƽlޮ�ia���Ҍ�3Έ�p���u������BH˽��߽B���@�L��uؽw1��D���z���rg��s>���L���2꼳�Ӽ:Ƽ0������
A¼R�̼��޼qW���^���.��-T�R΀�j���z���b�ν��U��ｎ����Խ�g��:���g񔽝]��Lʉ��R��|)��
̻�Ѣҽ��9+���w�Kѽ��������ꑃ��X�~�2�/��V�����rμg1ü�H���⾼�ż:�Ѽ�I缌����v:�(�b��,��K���!]��+ֽx��
 �t���Ὁ�ͽ}�������~j��2
��Pꋽꁘ�rg����ý�{ٽTv�|S�����޽ʁɽ����������v��:K���'�@3�K)��1Jڼ��ɼ�����꽼T��	�ȼ�
ؼ�𼪷
���$��  �  �DF���o�:㏽1ɩ�z�½MAؽ�l��뽎��X�ֽ>½Jn��i����W��)o��䈌��}���c��{ǽ��ڽ���p���佱Խ��������N��	�e�d(>�����V��s��׼�4ɼ|#¼����LżQ�ϼ�S�"c��n�//��)S� �j���e����ʽ��ݽ��TV�~��bн�{���?���2��臽�X�����������νS�߽���8��ڑ߽ͽ�6���D��g ����W���2����D�伉~Ѽ�	Ƽ^��������ȼ�ռ�d�-$�����9:���`�"�������Һ��ѽ��o��tr�ҍܽ�eɽ�ܲ������������`�����I�������b�Խ�@�.���j�X6ڽ��Žk��������t��mJ�I(��I�]��hݼ��̼{�ü�����ü��˼�(ۼE����q %��8F�T�o��ݏ��é��½�;ؽaf���z��ֽ?
½�d��3|��,M��_d��~��]s��|Y����ƽ��ڽ���?��}�Խ����E����I����e��>�ƾ��M��_�W׼ɼ�¼����2ż��ϼJ:�gJ��!b��#/�(S���~��e��pa����ʽl�ݽ	�T�H|ὓaн{��X?���2��/釽�Y��̟��������.ν�߽�������߽�ͽ�<��NK��8'���W���2�l�)�����Ѽ�(Ƽ���3����ȼ;,ռ_}��/����,D:��`�C������:غ�F�ѽ������z���ܽ`oɽ�沽x���̍�����Ik��O�������������ԽnH���6q�H<ڽR�Ž���w���d�t��zJ�$W(��X�&9��a�ݼͼw�üû��j7ü0�˼�Hۼ������%��  �  x�E���j�Y܊�h���yp��#m˽6ؽGܽ��ֽ1Wɽ(P��	���KH��f'���� ,���풽��L׺�o�̽��ؽ�۽D�ս��ǽ裳�+̜������a�x.>���!�-�������K���Ҽ�.˼��ɼ3�μ��ټ)�켼�|"���0� Q��qx��x�������J���sнqaڽQ۽�ӽFlýS[������b���耽Ad���툽�ܘ����	U��l�ѽU�ڽ��ڽe�ѽNt��?)����� }��U���3�ߑ����K)���ۼ%gϼ��ɼ��ʼ��Ѽ�8߼B�����	������:��]�.g��1���*���Ž�Խ��۽�ٽu�ν����^���ϔ��J���]�#C�������J�������gǽ9�սX�۽�ؽ+ͽW���Æ��]��'o�NAI��O*�
X�� �j��Ŷּ��̼V�ɼ�5̼sHռ�t弳�����qO'�vE�s�j��֊��k��ig˽ؽ�
ܽF�ֽOɽLG������C>�� �����!��7㒽+���ͺ���̽�ؽ	�۽�ս�ǽ����ǜ��ۅ�z�a�&>���!����z���]6�ȱҼ\˼üɼ�μ6�ټ���0�[�m�0�9Q�sgx��s��n����F��spн�^ڽ�N۽�ӽ�jý~Z��b���0b���逽se��b�ޘ����BX��$�ѽ��ڽQ�ڽ��ѽ�y��Q/��c
���-}��,U���3�Z��c��-I�Σۼ��ϼ�ʼ�ʼ�ѼS߼���,�	�����:��]�<l��S6��^0����Ž��Խw�۽+�ٽk�νJ���h��|ڔ��U��&s��M������-T������oǽ��ս:�۽x�ؽ1ͽ!Ǻ�����c���3o��NI��]*�\g�K� �l����ּ�ͼ�ɼ"Y̼�jռw�弁���	#��\'��  �  8uG�rTf��Ʉ�8����Ʃ�h���.ý�ƽ�<��Me��#פ��В�e낽�p��fj��6t�����Ö�Oƨ�A�����½W#ƽ������5䥽�_�������	_�GGA���(�	����+��n@伣�ۼ(ڼT�߼3�Q �6��;b�8�5��,Q�V�q�J���̝�+Q���&����Ľ�SŽ�����<���˞����)L}�g�l���k���z��@���Ĝ�\j��)���}�ĽahŽ�V������ӟ�����xu��}T�>r8�Ə!�pg�?V�F��p�B'ڼ��ڼ�⼂��'��c>&��A>�As[�f}�>A���⣽�s�������Ž��ý����੪�;�������Z)v�A�j�Z o�hd��7א�"Ϣ����y4��l�Ž�ý.���u���գ���҆��j���J�H0��	�fN
�����_�輼�ݼ7�ټL�ܼ缔���9��{��*�-��hG��Hf�)Ą�ǌ��S������v(ýQƽa5��V]��~Τ�Mǒ��Ⴝ��p�]Rj�v"t����8���M���򀸽&�½�ƽ }������ߥ�@[��}����_�	?A���(���������)�zۼ��ټ)g߼��6 �_���U�e�5��!Q���q������ǝ�WM���#����Ľ�QŽ��*;��˞�2���L}���l��k�>�z��B���ǜ��m��綼���ĽmŽ\��z���ٟ�;����u�%�T�|�8��!�~w�vf������^Fڼ�ۼ���L�34�""�?I&��K>�*}[��o}�UF��%製�y��e���� ƽy�ý���1���Ę��ć�)>v��j��4o�Dn�������ע�5����;��J�Ž{�ý<���[���©���؆��j�[�J��V0���0_
������輛�ݼ�ټ��ܼR2�6�����?�Һ-��  �  ��O�*Bg�Nq���ʍ�׌��� ���«�j���f>������>��.N��Mh���V��Q�u�Y�F�m�M���}��������ϩ�G=��̶�����Kח��ӊ�F{���a�GK���6��%����?	�<M�����
��s}���f�p�����H�.���A��aW���o�ބ�x+���d���ا� Ϭ����_��_����9���y��8a���S�<�R�Q_�Cv�2����7��dI�������������엟�M���7T���Wr�n�Y�+�C�8�0�������m�s���0��F��[�������#�@#�ڻ4���H��%_��x��R��Ho��K����8��*u��e���B��2���@p��M[���Q��xU���e�YU���������fT�����)�����؛�I>���䁽,�i��PR��C=��*�ċ�����M����,����KZ�Z��4����(��;���O�6g��k��Gō�X���B��߼������K7�����`6��@E��@:h�"�V�A|Q���Y�*{m�(����{������_ȩ��6��2����	���җ�xϊ�� {���a�;K��6�y%������\5���}�����b��Y���f����.�[�A�VW���o�%ل�'���`���է�6̬����^������9��y��8a��S���R��!_��v�񍉽);��)M�����v���������������Z��fr�U�Y��D�E�0���a-�F~����������U���*���0��K#���4��H�c/_�j$x�iW��vt��������m?���|������.���;���Tp��a[��Q�S�U���e��g�)��������[���ì��/�����ޛ�eD��끽�j�M_R�vS=�m�*�J��1���`��?��fS�C���l�њ�����(��#;��  �  �>b�d�q�7w��-���?K���K��k���鏔�Uf������Tjv��x^���I��;�Ɣ7��>��M�ׯc���{�ʈ��䐽	)���r���^�����+��d�}�Zn��^��N���=�g]-��W����y��'
����#���h&�nr6�D(G�Q�W�Mtg�t�v��킽I��j+��m�������E���̌�$�jSn���V���C�P9�!�8�}KB�l�T���k�����<׋����⥕�ӷ��绐�����<����|x�? i��QY�~�H�z:8�V(�j�����P
���
��l������+���;�~�L���\�(�l���{�Z���7��ؑ�<<���[��f���JӉ��B~��Cf���O�-F?�X�7���:�F�G���[���s� Z�����})��/���(����뎽���{E���ns���c�R�S�gfC�`�2��#�9���(���	�M��ɹ�%j!���0��A��!R�1b���q�iq�������E��F��{�������n_��9���<Zv��g^���I�e�;��7���=���M���c�]�{���7ސ�#���m��2Z���댽H'���}��Rn��^��~N���=�S-��L��x��l��
�ɫ����Z&��d6�G���W�~hg���v��肽���e'���i������}C���ʌ������Qn�"�V�;�C��9���8��NB��T�+�k�ݳ��ۋ�f�������-�������Ǌ�����x�y/i��aY��I�LK8�Y(�i��ɔ��`
�b
�k{�S��l�+�s<�<�L���\���l�'�{�(_���<��aݑ�B��ab������'ۉ��S~��Uf���O�QY?���7���:���G�I�[�>�s��a��e���N0���ĕ�g���,�f���L���|s� d��T��wC���2�#��"=���	������`|!���0���A��0R��  �  G(��?��䓆�e���[���q|��e��Z��x6s�3�b���O���<���,��8"��\�#�� 0�]A��?T��f��\v�{���侄��ӆ�H����s��G/�������}�Ŷp���_���L���9�l�*�R"!�VW�\�%�ی2��)D�oW�W�i�<�x�F���0���������!P��mօ�%߂���{��n��\�xsI�b7�(�S? ����%9'��45��LG���Z��Jl�c�z�.j��A���/0��+���� ���o���-���y��\k��{Y�x5F��C4�/�&�N���z �")� 8�րJ���]�4�n���|���:��Z��,�����F���x����w�F�h��SV��C��1�|�$�A,�}i!��<+�@�:���M��`�؂q��~�����D��#x��$���R���!���󮀽o�u�D�e��S�%�?�/�$m#�@��n�"���-���=�\�P���c��s�T!���8����������ш���v�������)s���b�(�O�`�<�{�,�"'"�O���#���/�'�@��0T�P�f�%Pv�������Qφ�����qp���+��|��Z�}�_�p�Y�_�(�L��9�Ѕ*��!�AI��t%�<~2�D��`W���i�5�x�*���q*�����S����K���҅�܂���{��n�&�\��qI��7�J(��@ �A���<'�95�\RG�4�Z��Rl�$�z�o������!6�������'���v��v5��c�y�ymk��Y��FF�NU4�m�&���� �>1)�*8�čJ���]�� o�[�|��������A_��ʬ����������~��"�w��h��cV��!C�Ҳ1���$��>��{!��N+�J�:���M�X�`�7�q�y�~�����K���~������7���~���඀��u���e�I.S�a@��./�K�#�_�-�"���-���=�?Q�|�c�:t��  �  ;���c������F���[�������p�y]a��FQ��@�k0�� ��5�pH���	�	������#���3�gdD���T���d��Tt�Դ���爽GB��瓽�ƕ�����&��Ȅ�.br��Z��F�#G:���7�8
@��Q���g����`]��_���Pw���"��˖��Jދ�����{���k��	\���K�2;�Ұ*���f��F�
�{
����d��|�(�m-9��I��:Z�\ j�]Vy�� ��������vڔ�s���}q���V��S���@j��JS��xA��>8��n9��D�X�o�o�L���N@��
��������@��Tݏ�æ��W���s�u���f��V�Q2F��|5���%����E��
�]�� �v��5.���>�fO��_��*o��b~�D����B����������* ������.5���Sz�$Kb�ݖL�!P=��r7�s(<��J��_���w���������ӡ���������wU��'��/�p�XQa�	:Q��@��0�O� �b%��7�+�	���������#�l�3��WD�+�T���d��Kt����L䈽?���㓽�Õ�o����"��SÄ��Wr�=�Z��F�;9:���7�3�?���P���g���EV���ّ��p�����u���~ً�����l{���k�n\���K�8
;��*��������
�w}
�����(�49���I��CZ�L
j�bay��&��%���
��┽m����y���_��4���Rj��\S���A��O8�S9���D��*X���o�6����E��Շ��3ƕ�(E��}ᏽ��������v��f�ĶV�=@F���5��%����+W�c
�ļ�	���UE.�{�>�HtO���_��7o��o~�Б��zI��ޝ��_���x�������>���gz�d`b�¬L�Uf=�
�7�0><��J��_�H�w�����ʏ��  �  P��m�������ᙽ����j���e�o�N��:�/�'��$���
��� ������[�=�����l��4r���+�l>���S�pdk�B�������w���ی���]��c���z⦽����#�����}�͡d���T��Q��B\�ѻq�C���畽Ȕ���ɪ�n6�������`��н������?�v�:�]��{G��3�3]"�e��.��������6�h���!���� ���1�"E��1[���s�����L���/�������NR��b����n��̰��ݑt� ^��kR���S��Ib��z�~���z��L⥽6A��$���:l���ĝ��p�����3&n�EV��@�7�-������������ e������ ��	�{��%���7�%4L��#c�r|�
����P���	���=-��li��,����䵃�ul���X��iQ�/^W�9~i����w������n���������蚤�(ܙ� ���_�K�e���N�Z:���'�`��
�� ����6<�������1��e��+��a>���S�~\k�ͣ�����������Z��ؙ��cަ�/񛽺���_�}�t�d���T���Q�3\��q�t���ߕ�o����ª��/������?[��ḕ�b�����v���]��vG��3�(Z"�c�.� ���7���
o�������g� ���1� +E��;[��s���pS���6���������Z��B����w�����X�t�;(^�F}R���S��Yb���z�!��π���祽�E��h���:p��sȝ�	u��#���/n��!V��@�R�-��$������������3���� ���	�m���&��7��AL��0c�3|�����������5���r��3������ ���Y5l�*�X�ӀQ��tW��i���,���Þ������  �  ?(ƽX�½ya��iѨ�����Ã�o|d���E��r,�����������m�{�ܼ^�ټ�޼��鼧W��z0�m&���1�(AL�5�k�)���G�������7��.2Ľ��Ž�����ಽ-ա��鏽������n���j�Nw�Z���������x����ĽW�Ž������`䢽n6��l{�=�Y���<�k%�+��t����#?���ڼ�]ڼ���
��Q�K�"�b�9�e5V�ow�����נ��뱽�羽�Ž��ĽK��Mz��ٽ���V��.�y�:sk�hBm�\�~� ���˟����f���.�Ž��Ľ񄼽oj��.Ü��q�o�
O�Q4�B��������A8��޼'�ټq�ۼ��伳+��o_����)�0�B���`������f���٦�#ֶ�����#ƽ��½Ǽ���§�����;��-s�y<j�=jq���������p˥�c+������� ƽu�½/[���˨�|���l���Aqd�
�E��f,����)���o���O�Inܼ'�ټ�޼ ���<��$�M��1��8L���k�݇�w���ޕ��c4��2/Ľ��Ž�����۲��ϡ��㏽����>vn�N�j�>w�@���ﺙ����謺��Ľ��Ž����睳�Sߢ��1��Xd{���Y���<�/%�d(��r����?�h�ڼdbڼ�%��n��X�3�"�k�9��?V�]zw�����ޠ�󱽡ﾽa�Žc�Ľ[������KǛ�`��֗y�V�k��Sm���~�u��Sҟ��#������чŽ��Ľǈ��(n���Ɯ���l�o��O�C\4�kN�f�������V뼼߼W�ټ��ۼ{�伳J��kn�v���)���B���`�/���~m���ঽ�ݶ�=���,ƽ��½1Ƿ��ͧ��ŕ�hG��Es�xTj�q�װ���˓�xե��4������  �  �ܽ�׽ȃʽGA��⭠�6���=nh��C���%��K[���y�%�ԼR̼*�ɼWeͼ"�׼p	�3w�ю���+��:K�\|q�Ʀ��:ԥ��컽�	ν�Tٽ��۽�սtƽ�ٲ�j8������2遽A�����ԕ������#���iϽ��ٽ.�۽�
Խ��Ľ_�D蘽a1���d[�D�8����K���S�fN޼B Ѽyʼ�!ʼ'�ϼrܼM�������z5� /W�ׄ�uM��yj����½��ҽ�)۽{�ڽJ�н�A���׫�З�8��Y(��{1��z ��������foĽ��ӽҁ۽�ڽ)�Ͻ|-��J`��#0��ev�)O���.�'��W'�Q]��
ټ�μJ�ɼ�W˼,OӼ�;⼂$��!����"���?���c�(�����QԴ�ÚȽ8sֽ�ܽTHؽ�̽�����ꤽ�����
�~�⒃�Z��餢��j��8;ʽP׽5ܽ�׽j}ʽa;��G�������-ch���C���%�m���@��^�t�Լ,�˼�ɼ�Hͼ�{׼���nk�F��u�+��2K��uq�ݣ���ѥ�껽ν�Qٽ��۽�սRoƽQԲ�!2�������ၽb���醽}̕�q������#bϽ?�ٽT�۽mԽĝĽ:믽�㘽s-��H^[���8�d}�$���O�L޼� Ѽ�{ʼ�&ʼ(�ϼ7{ܼ���l����܃5�@9W�A���S��Uq���½�ҽ�1۽W�ڽ�нK��"᫽�ٗ��A���1��C:���(��c��߈��euĽ��ӽf�۽�ڽޭϽ1���c��4���v��'O��/���Z4�Ly�S(ټx3μ��ɼ9w˼/nӼ�Y��A��]���#��?��d�������۴���Ƚ�{ֽ�ܽQRؽf̽����m������������������*��揤�t���Dʽ�X׽�  �  �$�彌;׽�����V���{���m�4D��r#���
�Y/�G2ڼa	˼��¼>���"/ļ��ͼ&�޼�������j*�ӜL��;w�G"�����O�ƽv/۽h����꽏��:�ӽ�K���ʧ���l��������u��*����'��E�ʽ�uݽ�轴}�b���н�q��֠��N/��J�^�^T8�$R�����S/Լ��Ǽ:{��+����ƼscҼO.����u���4�9�Y��v��"�������UEν^�z��4��X߽��̽x���UР��؏�����7����Hf��۽���}ѽ58�k��5��wݽ\gɽ����`���tb|���P��h-�D�=x��m�!ϼC�ļ����EH¼%�ɼ! ؼ���7h��C �Q@�&h����1j��x��ս;�佫 �罔�ٽ[�ŽN���l���勽W��F͊�.q��
���JHý��׽�
�C���!5׽����Q��v���m��(D��f#���
�/� ڼI�ʼD�¼գ��Zļ�ͼ:�޼����W����)�:�L�E5w��������ƽ -۽��罂�꽓��x�ӽfF��}ħ�ջ������ȸ���m������I���ʽ nݽ����v����M�н�l��@���V+����^��N8��M������}-Լa�Ǽ�}���/����Ƽ�lҼ�9漼��}�ė4���Y��|��v��������Lνf���&�齥&߽#�̽0���ڠ��⏽>!��z@��i
���m���Ļ��ѽq=����4��ݽ�jɽ{�������j|���P�Xs-��#��������=ϼA�ļG���g¼��ɼؼ��Vv��Q ��'@�w3h�ӱ��8q�������ս��
�G!�z�ٽ��Žc$��y��K򋽢c���ي�}��?����RýI�׽���  �  ~
���Ɔ��{� a���A���!�����ռqխ��v���2x�W�]���M���E��C�� G���P��|b�����&��Lµ��	༑_
���(��H�aog��2������扽����)�w���]�}VB�l�*��d�����,#��"7�:nQ���l�ρ�д��墉�&X��Zps���V�P7�y��3��8#ǼQݢ�������m��W��:J��D��CD��BI�_6U�&�j��M���o��3�¼�c���'b3��dS���p�A_��)Q��$���̂���o�ErT���9�6�$�b�ch�1�(��c?���Z�u�⯄����������P���j�PoL�	K,����U弢׹�����ꁼu�d���Q���G�B�C��?E�?SL�%[��dt�����d���ءм��<D�c(>�ע]���x�V���􉽱�����G�f�=K��1����}���vz/��6H�t�c�)�|������������~{���`�!�A���!�W�q�ռ�����]����w��e]���M�b�E��C���F��OP��Kb����%�������߼�X
���(���H��ig��/�����<㉽]�����w��]�JJB��*��V����+#�]7��^Q���l��ǁ�쭈�s���2R���es���V���6��q��&���Ǽ(բ�������m�*W��;J�8�D�OMD�UPI�!HU�$�j�[���~����¼Kw� �#n3��qS���p��f��$Y������Ղ���o�o�T���9�7�$���/y��(�hr?��Z� u�C���˸������T��͏j�%wL�;S,�Ŗ�6i��칼�+����$e�R���G��D��{E��L��_[�@�t�ˍ����ݼмn��Q�}6>���]�@�x��
������h���r4��f��SK�M2�� ��)�)����/�'LH�`�c���|�S���  �  ᆽ���#v�Ӊ\��o>�c�����ռ�r���ܑ�F�{��'a�g�P���H�òF��J�V�S��f�����j���"���߼����O&��OE�þb���z�$����"���:r�{�X��N>�~�'�Yd�3��f���i3�n�L�N�g�p�}�����~��7g��rRn���R��4�|���v����Ƽ�ʣ�B���_q���Z�(NM�$NG� G��JL�p�X��:n��臼�t���}¼���jX�U�0�riO�}k�'w��50������Ψ�m;j�v�O���5��!���(n� q%�tp;�i�U��o���������n����|��e�S�H�в)�y�F+����D��𗃼"�h��+U��J�<�F��H��}O�̪^���w�
$��󰪼'мY���+���:��JY�q�s����ĕ�2���_y���a��F��U.�b��M(�ߍ���+�QD���^�+w��能Fن����v��}\�d>��������Լ�Z���Ñ�<{���`�L�P��H�U{F�S�I�4�S�p�e�B���sU��J��\�޼����I&��IE��b���z��q����z���0r���X��B>�0�'�V�C��
��Z3�
�L�Fxg���}�9���`x��Ia���Gn�C�R�e 4����i��C�Ƽ�£�<���Wq�d�Z�OM�BSG�c	G�+XL�/�X��Pn����� ���C�¼d��Jc�K�0�xvO�'�k��~��+8�����)��BMj���O��	6��!�0#��~�Ȁ%�;���U��o����Տ��Ms�� }���e�9�H��)�`��>�,��\��;����h��dU���J�"�F��IH���O���^�U'x�+@��n̪�&BмG����8���:�vYY��s�	
��jՆ�ݏ���sy�y�a��G��l.�����?�Ϥ�,�nD���^��#w�B��  �  ��{��v��g��;P�U5���� ��HԼ�3��M���������l�g[�;2R��O��S��|^�0�q�J���훼�:���Mݼ������z;�b�U��Ck�^�x���{��s���b��]K��2�������5W�L��b�(�JW@�!�X�m��zy��]{��`r��`��G��,�{��;��<�Ǽ%g��܉����|�G�e��XW�OP�I$P��6V���c���y�2L���Q��^vü&��)����(�<D���]���p��z�+z�t�n�73[�]C�<++��p���g������40�T�H�/%`�g@r�'O{�X�y��-m�"qX���>���"�pB�X��"ӻ�/����'���t�o�_��<T�آO��_Q��Y�j�i����(��Z���C�ϼ�����k12�TM�X�d��8u�<�{���w��i�~mS�B�:�$$�0�������X�!�!8���P���f�9ev���{�|v��
g��/P��I5����= �~1ԼK������{���Wl��.[�p�Q���O�rhS�@G^��fq��2��K؛��'���<ݼU|�)���s;�z�U�w=k�ңx�A�{��s��b�SK���2�T��t��qH� ���(�H@�I�X��m�omy��P{��Tr��`�s{G� ,�������|Ǽ_��󃏼�|���e��YW�q�P��-P�DV�M�c���y�DY���`����ü��������(�-�D���]���p���z��;z���n��D[�MC�6=+����;����d�C0���H�01`�-Kr��X{�*�y�6m�"yX���>�H�"��K�Q��黼����A���Mt�D/`��xT���O�ޜQ��Z�8j�؁�E���ڭ�V�ϼ�������a?2��bM���d�:Iu��{���w��-i�؂S�|�:��:$�I$�������3
"��-8��P�g��uv��  �  S	b�^�˟Q��?��1)���Z>��w�ּ黸����;Ŏ��	���o�#%d�'a��e���r������l���ӥ�nԾ��F޼f�.���2.�ŖC�M�T��_�V�a�'oZ�(FK��7�}�!�rp��X���U	����~t-���B�A�T�4�_�˰a��Z��K���7�D�!�Da�O�˼���FX��Y���~�z��Sj�4b�ʬa���h��ax�����7���^���rȼ��I�����5���I�xYY��Ja�4.`��V���D���/����Ц
� ��9����_d�
�4��+I��Y�Ea�4P`���V�ǾE���0����W�	⼦����7���;��|	��J;t��f�a�?0c�|+m�VP��ꌼ���q�����ҼT���1-���&�Ӷ<���O���\�]�a�R�]��Q�>�̟(����@��`c���5���D&��;��&O�w�\�F�a�=�]���Q��	?�&)����O'����ּ4�������+����퀼��n���c���`���e�%Tr�d���6T������~����4޼��*��8,.���C��T�M�_��a��fZ��<K��7���!�yc�*������F	�����e-���B�={T��~_�S�a���Z���K�<�7��!�Z��B�˼���qR������H�z��Tj�[!b��a�:i�:sx�����D���m����ȼ
-�	�W�ؓ5�`�I�5hY�'Za��>`��%V�3�D�h�/���P�
�1��I�*���r�9�4��7I�lY��Na�*Y`��V��E��0�Q�a��/�f ¼�P���V���%���vt���f��La��nc��im�,��!���Ȟ�=ϵ��Ӽ&����:�m�&�3�<�2�O��]��b���]��Q��'>�{�(��������y�)����8Y&�B�;��8O���\��  �  �DD�u`B�� :��=-������w���	���ȼĵ��j���kk�����:����|�V��H<��%|���R���$��l�ͼ���̪��C�"X!��d0�:l<�aC��C���<�m�/���PL��[��j�N�开>����	���(�I�7�t�A�eD��=@��96��@(��g�.q��󼳁ؼ�Z���B���������.����}�$M}��X���Ì�/K���*���ڶռ���R��s��I�&�4�4�U?��5D�T'B�o9��*����u��h���C�G�v}���`�j��.'.�y�;��DC���C��s=���1�2#����N���Qgм=P��+��4����F���ہ�T|�HG�����}֐������o���-ƼF޼�d��K��M��e�+��8���A��XD���?���4���$�!�ê�T�P
�6F�Y�����"�s43���>��5D��RB�A:��1-����,��(�����༞�ȼ,����j��UN����������R|� 8��D���`���8����>�ͼ���i��I<�;Q!�,^0��e<�(ZC���C�U�<���/����@��B���N�
��!�A�(��~�(���7�x~A�SYD��2@�a/6�m7(�_�j�{�wؼS���<����:��/���}�uV}��_���̌�V��t7��������ռ��������&���4��c?�ED�d7B�09�,�*�����[���
e�f7�ۛ��o�w�3.�I�;�eNC���C��|=�]�1��#����X����+м1j���F������e��y���	�|���������������򌱼JƼ,޼|�������y�+���8�M�A��iD���?�!�4���$��Q���6��5��p�+�D&�'�"��E3��?��  �  �+'�U9(�O%����o�������4���ϓ��Ѽ¤��򳫼=������e�����a��iw�����)wռ���:�������;���u ��&��_(��F&�]��0�._��u�k�ؼ�ɼ��Ƽ��м��~����?�b����#��(���'�F#��Y�p�������:2�޼	{ʼgS���P��o���T���񑼻R��F���D���Dȼ��ۼ��� �3
�9��~m�d�"��5'��"(�p$����k��׀����pQҼd5Ǽ3�ȼWQּDf���7��uF�g�%�_W(�	~&��-!�������{�����Y�׼��ü�H���n��[R��le���N��*͛�#é��k����μT��S�������`��]��x$��(��v'�Y%"�rB���s���ݣ߼hRͼ^?Ƽy�˼�&ݼ�m��ف	����B!�T'�,(��%�����������i���y�e�мՇ�����������E���t���IZ������%^ռ@�����������о��n ��&�^X(�?&��T�~'��T��^�ؼ��ɼ>�Ƽ��м���T����1���&�#���'���'�<#��P�m������v(��	޼kuʼ�O��fO���o��XW��@���nY������N���Qȼ��ۼ�（� ��
����y�Ȝ"�D'��1(��$�:� ��Ǒ�����rҼVǼ��ȼ'oּ*������MQ�d�%��`(��&��6!�ʲ�?�6����=�꼨�׼4ļ�g�� ����s�����Qp��%4㩼����.�μrp�2o����������7�$� (�ֆ'��6"��T�7)�Ұ��T�߼f|ͼFiƼ�̼�Nݼ���֓	����,R!��  �  �m��>����,��#����������������㼒ͼ ������ʩ�񓯼�ƽ���Ѽ��ԝ������d�����G�>��!���[��6��R��U�߼��ɼ�Z���2�����a������ЎռQg��� �H�	��E�X�P���C����<������F��!��=�ۼ�Ƽ�ᴼ��������_��9�ü�=ټ��ђ�����g��X���:������_��T�
�������׼y�¼>����O���a�������'ǼDݼ���P(��=�����;�����=��j��&����?d	��b ���:Լ����٣���թ�-}�����ʼ��༴p��X���V������e�o-�($�L��S�h��V��':缞�м<����ޮ�E����ԭ�pź��μͬ�0�����_��1�Q��O �:�=�����
����Z����h��̼\߹�x^��9����r��9���$�Ѽ��*������Z���/?�6�����~�kT�"��e-��?����߼�pɼ�B��K�������E��^����sռ�L�� ��	��:�eM��y��:���m���:����������ۼ�Ƽ<ⴼq"��,���Ff����üBHټN#�1��,�7�������%G�B���������
���~�ؼ��¼񻲼�o��R�������7CǼ� ݼ��/3�H�"���D�(��2G��t��1�� ��q	�`q ��-뼛ZԼqƿ��ư��������.<���ʼ7��������Zd�@����r��:�2� �����-z��W_�M�м�ϼ����v���h����뺼@Cμz�伛"���,��  �  ����Z��ǘ�u`��K�,Y%�MH(���&�}� �mN����Y��dܼtq˼�vƼ�9μ
�p?�����o��C�"�H�'���'�:$�����w���u��^���W�2�ͼ�x�������E��^��g����ᖼ�K���Y��nż��ؼ���ǳ��&�����!��!��&�zT(��o%�{����������Tռ�Hȼ��ǼASӼ|�PT��|�Η�	�$��6(�x'�9"�&��}��~	��R ���!�ڼ$Ǽ�6���£�����v����������� ��"P��6�˼߼!7�sg�ڋ�(x�5���#���'���'�y`#�1�o��D��Đ�D�ϼ~�Ƽ� ʼ��ټi��/����Z��5z&�P(���%� 	 ��D���z�#���1��AԼ���b`��e0�����V9���F��ȝ�#������|Ҽ/��|q���u�Ɍ��T�(@�M%�'<(���&��� ��?�$������B�ۼyN˼XSƼ�μ������o��D��\�"���'�}�'��0$�x���o����m��N��"F�O�ͼd���ᨼ�-������}���ǖ�1��9?����ļ��ؼ��{����~�%����F�!�K�&��N(�k%�˺�K������뼨Tռ�Kȼd�Ǽ�YӼ"#鼣Y������T�$�@(��'�=D"�7�����	�>a �8�H�ڼ�CǼ�V��㣼�ߗ��ڑ����)���;��Ui����˼�3߼�K�>q�x����Z��ĝ#�E�'�v�'�vn#�3@�J�g��F�㼑�ϼ�Ƽ�Dʼ��ټ{��o/���������&�R](���%�� ��Q�[��F��0���%���bԼ����j���pV��-.���_���l���일k���b����1ҼP���  �  �|�`��<����5.�ù:���B��)D�?�>�bu2��!�{-��e ����YG��(�=����{�%��5�e@�3qD��gA��>8�9�*�s�������$�ܼ�ż0u�����
8��a�����B�|�K�������ܗ�':��m���x�Ѽ�]�2+����.�#�N�2�1�=��C��
C�O;��H-�S �D{
�A8����缇��Ь��������v+�%�9��yB�)!D���>��4��%�u�����QUԼu���{��Kg��b���肼��|��~�֑��F���d✼�D����¼ �ټr����K	��I�6)�6�6���@�}eD��#A��
7�U�'�X���'�Q�Ho弬��B���1������0�~m=���C��C���;��/��k ��T�� ��P弌{̼趼�<��˒��芈�怼�=|��X���v���
��W�����w�ɼ�b�@G��p�������-��:�b�B�sD�0{>�Kf2���!�v��S �fy�{"� �]}���V�%��5�pW@��dD��\A�58�.�*���
�������ܼ>�ļZb������Q"��N}��$�~��|�k1��;܊�R×�!!��Dm��p�ѼMH�!������#�ڝ2���=���C�4C��;�/F-�����z
��8��F��,��q���?�����|+�e�9�6�B�T*D� �>�4�Ȱ%�-����xm�(sԼ�׽��;��ц���3�����5}��S~���֎�U���\��ޜ¼��ټs����U	��S��)���6��@��rD��2A��7�D�'�.�:�2�2��$꼼����B�^ ���0�4|=���C��*C�L�;�k�/�Mx ��a��� ��m�<�̼����^��Q���h������ԇ|�}��b����,��<w��Gϴ��
ʼ�  �  גؼ�t�����?s*��:@�R��v^���a��B\�CN��:�-%�g�V�����x�"���)�sN?���Q�wP^�� b�z\�5�N���;��i%��������;Ѽ�Y��Ť���'��JE~�r�l��c�gWa��[g�wcu�#ׅ��F��⊩���ü�伏��aT���1���F�HHW��`�]a�G`X��"H�'p3��M�A������b�~i��;1���E���V���`��a�B�X�S�H��O4�������
輛�Ƽ>��w(��q8���8w�xIh��ga��Db�Y�j��{�i��3a���v���ͼ�a𼩏���"��,9�~�L�3H[���a�u_�j�S���A�E4,�_�����ϟ�\�A?�?�"��28��;L��[��a�@_�-#T��pB��,��R��� �BܼS,�� ���D_��邼�^q�j$e���`��Gd���o�b���ʋ�������yؼu\��9���g*�4/@�PsR�Zj^�1�a�B4\��3N�`�:�x%��6C�wq��e����?�)��=?���Q�)B^�	�a�un\���N��;��`%�)��_����*Ѽ5H���������~~�/il���b�u&a�*g�F1u�>����.��Ws��|ü�
伶x�UK���1���F��AW���`��
a��\X�* H��n3�GM������e��l�f�
1���E�*�V�%�`��!a�B�X�6�H��[4�1��h��&輥�Ƽ1"��G��\W��Yvw���h�M�a��~b��%k�`�{�Ɂ��sx�������ͼ�u�ϙ�)�"��79�C�L�U[���a��-_��S��A��F,������_��[o��Q�/�"��C8��KL��[���a�1M_��/T��|B�z�,��_��� �^ܼ�I��S���/���\���q��ke�D"a��d��o�F������{;��o;���  �  m�ּ�n��:���6�U�Q�<,h��w��{��u���e�?yO��6�~� ��Z����^���Y%�?<���T�53j� x��{���t���c���K�N�0��@�_G����ͼl2��O��
���+	i�!LY��IQ�k�O���T�y�`���u�[:��}	�����P���	�ZU$��@���Y��n���y�{��xq��^��6G�P�.�����?���N�)o,��pD�){\�[�o�Y�z��z���o�PR\�� C��\'�~v��	�.z��Ϣ�?1��'Fx�A�b�КU��O��P��W���f��~~�\�����ʋɼH�"F�ӏ-�;�H��Ma��s���{��y�Fl�SaW�'�>�֔'���E�?�#���4�׮L��c�0tt�b�{��#x��7j��_T���9��5�Y�F�ڼ�T��m|���8��p�9n]���R��xO��DR���[���m��^���◼	Ѳ�.gּ�b�p/�|�6��Q�e h�w���{�j�u���e�PhO���6��� �G�M��ɷ��F%��,<���T�	#j�Ix���{���t��c�)�K�;�0�8�s6��^�ͼ� ������值��h��Y�CQ�a�O���T�J�`��nu�z"��h����I;�K�	�uL$���?���Y��n�r�y��{�uq���^�`5G���.�;�l������Q�os,�vD�]�\���o�r�z��z���o�]\�|C��h'����O%�ז���좼eO���x�*�b��U�l#P���P��X���f��~���������ɼ�%�wP�x�-�xI��Ya�*s��{�^y�7.l�esW�'�>�~�'��2�M3��R�B��	-4��L�7�c�+�t�T�{��0x�Dj��kT��9��A�@&�wۼ�q��ߚ���X���Pp���]��@S� �O�o�R�b&\��m��|��g����벼�  �  a�׼Ml��<!�H)@�*^�Yw���y߆�I����u��s]��B��*���2M���O�/�цH��Ic�?�z�`ׄ�!ǆ������Xr���W��>9��������ͼ����E����bv�@�]�O�X H���F��K��%V��j�ѳ���ԛ��1����漙���k+��gJ��6g�:~�����n���<��]Rn��vT��:�Vz$�%��b�	�"�
W7�<rQ�2�k��Q��* �� ��n���j���M�R�.���r�EO��=Ԟ�v����l��W�o�K�M�F��dG�3�M�`[���r��j��Js��42ɼ�@���:�#�5��jT�x�o��с�S���IR��צ|��f�nK��2�F��r������(���?�VkZ�5os��ۂ�xǆ�{���q�y�u-a��C�ߒ$�$g��jܼ���pᕼ������d�#�R�#rI�lF�H�H��iQ��b��P}�z��"9��oj׼y`�?1!�	@��^�7Mw�����؆�铃�"�u��b]���B���*����39�'��ɐ/�	tH�8c��z��τ�H��������Mr���W��59�P��y�����ͼ�쨼�⍼);v�;�]���N�G�G��F�V�J� �U���i�=���ڽ����6��	���b+��_J��/g���}�奅��k��2;���On�HuT�N:��z$�}�'e�T�"�M[7�wwQ�b�k�OU��3$���������j�)�M���.����5켰k����V߆�_�l�r�W��K��G�Z�G�w�M�	�[��s����N���cGɼ�U��LE���5�FvT�ȳo�:؁�����FZ���|�$f�_�K��%2��2��������(��?��|Z�os�'ソtΆ����ڱy��9a��C��$��s�K�ܼ�-��V��������d�ZS�X�I�İF��I�s�Q��Xb��}��6���S���  �  E=ؼܧ��#���C�7�b���|����G	��毆��{��`b��F��`.����7��� ��B3���L�?bh��,���􇽪����|�w��\�i<�������9Hμ�7��y��[�r��?Z�@�K��5E��D�x$H���R�aqf��
���������輑0��.��3N��l�|܁��È�e����?��R�s�� Y�9�=���'����U���%��,;�-V���p��M���F��L'��:₽,
o�T�Q���1��l�ό�C���Ý��!���i�%>T�t�H��D��D�;�J��X��To��ቼ9����pɼZ���%���8��X�-�t��Ƅ�����ds��=@��a?k���O���5��G"��^����,���C��A_�ey��ꅽi�q���y/���e��G���&�����Pݼ��������د}���`�l�O���F���C���E��-N��^���y�ȼ������l$ؼ���y#�V�C�Җb���|����v�������{�vOb���F�]M.�����#�ŷ ��.3���L�^Ph�w$��S퇽�牽����X�w���[��_<���b���6μ�%��Of����r��Z�1�K�
E���C�X�G�<�R�mAf�]�헚�m�V�
'�(.��+N��
l�^ف�����1���+>��̻s�mY���=���'��	��W��%��0;�fV��p�\Q���J���+��(炽�o�ܴQ�I�1��y����_��᝼�?���Oi�JzT���H��JD�n�D�\�J��8X�{�o�����@���0�ɼ0,��0���8���X���t�Ÿ́�É�m{���H���Qk�.�O���5�\"�Is�����,�%�C�\S_��y�l�g��������;���e��&G� '�M��kݼ��������G�}��<a�9�O�L�F���C��<F��nN���^�Zz��ؑ�ů��  �  a�׼Ml��<!�H)@�*^�Yw���y߆�I����u��s]��B��*���2M���O�/�цH��Ic�?�z�`ׄ�!ǆ������Xr���W��>9��������ͼ����E����bv�@�]�O�X H���F��K��%V��j�ѳ���ԛ��1����漙���k+��gJ��6g�:~�����n���<��]Rn��vT��:�Vz$�%��b�	�"�
W7�<rQ�2�k��Q��* �� ��n���j���M�R�.���r�EO��=Ԟ�v����l��W�o�K�M�F��dG�3�M�`[���r��j��Js��42ɼ�@���:�#�5��jT�x�o��с�S���IR��צ|��f�nK��2�F��r������(���?�VkZ�5os��ۂ�xǆ�{���q�y�u-a��C�ߒ$�$g��jܼ���pᕼ������d�#�R�#rI�lF�H�H��iQ��b��P}�z��"9��oj׼y`�?1!�	@��^�7Mw�����؆�铃�"�u��b]���B���*����39�'��ɐ/�	tH�8c��z��τ�H��������Mr���W��59�P��y�����ͼ�쨼�⍼);v�;�]���N�G�G��F�V�J� �U���i�=���ڽ����6��	���b+��_J��/g���}�奅��k��2;���On�HuT�N:��z$�}�'e�T�"�M[7�wwQ�b�k�OU��3$���������j�)�M���.����5켰k����V߆�_�l�r�W��K��G�Z�G�w�M�	�[��s����N���cGɼ�U��LE���5�FvT�ȳo�:؁�����FZ���|�$f�_�K��%2��2��������(��?��|Z�os�'ソtΆ����ڱy��9a��C��$��s�K�ܼ�-��V��������d�ZS�X�I�İF��I�s�Q��Xb��}��6���S���  �  m�ּ�n��:���6�U�Q�<,h��w��{��u���e�?yO��6�~� ��Z����^���Y%�?<���T�53j� x��{���t���c���K�N�0��@�_G����ͼl2��O��
���+	i�!LY��IQ�k�O���T�y�`���u�[:��}	�����P���	�ZU$��@���Y��n���y�{��xq��^��6G�P�.�����?���N�)o,��pD�){\�[�o�Y�z��z���o�PR\�� C��\'�~v��	�.z��Ϣ�?1��'Fx�A�b�КU��O��P��W���f��~~�\�����ʋɼH�"F�ӏ-�;�H��Ma��s���{��y�Fl�SaW�'�>�֔'���E�?�#���4�׮L��c�0tt�b�{��#x��7j��_T���9��5�Y�F�ڼ�T��m|���8��p�9n]���R��xO��DR���[���m��^���◼	Ѳ�.gּ�b�p/�|�6��Q�e h�w���{�j�u���e�PhO���6��� �G�M��ɷ��F%��,<���T�	#j�Ix���{���t��c�)�K�;�0�8�s6��^�ͼ� ������值��h��Y�CQ�a�O���T�J�`��nu�z"��h����I;�K�	�uL$���?���Y��n�r�y��{�uq���^�`5G���.�;�l������Q�os,�vD�]�\���o�r�z��z���o�]\�|C��h'����O%�ז���좼eO���x�*�b��U�l#P���P��X���f��~���������ɼ�%�wP�x�-�xI��Ya�*s��{�^y�7.l�esW�'�>�~�'��2�M3��R�B��	-4��L�7�c�+�t�T�{��0x�Dj��kT��9��A�@&�wۼ�q��ߚ���X���Pp���]��@S� �O�o�R�b&\��m��|��g����벼�  �  גؼ�t�����?s*��:@�R��v^���a��B\�CN��:�-%�g�V�����x�"���)�sN?���Q�wP^�� b�z\�5�N���;��i%��������;Ѽ�Y��Ť���'��JE~�r�l��c�gWa��[g�wcu�#ׅ��F��⊩���ü�伏��aT���1���F�HHW��`�]a�G`X��"H�'p3��M�A������b�~i��;1���E���V���`��a�B�X�S�H��O4�������
輛�Ƽ>��w(��q8���8w�xIh��ga��Db�Y�j��{�i��3a���v���ͼ�a𼩏���"��,9�~�L�3H[���a�u_�j�S���A�E4,�_�����ϟ�\�A?�?�"��28��;L��[��a�@_�-#T��pB��,��R��� �BܼS,�� ���D_��邼�^q�j$e���`��Gd���o�b���ʋ�������yؼu\��9���g*�4/@�PsR�Zj^�1�a�B4\��3N�`�:�x%��6C�wq��e����?�)��=?���Q�)B^�	�a�un\���N��;��`%�)��_����*Ѽ5H���������~~�/il���b�u&a�*g�F1u�>����.��Ws��|ü�
伶x�UK���1���F��AW���`��
a��\X�* H��n3�GM������e��l�f�
1���E�*�V�%�`��!a�B�X�6�H��[4�1��h��&輥�Ƽ1"��G��\W��Yvw���h�M�a��~b��%k�`�{�Ɂ��sx�������ͼ�u�ϙ�)�"��79�C�L�U[���a��-_��S��A��F,������_��[o��Q�/�"��C8��KL��[���a�1M_��/T��|B�z�,��_��� �^ܼ�I��S���/���\���q��ke�D"a��d��o�F������{;��o;���  �  �|�`��<����5.�ù:���B��)D�?�>�bu2��!�{-��e ����YG��(�=����{�%��5�e@�3qD��gA��>8�9�*�s�������$�ܼ�ż0u�����
8��a�����B�|�K�������ܗ�':��m���x�Ѽ�]�2+����.�#�N�2�1�=��C��
C�O;��H-�S �D{
�A8����缇��Ь��������v+�%�9��yB�)!D���>��4��%�u�����QUԼu���{��Kg��b���肼��|��~�֑��F���d✼�D����¼ �ټr����K	��I�6)�6�6���@�}eD��#A��
7�U�'�X���'�Q�Ho弬��B���1������0�~m=���C��C���;��/��k ��T�� ��P弌{̼趼�<��˒��芈�怼�=|��X���v���
��W�����w�ɼ�b�@G��p�������-��:�b�B�sD�0{>�Kf2���!�v��S �fy�{"� �]}���V�%��5�pW@��dD��\A�58�.�*���
�������ܼ>�ļZb������Q"��N}��$�~��|�k1��;܊�R×�!!��Dm��p�ѼMH�!������#�ڝ2���=���C�4C��;�/F-�����z
��8��F��,��q���?�����|+�e�9�6�B�T*D� �>�4�Ȱ%�-����xm�(sԼ�׽��;��ц���3�����5}��S~���֎�U���\��ޜ¼��ټs����U	��S��)���6��@��rD��2A��7�D�'�.�:�2�2��$꼼����B�^ ���0�4|=���C��*C�L�;�k�/�Mx ��a��� ��m�<�̼����^��Q���h������ԇ|�}��b����,��<w��Gϴ��
ʼ�  �  ����Z��ǘ�u`��K�,Y%�MH(���&�}� �mN����Y��dܼtq˼�vƼ�9μ
�p?�����o��C�"�H�'���'�:$�����w���u��^���W�2�ͼ�x�������E��^��g����ᖼ�K���Y��nż��ؼ���ǳ��&�����!��!��&�zT(��o%�{����������Tռ�Hȼ��ǼASӼ|�PT��|�Η�	�$��6(�x'�9"�&��}��~	��R ���!�ڼ$Ǽ�6���£�����v����������� ��"P��6�˼߼!7�sg�ڋ�(x�5���#���'���'�y`#�1�o��D��Đ�D�ϼ~�Ƽ� ʼ��ټi��/����Z��5z&�P(���%� 	 ��D���z�#���1��AԼ���b`��e0�����V9���F��ȝ�#������|Ҽ/��|q���u�Ɍ��T�(@�M%�'<(���&��� ��?�$������B�ۼyN˼XSƼ�μ������o��D��\�"���'�}�'��0$�x���o����m��N��"F�O�ͼd���ᨼ�-������}���ǖ�1��9?����ļ��ؼ��{����~�%����F�!�K�&��N(�k%�˺�K������뼨Tռ�Kȼd�Ǽ�YӼ"#鼣Y������T�$�@(��'�=D"�7�����	�>a �8�H�ڼ�CǼ�V��㣼�ߗ��ڑ����)���;��Ui����˼�3߼�K�>q�x����Z��ĝ#�E�'�v�'�vn#�3@�J�g��F�㼑�ϼ�Ƽ�Dʼ��ټ{��o/���������&�R](���%�� ��Q�[��F��0���%���bԼ����j���pV��-.���_���l���일k���b����1ҼP���  �  �m��>����,��#����������������㼒ͼ ������ʩ�񓯼�ƽ���Ѽ��ԝ������d�����G�>��!���[��6��R��U�߼��ɼ�Z���2�����a������ЎռQg��� �H�	��E�X�P���C����<������F��!��=�ۼ�Ƽ�ᴼ��������_��9�ü�=ټ��ђ�����g��X���:������_��T�
�������׼y�¼>����O���a�������'ǼDݼ���P(��=�����;�����=��j��&����?d	��b ���:Լ����٣���թ�-}�����ʼ��༴p��X���V������e�o-�($�L��S�h��V��':缞�м<����ޮ�E����ԭ�pź��μͬ�0�����_��1�Q��O �:�=�����
����Z����h��̼\߹�x^��9����r��9���$�Ѽ��*������Z���/?�6�����~�kT�"��e-��?����߼�pɼ�B��K�������E��^����sռ�L�� ��	��:�eM��y��:���m���:����������ۼ�Ƽ<ⴼq"��,���Ff����üBHټN#�1��,�7�������%G�B���������
���~�ؼ��¼񻲼�o��R�������7CǼ� ݼ��/3�H�"���D�(��2G��t��1�� ��q	�`q ��-뼛ZԼqƿ��ư��������.<���ʼ7��������Zd�@����r��:�2� �����-z��W_�M�м�ϼ����v���h����뺼@Cμz�伛"���,��  �  �+'�U9(�O%����o�������4���ϓ��Ѽ¤��򳫼=������e�����a��iw�����)wռ���:�������;���u ��&��_(��F&�]��0�._��u�k�ؼ�ɼ��Ƽ��м��~����?�b����#��(���'�F#��Y�p�������:2�޼	{ʼgS���P��o���T���񑼻R��F���D���Dȼ��ۼ��� �3
�9��~m�d�"��5'��"(�p$����k��׀����pQҼd5Ǽ3�ȼWQּDf���7��uF�g�%�_W(�	~&��-!�������{�����Y�׼��ü�H���n��[R��le���N��*͛�#é��k����μT��S�������`��]��x$��(��v'�Y%"�rB���s���ݣ߼hRͼ^?Ƽy�˼�&ݼ�m��ف	����B!�T'�,(��%�����������i���y�e�мՇ�����������E���t���IZ������%^ռ@�����������о��n ��&�^X(�?&��T�~'��T��^�ؼ��ɼ>�Ƽ��м���T����1���&�#���'���'�<#��P�m������v(��	޼kuʼ�O��fO���o��XW��@���nY������N���Qȼ��ۼ�（� ��
����y�Ȝ"�D'��1(��$�:� ��Ǒ�����rҼVǼ��ȼ'oּ*������MQ�d�%��`(��&��6!�ʲ�?�6����=�꼨�׼4ļ�g�� ����s�����Qp��%4㩼����.�μrp�2o����������7�$� (�ֆ'��6"��T�7)�Ұ��T�߼f|ͼFiƼ�̼�Nݼ���֓	����,R!��  �  �DD�u`B�� :��=-������w���	���ȼĵ��j���kk�����:����|�V��H<��%|���R���$��l�ͼ���̪��C�"X!��d0�:l<�aC��C���<�m�/���PL��[��j�N�开>����	���(�I�7�t�A�eD��=@��96��@(��g�.q��󼳁ؼ�Z���B���������.����}�$M}��X���Ì�/K���*���ڶռ���R��s��I�&�4�4�U?��5D�T'B�o9��*����u��h���C�G�v}���`�j��.'.�y�;��DC���C��s=���1�2#����N���Qgм=P��+��4����F���ہ�T|�HG�����}֐������o���-ƼF޼�d��K��M��e�+��8���A��XD���?���4���$�!�ê�T�P
�6F�Y�����"�s43���>��5D��RB�A:��1-����,��(�����༞�ȼ,����j��UN����������R|� 8��D���`���8����>�ͼ���i��I<�;Q!�,^0��e<�(ZC���C�U�<���/����@��B���N�
��!�A�(��~�(���7�x~A�SYD��2@�a/6�m7(�_�j�{�wؼS���<����:��/���}�uV}��_���̌�V��t7��������ռ��������&���4��c?�ED�d7B�09�,�*�����[���
e�f7�ۛ��o�w�3.�I�;�eNC���C��|=�]�1��#����X����+м1j���F������e��y���	�|���������������򌱼JƼ,޼|�������y�+���8�M�A��iD���?�!�4���$��Q���6��5��p�+�D&�'�"��E3��?��  �  S	b�^�˟Q��?��1)���Z>��w�ּ黸����;Ŏ��	���o�#%d�'a��e���r������l���ӥ�nԾ��F޼f�.���2.�ŖC�M�T��_�V�a�'oZ�(FK��7�}�!�rp��X���U	����~t-���B�A�T�4�_�˰a��Z��K���7�D�!�Da�O�˼���FX��Y���~�z��Sj�4b�ʬa���h��ax�����7���^���rȼ��I�����5���I�xYY��Ja�4.`��V���D���/����Ц
� ��9����_d�
�4��+I��Y�Ea�4P`���V�ǾE���0����W�	⼦����7���;��|	��J;t��f�a�?0c�|+m�VP��ꌼ���q�����ҼT���1-���&�Ӷ<���O���\�]�a�R�]��Q�>�̟(����@��`c���5���D&��;��&O�w�\�F�a�=�]���Q��	?�&)����O'����ּ4�������+����퀼��n���c���`���e�%Tr�d���6T������~����4޼��*��8,.���C��T�M�_��a��fZ��<K��7���!�yc�*������F	�����e-���B�={T��~_�S�a���Z���K�<�7��!�Z��B�˼���qR������H�z��Tj�[!b��a�:i�:sx�����D���m����ȼ
-�	�W�ؓ5�`�I�5hY�'Za��>`��%V�3�D�h�/���P�
�1��I�*���r�9�4��7I�lY��Na�*Y`��V��E��0�Q�a��/�f ¼�P���V���%���vt���f��La��nc��im�,��!���Ȟ�=ϵ��Ӽ&����:�m�&�3�<�2�O��]��b���]��Q��'>�{�(��������y�)����8Y&�B�;��8O���\��  �  ��{��v��g��;P�U5���� ��HԼ�3��M���������l�g[�;2R��O��S��|^�0�q�J���훼�:���Mݼ������z;�b�U��Ck�^�x���{��s���b��]K��2�������5W�L��b�(�JW@�!�X�m��zy��]{��`r��`��G��,�{��;��<�Ǽ%g��܉����|�G�e��XW�OP�I$P��6V���c���y�2L���Q��^vü&��)����(�<D���]���p��z�+z�t�n�73[�]C�<++��p���g������40�T�H�/%`�g@r�'O{�X�y��-m�"qX���>���"�pB�X��"ӻ�/����'���t�o�_��<T�آO��_Q��Y�j�i����(��Z���C�ϼ�����k12�TM�X�d��8u�<�{���w��i�~mS�B�:�$$�0�������X�!�!8���P���f�9ev���{�|v��
g��/P��I5����= �~1ԼK������{���Wl��.[�p�Q���O�rhS�@G^��fq��2��K؛��'���<ݼU|�)���s;�z�U�w=k�ңx�A�{��s��b�SK���2�T��t��qH� ���(�H@�I�X��m�omy��P{��Tr��`�s{G� ,�������|Ǽ_��󃏼�|���e��YW�q�P��-P�DV�M�c���y�DY���`����ü��������(�-�D���]���p���z��;z���n��D[�MC�6=+����;����d�C0���H�01`�-Kr��X{�*�y�6m�"yX���>�H�"��K�Q��黼����A���Mt�D/`��xT���O�ޜQ��Z�8j�؁�E���ڭ�V�ϼ�������a?2��bM���d�:Iu��{���w��-i�؂S�|�:��:$�I$�������3
"��-8��P�g��uv��  �  ᆽ���#v�Ӊ\��o>�c�����ռ�r���ܑ�F�{��'a�g�P���H�òF��J�V�S��f�����j���"���߼����O&��OE�þb���z�$����"���:r�{�X��N>�~�'�Yd�3��f���i3�n�L�N�g�p�}�����~��7g��rRn���R��4�|���v����Ƽ�ʣ�B���_q���Z�(NM�$NG� G��JL�p�X��:n��臼�t���}¼���jX�U�0�riO�}k�'w��50������Ψ�m;j�v�O���5��!���(n� q%�tp;�i�U��o���������n����|��e�S�H�в)�y�F+����D��𗃼"�h��+U��J�<�F��H��}O�̪^���w�
$��󰪼'мY���+���:��JY�q�s����ĕ�2���_y���a��F��U.�b��M(�ߍ���+�QD���^�+w��能Fن����v��}\�d>��������Լ�Z���Ñ�<{���`�L�P��H�U{F�S�I�4�S�p�e�B���sU��J��\�޼����I&��IE��b���z��q����z���0r���X��B>�0�'�V�C��
��Z3�
�L�Fxg���}�9���`x��Ia���Gn�C�R�e 4����i��C�Ƽ�£�<���Wq�d�Z�OM�BSG�c	G�+XL�/�X��Pn����� ���C�¼d��Jc�K�0�xvO�'�k��~��+8�����)��BMj���O��	6��!�0#��~�Ȁ%�;���U��o����Տ��Ms�� }���e�9�H��)�`��>�,��\��;����h��dU���J�"�F��IH���O���^�U'x�+@��n̪�&BмG����8���:�vYY��s�	
��jՆ�ݏ���sy�y�a��G��l.�����?�Ϥ�,�nD���^��#w�B��  �  �������F�:)��M��e���R�o� �5����һ%������j�����t���q�ƨv�������� ���?޻����A���~��٢���ȼ+���$��k�N��{��-- �ܛ��.��A���#S������Y���9Ӽ�P��-�9L�
W�
�"����1ټA���D����	[��7%��������T��������4{��3r�b�q��y��ˆ��|��!���� ����HT�򊊼|E��ռ�o��:��������S�o���g�ּ���*O���s�����e�$����ݼx#����
��q����s�ke��̼��ϙG��A��c�\���-��Mރ�#�v��q��+s�8|~�/��S����̻���E�/���h�x�������#ἠ� ���ܶ������LB�§˼x��������W���閼�۪�HȼX�輵��G�W������9�V��5��
�����o��5�i���ѻ&���
���F��N�s���p��u�����Z���&`��L�ݻ۟��vA��f~��ˢ�W�ȼ"��4��d����؍��# �~��m��w��d8���鐼h=��Qֳ���Ҽ�4�m ��?�!K�
�����ټ>���\z��c�Z��$%����ƃ��+����|���8{��Gr���q�E�y��톻צ��K����Z�� ��mT�����\���ռ+���X���������c�����=�ּ�#���p������_<�����aŽ�/�ݼy;��|�
��{��
��|��v���̼������+�G�Bm���以�G|��5M���w���q��t��f�{��Hm���q̻����&0���h�򓖼���[A�� ��R���0��Lk�>�˼�譼����m�����\��T=ȼ<��s,�-X��  �  ��fV	�����߼F9��)㗼��l���4�6V	��tԻL��䎑�;o����y�W@v���{�х����<����V����-*@���z��П��Tļ�����n�
����H �������ۼ�l�������ΐ�T���Ǜ�����f�ͼ�,������������b����<Լ��r7���X���$�9���FĻ`����|��m5����v��Hv���~��������P��ʷ�.��a4R��]��5ʫ�\6мtj�h�M:�L�R��JT�:/Ѽ|���6������A������T����Tؼҷ��� �����T������Nȼ�ã������E��8�WS��p���+��	���n�{�7�u��w�����
��7{λG�X/�k�e�4ߓ�x���ۼ����n�����\
� ��P�ÛƼ\���$┼v�Q������\"ü*�����h�	�K�IH	�o���?�߼f!���˗��l�=�4��%	��Իך���$�����x��gu���z��j��w����R��+�Ⱥ��@���z�y�pGļ{�(��P�
�$���������p�ۼ�U��cw�������}��]��fq���ͼO�H��O�������U����*Լ�௼�)����X�6�$�����Z0ĻB����v��w7����v��lv���~�%߉�����.������J���YR�Nr���ૼ�Nмۄ��v�1I�������u��PѼX���ã��S$��߿��� ������nؼ��������^���԰�Y_ȼ�գ����SF�hd�����ն�e����*����|��lv�8�x��d��B����|��>�λFN��L/��f������'��mܼ� ��L���o
�3��y��Ƽ����������|��dߦ�?Jü��^���״	��  �  ���Ά���!��
ѼO@��-Ɛ� �e�@3�e��2�ݻ�����9���֌�焻�͂�M!�������u��/��K��;�=��Rr�ܗ������׼��� �_n�����c�O�˼��l6���͆�hۃ�����m���⾼|�ۼ��+�*,�w������>�ƼD��xU��Z�S���$��� � hλ󴫻̕�`#��Z>���킻�"��<铻U���Ŧɻ���V ���M��Ⴜk����ü�༾��w��>�������޼V¼�Υ�ɶ���:������ړ�Lī�a�ȼ̓�;���4�<�<S�¹ڼ�
���a���x�3�B�r��_����������h���r��-����+��v������pػ��s.�i_��,��g���s�ͼS_�$���z�r ��sռ�J��.���ъ��=������d���GҼ���������j��e�"�мq(������<�e�a3�X���`ݻ򋵻�͛��h��=x���_��7����!�����������Zq��f=��2r�s͗��q���׼�́ ��f�����SP��˼�֮�w������쿃��ݍ�����ƾ��ۼ���4�i ��r�����\�Ƽ74���G����S���$��� �Rλ����ƕ�w%��rH�������<��B��Uè���ɻ2��T9 ���M�v���㢢�T3ü[�༻���A�����%����޼�&¼�؏�I[��iՅ�����Rૼd�ȼ���-���)>���e�6�ڼ]��t����x���B�'�����`��!������܆��邻�g��������
{��/�ػW��Q.�<�_��G��e�����ͼ�}鼁��K��� ��>�L�ռ�t��쮝����"h��SE�����?��?mҼ���y����  �  h�hἯ�Ҽ����¢��G����_��5�����pͻ7���͟��N���[��U���.���\����Իy��0��H.>���i����������O�ּng㼊���ݼ#�˼,��kΚ�|E����o���j��0|�o|��%���{����ּ�������jݼ��˼�8���͙��w�ˇP��@)�i6
�j[�{�»�Ū�� ��� ��԰��}ҙ�����G���t�໡(��K%�a�K�.�y�r�3E���gɼ%�ۼbY�)O�l�ؼVļk��rؒ��0��0k�z�m�q4��
��_%��}sɼjܼu��V)�Qkؼ	}ļ"����쐼Bo�~B�&����)�ػ;���g���������"��D˝�5��AsɻT|�-X�/1�=EZ�:R��J���lȹ��^м��ZC�=���ҼeU����K����.v��vi�9�s� `��*��_���I~мXc�VJ�bLἶ�Ҽk������n0���V_��\5�9���f�ͻ򯱻�\���ܔ�Oꑻ����l¢������Իû���p��	>���i�{������7���I�ּ�X㼲�弒�ݼ��˼���x����,���o�m[j�f�{��`����������,�ּ�㼯��_Uݼb�˼�&�����v\��pP�~-)�t'
��E廮�»����%#��+����|왻����!ѿ�; �{E�`l%�%�K���y��ؖ�b]����ɼ��ۼ�v��m�'�ؼ�vļ"�������ur��pk�~n��Q���%��6?��X�ɼ`2ܼ¡�W<�{}ؼ�ļ0�������4o�ΨB�<'�}����ػ�)������������������D�������ɻ;��ď��e1�U{Z�im��͟�$幼�|мT8�e������Ҽ�|�����#ɋ�{�v�>�i�Dt�R����P�� �����м`���  �  �üަ���ƶ�y��k9��EY��a��:A�'�%���������H׻ڟ����������o^��*Ļ�ݻ����ѐ��+���G�Z�h�}~���e���3���������ɀ¼mͺ�ɼ��_◼� ���sb��KL�)H�_�V���t�B{��5L���䴼���i(ü�����I����َ��Wx���U�?7������"뻁)λsS�������U��Ņ���X˻[o绡y���5M4�]R��0t�橌��p���[��U��¼����_`��5[��ƴ����x��Y��H�c�J��_������r��џ��b��t���G¼�������g��C���cl��,K��X.�����:�,�໎!ƻOI���g���u���
����ӻ�l�[2��"�o�=�o]�C1��A��Eq���1���ǿ�� ü�,���Y��ö��������l�ޜQ��G�ԋO��0i��h��em��O������z�¼��������`���!���A��c�`��	A�b�%�����P�� �ֻ�+��@��#9���겻�û:ݻSZ��Wb��n+���G�D�h�hn���V��b%��0r�������p¼��������z͗��邼fCb��L�2�G�EeV�b�t�L`���1��+˴�����ü����	���y���ʎ��<x�ѺU��l7�b�������#λ�U�����g�������z˻��b�����m4��?R��Xt���������]u���	����¼�������<{��CՐ�*y�LY�M�H�p�J�.<_�#π�}�������x���¼ZZ¼�ƺ�6���z������w�l�YK��.�^��q����Йƻ�Ĵ��䬻`�$����AԻ���l�""#�2�=�pH]�AL��� ������<O���濼jAü�O��[~��"ݞ�v݉��7m�"�Q��mG���O�ni�����#���祯�
>���  �  Ū��̱��ٝ�s�����ڷ���ip�;D[���E�BT0����q����%ڻDԻR�ݻc(��Б�����#5��J���_�Bu����3���N��4��a桼����ޗ�O���<v�$FU�o9�m(���$�8-0���G��Wg��>�����ޜ�v����ڠ������h��i����U~�"Bi��T���>�� )�
��q�0,�ֻ�ջ��㻠��u��j�&�<���Q���f���{��[��I��%Ě�e_�����t��������ⅼ��j���J��2�#%��&�۲6���Q��Ur�Y[��/���p ��Hڡ������"���7��/��0Gw�9)b���L��W7���!�ru����)߻[�ӻ�1ػ�o��4�����-� PC���X���m��t��5ʋ��_�����Fa���2�������M���/�_�яA��;,�m$�c�*��>�)\�dp}�3��"���.������������Z���錼����9p�g[�ݷE��0�/���6�He�ٻʈӻ�ݻ����Y��}���4���J���_��t�����#���?��!����֡������̗�A��sv��U��?9���'�=�$�~�/�˴G�y#g�%��E���wƜ�W{��GƠ�ʔ���W��Z����;~��+i� �S�A�>�h�(�h��n��.�Rֻ�.ջ`��F@��,���&��:<� �Q��f��|�^q���`��vݚ�Pz��l������������k��"K��G2�a%��	'�%�6���Q�Y�r��r��0������������5��OK��w1��crw��Wb�M�m�7�"��������9�߻�OԻX�ػ���Ms�:����-�ȈC���X��n�l���7勼�{���.�����~�����ݏ�n���`���A�8�,��V$���*�
�>�7r\�׵}��S������  �  �|���숼����4I��/@�� ߋ�����h�� �u��_�/qF�.�,�;���xd��� l�n2�d7L�k�d�Ƽy�m��������N��6[��#��{w���ꇼ*ぼ|1r�'�[��B�	�(�v��%�e��h ����Ւ6� oP���h�Ğ|�k���c#������q\��=猼�����������n��bW���=��$�n�:���;�H_�S"��:���T��0l��B��h����������I�������f�����>H~�%�j�S��-9��� ��s�P��������&�b�>���X���o�#���bO��n��x�Q���k��牼�+��؇{��Hg�t�N���4��v�,3�ZV��g�����)��NC���\�v#s��5�����܄��`���>�����_D������|x� jc��J�V�0��&
���"��o���.��G�"�`�fv�a��T҈��䋼1��n(��Bǋ�=���	���Wu�}_��6F�U�,����Qm��$�l�
��.�32���K���d�H�y��}��߀���<��vJ��0���g���ڇ��ҁ�,r�/v[���A�?�(������~� ��O���_6�==P��|h��p|��w��`��Yy���K��،����|���ۘn�gXW��=�h�$���`���D�+l��c"���:�-�T��Ll��b��z��ת��>ǌ��`��嵌�v����0��e�~�D$k��ES�l9��=!�}����X��%�G&��.?���X���o����Oc���/�����e��%�������D��+�{���g�O�]<5����u�}��n��f�J>*���C�Y]��\s�KQ��l2��b����,���Y���8���a���;��ٽx���c���J�s1��R��r
��[��>	��%��L.�c�G��a���v��  �  �s\�w�q��L��
���2햼�*���š��q������������{��Z���=��)*�hd$�[e-�JXC���a�U�������ړ���6���[��NМ�8����P��3�����l���W��IB�Ю,�����i��g�1�׻mgԻ�~�o��<��'#�r�8��/N�hnc���x�����Ȑ�v����ɟ��ܡ�մ��$��<���Čp��P�@�5��l&���%�*>3�&�L��l��̆�!�������񹡼>.���]��BÑ��Ǉ��z���e�-WP���:��I%����"���F�ӍԻ�UֻK绒M�"!�� *���?��-U�^`j�'r�
��㓼V��������e��o`��'񑼓E���Pe�:&F���.��e$��(�$�:���V�T�w�oҋ�[���ٟ��ȡ�󬞼Aė������\���s�U�^�HI��3��G��C
�� �^ܻ.eӻ3fڻ��ﻃ4�o���L1���F�}=\��cq�[4��x��{Ֆ����ˬ��
X��|v��Hm��|�{�dZ��G=���)��!$�U#-��C��a�#z��w~���z������F��E����攼�?���䀼�l���W�h&B���,��g��>���3�׻pԻ��I�������"��}8�N�lDc��_x����V����������ҡ�����*���)���p�p�m P���5��q&���%�K3�ѱL���l��؆�$�������ˡ��A��s��6ڑ�=�����z�]�e�>�P�w;��%����~���O�⻿ջ��ֻ���-���R��O*���?��WU��j���61������[��|��I���{��l���d��ّe��iF��A/�m�$��(���:��W��&x������w��I���z㡼;Ǟ�mޗ�:���
x��
�s�!�^��I��3����;�
���7�ܻ��ӻ��ڻ�j��x��6���1��G��  �  �B���b�>b��$F��Gl���|��Y���a ü���������g���h����g�t�N�.�G��S�#o���������_���ʾ�%Eü=y�����&���>��Ă~��b[��R<��!��8���� �һ�f���^��-묻j`��T�ǻ��_j��8�)�/���L�kn�C���$v���ۭ��S��p�¼ܿ��-�������VP��~S���]��'J��I���Z��{�Iz��`0�������¼�h�������m������D-r��KP�#�2����R�S����ɻP����嬻�$�����Vhϻ��������9�M�W�tMz��ߏ�i����಼�|���%ü*���E������07��c�r��!U��G�j�L�!�c���P�������Y��N�¼ׂ��#ø�N3���E��7]����f�F��)����<�� �ۻ4z»�2�����"����5���Xػd=��
���'���B�!�b��I��f.���T���d��Y����¼؏������H�� H��;kg���N��:G���R��n��㊼5ޟ�+C������"-ü`c��%t���|������&a~�}A[��0<�]�!������]Uһ���������=����TǻZ#�';�S���/���L��Dn�����Ff��ͭ��G���u¼$���Q�������>M��Q��]��,J��I�b�Z�g{�I���W���I>���(��,�¼�{������>��������`r���P�5�2����,�����OʻA���~Z��ݕ������*�ϻ3�~��>�L+9�k�W�Fvz�W�����l���\���E@ü��������:��Y��bs��hU���G��%M��1d��%���������/w��1�¼����3ݸ�M��|_���w����f�k?F��-*��^������ܻAû>���'���튱�����ػ�������'P'��  �  l�7��b�͸��'>��������Ӽ���|\�6�߼�~ϼ�Q��ힼo����r���i�5�w������ؽ���Ӽ2=��Q��߼"^ϼ}��;L�������W�hO/����s컐Ȼ�`��oj��\,���{���_��eե�t����ڻ&������D���q��k�����z�żUټ���0U�aRۼ�>ȼ7į��Ŗ�Q��]"m�S�k�@����+��嬼�ż͎ټX�优弣�ڼ�2ȼ�կ��G��w�cBI��\#�6��e�޻����k^��_��NW��'4��ˠ�������dĻ�{绯���'+�#�R�L���@��x���zͼ�޼����㼠�ռ*j��&0��k*��cpz�<j�Gop�y.������a���ͼQa޼y�*���ռԐ�����3��� g���;�o��)��̍һ����Ρ�s���Б��0��B���費�λ����yB�5y7���a�̠���&��'彼ŐӼM���A���߼�`ϼ�1���˞�oL����r��i�,�w�7̌�+_��j����Ӽ�!��8�Dy߼ZIϼ�i��C:���냼��W��,/�&���'�3�ǻ�����Iѓ�;��� ��v�����enڻ���v����D�w�q�hZ���󬼓�ż�HټD�优L张Kۼ�9ȼ.����Ė��Q���'m�T�k������3��5לּ�ż��ټ���/��ۼ�GȼT쯼�_���:w�{wI�:�#�)����޻�n��_ԧ�R���ʒ�����6��]��Q�Ļ�������R+��S�.���U������ͼ.1޼��F;��ռx���	S��xN��׹z��Oj�L�p�#R��!0������.ͼ�~޼w-�����ռH���~4��<���Jg�<�������ӻ���V��ג��R[����������|i��Iϻ�T���y��  �  x�5���h�������X�Ҽ�i�8�����f ���o뼲�м�����֙������u���y��y ������*׼�q��d �X{�$5������˼ƫ�t���b�\���+��7�U�ջi����򊻕���ۂ�!����������nlû�񻝼���E���{�5��۽��Nܼ�s��G��������AǼvN��^Ԓ��V�����������R���ü%.༤�����f������hN߼�W��N���4��Y�J����e���!KǻX��4䒻Ņ�������@��L|��ǖ�������лb��d�&��yV�������iȼ9弘c���A�� ����"ڼ_(��������������a=��^E���_��fvͼ��3u���t��3 ������ռɛ�������n�{�:��c�!������=���X��N��+I�����9���㜻:Q����$z��5��h��q��������ҼPQ�6���������P�E�м����+���@u��<Q���U���ܞ�W칼

׼+S��V �xn������:�˼�����t���m\�ø+���>�ջ�c��F���_���ش����������Q���R���ûpn�˒�3bE���{�$���˽�=Aܼ�g���A�t�c�����C�ƼVM��Ւ�<Y��:����ǐ��Z����ü:�g�����������c߼�m���Ӡ�%M���K������
�ǻ�w���X��8���Q��쮃��扻�������	ѻ���.%'���V�����"����ȼQ�w}���O�� �����DڼL������Y!�������b���i��󂰼��ͼk���������@ �B��# ּ񴶼����)o���:���������]���=ގ�#Յ�NЂ��6�������`���ɷ�`��Y���  �  l�7�adp�+ܙ�FB����ă��:�	����O	�~@��CD����󀥼�9*��H㕼�����ȼN,����
�O���	�R���ڼ�������b�.�,��K��#̻����}n��Ɂ��*x��Hv��}�����v����Ը����7��I��₼�ͥ��Tʼ�c���<��i��s��3����ּ=h��䝼[7���h��0����*���Ӽ���&k�;�Q����n�＃=μ.é��}���O�m'�?!��ݼ����Uˈ���}���u�ѻv�E{��p7��H����ƻz���.5'���[�`�����$ּ�\���%���K����i�#�˼������JH��J��=������ݼO;��Yh�����e
��;;�v:¼�����<w�d=��|�8�ܻY>��q������z��=u�V
y�7���?-��mh��J�ֻ�6��[7��3p��ę��*��h��mk��u�	��2A	��!��w#�gl��]��Q�����L�������aȼ,輅��ȳ
�2���������ڼ5�����b�r,��'���˻�a��,��<s��yw�e�u��c|��^���a��{���v��t��H��Ђ�㼥�FEʼOV����#��2��"�K.���ּ!g���䝼�9��Bm�������2���Ӽ�
�r��B���S����＝Sμ�ک������<O��]����O��z���>����~�ܣv���w��䀻����z�� ǻ��`'�
\��,������;ּdu��:�Q��[�!����[	̼<������in���o���ݢ�j$����ݼ[��Hw���s
��%�DT�eS¼
֝�qw��G=����ZQݻ����~�x9���{��Gv�z����r���W߬�_Y׻"l��  �  ?�8�5�s�����i¼����:X�������&r��缎uƼ����T��	���+���xb��֜ͼ�*��A��m����T������@B߼��������[e�X-����y�ɻ򝢻�h���:~���s��q��x�ل�����o���G�综��L�J��ۄ������μ�9�u��J�SQ�A
�����ܼC��dɡ�R����ۑ�x��`����iؼAG�����f��޾�:M�2�����Ҽc+��Y���_ Q� j��r���똻8߅�ڐx��<q�z!r�׵{�X9�����Ļ�\��,�'��Y^�z��y���,,ۼy����
��q������2�� Ѽ�G���@��ﲐ��Ҕ�¦��¼�Q㼈� ��m��E
��h���Y�Ƽ&�����z�f>��P��ڻ�E���[��(遻X1u�?�p��Et�gÀ� ��?e����Ի!�
��}8��\s�l����R¼������qK�0��m���b�����RƼy���/���m���g��>���yͼa	�*2�A_�ŧ�O������.߼IṼ�y���8e��4-�Ɲ�|Qɻ}O�����f�}�>�r��q��ew��|��LG������组��c�J��Ʉ�����i�μG,��kE�M��	
�M����ܼ)��'ʡ�󲒼(���p~�������sؼ'S�����$��y���V������Ӽ�B��/���h4Q���8��V����^��^R��Auy��r���r���|�v����b��4_Ļ����$�'��^�d���b���+Cۼ����1�
���O�������;ѼRm���f��8ِ������榼u�¼�s�p� ���������u����4�ƼY̠���z��>�4��p'ۻO���jۑ��k��:v�"�q�VKu�NC�������۩�Pջ���  �  l�7�adp�+ܙ�FB����ă��:�	����O	�~@��CD����󀥼�9*��H㕼�����ȼN,����
�O���	�R���ڼ�������b�.�,��K��#̻����}n��Ɂ��*x��Hv��}�����v����Ը����7��I��₼�ͥ��Tʼ�c���<��i��s��3����ּ=h��䝼[7���h��0����*���Ӽ���&k�;�Q����n�＃=μ.é��}���O�m'�?!��ݼ����Uˈ���}���u�ѻv�E{��p7��H����ƻz���.5'���[�`�����$ּ�\���%���K����i�#�˼������JH��J��=������ݼO;��Yh�����e
��;;�v:¼�����<w�d=��|�8�ܻY>��q������z��=u�V
y�7���?-��mh��J�ֻ�6��[7��3p��ę��*��h��mk��u�	��2A	��!��w#�gl��]��Q�����L�������aȼ,輅��ȳ
�2���������ڼ5�����b�r,��'���˻�a��,��<s��yw�e�u��c|��^���a��{���v��t��H��Ђ�㼥�FEʼOV����#��2��"�K.���ּ!g���䝼�9��Bm�������2���Ӽ�
�r��B���S����＝Sμ�ک������<O��]����O��z���>����~�ܣv���w��䀻����z�� ǻ��`'�
\��,������;ּdu��:�Q��[�!����[	̼<������in���o���ݢ�j$����ݼ[��Hw���s
��%�DT�eS¼
֝�qw��G=����ZQݻ����~�x9���{��Gv�z����r���W߬�_Y׻"l��  �  x�5���h�������X�Ҽ�i�8�����f ���o뼲�м�����֙������u���y��y ������*׼�q��d �X{�$5������˼ƫ�t���b�\���+��7�U�ջi����򊻕���ۂ�!����������nlû�񻝼���E���{�5��۽��Nܼ�s��G��������AǼvN��^Ԓ��V�����������R���ü%.༤�����f������hN߼�W��N���4��Y�J����e���!KǻX��4䒻Ņ�������@��L|��ǖ�������лb��d�&��yV�������iȼ9弘c���A�� ����"ڼ_(��������������a=��^E���_��fvͼ��3u���t��3 ������ռɛ�������n�{�:��c�!������=���X��N��+I�����9���㜻:Q����$z��5��h��q��������ҼPQ�6���������P�E�м����+���@u��<Q���U���ܞ�W칼

׼+S��V �xn������:�˼�����t���m\�ø+���>�ջ�c��F���_���ش����������Q���R���ûpn�˒�3bE���{�$���˽�=Aܼ�g���A�t�c�����C�ƼVM��Ւ�<Y��:����ǐ��Z����ü:�g�����������c߼�m���Ӡ�%M���K������
�ǻ�w���X��8���Q��쮃��扻�������	ѻ���.%'���V�����"����ȼQ�w}���O�� �����DڼL������Y!�������b���i��󂰼��ͼk���������@ �B��# ּ񴶼����)o���:���������]���=ގ�#Յ�NЂ��6�������`���ɷ�`��Y���  �  l�7��b�͸��'>��������Ӽ���|\�6�߼�~ϼ�Q��ힼo����r���i�5�w������ؽ���Ӽ2=��Q��߼"^ϼ}��;L�������W�hO/����s컐Ȼ�`��oj��\,���{���_��eե�t����ڻ&������D���q��k�����z�żUټ���0U�aRۼ�>ȼ7į��Ŗ�Q��]"m�S�k�@����+��嬼�ż͎ټX�优弣�ڼ�2ȼ�կ��G��w�cBI��\#�6��e�޻����k^��_��NW��'4��ˠ�������dĻ�{绯���'+�#�R�L���@��x���zͼ�޼����㼠�ռ*j��&0��k*��cpz�<j�Gop�y.������a���ͼQa޼y�*���ռԐ�����3��� g���;�o��)��̍һ����Ρ�s���Б��0��B���費�λ����yB�5y7���a�̠���&��'彼ŐӼM���A���߼�`ϼ�1���˞�oL����r��i�,�w�7̌�+_��j����Ӽ�!��8�Dy߼ZIϼ�i��C:���냼��W��,/�&���'�3�ǻ�����Iѓ�;��� ��v�����enڻ���v����D�w�q�hZ���󬼓�ż�HټD�优L张Kۼ�9ȼ.����Ė��Q���'m�T�k������3��5לּ�ż��ټ���/��ۼ�GȼT쯼�_���:w�{wI�:�#�)����޻�n��_ԧ�R���ʒ�����6��]��Q�Ļ�������R+��S�.���U������ͼ.1޼��F;��ռx���	S��xN��׹z��Oj�L�p�#R��!0������.ͼ�~޼w-�����ռH���~4��<���Jg�<�������ӻ���V��ג��R[����������|i��Iϻ�T���y��  �  �B���b�>b��$F��Gl���|��Y���a ü���������g���h����g�t�N�.�G��S�#o���������_���ʾ�%Eü=y�����&���>��Ă~��b[��R<��!��8���� �һ�f���^��-묻j`��T�ǻ��_j��8�)�/���L�kn�C���$v���ۭ��S��p�¼ܿ��-�������VP��~S���]��'J��I���Z��{�Iz��`0�������¼�h�������m������D-r��KP�#�2����R�S����ɻP����嬻�$�����Vhϻ��������9�M�W�tMz��ߏ�i����಼�|���%ü*���E������07��c�r��!U��G�j�L�!�c���P�������Y��N�¼ׂ��#ø�N3���E��7]����f�F��)����<�� �ۻ4z»�2�����"����5���Xػd=��
���'���B�!�b��I��f.���T���d��Y����¼؏������H�� H��;kg���N��:G���R��n��㊼5ޟ�+C������"-ü`c��%t���|������&a~�}A[��0<�]�!������]Uһ���������=����TǻZ#�';�S���/���L��Dn�����Ff��ͭ��G���u¼$���Q�������>M��Q��]��,J��I�b�Z�g{�I���W���I>���(��,�¼�{������>��������`r���P�5�2����,�����OʻA���~Z��ݕ������*�ϻ3�~��>�L+9�k�W�Fvz�W�����l���\���E@ü��������:��Y��bs��hU���G��%M��1d��%���������/w��1�¼����3ݸ�M��|_���w����f�k?F��-*��^������ܻAû>���'���튱�����ػ�������'P'��  �  �s\�w�q��L��
���2햼�*���š��q������������{��Z���=��)*�hd$�[e-�JXC���a�U�������ړ���6���[��NМ�8����P��3�����l���W��IB�Ю,�����i��g�1�׻mgԻ�~�o��<��'#�r�8��/N�hnc���x�����Ȑ�v����ɟ��ܡ�մ��$��<���Čp��P�@�5��l&���%�*>3�&�L��l��̆�!�������񹡼>.���]��BÑ��Ǉ��z���e�-WP���:��I%����"���F�ӍԻ�UֻK绒M�"!�� *���?��-U�^`j�'r�
��㓼V��������e��o`��'񑼓E���Pe�:&F���.��e$��(�$�:���V�T�w�oҋ�[���ٟ��ȡ�󬞼Aė������\���s�U�^�HI��3��G��C
�� �^ܻ.eӻ3fڻ��ﻃ4�o���L1���F�}=\��cq�[4��x��{Ֆ����ˬ��
X��|v��Hm��|�{�dZ��G=���)��!$�U#-��C��a�#z��w~���z������F��E����攼�?���䀼�l���W�h&B���,��g��>���3�׻pԻ��I�������"��}8�N�lDc��_x����V����������ҡ�����*���)���p�p�m P���5��q&���%�K3�ѱL���l��؆�$�������ˡ��A��s��6ڑ�=�����z�]�e�>�P�w;��%����~���O�⻿ջ��ֻ���-���R��O*���?��WU��j���61������[��|��I���{��l���d��ّe��iF��A/�m�$��(���:��W��&x������w��I���z㡼;Ǟ�mޗ�:���
x��
�s�!�^��I��3����;�
���7�ܻ��ӻ��ڻ�j��x��6���1��G��  �  �|���숼����4I��/@�� ߋ�����h�� �u��_�/qF�.�,�;���xd��� l�n2�d7L�k�d�Ƽy�m��������N��6[��#��{w���ꇼ*ぼ|1r�'�[��B�	�(�v��%�e��h ����Ւ6� oP���h�Ğ|�k���c#������q\��=猼�����������n��bW���=��$�n�:���;�H_�S"��:���T��0l��B��h����������I�������f�����>H~�%�j�S��-9��� ��s�P��������&�b�>���X���o�#���bO��n��x�Q���k��牼�+��؇{��Hg�t�N���4��v�,3�ZV��g�����)��NC���\�v#s��5�����܄��`���>�����_D������|x� jc��J�V�0��&
���"��o���.��G�"�`�fv�a��T҈��䋼1��n(��Bǋ�=���	���Wu�}_��6F�U�,����Qm��$�l�
��.�32���K���d�H�y��}��߀���<��vJ��0���g���ڇ��ҁ�,r�/v[���A�?�(������~� ��O���_6�==P��|h��p|��w��`��Yy���K��،����|���ۘn�gXW��=�h�$���`���D�+l��c"���:�-�T��Ll��b��z��ת��>ǌ��`��嵌�v����0��e�~�D$k��ES�l9��=!�}����X��%�G&��.?���X���o����Oc���/�����e��%�������D��+�{���g�O�]<5����u�}��n��f�J>*���C�Y]��\s�KQ��l2��b����,���Y���8���a���;��ٽx���c���J�s1��R��r
��[��>	��%��L.�c�G��a���v��  �  Ū��̱��ٝ�s�����ڷ���ip�;D[���E�BT0����q����%ڻDԻR�ݻc(��Б�����#5��J���_�Bu����3���N��4��a桼����ޗ�O���<v�$FU�o9�m(���$�8-0���G��Wg��>�����ޜ�v����ڠ������h��i����U~�"Bi��T���>�� )�
��q�0,�ֻ�ջ��㻠��u��j�&�<���Q���f���{��[��I��%Ě�e_�����t��������ⅼ��j���J��2�#%��&�۲6���Q��Ur�Y[��/���p ��Hڡ������"���7��/��0Gw�9)b���L��W7���!�ru����)߻[�ӻ�1ػ�o��4�����-� PC���X���m��t��5ʋ��_�����Fa���2�������M���/�_�яA��;,�m$�c�*��>�)\�dp}�3��"���.������������Z���錼����9p�g[�ݷE��0�/���6�He�ٻʈӻ�ݻ����Y��}���4���J���_��t�����#���?��!����֡������̗�A��sv��U��?9���'�=�$�~�/�˴G�y#g�%��E���wƜ�W{��GƠ�ʔ���W��Z����;~��+i� �S�A�>�h�(�h��n��.�Rֻ�.ջ`��F@��,���&��:<� �Q��f��|�^q���`��vݚ�Pz��l������������k��"K��G2�a%��	'�%�6���Q�Y�r��r��0������������5��OK��w1��crw��Wb�M�m�7�"��������9�߻�OԻX�ػ���Ms�:����-�ȈC���X��n�l���7勼�{���.�����~�����ݏ�n���`���A�8�,��V$���*�
�>�7r\�׵}��S������  �  �üަ���ƶ�y��k9��EY��a��:A�'�%���������H׻ڟ����������o^��*Ļ�ݻ����ѐ��+���G�Z�h�}~���e���3���������ɀ¼mͺ�ɼ��_◼� ���sb��KL�)H�_�V���t�B{��5L���䴼���i(ü�����I����َ��Wx���U�?7������"뻁)λsS�������U��Ņ���X˻[o绡y���5M4�]R��0t�橌��p���[��U��¼����_`��5[��ƴ����x��Y��H�c�J��_������r��џ��b��t���G¼�������g��C���cl��,K��X.�����:�,�໎!ƻOI���g���u���
����ӻ�l�[2��"�o�=�o]�C1��A��Eq���1���ǿ�� ü�,���Y��ö��������l�ޜQ��G�ԋO��0i��h��em��O������z�¼��������`���!���A��c�`��	A�b�%�����P�� �ֻ�+��@��#9���겻�û:ݻSZ��Wb��n+���G�D�h�hn���V��b%��0r�������p¼��������z͗��邼fCb��L�2�G�EeV�b�t�L`���1��+˴�����ü����	���y���ʎ��<x�ѺU��l7�b�������#λ�U�����g�������z˻��b�����m4��?R��Xt���������]u���	����¼�������<{��CՐ�*y�LY�M�H�p�J�.<_�#π�}�������x���¼ZZ¼�ƺ�6���z������w�l�YK��.�^��q����Йƻ�Ĵ��䬻`�$����AԻ���l�""#�2�=�pH]�AL��� ������<O���濼jAü�O��[~��"ݞ�v݉��7m�"�Q��mG���O�ni�����#���祯�
>���  �  h�hἯ�Ҽ����¢��G����_��5�����pͻ7���͟��N���[��U���.���\����Իy��0��H.>���i����������O�ּng㼊���ݼ#�˼,��kΚ�|E����o���j��0|�o|��%���{����ּ�������jݼ��˼�8���͙��w�ˇP��@)�i6
�j[�{�»�Ū�� ��� ��԰��}ҙ�����G���t�໡(��K%�a�K�.�y�r�3E���gɼ%�ۼbY�)O�l�ؼVļk��rؒ��0��0k�z�m�q4��
��_%��}sɼjܼu��V)�Qkؼ	}ļ"����쐼Bo�~B�&����)�ػ;���g���������"��D˝�5��AsɻT|�-X�/1�=EZ�:R��J���lȹ��^м��ZC�=���ҼeU����K����.v��vi�9�s� `��*��_���I~мXc�VJ�bLἶ�Ҽk������n0���V_��\5�9���f�ͻ򯱻�\���ܔ�Oꑻ����l¢������Իû���p��	>���i�{������7���I�ּ�X㼲�弒�ݼ��˼���x����,���o�m[j�f�{��`����������,�ּ�㼯��_Uݼb�˼�&�����v\��pP�~-)�t'
��E廮�»����%#��+����|왻����!ѿ�; �{E�`l%�%�K���y��ؖ�b]����ɼ��ۼ�v��m�'�ؼ�vļ"�������ur��pk�~n��Q���%��6?��X�ɼ`2ܼ¡�W<�{}ؼ�ļ0�������4o�ΨB�<'�}����ػ�)������������������D�������ɻ;��ď��e1�U{Z�im��͟�$幼�|мT8�e������Ҽ�|�����#ɋ�{�v�>�i�Dt�R����P�� �����м`���  �  ���Ά���!��
ѼO@��-Ɛ� �e�@3�e��2�ݻ�����9���֌�焻�͂�M!�������u��/��K��;�=��Rr�ܗ������׼��� �_n�����c�O�˼��l6���͆�hۃ�����m���⾼|�ۼ��+�*,�w������>�ƼD��xU��Z�S���$��� � hλ󴫻̕�`#��Z>���킻�"��<铻U���Ŧɻ���V ���M��Ⴜk����ü�༾��w��>�������޼V¼�Υ�ɶ���:������ړ�Lī�a�ȼ̓�;���4�<�<S�¹ڼ�
���a���x�3�B�r��_����������h���r��-����+��v������pػ��s.�i_��,��g���s�ͼS_�$���z�r ��sռ�J��.���ъ��=������d���GҼ���������j��e�"�мq(������<�e�a3�X���`ݻ򋵻�͛��h��=x���_��7����!�����������Zq��f=��2r�s͗��q���׼�́ ��f�����SP��˼�֮�w������쿃��ݍ�����ƾ��ۼ���4�i ��r�����\�Ƽ74���G����S���$��� �Rλ����ƕ�w%��rH�������<��B��Uè���ɻ2��T9 ���M�v���㢢�T3ü[�༻���A�����%����޼�&¼�؏�I[��iՅ�����Rૼd�ȼ���-���)>���e�6�ڼ]��t����x���B�'�����`��!������܆��邻�g��������
{��/�ػW��Q.�<�_��G��e�����ͼ�}鼁��K��� ��>�L�ռ�t��쮝����"h��SE�����?��?mҼ���y����  �  ��fV	�����߼F9��)㗼��l���4�6V	��tԻL��䎑�;o����y�W@v���{�х����<����V����-*@���z��П��Tļ�����n�
����H �������ۼ�l�������ΐ�T���Ǜ�����f�ͼ�,������������b����<Լ��r7���X���$�9���FĻ`����|��m5����v��Hv���~��������P��ʷ�.��a4R��]��5ʫ�\6мtj�h�M:�L�R��JT�:/Ѽ|���6������A������T����Tؼҷ��� �����T������Nȼ�ã������E��8�WS��p���+��	���n�{�7�u��w�����
��7{λG�X/�k�e�4ߓ�x���ۼ����n�����\
� ��P�ÛƼ\���$┼v�Q������\"ü*�����h�	�K�IH	�o���?�߼f!���˗��l�=�4��%	��Իך���$�����x��gu���z��j��w����R��+�Ⱥ��@���z�y�pGļ{�(��P�
�$���������p�ۼ�U��cw�������}��]��fq���ͼO�H��O�������U����*Լ�௼�)����X�6�$�����Z0ĻB����v��w7����v��lv���~�%߉�����.������J���YR�Nr���ૼ�Nмۄ��v�1I�������u��PѼX���ã��S$��߿��� ������nؼ��������^���԰�Y_ȼ�գ����SF�hd�����ն�e����*����|��lv�8�x��d��B����|��>�λFN��L/��f������'��mܼ� ��L���o
�3��y��Ƽ����������|��dߦ�?Jü��^���״	��  �  �Iw���m�h�T�VV0����bܴ���L�
����I�9�ģ:,X�:��;�;�;�n;��;56;R;�C�:��:�\�7�H˺xwm���ǻ<W�F+9��[��uq�K�v��-k�a�P�`s,��b�N̻�Z��#����붻U���J�:>A��`���s�� v�"g�8�I��d"�N��P6��3���F�5j0:���:5�:e@
;�;��;1;g;�.;]��:��:�O:1T���s�����u���E��Nd���t���t��}c���D��U�����G������b��ƻ�/�,�'�P�L�h�h�?Sv���r�~�^�_W=����л��}�� 庐3��X�:���:iX;�;��;
J;;qV;�;af�:�ί:9��9�{�R<�E2���� �Ғ+�-$Q�I�k���v� �p�u�Z��8�͓��*߻�᭻����)��tػ�c��4�QW��o��w���m�J�T��#0��u��|��B�K��4��of�9#U�:���:�|;�;$�;IA;"�;��;��;���:ta�:��7�+ʺ��l�cǻ�9�d9���[�MWq���v��
k��cP��I,��5�i�˻����mT��D���Oh�^�A���`���s���u�A�f��I�NC"����v��e��$�_N1:�O�:di�:0K
;��;��;(�;%�;�
;�:B�:9JM:`D���oZ��;仵��J�E�ƃd�a-u���t�V�c�6E����G���Ż�����ڡ��}ƻf�H0(���L���h��|v���r��^�#|=��/�9.ѻ/i~�ao�&�
����:�j�:L�;|�;�;Be;v!;p;d�;��:��:��9�t~�-�<�n����� �-�+�!aQ�X�k�zw�q���Z�~/9���� �߻����V����˪��ٻ���P 5�a�W��Go��  �  n�n���e��KM���)�e� �K���=D�#4��xk�9ė�:���:�;E�;�;g�;��;'�
;�m;��:�r�:$%8 ºd�����
�r2���S�:�h�N2n���b�]�H���%��� �{1û�M��┻�`�����zG��!:�/�X�bk�Hm���^�EeB�}s���%O��@$�_
�g0:�4�:���:X�;I�;�;� ;[�;�	;OS�:�:��M:��ѹo��u��^ۻ<��$]>��#\��Cl�R�k�Z[��=�C3���Y�����f��������R�!�.@E�Zm`�d�m�`(j��V��x6�4���ɻ��s���ں�_θT̀:���:T�;j#;p;�];�;R;�;��:6g�:���9z�m�A^4�����\���BO%�T�I��Hc�n�2h�;�R�2�<��:�ջ�����,����ϻ����-��O�c�f��Ln�iKe��M�"�)��� �������C�)���U��9F)�:��:R�;��;�;V;J�;��;�-;m�:�Ì:�:8A�����c��ۿ�6�	�U2�K�S���h��n�W�b���H�)�%��� ��»�電�z��n���Bc�0���9��X���j�.m�I�^�@B��Q�&��i��P������0:���:(�:�;��;��;��;�;vz	;%��:�S�:B$L:�չ���qÊ�R�ۻj����>�fX\�>{l��0l���[���=�7r�����H&���ޙ������'��_�!��oE���`���m��Oj���V��6�@���Qɻ�rt�Z<ܺ:���~:(@�:-� ;�G
;\�;
x;*&;6;`3;5>�:o��:D�9'q�85�������|�%� �I�c�X_n��xh�cS�,P2����+ֻ�5��QГ�ݓ���ϻw	��?.��O�W�f��  �  ��U���M�
8��T�%��HP���1��������99��:J��:9|�:��;�3
;9;G�	; O;.��:���:��:f@�7���/XM�K���.�����[�=���P�J�U��+K��3�Ԉ��%�ra��V~���G}�,���nǻ?�&�zB��R���T�B�G�R@.�LE���ͻzj��NX���� :fð:��:�s;x�;Tr;#�;ac	;��;�N�:�L�:S<:<���F6����x���Ļ(�d�*�WE���S�_S��XD�qL)����9�ͻ����~��Ȃ�=����ۻ=��s+0���H�� U��Q�"q@�K�#�8����t���Z[���ź񨾸�l:՞�:q��:je;
<
;��;�P;�;�n ;���:ڟ:���9�{W�׃"��ꓻ�޻�/�;�4��K��|U��P��y<���������B�����z������=���j�X��!�9���N�:�U���M�C�7�t"����^�<M0��>��Y�9�,�:�*�:�$�:�z;�;*�;.
;[;~�:��:�*�:r�"8'q����L�C���l�������=��P�loU�YK��p3�J_���⻹�����z|��Õ� ǻH�|�%���A���R��T��G�m.�$��Hͻ7��� �.o�Wh!:��:���:�~;��;z^;w;21	;>Y;��:���:+]::b�¹O���y��-Ż3���*���E�9T�I�S���D� �)�v��λ�������?��@*��ܻ��[0�(I�/*U��R��@���#� ������[�i'Ǻ�`ո1i:d�:)�:�;[W	;&;�f
;A3;��:���:��:W �9#�Z��]#��X��،޻�i���4�UL���U��VP��<�G��c����㺻N����S{�+K���ش�o �%���9���N��  �  ��1�y{+�n��� ��*Ļz`��;��XS����r8Z/Y:켯:���:SZ�:2� ;��;��:R��:�1�:�G�:��2:��!��ī��6������ѻ�F������-��o1�aE(�����e�q����~�G���;��d�P��C�ջ�.�g ���.��0�n�&�Q��c|�p����g�8(��CN"��l�9*v�:aQ�:'�:�x�:d�;
�;VS�:o�:���:�Ϗ:��99 ��͈Z�uS���������$�K;0� �/�_U"���
��ܻ*����Sk�'�<��B�u;|��Ү��o黲���Z&��0�h�.��� �q+	� Iػ� ���YB�����#���#!:�$�:���:�:1��:�m;_	;�?�:�7�:D�:�n:cf39
ze����r���鼻IT����&�)�b|1���,�T��Z���LȻ`ȑ��MV���8��uP�%������~���
��/+�ߓ1�D+��������B�ûE ��z��0̄�cj�8vf\:�c�:���:�:w�;�x;�` ;�l�:��:�¤:�|5:[��f���`o6��S��Άѻ�(�br�F�-��N1��!(�����/��f���t�F�^�:�M�c��蜻(}ջ���}7 �7�.�'�0��|&����:컼5���:g�B{��E1!��,�9�Ǉ:���:�;�:!o�:z{;�;$��:���:T�:��:�c�9��^1�	#[�����V������$�+r0�X�/���"��9�S�ܻg#���Jl���=�M�C�o}�4>��-���)�&��1��.�� �SQ	���ػdO��"�B��e������+:i��:x��:Z@�:W��:��;;e�:�b�:�v�:lk:��%9��h��y�,���?Y������mV��*���1���,�o��V���Ȼ5f��3�W���9�;�Q�� ��;`»���M�jn+��  �  ���x��%��9λ�����xq�D !������}���69��<:V�:Di�:eQ�:���:�:q�:�܊:��:�{87�ZsӺ�2�Q,�������ֻ,�����x���e����ݻ!/��m���,����U޺"���W��q��T_ʻ�8�\m�'L����y组\���;���5U���	���iz���9�9��g:⪦:-;�:�l�:���:���:���:�u:7	�9�:���}��#���K�<��;\�����sU ������a\����λ<k����`��q���ߺ���If$���t��j����ػ0��vZ�}�\����ڻ������r":�l��bL�S�? ::0��:_f�:^u�:r�:���:>)�:S3N:�ǅ9aEݹ��i���Mg�����GSɻP9�S���Z�JO�` �?���;��,�D����BٺdN �h&<��䉻S{������)�
I���������ͻ3�����p��= �����O�B�C9�"@:��:-�:��:��:���:�"�:�|�:?�":nx;8�e4�|8ҺZv1��聻�U��6�ֻ�\��h���I��#Oݻ.ݯ���~��,�(��]�ܺ!O�W������ɻ���@�"����������u��j�T�ř�`"��*���\{�9N�g:��:>1�:�D�:�N�:��:�>�:E�s:��9�fA�K��� �4L��l������w)�� ��m;������]ϻ$埻��a�-e�#��)�뺟E%�Pmu�qϪ��ٻv��q���+����R(ۻg��������:��j�qcO��+'�y�:���:�'�:��:\��:��:L�:�K�:�J:C}9*C么�����~'h��*��h�ɻ���)�����V�껾L��ҏ�^ F��V���ۺ����P=��t�����.��xg��  �  �������P��u��ݥ���Zr��jC�,����Һ��w����Xݚ9a�O:��:���:�Ë:�6:p�09&0����P溇��ĹM�!�|�����1Ū�κ��g»��� |����O^��[������5-����H�w�JH�G�<������c�������6»WP�������P��¯���$b�!�3��T�������<�3���l��9�-u:a8�:��:Q�:��:�̅��(�?-��y� �A.��c\�<Ʌ����v\��W��»{9��ꥻ�	���D��B��ޥ���M�^���D����
�h3U��Ŏ�����?���P»;ٻ�ו��3◻g����FR�"$�g���^H��%�8(,:���:9�:!�:��_:ٱ�9>ke�V/a��JǺz��-s=�?Jl�����ɣ�W⵻�������p괻!���\v��+�d˺��Q��*�D�B������"��,n�Ug���ϲ��F��HF��q���a��yD��ǘq�k�B�6���%Ѻtwt�w������9��S:�Ĕ:ݐ�:`��:ң9:�X>9��Ṱ���m���%��!M��A|��i������ ����&»�u���4���v����]����X��A*����ot�5��n�;��3�����˧��������@R����?w��W�a�93������I�;����X��9�u:2�:�؝:�:��:b����*�����x�Պ.�[�\����t�$����X���y» ���j]������E�p$��c���W��uM#�����~���U��#������d�����»�(��嬻�2������R��$��0�6���,�����8�b(:\��:'�:��:=\:�9fNt���d��ɺ*���L>��"m����t8��mU�����w���m��RE���xw�}6,�;�ͺ��V���
�ЖG�I��I�#�f9o��晻H���  �  �z�L+�� ����9��0&���@��欇�1yx��%V��(�Up溔�o�à8�坥9n�99"u9+���Oݏ�.��5�3�3�^�r�~�����%���Y���Ґ��`������ds��O�h	 ��`ӺkK�����X��9b�9Ay-9�&�誡�yd�WN;���d�]-��5���ڑ��,I��O���K���6��=�m�e�G�%��N쿺Y'��58��9Y��9���8
�����R��*WB���i��ɂ��]������q���Ǝ����=��*�g���?����K;��#a���9�v�9C�9Ǔ�6'{1�%�źÙ���I�6Yo�0���0���O�� ��*;������=K���b�2)8�&���9��F�ʹmS9]��9�¿9u���T�?#غX."���P�/ct��@���R��瓐���֎�����]3|��[��
0�����|����N�����9���9}9�9�jM�lmw�.��̓*�TzW�[2y�6���P���֐��Đ�xߍ��I���w�=RU�:�'�:��W�k�n�)�+<�9O�9"�9qO�����p��W�2��^���}�c0���ێ�&��֏��/���ͅ���r�0�N��q�Һ*�H�ئx����9���9��99�߹�,����a�:���c��܀�(H���L���
�����s��X���m��cG�C������Y'���8���9���9⭺8�������(�7�B��9j����̨��T���U��3폻�W���}���h�Ms@�"l�3����]�8
>�9 �9i�޶��4�Ǻ�T�tsJ�p�`���	Ќ�����%s������[��=���1�b�\9�>�����M�ҹ]{C9Գ�9f��9D�4�W��ں�#���Q��@u�������������_���������'}���\��1��'������b����9���91�9�_�ް{����~�+��eX��  �  aO��F�|�t�푻 ������r���zJ���%��{*��.
k�]��y���?v@�@�&K^�ywԺ�K0�ir{�}ٞ�+a��0���ɶ��Il������Y����Xj�@�;�!�h�ú�yZ�d�L�o��9k�b:�ʗ:;&�:���:":���8F���蜺xp���
'�U5U��.��b?��縭�%����w»��Xj�����+MQ�[��d������	�����D����H�) ���|������7»{���m���b���u����Y�~Q+�����&ۤ���2��7��:��:J��:ٛ:�&q:���9
Z�q�D�%ٸ�0��]�5���d��ډ�`Z���V��$���f���qܷ�����G����7��ຨ]k�r�	�7�/�������Ϳa�^1��\���꾻V����Ź�m\�����bsy��\J��u��ߺ�p��WιH[b9)�@:�Ï:��:[W�:��M:�X�9�@���}���պ�t�;4E�{6t�����0��+P��F����⿻ι�������j����L���`�<��L��bZ�U�Һ�`/��z��p�������Z��~c����6���!x��e�i��;������ºvX�j�B����9��e:�5�:L��:�q�:�q%:��8������y!�!m&�x�T�l끻I��q����d�� O»g��� P�������5Q�V��o�������扺�����H��N�������X���{»sŽ�Ӿ��ǹ���҄�
tZ�� ,��T������ �!� F7h�:?�:ҝ:c�:�m:q�9�����G��<��;	���6�+)e��-��ɯ��$����￻�3»pG�����A���]�8���⺡zo�7����3�p�����b�����6ϯ��Y���X»T0���Ʃ��|��Pz�AK��c��ấu��ifֹQ9�u<:ы�:���:�&�:�{I:��9i3��uŀ�x�׺�  �  �˽�8>%��1v�h��pл7���n�Ak�J��,Z�W���Ƈ��9�Bn��`�ۺ7���`J��x��D�»��������%�����wmǻ*����Xc�h�"�����̹���9g,R:EU�:�T�:�h�:���:��:Z��:1��:�Q
:c����_Z��H���>��1��]���
ݻg���V�D%�"����sֻ�ܧ���o�?'!������⺡$�"�e��R����ѻ�:���m����m��H���������G����;p�q9��#�9Qy|:���:��:��:�t�:�A�:�Ԥ:�1b:+ʸ9<���}Β����Y�Y�����»q�軘A��F�m����_�ǻ�`��bzR�\��|ۺ�+���/����(�� ~߻�9 ����������iԻת��~�x�,���ʺY�'�4�8s�*:q��:0z�:�0�:��:�T�:ot�:�2�:�_9:�� 9Y������p$��ju�����л�r�?<��6�c��5���޷�J���8��e���ٺx��dI�����Qg»�5����c��]����h"ǻ�c���b�Z���h��33ȹLL�9��T:ן�:a��:���:9�:�0�:��:��:~:����W���J>��`\����ܻ����B���1���,aֻOѧ��o�-!�m����V�f��y���ѻ�o����E��ö��g%�%\��"��w�G�߮����s����� �9��x:6�:U��:<��:���:���:m?�:Y)_:���9{��&��Y�>.Z�+ٗ�.�»O!�Er�zz���5����ǻrᗻ0�S��j�M�ݺIJ���0�����������߻�s ��)�E9�����ԻA��L��y�-��X̺8�+�8Ԏ87�&:=��:EX�:;	�:���:4�:�_�:�.�:�5:��9���  �  ����%�b���F�ǻ�����C%,���1�b�*�r��T�����[�����N��:�H�Z����a$̻��6��[-�V�1��?)�� �[y��Eڹ��{�ν��V���[9y�t:���:߅�:���:��;d�;��:���:�f�:3��:[�:y����ȺR�H�B~����ۻ�
�4�!��E/���0�c|%�����I�?m9x��RA��K>���o��ѥ� �߻ɑ�>q#�-�/��/�c�#�}�:1��줻4BT��ۺh߹�:A�:ˑ�:x�:���:`P;��;n8�:�4�:qW�:S��:�p�9��1�3�H�m�w�����((�i'��1�1>.����w��6һ���E`���9�
�H����N4���K�7��(�g1�q+-��@�;��5λ�搻X0�B���
"��@:P�:��:_��:�� ;��;�^;�-�:,��:ϊ�:�WS:���7b獺H�$��H��\5ǻ*v�J��P�+�t�1��{*��������,���6	����M�r�8��Y�������˻-Y����s'-��l1��)����,�����j�z�
2��rT���d9�v:��:���:,�:�>;Bc;���:.��:��:$ �:Y: s��Q~Ǻ�%H�0=���ۻ��
��!��1/�<�0��o%�\��Z>�꫻r?x�9gA��n>��o�����߻Ѩ�Ë#�!0�^0���#��������G���U�]ݺ���f�9�W�:���:R��:y�:t;W�;]��:��:ֽ:ȅ�:q�9��4�����]n��
��a��3W��'�M1��v.� \�O���һL����[a��;�C�I�뛅��������dS��&)���1��a-��u�`���oλ9Q���21�	l���ԸF<:JU�:��:���:��:/�;IU ;<&�:G��:��:��O:��6�  �  �č�Y8��X���"뻬E�֋9�
�N���U�k�M�!S8�C�?B��䱻B����{�hi����!?��� � %>�>Q���U�K�^N3�/d��Eڻ�N���s�4XE����9��:=��:/\ ;i�;ƽ
;�?;�p	;�f;��:f/�:��^:��+�UvҺ�c�8���V���n%�=�A�"�R�H�T�&�G��.���?ػqf�����@C�������<ѻ��	�u+���E�o�S�uS�/D���(���������Lq�K{麻N���I:n��:6��:];�	;Q�;[�;x�;�7;���:} �:��:�K�����(����ѻ6���/���H�p�T�:
R��@��$�7'���û}�����{�iX��C���:`�p<���4���K���U���O��E<����"%���UoE�ח����8�:q��:���:H�;W�
;p;	;xD;m��:A~�:�N�:[�n9�#���B7�%���t��3�VZ9��kN�%�U��M��8������>_��0��zz�bᏻ�n������=q �u�=��P��`U�*�J��#3��<�,�ٻ������� C�z.�9�>�:��:7� ;U[;�j;3�;�"
;�;�W�:��:D1a:��!�EKѺzb��s��)���T%�b�A��}R�&�T�z�G���.�n���:ػ�i��T���T��)����\ѻL�	�g5+��E�>T�7�S�sSD�I
)�%����r�B�!͞�R-F:�߻:
 �:�~;�	;Z;P�
;�#;/p;p�:�:H4:� ��B�c~��.�ѻ�c��0���H��#U�%DR���@�mN$��j��PĻ�B����|�K冻k;��O���|�K;5��-L�
�U��(P�{z<�r����}��SFF��T���8	�:���:���:Ǖ;2�	;[;�
;�E;���:��:���:�
a9�  �  `k���ML�O������,���N�of�v�n�N�e�(N�F1,�e��wj̻�ߠ��> ���ٻq&��K4�ˇT�_5i��-n��ob��H�+H#��E󻇔��n�-��MY�C2:��:'�:��;u�;�q;n�;e�;�?
;�T ;�R�:�Ss:I�:�~��&Z|���ͻ��َ8��-X���j�iYm�?O_�߀C���C������Ө���N���xb�ʹ?��\��}l���k�h�Z��m<�Rp���ֻ92�� \��C��O\:�{�:���:�d
;�Q;�v;LN;q�;��;/�: `�:p_":�)�6"�����~�黯��-D�#�_��ym�Q[j�BW�H 8�_�*�߻ܼ������B����Ż��x�'��J��c�|,n��g�K	R��,0����1��[[��³�H��8+�:u��:%;�;\�;v;��;��;u_;���:���:�ȃ9�͚�'�K������B�+�A�N��;f��Rn���e�:�M�q�+���R�˻V���d��c�����ػ;���4�AMT���h��m�EAb���G�& #�5��L��'�,��W��v:0�:�]�:�;>F; ;Jd;�i;N�
;�;>��:��u:�0�����{�5�ͻ���t8��X�&�j�aIm��B_��wC�p��<�����P���G����g��f���u���?�;�\���l���k���Z�/�<�����׻#����"�����0�X:U��:�
�:�	;:v;t�;�z;��;�;��:�:��:	�,�����ח���黙���]D��+`��m���j�Y�W��A8��G��g��K�����hН�pFƻ���m(��J�'�c��dn�'%h��=R�`0�]��Й���/\�nz����8-	�: �:�;�;��;@r;��;��;�j;s�:&7�:�z9�  �  \Y��9�T�?������2��V�/�n�}Iw�Un�c�U���2����ջ
�����~��":㻐���:;��r\���q���v�r�j�,�O��w)����������4���e�K' :sd�:���:]{;��;�j;\�;q�;H�;S ;�p�:��u:ǞU���N��V�ջH��?��5`��{s�yv���g���J��%��N �	qû�|���������.����!��G�@�d�X.u���t�o�b��C�o"��߻ܡ��1�q���]:�z�:�;�;�n;�f;zC;�;�
;���:q�:�B": �4���$�,�������$���K�CCh��4v�*�r�DD_�9?����v��8��ԛ�TX���λ>6��b.��$R��l���v�H}p���Y���6������»qod�ѓ��pz�8J��:a1�:f�;`;�;�`;��;x�;?�;�>�:��:{9󼢺DT�*'��t���d2�fV���n�vw�-n�[�U���2�
V��?ջ����H7��f���{��	��'�:��7\��q�ӹv���j��TO�_O)��X��V���;\4�0�c�@l:���:���:?	;H{;�;�Q;n;T;��;���:�'x:��K�jl�	��ʈջfb�f?�`��hs�{ v��g���J���%��L �+tû놠�����$������i�!��G��e�
Lu���t��c�)�C��L��l߻� ��c��Pό�Z:	��:/5 ;��
;��;��;3p;�;�X	;��:���:*{:��7�\�%��睻e����$�7�K��vh�lv�4s�Ă_�O?�u;��S껏Ǵ�#d��"祻�wϻz���.��bR��Ol�R$w�b�p�EZ�?7�7���»�Ce��I����8Sϒ:I�:]�;`;_�;D^;��;��;�;Ai�:�C�:��m9�  �  `k���ML�O������,���N�of�v�n�N�e�(N�F1,�e��wj̻�ߠ��> ���ٻq&��K4�ˇT�_5i��-n��ob��H�+H#��E󻇔��n�-��MY�C2:��:'�:��;u�;�q;n�;e�;�?
;�T ;�R�:�Ss:I�:�~��&Z|���ͻ��َ8��-X���j�iYm�?O_�߀C���C������Ө���N���xb�ʹ?��\��}l���k�h�Z��m<�Rp���ֻ92�� \��C��O\:�{�:���:�d
;�Q;�v;LN;q�;��;/�: `�:p_":�)�6"�����~�黯��-D�#�_��ym�Q[j�BW�H 8�_�*�߻ܼ������B����Ż��x�'��J��c�|,n��g�K	R��,0����1��[[��³�H��8+�:u��:%;�;\�;v;��;��;u_;���:���:�ȃ9�͚�'�K������B�+�A�N��;f��Rn���e�:�M�q�+���R�˻V���d��c�����ػ;���4�AMT���h��m�EAb���G�& #�5��L��'�,��W��v:0�:�]�:�;>F; ;Jd;�i;N�
;�;>��:��u:�0�����{�5�ͻ���t8��X�&�j�aIm��B_��wC�p��<�����P���G����g��f���u���?�;�\���l���k���Z�/�<�����׻#����"�����0�X:U��:�
�:�	;:v;t�;�z;��;�;��:�:��:	�,�����ח���黙���]D��+`��m���j�Y�W��A8��G��g��K�����hН�pFƻ���m(��J�'�c��dn�'%h��=R�`0�]��Й���/\�nz����8-	�: �:�;�;��;@r;��;��;�j;s�:&7�:�z9�  �  �č�Y8��X���"뻬E�֋9�
�N���U�k�M�!S8�C�?B��䱻B����{�hi����!?��� � %>�>Q���U�K�^N3�/d��Eڻ�N���s�4XE����9��:=��:/\ ;i�;ƽ
;�?;�p	;�f;��:f/�:��^:��+�UvҺ�c�8���V���n%�=�A�"�R�H�T�&�G��.���?ػqf�����@C�������<ѻ��	�u+���E�o�S�uS�/D���(���������Lq�K{麻N���I:n��:6��:];�	;Q�;[�;x�;�7;���:} �:��:�K�����(����ѻ6���/���H�p�T�:
R��@��$�7'���û}�����{�iX��C���:`�p<���4���K���U���O��E<����"%���UoE�ח����8�:q��:���:H�;W�
;p;	;xD;m��:A~�:�N�:[�n9�#���B7�%���t��3�VZ9��kN�%�U��M��8������>_��0��zz�bᏻ�n������=q �u�=��P��`U�*�J��#3��<�,�ٻ������� C�z.�9�>�:��:7� ;U[;�j;3�;�"
;�;�W�:��:D1a:��!�EKѺzb��s��)���T%�b�A��}R�&�T�z�G���.�n���:ػ�i��T���T��)����\ѻL�	�g5+��E�>T�7�S�sSD�I
)�%����r�B�!͞�R-F:�߻:
 �:�~;�	;Z;P�
;�#;/p;p�:�:H4:� ��B�c~��.�ѻ�c��0���H��#U�%DR���@�mN$��j��PĻ�B����|�K冻k;��O���|�K;5��-L�
�U��(P�{z<�r����}��SFF��T���8	�:���:���:Ǖ;2�	;[;�
;�E;���:��:���:�
a9�  �  ����%�b���F�ǻ�����C%,���1�b�*�r��T�����[�����N��:�H�Z����a$̻��6��[-�V�1��?)�� �[y��Eڹ��{�ν��V���[9y�t:���:߅�:���:��;d�;��:���:�f�:3��:[�:y����ȺR�H�B~����ۻ�
�4�!��E/���0�c|%�����I�?m9x��RA��K>���o��ѥ� �߻ɑ�>q#�-�/��/�c�#�}�:1��줻4BT��ۺh߹�:A�:ˑ�:x�:���:`P;��;n8�:�4�:qW�:S��:�p�9��1�3�H�m�w�����((�i'��1�1>.����w��6һ���E`���9�
�H����N4���K�7��(�g1�q+-��@�;��5λ�搻X0�B���
"��@:P�:��:_��:�� ;��;�^;�-�:,��:ϊ�:�WS:���7b獺H�$��H��\5ǻ*v�J��P�+�t�1��{*��������,���6	����M�r�8��Y�������˻-Y����s'-��l1��)����,�����j�z�
2��rT���d9�v:��:���:,�:�>;Bc;���:.��:��:$ �:Y: s��Q~Ǻ�%H�0=���ۻ��
��!��1/�<�0��o%�\��Z>�꫻r?x�9gA��n>��o�����߻Ѩ�Ë#�!0�^0���#��������G���U�]ݺ���f�9�W�:���:R��:y�:t;W�;]��:��:ֽ:ȅ�:q�9��4�����]n��
��a��3W��'�M1��v.� \�O���һL����[a��;�C�I�뛅��������dS��&)���1��a-��u�`���oλ9Q���21�	l���ԸF<:JU�:��:���:��:/�;IU ;<&�:G��:��:��O:��6�  �  �˽�8>%��1v�h��pл7���n�Ak�J��,Z�W���Ƈ��9�Bn��`�ۺ7���`J��x��D�»��������%�����wmǻ*����Xc�h�"�����̹���9g,R:EU�:�T�:�h�:���:��:Z��:1��:�Q
:c����_Z��H���>��1��]���
ݻg���V�D%�"����sֻ�ܧ���o�?'!������⺡$�"�e��R����ѻ�:���m����m��H���������G����;p�q9��#�9Qy|:���:��:��:�t�:�A�:�Ԥ:�1b:+ʸ9<���}Β����Y�Y�����»q�軘A��F�m����_�ǻ�`��bzR�\��|ۺ�+���/����(�� ~߻�9 ����������iԻת��~�x�,���ʺY�'�4�8s�*:q��:0z�:�0�:��:�T�:ot�:�2�:�_9:�� 9Y������p$��ju�����л�r�?<��6�c��5���޷�J���8��e���ٺx��dI�����Qg»�5����c��]����h"ǻ�c���b�Z���h��33ȹLL�9��T:ן�:a��:���:9�:�0�:��:��:~:����W���J>��`\����ܻ����B���1���,aֻOѧ��o�-!�m����V�f��y���ѻ�o����E��ö��g%�%\��"��w�G�߮����s����� �9��x:6�:U��:<��:���:���:m?�:Y)_:���9{��&��Y�>.Z�+ٗ�.�»O!�Er�zz���5����ǻrᗻ0�S��j�M�ݺIJ���0�����������߻�s ��)�E9�����ԻA��L��y�-��X̺8�+�8Ԏ87�&:=��:EX�:;	�:���:4�:�_�:�.�:�5:��9���  �  aO��F�|�t�푻 ������r���zJ���%��{*��.
k�]��y���?v@�@�&K^�ywԺ�K0�ir{�}ٞ�+a��0���ɶ��Il������Y����Xj�@�;�!�h�ú�yZ�d�L�o��9k�b:�ʗ:;&�:���:":���8F���蜺xp���
'�U5U��.��b?��縭�%����w»��Xj�����+MQ�[��d������	�����D����H�) ���|������7»{���m���b���u����Y�~Q+�����&ۤ���2��7��:��:J��:ٛ:�&q:���9
Z�q�D�%ٸ�0��]�5���d��ډ�`Z���V��$���f���qܷ�����G����7��ຨ]k�r�	�7�/�������Ϳa�^1��\���꾻V����Ź�m\�����bsy��\J��u��ߺ�p��WιH[b9)�@:�Ï:��:[W�:��M:�X�9�@���}���պ�t�;4E�{6t�����0��+P��F����⿻ι�������j����L���`�<��L��bZ�U�Һ�`/��z��p�������Z��~c����6���!x��e�i��;������ºvX�j�B����9��e:�5�:L��:�q�:�q%:��8������y!�!m&�x�T�l끻I��q����d�� O»g��� P�������5Q�V��o�������扺�����H��N�������X���{»sŽ�Ӿ��ǹ���҄�
tZ�� ,��T������ �!� F7h�:?�:ҝ:c�:�m:q�9�����G��<��;	���6�+)e��-��ɯ��$����￻�3»pG�����A���]�8���⺡zo�7����3�p�����b�����6ϯ��Y���X»T0���Ʃ��|��Pz�AK��c��ấu��ifֹQ9�u<:ы�:���:�&�:�{I:��9i3��uŀ�x�׺�  �  �z�L+�� ����9��0&���@��欇�1yx��%V��(�Up溔�o�à8�坥9n�99"u9+���Oݏ�.��5�3�3�^�r�~�����%���Y���Ґ��`������ds��O�h	 ��`ӺkK�����X��9b�9Ay-9�&�誡�yd�WN;���d�]-��5���ڑ��,I��O���K���6��=�m�e�G�%��N쿺Y'��58��9Y��9���8
�����R��*WB���i��ɂ��]������q���Ǝ����=��*�g���?����K;��#a���9�v�9C�9Ǔ�6'{1�%�źÙ���I�6Yo�0���0���O�� ��*;������=K���b�2)8�&���9��F�ʹmS9]��9�¿9u���T�?#غX."���P�/ct��@���R��瓐���֎�����]3|��[��
0�����|����N�����9���9}9�9�jM�lmw�.��̓*�TzW�[2y�6���P���֐��Đ�xߍ��I���w�=RU�:�'�:��W�k�n�)�+<�9O�9"�9qO�����p��W�2��^���}�c0���ێ�&��֏��/���ͅ���r�0�N��q�Һ*�H�ئx����9���9��99�߹�,����a�:���c��܀�(H���L���
�����s��X���m��cG�C������Y'���8���9���9⭺8�������(�7�B��9j����̨��T���U��3폻�W���}���h�Ms@�"l�3����]�8
>�9 �9i�޶��4�Ǻ�T�tsJ�p�`���	Ќ�����%s������[��=���1�b�\9�>�����M�ҹ]{C9Գ�9f��9D�4�W��ں�#���Q��@u�������������_���������'}���\��1��'������b����9���91�9�_�ް{����~�+��eX��  �  �������P��u��ݥ���Zr��jC�,����Һ��w����Xݚ9a�O:��:���:�Ë:�6:p�09&0����P溇��ĹM�!�|�����1Ū�κ��g»��� |����O^��[������5-����H�w�JH�G�<������c�������6»WP�������P��¯���$b�!�3��T�������<�3���l��9�-u:a8�:��:Q�:��:�̅��(�?-��y� �A.��c\�<Ʌ����v\��W��»{9��ꥻ�	���D��B��ޥ���M�^���D����
�h3U��Ŏ�����?���P»;ٻ�ו��3◻g����FR�"$�g���^H��%�8(,:���:9�:!�:��_:ٱ�9>ke�V/a��JǺz��-s=�?Jl�����ɣ�W⵻�������p괻!���\v��+�d˺��Q��*�D�B������"��,n�Ug���ϲ��F��HF��q���a��yD��ǘq�k�B�6���%Ѻtwt�w������9��S:�Ĕ:ݐ�:`��:ң9:�X>9��Ṱ���m���%��!M��A|��i������ ����&»�u���4���v����]����X��A*����ot�5��n�;��3�����˧��������@R����?w��W�a�93������I�;����X��9�u:2�:�؝:�:��:b����*�����x�Պ.�[�\����t�$����X���y» ���j]������E�p$��c���W��uM#�����~���U��#������d�����»�(��嬻�2������R��$��0�6���,�����8�b(:\��:'�:��:=\:�9fNt���d��ɺ*���L>��"m����t8��mU�����w���m��RE���xw�}6,�;�ͺ��V���
�ЖG�I��I�#�f9o��晻H���  �  ���x��%��9λ�����xq�D !������}���69��<:V�:Di�:eQ�:���:�:q�:�܊:��:�{87�ZsӺ�2�Q,�������ֻ,�����x���e����ݻ!/��m���,����U޺"���W��q��T_ʻ�8�\m�'L����y组\���;���5U���	���iz���9�9��g:⪦:-;�:�l�:���:���:���:�u:7	�9�:���}��#���K�<��;\�����sU ������a\����λ<k����`��q���ߺ���If$���t��j����ػ0��vZ�}�\����ڻ������r":�l��bL�S�? ::0��:_f�:^u�:r�:���:>)�:S3N:�ǅ9aEݹ��i���Mg�����GSɻP9�S���Z�JO�` �?���;��,�D����BٺdN �h&<��䉻S{������)�
I���������ͻ3�����p��= �����O�B�C9�"@:��:-�:��:��:���:�"�:�|�:?�":nx;8�e4�|8ҺZv1��聻�U��6�ֻ�\��h���I��#Oݻ.ݯ���~��,�(��]�ܺ!O�W������ɻ���@�"����������u��j�T�ř�`"��*���\{�9N�g:��:>1�:�D�:�N�:��:�>�:E�s:��9�fA�K��� �4L��l������w)�� ��m;������]ϻ$埻��a�-e�#��)�뺟E%�Pmu�qϪ��ٻv��q���+����R(ۻg��������:��j�qcO��+'�y�:���:�'�:��:\��:��:L�:�K�:�J:C}9*C么�����~'h��*��h�ɻ���)�����V�껾L��ҏ�^ F��V���ۺ����P=��t�����.��xg��  �  ��1�y{+�n��� ��*Ļz`��;��XS����r8Z/Y:켯:���:SZ�:2� ;��;��:R��:�1�:�G�:��2:��!��ī��6������ѻ�F������-��o1�aE(�����e�q����~�G���;��d�P��C�ջ�.�g ���.��0�n�&�Q��c|�p����g�8(��CN"��l�9*v�:aQ�:'�:�x�:d�;
�;VS�:o�:���:�Ϗ:��99 ��͈Z�uS���������$�K;0� �/�_U"���
��ܻ*����Sk�'�<��B�u;|��Ү��o黲���Z&��0�h�.��� �q+	� Iػ� ���YB�����#���#!:�$�:���:�:1��:�m;_	;�?�:�7�:D�:�n:cf39
ze����r���鼻IT����&�)�b|1���,�T��Z���LȻ`ȑ��MV���8��uP�%������~���
��/+�ߓ1�D+��������B�ûE ��z��0̄�cj�8vf\:�c�:���:�:w�;�x;�` ;�l�:��:�¤:�|5:[��f���`o6��S��Άѻ�(�br�F�-��N1��!(�����/��f���t�F�^�:�M�c��蜻(}ջ���}7 �7�.�'�0��|&����:컼5���:g�B{��E1!��,�9�Ǉ:���:�;�:!o�:z{;�;$��:���:T�:��:�c�9��^1�	#[�����V������$�+r0�X�/���"��9�S�ܻg#���Jl���=�M�C�o}�4>��-���)�&��1��.�� �SQ	���ػdO��"�B��e������+:i��:x��:Z@�:W��:��;;e�:�b�:�v�:lk:��%9��h��y�,���?Y������mV��*���1���,�o��V���Ȼ5f��3�W���9�;�Q�� ��;`»���M�jn+��  �  ��U���M�
8��T�%��HP���1��������99��:J��:9|�:��;�3
;9;G�	; O;.��:���:��:f@�7���/XM�K���.�����[�=���P�J�U��+K��3�Ԉ��%�ra��V~���G}�,���nǻ?�&�zB��R���T�B�G�R@.�LE���ͻzj��NX���� :fð:��:�s;x�;Tr;#�;ac	;��;�N�:�L�:S<:<���F6����x���Ļ(�d�*�WE���S�_S��XD�qL)����9�ͻ����~��Ȃ�=����ۻ=��s+0���H�� U��Q�"q@�K�#�8����t���Z[���ź񨾸�l:՞�:q��:je;
<
;��;�P;�;�n ;���:ڟ:���9�{W�׃"��ꓻ�޻�/�;�4��K��|U��P��y<���������B�����z������=���j�X��!�9���N�:�U���M�C�7�t"����^�<M0��>��Y�9�,�:�*�:�$�:�z;�;*�;.
;[;~�:��:�*�:r�"8'q����L�C���l�������=��P�loU�YK��p3�J_���⻹�����z|��Õ� ǻH�|�%���A���R��T��G�m.�$��Hͻ7��� �.o�Wh!:��:���:�~;��;z^;w;21	;>Y;��:���:+]::b�¹O���y��-Ż3���*���E�9T�I�S���D� �)�v��λ�������?��@*��ܻ��[0�(I�/*U��R��@���#� ������[�i'Ǻ�`ո1i:d�:)�:�;[W	;&;�f
;A3;��:���:��:W �9#�Z��]#��X��،޻�i���4�UL���U��VP��<�G��c����㺻N����S{�+K���ش�o �%���9���N��  �  n�n���e��KM���)�e� �K���=D�#4��xk�9ė�:���:�;E�;�;g�;��;'�
;�m;��:�r�:$%8 ºd�����
�r2���S�:�h�N2n���b�]�H���%��� �{1û�M��┻�`�����zG��!:�/�X�bk�Hm���^�EeB�}s���%O��@$�_
�g0:�4�:���:X�;I�;�;� ;[�;�	;OS�:�:��M:��ѹo��u��^ۻ<��$]>��#\��Cl�R�k�Z[��=�C3���Y�����f��������R�!�.@E�Zm`�d�m�`(j��V��x6�4���ɻ��s���ں�_θT̀:���:T�;j#;p;�];�;R;�;��:6g�:���9z�m�A^4�����\���BO%�T�I��Hc�n�2h�;�R�2�<��:�ջ�����,����ϻ����-��O�c�f��Ln�iKe��M�"�)��� �������C�)���U��9F)�:��:R�;��;�;V;J�;��;�-;m�:�Ì:�:8A�����c��ۿ�6�	�U2�K�S���h��n�W�b���H�)�%��� ��»�電�z��n���Bc�0���9��X���j�.m�I�^�@B��Q�&��i��P������0:���:(�:�;��;��;��;�;vz	;%��:�S�:B$L:�չ���qÊ�R�ۻj����>�fX\�>{l��0l���[���=�7r�����H&���ޙ������'��_�!��oE���`���m��Oj���V��6�@���Qɻ�rt�Z<ܺ:���~:(@�:-� ;�G
;\�;
x;*&;6;`3;5>�:o��:D�9'q�85�������|�%� �I�c�X_n��xh�cS�,P2����+ֻ�5��QГ�ݓ���ϻw	��?.��O�W�f��  �  'R)��-���K8��c�:O�=;�׉;�g�;���;h��;��;��;�;Դ�;O��;� �;7��;�N�;l�;���;�ս;R�;��;��(;"�:VPǹ��к�E�e�(�����͠���T8N�:q�';�qV;�^_;7�@;Ug ;�N-:�3�@�xY!��%���g	{����9���:)�\;�u�;f�;!1�;�+�;e"�;�R�;6��;i��;�y�;qD�;��;�)�;���;���;9�;@��;��f;Gq	;1�:��S��F��92#�W#������T�W�:)�:e�;;��^;<Z;}G/;���:5�_9�}�����P�&�3%� A޺���ѐp:��;Xpy;ȿ�;���;�<�; ��;���;fy�;���;�e�;���;�8�;��;E�;�	�;�;�ޮ;��;��H;]��:Q{�8ጟ��l���'��<��κ�ʹ!�:��;|�K;߼a;��O;��;�~�:��y�[����V��e(��M�MC��8O{�$��:o>;�8�;�ȫ;K=�;m9�;�(�;7A�;��;��;qU�;���;c �;֬�;���;KM�;�$�;0�;�H�;�F); �:�lù��Ϻ���(�@A�󛟺Yc}8���:�X(;'.W;{ `;^vA;�+;|U0:m�0�7��e� �wW%�&h�u�x���9[��:��\;ў�;���;�K�;A?�;o.�;IW�;��;���;�h�;A,�;?��;J�;ݠ�;���;-��;bJ�;6f;=�;�B:E�V�x���F$���#� J����X�)=:�N�:�:;	�];�XY;l.;t��:�S9m���O��ŗ'�_��x{ߺt^��"n:�;��x;�i�;;��;���;9#�;�z�;��;�[�;���;���;���;��;_��;��;���;�q�;��;*�G;Z��:Ӈ�8Fm��*g�K�(�N�.�кFGӹ�'{:m�;�eJ;և`;��N;��;�=�:�l��'����P��  �  l��^������#;&9��:F;���;ܬ;R{�;��;M��;�,�;4��;�w�;���;���;�C�;��;��;Z<�;n��;���;� �;F�1;�,�:��:����D�?@��	����|��g�9pF�:[�1;"__;�h;!!J;f;��b:T��qDǺX����<qߺ�6��s%:��;�c;��;\��;��;�P�;XQ�;��;9(�;�^�;�G�;��;t��;�]�;���;�.�;`B�;ע�;w�m;m�;әQ:���pҺ���J��FҺb�Ͳ?:��;.zE;�g;c;,!9;��:
b�9*Y�&��ح�j

�F︺o̐���:�!(;[�;鑣;�м;+��;��;l"�;��;v��;^7�;���;���;`�;}l�;7�;{��;�6�;��;V�P;�|�:�l�9�x����Ӄ��y�[���l��l��:Yn;z�T;#pj;�Y;$;S��:�iŶ;���O����O��k��I39��:��F;��;i=�;���;m�;RM�;m��;��;b��;�'�;BA�;&��;���;��;��;��;��;?F�;/]2;�*�:A�	�����8��Ÿ�a���=z��~�9q��:�[2;O`;��h;��J;�);��e:*�ํ�ź`��[
�D޺Փ4�f':'�;y0d;!ؘ;&��;���;d�;Z]�;ο�;�%�;�T�;�6�;���;g�;-7�;L��;���;��;
`�;.m;�;#�N:>o���Ӻ���F����ӺO �<:�;O�D;6�f;D5b;F8;�^�:�&�9T\�R��hW�ˬ
�[*�������ސ:��';4;�;�;�u�;�*�;�C�;���; ��;��;���;+K�;Va�;��;���;X��;�8�;�ɯ;���;��O;<��:�2�9�>|�7������ˉ��Ȭ��C.��6�:<;��S;<i;��W;��";uO�:a:�����v���  �  �����9���k��"�O:�;e�[;��;���;EO�;���;d��;d��;���;#N�;���;��;�T�;��;�>�;$�;׿;:b�;|�;��I;C�:�
:S�
�.s��Nf��8G���g��m:7
;c�M;Vx;Z=�;��d;�*;,`�:�օ9 �=�����k��Fmg����7���:� %;�v;$��;;��;_��;���;�@�;�m�;T��;�Q�;�A�;~|�;DQ�;�^�;���;1e�;4�;���;~�;��.;���:p%9O��J���¬��%Q��a9�o�:��#;�N`;,�;�{;��T;�8;���:h;ʸ�{����d��^�!�c�9�h�:�KA;�Ӈ;S��;�E�;҉�;$U�;yL�;c��;s/�;.;�;��;�&�;���;�=�;���;�M�;��;)�;@�e;l;�vw:|Q��慺S´�ȩ��G�	�j�:�-�:	O:;�n;�Z�;�r;rbA;Đ�:}�*:޹*薺�ǵ��|���ʢ�-S:��;��\;�w�;�[�;���; 3�;Y�;� �;T�;ݷ�;�-�;��;���;+2�;��;6z�;�'�;���;�;�rJ;�D�:�	:މ��n��gV���'���u]�"�o:��
;��N;�y;7��;,Te;8M+;�߾:C��9�
;�SĨ�|)��2e�A(8�:�n%;�w;�%�;��;��;��;�L�;�r�;ʟ�;�G�;�0�;Ud�;�1�;V8�;�k�;�0�;l��;�G�;�;Q^.;&�:w�9�"R�3ꭺ�t����T�8�	9���:��";	d_;�;��z;��S;�g;��:A��>m~��Ӵ����.$��)�9�-�:��@;I��;�a�;��;)�;���;���;!��;w��;j��;{,�;���;r�;=��;r��;���;���;�;0�d;	�;>�s:E�_��և��Ƕ��ş�*�	:y��:�9;FYm;���;�Sq;<@;�V�:r]&:��ט��  �  f��$?�8�&G:�g�:�P2;зv;^��;eJ�;�k�;c��;� �;�~�;tl�;~��;���;�;p��;\�;|�;y1�;�{�;���;�k�;kh;T�";߾:�
:�� 8������=9V;f:��:�^<;�"w;M�;ر�;]x�;�sX;6�;�N�:���9P�������f�9<9�:@{;��I;�E�;/��;�·;u|�;��;r �;��;���;�/�;u,�;���;C��;pf�;���;���;�չ;���;���;�<R;��;4��:*��96�b���`�)��92>�:6;��R;���;Ԅ�;2��;	P};�YD;� ;�%�:28�9��͸���5�c:���:W�;�a;7��;��;�9�;D��;�}�;���;���;1��;�8�;0]�;���;���;N��;Z��;�0�;I߳;�;p�~;,�:;1��:!`b:�'D9�p�rl88,�":�B�:��&;�:f;���;C��;���;H`l;�b.;���:s9:V�8v�l9�rJ:M��:3;�{w;#�;��;4��;�)�;Q��;���;���;<a�;�/�;Fw�;���;^��;���;���;6ξ;���;x��;q�h;�e#;R�:[:q�!8j��S�F9�h:�W�:	=;.�w;�{�;��;L؅;�3Y;��;5��:S2�90�������9AH�:��;fjJ;eu�;���;=�;���;�;<,�;���;���;&�;�;�~�;��;@�;p�;%��;5��;LC�;���;h�Q;�	;�2�:�q�9$��!B��^��9�u�:8N;r�Q;a4�;C�;TG�;�w|;O�C;& ;�[:G{9�F�h����:࿰:�;�x`;!+�;�9�;�ۼ;�J�;T�;@�;w��;G�;b��;���;�^�;���;�c�;;s�;@��;�q�;;��};i
:;�
�:k�^:��49� ����7:A:~�:P�%;�e;J�;!�; �;>k;�I-;���:5:=r�8�  �  f�:\��:;��:B");ҲY;@(�;Sښ;+<�;��;h��;~}�;�;N%�;��;���;>`�;5��;/��;�`�;'��;���;�̨;�c�;=�;<�N;;@<�:4��:稯:�:�s;�	@;�v;��;y�;��;��;���;��X;��";���:A�:X�:{��:t<;]9;��j;<�;�j�;6;�;��;�!�;�K�;v��;��;�1�;�C�;�N�;�6�;���;���;!��;��;נ�;.��;3�p;�\?;̃;�1�:�=�:鱷:���:f$;o>S;([�;��;�;�s�;��;$8};=�F;�7;~��:�[�:$ĸ:c�:V�;�I;_${;)c�;pR�;��;r~�;r/�;9��;-��;b��;�o�;(�;c��;BN�;7u�;��;ꁺ;sJ�;�m�;�%�;0`;y,/;��;���:s��:|�:���:��.;<xe;5K�;��;��;��;mǎ;܁k;c�4;a�;�?�:6��:���:1R�:��); yZ;n��;�<�;柬;IU�;v
�;���;���;1��;k	�;�m�;W��;j�;o �;���;.Y�;ֶ;X�;���;�6�;ARO;��;8B�:n�:B��:n.�:;��@;�Lw;�g�;�q�;kY�;?s�;R�;�;Y;��#;��:W��:��:״�:�;��9;k;&4�;���;'\�;���;V4�;QW�;���;��;�'�;�2�;�6�;��;���;���;�u�;���;�^�;�s�;	p;�>;!�;A��:0��:��:���:�B;rYR;��;@>�;�y�;J�;�6�;/j|;z
F;~|;]L�:��:�y�:���:m;GBI; }z;�;��;�/�;H�;y��;�O�;Uc�;�;�;���;��;@\�;R��;�;�e�;��;�ܭ;} �;Q��;�)_;tJ.;��;���:��:�p�:���:)�-;hXd;ɸ�;|$�;]N�;��;9�;�mj;�3;ڄ;>]�:�  �  ,}3;��5;�C;Z9X;jq;��;$�;��;�m�;�w�;a0�;>S�;7�;tc�;,��;A��;���;���;�G�;�~�;2[�;:{�;�^�;�;ڼk;,S;�e?;�#4;�5;JrD;�2a;���;h�;�z�;���;���;Hi�;7M�;��;�[q;z�O;�A:;�3;JQ9;��I;��`;��z;*.�;��;�V�;�é;s��;~L�;O�;�#�;���;��;���;���;=Q�;�̳;D�;]��;�a�;R͋;�~;�&d;��L;�m;;?�3;��9; �M;-n;�݊;w��;=}�;�ƶ;;��;Hz�;m�;�6�;+�e;��G;y�6;�+4;F;>;�@Q;kyi;�ǁ;�_�;۩�;���;��;W��;a&�;�y�;m��;d�;�(�;�"�;q��;���;��;��;DL�;���;���;�"u;J�[;��E;�f7;��3;*r>;�W;�z;���;X��;�1�;Zz�;;�;`g�;Eܓ;);*�Z;{}@;>_4;_6;��C; Y;,0r;��;hT�;&�;?զ;��; ��;Z��; ~�;���;H�;��;4'�;i�;���;�ܭ;���;�͚;8��;2�;Hl;�S;6�?;̪4;��5;�E;B�a;=�;�8�;uѩ;Z�;\�;�ů;ͩ�;l�;�r;4�P;)�:;��3;{�9;.ZJ;~9a;}{;l\�;�;cw�;>ݩ;�Ĳ;�W�;��;� �;�z�;��;���;���;)+�;���;T��;�a�;G �;M��;�q};x}c;L;5�:;�3;Ǵ8;"�L;�(m;�l�;�A�;�;W�;�C�;V�;�;EՅ;��d;�F;�6;�3;c�=;ÜP;�h;+r�;g�;�K�;�I�;�|�;VN�;��;��;�@�;���;l��;U��;p(�;!�;ir�;]s�;�ݝ;r3�;�"�;MGt;��Z;R
E;=y6;��2;r=;V;�y;&�;`�;j��;��;ڬ�;5ܥ;AU�;5 ~;e�Y;B�?;�  �  ���;;x;�Ps;&q;�6q;3�s;+�x;F��;cu�;��;��;Sͭ;��;v��;�e�;���;�y�;5ͪ;��;�x�;m��;�e;c>w;��r;q;׌q;YKt;�y;2�;��;#6�;�{�;��;~��;��;IR�;1��;���;⧨;��;��;TO�;� ~;��v;��r;'Yq;V)r;@Wu;j�{;�Z�;8�;B�;}��;Vu�;�z�;���;�.�;R}�;��;���;�;�?�;V�;�};EYv;��r;��q;*s;��v;��};�؄;=�;$�;���;�´;:�;6�;���;-#�;�;^�;��;l��;��;It{;�Yu;wTr;f�q;�/s;�Fw;J�~;���;��;���;���;?��;3V�;?��;�
�;���;ɾ�;L�;�ߔ;��;^�;�?z;m�t;**r;$�q;��s;�^x;�i�;m�;ꑑ;sH�;��;'��;���;~��;:0�;}Ϲ;拭;�ʟ;ޒ;�d�;��;\y;{t;��q;��q;&Lt;miy;�V�;lވ;��; ��;F?�;�Y�;Xr�;Y��;��;��;�9�;Uu�;�ڐ;I��;��;�w;�ss;��q;�r;��t;�z;)U�;�e�;���;�ʢ;Io�;"	�;\H�;R��;�;A�;^�;RN�;<�;���;×~;�&w;�7s;�q;��r;b�u;%�{;�z�;`�;v��;��;�y�;�w�;���;��;[e�;�˳;�y�;C�;,�;��;É|;m�u;yRr;IFq;jgr;@�u;��|;q�;L��;�|�;^�;�R�;î�;"�;�^�;���;��;��;䑖;2,�;�Â;0�z;ȳt;��q;J�p;�r;�v;�6~;���;�4�;b��;F�;1�;�ۿ;HG�;w��;y�;�E�;���;l�;b|�;���;�ey;��s;�Pq;� q;A�r;-vw;��;��;`�;�;ル;��;Y��;Od�;���;�G�;
�;�K�;?d�;,��;�  �  O,�;�I�;��;�o;��V;�B;g5;��3;"�@;i[;O"�;�y�;ɦ;�/�;��;��;��;���;o{w;lT;H�<;N�2;�%7;Z:F;�T\;w�u;��;��;���;e�;�
�;ഹ;���;��;���;��;+�;q��;h�;���;Q%�;��;c��;��;C�;�g;��O;k'=;��3;[7;U�H;Cjg;_2�;�T�;#�;�ӵ;W`�;���;.��;ݑ�; �k;�K;��8;��3;<;��M;��e;��;��;7�;=�;��;�i�;H�;Dx�;��;7��;?��;��;���;���;iY�;�d�;x�;Yv�;̞�;�jy;��_;�I;�9;Ԃ3;C�;;��Q;t;�-�;���;g�;�8�;���;��;D+�;�ւ;�`;2�C;`5;�&5;C�@;�!U;��m;���;�h�;rv�;�M�;&o�;9�;��;^��;�\�;�+�;)��;:8�;T`�;�,�;Fk�;&W�;���;��;�i�;��p;a�W;w�B;[�5;�4;��A;�E\;��;��; @�;��;`�;���;��;�k�;�Qx;�6U;�S=;c�3;#�7;��F;��\;�qv;�1�;N0�;}ʞ;�W�;�U�;0�;* �;i�;�H�;>�;��;K%�;���;O�;�w�;�:�;t*�;͍;�&�;9h;�+P;0�=;74;�@7;��H;�g;]=�;�X�;.�;�ɵ;gO�;���;Ua�;l�;�Wk;YzK;�+8;�N3;W�;;NM;P�d;��~;�)�;��; ס;�!�;���;�|�;&
�;��;���;�(�;G��;�u�;���;���;h�;���;�!�;�J�;��x;+_;�\H;	Q8;ʻ2;Y�:;Q;�+s;���;)'�;(�;���;�;9��;¯�;_^�;�_;�C;d�4;RL4;$@;tJT;
m;���;���;� �;�Ӥ;��;ݶ�;���;��;'��;:��;1�;ͳ�;�߿;���;��;��;�  �  ;a�;s��;ك;��V;��&;ɥ�:|��:)�:��:�;��6;[}m;Yv�;v<�;rG�;l�;W{�;�ba;�+;��:�p�:���:�y�:�A;�1;.b;��;&�;��;\��;M��;c^�;W"�;��;S��;��;�K�;�c�;Z?�;��;p;;h��;�4�;�;�)x;U�F;�
;�:�ȶ:�в:ۈ�:d�;�I;�;}��;���;�n�;���;�ɂ;w�O;};B�:�ߵ:� �:�.�:z�;B;scs;���;Щ�;��;0A�;�b�;�7�;w��;
��;*r�;�Q�;�&�;���;�3�;���;%�;���;.��;��;/h;�7;�W
;t�:��:��:���:UD&;<\;{Z�;�N�;.��;_�;�N�;�ot;��=;�;Is�:�|�:�8�:�c�:H";e<R;f��;U�;��;ʋ�;���;i�;�d�;�C�; ��;t}�;?	�;���;���;ҫ�;#��;�ø;�̫;_%�;>�;}�W;�V';�4�:G�:��:S��:��;5�7;Uln;a��;�;å;o�;��;6Jb;��+;�B�:n��:���:K��:��;��1;Ӣb;�Z�;}l�;�;��;E*�;��;�r�;6��;�1�;�m�;-��;��;H��;���;F�;���;O}�;�N�;G�x;�WG;�o;��:`�:�M�:���:��;��I;��;q~�;���;�]�;�u�;˪�;I�O;��;�u�:b��:� �:��:�0;�fA;��r;���;�H�;6I�;5ٽ;"��;���;��;��;-�;���;[��;p�;C��;���;Ļ;+E�;�2�;���;z�g;pR6;��	;���:}�:�d�:V�:W%;�E[;�ۇ;�͛;0	�;�l�;�Α;zts;9�<;�
;��:ܽ�:���:��:ur!;�eQ;22�;\x�;w��;g�;k^�;_��;���;v��;�f�;D��;k��;9 �;�H�;92�;37�;�S�;�  �  �(�; �;�s;Om.;
!�:^�;:Y��8/���G�8��@:}6�:�1;�Jn;j݋;]�;d�;��a;`";���:j�:��7ay�<�T9�fk:T��:�>;�Ӏ;w%�;P��;^�;u��;���;ا�;v�;2�;���;WB�;:��;�V�;��;���;�/�; #�;[��;�];M�;���:���9:o����ŸJ��9��:�E;D�G;��;��;���;J�;[�N;�;�ؔ:4&�9ڐ�{17�}��9�:�~;V;��;��;hѺ;�_�;���;���;�;���;xP�;0[�;3��;��;:,�;���;�	�;��;TP�;̫�;spF;#
;���:��9lļ��~h�ID:曰:q;/\;��;NN�;6ٍ;Qu;`x9;b�:Ծ\:Ϻ+9�Q�F�8؉(:�Q�:�r';�ul;x`�;�D�;�;��;��;���;(��;}��;�=�;)t�;$��;9��;^l�;*��;R!�;ђ�;�|�;9�s;3/;B��:��>:�i�8j��|��8�zD:�:;2;+Do;�[�;���;t�;��b;��";+��:�:-�7�۸?�_9��m:l��:�>;��;�l�;�ܴ;��;7+�;���;���;���;TW�;p=�;Z��;��;��;DZ�;eJ�;�{�;�j�; ��;�]; 
;�g�:���9v)~��轸#2�9WW�:[;ϛG;h�;��;�;I2�;
�N;��;(�:*��9�.���W�%��9�:*�;�eU;�V�;��;�m�; ��;s��;b0�;ϫ�;�J�;���;g��;b�;Ƥ�;H��;t�;���;���;V��;�U�;��E;�U ;�:(؉9S�ָ[eⷙI�9���:Au;c|[;e�;�ɑ;.U�;�t;wy8;��:��X:�@9>,�z�M8�1%:���:7�&;z�k;Q�;)ӭ;�2�;���;L��;�[�;�q�;��;G��;��;vj�;�p�;��;<_�;۲�;�  �  ���;f5�;�wW;uM;�->:,fŹ� ��9���H
����ʹ#�7:��:��C;"8s;���;Ik;V�5;�>�:���9��Ϋ��Oµ�����l"�DR�:�s;
\i;(��;R�;)��;���;���;�z�;���;>=�;0��;���;���;l�;p��;:��;5�;��;���;e<;Ny�:'��90�.�ߓ���Ͳ�J�r�;3��Ǒ:� ;�sW;R�|;��~;g7];�A;�: ~�8�]�������VjD�
�d9�ȼ:@�3;9�;�6�;]�;�;C��;|}�;�[�;���;I_�;���;���;ϩ�;M_�;��;r�;��;k�;��r;ؕ ;N	�:p��N�o��䱺����R�/���9��:/;k�g;��;��w;#oK;b�;o�^: ����.�����u�\d���:n �:q1O;�ʍ;�5�;&�;N�;]��;�7�;��;
��;G:�;��;z�;o�;k�;=��;���;��;Y��;?X;�;�CA:"��B�����'O��ˡùƑ;:�:�D;�8t;V5�;VHl;j�6;�"�:=9�9��9���@��󨁺O�����:�
;��i;��;:�;���;9�;�B�;���;	�;{��;�C�;�L�;I�;�b�;�<�;��;_�;KK�;��;��<;lV�:���9�v-������S���/r��w*���:8;nmW;:�|;ޘ~;�];};�J�:<{�8ݳ^���������5�F�]�[9@��:3;]��;�ע;C��;3��;#��;��;j��;��;���;��;}�;>H�;� �;n~�;�;�\�;��;8�q;$�;S��:�u$���r�Ҍ��vI��uC3�R>�98��:.;�f;N]�;ّv;SgJ;��;I�Z:�F��> ���O���v�����[�:�z�:V\N;^�;�ū;Ȳ�;j��;S�;̺�;�/�;�z�;��;W�;t��;��;ˎ�;�e�;�v�;�  �  S�;}i�;� A;���:\��8ٕ�c��C�����\��4	U8Gܳ:a�&;�Y;6i;G_Q;�\;Qˍ:�$w������)	����U�8k����9#��:|�T;2��;(L�;c%�;:�;�;���;�Z�;�V�; ��;�Q�;>��;���;qA�;4��;���;!��;��z;��";Z�:���	$��c��7@��亹vI�aJ:*J�:�;;?�c;�1f;�+B;H4�:��*:,&���غ�2�����3̺����Tf:��;�sr;��;���;+��;*D�;9r�;%��;���;0b�;ϓ�;|p�;��;�w�;�,�;��;<Y�;+�;�Q_;_�;1:�~F�C-�
��h�%|��H+���y:@L;�M;si;��^;��.;��:��]9݄��h��/��}��kV����f�w%�:|�7;���;���;��;M"�;��;l��;c��;@6�;�3�;x�;pF�;_��;�D�;�	�;���;���;�Ί;.�A;i�:�=�8mG���� �6(�� �,���f��8ϵ: �';s�Z;�"j;�aR;�Y;O��:|h��Y��;����A�h�6��9W��:X�U;O��;&��;Dn�;���;�j�;m:�;���;���;�A�;��;')�;�C�;��;
�;�̻;P��;�t{;�*#;
�:����w���y�q��R�k�H���:�X�:��;;�c; f;f�A;��:��):ċ'��xٺ���3~��Hͺ�/�)�c:?9;վq;h!�;l)�;��;���;E	�;��;���;���;n-�;��;\��;��;��;���;��;y��;��^;��;SQ:�I�w��4��cJ��X��'�Ĺ�u:�B;wL;�ch;�~];��-;
��:�DN9"��;��N�����I ��ߪ����:��6;��;�'�;a��;���;ȝ�;�q�;��;c��;״�;׆�;��;B�;%��;c��;���;�  �  �ϩ;���;�v8; ��:�������Tf�ZW)�e!�T���޾;���:q;��P;�h`;LH;��;�g:����׺���X(�˳������09P�:�*M;�=�;U�;&��;]�;#��;���;ڽ�;���;��;��;�Z�;���;� �;�o�;
��;�̟;�yt;=;:�Y:�;�έ�����x&�j]�^d���f�9��:$02;�%[;Xh];X�8;��:Q��9[h�YP��OX$��8"�+�BNA��t0: �;�k;�{�;#��;8��;J"�;l;�;w�;:E�;Ӓ�;���;G��;���;)K�;'�;���;9*�;{��;]�W;Η�:���9갅�os��H&��Z��;�9m��D:^k;'D;�`;��U;��$;3\�:!ra��������:1(�ȴ�Y�Ǻ���{�:�.;��;���;�H�;���;���;h��;�;�x�;Ha�;�B�;G��;�j�;5!�;���;.M�;*8�;��;=9;M��:����b�������(�B��Է�D�,���:q;?�Q;Qna;�!I;ʯ;�k:���8ֺ-�
�'���
�M���:94��:�M;��;eJ�;��;�Y�;�A�;���;��;>��;7q�;��;F��;2�;$q�;w��;'�;��;|�t;Ņ;�x[:ɳ������;&��-����O�9'�:�)2;�[;�F];�X8;��:���9p�i�E���$��"��?��C� �-:�3;��j;9�;	,�;')�;���;���;#��;*��;�*�;jb�;si�;}<�;���;���;�6�;�Ҳ;�F�;�(W;R3�:f�9�2���>��'��= �溫U"��@:�`;9C;��_;3�T;>�#;�S�:��z���I��w)�َ��ɺY��,ٗ:��-;k5�;4��;�־;�m�;]|�;
)�;���;M��;���;���;I;�;���;��;wb�;'��;�  �  S�;}i�;� A;���:\��8ٕ�c��C�����\��4	U8Gܳ:a�&;�Y;6i;G_Q;�\;Qˍ:�$w������)	����U�8k����9#��:|�T;2��;(L�;c%�;:�;�;���;�Z�;�V�; ��;�Q�;>��;���;qA�;4��;���;!��;��z;��";Z�:���	$��c��7@��亹vI�aJ:*J�:�;;?�c;�1f;�+B;H4�:��*:,&���غ�2�����3̺����Tf:��;�sr;��;���;+��;*D�;9r�;%��;���;0b�;ϓ�;|p�;��;�w�;�,�;��;<Y�;+�;�Q_;_�;1:�~F�C-�
��h�%|��H+���y:@L;�M;si;��^;��.;��:��]9݄��h��/��}��kV����f�w%�:|�7;���;���;��;M"�;��;l��;c��;@6�;�3�;x�;pF�;_��;�D�;�	�;���;���;�Ί;.�A;i�:�=�8mG���� �6(�� �,���f��8ϵ: �';s�Z;�"j;�aR;�Y;O��:|h��Y��;����A�h�6��9W��:X�U;O��;&��;Dn�;���;�j�;m:�;���;���;�A�;��;')�;�C�;��;
�;�̻;P��;�t{;�*#;
�:����w���y�q��R�k�H���:�X�:��;;�c; f;f�A;��:��):ċ'��xٺ���3~��Hͺ�/�)�c:?9;վq;h!�;l)�;��;���;E	�;��;���;���;n-�;��;\��;��;��;���;��;y��;��^;��;SQ:�I�w��4��cJ��X��'�Ĺ�u:�B;wL;�ch;�~];��-;
��:�DN9"��;��N�����I ��ߪ����:��6;��;�'�;a��;���;ȝ�;�q�;��;c��;״�;׆�;��;B�;%��;c��;���;�  �  ���;f5�;�wW;uM;�->:,fŹ� ��9���H
����ʹ#�7:��:��C;"8s;���;Ik;V�5;�>�:���9��Ϋ��Oµ�����l"�DR�:�s;
\i;(��;R�;)��;���;���;�z�;���;>=�;0��;���;���;l�;p��;:��;5�;��;���;e<;Ny�:'��90�.�ߓ���Ͳ�J�r�;3��Ǒ:� ;�sW;R�|;��~;g7];�A;�: ~�8�]�������VjD�
�d9�ȼ:@�3;9�;�6�;]�;�;C��;|}�;�[�;���;I_�;���;���;ϩ�;M_�;��;r�;��;k�;��r;ؕ ;N	�:p��N�o��䱺����R�/���9��:/;k�g;��;��w;#oK;b�;o�^: ����.�����u�\d���:n �:q1O;�ʍ;�5�;&�;N�;]��;�7�;��;
��;G:�;��;z�;o�;k�;=��;���;��;Y��;?X;�;�CA:"��B�����'O��ˡùƑ;:�:�D;�8t;V5�;VHl;j�6;�"�:=9�9��9���@��󨁺O�����:�
;��i;��;:�;���;9�;�B�;���;	�;{��;�C�;�L�;I�;�b�;�<�;��;_�;KK�;��;��<;lV�:���9�v-������S���/r��w*���:8;nmW;:�|;ޘ~;�];};�J�:<{�8ݳ^���������5�F�]�[9@��:3;]��;�ע;C��;3��;#��;��;j��;��;���;��;}�;>H�;� �;n~�;�;�\�;��;8�q;$�;S��:�u$���r�Ҍ��vI��uC3�R>�98��:.;�f;N]�;ّv;SgJ;��;I�Z:�F��> ���O���v�����[�:�z�:V\N;^�;�ū;Ȳ�;j��;S�;̺�;�/�;�z�;��;W�;t��;��;ˎ�;�e�;�v�;�  �  �(�; �;�s;Om.;
!�:^�;:Y��8/���G�8��@:}6�:�1;�Jn;j݋;]�;d�;��a;`";���:j�:��7ay�<�T9�fk:T��:�>;�Ӏ;w%�;P��;^�;u��;���;ا�;v�;2�;���;WB�;:��;�V�;��;���;�/�; #�;[��;�];M�;���:���9:o����ŸJ��9��:�E;D�G;��;��;���;J�;[�N;�;�ؔ:4&�9ڐ�{17�}��9�:�~;V;��;��;hѺ;�_�;���;���;�;���;xP�;0[�;3��;��;:,�;���;�	�;��;TP�;̫�;spF;#
;���:��9lļ��~h�ID:曰:q;/\;��;NN�;6ٍ;Qu;`x9;b�:Ծ\:Ϻ+9�Q�F�8؉(:�Q�:�r';�ul;x`�;�D�;�;��;��;���;(��;}��;�=�;)t�;$��;9��;^l�;*��;R!�;ђ�;�|�;9�s;3/;B��:��>:�i�8j��|��8�zD:�:;2;+Do;�[�;���;t�;��b;��";+��:�:-�7�۸?�_9��m:l��:�>;��;�l�;�ܴ;��;7+�;���;���;���;TW�;p=�;Z��;��;��;DZ�;eJ�;�{�;�j�; ��;�]; 
;�g�:���9v)~��轸#2�9WW�:[;ϛG;h�;��;�;I2�;
�N;��;(�:*��9�.���W�%��9�:*�;�eU;�V�;��;�m�; ��;s��;b0�;ϫ�;�J�;���;g��;b�;Ƥ�;H��;t�;���;���;V��;�U�;��E;�U ;�:(؉9S�ָ[eⷙI�9���:Au;c|[;e�;�ɑ;.U�;�t;wy8;��:��X:�@9>,�z�M8�1%:���:7�&;z�k;Q�;)ӭ;�2�;���;L��;�[�;�q�;��;G��;��;vj�;�p�;��;<_�;۲�;�  �  ;a�;s��;ك;��V;��&;ɥ�:|��:)�:��:�;��6;[}m;Yv�;v<�;rG�;l�;W{�;�ba;�+;��:�p�:���:�y�:�A;�1;.b;��;&�;��;\��;M��;c^�;W"�;��;S��;��;�K�;�c�;Z?�;��;p;;h��;�4�;�;�)x;U�F;�
;�:�ȶ:�в:ۈ�:d�;�I;�;}��;���;�n�;���;�ɂ;w�O;};B�:�ߵ:� �:�.�:z�;B;scs;���;Щ�;��;0A�;�b�;�7�;w��;
��;*r�;�Q�;�&�;���;�3�;���;%�;���;.��;��;/h;�7;�W
;t�:��:��:���:UD&;<\;{Z�;�N�;.��;_�;�N�;�ot;��=;�;Is�:�|�:�8�:�c�:H";e<R;f��;U�;��;ʋ�;���;i�;�d�;�C�; ��;t}�;?	�;���;���;ҫ�;#��;�ø;�̫;_%�;>�;}�W;�V';�4�:G�:��:S��:��;5�7;Uln;a��;�;å;o�;��;6Jb;��+;�B�:n��:���:K��:��;��1;Ӣb;�Z�;}l�;�;��;E*�;��;�r�;6��;�1�;�m�;-��;��;H��;���;F�;���;O}�;�N�;G�x;�WG;�o;��:`�:�M�:���:��;��I;��;q~�;���;�]�;�u�;˪�;I�O;��;�u�:b��:� �:��:�0;�fA;��r;���;�H�;6I�;5ٽ;"��;���;��;��;-�;���;[��;p�;C��;���;Ļ;+E�;�2�;���;z�g;pR6;��	;���:}�:�d�:V�:W%;�E[;�ۇ;�͛;0	�;�l�;�Α;zts;9�<;�
;��:ܽ�:���:��:ur!;�eQ;22�;\x�;w��;g�;k^�;_��;���;v��;�f�;D��;k��;9 �;�H�;92�;37�;�S�;�  �  O,�;�I�;��;�o;��V;�B;g5;��3;"�@;i[;O"�;�y�;ɦ;�/�;��;��;��;���;o{w;lT;H�<;N�2;�%7;Z:F;�T\;w�u;��;��;���;e�;�
�;ഹ;���;��;���;��;+�;q��;h�;���;Q%�;��;c��;��;C�;�g;��O;k'=;��3;[7;U�H;Cjg;_2�;�T�;#�;�ӵ;W`�;���;.��;ݑ�; �k;�K;��8;��3;<;��M;��e;��;��;7�;=�;��;�i�;H�;Dx�;��;7��;?��;��;���;���;iY�;�d�;x�;Yv�;̞�;�jy;��_;�I;�9;Ԃ3;C�;;��Q;t;�-�;���;g�;�8�;���;��;D+�;�ւ;�`;2�C;`5;�&5;C�@;�!U;��m;���;�h�;rv�;�M�;&o�;9�;��;^��;�\�;�+�;)��;:8�;T`�;�,�;Fk�;&W�;���;��;�i�;��p;a�W;w�B;[�5;�4;��A;�E\;��;��; @�;��;`�;���;��;�k�;�Qx;�6U;�S=;c�3;#�7;��F;��\;�qv;�1�;N0�;}ʞ;�W�;�U�;0�;* �;i�;�H�;>�;��;K%�;���;O�;�w�;�:�;t*�;͍;�&�;9h;�+P;0�=;74;�@7;��H;�g;]=�;�X�;.�;�ɵ;gO�;���;Ua�;l�;�Wk;YzK;�+8;�N3;W�;;NM;P�d;��~;�)�;��; ס;�!�;���;�|�;&
�;��;���;�(�;G��;�u�;���;���;h�;���;�!�;�J�;��x;+_;�\H;	Q8;ʻ2;Y�:;Q;�+s;���;)'�;(�;���;�;9��;¯�;_^�;�_;�C;d�4;RL4;$@;tJT;
m;���;���;� �;�Ӥ;��;ݶ�;���;��;'��;:��;1�;ͳ�;�߿;���;��;��;�  �  ���;;x;�Ps;&q;�6q;3�s;+�x;F��;cu�;��;��;Sͭ;��;v��;�e�;���;�y�;5ͪ;��;�x�;m��;�e;c>w;��r;q;׌q;YKt;�y;2�;��;#6�;�{�;��;~��;��;IR�;1��;���;⧨;��;��;TO�;� ~;��v;��r;'Yq;V)r;@Wu;j�{;�Z�;8�;B�;}��;Vu�;�z�;���;�.�;R}�;��;���;�;�?�;V�;�};EYv;��r;��q;*s;��v;��};�؄;=�;$�;���;�´;:�;6�;���;-#�;�;^�;��;l��;��;It{;�Yu;wTr;f�q;�/s;�Fw;J�~;���;��;���;���;?��;3V�;?��;�
�;���;ɾ�;L�;�ߔ;��;^�;�?z;m�t;**r;$�q;��s;�^x;�i�;m�;ꑑ;sH�;��;'��;���;~��;:0�;}Ϲ;拭;�ʟ;ޒ;�d�;��;\y;{t;��q;��q;&Lt;miy;�V�;lވ;��; ��;F?�;�Y�;Xr�;Y��;��;��;�9�;Uu�;�ڐ;I��;��;�w;�ss;��q;�r;��t;�z;)U�;�e�;���;�ʢ;Io�;"	�;\H�;R��;�;A�;^�;RN�;<�;���;×~;�&w;�7s;�q;��r;b�u;%�{;�z�;`�;v��;��;�y�;�w�;���;��;[e�;�˳;�y�;C�;,�;��;É|;m�u;yRr;IFq;jgr;@�u;��|;q�;L��;�|�;^�;�R�;î�;"�;�^�;���;��;��;䑖;2,�;�Â;0�z;ȳt;��q;J�p;�r;�v;�6~;���;�4�;b��;F�;1�;�ۿ;HG�;w��;y�;�E�;���;l�;b|�;���;�ey;��s;�Pq;� q;A�r;-vw;��;��;`�;�;ル;��;Y��;Od�;���;�G�;
�;�K�;?d�;,��;�  �  ,}3;��5;�C;Z9X;jq;��;$�;��;�m�;�w�;a0�;>S�;7�;tc�;,��;A��;���;���;�G�;�~�;2[�;:{�;�^�;�;ڼk;,S;�e?;�#4;�5;JrD;�2a;���;h�;�z�;���;���;Hi�;7M�;��;�[q;z�O;�A:;�3;JQ9;��I;��`;��z;*.�;��;�V�;�é;s��;~L�;O�;�#�;���;��;���;���;=Q�;�̳;D�;]��;�a�;R͋;�~;�&d;��L;�m;;?�3;��9; �M;-n;�݊;w��;=}�;�ƶ;;��;Hz�;m�;�6�;+�e;��G;y�6;�+4;F;>;�@Q;kyi;�ǁ;�_�;۩�;���;��;W��;a&�;�y�;m��;d�;�(�;�"�;q��;���;��;��;DL�;���;���;�"u;J�[;��E;�f7;��3;*r>;�W;�z;���;X��;�1�;Zz�;;�;`g�;Eܓ;);*�Z;{}@;>_4;_6;��C; Y;,0r;��;hT�;&�;?զ;��; ��;Z��; ~�;���;H�;��;4'�;i�;���;�ܭ;���;�͚;8��;2�;Hl;�S;6�?;̪4;��5;�E;B�a;=�;�8�;uѩ;Z�;\�;�ů;ͩ�;l�;�r;4�P;)�:;��3;{�9;.ZJ;~9a;}{;l\�;�;cw�;>ݩ;�Ĳ;�W�;��;� �;�z�;��;���;���;)+�;���;T��;�a�;G �;M��;�q};x}c;L;5�:;�3;Ǵ8;"�L;�(m;�l�;�A�;�;W�;�C�;V�;�;EՅ;��d;�F;�6;�3;c�=;ÜP;�h;+r�;g�;�K�;�I�;�|�;VN�;��;��;�@�;���;l��;U��;p(�;!�;ir�;]s�;�ݝ;r3�;�"�;MGt;��Z;R
E;=y6;��2;r=;V;�y;&�;`�;j��;��;ڬ�;5ܥ;AU�;5 ~;e�Y;B�?;�  �  f�:\��:;��:B");ҲY;@(�;Sښ;+<�;��;h��;~}�;�;N%�;��;���;>`�;5��;/��;�`�;'��;���;�̨;�c�;=�;<�N;;@<�:4��:稯:�:�s;�	@;�v;��;y�;��;��;���;��X;��";���:A�:X�:{��:t<;]9;��j;<�;�j�;6;�;��;�!�;�K�;v��;��;�1�;�C�;�N�;�6�;���;���;!��;��;נ�;.��;3�p;�\?;̃;�1�:�=�:鱷:���:f$;o>S;([�;��;�;�s�;��;$8};=�F;�7;~��:�[�:$ĸ:c�:V�;�I;_${;)c�;pR�;��;r~�;r/�;9��;-��;b��;�o�;(�;c��;BN�;7u�;��;ꁺ;sJ�;�m�;�%�;0`;y,/;��;���:s��:|�:���:��.;<xe;5K�;��;��;��;mǎ;܁k;c�4;a�;�?�:6��:���:1R�:��); yZ;n��;�<�;柬;IU�;v
�;���;���;1��;k	�;�m�;W��;j�;o �;���;.Y�;ֶ;X�;���;�6�;ARO;��;8B�:n�:B��:n.�:;��@;�Lw;�g�;�q�;kY�;?s�;R�;�;Y;��#;��:W��:��:״�:�;��9;k;&4�;���;'\�;���;V4�;QW�;���;��;�'�;�2�;�6�;��;���;���;�u�;���;�^�;�s�;	p;�>;!�;A��:0��:��:���:�B;rYR;��;@>�;�y�;J�;�6�;/j|;z
F;~|;]L�:��:�y�:���:m;GBI; }z;�;��;�/�;H�;y��;�O�;Uc�;�;�;���;��;@\�;R��;�;�e�;��;�ܭ;} �;Q��;�)_;tJ.;��;���:��:�p�:���:)�-;hXd;ɸ�;|$�;]N�;��;9�;�mj;�3;ڄ;>]�:�  �  f��$?�8�&G:�g�:�P2;зv;^��;eJ�;�k�;c��;� �;�~�;tl�;~��;���;�;p��;\�;|�;y1�;�{�;���;�k�;kh;T�";߾:�
:�� 8������=9V;f:��:�^<;�"w;M�;ر�;]x�;�sX;6�;�N�:���9P�������f�9<9�:@{;��I;�E�;/��;�·;u|�;��;r �;��;���;�/�;u,�;���;C��;pf�;���;���;�չ;���;���;�<R;��;4��:*��96�b���`�)��92>�:6;��R;���;Ԅ�;2��;	P};�YD;� ;�%�:28�9��͸���5�c:���:W�;�a;7��;��;�9�;D��;�}�;���;���;1��;�8�;0]�;���;���;N��;Z��;�0�;I߳;�;p�~;,�:;1��:!`b:�'D9�p�rl88,�":�B�:��&;�:f;���;C��;���;H`l;�b.;���:s9:V�8v�l9�rJ:M��:3;�{w;#�;��;4��;�)�;Q��;���;���;<a�;�/�;Fw�;���;^��;���;���;6ξ;���;x��;q�h;�e#;R�:[:q�!8j��S�F9�h:�W�:	=;.�w;�{�;��;L؅;�3Y;��;5��:S2�90�������9AH�:��;fjJ;eu�;���;=�;���;�;<,�;���;���;&�;�;�~�;��;@�;p�;%��;5��;LC�;���;h�Q;�	;�2�:�q�9$��!B��^��9�u�:8N;r�Q;a4�;C�;TG�;�w|;O�C;& ;�[:G{9�F�h����:࿰:�;�x`;!+�;�9�;�ۼ;�J�;T�;@�;w��;G�;b��;���;�^�;���;�c�;;s�;@��;�q�;;��};i
:;�
�:k�^:��49� ����7:A:~�:P�%;�e;J�;!�; �;>k;�I-;���:5:=r�8�  �  �����9���k��"�O:�;e�[;��;���;EO�;���;d��;d��;���;#N�;���;��;�T�;��;�>�;$�;׿;:b�;|�;��I;C�:�
:S�
�.s��Nf��8G���g��m:7
;c�M;Vx;Z=�;��d;�*;,`�:�օ9 �=�����k��Fmg����7���:� %;�v;$��;;��;_��;���;�@�;�m�;T��;�Q�;�A�;~|�;DQ�;�^�;���;1e�;4�;���;~�;��.;���:p%9O��J���¬��%Q��a9�o�:��#;�N`;,�;�{;��T;�8;���:h;ʸ�{����d��^�!�c�9�h�:�KA;�Ӈ;S��;�E�;҉�;$U�;yL�;c��;s/�;.;�;��;�&�;���;�=�;���;�M�;��;)�;@�e;l;�vw:|Q��慺S´�ȩ��G�	�j�:�-�:	O:;�n;�Z�;�r;rbA;Đ�:}�*:޹*薺�ǵ��|���ʢ�-S:��;��\;�w�;�[�;���; 3�;Y�;� �;T�;ݷ�;�-�;��;���;+2�;��;6z�;�'�;���;�;�rJ;�D�:�	:މ��n��gV���'���u]�"�o:��
;��N;�y;7��;,Te;8M+;�߾:C��9�
;�SĨ�|)��2e�A(8�:�n%;�w;�%�;��;��;��;�L�;�r�;ʟ�;�G�;�0�;Ud�;�1�;V8�;�k�;�0�;l��;�G�;�;Q^.;&�:w�9�"R�3ꭺ�t����T�8�	9���:��";	d_;�;��z;��S;�g;��:A��>m~��Ӵ����.$��)�9�-�:��@;I��;�a�;��;)�;���;���;!��;w��;j��;{,�;���;r�;=��;r��;���;���;�;0�d;	�;>�s:E�_��և��Ƕ��ş�*�	:y��:�9;FYm;���;�Sq;<@;�V�:r]&:��ט��  �  l��^������#;&9��:F;���;ܬ;R{�;��;M��;�,�;4��;�w�;���;���;�C�;��;��;Z<�;n��;���;� �;F�1;�,�:��:����D�?@��	����|��g�9pF�:[�1;"__;�h;!!J;f;��b:T��qDǺX����<qߺ�6��s%:��;�c;��;\��;��;�P�;XQ�;��;9(�;�^�;�G�;��;t��;�]�;���;�.�;`B�;ע�;w�m;m�;әQ:���pҺ���J��FҺb�Ͳ?:��;.zE;�g;c;,!9;��:
b�9*Y�&��ح�j

�F︺o̐���:�!(;[�;鑣;�м;+��;��;l"�;��;v��;^7�;���;���;`�;}l�;7�;{��;�6�;��;V�P;�|�:�l�9�x����Ӄ��y�[���l��l��:Yn;z�T;#pj;�Y;$;S��:�iŶ;���O����O��k��I39��:��F;��;i=�;���;m�;RM�;m��;��;b��;�'�;BA�;&��;���;��;��;��;��;?F�;/]2;�*�:A�	�����8��Ÿ�a���=z��~�9q��:�[2;O`;��h;��J;�);��e:*�ํ�ź`��[
�D޺Փ4�f':'�;y0d;!ؘ;&��;���;d�;Z]�;ο�;�%�;�T�;�6�;���;g�;-7�;L��;���;��;
`�;.m;�;#�N:>o���Ӻ���F����ӺO �<:�;O�D;6�f;D5b;F8;�^�:�&�9T\�R��hW�ˬ
�[*�������ސ:��';4;�;�;�u�;�*�;�C�;���; ��;��;���;+K�;Va�;��;���;X��;�8�;�ɯ;���;��O;<��:�2�9�>|�7������ˉ��Ȭ��C.��6�:<;��S;<i;��W;��";uO�:a:�����v���  �  >?�;ا;,��;���;w��;�A<lM<��<��<��<�<!E<�c<�N<�<�<�<��<܍<-�<6_<�< <)u <p��;c��;TB�;:��;Vu�;���;��;��;b��;�<<�<=\	<]�<�;k�;d��;�ѯ;�y�;4_�;բ�;�A�;��;1X�;0a<c<m�<t�<�w<�X<�l<��<m<m�<D�<�!<�<T^<q�<�e<�c<^�<��;6*�;�1�;H��;=V�;�(�;�Y�;Y��;���;���;�E<�W	<گ<�l<%��;�;Sq�;BӪ;��;lʤ;yt�;u�;��;�U�;
 <��<�0<@�<�<8t<��<�<�<�^<�Q<v&<w�<	�<`a<�<��<��<`y�;��;�|�;���;B�;��;�6�;9��;���;�J�;��<j�	<�0<���;�\�;���;b�;��;k��;G�;��;w�;�a�;�r<b~<�'<#<��<8@<	x<��<�<��<��<b-<s<h�<��<G�<Ǽ<D<�� <'�;;�;��;Eť;���;�F�;���;�%�;���;�g<h;<��	<	<m�;���;�A�;�%�;�ɣ;s��;��;ԁ�;�;���;�w<7v<4�<԰<��<2^<�n<;�<�<5�<�t<�<\<�H<J�<iI<�C<v�<
O�;*��;���;(c�;B��;�¢;�;�?�;|��;���;9<� 	<�y<U8<�:�;���;�;�y�;���;Rw�;6#�;�$�;���;��;��
<��<�<��<X�<�@<�K<��<�<h'<�<��<3�<%�<�*<��<�S<��<P	�;��;3�;;�;Dd�;`�;ʮ�;.0�;I��;���;vE<h	<��<�;��;� �;��;O<�;�  �  �#�;\��;���;6�;y��;��<�,<��<�S<I�<l<��<c <a<lk<n]<V�<�a<��<�<��<7<<��<��;���;��;�\�;cQ�;�y�;�y�;3��;h��;�<T1	<�w
<D< �;��;�a�;��;T6�;_G�;	P�;�V�;�;���;1�<6%<�O<��<;�<�<��<b<z�<˽<+<Z�<�<�<�,<��<�<��	<μ�;I�;�0�;�`�;�<�;��;͢�;M:�;���;��;?�<�t
<��	<f�<���;���;,�;�>�;�ާ;���;b��;IG�;��;� <� <�<Ǟ<�?<�O<
�<"<��<*�<�<
�<��<j_<�<��<DU<�_<�<���;E}�;���;wx�;!ʧ;9A�;OF�;�;��;��;�</�
<cY<� <!��; ��;(]�;GN�;�;B�;Fe�;���;���;��<�]<ø<t�<J.<��<��<�3<�:<'�<@�<��<��<�<*=<+�<]<29<�<���;��;��;#��;���;
®;�ſ;�(�;p�;'�<�]	<�
<�G<�Z�;�k�;��;k\�;*��;v��;̕�;���;�I�;���;��<W8<�_<<+�<��<��<�`<��<��<a<O�<�m<�<�<�<%�<�	<�p�;!��;L��;��;ۨ;戨;)9�;���;rA�; ��;�I<�=
<�	<�<�a�;���;���;K�;���;cW�; ��;���;ܴ�;�v <�<�y<�p<�<�<e�<��<m�<�q<��<2�<m<(<��<�<�<%)<��<���;�
�;�C�;=��;iK�;潪;���;]y�;t�;ӄ�;�q<_�
<f<�` <�7�;�2�;޺;�ԫ;�  �  ���;ν;���;���;:�;��<wa<��<�)<�<I<�<��<@�<�m<�9<�<m�<��<��<c�<��<��<�<��;��;���;��;�·;��;��;�4�;���;w+<�H<�u<q	<i<)e�;�;���;�W�;/θ;��;^�;p��;�� <��<�<o<[�<u�<t�<�K<i<s�<L�<��<�<3�<r<��<��<L�<��<�<���;q��;��;���;�(�;���;D�;IC�;�. <-�<�v<��<@<���;b�;v��;���;WA�;#�;�G�;���;t��;��<�<x:<]�<��<�<P�<�<��<�<�	<%�<�<�D<��<L�<w�<�v<�X	<�F�;՞�; 9�;P��;�R�;&�;���;�&�;��;p<��
<*�<��<�s<�Q�;��;bs�;��;h�;�<�;��;�	�;?��;F*<��<�<R[<<�<	|<�)<l�<�$<�<%l<�I<��<��<��<#�<�<&�<߸<�?�;e��;��;w��;=�;7�;Af�;��;�.�;]V<u<��<V�	<�F<��;�]�;�;릹;��;,`�;���;���;,� <��< <�~<��<Y�<�<�M<	<��<�<�<� <�n<P\<��<B�<��<ԑ<��<�0�;��;E��;:[�;ø;i%�;h��;���;��;��<4@<�<�<�<�;E��;Q2�;;/�;R�;���;���;y9�;�O�;W<.�<�<�e<��<7�<+�<>X<b<+s<��<�`<��<H<Ț<�W<�_<�?<�!	<4��;�,�;q��;��;�Է;���;��;%��;XE�;-(<��
<�<=><�-<���;x�;#��;���;�  �  ,��;z	�;$��;��;*<�4<��<��<��<!�<d�<K<h�<n< <t�<��<�<(H<]<+*< <mH<EI
<�� <۹�;�N�;�B�;��;:��;�5�;���;�<�L<Յ<?�<�<L�<�}�;���;,u�;I��;w��;��;��;BS�;�L<G<'�<N0<Q<��<�<B�<hN<�_<ST<i/<�<�u<��<�-<M�<��<�<3x<���;�D�;�Z�;���;���;n��;*$�;���;;<ީ<^�<<f?<U7<�_�;VP�;��;,�;���;��;��;���;�p	<��<z�<?<:<}�<v<*Y<u�< M<S�<��<{P<�<�$<>�<��<��<QZ<�I<�J�;J��;ݍ�;�Y�;�t�;Ԭ�;'�;� <��<�h<��<c�<��	<�<I�;G:�;92�;�$�;Hw�;���;�,�;F5<tf<�<M<ĺ<�.<�+<2<��<��<@E<��<�'<N�<Tv<F7<�S<a'<�m<�l
<N<#��;��;���;��;���;s��;�4�;�,<2w<��<ĳ<rD<�'<���;P�;���;�B�;Z�;���;�O�;H��;(f<s(<�<�?<�<��<N�<E�<M<&[<L<�#<�<pc<��<�<}<Dx<�<�R<�p�;���;���;�>�;�~�;�; ��;�S�;2<s<Y<��<�<<&��;e��;0��;���;�o�;s��;��;"��;�F	<|<P{<$�<�<]j<��<�"<˽<�<}W<�r<�<��<�<:�<QR<s<o#<F<c��;�7�;m�;���;���;�'�;:}�;���;��<D!<t�<ڞ<��	<r� <<��;I��;��;�  �  �;I��;E �;�/<[ 	<t<n�<ZI<�3<��<Ӄ<y�<Z4<��<�<E�<�W<w<؟<e�<�<��<�<�<7�<8� <4��;��;��;$��;�f�;l�<�]
<��<��<ʣ<��<ap<_M<>!�;�{�;4�;���;Q��;{�;��<Y<
|<�6<�:<��<��<�x<��<�-<��<��<N$<��<�r<&�<��<��<��<�4<�5<�r<X��;R��;$��;8�;���;�;G�<��<_�<ܴ<�N<��<,V<}�<w�;���;�|�;�`�;C��;�/ <��<Γ<�L<sw<��<t�<��<�O<��<�<_�<��<�\<=<i�<� <��<��<�d<uP<��	<l$<���;�)�;��;�9�;��;�� <� <`
<%<��<Wg<�<]�<�<�2�;x��;tv�;7]�;_i�;c<u2	<��<�<c{<�f<K�<4�<�<�i<)�<0�<�<ي<�8<,�<m�<�<��<@�<�B<;�<o� <*��;���;[�;��;��;�$<��
<��<�<��<�!<o�<�x<�u�;F��;�R�;�"�;$��;�M�;ק<<r<��<eI<�I<��<c�<�}<��<3,<��<��<�<ͱ<�`<��<��<mp<i�</<9<�J<*d�;��;53�;:��;$v�;��;iw<��<u<<�<]<I$<\�<˹�;���; &�;��;C��;= <�<�h<� <hI<t�<P�<ʩ<�<	i<'�<�<�<#<��<�s<��<=R<��<�-<�<��	<�<C:�;���;�"�;ú�;��;X� <#�<��<߿<��<�!<r<�<�N<P��;$S�;�  �  ҝ<}�<+�<�%	<4�<n<˵<\�<�<%<��<��<.�<a<+<<<jq< �<w�<��<��<xO<*0<�T<,�<�i<Q<�9<o�<3%<5v<�<�<<J<��<+�<5<�W<Zl	<�o<?"<]�<H<�<m
<��<<<;Q<W�<��<�o<�E<��<Y<C`<<Jd<w�<��<��<=�<"�<*�<Hu<h�
<��<��<�<z/<RG<$	<K�<��<��<��<ר<><,�<G�< <��<�<�;<Z,<�0<��<"<�<�H<�<�<�<��<5�<�-<Ft<�Y<'�<�*<�P<�h<�c<�<,<�<G<
�	<�q<��<��<�<oZ<J�
<��<0[<q�<*<3	<��<�1<+<��<Z�<��<p�<^<uX	<J�<:3<��<��<�?<}J<�3<<��<;M<�r<�6<�<��<&�<�<��<�x<`W<z< <Ќ<�s<�\<��<I<ʛ<�<<D<ɨ<�t<! <�(<n`<<�<�	<��<cH<H�<�i<�#<ֈ
<�<�0<>�<w`<H�<��<�t<�G<@�<GT<X<��<`U<:�<#�<̦<>t<��<�e<P<d�
<�\<ƅ<�<�<8<��<�<F�<�<��<�t<>�<��<n�<��<\i<��<B<q<�<#�<k�<i�<�<�<��<��<<u\<��<�9<�<��<��<*<40<<,<��<n�<yU<<=�	<{8<�<-�<�`<<4`
<`<�<��<g�<%�<�<��<	�
<�<�<�  �  �W<X�<E�<�<z�<��<�<�c<T|<�[<��<��<W-<�<�m<��<ݪ<g
<1G<��<�.<�@<��<��<D�<��<��<�<��<E�<��<}b<*<��<Y%<r<�l<GT<u�<V�<{�<�<c<<��<��<&�<g�<��<2'<��<))<�H<'�<��<�<(f<{<�A<&<�M<��<0o<� <�L<�<�<N<�	<<h[<"<5�<$�<��<F?<�n<3�<<o<% <��<X�<~8<?"<_�<?3<� <��<��<�<�<�^<B;<Q�<�1<U�<��<O�<��<5C<R�<0<_g<L�<!�<�<�)<�<�<S�<��<%<�}<x<L8<�<�n<<
<K�</�<r<CK<�<��<8u<��<B�<�<�<��<��<��<i<�<f�<�< <��<He<R <��<��<��<�><Uy<N<�[<ak<<��<��<B�<��<�%<�<��<�<8�<R<��<lO<(�<m�<�~<g�</<��<2<�_<�<;<��<��<�<t9<��<�4<KQ<T�<f�<?<La<�r<H6<G�<�;<=�<�V<��<�-<��<��<��<|�<N�<s,<@�<�d<l�<mR<N
<�9<�b<�;<��<ur<̭<{
<��<�<�<��<�<��<�<��<o.<�<��<�<ʹ<|e<%r<�f<C<�j<�<<-<.�<�<�x<D�<g�<y�<�<h�<`�<B<�:<5�<+g<�,<?�<�<�j<��<�	<}<�<�9<He<�  �  )�<��<��< }<��<�<�p<I�<s�<�<�4<�:<�<*�<��<Eb<G�<�< "
<��<�N<g�<��<l<q�	<�K<A�<U <i�<�H<�J<v1<k
<5�<�2<�H<��<d<'�<7�<j�<#�<�<q�<��<�i<O�<��<8<��<��<�A<�<.<x3<�<y�<ڗ<��<"�<@�<f<�<�<�<�<.(<$�<�<1
<?�<+�<�<^�<�<D"<�u<�i<E�<�M<�u<�<��<�M<c�<�<1�<PO
<��<�B<��<�T<R�<�	<��<��<KQ<�	<�]<�v<J<��<�h<B/<��<�y<z�<��<�L<߰<I�<b�<�<�%<�<�<��<�C<z<�N<L�<T	<�+<�@<.2<��<��<C<}�<�&	<�<w�<��<8�<0�<l<Gs<?<�!<N<��<�<�S<�U
<�<x}<[�<�<\�< �	<�o<׭<�C<<m<�o<�W<2<��<\<�r<�(<�<^�<Y�<�<�<�7<��<w�<�<r<<?,<��<I�<�I<�	<�<�1<>�<D�<T�<ł<�<�<��<-�<�<Y�<{�<� <;}<ɇ<��<�}<L�<m�<{}<�L<��< B<�6<J�<E<�F<a<d<`"<sZ<��<�<P#
<k�<s<��<!<�<�	<�<�b<�<��<� <:<[�<��</<��<1�<�B<Cm<z�<E<Iy<kK<�`<��<�<B�<c�<v<<-8<X<.�<��<��<�<��<�  �  2 <
r<�<d�<��<f�;��;���;���;z[�;u�<�	<|�<S<ư<-�< q<ox<?$ <���;Z��;1J�;f,�;���;CU<(
<jv<u<��<�l<�<Ty<X�<�)<��<��<w�<,�<�5<$�<f�< �<N/<��<'%<�r<��;�7�;���;�n�;�7�;���;oQ<��<!�<oV<i�<T<3r<�0<�.�;E�;���;&��;g�;b�;�<�<��<��< �<6�<l�<�y<a�<�/<w�<��<>H<'�<��<��<��<�,<�<�?<�<>@<_��;h�;��;�w�;RI�;�.�;��<��<�]<��<z�<a�<�%
<��<H�;5��; g�;�P�;K��;�I<T<�<#<�<�2<�<��<a7<��<�<��<'�<x<e#<��<��<X<V<X�<Q<��<�<���;��;�f�;[�;7��;��<T	<�<܍<��<D�< �<��<6Y <�]�;���;j��;|��;N?�;�{<M
<�<ʘ<��<>�<C�<��<��<R<��<�<�<c�<K^<��<r�<h�<�Q<�<�B<��<*��;�a�;��;H��;�N�;/��;rV<=�<��<�Q<5�<�H<jc<�<)�;=�;���;x�;$�;^�; �<ej<�X<��<6�<�<��<SF<��<��<1�<K�<�<޷<�d<A�<r�<� <}�<�<�
<�<8�;��;i��;��;T��;���;��<8�<�<ş<L�<�k<��	<�<΢�;vW�;���;s��;83�;</�<�m<�<��<��<p�<��<�<�I<��<�<9�<"9<��<�<��<P <�  �  ޯ< d<޹<�y<���;��;���;Ч�;|)�;1��;̠�;we<4
<��<j�<��<xK<ŏ�;���;7s�;f��;��;M��;�+�;���;�<�<��<��<��<_�<��<<m<7]<U(<k�<�K<�<y�<�<��<{L<�*<K�<)��;$��;�0�;	G�;9%�;�q�;��;iJ�;|�<A�<{<z^<�><�<���;��;}��;���;���;���;�0�;���;��<<��<y�<8@<��< m<P�<�/<a<]z<�s<|<7�<�<z<<��<ʳ< �<bn�;�T�;�F�;$��;y�;�n�;���;���;Ş<p�<��<!�<�<�<�2�;���;���;��;��;�p�;@�;g�<�
<��<do<x<�><Ql<��<<M�<�J<��<��<6�<�D<�7<�<2�<ۗ<��<��<� �;��;g��;��;n��;O�;��;�<�B
<y<Q�<�<��<t �;	��;m��;&�;�i�;1�;�}�;�G�;u�<f�<��<�<W�<�<��<�3<F�<��</Q<Y<�t<�3<c�<@<h<?n<:J<Q�<���;K�;NZ�;Qj�;QB�;���;$�;JT�;(�<��<�<GV<}3<��<c�;y��;֖�;�c�;��;��;^��;t��;��<�S<0�<"�<f<��<D:</y<��<H.<JH<�B<��<|�<�<��<K�<[x<K�<�<��;���;���;�b�;��;���;U��;"k�;a<�R<��<F</�
<op<^��;;>�;N�;g��;d��;�;&��;�c<��
<��<�6<�=<?<K/<k�<�<ߎ<�<�u<�<�`<�	<��<�p<�  �  8�<y�<S`<P��;=_�;[��;�9�;:��;��;��;�V�;��;�<��<��<�a
<1�<��;�q�;�1�;6E�;+�;_ǿ;L��;ʈ�;�9�;־	<o�<��<x<b�<f�<#�<<S<5�<4�<�<�<��<�<I�<R<��<W<��<�,�;M6�;$D�;��;�D�;g�;ŀ�;�2�;���;��<�<A<Bn<��;���;h��;k��;Ѹ;���;���;��;���;��<6?<�D<>&<q�<9k<�n<�<��<L�<��<YI<�<��<q�<�<pI<3�<�<� <ew�;Hq�;D��;uθ;(�;���;o��;���;��<��	<��<�@<��<4�;�O�;�l�;_��;,�;ދ�;	 �;\D�;^��;[_<�1<P3<~<�<��<U�<2<`<@�<�;<�<^Q<t�<M�<�B<�<�<ؒ<OK�;:��;\�;���;�	�;n��;Ad�;��;3��;L�<i�<��<��
<6�<%��;��;��;���;�e�;��;�9�;���;Ӆ�;��	<��<��<��<r�<?"<��<�z<L�<��<��< �<u"<!7<c�<|u<�<�><S�<�`�;e�;!m�;��;qa�; +�;���;�<�;Ъ�;�<-�<�8<�b<O��;���;)��;�z�;t��;Y��;z��;���;���;��<�<�<>�<��<�9<Q<<W�<ɴ<�<��<�<�P<�<{<��<�<��<��
<���;�;~�;K/�;�f�;���;�p�;T�;Ą�;
�<�	<�w<� <v�<
��;.��;���;�;�;Y��;��;���;���;�<�;�)<2�<W�<�<;�<��<�Y<��<�!<�g<��<�<�<eb< �<v<�  �  P5<��<��<��;���;�ݼ;5�;��;�n�;���;��;m��;�� <�^<Ζ
<!<�i�;)�;9.�;Ƿ;aO�;~�;;ɯ;���;���;h�;v�<�<nr<9�<��<�<wR<j�<��<Շ<v�<K<m�<�J<| <�V<�-<�z<���;�i�;���;�޶;w�;�;	�;n<�;Q;�;���;�<��	<�;
<_�<؈�;Y �;���;Ϧ�;z��;D�;c6�;>p�;9��;(+�;x
<��<<=A<p�<-h<��<&<�<��<��<,-<��<��<��<G"< �<D�<oL�;���;�K�;U��;F�;�ܩ;<C�;���;���;э�;��<ֻ
<�$	<�9<��;6��;/��;%�;���;�>�;:�;j�;��;M�<2�<?�<�!<D<G <�p<x�<}<��<�T<�\<�<��<�9<�h<�i<��<<�y�;|1�;�B�;ij�;ֈ�;Eܬ;�j�;S�;��;9+<��<,�
<�]<���;ޏ�;u��;1�;ͳ�;�ܧ;_"�;���;o��;�X�;��<v�<��<��<�
<�8<y<��<�<
�<��<7=<�<2q<TE<�y< O<��<���;��;	 �;��;O;�;��;���;�L�;E�;���;�<��	<�3
<��<qk�;���;Ϩ�;fv�;�T�;�B�;6��;�(�;_o�;v��;nM
<�_<K�<<y<6<#a<��<�<�<�b<��<K�<��<�<h�<V�<Y�<��;�l�;��;�R�;�ݧ;�n�;�е;p��;�R�;��;�i<^{
<��<D�<.Q�;OY�;�7�;���;�&�;zѫ;ح�;���;��;��<ȗ<��<�<�	<��<4<�g<A<e< <) <��<5�<�<S2<�  �  ��<��<Ў<�s�;D8�;���;�2�;�;�;cݦ;	�;q�;;B�;�)�;�7<�|	<g�<ݕ�;C��;g��;B��;���;��;�;�O�;�*�;;��;+T<��<��<MP<��<��<`�<4<k%<*�<	<ǅ<t|<q�<��<s�<w�<Vt
<���;�s�;���;[S�;C6�;��;�}�;���;[�;���;)�<��<@	<�<�;W�;�9�;�T�;���;���;{��;�{�;���;Z�;'f	<��<�<��<1T<O�<�<�r<<84<��<&�<Ɛ<��<E�<ӡ<J�<��<���;���;\,�;~�;m^�;�%�;P�;���;�1�;��;�v<�	<7<�� <��;���;�ҹ;]��;��;g�;ѭ�;��;W��;�X<��<�#<�<��<�<��<<y�<d�<�<��<A�<�e<��<b<,�<�<"�<O��;:��;��;��;쥡;�J�;-z�;���;���;���;Ju<4�	<f/<{�;^
�;I�;��;u�; ��;�d�;K��;�z�;���;Iy<@<�<�t<��<H�<��<l,<5M<I�<71<��<��<�<B�<�	<��<G�
<��;��;="�;|�;Y�;J5�;b��;Ҝ�;�d�;���;��<��<	<s�<�a�;43�;k�;u$�;R��;)]�;]Z�;24�;�]�;���;$;	<��<+y<��<�"<Q�<x�<O@<�<�<2�<�y<`b</n<�w<�u<��<��<v��;x%�;�̾;���;���;з�;t��;��;k��;�*�;�6<r`	<��<%� <��;�J�;\�;/�;H�;���;|B�;�Q�;8[�;*#<E�<u�<W�<��<�i<3�<��<��<��<�_<6�<:l<,<�<O�<�  �  P5<��<��<��;���;�ݼ;5�;��;�n�;���;��;m��;�� <�^<Ζ
<!<�i�;)�;9.�;Ƿ;aO�;~�;;ɯ;���;���;h�;v�<�<nr<9�<��<�<wR<j�<��<Շ<v�<K<m�<�J<| <�V<�-<�z<���;�i�;���;�޶;w�;�;	�;n<�;Q;�;���;�<��	<�;
<_�<؈�;Y �;���;Ϧ�;z��;D�;c6�;>p�;9��;(+�;x
<��<<=A<p�<-h<��<&<�<��<��<,-<��<��<��<G"< �<D�<oL�;���;�K�;U��;F�;�ܩ;<C�;���;���;э�;��<ֻ
<�$	<�9<��;6��;/��;%�;���;�>�;:�;j�;��;M�<2�<?�<�!<D<G <�p<x�<}<��<�T<�\<�<��<�9<�h<�i<��<<�y�;|1�;�B�;ij�;ֈ�;Eܬ;�j�;S�;��;9+<��<,�
<�]<���;ޏ�;u��;1�;ͳ�;�ܧ;_"�;���;o��;�X�;��<v�<��<��<�
<�8<y<��<�<
�<��<7=<�<2q<TE<�y< O<��<���;��;	 �;��;O;�;��;���;�L�;E�;���;�<��	<�3
<��<qk�;���;Ϩ�;fv�;�T�;�B�;6��;�(�;_o�;v��;nM
<�_<K�<<y<6<#a<��<�<�<�b<��<K�<��<�<h�<V�<Y�<��;�l�;��;�R�;�ݧ;�n�;�е;p��;�R�;��;�i<^{
<��<D�<.Q�;OY�;�7�;���;�&�;zѫ;ح�;���;��;��<ȗ<��<�<�	<��<4<�g<A<e< <) <��<5�<�<S2<�  �  8�<y�<S`<P��;=_�;[��;�9�;:��;��;��;�V�;��;�<��<��<�a
<1�<��;�q�;�1�;6E�;+�;_ǿ;L��;ʈ�;�9�;־	<o�<��<x<b�<f�<#�<<S<5�<4�<�<�<��<�<I�<R<��<W<��<�,�;M6�;$D�;��;�D�;g�;ŀ�;�2�;���;��<�<A<Bn<��;���;h��;k��;Ѹ;���;���;��;���;��<6?<�D<>&<q�<9k<�n<�<��<L�<��<YI<�<��<q�<�<pI<3�<�<� <ew�;Hq�;D��;uθ;(�;���;o��;���;��<��	<��<�@<��<4�;�O�;�l�;_��;,�;ދ�;	 �;\D�;^��;[_<�1<P3<~<�<��<U�<2<`<@�<�;<�<^Q<t�<M�<�B<�<�<ؒ<OK�;:��;\�;���;�	�;n��;Ad�;��;3��;L�<i�<��<��
<6�<%��;��;��;���;�e�;��;�9�;���;Ӆ�;��	<��<��<��<r�<?"<��<�z<L�<��<��< �<u"<!7<c�<|u<�<�><S�<�`�;e�;!m�;��;qa�; +�;���;�<�;Ъ�;�<-�<�8<�b<O��;���;)��;�z�;t��;Y��;z��;���;���;��<�<�<>�<��<�9<Q<<W�<ɴ<�<��<�<�P<�<{<��<�<��<��
<���;�;~�;K/�;�f�;���;�p�;T�;Ą�;
�<�	<�w<� <v�<
��;.��;���;�;�;Y��;��;���;���;�<�;�)<2�<W�<�<;�<��<�Y<��<�!<�g<��<�<�<eb< �<v<�  �  ޯ< d<޹<�y<���;��;���;Ч�;|)�;1��;̠�;we<4
<��<j�<��<xK<ŏ�;���;7s�;f��;��;M��;�+�;���;�<�<��<��<��<_�<��<<m<7]<U(<k�<�K<�<y�<�<��<{L<�*<K�<)��;$��;�0�;	G�;9%�;�q�;��;iJ�;|�<A�<{<z^<�><�<���;��;}��;���;���;���;�0�;���;��<<��<y�<8@<��< m<P�<�/<a<]z<�s<|<7�<�<z<<��<ʳ< �<bn�;�T�;�F�;$��;y�;�n�;���;���;Ş<p�<��<!�<�<�<�2�;���;���;��;��;�p�;@�;g�<�
<��<do<x<�><Ql<��<<M�<�J<��<��<6�<�D<�7<�<2�<ۗ<��<��<� �;��;g��;��;n��;O�;��;�<�B
<y<Q�<�<��<t �;	��;m��;&�;�i�;1�;�}�;�G�;u�<f�<��<�<W�<�<��<�3<F�<��</Q<Y<�t<�3<c�<@<h<?n<:J<Q�<���;K�;NZ�;Qj�;QB�;���;$�;JT�;(�<��<�<GV<}3<��<c�;y��;֖�;�c�;��;��;^��;t��;��<�S<0�<"�<f<��<D:</y<��<H.<JH<�B<��<|�<�<��<K�<[x<K�<�<��;���;���;�b�;��;���;U��;"k�;a<�R<��<F</�
<op<^��;;>�;N�;g��;d��;�;&��;�c<��
<��<�6<�=<?<K/<k�<�<ߎ<�<�u<�<�`<�	<��<�p<�  �  2 <
r<�<d�<��<f�;��;���;���;z[�;u�<�	<|�<S<ư<-�< q<ox<?$ <���;Z��;1J�;f,�;���;CU<(
<jv<u<��<�l<�<Ty<X�<�)<��<��<w�<,�<�5<$�<f�< �<N/<��<'%<�r<��;�7�;���;�n�;�7�;���;oQ<��<!�<oV<i�<T<3r<�0<�.�;E�;���;&��;g�;b�;�<�<��<��< �<6�<l�<�y<a�<�/<w�<��<>H<'�<��<��<��<�,<�<�?<�<>@<_��;h�;��;�w�;RI�;�.�;��<��<�]<��<z�<a�<�%
<��<H�;5��; g�;�P�;K��;�I<T<�<#<�<�2<�<��<a7<��<�<��<'�<x<e#<��<��<X<V<X�<Q<��<�<���;��;�f�;[�;7��;��<T	<�<܍<��<D�< �<��<6Y <�]�;���;j��;|��;N?�;�{<M
<�<ʘ<��<>�<C�<��<��<R<��<�<�<c�<K^<��<r�<h�<�Q<�<�B<��<*��;�a�;��;H��;�N�;/��;rV<=�<��<�Q<5�<�H<jc<�<)�;=�;���;x�;$�;^�; �<ej<�X<��<6�<�<��<SF<��<��<1�<K�<�<޷<�d<A�<r�<� <}�<�<�
<�<8�;��;i��;��;T��;���;��<8�<�<ş<L�<�k<��	<�<΢�;vW�;���;s��;83�;</�<�m<�<��<��<p�<��<�<�I<��<�<9�<"9<��<�<��<P <�  �  )�<��<��< }<��<�<�p<I�<s�<�<�4<�:<�<*�<��<Eb<G�<�< "
<��<�N<g�<��<l<q�	<�K<A�<U <i�<�H<�J<v1<k
<5�<�2<�H<��<d<'�<7�<j�<#�<�<q�<��<�i<O�<��<8<��<��<�A<�<.<x3<�<y�<ڗ<��<"�<@�<f<�<�<�<�<.(<$�<�<1
<?�<+�<�<^�<�<D"<�u<�i<E�<�M<�u<�<��<�M<c�<�<1�<PO
<��<�B<��<�T<R�<�	<��<��<KQ<�	<�]<�v<J<��<�h<B/<��<�y<z�<��<�L<߰<I�<b�<�<�%<�<�<��<�C<z<�N<L�<T	<�+<�@<.2<��<��<C<}�<�&	<�<w�<��<8�<0�<l<Gs<?<�!<N<��<�<�S<�U
<�<x}<[�<�<\�< �	<�o<׭<�C<<m<�o<�W<2<��<\<�r<�(<�<^�<Y�<�<�<�7<��<w�<�<r<<?,<��<I�<�I<�	<�<�1<>�<D�<T�<ł<�<�<��<-�<�<Y�<{�<� <;}<ɇ<��<�}<L�<m�<{}<�L<��< B<�6<J�<E<�F<a<d<`"<sZ<��<�<P#
<k�<s<��<!<�<�	<�<�b<�<��<� <:<[�<��</<��<1�<�B<Cm<z�<E<Iy<kK<�`<��<�<B�<c�<v<<-8<X<.�<��<��<�<��<�  �  �W<X�<E�<�<z�<��<�<�c<T|<�[<��<��<W-<�<�m<��<ݪ<g
<1G<��<�.<�@<��<��<D�<��<��<�<��<E�<��<}b<*<��<Y%<r<�l<GT<u�<V�<{�<�<c<<��<��<&�<g�<��<2'<��<))<�H<'�<��<�<(f<{<�A<&<�M<��<0o<� <�L<�<�<N<�	<<h[<"<5�<$�<��<F?<�n<3�<<o<% <��<X�<~8<?"<_�<?3<� <��<��<�<�<�^<B;<Q�<�1<U�<��<O�<��<5C<R�<0<_g<L�<!�<�<�)<�<�<S�<��<%<�}<x<L8<�<�n<<
<K�</�<r<CK<�<��<8u<��<B�<�<�<��<��<��<i<�<f�<�< <��<He<R <��<��<��<�><Uy<N<�[<ak<<��<��<B�<��<�%<�<��<�<8�<R<��<lO<(�<m�<�~<g�</<��<2<�_<�<;<��<��<�<t9<��<�4<KQ<T�<f�<?<La<�r<H6<G�<�;<=�<�V<��<�-<��<��<��<|�<N�<s,<@�<�d<l�<mR<N
<�9<�b<�;<��<ur<̭<{
<��<�<�<��<�<��<�<��<o.<�<��<�<ʹ<|e<%r<�f<C<�j<�<<-<.�<�<�x<D�<g�<y�<�<h�<`�<B<�:<5�<+g<�,<?�<�<�j<��<�	<}<�<�9<He<�  �  ҝ<}�<+�<�%	<4�<n<˵<\�<�<%<��<��<.�<a<+<<<jq< �<w�<��<��<xO<*0<�T<,�<�i<Q<�9<o�<3%<5v<�<�<<J<��<+�<5<�W<Zl	<�o<?"<]�<H<�<m
<��<<<;Q<W�<��<�o<�E<��<Y<C`<<Jd<w�<��<��<=�<"�<*�<Hu<h�
<��<��<�<z/<RG<$	<K�<��<��<��<ר<><,�<G�< <��<�<�;<Z,<�0<��<"<�<�H<�<�<�<��<5�<�-<Ft<�Y<'�<�*<�P<�h<�c<�<,<�<G<
�	<�q<��<��<�<oZ<J�
<��<0[<q�<*<3	<��<�1<+<��<Z�<��<p�<^<uX	<J�<:3<��<��<�?<}J<�3<<��<;M<�r<�6<�<��<&�<�<��<�x<`W<z< <Ќ<�s<�\<��<I<ʛ<�<<D<ɨ<�t<! <�(<n`<<�<�	<��<cH<H�<�i<�#<ֈ
<�<�0<>�<w`<H�<��<�t<�G<@�<GT<X<��<`U<:�<#�<̦<>t<��<�e<P<d�
<�\<ƅ<�<�<8<��<�<F�<�<��<�t<>�<��<n�<��<\i<��<B<q<�<#�<k�<i�<�<�<��<��<<u\<��<�9<�<��<��<*<40<<,<��<n�<yU<<=�	<{8<�<-�<�`<<4`
<`<�<��<g�<%�<�<��<	�
<�<�<�  �  �;I��;E �;�/<[ 	<t<n�<ZI<�3<��<Ӄ<y�<Z4<��<�<E�<�W<w<؟<e�<�<��<�<�<7�<8� <4��;��;��;$��;�f�;l�<�]
<��<��<ʣ<��<ap<_M<>!�;�{�;4�;���;Q��;{�;��<Y<
|<�6<�:<��<��<�x<��<�-<��<��<N$<��<�r<&�<��<��<��<�4<�5<�r<X��;R��;$��;8�;���;�;G�<��<_�<ܴ<�N<��<,V<}�<w�;���;�|�;�`�;C��;�/ <��<Γ<�L<sw<��<t�<��<�O<��<�<_�<��<�\<=<i�<� <��<��<�d<uP<��	<l$<���;�)�;��;�9�;��;�� <� <`
<%<��<Wg<�<]�<�<�2�;x��;tv�;7]�;_i�;c<u2	<��<�<c{<�f<K�<4�<�<�i<)�<0�<�<ي<�8<,�<m�<�<��<@�<�B<;�<o� <*��;���;[�;��;��;�$<��
<��<�<��<�!<o�<�x<�u�;F��;�R�;�"�;$��;�M�;ק<<r<��<eI<�I<��<c�<�}<��<3,<��<��<�<ͱ<�`<��<��<mp<i�</<9<�J<*d�;��;53�;:��;$v�;��;iw<��<u<<�<]<I$<\�<˹�;���; &�;��;C��;= <�<�h<� <hI<t�<P�<ʩ<�<	i<'�<�<�<#<��<�s<��<=R<��<�-<�<��	<�<C:�;���;�"�;ú�;��;X� <#�<��<߿<��<�!<r<�<�N<P��;$S�;�  �  ,��;z	�;$��;��;*<�4<��<��<��<!�<d�<K<h�<n< <t�<��<�<(H<]<+*< <mH<EI
<�� <۹�;�N�;�B�;��;:��;�5�;���;�<�L<Յ<?�<�<L�<�}�;���;,u�;I��;w��;��;��;BS�;�L<G<'�<N0<Q<��<�<B�<hN<�_<ST<i/<�<�u<��<�-<M�<��<�<3x<���;�D�;�Z�;���;���;n��;*$�;���;;<ީ<^�<<f?<U7<�_�;VP�;��;,�;���;��;��;���;�p	<��<z�<?<:<}�<v<*Y<u�< M<S�<��<{P<�<�$<>�<��<��<QZ<�I<�J�;J��;ݍ�;�Y�;�t�;Ԭ�;'�;� <��<�h<��<c�<��	<�<I�;G:�;92�;�$�;Hw�;���;�,�;F5<tf<�<M<ĺ<�.<�+<2<��<��<@E<��<�'<N�<Tv<F7<�S<a'<�m<�l
<N<#��;��;���;��;���;s��;�4�;�,<2w<��<ĳ<rD<�'<���;P�;���;�B�;Z�;���;�O�;H��;(f<s(<�<�?<�<��<N�<E�<M<&[<L<�#<�<pc<��<�<}<Dx<�<�R<�p�;���;���;�>�;�~�;�; ��;�S�;2<s<Y<��<�<<&��;e��;0��;���;�o�;s��;��;"��;�F	<|<P{<$�<�<]j<��<�"<˽<�<}W<�r<�<��<�<:�<QR<s<o#<F<c��;�7�;m�;���;���;�'�;:}�;���;��<D!<t�<ڞ<��	<r� <<��;I��;��;�  �  ���;ν;���;���;:�;��<wa<��<�)<�<I<�<��<@�<�m<�9<�<m�<��<��<c�<��<��<�<��;��;���;��;�·;��;��;�4�;���;w+<�H<�u<q	<i<)e�;�;���;�W�;/θ;��;^�;p��;�� <��<�<o<[�<u�<t�<�K<i<s�<L�<��<�<3�<r<��<��<L�<��<�<���;q��;��;���;�(�;���;D�;IC�;�. <-�<�v<��<@<���;b�;v��;���;WA�;#�;�G�;���;t��;��<�<x:<]�<��<�<P�<�<��<�<�	<%�<�<�D<��<L�<w�<�v<�X	<�F�;՞�; 9�;P��;�R�;&�;���;�&�;��;p<��
<*�<��<�s<�Q�;��;bs�;��;h�;�<�;��;�	�;?��;F*<��<�<R[<<�<	|<�)<l�<�$<�<%l<�I<��<��<��<#�<�<&�<߸<�?�;e��;��;w��;=�;7�;Af�;��;�.�;]V<u<��<V�	<�F<��;�]�;�;릹;��;,`�;���;���;,� <��< <�~<��<Y�<�<�M<	<��<�<�<� <�n<P\<��<B�<��<ԑ<��<�0�;��;E��;:[�;ø;i%�;h��;���;��;��<4@<�<�<�<�;E��;Q2�;;/�;R�;���;���;y9�;�O�;W<.�<�<�e<��<7�<+�<>X<b<+s<��<�`<��<H<Ț<�W<�_<�?<�!	<4��;�,�;q��;��;�Է;���;��;%��;XE�;-(<��
<�<=><�-<���;x�;#��;���;�  �  �#�;\��;���;6�;y��;��<�,<��<�S<I�<l<��<c <a<lk<n]<V�<�a<��<�<��<7<<��<��;���;��;�\�;cQ�;�y�;�y�;3��;h��;�<T1	<�w
<D< �;��;�a�;��;T6�;_G�;	P�;�V�;�;���;1�<6%<�O<��<;�<�<��<b<z�<˽<+<Z�<�<�<�,<��<�<��	<μ�;I�;�0�;�`�;�<�;��;͢�;M:�;���;��;?�<�t
<��	<f�<���;���;,�;�>�;�ާ;���;b��;IG�;��;� <� <�<Ǟ<�?<�O<
�<"<��<*�<�<
�<��<j_<�<��<DU<�_<�<���;E}�;���;wx�;!ʧ;9A�;OF�;�;��;��;�</�
<cY<� <!��; ��;(]�;GN�;�;B�;Fe�;���;���;��<�]<ø<t�<J.<��<��<�3<�:<'�<@�<��<��<�<*=<+�<]<29<�<���;��;��;#��;���;
®;�ſ;�(�;p�;'�<�]	<�
<�G<�Z�;�k�;��;k\�;*��;v��;̕�;���;�I�;���;��<W8<�_<<+�<��<��<�`<��<��<a<O�<�m<�<�<�<%�<�	<�p�;!��;L��;��;ۨ;戨;)9�;���;rA�; ��;�I<�=
<�	<�<�a�;���;���;K�;���;cW�; ��;���;ܴ�;�v <�<�y<�p<�<�<e�<��<m�<�q<��<2�<m<(<��<�<�<%)<��<���;�
�;�C�;=��;iK�;潪;���;]y�;t�;ӄ�;�q<_�
<f<�` <�7�;�2�;޺;�ԫ;�  �  ��<؝<pn<3%<\�,<��3<�8<�N;<��;< �9<�j6<î2<�T/<�-<Vo,<�w-<� 0<��3<[77<�7:<��;<��:<�7<�+2<+<ɝ#<21<��<��<��<��<Q�%<_@-<ı3<�7<��8<�5<$X0<M")<ܾ!<�<'E<�<
<u� <��'<�;/<��5<��9<7�;<�9;<g�8<�S5<�1<�.<.�,<��,<nW.<�G1<]�4<��8<R;<��;<\:<@Q6<2$0<��(<�!<�<zg<�B<,_<,,!<�|(<�/<��5<I�8<�.8<�w4<�9.<.�&<��<O\<*�<�<��<��"<Z`*<��1<*^7<y�:<��;<��:<��7<�4<��0<��-<u�,<N&-<:/<x|2<w86<=�9<s�;<��;<D9<�o4<��-<�<&<�S<�?<��<j�<K<9}#<��*<(�1<��6<l�8<�I7<�2<��+<�J$<��<}7<��<��<��<�f%<��,<^�3<?�8<�;<�;<��9<��6<�2<'�/<�J-<�,<��-<00<��3<�c7< b:<�;<�;<��7<�O2<�1+<�#<8S<S<��<�<'�<�%<nh-<��3<�7<�8<�6<��0<�K)<[�!<��<9j<�0<}*<9� <��'<�S/<��5<� :<��;<3E;<��8<�X5<��1<s�.<x�,<��,<:L.<B91<��4<�s8<];<��;<>:<006<B 0<8�(<�[!<:�<v9<�<�-<=� <�H(<��/<�\5<-`8<j�7<�E4<�.<��&<�y<�/<��<�<!�<\�"<�6*<Ln1<�27<�:<۲;<3v:<(�7<��3<�Y0<c�-<Zv,<��,<Q/<�E2<�6<�W9<.d;<�q;<�9<�84<؁-<�&<�<�<�<Ū<��<9:#<��*<�1<M�6<�8<>7<�Z2<�+<$<f<�<�  �  nV<K<1  <Ò&<��-<!j4<�D9<��;<��;<:<n�6<;M3<N
0<&�-<�:-<�;.<P�0<�4<�7<Y�:<�<<Ot;<<e8< 3<1=,<�	%<9�<��<�a<uP<E <��&<,.<TO4<48<B�8<f6<<1<�*<f�"<B+<I�<��<�<�$"<�)<+D0<c6<e�:<�9<<��;<
N9<��5<]H2<6S/<��-<��-<�/<��1<�5<49<��;<�Z<<E�:<'7<�$1<#	*<�#<Y<�<��<�<�m"<W~)<��0<\6<�9<��8<5<�	/<Z�'<�� <��<�<Q�<f\< m$<�+<�2<�8<�f;<:S<<�;<6J8<��4<a<1<�.<�w-<�-<�/<�3<u�6<T:<:
<<�!<<��9<�C5<3�.<̕'<�� <�<�<$�<�n<��$<��+<l�2<vk7<�B9< �7<�F3<��,<Vp%<< �<w�<��<E5 <S�&<+.<՛4<-v9<-�;<$<<DN:<�$7<�3<�<0<c.<ll-<dl.<��0<J4<��7<��:<�E<<�;<R�8<�93<�_,<,%<N�<��<��<�t<�D <g '<0?.<tx4<^8<�9<��6<�>1<}F*<�!#<$R<J<��<k�<dB"<�1)<"\0<	x6<;�:<vH<<�;<QV9<��5<)J2<�Q/<��-<ƅ-<�
/<X�1<Et5<f�8<�t;<�?<<2�:<�6<� 1<w�)<Z�"<b-<��<�<}�<�:"<�J)<LZ0<��5<��8<Yp8<��4<��.<٤'<�� <d�<�l<V<�2<�C$<yl+<�_2<K�7<�9;<�$<<��:<�8<��4<�1<zo.<�A-<R�-<*�/<��2<��6<��9<��;<>�;<�9<5<��.<]'<�� <8�<ed<�A<t-<�f$<��+<z\2<'&7<��8<��7<�3<�q,<�0%<��<؎<�  �  �<8�<{X$<JS*<��0<�6<��:<��<<��<<�<;<qL8<N�4<��1<Y
0<�v/</]0<��2<c�5<9<��;<�+=<��<<E:<4}5<k/<V�(<S=#<�]<�<$�<�#<p�)<e0<+�5<�j9<L:<��7<d3<z�,<$m&<�F!<at<�|<L!<�O&<:�,<�3<\c8<��;<dV=<�<<s~:<^U7<
4<�\1<G�/<��/<&1</�3<17<�;:<�<<�r=<+K<</�8<��3<4w-<L'<�!<)�<�}<g!<.�%<�I,<~�2<)�7<):<�9<��6<0C1<��*<�$<�* <A<]<<%�"<ue(<��.<�5<��9<�<<�d=<�,<<��9<�B6<=3<��0<O�/<�0<��1<�4<�$8<�*;<+=<DJ=<.i;<l7<��1< B+<�*%<ݔ <#]<��<0h"<�'<�s.<]{4<��8<h`:<�9</5<D*/<��(<��"<@;<�G<�1 <r�$<̆*<O1<��6<;<q,=<U0=<�n;<�~8<'5<�02<�<0<٨/<�0<�2<�5<�19<��;<�T=<��<<�B:<8�5<	�/<�)<�_#<-�<4<[�<h$<*<��0<!6<��9<�>:<�7<v=3<��,<V�&<�m!</�<"�<Dl!<wm&<�,<�3<4x8<{ <<e=<��<<��:<aZ7<�4<t[1<��/<��/<�1<Ŭ3<��6<�&:<��<<�W=<(-<<:�8<�3<�P-<"�&<t�!<]�<�M<� <��%<V,<ll2< d7<+�9<�9<pt6<X1<_�*<x$<�<�<	<g�"<�;(<��.<4�4<L�9<�<<�5=<��;<�\9<N6<t�2<ċ0<�|/<��/<x�1<�4<��7<�:<��<<�=<�2;<*57<�1<�	+<��$<EY <�<��<J'"<��'<�/.<�64<�y8<�:<��8<Q�4<��.<�f(<��"<= <�  �  O�$<��&<�|*<({/<��4<Jj9<�<<�+><��=<�h<<��9<27<2�4<0&3<��2<�g3<E/5<T�7<f�:<��<<�-><S�=<<<�8</�3<W.<8�)<2&<�$<H&<2])<�=.<Ǝ3<�8< �:<,z;<��9<+�5<��0<�k+<fK'<�&%<�c%<��'<v(,<�^1<�6<<�:<3z=<[k><��=<s�;<z9<�e6<�;4<w3<f�2<%4<'6<A�8<��;<A�=<��><�=<�G;<!67<U2<V�,<4t(<�%<�;%<� '<1+<�;0<�k5<	{9<œ;<�M;<0�8<�L4<� /<�*<�t&<�%<&<v?)<�-<83<�,8<�;<�
><j><�A=<��:<�<8<�5<-�3<��2<hA3<K�4<�	7<#�9<i`<<$><�p><|=<�:<ӎ5<I0<v6+< J'<�C%<��%<D8(<ڰ,<��1<h�6<�k:<��;<v�:<Sh7<M�2<�A-<�(<��%<�+%<!�&<��*<��/<�4<!�9<��<<a]><�0><�<<o:<uR7<��4<}Y3<��2<�3<`5<��7<��:<�	=<TW><'><x=<<h�8<��3<�y.<��)<�T&<i%<�+&<��)<Gd.<v�3<�E8<�;<�;<��9<��5<��0<��+<�q'<"K%<&�%<�(<�E,<@y1<��6<��:<؋=<�y><��=<��;<q#9<�g6<:4<�3<p�2<�4<�6<��8<�};<j�=<f><�=<';<u7<��1<`�,<�H(<Z�%<V%<��&<��*<L0<�75<4G9<=`;<�;<R�8<�4<��.<�)<bH&<\�$<��%<�)<5�-<�3<8<��;<�=<�:><=<6�:<�8<�n5<��3<[�2<�	3<�{4<G�6<ӗ9<t)<<��=<:><�<<��9<nW5<�0<��*<�'<�%<�S%<��'<o,<��1<��6<j':<�|;<$k:< &7<�T2<�-<�e(<�%<�  �  ��,<�A.<o1<��4<Ӄ8<��;<�=<�><�'><N�<<-;<#9<�7<$�6<YG6<e�6<�7<�9<�~;<7<=<�T><�o><pX=<H
;<��7<{�3<�n0<j�-< �,<?F-<̈́/<Z�2<��6<�:<'*<<E�<<84;<p^8<ܫ4<��0<S.<e�,<�+-<�./<kc2<�'6<	�9<��<<�6><5�><��=<�t<<+�:<��8<)M7<��6<V�6<�37<��8<a:<�P<<!�=<M�><�j><`�<<,>:<�6<��2<X�/<[|-<\�,<M.<��0<�n4<O-8<�$;<p�<<5{<<x�:<W[7<ڊ3<�0<5�-<��,<��-<=0<\�3<�|7<�:<�O=<Q�><e�><H�=<��;<a�9<@:8<�7<܁6<��6<'�7<�'9<�;<��<<�C><n�><
><D<<a9<�i5<U�1<f�.<�-<g-<k�.<��1<ӱ5<�E9<�;<��<<Y<<3�9<�6<�L2<�/<�)-<��,<�w.<�S1<��4<?�8<��;<��=<��><Z><O=<�B;<W9<(�7<J�6<{6<U�6<�8<3�9<��;<�h=<4><<�>< =<k/;<��7<�4<ɑ0<c�-<x�,<�j-<�/<�3<.�6<?:<AS<<ɹ<<�];<��8<^�4<C1<:C.<{�,<�M-<EN/<x�2<CB6<��9<w�<<KH><��><�=<�|<<�:<E�8<�K7<2�6<a|6<�(7<P8<�O:<�;<<_�=<�><.M><��<<�:<��6<@�2<Gz/<&O-<D�,<��-<ޓ0<�;4<�7<C�:<Q|<<�H<<�`:<�*7<�[3<��/<�n-<p�,<-�-<�0<!�3<R7<��:<-#=<^><zc><�c=</�;<u�9<8<;�6<�I6<5}6<�f7<[�8<��:<��<<�><ڂ><��=<��;<7�8<�15<&~1<ʁ.<y�,<��,<�.<��1<�o5<%9<�;<ی<<��;<�\9<��5<�2<��.<��,<�  �  �4<�&5<G�6<��8<��:<tP<<�=<a0=<��<<b<<�$;<|]:<}�9<�9<f�9<�9<��9<��:<@W;<�5<<Y�<< :=<��<<�<<�:<�8<Y�6<��4< 4<�4<n/5<W7<�D9<�B;<�<<*�<<��;<9:<�8<P�5<�}4<��3<kn4<��5<��7<��9<��;<0�<<eM=<�:=<ͮ<<P�;<�;<�O:<��9<�9<T�9<��9<�G:<{�:<;�;<�<<�E=<ck=<��<<5�;<:<�8<96<�4<.!4<��4<��5<t�7<�.:<o�;<$�<<��<<*�;<#�9<�w7<e�5<�S4<�4<>�4<_v6<�x8<�|:<�<<N=<�g=<�&=<�}<<�;<C�:<D1:<K�9<G�9<t�9<n:<6�:<XD;<�"<<��<<%`=<�R=<@�<<K;<:i9<lX7<�5<N_4<s4<�4<ތ6<��8<��:<hf<<=<�<<;<��8<Q�6<	5<:'4<3J4<R\5<�7<�,9<�;<��<<�D=<�b=<��<<8<<Y;<O�:<�
:<�9<,�9<	�9<� :<�:<Ά;</c<<�=<�c=<"=<�9<<��:<ů8<��6<�5<�$4<&<4<�T5<57<�k9<�j;<��<<0�<<�<<�a:<�48<,6<,�4<�4<��4<��5<l�7<��9<*�;<��<<�^=<!I=<��<<T�;<�;<:Q:<k�9<L�9<_�9<��9<f9:<�:<��;<m�<<&+=<�M=<\�<<�;<�9<d�7<�5<�4<��3<M_4<1�5<%�7<��9<��;<~�<<Ԝ<<o;<9<�H7<�X5<'4<�3<g�4<�K6<�M8<~Q:<��;<��<<�8=<3�<<�J<<�n;<_�:<�9<�9<j�9<K�9<M�9<aJ:< ;<:�;<��<<g)=<V=<�l<<;<�19<�7<O5<�#4<s�3<��4<�L6<�t8<��:<R$<<��<<�C<<��:<��8<�6<��4<��3<�  �  L�9<�D:<s�:<�;<@;<��:<�=:<��9<7d9<�`9<g�9<�U:<�
;<��;<��;<;<��:<�/:<��9<
[9<Hs9<��9<�a:<��:<,;<�;<Ը:<>0:<Ʊ9<i9<�u9<6�9<Ӂ:<55;<�;<��;<�y;<{�:<�$:<��9<�j9<�9<��9<��:<�;<TD;<5$;<��:<�.:<�9<�{9<T�9<:<ֹ:<Gj;<��;<��;<�;<t�:<�):<�9<'�9<��9<>8:<��:<7:;<&g;<�7;<B�:<y8:<��9<
�9<��9<8B:<��:<�;<l�;<�;<�t;<t�:<G:<��9<��9<E�9<wH:<f�:<�;;<$X;<�;<h�:<�:<
�9<-�9<��9<�R:<4;<��;<��;<��;<�V;<Т:<��9<��9<�9<��9<]c:<��:<�J;< X;<�;<�:<�:<ܤ9<}�9<��9<�s:<=);<��;<�<<��;<r<;<r�:<��9<Q�9<y�9<2�9<�y:<j�:<�Q;<�N;<��:<Tp:<p�9<ė9<�9<��9<t�:<�@;<��;<��;<G�;<�;<Cb:<Z�9<��9<ϟ9<�:<,�:<@
;<UQ;<�>;<��:<�S:<��9<h�9<��9<(:<��:<�\;<6�;<,�;<{�;<��:<\L:<�9<��9<�9<!:<h�:<+%;<^;<+;;<��:<�?:< �9<��9<?�9<�:<p�:<�h;<�;<�;<�t;<+�:<2:<i�9<�t9<<�9<�:<F�:<-;<�A;<�;<�:<:<��9<Nh9<��9<p:<��:<�g;<E�;<m�;<�C;<��:<��9<y9<Nb9<��9<i:<��:<�;<^,;<��:<*o:<��9<Qy9<�W9<X�9<�:<��:<ap;< �;<��;<�;<Ei:<��9<je9<�^9<��9<�,:<3�:<�;<� ;<��:<�Q:<0�9<�h9<�U9<��9<�3:<��:<߀;<��;<��;<.�:<�H:<L�9<�[9<�d9<�  �  �0=<=<�?<<��:<��8<��6<45<�4<��3<�4<U�6<��8<��:<�U<<��<<�<<�}:<�Z8<�66<��4<�3<664<[m5<'E7<�W9<;5;<x�<<L,=<�1=<��<<��;<�;<�O:<O�9<&�9<B�9<B�9<�:<~�:<9�;<�i<<t=<<M=<�<<��;<�M:<�G8<J6<s�4<�4<1L4<��5<Ӄ7<��9<��;<��<<G�<<�;<��9<��7<��5<�u4<54<��4<w26<=+8<O8:<��;<�=<[t=<yI=<��<<J�;<a�:<�P:<e�9<|�9<��9<��9<oj:<� ;<��;<��<<�Q=<c\=<��<<�;<R�9<��7<@�5<}4<�4<߭4<U56<R8<�}:<�.<<��<<_�<<�U;<fQ9<�7<ZE5<�:4<�24<� 5<'�6<��8<�:<�S<<�2=<uk=<�=<�_<<��;<��:<�!:<>�9<f�9<)�9<�:<��:<di;<�G<<[=<7g=<�?=<�s<<� ;<�9<L 7<�E5<?4<�)4<5<<�6<>9<�;<�<<��<<�N<<ǲ:<F�8<�h6<I�4<�4<�a4<��5<�l7<�}9<Z;<��<<P=<�U=<�<<�<<~3;<Gv:<��9<��9<=�9<2�9<7::<P�:<��;<M�<<4=<�m=<u=<�<<g:<�^8<�]6<g�4<�4<W4<T�5<��7<�9<�;<�<<S�<<��;<��9<A�7<V�5<G^4<��3<l�4<Y6<n8<�:<��;<��<<YH=<�=<�}<<ߤ;< �:<�:<��9<Ր9<Δ9<��9<;:<��:<��;<��<<�%=< 1=<K�<<�_;<��9<}7<;�5<IL4<N�3<Oy4<��5<8<JD:<��;<˾<<fo<<!;<#9<V�6<�5<4<��3<Q�4<�6<��8<^�:<b<<i�<<�1=<��<<n#<<�D;<�u:<J�9<y�9<�|9<�9<Z�9<�c:<�-;<�<<`�<<�  �  �z><��=<:z;<Q8<�4<��0<^#.<3�,<-<��.<F2<>6<ʋ9<��;<!�<<{;<��8<�>5<�x1<Bm.<��,<
�,<��.<$�1<Aq5<�9<l<<��=<N�><><��<<y�:<��8<3d7<�6<�\6<��6<M+8<��9<��;<�=<><j><=<?�:<.47<�k3<" 0<��-<c�,<T�-<Q0<B�3<�{7<أ:<v<<�<<��:<,�7<�&4<χ0<�-<��,<s�-<��/<� 3<��6<�l:< =<�}><��><B�=<|C<<T:<��8<y67<��6<��6<Yo7<��8<6�:<��<<�><S�><>:><��<<��9<�6<dH2<�"/<7-<�,<�^.<#K1<N	5<ܶ8<�|;<��<<:C<<�:<�6<��2<6�/<�]-<Y�,<�.<��0<yY4<�8<�`;</�=<��><t~><�[=<ٙ;<d�9<��7<#�6<��6<��6<W�7<�u9<lb;<e/=<~h><y�><�=<��;<��8<��4<#1<LV.<��,<�6-<J4/<�|2<�N6<��9<!<<5�<<|�;<9<�s5<��1<�.<�,<T-<��.<R�1<Η5<(E9<�:<<�><`�><i/><q�<<�:<�
9<�7<]�6<+�6<E7<TR8<<:<3<<�=<+�><6�><<=<�:<PM7<!�3<�0<��-<6�,<!�-<&0<�3<}7<3�:<Jq<<(�<<��:<��7<�4<ss0<��-<��,<Gk-<��/<��2<��6< E:<v�<<R><E�><t�=<�<<T#:<dU8<7<�`6<Dt6<\?7<ү8<�:<�r<<m�=<��><�><<W<<�|9<	�5<@2<6�.<y-<��,<0).<�1<Z�4<�|8<|A;<5�<<g<<&�9< �6<կ2<N/<�%-<�,<M�-<ӑ0<k#4<��7<�);<Lh=<|n><&D><^ =<];<�l9<v�7<r�6<�A6<n�6<�7<�99<�';<p�<<)1><�  �   ><��<<�/9<�~4<�//<�=*<��&<��$<��%<\�(<�O-<Ϣ2<�d7<)�:<J~;<�:<7r6<tv1<-,<��'<&F%<%<dC'<�G+<�e0<��5<�:<�=<�K><��=<3<<�}9<�6<o4<�3<��2<α3<g�5<�B8<Q;<�==<U><�=<í;<��7<��2<�-<$�(<��%<�%<�&<�/*<�9/<�4<��8<QM;<Eq;<,99<25<��/<��*<��&<'%<M�%<u�(<J-<�c2<�y7<1z;<U�=<i�><��=<W{;<x�8<�6<�
4<�3<�#3<�f4<P�6<LX9<j�;<��=<�{><ur=<H�:<�^6<)1<��+<[�'<�m%<hU%<�'<w�+<G1<R,6<��9<ڮ;<";<�8<Ur3<.<pM)<J&<�%<K�&<�)<|�.<�4<��8<�m<<&>><�V><t�<<��:<N�7<H5<�3<��2<Rn3<55<y}7<lE:<_�<<#@><cU><׶<<�b9<��4<*b/<ep*<�&<� %<��%<��(<�-<
�2<��7<P�:<I�;<E@:<}�6<3�1<�`,<p�'<�u%<'I%<9n'<�p+<�0<]�5<h>:<#5=<�o><� ><;<< �9<��6<��4<�33<��2<��3<��5<�h8<*;<aa=<�v><��=<z�;<��7<|�2<R�-<�)<��%<T%<Ò&<�7*<i>/<��4<��8<�H;<Ri;<.9<5<q�/<r�*<��&<�%<A�%<��(<��,<�>2<�R7<�P;<�=<iZ><k=<�K;< �8<��5<��3<��2<��2<O74<xm6<Y*9<U�;<��=<�O><�F=<�:<W26<��0<B�+< �'<{;%<"!%<�f'<O�+<z�0<5�5<ȹ9<Vr;<��:<��7<�63<��-<�)<��%<��$<�I&<�)<��.<��3<R�8<i6<<�><B><��<<W:<{�7<�
5<YQ3<׫2<13<��4<AB7<�:<�<<]	><�  �  ��<<�:<?\6<�w0<��)<�$<0�<N
<�%<M�"<S�(<�G/<5<n�8<�:<HR8<��3<��-<_'<��!<��<N4<K� <HH%<<o+<��1<j�7<g;<3*=<�<<��:<��7<Ow4<?�1<F�/<&�/<�0<�3<uQ6<_�9<�,<<MN=<F�<<�9<�4<�j.<D�'<��"<d
<�7<�H <y�$<�+<M�1<@�6<�9<�:<�K7<p92<��+<}�%<D� <�b<��<�!"<�m'<0�-<R!4<@>9<�o<<�{=<g�<<�:<��6<��3<�1<��/<�/<�1<JH4<��7<�:<��<<�b=<^�;<�58<\�2<T,<�&<�.!<t�<n�<��!<��&<�X-<3<�/8<_K:<�x9<!�5<�80<�)<��#<c�<�;<�<��#<�u)<��/<I�5<q:<��<<U=<��;<�9<q�5<��2<0<h�/<�U0<\Z2<2Z5<�8<��;<�?=<�=<��:<2�6<��0<5**<�@$<� <�><�Z<�/#< �(<��/<�Q5<A09<GV:<`�8<�'4<^.<��'<
"<�<�a<�� <�q%<��+<�2<�7<��;<{N=<o�<<o ;< �7<�4<��1<�0<�/<��0<%D3<�v6<Ͽ9<�O<<�o=<۟<<��9<C�4<;�.<\(<��"<�< E<WS <�$<9+<��1<��6<=�9<��9<�@7<G+2<p�+<=~%<� <�H<�<�"<�K'<q�-<E�3<9<�D<<�N=<G_<<��9<�6<o3<#�0<M�/<��/<�^1<�4<.i7<�:<��<<7=<��;<�	8<��2<g&,<o�%<�� <�S<�u<�n!<ѯ&<M-<�Q3<�7<>:<v;9<g�5<��/<'{)<�#<�q<<vy<�y#<@@)<�/<#�5<�H:<��<<=<��;<��8<N|5<�h2<
B0<jp/<<0<�2<�5<�w8<�\;<?	=<�  �  p�;<J9<�4< j-<|-&<��<^<�S<?�<^<˘%<�,<X3<`�7<E�8<��6<
2<B+<�	$<�<�&<�w<��<�!<��'<�/<ig5<��9<�<<�;<ȳ9<�e6<��2<2�/<9�-<�W-<��.<�F1<�4<�Z8<b;<�;<<40;<O�7<�2<�+<;�#<<kM<�<J<�<!<�((<�V/<XA5<��8<��8<��5<�0<1)<� "<�<��<�(<%�<a[#<�n*<�1<TZ7<�;<�e<<�|;<��8<_5<��1<"/<��-<��-<��/<Ҋ2<s(6<��9<$�;<�C<<�i:<�+6<��/<��(<��!<��<��<q<��<h#<6�*<M�1<��6<�+9<�=8<514<��-<�&<��<L<׉<��<�C<r�%<"�,<p�3<m�8<��;<
G<<<�:<�7<+4<��0<oZ.<�p-<W,.<;j0<&�3<�Z7<v:<�2<<1�;<�@9<�G4<��-<�_&<r�<�O<Y�<��<EQ<��%<4-<��3<��7<j89<h27<�D2<y+<�>$<�<'W<ʥ<Z<B/!<��'<�-/<��5<D
:<.)<<m�;<|�9<��6<w�2<R�/<��-<!~-<�.<�l1<Z�4< 8<E<;<6]<<�O;<��7<�52< 5+<:$<�<�]<��<�<TD!<\-(<!X/<�?5<ץ8<�8<��5<y0<��(<c�!<�u<��<�<�t<.9#<�I*<+]1<L17<��:<9<<�N;<�8<>/5<D�1<��.<Rd-<��-<CX/<M\2<��5<�]9<դ;<�<<�=:<��5<��/<��(<D�!<�^<��<<�<b[<6F#<Yr*< \1<��6<]�8<i 8<'�3<��-<�d&<��<\<KR<3�<�<�b%<��,<�e3<̘8<��;<d<<v�:<�7<u�3<3�0<�.<04-<<�-<�.0<�|3<�!7<�>:<��;<�  �  8;<�h8<�53<�F,<��$<�<in<ɧ<�)<�<�v$<��+<�2<�57<K�8<u6<qY1<UR*<��"<~~<�<��<$C<�z<Aw&<��-<��4<�K9<j�;<J_;<�;9<��5<H 2<,�.<�,<��,<Y�-<��0<�34<u�7<3�:<n�;<5�:<�7<�%1<&�)<�"<d<�<j�<H�<$�<@'<)�.<��4<78<�j8<�:5<�W/<��'<�� <0<�!<7x<|�<h�!<�-)<8�0<��6<~�:<�;<;<gf8<2�4<&1<�F.<�,<�,<A�.<��1<��5<�9<Ta;<N�;<��9<b5<��.<�w'<�] <��<<$�<Q!<tH"<Q�)<��0<�B6<�8<H�7<�3<�-<�%<֞<)�<��<�I<{�<G/$<��+<��2<�$8<�<;<�;<�H:<�97<r�3<v0<�-<1�,<sf-<ϵ/<�3<A�6<T:<��;<�l;</�8<�h3<Iy,<��$<�M<ޡ<E�<i_<�<�$<3,<��2<p7<��8<Ǯ6<�1<o�*<�#<x�<��<�<�n<��<�&<&.<�4<]p9<ư;<��;<�`9<��5<�E2<?/<t-<�,<�.<��0<�X4<��7<�:<��;<��:<&"7<�@1<��)<�"<]w<��<��<ڎ<��<� '<��.<
�4<K28<�b8<�/5<�I/<��'<�� <�<�<X[<��<=�!<?	)<S`0<�t6<�]:<��;<2�:<p78<q�4<��0<T.<ә,<��,<�.<'�1<m5<��8<5;<c�;<Ĩ9<�55<�.<�I'<s. <��<��<�L<��<"<P{)<1�0<�6<G�8<��7<�S3<N�,<�I%<�d<g�<��<<�u<��#<p+<!2<]�7<g;<��;<8:<8�6<�G3<G�/<xY-<�h,<|*-<�z/<��2<s�6<��9<��;<�  �  p�;<J9<�4< j-<|-&<��<^<�S<?�<^<˘%<�,<X3<`�7<E�8<��6<
2<B+<�	$<�<�&<�w<��<�!<��'<�/<ig5<��9<�<<�;<ȳ9<�e6<��2<2�/<9�-<�W-<��.<�F1<�4<�Z8<b;<�;<<40;<O�7<�2<�+<;�#<<kM<�<J<�<!<�((<�V/<XA5<��8<��8<��5<�0<1)<� "<�<��<�(<%�<a[#<�n*<�1<TZ7<�;<�e<<�|;<��8<_5<��1<"/<��-<��-<��/<Ҋ2<s(6<��9<$�;<�C<<�i:<�+6<��/<��(<��!<��<��<q<��<h#<6�*<M�1<��6<�+9<�=8<514<��-<�&<��<L<׉<��<�C<r�%<"�,<p�3<m�8<��;<
G<<<�:<�7<+4<��0<oZ.<�p-<W,.<;j0<&�3<�Z7<v:<�2<<1�;<�@9<�G4<��-<�_&<r�<�O<Y�<��<EQ<��%<4-<��3<��7<j89<h27<�D2<y+<�>$<�<'W<ʥ<Z<B/!<��'<�-/<��5<D
:<.)<<m�;<|�9<��6<w�2<R�/<��-<!~-<�.<�l1<Z�4< 8<E<;<6]<<�O;<��7<�52< 5+<:$<�<�]<��<�<TD!<\-(<!X/<�?5<ץ8<�8<��5<y0<��(<c�!<�u<��<�<�t<.9#<�I*<+]1<L17<��:<9<<�N;<�8<>/5<D�1<��.<Rd-<��-<CX/<M\2<��5<�]9<դ;<�<<�=:<��5<��/<��(<D�!<�^<��<<�<b[<6F#<Yr*< \1<��6<]�8<i 8<'�3<��-<�d&<��<\<KR<3�<�<�b%<��,<�e3<̘8<��;<d<<v�:<�7<u�3<3�0<�.<04-<<�-<�.0<�|3<�!7<�>:<��;<�  �  ��<<�:<?\6<�w0<��)<�$<0�<N
<�%<M�"<S�(<�G/<5<n�8<�:<HR8<��3<��-<_'<��!<��<N4<K� <HH%<<o+<��1<j�7<g;<3*=<�<<��:<��7<Ow4<?�1<F�/<&�/<�0<�3<uQ6<_�9<�,<<MN=<F�<<�9<�4<�j.<D�'<��"<d
<�7<�H <y�$<�+<M�1<@�6<�9<�:<�K7<p92<��+<}�%<D� <�b<��<�!"<�m'<0�-<R!4<@>9<�o<<�{=<g�<<�:<��6<��3<�1<��/<�/<�1<JH4<��7<�:<��<<�b=<^�;<�58<\�2<T,<�&<�.!<t�<n�<��!<��&<�X-<3<�/8<_K:<�x9<!�5<�80<�)<��#<c�<�;<�<��#<�u)<��/<I�5<q:<��<<U=<��;<�9<q�5<��2<0<h�/<�U0<\Z2<2Z5<�8<��;<�?=<�=<��:<2�6<��0<5**<�@$<� <�><�Z<�/#< �(<��/<�Q5<A09<GV:<`�8<�'4<^.<��'<
"<�<�a<�� <�q%<��+<�2<�7<��;<{N=<o�<<o ;< �7<�4<��1<�0<�/<��0<%D3<�v6<Ͽ9<�O<<�o=<۟<<��9<C�4<;�.<\(<��"<�< E<WS <�$<9+<��1<��6<=�9<��9<�@7<G+2<p�+<=~%<� <�H<�<�"<�K'<q�-<E�3<9<�D<<�N=<G_<<��9<�6<o3<#�0<M�/<��/<�^1<�4<.i7<�:<��<<7=<��;<�	8<��2<g&,<o�%<�� <�S<�u<�n!<ѯ&<M-<�Q3<�7<>:<v;9<g�5<��/<'{)<�#<�q<<vy<�y#<@@)<�/<#�5<�H:<��<<=<��;<��8<N|5<�h2<
B0<jp/<<0<�2<�5<�w8<�\;<?	=<�  �   ><��<<�/9<�~4<�//<�=*<��&<��$<��%<\�(<�O-<Ϣ2<�d7<)�:<J~;<�:<7r6<tv1<-,<��'<&F%<%<dC'<�G+<�e0<��5<�:<�=<�K><��=<3<<�}9<�6<o4<�3<��2<α3<g�5<�B8<Q;<�==<U><�=<í;<��7<��2<�-<$�(<��%<�%<�&<�/*<�9/<�4<��8<QM;<Eq;<,99<25<��/<��*<��&<'%<M�%<u�(<J-<�c2<�y7<1z;<U�=<i�><��=<W{;<x�8<�6<�
4<�3<�#3<�f4<P�6<LX9<j�;<��=<�{><ur=<H�:<�^6<)1<��+<[�'<�m%<hU%<�'<w�+<G1<R,6<��9<ڮ;<";<�8<Ur3<.<pM)<J&<�%<K�&<�)<|�.<�4<��8<�m<<&>><�V><t�<<��:<N�7<H5<�3<��2<Rn3<55<y}7<lE:<_�<<#@><cU><׶<<�b9<��4<*b/<ep*<�&<� %<��%<��(<�-<
�2<��7<P�:<I�;<E@:<}�6<3�1<�`,<p�'<�u%<'I%<9n'<�p+<�0<]�5<h>:<#5=<�o><� ><;<< �9<��6<��4<�33<��2<��3<��5<�h8<*;<aa=<�v><��=<z�;<��7<|�2<R�-<�)<��%<T%<Ò&<�7*<i>/<��4<��8<�H;<Ri;<.9<5<q�/<r�*<��&<�%<A�%<��(<��,<�>2<�R7<�P;<�=<iZ><k=<�K;< �8<��5<��3<��2<��2<O74<xm6<Y*9<U�;<��=<�O><�F=<�:<W26<��0<B�+< �'<{;%<"!%<�f'<O�+<z�0<5�5<ȹ9<Vr;<��:<��7<�63<��-<�)<��%<��$<�I&<�)<��.<��3<R�8<i6<<�><B><��<<W:<{�7<�
5<YQ3<׫2<13<��4<AB7<�:<�<<]	><�  �  �z><��=<:z;<Q8<�4<��0<^#.<3�,<-<��.<F2<>6<ʋ9<��;<!�<<{;<��8<�>5<�x1<Bm.<��,<
�,<��.<$�1<Aq5<�9<l<<��=<N�><><��<<y�:<��8<3d7<�6<�\6<��6<M+8<��9<��;<�=<><j><=<?�:<.47<�k3<" 0<��-<c�,<T�-<Q0<B�3<�{7<أ:<v<<�<<��:<,�7<�&4<χ0<�-<��,<s�-<��/<� 3<��6<�l:< =<�}><��><B�=<|C<<T:<��8<y67<��6<��6<Yo7<��8<6�:<��<<�><S�><>:><��<<��9<�6<dH2<�"/<7-<�,<�^.<#K1<N	5<ܶ8<�|;<��<<:C<<�:<�6<��2<6�/<�]-<Y�,<�.<��0<yY4<�8<�`;</�=<��><t~><�[=<ٙ;<d�9<��7<#�6<��6<��6<W�7<�u9<lb;<e/=<~h><y�><�=<��;<��8<��4<#1<LV.<��,<�6-<J4/<�|2<�N6<��9<!<<5�<<|�;<9<�s5<��1<�.<�,<T-<��.<R�1<Η5<(E9<�:<<�><`�><i/><q�<<�:<�
9<�7<]�6<+�6<E7<TR8<<:<3<<�=<+�><6�><<=<�:<PM7<!�3<�0<��-<6�,<!�-<&0<�3<}7<3�:<Jq<<(�<<��:<��7<�4<ss0<��-<��,<Gk-<��/<��2<��6< E:<v�<<R><E�><t�=<�<<T#:<dU8<7<�`6<Dt6<\?7<ү8<�:<�r<<m�=<��><�><<W<<�|9<	�5<@2<6�.<y-<��,<0).<�1<Z�4<�|8<|A;<5�<<g<<&�9< �6<կ2<N/<�%-<�,<M�-<ӑ0<k#4<��7<�);<Lh=<|n><&D><^ =<];<�l9<v�7<r�6<�A6<n�6<�7<�99<�';<p�<<)1><�  �  �0=<=<�?<<��:<��8<��6<45<�4<��3<�4<U�6<��8<��:<�U<<��<<�<<�}:<�Z8<�66<��4<�3<664<[m5<'E7<�W9<;5;<x�<<L,=<�1=<��<<��;<�;<�O:<O�9<&�9<B�9<B�9<�:<~�:<9�;<�i<<t=<<M=<�<<��;<�M:<�G8<J6<s�4<�4<1L4<��5<Ӄ7<��9<��;<��<<G�<<�;<��9<��7<��5<�u4<54<��4<w26<=+8<O8:<��;<�=<[t=<yI=<��<<J�;<a�:<�P:<e�9<|�9<��9<��9<oj:<� ;<��;<��<<�Q=<c\=<��<<�;<R�9<��7<@�5<}4<�4<߭4<U56<R8<�}:<�.<<��<<_�<<�U;<fQ9<�7<ZE5<�:4<�24<� 5<'�6<��8<�:<�S<<�2=<uk=<�=<�_<<��;<��:<�!:<>�9<f�9<)�9<�:<��:<di;<�G<<[=<7g=<�?=<�s<<� ;<�9<L 7<�E5<?4<�)4<5<<�6<>9<�;<�<<��<<�N<<ǲ:<F�8<�h6<I�4<�4<�a4<��5<�l7<�}9<Z;<��<<P=<�U=<�<<�<<~3;<Gv:<��9<��9<=�9<2�9<7::<P�:<��;<M�<<4=<�m=<u=<�<<g:<�^8<�]6<g�4<�4<W4<T�5<��7<�9<�;<�<<S�<<��;<��9<A�7<V�5<G^4<��3<l�4<Y6<n8<�:<��;<��<<YH=<�=<�}<<ߤ;< �:<�:<��9<Ր9<Δ9<��9<;:<��:<��;<��<<�%=< 1=<K�<<�_;<��9<}7<;�5<IL4<N�3<Oy4<��5<8<JD:<��;<˾<<fo<<!;<#9<V�6<�5<4<��3<Q�4<�6<��8<^�:<b<<i�<<�1=<��<<n#<<�D;<�u:<J�9<y�9<�|9<�9<Z�9<�c:<�-;<�<<`�<<�  �  L�9<�D:<s�:<�;<@;<��:<�=:<��9<7d9<�`9<g�9<�U:<�
;<��;<��;<;<��:<�/:<��9<
[9<Hs9<��9<�a:<��:<,;<�;<Ը:<>0:<Ʊ9<i9<�u9<6�9<Ӂ:<55;<�;<��;<�y;<{�:<�$:<��9<�j9<�9<��9<��:<�;<TD;<5$;<��:<�.:<�9<�{9<T�9<:<ֹ:<Gj;<��;<��;<�;<t�:<�):<�9<'�9<��9<>8:<��:<7:;<&g;<�7;<B�:<y8:<��9<
�9<��9<8B:<��:<�;<l�;<�;<�t;<t�:<G:<��9<��9<E�9<wH:<f�:<�;;<$X;<�;<h�:<�:<
�9<-�9<��9<�R:<4;<��;<��;<��;<�V;<Т:<��9<��9<�9<��9<]c:<��:<�J;< X;<�;<�:<�:<ܤ9<}�9<��9<�s:<=);<��;<�<<��;<r<;<r�:<��9<Q�9<y�9<2�9<�y:<j�:<�Q;<�N;<��:<Tp:<p�9<ė9<�9<��9<t�:<�@;<��;<��;<G�;<�;<Cb:<Z�9<��9<ϟ9<�:<,�:<@
;<UQ;<�>;<��:<�S:<��9<h�9<��9<(:<��:<�\;<6�;<,�;<{�;<��:<\L:<�9<��9<�9<!:<h�:<+%;<^;<+;;<��:<�?:< �9<��9<?�9<�:<p�:<�h;<�;<�;<�t;<+�:<2:<i�9<�t9<<�9<�:<F�:<-;<�A;<�;<�:<:<��9<Nh9<��9<p:<��:<�g;<E�;<m�;<�C;<��:<��9<y9<Nb9<��9<i:<��:<�;<^,;<��:<*o:<��9<Qy9<�W9<X�9<�:<��:<ap;< �;<��;<�;<Ei:<��9<je9<�^9<��9<�,:<3�:<�;<� ;<��:<�Q:<0�9<�h9<�U9<��9<�3:<��:<߀;<��;<��;<.�:<�H:<L�9<�[9<�d9<�  �  �4<�&5<G�6<��8<��:<tP<<�=<a0=<��<<b<<�$;<|]:<}�9<�9<f�9<�9<��9<��:<@W;<�5<<Y�<< :=<��<<�<<�:<�8<Y�6<��4< 4<�4<n/5<W7<�D9<�B;<�<<*�<<��;<9:<�8<P�5<�}4<��3<kn4<��5<��7<��9<��;<0�<<eM=<�:=<ͮ<<P�;<�;<�O:<��9<�9<T�9<��9<�G:<{�:<;�;<�<<�E=<ck=<��<<5�;<:<�8<96<�4<.!4<��4<��5<t�7<�.:<o�;<$�<<��<<*�;<#�9<�w7<e�5<�S4<�4<>�4<_v6<�x8<�|:<�<<N=<�g=<�&=<�}<<�;<C�:<D1:<K�9<G�9<t�9<n:<6�:<XD;<�"<<��<<%`=<�R=<@�<<K;<:i9<lX7<�5<N_4<s4<�4<ތ6<��8<��:<hf<<=<�<<;<��8<Q�6<	5<:'4<3J4<R\5<�7<�,9<�;<��<<�D=<�b=<��<<8<<Y;<O�:<�
:<�9<,�9<	�9<� :<�:<Ά;</c<<�=<�c=<"=<�9<<��:<ů8<��6<�5<�$4<&<4<�T5<57<�k9<�j;<��<<0�<<�<<�a:<�48<,6<,�4<�4<��4<��5<l�7<��9<*�;<��<<�^=<!I=<��<<T�;<�;<:Q:<k�9<L�9<_�9<��9<f9:<�:<��;<m�<<&+=<�M=<\�<<�;<�9<d�7<�5<�4<��3<M_4<1�5<%�7<��9<��;<~�<<Ԝ<<o;<9<�H7<�X5<'4<�3<g�4<�K6<�M8<~Q:<��;<��<<�8=<3�<<�J<<�n;<_�:<�9<�9<j�9<K�9<M�9<aJ:< ;<:�;<��<<g)=<V=<�l<<;<�19<�7<O5<�#4<s�3<��4<�L6<�t8<��:<R$<<��<<�C<<��:<��8<�6<��4<��3<�  �  ��,<�A.<o1<��4<Ӄ8<��;<�=<�><�'><N�<<-;<#9<�7<$�6<YG6<e�6<�7<�9<�~;<7<=<�T><�o><pX=<H
;<��7<{�3<�n0<j�-< �,<?F-<̈́/<Z�2<��6<�:<'*<<E�<<84;<p^8<ܫ4<��0<S.<e�,<�+-<�./<kc2<�'6<	�9<��<<�6><5�><��=<�t<<+�:<��8<)M7<��6<V�6<�37<��8<a:<�P<<!�=<M�><�j><`�<<,>:<�6<��2<X�/<[|-<\�,<M.<��0<�n4<O-8<�$;<p�<<5{<<x�:<W[7<ڊ3<�0<5�-<��,<��-<=0<\�3<�|7<�:<�O=<Q�><e�><H�=<��;<a�9<@:8<�7<܁6<��6<'�7<�'9<�;<��<<�C><n�><
><D<<a9<�i5<U�1<f�.<�-<g-<k�.<��1<ӱ5<�E9<�;<��<<Y<<3�9<�6<�L2<�/<�)-<��,<�w.<�S1<��4<?�8<��;<��=<��><Z><O=<�B;<W9<(�7<J�6<{6<U�6<�8<3�9<��;<�h=<4><<�>< =<k/;<��7<�4<ɑ0<c�-<x�,<�j-<�/<�3<.�6<?:<AS<<ɹ<<�];<��8<^�4<C1<:C.<{�,<�M-<EN/<x�2<CB6<��9<w�<<KH><��><�=<�|<<�:<E�8<�K7<2�6<a|6<�(7<P8<�O:<�;<<_�=<�><.M><��<<�:<��6<@�2<Gz/<&O-<D�,<��-<ޓ0<�;4<�7<C�:<Q|<<�H<<�`:<�*7<�[3<��/<�n-<p�,<-�-<�0<!�3<R7<��:<-#=<^><zc><�c=</�;<u�9<8<;�6<�I6<5}6<�f7<[�8<��:<��<<�><ڂ><��=<��;<7�8<�15<&~1<ʁ.<y�,<��,<�.<��1<�o5<%9<�;<ی<<��;<�\9<��5<�2<��.<��,<�  �  O�$<��&<�|*<({/<��4<Jj9<�<<�+><��=<�h<<��9<27<2�4<0&3<��2<�g3<E/5<T�7<f�:<��<<�-><S�=<<<�8</�3<W.<8�)<2&<�$<H&<2])<�=.<Ǝ3<�8< �:<,z;<��9<+�5<��0<�k+<fK'<�&%<�c%<��'<v(,<�^1<�6<<�:<3z=<[k><��=<s�;<z9<�e6<�;4<w3<f�2<%4<'6<A�8<��;<A�=<��><�=<�G;<!67<U2<V�,<4t(<�%<�;%<� '<1+<�;0<�k5<	{9<œ;<�M;<0�8<�L4<� /<�*<�t&<�%<&<v?)<�-<83<�,8<�;<�
><j><�A=<��:<�<8<�5<-�3<��2<hA3<K�4<�	7<#�9<i`<<$><�p><|=<�:<ӎ5<I0<v6+< J'<�C%<��%<D8(<ڰ,<��1<h�6<�k:<��;<v�:<Sh7<M�2<�A-<�(<��%<�+%<!�&<��*<��/<�4<!�9<��<<a]><�0><�<<o:<uR7<��4<}Y3<��2<�3<`5<��7<��:<�	=<TW><'><x=<<h�8<��3<�y.<��)<�T&<i%<�+&<��)<Gd.<v�3<�E8<�;<�;<��9<��5<��0<��+<�q'<"K%<&�%<�(<�E,<@y1<��6<��:<؋=<�y><��=<��;<q#9<�g6<:4<�3<p�2<�4<�6<��8<�};<j�=<f><�=<';<u7<��1<`�,<�H(<Z�%<V%<��&<��*<L0<�75<4G9<=`;<�;<R�8<�4<��.<�)<bH&<\�$<��%<�)<5�-<�3<8<��;<�=<�:><=<6�:<�8<�n5<��3<[�2<�	3<�{4<G�6<ӗ9<t)<<��=<:><�<<��9<nW5<�0<��*<�'<�%<�S%<��'<o,<��1<��6<j':<�|;<$k:< &7<�T2<�-<�e(<�%<�  �  �<8�<{X$<JS*<��0<�6<��:<��<<��<<�<;<qL8<N�4<��1<Y
0<�v/</]0<��2<c�5<9<��;<�+=<��<<E:<4}5<k/<V�(<S=#<�]<�<$�<�#<p�)<e0<+�5<�j9<L:<��7<d3<z�,<$m&<�F!<at<�|<L!<�O&<:�,<�3<\c8<��;<dV=<�<<s~:<^U7<
4<�\1<G�/<��/<&1</�3<17<�;:<�<<�r=<+K<</�8<��3<4w-<L'<�!<)�<�}<g!<.�%<�I,<~�2<)�7<):<�9<��6<0C1<��*<�$<�* <A<]<<%�"<ue(<��.<�5<��9<�<<�d=<�,<<��9<�B6<=3<��0<O�/<�0<��1<�4<�$8<�*;<+=<DJ=<.i;<l7<��1< B+<�*%<ݔ <#]<��<0h"<�'<�s.<]{4<��8<h`:<�9</5<D*/<��(<��"<@;<�G<�1 <r�$<̆*<O1<��6<;<q,=<U0=<�n;<�~8<'5<�02<�<0<٨/<�0<�2<�5<�19<��;<�T=<��<<�B:<8�5<	�/<�)<�_#<-�<4<[�<h$<*<��0<!6<��9<�>:<�7<v=3<��,<V�&<�m!</�<"�<Dl!<wm&<�,<�3<4x8<{ <<e=<��<<��:<aZ7<�4<t[1<��/<��/<�1<Ŭ3<��6<�&:<��<<�W=<(-<<:�8<�3<�P-<"�&<t�!<]�<�M<� <��%<V,<ll2< d7<+�9<�9<pt6<X1<_�*<x$<�<�<	<g�"<�;(<��.<4�4<L�9<�<<�5=<��;<�\9<N6<t�2<ċ0<�|/<��/<x�1<�4<��7<�:<��<<�=<�2;<*57<�1<�	+<��$<EY <�<��<J'"<��'<�/.<�64<�y8<�:<��8<Q�4<��.<�f(<��"<= <�  �  nV<K<1  <Ò&<��-<!j4<�D9<��;<��;<:<n�6<;M3<N
0<&�-<�:-<�;.<P�0<�4<�7<Y�:<�<<Ot;<<e8< 3<1=,<�	%<9�<��<�a<uP<E <��&<,.<TO4<48<B�8<f6<<1<�*<f�"<B+<I�<��<�<�$"<�)<+D0<c6<e�:<�9<<��;<
N9<��5<]H2<6S/<��-<��-<�/<��1<�5<49<��;<�Z<<E�:<'7<�$1<#	*<�#<Y<�<��<�<�m"<W~)<��0<\6<�9<��8<5<�	/<Z�'<�� <��<�<Q�<f\< m$<�+<�2<�8<�f;<:S<<�;<6J8<��4<a<1<�.<�w-<�-<�/<�3<u�6<T:<:
<<�!<<��9<�C5<3�.<̕'<�� <�<�<$�<�n<��$<��+<l�2<vk7<�B9< �7<�F3<��,<Vp%<< �<w�<��<E5 <S�&<+.<՛4<-v9<-�;<$<<DN:<�$7<�3<�<0<c.<ll-<dl.<��0<J4<��7<��:<�E<<�;<R�8<�93<�_,<,%<N�<��<��<�t<�D <g '<0?.<tx4<^8<�9<��6<�>1<}F*<�!#<$R<J<��<k�<dB"<�1)<"\0<	x6<;�:<vH<<�;<QV9<��5<)J2<�Q/<��-<ƅ-<�
/<X�1<Et5<f�8<�t;<�?<<2�:<�6<� 1<w�)<Z�"<b-<��<�<}�<�:"<�J)<LZ0<��5<��8<Yp8<��4<��.<٤'<�� <d�<�l<V<�2<�C$<yl+<�_2<K�7<�9;<�$<<��:<�8<��4<�1<zo.<�A-<R�-<*�/<��2<��6<��9<��;<>�;<�9<5<��.<]'<�� <8�<ed<�A<t-<�f$<��+<z\2<'&7<��8<��7<�3<�q,<�0%<��<؎<�  �  kg><�?<�uB<;XF<�fJ<+�M<^�O<��O<D3N<�?K<R�G<Y�C<|@<:k><��=<>�><�A<�D<mbH<GL<H�N<X�O<�[O<zM<��I<�vE<�A<1:?<Zq><%�?<�{B<��F<�:K<QHO<z�Q<_R<}�P<**M<T�H<>D<��@<U�><�><�@<V�C<��G<ҾK<ئN< �O<��O<zM<�1J<\F<�B<��?<I5><� ><[�?<1VB<�E<��I<�:M<t{O< P<Y�N<X?L<�lH<0ZD<N�@<!�><��><�@<��C<f]H<"�L<ȉP<�xR<>7R<��O<��K<�OG<-C<��?<K�><�3?<8�A<�+E<�EI<��L<�YO<CP<�O<m�L<�H<� E<ܥA<�'?<><q{><�e@<u�C<UJG<�K<3#N<��O<x�O<�7N<�K<DG<C<N@<[�><+?<,�A<WE<��I<D;N<�eQ<�R<��Q<&�N<�eJ<��E<J�A<�U?<��><S�?<��B<ŋF<c�J<�M<��O<4�O<�dN<0qK<ԵG<��C<��@<m�><a><�><�LA<e�D<^�H<�+L<��N<sP<{�O<�?M<�I<��E<��A<$]?<��><9�?<��B<��F<^aK<�oO<ZR<6�R<��P<�QM<$�H<�cD<��@<��><t�><%�@<	�C<��G<1�K<f�N<�P<l�O<ÄM<�9J<�`F<��B<q�?<�0><)><��?<ZHB<)�E<�I<�#M<�aO<xP<��N<RL<;HH</3D<�@<��><~�><Rd@<��C<�,H<��L<'XP<GR<,R<a�O<W�K<<!G<��B<��?<v><,	?<bA<�E<�I<��L<�-O<F�O<v�N<�ZL<�H<��D<^rA<<�><��=<�E><�/@<tKC<[G<
�J<S�M<��O<L�O<?N<U�J<�F<��B<��?<%p><g�><GA<�E<��I<J�M<�#Q<�_R<bQ<�gN<�&J<5�E<n�A<�?<�  �  �b?<�@<�eC<�.G<�K<0JN<�P<?)P<�N<��K<�H<�KD<#(A<�"?<�><4x?<I�A<�E<��H<�kL<BO<�NP<��O<�M<�KJ<7SF<�B< 8@<xj?< z@<<?C<�9G<��K<�{O<��Q<�kR<d�P<SxM<�2I<��D<3�A<ڲ?<��?<'zA<��D<H�H<�gL<N.O<�kP<@�O<��M<m�J<��F<�LC<�}@<��><��><�D@<8�B<+�F<�NJ<ğM<��O<��P<{�O<9�L<�4I<�?E<�A<��?<�?<oA<�D<E�H<�5M<��P<?�R<HR<*P< DL<��G<%�C<��@<�?<�1@<��B<jF<JJ<'�M<��O<'�P<�uO<��L<Y{I<H�E<FLB<��?<s�><�3?<�A<D<�G<.�K<��N<EP<�`P<5�N<i�K<�G<y D<vA<��?<$@<�VB<��E<�XJ<Y~N<ӀQ<խR<��Q<��N<�J<0sF<��B<)A@<�?<I�@<��C<bG<*NK<|N<EP<�ZP<X�N<��K<09H<?}D<�YA<,T?<�><+�?<+�A<$GE<�I<�L<;O<�uP<��O<}�M<�oJ<GvF<��B<[@<�?<4�@<"dC<^_G<+�K<�O<gR<��R<\�P<ܟM<YYI<GE<[�A<>�?<��?<B�A<S�D<X�H<�}L<�AO<w|P<��O<_�M<�J<G�F<xNC<n|@<��><��>< :@<b�B<MuF<�:J<�M<��O<oP<&bO<9�L<I<�E<��A<��?<�?<b@A<7}D<{�H<2M<�}P<�TR<R<��O<�L<I�G<�C<��@<�m?<@@<�WB<I�E<��I<"_M<٫O<UP<QGO<+�L<2JI<ԀE<�B<+�?<0�><�><��@<��C<�G<9LK<�NN<&P<�*P<��N<#�K<�G< �C<��@<dl?<��?<�B<^�E<�J<<N<�>Q<�kR<>zQ<9�N<�J<�5F<�qB<?@<�  �  �(B<�bC<�F<��I<n	M<C�O<tEQ<N*Q<��O<��L<glI<�E<�C<�/A<ɣ@<�~A<2�C<�F<�5J<��M<ZP<�VQ<�Q<QO<�PL<��H<�`E<BC<p)B<��B<\E<�H<.�L<��O<�R<�}R<$Q<=N<F�J<R�F<
�C<�\B<�{B<�:D<Z;G<��J<�1N<�P<ÈQ<��P<�N<Q�K<WcH<�E<�sB<RA<��@<P?B<�D<�
H<��K<ӪN<U�P<y�Q<V�P<Y�N<�[K<��G<��D<)�B<�tB<��C<�F<JJ<E	N<|Q<��R<�eR<�tP<E7M<�gI<@�E<�WC<�SB<��B<
5E<{H<�L<�1O<�"Q<�Q<pP<GN<,�J<�GG<D D<��A<��@<�CA<0�B<��E<!=I<�L<��O<�CQ<s�Q<~AP<�M<B J<řF<��C<qB<R�B<�D<��G<ÍK<�$O<�Q<��R<"�Q<�}O<E�K<*H<��D<��B<�`B<�C<<;F<�I<�;M<+P<wQ<�[Q<�O<�M<<�I<(F<�?C<LaA<��@<�A<o�C<�F<gbJ<w�M<u6P<(~Q<�>Q<�uO<�tL<��H<��E<S(C<�LB<�!C<�E<��H<��L<	 P<9=R<��R<�BQ<_dN<ٯJ<��F<D<:B<�B<�XD<�VG<��J<�GN<��P<X�Q<��P<��N<��K<�gH<YE<>rB<��@<�@<�4B<�D<��G<�yK<	�N<��P<��Q<�P<k�N<7K<�G<nD<�B<	HB<�C<IpF<bJ<�M<�P<PiR<�4R<`DP<�M<�9I<
�E<�+C<L(B<��B<�
E<�PH<[�K<vO<l�P<�aQ<oAP<6�M<��J<�G<Z�C<�A<f�@<�A<��B<��E<�I<�vL<�OO<�Q<EUQ<�
P<�cM<1�I<�`F<*�C<&5B< xB<:[D<�G<�LK<]�N<.zQ<
{R<�Q<�=O<u�K<��G<�D< �B<�  �  �3F<�qG<��I<M�L<��O<��Q<4�R<^R<)�P<}LN<�QK<CUH<��E<%>D<��C<��D<tTF<��H<5L<I�N< >Q<G�R<-�R<�oQ<yO<�!L<�>I<$G<�(F<��F<-SH<��J<�M<�tP<R<aR<�SQ<gO<�EL<SoI<JBG<>9F<��F<�9H<y�J<��M<|�P<y_R<s�R<eR<�,P<~yM<pqJ<t�G<�XE<mD<�D<�,E<�PG<O&J<[3M<:�O<PR<r�R<f�R<J�P<!ZN<�TK< �H<�F<�ZF<Q@G<1SI<ML<�O<�OQ<<�R<�YR<��P<�^N<pK<e�H<A�F<�KF<G<�I<W�K<�N<xbQ<��R<��R<*�Q<�eO<%�L<I<�F<��D<mD<nWD<T�E<�;H<20K<-1N<S�P<^tR<��R<,R<�(P<.UM<�UJ<��G<�F<�zF< �G<X/J<CM<u�O<^�Q<l�R<��Q<�P<�iM<}J<	H<h�F<�kF<��G<vJ<��L<)�O<��Q<��R<��R<��P<z~N<�K<��H</	F<JpD<[�C<}�D<A�F<(I<*.L<�O<�gQ<=�R<��R<�Q<�<O<IEL<�aI<Y=G<ELF<��F<�wH<5K<nN<��P<�9R<��R<{Q<}FO<�kL<��I<fG<<[F<��F<ZWH<��J<��M<��P<�rR<��R<�$R<V7P<�M<�uJ<�G<+WE<�D<+D<�!E<�BG<}J<�M<~�O<��Q<�R<9zR<y�P<�5N<�-K<wH<,�F</.F<G<�#I<��K<��N<�Q<,QR<;)R<��P<�/N<�AK<A�H<�F<1 F<J�F<=�H<��K<6�N<�6Q<�R<�R<pQ<'5O<2VL<�KI<��F<R�D<h�C<� D<��E<�H<��J<��M<)�P<E>R<��R<��Q<��O<QM<�J<��G<hDF<�=F<�G<��I<��L<��O<-�Q<`ZR<
�Q<C�O<�+M<E@J<��G<UF<�  �  ;�J<p�K<��M<�:P<�AR<�S<��S<�5S<ٳQ<O�O<�6M<��J<WI<��G<�uG<QH<<`I<CeK<��M<cP<#R<�sS<�S<X^S<�Q<��O<~M<էK<b�J<ɎJ<�qK<+M<3�N<��P<;�Q<=�Q<Q<��O<5�M<�L<Z�J<�J<= K<��L<q�N<Q<w�R<o�S<*�S<��R<�/Q<��N<�L<[J<��H<Y�G<�G<��H<�*J<XL<g�N<]Q<��R<��S<]T<�+S<mQ<�0O<�M<�hK<��J<�J<�L<d�M<�O<)+Q<��Q<��Q<!�P<�BO<sdM<��K<��J<��J<d�K<kM<��O<��Q<�hS<>T<��S<�yR<��P<�7N<2�K<g�I<MSH<��G<*�G<�I<f�J<�(M<8�O<��Q<QIS<�T<��S<��R< �P<�gN<�^L<	K<��J<�:K<Y�L<qN<9P<%�Q<	R<��Q<'eP<ťN<��L<rXK<�J<}�J<(,L<&N<)nP<qtR<��S<�T<hgS<��Q<��O<�iM<�K<U4I<�H<Y�G<�2H<ŐI<y�K<��M<bHP<fFR<�S< T< �S<�R<l�O<�M<8�K<�J<�J<N�K<�+M<\	O<D�P<c�Q<��Q<�DQ<��O<$N<�?L<�K<��J<�?K<|�L<��N<�)Q<m�R<��S<��S<.�R<%:Q<z�N<f�L<�\J<��H<��G<g�G<ǁH<�J<IGL<��N<��P<�R<d�S<P�S<A
S<�HQ<
O<��L<@>K<�J<(�J<��K<Z�M<M}O<S�P<��Q<G�Q<d�P<�O<r6M<ԓK<W�J<��J<}{K<[@M<�|O<��Q<�<S<<�S<T�S<�IR<�YP<�N<H�K<W�I<TH<WyG<'�G<��H<P�J<��L<�VO<=}Q<S<y�S<y�S<pR<gxP<&/N<�$L<�J<pgJ<\�J<�_L<1N<��O<�AQ<��Q<�ZQ<A&P<hN<��L<�K< nJ<�  �  �N<�P<�Q<��R<T<dcT<�T<HS<��Q<a3P<��N<E#M<��K<KK<~K<�hK<N7L<rqM<��N<��P<�R<�bS<�2T<�dT<��S<g�R<�7Q<��O<~�N<�N<]	N<�~N<�6O<��O<�`P<�wP<�*P<�O<��N<C7N<�N<�XN<�?O<b�P<t#R<��S<TVT<wT<��S<��R<.fQ<�O< :N<v�L<��K<~TK<�NK<��K<u�L<�N<�O<�JQ<��R<�S<��T<V�T<H�S<8qR<��P<��O<��N<0N<�WN<��N<K�O<�IP<��P<$�P<�'P<�wO<f�N<�:N<	/N<��N<��O<�3Q<��R<��S<�T<�kT<'�S<�sR<z�P<RO<��M<4�L<��K<vPK<�uK<L<5M<$�N<W;P<[�Q<�2S<�-T<�T<JNT<7VS<��Q<{cP<b!O<H[N<�'N<8yN<�"O<�O<�nP<<�P<�yP<��O<t7O<�N<�)N<�LN<�O<79P<�Q<�/S<�8T<��T<�>T<QS<�Q<MfP<��N<�VM<�2L<�~K<�JK<�K<�hL<��M<M!O<O�P<�GR<݋S<HZT<�T<�T<��R<�[Q<��O<<�N<�1N<
.N<�N<�\O<7P<m�P<�P<oQP<δO<p�N<�[N<�%N< zN<Z_O<��P<T>R<�S<lT<"�T<��S<�R<�pQ<��O<p>N<��L<��K<�OK<�FK<�K<��L<
N<m�O<a4Q<F�R<��S<�jT<�^T<S�S<�JR<�P<�^O<�hN<kN<�(N<�N<wO<�P<@qP<eP<f�O<�HO<��N<�N<�N<5�N<��O<	Q<{�R<A�S<r\T<>T<A~S<�CR<��P<�O<)�M<dTL<�xK<#K<>K<Y�K<s�L<�jN<aP<��Q<V�R<��S<�`T<�T<�S<��Q<K*P<�N<�N<�M<O;N<�N<��O<8/P<�gP<�:P<��O<�N<WLN<��M<�N<�  �  ��Q<|�R<|�S<VT<RT<ƽS<��R<x�Q<�P<H�O<�O<ݖN< UN<5N<�,N<B:N<FaN<<�N<�(O<�O<��P<�Q<1	S<k�S<�gT<�JT<��S<+�R<��Q<C{P<��O<3�N<��N<\N<	AN<=N<�NN<X{N<�N<�TO<�P<1Q<�2R<�GS<L T<�T<LT<��S<��R<�nQ<iP<��O<� O<L�N<soN<tYN<�YN<LpN<i�N<��N<ڏO<�_P<�cQ<��R<n�S<<ZT<�T<nTT<��S<�yR<�]Q<�]P<!�O<�O<n�N<,N<�jN<lN<��N<��N<qO<�O<��P<��Q<�R<ܱS<gT<t�T<�-T<3RS<�=R<!$Q<�,P<
mO<��N<8�N<�sN<�dN<�jN<��N<*�N<�.O<��O<��P<%�Q<��R<��S<�|T<C�T<�T<�*S<>R<�P<�P<QWO<0�N<y�N<�rN<�fN<&pN<e�N<��N<PFO<x�O<��P<�Q<�S<j�S<)�T<��T<	�S<��R<�Q<��P<��O<�:O<-�N<��N<{iN<�`N<�mN<��N<6�N<2XO<�P<�Q<R<�1S<AT<�T<^oT<��S<��R<��Q<h�P<+�O<X"O<��N<'�N<|gN<�cN<�tN<5�N<�N<�xO<v<P<7Q<�QR<}dS<�:T<��T<�aT<��S<њR<�{Q<SsP<��O<�O<��N<�mN<�TN<*RN<�eN<��N<��N<:|O<NIP<�JQ<fR<�rS<�8T<4T<f.T<[`S<�OR<�1Q<�0P<�dO<q�N<�N< ON<�:N<V<N<wTN<�N<��N<�O<\P<�dQ<�R<��S<�;T<eiT<� T<$S<R<�P<��O<�8O<%�N<�fN<L<N<�,N<d2N<_ON<��N<��N<]�O<�|P<��Q<��R<T�S<XFT<P[T<I�S<V�R<��Q<.�P<��O<?O<J�N<YN<4N<c(N<2N<TN<Z�N<wO<�O<�P<�  �  �-S<\T<^bT<;�S<7�R<�pQ<�O<ֿN<�N<b�M<xWN<�O<��O<�CP<�kP<.P<"�O<�N<	:N<��M<�-N<��N< GP<%�Q<�9S<c*T<�iT<8�S<��R<r�Q<5�O<�bN<}�L<��K<�GK<+K<��K<huL<��M<WHO<��P<�kR<C�S<{YT<�nT<1�S<R�R<8Q<�O<3�N<�N<�,N<��N<�oO<{P<8�P<w�P<�1P<��O<��N<�DN<(&N<�N<��O<��P<��R<��S<��T<!�T<��S<G�R</?Q<��O<�N<2�L<��K<�\K<SjK<��K<� M<caN<C�O<m�Q<]�R<6
T<ƍT<�cT<�S<H%R<��P<MKO<�mN<S"N<�_N<m�N<��O<�XP<
�P<օP<P<VVO<<�N<�0N<�<N<��N<$�O<QyQ<X�R<ET<H�T<[T<��S<q;R<D�P<XO<,�M<%aL<��K<PK<׊K<�DL<9nM<��N<��P<�R<�cS<IT<�T</.T<�S<	�Q<�#P<��N<KDN<b(N<�N<�=O<��O<*yP<��P<RbP<]�O<O<XjN<RN<�ZN<n(O<pP<��Q<�_S<|OT<�T<DT<�S<��Q<�P<��N<�M<�L<nK<7QK<��K<ԚL<+�M<�kO<�	Q<�R<�S<vT<��T<�S<��R<�Q<�O<O�N<$N<4N<ضN<qO<�P<��P<P<�&P<�~O<3�N<1N<�N<�{N<�vO<[�P<~bR<u�S<�aT<BaT<ʹS<܏R<YQ<�sO<�M<ВL<'�K< -K< ;K<��K<��L<�3N<��O<UbQ<��R<��S<WbT<�7T<�YS<��Q<�nP<O<<N<��M<�*N< �N<:�O<� P<1iP<�LP<	�O<�O<�gN<�M<�N<M�N<��O<4CQ<�R<��S<^T<�"T<�KS<AR<tP<�N<&XM<�#L<�[K<aK<�MK<�L<�2M<ܪN<�GP<��Q<�  �  jCS<��S<�S<�(R<�P<��M<=�K<�J<�sJ<�0K</�L<�N<�?P<GjQ<�Q<*9Q<:�O<ZN<NL<y�J<8mJ<��J<FL<�WN<�P<�R<ѶS<�S<=S<nQ<NBO<I�L<��J<�H<�G<��G<�=H<��I<��K<�9N<�P<�tR<�S<�S<�AS<T�Q<asO<�:M<��K<ܞJ<}�J<A�K<lM<�IO<#�P<��Q<��Q<�Q<X�O<��M<�K<��J<,�J<�rK<%M<TNO<~�Q<X@S<T<��S<��R<��P<R�N<jDL<J<�H<i�G<��G<m�H<��J<p�L<�(O<�^Q<�S<�S<��S<p�R<&	Q<�N<;�L<-K<�J<jK<TTL<�N<��O<�TQ<��Q<��Q<ѢP<��N<�M<p�K<ͳJ<��J<h�K<z�M<\P<�)R<��S<�T<�S< 6R<0P<��M<|K<PI<�+H<A�G<�H<�OI<=K<��M<|�O<�R<�xS<OT<e�S<�[R<kMP<XN<�L<O�J<��J<1eK<Z�L<��N<�uP<U�Q<��Q<EnQ<RP<ON<-L<�$K<��J<&K<�oL<�N<��P<n�R<��S<OT<V1S<>�Q<�fO<M<̾J<�H<��G<\�G<cH<��I<�K<!]N<��P<�R<��S<iT<�[S<�Q<��O<mMM<h�K<ګJ<��J<x�K<UpM<5KO<n�P<��Q<?�Q<��P<�vO<�M<��K<~�J<
�J<�VK<��L<^-O<)fQ<�S<��S<-�S<l�R<+�P<�{N<�L<�I<�[H<(�G<��G<�H<�[J<(�L< �N<z2Q<��R<��S<9�S<N�R<=�P<�N<�wL<6�J<�kJ<I�J<�L<��M<x�O<�Q<5�Q<�~Q<.iP<��N<��L<fRK<s|J<��J<"�K<t�M<U�O<V�Q<$dS<�S<j^S<z�Q<��O<\�M<�?K<�BI<��G<ipG<W�G<KI<`K<DVM<T�O<��Q<�  �  1jR<[�R<޳Q<݄O<ҜL<?�I<�XG<�-F<{cF<��G<8kJ<�XM<wP<��Q<]R<D�Q<P|O<��L<5�I<�{G<�;F<�VF<A�G<!NJ<�QM<P<R<A�R<59R<�xP<��M<��J<��G<f�E<�#D<��C<��D<*�F<�I<�L<�mO<�Q<��R<��R<�0Q<��N<!�K<��H<��F<�8F<��F<��H<�K<�sN<��P<qRR<�gR<�#Q<B�N<��K<Z!I<�G<NF<�F<p�H<m{K<[�N<FQ<�R<1�R<��Q<��O<cM<�J<<;G<�$E<D<V8D<��E<��G<x�J<;�M<{`P<~=R<w�R<qbR<��P<�M<y�J<�4H<a�F< ^F<�{G<9�I<L�L<�kO<�Q<��R<.R<-�P<h�M<��J<�^H<�F<�WF<x\G<��I<lyL<RlO<U�Q<��R<иR<�TQ<�N<r
L<I<�jF<ԦD<��C</�D<B,F<9�H<$�K<X�N<�Q<\�R<y�R<(�Q<��O<P�L<��I<��G<caF<��F<�H<�J<ώM<<P<�
R<��R<�Q<(�O<�L<J<��G<�iF<�F<|�G<�vJ<�xM<�DP<9R<��R<g]R<�P<7N<P K< H<��E<ID<(D<��D<��F<�I<жL<�O<˼Q<��R<��R<}JQ<%�N<�K<�H<f�F<�EF<��F<�H<M�K<$uN<��P<�MR<�_R<�Q<��N<
�K<�I<?G<5F<Z�F<�H<�ZK<1_N<��P<�R<��R<$�Q<z�O<�L<x�I<�G<��D<�C<�	D<oUE<֛G<W�J<��M<o4P<�R<��R<�6R<$aP<٤M<�J< H<�mF<+F<GG<�I<�]L<�2O<CZQ<�UR<��Q<FP<��M<лJ<Y&H<�~F<!F<.&G<�YI<�CL<I6O<ـQ<өR<̀R<�Q<3�N<��K<��H<�.F<�jD<��C<wID<@�E<-zH<=zK<�qN<i�P<�  �  �4Q<�9Q<��O<�L<�MI<"�E<
HC<s%B<"�B<�D<'$H<��K<�lO<^�Q<7}R<�cQ<��N<K<WG<)=D<�oB<�EB<x�C<�F<t%J<M<�1P<�fQ<�	Q<:O<sUL<�H<9yE<�B<�A<k�@<�A<�%D<�WG<��J<�N<	oP<&{Q<�P<-�N<��K<�5H<��D<%�B<�DB<]`C<��E<|�I<XM<&�P<�aR<�|R<��P<��M<ZJ<>bF<ܩC<cB<�B<~�D<c�G<��K<S�N<��P<�Q<��P<V�N<<hK<��G<�D<Z3B<��@<�A<�B<JE<�H<� L<�O<�Q<A�Q<Z�P<yN<*�J<�#G<g3D<��B<��B<4+D<�(G<�J<��N</cQ<��R<@-R<^�O<��L<�H<]E<C<pUB<�HC<��E<3I<�L<Q�O<�UQ<R~Q<A"P<��M<F8J<U�F<��C<?�A<1�@<�xA<�gC<2[F<�I<d4M<��O<piQ<�mQ<��O<�M<�I<�F<{C<YB<��B<bE<;ZH<w*L<�O<��Q<=�R<-�Q<��N<PK<��G<�mD<t�B<UrB<�C<��F<�LJ<��M<�VP<��Q<�-Q<8^O<�yL<�I<�E<�B<33A<��@<��A<�ID<q{G<Z�J<5N<��P<��Q<�Q<�O<��K<�JH<0E<��B<�QB<\jC<�E<��I<UYM<h�P<�\R<IuR<;�P<D�M<��I<�NF<��C<"JB<ԮB<@�D<��G<�iK<�N<��P<�}Q<�P<aaN</;K<�G<�tD<�B<��@<.�@<�tB<�E<zH<<�K<��N<��P<mQ<QdP<��M<��J<$�F<7D</ZB<TB<��C<��F<ԭJ<�[N< )Q<�sR<{�Q<��O<�^L<��H<~$E<M�B<�B<mC<��E<}�H<7xL<kO<�Q<�FQ<��O<SM< �I<\F<LuC<�dA<��@<�=A<Q-C<�!F<��I<"�L<ۯO<�  �  �1P<�P<($N<-�J<7�F<�5C<}@<�`?<v @<p�B<�tF<z�J<a�N<��Q<�mR<�#Q<AN<G�I<ǈE<��A<��?<�{?<��@<hD<��G<�K<��N<@P<OP<Q7N<�'K<qG<��C<��@<K�><��><�?<UB<��E<�I</M<3uO<8lP<�O<8JM<��I<��E<qEB<W@<ƌ?<0�@<��C<FH<�lL<�P<�FR<�fR<3uP<?�L<R�H<hD<�>A<(�?<��?<$B<gqE<'kI<�M<��O<��P<��O<�M<�%J<B]F<��B<m6@<��><�?<~�@<��C<@.G<+�J<6N<9P<+yP<�$O<�LL<t�H<Q�D<qA<��?<��?<Q�A<�KE<��I<�M<�Q< �R<R<�wO< �K<�'G<�9C<�@<��?<*|@<�C<�F<k�J<
N<�P<�wP<6&O<apL<��H<�E<s�A<��?<�><"m?<��A<�D<�rH<�L<'�N<�fP<�7P<5WN<�K<�'G<�hC<7�@<��?<U@<��B<�F<|K<�O<!�Q<�R<lZQ<	BN<�J<��E<�$B<��?<��?<y(A<�+D<
H<2�K<��N<�dP<�0P<�[N<�KK<��G<��C<��@<g"?<��><��?<KyB<&�E<k�I<=#M<��O<�P<��O<�cM<��I<��E<�WB<�@<��?<$�@<��C<oH<�mL<�P<�AR<�^R<�jP<��L<̓H<�TD<�(A<4�?</�?<��A<�PE<2HI<��L<�wO<�iP<W�O<6TM<��I<�/F<��B<�@<��><h�><��@<`C<OG<��J<0�M<m�O<YMP<��N<�L<�RH<bgD<�@A<�?<)�?<ȠA<wE<m_I<\�M<!�P<cR<�Q<�<O<�RK<+�F<� C<9R@<�]?<�E@<�B<y�F<�xJ<u�M<��O<�@P<��N<@7L<	�H<
�D<W�A<_\?<ǅ><I2?<sJA<�zD<�:H<��K<S�N<�  �  ��O<O�O<H�M<k/J<%F<�DB<�?<f><"6?<�A<��E<"kJ<v�N<��Q<�aR<�Q<*�M<sfI<��D<� A<p�><>><�@<"C<zG<K</N<��O<��O<��M<U�J<?�F<J'C< @<�D><m�=<�?<ȯA<�6E< I<��L<\O<�P<�+O<�L<Z�H<��D<�NA<??<ϕ><
@<3C<�}G<1L<��O<�6R<:XR<`MP<�L<�H<�C<a@<Ѻ><��><�A<Z�D<8�H<�oL<O<(P<�lO<M<ìI<��E<�5B<C�?<�'><�R><9�?<��B<�F<�wJ<@�M<c�O<[
P<��N<�K<�G<��C<lv@<y�><��><��@<��D<�I<��M<��P<��R<��Q<BO<i&K<f�F<�sB<��?<ʚ><c~?<�B<��E<��I<�rM<�O<oP<�N<�L<2_H<��D<*A<"�><r><��><X�@<�D<��G<�K<��N<�P<	�O<N�M<bJ<�OF<xwB<�?<�><�j?<�B<]F<=�J<�N<b�Q</�R<�=Q<�M<�I<�E<�QA<z?<;�><�,@<R?C<9G<l6K<nTN<}�O<��O<��M<��J<�G<LC<?@<�i><i><gC?<��A<$ZE<P9I<��L<�4O<8!P<eGO<��L<�I<w�D<aA<�?<��><�@<':C<#�G<fL<��O<�1R<�PR<�BP<y�L<�G<��C<�J@<�><2�><��@<�lD<J�H<�JL<��N<?�O<_BO<W�L<�I<�E<�B<�T?<�=<G$><H�?<V�B<xF<`KJ<;�M<��O<��O<ioN<uK<T�G<�}C<�E@<P�><��><2�@<IfD<��H<�RM<�P<�VR<��Q<+O<	�J<�TF<	;B<�j?<�c><H?<��A<a�E<:�I<�<M<wgO<#�O<ލN<��K<[%H<4JD<�@<�><T�=<{><G�@<��C<��G<nK<�QN<�  �  �1P<�P<($N<-�J<7�F<�5C<}@<�`?<v @<p�B<�tF<z�J<a�N<��Q<�mR<�#Q<AN<G�I<ǈE<��A<��?<�{?<��@<hD<��G<�K<��N<@P<OP<Q7N<�'K<qG<��C<��@<K�><��><�?<UB<��E<�I</M<3uO<8lP<�O<8JM<��I<��E<qEB<W@<ƌ?<0�@<��C<FH<�lL<�P<�FR<�fR<3uP<?�L<R�H<hD<�>A<(�?<��?<$B<gqE<'kI<�M<��O<��P<��O<�M<�%J<B]F<��B<m6@<��><�?<~�@<��C<@.G<+�J<6N<9P<+yP<�$O<�LL<t�H<Q�D<qA<��?<��?<Q�A<�KE<��I<�M<�Q< �R<R<�wO< �K<�'G<�9C<�@<��?<*|@<�C<�F<k�J<
N<�P<�wP<6&O<apL<��H<�E<s�A<��?<�><"m?<��A<�D<�rH<�L<'�N<�fP<�7P<5WN<�K<�'G<�hC<7�@<��?<U@<��B<�F<|K<�O<!�Q<�R<lZQ<	BN<�J<��E<�$B<��?<��?<y(A<�+D<
H<2�K<��N<�dP<�0P<�[N<�KK<��G<��C<��@<g"?<��><��?<KyB<&�E<k�I<=#M<��O<�P<��O<�cM<��I<��E<�WB<�@<��?<$�@<��C<oH<�mL<�P<�AR<�^R<�jP<��L<̓H<�TD<�(A<4�?</�?<��A<�PE<2HI<��L<�wO<�iP<W�O<6TM<��I<�/F<��B<�@<��><h�><��@<`C<OG<��J<0�M<m�O<YMP<��N<�L<�RH<bgD<�@A<�?<)�?<ȠA<wE<m_I<\�M<!�P<cR<�Q<�<O<�RK<+�F<� C<9R@<�]?<�E@<�B<y�F<�xJ<u�M<��O<�@P<��N<@7L<	�H<
�D<W�A<_\?<ǅ><I2?<sJA<�zD<�:H<��K<S�N<�  �  �4Q<�9Q<��O<�L<�MI<"�E<
HC<s%B<"�B<�D<'$H<��K<�lO<^�Q<7}R<�cQ<��N<K<WG<)=D<�oB<�EB<x�C<�F<t%J<M<�1P<�fQ<�	Q<:O<sUL<�H<9yE<�B<�A<k�@<�A<�%D<�WG<��J<�N<	oP<&{Q<�P<-�N<��K<�5H<��D<%�B<�DB<]`C<��E<|�I<XM<&�P<�aR<�|R<��P<��M<ZJ<>bF<ܩC<cB<�B<~�D<c�G<��K<S�N<��P<�Q<��P<V�N<<hK<��G<�D<Z3B<��@<�A<�B<JE<�H<� L<�O<�Q<A�Q<Z�P<yN<*�J<�#G<g3D<��B<��B<4+D<�(G<�J<��N</cQ<��R<@-R<^�O<��L<�H<]E<C<pUB<�HC<��E<3I<�L<Q�O<�UQ<R~Q<A"P<��M<F8J<U�F<��C<?�A<1�@<�xA<�gC<2[F<�I<d4M<��O<piQ<�mQ<��O<�M<�I<�F<{C<YB<��B<bE<;ZH<w*L<�O<��Q<=�R<-�Q<��N<PK<��G<�mD<t�B<UrB<�C<��F<�LJ<��M<�VP<��Q<�-Q<8^O<�yL<�I<�E<�B<33A<��@<��A<�ID<q{G<Z�J<5N<��P<��Q<�Q<�O<��K<�JH<0E<��B<�QB<\jC<�E<��I<UYM<h�P<�\R<IuR<;�P<D�M<��I<�NF<��C<"JB<ԮB<@�D<��G<�iK<�N<��P<�}Q<�P<aaN</;K<�G<�tD<�B<��@<.�@<�tB<�E<zH<<�K<��N<��P<mQ<QdP<��M<��J<$�F<7D</ZB<TB<��C<��F<ԭJ<�[N< )Q<�sR<{�Q<��O<�^L<��H<~$E<M�B<�B<mC<��E<}�H<7xL<kO<�Q<�FQ<��O<SM< �I<\F<LuC<�dA<��@<�=A<Q-C<�!F<��I<"�L<ۯO<�  �  1jR<[�R<޳Q<݄O<ҜL<?�I<�XG<�-F<{cF<��G<8kJ<�XM<wP<��Q<]R<D�Q<P|O<��L<5�I<�{G<�;F<�VF<A�G<!NJ<�QM<P<R<A�R<59R<�xP<��M<��J<��G<f�E<�#D<��C<��D<*�F<�I<�L<�mO<�Q<��R<��R<�0Q<��N<!�K<��H<��F<�8F<��F<��H<�K<�sN<��P<qRR<�gR<�#Q<B�N<��K<Z!I<�G<NF<�F<p�H<m{K<[�N<FQ<�R<1�R<��Q<��O<cM<�J<<;G<�$E<D<V8D<��E<��G<x�J<;�M<{`P<~=R<w�R<qbR<��P<�M<y�J<�4H<a�F< ^F<�{G<9�I<L�L<�kO<�Q<��R<.R<-�P<h�M<��J<�^H<�F<�WF<x\G<��I<lyL<RlO<U�Q<��R<иR<�TQ<�N<r
L<I<�jF<ԦD<��C</�D<B,F<9�H<$�K<X�N<�Q<\�R<y�R<(�Q<��O<P�L<��I<��G<caF<��F<�H<�J<ώM<<P<�
R<��R<�Q<(�O<�L<J<��G<�iF<�F<|�G<�vJ<�xM<�DP<9R<��R<g]R<�P<7N<P K< H<��E<ID<(D<��D<��F<�I<жL<�O<˼Q<��R<��R<}JQ<%�N<�K<�H<f�F<�EF<��F<�H<M�K<$uN<��P<�MR<�_R<�Q<��N<
�K<�I<?G<5F<Z�F<�H<�ZK<1_N<��P<�R<��R<$�Q<z�O<�L<x�I<�G<��D<�C<�	D<oUE<֛G<W�J<��M<o4P<�R<��R<�6R<$aP<٤M<�J< H<�mF<+F<GG<�I<�]L<�2O<CZQ<�UR<��Q<FP<��M<лJ<Y&H<�~F<!F<.&G<�YI<�CL<I6O<ـQ<өR<̀R<�Q<3�N<��K<��H<�.F<�jD<��C<wID<@�E<-zH<=zK<�qN<i�P<�  �  jCS<��S<�S<�(R<�P<��M<=�K<�J<�sJ<�0K</�L<�N<�?P<GjQ<�Q<*9Q<:�O<ZN<NL<y�J<8mJ<��J<FL<�WN<�P<�R<ѶS<�S<=S<nQ<NBO<I�L<��J<�H<�G<��G<�=H<��I<��K<�9N<�P<�tR<�S<�S<�AS<T�Q<asO<�:M<��K<ܞJ<}�J<A�K<lM<�IO<#�P<��Q<��Q<�Q<X�O<��M<�K<��J<,�J<�rK<%M<TNO<~�Q<X@S<T<��S<��R<��P<R�N<jDL<J<�H<i�G<��G<m�H<��J<p�L<�(O<�^Q<�S<�S<��S<p�R<&	Q<�N<;�L<-K<�J<jK<TTL<�N<��O<�TQ<��Q<��Q<ѢP<��N<�M<p�K<ͳJ<��J<h�K<z�M<\P<�)R<��S<�T<�S< 6R<0P<��M<|K<PI<�+H<A�G<�H<�OI<=K<��M<|�O<�R<�xS<OT<e�S<�[R<kMP<XN<�L<O�J<��J<1eK<Z�L<��N<�uP<U�Q<��Q<EnQ<RP<ON<-L<�$K<��J<&K<�oL<�N<��P<n�R<��S<OT<V1S<>�Q<�fO<M<̾J<�H<��G<\�G<cH<��I<�K<!]N<��P<�R<��S<iT<�[S<�Q<��O<mMM<h�K<ګJ<��J<x�K<UpM<5KO<n�P<��Q<?�Q<��P<�vO<�M<��K<~�J<
�J<�VK<��L<^-O<)fQ<�S<��S<-�S<l�R<+�P<�{N<�L<�I<�[H<(�G<��G<�H<�[J<(�L< �N<z2Q<��R<��S<9�S<N�R<=�P<�N<�wL<6�J<�kJ<I�J<�L<��M<x�O<�Q<5�Q<�~Q<.iP<��N<��L<fRK<s|J<��J<"�K<t�M<U�O<V�Q<$dS<�S<j^S<z�Q<��O<\�M<�?K<�BI<��G<ipG<W�G<KI<`K<DVM<T�O<��Q<�  �  �-S<\T<^bT<;�S<7�R<�pQ<�O<ֿN<�N<b�M<xWN<�O<��O<�CP<�kP<.P<"�O<�N<	:N<��M<�-N<��N< GP<%�Q<�9S<c*T<�iT<8�S<��R<r�Q<5�O<�bN<}�L<��K<�GK<+K<��K<huL<��M<WHO<��P<�kR<C�S<{YT<�nT<1�S<R�R<8Q<�O<3�N<�N<�,N<��N<�oO<{P<8�P<w�P<�1P<��O<��N<�DN<(&N<�N<��O<��P<��R<��S<��T<!�T<��S<G�R</?Q<��O<�N<2�L<��K<�\K<SjK<��K<� M<caN<C�O<m�Q<]�R<6
T<ƍT<�cT<�S<H%R<��P<MKO<�mN<S"N<�_N<m�N<��O<�XP<
�P<օP<P<VVO<<�N<�0N<�<N<��N<$�O<QyQ<X�R<ET<H�T<[T<��S<q;R<D�P<XO<,�M<%aL<��K<PK<׊K<�DL<9nM<��N<��P<�R<�cS<IT<�T</.T<�S<	�Q<�#P<��N<KDN<b(N<�N<�=O<��O<*yP<��P<RbP<]�O<O<XjN<RN<�ZN<n(O<pP<��Q<�_S<|OT<�T<DT<�S<��Q<�P<��N<�M<�L<nK<7QK<��K<ԚL<+�M<�kO<�	Q<�R<�S<vT<��T<�S<��R<�Q<�O<O�N<$N<4N<ضN<qO<�P<��P<P<�&P<�~O<3�N<1N<�N<�{N<�vO<[�P<~bR<u�S<�aT<BaT<ʹS<܏R<YQ<�sO<�M<ВL<'�K< -K< ;K<��K<��L<�3N<��O<UbQ<��R<��S<WbT<�7T<�YS<��Q<�nP<O<<N<��M<�*N< �N<:�O<� P<1iP<�LP<	�O<�O<�gN<�M<�N<M�N<��O<4CQ<�R<��S<^T<�"T<�KS<AR<tP<�N<&XM<�#L<�[K<aK<�MK<�L<�2M<ܪN<�GP<��Q<�  �  ��Q<|�R<|�S<VT<RT<ƽS<��R<x�Q<�P<H�O<�O<ݖN< UN<5N<�,N<B:N<FaN<<�N<�(O<�O<��P<�Q<1	S<k�S<�gT<�JT<��S<+�R<��Q<C{P<��O<3�N<��N<\N<	AN<=N<�NN<X{N<�N<�TO<�P<1Q<�2R<�GS<L T<�T<LT<��S<��R<�nQ<iP<��O<� O<L�N<soN<tYN<�YN<LpN<i�N<��N<ڏO<�_P<�cQ<��R<n�S<<ZT<�T<nTT<��S<�yR<�]Q<�]P<!�O<�O<n�N<,N<�jN<lN<��N<��N<qO<�O<��P<��Q<�R<ܱS<gT<t�T<�-T<3RS<�=R<!$Q<�,P<
mO<��N<8�N<�sN<�dN<�jN<��N<*�N<�.O<��O<��P<%�Q<��R<��S<�|T<C�T<�T<�*S<>R<�P<�P<QWO<0�N<y�N<�rN<�fN<&pN<e�N<��N<PFO<x�O<��P<�Q<�S<j�S<)�T<��T<	�S<��R<�Q<��P<��O<�:O<-�N<��N<{iN<�`N<�mN<��N<6�N<2XO<�P<�Q<R<�1S<AT<�T<^oT<��S<��R<��Q<h�P<+�O<X"O<��N<'�N<|gN<�cN<�tN<5�N<�N<�xO<v<P<7Q<�QR<}dS<�:T<��T<�aT<��S<њR<�{Q<SsP<��O<�O<��N<�mN<�TN<*RN<�eN<��N<��N<:|O<NIP<�JQ<fR<�rS<�8T<4T<f.T<[`S<�OR<�1Q<�0P<�dO<q�N<�N< ON<�:N<V<N<wTN<�N<��N<�O<\P<�dQ<�R<��S<�;T<eiT<� T<$S<R<�P<��O<�8O<%�N<�fN<L<N<�,N<d2N<_ON<��N<��N<]�O<�|P<��Q<��R<T�S<XFT<P[T<I�S<V�R<��Q<.�P<��O<?O<J�N<YN<4N<c(N<2N<TN<Z�N<wO<�O<�P<�  �  �N<�P<�Q<��R<T<dcT<�T<HS<��Q<a3P<��N<E#M<��K<KK<~K<�hK<N7L<rqM<��N<��P<�R<�bS<�2T<�dT<��S<g�R<�7Q<��O<~�N<�N<]	N<�~N<�6O<��O<�`P<�wP<�*P<�O<��N<C7N<�N<�XN<�?O<b�P<t#R<��S<TVT<wT<��S<��R<.fQ<�O< :N<v�L<��K<~TK<�NK<��K<u�L<�N<�O<�JQ<��R<�S<��T<V�T<H�S<8qR<��P<��O<��N<0N<�WN<��N<K�O<�IP<��P<$�P<�'P<�wO<f�N<�:N<	/N<��N<��O<�3Q<��R<��S<�T<�kT<'�S<�sR<z�P<RO<��M<4�L<��K<vPK<�uK<L<5M<$�N<W;P<[�Q<�2S<�-T<�T<JNT<7VS<��Q<{cP<b!O<H[N<�'N<8yN<�"O<�O<�nP<<�P<�yP<��O<t7O<�N<�)N<�LN<�O<79P<�Q<�/S<�8T<��T<�>T<QS<�Q<MfP<��N<�VM<�2L<�~K<�JK<�K<�hL<��M<M!O<O�P<�GR<݋S<HZT<�T<�T<��R<�[Q<��O<<�N<�1N<
.N<�N<�\O<7P<m�P<�P<oQP<δO<p�N<�[N<�%N< zN<Z_O<��P<T>R<�S<lT<"�T<��S<�R<�pQ<��O<p>N<��L<��K<�OK<�FK<�K<��L<
N<m�O<a4Q<F�R<��S<�jT<�^T<S�S<�JR<�P<�^O<�hN<kN<�(N<�N<wO<�P<@qP<eP<f�O<�HO<��N<�N<�N<5�N<��O<	Q<{�R<A�S<r\T<>T<A~S<�CR<��P<�O<)�M<dTL<�xK<#K<>K<Y�K<s�L<�jN<aP<��Q<V�R<��S<�`T<�T<�S<��Q<K*P<�N<�N<�M<O;N<�N<��O<8/P<�gP<�:P<��O<�N<WLN<��M<�N<�  �  ;�J<p�K<��M<�:P<�AR<�S<��S<�5S<ٳQ<O�O<�6M<��J<WI<��G<�uG<QH<<`I<CeK<��M<cP<#R<�sS<�S<X^S<�Q<��O<~M<էK<b�J<ɎJ<�qK<+M<3�N<��P<;�Q<=�Q<Q<��O<5�M<�L<Z�J<�J<= K<��L<q�N<Q<w�R<o�S<*�S<��R<�/Q<��N<�L<[J<��H<Y�G<�G<��H<�*J<XL<g�N<]Q<��R<��S<]T<�+S<mQ<�0O<�M<�hK<��J<�J<�L<d�M<�O<)+Q<��Q<��Q<!�P<�BO<sdM<��K<��J<��J<d�K<kM<��O<��Q<�hS<>T<��S<�yR<��P<�7N<2�K<g�I<MSH<��G<*�G<�I<f�J<�(M<8�O<��Q<QIS<�T<��S<��R< �P<�gN<�^L<	K<��J<�:K<Y�L<qN<9P<%�Q<	R<��Q<'eP<ťN<��L<rXK<�J<}�J<(,L<&N<)nP<qtR<��S<�T<hgS<��Q<��O<�iM<�K<U4I<�H<Y�G<�2H<ŐI<y�K<��M<bHP<fFR<�S< T< �S<�R<l�O<�M<8�K<�J<�J<N�K<�+M<\	O<D�P<c�Q<��Q<�DQ<��O<$N<�?L<�K<��J<�?K<|�L<��N<�)Q<m�R<��S<��S<.�R<%:Q<z�N<f�L<�\J<��H<��G<g�G<ǁH<�J<IGL<��N<��P<�R<d�S<P�S<A
S<�HQ<
O<��L<@>K<�J<(�J<��K<Z�M<M}O<S�P<��Q<G�Q<d�P<�O<r6M<ԓK<W�J<��J<}{K<[@M<�|O<��Q<�<S<<�S<T�S<�IR<�YP<�N<H�K<W�I<TH<WyG<'�G<��H<P�J<��L<�VO<=}Q<S<y�S<y�S<pR<gxP<&/N<�$L<�J<pgJ<\�J<�_L<1N<��O<�AQ<��Q<�ZQ<A&P<hN<��L<�K< nJ<�  �  �3F<�qG<��I<M�L<��O<��Q<4�R<^R<)�P<}LN<�QK<CUH<��E<%>D<��C<��D<tTF<��H<5L<I�N< >Q<G�R<-�R<�oQ<yO<�!L<�>I<$G<�(F<��F<-SH<��J<�M<�tP<R<aR<�SQ<gO<�EL<SoI<JBG<>9F<��F<�9H<y�J<��M<|�P<y_R<s�R<eR<�,P<~yM<pqJ<t�G<�XE<mD<�D<�,E<�PG<O&J<[3M<:�O<PR<r�R<f�R<J�P<!ZN<�TK< �H<�F<�ZF<Q@G<1SI<ML<�O<�OQ<<�R<�YR<��P<�^N<pK<e�H<A�F<�KF<G<�I<W�K<�N<xbQ<��R<��R<*�Q<�eO<%�L<I<�F<��D<mD<nWD<T�E<�;H<20K<-1N<S�P<^tR<��R<,R<�(P<.UM<�UJ<��G<�F<�zF< �G<X/J<CM<u�O<^�Q<l�R<��Q<�P<�iM<}J<	H<h�F<�kF<��G<vJ<��L<)�O<��Q<��R<��R<��P<z~N<�K<��H</	F<JpD<[�C<}�D<A�F<(I<*.L<�O<�gQ<=�R<��R<�Q<�<O<IEL<�aI<Y=G<ELF<��F<�wH<5K<nN<��P<�9R<��R<{Q<}FO<�kL<��I<fG<<[F<��F<ZWH<��J<��M<��P<�rR<��R<�$R<V7P<�M<�uJ<�G<+WE<�D<+D<�!E<�BG<}J<�M<~�O<��Q<�R<9zR<y�P<�5N<�-K<wH<,�F</.F<G<�#I<��K<��N<�Q<,QR<;)R<��P<�/N<�AK<A�H<�F<1 F<J�F<=�H<��K<6�N<�6Q<�R<�R<pQ<'5O<2VL<�KI<��F<R�D<h�C<� D<��E<�H<��J<��M<)�P<E>R<��R<��Q<��O<QM<�J<��G<hDF<�=F<�G<��I<��L<��O<-�Q<`ZR<
�Q<C�O<�+M<E@J<��G<UF<�  �  �(B<�bC<�F<��I<n	M<C�O<tEQ<N*Q<��O<��L<glI<�E<�C<�/A<ɣ@<�~A<2�C<�F<�5J<��M<ZP<�VQ<�Q<QO<�PL<��H<�`E<BC<p)B<��B<\E<�H<.�L<��O<�R<�}R<$Q<=N<F�J<R�F<
�C<�\B<�{B<�:D<Z;G<��J<�1N<�P<ÈQ<��P<�N<Q�K<WcH<�E<�sB<RA<��@<P?B<�D<�
H<��K<ӪN<U�P<y�Q<V�P<Y�N<�[K<��G<��D<)�B<�tB<��C<�F<JJ<E	N<|Q<��R<�eR<�tP<E7M<�gI<@�E<�WC<�SB<��B<
5E<{H<�L<�1O<�"Q<�Q<pP<GN<,�J<�GG<D D<��A<��@<�CA<0�B<��E<!=I<�L<��O<�CQ<s�Q<~AP<�M<B J<řF<��C<qB<R�B<�D<��G<ÍK<�$O<�Q<��R<"�Q<�}O<E�K<*H<��D<��B<�`B<�C<<;F<�I<�;M<+P<wQ<�[Q<�O<�M<<�I<(F<�?C<LaA<��@<�A<o�C<�F<gbJ<w�M<u6P<(~Q<�>Q<�uO<�tL<��H<��E<S(C<�LB<�!C<�E<��H<��L<	 P<9=R<��R<�BQ<_dN<ٯJ<��F<D<:B<�B<�XD<�VG<��J<�GN<��P<X�Q<��P<��N<��K<�gH<YE<>rB<��@<�@<�4B<�D<��G<�yK<	�N<��P<��Q<�P<k�N<7K<�G<nD<�B<	HB<�C<IpF<bJ<�M<�P<PiR<�4R<`DP<�M<�9I<
�E<�+C<L(B<��B<�
E<�PH<[�K<vO<l�P<�aQ<oAP<6�M<��J<�G<Z�C<�A<f�@<�A<��B<��E<�I<�vL<�OO<�Q<EUQ<�
P<�cM<1�I<�`F<*�C<&5B< xB<:[D<�G<�LK<]�N<.zQ<
{R<�Q<�=O<u�K<��G<�D< �B<�  �  �b?<�@<�eC<�.G<�K<0JN<�P<?)P<�N<��K<�H<�KD<#(A<�"?<�><4x?<I�A<�E<��H<�kL<BO<�NP<��O<�M<�KJ<7SF<�B< 8@<xj?< z@<<?C<�9G<��K<�{O<��Q<�kR<d�P<SxM<�2I<��D<3�A<ڲ?<��?<'zA<��D<H�H<�gL<N.O<�kP<@�O<��M<m�J<��F<�LC<�}@<��><��><�D@<8�B<+�F<�NJ<ğM<��O<��P<{�O<9�L<�4I<�?E<�A<��?<�?<oA<�D<E�H<�5M<��P<?�R<HR<*P< DL<��G<%�C<��@<�?<�1@<��B<jF<JJ<'�M<��O<'�P<�uO<��L<Y{I<H�E<FLB<��?<s�><�3?<�A<D<�G<.�K<��N<EP<�`P<5�N<i�K<�G<y D<vA<��?<$@<�VB<��E<�XJ<Y~N<ӀQ<խR<��Q<��N<�J<0sF<��B<)A@<�?<I�@<��C<bG<*NK<|N<EP<�ZP<X�N<��K<09H<?}D<�YA<,T?<�><+�?<+�A<$GE<�I<�L<;O<�uP<��O<}�M<�oJ<GvF<��B<[@<�?<4�@<"dC<^_G<+�K<�O<gR<��R<\�P<ܟM<YYI<GE<[�A<>�?<��?<B�A<S�D<X�H<�}L<�AO<w|P<��O<_�M<�J<G�F<xNC<n|@<��><��>< :@<b�B<MuF<�:J<�M<��O<oP<&bO<9�L<I<�E<��A<��?<�?<b@A<7}D<{�H<2M<�}P<�TR<R<��O<�L<I�G<�C<��@<�m?<@@<�WB<I�E<��I<"_M<٫O<UP<QGO<+�L<2JI<ԀE<�B<+�?<0�><�><��@<��C<�G<9LK<�NN<&P<�*P<��N<#�K<�G< �C<��@<dl?<��?<�B<^�E<�J<<N<�>Q<�kR<>zQ<9�N<�J<�5F<�qB<?@<�  �  )lR<�8S<��T<@W<�WY<��Z<)�Z<�Y<�W<#�T<� Q<(�M<�J<XI<��H<gI<DxK<AsN<��Q<�_U<�LX<FZ<�[<��Z<O�X<��V<�T<��R<�tR<=(S<��T<B�W<ˆZ<<]<�^<�_<��]<��[<��X<�V<��S<�R<��R<u�S<��U<DX<�Z<h
[<��Z<�mY<�V<��S<P<#�L<UJ<c�H<`�H<�!J<��L<-�O<�GS<��V<mEY<�Z<�.[<JZ<�wX<�6V<s'T<z�R<�R<��S<+�U<��X<�[<��]<�$_<��^<}]<�[<�X<"jU<�wS<�R<�S<v�T<��V<5�X<n�Z<�0[<��Z<=�X<;�U<�R<PO<��K<��I<�H<�-I<�J<��M<��P<�sT<�W<��Y<�[<��Z<��Y<�W<tU<�S<+�R<c�R<rT<��V<�Y<�{\<^x^<|>_<�^<Ϳ\<�Z<�(W<=�T<DS<T�R<�nS<4U<lsW<D�Y<a�Z<�$[<�Z< �W<!�T<�QQ<	�M<�K<�JI<P�H<�I<J�K<�N<sR<��U<�uX<smZ<�+[<�Z<Y<9�V<-�T< S<L�R<LS<<"U<�W<�Z<�:]<��^<�+_<=^<�[<�Y<�@V<YT<9�R<��R<��S<m�U<�2X<�Z<�[<`�Z<fzY<�V<ϤS<AP<m�L<aSJ<��H<��H<�J<y�L<�O<�4S<�V<�,Y<��Z<[<�)Z<�TX<V<y T<��R<L�R<խS<��U<��X<t[<ɿ]<��^<��^<�N]<�Z<��W<�=U<LS<�uR<��R<�XT<,�V<_�X<`Z<�[<�iZ<�X<ùU<�NR<��N<�K<��I<ڗH<�H<�J<�_M<u�P<~>T<}eW<c�Y<��Z<��Z<ՈY<qW<�;U<m_S<hrR<t�R<5T<�V<>Y<i<\<�8^<2�^<5`^<Ɂ\<��Y<4�V<qT<��R<�  �  �S<!�S<��U<�W<3�Y<�[<�H[<�8Z<"X<��T<��Q<h>N<��K<A�I<�8I<J<qL<�N<�SR<�U<��X<b�Z<k^[<��Z<PqY<�WW<y3U<^�S<�S<W�S<�jU<;�W<w�Z<K]<��^<��^<W�]<m�[<+!Y<zV<aT<\@S<�KS<NwT<�nV<w�X<4vZ<�i[<|0[<F�Y<�4W<
�S<͍P<dM<��J<f�I<ށI<@�J<�M<�8P<&�S<a�V<%�Y<�,[<p�[<0�Z<m�X<H�V<��T<-�S<ZS<�\T<�_V<e�X<}�[<.�]<B_<B�^<p]<%[<�[X<�U<� T<�>S<��S<�$U<|@W<xcY<�Z<��[<��Z<�Y<�>V<=�R<pO<�L<�eJ<ErI<��I<�tK<~N<-`Q<o�T<��W<�;Z<�n[<4c[<�6Z<�BX<�V<�=T<�OS<8�S<��T<�/W<��Y<J|\<�^^<�_<@�^<��\<�2Z<[xW< U<��S<�DS<�T<�U<\X<�Z<�K[<z[<jZ<65X<�*U<��Q<\oN<��K<��I<�hI<27J<�9L<�O<mR<N�U<��X<ԻZ<��[<�[<��Y<:{W<�VU<��S<k7S<'�S<F�U<	X<��Z<�0]<߻^<�_<�^<��[<nEY<@�V<̂T<l`S<�iS<a�T<��V<ݹX<�Z<|[<@[<	�Y<�>W<T<��P<UeM<+�J<׎I<dzI<ݴJ<�M<~(P<-�S<��V<�yY<|[<�n[<�Z<��X<l�V<��T<S\S<�/S<�0T<s2V<E�X<��[<�]<�^<R�^<�A]<:�Z<[.X<��U<2�S<�S<@�S<h�T<�W<�8Y<��Z<�^[<u�Z<4�X<�V<��R<�MO<-SL<�1J<�=I<؜I<�?K<8�M<�*Q<�T<G�W<SZ<9[<-[<��Y<7X<�U<iT<�S<]NS<��T<��V<�Y<!=\<G^<j�^<�D^<�~\<��Y<�<W<��T<iS<�  �  ��T<0�U<]WW<\ZY<z"[<21\<[3\<�[<�X<��U<B�R<&�O<X-M<��K<�K<L�K<�M<J[P<�}S<��V<�rY<�k[<MQ\<�\<�Z<��X<y�V<�oU<o�T<3U<��V<5�X<]�Z<��\<L/^<jp^<ǔ]<��[<T�Y<UmW<��U<�T<NU<�@V<X<�Z<:�[<=p\<�\<^�Z<KX<HU<M�Q<��N<-�L<ChK<XK<�}L<��N<�Q<��T<��W<�fZ<@
\<��\<��[<�nZ<�uX<-�V<�NU<qU<��U<7_W<��Y<�[<��]<Б^<�p^<�<]<+E[<��X<�V<>wU<��T<�xU<I�V<��X<��Z<� \<��\<�[<:�Y<�.W<	T<�P< "N<�+L<YJK<��K<[&M<�O<ߞR<��U<C�X<F[<�U\<�t\<�[<��Y<��W<
V<�U<�U<H0V<!	X<(GZ<�o\<�^<<�^<�%^<~�\<��Z<�DX<�ZV<0U<�U<��U<��W<��Y<�T[<c\<�d\<?[<=Y<�)V<y�R<Q�O<Y^M<��K<AK<� L<K�M<��P<թS<'�V<��Y<��[<�w\<A5\<��Z<_Y<�W<
�U<��T<�VU<<�V<��X<� [<�]<U^<2�^<J�]<��[<u�Y<V�W<3�U<�U<]1U<�\V<�4X<�2Z<�[<m�\<l \<�Z<4#X<VU<y�Q<��N<��L<�cK<�PK<esL<I�N<�{Q<��T<��W<"NZ<!�[<�o\<]�[<hLZ<�PX<QkV<�%U< �T<��U<!2W<�YY<o�[<�i]<�b^<�A^<M]<S[<��X<��V<}KU<��T<�MU<��V<#�X<��Z<I�[<$V\<��[<��Y<&�V<�S<��P<��M<��K<�K<�mK<�L<�bO<diR<��U<ēX<��Z< \<v>\<`J[<D�Y<��W<��U<\�T<�T<��U<x�W<�Z<�0\<��]<Pg^<_�]<�g\<[JZ<o	X<� V<��T<�  �  ZCW<L<X<�Y<܌[<A�\<�]<^p]<q.\<EZ<KjW<��T<��Q<�O<9=N<��M<�yN<�P<zqR<54U<zX<�Z<�\<R�]<m�]<��\<4[<�uY< X<L4W<F>W<�X<�lY<<[<�u\<.f]<ڕ]<��\<4�[<�%Z<E�X<��W<~(W<��W<�X<2~Z<<1\<�l]<0�]<�?]<��[<�\Y<ΚV<��S<6Q<�<O<E#N<WN<�O<��P<�S<WV<n"Y<Q�[<;5]<{�]<�]<�z\<P�Z<�Y<��W<sQW<w�W<��X<$#Z<��[< ]<��]<y�]<`�\<t[[<��Y<PYX<�tW<�RW<EX<�mY<�*[<��\<"�]<s�]<��\<�
[<�X<A�U<0�R<��P<��N<�
N<JXN<��O<J�Q<AuT<�NW<� Z<�0\<��]<o�]<FO]<��[<;6Z<0�X<��W<iOW<��W<�Y<B�Z<u0\<$T]<O�]<�j]<�V\<�Z<�AY<��W<CTW<zW<�qX<>Z<�[<�-]<��]<��]<�_\<�CZ<��W<8�T<fR<E�O<JnN<�N<��N<ZHP<#�R<�`U<c6X<w�Z<�\<	�]<��]<]�\<X[<?�Y<|#X<�WW<bW<,3X<g�Y<X)[<��\<͋]<p�]<0]<��[<sIZ<�X<�W<@HW<��W<��X<ǗZ<pH\<��]<I�]<O]<g�[<bfY<ҡV< �S<V7Q<0;O<�N<�N<GO<J�P<drS<DV<�Y<�p[<,]<��]<�]<X\<��Z<&�X<�W<.'W<�uW<�{X<V�Y<'�[<;�\<"�]<�r]<�\<�-[<��Y<�,X<$IW<|'W<l�W<�BY<��Z<��\<F�]<��]<ܶ\<��Z<�WX<�U<��R<SP<?�N<�M<�"N< uO<��Q<�?T<W<"�Y< �[<�W]<R�]<�]<G�[<�Y<aX<pSW<W<F�W<Q�X<HjZ<�[<�]<҉]<�,]<�\<ȘZ<�Y<=�W<W<�  �  ��Y<��Z<Sq\<v�]<��^<a#_<��^<�9]<�C[<K�X<��V<�aT<P�R<�jQ<�Q<"�Q<k�R<'�T<W<�Y<^�[<z�]<#�^<�+_<G�^<d�]<�%\<��Z<	�Y<�QY<�xY<�Z<}�Z<9�[<{\<4\<��[<�6[<�iZ<��Y<+[Y<I�Y<�HZ<9�[<j
]<�\^<;&_<�)_<�T^<�\<ͦZ<'MX<��U<N�S<�CR<�\Q<�QQ<6$R<ıS<g�U<�X<NvZ<�\<�F^<�5_<�L_<��^<�T]<��[<��Z<}�Y<"�Y<S�Y<;~Z<L[<1�[<_[\<N\<��[<�[<7LZ<ȭY<�wY<j�Y<��Z<�"\<��]<��^<FR_<D_<��]<�(\<��Y<ȐW<�GU<SS<.�Q<eKQ<ۊQ<7�R<�]T<ΈV<k�X<�9[<�<]<�^<�R_<�!_<%5^<�\<FZ[<?0Z<��Y<&�Y<��Y<��Z<މ[<�$\<�b\<�0\<�[<��Z<kZ<��Y<��Y<?Z<2[<g�\<�^<\_<]U_<T�^<8k]<Cu[<(Y<��V<��T<,�R<7�Q<�CQ<�Q<�S<aU<�IW<-�Y<R�[<��]<E�^<rQ_<>�^<��]<iI\<J�Z<��Y<�uY<�Y<2Z<r�Z<z�[<�?\<hY\< \<3[[<��Z<��Y<P|Y<ͤY<<fZ<ק[<�#]<�s^<�:_<�;_<)d^<��\<��Z<TX<��U<��S<�AR<KXQ<9JQ<�R<��S<S�U<�X<�`Z<��\<�+^<_<�,_<Ww^<F0]<Q�[<dZ<p�Y<�UY<��Y<�PZ<�[<��[<�,\<�\<v�[<]�Z<EZ<x�Y<'LY<+�Y<ܘZ<�[<�p]<�^<&_<-�^<��]<b�[<��Y<�^W<�U< S<h�Q<Q<UQ<7jR<v'T<�RV<��X<+[<]<Hv^<�_<^�^<�]<9�\<~![<t�Y<�UY<OMY<��Y<.�Z<�K[<��[<�$\<,�[<+a[<;�Z<��Y<UVY<'OY<�  �  �\< S]<P�^<��_<�*`<��_<�"_<��]<\<�-Z<eX<��V<t�U<k�T<�mT<��T<��U<w"W<n�X<�Z<�m\<-^<^f_<�`<�#`<�_<_d^<X]<<�[< �Z<fZ<='Z<�Z<o'Z<�3Z<�5Z<q/Z<,#Z<�"Z<mHZ<g�Z<�t[<-�\<��]<^_<Z`<\L`<��_<@�^<ZP]<͉[<K�Y<�W<>yV<�SU<�T<��T<�>U<�ZV<F�W<}�Y<f[<T3]<��^<P�_<Ne`<1`<4__<�'^<��\<߶[<��Z<�yZ<�NZ<MZ<aYZ<�`Z<D_Z<�SZ<�FZ<|MZ<��Z<I[<��[<k]<,h^<ҏ_<�B`<TQ`<!�_<�p^<�\< �Z<h,Y<��W<�V<}U<��T<�T<��U<��V<;jX<!/Z<k\<s�]<�5_<C"`<�c`<��_<K�^<�]<~i\<	c[<ݶZ<'`Z<�FZ<�MZ<�ZZ<o_Z<�[Z<�NZ<�EZ<�YZ<<�Z<J[<�F\<�]<:�^<��_<k]`<�/`<�T_<h�]<6\<`Z<p�X<j�V<�U<��T<\�T<�U<��U<ZQW<��X<,�Z<�\<7B^<��_<D`<RI`<��_<b�^<7]<� \<�[<5�Z<�KZ<�@Z<vLZ<�XZ<�ZZ<-TZ<UGZ<�EZ<�jZ<?�Z<�[<��\<�]<�8_<8`<�``<��_<u�^<�\]<��[<3�Y<-�W<nzV<�QU<m�T<�T</4U<�MV<<�W<�|Y<oP[<]<�^<��_<vE`<�`<�:_<J^<��\<�[<��Z<oMZ<p!Z<:Z<'+Z<�2Z<1Z<�%Z<[Z<� Z<JXZ<��Z<��[<Z�\<=^<�d_</`<�$`<��_<"B^</�\<��Z<�X<MW<��U<%�T<�oT<��T<�cU<�V<�3X<��Y<x�[<��]<��^<J�_<A-`<ھ_<��^<�w]<)0\<�([<�{Z<	$Z<
Z<XZ<jZ<*"Z<�Z<|Z<�
Z<�Z<xoZ<�[<�  �  :p]<��^<}�_<�}`<{y`<��_<��^<�]]<w�[<��Z<@�Y<	�X<�X<̩W<�W<��W<�8X<��X<�Y<?�Z<�K\<Ʊ]<._<`<�`<q`<$�_<�^<�,]<�[<�Z<�Y<�X<X<�W<�W<N�W<�cX<w%Y<�Z<�D[<W�\<��]<�L_<LA`<��`<Hp`<O�_<�h^<B]<��[<�xZ<�vY<��X<:X<˽W<��W<�	X<3�X<�gY<�fZ<p�[<��\<�X^<��_<�{`<��`<�t`<.�_<�K^<h�\<��[<AcZ<\hY<�X<X<�W<q�W<W*X<D�X<̕Y<��Z<I�[<�,]<&�^<��_<w�`<\�`<rN`<7U_<�^<c�\<tQ[<(-Z<�;Y<�~X<#�W<N�W<�W<�=X<p�X<��Y<��Z<�
\<�j]<g�^<i�_<c�`<R�`<1`<�%_< �]<�j\<![<�Z<�Y<�gX<��W<��W<�W<�VX<jY<��Y<�Z<|C\<�]<b _<7`<ʰ`<�`<�	`<��^<�]<�-\<�Z<�Y<�X<�IX<��W<v�W<]�W<�iX<� Y<WZ<�*[<�v\<e�]<W/_<�4`<ѵ`<�`<h�_<Ѱ^<ZP]<��[<�Z<H�Y<��X<�2X<��W<��W<� X<��X<rHY<r=Z<e[<G�\<�^<h_<GZ`<��`<��`<�_<�w^<�]<:�[<�Z<�zY<��X<�X<2�W<4�W<g�W<�X<�WY<TZ<�[<��\<�=^<]~_<�[`<��`<�P`<j_<�#^<�\<�e[<47Z<l;Y<�sX<+�W<�W<��W<��W<�X<!iY<�nZ<��[<t]<�c^<��_<�``<6�`<|!`<<'_<��]<�p\<�[<$�Y<Y<gIX<.�W<ʉW<3�W<�X<��X<��Y<��Z<��[<�4]<��^<��_<@m`<��`<��_<��^<H�]<71\<^�Z<y�Y<��X< +X<ӲW<+�W<�W<!X<��X<P�Y<��Z<w\<�  �  b�]<�1_<V`<�'`<#�_<��^<^A]<�\<I	[<�kZ<~ Z<Z<�Z<p#Z<�&Z<�!Z<�Z<Z<&-Z<k�Z<<[<�H\<��]<3�^<k�_<28`<��_<M�^<��]<��[<��Y<h)X<�V<�cU<U�T<��T<��T<�V<9uW<�%Y<V�Z<��\<}k^<�_<R>`<�'`<fm_<3B^<'�\<��[<U�Z<�mZ<:Z<V5Z<�BZ<NNZ<$PZ<�HZ<�=Z<BZ<�qZ<�Z<(�[<��\<�5^<�k_<&8`<�d`<;�_< �^<�"]<�U[<i�Y<I�W<]VV<�AU<��T<��T<rU<�V<D#X<��Y<$�[<�z]<I�^<5`<�a`<�`<!'_<'�]<��\<߄[<��Z< fZ<�DZ<`HZ<VZ<�\Z<[Z<POZ<�DZ<�RZ<�Z<�([<\<�P]<��^<�_<aU`<6F`<چ_<4^<?�\<T�Z<B�X<�BW<��U<��T<4�T<��T<&�U<W<u�X<J}Z<CR\<�^<bf_<�7`<�Z`<��_<��^<�s]<G4\<�;[<��Z<�SZ<�AZ<�JZ<�VZ<�YZ<TZ<jFZ<m@Z<\Z<ҶZ<�g[<�r\<b�]<�_<��_<g]`<c`<d_<�]<��[<�Z<�MX<]�V<L�U<��T<g�T<�#U<E+V<ݗW<9GY<�[<��\<Z�^<��_<W`<>`<{�_<�S^<  ]<��[<��Z<TtZ<>Z<u6Z<#AZ<�IZ<�HZ<{>Z<�0Z<2Z<_Z<��Z<�[<B�\<�^<7L_<U`<�@`<U�_<Q�^<��\<�*[<�UY<��W<!)V<�U<�T<B�T<�DU<qV<��W<�Y<x�[<�O]<��^<��_<6`<?�_<��^<��]<Mi\<�S[<<�Z<^2Z<�Z<�Z<�Z<�%Z<�#Z<�Z<�Z<�Z<�^Z<e�Z<�[<�]<�k^<�_<`<Z`<LO_<��]<M\<ExZ<q�X<W<�U<��T<ShT<g�T<P�U<��V<�zX<�EZ<�\<�  �  �O]<��^<#$_<��^<��]<�\\<F�Z<c�Y<�MY<4]Y<n�Y<�Z<�n[<��[<�(\<1�[<�F[<Z{Z<&�Y<�PY<�aY<[Z<=[<�\<_^<T�^<�#_<�q^<W�\<��Z<]�X<v?V<VT<dR<�ZQ<)Q<�Q<�HS<VEU<=�W<Y�Y<*\<��]<��^<J9_<B�^<�s]<a�[<'�Z<�Y<eY<)�Y<�DZ<l[<��[<@@\<�G\<��[<�1[<(eZ<i�Y<�uY<-�Y<D�Z<��[<of]<y�^<�R_<�1_<[9^<�\<�^Z<��W<_�U<��S<�!R<\Q<�tQ<TgR<�T<�'V<�X<U�Z<��\<�y^<�C_<E5_<�c^<�]<��[<�UZ<��Y<�|Y<��Y<ŘZ<�f[<�\<S]\<U>\<͹[<p�Z<-Z<Q�Y<!~Y<�Y<Z�Z<?f\<q�]<��^<�Y_<��^<O�]<�[<��Y<�/W<0�T< S<N�Q<cHQ<��Q<��R<��T<W�V<�LY<~�[<�]<'�^<�W_<�_<��]<�\<�[<Z<̀Y<��Y<=Z<6�Z<�[<�0\<E\\<H\<�x[<U�Z<��Y<�~Y<�Y<6Z<Nf[<��\<�>^<�"_<�H_<�^<Q]<�[<Q�X<�cV<�=T<ֈR<QQ<=MQ<��Q<lS<�gU<z�W<BZ<mH\<�	^<�_<�Q_<��^<��]<�\<�Z<�Y<�nY<�Y<�HZ<�[<��[<�;\<\@\<��[<q$[<:UZ<��Y<$`Y<(�Y<�zZ<��[<G]<υ^<�._<�_<�^<�_\<�4Z<O�W<�U<�xS<��Q<�.Q<7GQ<-:R<��S<*�U<UX<��Z<�\<N^<�_<+	_<�6^<��\<�b[<�%Z<;kY<
JY<��Y<`cZ<_0[<��[<�%\<k\<߁[<��Z<��Y<VfY<�GY<�Y<}�Z<�0\<��]<��^<K#_<X�^<g|]<P�[<yWY<U�V<d�T<��R<��Q<(Q<�qQ<d�R<M{T<�V<�Y<I`[<�  �  �D\<�y]<9�]<��\<u[<�Y<�*X<=W<J"W<;�W<�Y<ɲZ<N0\<D;]<N�]<K]<M�[<!YZ<�X<ҟW<�W<�dW<
}X<�Z<��[<1]<e�]<�U]<r�[<��Y<z�V<%T<��Q<�jO<�&N<��M<8�N<n�P<U�R<�U<ϑX<W[<6�\<r�]<��]<��\<��Z<%CY<B�W<�<W<�jW<oXX<��Y<y_[<�\<��]<�]<[�\<��[<7�Y<o�X<��W<�IW<��W<�-Y<�Z<>�\<��]<��]<�(]<�r[<�Y<9V<hS<Q�P<�O<]N<i<N<�dO<|hQ<��S<>�V<��Y<��[<ib]<`�]<�u]<:2\<�}Z<G�X<4�W<�FW<Y�W<��X<T`Z<��[<~+]<��]<P�]<�\<�[<�Y<9)X<�bW<�dW<�;X< �Y<�x[<P�\<G�]<��]<ר\<�Z<xX<0?U<'�R<D2P<d�N<�N<=�N<��O<98R<��T<��W<�hZ<�y\<��]<w�]<L]<�[<H�Y<`]X<�oW<�UW<�X<5SY<U�Z<e\<�o]<��]<�A]<\<��Z<D�X<f�W<�EW<�W<��X<�GZ<c\<�V]<\�]<Mz]<�\<��Y<c!W<IT<�Q<�O<�JN<�N<��N<T�P<bS<�U<x�X<y-[<��\<��]<��]<ˮ\<�[<zTY<�W<�HW<tW<_X<��Y<�`[<G�\<�]<i�]<�\<t�[<Q�Y<�vX<;wW<�1W<m�W<�Y<��Z<�l\<�]<	�]<�]<�I[<��X<�V<	<S<��P<��N<%�M<=N<�7O<�;Q<��S<Q�V<�gY<"�[<�6]<��]<�I]<%\<�OZ<�X<�xW<�W<��W<*�X<l*Z<��[<��\<��]<�M]<�T\<x�Z<MIY<�W<�+W<f.W<X<q�Y<�B[<o�\< �]<$�]<Rq\<�tZ<s�W<}U<�FR<��O<�dN<(�M<�FN<��O<N�Q<�T<��W<�2Z<�  �  �#[<�9\<�'\<�[<�=Y<d<W<��U<��T<�U<_:V<(+X<�mZ<�\<��]<cj^<��]<6\<��Y<��W<�U<F�T</�T<D�U<c�W<Q�Y<�g[<�N\<� \<�Z<~yX<N~U<yIR<
IO<�L<
pK<*K<�L<�"N<��P<hT<�<W<d�Y<��[<nm\<��[<�Z<e�X<`�V<�WU<��T<tU<>�V<�Y<"R[<�A]<h^<�y^<�r]<�[<�XY<6W<2�U<
�T<SU<8�V<��X<q�Z<\<,�\<o�[<�NZ<�W<`�T<lQ<o�N<ttL<�_K<��K<��L<�$O<nR<�LU<�SX<ȽZ<�1\<w�\<N�[<�Z<XX<nEV<@&U<�U<I�U<��W<<�Y<�\<�]<ќ^<tL^<��\<��Z<�X<��V<�PU<$�T<�U<E:W<58Y<�[<RH\<�z\<9�[<��Y<@�V<D�S<ZeP<�M<&�K<EK<��K<��M<3P<�'S<YV<I8Y<�X[<�m\<�Z\<3?[<TpY<�nW<G�U<��T<o7U<gnV<�_X<��Z<��\<�.^<�^<��]<fM\<�Z<8�W<V<�U<�U<9V<��W<j�Y<�[< t\<+E\<-�Z<k�X<0�U<emR<mO<M<��K<�MK<�@L<cEN<�Q<.9T<Y\W<XZ<��[<Ç\<\<��Z<�X<��V<ofU<��T<l}U<��V<�Y<,S[<@]<zc^<@r^<�h]<��[<�HY<�#W<�U<"�T<�8U<U�V<�oX<fZ<��[<�k\<R�[<A&Z<�W<WqT<8@Q<�fN<�GL<�2K<�UK<�L<"�N<<�Q<� U<�'X<=�Z<!\<�U\<Њ[<��Y<�W<�V<Y�T<��T<��U<�wW<�Y<X�[<�]<Qd^<�^<�\<>�Z<�hX<IiV<U<��T</uU<�W<�Y<��Z<@\<BD\< O[<�HY<�xV<�IS<�+P<�M<ιK<�
K<��K<BHM<��O<��R<w"V<�Y<�  �  eNZ<M[<�[<շY<{�W<��U<[�S<US<1yS<�U<eW<�Z<�\<�Y^<7�^<7^<� \<��Y<�V<��T<-JS<\"S<�!T<�U<s3X<� Z<B@[<h;[<��Y<��W<�vT<rQ<A�M<;/K<۝I<�RI<BYJ<ۉL<��O<;�R<�NV<�Y<��Z<�s[<�Z<D3Y<�W<��T<ӋS<Z/S<*T<-�U<8pX<L*[<Zy]<a�^<��^<Y�]<l{[<��X<�0V<c;T<�JS<��S<��T<��V<Y<��Z<|�[<�"[<�yY<��V<��S<
P<u M<ʳJ<�I<b�I<�K<F�M<b�P<M?T<�pW<��Y<�O[<}x[<wZ<��X<�hV<6{T<	`S<�gS<�T<�V<�lY<m\<J^<�_<#�^<w]<w�Z<L�W<�vU< �S<�>S<��S<�zU<�W<�Y<�'[<�[<P�Z<��X<��U<�UR<o�N<�L<0)J<�lI<�J<��K<��N<�Q<�\U<T]X<�Z<Ȁ[<�@[<w�Y<��W<�U<�S<s?S<լS<09U<ÙW<�TZ<A�\<�^<4_<�D^<vT\<��Y<\W<�T<�wS<2NS<�KT<�'V<�ZX<�FZ<{e[<�_[<Z<�W<ԚT<R+Q<+�M<&SK<��I<vI<r|J<k�L<��O<�S<,nV<k1Y<��Z<�[<4�Z<>IY<:!W<	U<z�S<b;S<�T<��U<tX<R+[<�w]<��^<c�^<�]<Un[<ɸX<
V<&T<�2S<%nS<��T<��V<��X<Y�Z<,m[<��Z<hQY<�V<�WS<G�O<�L<�J<,\I<{�I<��J<�qM<>�P<sT<�DW<5�Y<)$[<yL[<vJZ<BnX<D:V<}KT<�.S<5S<�eT<��V<k6Y<��[<�]<,�^<:x^<��\<�kZ<7�W<j?U<6�S<KS<��S<=EU<]mW<x�Y<��Z<�S[<FxZ<�oX<��U<{R<ڿN<��K<�I<�2I<D�I<��K<BgN<��Q<F&U<�'X<�  �  � Z<��Z<�Z<?=Y<tW<��T<�&S<WkR<��R<�T<�W<��Y<Ҧ\<4v^<�_<�(^<M\<d[Y<y}V<iT<�R<WR<�|S<jcU<ǨW<�Y<��Z<��Z<�Y<\IW<zT<��P<�AM<ڕJ<��H<��H<�I<��K<UO<��R<E�U<��X<Q�Z<�[<RdZ<�X<�xV<�UT<�R<�R<�zS<WzU<2X<K[<Շ]<b�^<�
_<��]<�l[<��X<��U<�S<��R<��R<�:T<{SV<f�X<�^Z<�5[<��Z<-Y<�zV<2 S<%�O<ZrL<�J<a�H<�	I<��J<lM<�[P<��S<yW<�Y<��Z< [<~Z<\X<��U<�S<[�R<r�R<8T<�eV<�=Y<�\<�3^<k3_<��^<�]<��Z<��W<�U<�@S<ߞR<8S<��T<�W<-;Y<D�Z<2[<4aZ<iYX<�bU<\�Q<qxN<S�K<��I<F�H<VaI<AK<ZN<z�Q<�U<�X<R5Z<y*[<#�Z<�oY<�QW<fU<�YS<~�R<�S<4�T<sLW<(4Z<;�\<��^<7_<E]^<�Q\<ōY<n�V<�NT<��R<B�R<��S<�U<�W<�Y<:[<�[<;�Y<LmW<U>T<��P<�eM<��J<�I<�H<)�I<=L<4O<Q�R<�V<Q�X<j�Z<�2[<z|Z<��X<��V<)gT<"�R<��R<�S<�U<�5X<P[<�]<��^<s_<g�]<�_[<�X<d�U<��S<��R<$�R<�T<U4V<sX<e;Z<s[<ϫZ<�Y<�PV<R�R<mpO<FL<�I<~�H<��H<�UJ<��L<�/P<�S<��V<�qY<��Z<�Z<��Y<��W<N�U<S�S</�R<ѝR<%�S<}0V<>Y<F�[<e�]<��^<��^<��\<�OZ<�gW<N�T<�	S<�hR< S<5�T<T�V<�Y<_�Z<��Z<;*Z<�!X<:*U<c�Q<�>N<|NK<�MI<d�H<�'I<�K<�M<!PQ<]�T<-�W<�  �  eNZ<M[<�[<շY<{�W<��U<[�S<US<1yS<�U<eW<�Z<�\<�Y^<7�^<7^<� \<��Y<�V<��T<-JS<\"S<�!T<�U<s3X<� Z<B@[<h;[<��Y<��W<�vT<rQ<A�M<;/K<۝I<�RI<BYJ<ۉL<��O<;�R<�NV<�Y<��Z<�s[<�Z<D3Y<�W<��T<ӋS<Z/S<*T<-�U<8pX<L*[<Zy]<a�^<��^<Y�]<l{[<��X<�0V<c;T<�JS<��S<��T<��V<Y<��Z<|�[<�"[<�yY<��V<��S<
P<u M<ʳJ<�I<b�I<�K<F�M<b�P<M?T<�pW<��Y<�O[<}x[<wZ<��X<�hV<6{T<	`S<�gS<�T<�V<�lY<m\<J^<�_<#�^<w]<w�Z<L�W<�vU< �S<�>S<��S<�zU<�W<�Y<�'[<�[<P�Z<��X<��U<�UR<o�N<�L<0)J<�lI<�J<��K<��N<�Q<�\U<T]X<�Z<Ȁ[<�@[<w�Y<��W<�U<�S<s?S<լS<09U<ÙW<�TZ<A�\<�^<4_<�D^<vT\<��Y<\W<�T<�wS<2NS<�KT<�'V<�ZX<�FZ<{e[<�_[<Z<�W<ԚT<R+Q<+�M<&SK<��I<vI<r|J<k�L<��O<�S<,nV<k1Y<��Z<�[<4�Z<>IY<:!W<	U<z�S<b;S<�T<��U<tX<R+[<�w]<��^<c�^<�]<Un[<ɸX<
V<&T<�2S<%nS<��T<��V<��X<Y�Z<,m[<��Z<hQY<�V<�WS<G�O<�L<�J<,\I<{�I<��J<�qM<>�P<sT<�DW<5�Y<)$[<yL[<vJZ<BnX<D:V<}KT<�.S<5S<�eT<��V<k6Y<��[<�]<,�^<:x^<��\<�kZ<7�W<j?U<6�S<KS<��S<=EU<]mW<x�Y<��Z<�S[<FxZ<�oX<��U<{R<ڿN<��K<�I<�2I<D�I<��K<BgN<��Q<F&U<�'X<�  �  �#[<�9\<�'\<�[<�=Y<d<W<��U<��T<�U<_:V<(+X<�mZ<�\<��]<cj^<��]<6\<��Y<��W<�U<F�T</�T<D�U<c�W<Q�Y<�g[<�N\<� \<�Z<~yX<N~U<yIR<
IO<�L<
pK<*K<�L<�"N<��P<hT<�<W<d�Y<��[<nm\<��[<�Z<e�X<`�V<�WU<��T<tU<>�V<�Y<"R[<�A]<h^<�y^<�r]<�[<�XY<6W<2�U<
�T<SU<8�V<��X<q�Z<\<,�\<o�[<�NZ<�W<`�T<lQ<o�N<ttL<�_K<��K<��L<�$O<nR<�LU<�SX<ȽZ<�1\<w�\<N�[<�Z<XX<nEV<@&U<�U<I�U<��W<<�Y<�\<�]<ќ^<tL^<��\<��Z<�X<��V<�PU<$�T<�U<E:W<58Y<�[<RH\<�z\<9�[<��Y<@�V<D�S<ZeP<�M<&�K<EK<��K<��M<3P<�'S<YV<I8Y<�X[<�m\<�Z\<3?[<TpY<�nW<G�U<��T<o7U<gnV<�_X<��Z<��\<�.^<�^<��]<fM\<�Z<8�W<V<�U<�U<9V<��W<j�Y<�[< t\<+E\<-�Z<k�X<0�U<emR<mO<M<��K<�MK<�@L<cEN<�Q<.9T<Y\W<XZ<��[<Ç\<\<��Z<�X<��V<ofU<��T<l}U<��V<�Y<,S[<@]<zc^<@r^<�h]<��[<�HY<�#W<�U<"�T<�8U<U�V<�oX<fZ<��[<�k\<R�[<A&Z<�W<WqT<8@Q<�fN<�GL<�2K<�UK<�L<"�N<<�Q<� U<�'X<=�Z<!\<�U\<Њ[<��Y<�W<�V<Y�T<��T<��U<�wW<�Y<X�[<�]<Qd^<�^<�\<>�Z<�hX<IiV<U<��T</uU<�W<�Y<��Z<@\<BD\< O[<�HY<�xV<�IS<�+P<�M<ιK<�
K<��K<BHM<��O<��R<w"V<�Y<�  �  �D\<�y]<9�]<��\<u[<�Y<�*X<=W<J"W<;�W<�Y<ɲZ<N0\<D;]<N�]<K]<M�[<!YZ<�X<ҟW<�W<�dW<
}X<�Z<��[<1]<e�]<�U]<r�[<��Y<z�V<%T<��Q<�jO<�&N<��M<8�N<n�P<U�R<�U<ϑX<W[<6�\<r�]<��]<��\<��Z<%CY<B�W<�<W<�jW<oXX<��Y<y_[<�\<��]<�]<[�\<��[<7�Y<o�X<��W<�IW<��W<�-Y<�Z<>�\<��]<��]<�(]<�r[<�Y<9V<hS<Q�P<�O<]N<i<N<�dO<|hQ<��S<>�V<��Y<��[<ib]<`�]<�u]<:2\<�}Z<G�X<4�W<�FW<Y�W<��X<T`Z<��[<~+]<��]<P�]<�\<�[<�Y<9)X<�bW<�dW<�;X< �Y<�x[<P�\<G�]<��]<ר\<�Z<xX<0?U<'�R<D2P<d�N<�N<=�N<��O<98R<��T<��W<�hZ<�y\<��]<w�]<L]<�[<H�Y<`]X<�oW<�UW<�X<5SY<U�Z<e\<�o]<��]<�A]<\<��Z<D�X<f�W<�EW<�W<��X<�GZ<c\<�V]<\�]<Mz]<�\<��Y<c!W<IT<�Q<�O<�JN<�N<��N<T�P<bS<�U<x�X<y-[<��\<��]<��]<ˮ\<�[<zTY<�W<�HW<tW<_X<��Y<�`[<G�\<�]<i�]<�\<t�[<Q�Y<�vX<;wW<�1W<m�W<�Y<��Z<�l\<�]<	�]<�]<�I[<��X<�V<	<S<��P<��N<%�M<=N<�7O<�;Q<��S<Q�V<�gY<"�[<�6]<��]<�I]<%\<�OZ<�X<�xW<�W<��W<*�X<l*Z<��[<��\<��]<�M]<�T\<x�Z<MIY<�W<�+W<f.W<X<q�Y<�B[<o�\< �]<$�]<Rq\<�tZ<s�W<}U<�FR<��O<�dN<(�M<�FN<��O<N�Q<�T<��W<�2Z<�  �  �O]<��^<#$_<��^<��]<�\\<F�Z<c�Y<�MY<4]Y<n�Y<�Z<�n[<��[<�(\<1�[<�F[<Z{Z<&�Y<�PY<�aY<[Z<=[<�\<_^<T�^<�#_<�q^<W�\<��Z<]�X<v?V<VT<dR<�ZQ<)Q<�Q<�HS<VEU<=�W<Y�Y<*\<��]<��^<J9_<B�^<�s]<a�[<'�Z<�Y<eY<)�Y<�DZ<l[<��[<@@\<�G\<��[<�1[<(eZ<i�Y<�uY<-�Y<D�Z<��[<of]<y�^<�R_<�1_<[9^<�\<�^Z<��W<_�U<��S<�!R<\Q<�tQ<TgR<�T<�'V<�X<U�Z<��\<�y^<�C_<E5_<�c^<�]<��[<�UZ<��Y<�|Y<��Y<ŘZ<�f[<�\<S]\<U>\<͹[<p�Z<-Z<Q�Y<!~Y<�Y<Z�Z<?f\<q�]<��^<�Y_<��^<O�]<�[<��Y<�/W<0�T< S<N�Q<cHQ<��Q<��R<��T<W�V<�LY<~�[<�]<'�^<�W_<�_<��]<�\<�[<Z<̀Y<��Y<=Z<6�Z<�[<�0\<E\\<H\<�x[<U�Z<��Y<�~Y<�Y<6Z<Nf[<��\<�>^<�"_<�H_<�^<Q]<�[<Q�X<�cV<�=T<ֈR<QQ<=MQ<��Q<lS<�gU<z�W<BZ<mH\<�	^<�_<�Q_<��^<��]<�\<�Z<�Y<�nY<�Y<�HZ<�[<��[<�;\<\@\<��[<q$[<:UZ<��Y<$`Y<(�Y<�zZ<��[<G]<υ^<�._<�_<�^<�_\<�4Z<O�W<�U<�xS<��Q<�.Q<7GQ<-:R<��S<*�U<UX<��Z<�\<N^<�_<+	_<�6^<��\<�b[<�%Z<;kY<
JY<��Y<`cZ<_0[<��[<�%\<k\<߁[<��Z<��Y<VfY<�GY<�Y<}�Z<�0\<��]<��^<K#_<X�^<g|]<P�[<yWY<U�V<d�T<��R<��Q<(Q<�qQ<d�R<M{T<�V<�Y<I`[<�  �  b�]<�1_<V`<�'`<#�_<��^<^A]<�\<I	[<�kZ<~ Z<Z<�Z<p#Z<�&Z<�!Z<�Z<Z<&-Z<k�Z<<[<�H\<��]<3�^<k�_<28`<��_<M�^<��]<��[<��Y<h)X<�V<�cU<U�T<��T<��T<�V<9uW<�%Y<V�Z<��\<}k^<�_<R>`<�'`<fm_<3B^<'�\<��[<U�Z<�mZ<:Z<V5Z<�BZ<NNZ<$PZ<�HZ<�=Z<BZ<�qZ<�Z<(�[<��\<�5^<�k_<&8`<�d`<;�_< �^<�"]<�U[<i�Y<I�W<]VV<�AU<��T<��T<rU<�V<D#X<��Y<$�[<�z]<I�^<5`<�a`<�`<!'_<'�]<��\<߄[<��Z< fZ<�DZ<`HZ<VZ<�\Z<[Z<POZ<�DZ<�RZ<�Z<�([<\<�P]<��^<�_<aU`<6F`<چ_<4^<?�\<T�Z<B�X<�BW<��U<��T<4�T<��T<&�U<W<u�X<J}Z<CR\<�^<bf_<�7`<�Z`<��_<��^<�s]<G4\<�;[<��Z<�SZ<�AZ<�JZ<�VZ<�YZ<TZ<jFZ<m@Z<\Z<ҶZ<�g[<�r\<b�]<�_<��_<g]`<c`<d_<�]<��[<�Z<�MX<]�V<L�U<��T<g�T<�#U<E+V<ݗW<9GY<�[<��\<Z�^<��_<W`<>`<{�_<�S^<  ]<��[<��Z<TtZ<>Z<u6Z<#AZ<�IZ<�HZ<{>Z<�0Z<2Z<_Z<��Z<�[<B�\<�^<7L_<U`<�@`<U�_<Q�^<��\<�*[<�UY<��W<!)V<�U<�T<B�T<�DU<qV<��W<�Y<x�[<�O]<��^<��_<6`<?�_<��^<��]<Mi\<�S[<<�Z<^2Z<�Z<�Z<�Z<�%Z<�#Z<�Z<�Z<�Z<�^Z<e�Z<�[<�]<�k^<�_<`<Z`<LO_<��]<M\<ExZ<q�X<W<�U<��T<ShT<g�T<P�U<��V<�zX<�EZ<�\<�  �  :p]<��^<}�_<�}`<{y`<��_<��^<�]]<w�[<��Z<@�Y<	�X<�X<̩W<�W<��W<�8X<��X<�Y<?�Z<�K\<Ʊ]<._<`<�`<q`<$�_<�^<�,]<�[<�Z<�Y<�X<X<�W<�W<N�W<�cX<w%Y<�Z<�D[<W�\<��]<�L_<LA`<��`<Hp`<O�_<�h^<B]<��[<�xZ<�vY<��X<:X<˽W<��W<�	X<3�X<�gY<�fZ<p�[<��\<�X^<��_<�{`<��`<�t`<.�_<�K^<h�\<��[<AcZ<\hY<�X<X<�W<q�W<W*X<D�X<̕Y<��Z<I�[<�,]<&�^<��_<w�`<\�`<rN`<7U_<�^<c�\<tQ[<(-Z<�;Y<�~X<#�W<N�W<�W<�=X<p�X<��Y<��Z<�
\<�j]<g�^<i�_<c�`<R�`<1`<�%_< �]<�j\<![<�Z<�Y<�gX<��W<��W<�W<�VX<jY<��Y<�Z<|C\<�]<b _<7`<ʰ`<�`<�	`<��^<�]<�-\<�Z<�Y<�X<�IX<��W<v�W<]�W<�iX<� Y<WZ<�*[<�v\<e�]<W/_<�4`<ѵ`<�`<h�_<Ѱ^<ZP]<��[<�Z<H�Y<��X<�2X<��W<��W<� X<��X<rHY<r=Z<e[<G�\<�^<h_<GZ`<��`<��`<�_<�w^<�]<:�[<�Z<�zY<��X<�X<2�W<4�W<g�W<�X<�WY<TZ<�[<��\<�=^<]~_<�[`<��`<�P`<j_<�#^<�\<�e[<47Z<l;Y<�sX<+�W<�W<��W<��W<�X<!iY<�nZ<��[<t]<�c^<��_<�``<6�`<|!`<<'_<��]<�p\<�[<$�Y<Y<gIX<.�W<ʉW<3�W<�X<��X<��Y<��Z<��[<�4]<��^<��_<@m`<��`<��_<��^<H�]<71\<^�Z<y�Y<��X< +X<ӲW<+�W<�W<!X<��X<P�Y<��Z<w\<�  �  �\< S]<P�^<��_<�*`<��_<�"_<��]<\<�-Z<eX<��V<t�U<k�T<�mT<��T<��U<w"W<n�X<�Z<�m\<-^<^f_<�`<�#`<�_<_d^<X]<<�[< �Z<fZ<='Z<�Z<o'Z<�3Z<�5Z<q/Z<,#Z<�"Z<mHZ<g�Z<�t[<-�\<��]<^_<Z`<\L`<��_<@�^<ZP]<͉[<K�Y<�W<>yV<�SU<�T<��T<�>U<�ZV<F�W<}�Y<f[<T3]<��^<P�_<Ne`<1`<4__<�'^<��\<߶[<��Z<�yZ<�NZ<MZ<aYZ<�`Z<D_Z<�SZ<�FZ<|MZ<��Z<I[<��[<k]<,h^<ҏ_<�B`<TQ`<!�_<�p^<�\< �Z<h,Y<��W<�V<}U<��T<�T<��U<��V<;jX<!/Z<k\<s�]<�5_<C"`<�c`<��_<K�^<�]<~i\<	c[<ݶZ<'`Z<�FZ<�MZ<�ZZ<o_Z<�[Z<�NZ<�EZ<�YZ<<�Z<J[<�F\<�]<:�^<��_<k]`<�/`<�T_<h�]<6\<`Z<p�X<j�V<�U<��T<\�T<�U<��U<ZQW<��X<,�Z<�\<7B^<��_<D`<RI`<��_<b�^<7]<� \<�[<5�Z<�KZ<�@Z<vLZ<�XZ<�ZZ<-TZ<UGZ<�EZ<�jZ<?�Z<�[<��\<�]<�8_<8`<�``<��_<u�^<�\]<��[<3�Y<-�W<nzV<�QU<m�T<�T</4U<�MV<<�W<�|Y<oP[<]<�^<��_<vE`<�`<�:_<J^<��\<�[<��Z<oMZ<p!Z<:Z<'+Z<�2Z<1Z<�%Z<[Z<� Z<JXZ<��Z<��[<Z�\<=^<�d_</`<�$`<��_<"B^</�\<��Z<�X<MW<��U<%�T<�oT<��T<�cU<�V<�3X<��Y<x�[<��]<��^<J�_<A-`<ھ_<��^<�w]<)0\<�([<�{Z<	$Z<
Z<XZ<jZ<*"Z<�Z<|Z<�
Z<�Z<xoZ<�[<�  �  ��Y<��Z<Sq\<v�]<��^<a#_<��^<�9]<�C[<K�X<��V<�aT<P�R<�jQ<�Q<"�Q<k�R<'�T<W<�Y<^�[<z�]<#�^<�+_<G�^<d�]<�%\<��Z<	�Y<�QY<�xY<�Z<}�Z<9�[<{\<4\<��[<�6[<�iZ<��Y<+[Y<I�Y<�HZ<9�[<j
]<�\^<;&_<�)_<�T^<�\<ͦZ<'MX<��U<N�S<�CR<�\Q<�QQ<6$R<ıS<g�U<�X<NvZ<�\<�F^<�5_<�L_<��^<�T]<��[<��Z<}�Y<"�Y<S�Y<;~Z<L[<1�[<_[\<N\<��[<�[<7LZ<ȭY<�wY<j�Y<��Z<�"\<��]<��^<FR_<D_<��]<�(\<��Y<ȐW<�GU<SS<.�Q<eKQ<ۊQ<7�R<�]T<ΈV<k�X<�9[<�<]<�^<�R_<�!_<%5^<�\<FZ[<?0Z<��Y<&�Y<��Y<��Z<މ[<�$\<�b\<�0\<�[<��Z<kZ<��Y<��Y<?Z<2[<g�\<�^<\_<]U_<T�^<8k]<Cu[<(Y<��V<��T<,�R<7�Q<�CQ<�Q<�S<aU<�IW<-�Y<R�[<��]<E�^<rQ_<>�^<��]<iI\<J�Z<��Y<�uY<�Y<2Z<r�Z<z�[<�?\<hY\< \<3[[<��Z<��Y<P|Y<ͤY<<fZ<ק[<�#]<�s^<�:_<�;_<)d^<��\<��Z<TX<��U<��S<�AR<KXQ<9JQ<�R<��S<S�U<�X<�`Z<��\<�+^<_<�,_<Ww^<F0]<Q�[<dZ<p�Y<�UY<��Y<�PZ<�[<��[<�,\<�\<v�[<]�Z<EZ<x�Y<'LY<+�Y<ܘZ<�[<�p]<�^<&_<-�^<��]<b�[<��Y<�^W<�U< S<h�Q<Q<UQ<7jR<v'T<�RV<��X<+[<]<Hv^<�_<^�^<�]<9�\<~![<t�Y<�UY<OMY<��Y<.�Z<�K[<��[<�$\<,�[<+a[<;�Z<��Y<UVY<'OY<�  �  ZCW<L<X<�Y<܌[<A�\<�]<^p]<q.\<EZ<KjW<��T<��Q<�O<9=N<��M<�yN<�P<zqR<54U<zX<�Z<�\<R�]<m�]<��\<4[<�uY< X<L4W<F>W<�X<�lY<<[<�u\<.f]<ڕ]<��\<4�[<�%Z<E�X<��W<~(W<��W<�X<2~Z<<1\<�l]<0�]<�?]<��[<�\Y<ΚV<��S<6Q<�<O<E#N<WN<�O<��P<�S<WV<n"Y<Q�[<;5]<{�]<�]<�z\<P�Z<�Y<��W<sQW<w�W<��X<$#Z<��[< ]<��]<y�]<`�\<t[[<��Y<PYX<�tW<�RW<EX<�mY<�*[<��\<"�]<s�]<��\<�
[<�X<A�U<0�R<��P<��N<�
N<JXN<��O<J�Q<AuT<�NW<� Z<�0\<��]<o�]<FO]<��[<;6Z<0�X<��W<iOW<��W<�Y<B�Z<u0\<$T]<O�]<�j]<�V\<�Z<�AY<��W<CTW<zW<�qX<>Z<�[<�-]<��]<��]<�_\<�CZ<��W<8�T<fR<E�O<JnN<�N<��N<ZHP<#�R<�`U<c6X<w�Z<�\<	�]<��]<]�\<X[<?�Y<|#X<�WW<bW<,3X<g�Y<X)[<��\<͋]<p�]<0]<��[<sIZ<�X<�W<@HW<��W<��X<ǗZ<pH\<��]<I�]<O]<g�[<bfY<ҡV< �S<V7Q<0;O<�N<�N<GO<J�P<drS<DV<�Y<�p[<,]<��]<�]<X\<��Z<&�X<�W<.'W<�uW<�{X<V�Y<'�[<;�\<"�]<�r]<�\<�-[<��Y<�,X<$IW<|'W<l�W<�BY<��Z<��\<F�]<��]<ܶ\<��Z<�WX<�U<��R<SP<?�N<�M<�"N< uO<��Q<�?T<W<"�Y< �[<�W]<R�]<�]<G�[<�Y<aX<pSW<W<F�W<Q�X<HjZ<�[<�]<҉]<�,]<�\<ȘZ<�Y<=�W<W<�  �  ��T<0�U<]WW<\ZY<z"[<21\<[3\<�[<�X<��U<B�R<&�O<X-M<��K<�K<L�K<�M<J[P<�}S<��V<�rY<�k[<MQ\<�\<�Z<��X<y�V<�oU<o�T<3U<��V<5�X<]�Z<��\<L/^<jp^<ǔ]<��[<T�Y<UmW<��U<�T<NU<�@V<X<�Z<:�[<=p\<�\<^�Z<KX<HU<M�Q<��N<-�L<ChK<XK<�}L<��N<�Q<��T<��W<�fZ<@
\<��\<��[<�nZ<�uX<-�V<�NU<qU<��U<7_W<��Y<�[<��]<Б^<�p^<�<]<+E[<��X<�V<>wU<��T<�xU<I�V<��X<��Z<� \<��\<�[<:�Y<�.W<	T<�P< "N<�+L<YJK<��K<[&M<�O<ߞR<��U<C�X<F[<�U\<�t\<�[<��Y<��W<
V<�U<�U<H0V<!	X<(GZ<�o\<�^<<�^<�%^<~�\<��Z<�DX<�ZV<0U<�U<��U<��W<��Y<�T[<c\<�d\<?[<=Y<�)V<y�R<Q�O<Y^M<��K<AK<� L<K�M<��P<թS<'�V<��Y<��[<�w\<A5\<��Z<_Y<�W<
�U<��T<�VU<<�V<��X<� [<�]<U^<2�^<J�]<��[<u�Y<V�W<3�U<�U<]1U<�\V<�4X<�2Z<�[<m�\<l \<�Z<4#X<VU<y�Q<��N<��L<�cK<�PK<esL<I�N<�{Q<��T<��W<"NZ<!�[<�o\<]�[<hLZ<�PX<QkV<�%U< �T<��U<!2W<�YY<o�[<�i]<�b^<�A^<M]<S[<��X<��V<}KU<��T<�MU<��V<#�X<��Z<I�[<$V\<��[<��Y<&�V<�S<��P<��M<��K<�K<�mK<�L<�bO<diR<��U<ēX<��Z< \<v>\<`J[<D�Y<��W<��U<\�T<�T<��U<x�W<�Z<�0\<��]<Pg^<_�]<�g\<[JZ<o	X<� V<��T<�  �  �S<!�S<��U<�W<3�Y<�[<�H[<�8Z<"X<��T<��Q<h>N<��K<A�I<�8I<J<qL<�N<�SR<�U<��X<b�Z<k^[<��Z<PqY<�WW<y3U<^�S<�S<W�S<�jU<;�W<w�Z<K]<��^<��^<W�]<m�[<+!Y<zV<aT<\@S<�KS<NwT<�nV<w�X<4vZ<�i[<|0[<F�Y<�4W<
�S<͍P<dM<��J<f�I<ށI<@�J<�M<�8P<&�S<a�V<%�Y<�,[<p�[<0�Z<m�X<H�V<��T<-�S<ZS<�\T<�_V<e�X<}�[<.�]<B_<B�^<p]<%[<�[X<�U<� T<�>S<��S<�$U<|@W<xcY<�Z<��[<��Z<�Y<�>V<=�R<pO<�L<�eJ<ErI<��I<�tK<~N<-`Q<o�T<��W<�;Z<�n[<4c[<�6Z<�BX<�V<�=T<�OS<8�S<��T<�/W<��Y<J|\<�^^<�_<@�^<��\<�2Z<[xW< U<��S<�DS<�T<�U<\X<�Z<�K[<z[<jZ<65X<�*U<��Q<\oN<��K<��I<�hI<27J<�9L<�O<mR<N�U<��X<ԻZ<��[<�[<��Y<:{W<�VU<��S<k7S<'�S<F�U<	X<��Z<�0]<߻^<�_<�^<��[<nEY<@�V<̂T<l`S<�iS<a�T<��V<ݹX<�Z<|[<@[<	�Y<�>W<T<��P<UeM<+�J<׎I<dzI<ݴJ<�M<~(P<-�S<��V<�yY<|[<�n[<�Z<��X<l�V<��T<S\S<�/S<�0T<s2V<E�X<��[<�]<�^<R�^<�A]<:�Z<[.X<��U<2�S<�S<@�S<h�T<�W<�8Y<��Z<�^[<u�Z<4�X<�V<��R<�MO<-SL<�1J<�=I<؜I<�?K<8�M<�*Q<�T<G�W<SZ<9[<-[<��Y<7X<�U<iT<�S<]NS<��T<��V<�Y<!=\<G^<j�^<�D^<�~\<��Y<�<W<��T<iS<�  �  �0\<�\<�]<��^<3�_<�!`<��_<
8^<h\<�\Y<�uV<�S<pQ<7�O</�O<8P<L�Q<hIT<�W<� Z<4�\<e�^<��_<�'`<1�_<��^<��]<��\<:9\<�\<��]<�|_<Ia<F�b<��c<��c<sZc<�	b<�P`<�^<� ]<3[\<a\<r]<!>^<�`_<u`<=,`<X]_<x�]<�T[<ĈX<y�U<S<��P<+�O<��O<y�P<z�R<�^U<�BX<�[<\�]<yM_<K8`<)E`<+�_<f^<tZ]<�\<�v\<X(]<��^<SF`<7b<�fc<d<�d<I"c<y�a<S�_<0&^<�\<#c\<9�\<Ս]<��^<��_<M`<7`<��^<J	]<:}Z<h�W<��T<OR<��P<��O<�P<DnQ<2�S<WV<?Y<��[<87^<ݴ_<�R`<�`<�?_<^<�]<Wn\<ϖ\<��]<�_<��`<M�b<ӷc<�,d<��c<��b<|a<-B_<��]<$�\<�f\<�\<�]<�_<r`<�S`<��_<�h^<?\<��Y<�V<;�S<��Q<�)P<�O<�fP<�R<�uT<�GW<�*Z<��\<��^<�_<M`<��_<t�^<�]<�\<�\\<U�\<��]<��_<ma<�b<��c<�d<~c<�,b<s`<�^<�@]<:y\<?}\<�6]<JV^<kv_<�2`<P=`<�k_<c�]<^[<Q�X<J�U<S<:�P<��O<��O<v�P<��R<OU<�0X<[<r]<�3_<�`<�&`<Nx_<p\^<�5]<;j\<�N\<��\<�[^<�`<��a<�9c<�c<y�c<f�b<�va<3�_<��]<ڼ\<D8\<�}\<>c]<��^<��_<{!`<��_<��^<#�\<NZ<=nW<m�T<R<�ZP<L�O<�O<:Q<�iS<w"V<Q
Y<�[<0^<�_<`<��_<�_<d�]<E�\<�4\<{\\<�M]<��^<�`<kKb<�zc< �c<,�c<.ub<��`<N_<�s]<�n\<�  �  ��\<�#]<�,^<�R_<1`<�s`<�_<�~^<�W\<��Y<!�V<$T<+�Q<�~P<�P<�P<[XR<b�T<lvW<POZ<s�\<�^<�`<�{`<�`<w_<�]<]<��\<z�\<� ^<�_<�;a<�b<'�c<��c<#0c<��a<�R`<;�^<i`]<9�\<��\< �]<S�^<��_<\x`<�z`<?�_<t�]<%�[<��X<�V<�sS<m|Q<pcP<�UP<NUQ<�9S<��U<I�X<�d[<��]<��_<��`<ʜ`<\�_<��^<6�]<��\<.�\<'k]<#�^<QK`<��a<>c<m�c<6�c<�b<F�a<�_<�P^<k1]<��\<�]<��]<�$_<�$`<\�`<1^`<�=_<3Q]<�Z<��W<,U<��R<*Q<3KP<��P<��Q<�
T<G�V<�Y<�D\<�}^<��_<o�`<dv`<U�_<m�^<�s]<��\<&�\<q�]<H+_<+�`<Rkb<��c<E�c<(�c<��b<a<3X_<��]<��\<��\<�X]<�`^<Ʌ_<Kc`<m�`<P`<��^<x�\<E�Y<�W<bNT<"R<�P<�BP<H�P<��R<��T<��W<CyZ<(]<�_<0E`<*�`<C6`<l@_<�^<g$]<�\<�]<�$^<��_<�_a<�b<V�c<��c<�Sc<�b<�t`<,�^<�]<8�\<
�\<a�]<v�^<��_<�`<�`<ó_<\^<d�[<z�X<�	V<�tS<�zQ<�^P<NNP<KKQ<-S<-�U<%�X<,P[<F�]<{_<�i`<+~`<��_<��^<R�]<�\<�\<A]<Q^<�`<)�a<'c<]�c<)�c<%�b<�fa<��_<�$^<1]<��\<U�\<��]<��^<n�_<�v`<�1`<o_<�"]<ԛZ<a�W<��T<��R<X�P<�P<dP<��Q<v�S<��V<.\Y<\<�H^<��_<�m`<2@`<o_<�L^<o;]<C�\<�\<Q�]<j�^<��`<�.b<�Mc<z�c<�cc<�Ub<*�`<c_<K�]<��\<�  �  ��]<%R^<!\_<nn`<�.a<Ta<��`<DA_<#]<��Z<��W<+PU<�BS<W�Q<̐Q<&+R<�S<��U<wuX<�,[<�]<�_<�`<;ba<}a<�=`<R&_<,^<��]<�]<{^<��_<�a<dAb<yc<�,c<��b<ڢa<2N`< _<�^<Ф]<X�]<4�^<��_<�`<�ka<�Ra<<k`<.�^<$r\<��Y<.W<(�T<��R<n�Q<��Q<�R<�~T<��V<�Y<y9\<�^<�Y`<$[a<ތa<(a<�`<��^<^<I�]<b^<�_<�O`<��a<߾b<�Pc<=c<ևb<�Za<��_<
�^<��]<��]<�=^</_<TH`<�,a<�a<�.a<Q`<^<c�[<��X<�OV<nT<�|R<��Q<�R<�FS<�AU<��W<^xZ<\]<�@_<��`<��a<�pa<پ`<�_<O�^<��]<��]<�W^<$j_<��`<Eb<��b<!\c<c< .b<��`<3�_<o^<Q�]<��]<�^< �_<h�`<&aa<��a<��`<Br_<�S]<3�Z<z
X<��U<�rS<#R<��Q<�YR<��S<MV<נX<�V[<b�]<��_<�a<��a<-;a<�a`<�I_<{O^<��]<x�]<��^<]�_<�/a<�eb<�*c<�Pc<#�b<��a<)p`<� _<u(^<��]<z^<a�^<��_<��`<Ia<�ca<�y`<�^<\{\<C�Y<�W<4�T<(�R<��Q<]�Q<�R<�qT<�V<�xY<�$\<�}^<@`<�>a<Jna<\�`<�_<��^<w�]<�]<��]<�^<6$`<j|a<�b<�#c<c<[b<X.a<��_<i�^<��]<�]<�^<u_<`<�a<X`a<Oa<��_<��]<�u[<*�X<[V<.�S<�IR<F�Q<��Q<&S<UU<�W<�CZ<q�\<�_<H�`<Ka<�:a<�`<�z_<�j^<��]<��]<�^<x._<L�`<��a<C�b<�c<��b<��a< �`<�S_<�6^<
�]<�  �  l_<��_<��`<|�a<��b<6�b<�a<�L`<�@^<8�[<�_Y<BW<RHU<� T<��S<�QT<��U<�W<��Y<�i\<��^<'�`<�b<@�b<�zb<��a<W�`<O�_<�_<��^<_<L�_<U�`<�wa<�b<Ub<j�a<#a<)`<k\_<W�^<�^<n_<u]`<vma<1Nb<��b<�vb<�xa<��_<��]<m'[<��X<�V<m�T<�T<pT<M�T<ddV<X<4�Z<ig]<T�_<@fa<�{b<��b<�}b<�a<��`<�_<�_<H_<jq_<�8`<*a<��a<�Cb<p5b<J�a<�`<�`<�H_<��^<9!_<N�_<��`<��a<A�b<��b<0Ib<�a<�,_<��\<�aZ<�X<�V< �T<� T<�?T<�QU<�W<OY<\�[<�3^<M`<�a<��b<9�b<�>b<oNa<�@`<"d_<��^<�_<�_<x�`<�`a<	b<�Kb<�b<�va<<�`<��_<� _<��^<QP_<x"`<S.a<h%b<��b<�b<b�a<�}`<�q^<\<z�Y<�IW<�xU<�PT<a�S<��T<w�U<��W<LZ<F�\<��^<�`<I+b<��b<ٟb<��a<�`<��_<>*_<E�^<�4_<�_<D�`<��a<�&b<Bb<��a<�-a<�J`<}_<�_<�_<�_<�w`<m�a<�cb<��b<ȇb<*�a<��_<��]<�-[<X�X<�V<��T<	T<0 T<M�T<�WV<pX<�Z<�R]<�_<yLa<y_b<2�b<�\b<D�a<�w`<��_<��^<��^<�F_<`<��`<�a<�b<�b<��a<��`<��_< _<\�^<P�^<��_<�`<��a<�jb<�b<vb<$�`<Y�^<��\<(1Z<F�W<U�U<�lT<��S<NT<>U<��V<)Y<k�[<��]<�`<Ρa<wb<+�b<�b<a<|`<)+_<��^<�^<�m_<�E`<�$a<��a<Ib<��a<~;a<�_`<Q�_<B�^<x�^<�  �  ��`<>�a<�b<�vc<<�c<l�c</�b<\Ra<Ug_<~A]<�[<�2Y<ܰW<�V<7wV<d�V<~�W<ؙY<��[<:�]<=�_<�a<$c<%�c<&�c<Wc<�mb<�]a<i`<g�_<=�_<��_<��_<�C`<&�`<u�`<�h`<�`<D�_<��_<�_<�`<��`<Wb<v	c<#�c<m�c<N�c<{b<��`<v�^<W�\<��Z<5�X<0tW<�V<)�V<c[W<��X<�fZ<�y\<-�^<m�`<hb<`�c<�d<�c<�Ac<!Db<6a<kW`<��_<�_<a�_<�3`<T�`<ټ`<U�`<�v`<`<�_<M�_<7�_<z`<
ha<nxb<�ic<@�c<�c<�Vc<5b<ME`<�,^<j\<�Y<�UX<�/W<�V<#�V<�W<&6Y<�[<�7]< `_<�Ta<��b<P�c<d<��c<��b<1�a<��`<�`<�_<Ѵ_<`�_<�O`<�`<&�`<�`<Y`<)�_<9�_<��_<4
`<L�`<��a<��b<��c<ud<-�c<��b<��a<��_<�r]<�N[<�cY<��W<��V<'�V<�W<�*X<%�Y<��[<�]<�`<6�a<=6c<,�c<E�c<{{c<�b<a�a<~�`<��_<ʦ_<I�_<m`<ug`<�`<�`<�`<G7`<��_<u�_<�_<}<`<qa<@b<K!c<��c<�d<)�c<]�b<^�`<��^<ʰ\<v�Z<6�X<rrW<e�V<�V<eQW<�X<~WZ<�g\<��^<3�`<MNb<Csc<��c<��c<4c<�b<�a<�/`<l�_<��_<�_<�`<�]`<2�`<��`<�I`<��_<#�_<�~_<�_<,O`<8=a<�Mb<h>c<��c<��c<�)c<D�a<V`<��]<X�[< �Y<#X<J�V<�yV<|�V<3�W<Y<��Z<�]<+_<xa<E�b<��c<'�c<,�c<p�b<T�a<=�`<�_<�~_<�y_<�_<�`<�b`<V�`<�i`<5`<'�_<1_<{_<g�_<�  �  ��a<M�b<d�c<q�d<D�d<�ed<Roc<b<LK`<�~^<��\<�R[<�2Z<�Y<�OY<[�Y<�jZ<�[<�)]<Z�^<1�`<�_b<�c<ӏd<N�d<'�d<��c<W�b<�ta<�g`<|�_<e_<��^<ޛ^<j�^<Ґ^<̖^<��^<�^<�Y_<�`<�a<�'b<fQc<�Fd<�d<�d<�@d<.c<\�a<��_<^<�h\<y[<�Z<�Y<��Y<��Y<H�Z<�G\<��]<��_<swa<�c<s>d<�d<�d<{d<7�c<�lb<�Da<�I`<g�_<�_<H�^<��^<��^<�^<�^<��^<�+_<*�_<@u`<a|a<�b<��c<��d<��d<��d<>d<+�b<�a<jI_<;�]<�[<��Z<�Y<��Y<�Y<�MZ<Ib[<��\<р^<lL`<Ib<�c<��d<�d<��d<�2d<�.c<b</�`<��_<a__< �^<��^<
�^<��^<	�^<��^<��^<�P_<��_<<�`<+�a<�c<�d<;�d<{�d<��d<�c<�3b<�|`<>�^<�\<�[<dZ<�Y<
�Y<�Y<ʙZ<��[<OV]<�_<6�`<[�b<��c<0�d<��d<˧d<��c<�b<p�a<'�`<��_< 2_<F�^<��^<�^<+�^<��^<6�^<v_<z_<q*`<�a<�Cb< kc<P^d<��d<B�d<JQd<p-c<�a<��_<t^<Rl\<t[<�Z<`�Y<�|Y<��Y<��Z<h8\<��]<Y�_<I`a<�b<m"d<��d<��d<�Xd<�lc<mFb<9a<� `<:g_<��^<��^<g�^<�^<�^<��^<��^<��^<��_<J`<gQa< }b<��c<Hod<��d<��d<��c<݈b<��`<�_<�W]<��[<A�Z<��Y<�PY<
uY<�Z<�,[<d�\<�K^<*`<�a<�Jc<,Pd<?�d<p�d<�c<H�b<��a<�`<$�_<�$_< �^<;�^<��^<7}^<�^<��^<L�^<._<�_<��`<�  �  �4b<�c<އd<5e<be<}d<'vc<L"b<��`<�V_<M)^<�8]<��\<�)\<�\<�:\<��\<2j]<�i^<�_<;a<=vb<c�c<&�d<q#e<�e<�ad<MKc<<�a<��`<�,_<5	^<�$]<ۅ\<�.\<�\<9X\<��\<y�]<�^<y�_<qWa<��b<C d<��d<O<e<)	e<UNd<c)c<L�a<�\`<�_<o�]<�]<��\<P@\<�=\<�\<]<��]<�^<%E`<Ʊa<%c<�Id<�e<2Ze<�e<=?d<c<�a<;`</�^<��]<�]<�\<�K\<�R\<��\<V8]< ^<�1_<˂`<~�a<.Oc<pd<�$e</Qe<9�d<�	d<;�b<<_a<[�_<_�^<�]<��\<vw\<D\<�W\<�\<[W]<.@^<fg_<ۿ`<D.b<m�c<B�d<79e<�Me<��d<'�c<Ӓb<y%a<��_<��^<��]<��\<;l\<�D\<�c\<|�\<Rz]<�m^<��_<��`<�ib<M�c<C�d<�De<�@e<��d<اc<�Sb<P�`<��_< [^<�j]<h�\<Z[\<�?\<�j\<�\<��]<ʖ^<��_<�2a<f�b<F�c<��d<)Ie<�,e<��d<#oc<�b<	�`<9P_<�,^<:H]<b�\<�Q\<�B\<�z\<��\<��]<��^<#`<�ta<h�b<�d<S�d<�Qe<2e<�^d<�7c<��a<�e`<�_<�]<�]<��\<�;\<�6\<y\<h]<��]<"�^<�0`<��a<��b<�-d<s�d<�9e<T�d<�d< �b<u}a<1`<>�^<�]<q�\<�_\<\\<b&\<�u\<]]<M�]<V_<�W`<y�a<+$c<�Dd<f�d<%e<m�d<#�c<��b<s/a<u�_<d�^<	�]<Ⱦ\<�B\<\<L"\<@~\<�!]<�
^<�1_<s�`<��a<Rc<�cd<�e<we<�d<�c<�Zb<��`<��_<�S^<2X]<�\<V1\<�	\<�)\<��\<8A]<�5^<�f_<��`<�  �   b<Tc<�nd<�d<Ǒd<�c<�b<��a<��`<3�_<x_<�^<ԑ^<Ѓ^<��^<�^<K�^<��^<E2_<��_<��`<(�a<}c<�d<O�d<��d<�Od<PCc<A�a<�	`<-?^<[�\<�([<�Z<�~Y<kbY<>�Y<v�Z<��[<�]<pE_<�a<�b<j�c<��d<�d<�|d<!�c<�b<�Ya<V`<B�_<�_<��^<5�^<�^<�^<��^<��^<_<��_<WL`<�La<Gwb<�c<�d<��d<\�d<�4d<�b<gfa<d�_<�]<�>\<O�Z<Z<�Y<�Y<],Z<�.[<��\<�5^<_�_<�a<�Ec<ad<W�d<E�d<DSd<.[c<2b<6a<c`<Sr_<�_<N�^<�^<�^<O�^<|�^<��^<�<_<�_<��`<�a<G�b<S�c<�d<< e<M�d<��c<�yb<�`< _<yE]<��[<��Z<��Y<��Y<e�Y<�uZ<��[<`]<r�^<��`<Lb<X�c<�d<��d<��d<�	d<��b<��a<��`<I�_<�F_<Q�^<�^<��^<-�^<��^<A�^<��^<�__</`<��`<�b<�7c< 8d<W�d<��d<td<Jgc<��a<!-`<�b^<Ƕ\<KL[<.>Z<�Y<L�Y<��Y</�Z<\\<��]<�c_<�-a<I�b<�d<��d<G�d<x�d<��c<��b<*ea<�^`<��_<._<��^<i�^<~�^<ԣ^<��^<;�^<�_<�|_<�7`<z5a<�]b<A�c<ed<��d<"�d<vd<F�b<?a<�u_<W�]<\<	�Z<I�Y<dY<�qY<\ Z<�[<&d\<>
^<6�_<�a<�c<�5d<��d<�d<)&d<#-c<�b<��`<	�_<�?_<	�^<��^<�^<�^<l�^<s�^<��^<_<_�_<i`<�ya<�b<�c<a�d<X�d<�~d<�c<Bb<ܓ`<&�^<�]<��[<SWZ<��Y<{JY<�Y<_<Z<�a[<��\<��^<�b`<�  �  ia<��b<�c<�c<Ymc<x�b<�a<w�`<��_<z{_<}�_<L�_<�&`<�p`<}�`<kd`<`<
�_<8~_<)�_<��_<.�`<��a<��b<Ϙc<^�c<#�c<,�b<�a<5_<|�\<
�Z<�X<�W<�V<�V<�W<�HX<K�Y<�\<J.^<�E`<ab<?Lc<]�c<��c<xIc<�Ub<@Fa<~\`<Z�_<�_<��_<�`<j`<̦`<��`<w`<f `<��_< �_<|�_<tY`<>a<�Nb<�Kc<��c<�d<��c<�Xb<E�`<S�^<qe\<WZ<��X<�[W<һV<y�V<ȓW<��X<K�Z<��\<_<�a<�b<^�c<d<��c<�c<�b<a<�2`<�_<Ϭ_<��_<�=`<��`<|�`<��`<|f`<�
`<Z�_<��_<��_<��`< �a<��b<?�c<�	d<��c<n.c<B�a<'�_<��]<��[<��Y<�X<�W<k�V<~�V<�W<��Y<�o[<`�]<0�_<��a<tc<2�c<�d<��c<x�b<�a<~�`< `<ݭ_<�_<��_<xY`<�`<w�`<��`<�D`<u�_<k�_<�_<3`<8�`<q�a<.�b<!�c<�d<˼c<H�b<T5a<�<_<�]<a�Z<]Y<2�W<�V<ǮV<;W<jX<�Z<Y!\<}L^<�b`<g&b<lec<�d<��c<B\c<fb<<Ta<�g`<<�_<_�_<��_<�`<Eh`<E�`<S�`<#m`<�`<>�_<�_<�_<{B`<�$a<3b<�-c<n�c<��c<�bc<�2b<-z`<�h^<�;\<�,Z<�oX<0W<	�V<��V<�gW<5�X<˖Z<��\<��^<��`<�vb<�c<&�c< �c<:�b<^�a<��`<`<W�_<�y_<��_<�`<;\`<��`<hu`<0`<��_<*�_<�w_<̾_<:i`<�aa<=rb<�Wc<5�c<��c<��b<	�a<L�_<z�]<zr[<?zY<��W<��V<�qV<�V<#�W<fHY<D8[<�]]<��_<�  �  [d`<|�a<��b<i�b<��a<�`<��_<i_<O�^<��^<?�_<�o`<Ja<�a</b<��a<ja<�>`<ni_<��^<D�^<Y<_<�`<�.a<b<2�b<�zb<e�a<�`<��]<�{[<dY<��V<uU<"T<��S<�T<	�U<�X<�fZ<�\<�/_<t	a<]=b<�b<hyb<ֵa<�`<Ȱ_<�_<��^<�>_<k�_<E�`<έa<�(b<�0b<z�a<�a<`<�\_<y�^<}_<*�_<ݦ`<:�a<t�b<��b<ktb<�Va<"�_<�M]<��Z<[jX<�VV<P�T<�T<P)T<3U<"�V<:�X<�\[<o�]<��_<}�a<�b<��b<^[b<ywa<�h`<�~_<��^<�_<;�_<RX`<4;a<��a<~Fb<�$b<[�a<9�`<��_<;3_<J�^<%8_<��_<~a<�b<j�b<"�b<�$b<��`<��^<+x\<!�Y<��W<;�U<SyT<��S<�`T<�U<�kW<G�Y<21\<�^<͘`<(b<��b<�b<�b<a<�`<�E_<��^<g#_<�_<ۢ`<}a<�b<�Eb<T�a<VOa<gn`<�_<�
_<�^<�f_<�G`<\Va<�Bb<��b<m�b<��a<�,`<T^<��[<�(Y<�V<�:U<�3T<IT<�T<QV<�"X<ӅZ<�]<�L_<P$a<dVb<��b<T�b<��a<C�`<��_<�_<��^<!E_<��_<%�`<��a<)$b<�)b<��a<��`<�`<�J_<�^<��^<Փ_<3�`<V�a<veb<��b<�Pb<.1a<3h_<�%]<~�Z<+@X<,V<��T<P�S<��S<��T<��V<ϾX<x1[<G�]<j�_<2ta<hb<��b<�.b<�Ia<:`<O_<��^<^�^<�S_<$`<a<غa<&b<O�a<�^a<��`<8�_<�^<t�^<�_<��_<3�`<~�a<�wb<9�b<j�a<��`<h�^<@\<~�Y<~oW<�U<�?T<K�S<�'T<eZU<�3W<<Y<�[<�^^<�  �  Y_<Ӿ`<-Va<U'a<�``<�L_<�F^<�]<a�]<�E^<�h_<��`<�b<\�b<5#c<D�b<L�a<sx`<�"_<�^<�]<��]<��^<%�_<b�`<	Ja<�Pa<��`<�^<��\<�)Z<RtW<��T<�	S<j�Q<n�Q<#kR<#T<eSV<�X<�[<�^<�_<�!a<ua<�a<%`<a_<	 ^<��]<!�]<g�^<�_<\a<`�b<�1c<�<c<�b< �a</`<��^<	^<�]<� ^<~_<i `<)a<O�a<nUa<}J`<�}^<;\<nY<q�V<�mT<��R<>�Q<�Q<
S<��T<�QW<FZ<:�\<��^<i�`<na<�}a<:�`<��_<T�^<��]<��]<�2^<v2_<��`<��a<��b<�Uc<'c<�Zb<(!a<��_<k�^<��]<�]<0b^<�`_<�w`<CKa<2�a<�a<`�_<��]<�7[<�X<0�U<R�S<jPR<�Q<�4R<�S<ۥU<�3X<9�Z<�w]<X�_<`�`<�a<�Ya<Ԓ`<�~_<�x^<[�]<��]<�x^<ڛ_<��`<?9b<zc<�Uc<a�b<��a<��`<�Q_<mE^<-�]<�]<�^<�_<(�`<�oa<�ua<
�`<�_<?�\<�LZ<��W<�U<�,S<R<��Q<��R<C-T<�sV<?Y<��[<�8^<�`<�:a< �a<�"a<�7`<�_<�-^<޼]<��]<��^<�`<�\a<��b<8-c<c5c<��b<�{a<�`<��^<��]<>�]<\^<��^<�`<?�`<ona<�1a<&%`<�V^<%�[<�DY<f�V<�BT<Q�R<ƭQ<��Q<s�R<U�T<0&W<�Y<}\<��^<f`<kBa<_Qa<E�`<��_<p�^<w�]<��]<s ^<��^<%P`<9�a<Y�b<Sc<"�b<�#b<R�`<7�_<$`^<ҫ]<q�]<�,^<�+_<�B`<�a<qXa<P�`<��_<��]< [<�HX<r�U<Q�S<RR<�Q<��Q<�WS<OnU<,�W<F�Z<�B]<�  �  \�^<��_<^t`<�'`<}C_<�^<�]<r�\<��\<_�]<8_<�`<zlb<�qc<��c<�Fc<�b<s�`<��^<�|]<��\<<�\<�P]<-f^<\�_<mQ`<�t`<��_<9^<5�[<c@Y<�eV<��S<Y�Q<�gP<;+P<�P<��R<J2U<jX<r�Z<zV]<K:_<P`<ω`<�`<? _<��]<��\<�\<+]<�R^<j�_<a�a<�b<��c<|�c<�c< �a<�%`<��^<nS]<��\<h�\<��]<J�^<�`<¡`<e�`<�_<��]<EG[<FyX<�U<q&S<@NQ<�]P<�{P<2�Q<ѥS<�>V<XY<r�[<Y)^<��_<�`<��`<��_<v�^<��]<�\<��\<�]<��^<��`<m+b<Bcc<F�c<��c<��b<CMa<��_<�^<3]<��\<06]<0^<�W_<H`<2�`<A`<V�^<�\<�XZ<�W<1�T<]oR<��P<�FP<��P<8R<vT<9.W<�Z<R�\<��^<�&`<C�`<.Z`<�u_<!O^<K]<��\<{�\<\�]<�k_<}a<�b<(�c<��c<)yc<@Qb<ߺ`<
_<��]<�\<�\<z]<F�^<B�_<Kw`<��`<�_<]^<�\<�cY<�V<��S<9�Q<P�P<{MP<� Q<��R<mRU<w X<7�Z<�r]<�T_<�h`<��`<�`<�_<��]<�]<i�\<�3]<Y^<��_<:�a<A�b<U�c<>�c<�c<��a<�`<)w^<?]<ְ\<'�\<H�]<��^<�_<�`<�]`<�`_<��]<D[<1PX<#|U<��R<)#Q<]2P<6PP<�wQ<azS<5V<#�X<K�[<$�]<s�_<Si`<7\`<x�_<}�^<�i]<ް\<T�\<T\]<�^</Y`<��a<�,c<x�c<{�c<k�b<La<�f_<*�]<4�\<ߐ\<� ]<��]<�"_<�`<�s`<	`<��^<�\<7!Z<�GW<��T<�6R<�P<P<9�P< R<�>T<��V<+�Y<Wx\<�  �  �O^<��_<�!`<,�_<�^<�]<b�\<j0\<z\<܉]<$_<��`<ʌb<Рc<s�c<Gsc<};b<K�`<��^<=B]<\\<<@\<<�\<�]<&!_<��_<�$`<
{_<j�]<�[<��X<�V<TS<�.Q<U�O<�O<G~P< MR<��T<��W<�Z<�]<H�^<�`<�3`<��_<��^<k]<��\<�R\<K�\<3*^<b�_<��a<G"c<��c<�d<�Gc<j�a<`<�c^<�]<Zj\<��\<d]<,�^<R�_<�J`< 4`<�>_<Bq]<��Z</#X<'BU<O�R<��P<��O<��O<`&Q<�6S<��U<��X<s�[<w�]<��_<�E`</`<�i_<�E^<)]<�w\<�~\<-Q]<K�^<͍`<�Db<`�c<�%d<��c<��b<)Ya<��_<��]<�\<:c\<Y�\<��]<J�^<5�_<�U`<e�_<��^<y�\<�	Z<J%W<bVT<x�Q<�[P<	�O<�<P<��Q<�T<S�V<��Y<=d\<��^<�_<�T`<��_<H_<�]<��\<�b\<8�\<�]<eW_<o$a<S�b<2�c<u&d<��c<mb<ɽ`<��^<p]<��\<+k\<�
]<* ^<H_<�`<�I`<m�_<P^<v�[<GY<	*V<wS<�QQ<�P<�O<��P<�mR<��T<��W<ڥZ<+]<�_<�`<�J`<Z�_<��^<B{]<[�\<�]\<�\<\0^<��_<Ѫa<o c<�c<�d<�=c<��a<�`<�Q^<��\<�S\<�w\<wH]<io^<y�_<�(`<�`<Y_<�J]<��Z<"�W<<U<��R<��P<l�O<9�O<��P<QS<��U<��X<La[<@�]<MW_<4`<�`<q<_<�^<�\<�G\<nM\<]<v�^<�X`<b<�Wc<��c<t�c<вb<&"a<�U_<G�]<�\<�-\<��\<a�]<�^<ܳ_< `<_�_<-^<kr\<�Y<5�V<�T<��Q<�"P<T�O<BP<��Q<f�S<V<��Y<M/\<�  �  \�^<��_<^t`<�'`<}C_<�^<�]<r�\<��\<_�]<8_<�`<zlb<�qc<��c<�Fc<�b<s�`<��^<�|]<��\<<�\<�P]<-f^<\�_<mQ`<�t`<��_<9^<5�[<c@Y<�eV<��S<Y�Q<�gP<;+P<�P<��R<J2U<jX<r�Z<zV]<K:_<P`<ω`<�`<? _<��]<��\<�\<+]<�R^<j�_<a�a<�b<��c<|�c<�c< �a<�%`<��^<nS]<��\<h�\<��]<J�^<�`<¡`<e�`<�_<��]<EG[<FyX<�U<q&S<@NQ<�]P<�{P<2�Q<ѥS<�>V<XY<r�[<Y)^<��_<�`<��`<��_<v�^<��]<�\<��\<�]<��^<��`<m+b<Bcc<F�c<��c<��b<CMa<��_<�^<3]<��\<06]<0^<�W_<H`<2�`<A`<V�^<�\<�XZ<�W<1�T<]oR<��P<�FP<��P<8R<vT<9.W<�Z<R�\<��^<�&`<C�`<.Z`<�u_<!O^<K]<��\<{�\<\�]<�k_<}a<�b<(�c<��c<)yc<@Qb<ߺ`<
_<��]<�\<�\<z]<F�^<B�_<Kw`<��`<�_<]^<�\<�cY<�V<��S<9�Q<P�P<{MP<� Q<��R<mRU<w X<7�Z<�r]<�T_<�h`<��`<�`<�_<��]<�]<i�\<�3]<Y^<��_<:�a<A�b<U�c<>�c<�c<��a<�`<)w^<?]<ְ\<'�\<H�]<��^<�_<�`<�]`<�`_<��]<D[<1PX<#|U<��R<)#Q<]2P<6PP<�wQ<azS<5V<#�X<K�[<$�]<s�_<Si`<7\`<x�_<}�^<�i]<ް\<T�\<T\]<�^</Y`<��a<�,c<x�c<{�c<k�b<La<�f_<*�]<4�\<ߐ\<� ]<��]<�"_<�`<�s`<	`<��^<�\<7!Z<�GW<��T<�6R<�P<P<9�P< R<�>T<��V<+�Y<Wx\<�  �  Y_<Ӿ`<-Va<U'a<�``<�L_<�F^<�]<a�]<�E^<�h_<��`<�b<\�b<5#c<D�b<L�a<sx`<�"_<�^<�]<��]<��^<%�_<b�`<	Ja<�Pa<��`<�^<��\<�)Z<RtW<��T<�	S<j�Q<n�Q<#kR<#T<eSV<�X<�[<�^<�_<�!a<ua<�a<%`<a_<	 ^<��]<!�]<g�^<�_<\a<`�b<�1c<�<c<�b< �a</`<��^<	^<�]<� ^<~_<i `<)a<O�a<nUa<}J`<�}^<;\<nY<q�V<�mT<��R<>�Q<�Q<
S<��T<�QW<FZ<:�\<��^<i�`<na<�}a<:�`<��_<T�^<��]<��]<�2^<v2_<��`<��a<��b<�Uc<'c<�Zb<(!a<��_<k�^<��]<�]<0b^<�`_<�w`<CKa<2�a<�a<`�_<��]<�7[<�X<0�U<R�S<jPR<�Q<�4R<�S<ۥU<�3X<9�Z<�w]<X�_<`�`<�a<�Ya<Ԓ`<�~_<�x^<[�]<��]<�x^<ڛ_<��`<?9b<zc<�Uc<a�b<��a<��`<�Q_<mE^<-�]<�]<�^<�_<(�`<�oa<�ua<
�`<�_<?�\<�LZ<��W<�U<�,S<R<��Q<��R<C-T<�sV<?Y<��[<�8^<�`<�:a< �a<�"a<�7`<�_<�-^<޼]<��]<��^<�`<�\a<��b<8-c<c5c<��b<�{a<�`<��^<��]<>�]<\^<��^<�`<?�`<ona<�1a<&%`<�V^<%�[<�DY<f�V<�BT<Q�R<ƭQ<��Q<s�R<U�T<0&W<�Y<}\<��^<f`<kBa<_Qa<E�`<��_<p�^<w�]<��]<s ^<��^<%P`<9�a<Y�b<Sc<"�b<�#b<R�`<7�_<$`^<ҫ]<q�]<�,^<�+_<�B`<�a<qXa<P�`<��_<��]< [<�HX<r�U<Q�S<RR<�Q<��Q<�WS<OnU<,�W<F�Z<�B]<�  �  [d`<|�a<��b<i�b<��a<�`<��_<i_<O�^<��^<?�_<�o`<Ja<�a</b<��a<ja<�>`<ni_<��^<D�^<Y<_<�`<�.a<b<2�b<�zb<e�a<�`<��]<�{[<dY<��V<uU<"T<��S<�T<	�U<�X<�fZ<�\<�/_<t	a<]=b<�b<hyb<ֵa<�`<Ȱ_<�_<��^<�>_<k�_<E�`<έa<�(b<�0b<z�a<�a<`<�\_<y�^<}_<*�_<ݦ`<:�a<t�b<��b<ktb<�Va<"�_<�M]<��Z<[jX<�VV<P�T<�T<P)T<3U<"�V<:�X<�\[<o�]<��_<}�a<�b<��b<^[b<ywa<�h`<�~_<��^<�_<;�_<RX`<4;a<��a<~Fb<�$b<[�a<9�`<��_<;3_<J�^<%8_<��_<~a<�b<j�b<"�b<�$b<��`<��^<+x\<!�Y<��W<;�U<SyT<��S<�`T<�U<�kW<G�Y<21\<�^<͘`<(b<��b<�b<�b<a<�`<�E_<��^<g#_<�_<ۢ`<}a<�b<�Eb<T�a<VOa<gn`<�_<�
_<�^<�f_<�G`<\Va<�Bb<��b<m�b<��a<�,`<T^<��[<�(Y<�V<�:U<�3T<IT<�T<QV<�"X<ӅZ<�]<�L_<P$a<dVb<��b<T�b<��a<C�`<��_<�_<��^<!E_<��_<%�`<��a<)$b<�)b<��a<��`<�`<�J_<�^<��^<Փ_<3�`<V�a<veb<��b<�Pb<.1a<3h_<�%]<~�Z<+@X<,V<��T<P�S<��S<��T<��V<ϾX<x1[<G�]<j�_<2ta<hb<��b<�.b<�Ia<:`<O_<��^<^�^<�S_<$`<a<غa<&b<O�a<�^a<��`<8�_<�^<t�^<�_<��_<3�`<~�a<�wb<9�b<j�a<��`<h�^<@\<~�Y<~oW<�U<�?T<K�S<�'T<eZU<�3W<<Y<�[<�^^<�  �  ia<��b<�c<�c<Ymc<x�b<�a<w�`<��_<z{_<}�_<L�_<�&`<�p`<}�`<kd`<`<
�_<8~_<)�_<��_<.�`<��a<��b<Ϙc<^�c<#�c<,�b<�a<5_<|�\<
�Z<�X<�W<�V<�V<�W<�HX<K�Y<�\<J.^<�E`<ab<?Lc<]�c<��c<xIc<�Ub<@Fa<~\`<Z�_<�_<��_<�`<j`<̦`<��`<w`<f `<��_< �_<|�_<tY`<>a<�Nb<�Kc<��c<�d<��c<�Xb<E�`<S�^<qe\<WZ<��X<�[W<һV<y�V<ȓW<��X<K�Z<��\<_<�a<�b<^�c<d<��c<�c<�b<a<�2`<�_<Ϭ_<��_<�=`<��`<|�`<��`<|f`<�
`<Z�_<��_<��_<��`< �a<��b<?�c<�	d<��c<n.c<B�a<'�_<��]<��[<��Y<�X<�W<k�V<~�V<�W<��Y<�o[<`�]<0�_<��a<tc<2�c<�d<��c<x�b<�a<~�`< `<ݭ_<�_<��_<xY`<�`<w�`<��`<�D`<u�_<k�_<�_<3`<8�`<q�a<.�b<!�c<�d<˼c<H�b<T5a<�<_<�]<a�Z<]Y<2�W<�V<ǮV<;W<jX<�Z<Y!\<}L^<�b`<g&b<lec<�d<��c<B\c<fb<<Ta<�g`<<�_<_�_<��_<�`<Eh`<E�`<S�`<#m`<�`<>�_<�_<�_<{B`<�$a<3b<�-c<n�c<��c<�bc<�2b<-z`<�h^<�;\<�,Z<�oX<0W<	�V<��V<�gW<5�X<˖Z<��\<��^<��`<�vb<�c<&�c< �c<:�b<^�a<��`<`<W�_<�y_<��_<�`<;\`<��`<hu`<0`<��_<*�_<�w_<̾_<:i`<�aa<=rb<�Wc<5�c<��c<��b<	�a<L�_<z�]<zr[<?zY<��W<��V<�qV<�V<#�W<fHY<D8[<�]]<��_<�  �   b<Tc<�nd<�d<Ǒd<�c<�b<��a<��`<3�_<x_<�^<ԑ^<Ѓ^<��^<�^<K�^<��^<E2_<��_<��`<(�a<}c<�d<O�d<��d<�Od<PCc<A�a<�	`<-?^<[�\<�([<�Z<�~Y<kbY<>�Y<v�Z<��[<�]<pE_<�a<�b<j�c<��d<�d<�|d<!�c<�b<�Ya<V`<B�_<�_<��^<5�^<�^<�^<��^<��^<_<��_<WL`<�La<Gwb<�c<�d<��d<\�d<�4d<�b<gfa<d�_<�]<�>\<O�Z<Z<�Y<�Y<],Z<�.[<��\<�5^<_�_<�a<�Ec<ad<W�d<E�d<DSd<.[c<2b<6a<c`<Sr_<�_<N�^<�^<�^<O�^<|�^<��^<�<_<�_<��`<�a<G�b<S�c<�d<< e<M�d<��c<�yb<�`< _<yE]<��[<��Z<��Y<��Y<e�Y<�uZ<��[<`]<r�^<��`<Lb<X�c<�d<��d<��d<�	d<��b<��a<��`<I�_<�F_<Q�^<�^<��^<-�^<��^<A�^<��^<�__</`<��`<�b<�7c< 8d<W�d<��d<td<Jgc<��a<!-`<�b^<Ƕ\<KL[<.>Z<�Y<L�Y<��Y</�Z<\\<��]<�c_<�-a<I�b<�d<��d<G�d<x�d<��c<��b<*ea<�^`<��_<._<��^<i�^<~�^<ԣ^<��^<;�^<�_<�|_<�7`<z5a<�]b<A�c<ed<��d<"�d<vd<F�b<?a<�u_<W�]<\<	�Z<I�Y<dY<�qY<\ Z<�[<&d\<>
^<6�_<�a<�c<�5d<��d<�d<)&d<#-c<�b<��`<	�_<�?_<	�^<��^<�^<�^<l�^<s�^<��^<_<_�_<i`<�ya<�b<�c<a�d<X�d<�~d<�c<Bb<ܓ`<&�^<�]<��[<SWZ<��Y<{JY<�Y<_<Z<�a[<��\<��^<�b`<�  �  �4b<�c<އd<5e<be<}d<'vc<L"b<��`<�V_<M)^<�8]<��\<�)\<�\<�:\<��\<2j]<�i^<�_<;a<=vb<c�c<&�d<q#e<�e<�ad<MKc<<�a<��`<�,_<5	^<�$]<ۅ\<�.\<�\<9X\<��\<y�]<�^<y�_<qWa<��b<C d<��d<O<e<)	e<UNd<c)c<L�a<�\`<�_<o�]<�]<��\<P@\<�=\<�\<]<��]<�^<%E`<Ʊa<%c<�Id<�e<2Ze<�e<=?d<c<�a<;`</�^<��]<�]<�\<�K\<�R\<��\<V8]< ^<�1_<˂`<~�a<.Oc<pd<�$e</Qe<9�d<�	d<;�b<<_a<[�_<_�^<�]<��\<vw\<D\<�W\<�\<[W]<.@^<fg_<ۿ`<D.b<m�c<B�d<79e<�Me<��d<'�c<Ӓb<y%a<��_<��^<��]<��\<;l\<�D\<�c\<|�\<Rz]<�m^<��_<��`<�ib<M�c<C�d<�De<�@e<��d<اc<�Sb<P�`<��_< [^<�j]<h�\<Z[\<�?\<�j\<�\<��]<ʖ^<��_<�2a<f�b<F�c<��d<)Ie<�,e<��d<#oc<�b<	�`<9P_<�,^<:H]<b�\<�Q\<�B\<�z\<��\<��]<��^<#`<�ta<h�b<�d<S�d<�Qe<2e<�^d<�7c<��a<�e`<�_<�]<�]<��\<�;\<�6\<y\<h]<��]<"�^<�0`<��a<��b<�-d<s�d<�9e<T�d<�d< �b<u}a<1`<>�^<�]<q�\<�_\<\\<b&\<�u\<]]<M�]<V_<�W`<y�a<+$c<�Dd<f�d<%e<m�d<#�c<��b<s/a<u�_<d�^<	�]<Ⱦ\<�B\<\<L"\<@~\<�!]<�
^<�1_<s�`<��a<Rc<�cd<�e<we<�d<�c<�Zb<��`<��_<�S^<2X]<�\<V1\<�	\<�)\<��\<8A]<�5^<�f_<��`<�  �  ��a<M�b<d�c<q�d<D�d<�ed<Roc<b<LK`<�~^<��\<�R[<�2Z<�Y<�OY<[�Y<�jZ<�[<�)]<Z�^<1�`<�_b<�c<ӏd<N�d<'�d<��c<W�b<�ta<�g`<|�_<e_<��^<ޛ^<j�^<Ґ^<̖^<��^<�^<�Y_<�`<�a<�'b<fQc<�Fd<�d<�d<�@d<.c<\�a<��_<^<�h\<y[<�Z<�Y<��Y<��Y<H�Z<�G\<��]<��_<swa<�c<s>d<�d<�d<{d<7�c<�lb<�Da<�I`<g�_<�_<H�^<��^<��^<�^<�^<��^<�+_<*�_<@u`<a|a<�b<��c<��d<��d<��d<>d<+�b<�a<jI_<;�]<�[<��Z<�Y<��Y<�Y<�MZ<Ib[<��\<р^<lL`<Ib<�c<��d<�d<��d<�2d<�.c<b</�`<��_<a__< �^<��^<
�^<��^<	�^<��^<��^<�P_<��_<<�`<+�a<�c<�d<;�d<{�d<��d<�c<�3b<�|`<>�^<�\<�[<dZ<�Y<
�Y<�Y<ʙZ<��[<OV]<�_<6�`<[�b<��c<0�d<��d<˧d<��c<�b<p�a<'�`<��_< 2_<F�^<��^<�^<+�^<��^<6�^<v_<z_<q*`<�a<�Cb< kc<P^d<��d<B�d<JQd<p-c<�a<��_<t^<Rl\<t[<�Z<`�Y<�|Y<��Y<��Z<h8\<��]<Y�_<I`a<�b<m"d<��d<��d<�Xd<�lc<mFb<9a<� `<:g_<��^<��^<g�^<�^<�^<��^<��^<��^<��_<J`<gQa< }b<��c<Hod<��d<��d<��c<݈b<��`<�_<�W]<��[<A�Z<��Y<�PY<
uY<�Z<�,[<d�\<�K^<*`<�a<�Jc<,Pd<?�d<p�d<�c<H�b<��a<�`<$�_<�$_< �^<;�^<��^<7}^<�^<��^<L�^<._<�_<��`<�  �  ��`<>�a<�b<�vc<<�c<l�c</�b<\Ra<Ug_<~A]<�[<�2Y<ܰW<�V<7wV<d�V<~�W<ؙY<��[<:�]<=�_<�a<$c<%�c<&�c<Wc<�mb<�]a<i`<g�_<=�_<��_<��_<�C`<&�`<u�`<�h`<�`<D�_<��_<�_<�`<��`<Wb<v	c<#�c<m�c<N�c<{b<��`<v�^<W�\<��Z<5�X<0tW<�V<)�V<c[W<��X<�fZ<�y\<-�^<m�`<hb<`�c<�d<�c<�Ac<!Db<6a<kW`<��_<�_<a�_<�3`<T�`<ټ`<U�`<�v`<`<�_<M�_<7�_<z`<
ha<nxb<�ic<@�c<�c<�Vc<5b<ME`<�,^<j\<�Y<�UX<�/W<�V<#�V<�W<&6Y<�[<�7]< `_<�Ta<��b<P�c<d<��c<��b<1�a<��`<�`<�_<Ѵ_<`�_<�O`<�`<&�`<�`<Y`<)�_<9�_<��_<4
`<L�`<��a<��b<��c<ud<-�c<��b<��a<��_<�r]<�N[<�cY<��W<��V<'�V<�W<�*X<%�Y<��[<�]<�`<6�a<=6c<,�c<E�c<{{c<�b<a�a<~�`<��_<ʦ_<I�_<m`<ug`<�`<�`<�`<G7`<��_<u�_<�_<}<`<qa<@b<K!c<��c<�d<)�c<]�b<^�`<��^<ʰ\<v�Z<6�X<rrW<e�V<�V<eQW<�X<~WZ<�g\<��^<3�`<MNb<Csc<��c<��c<4c<�b<�a<�/`<l�_<��_<�_<�`<�]`<2�`<��`<�I`<��_<#�_<�~_<�_<,O`<8=a<�Mb<h>c<��c<��c<�)c<D�a<V`<��]<X�[< �Y<#X<J�V<�yV<|�V<3�W<Y<��Z<�]<+_<xa<E�b<��c<'�c<,�c<p�b<T�a<=�`<�_<�~_<�y_<�_<�`<�b`<V�`<�i`<5`<'�_<1_<{_<g�_<�  �  l_<��_<��`<|�a<��b<6�b<�a<�L`<�@^<8�[<�_Y<BW<RHU<� T<��S<�QT<��U<�W<��Y<�i\<��^<'�`<�b<@�b<�zb<��a<W�`<O�_<�_<��^<_<L�_<U�`<�wa<�b<Ub<j�a<#a<)`<k\_<W�^<�^<n_<u]`<vma<1Nb<��b<�vb<�xa<��_<��]<m'[<��X<�V<m�T<�T<pT<M�T<ddV<X<4�Z<ig]<T�_<@fa<�{b<��b<�}b<�a<��`<�_<�_<H_<jq_<�8`<*a<��a<�Cb<p5b<J�a<�`<�`<�H_<��^<9!_<N�_<��`<��a<A�b<��b<0Ib<�a<�,_<��\<�aZ<�X<�V< �T<� T<�?T<�QU<�W<OY<\�[<�3^<M`<�a<��b<9�b<�>b<oNa<�@`<"d_<��^<�_<�_<x�`<�`a<	b<�Kb<�b<�va<<�`<��_<� _<��^<QP_<x"`<S.a<h%b<��b<�b<b�a<�}`<�q^<\<z�Y<�IW<�xU<�PT<a�S<��T<w�U<��W<LZ<F�\<��^<�`<I+b<��b<ٟb<��a<�`<��_<>*_<E�^<�4_<�_<D�`<��a<�&b<Bb<��a<�-a<�J`<}_<�_<�_<�_<�w`<m�a<�cb<��b<ȇb<*�a<��_<��]<�-[<X�X<�V<��T<	T<0 T<M�T<�WV<pX<�Z<�R]<�_<yLa<y_b<2�b<�\b<D�a<�w`<��_<��^<��^<�F_<`<��`<�a<�b<�b<��a<��`<��_< _<\�^<P�^<��_<�`<��a<�jb<�b<vb<$�`<Y�^<��\<(1Z<F�W<U�U<�lT<��S<NT<>U<��V<)Y<k�[<��]<�`<Ρa<wb<+�b<�b<a<|`<)+_<��^<�^<�m_<�E`<�$a<��a<Ib<��a<~;a<�_`<Q�_<B�^<x�^<�  �  ��]<%R^<!\_<nn`<�.a<Ta<��`<DA_<#]<��Z<��W<+PU<�BS<W�Q<̐Q<&+R<�S<��U<wuX<�,[<�]<�_<�`<;ba<}a<�=`<R&_<,^<��]<�]<{^<��_<�a<dAb<yc<�,c<��b<ڢa<2N`< _<�^<Ф]<X�]<4�^<��_<�`<�ka<�Ra<<k`<.�^<$r\<��Y<.W<(�T<��R<n�Q<��Q<�R<�~T<��V<�Y<y9\<�^<�Y`<$[a<ތa<(a<�`<��^<^<I�]<b^<�_<�O`<��a<߾b<�Pc<=c<ևb<�Za<��_<
�^<��]<��]<�=^</_<TH`<�,a<�a<�.a<Q`<^<c�[<��X<�OV<nT<�|R<��Q<�R<�FS<�AU<��W<^xZ<\]<�@_<��`<��a<�pa<پ`<�_<O�^<��]<��]<�W^<$j_<��`<Eb<��b<!\c<c< .b<��`<3�_<o^<Q�]<��]<�^< �_<h�`<&aa<��a<��`<Br_<�S]<3�Z<z
X<��U<�rS<#R<��Q<�YR<��S<MV<נX<�V[<b�]<��_<�a<��a<-;a<�a`<�I_<{O^<��]<x�]<��^<]�_<�/a<�eb<�*c<�Pc<#�b<��a<)p`<� _<u(^<��]<z^<a�^<��_<��`<Ia<�ca<�y`<�^<\{\<C�Y<�W<4�T<(�R<��Q<]�Q<�R<�qT<�V<�xY<�$\<�}^<@`<�>a<Jna<\�`<�_<��^<w�]<�]<��]<�^<6$`<j|a<�b<�#c<c<[b<X.a<��_<i�^<��]<�]<�^<u_<`<�a<X`a<Oa<��_<��]<�u[<*�X<[V<.�S<�IR<F�Q<��Q<&S<UU<�W<�CZ<q�\<�_<H�`<Ka<�:a<�`<�z_<�j^<��]<��]<�^<x._<L�`<��a<C�b<�c<��b<��a< �`<�S_<�6^<
�]<�  �  ��\<�#]<�,^<�R_<1`<�s`<�_<�~^<�W\<��Y<!�V<$T<+�Q<�~P<�P<�P<[XR<b�T<lvW<POZ<s�\<�^<�`<�{`<�`<w_<�]<]<��\<z�\<� ^<�_<�;a<�b<'�c<��c<#0c<��a<�R`<;�^<i`]<9�\<��\< �]<S�^<��_<\x`<�z`<?�_<t�]<%�[<��X<�V<�sS<m|Q<pcP<�UP<NUQ<�9S<��U<I�X<�d[<��]<��_<��`<ʜ`<\�_<��^<6�]<��\<.�\<'k]<#�^<QK`<��a<>c<m�c<6�c<�b<F�a<�_<�P^<k1]<��\<�]<��]<�$_<�$`<\�`<1^`<�=_<3Q]<�Z<��W<,U<��R<*Q<3KP<��P<��Q<�
T<G�V<�Y<�D\<�}^<��_<o�`<dv`<U�_<m�^<�s]<��\<&�\<q�]<H+_<+�`<Rkb<��c<E�c<(�c<��b<a<3X_<��]<��\<��\<�X]<�`^<Ʌ_<Kc`<m�`<P`<��^<x�\<E�Y<�W<bNT<"R<�P<�BP<H�P<��R<��T<��W<CyZ<(]<�_<0E`<*�`<C6`<l@_<�^<g$]<�\<�]<�$^<��_<�_a<�b<V�c<��c<�Sc<�b<�t`<,�^<�]<8�\<
�\<a�]<v�^<��_<�`<�`<ó_<\^<d�[<z�X<�	V<�tS<�zQ<�^P<NNP<KKQ<-S<-�U<%�X<,P[<F�]<{_<�i`<+~`<��_<��^<R�]<�\<�\<A]<Q^<�`<)�a<'c<]�c<)�c<%�b<�fa<��_<�$^<1]<��\<U�\<��]<��^<n�_<�v`<�1`<o_<�"]<ԛZ<a�W<��T<��R<X�P<�P<dP<��Q<v�S<��V<.\Y<\<�H^<��_<�m`<2@`<o_<�L^<o;]<C�\<�\<Q�]<j�^<��`<�.b<�Mc<z�c<�cc<�Ub<*�`<c_<K�]<��\<�  �  �`<�`<)Ya<��a<�b<��a<�(a<�_<<�]<��[<��Y<{yW<�U<N�T<�wT<��T<Q"V<��W<�Z<�R\<�o^<@.`<�fa<�b<�b<��a<�Ca<��`<6�`<��`<lla<db<�wc<=id<Ue<x e<Ǽd<��c<1�b<'�a<sa<*�`<��`<*a<��a<�b<~7b<��a<~�`<�__<yh]<1[<�X< W<��U<�T<:�T<�kU<��V<�X<��Z<X:]<>_<#�`<��a<�Lb<�9b<+�a<�Ea<M�`<l�`<!a<3�a<A�b<��c<w�d<�Ce<�4e<̧d<޽c<��b<��a<��`<�`<-�`<�\a<O�a<}Ab<=;b<l�a<�`<��^<Ѿ\<�~Z<=SX<?~V<q:U<��T<��T<8�U<4vW<��Y<a�[<��]<��_<�=a<Sb<LRb<�b<�a<�a<��`<
�`<�Ta<q5b<_Fc<�Id<Je<�Le<Ee<Pbd<Ddc<sQb<0ha<��`<(�`<ca<��a<#b<�Nb<�b<�Ya<�`<z*^<� \<b�Y<��W<?�U<��T<��T<�U<�NV<UX<y;Z<M|\<
�^<�U`</�a<j.b<�Bb<��a<�ga<�`<C�`<��`<a�a<�b<ݚc<�d<�$e<�Be<��d<�d<Yc</�a<(+a<Z�`<�`<�0a<;�a<7*b<�Ib<��a<�`<�j_<q]<(7[<��X<� W<��U<�T<1�T<�aU<K�V<.�X<��Z<}&]<�'_<z�`<��a<�/b<vb<��a<�"a<��`<-�`<��`<|�a<��b<9�c<��d<�e<?	e<o|d<��c<vb<��a<:�`<p�`<ý`</2a<��a<gb<�b<&~a<V`<ܤ^<�\<=OZ<�"X<�LV<U<zT<�T<ߧU<�BW<�OY<Z�[<��]<=�_<�a<<�a<�b<��a<Pga<��`<��`<-�`<Ca<W�a<�c<�d<h�d<e<��d<v(d<"+c<.b<�0a<��`<�  �  �`<�a<=�a<z#b<�bb<T-b<�ga<A`<�:^<F\<�Y<��W<�(V<�!U<��T<=MU<{V<G<X<�ZZ<w�\<U�^<Yl`<<�a<|Kb<�db<�b<��a<		a<�`<��`<mxa<�[b<n]c<�@d<U�d<��d<�d<��c<~�b<�a<�$a< �`<<�`<�[a<��a<�]b<�{b<Kb<�"a<_�_<�]<�w[< FY<�UW<��U<�U<gU<.�U<,W<�Y<?D[<f|]<}_<da<�b<��b<��b<Nb<r�a<na<�`<�:a<Y�a<��b<��c<��d<xe<�e<Q~d<��c<�b<6�a<�a<�`<)%a<��a<�-b<��b<-~b<�a<I�`<;_<]<��Z<��X<r�V<�U<�
U<�AU<v5V<\�W<�Y<�\<�3^<	`<:|a<�Rb<��b<�cb<��a<�[a<Q�`<U�`<�ga<�3b<�1c<M%d<��d<�e<��d<�<d<�Mc<Mb<�xa<�`<D�`<La<��a<
Vb<��b<�^b<��a<�?`<�j^<NE\<�
Z<Q�W<XV<kPU<�U<�zU<��V<�gX<+�Z<�\<��^<��`<��a<�pb<H�b<�6b<N�a<I,a< �`<�
a<a�a<�~b<^�c<�cd<��d<	e<̱d<��c<��b<�a<mBa<J�`<�a<hta<Gb<crb<"�b<F)b<t0a<}�_<��]<�}[<�IY<�VW<��U<�U<_U<��U<�W<(Y<�2[<�h]<�f_<��`<� b<�sb<Vbb<�a<jga<��`<��`<a<��a<�b<��c<�{d<F�d<��d<�Rd<Wvc<�tb<e�a<��`<��`<��`<=xa<�b<�]b<�Rb<Ͻa<5�`<N�^<3�\<�Z<wsX<$�V<�dU<@�T<�U<V<��W<0�Y<��[<}�]<��_<�Ga<�b<bb<�-b<�a<9$a<5�`<��`<'.a<��a<�b<��c<��d<�d<[�d<�d<kc<Eb<�Aa<��`<�  �  KQa<��a<�`b<�b<c<��b<�b<��`<��^<��\<�Z<��X<O'W<�.V<��U<5WV<yuW<!Y<�([<HQ]<]_<Za<Rb<��b<�!c<��b<�Gb<H�a<�La<�<a<i�a<q=b<�
c<3�c<�>d<`Vd<Jd<Fgc<�b<�a<aa<�Da<��a<@b<�b<�c<4c<��b<i�a<�H`<^^<�<\<� Z<GX<��V<�(V< V<��V<�X<�Y<[\<�1^<&(`<��a<`�b<�Gc<�@c<��b<�Bb<��a<�ja<}a<��a<جb<Byc<�!d<�zd<�nd<��c<�Ic<i{b<��a<Fia<
na<U�a<�^b<��b<�Fc<i3c<.�b<aja<�_<$�]<��[<f�Y<��W<��V<�V<�OV<�5W<ӶX<��Z<s�\<��^<��`<�&b<�c<�Qc<�$c<Ȧb<�b<ґa<�aa<*�a<�(b<a�b<�c<�Hd<��d<�Sd<U�c<�c<�;b<�a<�`a<t�a<��a<�b<�c<�Oc<�c<�Cb</�`<�_<]<��Z<K�X<�VW<v]V<V<҄V<C�W<�LY<mS[< {]<��_<�<a<�xb<C%c<�Fc<��b<�kb<��a<�oa<�_a<Y�a<_`b<�-c<��c<ad<�xd<�)d<?�c<�b<�a<�~a<�`a<%�a<�*b<|�b<g2c<YFc<��b<��a<�S`<�f^<�B\<($Z<�GX<��V<y$V<V<�V<`X<F�Y<�[<'^<�`<��a<w�b<�*c<�!c<��b<�b<�a<�Da<�Ua<�a<J�b<�Nc<�c<�Od<QCd<��c<�c<gPb<Ƞa<�>a<�Ca<�a<4b<��b<�c<�c<�jb<0=a<�_<4�]<�c[<�UY<J�W<dmV<�U<�V<mW<�X<�qZ<W�\<��^<5�`<��a<��b<[c<��b<(pb<j�a<�Ya<�(a<�]a<��a<�b<}{c<�d<�Fd<Ud<��c<��b<�b<�ja<q*a<�  �  �b<�b<�bc<>�c<�d<!�c<��b<��a<��_<*�]<��[<�Z<˪X<��W<��W<��W<��X<�sZ<�R\<AW^< J`<��a<�4c<l�c<]d<2�c<�Gc<G�b<6b<��a<��a<�a<cwb<��b<Gc<"Xc<�!c<@�b<�4b<#�a<'�a<��a<^b<�	c</�c<Zd<�'d<*�c<άb</a<cW_<�U]<�`[<��Y<:uX<�W<b�W<�^X<��Y<�5[<�(]<+._<�a<�b<��c<+:d<1@d<_�c<�<c<�b<mb<��a<��a<�Mb<\�b<�?c<�}c<�tc<�'c<$�b<G/b<��a<��a<kb<#�b<�\c<J�c<�Cd<�"d<�zc<�Kb<P�`<�^<z�\<��Z<�EY<�7X<��W<�W<��X<�Z<��[<��]<��_<��a<\c<�c<�Hd<'d<ԩc<@�b<�Zb<��a<��a<�b<<ub<��b<�Yc<��c<yac<�c<�b<�b<d�a<:�a<�Ib<��b<5�c<�d<rHd<~�c<�$c<3�a<Y`<n^<�\<�BZ<R�X<��W<��W<�X<�Y<��Z<�}\<5�^<�r`<�b<�[c<(d<GBd<o�c<�kc<��b<S&b<��a<��a<�b<8�b<dc<�ic<?zc<dCc<�b<�Tb<��a<��a<��a<exb<>"c<��c<�2d</:d<�c<O�b<(:a<�__<�[]<ld[<ɱY<psX<��W<Z�W<UX<��Y<('[<9]<]_<��`<n�b<��c< d<!d<K�c<�c<�lb<\�a<&�a<�a<_$b<1�b<�c<�Rc<�Ic<��b<�b<Sb<׭a<-�a<��a<��b<X2c<h�c<od<��c<Nc<3b<|`<��^<p�\<�Z<SY<YX<ΐW<��W<։X<��Y<ި[<��]<��_<ma<��b<��c<_d<*�c<Usc<�b<	#b<�a<b�a<��a<';b<��b<�c<�Gc<�'c<H�b<*Jb<�a<k�a<:�a<�  �  ��b<��c<�dd<��d<fe<��d<�c<j|b<��`<�_<4B]<��[<%�Z<6�Y<+�Y<��Y<�Z<�\<j�]<js_<�=a<��b<�d<l�d<	e<��d<hGd<��c<�b<�
b<�a<�a<
�a<��a<n�a<��a<5�a<��a<��a<R�a<8�a<mb<@0c<Cd<!�d<�e<e<��d<��c<�b<Z_`<��^<��\<�f[<_Z<��Y<��Y<UMZ<cJ[<��\<�h^<�:`< �a<]vc<U�d<S#e<�9e<$�d<�6d<�hc<|�b<�b<(�a<��a<��a<w�a<�b<b<�a<��a<)�a<��a<&#b<f�b<�c<�Zd<��d<g:e<�e<Ud<5(c<�a<�_<�^<�`\<r[<p/Z<��Y<��Y<x�Z<�[<�E]<B_<�`<��b<q�c<[�d<�7e<*%e<��d<��c<� c<Ngb<�a<I�a<2�a<��a<>
b<b<�b<�a<�a<U�a<V�a<mTb<�c<��c<ɗd<e<B9e<c�d<�c<6�b<�a<9_<�r]<��[<��Z<��Y<
�Y<0Z<B�Z<
3\<��]<��_<�fa<��b<r5d<`�d<"7e<��d<=kd<�c<-�b<�-b<��a<��a<ɻa<��a<�b<�b<��a<>�a<z�a<��a<��a<�b<pJc<�d<��d<.e<)%e<Λd<��c<�!b<�g`<|�^<��\<rg[<6]Z<R�Y<��Y<�CZ<*>[<̤\<_W^<'`<��a<�]c<�pd<Ze<�e<(�d<�d<%Dc<�}b<��a<ʔa<��a<��a<��a<��a<	�a<��a<��a<Da<ؘa<��a<��b<_fc<B0d<��d<�e<��d<C(d<��b<�la<��_<��]<w/\<}�Z<��Y<}�Y<��Y<�iZ<΋[<Y]<��^<��`<Pb<��c<^�d<Ae<_�d<�ud<��c<��b</b<I�a<�ua<o|a<ɥa<+�a<�a<��a<c�a<��a<�ta<��a<�b<�  �  �Yc<PVd<�%e<֢e<��e<�Ee<�dd<�$c<o�a<5`<�^<oh]<��\<��[<g�[<�\<��\<0�]<��^<]t`<b<:wc<¥d<�ne<z�e<��e<|e<�+d<�+c<�/b<�[a<�`<�k`<�B`<�4`<e3`<<`<�X`<��`<$a<��a<��b<o�c<h�d<&te<��e<,�e<$e<G!d<'�b<�Ca<��_<T^<6]<�q\<�\<�
\<f\<?"]<�9^<Қ_<�%a<��b<�d<�"e<��e<%�e<��e<��d<�d<�c<b<Oa<r�`<o�`<Ge`<�[`<�[`<�g`<2�`<��`<�oa<B=b<56c<�7d<,e<��e<�e<�e<w�d<��c<p\b<��`<wK_<^�]<��\<�R\<�\<)\<r�\<�}]<�^<"!`<��a<b0c<�xd<
fe<��e<��e<#me<��d<��c<��b<x�a<La<��`<�t`<�^`<�Y`<y]`<op`<��`<A	a<B�a<�b<E�c<"�d<�Xe<;�e<q�e<<we<�d<�Uc<;�a<�I`<s�^<՘]<Գ\<�.\<�	\<`C\<o�\< �]<Y_<��`<y-b<��c<��d<�e<��e<�e<u+e<,Od<�Nc<�Rb<�~a<��`<��`<e`<�V`<4U`<A]`<y`<&�`<�6a<��a<7�b<x�c<��d<m�e<�e<0�e<�3e<�.d<�b<La<�_<vW^<�6]<'p\<
\<�\<r\\<]<�*^<��_<8a<��b<�c<e<��e<3�e<�e<��d<��c<��b<��a<�&a<R�`<�Z`<�:`<�0`<�0`<�<`<Eb`<-�`<Ea<�b<�c<`d<\�d<��e<k�e<�{e<o�d<ܚc<�-b<%�`<�_<��]<��\< \<�[<-�[<Ho\<�I]<�z^<��_<){a<��b<DDd<1e<X�e<�e<�6e<�nd<Luc<�rb<��a<L�`<Jr`<�:`< %`<�`<:$`<�7`<uj`<��`<�wa<sXb<�  �  �~c<��d<Oye<��e<��e<lpe<:�d<oc<�*b<��`<�_< _<�w^<r*^<�^<07^<:�^< 0_<�`<�3a<Mwb<�c<n�d<n�e<��e<��e<�Ze<=pd<�Dc<�a<��`<S�_<��^<�s^<71^<"&^<Q^<��^<#a_<5P`<
ya<u�b<T�c<�e<��e<3f<��e<�Me<Vd<�#c<N�a<��`<��_<�^<k|^<�C^<PB^<.w^<#�^<��_<ǘ`<Z�a<Yc<
Jd<�Le<)�e<b0f<_�e<�Ce<0?d<Rc<=�a<��`<E�_<��^<��^<�O^<U^<e�^<c_<W�_<��`<�b<�Hc<Nyd<pme<jf<s)f<�e<�e<d<9�b<�a<m``<tv_<��^<�p^<�I^<�X^<��^<�%_<��_<�`<�9b<�c<5�d<
�e<�f<�&f<�e<��d<9�c<��b<Ta<�7`<�X_<f�^<:h^<XJ^<�a^<D�^<C_<�`<1a<pb<p�c<?�d<B�e<f<kf<�e<x�d<4�c<�[b<}a<�	`<�5_<
�^<�Z^<�E^<.f^<i�^<;]_<�?`<�^a<#�b<��c<��d<��e<"f<h
f<e<ߓd<�gc<"b<j�`<�_<_<U�^<ES^<�G^</r^<I�^<��_<~n`<�a<��b<4d<�#e<$�e<I(f<|�e<`]e<^cd<�.c<��a<�`<��_<��^<�z^<�?^<H;^<�m^<��^<��_<��`<��a<D�b<�1d<�1e<\�e<�f<��e<`!e<d<��b<P�a<}k`<Su_<-�^<NV^<%^<N*^<�f^<��^<��_<�`<��a<c<�Nd<�Be<�e<��e<��e<8�d<��c<�b<�Ta<i/`<�D_<��^<0=^<�^<u$^<k^<�^<A�_<c�`<.b<�Jc<xtd<%[e<]�e<�e< �e<~�d<2�c<�]b<�a<	�_<�_</�^<�.^<2^<)^<�y^<�_<��_<��`<�:b<�  �  �6c<sd<GNe<��e<Ξe<�e<:Jd<�Lc<�Lb<yoa<|�`<�i`<�9`<�'`<�$`<�*`<EB`<�|`<�`<"�a<ևb<f�c<ԃd<�He<V�e<��e<'1e<�>d<��b<�pa<��_<�t^<�H]<[t\<, \<��[<�6\<_�\<�]<OA_<��`<MVb<�c<�d<��e<��e<X�e<��d<�d<c<-b<kTa<��`<_y`<�V`<L`<�L`<eX`<Hz`<a�`<�Ma<�b<�	c<�d<r�d<��e<��e<K�e<�e<�d<d�b<a<��_<a3^<�!]<l\<�\<� \<P�\<IT]<nw^<�_<la<��b<�Ed<�Ce<V�e<_�e<�e<n�d<��c<��b<��a<
/a<`�`<xx`<�^`<�W`<Z`<fj`<\�`<g�`<d�a<�eb<Ecc<cd<e<e<�e<_�e<דe<u�d<4�c<Qb<W�`<{_<��]<��\<�B\<2\<,8\<�\<ث]<�^<�b`<��a<1kc<��d<�e<�e<��e<aNe<�{d<�}c<~b<��a<��`<֚`<�j`<TX`<�T`<Z`<�p`<Q�`<a<��a<�b<g�c<��d<Moe<!�e<��e<nUe<�bd<Rc<�a<a`<��^<Uk]<��\<"\<N\<�W\<�]<D
^<g__<��`<�qb<��c<�d<��e<��e<)�e<y
e<�#d<�c<�&b<FZa<��`<z`<�T`<�G`<�E`<�N`<n`<��`<�<a<��a<��b<0�c<��d<�e<8�e<��e<s�d<��c<�}b<[�`<�g_<�
^<W�\<B\<Z�[<,�[<�_\<�)]<�L^<r�_<�Aa<�b<d<�e<ܥe<S�e<EWe<ۚd<b�c<@�b<�a<��`<�`<qE`<+`<�#`<�%`<�5`<�a`<��`<�Ya<1b<�.c<P.d<�e<�e<�e<^e<<�d<u\c<	�a<�W`<<�^<?�]<"�\<
\<t�[<��[<"�\<ut]<r�^<�,`<r�a<�  �  �b<`�c<ڲd<ye<��d<�[d<��c<.�b<b<z�a<�va<ƅa<��a<��a<q�a<'�a<��a<��a<�}a<.�a<P?b<��b<4�c<*�d<��d<}	e<ߗd<��c<nEb<]�`<��^<�]<��[<+kZ<i�Y<֮Y<Z<1�Z<rV\<�^<�_<��a<�!c<�Id<��d<�#e<��d<v<d<�qc<C�b<�	b<��a<[�a<Q�a<7�a<�b<�b<�a<�a<2�a<)�a<~
b<�b<fnc<c=d<V�d<z;e<�e<X�d<�hc<\�a<R)`<�X^<2�\<�E[<YPZ<��Y<�Y<\zZ<�[<��\<ź^<$�`<p@b<۫c<��d<n,e<�-e<�d<�d<�?c<�b<��a<*�a<0�a<��a<!b<_b<�b<��a<�a<��a<�a<�;b<�b<��c<�{d<�e<�=e<��d<�-d<��b<Ua<9�_<a�]<P$\<�Z<�Z<a�Y<�	Z<��Z<@�[<�]<�U_<�"a<(�b<�d<��d<�:e<�e<_�d<��c<��b<wIb<��a<1�a<"�a<��a<�
b<�b<�b<��a<��a<v�a<��a<�ib<G%c<W�c<1�d<�"e<�.e<L�d<��c<�hb<k�`<{�^<i)]<�[<D�Z<*�Y<#�Y<�6Z<$[<xu\<�^<��_<�a<q;c<�ad<�e<e7e<��d<�Kd<c<�b<b<��a<��a<	�a<\�a<b<�b<y�a<޶a<��a<��a<��a<�b<Vc<�"d<��d<�e<A�d<`d<�Dc<�a<�`<A1^<�\<K[<}&Z<��Y<��Y<�OZ<|^[<�\<3�^<�``<�b<�c<r�d<� e<Te<�d<��c<c<\Pb<��a<sa<�|a<S�a<�a<��a<��a<�a<�a<�ta<'�a<�b<Q�b<:�c<Gd<��d<�e<Z�d<��c<p�b<a<�R_<|�]<�[<��Z<"�Y<�Y<��Y<F�Z<1�[<�W]< _<��`<�  �  �a<;c<9�c<�d<��c<�Zc<F�b<mb<��a<8�a<L�a<�Tb<^�b<0/c<�Kc<= c<@�b<�9b<$�a<n�a<��a<�2b<�b<��c<�c<�d<(�c<��b<gaa<#�_<=�]<֚[<*�Y<шX<��W<��W<� X<8Y<O�Z<��\<ý^<Ψ`<Fb<ioc<1d</,d<��c<z?c<��b<kb<�a< �a<_$b<��b<c<Qgc<�lc<%,c<�b<;b<�a<-�a<�	b<�b<PBc<��c<_Bd<X7d<�c<čb<^�`<�_<h]<�&[<��Y<%_X<��W<<�W<�X<��Y<��[<'�]<��_<Za<u�b<P�c<�@d<�1d<e�c<�c<�pb<r�a<��a<��a<e]b<�b<�Jc<L~c<jc<[c<��b<b<�a<?�a<�3b<��b<�{c<�
d<�Id<�d<MTc<Eb<L_`<k^<�g\<��Z<�Y<}X<��W<�	X<��X<�]Z<�/\<�0^<])`<��a<{5c<�d<�Hd<�d<,�c<��b<�?b<&�a<��a<�b<:�b<�c<d`c<�|c<_Pc<��b<+hb<n�a<��a<p�a<c\b<kc<۫c<F%d<�@d<��c<��b<ڄa<6�_<�]<]�[<r�Y<ϪX<��W<��W<AX<�WY<.�Z<��\<A�^<��`<_b<�c<�&d<�?d<0�c<�Nc<��b<"b<G�a<��a<�'b<L�b<9c<�bc<�ec<�"c<ʭb<\,b<��a<��a<��a<�{b<�'c<��c<�#d<�d<��c<�ib<)�`<�^<��\<n�Z<�\Y<m5X<��W<�W<qhX<8�Y<b[<�Y]<�Z_<c/a<��b<
�c<�d<7d<:�c<��b<�Ab<l�a<{�a<��a<�*b<p�b<Uc<�Ic<�4c<�b<Abb<��a<�a<I�a<��a<�b<�Fc<��c<�d<,�c<~c<�a<�(`<�3^<>0\<�UZ<��X<W�W<��W<��W<��X<�&Z<|�[<�]<��_<�  �  ��`<� b<��b<Rc<T�b<�Xb<��a<PNa<-a<�sa<�b<x�b<�c<�"d<�Jd<�d<�vc<D�b<��a<�^a<l0a<�fa<��a<�b<�b<T%c<��b<-�a<�|`<��^<�\<caZ<xX<��V<�#V<�U<�V<4�W<~�Y<=�[<޼]<��_<Bea<��b<!!c<�.c<��b<*Bb<�a<�Xa</Za<��a<6ub<Dc<��c<bd<6id<�d<�`c<C�b<�a<�oa<ea<�a<Gb<��b<�Cc<�Ec<�b<&�a<�`<^<�[<��Y<X<��V<�)V<�=V<�W<�nX<�NZ<m\<��^<�t`<�a<Q�b<Lc<�0c<{�b<�#b<R�a<�`a<��a<�b<6�b<�c<h3d<$}d<r`d<$�c<'c<�Zb<��a<�ca<�ya<��a<{b<bc<Oc<�&c<rb<M.a<q_<c]<�;[<Z8Y<
�W<UV<=V<4kV<HmW<�Y<��Z<V%]<�8_<Za<�Sb<}c<}Oc</c<\�b<9�a<�a<�^a<[�a<�Bb<Lc<��c<�Sd<�{d<!=d<J�c<��b<�b<J�a<�[a<��a<`b<��b<}#c<�Jc<d�b<.b<u�`<
�^<٥\<�Z<=�X<p!W<sEV<V<}�V<��W<>�Y<�[<@�]<��_<�~a<B�b<�6c<^Bc<t�b<�Qb<-�a<Vca<mba<��a<sxb<�Dc<��c<�]d</bd<Dd<�Tc<��b<��a<9\a<Oa<�a<�,b<J�b<%c<J%c<��b<v�a<��_<��]<��[<=�Y< �W<��V<��U<bV<��V<�DX<$Z<�B\<
c^<�I`<�a<��b<$ c<Hc<)�b<��a<pa<J0a<BSa<z�a<�b<�`c<��c<)Hd<*+d<��c<��b<T%b<s�a<�.a<Ea<�a<>Fb<��b<c<<�b<r<b<6�`<�:_< ,]<+[<� Y</\W<nGV<r�U<�3V<-6W<�X<�Z<�\<z_<�  �  T$`<�ua<'3b<zab<�b<͙a<*a<]�`<��`<�Ma<�%b<�%c<d<��d<��d<^�d<��c<p�b<��a<,a<!�`<��`<p3a<��a<*<b<�kb<�b<Ba<*�_<�]<e�[<��Y<g�W<:�U<RU<~�T<I�U<1�V<��X<��Z<�]<g_<C�`<U�a<kb<Rpb<�b<�a<�a<;�`<�a<�a<˜b<\�c<�wd<�d<M�d<$�d<=�c<��b<c�a<%*a<��`<�a<��a<b<p�b<��b<�b<�a<Hi_<�e]<�-[<Y<F W<,�U<�U<.U<�V<�~W<1uY<4�[<[�]<T�_<kHa<�7b<M�b<�pb<��a<sna<�a<��`<kKa<
b<�c<��c<��d<�e<��d<.]d< wc<�ub<m�a<�a<��`<9a<$�a<bDb<4�b<�rb<�a<#�`<��^<8�\<lZ<RX<x�V<htU<�U<�^U<�oV<�X<-Z<�g\<��^<X`<��a<�eb<��b<qOb<}�a<�Ca<	�`<� a<�a<�Wb<�Wc<�Cd<-�d<e<��d<_d<>c<s b<�Xa<_�`<��`<(\a<�a<�bb<�b<�Db<fa<��_</^<(�[<�Y<��W< V<�6U<|U<��U<��V</�X<C�Z<!]<H-_<��`<��a<(�b<��b<}#b<m�a<�a<��`<�a<��a<�b<
�c<�ud<��d<G�d<��d<�c<>�b<H�a<�a<��`<��`<?sa<��a<�eb<�nb<��a<R�`<:D_<S?]<M[<��X<H�V<��U<��T<�U<v�U<~TW<�JY<�~[<ů]<��_<ja<b<^gb<�Cb<�a<@a<��`<��`<a<��a<x�b<��c<��d<��d<�d<�'d<tAc<e@b<&aa<��`<ջ`<8a<f�a<�b<>]b<=b<��a<'O`<R�^<`p\<�4Z<�X<�`V<�<U<Z�T<h'U<�8V<x�W<G�Y<w2\<%U^<�  �  /�_<�6a<A�a<vb<��a<Ra<�`<�`<��`<,>a<�*b<�=c<U8d<|�d<�e<��d<d<0c<A�a<a<��`<��`<>�`<�wa<��a<n&b<��a<ua<��_<'�]<�{[<�=Y<�5W<ͣU<��T<:�T<&U<itV<6QX<@�Z<��\<�^<~`<��a<c(b<�(b<��a<nAa<H�`<ݪ`<��`<T�a<s�b<��c<�d<�(e<�1e<R�d<�c<��b<�a<�a<��`<�`<�Ha<��a<�<b<[Kb<��a<��`<2*_<H#]<��Z<��X<J�V<LiU<��T<�T<�U<�)W<�'Y<�b[<��]<��_<�	a<��a<�Nb<6(b<��a<T+a< �`<��`<I5a<Rb<�c<�d<��d<�Ge<1#e<Ԅd<��c<%}b<G�a<��`<�`<"�`<va<G�a<�Kb<g0b<Ԇa<G`<ڂ^<;c\<�!Z< X<Z?V<|U<��T<|U<V<��W<�Y<#\<\I^<�`<�ia<�#b<�Mb<ub<��a<�a<��`<h�`<pa<�\b<�oc<:jd<!e<$Ge<5�d<�6d<1c<!b<�Da<+�`<��`<a<H�a<	b<�Kb<b<�'a<<�_<A�]<��[<M`Y<XW<��U<�T<3�T<fFU<��V<�oX<ϞZ<,�\<��^<_�`<�a<>b<�<b<K�a<�Pa<L�`<��`<�`<�a<��b<-�c< �d<y$e<�*e<��d<��c<��b<��a<�`<�`<��`<[.a<\�a<Eb<+b<±a<�`<)_< �\<��Z<j�X<Q�V<�?U<��T<�T<�}U<2�V<�X<g8[<fn]<�`_<��`<J�a<�"b<��a<#�a<��`<��`<z�`<�a<��a<1�b<}�c<:�d<�e<��d<?Od<[c<�Gb<�Sa<͵`<%�`<X�`<GAa<}�a<�b<3�a<IQa<`<yL^<n,\<��Y<��W<�V<��T<rT<*�T<5�U<��W<F�Y<��[<�^<�  �  T$`<�ua<'3b<zab<�b<͙a<*a<]�`<��`<�Ma<�%b<�%c<d<��d<��d<^�d<��c<p�b<��a<,a<!�`<��`<p3a<��a<*<b<�kb<�b<Ba<*�_<�]<e�[<��Y<g�W<:�U<RU<~�T<I�U<1�V<��X<��Z<�]<g_<C�`<U�a<kb<Rpb<�b<�a<�a<;�`<�a<�a<˜b<\�c<�wd<�d<M�d<$�d<=�c<��b<c�a<%*a<��`<�a<��a<b<p�b<��b<�b<�a<Hi_<�e]<�-[<Y<F W<,�U<�U<.U<�V<�~W<1uY<4�[<[�]<T�_<kHa<�7b<M�b<�pb<��a<sna<�a<��`<kKa<
b<�c<��c<��d<�e<��d<.]d< wc<�ub<m�a<�a<��`<9a<$�a<bDb<4�b<�rb<�a<#�`<��^<8�\<lZ<RX<x�V<htU<�U<�^U<�oV<�X<-Z<�g\<��^<X`<��a<�eb<��b<qOb<}�a<�Ca<	�`<� a<�a<�Wb<�Wc<�Cd<-�d<e<��d<_d<>c<s b<�Xa<_�`<��`<(\a<�a<�bb<�b<�Db<fa<��_</^<(�[<�Y<��W< V<�6U<|U<��U<��V</�X<C�Z<!]<H-_<��`<��a<(�b<��b<}#b<m�a<�a<��`<�a<��a<�b<
�c<�ud<��d<G�d<��d<�c<>�b<H�a<�a<��`<��`<?sa<��a<�eb<�nb<��a<R�`<:D_<S?]<M[<��X<H�V<��U<��T<�U<v�U<~TW<�JY<�~[<ů]<��_<ja<b<^gb<�Cb<�a<@a<��`<��`<a<��a<x�b<��c<��d<��d<�d<�'d<tAc<e@b<&aa<��`<ջ`<8a<f�a<�b<>]b<=b<��a<'O`<R�^<`p\<�4Z<�X<�`V<�<U<Z�T<h'U<�8V<x�W<G�Y<w2\<%U^<�  �  ��`<� b<��b<Rc<T�b<�Xb<��a<PNa<-a<�sa<�b<x�b<�c<�"d<�Jd<�d<�vc<D�b<��a<�^a<l0a<�fa<��a<�b<�b<T%c<��b<-�a<�|`<��^<�\<caZ<xX<��V<�#V<�U<�V<4�W<~�Y<=�[<޼]<��_<Bea<��b<!!c<�.c<��b<*Bb<�a<�Xa</Za<��a<6ub<Dc<��c<bd<6id<�d<�`c<C�b<�a<�oa<ea<�a<Gb<��b<�Cc<�Ec<�b<&�a<�`<^<�[<��Y<X<��V<�)V<�=V<�W<�nX<�NZ<m\<��^<�t`<�a<Q�b<Lc<�0c<{�b<�#b<R�a<�`a<��a<�b<6�b<�c<h3d<$}d<r`d<$�c<'c<�Zb<��a<�ca<�ya<��a<{b<bc<Oc<�&c<rb<M.a<q_<c]<�;[<Z8Y<
�W<UV<=V<4kV<HmW<�Y<��Z<V%]<�8_<Za<�Sb<}c<}Oc</c<\�b<9�a<�a<�^a<[�a<�Bb<Lc<��c<�Sd<�{d<!=d<J�c<��b<�b<J�a<�[a<��a<`b<��b<}#c<�Jc<d�b<.b<u�`<
�^<٥\<�Z<=�X<p!W<sEV<V<}�V<��W<>�Y<�[<@�]<��_<�~a<B�b<�6c<^Bc<t�b<�Qb<-�a<Vca<mba<��a<sxb<�Dc<��c<�]d</bd<Dd<�Tc<��b<��a<9\a<Oa<�a<�,b<J�b<%c<J%c<��b<v�a<��_<��]<��[<=�Y< �W<��V<��U<bV<��V<�DX<$Z<�B\<
c^<�I`<�a<��b<$ c<Hc<)�b<��a<pa<J0a<BSa<z�a<�b<�`c<��c<)Hd<*+d<��c<��b<T%b<s�a<�.a<Ea<�a<>Fb<��b<c<<�b<r<b<6�`<�:_< ,]<+[<� Y</\W<nGV<r�U<�3V<-6W<�X<�Z<�\<z_<�  �  �a<;c<9�c<�d<��c<�Zc<F�b<mb<��a<8�a<L�a<�Tb<^�b<0/c<�Kc<= c<@�b<�9b<$�a<n�a<��a<�2b<�b<��c<�c<�d<(�c<��b<gaa<#�_<=�]<֚[<*�Y<шX<��W<��W<� X<8Y<O�Z<��\<ý^<Ψ`<Fb<ioc<1d</,d<��c<z?c<��b<kb<�a< �a<_$b<��b<c<Qgc<�lc<%,c<�b<;b<�a<-�a<�	b<�b<PBc<��c<_Bd<X7d<�c<čb<^�`<�_<h]<�&[<��Y<%_X<��W<<�W<�X<��Y<��[<'�]<��_<Za<u�b<P�c<�@d<�1d<e�c<�c<�pb<r�a<��a<��a<e]b<�b<�Jc<L~c<jc<[c<��b<b<�a<?�a<�3b<��b<�{c<�
d<�Id<�d<MTc<Eb<L_`<k^<�g\<��Z<�Y<}X<��W<�	X<��X<�]Z<�/\<�0^<])`<��a<{5c<�d<�Hd<�d<,�c<��b<�?b<&�a<��a<�b<:�b<�c<d`c<�|c<_Pc<��b<+hb<n�a<��a<p�a<c\b<kc<۫c<F%d<�@d<��c<��b<ڄa<6�_<�]<]�[<r�Y<ϪX<��W<��W<AX<�WY<.�Z<��\<A�^<��`<_b<�c<�&d<�?d<0�c<�Nc<��b<"b<G�a<��a<�'b<L�b<9c<�bc<�ec<�"c<ʭb<\,b<��a<��a<��a<�{b<�'c<��c<�#d<�d<��c<�ib<)�`<�^<��\<n�Z<�\Y<m5X<��W<�W<qhX<8�Y<b[<�Y]<�Z_<c/a<��b<
�c<�d<7d<:�c<��b<�Ab<l�a<{�a<��a<�*b<p�b<Uc<�Ic<�4c<�b<Abb<��a<�a<I�a<��a<�b<�Fc<��c<�d<,�c<~c<�a<�(`<�3^<>0\<�UZ<��X<W�W<��W<��W<��X<�&Z<|�[<�]<��_<�  �  �b<`�c<ڲd<ye<��d<�[d<��c<.�b<b<z�a<�va<ƅa<��a<��a<q�a<'�a<��a<��a<�}a<.�a<P?b<��b<4�c<*�d<��d<}	e<ߗd<��c<nEb<]�`<��^<�]<��[<+kZ<i�Y<֮Y<Z<1�Z<rV\<�^<�_<��a<�!c<�Id<��d<�#e<��d<v<d<�qc<C�b<�	b<��a<[�a<Q�a<7�a<�b<�b<�a<�a<2�a<)�a<~
b<�b<fnc<c=d<V�d<z;e<�e<X�d<�hc<\�a<R)`<�X^<2�\<�E[<YPZ<��Y<�Y<\zZ<�[<��\<ź^<$�`<p@b<۫c<��d<n,e<�-e<�d<�d<�?c<�b<��a<*�a<0�a<��a<!b<_b<�b<��a<�a<��a<�a<�;b<�b<��c<�{d<�e<�=e<��d<�-d<��b<Ua<9�_<a�]<P$\<�Z<�Z<a�Y<�	Z<��Z<@�[<�]<�U_<�"a<(�b<�d<��d<�:e<�e<_�d<��c<��b<wIb<��a<1�a<"�a<��a<�
b<�b<�b<��a<��a<v�a<��a<�ib<G%c<W�c<1�d<�"e<�.e<L�d<��c<�hb<k�`<{�^<i)]<�[<D�Z<*�Y<#�Y<�6Z<$[<xu\<�^<��_<�a<q;c<�ad<�e<e7e<��d<�Kd<c<�b<b<��a<��a<	�a<\�a<b<�b<y�a<޶a<��a<��a<��a<�b<Vc<�"d<��d<�e<A�d<`d<�Dc<�a<�`<A1^<�\<K[<}&Z<��Y<��Y<�OZ<|^[<�\<3�^<�``<�b<�c<r�d<� e<Te<�d<��c<c<\Pb<��a<sa<�|a<S�a<�a<��a<��a<�a<�a<�ta<'�a<�b<Q�b<:�c<Gd<��d<�e<Z�d<��c<p�b<a<�R_<|�]<�[<��Z<"�Y<�Y<��Y<F�Z<1�[<�W]< _<��`<�  �  �6c<sd<GNe<��e<Ξe<�e<:Jd<�Lc<�Lb<yoa<|�`<�i`<�9`<�'`<�$`<�*`<EB`<�|`<�`<"�a<ևb<f�c<ԃd<�He<V�e<��e<'1e<�>d<��b<�pa<��_<�t^<�H]<[t\<, \<��[<�6\<_�\<�]<OA_<��`<MVb<�c<�d<��e<��e<X�e<��d<�d<c<-b<kTa<��`<_y`<�V`<L`<�L`<eX`<Hz`<a�`<�Ma<�b<�	c<�d<r�d<��e<��e<K�e<�e<�d<d�b<a<��_<a3^<�!]<l\<�\<� \<P�\<IT]<nw^<�_<la<��b<�Ed<�Ce<V�e<_�e<�e<n�d<��c<��b<��a<
/a<`�`<xx`<�^`<�W`<Z`<fj`<\�`<g�`<d�a<�eb<Ecc<cd<e<e<�e<_�e<דe<u�d<4�c<Qb<W�`<{_<��]<��\<�B\<2\<,8\<�\<ث]<�^<�b`<��a<1kc<��d<�e<�e<��e<aNe<�{d<�}c<~b<��a<��`<֚`<�j`<TX`<�T`<Z`<�p`<Q�`<a<��a<�b<g�c<��d<Moe<!�e<��e<nUe<�bd<Rc<�a<a`<��^<Uk]<��\<"\<N\<�W\<�]<D
^<g__<��`<�qb<��c<�d<��e<��e<)�e<y
e<�#d<�c<�&b<FZa<��`<z`<�T`<�G`<�E`<�N`<n`<��`<�<a<��a<��b<0�c<��d<�e<8�e<��e<s�d<��c<�}b<[�`<�g_<�
^<W�\<B\<Z�[<,�[<�_\<�)]<�L^<r�_<�Aa<�b<d<�e<ܥe<S�e<EWe<ۚd<b�c<@�b<�a<��`<�`<qE`<+`<�#`<�%`<�5`<�a`<��`<�Ya<1b<�.c<P.d<�e<�e<�e<^e<<�d<u\c<	�a<�W`<<�^<?�]<"�\<
\<t�[<��[<"�\<ut]<r�^<�,`<r�a<�  �  �~c<��d<Oye<��e<��e<lpe<:�d<oc<�*b<��`<�_< _<�w^<r*^<�^<07^<:�^< 0_<�`<�3a<Mwb<�c<n�d<n�e<��e<��e<�Ze<=pd<�Dc<�a<��`<S�_<��^<�s^<71^<"&^<Q^<��^<#a_<5P`<
ya<u�b<T�c<�e<��e<3f<��e<�Me<Vd<�#c<N�a<��`<��_<�^<k|^<�C^<PB^<.w^<#�^<��_<ǘ`<Z�a<Yc<
Jd<�Le<)�e<b0f<_�e<�Ce<0?d<Rc<=�a<��`<E�_<��^<��^<�O^<U^<e�^<c_<W�_<��`<�b<�Hc<Nyd<pme<jf<s)f<�e<�e<d<9�b<�a<m``<tv_<��^<�p^<�I^<�X^<��^<�%_<��_<�`<�9b<�c<5�d<
�e<�f<�&f<�e<��d<9�c<��b<Ta<�7`<�X_<f�^<:h^<XJ^<�a^<D�^<C_<�`<1a<pb<p�c<?�d<B�e<f<kf<�e<x�d<4�c<�[b<}a<�	`<�5_<
�^<�Z^<�E^<.f^<i�^<;]_<�?`<�^a<#�b<��c<��d<��e<"f<h
f<e<ߓd<�gc<"b<j�`<�_<_<U�^<ES^<�G^</r^<I�^<��_<~n`<�a<��b<4d<�#e<$�e<I(f<|�e<`]e<^cd<�.c<��a<�`<��_<��^<�z^<�?^<H;^<�m^<��^<��_<��`<��a<D�b<�1d<�1e<\�e<�f<��e<`!e<d<��b<P�a<}k`<Su_<-�^<NV^<%^<N*^<�f^<��^<��_<�`<��a<c<�Nd<�Be<�e<��e<��e<8�d<��c<�b<�Ta<i/`<�D_<��^<0=^<�^<u$^<k^<�^<A�_<c�`<.b<�Jc<xtd<%[e<]�e<�e< �e<~�d<2�c<�]b<�a<	�_<�_</�^<�.^<2^<)^<�y^<�_<��_<��`<�:b<�  �  �Yc<PVd<�%e<֢e<��e<�Ee<�dd<�$c<o�a<5`<�^<oh]<��\<��[<g�[<�\<��\<0�]<��^<]t`<b<:wc<¥d<�ne<z�e<��e<|e<�+d<�+c<�/b<�[a<�`<�k`<�B`<�4`<e3`<<`<�X`<��`<$a<��a<��b<o�c<h�d<&te<��e<,�e<$e<G!d<'�b<�Ca<��_<T^<6]<�q\<�\<�
\<f\<?"]<�9^<Қ_<�%a<��b<�d<�"e<��e<%�e<��e<��d<�d<�c<b<Oa<r�`<o�`<Ge`<�[`<�[`<�g`<2�`<��`<�oa<B=b<56c<�7d<,e<��e<�e<�e<w�d<��c<p\b<��`<wK_<^�]<��\<�R\<�\<)\<r�\<�}]<�^<"!`<��a<b0c<�xd<
fe<��e<��e<#me<��d<��c<��b<x�a<La<��`<�t`<�^`<�Y`<y]`<op`<��`<A	a<B�a<�b<E�c<"�d<�Xe<;�e<q�e<<we<�d<�Uc<;�a<�I`<s�^<՘]<Գ\<�.\<�	\<`C\<o�\< �]<Y_<��`<y-b<��c<��d<�e<��e<�e<u+e<,Od<�Nc<�Rb<�~a<��`<��`<e`<�V`<4U`<A]`<y`<&�`<�6a<��a<7�b<x�c<��d<m�e<�e<0�e<�3e<�.d<�b<La<�_<vW^<�6]<'p\<
\<�\<r\\<]<�*^<��_<8a<��b<�c<e<��e<3�e<�e<��d<��c<��b<��a<�&a<R�`<�Z`<�:`<�0`<�0`<�<`<Eb`<-�`<Ea<�b<�c<`d<\�d<��e<k�e<�{e<o�d<ܚc<�-b<%�`<�_<��]<��\< \<�[<-�[<Ho\<�I]<�z^<��_<){a<��b<DDd<1e<X�e<�e<�6e<�nd<Luc<�rb<��a<L�`<Jr`<�:`< %`<�`<:$`<�7`<uj`<��`<�wa<sXb<�  �  ��b<��c<�dd<��d<fe<��d<�c<j|b<��`<�_<4B]<��[<%�Z<6�Y<+�Y<��Y<�Z<�\<j�]<js_<�=a<��b<�d<l�d<	e<��d<hGd<��c<�b<�
b<�a<�a<
�a<��a<n�a<��a<5�a<��a<��a<R�a<8�a<mb<@0c<Cd<!�d<�e<e<��d<��c<�b<Z_`<��^<��\<�f[<_Z<��Y<��Y<UMZ<cJ[<��\<�h^<�:`< �a<]vc<U�d<S#e<�9e<$�d<�6d<�hc<|�b<�b<(�a<��a<��a<w�a<�b<b<�a<��a<)�a<��a<&#b<f�b<�c<�Zd<��d<g:e<�e<Ud<5(c<�a<�_<�^<�`\<r[<p/Z<��Y<��Y<x�Z<�[<�E]<B_<�`<��b<q�c<[�d<�7e<*%e<��d<��c<� c<Ngb<�a<I�a<2�a<��a<>
b<b<�b<�a<�a<U�a<V�a<mTb<�c<��c<ɗd<e<B9e<c�d<�c<6�b<�a<9_<�r]<��[<��Z<��Y<
�Y<0Z<B�Z<
3\<��]<��_<�fa<��b<r5d<`�d<"7e<��d<=kd<�c<-�b<�-b<��a<��a<ɻa<��a<�b<�b<��a<>�a<z�a<��a<��a<�b<pJc<�d<��d<.e<)%e<Λd<��c<�!b<�g`<|�^<��\<rg[<6]Z<R�Y<��Y<�CZ<*>[<̤\<_W^<'`<��a<�]c<�pd<Ze<�e<(�d<�d<%Dc<�}b<��a<ʔa<��a<��a<��a<��a<	�a<��a<��a<Da<ؘa<��a<��b<_fc<B0d<��d<�e<��d<C(d<��b<�la<��_<��]<w/\<}�Z<��Y<}�Y<��Y<�iZ<΋[<Y]<��^<��`<Pb<��c<^�d<Ae<_�d<�ud<��c<��b</b<I�a<�ua<o|a<ɥa<+�a<�a<��a<c�a<��a<�ta<��a<�b<�  �  �b<�b<�bc<>�c<�d<!�c<��b<��a<��_<*�]<��[<�Z<˪X<��W<��W<��W<��X<�sZ<�R\<AW^< J`<��a<�4c<l�c<]d<2�c<�Gc<G�b<6b<��a<��a<�a<cwb<��b<Gc<"Xc<�!c<@�b<�4b<#�a<'�a<��a<^b<�	c</�c<Zd<�'d<*�c<άb</a<cW_<�U]<�`[<��Y<:uX<�W<b�W<�^X<��Y<�5[<�(]<+._<�a<�b<��c<+:d<1@d<_�c<�<c<�b<mb<��a<��a<�Mb<\�b<�?c<�}c<�tc<�'c<$�b<G/b<��a<��a<kb<#�b<�\c<J�c<�Cd<�"d<�zc<�Kb<P�`<�^<z�\<��Z<�EY<�7X<��W<�W<��X<�Z<��[<��]<��_<��a<\c<�c<�Hd<'d<ԩc<@�b<�Zb<��a<��a<�b<<ub<��b<�Yc<��c<yac<�c<�b<�b<d�a<:�a<�Ib<��b<5�c<�d<rHd<~�c<�$c<3�a<Y`<n^<�\<�BZ<R�X<��W<��W<�X<�Y<��Z<�}\<5�^<�r`<�b<�[c<(d<GBd<o�c<�kc<��b<S&b<��a<��a<�b<8�b<dc<�ic<?zc<dCc<�b<�Tb<��a<��a<��a<exb<>"c<��c<�2d</:d<�c<O�b<(:a<�__<�[]<ld[<ɱY<psX<��W<Z�W<UX<��Y<('[<9]<]_<��`<n�b<��c< d<!d<K�c<�c<�lb<\�a<&�a<�a<_$b<1�b<�c<�Rc<�Ic<��b<�b<Sb<׭a<-�a<��a<��b<X2c<h�c<od<��c<Nc<3b<|`<��^<p�\<�Z<SY<YX<ΐW<��W<։X<��Y<ި[<��]<��_<ma<��b<��c<_d<*�c<Usc<�b<	#b<�a<b�a<��a<';b<��b<�c<�Gc<�'c<H�b<*Jb<�a<k�a<:�a<�  �  KQa<��a<�`b<�b<c<��b<�b<��`<��^<��\<�Z<��X<O'W<�.V<��U<5WV<yuW<!Y<�([<HQ]<]_<Za<Rb<��b<�!c<��b<�Gb<H�a<�La<�<a<i�a<q=b<�
c<3�c<�>d<`Vd<Jd<Fgc<�b<�a<aa<�Da<��a<@b<�b<�c<4c<��b<i�a<�H`<^^<�<\<� Z<GX<��V<�(V< V<��V<�X<�Y<[\<�1^<&(`<��a<`�b<�Gc<�@c<��b<�Bb<��a<�ja<}a<��a<جb<Byc<�!d<�zd<�nd<��c<�Ic<i{b<��a<Fia<
na<U�a<�^b<��b<�Fc<i3c<.�b<aja<�_<$�]<��[<f�Y<��W<��V<�V<�OV<�5W<ӶX<��Z<s�\<��^<��`<�&b<�c<�Qc<�$c<Ȧb<�b<ґa<�aa<*�a<�(b<a�b<�c<�Hd<��d<�Sd<U�c<�c<�;b<�a<�`a<t�a<��a<�b<�c<�Oc<�c<�Cb</�`<�_<]<��Z<K�X<�VW<v]V<V<҄V<C�W<�LY<mS[< {]<��_<�<a<�xb<C%c<�Fc<��b<�kb<��a<�oa<�_a<Y�a<_`b<�-c<��c<ad<�xd<�)d<?�c<�b<�a<�~a<�`a<%�a<�*b<|�b<g2c<YFc<��b<��a<�S`<�f^<�B\<($Z<�GX<��V<y$V<V<�V<`X<F�Y<�[<'^<�`<��a<w�b<�*c<�!c<��b<�b<�a<�Da<�Ua<�a<J�b<�Nc<�c<�Od<QCd<��c<�c<gPb<Ƞa<�>a<�Ca<�a<4b<��b<�c<�c<�jb<0=a<�_<4�]<�c[<�UY<J�W<dmV<�U<�V<mW<�X<�qZ<W�\<��^<5�`<��a<��b<[c<��b<(pb<j�a<�Ya<�(a<�]a<��a<�b<}{c<�d<�Fd<Ud<��c<��b<�b<�ja<q*a<�  �  �`<�a<=�a<z#b<�bb<T-b<�ga<A`<�:^<F\<�Y<��W<�(V<�!U<��T<=MU<{V<G<X<�ZZ<w�\<U�^<Yl`<<�a<|Kb<�db<�b<��a<		a<�`<��`<mxa<�[b<n]c<�@d<U�d<��d<�d<��c<~�b<�a<�$a< �`<<�`<�[a<��a<�]b<�{b<Kb<�"a<_�_<�]<�w[< FY<�UW<��U<�U<gU<.�U<,W<�Y<?D[<f|]<}_<da<�b<��b<��b<Nb<r�a<na<�`<�:a<Y�a<��b<��c<��d<xe<�e<Q~d<��c<�b<6�a<�a<�`<)%a<��a<�-b<��b<-~b<�a<I�`<;_<]<��Z<��X<r�V<�U<�
U<�AU<v5V<\�W<�Y<�\<�3^<	`<:|a<�Rb<��b<�cb<��a<�[a<Q�`<U�`<�ga<�3b<�1c<M%d<��d<�e<��d<�<d<�Mc<Mb<�xa<�`<D�`<La<��a<
Vb<��b<�^b<��a<�?`<�j^<NE\<�
Z<Q�W<XV<kPU<�U<�zU<��V<�gX<+�Z<�\<��^<��`<��a<�pb<H�b<�6b<N�a<I,a< �`<�
a<a�a<�~b<^�c<�cd<��d<	e<̱d<��c<��b<�a<mBa<J�`<�a<hta<Gb<crb<"�b<F)b<t0a<}�_<��]<�}[<�IY<�VW<��U<�U<_U<��U<�W<(Y<�2[<�h]<�f_<��`<� b<�sb<Vbb<�a<jga<��`<��`<a<��a<�b<��c<�{d<F�d<��d<�Rd<Wvc<�tb<e�a<��`<��`<��`<=xa<�b<�]b<�Rb<Ͻa<5�`<N�^<3�\<�Z<wsX<$�V<�dU<@�T<�U<V<��W<0�Y<��[<}�]<��_<�Ga<�b<bb<�-b<�a<9$a<5�`<��`<'.a<��a<�b<��c<��d<�d<[�d<�d<kc<Eb<�Aa<��`<�  �  CDb<tlb<��b<�b<}�b<�Yb<h�a<�h`<k�^< H]<�[<�Z<	�X<�5X< X<�TX<+Y<�mZ<_�[<*�]<�L_<��`<)�a<
b<��b<��b<-�b<�kb<lLb<�[b<U�b<c<|�c<7d<��d<Z�d<�gd<��c<rcc<��b<~b<Wb<fb<J�b<��b<O�b<o�b<q?b<VWa<6`<!�^<��\<�7[<"�Y<�X<b9X<�2X<��X<��Y<3[<j�\<gd^<��_<mJa<�?b<W�b<mc<��b<��b<ʉb<�wb<s�b<�b<*xc<*
d<H�d<>�d<O�d<�jd<��c<�Tc<��b<'�b<�rb<��b<��b<D�b<��b<��b<�b<�a<�_<^<�X\<{�Z<%yY<�X<3X<�YX<�Y<�'Z<p�[<#J]<[�^<u`<�a<|b<��b<�c<��b<ǧb<�|b<�yb<Y�b<�c<b�c<�5d<\�d<+�d<]�d<RCd<'�c<['c<��b<�{b<�xb<��b<��b<�b<��b<̊b<��a<�`<#_<jw]<7�[<JKZ<fY<dcX<\-X<A�X<�VY<��Z<n&\<?�]<�t_<��`<Z�a<a�b<w�b<�b<��b<Ǝb<ob<.~b<��b<#@c<]�c<�Xd<��d<$�d<��d<>d<�c<G�b<�b<�qb<	b<y�b<�b<��b<��b<qNb<da<�`<&�^<;�\<�:[<��Y<0�X<5X<+,X<B�X<0�Y<�[<ɣ\<jQ^<]�_<�2a<>&b<��b<��b<�b<W�b<�fb<Sb<�sb<@�b<jPc<��c<-Zd<��d<��d<�@d<۽c<�*c<Ǭb<4^b<�Hb<�cb<H�b<��b<
�b<D�b<��a<#�`<nv_<4�]<�)\<��Z<�HY<�dX<_X<�'X<�X< �Y<[n[<�]<��^<;A`<�ta<�Gb<յb<w�b<��b<fqb<�Eb<\Bb<Pwb<2�b<�nc<��c<Vfd<F�d<�nd<0d<�c<��b<��b<QFb<�  �  �[b<��b<��b<��b<��b<�b<6�a<��`<Z_<x]<��[<�UZ<�-Y<kvX<�AX<�X<�gY<E�Z<�/\<{�]<y_</�`<��a<:�b<Z�b<��b<��b<=�b<�ab<@fb<��b<+c<��c<�d<�dd<-ud<:@d<_�c<$Oc<a�b<B�b<�gb<��b<��b<��b<mc<��b<�hb<J�a<�<`<��^<
]<n[<Z<Y<�zX<�tX<��X<_�Y<�K[<S�\<��^<2$`<vta<^ib<��b<�,c<�c<��b<\�b<x�b<�b<��b<)ec<��c<�\d<&�d<��d<pEd<��c<�Dc<��b<f�b<҆b<��b<��b< c<p$c<��b<�9b<C0a<�_<u6^<ԋ\<F�Z<��Y< �X<�tX<ܚX<�DY<�aZ<��[<�z]<�!_<�`<��a<I�b<c<�+c<�c<��b<9�b<;�b<��b<c<\�c<d<�vd<ĝd<0~d<� d<ўc<^c<��b<��b<ߏb<�b<u�b<�'c<Pc<��b<��a<��`<L_<v�]<� \<��Z<J\Y<V�X<oX<��X<ޓY<M�Z<�Y\<�^<%�_<U	a<b<��b<�c<�c<[�b<@�b<M�b<��b<��b<=1c<u�c<=4d<ƅd<�d<a`d<��c<�mc<��b<B�b<m�b<��b<��b<�c<�&c<��b<�wb<�a<�F`<�^<�]</q[<�Z<HY<�vX<�mX<��X<��Y<�=[<��\<�^<�`<�\a<�Ob<��b<�c<F�b<>�b<k�b<eb<Uzb<�b<n=c<?�c<�3d<�od<�fd<}d<��c<�c<��b<sgb<�\b<|�b<o�b<��b<�b<��b<pb<za<��_<"^<�\\<k�Z< �Y<��X<�BX<�hX<bY<	/Z<}�[<KG]<�^<Al`<Ȟa<�pb<>�b<L�b<��b<C�b<K^b<�Pb<�yb<��b<�Wc<�c<�=d<�dd<�Ed<��c<Qgc<��b<��b<mSb<�  �  �b<�b<2c<ec<Zc<�b<�0b<�
a<S�_<^<�h\<��Z<��Y<2Y<��X<+OY<#Z<�H[<��\<�`^<�_<nXa<Skb<c<kc<�fc<�+c<N�b<��b<�b<��b<��b<gCc<5�c<A�c<�c<,�c<�tc<�c<>�b<\�b<&�b<w�b<�c<�ac<��c<]_c<��b<i�a<|�`<C4_<t�]<
\<��Z<n�Y<#8Y</2Y<b�Y<^�Z<��[<Du]<_<ϝ`<��a<��b<Dmc<<�c<��c<�>c<��b<�b<�b<��b<�)c<)�c<u�c<od<ld<��c<�uc<"c<��b<N�b<��b<<�b<�Jc<*�c<ޖc<�Rc< �b<B�a<\K`<��^<]<T�[<�dZ<��Y<�2Y<KWY<��Y<X	[<Go\<^<��_<�a<�Gb<Pc<c�c<��c<^nc<"c<��b<g�b<��b<�b<Ic<N�c<H�c<�d<>d<E�c<�Sc<9�b<R�b<�b<K�b<xc<�dc<�c<|�c<�'c<Xab<�:a<�_<�0^<̗\<|*[<
Z<%`Y<T-Y<�{Y<'DZ<�s[<��\<�^<K`<�a<��b<�Ac<��c<��c<Oc<Y c<��b<��b<3�b<�c<=ec<��c<vd<�d<E�c<�c<*.c<z�b<M�b<��b<W�b<�.c<wc<˗c<�pc<��b<b<ݿ`<C<_<�]<6\<C�Z<��Y<�3Y<[+Y<�Y<��Z<n�[<�d]<_<��`<P�a<��b<�Qc<��c<edc<6c<��b<��b<e�b<�b<c<�fc<m�c<��c<��c<��c< Lc<&�b<˛b<[~b<��b<'�b<� c<�_c<�kc<F'c<ׁb<cya<�`<�^<��\<_n[<�3Z<[^Y<Y<%Y<P�Y<m�Z<<\<��]<m_<��`<�b<��b<�Rc<Nfc<�8c<��b<��b<wb<�|b<³b<nc<zuc<l�c<>�c<��c<I�c<dc<��b<g�b<�ub<�  �  ��b<�[c<��c<+�c<��c<��c<�b<Ȱa<hN`<�^<�K]<��[<
�Z<)VZ<(Z<�pZ<)[<�@\<��]<x$_<r�`<S�a<�	c<ιc<1d<�c<k�c<:Nc<��b<E�b<s|b<)�b<h�b<(�b<c<!c<�c<_�b<��b<\�b<x�b<S�b<+c<��c<r�c<X d<��c<�zc<'�b<f_a<��_<�h^<�\<��[<��Z<�^Z<]YZ<��Z<�[<��\<UI^<��_<-Ia</�b<U{c<�
d<f:d<�d<��c<_Vc<[�b<%�b<#�b<Q�b<��b<�'c<8Fc<�Ac<�c<��b<�b<ʢb<��b<�c<�ic<}�c<�!d<�3d<��c<\Lc<dIb<-�`<�|_<9�]<��\<<s[<�Z<�ZZ<x|Z<�[<�
\<ZU]<��^<�V`<�a<>�b<�c<�$d<56d<��c<�c<�1c<��b<�b<�b<��b<�c<$4c<Hc<�7c<>
c<��b<z�b<��b<��b<%c<3�c<��c<%1d<�(d<��c<� c<��a<K~`<��^<�z]<�(\<�$[<^�Z<�UZ<ٝZ<FU[<2l\<��]<�M_<��`<�#b<E0c<`�c<�,d<9#d<��c<Qqc<H
c<��b<��b</�b<4�b<�c<:9c<�Ac<�&c<��b<Ҿb<��b<T�b<��b<�Cc<��c<�
d<�3d<d<��c<ңb<�ia<��_<=n^<7�\<%�[<��Z<fZZ<�RZ<6�Z<"�[<v�\<�8^<��_<�3a<�sb<�ac<(�c<�d<y�c<��c<�3c<�b<��b<{�b<��b<*�b<��b<�c<�c<��b<��b<*�b<�xb<��b<��b<e?c<)�c< �c<�d<�c< c<bb<e�`<bN_<��]<lc\<iB[<�~Z<�(Z<JZ<��Z<��[<"]<q�^<+#`<�a<+�b<��c<�c<d<6�c<�fc<��b<b�b<Xsb<�pb<m�b< �b<z�b<�c<��b<p�b<��b<�sb<�qb<ܜb<�  �  �>c<m�c<�Pd<әd<��d<2d<�qc<�^b<�a<q�_<!Z^<�1]<`P\<��[<�[<��[<�|\<�o]<�^<�`<�da<ͦb<�c<gWd<>�d<H�d<�Ad<J�c<�)c<ɣb<�?b<+b<��a<��a<�a<��a< �a<,�a<S�a<�'b<K{b<��b<X�c<@d<�d<s�d<W�d<d<�;c<�b<ʽ`<.\_<�^<� ]<2<\<��[<��[<�/\<@�\<��]<CA_<`�`<% b<1c<d<4�d<��d<ծd<�Ed<e�c<&c<_�b<(Rb<~#b<Mb<b<�$b<b#b<�b<"b<�&b<^b<ҽb<Ac<��c<�\d<�d<��d<M�d<(�c<i�b<��a<�W`<Y�^<7�]<v�\<8\<��[<�[<Vn\<G]<�h^<��_<4a<%ob<ˉc<�Td<�d<Z�d<6�d<�d<��c<h�b<m�b<
<b<�b<�b<�b<�$b<t b<�b<�b<}5b<>zb<��b<�rc<�d<>�d<��d<�d<ocd<E�c<3�b<�Ca<5�_<��^<�`]<@\<F�[<��[<\<!�\<��]<��^<h,`<(�a<j�b<��c<$}d<+�d<��d<�ed<q�c<�Lc<B�b<�ab<'&b<pb<Rb<b<�b<b<Gb<zb<�Db<
�b<�c<�c<80d<�d<��d<a�d<�'d<{Hc<Gb<��`<�a_<�^<�]<W:\<��[<��[<L&\<�\<��]<�0_<u�`<��a<�c<s d<��d<&�d<d�d<g$d<��c<�c<�b<�+b<�a<�a<>�a<��a<��a<��a<E�a<�a<4b<�b<
c<Z�c<M2d<_�d<��d<�bd<��c<9�b<��a<�(`<��^<ލ]<k�\<��[<Ѡ[<w�[<h;\<�]<M5^<$�_<��`<G;b<�Uc<u d<Y�d<I�d<�Zd<��c<�Mc<^�b<�Mb<!b<��a<K�a<Q�a<��a<s�a<W�a<��a<%�a<�Db<,�b<�  �  ?gc<�#d<��d<�
e<�e<�d<z�c<��b<��a<Z�`< r_<��^<n�]<c]<4E]<�t]<��]<O�^<��_<��`<�b<�1c<9$d<�d<e<De<[�d<!d< Gc<A�b<�a<[La<^�`<&�`<{�`<�`<��`<_�`<�"a<^�a<{:b<m�b<|�c<�sd<I�d<�.e<Qe<k�d<νc<��b<Ya<�O`<�=_<�`^<��]<�u]<�r]<�]<1R^<+_<�:`<ka<s�b<�c<.�d<4e<Ie<$e<�d<+�c<\0c<�pb<�a<Ra<a<��`<��`<��`<��`<Ja<�fa<��a<i�b<Xc<Wd<�d<|)e<�Ce<�e<ped<E{c<]b<)a<K�_<�^<�2^<��]<�w]<��]<��]<˛^<6�_<}�`<�a<(c<d<��d<�4e<�Be<��d<_kd<M�c<�b<�3b<e�a<<0a<��`<��`<v�`<�`<�`<\&a<m�a<4 b<p�b<#�c<�Vd<2�d<�<e<9e<��d<d<% c<��a<J�`<ء_<�^<��]<ȑ]<`s]<l�]<g^<3�^<��_<oa<�7b<�Yc<Kd<�d<7=e<�,e<�d<\*d<�ic<��b<8�a<Lna<a<}�`<j�`<Y�`<_�`<X�`<�@a<D�a<Vb<�c<�c<׊d<Je<�Ae<He<8�d<^�c<�b<@�a</U`<�@_<$a^<�]<pq]<�k]<ĳ]<sF^<�_<1*`<"Xa<G�b<��c<�wd<��d<�+e<��d<ցd<��c<Mc<WKb<�a<�*a<��`<�`<��`<�`<��`<�`<�<a<��a<xkb<.c< �c<��d<��d<}e<��d<�8d<�Mc<�.b<�`<u�_<m�^<�^<�}]<�E]<�Z]<Ѽ]<oh^<�S_<�o`<S�a<@�b<
�c<��d<H e<�e<M�d<�5d<�{c<P�b<e�a<�ea<N�`<��`<h�`<w�`<S�`<ɯ`<��`<PXa<��a<ˠb<�  �  Tc<4d<{�d<X4e<�1e<��d<�)d<Hc<dLb<kSa<Nw`<��_<�L_<�_<��^<w_<�d_<s�_<I�`<m�a<�b<j�c<t[d<��d<aBe<�0e<P�d<�d<{)c<�,b<�7a<�b`<�_<�J_<�_<�_<E+_<��_<�`<��`<�a<��b<�c<5�d<9e<�Xe<8e<8�d<d<qc<�b<�&a<xY`<��_<�S_< _<�_<TO_<ٳ_<\N`<a<�	b<	c<;�c<D�d<0Fe<#se<�Be<7�d<��c<�c<�b<Ha<KO`<�_<\X_<l+_<n0_<�g_<g�_<�t`<�Da<�7b<%5c<� d<m�d<�Qe<<ne< .e<�d<^�c<)�b<n�a<g�`<M.`<T�_<J_<,&_<4_<�t_<��_<(�`<�ka<�bb<�_c<�Ed<j�d<1_e<Ile<te<P~d<��c<[�b<1�a<��`<_`<2�_<RB_<�&_<�<_<|�_<�`<w�`<y�a<�b<c<gd<�e<3fe<Zce<�e<�Zd<�xc<�|b<��a<>�`<��_<|_<�5_<,"_<M@_<_<�`<��`<��a<G�b<��c<��d<�e<�ge<qUe<+�d<M4d<YLc<^Ob<�Ya<��`<��_<�k_<�._<�#_<�J_<w�_<�5`<��`<��a<��b<}�c<��d< 1e<�ke<�He<��d<�d<�c<yb<,a<�\`<N�_<�Q_<�_<�_<F_<�_<7@`<�a<��a<��b<��c<ͩd<�*e<�Ue<�#e<@�d<)�c<��b<��a<��`<(`<�_<�/_<a_<_<9>_<��_<�J`<�a<�b<c<s�c<ٲd<�&e<�Be<�e<6nd<��c<��b<$�a<L�`<m�_<�o_<�_<��^<_<UA_<q�_<y``<8a</b<�+c<�d<%�d<�*e<q7e<;�d<�Hd<�mc<�sb<4xa<��`<��_<iY_<�
_<��^<_<yN_<�_<�`<L^a<�Xb<�  �  ��b<��c<�d<
e<�e<��d<#d<�]c<�b<�a<=Ta<e�`<�`<\�`<	�`<��`<�`<a<Ssa<�b<^�b<��c<�Fd<
�d<�e<ye<5�d<��c<��b<�a<�k`<@R_<�j^<��]<gf]<�U]<��]<�^<��^<��_<la<cRb<�oc<�Wd<��d<s.e<Be<�d<��c<M:c<�xb<��a<�Oa<9�`<�`<�`<B�`<6�`<u�`<�La<��a<�rb<�4c<��c<ŧd<�e<�He<ze<7�d<Ϋc<R�b<�aa<�3`<"(_<�S^<��]<�~]<�]<�]<c{^<�\_<�q`<��a<��b<�c<X�d<@'e<wDe<�e<8�d<8�c<S
c<�Mb<b�a<D=a<��`<��`<<�`<��`<��`<�a<�ya<0b<͵b<�zc<j:d<��d<46e<�Ae<��d<�Ed<Qc<�,b<~�`<�_<^�^<�^<Ϣ]<�w]<	�]<�^<y�^<�_<��`<�	b<S1c<�,d<j�d<�;e<:e<��d<�Kd<c�c<��b<mb<e�a<Ya<��`<��`<ѹ`<��`<O�`<�/a<�a<7b<��b<�c<Ond<e�d<>e<"+e<.�d<E�c<��b<��a<Ս`<t_<B�^<��]<�]<v]<s�]<0:^<;_<�`<�8a<Mlb<@�c<Qnd<ce<OAe<!e<��d<�d<wDc<Ȁb<N�a<�Ra<��`<*�`<��`<o�`<�`<��`<�>a<j�a<�_b<�c<F�c<]�d<�e<�+e<M�d<Yid<d�c<�pb<�<a<�`<_<,^<f�]<�U]<�]]<��]<�Q^<�2_<�G`<�xa<��b<��c<��d<$�d<�e<g�d<,Wd<]�c<��b<db<�a<a<��`</�`<O�`<��`</�`<��`<�Ea<I�a<ہb<�Fc<Sd<f�d<�e<(e<��d<ld<0c<��a<��`<�_<
�^<z�]<Pk]<W@]<�b]<��]<A�^<N~_<ɠ`<��a<�  �  dnb<�}c<�9d<�d<͗d<oKd<��c<�7c<+�b<Bb<H�a<O�a<Y�a<��a<��a<��a<a�a<=�a<hb<�Yb<��b<�]c<��c<�hd<�d<��d<�!d<�Rc<5b<��`<	�_<�0^<[]<@\<�[<��[<] \<Ү\<�]<@�^<�N`<E�a<u�b<�c<@}d<��d<p�d<�Ad<�c<c&c<h�b<hHb< b<�b<zb<�b<�b<Ub<b<�b<Lb<
�b<	'c<Q�c< Id< �d<D�d<?�d<ud<�&c<��a<Q�`<B7_<�]<.�\<x4\<�[<��[<7T\<f]<�4^<��_<��`<�8b<^c<q7d<l�d<��d<<�d<#+d<��c<.
c</�b<Cb<tb<�b<\b<�"b<U b<�b<Tb<c-b<�kb<��b<�Zc<��c<Ard<��d<��d<�|d<��c<`�b<T�a<�`<��^<ő]<Y�\<
\<7�[<��[<��\</s]<Ǟ^<z�_<�Xa<աb<q�c<ld<��d<0�d<�|d<w�c<�hc<��b<�rb<�/b<~b<Fb<�b< b<0b<b<b<A9b<��b<��b<��c<Gd<?�d<��d<V�d<�Ed</vc<	Xb<^a<1�_<uR^<�4]<a\<��[<��[<�\<_�\<��]<�
_<	j`<�a<� c<��c<��d<|�d<,�d<[Pd<P�c<�0c<1�b<�Mb<b<8b<�	b<Zb<�b<b<X b<�b<�;b<@�b<�c<�c<�/d<��d<��d<'�d<��c<;c<F�a<]s`<9_<��]<u�\<#\<C�[<��[<�*\<��\<�
^<-W_<��`<�b<�3c<�d<2�d<æd<�pd<��c<�lc<?�b<dcb<yb<�a<��a<��a<��a<��a<6�a<i�a<e�a<�7b<��b<�&c<��c<>d<s�d<D�d<�Gd<��c<��b<:Ja<C�_<.�^<�Z]<)l\<��[< �[<��[<W\<7=]<bi^<��_<�$a<�  �  1�a<S�b<�c<��c<z�c<��c<�Vc<�b<7�b<sb<xb<��b<�b<bc<�c<N�b<G�b<z�b<1vb<}{b<��b<(c<�tc<]�c<hd<9�c<Ѓc<��b<׃a<�`<&�^<]<�[<��Z<�SZ<�9Z<��Z<�`[<φ\<��]<^v_<X�`<f@b<�?c<��c<�d<�	d<�c<Pc<�b<٨b<5�b<F�b<K�b<�c<�3c<7c<�c<�b<Ĳb<�b<�b<��b<�Vc<��c<cd<�9d<�d<psc<�b<�;a<��_<�<^<��\<��[<�Z<$dZ<qZ<$�Z<��[<T]<��^<;`<��a<�b<=�c<*d<�6d<�	d<<�c<@c<R�b<\�b<%�b<��b<G�b<�+c<�Ec<y;c<�c<��b<e�b<��b<��b<pc<�}c<��c<1,d<�1d<��c<;*c<�b<��`<<>_<�]<:`\<�M[<ڛZ<�YZ<��Z<�4[<W=\<O�]<�_<G�`<��a<c<H�c<�+d<�.d<��c<��c<�c<��b<��b<��b<�b<2	c<-5c<4Cc<-c<9�b<��b<J�b<��b<x�b< 1c<��c<�c<01d<(d< �c<5�b<٦a<`<`<L�^<�<]<~�[<�[<VtZ<�YZ<ܵZ<[<I�\<�^<x�_<a<�Xb<-Vc<h�c<�1d<hd<x�c<w\c<)�b<��b<��b<@�b<��b<�c<X/c<>0c<�c<R�b<��b<|�b<%�b<��b<�?c<��c<�c<ld<��c<�Rc<�]b<�a<��_<	^<%�\<"z[<ȤZ<p;Z<HZ<��Z<s�[<��\<�e^<H�_<W[a<��b<gnc<��c<�
d<��c<�~c<�c<0�b<Z}b<Ksb<��b<��b<��b<7c<�c<�b<��b<Gzb<�pb<z�b<Z�b<{Ic<\�c<��c<*�c<��c<�b<T�a<��`<�_<y�]<j)\<�[<�dZ<�"Z<XZ<[�Z<�\<]]<^�^<Sa`<�  �  �a<^=b<d�b<�\c<�cc<�.c<��b<\�b<3wb<�b<��b<R%c<�c<��c<r�c<��c<�uc<�c<��b<��b<gb<ͬb<o�b<�Dc<^pc<�Xc<,�b<�b<��`<�b_<�]<�3\<X�Z<g�Y<Z.Y<)Y<wY<VSZ<C�[<]<M�^<�E`<ԝa<��b<Bc<-�c<�rc<�2c<��b<�b<��b<Y�b<gc<Ikc<H�c<+d<�	d<��c<}c<c<]�b<��b<�b<I�b<�>c<��c<3�c<ic<��b<��a<X�`<�_<Xg]<_�[<ؖZ<�Y<�<Y<�JY<��Y<`�Z<�/\<ٿ]<�\_<R�`<�b<��b<�yc<U�c<�vc<-c<��b<��b<{�b<^�b<�5c<�c<��c<�d<�	d<+�c<#dc<�c<��b<v�b<{�b<�
c<�Yc<+�c<`�c<�@c<}�b<Xta<.`<y^<h�\<xf[<u;Z<RyY<f1Y<�jY< Z<i@[<��\<#J^<
�_<Oa<pb<�0c<@�c<�c<�_c<�c<=�b<�b<��b<��b<�Uc<T�c<�d<�d<��c<��c<�=c<��b<�b<��b<��b<X c<�kc<D�c<�}c<o
c<^3b<	�`<D�_<4�]<`U\<��Z<U�Y<�NY<2Y<0�Y<�qZ<��[<_3]<Q�^<#_`<�a<�b<�Vc<Ӕc<c�c<Ac<�b<��b<R�b<��b<\c<�kc<^�c<� d<�d<��c<eqc<�
c<�b<�b<�b<�b<�%c<Ric<�c<Jc<�b<Իa<�k`<��^<~A]<��[<PoZ<ˆY<Y<�!Y<_�Y<�Z<+\<�]<3_<#�`<,�a<��b<HNc<Noc<�Ic<z�b<S�b<��b<P}b<X�b<0c<�ic<�c<e�c<�c<�c<�/c<��b<ȉb<Nub<]�b<��b<d%c<�^c<�_c<>c<qVb<�>a<k�_<�B^< �\<�/[<�Z<�BY<��X<�4Y<��Y<�
[<�{\<�^<3�_<�  �  �`<��a<j�b<w�b<��b<	�b<<�b<c[b<�Vb<6�b<!�b<rc<��c<3Md<
id<�>d<��c<�Uc<j�b<�|b<VWb<hb<�b<��b< c<J�b<rb<�a<d`<"�^<�;]<#�[<*Z<�Y<�qX<$TX<�X<+�Y<�Z<��\<�1^<��_<(a<D-b<Y�b<�c<<c<0�b<[�b<psb<��b<*�b<�:c<��c<=;d<Ӄd<�d<�Id<��c<lRc<N�b<��b<��b<g�b< �b<�c<\+c<U�b<,ab<nha<K`<��^<��\<�@[<�Y<��X<�~X<��X<�!Y<�,Z<��[<83]<N�^<�c`<��a<��b<9c<�*c<Gc<��b<N�b<��b<|�b<��b<fwc<i�c<hd<`�d<��d<p2d<��c<N/c<}�b<��b<��b<��b<:�b<�$c<~!c<	�b<�b<��`<��_<�]<�H\< �Z<��Y<��X<sX<�X<�mY<c�Z<|\<��]<�d_<�`<[�a<��b<.c<&c<2�b<>�b<P�b<q�b<�b<�c<��c<#d<J}d<��d<�md<�d<0�c<�c<��b<��b< �b<��b<�c<&c<a
c<h�b<��a<�`<�_<^]<߻[<gKZ<�4Y<�X<�sX<3�X<w�Y<q[<��\<�L^<J�_<@a<�Cb<��b<�"c<�c<��b<��b<w}b<\�b<��b<�=c<H�c<Q9d<td<@�d<�@d<H�c<ZDc<��b<ہb<�mb<A�b<��b<��b<6c<g�b<�@b<PFa<��_<�]^<��\<[<��Y<��X<7VX<�dX<��X<"Z<�j[<u	]<[�^<�9`<'za<�\b<��b<s�b<v�b<�b<�jb<%Ub<6tb<��b<{Ec<��c<�4d<�fd<�Rd<F�c<U�c<�b<>�b<�Xb<oWb<��b<�b<��b<�b<[�b<��a<�`<�[_<�]<~\<|�Z<�SY<�X<�<X<2yX<�7Y<�eZ<��[<k�]<�0_<�  �  'z`<�a<Dab<�b<+�b<��b<�jb<�Db<Jb<݈b<��b<
�c<�d<�vd<\�d<�fd<��c<lc<F�b<�yb<UHb<Ob<�|b<7�b<#�b<�b<�Hb<qa<�8`<��^<2]<�d[<��Y<Q�X<|0X<�X<;~X<iY<��Z<S\<9^<Ξ_<��`<�b<�b<��b<��b<X�b<Axb<�_b<yb<#�b<�Kc<~�c<�`d<��d<�d<5pd<��c<�dc<��b<L�b<pb<K�b<�b<��b<c< �b<�7b<Q>a<��_<:T^<b�\<�	[<i�Y<c�X<9=X<0LX<��X<��Y<�^[<]<��^<}8`<�za<J^b<��b<�c<��b<Ϯb<`b<Utb<�b<'c<k�c<rd<��d<��d<��d<hVd<��c<y=c<��b<��b<�ub<Зb<9�b<��b<�b<ۣb<�a</�`<e_<~�]<	\<e�Z<_MY<~X<c1X<�nX<40Y<>bZ<3�[<�]<�7_<O�`<��a<b�b<��b<��b<��b<��b<�ub<{b<��b<�+c<��c<*Fd<��d<�d<�d<)d<��c<�c<�b<�rb<Bxb<��b<1�b<"�b<��b<.mb<��a< \`<N�^<U-]<n�[<@Z<3�X<�PX<\2X<U�X<R�Y<��Z<Po\<,^<Z�_<�a<b<��b<(�b<�b<ѻb<��b<�ib<b<|�b<�Nc<�c<�^d<6�d<>�d<�fd<!�c<�Vc<K�b<�zb<[b<&ob<��b<S�b<��b<�b<b<6a<%�_<�/^<�\<�Z<�Y<M�X<�X<A#X<��X<l�Y<�4[<D�\<��^<I`<=Pa<V3b<c�b<g�b<��b<(�b<�Pb<�Db<�ob<��b<wZc<��c<r\d<��d<�|d<6"d<��c<+	c<W�b<_Mb<�Ab<�cb<�b<T�b<��b<2ob<+�a<�`<b/_<��]<��[<�SZ<�Y<wGX<��W<m8X<K�X<�,Z<E�[<�]]<�_<�  �  �`<��a<j�b<w�b<��b<	�b<<�b<c[b<�Vb<6�b<!�b<rc<��c<3Md<
id<�>d<��c<�Uc<j�b<�|b<VWb<hb<�b<��b< c<J�b<rb<�a<d`<"�^<�;]<#�[<*Z<�Y<�qX<$TX<�X<+�Y<�Z<��\<�1^<��_<(a<D-b<Y�b<�c<<c<0�b<[�b<psb<��b<*�b<�:c<��c<=;d<Ӄd<�d<�Id<��c<lRc<N�b<��b<��b<g�b< �b<�c<\+c<U�b<,ab<nha<K`<��^<��\<�@[<�Y<��X<�~X<��X<�!Y<�,Z<��[<83]<N�^<�c`<��a<��b<9c<�*c<Gc<��b<N�b<��b<|�b<��b<fwc<i�c<hd<`�d<��d<p2d<��c<N/c<}�b<��b<��b<��b<:�b<�$c<~!c<	�b<�b<��`<��_<�]<�H\< �Z<��Y<��X<sX<�X<�mY<c�Z<|\<��]<�d_<�`<[�a<��b<.c<&c<2�b<>�b<P�b<q�b<�b<�c<��c<#d<J}d<��d<�md<�d<0�c<�c<��b<��b< �b<��b<�c<&c<a
c<h�b<��a<�`<�_<^]<߻[<gKZ<�4Y<�X<�sX<3�X<w�Y<q[<��\<�L^<J�_<@a<�Cb<��b<�"c<�c<��b<��b<w}b<\�b<��b<�=c<H�c<Q9d<td<@�d<�@d<H�c<ZDc<��b<ہb<�mb<A�b<��b<��b<6c<g�b<�@b<PFa<��_<�]^<��\<[<��Y<��X<7VX<�dX<��X<"Z<�j[<u	]<[�^<�9`<'za<�\b<��b<s�b<v�b<�b<�jb<%Ub<6tb<��b<{Ec<��c<�4d<�fd<�Rd<F�c<U�c<�b<>�b<�Xb<oWb<��b<�b<��b<�b<[�b<��a<�`<�[_<�]<~\<|�Z<�SY<�X<�<X<2yX<�7Y<�eZ<��[<k�]<�0_<�  �  �a<^=b<d�b<�\c<�cc<�.c<��b<\�b<3wb<�b<��b<R%c<�c<��c<r�c<��c<�uc<�c<��b<��b<gb<ͬb<o�b<�Dc<^pc<�Xc<,�b<�b<��`<�b_<�]<�3\<X�Z<g�Y<Z.Y<)Y<wY<VSZ<C�[<]<M�^<�E`<ԝa<��b<Bc<-�c<�rc<�2c<��b<�b<��b<Y�b<gc<Ikc<H�c<+d<�	d<��c<}c<c<]�b<��b<�b<I�b<�>c<��c<3�c<ic<��b<��a<X�`<�_<Xg]<_�[<ؖZ<�Y<�<Y<�JY<��Y<`�Z<�/\<ٿ]<�\_<R�`<�b<��b<�yc<U�c<�vc<-c<��b<��b<{�b<^�b<�5c<�c<��c<�d<�	d<+�c<#dc<�c<��b<v�b<{�b<�
c<�Yc<+�c<`�c<�@c<}�b<Xta<.`<y^<h�\<xf[<u;Z<RyY<f1Y<�jY< Z<i@[<��\<#J^<
�_<Oa<pb<�0c<@�c<�c<�_c<�c<=�b<�b<��b<��b<�Uc<T�c<�d<�d<��c<��c<�=c<��b<�b<��b<��b<X c<�kc<D�c<�}c<o
c<^3b<	�`<D�_<4�]<`U\<��Z<U�Y<�NY<2Y<0�Y<�qZ<��[<_3]<Q�^<#_`<�a<�b<�Vc<Ӕc<c�c<Ac<�b<��b<R�b<��b<\c<�kc<^�c<� d<�d<��c<eqc<�
c<�b<�b<�b<�b<�%c<Ric<�c<Jc<�b<Իa<�k`<��^<~A]<��[<PoZ<ˆY<Y<�!Y<_�Y<�Z<+\<�]<3_<#�`<,�a<��b<HNc<Noc<�Ic<z�b<S�b<��b<P}b<X�b<0c<�ic<�c<e�c<�c<�c<�/c<��b<ȉb<Nub<]�b<��b<d%c<�^c<�_c<>c<qVb<�>a<k�_<�B^< �\<�/[<�Z<�BY<��X<�4Y<��Y<�
[<�{\<�^<3�_<�  �  1�a<S�b<�c<��c<z�c<��c<�Vc<�b<7�b<sb<xb<��b<�b<bc<�c<N�b<G�b<z�b<1vb<}{b<��b<(c<�tc<]�c<hd<9�c<Ѓc<��b<׃a<�`<&�^<]<�[<��Z<�SZ<�9Z<��Z<�`[<φ\<��]<^v_<X�`<f@b<�?c<��c<�d<�	d<�c<Pc<�b<٨b<5�b<F�b<K�b<�c<�3c<7c<�c<�b<Ĳb<�b<�b<��b<�Vc<��c<cd<�9d<�d<psc<�b<�;a<��_<�<^<��\<��[<�Z<$dZ<qZ<$�Z<��[<T]<��^<;`<��a<�b<=�c<*d<�6d<�	d<<�c<@c<R�b<\�b<%�b<��b<G�b<�+c<�Ec<y;c<�c<��b<e�b<��b<��b<pc<�}c<��c<1,d<�1d<��c<;*c<�b<��`<<>_<�]<:`\<�M[<ڛZ<�YZ<��Z<�4[<W=\<O�]<�_<G�`<��a<c<H�c<�+d<�.d<��c<��c<�c<��b<��b<��b<�b<2	c<-5c<4Cc<-c<9�b<��b<J�b<��b<x�b< 1c<��c<�c<01d<(d< �c<5�b<٦a<`<`<L�^<�<]<~�[<�[<VtZ<�YZ<ܵZ<[<I�\<�^<x�_<a<�Xb<-Vc<h�c<�1d<hd<x�c<w\c<)�b<��b<��b<@�b<��b<�c<X/c<>0c<�c<R�b<��b<|�b<%�b<��b<�?c<��c<�c<ld<��c<�Rc<�]b<�a<��_<	^<%�\<"z[<ȤZ<p;Z<HZ<��Z<s�[<��\<�e^<H�_<W[a<��b<gnc<��c<�
d<��c<�~c<�c<0�b<Z}b<Ksb<��b<��b<��b<7c<�c<�b<��b<Gzb<�pb<z�b<Z�b<{Ic<\�c<��c<*�c<��c<�b<T�a<��`<�_<y�]<j)\<�[<�dZ<�"Z<XZ<[�Z<�\<]]<^�^<Sa`<�  �  dnb<�}c<�9d<�d<͗d<oKd<��c<�7c<+�b<Bb<H�a<O�a<Y�a<��a<��a<��a<a�a<=�a<hb<�Yb<��b<�]c<��c<�hd<�d<��d<�!d<�Rc<5b<��`<	�_<�0^<[]<@\<�[<��[<] \<Ү\<�]<@�^<�N`<E�a<u�b<�c<@}d<��d<p�d<�Ad<�c<c&c<h�b<hHb< b<�b<zb<�b<�b<Ub<b<�b<Lb<
�b<	'c<Q�c< Id< �d<D�d<?�d<ud<�&c<��a<Q�`<B7_<�]<.�\<x4\<�[<��[<7T\<f]<�4^<��_<��`<�8b<^c<q7d<l�d<��d<<�d<#+d<��c<.
c</�b<Cb<tb<�b<\b<�"b<U b<�b<Tb<c-b<�kb<��b<�Zc<��c<Ard<��d<��d<�|d<��c<`�b<T�a<�`<��^<ő]<Y�\<
\<7�[<��[<��\</s]<Ǟ^<z�_<�Xa<աb<q�c<ld<��d<0�d<�|d<w�c<�hc<��b<�rb<�/b<~b<Fb<�b< b<0b<b<b<A9b<��b<��b<��c<Gd<?�d<��d<V�d<�Ed</vc<	Xb<^a<1�_<uR^<�4]<a\<��[<��[<�\<_�\<��]<�
_<	j`<�a<� c<��c<��d<|�d<,�d<[Pd<P�c<�0c<1�b<�Mb<b<8b<�	b<Zb<�b<b<X b<�b<�;b<@�b<�c<�c<�/d<��d<��d<'�d<��c<;c<F�a<]s`<9_<��]<u�\<#\<C�[<��[<�*\<��\<�
^<-W_<��`<�b<�3c<�d<2�d<æd<�pd<��c<�lc<?�b<dcb<yb<�a<��a<��a<��a<��a<6�a<i�a<e�a<�7b<��b<�&c<��c<>d<s�d<D�d<�Gd<��c<��b<:Ja<C�_<.�^<�Z]<)l\<��[< �[<��[<W\<7=]<bi^<��_<�$a<�  �  ��b<��c<�d<
e<�e<��d<#d<�]c<�b<�a<=Ta<e�`<�`<\�`<	�`<��`<�`<a<Ssa<�b<^�b<��c<�Fd<
�d<�e<ye<5�d<��c<��b<�a<�k`<@R_<�j^<��]<gf]<�U]<��]<�^<��^<��_<la<cRb<�oc<�Wd<��d<s.e<Be<�d<��c<M:c<�xb<��a<�Oa<9�`<�`<�`<B�`<6�`<u�`<�La<��a<�rb<�4c<��c<ŧd<�e<�He<ze<7�d<Ϋc<R�b<�aa<�3`<"(_<�S^<��]<�~]<�]<�]<c{^<�\_<�q`<��a<��b<�c<X�d<@'e<wDe<�e<8�d<8�c<S
c<�Mb<b�a<D=a<��`<��`<<�`<��`<��`<�a<�ya<0b<͵b<�zc<j:d<��d<46e<�Ae<��d<�Ed<Qc<�,b<~�`<�_<^�^<�^<Ϣ]<�w]<	�]<�^<y�^<�_<��`<�	b<S1c<�,d<j�d<�;e<:e<��d<�Kd<c�c<��b<mb<e�a<Ya<��`<��`<ѹ`<��`<O�`<�/a<�a<7b<��b<�c<Ond<e�d<>e<"+e<.�d<E�c<��b<��a<Ս`<t_<B�^<��]<�]<v]<s�]<0:^<;_<�`<�8a<Mlb<@�c<Qnd<ce<OAe<!e<��d<�d<wDc<Ȁb<N�a<�Ra<��`<*�`<��`<o�`<�`<��`<�>a<j�a<�_b<�c<F�c<]�d<�e<�+e<M�d<Yid<d�c<�pb<�<a<�`<_<,^<f�]<�U]<�]]<��]<�Q^<�2_<�G`<�xa<��b<��c<��d<$�d<�e<g�d<,Wd<]�c<��b<db<�a<a<��`</�`<O�`<��`</�`<��`<�Ea<I�a<ہb<�Fc<Sd<f�d<�e<(e<��d<ld<0c<��a<��`<�_<
�^<z�]<Pk]<W@]<�b]<��]<A�^<N~_<ɠ`<��a<�  �  Tc<4d<{�d<X4e<�1e<��d<�)d<Hc<dLb<kSa<Nw`<��_<�L_<�_<��^<w_<�d_<s�_<I�`<m�a<�b<j�c<t[d<��d<aBe<�0e<P�d<�d<{)c<�,b<�7a<�b`<�_<�J_<�_<�_<E+_<��_<�`<��`<�a<��b<�c<5�d<9e<�Xe<8e<8�d<d<qc<�b<�&a<xY`<��_<�S_< _<�_<TO_<ٳ_<\N`<a<�	b<	c<;�c<D�d<0Fe<#se<�Be<7�d<��c<�c<�b<Ha<KO`<�_<\X_<l+_<n0_<�g_<g�_<�t`<�Da<�7b<%5c<� d<m�d<�Qe<<ne< .e<�d<^�c<)�b<n�a<g�`<M.`<T�_<J_<,&_<4_<�t_<��_<(�`<�ka<�bb<�_c<�Ed<j�d<1_e<Ile<te<P~d<��c<[�b<1�a<��`<_`<2�_<RB_<�&_<�<_<|�_<�`<w�`<y�a<�b<c<gd<�e<3fe<Zce<�e<�Zd<�xc<�|b<��a<>�`<��_<|_<�5_<,"_<M@_<_<�`<��`<��a<G�b<��c<��d<�e<�ge<qUe<+�d<M4d<YLc<^Ob<�Ya<��`<��_<�k_<�._<�#_<�J_<w�_<�5`<��`<��a<��b<}�c<��d< 1e<�ke<�He<��d<�d<�c<yb<,a<�\`<N�_<�Q_<�_<�_<F_<�_<7@`<�a<��a<��b<��c<ͩd<�*e<�Ue<�#e<@�d<)�c<��b<��a<��`<(`<�_<�/_<a_<_<9>_<��_<�J`<�a<�b<c<s�c<ٲd<�&e<�Be<�e<6nd<��c<��b<$�a<L�`<m�_<�o_<�_<��^<_<UA_<q�_<y``<8a</b<�+c<�d<%�d<�*e<q7e<;�d<�Hd<�mc<�sb<4xa<��`<��_<iY_<�
_<��^<_<yN_<�_<�`<L^a<�Xb<�  �  ?gc<�#d<��d<�
e<�e<�d<z�c<��b<��a<Z�`< r_<��^<n�]<c]<4E]<�t]<��]<O�^<��_<��`<�b<�1c<9$d<�d<e<De<[�d<!d< Gc<A�b<�a<[La<^�`<&�`<{�`<�`<��`<_�`<�"a<^�a<{:b<m�b<|�c<�sd<I�d<�.e<Qe<k�d<νc<��b<Ya<�O`<�=_<�`^<��]<�u]<�r]<�]<1R^<+_<�:`<ka<s�b<�c<.�d<4e<Ie<$e<�d<+�c<\0c<�pb<�a<Ra<a<��`<��`<��`<��`<Ja<�fa<��a<i�b<Xc<Wd<�d<|)e<�Ce<�e<ped<E{c<]b<)a<K�_<�^<�2^<��]<�w]<��]<��]<˛^<6�_<}�`<�a<(c<d<��d<�4e<�Be<��d<_kd<M�c<�b<�3b<e�a<<0a<��`<��`<v�`<�`<�`<\&a<m�a<4 b<p�b<#�c<�Vd<2�d<�<e<9e<��d<d<% c<��a<J�`<ء_<�^<��]<ȑ]<`s]<l�]<g^<3�^<��_<oa<�7b<�Yc<Kd<�d<7=e<�,e<�d<\*d<�ic<��b<8�a<Lna<a<}�`<j�`<Y�`<_�`<X�`<�@a<D�a<Vb<�c<�c<׊d<Je<�Ae<He<8�d<^�c<�b<@�a</U`<�@_<$a^<�]<pq]<�k]<ĳ]<sF^<�_<1*`<"Xa<G�b<��c<�wd<��d<�+e<��d<ցd<��c<Mc<WKb<�a<�*a<��`<�`<��`<�`<��`<�`<�<a<��a<xkb<.c< �c<��d<��d<}e<��d<�8d<�Mc<�.b<�`<u�_<m�^<�^<�}]<�E]<�Z]<Ѽ]<oh^<�S_<�o`<S�a<@�b<
�c<��d<H e<�e<M�d<�5d<�{c<P�b<e�a<�ea<N�`<��`<h�`<w�`<S�`<ɯ`<��`<PXa<��a<ˠb<�  �  �>c<m�c<�Pd<әd<��d<2d<�qc<�^b<�a<q�_<!Z^<�1]<`P\<��[<�[<��[<�|\<�o]<�^<�`<�da<ͦb<�c<gWd<>�d<H�d<�Ad<J�c<�)c<ɣb<�?b<+b<��a<��a<�a<��a< �a<,�a<S�a<�'b<K{b<��b<X�c<@d<�d<s�d<W�d<d<�;c<�b<ʽ`<.\_<�^<� ]<2<\<��[<��[<�/\<@�\<��]<CA_<`�`<% b<1c<d<4�d<��d<ծd<�Ed<e�c<&c<_�b<(Rb<~#b<Mb<b<�$b<b#b<�b<"b<�&b<^b<ҽb<Ac<��c<�\d<�d<��d<M�d<(�c<i�b<��a<�W`<Y�^<7�]<v�\<8\<��[<�[<Vn\<G]<�h^<��_<4a<%ob<ˉc<�Td<�d<Z�d<6�d<�d<��c<h�b<m�b<
<b<�b<�b<�b<�$b<t b<�b<�b<}5b<>zb<��b<�rc<�d<>�d<��d<�d<ocd<E�c<3�b<�Ca<5�_<��^<�`]<@\<F�[<��[<\<!�\<��]<��^<h,`<(�a<j�b<��c<$}d<+�d<��d<�ed<q�c<�Lc<B�b<�ab<'&b<pb<Rb<b<�b<b<Gb<zb<�Db<
�b<�c<�c<80d<�d<��d<a�d<�'d<{Hc<Gb<��`<�a_<�^<�]<W:\<��[<��[<L&\<�\<��]<�0_<u�`<��a<�c<s d<��d<&�d<d�d<g$d<��c<�c<�b<�+b<�a<�a<>�a<��a<��a<��a<E�a<�a<4b<�b<
c<Z�c<M2d<_�d<��d<�bd<��c<9�b<��a<�(`<��^<ލ]<k�\<��[<Ѡ[<w�[<h;\<�]<M5^<$�_<��`<G;b<�Uc<u d<Y�d<I�d<�Zd<��c<�Mc<^�b<�Mb<!b<��a<K�a<Q�a<��a<s�a<W�a<��a<%�a<�Db<,�b<�  �  ��b<�[c<��c<+�c<��c<��c<�b<Ȱa<hN`<�^<�K]<��[<
�Z<)VZ<(Z<�pZ<)[<�@\<��]<x$_<r�`<S�a<�	c<ιc<1d<�c<k�c<:Nc<��b<E�b<s|b<)�b<h�b<(�b<c<!c<�c<_�b<��b<\�b<x�b<S�b<+c<��c<r�c<X d<��c<�zc<'�b<f_a<��_<�h^<�\<��[<��Z<�^Z<]YZ<��Z<�[<��\<UI^<��_<-Ia</�b<U{c<�
d<f:d<�d<��c<_Vc<[�b<%�b<#�b<Q�b<��b<�'c<8Fc<�Ac<�c<��b<�b<ʢb<��b<�c<�ic<}�c<�!d<�3d<��c<\Lc<dIb<-�`<�|_<9�]<��\<<s[<�Z<�ZZ<x|Z<�[<�
\<ZU]<��^<�V`<�a<>�b<�c<�$d<56d<��c<�c<�1c<��b<�b<�b<��b<�c<$4c<Hc<�7c<>
c<��b<z�b<��b<��b<%c<3�c<��c<%1d<�(d<��c<� c<��a<K~`<��^<�z]<�(\<�$[<^�Z<�UZ<ٝZ<FU[<2l\<��]<�M_<��`<�#b<E0c<`�c<�,d<9#d<��c<Qqc<H
c<��b<��b</�b<4�b<�c<:9c<�Ac<�&c<��b<Ҿb<��b<T�b<��b<�Cc<��c<�
d<�3d<d<��c<ңb<�ia<��_<=n^<7�\<%�[<��Z<fZZ<�RZ<6�Z<"�[<v�\<�8^<��_<�3a<�sb<�ac<(�c<�d<y�c<��c<�3c<�b<��b<{�b<��b<*�b<��b<�c<�c<��b<��b<*�b<�xb<��b<��b<e?c<)�c< �c<�d<�c< c<bb<e�`<bN_<��]<lc\<iB[<�~Z<�(Z<JZ<��Z<��[<"]<q�^<+#`<�a<+�b<��c<�c<d<6�c<�fc<��b<b�b<Xsb<�pb<m�b< �b<z�b<�c<��b<p�b<��b<�sb<�qb<ܜb<�  �  �b<�b<2c<ec<Zc<�b<�0b<�
a<S�_<^<�h\<��Z<��Y<2Y<��X<+OY<#Z<�H[<��\<�`^<�_<nXa<Skb<c<kc<�fc<�+c<N�b<��b<�b<��b<��b<gCc<5�c<A�c<�c<,�c<�tc<�c<>�b<\�b<&�b<w�b<�c<�ac<��c<]_c<��b<i�a<|�`<C4_<t�]<
\<��Z<n�Y<#8Y</2Y<b�Y<^�Z<��[<Du]<_<ϝ`<��a<��b<Dmc<<�c<��c<�>c<��b<�b<�b<��b<�)c<)�c<u�c<od<ld<��c<�uc<"c<��b<N�b<��b<<�b<�Jc<*�c<ޖc<�Rc< �b<B�a<\K`<��^<]<T�[<�dZ<��Y<�2Y<KWY<��Y<X	[<Go\<^<��_<�a<�Gb<Pc<c�c<��c<^nc<"c<��b<g�b<��b<�b<Ic<N�c<H�c<�d<>d<E�c<�Sc<9�b<R�b<�b<K�b<xc<�dc<�c<|�c<�'c<Xab<�:a<�_<�0^<̗\<|*[<
Z<%`Y<T-Y<�{Y<'DZ<�s[<��\<�^<K`<�a<��b<�Ac<��c<��c<Oc<Y c<��b<��b<3�b<�c<=ec<��c<vd<�d<E�c<�c<*.c<z�b<M�b<��b<W�b<�.c<wc<˗c<�pc<��b<b<ݿ`<C<_<�]<6\<C�Z<��Y<�3Y<[+Y<�Y<��Z<n�[<�d]<_<��`<P�a<��b<�Qc<��c<edc<6c<��b<��b<e�b<�b<c<�fc<m�c<��c<��c<��c< Lc<&�b<˛b<[~b<��b<'�b<� c<�_c<�kc<F'c<ׁb<cya<�`<�^<��\<_n[<�3Z<[^Y<Y<%Y<P�Y<m�Z<<\<��]<m_<��`<�b<��b<�Rc<Nfc<�8c<��b<��b<wb<�|b<³b<nc<zuc<l�c<>�c<��c<I�c<dc<��b<g�b<�ub<�  �  �[b<��b<��b<��b<��b<�b<6�a<��`<Z_<x]<��[<�UZ<�-Y<kvX<�AX<�X<�gY<E�Z<�/\<{�]<y_</�`<��a<:�b<Z�b<��b<��b<=�b<�ab<@fb<��b<+c<��c<�d<�dd<-ud<:@d<_�c<$Oc<a�b<B�b<�gb<��b<��b<��b<mc<��b<�hb<J�a<�<`<��^<
]<n[<Z<Y<�zX<�tX<��X<_�Y<�K[<S�\<��^<2$`<vta<^ib<��b<�,c<�c<��b<\�b<x�b<�b<��b<)ec<��c<�\d<&�d<��d<pEd<��c<�Dc<��b<f�b<҆b<��b<��b< c<p$c<��b<�9b<C0a<�_<u6^<ԋ\<F�Z<��Y< �X<�tX<ܚX<�DY<�aZ<��[<�z]<�!_<�`<��a<I�b<c<�+c<�c<��b<9�b<;�b<��b<c<\�c<d<�vd<ĝd<0~d<� d<ўc<^c<��b<��b<ߏb<�b<u�b<�'c<Pc<��b<��a<��`<L_<v�]<� \<��Z<J\Y<V�X<oX<��X<ޓY<M�Z<�Y\<�^<%�_<U	a<b<��b<�c<�c<[�b<@�b<M�b<��b<��b<=1c<u�c<=4d<ƅd<�d<a`d<��c<�mc<��b<B�b<m�b<��b<��b<�c<�&c<��b<�wb<�a<�F`<�^<�]</q[<�Z<HY<�vX<�mX<��X<��Y<�=[<��\<�^<�`<�\a<�Ob<��b<�c<F�b<>�b<k�b<eb<Uzb<�b<n=c<?�c<�3d<�od<�fd<}d<��c<�c<��b<sgb<�\b<|�b<o�b<��b<�b<��b<pb<za<��_<"^<�\\<k�Z< �Y<��X<�BX<�hX<bY<	/Z<}�[<KG]<�^<Al`<Ȟa<�pb<>�b<L�b<��b<C�b<K^b<�Pb<�yb<��b<�Wc<�c<�=d<�dd<�Ed<��c<Qgc<��b<��b<mSb<�  �  ͷb<��b<��b<��b<��b<_Cb<�a<^�`<|�_<�K^<�]<\<�2[<R�Z<ʈZ<x�Z<;][<PB\<�]]</�^<��_<��`<��a<�gb<��b<��b<:�b<J�b<l�b<��b<k�b<S
c<>Hc<�c<�c<��c<?�c< gc<x*c<��b<��b<��b<�b<��b<V�b<�b<7�b<],b<�fa<�e`<<_<�^<��\<l�[<�[<,�Z<�Z<�[<��[<��\<b�]< '_<V`<_a<�-b<y�b<�c<�c<�c<g�b<��b<.�b<�c<�Fc<��c<)�c<��c<2�c<��c<(uc<�6c<c<��b<��b<��b<�c<�c<��b<��b<�b<)a<�`<6�^<y�]<�\<��[< [<1�Z<r�Z<&P[<�\<�)]<LZ^<M�_<a�`<�a<�eb<��b<gc<c<�c<��b<��b<C�b<sc<8Zc<ߖc<��c<��c<�c<ڜc<�`c<�$c<��b<#�b<=�b<� c<c<Bc<��b<�sb<��a<��`<��_<�z^<dG]<6\<_`[<m�Z<R�Z<X�Z<`�[<�l\<k�]<ƽ^<Q�_<N	a<��a<�b<)�b<>c<`c<��b<��b<��b<��b<�+c< ic<��c<�c<�c<��c<�c<bGc<]c<?�b<��b<��b<�c<ic<Dc<e�b<v:b<�ra<�o`<�C_<�^<��\<��[<�[<�Z<`�Z<�
[<��[<�\<r�]<�_<�A`<�Ha<cb<��b<��b<��b<��b<�b<�b<0�b<��b<� c<�]c<��c<��c<Ϊc<�c<ILc<�c<��b<{�b<��b<�b<��b<b�b<:�b<zsb<�a<��`<��_<t�^<~]<�]\<�q[<��Z<S�Z<"�Z<u[<��[<R�\<�'^<z`_<K�`<za<2b<Хb<��b<2�b<��b<ȸb<��b<��b<p�b<�"c<}_c<$�c<a�c<�c<=fc<�*c<�b<��b<��b<�  �  �b<�b<��b<R�b<�b<�[b<��a<��`<ȡ_<?m^<C>]<�0\<\^[<�Z<öZ<��Z<�[<%j\<l�]<�^<?�_<��`<&�a<#�b<��b<gc<r�b<H�b<�b<W�b<��b<��b<Q1c<=fc<��c<w�c<�{c<oMc<�c<U�b<��b<��b<f�b<R�b<�c<Cc<��b<Eb<�a<L�`<d[_<�&^<j ]<�\<SL[<�Z<��Z<_@[<��[<^�\<�^<�F_<�r`<aya<�Fb<U�b<fc<�-c<�c<uc<R�b<.�b<Ec<�4c<vkc<כc<n�c<��c<1�c<y]c<l&c<�b<|�b<��b<c<n c</*c<�c<��b<b<�Ca<$4`<�_<��]<��\<�[<?-[<%�Z<>[<(|[<�F\<UO]<S|^<�_<<�`<g�a<)~b<W�b<&c<9+c<�c<��b<�b<b�b<bc<�Ec<�{c<�c<;�c<5�c<&�c<>Kc<�c<��b<p�b<z�b<�c<�'c<�&c<��b<�b<��a<x�`<��_<�^<�l]<�^\<��[<)	[<R�Z<�[<<�[<��\<�]<��^<�`<c$a<b<E�b<Mc<#%c<�c<�c<\�b<9�b<G�b<�c<1Rc<��c<��c<�c<<�c<Pkc<m4c<c<V�b<��b<��b<-c<'c<mc<�b<*Sb<��a<�`<�b_<�+^<A]<m\<rJ[<��Z<<�Z<a7[<d�[<��\<��]<m4_<i^`<�ba<@.b<Ҷb<�b<�c<��b<�b<��b<2�b</�b<�c<�Dc<\tc<p�c<!�c<�hc<�4c<j�b<^�b<<�b<u�b<t�b<��b<��b<(�b<��b<D�a<�a<`<��^<�]<z�\<E�[<��Z<A�Z<��Z<qJ[<�\<]<�I^<_<%�`<�a<wJb<I�b<��b<T�b<M�b<��b<ϲb<��b<g�b<mc<zDc<�oc< �c<<sc<�Jc<(c<�b<��b<M�b<�  �  �b<c<)c<q0c<ac<s�b<z�a<�a<��_<
�^<^�]<��\<�[<6a[<q=[<,v[<�\<�\<��]<_<H;`<AIa<
&b<�b<Sc<	;c<�,c<c<�b<�b<��b<��b<��b<Cc<�)c<|/c<6c<��b<��b<��b<�b<��b<�b<�+c<3Ic<gCc<ic<�b<h�a<��`<`�_<��^<dn]<z}\<��[<(o[<9k[<��[<ll\<�Y]<Ds^<��_<�`<I�a<A�b<$c<Xc<ec<-Lc<�!c<��b<��b<�b<-�b<c<�@c<�Sc<�Pc<�8c<�c<��b<��b<��b<��b<)(c<vPc<cc<�Kc<]�b<ydb<�a<W�`<�__<�6^<i&]<�G\<�[<�n[<�[<��[< �\<ɺ]<^�^<�`<!a<�b<R�b<2c<�ac<k_c<>c<tc<��b<6�b<&�b<�c<$*c<�Hc<�Tc<�Jc<|-c<�	c<��b<��b<��b<~c<�7c<[c<�ac<<8c<��b<i$b<�;a<�%`<��^<��]<��\<�
\<m�[<j[<+�[<#0\<y]<�^<�:_<c`<$pa<Lb<O�b<�Ac<�^c<�Oc<�(c<b�b<��b<�b<��b<uc<�/c<�Ic<�Nc<�=c<ic<|�b<G�b<��b<��b<�c<pAc<<]c<�Uc<�c<.�b<U�a<p�`<׺_<�^<:q]<�}\<��[<�j[<�d[<��[<a\<�K]<Vc^<m�_<��`<Ьa<�sb<��b<�;c<�Fc<f,c<� c<,�b<�b< �b</�b<��b<:c<�+c<n(c<c<��b<��b<}�b<@�b<[�b<��b<�&c<�8c<!c<(�b<�8b<�ba<2Y`<�1_<T^<+�\<\<��[<�=[<zW[<*�[<�\<k�]<��^<�_<��`<`�a<��b<��b<-c<�*c<�c<��b<��b<��b<@�b<��b<��b<Bc<�c<�c<��b<��b<T�b<0�b<ɷb<�  �  N�b<�8c<�nc<y�c<�_c<��b<�Yb<%{a<�s`<sZ_<�I^<1Z]<&�\<�/\<6\<�B\<��\<d�]<�^<z�_<�`<�a<��b<
 c<)tc<�c<�nc<�4c<�b<ƴb<�b<�wb<~wb<��b<d�b<M�b<@�b<�~b<n{b<�b<l�b<�b<#c<�ec<�c<�c<�ac<��b<�2b<Ea<�5`<�_<O^<�7]<�\<�?\<Y<\<�\<l(]<�^<�	_<�#`<�7a<�,b<e�b<nc<��c<=�c<S�c<�Hc<�c<(�b<�b<��b<��b<��b<�b<{�b<ǧb<�b<1�b<$�b<��b<nc<lTc<��c<�c<�c<�Uc<U�b<��a<��`< �_<��^<��]<]<�|\<�@\<TX\<��\<�s]<u^^<�l_<��`<��a<�ub<M!c<�c<ٳc<a�c<�sc<�0c<��b<��b<j�b<�b<��b<�b<�b<ڮb<Z�b<��b<�b<t�b<#�b<�'c<Kkc<��c<۲c<|�c<.c<ŉb<��a<�`<d�_<dx^<p�]<��\<]\<�;\<o\<D�\<��]<ΰ^<Q�_<��`<��a<ïb<TEc<��c<ܭc<ّc<�Wc<Xc<��b<��b<�b<P�b<W�b<M�b<��b<ܦb<��b<9�b<Ţb<��b<�b<�:c<�{c<�c<6�c<�qc<��b<�>b<�Na<F=`<�"_<!^<+8]<�\<�;\<�5\<�\<]<�]<��^<�`<�#a<b<��b<�Sc<E�c<'�c<�hc<�'c<��b<E�b<��b<�xb<�zb<)�b<�b</�b<0b<Lub<9tb<�b<G�b<�b<�*c<�fc<��c<(wc<q*c<p�b<�a<H�`<&�_<I�^<t�]<~�\<CL\<�\<�&\<��\<yA]<,^<1:_<�S`<o^a<�Bb<��b<�Vc<|c<�qc<�>c<��b<��b<'�b<�lb<fb<�lb<�vb<|b<xb<�mb<�fb<�kb<Ʉb<&�b<�  �  �c<�ec<��c<��c<�c<�`c<��b<��a<�a<�`<m_<M:^<͗]<�4]<�]<�E]<'�]<�g^<�F_<A`<�@a<�.b<��b<a�c<��c<T�c<��c<\c<��b<q�b<)@b<��a<�a<�a<D�a<��a<P�a<��a<��a<�'b<vb<U�b<�=c<��c<[�c<��c<!�c<�Pc<��b<��a<��`<�_<�^<	 ^<��]<�G]<�D]<W�]<b^<]�^<i�_<ʿ`<�a</�b<�Tc<s�c<�d<�c<��c<wfc<� c<��b<LQb<�b<�a<	�a<��a<�a<��a<x�a<	 b<*^b<��b<.c<�xc<��c<��c<Q�c<7�c<Q1c<�qb<0�a<��`<��_<��^<��]<j~]<0J]<�^]<\�]<�V^<;'_<T`<4a<Kb<�b<��c<S�c<.d<�c<l�c<�Cc<��b<R�b<&:b<Xb<0�a<��a<��a<��a<��a<�b<�2b<Qxb<��b<7c<-�c<s�c<�d<��c<^�c<��b<�'b<�3a<�3`<+>_<�h^<��]<lb]<�E]<�q]<��]<��^<�p_<j`<�ha<�Ub<c<̦c<5�c<D�c<��c<�~c<$c<Y�b<�ab<� b<��a<k�a<�a<��a<��a<R�a<�b<�Cb<V�b<=�b<�Tc<M�c<G�c<�c<0�c<�^c<��b<��a<C�`<!�_<��^< ^<��]<fC]<9>]<\�]<^<��^<��_<��`<��a<ĉb<S<c<
�c<X�c<��c<ןc<HEc<\�b<�|b<e,b<��a<r�a<��a<ݱa<رa<r�a<��a<�a<5b<B�b<��b<�Nc<��c<z�c<y�c<Ҋc<Mc</Eb<�Za<�[`<�__<"}^<t�]<�M]<�]<-]<[�]<Z$^<��^<��_<C�`<&�a<��b<�Qc<a�c<��c<j�c<Tnc<:c<�b<
Lb<�b<��a<C�a<��a<¡a<�a<^�a<��a<��a<�Cb<�b<�  �  ��b<�yc<A�c<�d<�c<j�c<W%c<�jb<$�a<ϴ`<��_<�0_<��^<�Y^<�B^<kg^<��^<-W_<�`<9�`<��a<M�b<�Nc<D�c<Vd<�d<�c<�ic<q�b<kXb<O�a<:ba<}a<��`<Ǳ`<�`<��`<��`<�=a<�a<,$b<R�b<�=c<�c<�
d<)d<Pd<��c<�c<�Bb<ha<�`<�_<� _<Ĭ^<�o^<�m^<��^<�_<S�_<_�`<�\a<�:b<yc<��c<�d<�@d<g+d<��c<�ic<Y�b<�Sb<��a<Vja<Ja<�`<��`<�`<��`<^)a</}a<��a<eob<��b<�c<��c<�2d<;d<d<�c<�b<�b<�.a<�V`<p�_<C_<��^<=t^<�^<�^<�P_<w�_<]�`<^�a<��b<�Dc<I�c<?,d<�@d<�d<�c<8<c<�b<�%b<\�a<�Ka<Xa<v�`<;�`<^�`<a<?Ba<��a<6b<��b<�+c<��c<d<=d<�/d<��c<gUc<C�b<��a<��`<f`<j__<��^<h�^<p^<��^<[�^<2�_<�<`<sa<��a<��b<Muc<��c<4d<�2d<n�c<��c<�c<Wzb<��a<\�a<7,a<?�`<��`<3�`<_�`<ca<Za<��a<c>b<"�b<�Tc<��c<�d<�:d<Pd<��c<�c<�Lb<ooa<�`<��_<d!_<۪^<lk^<g^<��^<B_<��_<~p`<�Ja<�&b<�b<��c<U�c<�$d<pd<�c<�Hc<ݽb<)0b<��a<�Da<��`<��`<�`<�`<6�`<� a<ITa<��a<%Fb<�b<dYc<��c<Hd<d<}�c<�]c<8�b<"�a<C a<�'`<�h_<��^<�m^<�B^<S^<��^<z_<��_<��`<^ya<�Rb<�c<��c<[�c<Md</�c<�c<�c<�yb<x�a<�ua</a<��`<��`<��`<�`<�`<�a<�ja<��a<�jb<�  �  ��b<Ahc<��c<�d<d<p�c<jac<��b<jb<�Va<�`<�'`<��_<d�_<av_<��_<<�_<JE`<��`<��a<�9b<��b<L�c<�c<�)d<�d<��c<zRc<�b<v�a<�Da<�`<� `<�_<��_<υ_<��_<��_<�j`<@a<&�a<�hb<�c<��c<�d<�>d<A(d<��c<~Lc<T�b<Y�a<7=a<�`< $`<��_</�_<�_<D�_<s`<ߙ`<}5a<g�a<�b<�Lc<�c<�7d<�Wd<�5d<��c<�Hc<'�b<��a<&5a<U�`<$`<@�_<<�_<װ_<��_<�9`<��`<�Wa<�
b<��b<�hc<��c<�@d<�Td<a'd<O�c<�)c<�yb<��a<a<U�`<�`<(�_<��_<<�_<��_<L`<�`< ua<�)b<��b<u�c<�d<�Jd<�Sd<3d<t�c<�c<�]b<�a<��`<�n`<r`<��_<	�_<��_<��_<p``<��`<X�a<KHb<��b<��c<�d<�Nd<�Ld<�
d<��c<��b<�;b<	�a<&�`<]V`<`�_<V�_<ˣ_<r�_<L`<�p`<� a<(�a<bb<Vc<�c<�d<�Nd<Bd<P�c<buc<F�b<db<efa<��`<3A`<H�_<��_<ݤ_<
�_<"`<�`<�a<B�a<��b<�/c<:�c<�'d<�Pd<18d<��c<CXc<�b<��a<JBa<ǣ`<n$`<��_<�_<R�_<K�_<'`<G�`<�%a<S�a<ϋb<�6c<��c<�d<�;d<d<	�c<�'c<�yb<6�a<qa<�v`<��_<#�_<��_<ň_<2�_</`<��`<�.a<C�a<~�b<�>c<d�c<d<�)d<��c<��c<��b</Lb<)�a<��`<fR`<"�_<�_<v_<<�_<8�_<u`<D�`<5Ba<��a<e�b<Pc<]�c<�d<�d<��c<�vc<��b<5(b<qa<w�`<k8`<��_<%�_<�q_<��_<��_<+`<Ѷ`<!^a<�b<�  �  Otb<^-c<ʵc<>d<�
d<��c<"tc<}�b<eb<�a<�ga<�a<��`<§`<>�`<<�`<�`<�a<T�a<x�a<Јb<
c<h�c<��c<d<��c<?�c<�c<,Rb<�xa<ԛ`<	�_<y#_<>�^<'_^<�R^<��^<8�^<)�_<�D`<�a<��a<��b<}yc<z�c<�%d<6d<H�c<�hc<�b<�Ub<��a<6ga<�a<D�`<��`<��`<��`<ma<5ea<\�a<�Sb<��b<Zlc<��c<u,d<@d<�d<M�c<� c<�4b<�Wa<t}`<[�_<7_<S�^<�y^<�^<��^<�8_<��_<�`<r�a<�ab<]&c<6�c<} d<�?d<ed<�c<`Pc<��b<t9b<ϼa<�Wa<�a<��`<`�`<t�`<��`<�4a<؍a<� b<��b<5c<3�c<d<�:d<k8d<��c<�rc<��b<��a<�a<7`<=~_<��^<2�^<Ft^<~�^<��^<�k_<D `<��`<��a<,�b<�_c<��c<�2d<�;d< d<P�c<i"c<��b<�b<��a<�:a<~�`<��`<��`<B�`<_a<Ka<�a<''b<��b<�=c<4�c<|d<;d<7#d<��c<�5c<�tb<��a<T�`<�_<D_<c�^<�~^<�q^<ş^<�_<��_<�_`<�8a<Sb<�b<�c<+d<�7d<+d<�c<Ytc<��b<]b<��a<�ia<a<W�`<��`<=�`<��`<$	a<�Wa<��a<�Ab<��b<Vc<n�c<5d<�#d<�c<ۅc<��b<�b<%4a<�X`<Γ_<��^<O�^<�Q^<�W^<��^<_<�_<	�`<1]a<8b<��b<�c<��c<cd<��c<��c<.#c<�b<�
b<]�a<�'a<9�`<n�`<��`<F�`<}�`<a<�Za<��a<gTb<��b<�ec<��c<�d<`d<,�c<>c<��b<%�a<9�`<,`<H_<��^<�^^<'>^<�X^<1�^<y6_<��_<��`<��a<�  �  b<��b<�fc<޼c<P�c<��c<�ac<��b<��b<�Ab<�a<"�a<��a<��a<C�a<�a<˺a<z�a<?b<]Wb<��b<c<6{c<��c<��c<i�c<�Tc<رb<d�a<��`<��_<��^<�'^<x�]<�8]<)]<Qb]<K�]<q�^<�~_<|`<�za<"db<�!c<l�c<��c<:�c<j�c<�_c<��b<q�b<�Hb<�b<��a<�a<v�a<O�a<,�a< �a<�b<�Kb<��b<* c<�fc<W�c<�c<% d<��c<:Oc<�b<A�a<ڸ`<]�_<X�^<R^<�]<NP]<X]<��]<d9^<�_<�_<�`<��a<t�b<Qmc<��c<Pd<��c<(�c<LRc<_�b<,�b<�Bb<b<�a<}�a<F�a<Q�a<��a<4�a<�(b<"kb<�b<�&c<ۉc<��c<fd<�c<�c<�c<�Ob<�`a<�a`<�h_<�^<��]<cr]<�I]<0j]<��]<�v^<	N_<xD`<Da<�5b<�c<��c<�c<(d<x�c<�c<�/c<e�b<Pqb<q,b<@�a<��a<�a<�a<Q�a<S�a<3b<8b<B�b<��b<oCc<.�c<��c<�c<��c<dxc<��b<��a<�a<``<�_<*H^<��]<X]<�G]<s�]<��]<��^<�_<�`<��a<${b<B7c<�c<��c<�c<3�c<�kc<^c<��b<�Mb<bb<X�a<�a<.�a<��a<6�a<��a<Nb<*<b<��b<��b<�Pc<�c<��c<�c<&�c<�/c<8xb<	�a<j�`<ؖ_<�^<�]<�i]<�(]<.0]<o]<�^<�^<�_<��`<m�a<��b<Cc<9�c<�c<��c<��c<�$c<?�b<G_b<�b<��a<�a<��a<K�a<��a<��a<]�a<��a<8b<�b<A�b<vVc<	�c<��c<�c<�rc<�b<�b<�+a<,`<%3_<�V^<��]<]<]<�]<�4]<��]<�A^<�_<�`<�a<�  �  7�a<rcb<>c<�bc<ׁc<�lc<$6c<�b<��b<+�b<�mb<4jb<+rb<�|b<��b<Q{b<]qb<�kb<�sb<�b<�b<[c<7Jc<!|c<�c<u\c< �b<�Ab<�[a<P`<�6_<�*^<WC]<��\<�1\<�\<�a\<��\<;�]<��^<��_<��`<��a<��b<�Dc<-�c< �c<�yc<O=c<2�b<��b<a�b<C�b<��b<9�b<V�b<�b<>�b<��b<W�b<��b<��b<�c<�Gc<݇c<m�c<t�c<�ic<%�b<{$b</a<_`<<_< ^<�(]<��\<pG\<�P\<��\<[R]<�4^<%>_<tW`<7fa<*Rb<�c<|c<(�c<��c<�{c<�9c<y�b<%�b<^�b<�b<?�b<Ūb<g�b<�b<�b<��b<��b<��b<%�b<�c<+ac<z�c<L�c<��c<�Dc<��b<��a<��`<t�_<��^<Ұ]<*�\<�n\<
@\<ge\<0�\<ŗ]<��^<n�_<c�`<�a<��b<�5c<�c<��c<q�c<mfc<"c<��b<�b<3�b<y�b<�b<(�b<��b<��b<�b<��b<ݞb<�b<5�b<s.c<Uqc<M�c<3�c<�c<�c<eb<,~a<r`<oX_<�K^<�c]<õ\<JQ\<�>\<�\<�]<m�]<��^<��_<a<�b<��b<Xc<�c<�c<j�c<�Hc<�c<�b<b�b<��b<��b<G�b<�b<|�b<I�b<T�b<Ɇb<��b<ζb<z�b<V1c<�oc<D�c<y�c<5Lc<��b<�b<�a<�_<��^<��]<�]<�j\< \<�(\<Ã\<�)]<�^<$_<1.`<�<a<B(b<K�b<JQc<ăc<}c<�Nc<=c<2�b<�b<�tb<�jb<ob<yb<Db<f|b<Rrb<�ib<�kb<|�b<�b<�b<�-c<�fc<��c<hc<�c<Lwb<�a<��`<�_<r^<{]<R�\<�8\<R
\<�/\<�\< c]<uU^<�g_<,�`<�  �  �a<��a<L�b<�
c<N1c<;(c<�c<b�b<v�b<��b<i�b<�b<v�b<c<"c<�c<O�b<��b<_�b<��b<G�b<��b<7c<Y4c<v5c<+c<��b<E�a<z�`<`�_<|�^<�]<�\<��[<!b[<@N[<��[<�2\<�]<�)^<zT_<c{`<��a<MVb<��b<t8c<�Mc<|:c<bc<9�b<��b<��b<��b<�c<0+c<Cc<�Ec<M2c<�c<��b<�b<��b<�b<Mc<�Jc<wcc<yUc<�c<��b<��a<`�`<�_<tk^<�T]<l\<��[<v[<�[<n�[<�\<��]<��^<��_<��`<}�a<��b<8"c<�[c<k`c<�Bc<Dc<(�b<��b<��b<2�b<"c<�Bc<�Rc<�Lc<.2c<&c<k�b< �b<k�b<Kc<(1c<�Wc<�dc<�Dc<��b<�Gb<hha<Y`<�/_<L	^<C�\<@+\<v�[<n[<)�[<�\<4�\<N�]<�_<8`<HKa<�0b<��b<)<c<'bc<�Xc<4c<�c<m�b<]�b<�b<�c<�+c<�Gc<@Pc<nBc</#c<��b<��b<��b<��b<�c<q:c<�Zc<�Zc<�'c<r�b<f�a<a<]�_<��^<�]<l�\<��[<��[<�l[<~�[<P\<!2]<�D^<>n_<œ`<ٙa<�kb<�b< Jc<�]c<2Hc<�c<��b< �b<��b<��b<c<=)c<�>c<�>c<Y)c<�c<W�b<;�b<��b<��b<	c<k2c<XIc<�9c<��b<Efb<�a<I�`<�r_<G^<�/]<�E\<ՠ[<�N[<PX[<E�[<�p\<�d]<��^<��_<�`<��a<=}b<X�b<v0c<K4c<�c<��b<��b<��b<�b<��b<<�b<�c<� c<c<P�b<�b<B�b<�b<"�b<��b<��b<$c<1c<�c<��b<Eb<�3a<#$`<��^<��]<��\<��[<�k[<�8[<�a[<��[<��\< �]<@�^<�`<�  �  �`<��a<�bb<��b<��b<��b<��b<L�b<-�b<��b<��b<uc<�Pc<�xc<S�c<�rc<�Fc<c<0�b<N�b<I�b<��b<�b<��b<G�b<F�b<?Lb<��a<I�`<�y_<�D^<�]<\<cO[<e�Z<��Z<[<��[<�\<+�]<��^<�)`<58a<$b<3�b<��b<�c<c<(�b<h�b<�b<�b<�c<�Pc<b�c< �c<��c<Ќc<�\c<'c<��b<s�b<a�b<��b<_c<�+c<kc<��b<�?b<hpa<�h`<�<_<^<��\<��[<�D[<��Z<�Z<Uc[<!\<[ ]<�H^<z~_<��`<e�a<�bb<��b<$c<�*c<'c<��b<��b<�b<!	c<e:c<bqc<��c<�c<e�c<l�c<�Sc<&c<��b<��b<A�b<�c<�%c<�*c<c<q�b<t b<Za<�`<
�^<�]<��\<ܭ[<�[<O�Z<[<e�[<�o\<�]<��^<��_<��`<�a<P�b<�b<e'c<&c<�c<w�b<1�b<��b<3c<�Jc<%�c<��c<��c<u�c<�sc<?=c<s
c<��b<��b<�b<Qc<�%c<�c<��b<pb<ҵa<վ`<�_<Yf^<�:]<�5\<Xo[<��Z<^�Z<1[<��[<��\<$�]<�_<B`<Oa<\%b<��b<|c<7%c<�c<��b<��b<G�b<�b<]c<�Pc<n�c<��c<^�c<݃c<wQc<�c<�b<y�b<C�b<��b</c<�c<�b<�b<� b<�Oa<�F`<<_<��]<��\<��[<&[<I�Z<J�Z<2;[<��[<��\<�^<5U_<{`<qwa<m8b<�b<��b<��b<?�b<��b<��b<ȼb<�b<�	c<
@c<�mc<��c<�zc<}Uc<� c<��b<��b<O�b<�b<,�b<\�b<�b<>�b<fpb<%�a<��`<��_<�^<�k]<.V\<?x[<8�Z<ұZ<��Z<nd[<�:\<�K]<%|^<}�_<�  �  ��`<R�a<nJb<��b<1�b<��b<��b<l�b<G�b<��b<��b<91c<�lc<ݘc<��c<	�c<�ac<=%c<��b<��b<��b<r�b<�b<V�b<q�b<��b<�3b<�xa<O�`<*[_<�"^<�\<�[<8#[<��Z<��Z<��Z<X�[<�}\<O�]<��^<�`<�a<��a<(�b<�b<c<b�b<�b<��b<��b<%�b<�)c<�hc<��c<��c<��c<�c<vuc<�8c<�c<��b<}�b<l�b<c<�c<� c<��b<�&b<�Ua<�K`<�_<��]<��\<��[<�[<��Z<5�Z<�6[<��[<�\<,&^<[__<k�`<J�a<4Jb<U�b<	c<Ac<�c<��b<��b<p�b<�c<�Mc<h�c<��c<M�c<��c<�c<`jc<h-c<7�b<��b</�b<G�b<uc<�c<��b<5�b<��a<)a<��_<�^<S|]<�c\<Ђ[<K�Z<L�Z<j�Z<�m[<(G\<�Z]<c�^<i�_<�`<\�a<|b<��b<
c<`c< �b<��b<N�b<��b<�$c<�`c<-�c<��c<��c<��c<��c<nQc<c<��b<�b<��b<f c<�c<�c<[�b<�Wb<ޛa<ܢ`<)}_<!D^<]<�\<+C[<��Z<r�Z<�[<i�[<��\<E�]<��^<�$`<[4a<0b<��b<��b<�c<c<��b<@�b<��b<�b<X,c<�hc<	�c<{�c<W�c<�c<5jc<R+c<
�b<�b<a�b<=�b<��b<��b<��b<��b<�b<=5a<�)`<s�^<V�]<��\<��[<1�Z<h�Z<u�Z<�[<>�[<d�\<0�]<6_<�^`<T]a<�b<g�b<��b<�b<��b<��b<"�b<(�b<��b<c<	Zc<��c<�c<	�c<rc<@7c<.�b<��b<G�b<յb<��b<��b<�b<�b<-Xb<��a<��`<ڲ_<�|^<�F]<1.\<;M[<��Z<փZ<,�Z<9[<�\<�&]<�Z^<Z�_<�  �  �`<��a<�bb<��b<��b<��b<��b<L�b<-�b<��b<��b<uc<�Pc<�xc<S�c<�rc<�Fc<c<0�b<N�b<I�b<��b<�b<��b<G�b<F�b<?Lb<��a<I�`<�y_<�D^<�]<\<cO[<e�Z<��Z<[<��[<�\<+�]<��^<�)`<58a<$b<3�b<��b<�c<c<(�b<h�b<�b<�b<�c<�Pc<b�c< �c<��c<Ќc<�\c<'c<��b<s�b<a�b<��b<_c<�+c<kc<��b<�?b<hpa<�h`<�<_<^<��\<��[<�D[<��Z<�Z<Uc[<!\<[ ]<�H^<z~_<��`<e�a<�bb<��b<$c<�*c<'c<��b<��b<�b<!	c<e:c<bqc<��c<�c<e�c<l�c<�Sc<&c<��b<��b<A�b<�c<�%c<�*c<c<q�b<t b<Za<�`<
�^<�]<��\<ܭ[<�[<O�Z<[<e�[<�o\<�]<��^<��_<��`<�a<P�b<�b<e'c<&c<�c<w�b<1�b<��b<3c<�Jc<%�c<��c<��c<u�c<�sc<?=c<s
c<��b<��b<�b<Qc<�%c<�c<��b<pb<ҵa<վ`<�_<Yf^<�:]<�5\<Xo[<��Z<^�Z<1[<��[<��\<$�]<�_<B`<Oa<\%b<��b<|c<7%c<�c<��b<��b<G�b<�b<]c<�Pc<n�c<��c<^�c<݃c<wQc<�c<�b<y�b<C�b<��b</c<�c<�b<�b<� b<�Oa<�F`<<_<��]<��\<��[<&[<I�Z<J�Z<2;[<��[<��\<�^<5U_<{`<qwa<m8b<�b<��b<��b<?�b<��b<��b<ȼb<�b<�	c<
@c<�mc<��c<�zc<}Uc<� c<��b<��b<O�b<�b<,�b<\�b<�b<>�b<fpb<%�a<��`<��_<�^<�k]<.V\<?x[<8�Z<ұZ<��Z<nd[<�:\<�K]<%|^<}�_<�  �  �a<��a<L�b<�
c<N1c<;(c<�c<b�b<v�b<��b<i�b<�b<v�b<c<"c<�c<O�b<��b<_�b<��b<G�b<��b<7c<Y4c<v5c<+c<��b<E�a<z�`<`�_<|�^<�]<�\<��[<!b[<@N[<��[<�2\<�]<�)^<zT_<c{`<��a<MVb<��b<t8c<�Mc<|:c<bc<9�b<��b<��b<��b<�c<0+c<Cc<�Ec<M2c<�c<��b<�b<��b<�b<Mc<�Jc<wcc<yUc<�c<��b<��a<`�`<�_<tk^<�T]<l\<��[<v[<�[<n�[<�\<��]<��^<��_<��`<}�a<��b<8"c<�[c<k`c<�Bc<Dc<(�b<��b<��b<2�b<"c<�Bc<�Rc<�Lc<.2c<&c<k�b< �b<k�b<Kc<(1c<�Wc<�dc<�Dc<��b<�Gb<hha<Y`<�/_<L	^<C�\<@+\<v�[<n[<)�[<�\<4�\<N�]<�_<8`<HKa<�0b<��b<)<c<'bc<�Xc<4c<�c<m�b<]�b<�b<�c<�+c<�Gc<@Pc<nBc</#c<��b<��b<��b<��b<�c<q:c<�Zc<�Zc<�'c<r�b<f�a<a<]�_<��^<�]<l�\<��[<��[<�l[<~�[<P\<!2]<�D^<>n_<œ`<ٙa<�kb<�b< Jc<�]c<2Hc<�c<��b< �b<��b<��b<c<=)c<�>c<�>c<Y)c<�c<W�b<;�b<��b<��b<	c<k2c<XIc<�9c<��b<Efb<�a<I�`<�r_<G^<�/]<�E\<ՠ[<�N[<PX[<E�[<�p\<�d]<��^<��_<�`<��a<=}b<X�b<v0c<K4c<�c<��b<��b<��b<�b<��b<<�b<�c<� c<c<P�b<�b<B�b<�b<"�b<��b<��b<$c<1c<�c<��b<Eb<�3a<#$`<��^<��]<��\<��[<�k[<�8[<�a[<��[<��\< �]<@�^<�`<�  �  7�a<rcb<>c<�bc<ׁc<�lc<$6c<�b<��b<+�b<�mb<4jb<+rb<�|b<��b<Q{b<]qb<�kb<�sb<�b<�b<[c<7Jc<!|c<�c<u\c< �b<�Ab<�[a<P`<�6_<�*^<WC]<��\<�1\<�\<�a\<��\<;�]<��^<��_<��`<��a<��b<�Dc<-�c< �c<�yc<O=c<2�b<��b<a�b<C�b<��b<9�b<V�b<�b<>�b<��b<W�b<��b<��b<�c<�Gc<݇c<m�c<t�c<�ic<%�b<{$b</a<_`<<_< ^<�(]<��\<pG\<�P\<��\<[R]<�4^<%>_<tW`<7fa<*Rb<�c<|c<(�c<��c<�{c<�9c<y�b<%�b<^�b<�b<?�b<Ūb<g�b<�b<�b<��b<��b<��b<%�b<�c<+ac<z�c<L�c<��c<�Dc<��b<��a<��`<t�_<��^<Ұ]<*�\<�n\<
@\<ge\<0�\<ŗ]<��^<n�_<c�`<�a<��b<�5c<�c<��c<q�c<mfc<"c<��b<�b<3�b<y�b<�b<(�b<��b<��b<�b<��b<ݞb<�b<5�b<s.c<Uqc<M�c<3�c<�c<�c<eb<,~a<r`<oX_<�K^<�c]<õ\<JQ\<�>\<�\<�]<m�]<��^<��_<a<�b<��b<Xc<�c<�c<j�c<�Hc<�c<�b<b�b<��b<��b<G�b<�b<|�b<I�b<T�b<Ɇb<��b<ζb<z�b<V1c<�oc<D�c<y�c<5Lc<��b<�b<�a<�_<��^<��]<�]<�j\< \<�(\<Ã\<�)]<�^<$_<1.`<�<a<B(b<K�b<JQc<ăc<}c<�Nc<=c<2�b<�b<�tb<�jb<ob<yb<Db<f|b<Rrb<�ib<�kb<|�b<�b<�b<�-c<�fc<��c<hc<�c<Lwb<�a<��`<�_<r^<{]<R�\<�8\<R
\<�/\<�\< c]<uU^<�g_<,�`<�  �  b<��b<�fc<޼c<P�c<��c<�ac<��b<��b<�Ab<�a<"�a<��a<��a<C�a<�a<˺a<z�a<?b<]Wb<��b<c<6{c<��c<��c<i�c<�Tc<رb<d�a<��`<��_<��^<�'^<x�]<�8]<)]<Qb]<K�]<q�^<�~_<|`<�za<"db<�!c<l�c<��c<:�c<j�c<�_c<��b<q�b<�Hb<�b<��a<�a<v�a<O�a<,�a< �a<�b<�Kb<��b<* c<�fc<W�c<�c<% d<��c<:Oc<�b<A�a<ڸ`<]�_<X�^<R^<�]<NP]<X]<��]<d9^<�_<�_<�`<��a<t�b<Qmc<��c<Pd<��c<(�c<LRc<_�b<,�b<�Bb<b<�a<}�a<F�a<Q�a<��a<4�a<�(b<"kb<�b<�&c<ۉc<��c<fd<�c<�c<�c<�Ob<�`a<�a`<�h_<�^<��]<cr]<�I]<0j]<��]<�v^<	N_<xD`<Da<�5b<�c<��c<�c<(d<x�c<�c<�/c<e�b<Pqb<q,b<@�a<��a<�a<�a<Q�a<S�a<3b<8b<B�b<��b<oCc<.�c<��c<�c<��c<dxc<��b<��a<�a<``<�_<*H^<��]<X]<�G]<s�]<��]<��^<�_<�`<��a<${b<B7c<�c<��c<�c<3�c<�kc<^c<��b<�Mb<bb<X�a<�a<.�a<��a<6�a<��a<Nb<*<b<��b<��b<�Pc<�c<��c<�c<&�c<�/c<8xb<	�a<j�`<ؖ_<�^<�]<�i]<�(]<.0]<o]<�^<�^<�_<��`<m�a<��b<Cc<9�c<�c<��c<��c<�$c<?�b<G_b<�b<��a<�a<��a<K�a<��a<��a<]�a<��a<8b<�b<A�b<vVc<	�c<��c<�c<�rc<�b<�b<�+a<,`<%3_<�V^<��]<]<]<�]<�4]<��]<�A^<�_<�`<�a<�  �  Otb<^-c<ʵc<>d<�
d<��c<"tc<}�b<eb<�a<�ga<�a<��`<§`<>�`<<�`<�`<�a<T�a<x�a<Јb<
c<h�c<��c<d<��c<?�c<�c<,Rb<�xa<ԛ`<	�_<y#_<>�^<'_^<�R^<��^<8�^<)�_<�D`<�a<��a<��b<}yc<z�c<�%d<6d<H�c<�hc<�b<�Ub<��a<6ga<�a<D�`<��`<��`<��`<ma<5ea<\�a<�Sb<��b<Zlc<��c<u,d<@d<�d<M�c<� c<�4b<�Wa<t}`<[�_<7_<S�^<�y^<�^<��^<�8_<��_<�`<r�a<�ab<]&c<6�c<} d<�?d<ed<�c<`Pc<��b<t9b<ϼa<�Wa<�a<��`<`�`<t�`<��`<�4a<؍a<� b<��b<5c<3�c<d<�:d<k8d<��c<�rc<��b<��a<�a<7`<=~_<��^<2�^<Ft^<~�^<��^<�k_<D `<��`<��a<,�b<�_c<��c<�2d<�;d< d<P�c<i"c<��b<�b<��a<�:a<~�`<��`<��`<B�`<_a<Ka<�a<''b<��b<�=c<4�c<|d<;d<7#d<��c<�5c<�tb<��a<T�`<�_<D_<c�^<�~^<�q^<ş^<�_<��_<�_`<�8a<Sb<�b<�c<+d<�7d<+d<�c<Ytc<��b<]b<��a<�ia<a<W�`<��`<=�`<��`<$	a<�Wa<��a<�Ab<��b<Vc<n�c<5d<�#d<�c<ۅc<��b<�b<%4a<�X`<Γ_<��^<O�^<�Q^<�W^<��^<_<�_<	�`<1]a<8b<��b<�c<��c<cd<��c<��c<.#c<�b<�
b<]�a<�'a<9�`<n�`<��`<F�`<}�`<a<�Za<��a<gTb<��b<�ec<��c<�d<`d<,�c<>c<��b<%�a<9�`<,`<H_<��^<�^^<'>^<�X^<1�^<y6_<��_<��`<��a<�  �  ��b<Ahc<��c<�d<d<p�c<jac<��b<jb<�Va<�`<�'`<��_<d�_<av_<��_<<�_<JE`<��`<��a<�9b<��b<L�c<�c<�)d<�d<��c<zRc<�b<v�a<�Da<�`<� `<�_<��_<υ_<��_<��_<�j`<@a<&�a<�hb<�c<��c<�d<�>d<A(d<��c<~Lc<T�b<Y�a<7=a<�`< $`<��_</�_<�_<D�_<s`<ߙ`<}5a<g�a<�b<�Lc<�c<�7d<�Wd<�5d<��c<�Hc<'�b<��a<&5a<U�`<$`<@�_<<�_<װ_<��_<�9`<��`<�Wa<�
b<��b<�hc<��c<�@d<�Td<a'd<O�c<�)c<�yb<��a<a<U�`<�`<(�_<��_<<�_<��_<L`<�`< ua<�)b<��b<u�c<�d<�Jd<�Sd<3d<t�c<�c<�]b<�a<��`<�n`<r`<��_<	�_<��_<��_<p``<��`<X�a<KHb<��b<��c<�d<�Nd<�Ld<�
d<��c<��b<�;b<	�a<&�`<]V`<`�_<V�_<ˣ_<r�_<L`<�p`<� a<(�a<bb<Vc<�c<�d<�Nd<Bd<P�c<buc<F�b<db<efa<��`<3A`<H�_<��_<ݤ_<
�_<"`<�`<�a<B�a<��b<�/c<:�c<�'d<�Pd<18d<��c<CXc<�b<��a<JBa<ǣ`<n$`<��_<�_<R�_<K�_<'`<G�`<�%a<S�a<ϋb<�6c<��c<�d<�;d<d<	�c<�'c<�yb<6�a<qa<�v`<��_<#�_<��_<ň_<2�_</`<��`<�.a<C�a<~�b<�>c<d�c<d<�)d<��c<��c<��b</Lb<)�a<��`<fR`<"�_<�_<v_<<�_<8�_<u`<D�`<5Ba<��a<e�b<Pc<]�c<�d<�d<��c<�vc<��b<5(b<qa<w�`<k8`<��_<%�_<�q_<��_<��_<+`<Ѷ`<!^a<�b<�  �  ��b<�yc<A�c<�d<�c<j�c<W%c<�jb<$�a<ϴ`<��_<�0_<��^<�Y^<�B^<kg^<��^<-W_<�`<9�`<��a<M�b<�Nc<D�c<Vd<�d<�c<�ic<q�b<kXb<O�a<:ba<}a<��`<Ǳ`<�`<��`<��`<�=a<�a<,$b<R�b<�=c<�c<�
d<)d<Pd<��c<�c<�Bb<ha<�`<�_<� _<Ĭ^<�o^<�m^<��^<�_<S�_<_�`<�\a<�:b<yc<��c<�d<�@d<g+d<��c<�ic<Y�b<�Sb<��a<Vja<Ja<�`<��`<�`<��`<^)a</}a<��a<eob<��b<�c<��c<�2d<;d<d<�c<�b<�b<�.a<�V`<p�_<C_<��^<=t^<�^<�^<�P_<w�_<]�`<^�a<��b<�Dc<I�c<?,d<�@d<�d<�c<8<c<�b<�%b<\�a<�Ka<Xa<v�`<;�`<^�`<a<?Ba<��a<6b<��b<�+c<��c<d<=d<�/d<��c<gUc<C�b<��a<��`<f`<j__<��^<h�^<p^<��^<[�^<2�_<�<`<sa<��a<��b<Muc<��c<4d<�2d<n�c<��c<�c<Wzb<��a<\�a<7,a<?�`<��`<3�`<_�`<ca<Za<��a<c>b<"�b<�Tc<��c<�d<�:d<Pd<��c<�c<�Lb<ooa<�`<��_<d!_<۪^<lk^<g^<��^<B_<��_<~p`<�Ja<�&b<�b<��c<U�c<�$d<pd<�c<�Hc<ݽb<)0b<��a<�Da<��`<��`<�`<�`<6�`<� a<ITa<��a<%Fb<�b<dYc<��c<Hd<d<}�c<�]c<8�b<"�a<C a<�'`<�h_<��^<�m^<�B^<S^<��^<z_<��_<��`<^ya<�Rb<�c<��c<[�c<Md</�c<�c<�c<�yb<x�a<�ua</a<��`<��`<��`<�`<�`<�a<�ja<��a<�jb<�  �  �c<�ec<��c<��c<�c<�`c<��b<��a<�a<�`<m_<M:^<͗]<�4]<�]<�E]<'�]<�g^<�F_<A`<�@a<�.b<��b<a�c<��c<T�c<��c<\c<��b<q�b<)@b<��a<�a<�a<D�a<��a<P�a<��a<��a<�'b<vb<U�b<�=c<��c<[�c<��c<!�c<�Pc<��b<��a<��`<�_<�^<	 ^<��]<�G]<�D]<W�]<b^<]�^<i�_<ʿ`<�a</�b<�Tc<s�c<�d<�c<��c<wfc<� c<��b<LQb<�b<�a<	�a<��a<�a<��a<x�a<	 b<*^b<��b<.c<�xc<��c<��c<Q�c<7�c<Q1c<�qb<0�a<��`<��_<��^<��]<j~]<0J]<�^]<\�]<�V^<;'_<T`<4a<Kb<�b<��c<S�c<.d<�c<l�c<�Cc<��b<R�b<&:b<Xb<0�a<��a<��a<��a<��a<�b<�2b<Qxb<��b<7c<-�c<s�c<�d<��c<^�c<��b<�'b<�3a<�3`<+>_<�h^<��]<lb]<�E]<�q]<��]<��^<�p_<j`<�ha<�Ub<c<̦c<5�c<D�c<��c<�~c<$c<Y�b<�ab<� b<��a<k�a<�a<��a<��a<R�a<�b<�Cb<V�b<=�b<�Tc<M�c<G�c<�c<0�c<�^c<��b<��a<C�`<!�_<��^< ^<��]<fC]<9>]<\�]<^<��^<��_<��`<��a<ĉb<S<c<
�c<X�c<��c<ןc<HEc<\�b<�|b<e,b<��a<r�a<��a<ݱa<رa<r�a<��a<�a<5b<B�b<��b<�Nc<��c<z�c<y�c<Ҋc<Mc</Eb<�Za<�[`<�__<"}^<t�]<�M]<�]<-]<[�]<Z$^<��^<��_<C�`<&�a<��b<�Qc<a�c<��c<j�c<Tnc<:c<�b<
Lb<�b<��a<C�a<��a<¡a<�a<^�a<��a<��a<�Cb<�b<�  �  N�b<�8c<�nc<y�c<�_c<��b<�Yb<%{a<�s`<sZ_<�I^<1Z]<&�\<�/\<6\<�B\<��\<d�]<�^<z�_<�`<�a<��b<
 c<)tc<�c<�nc<�4c<�b<ƴb<�b<�wb<~wb<��b<d�b<M�b<@�b<�~b<n{b<�b<l�b<�b<#c<�ec<�c<�c<�ac<��b<�2b<Ea<�5`<�_<O^<�7]<�\<�?\<Y<\<�\<l(]<�^<�	_<�#`<�7a<�,b<e�b<nc<��c<=�c<S�c<�Hc<�c<(�b<�b<��b<��b<��b<�b<{�b<ǧb<�b<1�b<$�b<��b<nc<lTc<��c<�c<�c<�Uc<U�b<��a<��`< �_<��^<��]<]<�|\<�@\<TX\<��\<�s]<u^^<�l_<��`<��a<�ub<M!c<�c<ٳc<a�c<�sc<�0c<��b<��b<j�b<�b<��b<�b<�b<ڮb<Z�b<��b<�b<t�b<#�b<�'c<Kkc<��c<۲c<|�c<.c<ŉb<��a<�`<d�_<dx^<p�]<��\<]\<�;\<o\<D�\<��]<ΰ^<Q�_<��`<��a<ïb<TEc<��c<ܭc<ّc<�Wc<Xc<��b<��b<�b<P�b<W�b<M�b<��b<ܦb<��b<9�b<Ţb<��b<�b<�:c<�{c<�c<6�c<�qc<��b<�>b<�Na<F=`<�"_<!^<+8]<�\<�;\<�5\<�\<]<�]<��^<�`<�#a<b<��b<�Sc<E�c<'�c<�hc<�'c<��b<E�b<��b<�xb<�zb<)�b<�b</�b<0b<Lub<9tb<�b<G�b<�b<�*c<�fc<��c<(wc<q*c<p�b<�a<H�`<&�_<I�^<t�]<~�\<CL\<�\<�&\<��\<yA]<,^<1:_<�S`<o^a<�Bb<��b<�Vc<|c<�qc<�>c<��b<��b<'�b<�lb<fb<�lb<�vb<|b<xb<�mb<�fb<�kb<Ʉb<&�b<�  �  �b<c<)c<q0c<ac<s�b<z�a<�a<��_<
�^<^�]<��\<�[<6a[<q=[<,v[<�\<�\<��]<_<H;`<AIa<
&b<�b<Sc<	;c<�,c<c<�b<�b<��b<��b<��b<Cc<�)c<|/c<6c<��b<��b<��b<�b<��b<�b<�+c<3Ic<gCc<ic<�b<h�a<��`<`�_<��^<dn]<z}\<��[<(o[<9k[<��[<ll\<�Y]<Ds^<��_<�`<I�a<A�b<$c<Xc<ec<-Lc<�!c<��b<��b<�b<-�b<c<�@c<�Sc<�Pc<�8c<�c<��b<��b<��b<��b<)(c<vPc<cc<�Kc<]�b<ydb<�a<W�`<�__<�6^<i&]<�G\<�[<�n[<�[<��[< �\<ɺ]<^�^<�`<!a<�b<R�b<2c<�ac<k_c<>c<tc<��b<6�b<&�b<�c<$*c<�Hc<�Tc<�Jc<|-c<�	c<��b<��b<��b<~c<�7c<[c<�ac<<8c<��b<i$b<�;a<�%`<��^<��]<��\<�
\<m�[<j[<+�[<#0\<y]<�^<�:_<c`<$pa<Lb<O�b<�Ac<�^c<�Oc<�(c<b�b<��b<�b<��b<uc<�/c<�Ic<�Nc<�=c<ic<|�b<G�b<��b<��b<�c<pAc<<]c<�Uc<�c<.�b<U�a<p�`<׺_<�^<:q]<�}\<��[<�j[<�d[<��[<a\<�K]<Vc^<m�_<��`<Ьa<�sb<��b<�;c<�Fc<f,c<� c<,�b<�b< �b</�b<��b<:c<�+c<n(c<c<��b<��b<}�b<@�b<[�b<��b<�&c<�8c<!c<(�b<�8b<�ba<2Y`<�1_<T^<+�\<\<��[<�=[<zW[<*�[<�\<k�]<��^<�_<��`<`�a<��b<��b<-c<�*c<�c<��b<��b<��b<@�b<��b<��b<Bc<�c<�c<��b<��b<T�b<0�b<ɷb<�  �  �b<�b<��b<R�b<�b<�[b<��a<��`<ȡ_<?m^<C>]<�0\<\^[<�Z<öZ<��Z<�[<%j\<l�]<�^<?�_<��`<&�a<#�b<��b<gc<r�b<H�b<�b<W�b<��b<��b<Q1c<=fc<��c<w�c<�{c<oMc<�c<U�b<��b<��b<f�b<R�b<�c<Cc<��b<Eb<�a<L�`<d[_<�&^<j ]<�\<SL[<�Z<��Z<_@[<��[<^�\<�^<�F_<�r`<aya<�Fb<U�b<fc<�-c<�c<uc<R�b<.�b<Ec<�4c<vkc<כc<n�c<��c<1�c<y]c<l&c<�b<|�b<��b<c<n c</*c<�c<��b<b<�Ca<$4`<�_<��]<��\<�[<?-[<%�Z<>[<(|[<�F\<UO]<S|^<�_<<�`<g�a<)~b<W�b<&c<9+c<�c<��b<�b<b�b<bc<�Ec<�{c<�c<;�c<5�c<&�c<>Kc<�c<��b<p�b<z�b<�c<�'c<�&c<��b<�b<��a<x�`<��_<�^<�l]<�^\<��[<)	[<R�Z<�[<<�[<��\<�]<��^<�`<c$a<b<E�b<Mc<#%c<�c<�c<\�b<9�b<G�b<�c<1Rc<��c<��c<�c<<�c<Pkc<m4c<c<V�b<��b<��b<-c<'c<mc<�b<*Sb<��a<�`<�b_<�+^<A]<m\<rJ[<��Z<<�Z<a7[<d�[<��\<��]<m4_<i^`<�ba<@.b<Ҷb<�b<�c<��b<�b<��b<2�b</�b<�c<�Dc<\tc<p�c<!�c<�hc<�4c<j�b<^�b<<�b<u�b<t�b<��b<��b<(�b<��b<D�a<�a<`<��^<�]<z�\<E�[<��Z<A�Z<��Z<qJ[<�\<]<�I^<_<%�`<�a<wJb<I�b<��b<T�b<M�b<��b<ϲb<��b<g�b<mc<zDc<�oc< �c<<sc<�Jc<(c<�b<��b<M�b<�  �  �b<[�b<(�b<��b<)hb<�b<X{a<�`<��_<�_<2^<n]<��\<Vw\<�\\<Y�\<l�\<p�]<�d^<�E_<.'`<��`<��a<�(b<)b<t�b<^�b<��b<"�b</�b<��b<)�b<��b<�b<��b<��b<��b<2�b<��b<)�b<]�b<��b<�b<{�b<y�b<��b<=hb<F�a<�_a<��`<��_<��^<_^<W]<O�\<��\<G�\<��\<_K]<L�]<`�^<Z�_<?�`<1]a<s�a<�sb<��b<�b<��b<��b<��b<q�b<)�b<��b<
�b< c<�c<�c<c<D�b<��b<9�b<��b<�b<��b<M�b<��b<�b<]b<��a<�5a<j`<u�_<�^<L�]<�1]<v�\<��\<<�\<��\<ϊ]<K^<'_<!
`<�`<��a<�,b<��b<��b<��b<��b<a�b<Y�b<�b<��b<��b<c<�c<�c<3c<'c<��b<��b<��b<��b<��b<J�b<~�b<��b<i�b<]8b<��a<��`<l `<�=_<�_^<h�]<�]<��\<z�\<{�\<�]<�]<��^<�m_<dN`<�a<�a<zMb<7�b<��b<'�b<��b<��b<x�b<Z�b<��b<��b<�c<fc<�c<[c<��b<�b<��b<��b<V�b<>�b<*�b<q�b<ºb<~wb<�b<�ja<��`<��_<��^<�^<kW]<c�\<΅\<ր\<��\<s@]<+�]<�^<�_<��`<�Ga<��a<-Zb<x�b<-�b<��b<��b<S�b<��b<��b<�b<��b<�b<8�b<��b<��b<y�b<��b<�b<V�b<Y�b<�b<�b<٬b<σb<X2b<Y�a<�	a<�=`<G]_<A{^<۫]<�]<�\<�\\<�o\<��\<�Y]<�^<N�^<�_<��`<�ga<�a<�^b<ߗb<��b<q�b<��b<;�b<��b<ӟb<��b< �b<�b<��b<��b<��b<��b<Y�b<�b<d�b<�  �  ��b< �b<��b<ƨb<�ub<�b<g�a<��`<�`<+'_<�L^<��]<��\<ї\<q}\<��\<�]<�]<�~^<�\_<�;`<�a<"�a<�7b<��b<��b<m�b<��b<��b<֝b<Ȝb<��b<T�b<Q�b<��b<~�b<��b<�b<´b<K�b<��b<ϭb<��b<X�b<��b<5�b<�vb<2
b<nqa<<�`<��_<?�^<�(^<�t]<�\<��\<�\<s�\< i]<�^<4�^<�_</�`<oa<�b<�b<f�b<x�b</�b<[�b<U�b<Q�b<��b<G�b<Z�b<t�b<�c<c<��b<��b<��b<��b<��b<�b<d�b<�b<��b<7�b<�kb<�a<�Ga<�~`<0�_<��^<��]<P]<��\<~�\<��\<�]<�]<�e^<�>_<p`<�`<�a<�<b<�b<��b<J�b<��b<v�b<��b<�b<|�b<��b<2�b<��b<_c<��b<��b<9�b<�b<0�b<C�b<7�b<�b<�b<��b<=�b<�Gb<��a<�a<�5`<QU_<`z^<P�]<�!]</�\<=�\<��\<e=]<��]<k�^<��_<	c`<a/a<��a<\b<��b<�b<8�b<��b<a�b<�b<��b<��b<D�b<��b<��b<��b<j�b<��b<M�b<��b<ѽb<��b<G�b<�b<��b<Z�b<�b<xb<�|a<]�`<��_<
_<J+^<�t]<�\<a�\<z�\<��\<4^]<�^<��^<�_<��`<�Ya<�a<�hb<B�b<��b<��b<y�b<�b<ޡb<?�b<ǯb<�b<n�b<1�b<�b<u�b<��b<��b<��b<i�b<I�b<U�b<��b<ڷb<��b<-Ab<��a<�a<�Q`<�s_<ה^<�]<� ]< �\<i}\<?�\<�\<�v]<^4^<+_<Y�_<��`<Eya<�	b<�lb<��b<L�b<��b<��b<w�b<��b<ӓb<֣b<D�b<��b<��b<0�b<��b<k�b<ѕb<q�b<�b<�  �  Φb<��b<l�b<n�b<�b<eBb<�a<�a<�B`<�j_<��^<��]<O]<��\<�\<�]<�k]<^<{�^<Y�_<v`<�<a<f�a< ab<s�b<��b<b�b<��b<�b<��b<;�b<6~b<��b<�b<��b<ܗb<m�b<S�b<�b<�b<��b<S�b<"�b<F�b<��b<��b<�b<#6b<��a<d�`<�`<zB_<{w^<��]<LM]<�	]<q]<;F]<��]<�j^<^5_<�`<�`<�a<�:b<��b<��b<hc<%�b<��b<M�b<�b<"�b<�b<��b<��b<R�b<T�b<²b<d�b<��b<��b<�b<��b<\�b< c<( c<��b<ޔb<�b<�za<�`<�_<�_< H^<e�]<v<]<;]<�]<r]<��]<в^<]�_<(\`<�)a<��a<zgb<i�b<��b<�c<��b<��b<�b<��b<�b<�b<�b<ݷb<��b<w�b<��b<-�b<�b<�b<3�b<N�b<��b<�c<0�b<-�b<,rb<E�a<�<a<kq`<ʘ_<W�^<3^<�{]<�"]<�]<�0]<�]<�0^<u�^<}�_<j�`<!ca<	b<��b<��b<V�b<4�b<�b<��b<ܳb<�b<��b<s�b<��b<u�b<�b<Ұb<קb<��b<l�b<�b<�b<d�b<��b<��b<��b<B�b<eCb<�a<��`<� `<BG_<z^<�]<_K]<�]< ]<�=]<�]<v]^<&_<-�_<��`<e�a<�#b<��b<t�b<��b<��b<��b<�b<��b<��b<��b<g�b<��b<��b<E�b<N�b<��b<�{b<c~b<��b<,�b<J�b<��b<Y�b<M�b<jb<b�a<Oa<}�`<ʹ_<��^<z^<Iy]<�]<�\<1�\<A]<F�]<=�^<�Q_<*`<u�`<Z�a<�4b<(�b<R�b<��b<M�b<1�b<�b<Uxb<Uob<Jqb<0yb<�b<҅b<��b<�zb<orb<�ob<mwb<�b<�  �  �b<X�b<��b<.�b<��b<~b<	 b<R[a<��`<��_<s_<-`^<`�]<�]<�r]<ԗ]<1�]<��^<\9_<�`<6�`<ׇa<�%b<�b<��b<� c< �b<��b<�b<{b<�Sb<t8b</)b<�"b< "b<�"b<T$b<8)b<�5b<�Lb<qb<+�b<��b<��b<8c<jc<��b<�tb<��a<O;a<w`<<�_<�^<9P^<X�]<��]<y�]<�]<�F^<��^<��_<Km`<:5a<��a<^zb<c�b<c<�*c<Dc<+�b<r�b<ܔb<�pb<Yb<`Lb<�Gb<eFb<;Fb<#Gb<�Lb<`[b<�ub<��b<��b<��b<bc<�(c<�c<�b<,^b<,�a<�a<�C`<?{_<+�^<�1^<��]<¢]<̳]<s�]<k^<`(_<�_<�`<fxa<!b< �b<6�b<�%c<�(c<�c<+�b<�b<ˆb<�fb<Sb<nIb<�Fb<Fb<RFb<uHb<Qb<$cb<��b<��b<��b<2c<@%c<�%c<# c<٭b<g/b<M�a<\�`<�_<T:_<��^<h^<s�]<��]<+�]<� ^<��^<qb_<�)`<��`<a�a<dKb<��b<�c<-$c<�c<:�b<��b<Q�b<�tb<�Xb<Ib<?Bb<�@b<�@b<�Ab<�Eb<,Qb<Ugb<#�b<�b<��b<yc<$c<�c<��b<ǁb<��a<hDa<~`<�_<��^<�P^<i�]<z�]<�]<d�]<�;^<��^<i�_<�[`<�!a<r�a<�bb<�b<��b<$c<��b<Z�b<I�b<{rb<.Mb<�4b< 'b<�!b<�b<6b<�b<=%b<Z3b<9Mb<osb<�b<��b<��b<�b<��b<7�b<�2b<!�a<;�`<�`<AM_<��^<k^</�]<�r]<%�]<m�]<N^<��^<2�_<]�`<Fa<a�a<qb<��b<
�b<��b<��b<��b<�|b<�Qb<%1b<pb<�b<�b<jb<�b<eb<ab<�.b<Nb<�xb<�  �  àb<�b<Rc<�c<`c<ֽb<�Jb<��a<Oa<EL`<r�_<�_<��^<�D^<�0^<:Q^<e�^<i#_<�_<�x`<�0a<�a<�mb<u�b<�c<�(c<c<i�b<1�b<�Rb<�b<Z�a<9�a<f�a<��a<.�a<N�a<��a<��a<��a<<b<�b<��b<�c<T3c<�5c<hc<ڷb<�8b<�a<��`<8/`<p�_<��^<��^<�[^<�Y^<y�^<��^<"|_<�%`<�`<��a<�9b<Ծb<Cc<�Jc<yNc<�-c<��b<�b<�bb<�!b<��a<��a<�a<$�a<��a<͵a<c�a<&�a<"-b<apb<-�b<��b<�5c<zOc<Cc<Y
c<<�b<�b<�oa<��`<�`<�`_<d�^<��^<�`^<�o^<$�^<7#_<��_<�h`<!a<}�a<Vmb<��b<�1c<UQc<~Gc<�c<O�b<��b<<Kb<�b<�a<{�a<�a<�a<��a<��a<G�a<Fb<�Bb<Q�b<#�b<�c<�Bc<cPc<�5c<��b<Vzb<��a<�2a<�z`<l�_<�/_<��^<�q^<�\^<�|^<.�^<pM_<G�_<�`<tXa<�b<��b<x�b<!;c<Lc<6c<�c<��b<�sb<l/b<��a<�a<��a<l�a<>�a<��a<��a<�a<Ab<	Ub<��b<��b<"c<.Fc<�Fc<�c<�b< Db<��a<��`<�3`<��_<�^<��^<jW^<nS^<˃^<�^<o_<�`<��`<�a<$b<k�b<�c<|/c<�1c<�c<��b<��b<�@b<g�a<a�a<��a<�a<��a<�a<m�a<��a<&�a<�b<�Gb<_�b<��b<4c<�%c<�c<l�b<�yb<��a<Ca<��`<��_<?2_<�^<�V^<�0^<�>^<�^<��^<�_<�6`<��`<�a<�:b<�b<��b<�c<�c<j�b<ʧb<�]b<b<��a<��a<߉a<Zxa<�ra<Twa<��a<��a<:�a<nb<]Vb<�  �  څb<R�b<# c<�<c</c<��b<Ɏb<	b<�na<u�`<�6`<Ŵ_<�R_<+_<�_<�!_<�f_<T�_<�Y`<P�`<T�a<<.b<^�b<�c<�=c<�Bc<<c<��b<�{b<�b<ױa<�Ya<�a<��`<��`<��`<��`<� a<#>a<�a<!�a<"Yb<�b<�c<EGc<)Wc<;c<��b<�b<��a<�Wa<ݹ`<)`<~�_<�\_<0_<�._<Y_< �_<e"`<;�`<�Ra<��a<��b<g�b<RJc<Wmc<dc<�2c<��b<T�b<�b<7�a<aga<l(a<��`<%�`<E�`<Qa<:3a<eva<��a< 0b<��b<
�b<�>c<Thc<�hc<F<c<&�b<2hb<�a<3a<�`<�`<͞_<�U_<�6_<�B_<z_<��_<�W`<��`<��a<*b<�b<c<�\c<�oc<�Wc<c<�b<__b<�a<֛a<IOa<�a<g�`<�`<��`<Qa<�Ga<��a<E�a<�Rb<$�b<c<VQc<�mc<L_c<w#c<:�b<#8b<e�a<��`<�d`<}�_<�_<�C_<�2_<9M_<��_<��_<<�`<�a< �a<	Ub<P�b<�0c<5bc<�fc<7Ac<A�b<c�b<�6b<��a<Vza<�4a<=a<��`<��`<��`<�a<uYa<&�a<
b<�pb<$�b<%c<Zc<)hc<<Jc<�b<1�b<��a<�^a<��`<�+`<˱_<�Z_<�+_<g(_<ZP_<�_<N`<��`<8Aa<S�a</ob<�b<1c<URc<SGc<�c<��b<Iab<?�a<�a<Ca<Na<�`<��`<Z�`<��`<�a<kNa<��a<xb<�mb<��b<ec<[>c<N>c<Ac<��b<�;b<�a<ta<�h`<��_<To_<�%_<%_<�_<�H_<��_<�%`<�`<�[a<��a<M�b<=�b<�)c<�<c<<$c<��b<��b<�*b<!�a<�fa<�a<�`<��`<˳`<��`<��`<#a<�]a<߹a< b<�  �  �Tb<N�b<Kc<�Cc<�Bc<Nc<��b<�Ob<<�a<4Ja<�`<zi`<�`<_�_<��_<j�_<R-`<Z�`<��`<�ja<��a<�ob<��b<�)c<�Nc<�Fc<�c<+�b<�Db<��a<@a<�`< g`<� `<$�_<��_<'`<�G`<��`<a<��a<Wb<>�b<��b<�Dc<fbc<4Sc<�c<l�b<HCb<��a<t?a<��`<rn`<l-`<�`<#`<}+`<~k`<j�`<<a<��a<�Cb<2�b<#c<�cc<�yc<�bc<X!c<Q�b<�Bb<L�a<�=a<U�`<r`<�4`<3`<�`<�>`<l�`<$�`<qWa<��a<�\b<��b<�1c<�jc<Oxc<%Yc<�c<v�b<�)b<l�a<�&a<׸`<Tc`<�+`<�`<,`<CG`<)�`<a�`<�la<��a<sb<�b<w?c<�qc<*xc<�Qc<c<��b<b<��a<�a<t�`<�Y`<�&`<4`<�"`<R`<��`<ga<K�a<ib<�b<��b<sIc<otc<�rc<&Ec<Q�b<�~b<�a<�xa<H�`<V�`<K`<[`<$`<>$`<tX`<��`<5a<`�a<�b<��b<�c<<Oc<+sc<[jc<�5c<��b<�fb<�a<�`a<l�`<͆`<�?`<�`<r`<K*`<�c`<�`<2*a<|�a<�-b<D�b<mc<WWc<Xsc<Ebc<�%c<��b<KLb<k�a<+Da<w�`<�n`<y+`<�`<�`<�"`<�``<V�`<�,a<(�a<�0b<ɩb<�c<�Jc<�^c<KFc<'c<��b<�!b<�a<ya<�`<�L`<`<��_<��_<�`<�Z`<1�`<3/a</�a< 4b<��b<�c<�@c<�Mc<.c<��b<{b<��a<�wa<U�`<͉`<�3`<o�_<#�_<'�_<�`<�^`<��`<�:a<h�a<�@b<a�b<�c<�>c<�Dc<'c<%�b<nab<��a<�\a<��`<Au`<B$`<��_<�_<�_<i`<Tk`<��`<Oa<��a<�  �  �b<A�b<t�b<�0c<�<c<
c<��b<�b<1b<ɶa<�[a<�a<��`<��`<`�`</�`<��`<i#a<�qa<V�a<�7b<��b<3�b<1/c<�Ec<�0c<{�b<�b<k�a<^a<Y�`<�*`<�_<�R_<}_<�_<[8_<��_<=�_<*�`<�a<��a<AVb<��b<�(c<�Sc<�Qc<J'c<��b<y~b<�b<��a<�aa<� a<��`<��`<��`<��`<x a<�aa<��a<�b<�b<�b<p3c<dc<�lc<wHc<��b<��b<��a<�Pa<�`<�$`<0�_<la_<�:_<-?_<�n_<��_<�@`<z�`<xra<�b<��b<�c<VSc<�mc<�\c<?%c<��b<}nb<�b<�a<�Xa<�a<�`<a�`<��`<�
a<�<a<��a<�a<�Ab<h�b<�c<Jc<Cmc<�fc<�2c<��b<�Rb<Ӻa<xa<a�`<��_<��_< O_<�6_<J_<�_<�_<�o`<a<3�a<�Ab<��b<�(c<rac<�lc<�Mc<�c<)�b<!Kb<o�a<?�a<�@a<ma<��`<��`<1�`<Ca<�Ma<e�a<8�a<�_b<��b<lc<�Tc<Fjc<�Tc<�c<��b<Pb<�a<+�`<9K`<��_<�q_<=_<�3_<lU_<��_<g`<4�`<�8a<`�a<5lb<��b<Q;c<�dc<�`c<\4c<��b<t�b<db<@�a<\da<� a<��`<��`<H�`<��`<�a<�Ta<��a<�b<�nb<��b<"c<�Jc<�Qc<�+c<��b<�ab<��a<�.a<�`<� `<8�_<�;_<P_<b_<�G_<*�_<�`<?�`<�Ia<�a<~sb<��b<8)c<CCc<�1c<b�b<3�b<GAb<��a<�ya<�)a<��`<��`<��`<u�`<C�`<�
a<�Qa<��a<�b<�ub<��b<-c<3:c<:3c<��b<
�b<�b<c�a<��`<~K`<��_<x\_<_<�_<X_<tS_<	�_<�;`<��`<�ua<�  �  Y�a<BQb<P�b<�c< c<c<��b<B�b<+Tb<"b<�a<�a<�a<�za<wa<�}a<��a<��a<��a<� b<ib<O�b<��b<�c<K&c<c<��b<�=b<֡a<b�`<�8`<u�_<��^<؉^<K^<&@^<�i^<C�^<K_<��_<e�`<&_a<,b<��b<{�b<�.c<�9c<c<�b<��b<�Zb<�b<F�a<�a<�a<ța<e�a<ça<��a<]�a<{b<y_b<0�b<��b<B-c<�Mc<�Hc<�c<B�b<`5b<e�a<��`<6$`< }_< �^<�^<\e^<�j^<��^<_<��_<<J`<�a<�a<wTb<L�b<c&c<8Mc<�Ic<~#c<��b<�b<�Tb<jb<�a<�a<��a<�a<�a<?�a<��a<j�a<8b<R}b<��b<�c<�=c<Rc<�>c<��b<��b<� b<Ta<K�`<�_<�J_<+�^<~^<�`^<x^<��^<W:_<��_<�`<?a<a�a<˂b<a�b<j8c<PPc<�?c<}c<��b<0�b<�<b<�b<�a<ȷa<!�a<֣a<�a<�a<A�a<�b<�Ib<9�b<��b<�c<?Cc<�Jc< )c<��b<`b<��a<�a<�Y`<��_<m_<��^<�i^<�]^<��^<\�^<)f_<�
`<�`<�va<b<�b<
c<�?c<�Hc<",c<�b<{�b<yab<db<��a<^�a<�a<��a<��a<�a<��a<O�a<Gb<+Nb<Ԗb<w�b<�c<�4c<.c<�b</�b<�b<�oa<��`<`<�X_<�^<wn^<#?^<6D^<p}^<��^<�v_<"`<E�`<<�a<2+b<��b<3�b<}"c<mc<��b<B�b<�ob<�&b<��a<��a<�a<~a<va<�xa<��a<ءa<_�a<�b<�Jb<�b<3�b<c<c<�c<"�b<�^b<��a<�a<�g`<F�_<�_<=�^<.I^<,^<�C^<R�^<h_<��_<T`<za<�  �  �ca<	b<$�b<��b<>�b<��b<3�b<ާb<�wb<eNb<o0b<�b<�b<�b<�b<�b<Vb<�#b<�8b<WZb<��b<Էb<��b<��b<��b<��b<�tb<��a<�Fa<ф`<.�_<F�^<S^<��]<��]<A�]<��]<i^<m�^<#i_<n3`</�`<A�a<JMb<޻b<V�b<c<�c<��b<��b<Їb<�bb< Jb<�<b<A8b<G8b<d9b<�;b<�Ab<Pb<�ib<Ïb<
�b<�b<�c<C)c<�c<�b<vb<��a<!0a<�h`<�_<h�^<�I^<�]<��]<8�]<��]<xg^<1
_<T�_<0�`<vXa<b<��b<0�b<�c<~(c<�c<�b<ѷb<U�b<.ib<�Sb<�Hb<XEb<�Db<!Eb<�Fb<jNb<_b<�{b<4�b<��b<Hc<#c<�)c<c<��b<�Ib<u�a<N�`<�#`<]_<��^<^<�]<��]<[�]<^<p�^<xG_<�`<Y�`<��a<�8b<,�b<~c<{&c<}#c<�c<6�b<��b<:}b<�^b<Mb<�Db<ZBb<�Ab<$Bb<�Db<�Nb<�bb<��b<�b<2�b<?
c<�#c<�c<��b<:�b<b<�ha</�`<��_<�_<�r^<��]<k�]<��]<��]<r5^<r�^<	�_<L`<|a<�a<�ab<q�b<"c<�"c<�c<��b<o�b<��b<Ygb<xLb<0=b<I6b<4b<�2b<�2b<�6b<
Cb<qZb<y~b<��b<��b<s c</c<��b<��b<Xb<y�a<Wa<�F`<�{_<e�^<�$^<��]<��]<��]<��]<�?^<Q�^<�_<�k`<�/a<��a<�eb<��b<��b<�b<��b<R�b<\�b<.]b<Y:b<H$b<�b<�b<�b<�b<7b<}b<�,b<gIb<�qb<p�b<��b<B�b<��b<��b<+�b<�b<�va<�`<��_<~(_<�v^<@�]<W�]<�m]<�]<��]<�e^<_<��_<�`<�  �  �a<c�a<�Gb<T�b<��b<��b<d�b<��b<��b<yb<grb<�ub<�~b<Z�b<@�b<{�b<~b<�vb<�ub<�b<��b<n�b<��b<u�b<��b<��b<8b<�a<��`<�)`<�Q_<��^<��]<�H]<��\<��\<� ]<ݐ]<4^<~�^<x�_<�`<�ka<kb<'�b<h�b<��b<C�b<��b<�b<2�b<.�b<~�b<Q�b<|�b<��b<�b<��b<!�b<��b<��b<��b<��b<��b<��b< c<��b<6�b<)6b<R�a<J�`<]	`<�1_<�i^<\�]<�L]<�]<�]<Qa]<��]<U�^<T__<�7`<(a<��a<�Qb<�b<��b<�c<'�b<��b<A�b<f�b<��b<^�b<�b<�b<�b<f�b<�b<ħb<��b<�b<��b<��b<7�b<�c<;�b<H�b<*�b<�b<�^a<n�`<�_<`�^<;,^<,�]<�1]<�]<'*]<�]<�^<@�^<�_<`<�Ha<��a<�xb<��b<5�b<�c<�b<�b<Һb<�b<
�b<R�b<��b<�b<G�b<�b<©b<��b<ݟb<%�b<�b<��b<(�b<  c<}�b<��b<N[b<��a<�a<(K`<�r_<9�^<3�]<�g]</]<�
]<�=]<٬]<O^<W_<�_<Z�`<s�a<� b<��b<,�b<��b<=�b<��b<��b<��b<әb<�b<��b<��b<]�b<��b<S�b<D�b<�b<��b<b�b<\�b<>�b<��b<�b<��b<Éb<+b<�{a<��`<m�_<�_<�E^<��]<D']<c�\<��\<6:]<�]<yj^< 7_<(`<=�`<A�a<�'b<΍b<��b<V�b<�b<�b<��b<&�b<�tb<�tb<�{b<b�b<��b<�b<�~b<�ub<aqb<�vb<�b<[�b<��b<��b<C�b<�b<�Rb< �a<�*a<Pc`<��_<޶^<��]<}_]<��\<N�\<��\<R]<��]<�^<?t_<�L`<�  �  @�`<#�a<�b<�yb<��b<m�b<i�b<8�b<��b<�b<T�b<��b<d�b<��b<��b<��b<��b<��b<b�b<L�b<9�b<F�b<X�b<��b<��b< rb<�b<�za<��`<��_<�_<�5^<�z]<o�\<��\<9�\<<�\<�8]<'�]<�^<�_<�o`<�8a<�a<Zb<a�b<��b<��b<C�b<��b<�b<I�b<E�b<�b<�b<��b<h�b<l�b<!�b<L�b<��b<�b<��b<y�b<8�b<��b<?�b<~b<i	b<0ia<�`<��_<�^<h^<k]<��\<�\<R�\<U]<ی]<D^<�_<��_<]�`<��a<&b<��b<L�b<�b<��b<G�b<��b<4�b<��b<��b<\�b<��b<�c<�b<?�b<��b<#�b<��b<��b<��b<k�b<*�b<��b<�b<r\b<�a<�*a<�\`<�}_<ڠ^<��]<�:]<C�\< �\<��\< ,]<1�]<��^<d_<�C`<!a<��a<�Nb<9�b<��b<[�b<�b<��b<��b<ۿb<�b<�b<l�b<u�b< c<i�b<W�b<��b<��b<��b<��b<��b<��b<>�b<��b<�b<(0b<F�a<��`<`<�-_<�U^<5�]<~]<�\<�\<�\<�T]<�]<��^<��_<2�`<�Na<N�a<mb<�b<��b<��b<8�b<��b<��b<�b<��b<Q�b<�b<R�b<��b<��b<E�b<C�b<Z�b<��b<��b<.�b<�b<��b<w�b<�ab<p�a<�Ia<;�`<�_<�^<y�]<[F]<<�\<͌\<��\<?�\<^e]<-^<_�^<=�_<p�`<Oea<G�a<�fb<g�b<��b<��b<d�b<�b<�b<��b<1�b<%�b<D�b<��b<��b<n�b<�b<�b<J�b<��b<Z�b<¯b<_�b<��b<�b<)b<��a<��`<�(`<|I_<hl^<��]<]<��\<�x\<?�\<��\<��]<}U^<C1_<8`<�  �  ��`<=�a<ub<�kb<�b<�b<۫b<�b<�b<Ęb<!�b<@�b<��b<K�b<F�b<&�b<0�b<*�b<�b<�b<��b<�b<��b<��b<��b<�cb<+�a<9ia<s�`<>�_<��^<�^<U]]<�\<.{\<zl\<�\<�]<�]<��^<�{_<�[`<�&a<��a<�Kb<S�b<��b< �b<�b<�b<�b<ڻb<��b<�b<P�b<Tc<\c<�c<��b<R�b<��b<��b<��b<��b<��b<(�b<_�b<bob<6�a<*Wa<ܐ`<��_<�^<��]<:M]<��\<5�\<��\<��\<jo]<�(^<C_<�_<�`<}a<=b<��b<��b< �b<$�b<{�b<��b<<�b<��b<��b<��b<c<c<c<�c<��b<w�b<�b<�b< �b<K�b<��b<C�b<��b<WMb<d�a<a<�G`<�f_<Ɇ^<�]<]<ڲ\<_�\<	�\<]<d�]<_n^<�L_<�.`<aa<��a<p?b<��b<C�b<��b<��b<S�b<A�b<��b<��b<��b<�c<�c<dc<�c<�b<?�b<Y�b<Q�b<1�b<v�b<��b<\�b<��b<�b<~ b<ۋa<o�`<��_<�_<�:^<�|]<�\<��\<$�\<�\<�6]<��]<W�^<�_<�r`<�<a<��a<>^b<�b<��b<�b<
�b<��b<�b<|�b<*�b<L�b<U�b<c<�c<H�b<��b<J�b<v�b<��b<��b<{�b<��b< �b<��b<�Rb<@�a<�7a<'p`<��_<�^<��]<y(]<4�\<l\<!s\<��\<�G]<� ^<�^<��_<��`<�Sa<n�a<]Xb<�b<x�b<�b<��b<�b<�b<�b<B�b<l�b<Q�b<��b<��b<�b<�b<@�b<��b<��b<��b<��b<.�b<Q�b<qrb<�b<ѓa<D�`<�`<Y2_<\R^<e�]<y�\<I~\<�W\<�v\< �\<�t]<";^<�_<F�_<�  �  @�`<#�a<�b<�yb<��b<m�b<i�b<8�b<��b<�b<T�b<��b<d�b<��b<��b<��b<��b<��b<b�b<L�b<9�b<F�b<X�b<��b<��b< rb<�b<�za<��`<��_<�_<�5^<�z]<o�\<��\<9�\<<�\<�8]<'�]<�^<�_<�o`<�8a<�a<Zb<a�b<��b<��b<C�b<��b<�b<I�b<E�b<�b<�b<��b<h�b<l�b<!�b<L�b<��b<�b<��b<y�b<8�b<��b<?�b<~b<i	b<0ia<�`<��_<�^<h^<k]<��\<�\<R�\<U]<ی]<D^<�_<��_<]�`<��a<&b<��b<L�b<�b<��b<G�b<��b<4�b<��b<��b<\�b<��b<�c<�b<?�b<��b<#�b<��b<��b<��b<k�b<*�b<��b<�b<r\b<�a<�*a<�\`<�}_<ڠ^<��]<�:]<C�\< �\<��\< ,]<1�]<��^<d_<�C`<!a<��a<�Nb<9�b<��b<[�b<�b<��b<��b<ۿb<�b<�b<l�b<u�b< c<i�b<W�b<��b<��b<��b<��b<��b<��b<>�b<��b<�b<(0b<F�a<��`<`<�-_<�U^<5�]<~]<�\<�\<�\<�T]<�]<��^<��_<2�`<�Na<N�a<mb<�b<��b<��b<8�b<��b<��b<�b<��b<Q�b<�b<R�b<��b<��b<E�b<C�b<Z�b<��b<��b<.�b<�b<��b<w�b<�ab<p�a<�Ia<;�`<�_<�^<y�]<[F]<<�\<͌\<��\<?�\<^e]<-^<_�^<=�_<p�`<Oea<G�a<�fb<g�b<��b<��b<d�b<�b<�b<��b<1�b<%�b<D�b<��b<��b<n�b<�b<�b<J�b<��b<Z�b<¯b<_�b<��b<�b<)b<��a<��`<�(`<|I_<hl^<��]<]<��\<�x\<?�\<��\<��]<}U^<C1_<8`<�  �  �a<c�a<�Gb<T�b<��b<��b<d�b<��b<��b<yb<grb<�ub<�~b<Z�b<@�b<{�b<~b<�vb<�ub<�b<��b<n�b<��b<u�b<��b<��b<8b<�a<��`<�)`<�Q_<��^<��]<�H]<��\<��\<� ]<ݐ]<4^<~�^<x�_<�`<�ka<kb<'�b<h�b<��b<C�b<��b<�b<2�b<.�b<~�b<Q�b<|�b<��b<�b<��b<!�b<��b<��b<��b<��b<��b<��b< c<��b<6�b<)6b<R�a<J�`<]	`<�1_<�i^<\�]<�L]<�]<�]<Qa]<��]<U�^<T__<�7`<(a<��a<�Qb<�b<��b<�c<'�b<��b<A�b<f�b<��b<^�b<�b<�b<�b<f�b<�b<ħb<��b<�b<��b<��b<7�b<�c<;�b<H�b<*�b<�b<�^a<n�`<�_<`�^<;,^<,�]<�1]<�]<'*]<�]<�^<@�^<�_<`<�Ha<��a<�xb<��b<5�b<�c<�b<�b<Һb<�b<
�b<R�b<��b<�b<G�b<�b<©b<��b<ݟb<%�b<�b<��b<(�b<  c<}�b<��b<N[b<��a<�a<(K`<�r_<9�^<3�]<�g]</]<�
]<�=]<٬]<O^<W_<�_<Z�`<s�a<� b<��b<,�b<��b<=�b<��b<��b<��b<әb<�b<��b<��b<]�b<��b<S�b<D�b<�b<��b<b�b<\�b<>�b<��b<�b<��b<Éb<+b<�{a<��`<m�_<�_<�E^<��]<D']<c�\<��\<6:]<�]<yj^< 7_<(`<=�`<A�a<�'b<΍b<��b<V�b<�b<�b<��b<&�b<�tb<�tb<�{b<b�b<��b<�b<�~b<�ub<aqb<�vb<�b<[�b<��b<��b<C�b<�b<�Rb< �a<�*a<Pc`<��_<޶^<��]<}_]<��\<N�\<��\<R]<��]<�^<?t_<�L`<�  �  �ca<	b<$�b<��b<>�b<��b<3�b<ާb<�wb<eNb<o0b<�b<�b<�b<�b<�b<Vb<�#b<�8b<WZb<��b<Էb<��b<��b<��b<��b<�tb<��a<�Fa<ф`<.�_<F�^<S^<��]<��]<A�]<��]<i^<m�^<#i_<n3`</�`<A�a<JMb<޻b<V�b<c<�c<��b<��b<Їb<�bb< Jb<�<b<A8b<G8b<d9b<�;b<�Ab<Pb<�ib<Ïb<
�b<�b<�c<C)c<�c<�b<vb<��a<!0a<�h`<�_<h�^<�I^<�]<��]<8�]<��]<xg^<1
_<T�_<0�`<vXa<b<��b<0�b<�c<~(c<�c<�b<ѷb<U�b<.ib<�Sb<�Hb<XEb<�Db<!Eb<�Fb<jNb<_b<�{b<4�b<��b<Hc<#c<�)c<c<��b<�Ib<u�a<N�`<�#`<]_<��^<^<�]<��]<[�]<^<p�^<xG_<�`<Y�`<��a<�8b<,�b<~c<{&c<}#c<�c<6�b<��b<:}b<�^b<Mb<�Db<ZBb<�Ab<$Bb<�Db<�Nb<�bb<��b<�b<2�b<?
c<�#c<�c<��b<:�b<b<�ha</�`<��_<�_<�r^<��]<k�]<��]<��]<r5^<r�^<	�_<L`<|a<�a<�ab<q�b<"c<�"c<�c<��b<o�b<��b<Ygb<xLb<0=b<I6b<4b<�2b<�2b<�6b<
Cb<qZb<y~b<��b<��b<s c</c<��b<��b<Xb<y�a<Wa<�F`<�{_<e�^<�$^<��]<��]<��]<��]<�?^<Q�^<�_<�k`<�/a<��a<�eb<��b<��b<�b<��b<R�b<\�b<.]b<Y:b<H$b<�b<�b<�b<�b<7b<}b<�,b<gIb<�qb<p�b<��b<B�b<��b<��b<+�b<�b<�va<�`<��_<~(_<�v^<@�]<W�]<�m]<�]<��]<�e^<_<��_<�`<�  �  Y�a<BQb<P�b<�c< c<c<��b<B�b<+Tb<"b<�a<�a<�a<�za<wa<�}a<��a<��a<��a<� b<ib<O�b<��b<�c<K&c<c<��b<�=b<֡a<b�`<�8`<u�_<��^<؉^<K^<&@^<�i^<C�^<K_<��_<e�`<&_a<,b<��b<{�b<�.c<�9c<c<�b<��b<�Zb<�b<F�a<�a<�a<ța<e�a<ça<��a<]�a<{b<y_b<0�b<��b<B-c<�Mc<�Hc<�c<B�b<`5b<e�a<��`<6$`< }_< �^<�^<\e^<�j^<��^<_<��_<<J`<�a<�a<wTb<L�b<c&c<8Mc<�Ic<~#c<��b<�b<�Tb<jb<�a<�a<��a<�a<�a<?�a<��a<j�a<8b<R}b<��b<�c<�=c<Rc<�>c<��b<��b<� b<Ta<K�`<�_<�J_<+�^<~^<�`^<x^<��^<W:_<��_<�`<?a<a�a<˂b<a�b<j8c<PPc<�?c<}c<��b<0�b<�<b<�b<�a<ȷa<!�a<֣a<�a<�a<A�a<�b<�Ib<9�b<��b<�c<?Cc<�Jc< )c<��b<`b<��a<�a<�Y`<��_<m_<��^<�i^<�]^<��^<\�^<)f_<�
`<�`<�va<b<�b<
c<�?c<�Hc<",c<�b<{�b<yab<db<��a<^�a<�a<��a<��a<�a<��a<O�a<Gb<+Nb<Ԗb<w�b<�c<�4c<.c<�b</�b<�b<�oa<��`<`<�X_<�^<wn^<#?^<6D^<p}^<��^<�v_<"`<E�`<<�a<2+b<��b<3�b<}"c<mc<��b<B�b<�ob<�&b<��a<��a<�a<~a<va<�xa<��a<ءa<_�a<�b<�Jb<�b<3�b<c<c<�c<"�b<�^b<��a<�a<�g`<F�_<�_<=�^<.I^<,^<�C^<R�^<h_<��_<T`<za<�  �  �b<A�b<t�b<�0c<�<c<
c<��b<�b<1b<ɶa<�[a<�a<��`<��`<`�`</�`<��`<i#a<�qa<V�a<�7b<��b<3�b<1/c<�Ec<�0c<{�b<�b<k�a<^a<Y�`<�*`<�_<�R_<}_<�_<[8_<��_<=�_<*�`<�a<��a<AVb<��b<�(c<�Sc<�Qc<J'c<��b<y~b<�b<��a<�aa<� a<��`<��`<��`<��`<x a<�aa<��a<�b<�b<�b<p3c<dc<�lc<wHc<��b<��b<��a<�Pa<�`<�$`<0�_<la_<�:_<-?_<�n_<��_<�@`<z�`<xra<�b<��b<�c<VSc<�mc<�\c<?%c<��b<}nb<�b<�a<�Xa<�a<�`<a�`<��`<�
a<�<a<��a<�a<�Ab<h�b<�c<Jc<Cmc<�fc<�2c<��b<�Rb<Ӻa<xa<a�`<��_<��_< O_<�6_<J_<�_<�_<�o`<a<3�a<�Ab<��b<�(c<rac<�lc<�Mc<�c<)�b<!Kb<o�a<?�a<�@a<ma<��`<��`<1�`<Ca<�Ma<e�a<8�a<�_b<��b<lc<�Tc<Fjc<�Tc<�c<��b<Pb<�a<+�`<9K`<��_<�q_<=_<�3_<lU_<��_<g`<4�`<�8a<`�a<5lb<��b<Q;c<�dc<�`c<\4c<��b<t�b<db<@�a<\da<� a<��`<��`<H�`<��`<�a<�Ta<��a<�b<�nb<��b<"c<�Jc<�Qc<�+c<��b<�ab<��a<�.a<�`<� `<8�_<�;_<P_<b_<�G_<*�_<�`<?�`<�Ia<�a<~sb<��b<8)c<CCc<�1c<b�b<3�b<GAb<��a<�ya<�)a<��`<��`<��`<u�`<C�`<�
a<�Qa<��a<�b<�ub<��b<-c<3:c<:3c<��b<
�b<�b<c�a<��`<~K`<��_<x\_<_<�_<X_<tS_<	�_<�;`<��`<�ua<�  �  �Tb<N�b<Kc<�Cc<�Bc<Nc<��b<�Ob<<�a<4Ja<�`<zi`<�`<_�_<��_<j�_<R-`<Z�`<��`<�ja<��a<�ob<��b<�)c<�Nc<�Fc<�c<+�b<�Db<��a<@a<�`< g`<� `<$�_<��_<'`<�G`<��`<a<��a<Wb<>�b<��b<�Dc<fbc<4Sc<�c<l�b<HCb<��a<t?a<��`<rn`<l-`<�`<#`<}+`<~k`<j�`<<a<��a<�Cb<2�b<#c<�cc<�yc<�bc<X!c<Q�b<�Bb<L�a<�=a<U�`<r`<�4`<3`<�`<�>`<l�`<$�`<qWa<��a<�\b<��b<�1c<�jc<Oxc<%Yc<�c<v�b<�)b<l�a<�&a<׸`<Tc`<�+`<�`<,`<CG`<)�`<a�`<�la<��a<sb<�b<w?c<�qc<*xc<�Qc<c<��b<b<��a<�a<t�`<�Y`<�&`<4`<�"`<R`<��`<ga<K�a<ib<�b<��b<sIc<otc<�rc<&Ec<Q�b<�~b<�a<�xa<H�`<V�`<K`<[`<$`<>$`<tX`<��`<5a<`�a<�b<��b<�c<<Oc<+sc<[jc<�5c<��b<�fb<�a<�`a<l�`<͆`<�?`<�`<r`<K*`<�c`<�`<2*a<|�a<�-b<D�b<mc<WWc<Xsc<Ebc<�%c<��b<KLb<k�a<+Da<w�`<�n`<y+`<�`<�`<�"`<�``<V�`<�,a<(�a<�0b<ɩb<�c<�Jc<�^c<KFc<'c<��b<�!b<�a<ya<�`<�L`<`<��_<��_<�`<�Z`<1�`<3/a</�a< 4b<��b<�c<�@c<�Mc<.c<��b<{b<��a<�wa<U�`<͉`<�3`<o�_<#�_<'�_<�`<�^`<��`<�:a<h�a<�@b<a�b<�c<�>c<�Dc<'c<%�b<nab<��a<�\a<��`<Au`<B$`<��_<�_<�_<i`<Tk`<��`<Oa<��a<�  �  څb<R�b<# c<�<c</c<��b<Ɏb<	b<�na<u�`<�6`<Ŵ_<�R_<+_<�_<�!_<�f_<T�_<�Y`<P�`<T�a<<.b<^�b<�c<�=c<�Bc<<c<��b<�{b<�b<ױa<�Ya<�a<��`<��`<��`<��`<� a<#>a<�a<!�a<"Yb<�b<�c<EGc<)Wc<;c<��b<�b<��a<�Wa<ݹ`<)`<~�_<�\_<0_<�._<Y_< �_<e"`<;�`<�Ra<��a<��b<g�b<RJc<Wmc<dc<�2c<��b<T�b<�b<7�a<aga<l(a<��`<%�`<E�`<Qa<:3a<eva<��a< 0b<��b<
�b<�>c<Thc<�hc<F<c<&�b<2hb<�a<3a<�`<�`<͞_<�U_<�6_<�B_<z_<��_<�W`<��`<��a<*b<�b<c<�\c<�oc<�Wc<c<�b<__b<�a<֛a<IOa<�a<g�`<�`<��`<Qa<�Ga<��a<E�a<�Rb<$�b<c<VQc<�mc<L_c<w#c<:�b<#8b<e�a<��`<�d`<}�_<�_<�C_<�2_<9M_<��_<��_<<�`<�a< �a<	Ub<P�b<�0c<5bc<�fc<7Ac<A�b<c�b<�6b<��a<Vza<�4a<=a<��`<��`<��`<�a<uYa<&�a<
b<�pb<$�b<%c<Zc<)hc<<Jc<�b<1�b<��a<�^a<��`<�+`<˱_<�Z_<�+_<g(_<ZP_<�_<N`<��`<8Aa<S�a</ob<�b<1c<URc<SGc<�c<��b<Iab<?�a<�a<Ca<Na<�`<��`<Z�`<��`<�a<kNa<��a<xb<�mb<��b<ec<[>c<N>c<Ac<��b<�;b<�a<ta<�h`<��_<To_<�%_<%_<�_<�H_<��_<�%`<�`<�[a<��a<M�b<=�b<�)c<�<c<<$c<��b<��b<�*b<!�a<�fa<�a<�`<��`<˳`<��`<��`<#a<�]a<߹a< b<�  �  àb<�b<Rc<�c<`c<ֽb<�Jb<��a<Oa<EL`<r�_<�_<��^<�D^<�0^<:Q^<e�^<i#_<�_<�x`<�0a<�a<�mb<u�b<�c<�(c<c<i�b<1�b<�Rb<�b<Z�a<9�a<f�a<��a<.�a<N�a<��a<��a<��a<<b<�b<��b<�c<T3c<�5c<hc<ڷb<�8b<�a<��`<8/`<p�_<��^<��^<�[^<�Y^<y�^<��^<"|_<�%`<�`<��a<�9b<Ծb<Cc<�Jc<yNc<�-c<��b<�b<�bb<�!b<��a<��a<�a<$�a<��a<͵a<c�a<&�a<"-b<apb<-�b<��b<�5c<zOc<Cc<Y
c<<�b<�b<�oa<��`<�`<�`_<d�^<��^<�`^<�o^<$�^<7#_<��_<�h`<!a<}�a<Vmb<��b<�1c<UQc<~Gc<�c<O�b<��b<<Kb<�b<�a<{�a<�a<�a<��a<��a<G�a<Fb<�Bb<Q�b<#�b<�c<�Bc<cPc<�5c<��b<Vzb<��a<�2a<�z`<l�_<�/_<��^<�q^<�\^<�|^<.�^<pM_<G�_<�`<tXa<�b<��b<x�b<!;c<Lc<6c<�c<��b<�sb<l/b<��a<�a<��a<l�a<>�a<��a<��a<�a<Ab<	Ub<��b<��b<"c<.Fc<�Fc<�c<�b< Db<��a<��`<�3`<��_<�^<��^<jW^<nS^<˃^<�^<o_<�`<��`<�a<$b<k�b<�c<|/c<�1c<�c<��b<��b<�@b<g�a<a�a<��a<�a<��a<�a<m�a<��a<&�a<�b<�Gb<_�b<��b<4c<�%c<�c<l�b<�yb<��a<Ca<��`<��_<?2_<�^<�V^<�0^<�>^<�^<��^<�_<�6`<��`<�a<�:b<�b<��b<�c<�c<j�b<ʧb<�]b<b<��a<��a<߉a<Zxa<�ra<Twa<��a<��a<:�a<nb<]Vb<�  �  �b<X�b<��b<.�b<��b<~b<	 b<R[a<��`<��_<s_<-`^<`�]<�]<�r]<ԗ]<1�]<��^<\9_<�`<6�`<ׇa<�%b<�b<��b<� c< �b<��b<�b<{b<�Sb<t8b</)b<�"b< "b<�"b<T$b<8)b<�5b<�Lb<qb<+�b<��b<��b<8c<jc<��b<�tb<��a<O;a<w`<<�_<�^<9P^<X�]<��]<y�]<�]<�F^<��^<��_<Km`<:5a<��a<^zb<c�b<c<�*c<Dc<+�b<r�b<ܔb<�pb<Yb<`Lb<�Gb<eFb<;Fb<#Gb<�Lb<`[b<�ub<��b<��b<��b<bc<�(c<�c<�b<,^b<,�a<�a<�C`<?{_<+�^<�1^<��]<¢]<̳]<s�]<k^<`(_<�_<�`<fxa<!b< �b<6�b<�%c<�(c<�c<+�b<�b<ˆb<�fb<Sb<nIb<�Fb<Fb<RFb<uHb<Qb<$cb<��b<��b<��b<2c<@%c<�%c<# c<٭b<g/b<M�a<\�`<�_<T:_<��^<h^<s�]<��]<+�]<� ^<��^<qb_<�)`<��`<a�a<dKb<��b<�c<-$c<�c<:�b<��b<Q�b<�tb<�Xb<Ib<?Bb<�@b<�@b<�Ab<�Eb<,Qb<Ugb<#�b<�b<��b<yc<$c<�c<��b<ǁb<��a<hDa<~`<�_<��^<�P^<i�]<z�]<�]<d�]<�;^<��^<i�_<�[`<�!a<r�a<�bb<�b<��b<$c<��b<Z�b<I�b<{rb<.Mb<�4b< 'b<�!b<�b<6b<�b<=%b<Z3b<9Mb<osb<�b<��b<��b<�b<��b<7�b<�2b<!�a<;�`<�`<AM_<��^<k^</�]<�r]<%�]<m�]<N^<��^<2�_<]�`<Fa<a�a<qb<��b<
�b<��b<��b<��b<�|b<�Qb<%1b<pb<�b<�b<jb<�b<eb<ab<�.b<Nb<�xb<�  �  Φb<��b<l�b<n�b<�b<eBb<�a<�a<�B`<�j_<��^<��]<O]<��\<�\<�]<�k]<^<{�^<Y�_<v`<�<a<f�a< ab<s�b<��b<b�b<��b<�b<��b<;�b<6~b<��b<�b<��b<ܗb<m�b<S�b<�b<�b<��b<S�b<"�b<F�b<��b<��b<�b<#6b<��a<d�`<�`<zB_<{w^<��]<LM]<�	]<q]<;F]<��]<�j^<^5_<�`<�`<�a<�:b<��b<��b<hc<%�b<��b<M�b<�b<"�b<�b<��b<��b<R�b<T�b<²b<d�b<��b<��b<�b<��b<\�b< c<( c<��b<ޔb<�b<�za<�`<�_<�_< H^<e�]<v<]<;]<�]<r]<��]<в^<]�_<(\`<�)a<��a<zgb<i�b<��b<�c<��b<��b<�b<��b<�b<�b<�b<ݷb<��b<w�b<��b<-�b<�b<�b<3�b<N�b<��b<�c<0�b<-�b<,rb<E�a<�<a<kq`<ʘ_<W�^<3^<�{]<�"]<�]<�0]<�]<�0^<u�^<}�_<j�`<!ca<	b<��b<��b<V�b<4�b<�b<��b<ܳb<�b<��b<s�b<��b<u�b<�b<Ұb<קb<��b<l�b<�b<�b<d�b<��b<��b<��b<B�b<eCb<�a<��`<� `<BG_<z^<�]<_K]<�]< ]<�=]<�]<v]^<&_<-�_<��`<e�a<�#b<��b<t�b<��b<��b<��b<�b<��b<��b<��b<g�b<��b<��b<E�b<N�b<��b<�{b<c~b<��b<,�b<J�b<��b<Y�b<M�b<jb<b�a<Oa<}�`<ʹ_<��^<z^<Iy]<�]<�\<1�\<A]<F�]<=�^<�Q_<*`<u�`<Z�a<�4b<(�b<R�b<��b<M�b<1�b<�b<Uxb<Uob<Jqb<0yb<�b<҅b<��b<�zb<orb<�ob<mwb<�b<�  �  ��b< �b<��b<ƨb<�ub<�b<g�a<��`<�`<+'_<�L^<��]<��\<ї\<q}\<��\<�]<�]<�~^<�\_<�;`<�a<"�a<�7b<��b<��b<m�b<��b<��b<֝b<Ȝb<��b<T�b<Q�b<��b<~�b<��b<�b<´b<K�b<��b<ϭb<��b<X�b<��b<5�b<�vb<2
b<nqa<<�`<��_<?�^<�(^<�t]<�\<��\<�\<s�\< i]<�^<4�^<�_</�`<oa<�b<�b<f�b<x�b</�b<[�b<U�b<Q�b<��b<G�b<Z�b<t�b<�c<c<��b<��b<��b<��b<��b<�b<d�b<�b<��b<7�b<�kb<�a<�Ga<�~`<0�_<��^<��]<P]<��\<~�\<��\<�]<�]<�e^<�>_<p`<�`<�a<�<b<�b<��b<J�b<��b<v�b<��b<�b<|�b<��b<2�b<��b<_c<��b<��b<9�b<�b<0�b<C�b<7�b<�b<�b<��b<=�b<�Gb<��a<�a<�5`<QU_<`z^<P�]<�!]</�\<=�\<��\<e=]<��]<k�^<��_<	c`<a/a<��a<\b<��b<�b<8�b<��b<a�b<�b<��b<��b<D�b<��b<��b<��b<j�b<��b<M�b<��b<ѽb<��b<G�b<�b<��b<Z�b<�b<xb<�|a<]�`<��_<
_<J+^<�t]<�\<a�\<z�\<��\<4^]<�^<��^<�_<��`<�Ya<�a<�hb<B�b<��b<��b<y�b<�b<ޡb<?�b<ǯb<�b<n�b<1�b<�b<u�b<��b<��b<��b<i�b<I�b<U�b<��b<ڷb<��b<-Ab<��a<�a<�Q`<�s_<ה^<�]<� ]< �\<i}\<?�\<�\<�v]<^4^<+_<Y�_<��`<Eya<�	b<�lb<��b<L�b<��b<��b<w�b<��b<ӓb<֣b<D�b<��b<��b<0�b<��b<k�b<ѕb<q�b<�b<�  �  mgb<�nb<Xlb<�Wb<�(b<-�a<na< �`<�G`<L�_<�_<t^<�^<�]<��]<��]<^<R�^<'_<��_<lp`<�
a<��a<"�a<y=b<�fb<�wb<Ixb<�pb<�hb<�db<�fb<Dnb<�vb<Z}b<.b<;|b<�ub<�nb<�kb<ob<vwb<��b<[�b<��b<�db<�,b<��a<d_a<s�`<�.`<b�_<N�^<l^<�^<A�]<��]<�^<e^<�^<\�_<�(`<s�`<�`a<%�a<9b<vb<��b<�b<��b<
�b<��b<�b<P�b<�b<Q�b<~�b<Ġb<H�b<#�b<��b<{�b<-�b<V�b<��b<�b<��b<�jb<�'b<��a<Da<n�`<`<Gd_<��^<1U^<�^<��]<��]<�+^<c�^<Q _<߿_<�e`<�a<��a<�b<8Sb<��b<D�b<��b<X�b<Q�b<�b<G�b<��b<��b<=�b<�b<��b<�b<ېb<݊b<��b<K�b<�b<�b<�b<��b<dXb<P
b<ǜa<Ga<�u`<��_<�._<��^<�2^<��]<��]<)�]<�F^<X�^<dO_<:�_<�`<�0a<�a<�b<!ab<ډb<-�b<
�b< �b<g�b< �b<p�b<S�b<a�b<*�b<D�b<�b<.�b<H�b<%�b<�b<�b<��b<��b<��b<�tb<`;b<�a<�ia<�`<s5`<Ԏ_<��^<Kl^<�
^<%�]<K�]<V�]<zZ^<c�^<�s_<�`<��`<*La<��a<� b<\b<�zb<b<
b<+ub<zlb<�hb<2kb<�qb<�xb<&|b<�zb<�tb<^lb<�db<bb<deb<9mb<$ub<vb<ygb<1Ab<q�a<ڙa<�a<w�`<��_<7_<�^<�&^<��]<U�]<�]<��]<�d^<��^<ӎ_<�4`<J�`<_a<��a<� b<�Rb<'jb<+nb<�gb<J^b<�Wb<�Vb<�[b<�cb<�jb<amb<Pkb<
eb<6]b<�Wb<�Wb<^b<�  �  Mgb<rqb<=qb<E^b<1b<,�a<�ya<��`<�V`<�_<l_<܈^<�^<s�]<��]<�]<3^<��^<b9_<��_<�~`<Ta<1�a<��a<xEb<Amb<H|b<ozb<pb<�db<\]b<\b<�_b<Ffb<�kb<cmb<kb<Efb<�bb<�bb<dib<$ub<��b<�b<:�b<lb<�5b<�a<hka<��`<J>`<��_<�_<f�^<:#^<��]<@�]<�^<|z^<��^<�_<F8`<%�`<�la<��a<Bb<�}b<X�b<��b<ܞb<�b<@�b<U�b<O�b<��b<Q�b<��b<�b<z�b<v�b<��b<��b<��b<?�b<z�b<(�b<�b<�rb<1b<��a<�Pa<��`<`<Qv_<��^<	k^<�^<i�]<[^<>B^<]�^<Z3_<��_<�t`<�a<��a<�b<�[b<|�b<^�b<��b<��b<C�b<��b<��b<K�b<v�b<��b<�b<+�b<Ĉb<9�b<̀b<�b<�b<��b<��b<֡b<[�b<�`b<Ob<P�a<2 a<��`<\�_<zA_<y�^<I^<^<��]<p^<�\^<��^<�a_<n`<s�`<?=a<T�a<$b<"ib<>�b<��b<2�b<J�b<\�b<�}b<�{b<�~b<��b<��b<w�b<^�b<��b<�|b<,|b<[�b<��b<��b<~�b<0�b<I|b<3Db<��a<�ua<��`<�D`<�_<5_<��^<E!^<��]<��]<3^<�o^<6�^<1�_<�'`<o�`<XXa<k�a<�)b<�cb<��b<��b<N�b<>sb<0gb<0`b<4_b<�bb<�gb<djb<4ib<db<�]b<nYb<&Zb<�`b<"lb<wb<Nzb<�mb<	Ib<�b<�a<(%a<��`<��_<#I_<$�^<�<^<��]<�]<��]<#^<�y^<�_<��_<�C`<\�`<�ja<��a<4)b<�Yb<Cob<'qb<�gb<>[b<UQb<Mb<�Nb<�Sb<DYb<�[b<�Yb<�Tb<�Ob<�Mb<:Qb<�Zb<�  �  Yeb<wb<!~b<�pb<FHb<� b<w�a<�a<.�`<H�_<�J_<��^<�]^<^<�^<)^<�r^<��^<tn_<
`<��`<;a<�a</b<�[b<�~b<ćb<�~b<&lb<MWb<�Eb<�:b<6b<�5b<37b<8b<�8b<$9b<f=b<6Gb<�Wb<mb<`�b<N�b<�b<J�b<VNb<��a<Ќa<�a<�j`<�_<Z;_<&�^<"e^<5^<�3^<�`^<��^<�3_<��_<ne`<xa<�a<:b<[b<R�b<̫b<ܭb<��b<�b<�wb<�gb<$^b<BZb<(Zb<�Zb<>Zb<OYb<�Yb<e^b<
ib<4zb<M�b<�b<�b<��b<��b<-Kb<$�a<�sa<,�`<�F`<��_<>_<V�^<�\^<�:^<5H^<f�^<�^<�j_<�`<�`<�7a<�a<�'b<Nsb<��b<�b<k�b<��b<�b<|qb<�cb<#\b<�Yb<cZb<�Zb<DZb<oYb<[b<�ab<�nb<��b<��b<��b<��b<�b<�wb<�/b<.�a<&Ea<�`<�`<�w_<��^<̉^<�I^<7^<�S^<��^<�_<˖_<�1`<��`<aa<>�a<�>b<qb<��b<$�b<��b<\�b<�wb<fb<�Zb<Ub<,Tb<�Tb<&Ub<�Tb<wTb<�Wb<c`b<�ob<��b<��b<�b< �b<�b<�\b<r	b<a�a<:a<Uq`<u�_<�=_<V�^<-c^<�0^<Q-^<mX^<8�^<M'_<3�_<�T`<��`<Pza<��a<�Bb<Xxb<3�b<��b<�b<Clb<�Vb<~Eb<;b<R6b<z5b<05b<_4b<�2b<�2b<G7b<�Ab<kRb<.gb<�zb<�b<p~b<�^b<� b<N�a<IHa<(�`<�`<}_<q�^<�{^<�-^<�^<s^<BS^<��^<�9_<��_<�n`<�a<�a<��a<�@b<�lb<�|b<xb<�fb<Qb<D=b<//b<�'b<;%b<�%b<$&b<&b<|%b<�'b<�.b<<b<qOb<�  �  �^b<F}b<b�b<��b<�hb<�'b<��a<sMa<��`<-`<͞_<O"_<��^<χ^<8w^<$�^<��^<�=_<,�_<qQ`<C�`<�oa<��a<@b<rzb<��b<ԕb<��b<|bb<?b<b<�b<_�a<��a<��a<��a<��a<j�a<��a<Ob<~8b<#]b<�b<ɜb<`�b<��b<qb<�&b<ؽa<=a<��`<=`<~�_<d_<�^<��^<a�^<f�^<�_<#�_<E`<W�`<�;a<��a<�.b<�~b<o�b<�b<y�b<��b<�}b<Zb<o:b<"b<�b<Gb<Vb<�b<-	b<�b<v%b<|?b<B`b<�b<�b<�b<޽b<�b<Lpb<b<��a<�a<�`<l�_<�w_<[_<O�^<�^<Y�^<-�^<oE_<��_<�L`<��`<oa<=�a<�Ob<o�b<,�b<(�b<j�b<`�b<�qb<�Nb<31b<�b<�b<kb<	b<�b<@b<-b<�-b<WJb<�lb<g�b<Z�b<�b<��b<;�b<Wb<��a<�{a<��`<�Z`<��_<O_<��^<��^<f�^<��^<e _<+g_<��_<y`<a<ؕa<b<~db<1�b<��b<<�b<ƣb<��b<�_b<<>b<2#b<gb<�b<��a<��a<!b<�
b<'b<s1b<ePb<�sb<5�b<X�b<J�b<��b<yb<3b<d�a<�Ea<�`<�`<Δ_<�_<'�^<��^<�^< �^<l_<�_<�`<��`<)a<D�a<b<^fb<z�b<y�b<b�b<2�b<�]b<9b<Yb<�a<��a<��a<�a<��a<��a<��a<[�a<	b<y8b<�[b<a|b<��b<��b<�|b<�Eb<8�a<"|a<t�`<6``<!�_<�I_<��^<_�^<�v^<��^<��^<�_<��_<�`<B�`<s=a<Z�a<�b<�ab<p�b<�b<b<�ab<�=b<�b<��a<%�a<3�a<��a<��a<��a<a�a<��a<��a<�b<�:b<�  �  Ob<@}b<��b<��b<.�b<�Rb<��a<_�a<a<o�`<(`<ɗ_<�B_<G_<��^<|_<bT_<��_<}%`<��`<�.a<3�a<&b<�hb<�b<��b<S�b<�~b<�Nb<
b<��a<c�a<.�a<|a<�oa<Bna<-wa<Ƌa<īa<��a<�	b<~Ab<�vb<p�b<}�b<նb<ɕb<�Tb<7�a<�a<��`<fz`<d�_<Ș_<�N_<w'_<w&_<�K_<��_<{�_<�u`<��`<$�a<v�a<�]b<E�b<��b<e�b<��b</�b<db<�-b<��a<��a<��a<k�a<��a<ޑa<x�a<ϴa<9�a<b<%8b<�nb<�b<��b<��b<��b<�b<iKb<��a<�ga<��`<P_`<��_<B�_<!J_<�._<g9_<j_<U�_<�)`<Ĩ`<�.a<T�a<)"b<�{b< �b<C�b<��b<�b<f�b<�Qb<�b<�a<��a<�a<��a<2�a<��a<8�a<e�a<�a<^b<�Jb<��b<J�b<$�b<��b<ƹb<�b<Q+b<��a<;a<�`<a4`<��_<�n_<:_<+_<(B_<c~_<��_<N`<x�`<�Ua<R�a<y=b<W�b<��b<��b<��b<��b<-pb<�9b<
b<��a<0�a<s�a<g�a<>�a<V�a<�a<��a<��a<�!b<Xb<�b<��b<]�b<��b< �b<�`b<� b<��a<a<�~`<�`<��_<�L_<Z#_<4 _<SC_<��_<��_<Ig`<,�`<wna<��a<#Gb<�b<Ȱb<۶b<��b<�xb<IDb<�b<��a<֬a<��a<�ua<�ka<la<.wa<�a<"�a<��a<[b<rFb<bwb<�b<R�b<�b<�mb<s b<@�a<�;a<�`<�1`<�_<�[_<_<*�^<�	_<�9_<��_<��_<�w`<8�`<�~a<G�a<�Ib<��b<��b<��b<��b<�Sb<b<��a<޶a<L�a<�ra<�aa<�[a<�`a<rpa<��a<}�a<��a<�b<�  �  �2b<1rb<��b<t�b<�b<bxb<f.b<��a<�\a<`�`<�y`<�`<;�_<F�_<�_<�_<}�_<=0`<C�`<�a<�za<l�a<)Gb<��b<;�b<��b<��b<
pb<{.b<��a<ɚa<*Xa<
"a<{�`<6�`<��`<��`<za<�Ca<ׂa< �a<qb<�`b<l�b<�b<b�b< �b<~b<[,b<��a<Ta<L�`<�w`<X `<��_<��_<I�_<��_<�`<�t`<��`<FSa<��a<2b<��b<��b<p�b<I�b<'�b<ۂb<#=b<�a<P�a<�ia<�7a<3a<�a<�a<�a<�@a<�ua<��a<Yb<Lb<p�b<��b<|�b<+�b< �b<$yb<�b<�a<>a<@�`<�f`<$`<�_<��_<�_<�_<�@`<�`<�a<V�a<��a<kUb<��b<��b<A�b<Y�b<��b<mb<S$b<�a<��a<CWa<�*a<�a<na<�a<A&a<Qa<Ίa<�a<�b<9db<.�b<t�b<}�b<{�b<��b<0]b<X�a<�a<a<�`<�G`<��_<;�_<z�_<��_<�`<�Y`<�`<�-a<�a<�b<�lb<��b<�b<��b<5�b<�b<�Ob<Lb<�a<�wa<Aa<�a<�a<��`<a<�-a<�]a<��a<��a<�.b<�ub<�b<��b<~�b<o�b<��b<�6b<B�a<�Za<��`<
z`<� `<��_<Ӽ_<�_<Z�_<�`<h`<1�`<�Ba<��a<zb<rb<��b<��b<ɿb<%�b<pdb<jb<�a<S�a<�Fa<a<��`<��`<��`<_�`<a<�Na<!�a<��a<�#b<�fb<�b<�b<>�b<��b<Nb<��a<Ӆa<%a<`<�8`<��_<�_<h�_<�_<��_<@`<.m`<��`<�Na<�a<�#b<ypb<��b<��b<m�b<Nwb<�9b<��a<$�a<�^a<#a<B�`<q�`<L�`<��`<��`<�a<�Wa<��a<��a<�  �  Kb<@Yb<Z�b<E�b<��b<l�b<VVb<�b<s�a<�Fa<��`<۟`<Qf`<�C`<<:`<LJ`<�r`<��`<�a<�_a<(�a<�b<�kb<$�b<W�b<۷b<.�b<vSb<��a<סa<2Ba<'�`< `<_k`<|M`<�H`<8]`<�`<��`<� a<�a<�a<I<b<��b<ɺb<0�b<��b<��b<YYb<�b<A�a<�Fa<��`<��`<�y`<-``<�_`<y`<ܩ`<
�`<Fa<��a<�b<�`b<~�b<��b<��b<e�b<��b<p`b<�b<�a<~Ia<��`<��`<{�`<�k`<_n`</�`<��`<^a<�\a<8�a<2b<qb<�b<d�b<�b<��b<k�b<Qb<Z�a<�a<�8a<|�`<�`<�{`<+i`<p`<��`<	�`<.a<�la<$�a<z+b<b<�b<��b<U�b<)�b<8�b<�Db<`�a<��a<�+a<��`<��`< x`<�i`<u`<ݘ`<��`<_!a<E|a<��a<�9b<0�b<��b<J�b<2�b<��b<)�b<O3b<��a<�ta<a<��`<�`<p`<�e`<;u`<�`<%�`<j+a<�a<S�a<�Cb<p�b<��b<N�b<�b<��b<^ub<!b<��a<Tba<�	a<��`<��`<k`<ge`<Ey`<�`<��`<�9a<\�a<s�a<?Qb<�b<��b<B�b<�b<��b<�cb<b<��a<Ka<C�`<�`<�w`<\`<�Y`<�p`<Z�`<r�`<�7a<��a<��a<9Lb<�b<��b<��b<�b<�b<Bb<1�a<0�a<�'a<�`<8�`<�]`<�F`<�H`<�c`<ۖ`<P�`<$5a<l�a<�a<pHb<ߊb<�b<�b<n�b<Iqb<I%b<��a<�ha<�
a<J�`<&w`<CL`<x9`<f@`<$``<J�`<,�`<[;a<��a<��a< Mb<�b<��b<��b<M�b<`b<6b<��a<�Sa<��`<ۧ`<�j`<�C`<�5`<4A`<Te`<|�`<��`<�Ia<ުa<�  �  S�a<2b<	{b<2�b<r�b<��b<)pb<R0b<��a<ܛa<Wa< a<N�`<��`<��`<k�`<��`<�+a<jha<�a<��a< Eb<@�b<��b<��b<0�b<�vb<)b<��a<�Sa<<�`<t`<�`<3�_<�_<��_<Y�_<�_<KN`<��`<�(a<��a<�
b<Ceb<��b<�b<��b<\�b<�xb<�5b<��a<ޢa<cba</a<�a<��`<��`<(a<�/a<�ca<
�a<R�a<�;b<"�b<˹b<��b<��b<��b< �b<�0b<��a<�Sa<��`<�x`<�#`<��_<��_<H�_<��_<�3`<-�`<Q�`<*la<Y�a<�Db<.�b<�b<�b<�b<�b<|vb<�.b<��a<�a<�^a<e/a<�a<�a< 	a< a<gHa<�a<�a<�b<Yb<��b<��b<��b<��b<8�b<�mb<fb<�a<q,a<��`<~Y`<�`<C�_<T�_<��_<^`<OO`<��`<�a<0�a<�b<cb<x�b<2�b<	�b<��b<�b<�^b<�b<��a<��a<=Ka<� a<�a<� a<|a<	(a<bUa<U�a<�a<-#b<ukb<�b<[�b<��b<~�b<��b<�Jb<:�a<�ta<^ a<��`<�7`<~�_<}�_<]�_<Y�_<$`<Vh`<��`<�@a<N�a<�b<�xb<v�b<�b<��b<��b<9�b<>b<�a<;�a<�da<A/a<�	a<��`<��`<�a<P%a<Wa<g�a<��a<
)b<�mb<n�b<��b<��b<F�b<5jb<fb<9�a<�2a<ľ`<�U`<��_<#�_<ʦ_<��_<z�_< `<$f`<��`<^Da<(�a<Ob<!mb<��b<�b<c�b<�b<�Jb<|b<��a<Mna<<0a<� a<w�`<��`<��`<��`<�a<Oa<��a<B�a<k'b<�hb<ʘb<��b<��b<l�b<�:b<�a<dma<��`<�`<�%`<��_<H�_<v�_<ޣ_<��_<:`<�|`<v�`<_aa<�  �  ��a<� b<Vb<�b<T�b< �b<|b<�Mb<�b<L�a<ղa<V�a<�ra<da<o`a<ga<Eya<��a<��a<w�a<;(b<.^b<��b<�b<ߧb<��b<TOb<�a<тa<Ua<T|`<��_<��_<�C_<_<X_<�,_<�o_<M�_<�I`<��`<�Ta<��a<M8b<V�b<z�b<��b<Y�b<6�b<:Yb<�#b<��a<�a<�a<2�a<�a<��a<��a<��a<��a<*�a<�)b<kab<p�b<^�b<6�b<G�b<y�b<w[b<T�a<[a<�`<�v`<R�_<�_<T_<�1_<�5_<!`_<�_<�`<g�`<�a<��a<�b<Rmb<ҭb<$�b<<�b<
�b<b<3Yb<�"b<��a<��a<��a<��a<R�a<9�a<�a<��a<7�a<�b<
Bb<�xb<c�b<��b<.�b<��b<\�b<�=b<D�a<�Sa<D�`<L`<��_<�~_<#D_<�._<�?_<9v_<!�_<�=`<��`<EDa<��a<�1b<k�b<�b<��b<[�b<��b<8|b<�Eb<:b<l�a<��a<��a<b�a<:�a<O�a<Σa<��a<��a<�b<�Ob<��b<u�b<��b<��b<�b<�qb<b<(�a<"a<u�`<`<j�_<b_<�3_<"+_<�H_<��_<I�_<�b`<L�`<�ja<��a<�Kb<	�b<w�b<��b<��b<��b<�ab<�)b<��a<S�a<6�a<5�a<�a<l~a<\�a<�a<��a<��a<b<�Nb<�b<	�b<�b<�b<�b<�>b<�a<�_a<V�`<�T`<��_<Iv_<�/_<�_<S_<�9_<M�_<��_<�j`<��`<Wra<��a<:Db<<�b<�b<��b<��b<�ab<�,b<��a<!�a<{�a<�za<6ga<j_a<�aa<zoa<��a<�a<��a<�b<�Fb<~vb<��b<�b<�b<�\b<�
b<�a<o a<��`<X`<�_<�J_<H_<�^<1_<�B_<(�_<*`<|�`<�a<�  �  OSa<��a<�+b<kb<ϊb<��b<�|b<Y^b<t:b<Db<��a<��a<t�a<`�a<%�a<�a<�a<��a<�b</#b<�Fb<'kb<a�b<ޖb<3�b<�hb<�"b<��a<�@a<��`<�`<�_<�_<��^<؎^<��^<��^<��^<�`_<��_<�y`<7a<r�a<�b<*]b<��b<V�b< �b<�b<�ob<�Lb<-b<Mb<�b<p�a<��a<��a<�a<�b<�b<�3b<Ub<�yb<�b<n�b<.�b<k�b<D|b<�+b<�a<A9a<��`<,`<0�_<�_<H�^<��^<Q�^<��^<4_<��_<4`<h�`<HWa<��a<�?b<��b<v�b<ֿb<:�b< �b<�ub<�Rb<�3b<b<b<�b<	b<:b<
b<b<v)b<Eb<gb<#�b<ڪb<��b<��b<��b<fb<�
b<)�a<w	a<v`<��_<xe_<4 _<h�^<4�^<q�^<��^<BX_<�_<�d`<s�`<��a<��a<\b<�b<g�b<Ͻb<իb<�b<�hb<BFb<�)b<8b<Xb<�b< b<bb<�	b<�b<�-b<�Kb<tnb<ϑb<1�b<ۻb<c�b<��b<�Eb<��a<Cba<Y�`<�?`<m�_<�:_<��^<]�^<��^<u�^<�_<�z_<��_<S�`<v#a<C�a<�b<�nb<��b<��b<P�b<u�b<#xb<+Sb<i1b<�b<�b<q�a<��a<��a<��a<c�a<4b<*%b<eDb<\gb<��b<�b<�b<��b<�`b<�b<ҟa<�a< �`<d�_<rk_<&�^<�^<��^<��^<ڷ^<�_<��_<�`<��`</a<%�a<�b<`b<H�b<�b<وb<�lb<KIb<O%b<�b<��a<�a<c�a<
�a<��a<^�a<�a<E�a<�b<s5b<hYb<�xb<s�b<q�b<ob<S3b<��a<aa<!�`<�B`<H�_<�1_<j�^<��^<�r^<��^<~�^<_%_<��_<�2`<��`<�  �  /a<�a<�b<Kb<rrb<�~b<�wb<�eb<0Pb<r=b<�0b<{*b<)b<*b<�*b<�*b<�*b<�-b<�5b<�Db<YYb<�ob<��b<�b<0tb<�Fb<��a<َa<�a<�q`<
�_<a>_<:�^<u\^<�$^<�^<+@^<-�^<�_<��_<4`<g�`<ba<�a<|8b</ub<��b<��b<�b<�{b<�gb<�Wb<Nb<_Jb<Kb<�Lb<�Mb<zNb<�Ob<	Ub<`b<�qb<��b<7�b<.�b<m�b<֏b<WXb<b<��a<c�`<-c`<,�_<e5_<
�^<bh^<�>^<�C^<Dw^<R�^<�R_<d�_<6�`<Ya<B�a<�b<^gb<��b<�b<e�b<�b<Άb<�rb<�cb<a[b<uXb<�Xb<pYb<lYb<�Xb<Zb<�_b<lb<u~b<�b<�b<�b<8�b<_�b<�?b<��a<�^a<��`<.`<��_<�	_<�^<U^<�:^<�O^<�^<W�^<��_<�`<��`<bNa<��a<5b<{b<
�b<�b<��b<N�b<�~b<}kb<�^b<�Wb<Vb<�Vb<�Vb<Vb<JUb<�Wb<5_b<Mmb<�b<H�b<��b<�b<m�b<qjb<>b<�a<C*a<J�`<*�_<�]_<�^<�z^<B^<�7^<	\^<�^<� _<k�_<�K`<��`<�va<`�a<Jb<�b<סb<�b<M�b<'�b<�mb<�[b<@Pb<Jb<Ib<�Hb<�Gb<Fb<HEb<yHb<lQb<�`b<�tb<��b<�b<_�b<vb<=b<C�a<fma<��`<�B`<m�_<�_<z�^<D^<�^<=^<,Q^<ĭ^<�+_<��_<g]`<�`<�~a<��a<�=b<nnb<?�b<�b<�ob<Zb<IEb<�5b<�,b<S)b<U)b<_)b<�(b<(b<
)b<�.b<�:b<�Lb<Ibb<"ub<�}b<�sb<�Ob<b<ªa<�+a<N�`<��_<`_<��^<]h^<p!^<L^<g^<�^^<��^<1P_<��_<�`<�  �  ��`<Ha<��a<!4b<%`b<Jrb<'rb<hb<�[b<7Sb<[Pb<Sb<�Xb< ^b<�_b<�]b<�Xb<8Tb<[Sb<`Xb<�bb<pb<qyb<,wb<�`b</b<Z�a<<na<�`<�E`<��_<�_<B�^< ^<��]<s�]<~�]<)R^<��^<�b_<�`<&�`<??a<�a<�b<�_b<;�b<D�b<ϋb<6�b<�vb<�pb<�pb<�ub<l|b<��b<�b<d�b<�{b<�xb<.zb<��b<��b<��b<��b<��b<�zb<?b<y�a<Uia<��`<�5`<͒_<��^<~^<�%^<L�]<��]<�5^<Ӗ^<�_<\�_<Y`<��`<#�a<)�a<Ob<��b<��b<e�b<��b<k�b<�b<�b<�b<�b<͋b<юb<ݍb<�b<��b<��b<��b<N�b<y�b<=�b<�b<��b<�kb<%b<v�a<�:a<��`<��_<^_<F�^<\^<�^<R�]<;^<hQ^<w�^<~L_<��_<D�`<�)a<�a<�b<db<��b<��b<�b<Öb<P�b<K�b<~b<k�b<��b<��b<��b<S�b<��b<H~b<�|b<ـb<��b<ܖb<\�b<A�b<
�b<�Rb<b<J�a<pa<�f`<��_<d&_<�^<Q9^<,�]<&�]<W^<m^<��^<a{_<z`<W�`<Ta<@�a<H0b<�ob<]�b<��b<,�b<��b<�|b<�tb<�rb<�ub<lzb<�}b<�|b<xb<Jqb<"lb<�kb<qb<o{b<��b<L�b<��b<ab<�#b<��a<%Ka<C�`<`<q_<L�^<�Z^<�^<T�]<�]<t^<Gp^<��^<��_<21`<��`<s]a<��a<e%b<yZb<�sb<�wb<�ob<�bb<�Wb<Rb<jRb<�Vb<!\b<�^b<c]b<EXb<�Rb<]Ob<�Qb<�Yb<�eb<Vpb<�qb<Ebb<n9b<e�a<��a<�a<�n`<'�_<�*_<��^<e(^</�]<��]<��]<T^<��^<_<��_<�]`<�  �  ��`<�sa<��a<�+b<�Yb<�mb<�ob<ahb<�_b<'Zb<�Zb<�`b<ib<�ob<�qb</ob<�hb<>ab<�\b<�^b<�eb<�ob<Pvb<�qb<�Yb<�&b<�a<vba<��`<�6`<��_<��^<1k^<�^<$�]<��]<l�]<k<^<Ӹ^<�P_<�_<%�`<�2a<��a<`b<�Wb<'}b<,�b<�b<��b<Q{b<�xb<
|b<e�b<I�b<g�b<ǔb<U�b<�b<x�b<��b<��b<��b<��b<��b<��b<'sb<�5b<��a<]a<��`<�%`<#�_<	�^<�h^<^<��]<�]<�^<��^<Z_<2�_<�I`<��`<6za<��a<ZFb<s}b<#�b<�b<�b<�b<�b<?�b<��b<��b<��b<��b<m�b<��b<��b<;�b<Q�b<.�b<	�b<��b<z�b<	�b<�cb<\b<&�a<#.a<��`<E�_<�K_<��^<�E^<v�]<��]<��]<*;^<Ȫ^<�9_<#�_<��`<�a<��a<b<�[b< �b<ǜb<��b<�b<�b<=�b<Z�b<=�b<�b<)�b<؝b<��b<��b<S�b<)�b<�b<��b<q�b<?�b<�b<�}b<Jb<��a<��a<F�`<�W`<ֱ_<8_<�^<�"^<��]<]�]<C^<RW^<��^<zi_<�`<U�`<�Ga<9�a<�&b<�gb<G�b<s�b<u�b<�b<��b<�|b<E~b<��b<I�b<E�b<��b<�b<h�b<�wb<�sb<#vb<%}b<�b<k�b<�{b<qYb<�b<ͻa<�>a<w�`<W`<k__<[�^<dE^<��]<��]<��]<��]<[^<_�^<�|_<�!`<P�`<�Qa<~�a<�b<0Sb<Hnb<�tb<�nb<'eb<�]b<0[b<_b<�fb<Omb<�pb<�nb<�hb<�`b<�Yb<�Xb<�]b<Hfb<nb<kmb<�[b<\1b<��a<T�a<�`<T``<�_<2_<%�^<R^<��]<�]<�]<^<x^<y_<"�_<	O`<�  �  ��`<Ha<��a<!4b<%`b<Jrb<'rb<hb<�[b<7Sb<[Pb<Sb<�Xb< ^b<�_b<�]b<�Xb<8Tb<[Sb<`Xb<�bb<pb<qyb<,wb<�`b</b<Z�a<<na<�`<�E`<��_<�_<B�^< ^<��]<s�]<~�]<)R^<��^<�b_<�`<&�`<??a<�a<�b<�_b<;�b<D�b<ϋb<6�b<�vb<�pb<�pb<�ub<l|b<��b<�b<d�b<�{b<�xb<.zb<��b<��b<��b<��b<��b<�zb<?b<y�a<Uia<��`<�5`<͒_<��^<~^<�%^<L�]<��]<�5^<Ӗ^<�_<\�_<Y`<��`<#�a<)�a<Ob<��b<��b<e�b<��b<k�b<�b<�b<�b<�b<͋b<юb<ݍb<�b<��b<��b<��b<N�b<y�b<=�b<�b<��b<�kb<%b<v�a<�:a<��`<��_<^_<F�^<\^<�^<R�]<;^<hQ^<w�^<~L_<��_<D�`<�)a<�a<�b<db<��b<��b<�b<Öb<P�b<K�b<~b<k�b<��b<��b<��b<S�b<��b<H~b<�|b<ـb<��b<ܖb<\�b<A�b<
�b<�Rb<b<J�a<pa<�f`<��_<d&_<�^<Q9^<,�]<&�]<W^<m^<��^<a{_<z`<W�`<Ta<@�a<H0b<�ob<]�b<��b<,�b<��b<�|b<�tb<�rb<�ub<lzb<�}b<�|b<xb<Jqb<"lb<�kb<qb<o{b<��b<L�b<��b<ab<�#b<��a<%Ka<C�`<`<q_<L�^<�Z^<�^<T�]<�]<t^<Gp^<��^<��_<21`<��`<s]a<��a<e%b<yZb<�sb<�wb<�ob<�bb<�Wb<Rb<jRb<�Vb<!\b<�^b<c]b<EXb<�Rb<]Ob<�Qb<�Yb<�eb<Vpb<�qb<Ebb<n9b<e�a<��a<�a<�n`<'�_<�*_<��^<e(^</�]<��]<��]<T^<��^<_<��_<�]`<�  �  /a<�a<�b<Kb<rrb<�~b<�wb<�eb<0Pb<r=b<�0b<{*b<)b<*b<�*b<�*b<�*b<�-b<�5b<�Db<YYb<�ob<��b<�b<0tb<�Fb<��a<َa<�a<�q`<
�_<a>_<:�^<u\^<�$^<�^<+@^<-�^<�_<��_<4`<g�`<ba<�a<|8b</ub<��b<��b<�b<�{b<�gb<�Wb<Nb<_Jb<Kb<�Lb<�Mb<zNb<�Ob<	Ub<`b<�qb<��b<7�b<.�b<m�b<֏b<WXb<b<��a<c�`<-c`<,�_<e5_<
�^<bh^<�>^<�C^<Dw^<R�^<�R_<d�_<6�`<Ya<B�a<�b<^gb<��b<�b<e�b<�b<Άb<�rb<�cb<a[b<uXb<�Xb<pYb<lYb<�Xb<Zb<�_b<lb<u~b<�b<�b<�b<8�b<_�b<�?b<��a<�^a<��`<.`<��_<�	_<�^<U^<�:^<�O^<�^<W�^<��_<�`<��`<bNa<��a<5b<{b<
�b<�b<��b<N�b<�~b<}kb<�^b<�Wb<Vb<�Vb<�Vb<Vb<JUb<�Wb<5_b<Mmb<�b<H�b<��b<�b<m�b<qjb<>b<�a<C*a<J�`<*�_<�]_<�^<�z^<B^<�7^<	\^<�^<� _<k�_<�K`<��`<�va<`�a<Jb<�b<סb<�b<M�b<'�b<�mb<�[b<@Pb<Jb<Ib<�Hb<�Gb<Fb<HEb<yHb<lQb<�`b<�tb<��b<�b<_�b<vb<=b<C�a<fma<��`<�B`<m�_<�_<z�^<D^<�^<=^<,Q^<ĭ^<�+_<��_<g]`<�`<�~a<��a<�=b<nnb<?�b<�b<�ob<Zb<IEb<�5b<�,b<S)b<U)b<_)b<�(b<(b<
)b<�.b<�:b<�Lb<Ibb<"ub<�}b<�sb<�Ob<b<ªa<�+a<N�`<��_<`_<��^<]h^<p!^<L^<g^<�^^<��^<1P_<��_<�`<�  �  OSa<��a<�+b<kb<ϊb<��b<�|b<Y^b<t:b<Db<��a<��a<t�a<`�a<%�a<�a<�a<��a<�b</#b<�Fb<'kb<a�b<ޖb<3�b<�hb<�"b<��a<�@a<��`<�`<�_<�_<��^<؎^<��^<��^<��^<�`_<��_<�y`<7a<r�a<�b<*]b<��b<V�b< �b<�b<�ob<�Lb<-b<Mb<�b<p�a<��a<��a<�a<�b<�b<�3b<Ub<�yb<�b<n�b<.�b<k�b<D|b<�+b<�a<A9a<��`<,`<0�_<�_<H�^<��^<Q�^<��^<4_<��_<4`<h�`<HWa<��a<�?b<��b<v�b<ֿb<:�b< �b<�ub<�Rb<�3b<b<b<�b<	b<:b<
b<b<v)b<Eb<gb<#�b<ڪb<��b<��b<��b<fb<�
b<)�a<w	a<v`<��_<xe_<4 _<h�^<4�^<q�^<��^<BX_<�_<�d`<s�`<��a<��a<\b<�b<g�b<Ͻb<իb<�b<�hb<BFb<�)b<8b<Xb<�b< b<bb<�	b<�b<�-b<�Kb<tnb<ϑb<1�b<ۻb<c�b<��b<�Eb<��a<Cba<Y�`<�?`<m�_<�:_<��^<]�^<��^<u�^<�_<�z_<��_<S�`<v#a<C�a<�b<�nb<��b<��b<P�b<u�b<#xb<+Sb<i1b<�b<�b<q�a<��a<��a<��a<c�a<4b<*%b<eDb<\gb<��b<�b<�b<��b<�`b<�b<ҟa<�a< �`<d�_<rk_<&�^<�^<��^<��^<ڷ^<�_<��_<�`<��`</a<%�a<�b<`b<H�b<�b<وb<�lb<KIb<O%b<�b<��a<�a<c�a<
�a<��a<^�a<�a<E�a<�b<s5b<hYb<�xb<s�b<q�b<ob<S3b<��a<aa<!�`<�B`<H�_<�1_<j�^<��^<�r^<��^<~�^<_%_<��_<�2`<��`<�  �  ��a<� b<Vb<�b<T�b< �b<|b<�Mb<�b<L�a<ղa<V�a<�ra<da<o`a<ga<Eya<��a<��a<w�a<;(b<.^b<��b<�b<ߧb<��b<TOb<�a<тa<Ua<T|`<��_<��_<�C_<_<X_<�,_<�o_<M�_<�I`<��`<�Ta<��a<M8b<V�b<z�b<��b<Y�b<6�b<:Yb<�#b<��a<�a<�a<2�a<�a<��a<��a<��a<��a<*�a<�)b<kab<p�b<^�b<6�b<G�b<y�b<w[b<T�a<[a<�`<�v`<R�_<�_<T_<�1_<�5_<!`_<�_<�`<g�`<�a<��a<�b<Rmb<ҭb<$�b<<�b<
�b<b<3Yb<�"b<��a<��a<��a<��a<R�a<9�a<�a<��a<7�a<�b<
Bb<�xb<c�b<��b<.�b<��b<\�b<�=b<D�a<�Sa<D�`<L`<��_<�~_<#D_<�._<�?_<9v_<!�_<�=`<��`<EDa<��a<�1b<k�b<�b<��b<[�b<��b<8|b<�Eb<:b<l�a<��a<��a<b�a<:�a<O�a<Σa<��a<��a<�b<�Ob<��b<u�b<��b<��b<�b<�qb<b<(�a<"a<u�`<`<j�_<b_<�3_<"+_<�H_<��_<I�_<�b`<L�`<�ja<��a<�Kb<	�b<w�b<��b<��b<��b<�ab<�)b<��a<S�a<6�a<5�a<�a<l~a<\�a<�a<��a<��a<b<�Nb<�b<	�b<�b<�b<�b<�>b<�a<�_a<V�`<�T`<��_<Iv_<�/_<�_<S_<�9_<M�_<��_<�j`<��`<Wra<��a<:Db<<�b<�b<��b<��b<�ab<�,b<��a<!�a<{�a<�za<6ga<j_a<�aa<zoa<��a<�a<��a<�b<�Fb<~vb<��b<�b<�b<�\b<�
b<�a<o a<��`<X`<�_<�J_<H_<�^<1_<�B_<(�_<*`<|�`<�a<�  �  S�a<2b<	{b<2�b<r�b<��b<)pb<R0b<��a<ܛa<Wa< a<N�`<��`<��`<k�`<��`<�+a<jha<�a<��a< Eb<@�b<��b<��b<0�b<�vb<)b<��a<�Sa<<�`<t`<�`<3�_<�_<��_<Y�_<�_<KN`<��`<�(a<��a<�
b<Ceb<��b<�b<��b<\�b<�xb<�5b<��a<ޢa<cba</a<�a<��`<��`<(a<�/a<�ca<
�a<R�a<�;b<"�b<˹b<��b<��b<��b< �b<�0b<��a<�Sa<��`<�x`<�#`<��_<��_<H�_<��_<�3`<-�`<Q�`<*la<Y�a<�Db<.�b<�b<�b<�b<�b<|vb<�.b<��a<�a<�^a<e/a<�a<�a< 	a< a<gHa<�a<�a<�b<Yb<��b<��b<��b<��b<8�b<�mb<fb<�a<q,a<��`<~Y`<�`<C�_<T�_<��_<^`<OO`<��`<�a<0�a<�b<cb<x�b<2�b<	�b<��b<�b<�^b<�b<��a<��a<=Ka<� a<�a<� a<|a<	(a<bUa<U�a<�a<-#b<ukb<�b<[�b<��b<~�b<��b<�Jb<:�a<�ta<^ a<��`<�7`<~�_<}�_<]�_<Y�_<$`<Vh`<��`<�@a<N�a<�b<�xb<v�b<�b<��b<��b<9�b<>b<�a<;�a<�da<A/a<�	a<��`<��`<�a<P%a<Wa<g�a<��a<
)b<�mb<n�b<��b<��b<F�b<5jb<fb<9�a<�2a<ľ`<�U`<��_<#�_<ʦ_<��_<z�_< `<$f`<��`<^Da<(�a<Ob<!mb<��b<�b<c�b<�b<�Jb<|b<��a<Mna<<0a<� a<w�`<��`<��`<��`<�a<Oa<��a<B�a<k'b<�hb<ʘb<��b<��b<l�b<�:b<�a<dma<��`<�`<�%`<��_<H�_<v�_<ޣ_<��_<:`<�|`<v�`<_aa<�  �  Kb<@Yb<Z�b<E�b<��b<l�b<VVb<�b<s�a<�Fa<��`<۟`<Qf`<�C`<<:`<LJ`<�r`<��`<�a<�_a<(�a<�b<�kb<$�b<W�b<۷b<.�b<vSb<��a<סa<2Ba<'�`< `<_k`<|M`<�H`<8]`<�`<��`<� a<�a<�a<I<b<��b<ɺb<0�b<��b<��b<YYb<�b<A�a<�Fa<��`<��`<�y`<-``<�_`<y`<ܩ`<
�`<Fa<��a<�b<�`b<~�b<��b<��b<e�b<��b<p`b<�b<�a<~Ia<��`<��`<{�`<�k`<_n`</�`<��`<^a<�\a<8�a<2b<qb<�b<d�b<�b<��b<k�b<Qb<Z�a<�a<�8a<|�`<�`<�{`<+i`<p`<��`<	�`<.a<�la<$�a<z+b<b<�b<��b<U�b<)�b<8�b<�Db<`�a<��a<�+a<��`<��`< x`<�i`<u`<ݘ`<��`<_!a<E|a<��a<�9b<0�b<��b<J�b<2�b<��b<)�b<O3b<��a<�ta<a<��`<�`<p`<�e`<;u`<�`<%�`<j+a<�a<S�a<�Cb<p�b<��b<N�b<�b<��b<^ub<!b<��a<Tba<�	a<��`<��`<k`<ge`<Ey`<�`<��`<�9a<\�a<s�a<?Qb<�b<��b<B�b<�b<��b<�cb<b<��a<Ka<C�`<�`<�w`<\`<�Y`<�p`<Z�`<r�`<�7a<��a<��a<9Lb<�b<��b<��b<�b<�b<Bb<1�a<0�a<�'a<�`<8�`<�]`<�F`<�H`<�c`<ۖ`<P�`<$5a<l�a<�a<pHb<ߊb<�b<�b<n�b<Iqb<I%b<��a<�ha<�
a<J�`<&w`<CL`<x9`<f@`<$``<J�`<,�`<[;a<��a<��a< Mb<�b<��b<��b<M�b<`b<6b<��a<�Sa<��`<ۧ`<�j`<�C`<�5`<4A`<Te`<|�`<��`<�Ia<ުa<�  �  �2b<1rb<��b<t�b<�b<bxb<f.b<��a<�\a<`�`<�y`<�`<;�_<F�_<�_<�_<}�_<=0`<C�`<�a<�za<l�a<)Gb<��b<;�b<��b<��b<
pb<{.b<��a<ɚa<*Xa<
"a<{�`<6�`<��`<��`<za<�Ca<ׂa< �a<qb<�`b<l�b<�b<b�b< �b<~b<[,b<��a<Ta<L�`<�w`<X `<��_<��_<I�_<��_<�`<�t`<��`<FSa<��a<2b<��b<��b<p�b<I�b<'�b<ۂb<#=b<�a<P�a<�ia<�7a<3a<�a<�a<�a<�@a<�ua<��a<Yb<Lb<p�b<��b<|�b<+�b< �b<$yb<�b<�a<>a<@�`<�f`<$`<�_<��_<�_<�_<�@`<�`<�a<V�a<��a<kUb<��b<��b<A�b<Y�b<��b<mb<S$b<�a<��a<CWa<�*a<�a<na<�a<A&a<Qa<Ίa<�a<�b<9db<.�b<t�b<}�b<{�b<��b<0]b<X�a<�a<a<�`<�G`<��_<;�_<z�_<��_<�`<�Y`<�`<�-a<�a<�b<�lb<��b<�b<��b<5�b<�b<�Ob<Lb<�a<�wa<Aa<�a<�a<��`<a<�-a<�]a<��a<��a<�.b<�ub<�b<��b<~�b<o�b<��b<�6b<B�a<�Za<��`<
z`<� `<��_<Ӽ_<�_<Z�_<�`<h`<1�`<�Ba<��a<zb<rb<��b<��b<ɿb<%�b<pdb<jb<�a<S�a<�Fa<a<��`<��`<��`<_�`<a<�Na<!�a<��a<�#b<�fb<�b<�b<>�b<��b<Nb<��a<Ӆa<%a<`<�8`<��_<�_<h�_<�_<��_<@`<.m`<��`<�Na<�a<�#b<ypb<��b<��b<m�b<Nwb<�9b<��a<$�a<�^a<#a<B�`<q�`<L�`<��`<��`<�a<�Wa<��a<��a<�  �  Ob<@}b<��b<��b<.�b<�Rb<��a<_�a<a<o�`<(`<ɗ_<�B_<G_<��^<|_<bT_<��_<}%`<��`<�.a<3�a<&b<�hb<�b<��b<S�b<�~b<�Nb<
b<��a<c�a<.�a<|a<�oa<Bna<-wa<Ƌa<īa<��a<�	b<~Ab<�vb<p�b<}�b<նb<ɕb<�Tb<7�a<�a<��`<fz`<d�_<Ș_<�N_<w'_<w&_<�K_<��_<{�_<�u`<��`<$�a<v�a<�]b<E�b<��b<e�b<��b</�b<db<�-b<��a<��a<��a<k�a<��a<ޑa<x�a<ϴa<9�a<b<%8b<�nb<�b<��b<��b<��b<�b<iKb<��a<�ga<��`<P_`<��_<B�_<!J_<�._<g9_<j_<U�_<�)`<Ĩ`<�.a<T�a<)"b<�{b< �b<C�b<��b<�b<f�b<�Qb<�b<�a<��a<�a<��a<2�a<��a<8�a<e�a<�a<^b<�Jb<��b<J�b<$�b<��b<ƹb<�b<Q+b<��a<;a<�`<a4`<��_<�n_<:_<+_<(B_<c~_<��_<N`<x�`<�Ua<R�a<y=b<W�b<��b<��b<��b<��b<-pb<�9b<
b<��a<0�a<s�a<g�a<>�a<V�a<�a<��a<��a<�!b<Xb<�b<��b<]�b<��b< �b<�`b<� b<��a<a<�~`<�`<��_<�L_<Z#_<4 _<SC_<��_<��_<Ig`<,�`<wna<��a<#Gb<�b<Ȱb<۶b<��b<�xb<IDb<�b<��a<֬a<��a<�ua<�ka<la<.wa<�a<"�a<��a<[b<rFb<bwb<�b<R�b<�b<�mb<s b<@�a<�;a<�`<�1`<�_<�[_<_<*�^<�	_<�9_<��_<��_<�w`<8�`<�~a<G�a<�Ib<��b<��b<��b<��b<�Sb<b<��a<޶a<L�a<�ra<�aa<�[a<�`a<rpa<��a<}�a<��a<�b<�  �  �^b<F}b<b�b<��b<�hb<�'b<��a<sMa<��`<-`<͞_<O"_<��^<χ^<8w^<$�^<��^<�=_<,�_<qQ`<C�`<�oa<��a<@b<rzb<��b<ԕb<��b<|bb<?b<b<�b<_�a<��a<��a<��a<��a<j�a<��a<Ob<~8b<#]b<�b<ɜb<`�b<��b<qb<�&b<ؽa<=a<��`<=`<~�_<d_<�^<��^<a�^<f�^<�_<#�_<E`<W�`<�;a<��a<�.b<�~b<o�b<�b<y�b<��b<�}b<Zb<o:b<"b<�b<Gb<Vb<�b<-	b<�b<v%b<|?b<B`b<�b<�b<�b<޽b<�b<Lpb<b<��a<�a<�`<l�_<�w_<[_<O�^<�^<Y�^<-�^<oE_<��_<�L`<��`<oa<=�a<�Ob<o�b<,�b<(�b<j�b<`�b<�qb<�Nb<31b<�b<�b<kb<	b<�b<@b<-b<�-b<WJb<�lb<g�b<Z�b<�b<��b<;�b<Wb<��a<�{a<��`<�Z`<��_<O_<��^<��^<f�^<��^<e _<+g_<��_<y`<a<ؕa<b<~db<1�b<��b<<�b<ƣb<��b<�_b<<>b<2#b<gb<�b<��a<��a<!b<�
b<'b<s1b<ePb<�sb<5�b<X�b<J�b<��b<yb<3b<d�a<�Ea<�`<�`<Δ_<�_<'�^<��^<�^< �^<l_<�_<�`<��`<)a<D�a<b<^fb<z�b<y�b<b�b<2�b<�]b<9b<Yb<�a<��a<��a<�a<��a<��a<��a<[�a<	b<y8b<�[b<a|b<��b<��b<�|b<�Eb<8�a<"|a<t�`<6``<!�_<�I_<��^<_�^<�v^<��^<��^<�_<��_<�`<B�`<s=a<Z�a<�b<�ab<p�b<�b<b<�ab<�=b<�b<��a<%�a<3�a<��a<��a<��a<a�a<��a<��a<�b<�:b<�  �  Yeb<wb<!~b<�pb<FHb<� b<w�a<�a<.�`<H�_<�J_<��^<�]^<^<�^<)^<�r^<��^<tn_<
`<��`<;a<�a</b<�[b<�~b<ćb<�~b<&lb<MWb<�Eb<�:b<6b<�5b<37b<8b<�8b<$9b<f=b<6Gb<�Wb<mb<`�b<N�b<�b<J�b<VNb<��a<Ќa<�a<�j`<�_<Z;_<&�^<"e^<5^<�3^<�`^<��^<�3_<��_<ne`<xa<�a<:b<[b<R�b<̫b<ܭb<��b<�b<�wb<�gb<$^b<BZb<(Zb<�Zb<>Zb<OYb<�Yb<e^b<
ib<4zb<M�b<�b<�b<��b<��b<-Kb<$�a<�sa<,�`<�F`<��_<>_<V�^<�\^<�:^<5H^<f�^<�^<�j_<�`<�`<�7a<�a<�'b<Nsb<��b<�b<k�b<��b<�b<|qb<�cb<#\b<�Yb<cZb<�Zb<DZb<oYb<[b<�ab<�nb<��b<��b<��b<��b<�b<�wb<�/b<.�a<&Ea<�`<�`<�w_<��^<̉^<�I^<7^<�S^<��^<�_<˖_<�1`<��`<aa<>�a<�>b<qb<��b<$�b<��b<\�b<�wb<fb<�Zb<Ub<,Tb<�Tb<&Ub<�Tb<wTb<�Wb<c`b<�ob<��b<��b<�b< �b<�b<�\b<r	b<a�a<:a<Uq`<u�_<�=_<V�^<-c^<�0^<Q-^<mX^<8�^<M'_<3�_<�T`<��`<Pza<��a<�Bb<Xxb<3�b<��b<�b<Clb<�Vb<~Eb<;b<R6b<z5b<05b<_4b<�2b<�2b<G7b<�Ab<kRb<.gb<�zb<�b<p~b<�^b<� b<N�a<IHa<(�`<�`<}_<q�^<�{^<�-^<�^<s^<BS^<��^<�9_<��_<�n`<�a<�a<��a<�@b<�lb<�|b<xb<�fb<Qb<D=b<//b<�'b<;%b<�%b<$&b<&b<|%b<�'b<�.b<<b<qOb<�  �  Mgb<rqb<=qb<E^b<1b<,�a<�ya<��`<�V`<�_<l_<܈^<�^<s�]<��]<�]<3^<��^<b9_<��_<�~`<Ta<1�a<��a<xEb<Amb<H|b<ozb<pb<�db<\]b<\b<�_b<Ffb<�kb<cmb<kb<Efb<�bb<�bb<dib<$ub<��b<�b<:�b<lb<�5b<�a<hka<��`<J>`<��_<�_<f�^<:#^<��]<@�]<�^<|z^<��^<�_<F8`<%�`<�la<��a<Bb<�}b<X�b<��b<ܞb<�b<@�b<U�b<O�b<��b<Q�b<��b<�b<z�b<v�b<��b<��b<��b<?�b<z�b<(�b<�b<�rb<1b<��a<�Pa<��`<`<Qv_<��^<	k^<�^<i�]<[^<>B^<]�^<Z3_<��_<�t`<�a<��a<�b<�[b<|�b<^�b<��b<��b<C�b<��b<��b<K�b<v�b<��b<�b<+�b<Ĉb<9�b<̀b<�b<�b<��b<��b<֡b<[�b<�`b<Ob<P�a<2 a<��`<\�_<zA_<y�^<I^<^<��]<p^<�\^<��^<�a_<n`<s�`<?=a<T�a<$b<"ib<>�b<��b<2�b<J�b<\�b<�}b<�{b<�~b<��b<��b<w�b<^�b<��b<�|b<,|b<[�b<��b<��b<~�b<0�b<I|b<3Db<��a<�ua<��`<�D`<�_<5_<��^<E!^<��]<��]<3^<�o^<6�^<1�_<�'`<o�`<XXa<k�a<�)b<�cb<��b<��b<N�b<>sb<0gb<0`b<4_b<�bb<�gb<djb<4ib<db<�]b<nYb<&Zb<�`b<"lb<wb<Nzb<�mb<	Ib<�b<�a<(%a<��`<��_<#I_<$�^<�<^<��]<�]<��]<#^<�y^<�_<��_<�C`<\�`<�ja<��a<4)b<�Yb<Cob<'qb<�gb<>[b<UQb<Mb<�Nb<�Sb<DYb<�[b<�Yb<�Tb<�Ob<�Mb<:Qb<�Zb<�  �  4b<�8b<�3b<Zb<��a<��a<�ea<q�`<Չ`<!`<D�_<�4_<��^<#�^<_�^<ֽ^<H�^<�K_<K�_<�.`<�`<a<3�a<��a<a
b<.b<�?b<�Bb<D>b<h6b<k/b<+b<�)b<�*b<$,b<?-b<F-b<�-b<r/b<4b<�;b< Eb<vMb<#Pb<*Gb<�-b<��a<պa<�`a<J�`<�~`<[`<�_< 7_<�^<��^<��^<��^<I3_<��_<�`<�|`<�`<4ea<C�a<�b<�>b<�[b<)hb<�gb<Mab<Yb<sRb<xNb<�Mb<�Mb<�Nb<,Nb<3Mb<�Lb<;Nb<�Rb<�Yb<Hbb<hb<tfb<9Wb<X6b<��a<U�a<�Pa<��`<�f`<��_<U�_<~*_<"�^<:�^<s�^<�_<Y_<ν_<�1`<߫`<�!a<"�a<��a<�"b<Mb<�cb<�jb<?gb<:_b<Wb<$Qb<6Nb<�Mb<JNb<�Nb<5Nb<�Mb<�Mb<�Ob<aUb<B]b<Teb<.ib<�cb<�Nb<�&b<;�a<��a<,a<	�`<�<`<��_<�`_<_<�^<��^<��^<U_<At_<��_<�U`<-�`<kAa<פa<h�a<�-b<�Pb<�ab<7db<�^b<qVb<�Nb<�Ib<'Hb<1Hb<�Hb<PIb<{Hb<Hb<�Hb<2Lb<qRb<�Zb<�ab<�bb<9Xb<+=b<}b<��a<�ja<[�`<Ȅ`<z
`<
�_<17_<��^<��^<��^<��^<)_<��_<��_<�l`<�`<cQa<��a<P�a<�%b<wAb<1Lb<�Jb<�Bb<D9b<�1b<�,b<�*b<H*b<T*b<e)b<�'b<''b< (b<,b<�2b<�:b<B@b<1>b<�.b<&b<��a<�a<&a<~�`<�:`<t�_<JU_<��^<�^<��^<��^<w�^<g)_<Ӎ_<�`<M{`<��`<Za<r�a<6�a<b<[1b<8b<y4b<9,b<�#b<�b<�b<ab<�b<�b<b<�b<b<�b<�#b<�+b<�  �  3b<E9b<�5b<F#b<�a<^�a<�ma<?a<I�`<4`<�_<�C_<��^<��^<n�^<��^<O_<�Z_<��_<:`<�`<�$a<�a<��a<Bb<�1b<qAb<�Bb<]<b<U2b<�(b<G"b<�b< b<�b<�b<c b<"b<�%b<,b<p6b<SBb<�Lb<+Qb<Jb<2b<Pb< �a<�ha<t�`<��`<�`<2�_<�F_<�_<��^<��^<R _<C_<+�_<�`<�`<a�`<gma<��a<8b<@Cb<_b<^ib<]gb<�^b</Tb<Kb<�Db<�Ab<�@b<�@b<�@b<�@b<�Ab<<Eb<Lb<�Ub<7`b<�gb<	hb<�Zb<;b<�b<�a<SYa<��`<r`<��_<�_<y:_<��^<H�^<[�^<_<\h_<��_<$>`<��`<�*a<�a<��a<(b<Qb<fb<+kb<fb<\b<sQb<Ib<�Cb<�Ab<3Ab<\Ab<Ab<JAb<Cb<�Gb<�Ob<�Yb<�cb<�ib<�eb<�Rb<�+b<��a<��a<�4a<�`<�H`<<�_<�o_<I!_<��^<��^<E�^<`/_<(�_<+�_<ia`<+�`<�Ia<��a<��a<v2b<4Tb<Ncb<6db<�\b<^Rb<hHb< Ab<=b<�;b<�;b<�;b<�;b<J<b<�>b<�Db<QMb<�Wb<�`b<�cb<"[b<wAb<�b<��a<�ra<�a<Ϗ`<`<M�_<�F_<� _<��^<��^</�^<�8_<��_<b`<�w`<h�`<�Ya<��a<��a<O*b<�Db<gMb<Jb<7@b<d4b<A*b< #b<6b<yb<�b<�b<Jb<�b<b<]%b<�.b<�8b<@b<�?b<�1b<�b<��a<��a<�.a<9�`<)F`<}�_<	d_<�_<��^<÷^<k�^<��^<�8_<��_<�`<�`<��`<�aa<8�a<h�a<b<�3b<�8b<>3b<)b<Bb<�b<�b<Pb<�b<b<�b<lb<�b<�b<�b<�(b<�  �  .b<>:b<�;b<�-b<Vb<n�a<q�a<F!a<β`<;?`<0�_<4o_<c$_<��^<��^<��^</4_<K�_<��_<�\`<��`<�=a<�a<��a<�b<@;b<]Fb<�Bb<�5b<%b<�b<�b<�a<�a<��a<(�a<��a<��a<�b<�b</&b<�8b<�Ib<�Sb<�Qb<�=b<�b<f�a<;�a<a<ɩ`<Q7`<��_<As_<(2_<�_<_<�/_<�o_<P�_<_4`<��`<pa<�a<c�a<&"b<�Ob<*gb<�lb<eb<Vb<�Db<�4b<�(b<Y b<�b<�b<�b<+b<>!b<5*b<<7b<�Gb<�Xb<gb<plb<�cb<0Hb<wb<��a<�qa<�a<Ǔ`<�!`<5�_<h_<�/_<}_<!_<�K_<$�_<n�_<�a`<��`<FEa<t�a<�a<�6b<�[b<�lb<�lb<�ab<Qb<�?b<�0b<�%b<�b< b<�b<�b<�b<O$b<�.b<�<b<Nb<�^b<�jb<�kb<']b<C:b<� b<��a<�Na<	�`<l`<��_<"�_<�O_<m!_<�_<x(_<J]_<��_<�`<��`<��`<ca<��a<�b<�?b<�]b<?hb<�cb<�Vb< Eb<b4b<�&b<;b<�b<�b<4b<b<=b<�!b<�-b<=b<iNb<�]b<yfb<�bb<JMb<�"b<;�a<3�a<"a<�`<n;`<��_<Qs_<,0_<�_<�_<�'_<�e_<%�_<:&`<w�`<x	a<Pqa<��a<�
b<�6b<�Lb<�Pb<�Gb<�7b<�$b<b<�b<��a<F�a<^�a<��a<��a<u�a<�b<�b<� b<�1b<'?b<(Db<;b<�b<��a<E�a<(Ga<D�`<�g`<c�_<�_<w:_<�_<��^<�^<�_<td_<l�_<V1`<��`<la<Uxa<��a<b<*b<^:b<5:b<�.b<b<zb<h�a<d�a<h�a<��a<b�a<|�a<�a<��a<x�a<;b<�b<�  �  �#b<9b<�Bb<u;b<�b<��a<��a<YHa<��`<�t`<2`<Ͳ_<m_<�B_<7_<�J_<9|_<��_<Y&`<F�`<��`<;ca<��a<� b<�/b<kGb<rKb<�?b<�)b<�b<��a<i�a<��a<��a<��a<2�a<B�a<;�a<	�a<��a<#b<�'b<�Bb<hUb<�Zb<�Mb<D+b<i�a<��a<WCa<��`<zo`<+`<ڸ_<�|_<�\_<6\_<�z_<+�_<T	`<_m`<��`<�Ea<J�a<�a<99b<`b<�pb<ob<_b<QFb<�*b<=b<��a<b�a<��a<��a<�a<'�a<��a<��a< b<0b<�Kb<cb<�pb<5ob<CZb<�.b<��a<ϖa<@2a<��`<�\`<��_<��_<n{_<�d_<�m_<��_<w�_<;1`<�`<a<ma<Q�a<�b<�Kb<jjb<tb<^lb<�Xb<�=b<2"b<�b<�a<~�a<��a<��a<��a<��a<��a<Vb<Vb<�9b<�Tb<Sib<{rb<�jb<Nb< b<��a<va<�a<��`<�9`<��_<��_<�m_<�a_<kt_<e�_<��_<N`<J�`<#a<��a<G�a<�$b<�Rb<�ib<Zmb<�`b<7Jb<�.b<`b<?�a<��a<A�a<g�a<8�a<l�a<r�a<8�a<�b<�!b<�=b<�Vb<hb<�kb<(]b<�8b<:�a<��a<cKa<�`<�s`<B`<�_<�z_<�X_<V_<�r_<�_<*�_<<_`<��`<�3a<�a<r�a<�!b<0Gb<�Vb<"Sb<�Ab<�'b<�
b<j�a<�a<��a<2�a<��a<Z�a<ߺa<7�a<Y�a<^�a<�b<$b<%;b<fHb<rFb<1b<b<2�a<�ka<�a<��`<0`<��_<�_<GM_<\6_<�>_<"f_<��_<2`<�g`<��`<A<a<3�a<��a<b<�8b<�Ab<�9b<�%b<b<�a<S�a<��a< �a<F�a<S�a<Ҩa<$�a<;�a<?�a<��a<�b<�  �  9b<�2b<�Fb<dHb<T4b<�	b<��a<�va<�a<�`<�Y`<7`<)�_<�_<��_<�_<��_<	`<�p`<b�`<�2a<��a<��a<	b<�Bb<�Rb<kMb<7b<1b<f�a<s�a<'�a<�a<poa<qda<(ca<_ka<�}a<��a<��a<�a<	b<5b<�Rb<
bb<Q]b<�Bb<�b<��a<�ta<�a<W�`<�[`<�`</�_<�_<q�_<��_<`<�Y`<U�`<>a<xa<t�a<zb<�Qb<{pb<>yb<�mb<�Rb<�-b<b<X�a<��a<��a<A�a<��a<��a<�a<R�a<��a<�a<Lb<�5b<*Yb<�qb<yyb<rlb<*Ib<�b<%�a<&ga<�a<ѥ`<gO`<.
`<~�_<y�_<\�_<��_<�.`<�~`<��`<u=a<��a<��a<�3b<]ab<.xb<@yb<Qgb<-Hb< !b<�a<j�a<	�a<Řa<��a<E�a<c�a<C�a<n�a<��a<��a<ub<�Bb<cb<�vb<�wb<Acb<8b<��a<x�a<Fa<�`<�`<B4`<��_<*�_<�_<��_<� `<�C`<`�`<z�`<Ya<�a<�b<@b<�eb<1ub<[ob<XXb<�5b<tb<��a<��a<O�a<�a<9�a<%a<��a<��a<��a<��a<��a<�#b<"Ib<[eb<sb<�lb<?Pb<�b<��a<�|a<�a<p�`<�]`<`<0�_<�_<Z�_<��_<�`<�M`<5�`</a<*fa<��a<�b<G:b<�Wb<�^b<�Qb<c5b<=b<b�a<��a<��a<}a<�ia<�`a<�`a<�ja<�~a<Úa<l�a<A�a<_b<I1b<:Ib<�Pb<'Cb<Xb<��a<4�a<�;a<��`<'y`<1"`<r�_<F�_<Θ_<I�_<r�_<�_<�N`<K�`<�a<�ka<d�a<Ob<�/b<KFb<Gb<�4b<�b<'�a<�a<=�a<�}a<{ea<[Va<#Qa<pUa<�ca<{a<Úa<.�a<E�a<�  �  �a<f%b<GDb<8Pb<�Eb<E$b<��a<2�a<�Ta<=�`<=�`<Mh`<�2`<�`<�	`<�`<�>`<�x`<^�`<�a<�ka<~�a<xb<�4b<�Qb<,Xb<xHb<�&b<��a<��a<ϊa<?Xa<I.a< a<u�`<��`<	a<�"a<�Ia<cza<��a<��a<Eb<Ib<cb<whb<Wb</b<�a<`�a<�Ua<�a<t�`<\t`<DF`<].`<.`<�E`<~s`<��`<�a<�Wa<��a<��a<�:b<�fb<�|b<a{b<eb<G>b<�b<Y�a<˝a<(ma<Fa<�+a<�a<3 a<�/a<+Ma<�va<̨a<��a<b<�Gb<zkb< ~b<�zb<�`b<�0b<��a<؞a<�Ia<Z�`<�`<�p`<�H`<p7`<Q>`<~\`<'�`<��`<%%a<�za<W�a<~b<�Ob<�sb<�b<�wb<[b<j/b<<�a<C�a<�a<2_a<�;a<�%a<�a<9$a<�8a<4Za<Նa<R�a<�a<�(b<�Ub<tb<�b<�tb<�Rb<�b<��a<݁a<2,a<��`<k�`<�^`<�=`< 4`<�B`<�g`<��`<N�`< =a< �a<!�a<U&b<�Xb<1ub<�zb<qjb<CHb<�b<��a<@�a<wa<uLa<�-a<5a<�a<-$a<
=a<�ba<]�a<p�a<��a<N3b<�[b<�sb<�wb<�db<�:b<�a<d�a<�[a<�a<��`<ht`<ED`<R*`<�'`<p=`<Xi`<Ч`<��`<�Ga<�a< �a<$%b<�Ob<�cb<�`b<%Ib<!b<R�a<��a<}a<pKa<t#a<7a<��`<��`<�
a<o'a<VPa<,�a<�a<��a<�b< Cb<*Ub<lQb<�6b<b<��a<@sa<�a<��`<�~`<�B`<K`<�`<,`<�,`<S``<��`<��`<Ja<u�a<_�a<(b<Bb<<Ob<�Eb<�(b<��a<u�a<O�a<�Ya<,a<�a<��`<��`<]�`<�a<�'a<�Ta<ĉa<��a<�  �  A�a<�b<v9b<Pb<�Ob<;8b<&b<%�a<�a<Ga<Aa<��`<[�`<��`<~`<��`<
�`<��`<Ta<|Za<,�a<��a<Zb<=Fb<�Yb<�Ub<3;b<�b<�a<��a<OFa<7a<5�`<��`<��`<�`<�`<�`<��`<6/a<�ua<s�a< b<�6b<�[b<�kb<Fdb<�Fb<�b<��a<ݓa<FNa<�a<g�`<l�`<M�`<>�`<��`<��`<�a<?Pa<��a<��a<�b<�Sb</ub<�b<;ub<�Sb<� b<@�a<
�a<5Ta<|a<-�`<�`<ȭ`<�`<��`<��`<�!a<�ba</�a<��a<�,b<�\b<[zb<��b<Dqb<)Lb<�b<��a<��a<�Ga<�
a<��`<�`<�`<��`<��`<��`<d,a<�na<׵a<��a<`7b<�db<�~b<�b<'nb<�Eb<b<��a<΂a<�>a<"a<��`<��`<��`<B�`<F�`<��`<�6a<0za<-�a<�b<"?b<8ib<ub<�~b<�fb<J;b<��a<}�a<#ta<�0a<��`<�`<ð`<Ψ`<��`<}�`<�a<^=a<āa<��a<Wb<LCb<kjb<}b<jxb<7]b</b<��a<��a<�ea<$a<[�`<u�`<V�`<ԧ`<��`<��`<�	a<%Ga<f�a<��a<b<*Ib<�lb<{b<�qb<{Rb<� b<��a<�a<YRa<a<q�`<k�`<A�`<'�`<k�`<��`<�a<$Ba<{�a<��a<b<>b<�]b<>hb<�Zb<8b<Mb<��a<gza<3a<��`<��`<��`<��`<F�`<��`<�`<��`<�;a<"�a<0�a<b<�4b<{Qb<&Xb<TGb<�!b<��a<#�a<�`a<a<n�`<�`<��`</}`<�`<^�`<�`<8�`<B>a<,�a<��a<@b<Q3b<'Mb<JPb<<b<�b<��a<;�a<�Oa<�a<�`<��`<��`<�y`<�`<��`<��`<a<�Ha<�a<�  �  �a<�a<&b<�Fb<YPb<�Cb<L$b<��a<��a<�a<�Ta<�(a<a<��`<-�`<��`<�a<4a<�ba<�a<��a<b<�2b<BOb<Xb<Jb<j%b<�a<��a<�Pa<��`<�`<�i`<)8`< `<}`<�*`<U`<��`<��`<j3a<Y�a< �a<�b<�Kb<�eb<�hb<�Ub<.2b<�b<��a<S�a<Rda<a<a<� a<�a<�a<�!a<�=a<�fa<��a<��a<�	b<�<b<db<�zb<|b<Sfb<D:b<��a<��a<OYa<a<ܸ`<bz`<�N`<y9`<<`<2V`<K�`<#�`<�a<�ka<�a<
b<�Eb<�mb<�~b<1yb<F_b<�5b<�b<��a<�a<�da<�?a<�'a<a<e!a<�3a<eSa<�~a<^�a<,�a<� b<�Ob<Qqb<��b<�yb<�[b<P(b<1�a<��a<==a<��`<n�`<�i`<BE`<�7`<yB`<<d`<ƚ`<��`<3a<Q�a<��a<4 b<�Ub<�ub<Eb<1rb<wRb<�$b<7�a<�a<��a<#Ua<�3a<�a<�a<�"a<@9a<�\a<�a<e�a<2�a<�,b<�Wb<�sb<�{b<�lb<yGb<zb<��a<�pa<ma<��`<�`<�U`<�8`<_3`<�E`<o`<��`<n�`<Ja<��a<��a<;.b<�\b<�tb<vb<�ab<<b<�	b<��a<b�a<`fa<i<a<�a<�a<�a<�a<�3a<�Za<܊a<��a<��a<)b<�Nb<|cb<9cb<�Kb<wb<��a<8�a<�9a<[�`<9�`<�W`<f+`<{`<y`<1`<�``<��`<�`<�Da<��a<$�a<�b<�Db<gUb<2Ob<�4b<�
b<�a<��a<ga<?7a<�a<�`<2�`<�`<	a<r#a<sNa<�a<y�a<��a<�b<�?b<Ob<�Gb<�)b<�a<ða<�_a<u
a<׷`<to`<�6`<O`<�`<�`<�1`<�h`<��`<�a<OWa<�  �  <za<��a<�b<�5b<Ib<�Fb<d2b<�b<��a<D�a<��a<�|a<fa<�Xa<�Ua<�[a<�ka<�a<i�a<��a<|�a<b<N>b<Pb<�Nb<;7b< 	b<��a<�qa<�a<ر`<.V`<`<7�_<�_<��_<)�_<5�_<�6`<ˎ`<��`<jRa<ܭa<��a<�4b<�Wb<�db<�\b<aDb<u!b<��a<c�a<��a<'�a<G�a<?xa<�xa<�a<ܖa<i�a<��a<� b<�*b<_Pb<�kb<�wb<Gob<lPb<pb<��a<xa<.a<��`<!^`<v`<��_<��_<��_<s�_<e#`<p`<$�`<_,a<N�a<d�a<|(b<�Yb<Jtb<�xb<�ib<iLb<&b<:�a<��a<n�a<�a<C�a<��a<>�a<��a<��a<��a<>�a<�b<T=b<`_b<�ub<ezb<�ib<�Bb<b<��a<�Xa<�`<�`<�C`<	`<W�_<��_<�_<��_<,;`<��`<��`<1Ma<ƪa<��a<�;b< eb<�wb<[ub<�`b<x?b<_b<f�a<O�a<
�a<�a<a�a<�a<�a<��a<�a<��a<e�a<,b<�Db<gcb<]tb<rb<
Zb<+b<��a<K�a<�2a<I�`<�t`<6&`<��_<��_<~�_<!�_<8	`<�O`<��`<�a<�ga<��a<Db<�Eb<gb<%rb<Jhb<;Nb<j)b<��a<o�a<��a<-�a<Da<1ta<�ra<�za<��a<I�a<��a<��a<�b<�<b<nVb<�`b<�Vb<6b<��a<��a<�Ya<��`<�`<�<`<��_<G�_<ť_<$�_<L�_<��_<�I`<��`<Pa<�da<l�a< b<�0b<�Jb<�Nb<?b</!b<K�a<��a<�a<�a<�la<�[a<�Ta<�Va<�ba<�xa<��a<��a<B�a<fb<@.b<RDb<�Hb<8b<�b<��a<9�a<O&a<[�`<Me`<`<"�_<|�_<�_<��_<o�_<	`<�[`<+�`<>a<�  �  RLa<�a<o�a<}!b<�<b<(Cb<*9b<�#b<�b<z�a<��a<{�a<�a<��a<ƪa<u�a<�a<o�a<��a<7�a<�b<�.b<�Bb<LJb<O@b<,!b<��a<ڞa<�Aa<��`<�m`<8`<O�_<�p_<_K_<;E_<f^_<�_<��_<:F`<��`<"a<�a<��a<b<)Fb<�Zb<X\b<�Nb<�7b<%b<b<��a<S�a<��a<��a<��a<��a<�a<��a<�	b<�%b<iBb<\b<�lb<ob<g^b<�7b<r�a<�a<�Da<��`<$o`<�`<�_<C�_<dg_<�j_<>�_<��_<!`<م`<_�`<N[a<��a<m	b<�Bb<Ceb<rb<�lb<�Zb<�@b<%b<b<��a<+�a<~�a<��a<H�a<��a<��a<|b< b<�5b<Qb<agb<sb<�nb<UVb< 'b<E�a<��a<F"a<J�`<OM`<��_<N�_<�v_<,e_<�r_<]�_<*�_<�A`<��`<~a<�|a<#�a<b<�Pb<}kb<�qb<`gb<�Qb<y6b<�b<�b<��a<�a<�a<��a<��a<��a<{�a<b<�b<e:b<�Tb<�gb<�nb<�cb<Db<�b<I�a<Tba<�`<#�`< '`<i�_<��_< h_<a_<Vy_<	�_<p�_<	^`</�`<j3a<��a<K�a<�+b<WUb<[hb<hb<�Xb<�?b<'#b<b<��a<X�a<��a<��a<��a<��a<��a<��a<��a<�b<�0b<lHb<TWb<�Wb<�Eb<Jb<��a<��a<z&a<i�`<�N`<f�_<��_<	`_<vC_</F_<h_<�_<��_<>_`<P�`<�3a<a<��a<�b<�;b<Hb<EBb<|/b<�b<��a<��a<�a<�a<߭a<��a<۪a<ѱa<��a<-�a<v�a<�b< b<A6b<�Ab<==b<�$b<6�a<'�a<[Va<��`<��`<�`<�_<{s_<�C_<�2_<{@_<m_<.�_<�`<Sx`<��`<�  �  �%a<Q�a<��a<�b<D/b<�<b<�:b<�.b<�b<�b<��a<}�a<j�a<]�a<��a<��a<��a<��a<Mb<b<&&b<?7b<�Bb<cBb<�1b<�b<��a<�}a<[a<��`<�6`<�_<�l_<�&_<��^<��^<�_<�M_<]�_<�`<=`<��`<�^a<M�a<b<|4b<�Ob<�Xb<bSb<�Eb<F5b<�%b<�b< b<�b<zb<mb<�b<�b<. b<�-b<�>b<�Qb<�ab<�ib<�db<jMb< b<v�a<t�a<Za<j�`<�5`<��_<�u_<8_<_<�_<�B_<l�_<�_<N`<��`<[2a<��a<��a<�,b<�Ub<uib<�kb<Ubb<YRb<�@b<k1b<�%b<cb<Wb<�b<ub<�b<�"b<w,b<i:b<hKb<�\b<�ib<�mb<3bb<3Cb<�b<A�a<�ba<��`<�`<e`<<�_<�]_<�*_<�_<�&_<tV_<ڢ_<�`<�t`<�`<Va<c�a<5b<�<b<0^b<qkb<ib<�\b<?Kb<�9b<`+b<� b<tb<�b<�b<b<�b<�!b<�,b<�;b<�Lb<C]b<�gb<�fb<%Ub<�.b<��a<�a<!:a<�`<OV`<��_<Ǌ_<D_<>_<�_<�-_<�g_<G�_<�#`<Ε`<8a<�ra<��a<�b<�Cb<X]b<1db<4]b<�Mb<F;b<�)b<�b<b<�b<kb<Vb<�b<pb<b<�b<�.b<�?b<�Mb<fTb<�Mb<�4b<�b<��a<afa<�`<�`< `<�_<S_<�_<0�^<=�^<�_<�`_<��_<�'`<��`<�
a<�pa<<�a<�b<3,b<R?b<+Ab<�6b<h&b<?b<Kb<>�a<0�a<��a<��a<��a<��a<|�a< �a<�	b<�b<�+b<�8b<M<b<�0b<�b<��a<,�a<i0a<+�`<�O`<��_<|z_<(+_<��^<
�^<5�^<?$_<�p_<Q�_<PC`<>�`<�  �  �a<�qa<��a<��a< %b<#7b<(:b<4b<�)b<�b<�b<�b<�b<�b<ub<�b<�b<rb<Ob<g%b<�0b<:;b<�@b<�;b<Q&b<��a<�a<ga<��`<��`<(`<
�_<�@_<��^<��^<��^<�^< _<�y_<T�_<�]`<+�`<SFa<�a<x�a<�'b<Gb<kTb<�Tb<�Mb<�Cb<;b<H5b<�2b<�2b<�3b<�4b<�5b<�7b<)<b<�Cb<Nb<�Yb<}cb<Ffb<�\b<�@b<�b<o�a<|ka<�`<~�`<�`<)�_<hH_<q_<�^<��^<�_<Z_<��_<�)`<ˡ`<a<��a<��a<�b<*Jb<,bb<�ib<�eb<6\b<tQb<�Hb<'Cb<�@b<@b<V@b<F@b<�@b<2Bb<�Fb<Nb<FXb<�bb<�ib<hhb<bXb<z5b<\�a<��a<VIa<��`<�_`<��_<x�_<�/_<>�^<f�^<-�^<(_<�w_<��_<�Q`<��`<I<a<��a<Y�a<�.b<�Sb<�eb<ehb<�ab<ZWb<�Lb<�Db< @b<�=b<�=b<�=b<=b<�=b<�?b<�Db<Mb<�Wb<Gab<�eb<`b<�Ib<�b<�a<�a<\a<ɪ`<�2`<��_<�^_<"_<u�^<{�^<��^<o:_<h�_<�_<`t`<g�`<*Za<C�a<Bb<�6b<Tb<`b<k^b<oUb<�Ib<?b<O7b<�2b<�0b<�/b<�.b<�-b<�-b<0b<�5b<>b<Hb<�Ob<�Pb<cEb<3(b<��a<��a<mNa<��`<h`<�_<��_<&_<A�^<�^<W�^<��^<m4_<��_<[`<�z`<��`<�Ya<�a<��a<� b<8b<�>b<L:b<=0b<�$b<�b<pb<sb<`b<5b<�b<�b<b<&b<�b<�'b<�1b<�8b<7b<�&b<�b<~�a<�za<a<e�`<4-`<�_<�O_< �^<��^<Գ^<��^<��^<�E_<@�_<� `<��`<�  �  a<�ia<&�a<r�a<"!b<�4b<�9b<�5b<b-b<�%b<C b<%b<:b<b< b<�b<�b<� b<9$b<�*b<�3b<X<b<�?b<9b<2"b<��a<�a<_a<��`<�`<�`< �_<^1_<��^<�^<��^<��^<�_<�j_<_�_<bR`<��`<�=a<d�a<��a<�"b<�Cb<�Rb<�Tb<�Ob<'Hb<�Ab<c>b<>b<??b<Ab<JBb<�Bb<hCb<�Eb<�Jb<�Rb<J\b<�cb<�db<FYb<h<b<M
b<�a<:ca<��`<5|`<�`<��_<�8_<��^<��^<��^<Z_<�J_<|�_<y`<ٖ`<�a<�ya<��a<<b<�Eb<d_b<�hb<�fb<_b<�Vb<tPb<Mb<�Lb<Mb<�Mb<�Mb<�Lb<Mb< Ob<gTb<5\b<�db<�ib<|fb<�Tb<�0b<�a<9�a<�@a<��`<�S`<l�_<s_<�_<z�^<R�^<Z�^<�_<�h_<K�_<�E`<s�`<�3a<ؙa<��a<�)b<Pb<�cb<hb<cb<�Zb<�Rb<)Mb<�Jb<OJb<�Jb<!Kb<)Jb<�Ib<�Ib<�Lb<�Rb<�Zb<hbb<=eb<y]b<�Eb<�b<D�a<|�a<^a<
�`<I&`<�_<rO_<�_<��^<o�^<e�^<�*_<��_<!�_<�h`<��`<�Qa<��a<`�a<2b<Qb<�^b<�^b<�Wb<%Nb<�Eb<j@b<>b<:=b<=b<3<b<m:b<H9b<j9b<�<b<�Bb<pJb<QPb<�Ob<*Bb<�#b<�a<Z�a<,Fa<N�`<�\`<4�_<s_<1_<��^<�^<d�^<?�^<�$_<[�_<��_<�o`<m�`<�Qa<��a<1�a<Xb<85b<�=b<0;b<3b<*b<H#b<Ub<Xb<Pb<�b<b<$b<�b<�b<�#b<n+b<�3b<�8b<-5b<+#b<��a<*�a<,sa<ya<I�`<h!`<Ȫ_<�@_<�^<Ѷ^<Ţ^<��^<��^<�6_<��_<�`<��`<�  �  �a<�qa<��a<��a< %b<#7b<(:b<4b<�)b<�b<�b<�b<�b<�b<ub<�b<�b<rb<Ob<g%b<�0b<:;b<�@b<�;b<Q&b<��a<�a<ga<��`<��`<(`<
�_<�@_<��^<��^<��^<�^< _<�y_<T�_<�]`<+�`<SFa<�a<x�a<�'b<Gb<kTb<�Tb<�Mb<�Cb<;b<H5b<�2b<�2b<�3b<�4b<�5b<�7b<)<b<�Cb<Nb<�Yb<}cb<Ffb<�\b<�@b<�b<o�a<|ka<�`<~�`<�`<)�_<hH_<q_<�^<��^<�_<Z_<��_<�)`<ˡ`<a<��a<��a<�b<*Jb<,bb<�ib<�eb<6\b<tQb<�Hb<'Cb<�@b<@b<V@b<F@b<�@b<2Bb<�Fb<Nb<FXb<�bb<�ib<hhb<bXb<z5b<\�a<��a<VIa<��`<�_`<��_<x�_<�/_<>�^<f�^<-�^<(_<�w_<��_<�Q`<��`<I<a<��a<Y�a<�.b<�Sb<�eb<ehb<�ab<ZWb<�Lb<�Db< @b<�=b<�=b<�=b<=b<�=b<�?b<�Db<Mb<�Wb<Gab<�eb<`b<�Ib<�b<�a<�a<\a<ɪ`<�2`<��_<�^_<"_<u�^<{�^<��^<o:_<h�_<�_<`t`<g�`<*Za<C�a<Bb<�6b<Tb<`b<k^b<oUb<�Ib<?b<O7b<�2b<�0b<�/b<�.b<�-b<�-b<0b<�5b<>b<Hb<�Ob<�Pb<cEb<3(b<��a<��a<mNa<��`<h`<�_<��_<&_<A�^<�^<W�^<��^<m4_<��_<[`<�z`<��`<�Ya<�a<��a<� b<8b<�>b<L:b<=0b<�$b<�b<pb<sb<`b<5b<�b<�b<b<&b<�b<�'b<�1b<�8b<7b<�&b<�b<~�a<�za<a<e�`<4-`<�_<�O_< �^<��^<Գ^<��^<��^<�E_<@�_<� `<��`<�  �  �%a<Q�a<��a<�b<D/b<�<b<�:b<�.b<�b<�b<��a<}�a<j�a<]�a<��a<��a<��a<��a<Mb<b<&&b<?7b<�Bb<cBb<�1b<�b<��a<�}a<[a<��`<�6`<�_<�l_<�&_<��^<��^<�_<�M_<]�_<�`<=`<��`<�^a<M�a<b<|4b<�Ob<�Xb<bSb<�Eb<F5b<�%b<�b< b<�b<zb<mb<�b<�b<. b<�-b<�>b<�Qb<�ab<�ib<�db<jMb< b<v�a<t�a<Za<j�`<�5`<��_<�u_<8_<_<�_<�B_<l�_<�_<N`<��`<[2a<��a<��a<�,b<�Ub<uib<�kb<Ubb<YRb<�@b<k1b<�%b<cb<Wb<�b<ub<�b<�"b<w,b<i:b<hKb<�\b<�ib<�mb<3bb<3Cb<�b<A�a<�ba<��`<�`<e`<<�_<�]_<�*_<�_<�&_<tV_<ڢ_<�`<�t`<�`<Va<c�a<5b<�<b<0^b<qkb<ib<�\b<?Kb<�9b<`+b<� b<tb<�b<�b<b<�b<�!b<�,b<�;b<�Lb<C]b<�gb<�fb<%Ub<�.b<��a<�a<!:a<�`<OV`<��_<Ǌ_<D_<>_<�_<�-_<�g_<G�_<�#`<Ε`<8a<�ra<��a<�b<�Cb<X]b<1db<4]b<�Mb<F;b<�)b<�b<b<�b<kb<Vb<�b<pb<b<�b<�.b<�?b<�Mb<fTb<�Mb<�4b<�b<��a<afa<�`<�`< `<�_<S_<�_<0�^<=�^<�_<�`_<��_<�'`<��`<�
a<�pa<<�a<�b<3,b<R?b<+Ab<�6b<h&b<?b<Kb<>�a<0�a<��a<��a<��a<��a<|�a< �a<�	b<�b<�+b<�8b<M<b<�0b<�b<��a<,�a<i0a<+�`<�O`<��_<|z_<(+_<��^<
�^<5�^<?$_<�p_<Q�_<PC`<>�`<�  �  RLa<�a<o�a<}!b<�<b<(Cb<*9b<�#b<�b<z�a<��a<{�a<�a<��a<ƪa<u�a<�a<o�a<��a<7�a<�b<�.b<�Bb<LJb<O@b<,!b<��a<ڞa<�Aa<��`<�m`<8`<O�_<�p_<_K_<;E_<f^_<�_<��_<:F`<��`<"a<�a<��a<b<)Fb<�Zb<X\b<�Nb<�7b<%b<b<��a<S�a<��a<��a<��a<��a<�a<��a<�	b<�%b<iBb<\b<�lb<ob<g^b<�7b<r�a<�a<�Da<��`<$o`<�`<�_<C�_<dg_<�j_<>�_<��_<!`<م`<_�`<N[a<��a<m	b<�Bb<Ceb<rb<�lb<�Zb<�@b<%b<b<��a<+�a<~�a<��a<H�a<��a<��a<|b< b<�5b<Qb<agb<sb<�nb<UVb< 'b<E�a<��a<F"a<J�`<OM`<��_<N�_<�v_<,e_<�r_<]�_<*�_<�A`<��`<~a<�|a<#�a<b<�Pb<}kb<�qb<`gb<�Qb<y6b<�b<�b<��a<�a<�a<��a<��a<��a<{�a<b<�b<e:b<�Tb<�gb<�nb<�cb<Db<�b<I�a<Tba<�`<#�`< '`<i�_<��_< h_<a_<Vy_<	�_<p�_<	^`</�`<j3a<��a<K�a<�+b<WUb<[hb<hb<�Xb<�?b<'#b<b<��a<X�a<��a<��a<��a<��a<��a<��a<��a<�b<�0b<lHb<TWb<�Wb<�Eb<Jb<��a<��a<z&a<i�`<�N`<f�_<��_<	`_<vC_</F_<h_<�_<��_<>_`<P�`<�3a<a<��a<�b<�;b<Hb<EBb<|/b<�b<��a<��a<�a<�a<߭a<��a<۪a<ѱa<��a<-�a<v�a<�b< b<A6b<�Ab<==b<�$b<6�a<'�a<[Va<��`<��`<�`<�_<{s_<�C_<�2_<{@_<m_<.�_<�`<Sx`<��`<�  �  <za<��a<�b<�5b<Ib<�Fb<d2b<�b<��a<D�a<��a<�|a<fa<�Xa<�Ua<�[a<�ka<�a<i�a<��a<|�a<b<N>b<Pb<�Nb<;7b< 	b<��a<�qa<�a<ر`<.V`<`<7�_<�_<��_<)�_<5�_<�6`<ˎ`<��`<jRa<ܭa<��a<�4b<�Wb<�db<�\b<aDb<u!b<��a<c�a<��a<'�a<G�a<?xa<�xa<�a<ܖa<i�a<��a<� b<�*b<_Pb<�kb<�wb<Gob<lPb<pb<��a<xa<.a<��`<!^`<v`<��_<��_<��_<s�_<e#`<p`<$�`<_,a<N�a<d�a<|(b<�Yb<Jtb<�xb<�ib<iLb<&b<:�a<��a<n�a<�a<C�a<��a<>�a<��a<��a<��a<>�a<�b<T=b<`_b<�ub<ezb<�ib<�Bb<b<��a<�Xa<�`<�`<�C`<	`<W�_<��_<�_<��_<,;`<��`<��`<1Ma<ƪa<��a<�;b< eb<�wb<[ub<�`b<x?b<_b<f�a<O�a<
�a<�a<a�a<�a<�a<��a<�a<��a<e�a<,b<�Db<gcb<]tb<rb<
Zb<+b<��a<K�a<�2a<I�`<�t`<6&`<��_<��_<~�_<!�_<8	`<�O`<��`<�a<�ga<��a<Db<�Eb<gb<%rb<Jhb<;Nb<j)b<��a<o�a<��a<-�a<Da<1ta<�ra<�za<��a<I�a<��a<��a<�b<�<b<nVb<�`b<�Vb<6b<��a<��a<�Ya<��`<�`<�<`<��_<G�_<ť_<$�_<L�_<��_<�I`<��`<Pa<�da<l�a< b<�0b<�Jb<�Nb<?b</!b<K�a<��a<�a<�a<�la<�[a<�Ta<�Va<�ba<�xa<��a<��a<B�a<fb<@.b<RDb<�Hb<8b<�b<��a<9�a<O&a<[�`<Me`<`<"�_<|�_<�_<��_<o�_<	`<�[`<+�`<>a<�  �  �a<�a<&b<�Fb<YPb<�Cb<L$b<��a<��a<�a<�Ta<�(a<a<��`<-�`<��`<�a<4a<�ba<�a<��a<b<�2b<BOb<Xb<Jb<j%b<�a<��a<�Pa<��`<�`<�i`<)8`< `<}`<�*`<U`<��`<��`<j3a<Y�a< �a<�b<�Kb<�eb<�hb<�Ub<.2b<�b<��a<S�a<Rda<a<a<� a<�a<�a<�!a<�=a<�fa<��a<��a<�	b<�<b<db<�zb<|b<Sfb<D:b<��a<��a<OYa<a<ܸ`<bz`<�N`<y9`<<`<2V`<K�`<#�`<�a<�ka<�a<
b<�Eb<�mb<�~b<1yb<F_b<�5b<�b<��a<�a<�da<�?a<�'a<a<e!a<�3a<eSa<�~a<^�a<,�a<� b<�Ob<Qqb<��b<�yb<�[b<P(b<1�a<��a<==a<��`<n�`<�i`<BE`<�7`<yB`<<d`<ƚ`<��`<3a<Q�a<��a<4 b<�Ub<�ub<Eb<1rb<wRb<�$b<7�a<�a<��a<#Ua<�3a<�a<�a<�"a<@9a<�\a<�a<e�a<2�a<�,b<�Wb<�sb<�{b<�lb<yGb<zb<��a<�pa<ma<��`<�`<�U`<�8`<_3`<�E`<o`<��`<n�`<Ja<��a<��a<;.b<�\b<�tb<vb<�ab<<b<�	b<��a<b�a<`fa<i<a<�a<�a<�a<�a<�3a<�Za<܊a<��a<��a<)b<�Nb<|cb<9cb<�Kb<wb<��a<8�a<�9a<[�`<9�`<�W`<f+`<{`<y`<1`<�``<��`<�`<�Da<��a<$�a<�b<�Db<gUb<2Ob<�4b<�
b<�a<��a<ga<?7a<�a<�`<2�`<�`<	a<r#a<sNa<�a<y�a<��a<�b<�?b<Ob<�Gb<�)b<�a<ða<�_a<u
a<׷`<to`<�6`<O`<�`<�`<�1`<�h`<��`<�a<OWa<�  �  A�a<�b<v9b<Pb<�Ob<;8b<&b<%�a<�a<Ga<Aa<��`<[�`<��`<~`<��`<
�`<��`<Ta<|Za<,�a<��a<Zb<=Fb<�Yb<�Ub<3;b<�b<�a<��a<OFa<7a<5�`<��`<��`<�`<�`<�`<��`<6/a<�ua<s�a< b<�6b<�[b<�kb<Fdb<�Fb<�b<��a<ݓa<FNa<�a<g�`<l�`<M�`<>�`<��`<��`<�a<?Pa<��a<��a<�b<�Sb</ub<�b<;ub<�Sb<� b<@�a<
�a<5Ta<|a<-�`<�`<ȭ`<�`<��`<��`<�!a<�ba</�a<��a<�,b<�\b<[zb<��b<Dqb<)Lb<�b<��a<��a<�Ga<�
a<��`<�`<�`<��`<��`<��`<d,a<�na<׵a<��a<`7b<�db<�~b<�b<'nb<�Eb<b<��a<΂a<�>a<"a<��`<��`<��`<B�`<F�`<��`<�6a<0za<-�a<�b<"?b<8ib<ub<�~b<�fb<J;b<��a<}�a<#ta<�0a<��`<�`<ð`<Ψ`<��`<}�`<�a<^=a<āa<��a<Wb<LCb<kjb<}b<jxb<7]b</b<��a<��a<�ea<$a<[�`<u�`<V�`<ԧ`<��`<��`<�	a<%Ga<f�a<��a<b<*Ib<�lb<{b<�qb<{Rb<� b<��a<�a<YRa<a<q�`<k�`<A�`<'�`<k�`<��`<�a<$Ba<{�a<��a<b<>b<�]b<>hb<�Zb<8b<Mb<��a<gza<3a<��`<��`<��`<��`<F�`<��`<�`<��`<�;a<"�a<0�a<b<�4b<{Qb<&Xb<TGb<�!b<��a<#�a<�`a<a<n�`<�`<��`</}`<�`<^�`<�`<8�`<B>a<,�a<��a<@b<Q3b<'Mb<JPb<<b<�b<��a<;�a<�Oa<�a<�`<��`<��`<�y`<�`<��`<��`<a<�Ha<�a<�  �  �a<f%b<GDb<8Pb<�Eb<E$b<��a<2�a<�Ta<=�`<=�`<Mh`<�2`<�`<�	`<�`<�>`<�x`<^�`<�a<�ka<~�a<xb<�4b<�Qb<,Xb<xHb<�&b<��a<��a<ϊa<?Xa<I.a< a<u�`<��`<	a<�"a<�Ia<cza<��a<��a<Eb<Ib<cb<whb<Wb</b<�a<`�a<�Ua<�a<t�`<\t`<DF`<].`<.`<�E`<~s`<��`<�a<�Wa<��a<��a<�:b<�fb<�|b<a{b<eb<G>b<�b<Y�a<˝a<(ma<Fa<�+a<�a<3 a<�/a<+Ma<�va<̨a<��a<b<�Gb<zkb< ~b<�zb<�`b<�0b<��a<؞a<�Ia<Z�`<�`<�p`<�H`<p7`<Q>`<~\`<'�`<��`<%%a<�za<W�a<~b<�Ob<�sb<�b<�wb<[b<j/b<<�a<C�a<�a<2_a<�;a<�%a<�a<9$a<�8a<4Za<Նa<R�a<�a<�(b<�Ub<tb<�b<�tb<�Rb<�b<��a<݁a<2,a<��`<k�`<�^`<�=`< 4`<�B`<�g`<��`<N�`< =a< �a<!�a<U&b<�Xb<1ub<�zb<qjb<CHb<�b<��a<@�a<wa<uLa<�-a<5a<�a<-$a<
=a<�ba<]�a<p�a<��a<N3b<�[b<�sb<�wb<�db<�:b<�a<d�a<�[a<�a<��`<ht`<ED`<R*`<�'`<p=`<Xi`<Ч`<��`<�Ga<�a< �a<$%b<�Ob<�cb<�`b<%Ib<!b<R�a<��a<}a<pKa<t#a<7a<��`<��`<�
a<o'a<VPa<,�a<�a<��a<�b< Cb<*Ub<lQb<�6b<b<��a<@sa<�a<��`<�~`<�B`<K`<�`<,`<�,`<S``<��`<��`<Ja<u�a<_�a<(b<Bb<<Ob<�Eb<�(b<��a<u�a<O�a<�Ya<,a<�a<��`<��`<]�`<�a<�'a<�Ta<ĉa<��a<�  �  9b<�2b<�Fb<dHb<T4b<�	b<��a<�va<�a<�`<�Y`<7`<)�_<�_<��_<�_<��_<	`<�p`<b�`<�2a<��a<��a<	b<�Bb<�Rb<kMb<7b<1b<f�a<s�a<'�a<�a<poa<qda<(ca<_ka<�}a<��a<��a<�a<	b<5b<�Rb<
bb<Q]b<�Bb<�b<��a<�ta<�a<W�`<�[`<�`</�_<�_<q�_<��_<`<�Y`<U�`<>a<xa<t�a<zb<�Qb<{pb<>yb<�mb<�Rb<�-b<b<X�a<��a<��a<A�a<��a<��a<�a<R�a<��a<�a<Lb<�5b<*Yb<�qb<yyb<rlb<*Ib<�b<%�a<&ga<�a<ѥ`<gO`<.
`<~�_<y�_<\�_<��_<�.`<�~`<��`<u=a<��a<��a<�3b<]ab<.xb<@yb<Qgb<-Hb< !b<�a<j�a<	�a<Řa<��a<E�a<c�a<C�a<n�a<��a<��a<ub<�Bb<cb<�vb<�wb<Acb<8b<��a<x�a<Fa<�`<�`<B4`<��_<*�_<�_<��_<� `<�C`<`�`<z�`<Ya<�a<�b<@b<�eb<1ub<[ob<XXb<�5b<tb<��a<��a<O�a<�a<9�a<%a<��a<��a<��a<��a<��a<�#b<"Ib<[eb<sb<�lb<?Pb<�b<��a<�|a<�a<p�`<�]`<`<0�_<�_<Z�_<��_<�`<�M`<5�`</a<*fa<��a<�b<G:b<�Wb<�^b<�Qb<c5b<=b<b�a<��a<��a<}a<�ia<�`a<�`a<�ja<�~a<Úa<l�a<A�a<_b<I1b<:Ib<�Pb<'Cb<Xb<��a<4�a<�;a<��`<'y`<1"`<r�_<F�_<Θ_<I�_<r�_<�_<�N`<K�`<�a<�ka<d�a<Ob<�/b<KFb<Gb<�4b<�b<'�a<�a<=�a<�}a<{ea<[Va<#Qa<pUa<�ca<{a<Úa<.�a<E�a<�  �  �#b<9b<�Bb<u;b<�b<��a<��a<YHa<��`<�t`<2`<Ͳ_<m_<�B_<7_<�J_<9|_<��_<Y&`<F�`<��`<;ca<��a<� b<�/b<kGb<rKb<�?b<�)b<�b<��a<i�a<��a<��a<��a<2�a<B�a<;�a<	�a<��a<#b<�'b<�Bb<hUb<�Zb<�Mb<D+b<i�a<��a<WCa<��`<zo`<+`<ڸ_<�|_<�\_<6\_<�z_<+�_<T	`<_m`<��`<�Ea<J�a<�a<99b<`b<�pb<ob<_b<QFb<�*b<=b<��a<b�a<��a<��a<�a<'�a<��a<��a< b<0b<�Kb<cb<�pb<5ob<CZb<�.b<��a<ϖa<@2a<��`<�\`<��_<��_<n{_<�d_<�m_<��_<w�_<;1`<�`<a<ma<Q�a<�b<�Kb<jjb<tb<^lb<�Xb<�=b<2"b<�b<�a<~�a<��a<��a<��a<��a<��a<Vb<Vb<�9b<�Tb<Sib<{rb<�jb<Nb< b<��a<va<�a<��`<�9`<��_<��_<�m_<�a_<kt_<e�_<��_<N`<J�`<#a<��a<G�a<�$b<�Rb<�ib<Zmb<�`b<7Jb<�.b<`b<?�a<��a<A�a<g�a<8�a<l�a<r�a<8�a<�b<�!b<�=b<�Vb<hb<�kb<(]b<�8b<:�a<��a<cKa<�`<�s`<B`<�_<�z_<�X_<V_<�r_<�_<*�_<<_`<��`<�3a<�a<r�a<�!b<0Gb<�Vb<"Sb<�Ab<�'b<�
b<j�a<�a<��a<2�a<��a<Z�a<ߺa<7�a<Y�a<^�a<�b<$b<%;b<fHb<rFb<1b<b<2�a<�ka<�a<��`<0`<��_<�_<GM_<\6_<�>_<"f_<��_<2`<�g`<��`<A<a<3�a<��a<b<�8b<�Ab<�9b<�%b<b<�a<S�a<��a< �a<F�a<S�a<Ҩa<$�a<;�a<?�a<��a<�b<�  �  .b<>:b<�;b<�-b<Vb<n�a<q�a<F!a<β`<;?`<0�_<4o_<c$_<��^<��^<��^</4_<K�_<��_<�\`<��`<�=a<�a<��a<�b<@;b<]Fb<�Bb<�5b<%b<�b<�b<�a<�a<��a<(�a<��a<��a<�b<�b</&b<�8b<�Ib<�Sb<�Qb<�=b<�b<f�a<;�a<a<ɩ`<Q7`<��_<As_<(2_<�_<_<�/_<�o_<P�_<_4`<��`<pa<�a<c�a<&"b<�Ob<*gb<�lb<eb<Vb<�Db<�4b<�(b<Y b<�b<�b<�b<+b<>!b<5*b<<7b<�Gb<�Xb<gb<plb<�cb<0Hb<wb<��a<�qa<�a<Ǔ`<�!`<5�_<h_<�/_<}_<!_<�K_<$�_<n�_<�a`<��`<FEa<t�a<�a<�6b<�[b<�lb<�lb<�ab<Qb<�?b<�0b<�%b<�b< b<�b<�b<�b<O$b<�.b<�<b<Nb<�^b<�jb<�kb<']b<C:b<� b<��a<�Na<	�`<l`<��_<"�_<�O_<m!_<�_<x(_<J]_<��_<�`<��`<��`<ca<��a<�b<�?b<�]b<?hb<�cb<�Vb< Eb<b4b<�&b<;b<�b<�b<4b<b<=b<�!b<�-b<=b<iNb<�]b<yfb<�bb<JMb<�"b<;�a<3�a<"a<�`<n;`<��_<Qs_<,0_<�_<�_<�'_<�e_<%�_<:&`<w�`<x	a<Pqa<��a<�
b<�6b<�Lb<�Pb<�Gb<�7b<�$b<b<�b<��a<F�a<^�a<��a<��a<u�a<�b<�b<� b<�1b<'?b<(Db<;b<�b<��a<E�a<(Ga<D�`<�g`<c�_<�_<w:_<�_<��^<�^<�_<td_<l�_<V1`<��`<la<Uxa<��a<b<*b<^:b<5:b<�.b<b<zb<h�a<d�a<h�a<��a<b�a<|�a<�a<��a<x�a<;b<�b<�  �  3b<E9b<�5b<F#b<�a<^�a<�ma<?a<I�`<4`<�_<�C_<��^<��^<n�^<��^<O_<�Z_<��_<:`<�`<�$a<�a<��a<Bb<�1b<qAb<�Bb<]<b<U2b<�(b<G"b<�b< b<�b<�b<c b<"b<�%b<,b<p6b<SBb<�Lb<+Qb<Jb<2b<Pb< �a<�ha<t�`<��`<�`<2�_<�F_<�_<��^<��^<R _<C_<+�_<�`<�`<a�`<gma<��a<8b<@Cb<_b<^ib<]gb<�^b</Tb<Kb<�Db<�Ab<�@b<�@b<�@b<�@b<�Ab<<Eb<Lb<�Ub<7`b<�gb<	hb<�Zb<;b<�b<�a<SYa<��`<r`<��_<�_<y:_<��^<H�^<[�^<_<\h_<��_<$>`<��`<�*a<�a<��a<(b<Qb<fb<+kb<fb<\b<sQb<Ib<�Cb<�Ab<3Ab<\Ab<Ab<JAb<Cb<�Gb<�Ob<�Yb<�cb<�ib<�eb<�Rb<�+b<��a<��a<�4a<�`<�H`<<�_<�o_<I!_<��^<��^<E�^<`/_<(�_<+�_<ia`<+�`<�Ia<��a<��a<v2b<4Tb<Ncb<6db<�\b<^Rb<hHb< Ab<=b<�;b<�;b<�;b<�;b<J<b<�>b<�Db<QMb<�Wb<�`b<�cb<"[b<wAb<�b<��a<�ra<�a<Ϗ`<`<M�_<�F_<� _<��^<��^</�^<�8_<��_<b`<�w`<h�`<�Ya<��a<��a<O*b<�Db<gMb<Jb<7@b<d4b<A*b< #b<6b<yb<�b<�b<Jb<�b<b<]%b<�.b<�8b<@b<�?b<�1b<�b<��a<��a<�.a<9�`<)F`<}�_<	d_<�_<��^<÷^<k�^<��^<�8_<��_<�`<�`<��`<�aa<8�a<h�a<b<�3b<�8b<>3b<)b<Bb<�b<�b<Pb<�b<b<�b<lb<�b<�b<�b<�(b<�  �  �b<H
b<�b<y�a<�a<&�a<�`a<.a<|�`<�b`<�`<��_<_<�f_<�\_<m_<2�_<|�_<�"`<zz`<��`<�*a<Yva<^�a<��a<C b<Mb<�b<�b<�
b<b<n�a<��a<�a<'�a<��a<f�a<��a<�a<�b<�b<�b<�b<� b<�b<Db<?�a<��a<Yca<a<R�`<Ic`<x`<��_<+�_<�_<��_<��_<;�_<`<�b`<u�`<ya<�ia<d�a<��a<b<�+b<�7b<9b<�3b<�+b<4$b<gb<�b<b<b<b<[b<mb<bb<r%b<p-b<R5b<q9b<�6b<�(b<�b<W�a<��a<�[a<�a<�`<qV`<G`<w�_<X�_<�_<'�_<��_<Q�_<�2`<��`<<�`<�8a<�a<[�a<n�a<�b<�3b<�:b<�9b<�2b<Z*b<�"b<hb<�b<$b<�b<�b<�b<`b<N!b<�(b<�0b<�7b<�9b<�3b<&!b<Z b<��a<�a<#@a<�`<�`<@9`<#�_<s�_<֐_<��_<�_<��_<2�_<�I`<ɠ`<W�`<�Oa<x�a<��a<7b<E"b<�1b<b5b<�1b<*b<�!b<�b<$b<�b<b<�b<�b<Bb<Zb<�b<%b<y-b<3b<�2b<)(b<�b<3�a<�a<�la<�a<�`<g`<_`<��_<)�_<}_<�z_<�_<h�_<Z`<+U`<��`</a<�Va<��a< �a<�a<rb<�b<�b<lb<Ob<�b<��a<e�a<��a<��a<P�a<�a<��a<�a<��a<&b<�b<Bb<�b<c b<Y�a<6�a<�{a<�1a<��`<��`<�*`<��_<��_<o_< \_<�b_<p�_<l�_<y`<X`<m�`<�a<�Wa<��a<��a<��a<Cb<U	b<�b<� b<(�a<w�a<�a<3�a<��a<d�a<��a<�a<��a<�a<��a<Y b<�  �  �b<�	b<5b<��a<k�a<��a<-fa<ea<�`<�k`<�`<��_<q�_<�r_<i_</y_<ˡ_<D�_<�,`<��`<��`<�0a<�{a<y�a<��a<*b<�b<�b<�b<!b<��a<h�a<\�a<��a<4�a<��a<��a<�a<��a<� b<Ub<Fb<:b< b<(b<�b<��a<~�a<ia<�a<Y�`<jl`<�`<�_<�_<=�_<ь_<�_<��_<{`<l`<��`<&a<�oa<]�a<7�a<�b<S-b<7b<�7b<i1b<�'b<*b<�b<(b<|b<�
b<b<�b<�b<7b<�b<�)b<3b<J8b<�6b<C*b<�b<P�a<̪a<�aa<�a<g�`<�_`<�`< �_<e�_<�_<P�_<��_<k�_<�<`<s�`<��`<G?a<��a<��a<� b<:"b<�4b<e:b<�7b<�/b<�%b<+b<~b<wb<_b<b<b<�b<Sb<�b<�#b<�-b<�5b<'9b<S4b<]#b<�b<Z�a<��a<[Fa<��`<ԗ`<.C`<&�_<$�_<��_<��_<4�_<.�_<�`<�S`<K�`<�a<�Ua<͟a<��a<Eb<,$b<�1b<g4b<�/b<�&b<ub<�b<�b<{b<%b<�b< b<[
b<�b<�b<:!b<�*b<s1b<C2b<c)b<pb<��a<��a<sra<*!a<�`<?p`<�`<��_<�_<E�_<�_<�_<��_<�`<n^`<!�`<�a<u\a<��a<��a<��a<�b<�b<Ob<�b<B	b<x�a<M�a<��a<!�a<��a<G�a<��a<	�a<��a<��a<xb<Gb<b<b<"b<K�a<.�a<"�a<�7a<��`<�`<4`<��_<'�_<{_<@h_<#o_</�_<��_<�`<�``<$�`<1a<8]a<H�a<��a<�a<%b<�b<�b<��a<s�a<��a< �a<�a<	�a<E�a<��a<��a<��a<Z�a<��a<F�a<�  �  ��a<'b<xb<_�a<(�a<f�a<kua<�+a<�`<��`<�3`<[�_<�_<�_<��_<&�_<	�_<�_<>H`<��`<5�`<kBa<,�a<��a<��a<!b<$b<Ub<b<��a<v�a<��a<��a<o�a<?�a<T�a<��a<0�a<L�a<U�a<��a<b<�b<f b<�b<�b<��a<v�a<Uya<9-a<t�`<��`<<9`<G�_<T�_<��_<J�_<f�_<�_<S8`<��`<�`<51a<.�a<��a<M�a<�b<+1b<�7b<�3b<�(b<�b<cb<# b<��a<��a<��a<��a<^�a<�a<@b<b<�b<f+b<[5b<�7b<�.b<�b<#�a<��a<@sa<s#a<��`<V{`<s0`<�_<?�_<��_<��_<��_<!`<�Y`<�`<T�`<&Ra<*�a<�a<�	b<A(b</7b<k9b<2b<�%b<�b<�b<V�a<��a<��a<�a<P�a<��a<��a<�b<kb<#b<�/b<�7b<�6b<)b<eb<6�a<Ϣa<�Xa<�a<�`<�_`<�`<��_<4�_<T�_<3�_<s�_<�%`<Mo`<��`<�a<Mga<S�a<�a<Xb<')b<~3b<2b<�(b<�b<9b<��a<T�a<"�a<.�a<p�a<��a<r�a<��a<lb<zb<�!b<�,b<'2b<�,b<,b<��a<��a<a<�4a<.�`<��`<";`<;�_<S�_<��_<\�_<��_<E�_<�,`<y`<��`<�a<#ma<��a<��a<�b<�b<�b<Mb<Nb<�a<��a<{�a<	�a<-�a<��a<-�a<�a</�a<��a<D�a<U�a<�b<)b<0b<�b<	�a<��a<J�a<Ia<��`<P�`<{O`<`<(�_<�_<Ӌ_<r�_<�_<7�_<P*`<�z`<��`<"a<�la<��a<�a<"�a<�b<�b<A b<��a<��a<��a<��a<��a<��a<ٻa<J�a<�a<9�a<��a<��a<��a<�  �  �a<�b<H	b<�b<��a<1�a<�a<�Ga<D�`<�`<v``<�`<9�_<K�_<��_<�_<`�_<i.`<�s`<2�`<Oa<F]a<��a<j�a<)�a<Ub<�b<�b<$�a<��a<��a<�a<�a<��a<G�a<ڝa<Ӣa<%�a<��a<{�a<��a<��a<Ob<5b<O b<�b<�a<��a<��a<Ka<��`<��`<}g`<+`<b�_<\�_< �_<��_<:*`<g`<T�`<��`<�Oa</�a<��a<Yb<�&b<w5b<I6b<�+b<�b<�b<N�a<�a<
�a<��a<4�a<��a<�a<��a<��a<��a<L	b<?b<
/b<�7b<y4b<�"b<c b<��a<��a<Ca<��`<*�`<U``<(`<`<��_<�_<`<F`<��`<��`<4!a<�na<b�a<`�a<-b<-0b<�9b<�5b<(b<]b<�a<x�a<P�a<��a<v�a<w�a<��a<7�a<�a<��a<K�a<b<�$b<s3b<a8b<g0b<b<�a<s�a<�ta<�'a<(�`<-�`<�I`<�`<��_<b�_<,�_<�`<5V`<��`<��`<�6a<2�a<��a<��a<�b<b/b<�3b<f,b<2b<bb<��a<1�a<z�a<��a<3�a<�a<�a<b�a<��a<��a<��a<b<�$b<�/b<�0b<Q#b<�b<��a<,�a<�Ra<8a<��`<ai`<�*`<`�_<c�_<2�_<��_<i `<`[`<��`<E�`<O>a<&�a<��a<��a<�b<b<lb<�b<��a<)�a<��a<y�a<��a<��a<&�a<�a<1�a<Ȫa<_�a<��a<�a<��a<�b<	b<Pb<��a<5�a<0�a<Aca<6a<R�`<Dz`<�3`<�_<��_<��_<��_<��_<`<mW`<<�`<_�`<�>a<�a<ļa<Q�a<�a<?b<=b<O�a<f�a<a�a<=�a<�a<s�a<4�a<Q�a<��a<w�a<��a<z�a<��a<��a<�  �  ��a<��a<	b<�b<$�a<;�a<��a<�ia<�$a<�`<��`<]`<�/`<�`<N`<@`<�9`<�k`<D�`<��`<�8a<x}a<øa<��a<�b<�b<�b<�b<��a<H�a<��a<M�a<�ya<ia<�_a<�^a<�ea</ua<U�a<_�a<�a< �a<�b<�b<�"b<�b<�b<
�a<��a<Woa<w)a<;�`<ơ`<Ek`<(D`<�/`<{/`<�C`<k`<�`<��`<�,a<�ta<��a<��a<�b<10b<�8b<�1b<�b<hb<��a<(�a<��a<��a<��a<,a<�a<�a<˙a<��a<��a<��a<�
b<$b<�4b<9b<�-b<5b<V�a<�a<�ia<E"a<!�`<М`<j`<�G`<79`<?`<Y`<�`<��`<�a<mKa<v�a<��a<)b<4%b<�7b<F:b<r.b<|b<��a<��a<X�a<]�a<��a<σa<#a<��a<b�a<d�a<��a<I�a<d�a<tb<5+b<48b<A7b<`&b<b<�a<ɖa<8Qa<7	a<W�`<g�`<�Z`<B>`<6`<hB`<jb`<]�`<n�`<a<�^a<r�a<��a<r
b<�'b<�4b<2b<d"b<�	b<��a<w�a<d�a<`�a<��a<�{a<�ya<#�a<e�a<��a<j�a<��a<��a<�b<R*b<�2b<A,b<�b<9�a<$�a<�va<-/a<�`<��`<7k`<%B`<�+`<�)`< <`<Ea`<c�`<�`<a<oca<�a<��a<Lb<Cb<b<�b<�b<��a<L�a<��a<�a<>ta<?da<$\a<^\a<�da<�ta<��a<��a<E�a<�a<��a<,b<�b<b<��a<��a<��a<�>a<��`<-�`<Wp`<=`<�`<W`<�`<t*`<V`<B�`<�`<�a<\aa<g�a<��a<\�a<�b<�b<��a<��a<��a<v�a<+�a< ra<A^a<�Qa<Ma<�Pa<�\a<�oa<~�a<��a<�a<�  �  ��a<w�a<ab<b<{b<h�a<��a<}�a<}Qa<�a<K�`<��`<]|`<yd`<�]`<0i`<^�`<��`<��`<z$a<�ca<J�a<L�a<J�a<�b<pb<%
b<g�a<l�a<Ҩa<�a<�Ya<�9a<H"a<=a<ka<7a<�1a<�Oa<ua<�a<=�a<��a<db<� b<�#b<}b<��a<��a<�a<oYa<�a<[�`<+�`<i�`<ˀ`<ˀ`<��`<��`<��`<Ka<�]a<q�a<��a<Ib<T&b<97b<�7b<H(b<hb<��a<ݾa<�a<�pa<�Ra<9>a<�3a</5a<�Aa<yXa<Jxa<��a<��a<l�a<�b<v-b<�9b<�6b<�"b<�a<��a<��a<BUa<�a<	�`<�`<��`<��`<�`<\�`<��`<F�`<q:a<\ya<+�a<��a<Ab<^1b<<b<p6b<2"b<�b<��a<�a<ωa<�fa<mKa<4:a<�3a<�8a<�Ha<�ba<��a<��a<0�a<k�a<�b<q3b<�:b<�1b<=b<h�a<��a<!~a<?a<a<�`<>�`<׎`<��`<k�`<��`<t�`<4a<�Ja<��a<S�a<��a<�b<v1b<�6b<�+b<&b<��a<>�a<��a<�wa<�Va<�>a<1a<v.a<]7a<�Ja<�ga<�a<��a<��a<b< b<�0b<b2b<`#b<b<#�a<��a<"_a<�a<<�`<�`<e�`<�|`<�z`<��`<�`<��`<�a<Na<0�a<��a<��a<�b<Pb< b<wb<C�a<`�a<Q�a<Uva<bPa<M1a<�a<�a<�a<qa<�3a<�Ra<�xa<��a<��a<��a<�b<�b<�b<o�a<6�a<��a<�ha<�)a<��`<��`< �`<j`<�\`<�a`<�w`<��`<��`<�
a<~Ia<�a<��a<��a<� b<b<)b<��a<��a<˩a<�a<�Wa<�4a<@a<a<�a<�a<a<t1a<�Sa<�{a<�a<�  �  |�a<t�a<r�a<�
b<�
b<��a<h�a<U�a<�}a<8Ia<�a<��`<%�`<��`<�`<��`<��`<��`<(%a<�Xa<}�a<��a<��a<�b<b<Sb<E�a<0�a<�a<a<IKa<a<�`<��`<�`<\�`<��`<��`<�a<�;a<Wpa<a�a<F�a<��a<�b<�%b<X b<,b<E�a<=�a<�a<�Ua<�&a<��`<��`<��`<��`<��`<� a<)a</Ya<'�a<��a<p�a<�b<1b<�9b<h1b<db<��a<�a<z�a<�]a<2/a<�a<?�`<�`<��`<��`<a<�8a<�ha<��a<��a<��a<� b<�5b<$;b<O/b<gb<��a<b�a<G�a<	Ua<�'a<�a<��`<��`<F�`<��`<ma<�@a<ra<��a<�a<vb<�&b<k9b<�;b<e-b<0b<��a<h�a<�a<dNa<�!a<��`<��`<Y�`<�`<��`<a<yHa<rza<Ůa<W�a<�
b<})b<�9b<�8b<�'b<�b<f�a<3�a<ua<wCa<-a<�`<��`<��`<��`<q�`<�a<xLa<-a<W�a<�a<b<^)b<�6b<{3b<�b<��a<2�a<~�a<ja< 9a<ka<��`<��`<`�`<��`<��`<%a<�Ra<�a<۹a<a�a<(b<�)b<4b<6-b<Pb<��a<��a<��a<yYa<�(a<��`<��`<��`<��`<��`<�`<Ya<�Ka<�~a<~�a<r�a<�b<�b<�!b<b<��a<��a<��a<�ra<@>a<�a<5�`<��`<�`<�`<��`<E�`<[a<�Ba<�va<5�a<A�a<��a<�b<`b<b<��a<)�a<h�a<�\a<�(a<��`<��`<�`<�`<�`<�`<\�`<Ta<bBa<�va<��a<�a<��a<�b<�
b<'�a<��a<�a<��a<Oa<Za<��`<��`<ٶ`<h�`<O�`<�`<��`<a<�Ia<�~a<�  �  0�a<��a<��a<.b<Kb<#b<��a<��a<}�a< |a<�Ta<�2a<�a<K
a<a<�a<�a<
<a<�_a<��a<�a<J�a<�a<Lb<�b<�b<��a<5�a<��a<IQa<+a<"�`<ǧ`<?�`<�n`<Dk`<z`<S�`<�`<P�`<�=a<\}a<&�a<��a<�b<�!b<�$b<�b<(�a<B�a<~�a<�a<�fa<rHa<(3a<#(a<�(a<d4a<�Ja<Dja<��a<�a<��a<h
b<�&b<�6b<�6b<-&b<�b<��a<�a<;`a<S"a<-�`<�`<�`< �`<��`<}�`<��`<��`<�/a<na<a�a<��a<�b<�,b<�9b<�6b<�$b<�b<��a<��a<׎a<�ja<Na<S;a<3a<j6a<�Da<�]a<�~a<
�a<��a<��a<b<�1b<<b<�5b<mb<E�a<N�a<
�a<ILa<�a<'�`<)�`<A�`<�`<�`<�`<i�`<�a<�Da<C�a<�a<��a<�b<�2b<�:b<�1b<mb<
�a<4�a<S�a<y�a<_^a<�Da<�4a<0a<�6a<�Ha<!da<Z�a<��a<�a<u�a<�b<�1b<�6b<�*b<b< �a<��a<�pa<�1a<4�`<#�`<ݟ`<c�`<B�`<%�`<q�`<�`<Ba<�Sa<Αa<9�a<O�a<�b<0b<�1b<�#b<�b<��a<*�a<ҏa<�ha<_Ha<"1a<)$a<�"a<�,a<�@a<�^a<�a<w�a<��a<m�a<<b<U b<�b<�b<��a<��a<ƀa<�Aa<�a<��`<��`<�y`<i`<_j`<B}`<2�`<c�`<�	a<�Ga<��a<@�a<%�a<Db<!b<�b<��a<Y�a<ֵa<�a<�ba<->a<� a<�a<a<�a<a<h.a<YOa<`va<ןa<��a<��a<Pb<;b<�b<9�a<��a<��a<LYa<ia<��`<!�`<#~`<Hc`<?Y`<fa`<�z`<0�`<��`<�a<Sa<�  �  �ka<��a<��a<D�a<B	b<T	b<��a<~�a<3�a<"�a<��a<�qa<a_a<`Ta<~Qa<�Va<qda<ya<�a<Ųa<��a<��a<�b<�b<�b<4�a<��a<��a<gha<�"a<��`<��`<�_`<�5`<�`<�`<�*`<�N`<H�`<'�`<�a<Ta<��a<��a<��a<#b<�$b<n b<b</�a<��a<��a<(�a<-�a<�za<sa<�sa<u|a<�a<h�a<P�a<F�a<� b<_b<�/b<!7b<2/b<b<G�a<I�a<�ua<�.a<(�`<>�`<r`<�L`<�:`<�<`<sS`<p|`<��`<X�`<�>a<1�a<��a<}�a<%b<G4b<Y9b<�/b<b<E�a<A�a<��a<��a<-�a<W�a<z~a<��a<f�a<��a<��a<T�a<��a<�b<�(b<�7b<�9b<�+b<�b<;�a<��a<�_a<�a<R�`<��`<Od`<E`<�9`<�B`<�_`<�`<]�`<.a<�Va<��a<�a<�b<�'b<~7b<07b<.)b<�b<��a<��a<��a<l�a<t�a<�~a<�{a<d�a<E�a<E�a<Z�a<��a<��a<�b<D*b<T5b<�1b<qb<{�a<Y�a<��a<JBa<��`<�`<U}`<ZR`<r9`<�4`<�D`<�g`<R�`<�`<=!a<wha<˪a<�a<�b<�'b<_1b<�+b<\b<��a<`�a<U�a<�a<�a<�xa<!oa<�ma<�ta<L�a<��a<��a<��a<��a<h	b<b<� b<Zb<��a<��a<9�a<Xa<Ka<��`<��`<�P`<�*`<�`<;`<=/`<�W`<E�`<��`<La<e^a<��a<��a<��a<ob<�b<�b<��a<-�a<��a<��a<Dza<�da<�Va<^Pa<bRa<�\a<^na<��a<��a<��a<m�a<��a<fb<	b<��a<k�a<߭a<lra<�-a<	�`<j�`<�b`<[2`</`<�`<`<>.`<�\`<��`<��`<�&a<�  �  �Ja<n�a<4�a<Y�a<�b<�	b<]b<{�a<S�a<��a<�a<ݥa<r�a<o�a<��a<\�a<U�a<��a<y�a<)�a<��a<��a<�b<{b<�b<��a<��a<��a<WEa<6�`<��`<�_`<� `<��_<��_<X�_<��_<�`<3G`<��`<g�`<�-a<�xa<w�a<�a<ib<R b<�#b<mb<*b<��a<)�a<U�a<^�a<i�a<ݱa<��a<��a<�a<q�a<��a<��a<�b<�(b<�3b<�3b<'%b<Qb<��a<�a<;Pa<pa<d�`<�k`<�0`<�`<0�_<��_<�`<}<`<�z`<B�`<a<Qaa<l�a<��a<�b<�+b<v7b<�5b<W)b<Wb<� b<e�a<��a<��a<u�a<��a<D�a<�a<H�a<T�a<��a<�b<�"b<o2b<r9b<4b<�b<��a<��a<P�a<�7a<��`<6�`<(W`<!`<��_<��_<�_<]`<�O`<��`<��`<�-a<Gza<ͽa<1�a<�b<�0b<�7b<�1b<�"b<b<�a<�a<s�a<��a<�a<Ժa<�a<:�a<��a< �a<��a<�b<$b<21b<=4b<�)b<
b<S�a<��a<{ea<�a<o�`<�}`<�=`<+`<q�_<I�_<��_<&`<6_`<��`<�`<Ba<ʋa<
�a<*�a<�b<!-b<�.b<�$b<�b<��a<��a<.�a<H�a<b�a<�a<��a<��a<6�a<��a<[�a<3�a<�b<�b<Db<cb<Sb<�a<,�a<	}a<�2a<�`<�`<aK`<�`<U�_<H�_<�_<��_<�`<XU`<q�`<��`<�:a<�a<��a<��a<�b<b<�b<��a<3�a<��a<#�a<�a<=�a<��a<��a<��a<3�a<�a<ݳa<'�a<��a<e�a<b<�b<Ob<��a<��a<e�a<�Qa<�a<:�`<\i`<C%`<��_<��_<+�_<y�_<��_<�`<�a`<�`<��`<�  �  �.a<xa<��a<��a<��a<qb<�b<� b<��a<�a<��a<��a<G�a<�a<A�a<��a<%�a<B�a<��a<�a<b�a<Lb<�b<�b<��a<4�a<F�a<>sa<f(a<�`<��`<Z2`<��_<��_<%�_<d�_<M�_<B�_<�`< d`<��`<pa<�^a<ۤa</�a<�b<b<=$b<"b<�b<�b<�a<9�a<�a<u�a<�a<��a<��a<C�a<�a<�b<b<J$b<0b<5b</b<b<��a<��a<�a<�1a<l�`<t�`<�<`<��_<�_<I�_<�_<��_<�	`<�L`<��`<V�`<�Ca<P�a<��a<�b<�"b<!4b<F8b<+2b<`&b<�b<�	b<��a<��a<o�a<:�a<0�a<e�a<��a<�b<3b<� b<�.b<�7b<�8b<�-b<�b<��a<�a< ha<#a<��`<�o`<�&`<��_<��_<ٹ_<��_<b�_<�`<Ff`<˷`<�a<�^a<r�a<��a<�b<�)b<Q6b<t6b<�-b< b<�b<�b<r�a<s�a<��a<f�a<�a<�a<��a<b<�b<z!b<�-b<z4b<�1b<�!b<b<��a<�a<�Ha<��`<b�`<hP`<�`<��_<�_<Q�_<Q�_<M�_<�/`<�z`<d�`<�"a<�qa<i�a<8�a<6b<�'b<P/b<f+b<< b<Yb<�b<�a<��a<m�a<�a<��a<�a<x�a<c�a<�a<�b<b<b<f b<�b<Kb<��a<�a<�ca<Ia<�`<�i`<S`<0�_<�_<e�_<r�_<��_</�_<]'`<�u`<�`<�a< ia<��a<w�a<��a<�
b<?b<�b<2�a<�a<d�a<��a<��a<��a<�a<��a<{�a<��a<D�a<x�a<�a<X�a<[b<b<��a<��a<t�a<�~a<�6a<��`<<�`<�=`<��_<�_<ڕ_<)�_<E�_<�_<��_<�5`<X�`<��`<�  �  ta<ia<��a<`�a<+�a<`b<�
b<�b<��a<��a<��a<��a<C�a<��a<��a<��a<��a<,�a<x�a<��a<Mb<�b<�b<�
b<��a<��a<ߤa<vca<Ua<}�`<�g`<d`<��_<��_<�{_<�v_<��_<^�_<E�_<�H`<��`<��`<�Ma<�a<��a</�a<�b<X#b<O%b<� b<b<b<eb<b<�a<>�a<,�a<�b<�b<�b<b<"b<�,b<�3b<�4b<�*b<�b<��a<:�a<�na<Ea<��`<�n`<�`<��_<~�_<ė_<��_<Ķ_<��_<Y/`<q�`<m�`<W0a<.�a<��a<A�a<Pb<�0b<�8b<�6b<�/b<�%b<9b<Lb<�b<�b<�
b<b<�b<b<b<4"b<],b<a5b<�9b<�6b<d(b<�b<;�a<9�a<,Va<�a<3�`<�S`<�`<��_<��_<:�_<��_<��_<��_<J`<��`<�`<+La<`�a<��a<�b<h$b<A4b<#8b<&4b<h+b<!b<�b<Ab<ub<�b<�b<�b<�b<zb<b<s!b<k+b<�2b<;5b<�.b<�b<C�a<s�a<R�a<}5a<��`<��`<r3`<
�_<��_<��_<��_<��_<e�_<@`<�_`<]�`<"a<�`a<n�a<��a<�
b<o#b<j.b<�.b<(b<�b<�b<=	b<�b<�a<C�a<>�a<��a<��a<�b<�	b<�b<wb<� b<�b<�b<�a<c�a<��a<�Ra< a<]�`<!O`<N�_<��_<Z�_<�t_<w_<��_<�_<
`<�[`<�`<�	a<�Xa<��a<��a<f�a<db<�b<Wb<�b<�a<��a<s�a<��a<��a<l�a<��a<��a<��a<��a<w�a<g�a<6b<	b<eb<��a<��a< �a<�oa<�$a<�`<�w`<�!`<��_<��_<�r_<�d_<p_<~�_<��_<A`<Gn`<��`<�  �  Ma<�ca<��a<#�a<�a<�b<_b<	b<�b<��a<d�a<��a<|�a<��a<��a<��a<��a<��a<��a<,�a<b<nb<"b<�	b<�a<}�a<B�a<�]a<�a<��`<�^`<G`<��_<:�_<�o_<�j_<�_<�_<��_<�?`<f�`<��`<�Ga<��a<��a<N�a<�b<9#b<�&b<�"b<�b<�b<�b<�
b<�b<Ob<I	b<bb<ab<b<b<�%b</b<25b<�4b<u)b<b<��a<.�a<ia<�a<��`<Ee`<I`<x�_<~�_<��_<g�_<�_<��_< %`<ax`<w�`<�)a<�za<�a<��a<�b<�/b<�8b<�8b<|2b<:*b<�"b<�b<�b<\b<�b<b<�b<eb< b<�'b<�/b<�7b<�:b<�6b<k&b<b<�a<ۛa< Pa<`�`<��`<�I`<��_<�_<~�_<�_<{�_<�_<��_<#@`<�`<��`<Fa<�a<��a<�b<C"b<�3b<�8b<56b<�.b<&&b<ub<ab<�b<jb<�b<Nb<�b<Ob<�b<&b<<.b<�4b<�5b<�-b<.b<��a<��a<�~a</a<(�`<�}`<U)`<��_<ʪ_<f�_<��_<��_<��_<�`<ZV`<
�`<6a<�Za<D�a<��a<�b<�!b<K.b<�/b<s*b<�!b<�b<{b<�
b<�b<Tb<[b<�b<�b<Y	b<xb<�b<�b<B"b<�b<6b<I�a<��a<~�a<Ma<E�`<)�`<�E`<��_<&�_<\�_<�h_<�j_<��_<ҹ_<��_<�R`<'�`<a<7Sa<9�a<Z�a<��a<?b<�b<b<Fb<s�a<9�a<�a<��a<��a<��a<g�a<��a<(�a<��a<��a<��a<bb<g
b<�b<��a<��a<��a<�ja<�a<��`<�n`<`<��_<�_<�f_<sX_<�c_<ֈ_<��_<d`<�e`<��`<�  �  ta<ia<��a<`�a<+�a<`b<�
b<�b<��a<��a<��a<��a<C�a<��a<��a<��a<��a<,�a<x�a<��a<Mb<�b<�b<�
b<��a<��a<ߤa<vca<Ua<}�`<�g`<d`<��_<��_<�{_<�v_<��_<^�_<E�_<�H`<��`<��`<�Ma<�a<��a</�a<�b<X#b<O%b<� b<b<b<eb<b<�a<>�a<,�a<�b<�b<�b<b<"b<�,b<�3b<�4b<�*b<�b<��a<:�a<�na<Ea<��`<�n`<�`<��_<~�_<ė_<��_<Ķ_<��_<Y/`<q�`<m�`<W0a<.�a<��a<A�a<Pb<�0b<�8b<�6b<�/b<�%b<9b<Lb<�b<�b<�
b<b<�b<b<b<4"b<],b<a5b<�9b<�6b<d(b<�b<;�a<9�a<,Va<�a<3�`<�S`<�`<��_<��_<:�_<��_<��_<��_<J`<��`<�`<+La<`�a<��a<�b<h$b<A4b<#8b<&4b<h+b<!b<�b<Ab<ub<�b<�b<�b<�b<zb<b<s!b<k+b<�2b<;5b<�.b<�b<C�a<s�a<R�a<}5a<��`<��`<r3`<
�_<��_<��_<��_<��_<e�_<@`<�_`<]�`<"a<�`a<n�a<��a<�
b<o#b<j.b<�.b<(b<�b<�b<=	b<�b<�a<C�a<>�a<��a<��a<�b<�	b<�b<wb<� b<�b<�b<�a<c�a<��a<�Ra< a<]�`<!O`<N�_<��_<Z�_<�t_<w_<��_<�_<
`<�[`<�`<�	a<�Xa<��a<��a<f�a<db<�b<Wb<�b<�a<��a<s�a<��a<��a<l�a<��a<��a<��a<��a<w�a<g�a<6b<	b<eb<��a<��a< �a<�oa<�$a<�`<�w`<�!`<��_<��_<�r_<�d_<p_<~�_<��_<A`<Gn`<��`<�  �  �.a<xa<��a<��a<��a<qb<�b<� b<��a<�a<��a<��a<G�a<�a<A�a<��a<%�a<B�a<��a<�a<b�a<Lb<�b<�b<��a<4�a<F�a<>sa<f(a<�`<��`<Z2`<��_<��_<%�_<d�_<M�_<B�_<�`< d`<��`<pa<�^a<ۤa</�a<�b<b<=$b<"b<�b<�b<�a<9�a<�a<u�a<�a<��a<��a<C�a<�a<�b<b<J$b<0b<5b</b<b<��a<��a<�a<�1a<l�`<t�`<�<`<��_<�_<I�_<�_<��_<�	`<�L`<��`<V�`<�Ca<P�a<��a<�b<�"b<!4b<F8b<+2b<`&b<�b<�	b<��a<��a<o�a<:�a<0�a<e�a<��a<�b<3b<� b<�.b<�7b<�8b<�-b<�b<��a<�a< ha<#a<��`<�o`<�&`<��_<��_<ٹ_<��_<b�_<�`<Ff`<˷`<�a<�^a<r�a<��a<�b<�)b<Q6b<t6b<�-b< b<�b<�b<r�a<s�a<��a<f�a<�a<�a<��a<b<�b<z!b<�-b<z4b<�1b<�!b<b<��a<�a<�Ha<��`<b�`<hP`<�`<��_<�_<Q�_<Q�_<M�_<�/`<�z`<d�`<�"a<�qa<i�a<8�a<6b<�'b<P/b<f+b<< b<Yb<�b<�a<��a<m�a<�a<��a<�a<x�a<c�a<�a<�b<b<b<f b<�b<Kb<��a<�a<�ca<Ia<�`<�i`<S`<0�_<�_<e�_<r�_<��_</�_<]'`<�u`<�`<�a< ia<��a<w�a<��a<�
b<?b<�b<2�a<�a<d�a<��a<��a<��a<�a<��a<{�a<��a<D�a<x�a<�a<X�a<[b<b<��a<��a<t�a<�~a<�6a<��`<<�`<�=`<��_<�_<ڕ_<)�_<E�_<�_<��_<�5`<X�`<��`<�  �  �Ja<n�a<4�a<Y�a<�b<�	b<]b<{�a<S�a<��a<�a<ݥa<r�a<o�a<��a<\�a<U�a<��a<y�a<)�a<��a<��a<�b<{b<�b<��a<��a<��a<WEa<6�`<��`<�_`<� `<��_<��_<X�_<��_<�`<3G`<��`<g�`<�-a<�xa<w�a<�a<ib<R b<�#b<mb<*b<��a<)�a<U�a<^�a<i�a<ݱa<��a<��a<�a<q�a<��a<��a<�b<�(b<�3b<�3b<'%b<Qb<��a<�a<;Pa<pa<d�`<�k`<�0`<�`<0�_<��_<�`<}<`<�z`<B�`<a<Qaa<l�a<��a<�b<�+b<v7b<�5b<W)b<Wb<� b<e�a<��a<��a<u�a<��a<D�a<�a<H�a<T�a<��a<�b<�"b<o2b<r9b<4b<�b<��a<��a<P�a<�7a<��`<6�`<(W`<!`<��_<��_<�_<]`<�O`<��`<��`<�-a<Gza<ͽa<1�a<�b<�0b<�7b<�1b<�"b<b<�a<�a<s�a<��a<�a<Ժa<�a<:�a<��a< �a<��a<�b<$b<21b<=4b<�)b<
b<S�a<��a<{ea<�a<o�`<�}`<�=`<+`<q�_<I�_<��_<&`<6_`<��`<�`<Ba<ʋa<
�a<*�a<�b<!-b<�.b<�$b<�b<��a<��a<.�a<H�a<b�a<�a<��a<��a<6�a<��a<[�a<3�a<�b<�b<Db<cb<Sb<�a<,�a<	}a<�2a<�`<�`<aK`<�`<U�_<H�_<�_<��_<�`<XU`<q�`<��`<�:a<�a<��a<��a<�b<b<�b<��a<3�a<��a<#�a<�a<=�a<��a<��a<��a<3�a<�a<ݳa<'�a<��a<e�a<b<�b<Ob<��a<��a<e�a<�Qa<�a<:�`<\i`<C%`<��_<��_<+�_<y�_<��_<�`<�a`<�`<��`<�  �  �ka<��a<��a<D�a<B	b<T	b<��a<~�a<3�a<"�a<��a<�qa<a_a<`Ta<~Qa<�Va<qda<ya<�a<Ųa<��a<��a<�b<�b<�b<4�a<��a<��a<gha<�"a<��`<��`<�_`<�5`<�`<�`<�*`<�N`<H�`<'�`<�a<Ta<��a<��a<��a<#b<�$b<n b<b</�a<��a<��a<(�a<-�a<�za<sa<�sa<u|a<�a<h�a<P�a<F�a<� b<_b<�/b<!7b<2/b<b<G�a<I�a<�ua<�.a<(�`<>�`<r`<�L`<�:`<�<`<sS`<p|`<��`<X�`<�>a<1�a<��a<}�a<%b<G4b<Y9b<�/b<b<E�a<A�a<��a<��a<-�a<W�a<z~a<��a<f�a<��a<��a<T�a<��a<�b<�(b<�7b<�9b<�+b<�b<;�a<��a<�_a<�a<R�`<��`<Od`<E`<�9`<�B`<�_`<�`<]�`<.a<�Va<��a<�a<�b<�'b<~7b<07b<.)b<�b<��a<��a<��a<l�a<t�a<�~a<�{a<d�a<E�a<E�a<Z�a<��a<��a<�b<D*b<T5b<�1b<qb<{�a<Y�a<��a<JBa<��`<�`<U}`<ZR`<r9`<�4`<�D`<�g`<R�`<�`<=!a<wha<˪a<�a<�b<�'b<_1b<�+b<\b<��a<`�a<U�a<�a<�a<�xa<!oa<�ma<�ta<L�a<��a<��a<��a<��a<h	b<b<� b<Zb<��a<��a<9�a<Xa<Ka<��`<��`<�P`<�*`<�`<;`<=/`<�W`<E�`<��`<La<e^a<��a<��a<��a<ob<�b<�b<��a<-�a<��a<��a<Dza<�da<�Va<^Pa<bRa<�\a<^na<��a<��a<��a<m�a<��a<fb<	b<��a<k�a<߭a<lra<�-a<	�`<j�`<�b`<[2`</`<�`<`<>.`<�\`<��`<��`<�&a<�  �  0�a<��a<��a<.b<Kb<#b<��a<��a<}�a< |a<�Ta<�2a<�a<K
a<a<�a<�a<
<a<�_a<��a<�a<J�a<�a<Lb<�b<�b<��a<5�a<��a<IQa<+a<"�`<ǧ`<?�`<�n`<Dk`<z`<S�`<�`<P�`<�=a<\}a<&�a<��a<�b<�!b<�$b<�b<(�a<B�a<~�a<�a<�fa<rHa<(3a<#(a<�(a<d4a<�Ja<Dja<��a<�a<��a<h
b<�&b<�6b<�6b<-&b<�b<��a<�a<;`a<S"a<-�`<�`<�`< �`<��`<}�`<��`<��`<�/a<na<a�a<��a<�b<�,b<�9b<�6b<�$b<�b<��a<��a<׎a<�ja<Na<S;a<3a<j6a<�Da<�]a<�~a<
�a<��a<��a<b<�1b<<b<�5b<mb<E�a<N�a<
�a<ILa<�a<'�`<)�`<A�`<�`<�`<�`<i�`<�a<�Da<C�a<�a<��a<�b<�2b<�:b<�1b<mb<
�a<4�a<S�a<y�a<_^a<�Da<�4a<0a<�6a<�Ha<!da<Z�a<��a<�a<u�a<�b<�1b<�6b<�*b<b< �a<��a<�pa<�1a<4�`<#�`<ݟ`<c�`<B�`<%�`<q�`<�`<Ba<�Sa<Αa<9�a<O�a<�b<0b<�1b<�#b<�b<��a<*�a<ҏa<�ha<_Ha<"1a<)$a<�"a<�,a<�@a<�^a<�a<w�a<��a<m�a<<b<U b<�b<�b<��a<��a<ƀa<�Aa<�a<��`<��`<�y`<i`<_j`<B}`<2�`<c�`<�	a<�Ga<��a<@�a<%�a<Db<!b<�b<��a<Y�a<ֵa<�a<�ba<->a<� a<�a<a<�a<a<h.a<YOa<`va<ןa<��a<��a<Pb<;b<�b<9�a<��a<��a<LYa<ia<��`<!�`<#~`<Hc`<?Y`<fa`<�z`<0�`<��`<�a<Sa<�  �  |�a<t�a<r�a<�
b<�
b<��a<h�a<U�a<�}a<8Ia<�a<��`<%�`<��`<�`<��`<��`<��`<(%a<�Xa<}�a<��a<��a<�b<b<Sb<E�a<0�a<�a<a<IKa<a<�`<��`<�`<\�`<��`<��`<�a<�;a<Wpa<a�a<F�a<��a<�b<�%b<X b<,b<E�a<=�a<�a<�Ua<�&a<��`<��`<��`<��`<��`<� a<)a</Ya<'�a<��a<p�a<�b<1b<�9b<h1b<db<��a<�a<z�a<�]a<2/a<�a<?�`<�`<��`<��`<a<�8a<�ha<��a<��a<��a<� b<�5b<$;b<O/b<gb<��a<b�a<G�a<	Ua<�'a<�a<��`<��`<F�`<��`<ma<�@a<ra<��a<�a<vb<�&b<k9b<�;b<e-b<0b<��a<h�a<�a<dNa<�!a<��`<��`<Y�`<�`<��`<a<yHa<rza<Ůa<W�a<�
b<})b<�9b<�8b<�'b<�b<f�a<3�a<ua<wCa<-a<�`<��`<��`<��`<q�`<�a<xLa<-a<W�a<�a<b<^)b<�6b<{3b<�b<��a<2�a<~�a<ja< 9a<ka<��`<��`<`�`<��`<��`<%a<�Ra<�a<۹a<a�a<(b<�)b<4b<6-b<Pb<��a<��a<��a<yYa<�(a<��`<��`<��`<��`<��`<�`<Ya<�Ka<�~a<~�a<r�a<�b<�b<�!b<b<��a<��a<��a<�ra<@>a<�a<5�`<��`<�`<�`<��`<E�`<[a<�Ba<�va<5�a<A�a<��a<�b<`b<b<��a<)�a<h�a<�\a<�(a<��`<��`<�`<�`<�`<�`<\�`<Ta<bBa<�va<��a<�a<��a<�b<�
b<'�a<��a<�a<��a<Oa<Za<��`<��`<ٶ`<h�`<O�`<�`<��`<a<�Ia<�~a<�  �  ��a<w�a<ab<b<{b<h�a<��a<}�a<}Qa<�a<K�`<��`<]|`<yd`<�]`<0i`<^�`<��`<��`<z$a<�ca<J�a<L�a<J�a<�b<pb<%
b<g�a<l�a<Ҩa<�a<�Ya<�9a<H"a<=a<ka<7a<�1a<�Oa<ua<�a<=�a<��a<db<� b<�#b<}b<��a<��a<�a<oYa<�a<[�`<+�`<i�`<ˀ`<ˀ`<��`<��`<��`<Ka<�]a<q�a<��a<Ib<T&b<97b<�7b<H(b<hb<��a<ݾa<�a<�pa<�Ra<9>a<�3a</5a<�Aa<yXa<Jxa<��a<��a<l�a<�b<v-b<�9b<�6b<�"b<�a<��a<��a<BUa<�a<	�`<�`<��`<��`<�`<\�`<��`<F�`<q:a<\ya<+�a<��a<Ab<^1b<<b<p6b<2"b<�b<��a<�a<ωa<�fa<mKa<4:a<�3a<�8a<�Ha<�ba<��a<��a<0�a<k�a<�b<q3b<�:b<�1b<=b<h�a<��a<!~a<?a<a<�`<>�`<׎`<��`<k�`<��`<t�`<4a<�Ja<��a<S�a<��a<�b<v1b<�6b<�+b<&b<��a<>�a<��a<�wa<�Va<�>a<1a<v.a<]7a<�Ja<�ga<�a<��a<��a<b< b<�0b<b2b<`#b<b<#�a<��a<"_a<�a<<�`<�`<e�`<�|`<�z`<��`<�`<��`<�a<Na<0�a<��a<��a<�b<Pb< b<wb<C�a<`�a<Q�a<Uva<bPa<M1a<�a<�a<�a<qa<�3a<�Ra<�xa<��a<��a<��a<�b<�b<�b<o�a<6�a<��a<�ha<�)a<��`<��`< �`<j`<�\`<�a`<�w`<��`<��`<�
a<~Ia<�a<��a<��a<� b<b<)b<��a<��a<˩a<�a<�Wa<�4a<@a<a<�a<�a<a<t1a<�Sa<�{a<�a<�  �  ��a<��a<	b<�b<$�a<;�a<��a<�ia<�$a<�`<��`<]`<�/`<�`<N`<@`<�9`<�k`<D�`<��`<�8a<x}a<øa<��a<�b<�b<�b<�b<��a<H�a<��a<M�a<�ya<ia<�_a<�^a<�ea</ua<U�a<_�a<�a< �a<�b<�b<�"b<�b<�b<
�a<��a<Woa<w)a<;�`<ơ`<Ek`<(D`<�/`<{/`<�C`<k`<�`<��`<�,a<�ta<��a<��a<�b<10b<�8b<�1b<�b<hb<��a<(�a<��a<��a<��a<,a<�a<�a<˙a<��a<��a<��a<�
b<$b<�4b<9b<�-b<5b<V�a<�a<�ia<E"a<!�`<М`<j`<�G`<79`<?`<Y`<�`<��`<�a<mKa<v�a<��a<)b<4%b<�7b<F:b<r.b<|b<��a<��a<X�a<]�a<��a<σa<#a<��a<b�a<d�a<��a<I�a<d�a<tb<5+b<48b<A7b<`&b<b<�a<ɖa<8Qa<7	a<W�`<g�`<�Z`<B>`<6`<hB`<jb`<]�`<n�`<a<�^a<r�a<��a<r
b<�'b<�4b<2b<d"b<�	b<��a<w�a<d�a<`�a<��a<�{a<�ya<#�a<e�a<��a<j�a<��a<��a<�b<R*b<�2b<A,b<�b<9�a<$�a<�va<-/a<�`<��`<7k`<%B`<�+`<�)`< <`<Ea`<c�`<�`<a<oca<�a<��a<Lb<Cb<b<�b<�b<��a<L�a<��a<�a<>ta<?da<$\a<^\a<�da<�ta<��a<��a<E�a<�a<��a<,b<�b<b<��a<��a<��a<�>a<��`<-�`<Wp`<=`<�`<W`<�`<t*`<V`<B�`<�`<�a<\aa<g�a<��a<\�a<�b<�b<��a<��a<��a<v�a<+�a< ra<A^a<�Qa<Ma<�Pa<�\a<�oa<~�a<��a<�a<�  �  �a<�b<H	b<�b<��a<1�a<�a<�Ga<D�`<�`<v``<�`<9�_<K�_<��_<�_<`�_<i.`<�s`<2�`<Oa<F]a<��a<j�a<)�a<Ub<�b<�b<$�a<��a<��a<�a<�a<��a<G�a<ڝa<Ӣa<%�a<��a<{�a<��a<��a<Ob<5b<O b<�b<�a<��a<��a<Ka<��`<��`<}g`<+`<b�_<\�_< �_<��_<:*`<g`<T�`<��`<�Oa</�a<��a<Yb<�&b<w5b<I6b<�+b<�b<�b<N�a<�a<
�a<��a<4�a<��a<�a<��a<��a<��a<L	b<?b<
/b<�7b<y4b<�"b<c b<��a<��a<Ca<��`<*�`<U``<(`<`<��_<�_<`<F`<��`<��`<4!a<�na<b�a<`�a<-b<-0b<�9b<�5b<(b<]b<�a<x�a<P�a<��a<v�a<w�a<��a<7�a<�a<��a<K�a<b<�$b<s3b<a8b<g0b<b<�a<s�a<�ta<�'a<(�`<-�`<�I`<�`<��_<b�_<,�_<�`<5V`<��`<��`<�6a<2�a<��a<��a<�b<b/b<�3b<f,b<2b<bb<��a<1�a<z�a<��a<3�a<�a<�a<b�a<��a<��a<��a<b<�$b<�/b<�0b<Q#b<�b<��a<,�a<�Ra<8a<��`<ai`<�*`<`�_<c�_<2�_<��_<i `<`[`<��`<E�`<O>a<&�a<��a<��a<�b<b<lb<�b<��a<)�a<��a<y�a<��a<��a<&�a<�a<1�a<Ȫa<_�a<��a<�a<��a<�b<	b<Pb<��a<5�a<0�a<Aca<6a<R�`<Dz`<�3`<�_<��_<��_<��_<��_<`<mW`<<�`<_�`<�>a<�a<ļa<Q�a<�a<?b<=b<O�a<f�a<a�a<=�a<�a<s�a<4�a<Q�a<��a<w�a<��a<z�a<��a<��a<�  �  ��a<'b<xb<_�a<(�a<f�a<kua<�+a<�`<��`<�3`<[�_<�_<�_<��_<&�_<	�_<�_<>H`<��`<5�`<kBa<,�a<��a<��a<!b<$b<Ub<b<��a<v�a<��a<��a<o�a<?�a<T�a<��a<0�a<L�a<U�a<��a<b<�b<f b<�b<�b<��a<v�a<Uya<9-a<t�`<��`<<9`<G�_<T�_<��_<J�_<f�_<�_<S8`<��`<�`<51a<.�a<��a<M�a<�b<+1b<�7b<�3b<�(b<�b<cb<# b<��a<��a<��a<��a<^�a<�a<@b<b<�b<f+b<[5b<�7b<�.b<�b<#�a<��a<@sa<s#a<��`<V{`<s0`<�_<?�_<��_<��_<��_<!`<�Y`<�`<T�`<&Ra<*�a<�a<�	b<A(b</7b<k9b<2b<�%b<�b<�b<V�a<��a<��a<�a<P�a<��a<��a<�b<kb<#b<�/b<�7b<�6b<)b<eb<6�a<Ϣa<�Xa<�a<�`<�_`<�`<��_<4�_<T�_<3�_<s�_<�%`<Mo`<��`<�a<Mga<S�a<�a<Xb<')b<~3b<2b<�(b<�b<9b<��a<T�a<"�a<.�a<p�a<��a<r�a<��a<lb<zb<�!b<�,b<'2b<�,b<,b<��a<��a<a<�4a<.�`<��`<";`<;�_<S�_<��_<\�_<��_<E�_<�,`<y`<��`<�a<#ma<��a<��a<�b<�b<�b<Mb<Nb<�a<��a<{�a<	�a<-�a<��a<-�a<�a</�a<��a<D�a<U�a<�b<)b<0b<�b<	�a<��a<J�a<Ia<��`<P�`<{O`<`<(�_<�_<Ӌ_<r�_<�_<7�_<P*`<�z`<��`<"a<�la<��a<�a<"�a<�b<�b<A b<��a<��a<��a<��a<��a<��a<ٻa<J�a<�a<9�a<��a<��a<��a<�  �  �b<�	b<5b<��a<k�a<��a<-fa<ea<�`<�k`<�`<��_<q�_<�r_<i_</y_<ˡ_<D�_<�,`<��`<��`<�0a<�{a<y�a<��a<*b<�b<�b<�b<!b<��a<h�a<\�a<��a<4�a<��a<��a<�a<��a<� b<Ub<Fb<:b< b<(b<�b<��a<~�a<ia<�a<Y�`<jl`<�`<�_<�_<=�_<ь_<�_<��_<{`<l`<��`<&a<�oa<]�a<7�a<�b<S-b<7b<�7b<i1b<�'b<*b<�b<(b<|b<�
b<b<�b<�b<7b<�b<�)b<3b<J8b<�6b<C*b<�b<P�a<̪a<�aa<�a<g�`<�_`<�`< �_<e�_<�_<P�_<��_<k�_<�<`<s�`<��`<G?a<��a<��a<� b<:"b<�4b<e:b<�7b<�/b<�%b<+b<~b<wb<_b<b<b<�b<Sb<�b<�#b<�-b<�5b<'9b<S4b<]#b<�b<Z�a<��a<[Fa<��`<ԗ`<.C`<&�_<$�_<��_<��_<4�_<.�_<�`<�S`<K�`<�a<�Ua<͟a<��a<Eb<,$b<�1b<g4b<�/b<�&b<ub<�b<�b<{b<%b<�b< b<[
b<�b<�b<:!b<�*b<s1b<C2b<c)b<pb<��a<��a<sra<*!a<�`<?p`<�`<��_<�_<E�_<�_<�_<��_<�`<n^`<!�`<�a<u\a<��a<��a<��a<�b<�b<Ob<�b<B	b<x�a<M�a<��a<!�a<��a<G�a<��a<	�a<��a<��a<xb<Gb<b<b<"b<K�a<.�a<"�a<�7a<��`<�`<4`<��_<'�_<{_<@h_<#o_</�_<��_<�`<�``<$�`<1a<8]a<H�a<��a<�a<%b<�b<�b<��a<s�a<��a< �a<�a<	�a<E�a<��a<��a<��a<Z�a<��a<F�a<�  �  V�a<��a<p�a<J�a<�a<i�a<(^a<�#a<l�`<��`<�b`<�,`<`<b�_<��_<O�_<�`<�9`<Ts`<�`<��`<�6a<pa<��a<��a<(�a<��a<1�a<z�a<��a<��a<��a<��a<#�a<3�a<��a<��a<��a<��a<Z�a<��a<�a<��a<��a<7�a<.�a<��a<�a<+fa<**a<��`<�`<Gm`<~;`<|`<�`<�`<P`<�;`<�m`<��`<��`<x/a<na<��a<��a<��a<�b<�b<�b<�b<)b<��a<@�a<��a<��a<��a<��a<[�a<��a<��a<�b<�b<~b<Yb<Cb<rb<��a<��a<��a<!ea<&a<�`<��`<�i`<�;`<�`<�`<�`<�+`<-T`<��`<�`<
a<+Ka<��a<]�a<��a<h�a<b<�b<b<�b<Ib<��a<H�a<E�a<��a<��a<Y�a<x�a<+�a<�a<�b<�b<�b<�b<�b<@�a<��a<��a<݊a<Pa<Ha<�`<��`<W`<-`<�`<�`<�`<T4`< a`<��`<��`<�a<�Za<��a<��a<��a<��a<�
b<Mb<�b<rb< �a<�a<��a<�a<N�a<��a<Q�a<�a<A�a<��a<� b<�b<�b<�
b<�b<�a<2�a<��a<oa<Y1a<��`<��`<�n`<X;`<w`<� `<��_<�`<2`<�b`<��`<��`<�a<�[a<Őa<��a<��a<�a<��a<[�a<v�a<��a<�a<��a<)�a<_�a<��a<=�a<��a<��a<B�a<}�a<e�a<v�a<��a<A�a<��a<��a<'�a<�sa<�;a<�`<w�`<�x`<2>`<s`<V�_<��_<]�_<�_<
&`<1[`<W�`<��`<�a<Wa<��a<��a<�a<y�a<��a<�a<��a<�a<.�a<��a<��a<k�a<_�a<I�a<��a<��a<��a<��a<Q�a<�  �  p�a<��a<e�a<s�a<W�a<^�a<ba<j(a<��`<��`<5j`<z4`<�`<1�_<C�_<�_<�`<�A`<iz`<�`<��`<(;a<�sa<��a<��a<�a<��a<%�a<g�a<��a<K�a<4�a<��a<E�a<�a<H�a<��a<�a<3�a<N�a<B�a<��a<��a<-�a<��a<��a<l�a<R�a<Tja<,/a<`�`<��`<�t`<�C`<1 `<q`<g`< `<�C`<^u`<i�`<��`<�4a<Fra<�a<*�a<{�a<�b<4b<b<�b<�b<��a<��a<�a<��a<��a<��a<t�a<S�a<3�a<��a<�b<Ob<0b<b<4b<��a<k�a<��a<�ia<t+a<6�`<��`<�q`<�C`<�$`<H`<�`<i4`<.\`<�`<��`<�a<�Oa<��a<k�a<��a<��a<b<�b<3b<�
b<,b<6�a<T�a<��a<��a<I�a<9�a<��a<�a<��a<^ b<	b<�b<�b<�b<j�a<��a<�a<��a<�Ta<�a<`�`<-�`<�^`<�5`<�`</`<i`<�<`<�h`<Р`<��`<� a<t_a<`�a<f�a<��a<��a<j
b<Bb<�	b<gb<`�a<��a<]�a<-�a<�a<��a<G�a<h�a<��a<��a<A�a<Vb<[
b<#
b<�b<��a<��a<��a<Csa<Z6a<��`<5�`<lv`<hC`<,`<�	`<�`<j`<%:`<j`<D�`<��`<�#a<�_a<�a<��a<i�a<x�a<M�a<��a<�a<�a<'�a<��a<��a<c�a<�a<
�a<�a<Y�a<��a<��a<-�a<G�a<��a<�a<��a<��a<�a<{wa<�?a<Wa<��`<�`<�E`<�`<�_<C�_<)�_<�`<	.`<�b`<��`<��`<� a<[a<��a<�a<f�a<��a<�a<B�a<��a<��a<��a<��a<%�a<V�a<�a<,�a<ҹa<��a<W�a<l�a<��a<�  �  ��a<��a<��a<��a<��a<X�a<�la<�5a<��`<R�`<`<[K`<�#`<`<C`<�`<�,`<1X`<Ɏ`<��`<Ka<�Ga<�}a<�a<��a<��a<o�a<
�a<��a<��a<@�a<T�a<�a<��a<@�a<=�a<��a<C�a<�a<��a<�a<��a<M�a<��a<��a<��a<��a<8�a<�ua<@=a<, a<��`<^�`<�Z`<,9`<e'`<X'`<;9`<A[`<J�`<��`<�a<Ca<
~a<C�a<��a<��a<vb<'b<�b<�b<��a<��a<��a<��a<��a<��a<��a<��a<a�a<�a<Z�a<��a<fb<�b<�b<Pb<��a<��a<U�a<�ua<�:a<��`<Ͼ`<݇`<�[`<=>`<E1`<�6`<M`<?s`<.�`<(�`< a<Z]a<��a<��a<��a<b<�b<�b<�b<Rb<>�a<>�a<��a<K�a<2�a<*�a<��a<D�a<�a<^�a<�a<# b<�	b<Tb<(b<~b<��a<z�a<i�a<�aa<�$a<��`<�`<�u`<�M`<�5`<4.`<9`<�T`<I`<5�`<��`<R0a<la<z�a<��a<�a<b<<
b<)
b<Db<��a<V�a<��a<��a<l�a<Y�a<|�a<�a<��a<\�a<�a<
�a<_�a<�b<�b<1b<��a<.�a<ܰa<�~a<mDa<�a<v�`<�`<�Z`<&7`<~#`<�!`<�1`<�Q`<�`<Է`<��`<`2a<�ka<J�a<Q�a<��a<��a<C�a<��a<w�a<:�a<�a<"�a<!�a<D�a<��a<1�a<-�a<h�a<}�a<O�a<�a<\�a</�a<��a<��a<��a<�a<D�a<2La<`a<$�`<��`<1\`<�/`<�`<;`<	`<@`<E`<�w`<`�`<��`<.a<�ea<ڔa<˸a<��a<4�a<�a<��a<=�a<�a<�a<?�a<�a<�a<��a<��a<q�a<��a<�a<#�a<��a<�  �  ��a<K�a<A�a<c�a<��a<~�a<�|a<�Ia<xa<�`<��`<uo`<�J`<4`<�-`<|8`<$S`<�{`<l�`<��`<�"a<![a<(�a<)�a<��a<z�a<��a<��a<��a<��a<߸a<0�a<؛a<`�a<o�a<	�a<��a<��a<��a<v�a<q�a<F�a<	�a<�a<��a<��a<2�a<��a<[�a<�Ra<a<��`<�`<�`<M``<�O`<�O`<�``<��`<t�`<Z�`<&a<+Ya<�a<*�a<��a<g�a<	b<�
b<b<�a<��a<��a<�a<Q�a<��a<k�a<��a< �a<ûa<^�a<t�a<��a<��a<�b<xb<�b<1�a<`�a<8�a<��a<�Qa</a<	�`<ݪ`<��`<�e`<�Y`<�^`<�s`<��`<�`<X�`<�8a<!ra<4�a<G�a<S�a<]b<�b< b<\b<��a<�a<��a<��a<��a<��a<�a<�a<��a<��a<:�a<��a<��a<��a<
b<�b<Xb<��a<��a<��a<2va<\=a<�a<��`< �`<�t`<�]`<�V`<�``<�z`<��`<��`<xa<�Ga<za<ɰa<�a<�a<�b<�b<�b<9�a<]�a<��a<��a<�a<E�a<��a<E�a<��a<�a<D�a<��a<i�a<��a<d�a<b<8b<��a<~�a<P�a<G�a<Za<xa<r�`<ԭ`<�`<G^`<�K`<J`<�X`<(w`<�`<7�`<=a<�Ha<�}a<3�a<�a<Y�a<��a<�a<��a<��a<%�a<#�a<��a<٘a<_�a<_�a<=�a<��a<̗a<ڤa<j�a<&�a<��a<s�a<p�a<R�a<%�a<жa< �a< _a<y'a<�`<ղ`<(`<}U`<<9`<�,`<:1`< F`<�i`<��`<��`<�	a<�Ba<�va<q�a<A�a<�a<3�a<H�a<u�a<��a<Q�a<a�a<E�a<��a<z~a<�{a<~a<�a<�a<��a<�a<i�a<�  �  b�a<��a<�a<��a<��a<v�a< �a<�ba<�/a<*�`<��`<L�`<�{`<�g`<6b`<�k`<��`<k�`<��`<�
a<�?a<�ra<0�a<��a<a�a<��a<M�a<6�a<�a<�a<��a<'�a<�sa<=fa<�^a<&^a<da<�pa<��a<��a<�a<�a<��a<��a<��a<�a<��a<e�a<��a<�ma<a:a<�a<��`<M�`<��`<݃`<�`<+�`<P�`<��`<�	a<?a<�ta<ԥa<t�a<��a<b<f	b<Qb<q�a<�a<��a<��a<-�a<��a<k�a<�}a<M~a<��a<%�a<��a<ٻa<��a<F�a<��a<Kb<v
b<b<��a<��a<�a<.na<|9a<�a<A�`<(�`<��`<@�`<��`<��`<�`<��`<#a<�Wa<��a<�a<��a<��a<M	b<)b<Yb<��a<`�a<��a<{�a<�a<�a<��a<�}a<ǀa<D�a<��a<k�a<:�a<��a<��a<�b<i
b<�b<4�a<��a<ܼa<%�a<�[a<�&a<��`<��`<�`<B�`<<�`<.�`<«`<��`<�`<f0a<ea<5�a<��a<��a<��a<1b<"b<\�a<y�a<��a<�a<��a<e�a<�a<�ya<]xa<e}a<�a<˙a<Ѯa<��a<.�a<�a<��a<�b<��a<��a<�a<m�a<�ta<�?a<N
a<��`<&�`<��`<�`<;~`<��`<Ѧ`<d�`<��`<40a<�ca<��a<��a<*�a<�a<��a<u�a<H�a<��a<u�a<�a<��a<?oa<$ba<�[a<�[a<?ba<0oa<+�a<ϖa<�a<:�a<.�a<?�a<��a<�a<	�a<��a<9va<�Ca<�a<z�`<��`<�`<Kl`<&a`<	e`<�w`<ۗ`<d�`<?�`<�(a<V\a<{�a<��a<��a<�a<��a<��a<��a<[�a<{�a<Aa<�ja<�Za<oPa<�La<�Oa<�Ya<ia<8}a<Z�a<`�a<�  �  !�a<6�a<��a<��a<2�a<=�a<R�a<�}a<QQa<H#a<d�`<J�`<-�`<��`<ǝ`<4�`<?�`<R�`<�a<41a<�_a<:�a<�a<i�a<��a<r�a<��a<��a<�a<�a<�xa<�[a<{Ca<�1a<�'a<�&a<,.a<(>a<oUa<ra<Αa<n�a<�a<r�a<v�a<f�a<V�a<G�a<�a<��a<^a<01a<�a<��`<��`</�`<n�`<��`<?�`<�	a<�4a<�ca<?�a<�a<
�a<�a<b<�b<��a<��a<��a<��a<̐a<�ta<�]a<�Ma<Fa<�Fa<�Pa<Nba<�za<��a<��a<��a<�a<b<�	b<�b<o�a<��a<��a<u�a<h_a<M2a<�	a<�`<4�`<��`<��`<D�`<��`<7 a<�Ka<=za<R�a<��a<K�a<�b<2b<�b<X�a<E�a<��a<¦a<W�a<�ma<�Xa<*Ka<SFa<Ja<XVa<vja<��a<��a<`�a<>�a<��a<Ub<�	b<�b<c�a<�a<�a<A}a<�Na<y"a<��`<P�`<7�`<��`<��`< �`<�a<X*a<Wa<�a<��a<��a<f�a<�b<b<��a<��a<��a<׵a<��a<3ya<`a<sMa<�Ba<�@a<sGa<tVa<�la<-�a<��a<�a<W�a<X�a<� b<Eb<��a<��a<̻a<�a<wca<�4a<8	a<��`<��`<H�`<��`<�`<��`<��`<�'a<�Ta<��a<��a<�a<��a<�a<��a<��a<^�a<g�a<�a<?ra<5Ua<U=a<�,a<$a<D$a<@-a<\>a<Va<�ra<�a<��a<��a<�a<��a<��a<��a<��a<ߎa<8ca<�4a<a<��`<̼`<{�`<��`<�`<]�`<V�`<��`<"a<$Ka<�wa<c�a<x�a<��a<��a<C�a<��a<p�a<��a<�ua<)Wa<Z<a<X'a< a<Da<%a<�%a<:a<hTa<�ra<�a<�  �  -�a<��a<t�a<e�a<@�a<�a<*�a<��a<sa<RLa<W'a<ha<�`<j�`<^�`<��`<8�`<7a<32a<�Xa<�a<��a<;�a<��a<%�a<U�a<��a<��a<��a<�va<cPa<�,a<a<��`<,�`<w�`<��`<�a<U#a<�Fa<�ma<[�a<��a<8�a<H�a<!�a<��a<w�a<!�a<V�a<T�a<~\a<�9a<�a< a<��`<��`<?	a<�a<�<a<aa<��a<��a<��a<��a<b<�b<�b<)�a<��a<��a<{�a<!fa<JCa<�&a<�a<�a<5
a<Xa<P,a<�Ja<�na<b�a<$�a<��a<C�a<�b<�	b<� b<Q�a<0�a<��a<(�a<`a<�=a<�"a<ca<ya<�a<�a<[1a<�Pa<�ua<Ȝa<*�a<��a<��a<�b<^
b<��a<��a<�a<֧a<�a<;[a<
:a<�a<=a<�a<�a<Ka<M6a<�Va<�{a<��a<C�a<^�a<��a<Tb<�b<A�a<��a<�a<��a<�wa<wRa<2a<Ba<
a<�a<$a<(a<�7a<�Xa<�~a<1�a<�a<��a<��a<sb<�b<��a<��a<��a<t�a<yna<�Ia<�*a<�a<7a<�a<a<�a<�:a<�\a<˂a<��a<��a<�a<��a<�b<��a<�a<�a<y�a<��a<`a<];a<}a<a<��`<�`<�a<2a<�1a<�Sa<�ya<�a<��a<�a<��a<��a<�a<V�a<��a<2�a<oa<�Ga<�#a<:a<��`<��`<��`<�`<aa<"&a<�Ia<�oa<�a<�a<.�a<�a<c�a<R�a<�a<r�a<n�a<W[a<�4a<$a<I�`<��`<H�`<�`<��`<a<]"a<�Fa<�ma<Βa<�a<�a<��a< �a<�a<�a<N�a<�va<�Oa<*a<�a<��`<"�`<��`<�`<��`<�a<�&a<-La<Bsa<�  �  �~a<5�a<��a<��a<=�a<�a<�a<�a<�a<Hsa<�Ua<�;a<G(a<�a<�a<Ra<�-a<ZCa<�^a<�}a<W�a<P�a<��a<�a<��a<1�a<��a<��a<<�a<�Sa<;&a<~�`<�`<.�`<�`<�`<ߵ`<R�`<c�`<[a<�Ga<�va<`�a<�a<)�a<��a<��a<��a<��a<=�a<�a<��a<ja<�Ra<�Ba<Z:a<�:a<Da<�Ua<�ma<L�a<8�a<|�a<$�a<�a<�b<�b<5�a<��a<l�a<��a<�fa<�9a<a<��`<�`<u�`<��`<]�`<��`<�a<�Ca<�qa<�a<��a<{�a<��a</	b<�b<��a<�a<D�a<��a<�a<|pa<�Za<�Ka<�Ea<1Ha<SSa<pfa<�a<��a<��a<\�a<c�a<�b<Mb<ab<:�a<��a<I�a<\�a<Ya<^,a<�a<��`<��`<G�`<�`<��`<q a<'a<ISa<i�a<��a<��a<K�a<�b<�	b<1b<��a<u�a<�a<ߞa<��a<�fa<�Ra<cFa<�Ba<�Ga<�Ua<�ja<��a<�a<��a<��a<k�a<#b<�b<��a<��a<��a<��a<�ra<RDa<�a<��`<�`<�`<
�`<�`<��`<�a<m/a<u\a<+�a<��a<��a<��a<t�a<b<O�a<i�a<]�a<k�a<|�a<�ka<�Ra<�@a<r6a<5a<k<a<
La<�ba</~a<W�a<�a<��a<�a<��a<��a<��a<��a<S�a<Bxa<�Ia<a<��`<��`<ܴ`<|�`<B�`<�`<��`<X�`<�a<La<�xa<�a<a�a<;�a<�a<��a<��a<U�a<�a<�a<`a<�Da<#.a<a<�a<�a<Y%a<#8a<FQa<�na<��a<��a<��a<��a<H�a<)�a<��a<<�a<��a<yVa<(a<L�`<��`<��`<��`<V�`<K�`<��`<�`<�`<�#a<�Qa<�  �  da<_�a<��a<�a<[�a<n�a<M�a<��a<�a<S�a<�~a<2ka<]\a<tSa<1Qa<�Ua<�`a<lqa<��a<V�a<��a<M�a<.�a<"�a<N�a<��a<�a<K�a<=da<1a<��`<��`<W�`<l�`<�q`<^o`<�{`<��`<K�`<)�`<"a<�Wa<�a<l�a<��a<{�a<#�a<K�a<4�a<S�a<K�a<��a<k�a<�a<�wa<�qa<Sra<�ya<+�a<��a<��a<8�a<Y�a<��a<Ob<b<Kb<r�a<��a<�a<nva<"Ba<a<x�`<��`<M�`<��`<��`<?�`<x�`<��`<�a<9Na<P�a<��a<��a<��a<Fb<b<�b<P�a<��a<=�a<�a<�a<@�a<��a<N}a<Ga<Շa<r�a<٩a<��a<n�a<��a<f b<�
b<"b<��a<o�a<��a<u�a<�fa<2a<��`<��`<�`<�`<��`<:�`<��`<��`<��`<�+a<6`a<�a<	�a<��a<j�a<�b<�	b< b<(�a<��a<��a<�a<��a<��a<<}a<oza<K~a<ƈa<Ԙa<O�a<^�a<��a<��a< b<>b<�b<D�a<��a<��a<��a<�Oa<a<:�`<�`<@�`<�`<��`<
�`<�`<x�`<5a<�6a<Jka<[�a<B�a<�a<L�a<[b<��a<�a<p�a<��a<�a<�a<܃a<�ua<�ma<�la<�qa<�}a<��a<��a<Y�a<��a<[�a<i�a<��a<Q�a<�a<�a<Ջa<$Za<�$a<��`<�`<X�`<{`<m`<�m`<�}`<��`<�`<��`<�(a<;\a<�a<۱a<��a<�a<N�a<��a<}�a<h�a<T�a<�a<ra<�`a< Ua<Pa<�Qa<�Ya<ha<9{a<��a<J�a<~�a<��a<��a< �a<��a<�a<�a<�ha<6a<a<��`<|�`<}`<
f`<�]`<}d`<z`<Z�`<��`<��`<�0a<�  �  nKa<j~a<ݧa<!�a<E�a<��a<��a<i�a<X�a<2�a<̠a<��a<�a<Ła<!�a<��a<p�a<��a<`�a<Ѹa<��a<��a<w�a<W�a<�a<�a<�a<~a<cJa<�a<��`<ѡ`<�s`<xQ`<>`<;`<�H`<mf`<8�`<��`<  a<~;a<Tsa<E�a<��a<��a<��a<��a<��a<<�a<��a<��a<j�a<�a<g�a<l�a<�a<��a<��a<��a<d�a<��a<��a<� b<�b<Tb<K�a<�a<8�a<��a<�Za<� a<N�`<�`<Ӈ`<�i`<�Z`<�\`<�n`<j�`<��`<�`<I.a<�ga<ߜa<��a<i�a<vb<�b<nb<�b<��a<�a<�a<��a<��a<��a<?�a<ʭa<ѳa<O�a<��a<�a<��a<A�a<�	b<�b<�b<�a<L�a<N�a<n�a<xIa<�a<R�`<b�`<}`<�c`</Z`<�a`<7y`<�`<��`<�a<-Ba<pza<�a<%�a<�a<�b< b<�b<��a<d�a<��a<�a<O�a<B�a<��a<k�a<F�a<��a<"�a<'�a<��a<��a<1�a<Yb<{b<u�a<��a<��a<V�a<�ia<�0a<�`<-�`<^�`<Im`<Y`<'U`<b`<�~`<_�`<��`<�a<Oa<��a<�a<!�a<��a<b<`b<��a<V�a</�a<�a<�a<��a<]�a<��a<V�a<�a<	�a<A�a<J�a<��a<f�a<��a<��a<��a<U�a<��a<s�a<�ua<�>a<ha<��`<|�`<{g`<XH`<�8`< :`<�K`<�l`<��`<�`<�a<�Aa<Bva<o�a<��a<A�a<��a<�a<�a<��a<�a<��a<��a<�a<ςa<�~a<�a<Ņa<�a<�a<3�a<g�a<��a<�a<�a<��a<��a<�a<Ƃa<�Pa<�a<��`<W�`<_s`<L`<�2`<W)`<�0`<�H`<�n`<՟`<�`<�a<�  �  `7a<yna<�a<]�a<��a<��a<k�a<��a<��a<��a<,�a<�a<��a<d�a<^�a<�a<��a<n�a<��a<B�a<��a<��a< �a<�a<��a<V�a<<�a<?ma<b5a<��`<��`<��`<*O`<�*`<�`<|`<V!`<�@`<qn`<Ϧ`<�`<�$a<�`a<��a<M�a<��a<��a<@�a<��a< �a< �a<��a<M�a<��a<��a<q�a<=�a<`�a<��a<��a<�a<V�a<s�a<ab<{b<|b<[�a<�a<�a<�~a<bDa<+a<��`<��`<Ab`<#B`<32`<E4`<�G`<{k`<s�`<B�`<�a<hRa<��a<Y�a<S�a<��a<�
b<ub<�b<�b<��a<��a<�a<_�a<��a<�a<��a<��a<W�a<}�a<:�a<��a<	b<�b<<b<sb<��a<��a<ʣa<�ma<�1a<��`<n�`<̀`<�V`<�;`<�1`<�9`<�R`<{`<��`<"�`<�)a<]fa<�a<7�a<F�a</b<�b<;b<b<��a<h�a<n�a<��a<��a<?�a<��a<��a<��a<��a<y�a<^�a<2�a<Lb<�b<@b<��a<�a<3�a<}�a<�Ta<ba<��`<�`<�k`<nF`<�0`<�,`<�:`<�X`<��`<Ҽ`<��`<.8a<�ra<q�a<��a<O�a<��a<�b<�b<8�a<q�a<0�a<��a<��a<��a<��a<v�a<��a<(�a<��a<��a<z�a<��a<�a<��a<	�a<g�a<��a<M�a<tca< (a<��`<@�`<q`<�A`<� `<F`<�`<�$`<�G`<�w`<:�`<�`<P,a<�da<3�a<��a<G�a<�a< �a<��a<@�a<��a<Z�a<
�a<�a<��a<'�a<֢a<æa<��a<ӷa<N�a<|�a<��a<�a<q�a<w�a<��a<|�a<Gsa<=a<� a<��`<z�`<�O`<�%`<�
`<� `<�`<:"`<�J`<�`<y�`<��`<�  �  X*a<�ca<�a<ڸa<��a<��a<��a<��a<��a<4�a<��a<F�a<�a< �a<t�a<I�a<��a<�a<x�a<��a<?�a<��a<��a<E�a<�a<I�a<͓a<&ba<�'a<)�`<ʧ`<vk`<	8`<�`<��_<��_<�`<�(`<3X`<ْ`<��`<�a<~Ta<�a<;�a<��a<��a<��a<z�a<6�a<a�a<D�a<��a<��a<��a<R�a<+�a<o�a<��a<��a<��a<��a<�b<tb<_b<�b<��a<5�a<��a<�ra<�5a<��`<��`<|z`<�J`<�(`<@`<O`</`<-T`<�`<(�`<�a<�Da<8�a<��a<�a<��a<�	b<�b<db<�
b<^b<i�a<]�a<L�a<5�a<��a<K�a<��a<��a<7�a<�a<b<mb<�b<Eb<�b<��a<E�a<��a<aa<"a<��`<�`<,j`<�>`<"`<�`<�`<P:`<@d`<��`<��`<a<RYa<��a<_�a<��a<?�a<�b<�b<b<�b<��a<��a<�a<y�a<��a<��a<�a<��a<��a<N�a<�a<�b<�b<�b<tb<u�a<��a<Ǵa<f�a<QGa<�a<��`<Ј`<�T`<�-`<�`<�`<!`<�@`<To`<ڨ`<b�`<I)a<�fa<Μa<��a<��a<��a<eb<Ob<Nb<��a<��a<O�a<��a<��a<h�a<d�a<��a<��a<J�a<��a< �a<Q�a<3�a<�a<i�a<�a<ӹa<��a<�Wa<�a<��`<��`<[`<9*`<�`<U�_<��_<�`<G0`<tb`< �`<[�`<ga<�Ya<u�a<S�a<z�a<�a<��a<}�a<^�a<^�a<��a<V�a<ʾa<B�a<8�a<��a<k�a<p�a<��a<&�a<��a<
�a<��a<z�a<��a<V�a<�a<ia<c0a<Z�`<�`<�p`<69`<�`<$�_<��_</�_<�	`<	4`<�j`<:�`<��`<�  �  �%a<`a<0�a<��a<��a<��a<��a<��a<��a<��a<�a<a�a<��a<#�a<��a<Z�a<]�a<��a<��a<��a<��a<��a<w�a<'�a<��a<ܷa<��a<!^a<�"a<p�`<V�`<d`<�/`<P	`<�_<��_<!�_<� `<�P`<�`<��`<ua<)Pa<��a<��a<��a<��a<�a<��a<r�a<��a<�a<C�a<"�a<��a<��a<a�a<g�a<y�a<C�a<��a<nb<9	b<�b<�b<Vb<'�a<��a<U�a<Sna<�0a<��`<4�`<�r`<{B`< `<�`<�`<Z&`<L`<|`<��`<�`<�?a<|a<j�a<��a<)�a<�	b<�b<b<Yb<,b<��a<$�a<��a<C�a<��a<y�a<^�a<�a<��a<�b<b<qb<�b<hb<�b<`�a<j�a<̕a<�\a<�a<��`<Ú`<cb`<?6`<B`<�`<`<�1`<b\`<z�`<��`<�a<�Ta<��a<t�a<��a<&�a<�b<�b<b<�	b<Gb<I�a<:�a<M�a<�a<�a<!�a<��a<j�a<��a<"b<M	b<[b<fb<Wb<�a<��a<��a<b~a<�Ba<Aa<n�`<c�`<�L`<%`<`<
`<L`<�8`<�g`<�`<N�`<�#a<\ba<O�a<��a<��a<�a<�b<�b<�b<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<5�a<)�a<��a<JSa<Ya<��`<ŏ`<�S`<)"`<��_<��_<��_<`<7(`<[`<��`<��`<xa<zUa<B�a<бa<��a<��a<0�a<,�a<��a<+�a<��a<�a<o�a<N�a<��a<��a<G�a<��a<	�a<��a<��a<�a<��a<��a<��a<6�a<�a<Nea<�+a<��`<��`<�i`<o1`<N`<`�_<5�_<d�_<�`<-,`<�c`<��`<7�`<�  �  X*a<�ca<�a<ڸa<��a<��a<��a<��a<��a<4�a<��a<F�a<�a< �a<t�a<I�a<��a<�a<x�a<��a<?�a<��a<��a<E�a<�a<I�a<͓a<&ba<�'a<)�`<ʧ`<vk`<	8`<�`<��_<��_<�`<�(`<3X`<ْ`<��`<�a<~Ta<�a<;�a<��a<��a<��a<z�a<6�a<a�a<D�a<��a<��a<��a<R�a<+�a<o�a<��a<��a<��a<��a<�b<tb<_b<�b<��a<5�a<��a<�ra<�5a<��`<��`<|z`<�J`<�(`<@`<O`</`<-T`<�`<(�`<�a<�Da<8�a<��a<�a<��a<�	b<�b<db<�
b<^b<i�a<]�a<L�a<5�a<��a<K�a<��a<��a<7�a<�a<b<mb<�b<Eb<�b<��a<E�a<��a<aa<"a<��`<�`<,j`<�>`<"`<�`<�`<P:`<@d`<��`<��`<a<RYa<��a<_�a<��a<?�a<�b<�b<b<�b<��a<��a<�a<y�a<��a<��a<�a<��a<��a<N�a<�a<�b<�b<�b<tb<u�a<��a<Ǵa<f�a<QGa<�a<��`<Ј`<�T`<�-`<�`<�`<!`<�@`<To`<ڨ`<b�`<I)a<�fa<Μa<��a<��a<��a<eb<Ob<Nb<��a<��a<O�a<��a<��a<h�a<d�a<��a<��a<J�a<��a< �a<Q�a<3�a<�a<i�a<�a<ӹa<��a<�Wa<�a<��`<��`<[`<9*`<�`<U�_<��_<�`<G0`<tb`< �`<[�`<ga<�Ya<u�a<S�a<z�a<�a<��a<}�a<^�a<^�a<��a<V�a<ʾa<B�a<8�a<��a<k�a<p�a<��a<&�a<��a<
�a<��a<z�a<��a<V�a<�a<ia<c0a<Z�`<�`<�p`<69`<�`<$�_<��_</�_<�	`<	4`<�j`<:�`<��`<�  �  `7a<yna<�a<]�a<��a<��a<k�a<��a<��a<��a<,�a<�a<��a<d�a<^�a<�a<��a<n�a<��a<B�a<��a<��a< �a<�a<��a<V�a<<�a<?ma<b5a<��`<��`<��`<*O`<�*`<�`<|`<V!`<�@`<qn`<Ϧ`<�`<�$a<�`a<��a<M�a<��a<��a<@�a<��a< �a< �a<��a<M�a<��a<��a<q�a<=�a<`�a<��a<��a<�a<V�a<s�a<ab<{b<|b<[�a<�a<�a<�~a<bDa<+a<��`<��`<Ab`<#B`<32`<E4`<�G`<{k`<s�`<B�`<�a<hRa<��a<Y�a<S�a<��a<�
b<ub<�b<�b<��a<��a<�a<_�a<��a<�a<��a<��a<W�a<}�a<:�a<��a<	b<�b<<b<sb<��a<��a<ʣa<�ma<�1a<��`<n�`<̀`<�V`<�;`<�1`<�9`<�R`<{`<��`<"�`<�)a<]fa<�a<7�a<F�a</b<�b<;b<b<��a<h�a<n�a<��a<��a<?�a<��a<��a<��a<��a<y�a<^�a<2�a<Lb<�b<@b<��a<�a<3�a<}�a<�Ta<ba<��`<�`<�k`<nF`<�0`<�,`<�:`<�X`<��`<Ҽ`<��`<.8a<�ra<q�a<��a<O�a<��a<�b<�b<8�a<q�a<0�a<��a<��a<��a<��a<v�a<��a<(�a<��a<��a<z�a<��a<�a<��a<	�a<g�a<��a<M�a<tca< (a<��`<@�`<q`<�A`<� `<F`<�`<�$`<�G`<�w`<:�`<�`<P,a<�da<3�a<��a<G�a<�a< �a<��a<@�a<��a<Z�a<
�a<�a<��a<'�a<֢a<æa<��a<ӷa<N�a<|�a<��a<�a<q�a<w�a<��a<|�a<Gsa<=a<� a<��`<z�`<�O`<�%`<�
`<� `<�`<:"`<�J`<�`<y�`<��`<�  �  nKa<j~a<ݧa<!�a<E�a<��a<��a<i�a<X�a<2�a<̠a<��a<�a<Ła<!�a<��a<p�a<��a<`�a<Ѹa<��a<��a<w�a<W�a<�a<�a<�a<~a<cJa<�a<��`<ѡ`<�s`<xQ`<>`<;`<�H`<mf`<8�`<��`<  a<~;a<Tsa<E�a<��a<��a<��a<��a<��a<<�a<��a<��a<j�a<�a<g�a<l�a<�a<��a<��a<��a<d�a<��a<��a<� b<�b<Tb<K�a<�a<8�a<��a<�Za<� a<N�`<�`<Ӈ`<�i`<�Z`<�\`<�n`<j�`<��`<�`<I.a<�ga<ߜa<��a<i�a<vb<�b<nb<�b<��a<�a<�a<��a<��a<��a<?�a<ʭa<ѳa<O�a<��a<�a<��a<A�a<�	b<�b<�b<�a<L�a<N�a<n�a<xIa<�a<R�`<b�`<}`<�c`</Z`<�a`<7y`<�`<��`<�a<-Ba<pza<�a<%�a<�a<�b< b<�b<��a<d�a<��a<�a<O�a<B�a<��a<k�a<F�a<��a<"�a<'�a<��a<��a<1�a<Yb<{b<u�a<��a<��a<V�a<�ia<�0a<�`<-�`<^�`<Im`<Y`<'U`<b`<�~`<_�`<��`<�a<Oa<��a<�a<!�a<��a<b<`b<��a<V�a</�a<�a<�a<��a<]�a<��a<V�a<�a<	�a<A�a<J�a<��a<f�a<��a<��a<��a<U�a<��a<s�a<�ua<�>a<ha<��`<|�`<{g`<XH`<�8`< :`<�K`<�l`<��`<�`<�a<�Aa<Bva<o�a<��a<A�a<��a<�a<�a<��a<�a<��a<��a<�a<ςa<�~a<�a<Ņa<�a<�a<3�a<g�a<��a<�a<�a<��a<��a<�a<Ƃa<�Pa<�a<��`<W�`<_s`<L`<�2`<W)`<�0`<�H`<�n`<՟`<�`<�a<�  �  da<_�a<��a<�a<[�a<n�a<M�a<��a<�a<S�a<�~a<2ka<]\a<tSa<1Qa<�Ua<�`a<lqa<��a<V�a<��a<M�a<.�a<"�a<N�a<��a<�a<K�a<=da<1a<��`<��`<W�`<l�`<�q`<^o`<�{`<��`<K�`<)�`<"a<�Wa<�a<l�a<��a<{�a<#�a<K�a<4�a<S�a<K�a<��a<k�a<�a<�wa<�qa<Sra<�ya<+�a<��a<��a<8�a<Y�a<��a<Ob<b<Kb<r�a<��a<�a<nva<"Ba<a<x�`<��`<M�`<��`<��`<?�`<x�`<��`<�a<9Na<P�a<��a<��a<��a<Fb<b<�b<P�a<��a<=�a<�a<�a<@�a<��a<N}a<Ga<Շa<r�a<٩a<��a<n�a<��a<f b<�
b<"b<��a<o�a<��a<u�a<�fa<2a<��`<��`<�`<�`<��`<:�`<��`<��`<��`<�+a<6`a<�a<	�a<��a<j�a<�b<�	b< b<(�a<��a<��a<�a<��a<��a<<}a<oza<K~a<ƈa<Ԙa<O�a<^�a<��a<��a< b<>b<�b<D�a<��a<��a<��a<�Oa<a<:�`<�`<@�`<�`<��`<
�`<�`<x�`<5a<�6a<Jka<[�a<B�a<�a<L�a<[b<��a<�a<p�a<��a<�a<�a<܃a<�ua<�ma<�la<�qa<�}a<��a<��a<Y�a<��a<[�a<i�a<��a<Q�a<�a<�a<Ջa<$Za<�$a<��`<�`<X�`<{`<m`<�m`<�}`<��`<�`<��`<�(a<;\a<�a<۱a<��a<�a<N�a<��a<}�a<h�a<T�a<�a<ra<�`a< Ua<Pa<�Qa<�Ya<ha<9{a<��a<J�a<~�a<��a<��a< �a<��a<�a<�a<�ha<6a<a<��`<|�`<}`<
f`<�]`<}d`<z`<Z�`<��`<��`<�0a<�  �  �~a<5�a<��a<��a<=�a<�a<�a<�a<�a<Hsa<�Ua<�;a<G(a<�a<�a<Ra<�-a<ZCa<�^a<�}a<W�a<P�a<��a<�a<��a<1�a<��a<��a<<�a<�Sa<;&a<~�`<�`<.�`<�`<�`<ߵ`<R�`<c�`<[a<�Ga<�va<`�a<�a<)�a<��a<��a<��a<��a<=�a<�a<��a<ja<�Ra<�Ba<Z:a<�:a<Da<�Ua<�ma<L�a<8�a<|�a<$�a<�a<�b<�b<5�a<��a<l�a<��a<�fa<�9a<a<��`<�`<u�`<��`<]�`<��`<�a<�Ca<�qa<�a<��a<{�a<��a</	b<�b<��a<�a<D�a<��a<�a<|pa<�Za<�Ka<�Ea<1Ha<SSa<pfa<�a<��a<��a<\�a<c�a<�b<Mb<ab<:�a<��a<I�a<\�a<Ya<^,a<�a<��`<��`<G�`<�`<��`<q a<'a<ISa<i�a<��a<��a<K�a<�b<�	b<1b<��a<u�a<�a<ߞa<��a<�fa<�Ra<cFa<�Ba<�Ga<�Ua<�ja<��a<�a<��a<��a<k�a<#b<�b<��a<��a<��a<��a<�ra<RDa<�a<��`<�`<�`<
�`<�`<��`<�a<m/a<u\a<+�a<��a<��a<��a<t�a<b<O�a<i�a<]�a<k�a<|�a<�ka<�Ra<�@a<r6a<5a<k<a<
La<�ba</~a<W�a<�a<��a<�a<��a<��a<��a<��a<S�a<Bxa<�Ia<a<��`<��`<ܴ`<|�`<B�`<�`<��`<X�`<�a<La<�xa<�a<a�a<;�a<�a<��a<��a<U�a<�a<�a<`a<�Da<#.a<a<�a<�a<Y%a<#8a<FQa<�na<��a<��a<��a<��a<H�a<)�a<��a<<�a<��a<yVa<(a<L�`<��`<��`<��`<V�`<K�`<��`<�`<�`<�#a<�Qa<�  �  -�a<��a<t�a<e�a<@�a<�a<*�a<��a<sa<RLa<W'a<ha<�`<j�`<^�`<��`<8�`<7a<32a<�Xa<�a<��a<;�a<��a<%�a<U�a<��a<��a<��a<�va<cPa<�,a<a<��`<,�`<w�`<��`<�a<U#a<�Fa<�ma<[�a<��a<8�a<H�a<!�a<��a<w�a<!�a<V�a<T�a<~\a<�9a<�a< a<��`<��`<?	a<�a<�<a<aa<��a<��a<��a<��a<b<�b<�b<)�a<��a<��a<{�a<!fa<JCa<�&a<�a<�a<5
a<Xa<P,a<�Ja<�na<b�a<$�a<��a<C�a<�b<�	b<� b<Q�a<0�a<��a<(�a<`a<�=a<�"a<ca<ya<�a<�a<[1a<�Pa<�ua<Ȝa<*�a<��a<��a<�b<^
b<��a<��a<�a<֧a<�a<;[a<
:a<�a<=a<�a<�a<Ka<M6a<�Va<�{a<��a<C�a<^�a<��a<Tb<�b<A�a<��a<�a<��a<�wa<wRa<2a<Ba<
a<�a<$a<(a<�7a<�Xa<�~a<1�a<�a<��a<��a<sb<�b<��a<��a<��a<t�a<yna<�Ia<�*a<�a<7a<�a<a<�a<�:a<�\a<˂a<��a<��a<�a<��a<�b<��a<�a<�a<y�a<��a<`a<];a<}a<a<��`<�`<�a<2a<�1a<�Sa<�ya<�a<��a<�a<��a<��a<�a<V�a<��a<2�a<oa<�Ga<�#a<:a<��`<��`<��`<�`<aa<"&a<�Ia<�oa<�a<�a<.�a<�a<c�a<R�a<�a<r�a<n�a<W[a<�4a<$a<I�`<��`<H�`<�`<��`<a<]"a<�Fa<�ma<Βa<�a<�a<��a< �a<�a<�a<N�a<�va<�Oa<*a<�a<��`<"�`<��`<�`<��`<�a<�&a<-La<Bsa<�  �  !�a<6�a<��a<��a<2�a<=�a<R�a<�}a<QQa<H#a<d�`<J�`<-�`<��`<ǝ`<4�`<?�`<R�`<�a<41a<�_a<:�a<�a<i�a<��a<r�a<��a<��a<�a<�a<�xa<�[a<{Ca<�1a<�'a<�&a<,.a<(>a<oUa<ra<Αa<n�a<�a<r�a<v�a<f�a<V�a<G�a<�a<��a<^a<01a<�a<��`<��`</�`<n�`<��`<?�`<�	a<�4a<�ca<?�a<�a<
�a<�a<b<�b<��a<��a<��a<��a<̐a<�ta<�]a<�Ma<Fa<�Fa<�Pa<Nba<�za<��a<��a<��a<�a<b<�	b<�b<o�a<��a<��a<u�a<h_a<M2a<�	a<�`<4�`<��`<��`<D�`<��`<7 a<�Ka<=za<R�a<��a<K�a<�b<2b<�b<X�a<E�a<��a<¦a<W�a<�ma<�Xa<*Ka<SFa<Ja<XVa<vja<��a<��a<`�a<>�a<��a<Ub<�	b<�b<c�a<�a<�a<A}a<�Na<y"a<��`<P�`<7�`<��`<��`< �`<�a<X*a<Wa<�a<��a<��a<f�a<�b<b<��a<��a<��a<׵a<��a<3ya<`a<sMa<�Ba<�@a<sGa<tVa<�la<-�a<��a<�a<W�a<X�a<� b<Eb<��a<��a<̻a<�a<wca<�4a<8	a<��`<��`<H�`<��`<�`<��`<��`<�'a<�Ta<��a<��a<�a<��a<�a<��a<��a<^�a<g�a<�a<?ra<5Ua<U=a<�,a<$a<D$a<@-a<\>a<Va<�ra<�a<��a<��a<�a<��a<��a<��a<��a<ߎa<8ca<�4a<a<��`<̼`<{�`<��`<�`<]�`<V�`<��`<"a<$Ka<�wa<c�a<x�a<��a<��a<C�a<��a<p�a<��a<�ua<)Wa<Z<a<X'a< a<Da<%a<�%a<:a<hTa<�ra<�a<�  �  b�a<��a<�a<��a<��a<v�a< �a<�ba<�/a<*�`<��`<L�`<�{`<�g`<6b`<�k`<��`<k�`<��`<�
a<�?a<�ra<0�a<��a<a�a<��a<M�a<6�a<�a<�a<��a<'�a<�sa<=fa<�^a<&^a<da<�pa<��a<��a<�a<�a<��a<��a<��a<�a<��a<e�a<��a<�ma<a:a<�a<��`<M�`<��`<݃`<�`<+�`<P�`<��`<�	a<?a<�ta<ԥa<t�a<��a<b<f	b<Qb<q�a<�a<��a<��a<-�a<��a<k�a<�}a<M~a<��a<%�a<��a<ٻa<��a<F�a<��a<Kb<v
b<b<��a<��a<�a<.na<|9a<�a<A�`<(�`<��`<@�`<��`<��`<�`<��`<#a<�Wa<��a<�a<��a<��a<M	b<)b<Yb<��a<`�a<��a<{�a<�a<�a<��a<�}a<ǀa<D�a<��a<k�a<:�a<��a<��a<�b<i
b<�b<4�a<��a<ܼa<%�a<�[a<�&a<��`<��`<�`<B�`<<�`<.�`<«`<��`<�`<f0a<ea<5�a<��a<��a<��a<1b<"b<\�a<y�a<��a<�a<��a<e�a<�a<�ya<]xa<e}a<�a<˙a<Ѯa<��a<.�a<�a<��a<�b<��a<��a<�a<m�a<�ta<�?a<N
a<��`<&�`<��`<�`<;~`<��`<Ѧ`<d�`<��`<40a<�ca<��a<��a<*�a<�a<��a<u�a<H�a<��a<u�a<�a<��a<?oa<$ba<�[a<�[a<?ba<0oa<+�a<ϖa<�a<:�a<.�a<?�a<��a<�a<	�a<��a<9va<�Ca<�a<z�`<��`<�`<Kl`<&a`<	e`<�w`<ۗ`<d�`<?�`<�(a<V\a<{�a<��a<��a<�a<��a<��a<��a<[�a<{�a<Aa<�ja<�Za<oPa<�La<�Oa<�Ya<ia<8}a<Z�a<`�a<�  �  ��a<K�a<A�a<c�a<��a<~�a<�|a<�Ia<xa<�`<��`<uo`<�J`<4`<�-`<|8`<$S`<�{`<l�`<��`<�"a<![a<(�a<)�a<��a<z�a<��a<��a<��a<��a<߸a<0�a<؛a<`�a<o�a<	�a<��a<��a<��a<v�a<q�a<F�a<	�a<�a<��a<��a<2�a<��a<[�a<�Ra<a<��`<�`<�`<M``<�O`<�O`<�``<��`<t�`<Z�`<&a<+Ya<�a<*�a<��a<g�a<	b<�
b<b<�a<��a<��a<�a<Q�a<��a<k�a<��a< �a<ûa<^�a<t�a<��a<��a<�b<xb<�b<1�a<`�a<8�a<��a<�Qa</a<	�`<ݪ`<��`<�e`<�Y`<�^`<�s`<��`<�`<X�`<�8a<!ra<4�a<G�a<S�a<]b<�b< b<\b<��a<�a<��a<��a<��a<��a<�a<�a<��a<��a<:�a<��a<��a<��a<
b<�b<Xb<��a<��a<��a<2va<\=a<�a<��`< �`<�t`<�]`<�V`<�``<�z`<��`<��`<xa<�Ga<za<ɰa<�a<�a<�b<�b<�b<9�a<]�a<��a<��a<�a<E�a<��a<E�a<��a<�a<D�a<��a<i�a<��a<d�a<b<8b<��a<~�a<P�a<G�a<Za<xa<r�`<ԭ`<�`<G^`<�K`<J`<�X`<(w`<�`<7�`<=a<�Ha<�}a<3�a<�a<Y�a<��a<�a<��a<��a<%�a<#�a<��a<٘a<_�a<_�a<=�a<��a<̗a<ڤa<j�a<&�a<��a<s�a<p�a<R�a<%�a<жa< �a< _a<y'a<�`<ղ`<(`<}U`<<9`<�,`<:1`< F`<�i`<��`<��`<�	a<�Ba<�va<q�a<A�a<�a<3�a<H�a<u�a<��a<Q�a<a�a<E�a<��a<z~a<�{a<~a<�a<�a<��a<�a<i�a<�  �  ��a<��a<��a<��a<��a<X�a<�la<�5a<��`<R�`<`<[K`<�#`<`<C`<�`<�,`<1X`<Ɏ`<��`<Ka<�Ga<�}a<�a<��a<��a<o�a<
�a<��a<��a<@�a<T�a<�a<��a<@�a<=�a<��a<C�a<�a<��a<�a<��a<M�a<��a<��a<��a<��a<8�a<�ua<@=a<, a<��`<^�`<�Z`<,9`<e'`<X'`<;9`<A[`<J�`<��`<�a<Ca<
~a<C�a<��a<��a<vb<'b<�b<�b<��a<��a<��a<��a<��a<��a<��a<��a<a�a<�a<Z�a<��a<fb<�b<�b<Pb<��a<��a<U�a<�ua<�:a<��`<Ͼ`<݇`<�[`<=>`<E1`<�6`<M`<?s`<.�`<(�`< a<Z]a<��a<��a<��a<b<�b<�b<�b<Rb<>�a<>�a<��a<K�a<2�a<*�a<��a<D�a<�a<^�a<�a<# b<�	b<Tb<(b<~b<��a<z�a<i�a<�aa<�$a<��`<�`<�u`<�M`<�5`<4.`<9`<�T`<I`<5�`<��`<R0a<la<z�a<��a<�a<b<<
b<)
b<Db<��a<V�a<��a<��a<l�a<Y�a<|�a<�a<��a<\�a<�a<
�a<_�a<�b<�b<1b<��a<.�a<ܰa<�~a<mDa<�a<v�`<�`<�Z`<&7`<~#`<�!`<�1`<�Q`<�`<Է`<��`<`2a<�ka<J�a<Q�a<��a<��a<C�a<��a<w�a<:�a<�a<"�a<!�a<D�a<��a<1�a<-�a<h�a<}�a<O�a<�a<\�a</�a<��a<��a<��a<�a<D�a<2La<`a<$�`<��`<1\`<�/`<�`<;`<	`<@`<E`<�w`<`�`<��`<.a<�ea<ڔa<˸a<��a<4�a<�a<��a<=�a<�a<�a<?�a<�a<�a<��a<��a<q�a<��a<�a<#�a<��a<�  �  p�a<��a<e�a<s�a<W�a<^�a<ba<j(a<��`<��`<5j`<z4`<�`<1�_<C�_<�_<�`<�A`<iz`<�`<��`<(;a<�sa<��a<��a<�a<��a<%�a<g�a<��a<K�a<4�a<��a<E�a<�a<H�a<��a<�a<3�a<N�a<B�a<��a<��a<-�a<��a<��a<l�a<R�a<Tja<,/a<`�`<��`<�t`<�C`<1 `<q`<g`< `<�C`<^u`<i�`<��`<�4a<Fra<�a<*�a<{�a<�b<4b<b<�b<�b<��a<��a<�a<��a<��a<��a<t�a<S�a<3�a<��a<�b<Ob<0b<b<4b<��a<k�a<��a<�ia<t+a<6�`<��`<�q`<�C`<�$`<H`<�`<i4`<.\`<�`<��`<�a<�Oa<��a<k�a<��a<��a<b<�b<3b<�
b<,b<6�a<T�a<��a<��a<I�a<9�a<��a<�a<��a<^ b<	b<�b<�b<�b<j�a<��a<�a<��a<�Ta<�a<`�`<-�`<�^`<�5`<�`</`<i`<�<`<�h`<Р`<��`<� a<t_a<`�a<f�a<��a<��a<j
b<Bb<�	b<gb<`�a<��a<]�a<-�a<�a<��a<G�a<h�a<��a<��a<A�a<Vb<[
b<#
b<�b<��a<��a<��a<Csa<Z6a<��`<5�`<lv`<hC`<,`<�	`<�`<j`<%:`<j`<D�`<��`<�#a<�_a<�a<��a<i�a<x�a<M�a<��a<�a<�a<'�a<��a<��a<c�a<�a<
�a<�a<Y�a<��a<��a<-�a<G�a<��a<�a<��a<��a<�a<{wa<�?a<Wa<��`<�`<�E`<�`<�_<C�_<)�_<�`<	.`<�b`<��`<��`<� a<[a<��a<�a<f�a<��a<�a<B�a<��a<��a<��a<��a<%�a<V�a<�a<,�a<ҹa<��a<W�a<l�a<��a<�  �  ��a<8�a<y�a<o�a<ßa<��a<2]a<�1a<�a< �`<��`<F{`<�\`<SJ`<�E`<N`<]d`<��`<�`<��`<�a<�@a<Lla<͐a<��a<h�a<i�a<��a<��a<<�a<D�a<��a<0�a<3�a<U�a<��a<�a<��a<	�a<��a<��a<��a<�a<��a<��a<\�a<��a<��a<Oia<�<a<�a<��`<ñ`<��`<qs`<?f`<f`<�s`<ˎ`<ĳ`<��`<�a<RCa</ra<қa<��a<��a<v�a<��a<�a<~�a<��a<(�a<M�a<��a<��a<��a<:�a<��a<�a<��a<*�a<��a<R�a<K�a</�a<��a<��a<,�a<-�a<ma<>a<Fa<��`<D�`<x�`<>z`<�p`<�t`<�`<��`<��`<��`<r)a<�Ya<o�a<'�a<d�a<;�a<~�a<3�a<G�a<�a<��a<��a<��a<��a<(�a<�a<��a<��a<��a<$�a<A�a<��a<��a<B�a<�a<��a<��a<)�a<:�a<']a<�,a<��`<G�`<�`<@�`<s`<n`<�u`<k�`<�`<��`<�a<f5a<�da<R�a<�a<\�a<T�a<��a<?�a<��a<`�a<��a<_�a< �a<Z�a<��a<�a<��a<5�a<��a<9�a<��a<��a<��a<��a<k�a<��a<w�a<��a<�qa<�Ca<a<��`<Q�`<e�`<iq`<jb`<�``<�l`<��`<Ψ`<�`<Na<C3a<`a<��a<̨a<z�a<��a<��a<��a<�a<F�a<��a<��a<=�a<p�a<�a<d�a<�a<�a<F�a<��a<�a<��a<r�a<��a<ȿa<(�a<D�a<�na<Da<�a<L�`<M�`<O�`<f`<`N`<�D`<�G`<�X`<4v`<�`<��`<"�`<X+a<�Wa<~a<�a<��a<¾a<G�a<2�a<ڿa<q�a<&�a<k�a<,�a<ɢa<͡a<��a<�a<�a<��a<&�a<ſa<�  �  ��a<u�a<7�a<�a<�a<��a<�_a<�4a<�a<��`<M�`<��`<c`<�P`<�K`<hT`<Xj`<?�`<��`<��`<a<FDa<�na<��a<�a<��a<�a<��a<��a<��a<��a<y�a<z�a<�a<�a<N�a<ٯa<Ĵa<��a<��a<��a<f�a<��a<F�a<��a<;�a<0�a<��a<Ola<v@a<,a<O�`<:�`<o�`<�y`<Ol`<�l`<Pz`<��`<D�`<��`<�a<)Ga<Dua<�a<�a<��a<q�a<]�a<��a<4�a<��a<C�a<�a<��a<��a<��a<��a<i�a<C�a<��a<]�a<�a<:�a<-�a<��a<��a<��a<׻a<��a<Mpa<Ba<�a<��`<ڸ`<a�`<��`<�v`<�z`<*�`<S�`<�`<T�`<�-a<w]a<D�a<
�a<��a<��a<D�a<��a<��a<��a<R�a<��a<`�a<��a<��a<��a<��a<��a<2�a<�a<��a<��a<1�a<~�a<��a<1�a<��a<	�a<��a<�`a<�0a<i a<��`<ɪ`<`�`<jy`<�s`<|`<h�`<��`<��`<	a<x9a< ha<ϑa<�a<��a<��a<R�a<@�a<��a<��a<��a<+�a<j�a<:�a<_�a<��a<\�a<J�a<*�a<D�a<��a<S�a<F�a<��a<S�a<��a<�a<��a<�ta<AGa<>a<��`<ȸ`<3�`<�w`<zh`<�f`<�r`<m�`<N�`<��`<�a<7a<�ca<��a<P�a<o�a<��a<a�a<��a<��a<9�a<��a<h�a<]�a<E�a<��a<�a<�a<"�a<�a<�a<3�a<��a<T�a<~�a<�a<J�a<�a<qa<YGa<�a<��`<U�`<�`<�k`<�T`<�J`<N`<_`<�{`<b�`<M�`<N�`<�.a<nZa<�a<k�a<R�a<��a<��a<��a<Z�a<��a<�a<�a<)�a<��a<h�a<u�a<ՠa<��a<��a<��a<5�a<�  �  ��a<��a<��a<��a<��a<5�a<�ga<[>a<Na<�`<��`<ő`<�t`<�c`<�^`<@g`<�{`<ԛ`< �`<��`< a<CMa<va<��a<1�a<��a<�a<c�a<�a<��a<Y�a<E�a<K�a<�a<��a<��a<؟a<ԥa<��a<��a<��a<��a<7�a<X�a<��a<��a<~�a<�a<�ta<~Ja<Ka<c�`<D�`<��`<"�`<H`<s`<ٌ`<�`<s�`<��`<B"a<lQa<�}a<z�a<��a<7�a<��a<��a<��a<��a<=�a<S�a<�a<�a<��a<�a<^�a<��a<��a<Q�a<��a<�a<<�a<��a<��a<��a<��a<��a<��a<ya<�La<Xa<��`<Z�`<�`<l�`<؉`<��`<D�`<>�`<��`<�
a<_9a<ga<#�a<�a<��a<��a<��a<�a<��a<��a<��a<��a<��a<Z�a<��a<׻a<D�a<f�a<b�a<@�a<�a<��a<��a<��a<N�a<��a<��a<��a<��a<�ia<�<a<�a<�`<��`<T�`<^�`<�`<�`<�`<F�`<��`<	a<�Da<qa<�a<�a<��a<��a<T�a<��a<��a<��a<��a<��a<;�a<��a<�a<�a<Z�a<X�a<�a<�a<��a<��a<��a<��a<a�a<��a<8�a<�a<}a<HQa<]"a<��`<��`<\�`<�`<r{`<�y`<m�`<��`<~�`</�`<�a<^Aa<�ka<8�a<Үa<��a<�a<��a<R�a<Y�a<��a<��a<w�a<��a<W�a<ՙa<��a<;�a<��a<��a<��a<3�a<��a<��a<C�a<��a<Q�a<ۘa<xa<%Pa<f#a<Z�`< �`<`�`<s}`<�g`<�]`<a`<3q`<Ռ`<�`<��`<a<y8a<Mba<ͅa<M�a<"�a<0�a< �a<��a<L�a<��a<��a<Z�a<�a<e�a<��a<+�a<~�a<��a<ۡa<��a<�a<�  �  ��a<��a<T�a<n�a<٩a<��a<2sa<(Ma<Y#a<0�`<t�`</�`<,�`<ŀ`<Z|`<8�`<ؗ`<��`<)�`<�a<`1a<W[a<��a<W�a<��a<��a<��a<��a<Ƚa<��a<��a<#�a<��a<�a<��a<c�a<�a<+�a<�a<�a<�a<��a<��a<h�a<��a<~�a<��a<��a<0�a<ZZa<�0a<ma<��`<��`<��`<М`<�`<j�`<;�`<c�`<.
a<�5a<�aa<��a<s�a<%�a<��a<��a<�a<��a<8�a<��a<x�a<�a<��a<��a<ʠa<M�a<�a<߭a<Ӹa<��a<e�a<��a<e�a<��a<��a<��a<�a<7�a<Ԇa<�]a<�2a<�a<��`<��`<G�`<��`<�`<��`<��`<��`<l a<�Ka<2va<�a<��a<�a<��a<�a<P�a<u�a<��a<]�a<ҿa<��a<E�a<�a<��a<{�a<�a<�a<нa<�a<S�a<a�a<��a<��a<��a<��a<	�a<>�a<�xa<�Na<�"a<��`<	�`<��`<��`<��`<�`<�`<(�`<� a<�*a<�Ua<a<�a<��a<9�a<��a<)�a<*�a<��a<��a<�a<Եa<p�a<�a<�a<Лa<��a<��a<��a<ֻa<�a<��a<h�a<��a<G�a<��a<f�a<��a<��a<"aa<�5a<�	a<v�`<x�`<��`<��`<l�`<��`<�`<o�`<~�`<�'a<�Qa<�xa<4�a<`�a<J�a<Y�a<&�a<R�a<��a<>�a<ޤa<Q�a<+�a<0�a<�a<za<q�a<��a<�a<��a<��a<3�a<��a<��a<��a<Z�a<�a<��a<�]a<W4a<�a<��`<�`<(�`<^�`<8{`<_~`<�`<��`<�`<a�`<�a<�Ga<@na<��a<Ȧa<k�a<L�a<l�a<h�a<k�a<�a<v�a<K�a<�ya<�sa<fqa<isa<>ya<f�a<p�a<�a<��a<�  �  �a<2�a<`�a<ùa<��a<e�a<:�a<�_a<�9a<�a<��`<��`<��`<��`<Ţ`<ȩ`<̻`<��`<��`<Ma<�Fa<�la<��a<N�a<T�a<b�a<��a<)�a<��a<�a<C�a<f~a<!pa<�ea<�_a<�_a<rda<�na<�|a<9�a<�a<r�a<r�a<��a<�a<M�a<��a<��a<��a<,na<fHa<q"a<l�`<��`<��`<��`<O�`<��`<f�`<Ka<�&a<8Na<�ua<��a<�a<��a<��a<��a<��a<��a<p�a<@�a<��a<ߙa<H�a<��a<~a<�~a<v�a<!�a<��a<��a<��a<��a<z�a<��a<��a<	�a<��a<��a<�a<sa<�Ka<�%a<�a<_�`<��`<��`<�`<9�`<�`<�a<�;a<�ba<#�a<��a<��a<=�a<��a<��a<Y�a<	�a<�a<[�a<��a<{�a<��a<��a<�~a<��a<��a<q�a<�a<��a<L�a<n�a<4�a<�a<�a<f�a<��a<H�a<E�a<ea<�=a<&a<��`<��`<|�`<�`<��`<��`<5�`<�a<|Da<rka<��a<�a<��a< �a<Z�a<=�a<��a<��a<��a<��a<�a<�a<܀a<Gza<ya<�|a<�a<�a<��a<�a<V�a<�a<��a<��a<��a<}�a<��a<0�a<�ta<tMa<�%a<� a<R�`<��`<�`<��`<&�`<4�`<W�`<�a<�?a<�ea<�a<��a<�a<��a<Y�a<��a<s�a<�a<��a<�a<O{a<�la<Kba<�\a<�\a<�aa<la<�ya<��a<�a<��a<��a<5�a<��a<��a<��a<B�a<�na<yIa<�!a</�`<��`<�`<ϩ`<��`<Q�`<�`<��`<��`<�a<f4a<�Za<�|a<˘a<�a<:�a<Һa<z�a<�a<�a<�a<7va< fa<�Ya<lQa<�Na<�Pa<�Xa<�da<�ta<��a<��a<�  �  ��a<6�a<��a<��a<Ӵa<}�a<$�a<�sa<�Ra<	1a<�a<[�`<��`<��`<b�`<��`<|�`<h�`<�a<8<a<�^a<�a<ƛa<[�a<u�a<h�a<�a<�a<�a<��a<�sa<f^a<La<�>a<7a<p6a<M<a<�Ha<�Za<�pa<��a<i�a<��a<O�a<��a<9�a<��a<+�a<r�a<݃a<ca<@Ba<�#a<�	a<��`<k�`<��`<��`<a<�&a<�Fa<\ia<&�a<��a<�a<-�a<?�a<@�a<�a<��a<�a<��a<��a<^xa<ga<�Za<�Ta<�Ua<]a<�ja<-}a<�a<W�a<��a<��a<*�a<��a<��a<-�a<�a<K�a<h�a<[ha<(Ga<�(a<�a<~ a<��`<_�`<�a<�a<�9a<IZa<M|a<��a<�a<v�a<�a<��a<4�a<��a<&�a<�a<Ԟa<�a<�sa<�ca</Ya<�Ua<PXa<�aa<&qa<�a<��a<��a<��a<3�a<-�a<7�a<��a<��a<4�a<E�a<~a<�[a<�:a<Da<;a<��`<��`<v�`<�a<�"a<�@a<paa<f�a<��a<�a<��a<(�a<e�a<Y�a<x�a<�a<��a<h�a<{a<�ga<�Ya<dQa<�Oa<�Ta<p`a<qa<��a<Ϝa<I�a<O�a<~�a<��a<x�a<l�a<D�a<�a<��a<ha<�Ea<%a<�	a<��`<��`<8�`<y�`<�a<�a<C:a<�Za<|a<R�a<ղa<m�a<
�a<��a<-�a<Y�a<��a<�a<pa<�Ya<�Ga<Z:a<�3a<�3a<�:a<�Ga<zYa<�na<��a<O�a<��a<úa<�a<+�a<2�a<�a<A�a<�`a<F>a<�a<��`<E�`<��`<<�`<��`<��`<]�`<a<7,a<�Ma<oa<I�a<f�a<Ȳa<�a<��a<�a<&�a<ʅa<�na<�Wa<FCa<U3a<�(a<b%a<P(a<2a<�Aa<�Ua<~la<Ӄa<�  �  ��a<��a<��a<��a<s�a<��a<��a<��a<~la<�Oa<Q4a<�a<o
a<]�`<b�`<�a<xa<�#a<7=a<�Ya<Rwa<�a<�a<,�a<�a<Ϳa<�a<J�a<݌a<�qa<aUa<�:a<J$a<�a<E
a<$	a<na<�a<,5a<�Oa<&ma<��a<��a<��a<��a<}�a<�a<'�a<��a<ҙa<�~a<�ba<�Ha<s3a<&$a<Ma<�a<�%a<	6a<�La<�ga<p�a<��a<ؼa<��a<$�a<�a<��a<�a<�a<�a<��a<?ma<ISa<>a</a<�'a<�(a<�1a<vBa<Ya<�sa<Ȑa<۬a<k�a<i�a<��a<��a<b�a<��a<k�a<C�a<��a<>ia<�Oa<~;a<�-a<�'a<*a<�4a<�Fa< ^a<�ya<��a<c�a<<�a<+�a<?�a<��a<��a<�a<��a<�a<�a<�ea<Ma<�9a<�,a<(a<�+a<�7a<;Ja<^ba<~a<�a<��a<��a<D�a<��a<M�a<�a<��a<T�a<a<�za<�^a<�Fa<�3a<O(a<�$a<�)a<�6a<MJa<(ca</a<�a<]�a<E�a<��a<��a<��a<:�a<��a<��a<ԏa<�ra<�Wa<4@a<�.a<�$a<�"a<�(a<7a<�Ka<ea<A�a<��a<.�a<��a<|�a<��a<��a<<�a<)�a<��a<��a<�ea<aJa<43a<"a<va<(a<)a<�,a<�Aa<.[a<wa<��a<1�a<m�a<h�a<��a<?�a<$�a<�a<�a<&ma<�Oa<�4a<�a<�a<�a<�a<ha<]a<d5a<�Oa<�ka<�a<��a<��a<�a<-�a<`�a<A�a<Y�a<�xa<v[a<�>a<�$a<�a<�a<:�`<K�`<�a<
a<R0a<~Ka<Dha<ȃa<e�a<�a<��a<$�a<G�a<>�a<ĉa<�na<�Qa<�5a<�a<Y	a<��`<��`<��`<�a<�a<3a<Oa<9la<�  �  �sa<��a<�a<)�a<4�a<¶a<j�a<��a<j�a<uma<Wa<�Ca<�4a<�+a<�)a<.a<J9a<�Ia<�^a<bva<�a<��a<��a<�a<��a<Q�a<�a<�a<�wa<Wa<�5a<Ea<c�`<��`<��`<+�`<r�`<#�`<�a<.a<;Pa<;sa<ޓa</�a<��a<��a<��a<=�a<9�a<�a<h�a<�a</ma<�[a<fOa<]Ia<�Ia<Qa<�^a<pqa<�a<��a<r�a<��a<\�a<:�a<��a<��a<(�a<�a<��a<Cma<	La<6-a<�a<3a<��`<��`<�a<!a< 4a<�Sa<�ua<:�a<t�a<��a<��a<��a<��a<��a<��a<K�a<t�a<q�a<�ua<ea<�Ya<Ua<�Va<�_a< na<q�a<�a<8�a<K�a<��a<��a<��a<��a<��a<d�a<��a<�a<da<Ca<�%a<la<|�`<�`<F�`<a<2"a<�>a<�_a<z�a<4�a<z�a<�a<c�a<�a<:�a<��a<��a<��a<T�a<��a<�ma<b^a<�Ta<5Ra<�Ua<�`a<�pa<�a<��a<��a<x�a<��a<��a<_�a<Z�a<5�a<}�a<��a<7ua<BSa<�2a<Ka<�a<��`<��`<��`<�a<�$a<HCa<Pda<�a<e�a<U�a<��a<��a<B�a<P�a<��a<��a<r�a<d�a<�na<�[a<[Ma<�Ea<TDa<�Ia<�Ua<fa<={a<��a<k�a<Q�a<&�a<��a<��a<��a<?�a<��a<�sa<�Pa<�.a<�a<�`<��`<��`<��`<�`<
�`<Oa<�/a<�Pa<�qa<��a<Q�a<̷a<3�a<��a<6�a<ǣa<��a<Nwa<�_a<uJa<l9a<�-a<�(a<
*a<R2a<�@a<�Sa<�ia<ۀa<��a<��a<�a<M�a<Q�a<$�a<��a<�va<Va<�3a<�a<O�`<4�`<S�`<��`<\�`<L�`<��`<�a<�0a<�Ra<�  �  2`a<�a<�a<(�a<I�a<ٻa<��a<��a<w�a<ۇa<fva<&ga<�[a<�Ta<Sa<�Va<g_a<�la<<}a<��a<ѡa<!�a<��a<$�a<��a<2�a<�a<�a<ca<:=a<�a<��`<��`<�`<0�`<��`<Ҹ`<��`<y�`<�a<34a<!\a<a<<�a<��a<{�a<q�a<��a<j�a<��a</�a<F�a<�a<��a<�va<\ra<sa<�xa<Ճa<��a<��a<[�a<��a<��a<��a<��a<,�a<��a<��a<M�a<mxa<�Qa<d+a<ua<�`<��`<�`<U�`<��`<��`<a<P4a<8[a<Ӂa<�a<g�a<�a<�a<F�a<M�a<��a<��a<�a<K�a<ӗa<Њa<�a<B~a<�a<��a<�a<<�a<�a<��a<��a<�a<��a<8�a<T�a<r�a<K�a<r�a<�ma<�Fa<� a<��`<��`<x�`<d�`<�`<��`<��`<Ja<�Aa<�ha<|�a<دa<��a<a�a<#�a<S�a<��a<e�a<��a<��a<ݠa<)�a<+�a<�}a<�{a<l~a<��a<:�a<C�a<�a<x�a<�a<��a<��a<M�a<@�a<]�a<��a<�a<e[a<P4a<~a<m�`<�`<p�`<��`<=�`<U�`<��`< "a<EHa<�na<D�a<^�a<M�a<��a<�a<�a<��a<>�a<6�a<��a<q�a<?�a<�ta<�na<ima<{qa<�za<��a< �a<��a<��a<�a<r�a<��a< �a<8�a<֡a<$�a<]a<X5a<�a<��`<��`<��`<�`<��`<�`<��`<l�`<a<e6a<t\a<$a<��a< �a<��a<7�a<��a<űa<��a<ݏa<�}a<�la<,_a<�Ua<�Qa<�Ra<\Ya<vda<dsa<Ȅa<y�a<�a<��a<��a<��a<�a<՞a<��a<�ca<�=a<�a<��`<i�`<`�`<Y�`<_�`<?�`<1�`<q�`<�`<�a<:a<�  �  �Ma<ta<w�a<��a</�a<�a<f�a<�a<��a<��a<j�a<�a<Y|a<wa<�ua<�xa<�a<��a<<�a<L�a<�a<F�a<o�a<`�a<y�a<ˮa<��a<Lva<�Oa<&a<{�`<��`<3�`</�`<1�`<-�`<s�`<Q�`<�`<��`<%a<9Ga<�pa<��a<M�a<{�a<��a<��a<��a<k�a<�a<c�a<I�a<d�a<��a<�a<Õa<��a<	�a<z�a<:�a<��a<�a<`�a<��a<`�a<��a<��a<��a<�a<�ca<=9a<�a<W�`<��`<��`<˧`<:�`<��`<?�`<��`<�a<�Ca<=na<ŕa<��a<C�a<��a<�a<~�a<��a<K�a<S�a<��a<z�a<��a<�a<
�a<[�a<��a<6�a<��a<�a<��a<k�a<��a<O�a<��a<Q�a<@�a<�a<��a<Xa<�,a<a<]�`<r�`<̮`<�`<K�`<��`<P�`<�`<0'a<yRa<:|a<�a<�a<��a<	�a<��a<��a<��a<�a<u�a<�a<��a<�a<-�a<J�a<��a<ݦa<>�a<L�a<��a<��a<?�a<��a<��a<F�a<��a<��a<�a<�na<FDa<�a<��`<�`<E�`<n�`<��`<۫`<��`<`�`<a<3/a<Za<v�a<�a<��a<��a<_�a<��a<��a<'�a<�a<��a<Ϊa<"�a<��a<;�a<!�a<J�a<ڙa<��a<��a<K�a<�a<��a<��a<��a<}�a<f�a<�a<�qa<�Ha<�a<?�`<��`<M�`<G�`<ņ`<y�`<1�`<+�`<�`<<�`<�a<�Ha<�oa<!�a<D�a< �a<��a<��a<g�a<��a<�a<!�a<D�a<�~a<�wa<�ta<uua<^za<��a<�a<��a<C�a<ͳa<ݻa<C�a<S�a<�a<��a<Bwa<�Qa<(a<��`<��`<4�`<M�`<�~`<�w`<s}`<�`<ߪ`<��`<I�`<�#a<�  �  U?a<�ha<H�a<åa<n�a<��a<��a<��a<B�a<��a<�a<Z�a<��a<�a<��a<X�a<y�a<p�a<�a<��a<��a<8�a<��a<�a<�a<#�a<��a<+ja<�@a<ra<��`<��`<d�`<�|`<�m`<�k`<�v`<��`<��`<%�`< a<u6a<sca<��a<8�a<��a<��a<~�a<��a<T�a<��a<��a<��a<��a<o�a<&�a<�a<��a<X�a<x�a<��a<��a<k�a<*�a<�a<��a<%�a<4�a<Ҥa<�~a<�Sa<g%a<O�`<>�`<@�`<��`<'�`<��`<3�`<:�`<K�`<�a<�0a<�^a<N�a<2�a<B�a<��a<R�a<��a<)�a<��a<Y�a<L�a<�a<l�a<~�a<C�a<L�a<(�a<��a<��a<��a<��a<��a<K�a<D�a<$�a<��a<m�a<ߛa<bsa<�Fa<�a<��`<W�`<x�`<��`<5�`<�`<r�`< �`<}�`<&a<�@a<�ma<��a<ڸa<��a<H�a<�a<��a<X�a<��a<��a<��a<j�a<F�a<�a<��a<R�a<ھa</�a<*�a<�a<c�a<7�a<6�a<��a<��a<:�a<��a<Ήa<t_a<�1a<Ja<^�`<I�`<�`<	�`<ل`<�`<�`<��`<_�`<a<@Ia<�ta<��a<�a<��a<��a<��a<\�a<�a<��a<��a<y�a<=�a<c�a<O�a<B�a<V�a<)�a<��a<6�a<��a<j�a<��a<��a<;�a<��a<��a<�a<�da<18a<�a<��`<Ű`<ލ`<�u`<$i`<�i`<�w`<'�`<��`<U�`<�a</9a<aca<��a<@�a<4�a<9�a< �a<��a<ռa<�a<��a<��a<��a<\�a<��a<a�a<�a<R�a<١a<p�a<7�a<�a<t�a<9�a<�a<V�a<؍a<#la<�Ca<�a<��`<��`<4�`<Yu`<�a`<?Z`<L``<�r`<��`<S�`<C�`<a<�  �  6a< aa<ƅa</�a<��a<A�a<��a<�a<��a<o�a<�a<@�a<�a<D�a< a<}�a<��a<�a<��a<�a<��a<�a<H�a<K�a<�a<'�a<��a<3ba<�6a<�a<%�`<�`<l�`<�j`<�Z`<�X`<�c`<B|`<5�`<v�`<b�`<�+a<�Za<��a<h�a<��a<L�a<��a<��a<m�a<��a<0�a<��a<��a<.�a<��a<��a<��a<�a<I�a<��a<H�a<��a<4�a<��a<��a<y�a<��a<"�a<Pva<Ia<�a<��`<��`<�`<C�`<9w`<�x`<��`< �`<W�`<��`<�$a<�Ta<)�a<��a<�a<��a<`�a<��a<��a<E�a<U�a<��a<b�a<t�a<��a<�a<��a<��a<��a<��a<��a<I�a<-�a<x�a<(�a<��a<a�a<#�a<��a<Kja<k;a<�
a<��`<��`<`<�~`<Hw`<.}`<��`<=�`<+�`<�a<15a<Pda<
�a<W�a<e�a<��a<��a<��a<��a<�a<a�a<f�a<S�a<��a<]�a<R�a<{�a<�a<��a<��a<P�a<V�a<�a<��a<��a<��a<@�a<
�a<؁a<�Ua<�%a<��`<��`<O�`<��`<u`<�q`<\|`<��`<��`<��`<ka<�>a<;la<��a<�a<��a<��a<��a< �a<'�a<��a<w�a<�a<��a<!�a<�a<�a<5�a<׿a<[�a<�a<��a<��a<��a<z�a<��a<S�a<�a<D�a</\a<�-a<��`<a�`<��`<�|`<c`<7V`<W`<se`<�`<��`<`�`<��`<D/a<;[a<��a<�a<�a<E�a<�a<��a<��a<�a<׳a<#�a<��a<i�a<w�a<͟a<n�a<h�a<�a<{�a<�a<��a<��a<�a<��a<��a<��a<�da<p:a<ta<��`<}�`<��`<�c`<�N`<VG`<aM`<�``<�`<�`<�`<�a<�  �  �2a<r^a<�a<�a<��a<��a<Y�a<��a<M�a<	�a<�a<߭a<*�a<��a<&�a<��a<��a<Z�a<��a<F�a<�a<��a<��a<}�a<e�a<ȣa<ąa<T_a<?3a<ha<��`<��`<��`<}d`<�T`<�R`<�]`<`v`<��`<x�`<�`<�'a<�Wa<O�a<ƥa<��a<.�a<-�a<��a<��a<��a<�a<��a<��a<X�a<�a<��a<��a<��a<��a<��a<E�a<��a<x�a<�a<��a<z�a<�a<��a<.sa<9Ea<�a<��`<q�`<�`<�|`<9q`<�r`<��`<Z�`<��`<��`<T a<�Pa<3~a<
�a<��a<��a<��a<=�a<?�a<��a<��a<��a<��a<c�a<��a<b�a< �a<��a<��a< �a<V�a<��a<�a<g�a<w�a<��a<$�a<V�a<��a<�fa<Q7a<sa<k�`<�`<��`<~x`<Xq`<�v`<w�`<��`<��`<a a<1a<�`a<[�a<}�a<�a<h�a<�a<w�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<�a<��a<��a<��a<��a<4�a<�a<:�a<��a<#�a<�~a<)Ra<�!a<��`<7�`<��`<�`<�n`<�k`<�u`<č`<��`<��`<
a<�:a<�ha<i�a<q�a<��a<��a<7�a<J�a<K�a<��a<H�a<F�a<��a<K�a<:�a<D�a<b�a<��a<��a<��a<��a<��a<��a<��a<��a<T�a<��a<�a<Ya<�)a<E�`<{�`<��`<�v`<�\`<8P`<�P`<._`<Hz`<8�`<��`<�`<�+a<EXa<�a<��a<8�a<d�a<��a<�a<��a<V�a<շa<��a<��a<��a<Ԥa<�a<��a<�a<�a<0�a<��a<v�a<��a<m�a<k�a<��a<Ća<Aba<7a<[a<h�`<R�`<�}`<�]`<tH`<hA`<G`<�Z`<'z`<��`<��`<za<�  �  6a< aa<ƅa</�a<��a<A�a<��a<�a<��a<o�a<�a<@�a<�a<D�a< a<}�a<��a<�a<��a<�a<��a<�a<H�a<K�a<�a<'�a<��a<3ba<�6a<�a<%�`<�`<l�`<�j`<�Z`<�X`<�c`<B|`<5�`<v�`<b�`<�+a<�Za<��a<h�a<��a<L�a<��a<��a<m�a<��a<0�a<��a<��a<.�a<��a<��a<��a<�a<I�a<��a<H�a<��a<4�a<��a<��a<y�a<��a<"�a<Pva<Ia<�a<��`<��`<�`<C�`<9w`<�x`<��`< �`<W�`<��`<�$a<�Ta<)�a<��a<�a<��a<`�a<��a<��a<E�a<U�a<��a<b�a<t�a<��a<�a<��a<��a<��a<��a<��a<I�a<-�a<x�a<(�a<��a<a�a<#�a<��a<Kja<k;a<�
a<��`<��`<`<�~`<Hw`<.}`<��`<=�`<+�`<�a<15a<Pda<
�a<W�a<e�a<��a<��a<��a<��a<�a<a�a<f�a<S�a<��a<]�a<R�a<{�a<�a<��a<��a<P�a<V�a<�a<��a<��a<��a<@�a<
�a<؁a<�Ua<�%a<��`<��`<O�`<��`<u`<�q`<\|`<��`<��`<��`<ka<�>a<;la<��a<�a<��a<��a<��a< �a<'�a<��a<w�a<�a<��a<!�a<�a<�a<5�a<׿a<[�a<�a<��a<��a<��a<z�a<��a<S�a<�a<D�a</\a<�-a<��`<a�`<��`<�|`<c`<7V`<W`<se`<�`<��`<`�`<��`<D/a<;[a<��a<�a<�a<E�a<�a<��a<��a<�a<׳a<#�a<��a<i�a<w�a<͟a<n�a<h�a<�a<{�a<�a<��a<��a<�a<��a<��a<��a<�da<p:a<ta<��`<}�`<��`<�c`<�N`<VG`<aM`<�``<�`<�`<�`<�a<�  �  U?a<�ha<H�a<åa<n�a<��a<��a<��a<B�a<��a<�a<Z�a<��a<�a<��a<X�a<y�a<p�a<�a<��a<��a<8�a<��a<�a<�a<#�a<��a<+ja<�@a<ra<��`<��`<d�`<�|`<�m`<�k`<�v`<��`<��`<%�`< a<u6a<sca<��a<8�a<��a<��a<~�a<��a<T�a<��a<��a<��a<��a<o�a<&�a<�a<��a<X�a<x�a<��a<��a<k�a<*�a<�a<��a<%�a<4�a<Ҥa<�~a<�Sa<g%a<O�`<>�`<@�`<��`<'�`<��`<3�`<:�`<K�`<�a<�0a<�^a<N�a<2�a<B�a<��a<R�a<��a<)�a<��a<Y�a<L�a<�a<l�a<~�a<C�a<L�a<(�a<��a<��a<��a<��a<��a<K�a<D�a<$�a<��a<m�a<ߛa<bsa<�Fa<�a<��`<W�`<x�`<��`<5�`<�`<r�`< �`<}�`<&a<�@a<�ma<��a<ڸa<��a<H�a<�a<��a<X�a<��a<��a<��a<j�a<F�a<�a<��a<R�a<ھa</�a<*�a<�a<c�a<7�a<6�a<��a<��a<:�a<��a<Ήa<t_a<�1a<Ja<^�`<I�`<�`<	�`<ل`<�`<�`<��`<_�`<a<@Ia<�ta<��a<�a<��a<��a<��a<\�a<�a<��a<��a<y�a<=�a<c�a<O�a<B�a<V�a<)�a<��a<6�a<��a<j�a<��a<��a<;�a<��a<��a<�a<�da<18a<�a<��`<Ű`<ލ`<�u`<$i`<�i`<�w`<'�`<��`<U�`<�a</9a<aca<��a<@�a<4�a<9�a< �a<��a<ռa<�a<��a<��a<��a<\�a<��a<a�a<�a<R�a<١a<p�a<7�a<�a<t�a<9�a<�a<V�a<؍a<#la<�Ca<�a<��`<��`<4�`<Yu`<�a`<?Z`<L``<�r`<��`<S�`<C�`<a<�  �  �Ma<ta<w�a<��a</�a<�a<f�a<�a<��a<��a<j�a<�a<Y|a<wa<�ua<�xa<�a<��a<<�a<L�a<�a<F�a<o�a<`�a<y�a<ˮa<��a<Lva<�Oa<&a<{�`<��`<3�`</�`<1�`<-�`<s�`<Q�`<�`<��`<%a<9Ga<�pa<��a<M�a<{�a<��a<��a<��a<k�a<�a<c�a<I�a<d�a<��a<�a<Õa<��a<	�a<z�a<:�a<��a<�a<`�a<��a<`�a<��a<��a<��a<�a<�ca<=9a<�a<W�`<��`<��`<˧`<:�`<��`<?�`<��`<�a<�Ca<=na<ŕa<��a<C�a<��a<�a<~�a<��a<K�a<S�a<��a<z�a<��a<�a<
�a<[�a<��a<6�a<��a<�a<��a<k�a<��a<O�a<��a<Q�a<@�a<�a<��a<Xa<�,a<a<]�`<r�`<̮`<�`<K�`<��`<P�`<�`<0'a<yRa<:|a<�a<�a<��a<	�a<��a<��a<��a<�a<u�a<�a<��a<�a<-�a<J�a<��a<ݦa<>�a<L�a<��a<��a<?�a<��a<��a<F�a<��a<��a<�a<�na<FDa<�a<��`<�`<E�`<n�`<��`<۫`<��`<`�`<a<3/a<Za<v�a<�a<��a<��a<_�a<��a<��a<'�a<�a<��a<Ϊa<"�a<��a<;�a<!�a<J�a<ڙa<��a<��a<K�a<�a<��a<��a<��a<}�a<f�a<�a<�qa<�Ha<�a<?�`<��`<M�`<G�`<ņ`<y�`<1�`<+�`<�`<<�`<�a<�Ha<�oa<!�a<D�a< �a<��a<��a<g�a<��a<�a<!�a<D�a<�~a<�wa<�ta<uua<^za<��a<�a<��a<C�a<ͳa<ݻa<C�a<S�a<�a<��a<Bwa<�Qa<(a<��`<��`<4�`<M�`<�~`<�w`<s}`<�`<ߪ`<��`<I�`<�#a<�  �  2`a<�a<�a<(�a<I�a<ٻa<��a<��a<w�a<ۇa<fva<&ga<�[a<�Ta<Sa<�Va<g_a<�la<<}a<��a<ѡa<!�a<��a<$�a<��a<2�a<�a<�a<ca<:=a<�a<��`<��`<�`<0�`<��`<Ҹ`<��`<y�`<�a<34a<!\a<a<<�a<��a<{�a<q�a<��a<j�a<��a</�a<F�a<�a<��a<�va<\ra<sa<�xa<Ճa<��a<��a<[�a<��a<��a<��a<��a<,�a<��a<��a<M�a<mxa<�Qa<d+a<ua<�`<��`<�`<U�`<��`<��`<a<P4a<8[a<Ӂa<�a<g�a<�a<�a<F�a<M�a<��a<��a<�a<K�a<ӗa<Њa<�a<B~a<�a<��a<�a<<�a<�a<��a<��a<�a<��a<8�a<T�a<r�a<K�a<r�a<�ma<�Fa<� a<��`<��`<x�`<d�`<�`<��`<��`<Ja<�Aa<�ha<|�a<دa<��a<a�a<#�a<S�a<��a<e�a<��a<��a<ݠa<)�a<+�a<�}a<�{a<l~a<��a<:�a<C�a<�a<x�a<�a<��a<��a<M�a<@�a<]�a<��a<�a<e[a<P4a<~a<m�`<�`<p�`<��`<=�`<U�`<��`< "a<EHa<�na<D�a<^�a<M�a<��a<�a<�a<��a<>�a<6�a<��a<q�a<?�a<�ta<�na<ima<{qa<�za<��a< �a<��a<��a<�a<r�a<��a< �a<8�a<֡a<$�a<]a<X5a<�a<��`<��`<��`<�`<��`<�`<��`<l�`<a<e6a<t\a<$a<��a< �a<��a<7�a<��a<űa<��a<ݏa<�}a<�la<,_a<�Ua<�Qa<�Ra<\Ya<vda<dsa<Ȅa<y�a<�a<��a<��a<��a<�a<՞a<��a<�ca<�=a<�a<��`<i�`<`�`<Y�`<_�`<?�`<1�`<q�`<�`<�a<:a<�  �  �sa<��a<�a<)�a<4�a<¶a<j�a<��a<j�a<uma<Wa<�Ca<�4a<�+a<�)a<.a<J9a<�Ia<�^a<bva<�a<��a<��a<�a<��a<Q�a<�a<�a<�wa<Wa<�5a<Ea<c�`<��`<��`<+�`<r�`<#�`<�a<.a<;Pa<;sa<ޓa</�a<��a<��a<��a<=�a<9�a<�a<h�a<�a</ma<�[a<fOa<]Ia<�Ia<Qa<�^a<pqa<�a<��a<r�a<��a<\�a<:�a<��a<��a<(�a<�a<��a<Cma<	La<6-a<�a<3a<��`<��`<�a<!a< 4a<�Sa<�ua<:�a<t�a<��a<��a<��a<��a<��a<��a<K�a<t�a<q�a<�ua<ea<�Ya<Ua<�Va<�_a< na<q�a<�a<8�a<K�a<��a<��a<��a<��a<��a<d�a<��a<�a<da<Ca<�%a<la<|�`<�`<F�`<a<2"a<�>a<�_a<z�a<4�a<z�a<�a<c�a<�a<:�a<��a<��a<��a<T�a<��a<�ma<b^a<�Ta<5Ra<�Ua<�`a<�pa<�a<��a<��a<x�a<��a<��a<_�a<Z�a<5�a<}�a<��a<7ua<BSa<�2a<Ka<�a<��`<��`<��`<�a<�$a<HCa<Pda<�a<e�a<U�a<��a<��a<B�a<P�a<��a<��a<r�a<d�a<�na<�[a<[Ma<�Ea<TDa<�Ia<�Ua<fa<={a<��a<k�a<Q�a<&�a<��a<��a<��a<?�a<��a<�sa<�Pa<�.a<�a<�`<��`<��`<��`<�`<
�`<Oa<�/a<�Pa<�qa<��a<Q�a<̷a<3�a<��a<6�a<ǣa<��a<Nwa<�_a<uJa<l9a<�-a<�(a<
*a<R2a<�@a<�Sa<�ia<ۀa<��a<��a<�a<M�a<Q�a<$�a<��a<�va<Va<�3a<�a<O�`<4�`<S�`<��`<\�`<L�`<��`<�a<�0a<�Ra<�  �  ��a<��a<��a<��a<s�a<��a<��a<��a<~la<�Oa<Q4a<�a<o
a<]�`<b�`<�a<xa<�#a<7=a<�Ya<Rwa<�a<�a<,�a<�a<Ϳa<�a<J�a<݌a<�qa<aUa<�:a<J$a<�a<E
a<$	a<na<�a<,5a<�Oa<&ma<��a<��a<��a<��a<}�a<�a<'�a<��a<ҙa<�~a<�ba<�Ha<s3a<&$a<Ma<�a<�%a<	6a<�La<�ga<p�a<��a<ؼa<��a<$�a<�a<��a<�a<�a<�a<��a<?ma<ISa<>a</a<�'a<�(a<�1a<vBa<Ya<�sa<Ȑa<۬a<k�a<i�a<��a<��a<b�a<��a<k�a<C�a<��a<>ia<�Oa<~;a<�-a<�'a<*a<�4a<�Fa< ^a<�ya<��a<c�a<<�a<+�a<?�a<��a<��a<�a<��a<�a<�a<�ea<Ma<�9a<�,a<(a<�+a<�7a<;Ja<^ba<~a<�a<��a<��a<D�a<��a<M�a<�a<��a<T�a<a<�za<�^a<�Fa<�3a<O(a<�$a<�)a<�6a<MJa<(ca</a<�a<]�a<E�a<��a<��a<��a<:�a<��a<��a<ԏa<�ra<�Wa<4@a<�.a<�$a<�"a<�(a<7a<�Ka<ea<A�a<��a<.�a<��a<|�a<��a<��a<<�a<)�a<��a<��a<�ea<aJa<43a<"a<va<(a<)a<�,a<�Aa<.[a<wa<��a<1�a<m�a<h�a<��a<?�a<$�a<�a<�a<&ma<�Oa<�4a<�a<�a<�a<�a<ha<]a<d5a<�Oa<�ka<�a<��a<��a<�a<-�a<`�a<A�a<Y�a<�xa<v[a<�>a<�$a<�a<�a<:�`<K�`<�a<
a<R0a<~Ka<Dha<ȃa<e�a<�a<��a<$�a<G�a<>�a<ĉa<�na<�Qa<�5a<�a<Y	a<��`<��`<��`<�a<�a<3a<Oa<9la<�  �  ��a<6�a<��a<��a<Ӵa<}�a<$�a<�sa<�Ra<	1a<�a<[�`<��`<��`<b�`<��`<|�`<h�`<�a<8<a<�^a<�a<ƛa<[�a<u�a<h�a<�a<�a<�a<��a<�sa<f^a<La<�>a<7a<p6a<M<a<�Ha<�Za<�pa<��a<i�a<��a<O�a<��a<9�a<��a<+�a<r�a<݃a<ca<@Ba<�#a<�	a<��`<k�`<��`<��`<a<�&a<�Fa<\ia<&�a<��a<�a<-�a<?�a<@�a<�a<��a<�a<��a<��a<^xa<ga<�Za<�Ta<�Ua<]a<�ja<-}a<�a<W�a<��a<��a<*�a<��a<��a<-�a<�a<K�a<h�a<[ha<(Ga<�(a<�a<~ a<��`<_�`<�a<�a<�9a<IZa<M|a<��a<�a<v�a<�a<��a<4�a<��a<&�a<�a<Ԟa<�a<�sa<�ca</Ya<�Ua<PXa<�aa<&qa<�a<��a<��a<��a<3�a<-�a<7�a<��a<��a<4�a<E�a<~a<�[a<�:a<Da<;a<��`<��`<v�`<�a<�"a<�@a<paa<f�a<��a<�a<��a<(�a<e�a<Y�a<x�a<�a<��a<h�a<{a<�ga<�Ya<dQa<�Oa<�Ta<p`a<qa<��a<Ϝa<I�a<O�a<~�a<��a<x�a<l�a<D�a<�a<��a<ha<�Ea<%a<�	a<��`<��`<8�`<y�`<�a<�a<C:a<�Za<|a<R�a<ղa<m�a<
�a<��a<-�a<Y�a<��a<�a<pa<�Ya<�Ga<Z:a<�3a<�3a<�:a<�Ga<zYa<�na<��a<O�a<��a<úa<�a<+�a<2�a<�a<A�a<�`a<F>a<�a<��`<E�`<��`<<�`<��`<��`<]�`<a<7,a<�Ma<oa<I�a<f�a<Ȳa<�a<��a<�a<&�a<ʅa<�na<�Wa<FCa<U3a<�(a<b%a<P(a<2a<�Aa<�Ua<~la<Ӄa<�  �  �a<2�a<`�a<ùa<��a<e�a<:�a<�_a<�9a<�a<��`<��`<��`<��`<Ţ`<ȩ`<̻`<��`<��`<Ma<�Fa<�la<��a<N�a<T�a<b�a<��a<)�a<��a<�a<C�a<f~a<!pa<�ea<�_a<�_a<rda<�na<�|a<9�a<�a<r�a<r�a<��a<�a<M�a<��a<��a<��a<,na<fHa<q"a<l�`<��`<��`<��`<O�`<��`<f�`<Ka<�&a<8Na<�ua<��a<�a<��a<��a<��a<��a<��a<p�a<@�a<��a<ߙa<H�a<��a<~a<�~a<v�a<!�a<��a<��a<��a<��a<z�a<��a<��a<	�a<��a<��a<�a<sa<�Ka<�%a<�a<_�`<��`<��`<�`<9�`<�`<�a<�;a<�ba<#�a<��a<��a<=�a<��a<��a<Y�a<	�a<�a<[�a<��a<{�a<��a<��a<�~a<��a<��a<q�a<�a<��a<L�a<n�a<4�a<�a<�a<f�a<��a<H�a<E�a<ea<�=a<&a<��`<��`<|�`<�`<��`<��`<5�`<�a<|Da<rka<��a<�a<��a< �a<Z�a<=�a<��a<��a<��a<��a<�a<�a<܀a<Gza<ya<�|a<�a<�a<��a<�a<V�a<�a<��a<��a<��a<}�a<��a<0�a<�ta<tMa<�%a<� a<R�`<��`<�`<��`<&�`<4�`<W�`<�a<�?a<�ea<�a<��a<�a<��a<Y�a<��a<s�a<�a<��a<�a<O{a<�la<Kba<�\a<�\a<�aa<la<�ya<��a<�a<��a<��a<5�a<��a<��a<��a<B�a<�na<yIa<�!a</�`<��`<�`<ϩ`<��`<Q�`<�`<��`<��`<�a<f4a<�Za<�|a<˘a<�a<:�a<Һa<z�a<�a<�a<�a<7va< fa<�Ya<lQa<�Na<�Pa<�Xa<�da<�ta<��a<��a<�  �  ��a<��a<T�a<n�a<٩a<��a<2sa<(Ma<Y#a<0�`<t�`</�`<,�`<ŀ`<Z|`<8�`<ؗ`<��`<)�`<�a<`1a<W[a<��a<W�a<��a<��a<��a<��a<Ƚa<��a<��a<#�a<��a<�a<��a<c�a<�a<+�a<�a<�a<�a<��a<��a<h�a<��a<~�a<��a<��a<0�a<ZZa<�0a<ma<��`<��`<��`<М`<�`<j�`<;�`<c�`<.
a<�5a<�aa<��a<s�a<%�a<��a<��a<�a<��a<8�a<��a<x�a<�a<��a<��a<ʠa<M�a<�a<߭a<Ӹa<��a<e�a<��a<e�a<��a<��a<��a<�a<7�a<Ԇa<�]a<�2a<�a<��`<��`<G�`<��`<�`<��`<��`<��`<l a<�Ka<2va<�a<��a<�a<��a<�a<P�a<u�a<��a<]�a<ҿa<��a<E�a<�a<��a<{�a<�a<�a<нa<�a<S�a<a�a<��a<��a<��a<��a<	�a<>�a<�xa<�Na<�"a<��`<	�`<��`<��`<��`<�`<�`<(�`<� a<�*a<�Ua<a<�a<��a<9�a<��a<)�a<*�a<��a<��a<�a<Եa<p�a<�a<�a<Лa<��a<��a<��a<ֻa<�a<��a<h�a<��a<G�a<��a<f�a<��a<��a<"aa<�5a<�	a<v�`<x�`<��`<��`<l�`<��`<�`<o�`<~�`<�'a<�Qa<�xa<4�a<`�a<J�a<Y�a<&�a<R�a<��a<>�a<ޤa<Q�a<+�a<0�a<�a<za<q�a<��a<�a<��a<��a<3�a<��a<��a<��a<Z�a<�a<��a<�]a<W4a<�a<��`<�`<(�`<^�`<8{`<_~`<�`<��`<�`<a�`<�a<�Ga<@na<��a<Ȧa<k�a<L�a<l�a<h�a<k�a<�a<v�a<K�a<�ya<�sa<fqa<isa<>ya<f�a<p�a<�a<��a<�  �  ��a<��a<��a<��a<��a<5�a<�ga<[>a<Na<�`<��`<ő`<�t`<�c`<�^`<@g`<�{`<ԛ`< �`<��`< a<CMa<va<��a<1�a<��a<�a<c�a<�a<��a<Y�a<E�a<K�a<�a<��a<��a<؟a<ԥa<��a<��a<��a<��a<7�a<X�a<��a<��a<~�a<�a<�ta<~Ja<Ka<c�`<D�`<��`<"�`<H`<s`<ٌ`<�`<s�`<��`<B"a<lQa<�}a<z�a<��a<7�a<��a<��a<��a<��a<=�a<S�a<�a<�a<��a<�a<^�a<��a<��a<Q�a<��a<�a<<�a<��a<��a<��a<��a<��a<��a<ya<�La<Xa<��`<Z�`<�`<l�`<؉`<��`<D�`<>�`<��`<�
a<_9a<ga<#�a<�a<��a<��a<��a<�a<��a<��a<��a<��a<��a<Z�a<��a<׻a<D�a<f�a<b�a<@�a<�a<��a<��a<��a<N�a<��a<��a<��a<��a<�ia<�<a<�a<�`<��`<T�`<^�`<�`<�`<�`<F�`<��`<	a<�Da<qa<�a<�a<��a<��a<T�a<��a<��a<��a<��a<��a<;�a<��a<�a<�a<Z�a<X�a<�a<�a<��a<��a<��a<��a<a�a<��a<8�a<�a<}a<HQa<]"a<��`<��`<\�`<�`<r{`<�y`<m�`<��`<~�`</�`<�a<^Aa<�ka<8�a<Үa<��a<�a<��a<R�a<Y�a<��a<��a<w�a<��a<W�a<ՙa<��a<;�a<��a<��a<��a<3�a<��a<��a<C�a<��a<Q�a<ۘa<xa<%Pa<f#a<Z�`< �`<`�`<s}`<�g`<�]`<a`<3q`<Ռ`<�`<��`<a<y8a<Mba<ͅa<M�a<"�a<0�a< �a<��a<L�a<��a<��a<Z�a<�a<e�a<��a<+�a<~�a<��a<ۡa<��a<�a<�  �  ��a<u�a<7�a<�a<�a<��a<�_a<�4a<�a<��`<M�`<��`<c`<�P`<�K`<hT`<Xj`<?�`<��`<��`<a<FDa<�na<��a<�a<��a<�a<��a<��a<��a<��a<y�a<z�a<�a<�a<N�a<ٯa<Ĵa<��a<��a<��a<f�a<��a<F�a<��a<;�a<0�a<��a<Ola<v@a<,a<O�`<:�`<o�`<�y`<Ol`<�l`<Pz`<��`<D�`<��`<�a<)Ga<Dua<�a<�a<��a<q�a<]�a<��a<4�a<��a<C�a<�a<��a<��a<��a<��a<i�a<C�a<��a<]�a<�a<:�a<-�a<��a<��a<��a<׻a<��a<Mpa<Ba<�a<��`<ڸ`<a�`<��`<�v`<�z`<*�`<S�`<�`<T�`<�-a<w]a<D�a<
�a<��a<��a<D�a<��a<��a<��a<R�a<��a<`�a<��a<��a<��a<��a<��a<2�a<�a<��a<��a<1�a<~�a<��a<1�a<��a<	�a<��a<�`a<�0a<i a<��`<ɪ`<`�`<jy`<�s`<|`<h�`<��`<��`<	a<x9a< ha<ϑa<�a<��a<��a<R�a<@�a<��a<��a<��a<+�a<j�a<:�a<_�a<��a<\�a<J�a<*�a<D�a<��a<S�a<F�a<��a<S�a<��a<�a<��a<�ta<AGa<>a<��`<ȸ`<3�`<�w`<zh`<�f`<�r`<m�`<N�`<��`<�a<7a<�ca<��a<P�a<o�a<��a<a�a<��a<��a<9�a<��a<h�a<]�a<E�a<��a<�a<�a<"�a<�a<�a<3�a<��a<T�a<~�a<�a<J�a<�a<qa<YGa<�a<��`<U�`<�`<�k`<�T`<�J`<N`<_`<�{`<b�`<M�`<N�`<�.a<nZa<�a<k�a<R�a<��a<��a<��a<Z�a<��a<�a<�a<)�a<��a<h�a<u�a<ՠa<��a<��a<��a<5�a<�  �  �a<~�a<��a<�a<�a<�ya<{]a<�<a<�a<<�`<Z�`<;�`<��`<r�`<�`<O�`<ƥ`<]�`<��`<� a<�%a<�Ia<Uja<=�a<Λa<%�a<�a<׷a<Y�a<��a<�a<��a<��a<b�a<��a<�a<E�a<��a<Q�a<��a<�a<��a<�a<��a<�a<Ҳa<��a<�a<�la<FKa<�'a<9a<-�`<��`<ַ`<F�`<��`<ڸ`<��`<�`<g	a<�-a<�Ra<va<��a<��a<��a<0�a<�a</�a<O�a<��a<G�a<��a<��a<�a<_�a<��a<��a<�a<:�a<Z�a<	�a<I�a<��a<!�a<t�a<^�a<'�a<z�a<�sa<�Pa<v,a<�	a<7�`<Z�`<Y�`<q�`<5�`<�`<��`<��`<�a<uAa<�ea<'�a<d�a<��a<k�a<��a<��a<��a<��a<��a<Z�a<��a<	�a<׿a<��a<t�a<K�a<��a<�a<$�a<S�a<��a<��a<q�a<�a<B�a<��a<؈a<�ga<yCa<Pa<��`<_�`<��`<��`<��`<P�`</�`<(�`<�a<X%a<XIa<�la<ʌa< �a<޼a<��a<��a<��a<��a<�a<��a<��a<8�a<лa<4�a<��a<�a<X�a<�a<��a<Q�a<��a<��a<Z�a<�a<��a<جa<��a<�ta<�Qa<�,a<Ta<��`<��`<͵`<��`<#�`<��`<��`<t�`<!�`<�a<:Ca<ea<�a<}�a<n�a<Y�a<��a<Ͽa<üa<K�a<��a<֩a<�a<��a<%�a<��a<P�a<ơa<L�a<իa<�a<��a<��a<l�a<8�a<��a<��a<�ka<�Ka<�'a<$a<��`<�`<��`<.�`<ݍ`<=�`<��`<6�`<��`<>�`<�a<�7a<Ya<va<�a<��a< �a<��a<��a<Z�a<�a<ӝa</�a<��a<_�a<4�a<9�a<>�a<�a<��a<٣a<W�a<�  �  ��a<۬a<X�a<S�a<Ґa< {a<V_a<1?a<a<��`<)�`<[�`<z�`<"�`<��`<�`<8�`<~�`<Q�`<+a<�(a<�Ka<�ka<>�a<t�a<P�a<Գa<�a<˵a<ʱa<C�a<q�a<J�a<z�a<��a<ʛa<W�a<Ţa<�a<	�a<i�a<��a<��a<Z�a<ӽa<e�a<{�a<?�a<�na<�Ma<'+a<�a<(�`<�`<k�`<ٲ`<-�`<|�`<�`< �`<�a<�0a<�Ua<?xa<�a<n�a<��a<$�a<��a<�a<x�a<��a<W�a<<�a<�a<-�a<D�a<��a<	�a<^�a<�a<��a<��a<��a<��a<��a<��a<�a<�a<�a<va<�Sa<�/a<'a<O�`<��`<�`<��`<��`<��`<��`<}�`<� a<�Da<=ha<�a<��a<b�a<��a<��a<!�a<��a<��a<��a<]�a<;�a<#�a<�a<y�a<z�a<h�a<0�a<�a<��a<G�a<J�a<'�a<F�a<��a<��a<Ŧa<��a<$ja<�Fa<�"a<� a<��`< �`<B�`<!�`<�`<��`<K�`<za<�(a<eLa<oa<o�a<�a<��a<��a<}�a< �a<	�a<O�a<�a<x�a<��a<�a<-�a<y�a<�a<��a<��a<��a<��a<��a<��a<��a<��a<�a<��a<�a<�va<nTa<�/a<�a<��`<��`<a�`<�`<��`<F�`<�`<��`<� a<#a<
Fa<-ga<\�a<^�a<�a<M�a<��a<��a<�a<�a<��a<��a<X�a<��a<
�a<��a<`�a<�a<+�a<�a<��a<�a<��a<�a<N�a<A�a<ևa<Dma<�Ma<�*a<ja<X�`<�`<��`<�`<`�`<�`<:�`<R�`<~�`<��`<a<e:a<�Za<Awa<Սa<#�a<�a<�a<X�a<[�a<{�a<ؚa<��a<��a<k�a<�a<@�a<\�a<\�a<��a<:�a<L�a<�  �  R�a</�a<K�a<	�a<1�a< a<�da<Fa<�$a<ua<t�`<��`<��`<�`<Y�`<ʧ`<%�`<��`<?�`<�a<�0a<�Ra<Cqa<�a<��a<��a<|�a<��a<%�a<��a<D�a< �a<h�a<Ǒa<��a<��a<i�a<��a<�a<h�a<q�a<f�a<�a<F�a<U�a<��a<U�a<͏a<�ta<kUa<4a<
a<��`<��`<��`<��`<�`<�`<��`<��`<ma<	:a<%]a<l~a<��a<q�a<�a<��a<��a<u�a<Y�a<��a<��a<Z�a<��a<F�a<�a<{�a<=�a<T�a<�a<X�a<Y�a<��a<��a<X�a<��a<��a<��a<5�a<�|a<�[a<'9a<�a<\�`<��`<��`<��`<��`<��`<k�`<�
a<�*a<SMa<Poa<َa<ɩa<�a<��a<��a<��a<q�a<�a<��a<g�a<ݹa<��a<ݯa<?�a<n�a<زa<��a<�a<��a<f�a<��a<y�a<8�a<��a<[�a<Ūa<N�a<
qa<&Oa<�,a<a<��`<N�`<�`<��`<��`<��`<q�`<ka<;2a<�Ta<�ua<��a<��a<��a<�a<'�a<��a<d�a<�a<�a<�a<��a<5�a<�a<A�a<'�a<?�a<��a<��a<��a<��a< �a<��a<}�a<n�a<��a<t�a<�|a<�[a<�8a<$a<A�`<X�`<��`<�`<��`<��`<��`<V�`<'a<!,a<�Ma<Zma<�a<b�a<��a<	�a<��a<�a<εa<�a<+�a<��a<$�a<ُa<ٌa<��a<��a<�a<��a<Ӡa<B�a</�a<t�a<��a<p�a<*�a<F�a<fra<=Ta<�2a<�a<�`<�`<ѷ`<��`<-�`<��`<��`<��`<��`<��`<�a<xAa<�`a<u{a<c�a<�a<�a<��a<2�a<��a<�a<�a<U�a<%�a<i�a<�~a<7�a<σa<щa<b�a<��a<m�a<�  �  P�a<Υa<��a<ޡa<��a<ׄa<.ma<�Pa<�1a<a<�`<�`<L�`<V�`<=�`<�`<��`<��`<t�`<�a<e=a<�\a<�xa<*�a<I�a<��a<C�a<��a<�a<�a<S�a<��a<Q�a</a<�{a<�{a<Ba<��a<��a<Y�a<��a<}�a<��a<μa<��a<X�a<��a<}�a<�}a<aa<1Ba<R#a<a<��`<��`<S�`<��`<%�`<��`<`
a<�'a<dHa<ia<Ƈa<��a<�a<��a<m�a<��a<��a<��a<U�a<�a<L�a<�a<A�a<y�a<ݙa<��a<�a<�a<'�a<��a<��a<[�a<��a<��a<h�a<��a<��a<��a<�ga<Ha<�(a<;a<��`<�`<��`<3�`<��`<a<�a<�:a<�Za<nza<W�a<�a<��a<��a<��a<��a<��a<r�a<O�a<ϲa<>�a<��a<w�a<��a<��a<��a<ԧa<�a<i�a<��a<��a<�a<��a<j�a<��a<��a<��a<�{a<b\a<*<a<�a<=a<��`<�`<��`<�`<�`<�a<�"a<fAa<Baa<�a<z�a<��a<_�a<Y�a<��a<��a<��a<��a<�a<��a<��a<��a<|�a<��a<��a<u�a<^�a<�a<(�a<��a<��a<Z�a<��a<	�a<��a<!�a<օa<�ga<�Fa<k&a<{a<A�`<��`<��`<A�`<��`<��`<��`<�a<}:a<�Ya<�va<�a<ڣa<z�a<��a<��a<<�a<0�a<��a<e�a<��a<��a<�|a<Bya<�xa<�{a<ȁa<��a<��a<x�a<3�a<,�a<�a<��a<��a<H�a<�ya<6^a<&?a<�a<�`<��`<$�`<Ѽ`<�`<5�`<J�`<O�`<��`<va<=-a<�La<?ia<��a<	�a<�a<��a<u�a<{�a<�a<��a<Q�a<�ya<ra<ma<Qka<�la<�qa<ya<��a<%�a<��a<�  �  ��a<t�a<�a<R�a<k�a<�a<�wa<�^a<�Ba<�%a<�
a<��`<�`<�`<I�`<��`<�`<�`<\a<�/a<iMa<�ia<��a<��a<b�a<��a<��a<�a<�a<��a<'�a<Qya<{na<�fa<ba<ba<�ea<�ma<ya<ʆa<=�a<\�a<h�a<��a<Һa<�a<��a<��a<H�a<�oa<�Sa<8a<ja<<	a<�`<D�`<��`<]�`<�a<�!a<=a<jZa<xa<��a<(�a<Q�a<��a<��a<��a<e�a<��a<&�a<ءa<�a<��a<�a<�a<�a<��a<�a<7�a<��a<�a<�a<��a<��a<�a< �a<��a<�a<$�a<�wa<�Za<�>a<c%a<>a<ya<��`<��`<�
a<2a<�3a<�Na<�ka<w�a<�a<\�a<��a<��a<,�a<��a<X�a<~�a<*�a<��a<�a<c�a<�a<��a<E�a<7�a<p�a<u�a<�a<0�a<+�a<��a<��a<��a<��a<��a<�a<��a<ma<�Oa<-4a<0a<�	a<7�`<��`<��`<�a<�a<�8a<~Ta<Mqa<��a<�a<k�a<|�a<�a<N�a<��a<5�a<|�a<�a<W�a<��a<�a<�{a<�za<�}a<��a<��a<[�a<��a<��a<I�a< �a<��a<��a<��a<L�a<U�a</va<�Xa<5;a<�a<�a<��`<��`<@�`<'�`<�a<ca<�0a<�La<�ha<��a<��a<F�a<j�a<$�a<��a<�a<v�a<��a<-�a<Kwa<la<�ca<`_a<_a<ca<�ja<Jua<�a<�a<L�a<��a<�a<کa<V�a<g�a<�a<�ja<�Na<l1a<�a<�`<u�`<A�`<�`<��`<6�`<}�`<~a<�!a<F>a<�Za<ta<
�a<D�a<�a<C�a<��a<"�a<*�a<�}a<
pa<�ca<�Ya<{Sa<nQa<Sa<:Ya<�ba<�na<�|a<>�a<�  �  O�a<D�a<��a<�a<�a<L�a<ɂa<�ma<UUa<D<a<?$a<Za<��`<��`<��`<\�`<a<�a<v,a<�Ea<g_a<�wa<��a<�a< �a<��a<��a<Ξa<�a<�a<4qa<'aa<kSa<]Ia<�Ca<iCa<Ha<�Qa<�_a<[pa<w�a<��a<p�a<Ӱa<�a<�a<J�a<J�a<̕a<�a<�ga<�Oa<9a<V&a<)a<la<�a<�a<�(a<�<a<Ua<�na<��a<��a<9�a<s�a<H�a<��a<t�a<ݻa<��a<לa<a<�{a<�na<\ea<�`a<�aa<Qga<�qa<�a<D�a<��a<o�a<V�a<M�a<��a<W�a<��a<�a<�a<S�a<pa<eWa<�@a</a<#a<�a< a<P)a<�8a<�Ma<�ea<a<��a<ƭa<#�a<��a<��a<X�a<��a<z�a<Ϊa<v�a<L�a<�xa<�la<�da<�aa<da<qka<�va<�a<іa<�a<�a<��a<��a<��a<�a<�a<,�a<{�a<�a<ffa<�Ma<�8a<C(a</a<.a<va<�*a<�;a<�Qa<&ja<R�a<�a<��a<ܾa< �a<��a<F�a<ʽa<&�a<��a<��a<-}a<�na<�ca<X]a<\a<�_a<�ha<9ua<�a<ٕa<��a<N�a<Y�a<�a<��a<v�a<�a<םa<_�a<�la<�Ra<p:a<&a<a<�a<ra<sa< a<I2a<�Ha<�`a<?ya<~�a<��a<j�a<մa<��a<Y�a<��a<�a<9�a<oa<&^a<%Pa<�Ea<�@a<�@a<�Ea<\Oa<�\a<�la<�}a<ȍa<#�a<��a<J�a<��a<c�a<�a<�xa<m`a<�Fa<�-a<�a<>a<��`<P�`<��`<��`<a<� a<j8a<}Qa<�ia<�a<ѐa<+�a<�a<s�a<˗a<J�a<�{a<ja<�Xa<qIa<`=a<t5a<�2a<�4a<z<a<6Ha<fWa<�ha<'za<�  �  H|a<��a<�a<��a<��a< �a<Ǎa<�|a<�ha<^Sa<?a<R-a<�a<�a<ta<�a<�#a<43a<xFa<�[a<�qa<
�a<�a<�a<Ĩa<�a<�a<*�a<ނa<�na<Za<Fa<�5a<l)a<�"a<�!a<�'a<3a<vCa<�Wa<�ma<ăa<֗a<��a<��a<ĸa<S�a<��a<�a<��a<�|a<	ha<Ua<(Ea<�9a<94a<�4a<�;a<Ha<AYa<�ma<��a<ʙa<D�a<��a<��a<��a<��a<��a<��a<9�a<d�a<\sa<`a<Pa<�Da<w?a<;@a<6Ga<�Sa<�da<�xa<=�a<��a<7�a<N�a<��a<��a<+�a<��a<��a<W�a<��a<qa<�]a<�Na<mDa<�?a<�Aa<�Ia<Wa<�ha<A}a<�a<e�a<1�a<n�a<��a<��a<*�a<��a<�a<#�a<��a<�na<\a<nMa<Da<Z@a<*Ca<�Ka<�Ya<�ka<��a<��a<ީa<ܺa<��a<�a<��a<��a<+�a<��a<O�a<�}a<�ha<�Va<�Ha<�?a<(=a<�@a<gJa<!Ya<�ka<z�a<ӕa<L�a<��a<��a<��a<��a<��a<)�a<#�a<��a<�va<�ba<�Pa<�Ca<$<a<�:a<N?a<�Ia<Ya<la<�a<�a<��a<�a<��a<n�a<}�a<+�a<�a<��a<d�a<ka<sVa<�Da<�7a<t0a<H/a<l4a<"?a<�Na<�aa<va<M�a<8�a<e�a<�a<,�a<�a<z�a<g�a<��a<�la<�Va<hBa<�1a<�%a<Ha<La<�%a<[1a<�Aa<,Ua<$ja<M~a<�a<��a<a�a<ڦa<Сa<��a<8�a<kra<�\a<Ga<�3a<�#a<'a<?a<�a<Sa<X*a<�;a<�Oa<Qea<�ya<�a<�a<K�a<	�a<I�a<��a<�}a<�ia<;Ta<\?a<�,a<a<�a<a<a<�a<&+a<�=a<MRa<ha<�  �  ]ma<Ղa<q�a<�a<G�a<�a<��a<�a<{a<�ia<+Ya<�Ja<q?a<�8a<�6a<:a<Ca<�Oa<�_a<vqa<L�a<]�a<�a<ݧa<��a<��a<�a<��a<�ra<�Za<YBa<+a<Ta<�a<� a< a<ga<�a<�&a<2>a<�Wa<ra<`�a<�a<�a<��a<s�a<Ƕa<r�a<B�a<X�a<�a<Cpa<Nca<Za<�Ua<;Va<�[a<|fa<�ta<�a<$�a<�a<"�a<��a<~�a<�a<��a<��a<��a<�a<sa<_Za<yCa<�0a<�#a<�a<ma<�&a<�4a<�Ha<�`a<�ya<��a<.�a<N�a<��a<�a<��a<*�a<}�a<X�a<+�a<�a<Aza<�ma<	ea<taa<�ba<�ia<�ta<U�a<5�a<��a<,�a<��a<��a<��a<��a<�a<B�a<s�a<f�a<ma<�Ta<�>a<y-a<�"a<]a<�!a<�+a<<a<UQa<�ia<Ăa<�a<�a<T�a<��a<p�a<��a<�a<�a<��a<�a<�a<�sa<:ha<�`a<�^a<�aa<�ia<�ua<�a<�a<G�a<��a<��a<��a<��a<3�a<:�a<��a<A�a<{xa<#_a<Ga<�2a<S#a<[a<�a<a<?*a<;<a<�Ra<9ka<&�a<7�a<��a<��a<T�a<��a<c�a<y�a<��a<�a<�a<�qa<�ba<Xa<�Qa<�Pa<�Ta<�]a<9ja<�ya<A�a<n�a<�a<�a<z�a<��a<1�a<{�a<p�a<rqa<~Wa<�=a<�%a<Sa<�a<k�`<��`<�a<�a<�%a<=a<�Ua<�ma<��a<��a<��a<8�a<K�a<B�a<�a<f�a<�qa<`a<�Oa<�Ba<�9a<�5a<�6a<0=a<�Ga<CVa<�fa<xa<O�a<~�a<h�a<}�a<�a<(�a<?�a<Noa<%Wa<�=a<$%a<+a<�`</�`<&�`<t�`<��`<Qa<�"a<e;a<�Ta<�  �  �^a<�wa<R�a<֚a<̢a<i�a<�a<a�a<Z�a<2~a<�pa<#ea<J\a<�Va<�Ua<zXa<�_a<�ia<�va<�a<��a<��a<��a<q�a<3�a<��a<��a<�|a<|ca<�Ga<V+a<�a<��`<�`<��`<��`<��`<��`<@a<�%a<�Ba<�`a<�|a<N�a<��a<��a<:�a<u�a<A�a<�a<��a<[�a<�a<�~a<�wa<ta<�ta<�ya<:�a<ʍa<֛a<6�a<�a<h�a<��a<��a<d�a<��a<B�a<��a<�za<i^a<,Ba<j(a<ha<�a<]�`<I�`<ya<�a<^.a</Ia<�ea<��a<��a<�a<`�a<D�a<��a<.�a<��a<j�a<4�a<��a<�a<�a<�a<8�a<?�a<��a<��a<Z�a<��a<w�a<�a<n�a<��a<��a<��a<[�a<��a<#�a</ta<9Wa<9;a<�"a<Za<�a<�`<�a<Ra<�a<�7a<[Sa<(pa<<�a<��a<4�a<]�a<��a<3�a<��a<e�a<��a<c�a<��a<n�a<�a<a<�}a<�a<#�a<��a<!�a<��a<¶a<M�a<,�a<X�a<b�a<�a<@�a<��a<Ła<ea< Ha<�,a<�a<|a<F�`<c�`<��`<�a<� a<":a<&Va<�ra<��a<ʤa<Ѷa<R�a<_�a<�a<F�a<g�a<��a<o�a<L�a<y~a<~ua<Npa<Ooa<Rra<Rya<3�a<��a<U�a<��a<`�a<+�a<��a<��a<ئa<0�a<I|a<�`a<�Ba<�%a<�
a<��`<*�`<4�`<_�`<��`<��`<ta<�%a<�Aa<�]a<�wa< �a<�a<h�a<i�a<A�a<>�a<q�a<��a<�va<|ia<_a<�Wa<}Ta<$Ua<:Za<�ba<Dna<�{a<׈a<(�a<V�a<C�a<o�a<7�a<��a<�ya<aa<�Da<�'a<�a<?�`<�`<_�`<��`<��`<r�`<�`<O	a<2%a<JBa<�  �  /Qa<�ma<a�a<+�a<��a<r�a<��a<Y�a<ߘa<ώa<��a<�{a<�ta<pa<�oa<�qa<�wa<�a<�a<�a<y�a<"�a<S�a<ŭa<7�a<6�a<܉a<�qa<IUa<P6a<a<��`<D�`<�`<��`<��`<w�`<��`<?�`<a<G0a<Qa<rpa<I�a<Ǣa<,�a<�a<��a<�a<�a<��a<�a<ŝa<��a<{�a<�a<��a<��a<��a<��a<�a<2�a<��a<j�a<]�a<��a<A�a< �a<��a<��a<�ka<5La<�,a<�a<_�`<=�`<X�`<c�`<d�`<l�`<1a<�4a<bTa<#ta<��a<�a<��a<��a<��a<��a<w�a<��a<�a<i�a<��a<ơa<X�a< �a<	�a<I�a<U�a<��a<��a<a�a<e�a<\�a<�a<�a<��a<��a<ўa<��a<�ca<�Ca<(%a<
a<��`<
�`<
�`<��`<��`<�a<k!a<�?a<�_a<�~a<՚a<A�a<��a<��a<>�a<�a<`�a<�a<�a<o�a<�a<��a<Ҙa<p�a</�a<3�a<ѥa<B�a<��a<��a<x�a<��a<��a<k�a<��a<��a<��a<�sa<�Sa<�3a<�a<|�`<��`<{�`<X�`<!�`<V�`<�a<�$a<�Ca<8ca<C�a<Ûa<۰a<οa<7�a<Q�a<��a<}�a<Y�a<"�a<%�a<��a<o�a<,�a<1�a<n�a<��a<a�a<��a<Q�a< �a<c�a<Ӽa<�a<װa<<�a<��a<Cpa<UQa<�0a<Ta<�`<��`<��`<0�`<{�`<��`<%�`<H�`<a<H0a<wOa<Ula<!�a<;�a<�a<g�a<��a<��a<Şa<b�a<j�a<Ba<�va<�pa<`na<�na<�ra<�ya<k�a<��a<��a<��a<D�a<��a<��a<�a<�a<�oa<�Sa<�4a<�a<��`<��`<r�`<ȷ`<�`<�`<��`<O�`<�`<�a<�1a<�  �  tFa<�ea<�a<�a<ϡa<)�a<+�a<��a<�a<b�a<��a<�a<�a<��a<8�a<I�a<��a<M�a<T�a<�a<�a<��a<@�a<�a<�a<l�a<��a<ia<	Ja<�(a<a<�`<��`<S�`<n�`<�`<O�`<h�`<~�`<;�`<�!a<�Da<�fa<�a<�a<۰a<#�a<j�a<S�a<=�a<��a<e�a<{�a<M�a<C�a<��a<E�a<��a<%�a<�a<��a<u�a<�a<�a<X�a<?�a<;�a<f�a<}�a<�a<�_a<�=a<Ha<�`<=�`<&�`<��`<��`<��`<��`<a<`$a<uFa<�ha<��a<b�a<��a<y�a<��a<>�a<��a<��a<��a<��a<�a<��a<��a<��a<��a<ӱa<[�a<��a<��a<��a<��a<4�a<�a<��a<��a<K�a<�a<�xa<&Wa<�4a<�a<��`<?�`<��`<�`<��`<��`<��`<�a<40a<�Ra<�sa<��a<��a<u�a<��a<��a<��a<��a<��a<��a<h�a<ӵa<�a<S�a<�a<��a<<�a<W�a<��a<��a<��a<�a<��a<��a<;�a<�a<_�a<�a<Uha<9Fa<�#a<a<��`<��`<��`<��`<��`<�`<�`<�a<�4a<�Va<qwa<l�a<��a<{�a<D�a< �a<U�a<��a<I�a<w�a<ۮa<��a<6�a<ǝa<ǜa<\�a<>�a<R�a<C�a<��a<��a<�a<Ͽa<@�a<Ӯa<��a<o�a<�fa<JEa<#"a<��`<��`<��`<ʹ`<o�`<�`<�`<P�`<'�`<� a<["a<�Ca<kca<�~a<+�a<��a<<�a<H�a<G�a<קa<5�a<��a<��a<��a<7�a<�a<w�a<V�a<��a<��a<g�a<�a< �a<�a<��a<�a<��a<w�a<�ga<tIa<�'a<da<��`<��`<�`<y�`<��`<��`< �`<��`<{�`<a<�$a<�  �  �?a<�_a<�{a<��a</�a<I�a<�a<�a<רa<�a<Мa< �a<��a<	�a<o�a<H�a<��a<��a<3�a<B�a<~�a<Ĳa<��a<��a<�a<ʕa<Ma<:ca<�Ba<�a<�`<��`<&�`<�`<��`<�`<��`<��`<��`<��`<.a<�<a<>`a<�a<��a<�a<�a<��a<��a<$�a<�a<��a<(�a<d�a<�a<��a<s�a<r�a<R�a<��a<��a<#�a<�a<��a<�a<f�a<��a<H�a<��a<�ya<Xa<�4a<�a<7�`<��`<��`<��`<�`< �`<�`<h�`<,a<�=a<Gaa<��a<�a<��a<?�a<B�a<q�a<��a<E�a<��a<V�a<1�a<��a<��a<�a<��a<}�a<*�a< �a<��a<��a<p�a<+�a<R�a<�a<��a<��a<��a<�qa<�Na<+a<�a<��`<A�`<��`<P�`<��`<��`<W�`<�a<q&a<Ja<)ma</�a<��a<)�a<Y�a<�a<\�a<��a<{�a<W�a<��a<x�a<��a<d�a<B�a<��a<��a<��a<��a<�a<��a<"�a<N�a<��a<:�a<J�a<�a<D�a<.aa<x=a<�a<��`<\�`<T�`<�`<��`<H�`<J�`<�`<	a<+a<Oa<qa<_�a<��a<��a<9�a<��a<��a<��a<��a<��a<��a<�a<	�a<�a<��a<>�a<k�a<"�a<��a<D�a<��a<��a<��a<h�a<,�a<��a<�a<�`a<�=a<�a<(�`<��`<�`<(�`<��`<
�`<e�`<ǻ`<��`<��`<ua<�<a<t]a< za<d�a<\�a<Ԭa<y�a<*�a<A�a<H�a<Q�a<��a<	�a<+�a<*�a<��a<��a<Y�a<�a<N�a<8�a<��a<�a<�a<��a<ڒa<�}a<�ba<�Ba<�a<��`<��`<e�`<��`<��`<0�`<��`<�`<��`<G�`<S�`<Ca<�  �  ?=a<.^a<�za<�a<ܠa<z�a<��a<[�a<�a<¥a<֟a<��a<��a<�a<��a<;�a<�a<�a</�a<Ϫa<x�a<�a<$�a<ïa<�a<�a<~a<Caa<N@a<�a<��`<��`<
�`<h�`<��`<��`<�`<K�`<j�`<��`<�a<
:a<^a<[~a<��a<b�a<�a<T�a<��a<��a<\�a<��a<P�a<�a<�a<Ʊa<��a<W�a<�a<�a<��a<��a<��a<��a<��a<l�a<��a<a�a<%�a<�wa<8Ua<@1a<(a<!�`<J�`<��`<1�`<W�`<o�`<��`<z�`<�a<T:a<�^a<��a<��a<�a<��a<W�a<��a<��a<9�a<Q�a<Q�a<��a<��a<}�a<�a<��a<`�a<��a<0�a<e�a<�a<��a<��a<��a<��a<��a<��a<�a<�oa<�Ka<�'a<a<��`<��`<3�`<ֹ`<�`<T�`<6�`<� a<#a<�Fa<�ja<b�a<��a<w�a<�a<F�a<
�a<f�a<��a<��a<��a<
�a<`�a<`�a<^�a<�a<��a<�a<��a<��a<��a<g�a<��a<��a<��a<��a<۝a<M�a<�^a<E:a<da<��`<@�`<��`<x�`<+�`<��`<��`<�`<la<=(a< La<�na<эa<��a<�a</�a<��a<��a<9�a<�a<��a<��a<ǵa<��a< �a<�a<#�a<%�a<\�a<��a<��a<j�a<��a<��a<n�a<��a<��a<~a<U^a<�:a<�a<��`<��`<ε`<}�`<�`<r�`<գ`<��`<��`<)�`<9a<�9a<i[a<�xa<��a<Сa<�a<�a<`�a<3�a<ɩa<K�a<�a<�a<�a<K�a<��a<��a<��a<�a<�a<^�a<�a<ҭa<>�a<k�a<5�a<�|a<�`a<t@a<�a<m�`<��`<B�`<}�`<��`<��`<�`<��`<��`<~�`<��`<"a<�  �  �?a<�_a<�{a<��a</�a<I�a<�a<�a<רa<�a<Мa< �a<��a<	�a<o�a<H�a<��a<��a<3�a<B�a<~�a<Ĳa<��a<��a<�a<ʕa<Ma<:ca<�Ba<�a<�`<��`<&�`<�`<��`<�`<��`<��`<��`<��`<.a<�<a<>`a<�a<��a<�a<�a<��a<��a<$�a<�a<��a<(�a<d�a<�a<��a<s�a<r�a<R�a<��a<��a<#�a<�a<��a<�a<f�a<��a<H�a<��a<�ya<Xa<�4a<�a<7�`<��`<��`<��`<�`< �`<�`<h�`<,a<�=a<Gaa<��a<�a<��a<?�a<B�a<q�a<��a<E�a<��a<V�a<1�a<��a<��a<�a<��a<}�a<*�a< �a<��a<��a<p�a<+�a<R�a<�a<��a<��a<��a<�qa<�Na<+a<�a<��`<A�`<��`<P�`<��`<��`<W�`<�a<q&a<Ja<)ma</�a<��a<)�a<Y�a<�a<\�a<��a<{�a<W�a<��a<x�a<��a<d�a<B�a<��a<��a<��a<��a<�a<��a<"�a<N�a<��a<:�a<J�a<�a<D�a<.aa<x=a<�a<��`<\�`<T�`<�`<��`<H�`<J�`<�`<	a<+a<Oa<qa<_�a<��a<��a<9�a<��a<��a<��a<��a<��a<��a<�a<	�a<�a<��a<>�a<k�a<"�a<��a<D�a<��a<��a<��a<h�a<,�a<��a<�a<�`a<�=a<�a<(�`<��`<�`<(�`<��`<
�`<e�`<ǻ`<��`<��`<ua<�<a<t]a< za<d�a<\�a<Ԭa<y�a<*�a<A�a<H�a<Q�a<��a<	�a<+�a<*�a<��a<��a<Y�a<�a<N�a<8�a<��a<�a<�a<��a<ڒa<�}a<�ba<�Ba<�a<��`<��`<e�`<��`<��`<0�`<��`<�`<��`<G�`<S�`<Ca<�  �  tFa<�ea<�a<�a<ϡa<)�a<+�a<��a<�a<b�a<��a<�a<�a<��a<8�a<I�a<��a<M�a<T�a<�a<�a<��a<@�a<�a<�a<l�a<��a<ia<	Ja<�(a<a<�`<��`<S�`<n�`<�`<O�`<h�`<~�`<;�`<�!a<�Da<�fa<�a<�a<۰a<#�a<j�a<S�a<=�a<��a<e�a<{�a<M�a<C�a<��a<E�a<��a<%�a<�a<��a<u�a<�a<�a<X�a<?�a<;�a<f�a<}�a<�a<�_a<�=a<Ha<�`<=�`<&�`<��`<��`<��`<��`<a<`$a<uFa<�ha<��a<b�a<��a<y�a<��a<>�a<��a<��a<��a<��a<�a<��a<��a<��a<��a<ӱa<[�a<��a<��a<��a<��a<4�a<�a<��a<��a<K�a<�a<�xa<&Wa<�4a<�a<��`<?�`<��`<�`<��`<��`<��`<�a<40a<�Ra<�sa<��a<��a<u�a<��a<��a<��a<��a<��a<��a<h�a<ӵa<�a<S�a<�a<��a<<�a<W�a<��a<��a<��a<�a<��a<��a<;�a<�a<_�a<�a<Uha<9Fa<�#a<a<��`<��`<��`<��`<��`<�`<�`<�a<�4a<�Va<qwa<l�a<��a<{�a<D�a< �a<U�a<��a<I�a<w�a<ۮa<��a<6�a<ǝa<ǜa<\�a<>�a<R�a<C�a<��a<��a<�a<Ͽa<@�a<Ӯa<��a<o�a<�fa<JEa<#"a<��`<��`<��`<ʹ`<o�`<�`<�`<P�`<'�`<� a<["a<�Ca<kca<�~a<+�a<��a<<�a<H�a<G�a<קa<5�a<��a<��a<��a<7�a<�a<w�a<V�a<��a<��a<g�a<�a< �a<�a<��a<�a<��a<w�a<�ga<tIa<�'a<da<��`<��`<�`<y�`<��`<��`< �`<��`<{�`<a<�$a<�  �  /Qa<�ma<a�a<+�a<��a<r�a<��a<Y�a<ߘa<ώa<��a<�{a<�ta<pa<�oa<�qa<�wa<�a<�a<�a<y�a<"�a<S�a<ŭa<7�a<6�a<܉a<�qa<IUa<P6a<a<��`<D�`<�`<��`<��`<w�`<��`<?�`<a<G0a<Qa<rpa<I�a<Ǣa<,�a<�a<��a<�a<�a<��a<�a<ŝa<��a<{�a<�a<��a<��a<��a<��a<�a<2�a<��a<j�a<]�a<��a<A�a< �a<��a<��a<�ka<5La<�,a<�a<_�`<=�`<X�`<c�`<d�`<l�`<1a<�4a<bTa<#ta<��a<�a<��a<��a<��a<��a<w�a<��a<�a<i�a<��a<ơa<X�a< �a<	�a<I�a<U�a<��a<��a<a�a<e�a<\�a<�a<�a<��a<��a<ўa<��a<�ca<�Ca<(%a<
a<��`<
�`<
�`<��`<��`<�a<k!a<�?a<�_a<�~a<՚a<A�a<��a<��a<>�a<�a<`�a<�a<�a<o�a<�a<��a<Ҙa<p�a</�a<3�a<ѥa<B�a<��a<��a<x�a<��a<��a<k�a<��a<��a<��a<�sa<�Sa<�3a<�a<|�`<��`<{�`<X�`<!�`<V�`<�a<�$a<�Ca<8ca<C�a<Ûa<۰a<οa<7�a<Q�a<��a<}�a<Y�a<"�a<%�a<��a<o�a<,�a<1�a<n�a<��a<a�a<��a<Q�a< �a<c�a<Ӽa<�a<װa<<�a<��a<Cpa<UQa<�0a<Ta<�`<��`<��`<0�`<{�`<��`<%�`<H�`<a<H0a<wOa<Ula<!�a<;�a<�a<g�a<��a<��a<Şa<b�a<j�a<Ba<�va<�pa<`na<�na<�ra<�ya<k�a<��a<��a<��a<D�a<��a<��a<�a<�a<�oa<�Sa<�4a<�a<��`<��`<r�`<ȷ`<�`<�`<��`<O�`<�`<�a<�1a<�  �  �^a<�wa<R�a<֚a<̢a<i�a<�a<a�a<Z�a<2~a<�pa<#ea<J\a<�Va<�Ua<zXa<�_a<�ia<�va<�a<��a<��a<��a<q�a<3�a<��a<��a<�|a<|ca<�Ga<V+a<�a<��`<�`<��`<��`<��`<��`<@a<�%a<�Ba<�`a<�|a<N�a<��a<��a<:�a<u�a<A�a<�a<��a<[�a<�a<�~a<�wa<ta<�ta<�ya<:�a<ʍa<֛a<6�a<�a<h�a<��a<��a<d�a<��a<B�a<��a<�za<i^a<,Ba<j(a<ha<�a<]�`<I�`<ya<�a<^.a</Ia<�ea<��a<��a<�a<`�a<D�a<��a<.�a<��a<j�a<4�a<��a<�a<�a<�a<8�a<?�a<��a<��a<Z�a<��a<w�a<�a<n�a<��a<��a<��a<[�a<��a<#�a</ta<9Wa<9;a<�"a<Za<�a<�`<�a<Ra<�a<�7a<[Sa<(pa<<�a<��a<4�a<]�a<��a<3�a<��a<e�a<��a<c�a<��a<n�a<�a<a<�}a<�a<#�a<��a<!�a<��a<¶a<M�a<,�a<X�a<b�a<�a<@�a<��a<Ła<ea< Ha<�,a<�a<|a<F�`<c�`<��`<�a<� a<":a<&Va<�ra<��a<ʤa<Ѷa<R�a<_�a<�a<F�a<g�a<��a<o�a<L�a<y~a<~ua<Npa<Ooa<Rra<Rya<3�a<��a<U�a<��a<`�a<+�a<��a<��a<ئa<0�a<I|a<�`a<�Ba<�%a<�
a<��`<*�`<4�`<_�`<��`<��`<ta<�%a<�Aa<�]a<�wa< �a<�a<h�a<i�a<A�a<>�a<q�a<��a<�va<|ia<_a<�Wa<}Ta<$Ua<:Za<�ba<Dna<�{a<׈a<(�a<V�a<C�a<o�a<7�a<��a<�ya<aa<�Da<�'a<�a<?�`<�`<_�`<��`<��`<r�`<�`<O	a<2%a<JBa<�  �  ]ma<Ղa<q�a<�a<G�a<�a<��a<�a<{a<�ia<+Ya<�Ja<q?a<�8a<�6a<:a<Ca<�Oa<�_a<vqa<L�a<]�a<�a<ݧa<��a<��a<�a<��a<�ra<�Za<YBa<+a<Ta<�a<� a< a<ga<�a<�&a<2>a<�Wa<ra<`�a<�a<�a<��a<s�a<Ƕa<r�a<B�a<X�a<�a<Cpa<Nca<Za<�Ua<;Va<�[a<|fa<�ta<�a<$�a<�a<"�a<��a<~�a<�a<��a<��a<��a<�a<sa<_Za<yCa<�0a<�#a<�a<ma<�&a<�4a<�Ha<�`a<�ya<��a<.�a<N�a<��a<�a<��a<*�a<}�a<X�a<+�a<�a<Aza<�ma<	ea<taa<�ba<�ia<�ta<U�a<5�a<��a<,�a<��a<��a<��a<��a<�a<B�a<s�a<f�a<ma<�Ta<�>a<y-a<�"a<]a<�!a<�+a<<a<UQa<�ia<Ăa<�a<�a<T�a<��a<p�a<��a<�a<�a<��a<�a<�a<�sa<:ha<�`a<�^a<�aa<�ia<�ua<�a<�a<G�a<��a<��a<��a<��a<3�a<:�a<��a<A�a<{xa<#_a<Ga<�2a<S#a<[a<�a<a<?*a<;<a<�Ra<9ka<&�a<7�a<��a<��a<T�a<��a<c�a<y�a<��a<�a<�a<�qa<�ba<Xa<�Qa<�Pa<�Ta<�]a<9ja<�ya<A�a<n�a<�a<�a<z�a<��a<1�a<{�a<p�a<rqa<~Wa<�=a<�%a<Sa<�a<k�`<��`<�a<�a<�%a<=a<�Ua<�ma<��a<��a<��a<8�a<K�a<B�a<�a<f�a<�qa<`a<�Oa<�Ba<�9a<�5a<�6a<0=a<�Ga<CVa<�fa<xa<O�a<~�a<h�a<}�a<�a<(�a<?�a<Noa<%Wa<�=a<$%a<+a<�`</�`<&�`<t�`<��`<Qa<�"a<e;a<�Ta<�  �  H|a<��a<�a<��a<��a< �a<Ǎa<�|a<�ha<^Sa<?a<R-a<�a<�a<ta<�a<�#a<43a<xFa<�[a<�qa<
�a<�a<�a<Ĩa<�a<�a<*�a<ނa<�na<Za<Fa<�5a<l)a<�"a<�!a<�'a<3a<vCa<�Wa<�ma<ăa<֗a<��a<��a<ĸa<S�a<��a<�a<��a<�|a<	ha<Ua<(Ea<�9a<94a<�4a<�;a<Ha<AYa<�ma<��a<ʙa<D�a<��a<��a<��a<��a<��a<��a<9�a<d�a<\sa<`a<Pa<�Da<w?a<;@a<6Ga<�Sa<�da<�xa<=�a<��a<7�a<N�a<��a<��a<+�a<��a<��a<W�a<��a<qa<�]a<�Na<mDa<�?a<�Aa<�Ia<Wa<�ha<A}a<�a<e�a<1�a<n�a<��a<��a<*�a<��a<�a<#�a<��a<�na<\a<nMa<Da<Z@a<*Ca<�Ka<�Ya<�ka<��a<��a<ީa<ܺa<��a<�a<��a<��a<+�a<��a<O�a<�}a<�ha<�Va<�Ha<�?a<(=a<�@a<gJa<!Ya<�ka<z�a<ӕa<L�a<��a<��a<��a<��a<��a<)�a<#�a<��a<�va<�ba<�Pa<�Ca<$<a<�:a<N?a<�Ia<Ya<la<�a<�a<��a<�a<��a<n�a<}�a<+�a<�a<��a<d�a<ka<sVa<�Da<�7a<t0a<H/a<l4a<"?a<�Na<�aa<va<M�a<8�a<e�a<�a<,�a<�a<z�a<g�a<��a<�la<�Va<hBa<�1a<�%a<Ha<La<�%a<[1a<�Aa<,Ua<$ja<M~a<�a<��a<a�a<ڦa<Сa<��a<8�a<kra<�\a<Ga<�3a<�#a<'a<?a<�a<Sa<X*a<�;a<�Oa<Qea<�ya<�a<�a<K�a<	�a<I�a<��a<�}a<�ia<;Ta<\?a<�,a<a<�a<a<a<�a<&+a<�=a<MRa<ha<�  �  O�a<D�a<��a<�a<�a<L�a<ɂa<�ma<UUa<D<a<?$a<Za<��`<��`<��`<\�`<a<�a<v,a<�Ea<g_a<�wa<��a<�a< �a<��a<��a<Ξa<�a<�a<4qa<'aa<kSa<]Ia<�Ca<iCa<Ha<�Qa<�_a<[pa<w�a<��a<p�a<Ӱa<�a<�a<J�a<J�a<̕a<�a<�ga<�Oa<9a<V&a<)a<la<�a<�a<�(a<�<a<Ua<�na<��a<��a<9�a<s�a<H�a<��a<t�a<ݻa<��a<לa<a<�{a<�na<\ea<�`a<�aa<Qga<�qa<�a<D�a<��a<o�a<V�a<M�a<��a<W�a<��a<�a<�a<S�a<pa<eWa<�@a</a<#a<�a< a<P)a<�8a<�Ma<�ea<a<��a<ƭa<#�a<��a<��a<X�a<��a<z�a<Ϊa<v�a<L�a<�xa<�la<�da<�aa<da<qka<�va<�a<іa<�a<�a<��a<��a<��a<�a<�a<,�a<{�a<�a<ffa<�Ma<�8a<C(a</a<.a<va<�*a<�;a<�Qa<&ja<R�a<�a<��a<ܾa< �a<��a<F�a<ʽa<&�a<��a<��a<-}a<�na<�ca<X]a<\a<�_a<�ha<9ua<�a<ٕa<��a<N�a<Y�a<�a<��a<v�a<�a<םa<_�a<�la<�Ra<p:a<&a<a<�a<ra<sa< a<I2a<�Ha<�`a<?ya<~�a<��a<j�a<մa<��a<Y�a<��a<�a<9�a<oa<&^a<%Pa<�Ea<�@a<�@a<�Ea<\Oa<�\a<�la<�}a<ȍa<#�a<��a<J�a<��a<c�a<�a<�xa<m`a<�Fa<�-a<�a<>a<��`<P�`<��`<��`<a<� a<j8a<}Qa<�ia<�a<ѐa<+�a<�a<s�a<˗a<J�a<�{a<ja<�Xa<qIa<`=a<t5a<�2a<�4a<z<a<6Ha<fWa<�ha<'za<�  �  ��a<t�a<�a<R�a<k�a<�a<�wa<�^a<�Ba<�%a<�
a<��`<�`<�`<I�`<��`<�`<�`<\a<�/a<iMa<�ia<��a<��a<b�a<��a<��a<�a<�a<��a<'�a<Qya<{na<�fa<ba<ba<�ea<�ma<ya<ʆa<=�a<\�a<h�a<��a<Һa<�a<��a<��a<H�a<�oa<�Sa<8a<ja<<	a<�`<D�`<��`<]�`<�a<�!a<=a<jZa<xa<��a<(�a<Q�a<��a<��a<��a<e�a<��a<&�a<ءa<�a<��a<�a<�a<�a<��a<�a<7�a<��a<�a<�a<��a<��a<�a< �a<��a<�a<$�a<�wa<�Za<�>a<c%a<>a<ya<��`<��`<�
a<2a<�3a<�Na<�ka<w�a<�a<\�a<��a<��a<,�a<��a<X�a<~�a<*�a<��a<�a<c�a<�a<��a<E�a<7�a<p�a<u�a<�a<0�a<+�a<��a<��a<��a<��a<��a<�a<��a<ma<�Oa<-4a<0a<�	a<7�`<��`<��`<�a<�a<�8a<~Ta<Mqa<��a<�a<k�a<|�a<�a<N�a<��a<5�a<|�a<�a<W�a<��a<�a<�{a<�za<�}a<��a<��a<[�a<��a<��a<I�a< �a<��a<��a<��a<L�a<U�a</va<�Xa<5;a<�a<�a<��`<��`<@�`<'�`<�a<ca<�0a<�La<�ha<��a<��a<F�a<j�a<$�a<��a<�a<v�a<��a<-�a<Kwa<la<�ca<`_a<_a<ca<�ja<Jua<�a<�a<L�a<��a<�a<کa<V�a<g�a<�a<�ja<�Na<l1a<�a<�`<u�`<A�`<�`<��`<6�`<}�`<~a<�!a<F>a<�Za<ta<
�a<D�a<�a<C�a<��a<"�a<*�a<�}a<
pa<�ca<�Ya<{Sa<nQa<Sa<:Ya<�ba<�na<�|a<>�a<�  �  P�a<Υa<��a<ޡa<��a<ׄa<.ma<�Pa<�1a<a<�`<�`<L�`<V�`<=�`<�`<��`<��`<t�`<�a<e=a<�\a<�xa<*�a<I�a<��a<C�a<��a<�a<�a<S�a<��a<Q�a</a<�{a<�{a<Ba<��a<��a<Y�a<��a<}�a<��a<μa<��a<X�a<��a<}�a<�}a<aa<1Ba<R#a<a<��`<��`<S�`<��`<%�`<��`<`
a<�'a<dHa<ia<Ƈa<��a<�a<��a<m�a<��a<��a<��a<U�a<�a<L�a<�a<A�a<y�a<ݙa<��a<�a<�a<'�a<��a<��a<[�a<��a<��a<h�a<��a<��a<��a<�ga<Ha<�(a<;a<��`<�`<��`<3�`<��`<a<�a<�:a<�Za<nza<W�a<�a<��a<��a<��a<��a<��a<r�a<O�a<ϲa<>�a<��a<w�a<��a<��a<��a<ԧa<�a<i�a<��a<��a<�a<��a<j�a<��a<��a<��a<�{a<b\a<*<a<�a<=a<��`<�`<��`<�`<�`<�a<�"a<fAa<Baa<�a<z�a<��a<_�a<Y�a<��a<��a<��a<��a<�a<��a<��a<��a<|�a<��a<��a<u�a<^�a<�a<(�a<��a<��a<Z�a<��a<	�a<��a<!�a<օa<�ga<�Fa<k&a<{a<A�`<��`<��`<A�`<��`<��`<��`<�a<}:a<�Ya<�va<�a<ڣa<z�a<��a<��a<<�a<0�a<��a<e�a<��a<��a<�|a<Bya<�xa<�{a<ȁa<��a<��a<x�a<3�a<,�a<�a<��a<��a<H�a<�ya<6^a<&?a<�a<�`<��`<$�`<Ѽ`<�`<5�`<J�`<O�`<��`<va<=-a<�La<?ia<��a<	�a<�a<��a<u�a<{�a<�a<��a<Q�a<�ya<ra<ma<Qka<�la<�qa<ya<��a<%�a<��a<�  �  R�a</�a<K�a<	�a<1�a< a<�da<Fa<�$a<ua<t�`<��`<��`<�`<Y�`<ʧ`<%�`<��`<?�`<�a<�0a<�Ra<Cqa<�a<��a<��a<|�a<��a<%�a<��a<D�a< �a<h�a<Ǒa<��a<��a<i�a<��a<�a<h�a<q�a<f�a<�a<F�a<U�a<��a<U�a<͏a<�ta<kUa<4a<
a<��`<��`<��`<��`<�`<�`<��`<��`<ma<	:a<%]a<l~a<��a<q�a<�a<��a<��a<u�a<Y�a<��a<��a<Z�a<��a<F�a<�a<{�a<=�a<T�a<�a<X�a<Y�a<��a<��a<X�a<��a<��a<��a<5�a<�|a<�[a<'9a<�a<\�`<��`<��`<��`<��`<��`<k�`<�
a<�*a<SMa<Poa<َa<ɩa<�a<��a<��a<��a<q�a<�a<��a<g�a<ݹa<��a<ݯa<?�a<n�a<زa<��a<�a<��a<f�a<��a<y�a<8�a<��a<[�a<Ūa<N�a<
qa<&Oa<�,a<a<��`<N�`<�`<��`<��`<��`<q�`<ka<;2a<�Ta<�ua<��a<��a<��a<�a<'�a<��a<d�a<�a<�a<�a<��a<5�a<�a<A�a<'�a<?�a<��a<��a<��a<��a< �a<��a<}�a<n�a<��a<t�a<�|a<�[a<�8a<$a<A�`<X�`<��`<�`<��`<��`<��`<V�`<'a<!,a<�Ma<Zma<�a<b�a<��a<	�a<��a<�a<εa<�a<+�a<��a<$�a<ُa<ٌa<��a<��a<�a<��a<Ӡa<B�a</�a<t�a<��a<p�a<*�a<F�a<fra<=Ta<�2a<�a<�`<�`<ѷ`<��`<-�`<��`<��`<��`<��`<��`<�a<xAa<�`a<u{a<c�a<�a<�a<��a<2�a<��a<�a<�a<U�a<%�a<i�a<�~a<7�a<σa<щa<b�a<��a<m�a<�  �  ��a<۬a<X�a<S�a<Ґa< {a<V_a<1?a<a<��`<)�`<[�`<z�`<"�`<��`<�`<8�`<~�`<Q�`<+a<�(a<�Ka<�ka<>�a<t�a<P�a<Գa<�a<˵a<ʱa<C�a<q�a<J�a<z�a<��a<ʛa<W�a<Ţa<�a<	�a<i�a<��a<��a<Z�a<ӽa<e�a<{�a<?�a<�na<�Ma<'+a<�a<(�`<�`<k�`<ٲ`<-�`<|�`<�`< �`<�a<�0a<�Ua<?xa<�a<n�a<��a<$�a<��a<�a<x�a<��a<W�a<<�a<�a<-�a<D�a<��a<	�a<^�a<�a<��a<��a<��a<��a<��a<��a<�a<�a<�a<va<�Sa<�/a<'a<O�`<��`<�`<��`<��`<��`<��`<}�`<� a<�Da<=ha<�a<��a<b�a<��a<��a<!�a<��a<��a<��a<]�a<;�a<#�a<�a<y�a<z�a<h�a<0�a<�a<��a<G�a<J�a<'�a<F�a<��a<��a<Ŧa<��a<$ja<�Fa<�"a<� a<��`< �`<B�`<!�`<�`<��`<K�`<za<�(a<eLa<oa<o�a<�a<��a<��a<}�a< �a<	�a<O�a<�a<x�a<��a<�a<-�a<y�a<�a<��a<��a<��a<��a<��a<��a<��a<��a<�a<��a<�a<�va<nTa<�/a<�a<��`<��`<a�`<�`<��`<F�`<�`<��`<� a<#a<
Fa<-ga<\�a<^�a<�a<M�a<��a<��a<�a<�a<��a<��a<X�a<��a<
�a<��a<`�a<�a<+�a<�a<��a<�a<��a<�a<N�a<A�a<ևa<Dma<�Ma<�*a<ja<X�`<�`<��`<�`<`�`<�`<:�`<R�`<~�`<��`<a<e:a<�Za<Awa<Սa<#�a<�a<�a<X�a<[�a<{�a<ؚa<��a<��a<k�a<�a<@�a<\�a<\�a<��a<:�a<L�a<�  �  l�a<��a<v�a<��a<��a<�sa<^a<Fa<k+a<�a<��`<��`<2�`<Z�`<��`<��`<��`<�`<, a<la<�5a<Qa<�ia<�~a<X�a<@�a<��a<ϥa<��a<'�a<,�a<ƚa<��a<�a<�a<Y�a<C�a<�a<�a<��a<I�a<�a<�a<��a<ݬa<E�a<U�a<c�a<�oa<Wa<�<a<F#a<�a<��`<��`<��`<T�`<a�`<�`<_a<*(a<1Ca<_a<�ya<8�a</�a<!�a<��a<O�a<%�a<��a<r�a<ݼa<)�a<�a<&�a<��a<0�a<�a<f�a<Թa<�a<��a<��a<�a<��a<��a<�a<n�a<8�a<�ya<T_a<PDa<q*a<ja<a<��`<S�`<��`<�`<)a<Y a<z9a<4Ta<Loa<[�a<B�a<��a<ϼa<G�a<�a<r�a<��a<��a<��a<�a<�a<g�a<|�a< �a<H�a< �a<��a<t�a<��a<T�a<(�a<��a<��a<%�a<ܞa<1�a<[pa<GUa<S:a<� a<�
a</�`<��`<��`<0�`<��`<Ca<�$a<S>a<*Ya<�sa<f�a<��a<گa<�a<��a</�a<Q�a<�a<T�a<(�a<��a<٭a<իa<S�a<K�a<��a<�a<n�a<�a<��a<'�a<��a<r�a<p�a<�a<��a<zwa<-]a<[Aa<.&a<a<A�`<��`<.�`<��`<^�`<]�`<a<Ia<�5a<Pa<7ia<?a<ʑa<]�a<��a<��a<��a<�a<��a<�a<[�a<c�a<��a<��a<�a<�a<ݓa<��a<#�a<C�a<�a<��a<�a<�a<Îa<�~a<ja<Ra<'7a<�a<La<��`<�`<b�`<q�`<T�`<|�`<2�`<�`<�a<Y'a<-Ba<�Za<�pa<-�a<Ўa<�a<a<��a<U�a<	�a<�a<?�a<D�a<Ƀa<��a<��a<�a<��a<̎a<�a<r�a<�  �  1�a<��a<L�a<�a<3�a<�ta<�_a<�Ga<�-a<ra<��`<��`<y�`<��`<b�`<W�`<�`<2�`<�a<�a<�7a<vRa<�ja<�a<Џa<q�a<e�a<�a<^�a<r�a<.�a<��a<9�a<1�a<��a<ӏa<7�a<�a<T�a<Z�a<k�a<��a<�a<B�a<Ҭa<��a<��a<��a<!qa<�Xa<B?a<�%a<�a<��`<H�`<��`<�`<��`<0�`<la<�*a<�Ea<�`a<{a<b�a<ۥa<��a<��a<��a<4�a<X�a<��a<��a<��a<;�a<,�a<w�a<ˬa<�a<��a<��a<ۼa<��a<��a<I�a<��a<ӿa<T�a<!�a<i�a<{a<Saa<�Fa<5-a<�a<Ta<P�`<�`<A�`<k�`<Ia<@#a<<a<�Va<�pa<��a<-�a<��a</�a<*�a<��a<J�a<U�a<��a<r�a<E�a<��a<;�a<�a<ܮa<X�a<Q�a<M�a<��a<�a<�a<��a<��a<�a<��a<��a<u�a<�qa<�Wa<�<a<�#a<a<x�`<o�`<Q�`<��`<��`<`a<�'a<�@a<<[a<	ua<��a<��a<R�a<?�a<}�a<s�a<�a<\�a<V�a<�a<ήa<�a<z�a<ͧa<>�a<�a<O�a<;�a<%�a<
�a<%�a<3�a<f�a<�a<��a<��a<�xa<�^a<�Ca<�(a<a<g�`<>�`<��`<��`<��`<��`<%a<�a<98a<�Qa<�ja<j�a<v�a<Пa<��a<��a<��a<��a<Ȥa<ٞa<ؘa<��a<��a<�a<��a<-�a<�a<S�a<�a<��a<��a<Ƣa<��a<;�a<4�a<za<>ka<fSa<$9a<4a<a<��`<E�`<��`<+�`<��`<��`<R�`<��`<|a<�)a<�Ca<D\a<�qa<��a<0�a<��a<9�a<ՙa<Ɩa<%�a<Ìa<��a<S�a<��a<na<z�a<!�a<N�a<��a<�a<זa<�  �  ��a<��a<%�a<a�a<Ɇa<xwa<�ca<�La<�3a<�a<�a<��`<%�`<��`<U�`<+�`<��`<!�`<�
a<$a<�=a<[Wa<�na<�a<)�a<q�a<��a<}�a<��a<q�a<ݖa<?�a<�a<��a<��a<݆a<o�a<��a<��a<��a<ءa<F�a<ͬa<V�a<�a<|�a<��a<߉a<�ua<E^a<�Ea<{-a<ea<a<�`<��`<��`<~�`<�a<a<u2a<tLa<�fa<�a<ޕa<��a<��a<�a<�a<?�a<@�a<"�a<�a<�a<ڨa<j�a<��a<�a<^�a<r�a<.�a<i�a<��a<��a<��a<�a<��a<��a<��a</�a<�a<8ga<�Ma<5a<da<�a<!a<��`<%�`<%a<xa<�+a<hCa<�\a<va<�a<3�a<>�a<��a<&�a<_�a<��a<��a<�a<y�a<n�a<��a<c�a<��a<��a<ͨa<d�a<9�a<~�a<a�a<��a<G�a<]�a<=�a<E�a<��a<��a<wa<�]a<Da<�+a<4a<%a<U�`<G�`<��`<g	a<Qa<�/a<�Ga<@aa<�ya<��a<I�a<��a<@�a<�a<��a<S�a<[�a<�a<��a<��a<Q�a<��a<מa<u�a<��a<��a<|�a<��a<ʹa<�a<G�a<��a<��a<��a<�a<E}a<cda<oJa<b0a<�a<�a<�`<��`<��`<{�`<��`<�a<�&a< ?a<�Wa<oa<�a<��a<��a<��a<ªa<��a<��a<U�a<3�a<P�a<#�a<׆a<"�a<��a<��a<�a<�a<��a<Y�a<�a<�a<	�a<�a<k�a<�a<oa<*Xa<?a<5%a<�a<��`<��`<��`<�`<��`<��`<��`<T�`<�a<0a<�Ha<�`a<�ta<r�a<��a<��a<�a<}�a<=�a<G�a<ͅa<�a<�za<�wa<uva<�wa<�za<ca<t�a<��a<+�a<�  �  �a<�a<��a<��a<�a<�{a<�ia<�Ta<�=a<4&a<a<��`<s�`<��`<��`<��`<��`<a<�a<"/a<]Ga<_a<ta<��a<�a<E�a<��a<c�a<��a<;�a<�a<��a<Ia<bza<�wa<.xa<�za<6�a<��a<�a<Әa< �a<ȧa<o�a</�a<]�a<Ҝa<i�a<7|a<ga<Pa<�9a<�$a<�a<�a<�a<a<1	a<Ka<�(a<�>a<�Va<loa<��a<��a<�a<��a<O�a<p�a<l�a<P�a<O�a<��a<�a<��a<זa<єa<*�a<�a<u�a<m�a<L�a<Q�a<f�a<A�a<��a<H�a<�a<�a<\�a<M�a<upa<�Xa<�Aa<7-a<�a<�a<=a<a<�a<�%a<�8a< Oa<�fa<n~a<��a<n�a<��a<�a<��a<��a<|�a<2�a<y�a<n�a<��a<ța<��a<B�a<A�a<�a<͠a<�a<�a<��a<�a<��a<��a<u�a<~�a<��a<y�a<a<}ga<�Oa<9a<d%a<va<@a<�
a<]a<�a<F(a<N<a<Sa<�ja<��a<�a<�a<m�a<�a<�a<Ƽa<+�a<&�a<�a<
�a<ݙa<!�a<ڐa<'�a<Αa<;�a<y�a<Уa<��a<��a<�a<^�a<��a<��a<��a<��a<�a<ma<�Ta<�<a<&a<Na<�a<��`<��`<-a<�a<fa<�2a<gIa<n`a<va<��a<��a<١a<;�a<�a<ߤa<��a<��a<��a<G�a<�}a<Exa<pua<ua<)wa<�{a<A�a<��a<�a<q�a<��a<Ҝa<��a<�a<\�a<,ta<�_a<AHa<0a<�a<�a<��`<l�`<V�`<��`<��`<��`<�a<�"a<�9a<OQa<�fa<�xa<�a<�a<��a<��a<�a<��a<܂a<�za<Ksa<"ma<ia<�ga<�ha<�la<�ra<Aza<c�a<`�a<�  �  D�a<��a<�a<��a<��a<a<Yqa<�^a<Ja<�4a<� a<Xa<$a<�`< �`<#�`<8a<.a<(a<G=a<CSa<�ha<{a<n�a<�a<��a<��a<��a<-�a<g�a<�a<%va<na<ha<�da<�da<ha<�na<wa<��a<��a<��a<Πa<��a<k�a<0�a<X�a<t�a<��a<�qa<C]a<Ia<86a<�&a<�a<a<�a<"a<^)a<5:a<mNa<;da<�za<2�a<�a<֮a<��a<ֻa<?�a<��a</�a<��a<��a<ڑa<
�a<:�a<��a<��a<��a<"�a<��a<�a<:�a<ɲa<(�a<S�a<f�a<ιa<w�a<5�a<��a<|a<�fa<�Qa<&?a<80a<&a<�!a<�#a<W+a<g8a<�Ia<^a<psa<��a<כa<�a<��a<S�a<o�a<�a<��a<1�a<�a<��a<,�a<̉a<��a<��a<;�a<Ԉa<׏a<��a<;�a<H�a<&�a<M�a<!�a<n�a<�a<ܫa<�a<(�a<�sa<O^a<�Ia<�7a<,*a<�!a<a<�"a<,a<g:a<�La<;aa<�va<!�a<�a<��a<r�a<x�a<׺a<��a<ׯa<S�a<��a<��a<��a<΁a<�}a<�|a<a<��a<�a<��a<��a<8�a<�a<�a<��a<W�a<�a<��a<G�a<�wa<�aa<�Ka<{7a<8&a<�a<ca<>a<a<� a<�/a<�Ba<�Va<�ka<�~a<�a<u�a<��a<ĥa<�a<1�a<~�a<�a<�a<ua<Vla<�ea<.ba<�aa<�da<�ja<{ra<|a<؅a<Ԏa<��a<A�a<ɘa<��a<ɉa<{a<�ha<�Sa<�=a<�(a<�a<a<}�`<��`<@�`<��`<ia<�a<s1a<�Fa<�[a<zna<U~a<ԉa<Y�a<I�a<��a<��a<��a<{va<la<�ba<+[a<#Va<�Ta<�Ua<�Za<�aa<;ka<�ua<�a<�  �  �a<Z�a<r�a<@�a<�a<��a<�ya<ja<GXa<{Ea<�3a<m$a<�a<�a<�a<�a<�a<�)a<�:a<fMa<�`a<�ra<��a<�a<��a<��a<��a<z�a<�a<U|a<�oa<�ca<�Ya<BRa<3Na<Na<�Qa<YYa<�ca<�pa<�~a<a�a<K�a<��a<�a<ϧa<~�a<ߚa<��a<�}a<{la<[Za<�Ia<N<a<�2a<�-a<[.a<V4a<??a<*Na<`a<�sa<�a<ɘa<��a<L�a<��a<ɹa<�a<��a<'�a<��a<ߊa<�~a<�ta<$na<�ja<Bka<�oa<zwa<F�a<��a<Λa<U�a<��a<۹a<�a<V�a<��a<��a<��a<T�a<�va<da<�Sa<hFa<w=a<�9a<B;a<#Ba<�Ma<]a<�na<�a<:�a<��a<��a</�a<N�a<G�a<ҷa<��a<$�a<�a<3�a<�}a<Tta<Tna<la<�ma<5sa<�{a<G�a<�a<�a<��a<�a<��a<�a<f�a<�a<��a<R�a<,�a<�na<�\a<�La<�@a<J9a<�6a<:a<eBa<Oa<%_a<_qa<(�a<��a<�a<3�a<C�a<�a<��a<�a<��a<A�a<�a<_a<=ta<�ka<ga<�ea<�ha<Zoa<�xa<��a<9�a<ߝa<��a<p�a<��a<��a</�a<�a<��a<�a<�pa<@]a<2Ka<�;a<�0a< *a<�(a<S-a<�6a<�Ca<,Ta<Bfa<xa<L�a<a<�a<�a<��a<ʞa<�a<x�a<�|a<oa<4ba<LWa<�Oa<YKa<"Ka<�Na<�Ua<`a<�ka<lxa<_�a<6�a<Ɣa<w�a<-�a<�a<��a<�ra<aa<�Ma<�:a<�)a<Ka<�a<�a<�a<wa<�!a<�0a<MBa<-Ua<ga<Iwa<�a<f�a<V�a<$�a<��a<T�a<�ta<rga<�Za<�Na<�Ea<�?a<�=a<q?a<Ea<�Ma<�Ya<lfa<�sa<�  �  �ta<��a<��a<
�a<�a<1�a<E�a<lua<�fa<�Va<Ha<�:a<z0a<�*a<)a<a,a<�3a<�?a<2Na<6^a<�na<�}a<��a<m�a<&�a<��a<u�a<5�a<[|a<�ma<a^a<Pa<�Ca<j:a<�5a<;5a<�9a<RBa<Oa<(^a<�na<ma<t�a<#�a<��a<§a<��a<�a<j�a<|�a<�{a<�la<_a<Sa<�Ja<�Fa<sGa<�La<$Va<{ca<�ra<��a<ݓa<��a<S�a<̵a<�a<��a<�a<�a<z�a<�a<�xa<Rja<,^a<�Ua<�Qa<�Ra<�Wa<aa<$na<�|a<�a<Z�a<�a<s�a<��a<g�a<θa< �a<&�a<�a<�a<xwa<\ia<�]a<!Va<�Ra<6Ta<
Za<%da<�qa<��a<��a<�a<g�a<�a<��a<|�a<�a<��a<"�a<��a<��a<va<ha<�\a<�Ua<(Sa<MUa<�[a<@fa<�sa<�a<�a<��a<j�a<-�a<�a<��a<M�a<��a<��a<��a<m�a<qa<;ca<�Xa<2Ra<Pa<�Ra<�Ya<ea<�ra<6�a<�a<e�a<��a<��a<��a<��a<��a<��a<�a<֊a<�za<}ka<^a<%Ta<tNa<.Ma<�Pa<PXa<da< ra<h�a<�a<��a<�a<�a<�a<Y�a<P�a<�a<��a<�a<�oa<G`a<�Ra<�Ha<)Ca<Ba<�Ea<~Ma<7Ya<�fa<va<�a<�a<a�a<n�a<3�a<��a<��a<��a<�}a<Uma<�\a<�Ma<}@a<r7a<�2a<w2a<�6a<�?a<�Ka<"Za<�ia<bxa<��a<\�a<�a<;�a<�a<�a<f}a<�na<P^a<>Na<�?a<�3a<�+a<�'a<�(a<Z.a< 8a<KEa<Ta<da<�ra<	�a<|�a<�a<��a<��a<q�a<�ua<ga<�Va<mGa<|9a<P.a<h'a<�$a<'a<|-a<Q8a<-Fa<�Ua<�ea<�  �  �ia<�ya<��a<	�a<~�a<ԏa<�a<��a<�ta<�ga<�[a<uPa<Ha<Ca<�Aa<�Da<CKa<Ua<8aa<�na<#|a< �a<��a<k�a<Øa<��a<��a<I�a<ipa<�^a<lLa<p;a<-a<r"a<�a<a<!a<)+a<k9a<�Ja<g^a<�qa<6�a<��a<��a<�a<C�a<��a<E�a<��a<�a<�~a<Gsa<�ia<�ba<�_a<4`a<�da<�la<xa<�a<˒a<^�a<Ϋa<4�a<��a<n�a<��a<?�a<1�a<h�a<xa<�ea<�Ta<-Ga<�=a<�8a<�9a<�?a<oJa<2Ya<�ja<�}a<�a<Ѡa<f�a<��a<��a<{�a<��a<0�a<�a<�a<=�a<o~a<�ta<gna<�ka<�la<�qa<2za<b�a<�a<;�a<}�a<x�a<�a<y�a<ٻa<s�a<̨a<6�a<��a<�ta<.ba<Ra<eEa<'=a<�9a<m<a<�Ca<Pa<�_a<�qa<��a<c�a<*�a<&�a<�a<��a<�a<��a<�a<��a<k�a<��a<ya<7pa<�ja<�ha<5ka<+qa<\za<�a<��a<�a<Ϊa<��a<��a<X�a<ܴa<�a<��a<�a<�{a<�ha<�Va<�Ga<,<a<|5a<4a<8a<%Aa<ZNa<�^a<qa<x�a<l�a<ݢa<�a<�a<�a<߯a<�a<��a<i�a<��a<�ta<!ia<�`a<�[a<�Za<�]a<2da<�ma<%ya<\�a<d�a<T�a<C�a<e�a<��a<�a<�a<��a<�pa<[]a<�Ia<8a<�)a<�a<ua<ta<�a<�(a<7a<�Ga<PZa<la<G|a<M�a<�a<w�a<Õa<s�a<l�a<�{a<Nna<�`a<�Ta<�Ja<�Ca<�@a<oAa<!Fa<)Na<Ya<fea<Wra<[~a<�a<o�a<��a<�a<W�a<�za<�ja<	Ya<�Ea<�3a<{#a<�a<�a<�a<(a<�a<'"a<	2a<IDa<}Wa<�  �  �^a<Hqa<�a<܋a<��a<y�a<��a<?�a<_�a<jwa<Qma<zda<�]a<�Ya<�Xa<[a<�`a<�ha<�ra<n}a< �a<*�a<{�a<a�a<��a<H�a<�a<Uwa<�da<Pa<t;a<(a<�a<�a<�a<Ta<�	a<a<%a<�8a<�Na<�da<:za<��a<��a<��a<êa<S�a<ۧa<=�a<��a<�a<Ņa<H~a<�xa<Kva< wa<�za<ˁa<��a<��a<��a<>�a<��a<)�a<��a<^�a<Q�a<>�a<x�a<�}a<�ha<�Sa<�@a<51a<=&a<	!a<�!a<�(a<�4a<�Ea<mYa<�na<�a<��a<0�a<��a<2�a<�a<N�a<�a<��a<��a<Y�a<��a<�a<��a<��a<f�a<��a<~�a<o�a<ԡa<!�a<��a<d�a<��a<H�a<�a<��a<��a<��a<�ya<?da<�Oa<K=a<�.a<�%a<3"a<�$a<f-a<;a<�La<6aa<�va<a�a<̝a<�a<��a<v�a<��a<;�a<��a<N�a<�a<a�a<�a<�a<5�a<�a<��a<��a<؍a<;�a<z�a<a�a<ݳa<}�a<��a<7�a<)�a<�a<a<u�a<ma<�Wa<wCa<+2a<O%a<�a<Ca<� a<+a<:a<�La<Eaa<qva<m�a<��a<�a<��a<n�a<��a<��a<S�a<�a<��a<�a<�}a<�va<�ra<�qa<�sa<&ya<{�a<��a<Q�a<E�a<D�a<9�a<A�a<��a<G�a<�a<�xa<da<�Ma<8a<$a<�a<�a<�a<�a<�a<Qa<n#a<�6a<>Ka<`a<sa<�a<�a<��a<\�a<�a<�a<I�a<�|a<ra<�ga<�_a<Za<�Wa<Xa<�[a<rba<ka<2ua<<a<]�a<�a<m�a<��a<��a<��a<�ra<0`a<DKa<�5a<
!a<�a<o a<�`<��`<��`<P�`<,a<4a<�3a<_Ia<�  �  �Ta<�ia<�{a<i�a<(�a<A�a<�a<*�a<ˋa<)�a<w|a<ua<�oa<�la<la<�ma<�ra<3ya<&�a<��a<֑a<��a<d�a<��a<4�a<3�a<M�a<Zoa<PZa<RCa<j,a<�a<�a<��`<y�`<��`<��`<�a<Ka<�(a<�@a<|Ya<qa<�a<A�a<�a<ʫa<�a<�a<��a<��a<��a<��a<��a<@�a<��a<A�a<f�a<H�a<ۚa<f�a<6�a<9�a<D�a<2�a<�a<�a<S�a<Ǜa<��a<~ra<�Za<Da<%/a<a<Aa<{a<La<�a<�!a<M4a<"Ja<�aa<_ya<Z�a<J�a<X�a<��a<�a<��a<�a<%�a<��a<��a<2�a<ܛa<k�a<ȕa<��a<�a<��a<֦a<Ӯa<Ӷa<��a<�a<�a<ÿa<��a<�a<��a<�a<�ma<�Ua<?a<+a<ha<Ra<�a<ra<�a<�(a<3<a<�Ra<:ja<v�a<Z�a<��a<@�a<��a<^�a<��a<��a<��a<��a<��a<�a<�a<C�a<&�a<o�a<|�a<��a<ݥa<��a<<�a<E�a<j�a<�a<иa<�a<x�a<ɍa<xa<A`a<�Ha<]2a<ya<�a<Q	a<�a<�a<�a<5(a<�<a<�Sa<�ja<P�a<˔a<Ǥa<�a<t�a<;�a<��a<�a<8�a<x�a<�a<F�a<4�a<υa<�a<d�a<��a<��a<��a<Ȟa<A�a<̩a<C�a<��a<[�a<J�a<|�a<#pa<�Xa<B@a<B(a<ga<d a<��`<&�`<3�`<��`<y a<$a<X'a<9>a<dUa<�ja<-}a<��a<P�a<G�a<��a<<�a<֐a<�a<j�a<rxa<�qa<�la<�ja<"ka<(na<�sa<zza</�a<�a<��a<��a<��a< �a<Ήa<�|a<Ska<�Va<>?a<t'a<�a<��`<��`<��`<C�`<7�`<��`<��`<�a<D%a<=a<�  �  �La<da<�wa<O�a<�a<�a<��a<��a<��a<܍a<��a<�a<�}a<Y{a<�za<�|a<)�a<��a<�a< �a<N�a<��a<��a<ҝa<��a<��a< }a<ia<�Qa<b9a<� a<�	a<��`<S�`<|�`<��`<��`<��`<�a<Ra<6a<UPa<�ia<ڀa<�a<��a<C�a<b�a<��a<��a<@�a<˦a<{�a<��a<��a<<�a<��a<�a<x�a<Цa<ǭa<�a<
�a<��a<��a<��a<޴a<(�a<�a<��a<~ia<}Pa<�7a<}!a<:a<�a<Y�`<D�`<#a<va<�&a<>a<�Wa<�pa<܈a<֝a<��a<ºa<�a<��a<(�a<j�a<Ӻa<z�a<w�a<Y�a<�a<{�a<@�a<��a<i�a<T�a<��a<�a<��a<�a<��a<׿a<�a<#�a<�a<!}a<8da<�Ja<A2a<a<6a<{a<[�`<� a<t
a<�a<1/a<;Ga<�`a<}ya<��a<�a<%�a<��a<�a<r�a<N�a<��a<c�a<ذa<��a< �a<��a<ܡa<)�a<!�a<�a<Ӱa<�a<��a<��a<��a<'�a<C�a<��a<,�a<��a<�oa<RVa<�<a<%a<a<
a<S�`<|�`<��`<�a<qa< 0a<�Ha<�aa<�ya<��a<i�a<��a<�a<��a<7�a<��a<��a<��a<��a<S�a<��a<��a<��a<�a<ӗa<��a<�a<��a<�a<��a<ϭa<:�a<(�a<!�a<�a<ia<�Oa<�5a<�a<�a<��`<�`<�`<,�`<R�`<��`<�a<Ta<4a<�La<Nda<�xa<�a<��a<K�a<��a<Y�a<�a<�a<.�a<��a<%a<|{a<uya<�ya<A|a<X�a<��a<�a<�a<��a<��a<m�a<�a<��a<ya<�ea<�Na<�5a<@a<�a<��`<��`<
�`<�`<V�`<f�`<��`<�a<�a<�3a<�  �  �Ga<`a<
ua<Ʌa<ёa<,�a<�a<|�a<r�a<��a<��a<�a<h�a<<�a<��a<m�a<��a<^�a<��a<ɘa<ŝa<'�a<ˡa<a<�a<݊a<�ya<�da<�La<�2a<3a<Na<U�`<��`<��`<��`<�`<^�`<��`<�a<)/a<�Ja<ea<(}a<��a<f�a<��a<��a<T�a<m�a<{�a<K�a<٨a<��a<]�a<%�a<�a<��a<Ϩa<H�a<`�a<O�a<�a<��a<r�a<	�a<ܳa<��a<a�a<�|a<�ca<�Ia<�/a<�a<�a<��`<n�`<^�`<a�`<-
a<fa<�6a<�Pa<Nka<s�a<��a<��a<�a<��a<��a<Q�a<��a<x�a<H�a<)�a<ɱa<�a<t�a<(�a<��a<|�a<��a<��a<��a<_�a<��a<X�a<��a<x�a<y�a<�a<(xa<"^a<�Ca<.*a<a<�a<��`<f�`<��`<� a<ya<�&a<@a<cZa<ita<��a<6�a<��a<M�a<K�a<��a<��a<f�a<�a<��a<��a<��a<�a<תa<��a<��a<��a<��a<�a<1�a<��a<��a<�a<��a<Ūa<�a<?�a<Eja<�Oa<^5a<�a<�a<L�`<p�`<��`<�`<S�`<�a<P(a<�Aa<�[a<Gua<�a<�a<��a<2�a<"�a<��a<��a<��a<+�a<�a<��a<P�a<p�a<��a<��a<*�a<�a<��a<�a<�a<c�a<��a<��a<'�a<�a<|a<|da<$Ja<�.a<+a<�`<.�`<9�`<�`<G�`<��`<��`<=�`<�a<�-a<RGa<�_a<pua<�a<ٓa<�a<��a<�a<j�a<��a<��a<d�a<��a<D�a<l�a<��a<ۄa<j�a<.�a<O�a<��a<;�a<6�a<ǘa<��a<��a<eva<�aa<�Ia<�/a<!a<��`<��`<&�`<2�`<�`<u�`<��`<��`<Z�`<�a<G-a<�  �  Fa<�^a<7ta<C�a<��a<X�a<��a<��a<�a<�a<(�a<̌a<U�a<��a<A�a<��a<��a<�a<<�a<��a<Q�a<E�a<K�a<ٞa<��a<I�a<�xa<�ca<�Ja<�0a<�a<_�`<2�`<D�`<��`<��`<��`<(�`<��`<�a<�,a<�Ha<�ca<�{a<ߐa<��a<y�a<W�a</�a<Ƶa<B�a<f�a<9�a<��a<A�a<��a<Z�a<��a<��a<��a<��a<$�a<t�a<��a<��a<�a<i�a<K�a<5�a<�{a<�aa<Ga<B-a<�a<�a<`�`<��`<��`<�`<a<ga<�3a<�Na<�ia<"�a<{�a<�a<��a<��a<n�a<[�a<D�a<Y�a<~�a<Ÿa<��a<��a<��a<~�a<��a<8�a<ջa<��a<��a<��a<E�a<��a<��a<��a<��a<юa<�va<
\a<Aa<`'a<�a<j�`<�`<��`<�`<��`<\a<$$a<~=a<5Xa<�ra<>�a<d�a<�a<��a<w�a<m�a<�a<	�a<q�a<A�a<o�a<~�a<-�a<`�a<�a<��a<c�a<��a<¾a<��a<�a<X�a<0�a<]�a<1�a<�a<��a<�ha<�Ma<�2a<�a<�a<��`<��`<��`<��`<�`<�a<�%a<??a<�Ya<�sa<يa<b�a<�a< �a<��a<ҽa<ٻa<��a<F�a<x�a<[�a<4�a<ؠa<��a<��a<�a<~�a<��a<��a<~�a<L�a<�a<��a<��a<F�a<�za<"ca<EHa<e,a<�a<��`<��`<��`<b�`<��`<?�`<��`<>�`<.a<+a<�Ea<�^a<\ta<b�a<n�a<'�a<"�a<��a<�a<��a<.�a<��a<��a<X�a<�a<�a<Ƈa<%�a<v�a<G�a<��a<��a<�a<��a<Ña<�a<�ua<�`a<bHa<�-a<�a<��`<r�`<��`<��`<V�`<��`<�`<��`<��`<a<+a<�  �  �Ga<`a<
ua<Ʌa<ёa<,�a<�a<|�a<r�a<��a<��a<�a<h�a<<�a<��a<m�a<��a<^�a<��a<ɘa<ŝa<'�a<ˡa<a<�a<݊a<�ya<�da<�La<�2a<3a<Na<U�`<��`<��`<��`<�`<^�`<��`<�a<)/a<�Ja<ea<(}a<��a<f�a<��a<��a<T�a<m�a<{�a<K�a<٨a<��a<]�a<%�a<�a<��a<Ϩa<H�a<`�a<O�a<�a<��a<r�a<	�a<ܳa<��a<a�a<�|a<�ca<�Ia<�/a<�a<�a<��`<n�`<^�`<a�`<-
a<fa<�6a<�Pa<Nka<s�a<��a<��a<�a<��a<��a<Q�a<��a<x�a<H�a<)�a<ɱa<�a<t�a<(�a<��a<|�a<��a<��a<��a<_�a<��a<X�a<��a<x�a<y�a<�a<(xa<"^a<�Ca<.*a<a<�a<��`<f�`<��`<� a<ya<�&a<@a<cZa<ita<��a<6�a<��a<M�a<K�a<��a<��a<f�a<�a<��a<��a<��a<�a<תa<��a<��a<��a<��a<�a<1�a<��a<��a<�a<��a<Ūa<�a<?�a<Eja<�Oa<^5a<�a<�a<L�`<p�`<��`<�`<S�`<�a<P(a<�Aa<�[a<Gua<�a<�a<��a<2�a<"�a<��a<��a<��a<+�a<�a<��a<P�a<p�a<��a<��a<*�a<�a<��a<�a<�a<c�a<��a<��a<'�a<�a<|a<|da<$Ja<�.a<+a<�`<.�`<9�`<�`<G�`<��`<��`<=�`<�a<�-a<RGa<�_a<pua<�a<ٓa<�a<��a<�a<j�a<��a<��a<d�a<��a<D�a<l�a<��a<ۄa<j�a<.�a<O�a<��a<;�a<6�a<ǘa<��a<��a<eva<�aa<�Ia<�/a<!a<��`<��`<&�`<2�`<�`<u�`<��`<��`<Z�`<�a<G-a<�  �  �La<da<�wa<O�a<�a<�a<��a<��a<��a<܍a<��a<�a<�}a<Y{a<�za<�|a<)�a<��a<�a< �a<N�a<��a<��a<ҝa<��a<��a< }a<ia<�Qa<b9a<� a<�	a<��`<S�`<|�`<��`<��`<��`<�a<Ra<6a<UPa<�ia<ڀa<�a<��a<C�a<b�a<��a<��a<@�a<˦a<{�a<��a<��a<<�a<��a<�a<x�a<Цa<ǭa<�a<
�a<��a<��a<��a<޴a<(�a<�a<��a<~ia<}Pa<�7a<}!a<:a<�a<Y�`<D�`<#a<va<�&a<>a<�Wa<�pa<܈a<֝a<��a<ºa<�a<��a<(�a<j�a<Ӻa<z�a<w�a<Y�a<�a<{�a<@�a<��a<i�a<T�a<��a<�a<��a<�a<��a<׿a<�a<#�a<�a<!}a<8da<�Ja<A2a<a<6a<{a<[�`<� a<t
a<�a<1/a<;Ga<�`a<}ya<��a<�a<%�a<��a<�a<r�a<N�a<��a<c�a<ذa<��a< �a<��a<ܡa<)�a<!�a<�a<Ӱa<�a<��a<��a<��a<'�a<C�a<��a<,�a<��a<�oa<RVa<�<a<%a<a<
a<S�`<|�`<��`<�a<qa< 0a<�Ha<�aa<�ya<��a<i�a<��a<�a<��a<7�a<��a<��a<��a<��a<S�a<��a<��a<��a<�a<ӗa<��a<�a<��a<�a<��a<ϭa<:�a<(�a<!�a<�a<ia<�Oa<�5a<�a<�a<��`<�`<�`<,�`<R�`<��`<�a<Ta<4a<�La<Nda<�xa<�a<��a<K�a<��a<Y�a<�a<�a<.�a<��a<%a<|{a<uya<�ya<A|a<X�a<��a<�a<�a<��a<��a<m�a<�a<��a<ya<�ea<�Na<�5a<@a<�a<��`<��`<
�`<�`<V�`<f�`<��`<�a<�a<�3a<�  �  �Ta<�ia<�{a<i�a<(�a<A�a<�a<*�a<ˋa<)�a<w|a<ua<�oa<�la<la<�ma<�ra<3ya<&�a<��a<֑a<��a<d�a<��a<4�a<3�a<M�a<Zoa<PZa<RCa<j,a<�a<�a<��`<y�`<��`<��`<�a<Ka<�(a<�@a<|Ya<qa<�a<A�a<�a<ʫa<�a<�a<��a<��a<��a<��a<��a<@�a<��a<A�a<f�a<H�a<ۚa<f�a<6�a<9�a<D�a<2�a<�a<�a<S�a<Ǜa<��a<~ra<�Za<Da<%/a<a<Aa<{a<La<�a<�!a<M4a<"Ja<�aa<_ya<Z�a<J�a<X�a<��a<�a<��a<�a<%�a<��a<��a<2�a<ܛa<k�a<ȕa<��a<�a<��a<֦a<Ӯa<Ӷa<��a<�a<�a<ÿa<��a<�a<��a<�a<�ma<�Ua<?a<+a<ha<Ra<�a<ra<�a<�(a<3<a<�Ra<:ja<v�a<Z�a<��a<@�a<��a<^�a<��a<��a<��a<��a<��a<�a<�a<C�a<&�a<o�a<|�a<��a<ݥa<��a<<�a<E�a<j�a<�a<иa<�a<x�a<ɍa<xa<A`a<�Ha<]2a<ya<�a<Q	a<�a<�a<�a<5(a<�<a<�Sa<�ja<P�a<˔a<Ǥa<�a<t�a<;�a<��a<�a<8�a<x�a<�a<F�a<4�a<υa<�a<d�a<��a<��a<��a<Ȟa<A�a<̩a<C�a<��a<[�a<J�a<|�a<#pa<�Xa<B@a<B(a<ga<d a<��`<&�`<3�`<��`<y a<$a<X'a<9>a<dUa<�ja<-}a<��a<P�a<G�a<��a<<�a<֐a<�a<j�a<rxa<�qa<�la<�ja<"ka<(na<�sa<zza</�a<�a<��a<��a<��a< �a<Ήa<�|a<Ska<�Va<>?a<t'a<�a<��`<��`<��`<C�`<7�`<��`<��`<�a<D%a<=a<�  �  �^a<Hqa<�a<܋a<��a<y�a<��a<?�a<_�a<jwa<Qma<zda<�]a<�Ya<�Xa<[a<�`a<�ha<�ra<n}a< �a<*�a<{�a<a�a<��a<H�a<�a<Uwa<�da<Pa<t;a<(a<�a<�a<�a<Ta<�	a<a<%a<�8a<�Na<�da<:za<��a<��a<��a<êa<S�a<ۧa<=�a<��a<�a<Ņa<H~a<�xa<Kva< wa<�za<ˁa<��a<��a<��a<>�a<��a<)�a<��a<^�a<Q�a<>�a<x�a<�}a<�ha<�Sa<�@a<51a<=&a<	!a<�!a<�(a<�4a<�Ea<mYa<�na<�a<��a<0�a<��a<2�a<�a<N�a<�a<��a<��a<Y�a<��a<�a<��a<��a<f�a<��a<~�a<o�a<ԡa<!�a<��a<d�a<��a<H�a<�a<��a<��a<��a<�ya<?da<�Oa<K=a<�.a<�%a<3"a<�$a<f-a<;a<�La<6aa<�va<a�a<̝a<�a<��a<v�a<��a<;�a<��a<N�a<�a<a�a<�a<�a<5�a<�a<��a<��a<؍a<;�a<z�a<a�a<ݳa<}�a<��a<7�a<)�a<�a<a<u�a<ma<�Wa<wCa<+2a<O%a<�a<Ca<� a<+a<:a<�La<Eaa<qva<m�a<��a<�a<��a<n�a<��a<��a<S�a<�a<��a<�a<�}a<�va<�ra<�qa<�sa<&ya<{�a<��a<Q�a<E�a<D�a<9�a<A�a<��a<G�a<�a<�xa<da<�Ma<8a<$a<�a<�a<�a<�a<�a<Qa<n#a<�6a<>Ka<`a<sa<�a<�a<��a<\�a<�a<�a<I�a<�|a<ra<�ga<�_a<Za<�Wa<Xa<�[a<rba<ka<2ua<<a<]�a<�a<m�a<��a<��a<��a<�ra<0`a<DKa<�5a<
!a<�a<o a<�`<��`<��`<P�`<,a<4a<�3a<_Ia<�  �  �ia<�ya<��a<	�a<~�a<ԏa<�a<��a<�ta<�ga<�[a<uPa<Ha<Ca<�Aa<�Da<CKa<Ua<8aa<�na<#|a< �a<��a<k�a<Øa<��a<��a<I�a<ipa<�^a<lLa<p;a<-a<r"a<�a<a<!a<)+a<k9a<�Ja<g^a<�qa<6�a<��a<��a<�a<C�a<��a<E�a<��a<�a<�~a<Gsa<�ia<�ba<�_a<4`a<�da<�la<xa<�a<˒a<^�a<Ϋa<4�a<��a<n�a<��a<?�a<1�a<h�a<xa<�ea<�Ta<-Ga<�=a<�8a<�9a<�?a<oJa<2Ya<�ja<�}a<�a<Ѡa<f�a<��a<��a<{�a<��a<0�a<�a<�a<=�a<o~a<�ta<gna<�ka<�la<�qa<2za<b�a<�a<;�a<}�a<x�a<�a<y�a<ٻa<s�a<̨a<6�a<��a<�ta<.ba<Ra<eEa<'=a<�9a<m<a<�Ca<Pa<�_a<�qa<��a<c�a<*�a<&�a<�a<��a<�a<��a<�a<��a<k�a<��a<ya<7pa<�ja<�ha<5ka<+qa<\za<�a<��a<�a<Ϊa<��a<��a<X�a<ܴa<�a<��a<�a<�{a<�ha<�Va<�Ga<,<a<|5a<4a<8a<%Aa<ZNa<�^a<qa<x�a<l�a<ݢa<�a<�a<�a<߯a<�a<��a<i�a<��a<�ta<!ia<�`a<�[a<�Za<�]a<2da<�ma<%ya<\�a<d�a<T�a<C�a<e�a<��a<�a<�a<��a<�pa<[]a<�Ia<8a<�)a<�a<ua<ta<�a<�(a<7a<�Ga<PZa<la<G|a<M�a<�a<w�a<Õa<s�a<l�a<�{a<Nna<�`a<�Ta<�Ja<�Ca<�@a<oAa<!Fa<)Na<Ya<fea<Wra<[~a<�a<o�a<��a<�a<W�a<�za<�ja<	Ya<�Ea<�3a<{#a<�a<�a<�a<(a<�a<'"a<	2a<IDa<}Wa<�  �  �ta<��a<��a<
�a<�a<1�a<E�a<lua<�fa<�Va<Ha<�:a<z0a<�*a<)a<a,a<�3a<�?a<2Na<6^a<�na<�}a<��a<m�a<&�a<��a<u�a<5�a<[|a<�ma<a^a<Pa<�Ca<j:a<�5a<;5a<�9a<RBa<Oa<(^a<�na<ma<t�a<#�a<��a<§a<��a<�a<j�a<|�a<�{a<�la<_a<Sa<�Ja<�Fa<sGa<�La<$Va<{ca<�ra<��a<ݓa<��a<S�a<̵a<�a<��a<�a<�a<z�a<�a<�xa<Rja<,^a<�Ua<�Qa<�Ra<�Wa<aa<$na<�|a<�a<Z�a<�a<s�a<��a<g�a<θa< �a<&�a<�a<�a<xwa<\ia<�]a<!Va<�Ra<6Ta<
Za<%da<�qa<��a<��a<�a<g�a<�a<��a<|�a<�a<��a<"�a<��a<��a<va<ha<�\a<�Ua<(Sa<MUa<�[a<@fa<�sa<�a<�a<��a<j�a<-�a<�a<��a<M�a<��a<��a<��a<m�a<qa<;ca<�Xa<2Ra<Pa<�Ra<�Ya<ea<�ra<6�a<�a<e�a<��a<��a<��a<��a<��a<��a<�a<֊a<�za<}ka<^a<%Ta<tNa<.Ma<�Pa<PXa<da< ra<h�a<�a<��a<�a<�a<�a<Y�a<P�a<�a<��a<�a<�oa<G`a<�Ra<�Ha<)Ca<Ba<�Ea<~Ma<7Ya<�fa<va<�a<�a<a�a<n�a<3�a<��a<��a<��a<�}a<Uma<�\a<�Ma<}@a<r7a<�2a<w2a<�6a<�?a<�Ka<"Za<�ia<bxa<��a<\�a<�a<;�a<�a<�a<f}a<�na<P^a<>Na<�?a<�3a<�+a<�'a<�(a<Z.a< 8a<KEa<Ta<da<�ra<	�a<|�a<�a<��a<��a<q�a<�ua<ga<�Va<mGa<|9a<P.a<h'a<�$a<'a<|-a<Q8a<-Fa<�Ua<�ea<�  �  �a<Z�a<r�a<@�a<�a<��a<�ya<ja<GXa<{Ea<�3a<m$a<�a<�a<�a<�a<�a<�)a<�:a<fMa<�`a<�ra<��a<�a<��a<��a<��a<z�a<�a<U|a<�oa<�ca<�Ya<BRa<3Na<Na<�Qa<YYa<�ca<�pa<�~a<a�a<K�a<��a<�a<ϧa<~�a<ߚa<��a<�}a<{la<[Za<�Ia<N<a<�2a<�-a<[.a<V4a<??a<*Na<`a<�sa<�a<ɘa<��a<L�a<��a<ɹa<�a<��a<'�a<��a<ߊa<�~a<�ta<$na<�ja<Bka<�oa<zwa<F�a<��a<Λa<U�a<��a<۹a<�a<V�a<��a<��a<��a<T�a<�va<da<�Sa<hFa<w=a<�9a<B;a<#Ba<�Ma<]a<�na<�a<:�a<��a<��a</�a<N�a<G�a<ҷa<��a<$�a<�a<3�a<�}a<Tta<Tna<la<�ma<5sa<�{a<G�a<�a<�a<��a<�a<��a<�a<f�a<�a<��a<R�a<,�a<�na<�\a<�La<�@a<J9a<�6a<:a<eBa<Oa<%_a<_qa<(�a<��a<�a<3�a<C�a<�a<��a<�a<��a<A�a<�a<_a<=ta<�ka<ga<�ea<�ha<Zoa<�xa<��a<9�a<ߝa<��a<p�a<��a<��a</�a<�a<��a<�a<�pa<@]a<2Ka<�;a<�0a< *a<�(a<S-a<�6a<�Ca<,Ta<Bfa<xa<L�a<a<�a<�a<��a<ʞa<�a<x�a<�|a<oa<4ba<LWa<�Oa<YKa<"Ka<�Na<�Ua<`a<�ka<lxa<_�a<6�a<Ɣa<w�a<-�a<�a<��a<�ra<aa<�Ma<�:a<�)a<Ka<�a<�a<�a<wa<�!a<�0a<MBa<-Ua<ga<Iwa<�a<f�a<V�a<$�a<��a<T�a<�ta<rga<�Za<�Na<�Ea<�?a<�=a<q?a<Ea<�Ma<�Ya<lfa<�sa<�  �  D�a<��a<�a<��a<��a<a<Yqa<�^a<Ja<�4a<� a<Xa<$a<�`< �`<#�`<8a<.a<(a<G=a<CSa<�ha<{a<n�a<�a<��a<��a<��a<-�a<g�a<�a<%va<na<ha<�da<�da<ha<�na<wa<��a<��a<��a<Πa<��a<k�a<0�a<X�a<t�a<��a<�qa<C]a<Ia<86a<�&a<�a<a<�a<"a<^)a<5:a<mNa<;da<�za<2�a<�a<֮a<��a<ֻa<?�a<��a</�a<��a<��a<ڑa<
�a<:�a<��a<��a<��a<"�a<��a<�a<:�a<ɲa<(�a<S�a<f�a<ιa<w�a<5�a<��a<|a<�fa<�Qa<&?a<80a<&a<�!a<�#a<W+a<g8a<�Ia<^a<psa<��a<כa<�a<��a<S�a<o�a<�a<��a<1�a<�a<��a<,�a<̉a<��a<��a<;�a<Ԉa<׏a<��a<;�a<H�a<&�a<M�a<!�a<n�a<�a<ܫa<�a<(�a<�sa<O^a<�Ia<�7a<,*a<�!a<a<�"a<,a<g:a<�La<;aa<�va<!�a<�a<��a<r�a<x�a<׺a<��a<ׯa<S�a<��a<��a<��a<΁a<�}a<�|a<a<��a<�a<��a<��a<8�a<�a<�a<��a<W�a<�a<��a<G�a<�wa<�aa<�Ka<{7a<8&a<�a<ca<>a<a<� a<�/a<�Ba<�Va<�ka<�~a<�a<u�a<��a<ĥa<�a<1�a<~�a<�a<�a<ua<Vla<�ea<.ba<�aa<�da<�ja<{ra<|a<؅a<Ԏa<��a<A�a<ɘa<��a<ɉa<{a<�ha<�Sa<�=a<�(a<�a<a<}�`<��`<@�`<��`<ia<�a<s1a<�Fa<�[a<zna<U~a<ԉa<Y�a<I�a<��a<��a<��a<{va<la<�ba<+[a<#Va<�Ta<�Ua<�Za<�aa<;ka<�ua<�a<�  �  �a<�a<��a<��a<�a<�{a<�ia<�Ta<�=a<4&a<a<��`<s�`<��`<��`<��`<��`<a<�a<"/a<]Ga<_a<ta<��a<�a<E�a<��a<c�a<��a<;�a<�a<��a<Ia<bza<�wa<.xa<�za<6�a<��a<�a<Әa< �a<ȧa<o�a</�a<]�a<Ҝa<i�a<7|a<ga<Pa<�9a<�$a<�a<�a<�a<a<1	a<Ka<�(a<�>a<�Va<loa<��a<��a<�a<��a<O�a<p�a<l�a<P�a<O�a<��a<�a<��a<זa<єa<*�a<�a<u�a<m�a<L�a<Q�a<f�a<A�a<��a<H�a<�a<�a<\�a<M�a<upa<�Xa<�Aa<7-a<�a<�a<=a<a<�a<�%a<�8a< Oa<�fa<n~a<��a<n�a<��a<�a<��a<��a<|�a<2�a<y�a<n�a<��a<ța<��a<B�a<A�a<�a<͠a<�a<�a<��a<�a<��a<��a<u�a<~�a<��a<y�a<a<}ga<�Oa<9a<d%a<va<@a<�
a<]a<�a<F(a<N<a<Sa<�ja<��a<�a<�a<m�a<�a<�a<Ƽa<+�a<&�a<�a<
�a<ݙa<!�a<ڐa<'�a<Αa<;�a<y�a<Уa<��a<��a<�a<^�a<��a<��a<��a<��a<�a<ma<�Ta<�<a<&a<Na<�a<��`<��`<-a<�a<fa<�2a<gIa<n`a<va<��a<��a<١a<;�a<�a<ߤa<��a<��a<��a<G�a<�}a<Exa<pua<ua<)wa<�{a<A�a<��a<�a<q�a<��a<Ҝa<��a<�a<\�a<,ta<�_a<AHa<0a<�a<�a<��`<l�`<V�`<��`<��`<��`<�a<�"a<�9a<OQa<�fa<�xa<�a<�a<��a<��a<�a<��a<܂a<�za<Ksa<"ma<ia<�ga<�ha<�la<�ra<Aza<c�a<`�a<�  �  ��a<��a<%�a<a�a<Ɇa<xwa<�ca<�La<�3a<�a<�a<��`<%�`<��`<U�`<+�`<��`<!�`<�
a<$a<�=a<[Wa<�na<�a<)�a<q�a<��a<}�a<��a<q�a<ݖa<?�a<�a<��a<��a<݆a<o�a<��a<��a<��a<ءa<F�a<ͬa<V�a<�a<|�a<��a<߉a<�ua<E^a<�Ea<{-a<ea<a<�`<��`<��`<~�`<�a<a<u2a<tLa<�fa<�a<ޕa<��a<��a<�a<�a<?�a<@�a<"�a<�a<�a<ڨa<j�a<��a<�a<^�a<r�a<.�a<i�a<��a<��a<��a<�a<��a<��a<��a</�a<�a<8ga<�Ma<5a<da<�a<!a<��`<%�`<%a<xa<�+a<hCa<�\a<va<�a<3�a<>�a<��a<&�a<_�a<��a<��a<�a<y�a<n�a<��a<c�a<��a<��a<ͨa<d�a<9�a<~�a<a�a<��a<G�a<]�a<=�a<E�a<��a<��a<wa<�]a<Da<�+a<4a<%a<U�`<G�`<��`<g	a<Qa<�/a<�Ga<@aa<�ya<��a<I�a<��a<@�a<�a<��a<S�a<[�a<�a<��a<��a<Q�a<��a<מa<u�a<��a<��a<|�a<��a<ʹa<�a<G�a<��a<��a<��a<�a<E}a<cda<oJa<b0a<�a<�a<�`<��`<��`<{�`<��`<�a<�&a< ?a<�Wa<oa<�a<��a<��a<��a<ªa<��a<��a<U�a<3�a<P�a<#�a<׆a<"�a<��a<��a<�a<�a<��a<Y�a<�a<�a<	�a<�a<k�a<�a<oa<*Xa<?a<5%a<�a<��`<��`<��`<�`<��`<��`<��`<T�`<�a<0a<�Ha<�`a<�ta<r�a<��a<��a<�a<}�a<=�a<G�a<ͅa<�a<�za<�wa<uva<�wa<�za<ca<t�a<��a<+�a<�  �  1�a<��a<L�a<�a<3�a<�ta<�_a<�Ga<�-a<ra<��`<��`<y�`<��`<b�`<W�`<�`<2�`<�a<�a<�7a<vRa<�ja<�a<Џa<q�a<e�a<�a<^�a<r�a<.�a<��a<9�a<1�a<��a<ӏa<7�a<�a<T�a<Z�a<k�a<��a<�a<B�a<Ҭa<��a<��a<��a<!qa<�Xa<B?a<�%a<�a<��`<H�`<��`<�`<��`<0�`<la<�*a<�Ea<�`a<{a<b�a<ۥa<��a<��a<��a<4�a<X�a<��a<��a<��a<;�a<,�a<w�a<ˬa<�a<��a<��a<ۼa<��a<��a<I�a<��a<ӿa<T�a<!�a<i�a<{a<Saa<�Fa<5-a<�a<Ta<P�`<�`<A�`<k�`<Ia<@#a<<a<�Va<�pa<��a<-�a<��a</�a<*�a<��a<J�a<U�a<��a<r�a<E�a<��a<;�a<�a<ܮa<X�a<Q�a<M�a<��a<�a<�a<��a<��a<�a<��a<��a<u�a<�qa<�Wa<�<a<�#a<a<x�`<o�`<Q�`<��`<��`<`a<�'a<�@a<<[a<	ua<��a<��a<R�a<?�a<}�a<s�a<�a<\�a<V�a<�a<ήa<�a<z�a<ͧa<>�a<�a<O�a<;�a<%�a<
�a<%�a<3�a<f�a<�a<��a<��a<�xa<�^a<�Ca<�(a<a<g�`<>�`<��`<��`<��`<��`<%a<�a<98a<�Qa<�ja<j�a<v�a<Пa<��a<��a<��a<��a<Ȥa<ٞa<ؘa<��a<��a<�a<��a<-�a<�a<S�a<�a<��a<��a<Ƣa<��a<;�a<4�a<za<>ka<fSa<$9a<4a<a<��`<E�`<��`<+�`<��`<��`<R�`<��`<|a<�)a<�Ca<D\a<�qa<��a<0�a<��a<9�a<ՙa<Ɩa<%�a<Ìa<��a<S�a<��a<na<z�a<!�a<N�a<��a<�a<זa<�  �  P�a<9�a<ߋa<�a<�|a<�oa<�_a<�Ma<�9a<8&a<�a<a<#�`<��`<��`<��`<��`<�	a<�a<C.a<�Ba<#Wa<�ia<�ya<��a<�a<��a<U�a<��a<��a<��a<C�a<P�a<��a<&�a<��a<*�a<p�a<��a<4�a<�a<۠a<F�a<�a<P�a<��a<J�a<��a<�ra<i`a<Ma<I:a<.)a<a<Pa<a<�a<�a<�a<,-a<�?a<�Sa<�ha<�|a<��a<��a<��a<��a<��a<Ƿa<ٶa<(�a<��a<��a<Ʃa<C�a<~�a<��a<�a<"�a<��a<��a<p�a<D�a<�a<7�a<t�a<2�a<b�a<�a<l~a<�ja<�Va<�Ca<�2a<%a<a<�a<�a<� a<�,a<H<a<�Na<�ba<�va<��a< �a<ϧa<��a<�a<�a<��a<w�a<�a<$�a<N�a<�a<ݨa<F�a<��a<s�a<��a<)�a< �a<U�a<�a<�a<g�a<5�a<��a<>�a<�a<Twa<ca<�Na<<a<�+a<}a<�a<"a<�a<
!a<(.a<�>a<�Qa<xea<$ya<�a<l�a<��a<(�a<;�a<#�a<��a<ܲa<�a<�a<C�a<�a<`�a<��a<��a<ͤa<اa<n�a<�a<��a<�a<o�a<]�a<��a<��a<��a< za<<fa<YQa<=a<T*a<�a<Fa<ya<Ya<a<[a<3#a<4a<�Fa<EZa<�la<)}a<1�a<h�a</�a<\�a<��a<�a<&�a<��a<��a<܌a<}�a<�a<\�a<�a<Y�a<K�a<��a<��a<��a<*�a<ϓa<��a<��a<]ya<|ia<aWa<GCa<�.a<a<�	a<��`<@�`<��`<�`<��`<Ka<�a<�"a<�6a<�Ja<�\a<Ama<�za<f�a<��a<s�a<ߍa<��a<F�a<B�a<i�a<*}a<{a<�za<{a<}a<P�a<'�a<>�a<ًa<�  �  .�a<��a<��a<�a<}a<vpa<�`a<�Na<~;a<(a<�a<aa<e�`<��`<��`<��`<�`<�a<�a<0a<MDa<7Xa<�ja<Oza<�a<�a<j�a<��a<\�a<.�a< �a<v�a<+�a<Èa<��a<�a<�a<9�a<��a<��a<��a<��a<]�a<��a<4�a<�a<��a<��a<�sa<�aa<�Na<<a<g+a<ha<�a<a<�a<Xa< a<f/a<oAa<�Ua<ja<�}a<l�a<H�a<��a<��a<��a<�a<��a<ɲa<	�a<�a<��a<�a<£a<�a<�a<�a<�a<%�a<�a<�a<H�a<�a<x�a<i�a<ןa<��a<~a<Ela<�Xa<�Ea<�4a<H'a<�a<�a<�a<#a<�.a<t>a<�Pa<pda< xa<��a<ؚa<�a<��a<ڷa<��a<w�a<(�a<��a<v�a<\�a<רa<u�a<��a<(�a<?�a<��a<q�a<��a<��a<]�a<��a<�a<;�a<�a<�a<�a<sxa<�da<�Pa<4>a<:.a<�!a<�a<3a<Ra<I#a<l0a<�@a<eSa<�fa<8za<ދa<��a<צa<)�a<�a<z�a<n�a<��a<��a<9�a<�a<ݡa<̟a<;�a<@�a<��a<��a<ީa<��a<��a<�a<�a<A�a<ǥa<ښa<U�a<�za<xga<Sa<�>a<�,a<�a<�a<ta<]
a<�a<�a<m%a<�5a<�Ha<�[a<�ma<~a<��a<��a<!�a<�a<"�a<��a<Ƙa<�a<�a<��a<=�a<+�a<��a<υa<!�a<q�a<�a<d�a<��a<o�a<��a<��a<�a<�ya<rja<rXa<�Da<�0a<a<�a<��`<��`<��`<��`< �`<�a<�a<�$a<H8a<�Ka<�]a<�ma<{a<t�a<n�a<��a<Ɍa<a�a<Άa<��a<x~a<�za<�xa<�wa<�xa<�za<K~a<p�a<��a<��a<�  �  f�a<�a<��a<�a<~a<lra<�ca<�Ra<%@a<j-a<�a<3a<�a<��`<��`<��`<Ka<�a<�"a<J5a<�Ha<�[a<Rma<	|a<��a<��a</�a<��a<i�a<j�a<8�a<�a<��a<S�a<�a<?�a<{�a<�a<֋a<o�a<@�a<Y�a<��a<�a<��a<�a<ԑa<څa<�va<�ea<�Sa<�Aa<�1a<k$a<�a</a<�a<ya<1'a<�5a<Ga<�Za<.na<�a<�a<��a<#�a<�a<4�a<��a<i�a<��a<��a<U�a<;�a<��a<�a<e�a<{�a<��a<<�a<E�a<0�a<��a<�a<��a<$�a< �a<x�a<��a<��a<�pa<�]a<_Ka<�;a<l.a<�%a<�!a<�#a<9*a<�5a<�Da<Va<.ia<�{a<��a<�a<1�a<�a<��a<иa<ȷa<��a<*�a<�a<[�a<r�a<��a<՞a<��a<աa<q�a< �a<�a<p�a<��a<Ʒa<�a<K�a<�a<ܜa<ލa<1|a<]ia<2Va<LDa<5a<�(a<�!a<Oa<x"a<x*a<7a<�Fa<�Xa<hka<�}a<��a<��a<��a<�a<��a<t�a<|�a<��a<Ũa<��a<�a<n�a<+�a<��a<֙a<>�a<'�a<��a<V�a<>�a<��a<~�a<��a<,�a<�a<��a<,~a<}ka<
Xa<fDa<�2a<�#a<�a<�a<wa<�a<�a<�+a<�;a<�Ma<�_a<qa<��a<�a<
�a<��a<��a<��a<{�a<��a<�a<W�a<R�a<ـa<z~a<	~a<da<�a<ʅa<1�a<��a<��a<D�a<5�a<.�a<��a<r{a<%ma<�[a<	Ia<�5a<�"a<�a<a<��`<��`<�`<H�`<}
a<a<<*a<=a<�Oa<aa<pa<|a<��a<��a<@�a<�a<�a<S�a<5}a<yxa<�ta<(ra<!qa<ra<kta<8xa< }a</�a<��a<�  �  ݅a<�a<K�a<3�a<�a<`ua<-ha<�Xa<SGa<�5a<�%a<�a<a<�a<a<�a<�a<�a<	,a<�=a<�Oa<�aa<Gqa<�~a<�a<}�a<��a<S�a<��a<�a<��a<&�a<J{a<�wa<�ua<5va<xxa<�|a<��a<^�a<p�a<Жa<�a<��a<��a<�a<�a<7�a<�{a<&la<G[a<�Ja<;a<#/a<}&a<)"a<�"a</(a<2a<�?a<TPa<Uba<�ta<9�a<d�a<�a<תa<7�a<��a<��a<�a<�a<��a<+�a<@�a<��a<�a<g�a<��a<�a<\�a<��a<ƪa<��a<��a<δa<Ʋa<)�a<
�a<w�a<��a<dwa<�ea<�Ta<�Ea<�9a<�1a< .a<|/a<�5a<?@a<@Na<�^a<{pa<'�a<J�a< �a<ߪa<�a<ӵa<�a<p�a<ծa<�a<Ţa<�a<�a<�a<ɓa<��a<[�a<�a<��a<��a<l�a<	�a<ȴa<Ҵa<a�a<c�a<Пa<9�a<>�a<�pa<�^a<�Ma<f?a<k4a<�-a<^+a<D.a<�5a<9Aa<Pa<�`a<Yra<��a<��a<d�a<٨a<��a<�a<$�a<��a<r�a<D�a<�a<<�a<��a<(�a<��a<юa<%�a<�a<��a<��a<��a<��a<�a<��a<��a</�a<�a<)�a<�qa<�_a<�Ma<�<a<�.a<s$a<�a<ya<[!a<�)a<�5a<�Da<NUa<Afa<Ava<�a<*�a<��a<՚a<`�a<�a<$�a<�a<�a<.�a<Xza<�ua<ysa<sa<�ta<xa<�|a<��a<�a<��a<ɏa<d�a<ύa<��a<~a<�pa<uaa<�Oa<�=a<C,a<�a<)a<�a<�a<�a<�
a<�a<�"a<3a<RDa<�Ua<�ea<"sa<�}a<ބa<j�a<v�a<ąa<�a<;{a<�ta<oa<?ja<$ga<fa<ga<�ia<�na<�ta<�za<�a<�  �  �a<��a<�a<�a<]�a<Iya<�ma<`a<�Pa<�@a<2a<-%a<ka<�a<Xa<Ka<�a<*a<J8a<Ha<�Xa<�ha<}va<1�a<'�a<Ďa<��a<��a<�a<��a<�{a<`ta<bna<�ia<�ga<�ga<~ja<�oa<8va<�~a<E�a<f�a<j�a</�a<�a<^�a<l�a<��a<��a<9ta<ea<LVa<pHa<=a<
5a<F1a<�1a<�6a<@a<�La<\a<Qla<}a<��a<
�a<��a<c�a<�a<��a<m�a<إa<��a<Z�a<�a<�a<��a<��a<)�a<�a<�a<p�a<Q�a</�a<?�a<̮a<�a<رa</�a<?�a<�a<Z�a<�a<1pa<�`a<�Ra<�Ga<F@a<E=a<�>a<?Da<Na<�Za<ja<�ya<ˉa<
�a<�a<�a<��a<ʳa<�a<��a<�a<|�a<��a<H�a<��a<ֆa<t�a<k�a<�a<.�a<$�a<�a<i�a<��a<��a<��a<�a<-�a<��a<͗a<��a<�ya<�ia<qZa<Ma<�Ba<w<a<�:a<=a<Da<�Na<G\a<nka<4{a<��a<ؗa<ܢa< �a<�a<l�a<��a<�a<�a<,�a<#�a<S�a<�a<�a<2a<׀a<�a<��a<őa<W�a<H�a<�a<��a<$�a<	�a<��a<}�a<Q�a<
za<Tia<Ya<�Ia<�<a< 3a<�-a<�,a<�/a<�7a<�Ba<�Pa<J_a<�na<�|a<��a<��a<L�a<��a<�a<��a<�a<��a<V|a<�sa<7ma<�ga<,ea<�da<�fa<'ka<�pa<=xa<~a<��a<��a<��a<��a<��a<5�a<�ua<Hha<�Xa<"Ha<V8a<�)a<aa<pa<
a<�a<Ja<�"a<_/a<">a<�Ma<a]a<cka<=wa<�a<��a<c�a<u�a<�a<Cya<�qa<�ia<lba<�\a<Ya<�Wa<�Xa<}\a<�aa<*ia<5qa<�xa<�  �  �xa<�a<�a<o�a<�a<#}a<ta<Vha<?[a<MMa<,@a<�4a<G,a<'a<�%a<�(a<�/a<{9a<�Ea<'Ta<�ba<Qpa<U|a<u�a<d�a<��a<j�a<+�a<6�a<�xa<�oa<�fa<+_a<�Ya<�Va<�Va<�Ya<�_a<�ga<�qa<5|a<��a<ݏa<֖a<�a<��a<��a<x�a<�a<I}a<zpa< ca<)Wa<HMa<'Fa<�Ba<\Ca<�Ga<iPa<�[a<ia<�wa<f�a<��a<�a<"�a<��a<��a<��a< �a<O�a<�a<��a<΁a<Vza<Cua<�ra<sa<�va<�|a<��a<�a<�a<2�a<	�a<6�a<��a<<�a<@�a<"�a<�a<�a< |a<Lna<#ba<aXa<�Qa<�Na<Pa<1Ua<�]a<Bia<�va<لa<Z�a<��a<E�a<��a<ѱa<�a<?�a<��a<��a<��a<c�a<��a<�za<va<Gta<�ua<�ya<X�a<Ԉa<<�a<�a<��a<��a<��a<��a<խa<��a<�a<��a<|�a<va<�ha<�\a<�Sa<�Ma<-La<~Na<�Ta<^a<�ia<�wa<m�a<^�a<��a<#�a<`�a<��a<��a<��a<L�a<�a<�a<��a<ya<�ra<�na<na<Hpa<ua<1|a<�a<E�a<��a<��a<2�a<��a<a�a<�a<F�a<;�a<�a<�ta<�ea<NXa<�La<Da< ?a< >a<+Aa<Ha<�Qa<�]a<�ja<�wa<Ãa<��a<`�a<�a<��a<�a<W�a<e�a<!za<�oa<�ea<r]a<�Wa<Ta<�Sa<�Va<�[a<=ca<�ka<0ua<�}a<,�a<ɉa<��a<��a<3�a<�{a<�oa<rba<Ta<�Ea<$9a<�.a<�'a<�$a<b%a<8*a<�2a<�=a<�Ja<�Xa<�ea<�qa<h{a<��a<��a<��a<�a<�xa<pa<0fa<�\a<�Sa<�La<SHa<�Fa<Ha<`La<)Sa<�[a<�ea<toa<�  �  pa<�ya<��a<��a<��a<��a<}za<�pa<)fa<fZa<IOa<pEa<�=a<�9a<v8a<;a<�@a<�Ia<�Ta<�`a<!ma<pxa<8�a<��a<��a<:�a<��a<فa<Pxa<�ma<Yba<�Wa<�Na<Ha<�Da<eDa<�Ga<�Na<?Xa<�ca<Tpa<�|a<T�a<�a<:�a<��a<�a<.�a<)�a<��a< |a<�pa<�fa<^a<?Xa<kUa<Va<*Za<Maa<~ka<wa<̃a<�a<5�a<�a<��a<L�a<��a<�a<�a<��a<z�a<�|a<Sra<Gia<Mca<O`a<�`a<�da<�ka<�ua<��a<��a<�a<i�a<"�a<��a<�a<N�a<��a<۞a<:�a<��a<�|a<Nra<�ia<�ca<paa<�ba<
ga<�na<�xa<�a<�a<-�a<F�a<k�a<��a<7�a<�a<��a<V�a<|�a<��a<�{a<�qa<.ia<�ca<�aa<nca<3ha<pa<5za<��a<l�a<<�a<ǥa<)�a<��a<j�a<m�a<��a<��a<h�a<7�a<�wa<Wma<\ea<{`a<�^a<�`a<fa<`na<�xa<,�a<ݏa<��a<��a<q�a<~�a<��a<�a<��a<g�a<�a<�}a<�ra<�ha<"aa<�\a<�[a<C^a<�ca<�la<�va<b�a<��a<��a<J�a<@�a<f�a<D�a<��a<z�a<t�a<e�a<�sa<�ga<�]a<4Va<�Qa<�Pa<WSa<�Xa<�aa<�ka<�va<��a<?�a<��a<�a<8�a<3�a<O�a<�a<�za<na<�aa<[Va<dLa<�Ea<�Aa<�Aa<�Da<�Ja<Ta<�^a<ja<�ta<�~a<��a<��a<��a<>�a<'�a<�wa<�la<s`a<BTa<KIa<@a<:a<.7a<�7a<<a<<Ca<�La<�Wa<�ca<�na<�xa<�a<��a<��a<��a<5za<�pa<�ea<�Ya<#Na<�Ca<b;a<96a<24a<�5a<�:a<�Ba<BMa<�Xa<�da<�  �  �ga<�sa<�|a<�a<��a<��a<i�a<vya<�pa<1ga<�]a<�Ua<�Oa<�Ka<�Ja<+Ma<-Ra<�Ya<�ba<ma<Cwa<q�a<��a<׋a<�a<A�a<?�a<�za<\oa<{ba<�Ta<hHa<�=a< 6a<�1a<�1a<�5a<k=a<*Ha<JUa<da<�ra<��a<�a<O�a<�a<��a<d�a<�a<�a<i�a<y~a<va<�na<ja<�ga<Oha<la<Ira<�za<Єa<N�a<|�a<H�a<��a<�a<ҫa<ާa<��a<J�a<�a<x|a<�na<bba<RXa<Qa<�Ma<8Na<�Ra<�Za<�ea<�ra<0�a<َa<K�a<��a<��a<?�a<)�a<̬a<��a<'�a<��a<�a<�a<�za<
va<�sa<�ta<�xa<a<w�a<��a<Ԛa<��a<t�a<0�a<�a<��a<r�a<��a<�a<�a<�za<#ma<3aa<�Wa<�Qa<-Oa<�Pa<�Va<�_a<1ka<�xa<��a<œa<w�a<t�a<<�a<{�a<��a<z�a<!�a< �a<�a<\�a<�}a<�va<�ra<Eqa<sa<pwa<V~a<��a<u�a<�a<��a<��a<��a<�a<��a<Ңa<֘a<t�a<�~a<ipa<*ca<�Wa<6Oa<'Ja<Ia<�Ka<�Ra<r\a<zha<va<��a<%�a<ךa<S�a<��a<2�a</�a<A�a<��a<��a</�a<5wa<xna<ha<da<ca<Bea<�ia<�pa<Pya<J�a<��a<S�a<4�a<3�a<��a<��a<*�a<�~a<qa<~ba<�Sa<lFa<r;a<W3a</a<�.a<�2a<6:a<�Da<�Pa<~^a<�ka<lwa< �a<��a<��a<�a<2�a<ta<�va<ula<\ba<Ya<[Qa<)La<�Ia<'Ja<�Ma<�Sa<�[a<
ea<�na<�wa<�~a<T�a<��a<a<}a<-ta<yha<9[a<Ma<V?a<e3a<�)a<�#a<�!a<m#a<C)a<w2a<A>a<�Ka<1Za<�  �  z_a<uma<?ya<��a<D�a<��a<��a<�a<_za<�ra<Yka<�da<�_a<�\a<
\a<�]a<6ba<Cha<	pa<jxa<a�a<a�a<6�a<f�a<��a<J�a<�a<_ta<�fa<aWa<IHa<:a<�-a<'%a<s a<@ a<R$a<�,a<�8a<�Ga<8Xa<ia<ya<��a<p�a<�a<t�a<<�a<ٜa<�a<ؑa<ۊa<�a<m~a<pza<�xa<lya<�|a<��a<�a<`�a< �a<�a<q�a<��a<��a<�a<<�a<��a<�a<s�a<�pa<�aa<ZSa<�Ga<�?a<#<a<�<a<�Aa<�Ja<UWa<*fa<�ua<�a<z�a<�a<]�a<
�a<x�a<@�a<C�a<�a<��a<�a<}�a<Ȋa<��a< �a<��a<�a<(�a<��a<��a<��a<��a<ְa<��a<вa<��a<	�a<��a<-�a<�~a<�na<Z_a<�Qa<�Fa<@a<�=a<r?a<�Ea<�Oa<3]a<Dla<|a<��a<I�a<��a<��a<�a<�a<��a<��a<��a<ԛa<��a<��a<�a<��a<s�a<��a<}�a<�a<�a<כa<&�a<z�a<��a<�a<��a<��a<�a<7�a<ƃa<�sa<�ca<�Ta<�Ga<<>a<�8a<�7a<�:a<8Ba<@Ma<+[a<Cja<�ya<��a<S�a<s�a<��a<��a<�a<'�a<ݝa<�a<��a<�a<�}a<dxa<ua<0ta<�ua<�ya<�~a<��a<��a<d�a<}�a<C�a<��a<	�a<�a<�a<Iwa<�ga<�Va<�Fa<e7a<+a<"a<�a<da<�!a<!*a<�5a<Da<+Sa<�ba<�pa<}|a<\�a<~�a<b�a<��a<#�a<fa<�wa<Ooa<rga<Maa<�\a<�Za<[a<�]a<�ba<\ia<qa<�xa<<a<0�a<��a<ąa<k�a<�ya<9na<�`a<�Pa<�@a<�1a<�#a<;a<]a<a<�a<qa<�"a<G0a<�?a<�Oa<�  �   Xa<�ga<qua<�a<��a<��a<؉a<�a<y�a<�|a<�va<jqa<*ma<�ja<Yja<�ka<�oa<�ta<#{a<�a<�a<"�a<�a<L�a<��a<(�a<�{a<�na<�^a<�Ma<=a<>-a<* a<�a<fa< a<�a<�a<�+a<�;a<�Ma<l`a<Yra<�a<_�a<-�a<|�a<6�a<ˡa<�a<��a<7�a<�a<n�a<5�a<��a<��a<_�a<�a<�a<�a<�a< �a<��a<ίa<�a<p�a<k�a<Ėa<��a<xa<�fa<�Ua<=Fa<�9a<01a<�,a<�-a<,3a<�<a<oJa<�Za<3la<�}a<n�a<��a<��a<үa<$�a<�a<ײa<��a<�a<Ңa<�a<�a<��a<S�a<��a<��a<�a<��a<��a<�a<
�a<_�a<�a<l�a<:�a<q�a<g�a<�a<�ua<�ca<�Ra</Da<�8a<;1a<\.a<�0a<j7a<WBa<�Pa<daa<�ra<@�a<ɓa<�a<�a<~�a<m�a<�a<��a<��a<��a<@�a<[�a<��a<��a<Ɛa<ɑa<ؔa<|�a<7�a<S�a<�a<?�a<��a<�a<�a<x�a<P�a<a�a<	|a<?ja<�Xa< Ha<:a<�/a<�)a<F(a<�+a<4a<@a<+Oa<�_a<Eqa<��a<d�a<a�a<Фa<��a<��a<�a<��a<̞a<�a<�a<��a<)�a<[�a<y�a<��a<��a<�a<i�a<��a<��a<��a<q�a<0�a<_�a<�a<0�a<�pa<*_a<�La<�:a<J*a<�a<ta<ba<La<a<6a<�(a<�8a<�Ia<�Za<�ja<xa<��a<C�a<�a<I�a<��a<�a<�a<8za<�sa<�na<�ja<ia<Iia<�ka<�oa<
ua<{a<ـa<��a<��a<9�a<a�a<�a<va<�ha<lYa<�Ga<;6a<9%a<ha<�
a<�a<� a<a<
a<7a<�#a<�4a<}Fa<�  �  (Ra<�ca<�ra<o~a<��a<V�a<�a<��a<��a<�a<[a< {a<�wa<�ua<dua<�va<�ya<6~a<a�a<�a<ߍa<a�a<ʒa<\�a<��a<a�a<�xa<�ia<�Xa<�Fa<34a<�#a<�a<a<�a<�a<�	a<�a<�!a<�2a<�Ea<�Ya<�la<a~a<�a<<�a<�a< �a<\�a<�a<�a<��a<ޘa<A�a<�a<��a<��a<O�a<��a<%�a<ѣa<~�a<?�a<V�a<�a<��a<��a<�a<6�a<I�a<eqa<�^a<vLa<W<a<�.a<u%a<� a<�!a<�'a<O2a<�@a<�Qa<�da<�wa<��a<E�a<�a<`�a<�a<l�a<�a<1�a<�a<�a<=�a<5�a<��a<c�a<��a</�a<��a<Y�a<h�a<A�a<׶a<��a<��a<��a<��a<��a<W�a<7�a<�na<�[a<�Ia<:a<`-a<m%a<M"a<�$a<�+a<8a<*Ga<�Xa<�ka<F~a<��a<�a<��a<x�a<ʵa<��a<Z�a<Աa<��a<ŧa<��a<*�a<��a<ӛa<Ϝa<!�a<�a<w�a<\�a<��a<��a<;�a<�a<��a<��a<)�a<��a<�ua<�ba<�Oa<S>a<�/a<($a<�a<Ca<- a<�(a<	6a<�Ea< Xa<�ja<�|a<��a<�a<ޣa<+�a<�a<��a<ϩa<G�a<��a<��a<͔a<�a<V�a<w�a<}�a<��a<1�a<R�a<|�a<��a<c�a<��a<Ҝa<��a<��a<�|a<�ka<�Xa<�Da<|1a<e a<	a<�a<`a<Ya<ra<�a<Ba<�/a<
Ba<=Ta<�ea<�ta<��a<Љa<��a<ːa<ȏa<��a<Ňa<V�a<,}a<�xa<�ua<ta<Ota<)va<Yya<�}a<{�a<�a<i�a<��a<Ċa<��a<�~a<Psa<�da<�Sa<�@a<�-a<�a<Ba<��`<��`<��`<@�`<��`<�
a<Ca<=,a<b?a<�  �  vNa<�`a<�pa<|}a<��a<f�a<��a<�a<'�a<��a<ӄa<�a<~a<U|a<|a<g}a<4�a<,�a<��a<X�a<I�a<�a<v�a<1�a<p�a<@�a<nva<�fa<�Ta<�Aa<�.a<aa<�a<�a<n�`<��`<�a<�a<;a<�,a<�@a<nUa<yia<�{a<O�a<��a<U�a<��a<��a<�a<��a<�a<��a<��a<y�a<��a<e�a<��a<A�a<ߣa<ըa<��a<h�a<��a<_�a<�a<�a<��a<��a<�a<=ma<�Ya<�Fa<�5a<�'a<Qa<�a<�a<i a<V+a<m:a<.La<�_a<�sa<^�a<�a<Фa<�a<ӵa<	�a<w�a<��a<A�a<7�a<"�a<��a<!�a<�a<��a<��a<۪a<�a<#�a<��a<��a<��a<ʸa<��a<�a<�a<��a<�}a<#ja<dVa<�Ca<J3a<-&a<Ga<1a<�a<�$a<C1a<Aa<�Sa<+ga<�za<��a<'�a<��a<z�a<ڶa<Ըa</�a<o�a<��a<>�a<�a<��a<N�a<��a<J�a<��a<�a<Ьa<Ͱa<�a<$�a<�a<�a<z�a<��a<�a<��a<�qa<^a<MJa<#8a<�(a<a<�a<"a<a<�!a<}/a<@a<�Ra<Efa<ya<�a<N�a<2�a<��a<H�a<�a<�a<:�a<��a<��a<�a<m�a<�a<)�a<�a<ۖa<�a<W�a<��a<�a<��a<�a<W�a<�a<C�a<za<1ha<\Ta<�?a<�+a<�a<�
a<� a<D�`<B�`<Y a<�
a<�a<*a<'=a<DPa<{ba<�ra<�a<v�a<��a<g�a<Q�a<܏a<�a<��a<�a<a<5|a<�za<�za<�|a<�a<=�a<5�a<Ŋa<Q�a<�a<��a<��a<�}a<�qa<ba<Pa<x<a<�(a<�a<�a<s�`<��`<��`<"�`<��`<'a<5a<�&a<�:a<�  �  YMa<�_a<pa<3}a<��a<��a<K�a<��a<~�a<<�a<��a<(�a<Q�a<�~a<�~a<�a<f�a<�a<`�a<Ύa<��a<�a<�a<k�a<`�a<�a<�ua<�ea<�Sa<@a<�,a<.a<aa<�a<��`<��`<3 a<<
a<�a<�*a<?a<Ta<lha<�za<�a<a�a<T�a<ťa<[�a<V�a<U�a<h�a<g�a<��a<��a<Y�a<�a<�a<��a<��a<X�a<�a<��a<}�a<��a<�a<�a<A�a<ďa<�~a<�ka<Xa<�Da<�3a<u%a<�a<�a<�a<	a<�(a<58a<^Ja<^a<Yra<e�a<:�a<��a<�a<��a<o�a<l�a<ĸa<��a<ϱa<��a<ʪa<q�a<˧a<!�a<թa<��a<��a<��a<R�a<�a<1�a<�a<��a<تa<S�a<��a<�|a<�ha<�Ta<�Aa<1a<�#a<�a< a<�a<�"a<�.a< ?a<�Qa<�ea<vya<��a<��a<\�a<w�a<&�a<_�a<U�a<ƶa<�a<��a<�a<̧a<̥a<B�a<��a<��a<˪a<y�a<D�a<`�a<3�a<a�a<+�a<k�a<D�a<I�a<��a<�pa<i\a<vHa<�5a<O&a<�a<�a<a<�a<�a<9-a<>a<Qa<�da<xa<�a<�a<�a<��a<��a<��a< �a<��a<�a<��a<H�a<��a<��a<�a< �a<�a<ța<ٞa<�a<%�a<��a<G�a<]�a<�a<�a<2ya<1ga<
Sa<>a<�)a<�a<�a<�`<:�`<O�`<��`<2a<�a<J(a<k;a<Oa<�aa<�qa<�a<^�a<ޏa<̒a<E�a<�a<��a<1�a<�a<G�a<�~a<z}a<q}a<�~a<��a<�a<��a<!�a<��a<��a<<�a<��a<�}a<�pa<aa<�Na<�:a<�&a<�a<Da<6�`<��`<��`<m�`<@�`<�a<a<%a<-9a<�  �  vNa<�`a<�pa<|}a<��a<f�a<��a<�a<'�a<��a<ӄa<�a<~a<U|a<|a<g}a<4�a<,�a<��a<X�a<I�a<�a<v�a<1�a<p�a<@�a<nva<�fa<�Ta<�Aa<�.a<aa<�a<�a<n�`<��`<�a<�a<;a<�,a<�@a<nUa<yia<�{a<O�a<��a<U�a<��a<��a<�a<��a<�a<��a<��a<y�a<��a<e�a<��a<A�a<ߣa<ըa<��a<h�a<��a<_�a<�a<�a<��a<��a<�a<=ma<�Ya<�Fa<�5a<�'a<Qa<�a<�a<i a<V+a<m:a<.La<�_a<�sa<^�a<�a<Фa<�a<ӵa<	�a<w�a<��a<A�a<7�a<"�a<��a<!�a<�a<��a<��a<۪a<�a<#�a<��a<��a<��a<ʸa<��a<�a<�a<��a<�}a<#ja<dVa<�Ca<J3a<-&a<Ga<1a<�a<�$a<C1a<Aa<�Sa<+ga<�za<��a<'�a<��a<z�a<ڶa<Ըa</�a<o�a<��a<>�a<�a<��a<N�a<��a<J�a<��a<�a<Ьa<Ͱa<�a<$�a<�a<�a<z�a<��a<�a<��a<�qa<^a<MJa<#8a<�(a<a<�a<"a<a<�!a<}/a<@a<�Ra<Efa<ya<�a<N�a<2�a<��a<H�a<�a<�a<:�a<��a<��a<�a<m�a<�a<)�a<�a<ۖa<�a<W�a<��a<�a<��a<�a<W�a<�a<C�a<za<1ha<\Ta<�?a<�+a<�a<�
a<� a<D�`<B�`<Y a<�
a<�a<*a<'=a<DPa<{ba<�ra<�a<v�a<��a<g�a<Q�a<܏a<�a<��a<�a<a<5|a<�za<�za<�|a<�a<=�a<5�a<Ŋa<Q�a<�a<��a<��a<�}a<�qa<ba<Pa<x<a<�(a<�a<�a<s�`<��`<��`<"�`<��`<'a<5a<�&a<�:a<�  �  (Ra<�ca<�ra<o~a<��a<V�a<�a<��a<��a<�a<[a< {a<�wa<�ua<dua<�va<�ya<6~a<a�a<�a<ߍa<a�a<ʒa<\�a<��a<a�a<�xa<�ia<�Xa<�Fa<34a<�#a<�a<a<�a<�a<�	a<�a<�!a<�2a<�Ea<�Ya<�la<a~a<�a<<�a<�a< �a<\�a<�a<�a<��a<ޘa<A�a<�a<��a<��a<O�a<��a<%�a<ѣa<~�a<?�a<V�a<�a<��a<��a<�a<6�a<I�a<eqa<�^a<vLa<W<a<�.a<u%a<� a<�!a<�'a<O2a<�@a<�Qa<�da<�wa<��a<E�a<�a<`�a<�a<l�a<�a<1�a<�a<�a<=�a<5�a<��a<c�a<��a</�a<��a<Y�a<h�a<A�a<׶a<��a<��a<��a<��a<��a<W�a<7�a<�na<�[a<�Ia<:a<`-a<m%a<M"a<�$a<�+a<8a<*Ga<�Xa<�ka<F~a<��a<�a<��a<x�a<ʵa<��a<Z�a<Աa<��a<ŧa<��a<*�a<��a<ӛa<Ϝa<!�a<�a<w�a<\�a<��a<��a<;�a<�a<��a<��a<)�a<��a<�ua<�ba<�Oa<S>a<�/a<($a<�a<Ca<- a<�(a<	6a<�Ea< Xa<�ja<�|a<��a<�a<ޣa<+�a<�a<��a<ϩa<G�a<��a<��a<͔a<�a<V�a<w�a<}�a<��a<1�a<R�a<|�a<��a<c�a<��a<Ҝa<��a<��a<�|a<�ka<�Xa<�Da<|1a<e a<	a<�a<`a<Ya<ra<�a<Ba<�/a<
Ba<=Ta<�ea<�ta<��a<Љa<��a<ːa<ȏa<��a<Ňa<V�a<,}a<�xa<�ua<ta<Ota<)va<Yya<�}a<{�a<�a<i�a<��a<Ċa<��a<�~a<Psa<�da<�Sa<�@a<�-a<�a<Ba<��`<��`<��`<@�`<��`<�
a<Ca<=,a<b?a<�  �   Xa<�ga<qua<�a<��a<��a<؉a<�a<y�a<�|a<�va<jqa<*ma<�ja<Yja<�ka<�oa<�ta<#{a<�a<�a<"�a<�a<L�a<��a<(�a<�{a<�na<�^a<�Ma<=a<>-a<* a<�a<fa< a<�a<�a<�+a<�;a<�Ma<l`a<Yra<�a<_�a<-�a<|�a<6�a<ˡa<�a<��a<7�a<�a<n�a<5�a<��a<��a<_�a<�a<�a<�a<�a< �a<��a<ίa<�a<p�a<k�a<Ėa<��a<xa<�fa<�Ua<=Fa<�9a<01a<�,a<�-a<,3a<�<a<oJa<�Za<3la<�}a<n�a<��a<��a<үa<$�a<�a<ײa<��a<�a<Ңa<�a<�a<��a<S�a<��a<��a<�a<��a<��a<�a<
�a<_�a<�a<l�a<:�a<q�a<g�a<�a<�ua<�ca<�Ra</Da<�8a<;1a<\.a<�0a<j7a<WBa<�Pa<daa<�ra<@�a<ɓa<�a<�a<~�a<m�a<�a<��a<��a<��a<@�a<[�a<��a<��a<Ɛa<ɑa<ؔa<|�a<7�a<S�a<�a<?�a<��a<�a<�a<x�a<P�a<a�a<	|a<?ja<�Xa< Ha<:a<�/a<�)a<F(a<�+a<4a<@a<+Oa<�_a<Eqa<��a<d�a<a�a<Фa<��a<��a<�a<��a<̞a<�a<�a<��a<)�a<[�a<y�a<��a<��a<�a<i�a<��a<��a<��a<q�a<0�a<_�a<�a<0�a<�pa<*_a<�La<�:a<J*a<�a<ta<ba<La<a<6a<�(a<�8a<�Ia<�Za<�ja<xa<��a<C�a<�a<I�a<��a<�a<�a<8za<�sa<�na<�ja<ia<Iia<�ka<�oa<
ua<{a<ـa<��a<��a<9�a<a�a<�a<va<�ha<lYa<�Ga<;6a<9%a<ha<�
a<�a<� a<a<
a<7a<�#a<�4a<}Fa<�  �  z_a<uma<?ya<��a<D�a<��a<��a<�a<_za<�ra<Yka<�da<�_a<�\a<
\a<�]a<6ba<Cha<	pa<jxa<a�a<a�a<6�a<f�a<��a<J�a<�a<_ta<�fa<aWa<IHa<:a<�-a<'%a<s a<@ a<R$a<�,a<�8a<�Ga<8Xa<ia<ya<��a<p�a<�a<t�a<<�a<ٜa<�a<ؑa<ۊa<�a<m~a<pza<�xa<lya<�|a<��a<�a<`�a< �a<�a<q�a<��a<��a<�a<<�a<��a<�a<s�a<�pa<�aa<ZSa<�Ga<�?a<#<a<�<a<�Aa<�Ja<UWa<*fa<�ua<�a<z�a<�a<]�a<
�a<x�a<@�a<C�a<�a<��a<�a<}�a<Ȋa<��a< �a<��a<�a<(�a<��a<��a<��a<��a<ְa<��a<вa<��a<	�a<��a<-�a<�~a<�na<Z_a<�Qa<�Fa<@a<�=a<r?a<�Ea<�Oa<3]a<Dla<|a<��a<I�a<��a<��a<�a<�a<��a<��a<��a<ԛa<��a<��a<�a<��a<s�a<��a<}�a<�a<�a<כa<&�a<z�a<��a<�a<��a<��a<�a<7�a<ƃa<�sa<�ca<�Ta<�Ga<<>a<�8a<�7a<�:a<8Ba<@Ma<+[a<Cja<�ya<��a<S�a<s�a<��a<��a<�a<'�a<ݝa<�a<��a<�a<�}a<dxa<ua<0ta<�ua<�ya<�~a<��a<��a<d�a<}�a<C�a<��a<	�a<�a<�a<Iwa<�ga<�Va<�Fa<e7a<+a<"a<�a<da<�!a<!*a<�5a<Da<+Sa<�ba<�pa<}|a<\�a<~�a<b�a<��a<#�a<fa<�wa<Ooa<rga<Maa<�\a<�Za<[a<�]a<�ba<\ia<qa<�xa<<a<0�a<��a<ąa<k�a<�ya<9na<�`a<�Pa<�@a<�1a<�#a<;a<]a<a<�a<qa<�"a<G0a<�?a<�Oa<�  �  �ga<�sa<�|a<�a<��a<��a<i�a<vya<�pa<1ga<�]a<�Ua<�Oa<�Ka<�Ja<+Ma<-Ra<�Ya<�ba<ma<Cwa<q�a<��a<׋a<�a<A�a<?�a<�za<\oa<{ba<�Ta<hHa<�=a< 6a<�1a<�1a<�5a<k=a<*Ha<JUa<da<�ra<��a<�a<O�a<�a<��a<d�a<�a<�a<i�a<y~a<va<�na<ja<�ga<Oha<la<Ira<�za<Єa<N�a<|�a<H�a<��a<�a<ҫa<ާa<��a<J�a<�a<x|a<�na<bba<RXa<Qa<�Ma<8Na<�Ra<�Za<�ea<�ra<0�a<َa<K�a<��a<��a<?�a<)�a<̬a<��a<'�a<��a<�a<�a<�za<
va<�sa<�ta<�xa<a<w�a<��a<Ԛa<��a<t�a<0�a<�a<��a<r�a<��a<�a<�a<�za<#ma<3aa<�Wa<�Qa<-Oa<�Pa<�Va<�_a<1ka<�xa<��a<œa<w�a<t�a<<�a<{�a<��a<z�a<!�a< �a<�a<\�a<�}a<�va<�ra<Eqa<sa<pwa<V~a<��a<u�a<�a<��a<��a<��a<�a<��a<Ңa<֘a<t�a<�~a<ipa<*ca<�Wa<6Oa<'Ja<Ia<�Ka<�Ra<r\a<zha<va<��a<%�a<ךa<S�a<��a<2�a</�a<A�a<��a<��a</�a<5wa<xna<ha<da<ca<Bea<�ia<�pa<Pya<J�a<��a<S�a<4�a<3�a<��a<��a<*�a<�~a<qa<~ba<�Sa<lFa<r;a<W3a</a<�.a<�2a<6:a<�Da<�Pa<~^a<�ka<lwa< �a<��a<��a<�a<2�a<ta<�va<ula<\ba<Ya<[Qa<)La<�Ia<'Ja<�Ma<�Sa<�[a<
ea<�na<�wa<�~a<T�a<��a<a<}a<-ta<yha<9[a<Ma<V?a<e3a<�)a<�#a<�!a<m#a<C)a<w2a<A>a<�Ka<1Za<�  �  pa<�ya<��a<��a<��a<��a<}za<�pa<)fa<fZa<IOa<pEa<�=a<�9a<v8a<;a<�@a<�Ia<�Ta<�`a<!ma<pxa<8�a<��a<��a<:�a<��a<فa<Pxa<�ma<Yba<�Wa<�Na<Ha<�Da<eDa<�Ga<�Na<?Xa<�ca<Tpa<�|a<T�a<�a<:�a<��a<�a<.�a<)�a<��a< |a<�pa<�fa<^a<?Xa<kUa<Va<*Za<Maa<~ka<wa<̃a<�a<5�a<�a<��a<L�a<��a<�a<�a<��a<z�a<�|a<Sra<Gia<Mca<O`a<�`a<�da<�ka<�ua<��a<��a<�a<i�a<"�a<��a<�a<N�a<��a<۞a<:�a<��a<�|a<Nra<�ia<�ca<paa<�ba<
ga<�na<�xa<�a<�a<-�a<F�a<k�a<��a<7�a<�a<��a<V�a<|�a<��a<�{a<�qa<.ia<�ca<�aa<nca<3ha<pa<5za<��a<l�a<<�a<ǥa<)�a<��a<j�a<m�a<��a<��a<h�a<7�a<�wa<Wma<\ea<{`a<�^a<�`a<fa<`na<�xa<,�a<ݏa<��a<��a<q�a<~�a<��a<�a<��a<g�a<�a<�}a<�ra<�ha<"aa<�\a<�[a<C^a<�ca<�la<�va<b�a<��a<��a<J�a<@�a<f�a<D�a<��a<z�a<t�a<e�a<�sa<�ga<�]a<4Va<�Qa<�Pa<WSa<�Xa<�aa<�ka<�va<��a<?�a<��a<�a<8�a<3�a<O�a<�a<�za<na<�aa<[Va<dLa<�Ea<�Aa<�Aa<�Da<�Ja<Ta<�^a<ja<�ta<�~a<��a<��a<��a<>�a<'�a<�wa<�la<s`a<BTa<KIa<@a<:a<.7a<�7a<<a<<Ca<�La<�Wa<�ca<�na<�xa<�a<��a<��a<��a<5za<�pa<�ea<�Ya<#Na<�Ca<b;a<96a<24a<�5a<�:a<�Ba<BMa<�Xa<�da<�  �  �xa<�a<�a<o�a<�a<#}a<ta<Vha<?[a<MMa<,@a<�4a<G,a<'a<�%a<�(a<�/a<{9a<�Ea<'Ta<�ba<Qpa<U|a<u�a<d�a<��a<j�a<+�a<6�a<�xa<�oa<�fa<+_a<�Ya<�Va<�Va<�Ya<�_a<�ga<�qa<5|a<��a<ݏa<֖a<�a<��a<��a<x�a<�a<I}a<zpa< ca<)Wa<HMa<'Fa<�Ba<\Ca<�Ga<iPa<�[a<ia<�wa<f�a<��a<�a<"�a<��a<��a<��a< �a<O�a<�a<��a<΁a<Vza<Cua<�ra<sa<�va<�|a<��a<�a<�a<2�a<	�a<6�a<��a<<�a<@�a<"�a<�a<�a< |a<Lna<#ba<aXa<�Qa<�Na<Pa<1Ua<�]a<Bia<�va<لa<Z�a<��a<E�a<��a<ѱa<�a<?�a<��a<��a<��a<c�a<��a<�za<va<Gta<�ua<�ya<X�a<Ԉa<<�a<�a<��a<��a<��a<��a<խa<��a<�a<��a<|�a<va<�ha<�\a<�Sa<�Ma<-La<~Na<�Ta<^a<�ia<�wa<m�a<^�a<��a<#�a<`�a<��a<��a<��a<L�a<�a<�a<��a<ya<�ra<�na<na<Hpa<ua<1|a<�a<E�a<��a<��a<2�a<��a<a�a<�a<F�a<;�a<�a<�ta<�ea<NXa<�La<Da< ?a< >a<+Aa<Ha<�Qa<�]a<�ja<�wa<Ãa<��a<`�a<�a<��a<�a<W�a<e�a<!za<�oa<�ea<r]a<�Wa<Ta<�Sa<�Va<�[a<=ca<�ka<0ua<�}a<,�a<ɉa<��a<��a<3�a<�{a<�oa<rba<Ta<�Ea<$9a<�.a<�'a<�$a<b%a<8*a<�2a<�=a<�Ja<�Xa<�ea<�qa<h{a<��a<��a<��a<�a<�xa<pa<0fa<�\a<�Sa<�La<SHa<�Fa<Ha<`La<)Sa<�[a<�ea<toa<�  �  �a<��a<�a<�a<]�a<Iya<�ma<`a<�Pa<�@a<2a<-%a<ka<�a<Xa<Ka<�a<*a<J8a<Ha<�Xa<�ha<}va<1�a<'�a<Ďa<��a<��a<�a<��a<�{a<`ta<bna<�ia<�ga<�ga<~ja<�oa<8va<�~a<E�a<f�a<j�a</�a<�a<^�a<l�a<��a<��a<9ta<ea<LVa<pHa<=a<
5a<F1a<�1a<�6a<@a<�La<\a<Qla<}a<��a<
�a<��a<c�a<�a<��a<m�a<إa<��a<Z�a<�a<�a<��a<��a<)�a<�a<�a<p�a<Q�a</�a<?�a<̮a<�a<رa</�a<?�a<�a<Z�a<�a<1pa<�`a<�Ra<�Ga<F@a<E=a<�>a<?Da<Na<�Za<ja<�ya<ˉa<
�a<�a<�a<��a<ʳa<�a<��a<�a<|�a<��a<H�a<��a<ֆa<t�a<k�a<�a<.�a<$�a<�a<i�a<��a<��a<��a<�a<-�a<��a<͗a<��a<�ya<�ia<qZa<Ma<�Ba<w<a<�:a<=a<Da<�Na<G\a<nka<4{a<��a<ؗa<ܢa< �a<�a<l�a<��a<�a<�a<,�a<#�a<S�a<�a<�a<2a<׀a<�a<��a<őa<W�a<H�a<�a<��a<$�a<	�a<��a<}�a<Q�a<
za<Tia<Ya<�Ia<�<a< 3a<�-a<�,a<�/a<�7a<�Ba<�Pa<J_a<�na<�|a<��a<��a<L�a<��a<�a<��a<�a<��a<V|a<�sa<7ma<�ga<,ea<�da<�fa<'ka<�pa<=xa<~a<��a<��a<��a<��a<��a<5�a<�ua<Hha<�Xa<"Ha<V8a<�)a<aa<pa<
a<�a<Ja<�"a<_/a<">a<�Ma<a]a<cka<=wa<�a<��a<c�a<u�a<�a<Cya<�qa<�ia<lba<�\a<Ya<�Wa<�Xa<}\a<�aa<*ia<5qa<�xa<�  �  ݅a<�a<K�a<3�a<�a<`ua<-ha<�Xa<SGa<�5a<�%a<�a<a<�a<a<�a<�a<�a<	,a<�=a<�Oa<�aa<Gqa<�~a<�a<}�a<��a<S�a<��a<�a<��a<&�a<J{a<�wa<�ua<5va<xxa<�|a<��a<^�a<p�a<Жa<�a<��a<��a<�a<�a<7�a<�{a<&la<G[a<�Ja<;a<#/a<}&a<)"a<�"a</(a<2a<�?a<TPa<Uba<�ta<9�a<d�a<�a<תa<7�a<��a<��a<�a<�a<��a<+�a<@�a<��a<�a<g�a<��a<�a<\�a<��a<ƪa<��a<��a<δa<Ʋa<)�a<
�a<w�a<��a<dwa<�ea<�Ta<�Ea<�9a<�1a< .a<|/a<�5a<?@a<@Na<�^a<{pa<'�a<J�a< �a<ߪa<�a<ӵa<�a<p�a<ծa<�a<Ţa<�a<�a<�a<ɓa<��a<[�a<�a<��a<��a<l�a<	�a<ȴa<Ҵa<a�a<c�a<Пa<9�a<>�a<�pa<�^a<�Ma<f?a<k4a<�-a<^+a<D.a<�5a<9Aa<Pa<�`a<Yra<��a<��a<d�a<٨a<��a<�a<$�a<��a<r�a<D�a<�a<<�a<��a<(�a<��a<юa<%�a<�a<��a<��a<��a<��a<�a<��a<��a</�a<�a<)�a<�qa<�_a<�Ma<�<a<�.a<s$a<�a<ya<[!a<�)a<�5a<�Da<NUa<Afa<Ava<�a<*�a<��a<՚a<`�a<�a<$�a<�a<�a<.�a<Xza<�ua<ysa<sa<�ta<xa<�|a<��a<�a<��a<ɏa<d�a<ύa<��a<~a<�pa<uaa<�Oa<�=a<C,a<�a<)a<�a<�a<�a<�
a<�a<�"a<3a<RDa<�Ua<�ea<"sa<�}a<ބa<j�a<v�a<ąa<�a<;{a<�ta<oa<?ja<$ga<fa<ga<�ia<�na<�ta<�za<�a<�  �  f�a<�a<��a<�a<~a<lra<�ca<�Ra<%@a<j-a<�a<3a<�a<��`<��`<��`<Ka<�a<�"a<J5a<�Ha<�[a<Rma<	|a<��a<��a</�a<��a<i�a<j�a<8�a<�a<��a<S�a<�a<?�a<{�a<�a<֋a<o�a<@�a<Y�a<��a<�a<��a<�a<ԑa<څa<�va<�ea<�Sa<�Aa<�1a<k$a<�a</a<�a<ya<1'a<�5a<Ga<�Za<.na<�a<�a<��a<#�a<�a<4�a<��a<i�a<��a<��a<U�a<;�a<��a<�a<e�a<{�a<��a<<�a<E�a<0�a<��a<�a<��a<$�a< �a<x�a<��a<��a<�pa<�]a<_Ka<�;a<l.a<�%a<�!a<�#a<9*a<�5a<�Da<Va<.ia<�{a<��a<�a<1�a<�a<��a<иa<ȷa<��a<*�a<�a<[�a<r�a<��a<՞a<��a<աa<q�a< �a<�a<p�a<��a<Ʒa<�a<K�a<�a<ܜa<ލa<1|a<]ia<2Va<LDa<5a<�(a<�!a<Oa<x"a<x*a<7a<�Fa<�Xa<hka<�}a<��a<��a<��a<�a<��a<t�a<|�a<��a<Ũa<��a<�a<n�a<+�a<��a<֙a<>�a<'�a<��a<V�a<>�a<��a<~�a<��a<,�a<�a<��a<,~a<}ka<
Xa<fDa<�2a<�#a<�a<�a<wa<�a<�a<�+a<�;a<�Ma<�_a<qa<��a<�a<
�a<��a<��a<��a<{�a<��a<�a<W�a<R�a<ـa<z~a<	~a<da<�a<ʅa<1�a<��a<��a<D�a<5�a<.�a<��a<r{a<%ma<�[a<	Ia<�5a<�"a<�a<a<��`<��`<�`<H�`<}
a<a<<*a<=a<�Oa<aa<pa<|a<��a<��a<@�a<�a<�a<S�a<5}a<yxa<�ta<(ra<!qa<ra<kta<8xa< }a</�a<��a<�  �  .�a<��a<��a<�a<}a<vpa<�`a<�Na<~;a<(a<�a<aa<e�`<��`<��`<��`<�`<�a<�a<0a<MDa<7Xa<�ja<Oza<�a<�a<j�a<��a<\�a<.�a< �a<v�a<+�a<Èa<��a<�a<�a<9�a<��a<��a<��a<��a<]�a<��a<4�a<�a<��a<��a<�sa<�aa<�Na<<a<g+a<ha<�a<a<�a<Xa< a<f/a<oAa<�Ua<ja<�}a<l�a<H�a<��a<��a<��a<�a<��a<ɲa<	�a<�a<��a<�a<£a<�a<�a<�a<�a<%�a<�a<�a<H�a<�a<x�a<i�a<ןa<��a<~a<Ela<�Xa<�Ea<�4a<H'a<�a<�a<�a<#a<�.a<t>a<�Pa<pda< xa<��a<ؚa<�a<��a<ڷa<��a<w�a<(�a<��a<v�a<\�a<רa<u�a<��a<(�a<?�a<��a<q�a<��a<��a<]�a<��a<�a<;�a<�a<�a<�a<sxa<�da<�Pa<4>a<:.a<�!a<�a<3a<Ra<I#a<l0a<�@a<eSa<�fa<8za<ދa<��a<צa<)�a<�a<z�a<n�a<��a<��a<9�a<�a<ݡa<̟a<;�a<@�a<��a<��a<ީa<��a<��a<�a<�a<A�a<ǥa<ښa<U�a<�za<xga<Sa<�>a<�,a<�a<�a<ta<]
a<�a<�a<m%a<�5a<�Ha<�[a<�ma<~a<��a<��a<!�a<�a<"�a<��a<Ƙa<�a<�a<��a<=�a<+�a<��a<υa<!�a<q�a<�a<d�a<��a<o�a<��a<��a<�a<�ya<rja<rXa<�Da<�0a<a<�a<��`<��`<��`<��`< �`<�a<�a<�$a<H8a<�Ka<�]a<�ma<{a<t�a<n�a<��a<Ɍa<a�a<Άa<��a<x~a<�za<�xa<�wa<�xa<�za<K~a<p�a<��a<��a<�  �  ��a<��a<ςa<S~a<;wa<�ma<�aa<�Sa<8Ea<�6a<,)a<�a<�a<�a<4a<Sa<+a<H"a</a<�=a<�La<F\a<Oja<�va<m�a<��a<N�a<}�a<�a<x�a<`�a<��a<��a<߄a<�a<��a<4�a<�a<8�a</�a<�a<;�a<A�a<2�a<B�a<s�a<4�a<?�a<Eua<�ga<�Ya<La<w?a<G5a<0.a<�*a<+a<�/a<B8a<�Ca<�Qa<�`a<:pa<ma<�a<��a<��a<�a<��a<�a<o�a<��a<Ƨa<Ϥa<��a<��a<��a<ߟa<[�a<ãa<��a<�a<֬a<�a<{�a<!�a<��a<�a<F�a<��a<s�a<�sa<ea<�Va<GJa<V@a<�9a<}6a<�7a<.=a<�Ea<�Qa<g_a<na<�|a<�a<��a<ԡa<p�a<w�a<��a<%�a<��a<�a<ĩa<��a<J�a<Z�a<��a<�a<��a<�a<ܨa<�a<��a<%�a<ʯa<��a<רa<c�a<b�a<�a<�|a<�ma<_a<�Pa<�Da<�;a<�5a<�3a<v6a<�<a<BFa<iRa<�`a< oa<�}a<�a<Ŗa<ҟa<p�a<H�a<��a<d�a<6�a<W�a<բa<�a<\�a<��a<N�a<�a<ʝa<�a<͢a<��a<��a<]�a<�a<ңa<��a<�a<��a<I|a<8ma<�]a<�Na<�@a<�4a<',a<�&a<�%a<E)a<0a<:a<^Fa<Ta<'ba<�oa<4|a<��a<�a<P�a<��a<�a<9�a<?�a<�a<��a<`�a<��a<́a<@�a<��a<��a<υa<��a<Ҋa<g�a<H�a<\�a<=�a<?a<�ua<�ia<\a<�La<�=a<�.a<�!a<�a<ra<�a<�a<�a<Qa<�&a<54a<�Ba<GQa<,_a<yka<wua<�|a<Ła<ڃa<5�a<��a<�a<�|a<�ya<2wa<Rua<�ta<<ua<wa<�ya<�|a<�a<Âa<�  �  ȃa<E�a<��a<H~a<twa<na<hba<�Ta<�Fa<$8a<�*a<=a<�a<�a<ga<Ga<�a<�#a<t0a<	?a<3Na<E]a<ka<wa<��a<��a<�a<�a<�a<l�a< �a<a�a<�a<)�a<k�a<��a<z�a<L�a<�a<��a<��a<=�a<��a<�a<�a<��a<x�a<�a<2va<�ha<�Za<EMa<Aa<�6a<�/a<�,a<:-a<�1a<�9a<DEa<�Ra<ba<oqa<_�a<��a<�a<��a<�a<X�a<]�a<r�a<o�a<��a<~�a<Ša<Ϟa<�a<9�a<��a<�a<=�a<��a<ƫa<�a<��a<��a<{�a<M�a<��a<w�a<i�a<�ta<Xfa<*Xa<�Ka<�Aa<{;a<�8a<�9a<�>a<{Ga<Sa<�`a<\oa<!~a<�a</�a<�a<k�a<<�a<d�a<O�a<��a<�a<��a<M�a<��a<��a<�a<d�a<	�a<��a<��a<�a<��a<D�a<s�a<l�a<˨a<��a<ߗa<ϋa<�}a<!oa<I`a<^Ra<uFa<J=a<�7a<6a<j8a<E>a<�Ga<�Sa<�aa<Lpa<�~a<݋a<+�a<
�a<c�a<�a<G�a<k�a<+�a<�a<��a<F�a<��a<�a<��a<4�a<�a<��a<��a<u�a<��a<��a<ͦa<��a<��a<S�a<T�a<5}a<mna<_a<�Oa<Ba<[6a<�-a<)a<(a<+a<�1a<�;a<�Ga<dUa<\ca<�pa<�|a<Նa<;�a<(�a<g�a<C�a<<�a<*�a<F�a<@�a<��a<ʁa<�a<�a<D�a<��a<�a<I�a<a<f�a<ɋa<3�a<(�a<oa<=va<�ja<�\a<Na<�>a<O0a<�#a<"a<Ua<a<�a<�a<�a<((a<u5a<�Ca<iRa<`a<la<�ua<�|a<��a<��a<_�a<��a<�~a<m{a</xa<yua<�sa<sa<�sa<`ua<xa<^{a<�~a<��a<�  �  ��a<܂a<��a<V~a<?xa<uoa<tda<�Wa<�Ia<$<a<M/a<J$a<�a<a<�a<�a<�a<�(a<�4a<�Ba<�Qa<�_a< ma<Exa<E�a<�a<!�a<��a<��a<��a<d�a<<�a<P�a<F~a<h}a<�}a<�a<k�a<��a<��a<��a<��a<��a<��a<��a<�a<q�a<��a<rxa<�ka<�^a<{Qa<�Ea<�;a<H5a<2a<�2a<7a<�>a<Ja<'Wa<�ea<�ta<��a<q�a<�a<.�a<k�a<+�a<��a<��a<0�a<��a<3�a<��a<�a<ژa<.�a<��a<j�a<�a<ߤa<Ĩa<��a<a�a<�a<(�a<ڤa<��a<O�a<څa<?xa<4ja<�\a<�Pa<!Ga<�@a<�=a<L?a<(Da<�La<�Wa<�da<�ra<Հa<�a<��a<�a<��a<u�a<�a<<�a<�a<`�a<z�a<Ԡa<��a<��a<њa<l�a<�a<	�a<��a<J�a<ͪa<!�a<	�a<��a<ڨa<g�a<>�a<ڍa<��a<�ra<Ida<�Va<�Ka<�Ba<K=a<f;a<�=a<�Ca<�La<SXa<�ea<�sa<2�a<Ǎa<]�a<��a<1�a<�a<éa<&�a<M�a<\�a<g�a<��a<a<�a<k�a<G�a<&�a<B�a<��a<#�a<�a<��a<��a<�a<!�a<L�a<��a<ua<^qa<�ba<
Ta<�Fa<~;a<?3a<m.a<q-a<o0a<�6a<k@a<�Ka<"Ya<mfa<;sa<�~a<ևa<��a<��a<:�a<g�a<��a<�a<R�a<��a<�a<�|a<{a<�za<d{a<X}a<P�a<{�a<��a<�a<-�a<#�a<ԅa<�a<Zwa<dla<m_a<TQa<�Ba<�4a<}(a<ca<�a<qa<aa<�a<�!a<�,a<�9a<iGa<Ua<+ba<uma<�va<}a<Āa<<�a<L�a<�~a<L{a<]wa<�sa<�pa<�na<�ma<�na<tpa<�sa<Hwa<D{a<
a<�  �  ~a<Q�a<p�a<9~a<6ya<�qa<�ga<\a<MOa<�Ba<X6a<,a<K$a<�a<�a<9!a<J'a<V0a<�;a<Ia<�Va<�ca<
pa<Bza<��a<&�a<��a<��a<هa<��a<��a<�|a<ya<iva<)ua<sua<~wa<�za<�a<ӄa<R�a<p�a<i�a<��a<��a<�a<܍a<�a<|a<pa<Bda<6Xa<�La<Da<�=a<�:a<R;a<�?a<Ga<ZQa<�]a<{ka<Hya<v�a<�a<��a<|�a<��a<�a<y�a<פa<�a<��a<H�a<��a<ݑa<��a<�a<ђa<�a<R�a<��a<��a<ǧa<��a<&�a<��a<o�a<��a<;�a<�a<@}a<8pa<�ca<8Xa<^Oa<mIa<�Fa<�Ga<�La<bTa<�^a<;ka<Lxa<V�a<��a<�a<�a<��a<L�a<��a<Ϊa<V�a<ܢa<%�a<��a<��a<��a<��a<7�a<f�a<ߘa<�a<��a<�a<��a<}�a<J�a<��a<^�a<q�a<"�a<�a<�wa<�ja<^a<<Sa<	Ka<�Ea<5Da<`Fa<�Ka<TTa<Q_a<�ka<�xa<_�a<Ӑa<\�a<c�a<٥a<��a<��a<[�a<U�a<��a<Ėa<c�a<�a<Ìa<"�a<8�a<��a<D�a<o�a<ϛa<��a<��a<h�a<-�a<S�a<��a<��a<�a<va<Qha<�Za<Na<�Ca<�;a<+7a<46a<�8a<�>a<�Ga<�Ra<�^a<6ka<�va<=�a<g�a< �a<�a</�a<a�a<��a<��a<F�a<}a<axa<�ta<�ra<Kra<usa<va<�ya<�}a<��a<(�a<M�a<`�a<_�a<��a<8ya<Ooa<wca<TVa<�Ha<�;a<�/a<�&a<D a<;a<	a<["a<�)a<�3a<@a<�La<�Ya<�ea<�oa<�wa<}a<�a<�a<�}a<Rza<�ua<qa<�la<�ha<�fa<�ea<jfa<�ha<hla<�pa<�ua<Xza<�  �  xya<}a<�~a<�}a<cza<]ta<�ka<�aa<Va<�Ja<�?a<36a</a<�*a<�)a<-,a<�1a<U:a<�Da<�Pa<*]a<;ia<�sa<�|a<ła<��a<��a<$�a<�a</~a< ya<�sa<Woa<la<�ja<�ja<�la<�pa<Hva<�|a<^�a<ǉa<@�a<֒a<w�a<:�a<��a<3�a<��a<�va<vka<�`a<�Va<|Na<�Ha<�Ea<�Fa<pJa<�Qa<[a<�fa<�ra<�a<:�a<a�a<�a<âa<��a<��a<s�a<V�a<�a<��a<�a<��a<K�a<�a<I�a<`�a<J�a<[�a<D�a<*�a<��a<¦a<�a<�a<�a<ߠa<Иa<�a<��a<�wa<zla<ba<�Ya<[Ta<3Ra<Sa<`Wa<�^a<2ha<xsa<;a<&�a<a<Ξa<j�a<e�a<ժa<��a<S�a<]�a<��a<��a<:�a<؋a<݈a<߇a<��a<.�a<J�a<��a<Z�a<��a<�a<=�a<��a<n�a<��a<'�a<0�a<��a<�~a<�ra<Tga<q]a<�Ua<�Pa<�Oa<WQa<�Va<V^a<`ha<�sa<Ja<��a<��a<��a</�a<Q�a<��a<f�a<o�a<�a<��a<�a<��a<��a<�a<��a<��a<��a<��a<K�a<ٔa<�a<Z�a<��a<�a<r�a<k�a<��a<��a<)|a<�oa<Kca<�Wa<�Ma<�Fa<`Ba<Aa<�Ca<rIa<WQa<p[a<2fa<qqa<�{a<��a<P�a<I�a<�a<��a<[�a<#�a<܀a<Iza<�sa<una<Ija<ha<�ga<ia<:la<�pa<�ua<&{a<�a<��a<>�a<��a</�a<u{a<�ra<�ha<�\a<mPa<�Da<�9a<:1a<0+a<�(a<)a<-a<4a<H=a<DHa<�Sa<m_a<�ia<�ra<ya<�|a<&~a<�|a<gya<\ta<�na<�ha<"ca<�^a<�[a<�Za<�[a<�^a<�ba<Gha<Xna<7ta<�  �  �sa<ya<z|a<r}a<�{a<Pwa<wpa<�ga<^a<�Sa<.Ja<�Aa<~;a<�7a<�6a<9a<7>a<�Ea<9Oa<�Ya<�da<(oa<xa<4a<��a<��a<�a<Ła<�|a<�va<�oa<�ia<�ca<�_a<�]a<^a<�`a<2ea<�ka<sa<+{a<�a<�a<o�a<��a<e�a<_�a<a<ޅa<r}a<�sa<pja<�aa<\Za<QUa<�Ra<�Sa<5Wa<�]a<%fa<kpa<k{a<��a<��a<$�a<z�a<'�a<�a<a�a<v�a<˘a<�a<�a<{�a<�~a<	{a<0ya<�ya<3|a<׀a<��a<�a<��a<{�a<0�a</�a<ߧa<ۦa<<�a<��a<Ȕa<�a<��a<�va<wma<.fa<9aa<1_a<
`a<�ca<eja<�ra<�|a<_�a<��a<��a<�a<ݦa<%�a<��a<��a<Ƞa<R�a<�a<ŋa<:�a<�a<d|a< {a<�{a<)a<)�a<z�a<��a<Řa<5�a<:�a<R�a<��a<֥a<�a<��a<�a<��a<|a<�qa<
ia<Bba<�]a<�\a<>^a<�ba<�ia<�ra<�|a<�a<��a<�a<S�a<$�a<b�a<�a<�a<i�a<m�a<�a<��a<Q}a<exa<lua<�ta<Hva<�ya<Aa<��a<��a<^�a<-�a<F�a<@�a<��a<6�a<2�a<ߌa<��a<�wa<�la<�ba<�Ya<GSa<aOa<�Na<�Pa<iUa<w\a<@ea<�na<uxa<�a<K�a<L�a<��a<]�a<s�a<`�a<��a<�xa<�pa<Bia<�ba<^a<][a<�Za<�\a<�`a<;fa<�la<{sa<�ya<�~a<f�a<��a<��a<�}a<wa<Una<+da<NYa<�Na< Ea<i=a<8a<�5a<6a<�9a<�?a<Ha<�Qa<�[a<�ea<�na<�ua<�za<�|a<|a<�xa<�sa<Tma<fa<�^a<%Xa<�Ra<fOa<9Na<7Oa<�Ra<�Wa<=^a<�ea<ma<�  �  uma<�ta<�ya<�|a<�|a<@za<]ua<jna<afa<�]a<aUa<Na<�Ha<wEa<�Da<�Fa<0Ka<�Qa<%Za<bca<�la<Gua<�|a<��a<f�a<_�a<�a<�|a<$va<Tna<fa<2^a<rWa<�Ra<TPa<qPa<?Sa<PXa<�_a<|ha<!ra<�{a<b�a<��a<��a<@�a<�a<b�a<M�a<��a<�|a<�ta<3ma<�fa<�ba<�`a<raa<�da<7ja<�qa<�za<��a<̍a<5�a<��a<G�a<6�a<0�a<Ξa<��a<��a<<�a<��a<�xa<#ra<�ma<�ka<�ka<oa<1ta<�{a<��a<��a<��a<(�a< �a<a�a<Y�a<x�a<I�a<��a<Ȓa<!�a<^�a<}ya<sa<�na<ma<�ma<;qa<�va<I~a<��a<ۏa<J�a<��a<�a<�a<��a<=�a<��a<��a<�a<��a<�a<ya<�ra<oa<pma<�na<$ra<�wa<ua<�a<ʐa<�a<�a<��a<�a<�a<�a<Ǟa<n�a<��a<�a<}a<Qua<roa<�ka<�ja<la<�oa<�ua<�}a<-�a<ˎa<Ėa<k�a<͡a<գa<�a<�a<<�a<��a<�a<��a<\xa<�pa<Lka<�ga<ga<�ha<ma<bsa<{a<��a<�a<y�a<��a<*�a<u�a<לa<Ҙa<M�a<�a<ڀa<>wa<;na<`fa<�`a<6]a<U\a<^a<ba<>ha<�oa<�wa<�a<��a<"�a<�a<��a<x�a<�a<�a<Vya<�oa<\fa<�]a<Va<�Pa<�Ma<cMa<�Oa<"Ta<�Za<�ba<�ja<�ra<�ya<6a<�a<s�a<
�a<U{a<Ita<�ka<�ba<wYa<#Qa<EJa<�Ea<wCa<�Ca<�Fa<La<[Sa<�[a<ada<�la<�sa<�xa<�{a<|a<�ya<�ta<�ma<�ea<�\a<�Sa<La<�Ea<	Ba<�@a<�Aa<�Ea<rKa<;Sa<\a<ea<�  �  ga<�oa<
wa<�{a<�}a<�|a<�ya<�ta<ona<bga<v`a<dZa<�Ua<�Ra<qRa<(Ta<"Xa<�]a<�da<�la<_ta<H{a<��a<�a<�a<�a<�~a<�wa<^oa<�ea<�[a<�Ra<Ka<Ea<�Ba<�Ba<�Ea<�Ka<�Sa<�]a<�ha<ta<�~a<��a<��a<ݒa<��a<��a<q�a<��a<j�a<�~a<�xa<�sa<�oa<Yna<oa<�qa<wa<�}a<*�a<J�a<��a<��a<r�a<�a<�a<I�a<ښa<C�a<'�a<�a<va<�la<pea<,`a<�]a<)^a<�aa<�ga<�oa<�ya<3�a<��a<їa<�a<ڤa<��a<��a<#�a<��a<V�a<D�a<�a<n�a<�a<A|a<�za<[{a<Q~a<7�a<��a<��a<�a<�a<`�a<�a<A�a<��a<��a<��a<v�a<~�a<�a<�ua<�la<�ea<;aa<�_a<�`a< ea<�ka<Qta<A~a<��a<��a<�a<�a<(�a<ԧa<��a<>�a<؝a<�a<��a<3�a<��a<~|a<0ya<2xa<]ya<�|a<��a<\�a<}�a<��a<Ȝa<x�a<+�a<W�a<ʡa<��a<�a<�a<��a<�va<�la<gda<�]a<Za<CYa<M[a<8`a<kga<_pa<Hza<Y�a<��a<X�a<�a<�a<p�a<�a<p�a<�a<w�a<^�a<�ya<sa<�ma<�ja<�ia<Wka<�na<�sa<za<��a<�a<�a<��a<�a<��a<��a<�a<0|a<�qa<�fa<�[a<�Qa<OIa<-Ca<�?a<�?a<IBa<�Ga<6Oa<gXa<-ba<�ka<�ta<�{a<��a<��a<8�a<-a<za<^sa<�ka<da<]a<+Wa<Sa< Qa<fQa<Ta<�Xa<�^a<xea<�la<7sa<mxa<�{a<�|a<:{a<�va<0pa<�ga<�]a<Sa<�Ha<�?a<�8a<D4a<�2a<4a<f8a<6?a<Ha<ERa<�\a<�  �  �`a<Nka<.ta<qza<B~a<Wa<�}a<�za<�ua<6pa<�ja<�ea<�aa<}_a<-_a<�`a<da<�ha<�na<,ua<S{a<��a<Y�a<�a<	�a<��a<^{a<�ra<�ha<�]a<~Ra<�Ga<R?a<�8a<�5a<�5a<�8a<a?a<wHa<�Sa<`a<�la<�xa<r�a<A�a<*�a<ߕa<��a<!�a<ˑa<)�a<'�a<)�a<a<#|a<{a<�{a<8~a<��a<�a<��a<2�a<i�a<u�a<��a<��a<��a<3�a<��a<ˍa<
�a<bwa<2la<�aa<hYa<`Sa<�Pa<'Qa<�Ta<�[a<�da<*pa<�{a<؇a<��a<�a<(�a<��a<��a<��a<եa<%�a<��a<��a<9�a<��a<��a<v�a<�a<q�a<��a<��a<��a<��a<�a<��a<��a<�a<��a<��a<��a<p�a<ɂa<�va<�ka<raa<�Ya<PTa<�Ra<�Sa<�Xa<`a<�ia<ua<��a<P�a<t�a<�a<�a<k�a<"�a<V�a<��a<P�a<g�a<L�a<܌a<��a<Ʌa<�a<΅a<��a<�a<:�a<��a<��a<<�a</�a<8�a<|�a<C�a<b�a<#�a<V�a<Lya<wma<ba<�Xa<ZQa<Ma<FLa<wNa<Ta<!\a<Yfa<vqa<
}a<��a<E�a<ɘa<]�a<��a<�a<�a<T�a<5�a<��a<0�a<�~a<za<�wa<�va<�wa<jza<s~a<y�a<��a<Z�a<��a<��a<b�a<�a<~�a<�a<�va<�ja<&^a<�Qa<�Fa<I=a<b6a<�2a<�2a<�5a<�;a<?Da<�Na<�Ya<6ea<oa<@xa<�~a<��a<�a<��a<Za<+za<ta<�ma<�ga<�ba<j_a<�]a<^a< `a<�ca<�ha<xna<ta<+ya<�|a<i~a<�}a<2za<Sta<�ka<�aa<�Ua<�Ia<�>a<g4a<�,a<\'a<�%a<'a<�+a<�3a<�=a<Ia<�Ta<�  �  M[a<Yga<�qa<]ya<�~a<�a<B�a<Va<�{a<�wa</sa<.oa<�ka<#ja<�ia<<ka<na<Dra<$wa<O|a<5�a<�a<S�a<r�a< �a<�a<lxa<�na<�ba<�Va</Ja<�>a<�4a<".a<h*a<:*a<�-a<�4a<�>a<�Ja<wXa<_fa<�sa<�a<�a<��a<��a<Әa<�a<�a<ēa<��a<-�a<�a<��a<��a<i�a<Èa<x�a<?�a<��a<�a<Ӡa<i�a<��a<y�a<(�a<3�a<��a<�a<�|a<�oa<vca<�Wa<�Na<�Ha<bEa<�Ea<%Ja<vQa<|[a<�ga<�ta<́a<9�a<��a<��a<��a<��a<v�a<�a<�a<��a<��a<��a<ʕa<A�a<�a<��a<Ŕa<4�a<��a<:�a<�a<��a<+�a<{�a<��a<ҥa<��a<��a<�a<-|a<oa<rba<cWa<�Na<TIa<Ga<�Ha<�Ma<�Ua<�`a<ma<�ya<��a<}�a<c�a<ޣa<ʨa<�a<��a<^�a<��a<ʟa<�a<y�a<͒a<r�a<��a<x�a<Òa<V�a<��a<$�a<d�a<��a<,�a<��a<��a<Ξa<q�a<ҋa<ra<Kra<(ea<�Xa<NNa<�Fa<�Aa<�@a<�Ca<~Ia<GRa<}]a<�ia<�va<�a<Ía<��a<Ԝa<x�a<?�a<�a<��a<Зa<{�a<4�a<e�a<��a<#�a<L�a<�a<N�a<��a<b�a<R�a<Œa<�a<&�a<O�a<��a<�a<�}a<�qa<�da<�Va<8Ia<�<a<�2a<�+a<�'a<c'a<�*a<g1a<�:a<RFa<�Ra<*_a<�ja<,ua<+}a<��a<M�a<|�a<��a<�a<#{a<va</qa<�la<ja<xha<�ha<rja<�ma<�qa< va<eza<~a<7�a<S�a<8~a<Qya<�qa<�ga<&\a<9Oa<Ba<j5a<[*a<�!a<ca<Da<a<A!a<�)a<f4a<Aa<;Na<�  �  �Va<!da<koa<xxa<�~a<p�a<܃a<�a<��a<?}a<�ya<^va<�sa<Yra<ra<^sa<�ua<Yya<g}a<Áa<��a<v�a<��a<��a<�a<�~a<va<ka<`^a<Qa<�Ca<w7a<-a<�%a<�!a<q!a<W%a<�,a<@7a<Da<�Ra<kaa<�oa<}a<I�a<�a<)�a<��a<ۛa<��a<��a<ەa<��a<A�a<��a< �a<��a<ɐa<�a<�a<��a<$�a<ߤa<b�a<�a<"�a<ȡa<��a<�a<�a<�wa<-ja<�\a<�Pa<�Fa<�?a<�<a<C=a<�Aa<{Ia<YTa<aa<"oa<,}a<��a<}�a<2�a<`�a<��a<��a<H�a<@�a<��a<&�a<��a<S�a<V�a<a�a<�a<��a<t�a<�a<��a<˪a<{�a<�a<��a<תa<�a<w�a<��a<Ʉa<wa<�ha<p[a<�Oa<�Fa<�@a<M>a</@a<jEa<ANa<�Ya<�fa<�ta<`�a<E�a<?�a<��a<��a<<�a<H�a<��a<L�a<s�a<p�a<��a<��a<��a<�a<��a<]�a<m�a<ߠa<��a<�a<��a<��a<��a<��a<��a<�a<Y�a<�za<�la<�^a<�Qa<qFa<>a<P9a<8a<;a<JAa<�Ja<�Va<�ca<�qa<�~a<�a<ϔa<P�a<��a<�a<آa<}�a<�a<f�a<��a<��a<��a<l�a<��a<$�a<��a<t�a<b�a<��a<іa<�a<�a<��a<T�a<؅a<�za<na<�_a<�Pa<fBa<~5a<�*a<#a<�a<�a<N"a<m)a<�3a<�?a<Ma<�Za<jga<�ra<�{a<t�a<C�a<��a<Ɇa<B�a<�a<4|a<6xa<�ta<ra<�pa<�pa<Cra<�ta<'xa<�{a<Ma<��a<�a<ׁa<�~a<�xa<�oa<�da<�Wa<Ja<�;a<i.a<�"a<�a<�a<ua<wa<�a<�!a<`-a<�:a<�Ha<�  �  `Ta<ba<na<�wa<�~a<U�a<M�a<�a<e�a<�a<�}a<�za<�xa<Pwa<9wa<Rxa<�za<�}a<s�a<8�a<Q�a<��a<��a<B�a<݄a<�}a<�ta<�ha<�[a<�Ma<�?a<�2a<(a<P a<Ta<a<�a<['a<V2a<�?a<�Na<3^a<rma<I{a<4�a<��a<��a<Ûa<��a<Z�a<��a<��a<.�a<�a<v�a<�a<ȓa<��a<��a<d�a<w�a<V�a<S�a<0�a<�a<��a<M�a<��a<%�a<��a<�ta<gfa<LXa<�Ka<�Aa<�:a<G7a<�7a<N<a<ZDa<�Oa<�\a<ka<Jza<p�a<�a<>�a<
�a<T�a<��a<E�a<ͭa<X�a<,�a<��a<<�a<G�a<��a<�a<�a<�a<=�a<��a<��a<��a<_�a<�a<��a<_�a<:�a<��a<G�a<�sa<�da<�Va<�Ja<8Aa<Y;a<9a<�:a<@a<7Ia<�Ta<�ba<Cqa<�a<@�a<�a<7�a<��a<"�a<��a<&�a<�a<�a<��a<8�a<x�a<��a<�a<��a<M�a<ߡa<�a<�a<��a<	�a<۫a<m�a<U�a<��a<��a<9�a<'xa<Eia<}Za<�La<XAa<�8a<�3a<�2a<�5a<<a<�Ea<-Ra<$`a<{na<�|a<�a<��a<˛a<Z�a<.�a<��a<�a< �a<>�a<4�a<n�a<k�a<x�a<��a<�a<y�a<��a<O�a<��a<E�a<��a<G�a<i�a<ٍa<҄a<>ya<�ka<�\a<-Ma<>a<�0a<g%a<�a<xa<Ja<�a<L$a<�.a<t;a<xIa<�Wa<5ea<qa<�za<�a<ކa<��a<ƈa<Άa<݃a<9�a<�|a<iya<wa<�ua<�ua<*wa<fya<I|a<ta<�a<��a<l�a<ʂa<�~a<�wa<�na<�ba<iUa<�Fa<�7a<�)a<�a<<a<la<+a<a<�a<�a<�(a<�6a<�Ea<�  �  QSa<Eaa<�ma<~wa<�~a<��a<��a<�a<m�a<�a<a<a|a<]za<�xa<�xa<za<\|a<a<��a<c�a<O�a<O�a<F�a<{�a<ބa<�}a<�sa<ha<uZa<)La<D>a<01a<p&a<�a<?a<�a<a<�%a<�0a<?>a<qMa<�\a<|la<�za<��a<q�a<��a<�a<�a<Z�a<�a<�a<~�a<��a<2�a<��a<t�a<f�a<c�a<��a<��a<j�a<Q�a<Ωa<N�a<��a<+�a<=�a<v�a<Ɓa<�sa<ea<�Va<AJa<�?a<�8a<%5a<�5a<�:a<�Ba<Na<�[a<(ja<ya<��a<K�a<��a< �a<��a<6�a<�a<ˮa<z�a<c�a<I�a<��a< �a<I�a<��a<6�a<��a<��a<�a<��a<��a<ΰa<(�a<�a<'�a<Ϛa<ݎa<@�a<Wra<�ca<yUa<>Ia<�?a<_9a<�6a<�8a<�>a<�Ga<zSa<saa<�oa<�~a<h�a<s�a<��a<�a<`�a<�a<�a<�a<S�a<Ǧa<��a<0�a<K�a<Ǟa<E�a<
�a<6�a<'�a<;�a<��a<٬a<"�a<��a<V�a<z�a<�a<P�a<�va<�ga<=Ya<YKa<�?a<7a<�1a<�0a<�3a<�:a<kDa<�Pa<�^a<Ama<�{a<b�a<e�a<��a<s�a<V�a<	�a<�a<�a<u�a<��a<%�a<'�a< �a<W�a<��a<9�a<�a<��a<˘a<D�a<Y�a<z�a<��a<��a<��a<�xa<�ja<h[a<�Ka<�<a</a<�#a<�a<Wa<.a<=a<�"a<I-a<3:a<!Ha<sVa<Hda<|pa<�za<�a<�a<9�a<��a<ˇa<��a<p�a<�}a<){a<�xa<�wa<�wa<�xa<�za<�}a<��a<'�a<�a<ڄa<�a<�~a<�wa<+na<ba<bTa<fEa<�6a<t(a<:a<�a<sa<�	a<
a<�a<Ba<K'a<5a<;Da<�  �  `Ta<ba<na<�wa<�~a<U�a<M�a<�a<e�a<�a<�}a<�za<�xa<Pwa<9wa<Rxa<�za<�}a<s�a<8�a<Q�a<��a<��a<B�a<݄a<�}a<�ta<�ha<�[a<�Ma<�?a<�2a<(a<P a<Ta<a<�a<['a<V2a<�?a<�Na<3^a<rma<I{a<4�a<��a<��a<Ûa<��a<Z�a<��a<��a<.�a<�a<v�a<�a<ȓa<��a<��a<d�a<w�a<V�a<S�a<0�a<�a<��a<M�a<��a<%�a<��a<�ta<gfa<LXa<�Ka<�Aa<�:a<G7a<�7a<N<a<ZDa<�Oa<�\a<ka<Jza<p�a<�a<>�a<
�a<T�a<��a<E�a<ͭa<X�a<,�a<��a<<�a<G�a<��a<�a<�a<�a<=�a<��a<��a<��a<_�a<�a<��a<_�a<:�a<��a<G�a<�sa<�da<�Va<�Ja<8Aa<Y;a<9a<�:a<@a<7Ia<�Ta<�ba<Cqa<�a<@�a<�a<7�a<��a<"�a<��a<&�a<�a<�a<��a<8�a<x�a<��a<�a<��a<M�a<ߡa<�a<�a<��a<	�a<۫a<m�a<U�a<��a<��a<9�a<'xa<Eia<}Za<�La<XAa<�8a<�3a<�2a<�5a<<a<�Ea<-Ra<$`a<{na<�|a<�a<��a<˛a<Z�a<.�a<��a<�a< �a<>�a<4�a<n�a<k�a<x�a<��a<�a<y�a<��a<O�a<��a<E�a<��a<G�a<i�a<ٍa<҄a<>ya<�ka<�\a<-Ma<>a<�0a<g%a<�a<xa<Ja<�a<L$a<�.a<t;a<xIa<�Wa<5ea<qa<�za<�a<ކa<��a<ƈa<Άa<݃a<9�a<�|a<iya<wa<�ua<�ua<*wa<fya<I|a<ta<�a<��a<l�a<ʂa<�~a<�wa<�na<�ba<iUa<�Fa<�7a<�)a<�a<<a<la<+a<a<�a<�a<�(a<�6a<�Ea<�  �  �Va<!da<koa<xxa<�~a<p�a<܃a<�a<��a<?}a<�ya<^va<�sa<Yra<ra<^sa<�ua<Yya<g}a<Áa<��a<v�a<��a<��a<�a<�~a<va<ka<`^a<Qa<�Ca<w7a<-a<�%a<�!a<q!a<W%a<�,a<@7a<Da<�Ra<kaa<�oa<}a<I�a<�a<)�a<��a<ۛa<��a<��a<ەa<��a<A�a<��a< �a<��a<ɐa<�a<�a<��a<$�a<ߤa<b�a<�a<"�a<ȡa<��a<�a<�a<�wa<-ja<�\a<�Pa<�Fa<�?a<�<a<C=a<�Aa<{Ia<YTa<aa<"oa<,}a<��a<}�a<2�a<`�a<��a<��a<H�a<@�a<��a<&�a<��a<S�a<V�a<a�a<�a<��a<t�a<�a<��a<˪a<{�a<�a<��a<תa<�a<w�a<��a<Ʉa<wa<�ha<p[a<�Oa<�Fa<�@a<M>a</@a<jEa<ANa<�Ya<�fa<�ta<`�a<E�a<?�a<��a<��a<<�a<H�a<��a<L�a<s�a<p�a<��a<��a<��a<�a<��a<]�a<m�a<ߠa<��a<�a<��a<��a<��a<��a<��a<�a<Y�a<�za<�la<�^a<�Qa<qFa<>a<P9a<8a<;a<JAa<�Ja<�Va<�ca<�qa<�~a<�a<ϔa<P�a<��a<�a<آa<}�a<�a<f�a<��a<��a<��a<l�a<��a<$�a<��a<t�a<b�a<��a<іa<�a<�a<��a<T�a<؅a<�za<na<�_a<�Pa<fBa<~5a<�*a<#a<�a<�a<N"a<m)a<�3a<�?a<Ma<�Za<jga<�ra<�{a<t�a<C�a<��a<Ɇa<B�a<�a<4|a<6xa<�ta<ra<�pa<�pa<Cra<�ta<'xa<�{a<Ma<��a<�a<ׁa<�~a<�xa<�oa<�da<�Wa<Ja<�;a<i.a<�"a<�a<�a<ua<wa<�a<�!a<`-a<�:a<�Ha<�  �  M[a<Yga<�qa<]ya<�~a<�a<B�a<Va<�{a<�wa</sa<.oa<�ka<#ja<�ia<<ka<na<Dra<$wa<O|a<5�a<�a<S�a<r�a< �a<�a<lxa<�na<�ba<�Va</Ja<�>a<�4a<".a<h*a<:*a<�-a<�4a<�>a<�Ja<wXa<_fa<�sa<�a<�a<��a<��a<Әa<�a<�a<ēa<��a<-�a<�a<��a<��a<i�a<Èa<x�a<?�a<��a<�a<Ӡa<i�a<��a<y�a<(�a<3�a<��a<�a<�|a<�oa<vca<�Wa<�Na<�Ha<bEa<�Ea<%Ja<vQa<|[a<�ga<�ta<́a<9�a<��a<��a<��a<��a<v�a<�a<�a<��a<��a<��a<ʕa<A�a<�a<��a<Ŕa<4�a<��a<:�a<�a<��a<+�a<{�a<��a<ҥa<��a<��a<�a<-|a<oa<rba<cWa<�Na<TIa<Ga<�Ha<�Ma<�Ua<�`a<ma<�ya<��a<}�a<c�a<ޣa<ʨa<�a<��a<^�a<��a<ʟa<�a<y�a<͒a<r�a<��a<x�a<Òa<V�a<��a<$�a<d�a<��a<,�a<��a<��a<Ξa<q�a<ҋa<ra<Kra<(ea<�Xa<NNa<�Fa<�Aa<�@a<�Ca<~Ia<GRa<}]a<�ia<�va<�a<Ía<��a<Ԝa<x�a<?�a<�a<��a<Зa<{�a<4�a<e�a<��a<#�a<L�a<�a<N�a<��a<b�a<R�a<Œa<�a<&�a<O�a<��a<�a<�}a<�qa<�da<�Va<8Ia<�<a<�2a<�+a<�'a<c'a<�*a<g1a<�:a<RFa<�Ra<*_a<�ja<,ua<+}a<��a<M�a<|�a<��a<�a<#{a<va</qa<�la<ja<xha<�ha<rja<�ma<�qa< va<eza<~a<7�a<S�a<8~a<Qya<�qa<�ga<&\a<9Oa<Ba<j5a<[*a<�!a<ca<Da<a<A!a<�)a<f4a<Aa<;Na<�  �  �`a<Nka<.ta<qza<B~a<Wa<�}a<�za<�ua<6pa<�ja<�ea<�aa<}_a<-_a<�`a<da<�ha<�na<,ua<S{a<��a<Y�a<�a<	�a<��a<^{a<�ra<�ha<�]a<~Ra<�Ga<R?a<�8a<�5a<�5a<�8a<a?a<wHa<�Sa<`a<�la<�xa<r�a<A�a<*�a<ߕa<��a<!�a<ˑa<)�a<'�a<)�a<a<#|a<{a<�{a<8~a<��a<�a<��a<2�a<i�a<u�a<��a<��a<��a<3�a<��a<ˍa<
�a<bwa<2la<�aa<hYa<`Sa<�Pa<'Qa<�Ta<�[a<�da<*pa<�{a<؇a<��a<�a<(�a<��a<��a<��a<եa<%�a<��a<��a<9�a<��a<��a<v�a<�a<q�a<��a<��a<��a<��a<�a<��a<��a<�a<��a<��a<��a<p�a<ɂa<�va<�ka<raa<�Ya<PTa<�Ra<�Sa<�Xa<`a<�ia<ua<��a<P�a<t�a<�a<�a<k�a<"�a<V�a<��a<P�a<g�a<L�a<܌a<��a<Ʌa<�a<΅a<��a<�a<:�a<��a<��a<<�a</�a<8�a<|�a<C�a<b�a<#�a<V�a<Lya<wma<ba<�Xa<ZQa<Ma<FLa<wNa<Ta<!\a<Yfa<vqa<
}a<��a<E�a<ɘa<]�a<��a<�a<�a<T�a<5�a<��a<0�a<�~a<za<�wa<�va<�wa<jza<s~a<y�a<��a<Z�a<��a<��a<b�a<�a<~�a<�a<�va<�ja<&^a<�Qa<�Fa<I=a<b6a<�2a<�2a<�5a<�;a<?Da<�Na<�Ya<6ea<oa<@xa<�~a<��a<�a<��a<Za<+za<ta<�ma<�ga<�ba<j_a<�]a<^a< `a<�ca<�ha<xna<ta<+ya<�|a<i~a<�}a<2za<Sta<�ka<�aa<�Ua<�Ia<�>a<g4a<�,a<\'a<�%a<'a<�+a<�3a<�=a<Ia<�Ta<�  �  ga<�oa<
wa<�{a<�}a<�|a<�ya<�ta<ona<bga<v`a<dZa<�Ua<�Ra<qRa<(Ta<"Xa<�]a<�da<�la<_ta<H{a<��a<�a<�a<�a<�~a<�wa<^oa<�ea<�[a<�Ra<Ka<Ea<�Ba<�Ba<�Ea<�Ka<�Sa<�]a<�ha<ta<�~a<��a<��a<ݒa<��a<��a<q�a<��a<j�a<�~a<�xa<�sa<�oa<Yna<oa<�qa<wa<�}a<*�a<J�a<��a<��a<r�a<�a<�a<I�a<ښa<C�a<'�a<�a<va<�la<pea<,`a<�]a<)^a<�aa<�ga<�oa<�ya<3�a<��a<їa<�a<ڤa<��a<��a<#�a<��a<V�a<D�a<�a<n�a<�a<A|a<�za<[{a<Q~a<7�a<��a<��a<�a<�a<`�a<�a<A�a<��a<��a<��a<v�a<~�a<�a<�ua<�la<�ea<;aa<�_a<�`a< ea<�ka<Qta<A~a<��a<��a<�a<�a<(�a<ԧa<��a<>�a<؝a<�a<��a<3�a<��a<~|a<0ya<2xa<]ya<�|a<��a<\�a<}�a<��a<Ȝa<x�a<+�a<W�a<ʡa<��a<�a<�a<��a<�va<�la<gda<�]a<Za<CYa<M[a<8`a<kga<_pa<Hza<Y�a<��a<X�a<�a<�a<p�a<�a<p�a<�a<w�a<^�a<�ya<sa<�ma<�ja<�ia<Wka<�na<�sa<za<��a<�a<�a<��a<�a<��a<��a<�a<0|a<�qa<�fa<�[a<�Qa<OIa<-Ca<�?a<�?a<IBa<�Ga<6Oa<gXa<-ba<�ka<�ta<�{a<��a<��a<8�a<-a<za<^sa<�ka<da<]a<+Wa<Sa< Qa<fQa<Ta<�Xa<�^a<xea<�la<7sa<mxa<�{a<�|a<:{a<�va<0pa<�ga<�]a<Sa<�Ha<�?a<�8a<D4a<�2a<4a<f8a<6?a<Ha<ERa<�\a<�  �  uma<�ta<�ya<�|a<�|a<@za<]ua<jna<afa<�]a<aUa<Na<�Ha<wEa<�Da<�Fa<0Ka<�Qa<%Za<bca<�la<Gua<�|a<��a<f�a<_�a<�a<�|a<$va<Tna<fa<2^a<rWa<�Ra<TPa<qPa<?Sa<PXa<�_a<|ha<!ra<�{a<b�a<��a<��a<@�a<�a<b�a<M�a<��a<�|a<�ta<3ma<�fa<�ba<�`a<raa<�da<7ja<�qa<�za<��a<̍a<5�a<��a<G�a<6�a<0�a<Ξa<��a<��a<<�a<��a<�xa<#ra<�ma<�ka<�ka<oa<1ta<�{a<��a<��a<��a<(�a< �a<a�a<Y�a<x�a<I�a<��a<Ȓa<!�a<^�a<}ya<sa<�na<ma<�ma<;qa<�va<I~a<��a<ۏa<J�a<��a<�a<�a<��a<=�a<��a<��a<�a<��a<�a<ya<�ra<oa<pma<�na<$ra<�wa<ua<�a<ʐa<�a<�a<��a<�a<�a<�a<Ǟa<n�a<��a<�a<}a<Qua<roa<�ka<�ja<la<�oa<�ua<�}a<-�a<ˎa<Ėa<k�a<͡a<գa<�a<�a<<�a<��a<�a<��a<\xa<�pa<Lka<�ga<ga<�ha<ma<bsa<{a<��a<�a<y�a<��a<*�a<u�a<לa<Ҙa<M�a<�a<ڀa<>wa<;na<`fa<�`a<6]a<U\a<^a<ba<>ha<�oa<�wa<�a<��a<"�a<�a<��a<x�a<�a<�a<Vya<�oa<\fa<�]a<Va<�Pa<�Ma<cMa<�Oa<"Ta<�Za<�ba<�ja<�ra<�ya<6a<�a<s�a<
�a<U{a<Ita<�ka<�ba<wYa<#Qa<EJa<�Ea<wCa<�Ca<�Fa<La<[Sa<�[a<ada<�la<�sa<�xa<�{a<|a<�ya<�ta<�ma<�ea<�\a<�Sa<La<�Ea<	Ba<�@a<�Aa<�Ea<rKa<;Sa<\a<ea<�  �  �sa<ya<z|a<r}a<�{a<Pwa<wpa<�ga<^a<�Sa<.Ja<�Aa<~;a<�7a<�6a<9a<7>a<�Ea<9Oa<�Ya<�da<(oa<xa<4a<��a<��a<�a<Ła<�|a<�va<�oa<�ia<�ca<�_a<�]a<^a<�`a<2ea<�ka<sa<+{a<�a<�a<o�a<��a<e�a<_�a<a<ޅa<r}a<�sa<pja<�aa<\Za<QUa<�Ra<�Sa<5Wa<�]a<%fa<kpa<k{a<��a<��a<$�a<z�a<'�a<�a<a�a<v�a<˘a<�a<�a<{�a<�~a<	{a<0ya<�ya<3|a<׀a<��a<�a<��a<{�a<0�a</�a<ߧa<ۦa<<�a<��a<Ȕa<�a<��a<�va<wma<.fa<9aa<1_a<
`a<�ca<eja<�ra<�|a<_�a<��a<��a<�a<ݦa<%�a<��a<��a<Ƞa<R�a<�a<ŋa<:�a<�a<d|a< {a<�{a<)a<)�a<z�a<��a<Řa<5�a<:�a<R�a<��a<֥a<�a<��a<�a<��a<|a<�qa<
ia<Bba<�]a<�\a<>^a<�ba<�ia<�ra<�|a<�a<��a<�a<S�a<$�a<b�a<�a<�a<i�a<m�a<�a<��a<Q}a<exa<lua<�ta<Hva<�ya<Aa<��a<��a<^�a<-�a<F�a<@�a<��a<6�a<2�a<ߌa<��a<�wa<�la<�ba<�Ya<GSa<aOa<�Na<�Pa<iUa<w\a<@ea<�na<uxa<�a<K�a<L�a<��a<]�a<s�a<`�a<��a<�xa<�pa<Bia<�ba<^a<][a<�Za<�\a<�`a<;fa<�la<{sa<�ya<�~a<f�a<��a<��a<�}a<wa<Una<+da<NYa<�Na< Ea<i=a<8a<�5a<6a<�9a<�?a<Ha<�Qa<�[a<�ea<�na<�ua<�za<�|a<|a<�xa<�sa<Tma<fa<�^a<%Xa<�Ra<fOa<9Na<7Oa<�Ra<�Wa<=^a<�ea<ma<�  �  xya<}a<�~a<�}a<cza<]ta<�ka<�aa<Va<�Ja<�?a<36a</a<�*a<�)a<-,a<�1a<U:a<�Da<�Pa<*]a<;ia<�sa<�|a<ła<��a<��a<$�a<�a</~a< ya<�sa<Woa<la<�ja<�ja<�la<�pa<Hva<�|a<^�a<ǉa<@�a<֒a<w�a<:�a<��a<3�a<��a<�va<vka<�`a<�Va<|Na<�Ha<�Ea<�Fa<pJa<�Qa<[a<�fa<�ra<�a<:�a<a�a<�a<âa<��a<��a<s�a<V�a<�a<��a<�a<��a<K�a<�a<I�a<`�a<J�a<[�a<D�a<*�a<��a<¦a<�a<�a<�a<ߠa<Иa<�a<��a<�wa<zla<ba<�Ya<[Ta<3Ra<Sa<`Wa<�^a<2ha<xsa<;a<&�a<a<Ξa<j�a<e�a<ժa<��a<S�a<]�a<��a<��a<:�a<؋a<݈a<߇a<��a<.�a<J�a<��a<Z�a<��a<�a<=�a<��a<n�a<��a<'�a<0�a<��a<�~a<�ra<Tga<q]a<�Ua<�Pa<�Oa<WQa<�Va<V^a<`ha<�sa<Ja<��a<��a<��a</�a<Q�a<��a<f�a<o�a<�a<��a<�a<��a<��a<�a<��a<��a<��a<��a<K�a<ٔa<�a<Z�a<��a<�a<r�a<k�a<��a<��a<)|a<�oa<Kca<�Wa<�Ma<�Fa<`Ba<Aa<�Ca<rIa<WQa<p[a<2fa<qqa<�{a<��a<P�a<I�a<�a<��a<[�a<#�a<܀a<Iza<�sa<una<Ija<ha<�ga<ia<:la<�pa<�ua<&{a<�a<��a<>�a<��a</�a<u{a<�ra<�ha<�\a<mPa<�Da<�9a<:1a<0+a<�(a<)a<-a<4a<H=a<DHa<�Sa<m_a<�ia<�ra<ya<�|a<&~a<�|a<gya<\ta<�na<�ha<"ca<�^a<�[a<�Za<�[a<�^a<�ba<Gha<Xna<7ta<�  �  ~a<Q�a<p�a<9~a<6ya<�qa<�ga<\a<MOa<�Ba<X6a<,a<K$a<�a<�a<9!a<J'a<V0a<�;a<Ia<�Va<�ca<
pa<Bza<��a<&�a<��a<��a<هa<��a<��a<�|a<ya<iva<)ua<sua<~wa<�za<�a<ӄa<R�a<p�a<i�a<��a<��a<�a<܍a<�a<|a<pa<Bda<6Xa<�La<Da<�=a<�:a<R;a<�?a<Ga<ZQa<�]a<{ka<Hya<v�a<�a<��a<|�a<��a<�a<y�a<פa<�a<��a<H�a<��a<ݑa<��a<�a<ђa<�a<R�a<��a<��a<ǧa<��a<&�a<��a<o�a<��a<;�a<�a<@}a<8pa<�ca<8Xa<^Oa<mIa<�Fa<�Ga<�La<bTa<�^a<;ka<Lxa<V�a<��a<�a<�a<��a<L�a<��a<Ϊa<V�a<ܢa<%�a<��a<��a<��a<��a<7�a<f�a<ߘa<�a<��a<�a<��a<}�a<J�a<��a<^�a<q�a<"�a<�a<�wa<�ja<^a<<Sa<	Ka<�Ea<5Da<`Fa<�Ka<TTa<Q_a<�ka<�xa<_�a<Ӑa<\�a<c�a<٥a<��a<��a<[�a<U�a<��a<Ėa<c�a<�a<Ìa<"�a<8�a<��a<D�a<o�a<ϛa<��a<��a<h�a<-�a<S�a<��a<��a<�a<va<Qha<�Za<Na<�Ca<�;a<+7a<46a<�8a<�>a<�Ga<�Ra<�^a<6ka<�va<=�a<g�a< �a<�a</�a<a�a<��a<��a<F�a<}a<axa<�ta<�ra<Kra<usa<va<�ya<�}a<��a<(�a<M�a<`�a<_�a<��a<8ya<Ooa<wca<TVa<�Ha<�;a<�/a<�&a<D a<;a<	a<["a<�)a<�3a<@a<�La<�Ya<�ea<�oa<�wa<}a<�a<�a<�}a<Rza<�ua<qa<�la<�ha<�fa<�ea<jfa<�ha<hla<�pa<�ua<Xza<�  �  ��a<܂a<��a<V~a<?xa<uoa<tda<�Wa<�Ia<$<a<M/a<J$a<�a<a<�a<�a<�a<�(a<�4a<�Ba<�Qa<�_a< ma<Exa<E�a<�a<!�a<��a<��a<��a<d�a<<�a<P�a<F~a<h}a<�}a<�a<k�a<��a<��a<��a<��a<��a<��a<��a<�a<q�a<��a<rxa<�ka<�^a<{Qa<�Ea<�;a<H5a<2a<�2a<7a<�>a<Ja<'Wa<�ea<�ta<��a<q�a<�a<.�a<k�a<+�a<��a<��a<0�a<��a<3�a<��a<�a<ژa<.�a<��a<j�a<�a<ߤa<Ĩa<��a<a�a<�a<(�a<ڤa<��a<O�a<څa<?xa<4ja<�\a<�Pa<!Ga<�@a<�=a<L?a<(Da<�La<�Wa<�da<�ra<Հa<�a<��a<�a<��a<u�a<�a<<�a<�a<`�a<z�a<Ԡa<��a<��a<њa<l�a<�a<	�a<��a<J�a<ͪa<!�a<	�a<��a<ڨa<g�a<>�a<ڍa<��a<�ra<Ida<�Va<�Ka<�Ba<K=a<f;a<�=a<�Ca<�La<SXa<�ea<�sa<2�a<Ǎa<]�a<��a<1�a<�a<éa<&�a<M�a<\�a<g�a<��a<a<�a<k�a<G�a<&�a<B�a<��a<#�a<�a<��a<��a<�a<!�a<L�a<��a<ua<^qa<�ba<
Ta<�Fa<~;a<?3a<m.a<q-a<o0a<�6a<k@a<�Ka<"Ya<mfa<;sa<�~a<ևa<��a<��a<:�a<g�a<��a<�a<R�a<��a<�a<�|a<{a<�za<d{a<X}a<P�a<{�a<��a<�a<-�a<#�a<ԅa<�a<Zwa<dla<m_a<TQa<�Ba<�4a<}(a<ca<�a<qa<aa<�a<�!a<�,a<�9a<iGa<Ua<+ba<uma<�va<}a<Āa<<�a<L�a<�~a<L{a<]wa<�sa<�pa<�na<�ma<�na<tpa<�sa<Hwa<D{a<
a<�  �  ȃa<E�a<��a<H~a<twa<na<hba<�Ta<�Fa<$8a<�*a<=a<�a<�a<ga<Ga<�a<�#a<t0a<	?a<3Na<E]a<ka<wa<��a<��a<�a<�a<�a<l�a< �a<a�a<�a<)�a<k�a<��a<z�a<L�a<�a<��a<��a<=�a<��a<�a<�a<��a<x�a<�a<2va<�ha<�Za<EMa<Aa<�6a<�/a<�,a<:-a<�1a<�9a<DEa<�Ra<ba<oqa<_�a<��a<�a<��a<�a<X�a<]�a<r�a<o�a<��a<~�a<Ša<Ϟa<�a<9�a<��a<�a<=�a<��a<ƫa<�a<��a<��a<{�a<M�a<��a<w�a<i�a<�ta<Xfa<*Xa<�Ka<�Aa<{;a<�8a<�9a<�>a<{Ga<Sa<�`a<\oa<!~a<�a</�a<�a<k�a<<�a<d�a<O�a<��a<�a<��a<M�a<��a<��a<�a<d�a<	�a<��a<��a<�a<��a<D�a<s�a<l�a<˨a<��a<ߗa<ϋa<�}a<!oa<I`a<^Ra<uFa<J=a<�7a<6a<j8a<E>a<�Ga<�Sa<�aa<Lpa<�~a<݋a<+�a<
�a<c�a<�a<G�a<k�a<+�a<�a<��a<F�a<��a<�a<��a<4�a<�a<��a<��a<u�a<��a<��a<ͦa<��a<��a<S�a<T�a<5}a<mna<_a<�Oa<Ba<[6a<�-a<)a<(a<+a<�1a<�;a<�Ga<dUa<\ca<�pa<�|a<Նa<;�a<(�a<g�a<C�a<<�a<*�a<F�a<@�a<��a<ʁa<�a<�a<D�a<��a<�a<I�a<a<f�a<ɋa<3�a<(�a<oa<=va<�ja<�\a<Na<�>a<O0a<�#a<"a<Ua<a<�a<�a<�a<((a<u5a<�Ca<iRa<`a<la<�ua<�|a<��a<��a<_�a<��a<�~a<m{a</xa<yua<�sa<sa<�sa<`ua<xa<^{a<�~a<��a<�  �  �}a<�}a<m|a<$ya<�sa<�la<qca<^Ya<wNa<�Ca<�9a<M1a<�*a<'a<�&a<d(a<�-a<-5a<�>a<�Ia<HUa<�`a<fka<�ta<h|a<7�a<ʅa<��a<��a<�a<��a<��a<��a<�a<Y�a<�a<H�a<��a<Q�a<��a<��a<U�a<�a<%�a<�a<]�a<��a<��a<�wa<�ma<�ca<�Ya<`Pa<OIa<�Ca<�Aa<xBa<�Ea<_La<�Ta<]_a<�ja<�va<	�a<Z�a<?�a<%�a<I�a<��a<2�a<֤a<X�a<��a<�a<M�a<�a<A�a<|�a<̜a<��a<Πa<��a<��a<��a<�a<��a<I�a<B�a<��a<�a<�a<{a<8pa<�ea<4\a<�Ta<�Oa<Na<�Na<�Ra<=Ya<�aa<0la<wa<<�a<��a<>�a<�a<��a<��a<>�a<��a<]�a<m�a<�a<}�a<��a<�a<��a<ϝa<�a<ݠa<-�a<��a<c�a<��a<V�a<��a<�a<=�a<��a<5�a<��a<lva<rka<�`a<�Wa<Qa<�La<�Ka<�La<�Qa<�Xa<�aa<la<�va<ˁa<��a<~�a<B�a<]�a<8�a<Q�a<�a<#�a< �a<$�a<a<ؘa<\�a<��a<l�a<��a<p�a<ʜa<��a< �a<��a<��a<	�a<-�a<y�a<͈a<�~a<Bsa<�ga<\a<PQa<�Ha<�Aa<K>a<x=a<A?a<kDa<XKa<�Ta<�^a<�ha<sa<�{a<��a<;�a<(�a<��a<��a<M�a<Ċa<��a<��a<ށa<�a< ~a<�}a<!~a<-a<��a<�a<Y�a<��a<p�a<Ӄa<��a<{a<�sa<�ja<C`a<�Ta<tIa<Y>a<�4a<�,a<V'a<;%a<�%a<)a<N/a<}7a<�Aa<<La<1Wa<waa<�ja<?ra<�wa<�{a< }a<f}a<|a<za<�wa<ua<2sa<�qa<Rqa<�qa<0sa<ua<�wa<:za<P|a<�  �  #}a<�}a<3|a<ya<�sa<�la<da<7Za<tOa<�Da<�:a<~2a<4,a<c(a<�'a<�)a<�.a<j6a<�?a<�Ja<>Va<�aa<la<@ua<�|a<�a<~�a<'�a<?�a<?�a<��a<��a<݀a<�a<=a<�a<�a<^�a<S�a<��a<ڌa<��a<i�a<ܑa<��a<b�a<<�a<!�a<�xa<�na<�da<�Za<�Qa<dJa<XEa<�Ba<�Ca<&Ga<xMa<Va<``a<�ka<owa<��a<Ռa<��a<:�a<�a<��a<��a<"�a<��a<j�a<(�a<�a<��a<#�a<c�a<v�a<l�a<�a<��a< �a<Ǧa<~�a<��a<�a<k�a<�a<t�a<ʆa<�{a<qa<�fa<q]a<&Va<;Qa</Oa<Pa<�Sa<bZa<�ba<ma<xa<�a<e�a<��a<�a<��a<>�a<�a<�a<��a<��a<��a<n�a<C�a<ݜa<X�a<��a<ѝa<ȟa<1�a<��a<��a<�a<�a<e�a<�a<c�a<�a<یa<��a<iwa<Ola<�aa<Ya<SRa<Na<�La<RNa<�Ra<�Ya<�ba<�la<�wa<��a<=�a<˔a<j�a<+�a<�a<٣a<2�a<n�a<��a<;�a<��a<��a<@�a<וa<9�a<��a<q�a<��a<ʝa<k�a<�a<<�a<��a<2�a<��a<>�a<Ba<ta<sha<]a<�Ra<�Ia<QCa<u?a<�>a<�@a<�Ea<�La<�Ua<u_a<�ia<�sa<z|a<�a<Q�a<Ìa<]�a</�a<��a<��a<׆a<��a<��a<_~a<}a<y|a<�|a<~a<�a<ҁa<��a<̈́a<�a<��a<N�a<+{a<%ta<'ka<�`a<�Ua<NJa<l?a<�5a<.a<�(a<K&a<�&a<_*a<s0a<�8a<�Ba<5Ma<Xa< ba<ka<fra<�wa<A{a<�|a<�|a<\{a<(ya<�va<ta<�qa<�pa<%pa<�pa<�qa<ta<�va<Eya<�{a<�  �  c{a<g|a<�{a<ya<ata<�ma<�ea<\a<�Qa<�Ga<U>a<*6a<0a<�,a<�+a<.a<�2a<:a<FCa<�Ma<�Xa<fca<nma<va<�|a<�a<΄a<�a<i�a< �a<��a<�a<_}a<�{a<P{a<�{a<J}a<�a<�a<��a<v�a<��a<�a<�a<�a<��a<؈a<C�a<"za<�pa<4ga<�]a<EUa<Na<}Ia<(Ga<�Ga<YKa<'Qa<�Ya<�ca<fna<�ya<Y�a<�a<.�a<��a<��a<�a<0�a<3�a<@�a<n�a<��a<|�a<ٖa<�a<l�a<��a<�a<ʜa<��a<Ӣa<�a<1�a<�a<ͣa<ԟa<��a<ˑa<{�a<Y~a<�sa<�ia< aa<�Ya<wUa<CSa<ITa<�Wa<^a<wfa<pa<�za<	�a<�a<��a<��a<ţa<��a<�a<:�a<��a<�a<�a<�a<��a<�a<B�a<Șa<�a<_�a< �a<�a<��a<0�a<�a<ɥa<�a<�a<��a<Z�a<v�a<�ya<2oa<iea<�\a<<Va<?Ra<�Pa<�Ra<�Va<}]a<fa<�oa<3za<J�a<��a<��a<ڛa<	�a<<�a<��a<\�a<O�a<�a<&�a<"�a<��a<T�a<Ƒa<m�a<֓a<6�a<��a<f�a<u�a<|�a<k�a</�a<n�a<Q�a<`�a<ڀa<8va<ka<`a<6Va<�Ma<vGa<�Ca<�Ba<�Da<4Ia<EPa<�Xa<"ba<�ka<Sua<�}a<��a<��a<_�a<��a<��a<��a<��a<ۃa<o�a<}a<�za<�xa<�xa<�xa<�za<�|a<�~a<v�a<�a<��a<˂a<�a<�{a<�ta<~la<�ba<Xa<Ma<�Ba<s9a<�1a<�,a<^*a<+a<[.a<4a<9<a<zEa<�Oa<�Ya<�ca<la<�ra<�wa<�za<�{a<{a<\ya<�va<�sa<�pa<-na<�la<la<�la<na<�pa<�sa<�va<�ya<�  �  �xa<rza<|za<�xa<ua<�oa< ha<a_a<�Ua<qLa<�Ca<�;a<%6a<�2a<.2a</4a<�8a<�?a<]Ha<4Ra<�\a<�fa<�oa<�wa<o}a<��a<y�a<ԃa<��a<N�a<j}a<vza<�wa<va<Aua<�ua<xwa<za<�}a<�a<^�a<S�a<v�a<K�a<c�a<��a<ȉa<D�a<�|a<tta<�ka<�ba<�Za<Ta<�Oa<�Ma<)Na<eQa<8Wa<_a<qha<�ra<=}a<0�a<%�a<?�a<��a<�a<=�a<Ԡa<��a<6�a<��a<��a<�a<�a<�a<R�a<�a<P�a<��a<P�a<�a<�a<�a<}�a<h�a<&�a<��a<�a<��a<"�a<cxa<�na<�fa<`a<�[a<�Ya<�Za<�]a<�ca<�ka<�ta<�~a<j�a<��a<f�a<\�a<��a<��a<
�a<��a<�a<��a<%�a<��a<�a<�a<0�a<˒a<i�a<��a<;�a<��a<��a<��a<�a<��a<��a<��a<��a<�a<��a<�}a<�sa<�ja<�ba<F\a<�Xa<GWa<�Xa<�\a<ca<+ka<cta<~a<i�a<�a<�a<K�a<��a<�a<��a<��a<}�a<їa<�a<��a<�a<D�a<��a<��a<?�a<�a<�a<N�a<�a<�a<��a<~�a<p�a<A�a<`�a<��a<�ya<boa<ea<�[a<�Sa<|Ma<Ja<(Ia<�Ja<DOa<�Ua<�]a<�fa<�oa<+xa<�a<��a<��a<Ћa<�a<d�a<o�a<��a<ma<2{a<vwa<�ta<�ra<ira<Gsa<�ta<�wa<�za<�}a<�a<r�a<W�a<�a<�{a<2va<�na<�ea<�[a<�Qa<�Ga< ?a<�7a<3a<�0a<X1a<a4a<�9a<Aa<LJa<�Sa<^]a<Hfa<�ma<�sa<�wa<�ya<�ya<uxa<�ua<`ra<�na<Uka<�ha<�fa< fa<�fa<|ha<6ka<�na<]ra<�ua<�  �  Bua<�wa<2ya<�xa<�ua<kqa<ka<�ca<[a<�Ra<KJa<�Ca<Q>a<);a<�:a<j<a<�@a<'Ga<Oa<Xa<laa<|ja<yra<5ya<�}a<�a<߁a<�a<�~a<]{a<�wa<�sa<�pa<Dna<;ma<�ma<^oa<�ra<�va<�{a<�a<�a<M�a<�a<{�a<��a<�a<�a<J�a<ya<�pa<�ha<�aa<�[a<�Wa<�Ua<�Va<�Ya<&_a<5fa<�na<Mxa<�a<��a<x�a<��a<Ϝa<�a<'�a<ŝa<Қa<��a<�a<ʎa<j�a<
�a<�a<S�a<�a<��a<�a<��a<ޙa<�a<.�a<��a<¢a<��a<��a<��a<^�a<�a<~a<�ua<na<ha<�ca<@ba<�ba<)fa<�ka<�ra<�za<ڃa<��a<��a<e�a<]�a<r�a<��a<��a<I�a<��a<H�a<��a<��a<=�a<��a<E�a<��a<��a<a<��a<*�a<O�a<�a<w�a<b�a<k�a<h�a<��a<Փa<��a<�a<za<bqa<-ja<uda<�`a<�_a<�`a<�da<�ja<�qa<@za<��a<d�a<��a<Ęa<ۜa<*�a<O�a<͝a<ƚa<��a<!�a<j�a<Q�a<+�a<=�a<��a<��a<��a<�a<�a<��a<֕a<�a<u�a<��a<��a<��a<��a<�a<N~a<�ta<cka<�ba<d[a<�Ua<lRa<�Qa<Sa<2Wa<�\a<da<
la<;ta<�{a<�a<�a<�a<��a<ىa<U�a<L�a<d~a<[ya<Eta<�oa<�la<�ja<jja<\ka<�ma<�pa<�ta<�xa<|a<�~a<�a<a<N|a<�wa<Wqa<�ia<�`a<VWa<TNa<VFa<�?a<K;a<X9a<�9a<�<a<�Aa<NHa<vPa<Ya<�aa<\ia<�oa<�ta<�wa<�xa<�wa<ua<Cqa<�la<dha<1da<�`a<�^a<^a<�^a<�`a<da<7ha<�la<>qa<�  �  �pa<�ta<nwa<&xa<�va<�sa<�na<Pha<�`a<�Ya<YRa<La<~Ga<�Da<6Da<�Ea<�Ia<�Oa<�Va<�^a<ga<�na<�ua<,{a<�~a<C�a<�a<�}a<za<�ua<�pa<la<,ha<;ea<�ca<=da<#fa<�ia<�na<|ta<�za<�a<C�a<x�a<�a<Ǎa<��a<�a<;�a<!~a<wa<apa<�ia<�da<aa<�_a<)`a<ca<�ga<�na<qva<�~a<�a<Ԏa</�a<4�a<�a<�a<��a<ߙa<Еa<�a<��a<ʆa<ςa<�a<�~a<�~a<�a<��a<�a<i�a<�a<D�a<��a<��a<ۡa<'�a<r�a<��a<��a<v�a<��a<T}a<nva<�pa<Uma<�ka<�la<qoa<<ta<�za<'�a<̉a<��a<E�a<��a<��a</�a<�a<��a<��a<3�a<��a<8�a<^�a<d�a<��a<ˀa<h�a<��a<�a<&�a<{�a<ؖa<��a<F�a<��a<�a<g�a<Ŝa<R�a<��a<߈a<�a<rya<�ra<�ma<`ja<Tia<�ja<�ma<sa<�ya<�a<��a<܏a<�a<��a<��a<m�a<P�a<N�a<�a<ܐa<,�a<��a<�a<!}a<�za<Sza<E{a<~a<ځa<��a<͋a<��a<ڔa<՗a<8�a<��a<��a<2�a<�a<m�a<�za<�ra<�ja<da<_a< \a<([a<�\a<�_a<ea<�ka<Tra<xya<�a<քa<��a<$�a<ɉa<p�a<q�a<K~a<Xxa<ra<Fla<bga<�ca<�aa<aa<Eba<%ea< ia<�ma<�ra<Iwa<�za<w}a<$~a<�|a<�ya<Xta<�ma<%fa<�]a<Va<�Na<�Ha<�Da<�Ba<;Ca<�Ea<IJa<nPa<�Wa<�^a<�fa<�la<Ara<�ua<Zwa<�va<�ta<�pa<�ka<mfa<�`a<\a<Xa<pUa<�Ta<ZUa<�Wa<�[a<�`a<-fa<�ka<�  �  #la<}qa<lua<zwa<�wa<�ua<:ra<4ma<(ga<�`a<�Za<TUa<NQa<�Na<tNa<Pa<�Sa<�Xa<�^a<�ea<�la<�sa<ya<	}a<"a<Fa<�}a< za<$ua<Xoa<Wia<�ca<�^a<m[a<�Ya<�Ya<:\a<G`a<�ea<�la<�sa<M{a<�a<��a<��a<��a<��a<ߋa<E�a<p�a<�}a<�wa<�ra<na<ka<�ia<bja<ma<nqa<Twa< ~a<e�a<��a<��a<(�a<��a<��a<u�a<��a<ŕa<O�a<%�a<ރa<~a<Bya<�ua<Qta<�ta<wa<{a<��a<�a<��a<!�a<Ǚa<+�a<��a<i�a<#�a<��a<,�a<@�a<��a<F�a<ka<�za<�wa<va<�va<Qya<�}a<-�a<��a<7�a<��a<�a<(�a<\�a<��a<
�a<|�a<o�a<G�a<��a</�a<Wa<�za<�wa<mva<Swa<za<]~a<�a<D�a<ːa<�a<��a<��a<V�a< �a<�a<�a<��a<"�a<T�a<ׁa<�{a<vwa<�ta<�sa<�ta<�wa<|a<ʁa<�a<��a<|�a<O�a<��a<�a<q�a<�a<��a<�a<��a<��a<I}a<�wa<Ssa<�pa<�oa<Zqa<ita<ya<�~a<�a<�a<��a<��a<��a<]�a<�a<��a<��a<��a<��a<_za<�sa<�ma<ia<7fa<aea<�fa<{ia<�ma<Hsa<#ya<�~a<��a<Їa<�a<�a<W�a<��a<Xa<�xa<�qa<Oja<�ca<�]a<�Ya<4Wa<�Va<mXa<�[a<�`a<+fa<8la<&ra<3wa<{a<�|a<$}a<T{a<�wa<Vra<�ka<�da<^a<�Wa<�Ra<�Na<!Ma<vMa<�Oa<�Sa<�Xa<�^a<iea<�ka<�pa<�ta<�va<�va<ua<dqa<>la<fa<S_a<�Xa< Sa<]Na<jKa<DJa<HKa<Na<�Ra<~Xa<�^a<�ea<�  �  Pga<�ma<Gsa<�va<]xa<�wa<�ua<�qa<Dma<ha<�ba<^a<
[a<Ya<�Xa<Za<@]a<�aa<�fa<�la<�ra<xa<|a<�~a<�a<Y~a<{a<%va<pa<�ha<�aa<*[a<�Ua<�Qa<zOa<�Oa<Ra<�Va<�\a<�da<ma<�ua<�}a<c�a<��a<f�a<��a<e�a<�a<��a<O�a<�a<{a<�wa<�ta<ta<�ta<�va<�za<�a<ƅa<�a<��a<��a<Кa<�a<��a<	�a<�a<��a<Ɋa<H�a< |a<=ua<�oa<�ka<ja<�ja<!ma<�qa<�wa<\a<�a<�a<͕a<}�a<��a<��a<ˡa<�a<{�a<��a<��a</�a<P�a<M�a<r�a<i�a<�a<�a<Ԇa<}�a<�a<x�a<��a<��a<c�a<E�a<3�a<�a<��a<��a<>�a<��a<�|a<2va<�pa<vma<,la<ma<9pa<'ua<�{a<�a<��a<�a<[�a<v�a<��a<�a<�a<`�a<W�a<@�a<��a<�a<%�a<4�a<�~a<�}a<�~a<H�a<�a<ʉa<)�a<e�a<�a<`�a<f�a<o�a<��a<��a<ܒa<�a<�a<Q|a<�ta<Cna<nia<zfa<�ea<8ga<�ja<pa<�va<�}a<a�a<<�a<��a<�a<1�a<V�a<~�a<Ԓa<�a<*�a<�a<|a<�va<�ra<pa<�oa<tpa< sa<�va<�za<�a<S�a<��a<y�a<B�a<�a<�a<��a<{a<Fsa<�ja<�ba<�Za<CTa<�Oa<�La<�La<zNa<LRa<�Wa<�^a<�ea<�la<8sa<Sxa<�{a<j}a<�|a<�za<�va<�qa<�ka<�ea<�`a<)\a<�Xa<{Wa<�Wa<uYa<�\a<9aa<_fa<�ka<pa<Rta<�va<�wa<`va< sa<�ma<�ga<�_a<2Xa<�Pa<�Ia<�Da<9Aa<@a<Aa<VDa<pIa<)Pa<�Wa<�_a<�  �  �ba<uja<%qa<�ua<�xa<�ya<�xa<xva<�ra<�na<�ja<�fa<�ca<`ba<Eba<aca<	fa<�ia<lna<^sa<xa<A|a<
a<h�a<�a<"}a<�xa<mra<ka<�ba<�Za<�Ra<�La<9Ha<�Ea<Fa<�Ha<�Ma<�Ta<]a<|fa<*pa<bya<w�a<.�a<�a<ۏa<��a<ԏa<��a<,�a<��a<��a<�a<~a<_}a<~a<�a<��a<�a<�a<�a<�a<Қa<!�a<�a<��a<j�a<'�a<f�a<y�a<�|a<�ta<�la<�fa<dba<�`a<�`a<�ca<ia<�oa<xa<ڀa<։a<�a<��a<O�a<��a<=�a<��a<��a<$�a<��a<��a<f�a<�a<��a<܉a<@�a<�a<2�a<5�a<Зa<�a</�a<�a<S�a<�a<b�a<�a<��a<5�a<��a<�}a<ua<�ma<�ga<�ca<�ba<�ca<ga<�la<�sa<|a<Ԅa<p�a<�a<S�a<��a<b�a<�a<��a<ܞa<ǚa<]�a<��a<u�a<)�a<�a<k�a<��a<�a<=�a<F�a<��a<��a<2�a<P�a<��a<��a<Q�a<�a<%�a<�a<~a<ua<�la<�ea<`a<�\a</\a<�]a<�aa<�ga<oa<fwa<�a<��a<юa<D�a<��a<P�a<��a<��a<͒a<�a<�a<�a<ya<|a<�ya<ya<�ya<�{a<�~a<9�a<Ѕa<G�a<Ћa<ʌa<c�a<��a<N�a<�~a<�va<�ma<Zda<�Za<fRa<|Ka<Fa<gCa<Ca<Ea<�Ia<�Oa<JWa<{_a<�ga<Yoa<�ua<�za<m}a<k~a<I}a<�za<�va<)ra<Rma<�ha<�da<$ba<�`a<�`a<vba<:ea<�ha<Dma<Lqa<"ua<�wa<�xa<Exa<�ua<qa<�ja<ca<TZa<aQa<�Ha<hAa<�;a<�7a<w6a<�7a<6;a<�@a<(Ha<�Pa<�Ya<�  �  �^a<�ga<Hoa<ua<7ya<!{a<e{a<za<�wa<Zta<qa<na<�ka<lja<.ja<|ka<�ma<�pa<�ta<�xa<�|a<�a<b�a<|�a<�a<|a<�va<Eoa<�fa<�]a<yTa<'La<!Ea<@a<�=a<�=a<c@a<�Ea<XMa<Va<�`a<dka<�ua<�~a<��a<��a<��a<k�a<��a<v�a<I�a<��a<ǉa<g�a<��a<W�a<	�a<�a<�a<ˎa<�a<F�a<��a<ӝa<%�a<͞a<c�a<�a<őa<��a<ǀa<Xwa<na<�ea<�^a<6Za<Xa<�Xa<�[a<2aa<�ha<�qa<�{a<X�a<��a<ɖa<�a<��a<5�a<�a<ӣa<}�a<T�a<ٚa<v�a<��a<ϒa<Αa<K�a<�a<v�a<ҙa<t�a<��a<ڣa<��a<إa<e�a<��a<H�a<�a<+�a<��a<�wa<jna<=fa<�_a<�[a<Za<D[a<�^a<ea<�la<va<�a<G�a<�a<v�a<��a<��a<J�a<.�a<h�a<��a<�a<1�a<��a<�a<�a<W�a<�a<��a<]�a<��a<�a<,�a<��a<��a<�a<��a<=�a<�a<��a<��a<�xa<�na<�ea<�]a<�Wa<�Ta<�Sa<�Ua<�Ya<o`a<�ha<�qa<'{a<.�a<U�a<��a<U�a<�a<��a<n�a<��a<#�a<��a<��a<چa<��a<Ӂa<	�a<��a<�a<d�a<:�a<�a<X�a<юa<ώa<,�a<�a<Ճa<||a<Vsa<Fia<�^a<vTa<@Ka<�Ca<�=a<�:a<�:a<�<a<�Aa<�Ha<�Pa<)Za<[ca<la<�sa<Yya<k}a<ba<�a<�}a<#{a<�wa<�sa<�oa<sla<@ja<�ha<�ha<Hja<}la<�oa<�ra<,va<�xa<hza<_za<�xa<�ta<Toa<�ga<�^a<bUa<yKa<Ba<�9a<w3a<u/a<�-a<A/a<3a<^9a<pAa<�Ja<�Ta<�  �  C[a<ea<�ma<�ta<{ya<L|a<b}a<�|a<;{a<�xa< va<qsa<cqa<npa<@pa<gqa<Esa<>va<�ya<�|a<�a<�a<<�a<a�a<�a<?{a<�ta<�la<Nca<}Ya<�Oa<�Fa<;?a<:a<87a<'7a<J:a<�?a<�Ga<�Qa<R\a<�ga<�ra<�|a<Y�a<J�a<��a<�a<�a<��a<:�a<�a<��a<��a<��a<s�a<$�a<ݍa<��a<�a<s�a<H�a<*�a<#�a< a<N�a<>�a<Ζa<��a<ކa<!}a<�ra<ia<F`a<�Xa<&Ta<�Qa<+Ra<�Ua<6[a<lca<�la<Ewa<ցa<�a<הa<2�a<��a<��a<��a<H�a<�a<u�a<{�a<Üa<3�a<��a<�a<X�a<��a<��a<۞a<��a<Ťa<��a<��a<�a<��a<A�a<��a<��a< �a<�}a<sa<Fia<�`a<�Ya<zUa<�Sa<Ua<�Xa<Q_a<�ga<Tqa<�{a<�a<��a<̗a<]�a<��a<u�a<,�a<�a<9�a<)�a<"�a<�a<��a<�a<j�a<�a<S�a<��a<^�a</�a<��a<�a<��a<��a<ٞa<p�a<6�a<T�a<Ga<�ta<	ja<q`a<�Wa<�Qa<7Na<9Ma<gOa<�Sa<�Za<�ca<:ma<jwa<1�a<�a<n�a<�a<n�a<�a<��a<ʙa<�a<K�a<�a<o�a<��a<�a<#�a<b�a<��a<��a<��a<�a<��a<"�a<l�a<��a<Z�a<��a<Lza<tpa<�ea<\Za<�Oa<�Ea<q=a<�7a<�4a<F4a<�6a<�;a<[Ca<La<�Ua<�_a<Nia<�qa<txa<q}a<#�a<S�a<k�a<�~a<�{a<0xa<ua<	ra<pa<�na<oa<�oa<�qa<�ta<,wa<�ya<�{a<v|a<�{a<ya<qta<�ma<�ea<�[a<yQa<�Fa<�<a<C4a<j-a<C)a<{'a<)a<-a<�3a<@<a<Fa<�Pa<�  �  mYa<�ca<�la<ta<�ya<�|a<�~a<y~a<H}a<P{a<ya<�va<+ua<Qta<Tta<3ua<�va<�ya<�|a<{a<�a<��a<3�a<�a<�a<�za<�sa<ka<Taa<�Va<�La<=Ca<�;a<6a<3a<3a<6a<�;a<#Da<DNa<�Ya<Wea<�pa<i{a<��a<�a<<�a<��a<G�a<a�a<n�a<דa<�a<��a<��a<n�a<)�a<��a<&�a<1�a<l�a<��a<�a<��a<��a<��a<�a<$�a<\�a<;�a<�za<2pa<�ea<�\a<#Ua<�Oa<~Ma<�Ma<rQa<�Wa<�_a<�ia<�ta<�a<R�a<��a<��a<��a<u�a<��a<ۧa<ަa<�a<�a<�a<�a<x�a<�a<A�a<j�a<o�a<�a<��a<ߦa<x�a<�a<˧a<Фa<͟a<�a<$�a<?�a<G{a<Kpa<�ea<�\a<�Ua<;Qa<�Oa<�Pa<�Ta<�[a<Kda<xna<Nya<1�a<�a<�a<��a<�a<�a<M�a<ߦa<G�a<�a<3�a<��a<\�a<�a<�a<әa<�a<�a<j�a<��a<��a<��a<|�a<��a<��a<�a<.�a<ɇa<L}a<ra<ga<�\a<PTa<�Ma< Ja<"Ia<+Ka<	Pa<9Wa<H`a<xja<ua<�a<��a<��a<��a<��a<��a<��a<��a<G�a<<�a<�a<��a<~�a<�a<)�a<6�a<4�a<ʍa<��a<M�a<o�a<��a<*�a<�a<�a<
�a<ya<�na<bca<�Wa<YLa<Ba<�9a<�3a<d0a<0a<�2a<,8a<�?a<
Ia<JSa<�]a<�ga<�pa<�wa<=}a<��a</�a<��a<��a<~a<3{a<Ixa<�ua<�sa<�ra<�ra<�sa<uua<�wa<�ya<|a<k}a<�}a<R|a<*ya<�sa<�la<da<Za<
Oa<Da<�9a<�0a<�)a<%a<i#a<�$a< )a<�/a<�8a<3Ca<GNa<�  �  �Xa<�ba<ola<�sa<�ya<&}a<�~a<5a<�}a<M|a<za<�wa<{va<vua<ua<Yva<Bxa<�za<�}a<`�a<Ăa<o�a<}�a<9�a<�a<�za<Rsa<bja<x`a<�Ua<�Ka<Ba<n:a<�4a<�1a<�1a<�4a<�:a<�Ba<5Ma<�Xa<rda<>pa<�za<Q�a<��a<��a<��a<Ζa<�a<%�a<�a<��a<��a<ڐa<��a<D�a<��a<O�a<�a<��a<N�a<Ǡa<�a<ҡa<�a<ʛa<֕a<܍a<��a<za<Zoa<�da<Y[a<Ta<�Na<eLa<�La<Pa<tVa<�^a<�ha<�sa<�~a<��a<P�a<e�a<��a<ӥa<ԧa<�a<��a<��a<��a<�a<"�a<��a<�a<`�a<��a<��a<ݢa<��a<��a<8�a<]�a<�a<��a<��a<��a<��a<w�a<Lza<moa<�da<�[a<�Ta<�Oa<tNa<kOa<�Sa<mZa<,ca<�ma<Pxa<\�a<t�a<��a<��a<�a<O�a<��a<��a<��a<�a<*�a<��a<��a<'�a<��a<��a<R�a<�a<v�a<��a<a�a<e�a<Ǥa<Ԣa<Ğa<��a<ʐa<�a<q|a<"qa<+fa<�[a</Sa<�La<�Ha<Ha<�Ia<�Na<�Ua<9_a<�ia<4ta<�~a<3�a<f�a<��a< �a<�a<��a<b�a<��a<R�a<�a<"�a<Ҏa<�a<D�a<��a<]�a<��a<��a<�a<"�a<�a<|�a<h�a<�a<��a<�xa<na<�ba<�Va<SKa<�@a<�8a<<2a<K/a<�.a<l1a<7a<~>a<Ha<`Ra<�\a<ga<$pa<�wa<@}a<��a<y�a<��a<7�a<�~a<L|a<Mya<�va<ua<$ta<ta<ua<�va<�xa< {a<�|a<*~a<~a<�|a<Pya<�sa<�la<qca<MYa<Na<$Ca<x8a<Z/a<W(a<�#a<U"a<j#a<�'a<�.a<�7a<UBa<IMa<�  �  mYa<�ca<�la<ta<�ya<�|a<�~a<y~a<H}a<P{a<ya<�va<+ua<Qta<Tta<3ua<�va<�ya<�|a<{a<�a<��a<3�a<�a<�a<�za<�sa<ka<Taa<�Va<�La<=Ca<�;a<6a<3a<3a<6a<�;a<#Da<DNa<�Ya<Wea<�pa<i{a<��a<�a<<�a<��a<G�a<a�a<n�a<דa<�a<��a<��a<n�a<)�a<��a<&�a<1�a<l�a<��a<�a<��a<��a<��a<�a<$�a<\�a<;�a<�za<2pa<�ea<�\a<#Ua<�Oa<~Ma<�Ma<rQa<�Wa<�_a<�ia<�ta<�a<R�a<��a<��a<��a<u�a<��a<ۧa<ަa<�a<�a<�a<�a<x�a<�a<A�a<j�a<o�a<�a<��a<ߦa<x�a<�a<˧a<Фa<͟a<�a<$�a<?�a<G{a<Kpa<�ea<�\a<�Ua<;Qa<�Oa<�Pa<�Ta<�[a<Kda<xna<Nya<1�a<�a<�a<��a<�a<�a<M�a<ߦa<G�a<�a<3�a<��a<\�a<�a<�a<әa<�a<�a<j�a<��a<��a<��a<|�a<��a<��a<�a<.�a<ɇa<L}a<ra<ga<�\a<PTa<�Ma< Ja<"Ia<+Ka<	Pa<9Wa<H`a<xja<ua<�a<��a<��a<��a<��a<��a<��a<��a<G�a<<�a<�a<��a<~�a<�a<)�a<6�a<4�a<ʍa<��a<M�a<o�a<��a<*�a<�a<�a<
�a<ya<�na<bca<�Wa<YLa<Ba<�9a<�3a<d0a<0a<�2a<,8a<�?a<
Ia<JSa<�]a<�ga<�pa<�wa<=}a<��a</�a<��a<��a<~a<3{a<Ixa<�ua<�sa<�ra<�ra<�sa<uua<�wa<�ya<|a<k}a<�}a<R|a<*ya<�sa<�la<da<Za<
Oa<Da<�9a<�0a<�)a<%a<i#a<�$a< )a<�/a<�8a<3Ca<GNa<�  �  C[a<ea<�ma<�ta<{ya<L|a<b}a<�|a<;{a<�xa< va<qsa<cqa<npa<@pa<gqa<Esa<>va<�ya<�|a<�a<�a<<�a<a�a<�a<?{a<�ta<�la<Nca<}Ya<�Oa<�Fa<;?a<:a<87a<'7a<J:a<�?a<�Ga<�Qa<R\a<�ga<�ra<�|a<Y�a<J�a<��a<�a<�a<��a<:�a<�a<��a<��a<��a<s�a<$�a<ݍa<��a<�a<s�a<H�a<*�a<#�a< a<N�a<>�a<Ζa<��a<ކa<!}a<�ra<ia<F`a<�Xa<&Ta<�Qa<+Ra<�Ua<6[a<lca<�la<Ewa<ցa<�a<הa<2�a<��a<��a<��a<H�a<�a<u�a<{�a<Üa<3�a<��a<�a<X�a<��a<��a<۞a<��a<Ťa<��a<��a<�a<��a<A�a<��a<��a< �a<�}a<sa<Fia<�`a<�Ya<zUa<�Sa<Ua<�Xa<Q_a<�ga<Tqa<�{a<�a<��a<̗a<]�a<��a<u�a<,�a<�a<9�a<)�a<"�a<�a<��a<�a<j�a<�a<S�a<��a<^�a</�a<��a<�a<��a<��a<ٞa<p�a<6�a<T�a<Ga<�ta<	ja<q`a<�Wa<�Qa<7Na<9Ma<gOa<�Sa<�Za<�ca<:ma<jwa<1�a<�a<n�a<�a<n�a<�a<��a<ʙa<�a<K�a<�a<o�a<��a<�a<#�a<b�a<��a<��a<��a<�a<��a<"�a<l�a<��a<Z�a<��a<Lza<tpa<�ea<\Za<�Oa<�Ea<q=a<�7a<�4a<F4a<�6a<�;a<[Ca<La<�Ua<�_a<Nia<�qa<txa<q}a<#�a<S�a<k�a<�~a<�{a<0xa<ua<	ra<pa<�na<oa<�oa<�qa<�ta<,wa<�ya<�{a<v|a<�{a<ya<qta<�ma<�ea<�[a<yQa<�Fa<�<a<C4a<j-a<C)a<{'a<)a<-a<�3a<@<a<Fa<�Pa<�  �  �^a<�ga<Hoa<ua<7ya<!{a<e{a<za<�wa<Zta<qa<na<�ka<lja<.ja<|ka<�ma<�pa<�ta<�xa<�|a<�a<b�a<|�a<�a<|a<�va<Eoa<�fa<�]a<yTa<'La<!Ea<@a<�=a<�=a<c@a<�Ea<XMa<Va<�`a<dka<�ua<�~a<��a<��a<��a<k�a<��a<v�a<I�a<��a<ǉa<g�a<��a<W�a<	�a<�a<�a<ˎa<�a<F�a<��a<ӝa<%�a<͞a<c�a<�a<őa<��a<ǀa<Xwa<na<�ea<�^a<6Za<Xa<�Xa<�[a<2aa<�ha<�qa<�{a<X�a<��a<ɖa<�a<��a<5�a<�a<ӣa<}�a<T�a<ٚa<v�a<��a<ϒa<Αa<K�a<�a<v�a<ҙa<t�a<��a<ڣa<��a<إa<e�a<��a<H�a<�a<+�a<��a<�wa<jna<=fa<�_a<�[a<Za<D[a<�^a<ea<�la<va<�a<G�a<�a<v�a<��a<��a<J�a<.�a<h�a<��a<�a<1�a<��a<�a<�a<W�a<�a<��a<]�a<��a<�a<,�a<��a<��a<�a<��a<=�a<�a<��a<��a<�xa<�na<�ea<�]a<�Wa<�Ta<�Sa<�Ua<�Ya<o`a<�ha<�qa<'{a<.�a<U�a<��a<U�a<�a<��a<n�a<��a<#�a<��a<��a<چa<��a<Ӂa<	�a<��a<�a<d�a<:�a<�a<X�a<юa<ώa<,�a<�a<Ճa<||a<Vsa<Fia<�^a<vTa<@Ka<�Ca<�=a<�:a<�:a<�<a<�Aa<�Ha<�Pa<)Za<[ca<la<�sa<Yya<k}a<ba<�a<�}a<#{a<�wa<�sa<�oa<sla<@ja<�ha<�ha<Hja<}la<�oa<�ra<,va<�xa<hza<_za<�xa<�ta<Toa<�ga<�^a<bUa<yKa<Ba<�9a<w3a<u/a<�-a<A/a<3a<^9a<pAa<�Ja<�Ta<�  �  �ba<uja<%qa<�ua<�xa<�ya<�xa<xva<�ra<�na<�ja<�fa<�ca<`ba<Eba<aca<	fa<�ia<lna<^sa<xa<A|a<
a<h�a<�a<"}a<�xa<mra<ka<�ba<�Za<�Ra<�La<9Ha<�Ea<Fa<�Ha<�Ma<�Ta<]a<|fa<*pa<bya<w�a<.�a<�a<ۏa<��a<ԏa<��a<,�a<��a<��a<�a<~a<_}a<~a<�a<��a<�a<�a<�a<�a<Қa<!�a<�a<��a<j�a<'�a<f�a<y�a<�|a<�ta<�la<�fa<dba<�`a<�`a<�ca<ia<�oa<xa<ڀa<։a<�a<��a<O�a<��a<=�a<��a<��a<$�a<��a<��a<f�a<�a<��a<܉a<@�a<�a<2�a<5�a<Зa<�a</�a<�a<S�a<�a<b�a<�a<��a<5�a<��a<�}a<ua<�ma<�ga<�ca<�ba<�ca<ga<�la<�sa<|a<Ԅa<p�a<�a<S�a<��a<b�a<�a<��a<ܞa<ǚa<]�a<��a<u�a<)�a<�a<k�a<��a<�a<=�a<F�a<��a<��a<2�a<P�a<��a<��a<Q�a<�a<%�a<�a<~a<ua<�la<�ea<`a<�\a</\a<�]a<�aa<�ga<oa<fwa<�a<��a<юa<D�a<��a<P�a<��a<��a<͒a<�a<�a<�a<ya<|a<�ya<ya<�ya<�{a<�~a<9�a<Ѕa<G�a<Ћa<ʌa<c�a<��a<N�a<�~a<�va<�ma<Zda<�Za<fRa<|Ka<Fa<gCa<Ca<Ea<�Ia<�Oa<JWa<{_a<�ga<Yoa<�ua<�za<m}a<k~a<I}a<�za<�va<)ra<Rma<�ha<�da<$ba<�`a<�`a<vba<:ea<�ha<Dma<Lqa<"ua<�wa<�xa<Exa<�ua<qa<�ja<ca<TZa<aQa<�Ha<hAa<�;a<�7a<w6a<�7a<6;a<�@a<(Ha<�Pa<�Ya<�  �  Pga<�ma<Gsa<�va<]xa<�wa<�ua<�qa<Dma<ha<�ba<^a<
[a<Ya<�Xa<Za<@]a<�aa<�fa<�la<�ra<xa<|a<�~a<�a<Y~a<{a<%va<pa<�ha<�aa<*[a<�Ua<�Qa<zOa<�Oa<Ra<�Va<�\a<�da<ma<�ua<�}a<c�a<��a<f�a<��a<e�a<�a<��a<O�a<�a<{a<�wa<�ta<ta<�ta<�va<�za<�a<ƅa<�a<��a<��a<Кa<�a<��a<	�a<�a<��a<Ɋa<H�a< |a<=ua<�oa<�ka<ja<�ja<!ma<�qa<�wa<\a<�a<�a<͕a<}�a<��a<��a<ˡa<�a<{�a<��a<��a</�a<P�a<M�a<r�a<i�a<�a<�a<Ԇa<}�a<�a<x�a<��a<��a<c�a<E�a<3�a<�a<��a<��a<>�a<��a<�|a<2va<�pa<vma<,la<ma<9pa<'ua<�{a<�a<��a<�a<[�a<v�a<��a<�a<�a<`�a<W�a<@�a<��a<�a<%�a<4�a<�~a<�}a<�~a<H�a<�a<ʉa<)�a<e�a<�a<`�a<f�a<o�a<��a<��a<ܒa<�a<�a<Q|a<�ta<Cna<nia<zfa<�ea<8ga<�ja<pa<�va<�}a<a�a<<�a<��a<�a<1�a<V�a<~�a<Ԓa<�a<*�a<�a<|a<�va<�ra<pa<�oa<tpa< sa<�va<�za<�a<S�a<��a<y�a<B�a<�a<�a<��a<{a<Fsa<�ja<�ba<�Za<CTa<�Oa<�La<�La<zNa<LRa<�Wa<�^a<�ea<�la<8sa<Sxa<�{a<j}a<�|a<�za<�va<�qa<�ka<�ea<�`a<)\a<�Xa<{Wa<�Wa<uYa<�\a<9aa<_fa<�ka<pa<Rta<�va<�wa<`va< sa<�ma<�ga<�_a<2Xa<�Pa<�Ia<�Da<9Aa<@a<Aa<VDa<pIa<)Pa<�Wa<�_a<�  �  #la<}qa<lua<zwa<�wa<�ua<:ra<4ma<(ga<�`a<�Za<TUa<NQa<�Na<tNa<Pa<�Sa<�Xa<�^a<�ea<�la<�sa<ya<	}a<"a<Fa<�}a< za<$ua<Xoa<Wia<�ca<�^a<m[a<�Ya<�Ya<:\a<G`a<�ea<�la<�sa<M{a<�a<��a<��a<��a<��a<ߋa<E�a<p�a<�}a<�wa<�ra<na<ka<�ia<bja<ma<nqa<Twa< ~a<e�a<��a<��a<(�a<��a<��a<u�a<��a<ŕa<O�a<%�a<ރa<~a<Bya<�ua<Qta<�ta<wa<{a<��a<�a<��a<!�a<Ǚa<+�a<��a<i�a<#�a<��a<,�a<@�a<��a<F�a<ka<�za<�wa<va<�va<Qya<�}a<-�a<��a<7�a<��a<�a<(�a<\�a<��a<
�a<|�a<o�a<G�a<��a</�a<Wa<�za<�wa<mva<Swa<za<]~a<�a<D�a<ːa<�a<��a<��a<V�a< �a<�a<�a<��a<"�a<T�a<ׁa<�{a<vwa<�ta<�sa<�ta<�wa<|a<ʁa<�a<��a<|�a<O�a<��a<�a<q�a<�a<��a<�a<��a<��a<I}a<�wa<Ssa<�pa<�oa<Zqa<ita<ya<�~a<�a<�a<��a<��a<��a<]�a<�a<��a<��a<��a<��a<_za<�sa<�ma<ia<7fa<aea<�fa<{ia<�ma<Hsa<#ya<�~a<��a<Їa<�a<�a<W�a<��a<Xa<�xa<�qa<Oja<�ca<�]a<�Ya<4Wa<�Va<mXa<�[a<�`a<+fa<8la<&ra<3wa<{a<�|a<$}a<T{a<�wa<Vra<�ka<�da<^a<�Wa<�Ra<�Na<!Ma<vMa<�Oa<�Sa<�Xa<�^a<iea<�ka<�pa<�ta<�va<�va<ua<dqa<>la<fa<S_a<�Xa< Sa<]Na<jKa<DJa<HKa<Na<�Ra<~Xa<�^a<�ea<�  �  �pa<�ta<nwa<&xa<�va<�sa<�na<Pha<�`a<�Ya<YRa<La<~Ga<�Da<6Da<�Ea<�Ia<�Oa<�Va<�^a<ga<�na<�ua<,{a<�~a<C�a<�a<�}a<za<�ua<�pa<la<,ha<;ea<�ca<=da<#fa<�ia<�na<|ta<�za<�a<C�a<x�a<�a<Ǎa<��a<�a<;�a<!~a<wa<apa<�ia<�da<aa<�_a<)`a<ca<�ga<�na<qva<�~a<�a<Ԏa</�a<4�a<�a<�a<��a<ߙa<Еa<�a<��a<ʆa<ςa<�a<�~a<�~a<�a<��a<�a<i�a<�a<D�a<��a<��a<ۡa<'�a<r�a<��a<��a<v�a<��a<T}a<nva<�pa<Uma<�ka<�la<qoa<<ta<�za<'�a<̉a<��a<E�a<��a<��a</�a<�a<��a<��a<3�a<��a<8�a<^�a<d�a<��a<ˀa<h�a<��a<�a<&�a<{�a<ؖa<��a<F�a<��a<�a<g�a<Ŝa<R�a<��a<߈a<�a<rya<�ra<�ma<`ja<Tia<�ja<�ma<sa<�ya<�a<��a<܏a<�a<��a<��a<m�a<P�a<N�a<�a<ܐa<,�a<��a<�a<!}a<�za<Sza<E{a<~a<ځa<��a<͋a<��a<ڔa<՗a<8�a<��a<��a<2�a<�a<m�a<�za<�ra<�ja<da<_a< \a<([a<�\a<�_a<ea<�ka<Tra<xya<�a<քa<��a<$�a<ɉa<p�a<q�a<K~a<Xxa<ra<Fla<bga<�ca<�aa<aa<Eba<%ea< ia<�ma<�ra<Iwa<�za<w}a<$~a<�|a<�ya<Xta<�ma<%fa<�]a<Va<�Na<�Ha<�Da<�Ba<;Ca<�Ea<IJa<nPa<�Wa<�^a<�fa<�la<Ara<�ua<Zwa<�va<�ta<�pa<�ka<mfa<�`a<\a<Xa<pUa<�Ta<ZUa<�Wa<�[a<�`a<-fa<�ka<�  �  Bua<�wa<2ya<�xa<�ua<kqa<ka<�ca<[a<�Ra<KJa<�Ca<Q>a<);a<�:a<j<a<�@a<'Ga<Oa<Xa<laa<|ja<yra<5ya<�}a<�a<߁a<�a<�~a<]{a<�wa<�sa<�pa<Dna<;ma<�ma<^oa<�ra<�va<�{a<�a<�a<M�a<�a<{�a<��a<�a<�a<J�a<ya<�pa<�ha<�aa<�[a<�Wa<�Ua<�Va<�Ya<&_a<5fa<�na<Mxa<�a<��a<x�a<��a<Ϝa<�a<'�a<ŝa<Қa<��a<�a<ʎa<j�a<
�a<�a<S�a<�a<��a<�a<��a<ޙa<�a<.�a<��a<¢a<��a<��a<��a<^�a<�a<~a<�ua<na<ha<�ca<@ba<�ba<)fa<�ka<�ra<�za<ڃa<��a<��a<e�a<]�a<r�a<��a<��a<I�a<��a<H�a<��a<��a<=�a<��a<E�a<��a<��a<a<��a<*�a<O�a<�a<w�a<b�a<k�a<h�a<��a<Փa<��a<�a<za<bqa<-ja<uda<�`a<�_a<�`a<�da<�ja<�qa<@za<��a<d�a<��a<Ęa<ۜa<*�a<O�a<͝a<ƚa<��a<!�a<j�a<Q�a<+�a<=�a<��a<��a<��a<�a<�a<��a<֕a<�a<u�a<��a<��a<��a<��a<�a<N~a<�ta<cka<�ba<d[a<�Ua<lRa<�Qa<Sa<2Wa<�\a<da<
la<;ta<�{a<�a<�a<�a<��a<ىa<U�a<L�a<d~a<[ya<Eta<�oa<�la<�ja<jja<\ka<�ma<�pa<�ta<�xa<|a<�~a<�a<a<N|a<�wa<Wqa<�ia<�`a<VWa<TNa<VFa<�?a<K;a<X9a<�9a<�<a<�Aa<NHa<vPa<Ya<�aa<\ia<�oa<�ta<�wa<�xa<�wa<ua<Cqa<�la<dha<1da<�`a<�^a<^a<�^a<�`a<da<7ha<�la<>qa<�  �  �xa<rza<|za<�xa<ua<�oa< ha<a_a<�Ua<qLa<�Ca<�;a<%6a<�2a<.2a</4a<�8a<�?a<]Ha<4Ra<�\a<�fa<�oa<�wa<o}a<��a<y�a<ԃa<��a<N�a<j}a<vza<�wa<va<Aua<�ua<xwa<za<�}a<�a<^�a<S�a<v�a<K�a<c�a<��a<ȉa<D�a<�|a<tta<�ka<�ba<�Za<Ta<�Oa<�Ma<)Na<eQa<8Wa<_a<qha<�ra<=}a<0�a<%�a<?�a<��a<�a<=�a<Ԡa<��a<6�a<��a<��a<�a<�a<�a<R�a<�a<P�a<��a<P�a<�a<�a<�a<}�a<h�a<&�a<��a<�a<��a<"�a<cxa<�na<�fa<`a<�[a<�Ya<�Za<�]a<�ca<�ka<�ta<�~a<j�a<��a<f�a<\�a<��a<��a<
�a<��a<�a<��a<%�a<��a<�a<�a<0�a<˒a<i�a<��a<;�a<��a<��a<��a<�a<��a<��a<��a<��a<�a<��a<�}a<�sa<�ja<�ba<F\a<�Xa<GWa<�Xa<�\a<ca<+ka<cta<~a<i�a<�a<�a<K�a<��a<�a<��a<��a<}�a<їa<�a<��a<�a<D�a<��a<��a<?�a<�a<�a<N�a<�a<�a<��a<~�a<p�a<A�a<`�a<��a<�ya<boa<ea<�[a<�Sa<|Ma<Ja<(Ia<�Ja<DOa<�Ua<�]a<�fa<�oa<+xa<�a<��a<��a<Ћa<�a<d�a<o�a<��a<ma<2{a<vwa<�ta<�ra<ira<Gsa<�ta<�wa<�za<�}a<�a<r�a<W�a<�a<�{a<2va<�na<�ea<�[a<�Qa<�Ga< ?a<�7a<3a<�0a<X1a<a4a<�9a<Aa<LJa<�Sa<^]a<Hfa<�ma<�sa<�wa<�ya<�ya<uxa<�ua<`ra<�na<Uka<�ha<�fa< fa<�fa<|ha<6ka<�na<]ra<�ua<�  �  c{a<g|a<�{a<ya<ata<�ma<�ea<\a<�Qa<�Ga<U>a<*6a<0a<�,a<�+a<.a<�2a<:a<FCa<�Ma<�Xa<fca<nma<va<�|a<�a<΄a<�a<i�a< �a<��a<�a<_}a<�{a<P{a<�{a<J}a<�a<�a<��a<v�a<��a<�a<�a<�a<��a<؈a<C�a<"za<�pa<4ga<�]a<EUa<Na<}Ia<(Ga<�Ga<YKa<'Qa<�Ya<�ca<fna<�ya<Y�a<�a<.�a<��a<��a<�a<0�a<3�a<@�a<n�a<��a<|�a<ٖa<�a<l�a<��a<�a<ʜa<��a<Ӣa<�a<1�a<�a<ͣa<ԟa<��a<ˑa<{�a<Y~a<�sa<�ia< aa<�Ya<wUa<CSa<ITa<�Wa<^a<wfa<pa<�za<	�a<�a<��a<��a<ţa<��a<�a<:�a<��a<�a<�a<�a<��a<�a<B�a<Șa<�a<_�a< �a<�a<��a<0�a<�a<ɥa<�a<�a<��a<Z�a<v�a<�ya<2oa<iea<�\a<<Va<?Ra<�Pa<�Ra<�Va<}]a<fa<�oa<3za<J�a<��a<��a<ڛa<	�a<<�a<��a<\�a<O�a<�a<&�a<"�a<��a<T�a<Ƒa<m�a<֓a<6�a<��a<f�a<u�a<|�a<k�a</�a<n�a<Q�a<`�a<ڀa<8va<ka<`a<6Va<�Ma<vGa<�Ca<�Ba<�Da<4Ia<EPa<�Xa<"ba<�ka<Sua<�}a<��a<��a<_�a<��a<��a<��a<��a<ۃa<o�a<}a<�za<�xa<�xa<�xa<�za<�|a<�~a<v�a<�a<��a<˂a<�a<�{a<�ta<~la<�ba<Xa<Ma<�Ba<s9a<�1a<�,a<^*a<+a<[.a<4a<9<a<zEa<�Oa<�Ya<�ca<la<�ra<�wa<�za<�{a<{a<\ya<�va<�sa<�pa<-na<�la<la<�la<na<�pa<�sa<�va<�ya<�  �  #}a<�}a<3|a<ya<�sa<�la<da<7Za<tOa<�Da<�:a<~2a<4,a<c(a<�'a<�)a<�.a<j6a<�?a<�Ja<>Va<�aa<la<@ua<�|a<�a<~�a<'�a<?�a<?�a<��a<��a<݀a<�a<=a<�a<�a<^�a<S�a<��a<ڌa<��a<i�a<ܑa<��a<b�a<<�a<!�a<�xa<�na<�da<�Za<�Qa<dJa<XEa<�Ba<�Ca<&Ga<xMa<Va<``a<�ka<owa<��a<Ռa<��a<:�a<�a<��a<��a<"�a<��a<j�a<(�a<�a<��a<#�a<c�a<v�a<l�a<�a<��a< �a<Ǧa<~�a<��a<�a<k�a<�a<t�a<ʆa<�{a<qa<�fa<q]a<&Va<;Qa</Oa<Pa<�Sa<bZa<�ba<ma<xa<�a<e�a<��a<�a<��a<>�a<�a<�a<��a<��a<��a<n�a<C�a<ݜa<X�a<��a<ѝa<ȟa<1�a<��a<��a<�a<�a<e�a<�a<c�a<�a<یa<��a<iwa<Ola<�aa<Ya<SRa<Na<�La<RNa<�Ra<�Ya<�ba<�la<�wa<��a<=�a<˔a<j�a<+�a<�a<٣a<2�a<n�a<��a<;�a<��a<��a<@�a<וa<9�a<��a<q�a<��a<ʝa<k�a<�a<<�a<��a<2�a<��a<>�a<Ba<ta<sha<]a<�Ra<�Ia<QCa<u?a<�>a<�@a<�Ea<�La<�Ua<u_a<�ia<�sa<z|a<�a<Q�a<Ìa<]�a</�a<��a<��a<׆a<��a<��a<_~a<}a<y|a<�|a<~a<�a<ҁa<��a<̈́a<�a<��a<N�a<+{a<%ta<'ka<�`a<�Ua<NJa<l?a<�5a<.a<�(a<K&a<�&a<_*a<s0a<�8a<�Ba<5Ma<Xa< ba<ka<fra<�wa<A{a<�|a<�|a<\{a<(ya<�va<ta<�qa<�pa<%pa<�pa<�qa<ta<�va<Eya<�{a<�  �  :ya<Uya<>xa<�ua<�qa<Mla<�ea<.^a<�Ua<Na<�Fa<k@a<�;a<9a<9a<):a<;>a<�Ca<)Ka<qSa<*\a<�da<�la<2ta<�ya<�~a<R�a<܂a<A�a<��a<��a<d�a<1a<m~a<&~a<�~a<�a<�a<9�a<�a<X�a<��a<�a<R�a<��a<�a<�a<��a<Eza<*sa<wka<Gda<�]a<�Xa<�Ta<oSa< Ta<rVa<�[a<�aa<ja<�ra<�{a<U�a<=�a<�a<Z�a<m�a<��a<��a<x�a<R�a<*�a<S�a<�a<јa<s�a<��a<��a<+�a<�a<D�a<Ơa<:�a<��a<ۡa<�a<
�a<�a<��a<1�a<�a<�xa<qa<ja<�da<�`a<�_a<I`a<�ba<�ga<Mna<	va<)~a<��a<r�a<��a<R�a<ɟa<��a<�a<L�a<\�a<֡a<�a<�a<�a<@�a<�a<�a<�a<��a<Y�a<�a<t�a<_�a<0�a<̡a<��a<��a<Ԕa<��a<�a<N}a<ua<ma<nfa<Faa<^a<�]a< ^a<�aa<�fa<dma<ua<'}a<Q�a<��a<4�a<8�a<&�a<8�a<�a<��a<>�a<��a<o�a<f�a<ŕa<��a<G�a<|�a<~�a<͖a<��a<řa<�a<'�a<@�a<3�a<Q�a<)�a<��a<��a<=xa<&oa<�fa<a^a<�Wa<�Ra<�Oa<;Oa<Pa<�Sa<�Xa<�_a<�fa<tna<�ua<Z|a<�a<��a<݈a<��a<͉a<��a<e�a<A�a<w�a<$a<1}a<�{a<m{a<�{a<r|a<�}a<.a<�a<�a<��a<Sa<�|a<exa<�ra<�ka<�ca<][a<�Ra<eJa<�Ba<O=a<�8a<�7a<�7a<�9a<�>a<�Da<)La<Ta<W\a<�ca<�ja<Rpa<�ta<fwa<�xa<�xa<�wa<0va<hta<era<�pa<�oa<loa<�oa<�pa<pra<{ta<dva<xa<�  �  �xa<�xa<�wa<�ua<�qa<�la<�ea<�^a<�Va<�Na<�Ga<bAa<�<a<�9a<}9a<-;a<;?a<�Da<La<1Ta<�\a<iea<[ma<rta<za<K~a<��a<��a<ǂa<#�a<݀a<�a<[~a<�}a<T}a<�}a<a<�a<p�a<�a<��a<�a<��a<�a<.�a<��a<<�a<�a<�za<�sa<,la<ea<�^a<cYa<�Ua<Ta<�Ta<�Wa<�\a<�ba<�ja<^sa<H|a<ʄa<��a<E�a<z�a<�a<L�a<*�a<��a<��a<4�a<��a< �a<�a<��a<ӗa<Ęa<^�a<N�a<S�a<K�a<��a<:�a<��a<��a<0�a<O�a<��a<��a<��a<�ya<�qa<ka<�ea<�aa<l`a<aa<da<�ha<Boa<�va<�~a<+�a<�a<ܕa<��a<��a<a�a<ƣa<ɣa<�a<�a<-�a<<�a<��a<v�a<�a<=�a<4�a<��a<{�a<=�a<��a<ޢa<ڢa<y�a<�a<��a<!�a<!�a<a�a<�}a<�ua<na<fga<\ba<�^a<�]a<$_a<�ba<�ga<Ona<�ua<�}a<��a<
�a<u�a<c�a<�a<�a<��a<1�a<ǜa<��a<��a<��a<��a<ɓa<g�a<��a<��a<�a<��a<!�a<g�a<��a<��a<��a<i�a<]�a<�a<*�a<�xa<�oa<bga<e_a<�Xa<�Sa<�Pa<�Oa<EQa<�Ta<�Ya<Y`a<sga<oa<2va<�|a<�a<�a<��a<��a<V�a<�a<υa<K�a<��a<]~a<`|a< {a<�za<�za<�{a<�|a<>~a<�a<d�a<G�a<�~a<|a<�xa<!sa<Dla<wda< \a<dSa<IKa<�Ca<D>a<:a<*8a<u8a<";a<�?a<�Ea<�La<�Ta<�\a<Eda<ka<�pa<�ta<wa<Xxa<Bxa<Hwa<pua<�sa<�qa<�oa<�na<�na<�na<�oa<�qa<�sa<�ua<�wa<�  �  Qwa<2xa<~wa<�ua<ra<?ma<(ga<`a<�Xa<�Pa<Ja<Da<�?a<7=a<�<a<u>a<�Aa<Ga<zNa<HVa<�^a<�fa<sna<�ta<Qza<~a<��a<��a<C�a<{�a<�~a<F}a<�{a<�za<lza<�za<=|a<G~a<�a<܃a<�a<��a<Q�a<m�a<Ћa<�a<��a<�a<�{a<Uua<=na<Gga<+aa<�[a<�Xa<LWa<�Wa<�Za<(_a<�ea<ma<uua<�}a<�a<��a<��a<��a<śa<ȝa<��a<_�a<�a<��a<*�a<Y�a<#�a<��a<�a<�a<��a<�a<!�a<��a<.�a<3�a<�a<_�a<f�a<��a<�a<�a<��a<�{a<>ta<�ma<gha<6ea<�ca<Tda<ga<}ka<�qa<�xa<ڀa<��a<�a<��a<Лa<��a<��a<�a<m�a<H�a<)�a<�a<��a<јa<��a<�a<c�a<i�a<�a<4�a<B�a<^�a<u�a<�a<�a<Ϟa<��a<ƕa<O�a<ۇa<�a<�wa<�pa<ja<;ea<?ba<&aa<mba<bea<Sja<�pa<�wa<�a<$�a<#�a<�a<��a<��a<u�a<��a<��a<�a<��a<Q�a<�a<�a<��a<\�a<Ґa<��a<��a<a�a<T�a<Ϙa<r�a<Z�a<��a<��a<��a<��a<q�a<hza<�qa<�ia<ba<c[a<�Va<�Sa<Sa<vTa<iWa<}\a<�ba<�ia<�pa<�wa<�}a<{�a<?�a<5�a<�a<*�a<y�a<�a<�a<O~a<�{a<�ya<xa<�wa<�wa<�xa<�za<|a<�}a<�~a<?a<�~a<F|a<�xa<�sa<Nma<�ea<�]a<vUa<�Ma<�Fa<�@a<U=a<X;a<�;a<>a<2Ba<7Ha<Oa<�Va<P^a<~ea<�ka<�pa<�ta<�va<�wa<�va<�ua<�sa<Cqa<oa</ma<la<uka<la<.ma<oa<Vqa<�sa<�ua<�  �  Jua<�va<�va<zua<�ra<mna<�ha<�ba<�[a<~Ta<Na<wHa<$Da<�Aa<eAa<�Ba<vFa<�Ka<RRa<�Ya<�aa<ia<pa<�ua<�za<�}a<�a<�a<a<�}a<�{a<kya<�wa<mva<�ua<eva<�wa<�ya<�|a<]�a<ԃa<�a<}�a<�a<L�a<)�a<W�a<d�a<~a<�wa<vqa<�ja<Gea<�`a<?]a<�[a<�\a<,_a<�ca<�ia<�pa<�xa<��a<-�a<�a<|�a<��a<W�a<��a<6�a<�a<�a<��a<�a<�a<ϐa<%�a<r�a<��a<o�a<�a<�a<��a<�a<��a<�a<�a<��a<��a<��a<5�a<C�a<a<xa<�qa<�la<�ia<Wha<�ha<{ka<�oa<�ua<}|a<�a<+�a<��a<ݗa<h�a<��a<E�a<��a<|�a<��a<	�a<I�a<��a<��a<�a<��a<�a<�a<��a<|�a< �a<��a<m�a<��a<D�a<��a<��a<��a<�a<E�a<�a<l{a<�ta<|na<�ia<�fa<�ea<�fa<�ia<�na<�ta<U{a<��a<i�a<̏a<��a<�a<��a<|�a<�a<��a<<�a<c�a<v�a<��a<ōa<g�a<�a<k�a<��a<��a<�a<@�a<L�a<��a< �a<��a<��a<w�a<0�a<v�a<}a<%ua<'ma< fa<�_a<;[a<�Xa<�Wa<�Xa<�[a<�`a<<fa<�la<[sa<�ya</a<V�a<\�a<Ǉa<ʇa<c�a<�a<�a<�}a<?za<Pwa</ua<�sa<4sa<�sa<�ta<�va<�xa<�za<�|a<�}a<{}a<�{a<	ya<�ta<�na<ha<�`a<�Xa<kQa<�Ja<sEa<�Aa<@a<R@a<�Ba<�Fa<6La<�Ra<�Ya<�`a<Zga<ma<hqa<�ta<�ua<"va<�ta<�ra<epa<�ma<�ja<�ha<�ga<	ga<�ga<�ha<�ja<�ma<{pa<-sa<�  �  �ra<�ta<�ua<)ua<Csa<�oa<-ka<�ea<X_a<Ya<�Ra<Na<8Ja<�Ga<�Ga<Ia<vLa<1Qa<9Wa<$^a<ea<�ka<(ra<Uwa<{a<a}a<>~a<�}a<6|a<�ya<<wa<nta<+ra<�pa<�oa<Fpa<�qa<�ta<�wa<�{a<�a<��a<�a<V�a<{�a<�a<O�a<�a<��a<+{a<ua<�oa<bja<Ofa<_ca<?ba<�ba<Oea<�ia<�na<�ua<�|a<�a<Ɗa<ǐa<��a<ɘa<��a<ךa<�a<Ǘa<��a<�a<�a<��a<Ȋa<��a<>�a<��a<�a<��a<��a<ȗa<��a<]�a<��a<��a<��a<��a<��a<�a<Ɖa<a�a<�|a<Awa<�ra<�oa<�na<+oa<�qa<�ua<�za<7�a<Ňa<M�a<F�a<g�a<)�a<o�a<?�a<��a<ݝa<
�a<�a<��a<W�a<ڎa<�a<k�a<��a<Z�a<��a<��a<�a<��a<��a<��a<#�a<c�a<&�a<r�a<U�a<U�a<��a<�a<vya<
ta<�oa<ma<+la<ma<�oa<	ta<xya<�a<�a<X�a<ڑa<Y�a<m�a<�a<%�a<��a<��a<h�a<�a<x�a<`�a<�a<<�a<΅a<b�a<�a<Z�a<P�a<7�a<��a<5�a<C�a<+�a<��a<o�a<،a<�a<>�a<-ya<�qa<;ka<�ea<Zaa<�^a<�]a<�^a<�aa<�ea<ka<�pa<�va</|a<�a<f�a<j�a<�a<!�a<�a<�a<
}a<#ya<'ua<�qa<)oa<�ma<ma<�ma<Xoa<�qa<jta<wa<�ya<i{a<|a<h{a<Vya<�ua<�pa<�ja<da<5]a<PVa<0Pa<kKa<�Ga<SFa<�Fa<�Ha<ULa<5Qa<UWa<�]a<�ca<�ia<�na<*ra<Gta<�ta<4ta<Zra<toa<Fla<�ha<�ea<:ca<taa<�`a<caa<"ca<�ea<�ha<Lla<�oa<�  �  Foa<`ra<<ta<�ta<�sa<�qa<�ma<ia<�ca<H^a<�Xa<`Ta<�Pa<"Oa<�Na<APa<!Sa<�Wa<]a<"ca<Oia<Voa<�ta<�xa<�{a<�|a<�|a<<{a<�xa<�ua<ra<�na<�ka<�ia<�ha<Zia<�ja<�ma<�qa<Ava<${a<�a<�a<k�a<c�a<�a<L�a<�a<��a<a<za<.ua<�pa<�la<[ja<]ia<�ia<Zla<pa<&ua<6{a<��a<�a<�a<˒a<��a<טa<��a<�a<�a<�a<q�a<��a<��a<	�a<�a<�a<l�a<�a<��a<�a<1�a<}�a<Q�a<��a<�a<a<J�a<B�a<՗a<U�a<�a<@�a<��a<�}a<�ya<�va<�ua<Rva<ixa<|a<؀a<y�a<5�a<��a<�a<�a<�a<"�a<��a<{�a<��a<	�a<��a<؎a<�a<*�a<6�a<r�a<�a<��a<g�a<�a<�a<�a<h�a<9�a<ȝa<��a<ʜa<
�a<��a<�a<�a<8�a<sa<gza<�va</ta<Vsa<>ta<�va<`za<Pa<Ƅa<Q�a<��a<@�a<��a<ՙa<\�a<��a<g�a<�a<3�a<܋a<��a<�a<�a<la<�~a<�a<v�a<>�a<ća<��a<�a<*�a<V�a<�a<s�a<j�a<��a<��a<"�a<�}a<rwa<^qa<3la<Wha<�ea<ea<fa<Qha<�ka<�pa<�ua<�za<Ma<�a<|�a<y�a<�a<O�a<"�a<}a<�xa<�sa<oa<Hka<Oha<�fa</fa<�fa<�ha<�ka<oa<�ra<�ua<�xa<iza<�za<�ya<wa<sa<na<4ha<ba<\a<|Va<Ra<Oa<wMa<�Ma<oOa<�Ra<>Wa<�\a<ba<�ga<rla<Mpa<�ra<�sa<�sa<ra<!oa<tka<[ga<1ca<x_a<�\a<�Za<�Ya<�Za<o\a<[_a<	ca<Cga<�ka<�  �  �ka<�oa<�ra<Zta<�ta<#sa<�pa<�la<}ha<�ca<?_a<Y[a<TXa<�Va<eVa<�Wa<aZa<_^a< ca<gha<�ma<�ra<wa<za<�{a<|a<�za<oxa<�ta<�pa<\la<Zha<�da<oba<aaa<�aa<�ca<�fa</ka<Qpa<�ua<�{a<΀a<.�a<8�a<�a<3�a<�a<��a<�a<&a<�za<wa<�sa<�qa<�pa<�qa<�sa<7wa<�{a<��a<��a<�a<�a<�a<��a<�a<��a<�a<ӓa<�a<b�a<��a<��a<�~a<�|a<c{a<�{a<�}a<��a<ʄa<y�a<��a<z�a<��a<�a<��a<��a<��a<J�a<��a<Y�a<y�a<��a<]�a<��a<|~a<[}a<�}a<�a<�a<>�a<�a<�a<ʕa<�a<�a<��a<ܞa<��a<��a<)�a<��a<��a<Ɉa<u�a<�a<�~a<�}a<n~a<U�a<��a<ɇa<i�a<_�a<ѕa<��a<4�a<��a<d�a<��a<��a<��a<ۏa<��a<��a<c�a<�}a<�{a<�za<�{a<�}a<;�a<c�a<�a<��a<3�a<іa<�a<8�a<��a<ӗa<��a<W�a<~�a<7�a<e�a<!}a<�ya<�wa<)wa<+xa<Oza<�}a<Ӂa<d�a<�a<�a<�a<�a<l�a<R�a<ѐa<��a<.�a<Ԃa< }a<�wa<Rsa<�oa<�ma<�la<ma<yoa<�ra<qva<�za<�~a<o�a<!�a<��a<��a<�a<-�a<~a<�xa<xsa<�ma<�ha<1da<�`a<�^a<�^a<�_a<�aa<_ea<cia<�ma<ra<�ua<zxa<�ya<�ya<Yxa<�ua<{qa<�la<Jga<ba<H]a<?Ya<�Va<Ua<MUa<�Va<�Ya<�]a<ba<�fa<gka<Hoa<ra<�sa<�sa<;ra<�oa<�ka<ga<�aa<$]a<�Xa<IUa<1Sa<@Ra<Sa<!Ua<�Xa<�\a<�aa<�fa<�  �  	ha<ma<qa<�sa<�ta<�ta<4sa<tpa<ma<3ia<^ea<#ba<�_a<E^a<^a<A_a<�aa<�da<%ia<�ma<1ra<>va<�ya<{{a<|a<[{a<ya<�ua<qa<�ka<�fa<�aa<�]a<[a<�Ya<Za<\a<�_a<jda<ija<�pa<Fwa<�}a<Ȃa< �a<ȉa<
�a<�a<��a<�a<
�a<��a<d}a<�za<ya<�xa<Qya<&{a<E~a<2�a<҆a<��a<�a<�a<�a<��a<ɘa<z�a<��a<��a<��a<<�a<�a<�{a<�wa<ua<�sa<(ta<!va<�ya<A~a<׃a<��a<|�a<Ôa<�a<$�a<��a<̝a<��a<�a<��a<��a<��a<�a<�a<��a<�a<��a<#�a<�a<i�a<��a<Õa<}�a<��a<��a<,�a<k�a<�a<d�a<��a<	�a<O�a<��a<�}a<�ya<)wa<!va<�va<ya<�|a<��a<�a<��a<)�a<�a<��a<�a<֝a<L�a<^�a<:�a<m�a<%�a<ߋa<.�a<6�a<U�a<��a<B�a<�a<؇a<j�a<`�a<8�a<��a<=�a<��a<m�a<��a<��a<��a<t�a<��a<��a<�za<va<_ra<3pa<�oa<�pa<sa<�va<�{a<2�a<��a<��a<��a<��a<1�a<(�a<Βa<��a<�a<��a<�a<=~a<Lza<wa</ua<lta<�ta<�va<ya<G|a<�a<܂a<��a<8�a<z�a<l�a<�a<�a<�za<�ta<Sna<�ga<�aa<]a<}Ya<NWa<�Va<#Xa<�Za<�^a<�ca<�ha< na<�ra<xva<ya<�ya<�ya<�wa<�ta<�pa<�la<�ga<�ca<m`a<�]a<�\a<�\a<%^a<�`a<�ca<�ga<�ka<oa<ra<�sa<.ta<Dsa<�pa<�la<ha<wba<�\a<Wa<�Qa<Na<�Ka<�Ja<}Ka<�Ma<�Qa<�Va<o\a<Eba<�  �  �da<�ja<�oa<8sa<nua<+va<�ua<�sa<&qa<Gna<&ka<mha<[fa<ea<ea<fa<Iha<-ka<�na<�ra<)va<hya<�{a<�|a<S|a<�za<Iwa<�ra<Qma<nga<�aa<�[a<pWa<,Ta<�Ra<�Ra<�Ta<�Xa<#^a<�da<�ka<.sa<Bza<��a<ƅa<��a<ۋa<��a<L�a<��a<b�a<��a<]�a<_�a<�a<xa<,�a<�a<ӄa<4�a<;�a<�a<�a<��a<ۘa<��a<��a<V�a<��a<x�a<��a<��a<C{a<�ua<:qa<na<�la<	ma</oa<sa<%xa<r~a<�a<��a<ϑa<*�a<7�a<ǝa<�a<��a<�a<�a<n�a<9�a<	�a<��a<��a<�a<W�a<�a<D�a<B�a<��a<�a<��a<!�a< �a<ğa<��a<��a<�a<6�a<ȉa<A�a<�|a<9wa<�ra<�oa<�na<�oa<Bra<Xva<�{a<�a<P�a<��a<W�a<�a<q�a<Q�a<��a<��a<��a<��a<:�a<��a<y�a<�a<$�a<��a<�a<��a<�a<�a<=�a<2�a<˙a<S�a<��a<��a<.�a<4�a<�a<��a<�a<b{a<�ta<�oa<�ka<ia<gha<�ia<�la<�pa<3va<a|a<u�a<_�a<z�a<s�a<��a<��a<t�a<��a<ɏa<�a<:�a<5�a<ɀa<�}a<|a<H{a<�{a<}a<a<��a<5�a<��a<g�a<��a<k�a<P�a<ʂa<�}a<�wa<�pa<�ia<^ba<�[a<|Va<kRa<1Pa<�Oa<1Qa<cTa<�Xa<\^a<\da<Kja<�oa<�ta<xa<za<�za<�ya<�wa<�ta<<qa<�ma<�ia<ga<�da<�ca<�ca<�da<�fa<�ia<�la<�oa<�ra<�ta<Qua<�ta<�ra<_oa<�ja<�da<8^a<�Wa<$Qa<�Ka<QGa<uDa<�Ca<VDa<Ga<RKa<�Pa<OWa<�]a<�  �  �aa<Lha<na<�ra<�ua<Xwa<�wa<�va<�ta<}ra<pa<�ma< la<9ka<-ka<!la<�ma<jpa<�sa<�va<�ya<�{a<}}a<�}a<�|a<�ya<�ua<[pa<)ja<�ca<�\a<�Va<�Qa<Na<`La<�La<�Na<�Ra<�Xa<�_a<�ga<�oa<|wa<�~a<��a<M�a<w�a<1�a<|�a<��a<L�a<`�a<i�a<a<��a<��a<]�a<�a<@�a<H�a<��a<�a<�a<>�a<y�a<;�a<��a<;�a<��a<ϊa<9�a<T}a<cva<ppa<Uka<�ga<^fa<�fa<ia<Xma<sa<�ya<�a<q�a<`�a<��a<M�a<�a<͟a<[�a<��a<ݝa<~�a<טa<;�a<�a<Òa<%�a<��a<��a<��a<9�a<�a<��a<ӟa<9�a<h�a<8�a<�a<C�a<ғa<>�a<%�a<�~a<�wa<�qa<�la<�ia<�ha<~ia<1la<�pa<�va<Y}a<��a<��a<#�a<��a<ݛa<��a<�a<Ɵa<Y�a<1�a<q�a<��a<Ɠa<��a<L�a<��a<&�a<]�a<L�a<ɕa<Y�a<��a<`�a<7�a<��a<�a<a�a<��a<��a<��a<*~a<�va<�oa<�ia<hea<�ba<'ba<`ca<�fa<xka<Nqa<xa<�~a<��a<��a<>�a<��a<��a<��a<�a<ƒa<��a<��a<A�a<,�a<�a<7�a<x�a<��a<��a<"�a<)�a<-�a<��a<��a<��a<�a<1�a<��a<|a< ua<Xma<lea<]a<�Va<�Pa<DLa<�Ia<�Ia<Ka<�Na<�Sa<�Ya<]`a<ga<ima<�ra<.wa<<za<�{a<�{a<Rza<#xa<Jua</ra<"oa<�la<�ja<�ia<�ia<�ja<Mla<�na< qa<�sa<oua<�va<�va<<ua<Zra<�ma<lha<�aa<�Za<*Sa<;La<1Fa<MAa<M>a<>=a<+>a<Aa<�Ea<�Ka<�Ra<3Za<�  �  !_a<�fa<�la<)ra<�ua<+xa<+ya<�xa<�wa<�ua<�sa<�qa<qpa<�oa<�oa<�pa<2ra<�ta<wa<�ya<J|a<�}a<�~a<M~a<�|a<ya<eta<sna<�ga<n`a<6Ya<�Ra<>Ma<�Ia<�Ga<�Ga<eJa<tNa<�Ta<\a<Nda<�la<Tua<}a<��a<�a<ˌa<T�a</�a<�a<H�a<��a<^�a<��a<3�a<�a<Ȋa<P�a<��a<P�a<�a<�a<e�a< �a<��a<��a<e�a<X�a<.�a<��a<��a<za<�ra<<la<�fa<{ca<�aa<ba<�da<�ha<�na<
va<�}a<ޅa<c�a<�a<��a<�a<]�a<��a<l�a<l�a<��a<`�a<R�a<h�a<1�a<��a<��a<�a<əa<�a<1�a<��a<��a<آa<S�a<h�a<�a</�a<!�a<�a<E�a<T{a<�sa<qma<gha<Nea<�ca<�da<�ga<gla<�ra<�ya<��a<?�a<d�a<��a<b�a<͞a<��a<V�a<j�a<�a<��a<L�a<�a<�a<ʔa<'�a<��a<��a<h�a<d�a<u�a<U�a<G�a<��a<Z�a<�a<��a<R�a<��a<�a<{a<sa<�ka<rea<�`a<0^a<n]a<�^a<ba<3ga<�ma<�ta<E|a<o�a<�a<K�a<x�a<�a<�a<��a<�a<��a<�a<6�a<e�a<.�a<��a<�a<��a<Æa<*�a<��a<5�a<#�a<l�a<֋a<~�a<
�a<̀a<|za<�ra<�ja<ba<�Ya<fRa<La<�Ga<8Ea<�Da<�Fa<Ja<�Oa<�Ua</]a<�da<lka<�qa<rva<7za<&|a<}a<-|a<�za<`xa<�ua<8sa<�pa<Eoa<Cna<Rna<
oa<wpa<nra<Kta<mva<�wa<<xa<�wa<lua<�qa<�la<�fa<q_a<�Wa<�Oa<\Ha<�Aa<�<a<�9a<}8a<�9a<�<a<cAa<�Ga<COa<FWa<�  �  �]a<fea<]la<�qa<va<�xa<za<za<Bya<�wa<va<vta<;sa<�ra<�ra<xsa<ua<�va<Vya<�{a<�}a<6a<�a<�~a<�|a<�xa<�sa<6ma<fa<j^a<Wa<:Pa<�Ja<�Fa<�Da<�Da<'Ga<�Ka<�Qa<�Ya<<ba<7ka<�sa<|a<6�a<߈a<�a<ŏa<A�a<��a<��a<�a<��a<��a<�a<�a<ƍa<-�a<F�a<��a<O�a<Ҙa<��a<$�a</�a<�a<;�a<��a<=�a<_�a<�a<�wa<rpa<�ia<7da<F`a<s^a<�^a<�aa<9fa<_la<�sa<�{a<>�a< �a<Q�a<@�a<ȝa<��a<d�a<��a<�a<i�a<��a<a<9�a<�a<��a<��a<ښa<j�a<\�a<M�a<;�a<q�a<��a<Ģa<��a<ќa<��a<�a<��a<^�a<9ya<�qa<�ja<�ea<ba<�`a<�aa<�da<�ia<>pa<�wa<�a<ɇa<<�a<�a<�a<�a<%�a<,�a<١a<��a<��a<��a<��a<Иa<��a<8�a<�a<z�a<�a<��a<Y�a<�a<��a<^�a<ĝa<�a<n�a<��a<f�a<��a<ya<�pa<Eia<�ba<�]a<�Za<<Za<�[a<f_a<�da<=ka<�ra<|za<�a<��a<�a<G�a<&�a<��a<��a<��a<��a<%�a<��a<$�a<�a<��a<�a<ڈa<��a<��a<ŋa<�a<��a<��a<Q�a<͉a<�a<m�a<�ya<�qa<�ha<`a<�Wa<�Oa<yIa<�Da<Ba<�Aa<�Ca<�Ga<�La<�Sa<![a<�ba<(ja<�pa< va<za<�|a<�}a<q}a<H|a<3za<�wa<�ua<�sa<)ra<Qqa<5qa<�qa<sa<�ta<gva<xa<ya<%ya<�wa<�ua<�qa<cla<�ea<
^a<�Ua<�Ma<�Ea</?a<:a<�6a<X5a<S6a<�9a<�>a<lEa<#Ma<VUa<�  �  =]a<�da<la<�qa<+va<�xa<Xza<�za<�ya<yxa<�va<Kua<ta<[sa<�sa<?ta<�ua<�wa<@za<d|a<]~a<�a<�a<a<�|a<�xa<Lsa<�la<�ea<�]a<GVa<EOa<�Ia<�Ea<�Ca<+Da<Fa<�Ja<�Pa<�Xa<aa<�ja<�sa<�{a<��a<��a<Z�a<�a<��a<�a<w�a<אa<}�a<��a<�a<�a<��a<�a<�a<t�a<H�a<a�a<~�a<��a<~�a<C�a<�a<��a<Սa<�a<?a<0wa<�oa<�ha<Mca< _a<�]a<1^a<m`a<Tea<aka<sa<'{a<Ãa<��a<��a<�a<��a<�a<��a<)�a<�a<�a<��a<��a<�a<ۚa<��a<��a<��a<A�a<-�a<(�a<��a<�a<�a<�a<Ƞa<��a<i�a<��a<�a<��a<wxa<�pa<�ia<�da<aa<O`a<�`a<�ca<�ha<Poa<�va<a<Z�a<ˎa<��a<�a<�a<x�a<��a<Z�a<�a<n�a<o�a<[�a<��a<q�a< �a<G�a<W�a<��a<��a<�a<i�a<�a<��a<�a<�a<=�a<9�a<��a<�a<\xa<#pa<Pha<�aa<�\a<0Za<�Ya<�Za<v^a<�ca<Zja<�qa<�ya<��a<��a<��a<�a<v�a<��a< �a<%�a<"�a<�a<U�a<�a<�a<u�a<��a<��a<O�a<N�a<��a<x�a<<�a<�a<��a<"�a<��a</�a<$ya<qa<_ha<I_a<�Va<�Na<�Ha<�Ca<sAa<�@a<pBa<�Fa<�Ka<�Ra<kZa<gba<�ia<jpa<�ua<
za<�|a<�}a<�}a<�|a<�za<�xa<wva<�ta<�ra<5ra<ra<�ra<�sa<�ua<Bwa<�xa<�ya<|ya<Hxa<�ua<�qa<"la<,ea<�]a<'Ua<�La<Ea<2>a<9a<�5a<�4a<o5a<�8a<�=a<~Da<\La<�Ta<�  �  �]a<fea<]la<�qa<va<�xa<za<za<Bya<�wa<va<vta<;sa<�ra<�ra<xsa<ua<�va<Vya<�{a<�}a<6a<�a<�~a<�|a<�xa<�sa<6ma<fa<j^a<Wa<:Pa<�Ja<�Fa<�Da<�Da<'Ga<�Ka<�Qa<�Ya<<ba<7ka<�sa<|a<6�a<߈a<�a<ŏa<A�a<��a<��a<�a<��a<��a<�a<�a<ƍa<-�a<F�a<��a<O�a<Ҙa<��a<$�a</�a<�a<;�a<��a<=�a<_�a<�a<�wa<rpa<�ia<7da<F`a<s^a<�^a<�aa<9fa<_la<�sa<�{a<>�a< �a<Q�a<@�a<ȝa<��a<d�a<��a<�a<i�a<��a<a<9�a<�a<��a<��a<ښa<j�a<\�a<M�a<;�a<q�a<��a<Ģa<��a<ќa<��a<�a<��a<^�a<9ya<�qa<�ja<�ea<ba<�`a<�aa<�da<�ia<>pa<�wa<�a<ɇa<<�a<�a<�a<�a<%�a<,�a<١a<��a<��a<��a<��a<Иa<��a<8�a<�a<z�a<�a<��a<Y�a<�a<��a<^�a<ĝa<�a<n�a<��a<f�a<��a<ya<�pa<Eia<�ba<�]a<�Za<<Za<�[a<f_a<�da<=ka<�ra<|za<�a<��a<�a<G�a<&�a<��a<��a<��a<��a<%�a<��a<$�a<�a<��a<�a<ڈa<��a<��a<ŋa<�a<��a<��a<Q�a<͉a<�a<m�a<�ya<�qa<�ha<`a<�Wa<�Oa<yIa<�Da<Ba<�Aa<�Ca<�Ga<�La<�Sa<![a<�ba<(ja<�pa< va<za<�|a<�}a<q}a<H|a<3za<�wa<�ua<�sa<)ra<Qqa<5qa<�qa<sa<�ta<gva<xa<ya<%ya<�wa<�ua<�qa<cla<�ea<
^a<�Ua<�Ma<�Ea</?a<:a<�6a<X5a<S6a<�9a<�>a<lEa<#Ma<VUa<�  �  !_a<�fa<�la<)ra<�ua<+xa<+ya<�xa<�wa<�ua<�sa<�qa<qpa<�oa<�oa<�pa<2ra<�ta<wa<�ya<J|a<�}a<�~a<M~a<�|a<ya<eta<sna<�ga<n`a<6Ya<�Ra<>Ma<�Ia<�Ga<�Ga<eJa<tNa<�Ta<\a<Nda<�la<Tua<}a<��a<�a<ˌa<T�a</�a<�a<H�a<��a<^�a<��a<3�a<�a<Ȋa<P�a<��a<P�a<�a<�a<e�a< �a<��a<��a<e�a<X�a<.�a<��a<��a<za<�ra<<la<�fa<{ca<�aa<ba<�da<�ha<�na<
va<�}a<ޅa<c�a<�a<��a<�a<]�a<��a<l�a<l�a<��a<`�a<R�a<h�a<1�a<��a<��a<�a<əa<�a<1�a<��a<��a<آa<S�a<h�a<�a</�a<!�a<�a<E�a<T{a<�sa<qma<gha<Nea<�ca<�da<�ga<gla<�ra<�ya<��a<?�a<d�a<��a<b�a<͞a<��a<V�a<j�a<�a<��a<L�a<�a<�a<ʔa<'�a<��a<��a<h�a<d�a<u�a<U�a<G�a<��a<Z�a<�a<��a<R�a<��a<�a<{a<sa<�ka<rea<�`a<0^a<n]a<�^a<ba<3ga<�ma<�ta<E|a<o�a<�a<K�a<x�a<�a<�a<��a<�a<��a<�a<6�a<e�a<.�a<��a<�a<��a<Æa<*�a<��a<5�a<#�a<l�a<֋a<~�a<
�a<̀a<|za<�ra<�ja<ba<�Ya<fRa<La<�Ga<8Ea<�Da<�Fa<Ja<�Oa<�Ua</]a<�da<lka<�qa<rva<7za<&|a<}a<-|a<�za<`xa<�ua<8sa<�pa<Eoa<Cna<Rna<
oa<wpa<nra<Kta<mva<�wa<<xa<�wa<lua<�qa<�la<�fa<q_a<�Wa<�Oa<\Ha<�Aa<�<a<�9a<}8a<�9a<�<a<cAa<�Ga<COa<FWa<�  �  �aa<Lha<na<�ra<�ua<Xwa<�wa<�va<�ta<}ra<pa<�ma< la<9ka<-ka<!la<�ma<jpa<�sa<�va<�ya<�{a<}}a<�}a<�|a<�ya<�ua<[pa<)ja<�ca<�\a<�Va<�Qa<Na<`La<�La<�Na<�Ra<�Xa<�_a<�ga<�oa<|wa<�~a<��a<M�a<w�a<1�a<|�a<��a<L�a<`�a<i�a<a<��a<��a<]�a<�a<@�a<H�a<��a<�a<�a<>�a<y�a<;�a<��a<;�a<��a<ϊa<9�a<T}a<cva<ppa<Uka<�ga<^fa<�fa<ia<Xma<sa<�ya<�a<q�a<`�a<��a<M�a<�a<͟a<[�a<��a<ݝa<~�a<טa<;�a<�a<Òa<%�a<��a<��a<��a<9�a<�a<��a<ӟa<9�a<h�a<8�a<�a<C�a<ғa<>�a<%�a<�~a<�wa<�qa<�la<�ia<�ha<~ia<1la<�pa<�va<Y}a<��a<��a<#�a<��a<ݛa<��a<�a<Ɵa<Y�a<1�a<q�a<��a<Ɠa<��a<L�a<��a<&�a<]�a<L�a<ɕa<Y�a<��a<`�a<7�a<��a<�a<a�a<��a<��a<��a<*~a<�va<�oa<�ia<hea<�ba<'ba<`ca<�fa<xka<Nqa<xa<�~a<��a<��a<>�a<��a<��a<��a<�a<ƒa<��a<��a<A�a<,�a<�a<7�a<x�a<��a<��a<"�a<)�a<-�a<��a<��a<��a<�a<1�a<��a<|a< ua<Xma<lea<]a<�Va<�Pa<DLa<�Ia<�Ia<Ka<�Na<�Sa<�Ya<]`a<ga<ima<�ra<.wa<<za<�{a<�{a<Rza<#xa<Jua</ra<"oa<�la<�ja<�ia<�ia<�ja<Mla<�na< qa<�sa<oua<�va<�va<<ua<Zra<�ma<lha<�aa<�Za<*Sa<;La<1Fa<MAa<M>a<>=a<+>a<Aa<�Ea<�Ka<�Ra<3Za<�  �  �da<�ja<�oa<8sa<nua<+va<�ua<�sa<&qa<Gna<&ka<mha<[fa<ea<ea<fa<Iha<-ka<�na<�ra<)va<hya<�{a<�|a<S|a<�za<Iwa<�ra<Qma<nga<�aa<�[a<pWa<,Ta<�Ra<�Ra<�Ta<�Xa<#^a<�da<�ka<.sa<Bza<��a<ƅa<��a<ۋa<��a<L�a<��a<b�a<��a<]�a<_�a<�a<xa<,�a<�a<ӄa<4�a<;�a<�a<�a<��a<ۘa<��a<��a<V�a<��a<x�a<��a<��a<C{a<�ua<:qa<na<�la<	ma</oa<sa<%xa<r~a<�a<��a<ϑa<*�a<7�a<ǝa<�a<��a<�a<�a<n�a<9�a<	�a<��a<��a<�a<W�a<�a<D�a<B�a<��a<�a<��a<!�a< �a<ğa<��a<��a<�a<6�a<ȉa<A�a<�|a<9wa<�ra<�oa<�na<�oa<Bra<Xva<�{a<�a<P�a<��a<W�a<�a<q�a<Q�a<��a<��a<��a<��a<:�a<��a<y�a<�a<$�a<��a<�a<��a<�a<�a<=�a<2�a<˙a<S�a<��a<��a<.�a<4�a<�a<��a<�a<b{a<�ta<�oa<�ka<ia<gha<�ia<�la<�pa<3va<a|a<u�a<_�a<z�a<s�a<��a<��a<t�a<��a<ɏa<�a<:�a<5�a<ɀa<�}a<|a<H{a<�{a<}a<a<��a<5�a<��a<g�a<��a<k�a<P�a<ʂa<�}a<�wa<�pa<�ia<^ba<�[a<|Va<kRa<1Pa<�Oa<1Qa<cTa<�Xa<\^a<\da<Kja<�oa<�ta<xa<za<�za<�ya<�wa<�ta<<qa<�ma<�ia<ga<�da<�ca<�ca<�da<�fa<�ia<�la<�oa<�ra<�ta<Qua<�ta<�ra<_oa<�ja<�da<8^a<�Wa<$Qa<�Ka<QGa<uDa<�Ca<VDa<Ga<RKa<�Pa<OWa<�]a<�  �  	ha<ma<qa<�sa<�ta<�ta<4sa<tpa<ma<3ia<^ea<#ba<�_a<E^a<^a<A_a<�aa<�da<%ia<�ma<1ra<>va<�ya<{{a<|a<[{a<ya<�ua<qa<�ka<�fa<�aa<�]a<[a<�Ya<Za<\a<�_a<jda<ija<�pa<Fwa<�}a<Ȃa< �a<ȉa<
�a<�a<��a<�a<
�a<��a<d}a<�za<ya<�xa<Qya<&{a<E~a<2�a<҆a<��a<�a<�a<�a<��a<ɘa<z�a<��a<��a<��a<<�a<�a<�{a<�wa<ua<�sa<(ta<!va<�ya<A~a<׃a<��a<|�a<Ôa<�a<$�a<��a<̝a<��a<�a<��a<��a<��a<�a<�a<��a<�a<��a<#�a<�a<i�a<��a<Õa<}�a<��a<��a<,�a<k�a<�a<d�a<��a<	�a<O�a<��a<�}a<�ya<)wa<!va<�va<ya<�|a<��a<�a<��a<)�a<�a<��a<�a<֝a<L�a<^�a<:�a<m�a<%�a<ߋa<.�a<6�a<U�a<��a<B�a<�a<؇a<j�a<`�a<8�a<��a<=�a<��a<m�a<��a<��a<��a<t�a<��a<��a<�za<va<_ra<3pa<�oa<�pa<sa<�va<�{a<2�a<��a<��a<��a<��a<1�a<(�a<Βa<��a<�a<��a<�a<=~a<Lza<wa</ua<lta<�ta<�va<ya<G|a<�a<܂a<��a<8�a<z�a<l�a<�a<�a<�za<�ta<Sna<�ga<�aa<]a<}Ya<NWa<�Va<#Xa<�Za<�^a<�ca<�ha< na<�ra<xva<ya<�ya<�ya<�wa<�ta<�pa<�la<�ga<�ca<m`a<�]a<�\a<�\a<%^a<�`a<�ca<�ga<�ka<oa<ra<�sa<.ta<Dsa<�pa<�la<ha<wba<�\a<Wa<�Qa<Na<�Ka<�Ja<}Ka<�Ma<�Qa<�Va<o\a<Eba<�  �  �ka<�oa<�ra<Zta<�ta<#sa<�pa<�la<}ha<�ca<?_a<Y[a<TXa<�Va<eVa<�Wa<aZa<_^a< ca<gha<�ma<�ra<wa<za<�{a<|a<�za<oxa<�ta<�pa<\la<Zha<�da<oba<aaa<�aa<�ca<�fa</ka<Qpa<�ua<�{a<΀a<.�a<8�a<�a<3�a<�a<��a<�a<&a<�za<wa<�sa<�qa<�pa<�qa<�sa<7wa<�{a<��a<��a<�a<�a<�a<��a<�a<��a<�a<ӓa<�a<b�a<��a<��a<�~a<�|a<c{a<�{a<�}a<��a<ʄa<y�a<��a<z�a<��a<�a<��a<��a<��a<J�a<��a<Y�a<y�a<��a<]�a<��a<|~a<[}a<�}a<�a<�a<>�a<�a<�a<ʕa<�a<�a<��a<ܞa<��a<��a<)�a<��a<��a<Ɉa<u�a<�a<�~a<�}a<n~a<U�a<��a<ɇa<i�a<_�a<ѕa<��a<4�a<��a<d�a<��a<��a<��a<ۏa<��a<��a<c�a<�}a<�{a<�za<�{a<�}a<;�a<c�a<�a<��a<3�a<іa<�a<8�a<��a<ӗa<��a<W�a<~�a<7�a<e�a<!}a<�ya<�wa<)wa<+xa<Oza<�}a<Ӂa<d�a<�a<�a<�a<�a<l�a<R�a<ѐa<��a<.�a<Ԃa< }a<�wa<Rsa<�oa<�ma<�la<ma<yoa<�ra<qva<�za<�~a<o�a<!�a<��a<��a<�a<-�a<~a<�xa<xsa<�ma<�ha<1da<�`a<�^a<�^a<�_a<�aa<_ea<cia<�ma<ra<�ua<zxa<�ya<�ya<Yxa<�ua<{qa<�la<Jga<ba<H]a<?Ya<�Va<Ua<MUa<�Va<�Ya<�]a<ba<�fa<gka<Hoa<ra<�sa<�sa<;ra<�oa<�ka<ga<�aa<$]a<�Xa<IUa<1Sa<@Ra<Sa<!Ua<�Xa<�\a<�aa<�fa<�  �  Foa<`ra<<ta<�ta<�sa<�qa<�ma<ia<�ca<H^a<�Xa<`Ta<�Pa<"Oa<�Na<APa<!Sa<�Wa<]a<"ca<Oia<Voa<�ta<�xa<�{a<�|a<�|a<<{a<�xa<�ua<ra<�na<�ka<�ia<�ha<Zia<�ja<�ma<�qa<Ava<${a<�a<�a<k�a<c�a<�a<L�a<�a<��a<a<za<.ua<�pa<�la<[ja<]ia<�ia<Zla<pa<&ua<6{a<��a<�a<�a<˒a<��a<טa<��a<�a<�a<�a<q�a<��a<��a<	�a<�a<�a<l�a<�a<��a<�a<1�a<}�a<Q�a<��a<�a<a<J�a<B�a<՗a<U�a<�a<@�a<��a<�}a<�ya<�va<�ua<Rva<ixa<|a<؀a<y�a<5�a<��a<�a<�a<�a<"�a<��a<{�a<��a<	�a<��a<؎a<�a<*�a<6�a<r�a<�a<��a<g�a<�a<�a<�a<h�a<9�a<ȝa<��a<ʜa<
�a<��a<�a<�a<8�a<sa<gza<�va</ta<Vsa<>ta<�va<`za<Pa<Ƅa<Q�a<��a<@�a<��a<ՙa<\�a<��a<g�a<�a<3�a<܋a<��a<�a<�a<la<�~a<�a<v�a<>�a<ća<��a<�a<*�a<V�a<�a<s�a<j�a<��a<��a<"�a<�}a<rwa<^qa<3la<Wha<�ea<ea<fa<Qha<�ka<�pa<�ua<�za<Ma<�a<|�a<y�a<�a<O�a<"�a<}a<�xa<�sa<oa<Hka<Oha<�fa</fa<�fa<�ha<�ka<oa<�ra<�ua<�xa<iza<�za<�ya<wa<sa<na<4ha<ba<\a<|Va<Ra<Oa<wMa<�Ma<oOa<�Ra<>Wa<�\a<ba<�ga<rla<Mpa<�ra<�sa<�sa<ra<!oa<tka<[ga<1ca<x_a<�\a<�Za<�Ya<�Za<o\a<[_a<	ca<Cga<�ka<�  �  �ra<�ta<�ua<)ua<Csa<�oa<-ka<�ea<X_a<Ya<�Ra<Na<8Ja<�Ga<�Ga<Ia<vLa<1Qa<9Wa<$^a<ea<�ka<(ra<Uwa<{a<a}a<>~a<�}a<6|a<�ya<<wa<nta<+ra<�pa<�oa<Fpa<�qa<�ta<�wa<�{a<�a<��a<�a<V�a<{�a<�a<O�a<�a<��a<+{a<ua<�oa<bja<Ofa<_ca<?ba<�ba<Oea<�ia<�na<�ua<�|a<�a<Ɗa<ǐa<��a<ɘa<��a<ךa<�a<Ǘa<��a<�a<�a<��a<Ȋa<��a<>�a<��a<�a<��a<��a<ȗa<��a<]�a<��a<��a<��a<��a<��a<�a<Ɖa<a�a<�|a<Awa<�ra<�oa<�na<+oa<�qa<�ua<�za<7�a<Ňa<M�a<F�a<g�a<)�a<o�a<?�a<��a<ݝa<
�a<�a<��a<W�a<ڎa<�a<k�a<��a<Z�a<��a<��a<�a<��a<��a<��a<#�a<c�a<&�a<r�a<U�a<U�a<��a<�a<vya<
ta<�oa<ma<+la<ma<�oa<	ta<xya<�a<�a<X�a<ڑa<Y�a<m�a<�a<%�a<��a<��a<h�a<�a<x�a<`�a<�a<<�a<΅a<b�a<�a<Z�a<P�a<7�a<��a<5�a<C�a<+�a<��a<o�a<،a<�a<>�a<-ya<�qa<;ka<�ea<Zaa<�^a<�]a<�^a<�aa<�ea<ka<�pa<�va</|a<�a<f�a<j�a<�a<!�a<�a<�a<
}a<#ya<'ua<�qa<)oa<�ma<ma<�ma<Xoa<�qa<jta<wa<�ya<i{a<|a<h{a<Vya<�ua<�pa<�ja<da<5]a<PVa<0Pa<kKa<�Ga<SFa<�Fa<�Ha<ULa<5Qa<UWa<�]a<�ca<�ia<�na<*ra<Gta<�ta<4ta<Zra<toa<Fla<�ha<�ea<:ca<taa<�`a<caa<"ca<�ea<�ha<Lla<�oa<�  �  Jua<�va<�va<zua<�ra<mna<�ha<�ba<�[a<~Ta<Na<wHa<$Da<�Aa<eAa<�Ba<vFa<�Ka<RRa<�Ya<�aa<ia<pa<�ua<�za<�}a<�a<�a<a<�}a<�{a<kya<�wa<mva<�ua<eva<�wa<�ya<�|a<]�a<ԃa<�a<}�a<�a<L�a<)�a<W�a<d�a<~a<�wa<vqa<�ja<Gea<�`a<?]a<�[a<�\a<,_a<�ca<�ia<�pa<�xa<��a<-�a<�a<|�a<��a<W�a<��a<6�a<�a<�a<��a<�a<�a<ϐa<%�a<r�a<��a<o�a<�a<�a<��a<�a<��a<�a<�a<��a<��a<��a<5�a<C�a<a<xa<�qa<�la<�ia<Wha<�ha<{ka<�oa<�ua<}|a<�a<+�a<��a<ݗa<h�a<��a<E�a<��a<|�a<��a<	�a<I�a<��a<��a<�a<��a<�a<�a<��a<|�a< �a<��a<m�a<��a<D�a<��a<��a<��a<�a<E�a<�a<l{a<�ta<|na<�ia<�fa<�ea<�fa<�ia<�na<�ta<U{a<��a<i�a<̏a<��a<�a<��a<|�a<�a<��a<<�a<c�a<v�a<��a<ōa<g�a<�a<k�a<��a<��a<�a<@�a<L�a<��a< �a<��a<��a<w�a<0�a<v�a<}a<%ua<'ma< fa<�_a<;[a<�Xa<�Wa<�Xa<�[a<�`a<<fa<�la<[sa<�ya</a<V�a<\�a<Ǉa<ʇa<c�a<�a<�a<�}a<?za<Pwa</ua<�sa<4sa<�sa<�ta<�va<�xa<�za<�|a<�}a<{}a<�{a<	ya<�ta<�na<ha<�`a<�Xa<kQa<�Ja<sEa<�Aa<@a<R@a<�Ba<�Fa<6La<�Ra<�Ya<�`a<Zga<ma<hqa<�ta<�ua<"va<�ta<�ra<epa<�ma<�ja<�ha<�ga<	ga<�ga<�ha<�ja<�ma<{pa<-sa<�  �  Qwa<2xa<~wa<�ua<ra<?ma<(ga<`a<�Xa<�Pa<Ja<Da<�?a<7=a<�<a<u>a<�Aa<Ga<zNa<HVa<�^a<�fa<sna<�ta<Qza<~a<��a<��a<C�a<{�a<�~a<F}a<�{a<�za<lza<�za<=|a<G~a<�a<܃a<�a<��a<Q�a<m�a<Ћa<�a<��a<�a<�{a<Uua<=na<Gga<+aa<�[a<�Xa<LWa<�Wa<�Za<(_a<�ea<ma<uua<�}a<�a<��a<��a<��a<śa<ȝa<��a<_�a<�a<��a<*�a<Y�a<#�a<��a<�a<�a<��a<�a<!�a<��a<.�a<3�a<�a<_�a<f�a<��a<�a<�a<��a<�{a<>ta<�ma<gha<6ea<�ca<Tda<ga<}ka<�qa<�xa<ڀa<��a<�a<��a<Лa<��a<��a<�a<m�a<H�a<)�a<�a<��a<јa<��a<�a<c�a<i�a<�a<4�a<B�a<^�a<u�a<�a<�a<Ϟa<��a<ƕa<O�a<ۇa<�a<�wa<�pa<ja<;ea<?ba<&aa<mba<bea<Sja<�pa<�wa<�a<$�a<#�a<�a<��a<��a<u�a<��a<��a<�a<��a<Q�a<�a<�a<��a<\�a<Ґa<��a<��a<a�a<T�a<Ϙa<r�a<Z�a<��a<��a<��a<��a<q�a<hza<�qa<�ia<ba<c[a<�Va<�Sa<Sa<vTa<iWa<}\a<�ba<�ia<�pa<�wa<�}a<{�a<?�a<5�a<�a<*�a<y�a<�a<�a<O~a<�{a<�ya<xa<�wa<�wa<�xa<�za<|a<�}a<�~a<?a<�~a<F|a<�xa<�sa<Nma<�ea<�]a<vUa<�Ma<�Fa<�@a<U=a<X;a<�;a<>a<2Ba<7Ha<Oa<�Va<P^a<~ea<�ka<�pa<�ta<�va<�wa<�va<�ua<�sa<Cqa<oa</ma<la<uka<la<.ma<oa<Vqa<�sa<�ua<�  �  �xa<�xa<�wa<�ua<�qa<�la<�ea<�^a<�Va<�Na<�Ga<bAa<�<a<�9a<}9a<-;a<;?a<�Da<La<1Ta<�\a<iea<[ma<rta<za<K~a<��a<��a<ǂa<#�a<݀a<�a<[~a<�}a<T}a<�}a<a<�a<p�a<�a<��a<�a<��a<�a<.�a<��a<<�a<�a<�za<�sa<,la<ea<�^a<cYa<�Ua<Ta<�Ta<�Wa<�\a<�ba<�ja<^sa<H|a<ʄa<��a<E�a<z�a<�a<L�a<*�a<��a<��a<4�a<��a< �a<�a<��a<ӗa<Ęa<^�a<N�a<S�a<K�a<��a<:�a<��a<��a<0�a<O�a<��a<��a<��a<�ya<�qa<ka<�ea<�aa<l`a<aa<da<�ha<Boa<�va<�~a<+�a<�a<ܕa<��a<��a<a�a<ƣa<ɣa<�a<�a<-�a<<�a<��a<v�a<�a<=�a<4�a<��a<{�a<=�a<��a<ޢa<ڢa<y�a<�a<��a<!�a<!�a<a�a<�}a<�ua<na<fga<\ba<�^a<�]a<$_a<�ba<�ga<Ona<�ua<�}a<��a<
�a<u�a<c�a<�a<�a<��a<1�a<ǜa<��a<��a<��a<��a<ɓa<g�a<��a<��a<�a<��a<!�a<g�a<��a<��a<��a<i�a<]�a<�a<*�a<�xa<�oa<bga<e_a<�Xa<�Sa<�Pa<�Oa<EQa<�Ta<�Ya<Y`a<sga<oa<2va<�|a<�a<�a<��a<��a<V�a<�a<υa<K�a<��a<]~a<`|a< {a<�za<�za<�{a<�|a<>~a<�a<d�a<G�a<�~a<|a<�xa<!sa<Dla<wda< \a<dSa<IKa<�Ca<D>a<:a<*8a<u8a<";a<�?a<�Ea<�La<�Ta<�\a<Eda<ka<�pa<�ta<wa<Xxa<Bxa<Hwa<pua<�sa<�qa<�oa<�na<�na<�na<�oa<�qa<�sa<�ua<�wa<�  �  va<Xva<�ua<�sa<�pa<�la<�ga<Mba<?\a<QVa<�Pa<NLa<�Ha<Ga<�Fa<Ha<)Ka<[Oa<�Ta<0[a<�aa<�ha<�na<*ta<|xa<|a<w~a<�a<�a<�a<Ia<g~a<�}a<-}a<)}a<�}a<�~a<��a<S�a<��a<��a<]�a<��a<�a<~�a<��a<	�a<C�a<�|a<�wa<�qa<�la<�ga<,da<�aa<�`a<faa<�ca<Xga<Cla<�ra<�xa<�a<��a<��a<ˑa<ҕa<�a<�a<��a<��a<�a<�a<Řa<�a<��a<�a<�a<ɗa<�a<��a<2�a<�a<}�a<Ԟa<`�a<˜a<�a<L�a<��a<��a<�a<�a<za<�ta<�pa<na<*ma<�ma<�oa<Usa<xa<�}a<�a<m�a<4�a<��a<��a<�a<o�a<v�a<{�a<�a<מa<n�a<֛a<��a<��a<��a<��a<c�a<R�a<��a<�a<�a<��a<��a<��a<A�a<֘a<��a<H�a<w�a<�a<�|a<�va<�qa<�ma<zka<�ja<xka<na<�qa<�va<C|a<h�a<b�a<Ӎa<��a<H�a<7�a<ךa<Z�a<��a<��a<��a<�a<U�a<��a<�a<֒a<ǒa<��a<f�a<��a<��a<3�a<I�a<��a<͔a<͑a<׍a<ǈa<ɂa<l|a<Wua<�na<�ha<�ca<�_a<[]a<�\a<X]a<�_a<Xca<Fha<Zma<)sa<Rxa<%}a<�a<�a<�a<��a<d�a<Q�a<��a<ˁa<�a<�}a< |a<{a<zza<lza<{a<�{a<�|a<a}a<�}a<{}a<q|a<Kza<�va<�ra<fma<aga<�`a<%Za<Ta<MNa<Ja<�Fa<�Ea<�Ea<dGa<�Ja<"Oa<�Ta<�Za<�`a<<fa<]ka<hoa<�ra<�ta<�ua<�ua<�ta<�sa<pra<�pa<�oa<�na<�na<�na<�oa<�pa<�ra<ta<Lua<�  �  �ua<va<\ua<�sa<�pa<�la< ha<qba<�\a<�Va<�Qa<Ma<�Ia<�Ga<oGa<�Ha<�Ka<#Pa<�Ua<�[a<Oba<�ha<�na<Lta<�xa<|a<A~a<�a<�a<�a<�~a<�}a<�|a<�|a<t|a<}a<~a<�a<��a<�a<*�a<�a<Y�a<�a<g�a<�a<-�a<��a<�|a<�wa<cra<Uma<�ha<�da<}ba<caa<ba<]da<ha<ma<%sa<�ya<W�a<ǆa<�a<�a<�a<�a<��a<g�a<\�a<��a<h�a<�a< �a<e�a< �a<]�a<2�a<[�a<ՙa<��a<#�a<?�a<��a<-�a<Ŝa<,�a<h�a<đa<)�a<Z�a<W�a<�za<�ua<�qa<�na<�ma<Rna<�pa<ta<�xa<�~a<{�a<��a<x�a<Õa<��a<>�a<9�a<B�a<A�a<��a<D�a<��a<!�a<��a<�a<Øa<ݘa<��a<��a<�a<~�a<Ȟa<W�a<W�a<I�a<T�a<�a<Ӕa<��a<��a<l�a<I}a<�wa<�ra<�na<8la<_ka<Fla<�na<jra<\wa<�|a<Âa<��a<�a<Ȓa<��a<7�a<��a<+�a<��a<��a<��a<<�a<��a<]�a<a�a<	�a<(�a<Ԓa<��a<��a<�a<�a<
�a<g�a<��a<��a<��a<�a<�a<�|a<�ua<{oa<`ia<Uda<{`a<�]a<7]a<0^a<�`a<&da<�ha<�ma<osa<�xa<u}a<:�a<-�a<߅a<��a<'�a<�a<?�a<�a<�~a< }a<h{a<Pza<�ya<�ya<Cza<
{a<|a<}a<�}a<L}a<>|a<Eza<wa<�ra<�ma<�ga<Baa<�Za<�Ta<Oa<�Ja<�Ga<Fa<QFa<=Ha<sKa<�Oa<BUa<�Za<�`a<�fa<�ka<�oa<�ra<�ta<ua<gua<�ta<Lsa<�qa<%pa<oa<(na<�ma<*na<oa<8pa<�qa<sa<ua<�  �  �ta<�ua<�ta<�sa<qa<ima<�ha<�ca<0^a<�Xa<[Sa<�Na<�Ka<Ja<�Ia<'Ka<�Ma<	Ra<QWa<e]a<�ca<�ia<�oa<�ta<�xa<�{a<�}a<�~a<�~a<!~a<}a<|a<�za<wza<Hza<�za<�{a<�}a<�a<f�a<��a<҆a<g�a<\�a<�a<�a<k�a<:�a<�}a<ya<ta<�na<|ja<�fa<�da<�ca<]da<�fa<�ia<�na<�ta<,{a<��a<҇a<��a<,�a<�a<��a<-�a<��a<�a<�a<ܗa<t�a<�a<M�a<�a<(�a<�a<a�a<@�a<��a<��a<�a<�a<��a<z�a<S�a<ǖa<��a<H�a<��a<�a<P|a<wwa<�sa<0qa<pa<�pa<�ra<�ua<�za<�a<�a<֋a<v�a<K�a<0�a<%�a<Ԟa<��a<6�a<J�a<��a<*�a<d�a<�a<�a<��a<��a<��a<Әa<}�a<�a<l�a<D�a<��a<�a<0�a<J�a<U�a<��a<Ҋa<�a<�~a<@ya<bta<�pa<�na<�ma<�na<�pa<Pta<ya<y~a<8�a<��a<�a<4�a<��a<��a<:�a<r�a<��a<@�a<n�a<��a<��a<H�a<5�a<Ϗa<�a<ɐa<�a<m�a<��a<��a<�a<ߕa<Y�a<��a<9�a<��a<�a<�}a<�wa<qa<Aka<4fa<�ba<V`a<�_a<\`a<qba<fa<qja<�oa<�ta<�ya<(~a<�a<<�a<��a<�a<D�a<̓a<Ɂa<�a<:}a<�za<Pya<xa<�wa<�wa<Ixa<vya<�za<�{a<I|a<�|a<�{a<�ya<Ewa<0sa<na<�ha<�ba<]\a<KVa<Qa<�La<�Ia<uHa<�Ha<JJa<OMa<�Qa<�Va<�\a<ba<~ga<!la<�oa<�ra</ta<�ta<[ta<^sa<�qa<-pa<ina<�la<la<�ka<la<ma<ona<Ipa<�qa<�sa<�  �  Usa<@ta<Uta<jsa<cqa<;na<&ja<rea<C`a<[a<]Va<]Ra<HOa<�Ma<AMa<�Na<\Qa<eUa<IZa<�_a<�ea<�ka<�pa<�ua<'ya<�{a<}a<p}a<"}a<|a<�za<)ya<�wa<wa<�va<�wa<�xa<�za<�|a<�a<`�a<�a<�a<E�a<��a<�a<�a<�a<Oa<�za<8va<�qa<�ma<Jja<ha<.ga<�ga<�ia<zma<-ra<�wa<r}a<��a<X�a<�a<�a<'�a<�a<#�a<#�a<h�a<ؖa<�a<i�a<�a<Ґa<��a<Аa<��a<<�a<E�a<e�a<��a<s�a<��a<ܜa<�a<y�a<��a<��a<�a<��a<X�a<<a<�za<wa<�ta<�sa<ta<va<lya<�}a<��a<(�a<��a<��a<%�a<��a<
�a<C�a<~�a<ʝa<_�a<[�a<B�a<A�a<��a<��a<C�a<P�a<B�a<��a<��a<��a<p�a<՜a<z�a<C�a<�a<��a<'�a<��a<��a<�a<r�a<C|a<�wa<>ta<�qa<3qa<�qa<7ta<�wa<�{a<��a<<�a<a�a<	�a<��a<��a<��a<n�a<�a<�a<'�a<�a<��a<��a<�a<Ռa<��a<��a<��a<�a<��a<R�a<�a<��a<ɔa<ߓa<��a<ގa<��a<��a<�a<�ya<�sa<ena<�ia<fa<�ca<ca<�ca<�ea<Bia<?ma<�qa<�va<({a<a<4�a<I�a<�a<��a<�a<�a<�a<�|a</za<�wa<�ua<�ta<6ta<Pta<%ua<zva<�wa<tya<�za<({a<�za<�ya<kwa<�sa<}oa<Pja<�da<�^a<7Ya<STa<6Pa<XMa<�Ka<La<�Ma<�Pa<�Ta<wYa<�^a<�ca<�ha<�la<Opa<�ra<�sa<�sa<�ra<tqa<doa<Fma<Gka<�ia<�ha<vha<�ha<�ia<Nka<Zma<�oa<�qa<�  �  ?qa<�ra<�sa<:sa<�qa<Toa<�ka<�ga<ca<�^a<Za<cVa<�Sa<"Ra<�Qa<$Sa<�Ua<IYa<�]a<2ca<{ha<�ma<xra<vva<jya<U{a<|a<�{a<�za<!ya<Mwa<sua<�sa<�ra<`ra<�ra<'ta<}va<	ya</|a<Ta<��a<�a<��a<�a<�a<��a<^�a<U�a<m}a<Eya<Fua<eqa<yna<�la<�ka<ula<�na<�qa<�ua<({a<��a<�a<l�a<׏a<��a<-�a<��a<�a<K�a<�a<֓a<��a<��a<�a<u�a<�a<D�a<^�a<Q�a<��a<�a<��a<+�a<��a<Λa<ܛa<��a<r�a<�a<&�a<g�a<��a<�a<�~a<d{a<.ya<>xa<�xa<�za<�}a<r�a<E�a<�a<�a<��a<Q�a<(�a<�a<��a<�a<śa<��a<5�a<��a<g�a<��a<�a<��a<юa<�a<ґa<�a<T�a<��a<��a<ݛa<t�a<֛a<�a<A�a<u�a<��a<މa<��a<�a<�{a<�xa<�va<�ua<�va<�xa<�{a<�a<H�a<�a<��a<��a<��a<8�a<o�a<u�a<c�a<ӕa<?�a<��a<��a<��a<��a<M�a<�a<5�a<��a<�a<4�a<F�a<V�a<͒a<s�a<]�a<�a<~�a<�a<��a<K�a<�|a<kwa<*ra<�ma<�ja<mha<�ga<Sha<+ja<ma<�pa<�ta<2ya<;}a<e�a<�a<N�a<��a<ăa<�a<�a<�|a<rya<[va<�sa<yqa<6pa<�oa<pa<:qa<�ra<�ta<�va<lxa<gya<�ya<Zya<�wa<�ta<�pa<�la<Mga<
ba<�\a<(Xa<�Ta<�Qa<�Pa<�Pa</Ra<�Ta<zXa<]a<�aa<Wfa<�ja<&na<�pa<dra<�ra<1ra<�pa<�na<@la<�ia<nga<�ea<$da<�ca<!da<�ea<pga<�ia<Xla<�na<�  �  �na<qa<�ra<�ra<<ra<�pa<�ma<cja<xfa<\ba<�^a<R[a<�Xa<uWa<>Wa<kXa<�Za<4^a<;ba<�fa<�ka<Cpa<\ta<qwa<�ya<�za<�za<�ya</xa<�ua<�sa<qa<�na<�ma<Bma<�ma<oa<Oqa<eta<xa<�{a<�a<܂a<��a<3�a<؇a<b�a<�a<��a<J�a<�|a<4ya<va<jsa<�qa<%qa<�qa<�sa<�va<�za<'a<)�a<�a<��a<z�a<]�a<5�a<�a<��a<(�a<��a<k�a<��a<��a<̈a<o�a<ˆa<�a<F�a<D�a<�a<=�a<c�a<S�a<��a<��a<;�a<ؚa<X�a<�a<~�a<��a<E�a<�a<��a<`�a<p~a<�}a<~a<�a<p�a<��a<�a<~�a<��a<��a<��a<��a<��a<��a<r�a<L�a<��a<��a<��a<��a<^�a<��a<[�a<a<�a<�a<��a<��a<��a<)�a<O�a<p�a<~�a<��a<o�a<x�a<��a<<�a<��a<r�a<Āa<�}a<�{a<2{a<�{a<�}a<�a<�a<��a<(�a<�a<��a<�a<�a<�a<K�a<��a<�a<�a<ٌa<��a<��a<|�a<.�a<��a<-�a<b�a<v�a<�a<Ƌa<Z�a<��a<	�a<��a<�a<.�a<c�a<��a<'�a<V�a<Z{a<�va<�ra<�oa<�ma<�la<�ma<oa<�qa<�ta<�xa<!|a<ra<�a<��a<W�a<��a<g�a<�a<�|a<ya<pua<�qa<�na<sla<�ja<�ja<�ja<-la<Ana<�pa<Esa<�ua<�wa<�xa<�xa<�wa<�ua<�ra<�na<ija<�ea<aa<]a<Ya<)Wa<�Ua<Va<IWa<�Ya<]a<�`a<�da<�ha<�la<koa<Oqa<+ra<�qa<�pa<tna<�ka<�ha<�ea<�ba<o`a<_a<�^a<_a<d`a<�ba<�ea<�ha<�ka<�  �  �ka<oa<:qa<�ra<�ra<�qa<�oa<ma<ja<tfa<7ca<k`a<1^a< ]a<�\a<^a<`a<@ca<�fa<�ja<#oa<�ra<&va<xa<"za<Uza<sya<�wa<;ua<xra<(oa<dla<�ia<;ha<�ga<�ga<�ia<la<�oa<�sa<xa<p|a<G�a<ƃa<@�a<�a< �a<Y�a<��a<K�a<��a<q}a<�za<�xa<Ewa<�va<rwa<Gya<�{a<�a<t�a<��a<+�a<�a<�a<)�a<h�a<�a<��a<��a<�a<��a<#�a<I�a<��a<�a<�a<o�a<Ђa<-�a<]�a<ʋa<Ϗa<W�a<��a<�a<��a<9�a<R�a<��a<�a<�a<<�a<��a<��a<��a<�a<5�a<��a<�a<��a<��a<5�a<,�a<��a<��a<��a<J�a<��a<f�a<��a<��a<d�a<��a<�a<��a<��a<d�a<��a<'�a<��a<
�a<�a<��a<F�a<[�a<I�a<&�a<F�a<�a<��a<t�a<:�a<ِa<Όa< �a<ޅa<*�a<��a<Ӏa<��a<�a<��a<y�a<��a<��a<��a<S�a< �a<�a<q�a<וa<k�a< �a<��a<|�a<�a<��a<
a<�}a<�|a<�}a<a<��a<��a<�a<C�a<��a<G�a<��a< �a<�a<ێa<�a<(�a<�a<�a<�{a<xa<Cua<nsa<�ra<sa<^ta<�va<0ya<b|a<Ea<��a<��a<~�a<��a<�a<��a<q}a<�ya<]ua<�pa<ma<lia<�fa<9ea<�da<tea<ga<�ia<Sla<�oa<�ra<@ua<wa<!xa<)xa<�va<�ta<Hqa<�ma<�ia<�ea<ba<�^a<�\a<�[a<�[a<�\a<�^a<�aa<�da<�ha<�ka<�na<�pa<�qa<ra<�pa<�na<�ka<|ha<�da<�`a<�]a<[a<�Ya<�Xa<zYa<�Za<�]a<�`a<�da<�ha<�  �  ?ia<"ma<pa<ra<sa<sa<�qa<�oa<kma<�ja<�ga<Zea<�ca<�ba<�ba<�ca<kea<ha<gka<�na<Wra<tua<xa<�ya<2za<�ya<xa<�ua<era<�na< ka<�ga<�da<�ba<�aa<Bba<�ca<�fa<�ja<oa<ta<ya<�}a<�a<S�a<��a<ƈa<�a<�a<J�a<4�a<�a<�a<�}a<�|a<�|a<0}a<�~a<$�a<U�a<�a<��a<.�a<R�a<��a<�a<&�a<=�a<L�a<]�a<��a<ψa<Ȅa<Z�a<E~a<K|a<`{a<�{a<C}a<�a<��a<��a<�a<g�a<q�a<��a<�a<0�a<U�a<p�a<��a<�a<�a<-�a<J�a<�a<��a< �a<_�a<��a<��a<h�a<��a<��a<u�a<՚a<J�a<��a<�a<K�a<��a<�a<�a<��a<N�a<��a<��a<�~a<�}a<z~a<�a<�a<e�a<p�a<��a<��a<Y�a<��a<��a<`�a<��a<��a<�a<1�a<�a<ʍa<ϊa<��a<8�a<��a<�a<L�a<^�a<�a<��a<Ғa<K�a<5�a<#�a<�a<Ȗa<��a<W�a<J�a<�a<U�a<�a<s|a<�ya<�wa<Bwa<�wa<�ya<�|a<�a<�a<�a<��a<��a<��a<��a<��a<j�a<4�a<&�a<��a<�a<h�a<+}a<�za<"ya<fxa<�xa<�ya<k{a<�}a<�a<G�a<#�a<6�a<B�a<I�a<7�a<%a< {a<qva<�qa<�la<#ha<'da<Paa<�_a<(_a<�_a<�aa<�da<ha<�ka<�oa<sa<�ua<lwa<xa<�wa<Ova<�sa<�pa<�ma<#ja<�fa<"da<Zba<Vaa<Zaa</ba<�ca<nfa<Eia<la<�na<�pa< ra<\ra<�qa<�oa<�la</ia<�da<�`a<X\a<�Xa<�Ua<�Sa<!Sa<�Sa<�Ua<�Xa<6\a<v`a<�da<�  �  �fa<%ka<�na<�qa<zsa<ta<�sa<�ra<�pa<Zna<&la<Cja<�ha<�ga<�ga<�ha<�ja<�la<�oa<tra<[ua<�wa<�ya<�za<]za< ya<�va<�sa<�oa<Uka<-ga<ca<�_a<�]a<�\a<�\a<�^a<�aa<�ea<�ja<qpa<va<�{a<U�a<w�a<u�a<s�a<.�a<�a<*�a<�a<υa<�a<ڂa<ҁa<��a<c�a<уa<@�a<��a<��a<�a<�a<d�a<��a<��a<�a<q�a<��a<�a<��a<6�a<��a<�|a<Rya<wa<va<kva<#xa<{a<�~a<��a<��a<��a<M�a<0�a<K�a<E�a<:�a<��a<ۚa<�a<��a<M�a<��a<7�a<��a<E�a<y�a<��a<��a<��a<H�a<a<'�a<��a<k�a<+�a<��a<E�a<��a<��a<��a<Їa< �a<�~a<�{a<mya<�xa<*ya<	{a<~a< �a<��a<[�a<2�a<[�a<חa<R�a<��a<�a< �a<��a<M�a<��a<�a<��a<a<J�a<�a<�a<{�a< �a<J�a<��a<ؕa<��a<��a<�a</�a<>�a<2�a<@�a<��a<u�a<��a<�{a<�wa<rta<�ra<�qa<�ra<�ta<�wa<�{a<`�a<�a<F�a<Ռa<Ïa<��a<>�a<��a<$�a<�a<�a<�a<�a<<�a<�a<J~a<�}a<�}a<�~a<�a<��a<w�a<5�a<5�a<��a<�a<8�a<k�a<t}a<�xa<vsa<�ma<vha<Xca<4_a<\a<@Za<�Ya<�Za<�\a<`a<6da<oha<�la<�pa<=ta<�va<2xa<�xa<�wa<9va<�sa<qa<Bna<}ka<Ria<dga<�fa<rfa<Yga<�ha<�ja<ma<>oa<gqa<�ra<Bsa<�ra<Aqa<�na<ka<�fa<�aa<�\a<Xa<�Sa<�Pa<�Na<�Ma<�Na<�Pa<�Sa<�Wa<�\a<�aa<�  �  ada<oia<�ma<[qa<�sa<�ta<2ua<�ta<Tsa<�qa<�oa<"na<�la<Nla<�la<$ma<�na<�pa<sa<�ua<xa<�ya< {a<7{a<zza<�xa<�ua<�qa<:ma<\ha<�ca<H_a<�[a<.Ya<�Wa<KXa<'Za<u]a<�aa<Ega<7ma<msa<jya<�~a<��a<Q�a<��a<E�a<��a<��a<s�a<%�a<�a<ǆa<$�a<?�a<��a<*�a<5�a<��a<X�a<
�a<��a<4�a<&�a<
�a<�a<��a<8�a<�a<+�a<�a<}a<�xa<ua<�ra<iqa<�qa<�sa<�va<{a<�a<��a<�a<Q�a<�a<��a<W�a<ǜa<E�a<˜a<��a<��a<��a<Еa<A�a<�a<�a< �a<�a<u�a<q�a<��a<��a<R�a<4�a<\�a<f�a<t�a<D�a<�a<A�a<�a<n�a<La<�za<:wa<�ta<�sa<�ta<�va<za<G~a<:�a<��a<ݍa<��a<Ŗa<��a<��a<�a<a<Лa<�a<�a<��a<��a<�a<̐a<��a<��a<��a<��a<ǔa<��a<��a<��a<1�a<��a<M�a<��a<��a<\�a<!�a<|�a<�|a<�wa<fsa<�oa<�ma<Kma<3na<�pa<ta<Hxa<&}a<?�a<�a<_�a<�a<_�a<��a<Œa<�a<\�a<�a<I�a<��a<)�a<"�a<قa<+�a<��a<��a<Ƀa<�a<s�a<��a<�a<��a<`�a<(�a<��a<|a<�va<�pa<�ja<�da<�_a<�Za<�Wa<�Ua</Ua<KVa<�Xa<R\a<�`a<hea<Vja<�na<�ra<.va<Dxa<*ya<#ya<(xa<zva<ta<�qa<Uoa<[ma<�ka<6ka<�ja<�ka<�la<vna<Epa<ra<�sa<=ta<2ta<sa<�pa<�ma<^ia<nda< _a<~Ya<XTa<�Oa<PLa<�Ia<&Ia<�Ia<!La<�Oa<Ta<CYa<�^a<�  �  �ba<Lha<ma<qa<�sa<�ua<zva<va<Wua< ta<�ra<Aqa<Fpa<�oa<�oa<�pa<�qa<�sa<�ua<�wa<�ya<C{a<,|a<�{a<�za<xa<�ta<kpa<hka<<fa<�`a<<\a<EXa<�Ua<�Ta<�Ta<�Va<�Ya<�^a<ada<�ja<rqa<�wa<�}a<قa<0�a<!�a<5�a<�a<�a<��a<ȋa<�a<�a<��a<��a<B�a<��a<_�a<��a<�a<E�a<6�a<��a<)�a<|�a<�a<�a<N�a<s�a<8�a<�a<Aza<�ua<�qa<oa<�ma<Vna<6pa<bsa<xa<]}a<Z�a<?�a<�a<�a<�a<`�a<G�a<b�a<0�a<h�a<	�a<��a<�a<y�a<��a<$�a<d�a<P�a<��a<g�a<�a<��a<͞a<��a<�a<��a<3�a<y�a<�a<��a<݇a<��a<O|a<twa<�sa<jqa<vpa<"qa<+sa<�va<E{a<��a<�a<�a<��a<��a<��a<(�a<��a<
�a<C�a<�a<]�a<��a<��a<D�a<4�a<ʓa<�a<Дa<�a<��a<�a<d�a<�a<^�a<H�a<d�a<1�a<"�a<�a<O�a<\�a<Jza<�ta<�oa<�la<tja<�ia<�ja<ma<�pa<cua<�za<D�a<x�a<g�a<#�a<>�a<�a<��a<N�a<��a<#�a<�a<��a<P�a<��a<,�a<x�a<x�a<Ӆa<φa<̇a<��a<Q�a<f�a<��a<҆a<�a<�a<){a<7ua<�na<mha<�aa<N\a<pWa<$Ta<%Ra<�Qa<�Ra<LUa<7Ya<�]a<<ca<ha<�ma< ra<�ua<Lxa<�ya<?za<�ya<Gxa<pva<�ta<tra<�pa<?oa<wna<[na<�na<�oa<kqa<�ra<0ta<ua<�ua<�ta<Tsa<�pa<�la<Pha<�ba<�\a<Wa<\Qa<�La<�Ha<�Fa<�Ea<zFa<�Ha<CLa<Qa<�Va<�\a<�  �  eaa<Uga<�la<�pa<ta<va<wa<.wa<�va<�ua<Nta<sa<^ra<�qa<ra<�ra<�sa<ua<�wa<rya<8{a<I|a<�|a<'|a<�za<�wa<.ta<moa<&ja<�da<\_a<kZa<jVa<�Sa<3Ra<qRa<�Ta<Xa<�\a<�ba<<ia<pa<�va<}a<��a<�a<p�a<��a<�a<W�a<�a<Q�a<{�a<�a<��a<ˋa<|�a<��a<h�a<M�a<��a<��a<s�a<o�a<��a<ϗa<ڕa<��a<��a<c�a<�a<~a<�xa<�sa<�oa<�la<�ka<�ka<na<�qa<%va<�{a<��a<��a<�a<t�a<ޗa<g�a<��a<�a<(�a<��a<��a<"�a<��a<��a<��a<^�a<��a<g�a<x�a<��a<��a<�a<��a<?�a<��a<�a<��a<�a<�a<]�a<d�a<X�a<�za<�ua<�qa<oa<na<�na<-qa<�ta<�ya<a<��a<�a<��a<x�a<i�a<S�a<�a<��a<]�a<�a<�a<;�a<��a<\�a<Y�a<	�a<"�a<��a<җa<>�a<��a<��a<$�a<�a<��a<w�a<��a<��a<�a<�a<�~a<�xa<�ra<na<uja<ha<pga<�ha<!ka<�na<�sa<*ya<�~a<_�a<��a<ˍa<�a<:�a<&�a<�a<2�a<��a<u�a<>�a<P�a<��a<d�a<��a<��a<ۇa<d�a<V�a< �a<��a<A�a<5�a<%�a<��a<�a<mza<'ta<�ma<�fa<j`a<eZa<�Ua<�Qa<�Oa<fOa<�Pa<pSa<ZWa<P\a<�aa<>ga<�la<�qa<Xua<Sxa<za<�za<�za<�ya<�wa<va<ta<�ra<Yqa<�pa<�pa<qa<�qa<sa<Vta<�ua<6va<Hva<Wua<�sa<�pa<gla<bga<�aa<�[a<jUa<�Oa<�Ja<�Fa<EDa<TCa<%Da<�Fa<`Ja<cOa<Ua<@[a<�  �  Faa<ga<[la<�pa<ta<?va<Uwa<lwa<�va<-va<�ta<�sa<sa<�ra<�ra<Qsa<�ta<3va<3xa<�ya<y{a<�|a<�|a<S|a<}za<�wa<�sa<'oa<�ia<*da<�^a<�Ya<�Ua<�Ra<�Qa<�Qa<�Sa<HWa<�[a<%ba<�ha<�oa<�va<�|a<j�a<цa<x�a<׌a<�a<��a<o�a<��a<*�a<��a<?�a<��a<=�a<N�a<1�a<�a<G�a<%�a<��a<��a<֘a<חa<��a<��a<E�a<$�a<��a<}a<xa<�ra<�na<la< ka<Yka<:ma<�pa<Xua<,{a<3�a<Ǉa<��a<)�a<��a<9�a<ŝa<�a<g�a<��a<�a<Μa<N�a<I�a<D�a<.�a<C�a<�a<3�a<��a<6�a<g�a<4�a<r�a<��a<�a<��a<ߖa<֑a<8�a<�a<�a<�ya<�ta< qa<Wna<�ma<
na<bpa<�sa<�xa<t~a<��a<��a<C�a<F�a<+�a<H�a<.�a<�a<��a<ǝa<��a<�a<A�a<�a<
�a<ؖa<Ėa<��a<��a<�a<�a<��a<]�a<�a<ٚa<Q�a<ʔa<S�a<ϊa<߄a<J~a<xa<#ra<Nma<�ia<rga<�fa<�ga<Yja<	na<&sa<�xa<�~a<-�a<V�a<��a<ސa<B�a<W�a<G�a<q�a<�a<"�a<�a<�a<=�a<�a<s�a<"�a<��a<�a<�a<��a<Њa<{�a<g�a<.�a<ăa<�a< za<�sa<Yma<3fa<�_a<�Ya<�Ta<Qa<3Oa<�Na<�Oa<�Ra<�Va<�[a<aa<ga<Jla<5qa<1ua<%xa<'za<�za<�za<�ya<qxa<�va<�ta<asa<�qa<�qa<:qa<�qa<�ra<�sa<�ta<�ua<tva<zva<�ua<�sa<?pa<@la<ga<faa<$[a<�Ta<Oa<�Ia<Fa<~Ca<�Ba<cCa<�Ea<�Ia<�Na<~Ta<�Za<�  �  eaa<Uga<�la<�pa<ta<va<wa<.wa<�va<�ua<Nta<sa<^ra<�qa<ra<�ra<�sa<ua<�wa<rya<8{a<I|a<�|a<'|a<�za<�wa<.ta<moa<&ja<�da<\_a<kZa<jVa<�Sa<3Ra<qRa<�Ta<Xa<�\a<�ba<<ia<pa<�va<}a<��a<�a<p�a<��a<�a<W�a<�a<Q�a<{�a<�a<��a<ˋa<|�a<��a<h�a<M�a<��a<��a<s�a<o�a<��a<ϗa<ڕa<��a<��a<c�a<�a<~a<�xa<�sa<�oa<�la<�ka<�ka<na<�qa<%va<�{a<��a<��a<�a<t�a<ޗa<g�a<��a<�a<(�a<��a<��a<"�a<��a<��a<��a<^�a<��a<g�a<x�a<��a<��a<�a<��a<?�a<��a<�a<��a<�a<�a<]�a<d�a<X�a<�za<�ua<�qa<oa<na<�na<-qa<�ta<�ya<a<��a<�a<��a<x�a<i�a<S�a<�a<��a<]�a<�a<�a<;�a<��a<\�a<Y�a<	�a<"�a<��a<җa<>�a<��a<��a<$�a<�a<��a<w�a<��a<��a<�a<�a<�~a<�xa<�ra<na<uja<ha<pga<�ha<!ka<�na<�sa<*ya<�~a<_�a<��a<ˍa<�a<:�a<&�a<�a<2�a<��a<u�a<>�a<P�a<��a<d�a<��a<��a<ۇa<d�a<V�a< �a<��a<A�a<5�a<%�a<��a<�a<mza<'ta<�ma<�fa<j`a<eZa<�Ua<�Qa<�Oa<fOa<�Pa<pSa<ZWa<P\a<�aa<>ga<�la<�qa<Xua<Sxa<za<�za<�za<�ya<�wa<va<ta<�ra<Yqa<�pa<�pa<qa<�qa<sa<Vta<�ua<6va<Hva<Wua<�sa<�pa<gla<bga<�aa<�[a<jUa<�Oa<�Ja<�Fa<EDa<TCa<%Da<�Fa<`Ja<cOa<Ua<@[a<�  �  �ba<Lha<ma<qa<�sa<�ua<zva<va<Wua< ta<�ra<Aqa<Fpa<�oa<�oa<�pa<�qa<�sa<�ua<�wa<�ya<C{a<,|a<�{a<�za<xa<�ta<kpa<hka<<fa<�`a<<\a<EXa<�Ua<�Ta<�Ta<�Va<�Ya<�^a<ada<�ja<rqa<�wa<�}a<قa<0�a<!�a<5�a<�a<�a<��a<ȋa<�a<�a<��a<��a<B�a<��a<_�a<��a<�a<E�a<6�a<��a<)�a<|�a<�a<�a<N�a<s�a<8�a<�a<Aza<�ua<�qa<oa<�ma<Vna<6pa<bsa<xa<]}a<Z�a<?�a<�a<�a<�a<`�a<G�a<b�a<0�a<h�a<	�a<��a<�a<y�a<��a<$�a<d�a<P�a<��a<g�a<�a<��a<͞a<��a<�a<��a<3�a<y�a<�a<��a<݇a<��a<O|a<twa<�sa<jqa<vpa<"qa<+sa<�va<E{a<��a<�a<�a<��a<��a<��a<(�a<��a<
�a<C�a<�a<]�a<��a<��a<D�a<4�a<ʓa<�a<Дa<�a<��a<�a<d�a<�a<^�a<H�a<d�a<1�a<"�a<�a<O�a<\�a<Jza<�ta<�oa<�la<tja<�ia<�ja<ma<�pa<cua<�za<D�a<x�a<g�a<#�a<>�a<�a<��a<N�a<��a<#�a<�a<��a<P�a<��a<,�a<x�a<x�a<Ӆa<φa<̇a<��a<Q�a<f�a<��a<҆a<�a<�a<){a<7ua<�na<mha<�aa<N\a<pWa<$Ta<%Ra<�Qa<�Ra<LUa<7Ya<�]a<<ca<ha<�ma< ra<�ua<Lxa<�ya<?za<�ya<Gxa<pva<�ta<tra<�pa<?oa<wna<[na<�na<�oa<kqa<�ra<0ta<ua<�ua<�ta<Tsa<�pa<�la<Pha<�ba<�\a<Wa<\Qa<�La<�Ha<�Fa<�Ea<zFa<�Ha<CLa<Qa<�Va<�\a<�  �  ada<oia<�ma<[qa<�sa<�ta<2ua<�ta<Tsa<�qa<�oa<"na<�la<Nla<�la<$ma<�na<�pa<sa<�ua<xa<�ya< {a<7{a<zza<�xa<�ua<�qa<:ma<\ha<�ca<H_a<�[a<.Ya<�Wa<KXa<'Za<u]a<�aa<Ega<7ma<msa<jya<�~a<��a<Q�a<��a<E�a<��a<��a<s�a<%�a<�a<ǆa<$�a<?�a<��a<*�a<5�a<��a<X�a<
�a<��a<4�a<&�a<
�a<�a<��a<8�a<�a<+�a<�a<}a<�xa<ua<�ra<iqa<�qa<�sa<�va<{a<�a<��a<�a<Q�a<�a<��a<W�a<ǜa<E�a<˜a<��a<��a<��a<Еa<A�a<�a<�a< �a<�a<u�a<q�a<��a<��a<R�a<4�a<\�a<f�a<t�a<D�a<�a<A�a<�a<n�a<La<�za<:wa<�ta<�sa<�ta<�va<za<G~a<:�a<��a<ݍa<��a<Ŗa<��a<��a<�a<a<Лa<�a<�a<��a<��a<�a<̐a<��a<��a<��a<��a<ǔa<��a<��a<��a<1�a<��a<M�a<��a<��a<\�a<!�a<|�a<�|a<�wa<fsa<�oa<�ma<Kma<3na<�pa<ta<Hxa<&}a<?�a<�a<_�a<�a<_�a<��a<Œa<�a<\�a<�a<I�a<��a<)�a<"�a<قa<+�a<��a<��a<Ƀa<�a<s�a<��a<�a<��a<`�a<(�a<��a<|a<�va<�pa<�ja<�da<�_a<�Za<�Wa<�Ua</Ua<KVa<�Xa<R\a<�`a<hea<Vja<�na<�ra<.va<Dxa<*ya<#ya<(xa<zva<ta<�qa<Uoa<[ma<�ka<6ka<�ja<�ka<�la<vna<Epa<ra<�sa<=ta<2ta<sa<�pa<�ma<^ia<nda< _a<~Ya<XTa<�Oa<PLa<�Ia<&Ia<�Ia<!La<�Oa<Ta<CYa<�^a<�  �  �fa<%ka<�na<�qa<zsa<ta<�sa<�ra<�pa<Zna<&la<Cja<�ha<�ga<�ga<�ha<�ja<�la<�oa<tra<[ua<�wa<�ya<�za<]za< ya<�va<�sa<�oa<Uka<-ga<ca<�_a<�]a<�\a<�\a<�^a<�aa<�ea<�ja<qpa<va<�{a<U�a<w�a<u�a<s�a<.�a<�a<*�a<�a<υa<�a<ڂa<ҁa<��a<c�a<уa<@�a<��a<��a<�a<�a<d�a<��a<��a<�a<q�a<��a<�a<��a<6�a<��a<�|a<Rya<wa<va<kva<#xa<{a<�~a<��a<��a<��a<M�a<0�a<K�a<E�a<:�a<��a<ۚa<�a<��a<M�a<��a<7�a<��a<E�a<y�a<��a<��a<��a<H�a<a<'�a<��a<k�a<+�a<��a<E�a<��a<��a<��a<Їa< �a<�~a<�{a<mya<�xa<*ya<	{a<~a< �a<��a<[�a<2�a<[�a<חa<R�a<��a<�a< �a<��a<M�a<��a<�a<��a<a<J�a<�a<�a<{�a< �a<J�a<��a<ؕa<��a<��a<�a</�a<>�a<2�a<@�a<��a<u�a<��a<�{a<�wa<rta<�ra<�qa<�ra<�ta<�wa<�{a<`�a<�a<F�a<Ռa<Ïa<��a<>�a<��a<$�a<�a<�a<�a<�a<<�a<�a<J~a<�}a<�}a<�~a<�a<��a<w�a<5�a<5�a<��a<�a<8�a<k�a<t}a<�xa<vsa<�ma<vha<Xca<4_a<\a<@Za<�Ya<�Za<�\a<`a<6da<oha<�la<�pa<=ta<�va<2xa<�xa<�wa<9va<�sa<qa<Bna<}ka<Ria<dga<�fa<rfa<Yga<�ha<�ja<ma<>oa<gqa<�ra<Bsa<�ra<Aqa<�na<ka<�fa<�aa<�\a<Xa<�Sa<�Pa<�Na<�Ma<�Na<�Pa<�Sa<�Wa<�\a<�aa<�  �  ?ia<"ma<pa<ra<sa<sa<�qa<�oa<kma<�ja<�ga<Zea<�ca<�ba<�ba<�ca<kea<ha<gka<�na<Wra<tua<xa<�ya<2za<�ya<xa<�ua<era<�na< ka<�ga<�da<�ba<�aa<Bba<�ca<�fa<�ja<oa<ta<ya<�}a<�a<S�a<��a<ƈa<�a<�a<J�a<4�a<�a<�a<�}a<�|a<�|a<0}a<�~a<$�a<U�a<�a<��a<.�a<R�a<��a<�a<&�a<=�a<L�a<]�a<��a<ψa<Ȅa<Z�a<E~a<K|a<`{a<�{a<C}a<�a<��a<��a<�a<g�a<q�a<��a<�a<0�a<U�a<p�a<��a<�a<�a<-�a<J�a<�a<��a< �a<_�a<��a<��a<h�a<��a<��a<u�a<՚a<J�a<��a<�a<K�a<��a<�a<�a<��a<N�a<��a<��a<�~a<�}a<z~a<�a<�a<e�a<p�a<��a<��a<Y�a<��a<��a<`�a<��a<��a<�a<1�a<�a<ʍa<ϊa<��a<8�a<��a<�a<L�a<^�a<�a<��a<Ғa<K�a<5�a<#�a<�a<Ȗa<��a<W�a<J�a<�a<U�a<�a<s|a<�ya<�wa<Bwa<�wa<�ya<�|a<�a<�a<�a<��a<��a<��a<��a<��a<j�a<4�a<&�a<��a<�a<h�a<+}a<�za<"ya<fxa<�xa<�ya<k{a<�}a<�a<G�a<#�a<6�a<B�a<I�a<7�a<%a< {a<qva<�qa<�la<#ha<'da<Paa<�_a<(_a<�_a<�aa<�da<ha<�ka<�oa<sa<�ua<lwa<xa<�wa<Ova<�sa<�pa<�ma<#ja<�fa<"da<Zba<Vaa<Zaa</ba<�ca<nfa<Eia<la<�na<�pa< ra<\ra<�qa<�oa<�la</ia<�da<�`a<X\a<�Xa<�Ua<�Sa<!Sa<�Sa<�Ua<�Xa<6\a<v`a<�da<�  �  �ka<oa<:qa<�ra<�ra<�qa<�oa<ma<ja<tfa<7ca<k`a<1^a< ]a<�\a<^a<`a<@ca<�fa<�ja<#oa<�ra<&va<xa<"za<Uza<sya<�wa<;ua<xra<(oa<dla<�ia<;ha<�ga<�ga<�ia<la<�oa<�sa<xa<p|a<G�a<ƃa<@�a<�a< �a<Y�a<��a<K�a<��a<q}a<�za<�xa<Ewa<�va<rwa<Gya<�{a<�a<t�a<��a<+�a<�a<�a<)�a<h�a<�a<��a<��a<�a<��a<#�a<I�a<��a<�a<�a<o�a<Ђa<-�a<]�a<ʋa<Ϗa<W�a<��a<�a<��a<9�a<R�a<��a<�a<�a<<�a<��a<��a<��a<�a<5�a<��a<�a<��a<��a<5�a<,�a<��a<��a<��a<J�a<��a<f�a<��a<��a<d�a<��a<�a<��a<��a<d�a<��a<'�a<��a<
�a<�a<��a<F�a<[�a<I�a<&�a<F�a<�a<��a<t�a<:�a<ِa<Όa< �a<ޅa<*�a<��a<Ӏa<��a<�a<��a<y�a<��a<��a<��a<S�a< �a<�a<q�a<וa<k�a< �a<��a<|�a<�a<��a<
a<�}a<�|a<�}a<a<��a<��a<�a<C�a<��a<G�a<��a< �a<�a<ێa<�a<(�a<�a<�a<�{a<xa<Cua<nsa<�ra<sa<^ta<�va<0ya<b|a<Ea<��a<��a<~�a<��a<�a<��a<q}a<�ya<]ua<�pa<ma<lia<�fa<9ea<�da<tea<ga<�ia<Sla<�oa<�ra<@ua<wa<!xa<)xa<�va<�ta<Hqa<�ma<�ia<�ea<ba<�^a<�\a<�[a<�[a<�\a<�^a<�aa<�da<�ha<�ka<�na<�pa<�qa<ra<�pa<�na<�ka<|ha<�da<�`a<�]a<[a<�Ya<�Xa<zYa<�Za<�]a<�`a<�da<�ha<�  �  �na<qa<�ra<�ra<<ra<�pa<�ma<cja<xfa<\ba<�^a<R[a<�Xa<uWa<>Wa<kXa<�Za<4^a<;ba<�fa<�ka<Cpa<\ta<qwa<�ya<�za<�za<�ya</xa<�ua<�sa<qa<�na<�ma<Bma<�ma<oa<Oqa<eta<xa<�{a<�a<܂a<��a<3�a<؇a<b�a<�a<��a<J�a<�|a<4ya<va<jsa<�qa<%qa<�qa<�sa<�va<�za<'a<)�a<�a<��a<z�a<]�a<5�a<�a<��a<(�a<��a<k�a<��a<��a<̈a<o�a<ˆa<�a<F�a<D�a<�a<=�a<c�a<S�a<��a<��a<;�a<ؚa<X�a<�a<~�a<��a<E�a<�a<��a<`�a<p~a<�}a<~a<�a<p�a<��a<�a<~�a<��a<��a<��a<��a<��a<��a<r�a<L�a<��a<��a<��a<��a<^�a<��a<[�a<a<�a<�a<��a<��a<��a<)�a<O�a<p�a<~�a<��a<o�a<x�a<��a<<�a<��a<r�a<Āa<�}a<�{a<2{a<�{a<�}a<�a<�a<��a<(�a<�a<��a<�a<�a<�a<K�a<��a<�a<�a<ٌa<��a<��a<|�a<.�a<��a<-�a<b�a<v�a<�a<Ƌa<Z�a<��a<	�a<��a<�a<.�a<c�a<��a<'�a<V�a<Z{a<�va<�ra<�oa<�ma<�la<�ma<oa<�qa<�ta<�xa<!|a<ra<�a<��a<W�a<��a<g�a<�a<�|a<ya<pua<�qa<�na<sla<�ja<�ja<�ja<-la<Ana<�pa<Esa<�ua<�wa<�xa<�xa<�wa<�ua<�ra<�na<ija<�ea<aa<]a<Ya<)Wa<�Ua<Va<IWa<�Ya<]a<�`a<�da<�ha<�la<koa<Oqa<+ra<�qa<�pa<tna<�ka<�ha<�ea<�ba<o`a<_a<�^a<_a<d`a<�ba<�ea<�ha<�ka<�  �  ?qa<�ra<�sa<:sa<�qa<Toa<�ka<�ga<ca<�^a<Za<cVa<�Sa<"Ra<�Qa<$Sa<�Ua<IYa<�]a<2ca<{ha<�ma<xra<vva<jya<U{a<|a<�{a<�za<!ya<Mwa<sua<�sa<�ra<`ra<�ra<'ta<}va<	ya</|a<Ta<��a<�a<��a<�a<�a<��a<^�a<U�a<m}a<Eya<Fua<eqa<yna<�la<�ka<ula<�na<�qa<�ua<({a<��a<�a<l�a<׏a<��a<-�a<��a<�a<K�a<�a<֓a<��a<��a<�a<u�a<�a<D�a<^�a<Q�a<��a<�a<��a<+�a<��a<Λa<ܛa<��a<r�a<�a<&�a<g�a<��a<�a<�~a<d{a<.ya<>xa<�xa<�za<�}a<r�a<E�a<�a<�a<��a<Q�a<(�a<�a<��a<�a<śa<��a<5�a<��a<g�a<��a<�a<��a<юa<�a<ґa<�a<T�a<��a<��a<ݛa<t�a<֛a<�a<A�a<u�a<��a<މa<��a<�a<�{a<�xa<�va<�ua<�va<�xa<�{a<�a<H�a<�a<��a<��a<��a<8�a<o�a<u�a<c�a<ӕa<?�a<��a<��a<��a<��a<M�a<�a<5�a<��a<�a<4�a<F�a<V�a<͒a<s�a<]�a<�a<~�a<�a<��a<K�a<�|a<kwa<*ra<�ma<�ja<mha<�ga<Sha<+ja<ma<�pa<�ta<2ya<;}a<e�a<�a<N�a<��a<ăa<�a<�a<�|a<rya<[va<�sa<yqa<6pa<�oa<pa<:qa<�ra<�ta<�va<lxa<gya<�ya<Zya<�wa<�ta<�pa<�la<Mga<
ba<�\a<(Xa<�Ta<�Qa<�Pa<�Pa</Ra<�Ta<zXa<]a<�aa<Wfa<�ja<&na<�pa<dra<�ra<1ra<�pa<�na<@la<�ia<nga<�ea<$da<�ca<!da<�ea<pga<�ia<Xla<�na<�  �  Usa<@ta<Uta<jsa<cqa<;na<&ja<rea<C`a<[a<]Va<]Ra<HOa<�Ma<AMa<�Na<\Qa<eUa<IZa<�_a<�ea<�ka<�pa<�ua<'ya<�{a<}a<p}a<"}a<|a<�za<)ya<�wa<wa<�va<�wa<�xa<�za<�|a<�a<`�a<�a<�a<E�a<��a<�a<�a<�a<Oa<�za<8va<�qa<�ma<Jja<ha<.ga<�ga<�ia<zma<-ra<�wa<r}a<��a<X�a<�a<�a<'�a<�a<#�a<#�a<h�a<ؖa<�a<i�a<�a<Ґa<��a<Аa<��a<<�a<E�a<e�a<��a<s�a<��a<ܜa<�a<y�a<��a<��a<�a<��a<X�a<<a<�za<wa<�ta<�sa<ta<va<lya<�}a<��a<(�a<��a<��a<%�a<��a<
�a<C�a<~�a<ʝa<_�a<[�a<B�a<A�a<��a<��a<C�a<P�a<B�a<��a<��a<��a<p�a<՜a<z�a<C�a<�a<��a<'�a<��a<��a<�a<r�a<C|a<�wa<>ta<�qa<3qa<�qa<7ta<�wa<�{a<��a<<�a<a�a<	�a<��a<��a<��a<n�a<�a<�a<'�a<�a<��a<��a<�a<Ռa<��a<��a<��a<�a<��a<R�a<�a<��a<ɔa<ߓa<��a<ގa<��a<��a<�a<�ya<�sa<ena<�ia<fa<�ca<ca<�ca<�ea<Bia<?ma<�qa<�va<({a<a<4�a<I�a<�a<��a<�a<�a<�a<�|a</za<�wa<�ua<�ta<6ta<Pta<%ua<zva<�wa<tya<�za<({a<�za<�ya<kwa<�sa<}oa<Pja<�da<�^a<7Ya<STa<6Pa<XMa<�Ka<La<�Ma<�Pa<�Ta<wYa<�^a<�ca<�ha<�la<Opa<�ra<�sa<�sa<�ra<tqa<doa<Fma<Gka<�ia<�ha<vha<�ha<�ia<Nka<Zma<�oa<�qa<�  �  �ta<�ua<�ta<�sa<qa<ima<�ha<�ca<0^a<�Xa<[Sa<�Na<�Ka<Ja<�Ia<'Ka<�Ma<	Ra<QWa<e]a<�ca<�ia<�oa<�ta<�xa<�{a<�}a<�~a<�~a<!~a<}a<|a<�za<wza<Hza<�za<�{a<�}a<�a<f�a<��a<҆a<g�a<\�a<�a<�a<k�a<:�a<�}a<ya<ta<�na<|ja<�fa<�da<�ca<]da<�fa<�ia<�na<�ta<,{a<��a<҇a<��a<,�a<�a<��a<-�a<��a<�a<�a<ܗa<t�a<�a<M�a<�a<(�a<�a<a�a<@�a<��a<��a<�a<�a<��a<z�a<S�a<ǖa<��a<H�a<��a<�a<P|a<wwa<�sa<0qa<pa<�pa<�ra<�ua<�za<�a<�a<֋a<v�a<K�a<0�a<%�a<Ԟa<��a<6�a<J�a<��a<*�a<d�a<�a<�a<��a<��a<��a<Әa<}�a<�a<l�a<D�a<��a<�a<0�a<J�a<U�a<��a<Ҋa<�a<�~a<@ya<bta<�pa<�na<�ma<�na<�pa<Pta<ya<y~a<8�a<��a<�a<4�a<��a<��a<:�a<r�a<��a<@�a<n�a<��a<��a<H�a<5�a<Ϗa<�a<ɐa<�a<m�a<��a<��a<�a<ߕa<Y�a<��a<9�a<��a<�a<�}a<�wa<qa<Aka<4fa<�ba<V`a<�_a<\`a<qba<fa<qja<�oa<�ta<�ya<(~a<�a<<�a<��a<�a<D�a<̓a<Ɂa<�a<:}a<�za<Pya<xa<�wa<�wa<Ixa<vya<�za<�{a<I|a<�|a<�{a<�ya<Ewa<0sa<na<�ha<�ba<]\a<KVa<Qa<�La<�Ia<uHa<�Ha<JJa<OMa<�Qa<�Va<�\a<ba<~ga<!la<�oa<�ra</ta<�ta<[ta<^sa<�qa<-pa<ina<�la<la<�ka<la<ma<ona<Ipa<�qa<�sa<�  �  �ua<va<\ua<�sa<�pa<�la< ha<qba<�\a<�Va<�Qa<Ma<�Ia<�Ga<oGa<�Ha<�Ka<#Pa<�Ua<�[a<Oba<�ha<�na<Lta<�xa<|a<A~a<�a<�a<�a<�~a<�}a<�|a<�|a<t|a<}a<~a<�a<��a<�a<*�a<�a<Y�a<�a<g�a<�a<-�a<��a<�|a<�wa<cra<Uma<�ha<�da<}ba<caa<ba<]da<ha<ma<%sa<�ya<W�a<ǆa<�a<�a<�a<�a<��a<g�a<\�a<��a<h�a<�a< �a<e�a< �a<]�a<2�a<[�a<ՙa<��a<#�a<?�a<��a<-�a<Ŝa<,�a<h�a<đa<)�a<Z�a<W�a<�za<�ua<�qa<�na<�ma<Rna<�pa<ta<�xa<�~a<{�a<��a<x�a<Õa<��a<>�a<9�a<B�a<A�a<��a<D�a<��a<!�a<��a<�a<Øa<ݘa<��a<��a<�a<~�a<Ȟa<W�a<W�a<I�a<T�a<�a<Ӕa<��a<��a<l�a<I}a<�wa<�ra<�na<8la<_ka<Fla<�na<jra<\wa<�|a<Âa<��a<�a<Ȓa<��a<7�a<��a<+�a<��a<��a<��a<<�a<��a<]�a<a�a<	�a<(�a<Ԓa<��a<��a<�a<�a<
�a<g�a<��a<��a<��a<�a<�a<�|a<�ua<{oa<`ia<Uda<{`a<�]a<7]a<0^a<�`a<&da<�ha<�ma<osa<�xa<u}a<:�a<-�a<߅a<��a<'�a<�a<?�a<�a<�~a< }a<h{a<Pza<�ya<�ya<Cza<
{a<|a<}a<�}a<L}a<>|a<Eza<wa<�ra<�ma<�ga<Baa<�Za<�Ta<Oa<�Ja<�Ga<Fa<QFa<=Ha<sKa<�Oa<BUa<�Za<�`a<�fa<�ka<�oa<�ra<�ta<ua<gua<�ta<Lsa<�qa<%pa<oa<(na<�ma<*na<oa<8pa<�qa<sa<ua<�  �  �ta<�ta<ta<�ra<�pa<�ma<�ia<�ea<yaa<]a<Ya<�Ua<LSa<�Qa<�Qa<�Ra<0Ua<�Xa<�\a<�aa<�fa<�ka<npa<�ta</xa<�za<�|a<�}a<O~a<:~a<�}a<�}a<}a<�|a<�|a<�}a<S~a<�a<��a<P�a<�a<i�a<��a<'�a<��a<��a<لa<�a<�~a<4{a<wa<ysa<�oa<Rma<�ka<ka<�ka<�ma<|pa<ita<9ya<"~a<��a<��a</�a<O�a<��a<ɖa<��a<�a<�a<��a<$�a<l�a<Җa<��a<	�a<7�a<Ӗa<�a<%�a<J�a<V�a<!�a<��a<6�a<ךa<�a<;�a<��a<��a<�a<S�a<0�a<;}a<Aza<bxa<�wa<�wa<�ya<:|a<�a<6�a<ֈa<��a<ܑa<�a<1�a<��a<N�a<.�a<=�a<��a<Мa<ޛa<��a<�a<�a<ߘa<��a<��a<J�a<H�a<�a<ޜa<c�a<G�a<b�a<��a<<�a<��a<֐a<p�a<��a<؂a<o~a<�za<�wa<�ua<2ua<�ua<wa<@za<~a<�a<��a<�a<�a<ǒa<y�a<g�a<��a<�a<��a<חa<��a<��a<K�a<�a<G�a<�a<�a<��a<-�a<��a<q�a<єa<ٔa<H�a<��a<u�a<Z�a<[�a<��a<�a<|za<�ua<�pa<�la<�ia<�ga<�fa<�ga<ia<�ka<8oa<�ra<wa<�za<%~a<�a<�a<?�a<܄a<c�a<`�a< �a<p�a<�~a<L}a<�{a<�za<8za<za<�za<�za<l{a<�{a<�{a<�{a<�za<�xa<vva<9sa<oa<{ja<�ea<Y`a<�[a<_Wa<�Sa<�Qa<~Pa<�Pa<�Qa<,Ta<�Wa<�[a<�_a<rda<�ha<fla<zoa<�qa<Msa<ta<ta<dsa<�ra<�qa<npa<�oa<�na<�na<�na<�oa<�pa<�qa<�ra<�sa<�  �  [ta<vta<�sa<�ra<�pa<�ma<ja<�ea<�aa<q]a<�Ya<`Va<�Sa<�Ra<yRa<�Sa<�Ua<;Ya<Y]a<�aa<�fa<�ka<�pa<�ta<Gxa<�za<�|a<�}a<'~a<~a<z}a<�|a<`|a<>|a<J|a<�|a<�}a<>a<܀a<ςa<��a<W�a<b�a<�a<��a<؆a<̈́a<D�a<�~a<Q{a<xwa<�sa<�pa<na<Ola<�ka<^la<7na<-qa<ua<�ya<�~a<��a<��a<b�a<9�a<��a<Ȗa<:�a<�a<�a<y�a<��a<��a< �a<��a<i�a<��a<P�a<=�a<��a<ٙa<�a<��a<I�a<��a<�a<�a<!�a<��a<��a<B�a<a<��a<�}a<�za<ya</xa<�xa<4za<�|a<n�a<��a<�a<��a<�a<��a<8�a<a<0�a<��a<�a<��a<t�a<U�a<�a<.�a<j�a<@�a<?�a<ܘa<��a<��a<��a<ʜa<=�a<�a<?�a<Ța<D�a<��a<�a<��a<�a<4�a<�~a<>{a<Rxa<�va<�ua<vva<+xa<�za<�~a<�a<�a<+�a<E�a<��a<��a<�a<}�a<٘a<��a<��a<K�a<�a<��a<��a<��a<p�a<g�a<בa<u�a<_�a<&�a<��a<��a<�a<��a<��a<O�a<��a<�a<�a<�za<�ua<Dqa<^ma<Qja<fha<�ga<.ha<�ia<Vla<�oa<?sa<.wa<�za<X~a<��a<5�a<>�a<��a<5�a<M�a<��a<�a<~a<z|a<{a<5za<�ya<�ya<�ya<Oza<�za<�{a<�{a<�{a<�za<�xa<�va<sa<8oa<�ja<�ea<�`a<.\a<Xa<�Ta<ZRa<#Qa<6Qa<wRa<�Ta<Xa<�[a<7`a<�da<�ha<nla<�oa<�qa</sa<�sa<�sa<Rsa<#ra< qa<�oa<�na<-na<na<4na<�na<�oa<)qa<^ra<�sa<�  �  bsa<�sa<�sa<�ra<�pa<�ma<�ja<�fa<�ba<�^a<�Za<�Wa<]Ua<0Ta<Ta<Ua<JWa<�Za<�^a<7ca<ha<�la<Yqa< ua<]xa<�za<I|a<!}a<+}a<�|a<V|a<�{a<{a<�za<�za<L{a<q|a<�}a<�a<��a<s�a<F�a<��a<��a<u�a<ņa<�a<ʂa<�a<B|a<�xa<ua<�qa<toa<�ma<]ma<na<�oa<�ra<qva<�za<�a<��a<~�a<��a<z�a<��a<��a<ؗa<9�a< �a<E�a<��a<��a<��a<!�a<ʓa<�a<�a<ڕa<P�a<��a<�a<��a<��a<��a<��a< �a<j�a<r�a<r�a<N�a<	�a<ւa<Za<b|a<�za<�ya<6za<�{a<]~a<Ɓa<Ʌa<N�a<��a<֒a<d�a<[�a<��a<�a<��a<)�a<x�a<I�a<.�a<Ƙa<��a<�a<��a<��a<g�a<G�a<��a<��a<��a<D�a<��a<��a<��a<a�a<S�a<ˑa<w�a<�a<u�a<D�a<�|a<�ya<xa<~wa<�wa<�ya<l|a<�a<ăa<��a<�a<��a<��a<��a<U�a<(�a<D�a<��a<��a<(�a<��a</�a<�a<%�a<Ϗa<�a<n�a<:�a<:�a<�a<��a<�a<��a<h�a<��a<��a<	�a<��a<�a<|a<wa<�ra<�na<�ka<ja<Pia<�ia<Aka<�ma<�pa<�ta<!xa<�{a<�~a<>�a</�a<�a<3�a<��a<A�a<��a<�~a<�|a<{a<�ya<�xa<xa<(xa<]xa< ya<�ya<jza<�za<�za<8za<�xa<�va<gsa<�oa<jka<�fa<ba<h]a<}Ya<Va<�Sa<�Ra<�Ra<�Sa<OVa<lYa<(]a<kaa<}ea<~ia<�la<�oa<�qa<�ra<bsa<�ra<3ra<�pa<�oa<tna<oma<�la<lla<�la<~ma<�na<�oa<6qa<�ra<�  �  Tra<sa<3sa<jra<qa<�na<�ka<8ha<eda<�`a<(]a<CZa<Xa<�Va<�Va<�Wa<�Ya<]a<�`a<ea<�ia<na<ra<�ua<�xa<yza<�{a<1|a<|a<c{a<zza<iya<�xa<)xa<"xa<�xa<�ya<m{a<B}a<�a<ځa<�a<��a<φa<�a<��a<��a<i�a<΀a<�}a<Nza<*wa<3ta<�qa<�pa< pa<�pa<kra<0ua<�xa<�|a<m�a<)�a<��a<��a<&�a<��a<=�a<8�a<4�a<��a<��a<x�a<&�a<9�a<d�a<H�a<u�a<8�a<y�a<�a<Öa<m�a<ۙa<��a<�a<w�a<-�a<&�a<�a<��a<Ōa<Ĉa<
�a<��a<
a<7}a<v|a<�|a<]~a<׀a<�a<ԇa<Ӌa<��a<��a<!�a<Ǚa<v�a<��a<��a<�a<�a<��a<��a<b�a<?�a<I�a<�a<�a<�a<�a<Q�a<ۘa<4�a<5�a<��a<��a<m�a<��a<�a<��a<Ύa<��a<o�a<|�a<#a<{|a<�za< za<�za<G|a<�~a<�a<��a<w�a<S�a<��a<��a<˕a<�a<��a<T�a<w�a<��a<L�a<k�a<ʏa<x�a<��a<N�a<F�a<�a<ڎa<"�a<Z�a<Y�a<ݒa<�a<�a<h�a<�a<��a<ǆa<c�a<�}a<3ya<�ta<Xqa<�na<�la<�ka<bla<�ma< pa<�ra<"va<�ya<�|a<�a<�a< �a<��a<��a<~�a<��a<�~a<�|a<�za<�xa<wa<va<wua<vua<�ua<�va<�wa<�xa<�ya<�ya<�ya<�xa<�va<#ta<�pa<�la<Aha<�ca<�_a<�[a<�Xa<�Va<jUa<uUa<�Va<�Xa<�[a<3_a<�ba<�fa<eja<�ma<pa<�qa<�ra<�ra<�qa<�pa<Poa<�ma<la<�ja<ja<�ia<ja<�ja<#la<�ma<oa<qa<�  �  �pa<�qa<�ra<Ura<Hqa<�oa<�la<ja<�fa<Aca<�_a<']a<G[a<;Za<;Za<-[a<#]a<�_a<�ca<�ga<�ka<�oa<*sa<iva<�xa<Vza<{a<�za<aza<,ya<xa<�va<�ua<ua<�ta<xua<kva<^xa<\za<�|a<�a< �a<�a<��a<Ɔa<��a<�a<X�a<Q�a<�a<�|a<�ya<�va<ua<�sa<ksa<ta<�ua<:xa<�{a<�a<ƃa<(�a<9�a<��a<��a<��a<��a<'�a<��a<Ӕa<k�a<�a<=�a</�a<#�a<��a<5�a<�a<��a<!�a<H�a<.�a<�a<E�a<:�a<J�a<?�a<��a<%�a<a�a<Ўa<:�a<χa<��a<+�a<��a<�a<A�a<��a<ǃa<ʆa<n�a<��a<�a<�a<�a<�a<d�a<�a<v�a<��a<�a<2�a<K�a<{�a<&�a<��a<Őa<ΐa<Ña<��a<��a<h�a<�a<��a<j�a<�a<X�a<��a<ږa<��a<��a<��a<�a<E�a<�a<�a<#~a<�}a<
~a<sa<��a<��a<�a<��a<�a<Бa<d�a<�a<�a<�a<�a<Ĕa<ɒa<Ԑa<��a<݌a<V�a<K�a<��a<��a<��a<�a<��a<�a<h�a<a�a<͑a<��a<b�a<��a<��a<J�a<Z�a<�a<�{a<�wa<]ta<�qa<pa<aoa<�oa<�pa<�ra<�ua<{xa<�{a<i~a<��a<a�a<�a<m�a<��a<�a<a<�|a<5za<�wa<�ua<�sa<�ra<7ra<Jra<	sa<�sa<iua<�va<�wa<�xa<�xa<]xa<�va<�ta<�qa<Xna<Kja<>fa<_ba<�^a<�[a<�Ya<�Xa<�Xa<�Ya<�[a<o^a<�aa<ea<�ha<�ka<dna<]pa<�qa<ra<Zqa<gpa<�na<�la<�ja<)ia<�ga<�fa<�fa<�fa<�ga<;ia<
ka<ma<�na<�  �  �na<�pa<�qa<ra<�qa<qpa<mna<�ka<ia<	fa<Eca<�`a<_a<,^a<*^a<_a<�`a<�ca<�fa<Oja<�ma<rqa<�ta<,wa<�xa<�ya<za<�ya<Txa<�va<ua<rsa<�qa<<qa<�pa<fqa<�ra<�ta<�va<�ya<�|a<�a<��a<��a<�a<��a<��a<��a<΃a<��a<Qa<�|a<�za<�xa<�wa<mwa<xa<�ya<�{a<2a<��a<��a<1�a<��a<�a<!�a<��a<F�a<�a<E�a<��a<��a<�a<�a<X�a<s�a<�a<:�a<L�a<��a<�a<[�a<��a<�a<��a<&�a<��a<t�a<o�a<��a<�a<�a<�a<݊a<F�a<�a<t�a<�a<9�a<i�a<��a<9�a<B�a<��a<��a<��a<��a<x�a<+�a<�a<J�a<ǘa<��a<h�a<3�a<�a<G�a<6�a<��a< �a<�a<_�a<{�a<��a<��a<��a<9�a<�a<	�a<S�a<Ǘa<f�a<y�a<=�a<΋a<��a<Ӆa<|�a<�a<��a<�a<4�a<c�a<އa<ߊa<�a<��a<P�a<'�a<1�a<q�a<�a<��a<��a<K�a<�a<t�a<$�a<��a<d�a<�a<O�a<�a<��a<z�a<O�a<0�a<ҏa<��a<��a<Y�a<�a<ڌa<Ɖa<N�a<��a<�~a<P{a<"xa<�ua<ta<csa<�sa<�ta<�va<�xa<A{a<�}a<�a<ށa<�a<,�a<��a<n�a<�a<�|a<za<4wa<Lta<�qa<pa<�na<<na<�na<Boa<�pa<}ra<ta<�ua<5wa<�wa<�wa<�va<jua<sa<�oa<�la<	ia<lea<gba<�_a<�]a<�\a<�\a<�]a<�_a<�aa<�da<�ga<�ja<Ema<ooa<�pa<Mqa<qa<.pa<�na<fla<ja<�ga<�ea<�ca<�ba<�ba<�ba< da<�ea<�ga<9ja<�la<�  �  �la<(oa<�pa<�qa<�qa<Fqa<pa<�ma<�ka<ia<�fa<�da<.ca<sba<Uba<aca<�da<Xga<ja<Lma<�pa<asa<va<�wa<,ya<wya<ya<�wa<va<1ta<�qa<�oa<+na<&ma<�la<$ma<�na<�pa<isa<cva<	za<t}a<��a<W�a<B�a<��a<��a<��a<��a<��a<�a<�a<4~a<�|a<�{a<�{a<:|a<�}a<�a<ӂa<υa<f�a<��a<��a<	�a<��a<��a<��a<�a<X�a<X�a<�a<j�a<e�a<c�a<V�a<��a<�a<.�a<�a<_�a<��a<�a<��a<A�a<�a<<�a<��a<�a<�a<�a<��a<��a<%�a<�a<މa<ňa<�a<{�a<��a<X�a<��a<[�a<Z�a<ٕa<D�a<�a<ߚa<�a<>�a<�a<��a<J�a<k�a<��a<M�a<A�a<�a<k�a<܈a<܉a<��a<�a<{�a<I�a<��a<×a<�a<ؙa<��a<��a<��a<��a<�a<ގa<�a<��a<��a<^�a<��a<@�a<5�a<�a<;�a<ݍa<��a<��a<��a<ڕa<y�a<�a<�a<�a<}�a<΍a<��a<�a<V�a<t�a<7�a<��a<4�a<�a< �a<�a<��a<ڋa<эa<w�a<3�a<g�a<|�a<�a<��a<��a<z�a<�a<�~a<�{a<�ya<Dxa<�wa<�wa<}xa<"za<�{a<~a<�a<Ła<�a<n�a<M�a<�a<B�a<�}a<�za<Swa<�sa<�pa<�ma<�ka<yja<ja<mja<fka<.ma<oa<�qa<�sa<|ua<�va<Mwa<6wa<va<hta<�qa<oa<�ka<�ha<fa<�ca<ba<�`a<aa<�aa<Hca<^ea<�ga<vja<�la<�na<[pa<)qa<2qa<>pa<�na<xla<ja<ga<Uda<�aa<�_a<�^a<H^a<�^a<�_a<�aa<]da<!ga<*ja<�  �  �ja<�ma<�oa<�qa<;ra<9ra<�qa<pa<*na<;la<Mja<kha<8ga<�fa<�fa<|ga<�ha<�ja<�ma<:pa<�ra<yua<jwa<�xa<<ya<ya<xa<<va<�sa<mqa<�na<_la<eja<�ha<�ha<�ha<Uja<�la<�oa<#sa<wa<�za<�~a<�a<��a<t�a<��a<��a<b�a<@�a<��a<M�a<��a<z�a<�a<�a<o�a<�a<Ƀa<V�a<D�a<�a<�a<t�a<+�a<P�a<��a<�a<��a<z�a<�a<0�a<0�a<Åa<�a<�a<��a<ׁa<�a<�a<Їa<Պa<H�a<z�a<z�a<�a<ǘa<��a<ڙa<5�a<�a<��a<Γa<��a<��a<ߍa<��a<R�a<��a<��a<�a<K�a<��a<ϕa<�a<יa<ޚa<6�a<Śa<��a<t�a<��a<��a<h�a<?�a<��a<8�a<Ǆa<>�a<��a<ǅa<�a<v�a<p�a<��a<��a<6�a<F�a<��a<�a<��a<}�a<��a<\�a<�a<��a<N�a<��a<��a<�a<\�a<;�a<��a<ʎa<͐a<ߒa<ʔa<�a<��a<��a<��a<�a<a�a<V�a<�a<��a<`�a<��a<Fa<�}a<�}a<�}a</a<X�a<��a<��a<W�a<�a<1�a<��a<0�a<�a<��a<Z�a<�a<�a<U�a<n�a<�a<�}a<u|a<�{a<�{a<k|a<�}a<Ea<Àa<\�a<��a<#�a<�a<#�a<|�a<a<�{a<(xa<tta<}pa<#ma<�ia<�ga<Vfa<�ea<3fa<�ga<�ia<�ka<�na<Rqa<�sa<�ua<�va<1wa<�va<�ua<�sa<rqa<�na<?la<�ia<�ga<1fa<Bea<>ea<�ea<
ga<�ha<�ja<�la<�na<�pa<Uqa<�qa<�pa<�oa<Yma<�ja<hga<da<�`a<D^a<�[a<�Za<Za<�Za<�[a<2^a<�`a<da<{ga<�  �  �ha<la<oa<*qa<�ra<0sa<�ra<ra<�pa<oa<oma<la<ka<lja<�ja<7ka<�la<una<�pa<�ra<;ua<=wa<�xa<�ya<iya<�xa<�va<�ta<ra<�na<�ka<�ha<�fa<$ea<�da<ea<rfa<�ha<la<pa<Qta<�xa<}a<��a<�a<I�a<"�a<ֈa<��a<W�a<L�a<?�a<��a<F�a<��a<҃a<��a<��a<��a<��a<A�a<��a<�a<ܒa<B�a<��a<o�a<w�a<T�a<�a<ʋa<e�a<8�a<	�a<�a</~a<�}a<�}a<#a<Q�a<<�a<�a<��a<��a<��a<ޕa<Q�a<a<��a<S�a<��a<:�a<��a<Ŕa<��a<��a<��a<e�a<��a<t�a<Βa<u�a<z�a<G�a<�a<�a<�a<��a<{�a<��a<�a<��a<B�a<��a<�a<ʄa<t�a<��a<N�a<��a<��a<"�a<-�a<��a<�a<Ǒa<��a<f�a<-�a<C�a<��a<��a<��a<ʖa<۔a<ǒa<�a<|�a<X�a<�a<�a<�a<9�a<ߑa<��a<0�a<��a<:�a<��a<��a<7�a<ؒa<ُa<q�a<c�a<��a<�a<�}a<r{a<�ya<�ya<za<p{a<�}a<��a<΃a<�a<Y�a<��a<�a<�a<��a<�a<��a<�a<��a<G�a<��a<��a<��a<z�a<�a<�a<>�a<�a<A�a<f�a<~�a<�a<:�a<��a<
�a<�a<�}a<?za<va<�qa<�ma<jia<:fa<�ca<Uba<�aa<bba<�ca<fa<ia<
la<coa<8ra<�ta<bva<Ewa<�wa<�va<�ua<�sa<�qa<Qoa<ma<pka<�ia<Uia<ia<�ia<�ja<la<�ma<coa<�pa<�qa<Xra<�qa<�pa<�na<�ka<�ha<ea<Xaa<�]a<}Za</Xa<�Va<.Va<�Va<Xa<gZa<�]a<Saa< ea<�  �  ga<�ja<Zna<�pa<�ra<�sa<ta<�sa<�ra<�qa<*pa<�na<0na<�ma< na<�na<�oa<[qa<[sa<eua<Dwa<�xa<�ya<	za<xya<Kxa< va<Qsa<%pa<�la<@ia<fa<�ca<�aa<-aa<�aa<ca<�ea<'ia<_ma<�qa<�va<i{a<�a<q�a<>�a<T�a<��a<+�a<#�a<��a<��a<чa<A�a<��a<�a<ˇa<݈a<��a<��a<Ɏa<��a<�a<U�a<E�a<6�a<o�a<��a<O�a<U�a<ȉa<�a<��a<5a<�|a<�za<za<lza<�{a<O~a<r�a<N�a<U�a<��a<��a<��a<�a<˙a<�a<�a<�a<5�a<�a<b�a<ەa<Δa<ޓa<��a<̓a<��a<��a<:�a<�a<y�a<��a<p�a<��a<śa<N�a<
�a<̔a<7�a<)�a<�a<F�a<�a<Ea<}}a<�|a<;}a<�~a<@�a<d�a<�a<�a<��a<{�a<��a<�a<]�a<&�a<��a<=�a<�a<P�a<��a<ړa<��a<��a<k�a<j�a<1�a< �a<��a<��a<9�a<�a<p�a<�a<ǖa<�a<�a<w�a<��a<5�a<�a<~a<�za<8xa<�va<va<�va<Uxa<�za<�}a<`�a<�a<��a<��a<a�a<��a<Ӑa<��a<"�a<Ύa<�a<Ɗa<��a<��a<�a<��a<�a<Ԃa<E�a<ԃa<Ʉa<��a<[�a<��a<=�a<��a<
�a<p�a<�|a<�xa<ta<Hoa<�ja<�fa<+ca<�`a<�^a<o^a<!_a<�`a<Aca<ofa<�ia<qma<�pa<�sa<va<Mwa<xa<�wa< wa<�ua<�sa<�qa<�oa<�na<,ma<�la<`la<�la<�ma<�na<Npa<�qa<�ra<sa<sa<ra<rpa<na<�ja<ga<�ba<�^a<�Za<�Wa<Ua<ISa<�Ra<7Sa<�Ta<�Wa<�Za<�^a<�ba<�  �  �ea<ja<�ma<�pa<�ra<Cta<�ta<�ta</ta<Esa<ora<Zqa<�pa<Upa<}pa<3qa<Pra<�sa<�ua<	wa<�xa<�ya<�za<fza<�ya<�wa<kua<ara<�na<ka<-ga<�ca<(aa<0_a<�^a<�^a<k`a<ca<�fa<,ka<1pa<<ua<.za<�~a<��a<<�a<��a<B�a<$�a<N�a<�a<��a<.�a<��a<��a<��a<N�a<��a<��a<�a<Аa<��a<+�a<V�a<ڕa<��a<y�a<G�a<��a<'�a<R�a<`�a<S�a<�|a<za<(xa<swa<�wa< ya<�{a<6a<,�a<Ƈa<+�a<z�a<R�a<c�a<�a<d�a<8�a<�a<��a<��a<��a<>�a<;�a<��a<:�a<f�a<3�a< �a<��a<a<��a<՜a<^�a<�a<
�a< �a<E�a<�a<�a<��a<@�a<�a<�a<�|a<�za<*za<�za<|a<�~a<.�a<(�a<��a<��a<��a<�a<��a<��a<��a<�a<L�a<b�a<�a<ȗa<?�a<(�a<C�a<�a<�a<��a<��a<��a<��a<��a<�a<7�a<f�a<�a<o�a<N�a<��a<'�a<��a< �a<�{a<Sxa<~ua<�sa<msa<�sa<�ua<uxa<�{a<�a<��a<s�a<�a<��a<��a<�a<�a<�a<��a<n�a<��a<��a<��a<��a<G�a<��a<��a<��a<1�a<Іa<8�a<��a<��a<҆a<L�a<�a<�a<|a<twa<�ra<�ma<�ha<Uda<�`a<�]a<A\a<�[a<_\a<L^a<aa<Mda<@ha<la<�oa<�ra<rua<nwa<\xa<�xa<
xa<wa<�ua<ta<[ra<�pa<�oa<)oa<�na<qoa<pa<-qa<ra<sa<�sa<ta<�sa<Ura<Epa<Hma<�ia<�ea<naa<�\a<�Xa<GUa<SRa<�Pa<Pa<�Pa<4Ra<Ua<�Xa<�\a<daa<�  �  �da<[ia<;ma<�pa<sa<�ta<pua<�ua<Wua<mta<�sa<�ra<0ra<�qa<'ra<�ra<�sa<ua<�va<4xa<�ya<�za<�za<�za<�ya<�wa<�ta<�qa<�ma<�ia<�ea<�ba<�_a<�]a<�\a<J]a<�^a<�aa<tea<�ia<�na<8ta<Wya<K~a<r�a<,�a<ʈa<��a<ʋa<R�a<C�a<݋a<_�a<�a<��a<=�a<�a<��a<e�a<�a<��a<��a<3�a<�a<?�a<��a<w�a<�a<�a<W�a<Y�a<�a<a<�{a<�xa<�va<�ua<(va<�wa<Yza<�}a<�a<��a<7�a<��a<ӓa<0�a<�a<��a<��a<�a<��a<��a<��a<{�a<��a< �a<ݗa<�a<��a<z�a<��a<�a<!�a<ϝa<�a<_�a<0�a<	�a<�a<T�a<�a<��a<��a<ρa<~a<'{a<Iya<�xa<ya<�za<`}a<�a<�a<Z�a<��a<��a<��a<��a<��a<�a<j�a<G�a<��a<6�a<��a<��a<��a<Ǖa<��a<��a<�a<ʖa<ݗa<ʘa<��a<��a<��a<��a<
�a<F�a<ېa<��a<3�a<u�a<�~a<�za<�va<ta<Wra<�qa<|ra<Bta<	wa<~za<e~a<��a<��a<h�a<b�a<�a<I�a<�a<��a<��a<��a<�a<�a<]�a<��a<�a<=�a<�a<�a<e�a<��a<l�a<��a<5�a<8�a<�a<�a<za<x{a<�va<�qa<^la<fga<�ba<$_a<Q\a<�Za<+Za<�Za<�\a<�_a<ca<�fa<ka<�na<ura<?ua<�wa<�xa<ya<�xa<xa<�va<2ua<�sa<Zra<Nqa<�pa<�pa<�pa<gqa<Wra<Csa<<ta<�ta<�ta<�sa<{ra<.pa<�la<<ia<�da<R`a<�[a<�Wa<�Sa<�Pa<Oa<jNa<Oa<�Pa<�Sa<YWa<�[a<=`a<�  �  �da<"ia<Ima<�pa<�ra<�ta<�ua<�ua<oua<�ta<*ta<asa<�ra<\ra<�ra<"sa<}ta<�ua<3wa<�xa<�ya<�za<9{a<�za<�ya<�wa<�ta<eqa<�ma<�ia<�ea<�aa<_a<!]a<D\a<�\a<K^a<�`a<�da<�ia<|na<ta<>ya<~a<��a<�a<��a<�a<��a<r�a<�a<O�a<	�a<Ӌa<z�a<Ջa<��a<t�a<8�a<Ɛa<k�a<��a<I�a<2�a<��a<��a<\�a<�a<�a<4�a<6�a<��a<�~a<�za<�wa<va<%ua<}ua<wa<�ya<<}a<��a<5�a<�a<��a<��a<8�a<��a<��a<��a<�a<��a<�a<*�a<1�a<n�a<~�a<��a<�a<7�a<4�a<M�a<O�a<E�a<��a<*�a<��a<�a<��a<�a<!�a<�a<\�a<��a<R�a<c}a<{za<�xa<�wa<_xa<za<�|a<a�a<��a<�a<��a<��a<��a<��a<��a<�a<��a<n�a<��a<��a<��a<G�a<A�a<J�a<2�a<�a<Ֆa<|�a<d�a<$�a<əa<%�a<�a<ɘa<�a<D�a<Ȑa<��a<�a<0�a<r~a<�ya<3va<osa<�qa<&qa<�qa<�sa<]va<za<�}a<w�a<��a<0�a<{�a<ʏa<;�a<)�a<��a<�a<ُa<W�a<��a<-�a<{�a<}�a<ڇa<l�a<ڇa<�a<k�a<��a<��a<c�a<�a<z�a<��a<�a<B{a<�va<{qa<�ka<ga<Gba<q^a<�[a<�Ya<Ya<TZa<-\a<_a<�ba<�fa<�ja<�na<Sra<Hua<awa<�xa<Sya<ya<(xa<�va<�ua<Mta<!sa<�qa<oqa<qa<uqa<"ra<�ra<�sa<`ta<�ta<�ta<ta<`ra<pa<ma<ia<�da<`a<G[a<Wa<Sa<9Pa<lNa<�Ma<\Na<"Pa<�Ra<�Va</[a< `a<�  �  �da<[ia<;ma<�pa<sa<�ta<pua<�ua<Wua<mta<�sa<�ra<0ra<�qa<'ra<�ra<�sa<ua<�va<4xa<�ya<�za<�za<�za<�ya<�wa<�ta<�qa<�ma<�ia<�ea<�ba<�_a<�]a<�\a<J]a<�^a<�aa<tea<�ia<�na<8ta<Wya<K~a<r�a<,�a<ʈa<��a<ʋa<R�a<C�a<݋a<_�a<�a<��a<=�a<�a<��a<e�a<�a<��a<��a<3�a<�a<?�a<��a<w�a<�a<�a<W�a<Y�a<�a<a<�{a<�xa<�va<�ua<(va<�wa<Yza<�}a<�a<��a<7�a<��a<ӓa<0�a<�a<��a<��a<�a<��a<��a<��a<{�a<��a< �a<ݗa<�a<��a<z�a<��a<�a<!�a<ϝa<�a<_�a<0�a<	�a<�a<T�a<�a<��a<��a<ρa<~a<'{a<Iya<�xa<ya<�za<`}a<�a<�a<Z�a<��a<��a<��a<��a<��a<�a<j�a<G�a<��a<6�a<��a<��a<��a<Ǖa<��a<��a<�a<ʖa<ݗa<ʘa<��a<��a<��a<��a<
�a<F�a<ېa<��a<3�a<u�a<�~a<�za<�va<ta<Wra<�qa<|ra<Bta<	wa<~za<e~a<��a<��a<h�a<b�a<�a<I�a<�a<��a<��a<��a<�a<�a<]�a<��a<�a<=�a<�a<�a<e�a<��a<l�a<��a<5�a<8�a<�a<�a<za<x{a<�va<�qa<^la<fga<�ba<$_a<Q\a<�Za<+Za<�Za<�\a<�_a<ca<�fa<ka<�na<ura<?ua<�wa<�xa<ya<�xa<xa<�va<2ua<�sa<Zra<Nqa<�pa<�pa<�pa<gqa<Wra<Csa<<ta<�ta<�ta<�sa<{ra<.pa<�la<<ia<�da<R`a<�[a<�Wa<�Sa<�Pa<Oa<jNa<Oa<�Pa<�Sa<YWa<�[a<=`a<�  �  �ea<ja<�ma<�pa<�ra<Cta<�ta<�ta</ta<Esa<ora<Zqa<�pa<Upa<}pa<3qa<Pra<�sa<�ua<	wa<�xa<�ya<�za<fza<�ya<�wa<kua<ara<�na<ka<-ga<�ca<(aa<0_a<�^a<�^a<k`a<ca<�fa<,ka<1pa<<ua<.za<�~a<��a<<�a<��a<B�a<$�a<N�a<�a<��a<.�a<��a<��a<��a<N�a<��a<��a<�a<Аa<��a<+�a<V�a<ڕa<��a<y�a<G�a<��a<'�a<R�a<`�a<S�a<�|a<za<(xa<swa<�wa< ya<�{a<6a<,�a<Ƈa<+�a<z�a<R�a<c�a<�a<d�a<8�a<�a<��a<��a<��a<>�a<;�a<��a<:�a<f�a<3�a< �a<��a<a<��a<՜a<^�a<�a<
�a< �a<E�a<�a<�a<��a<@�a<�a<�a<�|a<�za<*za<�za<|a<�~a<.�a<(�a<��a<��a<��a<�a<��a<��a<��a<�a<L�a<b�a<�a<ȗa<?�a<(�a<C�a<�a<�a<��a<��a<��a<��a<��a<�a<7�a<f�a<�a<o�a<N�a<��a<'�a<��a< �a<�{a<Sxa<~ua<�sa<msa<�sa<�ua<uxa<�{a<�a<��a<s�a<�a<��a<��a<�a<�a<�a<��a<n�a<��a<��a<��a<��a<G�a<��a<��a<��a<1�a<Іa<8�a<��a<��a<҆a<L�a<�a<�a<|a<twa<�ra<�ma<�ha<Uda<�`a<�]a<A\a<�[a<_\a<L^a<aa<Mda<@ha<la<�oa<�ra<rua<nwa<\xa<�xa<
xa<wa<�ua<ta<[ra<�pa<�oa<)oa<�na<qoa<pa<-qa<ra<sa<�sa<ta<�sa<Ura<Epa<Hma<�ia<�ea<naa<�\a<�Xa<GUa<SRa<�Pa<Pa<�Pa<4Ra<Ua<�Xa<�\a<daa<�  �  ga<�ja<Zna<�pa<�ra<�sa<ta<�sa<�ra<�qa<*pa<�na<0na<�ma< na<�na<�oa<[qa<[sa<eua<Dwa<�xa<�ya<	za<xya<Kxa< va<Qsa<%pa<�la<@ia<fa<�ca<�aa<-aa<�aa<ca<�ea<'ia<_ma<�qa<�va<i{a<�a<q�a<>�a<T�a<��a<+�a<#�a<��a<��a<чa<A�a<��a<�a<ˇa<݈a<��a<��a<Ɏa<��a<�a<U�a<E�a<6�a<o�a<��a<O�a<U�a<ȉa<�a<��a<5a<�|a<�za<za<lza<�{a<O~a<r�a<N�a<U�a<��a<��a<��a<�a<˙a<�a<�a<�a<5�a<�a<b�a<ەa<Δa<ޓa<��a<̓a<��a<��a<:�a<�a<y�a<��a<p�a<��a<śa<N�a<
�a<̔a<7�a<)�a<�a<F�a<�a<Ea<}}a<�|a<;}a<�~a<@�a<d�a<�a<�a<��a<{�a<��a<�a<]�a<&�a<��a<=�a<�a<P�a<��a<ړa<��a<��a<k�a<j�a<1�a< �a<��a<��a<9�a<�a<p�a<�a<ǖa<�a<�a<w�a<��a<5�a<�a<~a<�za<8xa<�va<va<�va<Uxa<�za<�}a<`�a<�a<��a<��a<a�a<��a<Ӑa<��a<"�a<Ύa<�a<Ɗa<��a<��a<�a<��a<�a<Ԃa<E�a<ԃa<Ʉa<��a<[�a<��a<=�a<��a<
�a<p�a<�|a<�xa<ta<Hoa<�ja<�fa<+ca<�`a<�^a<o^a<!_a<�`a<Aca<ofa<�ia<qma<�pa<�sa<va<Mwa<xa<�wa< wa<�ua<�sa<�qa<�oa<�na<,ma<�la<`la<�la<�ma<�na<Npa<�qa<�ra<sa<sa<ra<rpa<na<�ja<ga<�ba<�^a<�Za<�Wa<Ua<ISa<�Ra<7Sa<�Ta<�Wa<�Za<�^a<�ba<�  �  �ha<la<oa<*qa<�ra<0sa<�ra<ra<�pa<oa<oma<la<ka<lja<�ja<7ka<�la<una<�pa<�ra<;ua<=wa<�xa<�ya<iya<�xa<�va<�ta<ra<�na<�ka<�ha<�fa<$ea<�da<ea<rfa<�ha<la<pa<Qta<�xa<}a<��a<�a<I�a<"�a<ֈa<��a<W�a<L�a<?�a<��a<F�a<��a<҃a<��a<��a<��a<��a<A�a<��a<�a<ܒa<B�a<��a<o�a<w�a<T�a<�a<ʋa<e�a<8�a<	�a<�a</~a<�}a<�}a<#a<Q�a<<�a<�a<��a<��a<��a<ޕa<Q�a<a<��a<S�a<��a<:�a<��a<Ŕa<��a<��a<��a<e�a<��a<t�a<Βa<u�a<z�a<G�a<�a<�a<�a<��a<{�a<��a<�a<��a<B�a<��a<�a<ʄa<t�a<��a<N�a<��a<��a<"�a<-�a<��a<�a<Ǒa<��a<f�a<-�a<C�a<��a<��a<��a<ʖa<۔a<ǒa<�a<|�a<X�a<�a<�a<�a<9�a<ߑa<��a<0�a<��a<:�a<��a<��a<7�a<ؒa<ُa<q�a<c�a<��a<�a<�}a<r{a<�ya<�ya<za<p{a<�}a<��a<΃a<�a<Y�a<��a<�a<�a<��a<�a<��a<�a<��a<G�a<��a<��a<��a<z�a<�a<�a<>�a<�a<A�a<f�a<~�a<�a<:�a<��a<
�a<�a<�}a<?za<va<�qa<�ma<jia<:fa<�ca<Uba<�aa<bba<�ca<fa<ia<
la<coa<8ra<�ta<bva<Ewa<�wa<�va<�ua<�sa<�qa<Qoa<ma<pka<�ia<Uia<ia<�ia<�ja<la<�ma<coa<�pa<�qa<Xra<�qa<�pa<�na<�ka<�ha<ea<Xaa<�]a<}Za</Xa<�Va<.Va<�Va<Xa<gZa<�]a<Saa< ea<�  �  �ja<�ma<�oa<�qa<;ra<9ra<�qa<pa<*na<;la<Mja<kha<8ga<�fa<�fa<|ga<�ha<�ja<�ma<:pa<�ra<yua<jwa<�xa<<ya<ya<xa<<va<�sa<mqa<�na<_la<eja<�ha<�ha<�ha<Uja<�la<�oa<#sa<wa<�za<�~a<�a<��a<t�a<��a<��a<b�a<@�a<��a<M�a<��a<z�a<�a<�a<o�a<�a<Ƀa<V�a<D�a<�a<�a<t�a<+�a<P�a<��a<�a<��a<z�a<�a<0�a<0�a<Åa<�a<�a<��a<ׁa<�a<�a<Їa<Պa<H�a<z�a<z�a<�a<ǘa<��a<ڙa<5�a<�a<��a<Γa<��a<��a<ߍa<��a<R�a<��a<��a<�a<K�a<��a<ϕa<�a<יa<ޚa<6�a<Śa<��a<t�a<��a<��a<h�a<?�a<��a<8�a<Ǆa<>�a<��a<ǅa<�a<v�a<p�a<��a<��a<6�a<F�a<��a<�a<��a<}�a<��a<\�a<�a<��a<N�a<��a<��a<�a<\�a<;�a<��a<ʎa<͐a<ߒa<ʔa<�a<��a<��a<��a<�a<a�a<V�a<�a<��a<`�a<��a<Fa<�}a<�}a<�}a</a<X�a<��a<��a<W�a<�a<1�a<��a<0�a<�a<��a<Z�a<�a<�a<U�a<n�a<�a<�}a<u|a<�{a<�{a<k|a<�}a<Ea<Àa<\�a<��a<#�a<�a<#�a<|�a<a<�{a<(xa<tta<}pa<#ma<�ia<�ga<Vfa<�ea<3fa<�ga<�ia<�ka<�na<Rqa<�sa<�ua<�va<1wa<�va<�ua<�sa<rqa<�na<?la<�ia<�ga<1fa<Bea<>ea<�ea<
ga<�ha<�ja<�la<�na<�pa<Uqa<�qa<�pa<�oa<Yma<�ja<hga<da<�`a<D^a<�[a<�Za<Za<�Za<�[a<2^a<�`a<da<{ga<�  �  �la<(oa<�pa<�qa<�qa<Fqa<pa<�ma<�ka<ia<�fa<�da<.ca<sba<Uba<aca<�da<Xga<ja<Lma<�pa<asa<va<�wa<,ya<wya<ya<�wa<va<1ta<�qa<�oa<+na<&ma<�la<$ma<�na<�pa<isa<cva<	za<t}a<��a<W�a<B�a<��a<��a<��a<��a<��a<�a<�a<4~a<�|a<�{a<�{a<:|a<�}a<�a<ӂa<υa<f�a<��a<��a<	�a<��a<��a<��a<�a<X�a<X�a<�a<j�a<e�a<c�a<V�a<��a<�a<.�a<�a<_�a<��a<�a<��a<A�a<�a<<�a<��a<�a<�a<�a<��a<��a<%�a<�a<މa<ňa<�a<{�a<��a<X�a<��a<[�a<Z�a<ٕa<D�a<�a<ߚa<�a<>�a<�a<��a<J�a<k�a<��a<M�a<A�a<�a<k�a<܈a<܉a<��a<�a<{�a<I�a<��a<×a<�a<ؙa<��a<��a<��a<��a<�a<ގa<�a<��a<��a<^�a<��a<@�a<5�a<�a<;�a<ݍa<��a<��a<��a<ڕa<y�a<�a<�a<�a<}�a<΍a<��a<�a<V�a<t�a<7�a<��a<4�a<�a< �a<�a<��a<ڋa<эa<w�a<3�a<g�a<|�a<�a<��a<��a<z�a<�a<�~a<�{a<�ya<Dxa<�wa<�wa<}xa<"za<�{a<~a<�a<Ła<�a<n�a<M�a<�a<B�a<�}a<�za<Swa<�sa<�pa<�ma<�ka<yja<ja<mja<fka<.ma<oa<�qa<�sa<|ua<�va<Mwa<6wa<va<hta<�qa<oa<�ka<�ha<fa<�ca<ba<�`a<aa<�aa<Hca<^ea<�ga<vja<�la<�na<[pa<)qa<2qa<>pa<�na<xla<ja<ga<Uda<�aa<�_a<�^a<H^a<�^a<�_a<�aa<]da<!ga<*ja<�  �  �na<�pa<�qa<ra<�qa<qpa<mna<�ka<ia<	fa<Eca<�`a<_a<,^a<*^a<_a<�`a<�ca<�fa<Oja<�ma<rqa<�ta<,wa<�xa<�ya<za<�ya<Txa<�va<ua<rsa<�qa<<qa<�pa<fqa<�ra<�ta<�va<�ya<�|a<�a<��a<��a<�a<��a<��a<��a<΃a<��a<Qa<�|a<�za<�xa<�wa<mwa<xa<�ya<�{a<2a<��a<��a<1�a<��a<�a<!�a<��a<F�a<�a<E�a<��a<��a<�a<�a<X�a<s�a<�a<:�a<L�a<��a<�a<[�a<��a<�a<��a<&�a<��a<t�a<o�a<��a<�a<�a<�a<݊a<F�a<�a<t�a<�a<9�a<i�a<��a<9�a<B�a<��a<��a<��a<��a<x�a<+�a<�a<J�a<ǘa<��a<h�a<3�a<�a<G�a<6�a<��a< �a<�a<_�a<{�a<��a<��a<��a<9�a<�a<	�a<S�a<Ǘa<f�a<y�a<=�a<΋a<��a<Ӆa<|�a<�a<��a<�a<4�a<c�a<އa<ߊa<�a<��a<P�a<'�a<1�a<q�a<�a<��a<��a<K�a<�a<t�a<$�a<��a<d�a<�a<O�a<�a<��a<z�a<O�a<0�a<ҏa<��a<��a<Y�a<�a<ڌa<Ɖa<N�a<��a<�~a<P{a<"xa<�ua<ta<csa<�sa<�ta<�va<�xa<A{a<�}a<�a<ށa<�a<,�a<��a<n�a<�a<�|a<za<4wa<Lta<�qa<pa<�na<<na<�na<Boa<�pa<}ra<ta<�ua<5wa<�wa<�wa<�va<jua<sa<�oa<�la<	ia<lea<gba<�_a<�]a<�\a<�\a<�]a<�_a<�aa<�da<�ga<�ja<Ema<ooa<�pa<Mqa<qa<.pa<�na<fla<ja<�ga<�ea<�ca<�ba<�ba<�ba< da<�ea<�ga<9ja<�la<�  �  �pa<�qa<�ra<Ura<Hqa<�oa<�la<ja<�fa<Aca<�_a<']a<G[a<;Za<;Za<-[a<#]a<�_a<�ca<�ga<�ka<�oa<*sa<iva<�xa<Vza<{a<�za<aza<,ya<xa<�va<�ua<ua<�ta<xua<kva<^xa<\za<�|a<�a< �a<�a<��a<Ɔa<��a<�a<X�a<Q�a<�a<�|a<�ya<�va<ua<�sa<ksa<ta<�ua<:xa<�{a<�a<ƃa<(�a<9�a<��a<��a<��a<��a<'�a<��a<Ӕa<k�a<�a<=�a</�a<#�a<��a<5�a<�a<��a<!�a<H�a<.�a<�a<E�a<:�a<J�a<?�a<��a<%�a<a�a<Ўa<:�a<χa<��a<+�a<��a<�a<A�a<��a<ǃa<ʆa<n�a<��a<�a<�a<�a<�a<d�a<�a<v�a<��a<�a<2�a<K�a<{�a<&�a<��a<Őa<ΐa<Ña<��a<��a<h�a<�a<��a<j�a<�a<X�a<��a<ږa<��a<��a<��a<�a<E�a<�a<�a<#~a<�}a<
~a<sa<��a<��a<�a<��a<�a<Бa<d�a<�a<�a<�a<�a<Ĕa<ɒa<Ԑa<��a<݌a<V�a<K�a<��a<��a<��a<�a<��a<�a<h�a<a�a<͑a<��a<b�a<��a<��a<J�a<Z�a<�a<�{a<�wa<]ta<�qa<pa<aoa<�oa<�pa<�ra<�ua<{xa<�{a<i~a<��a<a�a<�a<m�a<��a<�a<a<�|a<5za<�wa<�ua<�sa<�ra<7ra<Jra<	sa<�sa<iua<�va<�wa<�xa<�xa<]xa<�va<�ta<�qa<Xna<Kja<>fa<_ba<�^a<�[a<�Ya<�Xa<�Xa<�Ya<�[a<o^a<�aa<ea<�ha<�ka<dna<]pa<�qa<ra<Zqa<gpa<�na<�la<�ja<)ia<�ga<�fa<�fa<�fa<�ga<;ia<
ka<ma<�na<�  �  Tra<sa<3sa<jra<qa<�na<�ka<8ha<eda<�`a<(]a<CZa<Xa<�Va<�Va<�Wa<�Ya<]a<�`a<ea<�ia<na<ra<�ua<�xa<yza<�{a<1|a<|a<c{a<zza<iya<�xa<)xa<"xa<�xa<�ya<m{a<B}a<�a<ځa<�a<��a<φa<�a<��a<��a<i�a<΀a<�}a<Nza<*wa<3ta<�qa<�pa< pa<�pa<kra<0ua<�xa<�|a<m�a<)�a<��a<��a<&�a<��a<=�a<8�a<4�a<��a<��a<x�a<&�a<9�a<d�a<H�a<u�a<8�a<y�a<�a<Öa<m�a<ۙa<��a<�a<w�a<-�a<&�a<�a<��a<Ōa<Ĉa<
�a<��a<
a<7}a<v|a<�|a<]~a<׀a<�a<ԇa<Ӌa<��a<��a<!�a<Ǚa<v�a<��a<��a<�a<�a<��a<��a<b�a<?�a<I�a<�a<�a<�a<�a<Q�a<ۘa<4�a<5�a<��a<��a<m�a<��a<�a<��a<Ύa<��a<o�a<|�a<#a<{|a<�za< za<�za<G|a<�~a<�a<��a<w�a<S�a<��a<��a<˕a<�a<��a<T�a<w�a<��a<L�a<k�a<ʏa<x�a<��a<N�a<F�a<�a<ڎa<"�a<Z�a<Y�a<ݒa<�a<�a<h�a<�a<��a<ǆa<c�a<�}a<3ya<�ta<Xqa<�na<�la<�ka<bla<�ma< pa<�ra<"va<�ya<�|a<�a<�a< �a<��a<��a<~�a<��a<�~a<�|a<�za<�xa<wa<va<wua<vua<�ua<�va<�wa<�xa<�ya<�ya<�ya<�xa<�va<#ta<�pa<�la<Aha<�ca<�_a<�[a<�Xa<�Va<jUa<uUa<�Va<�Xa<�[a<3_a<�ba<�fa<eja<�ma<pa<�qa<�ra<�ra<�qa<�pa<Poa<�ma<la<�ja<ja<�ia<ja<�ja<#la<�ma<oa<qa<�  �  bsa<�sa<�sa<�ra<�pa<�ma<�ja<�fa<�ba<�^a<�Za<�Wa<]Ua<0Ta<Ta<Ua<JWa<�Za<�^a<7ca<ha<�la<Yqa< ua<]xa<�za<I|a<!}a<+}a<�|a<V|a<�{a<{a<�za<�za<L{a<q|a<�}a<�a<��a<s�a<F�a<��a<��a<u�a<ņa<�a<ʂa<�a<B|a<�xa<ua<�qa<toa<�ma<]ma<na<�oa<�ra<qva<�za<�a<��a<~�a<��a<z�a<��a<��a<ؗa<9�a< �a<E�a<��a<��a<��a<!�a<ʓa<�a<�a<ڕa<P�a<��a<�a<��a<��a<��a<��a< �a<j�a<r�a<r�a<N�a<	�a<ւa<Za<b|a<�za<�ya<6za<�{a<]~a<Ɓa<Ʌa<N�a<��a<֒a<d�a<[�a<��a<�a<��a<)�a<x�a<I�a<.�a<Ƙa<��a<�a<��a<��a<g�a<G�a<��a<��a<��a<D�a<��a<��a<��a<a�a<S�a<ˑa<w�a<�a<u�a<D�a<�|a<�ya<xa<~wa<�wa<�ya<l|a<�a<ăa<��a<�a<��a<��a<��a<U�a<(�a<D�a<��a<��a<(�a<��a</�a<�a<%�a<Ϗa<�a<n�a<:�a<:�a<�a<��a<�a<��a<h�a<��a<��a<	�a<��a<�a<|a<wa<�ra<�na<�ka<ja<Pia<�ia<Aka<�ma<�pa<�ta<!xa<�{a<�~a<>�a</�a<�a<3�a<��a<A�a<��a<�~a<�|a<{a<�ya<�xa<xa<(xa<]xa< ya<�ya<jza<�za<�za<8za<�xa<�va<gsa<�oa<jka<�fa<ba<h]a<}Ya<Va<�Sa<�Ra<�Ra<�Sa<OVa<lYa<(]a<kaa<}ea<~ia<�la<�oa<�qa<�ra<bsa<�ra<3ra<�pa<�oa<tna<oma<�la<lla<�la<~ma<�na<�oa<6qa<�ra<�  �  [ta<vta<�sa<�ra<�pa<�ma<ja<�ea<�aa<q]a<�Ya<`Va<�Sa<�Ra<yRa<�Sa<�Ua<;Ya<Y]a<�aa<�fa<�ka<�pa<�ta<Gxa<�za<�|a<�}a<'~a<~a<z}a<�|a<`|a<>|a<J|a<�|a<�}a<>a<܀a<ςa<��a<W�a<b�a<�a<��a<؆a<̈́a<D�a<�~a<Q{a<xwa<�sa<�pa<na<Ola<�ka<^la<7na<-qa<ua<�ya<�~a<��a<��a<b�a<9�a<��a<Ȗa<:�a<�a<�a<y�a<��a<��a< �a<��a<i�a<��a<P�a<=�a<��a<ٙa<�a<��a<I�a<��a<�a<�a<!�a<��a<��a<B�a<a<��a<�}a<�za<ya</xa<�xa<4za<�|a<n�a<��a<�a<��a<�a<��a<8�a<a<0�a<��a<�a<��a<t�a<U�a<�a<.�a<j�a<@�a<?�a<ܘa<��a<��a<��a<ʜa<=�a<�a<?�a<Ța<D�a<��a<�a<��a<�a<4�a<�~a<>{a<Rxa<�va<�ua<vva<+xa<�za<�~a<�a<�a<+�a<E�a<��a<��a<�a<}�a<٘a<��a<��a<K�a<�a<��a<��a<��a<p�a<g�a<בa<u�a<_�a<&�a<��a<��a<�a<��a<��a<O�a<��a<�a<�a<�za<�ua<Dqa<^ma<Qja<fha<�ga<.ha<�ia<Vla<�oa<?sa<.wa<�za<X~a<��a<5�a<>�a<��a<5�a<M�a<��a<�a<~a<z|a<{a<5za<�ya<�ya<�ya<Oza<�za<�{a<�{a<�{a<�za<�xa<�va<sa<8oa<�ja<�ea<�`a<.\a<Xa<�Ta<ZRa<#Qa<6Qa<wRa<�Ta<Xa<�[a<7`a<�da<�ha<nla<�oa<�qa</sa<�sa<�sa<Rsa<#ra< qa<�oa<�na<-na<na<4na<�na<�oa<)qa<^ra<�sa<�  �  �sa<�sa<�sa<sra<�pa<�na<�ka<	ia<�ea<�ba<�_a<P]a<�[a<�Za<�Za<�[a<`]a<�_a<Dca<�fa<�ja<�na<(ra<�ua<Wxa<vza<)|a<}a<n}a<w}a<q}a<5}a<}a<}a<(}a<�}a<�~a<�a<5�a<Ȃa<*�a<u�a<y�a<$�a<��a<>�a<�a<2�a<؀a<=~a<s{a<�xa<{va<�ta<�sa<Psa<�sa<tua<�wa<�za<�~a<t�a<��a<l�a<	�a<=�a<��a<��a<	�a<��a<��a<i�a<�a<z�a<�a<��a<a<�a<��a<]�a<>�a<?�a<�a<��a<�a<�a<�a<��a<u�a<��a<��a<]�a<�a<�a<��a<ҁa<Z�a<�a<�a<V�a<V�a<�a<_�a<��a<D�a<��a<��a<�a<ۚa<7�a<ٜa<Ӝa<d�a<ћa<�a<�a<��a<͘a<��a<��a<3�a<��a<y�a<)�a<��a<��a<�a<R�a<�a<	�a<��a<U�a<�a<h�a<��a<��a<��a<pa<	~a<�}a<�}a<'a<+�a<�a<��a<.�a<r�a<L�a<!�a<#�a<��a<��a<��a<S�a<��a<ƕa<��a<��a<ܒa<�a<ۑa<��a<�a<\�a<�a<?�a<w�a<`�a<�a<��a<��a<L�a<4�a<��a<��a<�~a<�za<wa<�sa<�qa<pa<Xoa<�oa<�pa<dra<�ta<rwa<Aza<�|a<aa<k�a<��a<��a<�a<R�a<p�a<5�a<�a<h~a<(}a<�{a<!{a<�za<dza<tza<�za<�za<{a<'{a<�za<za<�xa<�va<ta<�pa<9ma<jia<�ea<ba<�^a<\a<CZa<OYa<JYa<0Za<�[a<X^a<Waa<bda<�ga<�ja<�ma<�oa<�qa<�ra<Zsa<>sa<�ra<"ra<Tqa<kpa<�oa<2oa<9oa<8oa<�oa<�pa<�qa<hra<sa<�  �  �sa<�sa<bsa<vra<�pa<�na<Bla<<ia<	fa<�ba<`a<�]a<\a<,[a<[a<\a<�]a<f`a<}ca<)ga<�ja<�na<�ra<�ua<Zxa<rza<�{a<�|a<Y}a<j}a<}a<�|a<z|a<�|a<�|a<^}a<2~a<ea<րa<r�a<��a<o�a<N�a<��a<ۆa<P�a<�a<Q�a<
�a<k~a<�{a<ya<�va<ua<ta<�sa<qta<�ua<Dxa<K{a<�~a<��a<��a<��a<5�a<-�a<a<��a<Ŗa<]�a<��a<A�a<��a<%�a<��a<J�a<L�a<��a<�a<̖a<�a<�a<��a<��a<ޚa<��a<ߙa<�a<n�a<�a<ߐa<��a<G�a<�a<n�a<B�a<׀a<A�a<��a<ˁa<΃a<q�a<��a<�a<t�a<ȓa<��a<	�a<�a<�a<��a<��a<b�a<��a<��a<��a<��a<o�a<J�a<J�a<��a<<�a<�a<ܚa<��a<ޛa<��a<�a<�a<�a<��a<��a<B�a<��a<$�a<ބa<�a<�a<�~a<�}a<d~a<�a<��a< �a<3�a<h�a<��a<��a<"�a<%�a<��a<S�a<|�a<>�a<��a<m�a<X�a<*�a<U�a<��a<h�a<M�a<��a<��a<��a<�a<q�a<5�a<��a<x�a<��a<?�a<S�a<͆a<�a<�~a<	{a<�wa<tta<ra<�pa<�oa<pa<qa<�ra<ua<�wa<qza<#}a<�a<[�a<˂a<v�a<��a<)�a<g�a<�a<�a<~a<�|a<{{a<�za<za<�ya<�ya<Eza<�za<{a<{a<�za<�ya<�xa<�va<�sa<�pa<gma<�ia<�ea<5ba<$_a<�\a<�Za<�Ya<�Ya<�Za<W\a<�^a<�aa<�da<�ga<ka<�ma<�oa<�qa<�ra<&sa<sa<�ra<�qa<�pa<�oa<Poa<�na<�na<�na<aoa<pa<*qa<ra<sa<�  �  �ra<esa<$sa<wra<qa<oa<�la<�ia<�fa<�ca<!aa<�^a<"]a<[\a<K\a<@]a<�^a<�aa<�da<"ha<�ka<_oa<�ra<�ua<xxa<fza<�{a<u|a<�|a<�|a<|a<�{a<�{a<u{a<�{a<|a<}a<T~a<�a<w�a<�a<��a<��a<��a<��a<d�a<3�a<��a<��a<a<�|a<za<�wa<9va<,ua<�ta<�ua<wa<\ya<\|a<�a<��a<r�a<'�a<��a<]�a<ғa<m�a<v�a<Ԗa<Ӗa<Z�a<��a<+�a<��a<9�a<�a<b�a<�a<ϕa<��a<�a<�a<�a<o�a<d�a<ϙa<��a<��a<\�a<g�a<c�a<C�a<�a<��a<X�a<�a<q�a<́a<�a<�a<{�a<~�a<ލa<	�a<A�a<��a</�a<�a<כa<V�a<�a<��a<��a<��a<��a<�a<Z�a<��a<6�a<��a<B�a<$�a<�a<Кa<3�a<j�a<��a<�a<+�a<Օa<�a<Џa<��a<�a<�a<0�a<��a<�a<%a<�a<��a<��a<#�a<,�a<=�a<*�a<�a<P�a<D�a<~�a<�a<�a<��a<��a<q�a<k�a<0�a<I�a<��a<$�a<8�a<x�a<�a<��a<�a<��a<��a<X�a<T�a<ӏa<n�a<��a<V�a<��a<�a<�{a<�xa<�ua<1sa<�qa<�pa<&qa<*ra<�sa<va<�xa<3{a<�}a<�a<��a<܂a<Z�a<O�a<��a<��a<&�a<�~a<}a<�{a<kza<rya<�xa<�xa<�xa<Yya<�ya<$za<Wza<<za<�ya<sxa<�va<#ta<eqa<�ma<pja<�fa<;ca<?`a<�]a<�[a<�Za<�Za<�[a<r]a<�_a<vba<�ea<�ha<�ka<na<pa<�qa<ura<�ra<zra<�qa<�pa<pa<oa<=na<�ma<qma<�ma<Rna<!oa<0pa< qa<Ira<�  �  ra<�ra<�ra<Cra<Eqa<�oa<Xma<�ja<ha<Vea<�ba<�`a< _a<S^a<U^a<4_a<�`a<-ca<)fa<via<�la<\pa<|sa<kva<�xa<)za<?{a<�{a<�{a<Y{a<�za<.za<�ya<�ya<�ya<1za<{a<�|a<~a<�a<݁a<��a<��a<�a<k�a<<�a<��a<.�a<Z�a<)�a<�}a<�{a<�ya<xa<*wa<�va<�wa<ya<B{a<�}a<j�a<ڄa<{�a<��a<�a<ّa<��a<*�a<��a<�a<a</�a<V�a<`�a<Œa<;�a<#�a<g�a<�a<�a<6�a<��a<�a<�a<��a<�a<��a<��a<*�a<ޔa<X�a<s�a<��a<Éa<*�a<J�a<��a<s�a<ǃa<�a<��a<�a<�a<��a<�a<�a<��a<v�a<��a<y�a<��a<<�a<m�a<^�a<'�a<�a<�a<W�a<�a<0�a<��a<}�a<��a<��a<��a<V�a<a<��a<��a<`�a<i�a<��a<֐a<��a<��a<��a<��a<��a<��a<0�a<��a<��a<f�a<͆a<��a<P�a<'�a<��a<�a<Z�a<B�a<��a<g�a<��a<z�a</�a<��a<u�a<e�a<��a<;�a<8�a<��a<=�a<"�a<�a<��a<�a<͑a<�a<��a<ڍa</�a<�a<��a<
�a<�}a</za<jwa<0ua<�sa<sa<&sa<ta<}ua<�wa<�ya<<|a<�~a<l�a<�a<��a<�a<ӂa<�a<��a<�~a</}a<N{a<�ya<mxa<�wa<�va<�va<,wa<�wa<Uxa<�xa<Yya<�ya<(ya<3xa<�va<�ta<�qa<�na<ka<ha<�da<�aa<�_a<�]a<�\a<�\a<�]a<?_a<Vaa<�ca<�fa<�ia<2la<�na<\pa<yqa<ra<4ra<�qa<�pa<�oa<tna<Ama<gla<�ka<�ka<�ka<wla<\ma<�na<�oa<qa<�  �  �pa<�qa<Xra</ra<eqa<)pa<?na<?la<�ia<>ga<�da<�ba<�aa<�`a<�`a<�aa<Tca<nea<@ha<Ika<ina<�qa<Kta<�va<�xa<za<�za<�za<qza<�ya<ya<xa<�wa<wa<&wa<�wa<�xa<?za<�{a<~a<�a<�a<�a<�a<"�a<1�a<�a<Ԅa<g�a<��a<za<�}a<�{a<|za<�ya<wya<za<s{a<�}a<+�a<f�a<��a<��a<�a<ďa<7�a<��a<�a<�a<�a<b�a<k�a<h�a<?�a<��a<��a<��a<�a<��a<ӑa<�a<ʔa<1�a<��a<��a<B�a<_�a<��a<��a<��a<��a<��a<S�a<Ћa<f�a<��a<c�a<��a<?�a<Y�a<�a<9�a<�a<��a<��a<��a<�a<��a<��a<�a<��a<�a<ݘa<��a<�a<��a<��a<Ԓa<��a<��a<Y�a<F�a<w�a<ޖa<�a<,�a<��a<�a<��a<��a<�a<��a<E�a<6�a<u�a<��a<E�a<u�a<!�a<��a<�a<�a<��a<�a<U�a<׍a<~�a<q�a<a�a<g�a<�a<	�a<]�a<V�a<֒a<[�a<��a<5�a<�a<�a<ًa<��a<c�a<�a<&�a<,�a<�a<͐a<�a<��a<��a<'�a<Ջa<)�a<%�a<��a<�a<Z|a<�ya<�wa<-va<�ua<�ua<}va<�wa<�ya<�{a<�}a<�a<�a<e�a<��a<ւa<�a<Հa<+a<8}a<A{a<.ya<�wa<�ua<ua<�ta<hta<�ta<tua<~va<=wa<xa<xxa<xxa<xa<�va</ua<�ra<'pa<ma<�ia<�fa<da<	ba<J`a<�_a<m_a<1`a<�aa<vca<�ea<Hha<ka<$ma<#oa<�pa<jqa<�qa<9qa<�pa<9oa<�ma<kla<ka<ja<;ia<2ia<Bia<ja<&ka<�la<na<~oa<�  �  �oa<�pa<�qa<ra<�qa<�pa<_oa<�ma<xka<aia<Uga<�ea<ada<�ca<�ca<�da<fa<%ha<�ja<ema<)pa<�ra<_ua<twa<�xa<�ya<�ya<�ya<�xa<�wa<�va<�ua<�ta<Jta<9ta<�ta<�ua<lwa<|ya<�{a<~a<m�a<��a<E�a<��a<?�a<F�a<ƅa<��a<!�a<��a<�a<X~a<5}a<z|a<w|a<}a<d~a<f�a<҂a<��a<��a<��a<H�a<��a<��a<֓a<v�a<F�a<ܓa<��a<n�a<�a<Ԏa<��a<��a<��a<�a<͍a<�a<��a<�a<M�a< �a<��a<y�a<�a<�a<�a<��a<ٔa<��a<n�a<�a<�a<x�a<`�a<�a<8�a<)�a<a<Ía<�a<��a<�a<�a<ݘa<�a<��a<x�a<Йa<a<)�a<w�a<ɓa<,�a<�a<��a<��a<͏a<��a<��a<�a<��a<L�a<ɗa<ɘa<^�a<r�a<ۘa<��a<ƕa<��a<�a<��a<�a<��a<=�a<�a<��a<�a<އa<_�a<=�a<q�a<��a<��a<��a<�a<��a<Օa<C�a<Y�a<ݒa< �a<�a<9�a<��a<�a<+�a<��a<�a<��a<��a<ߋa<*�a<n�a<��a<
�a<;�a<��a<��a<ǌa<O�a<��a<ńa<��a<�~a<�|a<za<-ya<�xa<}xa<4ya<Wza<�{a<�}a<Ha<Ҁa<�a<Âa<��a<d�a< �a<�a<�}a<;{a<�xa<�va<�ta<+sa<
ra<�qa<�qa<+ra<sa<3ta<Yua<�va<ewa<�wa<�wa<�va<�ua<�sa<`qa<�na<la<6ia<�fa<�da<Gca<�ba<fba<ca<Jda< fa<ha<?ja<^la<Dna<�oa<�pa<Sqa<qa<Spa</oa<�ma<�ka<ja<}ha<@ga<efa<fa<efa<Hga<�ha<-ja<�ka<�ma<�  �  �ma<�oa<�pa<�qa<�qa<�qa<�pa<%oa<�ma<�ka<�ia<lha<hga<�fa<�fa<�ga<ia<�ja<#ma<�oa<ra<rta<�va<�wa<	ya<`ya<2ya<�xa<Fwa<va<]ta<sa<�qa<Cqa<+qa<�qa<�ra<Yta<�va<%ya<|a<�~a<8�a<q�a<�a<>�a<��a<��a<��a<߄a<��a<4�a<
�a<�a<�a<�a<D�a<��a<1�a<��a<�a<֊a<K�a<��a<��a<��a<ߓa<�a<��a<u�a<��a<r�a<��a<�a<��a<��a<��a<�a<Ǌa<�a<��a<�a<m�a<j�a<S�a<Ǘa<��a<�a<��a<ʗa<T�a<��a<��a<��a<�a<[�a<��a<�a<o�a<=�a<��a<c�a<f�a<��a<��a<X�a<��a<E�a<j�a<֙a<�a<6�a<X�a<B�a<+�a<O�a<Ѝa<��a<w�a<Ōa<{�a<Îa<}�a<m�a<v�a<1�a<̗a<��a<:�a<�a<I�a<�a<,�a<1�a<��a<��a<��a<E�a<U�a<ىa<+�a<͊a<#�a<ɍa<��a<��a<@�a<��a<s�a<וa<z�a<��a<)�a<-�a<$�a<��a<��a<��a<�a<�a<��a<�a<|�a<чa<E�a<�a<��a<�a<6�a<��a<��a<ێa<��a<��a<^�a<�a<"�a<��a<Qa<�}a<[|a<�{a<�{a<�{a<}a<A~a<�a<�a<=�a<�a<(�a<�a<сa<\�a<B~a<�{a<?ya<hva<�sa<�qa<)pa<�na<zna<�na<(oa<bpa<�qa<ysa<�ta< va<�va<@wa<wa<va<�ta<�ra<�pa<@na<�ka<�ia<�ga<�fa<�ea<�ea<fa<ga<�ha<]ja<`la<na<�oa<�pa<+qa<*qa<upa<eoa<�ma<�ka<�ia<{ga<�ea<*da<`ca<�ba<^ca<5da<�ea<�ga<�ia<�ka<�  �  Tla<�na<bpa<�qa<6ra<.ra<�qa<�pa<hoa<�ma<�la<Xka<zja< ja<ja<�ja<la<�ma<�oa<�qa<�sa<�ua<vwa<�xa<(ya<ya<xxa<$wa<�ua<�sa<
ra<apa<oa<*na<�ma<{na<�oa<~qa<�sa<�va<�ya<�|a<�a<d�a<��a<)�a<�a<P�a<B�a<��a<��a<��a<��a<�a<��a<��a<Z�a<��a<>�a<O�a<��a<Ȍa<�a<�a<h�a<��a<ғa<z�a<��a<�a<,�a<>�a<�a<M�a<Їa<a<k�a<��a<��a<I�a<R�a<��a<C�a<��a<�a<��a<I�a<�a<0�a<��a<Зa<U�a<ǔa<6�a<��a<q�a<��a<<�a<}�a<H�a<��a<�a<a<��a<2�a<{�a<;�a<��a<>�a<K�a<��a<��a<Y�a<��a<��a<��a<܊a<��a<[�a<��a<y�a<��a<�a<&�a<d�a<��a<��a<�a<�a<R�a<�a<�a<̖a<
�a<,�a<\�a<��a<W�a<`�a<��a<.�a<�a<��a<e�a<�a<^�a<Ŕa<��a<�a<��a<5�a<ܓa<̑a<��a<�a<`�a<�a<��a<��a<�a<��a<��a<��a<�a<Ća<߈a<Ɗa<��a<(�a<.�a<��a<W�a<P�a<�a<�a<ֈa<��a<a�a<X�a<��a<ka<�~a<�~a<a<�a<ʀa<Ɓa<тa<��a<a<��a<܂a<h�a<fa<�|a<�ya<wa<�sa<<qa<�na<�la<�ka<Ika<yka<ala<�ma<_oa<Oqa<sa<�ta<1va<�va< wa<�va<�ua<Uta<_ra<Zpa<Vna<ila<�ja<�ia<�ha<�ha<ia<	ja<Jka<�la<:na<�oa<�pa<Nqa<|qa<�pa<�oa<.na<la<�ia<Rga<�da<�ba<7aa<#`a<�_a<$`a<4aa<�ba<�da<iga<�ia<�  �  ka<ima<�oa<Bqa<lra<�ra<�ra<-ra<&qa<&pa<�na<�ma<Cma<�la<7ma<�ma<�na<Ipa<ra<�sa<�ua<Dwa<Vxa<4ya<7ya<�xa<�wa<va<;ta<�qa<�oa<�ma<Xla<Tka<�ja<zka<�la<�na<3qa<jta<�wa<!{a<�~a<[�a<$�a<�a<s�a<�a<Z�a< �a<��a<��a<"�a<Ʌa<l�a<��a<d�a<\�a<�a<��a<֌a<��a<��a<7�a<8�a<�a<��a<�a<��a<׏a<��a<!�a<�a<��a<�a<̓a<j�a<��a<Äa<��a<��a<��a<5�a<?�a<͓a<�a<�a<	�a<��a<��a<�a<�a<͖a<�a</�a<C�a<k�a<Y�a<f�a<�a</�a<f�a<�a<S�a<��a<z�a<��a<ۚa<�a<��a<��a<l�a<��a<ߎa<:�a<։a<�a<��a<X�a<��a<��a<H�a<v�a<�a<��a<U�a<l�a<n�a<��a<��a<��a<�a<5�a<Ȗa<_�a<��a<N�a<!�a<A�a<�a<�a<��a<��a<��a<��a<�a<�a<�a<��a<�a<ؔa<�a<��a<"�a<�a<;�a<U�a<�a<(�a<�a<�a<�a<�a<X�a<��a<��a<!�a<p�a<�a<��a<W�a<��a<�a<�a<��a<��a<�a<Ća<�a<q�a<h�a<ˁa<v�a<ځa<<�a<�a<��a<i�a<a<��a<�a<��a<�a<c~a<�{a<_xa<�ta<�qa<�na<&la< ja<�ha<Kha<�ha<�ia<ka<;ma<Aoa<�qa<�sa<Hua<�va<wa<Gwa<�va<�ua<ta<_ra<�pa<�na<�ma<Pla<�ka<�ka<�ka<�la<�ma<�na<	pa<"qa<�qa<ra<�qa<�pa<Poa<ma<�ja<�ga<4ea<�ba<*`a<u^a<(]a<�\a<(]a<p^a<+`a<�ba<Gea<ha<�  �  �ia<�la<3oa<(qa<�ra<]sa<�sa<Zsa<�ra<�qa<�pa</pa<�oa<eoa<�oa<)pa<=qa<{ra<ta<�ua<*wa<exa<Mya<�ya<Dya<�xa<wa<ua<�ra<Ipa<�ma<�ka<�ia<�ha<�ha<�ha<=ja<Ula<�na<`ra<�ua<�ya<M}a<��a<��a<�a<��a<وa<l�a<s�a<A�a<Ԉa<E�a<�a<�a<)�a<шa<ىa<Q�a<֌a<��a<��a< �a<G�a<�a<+�a<��a<��a<Ԑa<��a<�a<i�a<�a<k�a<��a<e�a<�a<=�a<X�a<.�a<��a<��a<��a<ďa<Ȓa<s�a<��a<�a<	�a<p�a<'�a<��a<��a<��a<]�a<��a<�a<��a<�a<��a<k�a<��a<Ԙa<�a<�a<��a<��a<��a<��a<4�a<��a<�a<�a<�a<!�a<��a<��a<U�a<σa<!�a<9�a<��a<Z�a<�a<��a<�a<��a<�a<��a<��a<!�a<�a<b�a<a�a<0�a<ȕa<��a<��a<ƒa<s�a<��a<�a<��a<��a<��a<��a<5�a<v�a<�a<�a<��a<u�a<��a<��a<j�a<N�a<4�a<��a<�~a<u}a<�|a<U}a<v~a<�a<�a<��a<��a<2�a<`�a<J�a<S�a<�a<ُa<-�a<�a<y�a<a<�a<`�a<�a<ބa<8�a<�a<�a<[�a<��a<��a<a<҅a<j�a<Z�a<��a<��a<�}a<yza<�va<7sa<�oa<Zla<�ia<�ga<Ifa<�ea<+fa<Fga<�ha<Eka<�ma<.pa<�ra<�ta<Lva<'wa<�wa<uwa<�va<�ua<(ta<�ra<qa<�oa<�na<>na<na<bna<�na<�oa<�pa<�qa<Zra<�ra<�ra<�qa<�pa<�na<Cla<}ia<dfa<[ca<s`a<�]a<�[a<�Za<OZa<�Za<�[a<�]a<k`a<cca<xfa<�  �  �ha<�ka<�na<�pa<�ra<�sa<Yta<=ta<�sa</sa<�ra<�qa<�qa<iqa<xqa<*ra<sa<=ta<�ua<�va<Qxa<5ya<�ya<�ya<tya<2xa<�va<Wta<�qa<(oa<gla<ja</ha<�fa<�fa<�fa<Dha<dja<\ma<�pa<�ta<�xa<b|a<�a<�a<�a<�a<N�a<"�a<t�a<s�a<*�a<	�a<ǉa<މa<"�a<Ċa<ԋa<�a<��a<�a<��a<
�a<��a<��a<k�a<��a<,�a<Z�a<͍a<�a<9�a<?�a<ςa<��a<ga<�~a<=a<Y�a<U�a<�a<��a<r�a<��a<�a<�a<F�a<@�a<Z�a<�a<�a<��a<a<��a<#�a<`�a<�a<��a<�a<n�a<*�a<7�a<�a<*�a<Лa<5�a<�a<3�a<a<��a<+�a<�a<�a<��a<y�a<܅a<��a<`�a<Áa<)�a<<�a<=�a<��a<��a<�a<�a<�a<X�a<i�a<әa<��a<a<E�a<��a<h�a<m�a<J�a<l�a<˔a<X�a<��a<ݔa<{�a<E�a<�a<×a<�a<�a<c�a<D�a<O�a<�a< �a<��a<I�a<��a<��a<�~a<�|a<y{a<�za<]{a<�|a<�~a<րa<��a<��a<G�a<�a<��a<W�a<#�a<M�a<�a<�a<��a<�a<��a<�a<�a<؆a<+�a<�a<߅a<%�a<_�a<��a<͆a<��a<�a<��a<Âa<�a<5}a<�ya<�ua<ra<na<�ja<�ga<�ea<Dda<�ca<-da<lea<Uga<�ia<~la<oa<�qa<$ta<�ua<Swa<�wa<xa<uwa<�va<Sua<ta<�ra<�qa<�pa<$pa<pa<Cpa<�pa<rqa<	ra<�ra<Jsa<ysa<sa<ra<�pa<>na<�ka<~ha<Rea<ba<�^a<0\a<Za<�Xa<CXa<�Xa<�Ya<!\a<�^a<�aa<cea<�  �  ha<yka<_na<�pa<�ra<ta<�ta<�ta<�ta<*ta<�sa<�ra<�ra<ra<�ra<@sa<"ta<4ua<�va<�wa<ya<�ya<9za<za<hya<
xa<3va<�sa<qa<:na<uka<ia<ga<�ea<Yea<�ea<ga<Nia<Bla<�oa<�sa<�wa<�{a<�a<��a<ׅa<��a<��a<��a<8�a<R�a<(�a<��a<Ŋa<�a<I�a<��a<�a<�a<��a<�a<��a<֓a<��a<֔a<��a<��a<��a<�a<A�a<G�a<@�a<>�a<��a<�a<D~a<�}a<~a<;a<9�a<�a<�a<��a<�a<��a<��a<�a</�a<��a<P�a<��a<i�a<��a<��a<�a<q�a<��a<�a<�a<{�a<#�a<'�a<�a<�a<��a<��a<8�a<<�a<��a<i�a<��a<��a<�a<��a<u�a<a<��a<0�a<��a<��a<&�a<%�a<��a<��a<�a<[�a<{�a<�a<D�a<יa<ǚa<�a<�a<j�a<c�a<d�a<D�a<y�a<�a<��a<��a<�a<s�a<?�a<�a<��a<��a<c�a<��a<8�a<&�a<��a<��a<�a<\�a<˃a<��a<�}a<�{a<Jza<�ya<2za<p{a<f}a<�a<Ăa<ąa<��a<u�a<��a<D�a<5�a<��a<W�a<��a<��a<�a<��a<�a<�a<��a<^�a<��a<�a<�a<^�a<��a<��a<�a<0�a<��a<��a<�a<�|a<ya<ua<qa<ma<�ia<�fa<xda<ca<�ba<ca<Qda<Ifa<�ha<�ka<una<Pqa<�sa<�ua<Awa<xa<Txa<xa<qwa<Eva<ua<�sa<�ra<�qa<oqa<1qa<Qqa<�qa<bra<sa<�sa<�sa<�sa<Ksa<$ra<bpa<
na<@ka<�ga<yda<
aa<�]a<[a<�Xa<�Wa<Wa<�Wa<�Xa<
[a<�]a<aa<�da<�  �  �ga<!ka<Qna<�pa<�ra<8ta<�ta<ua<�ta<xta<�sa<fsa<"sa<�ra<>sa<�sa<�ta<�ua<�va<xa<ya<�ya<rza<>za<^ya<xa<va<�sa<�pa<�ma<Ika<�ha<�fa<Uea<�da<Cea<�fa<�ha<�ka<�oa<vsa<�wa<�{a<ga<�a<ׅa<�a<Չa<��a<H�a<i�a<w�a<R�a<V�a<k�a<��a<k�a<^�a<��a<�a<l�a<��a<�a<��a<�a<��a<��a<�a<��a<�a<�a< �a<�a<N�a<4a<�}a<;}a<�}a<�~a<a<��a<Նa<7�a<ߍa<L�a<z�a<(�a<�a<��a<��a<��a<n�a<�a<P�a<��a<��a<b�a<^�a<f�a<�a<��a<��a<f�a<
�a<��a<��a<o�a<=�a<��a<f�a<b�a<T�a<ڍa<}�a<8�a<O�a< �a<��a<#�a<z�a<��a<��a<e�a<��a<Ìa<&�a<#�a<�a<C�a<ҙa<��a<E�a<�a<k�a<��a<��a<��a<�a<;�a<�a<��a<}�a<��a<��a<+�a<��a<ǘa<��a<��a<.�a<4�a<��a<D�a<Ԋa<�a<��a<4�a<J}a<({a<�ya<Kya<�ya<{a<�|a<�a<��a<��a<��a<*�a<��a<D�a<D�a<Րa<|�a<Əa<��a<e�a<�a<��a<p�a<n�a<҇a<x�a<p�a<r�a<��a<��a<��a<2�a<r�a<Ǆa<��a<�a<�|a<�xa<�ta<�pa<�la<>ia<Bfa<�ca<�ba<%ba<�ba<�ca<�ea<�ha<Bka<Hna<qa<�sa<�ua<0wa<.xa<�xa<1xa<vwa<�va<nua<0ta<Fsa<Era<�qa<�qa<�qa<.ra<�ra<[sa<�sa<ta<ta<�sa<$ra<_pa<na<�ja<�ga<:da<�`a<�]a<�Za<}Xa<Wa<�Va<Wa<nXa<�Za<v]a<�`a<?da<�  �  ha<yka<_na<�pa<�ra<ta<�ta<�ta<�ta<*ta<�sa<�ra<�ra<ra<�ra<@sa<"ta<4ua<�va<�wa<ya<�ya<9za<za<hya<
xa<3va<�sa<qa<:na<uka<ia<ga<�ea<Yea<�ea<ga<Nia<Bla<�oa<�sa<�wa<�{a<�a<��a<ׅa<��a<��a<��a<8�a<R�a<(�a<��a<Ŋa<�a<I�a<��a<�a<�a<��a<�a<��a<֓a<��a<֔a<��a<��a<��a<�a<A�a<G�a<@�a<>�a<��a<�a<D~a<�}a<~a<;a<9�a<�a<�a<��a<�a<��a<��a<�a</�a<��a<P�a<��a<i�a<��a<��a<�a<q�a<��a<�a<�a<{�a<#�a<'�a<�a<�a<��a<��a<8�a<<�a<��a<i�a<��a<��a<�a<��a<u�a<a<��a<0�a<��a<��a<&�a<%�a<��a<��a<�a<[�a<{�a<�a<D�a<יa<ǚa<�a<�a<j�a<c�a<d�a<D�a<y�a<�a<��a<��a<�a<s�a<?�a<�a<��a<��a<c�a<��a<8�a<&�a<��a<��a<�a<\�a<˃a<��a<�}a<�{a<Jza<�ya<2za<p{a<f}a<�a<Ăa<ąa<��a<u�a<��a<D�a<5�a<��a<W�a<��a<��a<�a<��a<�a<�a<��a<^�a<��a<�a<�a<^�a<��a<��a<�a<0�a<��a<��a<�a<�|a<ya<ua<qa<ma<�ia<�fa<xda<ca<�ba<ca<Qda<Ifa<�ha<�ka<una<Pqa<�sa<�ua<Awa<xa<Txa<xa<qwa<Eva<ua<�sa<�ra<�qa<oqa<1qa<Qqa<�qa<bra<sa<�sa<�sa<�sa<Ksa<$ra<bpa<
na<@ka<�ga<yda<
aa<�]a<[a<�Xa<�Wa<Wa<�Wa<�Xa<
[a<�]a<aa<�da<�  �  �ha<�ka<�na<�pa<�ra<�sa<Yta<=ta<�sa</sa<�ra<�qa<�qa<iqa<xqa<*ra<sa<=ta<�ua<�va<Qxa<5ya<�ya<�ya<tya<2xa<�va<Wta<�qa<(oa<gla<ja</ha<�fa<�fa<�fa<Dha<dja<\ma<�pa<�ta<�xa<b|a<�a<�a<�a<�a<N�a<"�a<t�a<s�a<*�a<	�a<ǉa<މa<"�a<Ċa<ԋa<�a<��a<�a<��a<
�a<��a<��a<k�a<��a<,�a<Z�a<͍a<�a<9�a<?�a<ςa<��a<ga<�~a<=a<Y�a<U�a<�a<��a<r�a<��a<�a<�a<F�a<@�a<Z�a<�a<�a<��a<a<��a<#�a<`�a<�a<��a<�a<n�a<*�a<7�a<�a<*�a<Лa<5�a<�a<3�a<a<��a<+�a<�a<�a<��a<y�a<܅a<��a<`�a<Áa<)�a<<�a<=�a<��a<��a<�a<�a<�a<X�a<i�a<әa<��a<a<E�a<��a<h�a<m�a<J�a<l�a<˔a<X�a<��a<ݔa<{�a<E�a<�a<×a<�a<�a<c�a<D�a<O�a<�a< �a<��a<I�a<��a<��a<�~a<�|a<y{a<�za<]{a<�|a<�~a<րa<��a<��a<G�a<�a<��a<W�a<#�a<M�a<�a<�a<��a<�a<��a<�a<�a<؆a<+�a<�a<߅a<%�a<_�a<��a<͆a<��a<�a<��a<Âa<�a<5}a<�ya<�ua<ra<na<�ja<�ga<�ea<Dda<�ca<-da<lea<Uga<�ia<~la<oa<�qa<$ta<�ua<Swa<�wa<xa<uwa<�va<Sua<ta<�ra<�qa<�pa<$pa<pa<Cpa<�pa<rqa<	ra<�ra<Jsa<ysa<sa<ra<�pa<>na<�ka<~ha<Rea<ba<�^a<0\a<Za<�Xa<CXa<�Xa<�Ya<!\a<�^a<�aa<cea<�  �  �ia<�la<3oa<(qa<�ra<]sa<�sa<Zsa<�ra<�qa<�pa</pa<�oa<eoa<�oa<)pa<=qa<{ra<ta<�ua<*wa<exa<Mya<�ya<Dya<�xa<wa<ua<�ra<Ipa<�ma<�ka<�ia<�ha<�ha<�ha<=ja<Ula<�na<`ra<�ua<�ya<M}a<��a<��a<�a<��a<وa<l�a<s�a<A�a<Ԉa<E�a<�a<�a<)�a<шa<ىa<Q�a<֌a<��a<��a< �a<G�a<�a<+�a<��a<��a<Ԑa<��a<�a<i�a<�a<k�a<��a<e�a<�a<=�a<X�a<.�a<��a<��a<��a<ďa<Ȓa<s�a<��a<�a<	�a<p�a<'�a<��a<��a<��a<]�a<��a<�a<��a<�a<��a<k�a<��a<Ԙa<�a<�a<��a<��a<��a<��a<4�a<��a<�a<�a<�a<!�a<��a<��a<U�a<σa<!�a<9�a<��a<Z�a<�a<��a<�a<��a<�a<��a<��a<!�a<�a<b�a<a�a<0�a<ȕa<��a<��a<ƒa<s�a<��a<�a<��a<��a<��a<��a<5�a<v�a<�a<�a<��a<u�a<��a<��a<j�a<N�a<4�a<��a<�~a<u}a<�|a<U}a<v~a<�a<�a<��a<��a<2�a<`�a<J�a<S�a<�a<ُa<-�a<�a<y�a<a<�a<`�a<�a<ބa<8�a<�a<�a<[�a<��a<��a<a<҅a<j�a<Z�a<��a<��a<�}a<yza<�va<7sa<�oa<Zla<�ia<�ga<Ifa<�ea<+fa<Fga<�ha<Eka<�ma<.pa<�ra<�ta<Lva<'wa<�wa<uwa<�va<�ua<(ta<�ra<qa<�oa<�na<>na<na<bna<�na<�oa<�pa<�qa<Zra<�ra<�ra<�qa<�pa<�na<Cla<}ia<dfa<[ca<s`a<�]a<�[a<�Za<OZa<�Za<�[a<�]a<k`a<cca<xfa<�  �  ka<ima<�oa<Bqa<lra<�ra<�ra<-ra<&qa<&pa<�na<�ma<Cma<�la<7ma<�ma<�na<Ipa<ra<�sa<�ua<Dwa<Vxa<4ya<7ya<�xa<�wa<va<;ta<�qa<�oa<�ma<Xla<Tka<�ja<zka<�la<�na<3qa<jta<�wa<!{a<�~a<[�a<$�a<�a<s�a<�a<Z�a< �a<��a<��a<"�a<Ʌa<l�a<��a<d�a<\�a<�a<��a<֌a<��a<��a<7�a<8�a<�a<��a<�a<��a<׏a<��a<!�a<�a<��a<�a<̓a<j�a<��a<Äa<��a<��a<��a<5�a<?�a<͓a<�a<�a<	�a<��a<��a<�a<�a<͖a<�a</�a<C�a<k�a<Y�a<f�a<�a</�a<f�a<�a<S�a<��a<z�a<��a<ۚa<�a<��a<��a<l�a<��a<ߎa<:�a<։a<�a<��a<X�a<��a<��a<H�a<v�a<�a<��a<U�a<l�a<n�a<��a<��a<��a<�a<5�a<Ȗa<_�a<��a<N�a<!�a<A�a<�a<�a<��a<��a<��a<��a<�a<�a<�a<��a<�a<ؔa<�a<��a<"�a<�a<;�a<U�a<�a<(�a<�a<�a<�a<�a<X�a<��a<��a<!�a<p�a<�a<��a<W�a<��a<�a<�a<��a<��a<�a<Ća<�a<q�a<h�a<ˁa<v�a<ځa<<�a<�a<��a<i�a<a<��a<�a<��a<�a<c~a<�{a<_xa<�ta<�qa<�na<&la< ja<�ha<Kha<�ha<�ia<ka<;ma<Aoa<�qa<�sa<Hua<�va<wa<Gwa<�va<�ua<ta<_ra<�pa<�na<�ma<Pla<�ka<�ka<�ka<�la<�ma<�na<	pa<"qa<�qa<ra<�qa<�pa<Poa<ma<�ja<�ga<4ea<�ba<*`a<u^a<(]a<�\a<(]a<p^a<+`a<�ba<Gea<ha<�  �  Tla<�na<bpa<�qa<6ra<.ra<�qa<�pa<hoa<�ma<�la<Xka<zja< ja<ja<�ja<la<�ma<�oa<�qa<�sa<�ua<vwa<�xa<(ya<ya<xxa<$wa<�ua<�sa<
ra<apa<oa<*na<�ma<{na<�oa<~qa<�sa<�va<�ya<�|a<�a<d�a<��a<)�a<�a<P�a<B�a<��a<��a<��a<��a<�a<��a<��a<Z�a<��a<>�a<O�a<��a<Ȍa<�a<�a<h�a<��a<ғa<z�a<��a<�a<,�a<>�a<�a<M�a<Їa<a<k�a<��a<��a<I�a<R�a<��a<C�a<��a<�a<��a<I�a<�a<0�a<��a<Зa<U�a<ǔa<6�a<��a<q�a<��a<<�a<}�a<H�a<��a<�a<a<��a<2�a<{�a<;�a<��a<>�a<K�a<��a<��a<Y�a<��a<��a<��a<܊a<��a<[�a<��a<y�a<��a<�a<&�a<d�a<��a<��a<�a<�a<R�a<�a<�a<̖a<
�a<,�a<\�a<��a<W�a<`�a<��a<.�a<�a<��a<e�a<�a<^�a<Ŕa<��a<�a<��a<5�a<ܓa<̑a<��a<�a<`�a<�a<��a<��a<�a<��a<��a<��a<�a<Ća<߈a<Ɗa<��a<(�a<.�a<��a<W�a<P�a<�a<�a<ֈa<��a<a�a<X�a<��a<ka<�~a<�~a<a<�a<ʀa<Ɓa<тa<��a<a<��a<܂a<h�a<fa<�|a<�ya<wa<�sa<<qa<�na<�la<�ka<Ika<yka<ala<�ma<_oa<Oqa<sa<�ta<1va<�va< wa<�va<�ua<Uta<_ra<Zpa<Vna<ila<�ja<�ia<�ha<�ha<ia<	ja<Jka<�la<:na<�oa<�pa<Nqa<|qa<�pa<�oa<.na<la<�ia<Rga<�da<�ba<7aa<#`a<�_a<$`a<4aa<�ba<�da<iga<�ia<�  �  �ma<�oa<�pa<�qa<�qa<�qa<�pa<%oa<�ma<�ka<�ia<lha<hga<�fa<�fa<�ga<ia<�ja<#ma<�oa<ra<rta<�va<�wa<	ya<`ya<2ya<�xa<Fwa<va<]ta<sa<�qa<Cqa<+qa<�qa<�ra<Yta<�va<%ya<|a<�~a<8�a<q�a<�a<>�a<��a<��a<��a<߄a<��a<4�a<
�a<�a<�a<�a<D�a<��a<1�a<��a<�a<֊a<K�a<��a<��a<��a<ߓa<�a<��a<u�a<��a<r�a<��a<�a<��a<��a<��a<�a<Ǌa<�a<��a<�a<m�a<j�a<S�a<Ǘa<��a<�a<��a<ʗa<T�a<��a<��a<��a<�a<[�a<��a<�a<o�a<=�a<��a<c�a<f�a<��a<��a<X�a<��a<E�a<j�a<֙a<�a<6�a<X�a<B�a<+�a<O�a<Ѝa<��a<w�a<Ōa<{�a<Îa<}�a<m�a<v�a<1�a<̗a<��a<:�a<�a<I�a<�a<,�a<1�a<��a<��a<��a<E�a<U�a<ىa<+�a<͊a<#�a<ɍa<��a<��a<@�a<��a<s�a<וa<z�a<��a<)�a<-�a<$�a<��a<��a<��a<�a<�a<��a<�a<|�a<чa<E�a<�a<��a<�a<6�a<��a<��a<ێa<��a<��a<^�a<�a<"�a<��a<Qa<�}a<[|a<�{a<�{a<�{a<}a<A~a<�a<�a<=�a<�a<(�a<�a<сa<\�a<B~a<�{a<?ya<hva<�sa<�qa<)pa<�na<zna<�na<(oa<bpa<�qa<ysa<�ta< va<�va<@wa<wa<va<�ta<�ra<�pa<@na<�ka<�ia<�ga<�fa<�ea<�ea<fa<ga<�ha<]ja<`la<na<�oa<�pa<+qa<*qa<upa<eoa<�ma<�ka<�ia<{ga<�ea<*da<`ca<�ba<^ca<5da<�ea<�ga<�ia<�ka<�  �  �oa<�pa<�qa<ra<�qa<�pa<_oa<�ma<xka<aia<Uga<�ea<ada<�ca<�ca<�da<fa<%ha<�ja<ema<)pa<�ra<_ua<twa<�xa<�ya<�ya<�ya<�xa<�wa<�va<�ua<�ta<Jta<9ta<�ta<�ua<lwa<|ya<�{a<~a<m�a<��a<E�a<��a<?�a<F�a<ƅa<��a<!�a<��a<�a<X~a<5}a<z|a<w|a<}a<d~a<f�a<҂a<��a<��a<��a<H�a<��a<��a<֓a<v�a<F�a<ܓa<��a<n�a<�a<Ԏa<��a<��a<��a<�a<͍a<�a<��a<�a<M�a< �a<��a<y�a<�a<�a<�a<��a<ٔa<��a<n�a<�a<�a<x�a<`�a<�a<8�a<)�a<a<Ía<�a<��a<�a<�a<ݘa<�a<��a<x�a<Йa<a<)�a<w�a<ɓa<,�a<�a<��a<��a<͏a<��a<��a<�a<��a<L�a<ɗa<ɘa<^�a<r�a<ۘa<��a<ƕa<��a<�a<��a<�a<��a<=�a<�a<��a<�a<އa<_�a<=�a<q�a<��a<��a<��a<�a<��a<Օa<C�a<Y�a<ݒa< �a<�a<9�a<��a<�a<+�a<��a<�a<��a<��a<ߋa<*�a<n�a<��a<
�a<;�a<��a<��a<ǌa<O�a<��a<ńa<��a<�~a<�|a<za<-ya<�xa<}xa<4ya<Wza<�{a<�}a<Ha<Ҁa<�a<Âa<��a<d�a< �a<�a<�}a<;{a<�xa<�va<�ta<+sa<
ra<�qa<�qa<+ra<sa<3ta<Yua<�va<ewa<�wa<�wa<�va<�ua<�sa<`qa<�na<la<6ia<�fa<�da<Gca<�ba<fba<ca<Jda< fa<ha<?ja<^la<Dna<�oa<�pa<Sqa<qa<Spa</oa<�ma<�ka<ja<}ha<@ga<efa<fa<efa<Hga<�ha<-ja<�ka<�ma<�  �  �pa<�qa<Xra</ra<eqa<)pa<?na<?la<�ia<>ga<�da<�ba<�aa<�`a<�`a<�aa<Tca<nea<@ha<Ika<ina<�qa<Kta<�va<�xa<za<�za<�za<qza<�ya<ya<xa<�wa<wa<&wa<�wa<�xa<?za<�{a<~a<�a<�a<�a<�a<"�a<1�a<�a<Ԅa<g�a<��a<za<�}a<�{a<|za<�ya<wya<za<s{a<�}a<+�a<f�a<��a<��a<�a<ďa<7�a<��a<�a<�a<�a<b�a<k�a<h�a<?�a<��a<��a<��a<�a<��a<ӑa<�a<ʔa<1�a<��a<��a<B�a<_�a<��a<��a<��a<��a<��a<S�a<Ћa<f�a<��a<c�a<��a<?�a<Y�a<�a<9�a<�a<��a<��a<��a<�a<��a<��a<�a<��a<�a<ݘa<��a<�a<��a<��a<Ԓa<��a<��a<Y�a<F�a<w�a<ޖa<�a<,�a<��a<�a<��a<��a<�a<��a<E�a<6�a<u�a<��a<E�a<u�a<!�a<��a<�a<�a<��a<�a<U�a<׍a<~�a<q�a<a�a<g�a<�a<	�a<]�a<V�a<֒a<[�a<��a<5�a<�a<�a<ًa<��a<c�a<�a<&�a<,�a<�a<͐a<�a<��a<��a<'�a<Ջa<)�a<%�a<��a<�a<Z|a<�ya<�wa<-va<�ua<�ua<}va<�wa<�ya<�{a<�}a<�a<�a<e�a<��a<ւa<�a<Հa<+a<8}a<A{a<.ya<�wa<�ua<ua<�ta<hta<�ta<tua<~va<=wa<xa<xxa<xxa<xa<�va</ua<�ra<'pa<ma<�ia<�fa<da<	ba<J`a<�_a<m_a<1`a<�aa<vca<�ea<Hha<ka<$ma<#oa<�pa<jqa<�qa<9qa<�pa<9oa<�ma<kla<ka<ja<;ia<2ia<Bia<ja<&ka<�la<na<~oa<�  �  ra<�ra<�ra<Cra<Eqa<�oa<Xma<�ja<ha<Vea<�ba<�`a< _a<S^a<U^a<4_a<�`a<-ca<)fa<via<�la<\pa<|sa<kva<�xa<)za<?{a<�{a<�{a<Y{a<�za<.za<�ya<�ya<�ya<1za<{a<�|a<~a<�a<݁a<��a<��a<�a<k�a<<�a<��a<.�a<Z�a<)�a<�}a<�{a<�ya<xa<*wa<�va<�wa<ya<B{a<�}a<j�a<ڄa<{�a<��a<�a<ّa<��a<*�a<��a<�a<a</�a<V�a<`�a<Œa<;�a<#�a<g�a<�a<�a<6�a<��a<�a<�a<��a<�a<��a<��a<*�a<ޔa<X�a<s�a<��a<Éa<*�a<J�a<��a<s�a<ǃa<�a<��a<�a<�a<��a<�a<�a<��a<v�a<��a<y�a<��a<<�a<m�a<^�a<'�a<�a<�a<W�a<�a<0�a<��a<}�a<��a<��a<��a<V�a<a<��a<��a<`�a<i�a<��a<֐a<��a<��a<��a<��a<��a<��a<0�a<��a<��a<f�a<͆a<��a<P�a<'�a<��a<�a<Z�a<B�a<��a<g�a<��a<z�a</�a<��a<u�a<e�a<��a<;�a<8�a<��a<=�a<"�a<�a<��a<�a<͑a<�a<��a<ڍa</�a<�a<��a<
�a<�}a</za<jwa<0ua<�sa<sa<&sa<ta<}ua<�wa<�ya<<|a<�~a<l�a<�a<��a<�a<ӂa<�a<��a<�~a</}a<N{a<�ya<mxa<�wa<�va<�va<,wa<�wa<Uxa<�xa<Yya<�ya<(ya<3xa<�va<�ta<�qa<�na<ka<ha<�da<�aa<�_a<�]a<�\a<�\a<�]a<?_a<Vaa<�ca<�fa<�ia<2la<�na<\pa<yqa<ra<4ra<�qa<�pa<�oa<tna<Ama<gla<�ka<�ka<�ka<wla<\ma<�na<�oa<qa<�  �  �ra<esa<$sa<wra<qa<oa<�la<�ia<�fa<�ca<!aa<�^a<"]a<[\a<K\a<@]a<�^a<�aa<�da<"ha<�ka<_oa<�ra<�ua<xxa<fza<�{a<u|a<�|a<�|a<|a<�{a<�{a<u{a<�{a<|a<}a<T~a<�a<w�a<�a<��a<��a<��a<��a<d�a<3�a<��a<��a<a<�|a<za<�wa<9va<,ua<�ta<�ua<wa<\ya<\|a<�a<��a<r�a<'�a<��a<]�a<ғa<m�a<v�a<Ԗa<Ӗa<Z�a<��a<+�a<��a<9�a<�a<b�a<�a<ϕa<��a<�a<�a<�a<o�a<d�a<ϙa<��a<��a<\�a<g�a<c�a<C�a<�a<��a<X�a<�a<q�a<́a<�a<�a<{�a<~�a<ލa<	�a<A�a<��a</�a<�a<כa<V�a<�a<��a<��a<��a<��a<�a<Z�a<��a<6�a<��a<B�a<$�a<�a<Кa<3�a<j�a<��a<�a<+�a<Օa<�a<Џa<��a<�a<�a<0�a<��a<�a<%a<�a<��a<��a<#�a<,�a<=�a<*�a<�a<P�a<D�a<~�a<�a<�a<��a<��a<q�a<k�a<0�a<I�a<��a<$�a<8�a<x�a<�a<��a<�a<��a<��a<X�a<T�a<ӏa<n�a<��a<V�a<��a<�a<�{a<�xa<�ua<1sa<�qa<�pa<&qa<*ra<�sa<va<�xa<3{a<�}a<�a<��a<܂a<Z�a<O�a<��a<��a<&�a<�~a<}a<�{a<kza<rya<�xa<�xa<�xa<Yya<�ya<$za<Wza<<za<�ya<sxa<�va<#ta<eqa<�ma<pja<�fa<;ca<?`a<�]a<�[a<�Za<�Za<�[a<r]a<�_a<vba<�ea<�ha<�ka<na<pa<�qa<ura<�ra<zra<�qa<�pa<pa<oa<=na<�ma<qma<�ma<Rna<!oa<0pa< qa<Ira<�  �  �sa<�sa<bsa<vra<�pa<�na<Bla<<ia<	fa<�ba<`a<�]a<\a<,[a<[a<\a<�]a<f`a<}ca<)ga<�ja<�na<�ra<�ua<Zxa<rza<�{a<�|a<Y}a<j}a<}a<�|a<z|a<�|a<�|a<^}a<2~a<ea<րa<r�a<��a<o�a<N�a<��a<ۆa<P�a<�a<Q�a<
�a<k~a<�{a<ya<�va<ua<ta<�sa<qta<�ua<Dxa<K{a<�~a<��a<��a<��a<5�a<-�a<a<��a<Ŗa<]�a<��a<A�a<��a<%�a<��a<J�a<L�a<��a<�a<̖a<�a<�a<��a<��a<ޚa<��a<ߙa<�a<n�a<�a<ߐa<��a<G�a<�a<n�a<B�a<׀a<A�a<��a<ˁa<΃a<q�a<��a<�a<t�a<ȓa<��a<	�a<�a<�a<��a<��a<b�a<��a<��a<��a<��a<o�a<J�a<J�a<��a<<�a<�a<ܚa<��a<ޛa<��a<�a<�a<�a<��a<��a<B�a<��a<$�a<ބa<�a<�a<�~a<�}a<d~a<�a<��a< �a<3�a<h�a<��a<��a<"�a<%�a<��a<S�a<|�a<>�a<��a<m�a<X�a<*�a<U�a<��a<h�a<M�a<��a<��a<��a<�a<q�a<5�a<��a<x�a<��a<?�a<S�a<͆a<�a<�~a<	{a<�wa<tta<ra<�pa<�oa<pa<qa<�ra<ua<�wa<qza<#}a<�a<[�a<˂a<v�a<��a<)�a<g�a<�a<�a<~a<�|a<{{a<�za<za<�ya<�ya<Eza<�za<{a<{a<�za<�ya<�xa<�va<�sa<�pa<gma<�ia<�ea<5ba<$_a<�\a<�Za<�Ya<�Ya<�Za<W\a<�^a<�aa<�da<�ga<ka<�ma<�oa<�qa<�ra<&sa<sa<�ra<�qa<�pa<�oa<Poa<�na<�na<�na<aoa<pa<*qa<ra<sa<�  �  �sa<�sa<�sa<�ra<�qa<pa<na<la<�ia<nga<2ea<�ca<Uba<�aa<�aa<}ba<da<fa<�ha<ska<3na<gqa< ta<�va<�xa<�za<�{a<�|a<c}a<j}a<�}a<M}a<d}a<�}a<�}a<o~a<Fa<U�a<Q�a<Ԃa<�a<:�a<�a<��a<߆a<m�a<��a<J�a<Ȃa<�a<a<V}a<�{a<�za<�ya<�ya<}za<�{a<�}a<	�a<�a<�a<�a<6�a<�a<��a<z�a<)�a<�a<��a<��a<͖a<��a<�a<��a<�a<ӕa<�a<��a<6�a<ۗa<�a<v�a<'�a<E�a<�a<��a<k�a<�a<ٔa<Ӓa<-�a<�a<��a<m�a<�a<��a<m�a<��a<��a<'�a<�a<��a<��a<��a<�a<\�a<N�a<Ěa<Ûa<�a<I�a<�a<o�a<��a<��a<��a<�a<��a<��a<b�a<��a<!�a<ۚa<(�a<}�a<=�a<Ϛa<ƙa<<�a<D�a<ݓa<~�a<��a<�a<p�a<h�a<��a<��a<4�a<M�a<U�a<ņa<��a<��a<!�a<��a<��a<��a<4�a<g�a<ޖa<��a<Жa<�a<w�a<\�a<��a<	�a<M�a<�a<�a<
�a<�a<��a<��a<ܒa<��a<�a<-�a<��a<��a<�a<Y�a<W�a</�a<-a<?|a<�ya<�wa<�va<�ua<�ua<�va<�wa<lya<D{a<$}a<a<��a<�a<�a<��a<^�a<��a<;�a<�a<�a<�~a<�}a<�|a<�{a<1{a<{a<�za<�za<-{a<{a<{a<�za<�ya<�xa<wa<ua<nra<�oa<�la<ja<6ga<�da<�ba<-aa<�`a<X`a<�`a<Cba<�ca<fa<Bha<�ja<�la<oa<�pa<ra<�ra<8sa<Osa<�ra<\ra<�qa<�pa<�pa<pa<pa<'pa<�pa<qa<�qa<�ra<6sa<�  �  ysa<�sa<|sa<�ra<�qa<Epa<Pna<*la<�ia<�ga<pea<�ca<�ba<�aa<ba<�ba<:da<Cfa<�ha<�ka<tna<�qa<Zta<�va<�xa<�za<�{a<�|a<}a<K}a<P}a<D}a<8}a<F}a<�}a<'~a<�~a<�a<R�a<��a<ރa<�a<�a<��a<��a<e�a<��a<~�a<��a<1�a<Va<�}a<�{a<�za<2za< za<�za<|a<�}a<W�a<!�a<1�a<J�a<Z�a<"�a<��a<��a<�a<�a<��a<��a<��a<j�a<�a<a<��a<��a<ѕa<N�a<�a<ٗa<��a<X�a<�a<-�a<�a<��a<r�a<�a<,�a<��a<q�a<�a<��a<��a<�a<�a<��a<�a<ԇa<R�a<M�a<��a<D�a<�a<W�a<��a<V�a<��a<��a<�a<��a<��a<6�a<��a<�a<F�a<טa<��a<��a<��a<~�a<�a<��a<��a<.�a<%�a<��a<��a<G�a<z�a<*�a<��a<ݎa<B�a<��a<��a<�a<Մa<\�a<��a<�a<��a<шa< �a<b�a<܏a<�a<�a<;�a<@�a<Жa<ޖa<��a<�a<.�a<S�a<q�a<��a<�a<��a<��a<ɑa<�a<a�a<��a<��a<x�a<�a< �a<��a<��a<E�a<��a<��a<n�a<ca<�|a<za<;xa<�va<?va<Hva<�va<xa<�ya<s{a<X}a<9a<րa<-�a<�a<`�a<_�a<ւa<�a<�a<�a<�~a<W}a<F|a<y{a<�za<�za<�za<�za<�za<�za<�za<�za<�ya<�xa<wa<5ua<�ra<pa<
ma<5ja<\ga<�da<�ba<�aa<�`a<�`a<@aa<nba<da<Ifa<�ha<�ja<1ma<=oa<�pa< ra<�ra<$sa<sa<�ra<#ra<�qa<�pa<9pa<�oa<�oa<�oa<Npa<�pa<�qa<mra<sa<�  �  
sa<�sa<Msa<�ra<�qa<Zpa<�na<~la<qja<<ha<Pfa<�da<�ca<ca<�ba<�ca<ea<+ga<�ia<:la<oa<�qa<�ta<�va<ya<�za<�{a<o|a<�|a<�|a<}|a<|a<N|a<I|a<�|a<1}a<~a<a<��a<Ɂa<B�a<��a<��a<_�a<��a<��a<��a<��a<I�a<��a<�a<7~a<�|a<�{a<5{a<	{a<�{a<}a<�~a<@�a<փa<Άa<ωa<��a<Z�a<��a<��a<�a<ؕa<9�a<H�a<�a<��a<D�a<Ȕa<��a<��a<�a<V�a<�a<�a<ėa<�a<g�a<�a<�a<t�a<��a<'�a<`�a<:�a<�a<��a<w�a<��a<�a<�a<z�a<�a<ǈa<-�a<.�a<`�a<�a<A�a<��a<��a<j�a<a<k�a<ۛa<��a<Q�a<��a<ƙa<�a<L�a<�a<��a<ۗa<��a<��a<D�a<ҙa<��a<��a<�a<w�a<��a<^�a<��a<n�a<��a<��a<�a<��a<p�a<ֆa<ۅa<9�a<��a<^�a<�a<��a<ŋa<�a<#�a<:�a<��a<]�a<:�a<��a<��a<�a<��a<[�a<��a<��a<��a<5�a<Ȑa<a<͐a<<�a<��a<�a<6�a<�a<Бa<ِa<��a<��a<}�a<وa<��a<�a<�a<r}a<�za<>ya<�wa<#wa<Qwa<�wa<�xa<Qza<|a<�}a<�a<�a<6�a<�a<>�a<&�a<�a<��a<e�a<�~a<�}a<]|a<^{a<�za<za<�ya<�ya<za<za<{za<^za<=za<�ya<�xa<<wa<?ua<�ra<Opa<�ma<�ja<(ha<�ea<�ca<�ba<�aa<�aa<3ba<Ica< ea<�fa<1ia<Qka<yma<]oa<�pa<ra<�ra<�ra<�ra<Gra<lqa<�pa<�oa<?oa<oa<�na<oa<Ooa<pa<�pa<�qa<�ra<�  �  gra<�ra<�ra<�ra<�qa<�pa<1oa<Xma<Nka<Iia<zga<�ea<�da<dda<xda<7ea<|fa<fha<�ja<9ma<�oa<�ra<ua<Hwa<ya<�za<9{a<�{a<�{a<�{a<�{a<E{a<{a<{a<D{a<�{a<�|a<�}a<Da<ǀa<I�a<��a<�a<̅a<S�a<p�a<�a<-�a<�a<x�a<�a<[a<~a<}a<||a<�|a<.}a<^~a<�a<b�a<��a<Ça<��a<a�a<ُa<ܑa<��a<��a<F�a<��a<o�a<�a<��a<	�a<�a<N�a<1�a<}�a<�a<ɔa<Օa<֖a<ܗa<��a<N�a<a�a<U�a<��a<r�a<�a<�a<�a<��a<��a<ˋa<N�a<l�a<�a<K�a<�a<}�a<T�a<v�a<Ƒa<�a<A�a<�a<��a<��a<�a<E�a<��a<[�a<��a<��a<Зa<�a<��a<J�a<l�a<��a<b�a<�a<ߘa<��a<�a<^�a<�a<��a<v�a<�a<�a<Ӓa<c�a<��a<��a<��a<'�a<;�a<Άa<�a<a<�a<ъa<Ōa<ގa<��a<ǒa<H�a<j�a<�a<"�a<�a<T�a<~�a<k�a<T�a<?�a<c�a<a<^�a<h�a<��a<��a<��a<��a<S�a<�a<<�a<��a<��a<�a<�a<��a<Άa<��a<1�a<�~a<R|a<�za<Nya<�xa<�xa<ya<za<v{a<}a<�~a<@�a<��a<l�a<�a<�a<��a<�a<��a<ga<�}a<|a<{a<za<ya<�xa<lxa<nxa<�xa<ya<uya<�ya<�ya<#ya<�xa<Bwa<�ua<~sa<qa<zna<�ka<Pia<ga<*ea<�ca<%ca<ca<�ca<�da<%fa<ha<ja<-la<na<�oa<qa<ra<Lra<ara<�qa<Rqa<upa<�oa<�na<�ma<�ma<ama<�ma<na<�na<�oa<�pa<�qa<�  �  �qa<Hra<�ra<�ra<ra<9qa<�oa<[na<tla<�ja<ia<�ga<�fa<3fa<qfa<�fa<nha<ja<7la<�na<qa<�sa<�ua<�wa<ya<Xza<�za<4{a<
{a<�za<+za<�ya<Vya<(ya<bya< za<�za<|a<�}a<8a<��a<��a<?�a<E�a<!�a<]�a<B�a<��a<��a<��a<%�a<�a<�a<�~a<N~a<y~a< a<'�a<	�a<
�a<��a<�a<��a<1�a<^�a<>�a<��a<��a<͔a<�a<n�a<ēa<�a<V�a<Ǒa<b�a<f�a<��a<+�a<�a<&�a<l�a<��a<��a<��a< �a<)�a<��a<ߗa<~�a<�a<��a<�a<)�a<{�a<B�a</�a<�a<'�a<��a<T�a<�a<��a<�a<(�a<��a<��a<��a<��a<ښa<��a<,�a<7�a<9�a<�a<�a<A�a<��a<��a<��a<�a<��a<�a<��a<i�a<I�a<��a<Йa<~�a<��a<o�a<��a<Փa<��a<n�a<D�a<��a<�a<
�a<Ȉa<̈a<��a<ъa<[�a<.�a<��a<�a<e�a<��a<l�a<��a<˕a<a�a<w�a<B�a<	�a<��a<��a<��a<�a<��a<z�a<ɍa<H�a<�a<��a<F�a<ːa<��a<o�a<��a<;�a<x�a<K�a<�a<<�a<a<7�a<3~a<W|a<<{a<�za<aza< {a<�{a<}a<S~a<�a<�a<�a<ςa<��a<�a<�a<7�a<�a<~a<l|a<�za<]ya<xa<Rwa<�va<�va<�va<wa<�wa<2xa<�xa<�xa<�xa<Xxa<6wa<�ua<ta<�qa<�oa<1ma<�ja<�ha<ga<�ea<ea<�da<eea<ofa<�ga<�ia<>ka<8ma<�na<Hpa<8qa<�qa<ra<�qa<3qa<.pa<'oa<�ma<ma<5la<�ka<�ka<�ka<Bla<"ma<$na<boa<xpa<�  �  fpa<xqa<6ra<�ra<Gra<�qa<�pa<joa<�ma<Yla<�ja<�ia<�ha<qha<�ha<?ia<wja<la<�ma<.pa<nra<�ta<uva<xa<Nya<'za<bza<Cza<�ya<Mya<rxa<�wa<_wa<wa<Cwa<�wa<�xa<za<�{a<m}a<�a<h�a<�a<��a<ƅa<h�a<��a<C�a<��a<̈́a<��a<��a<��a<Հa<��a<��a<?�a<j�a<��a<�a<3�a<��a<�a<3�a<��a<��a<��a<-�a<0�a<Փa<1�a<g�a<F�a<s�a<��a<<�a<3�a<�a<�a<"�a<T�a<��a<E�a<��a<��a<y�a<�a<��a</�a<,�a<�a<U�a<��a<�a<k�a<@�a<s�a<,�a<\�a< �a<B�a<��a<��a<^�a<C�a<՗a<�a<��a<x�a<n�a<��a<�a<��a<��a<F�a<,�a<0�a<��a<B�a<^�a<ݒa<��a<��a<�a<*�a<�a<�a<`�a<`�a<Әa<��a<��a<�a<��a<�a<�a<w�a<0�a<I�a<��a<�a<��a<��a<�a<��a<^�a<�a<�a<�a<��a<Ǖa<K�a<q�a<@�a<��a<P�a<�a<��a<k�a<��a<Y�a<Q�a<��a<b�a<&�a<=�a<
�a<��a<�a<�a<��a<}�a<
�a<G�a<"�a<��a<^�a<�a<#�a<�~a<a}a<�|a<�|a<�|a<�}a<�~a<�a<�a<�a<��a<�a<	�a<��a<�a<�a<w~a<�|a<�za<�xa<Pwa<�ua< ua<�ta<kta<�ta<Dua<�ua<�va<{wa<�wa<;xa<xa<_wa<Fva<�ta<sa<�pa<�na<�la<�ja<ia<�ga<Dga<ga<�ga<]ha<�ia<ka<�la<Sna<�oa<�pa<vqa<�qa<�qa<�pa<	pa<�na<�ma<0la<ka<%ja<�ia<Zia<�ia<0ja<1ka<Zla<�ma<9oa<�  �  7oa<�pa<�qa<Ira<tra<-ra<�qa<wpa<Xoa<na<�la<�ka<ka<�ja<�ja<�ka<�la</na<�oa<�qa<�sa<�ua<Pwa<�xa<kya<�ya<�ya<iya<�xa<�wa<�va<�ua<!ua<�ta<�ta<Tua<lva<�wa<�ya<�{a<�}a<�a<�a<��a<G�a<R�a<Ɔa<�a<��a<�a<6�a<V�a<��a<��a<҂a<��a<��a<��a<�a<�a<�a</�a<*�a<�a<��a<͒a<��a<��a<��a<ےa<Ցa<��a<��a<|�a<t�a<��a<a<�a<̍a<܎a<k�a<�a<��a<7�a<��a<ܗa<��a<֘a<��a<�a<�a<��a<@�a<ϒa<��a<c�a<ҏa<w�a<ďa<[�a<d�a<ْa<E�a<�a<W�a<��a<��a<0�a<N�a<�a<$�a<��a<��a<�a<u�a<�a<��a<5�a<Ώa<�a<��a<��a<ݒa<0�a<��a<�a<$�a<Θa<&�a< �a<c�a<p�a<�a<o�a<��a<&�a<��a<e�a<��a<9�a<m�a<�a<�a<�a<a�a<��a<�a<��a<��a<��a<i�a<��a<��a< �a<g�a<��a<��a<Z�a<*�a<c�a<�a<�a<p�a<d�a<a�a<��a<��a<��a<`�a<��a<x�a<��a<��a<.�a<>�a<M�a<,�a<;�a<H�a<ڀa<�a<a<�~a<a<�a<��a<r�a<8�a<��a<o�a<^�a<�a<�a<ۀa<"a<}a<{a<�xa<�va<
ua<�sa<�ra<:ra<,ra<�ra<[sa<5ta<Gua<-va<wa<�wa<�wa<vwa<�va<�ua<ta<=ra<apa<na<�la<=ka<Ija<�ia<�ia<�ia<ja<�ka<�la<5na<goa<�pa<Mqa<�qa<�qa<qa<Apa<�na<yma<�ka<`ja<�ha<�ga<9ga<�fa<@ga<�ga<
ia<�ja<la<�ma<�  �  -na<�oa<(qa<"ra<�ra<�ra<`ra<�qa<�pa<�oa<�na<�ma<\ma<'ma<Rma<�ma<�na<Cpa<�qa<�sa<@ua<�va<xa<ya<�ya<�ya<7ya<�xa<}wa<,va<�ta<�sa<�ra<�ra<|ra<sa<ta<�ua<�wa<�ya<5|a<�~a<!�a<�a<�a<>�a<6�a<��a<��a<=�a<҆a<�a<��a<B�a<�a<i�a<	�a<��a<f�a<�a<ǋa<ҍa<��a<�a<]�a<?�a<��a<f�a<Ēa<�a<��a<�a<��a<X�a<P�a<��a<m�a<��a<��a<��a<F�a<)�a<�a<�a<ٕa<9�a<B�a<�a<�a<��a<��a<�a<�a<��a<��a<��a<�a<�a<�a<��a<��a<��a<�a<t�a<��a<��a<=�a<��a<.�a<q�a<E�a<ۖa<�a<H�a<x�a<�a<��a<؍a<��a<��a<_�a<j�a<Րa<��a<5�a<��a<<�a<R�a<��a<B�a<��a<;�a<&�a<�a<r�a<�a<Ƒa<��a< �a<��a<��a<5�a<��a<�a<�a<1�a<�a<��a<�a<�a<0�a< �a<��a<�a<Վa<ڌa<��a<7�a<�a<��a<��a<��a<L�a<@�a<z�a<�a<_�a<��a<��a<4�a<d�a<.�a<W�a<�a<��a<�a<�a<(�a<��a<�a<,�a<��a<2�a<]�a<��a<B�a<�a<��a<�a<�a<Ѓa< �a<āa<�a<0~a<�{a<gya<wa<�ta<�ra<fqa<Ypa<�oa<�oa<\pa<6qa<kra<�sa<ua<2va<�va<pwa<�wa<-wa<?va<ua<�sa<ra<Fpa<�na<�ma<�la<�ka<�ka<	la<�la<�ma<�na<�oa<�pa<nqa<�qa<ra<�qa<�pa<coa<�ma<la<7ja<dha<�fa<�ea<�da<�da<�da<�ea<�fa<|ha<]ja<Ela<�  �  "ma< oa<�pa<�qa<�ra<5sa<6sa<�ra<ra<hqa<�pa<�oa<ooa<Foa<�oa<pa<�pa<,ra<�sa<ua<~va<�wa<�xa<uya<�ya<Pya<�xa<�wa<[va<�ta<esa<�qa<qa<bpa<Mpa<�pa<�qa<�sa<�ua<xa<�za<m}a<�a<t�a<��a<�a<y�a<�a<��a<z�a<&�a<чa<l�a<>�a<1�a<��a<6�a<�a<l�a<�a<��a<)�a<a<*�a<�a<��a<x�a<!�a<$�a<�a<W�a<��a<�a<o�a<\�a<e�a<M�a<��a<Q�a<Ȋa<i�a<��a<��a<�a<�a<��a<�a<�a<t�a<d�a<�a<K�a<e�a<d�a<{�a<��a<:�a<+�a<<�a<��a<��a<��a<��a<��a<Ǚa<{�a<��a<��a<��a<�a<��a<ԕa<��a<��a<��a<��a<��a<��a<]�a<i�a<D�a<}�a<�a<�a<̒a<Քa<p�a<�a<Øa<e�a<j�a<�a<W�a<5�a<�a<̔a<��a<Œa< �a<��a<ܑa<D�a<�a<��a<��a<o�a<1�a<u�a<v�a<�a<�a<��a<Ǒa<ʏa<i�a<D�a<�a<J�a<��a<˄a<y�a<s�a<R�a<Q�a<Ǉa<c�a<�a<��a<�a<�a<D�a<q�a<��a<!�a<όa<=�a<��a<��a<��a<:�a<T�a<��a<U�a<d�a<��a<�a<l�a<фa<	�a<��a<"�a<�a<�a<sa<,}a<�za<�wa<cua<�ra<�pa<#oa<:na<�ma<�ma<mna<Yoa<�pa<=ra<�sa<<ua<mva<1wa<�wa<�wa<�va<1va<�ta<�sa<ra<�pa<�oa<�na<Bna<�ma<!na<�na<Uoa<?pa<	qa<�qa<Ura<cra<-ra<Nqa<Fpa<�na<�la<�ja<�ha<�fa<�da<�ca<�ba<wba<�ba<�ca<�da<�fa<�ha<�ja<�  �  %la<Zna<?pa<�qa<sa<~sa<�sa<�sa<Ssa<�ra<,ra<�qa<=qa<1qa<[qa<�qa<�ra<�sa<ua<ava<�wa<�xa<aya<�ya<�ya<ya</xa<�va<Kua<�sa<�qa<apa<6oa<�na<mna<�na<pa<�qa<�sa<�va<Tya<R|a<<a<�a<3�a<,�a<��a<��a<;�a<e�a<p�a<C�a<�a<�a<�a<g�a<�a<�a<!�a<��a<
�a<|�a<��a<גa<d�a<��a<��a<��a<��a<�a<=�a<I�a<o�a<ňa<q�a<��a<Y�a<��a<y�a<�a<ϊa<�a<i�a<ԑa<!�a<(�a<��a<�a<��a<�a<יa<]�a<��a<��a<0�a<�a<*�a<�a<#�a<��a<E�a<+�a<�a<��a<��a<"�a<�a<ךa<�a<��a<�a<ޔa<��a<L�a<&�a<@�a<��a<Ήa<d�a<��a<W�a<��a<z�a<{�a<��a<דa<˕a<h�a<��a<��a<��a<��a<+�a<k�a<p�a<l�a<q�a<��a<�a<��a<͓a<�a<��a<F�a<�a<��a<��a<�a<��a<�a<��a<�a<�a<��a<6�a<��a<p�a<p�a<��a<�a<��a<��a<b�a<��a<;�a<�a<�a<ǋa<W�a<��a<Q�a<��a<G�a<ʎa<��a<��a<�a<��a<;�a<�a<*�a<��a<?�a<�a<O�a<��a<��a<ʅa<��a<�a<S�a<��a<�a<�~a<W|a<�ya<�va<�sa<<qa<oa<\ma<Fla<�ka<�ka<�la<�ma<Coa<qa<�ra<zta<�ua<�va<�wa<�wa<�wa<�va<�ua<�ta<�sa<qra<Xqa<�pa<pa<�oa<�oa<^pa<�pa<�qa<Bra<�ra<�ra<�ra<Vra<Eqa<�oa<na<�ka<�ia<=ga<ea</ca<�aa<�`a<~`a<�`a<�aa<0ca<"ea<Uga<�ia<�  �  Lka<�ma<�oa<�qa<sa<�sa<sta<Yta<Pta<�sa<Vsa<�ra<�ra<�ra<�ra<bsa<ta<$ua<6va<Xwa<�xa<?ya<�ya<�ya<�ya<�xa<�wa<=va<qta<�ra<�pa<;oa<�ma<5ma<�la<[ma<�na<Cpa<�ra<\ua<Yxa<|{a<r~a<_�a<�a<)�a<ɇa<
�a<щa<-�a<s�a<1�a<Y�a<;�a<b�a<ڊa<w�a<V�a<n�a<Ԏa<��a<|�a<��a<o�a<�a<�a<��a<|�a<�a<R�a<h�a<P�a<J�a<��a<�a<U�a<̈́a<#�a<2�a<��a<��a<��a<~�a< �a<z�a<��a<��a<�a<�a<��a<r�a<E�a<��a<��a<p�a<ȗa<��a<U�a<��a<ԗa<��a<`�a<�a<��a<T�a<��a<��a<�a<ۙa<@�a<U�a<
�a<��a<F�a<��a<�a<V�a<w�a<͇a<B�a<�a<o�a<O�a<o�a<̐a<��a<1�a<
�a<��a<��a<�a<N�a<ԙa<g�a<`�a<��a<��a<וa<|�a<�a<7�a<P�a<ߕa<]�a<�a<}�a<��a<��a<��a<#�a<��a<��a<l�a<ߍa<U�a<��a<J�a<�a<��a<z�a<�a<^�a<��a<x�a<�a<�a<�a<��a<͌a<7�a<N�a<��a<Џa<a�a<��a<��a<�a<�a<��a<j�a<��a<��a<��a<e�a<��a<y�a<��a<��a<O�a<��a<{�a<�a<ڀa<k~a<�{a<�xa<�ua<�ra<pa<�ma<la<�ja<Fja<�ja<2ka<�la<!na<pa<�qa<�sa<uua<�va<�wa<�wa<xa<�wa<�va<�ua<�ta<�sa<�ra<�qa<kqa<Rqa<=qa<�qa</ra<�ra<Fsa<dsa<�sa<+sa<ora<5qa<yoa<sma<ka<�ha<7fa<�ca<�aa<N`a<}_a<�^a<w_a<W`a<�aa<�ca<Ifa<�ha<�  �  �ja<~ma<�oa<�qa<sa<ta<�ta<�ta<�ta<xta<ta<�sa<sa<zsa<�sa<8ta<�ta<�ua<wa<
xa<�xa<�ya<#za<$za<�ya<�xa<�wa<�ua<ta<ra<!pa<[na<ma<@la<la<~la<�ma<moa<�qa<�ta<�wa<�za<.~a<*�a<�a<�a<އa<@�a<�a<��a<�a<�a<#�a<-�a<U�a<��a<^�a<A�a<d�a<��a<ސa<��a<�a<ēa<,�a<�a<l�a<s�a<�a<�a<ތa<��a<��a<��a<2�a<J�a<�a<7�a<3�a<��a<ňa<:�a<ߍa<��a<'�a<��a<��a<��a<�a<��a<՚a<��a<P�a<ڙa<E�a<Øa<g�a<O�a<p�a<Әa<q�a<&�a<њa<i�a<̛a<��a<��a<�a<��a<3�a<�a<��a<�a<��a<"�a<�a<t�a<h�a<�a<8�a<�a<��a<p�a<ȍa<#�a<��a<�a<��a<z�a<��a<K�a<��a<G�a<ҙa<&�a<_�a<��a<֖a<U�a<�a<�a<H�a<��a<4�a<��a<�a<��a<Зa<&�a<�a<��a<��a<�a<�a<��a< �a<i�a<A�a<��a<��a<�a<R�a<!�a<��a<M�a<l�a<��a<��a<��a</�a<(�a<֏a<�a<��a<��a<�a<�a<��a<|�a<^�a<�a<܇a<{�a<\�a<Y�a<Z�a<A�a<�a<��a<�a<��a<�a<рa<3~a<O{a<&xa<ua<�qa<,oa<�la<	ka<�ia<Zia<�ia<Xja<�ka<{ma<xoa<�qa<�sa<Bua<�va<�wa<&xa<Fxa<�wa<Mwa<pva<�ua<�ta<�sa<�ra<era<-ra<<ra<�ra<�ra<[sa<�sa<�sa<�sa<\sa<qra<qa<loa<8ma<�ja<ha<�ea<ca<aa<k_a<o^a<
^a<m^a<n_a<aa<ca<�ea<4ha<�  �  �ja<0ma<�oa<�qa<-sa<8ta<�ta<ua<�ta<�ta<0ta<�sa<�sa<�sa<	ta<zta<Oua<va<)wa<>xa<%ya<�ya<4za<Oza<�ya<�xa<gwa<�ua<�sa<�qa<�oa<na<�la<�ka<�ka<Hla<Rma<Loa<�qa<ota<�wa<�za<~a<߀a<��a<��a<�a<B�a<6�a<�a<�a<Y�a<"�a<_�a<��a<��a<��a<��a<��a<��a<�a<)�a<A�a<ߓa<+�a<,�a<a�a<T�a<��a<�a<��a<��a<b�a<k�a<�a<�a<��a<�a<�a<��a<x�a< �a<��a<c�a<�a<M�a<w�a<�a<@�a<��a<	�a<�a<��a< �a<H�a<
�a<��a<��a<��a<9�a<��a<2�a<�a<��a<�a<�a<ƛa<�a<��a<��a<��a<��a<Ԑa<��a<�a<�a<F�a<�a<Ɇa<�a<ۇa<b�a<7�a<��a<��a<��a<��a<ǖa<q�a<��a<n�a<��a<��a<��a<o�a<q�a<��a<>�a<��a<c�a<O�a<��a<ǖa<Q�a<Ηa<�a<>�a<��a<R�a<�a<{�a<R�a<ۏa<N�a<f�a<Ǉa<�a<�a<X�a<8�a<�a<�a< �a<E�a<&�a<H�a<G�a<��a<N�a<�a<�a< �a<�a<ŏa<>�a<&�a<.�a<��a<��a<��a<��a<!�a<؇a<��a<R�a<��a<l�a<P�a<��a<�a<��a<ւa<��a<�}a<*{a<�wa<�ta<�qa<�na<�la<�ja<�ia<ia<Dia<6ja<hka<Ama<0oa<Yqa<Jsa<ua<�va<�wa<Uxa<Qxa<xa<}wa<�va<�ua<�ta<�sa<!sa<�ra<hra<�ra<�ra<sa<�sa<�sa<(ta<�sa<psa<�ra<qa<8oa<�la<�ja<�ga<qea<�ba<�`a<>_a<^a<�]a<^a<1_a<�`a<�ba<�ea<�ga<�  �  �ja<~ma<�oa<�qa<sa<ta<�ta<�ta<�ta<xta<ta<�sa<sa<zsa<�sa<8ta<�ta<�ua<wa<
xa<�xa<�ya<#za<$za<�ya<�xa<�wa<�ua<ta<ra<!pa<[na<ma<@la<la<~la<�ma<moa<�qa<�ta<�wa<�za<.~a<*�a<�a<�a<އa<@�a<�a<��a<�a<�a<#�a<-�a<U�a<��a<^�a<A�a<d�a<��a<ސa<��a<�a<ēa<,�a<�a<l�a<s�a<�a<�a<ތa<��a<��a<��a<2�a<J�a<�a<7�a<3�a<��a<ňa<:�a<ߍa<��a<'�a<��a<��a<��a<�a<��a<՚a<��a<P�a<ڙa<E�a<Øa<g�a<O�a<p�a<Әa<q�a<&�a<њa<i�a<̛a<��a<��a<�a<��a<3�a<�a<��a<�a<��a<"�a<�a<t�a<h�a<�a<8�a<�a<��a<p�a<ȍa<#�a<��a<�a<��a<z�a<��a<K�a<��a<G�a<ҙa<&�a<_�a<��a<֖a<U�a<�a<�a<H�a<��a<4�a<��a<�a<��a<Зa<&�a<�a<��a<��a<�a<�a<��a< �a<i�a<A�a<��a<��a<�a<R�a<!�a<��a<M�a<l�a<��a<��a<��a</�a<(�a<֏a<�a<��a<��a<�a<�a<��a<|�a<^�a<�a<܇a<{�a<\�a<Y�a<Z�a<A�a<�a<��a<�a<��a<�a<рa<3~a<O{a<&xa<ua<�qa<,oa<�la<	ka<�ia<Zia<�ia<Xja<�ka<{ma<xoa<�qa<�sa<Bua<�va<�wa<&xa<Fxa<�wa<Mwa<pva<�ua<�ta<�sa<�ra<era<-ra<<ra<�ra<�ra<[sa<�sa<�sa<�sa<\sa<qra<qa<loa<8ma<�ja<ha<�ea<ca<aa<k_a<o^a<
^a<m^a<n_a<aa<ca<�ea<4ha<�  �  Lka<�ma<�oa<�qa<sa<�sa<sta<Yta<Pta<�sa<Vsa<�ra<�ra<�ra<�ra<bsa<ta<$ua<6va<Xwa<�xa<?ya<�ya<�ya<�ya<�xa<�wa<=va<qta<�ra<�pa<;oa<�ma<5ma<�la<[ma<�na<Cpa<�ra<\ua<Yxa<|{a<r~a<_�a<�a<)�a<ɇa<
�a<щa<-�a<s�a<1�a<Y�a<;�a<b�a<ڊa<w�a<V�a<n�a<Ԏa<��a<|�a<��a<o�a<�a<�a<��a<|�a<�a<R�a<h�a<P�a<J�a<��a<�a<U�a<̈́a<#�a<2�a<��a<��a<��a<~�a< �a<z�a<��a<��a<�a<�a<��a<r�a<E�a<��a<��a<p�a<ȗa<��a<U�a<��a<ԗa<��a<`�a<�a<��a<T�a<��a<��a<�a<ۙa<@�a<U�a<
�a<��a<F�a<��a<�a<V�a<w�a<͇a<B�a<�a<o�a<O�a<o�a<̐a<��a<1�a<
�a<��a<��a<�a<N�a<ԙa<g�a<`�a<��a<��a<וa<|�a<�a<7�a<P�a<ߕa<]�a<�a<}�a<��a<��a<��a<#�a<��a<��a<l�a<ߍa<U�a<��a<J�a<�a<��a<z�a<�a<^�a<��a<x�a<�a<�a<�a<��a<͌a<7�a<N�a<��a<Џa<a�a<��a<��a<�a<�a<��a<j�a<��a<��a<��a<e�a<��a<y�a<��a<��a<O�a<��a<{�a<�a<ڀa<k~a<�{a<�xa<�ua<�ra<pa<�ma<la<�ja<Fja<�ja<2ka<�la<!na<pa<�qa<�sa<uua<�va<�wa<�wa<xa<�wa<�va<�ua<�ta<�sa<�ra<�qa<kqa<Rqa<=qa<�qa</ra<�ra<Fsa<dsa<�sa<+sa<ora<5qa<yoa<sma<ka<�ha<7fa<�ca<�aa<N`a<}_a<�^a<w_a<W`a<�aa<�ca<Ifa<�ha<�  �  %la<Zna<?pa<�qa<sa<~sa<�sa<�sa<Ssa<�ra<,ra<�qa<=qa<1qa<[qa<�qa<�ra<�sa<ua<ava<�wa<�xa<aya<�ya<�ya<ya</xa<�va<Kua<�sa<�qa<apa<6oa<�na<mna<�na<pa<�qa<�sa<�va<Tya<R|a<<a<�a<3�a<,�a<��a<��a<;�a<e�a<p�a<C�a<�a<�a<�a<g�a<�a<�a<!�a<��a<
�a<|�a<��a<גa<d�a<��a<��a<��a<��a<�a<=�a<I�a<o�a<ňa<q�a<��a<Y�a<��a<y�a<�a<ϊa<�a<i�a<ԑa<!�a<(�a<��a<�a<��a<�a<יa<]�a<��a<��a<0�a<�a<*�a<�a<#�a<��a<E�a<+�a<�a<��a<��a<"�a<�a<ךa<�a<��a<�a<ޔa<��a<L�a<&�a<@�a<��a<Ήa<d�a<��a<W�a<��a<z�a<{�a<��a<דa<˕a<h�a<��a<��a<��a<��a<+�a<k�a<p�a<l�a<q�a<��a<�a<��a<͓a<�a<��a<F�a<�a<��a<��a<�a<��a<�a<��a<�a<�a<��a<6�a<��a<p�a<p�a<��a<�a<��a<��a<b�a<��a<;�a<�a<�a<ǋa<W�a<��a<Q�a<��a<G�a<ʎa<��a<��a<�a<��a<;�a<�a<*�a<��a<?�a<�a<O�a<��a<��a<ʅa<��a<�a<S�a<��a<�a<�~a<W|a<�ya<�va<�sa<<qa<oa<\ma<Fla<�ka<�ka<�la<�ma<Coa<qa<�ra<zta<�ua<�va<�wa<�wa<�wa<�va<�ua<�ta<�sa<qra<Xqa<�pa<pa<�oa<�oa<^pa<�pa<�qa<Bra<�ra<�ra<�ra<Vra<Eqa<�oa<na<�ka<�ia<=ga<ea</ca<�aa<�`a<~`a<�`a<�aa<0ca<"ea<Uga<�ia<�  �  "ma< oa<�pa<�qa<�ra<5sa<6sa<�ra<ra<hqa<�pa<�oa<ooa<Foa<�oa<pa<�pa<,ra<�sa<ua<~va<�wa<�xa<uya<�ya<Pya<�xa<�wa<[va<�ta<esa<�qa<qa<bpa<Mpa<�pa<�qa<�sa<�ua<xa<�za<m}a<�a<t�a<��a<�a<y�a<�a<��a<z�a<&�a<чa<l�a<>�a<1�a<��a<6�a<�a<l�a<�a<��a<)�a<a<*�a<�a<��a<x�a<!�a<$�a<�a<W�a<��a<�a<o�a<\�a<e�a<M�a<��a<Q�a<Ȋa<i�a<��a<��a<�a<�a<��a<�a<�a<t�a<d�a<�a<K�a<e�a<d�a<{�a<��a<:�a<+�a<<�a<��a<��a<��a<��a<��a<Ǚa<{�a<��a<��a<��a<�a<��a<ԕa<��a<��a<��a<��a<��a<��a<]�a<i�a<D�a<}�a<�a<�a<̒a<Քa<p�a<�a<Øa<e�a<j�a<�a<W�a<5�a<�a<̔a<��a<Œa< �a<��a<ܑa<D�a<�a<��a<��a<o�a<1�a<u�a<v�a<�a<�a<��a<Ǒa<ʏa<i�a<D�a<�a<J�a<��a<˄a<y�a<s�a<R�a<Q�a<Ǉa<c�a<�a<��a<�a<�a<D�a<q�a<��a<!�a<όa<=�a<��a<��a<��a<:�a<T�a<��a<U�a<d�a<��a<�a<l�a<фa<	�a<��a<"�a<�a<�a<sa<,}a<�za<�wa<cua<�ra<�pa<#oa<:na<�ma<�ma<mna<Yoa<�pa<=ra<�sa<<ua<mva<1wa<�wa<�wa<�va<1va<�ta<�sa<ra<�pa<�oa<�na<Bna<�ma<!na<�na<Uoa<?pa<	qa<�qa<Ura<cra<-ra<Nqa<Fpa<�na<�la<�ja<�ha<�fa<�da<�ca<�ba<wba<�ba<�ca<�da<�fa<�ha<�ja<�  �  -na<�oa<(qa<"ra<�ra<�ra<`ra<�qa<�pa<�oa<�na<�ma<\ma<'ma<Rma<�ma<�na<Cpa<�qa<�sa<@ua<�va<xa<ya<�ya<�ya<7ya<�xa<}wa<,va<�ta<�sa<�ra<�ra<|ra<sa<ta<�ua<�wa<�ya<5|a<�~a<!�a<�a<�a<>�a<6�a<��a<��a<=�a<҆a<�a<��a<B�a<�a<i�a<	�a<��a<f�a<�a<ǋa<ҍa<��a<�a<]�a<?�a<��a<f�a<Ēa<�a<��a<�a<��a<X�a<P�a<��a<m�a<��a<��a<��a<F�a<)�a<�a<�a<ٕa<9�a<B�a<�a<�a<��a<��a<�a<�a<��a<��a<��a<�a<�a<�a<��a<��a<��a<�a<t�a<��a<��a<=�a<��a<.�a<q�a<E�a<ۖa<�a<H�a<x�a<�a<��a<؍a<��a<��a<_�a<j�a<Րa<��a<5�a<��a<<�a<R�a<��a<B�a<��a<;�a<&�a<�a<r�a<�a<Ƒa<��a< �a<��a<��a<5�a<��a<�a<�a<1�a<�a<��a<�a<�a<0�a< �a<��a<�a<Վa<ڌa<��a<7�a<�a<��a<��a<��a<L�a<@�a<z�a<�a<_�a<��a<��a<4�a<d�a<.�a<W�a<�a<��a<�a<�a<(�a<��a<�a<,�a<��a<2�a<]�a<��a<B�a<�a<��a<�a<�a<Ѓa< �a<āa<�a<0~a<�{a<gya<wa<�ta<�ra<fqa<Ypa<�oa<�oa<\pa<6qa<kra<�sa<ua<2va<�va<pwa<�wa<-wa<?va<ua<�sa<ra<Fpa<�na<�ma<�la<�ka<�ka<	la<�la<�ma<�na<�oa<�pa<nqa<�qa<ra<�qa<�pa<coa<�ma<la<7ja<dha<�fa<�ea<�da<�da<�da<�ea<�fa<|ha<]ja<Ela<�  �  7oa<�pa<�qa<Ira<tra<-ra<�qa<wpa<Xoa<na<�la<�ka<ka<�ja<�ja<�ka<�la</na<�oa<�qa<�sa<�ua<Pwa<�xa<kya<�ya<�ya<iya<�xa<�wa<�va<�ua<!ua<�ta<�ta<Tua<lva<�wa<�ya<�{a<�}a<�a<�a<��a<G�a<R�a<Ɔa<�a<��a<�a<6�a<V�a<��a<��a<҂a<��a<��a<��a<�a<�a<�a</�a<*�a<�a<��a<͒a<��a<��a<��a<ےa<Ցa<��a<��a<|�a<t�a<��a<a<�a<̍a<܎a<k�a<�a<��a<7�a<��a<ܗa<��a<֘a<��a<�a<�a<��a<@�a<ϒa<��a<c�a<ҏa<w�a<ďa<[�a<d�a<ْa<E�a<�a<W�a<��a<��a<0�a<N�a<�a<$�a<��a<��a<�a<u�a<�a<��a<5�a<Ώa<�a<��a<��a<ݒa<0�a<��a<�a<$�a<Θa<&�a< �a<c�a<p�a<�a<o�a<��a<&�a<��a<e�a<��a<9�a<m�a<�a<�a<�a<a�a<��a<�a<��a<��a<��a<i�a<��a<��a< �a<g�a<��a<��a<Z�a<*�a<c�a<�a<�a<p�a<d�a<a�a<��a<��a<��a<`�a<��a<x�a<��a<��a<.�a<>�a<M�a<,�a<;�a<H�a<ڀa<�a<a<�~a<a<�a<��a<r�a<8�a<��a<o�a<^�a<�a<�a<ۀa<"a<}a<{a<�xa<�va<
ua<�sa<�ra<:ra<,ra<�ra<[sa<5ta<Gua<-va<wa<�wa<�wa<vwa<�va<�ua<ta<=ra<apa<na<�la<=ka<Ija<�ia<�ia<�ia<ja<�ka<�la<5na<goa<�pa<Mqa<�qa<�qa<qa<Apa<�na<yma<�ka<`ja<�ha<�ga<9ga<�fa<@ga<�ga<
ia<�ja<la<�ma<�  �  fpa<xqa<6ra<�ra<Gra<�qa<�pa<joa<�ma<Yla<�ja<�ia<�ha<qha<�ha<?ia<wja<la<�ma<.pa<nra<�ta<uva<xa<Nya<'za<bza<Cza<�ya<Mya<rxa<�wa<_wa<wa<Cwa<�wa<�xa<za<�{a<m}a<�a<h�a<�a<��a<ƅa<h�a<��a<C�a<��a<̈́a<��a<��a<��a<Հa<��a<��a<?�a<j�a<��a<�a<3�a<��a<�a<3�a<��a<��a<��a<-�a<0�a<Փa<1�a<g�a<F�a<s�a<��a<<�a<3�a<�a<�a<"�a<T�a<��a<E�a<��a<��a<y�a<�a<��a</�a<,�a<�a<U�a<��a<�a<k�a<@�a<s�a<,�a<\�a< �a<B�a<��a<��a<^�a<C�a<՗a<�a<��a<x�a<n�a<��a<�a<��a<��a<F�a<,�a<0�a<��a<B�a<^�a<ݒa<��a<��a<�a<*�a<�a<�a<`�a<`�a<Әa<��a<��a<�a<��a<�a<�a<w�a<0�a<I�a<��a<�a<��a<��a<�a<��a<^�a<�a<�a<�a<��a<Ǖa<K�a<q�a<@�a<��a<P�a<�a<��a<k�a<��a<Y�a<Q�a<��a<b�a<&�a<=�a<
�a<��a<�a<�a<��a<}�a<
�a<G�a<"�a<��a<^�a<�a<#�a<�~a<a}a<�|a<�|a<�|a<�}a<�~a<�a<�a<�a<��a<�a<	�a<��a<�a<�a<w~a<�|a<�za<�xa<Pwa<�ua< ua<�ta<kta<�ta<Dua<�ua<�va<{wa<�wa<;xa<xa<_wa<Fva<�ta<sa<�pa<�na<�la<�ja<ia<�ga<Dga<ga<�ga<]ha<�ia<ka<�la<Sna<�oa<�pa<vqa<�qa<�qa<�pa<	pa<�na<�ma<0la<ka<%ja<�ia<Zia<�ia<0ja<1ka<Zla<�ma<9oa<�  �  �qa<Hra<�ra<�ra<ra<9qa<�oa<[na<tla<�ja<ia<�ga<�fa<3fa<qfa<�fa<nha<ja<7la<�na<qa<�sa<�ua<�wa<ya<Xza<�za<4{a<
{a<�za<+za<�ya<Vya<(ya<bya< za<�za<|a<�}a<8a<��a<��a<?�a<E�a<!�a<]�a<B�a<��a<��a<��a<%�a<�a<�a<�~a<N~a<y~a< a<'�a<	�a<
�a<��a<�a<��a<1�a<^�a<>�a<��a<��a<͔a<�a<n�a<ēa<�a<V�a<Ǒa<b�a<f�a<��a<+�a<�a<&�a<l�a<��a<��a<��a< �a<)�a<��a<ߗa<~�a<�a<��a<�a<)�a<{�a<B�a</�a<�a<'�a<��a<T�a<�a<��a<�a<(�a<��a<��a<��a<��a<ښa<��a<,�a<7�a<9�a<�a<�a<A�a<��a<��a<��a<�a<��a<�a<��a<i�a<I�a<��a<Йa<~�a<��a<o�a<��a<Փa<��a<n�a<D�a<��a<�a<
�a<Ȉa<̈a<��a<ъa<[�a<.�a<��a<�a<e�a<��a<l�a<��a<˕a<a�a<w�a<B�a<	�a<��a<��a<��a<�a<��a<z�a<ɍa<H�a<�a<��a<F�a<ːa<��a<o�a<��a<;�a<x�a<K�a<�a<<�a<a<7�a<3~a<W|a<<{a<�za<aza< {a<�{a<}a<S~a<�a<�a<�a<ςa<��a<�a<�a<7�a<�a<~a<l|a<�za<]ya<xa<Rwa<�va<�va<�va<wa<�wa<2xa<�xa<�xa<�xa<Xxa<6wa<�ua<ta<�qa<�oa<1ma<�ja<�ha<ga<�ea<ea<�da<eea<ofa<�ga<�ia<>ka<8ma<�na<Hpa<8qa<�qa<ra<�qa<3qa<.pa<'oa<�ma<ma<5la<�ka<�ka<�ka<Bla<"ma<$na<boa<xpa<�  �  gra<�ra<�ra<�ra<�qa<�pa<1oa<Xma<Nka<Iia<zga<�ea<�da<dda<xda<7ea<|fa<fha<�ja<9ma<�oa<�ra<ua<Hwa<ya<�za<9{a<�{a<�{a<�{a<�{a<E{a<{a<{a<D{a<�{a<�|a<�}a<Da<ǀa<I�a<��a<�a<̅a<S�a<p�a<�a<-�a<�a<x�a<�a<[a<~a<}a<||a<�|a<.}a<^~a<�a<b�a<��a<Ça<��a<a�a<ُa<ܑa<��a<��a<F�a<��a<o�a<�a<��a<	�a<�a<N�a<1�a<}�a<�a<ɔa<Օa<֖a<ܗa<��a<N�a<a�a<U�a<��a<r�a<�a<�a<�a<��a<��a<ˋa<N�a<l�a<�a<K�a<�a<}�a<T�a<v�a<Ƒa<�a<A�a<�a<��a<��a<�a<E�a<��a<[�a<��a<��a<Зa<�a<��a<J�a<l�a<��a<b�a<�a<ߘa<��a<�a<^�a<�a<��a<v�a<�a<�a<Ӓa<c�a<��a<��a<��a<'�a<;�a<Άa<�a<a<�a<ъa<Ōa<ގa<��a<ǒa<H�a<j�a<�a<"�a<�a<T�a<~�a<k�a<T�a<?�a<c�a<a<^�a<h�a<��a<��a<��a<��a<S�a<�a<<�a<��a<��a<�a<�a<��a<Άa<��a<1�a<�~a<R|a<�za<Nya<�xa<�xa<ya<za<v{a<}a<�~a<@�a<��a<l�a<�a<�a<��a<�a<��a<ga<�}a<|a<{a<za<ya<�xa<lxa<nxa<�xa<ya<uya<�ya<�ya<#ya<�xa<Bwa<�ua<~sa<qa<zna<�ka<Pia<ga<*ea<�ca<%ca<ca<�ca<�da<%fa<ha<ja<-la<na<�oa<qa<ra<Lra<ara<�qa<Rqa<upa<�oa<�na<�ma<�ma<ama<�ma<na<�na<�oa<�pa<�qa<�  �  
sa<�sa<Msa<�ra<�qa<Zpa<�na<~la<qja<<ha<Pfa<�da<�ca<ca<�ba<�ca<ea<+ga<�ia<:la<oa<�qa<�ta<�va<ya<�za<�{a<o|a<�|a<�|a<}|a<|a<N|a<I|a<�|a<1}a<~a<a<��a<Ɂa<B�a<��a<��a<_�a<��a<��a<��a<��a<I�a<��a<�a<7~a<�|a<�{a<5{a<	{a<�{a<}a<�~a<@�a<փa<Άa<ωa<��a<Z�a<��a<��a<�a<ؕa<9�a<H�a<�a<��a<D�a<Ȕa<��a<��a<�a<V�a<�a<�a<ėa<�a<g�a<�a<�a<t�a<��a<'�a<`�a<:�a<�a<��a<w�a<��a<�a<�a<z�a<�a<ǈa<-�a<.�a<`�a<�a<A�a<��a<��a<j�a<a<k�a<ۛa<��a<Q�a<��a<ƙa<�a<L�a<�a<��a<ۗa<��a<��a<D�a<ҙa<��a<��a<�a<w�a<��a<^�a<��a<n�a<��a<��a<�a<��a<p�a<ֆa<ۅa<9�a<��a<^�a<�a<��a<ŋa<�a<#�a<:�a<��a<]�a<:�a<��a<��a<�a<��a<[�a<��a<��a<��a<5�a<Ȑa<a<͐a<<�a<��a<�a<6�a<�a<Бa<ِa<��a<��a<}�a<وa<��a<�a<�a<r}a<�za<>ya<�wa<#wa<Qwa<�wa<�xa<Qza<|a<�}a<�a<�a<6�a<�a<>�a<&�a<�a<��a<e�a<�~a<�}a<]|a<^{a<�za<za<�ya<�ya<za<za<{za<^za<=za<�ya<�xa<<wa<?ua<�ra<Opa<�ma<�ja<(ha<�ea<�ca<�ba<�aa<�aa<3ba<Ica< ea<�fa<1ia<Qka<yma<]oa<�pa<ra<�ra<�ra<�ra<Gra<lqa<�pa<�oa<?oa<oa<�na<oa<Ooa<pa<�pa<�qa<�ra<�  �  ysa<�sa<|sa<�ra<�qa<Epa<Pna<*la<�ia<�ga<pea<�ca<�ba<�aa<ba<�ba<:da<Cfa<�ha<�ka<tna<�qa<Zta<�va<�xa<�za<�{a<�|a<}a<K}a<P}a<D}a<8}a<F}a<�}a<'~a<�~a<�a<R�a<��a<ރa<�a<�a<��a<��a<e�a<��a<~�a<��a<1�a<Va<�}a<�{a<�za<2za< za<�za<|a<�}a<W�a<!�a<1�a<J�a<Z�a<"�a<��a<��a<�a<�a<��a<��a<��a<j�a<�a<a<��a<��a<ѕa<N�a<�a<ٗa<��a<X�a<�a<-�a<�a<��a<r�a<�a<,�a<��a<q�a<�a<��a<��a<�a<�a<��a<�a<ԇa<R�a<M�a<��a<D�a<�a<W�a<��a<V�a<��a<��a<�a<��a<��a<6�a<��a<�a<F�a<טa<��a<��a<��a<~�a<�a<��a<��a<.�a<%�a<��a<��a<G�a<z�a<*�a<��a<ݎa<B�a<��a<��a<�a<Մa<\�a<��a<�a<��a<шa< �a<b�a<܏a<�a<�a<;�a<@�a<Жa<ޖa<��a<�a<.�a<S�a<q�a<��a<�a<��a<��a<ɑa<�a<a�a<��a<��a<x�a<�a< �a<��a<��a<E�a<��a<��a<n�a<ca<�|a<za<;xa<�va<?va<Hva<�va<xa<�ya<s{a<X}a<9a<րa<-�a<�a<`�a<_�a<ւa<�a<�a<�a<�~a<W}a<F|a<y{a<�za<�za<�za<�za<�za<�za<�za<�za<�ya<�xa<wa<5ua<�ra<pa<
ma<5ja<\ga<�da<�ba<�aa<�`a<�`a<@aa<nba<da<Ifa<�ha<�ja<1ma<=oa<�pa< ra<�ra<$sa<sa<�ra<#ra<�qa<�pa<9pa<�oa<�oa<�oa<Npa<�pa<�qa<mra<sa<�  �  ita<%ta<ta<�sa<�ra<�qa<+pa<�na<�la<fka<�ia<�ha<�ga<gga<�ga<#ha<via<ka<�la</oa<_qa<�sa<�ua<(xa<�ya<u{a<>|a<(}a<�}a<�}a<$~a<�}a<)~a<d~a<�~a<wa<�a<!�a<
�a<O�a<e�a<��a<j�a<��a<'�a<�a<u�a<��a<��a<|�a<3�a<�a<�a<�a<�~a<#a<�a<��a<��a<?�a<��a<��a<e�a<�a<��a<�a<��a<&�a<��a<��a<ߖa<��a<��a<G�a<J�a< �a<Y�a<��a<�a<{�a<�a<��a<j�a<'�a<1�a<ߙa<Йa<˘a<ɗa<+�a<Ôa<��a<�a<>�a<ʍa<��a<ǋa<��a<ȋa<�a<Սa<�a<�a<Ւa<��a<��a<q�a<ҙa<�a<��a<ۛa<T�a<�a<��a<�a<a�a<�a<��a<��a<��a<��a<�a<_�a<�a<)�a<��a<	�a<��a<	�a<��a<V�a<|�a<��a<g�a<��a<u�a<�a<��a<��a<��a<r�a<=�a<9�a<{�a<>�a<ҏa<̑a<%�a<��a<��a<��a<��a<�a<��a<�a<��a<��a<�a<S�a<ڒa<��a<U�a<o�a<`�a<��a<��a<ؒa<��a<��a<,�a<͏a<2�a<1�a<�a<��a<-�a<҂a<{�a<�~a<�|a<�{a<Y{a<{a<�{a<&|a<;}a<r~a<�a<�a<�a<�a<��a<�a<d�a<I�a<��a<y�a<��a<=a<a~a<a}a<�|a<5|a<�{a<�{a<{a<�{a<�{a<�{a<{a<)za<�ya<�wa<jva<Gta<_ra<�oa<�ma<yka<�ia<%ha<�fa<Wfa<fa<xfa<ga<zha<#ja<�ka<�ma<)oa<�pa<�qa<�ra<xsa<�sa<�sa<tsa<sa<gra<�qa<�qa<=qa<Jqa<Fqa<�qa<ra<�ra<Ssa<�sa<�  �  �sa<5ta<	ta<�sa<�ra<�qa<Lpa<�na<ma<�ka<�ia<�ha<�ga<�ga<�ga<nha<{ia<*ka<ma<Zoa<�qa<ta<va<Dxa<�ya<A{a<N|a<}a<j}a<�}a<�}a<�}a<-~a<G~a<�~a<8a<�a<��a<�a<'�a<3�a<$�a< �a<��a<��a<׆a<��a<υa<ӄa<��a<f�a<B�a<5�a<na<a<Pa<�a<��a<y�a<z�a<��a<&�a<��a<	�a<.�a<6�a<��a<�a<ҕa<T�a<h�a<|�a<r�a<P�a<,�a<��a<$�a<e�a<˖a<y�a<�a<��a<6�a<��a<�a<��a<��a<͘a<�a<V�a<Ӕa<��a<9�a<y�a<��a<��a<�a<΋a<�a<��a<эa<X�a<0�a<�a<�a<ܖa<��a<�a<�a<��a<��a<�a<��a<E�a<Ԛa<c�a<ܙa<��a<X�a<b�a<��a<�a<U�a<��a<�a<#�a<�a<��a<�a<Θa<y�a<��a<a<��a<��a<��a<�a<��a<��a<��a<��a<B�a<c�a<��a<i�a<�a<בa<J�a<˔a<��a<j�a<��a<Жa<c�a<ݕa<M�a<��a<��a<6�a<��a<c�a</�a<H�a<g�a<�a<��a<m�a<X�a<ޑa<�a<��a<P�a<a�a<6�a<Շa<_�a<�a<��a<�~a<*}a< |a<{a<M{a<�{a<b|a<r}a<�~a<�a<6�a<9�a<#�a<y�a<��a<��a<�a<%�a<E�a<M�a<Ea<D~a<>}a<�|a<|a<�{a<�{a<�{a<|{a<W{a<%{a<�za<Bza<Qya<�wa<�va<rta<pra< pa<�ma<�ka<�ia<&ha<ga<tfa<Nfa<�fa<{ga<�ha<Kja<�ka<�ma<Goa<�pa<�qa<�ra<dsa<�sa<�sa<"sa<�ra<Sra<�qa<eqa<qa<qa<'qa<zqa<ra<�ra<sa<�sa<�  �  �sa<ta<�sa<�sa<�ra<�qa<�pa<oa<�ma<�ka<�ja<�ia<�ha<qha<Zha<Iia<.ja<�ka<�ma<�oa<ra<;ta<Yva<Exa<�ya<*{a<,|a<�|a<}a<�}a<E}a<U}a<^}a<�}a<�}a<{~a<Xa<&�a<Z�a<n�a<�a<�a<҅a<��a<̆a<�a<��a<��a<�a<��a<ׂa<��a<��a<�a<�a<�a<��a<܁a< �a<B�a<<�a<��a<��a<7�a<_�a<4�a<��a<��a<��a<�a<-�a<@�a<��a<��a<T�a<a�a<h�a<��a<�a<��a<g�a<�a<�a<]�a<ԙa<֙a<t�a<�a<�a<��a<�a<j�a<��a<�a<��a<j�a<�a<d�a<̌a<s�a<��a<�a<��a<��a<Z�a<�a<��a<�a<�a<l�a<՛a<��a<q�a<ؚa<%�a<��a<�a<�a<��a<ʘa<јa<=�a<��a</�a<��a<ǚa<�a<��a<�a<ؘa<��a<�a<�a<�a<�a<d�a<Ȍa<~�a<Ɗa<.�a<��a<��a< �a<Z�a<̎a<��a<�a<��a<̔a<ŕa<S�a<��a<��a<�a<��a<��a<�a<'�a<~�a<�a<��a<��a<t�a<��a<Ƒa<9�a<;�a<
�a<��a<ѐa<֏a<S�a<��a<i�a<.�a<хa<p�a<�a<aa<~a<�|a<&|a<4|a<?|a<)}a<�}a<a<P�a<e�a<j�a<"�a<��a<��a<p�a<ǂa<�a<	�a<�a<�~a<l}a<�|a<�{a<Y{a<{a<�za<�za<�za<3{a<�za<�za<za<+ya<xa<�va<�ta<�ra<�pa<Mna<Fla<�ja<�ha<�ga<
ga<ga<lga<*ha<nia<�ja<_la<�ma<�oa<�pa<ra<�ra<7sa<�sa<4sa<�ra<[ra<�qa<%qa<�pa<�pa<Dpa<�pa<�pa<Iqa<�qa<�ra<_sa<�  �  sa<�sa<�sa<�sa<�ra<"ra<qa<�oa<Ena<�la<�ka<sja<�ia<jia<�ia<0ja<0ka<�la<�na<�pa<�ra<�ta<�va<zxa<�ya<7{a<�{a<g|a<�|a<�|a<�|a<�|a<n|a<�|a<�|a<b}a<[~a<9a<��a<��a<	�a<;�a<P�a<�a<��a<�a<��a<Z�a<��a<��a<��a<��a<Ła<#�a<ހa<�a<��a<��a<1�a<�a<�a<l�a<��a<Ȏa<ΐa<H�a<͓a<��a<<�a<��a<��a<Y�a<�a<Ҕa<e�a<q�a<O�a<��a<8�a<��a<��a<W�a<)�a<˘a<X�a<y�a<��a<�a<�a<�a<��a<�a<x�a<ېa<��a<p�a<Ӎa<��a<ˍa<_�a<|�a<�a<q�a<B�a<��a<��a<��a<�a<��a<>�a<Q�a<�a<��a<�a<f�a<Ęa<)�a<ؗa<��a<��a<�a<X�a<�a<h�a<�a<B�a<m�a<C�a<�a<�a<͗a<`�a<��a<Ԓa<�a<9�a<��a<w�a<��a<V�a<��a<��a<��a<'�a<��a<1�a<��a<
�a<�a<ϕa<`�a<K�a< �a<��a<ٔa<��a<)�a<7�a<��a<��a<��a<��a<��a<ܐa<�a<\�a<��a<��a<@�a<��a<�a<e�a<�a<�a<ֈa<��a<C�a<K�a<m�a<�~a<�}a<;}a<}a<P}a<�}a<�~a<�a<��a<��a<قa<6�a<��a<��a<��a<H�a<?�a<"�a<�~a<�}a<}|a<�{a<�za<Fza<za<�ya<za< za<Jza<Iza<9za<�ya<7ya<xa<�va<-ua<Bsa<5qa<$oa<ma<`ka<�ia<�ha<0ha<ha<Wha<&ia<Cja<�ka<ma<�na<pa<9qa<ra<�ra<	sa<sa<�ra<1ra<�qa<�pa<Epa<�oa<poa</oa<yoa<�oa<dpa<qa<�qa<�ra<�  �  �ra<!sa<esa<asa<sa<�ra<dqa<Cpa<oa<�ma<�la<�ka<ka<�ja<ka<�ka<�la<na<�oa<�qa<vsa<Xua<+wa<�xa< za<�za<�{a<�{a<�{a<�{a<�{a<L{a<"{a<={a<r{a<�{a<�|a<�}a<6a<��a<�a<h�a<̈́a<΅a<}�a<ӆa<��a<��a<��a<J�a<��a<��a<�a<��a<A�a<��a<.�a<�a<��a<8�a<A�a<Q�a<J�a<9�a<$�a<��a<��a<��a<�a<�a<��a<k�a<��a<|�a<�a<�a<�a<+�a<��a<j�a<U�a<V�a<5�a<�a<Ԙa<,�a<K�a<�a<r�a<c�a<�a<Ȕa<��a<�a<ΐa<�a<+�a<�a<1�a<ȏa<ؐa<�a<��a<�a<��a<��a<g�a<A�a<��a<�a<�a<��a<a<�a<@�a<p�a<іa<P�a<�a<,�a<��a<�a<��a<r�a<�a<��a<�a<�a<��a<�a<;�a<��a<6�a<��a<�a<`�a<
�a<�a< �a<��a<یa<o�a<=�a<]�a<��a<�a<,�a<[�a<m�a<ەa<%�a< �a<��a<�a<�a<��a<�a<�a<,�a<��a<#�a<�a<5�a<��a<�a<j�a<��a<�a<�a<��a<��a<��a<F�a<^�a<z�a<|�a<}�a<s�a<؁a<N�a<Xa<�~a<m~a<�~a<a<�a<Ԁa<��a<g�a</�a<��a<��a<J�a<��a<��a<x�a<3a<�}a<r|a<-{a</za<Sya<�xa<�xa<�xa<�xa<ya<Vya<�ya<�ya<uya<ya<xa<wa<ua<�sa<�qa<-pa<Lna<�la<Oka<.ja<�ia<}ia<�ia<�ja<gka<�la<�ma<4oa<`pa<�qa<Qra<�ra<�ra<�ra<&ra<Oqa<�pa<�oa<�na<[na<�ma<�ma<�ma<sna<oa<�oa<�pa<�qa<�  �  �qa<�ra<sa<Hsa<Asa<�ra<ra<Hqa<,pa<oa<na<)ma<�la<qla<�la<<ma<*na<loa<qa<�ra<�ta<Jva<�wa<(ya<za<�za<,{a<0{a<�za<�za<Eza<�ya<�ya<�ya<�ya<gza<I{a<t|a<�}a<Da<	�a<��a<�a<I�a<'�a<Ԇa<;�a<	�a<Ɇa<V�a<��a<�a<R�a<�a<��a<�a<��a<҅a<�a<��a<��a<X�a<W�a<�a<��a<�a<��a</�a<w�a<0�a<�a<r�a<��a<�a<��a<X�a<O�a<��a<�a<��a<�a<�a<Q�a<5�a<�a<Øa<�a<�a<��a<�a<�a<��a<��a<f�a<5�a<]�a<�a<��a<Ґa<o�a<=�a<d�a<͔a<+�a<��a<��a<��a<l�a<��a<��a<X�a<��a<�a<�a<ߖa<��a<D�a<̔a<��a<��a<��a<��a<S�a<:�a<)�a<ǘa<c�a<��a<��a<B�a<|�a<m�a<;�a<��a<6�a<��a<p�a<�a<ǎa<q�a<��a<�a<��a<��a<Бa<	�a< �a<��a<��a<��a<�a<��a<�a<��a<�a<��a<~�a<v�a<��a<��a<��a<��a<a<�a<��a<\�a<ُa<#�a<j�a<+�a<��a<��a<��a<+�a<��a<��a<Æa<ׄa<;�a<�a<�a<S�a<*�a<"�a<��a<C�a<ہa<��a<;�a<��a<كa<��a<��a<3�a<�a<�a<;~a<x|a<{a<�ya<�xa<�wa<Dwa<wa<'wa<`wa<�wa<rxa<�xa<�xa<ya<�xa<0xa<[wa<	va<�ta<sa<:qa<�oa<na<�la<�ka<Gka<ka<gka<�ka<�la<�ma<oa<<pa<$qa<�qa<}ra<�ra<vra<ra<=qa<vpa<noa<_na<�ma<�la<ela<?la<mla<�la<�ma<�na<�oa<�pa<�  �  �pa<�qa<�ra<6sa<dsa<3sa<�ra<ra<Cqa<Gpa<�oa<�na<Sna<=na<Sna<oa<�oa<qa<�ra<�sa<�ua<wa<~xa<sya<>za<�za<�za<�za<za<�ya<�xa<�xa<xa<�wa<!xa<�xa<�ya<�za<T|a<�}a<�a<��a<1�a<˄a<�a<܆a<c�a<��a<��a<2�a<Æa<M�a<��a<��a<��a<�a<y�a<��a<��a<V�a<�a<��a<B�a<Ӑa<*�a<�a<Ǔa<��a<��a<��a<ߒa<�a<P�a<��a<��a<��a<��a<ԏa<r�a<M�a<��a<��a<�a<D�a<y�a<T�a<�a<"�a<��a<��a<Ǘa<ߖa<��a<Ӕa<�a<�a<��a<Y�a<��a<�a<�a<�a<�a<N�a<f�a<|�a<&�a<��a<��a<R�a<ԙa<Әa<̗a<��a<��a<|�a<��a<�a<��a<�a<A�a<�a<�a<ڕa<�a<�a<טa<D�a<��a<e�a<ߘa<*�a<�a<ӕa<n�a<U�a<�a<%�a<��a<*�a<Z�a<��a<X�a<3�a<�a<�a<�a<��a<��a<�a<Еa<5�a<X�a<�a<ȑa<_�a<'�a<ԍa<݌a<0�a<��a<ڋa<�a<��a<N�a<��a<Ύa<h�a<�a<�a<��a<�a<5�a<�a<a�a<��a<�a<��a<�a<��a<��a<�a<݁a<Ӂa<=�a<��a<�a<��a<�a<5�a<�a<��a<ła<��a<=�a<�~a<�|a<,{a<�ya<xa<�va<�ua<~ua<Yua<zua<va<~va<&wa<�wa<Zxa<�xa<�xa<Jxa<�wa<�va<bua< ta<ira<qa<�oa<pna<�ma<�la<�la<ma<�ma<fna<(oa<)pa<qa<�qa<ara<�ra<�ra<ra<�qa<ppa<Yoa<na<ma<�ka<ka<�ja<cja<�ja<(ka<la<9ma<Dna<�oa<�  �  	pa<9qa<Mra<sa<xsa<�sa<fsa<�ra<nra<�qa<�pa<dpa<pa<�oa<0pa<�pa<�qa<�ra<�sa<Oua<�va<�wa<�xa<�ya<Cza<~za<Aza<�ya<Jya<ixa<�wa<�va<eva<Eva<Vva<�va<�wa<ya<�za<�|a<v~a<��a<n�a<�a<��a<Ɔa<��a<�a<0�a<(�a<�a<��a<]�a<L�a<N�a<��a<E�a<0�a<j�a<��a<-�a<��a<@�a<y�a<��a<F�a<��a<̓a<Q�a<��a<�a<ِa<��a<�a<=�a<�a<ɍa<�a<Ǝa<��a<�a<l�a<ԓa<m�a<��a<��a<��a<�a<:�a<�a<��a<�a< �a<!�a<c�a<Ȕa<[�a<1�a<b�a<˔a<�a<\�a<c�a<��a<G�a<�a<��a<��a<��a<�a<�a<�a<Ėa<[�a<�a<˒a<�a<J�a<��a< �a<��a<X�a<l�a<��a<�a<-�a<�a<�a<g�a<y�a<F�a<��a<ڗa<��a<˕a<��a<��a<ڒa<Q�a<�a<�a<T�a<ؒa<��a<`�a<%�a<��a<.�a<J�a<�a<��a<��a<��a<C�a<��a<�a<��a<.�a<4�a<f�a<�a<�a<T�a<�a<�a<Ɍa<Ӎa<��a<?�a<��a<��a<I�a<��a<��a<W�a<�a<X�a<�a<��a<Z�a<|�a<كa<��a<��a<��a<��a<r�a<��a<��a<��a<4�a<��a<��a<�a<xa<�}a<�{a<�ya<�wa<Vva<4ua<;ta<�sa<�sa<�sa<[ta<5ua<�ua<�va<�wa<	xa<oxa<Fxa<�wa<7wa<va<ua<�sa<Zra<0qa<-pa<]oa<�na<�na<�na<(oa<�oa<}pa<`qa<�qa<wra<�ra<�ra<qra<�qa<�pa<�oa<Rna<�la<�ka<Nja<ria<�ha<�ha<�ha<�ia<fja<�ka<ma<�na<�  �  oa<�pa<ra<�ra<�sa<�sa<ta<�sa<Jsa<�ra<Qra<�qa<�qa<�qa<�qa<=ra<sa<ta<<ua<rva<�wa<�xa<�ya<za<Nza<Pza<�ya<ya<Axa<Twa<}va<�ua<ua<�ta<�ta<Tua<va<�wa<8ya<?{a<k}a<wa<��a<��a<k�a<��a<Շa<��a<��a<�a<��a<�a<Ɉa<��a<�a<;�a<׉a<͊a<Ջa<$�a<��a<ݏa<�a<L�a<�a<��a<��a<��a<�a<�a<ߐa<Џa<��a<��a<׌a<4�a<9�a<s�a<�a<B�a<��a<-�a<Œa<c�a<�a<p�a<��a<!�a<��a<��a<j�a<Ƙa<5�a<��a<Ԗa<B�a<�a<a<�a<g�a<��a<ėa<��a<c�a<3�a<��a<�a<ۚa<d�a<a<w�a<�a<��a<B�a<��a<c�a<]�a<��a<}�a<u�a<	�a<�a<�a<��a<Ҕa<*�a<k�a<��a<B�a<��a<��a<`�a<ǘa<ڗa<�a<�a<"�a<r�a<ؓa<��a<��a<ۓa<I�a<�a<��a<��a<��a<Öa<��a<*�a<z�a<j�a<ɒa<;�a<��a<�a<$�a<ˊa<��a<ǈa<~�a<Z�a<�a<��a<��a<��a<��a<ōa<��a<o�a<��a<��a<�a<Y�a<7�a<��a<��a<O�a<�a<��a<�a<k�a<%�a<�a<�a<@�a<`�a<r�a<{�a<"�a<��a<z�a<L�a<��a<�~a<�|a<�za<�xa<�va<�ta<vsa<�ra<ra<�qa<ora<�ra<�sa<�ta<�ua<�va<�wa<7xa<Ixa<.xa<�wa<wa<�ua<�ta<�sa<�ra<�qa<�pa<fpa<6pa<^pa<�pa<#qa<�qa<>ra<�ra<,sa<*sa<�ra<Pra<�qa<(pa<�na<2ma<�ka<0ja<�ha<�ga<4ga<+ga<=ga<�ga<ia<Kja<�ka<rma<�  �  zna<4pa<�qa<�ra<�sa<8ta<yta<ita<7ta<�sa<�sa<)sa<sa<sa< sa<�sa<gta<`ua<]va<jwa<gxa<Aya<�ya<Vza<�za<za<�ya<�xa<�wa<�va<Kua<bta<�sa<2sa<Nsa<�sa<�ta<!va<�wa<za<l|a<�~a<�a<K�a< �a<��a<�a<шa<{�a<��a<�a<�a<�a<�a<m�a<��a<F�a<N�a<#�a<z�a<��a<͐a<ܑa<Ғa<d�a<Гa<��a<#�a<��a<q�a<2�a<�a<m�a<Z�a<e�a<׊a<��a<��a<��a<׌a<Y�a<��a<�a<ēa<��a<�a<2�a<T�a<Йa<��a<�a<��a<+�a<��a<$�a<��a<j�a<)�a<i�a<Зa<D�a< �a<��a<U�a<ךa<8�a<7�a<�a<P�a<V�a<%�a<��a<�a<'�a<{�a<�a<�a<>�a<�a<�a<��a<��a<�a<f�a<�a<��a<�a<<�a<�a<ԙa<�a<˙a<\�a<ǘa<��a<>�a<s�a<ԕa<]�a<��a<�a<1�a<��a<�a<|�a<ޖa<�a<!�a<��a<a�a<9�a<�a<o�a<��a<��a<��a<��a<i�a<!�a<^�a<�a<�a<m�a<S�a<_�a<��a<�a<O�a<k�a<�a<��a<Ǐa<a�a<܎a<�a<�a<��a<��a<O�a<y�a<|�a<چa<��a<B�a<a�a<I�a<P�a<3�a< �a<p�a<��a<��a<�a<O�a<+~a<�{a<�ya<Jwa<Qua<}sa<ra<!qa<�pa<�pa<qa<�qa<�ra<ta<Aua<ava<\wa<�wa<{xa<oxa<xa<�wa<�va<�ua<�ta<�sa<�ra<kra<�qa<�qa<�qa<�qa<_ra<�ra<0sa<wsa<�sa<rsa<)sa<<ra<"qa<�oa<4na<xla<�ja<�ha<�ga<ufa<�ea<�ea<�ea<�fa<�ga<ia<�ja<�la<�  �  �ma<�oa<]qa<�ra<�sa<|ta<�ta<�ta<ua<�ta<Lta<ta<�sa<ta<6ta<�ta<Mua<=va<wa<6xa<.ya<�ya<qza<zza<xza<�ya<;ya<4xa<wa<�ua<mta<�sa<�ra<Kra<Kra<�ra<�sa<ua<-wa<8ya<�{a<~a<~�a<Ђa<�a<��a<�a<4�a<��a<V�a<ڊa<��a<ߊa<��a<P�a<��a<^�a<8�a<�a<D�a<H�a<��a<��a<O�a<Փa<͓a<��a<�a<�a<ߐa<��a<�a<��a<��a<V�a<��a<��a<��a<ъa<Ћa<��a<�a<!�a<�a<��a<��a< �a<E�a<�a<~�a<o�a<[�a<�a<T�a<��a<��a<n�a<@�a<}�a<��a<3�a<ʙa<^�a<4�a<\�a<��a<��a<�a<C�a<�a<��a<��a<:�a<M�a<��a<>�a<�a<T�a<��a<"�a<��a<��a<�a<��a<Z�a<��a<��a<��a<�a<˙a<(�a<Q�a<�a<��a<a<�a<]�a<��a<t�a<�a<'�a<�a<y�a<a<I�a<��a<��a<��a<�a<U�a<'�a<��a<�a<��a<��a<ًa<,�a<i�a<;�a<[�a<̅a<&�a<f�a<��a<��a<�a<e�a<��a<��a<�a<��a<��a<ŏa<Y�a<��a<ҍa<h�a<e�a<@�a<]�a<��a<�a<��a<1�a<,�a<��a<:�a<؆a<~�a<�a<��a<��a<ԁa<�a<�}a<I{a<�xa<va<�ta<ora<?qa<pa<�oa<�oa<�oa<qa<�qa<Asa<�ta<�ua<�va<�wa<lxa<�xa<�xa<	xa<{wa<�va<�ua<�ta<�sa<osa<�ra<�ra<�ra<�ra<(sa<xsa<ta<�sa<"ta<�sa<sa</ra<�pa<Woa<�ma<�ka<�ia<1ha<�fa<sea<�da<gda<�da<�ea<�fa<Mha<�ia<�ka<�  �  �ma<poa<Tqa<�ra<�sa<�ta<)ua<Hua<-ua< ua<�ta<�ta<�ta<�ta<�ta<lua<va<�va<�wa<�xa<Vya<za<�za<�za<kza<�ya<#ya<�wa<�va<Nua<	ta<�ra<�qa<pqa<�qa<ra<sa<qta<lva<�xa<*{a<�}a<L�a<��a<�a<��a<,�a<W�a<7�a<��a<�a<T�a<��a<̋a<��a<x�a<�a<؍a<�a<��a<��a<�a<��a<��a<��a<��a<��a<�a<�a<��a<+�a<��a<�a<Ǌa<��a<�a<�a<=�a<�a<&�a<ʌa<��a<��a<ƒa<��a<��a<�a<-�a<�a<��a<Úa<��a<Y�a<�a<��a<R�a<�a< �a< �a<q�a<��a<s�a<��a<U�a<��a<�a<��a<�a</�a<�a<d�a<��a<Óa<�a<�a<��a<-�a<}�a<-�a<R�a<،a<�a<j�a<,�a<�a<��a<S�a<�a<��a<љa<L�a<|�a<<�a<��a<I�a<��a<$�a<y�a<�a<Ζa<��a<�a<6�a<r�a<��a<Ηa<��a<ėa<4�a<H�a<�a<��a<��a<��a<��a<u�a<s�a<��a<_�a<��a<2�a<B�a<��a<��a<�a<|�a<��a<��a<��a<�a<y�a<�a<�a<��a<ʎa<��a<�a<�a<�a<�a<H�a<��a<0�a<
�a<ׇa<��a<m�a<�a<��a< �a<�a<m�a<ׁa<�a<k}a<�za<gxa<�ua<�sa<�qa<Ypa<eoa<�na<�na<Soa<Apa<qa<�ra<Cta<�ua<�va<�wa<Txa<�xa<�xa<\xa<�wa<wa<Cva<�ua<�ta<ta<�sa<jsa<hsa<�sa<�sa<ta</ta<Pta<Tta<�sa<-sa<ra<�pa<oa<Zma<Rka<qia<�ga<fa<�da<da<�ca<da<�da<fa<�ga<�ia<�ka<�  �  �ma<Ooa<4qa<�ra<�sa<�ta<!ua<�ua<pua<bua<�ta<�ta<�ta<�ta<:ua<�ua<Iva<�va<�wa<�xa<�ya<zza<sza<�za<�za<�ya<�xa<�wa<�va<ua<�sa<�ra<�qa<Mqa<Oqa<�qa<�ra<vta<5va<rxa<�za<r}a<6�a<g�a<˄a<��a<b�a<9�a<a�a<�a<6�a<��a<��a<Ջa<�a<��a<I�a<��a<�a<�a<:�a<�a<9�a<ʓa<ϓa<3�a<��a<�a<��a<��a<�a<i�a<�a<��a<ĉa<׈a<Јa<�a<Éa<<�a<��a<��a<{�a<��a<��a<e�a<��a<A�a<?�a<v�a<�a<�a<��a<,�a<��a<|�a<-�a<C�a<B�a<��a<��a<q�a<9�a<��a<*�a<�a<��a<K�a<'�a<��a<@�a<��a<��a<đa<ȏa<]�a<&�a<3�a<�a<�a<Ɍa<�a<'�a<�a<��a<��a<1�a<Зa<�a<��a<K�a<s�a<��a< �a<��a<��a<!�a<��a<-�a<�a<�a<�a<2�a<��a<�a<%�a<R�a<��a<P�a<c�a<�a<n�a<��a<��a<J�a<J�a<4�a<Ƈa<<�a<^�a<�a<��a<a<��a<ȇa<I�a<��a<m�a<��a<Ύa<v�a<�a<ʏa<a<I�a<.�a<X�a<�a<�a<#�a<s�a<݈a<O�a<"�a<Їa<�a<��a<��a<��a<ۅa<!�a<s�a<��a<ta<O}a<�za<3xa<�ua<�sa<�qa<pa<Boa<�na<�na<hoa<pa<Pqa<�ra< ta<�ua<�va<�wa<hxa<�xa<�xa<�xa<
xa<6wa<cva<xua<�ta<.ta<�sa<�sa<�sa<�sa<�sa<Sta<kta<�ta<[ta<�sa<\sa<ra<�pa<�na<Oma<ka<Iia<Jga<�ea<�da<�ca<�ca<�ca<�da<�ea<aga<pia<Cka<�  �  �ma<poa<Tqa<�ra<�sa<�ta<)ua<Hua<-ua< ua<�ta<�ta<�ta<�ta<�ta<lua<va<�va<�wa<�xa<Vya<za<�za<�za<kza<�ya<#ya<�wa<�va<Nua<	ta<�ra<�qa<pqa<�qa<ra<sa<qta<lva<�xa<*{a<�}a<L�a<��a<�a<��a<,�a<W�a<7�a<��a<�a<T�a<��a<̋a<��a<x�a<�a<؍a<�a<��a<��a<�a<��a<��a<��a<��a<��a<�a<�a<��a<+�a<��a<�a<Ǌa<��a<�a<�a<=�a<�a<&�a<ʌa<��a<��a<ƒa<��a<��a<�a<-�a<�a<��a<Úa<��a<Y�a<�a<��a<R�a<�a< �a< �a<q�a<��a<s�a<��a<U�a<��a<�a<��a<�a</�a<�a<d�a<��a<Óa<�a<�a<��a<-�a<}�a<-�a<R�a<،a<�a<j�a<,�a<�a<��a<S�a<�a<��a<љa<L�a<|�a<<�a<��a<I�a<��a<$�a<y�a<�a<Ζa<��a<�a<6�a<r�a<��a<Ηa<��a<ėa<4�a<H�a<�a<��a<��a<��a<��a<u�a<s�a<��a<_�a<��a<2�a<B�a<��a<��a<�a<|�a<��a<��a<��a<�a<y�a<�a<�a<��a<ʎa<��a<�a<�a<�a<�a<H�a<��a<0�a<
�a<ׇa<��a<m�a<�a<��a< �a<�a<m�a<ׁa<�a<k}a<�za<gxa<�ua<�sa<�qa<Ypa<eoa<�na<�na<Soa<Apa<qa<�ra<Cta<�ua<�va<�wa<Txa<�xa<�xa<\xa<�wa<wa<Cva<�ua<�ta<ta<�sa<jsa<hsa<�sa<�sa<ta</ta<Pta<Tta<�sa<-sa<ra<�pa<oa<Zma<Rka<qia<�ga<fa<�da<da<�ca<da<�da<fa<�ga<�ia<�ka<�  �  �ma<�oa<]qa<�ra<�sa<|ta<�ta<�ta<ua<�ta<Lta<ta<�sa<ta<6ta<�ta<Mua<=va<wa<6xa<.ya<�ya<qza<zza<xza<�ya<;ya<4xa<wa<�ua<mta<�sa<�ra<Kra<Kra<�ra<�sa<ua<-wa<8ya<�{a<~a<~�a<Ђa<�a<��a<�a<4�a<��a<V�a<ڊa<��a<ߊa<��a<P�a<��a<^�a<8�a<�a<D�a<H�a<��a<��a<O�a<Փa<͓a<��a<�a<�a<ߐa<��a<�a<��a<��a<V�a<��a<��a<��a<ъa<Ћa<��a<�a<!�a<�a<��a<��a< �a<E�a<�a<~�a<o�a<[�a<�a<T�a<��a<��a<n�a<@�a<}�a<��a<3�a<ʙa<^�a<4�a<\�a<��a<��a<�a<C�a<�a<��a<��a<:�a<M�a<��a<>�a<�a<T�a<��a<"�a<��a<��a<�a<��a<Z�a<��a<��a<��a<�a<˙a<(�a<Q�a<�a<��a<a<�a<]�a<��a<t�a<�a<'�a<�a<y�a<a<I�a<��a<��a<��a<�a<U�a<'�a<��a<�a<��a<��a<ًa<,�a<i�a<;�a<[�a<̅a<&�a<f�a<��a<��a<�a<e�a<��a<��a<�a<��a<��a<ŏa<Y�a<��a<ҍa<h�a<e�a<@�a<]�a<��a<�a<��a<1�a<,�a<��a<:�a<؆a<~�a<�a<��a<��a<ԁa<�a<�}a<I{a<�xa<va<�ta<ora<?qa<pa<�oa<�oa<�oa<qa<�qa<Asa<�ta<�ua<�va<�wa<lxa<�xa<�xa<	xa<{wa<�va<�ua<�ta<�sa<osa<�ra<�ra<�ra<�ra<(sa<xsa<ta<�sa<"ta<�sa<sa</ra<�pa<Woa<�ma<�ka<�ia<1ha<�fa<sea<�da<gda<�da<�ea<�fa<Mha<�ia<�ka<�  �  zna<4pa<�qa<�ra<�sa<8ta<yta<ita<7ta<�sa<�sa<)sa<sa<sa< sa<�sa<gta<`ua<]va<jwa<gxa<Aya<�ya<Vza<�za<za<�ya<�xa<�wa<�va<Kua<bta<�sa<2sa<Nsa<�sa<�ta<!va<�wa<za<l|a<�~a<�a<K�a< �a<��a<�a<шa<{�a<��a<�a<�a<�a<�a<m�a<��a<F�a<N�a<#�a<z�a<��a<͐a<ܑa<Ғa<d�a<Гa<��a<#�a<��a<q�a<2�a<�a<m�a<Z�a<e�a<׊a<��a<��a<��a<׌a<Y�a<��a<�a<ēa<��a<�a<2�a<T�a<Йa<��a<�a<��a<+�a<��a<$�a<��a<j�a<)�a<i�a<Зa<D�a< �a<��a<U�a<ךa<8�a<7�a<�a<P�a<V�a<%�a<��a<�a<'�a<{�a<�a<�a<>�a<�a<�a<��a<��a<�a<f�a<�a<��a<�a<<�a<�a<ԙa<�a<˙a<\�a<ǘa<��a<>�a<s�a<ԕa<]�a<��a<�a<1�a<��a<�a<|�a<ޖa<�a<!�a<��a<a�a<9�a<�a<o�a<��a<��a<��a<��a<i�a<!�a<^�a<�a<�a<m�a<S�a<_�a<��a<�a<O�a<k�a<�a<��a<Ǐa<a�a<܎a<�a<�a<��a<��a<O�a<y�a<|�a<چa<��a<B�a<a�a<I�a<P�a<3�a< �a<p�a<��a<��a<�a<O�a<+~a<�{a<�ya<Jwa<Qua<}sa<ra<!qa<�pa<�pa<qa<�qa<�ra<ta<Aua<ava<\wa<�wa<{xa<oxa<xa<�wa<�va<�ua<�ta<�sa<�ra<kra<�qa<�qa<�qa<�qa<_ra<�ra<0sa<wsa<�sa<rsa<)sa<<ra<"qa<�oa<4na<xla<�ja<�ha<�ga<ufa<�ea<�ea<�ea<�fa<�ga<ia<�ja<�la<�  �  oa<�pa<ra<�ra<�sa<�sa<ta<�sa<Jsa<�ra<Qra<�qa<�qa<�qa<�qa<=ra<sa<ta<<ua<rva<�wa<�xa<�ya<za<Nza<Pza<�ya<ya<Axa<Twa<}va<�ua<ua<�ta<�ta<Tua<va<�wa<8ya<?{a<k}a<wa<��a<��a<k�a<��a<Շa<��a<��a<�a<��a<�a<Ɉa<��a<�a<;�a<׉a<͊a<Ջa<$�a<��a<ݏa<�a<L�a<�a<��a<��a<��a<�a<�a<ߐa<Џa<��a<��a<׌a<4�a<9�a<s�a<�a<B�a<��a<-�a<Œa<c�a<�a<p�a<��a<!�a<��a<��a<j�a<Ƙa<5�a<��a<Ԗa<B�a<�a<a<�a<g�a<��a<ėa<��a<c�a<3�a<��a<�a<ۚa<d�a<a<w�a<�a<��a<B�a<��a<c�a<]�a<��a<}�a<u�a<	�a<�a<�a<��a<Ҕa<*�a<k�a<��a<B�a<��a<��a<`�a<ǘa<ڗa<�a<�a<"�a<r�a<ؓa<��a<��a<ۓa<I�a<�a<��a<��a<��a<Öa<��a<*�a<z�a<j�a<ɒa<;�a<��a<�a<$�a<ˊa<��a<ǈa<~�a<Z�a<�a<��a<��a<��a<��a<ōa<��a<o�a<��a<��a<�a<Y�a<7�a<��a<��a<O�a<�a<��a<�a<k�a<%�a<�a<�a<@�a<`�a<r�a<{�a<"�a<��a<z�a<L�a<��a<�~a<�|a<�za<�xa<�va<�ta<vsa<�ra<ra<�qa<ora<�ra<�sa<�ta<�ua<�va<�wa<7xa<Ixa<.xa<�wa<wa<�ua<�ta<�sa<�ra<�qa<�pa<fpa<6pa<^pa<�pa<#qa<�qa<>ra<�ra<,sa<*sa<�ra<Pra<�qa<(pa<�na<2ma<�ka<0ja<�ha<�ga<4ga<+ga<=ga<�ga<ia<Kja<�ka<rma<�  �  	pa<9qa<Mra<sa<xsa<�sa<fsa<�ra<nra<�qa<�pa<dpa<pa<�oa<0pa<�pa<�qa<�ra<�sa<Oua<�va<�wa<�xa<�ya<Cza<~za<Aza<�ya<Jya<ixa<�wa<�va<eva<Eva<Vva<�va<�wa<ya<�za<�|a<v~a<��a<n�a<�a<��a<Ɔa<��a<�a<0�a<(�a<�a<��a<]�a<L�a<N�a<��a<E�a<0�a<j�a<��a<-�a<��a<@�a<y�a<��a<F�a<��a<̓a<Q�a<��a<�a<ِa<��a<�a<=�a<�a<ɍa<�a<Ǝa<��a<�a<l�a<ԓa<m�a<��a<��a<��a<�a<:�a<�a<��a<�a< �a<!�a<c�a<Ȕa<[�a<1�a<b�a<˔a<�a<\�a<c�a<��a<G�a<�a<��a<��a<��a<�a<�a<�a<Ėa<[�a<�a<˒a<�a<J�a<��a< �a<��a<X�a<l�a<��a<�a<-�a<�a<�a<g�a<y�a<F�a<��a<ڗa<��a<˕a<��a<��a<ڒa<Q�a<�a<�a<T�a<ؒa<��a<`�a<%�a<��a<.�a<J�a<�a<��a<��a<��a<C�a<��a<�a<��a<.�a<4�a<f�a<�a<�a<T�a<�a<�a<Ɍa<Ӎa<��a<?�a<��a<��a<I�a<��a<��a<W�a<�a<X�a<�a<��a<Z�a<|�a<كa<��a<��a<��a<��a<r�a<��a<��a<��a<4�a<��a<��a<�a<xa<�}a<�{a<�ya<�wa<Vva<4ua<;ta<�sa<�sa<�sa<[ta<5ua<�ua<�va<�wa<	xa<oxa<Fxa<�wa<7wa<va<ua<�sa<Zra<0qa<-pa<]oa<�na<�na<�na<(oa<�oa<}pa<`qa<�qa<wra<�ra<�ra<qra<�qa<�pa<�oa<Rna<�la<�ka<Nja<ria<�ha<�ha<�ha<�ia<fja<�ka<ma<�na<�  �  �pa<�qa<�ra<6sa<dsa<3sa<�ra<ra<Cqa<Gpa<�oa<�na<Sna<=na<Sna<oa<�oa<qa<�ra<�sa<�ua<wa<~xa<sya<>za<�za<�za<�za<za<�ya<�xa<�xa<xa<�wa<!xa<�xa<�ya<�za<T|a<�}a<�a<��a<1�a<˄a<�a<܆a<c�a<��a<��a<2�a<Æa<M�a<��a<��a<��a<�a<y�a<��a<��a<V�a<�a<��a<B�a<Ӑa<*�a<�a<Ǔa<��a<��a<��a<ߒa<�a<P�a<��a<��a<��a<��a<ԏa<r�a<M�a<��a<��a<�a<D�a<y�a<T�a<�a<"�a<��a<��a<Ǘa<ߖa<��a<Ӕa<�a<�a<��a<Y�a<��a<�a<�a<�a<�a<N�a<f�a<|�a<&�a<��a<��a<R�a<ԙa<Әa<̗a<��a<��a<|�a<��a<�a<��a<�a<A�a<�a<�a<ڕa<�a<�a<טa<D�a<��a<e�a<ߘa<*�a<�a<ӕa<n�a<U�a<�a<%�a<��a<*�a<Z�a<��a<X�a<3�a<�a<�a<�a<��a<��a<�a<Еa<5�a<X�a<�a<ȑa<_�a<'�a<ԍa<݌a<0�a<��a<ڋa<�a<��a<N�a<��a<Ύa<h�a<�a<�a<��a<�a<5�a<�a<a�a<��a<�a<��a<�a<��a<��a<�a<݁a<Ӂa<=�a<��a<�a<��a<�a<5�a<�a<��a<ła<��a<=�a<�~a<�|a<,{a<�ya<xa<�va<�ua<~ua<Yua<zua<va<~va<&wa<�wa<Zxa<�xa<�xa<Jxa<�wa<�va<bua< ta<ira<qa<�oa<pna<�ma<�la<�la<ma<�ma<fna<(oa<)pa<qa<�qa<ara<�ra<�ra<ra<�qa<ppa<Yoa<na<ma<�ka<ka<�ja<cja<�ja<(ka<la<9ma<Dna<�oa<�  �  �qa<�ra<sa<Hsa<Asa<�ra<ra<Hqa<,pa<oa<na<)ma<�la<qla<�la<<ma<*na<loa<qa<�ra<�ta<Jva<�wa<(ya<za<�za<,{a<0{a<�za<�za<Eza<�ya<�ya<�ya<�ya<gza<I{a<t|a<�}a<Da<	�a<��a<�a<I�a<'�a<Ԇa<;�a<	�a<Ɇa<V�a<��a<�a<R�a<�a<��a<�a<��a<҅a<�a<��a<��a<X�a<W�a<�a<��a<�a<��a</�a<w�a<0�a<�a<r�a<��a<�a<��a<X�a<O�a<��a<�a<��a<�a<�a<Q�a<5�a<�a<Øa<�a<�a<��a<�a<�a<��a<��a<f�a<5�a<]�a<�a<��a<Ґa<o�a<=�a<d�a<͔a<+�a<��a<��a<��a<l�a<��a<��a<X�a<��a<�a<�a<ߖa<��a<D�a<̔a<��a<��a<��a<��a<S�a<:�a<)�a<ǘa<c�a<��a<��a<B�a<|�a<m�a<;�a<��a<6�a<��a<p�a<�a<ǎa<q�a<��a<�a<��a<��a<Бa<	�a< �a<��a<��a<��a<�a<��a<�a<��a<�a<��a<~�a<v�a<��a<��a<��a<��a<a<�a<��a<\�a<ُa<#�a<j�a<+�a<��a<��a<��a<+�a<��a<��a<Æa<ׄa<;�a<�a<�a<S�a<*�a<"�a<��a<C�a<ہa<��a<;�a<��a<كa<��a<��a<3�a<�a<�a<;~a<x|a<{a<�ya<�xa<�wa<Dwa<wa<'wa<`wa<�wa<rxa<�xa<�xa<ya<�xa<0xa<[wa<	va<�ta<sa<:qa<�oa<na<�la<�ka<Gka<ka<gka<�ka<�la<�ma<oa<<pa<$qa<�qa<}ra<�ra<vra<ra<=qa<vpa<noa<_na<�ma<�la<ela<?la<mla<�la<�ma<�na<�oa<�pa<�  �  �ra<!sa<esa<asa<sa<�ra<dqa<Cpa<oa<�ma<�la<�ka<ka<�ja<ka<�ka<�la<na<�oa<�qa<vsa<Xua<+wa<�xa< za<�za<�{a<�{a<�{a<�{a<�{a<L{a<"{a<={a<r{a<�{a<�|a<�}a<6a<��a<�a<h�a<̈́a<΅a<}�a<ӆa<��a<��a<��a<J�a<��a<��a<�a<��a<A�a<��a<.�a<�a<��a<8�a<A�a<Q�a<J�a<9�a<$�a<��a<��a<��a<�a<�a<��a<k�a<��a<|�a<�a<�a<�a<+�a<��a<j�a<U�a<V�a<5�a<�a<Ԙa<,�a<K�a<�a<r�a<c�a<�a<Ȕa<��a<�a<ΐa<�a<+�a<�a<1�a<ȏa<ؐa<�a<��a<�a<��a<��a<g�a<A�a<��a<�a<�a<��a<a<�a<@�a<p�a<іa<P�a<�a<,�a<��a<�a<��a<r�a<�a<��a<�a<�a<��a<�a<;�a<��a<6�a<��a<�a<`�a<
�a<�a< �a<��a<یa<o�a<=�a<]�a<��a<�a<,�a<[�a<m�a<ەa<%�a< �a<��a<�a<�a<��a<�a<�a<,�a<��a<#�a<�a<5�a<��a<�a<j�a<��a<�a<�a<��a<��a<��a<F�a<^�a<z�a<|�a<}�a<s�a<؁a<N�a<Xa<�~a<m~a<�~a<a<�a<Ԁa<��a<g�a</�a<��a<��a<J�a<��a<��a<x�a<3a<�}a<r|a<-{a</za<Sya<�xa<�xa<�xa<�xa<ya<Vya<�ya<�ya<uya<ya<xa<wa<ua<�sa<�qa<-pa<Lna<�la<Oka<.ja<�ia<}ia<�ia<�ja<gka<�la<�ma<4oa<`pa<�qa<Qra<�ra<�ra<�ra<&ra<Oqa<�pa<�oa<�na<[na<�ma<�ma<�ma<sna<oa<�oa<�pa<�qa<�  �  sa<�sa<�sa<�sa<�ra<"ra<qa<�oa<Ena<�la<�ka<sja<�ia<jia<�ia<0ja<0ka<�la<�na<�pa<�ra<�ta<�va<zxa<�ya<7{a<�{a<g|a<�|a<�|a<�|a<�|a<n|a<�|a<�|a<b}a<[~a<9a<��a<��a<	�a<;�a<P�a<�a<��a<�a<��a<Z�a<��a<��a<��a<��a<Ła<#�a<ހa<�a<��a<��a<1�a<�a<�a<l�a<��a<Ȏa<ΐa<H�a<͓a<��a<<�a<��a<��a<Y�a<�a<Ҕa<e�a<q�a<O�a<��a<8�a<��a<��a<W�a<)�a<˘a<X�a<y�a<��a<�a<�a<�a<��a<�a<x�a<ېa<��a<p�a<Ӎa<��a<ˍa<_�a<|�a<�a<q�a<B�a<��a<��a<��a<�a<��a<>�a<Q�a<�a<��a<�a<f�a<Ęa<)�a<ؗa<��a<��a<�a<X�a<�a<h�a<�a<B�a<m�a<C�a<�a<�a<͗a<`�a<��a<Ԓa<�a<9�a<��a<w�a<��a<V�a<��a<��a<��a<'�a<��a<1�a<��a<
�a<�a<ϕa<`�a<K�a< �a<��a<ٔa<��a<)�a<7�a<��a<��a<��a<��a<��a<ܐa<�a<\�a<��a<��a<@�a<��a<�a<e�a<�a<�a<ֈa<��a<C�a<K�a<m�a<�~a<�}a<;}a<}a<P}a<�}a<�~a<�a<��a<��a<قa<6�a<��a<��a<��a<H�a<?�a<"�a<�~a<�}a<}|a<�{a<�za<Fza<za<�ya<za< za<Jza<Iza<9za<�ya<7ya<xa<�va<-ua<Bsa<5qa<$oa<ma<`ka<�ia<�ha<0ha<ha<Wha<&ia<Cja<�ka<ma<�na<pa<9qa<ra<�ra<	sa<sa<�ra<1ra<�qa<�pa<Epa<�oa<poa</oa<yoa<�oa<dpa<qa<�qa<�ra<�  �  �sa<ta<�sa<�sa<�ra<�qa<�pa<oa<�ma<�ka<�ja<�ia<�ha<qha<Zha<Iia<.ja<�ka<�ma<�oa<ra<;ta<Yva<Exa<�ya<*{a<,|a<�|a<}a<�}a<E}a<U}a<^}a<�}a<�}a<{~a<Xa<&�a<Z�a<n�a<�a<�a<҅a<��a<̆a<�a<��a<��a<�a<��a<ׂa<��a<��a<�a<�a<�a<��a<܁a< �a<B�a<<�a<��a<��a<7�a<_�a<4�a<��a<��a<��a<�a<-�a<@�a<��a<��a<T�a<a�a<h�a<��a<�a<��a<g�a<�a<�a<]�a<ԙa<֙a<t�a<�a<�a<��a<�a<j�a<��a<�a<��a<j�a<�a<d�a<̌a<s�a<��a<�a<��a<��a<Z�a<�a<��a<�a<�a<l�a<՛a<��a<q�a<ؚa<%�a<��a<�a<�a<��a<ʘa<јa<=�a<��a</�a<��a<ǚa<�a<��a<�a<ؘa<��a<�a<�a<�a<�a<d�a<Ȍa<~�a<Ɗa<.�a<��a<��a< �a<Z�a<̎a<��a<�a<��a<̔a<ŕa<S�a<��a<��a<�a<��a<��a<�a<'�a<~�a<�a<��a<��a<t�a<��a<Ƒa<9�a<;�a<
�a<��a<ѐa<֏a<S�a<��a<i�a<.�a<хa<p�a<�a<aa<~a<�|a<&|a<4|a<?|a<)}a<�}a<a<P�a<e�a<j�a<"�a<��a<��a<p�a<ǂa<�a<	�a<�a<�~a<l}a<�|a<�{a<Y{a<{a<�za<�za<�za<3{a<�za<�za<za<+ya<xa<�va<�ta<�ra<�pa<Mna<Fla<�ja<�ha<�ga<
ga<ga<lga<*ha<nia<�ja<_la<�ma<�oa<�pa<ra<�ra<7sa<�sa<4sa<�ra<[ra<�qa<%qa<�pa<�pa<Dpa<�pa<�pa<Iqa<�qa<�ra<_sa<�  �  �sa<5ta<	ta<�sa<�ra<�qa<Lpa<�na<ma<�ka<�ia<�ha<�ga<�ga<�ga<nha<{ia<*ka<ma<Zoa<�qa<ta<va<Dxa<�ya<A{a<N|a<}a<j}a<�}a<�}a<�}a<-~a<G~a<�~a<8a<�a<��a<�a<'�a<3�a<$�a< �a<��a<��a<׆a<��a<υa<ӄa<��a<f�a<B�a<5�a<na<a<Pa<�a<��a<y�a<z�a<��a<&�a<��a<	�a<.�a<6�a<��a<�a<ҕa<T�a<h�a<|�a<r�a<P�a<,�a<��a<$�a<e�a<˖a<y�a<�a<��a<6�a<��a<�a<��a<��a<͘a<�a<V�a<Ӕa<��a<9�a<y�a<��a<��a<�a<΋a<�a<��a<эa<X�a<0�a<�a<�a<ܖa<��a<�a<�a<��a<��a<�a<��a<E�a<Ԛa<c�a<ܙa<��a<X�a<b�a<��a<�a<U�a<��a<�a<#�a<�a<��a<�a<Θa<y�a<��a<a<��a<��a<��a<�a<��a<��a<��a<��a<B�a<c�a<��a<i�a<�a<בa<J�a<˔a<��a<j�a<��a<Жa<c�a<ݕa<M�a<��a<��a<6�a<��a<c�a</�a<H�a<g�a<�a<��a<m�a<X�a<ޑa<�a<��a<P�a<a�a<6�a<Շa<_�a<�a<��a<�~a<*}a< |a<{a<M{a<�{a<b|a<r}a<�~a<�a<6�a<9�a<#�a<y�a<��a<��a<�a<%�a<E�a<M�a<Ea<D~a<>}a<�|a<|a<�{a<�{a<�{a<|{a<W{a<%{a<�za<Bza<Qya<�wa<�va<rta<pra< pa<�ma<�ka<�ia<&ha<ga<tfa<Nfa<�fa<{ga<�ha<Kja<�ka<�ma<Goa<�pa<�qa<�ra<dsa<�sa<�sa<"sa<�ra<Sra<�qa<eqa<qa<qa<'qa<zqa<ra<�ra<sa<�sa<�  �  ua<�ta<ua<�ta< ta<_sa<@ra<3qa<�oa<�na<�ma<�la<ula<"la<>la<�la<�ma<-oa<�pa<�ra<0ta<6va<�wa<�ya<�za<H|a<}a<�}a<h~a<�~a<�~a<a<Qa<�a<�a<��a<<�a</�a<�a<�a<�a<�a<ֆa<�a<��a<��a<��a<�a<|�a<��a<�a<I�a<��a<a�a<�a<Z�a<�a<��a<`�a<��a<��a<��a<q�a<|�a<>�a<�a<�a<a�a<ٕa<��a<�a<�a<�a<ʖa<�a<іa<�a<P�a<��a<0�a<��a<E�a<��a<2�a<G�a<+�a<�a<Y�a<Әa<��a<z�a<�a<ϓa<��a<o�a<��a<��a<ɏa<�a<��a<��a<��a<�a<N�a<�a<R�a<��a<��a<q�a<�a<�a<e�a<'�a<��a<y�a<�a<��a<x�a<~�a<_�a<z�a<��a<��a<b�a<y�a<��a<F�a<�a<~�a<{�a<��a<�a<��a<ۓa<~�a<ސa<ŏa<Ǝa<��a<��a<��a<J�a<�a<ُa<�a<-�a<��a<��a<̕a<E�a<��a<�a<�a<�a<k�a<�a<<�a<��a<�a<��a<v�a<�a<�a<��a<�a<�a<��a<��a<�a<��a<F�a<�a<y�a<��a<��a<Ƈa<��a<��a<��a<(�a<6�a<�a<Ua<�a<�a<��a<I�a<
�a<�a<��a<6�a<K�a<��a<��a<ƃa<�a<)�a<E�a<9�a<ya<�~a<~a<y}a<}a<�|a<�|a<�|a<\|a<3|a<�{a<�za<Xza<ya<�wa<:va<�ta<�ra< qa<Coa<�ma<�la<�ka<�ja<�ja<$ka<�ka<mla<�ma<�na<pa<Iqa<pra<;sa<�sa<jta<Xta<�ta<Cta<ta<�sa<sa<�ra<�ra<�ra<�ra<�ra<Nsa<�sa<Wta<�ta<�  �  �ta<ua<ua<�ta<ta<Rsa<Hra<Fqa<pa<�na<�ma<ma<ula<bla<�la< ma<�ma<Poa<�pa<�ra<ota<Iva<�wa<�ya<�za<>|a<$}a<�}a<~a<x~a<�~a<�~a<+a<sa<�a<f�a< �a<��a<�a<�a<�a<��a<��a<A�a<��a<��a<��a< �a<��a<݅a<�a<b�a<��a<Y�a<;�a<��a<!�a<�a<W�a<�a<ǉa<��a<��a<��a<H�a<�a< �a<M�a<��a<p�a<��a<Ȗa<ʖa<��a<��a<��a<ۖa<�a<��a<�a<��a<�a<��a<��a<A�a<F�a<�a<l�a<��a<��a<��a<?�a<��a<��a<��a<��a<7�a<�a<@�a<��a<��a<��a<'�a<��a<�a<X�a<��a<��a<v�a<�a<C�a<.�a<�a<a<Z�a<��a<��a<Z�a<0�a<=�a<^�a<��a<ߚa<+�a<E�a<c�a<h�a<�a<{�a<��a<y�a<�a<��a<�a<��a<�a<ُa<ǎa<9�a<ڍa<��a<D�a<�a<	�a<C�a<l�a<��a<��a<��a<_�a<��a<%�a<�a<��a<>�a<��a<#�a<��a<��a<��a<+�a<��a<�a<�a<�a<�a<��a<��a<�a<o�a<N�a<�a<��a<ˋa<�a<��a<�a<2�a<��a<L�a<i�a<�a<�a<�a<�a<��a<{�a<B�a<�a<��a<*�a<T�a<u�a<�a<��a<��a<�a<�a<*�a<Ia<w~a<�}a<D}a<�|a<�|a<�|a<a|a<1|a<�{a<�{a<{a<Lza<ya<�wa<Ava<�ta<�ra</qa<loa<�ma<�la<�ka<1ka<ka</ka<�ka<�la<�ma<�na<1pa<Pqa<gra<Jsa<�sa<gta<�ta<Yta<ta<�sa<isa<sa<�ra<�ra<kra<�ra<�ra<6sa<�sa<ta<pta<�  �  �ta<�ta<�ta<�ta<7ta<wsa<�ra<qqa<`pa<:oa<Ona<�ma<�la<�la<�la<�ma<una<�oa<7qa<�ra<�ta<rva<=xa<�ya<!{a<|a<�|a<�}a<�}a<a~a<S~a<�~a<�~a<�~a<Xa<�a<��a<p�a<��a<~�a<��a<��a<h�a<�a<k�a<��a<��a<I�a<��a<�a<l�a<��a<G�a<҃a<كa<	�a<��a<��a<φa<z�a<�a<�a<ٍa<��a<{�a<��a<A�a<�a<ٕa<;�a<y�a<��a<V�a<Y�a<#�a<D�a<N�a<��a<�a<m�a< �a<��a<q�a<��a<�a<�a<�a<��a<Иa<�a<��a<w�a<B�a<�a<�a<)�a<Аa<i�a<Đa<;�a<�a<6�a<j�a<��a<4�a<��a<ęa<Ěa<o�a<ƛa<�a<��a<ۛa<j�a<�a<��a<�a<�a<��a<��a<ԙa<�a<l�a<̚a<3�a<.�a<<�a<Ԛa<g�a<��a<��a<_�a<��a<m�a<ߒa<��a<Y�a<N�a<Ďa<>�a<��a<��a<��a<e�a<��a<��a<Гa<��a<ѕa<��a<Жa<�a<�a<{�a<'�a<Q�a<��a<��a<w�a< �a<��a<��a<\�a<��a<z�a<��a<��a<Q�a<�a<+�a<a�a<$�a<��a<��a<�a<I�a<X�a<��a<�a<�a<�a<>�a<"�a<�a<��a<��a<Áa<r�a<3�a<؃a<=�a<u�a<:�a<��a<`�a<��a<܁a<��a<�a<�~a<~a<>}a<�|a<l|a<|a<|a<�{a<|a<�{a<x{a<�za<za<Cya<�wa<�va<�ta<sa<sqa<�oa<ona<ma<Zla<�ka<�ka<�ka<Kla< ma<na<Goa<apa<�qa<�ra<bsa<�sa< ta<Yta<$ta<�sa<}sa<�ra<�ra<)ra<ra<�qa<ra<Hra<�ra<1sa<�sa<]ta<�  �  8ta<�ta<�ta<�ta<,ta<�sa<�ra<�qa<�pa<�oa<�na<=na<�ma<�ma<�ma<nna<Hoa<{pa<�qa<�sa<9ua<�va<~xa<�ya<{a<|a<�|a<>}a<�}a<�}a<�}a<�}a<�}a<1~a<�~a< a<�a<a<߁a<܂a<��a< �a<�a<҆a<l�a<��a<��a<��a<#�a<��a<�a<_�a<��a<��a<��a<�a<v�a<_�a<��a<�a<Ŋa<��a<a�a<"�a<��a<�a<;�a<�a<��a<�a< �a<ݕa<��a<��a<u�a<q�a<��a<Εa<?�a<Ŗa<��a<�a<��a<R�a<��a<�a<�a<��a<�a<(�a<"�a<�a<�a<��a<��a<��a<��a<N�a<��a< �a<ʒa<Γa<�a<p�a<��a<�a<��a<��a<m�a<Ǜa<ěa<��a<@�a<��a<I�a<љa<^�a<�a<�a<�a<�a<k�a<әa<'�a<��a<Ӛa<�a<њa<g�a<��a<Øa<��a<_�a<��a<��a<$�a<�a<�a<��a<'�a<B�a<��a<;�a<�a<4�a<7�a<D�a<9�a<�a<s�a<Жa<ϖa<��a<�a<m�a<��a<�a<O�a<��a<3�a<�a<��a<��a<֑a<ؑa<��a<�a<��a<��a<-�a<]�a<)�a<�a<Z�a<��a<�a<�a<Y�a<׃a<��a<��a<�a<Ԁa<ڀa</�a<��a<f�a<��a<��a<�a<I�a<o�a<8�a<��a<�a<.�a<�a<�a<a<	~a</}a<|a<�{a<�{a<s{a<z{a<R{a<T{a<S{a<{a<�za<za<2ya<xa<�va<Bua<�sa<ra<opa<oa<�ma<ma<{la<`la<�la<�la<�ma<�na<�oa<�pa<�qa<�ra<]sa<�sa< ta<ta<�sa<\sa<�ra<Yra<�qa<xqa<8qa<(qa<Aqa<�qa<ra<�ra<sa<�sa<�  �  �sa< ta<�ta<wta<Mta<�sa</sa<�ra<xqa<�pa<�oa<Hoa<�na<�na<�na<coa<^pa<{qa<�ra<Gta<�ua<vwa<�xa<*za<%{a<�{a<�|a<�|a<}a<�|a<}a<�|a<�|a<'}a<{}a<'~a<�~a<�a<ɀa<"�a<P�a<��a<��a<z�a<A�a<��a<�a<ׇa<��a<#�a<��a<5�a<Ʌa<��a<��a<�a<��a<^�a<��a<�a<��a<;�a<��a<��a<�a<E�a<'�a<�a<@�a<v�a<m�a<3�a<�a<��a<{�a<a�a<��a<Ôa<.�a<Õa<|�a<b�a<�a<̘a<G�a<��a<��a<��a<7�a<l�a<��a<��a<��a<��a<��a<�a<}�a<n�a<��a<�a<ݓa<��a<�a<��a<K�a<J�a<F�a<�a<L�a<��a<]�a<0�a<��a<�a<w�a<Ęa<i�a<��a<�a<ڗa<#�a<d�a<�a<~�a<ݙa<a�a<z�a<��a<B�a<șa<�a<��a<�a<��a<Y�a<�a<�a<,�a<�a<J�a<8�a<��a<:�a<��a<ߒa<ȓa<Քa<}�a<>�a<��a<��a<��a<�a<��a<��a<�a<�a<L�a<��a<#�a<�a<��a<��a<��a<�a<K�a<w�a<��a<Q�a<�a<A�a<f�a<6�a<ˌa</�a<r�a<�a<C�a<��a<��a<Âa<*�a<Ӂa<��a<�a<��a<��a<��a<�a<b�a<��a<[�a<�a<d�a<��a<��a<o�a<Xa<~a<}a< |a<�{a<�za<�za<qza<uza<�za<�za<�za<�za<nza<�ya<<ya<Zxa<wa<�ua<<ta<�ra<Tqa<
pa<oa<na<�ma<`ma<�ma<na<�na<�oa<`pa<xqa<Bra<sa<�sa<�sa<�sa<�sa<\sa<�ra<(ra<�qa<�pa<�pa<&pa<.pa<0pa<�pa<�pa<�qa<sra<sa<�  �  sa<�sa<6ta<ota<jta<ta<�sa<sa<Qra<�qa<�pa<Opa<pa<�oa<pa<�pa<zqa<�ra<�sa<#ua<�va<xa<5ya<Kza<={a<�{a<;|a<`|a<c|a<E|a<|a<�{a<�{a<�{a<D|a<�|a<�}a<�~a<�a<�a<m�a<ڃa<�a<*�a<�a<��a<	�a<�a<�a<�a<��a<,�a<ֆa<��a<Іa<�a<��a<��a<��a<�a<��a<&�a<��a<"�a<V�a<k�a<<�a<��a<�a<�a<��a<T�a<��a<��a<d�a<5�a<M�a<��a<�a<��a<x�a<X�a<D�a<�a<͘a<R�a<��a<��a<U�a<֘a<@�a<g�a<o�a<��a<��a<-�a<ȓa<��a<˓a<>�a<�a<Ǖa<Ζa<ٗa<�a<əa<v�a<�a<P�a<E�a<��a<��a<�a<%�a<m�a<��a<:�a<ʖa<��a<��a<��a<`�a<�a<��a<5�a<��a<�a<K�a<:�a<�a<A�a<~�a<��a<^�a<:�a<�a<�a<W�a<a<l�a<�a<Ǒa<@�a<��a<��a<��a<h�a<�a<_�a<��a<��a<>�a<��a<�a<�a<�a<�a<I�a<��a<�a<��a<u�a<��a<a<�a<h�a<ϐa<�a< �a<Ɛa<P�a<��a<x�a<I�a<�a<_�a<؈a<O�a<��a<�a<��a<[�a<�a<�a<#�a<��a<�a<W�a<��a<��a<��a<q�a<كa<�a<	�a<�a<�a<I~a<}a<�{a<�za<>za<�ya<mya<iya<rya<�ya<�ya<za<0za<za<�ya<Sya<xxa<twa<_va<ua<�sa<Xra<qa<pa<Roa<�na<�na<�na<oa<�oa<spa<@qa<ra<�ra<?sa<�sa<�sa<�sa<<sa<�ra<ra<8qa<}pa<�oa<Toa<�na<�na<�na<loa<�oa<�pa<zqa<`ra<�  �  _ra<Wsa<�sa<`ta<�ta<nta<9ta<�sa</sa<ra<ra<�qa<9qa<Eqa<jqa< ra<�ra<�sa<�ta<va<iwa<�xa<�ya<�za<Q{a<�{a<�{a<�{a<�{a<g{a<{a<�za<�za<�za<{a<�{a<V|a<L}a<�~a<�a<��a<�a<j�a<ǅa<��a<��a<,�a<��a<��a<��a<X�a<�a<�a<�a<�a<�a<�a<�a<�a<A�a<��a<��a<i�a<��a<ʒa<��a<B�a<p�a<��a<S�a<��a<p�a<�a<�a<�a<�a<��a<I�a<��a<m�a<e�a<L�a<f�a<\�a<L�a< �a<p�a<��a<��a<Y�a<��a<(�a<T�a<��a<�a<P�a<�a<�a<#�a<w�a<�a<�a<��a<��a<y�a<T�a<ؚa<+�a<D�a<��a<��a<Йa<$�a<2�a<c�a<��a<�a<��a<F�a<m�a<��a<)�a<��a<��a<e�a<��a<��a<��a<*�a<�a<��a<�a<�a<<�a<$�a<>�a<K�a<��a<�a<Ēa<֒a<�a<t�a<�a<��a<h�a<�a<|�a<��a<��a<m�a<�a</�a<*�a<-�a<�a<�a<�a<5�a<��a<H�a<0�a<8�a<��a<�a<}�a<
�a<R�a<��a<z�a<R�a<��a<�a<؍a<��a<5�a<��a<~�a<)�a<$�a<[�a<��a<Y�a<)�a<V�a<v�a<��a<�a<$�a<&�a<ӄa<w�a<��a<��a<y�a<*�a<�~a<@}a<�{a<�za<�ya<�xa<rxa<%xa<xa<_xa<�xa<	ya<]ya<�ya<�ya<�ya<`ya<�xa<�wa<�va<�ua<�ta<esa<Fra<<qa<�pa<pa<�oa<�oa<Jpa<�pa<[qa<ra<�ra<Lsa<�sa<�sa<�sa<Psa<�ra<�qa<Aqa<Fpa<toa<�na<�ma<�ma<�ma<�ma<na<�na<�oa<�pa<�qa<�  �  �qa<�ra<�sa<@ta<�ta<�ta<�ta<\ta<ta<zsa<sa<�ra<�ra<�ra<�ra<9sa<�sa<�ta<�ua<wa<4xa<1ya<za<�za<[{a<�{a<�{a<[{a<{a<�za<za<�ya<rya<tya<�ya<-za<{a<-|a<r}a<a<��a<Z�a<�a<H�a<��a<��a<T�a<݈a<#�a<@�a<7�a<#�a<�a<8�a<\�a<ĉa<b�a<-�a<@�a<]�a<��a<ݏa<$�a<5�a<#�a<Ǔa<;�a<I�a<�a<Γa<L�a<��a<��a<K�a<�a<��a<��a<�a<z�a<>�a<8�a<d�a<��a<Ŗa<��a<��a<N�a<��a<ՙa<��a<]�a<�a<C�a<��a<�a<��a<R�a<L�a<`�a<Ȗa<Z�a<��a<��a<��a<=�a<ƚa<*�a<C�a<,�a<��a<�a<T�a<Q�a<C�a<K�a<_�a<��a<5�a<�a<�a<n�a<��a<a<��a<��a<x�a<'�a<��a<
�a<�a<�a<m�a<̘a<�a< �a<E�a<��a<ߔa<Y�a<�a<�a<K�a<��a<�a<��a<3�a<��a<ۖa<�a<Ėa<M�a<��a<��a<��a<V�a<�a<�a<Ўa<��a<U�a<�a<�a<�a<h�a<	�a<��a<N�a<֏a<�a<L�a<H�a<؏a<<�a<Z�a<K�a<�a<ϊa<��a<}�a<m�a<��a<
�a<��a<��a<r�a<��a<��a<��a<��a<�a<�a<p�a<r�a<@�a<�a<za<�}a<K|a<�za<yya<hxa<�wa<wa<�va<�va<2wa<�wa<3xa<�xa<"ya<]ya<�ya<aya<�xa<Zxa<|wa<�va<rua<ita<isa<�ra<�qa<xqa<4qa<Hqa<�qa<�qa<]ra<�ra<jsa<�sa<�sa<�sa<�sa<sa<Tra<�qa<npa<Xoa<\na<sma<�la<_la<)la<gla<�la<�ma<�na<�oa<�pa<�  �  Eqa<Mra<isa<$ta<�ta<ua<ua<ua<�ta<xta<ta<�sa<�sa<�sa<ta<kta<*ua<�ua<�va<�wa<�xa<�ya<yza<{a<R{a<r{a<Q{a<�za<eza<�ya</ya<�xa<lxa<@xa<pxa< ya<�ya<{a<n|a<
~a<�a<��a<`�a<�a<m�a<��a<��a<.�a<��a<�a< �a<0�a<�a<C�a<��a<��a<��a<Y�a<S�a<^�a<��a<��a<ؑa<Òa<t�a<��a<$�a<$�a<Ɠa<F�a<��a<��a<��a<F�a<ݏa<d�a<l�a<��a<B�a<7�a<)�a<p�a<��a<�a<D�a<W�a<&�a<��a<�a<�a<��a<��a<'�a<��a<�a<Зa<��a<��a<��a<��a<^�a<�a<��a<=�a<�a<6�a<y�a<_�a<�a<��a<��a<��a<|�a<f�a<L�a<[�a<��a<�a<ϒa<͒a<E�a<�a<��a<��a<��a<ߗa<��a<~�a<�a<(�a<7�a<ڙa<|�a<��a<�a<Q�a<��a<�a<��a<n�a<B�a<x�a<��a< �a<��a<ؖa<:�a<6�a<1�a<��a<+�a<T�a<(�a<�a<s�a<.�a<Ўa<ʍa<ƌa<�a<ċa<��a<�a<e�a<�a<��a<�a<H�a<��a<-�a<0�a<�a<��a<ێa<��a<݌a<܋a<��a<��a<��a<؇a<H�a<φa<��a<r�a<��a<u�a<q�a<;�a<Ѕa<@�a<Y�a<N�a<�a<l�a<�~a<�|a<K{a<�ya<qxa<#wa<]va<�ua<�ua<�ua<"va<�va<Gwa<	xa<�xa<"ya<_ya<Uya<7ya<�xa<xa<;wa<Vva<qua<fta<�sa<sa<�ra<ira<tra<�ra<�ra<asa<�sa<ta<.ta<Ata<�sa<�sa<�ra<�qa<�pa<�oa<{na<^ma<nla<�ka<ka<ka<$ka<�ka<�la<�ma<�na<�oa<�  �  �pa<�qa<sa<ta<�ta<Jua<vua<�ua<Vua<ua<�ta<�ta<�ta<�ta<ua<�ua< va<�va<�wa<�xa<�ya<Iza<�za<R{a<r{a<A{a<�za<~za<�ya<"ya<exa<�wa<Vwa<5wa<nwa<�wa<�xa<�ya<~{a<'}a<#a<�a<؂a<��a<$�a<��a<��a<�a<�a<~�a<��a<ӊa<%�a<B�a<��a<�a<��a<h�a<N�a<k�a<Q�a<a�a<h�a<2�a<ɓa<#�a<1�a<�a<x�a<ǒa<�a<�a<�a<X�a<��a<f�a<\�a<��a<9�a<�a<A�a<��a<�a<t�a<֖a<�a<�a<əa<C�a<i�a<o�a<8�a<ҙa<s�a<+�a<ɘa<��a<��a<��a<��a<`�a<��a<b�a<�a<b�a<��a<��a<��a<��a<>�a<U�a<.�a<�a<��a<]�a<W�a<�a<��a<��a<Ցa<3�a<�a<ʓa<�a<&�a<M�a<W�a<-�a<Йa<M�a<q�a<D�a<�a<d�a<Řa<9�a<��a<	�a<��a<g�a<W�a<o�a<��a<�a<3�a<��a<��a<��a<g�a<ۖa<��a< �a<Ǔa<Y�a<�a<c�a<�a<��a<��a<�a<��a<��a<�a<t�a<"�a<�a<�a<��a<u�a<�a<.�a<,�a<ޏa<J�a<��a<��a<�a<��a<��a<��a<�a<K�a<݇a<��a<��a<9�a< �a<�a<��a<&�a<h�a<e�a<�a<��a<�a<~a<V|a<lza<�xa<Mwa<%va<Mua<�ta<�ta<�ta<;ua<�ua<�va<uwa<9xa<�xa<&ya<sya<dya<ya<�xa<�wa<wa<1va<}ua<�ta<"ta<�sa<{sa<xsa<�sa<�sa<ta<Qta<�ta<�ta<�ta<%ta<nsa<�ra<�qa<Zpa<oa<�ma<nla<kka<�ja<$ja<�ia<,ja<�ja<�ka<�la<�ma<Roa<�  �  8pa<�qa<�ra<ta<�ta<Rua<�ua<�ua<va<�ua<�ua<sua<nua<�ua<�ua<Uva<�va<�wa<Xxa<Fya<za<�za<0{a<Q{a<s{a<D{a<�za<&za<Pya<�xa<�wa<"wa<�va<tva<�va<�va<xa<,ya<�za<w|a<z~a<j�a<m�a<c�a<�a<��a<��a<��a<o�a<�a<o�a<v�a<ǋa<�a<`�a<Ȍa<c�a<8�a<��a<�a<��a<$�a<ܒa<��a<�a<%�a<9�a<ѓa<<�a<^�a<b�a<r�a<e�a<��a<�a<��a<z�a<ٍa<�a<_�a<��a<�a<��a<��a<v�a<ɗa<�a<ʙa<B�a<��a<Ěa<��a<��a<�a<ݙa<w�a<o�a<G�a<x�a<��a<
�a<��a<�a<��a<śa< �a<̛a<��a<�a<�a<�a<��a<e�a<�a<��a<��a<��a<=�a<��a<�a<d�a<<�a<+�a<N�a<��a<Җa<�a<�a<ޙa<M�a<y�a<��a<N�a<�a<i�a<јa<=�a<a<r�a<�a<,�a<�a<c�a<��a<��a<�a<�a<�a<g�a<ܖa<��a<ʔa<o�a<ۑa<W�a<��a<S�a<��a<��a<K�a<Éa<�a<�a<Ίa<r�a<t�a<^�a<U�a<9�a<ʏa<<�a<0�a<�a<��a<��a<L�a<"�a<@�a<1�a<q�a<��a<�a<��a<>�a<'�a<܇a<�a<u�a<�a<c�a<k�a<m�a<��a<a�a<�a<�}a<�{a<�ya<%xa<�va<rua<jta<ta<�sa<ta<�ta<7ua<#va<�va<�wa<�xa<$ya<tya<cya<Xya<�xa<exa<�wa<�va</va<bua<�ta<sta<Kta<5ta<<ta<xta<�ta<ua<�ta<�ta<�ta<%ta<�sa<zra<Sqa<�oa<�na<ma<�ka<�ja<�ia<hia<�ha<mia<�ia<�ja<�ka<Dma<�na<�  �  pa<jqa<�ra<�sa<�ta<�ua<�ua<va<va<%va<va<�ua<�ua<va<Qva<�va<Zwa<xa<�xa<�ya<#za<�za<V{a<�{a<u{a<.{a<�za<�ya<ya<:xa<mwa<�va<!va<�ua<"va<�va<}wa<�xa<Qza<%|a<5~a<5�a<G�a<�a<�a<n�a<ވa<׉a<��a<
�a<��a<�a<.�a<��a<݌a<S�a<�a<��a<��a<v�a<h�a<I�a<��a<��a<(�a<]�a<�a<��a<�a<:�a<0�a<-�a<�a<)�a<v�a<�a<	�a<[�a<�a<�a<�a<��a<.�a<a<F�a<��a<ۘa<��a<��a<ޚa<��a<Ϛa<˚a<��a<D�a<�a<ݙa<әa<��a<9�a<��a<��a<l�a<��a<�a<-�a<�a<��a<�a<�a<Øa<��a<�a<Ĕa<V�a<,�a<,�a<��a<]�a<��a<ސa<��a<a<�a<O�a<��a<ėa<�a<��a<f�a<��a<ɚa<��a<)�a<˙a<B�a<Ęa<K�a<�a<��a<��a<��a<՗a< �a<3�a<#�a<8�a<�a<��a<ޖa<�a<��a<2�a<��a< �a<k�a<όa<�a<g�a<ɉa<\�a<W�a<��a<G�a< �a</�a<)�a</�a<�a<��a<�a<a�a<6�a<ԏa<�a<j�a<��a<��a<ɋa<�a</�a<��a<&�a<Ԉa<��a<P�a<�a<��a<4�a<��a<��a<H�a<�a<'�a<`a<^}a<j{a<mya<�wa<
va<�ta<�sa<�sa<Msa<�sa<ta<�ta<�ua<�va<�wa<mxa<ya<kya<�ya<{ya<ya<sxa<�wa<Ewa<�va<�ua<eua<�ta<�ta<�ta<�ta<�ta<ua<ua<ua<%ua<�ta<Fta<[sa<]ra<qa<�oa<=na<�la<hka<@ja<Hia<�ha<�ha<�ha<Via<Xja<�ka<ma<{na<�  �  �oa<cqa<�ra<�sa<�ta<�ua<�ua<Nva<Jva<Zva<$va<va<va<=va<�va<�va<�wa<$xa<�xa<�ya<dza<{a<+{a<�{a<o{a<!{a<�za<�ya<ya<xa<Twa<iva<va<�ua<�ua<cva<Dwa<�xa<(za<|a<~a<�a<3�a<�a<�a<^�a<�a<��a<��a<^�a<��a<�a<A�a<��a<�a<��a<.�a<Ǝa<��a<��a<��a<m�a<M�a<�a<�a<r�a<�a<ϓa<��a<!�a<��a<��a<��a<��a<~�a<�a<ٌa<%�a<ƍa<�a<�a<��a<��a<��a<3�a<��a<Ԙa<��a<��a<��a<5�a<�a<��a<��a<U�a<4�a<��a<�a<(�a<U�a<��a<�a<��a<�a<;�a<�a< �a<��a<ƚa<�a<��a<|�a<ܕa<��a<"�a<�a<2�a<l�a<�a<F�a<�a<��a<��a<�a<	�a<��a<��a<��a<��a<l�a<��a<��a<��a<X�a< �a<^�a<ߘa<f�a<�a<��a<��a<ӗa<�a<"�a<k�a<d�a<p�a<�a<��a<ؖa<ٕa<��a<*�a<��a<ȏa<R�a<��a<|�a<U�a<��a<&�a<�a<��a<�a<��a<��a<�a<�a<�a<Ϗa<�a<q�a<�a<�a<j�a<��a<��a<��a<��a<�a<e�a<։a<;�a<�a<��a<y�a<,�a<�a<[�a<c�a<��a<=�a<��a< �a<Ga<&}a<9{a<Qya<mwa<va<�ta<�sa<Nsa<.sa<�sa<�sa<�ta<�ua<�va<�wa<jxa<ya<dya<�ya<Oya<Sya<�xa<*xa<jwa<�va<va<�ua<Jua<�ta<�ta<�ta<ua<Dua<Kua<gua<ua<�ta<Ota<Asa<rra< qa<�oa<�ma<�la<4ka<"ja<Oia<�ha<Uha<�ha<Yia<Aja<Oka<�la<5na<�  �  pa<jqa<�ra<�sa<�ta<�ua<�ua<va<va<%va<va<�ua<�ua<va<Qva<�va<Zwa<xa<�xa<�ya<#za<�za<V{a<�{a<u{a<.{a<�za<�ya<ya<:xa<mwa<�va<!va<�ua<"va<�va<}wa<�xa<Qza<%|a<5~a<5�a<G�a<�a<�a<n�a<ވa<׉a<��a<
�a<��a<�a<.�a<��a<݌a<S�a<�a<��a<��a<v�a<h�a<I�a<��a<��a<(�a<]�a<�a<��a<�a<:�a<0�a<-�a<�a<)�a<v�a<�a<	�a<[�a<�a<�a<�a<��a<.�a<a<F�a<��a<ۘa<��a<��a<ޚa<��a<Ϛa<˚a<��a<D�a<�a<ݙa<әa<��a<9�a<��a<��a<l�a<��a<�a<-�a<�a<��a<�a<�a<Øa<��a<�a<Ĕa<V�a<,�a<,�a<��a<]�a<��a<ސa<��a<a<�a<O�a<��a<ėa<�a<��a<f�a<��a<ɚa<��a<)�a<˙a<B�a<Ęa<K�a<�a<��a<��a<��a<՗a< �a<3�a<#�a<8�a<�a<��a<ޖa<�a<��a<2�a<��a< �a<k�a<όa<�a<g�a<ɉa<\�a<W�a<��a<G�a< �a</�a<)�a</�a<�a<��a<�a<a�a<6�a<ԏa<�a<j�a<��a<��a<ɋa<�a</�a<��a<&�a<Ԉa<��a<P�a<�a<��a<4�a<��a<��a<H�a<�a<'�a<`a<^}a<j{a<mya<�wa<
va<�ta<�sa<�sa<Msa<�sa<ta<�ta<�ua<�va<�wa<mxa<ya<kya<�ya<{ya<ya<sxa<�wa<Ewa<�va<�ua<eua<�ta<�ta<�ta<�ta<�ta<ua<ua<ua<%ua<�ta<Fta<[sa<]ra<qa<�oa<=na<�la<hka<@ja<Hia<�ha<�ha<�ha<Via<Xja<�ka<ma<{na<�  �  8pa<�qa<�ra<ta<�ta<Rua<�ua<�ua<va<�ua<�ua<sua<nua<�ua<�ua<Uva<�va<�wa<Xxa<Fya<za<�za<0{a<Q{a<s{a<D{a<�za<&za<Pya<�xa<�wa<"wa<�va<tva<�va<�va<xa<,ya<�za<w|a<z~a<j�a<m�a<c�a<�a<��a<��a<��a<o�a<�a<o�a<v�a<ǋa<�a<`�a<Ȍa<c�a<8�a<��a<�a<��a<$�a<ܒa<��a<�a<%�a<9�a<ѓa<<�a<^�a<b�a<r�a<e�a<��a<�a<��a<z�a<ٍa<�a<_�a<��a<�a<��a<��a<v�a<ɗa<�a<ʙa<B�a<��a<Ěa<��a<��a<�a<ݙa<w�a<o�a<G�a<x�a<��a<
�a<��a<�a<��a<śa< �a<̛a<��a<�a<�a<�a<��a<e�a<�a<��a<��a<��a<=�a<��a<�a<d�a<<�a<+�a<N�a<��a<Җa<�a<�a<ޙa<M�a<y�a<��a<N�a<�a<i�a<јa<=�a<a<r�a<�a<,�a<�a<c�a<��a<��a<�a<�a<�a<g�a<ܖa<��a<ʔa<o�a<ۑa<W�a<��a<S�a<��a<��a<K�a<Éa<�a<�a<Ίa<r�a<t�a<^�a<U�a<9�a<ʏa<<�a<0�a<�a<��a<��a<L�a<"�a<@�a<1�a<q�a<��a<�a<��a<>�a<'�a<܇a<�a<u�a<�a<c�a<k�a<m�a<��a<a�a<�a<�}a<�{a<�ya<%xa<�va<rua<jta<ta<�sa<ta<�ta<7ua<#va<�va<�wa<�xa<$ya<tya<cya<Xya<�xa<exa<�wa<�va</va<bua<�ta<sta<Kta<5ta<<ta<xta<�ta<ua<�ta<�ta<�ta<%ta<�sa<zra<Sqa<�oa<�na<ma<�ka<�ja<�ia<hia<�ha<mia<�ia<�ja<�ka<Dma<�na<�  �  �pa<�qa<sa<ta<�ta<Jua<vua<�ua<Vua<ua<�ta<�ta<�ta<�ta<ua<�ua< va<�va<�wa<�xa<�ya<Iza<�za<R{a<r{a<A{a<�za<~za<�ya<"ya<exa<�wa<Vwa<5wa<nwa<�wa<�xa<�ya<~{a<'}a<#a<�a<؂a<��a<$�a<��a<��a<�a<�a<~�a<��a<ӊa<%�a<B�a<��a<�a<��a<h�a<N�a<k�a<Q�a<a�a<h�a<2�a<ɓa<#�a<1�a<�a<x�a<ǒa<�a<�a<�a<X�a<��a<f�a<\�a<��a<9�a<�a<A�a<��a<�a<t�a<֖a<�a<�a<əa<C�a<i�a<o�a<8�a<ҙa<s�a<+�a<ɘa<��a<��a<��a<��a<`�a<��a<b�a<�a<b�a<��a<��a<��a<��a<>�a<U�a<.�a<�a<��a<]�a<W�a<�a<��a<��a<Ցa<3�a<�a<ʓa<�a<&�a<M�a<W�a<-�a<Йa<M�a<q�a<D�a<�a<d�a<Řa<9�a<��a<	�a<��a<g�a<W�a<o�a<��a<�a<3�a<��a<��a<��a<g�a<ۖa<��a< �a<Ǔa<Y�a<�a<c�a<�a<��a<��a<�a<��a<��a<�a<t�a<"�a<�a<�a<��a<u�a<�a<.�a<,�a<ޏa<J�a<��a<��a<�a<��a<��a<��a<�a<K�a<݇a<��a<��a<9�a< �a<�a<��a<&�a<h�a<e�a<�a<��a<�a<~a<V|a<lza<�xa<Mwa<%va<Mua<�ta<�ta<�ta<;ua<�ua<�va<uwa<9xa<�xa<&ya<sya<dya<ya<�xa<�wa<wa<1va<}ua<�ta<"ta<�sa<{sa<xsa<�sa<�sa<ta<Qta<�ta<�ta<�ta<%ta<nsa<�ra<�qa<Zpa<oa<�ma<nla<kka<�ja<$ja<�ia<,ja<�ja<�ka<�la<�ma<Roa<�  �  Eqa<Mra<isa<$ta<�ta<ua<ua<ua<�ta<xta<ta<�sa<�sa<�sa<ta<kta<*ua<�ua<�va<�wa<�xa<�ya<yza<{a<R{a<r{a<Q{a<�za<eza<�ya</ya<�xa<lxa<@xa<pxa< ya<�ya<{a<n|a<
~a<�a<��a<`�a<�a<m�a<��a<��a<.�a<��a<�a< �a<0�a<�a<C�a<��a<��a<��a<Y�a<S�a<^�a<��a<��a<ؑa<Òa<t�a<��a<$�a<$�a<Ɠa<F�a<��a<��a<��a<F�a<ݏa<d�a<l�a<��a<B�a<7�a<)�a<p�a<��a<�a<D�a<W�a<&�a<��a<�a<�a<��a<��a<'�a<��a<�a<Зa<��a<��a<��a<��a<^�a<�a<��a<=�a<�a<6�a<y�a<_�a<�a<��a<��a<��a<|�a<f�a<L�a<[�a<��a<�a<ϒa<͒a<E�a<�a<��a<��a<��a<ߗa<��a<~�a<�a<(�a<7�a<ڙa<|�a<��a<�a<Q�a<��a<�a<��a<n�a<B�a<x�a<��a< �a<��a<ؖa<:�a<6�a<1�a<��a<+�a<T�a<(�a<�a<s�a<.�a<Ўa<ʍa<ƌa<�a<ċa<��a<�a<e�a<�a<��a<�a<H�a<��a<-�a<0�a<�a<��a<ێa<��a<݌a<܋a<��a<��a<��a<؇a<H�a<φa<��a<r�a<��a<u�a<q�a<;�a<Ѕa<@�a<Y�a<N�a<�a<l�a<�~a<�|a<K{a<�ya<qxa<#wa<]va<�ua<�ua<�ua<"va<�va<Gwa<	xa<�xa<"ya<_ya<Uya<7ya<�xa<xa<;wa<Vva<qua<fta<�sa<sa<�ra<ira<tra<�ra<�ra<asa<�sa<ta<.ta<Ata<�sa<�sa<�ra<�qa<�pa<�oa<{na<^ma<nla<�ka<ka<ka<$ka<�ka<�la<�ma<�na<�oa<�  �  �qa<�ra<�sa<@ta<�ta<�ta<�ta<\ta<ta<zsa<sa<�ra<�ra<�ra<�ra<9sa<�sa<�ta<�ua<wa<4xa<1ya<za<�za<[{a<�{a<�{a<[{a<{a<�za<za<�ya<rya<tya<�ya<-za<{a<-|a<r}a<a<��a<Z�a<�a<H�a<��a<��a<T�a<݈a<#�a<@�a<7�a<#�a<�a<8�a<\�a<ĉa<b�a<-�a<@�a<]�a<��a<ݏa<$�a<5�a<#�a<Ǔa<;�a<I�a<�a<Γa<L�a<��a<��a<K�a<�a<��a<��a<�a<z�a<>�a<8�a<d�a<��a<Ŗa<��a<��a<N�a<��a<ՙa<��a<]�a<�a<C�a<��a<�a<��a<R�a<L�a<`�a<Ȗa<Z�a<��a<��a<��a<=�a<ƚa<*�a<C�a<,�a<��a<�a<T�a<Q�a<C�a<K�a<_�a<��a<5�a<�a<�a<n�a<��a<a<��a<��a<x�a<'�a<��a<
�a<�a<�a<m�a<̘a<�a< �a<E�a<��a<ߔa<Y�a<�a<�a<K�a<��a<�a<��a<3�a<��a<ۖa<�a<Ėa<M�a<��a<��a<��a<V�a<�a<�a<Ўa<��a<U�a<�a<�a<�a<h�a<	�a<��a<N�a<֏a<�a<L�a<H�a<؏a<<�a<Z�a<K�a<�a<ϊa<��a<}�a<m�a<��a<
�a<��a<��a<r�a<��a<��a<��a<��a<�a<�a<p�a<r�a<@�a<�a<za<�}a<K|a<�za<yya<hxa<�wa<wa<�va<�va<2wa<�wa<3xa<�xa<"ya<]ya<�ya<aya<�xa<Zxa<|wa<�va<rua<ita<isa<�ra<�qa<xqa<4qa<Hqa<�qa<�qa<]ra<�ra<jsa<�sa<�sa<�sa<�sa<sa<Tra<�qa<npa<Xoa<\na<sma<�la<_la<)la<gla<�la<�ma<�na<�oa<�pa<�  �  _ra<Wsa<�sa<`ta<�ta<nta<9ta<�sa</sa<ra<ra<�qa<9qa<Eqa<jqa< ra<�ra<�sa<�ta<va<iwa<�xa<�ya<�za<Q{a<�{a<�{a<�{a<�{a<g{a<{a<�za<�za<�za<{a<�{a<V|a<L}a<�~a<�a<��a<�a<j�a<ǅa<��a<��a<,�a<��a<��a<��a<X�a<�a<�a<�a<�a<�a<�a<�a<�a<A�a<��a<��a<i�a<��a<ʒa<��a<B�a<p�a<��a<S�a<��a<p�a<�a<�a<�a<�a<��a<I�a<��a<m�a<e�a<L�a<f�a<\�a<L�a< �a<p�a<��a<��a<Y�a<��a<(�a<T�a<��a<�a<P�a<�a<�a<#�a<w�a<�a<�a<��a<��a<y�a<T�a<ؚa<+�a<D�a<��a<��a<Йa<$�a<2�a<c�a<��a<�a<��a<F�a<m�a<��a<)�a<��a<��a<e�a<��a<��a<��a<*�a<�a<��a<�a<�a<<�a<$�a<>�a<K�a<��a<�a<Ēa<֒a<�a<t�a<�a<��a<h�a<�a<|�a<��a<��a<m�a<�a</�a<*�a<-�a<�a<�a<�a<5�a<��a<H�a<0�a<8�a<��a<�a<}�a<
�a<R�a<��a<z�a<R�a<��a<�a<؍a<��a<5�a<��a<~�a<)�a<$�a<[�a<��a<Y�a<)�a<V�a<v�a<��a<�a<$�a<&�a<ӄa<w�a<��a<��a<y�a<*�a<�~a<@}a<�{a<�za<�ya<�xa<rxa<%xa<xa<_xa<�xa<	ya<]ya<�ya<�ya<�ya<`ya<�xa<�wa<�va<�ua<�ta<esa<Fra<<qa<�pa<pa<�oa<�oa<Jpa<�pa<[qa<ra<�ra<Lsa<�sa<�sa<�sa<Psa<�ra<�qa<Aqa<Fpa<toa<�na<�ma<�ma<�ma<�ma<na<�na<�oa<�pa<�qa<�  �  sa<�sa<6ta<ota<jta<ta<�sa<sa<Qra<�qa<�pa<Opa<pa<�oa<pa<�pa<zqa<�ra<�sa<#ua<�va<xa<5ya<Kza<={a<�{a<;|a<`|a<c|a<E|a<|a<�{a<�{a<�{a<D|a<�|a<�}a<�~a<�a<�a<m�a<ڃa<�a<*�a<�a<��a<	�a<�a<�a<�a<��a<,�a<ֆa<��a<Іa<�a<��a<��a<��a<�a<��a<&�a<��a<"�a<V�a<k�a<<�a<��a<�a<�a<��a<T�a<��a<��a<d�a<5�a<M�a<��a<�a<��a<x�a<X�a<D�a<�a<͘a<R�a<��a<��a<U�a<֘a<@�a<g�a<o�a<��a<��a<-�a<ȓa<��a<˓a<>�a<�a<Ǖa<Ζa<ٗa<�a<əa<v�a<�a<P�a<E�a<��a<��a<�a<%�a<m�a<��a<:�a<ʖa<��a<��a<��a<`�a<�a<��a<5�a<��a<�a<K�a<:�a<�a<A�a<~�a<��a<^�a<:�a<�a<�a<W�a<a<l�a<�a<Ǒa<@�a<��a<��a<��a<h�a<�a<_�a<��a<��a<>�a<��a<�a<�a<�a<�a<I�a<��a<�a<��a<u�a<��a<a<�a<h�a<ϐa<�a< �a<Ɛa<P�a<��a<x�a<I�a<�a<_�a<؈a<O�a<��a<�a<��a<[�a<�a<�a<#�a<��a<�a<W�a<��a<��a<��a<q�a<كa<�a<	�a<�a<�a<I~a<}a<�{a<�za<>za<�ya<mya<iya<rya<�ya<�ya<za<0za<za<�ya<Sya<xxa<twa<_va<ua<�sa<Xra<qa<pa<Roa<�na<�na<�na<oa<�oa<spa<@qa<ra<�ra<?sa<�sa<�sa<�sa<<sa<�ra<ra<8qa<}pa<�oa<Toa<�na<�na<�na<loa<�oa<�pa<zqa<`ra<�  �  �sa< ta<�ta<wta<Mta<�sa</sa<�ra<xqa<�pa<�oa<Hoa<�na<�na<�na<coa<^pa<{qa<�ra<Gta<�ua<vwa<�xa<*za<%{a<�{a<�|a<�|a<}a<�|a<}a<�|a<�|a<'}a<{}a<'~a<�~a<�a<ɀa<"�a<P�a<��a<��a<z�a<A�a<��a<�a<ׇa<��a<#�a<��a<5�a<Ʌa<��a<��a<�a<��a<^�a<��a<�a<��a<;�a<��a<��a<�a<E�a<'�a<�a<@�a<v�a<m�a<3�a<�a<��a<{�a<a�a<��a<Ôa<.�a<Õa<|�a<b�a<�a<̘a<G�a<��a<��a<��a<7�a<l�a<��a<��a<��a<��a<��a<�a<}�a<n�a<��a<�a<ݓa<��a<�a<��a<K�a<J�a<F�a<�a<L�a<��a<]�a<0�a<��a<�a<w�a<Ęa<i�a<��a<�a<ڗa<#�a<d�a<�a<~�a<ݙa<a�a<z�a<��a<B�a<șa<�a<��a<�a<��a<Y�a<�a<�a<,�a<�a<J�a<8�a<��a<:�a<��a<ߒa<ȓa<Քa<}�a<>�a<��a<��a<��a<�a<��a<��a<�a<�a<L�a<��a<#�a<�a<��a<��a<��a<�a<K�a<w�a<��a<Q�a<�a<A�a<f�a<6�a<ˌa</�a<r�a<�a<C�a<��a<��a<Âa<*�a<Ӂa<��a<�a<��a<��a<��a<�a<b�a<��a<[�a<�a<d�a<��a<��a<o�a<Xa<~a<}a< |a<�{a<�za<�za<qza<uza<�za<�za<�za<�za<nza<�ya<<ya<Zxa<wa<�ua<<ta<�ra<Tqa<
pa<oa<na<�ma<`ma<�ma<na<�na<�oa<`pa<xqa<Bra<sa<�sa<�sa<�sa<�sa<\sa<�ra<(ra<�qa<�pa<�pa<&pa<.pa<0pa<�pa<�pa<�qa<sra<sa<�  �  8ta<�ta<�ta<�ta<,ta<�sa<�ra<�qa<�pa<�oa<�na<=na<�ma<�ma<�ma<nna<Hoa<{pa<�qa<�sa<9ua<�va<~xa<�ya<{a<|a<�|a<>}a<�}a<�}a<�}a<�}a<�}a<1~a<�~a< a<�a<a<߁a<܂a<��a< �a<�a<҆a<l�a<��a<��a<��a<#�a<��a<�a<_�a<��a<��a<��a<�a<v�a<_�a<��a<�a<Ŋa<��a<a�a<"�a<��a<�a<;�a<�a<��a<�a< �a<ݕa<��a<��a<u�a<q�a<��a<Εa<?�a<Ŗa<��a<�a<��a<R�a<��a<�a<�a<��a<�a<(�a<"�a<�a<�a<��a<��a<��a<��a<N�a<��a< �a<ʒa<Γa<�a<p�a<��a<�a<��a<��a<m�a<Ǜa<ěa<��a<@�a<��a<I�a<љa<^�a<�a<�a<�a<�a<k�a<әa<'�a<��a<Ӛa<�a<њa<g�a<��a<Øa<��a<_�a<��a<��a<$�a<�a<�a<��a<'�a<B�a<��a<;�a<�a<4�a<7�a<D�a<9�a<�a<s�a<Жa<ϖa<��a<�a<m�a<��a<�a<O�a<��a<3�a<�a<��a<��a<֑a<ؑa<��a<�a<��a<��a<-�a<]�a<)�a<�a<Z�a<��a<�a<�a<Y�a<׃a<��a<��a<�a<Ԁa<ڀa</�a<��a<f�a<��a<��a<�a<I�a<o�a<8�a<��a<�a<.�a<�a<�a<a<	~a</}a<|a<�{a<�{a<s{a<z{a<R{a<T{a<S{a<{a<�za<za<2ya<xa<�va<Bua<�sa<ra<opa<oa<�ma<ma<{la<`la<�la<�la<�ma<�na<�oa<�pa<�qa<�ra<]sa<�sa< ta<ta<�sa<\sa<�ra<Yra<�qa<xqa<8qa<(qa<Aqa<�qa<ra<�ra<sa<�sa<�  �  �ta<�ta<�ta<�ta<7ta<wsa<�ra<qqa<`pa<:oa<Ona<�ma<�la<�la<�la<�ma<una<�oa<7qa<�ra<�ta<rva<=xa<�ya<!{a<|a<�|a<�}a<�}a<a~a<S~a<�~a<�~a<�~a<Xa<�a<��a<p�a<��a<~�a<��a<��a<h�a<�a<k�a<��a<��a<I�a<��a<�a<l�a<��a<G�a<҃a<كa<	�a<��a<��a<φa<z�a<�a<�a<ٍa<��a<{�a<��a<A�a<�a<ٕa<;�a<y�a<��a<V�a<Y�a<#�a<D�a<N�a<��a<�a<m�a< �a<��a<q�a<��a<�a<�a<�a<��a<Иa<�a<��a<w�a<B�a<�a<�a<)�a<Аa<i�a<Đa<;�a<�a<6�a<j�a<��a<4�a<��a<ęa<Ěa<o�a<ƛa<�a<��a<ۛa<j�a<�a<��a<�a<�a<��a<��a<ԙa<�a<l�a<̚a<3�a<.�a<<�a<Ԛa<g�a<��a<��a<_�a<��a<m�a<ߒa<��a<Y�a<N�a<Ďa<>�a<��a<��a<��a<e�a<��a<��a<Гa<��a<ѕa<��a<Жa<�a<�a<{�a<'�a<Q�a<��a<��a<w�a< �a<��a<��a<\�a<��a<z�a<��a<��a<Q�a<�a<+�a<a�a<$�a<��a<��a<�a<I�a<X�a<��a<�a<�a<�a<>�a<"�a<�a<��a<��a<Áa<r�a<3�a<؃a<=�a<u�a<:�a<��a<`�a<��a<܁a<��a<�a<�~a<~a<>}a<�|a<l|a<|a<|a<�{a<|a<�{a<x{a<�za<za<Cya<�wa<�va<�ta<sa<sqa<�oa<ona<ma<Zla<�ka<�ka<�ka<Kla< ma<na<Goa<apa<�qa<�ra<bsa<�sa< ta<Yta<$ta<�sa<}sa<�ra<�ra<)ra<ra<�qa<ra<Hra<�ra<1sa<�sa<]ta<�  �  �ta<ua<ua<�ta<ta<Rsa<Hra<Fqa<pa<�na<�ma<ma<ula<bla<�la< ma<�ma<Poa<�pa<�ra<ota<Iva<�wa<�ya<�za<>|a<$}a<�}a<~a<x~a<�~a<�~a<+a<sa<�a<f�a< �a<��a<�a<�a<�a<��a<��a<A�a<��a<��a<��a< �a<��a<݅a<�a<b�a<��a<Y�a<;�a<��a<!�a<�a<W�a<�a<ǉa<��a<��a<��a<H�a<�a< �a<M�a<��a<p�a<��a<Ȗa<ʖa<��a<��a<��a<ۖa<�a<��a<�a<��a<�a<��a<��a<A�a<F�a<�a<l�a<��a<��a<��a<?�a<��a<��a<��a<��a<7�a<�a<@�a<��a<��a<��a<'�a<��a<�a<X�a<��a<��a<v�a<�a<C�a<.�a<�a<a<Z�a<��a<��a<Z�a<0�a<=�a<^�a<��a<ߚa<+�a<E�a<c�a<h�a<�a<{�a<��a<y�a<�a<��a<�a<��a<�a<ُa<ǎa<9�a<ڍa<��a<D�a<�a<	�a<C�a<l�a<��a<��a<��a<_�a<��a<%�a<�a<��a<>�a<��a<#�a<��a<��a<��a<+�a<��a<�a<�a<�a<�a<��a<��a<�a<o�a<N�a<�a<��a<ˋa<�a<��a<�a<2�a<��a<L�a<i�a<�a<�a<�a<�a<��a<{�a<B�a<�a<��a<*�a<T�a<u�a<�a<��a<��a<�a<�a<*�a<Ia<w~a<�}a<D}a<�|a<�|a<�|a<a|a<1|a<�{a<�{a<{a<Lza<ya<�wa<Ava<�ta<�ra</qa<loa<�ma<�la<�ka<1ka<ka</ka<�ka<�la<�ma<�na<1pa<Pqa<gra<Jsa<�sa<gta<�ta<Yta<ta<�sa<isa<sa<�ra<�ra<kra<�ra<�ra<6sa<�sa<ta<pta<�  �  va<va<va<�ua<�ua<(ua<>ta<�sa<�ra<�qa<qa<�pa<7pa<pa<Npa<�pa<�qa<�ra<�sa<`ua<�va<dxa<�ya<X{a<H|a<A}a<~a<�~a<Ia<�a<�a<5�a<��a<�a<P�a<�a<��a<h�a<9�a<�a<��a<��a<��a<��a<m�a<��a<ֈa<��a</�a<͇a<B�a<�a<��a<��a<��a<ӆa<i�a<Z�a<k�a<��a<J�a<��a<j�a< �a<}�a<�a<a<��a<b�a<�a<0�a<v�a<��a<��a<��a<��a<��a<�a<y�a<�a<]�a<ʙa<K�a<��a<��a<ǚa<��a<4�a<�a<��a<�a<�a<&�a<F�a<m�a<ܓa<��a<F�a<r�a<�a<��a<o�a<��a<��a<ǘa<̙a<�a<��a<�a<��a<��a<�a<��a<|�a<,�a<��a<��a<l�a<b�a<P�a<x�a<��a<��a<�a<�a<!�a<�a<��a<�a<��a<Ιa<��a<q�a<�a<�a<Гa<Ւa<�a<|�a<.�a<B�a<��a<��a<��a<��a<O�a<Q�a<�a<��a<@�a<��a<��a<��a<h�a<�a<{�a<��a<��a<�a<��a<J�a<�a<��a<֓a<��a<��a<c�a<#�a<��a<�a<��a<&�a<a<?�a<��a<�a<��a<
�a<Åa<��a<��a<%�a<�a<тa<��a<c�a<��a<C�a<��a<%�a<��a<N�a<@�a<�a<w�a<ǃa<�a<D�a<s�a<��a<�a<Ia<�~a<\~a<~a<�}a<�}a<l}a<}a<�|a<|a<O{a<^za<�ya<xa<�va<6ua<�sa<�ra<Bqa<Kpa<�oa<�na<�na<�na<Ooa<�oa<�pa<oqa<{ra<Ksa<:ta<�ta<ua<yua<�ua<�ua<`ua<ua<�ta<�ta<\ta<ta<(ta</ta<vta<�ta<ua<gua<�ua<�  �  �ua<-va< va<�ua<�ua<�ta<Gta<�sa<�ra<�qa<5qa<�pa<Npa<^pa<�pa<qa<�qa<�ra<ta<�ua<�va<xa<�ya<{a<O|a<[}a<$~a<�~a<5a<�a<�a<�a<P�a<a<%�a<��a<y�a<)�a<�a<�a<܅a<��a<}�a<�a<��a<��a<��a<p�a<B�a<�a<�a<�a<ǆa<��a<��a<�a<��a<��a<��a<�a<W�a<��a<��a<�a<d�a<��a<�a<ѕa<q�a<�a<(�a<Q�a<Z�a<f�a<i�a<��a<��a<�a<_�a<��a<;�a<��a<+�a<��a<Κa<Кa<��a<B�a<��a<�a<4�a<>�a<N�a<[�a<��a<�a<��a<��a<��a<
�a<Ɣa<��a<��a<a<�a<ڙa<��a<��a<6�a<��a<՜a<Ҝa<��a<b�a<�a<Ûa<��a<W�a<&�a<2�a<I�a<e�a<��a<͛a<��a<�a<�a<��a<7�a<|�a<��a<��a<��a<Q�a<�a<�a<�a<%�a<��a<p�a<r�a<��a<+�a<͒a<��a<��a<l�a<�a<��a<G�a<��a<��a<��a<T�a<�a<c�a<�a<G�a<�a<j�a<�a<��a<��a<��a<��a<��a<W�a<�a<��a<�a<�a<�a<��a<R�a<܋a<B�a<��a<6�a<�a<τa<�a<h�a<�a<��a<*�a<p�a<�a<i�a<Єa<�a<M�a<m�a<V�a<��a<z�a<��a<��a<�a<H�a<q�a<�a<a<�~a<B~a<�}a<�}a<v}a<K}a<�|a<�|a<|a<f{a<lza<Aya<xa<�va<dua<�sa<�ra<tqa<^pa<�oa<>oa<oa<oa<~oa<pa<�pa<�qa<�ra<Zsa<ta<�ta<8ua<�ua<�ua<�ua<Mua< ua<�ta<`ta<&ta<	ta<�sa<ta<Gta<�ta<�ta<Hua<�ua<�  �  �ua<�ua<�ua<�ua<�ua<ua<�ta<�sa<�ra<0ra<�qa<qa<�pa<�pa<�pa<dqa<ra<Hsa<Yta<�ua<$wa<�xa<za<5{a<o|a<A}a<�}a<�~a<�~a<Ya<�a<�a<�a<m�a<݀a<c�a<'�a<ɂa<΃a<��a<��a<��a<<�a<߇a<K�a<��a<Èa<��a<��a<�a<��a<G�a< �a<�a<�a<W�a<�a<׈a<�a<I�a<��a<5�a<��a<I�a<��a<Փa<�a<��a<?�a<��a<��a<	�a<�a<.�a<�a<I�a<`�a<��a<�a<]�a<�a<i�a<�a<G�a<��a<��a<��a<a�a<řa<D�a<[�a<f�a<��a<��a<�a<M�a<��a<Ɠa<�a<`�a<*�a<�a<ۖa<��a<��a<%�a<�a<��a<1�a<b�a<��a<��a<t�a<�a<ٛa<��a<#�a<�a<ٚa<�a<�a<"�a<h�a<��a<ɛa<ța<ța<r�a<+�a<��a<��a<�a<��a<��a<X�a<C�a<j�a<��a<�a<��a<��a<��a<��a<�a<�a<��a<��a<i�a<ږa<h�a<��a<y�a<r�a<�a<��a<�a<��a<��a<��a<!�a<Ɠa<��a<X�a<k�a<S�a<<�a<&�a<ےa<q�a<ˑa<�a<�a<�a<��a<�a<��a<�a<��a<H�a<!�a<?�a<��a<g�a<W�a<��a<��a<-�a<��a<�a<Z�a<m�a<�a<%�a<Ąa<;�a<��a<��a<ہa<�a<�a<~a<�~a<L~a<�}a<�}a<|}a<2}a<	}a<�|a<o|a<�{a<E{a<�za<gya<bxa<�va<�ua<?ta<�ra<�qa<�pa<pa<voa<[oa<foa<�oa<^pa<qa<�qa<�ra<�sa<>ta<�ta<3ua<Fua<dua<Aua<ua<�ta<sta< ta<�sa<�sa<�sa<�sa<�sa<Eta<�ta<ua<zua<�  �  ~ua<�ua<�ua<�ua<�ua<,ua<�ta<�sa<Rsa<�ra<ra<�qa<Lqa<Nqa<�qa<	ra<�ra<�sa<�ta<Lva<�wa<�xa<za<W{a<S|a<2}a<�}a<X~a<�~a<�~a<a<Ea<�a<�a<*�a<ˀa<V�a<S�a<0�a</�a<�a<�a< �a<·a<S�a<��a<ވa<��a<��a<d�a<#�a<�a<��a<��a<��a<�a<��a<y�a<q�a<��a<9�a<��a<�a<w�a<��a<��a<єa<��a<6�a<n�a<��a<��a<��a<��a<��a<|�a<Ėa<��a<O�a<�a<b�a<�a<y�a<��a<I�a<��a<��a<C�a<�a<7�a<��a<Ηa<�a<3�a<u�a<�a<��a<��a<��a<�a<��a<h�a<x�a<W�a<G�a</�a<��a<��a<�a<|�a<y�a<V�a<�a<��a<N�a<�a<��a<;�a<J�a<#�a<X�a<��a<֚a<�a<Z�a<��a<��a<��a<�a<��a<ҙa<�a<�a<�a<�a<Ŕa<ޓa<$�a<��a<l�a<f�a<��a<�a<��a<p�a<�a<Ǖa<a�a<��a<M�a<{�a<��a<4�a<Ԗa<E�a<��a<�a<��a<�a<n�a<.�a<Ғa<�a<͒a<Ւa<ƒa<��a<��a<_�a<ӑa<�a<.�a<�a<��a<O�a<�a<��a<�a<Ɇa<Åa<�a<c�a<
�a<؃a<�a<S�a<��a<�a<5�a<X�a<��a<]�a<�a<��a<��a<+�a<@�a<^�a<m�a<�a<�~a<-~a<�}a<2}a<}a<�|a<�|a<�|a<{|a<*|a<�{a<7{a<mza<�ya<Uxa<3wa<�ua<�ta<tsa<Jra<Sqa<�pa<<pa<pa<pa<Zpa<�pa<�qa<Dra<�ra<�sa<Ota<�ta<ua<_ua<Cua<ua<�ta<Cta<�sa<�sa<=sa<�ra<sa<sa<Vsa<�sa<#ta<�ta<ua<�  �  (ua<Tua<�ua<�ua<�ua<wua<�ta<�ta<�sa<6sa<�ra<Nra<
ra<�qa<Vra<�ra<zsa<eta<�ua<�va<�wa<uya<iza<�{a<k|a<}a<�}a<�}a<^~a<f~a<�~a<�~a<�~a<a<la<�a<��a<��a<Z�a<��a<��a<��a<��a<]�a<0�a<��a<�a<�a<�a<�a<��a<x�a<A�a<L�a<c�a<͈a<i�a<$�a<;�a<a�a<ȍa<��a<��a<�a<��a<#�a<Ԕa<��a<ҕa<�a<8�a<�a< �a<��a<��a<ŕa<�a<B�a<��a<3�a<��a<�a<��a<��a<�a<S�a<l�a<P�a<&�a<��a<!�a<>�a<m�a<іa<!�a<��a<E�a<P�a<]�a<a<b�a<�a<��a<��a<�a<��a<H�a<ӛa<�a<F�a<	�a<��a<��a<8�a<��a<�a<�a<�a<��a<e�a<��a<șa<+�a<��a<ޚa<=�a<*�a<M�a<�a<��a<�a<D�a<��a<L�a<_�a<l�a<��a<�a<Y�a<6�a<�a<P�a<��a<C�a<Ԕa<��a<b�a<��a<?�a<d�a<e�a<G�a<ϖa<|�a<a<9�a<L�a<��a<4�a<��a<}�a<�a<B�a<��a<O�a<U�a<[�a<C�a<�a<��a<�a<Q�a<3�a<�a<،a<G�a<�a<��a<��a<y�a<��a<%�a<��a<��a<��a<�a<��a<f�a<��a<��a<��a<`�a<
�a<W�a<��a<ςa<Ɂa<�a<�a<�~a<�}a<x}a<�|a<�|a<]|a<|a<H|a<|a<&|a<�{a<�{a<#{a<zza<�ya<�xa<�wa<cva<ua<ta<�ra<ra<Rqa< qa<�pa<�pa<qa<�qa<"ra<�ra<�sa<ta<�ta<�ta<ua<)ua<�ta<�ta<8ta<�sa<Nsa<�ra<�ra<2ra<bra<Era<�ra<�ra<xsa<"ta<�ta<�  �  �ta<)ua<�ua<�ua<�ua<�ua<Qua<�ta<kta<�sa<ysa< sa<�ra<�ra<9sa<�sa<hta<>ua<Iva<xwa<�xa<�ya<�za<�{a<||a<}a<x}a<�}a<�}a<�}a<�}a<�}a<�}a<0~a<s~a<a<�a<��a<��a<�a<��a<,�a<D�a<1�a<�a<��a<��a<X�a<X�a<J�a<L�a< �a<�a<)�a<S�a<��a<R�a<�a<$�a<9�a<s�a<̏a<��a<)�a<Y�a<�a<�a<l�a<��a<��a<��a<]�a<]�a<�a<�a<�a<�a<A�a<ĕa<X�a<��a<��a<J�a<�a<��a<�a<^�a<g�a<&�a<�a<Z�a<Řa<:�a<��a<��a<��a<D�a<2�a<X�a<��a<3�a<�a<��a<v�a<*�a<�a<~�a<қa<�a<�a<��a<��a<�a<d�a<��a<r�a<�a<��a<��a<w�a<��a<�a<u�a<ҙa<H�a<Ěa<��a<�a<�a<��a<B�a<��a<Řa<��a<�a<6�a<m�a<˔a<Z�a<�a<�a<?�a<��a<�a<��a<�a<��a<�a<H�a<u�a<]�a<�a<��a<��a<�a<k�a<��a<��a<Q�a<��a<r�a<5�a<O�a<W�a<��a<��a<ґa<�a<a<��a<�a<G�a<��a<h�a<5�a<�a<��a<��a<k�a<h�a<��a<�a<��a<��a<w�a<��a<Åa<΅a<�a<�a<��a<v�a<�a<%�a<J�a<F�a<�a< �a<�~a<~a<}a<p|a<�{a<�{a<�{a<q{a<~{a<j{a<�{a<�{a<b{a<{a<�za<�ya<ya<�wa<�va<�ua<�ta<�sa<sa<Qra<�qa<�qa<�qa<�qa<Sra<�ra<csa<�sa<jta<�ta<�ta<ua<�ta<�ta<Cta<�sa<sa<�ra<ra<�qa<Hqa<Lqa<Wqa<�qa<8ra<�ra<Nsa<�sa<�  �  ta<�ta<Dua<�ua<�ua<�ua<�ua<Iua<"ua<�ta<Gta<�sa<�sa<�sa<4ta<�ta<Dua<"va<wa<'xa<=ya<za<6{a<�{a<�|a<�|a<:}a<P}a<4}a<M}a<}a<
}a<�|a<0}a<�}a<~a<�~a<�a<ހa<�a<_�a<��a<��a<��a<��a<��a<�a<��a<��a<ԉa<�a<݉a<��a<��a<I�a<��a<L�a<�a<��a<�a<7�a<��a<��a<��a<��a<8�a<�a<�a<l�a<1�a<�a<�a<��a<D�a<�a<�a<�a<Z�a<Ȕa<X�a<(�a<�a<ٗa<y�a<6�a<ۙa<�a<n�a<R�a<R�a<��a<o�a<�a<K�a<ٗa<q�a<A�a<4�a<Z�a<��a<�a<��a<]�a</�a<��a<R�a<��a<�a<�a<ɛa<��a<�a<��a<ϙa<�a<��a< �a<��a<��a<��a<��a<"�a<��a<.�a<љa<�a<��a<՚a<�a<Ța<v�a<�a<:�a<��a<͗a<�a<K�a<��a<[�a<�a<�a<�a<m�a<Ǖa<M�a<ɖa<��a<��a<t�a<}�a<(�a<Жa<-�a<R�a<��a<��a<Ғa<��a<P�a<ِa<��a<W�a<N�a<{�a<��a<�a<A�a<L�a<��a<>�a<�a<a�a<Ϗa<ˎa<��a<Ča<w�a<f�a<@�a<^�a<��a<�a<��a<^�a<Y�a<P�a<z�a<e�a<L�a<O�a<υa<o�a<��a<�a<��a<��a<��a<Ca<&~a<}a<7|a<�{a<�za<�za<�za<�za<�za<�za<�za<{a<${a<�za<�za<�ya<oya<[xa<�wa<�va<�ua<�ta<�sa<Msa<�ra<�ra<�ra<�ra<&sa<�sa<ta<Wta<�ta<
ua<ua<ua<�ta<jta<�sa<+sa<mra<�qa<%qa<�pa<spa<Ypa<�pa<�pa<Eqa<�qa<�ra<�sa<�  �  �sa<nta<ua<�ua<�ua<va<va<�ua<�ua<Pua<ua<�ta<�ta<�ta<)ua<�ua<Iva<
wa<�wa<�xa<�ya<�za<r{a<|a<�|a<�|a<�|a<�|a<�|a<�|a<]|a<3|a<%|a<?|a<�|a<}a<�}a<�~a<�a<E�a<��a<��a<I�a<��a<��a<��a<[�a<ىa<8�a<w�a<p�a<��a<Ȋa<��a<?�a<��a<:�a< �a<��a<�a<�a<��a<(�a<�a<ݓa<��a<�a<��a<�a<˔a<{�a<2�a<��a<a�a<1�a<�a<�a<b�a<ԓa<��a<L�a<*�a<$�a<��a<Әa<��a<�a<{�a<��a<��a<X�a<��a<n�a<)�a<��a<w�a<�a<(�a<5�a<��a<�a<��a<�a<��a<L�a<��a<��a<�a<��a<��a<5�a<�a<ϙa<�a<R�a<��a<#�a<a<��a<��a<ܖa<B�a<їa<{�a<�a<��a<C�a<��a<ޚa<�a<��a<_�a<�a<&�a<y�a<ܗa<C�a<��a<3�a<
�a<�a< �a<U�a<��a<ۖa<M�a<��a<��a<×a<��a<�a<��a<Ǖa<הa<�a<�a<��a<�a<_�a<ڏa<~�a<X�a<w�a<��a<�a<W�a<��a<�a<4�a<�a<�a<��a<
�a<G�a<b�a<4�a<N�a<6�a<@�a<T�a<��a<��a<��a<^�a<-�a<+�a<�a<�a<ֆa<��a<�a<r�a<~�a<��a<V�a<�a<�a<~~a<D}a<:|a<8{a<�za<za<�ya<�ya<�ya<�ya<Eza<sza<�za<�za<�za<�za<Cza<�ya<�xa<!xa<wa<hva<�ua<�ta<*ta<�sa<�sa<�sa<�sa<�sa<Eta<�ta< ua</ua<Jua<>ua<�ta<�ta<�sa<6sa<wra<�qa<�pa<Bpa<�oa<uoa<]oa<�oa<�oa<fpa<qa<�qa<�ra<�  �  `sa<ta<�ta<�ua<�ua<Gva<>va<mva<1va<$va<�ua<�ua<�ua<�ua<>va<ova<7wa<�wa<�xa<�ya<Mza<{a<�{a<J|a<�|a<�|a<�|a<�|a<k|a<�{a<�{a<d{a<S{a<V{a<�{a<9|a<�|a<�}a<#a<��a<�a<w�a<�a<;�a<��a<��a<l�a<�a<��a<�a<&�a<|�a<b�a<ߋa<�a<��a<C�a<ۍa<�a<��a<Րa<��a<��a<k�a<�a<��a<Дa<�a<��a<��a<�a<c�a<�a<��a<@�a<�a<3�a<q�a<�a<��a<w�a<��a<a�a<��a<��a<I�a<�a<h�a<ƚa<��a<��a<��a<>�a<�a<]�a<h�a<�a<5�a<+�a<��a<Ιa<5�a<�a<B�a<ʛa<�a<1�a<�a<�a<��a<Ӛa<M�a<6�a<X�a<��a<ʖa<5�a<��a<��a<��a<�a<m�a<
�a<��a<r�a<u�a<�a<��a<ؚa<�a<�a<��a<^�a<��a<M�a<��a<��a<��a<$�a<�a<͖a<�a<��a<g�a<��a<ڗa<�a<�a<�a<��a<�a<Q�a<t�a<��a<6�a<B�a<-�a<J�a<v�a<�a<��a<[�a<��a<��a<6�a<��a<�a<��a<̐a<�a<�a<��a<E�a<��a<�a<�a<�a<ыa<!�a</�a<��a<��a<l�a<J�a<ɇa<�a<��a<��a<)�a<��a<3�a<\�a<��a<9�a<�a<��a<a<�}a<j|a<I{a<Aza<�ya<ya<�xa<�xa<�xa<Iya<�ya<za<fza<�za<�za<�za<gza<�ya<\ya<�xa<�wa<.wa<1va<�ua<ua<�ta<�ta<�ta<�ta<�ta<ua</ua<~ua<hua<�ua<Cua<�ta<rta<�sa<sa<�qa<�pa<*pa<hoa<�na<rna<yna<}na<�na<�oa<Xpa<:qa<$ra<�  �  �ra<�sa<�ta<uua<va<�va<�va<�va<�va<�va<�va<yva<rva<�va<�va<)wa<�wa<�xa<Aya<�ya<�za<v{a<	|a<z|a<�|a<�|a<s|a</|a<�{a<s{a<({a<�za<�za<�za<�za<w{a<@|a<0}a<{~a<�a<��a<�a<��a<�a<f�a<|�a<�a<b�a<֊a<X�a<��a<�a<2�a<��a<ʌa<^�a<��a<��a<��a<\�a<J�a<*�a<�a<��a<l�a<��a<̔a<Ӕa<j�a<�a<��a<�a<z�a<ݑa<y�a<d�a<q�a<��a<0�a<�a<ɓa<��a<��a<�a<�a<�a<�a<n�a<�a<!�a<�a<�a<��a<z�a<2�a<�a<��a<�a<�a<.�a<��a<�a<U�a<ěa<#�a<T�a<u�a<1�a<ћa<F�a<}�a<��a<Ęa<�a<�a<�a<w�a<�a<�a<�a<1�a<��a<f�a<Q�a<�a<טa<��a<<�a<��a<��a<-�a<��a<��a<=�a<��a<@�a<ǘa<L�a<�a<̗a<��a<��a<͗a<��a<�a<I�a<e�a<V�a< �a<��a<��a<	�a<�a<�a<ϒa<��a<~�a<��a<��a<,�a<ڍa<��a<��a<�a<��a<,�a<��a<&�a<}�a<�a<�a<ΐa<��a<�a<B�a<d�a<��a<��a<ًa<ߊa<F�a<��a< �a<��a<��a<d�a<"�a<�a<}�a<�a<I�a<X�a<Y�a<��a<��a<)�a<�~a<>}a<�{a<�za<�ya<�xa<Txa<xa<xa<?xa<�xa<ya<�ya<�ya<Lza<�za<�za<�za<>za<�ya<ya<^xa<�wa<wa<rva<�ua<�ua<Aua<2ua<Nua<aua<�ua<�ua<�ua<�ua<�ua<Xua<�ta<*ta<Hsa<era<mqa<�pa<�oa<�na<na<�ma<�ma<�ma<1na<�na<�oa<�pa<�qa<�  �  rra<�sa<�ta<}ua<va<qva<�va<�va<wa<wa<wa< wa<wa<;wa<{wa<�wa<`xa<ya<�ya<nza<({a<�{a<'|a<f|a<�|a<�|a<g|a<!|a<{a<{a<�za<>za<za<�ya<<za<�za<�{a<�|a<~a<Wa<
�a<��a<S�a<��a<>�a<��a<��a<]�a<�a<��a<�a<g�a<،a<�a<��a<�a<��a<Z�a<�a<�a<ȑa<��a<g�a<�a<r�a<��a<�a<��a<p�a<�a<)�a<��a<Ցa<r�a<��a<��a<��a< �a<��a<g�a<S�a<S�a<��a<��a< �a<��a<ՙa<��a<�a<8�a<S�a<V�a<&�a<��a<Кa<��a<��a<z�a<��a<Ԛa<�a<��a<͛a<5�a<`�a<��a<`�a<@�a<�a<(�a<��a<i�a<c�a<e�a<a�a<��a<ٔa<s�a< �a<R�a<��a<C�a<ޕa<��a<��a<��a<��a< �a<Śa<�a<�a</�a<�a<��a<,�a<ՙa<N�a<�a<��a<]�a<V�a<8�a<g�a<��a<��a<��a<��a<s�a<�a<��a<�a<��a<��a<��a<s�a<�a<�a<�a<�a<��a<�a<�a<-�a<��a<��a<��a<A�a<�a<��a<��a<�a<ڐa<��a<-�a<��a<ӎa<�a<F�a<E�a<��a<�a<S�a<�a<g�a<A�a<�a<��a<@�a<ća<�a<Q�a<y�a<3�a<��a<o�a<�a<A~a<�|a<U{a<�ya<�xa<xa<�wa<owa<�wa<�wa<xa<�xa<1ya<�ya<Eza<�za<�za<�za<Uza<�ya<zya<�xa<9xa<�wa<�va<�va<)va<�ua<�ua<�ua<�ua<�ua<"va<va<va<�ua<gua<�ta<ta<Msa< ra<qa<pa<�na<Jna<�ma<(ma<�la<4ma<�ma<gna<,oa<8pa<Vqa<�  �  ara<gsa<dta<^ua<%va<�va<wa<=wa<Uwa<Jwa<Kwa<Ewa<ewa<�wa<�wa<Hxa<�xa<Xya<�ya<�za<Y{a<�{a<_|a<�|a<�|a<�|a<*|a<�{a<m{a<�za<Qza<�ya<�ya<�ya<�ya<xza<G{a<@|a<�}a<a<ˀa<v�a<'�a<��a<�a<�a<��a<��a<_�a<ދa<U�a<��a<�a<S�a<ߍa<H�a<ގa<��a<V�a<:�a<�a<�a<��a<E�a<��a<�a<הa<��a<!�a<��a<�a<Y�a<��a<�a<��a<n�a<t�a<��a<:�a<�a<��a<�a<^�a<��a<��a<��a<��a<��a<�a<l�a<��a<��a<m�a<4�a<	�a<�a<�a<Ěa<�a<*�a<`�a<Ûa<�a<m�a<��a<ǜa<��a<U�a<Ǜa<��a<.�a<S�a<9�a<&�a<�a<C�a<y�a<$�a<�a<�a<3�a<ڔa<��a<�a<w�a<u�a<<�a<��a<��a<�a<V�a<j�a</�a<�a<s�a<	�a<��a<?�a<�a<��a<��a<��a<��a<��a<ۘa<�a<�a<��a<K�a<��a<іa<��a<��a<��a<9�a<�a<��a<��a<��a<:�a<یa<Ìa<όa<C�a<��a<s�a<�a<ŏa<6�a<��a<�a< �a<Ȑa<n�a<ȏa<�a<F�a<|�a<��a<�a<0�a<��a<;�a<��a<x�a<&�a<ۈa<s�a<�a<N�a<~�a<c�a<�a<��a<;�a<�a<~a<]|a<�za<�ya<�xa<�wa<cwa<wa<0wa<qwa<�wa<~xa<ya<�ya< za<mza<�za<�za<�za<3za<�ya<ya<sxa<�wa<Owa<�va<sva<Bva<.va<va<1va<?va<Zva<Tva<Fva<�ua<|ua<�ta<�sa<�ra<	ra<�pa<�oa<�na<�ma<ma<�la<�la<�la<2ma<�ma<�na<�oa<)qa<�  �  Fra<bsa<�ta<gua<va<�va<wa<Uwa<mwa<hwa<jwa<�wa<�wa<�wa<xa<Yxa<�xa<�ya<za<�za<j{a<	|a<G|a<�|a<�|a<�|a<W|a<�{a<O{a<�za<Eza<�ya<�ya<�ya<�ya<0za<{a<+|a<t}a<a<��a<L�a<�a<��a<c�a<l�a<��a<��a<O�a<�a<x�a<Ɍa<2�a<��a<��a<{�a<�a<��a<��a<a�a</�a<�a<��a<=�a<��a<єa<��a<̔a<4�a<��a<�a<!�a<��a<��a<s�a<D�a</�a<y�a<�a<ߑa<Ғa<�a<!�a<��a<��a<ۘa<�a<_�a<�a<U�a<��a<��a<��a<Z�a<<�a<�a<�a<��a<�a<N�a<��a<�a<-�a<��a<��a<��a<��a<;�a<śa<H�a<.�a<9�a<��a<�a<��a<�a<e�a<�a<��a<Ǔa<�a<��a<p�a<h�a<9�a<Z�a<7�a<;�a<��a<��a<J�a<R�a<G�a<��a<��a<(�a<ҙa<j�a<�a<�a<��a<Ϙa<ژa<ؘa<��a<��a<��a<��a<:�a<��a<�a<�a<��a<n�a<��a<ڐa<��a<�a<��a<�a<��a<��a<��a<�a<��a<E�a<�a<��a<A�a<�a<Րa<�a<��a<^�a<؏a<;�a<c�a<��a<܌a<�a<c�a<ъa<N�a<�a<��a<H�a<��a<}�a<��a<A�a<i�a<G�a<R�a<��a<*�a<|a<�}a<N|a<�za<|ya<zxa<�wa<wa<�va<	wa<Gwa<�wa<Axa<�xa<�ya<$za<�za<�za<�za<rza<Aza<�ya<:ya<�xa<xa<�wa<�va<�va<iva<Sva<[va<Ova<Xva<tva<lva<*va<�ua<bua<�ta<,ta<�ra<�qa<�pa<�oa<�na<�ma<ma<�la<rla<�la<ma<�ma<�na<�oa<�pa<�  �  ara<gsa<dta<^ua<%va<�va<wa<=wa<Uwa<Jwa<Kwa<Ewa<ewa<�wa<�wa<Hxa<�xa<Xya<�ya<�za<Y{a<�{a<_|a<�|a<�|a<�|a<*|a<�{a<m{a<�za<Qza<�ya<�ya<�ya<�ya<xza<G{a<@|a<�}a<a<ˀa<v�a<'�a<��a<�a<�a<��a<��a<_�a<ދa<U�a<��a<�a<S�a<ߍa<H�a<ގa<��a<V�a<:�a<�a<�a<��a<E�a<��a<�a<הa<��a<!�a<��a<�a<Y�a<��a<�a<��a<n�a<t�a<��a<:�a<�a<��a<�a<^�a<��a<��a<��a<��a<��a<�a<l�a<��a<��a<m�a<4�a<	�a<�a<�a<Ěa<�a<*�a<`�a<Ûa<�a<m�a<��a<ǜa<��a<U�a<Ǜa<��a<.�a<S�a<9�a<&�a<�a<C�a<y�a<$�a<�a<�a<3�a<ڔa<��a<�a<w�a<u�a<<�a<��a<��a<�a<V�a<j�a</�a<�a<s�a<	�a<��a<?�a<�a<��a<��a<��a<��a<��a<ۘa<�a<�a<��a<K�a<��a<іa<��a<��a<��a<9�a<�a<��a<��a<��a<:�a<یa<Ìa<όa<C�a<��a<s�a<�a<ŏa<6�a<��a<�a< �a<Ȑa<n�a<ȏa<�a<F�a<|�a<��a<�a<0�a<��a<;�a<��a<x�a<&�a<ۈa<s�a<�a<N�a<~�a<c�a<�a<��a<;�a<�a<~a<]|a<�za<�ya<�xa<�wa<cwa<wa<0wa<qwa<�wa<~xa<ya<�ya< za<mza<�za<�za<�za<3za<�ya<ya<sxa<�wa<Owa<�va<sva<Bva<.va<va<1va<?va<Zva<Tva<Fva<�ua<|ua<�ta<�sa<�ra<	ra<�pa<�oa<�na<�ma<ma<�la<�la<�la<2ma<�ma<�na<�oa<)qa<�  �  rra<�sa<�ta<}ua<va<qva<�va<�va<wa<wa<wa< wa<wa<;wa<{wa<�wa<`xa<ya<�ya<nza<({a<�{a<'|a<f|a<�|a<�|a<g|a<!|a<{a<{a<�za<>za<za<�ya<<za<�za<�{a<�|a<~a<Wa<
�a<��a<S�a<��a<>�a<��a<��a<]�a<�a<��a<�a<g�a<،a<�a<��a<�a<��a<Z�a<�a<�a<ȑa<��a<g�a<�a<r�a<��a<�a<��a<p�a<�a<)�a<��a<Ցa<r�a<��a<��a<��a< �a<��a<g�a<S�a<S�a<��a<��a< �a<��a<ՙa<��a<�a<8�a<S�a<V�a<&�a<��a<Кa<��a<��a<z�a<��a<Ԛa<�a<��a<͛a<5�a<`�a<��a<`�a<@�a<�a<(�a<��a<i�a<c�a<e�a<a�a<��a<ٔa<s�a< �a<R�a<��a<C�a<ޕa<��a<��a<��a<��a< �a<Śa<�a<�a</�a<�a<��a<,�a<ՙa<N�a<�a<��a<]�a<V�a<8�a<g�a<��a<��a<��a<��a<s�a<�a<��a<�a<��a<��a<��a<s�a<�a<�a<�a<�a<��a<�a<�a<-�a<��a<��a<��a<A�a<�a<��a<��a<�a<ڐa<��a<-�a<��a<ӎa<�a<F�a<E�a<��a<�a<S�a<�a<g�a<A�a<�a<��a<@�a<ća<�a<Q�a<y�a<3�a<��a<o�a<�a<A~a<�|a<U{a<�ya<�xa<xa<�wa<owa<�wa<�wa<xa<�xa<1ya<�ya<Eza<�za<�za<�za<Uza<�ya<zya<�xa<9xa<�wa<�va<�va<)va<�ua<�ua<�ua<�ua<�ua<"va<va<va<�ua<gua<�ta<ta<Msa< ra<qa<pa<�na<Jna<�ma<(ma<�la<4ma<�ma<gna<,oa<8pa<Vqa<�  �  �ra<�sa<�ta<uua<va<�va<�va<�va<�va<�va<�va<yva<rva<�va<�va<)wa<�wa<�xa<Aya<�ya<�za<v{a<	|a<z|a<�|a<�|a<s|a</|a<�{a<s{a<({a<�za<�za<�za<�za<w{a<@|a<0}a<{~a<�a<��a<�a<��a<�a<f�a<|�a<�a<b�a<֊a<X�a<��a<�a<2�a<��a<ʌa<^�a<��a<��a<��a<\�a<J�a<*�a<�a<��a<l�a<��a<̔a<Ӕa<j�a<�a<��a<�a<z�a<ݑa<y�a<d�a<q�a<��a<0�a<�a<ɓa<��a<��a<�a<�a<�a<�a<n�a<�a<!�a<�a<�a<��a<z�a<2�a<�a<��a<�a<�a<.�a<��a<�a<U�a<ěa<#�a<T�a<u�a<1�a<ћa<F�a<}�a<��a<Ęa<�a<�a<�a<w�a<�a<�a<�a<1�a<��a<f�a<Q�a<�a<טa<��a<<�a<��a<��a<-�a<��a<��a<=�a<��a<@�a<ǘa<L�a<�a<̗a<��a<��a<͗a<��a<�a<I�a<e�a<V�a< �a<��a<��a<	�a<�a<�a<ϒa<��a<~�a<��a<��a<,�a<ڍa<��a<��a<�a<��a<,�a<��a<&�a<}�a<�a<�a<ΐa<��a<�a<B�a<d�a<��a<��a<ًa<ߊa<F�a<��a< �a<��a<��a<d�a<"�a<�a<}�a<�a<I�a<X�a<Y�a<��a<��a<)�a<�~a<>}a<�{a<�za<�ya<�xa<Txa<xa<xa<?xa<�xa<ya<�ya<�ya<Lza<�za<�za<�za<>za<�ya<ya<^xa<�wa<wa<rva<�ua<�ua<Aua<2ua<Nua<aua<�ua<�ua<�ua<�ua<�ua<Xua<�ta<*ta<Hsa<era<mqa<�pa<�oa<�na<na<�ma<�ma<�ma<1na<�na<�oa<�pa<�qa<�  �  `sa<ta<�ta<�ua<�ua<Gva<>va<mva<1va<$va<�ua<�ua<�ua<�ua<>va<ova<7wa<�wa<�xa<�ya<Mza<{a<�{a<J|a<�|a<�|a<�|a<�|a<k|a<�{a<�{a<d{a<S{a<V{a<�{a<9|a<�|a<�}a<#a<��a<�a<w�a<�a<;�a<��a<��a<l�a<�a<��a<�a<&�a<|�a<b�a<ߋa<�a<��a<C�a<ۍa<�a<��a<Րa<��a<��a<k�a<�a<��a<Дa<�a<��a<��a<�a<c�a<�a<��a<@�a<�a<3�a<q�a<�a<��a<w�a<��a<a�a<��a<��a<I�a<�a<h�a<ƚa<��a<��a<��a<>�a<�a<]�a<h�a<�a<5�a<+�a<��a<Ιa<5�a<�a<B�a<ʛa<�a<1�a<�a<�a<��a<Ӛa<M�a<6�a<X�a<��a<ʖa<5�a<��a<��a<��a<�a<m�a<
�a<��a<r�a<u�a<�a<��a<ؚa<�a<�a<��a<^�a<��a<M�a<��a<��a<��a<$�a<�a<͖a<�a<��a<g�a<��a<ڗa<�a<�a<�a<��a<�a<Q�a<t�a<��a<6�a<B�a<-�a<J�a<v�a<�a<��a<[�a<��a<��a<6�a<��a<�a<��a<̐a<�a<�a<��a<E�a<��a<�a<�a<�a<ыa<!�a</�a<��a<��a<l�a<J�a<ɇa<�a<��a<��a<)�a<��a<3�a<\�a<��a<9�a<�a<��a<a<�}a<j|a<I{a<Aza<�ya<ya<�xa<�xa<�xa<Iya<�ya<za<fza<�za<�za<�za<gza<�ya<\ya<�xa<�wa<.wa<1va<�ua<ua<�ta<�ta<�ta<�ta<�ta<ua</ua<~ua<hua<�ua<Cua<�ta<rta<�sa<sa<�qa<�pa<*pa<hoa<�na<rna<yna<}na<�na<�oa<Xpa<:qa<$ra<�  �  �sa<nta<ua<�ua<�ua<va<va<�ua<�ua<Pua<ua<�ta<�ta<�ta<)ua<�ua<Iva<
wa<�wa<�xa<�ya<�za<r{a<|a<�|a<�|a<�|a<�|a<�|a<�|a<]|a<3|a<%|a<?|a<�|a<}a<�}a<�~a<�a<E�a<��a<��a<I�a<��a<��a<��a<[�a<ىa<8�a<w�a<p�a<��a<Ȋa<��a<?�a<��a<:�a< �a<��a<�a<�a<��a<(�a<�a<ݓa<��a<�a<��a<�a<˔a<{�a<2�a<��a<a�a<1�a<�a<�a<b�a<ԓa<��a<L�a<*�a<$�a<��a<Әa<��a<�a<{�a<��a<��a<X�a<��a<n�a<)�a<��a<w�a<�a<(�a<5�a<��a<�a<��a<�a<��a<L�a<��a<��a<�a<��a<��a<5�a<�a<ϙa<�a<R�a<��a<#�a<a<��a<��a<ܖa<B�a<їa<{�a<�a<��a<C�a<��a<ޚa<�a<��a<_�a<�a<&�a<y�a<ܗa<C�a<��a<3�a<
�a<�a< �a<U�a<��a<ۖa<M�a<��a<��a<×a<��a<�a<��a<Ǖa<הa<�a<�a<��a<�a<_�a<ڏa<~�a<X�a<w�a<��a<�a<W�a<��a<�a<4�a<�a<�a<��a<
�a<G�a<b�a<4�a<N�a<6�a<@�a<T�a<��a<��a<��a<^�a<-�a<+�a<�a<�a<ֆa<��a<�a<r�a<~�a<��a<V�a<�a<�a<~~a<D}a<:|a<8{a<�za<za<�ya<�ya<�ya<�ya<Eza<sza<�za<�za<�za<�za<Cza<�ya<�xa<!xa<wa<hva<�ua<�ta<*ta<�sa<�sa<�sa<�sa<�sa<Eta<�ta< ua</ua<Jua<>ua<�ta<�ta<�sa<6sa<wra<�qa<�pa<Bpa<�oa<uoa<]oa<�oa<�oa<fpa<qa<�qa<�ra<�  �  ta<�ta<Dua<�ua<�ua<�ua<�ua<Iua<"ua<�ta<Gta<�sa<�sa<�sa<4ta<�ta<Dua<"va<wa<'xa<=ya<za<6{a<�{a<�|a<�|a<:}a<P}a<4}a<M}a<}a<
}a<�|a<0}a<�}a<~a<�~a<�a<ހa<�a<_�a<��a<��a<��a<��a<��a<�a<��a<��a<ԉa<�a<݉a<��a<��a<I�a<��a<L�a<�a<��a<�a<7�a<��a<��a<��a<��a<8�a<�a<�a<l�a<1�a<�a<�a<��a<D�a<�a<�a<�a<Z�a<Ȕa<X�a<(�a<�a<ٗa<y�a<6�a<ۙa<�a<n�a<R�a<R�a<��a<o�a<�a<K�a<ٗa<q�a<A�a<4�a<Z�a<��a<�a<��a<]�a</�a<��a<R�a<��a<�a<�a<ɛa<��a<�a<��a<ϙa<�a<��a< �a<��a<��a<��a<��a<"�a<��a<.�a<љa<�a<��a<՚a<�a<Ța<v�a<�a<:�a<��a<͗a<�a<K�a<��a<[�a<�a<�a<�a<m�a<Ǖa<M�a<ɖa<��a<��a<t�a<}�a<(�a<Жa<-�a<R�a<��a<��a<Ғa<��a<P�a<ِa<��a<W�a<N�a<{�a<��a<�a<A�a<L�a<��a<>�a<�a<a�a<Ϗa<ˎa<��a<Ča<w�a<f�a<@�a<^�a<��a<�a<��a<^�a<Y�a<P�a<z�a<e�a<L�a<O�a<υa<o�a<��a<�a<��a<��a<��a<Ca<&~a<}a<7|a<�{a<�za<�za<�za<�za<�za<�za<�za<{a<${a<�za<�za<�ya<oya<[xa<�wa<�va<�ua<�ta<�sa<Msa<�ra<�ra<�ra<�ra<&sa<�sa<ta<Wta<�ta<
ua<ua<ua<�ta<jta<�sa<+sa<mra<�qa<%qa<�pa<spa<Ypa<�pa<�pa<Eqa<�qa<�ra<�sa<�  �  �ta<)ua<�ua<�ua<�ua<�ua<Qua<�ta<kta<�sa<ysa< sa<�ra<�ra<9sa<�sa<hta<>ua<Iva<xwa<�xa<�ya<�za<�{a<||a<}a<x}a<�}a<�}a<�}a<�}a<�}a<�}a<0~a<s~a<a<�a<��a<��a<�a<��a<,�a<D�a<1�a<�a<��a<��a<X�a<X�a<J�a<L�a< �a<�a<)�a<S�a<��a<R�a<�a<$�a<9�a<s�a<̏a<��a<)�a<Y�a<�a<�a<l�a<��a<��a<��a<]�a<]�a<�a<�a<�a<�a<A�a<ĕa<X�a<��a<��a<J�a<�a<��a<�a<^�a<g�a<&�a<�a<Z�a<Řa<:�a<��a<��a<��a<D�a<2�a<X�a<��a<3�a<�a<��a<v�a<*�a<�a<~�a<қa<�a<�a<��a<��a<�a<d�a<��a<r�a<�a<��a<��a<w�a<��a<�a<u�a<ҙa<H�a<Ěa<��a<�a<�a<��a<B�a<��a<Řa<��a<�a<6�a<m�a<˔a<Z�a<�a<�a<?�a<��a<�a<��a<�a<��a<�a<H�a<u�a<]�a<�a<��a<��a<�a<k�a<��a<��a<Q�a<��a<r�a<5�a<O�a<W�a<��a<��a<ґa<�a<a<��a<�a<G�a<��a<h�a<5�a<�a<��a<��a<k�a<h�a<��a<�a<��a<��a<w�a<��a<Åa<΅a<�a<�a<��a<v�a<�a<%�a<J�a<F�a<�a< �a<�~a<~a<}a<p|a<�{a<�{a<�{a<q{a<~{a<j{a<�{a<�{a<b{a<{a<�za<�ya<ya<�wa<�va<�ua<�ta<�sa<sa<Qra<�qa<�qa<�qa<�qa<Sra<�ra<csa<�sa<jta<�ta<�ta<ua<�ta<�ta<Cta<�sa<sa<�ra<ra<�qa<Hqa<Lqa<Wqa<�qa<8ra<�ra<Nsa<�sa<�  �  (ua<Tua<�ua<�ua<�ua<wua<�ta<�ta<�sa<6sa<�ra<Nra<
ra<�qa<Vra<�ra<zsa<eta<�ua<�va<�wa<uya<iza<�{a<k|a<}a<�}a<�}a<^~a<f~a<�~a<�~a<�~a<a<la<�a<��a<��a<Z�a<��a<��a<��a<��a<]�a<0�a<��a<�a<�a<�a<�a<��a<x�a<A�a<L�a<c�a<͈a<i�a<$�a<;�a<a�a<ȍa<��a<��a<�a<��a<#�a<Ԕa<��a<ҕa<�a<8�a<�a< �a<��a<��a<ŕa<�a<B�a<��a<3�a<��a<�a<��a<��a<�a<S�a<l�a<P�a<&�a<��a<!�a<>�a<m�a<іa<!�a<��a<E�a<P�a<]�a<a<b�a<�a<��a<��a<�a<��a<H�a<ӛa<�a<F�a<	�a<��a<��a<8�a<��a<�a<�a<�a<��a<e�a<��a<șa<+�a<��a<ޚa<=�a<*�a<M�a<�a<��a<�a<D�a<��a<L�a<_�a<l�a<��a<�a<Y�a<6�a<�a<P�a<��a<C�a<Ԕa<��a<b�a<��a<?�a<d�a<e�a<G�a<ϖa<|�a<a<9�a<L�a<��a<4�a<��a<}�a<�a<B�a<��a<O�a<U�a<[�a<C�a<�a<��a<�a<Q�a<3�a<�a<،a<G�a<�a<��a<��a<y�a<��a<%�a<��a<��a<��a<�a<��a<f�a<��a<��a<��a<`�a<
�a<W�a<��a<ςa<Ɂa<�a<�a<�~a<�}a<x}a<�|a<�|a<]|a<|a<H|a<|a<&|a<�{a<�{a<#{a<zza<�ya<�xa<�wa<cva<ua<ta<�ra<ra<Rqa< qa<�pa<�pa<qa<�qa<"ra<�ra<�sa<ta<�ta<�ta<ua<)ua<�ta<�ta<8ta<�sa<Nsa<�ra<�ra<2ra<bra<Era<�ra<�ra<xsa<"ta<�ta<�  �  ~ua<�ua<�ua<�ua<�ua<,ua<�ta<�sa<Rsa<�ra<ra<�qa<Lqa<Nqa<�qa<	ra<�ra<�sa<�ta<Lva<�wa<�xa<za<W{a<S|a<2}a<�}a<X~a<�~a<�~a<a<Ea<�a<�a<*�a<ˀa<V�a<S�a<0�a</�a<�a<�a< �a<·a<S�a<��a<ވa<��a<��a<d�a<#�a<�a<��a<��a<��a<�a<��a<y�a<q�a<��a<9�a<��a<�a<w�a<��a<��a<єa<��a<6�a<n�a<��a<��a<��a<��a<��a<|�a<Ėa<��a<O�a<�a<b�a<�a<y�a<��a<I�a<��a<��a<C�a<�a<7�a<��a<Ηa<�a<3�a<u�a<�a<��a<��a<��a<�a<��a<h�a<x�a<W�a<G�a</�a<��a<��a<�a<|�a<y�a<V�a<�a<��a<N�a<�a<��a<;�a<J�a<#�a<X�a<��a<֚a<�a<Z�a<��a<��a<��a<�a<��a<ҙa<�a<�a<�a<�a<Ŕa<ޓa<$�a<��a<l�a<f�a<��a<�a<��a<p�a<�a<Ǖa<a�a<��a<M�a<{�a<��a<4�a<Ԗa<E�a<��a<�a<��a<�a<n�a<.�a<Ғa<�a<͒a<Ւa<ƒa<��a<��a<_�a<ӑa<�a<.�a<�a<��a<O�a<�a<��a<�a<Ɇa<Åa<�a<c�a<
�a<؃a<�a<S�a<��a<�a<5�a<X�a<��a<]�a<�a<��a<��a<+�a<@�a<^�a<m�a<�a<�~a<-~a<�}a<2}a<}a<�|a<�|a<�|a<{|a<*|a<�{a<7{a<mza<�ya<Uxa<3wa<�ua<�ta<tsa<Jra<Sqa<�pa<<pa<pa<pa<Zpa<�pa<�qa<Dra<�ra<�sa<Ota<�ta<ua<_ua<Cua<ua<�ta<Cta<�sa<�sa<=sa<�ra<sa<sa<Vsa<�sa<#ta<�ta<ua<�  �  �ua<�ua<�ua<�ua<�ua<ua<�ta<�sa<�ra<0ra<�qa<qa<�pa<�pa<�pa<dqa<ra<Hsa<Yta<�ua<$wa<�xa<za<5{a<o|a<A}a<�}a<�~a<�~a<Ya<�a<�a<�a<m�a<݀a<c�a<'�a<ɂa<΃a<��a<��a<��a<<�a<߇a<K�a<��a<Èa<��a<��a<�a<��a<G�a< �a<�a<�a<W�a<�a<׈a<�a<I�a<��a<5�a<��a<I�a<��a<Փa<�a<��a<?�a<��a<��a<	�a<�a<.�a<�a<I�a<`�a<��a<�a<]�a<�a<i�a<�a<G�a<��a<��a<��a<a�a<řa<D�a<[�a<f�a<��a<��a<�a<M�a<��a<Ɠa<�a<`�a<*�a<�a<ۖa<��a<��a<%�a<�a<��a<1�a<b�a<��a<��a<t�a<�a<ٛa<��a<#�a<�a<ٚa<�a<�a<"�a<h�a<��a<ɛa<ța<ța<r�a<+�a<��a<��a<�a<��a<��a<X�a<C�a<j�a<��a<�a<��a<��a<��a<��a<�a<�a<��a<��a<i�a<ږa<h�a<��a<y�a<r�a<�a<��a<�a<��a<��a<��a<!�a<Ɠa<��a<X�a<k�a<S�a<<�a<&�a<ےa<q�a<ˑa<�a<�a<�a<��a<�a<��a<�a<��a<H�a<!�a<?�a<��a<g�a<W�a<��a<��a<-�a<��a<�a<Z�a<m�a<�a<%�a<Ąa<;�a<��a<��a<ہa<�a<�a<~a<�~a<L~a<�}a<�}a<|}a<2}a<	}a<�|a<o|a<�{a<E{a<�za<gya<bxa<�va<�ua<?ta<�ra<�qa<�pa<pa<voa<[oa<foa<�oa<^pa<qa<�qa<�ra<�sa<>ta<�ta<3ua<Fua<dua<Aua<ua<�ta<sta< ta<�sa<�sa<�sa<�sa<�sa<Eta<�ta<ua<zua<�  �  �ua<-va< va<�ua<�ua<�ta<Gta<�sa<�ra<�qa<5qa<�pa<Npa<^pa<�pa<qa<�qa<�ra<ta<�ua<�va<xa<�ya<{a<O|a<[}a<$~a<�~a<5a<�a<�a<�a<P�a<a<%�a<��a<y�a<)�a<�a<�a<܅a<��a<}�a<�a<��a<��a<��a<p�a<B�a<�a<�a<�a<ǆa<��a<��a<�a<��a<��a<��a<�a<W�a<��a<��a<�a<d�a<��a<�a<ѕa<q�a<�a<(�a<Q�a<Z�a<f�a<i�a<��a<��a<�a<_�a<��a<;�a<��a<+�a<��a<Κa<Кa<��a<B�a<��a<�a<4�a<>�a<N�a<[�a<��a<�a<��a<��a<��a<
�a<Ɣa<��a<��a<a<�a<ڙa<��a<��a<6�a<��a<՜a<Ҝa<��a<b�a<�a<Ûa<��a<W�a<&�a<2�a<I�a<e�a<��a<͛a<��a<�a<�a<��a<7�a<|�a<��a<��a<��a<Q�a<�a<�a<�a<%�a<��a<p�a<r�a<��a<+�a<͒a<��a<��a<l�a<�a<��a<G�a<��a<��a<��a<T�a<�a<c�a<�a<G�a<�a<j�a<�a<��a<��a<��a<��a<��a<W�a<�a<��a<�a<�a<�a<��a<R�a<܋a<B�a<��a<6�a<�a<τa<�a<h�a<�a<��a<*�a<p�a<�a<i�a<Єa<�a<M�a<m�a<V�a<��a<z�a<��a<��a<�a<H�a<q�a<�a<a<�~a<B~a<�}a<�}a<v}a<K}a<�|a<�|a<|a<f{a<lza<Aya<xa<�va<dua<�sa<�ra<tqa<^pa<�oa<>oa<oa<oa<~oa<pa<�pa<�qa<�ra<Zsa<ta<�ta<8ua<�ua<�ua<�ua<Mua< ua<�ta<`ta<&ta<	ta<�sa<ta<Gta<�ta<�ta<Hua<�ua<�  �  /wa<Nwa<]wa<<wa<wa<�va<+va<�ua<ua<�ta<#ta<�sa<�sa<�sa<�sa<<ta<�ta<�ua<�va<xa<4ya<�za<�{a<�|a<�}a<�~a<La<�a<Q�a<ŀa<#�a<��a<�a<0�a<��a<d�a<Ѓa<��a<r�a<4�a<�a<��a<[�a<��a<j�a<��a<�a<
�a<�a<Éa<i�a<i�a<I�a<?�a<��a<ˉa<]�a<A�a<&�a<S�a<��a<ďa<9�a<��a<��a<�a<��a<l�a<�a<s�a<��a<�a<3�a<b�a<}�a<��a<�a<&�a<[�a<љa<6�a<��a<�a<&�a<^�a<��a<`�a<5�a<��a<G�a<��a<�a<G�a<��a<�a<��a<\�a<B�a<f�a<Җa<O�a<
�a<טa<��a<��a<D�a<!�a<��a<�a<[�a<w�a<��a<i�a<K�a<"�a<�a<��a<s�a<��a<Y�a<l�a<��a<��a<��a<Ȝa<Ĝa<��a<p�a<�a<��a<��a<��a<.�a<�a<L�a<g�a<��a<��a<q�a<4�a<&�a<Z�a<��a<1�a<��a<P�a< �a<v�a<�a<O�a<e�a<x�a<J�a<	�a<��a<T�a<�a<w�a<�a<��a<k�a<�a<הa<��a<��a<\�a<�a<��a<P�a<��a<�a<*�a<�a<Ўa<��a<�a<�a<��a<~�a<��a<��a<+�a<�a<��a<��a<�a<�a<M�a<��a<��a<Ɇa<��a<I�a<��a<^�a<��a<,�a<`�a<��a<�a<0�a<΀a<=�a<�a<pa<#a<�~a<�~a<~a<�}a<D}a<�|a<�{a<{a<�ya<�xa<�wa<sva<nua<fta<�sa<�ra<qra<>ra<Xra<�ra<�ra<�sa<�sa<�ta<Fua<�ua<\va<�va<�va<�va<�va<�va<nva<Bva<va<�ua<�ua<�ua<�ua<�ua<8va<va<�va<�va<�  �  4wa<cwa<fwa<Zwa< wa<�va<-va<�ua<0ua<�ta<)ta<�sa<�sa<�sa<�sa<nta<ua<�ua<�va<xa<Mya<sza<�{a<�|a<�}a<�~a<Ka<�a<Y�a<��a<�a<f�a<��a<!�a<��a<�a<˃a<|�a<N�a<�a<�a<Ça<q�a<�a<z�a<щa<։a<�a<Ӊa<��a<��a<n�a<f�a<a�a<��a<�a<��a<\�a<C�a<r�a<��a<��a<8�a<o�a<��a<��a<��a<|�a<�a<��a<ݗa<�a<�a<B�a<P�a<��a<��a<�a<N�a<��a<�a<u�a<�a<8�a<v�a<|�a<p�a<<�a<��a<?�a<��a<�a<f�a<��a<8�a<��a<��a<|�a<��a<�a<p�a<�a<֘a<��a<��a<B�a<�a<��a<"�a<g�a<��a<��a<s�a<:�a<�a<��a<��a<`�a<;�a<A�a<N�a<[�a<��a<��a<Μa<ɜa<��a<y�a<$�a<}�a<a<��a<(�a<E�a<L�a<n�a<��a<�a<��a<c�a<X�a<s�a<єa<7�a<ϕa<j�a<�a<q�a<ۗa<G�a<y�a<w�a<`�a<�a<��a<<�a<˖a<A�a<�a<w�a<�a<�a<��a<��a<j�a<K�a< �a<ʓa<W�a<��a<�a<��a<�a<��a<��a<H�a<��a<ˉa<��a<��a<�a<p�a<�a<ʅa<مa<�a<!�a<L�a<o�a<��a<��a<��a<X�a<�a<v�a<ׄa<�a<D�a<��a<ǁa<+�a<��a<�a<�a<=a<a<�~a<~a</~a<�}a<?}a<�|a<�{a<�za<�ya<�xa<�wa<�va<uua<�ta<�sa<sa<�ra<|ra<mra<�ra<sa<�sa<&ta<�ta<Dua<�ua<8va<�va<�va<�va<�va<�va<^va<"va<�ua<�ua<�ua<�ua<�ua<�ua<va<cva<�va< wa<�  �  �va<?wa<@wa<Kwa<wa<�va<�va<�ua<cua<�ta<`ta<ta<�sa<�sa< ta<�ta<Iua<=va<!wa<Gxa<wya<�za<�{a<�|a<�}a<�~a<#a<�a<�a<��a<рa<5�a<m�a<�a<b�a<ނa<��a<3�a<�a<�a<��a<��a<3�a<؈a<S�a<̉a<�a<+�a<�a<Չa<Ӊa<��a<��a<��a<Ήa<D�a<Њa<��a<��a<��a<a<,�a<U�a<��a<�a<��a<��a<Y�a<�a<R�a<��a<ŗa<��a<�a<�a<U�a<o�a<��a<�a<^�a<�a<D�a<��a<��a<H�a<X�a<Y�a<<�a<ښa<��a<יa<8�a<��a<�a<|�a<��a<��a<��a<ۖa<�a<��a<P�a<��a<�a<��a<��a<(�a<��a<�a<<�a<k�a<O�a<D�a<��a<Ӝa<}�a<F�a<5�a<�a<�a<�a<�a<d�a<r�a<��a<��a<��a<S�a<�a<��a<��a<W�a<C�a<x�a<w�a<��a<��a<A�a<��a<��a<��a<��a<�a<j�a<��a<��a<�a<Ǘa< �a<O�a<g�a<O�a<5�a<ԗa<��a<�a<��a<�a<��a<H�a<�a<��a<l�a<_�a<A�a<�a<�a<��a<)�a<��a<��a<�a<2�a<�a<��a<�a<�a<�a<�a<�a<7�a<��a<3�a<�a<�a<
�a<Y�a<i�a<��a<ކa<��a<��a<6�a<Ʌa<=�a<��a<Ճa< �a<Z�a<~�a<��a<K�a<�a<ra<�~a<�~a<�~a<E~a<�}a<�}a<}a<�|a<�{a<�za<*za<�xa<�wa<�va<�ua<�ta<�sa<Ksa<�ra<�ra<�ra<�ra<@sa<�sa<Yta<�ta<�ua<�ua<Hva<�va<�va<�va<�va<qva<#va<�ua<�ua<pua<mua<Qua<|ua<�ua<�ua<3va<pva<�va<�  �  �va<#wa<Owa<2wa<wa<�va<wva<va<�ua<5ua<�ta<�ta<kta<qta<�ta<(ua<�ua<�va<�wa<�xa<�ya<�za<�{a<�|a<�}a<�~a<3a<�a<�a<I�a<��a<��a<�a<^�a<ρa<n�a<��a<�a<��a<��a<p�a<L�a<�a<ވa<b�a<��a<�a<�a<(�a<1�a<�a<
�a<��a<#�a<d�a<��a<J�a<!�a<�a<�a<;�a<d�a<��a<ɒa<֓a<�a<��a<g�a<��a<*�a<j�a<��a<��a<��a<×a<��a<��a<2�a<��a<�a<_�a<��a<n�a<Қa< �a<j�a<[�a<1�a<�a<{�a<�a<��a<�a<U�a<Ηa<{�a<F�a<)�a<S�a<��a<�a<��a<s�a<(�a<�a<��a<+�a<��a<��a<I�a<V�a<,�a<��a<��a<b�a<�a<�a<��a<��a<y�a<��a<Ûa<�a<#�a<W�a<i�a<y�a<a�a<��a<��a<�a<J�a<��a<��a<�a<�a<W�a<͕a<[�a<�a<�a<0�a<l�a<וa<T�a<ݖa<W�a<��a<&�a<N�a<_�a<_�a<�a<��a<@�a<��a<�a<��a<�a<��a<t�a< �a<!�a<��a<�a<˓a<��a<h�a</�a<��a<�a<5�a< �a<�a<��a<��a<��a<]�a<c�a<~�a<��a<�a<ˆa<��a<k�a<��a<��a<��a<Ɇa<Ɔa<ӆa<��a<C�a<؅a<�a<e�a<��a<΂a<ԁa<:�a<Y�a<�a<Ha<�~a<�~a<L~a<;~a<~a<�}a<{}a<-}a<�|a<�{a<{a<za<*ya<$xa<wa<va< ua<gta<�sa<Xsa<*sa<2sa<Rsa<�sa<ta<�ta<&ua<�ua<�ua<eva<�va<�va<�va<fva<)va<�ua<�ua<:ua<ua<�ta<�ta<�ta<,ua<iua<�ua<!va<�va<�  �  �va<�va<wa<"wa</wa<wa<�va<|va<�ua<�ua<Dua<ua<�ta<�ta<Iua<�ua<\va<wa<xa<ya<za<1{a<|a<}a<�}a<e~a<�~a<Da<�a<�a<1�a<1�a<��a<�a<G�a<�a<l�a<t�a< �a<'�a<�a<��a<͇a<��a<;�a<��a<:�a<D�a<k�a<��a<f�a<��a<s�a<��a<܊a<C�a<݋a<��a<��a<��a<a<Đa<�a<�a<�a<�a<��a<C�a<��a<�a<�a<�a<6�a<�a<N�a<(�a<r�a<��a<�a<��a<ؘa<��a<�a<��a<ɚa<�a<>�a<2�a<.�a<��a<f�a<ؙa<H�a<ݘa<O�a<�a<a<ʗa<ԗa<.�a<��a<-�a<�a<z�a<R�a<Ûa<]�a<Ӝa<�a<�a<��a<�a<��a<[�a<�a<|�a<q�a<�a<�a<�a<-�a</�a<r�a<қa<�a<$�a<�a<-�a<�a<��a<6�a<z�a<�a<�a<O�a<��a<ږa<V�a<ڕa<��a<��a<��a<�a<Z�a<��a<+�a<��a<�a<Q�a<N�a<E�a<�a<��a<e�a<a<a�a<��a<'�a<��a<-�a<�a<��a<��a<I�a<{�a<_�a<M�a<&�a<Ւa<��a<ܑa<Y�a<K�a<V�a<b�a<�a<�a<؊a<��a<��a<7�a<��a<C�a<�a<�a<
�a<��a<%�a<�a<�a<��a<|�a< �a<}�a<̄a<�a<"�a<b�a<B�a<ŀa<�a<Ma<�~a<_~a<0~a<�}a<�}a<�}a<z}a<#}a<�|a<o|a<�{a<I{a<Hza<�ya<yxa<twa<�va<�ua<�ta<Lta<�sa<�sa<�sa<�sa<ta<�ta<�ta<�ua<�ua<0va<}va<tva<�va<Hva<va<�ua<ua<ua<�ta<�ta<>ta<Zta<Nta<�ta<�ta<Aua<�ua<va<�  �  ?va<�va<�va<0wa<-wa<.wa< wa<�va<wva<va<�ua<�ua<�ua<�ua<�ua<]va< wa<�wa<�xa<�ya<{za<U{a<f|a<}a<�}a<g~a<�~a<a<Ua<Pa<�a<�a<�a<3�a<��a<,�a<сa<��a<��a<��a<n�a<��a<��a<\�a<�a<��a<"�a<��a<��a<Ŋa<�a<��a<�a<I�a<��a<�a<��a<I�a</�a<+�a<'�a<Q�a<O�a<U�a<d�a<��a<��a<#�a<p�a<��a<��a<��a<��a<�a<r�a<��a<��a<��a<_�a<��a<g�a< �a<o�a<+�a<��a<�a<5�a<F�a<$�a<�a<��a<9�a<יa<S�a<��a<��a<u�a<p�a<��a<�a<H�a<Ǚa<V�a<�a<v�a<�a<��a<ǜa<�a<�a<לa<��a<'�a<��a<t�a<�a<��a<k�a<U�a<J�a<h�a<��a<��a<1�a<r�a<ԛa<��a< �a<��a<��a<X�a<Қa<�a<��a<̘a<�a<��a< �a<��a<Y�a<H�a<d�a<��a<ߖa<G�a<��a<֗a<E�a<U�a<]�a<G�a<�a<��a<�a<G�a<��a<&�a<h�a<�a<z�a<3�a<�a<Ӓa<Вa<�a<ɒa<�a<�a<��a<W�a<�a<A�a<��a<��a<��a<��a<y�a<��a<��a<��a<��a<f�a<�a<��a<��a<o�a<}�a<d�a<U�a<T�a<�a<��a< �a<Q�a<��a<��a<��a<ҁa<΀a<�a<1a<�~a<~a<�}a<^}a<T}a<?}a<}a<"}a<�|a<�|a<f|a<�{a<?{a<�za<�ya<�xa<xa<wa<Lva<�ua< ua<�ta<ita<fta<�ta<�ta<ua<qua<�ua<va<gva<qva<�va<Zva<&va<�ua<Tua<�ta<�ta<ta<�sa<�sa<�sa<�sa<�sa<>ta<�ta</ua<�ua<�  �  �ua<qva<�va<"wa<Lwa<Ewa<Swa<wa<wa<�va<rva<Sva<Kva<ova<�va<(wa<�wa<gxa<#ya<za<{a<�{a<�|a<0}a<�}a<C~a<�~a<�~a<�~a<a<�~a<a<1a<�a<�a<c�a</�a<�a<�a<܃a<�a<7�a<�a<?�a<�a<ىa<8�a<Ȋa<�a<K�a<��a<s�a<ŋa<�a<Y�a<��a<H�a<�a<Ύa<ԏa<��a<��a<Ӓa<��a<��a<�a<ؕa<��a<U�a<A�a<Q�a<6�a<�a<�a<Õa<�a<��a<:�a<��a<�a<Ηa<O�a<9�a<��a<N�a<Κa<	�a<i�a<9�a<T�a<�a<Ța<R�a<ߙa<��a<K�a<E�a<#�a<M�a<��a<�a<h�a<њa<��a<�a<l�a<��a<�a<�a<��a<��a<&�a<�a<6�a<��a<W�a<�a<��a<��a<��a<��a<��a<G�a<��a<5�a<b�a<ƛa<ʛa<�a<ɛa<o�a<%�a<��a<�a<C�a<��a<*�a<��a<X�a<
�a<�a<�a<@�a<m�a<��a<+�a<<�a<��a<i�a<��a<$�a<ȗa<K�a<��a<�a<�a<��a<Ǔa<H�a<Œa<j�a<Q�a<�a<7�a<0�a<l�a<��a<t�a<��a<)�a<�a<W�a<ϐa<�a<�a<6�a<��a<*�a<#�a<s�a<��a<�a<��a<U�a<:�a<�a<�a<�a<��a<��a<��a<��a<ԅa<6�a<,�a<L�a<F�a<�a<9�a<:a<�~a<�}a<P}a<}a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<:|a<|a<T{a<�za<za<hya<~xa<�wa<�va<6va<�ua<Qua<$ua<ua<ua<Xua<~ua<va<&va<ova<�va<�va<�va<$va<�ua<aua<ua<Zta<�sa<zsa<sa<�ra<�ra<�ra<2sa<�sa<ta<�ta<gua<�  �  dua< va<�va<wa<_wa<ywa<�wa<�wa<@wa<.wa<#wa<�va<�va< wa<qwa<�wa<Yxa<ya<�ya<|za<V{a<+|a<�|a<c}a<�}a<,~a<|~a<�~a<j~a<�~a<k~a<x~a<�~a<�~a<'a<�a<_�a<E�a<H�a<T�a<��a<��a<��a<��a<Јa<��a<f�a<�a<Y�a<��a<ŋa<)�a<]�a<��a< �a<q�a<
�a<��a<z�a<h�a<g�a<)�a<:�a<�a<��a<E�a<��a<ޕa<�a<�a<̕a<��a<`�a<B�a<"�a<�a<B�a<��a<�a<~�a<%�a<͗a<��a<:�a<��a<��a<��a<U�a<h�a<s�a<]�a<�a<��a<��a<;�a<�a<�a<�a<��a<C�a<��a<�a<v�a<̛a<\�a<��a<ܜa<��a<ߜa<��a<^�a<��a<O�a<Ěa<,�a<��a<E�a<��a<Ϙa<֘a<�a<S�a<��a<)�a<��a<��a<v�a<��a<͛a<ܛa<��a<_�a<��a<V�a<ޙa<h�a<ɘa<a�a<
�a<ޗa<��a<��a<ۗa<)�a<2�a<t�a<��a<��a<��a<z�a<�a<��a<��a<"�a<z�a<��a<ޓa<+�a<��a<�a<��a<��a<}�a<��a<��a<�a<�a<�a<P�a<�a<�a<��a<�a<D�a<��a<q�a<��a<��a<ˋa<�a<e�a<ىa<f�a<�a<ψa<��a<V�a<N�a<�a<��a<*�a<��a<��a< �a<׃a<ǂa<��a<��a<�a<�~a<�}a<}a<�|a<L|a<|a<|a<|a<7|a<1|a<T|a<j|a<&|a<�{a<�{a<{a<wza<�ya<�xa<[xa<�wa<�va<rva<va<�ua<�ua<�ua<va<"va<;va<�va<�va<�va<�va<eva<va<�ua<�ta<|ta<�sa<Msa<�ra<pra<,ra<ra<;ra<�ra<�ra<�sa<(ta<�ta<�  �  <ua<�ua<�va<�va<Twa<�wa<�wa<�wa<�wa<�wa<�wa<�wa<�wa<�wa<*xa<lxa<-ya<�ya<^za<{a<�{a<v|a<�|a<�}a<�}a<<~a<=~a</~a<F~a<�}a<�}a<�}a<�}a<~a<i~a<a<�a<��a<��a<�a< �a<S�a<��a<��a<ވa<��a<t�a<�a<��a<�a<E�a<ƌa<Όa<d�a<��a<(�a<a<Z�a<V�a<ܐa<��a<��a<��a<=�a<ܔa<`�a<��a<�a<��a<��a<��a<�a<��a<��a<��a<k�a<��a<Ȕa<=�a<ԕa<�a<d�a<�a<�a<��a<U�a<�a<=�a<��a<��a<��a<~�a<R�a<$�a<��a<ښa<��a<��a<��a<��a<=�a<��a<�a<G�a<��a<՜a<�a<��a<Ԝa<��a<��a<��a<ܚa<9�a<��a<�a<��a<8�a<+�a<�a<`�a<��a<�a<��a<%�a<Кa<�a<��a<ța<Лa<Лa<��a<J�a<˚a<~�a<ۙa<i�a<#�a<��a<��a<W�a<��a<_�a<��a<Әa<ߘa<��a<٘a<ǘa<d�a<�a<j�a<��a<��a<�a<,�a<@�a<~�a<ۑa<O�a<�a<Ґa<ڐa<�a<9�a<[�a<��a<�a<�a<#�a<ӑa<��a<�a<v�a<ۏa<��a<O�a<2�a<��a<��a<�a<��a<�a<݉a<B�a<F�a<܈a<��a<=�a<̇a<E�a<y�a<Ѕa<��a<��a<��a<.�a<'�a<�~a<�}a<}a<h|a<�{a<�{a<t{a<l{a<�{a<�{a<|a<|a<|a<;|a<�{a<�{a<2{a<�za<za<~ya<�xa<xa<�wa<wa<�va<�va<�va<tva<qva<�va<�va<�va<�va<�va<�va<[va<va<Kua<�ta<	ta<]sa<�ra<*ra<�qa<qqa<wqa<~qa<�qa<Ora<�ra<�sa<Xta<�  �  �ta<�ua<[va<�va<gwa<�wa<	xa<xa<+xa<xa<xa<$xa<<xa<Rxa<�xa<�xa<�ya<!za<�za<v{a<%|a<�|a<X}a<�}a<�}a< ~a<~a<�}a<�}a<�}a<�}a<`}a<f}a<�}a<�}a<f~a<3a<�a<�a<Z�a<��a<��a<@�a<j�a<��a<��a<��a<f�a<�a<`�a<ǌa<(�a<X�a<�a<"�a<��a<F�a<�a<ΐa<l�a<i�a<,�a<�a<��a<6�a<��a<��a<ȕa<��a<e�a< �a<��a<q�a<�a<��a<�a<��a<C�a<a<U�a<�a<�a<��a<��a<o�a<*�a<�a<E�a<��a<��a<�a<ܛa<��a<��a<Q�a<Q�a<�a<1�a<9�a<s�a<ʛa<�a<f�a<a<��a<.�a<E�a<�a<Мa<p�a<̛a<<�a<��a<ҙa<�a<��a<�a<��a<��a<��a<ӗa<%�a<��a<=�a<ՙa<m�a<�a<m�a<��a<�a<�a<ܛa<��a<A�a<Κa<V�a<��a<��a<<�a<�a<�a<�a<��a<�a<-�a<C�a<?�a<7�a<�a<p�a<�a<:�a<m�a<��a<��a<��a<ƒa<��a<]�a<ΐa<l�a<U�a<R�a<e�a<��a<��a<T�a<��a<��a<��a<ґa<��a<l�a<ːa<-�a<s�a<��a<��a<"�a<;�a<��a<�a<��a<U�a<҉a<��a<Y�a< �a<��a<&�a<h�a<|�a<��a<p�a<P�a<�a<̀a<�a<i~a<u}a<�|a<�{a<Z{a<{a<�za<�za<'{a<S{a<�{a<�{a<�{a<|a<�{a<�{a<�{a< {a<|za<�ya<Iya<�xa<<xa<�wa<_wa<wa<�va<wa<�va<wa<1wa<2wa<0wa<wa<�va<Wva<�ua<ua<xta<�sa<�ra<@ra<�qa<<qa<�pa<�pa<�pa<Wqa<�qa<qra<<sa<ta<�  �  �ta<�ua<Dva<�va<|wa<�wa<'xa<<xa<sxa<mxa<�xa<}xa<�xa<�xa<"ya<�ya<�ya<�za<7{a<�{a<n|a<�|a<e}a<�}a<�}a<�}a<~a<�}a<�}a<k}a<}a< }a<�|a<
}a<o}a<�}a<�~a<�a<̀a<�a<Y�a<��a<�a<��a<��a<��a<��a<U�a<�a<��a<�a<q�a<ލa<*�a<��a<4�a<ŏa<��a<�a<�a<��a<g�a<%�a<��a<$�a<w�a<��a<��a<��a<A�a<ϔa<��a<��a<Ɠa<u�a<\�a<w�a<˓a<.�a<ݔa<��a<s�a<��a<N�a<d�a<6�a<��a<e�a<��a<��a<
�a<#�a<��a<�a<ʛa<��a<��a<��a<ϛa<��a<�a<��a<��a<�a<�a<O�a<7�a<�a<̜a<P�a<�a<��a<H�a<v�a<��a<)�a<��a<B�a<�a< �a<J�a<Ǘa<9�a<֘a<��a<&�a<��a<V�a<��a<��a<��a<��a<��a<��a<�a<Ԛa<T�a<�a<ؙa<��a<��a<_�a<g�a<��a<{�a<��a<b�a<E�a<�a<��a<ޗa<;�a<k�a<?�a<b�a<C�a<f�a<��a<ʐa<U�a<�a<ˏa<Ϗa<�a<;�a<��a<�a<h�a<ӑa<ˑa<�a<��a<[�a<��a<^�a<��a<��a<B�a<i�a<ڌa<'�a<��a</�a<��a<X�a<��a<��a<9�a<��a<�a<\�a<��a<v�a<��a<,�a<ʁa<��a<%a<~a<�|a<|a<S{a<�za<�za<|za<�za<�za<{a<E{a<�{a<�{a<�{a<|a<�{a<�{a<#{a<�za<*za<�ya<ya<�xa<?xa<�wa<�wa<ywa<Uwa<rwa<awa<swa<Uwa<Qwa<wa<�va<Sva<�ua<0ua<5ta<usa<�ra<�qa<Mqa<�pa<|pa<Npa<�pa<�pa<nqa<	ra<�ra<�sa<�  �  uta<Lua<va<�va<�wa<�wa<Mxa<xxa<�xa<�xa<�xa<�xa<�xa<ya<Xya<�ya<:za<�za<e{a<|a<�|a<}a<�}a<�}a<~a<�}a<�}a<�}a<q}a<8}a<�|a<�|a<�|a<�|a<:}a<�}a<t~a<Xa<��a<��a<%�a<��a<߅a<0�a<r�a<��a<��a<y�a<9�a<ǌa<C�a<��a<�a<j�a<�a<d�a<��a<��a<W�a<(�a<ےa<��a<X�a<�a<M�a<��a<��a<��a<W�a<�a<��a<K�a<Гa<��a<4�a<.�a<K�a<��a<��a<��a<q�a<N�a<L�a<8�a<�a<�a<��a<j�a<֛a< �a<F�a<V�a<<�a<�a<�a<�a<�a<؛a<��a</�a<Z�a<��a<�a<7�a<\�a<x�a<_�a<-�a<a<'�a<��a<ךa<�a<J�a<�a<�a<R�a<�a<זa<�a<�a<��a<�a<��a<e�a<	�a<��a<&�a<��a<�a<�a< �a<�a<��a<W�a<�a<��a<K�a<�a<řa<��a<��a<��a<��a<��a<��a<��a<i�a<�a<��a<͗a<��a<�a<*�a</�a<�a<.�a<N�a<��a< �a<a<��a<��a<ҏa<�a<��a<�a<8�a<��a<��a<�a<őa<�a<$�a<��a<�a<&�a<x�a<��a<�a<X�a<ȋa<^�a<ފa<��a<#�a<ԉa<m�a<�a<>�a<|�a<��a<g�a<8�a<�a<��a<\�a<�~a<�}a<�|a<�{a<'{a<�za<Vza<:za<^za<�za<�za<.{a<u{a<�{a<�{a<|a<�{a<�{a<_{a<�za<gza<�ya<Rya<�xa<lxa<xa<�wa<�wa<�wa<�wa<�wa<�wa<�wa<{wa<3wa<�va<Iva<�ua<�ta<ta<Gsa<nra<�qa<	qa<~pa<>pa<$pa<Ipa<�pa<*qa<�qa<�ra<�sa<�  �  }ta<Kua<Lva<�va<pwa<�wa<7xa<txa<�xa<�xa<�xa<�xa<ya<4ya<�ya<�ya<_za<�za<�{a<|a<�|a<}a<w}a<�}a<�}a<~a<~a<�}a<x}a<}a<�|a<�|a<�|a<�|a<�|a<}}a<M~a<?a<e�a<��a<��a<~�a<�a<;�a<��a<��a<��a<�a<#�a<��a<P�a<��a<2�a<��a<��a<��a<C�a<��a<��a<I�a<��a<��a<=�a<Ҕa<T�a<��a<��a<��a<j�a<�a<��a<�a<˓a<g�a<�a<�a<�a<T�a<�a<v�a<X�a<G�a<�a<@�a<)�a<�a<��a<H�a<ɛa<�a<4�a<<�a<K�a<<�a<+�a<�a<�a<'�a<#�a<A�a<��a<˜a<�a<7�a<W�a<c�a<_�a<�a<Ϝa<c�a<��a<�a<��a<=�a<y�a<ėa<;�a<Ӗa<��a<��a<��a<d�a<��a<��a<?�a<�a<��a<^�a<��a<�a<�a<
�a<�a<��a<l�a<�a<ƚa<d�a<�a<�a<Ùa<ęa<ҙa<әa<șa<��a<��a<W�a<�a<v�a<��a<0�a<$�a<1�a<��a<�a<�a<,�a<�a<��a<��a<n�a<w�a<��a<�a<Z�a<ڐa<K�a<��a<�a<ԑa<��a<��a<�a<}�a<��a<=�a<��a<ލa<�a<��a<�a<f�a<�a<��a<=�a<�a<R�a<҈a<D�a<j�a<|�a<��a<L�a<	�a<��a<.�a<�~a<�}a<�|a<�{a<�za<kza<;za<za<Dza<�za<�za<6{a<�{a<�{a<|a<�{a<�{a<�{a<N{a<�za<vza<�ya<{ya<�xa<txa<Uxa<�wa<�wa<�wa<�wa<�wa<�wa<�wa<ewa<3wa<�va<Vva<�ua<�ta< ta<*sa<bra<�qa<�pa<gpa<pa<�oa<pa<�pa<qa<�qa<�ra<rsa<�  �  uta<Lua<va<�va<�wa<�wa<Mxa<xxa<�xa<�xa<�xa<�xa<�xa<ya<Xya<�ya<:za<�za<e{a<|a<�|a<}a<�}a<�}a<~a<�}a<�}a<�}a<q}a<8}a<�|a<�|a<�|a<�|a<:}a<�}a<t~a<Xa<��a<��a<%�a<��a<߅a<0�a<r�a<��a<��a<y�a<9�a<ǌa<C�a<��a<�a<j�a<�a<d�a<��a<��a<W�a<(�a<ےa<��a<X�a<�a<M�a<��a<��a<��a<W�a<�a<��a<K�a<Гa<��a<4�a<.�a<K�a<��a<��a<��a<q�a<N�a<L�a<8�a<�a<�a<��a<j�a<֛a< �a<F�a<V�a<<�a<�a<�a<�a<�a<؛a<��a</�a<Z�a<��a<�a<7�a<\�a<x�a<_�a<-�a<a<'�a<��a<ךa<�a<J�a<�a<�a<R�a<�a<זa<�a<�a<��a<�a<��a<e�a<	�a<��a<&�a<��a<�a<�a< �a<�a<��a<W�a<�a<��a<K�a<�a<řa<��a<��a<��a<��a<��a<��a<��a<i�a<�a<��a<͗a<��a<�a<*�a</�a<�a<.�a<N�a<��a< �a<a<��a<��a<ҏa<�a<��a<�a<8�a<��a<��a<�a<őa<�a<$�a<��a<�a<&�a<x�a<��a<�a<X�a<ȋa<^�a<ފa<��a<#�a<ԉa<m�a<�a<>�a<|�a<��a<g�a<8�a<�a<��a<\�a<�~a<�}a<�|a<�{a<'{a<�za<Vza<:za<^za<�za<�za<.{a<u{a<�{a<�{a<|a<�{a<�{a<_{a<�za<gza<�ya<Rya<�xa<lxa<xa<�wa<�wa<�wa<�wa<�wa<�wa<�wa<{wa<3wa<�va<Iva<�ua<�ta<ta<Gsa<nra<�qa<	qa<~pa<>pa<$pa<Ipa<�pa<*qa<�qa<�ra<�sa<�  �  �ta<�ua<Dva<�va<|wa<�wa<'xa<<xa<sxa<mxa<�xa<}xa<�xa<�xa<"ya<�ya<�ya<�za<7{a<�{a<n|a<�|a<e}a<�}a<�}a<�}a<~a<�}a<�}a<k}a<}a< }a<�|a<
}a<o}a<�}a<�~a<�a<̀a<�a<Y�a<��a<�a<��a<��a<��a<��a<U�a<�a<��a<�a<q�a<ލa<*�a<��a<4�a<ŏa<��a<�a<�a<��a<g�a<%�a<��a<$�a<w�a<��a<��a<��a<A�a<ϔa<��a<��a<Ɠa<u�a<\�a<w�a<˓a<.�a<ݔa<��a<s�a<��a<N�a<d�a<6�a<��a<e�a<��a<��a<
�a<#�a<��a<�a<ʛa<��a<��a<��a<ϛa<��a<�a<��a<��a<�a<�a<O�a<7�a<�a<̜a<P�a<�a<��a<H�a<v�a<��a<)�a<��a<B�a<�a< �a<J�a<Ǘa<9�a<֘a<��a<&�a<��a<V�a<��a<��a<��a<��a<��a<��a<�a<Ԛa<T�a<�a<ؙa<��a<��a<_�a<g�a<��a<{�a<��a<b�a<E�a<�a<��a<ޗa<;�a<k�a<?�a<b�a<C�a<f�a<��a<ʐa<U�a<�a<ˏa<Ϗa<�a<;�a<��a<�a<h�a<ӑa<ˑa<�a<��a<[�a<��a<^�a<��a<��a<B�a<i�a<ڌa<'�a<��a</�a<��a<X�a<��a<��a<9�a<��a<�a<\�a<��a<v�a<��a<,�a<ʁa<��a<%a<~a<�|a<|a<S{a<�za<�za<|za<�za<�za<{a<E{a<�{a<�{a<�{a<|a<�{a<�{a<#{a<�za<*za<�ya<ya<�xa<?xa<�wa<�wa<ywa<Uwa<rwa<awa<swa<Uwa<Qwa<wa<�va<Sva<�ua<0ua<5ta<usa<�ra<�qa<Mqa<�pa<|pa<Npa<�pa<�pa<nqa<	ra<�ra<�sa<�  �  �ta<�ua<[va<�va<gwa<�wa<	xa<xa<+xa<xa<xa<$xa<<xa<Rxa<�xa<�xa<�ya<!za<�za<v{a<%|a<�|a<X}a<�}a<�}a< ~a<~a<�}a<�}a<�}a<�}a<`}a<f}a<�}a<�}a<f~a<3a<�a<�a<Z�a<��a<��a<@�a<j�a<��a<��a<��a<f�a<�a<`�a<ǌa<(�a<X�a<�a<"�a<��a<F�a<�a<ΐa<l�a<i�a<,�a<�a<��a<6�a<��a<��a<ȕa<��a<e�a< �a<��a<q�a<�a<��a<�a<��a<C�a<a<U�a<�a<�a<��a<��a<o�a<*�a<�a<E�a<��a<��a<�a<ܛa<��a<��a<Q�a<Q�a<�a<1�a<9�a<s�a<ʛa<�a<f�a<a<��a<.�a<E�a<�a<Мa<p�a<̛a<<�a<��a<ҙa<�a<��a<�a<��a<��a<��a<ӗa<%�a<��a<=�a<ՙa<m�a<�a<m�a<��a<�a<�a<ܛa<��a<A�a<Κa<V�a<��a<��a<<�a<�a<�a<�a<��a<�a<-�a<C�a<?�a<7�a<�a<p�a<�a<:�a<m�a<��a<��a<��a<ƒa<��a<]�a<ΐa<l�a<U�a<R�a<e�a<��a<��a<T�a<��a<��a<��a<ґa<��a<l�a<ːa<-�a<s�a<��a<��a<"�a<;�a<��a<�a<��a<U�a<҉a<��a<Y�a< �a<��a<&�a<h�a<|�a<��a<p�a<P�a<�a<̀a<�a<i~a<u}a<�|a<�{a<Z{a<{a<�za<�za<'{a<S{a<�{a<�{a<�{a<|a<�{a<�{a<�{a< {a<|za<�ya<Iya<�xa<<xa<�wa<_wa<wa<�va<wa<�va<wa<1wa<2wa<0wa<wa<�va<Wva<�ua<ua<xta<�sa<�ra<@ra<�qa<<qa<�pa<�pa<�pa<Wqa<�qa<qra<<sa<ta<�  �  <ua<�ua<�va<�va<Twa<�wa<�wa<�wa<�wa<�wa<�wa<�wa<�wa<�wa<*xa<lxa<-ya<�ya<^za<{a<�{a<v|a<�|a<�}a<�}a<<~a<=~a</~a<F~a<�}a<�}a<�}a<�}a<~a<i~a<a<�a<��a<��a<�a< �a<S�a<��a<��a<ވa<��a<t�a<�a<��a<�a<E�a<ƌa<Όa<d�a<��a<(�a<a<Z�a<V�a<ܐa<��a<��a<��a<=�a<ܔa<`�a<��a<�a<��a<��a<��a<�a<��a<��a<��a<k�a<��a<Ȕa<=�a<ԕa<�a<d�a<�a<�a<��a<U�a<�a<=�a<��a<��a<��a<~�a<R�a<$�a<��a<ښa<��a<��a<��a<��a<=�a<��a<�a<G�a<��a<՜a<�a<��a<Ԝa<��a<��a<��a<ܚa<9�a<��a<�a<��a<8�a<+�a<�a<`�a<��a<�a<��a<%�a<Кa<�a<��a<ța<Лa<Лa<��a<J�a<˚a<~�a<ۙa<i�a<#�a<��a<��a<W�a<��a<_�a<��a<Әa<ߘa<��a<٘a<ǘa<d�a<�a<j�a<��a<��a<�a<,�a<@�a<~�a<ۑa<O�a<�a<Ґa<ڐa<�a<9�a<[�a<��a<�a<�a<#�a<ӑa<��a<�a<v�a<ۏa<��a<O�a<2�a<��a<��a<�a<��a<�a<݉a<B�a<F�a<܈a<��a<=�a<̇a<E�a<y�a<Ѕa<��a<��a<��a<.�a<'�a<�~a<�}a<}a<h|a<�{a<�{a<t{a<l{a<�{a<�{a<|a<|a<|a<;|a<�{a<�{a<2{a<�za<za<~ya<�xa<xa<�wa<wa<�va<�va<�va<tva<qva<�va<�va<�va<�va<�va<�va<[va<va<Kua<�ta<	ta<]sa<�ra<*ra<�qa<qqa<wqa<~qa<�qa<Ora<�ra<�sa<Xta<�  �  dua< va<�va<wa<_wa<ywa<�wa<�wa<@wa<.wa<#wa<�va<�va< wa<qwa<�wa<Yxa<ya<�ya<|za<V{a<+|a<�|a<c}a<�}a<,~a<|~a<�~a<j~a<�~a<k~a<x~a<�~a<�~a<'a<�a<_�a<E�a<H�a<T�a<��a<��a<��a<��a<Јa<��a<f�a<�a<Y�a<��a<ŋa<)�a<]�a<��a< �a<q�a<
�a<��a<z�a<h�a<g�a<)�a<:�a<�a<��a<E�a<��a<ޕa<�a<�a<̕a<��a<`�a<B�a<"�a<�a<B�a<��a<�a<~�a<%�a<͗a<��a<:�a<��a<��a<��a<U�a<h�a<s�a<]�a<�a<��a<��a<;�a<�a<�a<�a<��a<C�a<��a<�a<v�a<̛a<\�a<��a<ܜa<��a<ߜa<��a<^�a<��a<O�a<Ěa<,�a<��a<E�a<��a<Ϙa<֘a<�a<S�a<��a<)�a<��a<��a<v�a<��a<͛a<ܛa<��a<_�a<��a<V�a<ޙa<h�a<ɘa<a�a<
�a<ޗa<��a<��a<ۗa<)�a<2�a<t�a<��a<��a<��a<z�a<�a<��a<��a<"�a<z�a<��a<ޓa<+�a<��a<�a<��a<��a<}�a<��a<��a<�a<�a<�a<P�a<�a<�a<��a<�a<D�a<��a<q�a<��a<��a<ˋa<�a<e�a<ىa<f�a<�a<ψa<��a<V�a<N�a<�a<��a<*�a<��a<��a< �a<׃a<ǂa<��a<��a<�a<�~a<�}a<}a<�|a<L|a<|a<|a<|a<7|a<1|a<T|a<j|a<&|a<�{a<�{a<{a<wza<�ya<�xa<[xa<�wa<�va<rva<va<�ua<�ua<�ua<va<"va<;va<�va<�va<�va<�va<eva<va<�ua<�ta<|ta<�sa<Msa<�ra<pra<,ra<ra<;ra<�ra<�ra<�sa<(ta<�ta<�  �  �ua<qva<�va<"wa<Lwa<Ewa<Swa<wa<wa<�va<rva<Sva<Kva<ova<�va<(wa<�wa<gxa<#ya<za<{a<�{a<�|a<0}a<�}a<C~a<�~a<�~a<�~a<a<�~a<a<1a<�a<�a<c�a</�a<�a<�a<܃a<�a<7�a<�a<?�a<�a<ىa<8�a<Ȋa<�a<K�a<��a<s�a<ŋa<�a<Y�a<��a<H�a<�a<Ύa<ԏa<��a<��a<Ӓa<��a<��a<�a<ؕa<��a<U�a<A�a<Q�a<6�a<�a<�a<Õa<�a<��a<:�a<��a<�a<Ηa<O�a<9�a<��a<N�a<Κa<	�a<i�a<9�a<T�a<�a<Ța<R�a<ߙa<��a<K�a<E�a<#�a<M�a<��a<�a<h�a<њa<��a<�a<l�a<��a<�a<�a<��a<��a<&�a<�a<6�a<��a<W�a<�a<��a<��a<��a<��a<��a<G�a<��a<5�a<b�a<ƛa<ʛa<�a<ɛa<o�a<%�a<��a<�a<C�a<��a<*�a<��a<X�a<
�a<�a<�a<@�a<m�a<��a<+�a<<�a<��a<i�a<��a<$�a<ȗa<K�a<��a<�a<�a<��a<Ǔa<H�a<Œa<j�a<Q�a<�a<7�a<0�a<l�a<��a<t�a<��a<)�a<�a<W�a<ϐa<�a<�a<6�a<��a<*�a<#�a<s�a<��a<�a<��a<U�a<:�a<�a<�a<�a<��a<��a<��a<��a<ԅa<6�a<,�a<L�a<F�a<�a<9�a<:a<�~a<�}a<P}a<}a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<:|a<|a<T{a<�za<za<hya<~xa<�wa<�va<6va<�ua<Qua<$ua<ua<ua<Xua<~ua<va<&va<ova<�va<�va<�va<$va<�ua<aua<ua<Zta<�sa<zsa<sa<�ra<�ra<�ra<2sa<�sa<ta<�ta<gua<�  �  ?va<�va<�va<0wa<-wa<.wa< wa<�va<wva<va<�ua<�ua<�ua<�ua<�ua<]va< wa<�wa<�xa<�ya<{za<U{a<f|a<}a<�}a<g~a<�~a<a<Ua<Pa<�a<�a<�a<3�a<��a<,�a<сa<��a<��a<��a<n�a<��a<��a<\�a<�a<��a<"�a<��a<��a<Ŋa<�a<��a<�a<I�a<��a<�a<��a<I�a</�a<+�a<'�a<Q�a<O�a<U�a<d�a<��a<��a<#�a<p�a<��a<��a<��a<��a<�a<r�a<��a<��a<��a<_�a<��a<g�a< �a<o�a<+�a<��a<�a<5�a<F�a<$�a<�a<��a<9�a<יa<S�a<��a<��a<u�a<p�a<��a<�a<H�a<Ǚa<V�a<�a<v�a<�a<��a<ǜa<�a<�a<לa<��a<'�a<��a<t�a<�a<��a<k�a<U�a<J�a<h�a<��a<��a<1�a<r�a<ԛa<��a< �a<��a<��a<X�a<Қa<�a<��a<̘a<�a<��a< �a<��a<Y�a<H�a<d�a<��a<ߖa<G�a<��a<֗a<E�a<U�a<]�a<G�a<�a<��a<�a<G�a<��a<&�a<h�a<�a<z�a<3�a<�a<Ӓa<Вa<�a<ɒa<�a<�a<��a<W�a<�a<A�a<��a<��a<��a<��a<y�a<��a<��a<��a<��a<f�a<�a<��a<��a<o�a<}�a<d�a<U�a<T�a<�a<��a< �a<Q�a<��a<��a<��a<ҁa<΀a<�a<1a<�~a<~a<�}a<^}a<T}a<?}a<}a<"}a<�|a<�|a<f|a<�{a<?{a<�za<�ya<�xa<xa<wa<Lva<�ua< ua<�ta<ita<fta<�ta<�ta<ua<qua<�ua<va<gva<qva<�va<Zva<&va<�ua<Tua<�ta<�ta<ta<�sa<�sa<�sa<�sa<�sa<>ta<�ta</ua<�ua<�  �  �va<�va<wa<"wa</wa<wa<�va<|va<�ua<�ua<Dua<ua<�ta<�ta<Iua<�ua<\va<wa<xa<ya<za<1{a<|a<}a<�}a<e~a<�~a<Da<�a<�a<1�a<1�a<��a<�a<G�a<�a<l�a<t�a< �a<'�a<�a<��a<͇a<��a<;�a<��a<:�a<D�a<k�a<��a<f�a<��a<s�a<��a<܊a<C�a<݋a<��a<��a<��a<a<Đa<�a<�a<�a<�a<��a<C�a<��a<�a<�a<�a<6�a<�a<N�a<(�a<r�a<��a<�a<��a<ؘa<��a<�a<��a<ɚa<�a<>�a<2�a<.�a<��a<f�a<ؙa<H�a<ݘa<O�a<�a<a<ʗa<ԗa<.�a<��a<-�a<�a<z�a<R�a<Ûa<]�a<Ӝa<�a<�a<��a<�a<��a<[�a<�a<|�a<q�a<�a<�a<�a<-�a</�a<r�a<қa<�a<$�a<�a<-�a<�a<��a<6�a<z�a<�a<�a<O�a<��a<ږa<V�a<ڕa<��a<��a<��a<�a<Z�a<��a<+�a<��a<�a<Q�a<N�a<E�a<�a<��a<e�a<a<a�a<��a<'�a<��a<-�a<�a<��a<��a<I�a<{�a<_�a<M�a<&�a<Ւa<��a<ܑa<Y�a<K�a<V�a<b�a<�a<�a<؊a<��a<��a<7�a<��a<C�a<�a<�a<
�a<��a<%�a<�a<�a<��a<|�a< �a<}�a<̄a<�a<"�a<b�a<B�a<ŀa<�a<Ma<�~a<_~a<0~a<�}a<�}a<�}a<z}a<#}a<�|a<o|a<�{a<I{a<Hza<�ya<yxa<twa<�va<�ua<�ta<Lta<�sa<�sa<�sa<�sa<ta<�ta<�ta<�ua<�ua<0va<}va<tva<�va<Hva<va<�ua<ua<ua<�ta<�ta<>ta<Zta<Nta<�ta<�ta<Aua<�ua<va<�  �  �va<#wa<Owa<2wa<wa<�va<wva<va<�ua<5ua<�ta<�ta<kta<qta<�ta<(ua<�ua<�va<�wa<�xa<�ya<�za<�{a<�|a<�}a<�~a<3a<�a<�a<I�a<��a<��a<�a<^�a<ρa<n�a<��a<�a<��a<��a<p�a<L�a<�a<ވa<b�a<��a<�a<�a<(�a<1�a<�a<
�a<��a<#�a<d�a<��a<J�a<!�a<�a<�a<;�a<d�a<��a<ɒa<֓a<�a<��a<g�a<��a<*�a<j�a<��a<��a<��a<×a<��a<��a<2�a<��a<�a<_�a<��a<n�a<Қa< �a<j�a<[�a<1�a<�a<{�a<�a<��a<�a<U�a<Ηa<{�a<F�a<)�a<S�a<��a<�a<��a<s�a<(�a<�a<��a<+�a<��a<��a<I�a<V�a<,�a<��a<��a<b�a<�a<�a<��a<��a<y�a<��a<Ûa<�a<#�a<W�a<i�a<y�a<a�a<��a<��a<�a<J�a<��a<��a<�a<�a<W�a<͕a<[�a<�a<�a<0�a<l�a<וa<T�a<ݖa<W�a<��a<&�a<N�a<_�a<_�a<�a<��a<@�a<��a<�a<��a<�a<��a<t�a< �a<!�a<��a<�a<˓a<��a<h�a</�a<��a<�a<5�a< �a<�a<��a<��a<��a<]�a<c�a<~�a<��a<�a<ˆa<��a<k�a<��a<��a<��a<Ɇa<Ɔa<ӆa<��a<C�a<؅a<�a<e�a<��a<΂a<ԁa<:�a<Y�a<�a<Ha<�~a<�~a<L~a<;~a<~a<�}a<{}a<-}a<�|a<�{a<{a<za<*ya<$xa<wa<va< ua<gta<�sa<Xsa<*sa<2sa<Rsa<�sa<ta<�ta<&ua<�ua<�ua<eva<�va<�va<�va<fva<)va<�ua<�ua<:ua<ua<�ta<�ta<�ta<,ua<iua<�ua<!va<�va<�  �  �va<?wa<@wa<Kwa<wa<�va<�va<�ua<cua<�ta<`ta<ta<�sa<�sa< ta<�ta<Iua<=va<!wa<Gxa<wya<�za<�{a<�|a<�}a<�~a<#a<�a<�a<��a<рa<5�a<m�a<�a<b�a<ނa<��a<3�a<�a<�a<��a<��a<3�a<؈a<S�a<̉a<�a<+�a<�a<Չa<Ӊa<��a<��a<��a<Ήa<D�a<Њa<��a<��a<��a<a<,�a<U�a<��a<�a<��a<��a<Y�a<�a<R�a<��a<ŗa<��a<�a<�a<U�a<o�a<��a<�a<^�a<�a<D�a<��a<��a<H�a<X�a<Y�a<<�a<ښa<��a<יa<8�a<��a<�a<|�a<��a<��a<��a<ۖa<�a<��a<P�a<��a<�a<��a<��a<(�a<��a<�a<<�a<k�a<O�a<D�a<��a<Ӝa<}�a<F�a<5�a<�a<�a<�a<�a<d�a<r�a<��a<��a<��a<S�a<�a<��a<��a<W�a<C�a<x�a<w�a<��a<��a<A�a<��a<��a<��a<��a<�a<j�a<��a<��a<�a<Ǘa< �a<O�a<g�a<O�a<5�a<ԗa<��a<�a<��a<�a<��a<H�a<�a<��a<l�a<_�a<A�a<�a<�a<��a<)�a<��a<��a<�a<2�a<�a<��a<�a<�a<�a<�a<�a<7�a<��a<3�a<�a<�a<
�a<Y�a<i�a<��a<ކa<��a<��a<6�a<Ʌa<=�a<��a<Ճa< �a<Z�a<~�a<��a<K�a<�a<ra<�~a<�~a<�~a<E~a<�}a<�}a<}a<�|a<�{a<�za<*za<�xa<�wa<�va<�ua<�ta<�sa<Ksa<�ra<�ra<�ra<�ra<@sa<�sa<Yta<�ta<�ua<�ua<Hva<�va<�va<�va<�va<qva<#va<�ua<�ua<pua<mua<Qua<|ua<�ua<�ua<3va<pva<�va<�  �  4wa<cwa<fwa<Zwa< wa<�va<-va<�ua<0ua<�ta<)ta<�sa<�sa<�sa<�sa<nta<ua<�ua<�va<xa<Mya<sza<�{a<�|a<�}a<�~a<Ka<�a<Y�a<��a<�a<f�a<��a<!�a<��a<�a<˃a<|�a<N�a<�a<�a<Ça<q�a<�a<z�a<щa<։a<�a<Ӊa<��a<��a<n�a<f�a<a�a<��a<�a<��a<\�a<C�a<r�a<��a<��a<8�a<o�a<��a<��a<��a<|�a<�a<��a<ݗa<�a<�a<B�a<P�a<��a<��a<�a<N�a<��a<�a<u�a<�a<8�a<v�a<|�a<p�a<<�a<��a<?�a<��a<�a<f�a<��a<8�a<��a<��a<|�a<��a<�a<p�a<�a<֘a<��a<��a<B�a<�a<��a<"�a<g�a<��a<��a<s�a<:�a<�a<��a<��a<`�a<;�a<A�a<N�a<[�a<��a<��a<Μa<ɜa<��a<y�a<$�a<}�a<a<��a<(�a<E�a<L�a<n�a<��a<�a<��a<c�a<X�a<s�a<єa<7�a<ϕa<j�a<�a<q�a<ۗa<G�a<y�a<w�a<`�a<�a<��a<<�a<˖a<A�a<�a<w�a<�a<�a<��a<��a<j�a<K�a< �a<ʓa<W�a<��a<�a<��a<�a<��a<��a<H�a<��a<ˉa<��a<��a<�a<p�a<�a<ʅa<مa<�a<!�a<L�a<o�a<��a<��a<��a<X�a<�a<v�a<ׄa<�a<D�a<��a<ǁa<+�a<��a<�a<�a<=a<a<�~a<~a</~a<�}a<?}a<�|a<�{a<�za<�ya<�xa<�wa<�va<uua<�ta<�sa<sa<�ra<|ra<mra<�ra<sa<�sa<&ta<�ta<Dua<�ua<8va<�va<�va<�va<�va<�va<^va<"va<�ua<�ua<�ua<�ua<�ua<�ua<va<cva<�va< wa<�  �  �xa<�xa<�xa<�xa<�xa<fxa<xa<�wa<Iwa<wa<�va<�va<�va<�va<�va<-wa<�wa<�xa<vya<eza<X{a<�|a<f}a<O~a<a<�a<��a< �a<��a<��a<��a<��a<7�a<��a<�a<τa<4�a<��a<��a<n�a<(�a<ۈa<��a<�a<��a<�a<(�a<^�a<x�a<��a<p�a<��a<��a<ɋa<�a<s�a<�a<��a<��a<|�a<��a<��a<Ւa<�a<�a<ƕa<��a<U�a<ؗa<J�a<��a<ܘa<�a<%�a<n�a<�a<�a<�a<S�a<��a< �a<��a<��a<�a<=�a<Z�a<W�a<�a<�a<��a<G�a<��a<-�a<əa<M�a< �a<Θa<�a<�a<H�a<��a<#�a<њa<Y�a<1�a<��a<D�a<��a<�a<T�a<i�a<m�a<U�a<@�a<�a<ȝa<��a<��a<��a<l�a<|�a<}�a<��a<��a<��a<��a<��a<o�a<�a<��a<�a<s�a<ޚa<�a<G�a<��a<�a<v�a<��a<�a<��a<�a<��a<S�a<��a<�a<��a<ܘa< �a<7�a<h�a<e�a<1�a<��a<��a<R�a<×a<p�a<��a<��a<~�a<�a<ߕa<��a<w�a<;�a<�a<��a<+�a<��a<�a<�a<<�a<A�a<;�a<�a<�a<�a<�a<&�a<r�a<�a<v�a<I�a<�a<�a<�a<"�a</�a<�a<�a<��a<��a<�a<��a<�a<M�a<��a<ڃa<N�a<��a<1�a<��a<�a<Ѐa<^�a<2�a<�a<ua<a<�~a<�}a<)}a<y|a<�{a<�za<�ya<�xa<�wa<wa<�va<�ua<�ua<Cua<Iua<Wua<�ua<�ua<Eva<�va<5wa<�wa<�wa<xa<;xa<7xa<(xa<xa<�wa<�wa<kwa<cwa<<wa<{wa<Owa<}wa<�wa<�wa<7xa<]xa<�  �  �xa<�xa<�xa<�xa<�xa<nxa<xa<�wa<gwa<wa<�va<�va<�va<�va<�va<Swa<�wa<�xa<ya<sza<l{a<_|a<i}a<_~a<.a<�a<��a<�a<��a<�a<`�a<��a<,�a<��a<��a<��a<2�a<�a<��a<[�a<�a<؈a<}�a<�a<��a<��a<1�a<d�a<f�a<z�a<��a<��a<��a<ڋa< �a<z�a<�a<Ӎa<��a<��a<��a<��a<˒a<Փa<�a<ҕa<��a<F�a<ٗa<B�a<��a<ؘa<�a<1�a<e�a<��a<��a<�a<Q�a<��a<�a<b�a<��a<�a<5�a<R�a<V�a<4�a<��a<��a< �a<��a<@�a<șa<`�a<(�a<��a<�a<�a<[�a<��a<9�a<Қa<}�a<�a<��a<H�a<��a<�a<;�a<j�a<c�a<V�a<%�a<��a<ҝa<��a<y�a<]�a<]�a<��a<��a<��a<��a<��a<��a<��a<V�a<�a<��a<!�a<k�a<��a<�a<J�a<��a<��a<��a<�a<ݖa<Ζa<�a<�a<\�a<��a<�a<v�a<��a<0�a<V�a<l�a<X�a<.�a<��a<��a<1�a<×a<e�a<��a<��a<7�a<��a<ڕa<��a<d�a<-�a<�a<��a<.�a<��a<��a<"�a<C�a</�a<+�a<!�a< �a<��a<�a<>�a<y�a<�a<��a<T�a<�a<�a<�a<�a<�a<�a<��a<Շa<t�a<�a<��a<�a<I�a<��a<�a<F�a<��a<��a<s�a<�a<Àa<c�a<�a<�a<qa<a<�~a<�}a<M}a<�|a<�{a<�za<�ya<�xa<�wa<*wa<�va<�ua<�ua<Wua<\ua<lua<�ua<�ua<iva<�va<)wa<�wa<�wa<xa<"xa<8xa<xa<xa<�wa<�wa<uwa<gwa<1wa<(wa<@wa<�wa<�wa<�wa<xa<bxa<�  �  fxa<�xa<�xa<�xa<�xa<uxa<1xa<�wa<�wa<3wa<wa<�va<�va<�va<wa<�wa<xa<�xa<�ya<�za<�{a<r|a<�}a<Z~a<*a<�a<��a<�a<p�a<�a<*�a<��a<�a<Z�a<ڃa<O�a<	�a<��a<r�a<.�a<�a<��a<X�a<�a<p�a<�a<'�a<��a<��a<��a<ċa<��a<�a<��a<H�a<��a<O�a<�a<Ŏa<׏a<ːa<��a<��a<��a<�a<ƕa<��a<0�a<їa<�a<l�a<��a<Ҙa<�a<�a<Z�a<z�a<̙a<�a<h�a<�a<-�a<��a<֛a<�a<F�a<C�a<1�a<�a<a<8�a<�a<n�a<��a<��a<@�a<:�a<#�a<O�a<�a<ޙa<~�a<��a<��a< �a<˜a<W�a<��a<�a<&�a<b�a<8�a<7�a<��a<؝a<��a<g�a<U�a<#�a<8�a<1�a<B�a<l�a<k�a<��a<�a<��a<?�a<�a<��a<'�a<��a<Śa<C�a<n�a<ݘa<%�a<��a<b�a<�a<�a<�a<B�a<��a<�a<S�a<��a<�a<+�a<R�a<]�a<I�a< �a<Ƙa<��a<��a<��a<�a<��a<g�a<��a<֕a<��a<l�a<6�a< �a<Ɣa<p�a<'�a<}�a<�a<�a<^�a<T�a<J�a<Z�a<-�a<>�a<-�a<f�a<��a<0�a<Ȉa<k�a<c�a<>�a<T�a<A�a<4�a<>�a<�a<هa<^�a<�a<b�a<Ņa<�a<b�a<��a<�a<l�a<Áa<Q�a<�a<x�a<@�a<�a<�a<@a<�~a<}~a<�}a<J}a<�|a<�{a<�za<�ya<ya<2xa<fwa<�va<>va<�ua<�ua<�ua<�ua<�ua<"va<�va<�va<Kwa<�wa<�wa<xa<xa<0xa<�wa<�wa<�wa<ywa<>wa<wa<wa<�va<wa<2wa<gwa<�wa<�wa<Fxa<�  �  Ixa<�xa<�xa<�xa<�xa<xa<Jxa<xa<�wa<hwa<Cwa<wa<wa<,wa<lwa<�wa<sxa<!ya<�ya<�za<�{a<�|a<�}a<i~a<4a<�a<`�a<�a<L�a<��a<��a<L�a<��a<��a<�a<�a<��a<]�a<#�a<�a<��a<��a<<�a<݉a<v�a<�a<:�a<��a<��a<ҋa<ыa<�a<�a<T�a<��a<�a<��a<R�a<.�a<�a<
�a<	�a<#�a<"�a<�a<ڕa<��a<5�a<��a<�a<W�a<m�a<��a<��a<Ҙa<��a<9�a<{�a<��a<(�a<��a<��a<\�a<��a<�a<�a<E�a<:�a<�a<ța<x�a<�a<��a<?�a<�a<��a<x�a<q�a<��a<�a<9�a<��a<1�a<Ǜa<m�a<�a<`�a<��a<�a<"�a<-�a<�a<	�a<��a<��a<T�a<�a<��a<�a<֜a<ݜa<�a<$�a<6�a<a�a<b�a<^�a<5�a<�a<��a<1�a<��a<�a<[�a<��a<�a<z�a<	�a<��a<h�a<U�a<h�a<��a<՗a<�a<t�a<Әa<�a<:�a<\�a<^�a<(�a<��a<��a<@�a<ɗa<S�a<ޖa<b�a<�a<ƕa<w�a<C�a<�a<��a<Ɣa<��a<T�a<�a<��a<�a<,�a<e�a<z�a<��a<g�a<l�a<y�a<��a<a<�a<�a<�a<Ԉa<��a<~�a<g�a<o�a<`�a<C�a<�a<Їa<c�a<نa<J�a<��a<߄a<$�a<g�a<��a<	�a<��a< �a<��a<8�a<�a<�a<ga<$a<�~a<W~a<�}a<S}a<�|a<�{a<	{a<za<7ya<txa<�wa<wa<|va<va<�ua<�ua<�ua<$va<Zva<�va< wa<mwa<�wa<�wa<xa<
xa<�wa<�wa<�wa<cwa<3wa<�va<�va<�va<�va<�va<�va<&wa<qwa<�wa<xa<�  �  "xa<Zxa<�xa<�xa<�xa<�xa<lxa<Pxa<�wa<�wa<�wa<xwa<�wa<�wa<�wa<Axa<�xa<}ya<Wza<1{a<|a<�|a<�}a<�~a</a<�a<P�a<��a<!�a<O�a<��a<�a<J�a<��a<�a<��a<&�a<�a<��a<��a<V�a<C�a<�a<��a<x�a<�a<`�a<��a<�a<�a<%�a<i�a<l�a<Ōa<
�a<��a<�a<��a<��a<`�a<�a<a�a<j�a<V�a<-�a<�a<��a<1�a<��a<՗a<�a<�a<>�a<L�a<{�a<{�a<ǘa< �a<Q�a<љa<%�a<��a<��a<��a<՛a<�a<<�a<2�a<,�a<ߛa<��a<P�a<��a<��a<:�a<*�a<�a<��a<�a<L�a<��a<
�a<��a<�a<��a<�a<��a<ϝa<��a<"�a<	�a<��a<��a<k�a<)�a<�a<��a<u�a<x�a<[�a<��a<��a<��a<�a<�a<;�a<5�a<1�a<��a<��a<U�a<Ǜa<P�a<��a<�a<n�a<ܘa<|�a<�a<�a<��a<�a<�a<5�a<|�a<��a<�a<'�a<c�a<X�a<X�a<�a<јa<w�a<�a<y�a<�a<��a<��a<��a<R�a<�a<�a<��a<��a<i�a<[�a<$�a<ѓa<��a<�a<R�a<��a<��a<ɏa<��a<�a<Ȍa<�a<)�a<��a<��a<}�a<G�a<�a<�a<��a<��a<��a<`�a<0�a<a<`�a<��a<�a<e�a<�a<΃a<�a<\�a<��a<�a<��a<�a<�a<�a<\a<	a<�~a<�~a<?~a<�}a<K}a<�|a<�{a<B{a<hza<�ya<�xa<xa<�wa<�va<�va<Sva<Lva<Tva<vva<�va<�va<awa<�wa<�wa<�wa<xa<	xa<�wa<�wa<^wa<wa<�va<�va<kva<-va<Cva<>va<�va<�va<wa<_wa<�wa<�  �  �wa<,xa<uxa<�xa<�xa<�xa<�xa<�xa<Wxa<(xa<xa<�wa<�wa<%xa<rxa<�xa<Mya<�ya<�za<z{a<\|a<*}a<�}a<�~a<0a<�a<<�a<��a<̀a<�a<C�a<��a<��a<�a<��a<�a<Ńa<h�a<H�a<7�a<�a<��a<ňa<��a<L�a<�a<R�a<ʋa<#�a<O�a<��a<��a<��a<-�a<��a<�a<��a<:�a<�a<�a<Ցa<��a<��a<��a<Y�a<��a<��a<
�a<u�a<��a<��a<ӗa<��a<�a<ܗa<�a<F�a<��a<ۘa<1�a<˙a<B�a<Úa<3�a<��a<��a<#�a<3�a<.�a<"�a<�a<��a<A�a< �a<��a<��a<j�a<z�a<��a<��a<�a<��a<�a<o�a<ޜa<]�a<��a<Ɲa<��a<��a<�a<��a<l�a< �a<Ӝa<j�a<+�a<�a<�a<��a<��a<�a<\�a<��a<ǜa<�a<�a<�a<��a<��a<q�a<�a<��a<��a<c�a<�a<T�a<�a<��a<o�a<J�a<C�a<g�a<��a<Ęa<�a<A�a<p�a<o�a<Y�a<D�a<�a<��a<"�a<��a<�a<��a<�a<��a<�a<Δa<��a<N�a<A�a<?�a<(�a<�a<ݓa<��a<X�a<�a<D�a<��a<�a<��a<�a<3�a<Q�a<j�a<��a<�a<�a<��a<��a<z�a<I�a<�a<��a<шa<��a<$�a<Ƈa<9�a<��a<څa<�a<E�a<q�a<��a<��a<#�a<��a<�a<�a<Aa<)a<�~a<�~a<�~a<g~a<4~a<�}a<K}a<�|a<1|a<w{a<�za<�ya<4ya<�xa<�wa<nwa<"wa<�va<�va<�va<�va<wa<[wa<�wa<�wa<�wa<�wa<xa<�wa<�wa<]wa<wa<�va<tva<va<�ua<�ua<�ua<�ua<�ua<2va<�va<wa<vwa<�  �  {wa<�wa<Axa<�xa<�xa<�xa<�xa<�xa<�xa<xxa<�xa<|xa<�xa<�xa<�xa<oya<�ya<�za<-{a<�{a<�|a<Z}a<~a<�~a<ba<�a<�a<P�a<x�a<��a<��a<�a<>�a<��a<��a<p�a<E�a<�a<�a<��a<��a<��a<��a<r�a<�a<�a<f�a<�a<J�a<��a<�a<�a<��a<��a<(�a<��a<�a<ݏa<��a<|�a<&�a<#�a<��a<��a<~�a<�a<Ŗa<��a<9�a<P�a<q�a<m�a<R�a<~�a<]�a<��a<��a<�a<b�a<��a<`�a<��a<m�a<ޚa<[�a<��a<�a<e�a<7�a<K�a<�a<�a<��a<m�a<Q�a<�a<�a<��a<�a<U�a<��a<�a<?�a<ٜa<�a<��a<��a<�a<	�a<Ɲa<��a<W�a<%�a<��a<U�a<�a<��a<��a<?�a<l�a<v�a<��a<�a<�a<y�a<��a<՜a<ٜa<��a<֜a<}�a<9�a<��a<d�a<��a<]�a<ߙa<x�a</�a<Ҙa<�a<˘a<��a<
�a< �a<s�a<q�a<��a<u�a<��a<)�a<ǘa<b�a<Ηa<U�a<��a<#�a<w�a<�a<��a<�a<�a<˓a<�a<��a<��a<Ǔa<��a<��a<(�a<�a<X�a<ɑa<�a<J�a<��a<|�a<ݍa<�a<F�a<��a<�a<��a<(�a<�a<��a<��a<G�a<��a<��a<3�a<�a<�a<p�a<��a<ʄa<ރa<�a<4�a<>�a<��a<�a<qa<)a<�~a<�~a<a~a<x~a<H~a<)~a<�}a<�}a<}}a<�|a<Y|a<�{a<{a<Gza<�ya<ya<gxa<xa<�wa<jwa<Uwa<Mwa<ywa<hwa<�wa<�wa<xa<xa<xa<xa<�wa<}wa<wa<�va<>va<�ua<�ua<Wua<Iua<
ua<Oua<wua<�ua<5va<�va<(wa<�  �  Ewa<�wa<7xa<}xa<�xa<�xa<ya<ya<ya<ya<�xa<�xa<ya<Cya<�ya<�ya<Vza<�za<�{a<X|a<}a<�}a<T~a<�~a<Pa<�a<�a<*�a<5�a<U�a<k�a<��a<��a<�a<w�a<�a<��a<d�a<X�a<I�a<>�a<V�a<S�a<G�a<�a<يa<��a<)�a<��a<�a<I�a<��a<�a<#�a<��a<#�a<��a<X�a<��a<�a<��a<��a<J�a<��a<��a<,�a<��a<Җa<�a<%�a<�a<�a<��a<�a<ܖa<�a</�a<l�a<×a<;�a<Ԙa<h�a<�a<��a<6�a<��a<�a<I�a<i�a<��a<Z�a<E�a<�a<�a<��a<��a<��a<��a<��a<ӛa<�a<z�a<͜a<*�a<r�a<��a<�a<��a<ٝa<��a<��a<&�a<��a<B�a<ߛa<u�a< �a<�a<ޚa<֚a<�a<�a<p�a<��a<�a<^�a<��a<Мa<Μa<ڜa<��a<k�a<�a<��a<A�a<Ϛa<E�a<��a<��a<��a<j�a<M�a<Z�a<��a<��a<��a<��a<˙a<��a<y�a<�a<��a<<�a<��a<�a<<�a<��a<�a<h�a<�a<��a<m�a<J�a<R�a<Q�a<P�a<n�a<k�a<[�a<�a<ڒa<x�a<�a<R�a<��a<ߏa<�a<G�a<a�a<��a<"�a<��a<�a<��a<p�a<*�a<�a<��a<>�a<�a<Z�a<Ça<�a<H�a<j�a<u�a<v�a<��a<��a<��a<�a<wa<�~a<�~a<K~a<3~a<~a<~a< ~a<~a<�}a<�}a<b}a<�|a<�|a<�{a<\{a<�za<'za<zya<�xa<�xa<8xa<�wa<�wa<�wa<�wa<�wa<xa<&xa<7xa<>xa<#xa<�wa<�wa<Zwa<�va<kva<�ua<�ua<ua<�ta<�ta<�ta<�ta<�ta<?ua<�ua<1va<�va<�  �  wa<�wa<xa<�xa<�xa<!ya<Aya<cya<Pya<Zya<Zya<vya<�ya<�ya<za<Qza<�za<h{a<|a<�|a<M}a<�}a<u~a<a<Ma<�a<�a<�a<�a<�a<�a<�a<J�a<��a<�a<��a<�a<�a<̓a<�a<�a<�a<�a<
�a<�a<يa<��a<4�a<ƌa<@�a<��a<��a<G�a<Ďa<�a<��a<6�a<Ɛa<��a<G�a<�a<��a<��a<>�a<ƕa<O�a<��a<ݖa<ߖa<�a<֖a<��a<��a<a�a<��a<p�a<��a<�a<H�a<їa<N�a<�a<��a<c�a<�a<~�a<��a<C�a<��a<��a<��a<��a<`�a<I�a<$�a< �a<�a<�a<�a<W�a<��a<Ԝa<,�a<i�a<ȝa<�a<�a<�a<ٝa<��a<?�a<�a<c�a<��a<z�a<��a<a<b�a<`�a<D�a<�a<��a< �a<l�a<��a<+�a<d�a<��a<ќa<�a<Ӝa<��a<d�a<�a<��a<,�a<ښa<��a<%�a<	�a<͙a<�a<ՙa<�a<�a<�a<
�a<�a<ԙa<v�a<�a<��a<�a<Z�a<��a<�a<�a<��a<�a<w�a<4�a<�a<��a<ƒa<��a<�a<�a<6�a<�a<�a<ڒa<��a<�a<��a<�a<�a<t�a<��a<�a<2�a<��a<�a<��a<D�a<ӊa<��a<�a<�a<|�a<��a<}�a<��a<�a<�a<0�a</�a< �a<3�a<�a<a�a<�a<�~a<h~a<~a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<[}a<'}a<�|a<4|a<�{a<{a<}za<�ya<�ya<�xa<�xa<kxa<Wxa<Sxa<@xa<Uxa<Uxa<{xa<mxa<Wxa<4xa<�wa<�wa<wa<�va<va<�ua<ua<�ta<nta<ta<,ta<(ta<�ta<�ta<Mua<�ua<bva<�  �  �va<jwa<�wa<xa<�xa<&ya<jya<�ya<�ya<�ya<�ya<�ya<�ya<&za<�za<�za<G{a<�{a<j|a<�|a<�}a<~a<�~a<a<[a<�a<�a<�a<�a<�a<�a<�a<�a<%�a<��a<��a<��a<��a<v�a<��a<��a<��a<�a<�a<�a<�a<��a<N�a<�a<y�a<��a<L�a<��a<�a<��a<�a<��a<>�a<�a<��a<i�a<�a<ߔa<n�a<�a<T�a<��a<��a<Ėa<��a<��a<T�a<1�a<�a<	�a<�a<*�a<{�a<��a<b�a<�a<��a<Q�a<�a<Úa<^�a<ڛa<P�a<��a<��a<ќa<�a<��a<��a<��a<y�a<t�a<��a<��a<��a<��a<A�a<}�a<ŝa<�a<�a<�a<�a<ܝa<��a<%�a<��a<$�a<��a<�a<��a<E�a<��a<ٙa<ܙa<	�a<B�a<��a<��a<u�a<�a<D�a<��a<Мa<�a<؜a<Ɯa<��a<L�a<�a<��a<:�a<ݚa<��a<��a<Q�a<>�a<A�a<I�a<B�a<W�a<2�a<�a<әa<��a< �a<r�a<˗a<�a<>�a<w�a<˔a<�a<��a<�a<��a<|�a<u�a<o�a<��a<��a<Ғa<��a<�a<��a<�a<��a<,�a<��a<)�a<v�a<ŏa<�a<V�a<��a<�a<��a<�a<��a<6�a<݊a<}�a<,�a<��a<�a<��a<·a<�a<��a<��a<�a<Ƃa<a<ƀa<�a<a<s~a< ~a<�}a<r}a<_}a<T}a<]}a<�}a<�}a<�}a<~}a<h}a<%}a<�|a<a|a<�{a<`{a<�za<[za<�ya<xya<2ya<�xa<�xa<�xa<�xa<�xa<�xa<�xa<�xa<cxa<<xa<�wa<nwa<�va<rva<�ua</ua<�ta<Ata<�sa<�sa<�sa<�sa<ta<hta<�ta<sua<$va<�  �  �va<Uwa<�wa<sxa<�xa<5ya<�ya<�ya<�ya<�ya<za<za<Bza<�za<�za<3{a<�{a<|a<�|a<.}a<�}a<8~a<�~a< a<ma<wa<�a<�a<xa<�a<la<�a<�a<�a<5�a<��a<p�a<'�a<6�a<D�a<p�a<��a<��a<�a<׉a<݊a<��a<u�a<�a<��a< �a<��a<�a<[�a<�a<e�a<�a<��a<4�a<�a<��a<\�a<��a<��a<�a<Q�a<��a<��a<��a<��a<c�a<;�a<�a<֕a<��a<��a<ܕa<$�a<��a<�a<ŗa<c�a<C�a<ߙa<��a<X�a<ța<d�a<��a<�a<�a<�a<��a<�a<ޜa<��a<Ҝa<��a<�a<�a<;�a<��a<��a<�a<�a<?�a<,�a<�a<ѝa<x�a<�a<k�a<�a<\�a<ߚa<O�a<ݙa<��a<��a<��a<��a<�a<k�a<Ěa<Y�a<��a<0�a<��a<Üa<�a<�a<��a<��a<��a<�a<�a<z�a<3�a< �a<��a<��a<��a<��a<��a<y�a<�a<P�a<E�a<ҙa<��a<�a<k�a<��a<ϖa<-�a<=�a<��a<��a<)�a<��a<b�a<=�a<�a<0�a<L�a<��a<��a<��a< �a<�a<ޒa<��a<T�a<בa<A�a<��a<��a<`�a<��a<�a<c�a<Ќa<d�a<ڋa<��a<�a<��a<B�a<ŉa<E�a<~�a<Їa<Άa<��a<ʄa<��a<��a<��a<��a<�a<�~a<%~a<�}a<I}a<}a<#}a<}a<N}a<H}a<m}a<�}a<m}a<}}a< }a<�|a<�|a<|a<�{a< {a<�za<za<�ya<hya<Dya<ya<�xa<�xa<�xa<�xa<�xa<�xa<xa<<xa<�wa<`wa<�va<&va<�ua<ua<�ta<�sa<�sa<vsa<Psa<�sa<�sa<ta<�ta<@ua<va<�  �  zva<2wa<�wa<sxa<�xa<Lya<�ya<�ya<za<za<1za<Zza<�za<�za<�za<W{a<�{a<P|a<�|a<Z}a<�}a<a~a<�~a<a<ia<{a<�a<ta<ia<aa<Ea<Ba<aa<�a<�a<w�a</�a<�a<��a<�a<?�a<k�a<��a<Ɉa<��a<ߊa<��a<�a<)�a<Ía<I�a<��a<)�a<��a<�a<��a<�a<ʑa<��a<+�a<֓a<��a<%�a<��a<�a<h�a<��a<��a<��a<f�a<8�a<�a<a<��a<��a<��a<��a<ޕa<Z�a<�a<��a<8�a<�a<ƙa<|�a<>�a<ϛa<_�a<��a<��a<�a<*�a< �a<�a<�a<�a<��a<��a<�a<S�a<��a<��a<�a<�a<E�a<K�a<>�a<�a<֝a<|�a<��a<Z�a<Λa<7�a<��a<�a<ƙa<t�a<L�a<S�a<��a<a<*�a<��a<�a<��a<�a<��a<Ĝa<��a<��a<��a<ۜa<��a<N�a<�a<��a<�a<$�a<�a<Ԛa<ݚa<��a<��a<��a<��a<y�a<M�a<�a<��a<��a<X�a<��a<��a<��a<�a<J�a<��a<�a<y�a<&�a<��a<��a<�a<�a<Q�a<��a<��a<ݒa<�a<��a<��a<]�a<�a<t�a<ߐa<.�a<��a<�a<3�a<��a<��a<��a<,�a<��a<J�a<�a<r�a<�a<M�a<��a<χa<چa<ԅa<��a<��a<x�a<T�a<H�a<ia<�~a<�}a<c}a<"}a<�|a<�|a<�|a<}a</}a<I}a<u}a<t}a<x}a<5}a<}a<�|a<A|a<�{a<J{a<�za<xza<�ya<�ya<hya<Sya<7ya<ya<ya<
ya<�xa<�xa<�xa<Ixa<�wa<cwa<�va<va<{ua<�ta<Dta<�sa<rsa<-sa<sa<7sa<�sa<�sa<xta<ua<�ua<�  �  �va<8wa<�wa<\xa<�xa<cya<�ya<�ya<�ya<4za<6za<Yza<�za<�za<A{a<`{a<�{a<E|a<�|a<r}a<�}a<j~a<�~a<.a<Ua<oa<�a<�a<�a<<a<Fa<-a<Ma<�a<�a<w�a<	�a<�a<�a<�a<-�a<c�a<��a<ňa<Љa<��a<ċa<��a<4�a<ōa<B�a<Ўa<#�a<��a<�a<��a<T�a<Ǒa<��a< �a<�a<��a<$�a<��a<�a<r�a<~�a<��a<��a<��a<<�a<�a<˕a<}�a<��a<c�a<��a<ؕa<D�a<Ԗa<i�a<=�a<�a<ٙa<��a<9�a<ƛa<F�a<��a<�a<�a<-�a<2�a<*�a<��a<�a<��a<C�a</�a<Q�a<��a<��a<	�a<�a<I�a<K�a<M�a<�a<��a<n�a<��a<��a<��a<+�a<��a<�a<��a<O�a<R�a<2�a<x�a<��a<�a<��a<�a<��a<�a<y�a<��a<�a<�a<��a<�a<��a<p�a<�a<��a<|�a<6�a<>�a<ݚa<ܚa<��a<Ěa<��a<��a<��a<J�a<�a<~�a<�a<R�a<��a<ؖa<ҕa<�a<5�a<��a<�a<k�a<'�a<֑a<�a<ܑa<�a<?�a<z�a<͒a<ْa<ݒa<��a<��a<e�a<��a<u�a<ؐa<I�a<~�a<�a<3�a<��a<4�a<��a<6�a<��a<`�a<�a<q�a<��a<O�a<��a<��a<͆a<ͅa<˄a<��a<e�a<\�a<3�a<`a<u~a<�}a<]}a<}a<�|a<�|a<�|a<�|a<C}a<X}a<o}a<k}a<^}a<N}a< }a<�|a<D|a<�{a<]{a<�za<|za<za<�ya<�ya<Pya<?ya<ya<2ya<�xa<�xa<�xa<�xa<Cxa<�wa<Vwa<�va<>va<dua<�ta<6ta<�sa<fsa<sa<sa<sa<{sa<�sa<eta<ua<�ua<�  �  zva<2wa<�wa<sxa<�xa<Lya<�ya<�ya<za<za<1za<Zza<�za<�za<�za<W{a<�{a<P|a<�|a<Z}a<�}a<a~a<�~a<a<ia<{a<�a<ta<ia<aa<Ea<Ba<aa<�a<�a<w�a</�a<�a<��a<�a<?�a<k�a<��a<Ɉa<��a<ߊa<��a<�a<)�a<Ía<I�a<��a<)�a<��a<�a<��a<�a<ʑa<��a<+�a<֓a<��a<%�a<��a<�a<h�a<��a<��a<��a<f�a<8�a<�a<a<��a<��a<��a<��a<ޕa<Z�a<�a<��a<8�a<�a<ƙa<|�a<>�a<ϛa<_�a<��a<��a<�a<*�a< �a<�a<�a<�a<��a<��a<�a<S�a<��a<��a<�a<�a<E�a<K�a<>�a<�a<֝a<|�a<��a<Z�a<Λa<7�a<��a<�a<ƙa<t�a<L�a<S�a<��a<a<*�a<��a<�a<��a<�a<��a<Ĝa<��a<��a<��a<ۜa<��a<N�a<�a<��a<�a<$�a<�a<Ԛa<ݚa<��a<��a<��a<��a<y�a<M�a<�a<��a<��a<X�a<��a<��a<��a<�a<J�a<��a<�a<y�a<&�a<��a<��a<�a<�a<Q�a<��a<��a<ݒa<�a<��a<��a<]�a<�a<t�a<ߐa<.�a<��a<�a<3�a<��a<��a<��a<,�a<��a<J�a<�a<r�a<�a<M�a<��a<χa<چa<ԅa<��a<��a<x�a<T�a<H�a<ia<�~a<�}a<c}a<"}a<�|a<�|a<�|a<}a</}a<I}a<u}a<t}a<x}a<5}a<}a<�|a<A|a<�{a<J{a<�za<xza<�ya<�ya<hya<Sya<7ya<ya<ya<
ya<�xa<�xa<�xa<Ixa<�wa<cwa<�va<va<{ua<�ta<Dta<�sa<rsa<-sa<sa<7sa<�sa<�sa<xta<ua<�ua<�  �  �va<Uwa<�wa<sxa<�xa<5ya<�ya<�ya<�ya<�ya<za<za<Bza<�za<�za<3{a<�{a<|a<�|a<.}a<�}a<8~a<�~a< a<ma<wa<�a<�a<xa<�a<la<�a<�a<�a<5�a<��a<p�a<'�a<6�a<D�a<p�a<��a<��a<�a<׉a<݊a<��a<u�a<�a<��a< �a<��a<�a<[�a<�a<e�a<�a<��a<4�a<�a<��a<\�a<��a<��a<�a<Q�a<��a<��a<��a<��a<c�a<;�a<�a<֕a<��a<��a<ܕa<$�a<��a<�a<ŗa<c�a<C�a<ߙa<��a<X�a<ța<d�a<��a<�a<�a<�a<��a<�a<ޜa<��a<Ҝa<��a<�a<�a<;�a<��a<��a<�a<�a<?�a<,�a<�a<ѝa<x�a<�a<k�a<�a<\�a<ߚa<O�a<ݙa<��a<��a<��a<��a<�a<k�a<Ěa<Y�a<��a<0�a<��a<Üa<�a<�a<��a<��a<��a<�a<�a<z�a<3�a< �a<��a<��a<��a<��a<��a<y�a<�a<P�a<E�a<ҙa<��a<�a<k�a<��a<ϖa<-�a<=�a<��a<��a<)�a<��a<b�a<=�a<�a<0�a<L�a<��a<��a<��a< �a<�a<ޒa<��a<T�a<בa<A�a<��a<��a<`�a<��a<�a<c�a<Ќa<d�a<ڋa<��a<�a<��a<B�a<ŉa<E�a<~�a<Їa<Άa<��a<ʄa<��a<��a<��a<��a<�a<�~a<%~a<�}a<I}a<}a<#}a<}a<N}a<H}a<m}a<�}a<m}a<}}a< }a<�|a<�|a<|a<�{a< {a<�za<za<�ya<hya<Dya<ya<�xa<�xa<�xa<�xa<�xa<�xa<xa<<xa<�wa<`wa<�va<&va<�ua<ua<�ta<�sa<�sa<vsa<Psa<�sa<�sa<ta<�ta<@ua<va<�  �  �va<jwa<�wa<xa<�xa<&ya<jya<�ya<�ya<�ya<�ya<�ya<�ya<&za<�za<�za<G{a<�{a<j|a<�|a<�}a<~a<�~a<a<[a<�a<�a<�a<�a<�a<�a<�a<�a<%�a<��a<��a<��a<��a<v�a<��a<��a<��a<�a<�a<�a<�a<��a<N�a<�a<y�a<��a<L�a<��a<�a<��a<�a<��a<>�a<�a<��a<i�a<�a<ߔa<n�a<�a<T�a<��a<��a<Ėa<��a<��a<T�a<1�a<�a<	�a<�a<*�a<{�a<��a<b�a<�a<��a<Q�a<�a<Úa<^�a<ڛa<P�a<��a<��a<ќa<�a<��a<��a<��a<y�a<t�a<��a<��a<��a<��a<A�a<}�a<ŝa<�a<�a<�a<�a<ܝa<��a<%�a<��a<$�a<��a<�a<��a<E�a<��a<ٙa<ܙa<	�a<B�a<��a<��a<u�a<�a<D�a<��a<Мa<�a<؜a<Ɯa<��a<L�a<�a<��a<:�a<ݚa<��a<��a<Q�a<>�a<A�a<I�a<B�a<W�a<2�a<�a<әa<��a< �a<r�a<˗a<�a<>�a<w�a<˔a<�a<��a<�a<��a<|�a<u�a<o�a<��a<��a<Ғa<��a<�a<��a<�a<��a<,�a<��a<)�a<v�a<ŏa<�a<V�a<��a<�a<��a<�a<��a<6�a<݊a<}�a<,�a<��a<�a<��a<·a<�a<��a<��a<�a<Ƃa<a<ƀa<�a<a<s~a< ~a<�}a<r}a<_}a<T}a<]}a<�}a<�}a<�}a<~}a<h}a<%}a<�|a<a|a<�{a<`{a<�za<[za<�ya<xya<2ya<�xa<�xa<�xa<�xa<�xa<�xa<�xa<�xa<cxa<<xa<�wa<nwa<�va<rva<�ua</ua<�ta<Ata<�sa<�sa<�sa<�sa<ta<hta<�ta<sua<$va<�  �  wa<�wa<xa<�xa<�xa<!ya<Aya<cya<Pya<Zya<Zya<vya<�ya<�ya<za<Qza<�za<h{a<|a<�|a<M}a<�}a<u~a<a<Ma<�a<�a<�a<�a<�a<�a<�a<J�a<��a<�a<��a<�a<�a<̓a<�a<�a<�a<�a<
�a<�a<يa<��a<4�a<ƌa<@�a<��a<��a<G�a<Ďa<�a<��a<6�a<Ɛa<��a<G�a<�a<��a<��a<>�a<ƕa<O�a<��a<ݖa<ߖa<�a<֖a<��a<��a<a�a<��a<p�a<��a<�a<H�a<їa<N�a<�a<��a<c�a<�a<~�a<��a<C�a<��a<��a<��a<��a<`�a<I�a<$�a< �a<�a<�a<�a<W�a<��a<Ԝa<,�a<i�a<ȝa<�a<�a<�a<ٝa<��a<?�a<�a<c�a<��a<z�a<��a<a<b�a<`�a<D�a<�a<��a< �a<l�a<��a<+�a<d�a<��a<ќa<�a<Ӝa<��a<d�a<�a<��a<,�a<ښa<��a<%�a<	�a<͙a<�a<ՙa<�a<�a<�a<
�a<�a<ԙa<v�a<�a<��a<�a<Z�a<��a<�a<�a<��a<�a<w�a<4�a<�a<��a<ƒa<��a<�a<�a<6�a<�a<�a<ڒa<��a<�a<��a<�a<�a<t�a<��a<�a<2�a<��a<�a<��a<D�a<ӊa<��a<�a<�a<|�a<��a<}�a<��a<�a<�a<0�a</�a< �a<3�a<�a<a�a<�a<�~a<h~a<~a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<[}a<'}a<�|a<4|a<�{a<{a<}za<�ya<�ya<�xa<�xa<kxa<Wxa<Sxa<@xa<Uxa<Uxa<{xa<mxa<Wxa<4xa<�wa<�wa<wa<�va<va<�ua<ua<�ta<nta<ta<,ta<(ta<�ta<�ta<Mua<�ua<bva<�  �  Ewa<�wa<7xa<}xa<�xa<�xa<ya<ya<ya<ya<�xa<�xa<ya<Cya<�ya<�ya<Vza<�za<�{a<X|a<}a<�}a<T~a<�~a<Pa<�a<�a<*�a<5�a<U�a<k�a<��a<��a<�a<w�a<�a<��a<d�a<X�a<I�a<>�a<V�a<S�a<G�a<�a<يa<��a<)�a<��a<�a<I�a<��a<�a<#�a<��a<#�a<��a<X�a<��a<�a<��a<��a<J�a<��a<��a<,�a<��a<Җa<�a<%�a<�a<�a<��a<�a<ܖa<�a</�a<l�a<×a<;�a<Ԙa<h�a<�a<��a<6�a<��a<�a<I�a<i�a<��a<Z�a<E�a<�a<�a<��a<��a<��a<��a<��a<ӛa<�a<z�a<͜a<*�a<r�a<��a<�a<��a<ٝa<��a<��a<&�a<��a<B�a<ߛa<u�a< �a<�a<ޚa<֚a<�a<�a<p�a<��a<�a<^�a<��a<Мa<Μa<ڜa<��a<k�a<�a<��a<A�a<Ϛa<E�a<��a<��a<��a<j�a<M�a<Z�a<��a<��a<��a<��a<˙a<��a<y�a<�a<��a<<�a<��a<�a<<�a<��a<�a<h�a<�a<��a<m�a<J�a<R�a<Q�a<P�a<n�a<k�a<[�a<�a<ڒa<x�a<�a<R�a<��a<ߏa<�a<G�a<a�a<��a<"�a<��a<�a<��a<p�a<*�a<�a<��a<>�a<�a<Z�a<Ça<�a<H�a<j�a<u�a<v�a<��a<��a<��a<�a<wa<�~a<�~a<K~a<3~a<~a<~a< ~a<~a<�}a<�}a<b}a<�|a<�|a<�{a<\{a<�za<'za<zya<�xa<�xa<8xa<�wa<�wa<�wa<�wa<�wa<xa<&xa<7xa<>xa<#xa<�wa<�wa<Zwa<�va<kva<�ua<�ua<ua<�ta<�ta<�ta<�ta<�ta<?ua<�ua<1va<�va<�  �  {wa<�wa<Axa<�xa<�xa<�xa<�xa<�xa<�xa<xxa<�xa<|xa<�xa<�xa<�xa<oya<�ya<�za<-{a<�{a<�|a<Z}a<~a<�~a<ba<�a<�a<P�a<x�a<��a<��a<�a<>�a<��a<��a<p�a<E�a<�a<�a<��a<��a<��a<��a<r�a<�a<�a<f�a<�a<J�a<��a<�a<�a<��a<��a<(�a<��a<�a<ݏa<��a<|�a<&�a<#�a<��a<��a<~�a<�a<Ŗa<��a<9�a<P�a<q�a<m�a<R�a<~�a<]�a<��a<��a<�a<b�a<��a<`�a<��a<m�a<ޚa<[�a<��a<�a<e�a<7�a<K�a<�a<�a<��a<m�a<Q�a<�a<�a<��a<�a<U�a<��a<�a<?�a<ٜa<�a<��a<��a<�a<	�a<Ɲa<��a<W�a<%�a<��a<U�a<�a<��a<��a<?�a<l�a<v�a<��a<�a<�a<y�a<��a<՜a<ٜa<��a<֜a<}�a<9�a<��a<d�a<��a<]�a<ߙa<x�a</�a<Ҙa<�a<˘a<��a<
�a< �a<s�a<q�a<��a<u�a<��a<)�a<ǘa<b�a<Ηa<U�a<��a<#�a<w�a<�a<��a<�a<�a<˓a<�a<��a<��a<Ǔa<��a<��a<(�a<�a<X�a<ɑa<�a<J�a<��a<|�a<ݍa<�a<F�a<��a<�a<��a<(�a<�a<��a<��a<G�a<��a<��a<3�a<�a<�a<p�a<��a<ʄa<ރa<�a<4�a<>�a<��a<�a<qa<)a<�~a<�~a<a~a<x~a<H~a<)~a<�}a<�}a<}}a<�|a<Y|a<�{a<{a<Gza<�ya<ya<gxa<xa<�wa<jwa<Uwa<Mwa<ywa<hwa<�wa<�wa<xa<xa<xa<xa<�wa<}wa<wa<�va<>va<�ua<�ua<Wua<Iua<
ua<Oua<wua<�ua<5va<�va<(wa<�  �  �wa<,xa<uxa<�xa<�xa<�xa<�xa<�xa<Wxa<(xa<xa<�wa<�wa<%xa<rxa<�xa<Mya<�ya<�za<z{a<\|a<*}a<�}a<�~a<0a<�a<<�a<��a<̀a<�a<C�a<��a<��a<�a<��a<�a<Ńa<h�a<H�a<7�a<�a<��a<ňa<��a<L�a<�a<R�a<ʋa<#�a<O�a<��a<��a<��a<-�a<��a<�a<��a<:�a<�a<�a<Ցa<��a<��a<��a<Y�a<��a<��a<
�a<u�a<��a<��a<ӗa<��a<�a<ܗa<�a<F�a<��a<ۘa<1�a<˙a<B�a<Úa<3�a<��a<��a<#�a<3�a<.�a<"�a<�a<��a<A�a< �a<��a<��a<j�a<z�a<��a<��a<�a<��a<�a<o�a<ޜa<]�a<��a<Ɲa<��a<��a<�a<��a<l�a< �a<Ӝa<j�a<+�a<�a<�a<��a<��a<�a<\�a<��a<ǜa<�a<�a<�a<��a<��a<q�a<�a<��a<��a<c�a<�a<T�a<�a<��a<o�a<J�a<C�a<g�a<��a<Ęa<�a<A�a<p�a<o�a<Y�a<D�a<�a<��a<"�a<��a<�a<��a<�a<��a<�a<Δa<��a<N�a<A�a<?�a<(�a<�a<ݓa<��a<X�a<�a<D�a<��a<�a<��a<�a<3�a<Q�a<j�a<��a<�a<�a<��a<��a<z�a<I�a<�a<��a<шa<��a<$�a<Ƈa<9�a<��a<څa<�a<E�a<q�a<��a<��a<#�a<��a<�a<�a<Aa<)a<�~a<�~a<�~a<g~a<4~a<�}a<K}a<�|a<1|a<w{a<�za<�ya<4ya<�xa<�wa<nwa<"wa<�va<�va<�va<�va<wa<[wa<�wa<�wa<�wa<�wa<xa<�wa<�wa<]wa<wa<�va<tva<va<�ua<�ua<�ua<�ua<�ua<2va<�va<wa<vwa<�  �  "xa<Zxa<�xa<�xa<�xa<�xa<lxa<Pxa<�wa<�wa<�wa<xwa<�wa<�wa<�wa<Axa<�xa<}ya<Wza<1{a<|a<�|a<�}a<�~a</a<�a<P�a<��a<!�a<O�a<��a<�a<J�a<��a<�a<��a<&�a<�a<��a<��a<V�a<C�a<�a<��a<x�a<�a<`�a<��a<�a<�a<%�a<i�a<l�a<Ōa<
�a<��a<�a<��a<��a<`�a<�a<a�a<j�a<V�a<-�a<�a<��a<1�a<��a<՗a<�a<�a<>�a<L�a<{�a<{�a<ǘa< �a<Q�a<љa<%�a<��a<��a<��a<՛a<�a<<�a<2�a<,�a<ߛa<��a<P�a<��a<��a<:�a<*�a<�a<��a<�a<L�a<��a<
�a<��a<�a<��a<�a<��a<ϝa<��a<"�a<	�a<��a<��a<k�a<)�a<�a<��a<u�a<x�a<[�a<��a<��a<��a<�a<�a<;�a<5�a<1�a<��a<��a<U�a<Ǜa<P�a<��a<�a<n�a<ܘa<|�a<�a<�a<��a<�a<�a<5�a<|�a<��a<�a<'�a<c�a<X�a<X�a<�a<јa<w�a<�a<y�a<�a<��a<��a<��a<R�a<�a<�a<��a<��a<i�a<[�a<$�a<ѓa<��a<�a<R�a<��a<��a<ɏa<��a<�a<Ȍa<�a<)�a<��a<��a<}�a<G�a<�a<�a<��a<��a<��a<`�a<0�a<a<`�a<��a<�a<e�a<�a<΃a<�a<\�a<��a<�a<��a<�a<�a<�a<\a<	a<�~a<�~a<?~a<�}a<K}a<�|a<�{a<B{a<hza<�ya<�xa<xa<�wa<�va<�va<Sva<Lva<Tva<vva<�va<�va<awa<�wa<�wa<�wa<xa<	xa<�wa<�wa<^wa<wa<�va<�va<kva<-va<Cva<>va<�va<�va<wa<_wa<�wa<�  �  Ixa<�xa<�xa<�xa<�xa<xa<Jxa<xa<�wa<hwa<Cwa<wa<wa<,wa<lwa<�wa<sxa<!ya<�ya<�za<�{a<�|a<�}a<i~a<4a<�a<`�a<�a<L�a<��a<��a<L�a<��a<��a<�a<�a<��a<]�a<#�a<�a<��a<��a<<�a<݉a<v�a<�a<:�a<��a<��a<ҋa<ыa<�a<�a<T�a<��a<�a<��a<R�a<.�a<�a<
�a<	�a<#�a<"�a<�a<ڕa<��a<5�a<��a<�a<W�a<m�a<��a<��a<Ҙa<��a<9�a<{�a<��a<(�a<��a<��a<\�a<��a<�a<�a<E�a<:�a<�a<ța<x�a<�a<��a<?�a<�a<��a<x�a<q�a<��a<�a<9�a<��a<1�a<Ǜa<m�a<�a<`�a<��a<�a<"�a<-�a<�a<	�a<��a<��a<T�a<�a<��a<�a<֜a<ݜa<�a<$�a<6�a<a�a<b�a<^�a<5�a<�a<��a<1�a<��a<�a<[�a<��a<�a<z�a<	�a<��a<h�a<U�a<h�a<��a<՗a<�a<t�a<Әa<�a<:�a<\�a<^�a<(�a<��a<��a<@�a<ɗa<S�a<ޖa<b�a<�a<ƕa<w�a<C�a<�a<��a<Ɣa<��a<T�a<�a<��a<�a<,�a<e�a<z�a<��a<g�a<l�a<y�a<��a<a<�a<�a<�a<Ԉa<��a<~�a<g�a<o�a<`�a<C�a<�a<Їa<c�a<نa<J�a<��a<߄a<$�a<g�a<��a<	�a<��a< �a<��a<8�a<�a<�a<ga<$a<�~a<W~a<�}a<S}a<�|a<�{a<	{a<za<7ya<txa<�wa<wa<|va<va<�ua<�ua<�ua<$va<Zva<�va< wa<mwa<�wa<�wa<xa<
xa<�wa<�wa<�wa<cwa<3wa<�va<�va<�va<�va<�va<�va<&wa<qwa<�wa<xa<�  �  fxa<�xa<�xa<�xa<�xa<uxa<1xa<�wa<�wa<3wa<wa<�va<�va<�va<wa<�wa<xa<�xa<�ya<�za<�{a<r|a<�}a<Z~a<*a<�a<��a<�a<p�a<�a<*�a<��a<�a<Z�a<ڃa<O�a<	�a<��a<r�a<.�a<�a<��a<X�a<�a<p�a<�a<'�a<��a<��a<��a<ċa<��a<�a<��a<H�a<��a<O�a<�a<Ŏa<׏a<ːa<��a<��a<��a<�a<ƕa<��a<0�a<їa<�a<l�a<��a<Ҙa<�a<�a<Z�a<z�a<̙a<�a<h�a<�a<-�a<��a<֛a<�a<F�a<C�a<1�a<�a<a<8�a<�a<n�a<��a<��a<@�a<:�a<#�a<O�a<�a<ޙa<~�a<��a<��a< �a<˜a<W�a<��a<�a<&�a<b�a<8�a<7�a<��a<؝a<��a<g�a<U�a<#�a<8�a<1�a<B�a<l�a<k�a<��a<�a<��a<?�a<�a<��a<'�a<��a<Śa<C�a<n�a<ݘa<%�a<��a<b�a<�a<�a<�a<B�a<��a<�a<S�a<��a<�a<+�a<R�a<]�a<I�a< �a<Ƙa<��a<��a<��a<�a<��a<g�a<��a<֕a<��a<l�a<6�a< �a<Ɣa<p�a<'�a<}�a<�a<�a<^�a<T�a<J�a<Z�a<-�a<>�a<-�a<f�a<��a<0�a<Ȉa<k�a<c�a<>�a<T�a<A�a<4�a<>�a<�a<هa<^�a<�a<b�a<Ņa<�a<b�a<��a<�a<l�a<Áa<Q�a<�a<x�a<@�a<�a<�a<@a<�~a<}~a<�}a<J}a<�|a<�{a<�za<�ya<ya<2xa<fwa<�va<>va<�ua<�ua<�ua<�ua<�ua<"va<�va<�va<Kwa<�wa<�wa<xa<xa<0xa<�wa<�wa<�wa<ywa<>wa<wa<wa<�va<wa<2wa<gwa<�wa<�wa<Fxa<�  �  �xa<�xa<�xa<�xa<�xa<nxa<xa<�wa<gwa<wa<�va<�va<�va<�va<�va<Swa<�wa<�xa<ya<sza<l{a<_|a<i}a<_~a<.a<�a<��a<�a<��a<�a<`�a<��a<,�a<��a<��a<��a<2�a<�a<��a<[�a<�a<؈a<}�a<�a<��a<��a<1�a<d�a<f�a<z�a<��a<��a<��a<ڋa< �a<z�a<�a<Ӎa<��a<��a<��a<��a<˒a<Փa<�a<ҕa<��a<F�a<ٗa<B�a<��a<ؘa<�a<1�a<e�a<��a<��a<�a<Q�a<��a<�a<b�a<��a<�a<5�a<R�a<V�a<4�a<��a<��a< �a<��a<@�a<șa<`�a<(�a<��a<�a<�a<[�a<��a<9�a<Қa<}�a<�a<��a<H�a<��a<�a<;�a<j�a<c�a<V�a<%�a<��a<ҝa<��a<y�a<]�a<]�a<��a<��a<��a<��a<��a<��a<��a<V�a<�a<��a<!�a<k�a<��a<�a<J�a<��a<��a<��a<�a<ݖa<Ζa<�a<�a<\�a<��a<�a<v�a<��a<0�a<V�a<l�a<X�a<.�a<��a<��a<1�a<×a<e�a<��a<��a<7�a<��a<ڕa<��a<d�a<-�a<�a<��a<.�a<��a<��a<"�a<C�a</�a<+�a<!�a< �a<��a<�a<>�a<y�a<�a<��a<T�a<�a<�a<�a<�a<�a<�a<��a<Շa<t�a<�a<��a<�a<I�a<��a<�a<F�a<��a<��a<s�a<�a<Àa<c�a<�a<�a<qa<a<�~a<�}a<M}a<�|a<�{a<�za<�ya<�xa<�wa<*wa<�va<�ua<�ua<Wua<\ua<lua<�ua<�ua<iva<�va<)wa<�wa<�wa<xa<"xa<8xa<xa<xa<�wa<�wa<uwa<gwa<1wa<(wa<@wa<�wa<�wa<�wa<xa<bxa<�  �  za<%za<Nza<Aza<za<�ya<�ya<�ya<_ya<`ya<ya<ya<ya<+ya<�ya<�ya<qza<�za<�{a<�|a<Y}a<O~a<�~a<�a<��a<_�a<�a<|�a<�a<<�a<�a<�a<��a<
�a<u�a<�a<��a<`�a<ׇa<Έa<D�a<�a<a<2�a<�a<�a<o�a<��a<�a< �a<;�a<��a<��a<�a<�a<Վa<q�a<��a<��a<h�a<��a<X�a<H�a<2�a<��a<זa<��a<Y�a<��a<;�a<��a<��a<#�a<
�a<r�a<��a<Қa<�a<d�a<��a<�a<��a<��a<�a<1�a<;�a<_�a<+�a<�a<��a<��a<3�a<��a<��a<E�a<9�a<�a<T�a<1�a<Y�a<��a<�a<��a<��a<��a<�a<a�a<��a<�a<]�a<Z�a<r�a<I�a<3�a<�a<͞a<՞a<��a<��a<v�a<��a<��a<��a<��a<��a<��a<��a<q�a<�a<��a<8�a<��a<J�a<��a<+�a<~�a< �a<��a<7�a<S�a<ۘa<��a<��a<K�a<��a<��a<�a<�a<@�a<Y�a<x�a<[�a</�a<�a<u�a<`�a<��a<r�a<�a<��a<m�a<
�a<��a<��a<��a<�a<�a<��a<�a<��a<�a<6�a<`�a<��a<��a<��a<��a<��a<$�a<7�a<ߋa<b�a<��a<y�a<�a<&�a<�a<ʉa<��a<m�a<H�a<��a<Ոa<-�a<Շa<9�a<j�a<�a<!�a<��a<��a<��a<��a<��a<3�a<��a<��a< �a<��a<n�a<�a<ta<�~a<~a<A}a<�|a<�{a<{a<^za<�ya<ya<kxa<rxa<�wa<�wa<�wa<�wa<Xxa<axa<�xa<�xa<,ya<bya<�ya<�ya<�ya<�ya<qya<Rya<:ya<�xa<�xa<�xa<�xa<�xa<ya<$ya<jya<�ya<�ya<�  �  �ya<za<"za<7za<>za<+za<�ya<�ya<wya<Fya<%ya<ya<)ya<-ya<vya<�ya<~za<{a<�{a<�|a<u}a<Q~a<%a<�a<��a<H�a<؁a<Y�a<�a<N�a<��a< �a<��a<�a<��a<�a<��a<V�a<�a<��a<P�a<	�a<��a<.�a<��a<"�a<��a<،a<�a<*�a<6�a<l�a<��a<��a<H�a<��a<2�a<�a<��a<�a<k�a<K�a<V�a<D�a<%�a<��a<��a<�a<��a<�a<x�a<��a<��a<�a<h�a<��a<ݚa<�a<`�a<��a<��a<Y�a<��a<�a<�a</�a<>�a<E�a<0�a<�a<��a<M�a<�a<��a<[�a<@�a<�a<�a<�a<|�a<˛a<#�a<��a<�a<��a<�a<��a<ߞa<�a<$�a<I�a<L�a<O�a<#�a<�a<�a<מa<��a<��a<��a<��a<��a<��a<��a<��a<��a<x�a<E�a<�a<Νa<j�a<לa<L�a<��a<�a<��a<�a<��a<9�a<�a<�a<
�a<�a<B�a<p�a<��a<�a<7�a<p�a<{�a<a�a<?�a<�a<�a<��a<2�a<͘a<z�a<�a<��a<u�a<�a<�a<��a<n�a<�a<��a<r�a<
�a<w�a<�a<Z�a<��a<��a<��a<��a<׎a<��a<5�a<j�a<��a<#�a<Ċa<��a<.�a<�a<ىa<׉a<��a<��a<k�a<�a<��a<0�a<��a<*�a<��a<�a<5�a<��a<�a<��a<�a<��a<4�a<Ɂa<x�a<�a<ƀa<I�a<�a<Ta<�~a<2~a<g}a<�|a<�{a<�za<Lza<�ya<ya<�xa<$xa<�wa<�wa<�wa<xa<7xa<sxa<�xa<ya<]ya<�ya<�ya<�ya<�ya<�ya<vya<Bya<,ya<ya<�xa<�xa<�xa<�xa<ya<=ya<fya<�ya<�ya<�  �  �ya<:za<6za<Cza<'za<	za<�ya<�ya<�ya<]ya<bya<3ya<Fya<�ya<�ya</za<�za<B{a<�{a<�|a<�}a<R~a<'a<�a<��a<G�a<��a<t�a<ła<K�a<��a<�a<Z�a<Єa<W�a<Ӆa<}�a<�a<Ӈa<q�a<D�a<�a<��a<e�a<��a<:�a<s�a<ƌa<��a<E�a<p�a<��a<�a<�a<��a<�a<u�a<;�a<Đa<őa<��a<~�a<z�a<A�a<�a<֖a<��a<�a<ݘa<	�a<S�a<��a<��a<�a<�a<h�a<��a<�a<-�a<x�a<�a<�a<��a<ɜa<�a<T�a<8�a<A�a<�a<�a<��a<|�a<
�a<ӛa<��a<I�a<a�a<I�a<n�a<��a<ޛa<c�a<��a<I�a<��a<�a<x�a<Ǟa<!�a<4�a<u�a<0�a<;�a<�a<�a<��a<��a<��a<a�a<h�a<V�a<j�a<}�a<x�a<��a<w�a<��a<Y�a<�a<��a<H�a<ڜa<P�a<ޛa<(�a<Ěa<(�a<șa<��a<>�a<@�a<�a<E�a<u�a<��a<�a<�a<9�a<H�a<n�a<`�a<_�a<&�a<��a<��a<��a<��a<:�a<ޗa<��a<0�a<��a<��a<��a<2�a<�a<��a<f�a<A�a<{�a<�a<:�a<�a<��a<ېa<�a<��a<6�a<<�a<��a<�a<f�a<�a<��a<u�a<2�a<�a<��a<��a<��a<H�a<�a<��a<e�a<��a<�a<{�a<��a<%�a<`�a<߃a<F�a<ւa<_�a<�a<��a<=�a<�a<��a<U�a<�a<Na<�~a<
~a<g}a<�|a<|a<!{a<{za<�ya<#ya<�xa<gxa<6xa<xa<xa<Fxa<Rxa<�xa<�xa<ya<Cya<jya<�ya<�ya<�ya<fya<bya<$ya< ya<�xa<�xa<�xa<�xa<�xa<�xa<ya<Cya<lya<�ya<�  �  �ya<�ya<za<?za<5za</za<za<�ya<�ya<�ya<�ya<wya<~ya<�ya<�ya<Hza<�za<v{a<'|a<�|a<�}a<~~a<Ua<�a<��a<H�a<��a<H�a<��a<�a<o�a<փa< �a<��a<�a<��a<M�a<ӆa<��a<W�a<�a<Ɖa<w�a<�a<��a<6�a<�a<��a<%�a<]�a<��a<Ía<�a<F�a<��a<�a<��a<G�a<	�a<�a<ƒa<��a<��a<k�a<N�a<�a<��a<�a<~�a<�a<4�a<t�a<��a<ؙa<�a<?�a<_�a<��a<�a<A�a<��a<�a<b�a<��a<�a<�a<9�a<I�a<"�a<�a<̜a<��a<<�a<��a<ƛa<��a<q�a<��a<��a<̛a<"�a<��a<�a<Y�a<Нa<@�a<��a<Ҟa<�a<�a<&�a<�a<�a<�a<��a<��a<U�a<P�a<.�a<3�a<&�a<-�a<T�a<^�a<n�a<`�a<\�a</�a<�a<ŝa<n�a<�a<{�a<�a<[�a<�a<l�a<�a<��a<��a<X�a<`�a<y�a<��a<ęa<��a</�a<g�a<h�a<w�a<a�a<�a<��a<��a<K�a<�a<��a< �a<��a<W�a<��a<ʖa<k�a<N�a<�a<ߕa<��a<R�a<�a<p�a<�a<F�a<��a<ϑa<��a<�a</�a<_�a<��a<��a<&�a<��a<!�a<͊a<��a<d�a<5�a<�a<�a<��a<T�a<�a<��a<�a<��a<�a<B�a<��a<�a<,�a<��a<�a<��a<9�a<��a<��a<'�a<ۀa<��a<.�a<�a<Na<�~a<$~a<�}a<�|a<|a<S{a<�za<za<hya<�xa<�xa<_xa<Cxa<Lxa<jxa<�xa<�xa<�xa<9ya<kya<uya<�ya<{ya<oya<Pya<4ya<ya<�xa<�xa<{xa<�xa<txa<�xa<�xa<�xa<ya<Rya<�ya<�  �  �ya<�ya<za<3za<@za<Eza<za<za<�ya<�ya<�ya<�ya<�ya<�ya<Xza<�za<D{a<�{a<d|a<;}a<�}a<�~a<Oa<�a<��a<I�a<��a<+�a<��a<Ԃa<&�a<v�a<�a<D�a<��a<E�a<ׅa<��a<R�a<�a<͈a<��a<^�a<�a<��a<�a<��a<��a<8�a<��a<ɍa<�a<0�a<��a<��a<x�a<�a<��a<��a<�a<�a<�a<��a<��a<P�a< �a<��a<&�a<r�a<՘a<�a<3�a<]�a<��a<��a<̙a<�a<D�a<��a<�a<U�a<��a<$�a<��a<֜a<�a<B�a<7�a<B�a<�a<�a<��a<��a<@�a<��a<�a<��a<�a<�a<6�a<��a<��a<F�a<��a<��a<D�a<��a<�a<
�a<!�a<�a<�a<̞a<��a<h�a<L�a<�a<ڝa<۝a<��a<؝a<��a<��a<�a<*�a<Q�a<?�a<3�a<�a<Нa<��a<�a<��a<�a<��a<�a<��a<l�a<��a<�a<��a<Йa<��a<ڙa<�a<#�a<S�a<a�a<��a<n�a<c�a<�a<ݙa<��a<�a<��a<#�a<ȗa<R�a<�a<��a<T�a<-�a<�a<Εa<��a<i�a<:�a<͔a<��a<�a<b�a<��a<�a<�a<K�a<��a<��a<��a< �a<��a<��a<|�a<K�a<Ċa<��a<s�a<7�a<��a<Éa<q�a<�a<��a<��a<p�a<��a< �a<M�a<��a<�a<C�a<��a<2�a<Ёa<��a< �a<߀a<��a<_�a<�a<�a<Wa<�~a<D~a<�}a<�|a<9|a<�{a<�za<2za<�ya<8ya<ya<�xa<�xa<�xa<�xa<�xa<�xa<$ya<=ya<zya<�ya<�ya<�ya<Uya<Bya<�xa<�xa<�xa<jxa<9xa<xa<!xa<xa<Sxa<�xa<�xa<ya<Qya<�  �  cya<�ya<�ya<za<Iza<Xza<Nza<Pza<0za<$za<za<za<'za<_za<�za<{a<z{a<|a<�|a<f}a<~a<�~a<za<4�a<��a<$�a<��a<��a<?�a<��a<�a<+�a<��a<�a<h�a<�a<��a<<�a<��a<��a<��a<]�a<�a<�a<��a<�a<��a<�a<z�a<ɍa<�a<a�a<��a<�a<Y�a<ޏa<n�a<�a<��a<z�a<b�a<�a<��a<��a<f�a<$�a<��a<��a<r�a<��a<Șa<�a<�a<&�a<P�a<|�a<��a<��a<H�a<��a<
�a<w�a<
�a<>�a<��a< �a<�a<8�a<c�a<9�a<)�a<�a<��a<��a<Y�a<:�a<1�a<H�a<Y�a<|�a<a<�a<~�a<Нa<9�a<��a<��a<��a<��a<�a< �a<��a<��a<p�a<�a<�a<��a<��a<w�a<t�a<v�a<��a<��a<��a<�a<�a<)�a<�a<��a<ٝa<��a<7�a<ߜa<_�a<�a<{�a<	�a<��a<k�a<F�a<�a<�a<�a<;�a<J�a<i�a<��a<��a<��a<o�a<>�a<�a<��a<7�a<�a<\�a<ؗa<i�a<��a<��a<F�a<�a<ԕa<��a<o�a<{�a<4�a<��a<͔a<Z�a<�a<~�a<Œa<#�a<`�a<��a<̏a<�a<.�a<{�a<�a<`�a<�a<��a<*�a<��a<��a<y�a<7�a<ىa<��a<�a<y�a<��a</�a<y�a<�a<�a<=�a<��a<�a<\�a<�a<z�a<$�a<Ԁa<��a<��a<�a<�a<�a<-a<�~a<e~a<�}a<+}a<z|a<�{a<J{a<�za<za<�ya<fya<!ya<�xa<�xa<�xa<ya<4ya<eya<{ya<�ya<�ya<wya<dya<Jya<�xa<�xa<�xa<+xa< xa<�wa<�wa<�wa<�wa<�wa<0xa<mxa<�xa<*ya<�  �  2ya<�ya<�ya<&za<Sza<hza<�za<mza<~za<dza<zza<�za<�za<�za<�za<�{a<�{a<|a<}a<�}a<]~a<�~a<�a<0�a<a<,�a<��a<߁a<	�a<^�a<��a<�a< �a<��a<��a<h�a</�a<Ѕa<��a<f�a<B�a<�a<�a<Ǌa<p�a<-�a<��a<2�a<��a<�a<V�a<��a<	�a<R�a<Ϗa<<�a<a<��a<�a<�a<��a<p�a<&�a<�a<��a<�a<��a<�a<F�a<p�a<��a<��a<��a<ܘa<�a< �a<1�a<��a<�a<<�a<Śa<�a<��a<�a<��a<֜a<�a<S�a<U�a<f�a<E�a<.�a<�a<ޜa<ʜa<��a<��a<��a<Ȝa<�a<(�a<��a<��a<�a<T�a<��a<מa<��a<�a<�a<؞a<��a<\�a<�a<͝a<��a<K�a<4�a<�a<�a<�a<:�a<b�a<�a<��a<ԝa<�a<�a<�a<�a<��a<l�a<��a<��a<0�a<ܛa<u�a<�a<��a<��a<��a<s�a<��a<��a<��a<��a<��a<��a<��a<��a<E�a<�a<��a<�a<��a<��a<��a<�a<��a<7�a<ŕa<��a<h�a<S�a<'�a<�a<�a<ʔa<��a<I�a<��a<x�a<�a<L�a<��a<ؐa<��a<]�a<��a<�a<F�a<��a<Z�a<��a<��a<6�a<��a<��a<^�a<�a<��a<�a<k�a<·a<�a<@�a<{�a<��a<�a<*�a<��a<�a<v�a<�a<��a<��a<8�a<!�a<�a<�a<}a</a<�~a<W~a<�}a<G}a<�|a<|a<�{a<{a<~za<%za<�ya<�ya<fya<Rya<cya<Wya<�ya<�ya<�ya<�ya<�ya<�ya<Nya<"ya<�xa<�xa<+xa<�wa<�wa<qwa<hwa<9wa<twa<�wa<�wa<)xa<sxa<�xa<�  �  ya<jya<�ya<za<Hza<�za<�za<�za<�za<�za<�za<�za<�za<4{a<z{a<�{a<O|a<�|a<R}a<~a<�~a<*a<�a<D�a<��a<'�a<l�a<��a<�a<�a<P�a<|�a<��a<�a<��a<#�a<��a<i�a<2�a<,�a<��a<�a<Љa<��a<��a<�a<��a<_�a<��a<$�a<��a<�a<Q�a<��a<.�a<��a<9�a<ݑa<��a<6�a<�a<Քa<\�a<�a<��a<!�a<��a<��a<�a<L�a<[�a<[�a<|�a<k�a<��a<��a<�a<%�a<q�a<ܙa<T�a<�a<Z�a<�a<[�a<��a<�a<=�a<f�a<��a<s�a<o�a<q�a<%�a<�a<�a<�a<�a<0�a<R�a<��a<ŝa<�a<t�a<��a<Ϟa<��a<�a<�a<�a<��a<s�a<�a<Ýa<|�a<"�a<ޜa<��a<��a<��a<��a<͜a<�a<;�a<r�a<��a<ϝa<��a<��a<؝a<ŝa<��a<0�a<��a<��a< �a<ћa<}�a<A�a<�a<�a<ۚa<Қa<Ța<��a<�a<ܚa<�a<��a<v�a<A�a<ԙa<f�a<�a<J�a<Ɨa<)�a<��a<#�a<˕a<��a<2�a<�a<�a<�a<Ôa<��a<��a<x�a<Y�a<�a<z�a<�a<i�a<��a<<�a<Y�a<��a<��a<P�a<��a<+�a<��a<K�a<�a<��a<c�a<ފa<�a<2�a<��a<�a<{�a<��a<�a<�a<)�a<k�a<��a<ɂa<�a<��a<�a<��a<X�a<�a<�a<�a<�a<�a<Za<0a<�~a<h~a<~a<u}a<�|a<�|a<�{a<V{a<�za<za<+za<�ya<�ya<�ya<�ya<�ya<�ya<�ya<�ya<�ya<�ya<qya<Mya<�xa<�xa<>xa<�wa<�wa<Awa<wa<�va<�va<�va<#wa<kwa<�wa</xa<�xa<�  �  �xa<:ya<�ya<za<dza<�za<�za<�za<�za<�za<{a<<{a<X{a<�{a<�{a<&|a<�|a<8}a<�}a<8~a<�~a<ua<�a<e�a<��a<�a<Z�a<s�a<��a<΁a<�a<�a<��a<̂a<%�a<ăa<C�a<5�a<ͅa<̆a<Ǉa<��a<��a<u�a<\�a<�a<ތa<d�a<��a<m�a<Վa<;�a<��a<�a<��a<��a<��a<0�a<�a<��a<@�a<�a<��a<F�a<��a<J�a<��a<ؗa< �a<�a<�a<'�a<$�a<�a<O�a<;�a<��a<��a<�a<��a<�a<��a<�a<��a<�a<��a<�a<F�a<��a<��a<��a<��a<��a<��a<~�a<k�a<S�a<l�a<w�a<��a<�a<�a<S�a<��a<՞a<��a<�a<�a<�a<Ҟa<w�a<8�a<ѝa<��a<�a<Ɯa<��a<E�a<V�a<*�a<j�a<}�a<��a<�a</�a<z�a<��a<�a<�a<��a<֝a<��a<{�a<�a<Ĝa<r�a<1�a<ۛa<��a<p�a<8�a<9�a<;�a<$�a<�a<�a<'�a<�a<Ԛa<��a<-�a<Ùa<%�a<��a<�a<��a<Öa<f�a<ڕa<]�a<!�a<��a<͔a<{�a<��a<��a<w�a<l�a<P�a<5�a<�a<��a<�a<��a<�a<W�a<��a<�a<W�a<��a<�a<��a<	�a<��a<=�a<ދa<��a<!�a<��a<1�a<��a< �a<T�a<��a<��a<̅a<��a<�a<�a<��a<��a<5�a<��a<N�a<$�a<�a<�a<�a<za<Va<Ka<a<�~a<�~a<~a<�}a<+}a<�|a<+|a<�{a<C{a<�za<�za<?za<#za<za<�ya<�ya<�ya<za<�ya<�ya<�ya<oya<4ya<�xa<nxa<�wa<�wa<7wa<�va<�va<yva<�va<�va<�va<wa<jwa< xa<Uxa<�  �  �xa<?ya<�ya<za<mza<�za<�za<�za<.{a<F{a<i{a<t{a<�{a<�{a</|a<�|a<�|a<s}a<~a<�~a<a<�a<�a<[�a<Ҁa<��a<O�a<k�a<��a<��a<��a<�a<�a<a�a<тa<i�a<��a<��a<��a<��a<z�a<w�a<u�a<{�a<>�a<&�a<ьa<e�a<�a<��a<�a<��a<�a<W�a<�a<e�a<�a<��a<�a<�a<��a<3�a<ʕa<`�a<ǖa<6�a<��a<��a<��a<��a<�a<�a<ߗa<ߗa<җa<�a<&�a<d�a<��a<3�a<řa<K�a<�a<z�a<	�a<��a<�a<_�a<~�a<��a<Нa<ڝa<֝a<ѝa<Ýa<��a<ʝa<��a<�a<�a<#�a<p�a<��a<ўa<�a<�a<�a<�a<��a<��a<}�a<�a<��a<:�a<ߜa<��a<9�a<��a<�a<ߛa<��a<.�a<p�a<��a<��a<S�a<��a<ɝa<�a<��a<ԝa<ǝa<��a<]�a<�a<̜a<i�a<2�a<��a<��a<��a<x�a<v�a<z�a<g�a<\�a<7�a<	�a<ʚa<��a<�a<��a<�a<}�a<җa<,�a<��a<��a<p�a<	�a<Ɣa<r�a<T�a<R�a<K�a<H�a<M�a<P�a<V�a<�a<��a<��a<�a<��a<)�a<��a<�a<U�a<��a<�a<o�a<ߍa<y�a<�a<��a<$�a<��a<L�a<يa<:�a<��a<�a<7�a<��a<��a<��a<��a<΃a<��a<�a<\�a<րa<Q�a<�a<�a<�a<ja<Za<Ra<Fa<Ca<�~a<�~a<�~a<(~a<�}a<d}a<�|a<x|a<|a<�{a<B{a<�za<�za<�za<Mza<Sza<@za<5za<za<za<�ya<�ya<tya<ya<�xa<Gxa<�wa<Zwa<�va<�va<_va<.va<7va<=va<zva<�va<6wa<�wa<$xa<�  �  �xa<ya<�ya< za<pza<�za<{a<{a<^{a<^{a<�{a<�{a<�{a<)|a<c|a<�|a< }a<�}a<%~a<�~a<9a<�a<J�a<o�a<؀a<�a<$�a<E�a<e�a<��a<��a<Ɓa<ׁa<@�a<��a<&�a<�a<v�a<v�a<\�a<I�a<o�a<K�a<J�a<(�a<�a<Ҍa<��a<6�a<��a<N�a<��a<;�a<��a<�a<��a<$�a<Œa<U�a<�a<��a<n�a<�a<{�a<#�a<>�a<��a<��a<̗a<̗a<�a<��a<��a<��a<��a<ڗa<�a<1�a<��a<�a<��a<�a<ǚa<`�a<�a<o�a<ݜa<c�a<��a<�a<�a<��a<�a<�a<��a<۝a<��a<��a< �a<7�a<^�a<��a<��a<�a<�a<E�a<@�a<�a<�a<��a<N�a<�a<��a<�a<��a<N�a<��a<��a<��a<a<a<�a<L�a<w�a<��a<&�a<v�a<��a<ܝa< �a<�a<�a<��a<��a<)�a<��a<��a<_�a<5�a<��a<�a<��a<��a<��a<��a<��a<K�a<]�a<ޚa<��a<�a<��a<��a<]�a<��a<��a<s�a<��a<N�a<ܔa<��a<d�a<�a<$�a<�a<�a<E�a<&�a<&�a< �a<�a<��a<q�a<ߒa<H�a<Бa<�a<��a<ȏa<7�a<��a<�a<��a<�a<όa<:�a<��a<j�a<�a<��a<��a<�a<)�a<U�a<g�a<��a<��a<��a<˂a<Ёa<Q�a<��a<�a<�a<ja<ha<5a<@a<8a<a<a<�~a<�~a<�~a<�~a<�}a<�}a<}a<�|a<7|a<�{a<t{a<{a<�za<�za<�za<�za<Uza<jza<4za<>za<za<�ya<iya<�xa<�xa<xa<�wa<%wa<�va<mva<va<va<�ua< va<>va<�va<wa<kwa<xa<�  �  �xa<ya<�ya<za<fza<�za<�za<9{a<h{a<�{a<�{a<�{a<|a<J|a<�|a<�|a<r}a<�}a<V~a<�~a<Qa<�a<�a<c�a<ƀa<�a<<�a<E�a<W�a<J�a<d�a<��a<ȁa<�a<U�a<�a<��a<n�a<4�a<.�a<"�a<A�a<H�a<K�a<O�a<�a<ڌa<��a<1�a<؎a<R�a<׏a<E�a<ϐa<F�a<בa<h�a<�a<��a<,�a<ޔa<t�a<�a<��a<�a<F�a<��a<їa<ӗa<Ηa<��a<��a<��a<n�a<��a<��a<��a<�a<f�a<�a<X�a<��a<��a<I�a<�a<��a<��a<L�a<��a<ҝa<��a<�a<�a<'�a<�a<.�a<�a<?�a<G�a<l�a<��a<��a<�a<�a<.�a<&�a<%�a<�a<��a<��a<M�a<�a<l�a<�a<��a< �a<�a<��a<s�a<n�a<��a<Λa<�a<`�a<��a<$�a<s�a<ɝa<�a<��a<�a<ߝa<ȝa<��a<Y�a<�a<ߜa<��a<W�a<?�a< �a<��a<ۛa<̛a<��a<��a<d�a</�a<Қa<��a<'�a<��a<��a<O�a<��a<ږa<1�a<��a<!�a<��a<>�a<
�a<�a<�a<�a<�a<�a<#�a<'�a<'�a<�a<��a<H�a<ڒa<o�a<ԑa<B�a<��a<
�a<h�a<�a<Z�a<̍a<a�a<یa<|�a<�a<��a<��a<b�a<��a<�a<M�a<\�a<i�a<k�a<W�a<r�a<��a<ˁa<��a<U�a<�a<�a<aa<"a<a<a<!a<$a<)a<a<�~a<�~a<Q~a<�}a<�}a<-}a<�|a<W|a<|a<�{a<\{a<{a<�za<�za<�za<�za<oza<Zza< za<�ya<�ya<zya<ya<�xa<xa<�wa<	wa<�va<?va<
va<�ua<�ua<�ua<$va<mva<�va<Twa<�wa<�  �  �xa<�xa<uya<�ya<sza<�za<{a<^{a<Z{a<�{a<�{a<�{a<|a<:|a<�|a<�|a<q}a<�}a<f~a<�~a<Ra<�a<)�a<��a<ʀa<�a<�a< �a<N�a<=�a<��a<y�a<��a<�a<o�a<-�a<q�a<j�a<�a<D�a<5�a<(�a<@�a<'�a<)�a<�a< �a<��a<V�a<�a<6�a<�a<2�a<ѐa<H�a<ʑa<]�a<�a<��a<�a<�a<V�a<�a<��a<�a<z�a<��a<��a<��a<��a<��a<��a<��a<W�a<��a<Z�a<�a<�a<5�a<՘a<K�a<�a<��a<>�a<Ǜa<Q�a<؜a<L�a<ǝa<ٝa<�a<'�a<�a<C�a<��a<3�a<�a<:�a<:�a<q�a<��a<��a<�a<��a<S�a<F�a<F�a<'�a<֞a<��a<"�a<�a<P�a<��a<��a<�a<қa<|�a<��a<f�a<��a<��a<�a<y�a<��a<"�a<H�a<��a<Νa<�a<�a<��a<�a<��a<{�a<�a<ʜa<��a<F�a<A�a<�a<��a<��a<ݛa<��a<��a<��a<<�a<�a<��a<�a<t�a<Ҙa<G�a<v�a<��a<'�a<��a<��a<��a<��a<�a<�a<Γa<�a<�a<��a<�a<�a<�a<ٓa<Ǔa<M�a<��a<��a<��a<p�a<��a<�a<j�a<Ԏa<N�a<Ǎa<h�a<ǌa<��a<�a<��a<"�a<`�a<�a<��a<*�a<3�a<Z�a<Z�a<g�a<��a<n�a<Ła<рa<��a<�a<ga<Pa<a<>a<a<a<a<�~a<�~a<�~a<�~a<X~a< ~a<�}a<(}a<�|a<<|a<|a<�{a<W{a<{a<�za<�za<�za<�za<`za<za<@za<za<�ya<Vya<�xa<kxa<xa<xwa<wa<�va<-va<�ua<�ua<va<�ua<va<]va<�va<mwa<�wa<�  �  �xa<ya<�ya<za<fza<�za<�za<9{a<h{a<�{a<�{a<�{a<|a<J|a<�|a<�|a<r}a<�}a<V~a<�~a<Qa<�a<�a<c�a<ƀa<�a<<�a<E�a<W�a<J�a<d�a<��a<ȁa<�a<U�a<�a<��a<n�a<4�a<.�a<"�a<A�a<H�a<K�a<O�a<�a<ڌa<��a<1�a<؎a<R�a<׏a<E�a<ϐa<F�a<בa<h�a<�a<��a<,�a<ޔa<t�a<�a<��a<�a<F�a<��a<їa<ӗa<Ηa<��a<��a<��a<n�a<��a<��a<��a<�a<f�a<�a<X�a<��a<��a<I�a<�a<��a<��a<L�a<��a<ҝa<��a<�a<�a<'�a<�a<.�a<�a<?�a<G�a<l�a<��a<��a<�a<�a<.�a<&�a<%�a<�a<��a<��a<M�a<�a<l�a<�a<��a< �a<�a<��a<s�a<n�a<��a<Λa<�a<`�a<��a<$�a<s�a<ɝa<�a<��a<�a<ߝa<ȝa<��a<Y�a<�a<ߜa<��a<W�a<?�a< �a<��a<ۛa<̛a<��a<��a<d�a</�a<Қa<��a<'�a<��a<��a<O�a<��a<ږa<1�a<��a<!�a<��a<>�a<
�a<�a<�a<�a<�a<�a<#�a<'�a<'�a<�a<��a<H�a<ڒa<o�a<ԑa<B�a<��a<
�a<h�a<�a<Z�a<̍a<a�a<یa<|�a<�a<��a<��a<b�a<��a<�a<M�a<\�a<i�a<k�a<W�a<r�a<��a<ˁa<��a<U�a<�a<�a<aa<"a<a<a<!a<$a<)a<a<�~a<�~a<Q~a<�}a<�}a<-}a<�|a<W|a<|a<�{a<\{a<{a<�za<�za<�za<�za<oza<Zza< za<�ya<�ya<zya<ya<�xa<xa<�wa<	wa<�va<?va<
va<�ua<�ua<�ua<$va<mva<�va<Twa<�wa<�  �  �xa<ya<�ya< za<pza<�za<{a<{a<^{a<^{a<�{a<�{a<�{a<)|a<c|a<�|a< }a<�}a<%~a<�~a<9a<�a<J�a<o�a<؀a<�a<$�a<E�a<e�a<��a<��a<Ɓa<ׁa<@�a<��a<&�a<�a<v�a<v�a<\�a<I�a<o�a<K�a<J�a<(�a<�a<Ҍa<��a<6�a<��a<N�a<��a<;�a<��a<�a<��a<$�a<Œa<U�a<�a<��a<n�a<�a<{�a<#�a<>�a<��a<��a<̗a<̗a<�a<��a<��a<��a<��a<ڗa<�a<1�a<��a<�a<��a<�a<ǚa<`�a<�a<o�a<ݜa<c�a<��a<�a<�a<��a<�a<�a<��a<۝a<��a<��a< �a<7�a<^�a<��a<��a<�a<�a<E�a<@�a<�a<�a<��a<N�a<�a<��a<�a<��a<N�a<��a<��a<��a<a<a<�a<L�a<w�a<��a<&�a<v�a<��a<ܝa< �a<�a<�a<��a<��a<)�a<��a<��a<_�a<5�a<��a<�a<��a<��a<��a<��a<��a<K�a<]�a<ޚa<��a<�a<��a<��a<]�a<��a<��a<s�a<��a<N�a<ܔa<��a<d�a<�a<$�a<�a<�a<E�a<&�a<&�a< �a<�a<��a<q�a<ߒa<H�a<Бa<�a<��a<ȏa<7�a<��a<�a<��a<�a<όa<:�a<��a<j�a<�a<��a<��a<�a<)�a<U�a<g�a<��a<��a<��a<˂a<Ёa<Q�a<��a<�a<�a<ja<ha<5a<@a<8a<a<a<�~a<�~a<�~a<�~a<�}a<�}a<}a<�|a<7|a<�{a<t{a<{a<�za<�za<�za<�za<Uza<jza<4za<>za<za<�ya<iya<�xa<�xa<xa<�wa<%wa<�va<mva<va<va<�ua< va<>va<�va<wa<kwa<xa<�  �  �xa<?ya<�ya<za<mza<�za<�za<�za<.{a<F{a<i{a<t{a<�{a<�{a</|a<�|a<�|a<s}a<~a<�~a<a<�a<�a<[�a<Ҁa<��a<O�a<k�a<��a<��a<��a<�a<�a<a�a<тa<i�a<��a<��a<��a<��a<z�a<w�a<u�a<{�a<>�a<&�a<ьa<e�a<�a<��a<�a<��a<�a<W�a<�a<e�a<�a<��a<�a<�a<��a<3�a<ʕa<`�a<ǖa<6�a<��a<��a<��a<��a<�a<�a<ߗa<ߗa<җa<�a<&�a<d�a<��a<3�a<řa<K�a<�a<z�a<	�a<��a<�a<_�a<~�a<��a<Нa<ڝa<֝a<ѝa<Ýa<��a<ʝa<��a<�a<�a<#�a<p�a<��a<ўa<�a<�a<�a<�a<��a<��a<}�a<�a<��a<:�a<ߜa<��a<9�a<��a<�a<ߛa<��a<.�a<p�a<��a<��a<S�a<��a<ɝa<�a<��a<ԝa<ǝa<��a<]�a<�a<̜a<i�a<2�a<��a<��a<��a<x�a<v�a<z�a<g�a<\�a<7�a<	�a<ʚa<��a<�a<��a<�a<}�a<җa<,�a<��a<��a<p�a<	�a<Ɣa<r�a<T�a<R�a<K�a<H�a<M�a<P�a<V�a<�a<��a<��a<�a<��a<)�a<��a<�a<U�a<��a<�a<o�a<ߍa<y�a<�a<��a<$�a<��a<L�a<يa<:�a<��a<�a<7�a<��a<��a<��a<��a<΃a<��a<�a<\�a<րa<Q�a<�a<�a<�a<ja<Za<Ra<Fa<Ca<�~a<�~a<�~a<(~a<�}a<d}a<�|a<x|a<|a<�{a<B{a<�za<�za<�za<Mza<Sza<@za<5za<za<za<�ya<�ya<tya<ya<�xa<Gxa<�wa<Zwa<�va<�va<_va<.va<7va<=va<zva<�va<6wa<�wa<$xa<�  �  �xa<:ya<�ya<za<dza<�za<�za<�za<�za<�za<{a<<{a<X{a<�{a<�{a<&|a<�|a<8}a<�}a<8~a<�~a<ua<�a<e�a<��a<�a<Z�a<s�a<��a<΁a<�a<�a<��a<̂a<%�a<ăa<C�a<5�a<ͅa<̆a<Ǉa<��a<��a<u�a<\�a<�a<ތa<d�a<��a<m�a<Վa<;�a<��a<�a<��a<��a<��a<0�a<�a<��a<@�a<�a<��a<F�a<��a<J�a<��a<ؗa< �a<�a<�a<'�a<$�a<�a<O�a<;�a<��a<��a<�a<��a<�a<��a<�a<��a<�a<��a<�a<F�a<��a<��a<��a<��a<��a<��a<~�a<k�a<S�a<l�a<w�a<��a<�a<�a<S�a<��a<՞a<��a<�a<�a<�a<Ҟa<w�a<8�a<ѝa<��a<�a<Ɯa<��a<E�a<V�a<*�a<j�a<}�a<��a<�a</�a<z�a<��a<�a<�a<��a<֝a<��a<{�a<�a<Ĝa<r�a<1�a<ۛa<��a<p�a<8�a<9�a<;�a<$�a<�a<�a<'�a<�a<Ԛa<��a<-�a<Ùa<%�a<��a<�a<��a<Öa<f�a<ڕa<]�a<!�a<��a<͔a<{�a<��a<��a<w�a<l�a<P�a<5�a<�a<��a<�a<��a<�a<W�a<��a<�a<W�a<��a<�a<��a<	�a<��a<=�a<ދa<��a<!�a<��a<1�a<��a< �a<T�a<��a<��a<̅a<��a<�a<�a<��a<��a<5�a<��a<N�a<$�a<�a<�a<�a<za<Va<Ka<a<�~a<�~a<~a<�}a<+}a<�|a<+|a<�{a<C{a<�za<�za<?za<#za<za<�ya<�ya<�ya<za<�ya<�ya<�ya<oya<4ya<�xa<nxa<�wa<�wa<7wa<�va<�va<yva<�va<�va<�va<wa<jwa< xa<Uxa<�  �  ya<jya<�ya<za<Hza<�za<�za<�za<�za<�za<�za<�za<�za<4{a<z{a<�{a<O|a<�|a<R}a<~a<�~a<*a<�a<D�a<��a<'�a<l�a<��a<�a<�a<P�a<|�a<��a<�a<��a<#�a<��a<i�a<2�a<,�a<��a<�a<Љa<��a<��a<�a<��a<_�a<��a<$�a<��a<�a<Q�a<��a<.�a<��a<9�a<ݑa<��a<6�a<�a<Քa<\�a<�a<��a<!�a<��a<��a<�a<L�a<[�a<[�a<|�a<k�a<��a<��a<�a<%�a<q�a<ܙa<T�a<�a<Z�a<�a<[�a<��a<�a<=�a<f�a<��a<s�a<o�a<q�a<%�a<�a<�a<�a<�a<0�a<R�a<��a<ŝa<�a<t�a<��a<Ϟa<��a<�a<�a<�a<��a<s�a<�a<Ýa<|�a<"�a<ޜa<��a<��a<��a<��a<͜a<�a<;�a<r�a<��a<ϝa<��a<��a<؝a<ŝa<��a<0�a<��a<��a< �a<ћa<}�a<A�a<�a<�a<ۚa<Қa<Ța<��a<�a<ܚa<�a<��a<v�a<A�a<ԙa<f�a<�a<J�a<Ɨa<)�a<��a<#�a<˕a<��a<2�a<�a<�a<�a<Ôa<��a<��a<x�a<Y�a<�a<z�a<�a<i�a<��a<<�a<Y�a<��a<��a<P�a<��a<+�a<��a<K�a<�a<��a<c�a<ފa<�a<2�a<��a<�a<{�a<��a<�a<�a<)�a<k�a<��a<ɂa<�a<��a<�a<��a<X�a<�a<�a<�a<�a<�a<Za<0a<�~a<h~a<~a<u}a<�|a<�|a<�{a<V{a<�za<za<+za<�ya<�ya<�ya<�ya<�ya<�ya<�ya<�ya<�ya<�ya<qya<Mya<�xa<�xa<>xa<�wa<�wa<Awa<wa<�va<�va<�va<#wa<kwa<�wa</xa<�xa<�  �  2ya<�ya<�ya<&za<Sza<hza<�za<mza<~za<dza<zza<�za<�za<�za<�za<�{a<�{a<|a<}a<�}a<]~a<�~a<�a<0�a<a<,�a<��a<߁a<	�a<^�a<��a<�a< �a<��a<��a<h�a</�a<Ѕa<��a<f�a<B�a<�a<�a<Ǌa<p�a<-�a<��a<2�a<��a<�a<V�a<��a<	�a<R�a<Ϗa<<�a<a<��a<�a<�a<��a<p�a<&�a<�a<��a<�a<��a<�a<F�a<p�a<��a<��a<��a<ܘa<�a< �a<1�a<��a<�a<<�a<Śa<�a<��a<�a<��a<֜a<�a<S�a<U�a<f�a<E�a<.�a<�a<ޜa<ʜa<��a<��a<��a<Ȝa<�a<(�a<��a<��a<�a<T�a<��a<מa<��a<�a<�a<؞a<��a<\�a<�a<͝a<��a<K�a<4�a<�a<�a<�a<:�a<b�a<�a<��a<ԝa<�a<�a<�a<�a<��a<l�a<��a<��a<0�a<ܛa<u�a<�a<��a<��a<��a<s�a<��a<��a<��a<��a<��a<��a<��a<��a<E�a<�a<��a<�a<��a<��a<��a<�a<��a<7�a<ŕa<��a<h�a<S�a<'�a<�a<�a<ʔa<��a<I�a<��a<x�a<�a<L�a<��a<ؐa<��a<]�a<��a<�a<F�a<��a<Z�a<��a<��a<6�a<��a<��a<^�a<�a<��a<�a<k�a<·a<�a<@�a<{�a<��a<�a<*�a<��a<�a<v�a<�a<��a<��a<8�a<!�a<�a<�a<}a</a<�~a<W~a<�}a<G}a<�|a<|a<�{a<{a<~za<%za<�ya<�ya<fya<Rya<cya<Wya<�ya<�ya<�ya<�ya<�ya<�ya<Nya<"ya<�xa<�xa<+xa<�wa<�wa<qwa<hwa<9wa<twa<�wa<�wa<)xa<sxa<�xa<�  �  cya<�ya<�ya<za<Iza<Xza<Nza<Pza<0za<$za<za<za<'za<_za<�za<{a<z{a<|a<�|a<f}a<~a<�~a<za<4�a<��a<$�a<��a<��a<?�a<��a<�a<+�a<��a<�a<h�a<�a<��a<<�a<��a<��a<��a<]�a<�a<�a<��a<�a<��a<�a<z�a<ɍa<�a<a�a<��a<�a<Y�a<ޏa<n�a<�a<��a<z�a<b�a<�a<��a<��a<f�a<$�a<��a<��a<r�a<��a<Șa<�a<�a<&�a<P�a<|�a<��a<��a<H�a<��a<
�a<w�a<
�a<>�a<��a< �a<�a<8�a<c�a<9�a<)�a<�a<��a<��a<Y�a<:�a<1�a<H�a<Y�a<|�a<a<�a<~�a<Нa<9�a<��a<��a<��a<��a<�a< �a<��a<��a<p�a<�a<�a<��a<��a<w�a<t�a<v�a<��a<��a<��a<�a<�a<)�a<�a<��a<ٝa<��a<7�a<ߜa<_�a<�a<{�a<	�a<��a<k�a<F�a<�a<�a<�a<;�a<J�a<i�a<��a<��a<��a<o�a<>�a<�a<��a<7�a<�a<\�a<ؗa<i�a<��a<��a<F�a<�a<ԕa<��a<o�a<{�a<4�a<��a<͔a<Z�a<�a<~�a<Œa<#�a<`�a<��a<̏a<�a<.�a<{�a<�a<`�a<�a<��a<*�a<��a<��a<y�a<7�a<ىa<��a<�a<y�a<��a</�a<y�a<�a<�a<=�a<��a<�a<\�a<�a<z�a<$�a<Ԁa<��a<��a<�a<�a<�a<-a<�~a<e~a<�}a<+}a<z|a<�{a<J{a<�za<za<�ya<fya<!ya<�xa<�xa<�xa<ya<4ya<eya<{ya<�ya<�ya<wya<dya<Jya<�xa<�xa<�xa<+xa< xa<�wa<�wa<�wa<�wa<�wa<0xa<mxa<�xa<*ya<�  �  �ya<�ya<za<3za<@za<Eza<za<za<�ya<�ya<�ya<�ya<�ya<�ya<Xza<�za<D{a<�{a<d|a<;}a<�}a<�~a<Oa<�a<��a<I�a<��a<+�a<��a<Ԃa<&�a<v�a<�a<D�a<��a<E�a<ׅa<��a<R�a<�a<͈a<��a<^�a<�a<��a<�a<��a<��a<8�a<��a<ɍa<�a<0�a<��a<��a<x�a<�a<��a<��a<�a<�a<�a<��a<��a<P�a< �a<��a<&�a<r�a<՘a<�a<3�a<]�a<��a<��a<̙a<�a<D�a<��a<�a<U�a<��a<$�a<��a<֜a<�a<B�a<7�a<B�a<�a<�a<��a<��a<@�a<��a<�a<��a<�a<�a<6�a<��a<��a<F�a<��a<��a<D�a<��a<�a<
�a<!�a<�a<�a<̞a<��a<h�a<L�a<�a<ڝa<۝a<��a<؝a<��a<��a<�a<*�a<Q�a<?�a<3�a<�a<Нa<��a<�a<��a<�a<��a<�a<��a<l�a<��a<�a<��a<Йa<��a<ڙa<�a<#�a<S�a<a�a<��a<n�a<c�a<�a<ݙa<��a<�a<��a<#�a<ȗa<R�a<�a<��a<T�a<-�a<�a<Εa<��a<i�a<:�a<͔a<��a<�a<b�a<��a<�a<�a<K�a<��a<��a<��a< �a<��a<��a<|�a<K�a<Ċa<��a<s�a<7�a<��a<Éa<q�a<�a<��a<��a<p�a<��a< �a<M�a<��a<�a<C�a<��a<2�a<Ёa<��a< �a<߀a<��a<_�a<�a<�a<Wa<�~a<D~a<�}a<�|a<9|a<�{a<�za<2za<�ya<8ya<ya<�xa<�xa<�xa<�xa<�xa<�xa<$ya<=ya<zya<�ya<�ya<�ya<Uya<Bya<�xa<�xa<�xa<jxa<9xa<xa<!xa<xa<Sxa<�xa<�xa<ya<Qya<�  �  �ya<�ya<za<?za<5za</za<za<�ya<�ya<�ya<�ya<wya<~ya<�ya<�ya<Hza<�za<v{a<'|a<�|a<�}a<~~a<Ua<�a<��a<H�a<��a<H�a<��a<�a<o�a<փa< �a<��a<�a<��a<M�a<ӆa<��a<W�a<�a<Ɖa<w�a<�a<��a<6�a<�a<��a<%�a<]�a<��a<Ía<�a<F�a<��a<�a<��a<G�a<	�a<�a<ƒa<��a<��a<k�a<N�a<�a<��a<�a<~�a<�a<4�a<t�a<��a<ؙa<�a<?�a<_�a<��a<�a<A�a<��a<�a<b�a<��a<�a<�a<9�a<I�a<"�a<�a<̜a<��a<<�a<��a<ƛa<��a<q�a<��a<��a<̛a<"�a<��a<�a<Y�a<Нa<@�a<��a<Ҟa<�a<�a<&�a<�a<�a<�a<��a<��a<U�a<P�a<.�a<3�a<&�a<-�a<T�a<^�a<n�a<`�a<\�a</�a<�a<ŝa<n�a<�a<{�a<�a<[�a<�a<l�a<�a<��a<��a<X�a<`�a<y�a<��a<ęa<��a</�a<g�a<h�a<w�a<a�a<�a<��a<��a<K�a<�a<��a< �a<��a<W�a<��a<ʖa<k�a<N�a<�a<ߕa<��a<R�a<�a<p�a<�a<F�a<��a<ϑa<��a<�a</�a<_�a<��a<��a<&�a<��a<!�a<͊a<��a<d�a<5�a<�a<�a<��a<T�a<�a<��a<�a<��a<�a<B�a<��a<�a<,�a<��a<�a<��a<9�a<��a<��a<'�a<ۀa<��a<.�a<�a<Na<�~a<$~a<�}a<�|a<|a<S{a<�za<za<hya<�xa<�xa<_xa<Cxa<Lxa<jxa<�xa<�xa<�xa<9ya<kya<uya<�ya<{ya<oya<Pya<4ya<ya<�xa<�xa<{xa<�xa<txa<�xa<�xa<�xa<ya<Rya<�ya<�  �  �ya<:za<6za<Cza<'za<	za<�ya<�ya<�ya<]ya<bya<3ya<Fya<�ya<�ya</za<�za<B{a<�{a<�|a<�}a<R~a<'a<�a<��a<G�a<��a<t�a<ła<K�a<��a<�a<Z�a<Єa<W�a<Ӆa<}�a<�a<Ӈa<q�a<D�a<�a<��a<e�a<��a<:�a<s�a<ƌa<��a<E�a<p�a<��a<�a<�a<��a<�a<u�a<;�a<Đa<őa<��a<~�a<z�a<A�a<�a<֖a<��a<�a<ݘa<	�a<S�a<��a<��a<�a<�a<h�a<��a<�a<-�a<x�a<�a<�a<��a<ɜa<�a<T�a<8�a<A�a<�a<�a<��a<|�a<
�a<ӛa<��a<I�a<a�a<I�a<n�a<��a<ޛa<c�a<��a<I�a<��a<�a<x�a<Ǟa<!�a<4�a<u�a<0�a<;�a<�a<�a<��a<��a<��a<a�a<h�a<V�a<j�a<}�a<x�a<��a<w�a<��a<Y�a<�a<��a<H�a<ڜa<P�a<ޛa<(�a<Ěa<(�a<șa<��a<>�a<@�a<�a<E�a<u�a<��a<�a<�a<9�a<H�a<n�a<`�a<_�a<&�a<��a<��a<��a<��a<:�a<ޗa<��a<0�a<��a<��a<��a<2�a<�a<��a<f�a<A�a<{�a<�a<:�a<�a<��a<ېa<�a<��a<6�a<<�a<��a<�a<f�a<�a<��a<u�a<2�a<�a<��a<��a<��a<H�a<�a<��a<e�a<��a<�a<{�a<��a<%�a<`�a<߃a<F�a<ւa<_�a<�a<��a<=�a<�a<��a<U�a<�a<Na<�~a<
~a<g}a<�|a<|a<!{a<{za<�ya<#ya<�xa<gxa<6xa<xa<xa<Fxa<Rxa<�xa<�xa<ya<Cya<jya<�ya<�ya<�ya<fya<bya<$ya< ya<�xa<�xa<�xa<�xa<�xa<�xa<ya<Cya<lya<�ya<�  �  �ya<za<"za<7za<>za<+za<�ya<�ya<wya<Fya<%ya<ya<)ya<-ya<vya<�ya<~za<{a<�{a<�|a<u}a<Q~a<%a<�a<��a<H�a<؁a<Y�a<�a<N�a<��a< �a<��a<�a<��a<�a<��a<V�a<�a<��a<P�a<	�a<��a<.�a<��a<"�a<��a<،a<�a<*�a<6�a<l�a<��a<��a<H�a<��a<2�a<�a<��a<�a<k�a<K�a<V�a<D�a<%�a<��a<��a<�a<��a<�a<x�a<��a<��a<�a<h�a<��a<ݚa<�a<`�a<��a<��a<Y�a<��a<�a<�a</�a<>�a<E�a<0�a<�a<��a<M�a<�a<��a<[�a<@�a<�a<�a<�a<|�a<˛a<#�a<��a<�a<��a<�a<��a<ߞa<�a<$�a<I�a<L�a<O�a<#�a<�a<�a<מa<��a<��a<��a<��a<��a<��a<��a<��a<��a<x�a<E�a<�a<Νa<j�a<לa<L�a<��a<�a<��a<�a<��a<9�a<�a<�a<
�a<�a<B�a<p�a<��a<�a<7�a<p�a<{�a<a�a<?�a<�a<�a<��a<2�a<͘a<z�a<�a<��a<u�a<�a<�a<��a<n�a<�a<��a<r�a<
�a<w�a<�a<Z�a<��a<��a<��a<��a<׎a<��a<5�a<j�a<��a<#�a<Ċa<��a<.�a<�a<ىa<׉a<��a<��a<k�a<�a<��a<0�a<��a<*�a<��a<�a<5�a<��a<�a<��a<�a<��a<4�a<Ɂa<x�a<�a<ƀa<I�a<�a<Ta<�~a<2~a<g}a<�|a<�{a<�za<Lza<�ya<ya<�xa<$xa<�wa<�wa<�wa<xa<7xa<sxa<�xa<ya<]ya<�ya<�ya<�ya<�ya<�ya<vya<Bya<,ya<ya<�xa<�xa<�xa<�xa<ya<=ya<fya<�ya<�ya<�  �  �{a<�{a<�{a<�{a<�{a<�{a<|{a<�{a<b{a<u{a<@{a<T{a<`{a<�{a<|a< |a<�|a<6}a<�}a<�~a<Ja<�a<��a<u�a<�a<͂a<i�a<ڃa<_�a<��a<F�a<��a<�a<��a<�a<m�a<��a<ψa<2�a<#�a<{�a<=�a<��a<p�a<)�a<_�a<͍a<�a<O�a<��a<�a<J�a<^�a<�a<�a<��a<T�a<��a<��a<-�a<'�a<�a<��a<k�a<)�a<��a<��a<`�a<��a<%�a<j�a<��a<"�a<�a<��a<��a<Λa<�a<s�a<Мa<��a<��a<{�a<��a<!�a<K�a<e�a<@�a<6�a<��a<�a<��a<��a<V�a<�a<�a<ڜa<,�a<�a<9�a<��a<˝a<[�a<��a<��a<5�a<��a<�a<'�a<t�a<\�a<s�a<;�a<3�a<@�a<�a<�a<��a<��a<��a<ڟa<��a<ǟa<��a<��a<şa<��a<��a<2�a<ߞa<{�a<��a<��a<&�a<՜a<8�a<ߛa<z�a<+�a<1�a<ʚa<�a<Ԛa<��a<*�a<5�a<O�a<[�a<��a<��a<��a<u�a<1�a<��a<t�a<e�a<ޙa<��a<A�a<˘a<|�a<1�a<�a<��a<��a<�a<ؖa<��a<�a<ѕa<�a<l�a<��a<ڒa<,�a<X�a<��a<��a<�a<=�a<̍a<U�a<��a<��a<��a<�a<��a<e�a<�a<׊a<��a<H�a<%�a<|�a<�a<o�a<��a<j�a<��a<+�a<q�a<߄a<a�a<
�a<��a<1�a<�a<]�a<8�a<ȁa<\�a<�a<5�a<�a<�~a<Q~a<�}a<}a<m|a<�{a<_{a<�za<�za<Qza<"za<2za<!za<oza<nza<�za<�za<�za<{a<{a<K{a<{a<{a<�za<�za<�za<�za<�za<jza<oza<zza<�za<�za<{a<${a</{a<�  �  r{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<i{a<U{a<G{a<U{a<s{a<�{a<�{a<5|a<�|a<G}a<�}a<�~a<Ra<�a<܀a<��a<"�a<��a<?�a<��a<D�a<��a<$�a<��a<��a<e�a<��a<��a<�a<��a<B�a<��a<��a<O�a<Ƌa<Y�a<�a<Y�a<׍a<2�a<~�a<��a<�a<:�a<w�a<֏a<3�a<��a<%�a<Бa<��a<G�a<�a<ߔa<��a<��a<Y�a<�a<��a<�a<��a<�a<m�a<��a<�a<!�a<b�a<��a<��a<0�a<b�a<��a<�a<Y�a<��a<�a<��a<(�a<3�a<G�a<C�a<,�a<��a<��a<y�a<T�a<%�a<�a<�a<�a<�a<T�a<��a<ڝa<=�a<��a<�a<m�a<��a<��a<�a<9�a<B�a<M�a<^�a<6�a<%�a<��a<ݟa<ɟa<��a<��a<��a<��a<��a<��a<��a<��a<u�a<X�a< �a<�a<��a<3�a<��a<,�a<��a<?�a<��a<��a<2�a<��a<ߚa<�a<�a<��a<�a<<�a<e�a<��a<��a<��a<c�a<K�a<	�a<�a<��a<C�a<�a<��a<"�a<��a<��a<3�a<�a<��a<s�a<#�a<�a<i�a< �a<��a<��a<v�a<ɓa<
�a<7�a<S�a<��a<Ïa<�a<Z�a<��a<&�a<��a<t�a<�a<�a<��a<r�a<E�a<�a<��a<D�a<��a<d�a<܈a<r�a<ˇa<7�a<��a<�a<m�a<
�a<��a<��a<��a<7�a<��a<��a<$�a<��a<9�a<��a<<�a<�a<a<j~a<�}a<�|a<k|a<�{a<a{a<�za<za<Pza<=za<.za<0za<Qza<kza<�za<�za< {a<{a<{a<{a<{a<�za<�za<�za<�za<�za<yza<rza<�za<�za<�za<�za<�za<{a<X{a<�  �  S{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<e{a<p{a<d{a<�{a<�{a<�{a<z|a<�|a<e}a<~a<�~a<qa<�a<̀a<_�a<-�a<��a<[�a<σa<%�a<��a<�a<}�a<څa<G�a<��a<B�a<�a<�a<M�a<��a<��a<8�a<��a<��a<�a<w�a<��a<�a<f�a<��a<�a<B�a<��a<Ϗa<n�a<אa<X�a<�a<��a<m�a<#�a<��a<ȕa<|�a<?�a<�a<��a<�a<��a<�a<S�a<��a<��a<,�a<:�a<|�a<��a<�a<F�a<��a<��a<�a<��a<ĝa<�a<N�a<8�a<\�a<"�a<�a<�a<ԝa<��a<f�a<F�a<�a<7�a<�a<Q�a<w�a<��a<�a<I�a<��a<�a<[�a<��a<�a<1�a<C�a<u�a<4�a<K�a<�a<��a<�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<g�a<3�a<ߞa<q�a<%�a<��a<V�a<Ŝa<h�a<�a<��a<o�a<�a<$�a<�a<�a<�a<&�a<\�a<V�a<~�a<n�a<��a<m�a<h�a<'�a<Ěa<��a<
�a<ԙa<g�a<�a<��a<Q�a<�a<Ηa<��a<:�a<�a<Җa<Z�a<3�a<��a<�a<X�a<��a<�a<:�a<w�a<��a<�a<	�a<��a<�a<Z�a<�a<j�a<>�a<�a<��a<{�a<+�a<�a<��a<g�a<߉a<��a<وa<X�a<̇a<��a<��a<܅a<S�a<��a<@�a<܃a<v�a</�a<��a<��a<�a<��a<`�a<��a<R�a<�a<a<T~a<�}a<}a<||a<�{a<\{a<!{a<�za<�za<_za<7za<^za<^za<�za<�za<�za<�za< {a<&{a<{a<4{a<�za<�za<�za<�za<�za<[za<Uza<Aza<bza<yza<�za<�za<�za<L{a<�  �  L{a<}{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<5|a<�|a<�|a<�}a<$~a<�~a<�a</�a<��a<��a<)�a<��a<(�a<��a<�a<��a<�a<L�a<��a<9�a<��a<�a<ׇa<Y�a<��a<��a<k�a<�a<��a<J�a<֌a<j�a<Սa<W�a<��a<��a<*�a<i�a<ȏa<�a<z�a<��a<��a<!�a<Ғa<��a<J�a<�a<�a<��a<��a<	�a<��a<�a<�a<�a<%�a<�a<��a<�a<�a<n�a<��a<ԛa<6�a<]�a<ɜa<�a<s�a<��a<��a<�a<6�a<R�a<R�a<Q�a<�a<�a<��a<��a<w�a<P�a<D�a<T�a<e�a<��a<ٝa<%�a<|�a<֞a<*�a<��a<ڟa<��a<�a<'�a<<�a<4�a<�a<�a<ٟa<��a<��a<��a<L�a<r�a<w�a<U�a<p�a<��a<��a<|�a<q�a<E�a<!�a<�a<��a<O�a<̝a<h�a<��a<��a<(�a<ța<��a<^�a<0�a<&�a<5�a<6�a<[�a<o�a<��a<��a<��a<��a<h�a<4�a<�a<��a<l�a<
�a<��a<+�a<��a<��a<#�a<�a<��a<d�a<,�a<��a<��a<]�a<�a<~�a<�a<u�a<�a< �a<_�a<��a<Ȑa<�a<R�a<��a<
�a<��a<�a<��a<j�a<�a<ڋa<��a<T�a</�a<��a<]�a<׉a<T�a<ֈa<*�a<��a<��a<T�a<��a<E�a<��a<%�a<̃a<>�a<��a<��a<U�a<�a<��a<%�a<��a<H�a<�a<>a<}~a<�}a<D}a<�|a<$|a<�{a<.{a<�za<�za<{za<vza<{za<�za<�za<�za<�za<{a<{a<{a<�za<�za<�za<�za<�za<kza<<za<Dza<;za<za<Eza<gza<hza<�za<�za<{a<�  �  C{a<\{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a< |a<|a<�|a<�|a<\}a<�}a<P~a<
a<�a<_�a<��a<��a<�a<a<,�a<��a<�a<H�a<��a<�a<{�a<ۅa<^�a<��a<x�a< �a<Ĉa<��a<6�a<܊a<��a<4�a<��a<T�a<эa<;�a<��a<	�a<K�a<��a<�a<m�a<��a<?�a<Αa<X�a<,�a<��a<��a<F�a<�a<��a<a�a<�a<��a<6�a<n�a<�a<�a<E�a<��a<��a<ޚa<�a<W�a<��a<֛a<8�a<��a<�a<2�a<��a<�a<�a<S�a<3�a<N�a<4�a<7�a<�a<�a<��a<��a<��a<{�a<��a<��a<�a< �a<@�a<��a<�a<Z�a<��a<̟a<�a<�a<D�a<�a<-�a<�a<ݟa<��a<|�a<[�a<7�a<9�a<�a<#�a<.�a<A�a<Z�a<L�a<s�a<P�a<]�a<'�a<ڞa<��a<A�a<�a<��a<3�a<��a<g�a<�a<��a<��a<g�a<��a<c�a<b�a<��a<��a<��a<��a<��a<v�a<�a<8�a<�a<��a<)�a<ܙa<m�a<�a<��a<F�a<�a<��a<o�a<,�a<�a<Ėa<v�a<[�a<ەa<��a<��a<p�a<ғa<(�a<��a<��a<�a<-�a<��a<�a<S�a<Ѝa<G�a<�a<��a<M�a<�a<ŋa<j�a<�a<��a<>�a<��a<C�a<ψa<�a<j�a<͆a<�a<��a<�a<h�a<�a<m�a<�a<��a<z�a<�a<ׁa<��a<!�a<Ԁa<(�a<�a<!a<�~a<~a<q}a<�|a<J|a<�{a<d{a</{a<�za<�za<�za<�za<�za<�za<�za<�za<{a<	{a<{a<{a<�za<�za<�za<rza<>za<za<�ya<�ya<�ya<�ya<za<@za<{za<�za<�za<�  �  {a<J{a<{a<�{a<�{a<�{a<�{a<|a<�{a<�{a<|a<|a<7|a<j|a<�|a<}a<�}a<~a<�~a<-a<�a<��a<�a<��a</�a<��a<�a<z�a<ʃa<)�a<{�a<τa<?�a<��a<�a<��a<*�a<߇a<��a<3�a<�a<��a<z�a<�a<Ɍa<V�a<�a<M�a<Ǝa<1�a<o�a<�a<2�a<��a<�a<��a<�a<��a<S�a< �a<˔a<j�a<=�a<�a<q�a<7�a<��a<�a<Q�a<��a<ݙa<�a<0�a<r�a<��a<��a<�a<S�a<��a<��a<L�a<��a<�a<`�a<��a<�a<(�a<P�a<v�a<E�a<`�a<8�a<�a<�a<�a<םa<ҝa<֝a<�a<�a<]�a<��a<��a<�a<��a<��a<ڟa<�a<�a<�a<�a<�a<��a<��a<[�a<J�a<�a<��a<�a<۞a<ݞa<��a<�a<�a<$�a<3�a<=�a<2�a<�a<�a<��a<\�a<*�a<��a<X�a<��a<��a<Q�a<�a<ڛa<��a<��a<��a<��a<��a<��a<כa<��a<a<��a<]�a<�a<Қa<h�a<	�a<��a<'�a<̘a<Q�a<�a<��a<\�a<.�a<��a<��a<��a<N�a<�a<ƕa<q�a<��a<��a<�a<R�a<��a<ߑa<B�a<~�a<ӏa<*�a<��a<	�a<��a<2�a<ьa<��a<$�a<��a<��a< �a<�a<K�a<Ɖa<&�a<��a<�a<C�a<y�a<�a<D�a<��a<!�a<��a<'�a<݂a<~�a<1�a<��a<��a<b�a<��a<��a<E�a<�a<2a<�~a<0~a<�}a<"}a<�|a< |a<�{a<e{a<){a<{a<�za<�za<�za<�za<!{a<{a<{a<3{a<{a<�za<�za<�za<^za<?za<�ya<�ya<�ya<�ya<�ya<�ya<�ya<za<-za<�za<�za<�  �  �za<={a<l{a<�{a<�{a<�{a<|a<|a<*|a<4|a<A|a<Y|a<||a<�|a<�|a<n}a<�}a<Q~a<�~a<ra<�a<��a<3�a<��a<*�a<��a<��a<j�a<��a<��a<=�a<��a<�a<Q�a<Ѕa<G�a<�a<��a<L�a< �a<щa<��a<`�a<�a<��a<Y�a<�a<l�a<��a<R�a<��a<�a<��a<Ԑa<V�a<֑a<]�a<��a<��a<R�a<��a<��a<^�a<�a<��a<#�a<��a<��a<G�a<��a<��a<�a<�a<.�a<=�a<��a<��a<�a<P�a<��a<�a<q�a<��a<@�a<��a<�a<)�a<N�a<g�a<{�a<�a<g�a<X�a<5�a</�a<�a<(�a< �a<K�a<h�a<��a<ܞa<�a<`�a<��a<ޟa<�a<�a<�a<�a<��a<ϟa<��a<g�a<"�a<��a<��a<��a<��a<��a<��a<��a<��a<ߞa<��a<�a<0�a<�a<�a<��a<a<��a<?�a<�a<��a<9�a<�a<��a<l�a<"�a<�a<�a<�a<�a<�a<�a<�a<�a<��a<��a<^�a<�a<��a<H�a<ܙa<[�a<�a<s�a<�a<��a<V�a<"�a<Жa<��a<}�a<_�a<-�a<�a<��a<`�a<��a<��a<�a<��a<Вa<&�a<q�a<ΐa<�a<}�a<�a<^�a<�a<l�a<#�a<��a<j�a<�a<Ëa<F�a<Պa<L�a<��a<�a<��a<��a<�a<K�a<��a<��a<[�a<Ńa<T�a<�a<��a<F�a<��a<a<��a<U�a<�a<��a<C�a<�a<ha<�~a<_~a<�}a<L}a<�|a<Y|a<|a<�{a<�{a<P{a<7{a<2{a<,{a<8{a<9{a<L{a<.{a<({a<{a<�za<�za<{za<9za<�ya<�ya<�ya<Yya<_ya<Bya<nya<zya<�ya<�ya<Fza<�za<�  �  �za<�za<g{a<�{a<�{a<|a<-|a<>|a<T|a<t|a<{|a<�|a<�|a<	}a<b}a<�}a<~a<�~a<a<�a<(�a<��a<?�a<��a<&�a<��a<�a<.�a<��a<��a<�a<N�a<��a<�a<t�a<��a<��a<J�a<��a<Ոa<��a<h�a<?�a<ދa<ˌa<[�a<�a<s�a<�a<s�a<�a<H�a<��a<3�a<��a<*�a<��a<:�a<�a<��a<)�a<�a<��a<$�a<��a<(�a<��a<�a<�a<n�a<��a<��a<ԙa<ܙa<�a<,�a<a�a<��a<��a<d�a<Ǜa<@�a<��a<"�a<u�a<Ɲa<9�a<I�a<y�a<��a<��a<��a<��a<j�a<x�a<k�a<b�a<��a<��a<��a<�a<�a<W�a<��a<��a<�a<��a<�a<�a<
�a<��a<��a<d�a<&�a<�a<��a<��a<Z�a<@�a<=�a<H�a<f�a<��a<��a<��a<��a<�a<�a< �a<��a<מa<��a<`�a<�a<ԝa<s�a<>�a<�a<��a<��a<V�a<A�a<=�a<�a<5�a<�a<�a<�a<̛a<��a<h�a<�a<��a<.�a<��a<&�a<��a<7�a<��a<\�a<
�a<̖a<��a<e�a<R�a<�a<�a<�a<��a<s�a< �a<��a<
�a<��a<�a<\�a<��a<�a<m�a<��a<>�a<��a<*�a<ύa<b�a<�a<��a<3�a<Ӌa<N�a<يa<L�a<҉a<�a<X�a<��a<Æa<�a<O�a<��a<�a<r�a<��a<��a<E�a<��a<ǁa<z�a<c�a<�a<׀a<��a<>�a<�a<wa<
a<�~a<~a<�}a<%}a<�|a<K|a<|a<�{a<�{a<�{a<j{a<k{a<c{a<Y{a<]{a<?{a<'{a<{a<�za<}za<cza<za<�ya<�ya<Lya<ya<ya<�xa<ya<8ya<yya<�ya<za<Zza<�  �  �za<�za<O{a<�{a<�{a</|a<@|a<||a<{|a<�|a<�|a<�|a<}a<J}a<�}a<�}a<_~a<�~a<\a<�a<P�a<��a<L�a<�a<1�a<��a<ӂa<�a<h�a<��a<ރa<��a<p�a<ńa<-�a<Ņa<D�a<"�a<��a<��a<d�a<=�a<�a<ϋa<��a<B�a<"�a<��a<4�a<��a<�a<��a<��a<o�a<ݑa<m�a<��a<��a<*�a<ǔa<{�a<�a<��a<Z�a<��a<\�a<��a<٘a<�a<B�a<l�a<y�a<��a<��a<��a<ۙa<*�a<f�a<��a<4�a<t�a<�a<q�a<��a<O�a<��a<�a<M�a<��a<��a<ٞa<��a<a<Þa<��a<��a<��a<ўa<֞a<�a<,�a<^�a<��a<��a<��a<�a<#�a<-�a<��a<�a<��a<��a<6�a<�a<��a<p�a<S�a<�a<�a<�a<�a<!�a<.�a<|�a<��a<Ԟa<؞a<�a<��a<�a<��a<��a<��a<>�a<�a<��a<r�a<+�a<�a<՜a<��a<��a<q�a<n�a<d�a<;�a<N�a<��a<��a<��a<=�a<��a<e�a<�a<h�a<��a<N�a<��a<��a<�a<Ԗa<u�a<q�a<!�a<�a<�a<וa<��a<v�a<G�a<�a<��a</�a<��a<"�a<{�a<�a<D�a<��a<�a<��a<��a<r�a<	�a<��a<@�a<Ɍa<`�a<	�a<n�a<�a<;�a<��a<�a<-�a<q�a<��a<؅a<	�a<��a<��a<;�a<��a<N�a<�a<��a<��a<S�a<=�a<��a<ŀa<��a<B�a<�a<�a<Ia<�~a<F~a<�}a<U}a<�|a<�|a<`|a<|a<�{a<�{a<�{a<�{a<�{a<�{a<u{a<c{a<E{a<�za<�za<gza<<za<�ya<�ya<2ya<ya<�xa<�xa<�xa<�xa<ya<4ya<hya<�ya<-za<�  �  oza<�za<W{a<�{a<�{a<|a<`|a<�|a<�|a<�|a<�|a<}a<i}a<�}a<�}a<M~a<�~a<a<�a<�a<~�a<�a<r�a<́a<7�a<��a<�a<�a<;�a<n�a<��a<܃a<%�a<z�a<�a<w�a<�a<Ća<��a<Q�a<8�a<�a<�a<�a<��a<b�a<�a<��a<C�a<��a<L�a<��a<3�a<��a<>�a<��a<-�a<�a<V�a<�a<��a<J�a<ǖa<d�a<Ηa<:�a<��a<ޘa<.�a<'�a<@�a<O�a<R�a<v�a<��a<��a<ݙa<�a<u�a<�a<[�a<̛a<S�a<ќa<L�a<͝a<�a<]�a<��a<��a<ܞa<۞a<�a<�a<ޞa<�a<�a<�a<!�a<P�a<P�a<��a<şa<�a<�a<"�a<�a<�a<�a<�a<��a<]�a<�a<Оa<w�a<=�a<��a<͝a<ĝa<��a<��a<�a<�a<F�a<w�a<��a<�a<	�a<�a<�a<�a<ܞa<��a<y�a<<�a<�a<��a<��a<A�a<�a<��a<ќa<��a<��a<��a<i�a<S�a<%�a<ܛa<��a<E�a<�a<f�a<ڙa<O�a<��a<4�a<��a<6�a<іa<��a<A�a<�a<��a<Εa<ŕa<��a<��a<��a<J�a<�a<��a<6�a<Γa<9�a<��a<�a<�a<Аa<e�a<��a<.�a<׎a<5�a<Սa<j�a<�a<{�a<�a<|�a<�a<[�a<��a<�a<�a<E�a<s�a<��a<�a<&�a<�a<�a<o�a<�a<Áa<��a<S�a<5�a<�a<�a<ހa<��a<R�a<�a<�a<Ka<�~a<x~a<�}a<�}a<6}a<�|a<{|a<Z|a<9|a<�{a<�{a<�{a<�{a<�{a<�{a<\{a<3{a<{a<�za<za<	za<�ya<fya<
ya<�xa<�xa<vxa<�xa<�xa<�xa<�xa<Gya<�ya<za<�  �  Mza<�za<{a<�{a<�{a<B|a<�|a<�|a<�|a<�|a<"}a<R}a<x}a<�}a<�}a<d~a<�~a<La<�a<$�a<��a<��a<��a<�a<H�a<q�a<��a<��a<�a<R�a<p�a<��a<�a<c�a<Մa<;�a<�a<��a<d�a<0�a<�a<��a<Ŋa<��a<x�a<m�a<�a<ގa<V�a<ڏa<z�a<��a<l�a<ˑa<N�a<Ēa<P�a<��a<��a<H�a<��a<u�a<�a<l�a<�a<?�a<��a<��a<�a<��a<$�a<'�a<+�a<H�a<=�a<��a<��a<�a<f�a<��a<=�a<��a<3�a<��a<�a<��a<�a<l�a<��a<��a<מa<�a<�a<��a<.�a<�a<�a<�a<;�a<^�a<��a<��a<ǟa<�a<�a<F�a<K�a<#�a<�a<��a<��a<6�a<	�a<��a<X�a<	�a<ǝa<��a<��a<��a<��a<��a<�a<�a<h�a<|�a<��a<Ξa<�a<�a<�a<�a<��a<��a<D�a<�a<ޝa<��a<^�a<!�a<�a<�a<�a<��a<��a<��a<P�a<`�a<��a<��a<.�a<��a<8�a<��a<3�a<��a<�a<p�a<�a<��a<J�a<3�a<ѕa<̕a<��a<��a<��a<h�a<Y�a<�a<�a<��a<u�a<�a<X�a<�a<�a<��a<�a<u�a<؏a<Q�a<�a<e�a<�a<j�a</�a<��a<�a<��a<�a<e�a<��a<Èa<�a<)�a<L�a<t�a<��a<��a<q�a<��a<V�a<��a<{�a<n�a<*�a<�a<�a<a<��a<r�a<a�a<�a<�a<Ga<	a<�~a<~a<�}a<X}a<	}a<�|a<t|a<G|a<,|a<|a<�{a<�{a<�{a<�{a<�{a<;{a<{a<�za<Sza<�ya<�ya</ya<�xa<�xa<cxa<ixa<?xa<rxa<�xa<�xa<&ya<wya<za<�  �  Zza<�za<A{a<�{a<�{a</|a<c|a<�|a<�|a<}a<>}a<a}a<�}a<�}a<P~a<~~a<�~a<Ja<�a<<�a<ƀa<�a<y�a<݁a<2�a<��a<ɂa<�a<�a<)�a<d�a<��a<ރa<:�a<��a<�a<��a<��a<C�a<#�a<�a<�a<ߊa<ŋa<��a<S�a< �a<��a<D�a<��a<w�a<��a<o�a<��a<k�a<	�a<��a<�a<��a<@�a<�a<r�a<�a<i�a<ޗa<>�a<��a<ۘa<�a<�a<�a<�a<&�a<%�a<G�a<T�a<}�a<əa<0�a<��a<�a<��a<�a<��a<2�a<��a<�a<Q�a<��a<Þa<�a<'�a<�a<0�a<&�a<1�a<8�a<t�a<p�a<~�a<��a<֟a<��a< �a<1�a<%�a<2�a<�a<	�a<ܟa<��a<D�a<�a<��a<;�a<�a<��a<|�a<^�a<^�a<��a<��a<ŝa<��a<>�a<��a<Ξa<�a<�a<�a< �a<ޞa<Ӟa<��a<r�a<6�a<�a<��a<��a<z�a<(�a<	�a<�a<�a<��a<��a<g�a<,�a<�a<��a<@�a<֚a<L�a<��a<
�a<��a<�a<j�a<��a<��a<%�a<�a<ٕa<��a<��a<��a<��a<��a<l�a<@�a<��a<��a<K�a<Гa<u�a<�a<Z�a<��a<-�a<��a<�a<��a<��a<��a<�a<��a<-�a<��a<�a<��a<��a<C�a<��a<ڈa<�a<�a<3�a<o�a<��a<�a<,�a<��a<�a<Ɓa<~�a<=�a< �a<�a<�a<ـa<��a<��a<F�a<�a<�a<Ya<a<�~a<G~a<�}a<z}a<!}a<}a<�|a<f|a<G|a<,|a<|a<�{a<�{a<�{a<r{a</{a<�za<�za<bza<�ya<�ya<ya<�xa<�xa<]xa<%xa<xa<1xa<uxa<�xa< ya<eya<�ya<�  �  Iza<�za<({a<�{a<�{a<e|a<�|a<�|a<�|a<}a<E}a<i}a<�}a<�}a<#~a<x~a<a<Ca<�a<2�a<��a<=�a<��a<�a<;�a<|�a<��a<��a<�a<-�a<��a<�a<�a<�a<��a<Q�a<��a<��a<'�a<"�a<�a<�a<��a<��a<��a<N�a<9�a<Ԏa<q�a<�a<T�a<+�a<h�a<�a<x�a<�a<q�a<�a<Ӕa<7�a<�a<R�a<�a<��a<��a<��a<��a<Ҙa<Ҙa<�a<�a<�a<*�a<	�a<R�a<>�a<��a<ڙa<�a<��a<��a<��a<�a<��a<�a<��a<�a<V�a<ٞa<ܞa<�a<�a<�a<Z�a<�a<`�a<5�a<I�a<_�a<��a<��a<ҟa<�a<��a<N�a<K�a<`�a<8�a<�a<˟a<m�a<.�a<ݞa<��a<;�a<�a<��a<i�a<��a<S�a<w�a<��a<��a<�a<4�a<x�a<��a<ڞa< �a<�a<5�a<�a<��a<��a<�a<=�a<��a<�a<y�a<M�a<"�a<=�a<�a<�a<��a<��a<��a<D�a<*�a<��a<9�a<��a<�a<��a<�a<��a<חa<r�a<ږa<��a<`�a<֕a<ەa<��a<��a<��a<|�a<d�a<8�a<3�a<�a<ؔa<k�a<��a<��a<Ēa<��a<��a<H�a<��a<��a<r�a<�a<��a<�a<܍a<�a<Ìa<J�a<��a<3�a<E�a<��a<��a<ۇa<�a<<�a<s�a<|�a<��a<�a<a<+�a<��a<��a<%�a<4�a<�a<�a<��a<��a<��a<K�a<G�a<�a<�a<a<�~a<p~a<�}a<�}a<}a<�|a<�|a<�|a<N|a<(|a<,|a<�{a<�{a<�{a<�{a<P{a<�za<�za<,za<�ya<{ya<7ya<�xa<vxa<Vxa<xa<Txa<'xa<gxa<�xa<�xa<�ya<�ya<�  �  Zza<�za<A{a<�{a<�{a</|a<c|a<�|a<�|a<}a<>}a<a}a<�}a<�}a<P~a<~~a<�~a<Ja<�a<<�a<ƀa<�a<y�a<݁a<2�a<��a<ɂa<�a<�a<)�a<d�a<��a<ރa<:�a<��a<�a<��a<��a<C�a<#�a<�a<�a<ߊa<ŋa<��a<S�a< �a<��a<D�a<��a<w�a<��a<o�a<��a<k�a<	�a<��a<�a<��a<@�a<�a<r�a<�a<i�a<ޗa<>�a<��a<ۘa<�a<�a<�a<�a<&�a<%�a<G�a<T�a<}�a<əa<0�a<��a<�a<��a<�a<��a<2�a<��a<�a<Q�a<��a<Þa<�a<'�a<�a<0�a<&�a<1�a<8�a<t�a<p�a<~�a<��a<֟a<��a< �a<1�a<%�a<2�a<�a<	�a<ܟa<��a<D�a<�a<��a<;�a<�a<��a<|�a<^�a<^�a<��a<��a<ŝa<��a<>�a<��a<Ξa<�a<�a<�a< �a<ޞa<Ӟa<��a<r�a<6�a<�a<��a<��a<z�a<(�a<	�a<�a<�a<��a<��a<g�a<,�a<�a<��a<@�a<֚a<L�a<��a<
�a<��a<�a<j�a<��a<��a<%�a<�a<ٕa<��a<��a<��a<��a<��a<l�a<@�a<��a<��a<K�a<Гa<u�a<�a<Z�a<��a<-�a<��a<�a<��a<��a<��a<�a<��a<-�a<��a<�a<��a<��a<C�a<��a<ڈa<�a<�a<3�a<o�a<��a<�a<,�a<��a<�a<Ɓa<~�a<=�a< �a<�a<�a<ـa<��a<��a<F�a<�a<�a<Ya<a<�~a<G~a<�}a<z}a<!}a<}a<�|a<f|a<G|a<,|a<|a<�{a<�{a<�{a<r{a</{a<�za<�za<bza<�ya<�ya<ya<�xa<�xa<]xa<%xa<xa<1xa<uxa<�xa< ya<eya<�ya<�  �  Mza<�za<{a<�{a<�{a<B|a<�|a<�|a<�|a<�|a<"}a<R}a<x}a<�}a<�}a<d~a<�~a<La<�a<$�a<��a<��a<��a<�a<H�a<q�a<��a<��a<�a<R�a<p�a<��a<�a<c�a<Մa<;�a<�a<��a<d�a<0�a<�a<��a<Ŋa<��a<x�a<m�a<�a<ގa<V�a<ڏa<z�a<��a<l�a<ˑa<N�a<Ēa<P�a<��a<��a<H�a<��a<u�a<�a<l�a<�a<?�a<��a<��a<�a<��a<$�a<'�a<+�a<H�a<=�a<��a<��a<�a<f�a<��a<=�a<��a<3�a<��a<�a<��a<�a<l�a<��a<��a<מa<�a<�a<��a<.�a<�a<�a<�a<;�a<^�a<��a<��a<ǟa<�a<�a<F�a<K�a<#�a<�a<��a<��a<6�a<	�a<��a<X�a<	�a<ǝa<��a<��a<��a<��a<��a<�a<�a<h�a<|�a<��a<Ξa<�a<�a<�a<�a<��a<��a<D�a<�a<ޝa<��a<^�a<!�a<�a<�a<�a<��a<��a<��a<P�a<`�a<��a<��a<.�a<��a<8�a<��a<3�a<��a<�a<p�a<�a<��a<J�a<3�a<ѕa<̕a<��a<��a<��a<h�a<Y�a<�a<�a<��a<u�a<�a<X�a<�a<�a<��a<�a<u�a<؏a<Q�a<�a<e�a<�a<j�a</�a<��a<�a<��a<�a<e�a<��a<Èa<�a<)�a<L�a<t�a<��a<��a<q�a<��a<V�a<��a<{�a<n�a<*�a<�a<�a<a<��a<r�a<a�a<�a<�a<Ga<	a<�~a<~a<�}a<X}a<	}a<�|a<t|a<G|a<,|a<|a<�{a<�{a<�{a<�{a<�{a<;{a<{a<�za<Sza<�ya<�ya</ya<�xa<�xa<cxa<ixa<?xa<rxa<�xa<�xa<&ya<wya<za<�  �  oza<�za<W{a<�{a<�{a<|a<`|a<�|a<�|a<�|a<�|a<}a<i}a<�}a<�}a<M~a<�~a<a<�a<�a<~�a<�a<r�a<́a<7�a<��a<�a<�a<;�a<n�a<��a<܃a<%�a<z�a<�a<w�a<�a<Ća<��a<Q�a<8�a<�a<�a<�a<��a<b�a<�a<��a<C�a<��a<L�a<��a<3�a<��a<>�a<��a<-�a<�a<V�a<�a<��a<J�a<ǖa<d�a<Ηa<:�a<��a<ޘa<.�a<'�a<@�a<O�a<R�a<v�a<��a<��a<ݙa<�a<u�a<�a<[�a<̛a<S�a<ќa<L�a<͝a<�a<]�a<��a<��a<ܞa<۞a<�a<�a<ޞa<�a<�a<�a<!�a<P�a<P�a<��a<şa<�a<�a<"�a<�a<�a<�a<�a<��a<]�a<�a<Оa<w�a<=�a<��a<͝a<ĝa<��a<��a<�a<�a<F�a<w�a<��a<�a<	�a<�a<�a<�a<ܞa<��a<y�a<<�a<�a<��a<��a<A�a<�a<��a<ќa<��a<��a<��a<i�a<S�a<%�a<ܛa<��a<E�a<�a<f�a<ڙa<O�a<��a<4�a<��a<6�a<іa<��a<A�a<�a<��a<Εa<ŕa<��a<��a<��a<J�a<�a<��a<6�a<Γa<9�a<��a<�a<�a<Аa<e�a<��a<.�a<׎a<5�a<Սa<j�a<�a<{�a<�a<|�a<�a<[�a<��a<�a<�a<E�a<s�a<��a<�a<&�a<�a<�a<o�a<�a<Áa<��a<S�a<5�a<�a<�a<ހa<��a<R�a<�a<�a<Ka<�~a<x~a<�}a<�}a<6}a<�|a<{|a<Z|a<9|a<�{a<�{a<�{a<�{a<�{a<�{a<\{a<3{a<{a<�za<za<	za<�ya<fya<
ya<�xa<�xa<vxa<�xa<�xa<�xa<�xa<Gya<�ya<za<�  �  �za<�za<O{a<�{a<�{a</|a<@|a<||a<{|a<�|a<�|a<�|a<}a<J}a<�}a<�}a<_~a<�~a<\a<�a<P�a<��a<L�a<�a<1�a<��a<ӂa<�a<h�a<��a<ރa<��a<p�a<ńa<-�a<Ņa<D�a<"�a<��a<��a<d�a<=�a<�a<ϋa<��a<B�a<"�a<��a<4�a<��a<�a<��a<��a<o�a<ݑa<m�a<��a<��a<*�a<ǔa<{�a<�a<��a<Z�a<��a<\�a<��a<٘a<�a<B�a<l�a<y�a<��a<��a<��a<ۙa<*�a<f�a<��a<4�a<t�a<�a<q�a<��a<O�a<��a<�a<M�a<��a<��a<ٞa<��a<a<Þa<��a<��a<��a<ўa<֞a<�a<,�a<^�a<��a<��a<��a<�a<#�a<-�a<��a<�a<��a<��a<6�a<�a<��a<p�a<S�a<�a<�a<�a<�a<!�a<.�a<|�a<��a<Ԟa<؞a<�a<��a<�a<��a<��a<��a<>�a<�a<��a<r�a<+�a<�a<՜a<��a<��a<q�a<n�a<d�a<;�a<N�a<��a<��a<��a<=�a<��a<e�a<�a<h�a<��a<N�a<��a<��a<�a<Ԗa<u�a<q�a<!�a<�a<�a<וa<��a<v�a<G�a<�a<��a</�a<��a<"�a<{�a<�a<D�a<��a<�a<��a<��a<r�a<	�a<��a<@�a<Ɍa<`�a<	�a<n�a<�a<;�a<��a<�a<-�a<q�a<��a<؅a<	�a<��a<��a<;�a<��a<N�a<�a<��a<��a<S�a<=�a<��a<ŀa<��a<B�a<�a<�a<Ia<�~a<F~a<�}a<U}a<�|a<�|a<`|a<|a<�{a<�{a<�{a<�{a<�{a<�{a<u{a<c{a<E{a<�za<�za<gza<<za<�ya<�ya<2ya<ya<�xa<�xa<�xa<�xa<ya<4ya<hya<�ya<-za<�  �  �za<�za<g{a<�{a<�{a<|a<-|a<>|a<T|a<t|a<{|a<�|a<�|a<	}a<b}a<�}a<~a<�~a<a<�a<(�a<��a<?�a<��a<&�a<��a<�a<.�a<��a<��a<�a<N�a<��a<�a<t�a<��a<��a<J�a<��a<Ոa<��a<h�a<?�a<ދa<ˌa<[�a<�a<s�a<�a<s�a<�a<H�a<��a<3�a<��a<*�a<��a<:�a<�a<��a<)�a<�a<��a<$�a<��a<(�a<��a<�a<�a<n�a<��a<��a<ԙa<ܙa<�a<,�a<a�a<��a<��a<d�a<Ǜa<@�a<��a<"�a<u�a<Ɲa<9�a<I�a<y�a<��a<��a<��a<��a<j�a<x�a<k�a<b�a<��a<��a<��a<�a<�a<W�a<��a<��a<�a<��a<�a<�a<
�a<��a<��a<d�a<&�a<�a<��a<��a<Z�a<@�a<=�a<H�a<f�a<��a<��a<��a<��a<�a<�a< �a<��a<מa<��a<`�a<�a<ԝa<s�a<>�a<�a<��a<��a<V�a<A�a<=�a<�a<5�a<�a<�a<�a<̛a<��a<h�a<�a<��a<.�a<��a<&�a<��a<7�a<��a<\�a<
�a<̖a<��a<e�a<R�a<�a<�a<�a<��a<s�a< �a<��a<
�a<��a<�a<\�a<��a<�a<m�a<��a<>�a<��a<*�a<ύa<b�a<�a<��a<3�a<Ӌa<N�a<يa<L�a<҉a<�a<X�a<��a<Æa<�a<O�a<��a<�a<r�a<��a<��a<E�a<��a<ǁa<z�a<c�a<�a<׀a<��a<>�a<�a<wa<
a<�~a<~a<�}a<%}a<�|a<K|a<|a<�{a<�{a<�{a<j{a<k{a<c{a<Y{a<]{a<?{a<'{a<{a<�za<}za<cza<za<�ya<�ya<Lya<ya<ya<�xa<ya<8ya<yya<�ya<za<Zza<�  �  �za<={a<l{a<�{a<�{a<�{a<|a<|a<*|a<4|a<A|a<Y|a<||a<�|a<�|a<n}a<�}a<Q~a<�~a<ra<�a<��a<3�a<��a<*�a<��a<��a<j�a<��a<��a<=�a<��a<�a<Q�a<Ѕa<G�a<�a<��a<L�a< �a<щa<��a<`�a<�a<��a<Y�a<�a<l�a<��a<R�a<��a<�a<��a<Ԑa<V�a<֑a<]�a<��a<��a<R�a<��a<��a<^�a<�a<��a<#�a<��a<��a<G�a<��a<��a<�a<�a<.�a<=�a<��a<��a<�a<P�a<��a<�a<q�a<��a<@�a<��a<�a<)�a<N�a<g�a<{�a<�a<g�a<X�a<5�a</�a<�a<(�a< �a<K�a<h�a<��a<ܞa<�a<`�a<��a<ޟa<�a<�a<�a<�a<��a<ϟa<��a<g�a<"�a<��a<��a<��a<��a<��a<��a<��a<��a<ߞa<��a<�a<0�a<�a<�a<��a<a<��a<?�a<�a<��a<9�a<�a<��a<l�a<"�a<�a<�a<�a<�a<�a<�a<�a<�a<��a<��a<^�a<�a<��a<H�a<ܙa<[�a<�a<s�a<�a<��a<V�a<"�a<Жa<��a<}�a<_�a<-�a<�a<��a<`�a<��a<��a<�a<��a<Вa<&�a<q�a<ΐa<�a<}�a<�a<^�a<�a<l�a<#�a<��a<j�a<�a<Ëa<F�a<Պa<L�a<��a<�a<��a<��a<�a<K�a<��a<��a<[�a<Ńa<T�a<�a<��a<F�a<��a<a<��a<U�a<�a<��a<C�a<�a<ha<�~a<_~a<�}a<L}a<�|a<Y|a<|a<�{a<�{a<P{a<7{a<2{a<,{a<8{a<9{a<L{a<.{a<({a<{a<�za<�za<{za<9za<�ya<�ya<�ya<Yya<_ya<Bya<nya<zya<�ya<�ya<Fza<�za<�  �  {a<J{a<{a<�{a<�{a<�{a<�{a<|a<�{a<�{a<|a<|a<7|a<j|a<�|a<}a<�}a<~a<�~a<-a<�a<��a<�a<��a</�a<��a<�a<z�a<ʃa<)�a<{�a<τa<?�a<��a<�a<��a<*�a<߇a<��a<3�a<�a<��a<z�a<�a<Ɍa<V�a<�a<M�a<Ǝa<1�a<o�a<�a<2�a<��a<�a<��a<�a<��a<S�a< �a<˔a<j�a<=�a<�a<q�a<7�a<��a<�a<Q�a<��a<ݙa<�a<0�a<r�a<��a<��a<�a<S�a<��a<��a<L�a<��a<�a<`�a<��a<�a<(�a<P�a<v�a<E�a<`�a<8�a<�a<�a<�a<םa<ҝa<֝a<�a<�a<]�a<��a<��a<�a<��a<��a<ڟa<�a<�a<�a<�a<�a<��a<��a<[�a<J�a<�a<��a<�a<۞a<ݞa<��a<�a<�a<$�a<3�a<=�a<2�a<�a<�a<��a<\�a<*�a<��a<X�a<��a<��a<Q�a<�a<ڛa<��a<��a<��a<��a<��a<��a<כa<��a<a<��a<]�a<�a<Қa<h�a<	�a<��a<'�a<̘a<Q�a<�a<��a<\�a<.�a<��a<��a<��a<N�a<�a<ƕa<q�a<��a<��a<�a<R�a<��a<ߑa<B�a<~�a<ӏa<*�a<��a<	�a<��a<2�a<ьa<��a<$�a<��a<��a< �a<�a<K�a<Ɖa<&�a<��a<�a<C�a<y�a<�a<D�a<��a<!�a<��a<'�a<݂a<~�a<1�a<��a<��a<b�a<��a<��a<E�a<�a<2a<�~a<0~a<�}a<"}a<�|a< |a<�{a<e{a<){a<{a<�za<�za<�za<�za<!{a<{a<{a<3{a<{a<�za<�za<�za<^za<?za<�ya<�ya<�ya<�ya<�ya<�ya<�ya<za<-za<�za<�za<�  �  C{a<\{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a< |a<|a<�|a<�|a<\}a<�}a<P~a<
a<�a<_�a<��a<��a<�a<a<,�a<��a<�a<H�a<��a<�a<{�a<ۅa<^�a<��a<x�a< �a<Ĉa<��a<6�a<܊a<��a<4�a<��a<T�a<эa<;�a<��a<	�a<K�a<��a<�a<m�a<��a<?�a<Αa<X�a<,�a<��a<��a<F�a<�a<��a<a�a<�a<��a<6�a<n�a<�a<�a<E�a<��a<��a<ޚa<�a<W�a<��a<֛a<8�a<��a<�a<2�a<��a<�a<�a<S�a<3�a<N�a<4�a<7�a<�a<�a<��a<��a<��a<{�a<��a<��a<�a< �a<@�a<��a<�a<Z�a<��a<̟a<�a<�a<D�a<�a<-�a<�a<ݟa<��a<|�a<[�a<7�a<9�a<�a<#�a<.�a<A�a<Z�a<L�a<s�a<P�a<]�a<'�a<ڞa<��a<A�a<�a<��a<3�a<��a<g�a<�a<��a<��a<g�a<��a<c�a<b�a<��a<��a<��a<��a<��a<v�a<�a<8�a<�a<��a<)�a<ܙa<m�a<�a<��a<F�a<�a<��a<o�a<,�a<�a<Ėa<v�a<[�a<ەa<��a<��a<p�a<ғa<(�a<��a<��a<�a<-�a<��a<�a<S�a<Ѝa<G�a<�a<��a<M�a<�a<ŋa<j�a<�a<��a<>�a<��a<C�a<ψa<�a<j�a<͆a<�a<��a<�a<h�a<�a<m�a<�a<��a<z�a<�a<ׁa<��a<!�a<Ԁa<(�a<�a<!a<�~a<~a<q}a<�|a<J|a<�{a<d{a</{a<�za<�za<�za<�za<�za<�za<�za<�za<{a<	{a<{a<{a<�za<�za<�za<rza<>za<za<�ya<�ya<�ya<�ya<za<@za<{za<�za<�za<�  �  L{a<}{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<5|a<�|a<�|a<�}a<$~a<�~a<�a</�a<��a<��a<)�a<��a<(�a<��a<�a<��a<�a<L�a<��a<9�a<��a<�a<ׇa<Y�a<��a<��a<k�a<�a<��a<J�a<֌a<j�a<Սa<W�a<��a<��a<*�a<i�a<ȏa<�a<z�a<��a<��a<!�a<Ғa<��a<J�a<�a<�a<��a<��a<	�a<��a<�a<�a<�a<%�a<�a<��a<�a<�a<n�a<��a<ԛa<6�a<]�a<ɜa<�a<s�a<��a<��a<�a<6�a<R�a<R�a<Q�a<�a<�a<��a<��a<w�a<P�a<D�a<T�a<e�a<��a<ٝa<%�a<|�a<֞a<*�a<��a<ڟa<��a<�a<'�a<<�a<4�a<�a<�a<ٟa<��a<��a<��a<L�a<r�a<w�a<U�a<p�a<��a<��a<|�a<q�a<E�a<!�a<�a<��a<O�a<̝a<h�a<��a<��a<(�a<ța<��a<^�a<0�a<&�a<5�a<6�a<[�a<o�a<��a<��a<��a<��a<h�a<4�a<�a<��a<l�a<
�a<��a<+�a<��a<��a<#�a<�a<��a<d�a<,�a<��a<��a<]�a<�a<~�a<�a<u�a<�a< �a<_�a<��a<Ȑa<�a<R�a<��a<
�a<��a<�a<��a<j�a<�a<ڋa<��a<T�a</�a<��a<]�a<׉a<T�a<ֈa<*�a<��a<��a<T�a<��a<E�a<��a<%�a<̃a<>�a<��a<��a<U�a<�a<��a<%�a<��a<H�a<�a<>a<}~a<�}a<D}a<�|a<$|a<�{a<.{a<�za<�za<{za<vza<{za<�za<�za<�za<�za<{a<{a<{a<�za<�za<�za<�za<�za<kza<<za<Dza<;za<za<Eza<gza<hza<�za<�za<{a<�  �  S{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<e{a<p{a<d{a<�{a<�{a<�{a<z|a<�|a<e}a<~a<�~a<qa<�a<̀a<_�a<-�a<��a<[�a<σa<%�a<��a<�a<}�a<څa<G�a<��a<B�a<�a<�a<M�a<��a<��a<8�a<��a<��a<�a<w�a<��a<�a<f�a<��a<�a<B�a<��a<Ϗa<n�a<אa<X�a<�a<��a<m�a<#�a<��a<ȕa<|�a<?�a<�a<��a<�a<��a<�a<S�a<��a<��a<,�a<:�a<|�a<��a<�a<F�a<��a<��a<�a<��a<ĝa<�a<N�a<8�a<\�a<"�a<�a<�a<ԝa<��a<f�a<F�a<�a<7�a<�a<Q�a<w�a<��a<�a<I�a<��a<�a<[�a<��a<�a<1�a<C�a<u�a<4�a<K�a<�a<��a<�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<g�a<3�a<ߞa<q�a<%�a<��a<V�a<Ŝa<h�a<�a<��a<o�a<�a<$�a<�a<�a<�a<&�a<\�a<V�a<~�a<n�a<��a<m�a<h�a<'�a<Ěa<��a<
�a<ԙa<g�a<�a<��a<Q�a<�a<Ηa<��a<:�a<�a<Җa<Z�a<3�a<��a<�a<X�a<��a<�a<:�a<w�a<��a<�a<	�a<��a<�a<Z�a<�a<j�a<>�a<�a<��a<{�a<+�a<�a<��a<g�a<߉a<��a<وa<X�a<̇a<��a<��a<܅a<S�a<��a<@�a<܃a<v�a</�a<��a<��a<�a<��a<`�a<��a<R�a<�a<a<T~a<�}a<}a<||a<�{a<\{a<!{a<�za<�za<_za<7za<^za<^za<�za<�za<�za<�za< {a<&{a<{a<4{a<�za<�za<�za<�za<�za<[za<Uza<Aza<bza<yza<�za<�za<�za<L{a<�  �  r{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<i{a<U{a<G{a<U{a<s{a<�{a<�{a<5|a<�|a<G}a<�}a<�~a<Ra<�a<܀a<��a<"�a<��a<?�a<��a<D�a<��a<$�a<��a<��a<e�a<��a<��a<�a<��a<B�a<��a<��a<O�a<Ƌa<Y�a<�a<Y�a<׍a<2�a<~�a<��a<�a<:�a<w�a<֏a<3�a<��a<%�a<Бa<��a<G�a<�a<ߔa<��a<��a<Y�a<�a<��a<�a<��a<�a<m�a<��a<�a<!�a<b�a<��a<��a<0�a<b�a<��a<�a<Y�a<��a<�a<��a<(�a<3�a<G�a<C�a<,�a<��a<��a<y�a<T�a<%�a<�a<�a<�a<�a<T�a<��a<ڝa<=�a<��a<�a<m�a<��a<��a<�a<9�a<B�a<M�a<^�a<6�a<%�a<��a<ݟa<ɟa<��a<��a<��a<��a<��a<��a<��a<��a<u�a<X�a< �a<�a<��a<3�a<��a<,�a<��a<?�a<��a<��a<2�a<��a<ߚa<�a<�a<��a<�a<<�a<e�a<��a<��a<��a<c�a<K�a<	�a<�a<��a<C�a<�a<��a<"�a<��a<��a<3�a<�a<��a<s�a<#�a<�a<i�a< �a<��a<��a<v�a<ɓa<
�a<7�a<S�a<��a<Ïa<�a<Z�a<��a<&�a<��a<t�a<�a<�a<��a<r�a<E�a<�a<��a<D�a<��a<d�a<܈a<r�a<ˇa<7�a<��a<�a<m�a<
�a<��a<��a<��a<7�a<��a<��a<$�a<��a<9�a<��a<<�a<�a<a<j~a<�}a<�|a<k|a<�{a<a{a<�za<za<Pza<=za<.za<0za<Qza<kza<�za<�za< {a<{a<{a<{a<{a<�za<�za<�za<�za<�za<yza<rza<�za<�za<�za<�za<�za<{a<X{a<�  �  �|a<}a<>}a<5}a<P}a<U}a<<}a<X}a<B}a<;}a</}a<Y}a<�}a<�}a<�}a<E~a<�~a<5a<�a<f�a< �a<��a<K�a<�a<��a<&�a<��a< �a<��a<��a<��a<�a<w�a<�a<O�a<ֈa<s�a<=�a<��a<Y�a<�a<m�a<$�a<��a<.�a<��a<�a<e�a<��a<0�a<e�a<��a<��a<��a<��a<Y�a<�a<��a<5�a<��a<}�a<;�a<�a<��a<S�a<�a<��a<)�a<��a<
�a<Q�a<��a<�a<�a<��a<��a<�a<1�a<��a<�a<��a<c�a<��a<�a<�a<G�a<V�a<Q�a<b�a<3�a<*�a<�a<�a<a<��a<��a<��a<��a<��a<��a<>�a<Q�a<��a<��a<f�a<��a<٠a<�a<&�a<^�a<\�a<u�a<C�a<G�a<?�a<�a<>�a<�a<ՠa<Рa<�a<Ӡa<Ԡa<ʠa<��a< a<��a<��a<5�a<�a<��a<N�a<�a<��a<4�a<��a<�a<7�a<�a<��a<��a<��a<s�a<t�a<��a<��a<��a<��a<��a<��a<��a<n�a<!�a<�a<��a<O�a<�a<��a<^�a<�a<��a<]�a<G�a<��a<��a<7�a<Ηa<��a<�a<��a<�a<��a<ܔa<,�a<��a<Òa<�a<?�a<̐a<"�a<w�a<��a<��a</�a<��a<f�a<�a<��a<��a<:�a<�a<��a<2�a<��a<@�a<��a<�a<��a<�a<��a<�a<X�a<�a<~�a<%�a<��a<M�a<уa<��a<�a<��a<>�a<��a<8�a<��a<�a<~a<�~a<C~a<�}a<g}a<�|a<�|a<_|a<R|a<H|a<|a<0|a<F|a<u|a<a|a<�|a<�|a<�|a<�|a<�|a<�|a<R|a<N|a<B|a<|a<K|a<
|a< |a<|a<a|a<T|a<}|a<�|a<�|a<�  �  �|a<	}a<)}a<8}a<G}a<S}a<b}a<D}a<@}a<I}a<[}a<b}a<}a<�}a<~a<g~a<�~a<Qa<�a<v�a<�a<��a<y�a<�a<��a<�a<��a<"�a<��a<�a<�a<�a<Q�a<·a<X�a<�a<d�a<�a<��a<:�a<�a<��a<�a<��a<"�a<��a<�a<��a<܏a< �a<|�a<Ԑa<0�a<��a<�a<s�a<��a<��a</�a<�a<��a<U�a<�a<̗a<�a<�a<��a<�a<��a<��a<_�a<��a<�a< �a<Y�a<��a<��a<:�a<p�a<��a<�a<Y�a<��a<�a<�a<3�a<D�a<X�a<R�a<f�a<7�a<�a<��a<�a<Ȟa<��a<��a<��a<�a<��a<7�a<��a<ßa<�a<P�a<��a<�a<
�a<3�a<M�a<Z�a<f�a<g�a<E�a<*�a<�a<�a<�a<�a<Ҡa<��a<��a<àa<Ơa<Πa<��a<��a<o�a<9�a<��a<��a<t�a<��a<��a<B�a<�a<��a<4�a<�a<˜a<��a<��a<��a<��a<��a<��a<��a<Ϝa<��a<��a<�a<]�a<"�a<��a<��a<K�a<�a<��a<=�a<��a<��a<M�a<��a<��a<x�a<3�a<�a<��a<�a<��a<�a<��a<��a<M�a<��a<ڒa<&�a<v�a<��a<�a<��a<�a<��a<)�a<܍a<��a<9�a<�a<��a<e�a<��a<��a<%�a<��a<2�a<��a<�a<��a<�a<T�a<ӆa<k�a<�a<g�a<��a<��a<D�a<�a<��a<�a<��a<,�a<��a<(�a<��a<�a<oa<�~a<k~a<�}a<f}a<}a<�|a<�|a<M|a<A|a<E|a<F|a<L|a<_|a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<v|a<L|a<-|a<
|a<�{a<|a<|a<|a<|a<9|a<m|a<�|a<�|a<�  �  �|a<}a<}a<K}a<]}a<A}a<]}a<D}a<k}a<P}a<i}a<t}a<�}a<�}a<~a<�~a<�~a<`a<�a<��a<2�a<��a<r�a<�a<��a<&�a<��a<'�a<��a<�a<Y�a<�a<Y�a<·a<=�a<��a<_�a<�a<��a<"�a<ċa<r�a<��a<��a<�a<��a<�a<v�a<ڏa<&�a<��a<ʐa<D�a<��a<�a<��a<	�a<��a<7�a<��a<��a<{�a<�a<ȗa<q�a<��a<��a<�a<��a<�a<J�a<��a<ța<?�a<O�a<��a<Ϝa<�a<r�a<��a<�a<5�a<��a<��a<�a<7�a<K�a<y�a<;�a<]�a<2�a<)�a<�a<�a<Ӟa<��a<ڞa<��a<��a<�a<C�a<��a<şa<1�a<O�a<��a<Ѡa<�a<I�a<@�a<d�a<@�a<O�a<'�a<#�a<*�a<�a<ݠa< a< a<��a<֠a< a<��a<��a<��a<��a<c�a<L�a<�a<��a<o�a<��a<ƞa<I�a<��a<��a<B�a<�a<Μa<Мa<��a<��a<��a<��a<��a<��a<ɜa<��a<��a<��a<]�a<(�a<̛a<��a<%�a<�a<��a<=�a<ڙa<��a<H�a<�a<ۘa<`�a<�a<ӗa<l�a<!�a<��a<5�a<�a<�a<J�a<��a<��a<�a<��a<Őa</�a<��a<�a<��a<0�a<�a<��a<_�a<�a<��a<X�a<�a<��a<%�a<��a<%�a<��a<�a<f�a<	�a<J�a<҆a<=�a<ąa<i�a<��a<��a<�a<Ճa<g�a<�a<��a<3�a<ցa<�a<��a<�a<�a<a<f~a<�}a<e}a</}a<�|a<�|a<]|a<M|a<W|a<G|a<w|a<^|a<�|a<�|a<�|a<�|a<�|a<�|a<]|a<]|a<-|a<&|a</|a<�{a<�{a<�{a<|a<|a<X|a<k|a<w|a<�|a<�  �  �|a<�|a<}a<1}a<b}a<h}a<`}a<e}a<j}a<l}a<�}a<�}a<�}a<�}a<0~a<�~a<a<�a<�a<��a<:�a<Ёa<o�a<�a<��a<�a<��a<�a<��a<�a<O�a<��a<!�a<��a<$�a<��a<4�a<ŉa<\�a<�a<��a<V�a<��a<��a<�a<��a<)�a<��a<�a<?�a<��a<�a<]�a<ˑa<4�a<��a<&�a<̓a<r�a<�a<��a<|�a<+�a<ڗa<��a<$�a<��a<�a<x�a<�a<0�a<�a<��a<�a<*�a<q�a<��a<��a<B�a<��a<ϝa<(�a<w�a<��a<�a<�a<7�a<[�a<l�a<_�a<I�a<9�a<$�a<�a<�a<�a<�a<�a<�a<=�a<}�a<��a<�a<+�a<n�a<��a<�a<&�a<)�a<6�a<B�a<J�a<.�a<�a<��a<٠a<Ǡa<��a<��a<��a<��a<��a<��a<��a<��a<��a<{�a<V�a<1�a<�a<ϟa<r�a<�a<Şa<e�a<�a<˝a<u�a<2�a<��a<��a<ɜa<Мa<��a<��a<ǜa<Ĝa<Ɯa<Ȝa<��a<s�a<D�a<	�a<ɛa<v�a<�a<��a<^�a<�a<��a<i�a<�a<Ϙa<��a<L�a<�a<��a<l�a<��a<��a<�a<��a<�a<Y�a<��a<��a<C�a<��a<�a<_�a<��a<7�a<Ўa<k�a<�a<��a<`�a<�a<��a<k�a<�a<��a<�a<��a<�a<��a<��a<V�a<��a<&�a<��a<#�a<��a<8�a<Ǆa<b�a<�a<��a<_�a<��a<��a<�a<��a<C�a<��a<!�a<�a<a<�~a<~a<�}a<D}a<�|a<�|a<�|a<�|a<n|a<e|a<q|a<}|a<�|a<�|a<�|a<�|a<~|a<r|a<f|a<=|a<%|a<|a<�{a<�{a<�{a<�{a<�{a<�{a<|a<@|a<o|a<�|a<�  �  �|a<�|a<5}a<>}a<?}a<i}a<p}a<�}a<t}a<�}a<�}a<�}a<�}a<'~a<z~a<�~a<'a<�a<7�a<ŀa<K�a<�a<v�a<�a<{�a<1�a<��a<�a<|�a<��a<=�a<��a<�a<h�a<�a<|�a<�a<��a<:�a<��a<��a<;�a<��a<g�a<>�a<��a<�a<��a<�a<g�a<��a<5�a<r�a<ڑa<N�a<�a<r�a<�a<��a<+�a<��a<��a<I�a<��a<~�a<%�a<��a<9�a<e�a<ߚa<�a<U�a<��a<ța<�a<,�a<��a<ɜa<�a<u�a<��a<�a<F�a<��a<�a<�a<_�a<?�a<u�a<_�a<y�a<M�a<?�a<9�a<�a<
�a<�a<6�a<H�a<W�a<��a<ȟa<"�a<8�a<��a<àa<�a<	�a<-�a<e�a<�a<G�a<�a<��a<ߠa<��a<��a<y�a<��a<c�a<e�a<n�a<t�a<��a<j�a<��a<X�a<{�a<?�a<��a<ϟa<��a<P�a<Оa<��a<4�a<؝a<��a<g�a<@�a<�a<�a<ܜa<�a<�a<؜a<��a<̜a<Ϝa<��a<��a<R�a<��a<śa<F�a<�a<��a<I�a<יa<��a<A�a<ژa<��a<`�a<5�a<�a<��a<e�a<ܖa<��a<
�a<��a<��a<u�a<ϓa<�a<��a<��a<�a<y�a<�a<��a<�a<��a<�a<�a<r�a<*�a<܌a<e�a<�a<��a<B�a<��a<�a<m�a<ˈa<D�a<��a<�a<_�a<��a<y�a<��a<��a<B�a<�a<��a<W�a<�a<��a<G�a<��a<K�a<��a<R�a<�a<.a<�~a<*~a<�}a<b}a<1}a<�|a<�|a<�|a<�|a<�|a<|a<�|a<�|a<�|a<�|a<�|a<�|a<O|a<d|a<|a<|a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<|a<W|a<q|a<�  �  �|a<�|a<}a<7}a<c}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<~a<a~a<�~a<a<`a<�a<^�a<�a<o�a<�a<��a</�a<��a<�a<t�a<�a<O�a<��a<
�a<]�a<ӆa<B�a<��a<8�a<̈a<l�a<#�a<��a<r�a<�a<ьa<\�a<�a<��a<1�a<��a<�a<v�a<ސa<B�a<��a<#�a<��a<�a<��a<3�a<ϔa<s�a<�a<��a<[�a<�a<��a<1�a<��a<�a<V�a<��a<��a<8�a<i�a<��a<֛a<�a<G�a<��a<ݜa<6�a<��a<��a<+�a<��a<Ҟa<��a<J�a<d�a<��a<t�a<��a<l�a<f�a<T�a<V�a<H�a<S�a<L�a<x�a<��a<ϟa<�a<5�a<k�a<��a<נa<�a<)�a<.�a<7�a<�a<�a<�a<ՠa<��a<��a<m�a<O�a<4�a<2�a<;�a<J�a<;�a<V�a<U�a<n�a<Q�a<K�a<8�a<�a<�a<��a<U�a<��a<��a<n�a<$�a<Нa<��a<W�a<O�a<&�a<�a<�a<�a<��a<��a<�a<�a<��a<��a<)�a<�a<��a<-�a<֚a<c�a<�a<��a<I�a<��a<��a<v�a<I�a<��a<×a<{�a<>�a<іa<��a<�a<��a<�a<��a<ޓa<<�a<��a<��a<[�a<��a<&�a<��a<7�a<Ȏa<c�a<��a<��a<=�a<�a<}�a<�a<��a<%�a<t�a<��a<M�a<��a<�a<s�a<цa<:�a<��a<6�a<Ԅa<x�a<�a<ʃa<q�a<,�a<ނa<q�a<1�a<��a<Z�a<ʀa<[�a<�a<Ua<�~a<n~a<�}a<�}a<G}a<}a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<|a<F|a<;|a<�{a<�{a<�{a<�{a<z{a<i{a<`{a<v{a<�{a<�{a<�{a<+|a<\|a<�  �  u|a<�|a<�|a<,}a<X}a<{}a<�}a<�}a<�}a<�}a<~a<#~a<J~a<�~a<�~a<Oa<�a<�a<��a<�a<��a<�a<��a< �a<��a<�a<p�a<ڄa<�a<��a<مa<9�a<��a<�a<��a<�a<��a<�a<��a<��a<X�a<��a<��a<l�a<�a<��a<&�a<��a<+�a<��a<�a<n�a<�a<D�a<Ӓa<E�a<ѓa<v�a<�a<��a<<�a<��a<v�a<�a<��a<)�a<��a<��a<b�a<��a<˚a<!�a<7�a<|�a<��a<�a<�a<W�a<��a<�a<Y�a<��a< �a<P�a<��a<��a<+�a<Y�a<{�a<��a<��a<��a<��a<�a<��a<i�a<��a<��a<��a<Οa<�a<0�a<c�a<��a<��a<��a<�a<�a<%�a<�a<�a<�a<ՠa<��a<w�a<]�a<�a<0�a<��a<�a<�a<�a<�a</�a<@�a<7�a<S�a<:�a<,�a<�a<�a<��a<e�a<7�a<�a<��a<I�a< �a<�a<��a<��a<L�a<Z�a<9�a<@�a<+�a<�a<	�a<՜a<��a<i�a<$�a<ۛa<d�a<"�a<��a<@�a<ʙa<t�a<!�a<Ƙa<��a<'�a<�a<ŗa<��a<V�a<�a<�a<|�a<�a<��a<+�a<��a<�a<}�a<��a<.�a<|�a<��a<c�a<�a<z�a<�a<��a<%�a<ލa<X�a<�a<��a<�a<��a<�a<��a<Չa<�a<��a<ԇa<E�a<��a<�a<��a<�a<��a<0�a<�a<��a<f�a<��a<a<q�a<�a<��a<Q�a<�a<p�a<�a<�a< a<�~a<~a<�}a<�}a<`}a<$}a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<d|a<M|a<|a<�{a<�{a<{{a<b{a<,{a<J{a<#{a<W{a<O{a<�{a<�{a<|a<G|a<�  �  e|a<�|a< }a<6}a<f}a<�}a<�}a<�}a<�}a<~a<)~a<h~a<�~a<�~a<a<na<�a<Y�a<��a<=�a<��a<I�a<��a<=�a<��a<�a<q�a<��a<	�a<X�a<��a<�a<j�a<ʆa<D�a<��a<a�a<��a<��a<[�a<�a<Ћa<��a<A�a<�a<��a<F�a<��a<L�a<��a<-�a<��a<�a<��a< �a<y�a<�a<��a<7�a<וa<q�a<�a<��a<A�a<��a<G�a<��a<�a<<�a<��a<��a<��a<
�a<@�a<n�a<��a<Λa<�a<n�a<˜a<)�a<}�a<ߝa<>�a<��a<�a<7�a<^�a<��a<��a<��a<��a<��a<��a<ɟa<��a<��a<ɟa<�a<�a<8�a<T�a<��a<��a<�a<�a<�a<2�a<0�a<+�a<��a<ܠa<��a<�a<P�a<'�a<��a<�a<��a<Οa<��a<ܟa<�a<��a<
�a<'�a<1�a<F�a<6�a<�a<�a<��a<��a<J�a<�a<��a<��a<I�a<�a<ӝa<��a<��a<��a<j�a<_�a<C�a<=�a< �a<�a<��a<v�a<%�a<��a<R�a<�a<w�a<�a<��a<9�a<��a<��a<K�a<	�a<ؗa<��a<k�a<1�a<�a<��a<��a<�a<��a<)�a<��a<)�a<��a<��a<W�a<Ƒa<+�a<��a<�a<��a<1�a<Ȏa<Z�a<�a<��a<$�a<��a<5�a<��a<�a<Z�a<��a<�a<V�a<��a<	�a<i�a<Յa<=�a<Ȅa<d�a<�a<��a<g�a<$�a<�a<��a<f�a<�a<��a<o�a<�a<��a<�a<�a<4a<�~a<m~a<~a<�}a<�}a<e}a<B}a<}a<}a<�|a<�|a<�|a<�|a<�|a<�|a<s|a<*|a<�{a<�{a<�{a<T{a<-{a<{a<{a<�za<{a<!{a<^{a<�{a<�{a<|a<�  �  a|a<�|a<�|a<}a<q}a<�}a<�}a<~a<~a<D~a<`~a<�~a<�~a<�~a<]a<�a<
�a<m�a<��a<h�a<сa<q�a<��a<h�a<��a<��a<R�a<��a<�a<%�a<��a<΅a<!�a<��a<�a<��a<�a<��a<m�a<D�a<�a<��a<��a<-�a<��a<�a<\�a<̏a<`�a<�a<G�a<ߑa<<�a<Βa<$�a<��a<G�a<��a<}�a<��a<��a<*�a<ʗa<\�a<��a<b�a<��a<��a<'�a<y�a<��a<��a<��a<��a<'�a<X�a<��a<��a<*�a<��a<�a<r�a<��a<1�a<��a<Оa<!�a<S�a<��a<��a<�a<ԟa<�a<�a<ޟa<��a<�a<�a<�a<8�a<m�a<��a< a<̠a<�a<�a<=�a<B�a<�a<�a<�a<נa<}�a<\�a<$�a<�a<��a<��a<��a<��a<��a<��a<��a<ޟa<ޟa<$�a<�a<,�a<�a<'�a<�a<ǟa<Ɵa<_�a<=�a<�a<��a<s�a<;�a<#�a<ܝa<ϝa<��a<��a<��a<^�a<f�a<
�a<�a<��a<Y�a<�a<��a<J�a<��a<h�a<ՙa<^�a<��a<��a<j�a<�a<Ǘa<��a<��a<C�a<�a<��a<��a<v�a<��a<וa<C�a<Дa<P�a<��a<1�a<��a<�a<O�a<ِa<X�a<��a<w�a<�a<��a<�a<��a<?�a<��a<P�a<~�a<�a<D�a<��a<�a<+�a<��a<Æa<"�a<��a<"�a<��a<!�a<Ńa<{�a<]�a<��a<؂a<��a<G�a<	�a<��a<��a<�a<��a<5�a<�a<oa<�~a<�~a<8~a<~a<�}a<�}a<w}a<K}a<D}a<}a<'}a<�|a<�|a<�|a<m|a<\|a<|a<�{a<�{a<c{a<({a<�za<�za<�za<�za<�za<�za<{a<`{a<�{a<�{a<�  �  /|a<�|a<�|a<5}a<^}a<�}a<�}a<~a<-~a<Z~a<�~a<�~a<�~a<9a<a<�a<0�a<��a<�a<��a<��a<t�a<ւa<6�a<��a<�a<S�a<��a<҄a<�a<X�a<��a<�a<q�a<܆a<W�a< �a<��a<^�a<�a<܊a<��a<c�a<0�a<�a<��a<2�a<Ϗa<k�a<�a<w�a<�a<[�a<ݒa<e�a<�a<v�a<�a<��a<�a<��a<V�a<ݗa<e�a<˘a<5�a<��a<��a<,�a<U�a<�a<��a<��a<�a<�a<=�a<g�a<��a<�a<w�a<Ϝa<,�a<��a<�a<p�a<֞a<1�a<X�a<��a<��a<�a<�a<�a<	�a<�a<�a<$�a<6�a<W�a<g�a<��a<��a<ՠa<��a<�a<%�a<)�a<%�a<)�a<�a<ؠa<��a<n�a<2�a<��a<֟a<��a<y�a<X�a<]�a<g�a<��a<��a<��a<ӟa<�a<
�a<*�a<6�a<�a<��a<�a<ȟa<��a<S�a<�a<՞a<��a<y�a<E�a<�a<��a<ϝa<��a<��a<��a<h�a<,�a<�a<��a<q�a<�a<��a<�a<��a<$�a<��a<V�a<ߘa<x�a<�a<�a<��a<��a<N�a<-�a<�a<Жa<��a<n�a<�a<��a<F�a<۔a<[�a<Փa<@�a<��a<�a<��a<�a<��a<�a<��a<	�a<��a<:�a<��a<H�a<��a<#�a<��a< �a<J�a<��a<҈a<�a<Z�a<��a<	�a<o�a<Մa<b�a<�a<��a<b�a<�a<�a<��a<}�a<M�a<�a<��a<a�a<�a<��a<S�a<�a<�a<a<�~a<y~a<1~a<�}a<�}a<�}a<p}a<W}a<>}a<*}a<}a<�|a<�|a<�|a<W|a<|a<�{a<~{a<8{a<�za<�za<�za<�za<�za<�za<�za<{a<={a<�{a<�{a<�  �  |a<�|a<�|a<5}a<w}a<�}a<�}a<
~a<N~a<b~a<�~a<�~a<a<Ua<�a<�a<Q�a<�a</�a<��a<�a<n�a<��a<A�a<��a<��a<8�a<��a<��a<�a<8�a<��a<܅a<:�a<ǆa<0�a<�a<g�a<2�a<�a<ъa<��a<N�a<)�a<��a<��a<D�a<�a<�a< �a<��a<��a<��a<
�a<��a<�a<��a<0�a<��a<p�a<Ζa<i�a<�a<r�a<�a<E�a<��a<řa<�a<B�a<h�a<��a<��a<Ța<՚a<�a<E�a<��a<ޛa<8�a<��a<�a<��a<�a<e�a<��a<�a<}�a<��a<�a<�a<�a<�a<!�a<Y�a<2�a<M�a<S�a<r�a<��a<��a<�a<ޠa<�a<�a<E�a<@�a<=�a<9�a<�a<ڠa<��a<i�a<�a<��a<��a<c�a<h�a<2�a<J�a<3�a<S�a<z�a<��a<џa<Οa<�a<��a<6�a<-�a<�a<�a<ğa<��a<[�a<E�a<�a<ɞa<��a<_�a<C�a<�a<#�a<�a<��a<��a<b�a<N�a<��a<͜a<]�a<�a<��a<��a<��a<�a<��a<�a<��a<c�a<��a<їa<q�a<X�a<(�a<#�a<�a<��a<��a<:�a<5�a<��a<h�a<�a<h�a<�a<O�a<�a<C�a<��a<"�a<��a<4�a<��a<`�a<��a<M�a<Սa<U�a<،a<4�a<��a<ϊa<:�a<y�a<��a<�a<2�a<��a<Ѕa<O�a<��a<K�a<ԃa<z�a<K�a<��a<�a<��a<r�a<6�a<��a<فa<n�a<6�a<��a<p�a<�a<�a<qa<�~a<�~a<N~a<~a<�}a<�}a<�}a<a}a<]}a<+}a<"}a<�|a<�|a<�|a<)|a<
|a<�{a<x{a<#{a<�za<�za<qza<�za<^za<�za<�za<�za<#{a<h{a<�{a<�  �  |a<�|a<�|a<}a<e}a<�}a<�}a</~a<f~a<�~a<�~a<�~a<a<ha<�a<�a<Y�a<��a<9�a<��a<0�a<��a<�a<L�a<��a<�a<G�a<��a<��a<�a<;�a<��a<҅a<)�a<��a<.�a<ʇa<g�a<'�a<�a<��a<s�a<S�a<4�a<؍a<��a<?�a<�a<~�a< �a<��a<�a<��a<�a<��a<.�a<��a</�a<��a<T�a<�a<��a<
�a<x�a<�a<D�a<��a<ޙa<*�a<H�a<T�a<z�a<��a<��a<Ϛa<�a<=�a<��a<˛a<0�a<��a<�a<}�a<�a<g�a<̞a<�a<e�a<��a<ԟa<�a<'�a<,�a<4�a<2�a<=�a<U�a<��a<��a<��a<��a<ݠa<�a</�a<C�a<=�a<B�a<0�a<�a<�a<ޠa<��a<F�a<�a<۟a<��a<a�a<G�a<-�a<.�a<)�a<A�a<o�a<��a<��a<Пa<�a<�a<�a<�a<�a<��a<�a<a<��a<D�a< �a<Ϟa<��a<��a<N�a<�a<��a<�a<ѝa<��a<��a<E�a<�a<��a<W�a<��a<��a<��a<�a<�a<��a<�a<��a<J�a<�a<��a<q�a<M�a<.�a<�a<Ԗa<��a<��a<R�a<�a<��a<c�a<�a<��a<�a<q�a<ڒa<F�a<��a<L�a<̐a<3�a<��a<D�a<֎a<e�a<�a<Z�a<ьa<2�a<��a<�a<H�a<~�a<��a<��a<;�a<��a<ʅa<5�a<��a<5�a<��a<r�a<7�a<��a<Âa<��a<s�a<D�a<��a<��a<u�a<)�a<܀a<��a<�a<�a<Ja<�~a<�~a<|~a<.~a<�}a<�}a<�}a<�}a<v}a<R}a<}a<�|a<�|a<�|a<8|a<|a<�{a<V{a<{a<�za<�za<nza<aza<Yza<rza<�za<�za<{a<^{a<�{a<�  �  !|a<^|a<�|a<$}a<d}a<�}a<�}a<6~a<B~a<�~a<�~a<�~a<Ta<da<�a<�a<��a<̀a<R�a<��a<�a<��a<�a<Z�a<��a<��a<6�a<c�a<ʄa<�a<#�a<U�a<ޅa<2�a<��a<�a<��a<f�a< �a<ɉa<��a<��a<B�a<�a<�a<��a<S�a<�a<��a< �a<��a<+�a<��a<?�a<��a<$�a<��a<<�a<��a<J�a<�a<z�a<�a<��a<��a<S�a<��a<�a<��a<0�a<e�a<a�a<w�a<��a<њa<��a<'�a<f�a<՛a<?�a<m�a<�a<i�a<��a<B�a<��a<!�a<P�a<��a<՟a<�a<�a<1�a<Q�a<7�a<��a<e�a<h�a<�a<àa<֠a<�a<�a<	�a<D�a<;�a<S�a<6�a<�a<��a<��a<��a<T�a<��a<��a<{�a<e�a<&�a<#�a<�a<+�a<2�a<F�a<{�a<��a<�a<�a<�a<$�a<�a<+�a<��a<�a<��a<��a<Q�a<�a<	�a<��a<s�a<Z�a<o�a<�a<�a<ԝa<��a<��a<G�a<�a<��a<a�a<�a<d�a<�a<t�a<�a<\�a<�a<��a<#�a<ܗa<��a<p�a<&�a<�a<�a<�a<��a<v�a<c�a<�a<͕a<y�a<��a<��a<�a<~�a<Ғa<x�a<ёa<B�a<��a<A�a<��a<;�a<�a<^�a<�a<h�a<ތa<A�a<��a<�a<�a<f�a<��a<ׇa<�a<R�a<̅a<&�a<��a<�a<̃a<��a<�a<܂a<��a<��a<O�a<*�a<	�a<��a<��a<*�a<�a<i�a< �a<�a<Oa<Aa<�~a<b~a<$~a<~a<�}a<�}a<�}a<O}a<S}a<}a<}a<�|a<�|a<F|a<�{a<�{a<c{a<{a<�za<�za<rza<@za<Pza<Sza<�za<�za<�za<Q{a<�{a<�  �  |a<�|a<�|a<}a<e}a<�}a<�}a</~a<f~a<�~a<�~a<�~a<a<ha<�a<�a<Y�a<��a<9�a<��a<0�a<��a<�a<L�a<��a<�a<G�a<��a<��a<�a<;�a<��a<҅a<)�a<��a<.�a<ʇa<g�a<'�a<�a<��a<s�a<S�a<4�a<؍a<��a<?�a<�a<~�a< �a<��a<�a<��a<�a<��a<.�a<��a</�a<��a<T�a<�a<��a<
�a<x�a<�a<D�a<��a<ޙa<*�a<H�a<T�a<z�a<��a<��a<Ϛa<�a<=�a<��a<˛a<0�a<��a<�a<}�a<�a<g�a<̞a<�a<e�a<��a<ԟa<�a<'�a<,�a<4�a<2�a<=�a<U�a<��a<��a<��a<��a<ݠa<�a</�a<C�a<=�a<B�a<0�a<�a<�a<ޠa<��a<F�a<�a<۟a<��a<a�a<G�a<-�a<.�a<)�a<A�a<o�a<��a<��a<Пa<�a<�a<�a<�a<�a<��a<�a<a<��a<D�a< �a<Ϟa<��a<��a<N�a<�a<��a<�a<ѝa<��a<��a<E�a<�a<��a<W�a<��a<��a<��a<�a<�a<��a<�a<��a<J�a<�a<��a<q�a<M�a<.�a<�a<Ԗa<��a<��a<R�a<�a<��a<c�a<�a<��a<�a<q�a<ڒa<F�a<��a<L�a<̐a<3�a<��a<D�a<֎a<e�a<�a<Z�a<ьa<2�a<��a<�a<H�a<~�a<��a<��a<;�a<��a<ʅa<5�a<��a<5�a<��a<r�a<7�a<��a<Âa<��a<s�a<D�a<��a<��a<u�a<)�a<܀a<��a<�a<�a<Ja<�~a<�~a<|~a<.~a<�}a<�}a<�}a<�}a<v}a<R}a<}a<�|a<�|a<�|a<8|a<|a<�{a<V{a<{a<�za<�za<nza<aza<Yza<rza<�za<�za<{a<^{a<�{a<�  �  |a<�|a<�|a<5}a<w}a<�}a<�}a<
~a<N~a<b~a<�~a<�~a<a<Ua<�a<�a<Q�a<�a</�a<��a<�a<n�a<��a<A�a<��a<��a<8�a<��a<��a<�a<8�a<��a<܅a<:�a<ǆa<0�a<�a<g�a<2�a<�a<ъa<��a<N�a<)�a<��a<��a<D�a<�a<�a< �a<��a<��a<��a<
�a<��a<�a<��a<0�a<��a<p�a<Ζa<i�a<�a<r�a<�a<E�a<��a<řa<�a<B�a<h�a<��a<��a<Ța<՚a<�a<E�a<��a<ޛa<8�a<��a<�a<��a<�a<e�a<��a<�a<}�a<��a<�a<�a<�a<�a<!�a<Y�a<2�a<M�a<S�a<r�a<��a<��a<�a<ޠa<�a<�a<E�a<@�a<=�a<9�a<�a<ڠa<��a<i�a<�a<��a<��a<c�a<h�a<2�a<J�a<3�a<S�a<z�a<��a<џa<Οa<�a<��a<6�a<-�a<�a<�a<ğa<��a<[�a<E�a<�a<ɞa<��a<_�a<C�a<�a<#�a<�a<��a<��a<b�a<N�a<��a<͜a<]�a<�a<��a<��a<��a<�a<��a<�a<��a<c�a<��a<їa<q�a<X�a<(�a<#�a<�a<��a<��a<:�a<5�a<��a<h�a<�a<h�a<�a<O�a<�a<C�a<��a<"�a<��a<4�a<��a<`�a<��a<M�a<Սa<U�a<،a<4�a<��a<ϊa<:�a<y�a<��a<�a<2�a<��a<Ѕa<O�a<��a<K�a<ԃa<z�a<K�a<��a<�a<��a<r�a<6�a<��a<فa<n�a<6�a<��a<p�a<�a<�a<qa<�~a<�~a<N~a<~a<�}a<�}a<�}a<a}a<]}a<+}a<"}a<�|a<�|a<�|a<)|a<
|a<�{a<x{a<#{a<�za<�za<qza<�za<^za<�za<�za<�za<#{a<h{a<�{a<�  �  /|a<�|a<�|a<5}a<^}a<�}a<�}a<~a<-~a<Z~a<�~a<�~a<�~a<9a<a<�a<0�a<��a<�a<��a<��a<t�a<ւa<6�a<��a<�a<S�a<��a<҄a<�a<X�a<��a<�a<q�a<܆a<W�a< �a<��a<^�a<�a<܊a<��a<c�a<0�a<�a<��a<2�a<Ϗa<k�a<�a<w�a<�a<[�a<ݒa<e�a<�a<v�a<�a<��a<�a<��a<V�a<ݗa<e�a<˘a<5�a<��a<��a<,�a<U�a<�a<��a<��a<�a<�a<=�a<g�a<��a<�a<w�a<Ϝa<,�a<��a<�a<p�a<֞a<1�a<X�a<��a<��a<�a<�a<�a<	�a<�a<�a<$�a<6�a<W�a<g�a<��a<��a<ՠa<��a<�a<%�a<)�a<%�a<)�a<�a<ؠa<��a<n�a<2�a<��a<֟a<��a<y�a<X�a<]�a<g�a<��a<��a<��a<ӟa<�a<
�a<*�a<6�a<�a<��a<�a<ȟa<��a<S�a<�a<՞a<��a<y�a<E�a<�a<��a<ϝa<��a<��a<��a<h�a<,�a<�a<��a<q�a<�a<��a<�a<��a<$�a<��a<V�a<ߘa<x�a<�a<�a<��a<��a<N�a<-�a<�a<Жa<��a<n�a<�a<��a<F�a<۔a<[�a<Փa<@�a<��a<�a<��a<�a<��a<�a<��a<	�a<��a<:�a<��a<H�a<��a<#�a<��a< �a<J�a<��a<҈a<�a<Z�a<��a<	�a<o�a<Մa<b�a<�a<��a<b�a<�a<�a<��a<}�a<M�a<�a<��a<a�a<�a<��a<S�a<�a<�a<a<�~a<y~a<1~a<�}a<�}a<�}a<p}a<W}a<>}a<*}a<}a<�|a<�|a<�|a<W|a<|a<�{a<~{a<8{a<�za<�za<�za<�za<�za<�za<�za<{a<={a<�{a<�{a<�  �  a|a<�|a<�|a<}a<q}a<�}a<�}a<~a<~a<D~a<`~a<�~a<�~a<�~a<]a<�a<
�a<m�a<��a<h�a<сa<q�a<��a<h�a<��a<��a<R�a<��a<�a<%�a<��a<΅a<!�a<��a<�a<��a<�a<��a<m�a<D�a<�a<��a<��a<-�a<��a<�a<\�a<̏a<`�a<�a<G�a<ߑa<<�a<Βa<$�a<��a<G�a<��a<}�a<��a<��a<*�a<ʗa<\�a<��a<b�a<��a<��a<'�a<y�a<��a<��a<��a<��a<'�a<X�a<��a<��a<*�a<��a<�a<r�a<��a<1�a<��a<Оa<!�a<S�a<��a<��a<�a<ԟa<�a<�a<ޟa<��a<�a<�a<�a<8�a<m�a<��a< a<̠a<�a<�a<=�a<B�a<�a<�a<�a<נa<}�a<\�a<$�a<�a<��a<��a<��a<��a<��a<��a<��a<ޟa<ޟa<$�a<�a<,�a<�a<'�a<�a<ǟa<Ɵa<_�a<=�a<�a<��a<s�a<;�a<#�a<ܝa<ϝa<��a<��a<��a<^�a<f�a<
�a<�a<��a<Y�a<�a<��a<J�a<��a<h�a<ՙa<^�a<��a<��a<j�a<�a<Ǘa<��a<��a<C�a<�a<��a<��a<v�a<��a<וa<C�a<Дa<P�a<��a<1�a<��a<�a<O�a<ِa<X�a<��a<w�a<�a<��a<�a<��a<?�a<��a<P�a<~�a<�a<D�a<��a<�a<+�a<��a<Æa<"�a<��a<"�a<��a<!�a<Ńa<{�a<]�a<��a<؂a<��a<G�a<	�a<��a<��a<�a<��a<5�a<�a<oa<�~a<�~a<8~a<~a<�}a<�}a<w}a<K}a<D}a<}a<'}a<�|a<�|a<�|a<m|a<\|a<|a<�{a<�{a<c{a<({a<�za<�za<�za<�za<�za<�za<{a<`{a<�{a<�{a<�  �  e|a<�|a< }a<6}a<f}a<�}a<�}a<�}a<�}a<~a<)~a<h~a<�~a<�~a<a<na<�a<Y�a<��a<=�a<��a<I�a<��a<=�a<��a<�a<q�a<��a<	�a<X�a<��a<�a<j�a<ʆa<D�a<��a<a�a<��a<��a<[�a<�a<Ћa<��a<A�a<�a<��a<F�a<��a<L�a<��a<-�a<��a<�a<��a< �a<y�a<�a<��a<7�a<וa<q�a<�a<��a<A�a<��a<G�a<��a<�a<<�a<��a<��a<��a<
�a<@�a<n�a<��a<Λa<�a<n�a<˜a<)�a<}�a<ߝa<>�a<��a<�a<7�a<^�a<��a<��a<��a<��a<��a<��a<ɟa<��a<��a<ɟa<�a<�a<8�a<T�a<��a<��a<�a<�a<�a<2�a<0�a<+�a<��a<ܠa<��a<�a<P�a<'�a<��a<�a<��a<Οa<��a<ܟa<�a<��a<
�a<'�a<1�a<F�a<6�a<�a<�a<��a<��a<J�a<�a<��a<��a<I�a<�a<ӝa<��a<��a<��a<j�a<_�a<C�a<=�a< �a<�a<��a<v�a<%�a<��a<R�a<�a<w�a<�a<��a<9�a<��a<��a<K�a<	�a<ؗa<��a<k�a<1�a<�a<��a<��a<�a<��a<)�a<��a<)�a<��a<��a<W�a<Ƒa<+�a<��a<�a<��a<1�a<Ȏa<Z�a<�a<��a<$�a<��a<5�a<��a<�a<Z�a<��a<�a<V�a<��a<	�a<i�a<Յa<=�a<Ȅa<d�a<�a<��a<g�a<$�a<�a<��a<f�a<�a<��a<o�a<�a<��a<�a<�a<4a<�~a<m~a<~a<�}a<�}a<e}a<B}a<}a<}a<�|a<�|a<�|a<�|a<�|a<�|a<s|a<*|a<�{a<�{a<�{a<T{a<-{a<{a<{a<�za<{a<!{a<^{a<�{a<�{a<|a<�  �  u|a<�|a<�|a<,}a<X}a<{}a<�}a<�}a<�}a<�}a<~a<#~a<J~a<�~a<�~a<Oa<�a<�a<��a<�a<��a<�a<��a< �a<��a<�a<p�a<ڄa<�a<��a<مa<9�a<��a<�a<��a<�a<��a<�a<��a<��a<X�a<��a<��a<l�a<�a<��a<&�a<��a<+�a<��a<�a<n�a<�a<D�a<Ӓa<E�a<ѓa<v�a<�a<��a<<�a<��a<v�a<�a<��a<)�a<��a<��a<b�a<��a<˚a<!�a<7�a<|�a<��a<�a<�a<W�a<��a<�a<Y�a<��a< �a<P�a<��a<��a<+�a<Y�a<{�a<��a<��a<��a<��a<�a<��a<i�a<��a<��a<��a<Οa<�a<0�a<c�a<��a<��a<��a<�a<�a<%�a<�a<�a<�a<ՠa<��a<w�a<]�a<�a<0�a<��a<�a<�a<�a<�a</�a<@�a<7�a<S�a<:�a<,�a<�a<�a<��a<e�a<7�a<�a<��a<I�a< �a<�a<��a<��a<L�a<Z�a<9�a<@�a<+�a<�a<	�a<՜a<��a<i�a<$�a<ۛa<d�a<"�a<��a<@�a<ʙa<t�a<!�a<Ƙa<��a<'�a<�a<ŗa<��a<V�a<�a<�a<|�a<�a<��a<+�a<��a<�a<}�a<��a<.�a<|�a<��a<c�a<�a<z�a<�a<��a<%�a<ލa<X�a<�a<��a<�a<��a<�a<��a<Չa<�a<��a<ԇa<E�a<��a<�a<��a<�a<��a<0�a<�a<��a<f�a<��a<a<q�a<�a<��a<Q�a<�a<p�a<�a<�a< a<�~a<~a<�}a<�}a<`}a<$}a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<d|a<M|a<|a<�{a<�{a<{{a<b{a<,{a<J{a<#{a<W{a<O{a<�{a<�{a<|a<G|a<�  �  �|a<�|a<}a<7}a<c}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<~a<a~a<�~a<a<`a<�a<^�a<�a<o�a<�a<��a</�a<��a<�a<t�a<�a<O�a<��a<
�a<]�a<ӆa<B�a<��a<8�a<̈a<l�a<#�a<��a<r�a<�a<ьa<\�a<�a<��a<1�a<��a<�a<v�a<ސa<B�a<��a<#�a<��a<�a<��a<3�a<ϔa<s�a<�a<��a<[�a<�a<��a<1�a<��a<�a<V�a<��a<��a<8�a<i�a<��a<֛a<�a<G�a<��a<ݜa<6�a<��a<��a<+�a<��a<Ҟa<��a<J�a<d�a<��a<t�a<��a<l�a<f�a<T�a<V�a<H�a<S�a<L�a<x�a<��a<ϟa<�a<5�a<k�a<��a<נa<�a<)�a<.�a<7�a<�a<�a<�a<ՠa<��a<��a<m�a<O�a<4�a<2�a<;�a<J�a<;�a<V�a<U�a<n�a<Q�a<K�a<8�a<�a<�a<��a<U�a<��a<��a<n�a<$�a<Нa<��a<W�a<O�a<&�a<�a<�a<�a<��a<��a<�a<�a<��a<��a<)�a<�a<��a<-�a<֚a<c�a<�a<��a<I�a<��a<��a<v�a<I�a<��a<×a<{�a<>�a<іa<��a<�a<��a<�a<��a<ޓa<<�a<��a<��a<[�a<��a<&�a<��a<7�a<Ȏa<c�a<��a<��a<=�a<�a<}�a<�a<��a<%�a<t�a<��a<M�a<��a<�a<s�a<цa<:�a<��a<6�a<Ԅa<x�a<�a<ʃa<q�a<,�a<ނa<q�a<1�a<��a<Z�a<ʀa<[�a<�a<Ua<�~a<n~a<�}a<�}a<G}a<}a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<|a<F|a<;|a<�{a<�{a<�{a<�{a<z{a<i{a<`{a<v{a<�{a<�{a<�{a<+|a<\|a<�  �  �|a<�|a<5}a<>}a<?}a<i}a<p}a<�}a<t}a<�}a<�}a<�}a<�}a<'~a<z~a<�~a<'a<�a<7�a<ŀa<K�a<�a<v�a<�a<{�a<1�a<��a<�a<|�a<��a<=�a<��a<�a<h�a<�a<|�a<�a<��a<:�a<��a<��a<;�a<��a<g�a<>�a<��a<�a<��a<�a<g�a<��a<5�a<r�a<ڑa<N�a<�a<r�a<�a<��a<+�a<��a<��a<I�a<��a<~�a<%�a<��a<9�a<e�a<ߚa<�a<U�a<��a<ța<�a<,�a<��a<ɜa<�a<u�a<��a<�a<F�a<��a<�a<�a<_�a<?�a<u�a<_�a<y�a<M�a<?�a<9�a<�a<
�a<�a<6�a<H�a<W�a<��a<ȟa<"�a<8�a<��a<àa<�a<	�a<-�a<e�a<�a<G�a<�a<��a<ߠa<��a<��a<y�a<��a<c�a<e�a<n�a<t�a<��a<j�a<��a<X�a<{�a<?�a<��a<ϟa<��a<P�a<Оa<��a<4�a<؝a<��a<g�a<@�a<�a<�a<ܜa<�a<�a<؜a<��a<̜a<Ϝa<��a<��a<R�a<��a<śa<F�a<�a<��a<I�a<יa<��a<A�a<ژa<��a<`�a<5�a<�a<��a<e�a<ܖa<��a<
�a<��a<��a<u�a<ϓa<�a<��a<��a<�a<y�a<�a<��a<�a<��a<�a<�a<r�a<*�a<܌a<e�a<�a<��a<B�a<��a<�a<m�a<ˈa<D�a<��a<�a<_�a<��a<y�a<��a<��a<B�a<�a<��a<W�a<�a<��a<G�a<��a<K�a<��a<R�a<�a<.a<�~a<*~a<�}a<b}a<1}a<�|a<�|a<�|a<�|a<�|a<|a<�|a<�|a<�|a<�|a<�|a<�|a<O|a<d|a<|a<|a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<|a<W|a<q|a<�  �  �|a<�|a<}a<1}a<b}a<h}a<`}a<e}a<j}a<l}a<�}a<�}a<�}a<�}a<0~a<�~a<a<�a<�a<��a<:�a<Ёa<o�a<�a<��a<�a<��a<�a<��a<�a<O�a<��a<!�a<��a<$�a<��a<4�a<ŉa<\�a<�a<��a<V�a<��a<��a<�a<��a<)�a<��a<�a<?�a<��a<�a<]�a<ˑa<4�a<��a<&�a<̓a<r�a<�a<��a<|�a<+�a<ڗa<��a<$�a<��a<�a<x�a<�a<0�a<�a<��a<�a<*�a<q�a<��a<��a<B�a<��a<ϝa<(�a<w�a<��a<�a<�a<7�a<[�a<l�a<_�a<I�a<9�a<$�a<�a<�a<�a<�a<�a<�a<=�a<}�a<��a<�a<+�a<n�a<��a<�a<&�a<)�a<6�a<B�a<J�a<.�a<�a<��a<٠a<Ǡa<��a<��a<��a<��a<��a<��a<��a<��a<��a<{�a<V�a<1�a<�a<ϟa<r�a<�a<Şa<e�a<�a<˝a<u�a<2�a<��a<��a<ɜa<Мa<��a<��a<ǜa<Ĝa<Ɯa<Ȝa<��a<s�a<D�a<	�a<ɛa<v�a<�a<��a<^�a<�a<��a<i�a<�a<Ϙa<��a<L�a<�a<��a<l�a<��a<��a<�a<��a<�a<Y�a<��a<��a<C�a<��a<�a<_�a<��a<7�a<Ўa<k�a<�a<��a<`�a<�a<��a<k�a<�a<��a<�a<��a<�a<��a<��a<V�a<��a<&�a<��a<#�a<��a<8�a<Ǆa<b�a<�a<��a<_�a<��a<��a<�a<��a<C�a<��a<!�a<�a<a<�~a<~a<�}a<D}a<�|a<�|a<�|a<�|a<n|a<e|a<q|a<}|a<�|a<�|a<�|a<�|a<~|a<r|a<f|a<=|a<%|a<|a<�{a<�{a<�{a<�{a<�{a<�{a<|a<@|a<o|a<�|a<�  �  �|a<}a<}a<K}a<]}a<A}a<]}a<D}a<k}a<P}a<i}a<t}a<�}a<�}a<~a<�~a<�~a<`a<�a<��a<2�a<��a<r�a<�a<��a<&�a<��a<'�a<��a<�a<Y�a<�a<Y�a<·a<=�a<��a<_�a<�a<��a<"�a<ċa<r�a<��a<��a<�a<��a<�a<v�a<ڏa<&�a<��a<ʐa<D�a<��a<�a<��a<	�a<��a<7�a<��a<��a<{�a<�a<ȗa<q�a<��a<��a<�a<��a<�a<J�a<��a<ța<?�a<O�a<��a<Ϝa<�a<r�a<��a<�a<5�a<��a<��a<�a<7�a<K�a<y�a<;�a<]�a<2�a<)�a<�a<�a<Ӟa<��a<ڞa<��a<��a<�a<C�a<��a<şa<1�a<O�a<��a<Ѡa<�a<I�a<@�a<d�a<@�a<O�a<'�a<#�a<*�a<�a<ݠa< a< a<��a<֠a< a<��a<��a<��a<��a<c�a<L�a<�a<��a<o�a<��a<ƞa<I�a<��a<��a<B�a<�a<Μa<Мa<��a<��a<��a<��a<��a<��a<ɜa<��a<��a<��a<]�a<(�a<̛a<��a<%�a<�a<��a<=�a<ڙa<��a<H�a<�a<ۘa<`�a<�a<ӗa<l�a<!�a<��a<5�a<�a<�a<J�a<��a<��a<�a<��a<Őa</�a<��a<�a<��a<0�a<�a<��a<_�a<�a<��a<X�a<�a<��a<%�a<��a<%�a<��a<�a<f�a<	�a<J�a<҆a<=�a<ąa<i�a<��a<��a<�a<Ճa<g�a<�a<��a<3�a<ցa<�a<��a<�a<�a<a<f~a<�}a<e}a</}a<�|a<�|a<]|a<M|a<W|a<G|a<w|a<^|a<�|a<�|a<�|a<�|a<�|a<�|a<]|a<]|a<-|a<&|a</|a<�{a<�{a<�{a<|a<|a<X|a<k|a<w|a<�|a<�  �  �|a<	}a<)}a<8}a<G}a<S}a<b}a<D}a<@}a<I}a<[}a<b}a<}a<�}a<~a<g~a<�~a<Qa<�a<v�a<�a<��a<y�a<�a<��a<�a<��a<"�a<��a<�a<�a<�a<Q�a<·a<X�a<�a<d�a<�a<��a<:�a<�a<��a<�a<��a<"�a<��a<�a<��a<܏a< �a<|�a<Ԑa<0�a<��a<�a<s�a<��a<��a</�a<�a<��a<U�a<�a<̗a<�a<�a<��a<�a<��a<��a<_�a<��a<�a< �a<Y�a<��a<��a<:�a<p�a<��a<�a<Y�a<��a<�a<�a<3�a<D�a<X�a<R�a<f�a<7�a<�a<��a<�a<Ȟa<��a<��a<��a<�a<��a<7�a<��a<ßa<�a<P�a<��a<�a<
�a<3�a<M�a<Z�a<f�a<g�a<E�a<*�a<�a<�a<�a<�a<Ҡa<��a<��a<àa<Ơa<Πa<��a<��a<o�a<9�a<��a<��a<t�a<��a<��a<B�a<�a<��a<4�a<�a<˜a<��a<��a<��a<��a<��a<��a<��a<Ϝa<��a<��a<�a<]�a<"�a<��a<��a<K�a<�a<��a<=�a<��a<��a<M�a<��a<��a<x�a<3�a<�a<��a<�a<��a<�a<��a<��a<M�a<��a<ڒa<&�a<v�a<��a<�a<��a<�a<��a<)�a<܍a<��a<9�a<�a<��a<e�a<��a<��a<%�a<��a<2�a<��a<�a<��a<�a<T�a<ӆa<k�a<�a<g�a<��a<��a<D�a<�a<��a<�a<��a<,�a<��a<(�a<��a<�a<oa<�~a<k~a<�}a<f}a<}a<�|a<�|a<M|a<A|a<E|a<F|a<L|a<_|a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<v|a<L|a<-|a<
|a<�{a<|a<|a<|a<|a<9|a<m|a<�|a<�|a<�  �  b~a<q~a<�~a<�~a<�~a<�~a<�~a<a<a< a<a<5a<va<�a<�a<;�a<��a<�a<��a<!�a<ւa<h�a<ʃa<��a<�a<��a<�a<v�a<��a<g�a<�a<^�a<�a<A�a<Éa<R�a<��a<|�a<�a<��a<2�a<��a<G�a<ώa<a�a<ڏa<c�a<��a<%�a<��a<ۑa<M�a<��a<��a<��a<�a<o�a<�a<��a<M�a<��a<��a<r�a<��a<{�a<0�a<��a<�a<��a<�a<C�a<��a<�a<<�a<��a<��a<�a<L�a<��a<��a<!�a<c�a<��a<џa<��a<+�a<K�a<k�a<��a<S�a<v�a<z�a<@�a<7�a<'�a<,�a<+�a<2�a<I�a<��a<��a<Рa<�a<R�a<��a<��a<��a<=�a<E�a<^�a<T�a<f�a<U�a<k�a<L�a<I�a</�a<�a<�a<�a<��a< �a<�a<�a<ơa<��a<��a<�a<S�a<1�a<�a<~�a<g�a<��a<��a<A�a<��a<˞a<o�a<J�a<$�a<�a<��a<��a<�a<	�a<�a<ȝa<�a<ŝa<��a<h�a<$�a<�a<��a<d�a<�a<כa<g�a<�a<Қa<b�a<E�a<�a<��a<K�a<Ԙa<��a<�a<��a<0�a<��a<�a<|�a<��a<)�a<��a<ܒa<3�a<��a<�a<��a<.�a<��a<[�a<
�a<��a<�a<
�a<��a<W�a<܌a<g�a<�a<i�a<�a<m�a<҉a<X�a<�a<9�a<·a<U�a<نa<��a<�a<��a<=�a<ׄa<h�a<�a<��a<*�a<��a<�a<��a<@�a<��a<�a<�a<Ga<�~a<�~a<W~a<G~a<~a<�}a<
~a<~a<2~a<~a<~a<0~a<~a<~a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<(~a<6~a<�  �  e~a<�~a<�~a<�~a<�~a<�~a<�~a<�~a<�~a<a<:a<Ga<la<�a<�a<N�a<��a<5�a<��a<2�a<��a<?�a<�a<r�a<�a<��a<�a<��a<��a<o�a<�a<I�a<��a<1�a<��a<6�a<Ċa<E�a<�a<��a<(�a<��a<V�a<�a<e�a<�a<G�a<��a<�a<j�a<��a<P�a<Ēa<�a<��a<�a<��a<�a<��a<n�a<�a<��a<0�a<�a<��a<�a<��a<$�a<��a< �a<L�a<��a<�a<*�a<[�a<��a<�a<8�a<{�a<��a<�a<^�a<��a<ݟa<�a<5�a<S�a<k�a<i�a<r�a<U�a<K�a<L�a<L�a<F�a<)�a<:�a<O�a<j�a<~�a<��a<��a<(�a<P�a<|�a<ʡa<��a<"�a<R�a<g�a<s�a<p�a<b�a<]�a<>�a<)�a<�a<�a<��a<�a<�a<ءa<ڡa<ޡa<Сa<��a<��a<��a<_�a<�a<ܠa<��a</�a<�a<��a<i�a<�a<��a<��a<b�a<8�a<�a<�a<�a<��a<�a<ڝa<�a<ϝa<��a<��a<n�a<>�a<��a<��a<`�a<�a<��a<V�a<
�a<��a<k�a<�a<әa<��a<A�a<�a<��a<(�a<��a<?�a<��a<�a<s�a<��a<.�a<��a<�a<H�a<��a<;�a<��a<7�a<��a<{�a<�a<��a<>�a<��a<��a<>�a<�a<m�a<��a<}�a<�a<g�a<ԉa<E�a<��a<:�a<��a<A�a<̆a<S�a<�a<��a<A�a<�a<��a<�a<��a<*�a<��a<+�a<��a<�a<��a<3�a<�a<Da<�~a<�~a<x~a<<~a<%~a<'~a<~a< ~a<�}a<~a<~a<~a<#~a<~a<~a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<~a<@~a<�  �  H~a<�~a<�~a<�~a<�~a<�~a<a<�~a<$a<a<a<Ka<ma<�a<�a<\�a<��a<8�a<��a<;�a<߂a<_�a<�a<j�a<�a<��a<��a<��a<�a<[�a<҇a<O�a<��a<:�a<��a<�a<ۊa<B�a<�a<��a<�a<��a<=�a<Վa<N�a<�a<C�a<ːa<B�a<��a<�a<0�a<��a<"�a<��a<�a<��a<"�a<��a<f�a<�a<ėa<Q�a<�a<��a<�a<��a<�a<��a<�a<=�a<��a<��a</�a<Y�a<ĝa<۝a<+�a<��a<��a<�a<N�a<��a<ğa<�a<)�a<K�a<u�a<^�a<��a<v�a<q�a<\�a<+�a<J�a<2�a<D�a<D�a<r�a<�a<��a<�a<�a<��a<��a<��a<�a<!�a<P�a<Q�a<n�a<S�a<Z�a<E�a<:�a<,�a<�a<�a<סa<�a<�a<ۡa<סa<ˡa<ơa<��a<��a<w�a<[�a<�a<۠a<��a<P�a<�a<��a<O�a<�a<a<��a<W�a<F�a<�a<�a<�a<�a<�a<��a<
�a<ȝa<ǝa<��a<]�a<4�a<ٜa<��a<P�a<	�a<��a<_�a<��a<��a<��a<�a<ԙa<��a<)�a<Ԙa<x�a<�a<��a<?�a<��a<$�a<��a<ߔa<]�a<w�a<��a<Z�a<��a<9�a<��a<;�a<Ώa<t�a<�a<ώa<_�a<�a<��a<6�a<�a<^�a<�a<i�a<ۊa<Q�a<͉a<J�a<��a<L�a<��a<4�a<چa<U�a<�a<��a<-�a<˄a<v�a<�a<��a<4�a<��a<H�a<��a<7�a<��a<�a<�a<Ma< a<�~a<�~a<=~a</~a<~a<�}a<6~a<~a<=~a<~a<~a<!~a<~a<	~a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<o}a<�}a<�}a<�}a<�}a<
~a<6~a<�  �  T~a<}~a<�~a<�~a<�~a<�~a<�~a<a<a<&a<Da<ya<�a<�a<�a<��a<�a<]�a<ǁa<H�a<؂a<n�a<��a<��a<�a<�a<�a<{�a<�a<T�a<ća<�a<��a<�a<��a<�a<��a<-�a<��a<h�a<
�a<��a<:�a<܎a<b�a<Ϗa<k�a<��a<2�a<��a<�a<m�a<Вa<K�a<��a<*�a<��a<Q�a<�a<��a< �a<��a<_�a<�a<y�a<9�a<��a<#�a<��a<�a<>�a<��a<˜a<��a<M�a<t�a<ҝa<�a<>�a<��a<�a<<�a<��a<ɟa<��a<9�a<J�a<f�a<��a<e�a<��a<o�a<_�a<]�a<j�a<g�a<m�a<j�a<��a<��a<�a<�a<;�a<t�a<��a<סa<��a<<�a<;�a<c�a<d�a<[�a<R�a<?�a<�a<�a<�a<֡a<ޡa<��a<��a<��a<��a<ša<��a<��a<��a<��a<G�a<,�a<�a<��a<d�a<�a<��a<t�a<=�a<��a<��a<}�a<k�a<R�a<>�a<�a<�a<�a<	�a<ߝa<�a<��a<��a<o�a<*�a<�a<��a<A�a<֛a<��a<�a<��a<��a<2�a<��a<��a<j�a<#�a<јa<u�a<#�a<��a<$�a<Öa<�a<��a<�a<Q�a<��a<�a<��a<�a<Q�a<ѐa<i�a<��a<��a<+�a<Ǝa<l�a<�a<��a<`�a<Ќa<m�a<��a<a�a<܊a<M�a<��a<�a<��a<��a<��a<�a<��a<F�a<҅a<��a<*�a<Єa<j�a<�a<��a<%�a<��a<�a<��a<6�a<��a<D�a<�a<�a<*a<�~a<�~a<s~a<Z~a<2~a<'~a<$~a<'~a<~a<~a<0~a<~a<~a<�}a<�}a<�}a<�}a<�}a<u}a<^}a<\}a<v}a<p}a<w}a<�}a<�}a<~a<-~a<�  �  D~a<L~a<�~a<�~a<�~a<�~a<�~a<,a< a<aa<ca<|a<�a<�a<E�a<��a<�a<\�a<�a<z�a<�a<��a<��a<��a<��a<��a<��a<N�a<نa<(�a<��a<��a<��a<�a<j�a<��a<k�a<2�a<��a<O�a<��a<��a<'�a<��a<c�a<a<x�a<ǐa<R�a<��a<�a<��a<�a<Q�a<Γa<P�a<ڔa<c�a<��a<��a<S�a<җa<t�a<#�a<��a<M�a<��a<&�a<m�a<̛a<�a<]�a<��a<ڜa<L�a<\�a<��a<�a<3�a<��a<��a<.�a<X�a<��a<ԟa<�a<O�a<V�a<��a<z�a<��a<~�a<��a<��a<g�a<q�a<��a<��a<��a<Ša<�a< �a<t�a<��a<̡a<�a<�a<<�a</�a<^�a<2�a<K�a<"�a<!�a<�a<��a<�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<k�a<��a<D�a<)�a<��a<��a<��a<�a<��a<��a<A�a<�a<՞a<��a<��a<[�a<>�a<I�a<A�a<�a<)�a<��a<��a<��a<��a<\�a<��a<Мa<e�a<0�a<��a<��a<�a<��a<w�a<�a<��a<��a<Q�a<��a<��a<b�a<��a<��a<�a<Жa< �a<��a<�a<]�a<�a<!�a<��a<��a<w�a<��a<{�a<�a<��a<^�a<ގa<��a<6�a<��a<t�a<Ča<p�a<ϋa<I�a<��a< �a<��a<��a<��a<�a<z�a<��a<��a<?�a<��a<v�a<��a<��a<A�a<��a<��a<�a<؂a<3�a<ށa<D�a<�a<v�a<�a<�a<?a<�~a<�~a<�~a<_~a<M~a<a~a<0~a<F~a<3~a</~a<0~a< ~a<~a<�}a<�}a<�}a<�}a<q}a<e}a<g}a<:}a<S}a<L}a<{}a<�}a<�}a<�}a<�}a<�  �  5~a<]~a<�~a<�~a<�~a<�~a<a<&a<]a<Xa<ua<�a<�a<$�a<P�a<Ȁa<*�a<��a<�a<��a<�a<��a<�a<��a<�a<~�a<�a<^�a<Æa<�a<��a<�a<H�a<Ոa<?�a<��a<g�a<ڊa<x�a<�a<͌a<v�a<%�a<��a<E�a<ۏa<[�a<�a<Z�a<Ǒa<P�a<��a<�a<��a<��a<v�a<��a<��a<5�a<ʖa<8�a<�a<��a<(�a<��a<&�a<��a<�a<i�a<̛a<�a<K�a<��a<��a<�a<U�a<x�a<ĝa<$�a<P�a<��a<�a<F�a<��a<�a<�a<C�a<e�a<}�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ڠa<��a<1�a<@�a<`�a<��a<̡a<��a<�a<4�a<D�a<C�a<@�a<@�a<�a<�a<ءa<��a<��a<��a<t�a<��a<x�a<p�a<v�a<��a<|�a<��a<|�a<g�a<P�a<'�a<��a<��a<{�a<U�a<�a<��a<��a<6�a<�a<��a<��a<��a<��a<J�a<W�a<D�a< �a<�a<�a<��a<��a<H�a<�a<��a<U�a<�a<��a<:�a<��a<��a<6�a<�a<��a<`�a<!�a<�a<��a<`�a<��a<��a<1�a<��a<<�a<��a<�a<��a<ɓa<Y�a<̒a</�a<��a<�a<��a<G�a<؏a<D�a<�a<��a<;�a<̍a<M�a<܌a<V�a<ˋa<I�a<��a<�a<r�a<Ոa<A�a<݇a<>�a<͆a<u�a<�a<��a<J�a<�a<��a<P�a<�a<��a<$�a<��a<Q�a<؁a<j�a<�a<k�a<0�a<�a<oa<	a<�~a<�~a<�~a<n~a<L~a<o~a<F~a<C~a<:~a<'~a<~a<�}a<�}a<�}a<�}a<u}a<H}a<+}a<}a<)}a<}a<3}a<C}a<]}a<�}a<�}a<�}a<�  �  �}a<^~a<y~a<�~a<�~a<a<9a<,a<va<ya<�a<�a<�a<_�a<��a<�a<*�a<ˁa<!�a<��a<(�a<��a<9�a<��a<�a<r�a<�a<P�a<��a<�a<I�a<Շa<�a<��a<"�a<��a<9�a<��a<u�a<�a<a<N�a<�a<��a</�a<�a<V�a<��a<i�a<ˑa<s�a<��a<N�a<��a<*�a<��a<+�a<a<.�a<��a<^�a<2�a<��a<.�a<Йa<"�a<��a<��a<v�a<��a<�a<J�a<J�a<��a<��a<�a<O�a<��a<�a<�a<��a<Þa<M�a<g�a<˟a<�a<2�a<{�a<{�a<��a<��a<��a<Ѡa<��a<ڠa<��a<�a<ܠa<�a<�a<<�a<}�a<��a<ۡa<ѡa<�a<+�a<5�a<K�a<0�a<G�a<�a<�a<�a<��a<��a<`�a<��a<L�a<h�a<2�a<[�a<Z�a<W�a<t�a<Q�a<|�a<X�a<O�a</�a<�a<�a<��a<n�a<�a<�a<��a<H�a<@�a<�a<�a<��a<��a<x�a<u�a<[�a<)�a<7�a<�a<ѝa<��a<G�a<��a<��a<W�a<Ǜa<��a<�a<��a<v�a<�a<ߙa<d�a<\�a<�a<ۘa<y�a</�a<�a<�a<?�a<��a<T�a<��a<�a<��a<�a<��a<ʒa<Y�a<ґa<J�a<ڐa<@�a<	�a<i�a<=�a<��a<A�a<�a<I�a<�a<>�a<׋a< �a<��a<�a<7�a<ӈa<�a<��a<�a<��a<7�a<��a<��a<�a<�a<n�a<8�a<�a<|�a<;�a<��a<v�a<�a<|�a<%�a<��a<X�a<�a<�a<>a< a<�~a<�~a<�~a<p~a<�~a<K~a<e~a<F~a<(~a<~a<�}a<�}a<�}a<�}a<S}a<'}a< }a<�|a<}a<�|a<}a<�|a<H}a<m}a<�}a<�}a<�  �  �}a<6~a<r~a<�~a<�~a<a<<a<ia<za<�a<�a<�a<8�a<z�a<��a<%�a<n�a<Ձa<H�a<ʂa<A�a<Ƀa<.�a<��a<�a<s�a<؅a<2�a<��a<��a<#�a<��a<�a<v�a<�a<Y�a<�a<��a<K�a<Ƌa<��a<@�a<�a<��a<3�a<ԏa<j�a<��a<��a<��a<j�a<�a<T�a<Ɠa<e�a<Δa<R�a<��a<g�a<��a<��a<-�a<Ęa<S�a<Ùa<:�a<��a<��a<V�a<��a<؛a<*�a<&�a<��a<��a<�a<�a<n�a<��a<�a<g�a<��a<*�a<c�a<��a<�a<6�a<o�a<��a<��a<ڠa<ڠa<�a<ݠa<�a<�a<�a<�a<,�a<U�a<c�a<��a<��a<ۡa<�a<&�a</�a<>�a<:�a<,�a< �a<��a<�a<��a<��a<��a<\�a<H�a<�a<,�a<%�a<?�a<�a<6�a<[�a<K�a<U�a<P�a<D�a<3�a<�a<�a<��a<r�a<B�a<��a<��a<��a<[�a<�a<�a<֞a<��a<��a<��a<t�a<d�a<-�a<��a<ȝa<��a<9�a<�a<|�a<9�a<��a<R�a<�a<��a<B�a<ؙa<��a<m�a<2�a<Șa<��a<k�a<'�a<ߗa<��a<)�a<a<L�a<ܕa<O�a<��a<1�a<��a<��a<��a<��a<q�a<�a<y�a<�a<��a<8�a<юa<f�a<ߍa<a�a<ڌa<B�a<��a<�a<v�a<�a<�a<��a<�a<s�a<��a<w�a<�a<��a<X�a<�a<τa<j�a<%�a<ڃa<�a<.�a<˂a<i�a<�a<��a<5�a<Āa<^�a<�a<�a<fa<9a<a<�~a<�~a<�~a<�~a<�~a<n~a<J~a<2~a<~a<�}a<�}a<�}a<h}a<3}a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<+}a<3}a<v}a<�}a<�  �  �}a<~a<|~a<�~a<�~a<&a<,a<{a<�a<�a<�a<4�a<h�a<��a<��a<3�a<��a<
�a<s�a<�a<K�a<ԃa<$�a<��a<��a<��a<Ʌa<%�a<��a<��a<:�a<r�a<чa<A�a<��a<H�a<Ӊa<e�a< �a<ԋa<x�a<�a<�a<z�a<W�a<��a<z�a<��a<x�a<�a<}�a<�a<k�a<�a<q�a<��a<��a<�a<��a<�a<ϗa<A�a<Ԙa<O�a<ʙa<Q�a<��a< �a<5�a<��a<��a<�a<=�a<D�a<��a<��a<�a<D�a<��a<ڝa<4�a<��a<�a<V�a<��a<�a<M�a<U�a<��a<��a<ߠa<�a<��a<	�a<�a<>�a<�a<H�a<S�a<v�a<��a<��a<�a<�a<!�a<�a<F�a<?�a<4�a<C�a<�a<�a<��a<��a<��a<C�a<*�a<�a<�a<��a<��a<��a<�a<9�a<!�a<P�a<>�a<Z�a<C�a<*�a<'�a<٠a<Рa<~�a<i�a<�a<��a<��a<y�a<\�a<�a<$�a<�a<ʞa<��a<~�a<o�a<"�a<�a<��a<��a<*�a<Ӝa<y�a<��a<��a<,�a<Úa<f�a<�a<Ǚa<y�a<.�a<�a<֘a<��a<H�a<)�a<��a<��a<�a<Җa<V�a<ϕa<d�a<˔a<^�a<��a<S�a<��a<&�a<��a<�a<Ӑa<)�a<ڏa<L�a<�a<a�a<�a<x�a<Ìa<j�a<��a<�a<X�a<��a<*�a<_�a<χa<F�a<ʆa<N�a<ޅa<y�a<%�a<��a<��a<\�a<�a<��a<��a<�a<�a<f�a<�a<��a<I�a<��a<��a<Y�a<�a<�a<aa<4a<a<�~a<�~a<�~a<�~a<^~a<a~a<3~a<~a<�}a<�}a<�}a<7}a<'}a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<%}a<x}a<�}a<�  �  �}a<~a<_~a<�~a<�~a<.a<[a<�a<�a<�a<�a<@�a<f�a<��a<�a<T�a<��a<�a<��a<�a<v�a<�a<U�a<��a<�a<~�a<��a<�a<a�a<��a<�a<X�a<ʇa<0�a<��a<�a<��a<[�a<�a<��a<N�a<�a<̍a<d�a<;�a<яa<t�a<�a<��a<,�a<��a<%�a<��a< �a<�a< �a<��a<�a<a<;�a<ޗa<o�a<��a<k�a<�a<M�a<��a<	�a<�a<y�a<��a<ӛa<	�a<A�a<u�a<��a<ٜa<�a<|�a<ԝa<�a<��a<ߞa<8�a<��a<͟a<E�a<c�a<��a<ܠa<�a<�a<�a<#�a<!�a<6�a<=�a<k�a<v�a<x�a<��a<ɡa< �a<�a<6�a<E�a<U�a<;�a<>�a<&�a<�a<�a<��a<�a<W�a<B�a<�a<��a<ݠa<�a<�a<�a<�a<��a<�a<4�a<-�a<=�a<I�a<+�a</�a<�a<�a<��a<��a<5�a<�a<��a<��a<��a<>�a<�a<��a<�a<͞a<��a<�a<T�a<�a<��a<��a<�a<��a<Y�a<�a<��a<�a<��a<U�a<�a<��a<d�a<$�a<�a<��a<g�a<7�a<�a<��a<��a<&�a<͖a<w�a<��a<�a<��a<l�a<ϓa<W�a<��a<G�a<Ǒa<-�a<Ԑa<I�a<�a<z�a<�a<~�a<�a<t�a<ьa<S�a<�a<��a<E�a<��a<��a<\�a<Ňa<4�a<��a<(�a<ͅa<r�a<�a<̄a<��a<?�a<��a<��a<��a<"�a<�a<��a<,�a<сa<q�a<
�a<��a<Q�a<�a<�a<�a<6a<'a<�~a<�~a<�~a<�~a<�~a<p~a</~a<~a<�}a<�}a<n}a<+}a<�|a<�|a<�|a<�|a<�|a<u|a<�|a<�|a<�|a<}a<>}a<�}a<�  �  �}a<7~a<T~a<�~a<�~a<a<ha<a<�a<�a<-�a<_�a<��a<�a<�a<��a<ցa<H�a<��a<�a<}�a<݃a<[�a<��a<�a<\�a<��a<(�a<O�a<Æa<Ԇa<9�a<��a<��a<��a<��a<��a<'�a<�a<k�a<P�a<�a<Ǎa<��a<�a<�a<r�a<�a<��a<)�a<��a<8�a<ɓa<+�a<̔a<3�a<��a<g�a<̖a<r�a<�a<r�a<�a<u�a<�a<A�a<��a<ޚa<G�a<z�a<��a<ڛa<Λa<$�a<D�a<}�a<��a<�a<I�a<��a<�a<I�a<�a<)�a<��a<�a<�a<|�a<��a<٠a<�a<�a<"�a<?�a<R�a<Q�a<��a<i�a<��a<��a<ˡa<��a<�a< �a<(�a<O�a<C�a<G�a<?�a<�a<�a<ԡa<��a<n�a<,�a<�a<�a<ܠa<��a<Ġa<��a<Ƞa<ʠa<�a<$�a< �a<V�a<2�a<>�a<=�a<�a<�a<Ԡa<��a<��a<\�a<$�a<��a<ǟa<y�a<��a<>�a<*�a< �a<Ҟa<��a<y�a<Z�a<�a<ԝa<k�a<�a<֜a<G�a< �a<Q�a<�a<��a<!�a<ۙa<v�a<8�a<�a<͘a<m�a<i�a<6�a<�a<֗a<c�a<;�a<ʖa<i�a<�a<|�a<��a<�a<�a<c�a<��a<Z�a<ґa<�a<ސa<��a<��a<}�a< �a<��a<�a<h�a<�a<(�a<��a<��a<:�a<��a<��a<@�a<��a<�a<��a<�a<��a<L�a<��a<��a<��a<0�a<�a<��a<f�a<;�a<ӂa<��a<,�a<Ձa<v�a<%�a<рa<k�a<G�a<�a<�a<{a<>a<%a<�~a<�~a<�~a<�~a<^~a<;~a<~a<�}a<�}a<]}a<5}a<�|a<�|a<�|a<a|a<b|a<N|a<s|a<}|a<�|a<�|a<#}a<�}a<�  �  �}a<~a<W~a<�~a<�~a<3a<pa<�a<�a<�a<.�a<[�a<��a<�a<7�a<��a<فa<E�a<��a<$�a<��a<��a<a�a<��a<�a<^�a<��a<��a<1�a<��a<�a<M�a<��a<��a<��a< �a<��a<�a<�a<��a<:�a<�a<��a<u�a<�a<܏a<|�a<�a<��a<>�a<a<G�a<��a<,�a<��a<B�a<ƕa<W�a<Ζa<k�a<��a<��a<�a<��a<�a<O�a<��a<�a<4�a<V�a<y�a<��a<�a<'�a<9�a<z�a<��a<�a<D�a<��a<�a<h�a<��a<�a<}�a<۟a< �a<|�a<��a<�a<	�a<�a<;�a<@�a<Q�a<T�a<u�a<��a<��a<��a<ġa<�a<�a<2�a<F�a<Y�a<V�a<N�a<7�a<�a<��a<��a<��a<k�a<M�a<�a<�a<Πa<��a<��a<��a<Ġa<�a<�a<��a<��a<-�a<6�a<<�a<B�a<4�a<�a<�a<ɠa<��a<^�a<�a<��a<͟a<��a<u�a<A�a<'�a<�a<�a<��a<��a<`�a<�a<ԝa<m�a<�a<��a<)�a<ɛa<l�a<�a<��a<�a<ԙa<�a<2�a<�a<ɘa<��a<S�a<�a<ߗa<��a<n�a<1�a<Ԗa<t�a<�a<��a<�a<��a<��a<d�a<�a<i�a<�a<o�a<��a<y�a<�a<��a<�a<��a<�a<v�a<�a<1�a<��a<ӊa<�a<~�a<ۈa<B�a<��a<�a<��a<�a<��a<;�a<�a<��a<`�a<�a<�a<��a<i�a<;�a<�a<��a<F�a<��a<��a<'�a<πa<o�a<1�a<�a<�a<ta<7a< a<a<�~a<�~a<�~a<q~a<A~a<~a<�}a<�}a<<}a<	}a<�|a<�|a<�|a<]|a<T|a<V|a<d|a<{|a<�|a<�|a<*}a<f}a<�  �  �}a<�}a<a~a<�~a<�~a<'a<Pa<�a<�a<�a<C�a<��a<��a<�a<T�a<}�a<��a<b�a<��a<4�a<y�a<�a<E�a<��a<�a<~�a<��a<��a<n�a<��a<�a<"�a<��a<�a<_�a<��a<�a<�a<Ċa<~�a<1�a<�a<��a<W�a<<�a<׏a<s�a<�a<��a<1�a<��a<K�a<ϓa<o�a<ǔa<Y�a<��a<Y�a<�a<}�a<��a<��a<��a<r�a<�a<F�a<��a<�a<�a<n�a<��a<��a<�a<�a<2�a<o�a<��a<�a<E�a<��a<�a<f�a<��a<E�a<�a<ԟa<?�a<o�a<��a<͠a<��a<�a<I�a<D�a<i�a<��a<h�a<��a<��a<ša<��a<�a<#�a<,�a<A�a<>�a<P�a<F�a<B�a<)�a<ۡa<�a<��a<W�a<.�a<��a<�a<��a<��a<��a<��a<��a<��a<֠a<�a<3�a<�a<@�a<N�a<6�a<(�a<��a<�a< a<��a<r�a<K�a<�a<ʟa<��a<h�a<e�a<C�a<�a<��a<��a<��a<D�a<�a<ɝa<��a<�a<��a<f�a<ɛa<d�a<ܚa<r�a<'�a<��a<_�a<%�a<�a<��a<��a<J�a<F�a<��a<��a<��a<,�a<˖a<g�a<��a<��a<�a<��a<�a<��a<��a<��a<��a<q�a<!�a<��a<�a<��a<�a<��a<��a<m�a<܌a<K�a<{�a<�a<W�a<z�a<Ոa<$�a<��a<��a<]�a<�a<��a<#�a<܄a<��a<\�a<L�a<�a<��a<��a<.�a<�a<��a<7�a<Ӂa<��a<*�a<�a<��a<%�a<�a<�a<�a<qa<8a<a<�~a<�~a<�~a<k~a<9~a<~a<�}a<w}a<j}a<&}a<�|a<�|a<m|a<b|a<>|a<B|a<F|a<�|a<�|a<�|a<}a<x}a<�  �  �}a<~a<W~a<�~a<�~a<3a<pa<�a<�a<�a<.�a<[�a<��a<�a<7�a<��a<فa<E�a<��a<$�a<��a<��a<a�a<��a<�a<^�a<��a<��a<1�a<��a<�a<M�a<��a<��a<��a< �a<��a<�a<�a<��a<:�a<�a<��a<u�a<�a<܏a<|�a<�a<��a<>�a<a<G�a<��a<,�a<��a<B�a<ƕa<W�a<Ζa<k�a<��a<��a<�a<��a<�a<O�a<��a<�a<4�a<V�a<y�a<��a<�a<'�a<9�a<z�a<��a<�a<D�a<��a<�a<h�a<��a<�a<}�a<۟a< �a<|�a<��a<�a<	�a<�a<;�a<@�a<Q�a<T�a<u�a<��a<��a<��a<ġa<�a<�a<2�a<F�a<Y�a<V�a<N�a<7�a<�a<��a<��a<��a<k�a<M�a<�a<�a<Πa<��a<��a<��a<Ġa<�a<�a<��a<��a<-�a<6�a<<�a<B�a<4�a<�a<�a<ɠa<��a<^�a<�a<��a<͟a<��a<u�a<A�a<'�a<�a<�a<��a<��a<`�a<�a<ԝa<m�a<�a<��a<)�a<ɛa<l�a<�a<��a<�a<ԙa<�a<2�a<�a<ɘa<��a<S�a<�a<ߗa<��a<n�a<1�a<Ԗa<t�a<�a<��a<�a<��a<��a<d�a<�a<i�a<�a<o�a<��a<y�a<�a<��a<�a<��a<�a<v�a<�a<1�a<��a<ӊa<�a<~�a<ۈa<B�a<��a<�a<��a<�a<��a<;�a<�a<��a<`�a<�a<�a<��a<i�a<;�a<�a<��a<F�a<��a<��a<'�a<πa<o�a<1�a<�a<�a<ta<7a< a<a<�~a<�~a<�~a<q~a<A~a<~a<�}a<�}a<<}a<	}a<�|a<�|a<�|a<]|a<T|a<V|a<d|a<{|a<�|a<�|a<*}a<f}a<�  �  �}a<7~a<T~a<�~a<�~a<a<ha<a<�a<�a<-�a<_�a<��a<�a<�a<��a<ցa<H�a<��a<�a<}�a<݃a<[�a<��a<�a<\�a<��a<(�a<O�a<Æa<Ԇa<9�a<��a<��a<��a<��a<��a<'�a<�a<k�a<P�a<�a<Ǎa<��a<�a<�a<r�a<�a<��a<)�a<��a<8�a<ɓa<+�a<̔a<3�a<��a<g�a<̖a<r�a<�a<r�a<�a<u�a<�a<A�a<��a<ޚa<G�a<z�a<��a<ڛa<Λa<$�a<D�a<}�a<��a<�a<I�a<��a<�a<I�a<�a<)�a<��a<�a<�a<|�a<��a<٠a<�a<�a<"�a<?�a<R�a<Q�a<��a<i�a<��a<��a<ˡa<��a<�a< �a<(�a<O�a<C�a<G�a<?�a<�a<�a<ԡa<��a<n�a<,�a<�a<�a<ܠa<��a<Ġa<��a<Ƞa<ʠa<�a<$�a< �a<V�a<2�a<>�a<=�a<�a<�a<Ԡa<��a<��a<\�a<$�a<��a<ǟa<y�a<��a<>�a<*�a< �a<Ҟa<��a<y�a<Z�a<�a<ԝa<k�a<�a<֜a<G�a< �a<Q�a<�a<��a<!�a<ۙa<v�a<8�a<�a<͘a<m�a<i�a<6�a<�a<֗a<c�a<;�a<ʖa<i�a<�a<|�a<��a<�a<�a<c�a<��a<Z�a<ґa<�a<ސa<��a<��a<}�a< �a<��a<�a<h�a<�a<(�a<��a<��a<:�a<��a<��a<@�a<��a<�a<��a<�a<��a<L�a<��a<��a<��a<0�a<�a<��a<f�a<;�a<ӂa<��a<,�a<Ձa<v�a<%�a<рa<k�a<G�a<�a<�a<{a<>a<%a<�~a<�~a<�~a<�~a<^~a<;~a<~a<�}a<�}a<]}a<5}a<�|a<�|a<�|a<a|a<b|a<N|a<s|a<}|a<�|a<�|a<#}a<�}a<�  �  �}a<~a<_~a<�~a<�~a<.a<[a<�a<�a<�a<�a<@�a<f�a<��a<�a<T�a<��a<�a<��a<�a<v�a<�a<U�a<��a<�a<~�a<��a<�a<a�a<��a<�a<X�a<ʇa<0�a<��a<�a<��a<[�a<�a<��a<N�a<�a<̍a<d�a<;�a<яa<t�a<�a<��a<,�a<��a<%�a<��a< �a<�a< �a<��a<�a<a<;�a<ޗa<o�a<��a<k�a<�a<M�a<��a<	�a<�a<y�a<��a<ӛa<	�a<A�a<u�a<��a<ٜa<�a<|�a<ԝa<�a<��a<ߞa<8�a<��a<͟a<E�a<c�a<��a<ܠa<�a<�a<�a<#�a<!�a<6�a<=�a<k�a<v�a<x�a<��a<ɡa< �a<�a<6�a<E�a<U�a<;�a<>�a<&�a<�a<�a<��a<�a<W�a<B�a<�a<��a<ݠa<�a<�a<�a<�a<��a<�a<4�a<-�a<=�a<I�a<+�a</�a<�a<�a<��a<��a<5�a<�a<��a<��a<��a<>�a<�a<��a<�a<͞a<��a<�a<T�a<�a<��a<��a<�a<��a<Y�a<�a<��a<�a<��a<U�a<�a<��a<d�a<$�a<�a<��a<g�a<7�a<�a<��a<��a<&�a<͖a<w�a<��a<�a<��a<l�a<ϓa<W�a<��a<G�a<Ǒa<-�a<Ԑa<I�a<�a<z�a<�a<~�a<�a<t�a<ьa<S�a<�a<��a<E�a<��a<��a<\�a<Ňa<4�a<��a<(�a<ͅa<r�a<�a<̄a<��a<?�a<��a<��a<��a<"�a<�a<��a<,�a<сa<q�a<
�a<��a<Q�a<�a<�a<�a<6a<'a<�~a<�~a<�~a<�~a<�~a<p~a</~a<~a<�}a<�}a<n}a<+}a<�|a<�|a<�|a<�|a<�|a<u|a<�|a<�|a<�|a<}a<>}a<�}a<�  �  �}a<~a<|~a<�~a<�~a<&a<,a<{a<�a<�a<�a<4�a<h�a<��a<��a<3�a<��a<
�a<s�a<�a<K�a<ԃa<$�a<��a<��a<��a<Ʌa<%�a<��a<��a<:�a<r�a<чa<A�a<��a<H�a<Ӊa<e�a< �a<ԋa<x�a<�a<�a<z�a<W�a<��a<z�a<��a<x�a<�a<}�a<�a<k�a<�a<q�a<��a<��a<�a<��a<�a<ϗa<A�a<Ԙa<O�a<ʙa<Q�a<��a< �a<5�a<��a<��a<�a<=�a<D�a<��a<��a<�a<D�a<��a<ڝa<4�a<��a<�a<V�a<��a<�a<M�a<U�a<��a<��a<ߠa<�a<��a<	�a<�a<>�a<�a<H�a<S�a<v�a<��a<��a<�a<�a<!�a<�a<F�a<?�a<4�a<C�a<�a<�a<��a<��a<��a<C�a<*�a<�a<�a<��a<��a<��a<�a<9�a<!�a<P�a<>�a<Z�a<C�a<*�a<'�a<٠a<Рa<~�a<i�a<�a<��a<��a<y�a<\�a<�a<$�a<�a<ʞa<��a<~�a<o�a<"�a<�a<��a<��a<*�a<Ӝa<y�a<��a<��a<,�a<Úa<f�a<�a<Ǚa<y�a<.�a<�a<֘a<��a<H�a<)�a<��a<��a<�a<Җa<V�a<ϕa<d�a<˔a<^�a<��a<S�a<��a<&�a<��a<�a<Ӑa<)�a<ڏa<L�a<�a<a�a<�a<x�a<Ìa<j�a<��a<�a<X�a<��a<*�a<_�a<χa<F�a<ʆa<N�a<ޅa<y�a<%�a<��a<��a<\�a<�a<��a<��a<�a<�a<f�a<�a<��a<I�a<��a<��a<Y�a<�a<�a<aa<4a<a<�~a<�~a<�~a<�~a<^~a<a~a<3~a<~a<�}a<�}a<�}a<7}a<'}a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<%}a<x}a<�}a<�  �  �}a<6~a<r~a<�~a<�~a<a<<a<ia<za<�a<�a<�a<8�a<z�a<��a<%�a<n�a<Ձa<H�a<ʂa<A�a<Ƀa<.�a<��a<�a<s�a<؅a<2�a<��a<��a<#�a<��a<�a<v�a<�a<Y�a<�a<��a<K�a<Ƌa<��a<@�a<�a<��a<3�a<ԏa<j�a<��a<��a<��a<j�a<�a<T�a<Ɠa<e�a<Δa<R�a<��a<g�a<��a<��a<-�a<Ęa<S�a<Ùa<:�a<��a<��a<V�a<��a<؛a<*�a<&�a<��a<��a<�a<�a<n�a<��a<�a<g�a<��a<*�a<c�a<��a<�a<6�a<o�a<��a<��a<ڠa<ڠa<�a<ݠa<�a<�a<�a<�a<,�a<U�a<c�a<��a<��a<ۡa<�a<&�a</�a<>�a<:�a<,�a< �a<��a<�a<��a<��a<��a<\�a<H�a<�a<,�a<%�a<?�a<�a<6�a<[�a<K�a<U�a<P�a<D�a<3�a<�a<�a<��a<r�a<B�a<��a<��a<��a<[�a<�a<�a<֞a<��a<��a<��a<t�a<d�a<-�a<��a<ȝa<��a<9�a<�a<|�a<9�a<��a<R�a<�a<��a<B�a<ؙa<��a<m�a<2�a<Șa<��a<k�a<'�a<ߗa<��a<)�a<a<L�a<ܕa<O�a<��a<1�a<��a<��a<��a<��a<q�a<�a<y�a<�a<��a<8�a<юa<f�a<ߍa<a�a<ڌa<B�a<��a<�a<v�a<�a<�a<��a<�a<s�a<��a<w�a<�a<��a<X�a<�a<τa<j�a<%�a<ڃa<�a<.�a<˂a<i�a<�a<��a<5�a<Āa<^�a<�a<�a<fa<9a<a<�~a<�~a<�~a<�~a<�~a<n~a<J~a<2~a<~a<�}a<�}a<�}a<h}a<3}a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<+}a<3}a<v}a<�}a<�  �  �}a<^~a<y~a<�~a<�~a<a<9a<,a<va<ya<�a<�a<�a<_�a<��a<�a<*�a<ˁa<!�a<��a<(�a<��a<9�a<��a<�a<r�a<�a<P�a<��a<�a<I�a<Շa<�a<��a<"�a<��a<9�a<��a<u�a<�a<a<N�a<�a<��a</�a<�a<V�a<��a<i�a<ˑa<s�a<��a<N�a<��a<*�a<��a<+�a<a<.�a<��a<^�a<2�a<��a<.�a<Йa<"�a<��a<��a<v�a<��a<�a<J�a<J�a<��a<��a<�a<O�a<��a<�a<�a<��a<Þa<M�a<g�a<˟a<�a<2�a<{�a<{�a<��a<��a<��a<Ѡa<��a<ڠa<��a<�a<ܠa<�a<�a<<�a<}�a<��a<ۡa<ѡa<�a<+�a<5�a<K�a<0�a<G�a<�a<�a<�a<��a<��a<`�a<��a<L�a<h�a<2�a<[�a<Z�a<W�a<t�a<Q�a<|�a<X�a<O�a</�a<�a<�a<��a<n�a<�a<�a<��a<H�a<@�a<�a<�a<��a<��a<x�a<u�a<[�a<)�a<7�a<�a<ѝa<��a<G�a<��a<��a<W�a<Ǜa<��a<�a<��a<v�a<�a<ߙa<d�a<\�a<�a<ۘa<y�a</�a<�a<�a<?�a<��a<T�a<��a<�a<��a<�a<��a<ʒa<Y�a<ґa<J�a<ڐa<@�a<	�a<i�a<=�a<��a<A�a<�a<I�a<�a<>�a<׋a< �a<��a<�a<7�a<ӈa<�a<��a<�a<��a<7�a<��a<��a<�a<�a<n�a<8�a<�a<|�a<;�a<��a<v�a<�a<|�a<%�a<��a<X�a<�a<�a<>a< a<�~a<�~a<�~a<p~a<�~a<K~a<e~a<F~a<(~a<~a<�}a<�}a<�}a<�}a<S}a<'}a< }a<�|a<}a<�|a<}a<�|a<H}a<m}a<�}a<�}a<�  �  5~a<]~a<�~a<�~a<�~a<�~a<a<&a<]a<Xa<ua<�a<�a<$�a<P�a<Ȁa<*�a<��a<�a<��a<�a<��a<�a<��a<�a<~�a<�a<^�a<Æa<�a<��a<�a<H�a<Ոa<?�a<��a<g�a<ڊa<x�a<�a<͌a<v�a<%�a<��a<E�a<ۏa<[�a<�a<Z�a<Ǒa<P�a<��a<�a<��a<��a<v�a<��a<��a<5�a<ʖa<8�a<�a<��a<(�a<��a<&�a<��a<�a<i�a<̛a<�a<K�a<��a<��a<�a<U�a<x�a<ĝa<$�a<P�a<��a<�a<F�a<��a<�a<�a<C�a<e�a<}�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ڠa<��a<1�a<@�a<`�a<��a<̡a<��a<�a<4�a<D�a<C�a<@�a<@�a<�a<�a<ءa<��a<��a<��a<t�a<��a<x�a<p�a<v�a<��a<|�a<��a<|�a<g�a<P�a<'�a<��a<��a<{�a<U�a<�a<��a<��a<6�a<�a<��a<��a<��a<��a<J�a<W�a<D�a< �a<�a<�a<��a<��a<H�a<�a<��a<U�a<�a<��a<:�a<��a<��a<6�a<�a<��a<`�a<!�a<�a<��a<`�a<��a<��a<1�a<��a<<�a<��a<�a<��a<ɓa<Y�a<̒a</�a<��a<�a<��a<G�a<؏a<D�a<�a<��a<;�a<̍a<M�a<܌a<V�a<ˋa<I�a<��a<�a<r�a<Ոa<A�a<݇a<>�a<͆a<u�a<�a<��a<J�a<�a<��a<P�a<�a<��a<$�a<��a<Q�a<؁a<j�a<�a<k�a<0�a<�a<oa<	a<�~a<�~a<�~a<n~a<L~a<o~a<F~a<C~a<:~a<'~a<~a<�}a<�}a<�}a<�}a<u}a<H}a<+}a<}a<)}a<}a<3}a<C}a<]}a<�}a<�}a<�}a<�  �  D~a<L~a<�~a<�~a<�~a<�~a<�~a<,a< a<aa<ca<|a<�a<�a<E�a<��a<�a<\�a<�a<z�a<�a<��a<��a<��a<��a<��a<��a<N�a<نa<(�a<��a<��a<��a<�a<j�a<��a<k�a<2�a<��a<O�a<��a<��a<'�a<��a<c�a<a<x�a<ǐa<R�a<��a<�a<��a<�a<Q�a<Γa<P�a<ڔa<c�a<��a<��a<S�a<җa<t�a<#�a<��a<M�a<��a<&�a<m�a<̛a<�a<]�a<��a<ڜa<L�a<\�a<��a<�a<3�a<��a<��a<.�a<X�a<��a<ԟa<�a<O�a<V�a<��a<z�a<��a<~�a<��a<��a<g�a<q�a<��a<��a<��a<Ša<�a< �a<t�a<��a<̡a<�a<�a<<�a</�a<^�a<2�a<K�a<"�a<!�a<�a<��a<�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<k�a<��a<D�a<)�a<��a<��a<��a<�a<��a<��a<A�a<�a<՞a<��a<��a<[�a<>�a<I�a<A�a<�a<)�a<��a<��a<��a<��a<\�a<��a<Мa<e�a<0�a<��a<��a<�a<��a<w�a<�a<��a<��a<Q�a<��a<��a<b�a<��a<��a<�a<Жa< �a<��a<�a<]�a<�a<!�a<��a<��a<w�a<��a<{�a<�a<��a<^�a<ގa<��a<6�a<��a<t�a<Ča<p�a<ϋa<I�a<��a< �a<��a<��a<��a<�a<z�a<��a<��a<?�a<��a<v�a<��a<��a<A�a<��a<��a<�a<؂a<3�a<ށa<D�a<�a<v�a<�a<�a<?a<�~a<�~a<�~a<_~a<M~a<a~a<0~a<F~a<3~a</~a<0~a< ~a<~a<�}a<�}a<�}a<�}a<q}a<e}a<g}a<:}a<S}a<L}a<{}a<�}a<�}a<�}a<�}a<�  �  T~a<}~a<�~a<�~a<�~a<�~a<�~a<a<a<&a<Da<ya<�a<�a<�a<��a<�a<]�a<ǁa<H�a<؂a<n�a<��a<��a<�a<�a<�a<{�a<�a<T�a<ća<�a<��a<�a<��a<�a<��a<-�a<��a<h�a<
�a<��a<:�a<܎a<b�a<Ϗa<k�a<��a<2�a<��a<�a<m�a<Вa<K�a<��a<*�a<��a<Q�a<�a<��a< �a<��a<_�a<�a<y�a<9�a<��a<#�a<��a<�a<>�a<��a<˜a<��a<M�a<t�a<ҝa<�a<>�a<��a<�a<<�a<��a<ɟa<��a<9�a<J�a<f�a<��a<e�a<��a<o�a<_�a<]�a<j�a<g�a<m�a<j�a<��a<��a<�a<�a<;�a<t�a<��a<סa<��a<<�a<;�a<c�a<d�a<[�a<R�a<?�a<�a<�a<�a<֡a<ޡa<��a<��a<��a<��a<ša<��a<��a<��a<��a<G�a<,�a<�a<��a<d�a<�a<��a<t�a<=�a<��a<��a<}�a<k�a<R�a<>�a<�a<�a<�a<	�a<ߝa<�a<��a<��a<o�a<*�a<�a<��a<A�a<֛a<��a<�a<��a<��a<2�a<��a<��a<j�a<#�a<јa<u�a<#�a<��a<$�a<Öa<�a<��a<�a<Q�a<��a<�a<��a<�a<Q�a<ѐa<i�a<��a<��a<+�a<Ǝa<l�a<�a<��a<`�a<Ќa<m�a<��a<a�a<܊a<M�a<��a<�a<��a<��a<��a<�a<��a<F�a<҅a<��a<*�a<Єa<j�a<�a<��a<%�a<��a<�a<��a<6�a<��a<D�a<�a<�a<*a<�~a<�~a<s~a<Z~a<2~a<'~a<$~a<'~a<~a<~a<0~a<~a<~a<�}a<�}a<�}a<�}a<�}a<u}a<^}a<\}a<v}a<p}a<w}a<�}a<�}a<~a<-~a<�  �  H~a<�~a<�~a<�~a<�~a<�~a<a<�~a<$a<a<a<Ka<ma<�a<�a<\�a<��a<8�a<��a<;�a<߂a<_�a<�a<j�a<�a<��a<��a<��a<�a<[�a<҇a<O�a<��a<:�a<��a<�a<ۊa<B�a<�a<��a<�a<��a<=�a<Վa<N�a<�a<C�a<ːa<B�a<��a<�a<0�a<��a<"�a<��a<�a<��a<"�a<��a<f�a<�a<ėa<Q�a<�a<��a<�a<��a<�a<��a<�a<=�a<��a<��a</�a<Y�a<ĝa<۝a<+�a<��a<��a<�a<N�a<��a<ğa<�a<)�a<K�a<u�a<^�a<��a<v�a<q�a<\�a<+�a<J�a<2�a<D�a<D�a<r�a<�a<��a<�a<�a<��a<��a<��a<�a<!�a<P�a<Q�a<n�a<S�a<Z�a<E�a<:�a<,�a<�a<�a<סa<�a<�a<ۡa<סa<ˡa<ơa<��a<��a<w�a<[�a<�a<۠a<��a<P�a<�a<��a<O�a<�a<a<��a<W�a<F�a<�a<�a<�a<�a<�a<��a<
�a<ȝa<ǝa<��a<]�a<4�a<ٜa<��a<P�a<	�a<��a<_�a<��a<��a<��a<�a<ԙa<��a<)�a<Ԙa<x�a<�a<��a<?�a<��a<$�a<��a<ߔa<]�a<w�a<��a<Z�a<��a<9�a<��a<;�a<Ώa<t�a<�a<ώa<_�a<�a<��a<6�a<�a<^�a<�a<i�a<ۊa<Q�a<͉a<J�a<��a<L�a<��a<4�a<چa<U�a<�a<��a<-�a<˄a<v�a<�a<��a<4�a<��a<H�a<��a<7�a<��a<�a<�a<Ma< a<�~a<�~a<=~a</~a<~a<�}a<6~a<~a<=~a<~a<~a<!~a<~a<	~a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<o}a<�}a<�}a<�}a<�}a<
~a<6~a<�  �  e~a<�~a<�~a<�~a<�~a<�~a<�~a<�~a<�~a<a<:a<Ga<la<�a<�a<N�a<��a<5�a<��a<2�a<��a<?�a<�a<r�a<�a<��a<�a<��a<��a<o�a<�a<I�a<��a<1�a<��a<6�a<Ċa<E�a<�a<��a<(�a<��a<V�a<�a<e�a<�a<G�a<��a<�a<j�a<��a<P�a<Ēa<�a<��a<�a<��a<�a<��a<n�a<�a<��a<0�a<�a<��a<�a<��a<$�a<��a< �a<L�a<��a<�a<*�a<[�a<��a<�a<8�a<{�a<��a<�a<^�a<��a<ݟa<�a<5�a<S�a<k�a<i�a<r�a<U�a<K�a<L�a<L�a<F�a<)�a<:�a<O�a<j�a<~�a<��a<��a<(�a<P�a<|�a<ʡa<��a<"�a<R�a<g�a<s�a<p�a<b�a<]�a<>�a<)�a<�a<�a<��a<�a<�a<ءa<ڡa<ޡa<Сa<��a<��a<��a<_�a<�a<ܠa<��a</�a<�a<��a<i�a<�a<��a<��a<b�a<8�a<�a<�a<�a<��a<�a<ڝa<�a<ϝa<��a<��a<n�a<>�a<��a<��a<`�a<�a<��a<V�a<
�a<��a<k�a<�a<әa<��a<A�a<�a<��a<(�a<��a<?�a<��a<�a<s�a<��a<.�a<��a<�a<H�a<��a<;�a<��a<7�a<��a<{�a<�a<��a<>�a<��a<��a<>�a<�a<m�a<��a<}�a<�a<g�a<ԉa<E�a<��a<:�a<��a<A�a<̆a<S�a<�a<��a<A�a<�a<��a<�a<��a<*�a<��a<+�a<��a<�a<��a<3�a<�a<Da<�~a<�~a<x~a<<~a<%~a<'~a<~a< ~a<�}a<~a<~a<~a<#~a<~a<~a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<~a<@~a<�  �  �a<�a<�a<!�a<E�a<k�a<u�a<��a<��a<��a<ˀa<�a<:�a<^�a<Ɂa<�a<y�a<��a<S�a<уa<V�a<	�a<]�a<��a<Z�a<�a<`�a<чa<P�a<ƈa<5�a<��a<3�a<��a<�a<��a<�a<��a<H�a<��a<c�a<��a<��a<��a<��a<��a<��a<�a<z�a<��a<0�a<��a<��a<~�a<��a<p�a<��a<�a<�a<��a<K�a<՘a<��a<&�a<��a<:�a<��a<-�a<{�a<�a<P�a<��a<ٝa<=�a<}�a<��a<�a<P�a<}�a<�a<�a<^�a<��a<Ԡa<�a<,�a<Y�a<^�a<��a<��a<��a<��a<��a<��a<p�a<��a<��a<��a<��a<�a<�a<&�a<s�a<��a<��a<��a<)�a<@�a<C�a<o�a<^�a<}�a<n�a<h�a<=�a<T�a</�a<�a<=�a<�a<��a<�a<ޢa<�a<٢a<Ϣa<��a<��a<X�a<3�a<�a<¡a<��a<2�a<��a<��a<N�a<3�a<�a<՟a<��a<��a<J�a<R�a<A�a<3�a<O�a<�a<�a<��a<��a<q�a<1�a<��a<��a<h�a<
�a<ݜa<e�a<"�a<�a<v�a<2�a<��a<��a<G�a<�a<��a<�a<Øa<+�a<җa<>�a<��a<<�a<p�a<�a<8�a<��a<(�a<��a<"�a<��a<>�a<��a<w�a<�a<͏a<f�a<�a<��a<�a<��a<�a<��a<3�a<��a<�a<��a<�a<��a<2�a<��a<$�a<�a<[�a< �a<��a<6�a<˅a<b�a< �a<{�a<,�a<��a<X�a<��a<=�a<ցa<P�a<�a<��a<y�a<+�a<	�a<�a<�a<�a<�a<�a<�a<�a<�a<{a<�a<`a<ma<Qa<Ba<a<,a<a<a<<a<a<,a<^a<Wa<�a<�a<�  �  �a< �a<�a<3�a<C�a<a�a<k�a<v�a<��a<��a<�a<�a<<�a<j�a<��a<�a<y�a<ނa<X�a<ԃa<F�a<Ʉa<X�a<�a<a�a<�a<l�a<�a<O�a<��a<)�a<��a<�a<��a<�a<��a<#�a<��a<B�a<ȍa<d�a<�a<��a<�a<��a<�a<��a<��a<V�a<Ēa<7�a<��a<�a<��a<�a<q�a<��a<��a<�a<��a<C�a<��a<l�a<��a<��a<�a<��a<*�a<��a<��a<I�a<��a<�a<5�a<g�a<a<��a<C�a<��a<ɟa<�a<R�a<��a<ՠa<�a<@�a<d�a<h�a<~�a<��a<~�a<}�a<��a<��a<��a<��a<��a<��a<��a<�a<�a<?�a<i�a<��a<��a<�a<�a<:�a<X�a<m�a<y�a<}�a<d�a<b�a<P�a<I�a<2�a<.�a<�a<�a<�a<��a<�a<�a<Ңa<Тa<��a<��a<k�a<1�a<�a<��a<l�a<0�a<��a<��a<k�a<4�a<�a<˟a<��a<��a<g�a<W�a<E�a<#�a<�a<�a<�a<Ǟa<��a<}�a<F�a<��a<��a<\�a<�a<��a<o�a< �a<a<��a<'�a<�a<��a<G�a<�a<��a</�a<��a<=�a<��a<3�a<��a<�a<w�a<�a<M�a<a<6�a<��a<!�a<��a<D�a<Րa<o�a<�a<��a<<�a<�a<|�a<�a<��a<6�a<��a<-�a<��a<�a<��a<�a<��a<�a<��a<4�a<��a<[�a<�a<��a<7�a<߅a<v�a<�a<��a<�a<��a<�a<��a<B�a<Ձa<k�a<�a<��a<r�a<0�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<|a<ma<Ga<<a<'a<"a<a<a<a<'a<3a<Ma<ga<�a<�a<�  �  �a<�a<�a<1�a<H�a<h�a<��a<��a<��a<��a<��a<�a<<�a<��a<a<�a<v�a<�a<S�a<�a<m�a<ׄa<~�a<�a<h�a<�a<H�a<Ňa<>�a<��a<�a<��a<�a<��a<�a<f�a<,�a<��a<+�a<��a<V�a<�a<o�a<��a<w�a<�a<��a<�a<�a<ْa<_�a<��a<!�a<��a<�a<|�a<��a<��a<�a<��a<B�a<�a<��a<!�a<��a<+�a<��a<�a<u�a<ٜa<:�a<��a<ӝa<%�a<`�a<˞a<�a<?�a<��a<��a<�a<D�a<��a<àa<�a<�a<H�a<q�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<աa<�a<�a<D�a<e�a<��a<¢a<�a<)�a<<�a<Y�a<H�a<_�a<_�a<e�a<U�a<K�a<3�a<&�a<7�a<�a<�a<��a<�a<�a<բa<Ңa<��a<��a<m�a<h�a<6�a<�a<ۡa<u�a<Z�a<��a<��a<u�a<4�a<�a<Οa<��a<��a<x�a<R�a<T�a<K�a<�a<(�a<�a<Ξa<��a<Y�a<%�a<�a<��a<P�a<�a<��a<s�a<�a<��a<��a< �a<ؚa<��a<:�a<�a<|�a<�a<��a<H�a<��a<Q�a<��a<�a<��a<ޔa<\�a<��a<8�a<��a<)�a<��a<@�a<�a<m�a<5�a<��a<a�a<	�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<��a<��a<��a<��a<=�a<��a<\�a<�a<��a<%�a<��a<O�a<�a<��a<�a<��a<-�a<̂a<\�a<сa<��a<�a<ʀa<y�a<G�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<ba<ba<Oa<Ha<.a<"a<a<a<$a<�~a<.a<*a<9a<da<ya<�a<�  �  �a<�a<�a<+�a<M�a<]�a<t�a<��a<��a<��a<��a<�a<O�a<��a<�a<+�a<��a<��a<{�a<�a<^�a<�a<]�a<�a<h�a<�a<m�a<Їa<E�a<��a<�a<{�a<�a<c�a<��a<x�a<�a<��a<�a<��a<C�a<�a<o�a<	�a<��a<�a<��a<�a<z�a<�a<I�a<˓a<6�a<��a<�a<��a<&�a<��a<0�a<̗a<j�a<�a<��a<#�a<��a<8�a<��a<,�a<��a<ݜa<A�a<�a<ǝa<�a<`�a<��a<�a<'�a<Z�a<a<��a<@�a<��a<ʠa<��a<>�a<X�a<k�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<֡a<�a<�a<%�a<_�a<��a<��a<֢a<��a<�a<G�a<Q�a<u�a<i�a<a�a<\�a<F�a<0�a<+�a<�a<��a<��a<�a<ܢa<�a<ʢa<ʢa<Ţa<��a<��a<��a<c�a<;�a<��a<��a<��a<B�a<�a<Рa<��a<G�a<�a<�a<��a<��a<��a<z�a<a�a<;�a<6�a<�a<��a<Ξa<��a<~�a</�a<�a<��a<J�a<�a<��a<C�a<�a<��a<L�a<�a<Ța<u�a<'�a<�a<{�a<%�a<Ƙa<9�a<Ηa</�a<��a<$�a<��a<	�a<p�a<Гa<J�a<Вa<S�a<͑a<Y�a<��a<��a<#�a<��a<c�a<�a<��a<�a<��a<.�a<��a<$�a<��a<��a<z�a<��a<\�a< �a<��a<�a<��a<=�a<�a<��a<,�a<ƅa<s�a<��a<��a<"�a<��a<B�a<a<]�a<��a<��a<*�a<Հa<��a<\�a<&�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<la<Qa<>a< a<a<a<�~a<�~a<�~a<�~a<a<9a<Ca<na<�a<�  �  �a<�a<	�a<�a<`�a<|�a<��a<��a<��a<��a<�a<5�a<q�a<��a< �a<;�a<��a<�a<��a<�a<c�a<�a<j�a<�a<o�a<چa<R�a<��a<0�a<��a<�a<_�a<�a<T�a<ъa<i�a<̋a<��a<��a<��a<-�a<ǎa<_�a<�a<��a<��a<��a<�a<��a<��a<R�a<�a<6�a<Ĕa<0�a<��a<0�a<��a<Y�a<Ηa<��a< �a<��a<=�a<��a<M�a<��a<�a<o�a<̜a<$�a<a�a<ʝa<�a<M�a<n�a<ўa<�a<I�a<��a<ҟa<C�a<^�a<��a<�a<�a<N�a<l�a<��a<��a<áa<��a<��a<áa<��a<ѡa<ǡa<�a<�a<#�a<E�a<^�a<��a<��a<��a<�a<1�a<\�a<@�a<a�a<K�a<W�a<6�a<@�a<#�a<�a<�a<آa<�a<âa<עa<ˢa<��a<ʢa<��a<��a<��a<��a<Q�a<N�a<�a<١a<��a<B�a<1�a<ՠa<��a<i�a<"�a<�a<˟a<��a<��a<��a<v�a<A�a<T�a<�a<�a<֞a<��a<c�a<�a<۝a<q�a<K�a<Мa<��a<3�a<�a<��a<2�a<�a<��a<v�a<�a<��a<k�a<
�a<��a<*�a<�a<D�a<іa<7�a<��a<�a<q�a<��a<d�a<ؒa<]�a<�a<��a<��a<��a<0�a<Ϗa<~�a<�a<��a<�a<��a<�a<��a<�a<l�a<�a<S�a<�a<G�a<�a<i�a<�a<��a<�a<�a<^�a<�a<��a<U�a<��a<��a<<�a<��a<`�a<ɂa<n�a<�a<��a<O�a<�a<��a<b�a<E�a<�a<�a<�a<�a<�a<�a<�a<�a<xa<{a<Na<Ga<a<a<�~a<�~a<�~a<�~a<�~a<�~a<a<a</a<na<va<�  �  �a<�a<�a<.�a<J�a<^�a<��a<��a<�a<��a<�a<_�a<��a<΁a<�a<i�a<Ȃa<=�a<��a<�a<��a<�a<��a<�a<n�a<�a<M�a<��a<,�a<��a<�a<^�a<��a<>�a<��a<*�a<ԋa<J�a<�a<��a< �a<Îa<`�a<��a<|�a<�a<��a<�a<��a<��a<��a<ܓa<c�a<ؔa<L�a<֕a<Z�a<ؖa<h�a<�a<x�a<.�a<��a<6�a<��a<'�a<��a<�a<t�a<Ϝa<�a<V�a<��a<�a<�a<s�a<��a<�a<=�a<o�a<ӟa<�a<X�a<��a<�a<�a<J�a<w�a<��a<��a<��a<͡a<ѡa<��a<�a<�a<�a<	�a<"�a<9�a<h�a<{�a<��a<�a<�a<�a<�a<<�a<Z�a<P�a<V�a<L�a<5�a<'�a<�a<�a<עa<٢a<��a<��a<��a<��a<��a<��a<��a<��a<��a<w�a<f�a<8�a<��a<�a<��a<��a<.�a<�a<Ơa<��a<R�a<#�a<��a<ןa<Ɵa<��a<��a<u�a<N�a<,�a<�a<՞a<��a<^�a<�a<֝a<s�a<�a<Μa<a�a<�a<Ǜa<h�a<:�a<֚a<��a<Z�a<�a<��a<l�a<�a<��a<N�a<��a<E�a<͖a<<�a<̕a<�a<��a<�a<�a<�a<��a<�a<��a<+�a<��a<^�a<ޏa<v�a<�a<��a<&�a<��a<�a<��a<�a<b�a<�a<N�a<��a<M�a<��a<C�a<�a<e�a<�a<��a<X�a<�a<��a<P�a<�a<��a<�a<a<Y�a<�a<��a<�a<Ɓa<c�a<�a<πa<��a<[�a<@�a<�a<�a<�a<�a<�a<�a<�a<�a<ka<Ya<<a<a<a<�~a<�~a<�~a<�~a<�~a<�~a<�~a<�~a<"a<Oa<va<�  �  {a<�a<�a<2�a<Y�a<t�a<��a<��a<��a<�a<X�a<{�a<��a<��a<(�a<��a<̂a<k�a<��a<!�a<��a<��a<��a<�a<��a<Նa<B�a<��a<��a<�a<��a<c�a<��a<�a<��a<�a<��a<�a<��a<b�a<�a<��a<6�a<��a<f�a<5�a<��a<'�a<��a<�a<��a<�a<��a<ޔa<i�a<��a<r�a<��a<o�a<H�a<��a<;�a<��a<>�a<՚a<)�a<ӛa<��a<v�a<��a<��a<H�a<v�a<��a<�a<I�a<��a<Ԟa<
�a<N�a<۟a<�a<Q�a<}�a<ڠa<�a<<�a<��a<��a<ȡa<��a<֡a<ߡa<�a<�a<�a<�a<�a<N�a<H�a<z�a<âa<��a<��a<�a<3�a<6�a<G�a<f�a<@�a<\�a<�a<(�a<��a<��a<�a<��a<��a<��a<��a<u�a<��a<��a<|�a<��a<p�a<��a<j�a<i�a<H�a<�a<�a<��a<��a<9�a<*�a<�a<��a<��a<5�a<(�a<۟a<��a<��a<��a<��a<E�a<M�a<��a<�a<��a<S�a<�a<��a<o�a<�a<Ԝa<K�a<�a<��a<K�a<�a<��a<��a<,�a<�a<��a<B�a<�a<��a<g�a<×a<d�a<ߖa<G�a<וa<+�a<�a<�a<��a<%�a<��a<)�a<��a<r�a<��a<k�a<�a<~�a<"�a<��a<C�a<~�a<�a<k�a<܋a<T�a<��a<]�a<��a<#�a<��a<2�a<��a<D�a<$�a<��a<Q�a<߅a<��a<K�a<�a<��a<�a<��a<S�a<��a<��a<2�a<��a<e�a<=�a<��a<��a<j�a<Q�a<T�a<�a<�a<�a<�a<�a<�a<�a<[a<_a<a<
a<�~a<�~a<�~a<�~a<�~a<�~a<�~a<�~a<�~a<a<!a<la<�  �  �a<�a<�a< �a<[�a<��a<��a<�a<�a<1�a<]�a<{�a<āa<�a<K�a<��a<��a<Z�a<ڃa<H�a<��a<+�a<��a<��a<z�a<ˆa<&�a<��a<�a<p�a<��a<�a<��a<��a<{�a<��a<��a<�a<��a<7�a<��a<��a<:�a<ڏa<f�a<�a<��a<'�a<��a<9�a<��a<$�a<��a<�a<��a<�a<��a<+�a<��a<:�a<ʘa<D�a<�a<^�a<Кa<<�a<��a<��a<X�a<��a<�a<<�a<V�a<��a<�a< �a<m�a<��a<�a<G�a<��a<ԟa<G�a<t�a<Ša<��a<3�a<��a<��a<ša<�a<�a<��a<�a<�a<�a<D�a<:�a<a�a<{�a<��a<��a<ܢa<��a<&�a<7�a<C�a<P�a<M�a<1�a<=�a<'�a<�a<�a<��a<Ƣa<��a<��a<~�a<v�a<m�a<{�a<^�a<q�a<��a<y�a<y�a<V�a<X�a<I�a< �a<��a<סa<��a<i�a</�a<�a<��a<��a<W�a<G�a<
�a<�a<ٟa<��a<��a<q�a<F�a<
�a<�a<��a<7�a<��a<��a<a�a<�a<��a<>�a<؛a<��a<;�a<�a<��a<f�a<�a<ݙa<��a<F�a<��a<��a<F�a<ԗa<d�a<�a<z�a<ޕa<a�a<ܔa<;�a<Γa<5�a<��a<U�a<đa<d�a<��a<u�a<�a<��a<�a<��a<%�a<�a<��a<g�a<΋a<G�a<��a<�a<��a<��a<��a<�a<��a<=�a<܆a<v�a<G�a<օa<��a<-�a<ڄa<��a</�a<݃a<|�a<�a<��a<[�a<�a<��a<c�a< �a<Ӏa<��a<b�a<Q�a<-�a<�a<�a<�a<�a<�a<�a<La<@a<a<�~a<�~a<�~a<�~a<�~a<z~a<|~a<�~a<�~a<�~a<�~a<a<\a<�  �  �a<�a<�a</�a<G�a<��a<��a<�a<��a<T�a<g�a<��a<�a<�a<��a<��a<4�a<��a<��a<]�a<��a<3�a<��a<�a<\�a<�a<6�a<��a<��a<-�a<��a<��a<t�a<�a<I�a<܊a<Y�a<�a<��a<@�a<܍a<w�a<C�a<��a<��a<�a<��a<+�a<��a<>�a<��a<M�a<��a<?�a<��a<2�a<��a<)�a<җa<:�a<�a<O�a<�a<Z�a<Κa<K�a<��a<�a<D�a<��a<՜a<�a<`�a<z�a<ӝa<��a<D�a<��a<؞a<0�a<i�a<؟a<�a<s�a<Ơa<��a<X�a<^�a<��a<��a<�a<�a<�a<.�a<)�a<P�a<<�a<x�a<w�a<��a<Ģa<âa<�a<��a<,�a<*�a<I�a<E�a<S�a<V�a<'�a<+�a<�a<�a<��a<��a<��a<_�a<j�a<F�a<U�a<M�a<Q�a<r�a<J�a<|�a<j�a<x�a<g�a<5�a<,�a<��a<�a<��a<��a<9�a<�a<�a<��a<��a<D�a<C�a<�a<�a<͟a<��a<y�a<;�a<�a<Þa<��a<G�a<��a<��a<�a<�a<j�a<�a<a<Y�a<�a<��a<��a<.�a<
�a<��a<p�a<O�a<ݘa<��a<4�a<ݗa<h�a<�a<�a<�a<��a<ڔa<v�a<֓a<b�a<�a<S�a<��a<d�a<�a<�a<�a<��a<�a<��a<�a<��a<�a<p�a<��a<�a<��a<�a<r�a<׈a<]�a<߇a<�a<&�a<��a<z�a<�a<Յa<��a<3�a<��a<{�a<C�a<ԃa<~�a<�a<Âa<v�a<	�a<́a<[�a<>�a<�a<��a<��a<U�a<X�a<�a<�a<�a<�a<�a<�a<qa<*a<a<�~a<�~a<�~a<k~a<i~a<L~a<i~a<\~a<�~a<�~a<�~a<a<a<�  �  da<�a<�a< �a<Y�a<��a<ƀa<��a<%�a<P�a<~�a<Ёa<��a<@�a<��a<Ղa<7�a<��a<��a<g�a<ۄa<>�a<��a<$�a<n�a<نa<�a<��a<ۇa<*�a<��a<��a<P�a<ŉa<C�a<ʊa<G�a<܋a<~�a<*�a<ˍa<n�a<&�a<��a<r�a<�a<��a<J�a<ƒa<R�a<ʓa<J�a<Ɣa<T�a<��a<L�a<Ԗa<<�a<�a<d�a<�a<n�a<��a<m�a<�a<Y�a<��a<�a<4�a<��a<ɜa<�a<G�a<w�a<��a<�a<7�a<{�a<��a<�a<k�a<ßa< �a<^�a<��a<�a<C�a<p�a<��a<ءa<�a<�a<�a<0�a<I�a<Z�a<Y�a<��a<��a<��a<ޢa<ܢa<�a<!�a<?�a<I�a<d�a<T�a<I�a<6�a<�a<�a<ޢa<Ѣa<��a<��a<e�a<N�a<M�a<7�a<3�a<;�a<K�a<W�a<I�a<Z�a<S�a<X�a<W�a<G�a<E�a<�a<�a<��a<��a<P�a<8�a<�a<Ša<��a<e�a<F�a<)�a<��a<ןa<��a<��a<X�a</�a<Ԟa<��a</�a<�a<��a<�a<Ԝa<l�a<��a<��a<T�a<�a<��a<g�a<*�a<��a<��a<h�a<3�a<Ϙa<��a<7�a<�a<��a<�a<��a<	�a<��a< �a<��a<�a<|�a<�a<g�a<�a<��a<�a<��a<5�a<��a<;�a<��a<�a<��a<֌a<U�a<��a<�a<�a<��a<I�a<Èa<Q�a<هa<d�a<��a<��a<f�a< �a<��a<z�a<�a<�a<��a<S�a<��a<��a<>�a<Ԃa<x�a<)�a<ׁa<x�a<M�a<	�a<ǀa<��a<n�a<U�a<6�a<�a<�a<�a<�a<�a<Qa<a<�~a<�~a<�~a<�~a<_~a<E~a<;~a<L~a<M~a<d~a<�~a<�~a<�~a<a<�  �  Na<�a<�a<�a<\�a<w�a<��a<�a<4�a<\�a<��a<ˁa<�a<l�a<{�a<�a<I�a<��a<�a<x�a<�a<>�a<��a<��a<x�a<͆a<4�a<��a<ɇa<C�a<t�a<�a<B�a<��a<*�a<��a<<�a<a<v�a<�a<эa<v�a<�a<ڏa<l�a<�a<��a<'�a<��a<K�a<ݓa<N�a<�a<N�a<��a<_�a<ؖa<��a<�a<z�a<�a<��a<��a<e�a<њa<7�a<��a<��a<^�a<��a<̜a<�a<!�a<m�a<��a<ڝa<�a<[�a<��a<�a<S�a<��a<�a<O�a<��a<�a<6�a<}�a<��a<ɡa<�a<�a<1�a<A�a<V�a<d�a<��a<p�a<��a<Тa<٢a<�a<�a<3�a<8�a<A�a<=�a<Q�a<H�a<7�a<6�a<��a<�a<��a<��a<x�a<O�a<C�a<*�a<,�a<�a<*�a<+�a<:�a<`�a<D�a<o�a<_�a<T�a<J�a<�a<
�a<�a<͡a<��a<r�a<3�a<�a<�a<��a<��a<X�a<0�a<�a<�a<��a<��a<O�a<�a<ޞa<��a<E�a<�a<s�a<3�a<��a<Q�a<�a<��a<;�a<�a<��a<N�a<#�a<Ιa<��a<p�a<!�a<��a<��a<@�a<ϗa<d�a<��a<��a<�a<��a<�a<��a<'�a<��a<�a<��a<�a<��a<�a<��a<.�a<��a<�a<��a<�a<��a<��a<M�a<��a< �a<Y�a<։a</�a<��a<)�a<��a<S�a<�a<��a<:�a<�a<��a<��a<;�a<ބa<��a<+�a<�a<��a<C�a<�a<��a<6�a<�a<��a<6�a<+�a<�a<��a<��a<]�a<H�a<�a<�a<�a<�a<a<Ra<9a<�~a<�~a<�~a<a~a<Q~a</~a<0~a<)~a<A~a<P~a<|~a<�~a<�~a<5a<�  �  Ca<�a<�a<�a<a�a<��a<݀a<�a<2�a<i�a<��a<߁a<�a<h�a<��a<�a<W�a<��a<�a<��a<�a<]�a<��a<�a<t�a<ˆa<#�a<h�a<��a<�a<w�a<ۈa<A�a<��a<�a<��a<,�a<ċa<^�a<�a<��a<P�a<��a<��a<b�a<�a<��a<N�a<�a<^�a<�a<_�a<�a<\�a<�a<d�a<�a<z�a<�a<��a<�a<��a<	�a<��a<��a<Z�a<��a<�a<9�a<l�a<��a<�a<#�a<W�a<��a<ҝa<�a<L�a<��a<��a<G�a<��a<�a<=�a<��a<�a<2�a<s�a<��a<�a<�a<�a<>�a<M�a<o�a<n�a<��a<��a<��a<Тa<�a<�a<�a<0�a<J�a<a�a<_�a<[�a<A�a<8�a<�a<�a<Ȣa<��a<��a<i�a<R�a<.�a<(�a<�a< �a<�a<-�a<6�a<7�a<9�a<M�a<Z�a<N�a<O�a<:�a<*�a<�a<ˡa<��a<t�a<F�a<�a<�a<��a<��a<f�a<I�a<�a<��a<��a<��a<h�a<'�a<ڞa<��a<5�a<ȝa<f�a<	�a<��a<L�a<�a<��a<&�a<ٚa<��a<P�a<�a<ҙa<��a<J�a<
�a<Иa<��a<5�a<�a<��a<!�a<��a<#�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<1�a<��a<@�a<ʏa<A�a<��a<�a<v�a<یa<,�a<��a<��a<Z�a<��a<3�a<��a< �a<��a<O�a<�a<��a<<�a<�a<��a<X�a<!�a<لa<��a<M�a<��a<��a<D�a<�a<��a<O�a<�a<��a<W�a<+�a<�a<��a<��a<j�a<F�a<)�a<�a<�a<�a<ya<Ra<a<�~a<�~a<�~a<f~a<B~a<2~a<~a<'~a<)~a<R~a<p~a<�~a<�~a<a<�  �  �a<�a<�a<�a<Q�a<��a<Àa<�a<;�a<o�a<��a<��a<�a<_�a<Ղa<��a<W�a<ʃa<�a<��a<�a<[�a<��a< �a<_�a<Նa<.�a<��a<��a<�a<��a<a<"�a<��a<�a<��a<"�a<ȋa<F�a<�a<��a<n�a<9�a<��a<z�a<��a<��a<8�a<͒a<]�a<�a<h�a<�a<|�a<וa<w�a<�a<f�a<�a<��a<�a<��a<�a<w�a<ۚa<Y�a<��a<�a<E�a<��a<ќa<�a<*�a<B�a<��a<ŝa<
�a<L�a<��a<�a<2�a<��a<�a<|�a<��a<��a<E�a<a�a<��a<ȡa<	�a<'�a<@�a<:�a<v�a<v�a<��a<Ţa<��a<Ƣa<�a<��a< �a<:�a<K�a<I�a<U�a<M�a<<�a<E�a<�a<'�a<Ӣa<��a<��a<L�a<Q�a<#�a<3�a<�a< �a<�a<�a<3�a<<�a<x�a<S�a<d�a<N�a<?�a<7�a<�a<�a<ԡa<��a<g�a<^�a<�a<�a<�a<��a<f�a<S�a<�a<��a<˟a<��a<L�a<+�a<ƞa<��a<?�a<�a<��a<�a<��a<3�a<̛a<��a<%�a<ߚa<��a<S�a<�a<ՙa<��a<g�a<E�a<٘a<��a<*�a<�a<u�a<�a<��a<'�a<��a<�a<��a<
�a<��a</�a<��a<1�a<��a<-�a<��a<C�a<��a<(�a<��a<�a<��a<�a<[�a<��a<�a<b�a<��a<1�a<��a<#�a<��a<B�a<ۆa<{�a<H�a<�a<ޅa<z�a<+�a<�a<~�a<O�a<��a<��a<M�a<�a<��a<V�a<�a<��a<��a<)�a<�a<ހa<��a<r�a<P�a<*�a<�a<�a<�a<ta<`a<a<a<�~a<�~a<]~a<%~a<1~a<~a<2~a<~a<Q~a<V~a<�~a<�~a<a<�  �  Ca<�a<�a<�a<a�a<��a<݀a<�a<2�a<i�a<��a<߁a<�a<h�a<��a<�a<W�a<��a<�a<��a<�a<]�a<��a<�a<t�a<ˆa<#�a<h�a<��a<�a<w�a<ۈa<A�a<��a<�a<��a<,�a<ċa<^�a<�a<��a<P�a<��a<��a<b�a<�a<��a<N�a<�a<^�a<�a<_�a<�a<\�a<�a<d�a<�a<z�a<�a<��a<�a<��a<	�a<��a<��a<Z�a<��a<�a<9�a<l�a<��a<�a<#�a<W�a<��a<ҝa<�a<L�a<��a<��a<G�a<��a<�a<=�a<��a<�a<2�a<s�a<��a<�a<�a<�a<>�a<M�a<o�a<n�a<��a<��a<��a<Тa<�a<�a<�a<0�a<J�a<a�a<_�a<[�a<A�a<8�a<�a<�a<Ȣa<��a<��a<i�a<R�a<.�a<(�a<�a< �a<�a<-�a<6�a<7�a<9�a<M�a<Z�a<N�a<O�a<:�a<*�a<�a<ˡa<��a<t�a<F�a<�a<�a<��a<��a<f�a<I�a<�a<��a<��a<��a<h�a<'�a<ڞa<��a<5�a<ȝa<f�a<	�a<��a<L�a<�a<��a<&�a<ٚa<��a<P�a<�a<ҙa<��a<J�a<
�a<Иa<��a<5�a<�a<��a<!�a<��a<#�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<1�a<��a<@�a<ʏa<A�a<��a<�a<v�a<یa<,�a<��a<��a<Z�a<��a<3�a<��a< �a<��a<O�a<�a<��a<<�a<�a<��a<X�a<!�a<لa<��a<M�a<��a<��a<D�a<�a<��a<O�a<�a<��a<W�a<+�a<�a<��a<��a<j�a<F�a<)�a<�a<�a<�a<ya<Ra<a<�~a<�~a<�~a<f~a<B~a<2~a<~a<'~a<)~a<R~a<p~a<�~a<�~a<a<�  �  Na<�a<�a<�a<\�a<w�a<��a<�a<4�a<\�a<��a<ˁa<�a<l�a<{�a<�a<I�a<��a<�a<x�a<�a<>�a<��a<��a<x�a<͆a<4�a<��a<ɇa<C�a<t�a<�a<B�a<��a<*�a<��a<<�a<a<v�a<�a<эa<v�a<�a<ڏa<l�a<�a<��a<'�a<��a<K�a<ݓa<N�a<�a<N�a<��a<_�a<ؖa<��a<�a<z�a<�a<��a<��a<e�a<њa<7�a<��a<��a<^�a<��a<̜a<�a<!�a<m�a<��a<ڝa<�a<[�a<��a<�a<S�a<��a<�a<O�a<��a<�a<6�a<}�a<��a<ɡa<�a<�a<1�a<A�a<V�a<d�a<��a<p�a<��a<Тa<٢a<�a<�a<3�a<8�a<A�a<=�a<Q�a<H�a<7�a<6�a<��a<�a<��a<��a<x�a<O�a<C�a<*�a<,�a<�a<*�a<+�a<:�a<`�a<D�a<o�a<_�a<T�a<J�a<�a<
�a<�a<͡a<��a<r�a<3�a<�a<�a<��a<��a<X�a<0�a<�a<�a<��a<��a<O�a<�a<ޞa<��a<E�a<�a<s�a<3�a<��a<Q�a<�a<��a<;�a<�a<��a<N�a<#�a<Ιa<��a<p�a<!�a<��a<��a<@�a<ϗa<d�a<��a<��a<�a<��a<�a<��a<'�a<��a<�a<��a<�a<��a<�a<��a<.�a<��a<�a<��a<�a<��a<��a<M�a<��a< �a<Y�a<։a</�a<��a<)�a<��a<S�a<�a<��a<:�a<�a<��a<��a<;�a<ބa<��a<+�a<�a<��a<C�a<�a<��a<6�a<�a<��a<6�a<+�a<�a<��a<��a<]�a<H�a<�a<�a<�a<�a<a<Ra<9a<�~a<�~a<�~a<a~a<Q~a</~a<0~a<)~a<A~a<P~a<|~a<�~a<�~a<5a<�  �  da<�a<�a< �a<Y�a<��a<ƀa<��a<%�a<P�a<~�a<Ёa<��a<@�a<��a<Ղa<7�a<��a<��a<g�a<ۄa<>�a<��a<$�a<n�a<نa<�a<��a<ۇa<*�a<��a<��a<P�a<ŉa<C�a<ʊa<G�a<܋a<~�a<*�a<ˍa<n�a<&�a<��a<r�a<�a<��a<J�a<ƒa<R�a<ʓa<J�a<Ɣa<T�a<��a<L�a<Ԗa<<�a<�a<d�a<�a<n�a<��a<m�a<�a<Y�a<��a<�a<4�a<��a<ɜa<�a<G�a<w�a<��a<�a<7�a<{�a<��a<�a<k�a<ßa< �a<^�a<��a<�a<C�a<p�a<��a<ءa<�a<�a<�a<0�a<I�a<Z�a<Y�a<��a<��a<��a<ޢa<ܢa<�a<!�a<?�a<I�a<d�a<T�a<I�a<6�a<�a<�a<ޢa<Ѣa<��a<��a<e�a<N�a<M�a<7�a<3�a<;�a<K�a<W�a<I�a<Z�a<S�a<X�a<W�a<G�a<E�a<�a<�a<��a<��a<P�a<8�a<�a<Ša<��a<e�a<F�a<)�a<��a<ןa<��a<��a<X�a</�a<Ԟa<��a</�a<�a<��a<�a<Ԝa<l�a<��a<��a<T�a<�a<��a<g�a<*�a<��a<��a<h�a<3�a<Ϙa<��a<7�a<�a<��a<�a<��a<	�a<��a< �a<��a<�a<|�a<�a<g�a<�a<��a<�a<��a<5�a<��a<;�a<��a<�a<��a<֌a<U�a<��a<�a<�a<��a<I�a<Èa<Q�a<هa<d�a<��a<��a<f�a< �a<��a<z�a<�a<�a<��a<S�a<��a<��a<>�a<Ԃa<x�a<)�a<ׁa<x�a<M�a<	�a<ǀa<��a<n�a<U�a<6�a<�a<�a<�a<�a<�a<Qa<a<�~a<�~a<�~a<�~a<_~a<E~a<;~a<L~a<M~a<d~a<�~a<�~a<�~a<a<�  �  �a<�a<�a</�a<G�a<��a<��a<�a<��a<T�a<g�a<��a<�a<�a<��a<��a<4�a<��a<��a<]�a<��a<3�a<��a<�a<\�a<�a<6�a<��a<��a<-�a<��a<��a<t�a<�a<I�a<܊a<Y�a<�a<��a<@�a<܍a<w�a<C�a<��a<��a<�a<��a<+�a<��a<>�a<��a<M�a<��a<?�a<��a<2�a<��a<)�a<җa<:�a<�a<O�a<�a<Z�a<Κa<K�a<��a<�a<D�a<��a<՜a<�a<`�a<z�a<ӝa<��a<D�a<��a<؞a<0�a<i�a<؟a<�a<s�a<Ơa<��a<X�a<^�a<��a<��a<�a<�a<�a<.�a<)�a<P�a<<�a<x�a<w�a<��a<Ģa<âa<�a<��a<,�a<*�a<I�a<E�a<S�a<V�a<'�a<+�a<�a<�a<��a<��a<��a<_�a<j�a<F�a<U�a<M�a<Q�a<r�a<J�a<|�a<j�a<x�a<g�a<5�a<,�a<��a<�a<��a<��a<9�a<�a<�a<��a<��a<D�a<C�a<�a<�a<͟a<��a<y�a<;�a<�a<Þa<��a<G�a<��a<��a<�a<�a<j�a<�a<a<Y�a<�a<��a<��a<.�a<
�a<��a<p�a<O�a<ݘa<��a<4�a<ݗa<h�a<�a<�a<�a<��a<ڔa<v�a<֓a<b�a<�a<S�a<��a<d�a<�a<�a<�a<��a<�a<��a<�a<��a<�a<p�a<��a<�a<��a<�a<r�a<׈a<]�a<߇a<�a<&�a<��a<z�a<�a<Յa<��a<3�a<��a<{�a<C�a<ԃa<~�a<�a<Âa<v�a<	�a<́a<[�a<>�a<�a<��a<��a<U�a<X�a<�a<�a<�a<�a<�a<�a<qa<*a<a<�~a<�~a<�~a<k~a<i~a<L~a<i~a<\~a<�~a<�~a<�~a<a<a<�  �  �a<�a<�a< �a<[�a<��a<��a<�a<�a<1�a<]�a<{�a<āa<�a<K�a<��a<��a<Z�a<ڃa<H�a<��a<+�a<��a<��a<z�a<ˆa<&�a<��a<�a<p�a<��a<�a<��a<��a<{�a<��a<��a<�a<��a<7�a<��a<��a<:�a<ڏa<f�a<�a<��a<'�a<��a<9�a<��a<$�a<��a<�a<��a<�a<��a<+�a<��a<:�a<ʘa<D�a<�a<^�a<Кa<<�a<��a<��a<X�a<��a<�a<<�a<V�a<��a<�a< �a<m�a<��a<�a<G�a<��a<ԟa<G�a<t�a<Ša<��a<3�a<��a<��a<ša<�a<�a<��a<�a<�a<�a<D�a<:�a<a�a<{�a<��a<��a<ܢa<��a<&�a<7�a<C�a<P�a<M�a<1�a<=�a<'�a<�a<�a<��a<Ƣa<��a<��a<~�a<v�a<m�a<{�a<^�a<q�a<��a<y�a<y�a<V�a<X�a<I�a< �a<��a<סa<��a<i�a</�a<�a<��a<��a<W�a<G�a<
�a<�a<ٟa<��a<��a<q�a<F�a<
�a<�a<��a<7�a<��a<��a<a�a<�a<��a<>�a<؛a<��a<;�a<�a<��a<f�a<�a<ݙa<��a<F�a<��a<��a<F�a<ԗa<d�a<�a<z�a<ޕa<a�a<ܔa<;�a<Γa<5�a<��a<U�a<đa<d�a<��a<u�a<�a<��a<�a<��a<%�a<�a<��a<g�a<΋a<G�a<��a<�a<��a<��a<��a<�a<��a<=�a<܆a<v�a<G�a<օa<��a<-�a<ڄa<��a</�a<݃a<|�a<�a<��a<[�a<�a<��a<c�a< �a<Ӏa<��a<b�a<Q�a<-�a<�a<�a<�a<�a<�a<�a<La<@a<a<�~a<�~a<�~a<�~a<�~a<z~a<|~a<�~a<�~a<�~a<�~a<a<\a<�  �  {a<�a<�a<2�a<Y�a<t�a<��a<��a<��a<�a<X�a<{�a<��a<��a<(�a<��a<̂a<k�a<��a<!�a<��a<��a<��a<�a<��a<Նa<B�a<��a<��a<�a<��a<c�a<��a<�a<��a<�a<��a<�a<��a<b�a<�a<��a<6�a<��a<f�a<5�a<��a<'�a<��a<�a<��a<�a<��a<ޔa<i�a<��a<r�a<��a<o�a<H�a<��a<;�a<��a<>�a<՚a<)�a<ӛa<��a<v�a<��a<��a<H�a<v�a<��a<�a<I�a<��a<Ԟa<
�a<N�a<۟a<�a<Q�a<}�a<ڠa<�a<<�a<��a<��a<ȡa<��a<֡a<ߡa<�a<�a<�a<�a<�a<N�a<H�a<z�a<âa<��a<��a<�a<3�a<6�a<G�a<f�a<@�a<\�a<�a<(�a<��a<��a<�a<��a<��a<��a<��a<u�a<��a<��a<|�a<��a<p�a<��a<j�a<i�a<H�a<�a<�a<��a<��a<9�a<*�a<�a<��a<��a<5�a<(�a<۟a<��a<��a<��a<��a<E�a<M�a<��a<�a<��a<S�a<�a<��a<o�a<�a<Ԝa<K�a<�a<��a<K�a<�a<��a<��a<,�a<�a<��a<B�a<�a<��a<g�a<×a<d�a<ߖa<G�a<וa<+�a<�a<�a<��a<%�a<��a<)�a<��a<r�a<��a<k�a<�a<~�a<"�a<��a<C�a<~�a<�a<k�a<܋a<T�a<��a<]�a<��a<#�a<��a<2�a<��a<D�a<$�a<��a<Q�a<߅a<��a<K�a<�a<��a<�a<��a<S�a<��a<��a<2�a<��a<e�a<=�a<��a<��a<j�a<Q�a<T�a<�a<�a<�a<�a<�a<�a<�a<[a<_a<a<
a<�~a<�~a<�~a<�~a<�~a<�~a<�~a<�~a<�~a<a<!a<la<�  �  �a<�a<�a<.�a<J�a<^�a<��a<��a<�a<��a<�a<_�a<��a<΁a<�a<i�a<Ȃa<=�a<��a<�a<��a<�a<��a<�a<n�a<�a<M�a<��a<,�a<��a<�a<^�a<��a<>�a<��a<*�a<ԋa<J�a<�a<��a< �a<Îa<`�a<��a<|�a<�a<��a<�a<��a<��a<��a<ܓa<c�a<ؔa<L�a<֕a<Z�a<ؖa<h�a<�a<x�a<.�a<��a<6�a<��a<'�a<��a<�a<t�a<Ϝa<�a<V�a<��a<�a<�a<s�a<��a<�a<=�a<o�a<ӟa<�a<X�a<��a<�a<�a<J�a<w�a<��a<��a<��a<͡a<ѡa<��a<�a<�a<�a<	�a<"�a<9�a<h�a<{�a<��a<�a<�a<�a<�a<<�a<Z�a<P�a<V�a<L�a<5�a<'�a<�a<�a<עa<٢a<��a<��a<��a<��a<��a<��a<��a<��a<��a<w�a<f�a<8�a<��a<�a<��a<��a<.�a<�a<Ơa<��a<R�a<#�a<��a<ןa<Ɵa<��a<��a<u�a<N�a<,�a<�a<՞a<��a<^�a<�a<֝a<s�a<�a<Μa<a�a<�a<Ǜa<h�a<:�a<֚a<��a<Z�a<�a<��a<l�a<�a<��a<N�a<��a<E�a<͖a<<�a<̕a<�a<��a<�a<�a<�a<��a<�a<��a<+�a<��a<^�a<ޏa<v�a<�a<��a<&�a<��a<�a<��a<�a<b�a<�a<N�a<��a<M�a<��a<C�a<�a<e�a<�a<��a<X�a<�a<��a<P�a<�a<��a<�a<a<Y�a<�a<��a<�a<Ɓa<c�a<�a<πa<��a<[�a<@�a<�a<�a<�a<�a<�a<�a<�a<�a<ka<Ya<<a<a<a<�~a<�~a<�~a<�~a<�~a<�~a<�~a<�~a<"a<Oa<va<�  �  �a<�a<	�a<�a<`�a<|�a<��a<��a<��a<��a<�a<5�a<q�a<��a< �a<;�a<��a<�a<��a<�a<c�a<�a<j�a<�a<o�a<چa<R�a<��a<0�a<��a<�a<_�a<�a<T�a<ъa<i�a<̋a<��a<��a<��a<-�a<ǎa<_�a<�a<��a<��a<��a<�a<��a<��a<R�a<�a<6�a<Ĕa<0�a<��a<0�a<��a<Y�a<Ηa<��a< �a<��a<=�a<��a<M�a<��a<�a<o�a<̜a<$�a<a�a<ʝa<�a<M�a<n�a<ўa<�a<I�a<��a<ҟa<C�a<^�a<��a<�a<�a<N�a<l�a<��a<��a<áa<��a<��a<áa<��a<ѡa<ǡa<�a<�a<#�a<E�a<^�a<��a<��a<��a<�a<1�a<\�a<@�a<a�a<K�a<W�a<6�a<@�a<#�a<�a<�a<آa<�a<âa<עa<ˢa<��a<ʢa<��a<��a<��a<��a<Q�a<N�a<�a<١a<��a<B�a<1�a<ՠa<��a<i�a<"�a<�a<˟a<��a<��a<��a<v�a<A�a<T�a<�a<�a<֞a<��a<c�a<�a<۝a<q�a<K�a<Мa<��a<3�a<�a<��a<2�a<�a<��a<v�a<�a<��a<k�a<
�a<��a<*�a<�a<D�a<іa<7�a<��a<�a<q�a<��a<d�a<ؒa<]�a<�a<��a<��a<��a<0�a<Ϗa<~�a<�a<��a<�a<��a<�a<��a<�a<l�a<�a<S�a<�a<G�a<�a<i�a<�a<��a<�a<�a<^�a<�a<��a<U�a<��a<��a<<�a<��a<`�a<ɂa<n�a<�a<��a<O�a<�a<��a<b�a<E�a<�a<�a<�a<�a<�a<�a<�a<�a<xa<{a<Na<Ga<a<a<�~a<�~a<�~a<�~a<�~a<�~a<a<a</a<na<va<�  �  �a<�a<�a<+�a<M�a<]�a<t�a<��a<��a<��a<��a<�a<O�a<��a<�a<+�a<��a<��a<{�a<�a<^�a<�a<]�a<�a<h�a<�a<m�a<Їa<E�a<��a<�a<{�a<�a<c�a<��a<x�a<�a<��a<�a<��a<C�a<�a<o�a<	�a<��a<�a<��a<�a<z�a<�a<I�a<˓a<6�a<��a<�a<��a<&�a<��a<0�a<̗a<j�a<�a<��a<#�a<��a<8�a<��a<,�a<��a<ݜa<A�a<�a<ǝa<�a<`�a<��a<�a<'�a<Z�a<a<��a<@�a<��a<ʠa<��a<>�a<X�a<k�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<֡a<�a<�a<%�a<_�a<��a<��a<֢a<��a<�a<G�a<Q�a<u�a<i�a<a�a<\�a<F�a<0�a<+�a<�a<��a<��a<�a<ܢa<�a<ʢa<ʢa<Ţa<��a<��a<��a<c�a<;�a<��a<��a<��a<B�a<�a<Рa<��a<G�a<�a<�a<��a<��a<��a<z�a<a�a<;�a<6�a<�a<��a<Ξa<��a<~�a</�a<�a<��a<J�a<�a<��a<C�a<�a<��a<L�a<�a<Ța<u�a<'�a<�a<{�a<%�a<Ƙa<9�a<Ηa</�a<��a<$�a<��a<	�a<p�a<Гa<J�a<Вa<S�a<͑a<Y�a<��a<��a<#�a<��a<c�a<�a<��a<�a<��a<.�a<��a<$�a<��a<��a<z�a<��a<\�a< �a<��a<�a<��a<=�a<�a<��a<,�a<ƅa<s�a<��a<��a<"�a<��a<B�a<a<]�a<��a<��a<*�a<Հa<��a<\�a<&�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<la<Qa<>a< a<a<a<�~a<�~a<�~a<�~a<a<9a<Ca<na<�a<�  �  �a<�a<�a<1�a<H�a<h�a<��a<��a<��a<��a<��a<�a<<�a<��a<a<�a<v�a<�a<S�a<�a<m�a<ׄa<~�a<�a<h�a<�a<H�a<Ňa<>�a<��a<�a<��a<�a<��a<�a<f�a<,�a<��a<+�a<��a<V�a<�a<o�a<��a<w�a<�a<��a<�a<�a<ْa<_�a<��a<!�a<��a<�a<|�a<��a<��a<�a<��a<B�a<�a<��a<!�a<��a<+�a<��a<�a<u�a<ٜa<:�a<��a<ӝa<%�a<`�a<˞a<�a<?�a<��a<��a<�a<D�a<��a<àa<�a<�a<H�a<q�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<աa<�a<�a<D�a<e�a<��a<¢a<�a<)�a<<�a<Y�a<H�a<_�a<_�a<e�a<U�a<K�a<3�a<&�a<7�a<�a<�a<��a<�a<�a<բa<Ңa<��a<��a<m�a<h�a<6�a<�a<ۡa<u�a<Z�a<��a<��a<u�a<4�a<�a<Οa<��a<��a<x�a<R�a<T�a<K�a<�a<(�a<�a<Ξa<��a<Y�a<%�a<�a<��a<P�a<�a<��a<s�a<�a<��a<��a< �a<ؚa<��a<:�a<�a<|�a<�a<��a<H�a<��a<Q�a<��a<�a<��a<ޔa<\�a<��a<8�a<��a<)�a<��a<@�a<�a<m�a<5�a<��a<a�a<	�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<��a<��a<��a<��a<=�a<��a<\�a<�a<��a<%�a<��a<O�a<�a<��a<�a<��a<-�a<̂a<\�a<сa<��a<�a<ʀa<y�a<G�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<ba<ba<Oa<Ha<.a<"a<a<a<$a<�~a<.a<*a<9a<da<ya<�a<�  �  �a< �a<�a<3�a<C�a<a�a<k�a<v�a<��a<��a<�a<�a<<�a<j�a<��a<�a<y�a<ނa<X�a<ԃa<F�a<Ʉa<X�a<�a<a�a<�a<l�a<�a<O�a<��a<)�a<��a<�a<��a<�a<��a<#�a<��a<B�a<ȍa<d�a<�a<��a<�a<��a<�a<��a<��a<V�a<Ēa<7�a<��a<�a<��a<�a<q�a<��a<��a<�a<��a<C�a<��a<l�a<��a<��a<�a<��a<*�a<��a<��a<I�a<��a<�a<5�a<g�a<a<��a<C�a<��a<ɟa<�a<R�a<��a<ՠa<�a<@�a<d�a<h�a<~�a<��a<~�a<}�a<��a<��a<��a<��a<��a<��a<��a<�a<�a<?�a<i�a<��a<��a<�a<�a<:�a<X�a<m�a<y�a<}�a<d�a<b�a<P�a<I�a<2�a<.�a<�a<�a<�a<��a<�a<�a<Ңa<Тa<��a<��a<k�a<1�a<�a<��a<l�a<0�a<��a<��a<k�a<4�a<�a<˟a<��a<��a<g�a<W�a<E�a<#�a<�a<�a<�a<Ǟa<��a<}�a<F�a<��a<��a<\�a<�a<��a<o�a< �a<a<��a<'�a<�a<��a<G�a<�a<��a</�a<��a<=�a<��a<3�a<��a<�a<w�a<�a<M�a<a<6�a<��a<!�a<��a<D�a<Րa<o�a<�a<��a<<�a<�a<|�a<�a<��a<6�a<��a<-�a<��a<�a<��a<�a<��a<�a<��a<4�a<��a<[�a<�a<��a<7�a<߅a<v�a<�a<��a<�a<��a<�a<��a<B�a<Ձa<k�a<�a<��a<r�a<0�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<|a<ma<Ga<<a<'a<"a<a<a<a<'a<3a<Ma<ga<�a<�a<�  �  ;�a<8�a<��a<��a<��a<߁a<�a<�a<�a<Z�a<u�a<��a<܂a<
�a<|�a<��a<$�a<o�a<��a<c�a<��a<Y�a<��a<V�a<��a<B�a<��a<�a<��a<�a<��a<Њa<g�a<ًa<R�a<܌a<_�a<�a<d�a<�a<��a<"�a<��a<�a<ˑa<&�a<ʒa<1�a<��a<�a<f�a<�a<R�a<�a<0�a<֖a<`�a<��a<v�a<ܘa<��a<��a<��a<,�a<��a<H�a<��a<#�a<\�a<�a<=�a<��a<�a<�a<p�a<��a<�a<E�a<��a<Рa<�a<e�a<��a<ϡa<�a<
�a<W�a<`�a<��a<��a<��a<��a<��a<Тa<��a<�a<��a<�a<	�a<&�a<Z�a<n�a<��a<��a<�a<�a<7�a<I�a<O�a<{�a<R�a<�a<n�a<w�a<O�a<J�a<F�a</�a</�a<�a<�a<�a<�a<�a<ߣa<ѣa<��a<��a<j�a<B�a<"�a<עa<��a<A�a<7�a<�a<��a<|�a<7�a<2�a<Πa<ޠa<��a<��a<��a<7�a<O�a<�a<�a<͟a<��a<b�a<*�a<�a<��a<��a<��a<Νa<w�a<"�a<ܜa<��a<>�a<ڛa<��a<I�a<�a<��a<�a<Ιa<5�a<�a<T�a<˗a<5�a<��a<8�a<��a<%�a<h�a<�a<��a<�a<��a< �a<ޑa<J�a<�a<��a<*�a<֏a<6�a<�a<9�a<�a<b�a<݌a<b�a<ċa<Z�a<؊a<l�a<�a<x�a<�a<��a<\�a<�a<��a<�a<��a<W�a<ׅa<��a<�a<��a<�a<̃a<u�a<��a<Ăa<:�a<3�a<فa<��a<��a<`�a<Y�a<�a<'�a<�a<�a<�a<�a<��a<��a<Ҁa<��a<��a<��a<��a<��a<}�a<��a<��a<��a<��a<��a<	�a<�a<�  �  5�a<`�a<��a<��a<��a<ǁa<�a<�a<.�a<D�a<l�a<��a<ׂa<�a<\�a<��a<�a<q�a<ބa<X�a<ۅa<X�a<��a<D�a<��a<E�a<��a<4�a<��a<�a<�a<��a<u�a<ߋa<c�a<ӌa<k�a<�a<��a<�a<��a<�a<��a<?�a<ȑa<9�a<��a<!�a<��a<�a<��a<�a<R�a<֕a<F�a<Öa<I�a<̗a<_�a<ߘa<}�a<�a<��a<)�a<��a<.�a<��a<$�a<��a<�a<-�a<��a<�a<5�a<y�a<��a<��a<H�a<��a<ݠa< �a<U�a<��a<áa<�a<2�a<\�a<m�a<��a<��a<��a<��a<��a<��a<��a<բa<עa<�a<��a<)�a<L�a<k�a<��a<ˣa<�a<�a<#�a<J�a<`�a<w�a<y�a<u�a<`�a<k�a<c�a<Y�a<=�a<:�a<�a<"�a<�a<�a<�a<��a<ԣa<ˣa<��a<��a<t�a<E�a<
�a<Ӣa<��a<l�a<!�a<�a<��a<w�a<5�a<�a<�a<Πa<��a<��a<v�a<g�a<M�a<�a< �a<ٟa<��a<~�a<I�a<��a<��a<l�a<)�a<ܝa<|�a<4�a<Ӝa<��a<>�a<��a<��a<F�a<ٚa<��a<2�a<ʙa<I�a<Ԙa<D�a<Ǘa<L�a<��a<&�a<��a<�a<~�a<��a<��a<�a<��a<"�a<Ǒa<`�a<�a<��a<�a<��a<J�a<�a<g�a<�a<R�a<ߌa<`�a<�a<b�a<�a<`�a<��a<��a<&�a<��a<L�a<�a<|�a<-�a<��a<\�a<�a<{�a<��a<��a<=�a<Ƀa<`�a<��a<��a<T�a<�a<ρa<��a<��a<]�a<F�a<A�a<4�a<�a<�a<�a<��a<�a<ހa<ǀa<��a<��a<��a<��a<�a<��a<z�a<��a<��a<Āa<܀a<��a<�a<�  �  /�a<Z�a<g�a<��a<��a<ԁa<��a<�a<;�a<=�a<��a<��a<�a<)�a<_�a<Ճa<�a<��a<��a<T�a<�a<D�a<چa<I�a<Їa<:�a<��a<#�a<��a<�a<g�a<��a<K�a<��a<`�a<Ȍa<^�a<Ía<u�a<��a<��a<�a<��a<>�a<��a<N�a<��a<<�a<��a<�a<��a<�a<��a<Еa<i�a<Жa<P�a<�a<[�a<�a<��a<�a<��a<$�a<��a<-�a<��a<�a<��a<ޝa<3�a<��a<Ǟa<+�a<M�a<��a<�a<>�a<u�a<��a<�a<>�a<��a<��a<��a<&�a<L�a<�a<��a<��a<��a<��a<��a<ʢa<ߢa<Тa<�a<��a<�a<=�a<L�a<��a<��a<֣a<�a<�a<5�a<O�a<m�a<Z�a<y�a<m�a<v�a<_�a<V�a<G�a<�a<9�a<�a<%�a<�a<��a<��a<�a<�a<ƣa<��a<��a<z�a<O�a<�a<�a<��a<y�a<�a< �a<��a<��a<V�a<�a<�a<͠a<��a<��a<q�a<o�a<:�a<5�a<�a<�a<��a<o�a<8�a<�a<Şa<S�a<"�a<��a<]�a<1�a<Ȝa<��a<�a<�a<��a<E�a<�a<��a<1�a<��a<^�a<јa<_�a<̗a<?�a<��a<'�a<��a<�a<��a<	�a<��a<.�a<��a<S�a<ˑa<c�a<��a<��a<6�a<��a<a�a<ʎa<a�a<ݍa<X�a<�a<E�a<܋a<7�a<׊a<U�a<�a<n�a<��a<��a<5�a<��a<z�a<�a<��a<L�a<��a<}�a<�a<��a<?�a<ȃa<o�a<�a<��a<��a<�a<�a<��a<��a<�a<B�a<L�a<&�a<)�a<�a<�a<�a<׀a<ހa<��a<��a<��a<��a<��a<X�a<��a<p�a<��a<y�a<��a<Հa<�a<�a<�  �  ,�a<K�a<{�a<��a<��a<сa<��a<�a<;�a<W�a<��a<��a<�a<*�a<z�a<ăa<%�a<��a<��a<h�a<��a<[�a<ֆa<@�a<��a<<�a<��a<�a<��a<�a<g�a<؊a<V�a<ʋa<?�a<Ɍa<M�a<ۍa<p�a<��a<z�a<�a<��a<'�a<��a<<�a<��a<3�a<��a<!�a<��a<��a<z�a<�a<]�a<�a<g�a<ߗa<l�a<��a<��a<�a<��a<*�a<��a<!�a<��a<�a<t�a<ޝa<0�a<y�a<ʞa<!�a<b�a<��a<�a<%�a<x�a<��a<��a<=�a<y�a<��a<��a<#�a<T�a<n�a<�a<��a<��a<��a<ɢa<Ѣa<Тa<�a<�a<�a<!�a<=�a<S�a<��a<��a<ӣa<��a<�a<0�a<:�a<\�a<n�a<d�a<k�a<_�a<N�a<G�a<I�a<-�a<�a<�a<�a<��a<��a<�a<գa<ʣa<£a<��a<��a<r�a<<�a<�a<�a<��a<y�a<5�a<��a<��a<��a<W�a<0�a<��a<ߠa<��a<��a<��a<l�a<Q�a<1�a<��a<ןa<��a<u�a<2�a<�a<��a<S�a<�a<��a<h�a<�a<Ȝa<x�a<-�a<�a<��a<,�a<ߚa<��a<�a<��a<L�a<Øa<V�a<˗a<O�a<��a</�a<��a<�a<��a<�a<��a<�a<��a<A�a<ґa<n�a<�a<��a<1�a<��a<J�a<َa<Q�a<ݍa<U�a<Ȍa<H�a<Ӌa<K�a<Ɋa<R�a<Ӊa<q�a<�a<��a<4�a<·a<v�a<�a<��a<U�a<�a<r�a<�a<��a<?�a<ۃa<v�a<�a<��a<k�a<4�a<�a<��a<��a<}�a<Y�a<I�a<<�a<"�a<�a<��a<��a<�a<ɀa<��a<��a<��a<��a<��a<o�a<m�a<w�a<{�a<��a<��a<��a<ڀa<��a<�  �  1�a<?�a<t�a<��a<��a<��a<��a<5�a<1�a<l�a<��a<҂a<�a</�a<��a<Ƀa<_�a<��a<�a<x�a<�a<o�a<͆a<\�a<��a<0�a<��a<�a<��a<܉a<x�a<��a<;�a<��a< �a<��a<"�a<a<3�a<�a<s�a<�a<��a<�a<��a<.�a<Ȓa<A�a<��a<9�a<��a<�a<u�a<�a<u�a<�a<v�a<�a<��a<�a<��a<&�a<��a<?�a<��a<@�a<��a<�a<f�a<ӝa<$�a<k�a<˞a<�a<N�a<~�a<ߟa<�a<X�a<��a<٠a<I�a<c�a<��a<�a<�a<M�a<l�a<��a<��a<Ǣa<âa<Ӣa<�a<�a<#�a<��a</�a<+�a<d�a<��a<��a<��a<Σa<�a<�a<?�a<R�a<N�a<m�a<Y�a<s�a<I�a<P�a<8�a<�a<�a<�a<�a<أa<�a<ңa<ѣa<ޣa<��a<ȣa<��a<��a<c�a<K�a<#�a<�a<΢a<o�a<I�a<�a<�a<��a<]�a<Q�a<�a<�a<ՠa<��a<��a<m�a<d�a<(�a<�a<ٟa<��a<l�a<+�a<��a<��a<d�a<�a<��a<K�a<�a<��a<M�a<�a<��a<��a<$�a<Қa<��a<�a<��a<>�a<�a<d�a<ۗa<g�a<ʖa<O�a<��a<R�a<��a<'�a<��a<-�a<�a<H�a<�a<x�a<�a<��a<8�a<Ώa<@�a<֎a<C�a<Ӎa<I�a<��a<J�a<��a<7�a<��a<G�a<��a<Q�a<��a<w�a<@�a<��a<u�a<�a<��a<M�a<�a<��a<�a<��a<F�a<�a<��a<)�a<��a<s�a<S�a<��a<�a<��a<|�a<q�a<E�a<U�a<#�a<"�a<�a<�a<�a<��a<ŀa<��a<��a<q�a<Q�a<W�a<@�a<r�a<O�a<t�a<��a<��a<�a<�a<�  �  �a<3�a<k�a<��a<��a<��a<�a<%�a<L�a<��a<��a<ɂa<�a<T�a<��a<�a<C�a<��a<)�a<��a<��a<g�a<�a<Y�a<Ça<8�a<��a<��a<}�a<�a<B�a<��a<*�a<��a<�a<��a<�a<��a<3�a<Ɏa<]�a< �a<��a<#�a<��a<=�a<��a<F�a<��a<1�a<��a<=�a<��a<�a<��a<�a<��a<�a<��a<�a<ƙa<8�a<��a<B�a<Ǜa<6�a<��a<�a<s�a<��a<�a<^�a<��a<�a<<�a<w�a<��a<�a<M�a<��a<Ѡa<�a<m�a<��a<Сa<�a<O�a<p�a<��a<��a<��a<ۢa<�a<�a<�a<�a< �a<G�a<K�a<f�a<w�a<��a<�a<�a<�a<1�a<B�a<N�a<]�a<`�a<S�a<R�a<K�a<+�a<$�a<�a<�a<�a<�a<ףa<ݣa<ˣa<��a<��a<��a<��a<��a<��a<q�a<K�a<#�a<��a<��a<��a<k�a<)�a<ءa<��a<��a<g�a<-�a<��a<Ѡa<ՠa<��a<��a<]�a<C�a<�a<ܟa<��a<m�a<�a<ޞa<��a<.�a<۝a<��a<B�a<�a<��a<H�a<
�a<��a<^�a<�a<˚a<d�a<�a<��a<L�a<֘a<i�a<�a<_�a<ߖa<q�a<��a<;�a<Ŕa<D�a<ϓa<S�a<̒a<[�a<�a<��a<�a<��a<B�a<ďa<O�a<Ўa<P�a<��a<A�a<��a<#�a<��a<&�a<��a< �a<��a<F�a<߈a<n�a<�a<a<f�a<�a<��a<O�a<�a<��a<+�a<��a<]�a<��a<��a<,�a<܂a<��a<k�a<�a<�a<��a<��a<��a<`�a<F�a<@�a<%�a<
�a<��a<݀a<��a<��a<��a<g�a<^�a<P�a<Q�a<=�a<A�a<N�a<p�a<�a<��a<��a<�a<�  �  ��a<A�a<`�a<��a<��a<�a<�a<&�a<q�a<{�a<Ăa<�a<3�a<u�a<��a<�a<d�a<ʄa<1�a<��a<�a<h�a<��a<N�a<Ňa<(�a<��a<�a<[�a<ىa<%�a<��a<�a<��a<�a<n�a<�a<��a<)�a<��a<I�a<��a<v�a<+�a<��a<8�a<��a<U�a<Ǔa<D�a<Ĕa<$�a<��a<'�a<��a<�a<��a<@�a<��a<=�a<��a<J�a<ؚa<G�a<ڛa<(�a<��a<��a<w�a<��a<�a<L�a<��a<۞a<�a<s�a<��a<�a<A�a<x�a<Ƞa<��a<[�a<��a<ܡa<�a<:�a<r�a<��a<ɢa<âa<��a<�a<�a<�a<"�a<J�a<<�a<k�a<��a<��a<ţa<ͣa<
�a<	�a<9�a<J�a<J�a<V�a<O�a<^�a<6�a<H�a<�a<�a<��a<�a<�a<��a<ƣa<��a<��a<��a<��a<��a<��a<��a<~�a<f�a<G�a<)�a<
�a<��a<��a<X�a<<�a<��a<ӡa<��a<X�a<U�a<�a<��a<ܠa<��a<��a<^�a<Q�a<
�a<ݟa<��a<h�a<�a<��a<��a<�a<ҝa<u�a</�a<Ҝa<n�a<C�a<ݛa<��a<I�a<��a<Ța<V�a<�a<��a<H�a<Ϙa<x�a<�a<r�a<��a<X�a<�a<]�a<�a<V�a<Փa<|�a<�a<��a< �a<��a<6�a<��a<U�a<��a<I�a<��a<T�a<��a<:�a<��a<	�a<��a<��a<��a<��a<��a<:�a<��a<e�a<�a<��a<L�a<��a<��a<:�a<�a<}�a<<�a<��a<}�a<��a<��a<[�a<��a<ǂa<`�a<;�a<�a<Ձa<��a<~�a<��a<I�a<H�a<-�a<�a<��a<̀a<Àa<��a<��a<P�a<L�a<7�a<*�a<2�a<�a<=�a<N�a<b�a<��a<��a<�a<�  �  �a<1�a<]�a<��a<Áa<�a<�a<H�a<x�a<��a<ςa<�a<S�a<��a<уa<%�a<��a<�a<B�a<��a<�a<��a<�a<a�a<ʇa<.�a<��a<�a<S�a<��a<=�a<��a<�a<h�a<�a<u�a<�a<l�a<��a<��a<?�a<ޏa<q�a<�a<��a<6�a<̒a<T�a<��a<X�a<Քa<C�a<��a<H�a<��a<>�a<��a<E�a<Әa<G�a<әa<\�a<�a<J�a<כa<D�a<��a<�a<d�a<��a<��a<;�a<��a<��a<��a<H�a<��a<Οa<�a<T�a<��a<�a<D�a<��a<֡a<�a<A�a<w�a<��a<��a<עa<��a<�a<�a<*�a<O�a<R�a<d�a<��a<��a<��a<ͣa<�a<�a<-�a<*�a<P�a<Z�a<V�a<V�a<P�a<4�a<&�a<�a<	�a<Уa<ȣa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<z�a<h�a<T�a<2�a<��a<�a<��a<s�a<G�a<�a<�a<��a<��a<`�a<I�a<�a<�a<��a<��a<y�a<G�a<�a<�a<��a<_�a<�a<��a<d�a<*�a<��a<O�a<�a<��a<t�a<�a<��a<t�a<M�a<�a<��a<Q�a<�a<��a<F�a<�a<w�a<�a<��a<�a<w�a<�a<�a<��a<v�a<��a<��a<�a<��a<�a<��a<A�a<��a<R�a<ҏa<L�a<Ďa<B�a<��a<�a<��a<�a<f�a<ߊa<o�a<��a<|�a<�a<��a<>�a<�a<��a<=�a<��a<��a<A�a<�a<��a<4�a<τa<��a<�a<��a<g�a<*�a<ςa<��a<S�a<'�a<�a<��a<��a<��a<n�a<9�a<2�a<�a<��a<Ҁa<��a<��a<k�a<[�a<C�a<�a<
�a<�a< �a<�a<,�a<;�a<|�a<��a<Āa<�  �  �a<�a<^�a<��a<��a<��a<�a<d�a<o�a<ǂa<��a<�a<X�a<��a<��a<'�a<��a<߄a<X�a<ąa<�a<��a<��a<n�a<��a<5�a<��a<�a<b�a<��a<�a<i�a<��a<a�a<ċa<\�a<a<��a<��a<��a<,�a<ʏa<v�a<�a<��a</�a<˒a<I�a<ޓa<d�a<ϔa<r�a<Õa<X�a<̖a<T�a<ߗa<N�a<�a<K�a<��a<b�a<�a<g�a<ɛa<H�a<��a<�a<V�a<��a<�a<+�a<z�a<��a<�a< �a<v�a<��a<�a<h�a<��a<�a<.�a<��a<��a<�a<M�a<h�a<��a<��a<��a<�a<�a<5�a<'�a<X�a<U�a<��a<��a<��a<ɣa<ߣa<!�a<�a<E�a<B�a<R�a<O�a<S�a<Y�a<5�a<>�a<�a<�a<�a<գa<ܣa<��a<��a<}�a<��a<��a<}�a<��a<t�a<��a<r�a<|�a<g�a<H�a<9�a<�a<��a<��a<��a<Y�a<$�a<��a<��a<��a<a�a<O�a<�a<�a<�a<��a<��a<K�a<*�a<ԟa<��a<[�a<��a<Þa<K�a<�a<��a<^�a<��a<��a<[�a<�a<��a<k�a<4�a<ޚa<��a<V�a<��a<��a<?�a<�a<l�a<�a<��a<�a<��a<��a<��a<�a<��a<�a<��a<$�a<��a<F�a<��a<I�a<Ґa<D�a<׏a<?�a<͎a<4�a<��a<�a<{�a<��a<W�a<��a<F�a<މa<_�a<��a<��a<'�a<�a<��a<H�a<�a<��a<M�a<߅a<��a<.�a<��a<��a<.�a<ڃa<e�a<3�a<҂a<��a<W�a<.�a< �a<сa<Ӂa<��a<��a<Q�a<5�a<�a<�a<րa<��a<��a<O�a<>�a<"�a<�a<�a<�a<
�a<�a<4�a<B�a<W�a<��a<��a<�  �  �a<�a<N�a<��a<Ła<��a<%�a<]�a<��a<��a<��a<=�a<n�a<��a<�a<T�a<��a<�a<f�a<Ņa<2�a<��a<��a<m�a<ɇa<�a<��a<�a<I�a<��a<��a<o�a<Ċa<?�a<��a<?�a<��a<N�a<ݍa<��a<#�a<��a<d�a<�a<��a<5�a<ђa<W�a<�a<j�a<�a<h�a<�a<o�a<�a<b�a<�a<p�a<��a<��a<��a<r�a<��a<t�a<؛a<K�a<��a<�a<S�a<��a<ݝa<!�a<[�a<��a<Ԟa<�a<c�a<��a<�a</�a<��a<Ѡa<%�a<w�a<��a<��a<-�a<u�a<��a<Ȣa<��a<�a<!�a<>�a<e�a<q�a<��a<��a<��a<ǣa<�a<��a<�a<"�a<>�a<I�a<[�a<]�a<N�a<B�a<>�a<+�a<�a<�a<أa<��a<��a<��a<��a<x�a<s�a<i�a<s�a<t�a<~�a<��a<y�a<k�a<[�a<V�a<A�a<�a<��a<Ţa<��a<n�a<K�a<�a<�a<��a<��a<g�a<K�a<�a<�a<��a<��a<V�a<)�a<�a<��a<K�a<��a<��a<K�a<�a<��a<+�a<ܜa<��a<?�a<�a<��a<S�a<�a<՚a<��a<D�a<��a<��a<E�a<�a<z�a<�a<��a<�a<��a<#�a<��a<%�a<��a<$�a<��a<7�a<Ēa<A�a<őa<T�a<ߐa<S�a<ُa<H�a<��a<0�a<��a<�a<p�a<ًa<J�a<��a<7�a<ˉa<V�a<�a<x�a<-�a<ȇa<z�a<0�a<Նa<��a<-�a<�a<��a<;�a<�a<��a<2�a<�a<��a<L�a<��a<��a<z�a<H�a< �a<�a<��a<��a<~�a<Y�a<>�a<�a<�a<��a<��a<}�a<T�a<-�a<�a<�a<�a<�a<�a<�a<�a<�a<L�a<x�a<��a<�  �  рa< �a<Q�a<��a<ˁa<�a<3�a<a�a<��a<Âa<�a<5�a<_�a<؃a<�a<l�a<��a<�a<q�a<ׅa<C�a<��a<�a<Z�a<ۇa<-�a<��a<�a<5�a<��a<�a<q�a<��a<A�a<��a<&�a<Ќa<<�a<�a<y�a<�a<��a<R�a<�a<��a<F�a<ǒa<\�a<�a<m�a<�a<g�a<�a<^�a<�a<v�a<�a<z�a<�a<��a<��a<��a<��a<s�a<�a<>�a<��a<��a<W�a<��a<՝a<�a<S�a<��a<Ğa<'�a<K�a<��a<�a<�a<��a<Ša<&�a<f�a<��a<�a<>�a<��a<��a<ߢa<��a<�a<8�a<A�a<g�a<W�a<��a<��a<Σa<��a<ݣa<�a<�a<J�a<B�a<S�a<Q�a<]�a<`�a<H�a<A�a<�a<�a<ڣa<ףa<��a<��a<��a<m�a<|�a<i�a<m�a<w�a<Z�a<~�a<g�a<}�a<o�a<p�a<[�a<0�a<$�a<��a<�a<��a<��a<D�a< �a<�a<��a<��a<O�a<K�a<�a<��a<Рa<��a<k�a<�a<�a<��a<Q�a<��a<��a<N�a<՝a<��a<�a<ޜa<}�a<&�a<��a<��a<c�a<�a<Ěa<��a<2�a<��a<��a<V�a<�a<�a<�a<��a<@�a<��a<<�a<��a<&�a<��a<-�a<��a<$�a<Ԓa<>�a<�a<X�a<ސa<_�a<̏a<_�a<��a<4�a<��a<��a<c�a<ыa<\�a<��a<M�a<��a<C�a<�a<g�a<3�a<��a<{�a<�a<؆a<��a<>�a<��a<��a<R�a<�a<��a<I�a<�a<��a<2�a<�a<��a<��a<;�a<�a<�a<Áa<��a<��a<b�a<3�a<�a<��a<ŀa<��a<c�a<U�a<�a<�a<�a<�a<�a<�a<�a<�a<!�a<Q�a<_�a<��a<�  �  �a<�a<G�a<��a<ȁa<�a<<�a<f�a<��a<ڂa<�a<R�a<��a<Ճa<�a<p�a<��a<&�a<��a<�a</�a<��a<�a<w�a<͇a<+�a<x�a<ֈa<C�a<��a<�a<K�a<��a<*�a<��a<!�a<��a<A�a<ʍa<n�a<�a<��a<a�a<�a<��a<2�a<ےa<g�a<��a<m�a<��a<�a<�a<��a<�a<��a<��a<��a<�a<��a<�a<��a<��a<��a<�a<V�a<��a<��a<8�a<��a<ߝa<�a<L�a<|�a<Ȟa<��a<E�a<��a<ҟa<&�a<h�a<Ǡa< �a<r�a<��a<�a<@�a<t�a<��a<ߢa<�a<�a<=�a<Z�a<t�a<�a<��a<��a<ͣa<ۣa<�a<�a<*�a<0�a<H�a<c�a<c�a<d�a<R�a<B�a<$�a<%�a<�a<�a<��a<��a<��a<q�a<j�a<X�a<`�a<X�a<\�a<a�a<q�a<y�a<d�a<d�a<c�a<Y�a<I�a<-�a< �a<Тa<��a<��a<`�a<$�a<�a<��a<��a<v�a<[�a</�a<��a<��a<��a<j�a<3�a<�a<��a<>�a<�a<��a<E�a<ٝa<v�a<"�a<ǜa<g�a<!�a<Λa<��a<?�a<�a<Ěa<��a<B�a<ޙa<��a<B�a<��a<��a<#�a<��a<*�a<��a<C�a<Õa<9�a<��a<8�a<Ǔa<R�a<ܒa<X�a<ܑa<T�a<�a<g�a<�a<G�a<��a<�a<��a<�a<`�a<ˋa<.�a<��a<#�a<��a<2�a<ˈa<n�a<�a<��a<u�a<+�a<Άa<}�a<@�a<�a<��a<Q�a<��a<��a<N�a<��a<��a<Z�a<�a<Ƃa<��a<\�a<:�a<�a<܁a<��a<��a<r�a<F�a< �a<�a<��a<��a<w�a<L�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<6�a<f�a<��a<�  �  ��a<�a<^�a<��a<��a<��a<�a<m�a<��a<�a<�a<G�a<��a<Ãa<�a<e�a<Ąa<�a<r�a<�a<?�a<��a<�a<{�a<��a<*�a<��a<؈a<1�a<r�a<��a<N�a<ϊa<"�a<��a<=�a<��a<U�a<ča<��a<�a<��a<d�a<�a<��a<&�a<Ւa<;�a<�a<z�a<��a<��a<�a<��a<��a<��a<�a<|�a<	�a<q�a<�a<��a<�a<t�a<��a<S�a<��a<�a<H�a<��a<��a<��a<e�a<y�a<ݞa<��a<_�a<��a<��a<<�a<g�a<٠a<��a<]�a<��a<��a<I�a<a�a<��a<��a<�a<�a<B�a<Q�a<Y�a<��a<��a<��a<��a<ڣa<��a<�a<>�a<:�a<R�a<A�a<N�a<a�a<I�a<U�a<&�a<'�a<٣a<�a<ͣa<��a<��a<a�a<��a<T�a<j�a<[�a<h�a<w�a<G�a<v�a<h�a<{�a<^�a<R�a<C�a<�a<�a<ۢa<ʢa<i�a<V�a<)�a<�a<ԡa<��a<~�a<H�a<�a<�a<ˠa<��a<@�a<7�a<џa<��a<O�a<�a<��a<�a<�a<y�a<5�a<��a<u�a<=�a<��a<��a<:�a<�a<��a<`�a<D�a<�a<��a<6�a<�a<^�a<�a<��a<)�a<��a<�a<��a<+�a<��a<E�a<��a<H�a<��a<]�a<ّa<b�a<ߐa<9�a<�a<5�a<Վa<%�a<��a<��a<O�a<�a<+�a<Ǌa<�a<Ɖa<D�a<��a<��a<�a<Їa<O�a<�a<цa<��a<I�a<؅a<��a<&�a< �a<��a<S�a<��a<��a<]�a<�a<тa<��a<[�a<-�a<�a<��a<��a<��a<P�a<1�a<�a<�a<Ҁa<��a<y�a<�a<+�a<�a<�a<�a<�a<�a<�a<�a<�a<A�a<|�a<{�a<�  �  �a<�a<G�a<��a<ȁa<�a<<�a<f�a<��a<ڂa<�a<R�a<��a<Ճa<�a<p�a<��a<&�a<��a<�a</�a<��a<�a<w�a<͇a<+�a<x�a<ֈa<C�a<��a<�a<K�a<��a<*�a<��a<!�a<��a<A�a<ʍa<n�a<�a<��a<a�a<�a<��a<2�a<ےa<g�a<��a<m�a<��a<�a<�a<��a<�a<��a<��a<��a<�a<��a<�a<��a<��a<��a<�a<V�a<��a<��a<8�a<��a<ߝa<�a<L�a<|�a<Ȟa<��a<E�a<��a<ҟa<&�a<h�a<Ǡa< �a<r�a<��a<�a<@�a<t�a<��a<ߢa<�a<�a<=�a<Z�a<t�a<�a<��a<��a<ͣa<ۣa<�a<�a<*�a<0�a<H�a<c�a<c�a<d�a<R�a<B�a<$�a<%�a<�a<�a<��a<��a<��a<q�a<j�a<X�a<`�a<X�a<\�a<a�a<q�a<y�a<d�a<d�a<c�a<Y�a<I�a<-�a< �a<Тa<��a<��a<`�a<$�a<�a<��a<��a<v�a<[�a</�a<��a<��a<��a<j�a<3�a<�a<��a<>�a<�a<��a<E�a<ٝa<v�a<"�a<ǜa<g�a<!�a<Λa<��a<?�a<�a<Ěa<��a<B�a<ޙa<��a<B�a<��a<��a<#�a<��a<*�a<��a<C�a<Õa<9�a<��a<8�a<Ǔa<R�a<ܒa<X�a<ܑa<T�a<�a<g�a<�a<G�a<��a<�a<��a<�a<`�a<ˋa<.�a<��a<#�a<��a<2�a<ˈa<n�a<�a<��a<u�a<+�a<Άa<}�a<@�a<�a<��a<Q�a<��a<��a<N�a<��a<��a<Z�a<�a<Ƃa<��a<\�a<:�a<�a<܁a<��a<��a<r�a<F�a< �a<�a<��a<��a<w�a<L�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<6�a<f�a<��a<�  �  рa< �a<Q�a<��a<ˁa<�a<3�a<a�a<��a<Âa<�a<5�a<_�a<؃a<�a<l�a<��a<�a<q�a<ׅa<C�a<��a<�a<Z�a<ۇa<-�a<��a<�a<5�a<��a<�a<q�a<��a<A�a<��a<&�a<Ќa<<�a<�a<y�a<�a<��a<R�a<�a<��a<F�a<ǒa<\�a<�a<m�a<�a<g�a<�a<^�a<�a<v�a<�a<z�a<�a<��a<��a<��a<��a<s�a<�a<>�a<��a<��a<W�a<��a<՝a<�a<S�a<��a<Ğa<'�a<K�a<��a<�a<�a<��a<Ša<&�a<f�a<��a<�a<>�a<��a<��a<ߢa<��a<�a<8�a<A�a<g�a<W�a<��a<��a<Σa<��a<ݣa<�a<�a<J�a<B�a<S�a<Q�a<]�a<`�a<H�a<A�a<�a<�a<ڣa<ףa<��a<��a<��a<m�a<|�a<i�a<m�a<w�a<Z�a<~�a<g�a<}�a<o�a<p�a<[�a<0�a<$�a<��a<�a<��a<��a<D�a< �a<�a<��a<��a<O�a<K�a<�a<��a<Рa<��a<k�a<�a<�a<��a<Q�a<��a<��a<N�a<՝a<��a<�a<ޜa<}�a<&�a<��a<��a<c�a<�a<Ěa<��a<2�a<��a<��a<V�a<�a<�a<�a<��a<@�a<��a<<�a<��a<&�a<��a<-�a<��a<$�a<Ԓa<>�a<�a<X�a<ސa<_�a<̏a<_�a<��a<4�a<��a<��a<c�a<ыa<\�a<��a<M�a<��a<C�a<�a<g�a<3�a<��a<{�a<�a<؆a<��a<>�a<��a<��a<R�a<�a<��a<I�a<�a<��a<2�a<�a<��a<��a<;�a<�a<�a<Áa<��a<��a<b�a<3�a<�a<��a<ŀa<��a<c�a<U�a<�a<�a<�a<�a<�a<�a<�a<�a<!�a<Q�a<_�a<��a<�  �  �a<�a<N�a<��a<Ła<��a<%�a<]�a<��a<��a<��a<=�a<n�a<��a<�a<T�a<��a<�a<f�a<Ņa<2�a<��a<��a<m�a<ɇa<�a<��a<�a<I�a<��a<��a<o�a<Ċa<?�a<��a<?�a<��a<N�a<ݍa<��a<#�a<��a<d�a<�a<��a<5�a<ђa<W�a<�a<j�a<�a<h�a<�a<o�a<�a<b�a<�a<p�a<��a<��a<��a<r�a<��a<t�a<؛a<K�a<��a<�a<S�a<��a<ݝa<!�a<[�a<��a<Ԟa<�a<c�a<��a<�a</�a<��a<Ѡa<%�a<w�a<��a<��a<-�a<u�a<��a<Ȣa<��a<�a<!�a<>�a<e�a<q�a<��a<��a<��a<ǣa<�a<��a<�a<"�a<>�a<I�a<[�a<]�a<N�a<B�a<>�a<+�a<�a<�a<أa<��a<��a<��a<��a<x�a<s�a<i�a<s�a<t�a<~�a<��a<y�a<k�a<[�a<V�a<A�a<�a<��a<Ţa<��a<n�a<K�a<�a<�a<��a<��a<g�a<K�a<�a<�a<��a<��a<V�a<)�a<�a<��a<K�a<��a<��a<K�a<�a<��a<+�a<ܜa<��a<?�a<�a<��a<S�a<�a<՚a<��a<D�a<��a<��a<E�a<�a<z�a<�a<��a<�a<��a<#�a<��a<%�a<��a<$�a<��a<7�a<Ēa<A�a<őa<T�a<ߐa<S�a<ُa<H�a<��a<0�a<��a<�a<p�a<ًa<J�a<��a<7�a<ˉa<V�a<�a<x�a<-�a<ȇa<z�a<0�a<Նa<��a<-�a<�a<��a<;�a<�a<��a<2�a<�a<��a<L�a<��a<��a<z�a<H�a< �a<�a<��a<��a<~�a<Y�a<>�a<�a<�a<��a<��a<}�a<T�a<-�a<�a<�a<�a<�a<�a<�a<�a<�a<L�a<x�a<��a<�  �  �a<�a<^�a<��a<��a<��a<�a<d�a<o�a<ǂa<��a<�a<X�a<��a<��a<'�a<��a<߄a<X�a<ąa<�a<��a<��a<n�a<��a<5�a<��a<�a<b�a<��a<�a<i�a<��a<a�a<ċa<\�a<a<��a<��a<��a<,�a<ʏa<v�a<�a<��a</�a<˒a<I�a<ޓa<d�a<ϔa<r�a<Õa<X�a<̖a<T�a<ߗa<N�a<�a<K�a<��a<b�a<�a<g�a<ɛa<H�a<��a<�a<V�a<��a<�a<+�a<z�a<��a<�a< �a<v�a<��a<�a<h�a<��a<�a<.�a<��a<��a<�a<M�a<h�a<��a<��a<��a<�a<�a<5�a<'�a<X�a<U�a<��a<��a<��a<ɣa<ߣa<!�a<�a<E�a<B�a<R�a<O�a<S�a<Y�a<5�a<>�a<�a<�a<�a<գa<ܣa<��a<��a<}�a<��a<��a<}�a<��a<t�a<��a<r�a<|�a<g�a<H�a<9�a<�a<��a<��a<��a<Y�a<$�a<��a<��a<��a<a�a<O�a<�a<�a<�a<��a<��a<K�a<*�a<ԟa<��a<[�a<��a<Þa<K�a<�a<��a<^�a<��a<��a<[�a<�a<��a<k�a<4�a<ޚa<��a<V�a<��a<��a<?�a<�a<l�a<�a<��a<�a<��a<��a<��a<�a<��a<�a<��a<$�a<��a<F�a<��a<I�a<Ґa<D�a<׏a<?�a<͎a<4�a<��a<�a<{�a<��a<W�a<��a<F�a<މa<_�a<��a<��a<'�a<�a<��a<H�a<�a<��a<M�a<߅a<��a<.�a<��a<��a<.�a<ڃa<e�a<3�a<҂a<��a<W�a<.�a< �a<сa<Ӂa<��a<��a<Q�a<5�a<�a<�a<րa<��a<��a<O�a<>�a<"�a<�a<�a<�a<
�a<�a<4�a<B�a<W�a<��a<��a<�  �  �a<1�a<]�a<��a<Áa<�a<�a<H�a<x�a<��a<ςa<�a<S�a<��a<уa<%�a<��a<�a<B�a<��a<�a<��a<�a<a�a<ʇa<.�a<��a<�a<S�a<��a<=�a<��a<�a<h�a<�a<u�a<�a<l�a<��a<��a<?�a<ޏa<q�a<�a<��a<6�a<̒a<T�a<��a<X�a<Քa<C�a<��a<H�a<��a<>�a<��a<E�a<Әa<G�a<әa<\�a<�a<J�a<כa<D�a<��a<�a<d�a<��a<��a<;�a<��a<��a<��a<H�a<��a<Οa<�a<T�a<��a<�a<D�a<��a<֡a<�a<A�a<w�a<��a<��a<עa<��a<�a<�a<*�a<O�a<R�a<d�a<��a<��a<��a<ͣa<�a<�a<-�a<*�a<P�a<Z�a<V�a<V�a<P�a<4�a<&�a<�a<	�a<Уa<ȣa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<z�a<h�a<T�a<2�a<��a<�a<��a<s�a<G�a<�a<�a<��a<��a<`�a<I�a<�a<�a<��a<��a<y�a<G�a<�a<�a<��a<_�a<�a<��a<d�a<*�a<��a<O�a<�a<��a<t�a<�a<��a<t�a<M�a<�a<��a<Q�a<�a<��a<F�a<�a<w�a<�a<��a<�a<w�a<�a<�a<��a<v�a<��a<��a<�a<��a<�a<��a<A�a<��a<R�a<ҏa<L�a<Ďa<B�a<��a<�a<��a<�a<f�a<ߊa<o�a<��a<|�a<�a<��a<>�a<�a<��a<=�a<��a<��a<A�a<�a<��a<4�a<τa<��a<�a<��a<g�a<*�a<ςa<��a<S�a<'�a<�a<��a<��a<��a<n�a<9�a<2�a<�a<��a<Ҁa<��a<��a<k�a<[�a<C�a<�a<
�a<�a< �a<�a<,�a<;�a<|�a<��a<Āa<�  �  ��a<A�a<`�a<��a<��a<�a<�a<&�a<q�a<{�a<Ăa<�a<3�a<u�a<��a<�a<d�a<ʄa<1�a<��a<�a<h�a<��a<N�a<Ňa<(�a<��a<�a<[�a<ىa<%�a<��a<�a<��a<�a<n�a<�a<��a<)�a<��a<I�a<��a<v�a<+�a<��a<8�a<��a<U�a<Ǔa<D�a<Ĕa<$�a<��a<'�a<��a<�a<��a<@�a<��a<=�a<��a<J�a<ؚa<G�a<ڛa<(�a<��a<��a<w�a<��a<�a<L�a<��a<۞a<�a<s�a<��a<�a<A�a<x�a<Ƞa<��a<[�a<��a<ܡa<�a<:�a<r�a<��a<ɢa<âa<��a<�a<�a<�a<"�a<J�a<<�a<k�a<��a<��a<ţa<ͣa<
�a<	�a<9�a<J�a<J�a<V�a<O�a<^�a<6�a<H�a<�a<�a<��a<�a<�a<��a<ƣa<��a<��a<��a<��a<��a<��a<��a<~�a<f�a<G�a<)�a<
�a<��a<��a<X�a<<�a<��a<ӡa<��a<X�a<U�a<�a<��a<ܠa<��a<��a<^�a<Q�a<
�a<ݟa<��a<h�a<�a<��a<��a<�a<ҝa<u�a</�a<Ҝa<n�a<C�a<ݛa<��a<I�a<��a<Ța<V�a<�a<��a<H�a<Ϙa<x�a<�a<r�a<��a<X�a<�a<]�a<�a<V�a<Փa<|�a<�a<��a< �a<��a<6�a<��a<U�a<��a<I�a<��a<T�a<��a<:�a<��a<	�a<��a<��a<��a<��a<��a<:�a<��a<e�a<�a<��a<L�a<��a<��a<:�a<�a<}�a<<�a<��a<}�a<��a<��a<[�a<��a<ǂa<`�a<;�a<�a<Ձa<��a<~�a<��a<I�a<H�a<-�a<�a<��a<̀a<Àa<��a<��a<P�a<L�a<7�a<*�a<2�a<�a<=�a<N�a<b�a<��a<��a<�a<�  �  �a<3�a<k�a<��a<��a<��a<�a<%�a<L�a<��a<��a<ɂa<�a<T�a<��a<�a<C�a<��a<)�a<��a<��a<g�a<�a<Y�a<Ça<8�a<��a<��a<}�a<�a<B�a<��a<*�a<��a<�a<��a<�a<��a<3�a<Ɏa<]�a< �a<��a<#�a<��a<=�a<��a<F�a<��a<1�a<��a<=�a<��a<�a<��a<�a<��a<�a<��a<�a<ƙa<8�a<��a<B�a<Ǜa<6�a<��a<�a<s�a<��a<�a<^�a<��a<�a<<�a<w�a<��a<�a<M�a<��a<Ѡa<�a<m�a<��a<Сa<�a<O�a<p�a<��a<��a<��a<ۢa<�a<�a<�a<�a< �a<G�a<K�a<f�a<w�a<��a<�a<�a<�a<1�a<B�a<N�a<]�a<`�a<S�a<R�a<K�a<+�a<$�a<�a<�a<�a<�a<ףa<ݣa<ˣa<��a<��a<��a<��a<��a<��a<q�a<K�a<#�a<��a<��a<��a<k�a<)�a<ءa<��a<��a<g�a<-�a<��a<Ѡa<ՠa<��a<��a<]�a<C�a<�a<ܟa<��a<m�a<�a<ޞa<��a<.�a<۝a<��a<B�a<�a<��a<H�a<
�a<��a<^�a<�a<˚a<d�a<�a<��a<L�a<֘a<i�a<�a<_�a<ߖa<q�a<��a<;�a<Ŕa<D�a<ϓa<S�a<̒a<[�a<�a<��a<�a<��a<B�a<ďa<O�a<Ўa<P�a<��a<A�a<��a<#�a<��a<&�a<��a< �a<��a<F�a<߈a<n�a<�a<a<f�a<�a<��a<O�a<�a<��a<+�a<��a<]�a<��a<��a<,�a<܂a<��a<k�a<�a<�a<��a<��a<��a<`�a<F�a<@�a<%�a<
�a<��a<݀a<��a<��a<��a<g�a<^�a<P�a<Q�a<=�a<A�a<N�a<p�a<�a<��a<��a<�a<�  �  1�a<?�a<t�a<��a<��a<��a<��a<5�a<1�a<l�a<��a<҂a<�a</�a<��a<Ƀa<_�a<��a<�a<x�a<�a<o�a<͆a<\�a<��a<0�a<��a<�a<��a<܉a<x�a<��a<;�a<��a< �a<��a<"�a<a<3�a<�a<s�a<�a<��a<�a<��a<.�a<Ȓa<A�a<��a<9�a<��a<�a<u�a<�a<u�a<�a<v�a<�a<��a<�a<��a<&�a<��a<?�a<��a<@�a<��a<�a<f�a<ӝa<$�a<k�a<˞a<�a<N�a<~�a<ߟa<�a<X�a<��a<٠a<I�a<c�a<��a<�a<�a<M�a<l�a<��a<��a<Ǣa<âa<Ӣa<�a<�a<#�a<��a</�a<+�a<d�a<��a<��a<��a<Σa<�a<�a<?�a<R�a<N�a<m�a<Y�a<s�a<I�a<P�a<8�a<�a<�a<�a<�a<أa<�a<ңa<ѣa<ޣa<��a<ȣa<��a<��a<c�a<K�a<#�a<�a<΢a<o�a<I�a<�a<�a<��a<]�a<Q�a<�a<�a<ՠa<��a<��a<m�a<d�a<(�a<�a<ٟa<��a<l�a<+�a<��a<��a<d�a<�a<��a<K�a<�a<��a<M�a<�a<��a<��a<$�a<Қa<��a<�a<��a<>�a<�a<d�a<ۗa<g�a<ʖa<O�a<��a<R�a<��a<'�a<��a<-�a<�a<H�a<�a<x�a<�a<��a<8�a<Ώa<@�a<֎a<C�a<Ӎa<I�a<��a<J�a<��a<7�a<��a<G�a<��a<Q�a<��a<w�a<@�a<��a<u�a<�a<��a<M�a<�a<��a<�a<��a<F�a<�a<��a<)�a<��a<s�a<S�a<��a<�a<��a<|�a<q�a<E�a<U�a<#�a<"�a<�a<�a<�a<��a<ŀa<��a<��a<q�a<Q�a<W�a<@�a<r�a<O�a<t�a<��a<��a<�a<�a<�  �  ,�a<K�a<{�a<��a<��a<сa<��a<�a<;�a<W�a<��a<��a<�a<*�a<z�a<ăa<%�a<��a<��a<h�a<��a<[�a<ֆa<@�a<��a<<�a<��a<�a<��a<�a<g�a<؊a<V�a<ʋa<?�a<Ɍa<M�a<ۍa<p�a<��a<z�a<�a<��a<'�a<��a<<�a<��a<3�a<��a<!�a<��a<��a<z�a<�a<]�a<�a<g�a<ߗa<l�a<��a<��a<�a<��a<*�a<��a<!�a<��a<�a<t�a<ޝa<0�a<y�a<ʞa<!�a<b�a<��a<�a<%�a<x�a<��a<��a<=�a<y�a<��a<��a<#�a<T�a<n�a<�a<��a<��a<��a<ɢa<Ѣa<Тa<�a<�a<�a<!�a<=�a<S�a<��a<��a<ӣa<��a<�a<0�a<:�a<\�a<n�a<d�a<k�a<_�a<N�a<G�a<I�a<-�a<�a<�a<�a<��a<��a<�a<գa<ʣa<£a<��a<��a<r�a<<�a<�a<�a<��a<y�a<5�a<��a<��a<��a<W�a<0�a<��a<ߠa<��a<��a<��a<l�a<Q�a<1�a<��a<ןa<��a<u�a<2�a<�a<��a<S�a<�a<��a<h�a<�a<Ȝa<x�a<-�a<�a<��a<,�a<ߚa<��a<�a<��a<L�a<Øa<V�a<˗a<O�a<��a</�a<��a<�a<��a<�a<��a<�a<��a<A�a<ґa<n�a<�a<��a<1�a<��a<J�a<َa<Q�a<ݍa<U�a<Ȍa<H�a<Ӌa<K�a<Ɋa<R�a<Ӊa<q�a<�a<��a<4�a<·a<v�a<�a<��a<U�a<�a<r�a<�a<��a<?�a<ۃa<v�a<�a<��a<k�a<4�a<�a<��a<��a<}�a<Y�a<I�a<<�a<"�a<�a<��a<��a<�a<ɀa<��a<��a<��a<��a<��a<o�a<m�a<w�a<{�a<��a<��a<��a<ڀa<��a<�  �  /�a<Z�a<g�a<��a<��a<ԁa<��a<�a<;�a<=�a<��a<��a<�a<)�a<_�a<Ճa<�a<��a<��a<T�a<�a<D�a<چa<I�a<Їa<:�a<��a<#�a<��a<�a<g�a<��a<K�a<��a<`�a<Ȍa<^�a<Ía<u�a<��a<��a<�a<��a<>�a<��a<N�a<��a<<�a<��a<�a<��a<�a<��a<Еa<i�a<Жa<P�a<�a<[�a<�a<��a<�a<��a<$�a<��a<-�a<��a<�a<��a<ޝa<3�a<��a<Ǟa<+�a<M�a<��a<�a<>�a<u�a<��a<�a<>�a<��a<��a<��a<&�a<L�a<�a<��a<��a<��a<��a<��a<ʢa<ߢa<Тa<�a<��a<�a<=�a<L�a<��a<��a<֣a<�a<�a<5�a<O�a<m�a<Z�a<y�a<m�a<v�a<_�a<V�a<G�a<�a<9�a<�a<%�a<�a<��a<��a<�a<�a<ƣa<��a<��a<z�a<O�a<�a<�a<��a<y�a<�a< �a<��a<��a<V�a<�a<�a<͠a<��a<��a<q�a<o�a<:�a<5�a<�a<�a<��a<o�a<8�a<�a<Şa<S�a<"�a<��a<]�a<1�a<Ȝa<��a<�a<�a<��a<E�a<�a<��a<1�a<��a<^�a<јa<_�a<̗a<?�a<��a<'�a<��a<�a<��a<	�a<��a<.�a<��a<S�a<ˑa<c�a<��a<��a<6�a<��a<a�a<ʎa<a�a<ݍa<X�a<�a<E�a<܋a<7�a<׊a<U�a<�a<n�a<��a<��a<5�a<��a<z�a<�a<��a<L�a<��a<}�a<�a<��a<?�a<ȃa<o�a<�a<��a<��a<�a<�a<��a<��a<�a<B�a<L�a<&�a<)�a<�a<�a<�a<׀a<ހa<��a<��a<��a<��a<��a<X�a<��a<p�a<��a<y�a<��a<Հa<�a<�a<�  �  5�a<`�a<��a<��a<��a<ǁa<�a<�a<.�a<D�a<l�a<��a<ׂa<�a<\�a<��a<�a<q�a<ބa<X�a<ۅa<X�a<��a<D�a<��a<E�a<��a<4�a<��a<�a<�a<��a<u�a<ߋa<c�a<ӌa<k�a<�a<��a<�a<��a<�a<��a<?�a<ȑa<9�a<��a<!�a<��a<�a<��a<�a<R�a<֕a<F�a<Öa<I�a<̗a<_�a<ߘa<}�a<�a<��a<)�a<��a<.�a<��a<$�a<��a<�a<-�a<��a<�a<5�a<y�a<��a<��a<H�a<��a<ݠa< �a<U�a<��a<áa<�a<2�a<\�a<m�a<��a<��a<��a<��a<��a<��a<��a<բa<עa<�a<��a<)�a<L�a<k�a<��a<ˣa<�a<�a<#�a<J�a<`�a<w�a<y�a<u�a<`�a<k�a<c�a<Y�a<=�a<:�a<�a<"�a<�a<�a<�a<��a<ԣa<ˣa<��a<��a<t�a<E�a<
�a<Ӣa<��a<l�a<!�a<�a<��a<w�a<5�a<�a<�a<Πa<��a<��a<v�a<g�a<M�a<�a< �a<ٟa<��a<~�a<I�a<��a<��a<l�a<)�a<ܝa<|�a<4�a<Ӝa<��a<>�a<��a<��a<F�a<ٚa<��a<2�a<ʙa<I�a<Ԙa<D�a<Ǘa<L�a<��a<&�a<��a<�a<~�a<��a<��a<�a<��a<"�a<Ǒa<`�a<�a<��a<�a<��a<J�a<�a<g�a<�a<R�a<ߌa<`�a<�a<b�a<�a<`�a<��a<��a<&�a<��a<L�a<�a<|�a<-�a<��a<\�a<�a<{�a<��a<��a<=�a<Ƀa<`�a<��a<��a<T�a<�a<ρa<��a<��a<]�a<F�a<A�a<4�a<�a<�a<�a<��a<�a<ހa<ǀa<��a<��a<��a<��a<�a<��a<z�a<��a<��a<Āa<܀a<��a<�a<�  �  ��a<��a<ۂa<�a<�a<D�a<L�a<]�a<{�a<كa<�a<9�a<g�a<��a<��a<%�a<��a<��a<c�a<نa<�a<��a<�a<��a<�a<��a<�a<d�a<��a<:�a<��a<�a<��a<�a<��a<�a<��a<&�a<��a<G�a<��a<M�a<��a<>�a<��a<P�a<�a<O�a<Ɣa<�a<��a<C�a<��a<7�a<w�a<�a<��a<�a<��a<�a<��a<�a<��a<&�a<��a<;�a<��a<&�a<]�a<�a<9�a<��a<�a<��a<i�a<��a<��a<<�a<}�a<��a<�a<l�a<x�a<ۢa<��a<�a<e�a<^�a<��a<��a<��a<��a<ۣa<�a<�a<�a<��a<9�a<5�a<V�a<��a<��a<Ҥa<��a<ޤa<�a<A�a<Z�a<X�a<{�a<S�a<��a<d�a<w�a<`�a<:�a<I�a<.�a<3�a<�a<�a<��a<��a<�a<Ѥa<��a<��a<��a<q�a<S�a</�a<�a<��a<c�a<a�a<�a<��a<��a<l�a<`�a<�a<�a<�a<��a<��a<L�a<D�a<)�a<#�a<ՠa<��a<q�a<3�a<�a<��a<��a<��a<��a<{�a<0�a<��a<�a<B�a<Ȝa<��a<D�a<�a<��a<�a<ۚa<A�a<�a<Z�a<ۘa<6�a<��a<o�a<Öa<m�a<��a<H�a<Ҕa<:�a<�a<h�a<�a<��a<�a<��a<J�a<��a<d�a<�a<s�a<'�a<��a<�a<��a<�a<��a<�a<��a<5�a<Êa<P�a<Ӊa<��a<�a<�a<k�a<��a<��a<+�a<�a<[�a<�a<t�a<D�a<�a<��a<R�a<̓a<��a<_�a<2�a<$�a<�a<߂a<��a<{�a<��a<��a<s�a<O�a<U�a<�a<H�a<�a<�a<��a<Ӂa<�a<ځa<��a<�a<�a<�a<)�a<e�a<`�a<�  �  ��a<��a<Ђa<�a<�a<'�a<Z�a<��a<��a<a<��a<�a<T�a<��a<�a<9�a<��a<�a<L�a<Ɇa<Y�a<ȇa<!�a<��a<�a<w�a<�a<i�a<Ίa<7�a<��a<1�a<��a<!�a<��a<�a<��a<4�a<��a<+�a<��a<:�a<Αa<Q�a<ْa<U�a<ۓa<E�a<ݔa<[�a<��a<!�a<��a<�a<��a<�a<��a<��a<��a< �a<��a<0�a<̛a<F�a<��a<+�a<��a<�a<l�a<͞a<�a<x�a<ȟa<%�a<~�a<��a<�a<=�a<��a<ڡa<�a<A�a<r�a<��a<�a<�a<?�a<e�a<��a<��a<Σa<�a<ԣa<ѣa<�a<�a<
�a<(�a<?�a<P�a<d�a<��a<��a<��a<�a<(�a<'�a<N�a<N�a<e�a<i�a<f�a<[�a<b�a<T�a<^�a<N�a<>�a<+�a<$�a<�a<�a<��a<�a<Ȥa<��a<��a<��a<c�a<N�a<�a<��a<ԣa<��a<J�a<�a<΢a<��a<z�a<N�a<!�a<�a<ˡa<��a<��a<��a<q�a<0�a<�a<٠a<��a<q�a<8�a<�a<��a<`�a<�a<ߞa<��a<2�a<ٝa<��a<P�a<��a<��a<=�a<ٛa<��a<�a<��a<F�a<ڙa<P�a<�a<x�a<�a<M�a<��a<8�a<��a<F�a<̔a<J�a<֓a<\�a<��a<��a<M�a<ّa<J�a<�a<n�a<��a<��a<�a<}�a<�a<��a<�a<��a< �a<��a<6�a<̊a<q�a<��a<��a<�a<��a<e�a<��a<��a<1�a<φa<c�a<�a<��a<=�a<τa<w�a<&�a<��a<��a<j�a<,�a<��a<ւa<Ȃa<ǂa<��a<��a<f�a<g�a<E�a<?�a<+�a<�a<��a<��a<�a<��a<�a<�a<�a<��a<�a<*�a<*�a<I�a<X�a<�  �  v�a<Ăa<ɂa<�a<�a<+�a<e�a<[�a<��a<��a<�a<+�a<g�a<��a<Ԅa<\�a<��a<�a<w�a<��a<9�a<��a<3�a<��a<�a<n�a<��a<u�a<Ŋa<f�a<��a<,�a<��a<��a<��a<�a<��a<��a<��a<�a<Аa<P�a<đa<l�a<��a<g�a<ѓa<[�a<ʔa<.�a<��a<�a<��a<�a<��a<�a<��a<*�a<��a<:�a<��a<�a<��a<)�a<��a<�a<��a<�a<��a<ɞa<(�a<��a<��a<!�a<=�a<��a<�a<:�a<j�a<��a<	�a<&�a<��a<��a<��a<)�a<2�a<z�a<z�a<��a<��a<��a<��a<�a<�a<�a</�a<�a<O�a<q�a<w�a<��a<��a<٤a<�a<'�a<1�a<L�a<[�a<Y�a<��a<[�a<~�a<a�a<>�a<Q�a< �a<:�a<�a<"�a<��a<�a<�a<�a<�a<��a<Ƥa<��a<h�a<P�a<�a<��a<��a<��a<>�a<:�a<�a<��a<��a<8�a<D�a<�a<�a<ԡa<��a<x�a<=�a<B�a<��a<�a<��a<x�a<D�a<�a<ʟa<L�a<�a<��a<_�a<*�a<ӝa<��a<�a<�a<w�a<S�a<�a<|�a<9�a<��a<X�a<Йa<e�a<ߘa<L�a<Ηa<E�a<�a<>�a<�a<H�a<ǔa<v�a<ԓa<��a<�a<��a<"�a<��a<c�a<ܐa<��a<�a<��a<�a<��a<&�a<o�a<�a<m�a<�a<��a<3�a<��a<9�a<��a<m�a<E�a<��a<m�a<�a<��a<F�a<a<w�a<�a<��a<&�a<�a<��a<&�a<�a<��a<z�a<M�a<	�a<�a<��a<��a<}�a<��a<q�a<d�a<R�a<3�a<K�a<
�a<!�a<��a<Ձa<�a<��a<�a<ہa<��a<�a<�a<�a<B�a<��a<�  �  y�a<��a<ła<��a<�a<A�a<h�a<y�a<��a<Ӄa< �a<$�a<l�a<��a<��a<K�a<��a<�a<e�a<܆a<[�a<��a<@�a<��a<�a<��a<�a<Z�a<Ŋa<9�a<��a<'�a<��a<*�a<}�a<�a<��a<�a<��a<$�a<��a<*�a<Ña<N�a<֒a<k�a<ʓa<n�a<єa<R�a<וa<,�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<I�a<ƛa<5�a<̜a<�a<��a<�a<e�a<Ğa<�a<n�a<��a<�a<T�a<��a<ՠa<�a<��a<��a<�a<6�a<t�a<��a<�a<�a<K�a<s�a<~�a<��a<��a<�a<�a<�a<�a<
�a<�a<8�a<I�a<g�a<}�a<��a<¤a< �a<�a<)�a<K�a<C�a<g�a<]�a<^�a<[�a<V�a<X�a<K�a<I�a<C�a<+�a<��a<�a<�a<��a<�a<�a<̤a<��a<��a<��a<w�a<D�a<,�a<�a<��a<��a<[�a<$�a<ߢa<��a<��a<^�a<4�a<�a<֡a<��a<��a<��a<V�a<O�a<�a<�a<��a<g�a<(�a<��a<��a<V�a<�a<��a<��a<�a<��a<��a<-�a<�a<��a<2�a<ɛa<z�a<�a<��a<\�a<șa<y�a<�a<p�a<��a<X�a<Жa<L�a<ѕa<Q�a<ڔa<b�a<�a<v�a<�a<��a<G�a<Ǒa<r�a<אa<��a<��a<{�a<��a<o�a<��a<��a<�a<��a<"�a<��a<�a<Պa<J�a<�a<}�a<�a<��a<W�a<�a<��a<?�a<Ɔa<��a<�a<��a<R�a<�a<��a<>�a<��a<��a<t�a<C�a<�a<�a<ςa<ӂa<��a<��a<��a<[�a<^�a<7�a< �a<�a<��a<�a<�a<�a<�a<ׁa<��a<�a<�a<�a<!�a<C�a<\�a<�  �  ��a<��a<ςa<�a<�a<D�a<A�a<��a<��a<ڃa<
�a<Q�a<��a<��a<!�a<<�a<Ӆa<�a<v�a<׆a<Z�a<��a<�a<��a<�a<�a<�a<a�a<ۊa<"�a<��a<�a<{�a<�a<n�a< �a<n�a<�a<u�a<#�a<��a<0�a<ڑa<G�a<ݒa<X�a<��a<[�a<��a<]�a<��a<D�a<��a<M�a<��a</�a<��a<�a<ϙa<'�a<��a<-�a<̛a<+�a<��a<3�a<��a<	�a<a�a<؞a<�a<h�a<��a<�a<S�a<��a<֠a<�a<^�a<��a<ޡa<>�a<a�a<��a<�a<�a<D�a<f�a<��a<��a<��a<�a<ޣa<��a<�a<A�a<�a<^�a<R�a<~�a<��a<��a<Ӥa<�a<�a<�a<E�a<M�a<V�a<g�a<X�a<s�a<J�a<\�a<B�a<�a<.�a<
�a<�a<�a<��a<Ӥa<ݤa<�a<��a<̤a<��a<��a<l�a<J�a</�a<ۣa<֣a<��a<b�a<.�a<�a<ڢa<��a<��a<%�a<;�a<��a<ҡa<��a<��a<h�a<*�a<�a<ڠa<��a<k�a</�a<��a<��a<]�a<�a<��a<a�a<�a<ŝa<`�a<)�a<��a<��a<-�a<Λa<��a<�a<��a<H�a<ߙa<f�a<Ҙa<{�a<ߗa<p�a<ݖa<��a<֕a<o�a<��a<_�a<"�a<��a<"�a<��a<M�a<��a<Z�a<�a<r�a<��a<w�a<�a<|�a<��a<��a<ߌa<��a<�a<��a<�a<��a<9�a<ˉa<��a<�a<a<d�a<��a<��a<2�a<݆a<f�a<�a<��a<G�a<��a<��a<v�a<�a<܃a<|�a<Z�a<=�a<��a<��a<Ăa<��a<r�a<��a<f�a<L�a<B�a<�a<#�a<�a<��a<فa<��a<΁a<��a<؁a<ǁa<�a<�a<�a<G�a<H�a<�  �  h�a<��a<͂a<�a<�a<E�a<g�a<��a<��a<�a<+�a<=�a<��a<Ȅa<#�a<e�a<ȅa<�a<��a<�a<O�a<a<5�a<��a<�a<�a<�a<E�a<��a<(�a<��a<�a<��a<ٌa<k�a<��a<L�a<��a<��a<�a<��a<$�a<��a<K�a<֒a<]�a<�a<^�a<ܔa<c�a<��a<f�a<a<8�a<��a<6�a<��a<1�a<��a<8�a<�a<*�a<қa<A�a<��a<6�a<��a<�a<i�a<��a<�a<[�a<��a<��a<H�a<]�a<۠a<�a<5�a<��a<�a< �a<c�a<��a<̢a<�a<B�a<k�a<��a<��a<ģa<ߣa<�a<'�a<�a<1�a<:�a<Y�a<f�a<��a<��a<ˤa<�a<�a<�a<,�a<C�a<V�a<Z�a<e�a<Y�a<J�a<M�a<;�a<9�a</�a<�a<�a<�a<�a<�a<�a<ݤa<��a<��a<��a<��a<��a<p�a<R�a<1�a<�a<գa<��a<u�a<N�a<��a<�a<��a<��a<M�a<1�a<�a< �a<��a<��a<k�a<D�a<�a<ߠa<��a<q�a<�a<͟a<��a<>�a<��a<��a<9�a<��a<ĝa<>�a<�a<ǜa<t�a<�a<Ûa<a�a<�a<��a<N�a<�a<i�a<�a<��a<ԗa<��a<�a<n�a<�a<v�a<��a<}�a<�a<��a<J�a<��a<S�a<ԑa<b�a<�a<v�a<��a<�a<�a<g�a<�a<k�a<�a<x�a<̋a<��a<�a<{�a<:�a<͉a<g�a<	�a<��a<@�a< �a<��a<7�a<߆a<y�a<�a<��a<N�a<$�a<��a<e�a<�a<׃a<��a<k�a<(�a<�a<��a<��a<��a<��a<��a<n�a<Q�a<?�a<�a<��a<��a<Ձa<Ёa<ǁa<��a<��a<сa<��a<ҁa<��a<�a< �a<N�a<�  �  g�a<��a<��a<�a<�a<:�a<y�a<��a<߃a<�a<)�a<V�a<��a<�a<"�a<��a<܅a<#�a<��a<�a<}�a<ʇa<F�a<��a<�a<x�a<݉a<R�a<��a<+�a<�a<�a<e�a<�a<L�a<ƍa<a�a<�a<c�a<��a<��a<6�a<��a<N�a<Òa<b�a<ړa<e�a<�a<s�a<�a<X�a<ϖa<R�a<ԗa<@�a<��a<Q�a<әa<K�a<Қa<U�a<�a<H�a<Ȝa<(�a<��a<��a<c�a<��a<�a<N�a<��a<ٟa<-�a<s�a<��a<�a<F�a<��a<ơa<�a<^�a<��a<Ңa<�a<9�a<s�a<��a<ãa<ͣa<�a<��a<�a<�a<C�a<]�a<\�a<{�a<��a<��a<Фa<�a<�a<&�a<>�a<>�a<M�a<Y�a<N�a<a�a<I�a<[�a<'�a<!�a<�a<�a<��a<ܤa<ݤa<ݤa<��a<¤a<��a<ˤa<��a<��a<z�a<j�a<L�a<%�a<�a<ۣa<ǣa<p�a<M�a<�a<��a<��a<��a<m�a<E�a<�a<�a<��a<��a<s�a<U�a<�a<�a<��a<[�a<!�a<ٟa<��a<(�a<ܞa<��a<D�a<��a<��a<T�a<�a<��a<b�a<�a<ԛa<b�a<�a<��a<S�a<ٙa<p�a<��a<��a<
�a<��a< �a<��a<�a<��a<�a<��a<'�a<��a<9�a<Ȓa<i�a<ۑa<o�a<�a<~�a<�a<y�a<�a<{�a<ލa<[�a<Ќa<]�a<�a<U�a<�a<��a<�a<��a<U�a<�a<��a<F�a<�a<��a<?�a<φa<��a<�a<݅a<c�a<�a<��a<w�a<4�a<ۃa<��a<��a<E�a<�a<�a<�a<Âa<��a<~�a<f�a<P�a<(�a<$�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<́a<́a<��a<�a<[�a<�  �  a�a<��a<Ƃa<�a<�a<P�a<n�a<��a<Ӄa<��a<D�a<��a<��a<�a<Z�a<x�a<�a<M�a<��a<�a<m�a<ʇa<?�a<��a<�a<�a<މa<C�a<��a<��a<��a<�a<I�a<όa<:�a<��a<>�a<юa<J�a<�a<n�a<�a<��a<:�a<Ӓa<Z�a<�a<x�a<ߔa<a�a<�a<j�a<�a<n�a<��a<l�a<�a<=�a<�a<g�a<�a<a�a<қa<D�a<Ӝa<6�a<��a<�a<S�a<��a< �a<)�a<��a<ğa<�a<R�a<��a<�a<,�a<k�a<��a<�a<%�a<��a<ʢa<�a<C�a<m�a<��a<��a<̣a<�a<�a<,�a<D�a<Y�a<J�a<��a<��a<��a<Ԥa<�a<��a<�a<�a</�a<T�a<S�a<X�a<^�a<P�a<C�a<,�a<�a<0�a<�a<��a<ڤa<ߤa<��a<Ǥa<��a<Ȥa<��a<��a<��a<��a<��a<n�a<R�a<;�a<�a<٣a<��a<��a<h�a<;�a<��a<Ƣa<��a<a�a<U�a<2�a<�a<ҡa<��a<s�a<N�a<"�a<�a<��a<[�a<�a<Οa<[�a<3�a<՞a<o�a<.�a<ϝa<��a<1�a<�a<��a<q�a<�a<��a<Z�a<�a<��a<K�a<�a<��a<��a<�a<�a<��a<�a<��a<��a<��a<7�a<��a<C�a<Óa<K�a<Ԓa<T�a<בa<y�a<�a<u�a<��a<i�a<ߎa<c�a<��a<j�a<��a<E�a<��a<M�a<܊a<r�a<�a<��a<b�a<̈a<��a<>�a<�a<��a<9�a<�a<��a<�a<˅a<t�a<)�a<ڄa<��a< �a<�a<��a<y�a<f�a<7�a<�a<�a<��a<��a<��a<l�a<O�a<8�a<�a<�a<ρa<��a<ǁa<��a<��a<��a<��a<��a<��a<��a<��a<�a<+�a<�  �  c�a<l�a<a<�a<�a<O�a<z�a<��a<ʃa<"�a<B�a<m�a<Ʉa<��a<`�a<��a<��a<8�a<��a<!�a<k�a<�a<<�a<��a<�a<x�a<��a<�a<��a<�a<o�a<ыa<]�a<��a<,�a<Ǎa<�a<�a<C�a<��a<h�a<�a<��a<,�a<Ӓa<U�a<�a<k�a<�a<��a<�a<��a<�a<p�a<�a<g�a<�a<b�a<��a<\�a<��a<k�a<�a<q�a<ɜa<<�a<��a<�a<I�a<��a<��a<(�a<��a<��a<(�a<1�a<��a<٠a<�a<��a<��a<��a<3�a<��a<��a<�a<<�a<h�a<��a<��a<��a<��a<"�a<=�a<2�a<j�a<j�a<��a<��a<��a<Ǥa<�a<�a<
�a<G�a<G�a<Q�a<T�a<R�a<Y�a<2�a<A�a<6�a<�a<�a<��a<��a<��a<ܤa<��a<Ĥa<��a<��a<��a<��a<��a<n�a<��a<h�a<P�a<:�a<�a<�a<��a<��a<e�a<'�a<�a<բa<Ģa<|�a<h�a<�a<�a<�a<��a<��a<K�a<$�a<ݠa<��a<]�a<�a<͟a<i�a<�a<��a<��a<�a<��a<��a<
�a< �a<��a<D�a<�a<��a<R�a<��a<��a<F�a<�a<v�a<�a<��a<�a<��a<�a<��a<#�a<��a<1�a<��a<K�a<��a<c�a<ޒa<m�a<�a<o�a<��a<q�a<��a<_�a<͎a<_�a<��a<A�a<��a<Y�a<��a<S�a<Ҋa<X�a<�a<��a<B�a<ڈa<��a<�a<�a<��a<4�a<�a<��a<J�a<Ӆa<��a<:�a<Ȅa<��a<@�a<�a<Ńa<��a<Y�a<4�a<&�a<܂a<�a<��a<��a<m�a<I�a<3�a<�a<�a<؁a<��a<��a<��a<��a<a�a<��a<v�a<��a<ǁa<ځa<��a<1�a<�  �  I�a<��a<��a<�a< �a<G�a<w�a<��a<�a<�a<S�a<��a<�a<�a<D�a<��a<�a<g�a<��a<�a<t�a<އa<C�a<��a<"�a<k�a<�a<?�a<��a<�a<[�a<ǋa<.�a<��a<�a<��a<"�a<��a<1�a<Ϗa<w�a<�a<��a<J�a<��a<c�a<�a<j�a<��a<p�a<��a<}�a<
�a<}�a<�a<p�a<�a<��a<��a<��a<��a<u�a<ޛa<`�a<˜a<<�a<��a<�a<d�a<��a<��a<A�a<k�a<��a<�a<8�a<}�a<��a<	�a<L�a<��a<�a<O�a<��a<��a<�a<)�a<~�a<��a<��a<�a<��a<&�a<@�a<_�a<r�a<��a<��a<��a<�a<�a< �a<�a<"�a</�a<B�a<K�a<Z�a<W�a<K�a<X�a<,�a<9�a<�a<��a<Ҥa<Τa<Ťa<��a<��a<��a<��a<��a<��a<��a<��a<��a<�a<c�a<X�a<2�a<�a<�a<ʣa<��a<v�a<N�a<5�a<�a<��a<��a<y�a<L�a<�a<�a<��a<��a<R�a<�a<�a<��a<j�a<�a<��a<|�a<�a<��a<T�a<�a<��a<g�a<�a<ɜa<r�a<3�a<��a<��a<L�a<�a<��a<S�a<�a<u�a<�a<��a<$�a<��a<;�a<��a<W�a<��a<4�a<�a<O�a<�a<_�a<�a<_�a<�a<r�a<��a<�a<ۏa<z�a<юa<Y�a<эa<,�a<��a< �a<��a</�a<��a<N�a<�a<��a<+�a<��a<��a<5�a<��a<}�a<J�a<�a<��a<2�a<҅a<��a<=�a<��a<��a<l�a<�a<փa<ăa<y�a<N�a< �a<��a<̂a<��a<��a<s�a<N�a<%�a<�a<ہa<܁a<��a<��a<k�a<m�a<q�a<r�a<��a<��a<��a<΁a<��a<6�a<�  �  -�a<��a<��a<�a<�a<O�a<��a<��a<
�a<�a<O�a<��a<a<(�a<c�a<Åa<��a<r�a<��a<+�a<��a<݇a<l�a<��a<�a<q�a<щa<;�a<v�a<�a<G�a<�a<%�a<��a< �a<��a<2�a<��a<T�a<ҏa<J�a<�a<��a<:�a<��a<i�a<֓a<��a<	�a<|�a<)�a<m�a<�a<i�a<��a<��a<�a<��a<�a<��a<�a<��a<�a<i�a<�a<$�a<��a<�a<U�a<��a<ўa<�a<d�a<ɟa<ٟa<H�a<f�a<��a<�a<A�a<��a<Сa<!�a<]�a<��a<��a</�a<w�a<��a<�a<�a<�a<A�a<.�a<l�a<V�a<��a<��a<��a<��a<�a<�a<	�a<O�a<.�a<_�a<W�a<E�a<`�a<?�a<N�a<�a<�a<�a<
�a<�a<��a<Ѥa<��a<��a<��a<��a<��a<{�a<��a<i�a<��a<l�a<o�a<I�a<:�a<4�a<�a<�a<��a<s�a<S�a<�a<�a<Ǣa<��a<Y�a<W�a<�a<��a<ۡa<��a<{�a<�a<�a<��a<O�a<
�a<��a<S�a<�a<Оa<K�a<�a<��a<G�a<$�a<��a<��a<6�a<͛a<��a<8�a<�a<��a<Z�a<ՙa<��a<�a<��a<N�a<��a<C�a<��a<6�a<͕a<R�a<͔a<9�a<�a<N�a<�a<t�a<��a<��a<�a<��a<ޏa<k�a<Ďa<4�a<��a<%�a<��a<	�a<��a<�a<��a<c�a<؉a<��a<�a<Ȉa<h�a<0�a<އa<��a<C�a<φa<��a<3�a<��a<��a<+�a<�a<��a<k�a< �a<�a<��a<u�a<P�a<�a<"�a<˂a<˂a<��a<^�a<W�a<�a<�a<��a<��a<��a<��a<��a<[�a<}�a<J�a<��a<��a<��a<�a<ہa<�a<�  �  d�a<��a<��a<�a<�a<R�a<��a<��a<݃a<#�a<]�a<��a<�a<+�a<o�a<ƅa<"�a<|�a<Æa<)�a<~�a<�a<M�a<��a<�a<w�a<ĉa<B�a<��a<	�a<U�a<��a<�a<��a<�a<��a<�a<��a<"�a<��a<b�a<�a<��a<&�a<Œa<S�a<�a<v�a<�a<{�a< �a<��a<�a<��a<�a<��a<
�a<��a<&�a<��a<�a<z�a<�a<j�a<Ӝa<8�a<��a<��a<=�a<��a<��a<)�a<Z�a<��a<ܟa<�a<p�a<��a<��a<7�a<��a<ۡa<9�a<��a<ʢa<�a<8�a<f�a<��a<ƣa<�a<�a<0�a<F�a<s�a<��a<��a<��a<ʤa<�a<�a<
�a<�a<�a<8�a<P�a<U�a<K�a<Q�a<F�a<=�a<F�a<5�a<�a<ۤa<Ǥa<��a<��a<��a<��a<��a<�a<y�a<��a<��a<��a<��a<k�a<h�a<G�a<>�a<�a<��a<ģa<��a<��a<m�a<4�a<�a<Ӣa<��a<��a<a�a< �a<��a<��a<��a<\�a<#�a<֠a<��a<B�a<�a<şa<m�a<��a<��a<;�a<�a<��a<Y�a<��a<��a<c�a<�a<�a<��a<e�a<�a<��a<D�a<�a<��a<�a<��a<%�a<��a<I�a<ۖa<P�a<͕a<O�a<ޔa<z�a<�a<i�a<�a<j�a<��a<z�a<��a<m�a<�a<S�a<�a<_�a<��a<�a<��a<�a<��a<"�a<��a<:�a<Ήa<m�a<"�a<��a<��a<?�a<̇a<��a<2�a<�a<��a<>�a<�a<��a<C�a<	�a<Ąa<p�a<(�a<��a<��a<��a<X�a<(�a<�a<Ղa<��a<��a<d�a<H�a<!�a< �a<��a<؁a<��a<r�a<_�a<T�a<\�a<b�a<l�a<w�a<��a<��a<�a<4�a<�  �  1�a<r�a<ǂa<�a<!�a<Z�a<r�a<�a<�a<D�a<U�a<��a<�a<#�a<x�a<��a<�a<T�a<ӆa<;�a<��a<�a<8�a<͈a<�a<��a<݉a<0�a<o�a<؊a<n�a<��a<D�a<��a<�a<��a<��a<Ďa<+�a<ӏa<c�a<ΐa<�a<�a<ܒa<M�a<	�a<n�a<�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<�a<g�a<+�a<��a<�a<��a<Ɯa<Y�a<��a<	�a<9�a<��a<��a<�a<{�a<��a<�a<�a<x�a<��a<�a<j�a<��a<��a<�a<K�a<��a<��a<D�a<e�a<��a<��a<�a<�a<;�a<_�a<H�a<��a<��a<��a<Ǥa<ޤa<�a<��a<C�a<$�a<h�a<E�a<W�a<g�a<M�a<d�a<3�a<�a<�a<�a<�a<ߤa<٤a<��a<��a<��a<��a<��a<��a<��a<b�a<l�a<t�a<��a<k�a<Y�a<E�a<�a<+�a<̣a<̣a<y�a<K�a<1�a<��a<ۢa<��a<��a<9�a</�a<�a<ơa<��a<G�a<>�a<ޠa<��a<Z�a<��a<��a<=�a<�a<��a<k�a<�a<��a<g�a<�a<��a<m�a<7�a<�a<m�a<7�a<�a<��a<=�a<�a<y�a<%�a<Ęa<-�a<ߗa<�a<��a<F�a<̕a<R�a<єa<`�a<Óa<��a<��a<��a<�a<m�a<�a<d�a<��a<N�a<��a<�a<��a<<�a<��a<C�a<}�a<)�a<��a<3�a<�a<v�a<A�a<��a<V�a<*�a<݇a<��a<1�a<�a<y�a<g�a<��a<��a<\�a<ބa<��a<`�a</�a<�a<��a<w�a<B�a<P�a<��a<�a<��a<��a<��a<D�a<?�a<��a<ǁa<��a<��a<��a<x�a<y�a<K�a<v�a<\�a<��a<��a<��a<��a<�a<�  �  d�a<��a<��a<�a<�a<R�a<��a<��a<݃a<#�a<]�a<��a<�a<+�a<o�a<ƅa<"�a<|�a<Æa<)�a<~�a<�a<M�a<��a<�a<w�a<ĉa<B�a<��a<	�a<U�a<��a<�a<��a<�a<��a<�a<��a<"�a<��a<b�a<�a<��a<&�a<Œa<S�a<�a<v�a<�a<{�a< �a<��a<�a<��a<�a<��a<
�a<��a<&�a<��a<�a<z�a<�a<j�a<Ӝa<8�a<��a<��a<=�a<��a<��a<)�a<Z�a<��a<ܟa<�a<p�a<��a<��a<7�a<��a<ۡa<9�a<��a<ʢa<�a<8�a<f�a<��a<ƣa<�a<�a<0�a<F�a<s�a<��a<��a<��a<ʤa<�a<�a<
�a<�a<�a<8�a<P�a<U�a<K�a<Q�a<F�a<=�a<F�a<5�a<�a<ۤa<Ǥa<��a<��a<��a<��a<��a<�a<y�a<��a<��a<��a<��a<k�a<h�a<G�a<>�a<�a<��a<ģa<��a<��a<m�a<4�a<�a<Ӣa<��a<��a<a�a< �a<��a<��a<��a<\�a<#�a<֠a<��a<B�a<�a<şa<m�a<��a<��a<;�a<�a<��a<Y�a<��a<��a<c�a<�a<�a<��a<e�a<�a<��a<D�a<�a<��a<�a<��a<%�a<��a<I�a<ۖa<P�a<͕a<O�a<ޔa<z�a<�a<i�a<�a<j�a<��a<z�a<��a<m�a<�a<S�a<�a<_�a<��a<�a<��a<�a<��a<"�a<��a<:�a<Ήa<m�a<"�a<��a<��a<?�a<̇a<��a<2�a<�a<��a<>�a<�a<��a<C�a<	�a<Ąa<p�a<(�a<��a<��a<��a<X�a<(�a<�a<Ղa<��a<��a<d�a<H�a<!�a< �a<��a<؁a<��a<r�a<_�a<T�a<\�a<b�a<l�a<w�a<��a<��a<�a<4�a<�  �  -�a<��a<��a<�a<�a<O�a<��a<��a<
�a<�a<O�a<��a<a<(�a<c�a<Åa<��a<r�a<��a<+�a<��a<݇a<l�a<��a<�a<q�a<щa<;�a<v�a<�a<G�a<�a<%�a<��a< �a<��a<2�a<��a<T�a<ҏa<J�a<�a<��a<:�a<��a<i�a<֓a<��a<	�a<|�a<)�a<m�a<�a<i�a<��a<��a<�a<��a<�a<��a<�a<��a<�a<i�a<�a<$�a<��a<�a<U�a<��a<ўa<�a<d�a<ɟa<ٟa<H�a<f�a<��a<�a<A�a<��a<Сa<!�a<]�a<��a<��a</�a<w�a<��a<�a<�a<�a<A�a<.�a<l�a<V�a<��a<��a<��a<��a<�a<�a<	�a<O�a<.�a<_�a<W�a<E�a<`�a<?�a<N�a<�a<�a<�a<
�a<�a<��a<Ѥa<��a<��a<��a<��a<��a<{�a<��a<i�a<��a<l�a<o�a<I�a<:�a<4�a<�a<�a<��a<s�a<S�a<�a<�a<Ǣa<��a<Y�a<W�a<�a<��a<ۡa<��a<{�a<�a<�a<��a<O�a<
�a<��a<S�a<�a<Оa<K�a<�a<��a<G�a<$�a<��a<��a<6�a<͛a<��a<8�a<�a<��a<Z�a<ՙa<��a<�a<��a<N�a<��a<C�a<��a<6�a<͕a<R�a<͔a<9�a<�a<N�a<�a<t�a<��a<��a<�a<��a<ޏa<k�a<Ďa<4�a<��a<%�a<��a<	�a<��a<�a<��a<c�a<؉a<��a<�a<Ȉa<h�a<0�a<އa<��a<C�a<φa<��a<3�a<��a<��a<+�a<�a<��a<k�a< �a<�a<��a<u�a<P�a<�a<"�a<˂a<˂a<��a<^�a<W�a<�a<�a<��a<��a<��a<��a<��a<[�a<}�a<J�a<��a<��a<��a<�a<ہa<�a<�  �  I�a<��a<��a<�a< �a<G�a<w�a<��a<�a<�a<S�a<��a<�a<�a<D�a<��a<�a<g�a<��a<�a<t�a<އa<C�a<��a<"�a<k�a<�a<?�a<��a<�a<[�a<ǋa<.�a<��a<�a<��a<"�a<��a<1�a<Ϗa<w�a<�a<��a<J�a<��a<c�a<�a<j�a<��a<p�a<��a<}�a<
�a<}�a<�a<p�a<�a<��a<��a<��a<��a<u�a<ޛa<`�a<˜a<<�a<��a<�a<d�a<��a<��a<A�a<k�a<��a<�a<8�a<}�a<��a<	�a<L�a<��a<�a<O�a<��a<��a<�a<)�a<~�a<��a<��a<�a<��a<&�a<@�a<_�a<r�a<��a<��a<��a<�a<�a< �a<�a<"�a</�a<B�a<K�a<Z�a<W�a<K�a<X�a<,�a<9�a<�a<��a<Ҥa<Τa<Ťa<��a<��a<��a<��a<��a<��a<��a<��a<��a<�a<c�a<X�a<2�a<�a<�a<ʣa<��a<v�a<N�a<5�a<�a<��a<��a<y�a<L�a<�a<�a<��a<��a<R�a<�a<�a<��a<j�a<�a<��a<|�a<�a<��a<T�a<�a<��a<g�a<�a<ɜa<r�a<3�a<��a<��a<L�a<�a<��a<S�a<�a<u�a<�a<��a<$�a<��a<;�a<��a<W�a<��a<4�a<�a<O�a<�a<_�a<�a<_�a<�a<r�a<��a<�a<ۏa<z�a<юa<Y�a<эa<,�a<��a< �a<��a</�a<��a<N�a<�a<��a<+�a<��a<��a<5�a<��a<}�a<J�a<�a<��a<2�a<҅a<��a<=�a<��a<��a<l�a<�a<փa<ăa<y�a<N�a< �a<��a<̂a<��a<��a<s�a<N�a<%�a<�a<ہa<܁a<��a<��a<k�a<m�a<q�a<r�a<��a<��a<��a<΁a<��a<6�a<�  �  c�a<l�a<a<�a<�a<O�a<z�a<��a<ʃa<"�a<B�a<m�a<Ʉa<��a<`�a<��a<��a<8�a<��a<!�a<k�a<�a<<�a<��a<�a<x�a<��a<�a<��a<�a<o�a<ыa<]�a<��a<,�a<Ǎa<�a<�a<C�a<��a<h�a<�a<��a<,�a<Ӓa<U�a<�a<k�a<�a<��a<�a<��a<�a<p�a<�a<g�a<�a<b�a<��a<\�a<��a<k�a<�a<q�a<ɜa<<�a<��a<�a<I�a<��a<��a<(�a<��a<��a<(�a<1�a<��a<٠a<�a<��a<��a<��a<3�a<��a<��a<�a<<�a<h�a<��a<��a<��a<��a<"�a<=�a<2�a<j�a<j�a<��a<��a<��a<Ǥa<�a<�a<
�a<G�a<G�a<Q�a<T�a<R�a<Y�a<2�a<A�a<6�a<�a<�a<��a<��a<��a<ܤa<��a<Ĥa<��a<��a<��a<��a<��a<n�a<��a<h�a<P�a<:�a<�a<�a<��a<��a<e�a<'�a<�a<բa<Ģa<|�a<h�a<�a<�a<�a<��a<��a<K�a<$�a<ݠa<��a<]�a<�a<͟a<i�a<�a<��a<��a<�a<��a<��a<
�a< �a<��a<D�a<�a<��a<R�a<��a<��a<F�a<�a<v�a<�a<��a<�a<��a<�a<��a<#�a<��a<1�a<��a<K�a<��a<c�a<ޒa<m�a<�a<o�a<��a<q�a<��a<_�a<͎a<_�a<��a<A�a<��a<Y�a<��a<S�a<Ҋa<X�a<�a<��a<B�a<ڈa<��a<�a<�a<��a<4�a<�a<��a<J�a<Ӆa<��a<:�a<Ȅa<��a<@�a<�a<Ńa<��a<Y�a<4�a<&�a<܂a<�a<��a<��a<m�a<I�a<3�a<�a<�a<؁a<��a<��a<��a<��a<a�a<��a<v�a<��a<ǁa<ځa<��a<1�a<�  �  a�a<��a<Ƃa<�a<�a<P�a<n�a<��a<Ӄa<��a<D�a<��a<��a<�a<Z�a<x�a<�a<M�a<��a<�a<m�a<ʇa<?�a<��a<�a<�a<މa<C�a<��a<��a<��a<�a<I�a<όa<:�a<��a<>�a<юa<J�a<�a<n�a<�a<��a<:�a<Ӓa<Z�a<�a<x�a<ߔa<a�a<�a<j�a<�a<n�a<��a<l�a<�a<=�a<�a<g�a<�a<a�a<қa<D�a<Ӝa<6�a<��a<�a<S�a<��a< �a<)�a<��a<ğa<�a<R�a<��a<�a<,�a<k�a<��a<�a<%�a<��a<ʢa<�a<C�a<m�a<��a<��a<̣a<�a<�a<,�a<D�a<Y�a<J�a<��a<��a<��a<Ԥa<�a<��a<�a<�a</�a<T�a<S�a<X�a<^�a<P�a<C�a<,�a<�a<0�a<�a<��a<ڤa<ߤa<��a<Ǥa<��a<Ȥa<��a<��a<��a<��a<��a<n�a<R�a<;�a<�a<٣a<��a<��a<h�a<;�a<��a<Ƣa<��a<a�a<U�a<2�a<�a<ҡa<��a<s�a<N�a<"�a<�a<��a<[�a<�a<Οa<[�a<3�a<՞a<o�a<.�a<ϝa<��a<1�a<�a<��a<q�a<�a<��a<Z�a<�a<��a<K�a<�a<��a<��a<�a<�a<��a<�a<��a<��a<��a<7�a<��a<C�a<Óa<K�a<Ԓa<T�a<בa<y�a<�a<u�a<��a<i�a<ߎa<c�a<��a<j�a<��a<E�a<��a<M�a<܊a<r�a<�a<��a<b�a<̈a<��a<>�a<�a<��a<9�a<�a<��a<�a<˅a<t�a<)�a<ڄa<��a< �a<�a<��a<y�a<f�a<7�a<�a<�a<��a<��a<��a<l�a<O�a<8�a<�a<�a<ρa<��a<ǁa<��a<��a<��a<��a<��a<��a<��a<��a<�a<+�a<�  �  g�a<��a<��a<�a<�a<:�a<y�a<��a<߃a<�a<)�a<V�a<��a<�a<"�a<��a<܅a<#�a<��a<�a<}�a<ʇa<F�a<��a<�a<x�a<݉a<R�a<��a<+�a<�a<�a<e�a<�a<L�a<ƍa<a�a<�a<c�a<��a<��a<6�a<��a<N�a<Òa<b�a<ړa<e�a<�a<s�a<�a<X�a<ϖa<R�a<ԗa<@�a<��a<Q�a<әa<K�a<Қa<U�a<�a<H�a<Ȝa<(�a<��a<��a<c�a<��a<�a<N�a<��a<ٟa<-�a<s�a<��a<�a<F�a<��a<ơa<�a<^�a<��a<Ңa<�a<9�a<s�a<��a<ãa<ͣa<�a<��a<�a<�a<C�a<]�a<\�a<{�a<��a<��a<Фa<�a<�a<&�a<>�a<>�a<M�a<Y�a<N�a<a�a<I�a<[�a<'�a<!�a<�a<�a<��a<ܤa<ݤa<ݤa<��a<¤a<��a<ˤa<��a<��a<z�a<j�a<L�a<%�a<�a<ۣa<ǣa<p�a<M�a<�a<��a<��a<��a<m�a<E�a<�a<�a<��a<��a<s�a<U�a<�a<�a<��a<[�a<!�a<ٟa<��a<(�a<ܞa<��a<D�a<��a<��a<T�a<�a<��a<b�a<�a<ԛa<b�a<�a<��a<S�a<ٙa<p�a<��a<��a<
�a<��a< �a<��a<�a<��a<�a<��a<'�a<��a<9�a<Ȓa<i�a<ۑa<o�a<�a<~�a<�a<y�a<�a<{�a<ލa<[�a<Ќa<]�a<�a<U�a<�a<��a<�a<��a<U�a<�a<��a<F�a<�a<��a<?�a<φa<��a<�a<݅a<c�a<�a<��a<w�a<4�a<ۃa<��a<��a<E�a<�a<�a<�a<Âa<��a<~�a<f�a<P�a<(�a<$�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<́a<́a<��a<�a<[�a<�  �  h�a<��a<͂a<�a<�a<E�a<g�a<��a<��a<�a<+�a<=�a<��a<Ȅa<#�a<e�a<ȅa<�a<��a<�a<O�a<a<5�a<��a<�a<�a<�a<E�a<��a<(�a<��a<�a<��a<ٌa<k�a<��a<L�a<��a<��a<�a<��a<$�a<��a<K�a<֒a<]�a<�a<^�a<ܔa<c�a<��a<f�a<a<8�a<��a<6�a<��a<1�a<��a<8�a<�a<*�a<қa<A�a<��a<6�a<��a<�a<i�a<��a<�a<[�a<��a<��a<H�a<]�a<۠a<�a<5�a<��a<�a< �a<c�a<��a<̢a<�a<B�a<k�a<��a<��a<ģa<ߣa<�a<'�a<�a<1�a<:�a<Y�a<f�a<��a<��a<ˤa<�a<�a<�a<,�a<C�a<V�a<Z�a<e�a<Y�a<J�a<M�a<;�a<9�a</�a<�a<�a<�a<�a<�a<�a<ݤa<��a<��a<��a<��a<��a<p�a<R�a<1�a<�a<գa<��a<u�a<N�a<��a<�a<��a<��a<M�a<1�a<�a< �a<��a<��a<k�a<D�a<�a<ߠa<��a<q�a<�a<͟a<��a<>�a<��a<��a<9�a<��a<ĝa<>�a<�a<ǜa<t�a<�a<Ûa<a�a<�a<��a<N�a<�a<i�a<�a<��a<ԗa<��a<�a<n�a<�a<v�a<��a<}�a<�a<��a<J�a<��a<S�a<ԑa<b�a<�a<v�a<��a<�a<�a<g�a<�a<k�a<�a<x�a<̋a<��a<�a<{�a<:�a<͉a<g�a<	�a<��a<@�a< �a<��a<7�a<߆a<y�a<�a<��a<N�a<$�a<��a<e�a<�a<׃a<��a<k�a<(�a<�a<��a<��a<��a<��a<��a<n�a<Q�a<?�a<�a<��a<��a<Ձa<Ёa<ǁa<��a<��a<сa<��a<ҁa<��a<�a< �a<N�a<�  �  ��a<��a<ςa<�a<�a<D�a<A�a<��a<��a<ڃa<
�a<Q�a<��a<��a<!�a<<�a<Ӆa<�a<v�a<׆a<Z�a<��a<�a<��a<�a<�a<�a<a�a<ۊa<"�a<��a<�a<{�a<�a<n�a< �a<n�a<�a<u�a<#�a<��a<0�a<ڑa<G�a<ݒa<X�a<��a<[�a<��a<]�a<��a<D�a<��a<M�a<��a</�a<��a<�a<ϙa<'�a<��a<-�a<̛a<+�a<��a<3�a<��a<	�a<a�a<؞a<�a<h�a<��a<�a<S�a<��a<֠a<�a<^�a<��a<ޡa<>�a<a�a<��a<�a<�a<D�a<f�a<��a<��a<��a<�a<ޣa<��a<�a<A�a<�a<^�a<R�a<~�a<��a<��a<Ӥa<�a<�a<�a<E�a<M�a<V�a<g�a<X�a<s�a<J�a<\�a<B�a<�a<.�a<
�a<�a<�a<��a<Ӥa<ݤa<�a<��a<̤a<��a<��a<l�a<J�a</�a<ۣa<֣a<��a<b�a<.�a<�a<ڢa<��a<��a<%�a<;�a<��a<ҡa<��a<��a<h�a<*�a<�a<ڠa<��a<k�a</�a<��a<��a<]�a<�a<��a<a�a<�a<ŝa<`�a<)�a<��a<��a<-�a<Λa<��a<�a<��a<H�a<ߙa<f�a<Ҙa<{�a<ߗa<p�a<ݖa<��a<֕a<o�a<��a<_�a<"�a<��a<"�a<��a<M�a<��a<Z�a<�a<r�a<��a<w�a<�a<|�a<��a<��a<ߌa<��a<�a<��a<�a<��a<9�a<ˉa<��a<�a<a<d�a<��a<��a<2�a<݆a<f�a<�a<��a<G�a<��a<��a<v�a<�a<܃a<|�a<Z�a<=�a<��a<��a<Ăa<��a<r�a<��a<f�a<L�a<B�a<�a<#�a<�a<��a<فa<��a<΁a<��a<؁a<ǁa<�a<�a<�a<G�a<H�a<�  �  y�a<��a<ła<��a<�a<A�a<h�a<y�a<��a<Ӄa< �a<$�a<l�a<��a<��a<K�a<��a<�a<e�a<܆a<[�a<��a<@�a<��a<�a<��a<�a<Z�a<Ŋa<9�a<��a<'�a<��a<*�a<}�a<�a<��a<�a<��a<$�a<��a<*�a<Ña<N�a<֒a<k�a<ʓa<n�a<єa<R�a<וa<,�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<I�a<ƛa<5�a<̜a<�a<��a<�a<e�a<Ğa<�a<n�a<��a<�a<T�a<��a<ՠa<�a<��a<��a<�a<6�a<t�a<��a<�a<�a<K�a<s�a<~�a<��a<��a<�a<�a<�a<�a<
�a<�a<8�a<I�a<g�a<}�a<��a<¤a< �a<�a<)�a<K�a<C�a<g�a<]�a<^�a<[�a<V�a<X�a<K�a<I�a<C�a<+�a<��a<�a<�a<��a<�a<�a<̤a<��a<��a<��a<w�a<D�a<,�a<�a<��a<��a<[�a<$�a<ߢa<��a<��a<^�a<4�a<�a<֡a<��a<��a<��a<V�a<O�a<�a<�a<��a<g�a<(�a<��a<��a<V�a<�a<��a<��a<�a<��a<��a<-�a<�a<��a<2�a<ɛa<z�a<�a<��a<\�a<șa<y�a<�a<p�a<��a<X�a<Жa<L�a<ѕa<Q�a<ڔa<b�a<�a<v�a<�a<��a<G�a<Ǒa<r�a<אa<��a<��a<{�a<��a<o�a<��a<��a<�a<��a<"�a<��a<�a<Պa<J�a<�a<}�a<�a<��a<W�a<�a<��a<?�a<Ɔa<��a<�a<��a<R�a<�a<��a<>�a<��a<��a<t�a<C�a<�a<�a<ςa<ӂa<��a<��a<��a<[�a<^�a<7�a< �a<�a<��a<�a<�a<�a<�a<ׁa<��a<�a<�a<�a<!�a<C�a<\�a<�  �  v�a<Ăa<ɂa<�a<�a<+�a<e�a<[�a<��a<��a<�a<+�a<g�a<��a<Ԅa<\�a<��a<�a<w�a<��a<9�a<��a<3�a<��a<�a<n�a<��a<u�a<Ŋa<f�a<��a<,�a<��a<��a<��a<�a<��a<��a<��a<�a<Аa<P�a<đa<l�a<��a<g�a<ѓa<[�a<ʔa<.�a<��a<�a<��a<�a<��a<�a<��a<*�a<��a<:�a<��a<�a<��a<)�a<��a<�a<��a<�a<��a<ɞa<(�a<��a<��a<!�a<=�a<��a<�a<:�a<j�a<��a<	�a<&�a<��a<��a<��a<)�a<2�a<z�a<z�a<��a<��a<��a<��a<�a<�a<�a</�a<�a<O�a<q�a<w�a<��a<��a<٤a<�a<'�a<1�a<L�a<[�a<Y�a<��a<[�a<~�a<a�a<>�a<Q�a< �a<:�a<�a<"�a<��a<�a<�a<�a<�a<��a<Ƥa<��a<h�a<P�a<�a<��a<��a<��a<>�a<:�a<�a<��a<��a<8�a<D�a<�a<�a<ԡa<��a<x�a<=�a<B�a<��a<�a<��a<x�a<D�a<�a<ʟa<L�a<�a<��a<_�a<*�a<ӝa<��a<�a<�a<w�a<S�a<�a<|�a<9�a<��a<X�a<Йa<e�a<ߘa<L�a<Ηa<E�a<�a<>�a<�a<H�a<ǔa<v�a<ԓa<��a<�a<��a<"�a<��a<c�a<ܐa<��a<�a<��a<�a<��a<&�a<o�a<�a<m�a<�a<��a<3�a<��a<9�a<��a<m�a<E�a<��a<m�a<�a<��a<F�a<a<w�a<�a<��a<&�a<�a<��a<&�a<�a<��a<z�a<M�a<	�a<�a<��a<��a<}�a<��a<q�a<d�a<R�a<3�a<K�a<
�a<!�a<��a<Ձa<�a<��a<�a<ہa<��a<�a<�a<�a<B�a<��a<�  �  ��a<��a<Ђa<�a<�a<'�a<Z�a<��a<��a<a<��a<�a<T�a<��a<�a<9�a<��a<�a<L�a<Ɇa<Y�a<ȇa<!�a<��a<�a<w�a<�a<i�a<Ίa<7�a<��a<1�a<��a<!�a<��a<�a<��a<4�a<��a<+�a<��a<:�a<Αa<Q�a<ْa<U�a<ۓa<E�a<ݔa<[�a<��a<!�a<��a<�a<��a<�a<��a<��a<��a< �a<��a<0�a<̛a<F�a<��a<+�a<��a<�a<l�a<͞a<�a<x�a<ȟa<%�a<~�a<��a<�a<=�a<��a<ڡa<�a<A�a<r�a<��a<�a<�a<?�a<e�a<��a<��a<Σa<�a<ԣa<ѣa<�a<�a<
�a<(�a<?�a<P�a<d�a<��a<��a<��a<�a<(�a<'�a<N�a<N�a<e�a<i�a<f�a<[�a<b�a<T�a<^�a<N�a<>�a<+�a<$�a<�a<�a<��a<�a<Ȥa<��a<��a<��a<c�a<N�a<�a<��a<ԣa<��a<J�a<�a<΢a<��a<z�a<N�a<!�a<�a<ˡa<��a<��a<��a<q�a<0�a<�a<٠a<��a<q�a<8�a<�a<��a<`�a<�a<ߞa<��a<2�a<ٝa<��a<P�a<��a<��a<=�a<ٛa<��a<�a<��a<F�a<ڙa<P�a<�a<x�a<�a<M�a<��a<8�a<��a<F�a<̔a<J�a<֓a<\�a<��a<��a<M�a<ّa<J�a<�a<n�a<��a<��a<�a<}�a<�a<��a<�a<��a< �a<��a<6�a<̊a<q�a<��a<��a<�a<��a<e�a<��a<��a<1�a<φa<c�a<�a<��a<=�a<τa<w�a<&�a<��a<��a<j�a<,�a<��a<ւa<Ȃa<ǂa<��a<��a<f�a<g�a<E�a<?�a<+�a<�a<��a<��a<�a<��a<�a<�a<�a<��a<�a<*�a<*�a<I�a<X�a<�  �  �a<�a<9�a<:�a<R�a<��a<��a<a<لa<+�a<R�a<��a<υa<�a<H�a<��a<�a<]�a<��a<&�a<k�a<��a<d�a<�a</�a<ˊa<C�a<��a<>�a<f�a<�a<_�a<ҍa<?�a<ʎa<j�a<��a<F�a<��a<t�a<ۑa<e�a<
�a<c�a<�a<W�a<��a<j�a<�a<B�a<��a<M�a<��a<K�a<��a<�a<��a<'�a<��a<�a<��a<�a<��a<+�a<��a<"�a<o�a<�a<S�a<ϟa<"�a<\�a<۠a<�a<L�a<��a<�a<0�a<`�a<��a<�a<S�a<X�a<ˣa<أa<�a<K�a<9�a<��a<��a<��a<��a<դa<��a<��a<$�a<�a</�a<<�a<z�a<��a<��a<ͥa<ɥa<�a<�a<,�a<=�a<D�a<{�a<P�a<��a<K�a<a�a<_�a<0�a<6�a<"�a<F�a<�a<�a<�a<��a<��a<��a<��a<��a<��a<f�a<5�a<�a<�a<��a<o�a<a�a<%�a<�a<̣a<~�a<^�a<0�a<(�a<��a<Тa<��a<`�a<V�a<+�a<�a<��a<��a<|�a< �a<�a<��a<x�a<�a<��a<d�a<%�a<��a<q�a</�a<ǝa<��a<2�a<ڜa<��a<�a<Лa<+�a<ښa<^�a<�a<Q�a<٘a<q�a<ܗa<��a<��a<a�a<�a<��a<&�a<��a<5�a<��a<4�a<�a<t�a<�a<v�a<;�a<��a<A�a<��a<(�a<ڎa<%�a<��a<<�a<��a<p�a<�a<��a<�a<�a<L�a<$�a<��a<K�a<�a<U�a<�a<��a<M�a<͆a<��a<E�a<�a<��a<G�a<�a<��a<��a<��a<E�a<1�a<�a<�a<ڃa<ăa<��a<��a<��a<l�a<��a<F�a<T�a<N�a<!�a<.�a<'�a<[�a<@�a<J�a<T�a<��a<��a<��a<�  �  Ӄa<�a< �a<8�a<r�a<}�a<��a<݄a<�a<#�a<K�a<��a<��a<�a<_�a<��a<�a<Q�a<��a<'�a<��a<�a<j�a<؉a<W�a<��a<+�a<��a<�a<z�a<�a<[�a<�a<V�a<��a<;�a<a<Y�a<֐a<L�a<ёa<[�a<ےa<d�a<��a<p�a<��a<d�a<�a<m�a<�a<:�a<��a<&�a<��a<.�a<��a<)�a<��a<%�a<��a<?�a<��a<3�a<��a<%�a<��a<��a<O�a<��a<
�a<Y�a<��a<�a<`�a<��a<ءa<�a<r�a<¢a<�a<-�a<g�a<��a<��a<�a<.�a<a�a<{�a<��a<��a<ؤa<�a<�a<��a<�a<0�a<E�a<]�a<j�a<��a<��a<��a<��a<�a<"�a<&�a<S�a<J�a<`�a<O�a<Y�a<X�a<Y�a<L�a<V�a<K�a<+�a<�a<�a<�a<�a<�a<�a<ɥa<��a<��a<��a<d�a<V�a<�a<��a<ͤa<��a<Y�a<�a<�a<��a<��a<u�a<K�a<�a<�a<��a<��a<��a<h�a<1�a<�a<�a<��a<e�a<�a<�a<��a<W�a<�a<՟a<{�a<�a<ɞa<�a<B�a<�a<��a<(�a<Мa<l�a<�a<��a<D�a<�a<Y�a<�a<|�a<��a<^�a<�a<\�a<�a<v�a< �a<��a<�a<��a<$�a<ѓa<d�a<�a<s�a<�a<��a<�a<��a<�a<��a<%�a<��a<?�a<Ӎa<J�a<Ќa<Z�a< �a<��a<$�a<��a<[�a<��a<��a<3�a<ӈa<~�a<�a<��a<\�a<�a<��a<3�a<��a<��a<\�a<�a<݄a<��a<j�a<F�a<"�a<!�a<�a<�a<��a<ăa<��a<��a<j�a<b�a<S�a<L�a<<�a<H�a<C�a<0�a<,�a<=�a<_�a<x�a<|�a<��a<��a<�  �  ƃa<�a<�a<9�a<s�a<r�a<��a<��a<��a<�a<q�a<��a<˅a<�a<9�a<��a<��a<t�a<̇a<�a<��a<݈a<��a<ĉa<e�a<��a<8�a<��a< �a<��a<یa<a�a<ʍa<G�a<Ύa<C�a<Џa<-�a<ސa<>�a<�a<x�a<ߒa<��a<ߓa<}�a<�a<i�a<ܕa<@�a<Ֆa<=�a<�a<0�a<��a<'�a<��a<8�a<��a<S�a<��a<3�a<��a<�a<��a<�a<��a<��a<s�a<��a<"�a<z�a<��a<�a<7�a<��a<�a<+�a<f�a<��a<��a<�a<��a<��a<�a<�a< �a<r�a<h�a<��a<��a<��a<פa<��a<�a<�a<:�a<'�a<_�a<v�a<��a<̥a<��a<�a<�a<"�a<!�a<O�a<Q�a<O�a<z�a<M�a<x�a<Z�a<E�a<N�a<�a<?�a<!�a<$�a<�a<�a<�a<ߥa<�a<��a<��a<��a<e�a<W�a<	�a<��a<��a<��a<S�a<D�a<�a<ȣa<��a<N�a<S�a<�a<�a<ݢa<��a<��a<=�a<G�a<�a<�a<��a<r�a<:�a<ڠa<àa<F�a<�a<��a<l�a<)�a<Ҟa<��a<�a<�a<t�a<>�a<�a<p�a<6�a<��a<P�a<Қa<^�a<ޙa<O�a<�a<a�a<�a<f�a<��a<o�a<�a<��a<	�a<ǔa<*�a<ēa<@�a<Ԓa<{�a<��a<��a<�a<��a<'�a<��a<F�a<��a<L�a<��a<P�a<،a<l�a<��a<~�a</�a<��a<��a<��a<��a<I�a<Ĉa<��a<�a<ća<5�a<�a<��a<H�a<�a<��a<f�a<��a<߄a<��a<}�a<p�a<�a<�a<Ճa<�a<��a<��a<��a<��a<��a<V�a<s�a<M�a<5�a<@�a<�a<C�a<6�a<P�a<:�a<i�a<w�a<��a<Ӄa<�  �  уa<�a<�a<N�a<_�a<�a<Äa<҄a<�a<4�a<Y�a<��a<ׅa<�a<j�a<��a<�a<Z�a<ˇa<6�a<��a<��a<��a<ωa<P�a<Êa<(�a<��a<�a<p�a<ތa<l�a<Ía<F�a<��a<+�a<��a<0�a<ʐa<K�a<ʑa<P�a<ؒa<l�a<�a<��a<�a<y�a<��a<b�a<�a<Z�a<��a<9�a<��a<7�a<��a<;�a<��a<+�a<��a<G�a<��a<;�a<��a<�a<��a<�a<U�a<��a<��a<S�a<��a<�a<:�a<��a<ȡa<�a<g�a<��a<��a<�a<_�a<��a<ƣa<�a<7�a<]�a<o�a<��a<��a<ݤa<�a<��a<��a< �a<;�a<T�a<c�a<~�a<��a<��a<եa< �a<�a<3�a</�a<=�a<b�a<R�a<]�a<Y�a<K�a<I�a<S�a<<�a<'�a<*�a<
�a<�a<��a<��a<��a<Хa<��a<��a<��a<��a<z�a<C�a<�a<	�a<äa<��a<j�a<,�a<��a<ԣa<��a<��a<T�a<'�a<�a<ܢa<��a<��a<X�a<P�a<��a<١a<��a<b�a<�a<۠a<��a<H�a<�a<��a<k�a<�a<��a<|�a<�a<۝a<��a<!�a<Ɯa<i�a<�a<��a<T�a<˚a<m�a<��a<q�a<�a<~�a<�a<o�a< �a<�a<�a<��a<�a<��a<@�a<ٓa<b�a<�a<��a<��a<��a<�a<��a<�a<��a<�a<��a<=�a<��a<I�a<��a<W�a<��a<z�a<3�a<��a<S�a<�a<��a<6�a<܈a<y�a<	�a<̇a<Q�a<	�a<��a<N�a<�a<��a<f�a<(�a<�a<��a<u�a<M�a<:�a<)�a<��a<��a<ǃa<��a<��a<��a<x�a<b�a<F�a<<�a<C�a<.�a< �a</�a< �a<=�a<C�a<[�a<��a<��a<��a<�  �  �a<�a<�a<9�a<^�a<��a<��a<�a<��a<5�a<k�a<��a<��a<�a<��a<��a<�a<e�a<؇a<%�a<��a<�a<g�a<�a<I�a<��a<$�a<��a<�a<m�a<ތa<9�a<��a<>�a<��a<2�a<��a<B�a<��a<@�a<͑a<`�a<�a<Z�a<�a<f�a<��a<s�a<�a<m�a<ɖa<e�a<ȗa<^�a<��a<D�a<ʙa<)�a<Ϛa<2�a<Λa<'�a<��a<+�a<��a<$�a<��a<��a<G�a<��a<�a<V�a<��a<ؠa<B�a<~�a<ʡa<�a<Z�a<��a<Ǣa<�a<\�a<��a<Σa<��a<3�a<U�a<��a<��a<��a<դa<֤a<�a<�a<2�a<�a<n�a<^�a<��a<��a<��a<ݥa<�a<�a<�a<@�a<@�a<I�a<Y�a<O�a<o�a<O�a<K�a<7�a<�a<:�a<�a<�a<��a<	�a<ڥa<ԥa<եa<��a<ͥa<��a<��a<e�a<B�a<0�a<�a<Ҥa<��a<k�a<=�a<�a<ݣa<��a<��a<9�a<6�a<��a<�a<��a<��a<e�a</�a<�a<ҡa<��a<^�a<�a<��a<��a<H�a<�a<��a<c�a<�a<��a<f�a<+�a<��a<v�a<$�a<՜a<��a<�a<��a<9�a<ښa<h�a<�a<|�a<�a<��a<��a<��a<�a<��a<�a<��a<6�a<��a<O�a<��a<c�a<�a<z�a<�a<��a<�a<��a<*�a<��a<"�a<��a<�a<��a<1�a<��a<L�a<�a<u�a<��a<��a<P�a<
�a<��a</�a<؈a<r�a<#�a<��a<V�a<�a<��a<]�a<�a<��a<J�a<B�a<߄a<��a<��a<`�a<B�a<�a<�a<݃a<؃a<��a<��a<��a<k�a<x�a<J�a<>�a<&�a<�a<3�a<�a<*�a<(�a<P�a<A�a<a�a<��a<��a<�  �  ��a<��a<�a<4�a<`�a<��a<��a<�a<
�a<9�a<��a<��a<��a<*�a<�a<��a<.�a<o�a<�a<0�a<��a<�a<�a<ۉa<P�a<��a<.�a<��a<�a<a�a<ӌa<K�a<a<�a<��a<4�a<��a<"�a<��a<<�a<��a<H�a<Вa<k�a<�a<l�a<�a<~�a<��a<��a<ۖa<l�a<ٗa<S�a<Ҙa<S�a<Йa<J�a<̚a<@�a<כa<<�a<՜a<@�a<��a<�a<��a<�a<W�a<��a<��a<F�a<��a<�a<.�a<^�a<͡a<�a<8�a<��a<ۢa<�a<K�a<��a<ѣa<
�a<"�a<_�a<x�a<��a<ʤa<�a<�a<�a<�a<A�a<E�a<d�a<|�a<��a<��a<ѥa<�a<�a<�a<*�a<9�a<F�a<H�a<T�a<`�a<=�a<B�a<;�a<;�a<.�a<�a<��a<�a<�a<ܥa<�a<ݥa<ťa<��a<��a<��a<��a<`�a<D�a<"�a<�a<ݤa<��a<p�a<T�a<�a<��a<��a<��a<\�a<K�a<�a<��a<��a<��a<u�a<F�a<�a<١a<��a<h�a<%�a<��a<��a<=�a<��a<��a<>�a<��a<a<F�a<�a<Ɲa<r�a<�a<��a<a�a<�a<��a<?�a<ךa<s�a<��a<��a<��a<��a<�a<��a<�a<��a<"�a<��a<3�a<��a<Y�a<͓a<x�a<��a<��a<�a<��a<�a<��a<�a<��a<�a<��a<$�a<��a<�a<Ča<C�a<Ƌa<z�a<�a<��a<>�a<ۉa<��a<<�a<ƈa<|�a<�a<Ƈa<k�a<�a<��a<l�a< �a<ʅa<q�a<8�a<��a<фa<��a<u�a<F�a<�a<�a<�a<уa<��a<��a<��a<{�a<F�a<>�a<.�a<*�a<�a<�a<��a<+�a<�a<#�a<L�a<j�a<|�a<��a<�  �  ��a<�a<��a<M�a<t�a<x�a<Ʉa<܄a<.�a<B�a<��a<��a<�a<B�a<��a<܆a<1�a<��a<�a<D�a<��a<�a<��a<͉a<i�a<��a<�a<��a<�a<o�a<��a<9�a<��a< �a<��a<�a<��a<�a<��a<%�a<��a<M�a<ʒa<j�a<ӓa<��a<�a<v�a<��a<x�a<��a<i�a<�a<\�a<�a<Z�a<ٙa<e�a<Ԛa<U�a<Лa<U�a<Μa<;�a<��a<�a<��a<ܞa<Q�a<��a<��a<C�a<��a<֠a<�a<s�a<��a<�a<B�a<w�a<Ţa<�a<W�a<��a<ãa<��a<&�a<}�a<k�a<��a<��a<�a<��a<�a<(�a<A�a<`�a<n�a<��a<��a<��a<إa<�a<�a<�a<7�a<+�a<M�a<f�a<7�a<\�a<9�a<Q�a</�a<+�a<�a<�a<�a<�a<�a<�a<̥a<ϥa<��a<ƥa<��a<��a<d�a<x�a<X�a<�a<�a<ͤa<Ĥa<x�a<[�a<�a<��a<Σa<��a<x�a<M�a<�a<��a<ɢa<��a<f�a<Q�a<��a<�a<��a<L�a<�a<Ǡa<��a<*�a<�a<��a<E�a<�a<��a<Y�a<��a<��a<[�a<�a<a<[�a<�a<��a<g�a<њa<j�a<��a<��a<�a<��a<�a<��a<'�a<��a<*�a<��a<;�a<ɔa<R�a<�a<r�a<�a<��a<��a<��a<�a<��a<�a<��a<�a<��a<�a<��a<%�a<��a<4�a<Ћa<X�a<��a<��a<K�a<�a<��a<&�a<ˈa<��a<�a<χa<`�a<�a<��a<b�a<�a<ʅa<��a<A�a<�a<؄a<��a<|�a<I�a<B�a<�a<��a<a<��a<��a<j�a<w�a<A�a<L�a<"�a<�a<�a<	�a<�a<�a<�a<)�a<3�a<[�a<k�a<��a<�  �  ��a<�a<	�a<5�a<_�a<��a<̄a<ބa<$�a<U�a<��a<υa<��a<;�a<��a<Άa<2�a<��a<��a<O�a<��a<
�a<��a<�a<I�a<��a< �a<��a<��a<H�a<��a<1�a<��a<�a<��a<�a<��a<�a<��a<1�a<��a<D�a<Ԓa<a�a<ݓa<t�a<�a<��a<�a<q�a<�a<x�a<��a<{�a<ݘa<m�a<��a<R�a<�a<k�a<�a<T�a<˜a<I�a<a<�a<��a<�a<O�a<��a<��a<-�a<��a<��a<�a<Y�a<��a<�a<0�a<l�a<��a<�a<3�a<��a<��a< �a<+�a<U�a<��a<��a<äa<�a<�a<&�a<@�a<J�a<N�a<��a<��a<��a<ӥa<�a<��a<�a<�a<=�a<J�a<?�a<M�a<G�a<P�a<I�a<6�a<�a<)�a<�a<�a<�a<�a<Хa<ݥa<��a<ǥa<��a<��a<��a<��a<x�a<a�a<C�a<0�a<�a<Ϥa<��a<��a<i�a<9�a<��a<ƣa<��a<i�a<N�a<4�a<	�a<Ԣa<��a<j�a<T�a<�a<ѡa<��a<Z�a<�a<Ԡa<l�a<)�a<ݟa<y�a<<�a<�a<��a<@�a<��a<��a<f�a<��a<��a<e�a<�a<��a<H�a<Ϛa<{�a<�a<��a<�a<��a<*�a<��a<�a<��a<G�a<��a<N�a<ޔa<e�a<�a<n�a<�a<��a<�a<��a<	�a<��a<�a<��a<��a<��a<��a<��a<�a<��a<,�a<��a<M�a<�a<��a<'�a<�a<��a<1�a<Јa<r�a<�a<чa<d�a<�a<��a<w�a<+�a<Ӆa<z�a<e�a<�a<фa<��a<��a<^�a<6�a<�a<�a<�a<��a<��a<z�a<k�a<R�a<2�a<�a<�a<�a<�a<�a<��a<��a<%�a<!�a<T�a<_�a<��a<�  �  ��a<΃a<�a<3�a<f�a<��a<��a<�a<(�a<c�a<��a<ƅa<%�a<T�a<��a<�a<[�a<��a<��a<^�a<��a<:�a<|�a<�a<H�a<��a<"�a<u�a<�a<6�a<��a<�a<��a<��a<o�a<�a<Z�a<�a<{�a<#�a<��a<6�a<��a<L�a<�a<i�a<��a<{�a<�a<��a<�a<��a<�a<{�a<��a<t�a<��a<p�a<��a<W�a<�a<c�a<�a<X�a<��a<(�a<��a<�a<<�a<��a<�a<�a<��a<��a<�a<4�a<��a<סa<�a<w�a<��a<��a<!�a<��a<��a<��a<+�a<P�a<��a<��a<�a<��a<�a<)�a<0�a<n�a<m�a<��a<��a<ƥa<ʥa<٥a<�a<�a<E�a<.�a<A�a<J�a<I�a<W�a<8�a<<�a<,�a<�a<�a<��a<��a<ƥa<��a<��a<ťa<��a<��a<��a<��a<��a<{�a<��a<_�a<J�a<.�a<�a<�a<��a<��a<^�a<0�a<"�a<�a<��a<��a<x�a<$�a<�a<�a<��a<��a<D�a<�a<ѡa<��a<\�a<�a<àa<Z�a<$�a<ʟa<��a<�a<˞a<��a<�a<��a<��a<Y�a<�a<��a<P�a<��a<��a<<�a<�a<o�a<	�a<��a<�a<��a<�a<��a<;�a<��a<F�a<̕a<\�a<ʔa<m�a<��a<��a<�a<��a<�a<��a<�a<��a<��a<��a<�a<��a<�a<��a<�a<��a<�a<��a<X�a<ފa<��a<�a<ډa<p�a<)�a<ψa<m�a<&�a<��a<��a<(�a<φa<z�a<�a<��a<��a<d�a<�a<��a<��a<~�a<h�a<@�a<9�a<�a<كa<��a<��a<��a<T�a<E�a<(�a<�a<�a<�a<�a<˂a<�a<݂a<�a< �a<?�a<Z�a<��a<�  �  ��a<�a<��a<7�a<x�a<��a<Ȅa<��a<'�a<`�a<��a<ޅa<�a<h�a<��a<�a<G�a<��a<�a<\�a<��a<#�a<��a<�a<b�a<��a<�a<��a<ًa<W�a<��a<�a<y�a<��a<o�a<��a<u�a<�a<s�a<�a<��a<=�a<��a<f�a<ԓa<r�a< �a<��a<��a<��a<�a<��a<�a<}�a<�a<{�a<��a<��a<�a<��a<�a<b�a<֜a<D�a<��a<+�a<��a<ٞa<M�a<��a<�a<7�a<x�a<��a<��a<J�a<��a<ϡa<�a<T�a<��a<��a<E�a<r�a<ȣa<��a<�a<l�a<��a<��a<Ѥa<�a<�a<7�a<T�a<Y�a<��a<��a<��a<ɥa<إa<
�a<�a<�a<*�a<4�a<C�a<U�a<N�a<;�a<Z�a<,�a<5�a< �a<
�a<�a<�a<ޥa<ӥa<ťa<��a<��a<��a<��a<��a<��a<��a<l�a<b�a<\�a<,�a<�a<�a<��a<��a<��a<H�a<�a<��a<��a<��a<c�a<D�a<�a<�a<��a<��a<R�a<�a<�a<��a<P�a<�a<��a<|�a<�a<��a<d�a<�a<˞a<��a<3�a<ݝa<��a<J�a< �a<��a<O�a<�a<��a<F�a<�a<w�a<��a<��a< �a<��a<K�a<��a<K�a<Öa<F�a<�a<X�a<��a<t�a<�a<z�a<��a<��a<�a<��a<��a<��a<�a<��a<�a<x�a<�a<m�a<��a<��a<�a<��a<5�a<͊a<��a<9�a<ˉa<��a<*�a<Èa<��a< �a<Їa<r�a<�a<̆a<��a<>�a<�a<��a<\�a<1�a<��a<��a<��a<h�a<A�a<�a<��a<ۃa<ƃa<��a<m�a<v�a<5�a<0�a<�a<��a<߂a<�a<�a<�a<�a< �a<�a</�a<]�a<��a<�  �  ��a<�a<��a<L�a<c�a<��a<�a<�a<X�a<k�a<��a<�a<�a<{�a<��a<�a<>�a<��a<�a<q�a<�a<�a<��a<�a<T�a<��a<�a<{�a<��a<A�a<��a<1�a<|�a<�a<h�a<͎a<v�a<��a<��a<
�a<��a<�a<��a<]�a<Гa<��a<�a<��a<�a<��a<3�a<~�a<�a<�a<�a<��a<�a<��a<�a<��a<�a<��a<��a<[�a<۝a<�a<��a<؞a<C�a<w�a<ȟa<#�a<g�a<Ҡa<�a<H�a<o�a<áa<�a<N�a<Ģa<֢a<.�a<P�a<��a<�a<*�a<f�a<{�a<դa<Ѥa<�a<*�a<*�a<h�a<U�a<��a<��a<¥a<ȥa<�a<��a<�a<G�a<&�a<U�a<P�a<B�a<e�a</�a<R�a<�a<�a<�a<�a<�a<٥a<ޥa<��a<ĥa<��a<��a<��a<��a<��a<i�a<��a<^�a<w�a<G�a<2�a<.�a<�a<�a<��a<x�a<S�a<�a<�a<ͣa<��a<Z�a<W�a<�a<��a<ڢa<z�a<p�a<�a<ݡa<��a<B�a<�a<��a<e�a<��a<ݟa<g�a<�a<Þa<[�a<4�a<ɝa<��a<@�a<�a<��a<2�a<�a<��a<Z�a<̚a<��a<�a<��a<L�a<��a<L�a<��a<K�a<ٖa<^�a<�a<U�a<�a<i�a<�a<��a<�a<��a<��a<��a<��a<��a<�a<e�a<�a<f�a<	�a<\�a<��a<g�a<�a<��a<.�a<��a<j�a<!�a<��a<p�a<�a<Έa<��a<�a<��a<s�a<D�a<�a<{�a<S�a<݅a<Åa<t�a<C�a<��a<ʄa<��a<k�a<q�a<�a<�a<�a<��a<��a<a�a<m�a<�a<�a<��a<��a<��a<тa<�a<��a<��a<�a<�a<@�a<F�a<{�a<�  �  ��a<؃a<��a<G�a<d�a<��a<��a<�a<2�a<v�a<��a<��a<4�a<g�a<��a<�a<l�a<Ça<	�a<i�a<ƈa<#�a<~�a<�a<J�a<Ċa<�a<}�a<�a<L�a<��a<�a<l�a<�a<g�a<�a<j�a<܏a<k�a<��a<��a<9�a<Œa<O�a<�a<v�a<��a<�a<��a<��a<�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<��a<h�a<�a<E�a<��a<*�a<��a<�a<8�a<��a<�a<-�a<]�a<��a<�a<:�a<��a<ơa<�a<B�a<��a<Ԣa<<�a<��a<��a<�a<8�a<Y�a<��a<��a<Ӥa<��a<�a<6�a<c�a<��a<��a<��a<��a<ۥa<��a<��a<�a<"�a<2�a<*�a<I�a<I�a<Y�a<A�a<=�a<>�a<7�a<�a<�a<�a<ѥa<ץa<ɥa<��a<��a<��a<��a<��a<��a<��a<��a<l�a<r�a<H�a<6�a<�a<�a<Ȥa<��a<|�a<e�a<1�a<�a<ãa<��a<��a<\�a<�a<�a<��a<��a<F�a<�a<ӡa<��a<B�a<	�a< a<q�a<��a<��a<W�a<
�a<Þa<t�a<(�a<ŝa<|�a<.�a<��a<��a<V�a<��a<��a<J�a<ܚa<s�a<��a<��a<&�a<��a<@�a<ۗa<T�a<˖a<V�a<�a<~�a<��a<w�a<��a<��a<��a<��a<�a<��a<�a<��a<�a<��a<��a<\�a<ݍa<W�a<�a<z�a<�a<��a<"�a<͊a<g�a<0�a<ىa<x�a<�a<݈a<v�a<)�a<ȇa<t�a<'�a<Նa<��a<N�a<�a<��a<l�a<-�a<�a<�a<��a<x�a<L�a<&�a<�a<��a<��a<��a<t�a<Y�a<G�a<2�a<�a<߂a<ւa<ʂa<܂a<߂a<�a<�a<�a<�a<N�a<��a<�  �  ��a<Ѓa<	�a<$�a<j�a<��a<��a<@�a<�a<��a<��a<څa<�a<n�a<݆a<��a<Y�a<��a<!�a<q�a<��a<_�a<~�a<�a<?�a<��a<�a<r�a<ŋa<#�a<��a<�a<��a<��a<J�a<юa<X�a<��a<o�a<�a<��a<�a<��a<M�a<�a<Q�a<�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<(�a<{�a< �a<o�a<"�a<f�a<��a<i�a<Ýa<J�a<o�a<�a<8�a<��a<��a<�a<l�a<��a<�a<3�a<n�a<��a<�a<g�a<��a<�a<�a<X�a<��a<�a<+�a<D�a<��a<��a<�a<��a<"�a<Z�a<B�a<o�a<x�a<ɥa<��a<åa<�a<�a<1�a<�a<j�a<6�a<a�a<V�a<2�a<O�a<5�a<)�a<��a<�a<��a<�a<�a<��a<��a<��a<��a<��a<��a<��a<p�a<�a<}�a<w�a<O�a<N�a<Q�a<�a<0�a<��a<��a<��a<D�a<�a<��a<�a<��a<u�a<7�a<2�a<��a<��a<��a<F�a<9�a<ȡa<��a<H�a<��a<��a<G�a<�a<��a<y�a<�a<��a<`�a<�a<�a<��a<@�a<�a<y�a<J�a<��a<��a<$�a<��a<��a<�a<Ùa<�a<ݘa<2�a<a<C�a<�a<y�a<וa<g�a<�a<��a<��a<��a<!�a<��a<3�a<u�a<�a<��a<��a<S�a<܎a<k�a<֍a<z�a<�a<f�a<�a<��a<H�a<Ŋa<|�a<
�a<��a<p�a<�a<Јa<a�a<E�a<Ƈa<��a<*�a<߆a<��a<,�a<��a<��a<��a<<�a<��a<ʄa<��a<��a<9�a<_�a<��a<��a<ǃa<��a<��a<P�a<2�a<��a<�a<�a<�a<��a<��a<ɂa<ǂa<��a<�a<'�a<U�a<W�a<�  �  ��a<؃a<��a<G�a<d�a<��a<��a<�a<2�a<v�a<��a<��a<4�a<g�a<��a<�a<l�a<Ça<	�a<i�a<ƈa<#�a<~�a<�a<J�a<Ċa<�a<}�a<�a<L�a<��a<�a<l�a<�a<g�a<�a<j�a<܏a<k�a<��a<��a<9�a<Œa<O�a<�a<v�a<��a<�a<��a<��a<�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<��a<h�a<�a<E�a<��a<*�a<��a<�a<8�a<��a<�a<-�a<]�a<��a<�a<:�a<��a<ơa<�a<B�a<��a<Ԣa<<�a<��a<��a<�a<8�a<Y�a<��a<��a<Ӥa<��a<�a<6�a<c�a<��a<��a<��a<��a<ۥa<��a<��a<�a<"�a<2�a<*�a<I�a<I�a<Y�a<A�a<=�a<>�a<7�a<�a<�a<�a<ѥa<ץa<ɥa<��a<��a<��a<��a<��a<��a<��a<��a<l�a<r�a<H�a<6�a<�a<�a<Ȥa<��a<|�a<e�a<1�a<�a<ãa<��a<��a<\�a<�a<�a<��a<��a<F�a<�a<ӡa<��a<B�a<	�a< a<q�a<��a<��a<W�a<
�a<Þa<t�a<(�a<ŝa<|�a<.�a<��a<��a<V�a<��a<��a<J�a<ܚa<s�a<��a<��a<&�a<��a<@�a<ۗa<T�a<˖a<V�a<�a<~�a<��a<w�a<��a<��a<��a<��a<�a<��a<�a<��a<�a<��a<��a<\�a<ݍa<W�a<�a<z�a<�a<��a<"�a<͊a<g�a<0�a<ىa<x�a<�a<݈a<v�a<)�a<ȇa<t�a<'�a<Նa<��a<N�a<�a<��a<l�a<-�a<�a<�a<��a<x�a<L�a<&�a<�a<��a<��a<��a<t�a<Y�a<G�a<2�a<�a<߂a<ւa<ʂa<܂a<߂a<�a<�a<�a<�a<N�a<��a<�  �  ��a<�a<��a<L�a<c�a<��a<�a<�a<X�a<k�a<��a<�a<�a<{�a<��a<�a<>�a<��a<�a<q�a<�a<�a<��a<�a<T�a<��a<�a<{�a<��a<A�a<��a<1�a<|�a<�a<h�a<͎a<v�a<��a<��a<
�a<��a<�a<��a<]�a<Гa<��a<�a<��a<�a<��a<3�a<~�a<�a<�a<�a<��a<�a<��a<�a<��a<�a<��a<��a<[�a<۝a<�a<��a<؞a<C�a<w�a<ȟa<#�a<g�a<Ҡa<�a<H�a<o�a<áa<�a<N�a<Ģa<֢a<.�a<P�a<��a<�a<*�a<f�a<{�a<դa<Ѥa<�a<*�a<*�a<h�a<U�a<��a<��a<¥a<ȥa<�a<��a<�a<G�a<&�a<U�a<P�a<B�a<e�a</�a<R�a<�a<�a<�a<�a<�a<٥a<ޥa<��a<ĥa<��a<��a<��a<��a<��a<i�a<��a<^�a<w�a<G�a<2�a<.�a<�a<�a<��a<x�a<S�a<�a<�a<ͣa<��a<Z�a<W�a<�a<��a<ڢa<z�a<p�a<�a<ݡa<��a<B�a<�a<��a<e�a<��a<ݟa<g�a<�a<Þa<[�a<4�a<ɝa<��a<@�a<�a<��a<2�a<�a<��a<Z�a<̚a<��a<�a<��a<L�a<��a<L�a<��a<K�a<ٖa<^�a<�a<U�a<�a<i�a<�a<��a<�a<��a<��a<��a<��a<��a<�a<e�a<�a<f�a<	�a<\�a<��a<g�a<�a<��a<.�a<��a<j�a<!�a<��a<p�a<�a<Έa<��a<�a<��a<s�a<D�a<�a<{�a<S�a<݅a<Åa<t�a<C�a<��a<ʄa<��a<k�a<q�a<�a<�a<�a<��a<��a<a�a<m�a<�a<�a<��a<��a<��a<тa<�a<��a<��a<�a<�a<@�a<F�a<{�a<�  �  ��a<�a<��a<7�a<x�a<��a<Ȅa<��a<'�a<`�a<��a<ޅa<�a<h�a<��a<�a<G�a<��a<�a<\�a<��a<#�a<��a<�a<b�a<��a<�a<��a<ًa<W�a<��a<�a<y�a<��a<o�a<��a<u�a<�a<s�a<�a<��a<=�a<��a<f�a<ԓa<r�a< �a<��a<��a<��a<�a<��a<�a<}�a<�a<{�a<��a<��a<�a<��a<�a<b�a<֜a<D�a<��a<+�a<��a<ٞa<M�a<��a<�a<7�a<x�a<��a<��a<J�a<��a<ϡa<�a<T�a<��a<��a<E�a<r�a<ȣa<��a<�a<l�a<��a<��a<Ѥa<�a<�a<7�a<T�a<Y�a<��a<��a<��a<ɥa<إa<
�a<�a<�a<*�a<4�a<C�a<U�a<N�a<;�a<Z�a<,�a<5�a< �a<
�a<�a<�a<ޥa<ӥa<ťa<��a<��a<��a<��a<��a<��a<��a<l�a<b�a<\�a<,�a<�a<�a<��a<��a<��a<H�a<�a<��a<��a<��a<c�a<D�a<�a<�a<��a<��a<R�a<�a<�a<��a<P�a<�a<��a<|�a<�a<��a<d�a<�a<˞a<��a<3�a<ݝa<��a<J�a< �a<��a<O�a<�a<��a<F�a<�a<w�a<��a<��a< �a<��a<K�a<��a<K�a<Öa<F�a<�a<X�a<��a<t�a<�a<z�a<��a<��a<�a<��a<��a<��a<�a<��a<�a<x�a<�a<m�a<��a<��a<�a<��a<5�a<͊a<��a<9�a<ˉa<��a<*�a<Èa<��a< �a<Їa<r�a<�a<̆a<��a<>�a<�a<��a<\�a<1�a<��a<��a<��a<h�a<A�a<�a<��a<ۃa<ƃa<��a<m�a<v�a<5�a<0�a<�a<��a<߂a<�a<�a<�a<�a< �a<�a</�a<]�a<��a<�  �  ��a<΃a<�a<3�a<f�a<��a<��a<�a<(�a<c�a<��a<ƅa<%�a<T�a<��a<�a<[�a<��a<��a<^�a<��a<:�a<|�a<�a<H�a<��a<"�a<u�a<�a<6�a<��a<�a<��a<��a<o�a<�a<Z�a<�a<{�a<#�a<��a<6�a<��a<L�a<�a<i�a<��a<{�a<�a<��a<�a<��a<�a<{�a<��a<t�a<��a<p�a<��a<W�a<�a<c�a<�a<X�a<��a<(�a<��a<�a<<�a<��a<�a<�a<��a<��a<�a<4�a<��a<סa<�a<w�a<��a<��a<!�a<��a<��a<��a<+�a<P�a<��a<��a<�a<��a<�a<)�a<0�a<n�a<m�a<��a<��a<ƥa<ʥa<٥a<�a<�a<E�a<.�a<A�a<J�a<I�a<W�a<8�a<<�a<,�a<�a<�a<��a<��a<ƥa<��a<��a<ťa<��a<��a<��a<��a<��a<{�a<��a<_�a<J�a<.�a<�a<�a<��a<��a<^�a<0�a<"�a<�a<��a<��a<x�a<$�a<�a<�a<��a<��a<D�a<�a<ѡa<��a<\�a<�a<àa<Z�a<$�a<ʟa<��a<�a<˞a<��a<�a<��a<��a<Y�a<�a<��a<P�a<��a<��a<<�a<�a<o�a<	�a<��a<�a<��a<�a<��a<;�a<��a<F�a<̕a<\�a<ʔa<m�a<��a<��a<�a<��a<�a<��a<�a<��a<��a<��a<�a<��a<�a<��a<�a<��a<�a<��a<X�a<ފa<��a<�a<ډa<p�a<)�a<ψa<m�a<&�a<��a<��a<(�a<φa<z�a<�a<��a<��a<d�a<�a<��a<��a<~�a<h�a<@�a<9�a<�a<كa<��a<��a<��a<T�a<E�a<(�a<�a<�a<�a<�a<˂a<�a<݂a<�a< �a<?�a<Z�a<��a<�  �  ��a<�a<	�a<5�a<_�a<��a<̄a<ބa<$�a<U�a<��a<υa<��a<;�a<��a<Άa<2�a<��a<��a<O�a<��a<
�a<��a<�a<I�a<��a< �a<��a<��a<H�a<��a<1�a<��a<�a<��a<�a<��a<�a<��a<1�a<��a<D�a<Ԓa<a�a<ݓa<t�a<�a<��a<�a<q�a<�a<x�a<��a<{�a<ݘa<m�a<��a<R�a<�a<k�a<�a<T�a<˜a<I�a<a<�a<��a<�a<O�a<��a<��a<-�a<��a<��a<�a<Y�a<��a<�a<0�a<l�a<��a<�a<3�a<��a<��a< �a<+�a<U�a<��a<��a<äa<�a<�a<&�a<@�a<J�a<N�a<��a<��a<��a<ӥa<�a<��a<�a<�a<=�a<J�a<?�a<M�a<G�a<P�a<I�a<6�a<�a<)�a<�a<�a<�a<�a<Хa<ݥa<��a<ǥa<��a<��a<��a<��a<x�a<a�a<C�a<0�a<�a<Ϥa<��a<��a<i�a<9�a<��a<ƣa<��a<i�a<N�a<4�a<	�a<Ԣa<��a<j�a<T�a<�a<ѡa<��a<Z�a<�a<Ԡa<l�a<)�a<ݟa<y�a<<�a<�a<��a<@�a<��a<��a<f�a<��a<��a<e�a<�a<��a<H�a<Ϛa<{�a<�a<��a<�a<��a<*�a<��a<�a<��a<G�a<��a<N�a<ޔa<e�a<�a<n�a<�a<��a<�a<��a<	�a<��a<�a<��a<��a<��a<��a<��a<�a<��a<,�a<��a<M�a<�a<��a<'�a<�a<��a<1�a<Јa<r�a<�a<чa<d�a<�a<��a<w�a<+�a<Ӆa<z�a<e�a<�a<фa<��a<��a<^�a<6�a<�a<�a<�a<��a<��a<z�a<k�a<R�a<2�a<�a<�a<�a<�a<�a<��a<��a<%�a<!�a<T�a<_�a<��a<�  �  ��a<�a<��a<M�a<t�a<x�a<Ʉa<܄a<.�a<B�a<��a<��a<�a<B�a<��a<܆a<1�a<��a<�a<D�a<��a<�a<��a<͉a<i�a<��a<�a<��a<�a<o�a<��a<9�a<��a< �a<��a<�a<��a<�a<��a<%�a<��a<M�a<ʒa<j�a<ӓa<��a<�a<v�a<��a<x�a<��a<i�a<�a<\�a<�a<Z�a<ٙa<e�a<Ԛa<U�a<Лa<U�a<Μa<;�a<��a<�a<��a<ܞa<Q�a<��a<��a<C�a<��a<֠a<�a<s�a<��a<�a<B�a<w�a<Ţa<�a<W�a<��a<ãa<��a<&�a<}�a<k�a<��a<��a<�a<��a<�a<(�a<A�a<`�a<n�a<��a<��a<��a<إa<�a<�a<�a<7�a<+�a<M�a<f�a<7�a<\�a<9�a<Q�a</�a<+�a<�a<�a<�a<�a<�a<�a<̥a<ϥa<��a<ƥa<��a<��a<d�a<x�a<X�a<�a<�a<ͤa<Ĥa<x�a<[�a<�a<��a<Σa<��a<x�a<M�a<�a<��a<ɢa<��a<f�a<Q�a<��a<�a<��a<L�a<�a<Ǡa<��a<*�a<�a<��a<E�a<�a<��a<Y�a<��a<��a<[�a<�a<a<[�a<�a<��a<g�a<њa<j�a<��a<��a<�a<��a<�a<��a<'�a<��a<*�a<��a<;�a<ɔa<R�a<�a<r�a<�a<��a<��a<��a<�a<��a<�a<��a<�a<��a<�a<��a<%�a<��a<4�a<Ћa<X�a<��a<��a<K�a<�a<��a<&�a<ˈa<��a<�a<χa<`�a<�a<��a<b�a<�a<ʅa<��a<A�a<�a<؄a<��a<|�a<I�a<B�a<�a<��a<a<��a<��a<j�a<w�a<A�a<L�a<"�a<�a<�a<	�a<�a<�a<�a<)�a<3�a<[�a<k�a<��a<�  �  ��a<��a<�a<4�a<`�a<��a<��a<�a<
�a<9�a<��a<��a<��a<*�a<�a<��a<.�a<o�a<�a<0�a<��a<�a<�a<ۉa<P�a<��a<.�a<��a<�a<a�a<ӌa<K�a<a<�a<��a<4�a<��a<"�a<��a<<�a<��a<H�a<Вa<k�a<�a<l�a<�a<~�a<��a<��a<ۖa<l�a<ٗa<S�a<Ҙa<S�a<Йa<J�a<̚a<@�a<כa<<�a<՜a<@�a<��a<�a<��a<�a<W�a<��a<��a<F�a<��a<�a<.�a<^�a<͡a<�a<8�a<��a<ۢa<�a<K�a<��a<ѣa<
�a<"�a<_�a<x�a<��a<ʤa<�a<�a<�a<�a<A�a<E�a<d�a<|�a<��a<��a<ѥa<�a<�a<�a<*�a<9�a<F�a<H�a<T�a<`�a<=�a<B�a<;�a<;�a<.�a<�a<��a<�a<�a<ܥa<�a<ݥa<ťa<��a<��a<��a<��a<`�a<D�a<"�a<�a<ݤa<��a<p�a<T�a<�a<��a<��a<��a<\�a<K�a<�a<��a<��a<��a<u�a<F�a<�a<١a<��a<h�a<%�a<��a<��a<=�a<��a<��a<>�a<��a<a<F�a<�a<Ɲa<r�a<�a<��a<a�a<�a<��a<?�a<ךa<s�a<��a<��a<��a<��a<�a<��a<�a<��a<"�a<��a<3�a<��a<Y�a<͓a<x�a<��a<��a<�a<��a<�a<��a<�a<��a<�a<��a<$�a<��a<�a<Ča<C�a<Ƌa<z�a<�a<��a<>�a<ۉa<��a<<�a<ƈa<|�a<�a<Ƈa<k�a<�a<��a<l�a< �a<ʅa<q�a<8�a<��a<фa<��a<u�a<F�a<�a<�a<�a<уa<��a<��a<��a<{�a<F�a<>�a<.�a<*�a<�a<�a<��a<+�a<�a<#�a<L�a<j�a<|�a<��a<�  �  �a<�a<�a<9�a<^�a<��a<��a<�a<��a<5�a<k�a<��a<��a<�a<��a<��a<�a<e�a<؇a<%�a<��a<�a<g�a<�a<I�a<��a<$�a<��a<�a<m�a<ތa<9�a<��a<>�a<��a<2�a<��a<B�a<��a<@�a<͑a<`�a<�a<Z�a<�a<f�a<��a<s�a<�a<m�a<ɖa<e�a<ȗa<^�a<��a<D�a<ʙa<)�a<Ϛa<2�a<Λa<'�a<��a<+�a<��a<$�a<��a<��a<G�a<��a<�a<V�a<��a<ؠa<B�a<~�a<ʡa<�a<Z�a<��a<Ǣa<�a<\�a<��a<Σa<��a<3�a<U�a<��a<��a<��a<դa<֤a<�a<�a<2�a<�a<n�a<^�a<��a<��a<��a<ݥa<�a<�a<�a<@�a<@�a<I�a<Y�a<O�a<o�a<O�a<K�a<7�a<�a<:�a<�a<�a<��a<	�a<ڥa<ԥa<եa<��a<ͥa<��a<��a<e�a<B�a<0�a<�a<Ҥa<��a<k�a<=�a<�a<ݣa<��a<��a<9�a<6�a<��a<�a<��a<��a<e�a</�a<�a<ҡa<��a<^�a<�a<��a<��a<H�a<�a<��a<c�a<�a<��a<f�a<+�a<��a<v�a<$�a<՜a<��a<�a<��a<9�a<ښa<h�a<�a<|�a<�a<��a<��a<��a<�a<��a<�a<��a<6�a<��a<O�a<��a<c�a<�a<z�a<�a<��a<�a<��a<*�a<��a<"�a<��a<�a<��a<1�a<��a<L�a<�a<u�a<��a<��a<P�a<
�a<��a</�a<؈a<r�a<#�a<��a<V�a<�a<��a<]�a<�a<��a<J�a<B�a<߄a<��a<��a<`�a<B�a<�a<�a<݃a<؃a<��a<��a<��a<k�a<x�a<J�a<>�a<&�a<�a<3�a<�a<*�a<(�a<P�a<A�a<a�a<��a<��a<�  �  уa<�a<�a<N�a<_�a<�a<Äa<҄a<�a<4�a<Y�a<��a<ׅa<�a<j�a<��a<�a<Z�a<ˇa<6�a<��a<��a<��a<ωa<P�a<Êa<(�a<��a<�a<p�a<ތa<l�a<Ía<F�a<��a<+�a<��a<0�a<ʐa<K�a<ʑa<P�a<ؒa<l�a<�a<��a<�a<y�a<��a<b�a<�a<Z�a<��a<9�a<��a<7�a<��a<;�a<��a<+�a<��a<G�a<��a<;�a<��a<�a<��a<�a<U�a<��a<��a<S�a<��a<�a<:�a<��a<ȡa<�a<g�a<��a<��a<�a<_�a<��a<ƣa<�a<7�a<]�a<o�a<��a<��a<ݤa<�a<��a<��a< �a<;�a<T�a<c�a<~�a<��a<��a<եa< �a<�a<3�a</�a<=�a<b�a<R�a<]�a<Y�a<K�a<I�a<S�a<<�a<'�a<*�a<
�a<�a<��a<��a<��a<Хa<��a<��a<��a<��a<z�a<C�a<�a<	�a<äa<��a<j�a<,�a<��a<ԣa<��a<��a<T�a<'�a<�a<ܢa<��a<��a<X�a<P�a<��a<١a<��a<b�a<�a<۠a<��a<H�a<�a<��a<k�a<�a<��a<|�a<�a<۝a<��a<!�a<Ɯa<i�a<�a<��a<T�a<˚a<m�a<��a<q�a<�a<~�a<�a<o�a< �a<�a<�a<��a<�a<��a<@�a<ٓa<b�a<�a<��a<��a<��a<�a<��a<�a<��a<�a<��a<=�a<��a<I�a<��a<W�a<��a<z�a<3�a<��a<S�a<�a<��a<6�a<܈a<y�a<	�a<̇a<Q�a<	�a<��a<N�a<�a<��a<f�a<(�a<�a<��a<u�a<M�a<:�a<)�a<��a<��a<ǃa<��a<��a<��a<x�a<b�a<F�a<<�a<C�a<.�a< �a</�a< �a<=�a<C�a<[�a<��a<��a<��a<�  �  ƃa<�a<�a<9�a<s�a<r�a<��a<��a<��a<�a<q�a<��a<˅a<�a<9�a<��a<��a<t�a<̇a<�a<��a<݈a<��a<ĉa<e�a<��a<8�a<��a< �a<��a<یa<a�a<ʍa<G�a<Ύa<C�a<Џa<-�a<ސa<>�a<�a<x�a<ߒa<��a<ߓa<}�a<�a<i�a<ܕa<@�a<Ֆa<=�a<�a<0�a<��a<'�a<��a<8�a<��a<S�a<��a<3�a<��a<�a<��a<�a<��a<��a<s�a<��a<"�a<z�a<��a<�a<7�a<��a<�a<+�a<f�a<��a<��a<�a<��a<��a<�a<�a< �a<r�a<h�a<��a<��a<��a<פa<��a<�a<�a<:�a<'�a<_�a<v�a<��a<̥a<��a<�a<�a<"�a<!�a<O�a<Q�a<O�a<z�a<M�a<x�a<Z�a<E�a<N�a<�a<?�a<!�a<$�a<�a<�a<�a<ߥa<�a<��a<��a<��a<e�a<W�a<	�a<��a<��a<��a<S�a<D�a<�a<ȣa<��a<N�a<S�a<�a<�a<ݢa<��a<��a<=�a<G�a<�a<�a<��a<r�a<:�a<ڠa<àa<F�a<�a<��a<l�a<)�a<Ҟa<��a<�a<�a<t�a<>�a<�a<p�a<6�a<��a<P�a<Қa<^�a<ޙa<O�a<�a<a�a<�a<f�a<��a<o�a<�a<��a<	�a<ǔa<*�a<ēa<@�a<Ԓa<{�a<��a<��a<�a<��a<'�a<��a<F�a<��a<L�a<��a<P�a<،a<l�a<��a<~�a</�a<��a<��a<��a<��a<I�a<Ĉa<��a<�a<ća<5�a<�a<��a<H�a<�a<��a<f�a<��a<߄a<��a<}�a<p�a<�a<�a<Ճa<�a<��a<��a<��a<��a<��a<V�a<s�a<M�a<5�a<@�a<�a<C�a<6�a<P�a<:�a<i�a<w�a<��a<Ӄa<�  �  Ӄa<�a< �a<8�a<r�a<}�a<��a<݄a<�a<#�a<K�a<��a<��a<�a<_�a<��a<�a<Q�a<��a<'�a<��a<�a<j�a<؉a<W�a<��a<+�a<��a<�a<z�a<�a<[�a<�a<V�a<��a<;�a<a<Y�a<֐a<L�a<ёa<[�a<ےa<d�a<��a<p�a<��a<d�a<�a<m�a<�a<:�a<��a<&�a<��a<.�a<��a<)�a<��a<%�a<��a<?�a<��a<3�a<��a<%�a<��a<��a<O�a<��a<
�a<Y�a<��a<�a<`�a<��a<ءa<�a<r�a<¢a<�a<-�a<g�a<��a<��a<�a<.�a<a�a<{�a<��a<��a<ؤa<�a<�a<��a<�a<0�a<E�a<]�a<j�a<��a<��a<��a<��a<�a<"�a<&�a<S�a<J�a<`�a<O�a<Y�a<X�a<Y�a<L�a<V�a<K�a<+�a<�a<�a<�a<�a<�a<�a<ɥa<��a<��a<��a<d�a<V�a<�a<��a<ͤa<��a<Y�a<�a<�a<��a<��a<u�a<K�a<�a<�a<��a<��a<��a<h�a<1�a<�a<�a<��a<e�a<�a<�a<��a<W�a<�a<՟a<{�a<�a<ɞa<�a<B�a<�a<��a<(�a<Мa<l�a<�a<��a<D�a<�a<Y�a<�a<|�a<��a<^�a<�a<\�a<�a<v�a< �a<��a<�a<��a<$�a<ѓa<d�a<�a<s�a<�a<��a<�a<��a<�a<��a<%�a<��a<?�a<Ӎa<J�a<Ќa<Z�a< �a<��a<$�a<��a<[�a<��a<��a<3�a<ӈa<~�a<�a<��a<\�a<�a<��a<3�a<��a<��a<\�a<�a<݄a<��a<j�a<F�a<"�a<!�a<�a<�a<��a<ăa<��a<��a<j�a<b�a<S�a<L�a<<�a<H�a<C�a<0�a<,�a<=�a<_�a<x�a<|�a<��a<��a<�  �  ,�a<�a<j�a<f�a<��a<˅a<�a<,�a<4�a<��a<��a<Ԇa<&�a<R�a<��a<�a<N�a<��a<�a<d�a<��a<S�a<��a<�a<g�a<؋a<c�a<��a<N�a<�a<�a<��a<��a<m�a<��a<��a<ېa<x�a<ޑa<t�a<�a<r�a<	�a<m�a<�a<`�a<��a<l�a<��a<g�a<̗a<f�a<Θa<<�a<��a<)�a<��a<*�a<��a<-�a<��a<�a<��a<,�a<��a<
�a<S�a<ԟa<1�a<��a<��a<<�a<��a<�a<F�a<q�a<�a<�a<G�a<��a<ѣa<�a<,�a<��a<��a<�a<�a<*�a<r�a<w�a<��a<��a<ɥa<�a<��a<�a<�a<6�a<M�a<{�a<��a<��a<զa<Φa<�a<�a< �a<'�a<!�a<R�a<.�a<b�a<.�a<R�a<@�a<1�a<4�a<!�a<H�a<�a<��a<�a<ܦa<ܦa<��a<��a<x�a<��a<A�a<(�a<�a<�a<Υa<|�a<i�a<6�a<�a<פa<��a<h�a<8�a<"�a<�a<ڣa<��a<p�a<n�a<�a<�a<��a<z�a<]�a<�a<�a<g�a<N�a<��a<��a<[�a<�a<�a<g�a<2�a<a<~�a< �a<a<v�a<��a<��a<�a<ʛa<L�a<�a<h�a<ۙa<��a<��a<r�a< �a<x�a<�a<��a<�a<��a<X�a<Ŕa<j�a<�a<~�a<�a<��a<*�a<��a<G�a<̐a<A�a<��a<T�a<��a<c�a<�a<��a<�a<Ìa<P�a<��a<h�a<A�a<Ċa<m�a<��a<��a<Y�a<߈a<��a<2�a<ԇa<��a<3�a<�a<��a<[�a<�a<��a<��a<��a<��a<K�a<I�a<"�a<�a<�a<Ąa<لa<��a<��a<}�a<��a<��a<w�a<��a<y�a<��a<��a<��a<��a<��a<�a<քa<�  �  �a<&�a<d�a<z�a<��a<ƅa<�a<�a<I�a<r�a<��a<�a<�a<o�a<��a<�a<M�a<��a<�a<m�a<Ήa<1�a<��a<�a<��a<�a<\�a<��a<4�a<��a<�a<}�a<��a<w�a<ۏa<M�a<ݐa<d�a<ݑa<l�a<�a<p�a<�a<u�a<�a<��a< �a<r�a<�a<g�a<�a<P�a<ۘa<A�a<��a<G�a<ƚa<5�a<��a<<�a<��a<4�a<��a<�a<��a<�a<x�a<۟a<7�a<��a<�a<D�a<��a<ܡa<4�a<y�a<��a<��a<Q�a<��a<ɣa<�a<K�a<��a<��a<�a<�a<S�a<`�a<y�a<��a<��a<إa<�a<�a<�a<3�a<V�a<j�a<t�a<��a<��a<��a<�a<�a<�a<�a<=�a<>�a<U�a<;�a<J�a<E�a<J�a<6�a<3�a</�a<�a<��a<��a<�a<�a<Ԧa<צa<��a<��a<��a<��a<V�a<D�a<�a<ߥa<��a<��a<[�a<3�a<��a<Ϥa<��a<��a<S�a< �a<��a<ѣa<��a<}�a<M�a<�a<��a<բa<��a<V�a<�a<Сa<��a<M�a<�a<��a<e�a<�a<��a<i�a<�a<��a<w�a<�a<��a<^�a<��a<��a<:�a<͛a<Q�a<ݚa<g�a<��a<l�a<�a<w�a<�a<��a<"�a<��a<$�a<ŕa<D�a<�a<j�a<�a<��a<�a<��a<0�a<��a<3�a<��a<I�a<֏a<O�a<�a<l�a<�a<}�a<$�a<��a<G�a<��a<��a<(�a<��a<j�a<	�a<��a<F�a<�a<��a<5�a<�a<��a<?�a<�a<��a<z�a<<�a<��a<ǅa<��a<v�a<b�a<:�a<�a<
�a<�a<�a<܄a<��a<��a<��a<��a<z�a<y�a<{�a<q�a<`�a<�a<��a<��a<��a<�a<�a<�  �  �a<E�a<N�a<m�a<��a<��a<�a<�a<]�a<h�a<��a<�a<�a<a�a<��a<��a<E�a<��a<��a<i�a<߉a<1�a<��a<��a<��a<׋a<S�a<֌a<+�a<��a<�a<��a<�a<o�a<��a<^�a<��a<O�a<�a<h�a<�a<x�a<�a<��a<�a<}�a<�a<{�a<��a<`�a<��a<?�a<��a<C�a<��a<8�a<��a</�a<��a<=�a<��a<9�a<��a<"�a<��a<��a<y�a<ßa<F�a<��a<�a<B�a<��a<�a<!�a<��a<��a<�a<S�a<��a<֣a<�a<S�a<�a<ɤa<�a<�a<P�a<N�a<��a<��a<åa<إa<֥a<�a<�a<)�a<5�a<Z�a<g�a<��a<��a<��a<��a<�a<�a<�a<5�a<2�a<:�a<V�a<A�a<R�a<5�a<9�a<2�a<�a<7�a<�a<"�a<�a<�a<ܦa<��a<Ȧa<��a<��a<l�a<H�a<<�a<�a<��a<��a<��a<Q�a<0�a<	�a<äa<��a<i�a<J�a<�a<��a<��a<��a<��a<M�a<B�a<�a<Ӣa<y�a<M�a<#�a<ǡa<��a<6�a<��a<��a<]�a< �a<��a<��a<	�a<˞a<s�a<�a<ȝa<_�a<�a<��a<5�a<��a<[�a<�a<a�a<�a<\�a<	�a<y�a<��a<��a<�a<��a<%�a<ƕa<.�a<�a<d�a<��a<��a<	�a<��a<�a<��a<;�a<Őa<F�a<̏a<Z�a<Ҏa<��a<��a<��a<&�a<��a<T�a<�a<��a<!�a<֊a<j�a<��a<��a<5�a<�a<��a<>�a<�a<v�a<A�a<�a<��a<Z�a<,�a<�a<υa<��a<k�a<u�a<5�a<6�a<	�a<��a<Մa<��a<ńa<��a<��a<|�a<|�a<w�a<c�a<��a<p�a<��a<��a<��a<��a<ʄa< �a<�  �  �a<.�a<W�a<z�a<��a<��a<��a<'�a<M�a<z�a<��a<�a<8�a<o�a<��a<�a<d�a<��a<�a<e�a<ډa<E�a<��a<�a<w�a<�a<Z�a<��a<-�a<��a<�a<��a<�a<I�a<��a<\�a<ːa<U�a<�a<l�a<ܒa<n�a<�a<y�a<��a<z�a<��a<b�a<��a<n�a<ޗa<`�a<ʘa<R�a<ՙa<N�a<ƚa<E�a<��a<+�a<��a<%�a<��a<.�a<��a<�a<k�a<ϟa<:�a<��a<�a<0�a<��a<�a<%�a<a�a<��a< �a<,�a<��a<٣a<�a<3�a<�a<��a<�a<�a<9�a<_�a<��a<��a<ĥa<˥a<�a<��a<+�a<7�a<P�a<k�a<��a<��a<��a<Φa<�a< �a<�a<�a</�a<9�a<B�a<D�a<F�a<:�a<1�a<A�a<2�a<�a<�a<�a<��a<٦a<�a<�a<��a<��a<��a<��a<u�a<U�a<2�a<��a<�a<ɥa<��a<d�a<0�a<�a<�a<��a<��a<V�a<8�a<��a<֣a<��a<��a<a�a<'�a<�a<��a<��a<T�a<�a<ʡa<r�a<5�a<�a<��a<7�a<�a<��a<W�a<�a<ʞa<v�a<�a<��a<]�a<�a<��a<2�a<ɛa<B�a<�a<n�a<�a<}�a<��a<��a<�a<��a<"�a<��a<7�a<��a<P�a<Ӕa<m�a<	�a<{�a<�a<��a<$�a<��a<2�a<��a<4�a<Ϗa<Y�a<֎a<T�a<�a<��a<��a<��a<W�a<�a<p�a<"�a<a<j�a<�a<��a<E�a<�a<��a<?�a<ևa<��a<9�a<�a<��a<u�a<=�a<�a<Ӆa<��a<��a<_�a<G�a</�a<��a<�a<݄a<Ʉa<��a<��a<��a<x�a<��a<x�a<\�a<h�a<v�a<{�a<s�a<��a<Ȅa<Ʉa<�a<�  �  �a<�a<_�a<z�a<��a<مa<�a<'�a<<�a<��a<��a<��a<<�a<^�a<ˇa<��a<p�a<��a<(�a<s�a<ωa<C�a<��a<*�a<x�a<�a<Y�a<��a<9�a<��a<�a<d�a<�a<k�a<֏a<[�a<Аa<i�a<đa<b�a<��a<o�a<�a<c�a<�a<u�a<�a<s�a<�a<v�a<ۗa<y�a<Ԙa<f�a<əa<?�a<��a<9�a<қa<7�a<Ҝa<(�a<��a<"�a<��a<�a<f�a<�a<(�a<��a<�a<6�a<��a<¡a<5�a<m�a<��a<��a<F�a<��a<��a<�a<@�a<��a<��a<�a<#�a<8�a<~�a<z�a<��a<��a<֥a<�a<�a<6�a<.�a<]�a<X�a<��a<��a<��a<�a<զa<�a<	�a<)�a<:�a<9�a<O�a<(�a<I�a<D�a<<�a<(�a<�a</�a<�a<�a<�a<��a<ߦa<Ʀa<ͦa<��a<��a<o�a<|�a<U�a<:�a<!�a<ݥa<ɥa<��a<y�a<E�a<�a<�a<��a<��a<I�a<C�a< �a<�a<��a<~�a<_�a<�a<�a<��a<��a<S�a<�a<֡a<��a<G�a<נa<��a<Y�a<��a<��a<\�a<"�a<��a<l�a<�a<��a<Z�a<�a<��a<-�a<ܛa<S�a<�a<w�a<�a<��a<��a<��a<�a<��a<�a<��a<K�a<��a<l�a<֔a<u�a<��a<��a<.�a<��a<=�a<��a<(�a<a<;�a<Ϗa<6�a<�a<`�a<�a<�a<�a<��a<,�a<�a<|�a<,�a<��a<a�a<�a<��a<e�a<�a<��a<8�a<�a<��a<@�a<�a<��a<��a<*�a<�a<��a<��a<��a<R�a<N�a< �a<�a<��a<܄a<քa<��a<��a<��a<��a<l�a<e�a<|�a<]�a<r�a<l�a<��a<��a<��a<ׄa<�a<�  �  ��a<:�a<U�a<q�a<��a<Ѕa<��a<$�a<f�a<��a<��a<�a<@�a<y�a<ʇa<�a<n�a<��a<�a<��a<�a<?�a<��a<�a<|�a<܋a<T�a<ǌa<"�a<��a< �a<m�a<��a<b�a<ŏa<>�a<Ԑa<F�a<Αa<V�a<Ԓa<g�a<�a<{�a<��a<t�a<�a<��a<�a<w�a<�a<g�a<�a<b�a<��a<U�a<њa<R�a<͛a<F�a<��a<P�a<��a<�a<��a<��a<k�a<՟a<8�a<��a<�a<-�a<��a<ϡa<�a<l�a<��a<�a<@�a<u�a<��a< �a<8�a<u�a<��a<�a<�a<?�a<\�a<��a<��a<ӥa<��a<��a<�a<2�a<I�a<a�a<s�a<��a<��a<æa<֦a<�a<�a<�a<2�a<*�a<1�a<@�a<K�a<:�a<>�a<'�a<(�a<�a<�a<�a<��a<�a<�a<Ԧa<Ȧa<��a<��a<��a<��a<s�a<L�a<0�a<�a<��a<ƥa<��a<v�a<G�a<�a<�a<��a<��a<d�a<B�a<�a<�a<ƣa<��a<[�a<=�a<��a<¢a<~�a<M�a<�a<��a<x�a</�a<�a<��a<P�a<�a<��a<`�a< �a<��a<`�a<�a<��a<Y�a<�a<��a<,�a<��a<r�a<��a<w�a<�a<��a<�a<��a<"�a<��a<.�a<��a<F�a<ϕa<V�a<��a<{�a<��a<��a<
�a<��a<*�a<��a<3�a<��a<1�a<��a<B�a<Ŏa<_�a<֍a<d�a<�a<��a<;�a<ۋa<u�a<�a<Êa<c�a<��a<��a<B�a<�a<��a<N�a< �a<��a<K�a<�a<ņa<��a<E�a<�a<߅a<��a<��a<��a<K�a<-�a<�a<�a<Ԅa<Ǆa<��a<��a<��a<n�a<k�a<_�a<[�a<`�a<_�a<k�a<��a<��a<��a<��a<�a<�  �  �a<:�a<>�a<��a<��a<��a<�a<�a<n�a<�a<цa<��a<C�a<��a<��a<,�a<g�a<ψa<"�a<�a<�a<0�a<a<��a<��a<ߋa<J�a<��a<�a<��a<�a<r�a<ˎa<R�a<Ǐa</�a<͐a</�a<Ցa<=�a<ܒa<^�a<ϓa<~�a<ٔa<��a<�a<��a<��a<j�a<�a<`�a<��a<X�a<�a<[�a<њa<e�a<��a<_�a<��a<Q�a<��a<!�a<��a<�a<��a<��a<:�a<v�a<Ԡa<8�a<h�a<աa<��a<e�a<��a<�a<7�a<^�a<��a<ߣa<D�a<Y�a<��a<�a<�a<]�a<N�a<��a<��a<ԥa<�a<��a</�a<)�a<^�a<X�a<��a<��a<��a<Ԧa<̦a<�a<�a<#�a<!�a<3�a<Q�a<&�a<O�a<�a<?�a< �a<�a<�a<��a<�a<ݦa<�a<զa<ɦa<Ȧa<��a<��a<{�a<��a<\�a<f�a<D�a<�a<�a<��a<��a<i�a<W�a<�a<��a<Фa<��a<~�a<;�a< �a<�a<��a<��a<K�a<F�a<�a<ޢa<��a<D�a<�a<��a<��a<�a<�a<~�a<A�a<�a<��a<Y�a<�a<��a<H�a<�a<��a<=�a<�a<{�a<O�a<��a<j�a<�a<j�a<�a<}�a<'�a<��a<5�a<��a<.�a<ϖa<9�a<�a<S�a<��a<r�a<��a<��a< �a<��a<
�a<��a<�a<��a<=�a<��a<H�a<��a<W�a<ʍa<f�a<	�a<��a<>�a<��a<��a<��a<��a<d�a<�a<Ɖa<5�a<	�a<��a<O�a<��a<��a<i�a<�a<ۆa<}�a<X�a< �a<�a<˅a<��a<��a<4�a<9�a<�a<��a<�a<��a<��a<z�a<��a<g�a<b�a<Z�a<K�a<_�a<G�a<k�a<o�a<��a<��a<��a<�a<�  �  ��a<*�a<M�a<r�a<��a<օa<�a<*�a<e�a<��a<φa<�a<U�a<��a<ׇa</�a<x�a<шa<0�a<��a<�a<M�a<��a<�a<u�a<ۋa<[�a<��a<�a<��a<�a<^�a<ˎa<G�a<��a<7�a<��a<9�a<��a<;�a<ޒa<^�a<ۓa<�a<�a<z�a<��a<��a<	�a<��a<��a<��a<��a<o�a<��a<\�a<ٚa<m�a<ڛa<Z�a<՜a<F�a<��a<6�a<��a<
�a<l�a<��a<>�a<y�a<٠a<7�a<j�a<��a<�a<Q�a<��a<٢a<&�a<e�a<��a<�a<C�a<i�a<��a<�a<�a<9�a<q�a<��a<��a<ۥa<�a<�a<(�a<?�a<e�a<j�a<��a<��a<��a<Ϧa<�a<��a<
�a<-�a</�a<)�a<6�a<5�a<C�a<.�a<8�a<)�a<�a<��a<�a<�a<�a<զa<֦a<��a<��a<��a<��a<��a<��a<k�a<M�a</�a<�a<�a<̥a<��a<}�a<U�a<*�a<�a<Ϥa<��a<��a<L�a<"�a<��a<��a<��a<h�a<@�a<�a<��a<}�a<T�a<��a<��a<��a<�a<Рa<}�a<6�a<ݟa<��a<D�a<�a<��a<F�a<�a<��a<I�a<�a<��a<2�a<ƛa<g�a<��a<��a<�a<��a<#�a<��a<=�a<��a<5�a<זa<S�a<�a<p�a<��a<��a<�a<��a<�a<��a<�a<��a<�a<��a<;�a<��a<.�a<��a<D�a<͍a<\�a<��a<��a<&�a<��a<�a<�a<��a<o�a<�a<��a<W�a<�a<��a<V�a<��a<��a<c�a<�a<�a<��a<V�a<2�a<��a<ƅa<��a<x�a<Q�a<D�a<�a<�a<لa<��a<��a<��a<��a<p�a<V�a<B�a<Q�a<F�a<P�a<T�a<p�a<q�a<��a<��a<�a<�  �  ��a<�a<\�a<y�a<��a<݅a<�a<B�a<l�a<��a<̆a<�a<h�a<��a<�a<*�a<��a<҈a<1�a<��a<��a<Z�a<��a<*�a<{�a<��a<J�a<��a<�a<i�a<��a<S�a<Ύa<=�a<��a<0�a<��a<>�a<��a<T�a<��a<L�a<ݓa<Z�a<
�a<s�a<�a<��a<�a<��a<�a<��a<�a<��a< �a<z�a<��a<p�a<��a<M�a<�a<O�a<Нa<%�a<��a<�a<e�a<�a<�a<|�a<Рa<�a<��a<��a<�a<5�a<��a<��a<�a<j�a<��a<��a<�a<l�a<��a<֤a<#�a<<�a<��a<��a<��a<�a<��a<�a<!�a<b�a<`�a<��a<��a<��a<̦a<ʦa< �a<�a<$�a<	�a<5�a<:�a<6�a<N�a<$�a<2�a<�a<�a<�a<��a<�a<Ҧa<�a<��a<Ҧa<��a<��a<��a<��a<��a<i�a<y�a<U�a<:�a<%�a<�a<�a<��a<��a<R�a<7�a<�a<Ԥa<��a<{�a<o�a<#�a<��a<գa<��a<u�a<!�a<�a<¢a<��a<C�a<�a<��a<Q�a<(�a<Ša<��a<,�a<ßa<��a<'�a<��a<��a<^�a<�a<��a<K�a<�a<��a<+�a<ޛa<a�a<�a<��a<�a<��a<�a<��a<B�a<ɗa<U�a<ږa<r�a<֕a<��a<��a<��a< �a<��a<1�a<��a<:�a<��a<!�a<��a<�a<��a<�a<��a<(�a<��a<E�a<�a<��a<�a<ҋa<P�a<�a<��a<R�a<�a<��a<g�a<�a<��a<^�a<�a<��a<[�a<;�a<܆a<��a<b�a<=�a<�a<��a<��a<��a<l�a< �a<!�a<��a<لa<Ԅa<��a<��a<g�a<c�a<c�a<>�a<P�a<+�a<T�a<:�a<m�a<p�a<��a<��a<��a<�  �  ��a<"�a<:�a<s�a<��a<؅a<�a<:�a<a�a<��a<�a<�a<A�a<��a<�a<2�a<�a<�a<F�a<��a<��a<V�a<��a<�a<|�a<�a</�a<��a<�a<u�a<�a<C�a<��a<C�a<��a<(�a<��a<1�a<��a<5�a<��a<P�a<�a<_�a<�a<u�a<��a<��a<	�a<��a<��a<��a<�a<��a<�a<|�a<��a<b�a<�a<q�a<�a<E�a<˝a<4�a<��a<�a<j�a<˟a<�a<��a<ˠa<�a<d�a<��a<��a<A�a<��a<Ӣa<�a<W�a<��a<�a<�a<b�a<��a<��a<�a<>�a<l�a<��a<��a<�a<��a<'�a<A�a<L�a<`�a<��a<��a<��a<˦a<�a<�a<��a<�a<$�a<6�a<0�a<3�a<*�a<2�a<4�a<%�a<�a<�a<�a<��a<�a<ئa<ʦa<̦a<��a<��a<��a<��a<��a<}�a<X�a<N�a<7�a<!�a<��a<ܥa<��a<��a<w�a<>�a<�a<�a<��a<��a<S�a<;�a<�a<ˣa<��a<r�a<<�a<�a<¢a<��a<)�a< �a<��a<]�a<�a<��a<q�a<1�a<ןa<��a<1�a<�a<��a<@�a<�a<��a<R�a<�a<��a<-�a<˛a<m�a<��a<��a<�a<��a<<�a<��a<-�a<̗a<S�a<̖a<d�a<��a<~�a<�a<��a<�a<��a<�a<��a< �a<��a<+�a<��a<�a<��a<�a<��a<4�a<��a<V�a<�a<}�a<�a<��a<V�a<�a<��a<=�a< �a<��a<R�a<�a<��a<[�a< �a<Ǉa<|�a<%�a<܆a<��a<n�a<�a<�a<�a<��a<s�a<`�a<;�a<!�a<��a<ׄa<��a<��a<��a<u�a<R�a<H�a<8�a<E�a<9�a<A�a<I�a<f�a<l�a<��a<��a<Єa<�  �  �a<2�a<;�a<��a<��a<υa<�a<4�a<~�a<��a<�a<�a<\�a<Ƈa<�a<\�a<��a<�a<@�a<��a<�a<S�a<ˊa<�a<x�a<�a<D�a<��a<�a<��a<ɍa<R�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<L�a<ԓa<z�a<ܔa<��a<�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<��a<��a<�a<q�a<�a<]�a<Нa<@�a<��a<��a<|�a<��a<2�a<w�a<Ġa<�a<C�a<��a<�a<0�a<n�a<��a<��a<J�a<��a<��a<4�a<T�a<��a<ڤa<	�a<?�a<d�a<��a<��a<�a<��a<$�a<C�a<H�a<��a<��a<��a<��a<Ʀa<�a<�a<�a<�a<:�a<,�a<$�a<E�a<$�a<J�a<�a<-�a<�a<�a<��a<ئa<զa<��a<��a<��a<��a<��a<��a<��a<x�a<��a<X�a<[�a<*�a<�a<�a<֥a<ƥa<��a<k�a<:�a<�a<�a<��a<��a<U�a<;�a<
�a<ѣa<��a<n�a<N�a<��a<��a<��a<=�a<�a<��a<u�a<��a<Ša<i�a<�a<ğa<f�a<#�a<Ҟa<��a<$�a<�a<��a<B�a<�a<}�a<D�a<��a<p�a<�a<��a<&�a<��a<:�a<��a<T�a<ؗa<[�a<��a<a�a<��a<|�a<
�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<"�a<}�a<#�a<��a<"�a<��a<@�a<Ќa<p�a<"�a<��a<p�a<��a<��a<V�a<��a<��a<J�a<�a<��a<h�a<	�a<Ňa<}�a<!�a<
�a<��a<��a<<�a< �a<�a<��a<��a<[�a<Q�a<�a<�a<�a<��a<��a<y�a<|�a<R�a<7�a<=�a<%�a<.�a<$�a<=�a<A�a<n�a<�a<��a<܄a<�  �  �a<�a<F�a<��a<��a<�a<��a<=�a<s�a<��a<܆a<'�a<q�a<��a<هa<=�a<��a<�a<?�a<��a<��a<[�a<��a</�a<��a<�a<D�a<��a<	�a<z�a<Ӎa<N�a<��a<'�a<��a<+�a<��a<�a<��a<,�a<��a<G�a<͓a<Y�a<�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<
�a<u�a<�a<{�a<��a<f�a<�a<\�a<Νa<2�a<��a<�a<z�a<˟a<�a<o�a<Ƞa<�a<Y�a<��a<�a<6�a<��a<ˢa<�a<F�a<��a<Σa<%�a<Z�a<��a<Ԥa<�a<E�a<�a<��a<��a<�a<
�a<&�a<9�a<^�a<p�a<t�a<��a<Ŧa<Ӧa<�a<�a<�a<�a<�a<7�a<6�a<H�a<3�a<%�a<�a<�a<�a< �a<�a<�a<ަa<ڦa<ʦa<��a<��a<��a<��a<��a<|�a<o�a<c�a<b�a<9�a<*�a<�a<ߥa<��a<��a<b�a<E�a<#�a<�a<��a<��a<l�a<8�a<	�a<�a<��a<w�a<4�a<�a<ɢa<��a<=�a<�a<��a<b�a<�a<��a<b�a<�a<՟a<��a<,�a<՞a<��a<7�a<�a<��a<;�a<�a<��a<D�a<ӛa<m�a<�a<��a<�a<��a</�a<Řa<M�a<ŗa<K�a<�a<u�a<�a<��a<
�a<��a<�a<��a<#�a<��a<!�a<��a<�a<��a<�a<��a<#�a<��a<)�a<a<O�a<ڌa<l�a<�a<��a<a�a<��a<��a<P�a<�a<��a<e�a<��a<��a<^�a<�a<Ǉa<s�a<7�a<�a<��a<k�a<I�a<�a<ׅa<��a<��a<e�a<2�a<"�a<��a<�a<��a<��a<z�a<i�a<X�a<D�a<9�a</�a<7�a<C�a<I�a<M�a<e�a<��a<��a<Ȅa<�  �  �a<�a<M�a<f�a<��a<�a<��a<V�a<T�a<��a<�a<'�a<j�a<��a<(�a<B�a<��a<�a<J�a<��a<�a<t�a<��a<-�a<e�a<ۋa<D�a<��a<�a<c�a<�a<G�a<��a<-�a<��a<�a<��a<�a<��a<;�a<��a<G�a<�a<X�a<��a<d�a<��a<��a<�a<��a<��a<��a<�a<��a<��a<��a<�a<r�a<
�a<l�a<��a<N�a<ݝa<B�a<��a<�a<T�a<՟a<�a<��a<Ǡa<�a<l�a<��a<�a<&�a<n�a<��a<�a<@�a<��a<�a<�a<\�a<��a<Фa<�a<%�a<{�a<��a<֥a<ߥa<�a</�a<9�a<p�a<p�a<��a<��a<��a<٦a<�a<	�a<�a<6�a<�a<A�a<%�a<$�a<A�a<%�a<@�a<
�a<�a<�a<�a<�a<¦a<��a<��a<��a<��a<��a<��a<{�a<��a<q�a<k�a<B�a<&�a<2�a<�a<��a<��a<��a<g�a<E�a<�a<�a<�a<��a<t�a<6�a<�a<�a<��a<��a<&�a<�a<��a<}�a<=�a<��a<��a<K�a<�a<��a<\�a<�a<��a<i�a<�a<Оa<��a<E�a<ݝa<��a<Y�a<�a<��a<�a<Ûa<m�a<��a<��a<�a<��a<8�a<јa<B�a<�a<{�a<ܖa<��a<��a<��a<��a<��a<�a<��a<�a<��a<*�a<��a<-�a<��a<�a<��a<�a<��a<�a<��a<2�a<ڌa<f�a<�a<Ëa<C�a<��a<��a<L�a<��a<��a<b�a<�a<ƈa<Z�a<�a<Їa<s�a<I�a<�a<ކa<��a<A�a<�a<ۅa<��a<h�a<~�a<3�a<-�a<�a<Ȅa<Ȅa<��a<��a<Z�a<S�a<L�a<,�a<2�a<�a<$�a<,�a<T�a<X�a<��a<��a<��a<�  �  �a<�a<F�a<��a<��a<�a<��a<=�a<s�a<��a<܆a<'�a<q�a<��a<هa<=�a<��a<�a<?�a<��a<��a<[�a<��a</�a<��a<�a<D�a<��a<	�a<z�a<Ӎa<N�a<��a<'�a<��a<+�a<��a<�a<��a<,�a<��a<G�a<͓a<Y�a<�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<
�a<u�a<�a<{�a<��a<f�a<�a<\�a<Νa<2�a<��a<�a<z�a<˟a<�a<o�a<Ƞa<�a<Y�a<��a<�a<6�a<��a<ˢa<�a<F�a<��a<Σa<%�a<Z�a<��a<Ԥa<�a<E�a<�a<��a<��a<�a<
�a<&�a<9�a<^�a<p�a<t�a<��a<Ŧa<Ӧa<�a<�a<�a<�a<�a<7�a<6�a<H�a<3�a<%�a<�a<�a<�a< �a<�a<�a<ަa<ڦa<ʦa<��a<��a<��a<��a<��a<|�a<o�a<c�a<b�a<9�a<*�a<�a<ߥa<��a<��a<b�a<E�a<#�a<�a<��a<��a<l�a<8�a<	�a<�a<��a<w�a<4�a<�a<ɢa<��a<=�a<�a<��a<b�a<�a<��a<b�a<�a<՟a<��a<,�a<՞a<��a<7�a<�a<��a<;�a<�a<��a<D�a<ӛa<m�a<�a<��a<�a<��a</�a<Řa<M�a<ŗa<K�a<�a<u�a<�a<��a<
�a<��a<�a<��a<#�a<��a<!�a<��a<�a<��a<�a<��a<#�a<��a<)�a<a<O�a<ڌa<l�a<�a<��a<a�a<��a<��a<P�a<�a<��a<e�a<��a<��a<^�a<�a<Ǉa<s�a<7�a<�a<��a<k�a<I�a<�a<ׅa<��a<��a<e�a<2�a<"�a<��a<�a<��a<��a<z�a<i�a<X�a<D�a<9�a</�a<7�a<C�a<I�a<M�a<e�a<��a<��a<Ȅa<�  �  �a<2�a<;�a<��a<��a<υa<�a<4�a<~�a<��a<�a<�a<\�a<Ƈa<�a<\�a<��a<�a<@�a<��a<�a<S�a<ˊa<�a<x�a<�a<D�a<��a<�a<��a<ɍa<R�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<L�a<ԓa<z�a<ܔa<��a<�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<��a<��a<�a<q�a<�a<]�a<Нa<@�a<��a<��a<|�a<��a<2�a<w�a<Ġa<�a<C�a<��a<�a<0�a<n�a<��a<��a<J�a<��a<��a<4�a<T�a<��a<ڤa<	�a<?�a<d�a<��a<��a<�a<��a<$�a<C�a<H�a<��a<��a<��a<��a<Ʀa<�a<�a<�a<�a<:�a<,�a<$�a<E�a<$�a<J�a<�a<-�a<�a<�a<��a<ئa<զa<��a<��a<��a<��a<��a<��a<��a<x�a<��a<X�a<[�a<*�a<�a<�a<֥a<ƥa<��a<k�a<:�a<�a<�a<��a<��a<U�a<;�a<
�a<ѣa<��a<n�a<N�a<��a<��a<��a<=�a<�a<��a<u�a<��a<Ša<i�a<�a<ğa<f�a<#�a<Ҟa<��a<$�a<�a<��a<B�a<�a<}�a<D�a<��a<p�a<�a<��a<&�a<��a<:�a<��a<T�a<ؗa<[�a<��a<a�a<��a<|�a<
�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<"�a<}�a<#�a<��a<"�a<��a<@�a<Ќa<p�a<"�a<��a<p�a<��a<��a<V�a<��a<��a<J�a<�a<��a<h�a<	�a<Ňa<}�a<!�a<
�a<��a<��a<<�a< �a<�a<��a<��a<[�a<Q�a<�a<�a<�a<��a<��a<y�a<|�a<R�a<7�a<=�a<%�a<.�a<$�a<=�a<A�a<n�a<�a<��a<܄a<�  �  ��a<"�a<:�a<s�a<��a<؅a<�a<:�a<a�a<��a<�a<�a<A�a<��a<�a<2�a<�a<�a<F�a<��a<��a<V�a<��a<�a<|�a<�a</�a<��a<�a<u�a<�a<C�a<��a<C�a<��a<(�a<��a<1�a<��a<5�a<��a<P�a<�a<_�a<�a<u�a<��a<��a<	�a<��a<��a<��a<�a<��a<�a<|�a<��a<b�a<�a<q�a<�a<E�a<˝a<4�a<��a<�a<j�a<˟a<�a<��a<ˠa<�a<d�a<��a<��a<A�a<��a<Ӣa<�a<W�a<��a<�a<�a<b�a<��a<��a<�a<>�a<l�a<��a<��a<�a<��a<'�a<A�a<L�a<`�a<��a<��a<��a<˦a<�a<�a<��a<�a<$�a<6�a<0�a<3�a<*�a<2�a<4�a<%�a<�a<�a<�a<��a<�a<ئa<ʦa<̦a<��a<��a<��a<��a<��a<}�a<X�a<N�a<7�a<!�a<��a<ܥa<��a<��a<w�a<>�a<�a<�a<��a<��a<S�a<;�a<�a<ˣa<��a<r�a<<�a<�a<¢a<��a<)�a< �a<��a<]�a<�a<��a<q�a<1�a<ןa<��a<1�a<�a<��a<@�a<�a<��a<R�a<�a<��a<-�a<˛a<m�a<��a<��a<�a<��a<<�a<��a<-�a<̗a<S�a<̖a<d�a<��a<~�a<�a<��a<�a<��a<�a<��a< �a<��a<+�a<��a<�a<��a<�a<��a<4�a<��a<V�a<�a<}�a<�a<��a<V�a<�a<��a<=�a< �a<��a<R�a<�a<��a<[�a< �a<Ǉa<|�a<%�a<܆a<��a<n�a<�a<�a<�a<��a<s�a<`�a<;�a<!�a<��a<ׄa<��a<��a<��a<u�a<R�a<H�a<8�a<E�a<9�a<A�a<I�a<f�a<l�a<��a<��a<Єa<�  �  ��a<�a<\�a<y�a<��a<݅a<�a<B�a<l�a<��a<̆a<�a<h�a<��a<�a<*�a<��a<҈a<1�a<��a<��a<Z�a<��a<*�a<{�a<��a<J�a<��a<�a<i�a<��a<S�a<Ύa<=�a<��a<0�a<��a<>�a<��a<T�a<��a<L�a<ݓa<Z�a<
�a<s�a<�a<��a<�a<��a<�a<��a<�a<��a< �a<z�a<��a<p�a<��a<M�a<�a<O�a<Нa<%�a<��a<�a<e�a<�a<�a<|�a<Рa<�a<��a<��a<�a<5�a<��a<��a<�a<j�a<��a<��a<�a<l�a<��a<֤a<#�a<<�a<��a<��a<��a<�a<��a<�a<!�a<b�a<`�a<��a<��a<��a<̦a<ʦa< �a<�a<$�a<	�a<5�a<:�a<6�a<N�a<$�a<2�a<�a<�a<�a<��a<�a<Ҧa<�a<��a<Ҧa<��a<��a<��a<��a<��a<i�a<y�a<U�a<:�a<%�a<�a<�a<��a<��a<R�a<7�a<�a<Ԥa<��a<{�a<o�a<#�a<��a<գa<��a<u�a<!�a<�a<¢a<��a<C�a<�a<��a<Q�a<(�a<Ša<��a<,�a<ßa<��a<'�a<��a<��a<^�a<�a<��a<K�a<�a<��a<+�a<ޛa<a�a<�a<��a<�a<��a<�a<��a<B�a<ɗa<U�a<ږa<r�a<֕a<��a<��a<��a< �a<��a<1�a<��a<:�a<��a<!�a<��a<�a<��a<�a<��a<(�a<��a<E�a<�a<��a<�a<ҋa<P�a<�a<��a<R�a<�a<��a<g�a<�a<��a<^�a<�a<��a<[�a<;�a<܆a<��a<b�a<=�a<�a<��a<��a<��a<l�a< �a<!�a<��a<لa<Ԅa<��a<��a<g�a<c�a<c�a<>�a<P�a<+�a<T�a<:�a<m�a<p�a<��a<��a<��a<�  �  ��a<*�a<M�a<r�a<��a<օa<�a<*�a<e�a<��a<φa<�a<U�a<��a<ׇa</�a<x�a<шa<0�a<��a<�a<M�a<��a<�a<u�a<ۋa<[�a<��a<�a<��a<�a<^�a<ˎa<G�a<��a<7�a<��a<9�a<��a<;�a<ޒa<^�a<ۓa<�a<�a<z�a<��a<��a<	�a<��a<��a<��a<��a<o�a<��a<\�a<ٚa<m�a<ڛa<Z�a<՜a<F�a<��a<6�a<��a<
�a<l�a<��a<>�a<y�a<٠a<7�a<j�a<��a<�a<Q�a<��a<٢a<&�a<e�a<��a<�a<C�a<i�a<��a<�a<�a<9�a<q�a<��a<��a<ۥa<�a<�a<(�a<?�a<e�a<j�a<��a<��a<��a<Ϧa<�a<��a<
�a<-�a</�a<)�a<6�a<5�a<C�a<.�a<8�a<)�a<�a<��a<�a<�a<�a<զa<֦a<��a<��a<��a<��a<��a<��a<k�a<M�a</�a<�a<�a<̥a<��a<}�a<U�a<*�a<�a<Ϥa<��a<��a<L�a<"�a<��a<��a<��a<h�a<@�a<�a<��a<}�a<T�a<��a<��a<��a<�a<Рa<}�a<6�a<ݟa<��a<D�a<�a<��a<F�a<�a<��a<I�a<�a<��a<2�a<ƛa<g�a<��a<��a<�a<��a<#�a<��a<=�a<��a<5�a<זa<S�a<�a<p�a<��a<��a<�a<��a<�a<��a<�a<��a<�a<��a<;�a<��a<.�a<��a<D�a<͍a<\�a<��a<��a<&�a<��a<�a<�a<��a<o�a<�a<��a<W�a<�a<��a<V�a<��a<��a<c�a<�a<�a<��a<V�a<2�a<��a<ƅa<��a<x�a<Q�a<D�a<�a<�a<لa<��a<��a<��a<��a<p�a<V�a<B�a<Q�a<F�a<P�a<T�a<p�a<q�a<��a<��a<�a<�  �  �a<:�a<>�a<��a<��a<��a<�a<�a<n�a<�a<цa<��a<C�a<��a<��a<,�a<g�a<ψa<"�a<�a<�a<0�a<a<��a<��a<ߋa<J�a<��a<�a<��a<�a<r�a<ˎa<R�a<Ǐa</�a<͐a</�a<Ցa<=�a<ܒa<^�a<ϓa<~�a<ٔa<��a<�a<��a<��a<j�a<�a<`�a<��a<X�a<�a<[�a<њa<e�a<��a<_�a<��a<Q�a<��a<!�a<��a<�a<��a<��a<:�a<v�a<Ԡa<8�a<h�a<աa<��a<e�a<��a<�a<7�a<^�a<��a<ߣa<D�a<Y�a<��a<�a<�a<]�a<N�a<��a<��a<ԥa<�a<��a</�a<)�a<^�a<X�a<��a<��a<��a<Ԧa<̦a<�a<�a<#�a<!�a<3�a<Q�a<&�a<O�a<�a<?�a< �a<�a<�a<��a<�a<ݦa<�a<զa<ɦa<Ȧa<��a<��a<{�a<��a<\�a<f�a<D�a<�a<�a<��a<��a<i�a<W�a<�a<��a<Фa<��a<~�a<;�a< �a<�a<��a<��a<K�a<F�a<�a<ޢa<��a<D�a<�a<��a<��a<�a<�a<~�a<A�a<�a<��a<Y�a<�a<��a<H�a<�a<��a<=�a<�a<{�a<O�a<��a<j�a<�a<j�a<�a<}�a<'�a<��a<5�a<��a<.�a<ϖa<9�a<�a<S�a<��a<r�a<��a<��a< �a<��a<
�a<��a<�a<��a<=�a<��a<H�a<��a<W�a<ʍa<f�a<	�a<��a<>�a<��a<��a<��a<��a<d�a<�a<Ɖa<5�a<	�a<��a<O�a<��a<��a<i�a<�a<ۆa<}�a<X�a< �a<�a<˅a<��a<��a<4�a<9�a<�a<��a<�a<��a<��a<z�a<��a<g�a<b�a<Z�a<K�a<_�a<G�a<k�a<o�a<��a<��a<��a<�a<�  �  ��a<:�a<U�a<q�a<��a<Ѕa<��a<$�a<f�a<��a<��a<�a<@�a<y�a<ʇa<�a<n�a<��a<�a<��a<�a<?�a<��a<�a<|�a<܋a<T�a<ǌa<"�a<��a< �a<m�a<��a<b�a<ŏa<>�a<Ԑa<F�a<Αa<V�a<Ԓa<g�a<�a<{�a<��a<t�a<�a<��a<�a<w�a<�a<g�a<�a<b�a<��a<U�a<њa<R�a<͛a<F�a<��a<P�a<��a<�a<��a<��a<k�a<՟a<8�a<��a<�a<-�a<��a<ϡa<�a<l�a<��a<�a<@�a<u�a<��a< �a<8�a<u�a<��a<�a<�a<?�a<\�a<��a<��a<ӥa<��a<��a<�a<2�a<I�a<a�a<s�a<��a<��a<æa<֦a<�a<�a<�a<2�a<*�a<1�a<@�a<K�a<:�a<>�a<'�a<(�a<�a<�a<�a<��a<�a<�a<Ԧa<Ȧa<��a<��a<��a<��a<s�a<L�a<0�a<�a<��a<ƥa<��a<v�a<G�a<�a<�a<��a<��a<d�a<B�a<�a<�a<ƣa<��a<[�a<=�a<��a<¢a<~�a<M�a<�a<��a<x�a</�a<�a<��a<P�a<�a<��a<`�a< �a<��a<`�a<�a<��a<Y�a<�a<��a<,�a<��a<r�a<��a<w�a<�a<��a<�a<��a<"�a<��a<.�a<��a<F�a<ϕa<V�a<��a<{�a<��a<��a<
�a<��a<*�a<��a<3�a<��a<1�a<��a<B�a<Ŏa<_�a<֍a<d�a<�a<��a<;�a<ۋa<u�a<�a<Êa<c�a<��a<��a<B�a<�a<��a<N�a< �a<��a<K�a<�a<ņa<��a<E�a<�a<߅a<��a<��a<��a<K�a<-�a<�a<�a<Ԅa<Ǆa<��a<��a<��a<n�a<k�a<_�a<[�a<`�a<_�a<k�a<��a<��a<��a<��a<�a<�  �  �a<�a<_�a<z�a<��a<مa<�a<'�a<<�a<��a<��a<��a<<�a<^�a<ˇa<��a<p�a<��a<(�a<s�a<ωa<C�a<��a<*�a<x�a<�a<Y�a<��a<9�a<��a<�a<d�a<�a<k�a<֏a<[�a<Аa<i�a<đa<b�a<��a<o�a<�a<c�a<�a<u�a<�a<s�a<�a<v�a<ۗa<y�a<Ԙa<f�a<əa<?�a<��a<9�a<қa<7�a<Ҝa<(�a<��a<"�a<��a<�a<f�a<�a<(�a<��a<�a<6�a<��a<¡a<5�a<m�a<��a<��a<F�a<��a<��a<�a<@�a<��a<��a<�a<#�a<8�a<~�a<z�a<��a<��a<֥a<�a<�a<6�a<.�a<]�a<X�a<��a<��a<��a<�a<զa<�a<	�a<)�a<:�a<9�a<O�a<(�a<I�a<D�a<<�a<(�a<�a</�a<�a<�a<�a<��a<ߦa<Ʀa<ͦa<��a<��a<o�a<|�a<U�a<:�a<!�a<ݥa<ɥa<��a<y�a<E�a<�a<�a<��a<��a<I�a<C�a< �a<�a<��a<~�a<_�a<�a<�a<��a<��a<S�a<�a<֡a<��a<G�a<נa<��a<Y�a<��a<��a<\�a<"�a<��a<l�a<�a<��a<Z�a<�a<��a<-�a<ܛa<S�a<�a<w�a<�a<��a<��a<��a<�a<��a<�a<��a<K�a<��a<l�a<֔a<u�a<��a<��a<.�a<��a<=�a<��a<(�a<a<;�a<Ϗa<6�a<�a<`�a<�a<�a<�a<��a<,�a<�a<|�a<,�a<��a<a�a<�a<��a<e�a<�a<��a<8�a<�a<��a<@�a<�a<��a<��a<*�a<�a<��a<��a<��a<R�a<N�a< �a<�a<��a<܄a<քa<��a<��a<��a<��a<l�a<e�a<|�a<]�a<r�a<l�a<��a<��a<��a<ׄa<�a<�  �  �a<.�a<W�a<z�a<��a<��a<��a<'�a<M�a<z�a<��a<�a<8�a<o�a<��a<�a<d�a<��a<�a<e�a<ډa<E�a<��a<�a<w�a<�a<Z�a<��a<-�a<��a<�a<��a<�a<I�a<��a<\�a<ːa<U�a<�a<l�a<ܒa<n�a<�a<y�a<��a<z�a<��a<b�a<��a<n�a<ޗa<`�a<ʘa<R�a<ՙa<N�a<ƚa<E�a<��a<+�a<��a<%�a<��a<.�a<��a<�a<k�a<ϟa<:�a<��a<�a<0�a<��a<�a<%�a<a�a<��a< �a<,�a<��a<٣a<�a<3�a<�a<��a<�a<�a<9�a<_�a<��a<��a<ĥa<˥a<�a<��a<+�a<7�a<P�a<k�a<��a<��a<��a<Φa<�a< �a<�a<�a</�a<9�a<B�a<D�a<F�a<:�a<1�a<A�a<2�a<�a<�a<�a<��a<٦a<�a<�a<��a<��a<��a<��a<u�a<U�a<2�a<��a<�a<ɥa<��a<d�a<0�a<�a<�a<��a<��a<V�a<8�a<��a<֣a<��a<��a<a�a<'�a<�a<��a<��a<T�a<�a<ʡa<r�a<5�a<�a<��a<7�a<�a<��a<W�a<�a<ʞa<v�a<�a<��a<]�a<�a<��a<2�a<ɛa<B�a<�a<n�a<�a<}�a<��a<��a<�a<��a<"�a<��a<7�a<��a<P�a<Ӕa<m�a<	�a<{�a<�a<��a<$�a<��a<2�a<��a<4�a<Ϗa<Y�a<֎a<T�a<�a<��a<��a<��a<W�a<�a<p�a<"�a<a<j�a<�a<��a<E�a<�a<��a<?�a<ևa<��a<9�a<�a<��a<u�a<=�a<�a<Ӆa<��a<��a<_�a<G�a</�a<��a<�a<݄a<Ʉa<��a<��a<��a<x�a<��a<x�a<\�a<h�a<v�a<{�a<s�a<��a<Ȅa<Ʉa<�a<�  �  �a<E�a<N�a<m�a<��a<��a<�a<�a<]�a<h�a<��a<�a<�a<a�a<��a<��a<E�a<��a<��a<i�a<߉a<1�a<��a<��a<��a<׋a<S�a<֌a<+�a<��a<�a<��a<�a<o�a<��a<^�a<��a<O�a<�a<h�a<�a<x�a<�a<��a<�a<}�a<�a<{�a<��a<`�a<��a<?�a<��a<C�a<��a<8�a<��a</�a<��a<=�a<��a<9�a<��a<"�a<��a<��a<y�a<ßa<F�a<��a<�a<B�a<��a<�a<!�a<��a<��a<�a<S�a<��a<֣a<�a<S�a<�a<ɤa<�a<�a<P�a<N�a<��a<��a<åa<إa<֥a<�a<�a<)�a<5�a<Z�a<g�a<��a<��a<��a<��a<�a<�a<�a<5�a<2�a<:�a<V�a<A�a<R�a<5�a<9�a<2�a<�a<7�a<�a<"�a<�a<�a<ܦa<��a<Ȧa<��a<��a<l�a<H�a<<�a<�a<��a<��a<��a<Q�a<0�a<	�a<äa<��a<i�a<J�a<�a<��a<��a<��a<��a<M�a<B�a<�a<Ӣa<y�a<M�a<#�a<ǡa<��a<6�a<��a<��a<]�a< �a<��a<��a<	�a<˞a<s�a<�a<ȝa<_�a<�a<��a<5�a<��a<[�a<�a<a�a<�a<\�a<	�a<y�a<��a<��a<�a<��a<%�a<ƕa<.�a<�a<d�a<��a<��a<	�a<��a<�a<��a<;�a<Őa<F�a<̏a<Z�a<Ҏa<��a<��a<��a<&�a<��a<T�a<�a<��a<!�a<֊a<j�a<��a<��a<5�a<�a<��a<>�a<�a<v�a<A�a<�a<��a<Z�a<,�a<�a<υa<��a<k�a<u�a<5�a<6�a<	�a<��a<Մa<��a<ńa<��a<��a<|�a<|�a<w�a<c�a<��a<p�a<��a<��a<��a<��a<ʄa< �a<�  �  �a<&�a<d�a<z�a<��a<ƅa<�a<�a<I�a<r�a<��a<�a<�a<o�a<��a<�a<M�a<��a<�a<m�a<Ήa<1�a<��a<�a<��a<�a<\�a<��a<4�a<��a<�a<}�a<��a<w�a<ۏa<M�a<ݐa<d�a<ݑa<l�a<�a<p�a<�a<u�a<�a<��a< �a<r�a<�a<g�a<�a<P�a<ۘa<A�a<��a<G�a<ƚa<5�a<��a<<�a<��a<4�a<��a<�a<��a<�a<x�a<۟a<7�a<��a<�a<D�a<��a<ܡa<4�a<y�a<��a<��a<Q�a<��a<ɣa<�a<K�a<��a<��a<�a<�a<S�a<`�a<y�a<��a<��a<إa<�a<�a<�a<3�a<V�a<j�a<t�a<��a<��a<��a<�a<�a<�a<�a<=�a<>�a<U�a<;�a<J�a<E�a<J�a<6�a<3�a</�a<�a<��a<��a<�a<�a<Ԧa<צa<��a<��a<��a<��a<V�a<D�a<�a<ߥa<��a<��a<[�a<3�a<��a<Ϥa<��a<��a<S�a< �a<��a<ѣa<��a<}�a<M�a<�a<��a<բa<��a<V�a<�a<Сa<��a<M�a<�a<��a<e�a<�a<��a<i�a<�a<��a<w�a<�a<��a<^�a<��a<��a<:�a<͛a<Q�a<ݚa<g�a<��a<l�a<�a<w�a<�a<��a<"�a<��a<$�a<ŕa<D�a<�a<j�a<�a<��a<�a<��a<0�a<��a<3�a<��a<I�a<֏a<O�a<�a<l�a<�a<}�a<$�a<��a<G�a<��a<��a<(�a<��a<j�a<	�a<��a<F�a<�a<��a<5�a<�a<��a<?�a<�a<��a<z�a<<�a<��a<ǅa<��a<v�a<b�a<:�a<�a<
�a<�a<�a<܄a<��a<��a<��a<��a<z�a<y�a<{�a<q�a<`�a<�a<��a<��a<��a<�a<�a<�  �  N�a<Z�a<��a<��a<�a<�a<�a<p�a<z�a<��a<܇a<�a<e�a<��a<��a<,�a<��a<��a<7�a<��a<�a<��a<��a<J�a<��a<��a<n�a<ԍa<T�a<��a</�a<��a<&�a<��a<��a<��a<�a<��a<��a<Z�a<�a<j�a<��a<q�a<��a<s�a<�a<h�a<��a<��a<Әa<d�a<��a<=�a<��a<-�a<��a<%�a<��a<
�a<��a<�a<��a<�a<f�a<��a<F�a<��a<�a<g�a<��a<�a<Z�a<��a<%�a<E�a<��a<�a<$�a<��a<��a<�a<�a<b�a<��a<��a<�a<�a<\�a<S�a<��a<��a<��a<Ӧa<Ϧa<
�a<�a<8�a<;�a<e�a<i�a<��a<��a<��a<��a<��a<�a<&�a<�a<�a<�a<3�a<�a<3�a<�a<+�a<�a<��a<�a<�a<�a<�a<��a<��a<��a<��a<h�a<R�a<*�a<*�a<�a<Ʀa<ɦa<x�a<R�a<�a<إa<ϥa<��a<u�a<8�a<�a<̤a<��a<��a<u�a<_�a<��a<�a<��a<a�a<,�a<�a<��a<b�a<&�a<ˡa<��a<C�a<��a<��a<A�a<�a<��a<<�a<��a<��a<D�a<۝a<{�a<�a<Ɯa<5�a<ڛa<t�a<ؚa<z�a<�a<s�a<��a<��a<�a<��a<4�a<��a<X�a<ѕa<��a<�a<�a<3�a<��a<*�a<��a<=�a<Ƒa<P�a<ʐa<g�a<�a<s�a<�a<��a<7�a<�a<a�a<�a<��a<J�a<֋a<��a<�a<̊a<��a<�a<ԉa<t�a<�a<��a<T�a</�a<ڇa<��a<Z�a<6�a<�a<цa<��a<��a<��a<Y�a<G�a<:�a<�a<�a<݅a<߅a<��a<Ʌa<��a<��a<��a<��a<ƅa<��a<̅a<�a<ޅa<�a<�a<�  �  O�a<m�a<��a<��a<Ɇa<�a<�a<<�a<r�a<��a<�a<"�a<i�a<��a<�a<3�a<��a<�a<A�a<��a<�a<O�a<Ƌa<'�a<��a<�a<��a<�a<R�a<��a<5�a<��a<�a<|�a<��a<n�a<�a<f�a<�a<y�a<��a<z�a<�a<~�a< �a<|�a<�a<l�a<�a<Q�a<֘a<Q�a<Ιa<P�a<͚a<;�a<��a<4�a<��a<"�a<��a<�a<y�a<�a<m�a<џa<K�a<��a<�a<y�a<ˡa<(�a<w�a<��a<��a<Q�a<��a<�a< �a<^�a<��a<�a<)�a<`�a<��a<ҥa<��a<�a<3�a<b�a<o�a<��a<��a<צa<��a<�a<�a<8�a<K�a<u�a<��a<��a<��a<��a<˧a<�a<��a<�a<!�a<,�a</�a<9�a<&�a<-�a<�a<�a<��a<�a<�a<�a<Χa<ϧa<��a<��a<��a<��a<{�a<a�a<?�a<�a<�a<Ʀa<��a<q�a<I�a<'�a<��a<ԥa<��a<p�a<@�a<"�a<��a<Ȥa<��a<\�a<)�a<
�a<ϣa<��a<v�a<>�a<��a<��a<n�a<-�a<ڡa<��a<7�a<�a<��a<Q�a<�a<��a<\�a<�a<��a<S�a<�a<��a<�a<��a<8�a<ěa<D�a<ۚa<g�a<��a<��a<�a<��a<�a<��a<=�a<��a<J�a<֕a<Z�a<�a<��a<
�a<��a<4�a<Œa<O�a<Бa<a�a<�a<d�a<�a<�a<
�a<��a<2�a<ōa<g�a<�a<��a<H�a<�a<��a<0�a<Ɗa<b�a<�a<��a<T�a<�a<Èa<y�a<4�a<�a<��a<i�a<F�a<�a<�a<��a<��a<a�a<N�a<1�a<�a<�a<�a<�a<�a<Ņa<ąa<��a<��a<��a<��a<��a<��a<��a<ׅa<�a<�a<%�a<�  �  3�a<]�a<{�a<��a<͆a<��a<:�a<=�a<��a<��a<�a<�a<T�a<��a<�a<:�a<�a<�a<;�a<��a<�a<V�a<�a<)�a<��a<�a<b�a<؍a<?�a<��a< �a<��a<�a<��a<�a<b�a<�a<k�a<�a<p�a<�a<m�a<�a<k�a<�a<��a<�a<��a<��a<_�a<��a<H�a<ҙa<B�a<��a<1�a<��a<-�a<��a<(�a<��a<1�a<��a<	�a<��a<Пa<S�a<��a<�a<_�a<��a<�a<j�a<��a<�a<k�a<��a<�a<5�a<f�a<��a<�a<�a<K�a<��a<��a<�a<�a<2�a<��a<}�a<��a<ʦa<Ѧa<��a<��a<�a<7�a<N�a<a�a<��a<��a<��a<�a<ϧa<�a<
�a<�a<�a<�a<�a<�a<$�a<�a<�a<�a<�a<�a<اa<�a<�a<ӧa<ħa<��a<��a<z�a<k�a<L�a<<�a<�a<��a<�a<��a<��a<L�a<%�a<��a<��a<��a<r�a<G�a<�a<��a<¤a<��a<y�a<0�a<+�a<ѣa<��a<j�a< �a<�a<��a<i�a<�a<ڡa<��a<H�a<��a<��a<k�a<��a<��a<R�a<�a<��a<:�a<֝a<v�a< �a<��a<T�a<ٛa<R�a< �a<^�a<��a<x�a<�a<��a<�a<��a<,�a<Ŗa<E�a<��a<m�a<�a<��a<	�a<��a<$�a<��a<5�a<��a<K�a<ېa<f�a<�a<��a<�a<��a<G�a<͍a<h�a<��a<��a<2�a<׋a<r�a<!�a<Ίa<a�a<4�a<��a<n�a< �a<��a<}�a< �a<�a<��a<m�a<2�a<�a<�a<��a<��a<e�a<j�a<D�a<�a<�a<�a<݅a<ʅa<Åa<��a<��a<��a<��a<ǅa<��a<хa<Ʌa<܅a<�a<��a<"�a<�  �  H�a<e�a<��a<��a<݆a< �a<�a<M�a<s�a<��a<��a<�a<e�a<��a<��a<:�a<��a<��a<Q�a<��a<��a<f�a<��a<B�a<��a<�a<y�a<��a<Y�a<��a<.�a<~�a<�a<v�a<�a<o�a<בa<x�a<�a<d�a<��a<{�a<��a<�a<��a<k�a<�a<d�a<�a<g�a<ؘa<f�a<ۙa<O�a<Ěa<E�a<��a<4�a<��a<,�a<��a<�a<��a<��a<_�a<�a<@�a<��a<�a<u�a<ѡa<�a<e�a<��a<�a<5�a<��a<أa<�a<u�a<��a<�a<#�a<j�a<��a<ĥa<�a<�a<S�a<H�a<��a<��a<��a<�a<�a<�a<!�a<E�a<Y�a<n�a<��a<��a<��a<��a<�a<�a<�a<%�a<�a<.�a<+�a<.�a<(�a<,�a<�a<�a<�a<�a<�a<ڧa<ۧa<ӧa<��a<��a<��a<��a<t�a<b�a<.�a<&�a<��a<��a<��a<q�a<V�a<3�a<�a<Хa<��a<|�a<G�a<!�a<�a<ؤa<��a<i�a<A�a<�a<�a<��a<i�a<6�a<�a<��a<k�a<&�a<��a<��a<1�a<�a<��a<5�a<�a<��a<F�a<��a<��a<K�a<�a<��a<
�a<Üa<1�a<ʛa<Z�a<ݚa<|�a<�a<��a<
�a<��a<'�a<��a<<�a<ɖa<c�a<ܕa<k�a<��a<w�a<+�a<��a</�a<��a<K�a<בa<V�a<Րa<V�a<��a<d�a<�a<��a<"�a<܍a<O�a<	�a<��a<Q�a<�a<��a<%�a<ϊa<��a<��a<��a<c�a<�a<Ԉa<t�a<2�a<�a<��a<x�a<?�a<�a<�a<��a<��a<u�a<M�a<@�a<8�a< �a<�a<�a<څa<ǅa<a<��a<��a<��a<��a<��a<��a<ąa<ۅa<ԅa<�a<&�a<�  �  B�a<K�a<��a<��a<Ԇa<�a<�a<p�a<r�a<a<�a<�a<p�a<��a<��a<1�a<��a<ۉa<M�a<��a<��a<��a<��a<H�a<��a<�a<z�a<Ǎa<J�a<��a<:�a<{�a<�a<t�a<�a<}�a<͑a<r�a<֒a<w�a<�a<\�a<�a<f�a<�a<a�a<�a<h�a<��a<}�a<٘a<q�a<ʙa<R�a<Śa<H�a<śa<0�a<��a<�a<��a<�a<��a<�a<a�a<��a</�a<��a<�a<d�a<��a<�a<u�a<��a<�a<.�a<��a<ףa<�a<s�a<��a<��a<��a<S�a<�a<åa<��a<�a<X�a<P�a<��a<��a<Ŧa<�a<�a<�a<�a<H�a<O�a<v�a<��a<��a<ɧa<��a<��a<�a<�a<�a<�a<4�a<�a<$�a<�a<(�a<�a<�a<�a<�a<�a<Χa<֧a<ŧa<��a<��a<|�a<��a<Y�a<f�a<0�a<�a< �a<Ħa<Ȧa<q�a<c�a<(�a<��a<ۥa<��a<�a<=�a<2�a<�a<Ԥa<��a<j�a<_�a<��a<�a<��a<p�a<7�a<٢a<��a<B�a<2�a<��a<��a</�a<�a<��a<+�a<��a<��a<Y�a<�a<��a<=�a<ѝa<��a<�a<Ŝa<4�a<ޛa<p�a<ޚa<��a<�a<��a<�a<��a<+�a<��a<A�a<��a<d�a<ݕa<��a<�a<z�a<2�a<��a<9�a<��a<:�a<��a<A�a<�a<J�a<��a<\�a<�a<��a<"�a<ڍa<I�a<�a<��a<;�a<ыa<��a<.�a<��a<��a<�a<ۉa<l�a<�a<ӈa<k�a<B�a<�a<��a<n�a<G�a<�a<ކa<Άa<��a<��a<R�a<>�a<2�a< �a<
�a<ͅa<Ѕa<��a<��a<��a<��a<��a<��a<��a<��a<��a<ͅa<ׅa<�a<�a<�  �  H�a<Y�a<|�a<��a<ʆa<��a<*�a<O�a<��a<��a<�a<7�a<m�a<��a<
�a<J�a<��a<��a<<�a<��a<�a<`�a<؋a<-�a<��a<�a<c�a<׍a<W�a<��a<�a<��a<�a<m�a<�a<V�a<�a<R�a<ڒa<i�a<ݓa<p�a<��a<j�a<��a<{�a<�a<y�a<�a<b�a<�a<P�a<�a<Z�a<Кa<R�a<͛a<@�a<��a<?�a<��a<'�a<��a<�a<|�a<ٟa<L�a<��a<��a<p�a<��a<�a<_�a<��a<�a<H�a<�a<ϣa<�a<C�a<��a<٤a<�a<a�a<��a<��a<��a<�a<:�a<s�a<�a<��a<̦a<̦a<�a<�a<0�a<U�a<e�a<v�a<��a<��a<��a<ߧa<ާa<��a<	�a<�a<�a<�a<�a<.�a<�a<�a<�a<��a<�a<��a<קa<�a<ŧa<��a<��a<��a<��a<��a<g�a<M�a<9�a<�a<��a<צa<��a<��a<S�a<(�a<�a<إa<��a<��a<W�a<'�a<�a<äa<��a<v�a<:�a<�a<գa<��a<q�a< �a<�a<��a<S�a<�a<ˡa<e�a<(�a<�a<��a<K�a<ߟa<��a<K�a<�a<��a<K�a<ԝa<{�a<�a<��a<E�a<қa<U�a<��a<f�a<�a<��a<�a<��a<4�a<��a<A�a<ܖa<E�a<�a<j�a<��a<��a<�a<��a<.�a<��a<F�a<Ǒa<@�a<Аa<S�a<׏a<v�a<��a<��a<$�a<��a<Y�a<��a<��a<H�a<ߋa<u�a<,�a<Ɋa<i�a<%�a<��a<k�a<"�a<��a<��a<6�a<��a<Ƈa<��a<G�a< �a<�a<��a<��a<s�a<^�a<D�a<�a<�a<�a<ۅa<څa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<�a<��a<�a<�  �  "�a<f�a<t�a<��a<цa<��a<8�a<J�a<��a<��a<�a<=�a<f�a<ˈa<�a<b�a<��a<�a<U�a<��a<�a<_�a<�a<'�a<��a< �a<m�a<�a<3�a<��a<��a<��a<��a<a�a<�a<M�a<�a<:�a<��a<Q�a<�a<i�a<ߔa<��a<�a<��a<�a<~�a<��a<n�a< �a<R�a<�a<M�a<ٚa<\�a<Λa<O�a<��a<c�a<��a<6�a<��a<�a<��a<ԟa<c�a<��a<�a<^�a<��a<�a<F�a<̢a<բa<A�a<y�a<Уa<�a<@�a<��a<��a<!�a<E�a<��a<��a<�a<4�a<2�a<~�a<��a<��a<ͦa<�a<'�a<�a<H�a<A�a<y�a<x�a<��a<Чa<��a<�a<ߧa<	�a<�a<�a<)�a<�a</�a<	�a<"�a< �a<�a<�a<ܧa<��a<ħa<ߧa<��a<��a<��a<��a<��a<i�a<u�a<E�a<:�a<�a<�a<�a<��a<��a<O�a<N�a<�a<ѥa<ťa<u�a<o�a<�a<�a<ܤa<��a<��a<9�a<)�a<ϣa<��a<e�a<*�a<�a<��a<j�a<��a<�a<m�a<�a<�a<x�a<C�a<ǟa<��a<4�a<�a<��a<+�a<�a<h�a<3�a<��a<K�a<ߛa<b�a<�a<h�a<4�a<��a<�a<��a<4�a<Ɨa<4�a<�a<P�a<��a<y�a<
�a<��a<�a<��a<�a<��a<4�a<��a<L�a<��a<x�a<��a<o�a<��a<��a<�a<��a<z�a<׌a<��a<,�a<��a<��a<�a<�a<a�a<0�a<��a<{�a<#�a<Јa<��a<(�a<�a<��a<��a<I�a<!�a<�a<��a<��a<u�a<n�a<A�a<#�a<�a<�a<�a<��a<��a<��a<��a<��a<w�a<��a<|�a<��a<��a<Ʌa<�a<��a<#�a<�  �  (�a<X�a<|�a<��a<Ԇa<��a<-�a<q�a<��a<Ǉa<�a<0�a<y�a<͈a< �a<h�a<��a<��a<c�a<��a<�a<��a<ыa<9�a<��a<�a<k�a<эa</�a<��a<��a<|�a<�a<^�a<ېa<\�a<ϑa<G�a<ےa<;�a<ޓa<Y�a<ܔa<w�a<�a<x�a< �a<r�a<�a<��a<�a<r�a<�a<W�a<�a<\�a<ћa<V�a<��a<@�a<��a<'�a<��a<�a<p�a<�a<K�a<��a<�a<T�a<��a<�a<5�a<��a<�a</�a<�a<£a< �a<K�a<��a<��a<�a<;�a<��a<��a<ܥa<�a<D�a<g�a<��a<��a<˦a<��a<�a<�a<P�a<M�a<x�a<��a<��a<��a<ͧa<קa<�a<��a<�a<�a<�a<�a<"�a<�a<�a<�a<�a<��a<�a<ߧa<�a<ɧa<��a<��a<��a<��a<��a<o�a<g�a<N�a<2�a<�a<��a<ڦa<ɦa<��a<h�a<I�a<�a<�a<ȥa<��a<u�a<2�a<�a<�a<��a<��a<^�a<�a<�a<��a<Z�a<(�a<�a<��a<\�a<��a<��a<q�a<�a<Рa<��a<,�a<ԟa<��a<�a<�a<��a<)�a<�a<q�a<�a<��a<>�a<�a<z�a<��a<��a<�a<��a<(�a<��a<8�a<͗a<H�a<ݖa<j�a<�a<��a<�a<��a< �a<��a<"�a<��a<*�a<��a<?�a<��a<T�a<͏a<^�a<��a<��a<�a<��a<P�a<֌a<��a<"�a<Ӌa<|�a<�a<͊a<s�a<�a<݉a<�a<!�a<�a<��a<@�a<�a<��a<��a<U�a<�a<�a<҆a<��a<��a<e�a<;�a<-�a<	�a<�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<Ņa<�a<�a<�  �  I�a<C�a<��a<��a<Άa<�a<�a<i�a<{�a<�a<��a<I�a<��a<��a<,�a<J�a<��a<��a<c�a<Ŋa<��a<v�a<ċa<N�a<��a<�a<b�a<ɍa<O�a<��a<�a<k�a<�a<Z�a<ɐa<R�a<��a<R�a<��a<X�a<Փa<`�a<��a<U�a<
�a<`�a<�a<��a<��a<z�a<�a<��a<ߙa<��a<ښa<h�a<�a<A�a<�a<4�a<ӝa<$�a<��a<�a<y�a<�a</�a<��a<�a<k�a<��a<��a<U�a<��a<�a<�a<w�a<��a<��a<?�a<v�a<٤a<��a<X�a<��a<��a<��a<�a<X�a<_�a<��a<��a<ۦa<�a<�a<9�a</�a<x�a<u�a<��a<��a<��a<�a<ŧa<��a<�a<�a<�a<�a<,�a<�a<0�a<�a<�a<��a<ߧa<�a<ħa<ѧa<��a<��a<��a<��a<��a<r�a<��a<R�a<Z�a<5�a<�a<�a<˦a<¦a<z�a<��a<6�a<�a<�a<��a<��a<W�a<J�a<�a<�a<��a<m�a<P�a<�a<��a<��a<x�a< �a<ۢa<��a<>�a<�a<��a<_�a<�a<��a<}�a<�a<��a<o�a<;�a<ޞa<��a<H�a<��a<��a<��a<��a<M�a<ԛa<m�a<�a<��a<�a<��a< �a<��a<M�a<��a<n�a<іa<��a<�a<|�a<	�a<��a<)�a<��a<A�a<��a<A�a<��a<1�a<Őa</�a<ҏa<M�a<�a<x�a<	�a<��a<6�a<��a<y�a<?�a<؋a<n�a<7�a<��a<��a<�a<Ήa<i�a<0�a<�a<��a<^�a<��a<�a<��a<`�a<;�a<�a<�a<��a<��a<T�a<S�a<*�a<�a<�a<ąa<܅a<��a<��a<��a<t�a<��a<k�a<��a<}�a<��a<��a<Ʌa<�a<��a<�  �  &�a<<�a<��a<��a<ˆa<�a<6�a<q�a<��a<߇a<��a<W�a<��a<ǈa<�a<X�a<��a<�a<V�a<ʊa<!�a<��a<�a<G�a<��a<�a<f�a<Ía<1�a<��a<�a<|�a<��a<S�a<ϐa<N�a<��a<F�a<Òa<Y�a<˓a<S�a<ߔa<M�a<�a<y�a<��a<��a<
�a<��a<�a<��a<�a<��a<ݚa<g�a<�a<H�a<�a<>�a<ĝa<<�a<��a<"�a<��a<�a<C�a<��a<�a<T�a<��a<�a<V�a<��a<ޢa<"�a<r�a<��a<��a<<�a<��a<ˤa<��a<?�a<w�a<��a< �a<�a<P�a<z�a<��a<Ħa<�a<�a<�a<?�a<;�a<f�a<x�a<��a<��a<��a<�a<�a<�a<�a<�a<�a<#�a<&�a<��a<�a<�a<��a<�a<�a<�a<Чa<ͧa<��a<��a<��a<��a<��a<s�a<m�a<K�a<U�a<@�a<�a<�a<�a<ɦa<��a<�a<5�a<.�a<��a<��a<��a<d�a<N�a<�a<ݤa<Ǥa<��a<]�a<$�a<�a<��a<}�a<#�a<բa<��a<:�a<�a<��a<^�a<�a<àa<y�a<�a<ӟa<|�a<;�a<Ԟa<�a<+�a<��a<��a<�a<��a<P�a<�a<��a<�a<��a<�a<��a<#�a<��a<I�a<��a<m�a<ۖa<v�a<�a<��a<�a<��a<�a<��a<9�a<��a<*�a<��a<,�a<ǐa<>�a<ɏa<Q�a<�a<w�a<�a<��a<H�a<�a<u�a<&�a<ɋa<m�a<8�a<��a<�a<,�a<܉a<��a<<�a<݈a<��a<d�a<�a<ׇa<��a<d�a<H�a<�a<�a<��a<��a<m�a<R�a<$�a<�a<��a<��a<��a<��a<��a<��a<y�a<}�a<x�a<��a<��a<��a<��a<хa<�a<��a<�  �  �a<i�a<x�a<��a<׆a<��a<0�a<[�a<��a<̇a<�a<S�a<��a<�a<�a<��a<��a<�a<i�a<��a<�a<s�a<ҋa<2�a<��a<��a<o�a<ۍa<"�a<��a<��a<p�a<ۏa<H�a<Ða<>�a<��a<3�a<ɒa<A�a<��a<\�a<ݔa<��a<��a<|�a<��a<p�a<��a<s�a<��a<}�a<��a<w�a<�a<u�a<�a<z�a<לa<R�a<ŝa<2�a<��a<
�a<s�a<ܟa<R�a<��a<�a<Y�a<��a<�a<:�a<��a<͢a<�a<^�a<��a<�a<1�a<|�a<��a<�a<4�a<��a<ťa<ޥa<"�a<@�a<h�a<��a<��a<ئa< �a<�a<4�a<o�a<U�a<��a<��a<��a<̧a<Чa<�a<�a< �a<�a<�a<�a<�a<1�a< �a<�a< �a<�a<�a<̧a<Χa<§a<��a<��a<��a<��a<��a<��a<]�a<w�a<J�a<4�a<�a<��a<ݦa<��a<��a<m�a<T�a<*�a<�a<�a<��a<��a<J�a< �a<�a<��a<��a<N�a<�a<ڣa<��a<\�a<-�a<�a<��a<_�a<�a<��a<X�a<�a<��a<i�a<�a<��a<��a<#�a<�a<��a<)�a<�a<f�a<�a<��a<<�a<֛a<f�a<�a<��a<#�a<��a<L�a<˘a<M�a<�a<a�a<�a<w�a<��a<|�a<�a<��a<�a<��a<�a<Œa</�a<��a<G�a<��a<>�a<��a<K�a<Ԏa<f�a<��a<��a<=�a<̌a<��a<�a<ًa<��a<�a<ӊa<o�a<�a<ˉa<�a<.�a<�a<��a<Y�a<8�a<Ƈa<��a<u�a<=�a<�a<Նa<��a<��a<f�a<=�a<*�a<�a<�a<��a<��a<��a<��a<��a<~�a<h�a<v�a<{�a<��a<��a<��a<Åa<ޅa<�a<�  �  �a<H�a<n�a<��a<ۆa<�a<A�a<u�a<��a<��a<�a<N�a<��a<ֈa<�a<o�a<��a<�a<g�a<Ίa<�a<��a<�a<E�a<��a<��a<[�a<��a<�a<��a<��a<o�a<�a<]�a<Ða<B�a<��a<G�a<Ēa<G�a<ȓa<F�a<̔a<h�a<�a<t�a<�a<��a<�a<��a<
�a<��a<��a<o�a<�a<n�a<�a<`�a<ќa<O�a<ԝa<F�a<��a<#�a<��a<�a<J�a<��a<��a<D�a<��a<�a<>�a<��a<�a< �a<f�a<��a<��a<@�a<z�a<��a<��a<(�a<r�a<��a<ݥa<�a<P�a<y�a<��a<Ħa<�a<�a<�a<.�a<T�a<d�a<��a<��a<��a<ʧa<�a<�a<�a<�a<�a<�a<�a<�a<�a<��a<��a<��a<��a<�a<�a<Ƨa<��a<��a<��a<��a<��a<��a<q�a<[�a<W�a<@�a</�a<$�a<�a<�a<ͦa<��a<��a<Q�a<%�a<�a<ѥa<��a<|�a<@�a<�a<�a<ʤa<��a<h�a<&�a<�a<��a<Z�a<�a<Ңa<}�a<<�a<�a<��a<c�a<�a<��a<m�a<�a<ԟa<}�a<)�a<Оa<q�a<�a<ҝa<i�a<�a<��a<^�a<�a<|�a<�a<��a< �a<��a<5�a<Ęa<K�a<ؗa<[�a<�a<��a<�a<��a<�a<��a<%�a<��a<�a<��a<�a<��a<&�a<��a<7�a<ˏa<O�a<ݎa<m�a<�a<��a<;�a<Ռa<w�a<�a<ŋa<n�a<�a<Њa<�a<*�a<�a<��a<B�a<�a<��a<S�a<�a<Շa<��a<c�a<6�a<�a<�a<��a<��a<v�a<X�a<3�a<�a<�a<υa<��a<��a<��a<��a<~�a<|�a<m�a<x�a<z�a<��a<��a<Ņa<مa<��a<�  �  H�a<B�a<��a<��a<Ɔa<��a<,�a<u�a<��a<�a<�a<i�a<��a<Јa<9�a<a�a<͉a<$�a<R�a<Њa<�a<��a<ыa<8�a<��a<�a<k�a<΍a<N�a<��a<�a<]�a<ɏa<G�a<��a<?�a<��a<B�a<��a<E�a<��a<g�a<�a<Y�a<�a<x�a<�a<�a<��a<��a<��a<�a<��a<��a<�a<y�a<�a<Y�a<��a<O�a<��a<5�a<��a<�a<�a<ߟa<H�a<��a<�a<`�a<��a<�a<G�a<o�a<٢a<�a<_�a<��a<�a<'�a<h�a<ˤa<�a<Y�a<��a<��a<�a<�a<D�a<k�a<��a<��a<�a<�a<*�a<R�a<E�a<��a<��a<��a<ʧa<��a<�a<�a<�a<��a<�a<
�a< �a<.�a<�a<2�a<�a<��a<�a<ħa<ާa<��a<ȧa<��a<��a<��a<��a<��a<~�a<��a<Q�a<\�a<D�a<�a<��a<٦a<Φa<��a<��a<A�a<@�a<�a<ʥa<��a<m�a<\�a<1�a<٤a<ͤa<�a<`�a<�a<�a<��a<|�a<(�a<�a<��a<;�a<�a<��a<F�a<�a<��a<i�a<�a<ϟa<[�a<'�a<ɞa<��a<>�a<Ýa<��a<�a<��a<K�a<ڛa<}�a< �a<��a<�a<˙a<8�a<Ϙa<Z�a<їa<��a<�a<n�a<��a<��a<�a<��a<�a<��a<A�a<��a<6�a<��a< �a<��a<�a<ďa<@�a<Վa<\�a<��a<��a<(�a<�a<s�a<@�a<ًa<p�a<8�a<Ɗa<s�a<�a<ىa<y�a<9�a<Ոa<��a<w�a<�a<�a<��a<s�a<R�a<��a<�a<��a<��a<c�a<F�a<�a<�a<�a<Ņa<ޅa<��a<��a<}�a<Y�a<z�a<g�a<��a<q�a<��a<��a<��a<ޅa<�a<�  �  �a<H�a<n�a<��a<ۆa<�a<A�a<u�a<��a<��a<�a<N�a<��a<ֈa<�a<o�a<��a<�a<g�a<Ίa<�a<��a<�a<E�a<��a<��a<[�a<��a<�a<��a<��a<o�a<�a<]�a<Ða<B�a<��a<G�a<Ēa<G�a<ȓa<F�a<̔a<h�a<�a<t�a<�a<��a<�a<��a<
�a<��a<��a<o�a<�a<n�a<�a<`�a<ќa<O�a<ԝa<F�a<��a<#�a<��a<�a<J�a<��a<��a<D�a<��a<�a<>�a<��a<�a< �a<f�a<��a<��a<@�a<z�a<��a<��a<(�a<r�a<��a<ݥa<�a<P�a<y�a<��a<Ħa<�a<�a<�a<.�a<T�a<d�a<��a<��a<��a<ʧa<�a<�a<�a<�a<�a<�a<�a<�a<�a<��a<��a<��a<��a<�a<�a<Ƨa<��a<��a<��a<��a<��a<��a<q�a<[�a<W�a<@�a</�a<$�a<�a<�a<ͦa<��a<��a<Q�a<%�a<�a<ѥa<��a<|�a<@�a<�a<�a<ʤa<��a<h�a<&�a<�a<��a<Z�a<�a<Ңa<}�a<<�a<�a<��a<c�a<�a<��a<m�a<�a<ԟa<}�a<)�a<Оa<q�a<�a<ҝa<i�a<�a<��a<^�a<�a<|�a<�a<��a< �a<��a<5�a<Ęa<K�a<ؗa<[�a<�a<��a<�a<��a<�a<��a<%�a<��a<�a<��a<�a<��a<&�a<��a<7�a<ˏa<O�a<ݎa<m�a<�a<��a<;�a<Ռa<w�a<�a<ŋa<n�a<�a<Њa<�a<*�a<�a<��a<B�a<�a<��a<S�a<�a<Շa<��a<c�a<6�a<�a<�a<��a<��a<v�a<X�a<3�a<�a<�a<υa<��a<��a<��a<��a<~�a<|�a<m�a<x�a<z�a<��a<��a<Ņa<مa<��a<�  �  �a<i�a<x�a<��a<׆a<��a<0�a<[�a<��a<̇a<�a<S�a<��a<�a<�a<��a<��a<�a<i�a<��a<�a<s�a<ҋa<2�a<��a<��a<o�a<ۍa<"�a<��a<��a<p�a<ۏa<H�a<Ða<>�a<��a<3�a<ɒa<A�a<��a<\�a<ݔa<��a<��a<|�a<��a<p�a<��a<s�a<��a<}�a<��a<w�a<�a<u�a<�a<z�a<לa<R�a<ŝa<2�a<��a<
�a<s�a<ܟa<R�a<��a<�a<Y�a<��a<�a<:�a<��a<͢a<�a<^�a<��a<�a<1�a<|�a<��a<�a<4�a<��a<ťa<ޥa<"�a<@�a<h�a<��a<��a<ئa< �a<�a<4�a<o�a<U�a<��a<��a<��a<̧a<Чa<�a<�a< �a<�a<�a<�a<�a<1�a< �a<�a< �a<�a<�a<̧a<Χa<§a<��a<��a<��a<��a<��a<��a<]�a<w�a<J�a<4�a<�a<��a<ݦa<��a<��a<m�a<T�a<*�a<�a<�a<��a<��a<J�a< �a<�a<��a<��a<N�a<�a<ڣa<��a<\�a<-�a<�a<��a<_�a<�a<��a<X�a<�a<��a<i�a<�a<��a<��a<#�a<�a<��a<)�a<�a<f�a<�a<��a<<�a<֛a<f�a<�a<��a<#�a<��a<L�a<˘a<M�a<�a<a�a<�a<w�a<��a<|�a<�a<��a<�a<��a<�a<Œa</�a<��a<G�a<��a<>�a<��a<K�a<Ԏa<f�a<��a<��a<=�a<̌a<��a<�a<ًa<��a<�a<ӊa<o�a<�a<ˉa<�a<.�a<�a<��a<Y�a<8�a<Ƈa<��a<u�a<=�a<�a<Նa<��a<��a<f�a<=�a<*�a<�a<�a<��a<��a<��a<��a<��a<~�a<h�a<v�a<{�a<��a<��a<��a<Åa<ޅa<�a<�  �  &�a<<�a<��a<��a<ˆa<�a<6�a<q�a<��a<߇a<��a<W�a<��a<ǈa<�a<X�a<��a<�a<V�a<ʊa<!�a<��a<�a<G�a<��a<�a<f�a<Ía<1�a<��a<�a<|�a<��a<S�a<ϐa<N�a<��a<F�a<Òa<Y�a<˓a<S�a<ߔa<M�a<�a<y�a<��a<��a<
�a<��a<�a<��a<�a<��a<ݚa<g�a<�a<H�a<�a<>�a<ĝa<<�a<��a<"�a<��a<�a<C�a<��a<�a<T�a<��a<�a<V�a<��a<ޢa<"�a<r�a<��a<��a<<�a<��a<ˤa<��a<?�a<w�a<��a< �a<�a<P�a<z�a<��a<Ħa<�a<�a<�a<?�a<;�a<f�a<x�a<��a<��a<��a<�a<�a<�a<�a<�a<�a<#�a<&�a<��a<�a<�a<��a<�a<�a<�a<Чa<ͧa<��a<��a<��a<��a<��a<s�a<m�a<K�a<U�a<@�a<�a<�a<�a<ɦa<��a<�a<5�a<.�a<��a<��a<��a<d�a<N�a<�a<ݤa<Ǥa<��a<]�a<$�a<�a<��a<}�a<#�a<բa<��a<:�a<�a<��a<^�a<�a<àa<y�a<�a<ӟa<|�a<;�a<Ԟa<�a<+�a<��a<��a<�a<��a<P�a<�a<��a<�a<��a<�a<��a<#�a<��a<I�a<��a<m�a<ۖa<v�a<�a<��a<�a<��a<�a<��a<9�a<��a<*�a<��a<,�a<ǐa<>�a<ɏa<Q�a<�a<w�a<�a<��a<H�a<�a<u�a<&�a<ɋa<m�a<8�a<��a<�a<,�a<܉a<��a<<�a<݈a<��a<d�a<�a<ׇa<��a<d�a<H�a<�a<�a<��a<��a<m�a<R�a<$�a<�a<��a<��a<��a<��a<��a<��a<y�a<}�a<x�a<��a<��a<��a<��a<хa<�a<��a<�  �  I�a<C�a<��a<��a<Άa<�a<�a<i�a<{�a<�a<��a<I�a<��a<��a<,�a<J�a<��a<��a<c�a<Ŋa<��a<v�a<ċa<N�a<��a<�a<b�a<ɍa<O�a<��a<�a<k�a<�a<Z�a<ɐa<R�a<��a<R�a<��a<X�a<Փa<`�a<��a<U�a<
�a<`�a<�a<��a<��a<z�a<�a<��a<ߙa<��a<ښa<h�a<�a<A�a<�a<4�a<ӝa<$�a<��a<�a<y�a<�a</�a<��a<�a<k�a<��a<��a<U�a<��a<�a<�a<w�a<��a<��a<?�a<v�a<٤a<��a<X�a<��a<��a<��a<�a<X�a<_�a<��a<��a<ۦa<�a<�a<9�a</�a<x�a<u�a<��a<��a<��a<�a<ŧa<��a<�a<�a<�a<�a<,�a<�a<0�a<�a<�a<��a<ߧa<�a<ħa<ѧa<��a<��a<��a<��a<��a<r�a<��a<R�a<Z�a<5�a<�a<�a<˦a<¦a<z�a<��a<6�a<�a<�a<��a<��a<W�a<J�a<�a<�a<��a<m�a<P�a<�a<��a<��a<x�a< �a<ۢa<��a<>�a<�a<��a<_�a<�a<��a<}�a<�a<��a<o�a<;�a<ޞa<��a<H�a<��a<��a<��a<��a<M�a<ԛa<m�a<�a<��a<�a<��a< �a<��a<M�a<��a<n�a<іa<��a<�a<|�a<	�a<��a<)�a<��a<A�a<��a<A�a<��a<1�a<Őa</�a<ҏa<M�a<�a<x�a<	�a<��a<6�a<��a<y�a<?�a<؋a<n�a<7�a<��a<��a<�a<Ήa<i�a<0�a<�a<��a<^�a<��a<�a<��a<`�a<;�a<�a<�a<��a<��a<T�a<S�a<*�a<�a<�a<ąa<܅a<��a<��a<��a<t�a<��a<k�a<��a<}�a<��a<��a<Ʌa<�a<��a<�  �  (�a<X�a<|�a<��a<Ԇa<��a<-�a<q�a<��a<Ǉa<�a<0�a<y�a<͈a< �a<h�a<��a<��a<c�a<��a<�a<��a<ыa<9�a<��a<�a<k�a<эa</�a<��a<��a<|�a<�a<^�a<ېa<\�a<ϑa<G�a<ےa<;�a<ޓa<Y�a<ܔa<w�a<�a<x�a< �a<r�a<�a<��a<�a<r�a<�a<W�a<�a<\�a<ћa<V�a<��a<@�a<��a<'�a<��a<�a<p�a<�a<K�a<��a<�a<T�a<��a<�a<5�a<��a<�a</�a<�a<£a< �a<K�a<��a<��a<�a<;�a<��a<��a<ܥa<�a<D�a<g�a<��a<��a<˦a<��a<�a<�a<P�a<M�a<x�a<��a<��a<��a<ͧa<קa<�a<��a<�a<�a<�a<�a<"�a<�a<�a<�a<�a<��a<�a<ߧa<�a<ɧa<��a<��a<��a<��a<��a<o�a<g�a<N�a<2�a<�a<��a<ڦa<ɦa<��a<h�a<I�a<�a<�a<ȥa<��a<u�a<2�a<�a<�a<��a<��a<^�a<�a<�a<��a<Z�a<(�a<�a<��a<\�a<��a<��a<q�a<�a<Рa<��a<,�a<ԟa<��a<�a<�a<��a<)�a<�a<q�a<�a<��a<>�a<�a<z�a<��a<��a<�a<��a<(�a<��a<8�a<͗a<H�a<ݖa<j�a<�a<��a<�a<��a< �a<��a<"�a<��a<*�a<��a<?�a<��a<T�a<͏a<^�a<��a<��a<�a<��a<P�a<֌a<��a<"�a<Ӌa<|�a<�a<͊a<s�a<�a<݉a<�a<!�a<�a<��a<@�a<�a<��a<��a<U�a<�a<�a<҆a<��a<��a<e�a<;�a<-�a<	�a<�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<Ņa<�a<�a<�  �  "�a<f�a<t�a<��a<цa<��a<8�a<J�a<��a<��a<�a<=�a<f�a<ˈa<�a<b�a<��a<�a<U�a<��a<�a<_�a<�a<'�a<��a< �a<m�a<�a<3�a<��a<��a<��a<��a<a�a<�a<M�a<�a<:�a<��a<Q�a<�a<i�a<ߔa<��a<�a<��a<�a<~�a<��a<n�a< �a<R�a<�a<M�a<ٚa<\�a<Λa<O�a<��a<c�a<��a<6�a<��a<�a<��a<ԟa<c�a<��a<�a<^�a<��a<�a<F�a<̢a<բa<A�a<y�a<Уa<�a<@�a<��a<��a<!�a<E�a<��a<��a<�a<4�a<2�a<~�a<��a<��a<ͦa<�a<'�a<�a<H�a<A�a<y�a<x�a<��a<Чa<��a<�a<ߧa<	�a<�a<�a<)�a<�a</�a<	�a<"�a< �a<�a<�a<ܧa<��a<ħa<ߧa<��a<��a<��a<��a<��a<i�a<u�a<E�a<:�a<�a<�a<�a<��a<��a<O�a<N�a<�a<ѥa<ťa<u�a<o�a<�a<�a<ܤa<��a<��a<9�a<)�a<ϣa<��a<e�a<*�a<�a<��a<j�a<��a<�a<m�a<�a<�a<x�a<C�a<ǟa<��a<4�a<�a<��a<+�a<�a<h�a<3�a<��a<K�a<ߛa<b�a<�a<h�a<4�a<��a<�a<��a<4�a<Ɨa<4�a<�a<P�a<��a<y�a<
�a<��a<�a<��a<�a<��a<4�a<��a<L�a<��a<x�a<��a<o�a<��a<��a<�a<��a<z�a<׌a<��a<,�a<��a<��a<�a<�a<a�a<0�a<��a<{�a<#�a<Јa<��a<(�a<�a<��a<��a<I�a<!�a<�a<��a<��a<u�a<n�a<A�a<#�a<�a<�a<�a<��a<��a<��a<��a<��a<w�a<��a<|�a<��a<��a<Ʌa<�a<��a<#�a<�  �  H�a<Y�a<|�a<��a<ʆa<��a<*�a<O�a<��a<��a<�a<7�a<m�a<��a<
�a<J�a<��a<��a<<�a<��a<�a<`�a<؋a<-�a<��a<�a<c�a<׍a<W�a<��a<�a<��a<�a<m�a<�a<V�a<�a<R�a<ڒa<i�a<ݓa<p�a<��a<j�a<��a<{�a<�a<y�a<�a<b�a<�a<P�a<�a<Z�a<Кa<R�a<͛a<@�a<��a<?�a<��a<'�a<��a<�a<|�a<ٟa<L�a<��a<��a<p�a<��a<�a<_�a<��a<�a<H�a<�a<ϣa<�a<C�a<��a<٤a<�a<a�a<��a<��a<��a<�a<:�a<s�a<�a<��a<̦a<̦a<�a<�a<0�a<U�a<e�a<v�a<��a<��a<��a<ߧa<ާa<��a<	�a<�a<�a<�a<�a<.�a<�a<�a<�a<��a<�a<��a<קa<�a<ŧa<��a<��a<��a<��a<��a<g�a<M�a<9�a<�a<��a<צa<��a<��a<S�a<(�a<�a<إa<��a<��a<W�a<'�a<�a<äa<��a<v�a<:�a<�a<գa<��a<q�a< �a<�a<��a<S�a<�a<ˡa<e�a<(�a<�a<��a<K�a<ߟa<��a<K�a<�a<��a<K�a<ԝa<{�a<�a<��a<E�a<қa<U�a<��a<f�a<�a<��a<�a<��a<4�a<��a<A�a<ܖa<E�a<�a<j�a<��a<��a<�a<��a<.�a<��a<F�a<Ǒa<@�a<Аa<S�a<׏a<v�a<��a<��a<$�a<��a<Y�a<��a<��a<H�a<ߋa<u�a<,�a<Ɋa<i�a<%�a<��a<k�a<"�a<��a<��a<6�a<��a<Ƈa<��a<G�a< �a<�a<��a<��a<s�a<^�a<D�a<�a<�a<�a<ۅa<څa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<�a<��a<�a<�  �  B�a<K�a<��a<��a<Ԇa<�a<�a<p�a<r�a<a<�a<�a<p�a<��a<��a<1�a<��a<ۉa<M�a<��a<��a<��a<��a<H�a<��a<�a<z�a<Ǎa<J�a<��a<:�a<{�a<�a<t�a<�a<}�a<͑a<r�a<֒a<w�a<�a<\�a<�a<f�a<�a<a�a<�a<h�a<��a<}�a<٘a<q�a<ʙa<R�a<Śa<H�a<śa<0�a<��a<�a<��a<�a<��a<�a<a�a<��a</�a<��a<�a<d�a<��a<�a<u�a<��a<�a<.�a<��a<ףa<�a<s�a<��a<��a<��a<S�a<�a<åa<��a<�a<X�a<P�a<��a<��a<Ŧa<�a<�a<�a<�a<H�a<O�a<v�a<��a<��a<ɧa<��a<��a<�a<�a<�a<�a<4�a<�a<$�a<�a<(�a<�a<�a<�a<�a<�a<Χa<֧a<ŧa<��a<��a<|�a<��a<Y�a<f�a<0�a<�a< �a<Ħa<Ȧa<q�a<c�a<(�a<��a<ۥa<��a<�a<=�a<2�a<�a<Ԥa<��a<j�a<_�a<��a<�a<��a<p�a<7�a<٢a<��a<B�a<2�a<��a<��a</�a<�a<��a<+�a<��a<��a<Y�a<�a<��a<=�a<ѝa<��a<�a<Ŝa<4�a<ޛa<p�a<ޚa<��a<�a<��a<�a<��a<+�a<��a<A�a<��a<d�a<ݕa<��a<�a<z�a<2�a<��a<9�a<��a<:�a<��a<A�a<�a<J�a<��a<\�a<�a<��a<"�a<ڍa<I�a<�a<��a<;�a<ыa<��a<.�a<��a<��a<�a<ۉa<l�a<�a<ӈa<k�a<B�a<�a<��a<n�a<G�a<�a<ކa<Άa<��a<��a<R�a<>�a<2�a< �a<
�a<ͅa<Ѕa<��a<��a<��a<��a<��a<��a<��a<��a<��a<ͅa<ׅa<�a<�a<�  �  H�a<e�a<��a<��a<݆a< �a<�a<M�a<s�a<��a<��a<�a<e�a<��a<��a<:�a<��a<��a<Q�a<��a<��a<f�a<��a<B�a<��a<�a<y�a<��a<Y�a<��a<.�a<~�a<�a<v�a<�a<o�a<בa<x�a<�a<d�a<��a<{�a<��a<�a<��a<k�a<�a<d�a<�a<g�a<ؘa<f�a<ۙa<O�a<Ěa<E�a<��a<4�a<��a<,�a<��a<�a<��a<��a<_�a<�a<@�a<��a<�a<u�a<ѡa<�a<e�a<��a<�a<5�a<��a<أa<�a<u�a<��a<�a<#�a<j�a<��a<ĥa<�a<�a<S�a<H�a<��a<��a<��a<�a<�a<�a<!�a<E�a<Y�a<n�a<��a<��a<��a<��a<�a<�a<�a<%�a<�a<.�a<+�a<.�a<(�a<,�a<�a<�a<�a<�a<�a<ڧa<ۧa<ӧa<��a<��a<��a<��a<t�a<b�a<.�a<&�a<��a<��a<��a<q�a<V�a<3�a<�a<Хa<��a<|�a<G�a<!�a<�a<ؤa<��a<i�a<A�a<�a<�a<��a<i�a<6�a<�a<��a<k�a<&�a<��a<��a<1�a<�a<��a<5�a<�a<��a<F�a<��a<��a<K�a<�a<��a<
�a<Üa<1�a<ʛa<Z�a<ݚa<|�a<�a<��a<
�a<��a<'�a<��a<<�a<ɖa<c�a<ܕa<k�a<��a<w�a<+�a<��a</�a<��a<K�a<בa<V�a<Րa<V�a<��a<d�a<�a<��a<"�a<܍a<O�a<	�a<��a<Q�a<�a<��a<%�a<ϊa<��a<��a<��a<c�a<�a<Ԉa<t�a<2�a<�a<��a<x�a<?�a<�a<�a<��a<��a<u�a<M�a<@�a<8�a< �a<�a<�a<څa<ǅa<a<��a<��a<��a<��a<��a<��a<ąa<ۅa<ԅa<�a<&�a<�  �  3�a<]�a<{�a<��a<͆a<��a<:�a<=�a<��a<��a<�a<�a<T�a<��a<�a<:�a<�a<�a<;�a<��a<�a<V�a<�a<)�a<��a<�a<b�a<؍a<?�a<��a< �a<��a<�a<��a<�a<b�a<�a<k�a<�a<p�a<�a<m�a<�a<k�a<�a<��a<�a<��a<��a<_�a<��a<H�a<ҙa<B�a<��a<1�a<��a<-�a<��a<(�a<��a<1�a<��a<	�a<��a<Пa<S�a<��a<�a<_�a<��a<�a<j�a<��a<�a<k�a<��a<�a<5�a<f�a<��a<�a<�a<K�a<��a<��a<�a<�a<2�a<��a<}�a<��a<ʦa<Ѧa<��a<��a<�a<7�a<N�a<a�a<��a<��a<��a<�a<ϧa<�a<
�a<�a<�a<�a<�a<�a<$�a<�a<�a<�a<�a<�a<اa<�a<�a<ӧa<ħa<��a<��a<z�a<k�a<L�a<<�a<�a<��a<�a<��a<��a<L�a<%�a<��a<��a<��a<r�a<G�a<�a<��a<¤a<��a<y�a<0�a<+�a<ѣa<��a<j�a< �a<�a<��a<i�a<�a<ڡa<��a<H�a<��a<��a<k�a<��a<��a<R�a<�a<��a<:�a<֝a<v�a< �a<��a<T�a<ٛa<R�a< �a<^�a<��a<x�a<�a<��a<�a<��a<,�a<Ŗa<E�a<��a<m�a<�a<��a<	�a<��a<$�a<��a<5�a<��a<K�a<ېa<f�a<�a<��a<�a<��a<G�a<͍a<h�a<��a<��a<2�a<׋a<r�a<!�a<Ίa<a�a<4�a<��a<n�a< �a<��a<}�a< �a<�a<��a<m�a<2�a<�a<�a<��a<��a<e�a<j�a<D�a<�a<�a<�a<݅a<ʅa<Åa<��a<��a<��a<��a<ǅa<��a<хa<Ʌa<܅a<�a<��a<"�a<�  �  O�a<m�a<��a<��a<Ɇa<�a<�a<<�a<r�a<��a<�a<"�a<i�a<��a<�a<3�a<��a<�a<A�a<��a<�a<O�a<Ƌa<'�a<��a<�a<��a<�a<R�a<��a<5�a<��a<�a<|�a<��a<n�a<�a<f�a<�a<y�a<��a<z�a<�a<~�a< �a<|�a<�a<l�a<�a<Q�a<֘a<Q�a<Ιa<P�a<͚a<;�a<��a<4�a<��a<"�a<��a<�a<y�a<�a<m�a<џa<K�a<��a<�a<y�a<ˡa<(�a<w�a<��a<��a<Q�a<��a<�a< �a<^�a<��a<�a<)�a<`�a<��a<ҥa<��a<�a<3�a<b�a<o�a<��a<��a<צa<��a<�a<�a<8�a<K�a<u�a<��a<��a<��a<��a<˧a<�a<��a<�a<!�a<,�a</�a<9�a<&�a<-�a<�a<�a<��a<�a<�a<�a<Χa<ϧa<��a<��a<��a<��a<{�a<a�a<?�a<�a<�a<Ʀa<��a<q�a<I�a<'�a<��a<ԥa<��a<p�a<@�a<"�a<��a<Ȥa<��a<\�a<)�a<
�a<ϣa<��a<v�a<>�a<��a<��a<n�a<-�a<ڡa<��a<7�a<�a<��a<Q�a<�a<��a<\�a<�a<��a<S�a<�a<��a<�a<��a<8�a<ěa<D�a<ۚa<g�a<��a<��a<�a<��a<�a<��a<=�a<��a<J�a<֕a<Z�a<�a<��a<
�a<��a<4�a<Œa<O�a<Бa<a�a<�a<d�a<�a<�a<
�a<��a<2�a<ōa<g�a<�a<��a<H�a<�a<��a<0�a<Ɗa<b�a<�a<��a<T�a<�a<Èa<y�a<4�a<�a<��a<i�a<F�a<�a<�a<��a<��a<a�a<N�a<1�a<�a<�a<�a<�a<�a<Ņa<ąa<��a<��a<��a<��a<��a<��a<��a<ׅa<�a<�a<%�a<�  �  L�a<n�a<��a<ȇa<��a<!�a</�a<��a<��a<׈a<
�a<@�a<��a<��a<<�a<M�a<��a<�a<i�a<��a<"�a<��a<ǌa<T�a<��a<�a<o�a<Ԏa<F�a<Əa<9�a<��a<0�a<��a<�a<o�a<�a<x�a<�a<^�a<��a<Z�a<ѕa<`�a<�a<`�a<�a<\�a<՘a<t�a<͙a<Q�a<��a<B�a<��a</�a<��a<�a<��a<�a<��a<��a<��a<ڟa<>�a<Ơa<�a<��a<ʡa<�a<~�a<�a</�a<��a<�a<�a<a�a<��a<��a<P�a<c�a<��a<�a<�a<A�a<~�a<Ħa<�a<�a<"�a<b�a<��a<��a<ħa<��a<��a<�a<<�a<.�a<D�a<c�a<o�a<��a<��a<Шa<��a<ڨa<��a<�a<��a<�a<�a<�a<�a<٨a<��a<�a<˨a<��a<��a<Ȩa<��a<~�a<��a<h�a<J�a<4�a<*�a<�a<��a<اa<��a<��a<Z�a<3�a<�a<Ӧa<��a<w�a<��a<�a<�a<��a<��a<y�a<Q�a<$�a<Τa<��a<��a<F�a<��a<��a<r�a<@�a<��a<��a<|�a<�a<��a<m�a<�a<ܠa<��a<�a<ڟa<d�a<��a<��a<]�a<�a<��a<�a<��a<[�a<ɛa<a�a<Ța<x�a<�a<��a< �a<��a<<�a<��a<Y�a<Ֆa<��a<��a<x�a<"�a<��a<-�a<��a<�a<��a<R�a<ґa<h�a<�a<��a<�a<��a<F�a<�a<a�a<�a<��a<>�a<֌a<��a<>�a<�a<��a<�a<��a<��a<1�a<��a<�a<g�a< �a<��a<��a<^�a<4�a<��a<�a<��a<��a<h�a<^�a<W�a<)�a<�a<��a<ކa<نa<�a<��a<݆a<نa<��a<��a<φa<��a<�a<��a<3�a<6�a<�  �  j�a<��a<��a<ʇa<݇a<�a<M�a<f�a<��a<шa<�a<H�a<��a<��a<�a<K�a<��a<�a<b�a<��a<�a<p�a<�a<>�a<��a<�a<��a<��a<_�a<Ǐa<,�a<��a<�a<w�a<�a<��a<��a<W�a<��a<m�a<�a<r�a< �a<w�a<�a<_�a<חa<a�a<Әa<F�a<��a<M�a<��a<9�a<��a<�a<��a<�a<��a<�a<��a<�a<Z�a<Οa<M�a<��a<�a<w�a<�a<N�a<��a<�a<9�a<��a<��a<$�a<w�a<��a<�a<+�a<��a<��a<�a<3�a<r�a<��a<��a<ܦa<�a<B�a<L�a<p�a<��a<��a<ǧa<�a<�a<�a<"�a<Q�a<c�a<~�a<��a<��a<��a<Ϩa<Өa<بa<�a<�a<�a<	�a<��a<��a<��a<�a<ɨa<�a<�a<٨a<��a<��a<��a<��a<r�a<i�a<S�a<)�a<�a<ߧa<ŧa<��a<x�a<T�a<-�a<�a<ۦa<��a<q�a<K�a<�a<�a<ϥa<��a<m�a<D�a<�a<�a<��a<l�a<C�a<�a<أa<��a<A�a<�a<��a<Y�a<�a<֡a<��a<0�a<��a<��a<*�a<ןa<}�a<-�a<Şa<R�a<�a<y�a<�a<��a<.�a<��a<]�a<�a<p�a<��a<y�a<�a<��a<,�a<��a<O�a<Öa<W�a<�a<��a< �a<��a< �a<��a<Q�a<Вa<V�a<ܑa<t�a<��a<��a<'�a<��a<4�a<Ўa<~�a<�a<��a<[�a<�a<��a<7�a<Ћa<{�a<8�a<ʊa<{�a<$�a<�a<��a<T�a< �a<ňa<��a<k�a<4�a<�a<߇a<��a<��a<�a<W�a<7�a<+�a<�a<�a<��a<�a<چa<҆a<φa<��a<߆a<�a<�a<Іa<��a<�a<%�a<A�a<�  �  P�a<v�a<��a<߇a<�a<�a<Y�a<j�a<��a<Ɉa<�a<=�a<��a<։a<�a<s�a<��a<�a<S�a<��a<4�a<t�a<��a<8�a<��a<#�a<v�a<��a<E�a<��a< �a<��a<�a<��a<�a<\�a<��a<]�a<�a<d�a<�a<]�a<ߕa<a�a<�a<��a<՗a<i�a<ߘa<[�a<�a<=�a<Śa<!�a<��a<+�a<��a<'�a<z�a<�a<r�a< �a<s�a<ԟa<T�a<��a<-�a<{�a<ҡa<,�a<��a<ޢa<+�a<��a<ƣa<'�a<O�a<��a<�a<0�a<��a<��a<�a<�a<S�a<��a<Ħa<�a<�a<K�a<O�a<��a<��a<��a<Чa<קa<�a<�a<8�a<Q�a<P�a<z�a<��a<èa<��a<ݨa<Ԩa<�a<�a<�a<�a<�a<�a<�a<��a<��a<̨a<�a<��a<˨a<��a<��a<��a<z�a<o�a<N�a<<�a<�a<'�a<�a<ħa<��a<}�a<y�a<%�a<�a<Цa<��a<��a<R�a<>�a<��a<ҥa<��a<r�a<d�a<�a< �a<��a<��a<N�a<��a<��a<p�a<:�a<�a<��a<^�a<�a<ǡa<Z�a</�a<��a<��a<!�a<ɟa<g�a<�a<��a<S�a<
�a<w�a<#�a<��a<B�a<ߛa<M�a<�a<W�a<�a<��a<�a<��a<�a<��a<:�a<�a<p�a<�a<��a<��a<��a<%�a<��a</�a<��a<H�a<ϑa<��a<�a<��a<��a<��a<@�a<Ԏa<��a<��a<��a<B�a<�a<��a<>�a<�a<t�a<A�a<͊a<��a<2�a<Չa<��a<C�a<'�a<шa<��a<k�a<!�a<�a<ԇa<ׇa<��a<��a<Y�a<?�a<I�a<�a<��a<�a<ۆa<Іa<نa<ֆa<��a<׆a<��a<�a<Ԇa<��a<�a<�a<=�a<�  �  j�a<��a<��a<��a<�a<�a<5�a<o�a<��a<Έa<�a<O�a<��a<ʉa<�a<b�a<��a<�a<i�a<��a<�a<y�a<ьa<N�a<��a<�a<��a<�a<_�a<̏a<A�a<��a<�a<��a<��a<��a<�a<p�a<�a<X�a<��a<p�a<�a<l�a<��a<Z�a<�a<\�a<͘a<N�a<řa<A�a<˚a<@�a<��a<$�a<��a<�a<��a<�a<z�a<�a<[�a<̟a<?�a<��a<�a<��a<ۡa<8�a<��a<��a<-�a<x�a<ףa<�a<m�a<��a<�a<2�a<W�a<��a<��a<0�a<Z�a<��a<��a<�a<�a<(�a<U�a<k�a<��a<��a<ԧa<�a<�a<�a</�a<J�a<k�a<��a<��a<��a<��a<��a<٨a<�a<�a<��a<��a<�a<��a<�a<Ԩa<�a<�a<Ѩa<רa<��a<��a<��a<x�a<��a<u�a<h�a<H�a<1�a<�a<�a<ѧa<��a<��a<Y�a<*�a<�a<�a<��a<��a<U�a<.�a<�a<٥a<��a<t�a<@�a<�a<ؤa<��a<{�a<<�a<�a<ãa<��a<E�a<�a<��a<^�a<�a<��a<�a< �a<Ӡa<t�a<�a<�a<z�a<�a<��a<`�a<�a<��a<�a<��a<5�a<��a<Q�a<�a<w�a<��a<��a<�a<��a<3�a<×a<A�a<ʖa<X�a<�a<y�a<�a<��a</�a<��a<;�a<˒a<_�a<Бa<Y�a<��a<��a<�a<��a<;�a<׎a<V�a<�a<��a<X�a<�a<��a<9�a<ڋa<��a<�a<ӊa<v�a<,�a<�a<��a<Y�a<�a<шa<��a<d�a<<�a<�a<ׇa<��a<��a<l�a<]�a<E�a<�a<�a<�a<��a<�a<�a<��a<Æa<Ɔa<a<چa<Іa<�a<�a<�a<4�a<D�a<�  �  n�a<n�a<��a<��a<�a<�a<G�a<��a<��a<�a<�a<L�a<��a<Ήa<'�a<^�a<Ɗa<��a<^�a<͋a<�a<��a<ڌa<T�a<��a<�a<��a<�a<\�a<��a<E�a<��a<$�a<p�a<�a<��a<Вa<w�a<�a<m�a<�a<Q�a<��a<X�a<��a<M�a<�a<Z�a<�a<c�a<Йa<]�a<��a<D�a<��a<2�a<��a<�a<��a<��a<��a<��a<n�a<��a<=�a<��a<��a<��a<ˡa<=�a<z�a<Ңa<A�a<x�a<ߣa< �a<n�a<��a<פa<F�a<`�a<åa<ǥa<"�a<Y�a<��a<��a<Цa<#�a<,�a<��a<q�a<��a<��a<��a<��a<��a<)�a<:�a<X�a<i�a<r�a<��a<��a<بa<Өa<بa<�a<ڨa<��a<�a<�a<Ϩa<��a<�a<�a<ߨa<��a<�a<��a<��a<��a<��a<��a<B�a<m�a<5�a<3�a<�a<�a<Χa<��a<��a<U�a<I�a<�a<ߦa<��a<��a<k�a<)�a<�a<ɥa<��a<��a<A�a<A�a<�a<��a<f�a<9�a<�a<��a<��a<�a<�a<��a<p�a<��a<��a<��a<�a<۠a<v�a<*�a<Ɵa<\�a<!�a<��a<d�a<՝a<��a<�a<Üa<J�a<̛a<m�a<Қa<z�a<��a<��a<�a<��a<;�a<��a<Z�a<ܖa<k�a<�a<w�a<�a<}�a<0�a<��a<@�a<��a<<�a<�a<Y�a<�a<g�a<�a<��a<%�a<�a<^�a< �a<��a<J�a<�a<��a<5�a<ċa<��a<"�a< �a<{�a<@�a<�a<��a<k�a<�a<�a<��a<r�a<:�a<��a<��a<��a<��a<��a<]�a<D�a<�a<�a<�a<�a<��a<چa<ʆa<ˆa<ņa<��a<�a<��a<܆a<��a<�a<.�a<�a<�  �  j�a<j�a<��a<؇a<��a<�a<I�a<i�a<��a<�a<�a<f�a<��a<Չa<!�a<l�a<��a<%�a<b�a<ˋa<�a<z�a<��a<H�a<��a<!�a<t�a<֎a<\�a<��a<(�a<��a<�a<�a<��a<Y�a<�a<g�a<ӓa<X�a<�a<c�a<�a<U�a<�a<o�a<�a<Y�a<�a<O�a<ݙa<P�a<˚a<E�a<��a<*�a<��a<*�a<��a<�a<��a<�a<`�a<�a<>�a<��a<�a<��a<ša<6�a<��a<�a<'�a<o�a<ʣa<�a<Q�a<��a<�a<,�a<_�a<��a<�a<&�a<O�a<}�a<Ǧa<�a<�a<0�a<[�a<v�a<��a<��a<�a<�a<�a<$�a<=�a<U�a<y�a<��a<��a<��a<��a<Ԩa<֨a<�a<��a<�a<�a<�a<�a<�a<�a<ըa<ۨa<Ԩa<��a<��a<��a<��a<��a<~�a<g�a<h�a<0�a<'�a< �a<��a<̧a<��a<|�a<\�a<B�a<�a<��a<��a<��a<e�a<8�a<�a<�a<��a<��a<K�a<�a<�a<��a<��a<M�a<��a<��a<��a<3�a<�a<��a<X�a<
�a<��a<W�a< �a<ʠa<e�a<�a<ɟa<m�a<�a<��a<W�a<��a<��a<�a<��a<6�a<ٛa<`�a<�a<|�a<�a<��a<�a<��a<5�a<ʗa<P�a<�a<]�a<��a<w�a<�a<��a<+�a<��a<9�a<��a<K�a<ˑa<O�a<�a<��a<�a<��a<9�a<юa<]�a<�a<��a<N�a<�a<��a<B�a<�a<��a<'�a<يa<��a<B�a<�a<��a<]�a<�a<݈a<��a<o�a<J�a<�a<�a<��a<��a<��a<[�a<K�a<;�a<�a<�a<��a<نa<цa<��a<��a<��a<Ɔa<��a<׆a<݆a<�a<��a<�a<6�a<�  �  C�a<��a<��a<��a<�a<�a<X�a<h�a<��a<ۈa<�a<]�a<��a<�a<�a<��a<��a<!�a<e�a<ʋa<3�a<w�a<��a<A�a<��a<
�a<�a<�a<:�a<ʏa<�a<��a<��a<q�a<��a<R�a<��a<D�a<�a<N�a<�a<b�a<ߕa<u�a<ݖa<`�a<�a<k�a<�a<R�a<�a<D�a<ߚa<;�a<ɛa<8�a<��a<;�a<��a<'�a<|�a<�a<h�a<�a<U�a<��a<�a<q�a<�a</�a<�a<�a<�a<��a<��a<�a<G�a<��a<�a<�a<q�a<��a<��a<�a<Z�a<��a<��a<�a<�a<M�a<Y�a<��a<��a<��a<�a<�a<,�a<�a<T�a<U�a<q�a<��a<��a<Ĩa<��a<ܨa<�a<ߨa<�a<�a<�a<�a<��a<�a<ۨa<�a<��a<ۨa<��a<Ĩa<��a<��a<��a<q�a<w�a<A�a<N�a<)�a<	�a<�a<֧a<��a<z�a<x�a<7�a<�a<�a<��a<��a<R�a<U�a<��a<�a<��a<��a<b�a<�a<��a<��a<w�a<5�a<�a<ţa<f�a<D�a<٢a<��a<J�a<��a<��a<P�a<(�a<��a<z�a<�a<˟a<l�a<�a<Þa<I�a<�a<��a<%�a<��a<:�a<�a<T�a<�a<q�a<�a<��a<�a<��a<&�a<חa<C�a<�a<d�a<��a<��a<
�a<��a<�a<��a<2�a<��a<Q�a<��a<e�a<ːa<��a<��a<��a<0�a<��a<p�a<��a<��a<5�a<�a<��a<.�a<֋a<~�a<C�a<׊a<��a<E�a<�a<��a<M�a<<�a<шa<��a<o�a<B�a<�a<�a<هa<��a<��a<h�a<>�a<'�a<�a<�a<چa<�a<Ɇa<��a<��a<��a<͆a<��a<܆a<Æa<�a<��a<�a<E�a<�  �  E�a<v�a<��a<͇a<�a<�a<;�a<��a<��a<�a<�a<\�a<��a<�a<�a<��a<ϊa<�a<k�a<ϋa<(�a<��a<׌a<K�a<��a<�a<q�a<�a<8�a<��a<#�a<��a<�a<n�a<�a<Y�a<ڒa<U�a<�a<U�a<��a<R�a<ߕa<W�a<�a<j�a<��a<X�a<�a<g�a<�a<W�a<ɚa<S�a<Λa<C�a<��a<9�a<��a<�a<��a<	�a<w�a<�a<;�a<��a<�a<|�a<ơa<0�a<t�a<ݢa<#�a<|�a<��a<
�a<E�a<��a<ڤa<!�a<]�a<��a<ߥa<
�a<X�a<|�a<æa<��a<�a<+�a<m�a<��a<��a<��a<֧a<�a<#�a<�a<V�a<e�a<{�a<��a<��a<��a<֨a<Ĩa<ڨa<��a<��a<�a<�a<�a<�a<�a<ըa<�a<¨a<��a<��a<��a<��a<��a<z�a<y�a<\�a<C�a<=�a<!�a<�a<�a<Чa<��a<��a<j�a<F�a<�a<�a<ɦa<��a<Y�a<N�a<�a<ߥa<��a<��a<X�a<0�a<ߤa<��a<��a<E�a<��a<��a<d�a<&�a<�a<��a<R�a<��a<��a<W�a<�a<��a<y�a<�a<şa<\�a<�a<��a<U�a<�a<��a<�a<��a<O�a<ߛa<g�a<�a<��a<�a<��a<$�a<��a<C�a<a<V�a<�a<t�a< �a<u�a<�a<��a<%�a<��a<3�a<��a<H�a<Ǒa<]�a<ڐa<p�a<�a<��a<)�a<Ǝa<\�a<��a<��a<2�a<�a<��a<=�a<�a<��a<"�a<�a<��a<E�a<��a<��a<q�a<3�a<؈a<��a<�a<L�a<�a<�a<ʇa<��a<s�a<_�a<U�a<2�a<�a<��a<܆a<φa<͆a<��a<ǆa<��a<��a<��a<��a<Ȇa<��a<�a<�a<+�a<�  �  s�a<t�a<��a<��a<�a<&�a<B�a<��a<��a<��a<!�a<s�a<��a<։a<P�a<d�a<׊a<'�a<y�a<֋a<
�a<��a<܌a<W�a<��a<�a<s�a<�a<[�a<��a<0�a<x�a<��a<p�a<�a<]�a<Ȓa<b�a<��a<Y�a<ܔa<P�a<�a<U�a<��a<K�a<�a<d�a<�a<a�a<ƙa<s�a<ʚa<l�a<��a<F�a<ɜa<!�a<��a<�a<��a<��a<i�a<�a<D�a<��a<��a<��a<ơa<J�a<}�a<Ӣa<+�a<W�a<ãa<��a<K�a<��a<֤a<�a<D�a<��a<ҥa<"�a<]�a<�a<æa<Ϧa<'�a<1�a<v�a<r�a<��a<Чa<�a<�a<�a<P�a<A�a<Z�a<��a<��a<��a<��a<֨a<Ψa<�a<�a<ڨa<��a<�a<�a<ڨa<�a<Ϩa<��a<Ҩa<��a<��a<��a<��a<��a<q�a<�a<S�a<q�a<:�a<%�a< �a<�a<ݧa<��a<��a<B�a<[�a<�a<�a<Ǧa<��a<��a<0�a<&�a<��a<��a<��a<:�a<=�a<�a<Ĥa<d�a<A�a<��a<��a<��a<�a<�a<��a<E�a<��a<��a<[�a<��a<Ša<O�a<�a<��a<Z�a</�a<��a<a�a<ӝa<��a<�a<��a<H�a<a<��a<�a<��a<�a<��a<9�a<��a<[�a<ȗa<p�a<֖a<f�a<�a<~�a<�a<|�a<1�a<��a<M�a<��a<>�a<Αa<8�a<�a<_�a<��a<��a<%�a<��a<C�a<�a<��a<J�a<�a<��a<=�a<Ëa<��a<'�a<�a<|�a<F�a<�a<��a<�a<�a<	�a<��a<s�a<d�a<�a<�a<��a<��a<~�a<k�a<>�a<�a<�a<�a<�a<Ća<цa<��a<��a<��a<��a<��a<��a<ӆa<ֆa<�a<�a<!�a<�  �  I�a<c�a<��a<Ǉa<�a<%�a<R�a<��a<��a<�a<�a<h�a<��a<�a<D�a<�a<Պa<!�a<b�a<�a<4�a<��a<�a<U�a<��a<�a<s�a<̎a<>�a<��a<�a<��a<��a<d�a<Ցa<O�a<͒a<O�a<ғa<O�a<Ȕa<G�a<ԕa<S�a<�a<d�a<�a<p�a<�a<t�a<��a<h�a<Śa<Y�a<ϛa<M�a<ʜa<;�a<��a<�a<��a<�a<��a<�a<Q�a<��a<�a<~�a<ȡa<�a<m�a<��a<�a<o�a<��a<��a<=�a<��a<Ϥa<�a<a�a<��a<ͥa<�a<=�a<��a<��a<ڦa<!�a<D�a<r�a<��a<§a<��a<�a<�a<"�a<J�a<Q�a<m�a<��a<x�a<��a<Ũa<֨a<٨a<�a<�a<�a<��a<ߨa<�a<ڨa<רa<ިa<ͨa<��a<��a<��a<��a<��a<��a<��a<c�a<W�a<H�a<*�a<'�a<�a<�a<ܧa<��a<��a<w�a<]�a<�a<��a<Ԧa<��a<��a<K�a<$�a<�a<��a<��a<d�a<8�a<��a<¤a<n�a<=�a<��a<��a<j�a<�a<Ѣa<��a<G�a<�a<��a<M�a<��a<��a<d�a<�a<��a<R�a<�a<��a<Y�a<�a<��a<*�a<��a<[�a<�a<x�a<�a<��a<�a<��a<:�a<��a<P�a<ȗa<^�a<��a<��a<�a<��a<�a<��a<(�a<��a< �a<��a<*�a<��a<O�a<ِa<^�a<�a<��a<�a<��a<_�a<�a<��a<4�a<ьa<��a<5�a<ϋa<��a<:�a<��a<��a<^�a<�a<��a<y�a<3�a<�a<��a<��a<T�a<�a<�a<ڇa<��a<��a<j�a<@�a<+�a<�a<�a<݆a<Ća<��a<��a<��a<��a<��a<��a<��a<ņa<݆a<��a<�a<%�a<�  �  E�a<��a<��a<Ǉa<�a<�a<G�a<u�a<��a<�a<>�a<m�a<��a<��a<�a<��a<��a<7�a<��a<ϋa<'�a<~�a<�a<E�a<͍a<	�a<s�a<�a<@�a<Əa<	�a<��a<ݐa<k�a<ݑa<R�a<�a<8�a<ϓa<=�a<Ҕa<j�a<Еa<r�a<Ӗa<u�a<�a<e�a<�a<_�a<�a<T�a<��a<T�a<כa<B�a<��a<D�a<��a<D�a<��a<�a<q�a<ޟa<I�a<��a<*�a<b�a<�a<�a<��a<Ԣa<�a<l�a<��a<
�a<E�a<��a<פa<��a<X�a<��a<�a<�a<S�a<��a<��a<�a<�a<8�a<]�a<��a<��a<Χa<�a<��a<3�a<$�a<^�a<g�a<��a<��a<��a<��a<��a<Шa<רa<��a<�a<ߨa<�a<�a<��a<Ѩa<Ȩa<èa<��a<èa<��a<��a<��a<z�a<s�a<^�a<x�a<C�a<P�a<�a<�a<�a<ɧa<��a<��a<q�a<B�a<8�a< �a<Ŧa<��a<_�a<_�a<�a<�a<̥a<��a<V�a<�a<�a<��a<��a<5�a<��a<ãa<k�a<?�a<̢a<��a<)�a<��a<��a<P�a<�a<��a<a�a<��a<��a<t�a<��a<��a<?�a<��a<��a< �a<��a<F�a<ޛa<d�a<�a<��a< �a<��a<!�a<Șa<B�a<��a<V�a<�a<m�a<��a<��a<�a<��a<�a<��a<#�a<��a<>�a<��a<M�a<��a<p�a<�a<��a<%�a<��a<W�a<�a<��a<=�a<�a<��a<%�a<��a<��a</�a<ۊa<��a<G�a< �a<Љa<e�a<C�a<݈a<ňa<��a<U�a<:�a<�a<чa<��a<�a<\�a<W�a<.�a< �a<�a<؆a<�a<��a<��a<��a<��a<��a<��a<��a<Æa<͆a<�a<��a<F�a<�  �  ?�a<}�a<��a<��a<�a<�a<`�a<��a<��a<�a<4�a<e�a<��a<	�a<N�a<��a<��a<0�a<��a<ڋa<2�a<��a<��a<H�a<��a<�a<q�a<ݎa<7�a<��a<�a<��a<�a<i�a<ʑa<E�a<��a<L�a<ēa<S�a<��a<K�a<͕a<k�a<ږa<]�a<�a<s�a<�a<x�a<�a<c�a<�a<O�a<̛a<[�a<՜a<>�a<��a<5�a<��a<�a<��a<��a<Y�a<��a<�a<i�a<ڡa<�a<o�a<��a<"�a<a�a<��a<�a<7�a<{�a<ˤa<�a<W�a<��a<ƥa<�a<G�a<��a<��a<�a<�a<Q�a<|�a<��a<��a<ԧa<��a<��a<5�a<U�a<l�a<\�a<�a<��a<��a<��a<ըa<�a<�a<�a<ިa<�a<��a<ݨa<ݨa<Шa<֨a<Ũa<èa<��a<��a<��a<��a<��a<}�a<a�a<R�a<=�a<C�a<�a<��a<��a<էa<ǧa<��a<t�a<M�a<.�a<��a<��a<��a<��a<d�a<�a<��a<ɥa<��a<b�a<:�a<�a<��a<{�a<1�a<��a<��a<c�a<�a<ۢa<��a<>�a<��a<��a<C�a<�a<��a<V�a<�a<��a<V�a<��a<��a<E�a<�a<��a<-�a<Ӝa<_�a<�a<s�a<�a<��a<�a<��a<E�a<Øa<:�a<�a<d�a<��a<��a<�a<��a<�a<��a<�a<��a<�a<��a<#�a<Ƒa<B�a<Ԑa<R�a<�a<x�a<�a<��a<U�a<��a<��a<+�a<یa<��a<&�a<׋a<��a<G�a<��a<��a<T�a<�a<ǉa<a�a<E�a<�a<ӈa<v�a<P�a<1�a<��a<Շa<��a<��a<h�a<J�a<�a<�a<�a<Ԇa<Ɔa<��a<��a<��a<��a<��a<��a<��a<Ɇa<Ԇa<�a<�a<!�a<�  �  X�a<]�a<��a<҇a<�a<�a<?�a<s�a<��a<��a<�a<��a<��a<�a<*�a<v�a<�a<9�a<g�a<�a<%�a<x�a<�a<S�a<��a<)�a<s�a<ʎa<]�a<��a<�a<s�a<��a<[�a<בa<p�a<��a<_�a<��a<a�a<Δa<e�a<�a<M�a<�a<j�a<�a<Y�a<Ϙa<X�a<�a<d�a<њa<t�a<ٛa<D�a<��a<A�a<ɝa<&�a<��a<�a<j�a<ʟa<=�a<��a<�a<��a<ša<,�a<��a<ʢa</�a<F�a<ţa<�a<U�a<��a<��a<�a<=�a<��a<ҥa</�a<B�a<�a<Ԧa<�a<�a<9�a<P�a<�a<��a<��a<��a<�a<�a<6�a<F�a<{�a<��a<��a<��a<��a<��a<Ũa<ըa<�a<��a<��a<Өa<��a<�a<ۨa<بa<��a<Ȩa<��a<Шa<��a<��a<x�a<x�a<j�a<]�a<W�a<#�a<0�a<�a<��a<ҧa<��a<��a<m�a<[�a<�a<�a<�a<��a<n�a<B�a<2�a<�a<��a<��a<U�a<�a<�a<��a<x�a<T�a<��a<��a<��a<�a<ܢa<|�a<A�a<�a<��a<n�a<�a<àa<@�a<�a<��a<o�a<�a<��a<[�a<�a<��a<�a<��a<@�a<�a<t�a<��a<��a<"�a<��a<0�a<Řa<c�a<֗a<^�a<�a<g�a<�a<w�a<�a<��a<0�a<��a</�a<Ȓa<4�a<ӑa<'�a<�a<H�a<�a<��a<	�a<��a<<�a<��a<��a<X�a<֌a<��a<N�a<׋a<��a</�a<Ίa<��a<Z�a<�a<Éa<��a<+�a<�a<��a<��a<r�a<�a<�a<Ӈa<��a<u�a<Y�a<K�a<5�a<�a<܆a<�a<ӆa<��a<��a<��a<��a<��a<҆a<��a<Ɔa<ˆa<�a<
�a<+�a<�  �  ?�a<}�a<��a<��a<�a<�a<`�a<��a<��a<�a<4�a<e�a<��a<	�a<N�a<��a<��a<0�a<��a<ڋa<2�a<��a<��a<H�a<��a<�a<q�a<ݎa<7�a<��a<�a<��a<�a<i�a<ʑa<E�a<��a<L�a<ēa<S�a<��a<K�a<͕a<k�a<ږa<]�a<�a<s�a<�a<x�a<�a<c�a<�a<O�a<̛a<[�a<՜a<>�a<��a<5�a<��a<�a<��a<��a<Y�a<��a<�a<i�a<ڡa<�a<o�a<��a<"�a<a�a<��a<�a<7�a<{�a<ˤa<�a<W�a<��a<ƥa<�a<G�a<��a<��a<�a<�a<Q�a<|�a<��a<��a<ԧa<��a<��a<5�a<U�a<l�a<\�a<�a<��a<��a<��a<ըa<�a<�a<�a<ިa<�a<��a<ݨa<ݨa<Шa<֨a<Ũa<èa<��a<��a<��a<��a<��a<}�a<a�a<R�a<=�a<C�a<�a<��a<��a<էa<ǧa<��a<t�a<M�a<.�a<��a<��a<��a<��a<d�a<�a<��a<ɥa<��a<b�a<:�a<�a<��a<{�a<1�a<��a<��a<c�a<�a<ۢa<��a<>�a<��a<��a<C�a<�a<��a<V�a<�a<��a<V�a<��a<��a<E�a<�a<��a<-�a<Ӝa<_�a<�a<s�a<�a<��a<�a<��a<E�a<Øa<:�a<�a<d�a<��a<��a<�a<��a<�a<��a<�a<��a<�a<��a<#�a<Ƒa<B�a<Ԑa<R�a<�a<x�a<�a<��a<U�a<��a<��a<+�a<یa<��a<&�a<׋a<��a<G�a<��a<��a<T�a<�a<ǉa<a�a<E�a<�a<ӈa<v�a<P�a<1�a<��a<Շa<��a<��a<h�a<J�a<�a<�a<�a<Ԇa<Ɔa<��a<��a<��a<��a<��a<��a<��a<Ɇa<Ԇa<�a<�a<!�a<�  �  E�a<��a<��a<Ǉa<�a<�a<G�a<u�a<��a<�a<>�a<m�a<��a<��a<�a<��a<��a<7�a<��a<ϋa<'�a<~�a<�a<E�a<͍a<	�a<s�a<�a<@�a<Əa<	�a<��a<ݐa<k�a<ݑa<R�a<�a<8�a<ϓa<=�a<Ҕa<j�a<Еa<r�a<Ӗa<u�a<�a<e�a<�a<_�a<�a<T�a<��a<T�a<כa<B�a<��a<D�a<��a<D�a<��a<�a<q�a<ޟa<I�a<��a<*�a<b�a<�a<�a<��a<Ԣa<�a<l�a<��a<
�a<E�a<��a<פa<��a<X�a<��a<�a<�a<S�a<��a<��a<�a<�a<8�a<]�a<��a<��a<Χa<�a<��a<3�a<$�a<^�a<g�a<��a<��a<��a<��a<��a<Шa<רa<��a<�a<ߨa<�a<�a<��a<Ѩa<Ȩa<èa<��a<èa<��a<��a<��a<z�a<s�a<^�a<x�a<C�a<P�a<�a<�a<�a<ɧa<��a<��a<q�a<B�a<8�a< �a<Ŧa<��a<_�a<_�a<�a<�a<̥a<��a<V�a<�a<�a<��a<��a<5�a<��a<ãa<k�a<?�a<̢a<��a<)�a<��a<��a<P�a<�a<��a<a�a<��a<��a<t�a<��a<��a<?�a<��a<��a< �a<��a<F�a<ޛa<d�a<�a<��a< �a<��a<!�a<Șa<B�a<��a<V�a<�a<m�a<��a<��a<�a<��a<�a<��a<#�a<��a<>�a<��a<M�a<��a<p�a<�a<��a<%�a<��a<W�a<�a<��a<=�a<�a<��a<%�a<��a<��a</�a<ۊa<��a<G�a< �a<Љa<e�a<C�a<݈a<ňa<��a<U�a<:�a<�a<чa<��a<�a<\�a<W�a<.�a< �a<�a<؆a<�a<��a<��a<��a<��a<��a<��a<��a<Æa<͆a<�a<��a<F�a<�  �  I�a<c�a<��a<Ǉa<�a<%�a<R�a<��a<��a<�a<�a<h�a<��a<�a<D�a<�a<Պa<!�a<b�a<�a<4�a<��a<�a<U�a<��a<�a<s�a<̎a<>�a<��a<�a<��a<��a<d�a<Ցa<O�a<͒a<O�a<ғa<O�a<Ȕa<G�a<ԕa<S�a<�a<d�a<�a<p�a<�a<t�a<��a<h�a<Śa<Y�a<ϛa<M�a<ʜa<;�a<��a<�a<��a<�a<��a<�a<Q�a<��a<�a<~�a<ȡa<�a<m�a<��a<�a<o�a<��a<��a<=�a<��a<Ϥa<�a<a�a<��a<ͥa<�a<=�a<��a<��a<ڦa<!�a<D�a<r�a<��a<§a<��a<�a<�a<"�a<J�a<Q�a<m�a<��a<x�a<��a<Ũa<֨a<٨a<�a<�a<�a<��a<ߨa<�a<ڨa<רa<ިa<ͨa<��a<��a<��a<��a<��a<��a<��a<c�a<W�a<H�a<*�a<'�a<�a<�a<ܧa<��a<��a<w�a<]�a<�a<��a<Ԧa<��a<��a<K�a<$�a<�a<��a<��a<d�a<8�a<��a<¤a<n�a<=�a<��a<��a<j�a<�a<Ѣa<��a<G�a<�a<��a<M�a<��a<��a<d�a<�a<��a<R�a<�a<��a<Y�a<�a<��a<*�a<��a<[�a<�a<x�a<�a<��a<�a<��a<:�a<��a<P�a<ȗa<^�a<��a<��a<�a<��a<�a<��a<(�a<��a< �a<��a<*�a<��a<O�a<ِa<^�a<�a<��a<�a<��a<_�a<�a<��a<4�a<ьa<��a<5�a<ϋa<��a<:�a<��a<��a<^�a<�a<��a<y�a<3�a<�a<��a<��a<T�a<�a<�a<ڇa<��a<��a<j�a<@�a<+�a<�a<�a<݆a<Ća<��a<��a<��a<��a<��a<��a<��a<ņa<݆a<��a<�a<%�a<�  �  s�a<t�a<��a<��a<�a<&�a<B�a<��a<��a<��a<!�a<s�a<��a<։a<P�a<d�a<׊a<'�a<y�a<֋a<
�a<��a<܌a<W�a<��a<�a<s�a<�a<[�a<��a<0�a<x�a<��a<p�a<�a<]�a<Ȓa<b�a<��a<Y�a<ܔa<P�a<�a<U�a<��a<K�a<�a<d�a<�a<a�a<ƙa<s�a<ʚa<l�a<��a<F�a<ɜa<!�a<��a<�a<��a<��a<i�a<�a<D�a<��a<��a<��a<ơa<J�a<}�a<Ӣa<+�a<W�a<ãa<��a<K�a<��a<֤a<�a<D�a<��a<ҥa<"�a<]�a<�a<æa<Ϧa<'�a<1�a<v�a<r�a<��a<Чa<�a<�a<�a<P�a<A�a<Z�a<��a<��a<��a<��a<֨a<Ψa<�a<�a<ڨa<��a<�a<�a<ڨa<�a<Ϩa<��a<Ҩa<��a<��a<��a<��a<��a<q�a<�a<S�a<q�a<:�a<%�a< �a<�a<ݧa<��a<��a<B�a<[�a<�a<�a<Ǧa<��a<��a<0�a<&�a<��a<��a<��a<:�a<=�a<�a<Ĥa<d�a<A�a<��a<��a<��a<�a<�a<��a<E�a<��a<��a<[�a<��a<Ša<O�a<�a<��a<Z�a</�a<��a<a�a<ӝa<��a<�a<��a<H�a<a<��a<�a<��a<�a<��a<9�a<��a<[�a<ȗa<p�a<֖a<f�a<�a<~�a<�a<|�a<1�a<��a<M�a<��a<>�a<Αa<8�a<�a<_�a<��a<��a<%�a<��a<C�a<�a<��a<J�a<�a<��a<=�a<Ëa<��a<'�a<�a<|�a<F�a<�a<��a<�a<�a<	�a<��a<s�a<d�a<�a<�a<��a<��a<~�a<k�a<>�a<�a<�a<�a<�a<Ća<цa<��a<��a<��a<��a<��a<��a<ӆa<ֆa<�a<�a<!�a<�  �  E�a<v�a<��a<͇a<�a<�a<;�a<��a<��a<�a<�a<\�a<��a<�a<�a<��a<ϊa<�a<k�a<ϋa<(�a<��a<׌a<K�a<��a<�a<q�a<�a<8�a<��a<#�a<��a<�a<n�a<�a<Y�a<ڒa<U�a<�a<U�a<��a<R�a<ߕa<W�a<�a<j�a<��a<X�a<�a<g�a<�a<W�a<ɚa<S�a<Λa<C�a<��a<9�a<��a<�a<��a<	�a<w�a<�a<;�a<��a<�a<|�a<ơa<0�a<t�a<ݢa<#�a<|�a<��a<
�a<E�a<��a<ڤa<!�a<]�a<��a<ߥa<
�a<X�a<|�a<æa<��a<�a<+�a<m�a<��a<��a<��a<֧a<�a<#�a<�a<V�a<e�a<{�a<��a<��a<��a<֨a<Ĩa<ڨa<��a<��a<�a<�a<�a<�a<�a<ըa<�a<¨a<��a<��a<��a<��a<��a<z�a<y�a<\�a<C�a<=�a<!�a<�a<�a<Чa<��a<��a<j�a<F�a<�a<�a<ɦa<��a<Y�a<N�a<�a<ߥa<��a<��a<X�a<0�a<ߤa<��a<��a<E�a<��a<��a<d�a<&�a<�a<��a<R�a<��a<��a<W�a<�a<��a<y�a<�a<şa<\�a<�a<��a<U�a<�a<��a<�a<��a<O�a<ߛa<g�a<�a<��a<�a<��a<$�a<��a<C�a<a<V�a<�a<t�a< �a<u�a<�a<��a<%�a<��a<3�a<��a<H�a<Ǒa<]�a<ڐa<p�a<�a<��a<)�a<Ǝa<\�a<��a<��a<2�a<�a<��a<=�a<�a<��a<"�a<�a<��a<E�a<��a<��a<q�a<3�a<؈a<��a<�a<L�a<�a<�a<ʇa<��a<s�a<_�a<U�a<2�a<�a<��a<܆a<φa<͆a<��a<ǆa<��a<��a<��a<��a<Ȇa<��a<�a<�a<+�a<�  �  C�a<��a<��a<��a<�a<�a<X�a<h�a<��a<ۈa<�a<]�a<��a<�a<�a<��a<��a<!�a<e�a<ʋa<3�a<w�a<��a<A�a<��a<
�a<�a<�a<:�a<ʏa<�a<��a<��a<q�a<��a<R�a<��a<D�a<�a<N�a<�a<b�a<ߕa<u�a<ݖa<`�a<�a<k�a<�a<R�a<�a<D�a<ߚa<;�a<ɛa<8�a<��a<;�a<��a<'�a<|�a<�a<h�a<�a<U�a<��a<�a<q�a<�a</�a<�a<�a<�a<��a<��a<�a<G�a<��a<�a<�a<q�a<��a<��a<�a<Z�a<��a<��a<�a<�a<M�a<Y�a<��a<��a<��a<�a<�a<,�a<�a<T�a<U�a<q�a<��a<��a<Ĩa<��a<ܨa<�a<ߨa<�a<�a<�a<�a<��a<�a<ۨa<�a<��a<ۨa<��a<Ĩa<��a<��a<��a<q�a<w�a<A�a<N�a<)�a<	�a<�a<֧a<��a<z�a<x�a<7�a<�a<�a<��a<��a<R�a<U�a<��a<�a<��a<��a<b�a<�a<��a<��a<w�a<5�a<�a<ţa<f�a<D�a<٢a<��a<J�a<��a<��a<P�a<(�a<��a<z�a<�a<˟a<l�a<�a<Þa<I�a<�a<��a<%�a<��a<:�a<�a<T�a<�a<q�a<�a<��a<�a<��a<&�a<חa<C�a<�a<d�a<��a<��a<
�a<��a<�a<��a<2�a<��a<Q�a<��a<e�a<ːa<��a<��a<��a<0�a<��a<p�a<��a<��a<5�a<�a<��a<.�a<֋a<~�a<C�a<׊a<��a<E�a<�a<��a<M�a<<�a<шa<��a<o�a<B�a<�a<�a<هa<��a<��a<h�a<>�a<'�a<�a<�a<چa<�a<Ɇa<��a<��a<��a<͆a<��a<܆a<Æa<�a<��a<�a<E�a<�  �  j�a<j�a<��a<؇a<��a<�a<I�a<i�a<��a<�a<�a<f�a<��a<Չa<!�a<l�a<��a<%�a<b�a<ˋa<�a<z�a<��a<H�a<��a<!�a<t�a<֎a<\�a<��a<(�a<��a<�a<�a<��a<Y�a<�a<g�a<ӓa<X�a<�a<c�a<�a<U�a<�a<o�a<�a<Y�a<�a<O�a<ݙa<P�a<˚a<E�a<��a<*�a<��a<*�a<��a<�a<��a<�a<`�a<�a<>�a<��a<�a<��a<ša<6�a<��a<�a<'�a<o�a<ʣa<�a<Q�a<��a<�a<,�a<_�a<��a<�a<&�a<O�a<}�a<Ǧa<�a<�a<0�a<[�a<v�a<��a<��a<�a<�a<�a<$�a<=�a<U�a<y�a<��a<��a<��a<��a<Ԩa<֨a<�a<��a<�a<�a<�a<�a<�a<�a<ըa<ۨa<Ԩa<��a<��a<��a<��a<��a<~�a<g�a<h�a<0�a<'�a< �a<��a<̧a<��a<|�a<\�a<B�a<�a<��a<��a<��a<e�a<8�a<�a<�a<��a<��a<K�a<�a<�a<��a<��a<M�a<��a<��a<��a<3�a<�a<��a<X�a<
�a<��a<W�a< �a<ʠa<e�a<�a<ɟa<m�a<�a<��a<W�a<��a<��a<�a<��a<6�a<ٛa<`�a<�a<|�a<�a<��a<�a<��a<5�a<ʗa<P�a<�a<]�a<��a<w�a<�a<��a<+�a<��a<9�a<��a<K�a<ˑa<O�a<�a<��a<�a<��a<9�a<юa<]�a<�a<��a<N�a<�a<��a<B�a<�a<��a<'�a<يa<��a<B�a<�a<��a<]�a<�a<݈a<��a<o�a<J�a<�a<�a<��a<��a<��a<[�a<K�a<;�a<�a<�a<��a<نa<цa<��a<��a<��a<Ɔa<��a<׆a<݆a<�a<��a<�a<6�a<�  �  n�a<n�a<��a<��a<�a<�a<G�a<��a<��a<�a<�a<L�a<��a<Ήa<'�a<^�a<Ɗa<��a<^�a<͋a<�a<��a<ڌa<T�a<��a<�a<��a<�a<\�a<��a<E�a<��a<$�a<p�a<�a<��a<Вa<w�a<�a<m�a<�a<Q�a<��a<X�a<��a<M�a<�a<Z�a<�a<c�a<Йa<]�a<��a<D�a<��a<2�a<��a<�a<��a<��a<��a<��a<n�a<��a<=�a<��a<��a<��a<ˡa<=�a<z�a<Ңa<A�a<x�a<ߣa< �a<n�a<��a<פa<F�a<`�a<åa<ǥa<"�a<Y�a<��a<��a<Цa<#�a<,�a<��a<q�a<��a<��a<��a<��a<��a<)�a<:�a<X�a<i�a<r�a<��a<��a<بa<Өa<بa<�a<ڨa<��a<�a<�a<Ϩa<��a<�a<�a<ߨa<��a<�a<��a<��a<��a<��a<��a<B�a<m�a<5�a<3�a<�a<�a<Χa<��a<��a<U�a<I�a<�a<ߦa<��a<��a<k�a<)�a<�a<ɥa<��a<��a<A�a<A�a<�a<��a<f�a<9�a<�a<��a<��a<�a<�a<��a<p�a<��a<��a<��a<�a<۠a<v�a<*�a<Ɵa<\�a<!�a<��a<d�a<՝a<��a<�a<Üa<J�a<̛a<m�a<Қa<z�a<��a<��a<�a<��a<;�a<��a<Z�a<ܖa<k�a<�a<w�a<�a<}�a<0�a<��a<@�a<��a<<�a<�a<Y�a<�a<g�a<�a<��a<%�a<�a<^�a< �a<��a<J�a<�a<��a<5�a<ċa<��a<"�a< �a<{�a<@�a<�a<��a<k�a<�a<�a<��a<r�a<:�a<��a<��a<��a<��a<��a<]�a<D�a<�a<�a<�a<�a<��a<چa<ʆa<ˆa<ņa<��a<�a<��a<܆a<��a<�a<.�a<�a<�  �  j�a<��a<��a<��a<�a<�a<5�a<o�a<��a<Έa<�a<O�a<��a<ʉa<�a<b�a<��a<�a<i�a<��a<�a<y�a<ьa<N�a<��a<�a<��a<�a<_�a<̏a<A�a<��a<�a<��a<��a<��a<�a<p�a<�a<X�a<��a<p�a<�a<l�a<��a<Z�a<�a<\�a<͘a<N�a<řa<A�a<˚a<@�a<��a<$�a<��a<�a<��a<�a<z�a<�a<[�a<̟a<?�a<��a<�a<��a<ۡa<8�a<��a<��a<-�a<x�a<ףa<�a<m�a<��a<�a<2�a<W�a<��a<��a<0�a<Z�a<��a<��a<�a<�a<(�a<U�a<k�a<��a<��a<ԧa<�a<�a<�a</�a<J�a<k�a<��a<��a<��a<��a<��a<٨a<�a<�a<��a<��a<�a<��a<�a<Ԩa<�a<�a<Ѩa<רa<��a<��a<��a<x�a<��a<u�a<h�a<H�a<1�a<�a<�a<ѧa<��a<��a<Y�a<*�a<�a<�a<��a<��a<U�a<.�a<�a<٥a<��a<t�a<@�a<�a<ؤa<��a<{�a<<�a<�a<ãa<��a<E�a<�a<��a<^�a<�a<��a<�a< �a<Ӡa<t�a<�a<�a<z�a<�a<��a<`�a<�a<��a<�a<��a<5�a<��a<Q�a<�a<w�a<��a<��a<�a<��a<3�a<×a<A�a<ʖa<X�a<�a<y�a<�a<��a</�a<��a<;�a<˒a<_�a<Бa<Y�a<��a<��a<�a<��a<;�a<׎a<V�a<�a<��a<X�a<�a<��a<9�a<ڋa<��a<�a<ӊa<v�a<,�a<�a<��a<Y�a<�a<шa<��a<d�a<<�a<�a<ׇa<��a<��a<l�a<]�a<E�a<�a<�a<�a<��a<�a<�a<��a<Æa<Ɔa<a<چa<Іa<�a<�a<�a<4�a<D�a<�  �  P�a<v�a<��a<߇a<�a<�a<Y�a<j�a<��a<Ɉa<�a<=�a<��a<։a<�a<s�a<��a<�a<S�a<��a<4�a<t�a<��a<8�a<��a<#�a<v�a<��a<E�a<��a< �a<��a<�a<��a<�a<\�a<��a<]�a<�a<d�a<�a<]�a<ߕa<a�a<�a<��a<՗a<i�a<ߘa<[�a<�a<=�a<Śa<!�a<��a<+�a<��a<'�a<z�a<�a<r�a< �a<s�a<ԟa<T�a<��a<-�a<{�a<ҡa<,�a<��a<ޢa<+�a<��a<ƣa<'�a<O�a<��a<�a<0�a<��a<��a<�a<�a<S�a<��a<Ħa<�a<�a<K�a<O�a<��a<��a<��a<Чa<קa<�a<�a<8�a<Q�a<P�a<z�a<��a<èa<��a<ݨa<Ԩa<�a<�a<�a<�a<�a<�a<�a<��a<��a<̨a<�a<��a<˨a<��a<��a<��a<z�a<o�a<N�a<<�a<�a<'�a<�a<ħa<��a<}�a<y�a<%�a<�a<Цa<��a<��a<R�a<>�a<��a<ҥa<��a<r�a<d�a<�a< �a<��a<��a<N�a<��a<��a<p�a<:�a<�a<��a<^�a<�a<ǡa<Z�a</�a<��a<��a<!�a<ɟa<g�a<�a<��a<S�a<
�a<w�a<#�a<��a<B�a<ߛa<M�a<�a<W�a<�a<��a<�a<��a<�a<��a<:�a<�a<p�a<�a<��a<��a<��a<%�a<��a</�a<��a<H�a<ϑa<��a<�a<��a<��a<��a<@�a<Ԏa<��a<��a<��a<B�a<�a<��a<>�a<�a<t�a<A�a<͊a<��a<2�a<Չa<��a<C�a<'�a<шa<��a<k�a<!�a<�a<ԇa<ׇa<��a<��a<Y�a<?�a<I�a<�a<��a<�a<ۆa<Іa<نa<ֆa<��a<׆a<��a<�a<Ԇa<��a<�a<�a<=�a<�  �  j�a<��a<��a<ʇa<݇a<�a<M�a<f�a<��a<шa<�a<H�a<��a<��a<�a<K�a<��a<�a<b�a<��a<�a<p�a<�a<>�a<��a<�a<��a<��a<_�a<Ǐa<,�a<��a<�a<w�a<�a<��a<��a<W�a<��a<m�a<�a<r�a< �a<w�a<�a<_�a<חa<a�a<Әa<F�a<��a<M�a<��a<9�a<��a<�a<��a<�a<��a<�a<��a<�a<Z�a<Οa<M�a<��a<�a<w�a<�a<N�a<��a<�a<9�a<��a<��a<$�a<w�a<��a<�a<+�a<��a<��a<�a<3�a<r�a<��a<��a<ܦa<�a<B�a<L�a<p�a<��a<��a<ǧa<�a<�a<�a<"�a<Q�a<c�a<~�a<��a<��a<��a<Ϩa<Өa<بa<�a<�a<�a<	�a<��a<��a<��a<�a<ɨa<�a<�a<٨a<��a<��a<��a<��a<r�a<i�a<S�a<)�a<�a<ߧa<ŧa<��a<x�a<T�a<-�a<�a<ۦa<��a<q�a<K�a<�a<�a<ϥa<��a<m�a<D�a<�a<�a<��a<l�a<C�a<�a<أa<��a<A�a<�a<��a<Y�a<�a<֡a<��a<0�a<��a<��a<*�a<ןa<}�a<-�a<Şa<R�a<�a<y�a<�a<��a<.�a<��a<]�a<�a<p�a<��a<y�a<�a<��a<,�a<��a<O�a<Öa<W�a<�a<��a< �a<��a< �a<��a<Q�a<Вa<V�a<ܑa<t�a<��a<��a<'�a<��a<4�a<Ўa<~�a<�a<��a<[�a<�a<��a<7�a<Ћa<{�a<8�a<ʊa<{�a<$�a<�a<��a<T�a< �a<ňa<��a<k�a<4�a<�a<߇a<��a<��a<�a<W�a<7�a<+�a<�a<�a<��a<�a<چa<҆a<φa<��a<߆a<�a<�a<Іa<��a<�a<%�a<A�a<�  �  m�a<~�a<̈a<ڈa<��a<$�a<8�a<��a<��a<�a<�a<]�a<��a<Պa<P�a<U�a<ۋa<�a<p�a<��a<!�a<��a<ύa<F�a<��a<(�a<��a<�a<J�a<��a<G�a<��a<�a<��a<ݒa<N�a<ߓa<u�a<єa<k�a<ݕa<Q�a<ϖa<@�a<�a<A�a<Řa<2�a<��a<@�a<��a<(�a<}�a</�a<�a<�a<��a<ڝa<��a<��a<U�a<��a<>�a<��a<��a<q�a<Сa<`�a<��a<��a<N�a<��a<�a<;�a<��a<ܤa<�a<W�a<��a<�a<&�a<��a<��a<�a<�a<U�a<��a<��a<ѧa<�a<$�a<E�a<X�a<��a<��a<רa<��a<�a<�a<�a<=�a<6�a<`�a<v�a<��a<z�a<��a<��a<��a<�a<��a<��a<��a<Щa<��a<��a<��a<��a<w�a<t�a<��a<s�a<[�a<g�a<2�a<'�a<�a<�a<ߨa<��a<��a<]�a<]�a<0�a<�a<˧a<��a<��a<O�a<W�a<�a<�a<��a<}�a<C�a<�a<�a<��a<{�a<9�a<�a<ۤa<��a<C�a<��a<ڣa<h�a<4�a<�a<x�a<#�a<�a<��a<?�a<�a<��a<=�a<��a<s�a<E�a<��a<T�a<ܝa<l�a<�a<��a<3�a<��a<e�a<˚a<|�a<�a<j�a<,�a<y�a<1�a<��a<T�a<̖a<O�a<�a<t�a<0�a<��a<&�a<��a<A�a<�a<M�a<��a<v�a<�a<��a<C�a<�a<^�a<)�a<��a<D�a<��a<��a<S�a<Ռa<��a<�a<�a<��a<5�a<��a<��a<��a<�a<�a<��a<u�a<S�a<�a<�a<Јa<��a<o�a<g�a<N�a<9�a<H�a<��a<��a<�a<��a<�a<ԇa<�a<͇a<��a<҇a<�a<�a<�a<K�a<E�a<�  �  y�a<��a<��a<Ĉa< �a<4�a<_�a<u�a<��a<�a<+�a<Q�a<��a<ӊa<�a<d�a<ŋa<�a<{�a<��a<�a<z�a<�a<S�a<��a<�a<r�a<�a<Z�a<Đa<&�a<��a<�a<�a<�a<}�a<��a<Y�a<֔a<I�a<ѕa<Z�a<ܖa<M�a<��a<A�a<ɘa<P�a<��a<-�a<��a<-�a<��a<�a<��a<�a<h�a<�a<h�a<ޞa<Z�a<��a<-�a<��a<�a<~�a<١a<0�a<��a<�a<V�a<��a<�a<D�a<��a<�a<>�a<��a<��a<�a<3�a<m�a<��a<�a<)�a<D�a<m�a<��a<ߧa<�a<�a<>�a<S�a<��a<��a<��a<��a<ިa<��a<�a<(�a<T�a<`�a<e�a<x�a<��a<��a<��a<��a<��a<ȩa<ѩa<Ωa<��a<��a<��a<��a<��a<��a<��a<z�a<o�a<\�a<K�a<G�a<4�a<�a<�a<ɨa<��a<��a<��a<G�a<#�a<�a<�a<��a<��a<L�a<%�a<�a<צa<��a<��a<A�a<�a<ߥa<��a<��a<H�a<��a<¤a<��a<S�a<�a<��a<s�a< �a<ݢa<��a<Q�a<��a<��a<D�a<�a<��a<F�a<�a<��a<�a<��a<Y�a<��a<��a<	�a<��a<7�a<ěa<I�a<Κa<P�a<�a<t�a<�a<��a<6�a<��a<C�a<Ֆa<t�a<��a<~�a<��a<��a<1�a<��a<>�a<��a<V�a<�a<��a<#�a<��a<<�a<ȏa<l�a<�a<��a<S�a<��a<��a<&�a<�a<��a<>�a<؋a<��a<0�a< �a<��a<i�a<�a<ۉa<��a<s�a<=�a<&�a<�a<��a<��a<��a<~�a<V�a<(�a<�a<�a<�a<��a<�a<ڇa<Շa<҇a<��a<��a<��a<�a<�a<�a<0�a<Y�a<�  �  ^�a<��a<��a<وa<�a<�a<W�a<r�a<ɉa<։a<)�a<K�a<��a<�a<!�a<��a<��a<�a<i�a<��a<?�a<q�a<�a<0�a<Îa<�a<�a<��a<C�a<̐a<�a<��a<
�a<~�a<�a<B�a<�a<K�a<��a<I�a<ܕa<M�a<ɖa<`�a<��a<a�a<��a<:�a<��a<B�a<��a<�a<��a<��a<��a<�a<��a<�a<K�a<�a<@�a<ɟa<K�a<��a<	�a<f�a<�a<,�a<��a<��a<F�a<��a<�a<f�a<��a<�a<	�a<e�a<��a<�a<T�a<Y�a<��a<٦a< �a<X�a<r�a<ŧa<��a<��a<�a<^�a<]�a<v�a<��a<��a<�a<�a<�a<'�a<�a<X�a<K�a<��a<{�a<��a<��a<��a<éa<��a<שa<��a<ʩa<��a<��a<ȩa<��a<��a<h�a<��a<w�a<~�a<h�a<=�a<H�a<�a<!�a<�a<ިa<Ȩa<��a<}�a<C�a<B�a<�a<�a<��a<��a<n�a<'�a<�a<Ŧa<��a<u�a<A�a<5�a<եa<��a<e�a<[�a<�a<Ϥa<��a<<�a<�a<��a<��a<(�a<ܢa<��a<�a<�a<��a<e�a<�a<��a<9�a<ڟa<��a<�a<Ӟa<K�a<�a<~�a<�a<��a<�a<̛a<.�a<�a<p�a<��a<��a<�a<��a<�a<a<a�a<Ζa<b�a<�a<��a<��a<��a<!�a<��a<I�a<��a<x�a<בa<��a<�a<��a<>�a<ʏa<��a<�a<��a<>�a<�a<��a<+�a<��a<q�a<1�a<΋a<��a<;�a<�a<��a<Q�a<D�a<�a<a<��a<3�a<*�a<߈a<߈a<��a<��a<[�a<X�a<F�a<�a<'�a<�a<��a<܇a<܇a<�a<̇a<߇a<��a<�a<�a<�a<#�a<"�a<Z�a<�  �  g�a<��a<��a<ψa<��a<+�a<Y�a<w�a<��a<݉a<*�a<o�a<��a<֊a<�a<h�a<��a<)�a<m�a<ǌa<"�a<�a<�a<D�a<��a<�a<~�a<ޏa<I�a<��a<)�a<��a<��a<��a<��a<o�a<��a<H�a<הa<N�a<ݕa<K�a<Ζa<E�a<Ɨa<E�a<Øa<N�a<��a<2�a<��a<�a<��a<�a<��a<��a<p�a<�a<k�a<�a<E�a<ɟa<3�a<��a<�a<r�a<ӡa<6�a<��a<��a<I�a<��a<�a<D�a<|�a<�a<+�a<x�a<¥a<�a<4�a<n�a<��a<ߦa<�a<P�a<w�a<��a<ϧa<�a< �a<?�a<g�a<|�a<��a<��a<ƨa<ܨa<��a<�a<D�a<S�a<P�a<}�a<z�a<��a<��a<��a<��a<��a<��a<��a<��a<ũa<��a<��a<��a<��a<��a<��a<~�a<e�a<X�a<S�a<8�a<!�a<�a<��a<Ԩa<��a<��a<~�a<H�a<3�a<��a<�a<§a<~�a<P�a<!�a<��a<Φa<��a<y�a<K�a<�a<�a<��a<y�a<C�a<�a<Τa<��a<B�a<��a<��a<q�a<�a<�a<��a<C�a<�a<��a<D�a<�a<��a<7�a<ߟa<x�a<�a<��a<R�a<��a<��a<�a<��a<!�a<ɛa<R�a<Қa<]�a<�a<y�a<�a<��a<!�a<��a<I�a<זa<s�a<�a<w�a<�a<��a<!�a<��a<F�a<a<U�a<Бa<��a<�a<��a<H�a<��a<l�a<�a<��a<D�a<�a<��a<0�a<ڌa<��a<B�a<ދa<��a<D�a<��a<��a<b�a<�a<ىa<��a<u�a<Y�a<%�a<�a<ֈa<��a<��a<s�a<P�a<6�a<%�a<�a<��a<�a<�a<Ӈa<ԇa<҇a<�a<�a<��a<��a<��a<�a<8�a<K�a<�  �  ��a<w�a<��a<Јa<��a</�a<P�a<��a<��a<�a<�a<\�a<��a<�a<B�a<u�a<Ӌa<�a<h�a<ߌa<�a<��a<ٍa<Q�a<��a<�a<~�a<ޏa<c�a<��a<2�a<��a<�a<n�a<�a<f�a<˓a<Y�a<ٔa<U�a<ȕa<G�a<�a<:�a<�a<>�a<͘a<<�a<��a</�a<��a<:�a<��a<&�a<��a<�a<��a<�a<z�a<͞a<`�a<˟a<'�a<��a<�a<��a<ϡa<S�a<��a<	�a<L�a<��a<��a<D�a<��a<ɤa<�a<`�a<��a<��a<0�a<{�a<��a<��a<�a<H�a<��a<��a<�a<�a<.�a<0�a<v�a<��a<��a<ɨa<Өa<�a<�a< �a<:�a<9�a<v�a<j�a<��a<��a<��a<��a<��a<ѩa<��a<کa<��a<��a<��a<��a<��a<��a<��a<p�a<u�a<u�a<\�a<V�a<&�a<=�a<��a<�a<ըa<��a<��a<u�a<V�a<�a<�a<ͧa<��a<��a<f�a<H�a<�a<�a<��a<u�a<c�a<	�a<�a<��a<��a<C�a<�a<Τa<��a<\�a<�a<ţa<k�a<.�a<̢a<}�a<:�a<աa<��a<F�a<�a<��a<3�a<��a<n�a<8�a<��a<\�a<�a<��a<�a<��a<D�a<��a<\�a<՚a<w�a<	�a<~�a<"�a<��a<<�a<×a<=�a<��a<Z�a<��a<s�a<"�a<��a<6�a<��a<+�a<̒a<V�a<�a<c�a<�a<��a<%�a<Տa<h�a<�a<��a<Y�a<�a<��a<C�a<ٌa<��a<&�a<�a<|�a<T�a<�a<��a<x�a<&�a<�a<��a<~�a<O�a<�a<
�a<Ĉa<��a<��a<s�a<X�a<4�a<8�a<��a<�a<߇a<�a<݇a<݇a<χa<��a<��a<·a<�a<�a<�a<;�a<9�a<�  �  d�a<��a<��a<҈a<�a<�a<M�a<��a<��a<��a<$�a<k�a<��a<�a<�a<|�a<Ëa<)�a<r�a<Ќa<&�a<��a<ԍa<O�a<��a<�a<��a<܏a<E�a<a<&�a<��a<�a<u�a<�a<W�a<ܓa<^�a<Ӕa<K�a<��a<F�a<Ȗa<C�a<՗a<H�a<ܘa<-�a<��a<<�a<��a</�a<��a< �a<��a<�a<��a<��a<n�a<�a<V�a<Ɵa<8�a<��a<��a<��a<ܡa<G�a<��a<�a<G�a<��a<�a<@�a<��a<פa<�a<h�a<��a<��a<"�a<o�a<��a<ܦa<�a<N�a<��a<��a<�a<�a<-�a<H�a<j�a<��a<��a<��a<ܨa<�a<�a<!�a<E�a<P�a<r�a<s�a<��a<��a<��a<ĩa<��a<��a<��a<��a<��a<ũa<��a<��a<��a<��a<��a<��a<y�a<k�a<D�a<P�a<9�a<�a<�a<��a<רa<Ψa<��a<s�a<_�a<+�a<�a<ާa<��a<��a<]�a<%�a<�a<զa<��a<~�a<S�a<�a<��a<��a<��a<V�a<�a<Фa<��a<>�a<	�a<��a<[�a<+�a<Ӣa<��a<+�a<�a<��a<@�a<�a<��a<2�a<ٟa<w�a<)�a<��a<k�a<םa<��a<�a<��a<:�a<ɛa<V�a<�a<m�a<��a<��a<�a<��a<2�a<��a<N�a<�a<M�a<�a<��a<�a<��a< �a<��a<H�a<��a<R�a<�a<r�a<��a<��a</�a<ҏa<Z�a<�a<��a<A�a<�a<��a<=�a<�a<��a<�a<�a<��a<G�a<��a<��a<g�a</�a<�a<��a<�a<Z�a<"�a<�a<̈a<��a<��a<]�a<h�a<;�a<'�a<�a<��a<�a<�a<Ǉa<҇a<ԇa<ևa<ɇa<�a<�a<�a< �a<5�a<L�a<�  �  Z�a<��a<��a<��a<�a<*�a<n�a<}�a<��a<�a<&�a<j�a<��a<�a<*�a<��a<��a<*�a<p�a<Ќa<*�a<��a<�a<H�a<��a<�a<�a<�a<8�a<��a<�a<��a<��a<g�a<�a<S�a<�a<9�a<֔a<@�a<Εa<A�a<Ɩa<[�a<˗a<.�a<��a<P�a<˙a<(�a<��a<#�a<��a<�a<��a<�a<��a<	�a<`�a<��a<J�a<џa<+�a<��a<�a<u�a<¡a<:�a<��a<�a<:�a<��a<ܣa<G�a<r�a<�a<�a<d�a<��a<ܥa<,�a<]�a<��a<ʦa<"�a<U�a<s�a<��a<اa<�a<!�a<C�a<m�a<��a<��a<��a<��a<�a<�a<�a<>�a<R�a<c�a<��a<}�a<��a<��a<��a<��a<��a<թa<��a<��a<��a<��a<��a<��a<��a<~�a<��a<]�a<g�a<N�a<B�a<7�a<�a<"�a<�a<Ǩa<��a<��a<��a<N�a<:�a<
�a<�a<��a<��a<|�a<0�a<+�a<ʦa<��a<}�a<S�a< �a<�a<Хa<~�a<0�a<��a<Ϥa<��a<1�a<�a<��a<e�a<�a<Ţa<��a<'�a<�a<w�a<C�a<ڠa<��a<-�a<ןa<��a<�a<��a<P�a<��a<��a<�a<��a<.�a<ћa<H�a<�a<v�a<��a<��a<�a<��a<&�a<ɗa<A�a<�a<t�a<�a<f�a<	�a<��a<�a<��a<9�a<��a<X�a<Ǒa<z�a<��a<��a<+�a<��a<d�a<��a<��a</�a<�a<��a<,�a<Ōa<��a<K�a<��a<��a<J�a<��a<��a<[�a<H�a<�a<ɉa<z�a<S�a<#�a<��a<܈a<��a<��a<u�a<C�a<&�a<�a<%�a<�a<�a<ۇa<ˇa<ԇa<��a<�a<Ƈa<�a<Շa<��a<	�a<'�a<J�a<�  �  i�a<{�a<��a<�a<��a</�a<Q�a<��a<ĉa<��a<�a<u�a<��a<��a<-�a<��a<ًa<(�a<p�a<�a<,�a<��a<�a<R�a<��a<(�a<d�a<ڏa<R�a<��a<'�a<��a<�a<j�a<ےa<N�a<ӓa<E�a<͔a<F�a<ȕa<I�a<Жa<,�a<ڗa<Q�a<Иa<C�a<ęa<:�a<ɚa<6�a<��a<-�a<��a<�a<��a<�a<�a<�a<^�a<ߟa<:�a<��a<�a<��a<ޡa<N�a<{�a<��a<E�a<��a<�a<;�a<��a<Фa<�a<Y�a<��a<�a<'�a<k�a<��a<�a<�a<4�a<��a<��a<�a<��a<$�a<G�a<��a<��a<��a<Ѩa<�a<�a<!�a</�a<O�a<H�a<q�a<��a<��a<��a<��a<��a<ȩa<��a<��a<��a<��a<��a<��a<��a<��a<��a<q�a<t�a<d�a<f�a<M�a<K�a<*�a<$�a<��a<�a<�a<��a<��a<v�a<X�a<=�a<�a<֧a<ȧa<��a<u�a<3�a<�a<�a<��a<}�a<e�a<"�a<�a<��a<��a<H�a<�a<��a<��a<K�a<�a<��a<d�a< �a<Ȣa<v�a<"�a<ݡa<��a<:�a<�a<��a<5�a<�a<`�a<.�a<Ğa<_�a<�a<��a<�a<��a<@�a<śa<c�a<�a<x�a<��a<��a<'�a<��a<:�a<חa<P�a<��a<d�a< �a<��a<�a<w�a<$�a<��a</�a<��a<M�a<ԑa<j�a<��a<��a<(�a<ŏa<_�a<�a<��a<G�a<�a<w�a<K�a<ߌa<��a<0�a<�a<��a<^�a<��a<��a<��a<:�a<��a<̉a<��a<d�a<�a<�a<�a<��a<��a<w�a<P�a<K�a<"�a<��a<��a<�a<݇a<̇a<҇a<��a<Ƈa<��a<҇a<܇a<��a<	�a<0�a<<�a<�  �  c�a<~�a<��a<Ԉa<��a<8�a<K�a<��a<��a<�a<3�a<|�a<��a<�a<C�a<r�a<Ջa<1�a<��a<ڌa<#�a<��a<Սa<b�a<��a<�a<y�a<܏a<D�a<��a<+�a<r�a<��a<d�a<�a<h�a<ɓa<W�a<��a<D�a<ҕa<1�a<Жa<:�a<ԗa<@�a<טa<=�a<͙a<M�a<��a<C�a<��a<1�a<��a<�a<��a<��a<��a<�a<j�a<ßa<C�a<��a<�a<��a<Ρa<F�a<��a<��a<1�a<��a<�a<�a<��a<¤a<#�a<b�a<��a<�a<�a<r�a<��a<צa<�a<F�a<��a<��a<�a<�a<B�a<E�a<n�a<��a<��a<̨a<Өa<�a<�a<)�a<T�a<Z�a<|�a<l�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ĩa<��a<��a<��a<��a<��a<{�a<o�a<R�a<?�a<T�a<�a<�a<�a<��a<ڨa<��a<��a<p�a<w�a<'�a<!�a<�a<ϧa<��a<\�a<J�a<�a<�a<¦a<��a<]�a<�a<�a<��a<��a<>�a<�a<ɤa<��a<=�a<�a<��a<L�a<�a<¢a<��a<<�a<ӡa<��a<�a<ޠa<��a<�a<�a<m�a<(�a<��a<f�a<�a<��a<*�a<��a<N�a<ћa<g�a<ޚa<v�a<�a<��a<(�a<��a<F�a<��a<Y�a<�a<_�a<
�a<s�a<�a<��a<#�a<��a<6�a<��a<1�a<�a<]�a<�a<��a<�a<Əa<H�a<�a<��a<;�a<�a<��a<<�a<Ԍa<��a<%�a<�a<��a<K�a<�a<Êa<{�a<'�a<�a<��a<��a<i�a<,�a<�a<ƈa<͈a<��a<y�a<W�a<8�a<(�a<��a<��a<чa<�a<��a<��a<̇a<Ça<݇a<هa<�a<�a<��a<9�a<.�a<�  �  U�a<��a<��a<Ԉa<��a<0�a<U�a<��a<��a<��a<0�a<h�a<��a<�a<H�a<��a<ԋa<+�a<y�a<�a<0�a<��a<��a<L�a<��a<�a<~�a<܏a<9�a<��a<�a<��a< �a<_�a<Вa<A�a<��a<A�a<Ԕa<;�a<Ǖa<@�a<Ėa<V�a<a<C�a<��a<H�a<��a<<�a<��a<7�a<��a<�a<��a<(�a<��a<�a<i�a<�a<^�a<ݟa<<�a<��a<�a<r�a<ӡa<5�a<��a<�a<@�a<��a<أa<=�a<|�a<��a<�a<I�a<��a<�a<(�a<M�a<��a<Ԧa<�a<T�a<y�a<��a<էa<��a<)�a<K�a<~�a<��a<��a<��a<�a<�a<*�a<>�a<=�a<^�a<t�a<}�a<��a<��a<��a<��a<��a<��a<ĩa<��a<��a<��a<��a<��a<��a<|�a<o�a<f�a<\�a<h�a<Q�a<1�a<0�a<�a<�a<�a<ڨa<��a<��a<z�a<\�a<8�a<�a<�a<��a<��a<��a<N�a<,�a<�a<��a<��a<f�a<&�a<�a<��a<��a<C�a<�a<Τa<��a<2�a<��a<��a<f�a<�a<��a<k�a<�a<ɡa<�a<A�a<ՠa<��a<,�a<՟a<��a<�a<��a<Q�a<�a<��a<�a<��a<B�a<՛a<P�a<�a<��a<�a<��a<�a<��a<:�a<՗a<R�a<ޖa<h�a<�a<x�a<�a<��a<�a<��a<2�a<��a<O�a<ёa<V�a<�a<}�a<�a<a<`�a<�a<��a<9�a<�a<��a<2�a<݌a<��a<0�a<�a<��a<[�a<�a<��a<m�a<T�a<�a<Չa<��a<S�a<0�a<�a<׈a<��a<��a<v�a<P�a<9�a<�a<�a<�a<�a<Їa<ʇa<Ӈa<��a<��a<��a<Ça<ԇa< �a<�a<�a<B�a<�  �  N�a<��a<��a<�a<��a<)�a<n�a<��a<҉a<�a<E�a<��a<��a<��a<�a<��a<Ћa<E�a<~�a<Ռa<9�a<��a<�a<?�a<��a<�a<g�a<ޏa<;�a<��a<�a<��a<ّa<s�a<�a<L�a<�a<-�a<͔a<5�a<��a<_�a<��a<D�a<��a<a�a<��a<U�a<șa<7�a<Κa<!�a<ԛa<#�a<��a<�a<|�a<�a<q�a<�a<N�a<�a<7�a<��a<%�a<i�a<�a<(�a<��a<ߢa<[�a<��a<ңa<<�a<`�a<�a<�a<^�a<��a<��a<,�a<J�a<��a<ߦa<�a<>�a<v�a<ça<ȧa<�a<$�a<P�a<z�a<��a<Шa<��a<�a<ۨa<!�a<5�a<P�a<z�a<^�a<��a<��a<��a<��a<��a<ʩa<��a<��a<��a<̩a<��a<��a<��a<��a<��a<u�a<��a<^�a<I�a<M�a<)�a<B�a<�a<
�a<٨a<�a<��a<��a<��a<R�a<K�a<�a<��a<էa<��a<y�a<�a<"�a<�a<צa<��a<Y�a</�a<�a<ӥa<t�a<U�a<	�a<��a<��a<4�a<�a<��a<l�a<��a<Ѣa<��a< �a<�a<j�a<;�a<Ϡa<��a<K�a<Ɵa<x�a<�a<Ԟa<I�a<��a<��a<�a<a<+�a<��a<Y�a<��a<t�a<��a<��a<�a<Ԙa<*�a<ڗa<M�a<�a<~�a<�a<��a<��a<��a<�a<��a<.�a<��a<M�a<��a<|�a<��a<��a<4�a<��a<e�a<�a<��a<D�a<�a<��a</�a<��a<{�a<O�a<�a<��a<W�a<��a<ߊa<n�a<F�a<؉a<̉a<��a<e�a<L�a<�a<�a<��a<��a<t�a<O�a<M�a<�a<	�a<߇a<��a<Ǉa<Ƈa<��a<��a<هa<��a<�a<ևa<�a<	�a<�a<U�a<�  �  S�a<��a<��a<ֈa<�a<%�a<f�a<��a<ωa<��a<4�a<t�a<��a<�a<S�a<��a<؋a<*�a<~�a<׌a<A�a<��a<�a<B�a<��a<�a<��a<�a<6�a<��a<�a<��a<�a<[�a<Œa<>�a<��a<G�a<��a<M�a<��a<>�a<��a<S�a<їa<K�a<��a<?�a<әa<K�a<ƚa<4�a<��a<&�a<��a<9�a<��a<�a<z�a<�a<]�a<ٟa<I�a<��a<�a<k�a<ڡa<C�a<��a<�a<;�a<|�a<�a<.�a<|�a<��a<��a<=�a<��a<եa<%�a<c�a<��a<Цa<�a<Y�a<~�a<��a<ϧa<�a<9�a<[�a<r�a<��a<��a<ͨa< �a<�a<9�a<8�a<F�a<`�a<o�a<��a<��a<��a<��a<��a<��a<ĩa<Ʃa<��a<��a<��a<��a<��a<��a<x�a<s�a<b�a<c�a<K�a<U�a<7�a<!�a<�a<�a<��a<ܨa<��a<��a<��a<m�a<H�a<�a<�a<ȧa<��a<��a<Y�a<4�a<�a<��a<��a<Z�a<7�a<�a<¥a<w�a<4�a<	�a<פa<��a</�a<�a<��a<f�a<�a<��a<`�a<�a<��a<��a<(�a<�a<t�a<*�a<Οa<��a<%�a<��a<G�a<�a<��a<(�a<��a<?�a<՛a<\�a<��a<��a<&�a<��a<"�a<��a<8�a<їa<_�a<�a<i�a<�a<�a<�a<��a<�a<��a<�a<��a<?�a<Бa<P�a<ߐa<p�a<�a<��a<]�a<��a<��a<4�a<�a<��a<7�a<Ԍa<��a<=�a<��a<��a<O�a<��a<��a<|�a<S�a<�a<�a<��a<[�a<1�a<�a<�a<Èa<��a<l�a<D�a<<�a<+�a<�a<�a<ۇa<̇a<Շa<��a<��a<��a<��a<��a<ۇa<�a<�a<�a<4�a<�  �  i�a<j�a<��a<̈a<�a<E�a<P�a<��a<��a<�a</�a<{�a<Ɋa<�a<#�a<��a<�a<(�a<��a<�a<3�a<��a<ٍa<r�a<��a<�a<n�a<��a<L�a<��a<�a<k�a<��a<\�a<��a<w�a<��a<c�a<��a<H�a<��a<H�a<Ɩa</�a<×a<>�a<�a<L�a<əa<=�a<��a<X�a<��a<@�a<��a<�a<y�a<
�a<��a<�a<��a<֟a<@�a<��a<�a<��a<ϡa<5�a<{�a<�a<K�a<��a<�a<	�a<��a<��a</�a<d�a<��a<�a<��a<_�a<��a<�a<��a<<�a<z�a<��a<��a<�a<*�a<Q�a<�a<��a<��a<�a<�a<�a<	�a<K�a<V�a<V�a<��a<u�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<m�a<��a<`�a<k�a<P�a<>�a<7�a<-�a<$�a<�a<�a<Ѩa<ƨa<��a<v�a<`�a<2�a<2�a<�a<ϧa<��a<]�a<*�a<�a<�a<��a<��a<l�a<)�a<�a<��a<��a<C�a<�a<��a<g�a<E�a<�a<��a<E�a<�a<��a<z�a<K�a<��a<��a<�a<�a<{�a<3�a<֟a<c�a<�a<��a<w�a<��a<��a<�a<��a<c�a<Ǜa<w�a<��a<i�a<�a<��a<<�a<��a<]�a<Ηa<V�a<�a<l�a<�a<t�a<�a<x�a<�a<��a< �a<��a<�a<�a<F�a<�a<��a<�a<Ώa<7�a<��a<��a<I�a<͍a<�a<3�a<ٌa<��a<(�a<�a<��a<\�a<�a<��a<��a<;�a<�a<��a<��a<k�a<(�a<#�a<ψa<��a<��a<��a<e�a</�a<�a<�a<��a<އa<̇a<ȇa<��a<χa<��a<�a<��a<�a<�a<��a<�a<@�a<�  �  S�a<��a<��a<ֈa<�a<%�a<f�a<��a<ωa<��a<4�a<t�a<��a<�a<S�a<��a<؋a<*�a<~�a<׌a<A�a<��a<�a<B�a<��a<�a<��a<�a<6�a<��a<�a<��a<�a<[�a<Œa<>�a<��a<G�a<��a<M�a<��a<>�a<��a<S�a<їa<K�a<��a<?�a<әa<K�a<ƚa<4�a<��a<&�a<��a<9�a<��a<�a<z�a<�a<]�a<ٟa<I�a<��a<�a<k�a<ڡa<C�a<��a<�a<;�a<|�a<�a<.�a<|�a<��a<��a<=�a<��a<եa<%�a<c�a<��a<Цa<�a<Y�a<~�a<��a<ϧa<�a<9�a<[�a<r�a<��a<��a<ͨa< �a<�a<9�a<8�a<F�a<`�a<o�a<��a<��a<��a<��a<��a<��a<ĩa<Ʃa<��a<��a<��a<��a<��a<��a<x�a<s�a<b�a<c�a<K�a<U�a<7�a<!�a<�a<�a<��a<ܨa<��a<��a<��a<m�a<H�a<�a<�a<ȧa<��a<��a<Y�a<4�a<�a<��a<��a<Z�a<7�a<�a<¥a<w�a<4�a<	�a<פa<��a</�a<�a<��a<f�a<�a<��a<`�a<�a<��a<��a<(�a<�a<t�a<*�a<Οa<��a<%�a<��a<G�a<�a<��a<(�a<��a<?�a<՛a<\�a<��a<��a<&�a<��a<"�a<��a<8�a<їa<_�a<�a<i�a<�a<�a<�a<��a<�a<��a<�a<��a<?�a<Бa<P�a<ߐa<p�a<�a<��a<]�a<��a<��a<4�a<�a<��a<7�a<Ԍa<��a<=�a<��a<��a<O�a<��a<��a<|�a<S�a<�a<�a<��a<[�a<1�a<�a<�a<Èa<��a<l�a<D�a<<�a<+�a<�a<�a<ۇa<̇a<Շa<��a<��a<��a<��a<��a<ۇa<�a<�a<�a<4�a<�  �  N�a<��a<��a<�a<��a<)�a<n�a<��a<҉a<�a<E�a<��a<��a<��a<�a<��a<Ћa<E�a<~�a<Ռa<9�a<��a<�a<?�a<��a<�a<g�a<ޏa<;�a<��a<�a<��a<ّa<s�a<�a<L�a<�a<-�a<͔a<5�a<��a<_�a<��a<D�a<��a<a�a<��a<U�a<șa<7�a<Κa<!�a<ԛa<#�a<��a<�a<|�a<�a<q�a<�a<N�a<�a<7�a<��a<%�a<i�a<�a<(�a<��a<ߢa<[�a<��a<ңa<<�a<`�a<�a<�a<^�a<��a<��a<,�a<J�a<��a<ߦa<�a<>�a<v�a<ça<ȧa<�a<$�a<P�a<z�a<��a<Шa<��a<�a<ۨa<!�a<5�a<P�a<z�a<^�a<��a<��a<��a<��a<��a<ʩa<��a<��a<��a<̩a<��a<��a<��a<��a<��a<u�a<��a<^�a<I�a<M�a<)�a<B�a<�a<
�a<٨a<�a<��a<��a<��a<R�a<K�a<�a<��a<էa<��a<y�a<�a<"�a<�a<צa<��a<Y�a</�a<�a<ӥa<t�a<U�a<	�a<��a<��a<4�a<�a<��a<l�a<��a<Ѣa<��a< �a<�a<j�a<;�a<Ϡa<��a<K�a<Ɵa<x�a<�a<Ԟa<I�a<��a<��a<�a<a<+�a<��a<Y�a<��a<t�a<��a<��a<�a<Ԙa<*�a<ڗa<M�a<�a<~�a<�a<��a<��a<��a<�a<��a<.�a<��a<M�a<��a<|�a<��a<��a<4�a<��a<e�a<�a<��a<D�a<�a<��a</�a<��a<{�a<O�a<�a<��a<W�a<��a<ߊa<n�a<F�a<؉a<̉a<��a<e�a<L�a<�a<�a<��a<��a<t�a<O�a<M�a<�a<	�a<߇a<��a<Ǉa<Ƈa<��a<��a<هa<��a<�a<ևa<�a<	�a<�a<U�a<�  �  U�a<��a<��a<Ԉa<��a<0�a<U�a<��a<��a<��a<0�a<h�a<��a<�a<H�a<��a<ԋa<+�a<y�a<�a<0�a<��a<��a<L�a<��a<�a<~�a<܏a<9�a<��a<�a<��a< �a<_�a<Вa<A�a<��a<A�a<Ԕa<;�a<Ǖa<@�a<Ėa<V�a<a<C�a<��a<H�a<��a<<�a<��a<7�a<��a<�a<��a<(�a<��a<�a<i�a<�a<^�a<ݟa<<�a<��a<�a<r�a<ӡa<5�a<��a<�a<@�a<��a<أa<=�a<|�a<��a<�a<I�a<��a<�a<(�a<M�a<��a<Ԧa<�a<T�a<y�a<��a<էa<��a<)�a<K�a<~�a<��a<��a<��a<�a<�a<*�a<>�a<=�a<^�a<t�a<}�a<��a<��a<��a<��a<��a<��a<ĩa<��a<��a<��a<��a<��a<��a<|�a<o�a<f�a<\�a<h�a<Q�a<1�a<0�a<�a<�a<�a<ڨa<��a<��a<z�a<\�a<8�a<�a<�a<��a<��a<��a<N�a<,�a<�a<��a<��a<f�a<&�a<�a<��a<��a<C�a<�a<Τa<��a<2�a<��a<��a<f�a<�a<��a<k�a<�a<ɡa<�a<A�a<ՠa<��a<,�a<՟a<��a<�a<��a<Q�a<�a<��a<�a<��a<B�a<՛a<P�a<�a<��a<�a<��a<�a<��a<:�a<՗a<R�a<ޖa<h�a<�a<x�a<�a<��a<�a<��a<2�a<��a<O�a<ёa<V�a<�a<}�a<�a<a<`�a<�a<��a<9�a<�a<��a<2�a<݌a<��a<0�a<�a<��a<[�a<�a<��a<m�a<T�a<�a<Չa<��a<S�a<0�a<�a<׈a<��a<��a<v�a<P�a<9�a<�a<�a<�a<�a<Їa<ʇa<Ӈa<��a<��a<��a<Ça<ԇa< �a<�a<�a<B�a<�  �  c�a<~�a<��a<Ԉa<��a<8�a<K�a<��a<��a<�a<3�a<|�a<��a<�a<C�a<r�a<Ջa<1�a<��a<ڌa<#�a<��a<Սa<b�a<��a<�a<y�a<܏a<D�a<��a<+�a<r�a<��a<d�a<�a<h�a<ɓa<W�a<��a<D�a<ҕa<1�a<Жa<:�a<ԗa<@�a<טa<=�a<͙a<M�a<��a<C�a<��a<1�a<��a<�a<��a<��a<��a<�a<j�a<ßa<C�a<��a<�a<��a<Ρa<F�a<��a<��a<1�a<��a<�a<�a<��a<¤a<#�a<b�a<��a<�a<�a<r�a<��a<צa<�a<F�a<��a<��a<�a<�a<B�a<E�a<n�a<��a<��a<̨a<Өa<�a<�a<)�a<T�a<Z�a<|�a<l�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ĩa<��a<��a<��a<��a<��a<{�a<o�a<R�a<?�a<T�a<�a<�a<�a<��a<ڨa<��a<��a<p�a<w�a<'�a<!�a<�a<ϧa<��a<\�a<J�a<�a<�a<¦a<��a<]�a<�a<�a<��a<��a<>�a<�a<ɤa<��a<=�a<�a<��a<L�a<�a<¢a<��a<<�a<ӡa<��a<�a<ޠa<��a<�a<�a<m�a<(�a<��a<f�a<�a<��a<*�a<��a<N�a<ћa<g�a<ޚa<v�a<�a<��a<(�a<��a<F�a<��a<Y�a<�a<_�a<
�a<s�a<�a<��a<#�a<��a<6�a<��a<1�a<�a<]�a<�a<��a<�a<Əa<H�a<�a<��a<;�a<�a<��a<<�a<Ԍa<��a<%�a<�a<��a<K�a<�a<Êa<{�a<'�a<�a<��a<��a<i�a<,�a<�a<ƈa<͈a<��a<y�a<W�a<8�a<(�a<��a<��a<чa<�a<��a<��a<̇a<Ça<݇a<هa<�a<�a<��a<9�a<.�a<�  �  i�a<{�a<��a<�a<��a</�a<Q�a<��a<ĉa<��a<�a<u�a<��a<��a<-�a<��a<ًa<(�a<p�a<�a<,�a<��a<�a<R�a<��a<(�a<d�a<ڏa<R�a<��a<'�a<��a<�a<j�a<ےa<N�a<ӓa<E�a<͔a<F�a<ȕa<I�a<Жa<,�a<ڗa<Q�a<Иa<C�a<ęa<:�a<ɚa<6�a<��a<-�a<��a<�a<��a<�a<�a<�a<^�a<ߟa<:�a<��a<�a<��a<ޡa<N�a<{�a<��a<E�a<��a<�a<;�a<��a<Фa<�a<Y�a<��a<�a<'�a<k�a<��a<�a<�a<4�a<��a<��a<�a<��a<$�a<G�a<��a<��a<��a<Ѩa<�a<�a<!�a</�a<O�a<H�a<q�a<��a<��a<��a<��a<��a<ȩa<��a<��a<��a<��a<��a<��a<��a<��a<��a<q�a<t�a<d�a<f�a<M�a<K�a<*�a<$�a<��a<�a<�a<��a<��a<v�a<X�a<=�a<�a<֧a<ȧa<��a<u�a<3�a<�a<�a<��a<}�a<e�a<"�a<�a<��a<��a<H�a<�a<��a<��a<K�a<�a<��a<d�a< �a<Ȣa<v�a<"�a<ݡa<��a<:�a<�a<��a<5�a<�a<`�a<.�a<Ğa<_�a<�a<��a<�a<��a<@�a<śa<c�a<�a<x�a<��a<��a<'�a<��a<:�a<חa<P�a<��a<d�a< �a<��a<�a<w�a<$�a<��a</�a<��a<M�a<ԑa<j�a<��a<��a<(�a<ŏa<_�a<�a<��a<G�a<�a<w�a<K�a<ߌa<��a<0�a<�a<��a<^�a<��a<��a<��a<:�a<��a<̉a<��a<d�a<�a<�a<�a<��a<��a<w�a<P�a<K�a<"�a<��a<��a<�a<݇a<̇a<҇a<��a<Ƈa<��a<҇a<܇a<��a<	�a<0�a<<�a<�  �  Z�a<��a<��a<��a<�a<*�a<n�a<}�a<��a<�a<&�a<j�a<��a<�a<*�a<��a<��a<*�a<p�a<Ќa<*�a<��a<�a<H�a<��a<�a<�a<�a<8�a<��a<�a<��a<��a<g�a<�a<S�a<�a<9�a<֔a<@�a<Εa<A�a<Ɩa<[�a<˗a<.�a<��a<P�a<˙a<(�a<��a<#�a<��a<�a<��a<�a<��a<	�a<`�a<��a<J�a<џa<+�a<��a<�a<u�a<¡a<:�a<��a<�a<:�a<��a<ܣa<G�a<r�a<�a<�a<d�a<��a<ܥa<,�a<]�a<��a<ʦa<"�a<U�a<s�a<��a<اa<�a<!�a<C�a<m�a<��a<��a<��a<��a<�a<�a<�a<>�a<R�a<c�a<��a<}�a<��a<��a<��a<��a<��a<թa<��a<��a<��a<��a<��a<��a<��a<~�a<��a<]�a<g�a<N�a<B�a<7�a<�a<"�a<�a<Ǩa<��a<��a<��a<N�a<:�a<
�a<�a<��a<��a<|�a<0�a<+�a<ʦa<��a<}�a<S�a< �a<�a<Хa<~�a<0�a<��a<Ϥa<��a<1�a<�a<��a<e�a<�a<Ţa<��a<'�a<�a<w�a<C�a<ڠa<��a<-�a<ןa<��a<�a<��a<P�a<��a<��a<�a<��a<.�a<ћa<H�a<�a<v�a<��a<��a<�a<��a<&�a<ɗa<A�a<�a<t�a<�a<f�a<	�a<��a<�a<��a<9�a<��a<X�a<Ǒa<z�a<��a<��a<+�a<��a<d�a<��a<��a</�a<�a<��a<,�a<Ōa<��a<K�a<��a<��a<J�a<��a<��a<[�a<H�a<�a<ɉa<z�a<S�a<#�a<��a<܈a<��a<��a<u�a<C�a<&�a<�a<%�a<�a<�a<ۇa<ˇa<ԇa<��a<�a<Ƈa<�a<Շa<��a<	�a<'�a<J�a<�  �  d�a<��a<��a<҈a<�a<�a<M�a<��a<��a<��a<$�a<k�a<��a<�a<�a<|�a<Ëa<)�a<r�a<Ќa<&�a<��a<ԍa<O�a<��a<�a<��a<܏a<E�a<a<&�a<��a<�a<u�a<�a<W�a<ܓa<^�a<Ӕa<K�a<��a<F�a<Ȗa<C�a<՗a<H�a<ܘa<-�a<��a<<�a<��a</�a<��a< �a<��a<�a<��a<��a<n�a<�a<V�a<Ɵa<8�a<��a<��a<��a<ܡa<G�a<��a<�a<G�a<��a<�a<@�a<��a<פa<�a<h�a<��a<��a<"�a<o�a<��a<ܦa<�a<N�a<��a<��a<�a<�a<-�a<H�a<j�a<��a<��a<��a<ܨa<�a<�a<!�a<E�a<P�a<r�a<s�a<��a<��a<��a<ĩa<��a<��a<��a<��a<��a<ũa<��a<��a<��a<��a<��a<��a<y�a<k�a<D�a<P�a<9�a<�a<�a<��a<רa<Ψa<��a<s�a<_�a<+�a<�a<ާa<��a<��a<]�a<%�a<�a<զa<��a<~�a<S�a<�a<��a<��a<��a<V�a<�a<Фa<��a<>�a<	�a<��a<[�a<+�a<Ӣa<��a<+�a<�a<��a<@�a<�a<��a<2�a<ٟa<w�a<)�a<��a<k�a<םa<��a<�a<��a<:�a<ɛa<V�a<�a<m�a<��a<��a<�a<��a<2�a<��a<N�a<�a<M�a<�a<��a<�a<��a< �a<��a<H�a<��a<R�a<�a<r�a<��a<��a</�a<ҏa<Z�a<�a<��a<A�a<�a<��a<=�a<�a<��a<�a<�a<��a<G�a<��a<��a<g�a</�a<�a<��a<�a<Z�a<"�a<�a<̈a<��a<��a<]�a<h�a<;�a<'�a<�a<��a<�a<�a<Ǉa<҇a<ԇa<ևa<ɇa<�a<�a<�a< �a<5�a<L�a<�  �  ��a<w�a<��a<Јa<��a</�a<P�a<��a<��a<�a<�a<\�a<��a<�a<B�a<u�a<Ӌa<�a<h�a<ߌa<�a<��a<ٍa<Q�a<��a<�a<~�a<ޏa<c�a<��a<2�a<��a<�a<n�a<�a<f�a<˓a<Y�a<ٔa<U�a<ȕa<G�a<�a<:�a<�a<>�a<͘a<<�a<��a</�a<��a<:�a<��a<&�a<��a<�a<��a<�a<z�a<͞a<`�a<˟a<'�a<��a<�a<��a<ϡa<S�a<��a<	�a<L�a<��a<��a<D�a<��a<ɤa<�a<`�a<��a<��a<0�a<{�a<��a<��a<�a<H�a<��a<��a<�a<�a<.�a<0�a<v�a<��a<��a<ɨa<Өa<�a<�a< �a<:�a<9�a<v�a<j�a<��a<��a<��a<��a<��a<ѩa<��a<کa<��a<��a<��a<��a<��a<��a<��a<p�a<u�a<u�a<\�a<V�a<&�a<=�a<��a<�a<ըa<��a<��a<u�a<V�a<�a<�a<ͧa<��a<��a<f�a<H�a<�a<�a<��a<u�a<c�a<	�a<�a<��a<��a<C�a<�a<Τa<��a<\�a<�a<ţa<k�a<.�a<̢a<}�a<:�a<աa<��a<F�a<�a<��a<3�a<��a<n�a<8�a<��a<\�a<�a<��a<�a<��a<D�a<��a<\�a<՚a<w�a<	�a<~�a<"�a<��a<<�a<×a<=�a<��a<Z�a<��a<s�a<"�a<��a<6�a<��a<+�a<̒a<V�a<�a<c�a<�a<��a<%�a<Տa<h�a<�a<��a<Y�a<�a<��a<C�a<ٌa<��a<&�a<�a<|�a<T�a<�a<��a<x�a<&�a<�a<��a<~�a<O�a<�a<
�a<Ĉa<��a<��a<s�a<X�a<4�a<8�a<��a<�a<߇a<�a<݇a<݇a<χa<��a<��a<·a<�a<�a<�a<;�a<9�a<�  �  g�a<��a<��a<ψa<��a<+�a<Y�a<w�a<��a<݉a<*�a<o�a<��a<֊a<�a<h�a<��a<)�a<m�a<ǌa<"�a<�a<�a<D�a<��a<�a<~�a<ޏa<I�a<��a<)�a<��a<��a<��a<��a<o�a<��a<H�a<הa<N�a<ݕa<K�a<Ζa<E�a<Ɨa<E�a<Øa<N�a<��a<2�a<��a<�a<��a<�a<��a<��a<p�a<�a<k�a<�a<E�a<ɟa<3�a<��a<�a<r�a<ӡa<6�a<��a<��a<I�a<��a<�a<D�a<|�a<�a<+�a<x�a<¥a<�a<4�a<n�a<��a<ߦa<�a<P�a<w�a<��a<ϧa<�a< �a<?�a<g�a<|�a<��a<��a<ƨa<ܨa<��a<�a<D�a<S�a<P�a<}�a<z�a<��a<��a<��a<��a<��a<��a<��a<��a<ũa<��a<��a<��a<��a<��a<��a<~�a<e�a<X�a<S�a<8�a<!�a<�a<��a<Ԩa<��a<��a<~�a<H�a<3�a<��a<�a<§a<~�a<P�a<!�a<��a<Φa<��a<y�a<K�a<�a<�a<��a<y�a<C�a<�a<Τa<��a<B�a<��a<��a<q�a<�a<�a<��a<C�a<�a<��a<D�a<�a<��a<7�a<ߟa<x�a<�a<��a<R�a<��a<��a<�a<��a<!�a<ɛa<R�a<Қa<]�a<�a<y�a<�a<��a<!�a<��a<I�a<זa<s�a<�a<w�a<�a<��a<!�a<��a<F�a<a<U�a<Бa<��a<�a<��a<H�a<��a<l�a<�a<��a<D�a<�a<��a<0�a<ڌa<��a<B�a<ދa<��a<D�a<��a<��a<b�a<�a<ىa<��a<u�a<Y�a<%�a<�a<ֈa<��a<��a<s�a<P�a<6�a<%�a<�a<��a<�a<�a<Ӈa<ԇa<҇a<�a<�a<��a<��a<��a<�a<8�a<K�a<�  �  ^�a<��a<��a<وa<�a<�a<W�a<r�a<ɉa<։a<)�a<K�a<��a<�a<!�a<��a<��a<�a<i�a<��a<?�a<q�a<�a<0�a<Îa<�a<�a<��a<C�a<̐a<�a<��a<
�a<~�a<�a<B�a<�a<K�a<��a<I�a<ܕa<M�a<ɖa<`�a<��a<a�a<��a<:�a<��a<B�a<��a<�a<��a<��a<��a<�a<��a<�a<K�a<�a<@�a<ɟa<K�a<��a<	�a<f�a<�a<,�a<��a<��a<F�a<��a<�a<f�a<��a<�a<	�a<e�a<��a<�a<T�a<Y�a<��a<٦a< �a<X�a<r�a<ŧa<��a<��a<�a<^�a<]�a<v�a<��a<��a<�a<�a<�a<'�a<�a<X�a<K�a<��a<{�a<��a<��a<��a<éa<��a<שa<��a<ʩa<��a<��a<ȩa<��a<��a<h�a<��a<w�a<~�a<h�a<=�a<H�a<�a<!�a<�a<ިa<Ȩa<��a<}�a<C�a<B�a<�a<�a<��a<��a<n�a<'�a<�a<Ŧa<��a<u�a<A�a<5�a<եa<��a<e�a<[�a<�a<Ϥa<��a<<�a<�a<��a<��a<(�a<ܢa<��a<�a<�a<��a<e�a<�a<��a<9�a<ڟa<��a<�a<Ӟa<K�a<�a<~�a<�a<��a<�a<̛a<.�a<�a<p�a<��a<��a<�a<��a<�a<a<a�a<Ζa<b�a<�a<��a<��a<��a<!�a<��a<I�a<��a<x�a<בa<��a<�a<��a<>�a<ʏa<��a<�a<��a<>�a<�a<��a<+�a<��a<q�a<1�a<΋a<��a<;�a<�a<��a<Q�a<D�a<�a<a<��a<3�a<*�a<߈a<߈a<��a<��a<[�a<X�a<F�a<�a<'�a<�a<��a<܇a<܇a<�a<̇a<߇a<��a<�a<�a<�a<#�a<"�a<Z�a<�  �  y�a<��a<��a<Ĉa< �a<4�a<_�a<u�a<��a<�a<+�a<Q�a<��a<ӊa<�a<d�a<ŋa<�a<{�a<��a<�a<z�a<�a<S�a<��a<�a<r�a<�a<Z�a<Đa<&�a<��a<�a<�a<�a<}�a<��a<Y�a<֔a<I�a<ѕa<Z�a<ܖa<M�a<��a<A�a<ɘa<P�a<��a<-�a<��a<-�a<��a<�a<��a<�a<h�a<�a<h�a<ޞa<Z�a<��a<-�a<��a<�a<~�a<١a<0�a<��a<�a<V�a<��a<�a<D�a<��a<�a<>�a<��a<��a<�a<3�a<m�a<��a<�a<)�a<D�a<m�a<��a<ߧa<�a<�a<>�a<S�a<��a<��a<��a<��a<ިa<��a<�a<(�a<T�a<`�a<e�a<x�a<��a<��a<��a<��a<��a<ȩa<ѩa<Ωa<��a<��a<��a<��a<��a<��a<��a<z�a<o�a<\�a<K�a<G�a<4�a<�a<�a<ɨa<��a<��a<��a<G�a<#�a<�a<�a<��a<��a<L�a<%�a<�a<צa<��a<��a<A�a<�a<ߥa<��a<��a<H�a<��a<¤a<��a<S�a<�a<��a<s�a< �a<ݢa<��a<Q�a<��a<��a<D�a<�a<��a<F�a<�a<��a<�a<��a<Y�a<��a<��a<	�a<��a<7�a<ěa<I�a<Κa<P�a<�a<t�a<�a<��a<6�a<��a<C�a<Ֆa<t�a<��a<~�a<��a<��a<1�a<��a<>�a<��a<V�a<�a<��a<#�a<��a<<�a<ȏa<l�a<�a<��a<S�a<��a<��a<&�a<�a<��a<>�a<؋a<��a<0�a< �a<��a<i�a<�a<ۉa<��a<s�a<=�a<&�a<�a<��a<��a<��a<~�a<V�a<(�a<�a<�a<�a<��a<�a<ڇa<Շa<҇a<��a<��a<��a<�a<�a<�a<0�a<Y�a<�  �  ��a<x�a<ȉa<׉a<�a<�a<;�a<��a<��a<�a<�a<^�a<��a<ʋa<@�a<V�a<ٌa<��a<W�a<��a<"�a<��a<Îa<1�a<��a<�a<~�a<Аa<c�a<�a<3�a<��a<��a<a�a<Ǔa<P�a<��a<U�a<��a<_�a<��a<(�a<Зa<�a<Ęa<�a<��a<��a<��a<�a<��a<��a<I�a<�a<R�a<ٝa<X�a<��a<C�a<~�a<�a<��a<��a<Z�a<��a<*�a<�a<�a<P�a<ˣa<�a<?�a<դa<�a<c�a<~�a<֥a<�a<]�a<��a<�a<L�a<A�a<��a<ݧa<�a<Q�a<C�a<��a<��a<ިa<�a<�a<3�a<;�a<��a<t�a<ȩa<��a<�a<��a<�a<#�a<3�a<U�a<C�a<N�a<]�a<x�a<��a<i�a<��a<c�a<z�a<��a<d�a<y�a<D�a<h�a<7�a<D�a<(�a<0�a<�a<ԩa<�a<��a<ϩa<��a<i�a<I�a<#�a<)�a<�a<Ǩa<��a<v�a<[�a<
�a<�a<��a<��a<R�a<,�a<�a<�a<��a<]�a<3�a<�a<ܥa<��a<F�a<,�a<��a<��a<2�a<�a<��a<:�a<��a<��a<o�a<�a<١a<@�a<��a<Ơa<4�a<�a<q�a<
�a<��a<;�a<ߝa<l�a<�a<h�a<'�a<��a<A�a<ٚa<D�a<��a<P�a<�a<��a<'�a<��a<&�a<Ɩa<E�a<�a<q�a<�a<��a<�a<ԓa<*�a<�a<I�a<�a<{�a<�a<ΐa<T�a<�a<u�a<X�a<�a<��a<E�a<��a<z�a<�a<ٌa<��a<5�a<�a<��a<��a<�a<�a<��a<��a<R�a<��a<��a<Ήa<��a<y�a<Y�a<B�a<<�a<B�a<��a<+�a<Ԉa<�a<��a<ˈa<�a<��a<�a<Ոa<��a< �a<,�a<>�a<'�a<�  �  a�a<p�a<��a<Ɖa<	�a<.�a<\�a<}�a<��a<�a<-�a<Z�a<��a<ыa<�a<j�a<Ȍa<�a<x�a<��a<�a<x�a<�a<E�a<��a<��a<_�a<��a<7�a<��a<�a<w�a<��a<a�a<�a<f�a<��a<C�a<��a<2�a<��a<'�a<��a<�a<��a<�a<��a<#�a<��a<�a<|�a<��a<o�a<�a<Z�a<��a<4�a<��a<1�a<��a<�a<��a<�a<h�a<ۡa<<�a<��a<�a<>�a<��a<��a<W�a<��a<�a<Q�a<��a<�a<3�a<d�a<��a<ߦa<(�a<c�a<��a<��a<��a<+�a<f�a<��a<Ǩa<ܨa<��a<�a<P�a<V�a<��a<��a<��a<��a<�a<�a<�a<!�a<+�a<A�a<_�a<j�a<y�a<l�a<t�a<f�a<u�a<z�a<z�a<u�a<j�a<j�a<[�a<q�a<K�a<9�a<,�a<�a<�a<��a<ܩa<��a<��a<��a<��a<e�a<D�a<�a<�a<ɨa<��a<s�a<Q�a<�a<�a<��a<��a<f�a<M�a<
�a<զa<��a<��a<F�a<�a<��a<~�a<*�a<�a<��a<z�a<%�a<�a<��a<U�a<�a<��a<]�a<��a<��a<Q�a<��a<��a<-�a<ןa<{�a<$�a<��a<O�a<ԝa<h�a<�a<��a<�a<��a<$�a<��a<S�a<�a<s�a<�a<��a<�a<��a<P�a<ؖa<Y�a<ەa<_�a<�a<��a<�a<��a</�a<Ԓa<[�a<	�a<��a<�a<��a<N�a<��a<��a<4�a<��a<t�a<�a<ԍa<��a<:�a<׌a<��a<8�a<�a<��a<m�a< �a<��a<��a<��a<H�a<&�a<�a<ŉa<��a<��a<u�a<^�a<0�a<�a<��a<�a<�a<�a<ڈa<шa<؈a<Ԉa<��a<�a<�a<�a<�a<3�a<G�a<�  �  N�a<��a<��a<ʉa<�a< �a<R�a<p�a<a<֊a<-�a<Q�a<��a<�a<�a<��a<��a<�a<j�a<��a<"�a<d�a<ێa<�a<��a<��a<��a<�a<(�a<ȑa<�a<��a<��a<`�a<ѓa<:�a<Ҕa<7�a<Еa<$�a<Ŗa<3�a<��a<Q�a<��a<*�a<��a<��a<z�a<��a<��a<�a<|�a<Μa<o�a<՝a<D�a<Ӟa<�a<��a<�a<��a<�a<L�a<��a<�a<��a<�a<z�a<��a<�a<v�a<��a<�a<C�a<��a<ʥa<�a<f�a<��a<��a<�a<��a<��a<ܧa<#�a<&�a<z�a<k�a<��a<Ǩa<��a<�a<:�a<_�a<a�a<��a<��a<թa<�a<�a<�a<
�a<B�a<6�a<P�a<>�a<n�a<q�a<x�a<��a<e�a<��a<�a<o�a<��a<c�a<g�a<=�a<L�a<5�a<:�a<�a<�a<�a<ɩa<�a<��a<��a<��a<7�a<:�a<�a<��a<��a<��a<i�a<L�a<4�a<�a<�a<��a<n�a<@�a<�a<�a<��a<u�a<�a<�a<��a<��a<X�a<�a<�a<f�a<8�a<�a<��a<D�a<�a<��a<P�a<�a<��a<k�a<�a<��a<m�a<ԟa<��a<�a<��a<2�a<ʝa<s�a<�a<��a<�a<��a<=�a<Śa<m�a<͙a<}�a<��a<��a<�a<��a<1�a<��a<l�a<ٕa<��a<��a<��a<8�a<��a<T�a<ǒa<h�a<�a<{�a< �a<��a<g�a<�a<��a<+�a<�a<��a<�a<�a<Y�a<*�a<a<��a<2�a<�a<��a<N�a<A�a<�a<��a<��a<9�a<.�a<މa<݉a<��a<��a<I�a<S�a<5�a< �a<3�a<�a<�a<�a<Ԉa<�a<Јa<߈a<ǈa<�a<�a<�a<�a<-�a<d�a<�  �  f�a<��a<��a<Љa<��a<%�a<k�a<}�a<Êa<�a<#�a<g�a<��a<ۋa<%�a<m�a<��a<!�a<a�a<��a<$�a<w�a<��a<<�a<��a<��a<b�a<ʐa<:�a<��a<�a<��a<�a<k�a<�a<D�a<ߔa<.�a<��a<0�a<��a<#�a<��a<�a<��a<%�a<��a<#�a<��a<�a<��a<��a<x�a<�a<Q�a<˝a<?�a<��a<1�a<��a<�a<��a<�a<f�a<ܡa<1�a<��a<�a<K�a<��a<��a<Y�a<��a<�a<8�a<��a<٥a<&�a<r�a<��a<�a<"�a<e�a<��a<ϧa<��a<+�a<l�a<��a<Шa<بa<�a<#�a<7�a<k�a<t�a<��a<��a<©a<ԩa<��a<�a<�a<F�a<@�a<k�a<i�a<p�a<t�a<p�a<v�a<{�a<y�a<z�a<}�a<e�a<_�a<t�a<K�a<[�a<6�a<�a<&�a<�a<��a<�a<éa<��a<��a<|�a<\�a<S�a<�a< �a<èa<��a<�a<D�a<�a<�a<§a<��a<{�a<6�a<�a<�a<��a<��a<>�a<�a<¥a<��a<@�a<�a<��a<r�a<9�a<գa<��a<U�a<�a<Ģa<H�a<�a<��a<R�a<�a<��a<:�a<՟a<��a<�a<��a<O�a<ӝa<x�a<��a<��a< �a<��a<3�a<��a<N�a<�a<�a<�a<��a<�a<��a<Q�a<͖a<b�a<ܕa<m�a<��a<��a<�a<��a<B�a<��a<t�a<�a<��a<-�a<��a<b�a<�a<��a<6�a<َa<{�a<�a<ۍa<}�a<C�a<ӌa<��a<>�a<�a<��a<a�a< �a<�a<��a<q�a<R�a<#�a<�a<�a<��a<��a<t�a<U�a<8�a<�a<�a<��a<�a<�a<�a<̈a<̈a<�a<Ԉa<��a<�a<��a<"�a<,�a<H�a<�  �  ��a<z�a<��a<̉a<�a<'�a<F�a<�a<��a<��a<�a<\�a<��a<�a<?�a<r�a<ˌa<�a<h�a<͍a<�a<z�a<͎a<<�a<��a<�a<k�a<Đa<O�a<��a<�a<z�a<�a<_�a<ғa<A�a<��a<<�a<��a<1�a<��a<(�a<��a<�a<��a<�a<��a<�a<��a<�a<w�a<�a<\�a<�a<S�a<ޝa<X�a<��a<;�a<��a<�a<��a<�a<]�a<��a<0�a<��a<�a<C�a<��a<�a<N�a<��a<��a<K�a<��a<ҥa<�a<a�a<��a<�a<&�a<T�a<��a<̧a< �a<H�a<Q�a<��a<��a<٨a<��a<(�a<B�a<S�a<��a<��a<ũa<̩a<ݩa<��a<��a<2�a<(�a<@�a<K�a<b�a<`�a<g�a<��a<m�a<��a<s�a<s�a<q�a<g�a<f�a<V�a<L�a<?�a<:�a<(�a<�a<�a<�a<��a<��a<ȩa<��a<o�a<^�a<.�a<�a<�a<بa<��a<u�a<O�a<#�a<�a<ȧa<��a<d�a<=�a<�a<Ҧa<��a<g�a<>�a<�a<ӥa<��a<:�a<�a<��a<x�a<(�a<�a<��a<E�a<�a<��a<V�a<��a<��a<L�a<��a<��a<.�a<��a<k�a<�a<��a<B�a<ӝa<c�a<
�a<z�a<&�a<��a<F�a<ٚa<O�a<�a<a�a<�a<��a<�a<��a<3�a<̖a<F�a<��a<d�a<
�a<��a<�a<��a<6�a<Βa<V�a<�a<��a<�a<��a<Q�a<��a<��a<H�a<׎a<}�a<;�a<��a<}�a<�a<Ԍa<}�a<C�a<�a<��a<r�a<%�a<�a<��a<z�a<N�a<�a<�a<a<��a<��a<m�a<E�a<+�a<;�a<��a<�a<�a<܈a<׈a<Έa<ӈa<ψa<ֈa<ވa<�a< �a<�a<,�a<@�a<�  �  W�a<��a<��a<��a<�a< �a<E�a<��a<��a<ߊa<&�a<h�a<��a<�a<�a<~�a<Ȍa<�a<l�a<��a<$�a<��a<͎a<<�a<��a<�a<e�a<Ӑa<)�a<��a<�a<x�a<�a<Q�a<ٓa<P�a<��a<0�a<��a<"�a<��a<!�a<��a<�a<��a<�a<��a<�a<��a<#�a<z�a<�a<y�a<�a<_�a<ѝa<C�a<��a<4�a<��a<�a<��a<	�a<n�a<��a<C�a<��a<�a<J�a<��a<��a<b�a<��a<�a<>�a<��a<�a<&�a<Z�a<��a<�a<�a<d�a<��a<Чa<��a<#�a<_�a<��a<��a<��a<
�a<�a<A�a<j�a<�a<��a<��a<ѩa<�a<��a<�a<�a</�a<g�a<J�a<Y�a<~�a<[�a<t�a<|�a<r�a<x�a<��a<f�a<r�a<Z�a<[�a<U�a<E�a<*�a<0�a<�a<�a<�a<ҩa<ͩa<��a<��a<��a<W�a<-�a<:�a<�a<��a<��a<��a<X�a<,�a<�a<ӧa<��a<t�a<B�a<�a<�a<Ŧa<g�a<>�a<�a<��a<��a<I�a<�a<��a<x�a<&�a<�a<��a<K�a<��a<��a<J�a<��a<��a<_�a<�a<��a<9�a<ӟa<m�a<)�a<��a<K�a<��a<f�a<��a<��a< �a<��a<9�a<Ěa<X�a<�a<��a<��a<��a<7�a<��a<3�a<ߖa<L�a<וa<k�a<��a<�a<$�a<��a<2�a<��a<Y�a<��a<��a<�a<��a<N�a<�a<��a<(�a<ڎa<z�a<�a<͍a<��a<�a<�a<��a<4�a<�a<��a<l�a<-�a<��a<��a<��a<S�a<$�a<�a<ɉa<͉a<��a<d�a<c�a<�a<�a<�a<��a<�a<�a<ˈa<؈a<ǈa<Ԉa<ވa<�a<�a<�a<
�a<6�a<F�a<�  �  [�a<��a<��a<߉a<�a<�a<[�a<|�a<��a<�a<:�a<q�a<��a<��a<(�a<��a<��a<.�a<s�a<ōa<�a<x�a<�a<4�a<��a<
�a<e�a<אa<0�a<��a<�a<��a<�a<R�a<ٓa<?�a<Ŕa<"�a<ȕa<$�a<��a<�a<��a<&�a<��a<-�a<��a<�a<��a<�a<��a<�a<��a<�a<b�a<ޝa<Q�a<ʞa<(�a<şa<�a<��a<�a<i�a<̡a<.�a<��a<�a<Q�a<��a<��a<Y�a<��a<�a<-�a<��a<ҥa< �a<Z�a<��a<��a<�a<`�a<��a<֧a<��a<8�a<t�a<��a<��a<ݨa<��a<%�a<A�a<|�a<n�a<��a<��a<ݩa<ܩa<�a<(�a< �a<7�a<B�a<`�a<`�a<v�a<��a<n�a<��a<r�a<t�a<p�a<u�a<y�a<H�a<b�a<@�a<M�a<�a<2�a<#�a<��a<�a<֩a<Щa<��a<��a<��a<V�a<C�a<�a<�a<ɨa<��a<��a<C�a<8�a<��a<ާa<��a<��a<H�a<�a<ަa<��a<��a<5�a<�a<Υa<��a<M�a<��a<��a<j�a<>�a<ڣa<��a<L�a<�a<��a<;�a<�a<��a<N�a<�a<��a<A�a<ڟa<��a<�a<��a<O�a<؝a<w�a<��a<��a<�a<��a<E�a<Қa<e�a<ݙa<��a<�a<��a<�a<��a<A�a<ʖa<g�a<�a<s�a<�a<��a<�a<��a<M�a<��a<\�a<�a<��a<�a<��a<g�a<�a<��a<-�a<�a<|�a<+�a<�a<x�a<1�a<ٌa<��a<@�a<�a<ɋa<[�a<:�a<�a<Ȋa<z�a<W�a<:�a<�a<щa<��a<��a<k�a<[�a<F�a<�a<�a<�a<�a<؈a<ڈa<��a<��a<ۈa<Ɉa<�a<ֈa<
�a<�a<$�a<B�a<�  �  ��a<v�a<��a<މa<�a<(�a<Y�a<w�a<��a<��a<"�a<p�a<��a<�a<<�a<��a<ǌa<&�a<f�a<ԍa<!�a<z�a<ݎa<7�a<��a<�a<\�a<Ða<S�a<��a<��a<y�a<�a<]�a<̓a<3�a<��a<0�a<��a<%�a<��a<.�a<��a<�a<��a<�a<��a<�a<��a<��a<��a<��a<s�a<�a<c�a<�a<]�a<Ǟa<8�a<��a<�a<��a<�a<c�a<ša<"�a<��a<�a<B�a<��a<�a<I�a<��a<��a<<�a<��a<ĥa<�a<\�a<��a<�a<�a<Q�a<��a<˧a<��a<F�a<S�a<��a<��a<�a< �a<5�a<=�a<k�a<~�a<��a<éa<ةa<ީa<�a<�a<1�a<<�a<<�a<]�a<d�a<U�a<|�a<v�a<k�a<��a<y�a<f�a<k�a<f�a<]�a<W�a<2�a<B�a<5�a<%�a<�a<��a<�a<��a<��a<��a<��a<c�a<_�a<A�a<�a<��a<ۨa<��a<��a<L�a<0�a<	�a<קa<��a<��a<<�a<!�a<�a<��a<w�a<8�a<�a<֥a<{�a<:�a<�a<��a<d�a<'�a<ۣa<��a<?�a<�a<��a<J�a<�a<��a<B�a<��a<��a<1�a<�a<s�a<�a<��a<I�a<ѝa<z�a<��a<��a<*�a<��a<P�a<ޚa<b�a<�a<z�a<�a<��a<�a<��a<:�a<��a<M�a<��a<c�a<�a<��a<�a<��a<7�a<��a<O�a<ۑa<y�a<�a<��a<R�a<�a<��a<M�a<֎a<q�a<9�a<��a<t�a<)�a<݌a<��a<P�a<�a<��a<k�a<4�a<��a<a<{�a<[�a<!�a<�a<։a<��a<��a<o�a<:�a<@�a<�a<��a<�a<�a<ψa<Јa<͈a<ʈa<Јa<��a<��a<�a<��a<�a<�a<C�a<�  �  _�a<v�a<��a<ĉa<��a<8�a<H�a<��a<��a<�a<)�a<j�a<��a<�a<3�a<�a<Ҍa<�a<s�a<ƍa<�a<��a<Ύa<Y�a<��a<��a<d�a<a<,�a<��a<�a<c�a<�a<M�a<˓a<Q�a<��a<8�a<��a<(�a<��a<�a<��a<�a<��a<
�a<��a<�a<��a<�a<{�a<�a<x�a<��a<d�a<ޝa<P�a<Ğa<E�a<��a<�a<��a<�a<l�a<��a<J�a<��a<�a<@�a<��a<�a<M�a<��a<ڤa<C�a<z�a<ݥa<�a<N�a<��a<ʦa<(�a<M�a<��a<ŧa<��a<,�a<S�a<��a<��a<��a<�a<$�a<L�a<f�a<��a<��a<��a<ҩa<�a<�a<�a<.�a<4�a<e�a<K�a<l�a<u�a<d�a<x�a<i�a<w�a<h�a<z�a<e�a<X�a<^�a<L�a<W�a<6�a</�a<�a<�a<�a<�a<کa<��a<��a<��a<{�a<o�a<0�a<7�a<�a<Ҩa<��a<��a<]�a<+�a< �a<ԧa<��a<u�a<I�a<�a<ݦa<Ȧa<i�a<Z�a<��a<��a<��a<8�a<��a<��a<{�a<�a<٣a<��a<=�a<��a<��a<R�a<�a<��a<O�a<�a<��a<.�a<ݟa<i�a<.�a<��a<K�a<�a<g�a<�a<��a<.�a<��a<F�a<њa<_�a<��a<�a<�a<��a<0�a<��a<6�a<�a<F�a<�a<b�a<��a<|�a<�a<��a<�a<ƒa<E�a<��a<��a<�a<��a<8�a<��a<��a<*�a<Ўa<y�a< �a<a<��a<�a<�a<��a<?�a<��a<��a<v�a<2�a<�a<��a<��a<Y�a<%�a<�a<ωa<ʉa<��a<v�a<Z�a<'�a< �a<��a<��a<وa<�a<ʈa<��a<ˈa<ňa<��a<Ոa<�a<��a<�a<1�a<6�a<�  �  \�a<��a<��a<щa<��a< �a<M�a<��a<��a<�a<<�a<`�a<��a<�a<3�a<��a<Ȍa<�a<}�a<͍a<"�a<�a<ڎa<6�a<��a<�a<p�a<��a<+�a<��a<�a<x�a<�a<E�a<��a<4�a<��a<'�a<��a<�a<��a<#�a<��a<7�a<��a<'�a<��a<�a<��a<�a<��a<��a<��a<�a<z�a<�a<W�a<��a</�a<��a<�a<��a<��a<g�a<ǡa<'�a<��a<�a<a�a<��a<��a<T�a<��a<��a<7�a<y�a<åa<
�a<J�a<��a<�a<�a<f�a<��a<٧a<�a<5�a<j�a<��a<��a<�a<�a<*�a<M�a<m�a<|�a<©a<��a<�a<��a<��a<%�a<(�a<@�a<L�a<Q�a<]�a<i�a<u�a<w�a<��a<s�a<}�a<h�a<a�a<n�a<P�a<F�a<?�a</�a<#�a<(�a<�a<��a<��a<שa<�a<��a<��a<y�a<W�a<5�a<�a<��a<Ѩa<��a<x�a<]�a<E�a< �a<�a<��a<v�a<R�a<�a<�a<��a<t�a<7�a<�a<ɥa<��a<V�a<��a<Ťa<h�a<&�a<٣a<z�a<2�a<�a<��a<A�a<�a<��a<M�a<�a<��a<R�a<ݟa<��a<�a<��a<J�a<ߝa<y�a<�a<��a<�a<ʛa<L�a<ؚa<{�a<�a<��a<�a<��a<%�a<��a<<�a<Öa<b�a<�a<��a<��a<��a<�a<��a<8�a<��a<D�a<ّa<q�a<�a<��a<P�a<�a<��a<(�a<�a<��a<(�a<ٍa<u�a<)�a<ތa<��a<E�a<��a<��a<i�a<T�a<�a<Ҋa<��a<M�a<7�a<��a<ډa<��a<��a<h�a<N�a<9�a<�a<#�a<�a<�a<шa<ƈa<Ոa<��a<��a<Ȉa<Έa<ۈa< �a<	�a<�a<N�a<�  �  L�a<��a<��a<܉a<�a<4�a<r�a<p�a<ۊa<�a<2�a<{�a<��a<��a<%�a<��a<Όa<7�a<n�a<֍a<9�a<l�a<�a<9�a<��a<��a<C�a<Đa<$�a<��a<�a<��a<͒a<[�a<ғa<4�a<̔a<�a<��a<�a<��a<�a<��a<�a<}�a<5�a<��a<:�a<��a<�a<��a<�a<��a<�a<o�a<ӝa<H�a<՞a<;�a<˟a<�a<��a<��a<h�a<�a<%�a<��a<Ӣa<D�a<��a<�a<K�a<��a<�a<�a<��a<ťa<�a<g�a<��a<�a<�a<b�a<��a<��a<�a<(�a<l�a<��a<�a<ըa<�a<>�a<A�a<��a<��a<��a<��a<֩a<�a<�a<!�a<�a<a�a<8�a<o�a<x�a<`�a<��a<S�a<y�a<a�a<|�a<_�a<k�a<]�a<I�a<b�a<7�a<J�a<%�a<�a<�a<�a<��a<ǩa<ȩa<��a<��a<r�a<k�a<Z�a<�a<�a<Ψa<��a<��a<X�a<6�a<�a<�a<��a<��a<C�a<"�a<��a<��a<��a<:�a<�a<åa<b�a<:�a<�a<¤a<T�a<1�a<��a<��a<E�a<�a<��a<+�a<��a<��a<B�a<�a<��a<:�a<��a<��a<
�a<՞a<S�a<֝a<��a<��a<��a<)�a<��a<;�a<ɚa<p�a<�a<��a<�a<��a<%�a<��a<h�a<��a<o�a<ƕa<e�a<�a<z�a<�a<��a<2�a<��a<d�a<ܑa<~�a<!�a<��a<W�a<ԏa<��a< �a<Ǝa<c�a<�a<ڍa<t�a<Z�a<Ќa<��a<Y�a<�a<ҋa<r�a<F�a<�a<��a<��a<e�a<3�a<�a<��a<��a<��a<��a<E�a<I�a<��a<
�a<߈a<�a<Ȉa<Јa<Ĉa<��a<ۈa<��a<�a<ވa<�a<�a<�a<M�a<�  �  \�a<��a<��a<��a<�a<!�a<>�a<��a<��a<��a<*�a<p�a<��a<��a<W�a<��a<׌a<�a<w�a<ˍa<"�a<v�a<Ɏa<8�a<��a<�a<o�a<Րa<.�a<��a<�a<x�a<ߒa<U�a<��a<0�a<��a<2�a<��a<4�a<��a<�a<��a<0�a<��a<�a<��a<�a<z�a<
�a<��a<�a<s�a<��a<j�a<��a<o�a<˞a<H�a<��a<"�a<��a<��a<O�a<��a<'�a<��a<��a<^�a<��a<��a<K�a<��a<�a<;�a<}�a<��a<��a<V�a<��a<ݦa<�a<S�a<��a<էa<�a<A�a<a�a<��a<��a<֨a<�a<)�a<N�a<c�a<��a<��a<ܩa<�a<�a<
�a<�a<1�a<@�a<J�a<=�a<[�a<b�a<�a<�a<��a<t�a<j�a<j�a<u�a<X�a<[�a<A�a<5�a<'�a</�a<�a<�a<��a<�a<שa<ѩa<��a<��a<q�a<X�a<&�a<�a<��a<بa<��a<��a<Z�a<8�a<$�a<֧a<��a<w�a<M�a<�a<�a<��a<d�a<:�a<��a<ҥa<��a<K�a<��a<��a<j�a<&�a<ңa<��a<#�a<ݢa<��a<L�a<�a<��a<E�a<�a<��a<L�a<�a<~�a<�a<��a<2�a<ܝa<v�a<
�a<��a<1�a<��a<^�a<�a<f�a<��a<x�a<�a<��a<$�a<��a<.�a<Öa<Z�a<�a<��a< �a<}�a<�a<��a<)�a<��a<H�a<ёa<b�a<�a<��a<L�a<�a<��a<*�a<ߎa<��a<4�a<Ѝa<x�a<�a<ьa<��a<C�a< �a<��a<}�a<5�a<�a<̊a<��a<_�a<$�a<�a<ډa<��a<s�a<f�a<G�a<C�a<'�a<�a<�a<ۈa<ӈa<ۈa<��a<Ɉa<��a<��a<ƈa<�a<��a<�a<#�a<6�a<�  �  r�a<j�a<��a<��a<�a<B�a<J�a<��a<��a<�a<@�a<m�a<��a<�a<M�a<j�a<�a<�a<��a<ƍa<�a<��a<̎a<a�a<��a<�a<T�a<��a<?�a<��a<	�a<P�a<�a<V�a<��a<U�a<��a<E�a<��a<�a<��a<(�a<��a<�a<��a<��a<��a<#�a<��a<*�a<k�a<*�a<t�a<�a<a�a<؝a<Q�a<��a<Y�a<��a<J�a<u�a<�a<��a<Сa<Q�a<{�a<�a<5�a<��a<�a<J�a<��a<Ǥa<L�a<j�a<ߥa<�a<Q�a<��a<��a<!�a<X�a<��a<��a<�a<'�a<_�a<��a<��a<�a<�a<�a<z�a<_�a<��a<��a<ʩa<ʩa<�a<�a<#�a<L�a<�a<w�a<T�a<|�a<~�a<Y�a<i�a<_�a<��a<w�a<g�a<R�a<J�a<l�a<1�a<Y�a<�a<:�a<�a<�a<��a<�a<�a<��a<��a<��a<��a<y�a<2�a<L�a<ըa<�a<��a<��a<b�a<$�a<�a<��a<��a<q�a<q�a<�a<Ѧa<ߦa<f�a<c�a<�a<��a<s�a<2�a<�a<��a<n�a<��a<ߣa<��a<*�a<�a<y�a<_�a<ϡa<��a<B�a<��a<��a<#�a<ܟa<^�a<6�a<��a<^�a<��a<W�a<0�a<��a<A�a<��a<@�a<Қa<U�a<�a<s�a<9�a<��a<9�a<ӗa<E�a<�a<A�a<��a<V�a<��a<��a<�a<��a<�a<Вa<5�a<��a<w�a<�a<��a<&�a<��a<��a<7�a<ʎa<f�a<�a<͍a<��a<�a<�a<��a<6�a<,�a<��a<��a<�a<�a<��a<��a<`�a<5�a< �a<��a<݉a<��a<��a<c�a<�a<�a<�a<�a<�a<Јa<��a<��a<وa<��a<�a<��a<�a<�a<�a<�a<@�a<�  �  \�a<��a<��a<��a<�a<!�a<>�a<��a<��a<��a<*�a<p�a<��a<��a<W�a<��a<׌a<�a<w�a<ˍa<"�a<v�a<Ɏa<8�a<��a<�a<o�a<Րa<.�a<��a<�a<x�a<ߒa<U�a<��a<0�a<��a<2�a<��a<4�a<��a<�a<��a<0�a<��a<�a<��a<�a<z�a<
�a<��a<�a<s�a<��a<j�a<��a<o�a<˞a<H�a<��a<"�a<��a<��a<O�a<��a<'�a<��a<��a<^�a<��a<��a<K�a<��a<�a<;�a<}�a<��a<��a<V�a<��a<ݦa<�a<S�a<��a<էa<�a<A�a<a�a<��a<��a<֨a<�a<)�a<N�a<c�a<��a<��a<ܩa<�a<�a<
�a<�a<1�a<@�a<J�a<=�a<[�a<b�a<�a<�a<��a<t�a<j�a<j�a<u�a<X�a<[�a<A�a<5�a<'�a</�a<�a<�a<��a<�a<שa<ѩa<��a<��a<q�a<X�a<&�a<�a<��a<بa<��a<��a<Z�a<8�a<$�a<֧a<��a<w�a<M�a<�a<�a<��a<d�a<:�a<��a<ҥa<��a<K�a<��a<��a<j�a<&�a<ңa<��a<#�a<ݢa<��a<L�a<�a<��a<E�a<�a<��a<L�a<�a<~�a<�a<��a<2�a<ܝa<v�a<
�a<��a<1�a<��a<^�a<�a<f�a<��a<x�a<�a<��a<$�a<��a<.�a<Öa<Z�a<�a<��a< �a<}�a<�a<��a<)�a<��a<H�a<ёa<b�a<�a<��a<L�a<�a<��a<*�a<ߎa<��a<4�a<Ѝa<x�a<�a<ьa<��a<C�a< �a<��a<}�a<5�a<�a<̊a<��a<_�a<$�a<�a<ډa<��a<s�a<f�a<G�a<C�a<'�a<�a<�a<ۈa<ӈa<ۈa<��a<Ɉa<��a<��a<ƈa<�a<��a<�a<#�a<6�a<�  �  L�a<��a<��a<܉a<�a<4�a<r�a<p�a<ۊa<�a<2�a<{�a<��a<��a<%�a<��a<Όa<7�a<n�a<֍a<9�a<l�a<�a<9�a<��a<��a<C�a<Đa<$�a<��a<�a<��a<͒a<[�a<ғa<4�a<̔a<�a<��a<�a<��a<�a<��a<�a<}�a<5�a<��a<:�a<��a<�a<��a<�a<��a<�a<o�a<ӝa<H�a<՞a<;�a<˟a<�a<��a<��a<h�a<�a<%�a<��a<Ӣa<D�a<��a<�a<K�a<��a<�a<�a<��a<ťa<�a<g�a<��a<�a<�a<b�a<��a<��a<�a<(�a<l�a<��a<�a<ըa<�a<>�a<A�a<��a<��a<��a<��a<֩a<�a<�a<!�a<�a<a�a<8�a<o�a<x�a<`�a<��a<S�a<y�a<a�a<|�a<_�a<k�a<]�a<I�a<b�a<7�a<J�a<%�a<�a<�a<�a<��a<ǩa<ȩa<��a<��a<r�a<k�a<Z�a<�a<�a<Ψa<��a<��a<X�a<6�a<�a<�a<��a<��a<C�a<"�a<��a<��a<��a<:�a<�a<åa<b�a<:�a<�a<¤a<T�a<1�a<��a<��a<E�a<�a<��a<+�a<��a<��a<B�a<�a<��a<:�a<��a<��a<
�a<՞a<S�a<֝a<��a<��a<��a<)�a<��a<;�a<ɚa<p�a<�a<��a<�a<��a<%�a<��a<h�a<��a<o�a<ƕa<e�a<�a<z�a<�a<��a<2�a<��a<d�a<ܑa<~�a<!�a<��a<W�a<ԏa<��a< �a<Ǝa<c�a<�a<ڍa<t�a<Z�a<Ќa<��a<Y�a<�a<ҋa<r�a<F�a<�a<��a<��a<e�a<3�a<�a<��a<��a<��a<��a<E�a<I�a<��a<
�a<߈a<�a<Ȉa<Јa<Ĉa<��a<ۈa<��a<�a<ވa<�a<�a<�a<M�a<�  �  \�a<��a<��a<щa<��a< �a<M�a<��a<��a<�a<<�a<`�a<��a<�a<3�a<��a<Ȍa<�a<}�a<͍a<"�a<�a<ڎa<6�a<��a<�a<p�a<��a<+�a<��a<�a<x�a<�a<E�a<��a<4�a<��a<'�a<��a<�a<��a<#�a<��a<7�a<��a<'�a<��a<�a<��a<�a<��a<��a<��a<�a<z�a<�a<W�a<��a</�a<��a<�a<��a<��a<g�a<ǡa<'�a<��a<�a<a�a<��a<��a<T�a<��a<��a<7�a<y�a<åa<
�a<J�a<��a<�a<�a<f�a<��a<٧a<�a<5�a<j�a<��a<��a<�a<�a<*�a<M�a<m�a<|�a<©a<��a<�a<��a<��a<%�a<(�a<@�a<L�a<Q�a<]�a<i�a<u�a<w�a<��a<s�a<}�a<h�a<a�a<n�a<P�a<F�a<?�a</�a<#�a<(�a<�a<��a<��a<שa<�a<��a<��a<y�a<W�a<5�a<�a<��a<Ѩa<��a<x�a<]�a<E�a< �a<�a<��a<v�a<R�a<�a<�a<��a<t�a<7�a<�a<ɥa<��a<V�a<��a<Ťa<h�a<&�a<٣a<z�a<2�a<�a<��a<A�a<�a<��a<M�a<�a<��a<R�a<ݟa<��a<�a<��a<J�a<ߝa<y�a<�a<��a<�a<ʛa<L�a<ؚa<{�a<�a<��a<�a<��a<%�a<��a<<�a<Öa<b�a<�a<��a<��a<��a<�a<��a<8�a<��a<D�a<ّa<q�a<�a<��a<P�a<�a<��a<(�a<�a<��a<(�a<ٍa<u�a<)�a<ތa<��a<E�a<��a<��a<i�a<T�a<�a<Ҋa<��a<M�a<7�a<��a<ډa<��a<��a<h�a<N�a<9�a<�a<#�a<�a<�a<шa<ƈa<Ոa<��a<��a<Ȉa<Έa<ۈa< �a<	�a<�a<N�a<�  �  _�a<v�a<��a<ĉa<��a<8�a<H�a<��a<��a<�a<)�a<j�a<��a<�a<3�a<�a<Ҍa<�a<s�a<ƍa<�a<��a<Ύa<Y�a<��a<��a<d�a<a<,�a<��a<�a<c�a<�a<M�a<˓a<Q�a<��a<8�a<��a<(�a<��a<�a<��a<�a<��a<
�a<��a<�a<��a<�a<{�a<�a<x�a<��a<d�a<ޝa<P�a<Ğa<E�a<��a<�a<��a<�a<l�a<��a<J�a<��a<�a<@�a<��a<�a<M�a<��a<ڤa<C�a<z�a<ݥa<�a<N�a<��a<ʦa<(�a<M�a<��a<ŧa<��a<,�a<S�a<��a<��a<��a<�a<$�a<L�a<f�a<��a<��a<��a<ҩa<�a<�a<�a<.�a<4�a<e�a<K�a<l�a<u�a<d�a<x�a<i�a<w�a<h�a<z�a<e�a<X�a<^�a<L�a<W�a<6�a</�a<�a<�a<�a<�a<کa<��a<��a<��a<{�a<o�a<0�a<7�a<�a<Ҩa<��a<��a<]�a<+�a< �a<ԧa<��a<u�a<I�a<�a<ݦa<Ȧa<i�a<Z�a<��a<��a<��a<8�a<��a<��a<{�a<�a<٣a<��a<=�a<��a<��a<R�a<�a<��a<O�a<�a<��a<.�a<ݟa<i�a<.�a<��a<K�a<�a<g�a<�a<��a<.�a<��a<F�a<њa<_�a<��a<�a<�a<��a<0�a<��a<6�a<�a<F�a<�a<b�a<��a<|�a<�a<��a<�a<ƒa<E�a<��a<��a<�a<��a<8�a<��a<��a<*�a<Ўa<y�a< �a<a<��a<�a<�a<��a<?�a<��a<��a<v�a<2�a<�a<��a<��a<Y�a<%�a<�a<ωa<ʉa<��a<v�a<Z�a<'�a< �a<��a<��a<وa<�a<ʈa<��a<ˈa<ňa<��a<Ոa<�a<��a<�a<1�a<6�a<�  �  ��a<v�a<��a<މa<�a<(�a<Y�a<w�a<��a<��a<"�a<p�a<��a<�a<<�a<��a<ǌa<&�a<f�a<ԍa<!�a<z�a<ݎa<7�a<��a<�a<\�a<Ða<S�a<��a<��a<y�a<�a<]�a<̓a<3�a<��a<0�a<��a<%�a<��a<.�a<��a<�a<��a<�a<��a<�a<��a<��a<��a<��a<s�a<�a<c�a<�a<]�a<Ǟa<8�a<��a<�a<��a<�a<c�a<ša<"�a<��a<�a<B�a<��a<�a<I�a<��a<��a<<�a<��a<ĥa<�a<\�a<��a<�a<�a<Q�a<��a<˧a<��a<F�a<S�a<��a<��a<�a< �a<5�a<=�a<k�a<~�a<��a<éa<ةa<ީa<�a<�a<1�a<<�a<<�a<]�a<d�a<U�a<|�a<v�a<k�a<��a<y�a<f�a<k�a<f�a<]�a<W�a<2�a<B�a<5�a<%�a<�a<��a<�a<��a<��a<��a<��a<c�a<_�a<A�a<�a<��a<ۨa<��a<��a<L�a<0�a<	�a<קa<��a<��a<<�a<!�a<�a<��a<w�a<8�a<�a<֥a<{�a<:�a<�a<��a<d�a<'�a<ۣa<��a<?�a<�a<��a<J�a<�a<��a<B�a<��a<��a<1�a<�a<s�a<�a<��a<I�a<ѝa<z�a<��a<��a<*�a<��a<P�a<ޚa<b�a<�a<z�a<�a<��a<�a<��a<:�a<��a<M�a<��a<c�a<�a<��a<�a<��a<7�a<��a<O�a<ۑa<y�a<�a<��a<R�a<�a<��a<M�a<֎a<q�a<9�a<��a<t�a<)�a<݌a<��a<P�a<�a<��a<k�a<4�a<��a<a<{�a<[�a<!�a<�a<։a<��a<��a<o�a<:�a<@�a<�a<��a<�a<�a<ψa<Јa<͈a<ʈa<Јa<��a<��a<�a<��a<�a<�a<C�a<�  �  [�a<��a<��a<߉a<�a<�a<[�a<|�a<��a<�a<:�a<q�a<��a<��a<(�a<��a<��a<.�a<s�a<ōa<�a<x�a<�a<4�a<��a<
�a<e�a<אa<0�a<��a<�a<��a<�a<R�a<ٓa<?�a<Ŕa<"�a<ȕa<$�a<��a<�a<��a<&�a<��a<-�a<��a<�a<��a<�a<��a<�a<��a<�a<b�a<ޝa<Q�a<ʞa<(�a<şa<�a<��a<�a<i�a<̡a<.�a<��a<�a<Q�a<��a<��a<Y�a<��a<�a<-�a<��a<ҥa< �a<Z�a<��a<��a<�a<`�a<��a<֧a<��a<8�a<t�a<��a<��a<ݨa<��a<%�a<A�a<|�a<n�a<��a<��a<ݩa<ܩa<�a<(�a< �a<7�a<B�a<`�a<`�a<v�a<��a<n�a<��a<r�a<t�a<p�a<u�a<y�a<H�a<b�a<@�a<M�a<�a<2�a<#�a<��a<�a<֩a<Щa<��a<��a<��a<V�a<C�a<�a<�a<ɨa<��a<��a<C�a<8�a<��a<ާa<��a<��a<H�a<�a<ަa<��a<��a<5�a<�a<Υa<��a<M�a<��a<��a<j�a<>�a<ڣa<��a<L�a<�a<��a<;�a<�a<��a<N�a<�a<��a<A�a<ڟa<��a<�a<��a<O�a<؝a<w�a<��a<��a<�a<��a<E�a<Қa<e�a<ݙa<��a<�a<��a<�a<��a<A�a<ʖa<g�a<�a<s�a<�a<��a<�a<��a<M�a<��a<\�a<�a<��a<�a<��a<g�a<�a<��a<-�a<�a<|�a<+�a<�a<x�a<1�a<ٌa<��a<@�a<�a<ɋa<[�a<:�a<�a<Ȋa<z�a<W�a<:�a<�a<щa<��a<��a<k�a<[�a<F�a<�a<�a<�a<�a<؈a<ڈa<��a<��a<ۈa<Ɉa<�a<ֈa<
�a<�a<$�a<B�a<�  �  W�a<��a<��a<��a<�a< �a<E�a<��a<��a<ߊa<&�a<h�a<��a<�a<�a<~�a<Ȍa<�a<l�a<��a<$�a<��a<͎a<<�a<��a<�a<e�a<Ӑa<)�a<��a<�a<x�a<�a<Q�a<ٓa<P�a<��a<0�a<��a<"�a<��a<!�a<��a<�a<��a<�a<��a<�a<��a<#�a<z�a<�a<y�a<�a<_�a<ѝa<C�a<��a<4�a<��a<�a<��a<	�a<n�a<��a<C�a<��a<�a<J�a<��a<��a<b�a<��a<�a<>�a<��a<�a<&�a<Z�a<��a<�a<�a<d�a<��a<Чa<��a<#�a<_�a<��a<��a<��a<
�a<�a<A�a<j�a<�a<��a<��a<ѩa<�a<��a<�a<�a</�a<g�a<J�a<Y�a<~�a<[�a<t�a<|�a<r�a<x�a<��a<f�a<r�a<Z�a<[�a<U�a<E�a<*�a<0�a<�a<�a<�a<ҩa<ͩa<��a<��a<��a<W�a<-�a<:�a<�a<��a<��a<��a<X�a<,�a<�a<ӧa<��a<t�a<B�a<�a<�a<Ŧa<g�a<>�a<�a<��a<��a<I�a<�a<��a<x�a<&�a<�a<��a<K�a<��a<��a<J�a<��a<��a<_�a<�a<��a<9�a<ӟa<m�a<)�a<��a<K�a<��a<f�a<��a<��a< �a<��a<9�a<Ěa<X�a<�a<��a<��a<��a<7�a<��a<3�a<ߖa<L�a<וa<k�a<��a<�a<$�a<��a<2�a<��a<Y�a<��a<��a<�a<��a<N�a<�a<��a<(�a<ڎa<z�a<�a<͍a<��a<�a<�a<��a<4�a<�a<��a<l�a<-�a<��a<��a<��a<S�a<$�a<�a<ɉa<͉a<��a<d�a<c�a<�a<�a<�a<��a<�a<�a<ˈa<؈a<ǈa<Ԉa<ވa<�a<�a<�a<
�a<6�a<F�a<�  �  ��a<z�a<��a<̉a<�a<'�a<F�a<�a<��a<��a<�a<\�a<��a<�a<?�a<r�a<ˌa<�a<h�a<͍a<�a<z�a<͎a<<�a<��a<�a<k�a<Đa<O�a<��a<�a<z�a<�a<_�a<ғa<A�a<��a<<�a<��a<1�a<��a<(�a<��a<�a<��a<�a<��a<�a<��a<�a<w�a<�a<\�a<�a<S�a<ޝa<X�a<��a<;�a<��a<�a<��a<�a<]�a<��a<0�a<��a<�a<C�a<��a<�a<N�a<��a<��a<K�a<��a<ҥa<�a<a�a<��a<�a<&�a<T�a<��a<̧a< �a<H�a<Q�a<��a<��a<٨a<��a<(�a<B�a<S�a<��a<��a<ũa<̩a<ݩa<��a<��a<2�a<(�a<@�a<K�a<b�a<`�a<g�a<��a<m�a<��a<s�a<s�a<q�a<g�a<f�a<V�a<L�a<?�a<:�a<(�a<�a<�a<�a<��a<��a<ȩa<��a<o�a<^�a<.�a<�a<�a<بa<��a<u�a<O�a<#�a<�a<ȧa<��a<d�a<=�a<�a<Ҧa<��a<g�a<>�a<�a<ӥa<��a<:�a<�a<��a<x�a<(�a<�a<��a<E�a<�a<��a<V�a<��a<��a<L�a<��a<��a<.�a<��a<k�a<�a<��a<B�a<ӝa<c�a<
�a<z�a<&�a<��a<F�a<ٚa<O�a<�a<a�a<�a<��a<�a<��a<3�a<̖a<F�a<��a<d�a<
�a<��a<�a<��a<6�a<Βa<V�a<�a<��a<�a<��a<Q�a<��a<��a<H�a<׎a<}�a<;�a<��a<}�a<�a<Ԍa<}�a<C�a<�a<��a<r�a<%�a<�a<��a<z�a<N�a<�a<�a<a<��a<��a<m�a<E�a<+�a<;�a<��a<�a<�a<܈a<׈a<Έa<ӈa<ψa<ֈa<ވa<�a< �a<�a<,�a<@�a<�  �  f�a<��a<��a<Љa<��a<%�a<k�a<}�a<Êa<�a<#�a<g�a<��a<ۋa<%�a<m�a<��a<!�a<a�a<��a<$�a<w�a<��a<<�a<��a<��a<b�a<ʐa<:�a<��a<�a<��a<�a<k�a<�a<D�a<ߔa<.�a<��a<0�a<��a<#�a<��a<�a<��a<%�a<��a<#�a<��a<�a<��a<��a<x�a<�a<Q�a<˝a<?�a<��a<1�a<��a<�a<��a<�a<f�a<ܡa<1�a<��a<�a<K�a<��a<��a<Y�a<��a<�a<8�a<��a<٥a<&�a<r�a<��a<�a<"�a<e�a<��a<ϧa<��a<+�a<l�a<��a<Шa<بa<�a<#�a<7�a<k�a<t�a<��a<��a<©a<ԩa<��a<�a<�a<F�a<@�a<k�a<i�a<p�a<t�a<p�a<v�a<{�a<y�a<z�a<}�a<e�a<_�a<t�a<K�a<[�a<6�a<�a<&�a<�a<��a<�a<éa<��a<��a<|�a<\�a<S�a<�a< �a<èa<��a<�a<D�a<�a<�a<§a<��a<{�a<6�a<�a<�a<��a<��a<>�a<�a<¥a<��a<@�a<�a<��a<r�a<9�a<գa<��a<U�a<�a<Ģa<H�a<�a<��a<R�a<�a<��a<:�a<՟a<��a<�a<��a<O�a<ӝa<x�a<��a<��a< �a<��a<3�a<��a<N�a<�a<�a<�a<��a<�a<��a<Q�a<͖a<b�a<ܕa<m�a<��a<��a<�a<��a<B�a<��a<t�a<�a<��a<-�a<��a<b�a<�a<��a<6�a<َa<{�a<�a<ۍa<}�a<C�a<ӌa<��a<>�a<�a<��a<a�a< �a<�a<��a<q�a<R�a<#�a<�a<�a<��a<��a<t�a<U�a<8�a<�a<�a<��a<�a<�a<�a<̈a<̈a<�a<Ԉa<��a<�a<��a<"�a<,�a<H�a<�  �  N�a<��a<��a<ʉa<�a< �a<R�a<p�a<a<֊a<-�a<Q�a<��a<�a<�a<��a<��a<�a<j�a<��a<"�a<d�a<ێa<�a<��a<��a<��a<�a<(�a<ȑa<�a<��a<��a<`�a<ѓa<:�a<Ҕa<7�a<Еa<$�a<Ŗa<3�a<��a<Q�a<��a<*�a<��a<��a<z�a<��a<��a<�a<|�a<Μa<o�a<՝a<D�a<Ӟa<�a<��a<�a<��a<�a<L�a<��a<�a<��a<�a<z�a<��a<�a<v�a<��a<�a<C�a<��a<ʥa<�a<f�a<��a<��a<�a<��a<��a<ܧa<#�a<&�a<z�a<k�a<��a<Ǩa<��a<�a<:�a<_�a<a�a<��a<��a<թa<�a<�a<�a<
�a<B�a<6�a<P�a<>�a<n�a<q�a<x�a<��a<e�a<��a<�a<o�a<��a<c�a<g�a<=�a<L�a<5�a<:�a<�a<�a<�a<ɩa<�a<��a<��a<��a<7�a<:�a<�a<��a<��a<��a<i�a<L�a<4�a<�a<�a<��a<n�a<@�a<�a<�a<��a<u�a<�a<�a<��a<��a<X�a<�a<�a<f�a<8�a<�a<��a<D�a<�a<��a<P�a<�a<��a<k�a<�a<��a<m�a<ԟa<��a<�a<��a<2�a<ʝa<s�a<�a<��a<�a<��a<=�a<Śa<m�a<͙a<}�a<��a<��a<�a<��a<1�a<��a<l�a<ٕa<��a<��a<��a<8�a<��a<T�a<ǒa<h�a<�a<{�a< �a<��a<g�a<�a<��a<+�a<�a<��a<�a<�a<Y�a<*�a<a<��a<2�a<�a<��a<N�a<A�a<�a<��a<��a<9�a<.�a<މa<݉a<��a<��a<I�a<S�a<5�a< �a<3�a<�a<�a<�a<Ԉa<�a<Јa<߈a<ǈa<�a<�a<�a<�a<-�a<d�a<�  �  a�a<p�a<��a<Ɖa<	�a<.�a<\�a<}�a<��a<�a<-�a<Z�a<��a<ыa<�a<j�a<Ȍa<�a<x�a<��a<�a<x�a<�a<E�a<��a<��a<_�a<��a<7�a<��a<�a<w�a<��a<a�a<�a<f�a<��a<C�a<��a<2�a<��a<'�a<��a<�a<��a<�a<��a<#�a<��a<�a<|�a<��a<o�a<�a<Z�a<��a<4�a<��a<1�a<��a<�a<��a<�a<h�a<ۡa<<�a<��a<�a<>�a<��a<��a<W�a<��a<�a<Q�a<��a<�a<3�a<d�a<��a<ߦa<(�a<c�a<��a<��a<��a<+�a<f�a<��a<Ǩa<ܨa<��a<�a<P�a<V�a<��a<��a<��a<��a<�a<�a<�a<!�a<+�a<A�a<_�a<j�a<y�a<l�a<t�a<f�a<u�a<z�a<z�a<u�a<j�a<j�a<[�a<q�a<K�a<9�a<,�a<�a<�a<��a<ܩa<��a<��a<��a<��a<e�a<D�a<�a<�a<ɨa<��a<s�a<Q�a<�a<�a<��a<��a<f�a<M�a<
�a<զa<��a<��a<F�a<�a<��a<~�a<*�a<�a<��a<z�a<%�a<�a<��a<U�a<�a<��a<]�a<��a<��a<Q�a<��a<��a<-�a<ןa<{�a<$�a<��a<O�a<ԝa<h�a<�a<��a<�a<��a<$�a<��a<S�a<�a<s�a<�a<��a<�a<��a<P�a<ؖa<Y�a<ەa<_�a<�a<��a<�a<��a</�a<Ԓa<[�a<	�a<��a<�a<��a<N�a<��a<��a<4�a<��a<t�a<�a<ԍa<��a<:�a<׌a<��a<8�a<�a<��a<m�a< �a<��a<��a<��a<H�a<&�a<�a<ŉa<��a<��a<u�a<^�a<0�a<�a<��a<�a<�a<�a<ڈa<шa<؈a<Ԉa<��a<�a<�a<�a<�a<3�a<G�a<�  �  ��a<o�a<��a<��a<݊a<�a<+�a<l�a<��a<�a<�a<?�a<��a<��a<7�a<I�a<��a<��a<S�a<��a<��a<S�a<��a<)�a<r�a<ܐa<P�a<��a<Q�a<X�a<�a<M�a<Гa<@�a<��a<@�a<��a<4�a<j�a<�a<f�a<��a<��a<�a<r�a<˙a<f�a<��a<F�a<��a<'�a<��a<(�a<��a<	�a<��a<	�a<`�a<�a<R�a<Πa<%�a<��a<�a<Y�a<�a<)�a<��a<��a<s�a<��a<�a<s�a<��a<�a<4�a<��a<Цa<�a<a�a<�a<�a<�a<s�a<��a<��a<�a<��a<M�a<@�a<��a<��a<ǩa<��a<�a<2�a<-�a<�a<m�a<��a<��a<��a<�a<̪a<�a<��a<	�a<�a<�a<1�a<,�a<j�a<�a<-�a<,�a<�a<?�a<��a<!�a<�a<�a<֪a<Ϫa<ƪa<��a<ժa<x�a<t�a<>�a<$�a<�a<کa<ȩa<��a<��a<O�a<!�a<�a<ʨa<Ψa<i�a<W�a<�a<��a<ça<��a<Q�a<�a<��a<��a<q�a<A�a<��a<�a<G�a<>�a<Ҥa<��a<N�a<��a<ɣa<K�a<-�a<��a<u�a<�a<��a<y�a<��a<��a<�a<ӟa<K�a<�a<��a<�a<��a<D�a<ڜa<[�a<��a<��a<�a<��a<2�a<͙a<F�a<��a<m�a<�a<��a<�a<��a<C�a<�a<p�a<͔a<��a<��a<��a<,�a<�a<f�a<��a<��a< �a<�a<M�a<E�a<��a<e�a<�a<��a<r�a<�a<��a<m�a<�a<ތa<��a<Y�a<��a<��a<��a<j�a<-�a<�a<��a<��a<��a<g�a<P�a<8�a<�a<�a<��a<&�a<ŉa<҉a<Ήa<��a<�a<��a<�a<ȉa< �a<�a<�a<'�a<�a<�  �  R�a<[�a<��a<��a<�a<�a<G�a<l�a<��a<Ջa<�a<H�a<��a<ǌa<�a<X�a<��a<��a<U�a<��a< �a<_�a<ɏa<�a<��a<ސa<J�a<��a<�a<{�a<��a<Q�a<֓a<>�a<��a<,�a<��a<�a<��a<�a<��a<��a<\�a<ޘa<i�a<�a<h�a<ߚa<\�a<ța<D�a<��a<3�a<��a<�a<��a<�a<t�a<�a<^�a<Ơa<>�a<��a<�a<~�a<�a<?�a<��a<�a<A�a<��a<�a<a�a<��a<��a<.�a<��a<ʦa<�a<_�a<��a<ܧa<�a<L�a<c�a<��a<ߨa<�a<=�a<k�a<��a<��a<ϩa<��a<�a</�a<A�a<h�a<u�a<��a<��a<Īa<Ҫa<�a<��a<�a<�a<%�a<#�a<,�a<�a<#�a<0�a<7�a<%�a<�a<$�a<��a<�a<�a<��a<ߪa<Ȫa<ɪa<��a<��a<d�a<h�a<G�a<5�a<�a<��a<ǩa<��a<}�a<Z�a<*�a<�a<Ѩa<��a<y�a<S�a<$�a<��a<��a<��a<\�a<2�a<�a<��a<s�a<;�a<ޥa<��a<i�a<6�a<פa<��a<L�a<�a<��a<I�a<�a<��a<g�a<�a<��a<:�a<�a<��a<.�a<֟a<m�a<�a<��a<)�a<��a<O�a<ڜa<l�a<��a<��a<�a<��a<>�a<ƙa<_�a<�a<��a<�a<��a<#�a<��a<5�a<��a<i�a<�a<��a<�a<��a<&�a<ђa<_�a<��a<��a<,�a<ݐa<n�a<�a<��a<_�a<	�a<��a<b�a<�a<��a<o�a<"�a<ߌa<��a<V�a<�a<ދa<��a<q�a<6�a<�a<�a<��a<��a<�a<_�a<G�a<#�a<�a<�a<މa<މa<܉a<ǉa<a<Ήa<��a<҉a<ĉa<�a<�a< �a<*�a<6�a<�  �  G�a<��a<��a<��a<�a<��a<H�a<Z�a<��a<ċa<�a<A�a<��a<ӌa<�a<d�a<��a<��a<K�a<��a<
�a<R�a<ˏa<��a<��a<Րa<Z�a<Ǒa<�a<��a<�a<\�a<Гa<8�a<��a<)�a<��a<�a<��a<�a<y�a<�a<i�a<�a<_�a<�a<I�a<Ԛa<R�a<��a<O�a<��a<4�a<��a<�a<��a<��a<w�a<֟a<_�a<��a<B�a<��a<�a<y�a<��a<H�a<��a<�a<X�a<��a<�a<E�a<��a<�a<@�a<��a<Цa<�a<V�a<��a<ça<�a<<�a<��a<ƨa<Өa<�a<�a<o�a<��a<��a<ϩa<�a<�a<�a<L�a<P�a<~�a<��a<��a<êa<��a<��a<�a<�a< �a<�a<"�a<)�a<K�a<�a<?�a<!�a<�a<.�a<�a<�a<�a<�a<�a<�a<ɪa<��a<��a<��a<��a<j�a<E�a<-�a<��a<��a<��a<��a<l�a<X�a<#�a<��a<ݨa<��a<��a<F�a<�a<�a<��a<��a<P�a<4�a<˦a<��a<j�a<K�a<�a<��a<z�a<�a<�a<��a<F�a<�a<��a<`�a<��a<Ģa<O�a<�a<��a<G�a<�a<��a<3�a<��a<a�a<��a<��a<4�a<��a<Q�a<ʜa<h�a<��a<��a<�a<��a<?�a<��a<c�a<ޘa<t�a<�a<x�a<,�a<��a<^�a<Еa<c�a<�a<l�a<�a<��a<8�a<Вa<f�a<��a<��a<<�a<Őa<|�a<�a<͏a<y�a<��a<��a<;�a<�a<��a<p�a<#�a<Ќa<��a<D�a<�a<ǋa<��a<g�a<,�a<�a<͊a<͊a<��a<�a<G�a<8�a<#�a<�a<�a<ډa<�a<ǉa<��a<҉a<��a<щa<҉a<މa<ډa<��a<�a<�a<I�a<�  �  \�a<m�a<{�a<��a<�a<�a<F�a<d�a<��a<Ћa<�a<L�a<��a<Ќa<�a<b�a<��a<��a<P�a<��a<�a<V�a<��a<!�a<��a<ؐa<-�a<��a<�a<y�a<�a<_�a<ēa<0�a<��a<�a<��a<�a<��a<�a<u�a<��a<r�a<ݘa<V�a<�a<g�a<ؚa<\�a<̛a<;�a<��a<*�a<��a<�a<��a<�a<w�a<�a<[�a<Ƞa<2�a<��a<�a<y�a<�a<J�a<��a<�a<T�a<��a<��a<U�a<��a<�a<9�a<��a<Цa<
�a<N�a<��a<ӧa<�a<B�a<x�a<��a<Ҩa<�a<@�a<b�a<��a<��a<ɩa<�a<�a<7�a<L�a<d�a<~�a<��a<��a<��a<ͪa<�a<�a<�a<�a<(�a<(�a<�a<#�a<5�a<'�a<$�a<0�a<�a<�a<�a<��a<��a<�a<۪a<٪a<��a<��a<��a<v�a<H�a<M�a<9�a<�a<��a<��a<��a<w�a<S�a<.�a<�a<٨a<��a<��a<_�a<$�a<�a<��a<��a<T�a<%�a<�a<��a<m�a<�a<��a<��a<h�a<+�a<�a<��a<?�a< �a<��a<U�a<��a<��a<`�a<��a<��a<P�a<�a<��a<8�a<ԟa<e�a<�a<��a< �a<��a<F�a<�a<l�a<��a<��a<�a<��a<;�a<Ǚa<S�a<�a<~�a<	�a<��a<.�a<��a<,�a<̕a<Z�a<�a<|�a<
�a<��a<1�a<˒a<f�a<��a<��a<3�a<Րa<k�a<�a<��a<I�a<��a<��a<e�a<�a<��a<}�a<�a<ڌa<��a<^�a<�a<ۋa<��a<t�a<>�a<	�a<܊a<��a<��a<��a<S�a<I�a<)�a<�a<�a<��a<Չa<ʉa<҉a<a<��a<Éa<��a<։a<؉a<�a<�a<�a<0�a<�  �  `�a<`�a<��a<ʊa<֊a<�a<.�a<r�a<��a<�a<�a<P�a<��a<��a<!�a<L�a<��a<��a<c�a<��a<��a<^�a<��a<(�a<f�a<��a<T�a<��a<�a<p�a<��a<N�a<֓a<;�a<��a<"�a<��a<$�a<��a<�a<��a<�a<r�a<�a<��a<יa<^�a<͚a<F�a<Λa<2�a<͜a<�a<��a<�a<��a<�a<s�a<��a<I�a<ߠa<-�a<��a<	�a<k�a<ߢa<-�a<ģa<��a<U�a<��a<�a<d�a<��a<�a<3�a<��a<ʦa<�a<a�a<��a<�a<�a<K�a<t�a<��a< �a<��a<C�a<U�a<��a<��a<ɩa<�a<�a<4�a<8�a<h�a<n�a<��a<��a<��a<�a<٪a<��a<��a<�a<�a<(�a<@�a<�a<7�a<�a</�a<'�a<�a<+�a<	�a<�a<��a<��a<�a<˪a<ªa<��a<��a<i�a<w�a<V�a<�a<�a<ݩa<Ωa<��a<��a<^�a<1�a<	�a<Ĩa<��a<m�a<[�a<�a<�a<§a<��a<\�a<�a<��a<��a<��a<E�a<�a<��a<_�a<3�a<Ԥa<��a<I�a<��a<��a<S�a<�a<��a<i�a<�a<��a<P�a<�a<��a<$�a<˟a<[�a<�a<��a<�a<Νa<9�a<�a<o�a<��a<��a<�a<��a<*�a<ޙa<M�a<�a<r�a<��a<��a<�a<֖a<:�a<̕a<_�a<�a<��a<�a<��a<*�a<Ȓa<_�a<��a<��a<%�a<�a<j�a<�a<��a<i�a<*�a<��a<i�a< �a<��a<p�a<�a<�a<��a<\�a<�a<ދa<��a<s�a<E�a<�a<��a<��a<��a<j�a<T�a<3�a<)�a<%�a<�a<�a<̉a<Չa<ʉa<a<Չa<��a<̉a<ωa<�a<�a<�a<"�a<&�a<�  �  T�a<{�a<��a<��a<��a<"�a<>�a<q�a<��a<׋a<�a<E�a<��a<ٌa<�a<k�a<��a<��a<X�a<��a<�a<`�a<ŏa<(�a<v�a<Ԑa<D�a<��a<�a<��a<�a<K�a<˓a<7�a<��a<�a<��a<�a<��a<�a<z�a<�a<v�a<��a<c�a<ՙa<a�a<�a<J�a<Ǜa<B�a<��a<0�a<��a<&�a<��a<�a<��a<�a<[�a<Рa<<�a<��a<	�a<��a<�a<3�a<��a<�a<^�a<��a<�a<I�a<��a<�a<8�a<~�a<��a<�a<S�a<��a<̧a<�a<=�a<��a<��a<Ԩa<�a<B�a<p�a<��a<��a<ԩa<��a<
�a<3�a<T�a<c�a<��a<��a<��a<Īa<ժa<�a<��a<�a<'�a<�a<�a<'�a<1�a</�a<+�a<,�a<�a< �a<�a<	�a<�a<�a<�a<ުa<��a<��a<��a<��a<��a<b�a<8�a<'�a<�a<�a<ͩa<��a<~�a<[�a<'�a<�a<�a<��a<��a<]�a<�a<��a<ħa<��a<]�a</�a<��a<��a<i�a<5�a<�a<��a<o�a<$�a<Ѥa<��a<E�a<�a<��a<V�a<��a<��a<L�a<�a<��a<T�a<��a<��a<!�a<Οa<v�a<��a<��a<(�a<��a<L�a<ڜa<x�a<��a<��a<)�a<��a<<�a<ϙa<]�a<�a<q�a<�a<��a<�a<��a<G�a<Օa<R�a<�a<q�a<�a<��a<0�a<Òa<V�a<��a<��a<'�a<ΐa<u�a<�a<Ïa<c�a<��a<��a<g�a<�a<��a<l�a<'�a<�a<��a<Z�a<!�a<ًa<��a<r�a<2�a<�a<�a<��a<��a<u�a<n�a<;�a<�a<�a<��a<�a<ىa<щa<��a<ĉa<��a<��a<ˉa<Ήa<܉a<�a<��a<�a<7�a<�  �  A�a<t�a<��a<ˊa<��a<�a<@�a<`�a<��a<׋a<�a<K�a<��a<݌a<�a<p�a<��a<	�a<O�a<��a<�a<N�a<��a<�a<��a<��a<9�a<��a<�a<��a<ޒa<Z�a<��a<=�a<��a<	�a<��a<��a<��a<�a<��a<�a<b�a<�a<S�a<�a<S�a<Ԛa<O�a<��a<W�a<��a<=�a<��a<-�a<��a<��a<��a<ߟa<j�a<��a<N�a<��a<�a<u�a<͢a<g�a<��a<��a<L�a<��a<�a<C�a<��a<ݥa<F�a<r�a<��a<�a<?�a<��a<��a<�a<4�a<u�a<��a<֨a<1�a<'�a<c�a<|�a<��a<�a<�a<�a<'�a<]�a<U�a<��a<��a<��a<Ȫa<Ъa<��a<�a<�a<�a<�a<;�a<�a<+�a<�a<2�a<)�a<�a<�a<
�a<�a<�a<��a<�a<Ӫa<Ūa<��a<��a<��a<|�a<T�a<X�a<7�a<�a<�a<��a<��a<�a<Z�a<,�a<�a<�a<��a<��a<P�a<.�a<�a<ϧa<��a<L�a<(�a<ݦa<Цa<u�a<+�a<�a<��a<~�a<�a<ߤa<��a<K�a<��a<��a<d�a<��a<��a<L�a<�a<��a<@�a<�a<}�a<U�a<��a<b�a<��a<��a<<�a<��a<Y�a<Ӝa<�a<��a<��a<0�a<��a<J�a<��a<o�a<��a<s�a<�a<��a<K�a<��a<:�a<Õa<Q�a<��a<k�a<�a<��a<>�a<��a<W�a< �a<��a<8�a<a<��a<�a<��a<Y�a< �a<֎a<M�a<�a<��a<t�a<8�a<֌a<��a<N�a<)�a<̋a<��a<w�a<6�a<�a<ߊa<Ҋa<��a<u�a<L�a<?�a<<�a<��a<��a<Ӊa<��a<ωa<��a<��a<��a<ȉa<��a<׉a<Չa<�a<��a<�a<@�a<�  �  Q�a<s�a<��a<��a<֊a<�a<J�a<s�a<��a<�a<�a<X�a<��a<Ռa<#�a<f�a<��a<	�a<L�a<��a<�a<e�a<ŏa<�a<p�a<�a<[�a<��a<�a<{�a<�a<R�a<��a<5�a<��a<�a<��a<	�a<y�a<��a<x�a<�a<j�a<��a<l�a<ؙa<U�a<ߚa<]�a<śa<K�a<��a<.�a<��a<!�a<��a<�a<~�a<�a<\�a<ˠa<B�a<��a<�a<��a<עa<4�a<��a<�a<L�a<��a<��a<Q�a<��a<�a<>�a<x�a<��a<�a<B�a<��a<˧a<�a<>�a<q�a<��a<�a< �a<8�a<n�a<��a<��a<ةa<�a<�a</�a<P�a<m�a<~�a<��a<��a<��a<ڪa<�a<��a<�a<�a<�a<�a<2�a<.�a<*�a<%�a<#�a< �a<�a<�a<�a< �a<��a<�a<̪a<Ȫa<��a<��a<��a<{�a<r�a<C�a<�a<�a<��a<ϩa<��a<��a<S�a<:�a<�a<ߨa<��a<��a<W�a</�a<�a<Χa<��a<c�a</�a<�a<��a<v�a<L�a<�a<��a<j�a<!�a<פa<��a<C�a<�a<��a<Z�a<�a<��a<Y�a<�a<��a<H�a<��a<��a<$�a<a<l�a<�a<��a<0�a<��a<J�a<�a<s�a<��a<��a<#�a<��a<=�a<˙a<b�a<�a<��a<�a<��a<�a<��a<I�a<Õa<Q�a<�a<y�a<�a<��a<5�a<��a<U�a<��a<��a<+�a<͐a<n�a<�a<��a<r�a<	�a<��a<]�a<�a<ƍa<n�a<,�a<Ԍa<��a<V�a<�a<�a<��a<v�a<I�a<	�a<�a<a<��a<��a<W�a</�a<�a<�a<��a<�a<Ӊa<ȉa<a<��a<a<ĉa<ŉa<҉a<މa<��a< �a<�a</�a<�  �  R�a<`�a<��a<��a<��a<#�a<0�a<��a<��a<�a<�a<\�a<��a<׌a<#�a<e�a<͍a<�a<`�a<��a<��a<l�a<��a<:�a<��a<ېa<@�a<��a<�a<m�a<��a<J�a<˓a<6�a<��a<�a<}�a<�a<o�a<	�a<k�a<�a<l�a<ܘa<o�a<͙a<��a<ߚa<O�a<՛a<C�a<Ӝa<+�a<��a<�a<��a<�a<y�a<�a<Y�a<�a<A�a<��a<�a<x�a<�a<+�a<��a<�a<M�a<��a<�a<_�a<��a<�a<*�a<|�a<��a<
�a<U�a<y�a<ܧa<��a<D�a<k�a<��a<ݨa<�a<]�a<W�a<��a<��a<�a<�a<�a<M�a<M�a<p�a<��a<��a<��a<ªa<�a<۪a<�a<��a<!�a<5�a<�a<1�a<�a<(�a<�a<&�a<*�a<�a<�a<�a<�a<֪a<�a<Ӫa<ͪa<��a<��a<��a<i�a<e�a<7�a<>�a< �a<ߩa<۩a<��a<��a<]�a<=�a<�a<�a<��a<��a<r�a<-�a<�a<ҧa<��a<j�a<�a<�a<��a<p�a<1�a<�a<��a<\�a<4�a<Ϥa<��a<D�a<�a<��a<@�a<�a<��a<e�a<��a<��a<J�a<�a<��a<�a<�a<l�a<��a<��a<)�a<ӝa<G�a<��a<q�a<�a<��a<�a<ɚa<:�a<�a<b�a<��a<z�a<�a<��a<�a<��a</�a<ŕa<\�a<ڔa<��a<�a<��a<"�a<��a<Q�a<��a<��a<�a<ސa<^�a<�a<��a<V�a<�a<��a<��a<�a<ča<o�a<4�a<�a<��a<t�a<�a<�a<��a<|�a<Q�a<�a<��a<��a<��a<n�a<i�a<W�a<�a<�a<�a<�a<ˉa<ˉa<͉a<��a<��a<��a<ˉa<��a<ډa<�a<�a<�a<&�a<�  �  E�a<y�a<��a<Ȋa<�a<��a<=�a<y�a<��a<݋a<$�a<T�a<��a<ތa<�a<j�a<��a<�a<d�a<��a<�a<j�a<��a<�a<��a<�a<?�a<��a<�a<u�a<ޒa<J�a<Óa<6�a<��a<�a<��a<�a<�a<��a<l�a<��a<k�a<�a<n�a<�a<O�a<Ěa<P�a<˛a<A�a<a<6�a<��a<"�a<��a<�a<��a<�a<a�a<Ԡa<7�a<��a<�a<e�a<͢a<J�a<��a<��a<V�a<��a<�a<I�a<��a<�a<3�a<x�a<��a<�a<L�a<��a<ŧa<��a<>�a<��a<��a<�a<�a<(�a<X�a<��a<��a<өa<��a<�a<.�a<O�a<e�a<��a<��a<��a<Ѫa<ުa<�a<��a<�a<��a<�a<+�a<+�a<*�a<�a<.�a<�a<�a<�a<�a<�a<��a<�a<�a<Ѫa<��a<��a<��a<��a<��a<c�a<T�a</�a<��a<�a<թa<��a<��a<k�a<5�a<�a<�a<��a<��a<T�a<-�a<�a<ŧa<��a<h�a<�a<צa<��a<��a<0�a<��a<��a<c�a<�a<Фa<��a<D�a<�a<��a<R�a<�a<��a<Q�a<��a<��a<J�a<�a<��a<:�a<��a<Q�a<��a<��a<&�a<Ýa<R�a<�a<t�a<�a<��a<%�a<��a<A�a<ԙa<X�a<�a<y�a<��a<��a<-�a<��a<>�a<Εa<_�a<ݔa<q�a<�a<��a<+�a<��a<V�a<�a<��a<$�a<ǐa<f�a<�a<Ïa<]�a<�a<��a<N�a<�a<ča<u�a<'�a<�a<��a<U�a<�a<ۋa<��a<m�a<A�a<�a<�a<��a<��a<y�a<B�a<8�a<,�a<�a<��a<ىa<܉a<a<��a<��a<a<��a<a<ȉa<��a<�a<��a<�a<4�a<�  �  <�a<}�a<z�a<��a<��a<�a<a�a<e�a<��a<׋a<�a<a�a<��a<�a<+�a<y�a<��a<�a<S�a<��a<�a<U�a<ޏa<�a<�a<ِa<5�a<��a<��a<��a<̒a<T�a<��a<(�a<��a<�a<��a<�a<z�a<�a<u�a<�a<e�a<��a<C�a<�a<R�a<��a<d�a<˛a<P�a<��a<D�a<��a<*�a<��a<�a<��a<�a<r�a<àa<E�a<��a<�a<��a<Ңa<I�a<~�a<��a<L�a<��a<�a<6�a<��a<ӥa<3�a<p�a<��a<��a<6�a<��a<��a<�a</�a<z�a<��a<Ϩa<�a<5�a<��a<��a<éa<թa<�a<+�a<,�a<]�a<w�a<��a<��a<��a<ɪa<Ҫa<��a<�a<%�a<$�a<�a<)�a<�a<7�a<�a</�a<�a<�a<�a<�a<�a<�a<�a<تa<Ǫa<êa<��a<��a<{�a<��a<G�a<L�a<'�a<�a<�a<��a<��a<�a<]�a<C�a<
�a<�a<¨a<��a<R�a<?�a<��a<ŧa<��a<S�a<H�a<�a<��a<n�a<'�a<��a<��a<x�a<�a<٤a<y�a<7�a<�a<��a<S�a<�a<��a<D�a<��a<��a<C�a<��a<l�a<:�a<��a<��a<�a<��a<5�a<��a<`�a<�a<|�a<�a<��a<*�a<��a<R�a<Ùa<f�a<�a<��a<'�a<��a<-�a<��a<@�a<ĕa<M�a<�a<^�a<�a<��a<+�a<��a<T�a<�a<z�a</�a<��a<{�a< �a<��a<W�a<��a<��a<[�a<1�a<��a<��a<(�a<ٌa<��a<S�a<)�a<�a<��a<t�a<N�a<�a<�a<Њa<��a<��a<k�a<3�a<*�a<�a<�a<Չa<݉a<��a<��a<��a<��a<��a<��a<͉a<͉a<ۉa<��a<�a<=�a<�  �  M�a<{�a<��a<Êa<�a<�a<(�a<s�a<��a<�a<�a<\�a<��a<͌a<+�a<[�a<ƍa<�a<^�a<��a<�a<V�a<��a<!�a<~�a<�a<K�a<��a<�a<z�a<�a<S�a<��a<3�a<��a<�a<��a<�a<~�a<��a<t�a<�a<s�a<�a<i�a<�a<`�a<Ԛa<>�a<؛a<D�a<̜a<1�a<��a<"�a<��a<�a<v�a<��a<]�a<ߠa<A�a<��a<��a<q�a<�a<@�a<��a<��a<[�a<��a<�a<I�a<��a<�a<,�a<~�a<��a<�a<E�a<��a<��a<�a<=�a<��a<��a<�a<�a<>�a<W�a<{�a<��a<�a<�a<�a<D�a<B�a<y�a<}�a<��a<��a<��a<�a<�a<��a<�a<�a<�a<+�a<)�a<4�a<&�a<"�a<�a<�a<�a<�a<��a<��a<�a<ުa<Ϫa<Ǫa<��a<��a<��a<��a<f�a<P�a<*�a<�a<שa<ϩa<��a<��a<Z�a<>�a<�a<רa<¨a<{�a<k�a<,�a< �a<٧a<��a<T�a<�a<�a<��a<��a<<�a<��a<��a<i�a<�a<٤a<��a<A�a<�a<��a<H�a<��a<��a<V�a<��a<��a<Q�a<��a<��a<2�a<Οa<a�a<�a<��a<)�a<͝a<M�a<�a<t�a<�a<��a<�a<��a<=�a<ޙa<a�a<��a<g�a< �a<��a<$�a<��a<B�a<ӕa<V�a<�a<q�a<�a<��a<$�a<a<T�a<�a<��a<-�a<a<o�a<�a<��a<f�a<�a<��a<c�a<�a<��a<}�a<6�a<�a<��a<k�a<�a<�a<��a<~�a<R�a<�a<��a<��a<��a<b�a<]�a<9�a<+�a<�a<�a<�a<Љa<a<��a<��a<��a<��a<ĉa<��a<Ӊa<�a<��a<�a<-�a<�  �  J�a<[�a<��a<��a<݊a<$�a<=�a<��a<��a<�a<�a<T�a<��a<Ҍa<>�a<Z�a<�a<��a<e�a<��a<��a<��a<Ïa<%�a<e�a<ސa<7�a<��a<�a<^�a<�a<F�a<��a<*�a<��a<+�a<n�a<�a<s�a<��a<f�a<�a<d�a<Ƙa<y�a<Йa<f�a<ݚa<a�a<��a<%�a<ۜa<#�a<ĝa<"�a<��a<%�a<}�a<�a<N�a<�a<�a<ġa<+�a<}�a<�a<*�a<��a<٣a<I�a<��a<�a<M�a<��a<�a<�a<��a<��a<��a<C�a<��a<ϧa<�a<7�a<m�a<��a<�a<��a<E�a<i�a<��a<��a<˩a<�a<��a<_�a<B�a<��a<��a<��a<��a<��a<�a<Ūa<:�a<�a< �a<�a<�a<2�a<�a<�a< �a<'�a<�a<�a<�a<�a<�a<ܪa<�a<Ȫa<��a<��a<��a<��a<d�a<f�a<>�a<$�a<!�a<�a<�a<��a<��a<_�a<6�a<*�a<ܨa<֨a<z�a<��a<�a<�a<ʧa<��a<��a<,�a<��a<��a<s�a<(�a<�a<��a<M�a<-�a<̤a<}�a<8�a<�a<��a<1�a< �a<��a<W�a<�a<��a<C�a<ˠa<��a<�a<ӟa<j�a<�a<��a<
�a<ܝa<?�a<��a<t�a<�a<��a<"�a<Ӛa<.�a<�a<@�a<�a<��a<�a<��a<�a<��a<�a<��a<M�a<Ӕa<u�a<��a<��a<�a<ɒa<M�a<�a<��a< �a<ѐa<Q�a<	�a<��a<H�a<�a<��a<j�a<�a<�a<r�a<�a<��a<��a<��a<�a<�a<��a<��a<K�a<�a< �a<��a<܊a<z�a<g�a<6�a<�a<�a<ډa<ډa<Ήa<̉a<��a<��a<��a<��a<߉a<��a<׉a<܉a<��a<�a<�a<�  �  M�a<{�a<��a<Êa<�a<�a<(�a<s�a<��a<�a<�a<\�a<��a<͌a<+�a<[�a<ƍa<�a<^�a<��a<�a<V�a<��a<!�a<~�a<�a<K�a<��a<�a<z�a<�a<S�a<��a<3�a<��a<�a<��a<�a<~�a<��a<t�a<�a<s�a<�a<i�a<�a<`�a<Ԛa<>�a<؛a<D�a<̜a<1�a<��a<"�a<��a<�a<v�a<��a<]�a<ߠa<A�a<��a<��a<q�a<�a<@�a<��a<��a<[�a<��a<�a<I�a<��a<�a<,�a<~�a<��a<�a<E�a<��a<��a<�a<=�a<��a<��a<�a<�a<>�a<W�a<{�a<��a<�a<�a<�a<D�a<B�a<y�a<}�a<��a<��a<��a<�a<�a<��a<�a<�a<�a<+�a<)�a<4�a<&�a<"�a<�a<�a<�a<�a<��a<��a<�a<ުa<Ϫa<Ǫa<��a<��a<��a<��a<f�a<P�a<*�a<�a<שa<ϩa<��a<��a<Z�a<>�a<�a<רa<¨a<{�a<k�a<,�a< �a<٧a<��a<T�a<�a<�a<��a<��a<<�a<��a<��a<i�a<�a<٤a<��a<A�a<�a<��a<H�a<��a<��a<V�a<��a<��a<Q�a<��a<��a<2�a<Οa<a�a<�a<��a<)�a<͝a<M�a<�a<t�a<�a<��a<�a<��a<=�a<ޙa<a�a<��a<g�a< �a<��a<$�a<��a<B�a<ӕa<V�a<�a<q�a<�a<��a<$�a<a<T�a<�a<��a<-�a<a<o�a<�a<��a<f�a<�a<��a<c�a<�a<��a<}�a<6�a<�a<��a<k�a<�a<�a<��a<~�a<R�a<�a<��a<��a<��a<b�a<]�a<9�a<+�a<�a<�a<�a<Љa<a<��a<��a<��a<��a<ĉa<��a<Ӊa<�a<��a<�a<-�a<�  �  <�a<}�a<z�a<��a<��a<�a<a�a<e�a<��a<׋a<�a<a�a<��a<�a<+�a<y�a<��a<�a<S�a<��a<�a<U�a<ޏa<�a<�a<ِa<5�a<��a<��a<��a<̒a<T�a<��a<(�a<��a<�a<��a<�a<z�a<�a<u�a<�a<e�a<��a<C�a<�a<R�a<��a<d�a<˛a<P�a<��a<D�a<��a<*�a<��a<�a<��a<�a<r�a<àa<E�a<��a<�a<��a<Ңa<I�a<~�a<��a<L�a<��a<�a<6�a<��a<ӥa<3�a<p�a<��a<��a<6�a<��a<��a<�a</�a<z�a<��a<Ϩa<�a<5�a<��a<��a<éa<թa<�a<+�a<,�a<]�a<w�a<��a<��a<��a<ɪa<Ҫa<��a<�a<%�a<$�a<�a<)�a<�a<7�a<�a</�a<�a<�a<�a<�a<�a<�a<�a<تa<Ǫa<êa<��a<��a<{�a<��a<G�a<L�a<'�a<�a<�a<��a<��a<�a<]�a<C�a<
�a<�a<¨a<��a<R�a<?�a<��a<ŧa<��a<S�a<H�a<�a<��a<n�a<'�a<��a<��a<x�a<�a<٤a<y�a<7�a<�a<��a<S�a<�a<��a<D�a<��a<��a<C�a<��a<l�a<:�a<��a<��a<�a<��a<5�a<��a<`�a<�a<|�a<�a<��a<*�a<��a<R�a<Ùa<f�a<�a<��a<'�a<��a<-�a<��a<@�a<ĕa<M�a<�a<^�a<�a<��a<+�a<��a<T�a<�a<z�a</�a<��a<{�a< �a<��a<W�a<��a<��a<[�a<1�a<��a<��a<(�a<ٌa<��a<S�a<)�a<�a<��a<t�a<N�a<�a<�a<Њa<��a<��a<k�a<3�a<*�a<�a<�a<Չa<݉a<��a<��a<��a<��a<��a<��a<͉a<͉a<ۉa<��a<�a<=�a<�  �  E�a<y�a<��a<Ȋa<�a<��a<=�a<y�a<��a<݋a<$�a<T�a<��a<ތa<�a<j�a<��a<�a<d�a<��a<�a<j�a<��a<�a<��a<�a<?�a<��a<�a<u�a<ޒa<J�a<Óa<6�a<��a<�a<��a<�a<�a<��a<l�a<��a<k�a<�a<n�a<�a<O�a<Ěa<P�a<˛a<A�a<a<6�a<��a<"�a<��a<�a<��a<�a<a�a<Ԡa<7�a<��a<�a<e�a<͢a<J�a<��a<��a<V�a<��a<�a<I�a<��a<�a<3�a<x�a<��a<�a<L�a<��a<ŧa<��a<>�a<��a<��a<�a<�a<(�a<X�a<��a<��a<өa<��a<�a<.�a<O�a<e�a<��a<��a<��a<Ѫa<ުa<�a<��a<�a<��a<�a<+�a<+�a<*�a<�a<.�a<�a<�a<�a<�a<�a<��a<�a<�a<Ѫa<��a<��a<��a<��a<��a<c�a<T�a</�a<��a<�a<թa<��a<��a<k�a<5�a<�a<�a<��a<��a<T�a<-�a<�a<ŧa<��a<h�a<�a<צa<��a<��a<0�a<��a<��a<c�a<�a<Фa<��a<D�a<�a<��a<R�a<�a<��a<Q�a<��a<��a<J�a<�a<��a<:�a<��a<Q�a<��a<��a<&�a<Ýa<R�a<�a<t�a<�a<��a<%�a<��a<A�a<ԙa<X�a<�a<y�a<��a<��a<-�a<��a<>�a<Εa<_�a<ݔa<q�a<�a<��a<+�a<��a<V�a<�a<��a<$�a<ǐa<f�a<�a<Ïa<]�a<�a<��a<N�a<�a<ča<u�a<'�a<�a<��a<U�a<�a<ۋa<��a<m�a<A�a<�a<�a<��a<��a<y�a<B�a<8�a<,�a<�a<��a<ىa<܉a<a<��a<��a<a<��a<a<ȉa<��a<�a<��a<�a<4�a<�  �  R�a<`�a<��a<��a<��a<#�a<0�a<��a<��a<�a<�a<\�a<��a<׌a<#�a<e�a<͍a<�a<`�a<��a<��a<l�a<��a<:�a<��a<ېa<@�a<��a<�a<m�a<��a<J�a<˓a<6�a<��a<�a<}�a<�a<o�a<	�a<k�a<�a<l�a<ܘa<o�a<͙a<��a<ߚa<O�a<՛a<C�a<Ӝa<+�a<��a<�a<��a<�a<y�a<�a<Y�a<�a<A�a<��a<�a<x�a<�a<+�a<��a<�a<M�a<��a<�a<_�a<��a<�a<*�a<|�a<��a<
�a<U�a<y�a<ܧa<��a<D�a<k�a<��a<ݨa<�a<]�a<W�a<��a<��a<�a<�a<�a<M�a<M�a<p�a<��a<��a<��a<ªa<�a<۪a<�a<��a<!�a<5�a<�a<1�a<�a<(�a<�a<&�a<*�a<�a<�a<�a<�a<֪a<�a<Ӫa<ͪa<��a<��a<��a<i�a<e�a<7�a<>�a< �a<ߩa<۩a<��a<��a<]�a<=�a<�a<�a<��a<��a<r�a<-�a<�a<ҧa<��a<j�a<�a<�a<��a<p�a<1�a<�a<��a<\�a<4�a<Ϥa<��a<D�a<�a<��a<@�a<�a<��a<e�a<��a<��a<J�a<�a<��a<�a<�a<l�a<��a<��a<)�a<ӝa<G�a<��a<q�a<�a<��a<�a<ɚa<:�a<�a<b�a<��a<z�a<�a<��a<�a<��a</�a<ŕa<\�a<ڔa<��a<�a<��a<"�a<��a<Q�a<��a<��a<�a<ސa<^�a<�a<��a<V�a<�a<��a<��a<�a<ča<o�a<4�a<�a<��a<t�a<�a<�a<��a<|�a<Q�a<�a<��a<��a<��a<n�a<i�a<W�a<�a<�a<�a<�a<ˉa<ˉa<͉a<��a<��a<��a<ˉa<��a<ډa<�a<�a<�a<&�a<�  �  Q�a<s�a<��a<��a<֊a<�a<J�a<s�a<��a<�a<�a<X�a<��a<Ռa<#�a<f�a<��a<	�a<L�a<��a<�a<e�a<ŏa<�a<p�a<�a<[�a<��a<�a<{�a<�a<R�a<��a<5�a<��a<�a<��a<	�a<y�a<��a<x�a<�a<j�a<��a<l�a<ؙa<U�a<ߚa<]�a<śa<K�a<��a<.�a<��a<!�a<��a<�a<~�a<�a<\�a<ˠa<B�a<��a<�a<��a<עa<4�a<��a<�a<L�a<��a<��a<Q�a<��a<�a<>�a<x�a<��a<�a<B�a<��a<˧a<�a<>�a<q�a<��a<�a< �a<8�a<n�a<��a<��a<ةa<�a<�a</�a<P�a<m�a<~�a<��a<��a<��a<ڪa<�a<��a<�a<�a<�a<�a<2�a<.�a<*�a<%�a<#�a< �a<�a<�a<�a< �a<��a<�a<̪a<Ȫa<��a<��a<��a<{�a<r�a<C�a<�a<�a<��a<ϩa<��a<��a<S�a<:�a<�a<ߨa<��a<��a<W�a</�a<�a<Χa<��a<c�a</�a<�a<��a<v�a<L�a<�a<��a<j�a<!�a<פa<��a<C�a<�a<��a<Z�a<�a<��a<Y�a<�a<��a<H�a<��a<��a<$�a<a<l�a<�a<��a<0�a<��a<J�a<�a<s�a<��a<��a<#�a<��a<=�a<˙a<b�a<�a<��a<�a<��a<�a<��a<I�a<Õa<Q�a<�a<y�a<�a<��a<5�a<��a<U�a<��a<��a<+�a<͐a<n�a<�a<��a<r�a<	�a<��a<]�a<�a<ƍa<n�a<,�a<Ԍa<��a<V�a<�a<�a<��a<v�a<I�a<	�a<�a<a<��a<��a<W�a</�a<�a<�a<��a<�a<Ӊa<ȉa<a<��a<a<ĉa<ŉa<҉a<މa<��a< �a<�a</�a<�  �  A�a<t�a<��a<ˊa<��a<�a<@�a<`�a<��a<׋a<�a<K�a<��a<݌a<�a<p�a<��a<	�a<O�a<��a<�a<N�a<��a<�a<��a<��a<9�a<��a<�a<��a<ޒa<Z�a<��a<=�a<��a<	�a<��a<��a<��a<�a<��a<�a<b�a<�a<S�a<�a<S�a<Ԛa<O�a<��a<W�a<��a<=�a<��a<-�a<��a<��a<��a<ߟa<j�a<��a<N�a<��a<�a<u�a<͢a<g�a<��a<��a<L�a<��a<�a<C�a<��a<ݥa<F�a<r�a<��a<�a<?�a<��a<��a<�a<4�a<u�a<��a<֨a<1�a<'�a<c�a<|�a<��a<�a<�a<�a<'�a<]�a<U�a<��a<��a<��a<Ȫa<Ъa<��a<�a<�a<�a<�a<;�a<�a<+�a<�a<2�a<)�a<�a<�a<
�a<�a<�a<��a<�a<Ӫa<Ūa<��a<��a<��a<|�a<T�a<X�a<7�a<�a<�a<��a<��a<�a<Z�a<,�a<�a<�a<��a<��a<P�a<.�a<�a<ϧa<��a<L�a<(�a<ݦa<Цa<u�a<+�a<�a<��a<~�a<�a<ߤa<��a<K�a<��a<��a<d�a<��a<��a<L�a<�a<��a<@�a<�a<}�a<U�a<��a<b�a<��a<��a<<�a<��a<Y�a<Ӝa<�a<��a<��a<0�a<��a<J�a<��a<o�a<��a<s�a<�a<��a<K�a<��a<:�a<Õa<Q�a<��a<k�a<�a<��a<>�a<��a<W�a< �a<��a<8�a<a<��a<�a<��a<Y�a< �a<֎a<M�a<�a<��a<t�a<8�a<֌a<��a<N�a<)�a<̋a<��a<w�a<6�a<�a<ߊa<Ҋa<��a<u�a<L�a<?�a<<�a<��a<��a<Ӊa<��a<ωa<��a<��a<��a<ȉa<��a<׉a<Չa<�a<��a<�a<@�a<�  �  T�a<{�a<��a<��a<��a<"�a<>�a<q�a<��a<׋a<�a<E�a<��a<ٌa<�a<k�a<��a<��a<X�a<��a<�a<`�a<ŏa<(�a<v�a<Ԑa<D�a<��a<�a<��a<�a<K�a<˓a<7�a<��a<�a<��a<�a<��a<�a<z�a<�a<v�a<��a<c�a<ՙa<a�a<�a<J�a<Ǜa<B�a<��a<0�a<��a<&�a<��a<�a<��a<�a<[�a<Рa<<�a<��a<	�a<��a<�a<3�a<��a<�a<^�a<��a<�a<I�a<��a<�a<8�a<~�a<��a<�a<S�a<��a<̧a<�a<=�a<��a<��a<Ԩa<�a<B�a<p�a<��a<��a<ԩa<��a<
�a<3�a<T�a<c�a<��a<��a<��a<Īa<ժa<�a<��a<�a<'�a<�a<�a<'�a<1�a</�a<+�a<,�a<�a< �a<�a<	�a<�a<�a<�a<ުa<��a<��a<��a<��a<��a<b�a<8�a<'�a<�a<�a<ͩa<��a<~�a<[�a<'�a<�a<�a<��a<��a<]�a<�a<��a<ħa<��a<]�a</�a<��a<��a<i�a<5�a<�a<��a<o�a<$�a<Ѥa<��a<E�a<�a<��a<V�a<��a<��a<L�a<�a<��a<T�a<��a<��a<!�a<Οa<v�a<��a<��a<(�a<��a<L�a<ڜa<x�a<��a<��a<)�a<��a<<�a<ϙa<]�a<�a<q�a<�a<��a<�a<��a<G�a<Օa<R�a<�a<q�a<�a<��a<0�a<Òa<V�a<��a<��a<'�a<ΐa<u�a<�a<Ïa<c�a<��a<��a<g�a<�a<��a<l�a<'�a<�a<��a<Z�a<!�a<ًa<��a<r�a<2�a<�a<�a<��a<��a<u�a<n�a<;�a<�a<�a<��a<�a<ىa<щa<��a<ĉa<��a<��a<ˉa<Ήa<܉a<�a<��a<�a<7�a<�  �  `�a<`�a<��a<ʊa<֊a<�a<.�a<r�a<��a<�a<�a<P�a<��a<��a<!�a<L�a<��a<��a<c�a<��a<��a<^�a<��a<(�a<f�a<��a<T�a<��a<�a<p�a<��a<N�a<֓a<;�a<��a<"�a<��a<$�a<��a<�a<��a<�a<r�a<�a<��a<יa<^�a<͚a<F�a<Λa<2�a<͜a<�a<��a<�a<��a<�a<s�a<��a<I�a<ߠa<-�a<��a<	�a<k�a<ߢa<-�a<ģa<��a<U�a<��a<�a<d�a<��a<�a<3�a<��a<ʦa<�a<a�a<��a<�a<�a<K�a<t�a<��a< �a<��a<C�a<U�a<��a<��a<ɩa<�a<�a<4�a<8�a<h�a<n�a<��a<��a<��a<�a<٪a<��a<��a<�a<�a<(�a<@�a<�a<7�a<�a</�a<'�a<�a<+�a<	�a<�a<��a<��a<�a<˪a<ªa<��a<��a<i�a<w�a<V�a<�a<�a<ݩa<Ωa<��a<��a<^�a<1�a<	�a<Ĩa<��a<m�a<[�a<�a<�a<§a<��a<\�a<�a<��a<��a<��a<E�a<�a<��a<_�a<3�a<Ԥa<��a<I�a<��a<��a<S�a<�a<��a<i�a<�a<��a<P�a<�a<��a<$�a<˟a<[�a<�a<��a<�a<Νa<9�a<�a<o�a<��a<��a<�a<��a<*�a<ޙa<M�a<�a<r�a<��a<��a<�a<֖a<:�a<̕a<_�a<�a<��a<�a<��a<*�a<Ȓa<_�a<��a<��a<%�a<�a<j�a<�a<��a<i�a<*�a<��a<i�a< �a<��a<p�a<�a<�a<��a<\�a<�a<ދa<��a<s�a<E�a<�a<��a<��a<��a<j�a<T�a<3�a<)�a<%�a<�a<�a<̉a<Չa<ʉa<a<Չa<��a<̉a<ωa<�a<�a<�a<"�a<&�a<�  �  \�a<m�a<{�a<��a<�a<�a<F�a<d�a<��a<Ћa<�a<L�a<��a<Ќa<�a<b�a<��a<��a<P�a<��a<�a<V�a<��a<!�a<��a<ؐa<-�a<��a<�a<y�a<�a<_�a<ēa<0�a<��a<�a<��a<�a<��a<�a<u�a<��a<r�a<ݘa<V�a<�a<g�a<ؚa<\�a<̛a<;�a<��a<*�a<��a<�a<��a<�a<w�a<�a<[�a<Ƞa<2�a<��a<�a<y�a<�a<J�a<��a<�a<T�a<��a<��a<U�a<��a<�a<9�a<��a<Цa<
�a<N�a<��a<ӧa<�a<B�a<x�a<��a<Ҩa<�a<@�a<b�a<��a<��a<ɩa<�a<�a<7�a<L�a<d�a<~�a<��a<��a<��a<ͪa<�a<�a<�a<�a<(�a<(�a<�a<#�a<5�a<'�a<$�a<0�a<�a<�a<�a<��a<��a<�a<۪a<٪a<��a<��a<��a<v�a<H�a<M�a<9�a<�a<��a<��a<��a<w�a<S�a<.�a<�a<٨a<��a<��a<_�a<$�a<�a<��a<��a<T�a<%�a<�a<��a<m�a<�a<��a<��a<h�a<+�a<�a<��a<?�a< �a<��a<U�a<��a<��a<`�a<��a<��a<P�a<�a<��a<8�a<ԟa<e�a<�a<��a< �a<��a<F�a<�a<l�a<��a<��a<�a<��a<;�a<Ǚa<S�a<�a<~�a<	�a<��a<.�a<��a<,�a<̕a<Z�a<�a<|�a<
�a<��a<1�a<˒a<f�a<��a<��a<3�a<Րa<k�a<�a<��a<I�a<��a<��a<e�a<�a<��a<}�a<�a<ڌa<��a<^�a<�a<ۋa<��a<t�a<>�a<	�a<܊a<��a<��a<��a<S�a<I�a<)�a<�a<�a<��a<Չa<ʉa<҉a<a<��a<Éa<��a<։a<؉a<�a<�a<�a<0�a<�  �  G�a<��a<��a<��a<�a<��a<H�a<Z�a<��a<ċa<�a<A�a<��a<ӌa<�a<d�a<��a<��a<K�a<��a<
�a<R�a<ˏa<��a<��a<Րa<Z�a<Ǒa<�a<��a<�a<\�a<Гa<8�a<��a<)�a<��a<�a<��a<�a<y�a<�a<i�a<�a<_�a<�a<I�a<Ԛa<R�a<��a<O�a<��a<4�a<��a<�a<��a<��a<w�a<֟a<_�a<��a<B�a<��a<�a<y�a<��a<H�a<��a<�a<X�a<��a<�a<E�a<��a<�a<@�a<��a<Цa<�a<V�a<��a<ça<�a<<�a<��a<ƨa<Өa<�a<�a<o�a<��a<��a<ϩa<�a<�a<�a<L�a<P�a<~�a<��a<��a<êa<��a<��a<�a<�a< �a<�a<"�a<)�a<K�a<�a<?�a<!�a<�a<.�a<�a<�a<�a<�a<�a<�a<ɪa<��a<��a<��a<��a<j�a<E�a<-�a<��a<��a<��a<��a<l�a<X�a<#�a<��a<ݨa<��a<��a<F�a<�a<�a<��a<��a<P�a<4�a<˦a<��a<j�a<K�a<�a<��a<z�a<�a<�a<��a<F�a<�a<��a<`�a<��a<Ģa<O�a<�a<��a<G�a<�a<��a<3�a<��a<a�a<��a<��a<4�a<��a<Q�a<ʜa<h�a<��a<��a<�a<��a<?�a<��a<c�a<ޘa<t�a<�a<x�a<,�a<��a<^�a<Еa<c�a<�a<l�a<�a<��a<8�a<Вa<f�a<��a<��a<<�a<Őa<|�a<�a<͏a<y�a<��a<��a<;�a<�a<��a<p�a<#�a<Ќa<��a<D�a<�a<ǋa<��a<g�a<,�a<�a<͊a<͊a<��a<�a<G�a<8�a<#�a<�a<�a<ډa<�a<ǉa<��a<҉a<��a<щa<҉a<މa<ډa<��a<�a<�a<I�a<�  �  R�a<[�a<��a<��a<�a<�a<G�a<l�a<��a<Ջa<�a<H�a<��a<ǌa<�a<X�a<��a<��a<U�a<��a< �a<_�a<ɏa<�a<��a<ސa<J�a<��a<�a<{�a<��a<Q�a<֓a<>�a<��a<,�a<��a<�a<��a<�a<��a<��a<\�a<ޘa<i�a<�a<h�a<ߚa<\�a<ța<D�a<��a<3�a<��a<�a<��a<�a<t�a<�a<^�a<Ơa<>�a<��a<�a<~�a<�a<?�a<��a<�a<A�a<��a<�a<a�a<��a<��a<.�a<��a<ʦa<�a<_�a<��a<ܧa<�a<L�a<c�a<��a<ߨa<�a<=�a<k�a<��a<��a<ϩa<��a<�a</�a<A�a<h�a<u�a<��a<��a<Īa<Ҫa<�a<��a<�a<�a<%�a<#�a<,�a<�a<#�a<0�a<7�a<%�a<�a<$�a<��a<�a<�a<��a<ߪa<Ȫa<ɪa<��a<��a<d�a<h�a<G�a<5�a<�a<��a<ǩa<��a<}�a<Z�a<*�a<�a<Ѩa<��a<y�a<S�a<$�a<��a<��a<��a<\�a<2�a<�a<��a<s�a<;�a<ޥa<��a<i�a<6�a<פa<��a<L�a<�a<��a<I�a<�a<��a<g�a<�a<��a<:�a<�a<��a<.�a<֟a<m�a<�a<��a<)�a<��a<O�a<ڜa<l�a<��a<��a<�a<��a<>�a<ƙa<_�a<�a<��a<�a<��a<#�a<��a<5�a<��a<i�a<�a<��a<�a<��a<&�a<ђa<_�a<��a<��a<,�a<ݐa<n�a<�a<��a<_�a<	�a<��a<b�a<�a<��a<o�a<"�a<ߌa<��a<V�a<�a<ދa<��a<q�a<6�a<�a<�a<��a<��a<�a<_�a<G�a<#�a<�a<�a<މa<މa<܉a<ǉa<a<Ήa<��a<҉a<ĉa<�a<�a< �a<*�a<6�a<�  �  /�a<H�a<��a<��a<ɋa<�a<�a<P�a<i�a<��a<�a<�a<i�a<��a<�a<%�a<��a<Ɏa<6�a<}�a<͏a<<�a<��a<��a<O�a<��a<%�a<k�a<��a<3�a<Ǔa<�a<��a<
�a<|�a<��a<Z�a<�a<4�a<×a<0�a<��a<%�a<��a<$�a<��a<+�a<��a<
�a<��a<�a<z�a<ܝa<N�a<Ğa<*�a<��a<�a<��a<��a<��a<Ρa<I�a<��a<�a<��a<̣a<<�a<��a<�a<A�a<��a<��a<+�a<��a<ئa<7�a<s�a<��a<��a<�a<��a<��a<ܨa<�a<Z�a<r�a<��a<�a<��a<8�a<F�a<i�a<��a<��a<Ϫa<۪a<��a<	�a<7�a<D�a<n�a<��a<t�a<��a<��a<��a<̫a<��a<֫a<ͫa<̫a<��a<ӫa<«a<��a<ɫa<��a<ȫa<��a<��a<y�a<h�a<k�a<6�a<8�a<�a<�a<٪a<۪a<��a<��a<w�a<9�a<1�a<�a<̩a<��a<k�a<H�a<�a<��a<��a<��a<h�a<-�a<�a<��a<��a<Y�a<�a<�a<��a<U�a<��a<ݥa<q�a<9�a<��a<��a<h�a<��a<£a<C�a<�a<��a<A�a<�a<��a<;�a< a<��a<�a<��a<C�a<��a<w�a<��a<��a<�a<��a<0�a<ʛa<^�a<�a<��a<�a<��a<;�a<��a<h�a<̗a<l�a<�a<��a<�a<��a<J�a<��a<x�a<��a<��a<4�a<˒a<h�a<�a<��a<-�a<ސa<~�a<>�a<͏a<~�a<B�a<Վa<��a<<�a<�a<ƍa<d�a<,�a<݌a<��a<e�a<F�a<�a<�a<ʋa<��a<�a<L�a<6�a<%�a<�a<�a<ӊa<��a<��a<��a<��a<��a<��a<��a<Ɗa<��a<Ǌa<Ċa<؊a<�a<��a<�  �  /�a<F�a<v�a<��a<��a<ߋa<�a<G�a<��a<��a<��a<)�a<n�a<��a<��a<@�a<��a<ӎa<�a<s�a<ۏa<.�a<��a<ސa<Q�a<��a<�a<q�a<�a<Q�a<Ɠa<&�a<��a<�a<d�a<ϕa<V�a<Ֆa<I�a<ȗa<@�a<Øa<&�a<��a<&�a<��a<�a<�a<��a<z�a<��a<Z�a<ڝa<T�a<Ӟa<A�a<��a<+�a<��a< �a<`�a<�a<H�a<��a<�a<z�a<�a<A�a<��a<�a<Y�a<��a<��a<A�a<��a<ئa<�a<X�a<��a<�a<3�a<}�a<��a<�a<�a<Q�a<z�a<��a<Ωa<��a<&�a<R�a<j�a<��a<��a<תa<�a<�a<%�a<@�a<O�a<\�a<c�a<��a<��a<��a<��a<��a<ʫa<ѫa<ɫa<Ϋa<۫a<׫a<ѫa<ƫa<��a<��a<��a<��a<��a<��a<z�a<k�a<V�a<9�a<�a<�a<�a<Ъa<��a<��a<o�a<W�a<�a<�a<ةa<��a<��a<]�a</�a<�a<ɨa<��a<^�a<;�a<��a<ʧa<��a<[�a<�a<�a<��a<`�a<�a<ۥa<��a<6�a<�a<��a<8�a<��a<��a<X�a<	�a<��a<`�a<�a<��a<=�a<ܠa<m�a< �a<��a<:�a<ڞa<W�a<��a<��a<'�a<��a<C�a<ڛa<b�a<�a<p�a<�a<��a<,�a<��a<L�a<�a<q�a< �a<��a<*�a<��a<H�a<єa<j�a<��a<}�a<�a<ǒa<]�a<�a<��a<F�a<�a<��a<5�a<֏a<��a<&�a<܎a<��a<G�a<�a<��a<j�a<3�a<�a<��a<��a<O�a<�a<�a<��a<��a<q�a<K�a<*�a<�a<�a<�a<Ίa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ϊa<�a<�a<�a<�  �  $�a<X�a<j�a<��a<��a<�a<(�a<.�a<��a<��a<��a<*�a<Y�a<��a<�a<5�a<}�a<ގa<0�a<��a<܏a<�a<��a<�a<X�a<��a<�a<~�a<ߒa<L�a<��a<-�a<��a<	�a<��a<�a<w�a<Ȗa<T�a<��a<(�a<��a<)�a<��a<�a<��a<�a<��a<�a<i�a<�a<a�a<�a<N�a<��a<2�a<��a<�a<��a<�a<j�a<�a<>�a<��a<.�a<r�a<�a<2�a<��a<�a<J�a<��a<�a<O�a<��a<�a<)�a<x�a<��a<�a<<�a<e�a<��a<�a<�a<K�a<w�a<��a<ͩa<�a<�a<O�a<|�a<��a<��a<Ȫa<�a<��a<�a<+�a<P�a<w�a<o�a<��a<��a<��a<��a<��a<ɫa<īa<ثa<ʫa<իa<��a<ͫa<̫a<��a<Ыa<��a<��a<��a<��a<x�a<M�a<P�a<.�a<+�a<�a<�a<˪a<��a<��a<U�a<_�a<�a<�a<٩a<��a<~�a<J�a<$�a<�a<Өa<��a<o�a<<�a<�a<�a<��a<b�a<�a<֦a<��a<U�a<�a<��a<��a<0�a<��a<��a<R�a<�a<��a<d�a<�a<��a<P�a<�a<��a<-�a<�a<d�a<�a<��a<*�a<�a<^�a<�a<��a<�a<��a<2�a<ʛa<Y�a<�a<y�a<$�a<��a<)�a<՘a<D�a<�a<b�a<�a<��a<�a<��a<>�a<ߔa<_�a<�a<��a<9�a<ђa<S�a<�a<��a<>�a<�a<��a</�a<ҏa<��a<%�a<��a<}�a<E�a<�a<��a<{�a<%�a<�a<��a<x�a<:�a<�a<��a<��a<��a<Y�a<_�a<;�a<	�a<�a<��a<ފa<��a<��a<��a<��a<��a<��a<��a<��a<ʊa<��a<Њa<�a<�a<�a<�  �  /�a<W�a<n�a<��a<a<�a<�a<J�a<s�a<��a<�a<�a<r�a<��a<��a<:�a<��a<Ǝa<3�a<t�a<ԏa<3�a<��a<��a<O�a<��a<�a<~�a<�a<J�a<��a<�a<��a<��a<m�a<��a<P�a<ٖa<?�a<ɗa<;�a<��a<6�a<��a<�a<��a<�a<��a<��a<��a<�a<p�a<ڝa<T�a<Ξa<E�a<��a<'�a<��a<��a<x�a<ѡa<N�a<��a<�a<��a<٣a<7�a<��a<��a<P�a<��a<��a<8�a<��a<Φa<�a<c�a<��a<��a<&�a<w�a<��a<�a<�a<K�a<{�a<��a<ߩa<��a<)�a<M�a<e�a<��a<��a<تa<�a<�a<$�a<?�a<D�a<c�a<|�a<�a<��a<��a<��a<ëa<��a<ȫa<ԫa<ӫa<ϫa<իa<ƫa<ëa<��a<��a<��a<��a<��a<��a<k�a<i�a<N�a<8�a<)�a<�a<�a<Ԫa<��a<��a<q�a<C�a<%�a<�a<ǩa<��a<��a<d�a<)�a<�a<��a<��a<_�a<3�a<�a<��a<��a<X�a<�a<զa<��a<]�a<�a<ӥa<y�a<A�a<�a<��a<I�a<�a<��a<N�a<
�a<��a<Q�a<��a<��a<0�a<Рa<z�a<�a<��a<A�a<a<m�a<��a<��a<"�a<��a<I�a<՛a<b�a<�a<��a<�a<��a<)�a<��a<V�a<ٗa<g�a< �a<��a<"�a<��a<K�a<Ȕa<o�a<�a<��a<$�a<��a<j�a<��a<��a<>�a<�a<��a</�a<׏a<��a<8�a<Ԏa<��a<C�a<�a<��a<_�a<5�a<�a<a<�a<N�a<�a<�a<Ëa<��a<w�a<K�a</�a<�a<��a<�a<ڊa<Ɗa<��a<��a<��a<��a<��a<��a<��a<��a<��a<Њa<ڊa<�a<�a<�  �  2�a<>�a<|�a<��a<��a<�a<�a<i�a<t�a<��a<�a<$�a<t�a<��a<�a<�a<��a<Ɏa<5�a<r�a<ڏa<L�a<x�a<��a<<�a<��a<�a<n�a<�a<=�a<̓a<�a<��a<��a<q�a<��a<H�a<�a<,�a<��a<8�a<��a<-�a<��a<0�a<��a<"�a<��a<��a<��a<�a<�a<ѝa<`�a<��a<5�a<��a<�a<��a<�a<��a<ˡa<^�a<��a<�a<��a<Σa<M�a<��a<�a<N�a<��a<��a<#�a<��a<ɦa<5�a<o�a<��a< �a<�a<��a<��a<�a<�a<E�a<��a<��a<�a<�a<<�a<X�a<c�a<��a<��a<�a<Ҫa<�a<�a<<�a<Q�a<V�a<�a<�a<��a<��a<��a<��a<īa<ثa<��a<ӫa<ƫa<߫a<��a<��a<ǫa<��a<ëa<��a<��a<{�a<c�a<v�a<B�a<;�a<�a<�a<�a<̪a<��a<��a<��a<D�a<%�a<��a<өa<��a<j�a<j�a<
�a<�a<��a<��a<]�a<:�a<�a<��a<��a<E�a<%�a<٦a<��a<]�a<�a<�a<j�a<B�a<�a<��a<f�a<�a<��a<;�a<�a<��a<O�a<��a<��a<H�a<Ǡa<��a< �a<��a<Y�a<a<{�a<�a<��a<�a<��a<?�a<��a<m�a<�a<��a<��a<��a<1�a<��a<a�a<Ηa<}�a<�a<��a< �a<��a<H�a<��a<y�a<�a<��a<0�a<��a<p�a<�a<��a</�a<�a<��a<)�a<�a<s�a<C�a<Ɏa<��a<N�a<�a<ƍa<^�a<?�a<Ԍa<Ìa<i�a<K�a<�a<ۋa<Ƌa<��a<��a<C�a<1�a<�a<��a<��a<��a<Ǌa<��a<��a<��a<��a<��a<��a<��a<��a<��a<Ɗa<ӊa<�a<�a<�  �  5�a<O�a<m�a<��a<��a<��a<#�a<4�a<|�a<��a<�a<'�a<g�a<��a<	�a<3�a<��a<Ԏa<,�a<��a<׏a<#�a<��a<�a<F�a<��a<�a<}�a<�a<C�a<��a<'�a<��a<��a<l�a<�a<S�a<Ɩa<Q�a<ȗa<)�a<��a</�a<��a<�a<��a<�a<��a<�a<s�a<��a<i�a<�a<U�a<a<K�a<a<�a<��a<�a<r�a<ޡa<D�a<��a<0�a<s�a<ޣa<=�a<��a<��a<J�a<��a<��a<K�a<��a<Ӧa<$�a<f�a<��a<�a<4�a<n�a<��a<�a<�a<H�a<��a<��a<֩a<�a<�a<L�a<s�a<��a<��a<תa<�a<!�a<&�a<4�a<R�a<n�a<x�a<��a<��a<��a<ūa<��a<ʫa<ȫa<ҫa<ثa<ƫa<��a<Ыa<īa<��a<��a<��a<��a<��a<��a<w�a<V�a<C�a<?�a<"�a<�a<��a<ªa<��a<��a<[�a<K�a<*�a<�a<֩a<��a<��a<o�a<#�a<�a<ʨa<��a<k�a<6�a<�a<اa<��a<P�a<#�a<֦a<��a<Z�a<
�a<ʥa<��a<2�a<�a<��a<Q�a<��a<��a<`�a<	�a<��a<L�a<��a<��a<6�a<Ԡa<d�a<#�a<��a<4�a<Ӟa<f�a<�a<��a<�a<��a<R�a<̛a<a�a<�a<��a<�a<��a<-�a<טa<F�a<ޗa<m�a<��a<��a<�a<��a<E�a<۔a<^�a<��a<��a<'�a<��a<Y�a<�a<��a<3�a<�a<��a<,�a<ݏa<��a</�a<��a<��a<B�a<��a<��a<l�a<4�a<�a<͌a<��a<C�a<�a<�a<��a<��a<`�a<Y�a<E�a<�a<�a<�a<؊a<ˊa<��a<��a<��a<��a<��a<��a<��a<��a<��a<̊a<�a<�a<�a<�  �  �a<]�a<[�a<��a<��a<ًa<(�a<<�a<��a<��a<�a<,�a<t�a<��a<�a<N�a<��a<�a<)�a<}�a<�a<'�a<��a<Аa<]�a<��a<�a<��a<Ԓa<_�a<��a<-�a<��a<�a<q�a<ԕa<d�a<��a<P�a<��a<=�a<��a<#�a<��a<�a<��a<��a<��a<	�a<z�a<�a<U�a<�a<K�a<۞a<B�a<��a<2�a<��a<�a<_�a<�a<R�a<��a<!�a<`�a<��a<�a<��a<�a<S�a<��a<ۥa<K�a<}�a<�a<�a<f�a<��a<�a<:�a<R�a<��a<بa<�a<K�a<f�a<éa<��a<�a<#�a<_�a<x�a<��a<ªa<˪a< �a<��a<)�a<G�a<O�a<s�a<g�a<��a<��a<��a<��a<��a<ѫa<��a<ޫa<��a<ݫa<īa<ūa<ūa<��a<��a<��a<��a<��a<��a<q�a<Q�a<^�a<(�a</�a<�a<�a<Ъa<��a<��a<d�a<c�a<�a<�a<۩a<��a<��a<H�a<=�a<��a<רa<��a<h�a<H�a<��a<ާa<v�a<f�a<
�a<Ӧa<��a<I�a<&�a<��a<��a<-�a<�a<��a<=�a<�a<��a<_�a<�a<��a<Z�a<�a<��a<�a<�a<W�a<�a<��a<;�a<�a<R�a<�a<��a</�a<��a<>�a<�a<W�a<�a<n�a<!�a<��a<1�a<Șa<2�a<��a<O�a<�a<��a<%�a<��a<(�a<۔a<T�a<�a<��a<'�a<Βa<P�a<	�a<��a<O�a<ڐa<��a</�a<��a<��a<�a<�a<��a<T�a< �a<��a<~�a<(�a<�a<��a<��a<V�a<�a<��a<��a<��a<h�a<_�a<*�a<�a<
�a<͊a<�a<��a<Êa<��a<��a<��a<��a<��a<��a<��a<��a<̊a<��a<�a<"�a<�  �  �a<X�a<z�a<��a<ɋa<�a<�a<R�a<w�a<��a<��a<-�a<j�a<��a<��a<=�a<��a<��a<8�a<x�a<ӏa<=�a<��a<�a<Q�a<��a<%�a<|�a<̒a<G�a<��a<'�a<��a<�a<q�a<��a<P�a<Ζa<=�a<��a<4�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<�a<r�a<�a<U�a<˞a<C�a<��a<%�a<��a<�a<}�a<ӡa<N�a<��a<�a<~�a<ߣa<5�a<��a<�a<A�a<��a<�a<9�a<��a<Φa<.�a<l�a<��a<�a<1�a<f�a<��a<Ҩa<�a<`�a<k�a<��a<کa<	�a<3�a<O�a<h�a<��a<ªa<ͪa<�a<�a<#�a<<�a<Q�a<p�a<{�a<��a<��a<��a<��a<ȫa<��a<ͫa<ثa<��a<˫a<ʫa<ƫa<��a<��a<��a<��a<��a<��a<y�a<q�a<_�a<H�a< �a<*�a<�a<�a<۪a<��a<��a<y�a<G�a<#�a<�a<ܩa<��a<��a<b�a<-�a<��a<ըa<��a<c�a<3�a<�a<ҧa<��a<[�a<�a<�a<��a<B�a<�a<ĥa<��a<3�a<ݤa<��a<_�a<�a<��a<L�a<��a<��a<G�a<�a<��a<3�a<֠a<t�a<
�a<��a<D�a<Ȟa<o�a<�a<��a< �a<��a<I�a<ӛa<c�a<�a<��a<�a<��a<5�a<��a<P�a<ޗa<e�a<�a<��a<�a<��a<8�a<ɔa<_�a<�a<��a<-�a<��a<Y�a< �a<��a<;�a<Ӑa<��a<D�a<Ǐa<��a<2�a<�a<��a<D�a<�a<a<~�a<*�a<��a<��a<~�a<K�a<�a<�a<a<��a<|�a<X�a<0�a<"�a<�a<�a<ފa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<Ŋa<��a<��a<�a<�  �  J�a<9�a<w�a<��a<ŋa<�a<�a<P�a<u�a<Όa<�a<,�a<p�a<��a<�a<0�a<��a<͎a<)�a<��a<ԏa<9�a<~�a<��a<I�a<��a<�a<j�a<��a<8�a<��a<�a<��a<��a<Y�a<�a<9�a<ٖa</�a<Ηa<!�a<��a<7�a<��a<1�a<��a<!�a<��a<�a<��a<�a<��a<̝a<n�a<ƞa<N�a<ǟa<�a<��a<�a<��a<סa<T�a<��a<�a<��a<ͣa<N�a<��a<��a<X�a<��a<�a<)�a<��a<��a<�a<U�a<��a<�a<�a<y�a<��a<��a<�a<?�a<��a<��a<�a<��a<0�a<P�a<}�a<��a<��a<�a<�a<)�a<%�a<;�a<\�a<V�a<��a<��a<��a<��a<��a<ȫa<��a<׫a<��a<�a<ʫa<��a<ɫa<��a<ūa<��a<��a<{�a<��a<t�a<h�a<V�a<B�a<S�a<�a<�a<�a<תa<��a<��a<w�a<D�a<B�a<��a<۩a<��a<��a<y�a< �a<�a<èa<��a<~�a<3�a<	�a<��a<��a<S�a<!�a<Ӧa<��a<s�a<��a<ϥa<m�a<4�a<�a<��a<P�a<ܣa<��a<>�a<�a<��a<W�a<��a<�a<H�a<àa<��a<�a<��a<K�a<ƞa<�a<�a<��a<�a<��a<W�a<ʛa<|�a<ښa<��a<	�a<��a<1�a<��a<_�a<̗a<~�a<�a<��a<*�a<��a<N�a<��a<j�a<ܓa<��a<�a<��a<a�a<�a<��a<+�a<��a<|�a<#�a<�a<x�a<B�a<юa<��a<F�a<�a<��a<_�a<I�a<�a<֌a<��a<K�a<#�a<ۋa<ۋa<��a<|�a<G�a<5�a<"�a<�a<�a<��a<݊a<��a<��a<��a<��a<��a<x�a<��a<��a<Ċa<��a<׊a<�a<�a<�  �  +�a<B�a<s�a<��a<��a<�a<#�a<M�a<��a<��a<�a<4�a<n�a<��a<��a<9�a<��a<܎a<0�a<��a<ۏa<:�a<��a<�a<G�a<��a<�a<p�a<�a<8�a<��a<�a<��a<��a<o�a<�a<V�a<͖a<1�a<ŗa<%�a<��a<%�a<��a<&�a<��a<�a<��a<�a<��a<��a<|�a<ݝa<f�a<Ǟa<>�a<��a<�a<��a< �a<��a<�a<S�a<��a<�a<y�a<ڣa<C�a<��a<�a<K�a<��a<��a</�a<��a<զa<#�a<g�a<��a<�a<#�a<m�a<��a<�a<�a<?�a<��a<��a<ԩa<�a<7�a<T�a<|�a<��a<��a<�a<�a<�a<$�a<<�a<`�a<c�a<��a<��a<��a<��a<��a<��a<ȫa<ϫa<��a<Ϋa<ƫa<��a<˫a<��a<��a<��a<��a<��a<��a<i�a<p�a<W�a<A�a<5�a<�a<
�a<�a<̪a<��a<��a<u�a<S�a<4�a<��a<�a<��a<��a<[�a<(�a<
�a<Ѩa<��a<w�a<;�a<
�a<ѧa<��a<Q�a<!�a<Ҧa<��a<W�a<��a<ɥa<x�a<'�a<�a<��a<R�a<��a<��a<@�a<�a<��a<L�a<�a<��a<=�a<Ѡa<p�a<�a<��a<F�a<֞a<y�a<��a<��a<�a<��a<?�a<͛a<r�a<�a<��a<�a<��a<:�a<Ƙa<K�a<ٗa<s�a<�a<��a<�a<��a<A�a<��a<_�a<��a<��a<(�a<��a<U�a<�a<��a<*�a<�a<�a<#�a<�a<�a<,�a<�a<��a<I�a<�a<��a<o�a<=�a<�a<��a<�a<L�a<'�a<�a<͋a<��a<{�a<Z�a<.�a<�a< �a<�a<Ŋa<a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ߊa<�a<�a<�  �  �a<\�a<k�a<��a<a<�a<$�a<C�a<��a<��a<��a<0�a<q�a<ˍa<��a<`�a<��a<�a<3�a<q�a<��a<2�a<��a<�a<S�a<��a<�a<��a<Òa<\�a<��a</�a<��a<�a<d�a<ϕa<J�a<��a<O�a<��a<@�a<��a<�a<��a<�a<��a<�a<��a<�a<�a<��a<i�a<��a<P�a<�a<R�a<��a<B�a<��a<�a<u�a<ݡa<L�a<��a<"�a<s�a<�a<2�a<��a<�a<?�a<��a<�a<M�a<~�a<ʦa<�a<X�a<��a<�a<<�a<]�a<��a<Ȩa<�a<W�a<n�a<��a<ѩa<�a<,�a<V�a<e�a<��a<Ǫa<Ъa<�a<�a<>�a<H�a<R�a<v�a<s�a<��a<��a<��a<��a<��a<ͫa<��a<�a<��a<ԫa<ȫa<̫a<«a<��a<��a<��a<��a<z�a<�a<z�a<T�a<Y�a<�a</�a<�a<�a<Ԫa<��a<��a<j�a<S�a<�a<�a<ߩa<��a<��a<_�a<O�a<��a<ިa<��a<\�a<@�a<�a<קa<��a<\�a<�a<�a<��a<9�a<#�a<��a<��a<1�a<֤a<��a<8�a<�a<��a<^�a<��a<��a<I�a<ޡa<��a<*�a<�a<j�a<�a<��a<?�a<Ԟa<f�a<�a<��a<5�a<Ĝa<Q�a<�a<b�a<�a<��a<�a<��a<.�a<ɘa<E�a<�a<b�a<�a<~�a<�a<��a<2�a<ޔa<U�a<�a<z�a<�a<��a<T�a<�a<��a<N�a<ʐa<��a<;�a<ʏa<��a<*�a<�a<��a<L�a<�a<��a<��a<-�a<�a<��a<��a<W�a<�a<��a<��a<��a<s�a<Z�a<-�a<�a<�a<܊a<�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ʊa<�a<�a<�a<�  �  +�a<H�a<c�a<��a<��a<�a<�a<P�a<��a<Ōa<��a<0�a<s�a<��a<�a<@�a<��a<�a<7�a<��a<�a<2�a<��a<��a<R�a<��a<	�a<p�a<ܒa<P�a<��a<�a<��a<�a<o�a<�a<W�a<͖a<;�a<��a<.�a<��a<%�a<��a<�a<��a<�a<��a<�a<��a<��a<}�a<�a<Z�a<Ԟa<5�a<��a<)�a<��a<
�a<��a<�a<Z�a<��a< �a<��a<�a<9�a<��a<�a<F�a<��a<إa<7�a<��a<٦a<�a<f�a<��a<�a<#�a<V�a<��a<ڨa<�a<=�a<x�a<��a<�a<�a<*�a<d�a<��a<��a<��a<ܪa<�a<��a<�a<E�a<U�a<p�a<��a<��a<��a<��a<��a<��a<ǫa<��a<˫a<ʫa<Ыa<��a<��a<��a<��a<��a<��a<��a<��a<{�a<^�a<G�a<Q�a<4�a<�a<��a<�a<Ҫa<��a<��a<w�a<Z�a<9�a<�a<ީa<��a<��a<K�a</�a<�a<רa<��a<y�a<G�a<�a<ȧa<��a<\�a<�a<Цa<��a<Q�a<�a<��a<u�a<0�a<�a<��a<L�a<��a<��a<K�a<�a<��a<K�a<�a<��a<.�a<ܠa<r�a<�a<��a<L�a<ݞa<z�a<�a<��a<(�a<��a<6�a<؛a<k�a<��a<��a<�a<��a<,�a<ǘa<R�a<�a<i�a<�a<��a<�a<��a<&�a<ǔa<_�a<��a<��a<'�a<Œa<X�a<�a<��a<D�a<ܐa<}�a<!�a<ԏa<��a<9�a<��a<��a<Y�a<�a<a<z�a<9�a<�a<��a<x�a<T�a<�a<��a<Ջa<��a<�a<K�a<<�a<�a< �a<׊a<ъa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<Ǌa<͊a<ފa<�a<�  �  2�a<A�a<|�a<��a<��a<��a<�a<N�a<k�a<Ča<�a<)�a<y�a<��a<�a<F�a<��a<юa<*�a<��a<ďa</�a<��a<��a<;�a<��a<�a<u�a<�a</�a<��a<#�a<~�a<��a<S�a<ҕa<F�a<ǖa<5�a<̗a<(�a<��a<7�a<��a<3�a<��a<�a<��a<��a<x�a<�a<��a<ӝa<g�a<מa<R�a<˟a<*�a<��a<��a<��a<աa<D�a<��a<#�a<{�a<ͣa<T�a<��a<��a<C�a<��a<��a<2�a<��a<ʦa<
�a<L�a<��a<ߧa<(�a<x�a<��a<�a<�a<D�a<��a<��a<�a<�a<'�a<B�a<s�a<��a<��a<�a<��a<-�a<0�a<J�a<U�a<[�a<��a<x�a<��a<��a<ɫa<��a<ȫa<׫a<«a<իa<��a<ʫa<ͫa<��a<��a<��a<��a<~�a<��a<n�a<s�a<f�a<8�a<;�a<�a<�a<��a<��a<Īa<��a<u�a<;�a<9�a<��a<ةa<��a<��a<}�a<6�a<�a<ƨa<��a<s�a<$�a<��a<̧a<��a<D�a<+�a<ئa<��a<`�a<��a<ѥa<��a<$�a<�a<�a<:�a<�a<��a<D�a<�a<��a<B�a<��a<��a<J�a<ʠa<j�a<�a<��a<9�a<ƞa<�a<�a<��a<+�a<Üa<Z�a<؛a<w�a<�a<��a<�a<��a<*�a<ʘa<M�a<͗a<��a<�a<��a<�a<��a<J�a<a<Z�a<�a<y�a<�a<��a<O�a<��a<��a<(�a<�a<��a<(�a<�a<q�a<9�a<�a<��a<8�a<��a<��a<e�a<L�a<��a<ٌa<��a<Y�a<�a<��a<Ջa<��a<w�a<E�a<H�a<�a<�a<�a<Ǌa<Ɋa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<�a<��a<��a<�  �  +�a<H�a<c�a<��a<��a<�a<�a<P�a<��a<Ōa<��a<0�a<s�a<��a<�a<@�a<��a<�a<7�a<��a<�a<2�a<��a<��a<R�a<��a<	�a<p�a<ܒa<P�a<��a<�a<��a<�a<o�a<�a<W�a<͖a<;�a<��a<.�a<��a<%�a<��a<�a<��a<�a<��a<�a<��a<��a<}�a<�a<Z�a<Ԟa<5�a<��a<)�a<��a<
�a<��a<�a<Z�a<��a< �a<��a<�a<9�a<��a<�a<F�a<��a<إa<7�a<��a<٦a<�a<f�a<��a<�a<#�a<V�a<��a<ڨa<�a<=�a<x�a<��a<�a<�a<*�a<d�a<��a<��a<��a<ܪa<�a<��a<�a<E�a<U�a<p�a<��a<��a<��a<��a<��a<��a<ǫa<��a<˫a<ʫa<Ыa<��a<��a<��a<��a<��a<��a<��a<��a<{�a<^�a<G�a<Q�a<4�a<�a<��a<�a<Ҫa<��a<��a<w�a<Z�a<9�a<�a<ީa<��a<��a<K�a</�a<�a<רa<��a<y�a<G�a<�a<ȧa<��a<\�a<�a<Цa<��a<Q�a<�a<��a<u�a<0�a<�a<��a<L�a<��a<��a<K�a<�a<��a<K�a<�a<��a<.�a<ܠa<r�a<�a<��a<L�a<ݞa<z�a<�a<��a<(�a<��a<6�a<؛a<k�a<��a<��a<�a<��a<,�a<ǘa<R�a<�a<i�a<�a<��a<�a<��a<&�a<ǔa<_�a<��a<��a<'�a<Œa<X�a<�a<��a<D�a<ܐa<}�a<!�a<ԏa<��a<9�a<��a<��a<Y�a<�a<a<z�a<9�a<�a<��a<x�a<T�a<�a<��a<Ջa<��a<�a<K�a<<�a<�a< �a<׊a<ъa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<Ǌa<͊a<ފa<�a<�  �  �a<\�a<k�a<��a<a<�a<$�a<C�a<��a<��a<��a<0�a<q�a<ˍa<��a<`�a<��a<�a<3�a<q�a<��a<2�a<��a<�a<S�a<��a<�a<��a<Òa<\�a<��a</�a<��a<�a<d�a<ϕa<J�a<��a<O�a<��a<@�a<��a<�a<��a<�a<��a<�a<��a<�a<�a<��a<i�a<��a<P�a<�a<R�a<��a<B�a<��a<�a<u�a<ݡa<L�a<��a<"�a<s�a<�a<2�a<��a<�a<?�a<��a<�a<M�a<~�a<ʦa<�a<X�a<��a<�a<<�a<]�a<��a<Ȩa<�a<W�a<n�a<��a<ѩa<�a<,�a<V�a<e�a<��a<Ǫa<Ъa<�a<�a<>�a<H�a<R�a<v�a<s�a<��a<��a<��a<��a<��a<ͫa<��a<�a<��a<ԫa<ȫa<̫a<«a<��a<��a<��a<��a<z�a<�a<z�a<T�a<Y�a<�a</�a<�a<�a<Ԫa<��a<��a<j�a<S�a<�a<�a<ߩa<��a<��a<_�a<O�a<��a<ިa<��a<\�a<@�a<�a<קa<��a<\�a<�a<�a<��a<9�a<#�a<��a<��a<1�a<֤a<��a<8�a<�a<��a<^�a<��a<��a<I�a<ޡa<��a<*�a<�a<j�a<�a<��a<?�a<Ԟa<f�a<�a<��a<5�a<Ĝa<Q�a<�a<b�a<�a<��a<�a<��a<.�a<ɘa<E�a<�a<b�a<�a<~�a<�a<��a<2�a<ޔa<U�a<�a<z�a<�a<��a<T�a<�a<��a<N�a<ʐa<��a<;�a<ʏa<��a<*�a<�a<��a<L�a<�a<��a<��a<-�a<�a<��a<��a<W�a<�a<��a<��a<��a<s�a<Z�a<-�a<�a<�a<܊a<�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ʊa<�a<�a<�a<�  �  +�a<B�a<s�a<��a<��a<�a<#�a<M�a<��a<��a<�a<4�a<n�a<��a<��a<9�a<��a<܎a<0�a<��a<ۏa<:�a<��a<�a<G�a<��a<�a<p�a<�a<8�a<��a<�a<��a<��a<o�a<�a<V�a<͖a<1�a<ŗa<%�a<��a<%�a<��a<&�a<��a<�a<��a<�a<��a<��a<|�a<ݝa<f�a<Ǟa<>�a<��a<�a<��a< �a<��a<�a<S�a<��a<�a<y�a<ڣa<C�a<��a<�a<K�a<��a<��a</�a<��a<զa<#�a<g�a<��a<�a<#�a<m�a<��a<�a<�a<?�a<��a<��a<ԩa<�a<7�a<T�a<|�a<��a<��a<�a<�a<�a<$�a<<�a<`�a<c�a<��a<��a<��a<��a<��a<��a<ȫa<ϫa<��a<Ϋa<ƫa<��a<˫a<��a<��a<��a<��a<��a<��a<i�a<p�a<W�a<A�a<5�a<�a<
�a<�a<̪a<��a<��a<u�a<S�a<4�a<��a<�a<��a<��a<[�a<(�a<
�a<Ѩa<��a<w�a<;�a<
�a<ѧa<��a<Q�a<!�a<Ҧa<��a<W�a<��a<ɥa<x�a<'�a<�a<��a<R�a<��a<��a<@�a<�a<��a<L�a<�a<��a<=�a<Ѡa<p�a<�a<��a<F�a<֞a<y�a<��a<��a<�a<��a<?�a<͛a<r�a<�a<��a<�a<��a<:�a<Ƙa<K�a<ٗa<s�a<�a<��a<�a<��a<A�a<��a<_�a<��a<��a<(�a<��a<U�a<�a<��a<*�a<�a<�a<#�a<�a<�a<,�a<�a<��a<I�a<�a<��a<o�a<=�a<�a<��a<�a<L�a<'�a<�a<͋a<��a<{�a<Z�a<.�a<�a< �a<�a<Ŋa<a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ߊa<�a<�a<�  �  J�a<9�a<w�a<��a<ŋa<�a<�a<P�a<u�a<Όa<�a<,�a<p�a<��a<�a<0�a<��a<͎a<)�a<��a<ԏa<9�a<~�a<��a<I�a<��a<�a<j�a<��a<8�a<��a<�a<��a<��a<Y�a<�a<9�a<ٖa</�a<Ηa<!�a<��a<7�a<��a<1�a<��a<!�a<��a<�a<��a<�a<��a<̝a<n�a<ƞa<N�a<ǟa<�a<��a<�a<��a<סa<T�a<��a<�a<��a<ͣa<N�a<��a<��a<X�a<��a<�a<)�a<��a<��a<�a<U�a<��a<�a<�a<y�a<��a<��a<�a<?�a<��a<��a<�a<��a<0�a<P�a<}�a<��a<��a<�a<�a<)�a<%�a<;�a<\�a<V�a<��a<��a<��a<��a<��a<ȫa<��a<׫a<��a<�a<ʫa<��a<ɫa<��a<ūa<��a<��a<{�a<��a<t�a<h�a<V�a<B�a<S�a<�a<�a<�a<תa<��a<��a<w�a<D�a<B�a<��a<۩a<��a<��a<y�a< �a<�a<èa<��a<~�a<3�a<	�a<��a<��a<S�a<!�a<Ӧa<��a<s�a<��a<ϥa<m�a<4�a<�a<��a<P�a<ܣa<��a<>�a<�a<��a<W�a<��a<�a<H�a<àa<��a<�a<��a<K�a<ƞa<�a<�a<��a<�a<��a<W�a<ʛa<|�a<ښa<��a<	�a<��a<1�a<��a<_�a<̗a<~�a<�a<��a<*�a<��a<N�a<��a<j�a<ܓa<��a<�a<��a<a�a<�a<��a<+�a<��a<|�a<#�a<�a<x�a<B�a<юa<��a<F�a<�a<��a<_�a<I�a<�a<֌a<��a<K�a<#�a<ۋa<ۋa<��a<|�a<G�a<5�a<"�a<�a<�a<��a<݊a<��a<��a<��a<��a<��a<x�a<��a<��a<Ċa<��a<׊a<�a<�a<�  �  �a<X�a<z�a<��a<ɋa<�a<�a<R�a<w�a<��a<��a<-�a<j�a<��a<��a<=�a<��a<��a<8�a<x�a<ӏa<=�a<��a<�a<Q�a<��a<%�a<|�a<̒a<G�a<��a<'�a<��a<�a<q�a<��a<P�a<Ζa<=�a<��a<4�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<�a<r�a<�a<U�a<˞a<C�a<��a<%�a<��a<�a<}�a<ӡa<N�a<��a<�a<~�a<ߣa<5�a<��a<�a<A�a<��a<�a<9�a<��a<Φa<.�a<l�a<��a<�a<1�a<f�a<��a<Ҩa<�a<`�a<k�a<��a<کa<	�a<3�a<O�a<h�a<��a<ªa<ͪa<�a<�a<#�a<<�a<Q�a<p�a<{�a<��a<��a<��a<��a<ȫa<��a<ͫa<ثa<��a<˫a<ʫa<ƫa<��a<��a<��a<��a<��a<��a<y�a<q�a<_�a<H�a< �a<*�a<�a<�a<۪a<��a<��a<y�a<G�a<#�a<�a<ܩa<��a<��a<b�a<-�a<��a<ըa<��a<c�a<3�a<�a<ҧa<��a<[�a<�a<�a<��a<B�a<�a<ĥa<��a<3�a<ݤa<��a<_�a<�a<��a<L�a<��a<��a<G�a<�a<��a<3�a<֠a<t�a<
�a<��a<D�a<Ȟa<o�a<�a<��a< �a<��a<I�a<ӛa<c�a<�a<��a<�a<��a<5�a<��a<P�a<ޗa<e�a<�a<��a<�a<��a<8�a<ɔa<_�a<�a<��a<-�a<��a<Y�a< �a<��a<;�a<Ӑa<��a<D�a<Ǐa<��a<2�a<�a<��a<D�a<�a<a<~�a<*�a<��a<��a<~�a<K�a<�a<�a<a<��a<|�a<X�a<0�a<"�a<�a<�a<ފa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<Ŋa<��a<��a<�a<�  �  �a<]�a<[�a<��a<��a<ًa<(�a<<�a<��a<��a<�a<,�a<t�a<��a<�a<N�a<��a<�a<)�a<}�a<�a<'�a<��a<Аa<]�a<��a<�a<��a<Ԓa<_�a<��a<-�a<��a<�a<q�a<ԕa<d�a<��a<P�a<��a<=�a<��a<#�a<��a<�a<��a<��a<��a<	�a<z�a<�a<U�a<�a<K�a<۞a<B�a<��a<2�a<��a<�a<_�a<�a<R�a<��a<!�a<`�a<��a<�a<��a<�a<S�a<��a<ۥa<K�a<}�a<�a<�a<f�a<��a<�a<:�a<R�a<��a<بa<�a<K�a<f�a<éa<��a<�a<#�a<_�a<x�a<��a<ªa<˪a< �a<��a<)�a<G�a<O�a<s�a<g�a<��a<��a<��a<��a<��a<ѫa<��a<ޫa<��a<ݫa<īa<ūa<ūa<��a<��a<��a<��a<��a<��a<q�a<Q�a<^�a<(�a</�a<�a<�a<Ъa<��a<��a<d�a<c�a<�a<�a<۩a<��a<��a<H�a<=�a<��a<רa<��a<h�a<H�a<��a<ާa<v�a<f�a<
�a<Ӧa<��a<I�a<&�a<��a<��a<-�a<�a<��a<=�a<�a<��a<_�a<�a<��a<Z�a<�a<��a<�a<�a<W�a<�a<��a<;�a<�a<R�a<�a<��a</�a<��a<>�a<�a<W�a<�a<n�a<!�a<��a<1�a<Șa<2�a<��a<O�a<�a<��a<%�a<��a<(�a<۔a<T�a<�a<��a<'�a<Βa<P�a<	�a<��a<O�a<ڐa<��a</�a<��a<��a<�a<�a<��a<T�a< �a<��a<~�a<(�a<�a<��a<��a<V�a<�a<��a<��a<��a<h�a<_�a<*�a<�a<
�a<͊a<�a<��a<Êa<��a<��a<��a<��a<��a<��a<��a<��a<̊a<��a<�a<"�a<�  �  5�a<O�a<m�a<��a<��a<��a<#�a<4�a<|�a<��a<�a<'�a<g�a<��a<	�a<3�a<��a<Ԏa<,�a<��a<׏a<#�a<��a<�a<F�a<��a<�a<}�a<�a<C�a<��a<'�a<��a<��a<l�a<�a<S�a<Ɩa<Q�a<ȗa<)�a<��a</�a<��a<�a<��a<�a<��a<�a<s�a<��a<i�a<�a<U�a<a<K�a<a<�a<��a<�a<r�a<ޡa<D�a<��a<0�a<s�a<ޣa<=�a<��a<��a<J�a<��a<��a<K�a<��a<Ӧa<$�a<f�a<��a<�a<4�a<n�a<��a<�a<�a<H�a<��a<��a<֩a<�a<�a<L�a<s�a<��a<��a<תa<�a<!�a<&�a<4�a<R�a<n�a<x�a<��a<��a<��a<ūa<��a<ʫa<ȫa<ҫa<ثa<ƫa<��a<Ыa<īa<��a<��a<��a<��a<��a<��a<w�a<V�a<C�a<?�a<"�a<�a<��a<ªa<��a<��a<[�a<K�a<*�a<�a<֩a<��a<��a<o�a<#�a<�a<ʨa<��a<k�a<6�a<�a<اa<��a<P�a<#�a<֦a<��a<Z�a<
�a<ʥa<��a<2�a<�a<��a<Q�a<��a<��a<`�a<	�a<��a<L�a<��a<��a<6�a<Ԡa<d�a<#�a<��a<4�a<Ӟa<f�a<�a<��a<�a<��a<R�a<̛a<a�a<�a<��a<�a<��a<-�a<טa<F�a<ޗa<m�a<��a<��a<�a<��a<E�a<۔a<^�a<��a<��a<'�a<��a<Y�a<�a<��a<3�a<�a<��a<,�a<ݏa<��a</�a<��a<��a<B�a<��a<��a<l�a<4�a<�a<͌a<��a<C�a<�a<�a<��a<��a<`�a<Y�a<E�a<�a<�a<�a<؊a<ˊa<��a<��a<��a<��a<��a<��a<��a<��a<��a<̊a<�a<�a<�a<�  �  2�a<>�a<|�a<��a<��a<�a<�a<i�a<t�a<��a<�a<$�a<t�a<��a<�a<�a<��a<Ɏa<5�a<r�a<ڏa<L�a<x�a<��a<<�a<��a<�a<n�a<�a<=�a<̓a<�a<��a<��a<q�a<��a<H�a<�a<,�a<��a<8�a<��a<-�a<��a<0�a<��a<"�a<��a<��a<��a<�a<�a<ѝa<`�a<��a<5�a<��a<�a<��a<�a<��a<ˡa<^�a<��a<�a<��a<Σa<M�a<��a<�a<N�a<��a<��a<#�a<��a<ɦa<5�a<o�a<��a< �a<�a<��a<��a<�a<�a<E�a<��a<��a<�a<�a<<�a<X�a<c�a<��a<��a<�a<Ҫa<�a<�a<<�a<Q�a<V�a<�a<�a<��a<��a<��a<��a<īa<ثa<��a<ӫa<ƫa<߫a<��a<��a<ǫa<��a<ëa<��a<��a<{�a<c�a<v�a<B�a<;�a<�a<�a<�a<̪a<��a<��a<��a<D�a<%�a<��a<өa<��a<j�a<j�a<
�a<�a<��a<��a<]�a<:�a<�a<��a<��a<E�a<%�a<٦a<��a<]�a<�a<�a<j�a<B�a<�a<��a<f�a<�a<��a<;�a<�a<��a<O�a<��a<��a<H�a<Ǡa<��a< �a<��a<Y�a<a<{�a<�a<��a<�a<��a<?�a<��a<m�a<�a<��a<��a<��a<1�a<��a<a�a<Ηa<}�a<�a<��a< �a<��a<H�a<��a<y�a<�a<��a<0�a<��a<p�a<�a<��a</�a<�a<��a<)�a<�a<s�a<C�a<Ɏa<��a<N�a<�a<ƍa<^�a<?�a<Ԍa<Ìa<i�a<K�a<�a<ۋa<Ƌa<��a<��a<C�a<1�a<�a<��a<��a<��a<Ǌa<��a<��a<��a<��a<��a<��a<��a<��a<��a<Ɗa<ӊa<�a<�a<�  �  /�a<W�a<n�a<��a<a<�a<�a<J�a<s�a<��a<�a<�a<r�a<��a<��a<:�a<��a<Ǝa<3�a<t�a<ԏa<3�a<��a<��a<O�a<��a<�a<~�a<�a<J�a<��a<�a<��a<��a<m�a<��a<P�a<ٖa<?�a<ɗa<;�a<��a<6�a<��a<�a<��a<�a<��a<��a<��a<�a<p�a<ڝa<T�a<Ξa<E�a<��a<'�a<��a<��a<x�a<ѡa<N�a<��a<�a<��a<٣a<7�a<��a<��a<P�a<��a<��a<8�a<��a<Φa<�a<c�a<��a<��a<&�a<w�a<��a<�a<�a<K�a<{�a<��a<ߩa<��a<)�a<M�a<e�a<��a<��a<تa<�a<�a<$�a<?�a<D�a<c�a<|�a<�a<��a<��a<��a<ëa<��a<ȫa<ԫa<ӫa<ϫa<իa<ƫa<ëa<��a<��a<��a<��a<��a<��a<k�a<i�a<N�a<8�a<)�a<�a<�a<Ԫa<��a<��a<q�a<C�a<%�a<�a<ǩa<��a<��a<d�a<)�a<�a<��a<��a<_�a<3�a<�a<��a<��a<X�a<�a<զa<��a<]�a<�a<ӥa<y�a<A�a<�a<��a<I�a<�a<��a<N�a<
�a<��a<Q�a<��a<��a<0�a<Рa<z�a<�a<��a<A�a<a<m�a<��a<��a<"�a<��a<I�a<՛a<b�a<�a<��a<�a<��a<)�a<��a<V�a<ٗa<g�a< �a<��a<"�a<��a<K�a<Ȕa<o�a<�a<��a<$�a<��a<j�a<��a<��a<>�a<�a<��a</�a<׏a<��a<8�a<Ԏa<��a<C�a<�a<��a<_�a<5�a<�a<a<�a<N�a<�a<�a<Ëa<��a<w�a<K�a</�a<�a<��a<�a<ڊa<Ɗa<��a<��a<��a<��a<��a<��a<��a<��a<��a<Њa<ڊa<�a<�a<�  �  $�a<X�a<j�a<��a<��a<�a<(�a<.�a<��a<��a<��a<*�a<Y�a<��a<�a<5�a<}�a<ގa<0�a<��a<܏a<�a<��a<�a<X�a<��a<�a<~�a<ߒa<L�a<��a<-�a<��a<	�a<��a<�a<w�a<Ȗa<T�a<��a<(�a<��a<)�a<��a<�a<��a<�a<��a<�a<i�a<�a<a�a<�a<N�a<��a<2�a<��a<�a<��a<�a<j�a<�a<>�a<��a<.�a<r�a<�a<2�a<��a<�a<J�a<��a<�a<O�a<��a<�a<)�a<x�a<��a<�a<<�a<e�a<��a<�a<�a<K�a<w�a<��a<ͩa<�a<�a<O�a<|�a<��a<��a<Ȫa<�a<��a<�a<+�a<P�a<w�a<o�a<��a<��a<��a<��a<��a<ɫa<īa<ثa<ʫa<իa<��a<ͫa<̫a<��a<Ыa<��a<��a<��a<��a<x�a<M�a<P�a<.�a<+�a<�a<�a<˪a<��a<��a<U�a<_�a<�a<�a<٩a<��a<~�a<J�a<$�a<�a<Өa<��a<o�a<<�a<�a<�a<��a<b�a<�a<֦a<��a<U�a<�a<��a<��a<0�a<��a<��a<R�a<�a<��a<d�a<�a<��a<P�a<�a<��a<-�a<�a<d�a<�a<��a<*�a<�a<^�a<�a<��a<�a<��a<2�a<ʛa<Y�a<�a<y�a<$�a<��a<)�a<՘a<D�a<�a<b�a<�a<��a<�a<��a<>�a<ߔa<_�a<�a<��a<9�a<ђa<S�a<�a<��a<>�a<�a<��a</�a<ҏa<��a<%�a<��a<}�a<E�a<�a<��a<{�a<%�a<�a<��a<x�a<:�a<�a<��a<��a<��a<Y�a<_�a<;�a<	�a<�a<��a<ފa<��a<��a<��a<��a<��a<��a<��a<��a<ʊa<��a<Њa<�a<�a<�a<�  �  /�a<F�a<v�a<��a<��a<ߋa<�a<G�a<��a<��a<��a<)�a<n�a<��a<��a<@�a<��a<ӎa<�a<s�a<ۏa<.�a<��a<ސa<Q�a<��a<�a<q�a<�a<Q�a<Ɠa<&�a<��a<�a<d�a<ϕa<V�a<Ֆa<I�a<ȗa<@�a<Øa<&�a<��a<&�a<��a<�a<�a<��a<z�a<��a<Z�a<ڝa<T�a<Ӟa<A�a<��a<+�a<��a< �a<`�a<�a<H�a<��a<�a<z�a<�a<A�a<��a<�a<Y�a<��a<��a<A�a<��a<ئa<�a<X�a<��a<�a<3�a<}�a<��a<�a<�a<Q�a<z�a<��a<Ωa<��a<&�a<R�a<j�a<��a<��a<תa<�a<�a<%�a<@�a<O�a<\�a<c�a<��a<��a<��a<��a<��a<ʫa<ѫa<ɫa<Ϋa<۫a<׫a<ѫa<ƫa<��a<��a<��a<��a<��a<��a<z�a<k�a<V�a<9�a<�a<�a<�a<Ъa<��a<��a<o�a<W�a<�a<�a<ةa<��a<��a<]�a</�a<�a<ɨa<��a<^�a<;�a<��a<ʧa<��a<[�a<�a<�a<��a<`�a<�a<ۥa<��a<6�a<�a<��a<8�a<��a<��a<X�a<	�a<��a<`�a<�a<��a<=�a<ܠa<m�a< �a<��a<:�a<ڞa<W�a<��a<��a<'�a<��a<C�a<ڛa<b�a<�a<p�a<�a<��a<,�a<��a<L�a<�a<q�a< �a<��a<*�a<��a<H�a<єa<j�a<��a<}�a<�a<ǒa<]�a<�a<��a<F�a<�a<��a<5�a<֏a<��a<&�a<܎a<��a<G�a<�a<��a<j�a<3�a<�a<��a<��a<O�a<�a<�a<��a<��a<q�a<K�a<*�a<�a<�a<�a<Ίa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ϊa<�a<�a<�a<�  �  ��a<�a<B�a<Q�a<��a<��a<�a<"�a<-�a<��a<Ǎa<�a<2�a<g�a<��a<��a<T�a<��a<�a<L�a<��a<�a<[�a<��a<�a<g�a<ؒa<*�a<��a<�a<q�a<֔a<_�a<��a<8�a<��a<�a<|�a<�a<s�a<�a<S�a<˙a<G�a<Κa<4�a<͛a<E�a<��a<'�a<��a</�a<~�a<��a<c�a<՟a<E�a<��a<3�a<��a<2�a<w�a<�a<^�a<��a<!�a<d�a<Ԥa<$�a<|�a<Υa<<�a<��a<֦a<%�a<^�a<ӧa<�a<3�a<��a<��a<��a<A�a<`�a<��a<�a<�a<:�a<v�a<��a<Ѫa<Ӫa<�a<N�a<;�a<m�a<}�a<��a<��a<ӫa<�a<�a<+�a<�a<>�a<K�a<U�a<c�a<M�a<h�a<Y�a<S�a<d�a<i�a<Y�a<n�a<F�a<J�a<b�a<;�a<�a<,�a<��a<��a<�a<��a<��a<��a<v�a<t�a<T�a<4�a<�a<ͪa<֪a<��a<g�a<I�a<�a<�a<��a<��a<W�a<T�a<�a<��a<��a<n�a<4�a<�a<��a<x�a<%�a<ڦa<��a<c�a<�a<�a<u�a<D�a<�a<��a<;�a<��a<��a<J�a<ۢa<�a<%�a<ԡa<a�a<�a<��a<T�a<��a<d�a<(�a<��a<1�a<��a<K�a<ۜa<n�a<�a<��a<P�a<��a<K�a<�a<|�a<�a<}�a<�a<��a<3�a<��a<j�a<��a<��a< �a<��a<h�a<��a<r�a<-�a<��a<X�a<�a<��a<;�a<�a<��a<@�a<��a<��a<h�a<��a<ʎa<��a<(�a<��a<��a<n�a<<�a<�a<ތa<��a<��a<O�a<K�a<(�a<�a<��a<��a<��a<��a<z�a<~�a<{�a<h�a<}�a<\�a<k�a<��a<��a<z�a<��a<��a<ŋa<ۋa<�  �  �a<+�a<7�a<e�a<��a<��a<֌a<�a<L�a<j�a<��a<�a<2�a<}�a<��a<�a<O�a<��a<ޏa<:�a<��a<�a<B�a<��a<�a<l�a<Ւa<H�a<��a<�a<a�a<�a<L�a<��a<,�a<��a<�a<z�a<�a<k�a<�a<k�a<�a<\�a<Śa<G�a<��a<"�a<��a<�a<��a<��a<t�a<�a<m�a<�a<V�a<Ġa<)�a<��a<��a<r�a<ߢa<:�a<��a<��a<w�a<Τa<6�a<��a<�a<5�a<z�a<�a<�a<s�a<��a<��a<A�a<��a<ͨa<�a<A�a<�a<��a<�a<�a<C�a<W�a<��a<��a<�a<�a<�a<@�a<e�a<��a<��a<��a<ҫa<�a<�a<��a<'�a<*�a<1�a<4�a<N�a<a�a<[�a<s�a<|�a<q�a<]�a<a�a<f�a<M�a<V�a<*�a<C�a<$�a<#�a<�a<�a<�a<�a<̫a<��a<��a<h�a<6�a<�a<�a<�a<��a<��a<k�a<I�a<'�a<��a<Ωa<��a<_�a<%�a<��a<ڨa<��a<V�a<�a<�a<��a<u�a<C�a<��a<��a<S�a<$�a<ҥa<��a<8�a<֤a<��a<9�a<��a<��a<C�a<�a<��a<:�a<ˡa<s�a<��a<��a<3�a<֟a<n�a<��a<��a<)�a<ĝa<\�a<�a<{�a<�a<��a<�a<��a<I�a<͙a<Y�a<�a<��a<�a<��a<T�a<ٖa<d�a<�a<��a<�a<��a<=�a<ޓa<��a<�a<ƒa<J�a<�a<��a<[�a<��a<��a<I�a<ߏa<��a<G�a<�a<��a<f�a<-�a<�a<a<��a<O�a<�a<یa<��a<v�a<h�a<6�a<�a<�a<ۋa<͋a<��a<��a<��a<��a<o�a<o�a<v�a<c�a<w�a<[�a<��a<��a<��a<��a<��a<�a<�  �  �a<�a<%�a<o�a<��a<��a<��a<��a<S�a<o�a<��a<��a<&�a<p�a<��a<��a<=�a<��a<�a<>�a<��a<ݐa<k�a<��a<�a<m�a<Òa<%�a<��a<	�a<^�a<�a<3�a<��a<=�a<��a<,�a<g�a<��a<l�a<�a<[�a<əa<G�a<��a<V�a<��a<N�a<��a<�a<��a<�a<��a<�a<i�a<ҟa<B�a<��a<"�a<��a<�a<~�a<ݢa<J�a<ˣa<�a<��a<��a<"�a<t�a<إa<3�a<y�a<ئa< �a<��a<��a<�a<J�a<j�a<Өa<�a<>�a<j�a<��a<ѩa<�a<H�a<e�a<��a<��a<�a<	�a<'�a<a�a<X�a<��a<��a<��a<ȫa<�a<
�a< �a</�a<�a<O�a<U�a<O�a<o�a<J�a<X�a<Z�a<d�a<_�a<j�a<Q�a<A�a<g�a<)�a<P�a<�a<�a<�a<�a<�a<īa<��a<��a<��a<g�a<Q�a<B�a<�a<�a<��a<��a<w�a<=�a<�a<�a<��a<��a<y�a<8�a<��a<ܨa<��a<�a<)�a<�a<��a<c�a< �a<�a<��a<P�a<.�a<��a<��a<I�a<ޤa<��a<&�a<�a<��a<D�a<�a<}�a<%�a<��a<��a<�a<àa<I�a<ҟa<}�a<��a<��a<&�a<��a<H�a<ٜa<v�a<��a<��a<!�a<a<G�a<ܙa<��a<�a<��a<	�a<��a<+�a<ɖa<b�a<�a<��a<��a<ʔa<I�a<�a<��a<�a<̒a<I�a<�a<��a<5�a<�a<��a<N�a<�a<��a<E�a<�a<a<x�a<N�a<�a<��a<s�a<A�a<
�a<�a<��a<y�a<p�a<+�a<-�a<�a<܋a<ۋa<��a<��a<��a<~�a<q�a<x�a<a�a<W�a<��a<Z�a<��a<x�a<��a<��a<��a<ߋa<�  �  �a<�a<T�a<Z�a<��a<��a<֌a<�a<8�a<�a<��a<ݍa<:�a<m�a<��a< �a<S�a<��a<�a<>�a<��a<��a<J�a<��a<��a<u�a<�a<:�a<��a<�a<t�a<ؔa<[�a<��a<�a<��a<�a<��a<��a<y�a<�a<]�a<ԙa<e�a<��a<9�a<��a<-�a<��a<!�a<��a<�a<t�a<�a<u�a<�a<V�a<ɠa<,�a<��a<�a<m�a<ܢa<E�a<��a<�a<j�a<�a<E�a<��a<ޥa<9�a<��a<֦a<2�a<a�a<��a<�a<:�a<��a<��a<�a<A�a<u�a<��a<��a<�a<3�a<c�a<��a<êa<تa< �a<.�a<0�a<j�a<��a<��a<��a<ܫa<ثa<��a<�a<�a<8�a<2�a<F�a<N�a<S�a<{�a<o�a<_�a<g�a<o�a<]�a<d�a<\�a<@�a<B�a<)�a</�a<(�a<�a<��a<�a<ɫa<��a<��a<�a<a�a<E�a<�a<�a<تa<Īa<��a<]�a<Q�a<�a<��a<éa<��a<N�a<:�a<��a<èa<��a<]�a<!�a<�a<��a<��a<5�a<�a<��a<f�a<�a<�a<��a<(�a<�a<��a<T�a<��a<��a<L�a<�a<��a<C�a<�a<f�a<�a<��a<8�a<ڟa<g�a<�a<��a<&�a<̝a<Z�a<�a<�a<�a<��a</�a<��a<F�a<יa<f�a<�a<��a</�a<ŗa<:�a<ϖa<g�a<��a<��a<-�a<��a<@�a<דa<y�a<-�a<��a<a�a<�a<��a<I�a<�a<��a<9�a<�a<��a<Z�a<��a<��a<~�a<�a<��a<��a<��a<C�a<�a<Ҍa<��a<��a<T�a<E�a<�a<��a<ۋa<��a<ˋa<��a<��a<��a<��a<k�a<s�a<r�a<a�a<s�a<o�a<��a<��a<��a<ɋa<�a<�  �  �a<�a<5�a<D�a<��a<��a<ʌa</�a<7�a<��a<��a<�a<G�a<]�a<̎a<�a<s�a<��a<��a<F�a<��a<
�a<7�a<a<�a<Y�a<Œa</�a<��a<��a<|�a<Ôa<R�a<��a<$�a<��a<��a<��a<ߗa<o�a<ܘa<c�a<�a<@�a<ǚa<0�a<ԛa<1�a<��a<3�a<��a<�a<p�a<�a<d�a<؟a<O�a<��a<N�a<��a<�a<i�a<�a<P�a<��a<+�a<g�a<Ȥa<�a<��a<�a< �a<��a<��a<7�a<\�a<ħa<��a<:�a<��a<��a<
�a<&�a<~�a<��a<Ωa<��a<:�a<��a<��a<Ѫa<�a<�a<6�a<;�a<��a<m�a<��a<��a<߫a<�a<�a<�a<�a<J�a<-�a<S�a<e�a<>�a<]�a<Z�a<u�a<_�a<d�a<R�a<R�a<e�a<7�a<]�a<&�a<6�a<�a<��a<��a<ګa<ޫa<��a<��a<i�a<v�a<W�a<�a<'�a<תa<Ūa<��a<r�a<^�a<�a<�a<��a<��a<Z�a<=�a<�a<ʨa<��a<J�a<>�a<�a<��a<e�a<*�a<��a<��a<n�a< �a<إa<��a<0�a<��a<��a<\�a<ԣa<��a<5�a<�a<��a<�a<͡a<]�a<%�a<��a<C�a<�a<^�a<�a<��a<E�a<��a<N�a<�a<h�a<&�a<��a<;�a<��a<X�a<�a<a�a<�a<��a<�a<��a<>�a<Ӗa<O�a<��a<g�a<2�a<��a<Z�a<�a<y�a<*�a<��a<f�a<�a<��a<A�a<��a<��a<@�a<�a<��a<g�a<�a<��a<��a<(�a<�a<��a<��a<5�a< �a<�a<��a<��a<O�a<W�a<
�a<�a<�a<��a<��a<��a<��a<y�a<v�a<`�a<b�a<{�a<X�a<��a<l�a<��a<��a<��a<ǋa<ыa<�  �  ��a<�a<:�a<t�a<��a<��a<�a< �a<K�a<{�a<��a<��a<-�a<l�a<Ɏa<�a<P�a<��a<�a<E�a<��a<�a<V�a<��a<�a<}�a<Ғa<.�a<��a<��a<p�a<�a<:�a<��a<'�a<��a<�a<~�a<��a<��a<ޘa<g�a<Ιa<M�a<Κa<V�a<��a</�a<��a<�a<��a<
�a<��a< �a<c�a<�a<X�a<��a<9�a<��a<�a<y�a<ݢa<?�a<��a<�a<~�a<פa<0�a<z�a<�a<)�a<��a<զa<�a<k�a<��a<��a<>�a<t�a<Ѩa<�a<.�a<w�a<��a<�a<�a<A�a<]�a<��a<��a<�a<�a<-�a<P�a<m�a<o�a<��a<��a<ͫa<�a<�a<�a<(�a<!�a<?�a<A�a<J�a<p�a<`�a<]�a<`�a<b�a<Y�a<x�a<V�a<N�a<L�a<9�a<5�a<"�a<�a<#�a<�a<ܫa<̫a<��a<��a<��a<b�a<B�a</�a<��a<�a<��a<��a<u�a<D�a<�a<�a<��a<��a<i�a<9�a<�a<Ҩa<��a<i�a<�a<�a<��a<r�a<(�a<�a<��a<b�a<0�a<��a<��a<3�a<�a<��a<=�a<�a<��a<8�a<�a<��a<+�a<ԡa<��a<��a<��a<=�a<ҟa<t�a<�a<��a<8�a<��a<Y�a<�a<k�a<�a<��a<,�a<��a<G�a<љa<k�a<�a<��a<"�a<��a<0�a<Ԗa<W�a<�a<��a<�a<��a<G�a<ޓa<}�a<�a<ʒa<a�a<�a<��a<=�a<�a<��a<G�a<�a<��a<E�a<�a<��a<}�a<=�a<��a<��a<��a<D�a<�a<�a<��a<��a<h�a<.�a<�a<�a<׋a<݋a<��a<��a<��a<|�a<k�a<��a<e�a<d�a<m�a<j�a<{�a<��a<��a<ŋa<��a<ԋa<�  �  �a<+�a<+�a<h�a<��a<��a<�a<�a<b�a<c�a<��a<�a<4�a<��a<��a<�a<G�a<��a<�a<5�a<��a<�a<j�a<��a<�a<l�a<Ғa<?�a<��a<�a<P�a<�a<8�a<��a<&�a<��a<�a<v�a<��a<a�a<ܘa<m�a<ƙa<l�a<��a<W�a<��a<@�a<��a<$�a<��a<��a<��a<�a<y�a<՟a<C�a<Ҡa<(�a<��a<��a<��a<�a<<�a<ãa<�a<��a<��a<C�a<u�a<�a<1�a<p�a<ۦa<�a<y�a<��a<�a<F�a<q�a<Ψa<�a<N�a<p�a<��a<�a<�a<R�a<T�a<��a<��a<��a<��a<"�a<P�a<`�a<��a<��a<��a<٫a<ݫa<�a<�a<;�a<(�a<L�a<H�a<U�a<h�a<L�a<|�a<T�a<~�a<O�a<_�a<W�a<I�a<[�a<*�a<@�a<"�a<�a<�a<ݫa<��a<��a<̫a<��a<��a<p�a<@�a<=�a<��a<�a<��a<��a<l�a<K�a<,�a<�a<کa<��a<j�a<6�a<��a<�a<��a<}�a<�a<��a<��a<s�a<9�a<�a<��a<B�a<%�a<��a<��a<2�a<Фa<��a<5�a<�a<��a<5�a<��a<z�a<I�a<��a<��a<�a<��a<=�a<ݟa<��a<�a<��a<%�a<Нa<K�a<ٜa<��a< �a<��a<�a<Śa<S�a<ϙa<��a<�a<��a<�a<×a<+�a<Ֆa<`�a<ߕa<��a<�a<��a<6�a<דa<��a<
�a<ǒa<?�a<�a<��a<E�a<��a<��a<X�a<ۏa<��a<E�a<�a<��a<s�a<=�a<�a<΍a<m�a<M�a<�a<׌a<Ìa<m�a<|�a<4�a<)�a<��a<�a<ԋa<��a<��a<|�a<��a<`�a<m�a<f�a<_�a<|�a<[�a<��a<��a<��a<��a<��a<��a<�  �  �a<�a<1�a<Y�a<��a<��a<یa<�a<?�a<y�a<ҍa<�a<1�a<y�a<��a<
�a<O�a<��a<�a<<�a<��a<�a<H�a<��a<#�a<c�a<ɒa<5�a<��a<	�a<j�a<ڔa<L�a<��a<$�a<��a<��a<��a<��a<p�a<�a<`�a<șa<V�a<��a<G�a<ɛa<:�a<��a<)�a<��a<�a<��a<�a<p�a<ޟa<Q�a<Ša<)�a<��a< �a<r�a<�a<>�a<��a<�a<{�a<��a<-�a<x�a<٥a</�a<��a<Ҧa<$�a<W�a<��a<��a<3�a<��a<��a<��a<;�a<e�a<��a<֩a<�a<T�a<o�a<��a<��a<�a<�a<G�a<L�a<h�a<��a<��a<��a<իa<ޫa<�a<�a<�a<1�a<8�a<K�a<d�a<X�a<W�a<i�a<P�a<g�a<`�a<_�a<W�a<N�a<7�a<K�a<%�a<�a<�a<	�a<�a<�a<��a<��a<��a<~�a<{�a<K�a<%�a<	�a<ߪa<��a<��a<j�a<I�a<#�a<�a<̩a<��a<i�a<S�a<��a<Өa<��a<\�a<*�a<�a<��a<j�a</�a<ݦa<��a<\�a<�a<ҥa<{�a<0�a<�a<{�a<D�a<�a<��a<=�a<�a<|�a<3�a<��a<t�a<�a<��a<8�a<�a<j�a<�a<��a<(�a<ǝa<T�a<�a<|�a<�a<��a<>�a<��a<S�a<љa<r�a<�a<��a<	�a<��a</�a<ʖa<]�a<�a<��a<�a<��a<O�a<�a<r�a<�a<��a<S�a<��a<��a<B�a<�a<��a<Z�a<��a<��a<M�a<�a<��a<��a<9�a<��a<��a<�a<K�a<�a<،a<ьa<��a<X�a<>�a<�a<��a<�a<ŋa<��a<��a<w�a<��a<q�a<m�a<f�a<d�a<X�a<|�a<k�a<�a<��a<��a<��a<ދa<�  �  �a<��a<H�a<j�a<o�a<��a<܌a<#�a<>�a<��a<��a<��a<B�a<l�a<َa<�a<h�a<��a<�a<C�a<��a<�a<E�a<��a<�a<��a<גa<'�a<��a<�a<z�a<ʔa<P�a<��a<�a<��a<�a<��a<�a<|�a<ߘa<c�a<�a<>�a<�a<;�a<��a<$�a<��a<.�a<��a<�a<h�a<�a<i�a<�a<c�a<��a<L�a<��a<�a<h�a<�a<J�a<��a<�a<i�a<�a<�a<��a<�a<"�a<��a<��a<=�a<R�a<��a<�a<7�a<��a<��a<�a<#�a<��a<��a<ݩa<&�a<(�a<i�a<��a<˪a<�a<�a<)�a<8�a<��a<t�a<��a<��a<ܫa<�a<�a<�a<�a<@�a<:�a<A�a<>�a<^�a<r�a<I�a<}�a<[�a<c�a<`�a<J�a<o�a<0�a<N�a<�a<=�a<�a<�a<��a<֫a<�a<��a<��a<��a<P�a<F�a<&�a<�a<ުa<̪a<��a<x�a<Y�a<�a<�a<��a<��a<^�a<.�a<�a<Ψa<��a<X�a<&�a<ѧa<ħa<w�a<"�a<�a<��a<l�a<�a<֥a<��a<!�a<�a<y�a<c�a<ۣa<��a<8�a<�a<��a<�a<�a<h�a< �a<��a<>�a<�a<`�a<�a<��a<E�a<��a<`�a<��a<q�a<$�a<�a<5�a<��a<T�a<ܙa<]�a<�a<��a<4�a<��a<D�a<֖a<P�a<��a<q�a<8�a<��a<F�a<Փa<v�a<)�a<��a<d�a<�a<��a<A�a<�a<��a<.�a<��a<��a<b�a<�a<��a<z�a<%�a<�a<��a<��a<C�a<�a<�a<��a<��a<X�a<L�a<�a<�a<ʋa<ʋa<Ëa<��a<��a<u�a<t�a<n�a<Y�a<��a<Q�a<�a<^�a<��a<��a<��a<a<͋a<�  �  ��a<�a<3�a<U�a<��a<όa<�a<�a<P�a<��a<��a<�a<;�a<l�a<��a<��a<^�a<��a<�a<U�a<��a<�a<]�a<Ǒa<�a<h�a<̒a<)�a<��a<��a<t�a<Քa<6�a<��a<#�a<��a<�a<~�a<ۗa<p�a<ژa<S�a<ٙa<L�a<��a<9�a<˛a<S�a<��a<'�a<��a<�a<��a<�a<i�a<ٟa<K�a<��a<G�a<��a<�a<��a<�a<K�a<ʣa<$�a<l�a<Ťa<&�a<��a<ҥa<#�a<��a<��a<�a<m�a<��a<��a<D�a<q�a<��a<�a<,�a<r�a<��a<שa<�a<5�a<��a<��a<��a<�a<�a<4�a<T�a<}�a<��a<��a<��a<ګa<��a<��a<�a<,�a</�a<E�a<k�a<W�a<M�a<X�a<[�a<l�a<V�a<\�a<a�a<=�a<S�a<C�a<@�a<)�a<*�a<��a<
�a<��a<ԫa<իa<��a<��a<z�a<f�a<f�a<2�a<�a<�a<ʪa<��a<��a<R�a<�a<��a<��a<��a<s�a<:�a<�a<Ҩa<��a<q�a<D�a<�a<��a<m�a<#�a<�a<��a<f�a<�a<��a<��a</�a<�a<��a<=�a<Уa<��a<3�a<ڢa<��a<)�a<ǡa<e�a<�a<Ƞa<F�a<��a<|�a<�a<��a<F�a<��a<O�a<�a<s�a<�a<��a<6�a<Śa<Q�a<ݙa<��a<�a<��a<�a<��a<8�a<Öa<Q�a<�a<k�a<�a<��a<J�a<�a<��a<�a<��a<^�a<�a<��a<:�a<�a<��a<;�a<�a<��a<S�a<
�a<юa<��a<B�a<�a<��a<��a<?�a<�a<��a<��a<��a<l�a<<�a<"�a<�a<�a<��a<��a<��a<��a<p�a<n�a<o�a<M�a<i�a<d�a<r�a<o�a<��a<}�a<��a<��a<ˋa<�  �  ߋa<0�a<?�a<]�a<��a<��a<֌a<	�a<L�a<r�a<̍a<�a<*�a<��a<��a<%�a<?�a<��a<��a<E�a<��a<�a<E�a<��a< �a<f�a<ߒa<C�a<��a<�a<[�a<�a<D�a<��a<�a<��a<�a<n�a<�a<g�a<�a<d�a<˙a<m�a<��a<O�a<��a<(�a<��a<�a<��a<�a<��a<�a<�a<�a<X�a<۠a<�a<��a<�a<}�a<ޢa<:�a<��a<�a<��a<Ĥa<I�a<��a<٥a<4�a<w�a<�a<�a<e�a<��a<�a<6�a<v�a<ͨa<�a<D�a<e�a<��a<��a<�a<R�a<W�a<��a<��a<�a<�a<-�a<M�a<S�a<��a<��a<ӫa<ԫa<׫a<�a<�a<'�a<)�a<1�a<;�a<W�a<]�a<b�a<~�a<K�a<q�a<X�a<^�a<e�a<<�a<@�a</�a<,�a<�a<�a<�a<�a<�a<��a<ѫa<��a<��a<u�a<8�a<�a< �a<�a<��a<��a<e�a<A�a<<�a<�a<�a<��a<f�a<A�a<�a<Ψa<��a<X�a<�a<�a<��a<��a<>�a<ۦa<��a<M�a<#�a<ɥa<v�a<*�a<֤a<��a<-�a<�a<��a<@�a<�a<~�a<K�a<ȡa<{�a<�a<��a<2�a<՟a<y�a<��a<��a<�a<֝a<c�a<�a<��a<�a<��a<#�a<��a<H�a<̙a<a�a<�a<��a<�a<ȗa<8�a<ʖa<b�a<�a<��a<�a<��a<7�a<ԓa<u�a<�a<ƒa<I�a<�a<��a<O�a<�a<��a<X�a<ޏa<��a<I�a<�a<Ǝa<~�a<:�a<�a<ݍa<w�a<a�a<�a<ьa<͌a<|�a<h�a<5�a<�a<�a<�a<ɋa<��a<��a<r�a<��a<i�a<l�a<t�a<R�a<a�a<`�a<r�a<u�a<��a<��a<��a<�a<�  �  �a<�a<%�a<_�a<��a<��a<��a<&�a<S�a<t�a<��a<��a<3�a<��a<��a<�a<K�a<��a<�a<C�a<��a<�a<^�a<��a<�a<d�a<��a<&�a<��a<�a<X�a<Ĕa<=�a<��a<,�a<��a<�a<z�a<�a<W�a<ޘa<c�a<șa<A�a<��a<I�a<��a<<�a<a<1�a<��a<�a<��a<��a<t�a<ܟa<J�a<͠a<4�a<��a<�a<��a<�a<b�a<��a<�a<x�a<��a<�a<v�a<ڥa<'�a<k�a<��a<�a<k�a<��a<��a<:�a<v�a<��a<�a<6�a<k�a<��a<˩a<��a<C�a<g�a<��a<تa<�a<�a<+�a<\�a<c�a<��a<��a<ūa<ԫa<�a<�a<�a<-�a<D�a<S�a<N�a<T�a<]�a<K�a<U�a<Z�a<n�a<U�a<K�a<O�a<O�a<P�a<B�a<9�a<#�a<�a<��a<�a<�a<ƫa<��a<��a<��a<m�a<K�a<@�a<�a<��a<��a<��a<}�a<J�a<2�a<�a<թa<��a<y�a<:�a<�a<ݨa<��a<q�a<$�a<�a<��a<\�a<!�a<�a<��a<J�a<�a<åa<}�a<8�a<�a<��a<9�a<�a<��a<7�a<�a<|�a<�a<��a<u�a<�a<��a<Y�a<�a<|�a<��a<��a<4�a<˝a<R�a<��a<��a<�a<��a<%�a<Úa<Y�a<��a<u�a<��a<��a<�a<��a<,�a<˖a<V�a<ڕa<u�a<�a<��a<J�a<�a<z�a<�a<��a<D�a<��a<��a<7�a<ܐa<��a<I�a<�a<��a<o�a<�a<Ďa<{�a<I�a<�a<ɍa<q�a<S�a<�a<�a<Ìa<~�a<m�a<Q�a<0�a<�a<�a<ʋa<��a<��a<��a<��a<g�a<Y�a<^�a<e�a<q�a<s�a<�a<��a<��a<��a<��a<��a<�  �  �a<�a<B�a<i�a<y�a<��a<ڌa<��a<I�a<��a<��a<�a<'�a<��a<�a<�a<E�a<��a<��a<O�a<��a<�a<D�a<��a<��a<�a<ݒa<B�a<��a<�a<��a<ߔa<D�a<��a<�a<��a<�a<��a<�a<��a<�a<P�a<�a<]�a<Ԛa<;�a<��a<3�a<��a<�a<��a<�a<��a<
�a<d�a<��a<q�a<��a<?�a<��a<�a<��a<֢a<A�a<��a<�a<e�a<ޤa<:�a<��a<֥a<0�a<��a<æa<�a<^�a<��a<�a<3�a<~�a<��a<�a<&�a<y�a<��a<�a<!�a<2�a<t�a<��a<��a<ܪa<�a<0�a<[�a<a�a<��a<ƫa<̫a<ȫa<�a<��a<�a<(�a<�a<4�a<Q�a<I�a<b�a<i�a<k�a<w�a<I�a<k�a<v�a<F�a<S�a<;�a<*�a<#�a<%�a<�a<�a<�a<ƫa<ޫa<��a<��a<��a<Z�a<R�a<#�a<�a<�a<ƪa<��a<��a<?�a<,�a<�a<ǩa<��a<�a<7�a<�a<Шa<��a<X�a<3�a<�a<§a<}�a<<�a<��a<��a<y�a<�a<ʥa<}�a<%�a<Фa<��a<B�a<ݣa<��a<E�a<آa<��a<:�a<ۡa<g�a<�a<��a<9�a<̟a<|�a<	�a<��a<A�a<��a<q�a<�a<p�a<�a<��a<.�a<Ța<@�a<ԙa<e�a<��a<�a<)�a<��a<Q�a<ǖa<_�a<�a<v�a<�a<��a<7�a<ԓa<s�a<�a<��a<t�a<�a<��a<V�a<��a<��a<8�a<��a<��a<I�a<�a<͎a<��a<H�a<�a<��a<��a<Y�a<	�a<��a<��a<��a<h�a<*�a<�a<�a<֋a<΋a<��a<��a<��a<c�a<}�a<��a<V�a<i�a<\�a<[�a<i�a<��a<��a<��a<ыa<��a<�  �  �a<�a<%�a<_�a<��a<��a<��a<&�a<S�a<t�a<��a<��a<3�a<��a<��a<�a<K�a<��a<�a<C�a<��a<�a<^�a<��a<�a<d�a<��a<&�a<��a<�a<X�a<Ĕa<=�a<��a<,�a<��a<�a<z�a<�a<W�a<ޘa<c�a<șa<A�a<��a<I�a<��a<<�a<a<1�a<��a<�a<��a<��a<t�a<ܟa<J�a<͠a<4�a<��a<�a<��a<�a<b�a<��a<�a<x�a<��a<�a<v�a<ڥa<'�a<k�a<��a<�a<k�a<��a<��a<:�a<v�a<��a<�a<6�a<k�a<��a<˩a<��a<C�a<g�a<��a<تa<�a<�a<+�a<\�a<c�a<��a<��a<ūa<ԫa<�a<�a<�a<-�a<D�a<S�a<N�a<T�a<]�a<K�a<U�a<Z�a<n�a<U�a<K�a<O�a<O�a<P�a<B�a<9�a<#�a<�a<��a<�a<�a<ƫa<��a<��a<��a<m�a<K�a<@�a<�a<��a<��a<��a<}�a<J�a<2�a<�a<թa<��a<y�a<:�a<�a<ݨa<��a<q�a<$�a<�a<��a<\�a<!�a<�a<��a<J�a<�a<åa<}�a<8�a<�a<��a<9�a<�a<��a<7�a<�a<|�a<�a<��a<u�a<�a<��a<Y�a<�a<|�a<��a<��a<4�a<˝a<R�a<��a<��a<�a<��a<%�a<Úa<Y�a<��a<u�a<��a<��a<�a<��a<,�a<˖a<V�a<ڕa<u�a<�a<��a<J�a<�a<z�a<�a<��a<D�a<��a<��a<7�a<ܐa<��a<I�a<�a<��a<o�a<�a<Ďa<{�a<I�a<�a<ɍa<q�a<S�a<�a<�a<Ìa<~�a<m�a<Q�a<0�a<�a<�a<ʋa<��a<��a<��a<��a<g�a<Y�a<^�a<e�a<q�a<s�a<�a<��a<��a<��a<��a<��a<�  �  ߋa<0�a<?�a<]�a<��a<��a<֌a<	�a<L�a<r�a<̍a<�a<*�a<��a<��a<%�a<?�a<��a<��a<E�a<��a<�a<E�a<��a< �a<f�a<ߒa<C�a<��a<�a<[�a<�a<D�a<��a<�a<��a<�a<n�a<�a<g�a<�a<d�a<˙a<m�a<��a<O�a<��a<(�a<��a<�a<��a<�a<��a<�a<�a<�a<X�a<۠a<�a<��a<�a<}�a<ޢa<:�a<��a<�a<��a<Ĥa<I�a<��a<٥a<4�a<w�a<�a<�a<e�a<��a<�a<6�a<v�a<ͨa<�a<D�a<e�a<��a<��a<�a<R�a<W�a<��a<��a<�a<�a<-�a<M�a<S�a<��a<��a<ӫa<ԫa<׫a<�a<�a<'�a<)�a<1�a<;�a<W�a<]�a<b�a<~�a<K�a<q�a<X�a<^�a<e�a<<�a<@�a</�a<,�a<�a<�a<�a<�a<�a<��a<ѫa<��a<��a<u�a<8�a<�a< �a<�a<��a<��a<e�a<A�a<<�a<�a<�a<��a<f�a<A�a<�a<Ψa<��a<X�a<�a<�a<��a<��a<>�a<ۦa<��a<M�a<#�a<ɥa<v�a<*�a<֤a<��a<-�a<�a<��a<@�a<�a<~�a<K�a<ȡa<{�a<�a<��a<2�a<՟a<y�a<��a<��a<�a<֝a<c�a<�a<��a<�a<��a<#�a<��a<H�a<̙a<a�a<�a<��a<�a<ȗa<8�a<ʖa<b�a<�a<��a<�a<��a<7�a<ԓa<u�a<�a<ƒa<I�a<�a<��a<O�a<�a<��a<X�a<ޏa<��a<I�a<�a<Ǝa<~�a<:�a<�a<ݍa<w�a<a�a<�a<ьa<͌a<|�a<h�a<5�a<�a<�a<�a<ɋa<��a<��a<r�a<��a<i�a<l�a<t�a<R�a<a�a<`�a<r�a<u�a<��a<��a<��a<�a<�  �  ��a<�a<3�a<U�a<��a<όa<�a<�a<P�a<��a<��a<�a<;�a<l�a<��a<��a<^�a<��a<�a<U�a<��a<�a<]�a<Ǒa<�a<h�a<̒a<)�a<��a<��a<t�a<Քa<6�a<��a<#�a<��a<�a<~�a<ۗa<p�a<ژa<S�a<ٙa<L�a<��a<9�a<˛a<S�a<��a<'�a<��a<�a<��a<�a<i�a<ٟa<K�a<��a<G�a<��a<�a<��a<�a<K�a<ʣa<$�a<l�a<Ťa<&�a<��a<ҥa<#�a<��a<��a<�a<m�a<��a<��a<D�a<q�a<��a<�a<,�a<r�a<��a<שa<�a<5�a<��a<��a<��a<�a<�a<4�a<T�a<}�a<��a<��a<��a<ګa<��a<��a<�a<,�a</�a<E�a<k�a<W�a<M�a<X�a<[�a<l�a<V�a<\�a<a�a<=�a<S�a<C�a<@�a<)�a<*�a<��a<
�a<��a<ԫa<իa<��a<��a<z�a<f�a<f�a<2�a<�a<�a<ʪa<��a<��a<R�a<�a<��a<��a<��a<s�a<:�a<�a<Ҩa<��a<q�a<D�a<�a<��a<m�a<#�a<�a<��a<f�a<�a<��a<��a</�a<�a<��a<=�a<Уa<��a<3�a<ڢa<��a<)�a<ǡa<e�a<�a<Ƞa<F�a<��a<|�a<�a<��a<F�a<��a<O�a<�a<s�a<�a<��a<6�a<Śa<Q�a<ݙa<��a<�a<��a<�a<��a<8�a<Öa<Q�a<�a<k�a<�a<��a<J�a<�a<��a<�a<��a<^�a<�a<��a<:�a<�a<��a<;�a<�a<��a<S�a<
�a<юa<��a<B�a<�a<��a<��a<?�a<�a<��a<��a<��a<l�a<<�a<"�a<�a<�a<��a<��a<��a<��a<p�a<n�a<o�a<M�a<i�a<d�a<r�a<o�a<��a<}�a<��a<��a<ˋa<�  �  �a<��a<H�a<j�a<o�a<��a<܌a<#�a<>�a<��a<��a<��a<B�a<l�a<َa<�a<h�a<��a<�a<C�a<��a<�a<E�a<��a<�a<��a<גa<'�a<��a<�a<z�a<ʔa<P�a<��a<�a<��a<�a<��a<�a<|�a<ߘa<c�a<�a<>�a<�a<;�a<��a<$�a<��a<.�a<��a<�a<h�a<�a<i�a<�a<c�a<��a<L�a<��a<�a<h�a<�a<J�a<��a<�a<i�a<�a<�a<��a<�a<"�a<��a<��a<=�a<R�a<��a<�a<7�a<��a<��a<�a<#�a<��a<��a<ݩa<&�a<(�a<i�a<��a<˪a<�a<�a<)�a<8�a<��a<t�a<��a<��a<ܫa<�a<�a<�a<�a<@�a<:�a<A�a<>�a<^�a<r�a<I�a<}�a<[�a<c�a<`�a<J�a<o�a<0�a<N�a<�a<=�a<�a<�a<��a<֫a<�a<��a<��a<��a<P�a<F�a<&�a<�a<ުa<̪a<��a<x�a<Y�a<�a<�a<��a<��a<^�a<.�a<�a<Ψa<��a<X�a<&�a<ѧa<ħa<w�a<"�a<�a<��a<l�a<�a<֥a<��a<!�a<�a<y�a<c�a<ۣa<��a<8�a<�a<��a<�a<�a<h�a< �a<��a<>�a<�a<`�a<�a<��a<E�a<��a<`�a<��a<q�a<$�a<�a<5�a<��a<T�a<ܙa<]�a<�a<��a<4�a<��a<D�a<֖a<P�a<��a<q�a<8�a<��a<F�a<Փa<v�a<)�a<��a<d�a<�a<��a<A�a<�a<��a<.�a<��a<��a<b�a<�a<��a<z�a<%�a<�a<��a<��a<C�a<�a<�a<��a<��a<X�a<L�a<�a<�a<ʋa<ʋa<Ëa<��a<��a<u�a<t�a<n�a<Y�a<��a<Q�a<�a<^�a<��a<��a<��a<a<͋a<�  �  �a<�a<1�a<Y�a<��a<��a<یa<�a<?�a<y�a<ҍa<�a<1�a<y�a<��a<
�a<O�a<��a<�a<<�a<��a<�a<H�a<��a<#�a<c�a<ɒa<5�a<��a<	�a<j�a<ڔa<L�a<��a<$�a<��a<��a<��a<��a<p�a<�a<`�a<șa<V�a<��a<G�a<ɛa<:�a<��a<)�a<��a<�a<��a<�a<p�a<ޟa<Q�a<Ša<)�a<��a< �a<r�a<�a<>�a<��a<�a<{�a<��a<-�a<x�a<٥a</�a<��a<Ҧa<$�a<W�a<��a<��a<3�a<��a<��a<��a<;�a<e�a<��a<֩a<�a<T�a<o�a<��a<��a<�a<�a<G�a<L�a<h�a<��a<��a<��a<իa<ޫa<�a<�a<�a<1�a<8�a<K�a<d�a<X�a<W�a<i�a<P�a<g�a<`�a<_�a<W�a<N�a<7�a<K�a<%�a<�a<�a<	�a<�a<�a<��a<��a<��a<~�a<{�a<K�a<%�a<	�a<ߪa<��a<��a<j�a<I�a<#�a<�a<̩a<��a<i�a<S�a<��a<Өa<��a<\�a<*�a<�a<��a<j�a</�a<ݦa<��a<\�a<�a<ҥa<{�a<0�a<�a<{�a<D�a<�a<��a<=�a<�a<|�a<3�a<��a<t�a<�a<��a<8�a<�a<j�a<�a<��a<(�a<ǝa<T�a<�a<|�a<�a<��a<>�a<��a<S�a<љa<r�a<�a<��a<	�a<��a</�a<ʖa<]�a<�a<��a<�a<��a<O�a<�a<r�a<�a<��a<S�a<��a<��a<B�a<�a<��a<Z�a<��a<��a<M�a<�a<��a<��a<9�a<��a<��a<�a<K�a<�a<،a<ьa<��a<X�a<>�a<�a<��a<�a<ŋa<��a<��a<w�a<��a<q�a<m�a<f�a<d�a<X�a<|�a<k�a<�a<��a<��a<��a<ދa<�  �  �a<+�a<+�a<h�a<��a<��a<�a<�a<b�a<c�a<��a<�a<4�a<��a<��a<�a<G�a<��a<�a<5�a<��a<�a<j�a<��a<�a<l�a<Ғa<?�a<��a<�a<P�a<�a<8�a<��a<&�a<��a<�a<v�a<��a<a�a<ܘa<m�a<ƙa<l�a<��a<W�a<��a<@�a<��a<$�a<��a<��a<��a<�a<y�a<՟a<C�a<Ҡa<(�a<��a<��a<��a<�a<<�a<ãa<�a<��a<��a<C�a<u�a<�a<1�a<p�a<ۦa<�a<y�a<��a<�a<F�a<q�a<Ψa<�a<N�a<p�a<��a<�a<�a<R�a<T�a<��a<��a<��a<��a<"�a<P�a<`�a<��a<��a<��a<٫a<ݫa<�a<�a<;�a<(�a<L�a<H�a<U�a<h�a<L�a<|�a<T�a<~�a<O�a<_�a<W�a<I�a<[�a<*�a<@�a<"�a<�a<�a<ݫa<��a<��a<̫a<��a<��a<p�a<@�a<=�a<��a<�a<��a<��a<l�a<K�a<,�a<�a<کa<��a<j�a<6�a<��a<�a<��a<}�a<�a<��a<��a<s�a<9�a<�a<��a<B�a<%�a<��a<��a<2�a<Фa<��a<5�a<�a<��a<5�a<��a<z�a<I�a<��a<��a<�a<��a<=�a<ݟa<��a<�a<��a<%�a<Нa<K�a<ٜa<��a< �a<��a<�a<Śa<S�a<ϙa<��a<�a<��a<�a<×a<+�a<Ֆa<`�a<ߕa<��a<�a<��a<6�a<דa<��a<
�a<ǒa<?�a<�a<��a<E�a<��a<��a<X�a<ۏa<��a<E�a<�a<��a<s�a<=�a<�a<΍a<m�a<M�a<�a<׌a<Ìa<m�a<|�a<4�a<)�a<��a<�a<ԋa<��a<��a<|�a<��a<`�a<m�a<f�a<_�a<|�a<[�a<��a<��a<��a<��a<��a<��a<�  �  ��a<�a<:�a<t�a<��a<��a<�a< �a<K�a<{�a<��a<��a<-�a<l�a<Ɏa<�a<P�a<��a<�a<E�a<��a<�a<V�a<��a<�a<}�a<Ғa<.�a<��a<��a<p�a<�a<:�a<��a<'�a<��a<�a<~�a<��a<��a<ޘa<g�a<Ιa<M�a<Κa<V�a<��a</�a<��a<�a<��a<
�a<��a< �a<c�a<�a<X�a<��a<9�a<��a<�a<y�a<ݢa<?�a<��a<�a<~�a<פa<0�a<z�a<�a<)�a<��a<զa<�a<k�a<��a<��a<>�a<t�a<Ѩa<�a<.�a<w�a<��a<�a<�a<A�a<]�a<��a<��a<�a<�a<-�a<P�a<m�a<o�a<��a<��a<ͫa<�a<�a<�a<(�a<!�a<?�a<A�a<J�a<p�a<`�a<]�a<`�a<b�a<Y�a<x�a<V�a<N�a<L�a<9�a<5�a<"�a<�a<#�a<�a<ܫa<̫a<��a<��a<��a<b�a<B�a</�a<��a<�a<��a<��a<u�a<D�a<�a<�a<��a<��a<i�a<9�a<�a<Ҩa<��a<i�a<�a<�a<��a<r�a<(�a<�a<��a<b�a<0�a<��a<��a<3�a<�a<��a<=�a<�a<��a<8�a<�a<��a<+�a<ԡa<��a<��a<��a<=�a<ҟa<t�a<�a<��a<8�a<��a<Y�a<�a<k�a<�a<��a<,�a<��a<G�a<љa<k�a<�a<��a<"�a<��a<0�a<Ԗa<W�a<�a<��a<�a<��a<G�a<ޓa<}�a<�a<ʒa<a�a<�a<��a<=�a<�a<��a<G�a<�a<��a<E�a<�a<��a<}�a<=�a<��a<��a<��a<D�a<�a<�a<��a<��a<h�a<.�a<�a<�a<׋a<݋a<��a<��a<��a<|�a<k�a<��a<e�a<d�a<m�a<j�a<{�a<��a<��a<ŋa<��a<ԋa<�  �  �a<�a<5�a<D�a<��a<��a<ʌa</�a<7�a<��a<��a<�a<G�a<]�a<̎a<�a<s�a<��a<��a<F�a<��a<
�a<7�a<a<�a<Y�a<Œa</�a<��a<��a<|�a<Ôa<R�a<��a<$�a<��a<��a<��a<ߗa<o�a<ܘa<c�a<�a<@�a<ǚa<0�a<ԛa<1�a<��a<3�a<��a<�a<p�a<�a<d�a<؟a<O�a<��a<N�a<��a<�a<i�a<�a<P�a<��a<+�a<g�a<Ȥa<�a<��a<�a< �a<��a<��a<7�a<\�a<ħa<��a<:�a<��a<��a<
�a<&�a<~�a<��a<Ωa<��a<:�a<��a<��a<Ѫa<�a<�a<6�a<;�a<��a<m�a<��a<��a<߫a<�a<�a<�a<�a<J�a<-�a<S�a<e�a<>�a<]�a<Z�a<u�a<_�a<d�a<R�a<R�a<e�a<7�a<]�a<&�a<6�a<�a<��a<��a<ګa<ޫa<��a<��a<i�a<v�a<W�a<�a<'�a<תa<Ūa<��a<r�a<^�a<�a<�a<��a<��a<Z�a<=�a<�a<ʨa<��a<J�a<>�a<�a<��a<e�a<*�a<��a<��a<n�a< �a<إa<��a<0�a<��a<��a<\�a<ԣa<��a<5�a<�a<��a<�a<͡a<]�a<%�a<��a<C�a<�a<^�a<�a<��a<E�a<��a<N�a<�a<h�a<&�a<��a<;�a<��a<X�a<�a<a�a<�a<��a<�a<��a<>�a<Ӗa<O�a<��a<g�a<2�a<��a<Z�a<�a<y�a<*�a<��a<f�a<�a<��a<A�a<��a<��a<@�a<�a<��a<g�a<�a<��a<��a<(�a<�a<��a<��a<5�a< �a<�a<��a<��a<O�a<W�a<
�a<�a<�a<��a<��a<��a<��a<y�a<v�a<`�a<b�a<{�a<X�a<��a<l�a<��a<��a<��a<ǋa<ыa<�  �  �a<�a<T�a<Z�a<��a<��a<֌a<�a<8�a<�a<��a<ݍa<:�a<m�a<��a< �a<S�a<��a<�a<>�a<��a<��a<J�a<��a<��a<u�a<�a<:�a<��a<�a<t�a<ؔa<[�a<��a<�a<��a<�a<��a<��a<y�a<�a<]�a<ԙa<e�a<��a<9�a<��a<-�a<��a<!�a<��a<�a<t�a<�a<u�a<�a<V�a<ɠa<,�a<��a<�a<m�a<ܢa<E�a<��a<�a<j�a<�a<E�a<��a<ޥa<9�a<��a<֦a<2�a<a�a<��a<�a<:�a<��a<��a<�a<A�a<u�a<��a<��a<�a<3�a<c�a<��a<êa<تa< �a<.�a<0�a<j�a<��a<��a<��a<ܫa<ثa<��a<�a<�a<8�a<2�a<F�a<N�a<S�a<{�a<o�a<_�a<g�a<o�a<]�a<d�a<\�a<@�a<B�a<)�a</�a<(�a<�a<��a<�a<ɫa<��a<��a<�a<a�a<E�a<�a<�a<تa<Īa<��a<]�a<Q�a<�a<��a<éa<��a<N�a<:�a<��a<èa<��a<]�a<!�a<�a<��a<��a<5�a<�a<��a<f�a<�a<�a<��a<(�a<�a<��a<T�a<��a<��a<L�a<�a<��a<C�a<�a<f�a<�a<��a<8�a<ڟa<g�a<�a<��a<&�a<̝a<Z�a<�a<�a<�a<��a</�a<��a<F�a<יa<f�a<�a<��a</�a<ŗa<:�a<ϖa<g�a<��a<��a<-�a<��a<@�a<דa<y�a<-�a<��a<a�a<�a<��a<I�a<�a<��a<9�a<�a<��a<Z�a<��a<��a<~�a<�a<��a<��a<��a<C�a<�a<Ҍa<��a<��a<T�a<E�a<�a<��a<ۋa<��a<ˋa<��a<��a<��a<��a<k�a<s�a<r�a<a�a<s�a<o�a<��a<��a<��a<ɋa<�a<�  �  �a<�a<%�a<o�a<��a<��a<��a<��a<S�a<o�a<��a<��a<&�a<p�a<��a<��a<=�a<��a<�a<>�a<��a<ݐa<k�a<��a<�a<m�a<Òa<%�a<��a<	�a<^�a<�a<3�a<��a<=�a<��a<,�a<g�a<��a<l�a<�a<[�a<əa<G�a<��a<V�a<��a<N�a<��a<�a<��a<�a<��a<�a<i�a<ҟa<B�a<��a<"�a<��a<�a<~�a<ݢa<J�a<ˣa<�a<��a<��a<"�a<t�a<إa<3�a<y�a<ئa< �a<��a<��a<�a<J�a<j�a<Өa<�a<>�a<j�a<��a<ѩa<�a<H�a<e�a<��a<��a<�a<	�a<'�a<a�a<X�a<��a<��a<��a<ȫa<�a<
�a< �a</�a<�a<O�a<U�a<O�a<o�a<J�a<X�a<Z�a<d�a<_�a<j�a<Q�a<A�a<g�a<)�a<P�a<�a<�a<�a<�a<�a<īa<��a<��a<��a<g�a<Q�a<B�a<�a<�a<��a<��a<w�a<=�a<�a<�a<��a<��a<y�a<8�a<��a<ܨa<��a<�a<)�a<�a<��a<c�a< �a<�a<��a<P�a<.�a<��a<��a<I�a<ޤa<��a<&�a<�a<��a<D�a<�a<}�a<%�a<��a<��a<�a<àa<I�a<ҟa<}�a<��a<��a<&�a<��a<H�a<ٜa<v�a<��a<��a<!�a<a<G�a<ܙa<��a<�a<��a<	�a<��a<+�a<ɖa<b�a<�a<��a<��a<ʔa<I�a<�a<��a<�a<̒a<I�a<�a<��a<5�a<�a<��a<N�a<�a<��a<E�a<�a<a<x�a<N�a<�a<��a<s�a<A�a<
�a<�a<��a<y�a<p�a<+�a<-�a<�a<܋a<ۋa<��a<��a<��a<~�a<q�a<x�a<a�a<W�a<��a<Z�a<��a<x�a<��a<��a<��a<ߋa<�  �  �a<+�a<7�a<e�a<��a<��a<֌a<�a<L�a<j�a<��a<�a<2�a<}�a<��a<�a<O�a<��a<ޏa<:�a<��a<�a<B�a<��a<�a<l�a<Ւa<H�a<��a<�a<a�a<�a<L�a<��a<,�a<��a<�a<z�a<�a<k�a<�a<k�a<�a<\�a<Śa<G�a<��a<"�a<��a<�a<��a<��a<t�a<�a<m�a<�a<V�a<Ġa<)�a<��a<��a<r�a<ߢa<:�a<��a<��a<w�a<Τa<6�a<��a<�a<5�a<z�a<�a<�a<s�a<��a<��a<A�a<��a<ͨa<�a<A�a<�a<��a<�a<�a<C�a<W�a<��a<��a<�a<�a<�a<@�a<e�a<��a<��a<��a<ҫa<�a<�a<��a<'�a<*�a<1�a<4�a<N�a<a�a<[�a<s�a<|�a<q�a<]�a<a�a<f�a<M�a<V�a<*�a<C�a<$�a<#�a<�a<�a<�a<�a<̫a<��a<��a<h�a<6�a<�a<�a<�a<��a<��a<k�a<I�a<'�a<��a<Ωa<��a<_�a<%�a<��a<ڨa<��a<V�a<�a<�a<��a<u�a<C�a<��a<��a<S�a<$�a<ҥa<��a<8�a<֤a<��a<9�a<��a<��a<C�a<�a<��a<:�a<ˡa<s�a<��a<��a<3�a<֟a<n�a<��a<��a<)�a<ĝa<\�a<�a<{�a<�a<��a<�a<��a<I�a<͙a<Y�a<�a<��a<�a<��a<T�a<ٖa<d�a<�a<��a<�a<��a<=�a<ޓa<��a<�a<ƒa<J�a<�a<��a<[�a<��a<��a<I�a<ߏa<��a<G�a<�a<��a<f�a<-�a<�a<a<��a<O�a<�a<یa<��a<v�a<h�a<6�a<�a<�a<ۋa<͋a<��a<��a<��a<��a<o�a<o�a<v�a<c�a<w�a<[�a<��a<��a<��a<��a<��a<�a<�  �  ��a<��a<�a<�a<:�a<{�a<��a<эa<ٍa<?�a<g�a<��a<�a<%�a<��a<��a<�a<N�a<��a<��a<-�a<��a<�a<o�a<��a< �a<d�a<ϓa<E�a<��a<0�a<q�a<��a<F�a<͖a<I�a<��a<#�a<��a<�a<��a<��a<v�a<Śa<y�a<Лa<_�a<֜a<?�a<��a<�a<��a<�a<��a<�a<o�a<�a<<�a<ܡa< �a<��a<�a<]�a<Уa<C�a<��a<�a<l�a<��a<�a<\�a<˦a<�a<I�a<��a<ܧa<E�a<��a<��a<�a<5�a<��a<ϩa<��a<�a<=�a<��a<��a<�a< �a<I�a<S�a<��a<��a<ͫa<�a<��a<3�a<C�a<W�a<|�a<y�a<��a<��a<��a<ˬa<�a<ݬa<֬a<��a<Ȭa<�a<��a<�a<ܬa<�a<Ӭa<Ǭa<Ӭa<��a<��a<��a<��a<��a<{�a<U�a<"�a<*�a<�a<�a<�a<��a<��a<M�a<X�a< �a<�a<تa<��a<��a<@�a<3�a<�a<̩a<��a<;�a<,�a<�a<ƨa<k�a<?�a<�a<��a<t�a<A�a<�a<��a<c�a<��a<��a<y�a<�a<ɤa<p�a<�a<�a<s�a<�a<��a<p�a<�a<��a<A�a<Πa<f�a<�a<��a<�a<ߞa<E�a<�a<}�a<��a<��a<%�a<ԛa<@�a<ךa<u�a<�a<��a<�a<Ϙa< �a<חa<i�a<�a<��a<�a<��a<D�a<��a<��a<�a<ȓa<T�a<�a<��a<M�a<�a<x�a<R�a<�a<��a<X�a<�a<��a<n�a<:�a<�a<a<\�a<?�a<��a<ƍa<��a<_�a<Q�a<��a<��a<׌a<Ča<��a<r�a<u�a<0�a<B�a<A�a<G�a<�a<'�a<�a<�a<2�a<%�a<0�a<[�a<U�a<��a<��a<�  �  ��a<�a<��a<�a<<�a<b�a<��a<Ía<�a<9�a<f�a<��a<ێa<$�a<m�a<��a<��a<L�a<��a<��a<Y�a<��a<�a<W�a<��a<$�a<��a<��a<C�a<��a<�a<��a<��a<j�a<֖a<1�a<Ɨa<5�a<��a<�a<��a<�a<��a<��a<n�a<ߛa<N�a<��a<4�a<��a<,�a<��a<�a<��a<�a<q�a<�a<G�a<��a<'�a<��a<��a<v�a<ţa<&�a<��a<��a<a�a<��a<#�a<P�a<��a<��a<n�a<��a< �a<,�a<|�a<Ϩa<�a<N�a<~�a<��a<�a<J�a<k�a<��a<Ūa<�a<�a<=�a<w�a<��a<��a<Ϋa<�a<�a<'�a<@�a<M�a<n�a<��a<��a<��a<��a<��a<Ȭa<٬a<�a<�a<�a<��a<ܬa<�a<ެa<�a<�a<�a<��a<̬a<��a<��a<��a<}�a<`�a<^�a<[�a<.�a<�a<�a<̫a<��a<��a<y�a<S�a< �a<��a<Ȫa<��a<|�a<J�a<�a<�a<��a<��a<h�a<�a<ިa<��a<x�a<C�a<�a<קa<q�a<+�a<�a<��a<f�a<�a<ƥa<a�a<3�a<ۤa<��a<�a<ˣa<^�a<)�a<̢a<d�a<��a<��a<'�a<àa<q�a< �a<��a<'�a<��a<J�a<�a<�a<�a<��a<,�a<��a<Q�a<�a<i�a<��a<��a<,�a<Řa<X�a<��a<]�a<�a<��a<A�a<͕a<h�a<�a<��a<3�a<ϓa<m�a< �a<��a<E�a<�a<��a<Q�a<��a<��a<D�a<��a<ȏa<o�a<%�a<�a<��a<i�a<2�a<��a<��a<��a<f�a<I�a<�a<�a<ʌa<��a<��a<~�a<o�a<m�a<N�a<%�a<,�a<�a<0�a<0�a<7�a<�a<A�a<L�a<_�a<[�a<u�a<��a<�  �  ��a<ӌa<،a<�a<A�a<n�a<��a<��a<
�a<"�a<p�a<��a<�a<3�a<`�a<ʏa<��a<g�a<��a<�a<\�a<��a<�a<]�a<Œa<�a<m�a<�a<>�a<Ŕa<�a<��a<ܕa<_�a<ۖa<3�a<a<	�a<��a< �a<��a<�a<n�a<�a<F�a<�a<T�a<ۜa<I�a<��a<2�a<��a</�a<��a<�a<j�a<ؠa<]�a<��a<G�a<��a<�a<r�a<ԣa<I�a<��a<	�a<9�a<��a<�a<c�a<ʦa<��a<i�a<��a<��a<1�a<��a<ʨa<�a<U�a<z�a<өa<�a<.�a<U�a<�a<Ѫa<�a<1�a<<�a<v�a<��a<��a<�a<�a< �a<�a<H�a<_�a<r�a<��a<��a<��a<��a<ڬa<٬a<߬a<�a<ͬa<�a<�a<��a<��a<�a<�a<ˬa<�a<��a<Ԭa<��a<��a<��a<��a<y�a<Q�a<F�a<�a<�a<��a<٫a<˫a<��a<~�a<;�a<*�a<�a<Ԫa<��a<n�a<d�a<�a<	�a<��a<��a<k�a<�a<�a<��a<��a<-�a<�a<��a<m�a<G�a<�a<��a<C�a<�a<˥a<c�a<.�a<��a<��a<�a<ߣa<w�a<�a<��a<=�a<�a<��a<F�a<נa<k�a<�a<��a<E�a<��a<`�a<�a<t�a<�a<��a<M�a<��a<W�a<�a<y�a<�a<��a<9�a<��a<G�a<ؗa<p�a<�a<��a<<�a<��a<g�a<�a<��a<-�a<��a<t�a<��a<��a<D�a<��a<��a<3�a<�a<��a<i�a<��a<ȏa<j�a<)�a<�a<��a<��a<%�a<�a<΍a<��a<w�a<0�a<$�a<�a<�a<��a<��a<��a<L�a<[�a<>�a<?�a<:�a<%�a<!�a<�a<9�a<�a<I�a<4�a<H�a<j�a<�a<��a<�  �  ��a<Ȍa<�a< �a<9�a<Z�a<��a<ȍa<��a<5�a<g�a<��a<�a<)�a<p�a<��a< �a<M�a<��a<��a<J�a<��a<��a<G�a<��a< �a<��a<ݓa<D�a<��a<�a<��a<��a<]�a<Ζa<P�a<��a<'�a<��a<�a<��a<�a<q�a<�a<v�a<ߛa<B�a<��a<7�a<��a<4�a<��a<�a<��a<��a<j�a<ܠa<M�a<��a<'�a<��a<
�a<h�a<ɣa</�a<��a<��a<c�a<��a<�a<d�a<��a<��a<d�a<��a<�a<E�a<��a<��a<�a<J�a<~�a<��a<��a<*�a<k�a<��a<Ūa<ܪa<�a<@�a<h�a<��a<��a<ͫa<�a<�a<(�a<A�a<^�a<d�a<��a<��a<��a<��a<��a<ìa<Ьa<�a<��a<�a<�a<�a<�a<�a<��a<ڬa<άa<۬a<��a<��a<��a<��a<|�a<n�a<[�a<;�a<>�a<�a<�a<īa<��a<��a<o�a<N�a<!�a<��a<תa<��a<�a<Q�a< �a<�a<��a<��a<Y�a<!�a<�a<��a<w�a<?�a<	�a<��a<s�a<3�a<�a<��a<^�a<
�a<��a<��a<�a<Τa<��a<�a<ȣa<x�a<�a<��a<l�a<��a<��a<,�a<Ơa<i�a<�a<��a<+�a<��a<T�a<�a<x�a<�a<��a<-�a<a<\�a<�a<n�a< �a<��a<+�a<Ƙa<P�a<֗a<q�a<��a<��a<8�a<ŕa<T�a<��a<��a<#�a<˓a<i�a<�a<��a<J�a<�a<��a<M�a<��a<��a<M�a<�a<��a<}�a<-�a<�a<��a<o�a<3�a<��a<͍a<��a<g�a<?�a<�a<��a<Ȍa<��a<��a<��a<|�a<N�a<G�a<;�a<&�a<&�a<2�a<�a<�a<:�a<.�a<?�a<]�a<e�a<t�a<��a<�  �  Ōa<a<�a<�a<U�a<}�a<��a<эa<�a<C�a<k�a<��a<�a<�a<~�a<��a<�a<G�a<��a<��a<;�a<��a<��a<r�a<͒a<�a<z�a<ޓa<X�a<��a<%�a<t�a<�a<d�a<Ėa<P�a<��a<9�a<��a< �a<}�a<��a<��a<�a<a�a<Λa<j�a<ќa<G�a<��a<!�a<��a<�a<��a<��a<n�a<�a<C�a<֡a<�a<��a<��a<i�a<ףa<7�a<��a<�a<M�a<��a<�a<e�a<��a<�a<E�a<��a<ާa<?�a<z�a<��a<�a<1�a<��a<��a<�a<-�a<]�a<��a<ͪa<�a<�a<M�a<^�a<��a<��a<ëa<�a<��a<9�a<7�a<_�a<w�a<��a<��a<��a<¬a<Ŭa<�a<�a<Ѭa<�a<߬a<�a<�a<�a<�a<٬a<�a<¬a<٬a<��a<��a<��a<��a<��a<_�a<n�a<5�a<*�a<��a<	�a<�a<��a<��a<\�a<\�a<%�a<��a<ުa<��a<��a<=�a<4�a<�a<éa<��a<J�a</�a<�a<ɨa<��a<,�a<��a<��a<��a<#�a<��a<��a<Z�a<�a<��a<�a<
�a<ߤa<h�a<2�a<��a<p�a<$�a<��a<X�a<�a<��a<<�a<֠a<j�a<��a<��a<!�a<՞a<P�a<�a<��a<�a<��a<!�a<ϛa<K�a<�a<|�a<�a<��a<"�a<��a<A�a<�a<r�a<��a<��a<�a<ҕa<F�a<��a<��a<$�a<̓a<P�a<�a<��a<Y�a<��a<��a<<�a<��a<��a<L�a<�a<��a<u�a<2�a<܎a<��a<^�a<E�a<�a<΍a<��a<g�a<R�a<�a<��a<ьa<Ča<��a<l�a<j�a<G�a<Y�a<,�a<+�a<*�a<�a<1�a<�a<9�a<!�a<M�a<I�a<_�a<|�a<��a<�  �  ��a<Όa<��a<�a<4�a<]�a<��a<��a< �a<5�a<m�a<��a<�a<*�a<w�a<��a<��a<O�a<��a<��a<N�a<��a<	�a<P�a<��a<�a<��a<ݓa<J�a<��a<�a<��a<�a<i�a<̖a<9�a<��a<*�a<��a<�a<��a<�a<j�a<��a<f�a<�a<H�a<��a<H�a<��a<2�a<��a<�a<��a<��a<r�a<�a<O�a<��a<!�a<��a<�a<j�a<գa<2�a<��a<��a<V�a<��a<�a<i�a<��a<�a<O�a<��a<�a<3�a<{�a<˨a< �a<H�a<��a<��a<��a<'�a<t�a<��a<��a<�a<"�a<@�a<n�a<��a<��a<˫a<�a<�a<3�a<A�a<[�a<i�a<��a<��a<��a<��a<Ԭa<Ĭa<Ӭa<�a<�a<�a<�a<��a<�a<�a<լa<�a<Ԭa<��a<¬a<��a<��a<��a<��a<v�a<R�a<A�a<6�a<�a<�a<ȫa<ëa<��a<u�a<N�a<'�a<��a<Ӫa<��a<��a<P�a<�a<�a<ɩa<��a<]�a<!�a<��a<��a<p�a<:�a<�a<��a<y�a<6�a<�a<��a<Q�a<�a<��a<i�a<�a<Фa<j�a<.�a<ʣa<y�a<�a<Ƣa<]�a<�a<��a<+�a<נa<d�a<�a<��a<%�a<��a<X�a<�a<��a<�a<��a<&�a<Лa<U�a<�a<y�a<�a<��a<-�a<��a<Z�a<՗a<v�a<�a<��a<"�a<��a<W�a<�a<��a</�a<��a<g�a<�a<��a<P�a<�a<��a<G�a<�a<��a<Z�a<�a<��a<s�a<9�a<�a<��a<n�a<?�a<��a<ʍa<��a<h�a<H�a<�a<�a<ߌa<��a<��a<��a<r�a<W�a<9�a<@�a<2�a<0�a<�a<(�a<$�a<�a<6�a<F�a<B�a<n�a<}�a<��a<�  �  ��a<��a<�a<�a<:�a<d�a<��a<��a<�a<�a<p�a<��a<�a<:�a<b�a<Ώa<��a<U�a<��a<�a<d�a<��a<�a<M�a<��a<�a<~�a<�a<8�a<Ŕa<�a<��a<�a<i�a<Җa<4�a<ȗa<�a<��a<	�a<~�a<�a<^�a<�a<R�a<�a<C�a<؜a<?�a<��a<5�a<��a<!�a<}�a<�a<p�a<ߠa<f�a<��a<6�a<��a<�a<l�a<ǣa<I�a<��a<�a<D�a<ƥa<��a<e�a<��a<��a<\�a<��a<�a<2�a<}�a<Шa<��a<M�a<l�a<ɩa<�a<,�a<k�a<��a<ƪa<�a<6�a<-�a<}�a<��a<��a<֫a<�a<'�a<�a<L�a<e�a<h�a<��a<��a<Ĭa<��a<άa<Ѭa<Ӭa<�a<ܬa<�a<֬a<�a<جa<�a<�a<լa<�a<��a<ͬa<��a<��a<��a<i�a<��a<A�a<S�a<!�a<
�a<�a<ϫa<īa<~�a<��a<5�a<*�a<��a<תa<��a<q�a<g�a<�a<��a<��a<�a<s�a<�a<�a<��a<u�a<.�a<��a<��a<g�a<G�a<զa<��a<K�a<�a<��a<d�a<5�a<Ĥa<z�a<�a<£a<��a<��a<Ӣa<I�a<�a<��a<C�a<͠a<d�a<	�a<��a<8�a<��a<h�a<�a<{�a<$�a<��a<<�a<��a<T�a<�a<k�a<�a<��a<3�a<��a<_�a<̗a<s�a<��a<��a<0�a<��a<k�a<�a<��a<4�a<��a<l�a<�a<��a<B�a<�a<��a<8�a<��a<��a<n�a<�a<Ϗa<j�a<*�a<��a<��a<��a<+�a<�a<ԍa<��a<s�a<,�a<3�a<�a<ڌa<��a<��a<{�a<[�a<k�a<,�a<P�a<�a<"�a<"�a<�a<4�a<�a<B�a<=�a<L�a<c�a<a�a<��a<�  �  ��a<ڌa<�a<�a<A�a<x�a<��a<ōa<�a<8�a<{�a<��a<�a<1�a<j�a<��a<�a<E�a<��a<��a<W�a<��a<�a<d�a<Ēa<�a<n�a<�a<A�a<��a< �a<|�a<�a<[�a<Ȗa<G�a<��a<�a<��a<�a<��a< �a<p�a<�a<X�a<ۛa<S�a<ޜa<=�a<��a</�a<��a<�a<��a<�a<o�a<�a<U�a<��a<)�a<��a<�a<u�a<ͣa<G�a<��a<��a<H�a<��a<
�a<`�a<��a<�a<G�a<��a<�a<=�a<|�a<��a<��a<:�a<��a<��a<�a<6�a<U�a<��a<˪a<��a<&�a<;�a<u�a<��a<��a<ƫa<��a<�a<%�a<E�a<g�a<k�a<��a<��a<��a<��a<Ĭa<�a<ݬa<ڬa<ެa<��a<�a<�a<�a<�a<ެa<֬a<Ѭa<Ϭa<��a<��a<��a<��a<�a<p�a<P�a<M�a<�a<�a<��a<�a<��a<��a<z�a<R�a<5�a<��a<ުa<��a<x�a<T�a<-�a<�a<ϩa<��a<e�a<�a<�a<��a<��a<1�a<�a<ça<p�a<5�a<�a<��a<M�a<�a<��a<v�a<�a<��a<k�a<+�a<ɣa<t�a<�a<��a<O�a<��a<��a<I�a<̠a<p�a<�a<��a<0�a<��a<`�a<�a<|�a<�a<��a</�a<̛a<V�a<�a<q�a<�a<��a<,�a<��a<H�a<ܗa<n�a<��a<��a<�a<��a<R�a<��a<��a<%�a<��a<Y�a<�a<��a<E�a<��a<��a<=�a<��a<��a<^�a<��a<Əa<v�a<>�a<��a<��a<q�a<1�a< �a<֍a<��a<y�a<C�a< �a<��a<όa<Ìa<��a<u�a<]�a<_�a<?�a<8�a<(�a<+�a<�a<�a<!�a<.�a<1�a<;�a<H�a<d�a<x�a<��a<�  �  ��a<Ōa<�a<,�a<-�a<i�a<��a<ލa<�a<;�a<g�a<��a<��a<�a<��a<��a<�a<H�a<��a<��a<E�a<��a<��a<^�a<��a<0�a<��a<��a<M�a<��a<'�a<y�a<��a<]�a<��a<L�a<��a<:�a<��a<�a<��a<�a<z�a<�a<}�a<�a<G�a<Ɯa<D�a<a<%�a<��a<�a<��a<��a<p�a<�a<E�a<ҡa<�a<��a<��a<r�a<أa</�a<��a<��a<o�a<��a<�a<\�a<��a<�a<B�a<��a<ݧa<>�a<v�a<��a<�a<7�a<��a<��a<��a<0�a<j�a<��a<��a<�a<�a<U�a<i�a<��a<��a<ƫa<�a<��a<>�a<:�a<f�a<s�a<|�a<��a<��a<ͬa<¬a<Ьa<ͬa<��a<��a<�a<��a<ڬa<��a<�a<جa<�a<��a<Ԭa<��a<��a<��a<��a<��a<W�a<`�a<8�a<=�a<%�a<�a<ԫa<��a<��a<b�a<U�a<!�a<��a<�a<��a<��a<B�a<7�a<�a<ͩa<��a<T�a<9�a<�a<��a<e�a<O�a<�a<��a<|�a<�a<��a<��a<^�a<�a<��a<|�a<�a<�a<c�a<$�a<ǣa<e�a<�a<��a<t�a< �a<��a<0�a<Ӡa<t�a<��a<��a<�a<Оa<Q�a<�a<��a<�a<��a<"�a<ڛa<M�a<�a<}�a< �a<��a<%�a<Ҙa<H�a<�a<i�a<��a<��a<�a<֕a<F�a<��a<��a< �a<ѓa<V�a<�a<��a<M�a<��a<��a<\�a<�a<��a<I�a<�a<��a<m�a<>�a<ߎa<a<^�a<I�a<��a<Սa<��a<a�a<M�a<�a<�a<Όa<��a<��a<��a<~�a<J�a<L�a<#�a<7�a<%�a<�a</�a<�a<4�a< �a<H�a<I�a<a�a<��a<|�a<�  �  ��a<Ɍa<ߌa<�a<H�a<}�a<��a<ˍa<��a<1�a<r�a<��a<�a<'�a<��a<��a<�a<f�a<��a<�a<S�a<��a<��a<o�a<��a<�a<o�a<Փa<G�a<��a<�a<}�a<�a<_�a<Ȗa<:�a<��a< �a<��a<�a<��a<��a<o�a<�a<O�a<ޛa<Z�a<Ԝa<?�a<��a<.�a<��a<!�a<��a<��a<z�a<�a<P�a<ȡa<:�a<��a<�a<n�a<̣a<>�a<��a<��a<B�a<��a<�a<]�a<��a<�a<N�a<��a<�a<1�a<v�a<��a<��a<?�a<~�a<��a<��a<!�a<W�a<��a<ƪa<�a<�a<B�a<s�a<��a<��a<�a<��a<	�a<>�a<C�a<\�a<{�a<��a<��a<��a<��a<Ĭa<�a<�a<�a<լa<�a<�a<�a<�a<�a<۬a<׬a<Ьa<Ȭa<��a<��a<��a<��a<��a<i�a<W�a<<�a<�a<�a<��a<�a<��a<��a<q�a<J�a<+�a<�a<תa<��a<��a<O�a<#�a<�a<©a<��a<b�a<&�a<�a<ƨa<|�a<+�a<�a<��a<v�a<0�a<�a<��a<H�a<�a<��a<i�a<�a<Ƥa<p�a<�a<ңa<n�a<�a<��a<F�a<��a<��a<?�a<Πa<j�a<�a<��a<8�a<̞a<T�a<��a<��a<�a<��a<@�a<��a<T�a<�a<q�a<�a<��a<*�a<��a<E�a<ԗa<k�a<�a<��a<!�a<��a<R�a<�a<��a<#�a<��a<^�a<�a<��a<K�a<�a<��a<6�a<��a<��a<T�a<�a<ďa<s�a<*�a< �a<��a<j�a<J�a<��a<ˍa<��a<t�a<A�a<�a<�a<όa<Ōa<��a<}�a<U�a<P�a<A�a<3�a<3�a<!�a<�a<�a< �a<(�a</�a<>�a<E�a<\�a<z�a<��a<�  �  ��a<�a<�a<�a<>�a<T�a<��a<Ía<�a<9�a<z�a<��a<�a<A�a<c�a<яa<�a<X�a<��a<�a<U�a<��a<�a<>�a<ɒa<�a<��a<�a<?�a<��a<�a<��a<�a<b�a<̖a<-�a<��a<�a<��a<�a<�a<�a<m�a<�a<`�a<�a<=�a<��a<B�a<��a<D�a<��a<*�a<r�a<
�a<v�a<�a<b�a<��a<@�a<��a<�a<l�a<Уa<1�a<}�a<	�a<R�a<ƥa<�a<g�a<��a<��a<p�a<��a<��a<*�a<w�a<Ȩa<��a<W�a<n�a<��a<��a<6�a<o�a<��a<ժa<Ӫa<!�a<>�a<r�a<��a<��a<�a<ګa<"�a<�a<U�a<[�a<b�a<��a<��a<��a<��a<ʬa<��a<Ӭa<�a<�a<�a<ݬa<��a<۬a<�a<�a<Ѭa<�a<��a<Ȭa<��a<��a<��a<o�a<z�a<F�a<W�a<,�a<�a<�a<��a<��a<��a<��a<R�a<3�a<��a<Ϫa<��a<r�a<j�a<�a<��a<��a<��a<c�a<�a<�a<��a<��a<<�a<�a<ʧa<m�a<7�a<֦a<��a<R�a<�a<��a<]�a<-�a<��a<��a<�a<ãa<y�a<�a<΢a<W�a<	�a<��a<+�a<Ѡa<c�a<�a<��a<A�a<��a<c�a<�a<|�a< �a<��a<F�a<��a<k�a<�a<t�a<�a<}�a<9�a<��a<_�a<ڗa<t�a< �a<��a<C�a<��a<c�a<�a<��a<+�a<��a<v�a<�a<��a<J�a<��a<��a<H�a<�a<��a<Y�a<�a<Ïa<��a<"�a<��a<��a<��a<*�a<�a<ʍa<��a<�a<C�a</�a<�a<֌a<��a<��a<��a<j�a<k�a<3�a<F�a<�a< �a<2�a<�a<2�a<�a<<�a<:�a<W�a<a�a<g�a<��a<�  �  ��a<��a<�a<�a<E�a<o�a<��a<͍a<�a<1�a<h�a<��a<��a<:�a<a�a<яa<�a<c�a<��a<��a<;�a<��a<�a<d�a<��a<�a<q�a<ؓa<E�a<��a<�a<}�a<�a<N�a<˖a<<�a<��a<�a<��a<�a<��a<�a<k�a<ݚa<_�a<ޛa<`�a<֜a<_�a<��a<.�a<��a<'�a<��a<�a<m�a<٠a<b�a<͡a<C�a<��a<�a<]�a<�a<D�a<��a<��a<P�a<��a<��a<j�a<��a<��a<N�a<��a<�a<7�a<|�a<��a< �a<<�a<��a<��a<��a<�a<T�a<��a<ƪa<��a<2�a<V�a<Y�a<��a<��a<�a<�a<'�a<�a<Q�a<j�a<��a<��a<��a<��a<��a<�a<٬a<�a<�a<�a<ݬa<�a<��a<�a<ެa<۬a<Ϭa<ɬa<ìa<��a<��a<��a<��a<��a<v�a<Q�a<2�a<!�a<�a<��a<ګa<Ыa<��a<h�a<J�a<!�a<�a<�a<��a<p�a<j�a<5�a<�a<��a<��a<I�a<1�a<�a<��a<y�a<8�a<�a<��a<s�a<3�a<�a<��a<R�a<��a<��a<k�a<�a<��a<p�a<�a<ģa<{�a<�a<��a<V�a<��a<��a<A�a<�a<a�a<�a<��a<=�a<Ϟa<f�a<�a<u�a< �a<��a<I�a<��a<W�a<ךa<��a<�a<��a<+�a<��a<:�a<Ηa<x�a<��a<��a<"�a<��a<L�a<�a<��a<�a<��a<[�a<�a<��a<Q�a<�a<��a<C�a<��a<��a<i�a<�a<��a<w�a<$�a<�a<��a<��a<(�a<�a<ٍa<��a<l�a<?�a<�a<�a<��a<��a<��a<~�a<c�a<E�a<=�a<B�a<,�a<�a<�a<�a<�a<#�a<)�a<0�a<H�a<Z�a<|�a<��a<�  �  ��a<ӌa<�a<�a<?�a<e�a<�a<ƍa<�a<Q�a<_�a<��a<׎a< �a<z�a<��a< �a<V�a<��a<�a<V�a<��a<ڑa<j�a<��a<�a<��a<�a<E�a<��a<)�a<t�a<��a<U�a<͖a<C�a<��a<:�a<��a<�a<z�a<�a<x�a<�a<y�a<ϛa<b�a<��a<5�a<��a<@�a<��a<
�a<��a<�a<|�a<�a<>�a<¡a<!�a<��a<�a<g�a<ʣa<�a<��a<�a<i�a<��a<
�a<N�a<��a<�a<I�a<��a<֧a<8�a<|�a<��a<�a<3�a<��a<��a<��a<*�a<m�a<��a<��a<�a<��a<E�a<p�a<��a<��a<ѫa<�a<�a<4�a<A�a<F�a<��a<t�a<��a<��a<��a<��a<��a<߬a<٬a<��a<�a<��a<ʬa<�a<�a<ެa<�a<��a<ڬa<��a<��a<��a<��a<��a<I�a<d�a<F�a<:�a<�a<�a<Ыa<��a<��a<��a<k�a<�a<�a<Īa<��a<��a<I�a<�a<��a<��a<��a<d�a<$�a<Ǩa<¨a<g�a<=�a<	�a<��a<t�a<�a<��a<��a<e�a<�a<��a<s�a<�a<�a<n�a<,�a<��a<Z�a<�a<��a<p�a<�a<��a<�a<Ġa<j�a<�a<��a<!�a<Ȟa<B�a<��a<��a<��a<��a<'�a<ƛa<j�a<�a<o�a<ޙa<��a<�a<̘a<V�a<ۗa<[�a<�a<��a<�a<ٕa<>�a<�a<��a<�a<ړa<R�a<�a<��a<K�a<�a<��a<O�a<�a<��a<-�a<�a<a<��a<'�a<�a<��a<f�a<?�a<��a<��a<��a<Z�a<]�a<*�a<�a<��a<��a<��a<t�a<{�a<Y�a<N�a<�a<.�a<+�a<�a<+�a<�a<:�a<)�a<D�a<O�a<`�a<��a<n�a<�  �  ��a<��a<�a<�a<E�a<o�a<��a<͍a<�a<1�a<h�a<��a<��a<:�a<a�a<яa<�a<c�a<��a<��a<;�a<��a<�a<d�a<��a<�a<q�a<ؓa<E�a<��a<�a<}�a<�a<N�a<˖a<<�a<��a<�a<��a<�a<��a<�a<k�a<ݚa<_�a<ޛa<`�a<֜a<_�a<��a<.�a<��a<'�a<��a<�a<m�a<٠a<b�a<͡a<C�a<��a<�a<]�a<�a<D�a<��a<��a<P�a<��a<��a<j�a<��a<��a<N�a<��a<�a<7�a<|�a<��a< �a<<�a<��a<��a<��a<�a<T�a<��a<ƪa<��a<2�a<V�a<Y�a<��a<��a<�a<�a<'�a<�a<Q�a<j�a<��a<��a<��a<��a<��a<�a<٬a<�a<�a<�a<ݬa<�a<��a<�a<ެa<۬a<Ϭa<ɬa<ìa<��a<��a<��a<��a<��a<v�a<Q�a<2�a<!�a<�a<��a<ګa<Ыa<��a<h�a<J�a<!�a<�a<�a<��a<p�a<j�a<5�a<�a<��a<��a<I�a<1�a<�a<��a<y�a<8�a<�a<��a<s�a<3�a<�a<��a<R�a<��a<��a<k�a<�a<��a<p�a<�a<ģa<{�a<�a<��a<V�a<��a<��a<A�a<�a<a�a<�a<��a<=�a<Ϟa<f�a<�a<u�a< �a<��a<I�a<��a<W�a<ךa<��a<�a<��a<+�a<��a<:�a<Ηa<x�a<��a<��a<"�a<��a<L�a<�a<��a<�a<��a<[�a<�a<��a<Q�a<�a<��a<C�a<��a<��a<i�a<�a<��a<w�a<$�a<�a<��a<��a<(�a<�a<ٍa<��a<l�a<?�a<�a<�a<��a<��a<��a<~�a<c�a<E�a<=�a<B�a<,�a<�a<�a<�a<�a<#�a<)�a<0�a<H�a<Z�a<|�a<��a<�  �  ��a<�a<�a<�a<>�a<T�a<��a<Ía<�a<9�a<z�a<��a<�a<A�a<c�a<яa<�a<X�a<��a<�a<U�a<��a<�a<>�a<ɒa<�a<��a<�a<?�a<��a<�a<��a<�a<b�a<̖a<-�a<��a<�a<��a<�a<�a<�a<m�a<�a<`�a<�a<=�a<��a<B�a<��a<D�a<��a<*�a<r�a<
�a<v�a<�a<b�a<��a<@�a<��a<�a<l�a<Уa<1�a<}�a<	�a<R�a<ƥa<�a<g�a<��a<��a<p�a<��a<��a<*�a<w�a<Ȩa<��a<W�a<n�a<��a<��a<6�a<o�a<��a<ժa<Ӫa<!�a<>�a<r�a<��a<��a<�a<ګa<"�a<�a<U�a<[�a<b�a<��a<��a<��a<��a<ʬa<��a<Ӭa<�a<�a<�a<ݬa<��a<۬a<�a<�a<Ѭa<�a<��a<Ȭa<��a<��a<��a<o�a<z�a<F�a<W�a<,�a<�a<�a<��a<��a<��a<��a<R�a<3�a<��a<Ϫa<��a<r�a<j�a<�a<��a<��a<��a<c�a<�a<�a<��a<��a<<�a<�a<ʧa<m�a<7�a<֦a<��a<R�a<�a<��a<]�a<-�a<��a<��a<�a<ãa<y�a<�a<΢a<W�a<	�a<��a<+�a<Ѡa<c�a<�a<��a<A�a<��a<c�a<�a<|�a< �a<��a<F�a<��a<k�a<�a<t�a<�a<}�a<9�a<��a<_�a<ڗa<t�a< �a<��a<C�a<��a<c�a<�a<��a<+�a<��a<v�a<�a<��a<J�a<��a<��a<H�a<�a<��a<Y�a<�a<Ïa<��a<"�a<��a<��a<��a<*�a<�a<ʍa<��a<�a<C�a</�a<�a<֌a<��a<��a<��a<j�a<k�a<3�a<F�a<�a< �a<2�a<�a<2�a<�a<<�a<:�a<W�a<a�a<g�a<��a<�  �  ��a<Ɍa<ߌa<�a<H�a<}�a<��a<ˍa<��a<1�a<r�a<��a<�a<'�a<��a<��a<�a<f�a<��a<�a<S�a<��a<��a<o�a<��a<�a<o�a<Փa<G�a<��a<�a<}�a<�a<_�a<Ȗa<:�a<��a< �a<��a<�a<��a<��a<o�a<�a<O�a<ޛa<Z�a<Ԝa<?�a<��a<.�a<��a<!�a<��a<��a<z�a<�a<P�a<ȡa<:�a<��a<�a<n�a<̣a<>�a<��a<��a<B�a<��a<�a<]�a<��a<�a<N�a<��a<�a<1�a<v�a<��a<��a<?�a<~�a<��a<��a<!�a<W�a<��a<ƪa<�a<�a<B�a<s�a<��a<��a<�a<��a<	�a<>�a<C�a<\�a<{�a<��a<��a<��a<��a<Ĭa<�a<�a<�a<լa<�a<�a<�a<�a<�a<۬a<׬a<Ьa<Ȭa<��a<��a<��a<��a<��a<i�a<W�a<<�a<�a<�a<��a<�a<��a<��a<q�a<J�a<+�a<�a<תa<��a<��a<O�a<#�a<�a<©a<��a<b�a<&�a<�a<ƨa<|�a<+�a<�a<��a<v�a<0�a<�a<��a<H�a<�a<��a<i�a<�a<Ƥa<p�a<�a<ңa<n�a<�a<��a<F�a<��a<��a<?�a<Πa<j�a<�a<��a<8�a<̞a<T�a<��a<��a<�a<��a<@�a<��a<T�a<�a<q�a<�a<��a<*�a<��a<E�a<ԗa<k�a<�a<��a<!�a<��a<R�a<�a<��a<#�a<��a<^�a<�a<��a<K�a<�a<��a<6�a<��a<��a<T�a<�a<ďa<s�a<*�a< �a<��a<j�a<J�a<��a<ˍa<��a<t�a<A�a<�a<�a<όa<Ōa<��a<}�a<U�a<P�a<A�a<3�a<3�a<!�a<�a<�a< �a<(�a</�a<>�a<E�a<\�a<z�a<��a<�  �  ��a<Ōa<�a<,�a<-�a<i�a<��a<ލa<�a<;�a<g�a<��a<��a<�a<��a<��a<�a<H�a<��a<��a<E�a<��a<��a<^�a<��a<0�a<��a<��a<M�a<��a<'�a<y�a<��a<]�a<��a<L�a<��a<:�a<��a<�a<��a<�a<z�a<�a<}�a<�a<G�a<Ɯa<D�a<a<%�a<��a<�a<��a<��a<p�a<�a<E�a<ҡa<�a<��a<��a<r�a<أa</�a<��a<��a<o�a<��a<�a<\�a<��a<�a<B�a<��a<ݧa<>�a<v�a<��a<�a<7�a<��a<��a<��a<0�a<j�a<��a<��a<�a<�a<U�a<i�a<��a<��a<ƫa<�a<��a<>�a<:�a<f�a<s�a<|�a<��a<��a<ͬa<¬a<Ьa<ͬa<��a<��a<�a<��a<ڬa<��a<�a<جa<�a<��a<Ԭa<��a<��a<��a<��a<��a<W�a<`�a<8�a<=�a<%�a<�a<ԫa<��a<��a<b�a<U�a<!�a<��a<�a<��a<��a<B�a<7�a<�a<ͩa<��a<T�a<9�a<�a<��a<e�a<O�a<�a<��a<|�a<�a<��a<��a<^�a<�a<��a<|�a<�a<�a<c�a<$�a<ǣa<e�a<�a<��a<t�a< �a<��a<0�a<Ӡa<t�a<��a<��a<�a<Оa<Q�a<�a<��a<�a<��a<"�a<ڛa<M�a<�a<}�a< �a<��a<%�a<Ҙa<H�a<�a<i�a<��a<��a<�a<֕a<F�a<��a<��a< �a<ѓa<V�a<�a<��a<M�a<��a<��a<\�a<�a<��a<I�a<�a<��a<m�a<>�a<ߎa<a<^�a<I�a<��a<Սa<��a<a�a<M�a<�a<�a<Όa<��a<��a<��a<~�a<J�a<L�a<#�a<7�a<%�a<�a</�a<�a<4�a< �a<H�a<I�a<a�a<��a<|�a<�  �  ��a<ڌa<�a<�a<A�a<x�a<��a<ōa<�a<8�a<{�a<��a<�a<1�a<j�a<��a<�a<E�a<��a<��a<W�a<��a<�a<d�a<Ēa<�a<n�a<�a<A�a<��a< �a<|�a<�a<[�a<Ȗa<G�a<��a<�a<��a<�a<��a< �a<p�a<�a<X�a<ۛa<S�a<ޜa<=�a<��a</�a<��a<�a<��a<�a<o�a<�a<U�a<��a<)�a<��a<�a<u�a<ͣa<G�a<��a<��a<H�a<��a<
�a<`�a<��a<�a<G�a<��a<�a<=�a<|�a<��a<��a<:�a<��a<��a<�a<6�a<U�a<��a<˪a<��a<&�a<;�a<u�a<��a<��a<ƫa<��a<�a<%�a<E�a<g�a<k�a<��a<��a<��a<��a<Ĭa<�a<ݬa<ڬa<ެa<��a<�a<�a<�a<�a<ެa<֬a<Ѭa<Ϭa<��a<��a<��a<��a<�a<p�a<P�a<M�a<�a<�a<��a<�a<��a<��a<z�a<R�a<5�a<��a<ުa<��a<x�a<T�a<-�a<�a<ϩa<��a<e�a<�a<�a<��a<��a<1�a<�a<ça<p�a<5�a<�a<��a<M�a<�a<��a<v�a<�a<��a<k�a<+�a<ɣa<t�a<�a<��a<O�a<��a<��a<I�a<̠a<p�a<�a<��a<0�a<��a<`�a<�a<|�a<�a<��a</�a<̛a<V�a<�a<q�a<�a<��a<,�a<��a<H�a<ܗa<n�a<��a<��a<�a<��a<R�a<��a<��a<%�a<��a<Y�a<�a<��a<E�a<��a<��a<=�a<��a<��a<^�a<��a<Əa<v�a<>�a<��a<��a<q�a<1�a< �a<֍a<��a<y�a<C�a< �a<��a<όa<Ìa<��a<u�a<]�a<_�a<?�a<8�a<(�a<+�a<�a<�a<!�a<.�a<1�a<;�a<H�a<d�a<x�a<��a<�  �  ��a<��a<�a<�a<:�a<d�a<��a<��a<�a<�a<p�a<��a<�a<:�a<b�a<Ώa<��a<U�a<��a<�a<d�a<��a<�a<M�a<��a<�a<~�a<�a<8�a<Ŕa<�a<��a<�a<i�a<Җa<4�a<ȗa<�a<��a<	�a<~�a<�a<^�a<�a<R�a<�a<C�a<؜a<?�a<��a<5�a<��a<!�a<}�a<�a<p�a<ߠa<f�a<��a<6�a<��a<�a<l�a<ǣa<I�a<��a<�a<D�a<ƥa<��a<e�a<��a<��a<\�a<��a<�a<2�a<}�a<Шa<��a<M�a<l�a<ɩa<�a<,�a<k�a<��a<ƪa<�a<6�a<-�a<}�a<��a<��a<֫a<�a<'�a<�a<L�a<e�a<h�a<��a<��a<Ĭa<��a<άa<Ѭa<Ӭa<�a<ܬa<�a<֬a<�a<جa<�a<�a<լa<�a<��a<ͬa<��a<��a<��a<i�a<��a<A�a<S�a<!�a<
�a<�a<ϫa<īa<~�a<��a<5�a<*�a<��a<תa<��a<q�a<g�a<�a<��a<��a<�a<s�a<�a<�a<��a<u�a<.�a<��a<��a<g�a<G�a<զa<��a<K�a<�a<��a<d�a<5�a<Ĥa<z�a<�a<£a<��a<��a<Ӣa<I�a<�a<��a<C�a<͠a<d�a<	�a<��a<8�a<��a<h�a<�a<{�a<$�a<��a<<�a<��a<T�a<�a<k�a<�a<��a<3�a<��a<_�a<̗a<s�a<��a<��a<0�a<��a<k�a<�a<��a<4�a<��a<l�a<�a<��a<B�a<�a<��a<8�a<��a<��a<n�a<�a<Ϗa<j�a<*�a<��a<��a<��a<+�a<�a<ԍa<��a<s�a<,�a<3�a<�a<ڌa<��a<��a<{�a<[�a<k�a<,�a<P�a<�a<"�a<"�a<�a<4�a<�a<B�a<=�a<L�a<c�a<a�a<��a<�  �  ��a<Όa<��a<�a<4�a<]�a<��a<��a< �a<5�a<m�a<��a<�a<*�a<w�a<��a<��a<O�a<��a<��a<N�a<��a<	�a<P�a<��a<�a<��a<ݓa<J�a<��a<�a<��a<�a<i�a<̖a<9�a<��a<*�a<��a<�a<��a<�a<j�a<��a<f�a<�a<H�a<��a<H�a<��a<2�a<��a<�a<��a<��a<r�a<�a<O�a<��a<!�a<��a<�a<j�a<գa<2�a<��a<��a<V�a<��a<�a<i�a<��a<�a<O�a<��a<�a<3�a<{�a<˨a< �a<H�a<��a<��a<��a<'�a<t�a<��a<��a<�a<"�a<@�a<n�a<��a<��a<˫a<�a<�a<3�a<A�a<[�a<i�a<��a<��a<��a<��a<Ԭa<Ĭa<Ӭa<�a<�a<�a<�a<��a<�a<�a<լa<�a<Ԭa<��a<¬a<��a<��a<��a<��a<v�a<R�a<A�a<6�a<�a<�a<ȫa<ëa<��a<u�a<N�a<'�a<��a<Ӫa<��a<��a<P�a<�a<�a<ɩa<��a<]�a<!�a<��a<��a<p�a<:�a<�a<��a<y�a<6�a<�a<��a<Q�a<�a<��a<i�a<�a<Фa<j�a<.�a<ʣa<y�a<�a<Ƣa<]�a<�a<��a<+�a<נa<d�a<�a<��a<%�a<��a<X�a<�a<��a<�a<��a<&�a<Лa<U�a<�a<y�a<�a<��a<-�a<��a<Z�a<՗a<v�a<�a<��a<"�a<��a<W�a<�a<��a</�a<��a<g�a<�a<��a<P�a<�a<��a<G�a<�a<��a<Z�a<�a<��a<s�a<9�a<�a<��a<n�a<?�a<��a<ʍa<��a<h�a<H�a<�a<�a<ߌa<��a<��a<��a<r�a<W�a<9�a<@�a<2�a<0�a<�a<(�a<$�a<�a<6�a<F�a<B�a<n�a<}�a<��a<�  �  Ōa<a<�a<�a<U�a<}�a<��a<эa<�a<C�a<k�a<��a<�a<�a<~�a<��a<�a<G�a<��a<��a<;�a<��a<��a<r�a<͒a<�a<z�a<ޓa<X�a<��a<%�a<t�a<�a<d�a<Ėa<P�a<��a<9�a<��a< �a<}�a<��a<��a<�a<a�a<Λa<j�a<ќa<G�a<��a<!�a<��a<�a<��a<��a<n�a<�a<C�a<֡a<�a<��a<��a<i�a<ףa<7�a<��a<�a<M�a<��a<�a<e�a<��a<�a<E�a<��a<ާa<?�a<z�a<��a<�a<1�a<��a<��a<�a<-�a<]�a<��a<ͪa<�a<�a<M�a<^�a<��a<��a<ëa<�a<��a<9�a<7�a<_�a<w�a<��a<��a<��a<¬a<Ŭa<�a<�a<Ѭa<�a<߬a<�a<�a<�a<�a<٬a<�a<¬a<٬a<��a<��a<��a<��a<��a<_�a<n�a<5�a<*�a<��a<	�a<�a<��a<��a<\�a<\�a<%�a<��a<ުa<��a<��a<=�a<4�a<�a<éa<��a<J�a</�a<�a<ɨa<��a<,�a<��a<��a<��a<#�a<��a<��a<Z�a<�a<��a<�a<
�a<ߤa<h�a<2�a<��a<p�a<$�a<��a<X�a<�a<��a<<�a<֠a<j�a<��a<��a<!�a<՞a<P�a<�a<��a<�a<��a<!�a<ϛa<K�a<�a<|�a<�a<��a<"�a<��a<A�a<�a<r�a<��a<��a<�a<ҕa<F�a<��a<��a<$�a<̓a<P�a<�a<��a<Y�a<��a<��a<<�a<��a<��a<L�a<�a<��a<u�a<2�a<܎a<��a<^�a<E�a<�a<΍a<��a<g�a<R�a<�a<��a<ьa<Ča<��a<l�a<j�a<G�a<Y�a<,�a<+�a<*�a<�a<1�a<�a<9�a<!�a<M�a<I�a<_�a<|�a<��a<�  �  ��a<Ȍa<�a< �a<9�a<Z�a<��a<ȍa<��a<5�a<g�a<��a<�a<)�a<p�a<��a< �a<M�a<��a<��a<J�a<��a<��a<G�a<��a< �a<��a<ݓa<D�a<��a<�a<��a<��a<]�a<Ζa<P�a<��a<'�a<��a<�a<��a<�a<q�a<�a<v�a<ߛa<B�a<��a<7�a<��a<4�a<��a<�a<��a<��a<j�a<ܠa<M�a<��a<'�a<��a<
�a<h�a<ɣa</�a<��a<��a<c�a<��a<�a<d�a<��a<��a<d�a<��a<�a<E�a<��a<��a<�a<J�a<~�a<��a<��a<*�a<k�a<��a<Ūa<ܪa<�a<@�a<h�a<��a<��a<ͫa<�a<�a<(�a<A�a<^�a<d�a<��a<��a<��a<��a<��a<ìa<Ьa<�a<��a<�a<�a<�a<�a<�a<��a<ڬa<άa<۬a<��a<��a<��a<��a<|�a<n�a<[�a<;�a<>�a<�a<�a<īa<��a<��a<o�a<N�a<!�a<��a<תa<��a<�a<Q�a< �a<�a<��a<��a<Y�a<!�a<�a<��a<w�a<?�a<	�a<��a<s�a<3�a<�a<��a<^�a<
�a<��a<��a<�a<Τa<��a<�a<ȣa<x�a<�a<��a<l�a<��a<��a<,�a<Ơa<i�a<�a<��a<+�a<��a<T�a<�a<x�a<�a<��a<-�a<a<\�a<�a<n�a< �a<��a<+�a<Ƙa<P�a<֗a<q�a<��a<��a<8�a<ŕa<T�a<��a<��a<#�a<˓a<i�a<�a<��a<J�a<�a<��a<M�a<��a<��a<M�a<�a<��a<}�a<-�a<�a<��a<o�a<3�a<��a<͍a<��a<g�a<?�a<�a<��a<Ȍa<��a<��a<��a<|�a<N�a<G�a<;�a<&�a<&�a<2�a<�a<�a<:�a<.�a<?�a<]�a<e�a<t�a<��a<�  �  ��a<ӌa<،a<�a<A�a<n�a<��a<��a<
�a<"�a<p�a<��a<�a<3�a<`�a<ʏa<��a<g�a<��a<�a<\�a<��a<�a<]�a<Œa<�a<m�a<�a<>�a<Ŕa<�a<��a<ܕa<_�a<ۖa<3�a<a<	�a<��a< �a<��a<�a<n�a<�a<F�a<�a<T�a<ۜa<I�a<��a<2�a<��a</�a<��a<�a<j�a<ؠa<]�a<��a<G�a<��a<�a<r�a<ԣa<I�a<��a<	�a<9�a<��a<�a<c�a<ʦa<��a<i�a<��a<��a<1�a<��a<ʨa<�a<U�a<z�a<өa<�a<.�a<U�a<�a<Ѫa<�a<1�a<<�a<v�a<��a<��a<�a<�a< �a<�a<H�a<_�a<r�a<��a<��a<��a<��a<ڬa<٬a<߬a<�a<ͬa<�a<�a<��a<��a<�a<�a<ˬa<�a<��a<Ԭa<��a<��a<��a<��a<y�a<Q�a<F�a<�a<�a<��a<٫a<˫a<��a<~�a<;�a<*�a<�a<Ԫa<��a<n�a<d�a<�a<	�a<��a<��a<k�a<�a<�a<��a<��a<-�a<�a<��a<m�a<G�a<�a<��a<C�a<�a<˥a<c�a<.�a<��a<��a<�a<ߣa<w�a<�a<��a<=�a<�a<��a<F�a<נa<k�a<�a<��a<E�a<��a<`�a<�a<t�a<�a<��a<M�a<��a<W�a<�a<y�a<�a<��a<9�a<��a<G�a<ؗa<p�a<�a<��a<<�a<��a<g�a<�a<��a<-�a<��a<t�a<��a<��a<D�a<��a<��a<3�a<�a<��a<i�a<��a<ȏa<j�a<)�a<�a<��a<��a<%�a<�a<΍a<��a<w�a<0�a<$�a<�a<�a<��a<��a<��a<L�a<[�a<>�a<?�a<:�a<%�a<!�a<�a<9�a<�a<I�a<4�a<H�a<j�a<�a<��a<�  �  ��a<�a<��a<�a<<�a<b�a<��a<Ía<�a<9�a<f�a<��a<ێa<$�a<m�a<��a<��a<L�a<��a<��a<Y�a<��a<�a<W�a<��a<$�a<��a<��a<C�a<��a<�a<��a<��a<j�a<֖a<1�a<Ɨa<5�a<��a<�a<��a<�a<��a<��a<n�a<ߛa<N�a<��a<4�a<��a<,�a<��a<�a<��a<�a<q�a<�a<G�a<��a<'�a<��a<��a<v�a<ţa<&�a<��a<��a<a�a<��a<#�a<P�a<��a<��a<n�a<��a< �a<,�a<|�a<Ϩa<�a<N�a<~�a<��a<�a<J�a<k�a<��a<Ūa<�a<�a<=�a<w�a<��a<��a<Ϋa<�a<�a<'�a<@�a<M�a<n�a<��a<��a<��a<��a<��a<Ȭa<٬a<�a<�a<�a<��a<ܬa<�a<ެa<�a<�a<�a<��a<̬a<��a<��a<��a<}�a<`�a<^�a<[�a<.�a<�a<�a<̫a<��a<��a<y�a<S�a< �a<��a<Ȫa<��a<|�a<J�a<�a<�a<��a<��a<h�a<�a<ިa<��a<x�a<C�a<�a<קa<q�a<+�a<�a<��a<f�a<�a<ƥa<a�a<3�a<ۤa<��a<�a<ˣa<^�a<)�a<̢a<d�a<��a<��a<'�a<àa<q�a< �a<��a<'�a<��a<J�a<�a<�a<�a<��a<,�a<��a<Q�a<�a<i�a<��a<��a<,�a<Řa<X�a<��a<]�a<�a<��a<A�a<͕a<h�a<�a<��a<3�a<ϓa<m�a< �a<��a<E�a<�a<��a<Q�a<��a<��a<D�a<��a<ȏa<o�a<%�a<�a<��a<i�a<2�a<��a<��a<��a<f�a<I�a<�a<�a<ʌa<��a<��a<~�a<o�a<m�a<N�a<%�a<,�a<�a<0�a<0�a<7�a<�a<A�a<L�a<_�a<[�a<u�a<��a<�  �  ��a<Q�a<��a<��a<؍a<%�a<,�a<��a<��a<Ԏa<�a<`�a<��a<��a<2�a<G�a<ǐa<�a<+�a<��a<ۑa<V�a<��a<�a<:�a<˓a<�a<s�a<�a<@�a<ѕa<�a<��a<�a<l�a<��a<7�a<��a<�a<��a<'�a<��a<,�a<F�a<	�a<K�a<�a<X�a<ǝa<G�a<��a<*�a<v�a<.�a<~�a<��a<m�a<ȡa<]�a<��a<�a<n�a<�a<Q�a<��a<&�a<P�a<�a<��a<��a<��a<9�a<��a<��a< �a<[�a<��a<��a<1�a<��a<��a<�a<.�a<��a<��a<��a<#�a<�a<��a<��a<ͫa<ثa<�a<�a<B�a<��a<w�a<��a<��a<ެa<�a<ܬa<�a<�a<L�a<2�a<Z�a<X�a<X�a<u�a<8�a<��a<n�a<|�a<i�a<P�a<X�a<G�a<_�a<:�a<.�a<�a<�a<�a<�a<�a<��a<��a<��a<c�a<h�a<"�a<'�a<׫a<ƫa<��a<��a<h�a<�a<�a<��a<ªa<o�a<'�a<�a<ǩa<��a<X�a<M�a<רa<ʨa<b�a<+�a<"�a<��a<��a<
�a<Ԧa<�a<B�a<��a<��a<L�a<٤a<��a<X�a<�a<��a<�a<�a<^�a<&�a<��a<N�a<�a<m�a<�a<��a<g�a<ٞa<u�a<�a<��a<G�a<��a<N�a<͛a<p�a<�a<��a<8�a<��a<b�a<��a<��a<�a<��a<6�a<��a<Z�a<�a<��a<)�a<��a<b�a<�a<��a<<�a<�a<��a<�a<��a<s�a<`�a<�a<��a<Q�a<�a<��a<��a<r�a<�a<�a<��a<w�a<Z�a<�a<�a<��a<��a<h�a<f�a<>�a<�a<�a<ˌa<!�a<�a<�a<ьa<��a<Ȍa<��a<�a<ٌa<�a<�a<�a<:�a<4�a<�  �  J�a<u�a<��a<��a<�a<�a<0�a<|�a<��a<�a<�a<K�a<��a<Ǐa<�a<T�a<��a<�a<O�a<��a<�a<R�a<��a<��a<J�a<Ǔa<%�a<�a<̔a<1�a<��a<�a<��a<�a<n�a<חa<R�a<��a<4�a<��a<�a<i�a<�a<�a<�a<^�a<�a<M�a<͝a<M�a<��a<<�a<��a<�a<x�a<�a<\�a<ɡa<5�a<��a<(�a<��a<��a<U�a<��a<�a<d�a<�a<1�a<��a<��a<*�a<��a<ԧa<$�a<v�a<��a<��a<J�a<��a<��a<�a<"�a<T�a<��a<�a<�a<+�a<m�a<��a<ͫa<�a<�a<;�a<G�a<d�a<��a<��a<��a<̬a<�a<�a<$�a<-�a<D�a<9�a<H�a<Z�a<^�a<w�a<i�a<a�a<I�a<p�a<h�a<k�a<^�a<W�a<N�a<?�a<5�a<+�a<�a<�a<ˬa<ʬa<��a<��a<��a<n�a<R�a<%�a<�a<��a<ثa<��a<z�a<J�a<!�a<��a<Ȫa<��a<k�a<J�a<�a<۩a<��a<\�a<2�a<�a<ƨa<��a<8�a<ݧa<��a<q�a<�a<�a<��a<D�a<�a<��a<O�a<��a<��a<J�a<̣a<��a<=�a<�a<q�a<�a<��a<T�a<��a<��a</�a<��a<?�a<Ӟa<k�a<��a<��a<�a<��a<_�a<�a<��a<
�a<��a<+�a<��a<Z�a<�a<n�a<ߗa<��a<-�a<Ŗa<^�a<��a<��a<+�a<ϔa<k�a<��a<��a<0�a<Βa<��a<F�a<��a<��a<F�a<�a<��a<d�a<(�a<��a<��a<H�a<�a<ӎa<��a<e�a<?�a<�a<��a<ƍa<��a<o�a<T�a<A�a<$�a<!�a<��a<�a<��a<یa<Ќa<Ԍa<͌a<ьa<،a<ތa<�a<�a<�a<(�a<�a<�  �  K�a<��a<��a<��a<�a<�a<J�a<\�a<��a<a<�a<L�a<��a<�a<��a<��a<��a<��a<E�a<��a<�a<6�a<��a<�a<g�a<��a<�a<��a<ߔa<m�a<��a<�a<��a<�a<d�a<ȗa<V�a<��a<B�a<��a<2�a<��a<�a<��a<؛a<n�a<��a<W�a<ʝa<&�a<��a<�a<��a<�a<��a<�a<Z�a<�a<0�a<��a<�a<w�a<Уa<G�a<��a<�a<}�a<��a<;�a<��a<�a<O�a<s�a<�a<	�a<t�a<��a<�a<<�a<p�a<ĩa<�a<[�a<o�a<��a<۪a<��a<L�a<g�a<��a<��a<ԫa<��a<$�a<S�a<]�a<��a<��a<Ҭa<ݬa<�a<�a<��a<%�a<�a<N�a<N�a<_�a<Y�a<Q�a<��a<`�a<��a<x�a<Y�a<q�a<I�a<X�a<<�a<A�a<%�a<+�a<�a<	�a<�a<ˬa<Ԭa<��a<��a<|�a<Q�a<@�a<��a<�a<��a<��a<{�a<Q�a<D�a<�a<��a<��a<t�a<@�a<��a<̩a<��a<x�a<)�a<�a<��a<p�a<F�a<�a<ҧa<`�a<�a<Цa<��a<:�a<ߥa<��a<4�a<
�a<��a<c�a<��a<��a<N�a<��a<��a<�a<��a<Q�a<Ҡa<~�a<�a<��a<:�a<��a<q�a<��a<��a<�a<Ȝa<:�a<֛a<Y�a<��a<��a<'�a<��a<3�a<�a<o�a<�a<��a<�a<іa<C�a<��a<{�a<�a<��a<Q�a<�a<��a<i�a<�a<��a<;�a<בa<��a<@�a<�a<��a<M�a<
�a<ɏa<��a<A�a<9�a<Ŏa<��a<v�a<9�a<�a<Ѝa<��a<��a<��a<Z�a<E�a<�a<��a<�a<�a<��a<�a<��a<ڌa<��a<ӌa<ƌa<��a<݌a<�a<�a<+�a<U�a<�  �  ]�a<o�a<��a<��a<ߍa<�a<E�a<k�a<��a<ڎa<�a<V�a<|�a<Џa<�a<Y�a<��a< �a<<�a<��a<��a<@�a<��a<�a<[�a<��a<�a<}�a<�a<?�a<��a<$�a<��a<��a<j�a<ڗa<S�a<��a<5�a<��a<�a<��a<�a<s�a<��a<q�a<֜a<T�a<̝a<B�a<Ȟa<�a<��a<�a<z�a<�a<d�a<ʡa<6�a<��a<�a<��a<�a<L�a<��a<�a<y�a<إa<'�a<��a<ڦa<!�a<v�a<֧a<�a<p�a<��a<��a<A�a<��a<ǩa<�a<)�a<s�a<��a<תa<�a<@�a<^�a<��a<��a<�a<�a<$�a<Z�a<_�a<��a<��a<��a<Ǭa<�a<�a<�a<@�a<3�a<H�a<J�a<Q�a<g�a<k�a<b�a<n�a<j�a<X�a<b�a<g�a<\�a<Z�a<K�a<D�a<2�a<#�a<�a<�a<�a<ݬa<��a<��a<��a<k�a<G�a<:�a<�a<�a<ͫa<��a<��a<B�a<+�a<��a<ͪa<��a<}�a<8�a<�a<�a<��a<s�a<"�a<��a<��a<s�a<6�a<��a<��a<W�a<&�a<٦a<��a<@�a<�a<��a<K�a<��a<��a<8�a<�a<��a<1�a<�a<��a<�a<��a<S�a<�a<��a<�a<��a<A�a<՞a<q�a<�a<��a< �a<Ĝa<E�a<�a<w�a<�a<��a<�a<��a<Q�a<טa<q�a<�a<��a< �a<ǖa<X�a<��a<��a<(�a<Ɣa<e�a<�a<��a<7�a<�a<��a<7�a<�a<��a<6�a<��a<��a<k�a<'�a<ɏa<��a<C�a<�a<؎a<��a<`�a<A�a<�a<�a<ٍa<��a<~�a<U�a<7�a<-�a<�a<��a<�a<݌a<Ìa<ʌa<Ќa<ˌa<Ԍa<Ռa<�a<�a<��a<
�a<�a<4�a<�  �  g�a<b�a<��a<��a<�a<�a<:�a<u�a<��a<؎a<�a<V�a<��a<ˏa<#�a<P�a<��a<��a<;�a<��a<�a<O�a<��a<��a<N�a<��a<�a<r�a<�a<<�a<Еa<�a<��a<��a<Y�a<ߗa<=�a<ǘa<�a<��a<�a<��a<�a<o�a<��a<]�a<�a<Q�a<ǝa<B�a<��a<&�a<��a<�a<y�a<��a<o�a<ơa<P�a<��a<�a<q�a<�a<K�a<��a<�a<f�a<ޥa<$�a<��a<֦a<-�a<��a<��a<%�a<_�a<��a<�a<9�a<��a<��a<�a<,�a<w�a<��a<ݪa<�a<1�a<p�a<��a<ƫa<ܫa< �a<*�a<R�a<x�a<{�a<��a<��a<լa<��a<��a<�a<�a<;�a<=�a<O�a<\�a<X�a<q�a<X�a<z�a<Z�a<|�a<x�a<I�a<e�a<G�a<Q�a</�a<7�a<�a<�a<�a<٬a<�a<��a<��a<��a<p�a<T�a</�a<�a<�a<ʫa<��a<��a<T�a<%�a<�a<Īa<��a<w�a<7�a<�a<ͩa<��a<f�a<4�a<�a<��a<|�a<+�a<��a<��a<��a<�a<Ѧa<��a</�a<��a<��a<V�a<ޤa<��a<P�a<�a<��a<-�a<�a<p�a<%�a<��a<N�a<�a<t�a<�a<��a<W�a<Ԟa<v�a<�a<��a<:�a<��a<N�a<Лa<q�a< �a<��a<1�a<��a<W�a<Ԙa<u�a<��a<��a<H�a<��a<_�a<�a<��a<�a<��a<b�a<��a<��a<:�a<�a<��a<=�a<�a<��a<I�a<�a<��a<U�a<�a<Ϗa<��a<\�a<�a<�a<��a<m�a<L�a<�a<�a<��a<��a<s�a<[�a<C�a<�a<�a<�a<��a<Όa<�a<��a<��a<Ԍa<��a<یa<Όa<�a<�a<�a<9�a<(�a<�  �  W�a<z�a<��a<��a<�a<�a<A�a<v�a<��a<ڎa<�a<H�a<��a<ԏa<
�a<j�a<��a<�a<O�a<��a<�a<O�a<��a<��a<^�a<��a<�a<x�a<�a<M�a<��a<�a<��a<�a<b�a<�a<8�a<Ƙa<,�a<��a<�a<��a< �a<��a<�a<f�a<�a<P�a<ҝa<H�a<��a<0�a<��a<
�a<��a<�a<[�a<סa<<�a<��a<#�a<}�a<�a<V�a<��a<�a<u�a<ɥa<,�a<{�a<ܦa<(�a<s�a<Χa<)�a<]�a<��a<��a<5�a<��a<��a<�a<7�a<s�a<��a<ڪa<�a<E�a<h�a<��a<ɫa<�a<�a<9�a<F�a<m�a<��a<��a<��a<�a<�a<�a<�a<#�a<:�a<J�a<F�a<\�a<V�a<b�a<q�a<m�a<i�a<f�a<Y�a<b�a<c�a<H�a<]�a<6�a<4�a<'�a<�a<��a<�a<׬a<ìa<��a<��a<w�a<J�a<7�a<�a<�a<ͫa<��a<v�a<\�a<.�a<�a<ުa<��a<i�a<J�a<�a<ީa<��a<c�a<+�a<��a<��a<{�a<1�a<��a<��a<_�a<�a<ڦa<��a<8�a<��a<��a<V�a<��a<��a<A�a<�a<��a<@�a<Ӣa<y�a<�a<��a<Y�a<��a<��a<#�a<��a<B�a<�a<h�a<��a<��a<&�a<��a<Z�a<ݛa<y�a<�a<��a<)�a<��a<B�a<ܘa<e�a<�a<��a<�a<��a<c�a<�a<��a<%�a<��a<e�a<��a<��a<E�a<�a<��a<:�a<ܑa<��a<@�a<�a<��a<f�a<�a<ޏa<��a<Q�a< �a<юa<��a<y�a<:�a<�a<�a<��a<��a<��a<R�a<C�a<�a<�a<�a<�a<݌a<ьa<��a<ˌa<Ҍa<Ìa<�a<Ռa<�a<��a<��a<�a<9�a<�  �  B�a<}�a<��a<̍a<�a<�a<F�a<[�a<��a<͎a<#�a<^�a<��a<Ώa<�a<^�a<��a<�a<M�a<��a<��a<2�a<��a<�a<l�a<��a<�a<��a<Ӕa<O�a<��a<4�a<��a<�a<g�a<ӗa<B�a<��a<G�a<��a<�a<��a<��a<��a<�a<��a<לa<Y�a<˝a<=�a<��a< �a<��a<�a<�a<��a<c�a<̡a<9�a<Ǣa<�a<��a<�a<I�a<��a<�a<��a<åa<1�a<|�a<�a</�a<}�a<�a<�a<a�a<��a<��a<7�a<z�a<ةa<�a<:�a<g�a<��a<ުa<	�a<T�a<`�a<��a<��a<�a<�a<1�a<h�a<e�a<��a<��a<¬a<Ҭa<��a<�a<	�a<.�a<$�a<J�a<M�a<_�a<q�a<]�a<p�a<W�a<r�a<^�a<n�a<t�a<M�a<Q�a<@�a<9�a<"�a<1�a<�a<�a<�a<¬a<Ǭa<��a<��a<}�a<K�a<;�a<��a<��a<��a<��a<��a<K�a<(�a<��a<Ҫa<��a<��a<H�a<�a<�a<��a<r�a<(�a<�a<��a<y�a<<�a<�a<��a<Y�a<6�a<٦a<��a<>�a<�a<��a<@�a<�a<��a<C�a<��a<��a<@�a<΢a<��a<�a<��a<R�a<�a<��a<�a<Пa<D�a<ڞa<r�a<�a<��a<#�a<לa<J�a<�a<w�a<��a<��a<�a<Йa<<�a<�a<f�a<	�a<��a<'�a<ٖa<N�a<�a<��a<$�a<��a<[�a<�a<��a<H�a<�a<��a<>�a<�a<��a<8�a<��a<��a<j�a<�a<֏a<��a<H�a<�a<؎a<��a<j�a<I�a<(�a<ۍa<Ǎa<��a<��a<Y�a<E�a<6�a<�a<�a<،a<�a<Ɍa<Ռa<݌a<��a<̌a<ˌa<،a<یa<�a<�a<�a<B�a<�  �  _�a<v�a<��a<Ía<ߍa<�a<@�a<q�a<��a<Ԏa<�a<W�a<��a<̏a<+�a<R�a<��a<��a<:�a<��a<�a<G�a<��a<��a<P�a<��a<�a<��a<�a<D�a<��a<�a<��a<��a<a�a<˗a<O�a<��a<$�a<��a<�a<��a<�a<v�a<�a<p�a<Ԝa<S�a<a<F�a<��a< �a<��a<�a<~�a<��a<o�a<ˡa<N�a<��a<�a<{�a<�a<E�a<��a<�a<w�a<ѥa<*�a<��a<�a<(�a<��a<ǧa<�a<l�a<��a<�a<@�a<u�a<��a<��a<2�a<u�a<��a<Ӫa<�a<8�a<b�a<��a<��a<�a<�a<"�a<N�a<{�a<{�a<��a<��a<֬a<��a<��a<�a<+�a<9�a<A�a<T�a<S�a<e�a<_�a<c�a<u�a<o�a<i�a<m�a<V�a<Y�a<[�a<;�a<@�a<2�a<�a<�a<��a<�a<߬a<��a<��a<��a<k�a<V�a<6�a<�a<�a<ƫa<��a<��a<X�a<&�a<�a<ƪa<��a<s�a<5�a<
�a<٩a<��a<t�a<*�a<�a<��a<n�a<>�a<��a<��a<h�a< �a<Φa<��a<8�a<�a<��a<H�a<�a<��a<A�a<��a<��a<4�a<آa<��a<�a<��a<I�a<�a<��a<�a<��a<S�a<ٞa<w�a<�a<��a<8�a<��a<C�a<ۛa<u�a<��a<��a<�a<��a<J�a<ژa<v�a<�a<��a<5�a<��a<S�a<��a<�a<�a<Ŕa<W�a<��a<��a<@�a<�a<��a<3�a<�a<��a<;�a<��a<��a<a�a<�a<Ǐa<��a<_�a<�a<�a<��a<o�a<F�a<	�a<�a<ča<��a<w�a<_�a<9�a<+�a<	�a<��a<��a<�a<Ԍa<Ԍa<��a<Ȍa<Ռa<Ōa<ߌa<�a<�a<�a<!�a<<�a<�  �  ]�a<q�a<��a<��a<��a<�a<,�a<��a<��a<�a<�a<C�a<��a<Ïa< �a<T�a<��a<ܐa<^�a<��a<ߑa<R�a<��a<�a<Q�a<��a<�a<w�a<�a<<�a<��a<�a<��a<�a<c�a<�a<6�a<Ƙa</�a<��a<�a<��a<	�a<w�a<��a<\�a<�a<W�a<ʝa<G�a<��a<G�a<��a<�a<��a<�a<f�a<͡a<H�a<��a<6�a<~�a<�a<R�a<��a<!�a<f�a<ڥa<(�a<��a<צa<�a<�a<ͧa<+�a<X�a<��a<��a<2�a<��a<��a<��a<&�a<r�a<��a<תa<�a<3�a<w�a<��a<ʫa<ݫa<�a<K�a<6�a<}�a<��a<��a<��a<ެa<�a<�a<3�a<�a<C�a<6�a<V�a<W�a<W�a<g�a<e�a<t�a<^�a<c�a<X�a<e�a<^�a<D�a<U�a<3�a</�a<&�a<�a<��a<ެa<ݬa<��a<��a<��a<l�a<]�a<!�a<$�a<߫a<�a<��a<r�a<]�a<�a<
�a<Ȫa<��a<Z�a<Y�a<�a<ʩa<��a<Y�a<<�a<�a<��a<w�a<0�a<��a<��a<e�a<�a<�a<��a<9�a<��a<��a<V�a<��a<��a<<�a<�a<��a<5�a<�a<o�a<"�a<��a<Q�a<�a<}�a<9�a<��a<N�a<۞a<o�a<�a<��a<2�a<��a<m�a<ݛa<r�a<�a<��a<3�a<��a<S�a<ؘa<l�a<��a<��a<)�a<��a<e�a<ߕa<��a<$�a<��a<k�a<��a<��a<4�a<�a<��a<7�a<�a<��a<O�a<�a<��a<V�a<#�a<�a<x�a<`�a<�a<�a<��a<w�a<:�a<�a<�a<��a<��a<l�a<a�a<=�a<�a<�a<��a<��a<ьa<Όa<��a<Όa<͌a<��a<��a<Ҍa<�a<��a<��a<�a<,�a<�  �  R�a<|�a<��a<��a<�a<�a<:�a<v�a<��a<Ύa<�a<Q�a<��a<؏a<�a<g�a<��a<��a<A�a<��a<�a<H�a<��a< �a<`�a<��a<�a<��a<��a<b�a<��a<�a<��a<�a<e�a<ӗa<=�a<��a<8�a<��a<'�a<��a<�a<�a<�a<m�a<�a<S�a<͝a<D�a<��a<�a<��a<�a<��a<��a<g�a<ۡa<C�a<��a<�a<u�a<�a<Q�a<��a<�a<y�a<ĥa<,�a<��a<�a<=�a<v�a<קa<�a<]�a<��a<��a<0�a<u�a<©a<�a<J�a<p�a<��a<٪a<�a<F�a<p�a<��a<«a<�a<��a<(�a<W�a<q�a<��a<��a<Ƭa<�a<�a<
�a<�a<�a<<�a<B�a<L�a<\�a<b�a<U�a<p�a<f�a<y�a<p�a<[�a<i�a<H�a<M�a<B�a<:�a<�a<(�a<
�a<�a<��a<Ҭa<Ƭa<��a<��a<t�a<V�a</�a<�a<�a<��a<��a<��a<[�a<3�a<�a<۪a<��a<|�a<=�a<��a<کa<��a<b�a<6�a<��a<��a<u�a<8�a<�a<Ƨa<b�a<!�a<Ѧa<y�a<;�a<�a<��a<;�a< �a<��a<X�a<��a<��a<=�a<͢a<��a<"�a<��a<T�a<�a<x�a<�a<��a<O�a<�a<w�a<�a<��a<-�a<Ɯa<E�a<՛a<s�a<�a<��a</�a<��a<=�a<ݘa<k�a<�a<��a< �a<Ȗa<J�a<�a<��a<#�a<��a<V�a<�a<��a<X�a<�a<��a<9�a<ݑa<��a<H�a<�a<��a<`�a<�a<͏a<��a<T�a<!�a<�a<��a<z�a<D�a<�a<؍a<��a<��a<x�a<X�a<C�a<'�a<��a<�a<�a<�a<یa<Ìa<ӌa<��a<Ȍa<̌a<ٌa<Ԍa<��a<�a<$�a<L�a<�  �  E�a<��a<��a<ˍa<؍a<�a<R�a<e�a<��a<ߎa<�a<W�a<��a<Տa<
�a<f�a<��a<	�a<:�a<��a<�a<<�a<��a<�a<T�a<��a<�a<��a<ʔa<G�a<��a<)�a<~�a< �a<r�a<a<h�a<��a<2�a<��a<	�a<y�a<��a<��a<�a<w�a<Μa<Z�a<ԝa<C�a<۞a<!�a<��a<�a<��a<�a<Y�a<ߡa<0�a<��a<�a<��a<�a<R�a<��a<��a<�a<ҥa<3�a<z�a<¦a< �a<l�a<٧a<�a<��a<��a<��a<M�a<o�a<˩a<�a<0�a<V�a<��a<۪a<�a<?�a<O�a<��a<��a<��a<#�a<#�a<d�a<Y�a<��a<��a<��a<լa<�a<�a<�a<I�a<1�a<U�a<F�a<K�a<p�a<^�a<v�a<\�a<a�a<U�a<g�a<`�a<N�a<r�a<*�a<W�a<'�a<�a<�a<�a<�a<Ŭa<̬a<��a<��a<c�a<G�a<G�a<	�a<�a<ѫa<��a<��a<N�a</�a<�a<ڪa<��a<��a<5�a< �a<�a<��a<��a<�a<�a<��a<x�a<>�a<ڧa<��a<O�a<+�a<ʦa<��a<H�a<٥a<��a<7�a<��a<��a<:�a<ۣa<��a<D�a<ۢa<��a<	�a<��a<Z�a<�a<��a<�a<��a<9�a<�a<l�a<��a<��a<�a<Ϝa<C�a<�a<w�a<�a<��a<�a<ęa<K�a<�a<d�a<�a<��a<�a<ɖa<E�a<
�a<z�a<'�a<Ҕa<P�a<�a<��a<>�a<Вa<��a<:�a<�a<��a<'�a<�a<��a<n�a<0�a<ȏa<��a<<�a<#�a<ώa<��a<m�a<@�a<�a<�a<�a<��a<��a<R�a<1�a<5�a<�a<	�a<݌a<Ԍa<��a<όa<Ɍa<��a<�a<��a<��a<��a<��a<�a<	�a<5�a<�  �  b�a<f�a<��a<��a<�a<�a<>�a<a�a<��a<�a<�a<\�a<��a<֏a<�a<d�a<��a< �a<K�a<��a<ˑa<=�a<��a<�a<U�a<��a<�a<v�a<�a<P�a<��a<�a<��a<�a<^�a<̗a<?�a<��a<%�a<��a<(�a<��a<�a<m�a<��a<V�a<�a<`�a<Νa<$�a<��a<2�a<��a<�a<��a<��a<g�a<�a<J�a<��a<�a<z�a<ɣa<P�a<��a<#�a<b�a<֥a<�a<��a<�a<<�a<��a<Ƨa<�a<]�a<��a<�a<0�a<t�a<��a<�a<=�a<|�a<��a<Ӫa<�a<6�a<|�a<��a<��a<ëa<�a<4�a<W�a<r�a<��a<��a<ɬa<�a<��a< �a<!�a<�a<"�a<D�a<[�a<f�a<T�a<e�a<Z�a<x�a<m�a<u�a<l�a<X�a<O�a<G�a<<�a<1�a<$�a<�a<�a<
�a<�a<�a<��a<��a<��a<w�a<a�a<3�a<�a<ҫa<ԫa<��a<��a<\�a<0�a<�a<تa<��a<}�a<G�a<�a<��a<��a<l�a<C�a<�a<��a<o�a<.�a<�a<��a<v�a<�a<Ѧa<}�a<5�a<�a<��a<?�a<�a<��a<Y�a<��a<��a<+�a<ߢa<h�a<)�a<��a<U�a<Ϡa<v�a<%�a<��a<U�a<�a<x�a<	�a<��a<4�a<��a<S�a<ٛa<R�a<�a<��a<5�a<��a<O�a<Ϙa<w�a<�a<��a<9�a<��a<K�a<�a<��a<�a<��a<V�a<��a<��a<K�a<��a<��a<3�a<�a<��a<U�a<��a<��a<;�a<�a<ُa<��a<V�a<�a<ߎa<��a<z�a<P�a<�a<�a<��a<��a<z�a<g�a<L�a<�a<�a<�a<��a<��a<�a<ӌa<��a<��a<a<ƌa<Ќa<܌a<�a<�a<,�a<=�a<�  �  i�a<c�a<��a<��a<�a<�a<!�a<��a<��a<��a<
�a<F�a<��a<ӏa<,�a<P�a<��a<�a<L�a<��a<��a<y�a<k�a<�a<K�a<��a<!�a<o�a<��a<0�a<��a<�a<��a<��a<_�a<�a<4�a<ژa<�a<��a<�a<��a<�a<j�a<�a<F�a<��a<4�a<םa<e�a<��a<B�a<��a<�a<x�a<��a<l�a<ǡa<E�a<��a<)�a<��a<	�a<h�a<��a<-�a<P�a<�a<"�a<��a<Ԧa<�a<|�a<��a<:�a<Y�a<��a<��a<7�a<��a<��a<��a<�a<x�a<��a<�a<�a<&�a<��a<a�a<�a<��a<�a<6�a<6�a<o�a<|�a<��a<Ǭa<Ьa<�a<�a<6�a<�a<g�a<3�a<@�a<i�a<C�a<��a<U�a<|�a<W�a<f�a<G�a<b�a<u�a<<�a<f�a<)�a<D�a<+�a<�a<��a<Ӭa<�a<��a<��a<z�a<x�a<Q�a<�a<I�a<�a<�a<��a<u�a<R�a<.�a<�a<Īa<��a<a�a<G�a<�a<�a<שa<7�a<D�a<�a<��a<�a<(�a<�a<��a<a�a<��a<�a<��a<6�a< �a<��a<i�a<�a<��a<>�a<�a<��a<(�a<��a<Y�a<2�a<��a<^�a<�a<��a<4�a<��a<O�a<Ӟa<x�a<�a<��a</�a<��a<`�a<�a<��a<�a<k�a<?�a<��a<^�a<Ҙa<t�a<��a<��a<&�a<��a<t�a<�a<��a<#�a<��a<{�a<ԓa<��a<*�a<�a<��a<@�a<�a<|�a<Z�a<��a<Րa<q�a<'�a<ۏa<y�a<S�a<�a<�a<��a<h�a<?�a<�a<�a<��a<̍a<i�a<L�a<O�a<	�a<*�a<�a<��a<ˌa<Ҍa<��a<ˌa<�a<��a<��a<Ȍa<��a<�a<�a<�a<"�a<�  �  b�a<f�a<��a<��a<�a<�a<>�a<a�a<��a<�a<�a<\�a<��a<֏a<�a<d�a<��a< �a<K�a<��a<ˑa<=�a<��a<�a<U�a<��a<�a<v�a<�a<P�a<��a<�a<��a<�a<^�a<̗a<?�a<��a<%�a<��a<(�a<��a<�a<m�a<��a<V�a<�a<`�a<Νa<$�a<��a<2�a<��a<�a<��a<��a<g�a<�a<J�a<��a<�a<z�a<ɣa<P�a<��a<#�a<b�a<֥a<�a<��a<�a<<�a<��a<Ƨa<�a<]�a<��a<�a<0�a<t�a<��a<�a<=�a<|�a<��a<Ӫa<�a<6�a<|�a<��a<��a<ëa<�a<4�a<W�a<r�a<��a<��a<ɬa<�a<��a< �a<!�a<�a<"�a<D�a<[�a<f�a<T�a<e�a<Z�a<x�a<m�a<u�a<l�a<X�a<O�a<G�a<<�a<1�a<$�a<�a<�a<
�a<�a<�a<��a<��a<��a<w�a<a�a<3�a<�a<ҫa<ԫa<��a<��a<\�a<0�a<�a<تa<��a<}�a<G�a<�a<��a<��a<l�a<C�a<�a<��a<o�a<.�a<�a<��a<v�a<�a<Ѧa<}�a<5�a<�a<��a<?�a<�a<��a<Y�a<��a<��a<+�a<ߢa<h�a<)�a<��a<U�a<Ϡa<v�a<%�a<��a<U�a<�a<x�a<	�a<��a<4�a<��a<S�a<ٛa<R�a<�a<��a<5�a<��a<O�a<Ϙa<w�a<�a<��a<9�a<��a<K�a<�a<��a<�a<��a<V�a<��a<��a<K�a<��a<��a<3�a<�a<��a<U�a<��a<��a<;�a<�a<ُa<��a<V�a<�a<ߎa<��a<z�a<P�a<�a<�a<��a<��a<z�a<g�a<L�a<�a<�a<�a<��a<��a<�a<ӌa<��a<��a<a<ƌa<Ќa<܌a<�a<�a<,�a<=�a<�  �  E�a<��a<��a<ˍa<؍a<�a<R�a<e�a<��a<ߎa<�a<W�a<��a<Տa<
�a<f�a<��a<	�a<:�a<��a<�a<<�a<��a<�a<T�a<��a<�a<��a<ʔa<G�a<��a<)�a<~�a< �a<r�a<a<h�a<��a<2�a<��a<	�a<y�a<��a<��a<�a<w�a<Μa<Z�a<ԝa<C�a<۞a<!�a<��a<�a<��a<�a<Y�a<ߡa<0�a<��a<�a<��a<�a<R�a<��a<��a<�a<ҥa<3�a<z�a<¦a< �a<l�a<٧a<�a<��a<��a<��a<M�a<o�a<˩a<�a<0�a<V�a<��a<۪a<�a<?�a<O�a<��a<��a<��a<#�a<#�a<d�a<Y�a<��a<��a<��a<լa<�a<�a<�a<I�a<1�a<U�a<F�a<K�a<p�a<^�a<v�a<\�a<a�a<U�a<g�a<`�a<N�a<r�a<*�a<W�a<'�a<�a<�a<�a<�a<Ŭa<̬a<��a<��a<c�a<G�a<G�a<	�a<�a<ѫa<��a<��a<N�a</�a<�a<ڪa<��a<��a<5�a< �a<�a<��a<��a<�a<�a<��a<x�a<>�a<ڧa<��a<O�a<+�a<ʦa<��a<H�a<٥a<��a<7�a<��a<��a<:�a<ۣa<��a<D�a<ۢa<��a<	�a<��a<Z�a<�a<��a<�a<��a<9�a<�a<l�a<��a<��a<�a<Ϝa<C�a<�a<w�a<�a<��a<�a<ęa<K�a<�a<d�a<�a<��a<�a<ɖa<E�a<
�a<z�a<'�a<Ҕa<P�a<�a<��a<>�a<Вa<��a<:�a<�a<��a<'�a<�a<��a<n�a<0�a<ȏa<��a<<�a<#�a<ώa<��a<m�a<@�a<�a<�a<�a<��a<��a<R�a<1�a<5�a<�a<	�a<݌a<Ԍa<��a<όa<Ɍa<��a<�a<��a<��a<��a<��a<�a<	�a<5�a<�  �  R�a<|�a<��a<��a<�a<�a<:�a<v�a<��a<Ύa<�a<Q�a<��a<؏a<�a<g�a<��a<��a<A�a<��a<�a<H�a<��a< �a<`�a<��a<�a<��a<��a<b�a<��a<�a<��a<�a<e�a<ӗa<=�a<��a<8�a<��a<'�a<��a<�a<�a<�a<m�a<�a<S�a<͝a<D�a<��a<�a<��a<�a<��a<��a<g�a<ۡa<C�a<��a<�a<u�a<�a<Q�a<��a<�a<y�a<ĥa<,�a<��a<�a<=�a<v�a<קa<�a<]�a<��a<��a<0�a<u�a<©a<�a<J�a<p�a<��a<٪a<�a<F�a<p�a<��a<«a<�a<��a<(�a<W�a<q�a<��a<��a<Ƭa<�a<�a<
�a<�a<�a<<�a<B�a<L�a<\�a<b�a<U�a<p�a<f�a<y�a<p�a<[�a<i�a<H�a<M�a<B�a<:�a<�a<(�a<
�a<�a<��a<Ҭa<Ƭa<��a<��a<t�a<V�a</�a<�a<�a<��a<��a<��a<[�a<3�a<�a<۪a<��a<|�a<=�a<��a<کa<��a<b�a<6�a<��a<��a<u�a<8�a<�a<Ƨa<b�a<!�a<Ѧa<y�a<;�a<�a<��a<;�a< �a<��a<X�a<��a<��a<=�a<͢a<��a<"�a<��a<T�a<�a<x�a<�a<��a<O�a<�a<w�a<�a<��a<-�a<Ɯa<E�a<՛a<s�a<�a<��a</�a<��a<=�a<ݘa<k�a<�a<��a< �a<Ȗa<J�a<�a<��a<#�a<��a<V�a<�a<��a<X�a<�a<��a<9�a<ݑa<��a<H�a<�a<��a<`�a<�a<͏a<��a<T�a<!�a<�a<��a<z�a<D�a<�a<؍a<��a<��a<x�a<X�a<C�a<'�a<��a<�a<�a<�a<یa<Ìa<ӌa<��a<Ȍa<̌a<ٌa<Ԍa<��a<�a<$�a<L�a<�  �  ]�a<q�a<��a<��a<��a<�a<,�a<��a<��a<�a<�a<C�a<��a<Ïa< �a<T�a<��a<ܐa<^�a<��a<ߑa<R�a<��a<�a<Q�a<��a<�a<w�a<�a<<�a<��a<�a<��a<�a<c�a<�a<6�a<Ƙa</�a<��a<�a<��a<	�a<w�a<��a<\�a<�a<W�a<ʝa<G�a<��a<G�a<��a<�a<��a<�a<f�a<͡a<H�a<��a<6�a<~�a<�a<R�a<��a<!�a<f�a<ڥa<(�a<��a<צa<�a<�a<ͧa<+�a<X�a<��a<��a<2�a<��a<��a<��a<&�a<r�a<��a<תa<�a<3�a<w�a<��a<ʫa<ݫa<�a<K�a<6�a<}�a<��a<��a<��a<ެa<�a<�a<3�a<�a<C�a<6�a<V�a<W�a<W�a<g�a<e�a<t�a<^�a<c�a<X�a<e�a<^�a<D�a<U�a<3�a</�a<&�a<�a<��a<ެa<ݬa<��a<��a<��a<l�a<]�a<!�a<$�a<߫a<�a<��a<r�a<]�a<�a<
�a<Ȫa<��a<Z�a<Y�a<�a<ʩa<��a<Y�a<<�a<�a<��a<w�a<0�a<��a<��a<e�a<�a<�a<��a<9�a<��a<��a<V�a<��a<��a<<�a<�a<��a<5�a<�a<o�a<"�a<��a<Q�a<�a<}�a<9�a<��a<N�a<۞a<o�a<�a<��a<2�a<��a<m�a<ݛa<r�a<�a<��a<3�a<��a<S�a<ؘa<l�a<��a<��a<)�a<��a<e�a<ߕa<��a<$�a<��a<k�a<��a<��a<4�a<�a<��a<7�a<�a<��a<O�a<�a<��a<V�a<#�a<�a<x�a<`�a<�a<�a<��a<w�a<:�a<�a<�a<��a<��a<l�a<a�a<=�a<�a<�a<��a<��a<ьa<Όa<��a<Όa<͌a<��a<��a<Ҍa<�a<��a<��a<�a<,�a<�  �  _�a<v�a<��a<Ía<ߍa<�a<@�a<q�a<��a<Ԏa<�a<W�a<��a<̏a<+�a<R�a<��a<��a<:�a<��a<�a<G�a<��a<��a<P�a<��a<�a<��a<�a<D�a<��a<�a<��a<��a<a�a<˗a<O�a<��a<$�a<��a<�a<��a<�a<v�a<�a<p�a<Ԝa<S�a<a<F�a<��a< �a<��a<�a<~�a<��a<o�a<ˡa<N�a<��a<�a<{�a<�a<E�a<��a<�a<w�a<ѥa<*�a<��a<�a<(�a<��a<ǧa<�a<l�a<��a<�a<@�a<u�a<��a<��a<2�a<u�a<��a<Ӫa<�a<8�a<b�a<��a<��a<�a<�a<"�a<N�a<{�a<{�a<��a<��a<֬a<��a<��a<�a<+�a<9�a<A�a<T�a<S�a<e�a<_�a<c�a<u�a<o�a<i�a<m�a<V�a<Y�a<[�a<;�a<@�a<2�a<�a<�a<��a<�a<߬a<��a<��a<��a<k�a<V�a<6�a<�a<�a<ƫa<��a<��a<X�a<&�a<�a<ƪa<��a<s�a<5�a<
�a<٩a<��a<t�a<*�a<�a<��a<n�a<>�a<��a<��a<h�a< �a<Φa<��a<8�a<�a<��a<H�a<�a<��a<A�a<��a<��a<4�a<آa<��a<�a<��a<I�a<�a<��a<�a<��a<S�a<ٞa<w�a<�a<��a<8�a<��a<C�a<ۛa<u�a<��a<��a<�a<��a<J�a<ژa<v�a<�a<��a<5�a<��a<S�a<��a<�a<�a<Ŕa<W�a<��a<��a<@�a<�a<��a<3�a<�a<��a<;�a<��a<��a<a�a<�a<Ǐa<��a<_�a<�a<�a<��a<o�a<F�a<	�a<�a<ča<��a<w�a<_�a<9�a<+�a<	�a<��a<��a<�a<Ԍa<Ԍa<��a<Ȍa<Ռa<Ōa<ߌa<�a<�a<�a<!�a<<�a<�  �  B�a<}�a<��a<̍a<�a<�a<F�a<[�a<��a<͎a<#�a<^�a<��a<Ώa<�a<^�a<��a<�a<M�a<��a<��a<2�a<��a<�a<l�a<��a<�a<��a<Ӕa<O�a<��a<4�a<��a<�a<g�a<ӗa<B�a<��a<G�a<��a<�a<��a<��a<��a<�a<��a<לa<Y�a<˝a<=�a<��a< �a<��a<�a<�a<��a<c�a<̡a<9�a<Ǣa<�a<��a<�a<I�a<��a<�a<��a<åa<1�a<|�a<�a</�a<}�a<�a<�a<a�a<��a<��a<7�a<z�a<ةa<�a<:�a<g�a<��a<ުa<	�a<T�a<`�a<��a<��a<�a<�a<1�a<h�a<e�a<��a<��a<¬a<Ҭa<��a<�a<	�a<.�a<$�a<J�a<M�a<_�a<q�a<]�a<p�a<W�a<r�a<^�a<n�a<t�a<M�a<Q�a<@�a<9�a<"�a<1�a<�a<�a<�a<¬a<Ǭa<��a<��a<}�a<K�a<;�a<��a<��a<��a<��a<��a<K�a<(�a<��a<Ҫa<��a<��a<H�a<�a<�a<��a<r�a<(�a<�a<��a<y�a<<�a<�a<��a<Y�a<6�a<٦a<��a<>�a<�a<��a<@�a<�a<��a<C�a<��a<��a<@�a<΢a<��a<�a<��a<R�a<�a<��a<�a<Пa<D�a<ڞa<r�a<�a<��a<#�a<לa<J�a<�a<w�a<��a<��a<�a<Йa<<�a<�a<f�a<	�a<��a<'�a<ٖa<N�a<�a<��a<$�a<��a<[�a<�a<��a<H�a<�a<��a<>�a<�a<��a<8�a<��a<��a<j�a<�a<֏a<��a<H�a<�a<؎a<��a<j�a<I�a<(�a<ۍa<Ǎa<��a<��a<Y�a<E�a<6�a<�a<�a<،a<�a<Ɍa<Ռa<݌a<��a<̌a<ˌa<،a<یa<�a<�a<�a<B�a<�  �  W�a<z�a<��a<��a<�a<�a<A�a<v�a<��a<ڎa<�a<H�a<��a<ԏa<
�a<j�a<��a<�a<O�a<��a<�a<O�a<��a<��a<^�a<��a<�a<x�a<�a<M�a<��a<�a<��a<�a<b�a<�a<8�a<Ƙa<,�a<��a<�a<��a< �a<��a<�a<f�a<�a<P�a<ҝa<H�a<��a<0�a<��a<
�a<��a<�a<[�a<סa<<�a<��a<#�a<}�a<�a<V�a<��a<�a<u�a<ɥa<,�a<{�a<ܦa<(�a<s�a<Χa<)�a<]�a<��a<��a<5�a<��a<��a<�a<7�a<s�a<��a<ڪa<�a<E�a<h�a<��a<ɫa<�a<�a<9�a<F�a<m�a<��a<��a<��a<�a<�a<�a<�a<#�a<:�a<J�a<F�a<\�a<V�a<b�a<q�a<m�a<i�a<f�a<Y�a<b�a<c�a<H�a<]�a<6�a<4�a<'�a<�a<��a<�a<׬a<ìa<��a<��a<w�a<J�a<7�a<�a<�a<ͫa<��a<v�a<\�a<.�a<�a<ުa<��a<i�a<J�a<�a<ީa<��a<c�a<+�a<��a<��a<{�a<1�a<��a<��a<_�a<�a<ڦa<��a<8�a<��a<��a<V�a<��a<��a<A�a<�a<��a<@�a<Ӣa<y�a<�a<��a<Y�a<��a<��a<#�a<��a<B�a<�a<h�a<��a<��a<&�a<��a<Z�a<ݛa<y�a<�a<��a<)�a<��a<B�a<ܘa<e�a<�a<��a<�a<��a<c�a<�a<��a<%�a<��a<e�a<��a<��a<E�a<�a<��a<:�a<ܑa<��a<@�a<�a<��a<f�a<�a<ޏa<��a<Q�a< �a<юa<��a<y�a<:�a<�a<�a<��a<��a<��a<R�a<C�a<�a<�a<�a<�a<݌a<ьa<��a<ˌa<Ҍa<Ìa<�a<Ռa<�a<��a<��a<�a<9�a<�  �  g�a<b�a<��a<��a<�a<�a<:�a<u�a<��a<؎a<�a<V�a<��a<ˏa<#�a<P�a<��a<��a<;�a<��a<�a<O�a<��a<��a<N�a<��a<�a<r�a<�a<<�a<Еa<�a<��a<��a<Y�a<ߗa<=�a<ǘa<�a<��a<�a<��a<�a<o�a<��a<]�a<�a<Q�a<ǝa<B�a<��a<&�a<��a<�a<y�a<��a<o�a<ơa<P�a<��a<�a<q�a<�a<K�a<��a<�a<f�a<ޥa<$�a<��a<֦a<-�a<��a<��a<%�a<_�a<��a<�a<9�a<��a<��a<�a<,�a<w�a<��a<ݪa<�a<1�a<p�a<��a<ƫa<ܫa< �a<*�a<R�a<x�a<{�a<��a<��a<լa<��a<��a<�a<�a<;�a<=�a<O�a<\�a<X�a<q�a<X�a<z�a<Z�a<|�a<x�a<I�a<e�a<G�a<Q�a</�a<7�a<�a<�a<�a<٬a<�a<��a<��a<��a<p�a<T�a</�a<�a<�a<ʫa<��a<��a<T�a<%�a<�a<Īa<��a<w�a<7�a<�a<ͩa<��a<f�a<4�a<�a<��a<|�a<+�a<��a<��a<��a<�a<Ѧa<��a</�a<��a<��a<V�a<ޤa<��a<P�a<�a<��a<-�a<�a<p�a<%�a<��a<N�a<�a<t�a<�a<��a<W�a<Ԟa<v�a<�a<��a<:�a<��a<N�a<Лa<q�a< �a<��a<1�a<��a<W�a<Ԙa<u�a<��a<��a<H�a<��a<_�a<�a<��a<�a<��a<b�a<��a<��a<:�a<�a<��a<=�a<�a<��a<I�a<�a<��a<U�a<�a<Ϗa<��a<\�a<�a<�a<��a<m�a<L�a<�a<�a<��a<��a<s�a<[�a<C�a<�a<�a<�a<��a<Όa<�a<��a<��a<Ԍa<��a<یa<Όa<�a<�a<�a<9�a<(�a<�  �  ]�a<o�a<��a<��a<ߍa<�a<E�a<k�a<��a<ڎa<�a<V�a<|�a<Џa<�a<Y�a<��a< �a<<�a<��a<��a<@�a<��a<�a<[�a<��a<�a<}�a<�a<?�a<��a<$�a<��a<��a<j�a<ڗa<S�a<��a<5�a<��a<�a<��a<�a<s�a<��a<q�a<֜a<T�a<̝a<B�a<Ȟa<�a<��a<�a<z�a<�a<d�a<ʡa<6�a<��a<�a<��a<�a<L�a<��a<�a<y�a<إa<'�a<��a<ڦa<!�a<v�a<֧a<�a<p�a<��a<��a<A�a<��a<ǩa<�a<)�a<s�a<��a<תa<�a<@�a<^�a<��a<��a<�a<�a<$�a<Z�a<_�a<��a<��a<��a<Ǭa<�a<�a<�a<@�a<3�a<H�a<J�a<Q�a<g�a<k�a<b�a<n�a<j�a<X�a<b�a<g�a<\�a<Z�a<K�a<D�a<2�a<#�a<�a<�a<�a<ݬa<��a<��a<��a<k�a<G�a<:�a<�a<�a<ͫa<��a<��a<B�a<+�a<��a<ͪa<��a<}�a<8�a<�a<�a<��a<s�a<"�a<��a<��a<s�a<6�a<��a<��a<W�a<&�a<٦a<��a<@�a<�a<��a<K�a<��a<��a<8�a<�a<��a<1�a<�a<��a<�a<��a<S�a<�a<��a<�a<��a<A�a<՞a<q�a<�a<��a< �a<Ĝa<E�a<�a<w�a<�a<��a<�a<��a<Q�a<טa<q�a<�a<��a< �a<ǖa<X�a<��a<��a<(�a<Ɣa<e�a<�a<��a<7�a<�a<��a<7�a<�a<��a<6�a<��a<��a<k�a<'�a<ɏa<��a<C�a<�a<؎a<��a<`�a<A�a<�a<�a<ٍa<��a<~�a<U�a<7�a<-�a<�a<��a<�a<݌a<Ìa<ʌa<Ќa<ˌa<Ԍa<Ռa<�a<�a<��a<
�a<�a<4�a<�  �  K�a<��a<��a<��a<�a<�a<J�a<\�a<��a<a<�a<L�a<��a<�a<��a<��a<��a<��a<E�a<��a<�a<6�a<��a<�a<g�a<��a<�a<��a<ߔa<m�a<��a<�a<��a<�a<d�a<ȗa<V�a<��a<B�a<��a<2�a<��a<�a<��a<؛a<n�a<��a<W�a<ʝa<&�a<��a<�a<��a<�a<��a<�a<Z�a<�a<0�a<��a<�a<w�a<Уa<G�a<��a<�a<}�a<��a<;�a<��a<�a<O�a<s�a<�a<	�a<t�a<��a<�a<<�a<p�a<ĩa<�a<[�a<o�a<��a<۪a<��a<L�a<g�a<��a<��a<ԫa<��a<$�a<S�a<]�a<��a<��a<Ҭa<ݬa<�a<�a<��a<%�a<�a<N�a<N�a<_�a<Y�a<Q�a<��a<`�a<��a<x�a<Y�a<q�a<I�a<X�a<<�a<A�a<%�a<+�a<�a<	�a<�a<ˬa<Ԭa<��a<��a<|�a<Q�a<@�a<��a<�a<��a<��a<{�a<Q�a<D�a<�a<��a<��a<t�a<@�a<��a<̩a<��a<x�a<)�a<�a<��a<p�a<F�a<�a<ҧa<`�a<�a<Цa<��a<:�a<ߥa<��a<4�a<
�a<��a<c�a<��a<��a<N�a<��a<��a<�a<��a<Q�a<Ҡa<~�a<�a<��a<:�a<��a<q�a<��a<��a<�a<Ȝa<:�a<֛a<Y�a<��a<��a<'�a<��a<3�a<�a<o�a<�a<��a<�a<іa<C�a<��a<{�a<�a<��a<Q�a<�a<��a<i�a<�a<��a<;�a<בa<��a<@�a<�a<��a<M�a<
�a<ɏa<��a<A�a<9�a<Ŏa<��a<v�a<9�a<�a<Ѝa<��a<��a<��a<Z�a<E�a<�a<��a<�a<�a<��a<�a<��a<ڌa<��a<ӌa<ƌa<��a<݌a<�a<�a<+�a<U�a<�  �  J�a<u�a<��a<��a<�a<�a<0�a<|�a<��a<�a<�a<K�a<��a<Ǐa<�a<T�a<��a<�a<O�a<��a<�a<R�a<��a<��a<J�a<Ǔa<%�a<�a<̔a<1�a<��a<�a<��a<�a<n�a<חa<R�a<��a<4�a<��a<�a<i�a<�a<�a<�a<^�a<�a<M�a<͝a<M�a<��a<<�a<��a<�a<x�a<�a<\�a<ɡa<5�a<��a<(�a<��a<��a<U�a<��a<�a<d�a<�a<1�a<��a<��a<*�a<��a<ԧa<$�a<v�a<��a<��a<J�a<��a<��a<�a<"�a<T�a<��a<�a<�a<+�a<m�a<��a<ͫa<�a<�a<;�a<G�a<d�a<��a<��a<��a<̬a<�a<�a<$�a<-�a<D�a<9�a<H�a<Z�a<^�a<w�a<i�a<a�a<I�a<p�a<h�a<k�a<^�a<W�a<N�a<?�a<5�a<+�a<�a<�a<ˬa<ʬa<��a<��a<��a<n�a<R�a<%�a<�a<��a<ثa<��a<z�a<J�a<!�a<��a<Ȫa<��a<k�a<J�a<�a<۩a<��a<\�a<2�a<�a<ƨa<��a<8�a<ݧa<��a<q�a<�a<�a<��a<D�a<�a<��a<O�a<��a<��a<J�a<̣a<��a<=�a<�a<q�a<�a<��a<T�a<��a<��a</�a<��a<?�a<Ӟa<k�a<��a<��a<�a<��a<_�a<�a<��a<
�a<��a<+�a<��a<Z�a<�a<n�a<ߗa<��a<-�a<Ŗa<^�a<��a<��a<+�a<ϔa<k�a<��a<��a<0�a<Βa<��a<F�a<��a<��a<F�a<�a<��a<d�a<(�a<��a<��a<H�a<�a<ӎa<��a<e�a<?�a<�a<��a<ƍa<��a<o�a<T�a<A�a<$�a<!�a<��a<�a<��a<یa<Ќa<Ԍa<͌a<ьa<،a<ތa<�a<�a<�a<(�a<�a<�  �  2�a<��a<6�a<I�a<u�a<��a<��a<�a<�a<~�a<��a<�a<*�a<H�a<��a<ؐa<I�a<��a<��a<*�a<e�a<ےa<�a<��a<ړa<Q�a<��a<�a<��a<��a<I�a<��a<�a<��a<�a<`�a<a<d�a<��a<:�a<��a<�a<��a<�a<��a<Ϝa<o�a<Ýa<8�a<��a<�a<��a<�a<��a<��a<h�a<ߡa<C�a<ɢa<�a<��a<ڣa<G�a<��a<�a<��a<Хa<[�a<��a<�a<b�a<��a<�a<=�a<��a<ɨa<�a<^�a<��a<��a<�a<z�a<��a<�a<�a<?�a<��a<��a<��a<�a<1�a<9�a<p�a<��a<��a<�a<�a<(�a<�a<L�a<j�a<`�a<��a<y�a<��a<��a<ͭa<ȭa<��a<�a<��a<!�a<έa<ҭa<ܭa<ʭa<�a<��a<��a<��a<��a<��a<��a<n�a<F�a<��a<�a<!�a<��a<ݬa<ڬa<��a<��a<F�a<M�a<�a<��a<ϫa<��a<��a<+�a<#�a<�a<��a<��a<1�a<�a<��a<ũa<Y�a<3�a<�a<��a<��a<�a<�a<��a<R�a<��a<��a<a�a<�a<�a<i�a<&�a<��a<n�a<;�a<��a<i�a<֢a<��a<�a<��a<U�a<ݠa<��a<�a<֟a<R�a<�a<��a<�a<��a<+�a<Ĝa<E�a<ݛa<{�a<��a<a<'�a<�a<I�a<�a<��a<�a<ȗa<G�a<��a<k�a<�a<��a<@�a<��a<��a<?�a<��a<��a<*�a<��a<��a<�a<��a<b�a<>�a<Րa<��a<M�a<�a<��a<��a<��a<$�a<
�a<�a<��a<��a<8�a<0�a<��a<��a<Սa<��a<��a<x�a<ȍa<h�a<c�a<j�a<Y�a<��a<W�a<g�a<j�a<��a<��a<��a<��a<��a<�  �  �a<��a<6�a<N�a<w�a<��a<Ԏa<�a</�a<z�a<��a<؏a<�a<h�a<��a<�a<0�a<��a<�a<9�a<r�a<�a<&�a<��a<ݓa<A�a<��a<��a<d�a<ɕa<D�a<��a<�a<u�a<�a<f�a<ɘa<9�a<��a<%�a<��a< �a<y�a<�a<{�a<ޜa<d�a<ʝa<U�a<��a<4�a<��a<�a<}�a<�a<i�a<סa<>�a<��a<&�a<��a<��a<W�a<Ѥa<�a<��a<٥a<F�a<��a<�a<7�a<��a<�a<8�a<��a<Ψa<'�a<j�a<��a<�a<'�a<j�a<��a<Ϫa<��a<C�a<x�a<��a<�a<��a<@�a<J�a<��a<��a<��a<Ҭa<�a<�a<2�a<>�a<Q�a<x�a<��a<��a<��a<��a<��a<ȭa<˭a<ޭa<ʭa<ԭa<ϭa<ۭa<֭a<ҭa<ȭa<��a<��a<��a<��a<��a<��a<s�a<R�a<@�a< �a< �a<��a<ެa<¬a<��a<��a<Y�a<I�a< �a<�a<��a<��a<s�a<@�a<
�a<�a<��a<��a<?�a<&�a<ԩa<��a<\�a<#�a<�a<��a<Z�a<�a<ߧa<��a<L�a<�a<��a<g�a<	�a<��a<b�a<�a<��a<S�a<��a<��a<X�a<�a<��a<#�a<աa<d�a<��a<��a<2�a<��a<J�a<�a<}�a<	�a<��a<?�a<לa<g�a<�a<��a<�a<��a<0�a<әa<T�a<�a<u�a<�a<��a<B�a<ؖa<p�a<�a<��a<@�a<�a<��a</�a<œa<j�a<
�a<Ēa<s�a<�a<ۑa<{�a<L�a<�a<��a<r�a<'�a<ڏa<��a<n�a<<�a<��a<Ȏa<��a<��a<Q�a<;�a<�a<�a<ԍa<��a<��a<��a<{�a<h�a<l�a<d�a<b�a<]�a<_�a<p�a<m�a<y�a<��a<��a<��a<ōa<�  �  ܍a<�a<%�a<R�a<��a<��a<ێa<�a<3�a<V�a<��a<ُa<�a<}�a<��a<
�a</�a<��a<Αa<�a<u�a<̒a<1�a<u�a<��a<;�a<��a<�a<d�a<��a</�a<��a<�a<u�a<��a<W�a<ژa</�a<��a<�a<��a<$�a<{�a<�a<_�a<�a<T�a<ŝa<N�a<��a<4�a<��a<�a<|�a<�a<d�a<ʡa<[�a<��a<)�a<q�a<��a<?�a<¤a<�a<v�a<�a</�a<��a<�a<U�a<��a<ڧa<K�a<z�a<ۨa<�a<i�a<��a<�a<4�a<U�a<Īa<۪a<�a<M�a<n�a<��a<ūa<�a<(�a<E�a<q�a<��a<��a<Ҭa<�a<��a<?�a<H�a<T�a<v�a<j�a<��a<��a<��a<��a<έa<խa<ǭa<�a<ɭa<��a<ڭa<ɭa<�a<��a<ϭa<��a<��a<��a<��a<y�a<j�a<��a<7�a<C�a<�a<��a<�a<��a<��a<q�a<]�a<%�a<�a<�a<��a<��a<I�a<]�a<�a<�a<��a<r�a<A�a<�a<ߩa<��a<t�a<�a<�a<��a<Y�a<C�a<˧a<��a<J�a<�a<��a<X�a<�a<��a<v�a<�a<ˤa<v�a<��a<��a<<�a<��a<��a<�a<Ρa<G�a< �a<v�a<2�a<��a<d�a<�a<p�a<&�a<��a<B�a<��a<_�a<՛a<��a<�a<��a<D�a<��a<l�a<�a<��a<2�a<��a<U�a<ϖa<~�a<�a<��a<D�a<�a<��a<�a<�a<u�a<#�a<Βa<i�a<1�a<��a<��a<4�a<�a<��a<S�a<'�a<ڏa<��a<O�a<H�a<�a<ʎa<��a<b�a<V�a<�a<�a<ݍa<ۍa<��a<��a<��a<p�a<��a<l�a<V�a<p�a<N�a<p�a<`�a<|�a<m�a<��a<��a<��a<��a<�  �  �a<�a<)�a<Q�a<��a<��a<ߎa<��a<H�a<v�a<��a<�a<�a<d�a<��a<�a<-�a<��a<͑a<6�a<��a<̒a<6�a<��a<�a<I�a<��a<	�a<j�a<ɕa<2�a<��a<�a<��a<��a<K�a<Ԙa<C�a<��a<*�a<��a<�a<��a<��a<p�a<�a<[�a<۝a<U�a<��a<G�a<��a<�a<��a<��a<e�a<աa<D�a<��a<#�a<��a<�a<b�a<̤a<*�a<��a<�a<>�a<��a<�a<<�a<��a<�a<B�a<��a<ڨa<�a<j�a<��a<�a<2�a<`�a<��a<ժa<�a<A�a<{�a<��a<۫a<�a<*�a<b�a<��a<��a<Ƭa<Ѭa<��a<�a<.�a<=�a<f�a<q�a<��a<��a<��a<��a<ŭa<ɭa<έa<ѭa<ۭa<׭a<Эa<˭a<ݭa<ѭa<έa<Эa<��a<��a<��a<��a<��a<`�a<N�a<E�a<0�a<�a<��a<�a<ɬa<��a<w�a<r�a<E�a<�a<��a<��a<��a<j�a<D�a<�a<�a<��a<��a<\�a<�a<�a<��a<d�a<+�a<�a<��a<_�a<�a<ͧa<��a<C�a<��a<��a<M�a<�a<��a<j�a<�a<��a<U�a<�a<��a<M�a<�a<��a<4�a<աa<b�a<�a<��a<,�a<��a<Q�a<�a<{�a<�a<��a<;�a<ɜa<r�a<��a<��a<�a<��a<7�a<˙a<R�a<�a<z�a<�a<��a<L�a<�a<}�a<�a<��a<P�a<�a<��a<%�a<Óa<p�a<�a<a<v�a<�a<֑a<��a<6�a<��a<��a<[�a<,�a<ُa<��a<l�a<7�a<��a<ݎa<��a<��a<g�a<'�a<�a<��a<Սa<��a<��a<��a<~�a<j�a<\�a<j�a<`�a<d�a<q�a<T�a<��a<��a<��a<��a<��a<a<�  �  ��a<��a<A�a<Q�a<q�a<��a<Ďa<�a<$�a<m�a<��a<�a< �a<^�a<��a<�a<A�a<��a<ؑa<'�a<m�a<Вa<!�a<��a<̓a<Q�a<��a<�a<|�a<˕a<[�a<��a<�a<��a<�a<[�a<Ęa<J�a<��a<<�a<��a<�a<��a<�a<��a<Ӝa<_�a<ȝa<:�a<��a<�a<��a<�a<��a<�a<l�a<ޡa<:�a<��a<�a<��a<�a<W�a<��a<�a<��a<ɥa<V�a<��a<��a<L�a<��a<�a<%�a<��a<Ϩa<�a<`�a<��a<�a<�a<��a<��a<�a<�a<J�a<��a<��a<�a<��a<&�a<G�a<r�a<��a<��a<�a<�a<!�a<.�a<E�a<f�a<i�a<��a<��a<��a<��a<��a<ĭa<ɭa<�a<ƭa<�a<ӭa<�a<�a<��a<խa<��a<��a<��a<��a<��a<��a<��a<Q�a<X�a<�a<+�a<��a<جa<ʬa<��a<��a<N�a<<�a<�a<��a<ūa<��a<~�a<:�a<�a<�a<��a<}�a<9�a<�a<Ωa<��a<K�a<3�a<�a<��a<q�a<�a<��a<��a<B�a<�a<��a<\�a<�a<ƥa<M�a<(�a<Ƥa<b�a<�a<��a<f�a<ڢa<��a<!�a<��a<`�a<�a<��a<%�a<ȟa<N�a<�a<��a<�a<��a<2�a<Ҝa<L�a<�a<x�a<�a<��a< �a<�a<R�a<��a<��a<�a<ʗa</�a<�a<r�a<�a<��a<L�a<�a<y�a<J�a<ɓa<��a<�a<˒a<��a<�a<�a<y�a<3�a<�a<��a<h�a<$�a<�a<��a<z�a<8�a<�a<ݎa<��a<~�a<B�a<1�a<��a<�a<Ѝa<��a<��a<�a<��a<m�a<��a<o�a<O�a<k�a<W�a<g�a<j�a<��a<��a<��a<Ѝa<ōa<�  �  �a<�a<&�a<E�a<��a<��a<Ǝa<�a<8�a<o�a<��a<Џa<+�a<k�a<��a<��a<A�a<p�a<Ցa<.�a<{�a<ߒa<!�a<��a<�a<<�a<��a<�a<s�a<ѕa<3�a<��a<!�a<��a<�a<m�a<Řa<M�a<��a<�a<��a<�a<��a<��a<n�a<ޜa<a�a<ϝa<?�a<��a<1�a<��a<	�a<��a<
�a<d�a<ϡa<Y�a<��a<�a<��a<�a<\�a<��a<�a<��a<ܥa<=�a<��a<�a<I�a<��a<ݧa<<�a<��a<ͨa<%�a<_�a<��a<��a<�a<\�a<��a<�a<�a<D�a<t�a<��a<ݫa<��a<2�a<S�a<|�a<��a<��a<�a<
�a<��a<4�a<R�a<O�a<n�a<��a<��a<��a<��a<��a<ԭa<ía<έa<׭a<�a<٭a<ӭa<��a<�a<ҭa<��a<ͭa<��a<��a<��a<g�a<j�a<Y�a<N�a<1�a<�a<�a<�a<Ȭa<��a<��a<b�a<>�a<�a<ܫa<Ыa<��a<W�a<P�a<�a<ͪa<��a<��a<H�a<�a<Ωa<��a<l�a<�a<ߨa<��a<h�a<�a<Χa<�a<U�a<��a<��a<o�a<�a<ɥa<m�a<��a<��a<c�a<�a<��a<K�a<�a<��a<(�a<��a<f�a<��a<��a<�a<��a<g�a<�a<u�a<%�a<��a<(�a<ʜa<]�a<�a<{�a<�a<��a<3�a<ʙa<_�a<�a<��a<�a<��a<F�a<�a<p�a<�a<��a<H�a<��a<�a<!�a<Γa<z�a< �a<Œa<n�a<%�a<ؑa<{�a<?�a<�a<��a<d�a<�a<�a<��a<X�a<=�a<�a<Ǝa<��a<�a<[�a<=�a<�a<�a<��a<��a<��a<��a<��a<s�a<e�a<K�a<r�a<g�a<R�a<}�a<d�a<��a<��a<��a<��a<̍a<�  �  �a<�a<%�a<R�a<w�a<��a<ߎa<��a<<�a<r�a<��a<ۏa<�a<l�a<��a<��a<&�a<��a<ؑa<2�a<|�a<̒a<8�a<��a<�a<>�a<��a<�a<b�a<��a<:�a<��a<�a<r�a<�a<\�a<͘a<)�a<��a<"�a<��a<�a<|�a<�a<c�a<�a<O�a<۝a<F�a<��a<=�a<��a< �a<y�a<��a<n�a<ܡa<F�a<��a<'�a<��a<��a<N�a<��a</�a<u�a<�a<1�a<��a<�a<=�a<��a<�a<B�a<u�a<Ҩa<�a<g�a<��a<۩a<4�a<c�a<��a<Ϊa<�a<M�a<o�a<��a<̫a<�a<$�a<O�a<��a<��a<Ĭa<Ǭa<��a<�a<6�a<:�a<T�a<}�a<��a<��a<��a<��a<��a<­a<խa<ͭa<�a<ҭa<ڭa<�a<׭a<ҭa<��a<ǭa<��a<��a<��a<��a<��a<u�a<^�a<=�a<<�a<�a<��a<ެa<��a<��a<y�a<f�a<A�a<�a<�a<��a<��a<r�a<G�a< �a<�a<��a<��a<H�a<�a<�a<��a<m�a< �a<�a<��a<X�a<*�a<էa<��a<:�a<�a<��a<]�a<�a<��a<m�a<�a<äa<Z�a<��a<��a<@�a<��a<��a<4�a<ǡa<T�a<�a<��a<4�a<��a<R�a<�a<��a<�a<��a<@�a<Ɯa<j�a<�a<~�a<!�a<��a<D�a<��a<k�a<�a<{�a<$�a<��a<L�a<ʖa<u�a<�a<��a<C�a<۔a<��a<(�a<ޓa<i�a<!�a<Βa<i�a<,�a<Ǒa<��a<0�a<�a<��a<d�a<*�a<Ϗa<��a<q�a<?�a<��a<ˎa<��a<|�a<_�a<&�a<�a<�a<΍a<��a<��a<��a<y�a<s�a<r�a<e�a<a�a<K�a<g�a<i�a<y�a<m�a<��a<��a<��a<ҍa<�  �  ��a<��a<3�a<]�a<m�a<��a<Ԏa<
�a<3�a<h�a<��a<�a<'�a<Z�a<��a<�a<E�a<��a<��a<$�a<~�a<ےa<,�a<��a<ۓa<P�a<��a< �a<w�a<ەa<?�a<��a<�a<��a<�a<F�a<ݘa<F�a<��a<%�a<��a<�a<��a<�a<t�a<�a<Y�a<Нa<F�a<��a<.�a<��a<�a<��a<��a<h�a<ޡa<A�a<��a<�a<}�a<�a<\�a<��a<#�a<��a<ޥa<B�a<��a<�a<I�a<��a<�a<)�a<��a<�a<�a<_�a<��a<�a<�a<f�a<��a<�a<�a<E�a<��a<��a<ԫa<�a<.�a<U�a<v�a<��a<Ǭa<�a<�a<+�a<)�a<L�a<o�a<_�a<}�a<��a<��a<��a<��a<��a<حa<ݭa<ʭa<�a<حa<ޭa<ԭa<��a<ѭa<έa<��a<��a<��a<|�a<�a<q�a<[�a<R�a<!�a<�a<�a<Ԭa<��a<��a<��a<]�a<7�a<��a< �a<˫a<��a<��a<4�a<�a<��a<��a<z�a<J�a<�a<کa<��a<Z�a<2�a<�a<��a<m�a<%�a<ڧa<��a<7�a<�a<��a<H�a<�a<¥a<P�a<�a<��a<b�a<	�a<��a<Q�a<�a<��a<*�a<ơa<e�a<��a<��a<!�a<͟a<R�a<�a<��a<�a<��a<6�a<��a<^�a<�a<��a<�a<��a<5�a<Ιa<X�a<�a<��a<�a<��a<3�a<�a<��a<�a<��a<Y�a<�a<�a<+�a<ӓa<}�a<�a<ƒa<|�a<�a<ϑa<��a<;�a<�a<��a<O�a<-�a<�a<��a<��a<2�a<
�a<�a<��a<t�a<Q�a<6�a<�a<�a<ɍa<Ía<��a<��a<��a<r�a<o�a<a�a<I�a<f�a<n�a<M�a<z�a<��a<y�a<��a<��a<΍a<�  �  �a<��a<6�a<D�a<}�a<��a<a<�a<,�a<��a<��a<ޏa<*�a<]�a<��a<�a<H�a<s�a<�a<=�a<x�a<�a<�a<��a<ݓa<C�a<��a<��a<n�a<a<?�a<��a<�a<{�a<�a<d�a<��a<F�a<��a<)�a<��a<�a<|�a<�a<}�a<˜a<n�a<ѝa<F�a<Ğa<+�a<a<�a<��a<��a<h�a<ڡa<E�a<��a<
�a<��a<��a<a�a<Ƥa<�a<��a<ȥa<H�a<��a<�a<C�a<��a<�a<5�a<��a<Ũa<#�a<c�a<��a<�a<"�a<k�a<��a<۪a<�a<@�a<z�a<��a<�a<�a<9�a<R�a<��a<��a<��a<�a<�a<�a<*�a<P�a<[�a<n�a<��a<��a<��a<��a<̭a<Эa<��a<�a<̭a<׭a<ȭa<׭a<խa<ڭa<έa<��a<ƭa<��a<��a<��a<{�a<m�a<I�a<F�a<"�a<!�a<�a<�a<׬a<��a<��a<V�a<Y�a<�a<�a<ϫa<��a<p�a<8�a<"�a<Ъa<��a<��a<D�a<#�a<ʩa<��a<\�a<%�a<�a<��a<c�a<�a<ڧa<��a<L�a<��a<��a<e�a< �a<¥a<c�a<�a<��a<X�a<��a<��a<Z�a<Ӣa<��a<*�a<ơa<j�a<��a<��a<�a<a<W�a<�a<��a<�a<��a<#�a<�a<`�a<��a<��a<�a<��a<�a<ՙa<R�a<�a<��a<
�a<��a<?�a<�a<h�a<�a<��a<E�a<�a<��a<0�a<��a<v�a<�a<��a<u�a<�a<�a<u�a<F�a<�a<��a<z�a<�a<�a<��a<n�a<3�a<�a<юa<��a<��a<L�a<@�a<�a<��a<܍a<��a<��a<��a<~�a<b�a<i�a<c�a<i�a<c�a<Z�a<v�a<i�a<~�a<��a<��a<��a<��a<�  �  ݍa<�a<2�a<W�a<z�a<��a<Ҏa<�a<+�a<_�a<��a<�a<%�a<u�a<��a<��a<@�a<��a<ߑa<�a<t�a<ђa</�a<��a<�a<F�a<��a<�a<f�a<�a<>�a<��a<�a<t�a<�a<X�a<̘a<4�a<��a<�a<��a<�a<��a<�a<s�a<�a<[�a<ȝa<C�a<��a<"�a<��a<�a<��a< �a<m�a<աa<N�a<��a<(�a<��a<�a<P�a<��a<�a<��a<�a<?�a<��a<��a<Q�a<��a<�a<>�a<��a<Ҩa<�a<]�a<��a<�a<*�a<g�a<��a<تa<!�a<Q�a<y�a<��a<٫a<�a<*�a<I�a<g�a<��a<��a<�a<�a<�a<?�a<M�a<]�a<}�a<{�a<��a<��a<��a<��a<ʭa<Эa<ۭa<�a<ϭa<�a<�a<̭a<ڭa<��a<­a<��a<��a<��a<��a<z�a<y�a<l�a<8�a<:�a<�a<�a<�a<��a<��a<��a<U�a<.�a<�a<�a<ɫa<��a<]�a<P�a<�a<�a<��a<q�a<A�a<�a<ݩa<��a<f�a<(�a<�a<��a<[�a<1�a<٧a<��a<I�a<�a<��a<Z�a<�a<��a<l�a<�a<Ȥa<n�a<�a<��a<P�a<�a<��a<!�a<áa<Z�a<�a<��a<3�a<��a<]�a<�a<{�a<�a<��a<A�a<ʜa<M�a<�a<��a<�a<��a<7�a<̙a<f�a<��a<��a<,�a<��a<H�a<Ֆa<u�a<�a<��a<C�a<�a<��a<,�a<�a<s�a<-�a<Ғa<t�a<"�a<ӑa<��a<7�a<�a<��a<l�a<%�a<�a<��a<^�a<H�a<
�a<Ԏa<��a<r�a<J�a<-�a<�a<�a<֍a<��a<��a<��a<v�a<��a<w�a<Z�a<i�a<Q�a<b�a<`�a<p�a<n�a<��a<��a<��a<��a<�  �  ܍a<�a<�a<b�a<v�a<��a<�a<��a<^�a<e�a<��a<��a<�a<o�a<��a< �a<+�a<��a<ɑa<.�a<��a<Ēa<D�a<y�a<�a<H�a<��a<�a<V�a<וa< �a<��a<�a<��a<��a<?�a<�a<4�a<��a<�a<��a<��a<��a<��a<_�a<��a<P�a<ٝa<I�a<��a<N�a<��a<#�a<��a<��a<m�a<ءa<L�a<��a<.�a<v�a<�a<d�a<��a<.�a<u�a<�a</�a<��a<�a</�a<��a<էa<B�a<}�a<�a<�a<a�a<��a<ݩa<0�a<J�a<��a<��a<�a<;�a<u�a<��a<ǫa<�a< �a<m�a<��a<��a<ͬa<ͬa<
�a<�a<:�a<=�a<e�a<v�a<z�a<��a<��a<��a<��a<��a<߭a<��a<ޭa<Эa<ӭa<ʭa<ѭa<̭a<��a<ܭa<��a<ǭa<��a<��a<��a<Y�a<V�a<7�a<8�a<�a<�a<ݬa<��a<��a<t�a<��a<5�a<�a<��a<��a<��a<j�a<S�a<�a<��a<��a<��a<i�a<�a<�a<��a<m�a<*�a<بa<��a<K�a<!�a<��a<��a<9�a<��a<��a<A�a<$�a<��a<l�a<��a<��a<O�a<�a<��a<<�a<��a<��a<3�a<ɡa<e�a<�a<��a<7�a<��a<U�a<�a<~�a<�a<��a<G�a<��a<x�a<��a<��a< �a<��a<E�a<��a<W�a<�a<m�a<�a<��a<L�a<Җa<��a<��a<��a<S�a<ݔa<��a<�a<֓a<[�a<&�a<��a<p�a<,�a<a<��a<-�a<	�a<��a<V�a<3�a<Տa<��a<j�a<C�a<��a<܎a<��a<r�a<{�a<%�a<�a<�a<ʍa<ˍa<��a<��a<w�a<l�a<[�a<_�a<[�a<S�a<|�a<?�a<��a<u�a<��a<��a<��a<ʍa<�  �  ��a<�a<-�a<M�a<v�a<��a<a<��a<.�a<t�a<��a<�a<�a<`�a<��a<�a<9�a<��a<ؑa<)�a<q�a<͒a<�a<��a<��a<G�a<��a<�a<v�a<ҕa<I�a<��a<�a<s�a<�a<Y�a<Øa<3�a<��a<2�a<��a<�a<��a<�a<x�a<ۜa<\�a<˝a<4�a<��a<#�a<��a<�a<��a<�a<s�a<�a<A�a<��a<�a<��a<�a<K�a<��a<�a<��a<إa<F�a<��a<�a<B�a<��a<��a<A�a<{�a<ʨa<�a<b�a<��a<ީa</�a<r�a<��a<�a<�a<A�a<�a<��a<�a<��a<"�a<F�a<t�a<��a<��a<٬a<��a<�a</�a<?�a<e�a<u�a<��a<��a<��a<��a<ía<ía<ȭa<ܭa<ӭa<�a<ϭa<�a<�a<έa<��a<��a<��a<��a<��a<��a<��a<|�a<S�a<W�a<0�a<�a<��a<ެa<ͬa<��a<}�a<W�a<C�a<�a<��a<��a<��a<z�a<A�a<�a<�a<��a<�a<=�a<�a<̩a<��a<_�a<)�a<�a<��a<k�a<�a<�a<��a<9�a<�a<��a<Z�a<�a<��a<k�a<�a<ɤa<Z�a<�a<��a<U�a<�a<��a<%�a<��a<S�a<�a<��a<(�a<şa<N�a<��a<��a<�a<��a<5�a<̜a<S�a<�a<q�a<�a<��a<.�a<әa<S�a<�a<��a<%�a<��a<K�a<Жa<m�a<�a<��a<=�a<ݔa<��a<7�a<ӓa<{�a<*�a<a<z�a<�a<ݑa<w�a<.�a<�a<��a<f�a< �a<�a<��a<y�a<8�a<��a<܎a<��a<��a<J�a<)�a<��a<��a<ύa<��a<��a<��a<��a<i�a<x�a<p�a<]�a<S�a<a�a<k�a<t�a<s�a<��a<��a<Ía<Ǎa<�  �  �a<�a<G�a<J�a<v�a<��a<a<K�a<�a<p�a<��a<�a<7�a<_�a<��a<�a<^�a<��a<�a<�a<y�a<�a<�a<��a<ғa<K�a<��a<��a<k�a<��a<L�a<��a<"�a<�a<ݗa<k�a<��a<O�a<��a<�a<��a<��a<��a<ٛa<��a<؜a<s�a<ŝa<Y�a<�a<�a<��a<�a<��a<�a<e�a<סa<=�a<Ңa<�a<��a<ߣa<|�a<�a<�a<��a<ҥa<]�a<{�a<�a<0�a<��a<�a<.�a<��a<̨a<%�a<\�a<��a<��a<�a<l�a<��a<Ԫa<�a<A�a<��a<��a<�a<�a<h�a<Z�a<h�a<��a<��a<�a<�a<�a<-�a<Q�a<h�a<o�a<��a<|�a<�a<��a<��a<έa<ŭa<��a<��a<�a<ía<߭a<��a<ѭa<׭a<��a<ͭa<��a<��a<��a<i�a<}�a<B�a<I�a<�a<1�a<��a<ݬa<ʬa<��a<ˬa<H�a<?�a<�a<�a<ܫa<��a<r�a<6�a<8�a<ުa<��a<u�a<E�a<Y�a<��a<��a<Q�a<-�a<�a<��a<a�a<�a<�a<�a<V�a<��a<��a<m�a<��a<˥a<Z�a<��a<��a<F�a<	�a<��a<p�a<�a<��a<�a<١a<��a<�a<��a<!�a<ןa<J�a<�a<}�a<�a<ĝa<7�a<�a<J�a<�a<��a<�a<Úa<)�a<�a<@�a<�a<n�a<�a<��a<8�a<�a<o�a<�a<��a<G�a<��a<{�a<1�a<��a<o�a<�a<a<��a<�a<�a<k�a<t�a<��a<��a<x�a<#�a<
�a<��a<s�a<6�a<�a<ߎa<��a<��a<;�a<y�a<	�a<�a<ڍa<��a<ȍa<m�a<��a<]�a<p�a<H�a<`�a<m�a<G�a<}�a<R�a<��a<��a<��a<ča<��a<�  �  ��a<�a<-�a<M�a<v�a<��a<a<��a<.�a<t�a<��a<�a<�a<`�a<��a<�a<9�a<��a<ؑa<)�a<q�a<͒a<�a<��a<��a<G�a<��a<�a<v�a<ҕa<I�a<��a<�a<s�a<�a<Y�a<Øa<3�a<��a<2�a<��a<�a<��a<�a<x�a<ۜa<\�a<˝a<4�a<��a<#�a<��a<�a<��a<�a<s�a<�a<A�a<��a<�a<��a<�a<K�a<��a<�a<��a<إa<F�a<��a<�a<B�a<��a<��a<A�a<{�a<ʨa<�a<b�a<��a<ީa</�a<r�a<��a<�a<�a<A�a<�a<��a<�a<��a<"�a<F�a<t�a<��a<��a<٬a<��a<�a</�a<?�a<e�a<u�a<��a<��a<��a<��a<ía<ía<ȭa<ܭa<ӭa<�a<ϭa<�a<�a<έa<��a<��a<��a<��a<��a<��a<��a<|�a<S�a<W�a<0�a<�a<��a<ެa<ͬa<��a<}�a<W�a<C�a<�a<��a<��a<��a<z�a<A�a<�a<�a<��a<�a<=�a<�a<̩a<��a<_�a<)�a<�a<��a<k�a<�a<�a<��a<9�a<�a<��a<Z�a<�a<��a<k�a<�a<ɤa<Z�a<�a<��a<U�a<�a<��a<%�a<��a<S�a<�a<��a<(�a<şa<N�a<��a<��a<�a<��a<5�a<̜a<S�a<�a<q�a<�a<��a<.�a<әa<S�a<�a<��a<%�a<��a<K�a<Жa<m�a<�a<��a<=�a<ݔa<��a<7�a<ӓa<{�a<*�a<a<z�a<�a<ݑa<w�a<.�a<�a<��a<f�a< �a<�a<��a<y�a<8�a<��a<܎a<��a<��a<J�a<)�a<��a<��a<ύa<��a<��a<��a<��a<i�a<x�a<p�a<]�a<S�a<a�a<k�a<t�a<s�a<��a<��a<Ía<Ǎa<�  �  ܍a<�a<�a<b�a<v�a<��a<�a<��a<^�a<e�a<��a<��a<�a<o�a<��a< �a<+�a<��a<ɑa<.�a<��a<Ēa<D�a<y�a<�a<H�a<��a<�a<V�a<וa< �a<��a<�a<��a<��a<?�a<�a<4�a<��a<�a<��a<��a<��a<��a<_�a<��a<P�a<ٝa<I�a<��a<N�a<��a<#�a<��a<��a<m�a<ءa<L�a<��a<.�a<v�a<�a<d�a<��a<.�a<u�a<�a</�a<��a<�a</�a<��a<էa<B�a<}�a<�a<�a<a�a<��a<ݩa<0�a<J�a<��a<��a<�a<;�a<u�a<��a<ǫa<�a< �a<m�a<��a<��a<ͬa<ͬa<
�a<�a<:�a<=�a<e�a<v�a<z�a<��a<��a<��a<��a<��a<߭a<��a<ޭa<Эa<ӭa<ʭa<ѭa<̭a<��a<ܭa<��a<ǭa<��a<��a<��a<Y�a<V�a<7�a<8�a<�a<�a<ݬa<��a<��a<t�a<��a<5�a<�a<��a<��a<��a<j�a<S�a<�a<��a<��a<��a<i�a<�a<�a<��a<m�a<*�a<بa<��a<K�a<!�a<��a<��a<9�a<��a<��a<A�a<$�a<��a<l�a<��a<��a<O�a<�a<��a<<�a<��a<��a<3�a<ɡa<e�a<�a<��a<7�a<��a<U�a<�a<~�a<�a<��a<G�a<��a<x�a<��a<��a< �a<��a<E�a<��a<W�a<�a<m�a<�a<��a<L�a<Җa<��a<��a<��a<S�a<ݔa<��a<�a<֓a<[�a<&�a<��a<p�a<,�a<a<��a<-�a<	�a<��a<V�a<3�a<Տa<��a<j�a<C�a<��a<܎a<��a<r�a<{�a<%�a<�a<�a<ʍa<ˍa<��a<��a<w�a<l�a<[�a<_�a<[�a<S�a<|�a<?�a<��a<u�a<��a<��a<��a<ʍa<�  �  ݍa<�a<2�a<W�a<z�a<��a<Ҏa<�a<+�a<_�a<��a<�a<%�a<u�a<��a<��a<@�a<��a<ߑa<�a<t�a<ђa</�a<��a<�a<F�a<��a<�a<f�a<�a<>�a<��a<�a<t�a<�a<X�a<̘a<4�a<��a<�a<��a<�a<��a<�a<s�a<�a<[�a<ȝa<C�a<��a<"�a<��a<�a<��a< �a<m�a<աa<N�a<��a<(�a<��a<�a<P�a<��a<�a<��a<�a<?�a<��a<��a<Q�a<��a<�a<>�a<��a<Ҩa<�a<]�a<��a<�a<*�a<g�a<��a<تa<!�a<Q�a<y�a<��a<٫a<�a<*�a<I�a<g�a<��a<��a<�a<�a<�a<?�a<M�a<]�a<}�a<{�a<��a<��a<��a<��a<ʭa<Эa<ۭa<�a<ϭa<�a<�a<̭a<ڭa<��a<­a<��a<��a<��a<��a<z�a<y�a<l�a<8�a<:�a<�a<�a<�a<��a<��a<��a<U�a<.�a<�a<�a<ɫa<��a<]�a<P�a<�a<�a<��a<q�a<A�a<�a<ݩa<��a<f�a<(�a<�a<��a<[�a<1�a<٧a<��a<I�a<�a<��a<Z�a<�a<��a<l�a<�a<Ȥa<n�a<�a<��a<P�a<�a<��a<!�a<áa<Z�a<�a<��a<3�a<��a<]�a<�a<{�a<�a<��a<A�a<ʜa<M�a<�a<��a<�a<��a<7�a<̙a<f�a<��a<��a<,�a<��a<H�a<Ֆa<u�a<�a<��a<C�a<�a<��a<,�a<�a<s�a<-�a<Ғa<t�a<"�a<ӑa<��a<7�a<�a<��a<l�a<%�a<�a<��a<^�a<H�a<
�a<Ԏa<��a<r�a<J�a<-�a<�a<�a<֍a<��a<��a<��a<v�a<��a<w�a<Z�a<i�a<Q�a<b�a<`�a<p�a<n�a<��a<��a<��a<��a<�  �  �a<��a<6�a<D�a<}�a<��a<a<�a<,�a<��a<��a<ޏa<*�a<]�a<��a<�a<H�a<s�a<�a<=�a<x�a<�a<�a<��a<ݓa<C�a<��a<��a<n�a<a<?�a<��a<�a<{�a<�a<d�a<��a<F�a<��a<)�a<��a<�a<|�a<�a<}�a<˜a<n�a<ѝa<F�a<Ğa<+�a<a<�a<��a<��a<h�a<ڡa<E�a<��a<
�a<��a<��a<a�a<Ƥa<�a<��a<ȥa<H�a<��a<�a<C�a<��a<�a<5�a<��a<Ũa<#�a<c�a<��a<�a<"�a<k�a<��a<۪a<�a<@�a<z�a<��a<�a<�a<9�a<R�a<��a<��a<��a<�a<�a<�a<*�a<P�a<[�a<n�a<��a<��a<��a<��a<̭a<Эa<��a<�a<̭a<׭a<ȭa<׭a<խa<ڭa<έa<��a<ƭa<��a<��a<��a<{�a<m�a<I�a<F�a<"�a<!�a<�a<�a<׬a<��a<��a<V�a<Y�a<�a<�a<ϫa<��a<p�a<8�a<"�a<Ъa<��a<��a<D�a<#�a<ʩa<��a<\�a<%�a<�a<��a<c�a<�a<ڧa<��a<L�a<��a<��a<e�a< �a<¥a<c�a<�a<��a<X�a<��a<��a<Z�a<Ӣa<��a<*�a<ơa<j�a<��a<��a<�a<a<W�a<�a<��a<�a<��a<#�a<�a<`�a<��a<��a<�a<��a<�a<ՙa<R�a<�a<��a<
�a<��a<?�a<�a<h�a<�a<��a<E�a<�a<��a<0�a<��a<v�a<�a<��a<u�a<�a<�a<u�a<F�a<�a<��a<z�a<�a<�a<��a<n�a<3�a<�a<юa<��a<��a<L�a<@�a<�a<��a<܍a<��a<��a<��a<~�a<b�a<i�a<c�a<i�a<c�a<Z�a<v�a<i�a<~�a<��a<��a<��a<��a<�  �  ��a<��a<3�a<]�a<m�a<��a<Ԏa<
�a<3�a<h�a<��a<�a<'�a<Z�a<��a<�a<E�a<��a<��a<$�a<~�a<ےa<,�a<��a<ۓa<P�a<��a< �a<w�a<ەa<?�a<��a<�a<��a<�a<F�a<ݘa<F�a<��a<%�a<��a<�a<��a<�a<t�a<�a<Y�a<Нa<F�a<��a<.�a<��a<�a<��a<��a<h�a<ޡa<A�a<��a<�a<}�a<�a<\�a<��a<#�a<��a<ޥa<B�a<��a<�a<I�a<��a<�a<)�a<��a<�a<�a<_�a<��a<�a<�a<f�a<��a<�a<�a<E�a<��a<��a<ԫa<�a<.�a<U�a<v�a<��a<Ǭa<�a<�a<+�a<)�a<L�a<o�a<_�a<}�a<��a<��a<��a<��a<��a<حa<ݭa<ʭa<�a<حa<ޭa<ԭa<��a<ѭa<έa<��a<��a<��a<|�a<�a<q�a<[�a<R�a<!�a<�a<�a<Ԭa<��a<��a<��a<]�a<7�a<��a< �a<˫a<��a<��a<4�a<�a<��a<��a<z�a<J�a<�a<کa<��a<Z�a<2�a<�a<��a<m�a<%�a<ڧa<��a<7�a<�a<��a<H�a<�a<¥a<P�a<�a<��a<b�a<	�a<��a<Q�a<�a<��a<*�a<ơa<e�a<��a<��a<!�a<͟a<R�a<�a<��a<�a<��a<6�a<��a<^�a<�a<��a<�a<��a<5�a<Ιa<X�a<�a<��a<�a<��a<3�a<�a<��a<�a<��a<Y�a<�a<�a<+�a<ӓa<}�a<�a<ƒa<|�a<�a<ϑa<��a<;�a<�a<��a<O�a<-�a<�a<��a<��a<2�a<
�a<�a<��a<t�a<Q�a<6�a<�a<�a<ɍa<Ía<��a<��a<��a<r�a<o�a<a�a<I�a<f�a<n�a<M�a<z�a<��a<y�a<��a<��a<΍a<�  �  �a<�a<%�a<R�a<w�a<��a<ߎa<��a<<�a<r�a<��a<ۏa<�a<l�a<��a<��a<&�a<��a<ؑa<2�a<|�a<̒a<8�a<��a<�a<>�a<��a<�a<b�a<��a<:�a<��a<�a<r�a<�a<\�a<͘a<)�a<��a<"�a<��a<�a<|�a<�a<c�a<�a<O�a<۝a<F�a<��a<=�a<��a< �a<y�a<��a<n�a<ܡa<F�a<��a<'�a<��a<��a<N�a<��a</�a<u�a<�a<1�a<��a<�a<=�a<��a<�a<B�a<u�a<Ҩa<�a<g�a<��a<۩a<4�a<c�a<��a<Ϊa<�a<M�a<o�a<��a<̫a<�a<$�a<O�a<��a<��a<Ĭa<Ǭa<��a<�a<6�a<:�a<T�a<}�a<��a<��a<��a<��a<��a<­a<խa<ͭa<�a<ҭa<ڭa<�a<׭a<ҭa<��a<ǭa<��a<��a<��a<��a<��a<u�a<^�a<=�a<<�a<�a<��a<ެa<��a<��a<y�a<f�a<A�a<�a<�a<��a<��a<r�a<G�a< �a<�a<��a<��a<H�a<�a<�a<��a<m�a< �a<�a<��a<X�a<*�a<էa<��a<:�a<�a<��a<]�a<�a<��a<m�a<�a<äa<Z�a<��a<��a<@�a<��a<��a<4�a<ǡa<T�a<�a<��a<4�a<��a<R�a<�a<��a<�a<��a<@�a<Ɯa<j�a<�a<~�a<!�a<��a<D�a<��a<k�a<�a<{�a<$�a<��a<L�a<ʖa<u�a<�a<��a<C�a<۔a<��a<(�a<ޓa<i�a<!�a<Βa<i�a<,�a<Ǒa<��a<0�a<�a<��a<d�a<*�a<Ϗa<��a<q�a<?�a<��a<ˎa<��a<|�a<_�a<&�a<�a<�a<΍a<��a<��a<��a<y�a<s�a<r�a<e�a<a�a<K�a<g�a<i�a<y�a<m�a<��a<��a<��a<ҍa<�  �  �a<�a<&�a<E�a<��a<��a<Ǝa<�a<8�a<o�a<��a<Џa<+�a<k�a<��a<��a<A�a<p�a<Ցa<.�a<{�a<ߒa<!�a<��a<�a<<�a<��a<�a<s�a<ѕa<3�a<��a<!�a<��a<�a<m�a<Řa<M�a<��a<�a<��a<�a<��a<��a<n�a<ޜa<a�a<ϝa<?�a<��a<1�a<��a<	�a<��a<
�a<d�a<ϡa<Y�a<��a<�a<��a<�a<\�a<��a<�a<��a<ܥa<=�a<��a<�a<I�a<��a<ݧa<<�a<��a<ͨa<%�a<_�a<��a<��a<�a<\�a<��a<�a<�a<D�a<t�a<��a<ݫa<��a<2�a<S�a<|�a<��a<��a<�a<
�a<��a<4�a<R�a<O�a<n�a<��a<��a<��a<��a<��a<ԭa<ía<έa<׭a<�a<٭a<ӭa<��a<�a<ҭa<��a<ͭa<��a<��a<��a<g�a<j�a<Y�a<N�a<1�a<�a<�a<�a<Ȭa<��a<��a<b�a<>�a<�a<ܫa<Ыa<��a<W�a<P�a<�a<ͪa<��a<��a<H�a<�a<Ωa<��a<l�a<�a<ߨa<��a<h�a<�a<Χa<�a<U�a<��a<��a<o�a<�a<ɥa<m�a<��a<��a<c�a<�a<��a<K�a<�a<��a<(�a<��a<f�a<��a<��a<�a<��a<g�a<�a<u�a<%�a<��a<(�a<ʜa<]�a<�a<{�a<�a<��a<3�a<ʙa<_�a<�a<��a<�a<��a<F�a<�a<p�a<�a<��a<H�a<��a<�a<!�a<Γa<z�a< �a<Œa<n�a<%�a<ؑa<{�a<?�a<�a<��a<d�a<�a<�a<��a<X�a<=�a<�a<Ǝa<��a<�a<[�a<=�a<�a<�a<��a<��a<��a<��a<��a<s�a<e�a<K�a<r�a<g�a<R�a<}�a<d�a<��a<��a<��a<��a<̍a<�  �  ��a<��a<A�a<Q�a<q�a<��a<Ďa<�a<$�a<m�a<��a<�a< �a<^�a<��a<�a<A�a<��a<ؑa<'�a<m�a<Вa<!�a<��a<̓a<Q�a<��a<�a<|�a<˕a<[�a<��a<�a<��a<�a<[�a<Ęa<J�a<��a<<�a<��a<�a<��a<�a<��a<Ӝa<_�a<ȝa<:�a<��a<�a<��a<�a<��a<�a<l�a<ޡa<:�a<��a<�a<��a<�a<W�a<��a<�a<��a<ɥa<V�a<��a<��a<L�a<��a<�a<%�a<��a<Ϩa<�a<`�a<��a<�a<�a<��a<��a<�a<�a<J�a<��a<��a<�a<��a<&�a<G�a<r�a<��a<��a<�a<�a<!�a<.�a<E�a<f�a<i�a<��a<��a<��a<��a<��a<ĭa<ɭa<�a<ƭa<�a<ӭa<�a<�a<��a<խa<��a<��a<��a<��a<��a<��a<��a<Q�a<X�a<�a<+�a<��a<جa<ʬa<��a<��a<N�a<<�a<�a<��a<ūa<��a<~�a<:�a<�a<�a<��a<}�a<9�a<�a<Ωa<��a<K�a<3�a<�a<��a<q�a<�a<��a<��a<B�a<�a<��a<\�a<�a<ƥa<M�a<(�a<Ƥa<b�a<�a<��a<f�a<ڢa<��a<!�a<��a<`�a<�a<��a<%�a<ȟa<N�a<�a<��a<�a<��a<2�a<Ҝa<L�a<�a<x�a<�a<��a< �a<�a<R�a<��a<��a<�a<ʗa</�a<�a<r�a<�a<��a<L�a<�a<y�a<J�a<ɓa<��a<�a<˒a<��a<�a<�a<y�a<3�a<�a<��a<h�a<$�a<�a<��a<z�a<8�a<�a<ݎa<��a<~�a<B�a<1�a<��a<�a<Ѝa<��a<��a<�a<��a<m�a<��a<o�a<O�a<k�a<W�a<g�a<j�a<��a<��a<��a<Ѝa<ōa<�  �  �a<�a<)�a<Q�a<��a<��a<ߎa<��a<H�a<v�a<��a<�a<�a<d�a<��a<�a<-�a<��a<͑a<6�a<��a<̒a<6�a<��a<�a<I�a<��a<	�a<j�a<ɕa<2�a<��a<�a<��a<��a<K�a<Ԙa<C�a<��a<*�a<��a<�a<��a<��a<p�a<�a<[�a<۝a<U�a<��a<G�a<��a<�a<��a<��a<e�a<աa<D�a<��a<#�a<��a<�a<b�a<̤a<*�a<��a<�a<>�a<��a<�a<<�a<��a<�a<B�a<��a<ڨa<�a<j�a<��a<�a<2�a<`�a<��a<ժa<�a<A�a<{�a<��a<۫a<�a<*�a<b�a<��a<��a<Ƭa<Ѭa<��a<�a<.�a<=�a<f�a<q�a<��a<��a<��a<��a<ŭa<ɭa<έa<ѭa<ۭa<׭a<Эa<˭a<ݭa<ѭa<έa<Эa<��a<��a<��a<��a<��a<`�a<N�a<E�a<0�a<�a<��a<�a<ɬa<��a<w�a<r�a<E�a<�a<��a<��a<��a<j�a<D�a<�a<�a<��a<��a<\�a<�a<�a<��a<d�a<+�a<�a<��a<_�a<�a<ͧa<��a<C�a<��a<��a<M�a<�a<��a<j�a<�a<��a<U�a<�a<��a<M�a<�a<��a<4�a<աa<b�a<�a<��a<,�a<��a<Q�a<�a<{�a<�a<��a<;�a<ɜa<r�a<��a<��a<�a<��a<7�a<˙a<R�a<�a<z�a<�a<��a<L�a<�a<}�a<�a<��a<P�a<�a<��a<%�a<Óa<p�a<�a<a<v�a<�a<֑a<��a<6�a<��a<��a<[�a<,�a<ُa<��a<l�a<7�a<��a<ݎa<��a<��a<g�a<'�a<�a<��a<Սa<��a<��a<��a<~�a<j�a<\�a<j�a<`�a<d�a<q�a<T�a<��a<��a<��a<��a<��a<a<�  �  ܍a<�a<%�a<R�a<��a<��a<ێa<�a<3�a<V�a<��a<ُa<�a<}�a<��a<
�a</�a<��a<Αa<�a<u�a<̒a<1�a<u�a<��a<;�a<��a<�a<d�a<��a</�a<��a<�a<u�a<��a<W�a<ژa</�a<��a<�a<��a<$�a<{�a<�a<_�a<�a<T�a<ŝa<N�a<��a<4�a<��a<�a<|�a<�a<d�a<ʡa<[�a<��a<)�a<q�a<��a<?�a<¤a<�a<v�a<�a</�a<��a<�a<U�a<��a<ڧa<K�a<z�a<ۨa<�a<i�a<��a<�a<4�a<U�a<Īa<۪a<�a<M�a<n�a<��a<ūa<�a<(�a<E�a<q�a<��a<��a<Ҭa<�a<��a<?�a<H�a<T�a<v�a<j�a<��a<��a<��a<��a<έa<խa<ǭa<�a<ɭa<��a<ڭa<ɭa<�a<��a<ϭa<��a<��a<��a<��a<y�a<j�a<��a<7�a<C�a<�a<��a<�a<��a<��a<q�a<]�a<%�a<�a<�a<��a<��a<I�a<]�a<�a<�a<��a<r�a<A�a<�a<ߩa<��a<t�a<�a<�a<��a<Y�a<C�a<˧a<��a<J�a<�a<��a<X�a<�a<��a<v�a<�a<ˤa<v�a<��a<��a<<�a<��a<��a<�a<Ρa<G�a< �a<v�a<2�a<��a<d�a<�a<p�a<&�a<��a<B�a<��a<_�a<՛a<��a<�a<��a<D�a<��a<l�a<�a<��a<2�a<��a<U�a<ϖa<~�a<�a<��a<D�a<�a<��a<�a<�a<u�a<#�a<Βa<i�a<1�a<��a<��a<4�a<�a<��a<S�a<'�a<ڏa<��a<O�a<H�a<�a<ʎa<��a<b�a<V�a<�a<�a<ݍa<ۍa<��a<��a<��a<p�a<��a<l�a<V�a<p�a<N�a<p�a<`�a<|�a<m�a<��a<��a<��a<��a<�  �  �a<��a<6�a<N�a<w�a<��a<Ԏa<�a</�a<z�a<��a<؏a<�a<h�a<��a<�a<0�a<��a<�a<9�a<r�a<�a<&�a<��a<ݓa<A�a<��a<��a<d�a<ɕa<D�a<��a<�a<u�a<�a<f�a<ɘa<9�a<��a<%�a<��a< �a<y�a<�a<{�a<ޜa<d�a<ʝa<U�a<��a<4�a<��a<�a<}�a<�a<i�a<סa<>�a<��a<&�a<��a<��a<W�a<Ѥa<�a<��a<٥a<F�a<��a<�a<7�a<��a<�a<8�a<��a<Ψa<'�a<j�a<��a<�a<'�a<j�a<��a<Ϫa<��a<C�a<x�a<��a<�a<��a<@�a<J�a<��a<��a<��a<Ҭa<�a<�a<2�a<>�a<Q�a<x�a<��a<��a<��a<��a<��a<ȭa<˭a<ޭa<ʭa<ԭa<ϭa<ۭa<֭a<ҭa<ȭa<��a<��a<��a<��a<��a<��a<s�a<R�a<@�a< �a< �a<��a<ެa<¬a<��a<��a<Y�a<I�a< �a<�a<��a<��a<s�a<@�a<
�a<�a<��a<��a<?�a<&�a<ԩa<��a<\�a<#�a<�a<��a<Z�a<�a<ߧa<��a<L�a<�a<��a<g�a<	�a<��a<b�a<�a<��a<S�a<��a<��a<X�a<�a<��a<#�a<աa<d�a<��a<��a<2�a<��a<J�a<�a<}�a<	�a<��a<?�a<לa<g�a<�a<��a<�a<��a<0�a<әa<T�a<�a<u�a<�a<��a<B�a<ؖa<p�a<�a<��a<@�a<�a<��a</�a<œa<j�a<
�a<Ēa<s�a<�a<ۑa<{�a<L�a<�a<��a<r�a<'�a<ڏa<��a<n�a<<�a<��a<Ȏa<��a<��a<Q�a<;�a<�a<�a<ԍa<��a<��a<��a<{�a<h�a<l�a<d�a<b�a<]�a<_�a<p�a<m�a<y�a<��a<��a<��a<ōa<�  �  m�a<��a<Ďa<ӎa<�a<&�a<=�a<��a<��a<��a<�a<e�a<��a<͐a<$�a<a�a<��a<�a<M�a<��a<�a<_�a<��a<�a<\�a<Ĕa<2�a<t�a<�a<7�a<ǖa<�a<��a<�a<\�a<טa<:�a<̙a<�a<��a<�a<q�a<��a<f�a<�a<E�a<ӝa<,�a<��a<*�a<��a<�a<p�a<�a<b�a<��a<-�a<��a<�a<|�a<�a<\�a<��a<�a<m�a<�a<0�a<��a<��a<N�a<��a<�a<[�a<��a<�a<1�a<~�a<éa<�a<Y�a<x�a<٪a<�a<7�a<h�a<��a<�a<��a<8�a<I�a<��a<��a<�a<��a<�a<C�a<T�a<q�a<y�a<��a<��a<ĭa<��a<�a<
�a< �a<�a</�a<*�a<M�a<3�a<8�a<%�a<J�a<=�a<&�a<F�a<�a<!�a<��a<�a<�a<�a<�a<��a<��a<��a<��a<^�a<L�a<%�a<�a<�a<��a<��a<k�a<S�a<8�a<�a<Ϋa<��a<}�a<G�a<�a<�a<��a<��a<"�a<�a<©a<��a<Z�a<��a<ƨa<j�a<L�a<�a<��a<n�a<�a<Ŧa<g�a<6�a<��a<��a<�a<��a<j�a<�a<ģa<C�a<��a<~�a<$�a<ˡa<c�a<��a<��a<*�a<��a<C�a<מa<z�a<�a<��a<6�a<Ҝa<_�a<�a<m�a<�a<��a<J�a<Йa<b�a<�a<��a<3�a<��a<m�a<�a<��a<%�a<Εa<s�a<�a<��a<7�a<�a<��a<P�a<��a<��a<Q�a<�a<a<l�a<3�a<ߐa<��a<k�a<"�a<�a<��a<��a<W�a<�a<�a<̎a<��a<}�a<n�a<\�a<8�a<>�a<�a< �a<��a<��a<�a<׍a<��a<ٍa<�a<�a<�a<�a<$�a<H�a<?�a<�  �  f�a<��a<��a<Ύa<��a<,�a<g�a<��a<��a<�a<(�a<h�a<��a<�a<4�a<w�a<��a<�a<N�a<��a<��a<W�a<��a<	�a<d�a<��a<$�a<�a<�a<U�a<��a<�a<��a<��a<c�a<՘a<>�a<��a< �a<��a<�a<��a<�a<h�a<לa<N�a<͝a<C�a<��a<#�a<��a<��a<��a<�a<]�a<ܡa<I�a<��a<�a<��a<ޣa<^�a<��a<-�a<��a<�a<<�a<��a<��a<J�a<��a<�a<N�a<��a<�a</�a<|�a<éa<�a<B�a<��a<ͪa<�a<;�a<n�a<��a<Ϋa<
�a<<�a<m�a<��a<��a<ܬa<�a<&�a<2�a<`�a<��a<��a<��a<��a<֭a<ޭa<��a<�a<%�a<&�a<'�a<,�a<4�a<;�a<4�a<E�a<C�a<:�a<.�a<'�a<%�a<$�a<�a< �a<�a<�a<׭a<ȭa<��a<��a<y�a<Y�a<C�a<+�a<�a<�a<ìa<��a<y�a<V�a<&�a<�a<ޫa<��a<m�a<M�a<�a<�a<��a<{�a<J�a<�a<ʩa<~�a<L�a<�a<Ĩa<��a<A�a<�a<��a<\�a<�a<æa<k�a<�a<ťa<t�a<&�a<ͤa<c�a<�a<��a<L�a<��a<��a<:�a<ġa<h�a<�a<��a<!�a<��a<`�a<�a<|�a<�a<��a<(�a<Ӝa<X�a<��a<��a<�a<��a<3�a<Ιa<]�a<��a<��a<&�a<��a<O�a<�a<��a<&�a<��a<\�a< �a<��a<Q�a<�a<��a<F�a<�a<��a<U�a<�a<��a<i�a<,�a<ِa<��a<Z�a<.�a<��a<ďa<��a<V�a<,�a<��a<׎a<��a<��a<y�a<U�a<9�a<%�a<�a<��a<�a<��a<�a<ލa<ލa<�a<��a<��a<��a<�a<%�a<?�a<\�a<�  �  _�a<��a<��a<��a<��a<�a<\�a<w�a<ҏa<�a<,�a<p�a<��a<�a<�a<{�a<��a<�a<K�a<��a<
�a<F�a<��a<�a<s�a<��a<&�a<��a<ܕa<]�a<��a<+�a<��a<��a<p�a<Șa<U�a<��a<?�a<��a<�a<��a<�a<~�a<Ӝa<i�a<��a<0�a<��a<�a<��a<�a<��a<�a<`�a<͡a<7�a<��a<�a<��a<գa<k�a<��a<�a<{�a<եa<V�a<��a<�a<S�a<��a< �a<=�a<��a<�a<E�a<u�a<ũa<�a<I�a<��a<��a<�a<4�a<��a<��a<իa<�a<"�a<e�a<��a<��a<ެa<�a<1�a<1�a<c�a<b�a<��a<��a<ŭa<�a<٭a<�a<��a<�a<�a<'�a<C�a<)�a<R�a<.�a<M�a<-�a<9�a<B�a<$�a<<�a<�a<(�a<��a<��a<�a<��a<ϭa<��a<��a<r�a<k�a<F�a<�a<�a<׬a<ݬa<��a<}�a<^�a<!�a<�a<��a<��a<m�a<Y�a<
�a<ߪa<��a<j�a<B�a<�a<ةa<��a<O�a<�a<��a<��a<'�a<��a<��a<c�a<�a<��a<��a<�a<�a<h�a<�a<Ѥa<c�a<#�a<��a<g�a<�a<��a<+�a<��a<y�a<�a<��a<%�a<��a<Q�a<�a<~�a<�a<��a<�a<��a<W�a<�a<{�a<�a<��a<3�a<�a<f�a<��a<��a<�a<՗a<Q�a< �a<��a<(�a<Εa<c�a<�a<��a<W�a<�a<��a<Q�a<�a<��a<;�a<�a<��a<v�a<.�a<אa<��a<Y�a<1�a<ۏa<��a<��a<]�a<6�a<�a<�a<��a<��a<_�a<U�a<P�a<�a<,�a<��a<	�a<��a<�a<�a<ۍa<��a<ݍa<�a<��a<�a<)�a<(�a<c�a<�  �  l�a<��a<��a<ώa<��a<)�a<Y�a<��a<��a<��a<�a<a�a<��a<�a<0�a<y�a<��a<�a<Q�a<��a<��a<T�a<��a<
�a<_�a<��a<�a<��a<�a<Q�a<��a<$�a<��a<�a<j�a<јa<D�a<��a<$�a<��a<�a<|�a<��a<j�a<ٜa<N�a<ѝa<9�a<��a<�a<��a<�a<y�a<�a<h�a<ϡa<@�a<��a<�a<�a<�a<P�a<��a<�a<}�a<�a<=�a<��a<��a<S�a<��a<��a<Q�a<��a<�a<2�a<{�a<ũa<��a<C�a<��a<˪a<�a<2�a<r�a<��a<ӫa<�a<=�a<_�a<��a<��a<֬a<��a<�a<<�a<e�a<|�a<��a<��a<��a<ǭa<�a<�a<�a<�a<�a<+�a<*�a<*�a<>�a<;�a<:�a<=�a<E�a<0�a<!�a<,�a<�a<�a<��a<�a<�a<׭a<��a<��a<��a<o�a<[�a<D�a<(�a<�a<�a<��a<��a<k�a<O�a<1�a<�a<ګa<��a<w�a<E�a<�a<�a<��a<x�a<;�a<�a<ĩa<��a<<�a<�a<��a<��a<>�a<��a<��a<O�a<�a<��a<r�a<�a<ɥa<|�a<�a<��a<k�a<�a<��a<L�a<��a<��a<*�a<��a<\�a<��a<��a<(�a<ǟa<S�a<�a<��a<�a<��a<8�a<Ŝa<Q�a<�a<~�a<�a<��a<9�a<͙a<f�a<�a<��a<*�a<��a<N�a<�a<��a<(�a<��a<]�a<�a<��a<N�a<�a<��a<<�a<�a<��a<V�a< �a<��a<h�a<&�a<�a<��a<d�a<3�a<��a<��a<��a<T�a<�a<�a<юa<��a<��a<r�a<Y�a<7�a<�a<�a<�a<��a<��a<�a<��a<؍a<�a<ߍa<��a<�a<�a</�a<?�a<Q�a<�  �  ��a<}�a<��a<Վa<��a<1�a<J�a<��a<��a<�a<(�a<b�a<��a<Րa<>�a<Z�a<��a<��a<^�a<��a<�a<e�a<��a<�a<Q�a<ϔa< �a<}�a<��a<D�a<��a<�a<��a<�a<f�a<�a<:�a<��a<�a<��a<�a<��a<�a<W�a<�a<B�a<՝a<9�a<��a<.�a<��a<$�a<t�a<�a<R�a<ѡa<F�a<��a<�a<v�a<�a<E�a<��a<%�a<y�a<��a<.�a<��a<�a<Z�a<��a<�a<O�a<��a<�a<)�a<��a<ȩa<��a<Q�a<z�a<Ҫa<��a<I�a<q�a<��a<�a<��a<M�a<O�a<��a<��a<٬a<	�a<�a<>�a<G�a<��a<��a<��a<��a<ϭa<��a<ݭa<�a<�a<$�a<#�a<*�a<K�a<'�a<P�a<7�a<;�a<0�a<0�a<0�a<"�a<2�a<�a<�a<��a<׭a<حa<��a<��a<��a<��a<`�a<7�a<0�a<��a<��a<��a<��a<y�a<P�a<%�a<�a<�a<��a<t�a<=�a<�a<�a<��a<��a<)�a<�a<��a<��a<I�a<�a<֨a<v�a<C�a<�a<��a<V�a<�a<Ӧa<h�a<&�a<��a<u�a<�a<Ĥa<z�a<��a<ƣa<@�a<��a<��a<.�a<Сa<K�a<�a<��a<*�a<��a<U�a<�a<k�a<�a<��a<N�a<��a<_�a<��a<y�a<)�a<��a<P�a<��a<m�a<��a<��a<'�a<��a<^�a<�a<��a<+�a<��a<k�a<��a<��a<A�a< �a<��a<<�a<�a<��a<g�a<�a<őa<g�a<(�a<�a<��a<f�a<�a<�a<��a<�a<V�a<%�a<�a<��a<ǎa<��a<w�a<Q�a<7�a<=�a<�a<�a<�a<�a<ߍa<�a<�a<�a<�a<��a<�a<�a<�a<@�a<K�a<�  �  k�a<��a<��a<ݎa<��a<-�a<K�a<��a<��a<�a<*�a<l�a<��a<�a<�a<o�a<Ƒa<�a<P�a<��a<��a<b�a<��a<�a<a�a<Δa<�a<��a<�a<J�a<��a<#�a<��a<��a<X�a<Ęa<D�a<��a<4�a<��a<�a<}�a<��a<_�a<�a<[�a<͝a<>�a<��a</�a<��a<
�a<��a<��a<^�a<Ρa<:�a<��a<"�a<��a<�a<X�a<Ǥa<)�a<��a<�a<G�a<��a<�a<Q�a<��a<��a<H�a<��a<�a<6�a<p�a<��a<�a<S�a<��a<Ǫa<��a<8�a<s�a<��a<�a<	�a<8�a<]�a<��a<��a<جa<��a<&�a<I�a<\�a<o�a<��a<��a<ʭa<׭a<߭a<��a<�a<�a<%�a<-�a<7�a<?�a</�a<8�a<;�a<B�a<2�a<A�a<+�a<#�a<�a<�a<�a<�a<�a<حa<��a<��a<��a<~�a<h�a<F�a<,�a<��a<�a<Ĭa<��a<{�a<Z�a</�a<�a<ȫa<��a<��a<P�a<�a<ݪa<��a<��a<5�a<�a<Ʃa<��a<G�a<
�a<¨a<|�a<?�a<��a<��a<d�a<�a<��a<q�a<�a<٥a<p�a< �a<��a<k�a<�a<��a<Y�a<��a<��a<1�a<Сa<b�a<��a<��a<2�a<��a<R�a<�a<{�a<�a<��a<6�a<Μa<i�a<��a<��a<�a<��a<>�a<Ǚa<d�a<��a<��a<!�a<ȗa<V�a<�a<}�a<�a<ʕa<m�a<
�a<��a<F�a<�a<��a<?�a<��a<��a<Q�a<��a<đa<p�a<(�a<��a<��a<q�a<+�a<�a<��a<��a<b�a<,�a<��a<׎a<��a<��a<x�a<Z�a<E�a<1�a<	�a< �a<��a<��a<�a<�a<�a<�a<��a<�a<�a<�a<"�a<@�a<P�a<�  �  _�a<��a<��a<͎a<��a<(�a<g�a<t�a<��a<�a<1�a<_�a<��a<��a<�a<��a<��a<�a<V�a<��a<��a<I�a<��a<��a<Z�a<��a<#�a<��a<ѕa<Y�a<��a<(�a<}�a<��a<n�a<ʘa<Z�a<��a</�a<��a<�a<t�a<�a<~�a<Ϝa<V�a<��a<E�a<��a<�a<��a<�a<��a<ݠa<h�a<֡a<?�a<��a<�a<��a<�a<`�a<��a<"�a<��a<ϥa<J�a<��a<�a<Q�a<��a<�a<G�a<��a<Ҩa<D�a<y�a<ɩa<
�a<7�a<��a<��a<�a<%�a<x�a<��a<ȫa<�a<(�a<x�a<��a<��a<�a<��a<'�a<'�a<u�a<m�a<��a<��a<��a<ݭa<�a<�a<�a<"�a<"�a<�a<(�a<-�a<O�a<1�a<:�a<C�a<9�a<5�a<�a<>�a<�a<&�a<��a<�a<�a<ҭa<­a<��a<��a<w�a<X�a<=�a<'�a<�a<Ԭa<ʬa<��a<��a<M�a<'�a<�a<ǫa<«a<g�a<K�a<�a<�a<��a<m�a<R�a<��a<��a<}�a<L�a<�a<��a<��a<2�a<��a<��a<]�a<�a<��a<��a<�a<ӥa<q�a<*�a<��a<g�a<#�a<��a<T�a<ߢa<��a<1�a<��a<m�a<�a<��a<�a<Ɵa<Z�a<�a<��a<��a<��a<2�a<՜a<M�a<�a<��a<�a<��a<)�a<ߙa<d�a<�a<��a<�a<Ǘa<>�a<��a<��a<,�a<Ǖa<Q�a<�a<��a<W�a<ܓa<��a<J�a<��a<��a<A�a<�a<��a<d�a<4�a<�a<��a<O�a<D�a<�a<ɏa<��a<L�a<2�a<��a<�a<��a<��a<u�a<M�a<5�a<�a<*�a<��a<��a<��a<�a<�a<֍a< �a<ߍa<�a<��a<�a<*�a<:�a<V�a<�  �  y�a<��a<��a<֎a<�a<)�a<N�a<��a<��a<��a<(�a<q�a<��a<ڐa<�a<q�a<��a<�a<Q�a<��a<��a<N�a<��a<�a<i�a<Ɣa<'�a<�a<�a<N�a<��a<!�a<��a<��a<d�a<̘a<D�a<��a<,�a<��a<�a<��a<��a<e�a<�a<T�a<ϝa<7�a<��a<#�a<��a<�a<��a<��a<g�a<ɡa<6�a<��a<�a<��a<�a<T�a<��a< �a<{�a<�a<F�a<��a<��a<Z�a<��a<��a<I�a<��a<�a<1�a<v�a<��a<�a<Q�a<��a<ªa<�a<B�a<s�a<��a<ܫa<�a<?�a<X�a<��a<��a<ݬa<��a<-�a<;�a<]�a<i�a<��a<��a<˭a<حa<�a<��a<�a<�a<�a<5�a</�a<8�a<1�a<K�a<:�a<5�a<2�a<;�a<7�a<$�a<�a<�a<�a<��a<�a<ʭa<��a<��a<��a<�a<a�a<N�a<(�a< �a<�a<��a<��a<z�a<`�a<.�a<��a<ǫa<��a<u�a<U�a<�a<�a<��a<q�a<1�a<�a<Ωa<��a<O�a<�a<ʨa<��a<2�a<��a<��a<^�a<�a<��a<q�a<(�a<Хa<p�a<�a<ɤa<u�a<
�a<��a<R�a<��a<��a<.�a<ša<\�a<��a<��a<2�a<Ɵa<M�a<��a<��a<�a<��a<5�a<ɜa<[�a<�a<|�a<�a<��a<@�a<̙a<m�a<�a<��a<"�a<��a<]�a<�a<��a<#�a<a<k�a<�a<��a<L�a<��a<��a<G�a<��a<��a<X�a<��a<��a<m�a<-�a<��a<��a<c�a<+�a<�a<��a<��a<c�a<-�a<�a<Ԏa<��a<��a<p�a<c�a<<�a<)�a<�a<�a<��a<�a<�a<�a<�a<�a<ߍa<��a<�a<�a<#�a<2�a<S�a<�  �  ��a<��a<��a<Ǝa<�a<4�a<H�a<��a<��a<��a<�a<f�a<��a<�a<A�a<l�a<��a<�a<Q�a<��a<��a<e�a<��a<�a<W�a<��a<$�a<��a<��a<3�a<͖a<�a<��a<�a<Y�a<�a<.�a<��a<�a<��a<�a<{�a<��a<X�a<��a<B�a<ڝa<2�a<��a<2�a<��a<�a<r�a<��a<X�a<ءa<J�a<��a<$�a<x�a<�a<M�a<¤a<(�a<t�a<��a<.�a<��a<�a<W�a<��a<�a<_�a<��a<�a<�a<��a<��a<��a<H�a<~�a<ުa<�a<F�a<r�a<��a<�a<��a<K�a<P�a<��a<��a<Ӭa<��a<�a<F�a<T�a<��a<��a<��a<ía<ĭa<�a<�a<�a<�a<#�a<5�a<�a<H�a<'�a<R�a<,�a<D�a<?�a<+�a<'�a<�a<0�a<��a<��a<�a<�a<�a<��a<��a<��a<��a<Q�a<H�a<3�a<��a<��a<��a<��a<l�a<T�a<'�a< �a<�a<��a<}�a<C�a<�a<ުa<��a<��a<+�a<�a<��a<��a<L�a<�a<רa<e�a<R�a<�a<��a<R�a<�a<Цa<[�a<�a<��a<��a<�a<��a<u�a<��a<ȣa<A�a<�a<��a<0�a<ӡa<W�a<�a<��a<4�a<��a<\�a<��a<s�a<�a<��a<>�a<Üa<d�a<��a<u�a<)�a<��a<Q�a<Ùa<j�a<��a<�a<8�a<��a<W�a<ٖa<��a<!�a<��a<c�a<��a<��a<3�a<��a<��a<C�a<��a<��a<d�a<�a<ʑa<m�a<"�a<�a<��a<n�a<"�a<�a<��a<��a<[�a<�a<�a<̎a<Ǝa<��a<v�a<c�a<-�a<9�a<�a<�a<�a<��a<�a<ۍa<ލa<эa<�a<�a<��a<�a<'�a<I�a<>�a<�  �  o�a<��a<��a<Ԏa<��a<�a<X�a<��a<��a<�a<2�a<b�a<��a<�a<�a<x�a<��a<�a<c�a<��a<��a<P�a<��a<��a<[�a<Ôa<�a<��a<�a<F�a<��a<�a<��a<��a<b�a<֘a<K�a<��a<#�a<��a<
�a<x�a<��a<g�a<�a<R�a<ŝa<7�a<��a<�a<��a<�a<~�a<�a<\�a<ҡa<?�a<��a<�a<��a<�a<W�a<��a<#�a<�a<�a<>�a<��a<��a<O�a<��a<��a<L�a<��a<�a<:�a<~�a<��a<�a<G�a<��a<Ǫa<��a<2�a<q�a<��a<߫a<�a<.�a<c�a<��a<��a<۬a<�a<�a<7�a<^�a<t�a<��a<��a<��a<ۭa<�a<��a<�a<�a<�a<$�a<.�a<:�a<:�a<=�a<9�a<:�a</�a<0�a<.�a<,�a< �a<�a<�a<�a<֭a<֭a<��a<��a<��a<|�a<_�a<?�a<�a<
�a<�a<ìa<��a<��a<P�a<�a<	�a<ʫa<��a<n�a<C�a<"�a<�a<��a<t�a<A�a<��a<��a<��a<F�a<�a<èa<y�a<?�a<�a<��a<e�a<�a<Ħa<x�a<�a<ǥa<v�a<�a<��a<k�a<�a<��a<P�a<�a<��a</�a<��a<c�a< �a<��a<$�a<��a<V�a<�a<|�a<�a<��a<=�a<͜a<S�a<�a<�a<�a<��a<E�a<̙a<b�a<�a<��a<%�a<��a<U�a<��a<��a<$�a<ʕa<a�a<��a<��a<F�a<�a<��a<@�a<��a<��a<G�a<�a<��a<k�a<*�a<�a<��a<_�a<-�a<�a<Ïa<y�a<T�a<1�a<�a<ڎa<��a<��a<e�a<R�a<;�a<+�a<�a<�a<��a<�a<ލa<�a<�a<�a<�a<��a<�a<�a<�a<>�a<P�a<�  �  ^�a<��a<��a<ڎa<�a<!�a<l�a<v�a<ˏa<ݏa</�a<m�a<��a<��a<�a<��a<��a<�a<T�a<��a<�a<E�a<a<��a<w�a<��a<�a<��a<ܕa<i�a<��a<-�a<��a<�a<f�a<��a<G�a<��a<8�a<��a<�a<��a<�a<j�a<ʜa<h�a<ĝa<M�a<��a<"�a<��a<��a<��a<�a<m�a<ѡa<<�a<��a<�a<��a<ޣa<_�a<��a<&�a<��a<ݥa<V�a<��a<��a<L�a<��a<�a<5�a<��a<ܨa<5�a<p�a<��a<�a<G�a<��a<��a<�a<.�a<r�a<��a<ҫa<�a<+�a<y�a<��a<ìa<լa<��a<6�a<:�a<o�a<l�a<��a<��a<ŭa<�a<ԭa<�a<��a<)�a<!�a<+�a<=�a<�a<A�a<.�a<O�a<5�a</�a<D�a<$�a<-�a<��a<�a<��a<�a<�a<ɭa<֭a<��a<��a<a�a<e�a<L�a< �a<�a<׬a<լa<��a<��a<[�a<)�a<�a<ƫa<��a<o�a<Y�a<�a<֪a<��a<h�a<U�a<��a<ܩa<��a<7�a<�a<��a<��a<)�a< �a<��a<W�a<�a<��a<u�a<�a<ܥa<d�a<'�a<Ȥa<d�a<�a<��a<f�a<�a<��a<:�a<áa<m�a<�a<��a<(�a<˟a<U�a<�a<��a<�a<��a<)�a<Ԝa<a�a<��a<��a<�a<��a<+�a<˙a<_�a<��a<��a<�a<ϗa<H�a<�a<}�a<$�a<��a<a�a<�a<��a<d�a<�a<��a<5�a<�a<��a<D�a<�a<��a<~�a<%�a<ܐa<��a<b�a<=�a<�a<̏a<��a<]�a<5�a<�a<�a<��a<��a<t�a<Y�a<J�a<�a<�a<��a<
�a<�a<ލa<�a<ۍa<�a<ύa<��a<��a<�a<$�a<1�a<j�a<�  �  q�a<��a<��a<֎a<��a<'�a<S�a<�a<Ïa<��a<(�a<]�a<��a<�a<2�a<o�a<��a<�a<W�a<��a<�a<J�a<��a<�a<^�a<��a<(�a<��a<�a<O�a<��a<!�a<��a<�a<m�a<ݘa<E�a<��a<.�a<��a<�a<y�a<��a<t�a<�a<S�a<��a<>�a<��a<(�a<��a<�a<}�a<�a<^�a<ӡa<A�a<��a<�a<��a<�a<]�a<��a<�a<��a<ڥa<=�a<��a<�a<[�a<��a<�a<;�a<��a<ݨa<2�a<��a<ͩa<�a<A�a<��a<��a<�a<8�a<�a<��a<ݫa<�a<1�a<c�a<��a<��a<�a<��a<�a<9�a<W�a<|�a<��a<��a<��a<ѭa<�a< �a<�a<�a<"�a<�a<3�a<8�a<H�a<@�a<7�a<;�a<2�a<8�a<#�a<*�a<&�a<�a<��a<��a<�a<ͭa<��a<��a<��a<}�a<a�a<<�a<&�a<�a<߬a<ͬa<��a<z�a<K�a<)�a<�a<ܫa<��a<r�a<B�a<�a<�a<��a<n�a<>�a< �a<éa<��a<P�a<�a<ƨa<��a<0�a<��a<��a<Y�a<�a<˦a<s�a<�a<ҥa<g�a<"�a<��a<r�a<�a<��a<R�a<�a<��a<'�a<ɡa<h�a<�a<��a<#�a<��a<W�a<�a<z�a<�a<��a<<�a<Ҝa<b�a<�a<��a<�a<��a<B�a<ٙa<o�a<�a<��a<�a<Ɨa<I�a<�a<��a<0�a<��a<[�a<�a<��a<P�a<�a<��a<I�a<��a<��a<J�a<�a<��a<w�a<2�a<�a<��a<a�a<&�a<��a<��a<��a<N�a<'�a<�a<��a<��a<��a<u�a<M�a<@�a<)�a<"�a<	�a<�a<�a<�a<�a<ڍa<�a<��a<��a<��a<�a<"�a<5�a<Q�a<�  �  v�a<u�a<��a<ێa<��a<:�a<I�a<��a<��a<��a<$�a<a�a<��a<Րa</�a<e�a<֑a<��a<^�a<��a<�a<N�a<��a<�a<Y�a<Ɣa<�a<r�a<�a<D�a<a<�a<��a< �a<N�a<ʘa<=�a<��a<$�a<��a<�a<~�a<��a<S�a<�a<F�a<ԝa<G�a<��a<"�a<��a<�a<l�a<�a<i�a<ԡa<A�a<��a<0�a<m�a<��a<I�a<��a<�a<��a<�a</�a<��a<�a<S�a<��a<�a<F�a<��a<�a<.�a<m�a<��a<
�a<I�a<y�a<ͪa< �a<@�a<d�a<��a<�a<��a<J�a<]�a<��a<��a<�a<	�a<�a<X�a<Q�a<|�a<��a<��a<ía<ʭa<��a<�a<�a<�a<2�a<+�a</�a<3�a< �a<H�a<2�a<G�a<,�a<2�a<5�a<�a<�a<��a<�a<�a<խa<ݭa<��a<��a<z�a<y�a<f�a<C�a<9�a<��a<�a<��a<��a<v�a<O�a<B�a<�a<٫a<��a<��a<8�a<�a<�a<��a<q�a<7�a<�a<��a<��a<A�a<��a<ɨa<w�a<F�a<�a<��a<g�a<��a<��a<k�a<#�a<ȥa<p�a<)�a<¤a<r�a<��a<��a<D�a<��a<��a<%�a<áa<P�a<�a<��a<<�a<ȟa<X�a<�a<~�a<(�a<��a<H�a<��a<U�a<�a<��a<"�a<��a<E�a<��a<f�a<��a<��a<�a<��a<Y�a<�a<z�a<�a<Ǖa<c�a<��a<��a<I�a<��a<��a<5�a<��a<��a<c�a<��a<��a<\�a<0�a<�a<��a<��a< �a<��a<��a<��a<[�a< �a<�a<a<��a<��a<��a<X�a<<�a<%�a<��a<�a<�a<��a<܍a<�a<�a<Ӎa<�a<ލa<�a<�a<�a<E�a<H�a<�  �  q�a<��a<��a<֎a<��a<'�a<S�a<�a<Ïa<��a<(�a<]�a<��a<�a<2�a<o�a<��a<�a<W�a<��a<�a<J�a<��a<�a<^�a<��a<(�a<��a<�a<O�a<��a<!�a<��a<�a<m�a<ݘa<E�a<��a<.�a<��a<�a<y�a<��a<t�a<�a<S�a<��a<>�a<��a<(�a<��a<�a<}�a<�a<^�a<ӡa<A�a<��a<�a<��a<�a<]�a<��a<�a<��a<ڥa<=�a<��a<�a<[�a<��a<�a<;�a<��a<ݨa<2�a<��a<ͩa<�a<A�a<��a<��a<�a<8�a<�a<��a<ݫa<�a<1�a<c�a<��a<��a<�a<��a<�a<9�a<W�a<|�a<��a<��a<��a<ѭa<�a< �a<�a<�a<"�a<�a<3�a<8�a<H�a<@�a<7�a<;�a<2�a<8�a<#�a<*�a<&�a<�a<��a<��a<�a<ͭa<��a<��a<��a<}�a<a�a<<�a<&�a<�a<߬a<ͬa<��a<z�a<K�a<)�a<�a<ܫa<��a<r�a<B�a<�a<�a<��a<n�a<>�a< �a<éa<��a<P�a<�a<ƨa<��a<0�a<��a<��a<Y�a<�a<˦a<s�a<�a<ҥa<g�a<"�a<��a<r�a<�a<��a<R�a<�a<��a<'�a<ɡa<h�a<�a<��a<#�a<��a<W�a<�a<z�a<�a<��a<<�a<Ҝa<b�a<�a<��a<�a<��a<B�a<ٙa<o�a<�a<��a<�a<Ɨa<I�a<�a<��a<0�a<��a<[�a<�a<��a<P�a<�a<��a<I�a<��a<��a<J�a<�a<��a<w�a<2�a<�a<��a<a�a<&�a<��a<��a<��a<N�a<'�a<�a<��a<��a<��a<u�a<M�a<@�a<)�a<"�a<	�a<�a<�a<�a<�a<ڍa<�a<��a<��a<��a<�a<"�a<5�a<Q�a<�  �  ^�a<��a<��a<ڎa<�a<!�a<l�a<v�a<ˏa<ݏa</�a<m�a<��a<��a<�a<��a<��a<�a<T�a<��a<�a<E�a<a<��a<w�a<��a<�a<��a<ܕa<i�a<��a<-�a<��a<�a<f�a<��a<G�a<��a<8�a<��a<�a<��a<�a<j�a<ʜa<h�a<ĝa<M�a<��a<"�a<��a<��a<��a<�a<m�a<ѡa<<�a<��a<�a<��a<ޣa<_�a<��a<&�a<��a<ݥa<V�a<��a<��a<L�a<��a<�a<5�a<��a<ܨa<5�a<p�a<��a<�a<G�a<��a<��a<�a<.�a<r�a<��a<ҫa<�a<+�a<y�a<��a<ìa<լa<��a<6�a<:�a<o�a<l�a<��a<��a<ŭa<�a<ԭa<�a<��a<)�a<!�a<+�a<=�a<�a<A�a<.�a<O�a<5�a</�a<D�a<$�a<-�a<��a<�a<��a<�a<�a<ɭa<֭a<��a<��a<a�a<e�a<L�a< �a<�a<׬a<լa<��a<��a<[�a<)�a<�a<ƫa<��a<o�a<Y�a<�a<֪a<��a<h�a<U�a<��a<ܩa<��a<7�a<�a<��a<��a<)�a< �a<��a<W�a<�a<��a<u�a<�a<ܥa<d�a<'�a<Ȥa<d�a<�a<��a<f�a<�a<��a<:�a<áa<m�a<�a<��a<(�a<˟a<U�a<�a<��a<�a<��a<)�a<Ԝa<a�a<��a<��a<�a<��a<+�a<˙a<_�a<��a<��a<�a<ϗa<H�a<�a<}�a<$�a<��a<a�a<�a<��a<d�a<�a<��a<5�a<�a<��a<D�a<�a<��a<~�a<%�a<ܐa<��a<b�a<=�a<�a<̏a<��a<]�a<5�a<�a<�a<��a<��a<t�a<Y�a<J�a<�a<�a<��a<
�a<�a<ލa<�a<ۍa<�a<ύa<��a<��a<�a<$�a<1�a<j�a<�  �  o�a<��a<��a<Ԏa<��a<�a<X�a<��a<��a<�a<2�a<b�a<��a<�a<�a<x�a<��a<�a<c�a<��a<��a<P�a<��a<��a<[�a<Ôa<�a<��a<�a<F�a<��a<�a<��a<��a<b�a<֘a<K�a<��a<#�a<��a<
�a<x�a<��a<g�a<�a<R�a<ŝa<7�a<��a<�a<��a<�a<~�a<�a<\�a<ҡa<?�a<��a<�a<��a<�a<W�a<��a<#�a<�a<�a<>�a<��a<��a<O�a<��a<��a<L�a<��a<�a<:�a<~�a<��a<�a<G�a<��a<Ǫa<��a<2�a<q�a<��a<߫a<�a<.�a<c�a<��a<��a<۬a<�a<�a<7�a<^�a<t�a<��a<��a<��a<ۭa<�a<��a<�a<�a<�a<$�a<.�a<:�a<:�a<=�a<9�a<:�a</�a<0�a<.�a<,�a< �a<�a<�a<�a<֭a<֭a<��a<��a<��a<|�a<_�a<?�a<�a<
�a<�a<ìa<��a<��a<P�a<�a<	�a<ʫa<��a<n�a<C�a<"�a<�a<��a<t�a<A�a<��a<��a<��a<F�a<�a<èa<y�a<?�a<�a<��a<e�a<�a<Ħa<x�a<�a<ǥa<v�a<�a<��a<k�a<�a<��a<P�a<�a<��a</�a<��a<c�a< �a<��a<$�a<��a<V�a<�a<|�a<�a<��a<=�a<͜a<S�a<�a<�a<�a<��a<E�a<̙a<b�a<�a<��a<%�a<��a<U�a<��a<��a<$�a<ʕa<a�a<��a<��a<F�a<�a<��a<@�a<��a<��a<G�a<�a<��a<k�a<*�a<�a<��a<_�a<-�a<�a<Ïa<y�a<T�a<1�a<�a<ڎa<��a<��a<e�a<R�a<;�a<+�a<�a<�a<��a<�a<ލa<�a<�a<�a<�a<��a<�a<�a<�a<>�a<P�a<�  �  ��a<��a<��a<Ǝa<�a<4�a<H�a<��a<��a<��a<�a<f�a<��a<�a<A�a<l�a<��a<�a<Q�a<��a<��a<e�a<��a<�a<W�a<��a<$�a<��a<��a<3�a<͖a<�a<��a<�a<Y�a<�a<.�a<��a<�a<��a<�a<{�a<��a<X�a<��a<B�a<ڝa<2�a<��a<2�a<��a<�a<r�a<��a<X�a<ءa<J�a<��a<$�a<x�a<�a<M�a<¤a<(�a<t�a<��a<.�a<��a<�a<W�a<��a<�a<_�a<��a<�a<�a<��a<��a<��a<H�a<~�a<ުa<�a<F�a<r�a<��a<�a<��a<K�a<P�a<��a<��a<Ӭa<��a<�a<F�a<T�a<��a<��a<��a<ía<ĭa<�a<�a<�a<�a<#�a<5�a<�a<H�a<'�a<R�a<,�a<D�a<?�a<+�a<'�a<�a<0�a<��a<��a<�a<�a<�a<��a<��a<��a<��a<Q�a<H�a<3�a<��a<��a<��a<��a<l�a<T�a<'�a< �a<�a<��a<}�a<C�a<�a<ުa<��a<��a<+�a<�a<��a<��a<L�a<�a<רa<e�a<R�a<�a<��a<R�a<�a<Цa<[�a<�a<��a<��a<�a<��a<u�a<��a<ȣa<A�a<�a<��a<0�a<ӡa<W�a<�a<��a<4�a<��a<\�a<��a<s�a<�a<��a<>�a<Üa<d�a<��a<u�a<)�a<��a<Q�a<Ùa<j�a<��a<�a<8�a<��a<W�a<ٖa<��a<!�a<��a<c�a<��a<��a<3�a<��a<��a<C�a<��a<��a<d�a<�a<ʑa<m�a<"�a<�a<��a<n�a<"�a<�a<��a<��a<[�a<�a<�a<̎a<Ǝa<��a<v�a<c�a<-�a<9�a<�a<�a<�a<��a<�a<ۍa<ލa<эa<�a<�a<��a<�a<'�a<I�a<>�a<�  �  y�a<��a<��a<֎a<�a<)�a<N�a<��a<��a<��a<(�a<q�a<��a<ڐa<�a<q�a<��a<�a<Q�a<��a<��a<N�a<��a<�a<i�a<Ɣa<'�a<�a<�a<N�a<��a<!�a<��a<��a<d�a<̘a<D�a<��a<,�a<��a<�a<��a<��a<e�a<�a<T�a<ϝa<7�a<��a<#�a<��a<�a<��a<��a<g�a<ɡa<6�a<��a<�a<��a<�a<T�a<��a< �a<{�a<�a<F�a<��a<��a<Z�a<��a<��a<I�a<��a<�a<1�a<v�a<��a<�a<Q�a<��a<ªa<�a<B�a<s�a<��a<ܫa<�a<?�a<X�a<��a<��a<ݬa<��a<-�a<;�a<]�a<i�a<��a<��a<˭a<حa<�a<��a<�a<�a<�a<5�a</�a<8�a<1�a<K�a<:�a<5�a<2�a<;�a<7�a<$�a<�a<�a<�a<��a<�a<ʭa<��a<��a<��a<�a<a�a<N�a<(�a< �a<�a<��a<��a<z�a<`�a<.�a<��a<ǫa<��a<u�a<U�a<�a<�a<��a<q�a<1�a<�a<Ωa<��a<O�a<�a<ʨa<��a<2�a<��a<��a<^�a<�a<��a<q�a<(�a<Хa<p�a<�a<ɤa<u�a<
�a<��a<R�a<��a<��a<.�a<ša<\�a<��a<��a<2�a<Ɵa<M�a<��a<��a<�a<��a<5�a<ɜa<[�a<�a<|�a<�a<��a<@�a<̙a<m�a<�a<��a<"�a<��a<]�a<�a<��a<#�a<a<k�a<�a<��a<L�a<��a<��a<G�a<��a<��a<X�a<��a<��a<m�a<-�a<��a<��a<c�a<+�a<�a<��a<��a<c�a<-�a<�a<Ԏa<��a<��a<p�a<c�a<<�a<)�a<�a<�a<��a<�a<�a<�a<�a<�a<ߍa<��a<�a<�a<#�a<2�a<S�a<�  �  _�a<��a<��a<͎a<��a<(�a<g�a<t�a<��a<�a<1�a<_�a<��a<��a<�a<��a<��a<�a<V�a<��a<��a<I�a<��a<��a<Z�a<��a<#�a<��a<ѕa<Y�a<��a<(�a<}�a<��a<n�a<ʘa<Z�a<��a</�a<��a<�a<t�a<�a<~�a<Ϝa<V�a<��a<E�a<��a<�a<��a<�a<��a<ݠa<h�a<֡a<?�a<��a<�a<��a<�a<`�a<��a<"�a<��a<ϥa<J�a<��a<�a<Q�a<��a<�a<G�a<��a<Ҩa<D�a<y�a<ɩa<
�a<7�a<��a<��a<�a<%�a<x�a<��a<ȫa<�a<(�a<x�a<��a<��a<�a<��a<'�a<'�a<u�a<m�a<��a<��a<��a<ݭa<�a<�a<�a<"�a<"�a<�a<(�a<-�a<O�a<1�a<:�a<C�a<9�a<5�a<�a<>�a<�a<&�a<��a<�a<�a<ҭa<­a<��a<��a<w�a<X�a<=�a<'�a<�a<Ԭa<ʬa<��a<��a<M�a<'�a<�a<ǫa<«a<g�a<K�a<�a<�a<��a<m�a<R�a<��a<��a<}�a<L�a<�a<��a<��a<2�a<��a<��a<]�a<�a<��a<��a<�a<ӥa<q�a<*�a<��a<g�a<#�a<��a<T�a<ߢa<��a<1�a<��a<m�a<�a<��a<�a<Ɵa<Z�a<�a<��a<��a<��a<2�a<՜a<M�a<�a<��a<�a<��a<)�a<ߙa<d�a<�a<��a<�a<Ǘa<>�a<��a<��a<,�a<Ǖa<Q�a<�a<��a<W�a<ܓa<��a<J�a<��a<��a<A�a<�a<��a<d�a<4�a<�a<��a<O�a<D�a<�a<ɏa<��a<L�a<2�a<��a<�a<��a<��a<u�a<M�a<5�a<�a<*�a<��a<��a<��a<�a<�a<֍a< �a<ߍa<�a<��a<�a<*�a<:�a<V�a<�  �  k�a<��a<��a<ݎa<��a<-�a<K�a<��a<��a<�a<*�a<l�a<��a<�a<�a<o�a<Ƒa<�a<P�a<��a<��a<b�a<��a<�a<a�a<Δa<�a<��a<�a<J�a<��a<#�a<��a<��a<X�a<Ęa<D�a<��a<4�a<��a<�a<}�a<��a<_�a<�a<[�a<͝a<>�a<��a</�a<��a<
�a<��a<��a<^�a<Ρa<:�a<��a<"�a<��a<�a<X�a<Ǥa<)�a<��a<�a<G�a<��a<�a<Q�a<��a<��a<H�a<��a<�a<6�a<p�a<��a<�a<S�a<��a<Ǫa<��a<8�a<s�a<��a<�a<	�a<8�a<]�a<��a<��a<جa<��a<&�a<I�a<\�a<o�a<��a<��a<ʭa<׭a<߭a<��a<�a<�a<%�a<-�a<7�a<?�a</�a<8�a<;�a<B�a<2�a<A�a<+�a<#�a<�a<�a<�a<�a<�a<حa<��a<��a<��a<~�a<h�a<F�a<,�a<��a<�a<Ĭa<��a<{�a<Z�a</�a<�a<ȫa<��a<��a<P�a<�a<ݪa<��a<��a<5�a<�a<Ʃa<��a<G�a<
�a<¨a<|�a<?�a<��a<��a<d�a<�a<��a<q�a<�a<٥a<p�a< �a<��a<k�a<�a<��a<Y�a<��a<��a<1�a<Сa<b�a<��a<��a<2�a<��a<R�a<�a<{�a<�a<��a<6�a<Μa<i�a<��a<��a<�a<��a<>�a<Ǚa<d�a<��a<��a<!�a<ȗa<V�a<�a<}�a<�a<ʕa<m�a<
�a<��a<F�a<�a<��a<?�a<��a<��a<Q�a<��a<đa<p�a<(�a<��a<��a<q�a<+�a<�a<��a<��a<b�a<,�a<��a<׎a<��a<��a<x�a<Z�a<E�a<1�a<	�a< �a<��a<��a<�a<�a<�a<�a<��a<�a<�a<�a<"�a<@�a<P�a<�  �  ��a<}�a<��a<Վa<��a<1�a<J�a<��a<��a<�a<(�a<b�a<��a<Րa<>�a<Z�a<��a<��a<^�a<��a<�a<e�a<��a<�a<Q�a<ϔa< �a<}�a<��a<D�a<��a<�a<��a<�a<f�a<�a<:�a<��a<�a<��a<�a<��a<�a<W�a<�a<B�a<՝a<9�a<��a<.�a<��a<$�a<t�a<�a<R�a<ѡa<F�a<��a<�a<v�a<�a<E�a<��a<%�a<y�a<��a<.�a<��a<�a<Z�a<��a<�a<O�a<��a<�a<)�a<��a<ȩa<��a<Q�a<z�a<Ҫa<��a<I�a<q�a<��a<�a<��a<M�a<O�a<��a<��a<٬a<	�a<�a<>�a<G�a<��a<��a<��a<��a<ϭa<��a<ݭa<�a<�a<$�a<#�a<*�a<K�a<'�a<P�a<7�a<;�a<0�a<0�a<0�a<"�a<2�a<�a<�a<��a<׭a<حa<��a<��a<��a<��a<`�a<7�a<0�a<��a<��a<��a<��a<y�a<P�a<%�a<�a<�a<��a<t�a<=�a<�a<�a<��a<��a<)�a<�a<��a<��a<I�a<�a<֨a<v�a<C�a<�a<��a<V�a<�a<Ӧa<h�a<&�a<��a<u�a<�a<Ĥa<z�a<��a<ƣa<@�a<��a<��a<.�a<Сa<K�a<�a<��a<*�a<��a<U�a<�a<k�a<�a<��a<N�a<��a<_�a<��a<y�a<)�a<��a<P�a<��a<m�a<��a<��a<'�a<��a<^�a<�a<��a<+�a<��a<k�a<��a<��a<A�a< �a<��a<<�a<�a<��a<g�a<�a<őa<g�a<(�a<�a<��a<f�a<�a<�a<��a<�a<V�a<%�a<�a<��a<ǎa<��a<w�a<Q�a<7�a<=�a<�a<�a<�a<�a<ߍa<�a<�a<�a<�a<��a<�a<�a<�a<@�a<K�a<�  �  l�a<��a<��a<ώa<��a<)�a<Y�a<��a<��a<��a<�a<a�a<��a<�a<0�a<y�a<��a<�a<Q�a<��a<��a<T�a<��a<
�a<_�a<��a<�a<��a<�a<Q�a<��a<$�a<��a<�a<j�a<јa<D�a<��a<$�a<��a<�a<|�a<��a<j�a<ٜa<N�a<ѝa<9�a<��a<�a<��a<�a<y�a<�a<h�a<ϡa<@�a<��a<�a<�a<�a<P�a<��a<�a<}�a<�a<=�a<��a<��a<S�a<��a<��a<Q�a<��a<�a<2�a<{�a<ũa<��a<C�a<��a<˪a<�a<2�a<r�a<��a<ӫa<�a<=�a<_�a<��a<��a<֬a<��a<�a<<�a<e�a<|�a<��a<��a<��a<ǭa<�a<�a<�a<�a<�a<+�a<*�a<*�a<>�a<;�a<:�a<=�a<E�a<0�a<!�a<,�a<�a<�a<��a<�a<�a<׭a<��a<��a<��a<o�a<[�a<D�a<(�a<�a<�a<��a<��a<k�a<O�a<1�a<�a<ګa<��a<w�a<E�a<�a<�a<��a<x�a<;�a<�a<ĩa<��a<<�a<�a<��a<��a<>�a<��a<��a<O�a<�a<��a<r�a<�a<ɥa<|�a<�a<��a<k�a<�a<��a<L�a<��a<��a<*�a<��a<\�a<��a<��a<(�a<ǟa<S�a<�a<��a<�a<��a<8�a<Ŝa<Q�a<�a<~�a<�a<��a<9�a<͙a<f�a<�a<��a<*�a<��a<N�a<�a<��a<(�a<��a<]�a<�a<��a<N�a<�a<��a<<�a<�a<��a<V�a< �a<��a<h�a<&�a<�a<��a<d�a<3�a<��a<��a<��a<T�a<�a<�a<юa<��a<��a<r�a<Y�a<7�a<�a<�a<�a<��a<��a<�a<��a<؍a<�a<ߍa<��a<�a<�a</�a<?�a<Q�a<�  �  _�a<��a<��a<��a<��a<�a<\�a<w�a<ҏa<�a<,�a<p�a<��a<�a<�a<{�a<��a<�a<K�a<��a<
�a<F�a<��a<�a<s�a<��a<&�a<��a<ܕa<]�a<��a<+�a<��a<��a<p�a<Șa<U�a<��a<?�a<��a<�a<��a<�a<~�a<Ӝa<i�a<��a<0�a<��a<�a<��a<�a<��a<�a<`�a<͡a<7�a<��a<�a<��a<գa<k�a<��a<�a<{�a<եa<V�a<��a<�a<S�a<��a< �a<=�a<��a<�a<E�a<u�a<ũa<�a<I�a<��a<��a<�a<4�a<��a<��a<իa<�a<"�a<e�a<��a<��a<ެa<�a<1�a<1�a<c�a<b�a<��a<��a<ŭa<�a<٭a<�a<��a<�a<�a<'�a<C�a<)�a<R�a<.�a<M�a<-�a<9�a<B�a<$�a<<�a<�a<(�a<��a<��a<�a<��a<ϭa<��a<��a<r�a<k�a<F�a<�a<�a<׬a<ݬa<��a<}�a<^�a<!�a<�a<��a<��a<m�a<Y�a<
�a<ߪa<��a<j�a<B�a<�a<ةa<��a<O�a<�a<��a<��a<'�a<��a<��a<c�a<�a<��a<��a<�a<�a<h�a<�a<Ѥa<c�a<#�a<��a<g�a<�a<��a<+�a<��a<y�a<�a<��a<%�a<��a<Q�a<�a<~�a<�a<��a<�a<��a<W�a<�a<{�a<�a<��a<3�a<�a<f�a<��a<��a<�a<՗a<Q�a< �a<��a<(�a<Εa<c�a<�a<��a<W�a<�a<��a<Q�a<�a<��a<;�a<�a<��a<v�a<.�a<אa<��a<Y�a<1�a<ۏa<��a<��a<]�a<6�a<�a<�a<��a<��a<_�a<U�a<P�a<�a<,�a<��a<	�a<��a<�a<�a<ۍa<��a<ݍa<�a<��a<�a<)�a<(�a<c�a<�  �  f�a<��a<��a<Ύa<��a<,�a<g�a<��a<��a<�a<(�a<h�a<��a<�a<4�a<w�a<��a<�a<N�a<��a<��a<W�a<��a<	�a<d�a<��a<$�a<�a<�a<U�a<��a<�a<��a<��a<c�a<՘a<>�a<��a< �a<��a<�a<��a<�a<h�a<לa<N�a<͝a<C�a<��a<#�a<��a<��a<��a<�a<]�a<ܡa<I�a<��a<�a<��a<ޣa<^�a<��a<-�a<��a<�a<<�a<��a<��a<J�a<��a<�a<N�a<��a<�a</�a<|�a<éa<�a<B�a<��a<ͪa<�a<;�a<n�a<��a<Ϋa<
�a<<�a<m�a<��a<��a<ܬa<�a<&�a<2�a<`�a<��a<��a<��a<��a<֭a<ޭa<��a<�a<%�a<&�a<'�a<,�a<4�a<;�a<4�a<E�a<C�a<:�a<.�a<'�a<%�a<$�a<�a< �a<�a<�a<׭a<ȭa<��a<��a<y�a<Y�a<C�a<+�a<�a<�a<ìa<��a<y�a<V�a<&�a<�a<ޫa<��a<m�a<M�a<�a<�a<��a<{�a<J�a<�a<ʩa<~�a<L�a<�a<Ĩa<��a<A�a<�a<��a<\�a<�a<æa<k�a<�a<ťa<t�a<&�a<ͤa<c�a<�a<��a<L�a<��a<��a<:�a<ġa<h�a<�a<��a<!�a<��a<`�a<�a<|�a<�a<��a<(�a<Ӝa<X�a<��a<��a<�a<��a<3�a<Ιa<]�a<��a<��a<&�a<��a<O�a<�a<��a<&�a<��a<\�a< �a<��a<Q�a<�a<��a<F�a<�a<��a<U�a<�a<��a<i�a<,�a<ِa<��a<Z�a<.�a<��a<ďa<��a<V�a<,�a<��a<׎a<��a<��a<y�a<U�a<9�a<%�a<�a<��a<�a<��a<�a<ލa<ލa<�a<��a<��a<��a<�a<%�a<?�a<\�a<�  �  Ԏa<�a<+�a<I�a<v�a<��a<��a<�a<1�a<q�a<��a<ʐa<�a<P�a<��a<ܑa<4�a<m�a<ڒa<"�a<p�a<ԓa<�a<b�a<Ӕa</�a<��a<�a<D�a<��a<'�a<��a<��a<d�a<Řa<Q�a<��a<)�a<w�a<��a<o�a<ӛa<M�a<̜a<J�a<��a<+�a<��a<�a<��a<��a<��a<Ѡa<I�a<��a<�a<��a<�a<l�a<ѣa<_�a<��a<$�a<}�a<ɥa<6�a<��a<��a<R�a<��a<�a<I�a<��a<بa<L�a<��a<ީa<�a<]�a<��a<̪a<�a<G�a<�a<��a<�a<1�a<]�a<}�a<��a<�a<�a<9�a<j�a<h�a<��a<��a<��a<ݭa<�a<�a<(�a<P�a<V�a<}�a<\�a<[�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<k�a<��a<U�a<g�a<M�a<2�a<+�a<�a<�a<�a<٭a<��a<��a<d�a<O�a<[�a<!�a<�a<جa<��a<��a<Q�a<�a<��a<ثa<��a<��a<D�a<	�a<�a<��a<I�a<"�a<�a<��a<\�a<�a<̨a<��a<@�a<�a<��a<_�a</�a<��a<��a<�a<˥a<t�a<�a<��a<g�a<�a<��a<L�a<٢a<��a<6�a<��a<m�a<�a<��a<�a<��a<:�a<۞a<k�a<��a<��a<5�a<Мa<Y�a<՛a<u�a<�a<��a<9�a<��a<N�a<�a<��a<�a<̗a<P�a<�a<��a<0�a<ܕa<_�a<�a<��a<O�a<��a<��a<c�a<�a<��a<e�a<5�a<�a<��a<n�a<
�a<ؐa<��a<P�a<#�a<��a<��a<��a<��a<R�a<F�a<��a<ˎa<Վa<��a<��a<��a<l�a<d�a<b�a<U�a<U�a<f�a<J�a<��a<X�a<��a<��a<��a<��a<��a<�  �  ��a<�a<�a<C�a<n�a<��a<Џa<ߏa<$�a<M�a<��a<Ԑa<�a<^�a<��a<�a<'�a<s�a<��a<�a<a�a<��a<*�a<s�a<Ӕa<%�a<��a<��a<f�a<ǖa< �a<��a<�a<[�a<ǘa<?�a<��a<�a<��a<�a<t�a<��a<d�a<ќa<0�a<��a<"�a<��a<
�a<i�a<�a<Z�a<۠a<L�a<áa</�a<��a<�a<q�a<ޣa<5�a<��a<��a<i�a<�a<4�a<��a<�a<O�a<��a<�a<U�a<��a<��a<6�a<��a<ϩa<�a<V�a<��a<�a<�a<b�a<��a<ͫa<�a<#�a<b�a<��a<Ȭa<Ǭa<��a<�a<A�a<p�a<��a<��a<Эa<�a<��a<�a<&�a<'�a<D�a<E�a<n�a<��a<z�a<��a<x�a<��a<��a<��a<��a<��a<��a<�a<s�a<u�a<_�a<V�a<H�a<D�a<#�a<'�a<�a<��a<��a<��a<��a<��a<g�a<$�a<�a<�a<ʬa<��a<{�a<_�a<0�a<�a<˫a<��a<_�a<)�a<��a<��a<��a<[�a<"�a<ةa<��a<h�a</�a<�a<��a<S�a<��a<��a<a�a<�a<Ŧa<p�a<)�a<ԥa<x�a<-�a<Ϥa<l�a<��a<��a<C�a<��a<�a<�a<��a<F�a<�a<��a<#�a<��a<K�a<�a<o�a<�a<��a<�a<��a<D�a<�a<t�a<�a<��a<5�a<әa<q�a<��a<��a<+�a<��a<S�a<�a<��a<)�a<��a<v�a<�a<Ĕa<r�a<�a<��a<U�a<�a<��a<��a<�a<Бa<��a<E�a<�a<Ԑa<��a<f�a<4�a<��a<ˏa<��a<\�a<@�a<�a<�a<�a<Ŏa<��a<��a<��a<��a<��a<[�a<b�a<Z�a<S�a<R�a<c�a<b�a<s�a<��a<��a<��a<؎a<�  �  юa<�a<�a<[�a<e�a<��a<͏a<��a<K�a<]�a<��a<ېa<��a<T�a<��a<ޑa<�a<��a<Ȓa<!�a<��a<��a<)�a<a�a<Дa<6�a<��a<�a<A�a<��a<	�a<��a<�a<o�a<͘a<'�a<��a<�a<��a<��a<[�a<қa<H�a<֜a<6�a<ŝa<�a<��a<�a<��a<�a<c�a<�a<9�a<��a<$�a<��a<��a<\�a<�a<=�a<Ĥa<�a<q�a<�a<&�a<��a<�a<P�a<��a<�a<=�a<��a<��a<,�a<��a<éa<�a<o�a<��a<�a<�a<K�a<z�a<��a<��a<,�a<b�a<u�a<Ǭa<ˬa<�a<=�a<O�a<��a<{�a<��a<ía<�a<�a<�a<7�a<4�a<k�a<J�a<k�a<}�a<n�a<��a<��a<��a<��a<��a<z�a<��a<��a<��a<��a<U�a<s�a<_�a<H�a<B�a<�a<�a<�a<��a<ƭa<ʭa<��a<�a<d�a<&�a<:�a<�a<ܬa<��a<h�a<U�a<$�a<��a<��a<��a<o�a<B�a<�a<��a<��a<H�a<�a<�a<��a<b�a<
�a<Ψa<z�a<V�a<��a<ħa<g�a<�a<ۦa<g�a<,�a<åa<`�a<�a<��a<q�a<��a<��a<7�a<��a<��a<"�a<סa<O�a<��a<r�a<�a<��a<>�a<Ӟa<Z�a<�a<��a<C�a<ɜa<L�a<�a<e�a<�a<��a<7�a<��a<J�a<�a<z�a<0�a<��a<j�a<�a<��a<B�a<��a<~�a<��a<��a<J�a< �a<��a<^�a<�a<��a<��a<�a<��a<��a<S�a<!�a<��a<��a<Y�a<*�a<�a<Ǐa<��a<i�a<g�a<�a<�a<�a<��a<Îa<��a<��a<e�a<f�a<J�a<^�a<[�a<X�a<l�a<C�a<v�a<{�a<��a<��a<��a<��a<�  �  ގa<�a< �a<G�a<s�a<��a<��a<�a<�a<Y�a<��a<ΐa<&�a<U�a<��a<�a<9�a<m�a<˒a<	�a<P�a<͓a<�a<w�a<Δa<.�a<��a<��a<R�a<ʖa<0�a<��a<��a<]�a<��a<8�a<��a<�a<�a<��a<��a<�a<W�a<ɜa<>�a<��a</�a<��a<�a<��a<��a<h�a<Ӡa<N�a<ȡa<(�a<��a<�a<x�a<ԣa<E�a<��a<�a<y�a<֥a<>�a<��a<�a<L�a<��a<��a<k�a<��a<�a<7�a<��a<Ωa<�a<W�a<��a<Ԫa<#�a<i�a<��a<ɫa<��a<-�a<Z�a<��a<��a<�a<��a<�a<U�a<g�a<��a<��a<ȭa<�a<�a<�a<"�a<8�a<1�a<h�a<]�a<{�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<t�a<p�a<\�a<X�a<M�a<3�a<@�a<"�a<��a<�a<έa<��a<��a<��a<R�a<K�a<��a<�a<Ϭa<��a<��a<V�a<'�a<��a<ݫa<��a<r�a<+�a<�a<٪a<��a<^�a<�a<�a<��a<f�a<�a<�a<��a<A�a<�a<��a<Z�a<�a<æa<p�a<�a<Υa<��a<#�a<��a<d�a<�a<��a<Q�a<�a<��a<&�a<��a<S�a<�a<��a<(�a<��a<D�a<�a<v�a<��a<��a<�a<��a<U�a<�a<~�a<�a<��a<2�a<˙a<a�a<�a<��a<�a<��a<R�a<�a<��a<*�a<Еa<g�a<�a<˔a<]�a<�a<��a<_�a<
�a<��a<n�a</�a<ʑa<��a<Y�a<	�a<�a<��a<]�a<,�a<�a<ďa<��a<m�a<-�a<1�a<��a<�a<юa<��a<��a<��a<t�a<v�a<z�a<V�a<T�a<U�a<S�a<^�a<_�a<t�a<��a<��a<Ŏa<ӎa<�  �  �a<��a<)�a<?�a<j�a<��a<��a<�a<�a<��a<��a<ːa<�a<B�a<��a<Αa<<�a<_�a<ǒa<*�a<`�a<ۓa<��a<��a<��a</�a<��a<�a<Z�a<��a<�a<|�a<�a<Y�a<͘a<P�a<��a<-�a<��a<��a<f�a<՛a<b�a<��a<S�a<��a<1�a<��a<�a<��a<�a<��a<��a<V�a<��a<+�a<��a<��a<��a<£a<Z�a<��a<�a<~�a<ɥa<A�a<��a<�a<E�a<��a<�a<A�a<��a<�a<R�a<v�a<�a<�a<M�a<��a<Ѫa<�a<A�a<��a<ǫa<��a<5�a<G�a<��a<��a<��a<�a<8�a<Y�a<Z�a<��a<��a<ܭa<حa<�a<�a<�a<^�a<<�a<x�a<X�a<z�a<~�a<x�a<��a<��a<��a<�a<��a<��a<��a<��a<n�a<��a<_�a<_�a<Z�a<*�a<"�a<��a<�a<�a<׭a<��a<��a<��a<H�a<X�a<�a<�a<Ȭa<��a<��a<C�a<<�a<�a<�a<��a<n�a<L�a<��a<�a<y�a<j�a<�a<�a<��a<_�a<#�a<èa<��a<<�a<�a<��a<g�a<.�a<��a<��a<'�a<ĥa<k�a<�a<ͤa<\�a<�a<��a<R�a<ޢa<��a<2�a<��a<n�a<Ҡa<��a<�a<��a<O�a<ўa<��a<�a<��a<)�a<ǜa<Z�a<՛a<��a<��a<��a<,�a<ϙa<U�a<�a<��a<#�a<җa<F�a<�a<��a< �a<�a<d�a<�a<��a<`�a<�a<��a<g�a<��a<͒a<Y�a<>�a<ۑa<��a<\�a<��a<�a<��a<r�a<�a<��a<Ǐa<��a<��a<9�a<A�a<�a<�a<Ɏa<��a<��a<~�a<��a<W�a<[�a<N�a<f�a<a�a<M�a<|�a<b�a<{�a<��a<��a<��a<��a<�  �  �a<��a<�a<T�a<h�a<��a<Ïa<�a<3�a<W�a<��a<�a<�a<P�a<��a<Ցa<&�a<��a<��a<�a<m�a<��a<�a<w�a<̔a<8�a<��a<�a<S�a<��a<'�a<��a<ߗa<[�a<Ҙa<&�a<��a<�a<��a<��a<{�a<�a<\�a<Üa<<�a<��a<'�a<��a<�a<|�a<��a<Z�a<ߠa<\�a<��a<.�a<��a<��a<z�a<�a<5�a<��a<�a<l�a<ѥa<7�a<��a<�a<E�a<��a<��a<X�a<��a<�a<(�a<��a<��a<�a<Z�a<��a<�a<�a<\�a<��a<ëa<�a<4�a<Z�a<��a<��a<׬a<�a<(�a<B�a<��a<��a<��a<׭a<�a<�a<+�a<#�a<.�a<R�a<T�a<d�a<r�a<x�a<��a<��a<��a<��a<��a<��a<��a<��a<w�a<��a<V�a<s�a<R�a<?�a<G�a<0�a<�a<�a<�a<ƭa<ía<��a<|�a<Y�a<3�a<#�a<�a<Ǭa<��a<u�a<Q�a<:�a<�a<ʫa<��a<_�a<4�a<�a<��a<��a<^�a<�a<�a<��a<]�a<�a<ިa<��a<S�a<�a<��a<l�a<�a<Ҧa<b�a<"�a<ͥa<��a<�a<Ǥa<^�a<�a<��a<H�a<�a<}�a<�a<��a<F�a<�a<��a<�a<��a<L�a<˞a<x�a<�a<��a<&�a<��a<G�a<ݛa<v�a<�a<��a<,�a<ʙa<`�a<��a<��a<$�a<��a<`�a<�a<��a<-�a<��a<t�a<�a<��a<_�a<�a<��a<f�a<�a<��a<g�a<�a<ޑa<��a<F�a<,�a<Ӑa<��a<m�a<)�a<�a<ߏa<��a<c�a<O�a<�a<��a<�a<a<��a<��a<��a<~�a<j�a<l�a<d�a<Q�a<K�a<j�a<E�a<v�a<n�a<y�a<��a<��a<ǎa<�  �  юa<�a<�a<M�a<t�a<��a<܏a<�a<@�a<K�a<��a<ѐa<�a<k�a<��a<��a<�a<~�a<��a<�a<r�a<��a<,�a<d�a<ܔa<.�a<��a< �a<G�a<ϖa<�a<��a<�a<]�a<ژa<%�a<Ǚa<��a<��a<�a<r�a<�a<P�a<؜a</�a<Ɲa<#�a<��a<�a<}�a<�a<T�a<�a<:�a<ǡa<*�a<��a<�a<Z�a<�a<0�a<��a<�a<u�a<�a<,�a<��a<�a<W�a<��a<��a<U�a<��a<��a<"�a<��a<��a<�a<_�a<��a<�a<�a<g�a<��a<Ыa<��a<(�a<m�a<{�a<Ŭa<׬a<�a<-�a<>�a<�a<w�a<Эa<��a<��a<��a<	�a<2�a<$�a<d�a<N�a<|�a<l�a<��a<��a<~�a<��a<��a<��a<��a<��a<��a<h�a<��a<V�a<|�a<E�a<I�a<9�a<�a<'�a<�a<��a<��a<��a<��a<o�a<s�a<-�a<0�a<�a<Ӭa<��a<r�a<l�a<�a<�a<��a<��a<b�a<2�a<�a<��a<��a<L�a<+�a<�a<��a<p�a<�a<�a<y�a<Q�a<�a<��a<t�a<�a<�a<Z�a</�a<��a<w�a<�a<��a<r�a<��a<��a<D�a<�a<��a<�a<ˡa<@�a<��a<s�a<&�a<��a<;�a<�a<X�a<�a<��a<5�a<��a<P�a<�a<l�a<�a<��a<>�a<ęa<[�a<��a<u�a<3�a<��a<n�a<�a<��a<3�a<��a<|�a<��a<ɔa<V�a<�a<��a<Z�a<�a<��a<�a<�a<�a<��a<B�a<!�a<��a<��a<K�a<>�a<�a<��a<��a<Y�a<a�a<�a<�a<܎a<ˎa<��a<��a<��a<i�a<u�a<W�a<S�a<[�a<<�a<u�a<D�a<~�a<a�a<��a<��a<��a<؎a<�  �  ֎a<��a<#�a<A�a<|�a<��a<ďa<��a<.�a<h�a<��a<ɐa<�a<b�a<��a<�a<�a<r�a<Βa<"�a<i�a<Ɠa<�a<m�a<֔a<'�a<��a<�a<L�a<��a<�a<��a<�a<O�a<ɘa<A�a<��a<�a<��a<�a<j�a<��a<N�a<a<A�a<��a<0�a<��a<�a<��a< �a<n�a<�a<9�a<��a<(�a<��a<�a<_�a<ߣa<G�a<��a<�a<w�a<Хa<;�a<��a<�a<E�a<��a<��a<H�a<��a<��a<@�a<t�a<ԩa<�a<J�a<��a<ݪa<
�a<S�a<��a<��a<��a<(�a<a�a<��a<��a<�a<�a<:�a<U�a<s�a<��a<��a<��a<�a<��a<�a<6�a<D�a<T�a<]�a<g�a<i�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<}�a<p�a<��a<^�a<O�a<c�a<.�a<�a<�a<��a<�a<ѭa<��a<��a<r�a<[�a<A�a<�a<��a<ެa<��a<|�a<b�a<�a<�a<��a<��a<t�a<D�a<�a<Ӫa<��a<T�a<%�a<کa<��a<Y�a<�a<ڨa<��a<E�a<�a<��a<d�a<�a<��a<s�a<6�a<��a<n�a<�a<��a<]�a<
�a<��a<Q�a<ޢa<��a<#�a<ġa<Z�a<�a<r�a<�a<��a<=�a<�a<]�a<�a<��a<4�a<a<R�a<ܛa<z�a<�a<��a<,�a<��a<W�a<�a<z�a</�a<��a<D�a<��a<��a<�a<ߕa<p�a<�a<��a<W�a<��a<��a<Z�a<�a<��a<h�a<+�a<ޑa<��a<Y�a<�a<Őa<��a<L�a<5�a<��a<��a<��a<y�a<P�a<&�a<�a<؎a<Վa<��a<��a<��a<l�a<o�a<\�a<M�a<q�a<P�a<O�a<p�a<a�a<k�a<��a<��a<��a<͎a<�  �  ��a<�a<0�a<?�a<i�a<��a<a<�a<�a<[�a<��a<�a<�a<R�a<��a<ґa<7�a<��a<��a<�a<Y�a<ѓa<�a<��a<��a</�a<��a<��a<m�a<��a<A�a<v�a<�a<]�a<��a<H�a<��a<+�a<r�a<�a<v�a<�a<l�a<��a<L�a<��a<6�a<��a<�a<��a<�a<c�a<Ҡa<c�a<��a<5�a<��a<��a<��a<٣a<@�a<��a<�a<{�a<ѥa<K�a<�a<��a<:�a<��a< �a<N�a<��a<Ԩa<L�a<x�a<کa<�a<S�a<��a<êa<5�a<I�a<��a<��a<�a<3�a<J�a<��a<��a<�a<��a<&�a<H�a<|�a<��a<��a<�a<�a<��a<,�a<�a<7�a<9�a<f�a<h�a<v�a<~�a<x�a<��a<t�a<��a<��a<��a<��a<t�a<��a<g�a<��a<Q�a<d�a<;�a<4�a<D�a<�a<�a<Эa<ޭa<��a<��a<��a<Y�a<K�a<�a<�a<��a<��a<��a<S�a<G�a<�a<۫a<��a<a�a<2�a<�a<ݪa<��a<g�a<�a<�a<��a<P�a<6�a<Ǩa<��a<6�a<��a<��a<Z�a<&�a<��a<��a<�a<ץa<{�a<�a<פa<O�a<�a<��a<W�a<�a<��a<!�a<��a<O�a<�a<��a<�a<��a<V�a<̞a<��a<�a<��a<�a<��a<V�a<ޛa<��a<��a<��a<!�a<ՙa<c�a<��a<��a<�a<̗a<H�a<��a<��a<'�a<ӕa<V�a<-�a<��a<r�a< �a<��a<e�a<��a<ϒa<f�a<4�a<Αa<��a<L�a<�a<�a<��a<|�a<-�a<��a<��a<��a<l�a<5�a</�a<�a<�a<Ȏa<��a<��a<l�a<��a<]�a<x�a<Z�a<A�a<f�a<E�a<q�a<T�a<��a<u�a<��a<Ɏa<��a<�  �  �a<��a<(�a<J�a<q�a<��a<ˏa<�a<:�a<y�a<��a<ېa<�a<J�a<��a<ݑa<)�a<q�a<Òa<1�a<u�a<��a<�a<r�a<ϔa<6�a<��a<�a<\�a<��a<�a<~�a<�a<o�a<˘a<5�a<��a<%�a<�a<��a<^�a<ӛa<^�a<Ȝa<B�a<��a<)�a<��a<�a<��a<�a<r�a<Ӡa<N�a<��a<%�a<��a<�a<o�a<Уa<M�a<ɤa<�a<z�a<ץa<8�a<��a<��a<I�a<��a<��a<;�a<��a<�a<C�a<��a<˩a<�a<f�a<��a<Ԫa<�a<<�a<��a<��a<��a<5�a<Z�a<��a<��a<߬a<�a<J�a<R�a<g�a<��a<��a<ʭa<٭a<��a<�a<#�a<P�a<^�a<[�a<q�a<t�a<��a<��a<��a<��a<��a<v�a<��a<��a<��a<��a<{�a<n�a<d�a<i�a<@�a<:�a<�a<��a<�a<߭a<֭a<��a<��a<{�a<a�a<:�a<*�a<�a<ʬa<��a<��a<K�a<)�a<��a<ͫa<��a<i�a<R�a<�a<ɪa<��a<Y�a<�a<�a<��a<U�a<%�a<��a<��a<>�a<��a<ħa<e�a<�a<ɦa<��a<�a<Υa<b�a<�a<ɤa<c�a<�a<��a<K�a<�a<��a<!�a<ӡa<^�a<�a<��a<�a<��a<D�a<؞a<m�a<��a<��a<G�a<��a<U�a<�a<w�a<�a<��a<0�a<̙a<W�a<�a<��a<�a<×a<Z�a<�a<��a<9�a<̕a<f�a<�a<��a<e�a<�a<��a<f�a<�a<��a<p�a<%�a<�a<��a<V�a<	�a<Ӑa<��a<`�a<�a<��a<Џa<��a<��a<[�a<$�a<�a<�a<ˎa<��a<��a<��a<��a<O�a<U�a<`�a<N�a<f�a<Y�a<\�a<g�a<��a<{�a<��a<��a<��a<�  �  Ɏa<�a< �a<@�a<��a<��a<ҏa<�a<%�a<K�a<��a<ѐa<�a<`�a<��a<��a<(�a<�a<ƒa< �a<d�a<��a<$�a<h�a<��a<�a<��a<�a<D�a<Ֆa<�a<��a<�a<H�a<Șa<0�a<��a<�a<��a<��a<��a<��a<F�a<ۜa<+�a<��a<$�a<��a<�a<o�a<�a<U�a<�a<?�a<ӡa<'�a<��a<�a<c�a<�a<3�a<��a<��a<j�a<إa<0�a<��a<�a<Y�a<��a<	�a<c�a<��a<��a<#�a<��a<ũa<�a<J�a<��a<�a<�a<p�a<��a<ƫa<�a<�a<m�a<��a<¬a<Ϭa<��a<�a<M�a<}�a<��a<ŭa<��a<�a<�a<�a<6�a<%�a<F�a<M�a<r�a<l�a<��a<��a<��a<��a<x�a<��a<��a<��a<��a<i�a<w�a<k�a<b�a<?�a<S�a<B�a<&�a<5�a<�a<�a<έa<��a<��a<s�a<i�a<,�a<�a<�a<۬a<��a<��a<a�a<�a<�a<̫a<��a<m�a<"�a<��a<��a<��a<O�a</�a<Ωa<��a<`�a<�a<��a<��a<V�a<��a<��a<c�a<�a<æa<]�a<.�a<ǥa<��a</�a<��a<v�a<��a<��a<E�a<�a<}�a<�a<��a<A�a<��a<x�a<2�a<��a<>�a<�a<a�a<�a<��a<�a<��a<E�a<�a<o�a<�a<��a<@�a<��a<l�a<�a<��a<4�a<��a<O�a<�a<��a<�a<��a<~�a<
�a<Ӕa<Z�a<�a<��a<K�a<�a<��a<}�a<�a<Бa<��a<Q�a<�a<ːa<��a<M�a<0�a<�a<a<��a<Z�a<B�a<�a<�a<܎a<֎a<��a<��a<��a<]�a<��a<g�a<_�a<b�a<<�a<V�a<Y�a<e�a<[�a<��a<��a<��a<�a<�  �  Ȏa<�a<+�a<G�a<j�a<��a<ӏa<�a<<�a<]�a<��a<ѐa<�a<P�a<��a<ڑa<&�a<}�a<͒a<�a<��a<ϓa<!�a<^�a<˔a<(�a<��a<�a<<�a<��a<�a<��a<��a<]�a<Ҙa<=�a<��a<�a<��a<�a<]�a<қa<@�a<ۜa<?�a<��a<�a<��a<�a<��a<�a<m�a<�a<A�a<��a<'�a<��a<�a<k�a<�a<J�a<��a<&�a<��a<إa<.�a<��a<�a<Z�a<��a<�a<;�a<��a<�a<9�a<��a<өa<�a<^�a<��a<۪a<
�a<E�a<s�a<«a<�a<%�a<Z�a<z�a<��a<�a<�a</�a<Y�a<{�a<��a<��a<ԭa<�a<��a<�a<5�a<;�a<^�a<o�a<t�a<h�a<w�a<��a<��a<��a<w�a<��a<��a<��a<��a<~�a<��a<w�a<m�a<R�a<G�a<2�a<�a<�a<�a<��a<ڭa<��a<��a<m�a<j�a<K�a<+�a<�a<ܬa<��a<~�a<Q�a<1�a<��a<ʫa<��a<t�a<4�a<�a<ܪa<��a<E�a<�a<۩a<��a<`�a<�a<̨a<}�a<G�a<�a<��a<l�a<�a<Ӧa<q�a< �a<��a<a�a<�a<��a<v�a<	�a<��a<A�a<�a<��a<6�a<ȡa<X�a<��a<{�a<�a<��a<F�a<؞a<i�a<�a<��a<3�a<Ҝa<[�a<�a<n�a<�a<��a<A�a<��a<E�a<��a<y�a<$�a<��a<d�a<��a<��a<1�a<͕a<m�a<�a<��a<C�a<�a<��a<W�a<�a<��a<x�a<4�a<�a<��a<]�a<�a<ѐa<��a<j�a<'�a<��a<a<��a<o�a<Z�a<7�a<�a<؎a<a<��a<��a<��a<]�a<d�a<Q�a<P�a<S�a<R�a<b�a<e�a<p�a<n�a<��a<��a<��a<��a<�  �  ��a<�a<�a<L�a<p�a<��a<ʏa<�a<&�a<f�a<��a<ܐa<!�a<G�a<��a<ӑa<:�a<q�a<��a<�a<a�a<��a<�a<y�a<Ԕa<8�a<u�a<�a<r�a<��a<4�a<��a<�a<b�a<��a<%�a<��a<�a<��a<�a<|�a<�a<d�a<��a<3�a<��a</�a<��a<�a<u�a<�a<m�a<ɠa<]�a<��a<.�a<��a<�a<��a<ǣa<I�a<��a<�a<n�a<�a<A�a<��a<�a<<�a<��a<
�a<[�a<��a<�a<5�a<��a<��a<�a<\�a<��a<Ѫa<0�a<X�a<��a<ëa<�a<0�a<a�a<��a<��a<լa<��a</�a<N�a<c�a<��a<��a<�a<ۭa<�a< �a<$�a<D�a<E�a<M�a<i�a<��a<�a<��a<z�a<��a<��a<��a<��a<��a<~�a<��a<v�a<a�a<a�a<b�a<=�a<E�a<7�a<�a<�a<ۭa<��a<��a<��a<��a<`�a</�a<�a<��a<ˬa<��a<��a<G�a<N�a<�a<ޫa<��a<g�a<9�a<��a<��a<��a<`�a<#�a<�a<��a<S�a<;�a<ިa<��a<C�a<��a<��a<Z�a<�a<��a<s�a<�a<�a<��a<)�a<Ϥa<X�a<��a<��a<P�a<�a<}�a<�a<��a<Y�a<ܠa<��a<�a<��a<R�a<ٞa<��a<�a<��a<%�a<��a<I�a<�a<��a<�a<��a<#�a<љa<m�a<�a<��a<�a<��a<S�a<�a<��a</�a<ɕa<d�a<(�a<��a<u�a<�a<��a<b�a<�a<ɒa<q�a<�a<ϑa<��a<R�a<�a<�a<��a<�a<!�a<�a<ԏa<��a<y�a<A�a<�a<�a<�a<Ɏa<��a<��a<~�a<��a<o�a<m�a<m�a<K�a<b�a<T�a<P�a<d�a<~�a<x�a<��a<��a<ʎa<�  �  Ȏa<�a<+�a<G�a<j�a<��a<ӏa<�a<<�a<]�a<��a<ѐa<�a<P�a<��a<ڑa<&�a<}�a<͒a<�a<��a<ϓa<!�a<^�a<˔a<(�a<��a<�a<<�a<��a<�a<��a<��a<]�a<Ҙa<=�a<��a<�a<��a<�a<]�a<қa<@�a<ۜa<?�a<��a<�a<��a<�a<��a<�a<m�a<�a<A�a<��a<'�a<��a<�a<k�a<�a<J�a<��a<&�a<��a<إa<.�a<��a<�a<Z�a<��a<�a<;�a<��a<�a<9�a<��a<өa<�a<^�a<��a<۪a<
�a<E�a<s�a<«a<�a<%�a<Z�a<z�a<��a<�a<�a</�a<Y�a<{�a<��a<��a<ԭa<�a<��a<�a<5�a<;�a<^�a<o�a<t�a<h�a<w�a<��a<��a<��a<w�a<��a<��a<��a<��a<~�a<��a<w�a<m�a<R�a<G�a<2�a<�a<�a<�a<��a<ڭa<��a<��a<m�a<j�a<K�a<+�a<�a<ܬa<��a<~�a<Q�a<1�a<��a<ʫa<��a<t�a<4�a<�a<ܪa<��a<E�a<�a<۩a<��a<`�a<�a<̨a<}�a<G�a<�a<��a<l�a<�a<Ӧa<q�a< �a<��a<a�a<�a<��a<v�a<	�a<��a<A�a<�a<��a<6�a<ȡa<X�a<��a<{�a<�a<��a<F�a<؞a<i�a<�a<��a<3�a<Ҝa<[�a<�a<n�a<�a<��a<A�a<��a<E�a<��a<y�a<$�a<��a<d�a<��a<��a<1�a<͕a<m�a<�a<��a<C�a<�a<��a<W�a<�a<��a<x�a<4�a<�a<��a<]�a<�a<ѐa<��a<j�a<'�a<��a<a<��a<o�a<Z�a<7�a<�a<؎a<a<��a<��a<��a<]�a<d�a<Q�a<P�a<S�a<R�a<b�a<e�a<p�a<n�a<��a<��a<��a<��a<�  �  Ɏa<�a< �a<@�a<��a<��a<ҏa<�a<%�a<K�a<��a<ѐa<�a<`�a<��a<��a<(�a<�a<ƒa< �a<d�a<��a<$�a<h�a<��a<�a<��a<�a<D�a<Ֆa<�a<��a<�a<H�a<Șa<0�a<��a<�a<��a<��a<��a<��a<F�a<ۜa<+�a<��a<$�a<��a<�a<o�a<�a<U�a<�a<?�a<ӡa<'�a<��a<�a<c�a<�a<3�a<��a<��a<j�a<إa<0�a<��a<�a<Y�a<��a<	�a<c�a<��a<��a<#�a<��a<ũa<�a<J�a<��a<�a<�a<p�a<��a<ƫa<�a<�a<m�a<��a<¬a<Ϭa<��a<�a<M�a<}�a<��a<ŭa<��a<�a<�a<�a<6�a<%�a<F�a<M�a<r�a<l�a<��a<��a<��a<��a<x�a<��a<��a<��a<��a<i�a<w�a<k�a<b�a<?�a<S�a<B�a<&�a<5�a<�a<�a<έa<��a<��a<s�a<i�a<,�a<�a<�a<۬a<��a<��a<a�a<�a<�a<̫a<��a<m�a<"�a<��a<��a<��a<O�a</�a<Ωa<��a<`�a<�a<��a<��a<V�a<��a<��a<c�a<�a<æa<]�a<.�a<ǥa<��a</�a<��a<v�a<��a<��a<E�a<�a<}�a<�a<��a<A�a<��a<x�a<2�a<��a<>�a<�a<a�a<�a<��a<�a<��a<E�a<�a<o�a<�a<��a<@�a<��a<l�a<�a<��a<4�a<��a<O�a<�a<��a<�a<��a<~�a<
�a<Ӕa<Z�a<�a<��a<K�a<�a<��a<}�a<�a<Бa<��a<Q�a<�a<ːa<��a<M�a<0�a<�a<a<��a<Z�a<B�a<�a<�a<܎a<֎a<��a<��a<��a<]�a<��a<g�a<_�a<b�a<<�a<V�a<Y�a<e�a<[�a<��a<��a<��a<�a<�  �  �a<��a<(�a<J�a<q�a<��a<ˏa<�a<:�a<y�a<��a<ېa<�a<J�a<��a<ݑa<)�a<q�a<Òa<1�a<u�a<��a<�a<r�a<ϔa<6�a<��a<�a<\�a<��a<�a<~�a<�a<o�a<˘a<5�a<��a<%�a<�a<��a<^�a<ӛa<^�a<Ȝa<B�a<��a<)�a<��a<�a<��a<�a<r�a<Ӡa<N�a<��a<%�a<��a<�a<o�a<Уa<M�a<ɤa<�a<z�a<ץa<8�a<��a<��a<I�a<��a<��a<;�a<��a<�a<C�a<��a<˩a<�a<f�a<��a<Ԫa<�a<<�a<��a<��a<��a<5�a<Z�a<��a<��a<߬a<�a<J�a<R�a<g�a<��a<��a<ʭa<٭a<��a<�a<#�a<P�a<^�a<[�a<q�a<t�a<��a<��a<��a<��a<��a<v�a<��a<��a<��a<��a<{�a<n�a<d�a<i�a<@�a<:�a<�a<��a<�a<߭a<֭a<��a<��a<{�a<a�a<:�a<*�a<�a<ʬa<��a<��a<K�a<)�a<��a<ͫa<��a<i�a<R�a<�a<ɪa<��a<Y�a<�a<�a<��a<U�a<%�a<��a<��a<>�a<��a<ħa<e�a<�a<ɦa<��a<�a<Υa<b�a<�a<ɤa<c�a<�a<��a<K�a<�a<��a<!�a<ӡa<^�a<�a<��a<�a<��a<D�a<؞a<m�a<��a<��a<G�a<��a<U�a<�a<w�a<�a<��a<0�a<̙a<W�a<�a<��a<�a<×a<Z�a<�a<��a<9�a<̕a<f�a<�a<��a<e�a<�a<��a<f�a<�a<��a<p�a<%�a<�a<��a<V�a<	�a<Ӑa<��a<`�a<�a<��a<Џa<��a<��a<[�a<$�a<�a<�a<ˎa<��a<��a<��a<��a<O�a<U�a<`�a<N�a<f�a<Y�a<\�a<g�a<��a<{�a<��a<��a<��a<�  �  ��a<�a<0�a<?�a<i�a<��a<a<�a<�a<[�a<��a<�a<�a<R�a<��a<ґa<7�a<��a<��a<�a<Y�a<ѓa<�a<��a<��a</�a<��a<��a<m�a<��a<A�a<v�a<�a<]�a<��a<H�a<��a<+�a<r�a<�a<v�a<�a<l�a<��a<L�a<��a<6�a<��a<�a<��a<�a<c�a<Ҡa<c�a<��a<5�a<��a<��a<��a<٣a<@�a<��a<�a<{�a<ѥa<K�a<�a<��a<:�a<��a< �a<N�a<��a<Ԩa<L�a<x�a<کa<�a<S�a<��a<êa<5�a<I�a<��a<��a<�a<3�a<J�a<��a<��a<�a<��a<&�a<H�a<|�a<��a<��a<�a<�a<��a<,�a<�a<7�a<9�a<f�a<h�a<v�a<~�a<x�a<��a<t�a<��a<��a<��a<��a<t�a<��a<g�a<��a<Q�a<d�a<;�a<4�a<D�a<�a<�a<Эa<ޭa<��a<��a<��a<Y�a<K�a<�a<�a<��a<��a<��a<S�a<G�a<�a<۫a<��a<a�a<2�a<�a<ݪa<��a<g�a<�a<�a<��a<P�a<6�a<Ǩa<��a<6�a<��a<��a<Z�a<&�a<��a<��a<�a<ץa<{�a<�a<פa<O�a<�a<��a<W�a<�a<��a<!�a<��a<O�a<�a<��a<�a<��a<V�a<̞a<��a<�a<��a<�a<��a<V�a<ޛa<��a<��a<��a<!�a<ՙa<c�a<��a<��a<�a<̗a<H�a<��a<��a<'�a<ӕa<V�a<-�a<��a<r�a< �a<��a<e�a<��a<ϒa<f�a<4�a<Αa<��a<L�a<�a<�a<��a<|�a<-�a<��a<��a<��a<l�a<5�a</�a<�a<�a<Ȏa<��a<��a<l�a<��a<]�a<x�a<Z�a<A�a<f�a<E�a<q�a<T�a<��a<u�a<��a<Ɏa<��a<�  �  ֎a<��a<#�a<A�a<|�a<��a<ďa<��a<.�a<h�a<��a<ɐa<�a<b�a<��a<�a<�a<r�a<Βa<"�a<i�a<Ɠa<�a<m�a<֔a<'�a<��a<�a<L�a<��a<�a<��a<�a<O�a<ɘa<A�a<��a<�a<��a<�a<j�a<��a<N�a<a<A�a<��a<0�a<��a<�a<��a< �a<n�a<�a<9�a<��a<(�a<��a<�a<_�a<ߣa<G�a<��a<�a<w�a<Хa<;�a<��a<�a<E�a<��a<��a<H�a<��a<��a<@�a<t�a<ԩa<�a<J�a<��a<ݪa<
�a<S�a<��a<��a<��a<(�a<a�a<��a<��a<�a<�a<:�a<U�a<s�a<��a<��a<��a<�a<��a<�a<6�a<D�a<T�a<]�a<g�a<i�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<}�a<p�a<��a<^�a<O�a<c�a<.�a<�a<�a<��a<�a<ѭa<��a<��a<r�a<[�a<A�a<�a<��a<ެa<��a<|�a<b�a<�a<�a<��a<��a<t�a<D�a<�a<Ӫa<��a<T�a<%�a<کa<��a<Y�a<�a<ڨa<��a<E�a<�a<��a<d�a<�a<��a<s�a<6�a<��a<n�a<�a<��a<]�a<
�a<��a<Q�a<ޢa<��a<#�a<ġa<Z�a<�a<r�a<�a<��a<=�a<�a<]�a<�a<��a<4�a<a<R�a<ܛa<z�a<�a<��a<,�a<��a<W�a<�a<z�a</�a<��a<D�a<��a<��a<�a<ߕa<p�a<�a<��a<W�a<��a<��a<Z�a<�a<��a<h�a<+�a<ޑa<��a<Y�a<�a<Őa<��a<L�a<5�a<��a<��a<��a<y�a<P�a<&�a<�a<؎a<Վa<��a<��a<��a<l�a<o�a<\�a<M�a<q�a<P�a<O�a<p�a<a�a<k�a<��a<��a<��a<͎a<�  �  юa<�a<�a<M�a<t�a<��a<܏a<�a<@�a<K�a<��a<ѐa<�a<k�a<��a<��a<�a<~�a<��a<�a<r�a<��a<,�a<d�a<ܔa<.�a<��a< �a<G�a<ϖa<�a<��a<�a<]�a<ژa<%�a<Ǚa<��a<��a<�a<r�a<�a<P�a<؜a</�a<Ɲa<#�a<��a<�a<}�a<�a<T�a<�a<:�a<ǡa<*�a<��a<�a<Z�a<�a<0�a<��a<�a<u�a<�a<,�a<��a<�a<W�a<��a<��a<U�a<��a<��a<"�a<��a<��a<�a<_�a<��a<�a<�a<g�a<��a<Ыa<��a<(�a<m�a<{�a<Ŭa<׬a<�a<-�a<>�a<�a<w�a<Эa<��a<��a<��a<	�a<2�a<$�a<d�a<N�a<|�a<l�a<��a<��a<~�a<��a<��a<��a<��a<��a<��a<h�a<��a<V�a<|�a<E�a<I�a<9�a<�a<'�a<�a<��a<��a<��a<��a<o�a<s�a<-�a<0�a<�a<Ӭa<��a<r�a<l�a<�a<�a<��a<��a<b�a<2�a<�a<��a<��a<L�a<+�a<�a<��a<p�a<�a<�a<y�a<Q�a<�a<��a<t�a<�a<�a<Z�a</�a<��a<w�a<�a<��a<r�a<��a<��a<D�a<�a<��a<�a<ˡa<@�a<��a<s�a<&�a<��a<;�a<�a<X�a<�a<��a<5�a<��a<P�a<�a<l�a<�a<��a<>�a<ęa<[�a<��a<u�a<3�a<��a<n�a<�a<��a<3�a<��a<|�a<��a<ɔa<V�a<�a<��a<Z�a<�a<��a<�a<�a<�a<��a<B�a<!�a<��a<��a<K�a<>�a<�a<��a<��a<Y�a<a�a<�a<�a<܎a<ˎa<��a<��a<��a<i�a<u�a<W�a<S�a<[�a<<�a<u�a<D�a<~�a<a�a<��a<��a<��a<؎a<�  �  �a<��a<�a<T�a<h�a<��a<Ïa<�a<3�a<W�a<��a<�a<�a<P�a<��a<Ցa<&�a<��a<��a<�a<m�a<��a<�a<w�a<̔a<8�a<��a<�a<S�a<��a<'�a<��a<ߗa<[�a<Ҙa<&�a<��a<�a<��a<��a<{�a<�a<\�a<Üa<<�a<��a<'�a<��a<�a<|�a<��a<Z�a<ߠa<\�a<��a<.�a<��a<��a<z�a<�a<5�a<��a<�a<l�a<ѥa<7�a<��a<�a<E�a<��a<��a<X�a<��a<�a<(�a<��a<��a<�a<Z�a<��a<�a<�a<\�a<��a<ëa<�a<4�a<Z�a<��a<��a<׬a<�a<(�a<B�a<��a<��a<��a<׭a<�a<�a<+�a<#�a<.�a<R�a<T�a<d�a<r�a<x�a<��a<��a<��a<��a<��a<��a<��a<��a<w�a<��a<V�a<s�a<R�a<?�a<G�a<0�a<�a<�a<�a<ƭa<ía<��a<|�a<Y�a<3�a<#�a<�a<Ǭa<��a<u�a<Q�a<:�a<�a<ʫa<��a<_�a<4�a<�a<��a<��a<^�a<�a<�a<��a<]�a<�a<ިa<��a<S�a<�a<��a<l�a<�a<Ҧa<b�a<"�a<ͥa<��a<�a<Ǥa<^�a<�a<��a<H�a<�a<}�a<�a<��a<F�a<�a<��a<�a<��a<L�a<˞a<x�a<�a<��a<&�a<��a<G�a<ݛa<v�a<�a<��a<,�a<ʙa<`�a<��a<��a<$�a<��a<`�a<�a<��a<-�a<��a<t�a<�a<��a<_�a<�a<��a<f�a<�a<��a<g�a<�a<ޑa<��a<F�a<,�a<Ӑa<��a<m�a<)�a<�a<ߏa<��a<c�a<O�a<�a<��a<�a<a<��a<��a<��a<~�a<j�a<l�a<d�a<Q�a<K�a<j�a<E�a<v�a<n�a<y�a<��a<��a<ǎa<�  �  �a<��a<)�a<?�a<j�a<��a<��a<�a<�a<��a<��a<ːa<�a<B�a<��a<Αa<<�a<_�a<ǒa<*�a<`�a<ۓa<��a<��a<��a</�a<��a<�a<Z�a<��a<�a<|�a<�a<Y�a<͘a<P�a<��a<-�a<��a<��a<f�a<՛a<b�a<��a<S�a<��a<1�a<��a<�a<��a<�a<��a<��a<V�a<��a<+�a<��a<��a<��a<£a<Z�a<��a<�a<~�a<ɥa<A�a<��a<�a<E�a<��a<�a<A�a<��a<�a<R�a<v�a<�a<�a<M�a<��a<Ѫa<�a<A�a<��a<ǫa<��a<5�a<G�a<��a<��a<��a<�a<8�a<Y�a<Z�a<��a<��a<ܭa<حa<�a<�a<�a<^�a<<�a<x�a<X�a<z�a<~�a<x�a<��a<��a<��a<�a<��a<��a<��a<��a<n�a<��a<_�a<_�a<Z�a<*�a<"�a<��a<�a<�a<׭a<��a<��a<��a<H�a<X�a<�a<�a<Ȭa<��a<��a<C�a<<�a<�a<�a<��a<n�a<L�a<��a<�a<y�a<j�a<�a<�a<��a<_�a<#�a<èa<��a<<�a<�a<��a<g�a<.�a<��a<��a<'�a<ĥa<k�a<�a<ͤa<\�a<�a<��a<R�a<ޢa<��a<2�a<��a<n�a<Ҡa<��a<�a<��a<O�a<ўa<��a<�a<��a<)�a<ǜa<Z�a<՛a<��a<��a<��a<,�a<ϙa<U�a<�a<��a<#�a<җa<F�a<�a<��a< �a<�a<d�a<�a<��a<`�a<�a<��a<g�a<��a<͒a<Y�a<>�a<ۑa<��a<\�a<��a<�a<��a<r�a<�a<��a<Ǐa<��a<��a<9�a<A�a<�a<�a<Ɏa<��a<��a<~�a<��a<W�a<[�a<N�a<f�a<a�a<M�a<|�a<b�a<{�a<��a<��a<��a<��a<�  �  ގa<�a< �a<G�a<s�a<��a<��a<�a<�a<Y�a<��a<ΐa<&�a<U�a<��a<�a<9�a<m�a<˒a<	�a<P�a<͓a<�a<w�a<Δa<.�a<��a<��a<R�a<ʖa<0�a<��a<��a<]�a<��a<8�a<��a<�a<�a<��a<��a<�a<W�a<ɜa<>�a<��a</�a<��a<�a<��a<��a<h�a<Ӡa<N�a<ȡa<(�a<��a<�a<x�a<ԣa<E�a<��a<�a<y�a<֥a<>�a<��a<�a<L�a<��a<��a<k�a<��a<�a<7�a<��a<Ωa<�a<W�a<��a<Ԫa<#�a<i�a<��a<ɫa<��a<-�a<Z�a<��a<��a<�a<��a<�a<U�a<g�a<��a<��a<ȭa<�a<�a<�a<"�a<8�a<1�a<h�a<]�a<{�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<t�a<p�a<\�a<X�a<M�a<3�a<@�a<"�a<��a<�a<έa<��a<��a<��a<R�a<K�a<��a<�a<Ϭa<��a<��a<V�a<'�a<��a<ݫa<��a<r�a<+�a<�a<٪a<��a<^�a<�a<�a<��a<f�a<�a<�a<��a<A�a<�a<��a<Z�a<�a<æa<p�a<�a<Υa<��a<#�a<��a<d�a<�a<��a<Q�a<�a<��a<&�a<��a<S�a<�a<��a<(�a<��a<D�a<�a<v�a<��a<��a<�a<��a<U�a<�a<~�a<�a<��a<2�a<˙a<a�a<�a<��a<�a<��a<R�a<�a<��a<*�a<Еa<g�a<�a<˔a<]�a<�a<��a<_�a<
�a<��a<n�a</�a<ʑa<��a<Y�a<	�a<�a<��a<]�a<,�a<�a<ďa<��a<m�a<-�a<1�a<��a<�a<юa<��a<��a<��a<t�a<v�a<z�a<V�a<T�a<U�a<S�a<^�a<_�a<t�a<��a<��a<Ŏa<ӎa<�  �  юa<�a<�a<[�a<e�a<��a<͏a<��a<K�a<]�a<��a<ېa<��a<T�a<��a<ޑa<�a<��a<Ȓa<!�a<��a<��a<)�a<a�a<Дa<6�a<��a<�a<A�a<��a<	�a<��a<�a<o�a<͘a<'�a<��a<�a<��a<��a<[�a<қa<H�a<֜a<6�a<ŝa<�a<��a<�a<��a<�a<c�a<�a<9�a<��a<$�a<��a<��a<\�a<�a<=�a<Ĥa<�a<q�a<�a<&�a<��a<�a<P�a<��a<�a<=�a<��a<��a<,�a<��a<éa<�a<o�a<��a<�a<�a<K�a<z�a<��a<��a<,�a<b�a<u�a<Ǭa<ˬa<�a<=�a<O�a<��a<{�a<��a<ía<�a<�a<�a<7�a<4�a<k�a<J�a<k�a<}�a<n�a<��a<��a<��a<��a<��a<z�a<��a<��a<��a<��a<U�a<s�a<_�a<H�a<B�a<�a<�a<�a<��a<ƭa<ʭa<��a<�a<d�a<&�a<:�a<�a<ܬa<��a<h�a<U�a<$�a<��a<��a<��a<o�a<B�a<�a<��a<��a<H�a<�a<�a<��a<b�a<
�a<Ψa<z�a<V�a<��a<ħa<g�a<�a<ۦa<g�a<,�a<åa<`�a<�a<��a<q�a<��a<��a<7�a<��a<��a<"�a<סa<O�a<��a<r�a<�a<��a<>�a<Ӟa<Z�a<�a<��a<C�a<ɜa<L�a<�a<e�a<�a<��a<7�a<��a<J�a<�a<z�a<0�a<��a<j�a<�a<��a<B�a<��a<~�a<��a<��a<J�a< �a<��a<^�a<�a<��a<��a<�a<��a<��a<S�a<!�a<��a<��a<Y�a<*�a<�a<Ǐa<��a<i�a<g�a<�a<�a<�a<��a<Îa<��a<��a<e�a<f�a<J�a<^�a<[�a<X�a<l�a<C�a<v�a<{�a<��a<��a<��a<��a<�  �  ��a<�a<�a<C�a<n�a<��a<Џa<ߏa<$�a<M�a<��a<Ԑa<�a<^�a<��a<�a<'�a<s�a<��a<�a<a�a<��a<*�a<s�a<Ӕa<%�a<��a<��a<f�a<ǖa< �a<��a<�a<[�a<ǘa<?�a<��a<�a<��a<�a<t�a<��a<d�a<ќa<0�a<��a<"�a<��a<
�a<i�a<�a<Z�a<۠a<L�a<áa</�a<��a<�a<q�a<ޣa<5�a<��a<��a<i�a<�a<4�a<��a<�a<O�a<��a<�a<U�a<��a<��a<6�a<��a<ϩa<�a<V�a<��a<�a<�a<b�a<��a<ͫa<�a<#�a<b�a<��a<Ȭa<Ǭa<��a<�a<A�a<p�a<��a<��a<Эa<�a<��a<�a<&�a<'�a<D�a<E�a<n�a<��a<z�a<��a<x�a<��a<��a<��a<��a<��a<��a<�a<s�a<u�a<_�a<V�a<H�a<D�a<#�a<'�a<�a<��a<��a<��a<��a<��a<g�a<$�a<�a<�a<ʬa<��a<{�a<_�a<0�a<�a<˫a<��a<_�a<)�a<��a<��a<��a<[�a<"�a<ةa<��a<h�a</�a<�a<��a<S�a<��a<��a<a�a<�a<Ŧa<p�a<)�a<ԥa<x�a<-�a<Ϥa<l�a<��a<��a<C�a<��a<�a<�a<��a<F�a<�a<��a<#�a<��a<K�a<�a<o�a<�a<��a<�a<��a<D�a<�a<t�a<�a<��a<5�a<әa<q�a<��a<��a<+�a<��a<S�a<�a<��a<)�a<��a<v�a<�a<Ĕa<r�a<�a<��a<U�a<�a<��a<��a<�a<Бa<��a<E�a<�a<Ԑa<��a<f�a<4�a<��a<ˏa<��a<\�a<@�a<�a<�a<�a<Ŏa<��a<��a<��a<��a<��a<[�a<b�a<Z�a<S�a<R�a<c�a<b�a<s�a<��a<��a<��a<؎a<�  �  3�a<\�a<��a<��a<ҏa<��a<!�a<}�a<~�a<Ԑa<�a<&�a<h�a<��a<�a<,�a<��a<��a<?�a<r�a<Гa<7�a<d�a<Ҕa<.�a<��a<�a<H�a<��a<�a<p�a<Ηa<W�a<��a<�a<��a<�a<��a<ؚa<O�a<��a<&�a<��a<�a<��a<�a<~�a<�a<d�a<��a<7�a<ՠa<�a<��a<�a<��a<��a<2�a<��a<�a<��a<�a<}�a<ʥa<�a<��a<ݦa<;�a<��a<�a<-�a<{�a<�a<*�a<��a<��a<�a<U�a<��a<��a<�a<^�a<��a<ūa<�a<B�a<l�a<��a<֬a<�a<?�a<^�a<n�a<��a<��a<ܭa<�a<(�a<4�a<3�a<P�a<x�a<��a<��a<Ȯa<��a<��a<ʮa<Ǯa<߮a<ծa<ͮa<ͮa<̮a<Үa<ˮa<�a<��a<Юa<��a<��a<��a<x�a<f�a<O�a<:�a<-�a<$�a<��a<�a<ía<��a<��a<W�a<S�a<,�a<�a<��a<��a<��a<3�a<�a<ʫa<ѫa<��a<U�a<0�a<ͪa<��a<j�a<!�a<�a<��a<T�a<�a<Ѩa<~�a<S�a<��a<��a<h�a<��a<ۦa<b�a<�a<��a<T�a<�a<��a<[�a<�a<��a<(�a<Ԣa<��a<��a<��a<-�a<Ϡa<I�a<�a<��a<�a<��a<?�a<�a<n�a<2�a<��a<*�a<ћa<^�a<��a<��a<�a<��a<0�a<�a<o�a<-�a<��a<P�a<��a<�a<:�a<��a<k�a<��a<��a<[�a<�a<��a<l�a< �a<��a<��a<K�a<�a<ёa<V�a<7�a<�a<֐a<��a<E�a<�a<�a<�a<��a<��a<c�a<?�a<-�a<	�a<�a<�a<ˎa<��a<��a<��a<��a<ӎa<��a<׎a<��a<�a<�a<�a<�a<�a<�  �  I�a<^�a<y�a<��a<ˏa<�a<%�a<E�a<}�a<��a<��a<:�a<��a<��a<�a<<�a<��a<Ԓa<#�a<[�a<ēa<	�a<x�a<ϔa<+�a<��a<�a<H�a<��a<!�a<v�a<�a<G�a<��a<!�a<��a<��a<o�a<�a<Z�a<ța<P�a<��a<�a<��a<�a<r�a<�a<O�a<ɟa<.�a<��a< �a<��a<�a<k�a<բa<T�a<Σa<�a<��a<ܤa<R�a<��a<'�a<y�a<�a<3�a<��a<�a<Y�a<��a<�a<:�a<�a<ĩa<�a<\�a<��a<ުa<-�a<^�a<��a<�a<�a<>�a<r�a<��a<Ϭa<�a<�a<J�a<[�a<��a<��a<�a<��a<�a<*�a<R�a<g�a<j�a<}�a<��a<��a<��a<Ʈa<®a<ծa<̮a<֮a<ޮa<�a<خa<�a<ɮa<ήa<��a<��a<��a<��a<��a<��a<o�a<n�a<P�a</�a<�a<�a<�a<ͭa<��a<s�a<V�a<4�a<�a<��a<٬a<��a<c�a<C�a<+�a<�a<��a<h�a<H�a<�a<�a<��a<g�a<*�a<�a<��a<r�a</�a<֨a<��a<C�a<��a<��a<c�a<�a<��a<j�a<�a<¥a<�a<�a<��a<K�a<��a<��a<:�a<��a<c�a<�a<��a<2�a<�a<o�a<��a<��a<.�a<ўa<M�a<�a<b�a<�a<��a<=�a<ěa<d�a<�a<��a<"�a<˙a<P�a<�a<�a<�a<��a<O�a<�a<��a<#�a<ӕa<j�a<�a<˔a<c�a<�a<��a<n�a<�a<Ԓa<r�a<7�a<ܑa<��a<q�a<I�a<��a<��a<��a<e�a<3�a<�a<ʏa<��a<r�a<_�a<N�a<%�a<�a<�a<�a<܎a<ݎa<��a<̎a<��a<��a<��a<Ďa<a<׎a<ގa<�a<�a<6�a<�  �  2�a<e�a<}�a<��a<��a<��a<2�a<T�a<��a<��a<��a<-�a<k�a<��a<��a<I�a<y�a<Ԓa<"�a<u�a<�a<�a<��a<��a<�a<��a<�a<C�a<��a<�a<h�a<��a<7�a<��a<+�a<��a<�a<`�a<�a<P�a<��a</�a<��a<%�a<��a<�a<^�a<��a<[�a<ߟa<\�a<��a<*�a<��a<�a<}�a<�a<Y�a<��a<*�a<��a<�a<n�a<��a<-�a<f�a<�a<7�a<��a<ߧa<6�a<��a<ܨa<@�a<q�a<ܩa<�a<_�a<��a<ͪa<6�a<N�a<��a<ūa<�a<D�a<t�a<��a<��a<�a<�a<s�a<{�a<��a<��a<ǭa<�a<�a<9�a<?�a<P�a<s�a<��a<��a<��a<��a<��a<��a<�a<Ϯa<�a<Ȯa<׮a<ͮa<�a<ɮa<Ǯa<ծa<��a<��a<��a<��a<��a<`�a<[�a<8�a<6�a<�a<�a<ʭa<ía<��a<��a<��a<=�a<�a<�a<��a<��a<x�a<Q�a<�a<�a<��a<��a<r�a<�a<�a<��a<[�a<.�a<�a<��a<T�a<�a<ɨa<��a<3�a<�a<��a<\�a<!�a<��a<n�a<�a<��a<^�a<��a<��a<N�a<�a<y�a<>�a<ˢa<y�a<�a<��a<<�a<��a<l�a<�a<��a<2�a<��a<W�a<�a<��a<#�a<��a<D�a<��a<i�a<�a<��a<�a<��a<>�a<טa<��a<�a<��a<H�a<�a<��a<�a<ݕa<[�a<�a<��a<Y�a<�a<��a<g�a<�a<�a<w�a<`�a<��a<��a<w�a<"�a<�a<Ða<��a<R�a<�a<��a<Џa<͏a<��a<l�a<G�a<�a<#�a<��a<��a<Ǝa<Ȏa<��a<Ȏa<��a<��a<̎a<��a<َa<׎a<؎a<�a<��a<$�a<�  �  E�a<b�a<��a<��a<Ϗa< �a<�a<k�a<s�a<��a<�a<3�a<w�a<��a<��a<6�a<��a<Вa<*�a<d�a<��a<#�a<g�a<הa<1�a<��a<�a<L�a<��a<!�a<��a<җa<A�a<��a< �a<��a<��a<{�a<ۚa<P�a<ԛa<D�a<��a<�a<��a<�a<{�a<�a<T�a<џa<'�a<��a<0�a<��a<�a<t�a<�a<L�a<��a<)�a<��a<٤a<T�a<��a<�a<��a<�a<4�a<��a<��a<M�a<��a<�a<.�a<��a<ɩa<�a<Z�a<��a<ܪa<�a<i�a<��a<ޫa<�a<=�a<m�a<��a<ܬa<��a<%�a<B�a<_�a<��a<��a<�a<�a<�a<*�a<G�a<_�a<�a<|�a<z�a<��a<��a<��a<Įa<ʮa<Ѯa<خa<�a<�a<�a<ɮa<Ϯa<Ԯa<��a<Юa<��a<��a<��a<s�a<��a<j�a<K�a<2�a<�a<��a<�a<̭a<��a<��a<L�a<5�a<)�a<�a<ͬa<��a<p�a<=�a<!�a<�a<��a<q�a<;�a<�a<Ϫa<��a<m�a<#�a<�a<��a<i�a<.�a<�a<��a<>�a< �a<��a<g�a<�a<ɦa<e�a<�a<Υa<s�a<�a<��a<M�a<�a<��a<3�a<Ģa<k�a<�a<��a<B�a<֠a<f�a<��a<��a<%�a<Þa<W�a<�a<_�a<	�a<��a<3�a<ћa<a�a<�a<��a<)�a<��a<Z�a<�a<s�a<�a<��a<M�a<�a<��a< �a<��a<v�a<#�a<Ôa<i�a<
�a<��a<q�a<%�a<ƒa<��a</�a<�a<��a<p�a<=�a<�a<��a<��a<Y�a<+�a<	�a<ɏa<��a<��a<V�a<I�a<'�a<�a<��a<�a<ގa<؎a<ӎa<��a<��a<��a<��a<׎a<��a<ގa<�a<�a<�a<3�a<�  �  G�a<W�a<��a<��a<Ϗa<�a<�a<m�a<{�a<ېa<�a<,�a<��a<��a<��a<3�a<��a<��a<#�a<��a<��a<1�a<_�a<ݔa<�a<��a<�a<B�a<��a<��a<~�a<ٗa<^�a<��a<�a<��a<�a<��a<ޚa<O�a<��a<!�a<��a<�a<��a<��a<��a<�a<]�a<۟a<F�a<Ҡa<�a<��a<�a<n�a<�a<H�a<̣a<�a<��a<��a<_�a<åa<�a<��a<Цa<K�a<��a<�a</�a<��a<�a<0�a<��a<��a<�a<X�a<��a<��a<�a<e�a<��a<̫a<�a<@�a<{�a<��a<�a<�a<7�a<G�a<��a<��a<��a<��a<�a<�a<$�a<P�a<[�a<[�a<��a<��a<��a<��a<Ǯa<ɮa<Ʈa<�a<̮a<�a<��a<ޮa<Юa<ڮa<׮a<��a<Ȯa<��a<��a<��a<~�a<w�a<D�a<M�a<(�a<'�a<��a<�a<ԭa<��a<��a<T�a<Z�a<
�a<�a<ݬa<��a<z�a<:�a<4�a<Ыa<��a<��a<?�a<)�a<Ǫa<��a<Y�a<,�a<�a<��a<c�a<	�a<ߨa<��a<[�a<��a<��a<h�a<�a<Ӧa<h�a<�a<��a<P�a<�a<��a<i�a<�a<��a<2�a<΢a<u�a<�a<��a<�a<ݠa<d�a<��a<��a<!�a<Ϟa<6�a<��a<��a<�a<��a<.�a<՛a<P�a<�a<z�a<�a<��a<6�a<�a<u�a<*�a<��a<O�a<�a<{�a<=�a<��a<q�a<��a<��a<]�a<�a<Óa<Y�a<)�a<��a<��a<4�a<�a<��a<W�a<Q�a<�a<ɐa<��a<c�a<'�a<�a<�a<��a<��a<Q�a<P�a<,�a<	�a<�a<ݎa<ߎa<��a<Ǝa<��a<��a<Îa<��a<ώa<��a<ێa<�a<�a<�a<�a<�  �  E�a<c�a<|�a<��a<ďa<��a<6�a<D�a<��a<Őa<�a<@�a<f�a<��a<�a<:�a<w�a<ܒa<�a<y�a<Ɠa<�a<��a<ؔa<�a<��a<�a<K�a<��a<�a<x�a<�a<;�a<��a</�a<��a<�a<c�a<ךa<V�a<ϛa<3�a<��a<�a<��a<��a<v�a<��a<`�a<ßa<I�a<��a<%�a<��a<��a<�a<�a<I�a<��a<(�a<��a<��a<M�a<��a<)�a<��a<զa<5�a<��a<�a<>�a<��a<�a<-�a<q�a<۩a<�a<b�a<��a<Ѫa< �a<d�a<��a<Ыa<�a<=�a<p�a<��a<۬a<�a<�a<G�a<{�a<��a<��a<˭a<�a<!�a<0�a<9�a<b�a<j�a<��a<��a<��a<��a<îa<��a<Ѯa<ˮa<خa<�a<ڮa<�a<ۮa<Įa<ʮa<ٮa<��a<Ʈa<��a<��a<��a<v�a<`�a<K�a<4�a<�a<�a<حa<̭a<��a<s�a<f�a<D�a<�a<��a<��a<��a<��a<A�a<�a<�a<��a<��a<K�a<�a<�a<��a<W�a<&�a<�a<��a<c�a<&�a<بa<��a<7�a<��a<��a<Y�a<"�a<��a<a�a<�a<ɥa<b�a<�a<��a<N�a<�a<��a<<�a<Тa<\�a<�a<��a<7�a<Ϡa<^�a<�a<��a<#�a<��a<U�a<�a<��a<�a<��a<?�a<̛a<U�a<�a<��a<�a<��a<S�a<�a<r�a<�a<��a<D�a<�a<��a<�a<ƕa<p�a<�a<��a<c�a<
�a<��a<\�a<%�a<ؒa<x�a<4�a<��a<��a<w�a<&�a<��a<ΐa<��a<K�a<.�a<�a<֏a<��a<s�a<o�a<K�a<!�a<�a<�a<�a<ߎa<ˎa<Ɏa<��a<��a<��a<Ўa<��a<�a<֎a<Ԏa<��a<�a<)�a<�  �  ,�a<u�a<p�a<��a<Տa<�a<<�a<A�a<��a<��a<�a<?�a<m�a<ʑa<֑a<Y�a<{�a<�a<�a<h�a<ٓa<�a<��a<��a<6�a<��a<ޕa<Y�a<��a<#�a<b�a<��a<L�a<��a<(�a<r�a<�a<`�a<��a<C�a<ƛa<@�a<��a<+�a<��a<�a<p�a<�a<g�a<̟a<Q�a<��a<>�a<��a<�a<q�a<Ӣa<i�a<��a<>�a<y�a<��a<[�a<��a<*�a<t�a<�a<,�a<��a<�a<E�a<��a<Ѩa<N�a<s�a<�a<��a<Z�a<��a<ܪa<7�a<G�a<��a<ɫa<�a<?�a<l�a<��a<��a<�a<�a<Z�a<s�a<��a<ҭa<˭a<�a<�a<9�a<H�a<a�a<��a<n�a<��a<��a<Ůa<��a<Ǯa<ڮa<��a<�a<ʮa<�a<ʮa<Ӯa<�a<��a<ݮa<��a<Ůa<��a<��a<��a<_�a<r�a<2�a<F�a<�a<�a<�a<��a<��a<p�a<x�a<-�a<%�a<��a<ìa<��a<Q�a<`�a<	�a<��a<��a<u�a<^�a<�a<�a<��a<r�a<'�a<ߩa<��a<S�a<1�a<èa<��a<I�a<�a<��a<A�a<-�a<��a<��a<�a<��a<n�a<�a<��a<D�a<��a<��a<6�a<עa<e�a<�a<��a<P�a<Ƞa<y�a<��a<��a<B�a<��a<k�a<ҝa<��a<�a<��a<A�a<��a<h�a<�a<��a<�a<��a<Q�a<͘a<��a<�a<ȗa<3�a<�a<��a< �a<ޕa<T�a<�a<��a<l�a<�a<��a<u�a<
�a<ܒa<z�a<G�a<��a<��a<��a<&�a<�a<��a<��a<Z�a<-�a<�a<��a<��a<s�a<w�a<7�a<+�a<�a<�a<��a<Ȏa<��a<��a<��a<̎a<��a<Ԏa<��a<�a<̎a<�a<��a<��a<;�a<�  �  0�a<p�a<��a<��a<ҏa<�a<*�a<X�a<��a<Đa<�a<#�a<r�a<ˑa<�a<U�a<��a<ɒa<'�a<|�a<ēa<#�a<u�a<Ŕa<)�a<��a<�a<Q�a<��a<�a<{�a<ٗa<L�a<��a<&�a<��a<��a<c�a<�a<L�a<˛a<-�a<��a<(�a<��a<��a<v�a<�a<b�a<Пa<N�a<��a<%�a<��a<�a<z�a<�a<^�a<��a< �a<��a<��a<X�a<��a<�a<|�a<Ԧa<>�a<��a<�a<4�a<��a<ߨa<7�a<y�a<ũa<�a<c�a<��a<ߪa<�a<^�a<��a<ëa<�a<H�a<n�a<��a<ʬa<��a<-�a<J�a<�a<��a<��a<ѭa<�a<�a<?�a<F�a<K�a<v�a<��a<��a<��a<��a<��a<Ǯa<��a<ܮa<�a<ɮa<ۮa<߮a<Ϯa<ۮa<��a<��a<ɮa<��a<��a<��a<y�a<v�a<_�a<6�a<A�a<�a<�a<�a<��a<��a<��a<g�a<C�a<!�a<�a<ɬa<��a<i�a<\�a<�a<۫a<��a<��a<I�a<�a<ݪa<��a<e�a<!�a<�a<��a<R�a<$�a<ܨa<��a<I�a<�a<��a<k�a<�a<��a<l�a<�a<ťa<[�a<�a<��a<]�a<�a<��a<2�a<Ңa<i�a<�a<��a<7�a<��a<r�a<�a<��a<7�a<��a<M�a<�a<��a<�a<��a<6�a<ƛa<T�a<��a<��a<�a<��a<N�a<ۘa<|�a<
�a<��a<S�a<�a<z�a<$�a<Õa<k�a<�a<��a<c�a<�a<��a<c�a<�a<ϒa<��a<7�a<�a<��a<j�a<,�a<�a<��a<��a<Y�a<�a< �a<Џa<��a<��a<f�a<@�a<*�a<�a<�a<��a<ǎa<̎a<ǎa<��a<��a<��a<��a<Ўa<Ɏa<Ȏa<�a<�a<�a<(�a<�  �  Y�a<J�a<��a<��a<ʏa<�a<�a<[�a<r�a<ǐa<��a<E�a<u�a<��a<�a<�a<��a<ڒa<�a<v�a<��a<#�a<h�a<�a<!�a<��a<�a<9�a<��a<�a<��a<ȗa<M�a<��a<�a<��a<��a<��a<��a<^�a<՛a<2�a<��a<�a<��a<��a<��a<�a<]�a<ȟa<0�a<��a<!�a<��a<��a<v�a<�a<<�a<ԣa<!�a<��a<�a<L�a<��a<�a<��a<Ϧa<F�a<��a<��a<B�a<��a<��a<�a<��a<éa<�a<R�a<��a<�a<�a<z�a<��a<߫a<�a<B�a<x�a<��a<�a<�a<,�a<7�a<n�a<��a<��a<�a<حa<�a<�a<B�a<o�a<i�a<��a<�a<��a<��a<Ʈa<Ǯa<Įa<�a<®a<�a<̮a<�a<Үa<��a<�a<��a<��a<��a<��a<��a<v�a<��a<N�a<`�a<�a<)�a<��a<ޭa<ӭa<��a<��a<K�a<E�a<�a<�a<ˬa<��a<��a<%�a<&�a<�a<��a<��a<1�a<�a<Ъa<��a<\�a<+�a<�a<��a<t�a<�a<�a<x�a<I�a<�a<��a<e�a<�a<ئa<K�a<!�a<ϥa<`�a<�a<��a<b�a<�a<��a<0�a<͢a<b�a<�a<��a<3�a<�a<\�a<��a<��a<�a<מa<O�a<�a<f�a< �a<��a<+�a<ڛa<O�a< �a<|�a<%�a<��a<T�a<�a<Z�a<%�a<��a<I�a<ݖa<��a</�a<��a<��a<�a<Ĕa<[�a<�a<��a<\�a<0�a<��a<��a<$�a<�a<��a<t�a<H�a<ڐa<ːa<z�a<U�a<;�a<�a<؏a<��a<��a<[�a<N�a<*�a<�a<�a<Ҏa<�a<��a<؎a<��a<��a<Ԏa<��a<Ǝa<��a<�a<َa<�a<(�a<�a<�  �  S�a<O�a<��a<��a<ʏa<��a<'�a<Z�a<��a<ϐa<�a<1�a<{�a<��a<�a<7�a<��a<ђa<�a<��a<ӓa<$�a<s�a<˔a<&�a<��a<�a<<�a<��a<��a<r�a<�a<P�a<��a<�a<��a<��a<v�a<ݚa<S�a<��a<+�a<��a<�a<��a<�a<t�a<�a<i�a<ޟa<W�a<��a<!�a<��a<�a<v�a<�a<O�a<£a< �a<��a<�a<g�a<ɥa<�a<|�a<�a<C�a<��a<�a<8�a<z�a<�a<6�a<��a<ǩa<�a<X�a<��a<�a<+�a<[�a<}�a<֫a<��a<B�a<r�a<��a<ͬa<��a<1�a<\�a<��a<��a<��a<�a<�a<�a<+�a<M�a<T�a<a�a<��a<��a<��a<��a<��a<��a<Ӯa<ݮa<ɮa<�a<Ȯa<̮a<�a<ͮa<Ԯa<��a<��a<��a<��a<��a<��a<f�a<G�a<Y�a< �a<!�a< �a<ޭa<ƭa<��a<��a<p�a<N�a<
�a<�a<Ҭa<��a<��a<>�a<!�a<�a<��a<��a<X�a<�a<۪a<��a<b�a<&�a<�a<��a<p�a<�a<Өa<��a<L�a<��a<��a<[�a<�a<Ŧa<g�a<�a<��a<Z�a<�a<��a<^�a<��a<��a<0�a<٢a<w�a<�a<��a<2�a<Ϡa<h�a<��a<��a<)�a<Şa<M�a<�a<��a<�a<��a<1�a<ƛa<b�a<��a<��a<�a<��a</�a<��a<z�a<�a<��a<F�a<�a<��a<+�a<ҕa<h�a<��a<��a<U�a<�a<��a<f�a<�a<ʒa<��a<I�a<�a<��a<o�a<@�a<��a<̐a<��a<_�a< �a<�a<�a<��a<��a<f�a<F�a<%�a<�a<�a<َa<�a<��a<��a<Ŏa<��a<��a<��a<��a<Îa<ێa<�a<�a<�a<�a<�  �  <�a<m�a<|�a<��a<ݏa<��a<)�a<G�a<��a<��a<	�a<'�a<w�a<Ña<��a<R�a<��a<Βa<,�a<g�a<��a<	�a<|�a<ɔa<<�a<k�a<�a<N�a<��a<3�a<v�a<�a<<�a<��a<,�a<��a<�a<[�a<�a<T�a<Λa<X�a<��a</�a<z�a<�a<y�a<�a<W�a<ğa<=�a<��a<<�a<��a<�a<y�a<�a<a�a<��a<5�a<��a<�a<N�a<��a<'�a<~�a<�a< �a<��a<�a<X�a<��a<�a<:�a<m�a<֩a<�a<b�a<��a<Ϊa<#�a<\�a<��a<ݫa<�a<I�a<X�a<��a<̬a<�a<�a<H�a<g�a<��a<��a<έa<
�a<�a<:�a<L�a<J�a<��a<t�a<��a<��a<��a<��a<ήa<��a<Ǯa<�a<Ϯa< �a<خa<׮a<Ϯa<��a<Ϯa<��a<��a<��a<��a<��a<o�a<��a<B�a<>�a<�a<�a<�a<��a<��a<v�a<a�a</�a<*�a<�a<ͬa<��a<q�a<Y�a<�a<�a<��a<u�a<F�a<�a<�a<��a<x�a<�a<�a<��a<i�a<@�a<רa<��a<9�a<��a<��a<`�a<�a<��a<o�a<�a<ȥa<��a< �a<��a<;�a<��a<��a<:�a<Ȣa<^�a<��a<��a<N�a<��a<v�a<�a<��a<:�a<��a<b�a<ܝa<q�a<�a<��a<>�a<ɛa<f�a<ٚa<��a<�a<ʙa<Y�a<�a<~�a<��a<��a<K�a<�a<��a<�a<ɕa<i�a<,�a<��a<^�a<�a<��a<{�a<�a<֒a<s�a<5�a<�a<��a<t�a<)�a<�a<��a<��a<_�a<�a<�a<��a<��a<s�a<_�a<C�a<1�a<�a<�a<��a<͎a<�a<��a<��a<��a<��a<Ǝa<Ŏa<׎a<͎a<ߎa<��a<�a<K�a<�  �  /�a<`�a<��a<��a<ԏa<��a<$�a<`�a<��a<��a<�a</�a<s�a<��a<��a<8�a<��a<͒a<2�a<s�a<ړa<�a<q�a<ǔa<2�a<��a<�a<B�a<��a<�a<s�a<ڗa<W�a<��a<�a<��a< �a<��a<ޚa<R�a<��a<1�a<��a<$�a<��a<�a<x�a<�a<c�a<�a<P�a<��a<1�a<��a<�a<y�a<�a<I�a<��a<,�a<��a<��a<r�a<ĥa<�a<{�a<�a<4�a<��a<ܧa<8�a<{�a<�a</�a<��a<ϩa<�a<S�a<��a<�a<�a<Z�a<��a<ȫa<��a<H�a<l�a<��a<ɬa<��a<-�a<g�a<x�a<��a<��a<ۭa<�a<�a<+�a<C�a<X�a<��a<��a<��a<��a<��a<��a<ɮa<ͮa<׮a<ٮa<Ʈa<׮a<®a<ծa<Ӯa<ޮa<��a<��a<��a<��a<��a<~�a<b�a<S�a<6�a<1�a<�a<��a<�a<��a<��a<��a<u�a<=�a<,�a<�a<ʬa<��a<v�a<?�a<�a<߫a<īa<��a<_�a<�a<٪a<��a<n�a<#�a<�a<��a<S�a<�a<Өa<��a<T�a<�a<��a<P�a<�a<Ѧa<g�a<�a<��a<`�a<��a<��a<P�a<��a<��a<1�a<Ӣa<��a<�a<��a<C�a<Πa<c�a<�a<��a<#�a<��a<Z�a<�a<��a<&�a<��a<4�a<ƛa<d�a<�a<��a<�a<��a<0�a<�a<s�a<%�a<��a<:�a<ޖa<��a<7�a<��a<g�a<��a<��a<S�a<�a<��a<q�a<�a<Ȓa<��a<T�a<��a<��a<q�a<6�a<�a<Ða<��a<U�a<$�a<�a<Ώa<��a<��a<a�a<=�a<,�a<�a<��a<�a<Ďa<Ȏa<��a<��a<��a<ˎa<��a<��a<Ǝa<�a<�a<�a<��a<�a<�  �  f�a<X�a<��a<��a<ʏa<�a<"�a<G�a<|�a<��a<�a<6�a<��a<��a<
�a<)�a<��a<̒a< �a<d�a<��a<�a<q�a<ڔa<#�a<��a<�a<J�a<Җa<�a<��a<�a<A�a<��a<,�a<��a<�a<p�a<Ěa<n�a<��a<I�a<��a<�a<��a<�a<u�a<�a<V�a<ßa<2�a<��a<�a<��a<��a<u�a<�a<@�a<֣a<�a<��a<ޤa<G�a<��a<�a<�a<ݦa<A�a<��a<��a<]�a<��a<�a<�a<��a<��a<(�a<i�a<��a<ݪa<�a<}�a<��a<��a<�a<6�a<u�a<��a<۬a<��a<�a<>�a<`�a<��a<��a<��a<�a<�a<#�a<O�a<c�a<_�a<z�a<��a<��a<��a<Įa<��a<Ѯa<֮a<ʮa<��a<߮a<ܮa<�a<��a<Ȯa<��a<ˮa<��a<��a<��a<��a<��a<V�a<l�a<(�a<�a<�a<ޭa<Эa<��a<v�a<U�a<4�a<�a<��a<ܬa<��a<��a<0�a<5�a<߫a<��a<q�a<>�a<	�a<٪a<��a<_�a<+�a<�a<��a<��a<�a<��a<��a<=�a<�a<��a<u�a<��a<��a<N�a<1�a<��a<x�a<!�a<��a<Z�a<��a<��a<2�a<Ǣa<\�a<��a<��a<-�a<�a<_�a<��a<��a<�a<ٞa<I�a<�a<d�a<��a<��a<1�a<ʛa<^�a<��a<|�a<-�a<ϙa<=�a<��a<b�a<�a<��a<\�a<��a<h�a<"�a<��a<��a<�a<�a<c�a<�a<��a<e�a<$�a<ɒa<z�a<+�a<�a<��a<l�a<T�a<�a<̐a<��a<b�a</�a<�a<Ǐa<��a<u�a<a�a<M�a<$�a<�a<��a<ڎa<��a<Ўa<Ďa<֎a<��a<��a<��a<Ҏa<��a<Ύa<ӎa<�a<�a<�a<�  �  /�a<`�a<��a<��a<ԏa<��a<$�a<`�a<��a<��a<�a</�a<s�a<��a<��a<8�a<��a<͒a<2�a<s�a<ړa<�a<q�a<ǔa<2�a<��a<�a<B�a<��a<�a<s�a<ڗa<W�a<��a<�a<��a< �a<��a<ޚa<R�a<��a<1�a<��a<$�a<��a<�a<x�a<�a<c�a<�a<P�a<��a<1�a<��a<�a<y�a<�a<I�a<��a<,�a<��a<��a<r�a<ĥa<�a<{�a<�a<4�a<��a<ܧa<8�a<{�a<�a</�a<��a<ϩa<�a<S�a<��a<�a<�a<Z�a<��a<ȫa<��a<H�a<l�a<��a<ɬa<��a<-�a<g�a<x�a<��a<��a<ۭa<�a<�a<+�a<C�a<X�a<��a<��a<��a<��a<��a<��a<ɮa<ͮa<׮a<ٮa<Ʈa<׮a<®a<ծa<Ӯa<ޮa<��a<��a<��a<��a<��a<~�a<b�a<S�a<6�a<1�a<�a<��a<�a<��a<��a<��a<u�a<=�a<,�a<�a<ʬa<��a<v�a<?�a<�a<߫a<īa<��a<_�a<�a<٪a<��a<n�a<#�a<�a<��a<S�a<�a<Өa<��a<T�a<�a<��a<P�a<�a<Ѧa<g�a<�a<��a<`�a<��a<��a<P�a<��a<��a<1�a<Ӣa<��a<�a<��a<C�a<Πa<c�a<�a<��a<#�a<��a<Z�a<�a<��a<&�a<��a<4�a<ƛa<d�a<�a<��a<�a<��a<0�a<�a<s�a<%�a<��a<:�a<ޖa<��a<7�a<��a<g�a<��a<��a<S�a<�a<��a<q�a<�a<Ȓa<��a<T�a<��a<��a<q�a<6�a<�a<Ða<��a<U�a<$�a<�a<Ώa<��a<��a<a�a<=�a<,�a<�a<��a<�a<Ďa<Ȏa<��a<��a<��a<ˎa<��a<��a<Ǝa<�a<�a<�a<��a<�a<�  �  <�a<m�a<|�a<��a<ݏa<��a<)�a<G�a<��a<��a<	�a<'�a<w�a<Ña<��a<R�a<��a<Βa<,�a<g�a<��a<	�a<|�a<ɔa<<�a<k�a<�a<N�a<��a<3�a<v�a<�a<<�a<��a<,�a<��a<�a<[�a<�a<T�a<Λa<X�a<��a</�a<z�a<�a<y�a<�a<W�a<ğa<=�a<��a<<�a<��a<�a<y�a<�a<a�a<��a<5�a<��a<�a<N�a<��a<'�a<~�a<�a< �a<��a<�a<X�a<��a<�a<:�a<m�a<֩a<�a<b�a<��a<Ϊa<#�a<\�a<��a<ݫa<�a<I�a<X�a<��a<̬a<�a<�a<H�a<g�a<��a<��a<έa<
�a<�a<:�a<L�a<J�a<��a<t�a<��a<��a<��a<��a<ήa<��a<Ǯa<�a<Ϯa< �a<خa<׮a<Ϯa<��a<Ϯa<��a<��a<��a<��a<��a<o�a<��a<B�a<>�a<�a<�a<�a<��a<��a<v�a<a�a</�a<*�a<�a<ͬa<��a<q�a<Y�a<�a<�a<��a<u�a<F�a<�a<�a<��a<x�a<�a<�a<��a<i�a<@�a<רa<��a<9�a<��a<��a<`�a<�a<��a<o�a<�a<ȥa<��a< �a<��a<;�a<��a<��a<:�a<Ȣa<^�a<��a<��a<N�a<��a<v�a<�a<��a<:�a<��a<b�a<ܝa<q�a<�a<��a<>�a<ɛa<f�a<ٚa<��a<�a<ʙa<Y�a<�a<~�a<��a<��a<K�a<�a<��a<�a<ɕa<i�a<,�a<��a<^�a<�a<��a<{�a<�a<֒a<s�a<5�a<�a<��a<t�a<)�a<�a<��a<��a<_�a<�a<�a<��a<��a<s�a<_�a<C�a<1�a<�a<�a<��a<͎a<�a<��a<��a<��a<��a<Ǝa<Ŏa<׎a<͎a<ߎa<��a<�a<K�a<�  �  S�a<O�a<��a<��a<ʏa<��a<'�a<Z�a<��a<ϐa<�a<1�a<{�a<��a<�a<7�a<��a<ђa<�a<��a<ӓa<$�a<s�a<˔a<&�a<��a<�a<<�a<��a<��a<r�a<�a<P�a<��a<�a<��a<��a<v�a<ݚa<S�a<��a<+�a<��a<�a<��a<�a<t�a<�a<i�a<ޟa<W�a<��a<!�a<��a<�a<v�a<�a<O�a<£a< �a<��a<�a<g�a<ɥa<�a<|�a<�a<C�a<��a<�a<8�a<z�a<�a<6�a<��a<ǩa<�a<X�a<��a<�a<+�a<[�a<}�a<֫a<��a<B�a<r�a<��a<ͬa<��a<1�a<\�a<��a<��a<��a<�a<�a<�a<+�a<M�a<T�a<a�a<��a<��a<��a<��a<��a<��a<Ӯa<ݮa<ɮa<�a<Ȯa<̮a<�a<ͮa<Ԯa<��a<��a<��a<��a<��a<��a<f�a<G�a<Y�a< �a<!�a< �a<ޭa<ƭa<��a<��a<p�a<N�a<
�a<�a<Ҭa<��a<��a<>�a<!�a<�a<��a<��a<X�a<�a<۪a<��a<b�a<&�a<�a<��a<p�a<�a<Өa<��a<L�a<��a<��a<[�a<�a<Ŧa<g�a<�a<��a<Z�a<�a<��a<^�a<��a<��a<0�a<٢a<w�a<�a<��a<2�a<Ϡa<h�a<��a<��a<)�a<Şa<M�a<�a<��a<�a<��a<1�a<ƛa<b�a<��a<��a<�a<��a</�a<��a<z�a<�a<��a<F�a<�a<��a<+�a<ҕa<h�a<��a<��a<U�a<�a<��a<f�a<�a<ʒa<��a<I�a<�a<��a<o�a<@�a<��a<̐a<��a<_�a< �a<�a<�a<��a<��a<f�a<F�a<%�a<�a<�a<َa<�a<��a<��a<Ŏa<��a<��a<��a<��a<Îa<ێa<�a<�a<�a<�a<�  �  Y�a<J�a<��a<��a<ʏa<�a<�a<[�a<r�a<ǐa<��a<E�a<u�a<��a<�a<�a<��a<ڒa<�a<v�a<��a<#�a<h�a<�a<!�a<��a<�a<9�a<��a<�a<��a<ȗa<M�a<��a<�a<��a<��a<��a<��a<^�a<՛a<2�a<��a<�a<��a<��a<��a<�a<]�a<ȟa<0�a<��a<!�a<��a<��a<v�a<�a<<�a<ԣa<!�a<��a<�a<L�a<��a<�a<��a<Ϧa<F�a<��a<��a<B�a<��a<��a<�a<��a<éa<�a<R�a<��a<�a<�a<z�a<��a<߫a<�a<B�a<x�a<��a<�a<�a<,�a<7�a<n�a<��a<��a<�a<حa<�a<�a<B�a<o�a<i�a<��a<�a<��a<��a<Ʈa<Ǯa<Įa<�a<®a<�a<̮a<�a<Үa<��a<�a<��a<��a<��a<��a<��a<v�a<��a<N�a<`�a<�a<)�a<��a<ޭa<ӭa<��a<��a<K�a<E�a<�a<�a<ˬa<��a<��a<%�a<&�a<�a<��a<��a<1�a<�a<Ъa<��a<\�a<+�a<�a<��a<t�a<�a<�a<x�a<I�a<�a<��a<e�a<�a<ئa<K�a<!�a<ϥa<`�a<�a<��a<b�a<�a<��a<0�a<͢a<b�a<�a<��a<3�a<�a<\�a<��a<��a<�a<מa<O�a<�a<f�a< �a<��a<+�a<ڛa<O�a< �a<|�a<%�a<��a<T�a<�a<Z�a<%�a<��a<I�a<ݖa<��a</�a<��a<��a<�a<Ĕa<[�a<�a<��a<\�a<0�a<��a<��a<$�a<�a<��a<t�a<H�a<ڐa<ːa<z�a<U�a<;�a<�a<؏a<��a<��a<[�a<N�a<*�a<�a<�a<Ҏa<�a<��a<؎a<��a<��a<Ԏa<��a<Ǝa<��a<�a<َa<�a<(�a<�a<�  �  0�a<p�a<��a<��a<ҏa<�a<*�a<X�a<��a<Đa<�a<#�a<r�a<ˑa<�a<U�a<��a<ɒa<'�a<|�a<ēa<#�a<u�a<Ŕa<)�a<��a<�a<Q�a<��a<�a<{�a<ٗa<L�a<��a<&�a<��a<��a<c�a<�a<L�a<˛a<-�a<��a<(�a<��a<��a<v�a<�a<b�a<Пa<N�a<��a<%�a<��a<�a<z�a<�a<^�a<��a< �a<��a<��a<X�a<��a<�a<|�a<Ԧa<>�a<��a<�a<4�a<��a<ߨa<7�a<y�a<ũa<�a<c�a<��a<ߪa<�a<^�a<��a<ëa<�a<H�a<n�a<��a<ʬa<��a<-�a<J�a<�a<��a<��a<ѭa<�a<�a<?�a<F�a<K�a<v�a<��a<��a<��a<��a<��a<Ǯa<��a<ܮa<�a<ɮa<ۮa<߮a<Ϯa<ۮa<��a<��a<ɮa<��a<��a<��a<y�a<v�a<_�a<6�a<A�a<�a<�a<�a<��a<��a<��a<g�a<C�a<!�a<�a<ɬa<��a<i�a<\�a<�a<۫a<��a<��a<I�a<�a<ݪa<��a<e�a<!�a<�a<��a<R�a<$�a<ܨa<��a<I�a<�a<��a<k�a<�a<��a<l�a<�a<ťa<[�a<�a<��a<]�a<�a<��a<2�a<Ңa<i�a<�a<��a<7�a<��a<r�a<�a<��a<7�a<��a<M�a<�a<��a<�a<��a<6�a<ƛa<T�a<��a<��a<�a<��a<N�a<ۘa<|�a<
�a<��a<S�a<�a<z�a<$�a<Õa<k�a<�a<��a<c�a<�a<��a<c�a<�a<ϒa<��a<7�a<�a<��a<j�a<,�a<�a<��a<��a<Y�a<�a< �a<Џa<��a<��a<f�a<@�a<*�a<�a<�a<��a<ǎa<̎a<ǎa<��a<��a<��a<��a<Ўa<Ɏa<Ȏa<�a<�a<�a<(�a<�  �  ,�a<u�a<p�a<��a<Տa<�a<<�a<A�a<��a<��a<�a<?�a<m�a<ʑa<֑a<Y�a<{�a<�a<�a<h�a<ٓa<�a<��a<��a<6�a<��a<ޕa<Y�a<��a<#�a<b�a<��a<L�a<��a<(�a<r�a<�a<`�a<��a<C�a<ƛa<@�a<��a<+�a<��a<�a<p�a<�a<g�a<̟a<Q�a<��a<>�a<��a<�a<q�a<Ӣa<i�a<��a<>�a<y�a<��a<[�a<��a<*�a<t�a<�a<,�a<��a<�a<E�a<��a<Ѩa<N�a<s�a<�a<��a<Z�a<��a<ܪa<7�a<G�a<��a<ɫa<�a<?�a<l�a<��a<��a<�a<�a<Z�a<s�a<��a<ҭa<˭a<�a<�a<9�a<H�a<a�a<��a<n�a<��a<��a<Ůa<��a<Ǯa<ڮa<��a<�a<ʮa<�a<ʮa<Ӯa<�a<��a<ݮa<��a<Ůa<��a<��a<��a<_�a<r�a<2�a<F�a<�a<�a<�a<��a<��a<p�a<x�a<-�a<%�a<��a<ìa<��a<Q�a<`�a<	�a<��a<��a<u�a<^�a<�a<�a<��a<r�a<'�a<ߩa<��a<S�a<1�a<èa<��a<I�a<�a<��a<A�a<-�a<��a<��a<�a<��a<n�a<�a<��a<D�a<��a<��a<6�a<עa<e�a<�a<��a<P�a<Ƞa<y�a<��a<��a<B�a<��a<k�a<ҝa<��a<�a<��a<A�a<��a<h�a<�a<��a<�a<��a<Q�a<͘a<��a<�a<ȗa<3�a<�a<��a< �a<ޕa<T�a<�a<��a<l�a<�a<��a<u�a<
�a<ܒa<z�a<G�a<��a<��a<��a<&�a<�a<��a<��a<Z�a<-�a<�a<��a<��a<s�a<w�a<7�a<+�a<�a<�a<��a<Ȏa<��a<��a<��a<̎a<��a<Ԏa<��a<�a<̎a<�a<��a<��a<;�a<�  �  E�a<c�a<|�a<��a<ďa<��a<6�a<D�a<��a<Őa<�a<@�a<f�a<��a<�a<:�a<w�a<ܒa<�a<y�a<Ɠa<�a<��a<ؔa<�a<��a<�a<K�a<��a<�a<x�a<�a<;�a<��a</�a<��a<�a<c�a<ךa<V�a<ϛa<3�a<��a<�a<��a<��a<v�a<��a<`�a<ßa<I�a<��a<%�a<��a<��a<�a<�a<I�a<��a<(�a<��a<��a<M�a<��a<)�a<��a<զa<5�a<��a<�a<>�a<��a<�a<-�a<q�a<۩a<�a<b�a<��a<Ѫa< �a<d�a<��a<Ыa<�a<=�a<p�a<��a<۬a<�a<�a<G�a<{�a<��a<��a<˭a<�a<!�a<0�a<9�a<b�a<j�a<��a<��a<��a<��a<îa<��a<Ѯa<ˮa<خa<�a<ڮa<�a<ۮa<Įa<ʮa<ٮa<��a<Ʈa<��a<��a<��a<v�a<`�a<K�a<4�a<�a<�a<حa<̭a<��a<s�a<f�a<D�a<�a<��a<��a<��a<��a<A�a<�a<�a<��a<��a<K�a<�a<�a<��a<W�a<&�a<�a<��a<c�a<&�a<بa<��a<7�a<��a<��a<Y�a<"�a<��a<a�a<�a<ɥa<b�a<�a<��a<N�a<�a<��a<<�a<Тa<\�a<�a<��a<7�a<Ϡa<^�a<�a<��a<#�a<��a<U�a<�a<��a<�a<��a<?�a<̛a<U�a<�a<��a<�a<��a<S�a<�a<r�a<�a<��a<D�a<�a<��a<�a<ƕa<p�a<�a<��a<c�a<
�a<��a<\�a<%�a<ؒa<x�a<4�a<��a<��a<w�a<&�a<��a<ΐa<��a<K�a<.�a<�a<֏a<��a<s�a<o�a<K�a<!�a<�a<�a<�a<ߎa<ˎa<Ɏa<��a<��a<��a<Ўa<��a<�a<֎a<Ԏa<��a<�a<)�a<�  �  G�a<W�a<��a<��a<Ϗa<�a<�a<m�a<{�a<ېa<�a<,�a<��a<��a<��a<3�a<��a<��a<#�a<��a<��a<1�a<_�a<ݔa<�a<��a<�a<B�a<��a<��a<~�a<ٗa<^�a<��a<�a<��a<�a<��a<ޚa<O�a<��a<!�a<��a<�a<��a<��a<��a<�a<]�a<۟a<F�a<Ҡa<�a<��a<�a<n�a<�a<H�a<̣a<�a<��a<��a<_�a<åa<�a<��a<Цa<K�a<��a<�a</�a<��a<�a<0�a<��a<��a<�a<X�a<��a<��a<�a<e�a<��a<̫a<�a<@�a<{�a<��a<�a<�a<7�a<G�a<��a<��a<��a<��a<�a<�a<$�a<P�a<[�a<[�a<��a<��a<��a<��a<Ǯa<ɮa<Ʈa<�a<̮a<�a<��a<ޮa<Юa<ڮa<׮a<��a<Ȯa<��a<��a<��a<~�a<w�a<D�a<M�a<(�a<'�a<��a<�a<ԭa<��a<��a<T�a<Z�a<
�a<�a<ݬa<��a<z�a<:�a<4�a<Ыa<��a<��a<?�a<)�a<Ǫa<��a<Y�a<,�a<�a<��a<c�a<	�a<ߨa<��a<[�a<��a<��a<h�a<�a<Ӧa<h�a<�a<��a<P�a<�a<��a<i�a<�a<��a<2�a<΢a<u�a<�a<��a<�a<ݠa<d�a<��a<��a<!�a<Ϟa<6�a<��a<��a<�a<��a<.�a<՛a<P�a<�a<z�a<�a<��a<6�a<�a<u�a<*�a<��a<O�a<�a<{�a<=�a<��a<q�a<��a<��a<]�a<�a<Óa<Y�a<)�a<��a<��a<4�a<�a<��a<W�a<Q�a<�a<ɐa<��a<c�a<'�a<�a<�a<��a<��a<Q�a<P�a<,�a<	�a<�a<ݎa<ߎa<��a<Ǝa<��a<��a<Îa<��a<ώa<��a<ێa<�a<�a<�a<�a<�  �  E�a<b�a<��a<��a<Ϗa< �a<�a<k�a<s�a<��a<�a<3�a<w�a<��a<��a<6�a<��a<Вa<*�a<d�a<��a<#�a<g�a<הa<1�a<��a<�a<L�a<��a<!�a<��a<җa<A�a<��a< �a<��a<��a<{�a<ۚa<P�a<ԛa<D�a<��a<�a<��a<�a<{�a<�a<T�a<џa<'�a<��a<0�a<��a<�a<t�a<�a<L�a<��a<)�a<��a<٤a<T�a<��a<�a<��a<�a<4�a<��a<��a<M�a<��a<�a<.�a<��a<ɩa<�a<Z�a<��a<ܪa<�a<i�a<��a<ޫa<�a<=�a<m�a<��a<ܬa<��a<%�a<B�a<_�a<��a<��a<�a<�a<�a<*�a<G�a<_�a<�a<|�a<z�a<��a<��a<��a<Įa<ʮa<Ѯa<خa<�a<�a<�a<ɮa<Ϯa<Ԯa<��a<Юa<��a<��a<��a<s�a<��a<j�a<K�a<2�a<�a<��a<�a<̭a<��a<��a<L�a<5�a<)�a<�a<ͬa<��a<p�a<=�a<!�a<�a<��a<q�a<;�a<�a<Ϫa<��a<m�a<#�a<�a<��a<i�a<.�a<�a<��a<>�a< �a<��a<g�a<�a<ɦa<e�a<�a<Υa<s�a<�a<��a<M�a<�a<��a<3�a<Ģa<k�a<�a<��a<B�a<֠a<f�a<��a<��a<%�a<Þa<W�a<�a<_�a<	�a<��a<3�a<ћa<a�a<�a<��a<)�a<��a<Z�a<�a<s�a<�a<��a<M�a<�a<��a< �a<��a<v�a<#�a<Ôa<i�a<
�a<��a<q�a<%�a<ƒa<��a</�a<�a<��a<p�a<=�a<�a<��a<��a<Y�a<+�a<	�a<ɏa<��a<��a<V�a<I�a<'�a<�a<��a<�a<ގa<؎a<ӎa<��a<��a<��a<��a<׎a<��a<ގa<�a<�a<�a<3�a<�  �  2�a<e�a<}�a<��a<��a<��a<2�a<T�a<��a<��a<��a<-�a<k�a<��a<��a<I�a<y�a<Ԓa<"�a<u�a<�a<�a<��a<��a<�a<��a<�a<C�a<��a<�a<h�a<��a<7�a<��a<+�a<��a<�a<`�a<�a<P�a<��a</�a<��a<%�a<��a<�a<^�a<��a<[�a<ߟa<\�a<��a<*�a<��a<�a<}�a<�a<Y�a<��a<*�a<��a<�a<n�a<��a<-�a<f�a<�a<7�a<��a<ߧa<6�a<��a<ܨa<@�a<q�a<ܩa<�a<_�a<��a<ͪa<6�a<N�a<��a<ūa<�a<D�a<t�a<��a<��a<�a<�a<s�a<{�a<��a<��a<ǭa<�a<�a<9�a<?�a<P�a<s�a<��a<��a<��a<��a<��a<��a<�a<Ϯa<�a<Ȯa<׮a<ͮa<�a<ɮa<Ǯa<ծa<��a<��a<��a<��a<��a<`�a<[�a<8�a<6�a<�a<�a<ʭa<ía<��a<��a<��a<=�a<�a<�a<��a<��a<x�a<Q�a<�a<�a<��a<��a<r�a<�a<�a<��a<[�a<.�a<�a<��a<T�a<�a<ɨa<��a<3�a<�a<��a<\�a<!�a<��a<n�a<�a<��a<^�a<��a<��a<N�a<�a<y�a<>�a<ˢa<y�a<�a<��a<<�a<��a<l�a<�a<��a<2�a<��a<W�a<�a<��a<#�a<��a<D�a<��a<i�a<�a<��a<�a<��a<>�a<טa<��a<�a<��a<H�a<�a<��a<�a<ݕa<[�a<�a<��a<Y�a<�a<��a<g�a<�a<�a<w�a<`�a<��a<��a<w�a<"�a<�a<Ða<��a<R�a<�a<��a<Џa<͏a<��a<l�a<G�a<�a<#�a<��a<��a<Ǝa<Ȏa<��a<Ȏa<��a<��a<̎a<��a<َa<׎a<؎a<�a<��a<$�a<�  �  I�a<^�a<y�a<��a<ˏa<�a<%�a<E�a<}�a<��a<��a<:�a<��a<��a<�a<<�a<��a<Ԓa<#�a<[�a<ēa<	�a<x�a<ϔa<+�a<��a<�a<H�a<��a<!�a<v�a<�a<G�a<��a<!�a<��a<��a<o�a<�a<Z�a<ța<P�a<��a<�a<��a<�a<r�a<�a<O�a<ɟa<.�a<��a< �a<��a<�a<k�a<բa<T�a<Σa<�a<��a<ܤa<R�a<��a<'�a<y�a<�a<3�a<��a<�a<Y�a<��a<�a<:�a<�a<ĩa<�a<\�a<��a<ުa<-�a<^�a<��a<�a<�a<>�a<r�a<��a<Ϭa<�a<�a<J�a<[�a<��a<��a<�a<��a<�a<*�a<R�a<g�a<j�a<}�a<��a<��a<��a<Ʈa<®a<ծa<̮a<֮a<ޮa<�a<خa<�a<ɮa<ήa<��a<��a<��a<��a<��a<��a<o�a<n�a<P�a</�a<�a<�a<�a<ͭa<��a<s�a<V�a<4�a<�a<��a<٬a<��a<c�a<C�a<+�a<�a<��a<h�a<H�a<�a<�a<��a<g�a<*�a<�a<��a<r�a</�a<֨a<��a<C�a<��a<��a<c�a<�a<��a<j�a<�a<¥a<�a<�a<��a<K�a<��a<��a<:�a<��a<c�a<�a<��a<2�a<�a<o�a<��a<��a<.�a<ўa<M�a<�a<b�a<�a<��a<=�a<ěa<d�a<�a<��a<"�a<˙a<P�a<�a<�a<�a<��a<O�a<�a<��a<#�a<ӕa<j�a<�a<˔a<c�a<�a<��a<n�a<�a<Ԓa<r�a<7�a<ܑa<��a<q�a<I�a<��a<��a<��a<e�a<3�a<�a<ʏa<��a<r�a<_�a<N�a<%�a<�a<�a<�a<܎a<ݎa<��a<̎a<��a<��a<��a<Ďa<a<׎a<ގa<�a<�a<6�a<�  �  ��a<��a<�a<�a<�a<[�a<_�a<��a<Ɛa<�a<3�a<x�a<��a<��a<��a<u�a<ڒa<�a<p�a<a<�a<v�a<��a<+�a<`�a<ʕa<:�a<��a<��a<H�a<ޗa< �a<��a<�a<b�a<�a<6�a<ʚa<�a<��a<��a<n�a<�a<m�a<��a<*�a<��a<1�a<��a<&�a<m�a<�a<F�a<�a<'�a<עa<R�a<n�a<
�a<C�a<ۤa<�a<��a<�a<T�a<¦a<��a<~�a<ۧa<*�a<q�a<��a<;�a<Y�a<ѩa<��a<O�a<��a<۪a<#�a<H�a<��a<��a<�a<F�a<��a<��a<Ŭa<�a<!�a<h�a<��a<��a<حa<ѭa< �a<�a<��a<k�a<k�a<��a<��a<ˮa<��a<��a<ڮa<�a<��a<�a<"�a<�a<�a<�a<�a<#�a<��a<�a<�a<�a<Ԯa<�a<®a<Ʈa<��a<��a<��a<o�a<f�a<&�a<�a<�a<˭a<٭a<��a<��a<A�a<#�a<��a<Ӭa<��a<k�a<W�a<�a<�a<��a<��a<_�a<�a<�a<��a<[�a<,�a<�a<��a<H�a<1�a<èa<��a<@�a<�a<��a<;�a<�a<��a<n�a<�a<��a<L�a<��a<��a<�a<գa<s�a<��a<��a<-�a<��a<W�a<�a<��a<b�a<�a<K�a<�a<u�a<:�a<��a<`�a<ٜa<r�a<�a<��a<A�a<ښa<f�a<�a<��a<C�a<��a<p�a<�a<��a<,�a<Жa<w�a<��a<ԕa<F�a<��a<��a<b�a<�a<��a<v�a<�a<גa<��a<@�a<�a<��a<��a<,�a<U�a<ܐa<��a<s�a<2�a<,�a<�a<�a<��a<��a<o�a<F�a<]�a<9�a</�a<�a<�a<�a<��a<�a<�a<�a<�a<9�a<(�a<O�a<h�a<f�a<�  �  ��a<��a<Ϗa<��a<#�a<H�a<k�a<��a<Ԑa<�a<D�a<��a<֑a<�a<0�a<z�a<�a<%�a<|�a<��a<�a<g�a<��a<�a<y�a<ؕa<1�a<��a<��a<g�a<a<!�a<��a<�a<m�a<��a<G�a<��a<�a<��a<�a<��a<�a<^�a<̝a<K�a<��a<7�a<��a<�a<z�a<�a<^�a<�a<H�a<��a<	�a<��a<�a<X�a<פa<*�a<��a<�a<c�a<��a<�a<l�a<̧a<�a<��a<ըa<�a<X�a<��a<	�a<U�a<��a<ߪa<�a<M�a<��a<ܫa<�a<;�a<v�a<��a<߬a<
�a<6�a<\�a<��a<��a<߭a<�a<)�a<"�a<5�a<K�a<��a<��a<��a<Ʈa<ɮa<�a<�a<��a<�a<�a<
�a<�a<�a<&�a<�a<�a<��a<�a<��a<�a<�a<�a<��a<��a<��a<��a<��a<k�a<R�a<A�a<$�a<�a<حa<ŭa<��a<��a<R�a<<�a<�a<��a<��a<o�a<k�a<&�a<��a<��a<��a<P�a<�a<ݪa<��a<i�a<#�a<ݩa<��a<g�a<�a<Ĩa<~�a<=�a<�a<��a<M�a<��a<��a<O�a<��a<��a<<�a<�a<��a<5�a<ԣa<y�a<�a<��a<;�a<�a<o�a<(�a<��a<(�a<��a<c�a<�a<��a<5�a<��a<U�a<ܜa<��a<�a<��a</�a<ʚa<W�a<�a<��a<%�a<��a<\�a<��a<��a<4�a<Ԗa<n�a<�a<��a<d�a<�a<��a<U�a<�a<��a<e�a<�a<̒a<��a<>�a<�a<��a<��a<7�a<��a<��a<��a<��a<B�a<'�a<�a<؏a<��a<��a<~�a<g�a<E�a<4�a<#�a<,�a<�a<�a<��a<�a<	�a<�a<�a</�a<'�a<G�a<[�a<��a<�  �  ~�a<ɏa<ɏa<��a<�a<>�a<��a<��a<�a<�a<C�a<u�a<��a<�a<D�a<��a<ǒa<�a<l�a<��a<�a<[�a<єa<
�a<|�a<̕a<?�a<��a<�a<f�a<��a<@�a<��a<��a<b�a<řa<H�a<��a<7�a<��a<�a<{�a<ܜa<~�a<Ɲa<W�a<��a<5�a<��a<�a<��a<�a<e�a<ša<P�a<��a<)�a<��a<�a<^�a<��a<8�a<��a<�a<h�a<��a<&�a<f�a<�a<�a<t�a<Ϩa<�a<��a<��a<
�a<=�a<��a<ܪa<�a<r�a<��a<ܫa< �a<K�a<��a<��a<�a<��a<H�a<S�a<��a<��a<˭a<�a<��a<K�a<P�a<t�a<��a<��a<��a<��a<ڮa<ծa<��a<�a< �a<�a<��a</�a<�a<�a<�a< �a<�a< �a<��a<�a<�a<ٮa<Ӯa<Ѯa<��a<��a<q�a<��a<L�a<B�a< �a<��a<�a<��a<��a<r�a<Q�a<!�a<�a<�a<��a<��a<E�a<�a<�a<��a<��a<C�a<)�a<Ϊa<��a<]�a<1�a<�a<��a<f�a< �a<�a<��a<7�a<�a<��a<N�a<��a<��a<R�a<��a<��a<6�a<	�a<��a<A�a<£a<w�a<�a<��a<P�a<֡a<v�a<��a<��a<H�a<ܟa<z�a<�a<��a< �a<ĝa<V�a<ߜa<��a<��a<��a<*�a<�a<V�a<�a<��a<$�a<Ԙa<T�a<��a<��a<#�a<іa<n�a<(�a<��a<c�a<��a<��a<i�a<��a<��a<R�a<+�a<a<��a<<�a<��a<��a<m�a<`�a<�a<�a<��a<f�a<E�a<�a<�a<ʏa<��a<��a<w�a<m�a<9�a<S�a<�a<$�a<�a<�a<�a<�a<�a<��a<�a<!�a<:�a<Z�a<J�a<��a<�  �  ��a<��a<Əa<��a<"�a<P�a<q�a<��a<Րa<	�a<P�a<��a<��a<��a<N�a<��a<ɒa</�a<s�a<��a<�a<_�a<��a<�a<|�a<a<'�a<��a<��a<U�a<��a<)�a<��a<�a<n�a<�a<C�a<��a<�a<��a<��a<|�a<�a<a�a<ŝa<F�a<��a<1�a<��a<�a<}�a<�a<v�a<ڡa<5�a<��a<$�a<��a<��a<s�a<Ǥa<(�a<��a<�a<[�a<��a<�a<g�a<̧a<&�a<|�a<Ĩa<�a<e�a<��a<�a<X�a<��a<ݪa<�a<V�a<��a<ͫa<�a<E�a<p�a<��a<�a<�a<2�a<W�a<��a<��a<ԭa<�a<
�a<&�a<S�a<b�a<m�a<��a<��a<��a<Ȯa<׮a<�a<��a<�a<�a< �a<�a<�a<�a<�a<�a<
�a<�a<��a<�a<�a<�a<Ǯa<��a<��a<��a<��a<p�a<I�a<5�a<#�a<	�a<ޭa<��a<��a<v�a<^�a<8�a<�a<Ԭa<��a<w�a<F�a<0�a<��a<��a<��a<G�a<�a<�a<��a<S�a<�a<�a<��a<U�a<�a<̨a<~�a<<�a<�a<��a<H�a<��a<��a<S�a<�a<��a<K�a<�a<��a<0�a<ԣa<s�a<�a<��a<>�a<١a<��a<�a<��a<?�a<ןa<]�a<�a<��a<%�a<��a<O�a<ܜa<z�a<�a<��a<+�a<˚a<c�a<��a<��a<'�a<��a<W�a<��a<��a<5�a<Ӗa<h�a<�a<��a<U�a<�a<��a<N�a<��a<��a<i�a<�a<ƒa<��a<;�a<�a<ϑa<x�a<;�a<�a<Ӑa<��a<}�a<V�a<�a<�a<̏a<��a<��a<}�a<\�a<;�a<9�a<0�a<�a<�a<�a<�a<�a<�a<�a<�a<,�a<-�a<J�a<S�a<w�a<�  �  ��a<��a<��a<��a<�a<F�a<g�a<��a<Аa<�a<7�a<��a<̑a<��a<M�a<��a<�a<�a<n�a<��a<�a<�a<��a<�a<p�a<�a<3�a<��a<�a<K�a<֗a<&�a<��a<��a<Y�a<�a<1�a<Ěa<�a<��a<�a<}�a<��a<I�a<�a<B�a<��a<"�a<��a<�a<{�a<��a<S�a<�a<J�a<��a<#�a<��a<�a<P�a<Ѥa<+�a<��a<�a<M�a<��a<�a<��a<��a<)�a<��a<Ȩa<1�a<[�a<ɩa<�a<U�a<��a<Ъa<(�a<Q�a<��a<īa<�a<:�a<r�a<��a<Ԭa<	�a<%�a<t�a<��a<��a<ԭa<�a<#�a<'�a<O�a<c�a<��a<��a<��a<Ȯa<Ǯa<�a<�a<��a<��a<	�a<#�a<��a<!�a<�a<�a<�a<�a<�a<�a<
�a<Ӯa<�a<ʮa<îa<��a<��a<��a<U�a<c�a<>�a<�a<��a<ԭa<׭a<��a<��a<F�a<0�a<�a<լa<��a<w�a<a�a<�a<�a<��a<�a<g�a<�a<۪a<��a<s�a<%�a<ҩa<��a<K�a<)�a<ɨa<��a<4�a<٧a<��a<7�a<�a<��a<`�a<��a<��a<O�a<դa<��a<+�a<ӣa<e�a<�a<��a<<�a<�a<d�a<�a<��a<@�a<֟a<j�a<�a<��a<0�a<��a<U�a<�a<k�a<�a<��a<K�a<��a<f�a<��a<��a<9�a<��a<h�a<�a<��a<%�a<Ɩa<|�a<�a<ȕa<L�a<�a<��a<Q�a<�a<��a<e�a<�a<�a<��a<@�a<�a<��a<��a<<�a<�a<Ԑa<��a<~�a<7�a<)�a<��a<�a<��a<��a<u�a<`�a<^�a<�a<3�a<�a<�a<�a<��a<�a<��a<%�a<�a<0�a<1�a<L�a<j�a<k�a<�  �  ��a<��a<ُa<��a<�a<F�a<|�a<��a<ϐa<�a<L�a<|�a<��a<�a<E�a<��a<͒a<�a<u�a<��a<�a<l�a<Ɣa<�a<q�a<ӕa<;�a<��a<��a<_�a<��a<�a<��a<��a<k�a<�a<H�a<��a< �a<��a<�a<v�a<�a<d�a<֝a<F�a<��a<+�a<��a<�a<��a<��a<m�a<͡a<F�a<��a<$�a<��a<�a<f�a<Ϥa<.�a<��a<�a<W�a<��a<�a<u�a<ѧa<(�a<u�a<ͨa<!�a<j�a<��a<�a<W�a<��a<תa<�a<S�a<��a<֫a<�a<J�a<~�a<��a<ڬa<
�a<8�a<g�a<��a<��a<խa<�a<�a<:�a<N�a<o�a<}�a<��a<��a<îa<Ǯa<�a<��a<��a<��a<�a<�a<�a<�a<�a<�a<�a<�a<�a<��a<�a<�a<ܮa<ɮa<��a<��a<��a<��a<o�a<\�a<5�a<�a< �a<�a<ŭa<��a<~�a<Z�a<'�a<��a<�a<��a<��a<J�a<�a<��a<��a<��a<U�a<�a<ܪa<��a<e�a<-�a<�a<��a<_�a<�a<¨a<��a<7�a<�a<��a<M�a<��a<��a<Q�a<��a<��a<I�a<�a<��a<0�a<ԣa<m�a<�a<��a<B�a<�a<~�a<�a<��a<B�a<ןa<m�a<��a<��a<.�a<��a<N�a<�a<v�a<�a<��a<8�a<Кa<d�a<�a<��a<)�a<��a<Z�a<��a<��a<1�a<͖a<n�a<
�a<��a<]�a<�a<��a<\�a<�a<��a<f�a<�a<גa<��a<?�a<�a<��a<y�a<P�a<�a<��a<��a<o�a<N�a<$�a<��a<Տa<��a<��a<v�a<Y�a<Q�a<<�a<&�a<�a<�a<�a<��a<�a<�a<�a<�a<%�a</�a<>�a<X�a<w�a<�  �  ��a<��a<ŏa<�a<'�a<<�a<w�a<��a<�a< �a<N�a<��a<��a<�a<*�a<��a<Βa<5�a<m�a<��a< �a<W�a<a<	�a<��a<ӕa<'�a<��a<�a<g�a<��a<6�a<��a<��a<h�a<��a<K�a<��a<=�a<��a<�a<��a<�a<_�a<ĝa<[�a<��a<$�a<��a<�a<��a<�a<|�a<ѡa<H�a<��a<�a<��a<�a<x�a<��a<4�a<��a<�a<R�a<��a<-�a<g�a<ǧa<�a<z�a<Ψa<�a<��a<��a<
�a<<�a<��a<٪a<�a<l�a<��a<ޫa<�a<@�a<n�a<��a<�a<��a<6�a<S�a<��a<��a<ɭa<�a<�a<8�a<5�a<i�a<~�a<��a<��a<��a<ݮa<ήa<�a<�a<�a<�a< �a<�a<�a<%�a<	�a<�a<�a< �a<	�a<خa<�a<֮a<ۮa<îa<��a<��a<s�a<p�a<H�a<E�a<(�a<��a<�a<��a<��a<l�a<\�a<8�a< �a<�a<��a<��a<L�a<6�a<�a<��a<��a<?�a<�a<ͪa<��a<d�a<�a<�a<��a<f�a<�a<٨a<��a<5�a<�a<��a<P�a<�a<��a<C�a<��a<��a<<�a<�a<�a<D�a<ˣa<f�a<�a<��a<N�a<ˡa<��a<
�a<��a<6�a<ǟa<n�a<��a<��a<�a<��a<N�a<ޜa<q�a<�a<��a<*�a<Śa<Y�a<��a<��a<�a<טa<L�a<��a<�a<(�a<ϖa<j�a<#�a<��a<e�a<��a<��a<L�a< �a<œa<U�a<�a<a<��a<=�a<��a<בa<v�a<N�a<��a<ڐa<��a<y�a<T�a<�a<�a<Ïa<��a<��a<}�a<m�a<;�a<<�a<�a<*�a<�a<�a<�a<�a<�a<�a< �a<�a<A�a<L�a<N�a<��a<�  �  ��a<��a<Ϗa<�a<�a<O�a<x�a<��a<ܐa<�a<=�a<��a<a<�a<R�a<��a<ђa<�a<n�a<a<�a<h�a<Ŕa< �a<q�a<ҕa<1�a<��a<��a<T�a<Ɨa</�a<��a<��a<p�a<ؙa<L�a<��a<$�a<��a<�a<t�a<��a<_�a<ӝa<E�a<��a<1�a<��a<�a<��a<��a<a�a<סa<F�a<��a<+�a<��a<��a<]�a<̤a<2�a<��a<��a<^�a<��a<�a<u�a<ʧa<.�a<v�a<˨a<"�a<q�a<��a<	�a<P�a<��a<֪a<�a<`�a<��a<ϫa<�a<L�a<w�a<��a<ڬa<�a<:�a<b�a<��a<��a<ҭa<�a<�a<3�a<Z�a<j�a<��a<��a<��a<��a<ծa<�a<�a< �a<�a<�a<�a<�a<�a<�a<�a<�a<�a<��a<�a<�a<�a<Үa<Ʈa<îa<��a<��a<��a<s�a<R�a<8�a<�a<�a<�a<­a<��a<x�a<L�a<+�a<�a<۬a<��a<��a<N�a<�a<�a<��a<��a<Q�a<�a<�a<��a<c�a<#�a<�a<��a<T�a<�a<Ҩa<z�a<3�a<�a<��a<Q�a<�a<��a<S�a<��a<��a<O�a<�a<��a<.�a<ңa<s�a<�a<��a<F�a<�a<r�a<�a<��a<C�a<ޟa<k�a<�a<��a<+�a<��a<L�a<�a<}�a<�a<��a<9�a<ɚa<k�a<��a<��a<+�a<Øa<O�a<��a<��a<4�a<˖a<e�a<�a<��a<W�a<�a<��a<U�a<�a<��a<j�a<�a<ђa<��a<B�a< �a<��a<�a<H�a<�a<ېa<��a<u�a<@�a<�a<��a<Տa<��a<��a<y�a<\�a<G�a<?�a<+�a<�a<�a<�a<��a<��a<�a<�a<�a<�a<,�a<L�a<_�a<j�a<�  �  ��a<��a<Ϗa<��a<$�a<T�a<_�a<��a<͐a<�a<K�a<��a<ʑa<�a<Z�a<z�a<�a<�a<z�a<ȓa<�a<s�a<��a<.�a<s�a<ѕa<.�a<��a<�a<R�a<ʗa<�a<��a<�a<e�a<יa<;�a<Ěa<�a<��a<�a<w�a<��a<N�a<ԝa<>�a<Ξa<$�a<��a<�a<w�a<
�a<[�a<�a<<�a<��a<%�a<~�a<�a<Q�a<ݤa<)�a<��a<��a<M�a<Φa<�a<u�a<��a<2�a<z�a<Ȩa<$�a<]�a<ʩa< �a<N�a<��a<ݪa<'�a<E�a<��a<ɫa<�a<E�a<p�a<��a<جa<�a<�a<i�a<��a<��a<�a<�a<#�a<�a<^�a<U�a<��a<��a<��a<Үa<��a<�a<ٮa<��a<�a<�a<�a<�a<,�a<�a<�a<�a<
�a<�a<��a<��a<�a<�a<Ϯa<��a<��a<��a<��a<^�a<R�a<5�a<%�a<�a<̭a<ҭa<��a<��a<Y�a<.�a<�a<Ŭa<ìa<p�a<b�a<�a<��a<ūa<��a<[�a<��a<�a<��a<b�a< �a<ݩa<��a<R�a<�a<��a<��a<>�a<�a<��a<@�a<�a<��a<T�a<��a<��a<Y�a<ڤa<��a<'�a<�a<f�a<	�a<��a<7�a<�a<l�a< �a<��a<8�a<؟a<Z�a<�a<��a<;�a<��a<Z�a<�a<l�a<"�a<��a<9�a<��a<n�a<��a<��a<,�a<��a<i�a<�a<��a<-�a<Җa<{�a<��a<��a<Q�a<�a<��a<N�a<�a<��a<z�a<�a<ؒa<��a<D�a<�a<��a<��a<4�a<�a<Ɛa<��a<�a<I�a<2�a<�a<�a<��a<��a<��a<[�a<G�a<(�a<?�a<�a<�a<�a<�a<�a< �a<�a<�a<0�a<5�a<9�a<b�a<k�a<�  �  ��a<��a<ُa<��a<�a<>�a<x�a<��a<ؐa<�a<J�a<z�a<ȑa<�a<R�a<��a<ܒa<�a<s�a<��a<�a<q�a<��a<�a<q�a<֕a<6�a<��a<�a<S�a<��a<7�a<��a<�a<f�a<ܙa<8�a<��a<7�a<��a< �a<~�a<�a<^�a<םa<L�a<��a<&�a<��a<�a<�a<��a<a�a<ѡa<K�a<��a<+�a<��a<��a<Z�a<Ȥa<)�a<��a<��a<W�a<��a<�a<v�a<̧a<�a<y�a<Ĩa<�a<�a<��a<��a<Q�a<��a<Ūa<�a<h�a<��a<̫a<	�a<=�a<}�a<��a<ڬa<��a<6�a<f�a<��a<��a<խa<�a<�a<.�a<\�a<m�a<��a<��a<��a<��a<ˮa<�a<�a<�a<��a<�a<�a<�a<�a<�a<�a<�a<�a<��a<��a<��a<�a<̮a<ٮa<Įa<��a<��a<{�a<h�a<\�a<@�a<�a<��a<�a<˭a<��a<r�a<X�a<&�a<�a<ݬa<��a<~�a<Y�a<!�a<��a<��a<��a<Y�a<�a<̪a<��a<g�a<(�a<ݩa<��a<R�a<�a<ڨa<��a<"�a<�a<��a<>�a<�a<��a<Q�a<�a<��a<>�a<�a<��a<5�a<£a<h�a<�a<��a<?�a<ݡa<r�a<
�a<��a<F�a<ޟa<k�a<��a<��a<'�a<��a<S�a<�a<v�a< �a<��a<:�a<˚a<X�a<��a<��a<$�a<јa<W�a<�a<��a<.�a<��a<r�a<�a<��a<S�a<��a<��a<[�a<�a<��a<V�a<�a<Ւa<��a<5�a<�a<��a<��a<C�a<�a<ސa<��a<q�a<K�a<�a<�a<ߏa<��a<��a<k�a<g�a<O�a<1�a<�a<�a<�a<�a<�a<��a< �a<�a<�a<�a<?�a<M�a<W�a<s�a<�  �  ��a<��a<Əa<��a<"�a<E�a<��a<��a<�a<��a<\�a<��a<��a<��a<3�a<��a<Вa<,�a<{�a<��a<�a<Y�a<ݔa<�a<��a<ϕa<-�a<��a<�a<f�a<��a<%�a<��a<�a<v�a<ڙa<]�a<��a<�a<��a<�a<��a<�a<r�a<��a<T�a<��a<@�a<��a<�a<��a<�a<�a<աa<K�a<��a<�a<��a<��a<x�a<Ĥa<5�a<��a<�a<r�a<��a<&�a<`�a<ܧa<�a<�a<Ѩa<�a<h�a<��a<�a<S�a<��a<�a<�a<X�a<��a<߫a<�a<E�a<|�a<��a<�a<��a<T�a<O�a<��a<��a<֭a<�a<�a<3�a<<�a<c�a<�a<��a<®a<��a<ܮa<Үa<��a< �a<��a<�a<�a<$�a<�a<�a<�a<�a<�a<��a<�a<�a<��a<׮a<��a<��a<��a<��a<w�a<}�a<I�a<>�a<#�a<��a<��a<��a<��a<h�a<j�a<4�a<�a<جa<��a<��a<M�a<.�a<��a<��a<��a<A�a<5�a<̪a<��a<`�a<�a<�a<��a<f�a<
�a<Ȩa<o�a<=�a<��a<��a<c�a<�a<��a<G�a<��a<��a<;�a<��a<{�a<=�a<ǣa<��a<�a<��a<M�a<ӡa<��a<�a<��a<2�a<şa<p�a<��a<��a<#�a<��a<H�a<ݜa<��a<�a<��a<#�a<ۚa<Y�a<��a<��a<�a<��a<C�a<�a<��a<:�a<֖a<[�a<�a<��a<g�a<�a<��a<[�a<��a<ēa<W�a<8�a<��a<��a<<�a<�a<ϑa<}�a<H�a<��a<Ԑa<��a<|�a<`�a<�a<�a<Ǐa<ŏa<��a<v�a<g�a<=�a<H�a<�a<$�a<	�a<�a<��a<��a<�a<
�a<'�a<�a<'�a<C�a<T�a<~�a<�  �  ��a<��a<ҏa<��a<$�a<F�a<s�a<��a<�a<�a<F�a<y�a<ʑa<�a<T�a<��a<�a<�a<r�a<��a<$�a<b�a<��a<�a<{�a<ؕa<4�a<��a<��a<S�a<ɗa<�a<��a<
�a<M�a<��a<6�a<ʚa<�a<��a<�a<x�a<�a<b�a<ӝa<I�a<��a<*�a<��a<�a<��a<��a<X�a<ءa<L�a<��a<(�a<��a<��a<N�a<ʤa<:�a<��a<�a<X�a<��a<�a<t�a<ԧa<�a<|�a<Ǩa<*�a<d�a<ѩa<��a<4�a<|�a<ݪa<1�a<Q�a<��a<ȫa<�a<9�a<��a<��a<�a<�a<4�a<V�a<��a<��a<ҭa<ޭa<�a<4�a<X�a<j�a<��a<��a<��a<��a<ݮa<�a<�a<��a<�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<߮a<Ѯa<�a<ٮa<��a<��a<��a<��a<d�a<U�a<@�a<%�a<��a<�a<��a<��a<|�a<T�a<$�a<�a<ܬa<��a<��a<^�a<�a<�a<��a<��a<K�a<�a<תa<��a<i�a<&�a<שa<��a<S�a<�a<¨a<��a<D�a<ͧa<��a<;�a<�a<��a<\�a<��a<��a<B�a<�a<��a<3�a<Σa<m�a<�a<��a<N�a<ߡa<i�a<�a<��a<E�a<۟a<o�a<�a<��a<(�a<Ɲa<^�a<ܜa<w�a<�a<��a<7�a<Қa<X�a<��a<��a<2�a<��a<p�a<�a<w�a<�a<Җa<��a<�a<��a<O�a<�a<��a<_�a<�a<��a<^�a<�a<Œa<��a<G�a< �a<��a<��a<I�a<�a<ېa<��a<r�a<D�a< �a<�a<Տa<��a<��a<�a<d�a<K�a<3�a<)�a<�a<�a<�a<�a<�a<��a<��a< �a<:�a<?�a<G�a<a�a<p�a<�  �  ��a<��a<�a<�a<�a<W�a<y�a<��a<ǐa<�a<K�a<z�a<ӑa<�a<U�a<t�a<�a<�a<��a<��a<�a<o�a<Ĕa<+�a<Y�a<˕a<<�a<��a<�a<B�a<Зa<�a<��a<�a<s�a<�a<(�a<Ěa<�a<��a<�a<��a<�a<N�a<�a</�a<��a<9�a<��a<�a<p�a<�a<S�a<�a<C�a<��a<!�a<��a<�a<N�a<�a<�a<��a<��a<g�a<��a<��a<�a<��a<�a<��a<��a<,�a<N�a<Ωa<�a<��a<��a<��a<�a<;�a<��a<��a<#�a<3�a<�a<��a<��a<�a<A�a<f�a<z�a<��a<�a<�a<(�a< �a<Z�a<_�a<��a<��a<��a<ٮa<��a<�a<�a<�a<��a<��a<!�a<��a<&�a<�a<�a<�a<�a<�a<�a<F�a<ݮa<Үa<��a<��a<��a<��a<��a<W�a<i�a<.�a<�a<�a<�a<ɭa<��a<��a<Y�a<%�a<�a<ˬa<��a<j�a<j�a<�a<�a<��a<y�a<W�a<�a<�a<��a<\�a<.�a<ҩa<��a<B�a<#�a<��a<��a<�a<�a<ܧa<.�a<�a<��a<Z�a<��a<��a<I�a<٤a<��a<�a<ңa<{�a<�a<��a<0�a<��a<d�a<�a<��a<=�a<ԟa<`�a<�a<��a<F�a<��a<J�a<�a<��a<�a<��a<B�a<��a<X�a<�a<�a<4�a<��a<m�a<ԗa<Ǘa<J�a<��a<s�a<�a<ɕa<A�a<�a<��a<]�a<�a<��a<s�a<$�a<Ւa<y�a<<�a<�a<��a<��a<5�a<�a<Аa<��a<v�a<E�a<:�a<�a<׏a<��a<��a<o�a<M�a<\�a<"�a<8�a<�a<�a<�a<�a<�a<��a<a�a<�a<�a<%�a<6�a<b�a<e�a<�  �  ��a<��a<ҏa<��a<$�a<F�a<s�a<��a<�a<�a<F�a<y�a<ʑa<�a<T�a<��a<�a<�a<r�a<��a<$�a<b�a<��a<�a<{�a<ؕa<4�a<��a<��a<S�a<ɗa<�a<��a<
�a<M�a<��a<6�a<ʚa<�a<��a<�a<x�a<�a<b�a<ӝa<I�a<��a<*�a<��a<�a<��a<��a<X�a<ءa<L�a<��a<(�a<��a<��a<N�a<ʤa<:�a<��a<�a<X�a<��a<�a<t�a<ԧa<�a<|�a<Ǩa<*�a<d�a<ѩa<��a<4�a<|�a<ݪa<1�a<Q�a<��a<ȫa<�a<9�a<��a<��a<�a<�a<4�a<V�a<��a<��a<ҭa<ޭa<�a<4�a<X�a<j�a<��a<��a<��a<��a<ݮa<�a<�a<��a<�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<߮a<Ѯa<�a<ٮa<��a<��a<��a<��a<d�a<U�a<@�a<%�a<��a<�a<��a<��a<|�a<T�a<$�a<�a<ܬa<��a<��a<^�a<�a<�a<��a<��a<K�a<�a<תa<��a<i�a<&�a<שa<��a<S�a<�a<¨a<��a<D�a<ͧa<��a<;�a<�a<��a<\�a<��a<��a<B�a<�a<��a<3�a<Σa<m�a<�a<��a<N�a<ߡa<i�a<�a<��a<E�a<۟a<o�a<�a<��a<(�a<Ɲa<^�a<ܜa<w�a<�a<��a<7�a<Қa<X�a<��a<��a<2�a<��a<p�a<�a<w�a<�a<Җa<��a<�a<��a<O�a<�a<��a<_�a<�a<��a<^�a<�a<Œa<��a<G�a< �a<��a<��a<I�a<�a<ېa<��a<r�a<D�a< �a<�a<Տa<��a<��a<�a<d�a<K�a<3�a<)�a<�a<�a<�a<�a<�a<��a<��a< �a<:�a<?�a<G�a<a�a<p�a<�  �  ��a<��a<Əa<��a<"�a<E�a<��a<��a<�a<��a<\�a<��a<��a<��a<3�a<��a<Вa<,�a<{�a<��a<�a<Y�a<ݔa<�a<��a<ϕa<-�a<��a<�a<f�a<��a<%�a<��a<�a<v�a<ڙa<]�a<��a<�a<��a<�a<��a<�a<r�a<��a<T�a<��a<@�a<��a<�a<��a<�a<�a<աa<K�a<��a<�a<��a<��a<x�a<Ĥa<5�a<��a<�a<r�a<��a<&�a<`�a<ܧa<�a<�a<Ѩa<�a<h�a<��a<�a<S�a<��a<�a<�a<X�a<��a<߫a<�a<E�a<|�a<��a<�a<��a<T�a<O�a<��a<��a<֭a<�a<�a<3�a<<�a<c�a<�a<��a<®a<��a<ܮa<Үa<��a< �a<��a<�a<�a<$�a<�a<�a<�a<�a<�a<��a<�a<�a<��a<׮a<��a<��a<��a<��a<w�a<}�a<I�a<>�a<#�a<��a<��a<��a<��a<h�a<j�a<4�a<�a<جa<��a<��a<M�a<.�a<��a<��a<��a<A�a<5�a<̪a<��a<`�a<�a<�a<��a<f�a<
�a<Ȩa<o�a<=�a<��a<��a<c�a<�a<��a<G�a<��a<��a<;�a<��a<{�a<=�a<ǣa<��a<�a<��a<M�a<ӡa<��a<�a<��a<2�a<şa<p�a<��a<��a<#�a<��a<H�a<ݜa<��a<�a<��a<#�a<ۚa<Y�a<��a<��a<�a<��a<C�a<�a<��a<:�a<֖a<[�a<�a<��a<g�a<�a<��a<[�a<��a<ēa<W�a<8�a<��a<��a<<�a<�a<ϑa<}�a<H�a<��a<Ԑa<��a<|�a<`�a<�a<�a<Ǐa<ŏa<��a<v�a<g�a<=�a<H�a<�a<$�a<	�a<�a<��a<��a<�a<
�a<'�a<�a<'�a<C�a<T�a<~�a<�  �  ��a<��a<ُa<��a<�a<>�a<x�a<��a<ؐa<�a<J�a<z�a<ȑa<�a<R�a<��a<ܒa<�a<s�a<��a<�a<q�a<��a<�a<q�a<֕a<6�a<��a<�a<S�a<��a<7�a<��a<�a<f�a<ܙa<8�a<��a<7�a<��a< �a<~�a<�a<^�a<םa<L�a<��a<&�a<��a<�a<�a<��a<a�a<ѡa<K�a<��a<+�a<��a<��a<Z�a<Ȥa<)�a<��a<��a<W�a<��a<�a<v�a<̧a<�a<y�a<Ĩa<�a<�a<��a<��a<Q�a<��a<Ūa<�a<h�a<��a<̫a<	�a<=�a<}�a<��a<ڬa<��a<6�a<f�a<��a<��a<խa<�a<�a<.�a<\�a<m�a<��a<��a<��a<��a<ˮa<�a<�a<�a<��a<�a<�a<�a<�a<�a<�a<�a<�a<��a<��a<��a<�a<̮a<ٮa<Įa<��a<��a<{�a<h�a<\�a<@�a<�a<��a<�a<˭a<��a<r�a<X�a<&�a<�a<ݬa<��a<~�a<Y�a<!�a<��a<��a<��a<Y�a<�a<̪a<��a<g�a<(�a<ݩa<��a<R�a<�a<ڨa<��a<"�a<�a<��a<>�a<�a<��a<Q�a<�a<��a<>�a<�a<��a<5�a<£a<h�a<�a<��a<?�a<ݡa<r�a<
�a<��a<F�a<ޟa<k�a<��a<��a<'�a<��a<S�a<�a<v�a< �a<��a<:�a<˚a<X�a<��a<��a<$�a<јa<W�a<�a<��a<.�a<��a<r�a<�a<��a<S�a<��a<��a<[�a<�a<��a<V�a<�a<Ւa<��a<5�a<�a<��a<��a<C�a<�a<ސa<��a<q�a<K�a<�a<�a<ߏa<��a<��a<k�a<g�a<O�a<1�a<�a<�a<�a<�a<�a<��a< �a<�a<�a<�a<?�a<M�a<W�a<s�a<�  �  ��a<��a<Ϗa<��a<$�a<T�a<_�a<��a<͐a<�a<K�a<��a<ʑa<�a<Z�a<z�a<�a<�a<z�a<ȓa<�a<s�a<��a<.�a<s�a<ѕa<.�a<��a<�a<R�a<ʗa<�a<��a<�a<e�a<יa<;�a<Ěa<�a<��a<�a<w�a<��a<N�a<ԝa<>�a<Ξa<$�a<��a<�a<w�a<
�a<[�a<�a<<�a<��a<%�a<~�a<�a<Q�a<ݤa<)�a<��a<��a<M�a<Φa<�a<u�a<��a<2�a<z�a<Ȩa<$�a<]�a<ʩa< �a<N�a<��a<ݪa<'�a<E�a<��a<ɫa<�a<E�a<p�a<��a<جa<�a<�a<i�a<��a<��a<�a<�a<#�a<�a<^�a<U�a<��a<��a<��a<Үa<��a<�a<ٮa<��a<�a<�a<�a<�a<,�a<�a<�a<�a<
�a<�a<��a<��a<�a<�a<Ϯa<��a<��a<��a<��a<^�a<R�a<5�a<%�a<�a<̭a<ҭa<��a<��a<Y�a<.�a<�a<Ŭa<ìa<p�a<b�a<�a<��a<ūa<��a<[�a<��a<�a<��a<b�a< �a<ݩa<��a<R�a<�a<��a<��a<>�a<�a<��a<@�a<�a<��a<T�a<��a<��a<Y�a<ڤa<��a<'�a<�a<f�a<	�a<��a<7�a<�a<l�a< �a<��a<8�a<؟a<Z�a<�a<��a<;�a<��a<Z�a<�a<l�a<"�a<��a<9�a<��a<n�a<��a<��a<,�a<��a<i�a<�a<��a<-�a<Җa<{�a<��a<��a<Q�a<�a<��a<N�a<�a<��a<z�a<�a<ؒa<��a<D�a<�a<��a<��a<4�a<�a<Ɛa<��a<�a<I�a<2�a<�a<�a<��a<��a<��a<[�a<G�a<(�a<?�a<�a<�a<�a<�a<�a< �a<�a<�a<0�a<5�a<9�a<b�a<k�a<�  �  ��a<��a<Ϗa<�a<�a<O�a<x�a<��a<ܐa<�a<=�a<��a<a<�a<R�a<��a<ђa<�a<n�a<a<�a<h�a<Ŕa< �a<q�a<ҕa<1�a<��a<��a<T�a<Ɨa</�a<��a<��a<p�a<ؙa<L�a<��a<$�a<��a<�a<t�a<��a<_�a<ӝa<E�a<��a<1�a<��a<�a<��a<��a<a�a<סa<F�a<��a<+�a<��a<��a<]�a<̤a<2�a<��a<��a<^�a<��a<�a<u�a<ʧa<.�a<v�a<˨a<"�a<q�a<��a<	�a<P�a<��a<֪a<�a<`�a<��a<ϫa<�a<L�a<w�a<��a<ڬa<�a<:�a<b�a<��a<��a<ҭa<�a<�a<3�a<Z�a<j�a<��a<��a<��a<��a<ծa<�a<�a< �a<�a<�a<�a<�a<�a<�a<�a<�a<�a<��a<�a<�a<�a<Үa<Ʈa<îa<��a<��a<��a<s�a<R�a<8�a<�a<�a<�a<­a<��a<x�a<L�a<+�a<�a<۬a<��a<��a<N�a<�a<�a<��a<��a<Q�a<�a<�a<��a<c�a<#�a<�a<��a<T�a<�a<Ҩa<z�a<3�a<�a<��a<Q�a<�a<��a<S�a<��a<��a<O�a<�a<��a<.�a<ңa<s�a<�a<��a<F�a<�a<r�a<�a<��a<C�a<ޟa<k�a<�a<��a<+�a<��a<L�a<�a<}�a<�a<��a<9�a<ɚa<k�a<��a<��a<+�a<Øa<O�a<��a<��a<4�a<˖a<e�a<�a<��a<W�a<�a<��a<U�a<�a<��a<j�a<�a<ђa<��a<B�a< �a<��a<�a<H�a<�a<ېa<��a<u�a<@�a<�a<��a<Տa<��a<��a<y�a<\�a<G�a<?�a<+�a<�a<�a<�a<��a<��a<�a<�a<�a<�a<,�a<L�a<_�a<j�a<�  �  ��a<��a<ŏa<�a<'�a<<�a<w�a<��a<�a< �a<N�a<��a<��a<�a<*�a<��a<Βa<5�a<m�a<��a< �a<W�a<a<	�a<��a<ӕa<'�a<��a<�a<g�a<��a<6�a<��a<��a<h�a<��a<K�a<��a<=�a<��a<�a<��a<�a<_�a<ĝa<[�a<��a<$�a<��a<�a<��a<�a<|�a<ѡa<H�a<��a<�a<��a<�a<x�a<��a<4�a<��a<�a<R�a<��a<-�a<g�a<ǧa<�a<z�a<Ψa<�a<��a<��a<
�a<<�a<��a<٪a<�a<l�a<��a<ޫa<�a<@�a<n�a<��a<�a<��a<6�a<S�a<��a<��a<ɭa<�a<�a<8�a<5�a<i�a<~�a<��a<��a<��a<ݮa<ήa<�a<�a<�a<�a< �a<�a<�a<%�a<	�a<�a<�a< �a<	�a<خa<�a<֮a<ۮa<îa<��a<��a<s�a<p�a<H�a<E�a<(�a<��a<�a<��a<��a<l�a<\�a<8�a< �a<�a<��a<��a<L�a<6�a<�a<��a<��a<?�a<�a<ͪa<��a<d�a<�a<�a<��a<f�a<�a<٨a<��a<5�a<�a<��a<P�a<�a<��a<C�a<��a<��a<<�a<�a<�a<D�a<ˣa<f�a<�a<��a<N�a<ˡa<��a<
�a<��a<6�a<ǟa<n�a<��a<��a<�a<��a<N�a<ޜa<q�a<�a<��a<*�a<Śa<Y�a<��a<��a<�a<טa<L�a<��a<�a<(�a<ϖa<j�a<#�a<��a<e�a<��a<��a<L�a< �a<œa<U�a<�a<a<��a<=�a<��a<בa<v�a<N�a<��a<ڐa<��a<y�a<T�a<�a<�a<Ïa<��a<��a<}�a<m�a<;�a<<�a<�a<*�a<�a<�a<�a<�a<�a<�a< �a<�a<A�a<L�a<N�a<��a<�  �  ��a<��a<ُa<��a<�a<F�a<|�a<��a<ϐa<�a<L�a<|�a<��a<�a<E�a<��a<͒a<�a<u�a<��a<�a<l�a<Ɣa<�a<q�a<ӕa<;�a<��a<��a<_�a<��a<�a<��a<��a<k�a<�a<H�a<��a< �a<��a<�a<v�a<�a<d�a<֝a<F�a<��a<+�a<��a<�a<��a<��a<m�a<͡a<F�a<��a<$�a<��a<�a<f�a<Ϥa<.�a<��a<�a<W�a<��a<�a<u�a<ѧa<(�a<u�a<ͨa<!�a<j�a<��a<�a<W�a<��a<תa<�a<S�a<��a<֫a<�a<J�a<~�a<��a<ڬa<
�a<8�a<g�a<��a<��a<խa<�a<�a<:�a<N�a<o�a<}�a<��a<��a<îa<Ǯa<�a<��a<��a<��a<�a<�a<�a<�a<�a<�a<�a<�a<�a<��a<�a<�a<ܮa<ɮa<��a<��a<��a<��a<o�a<\�a<5�a<�a< �a<�a<ŭa<��a<~�a<Z�a<'�a<��a<�a<��a<��a<J�a<�a<��a<��a<��a<U�a<�a<ܪa<��a<e�a<-�a<�a<��a<_�a<�a<¨a<��a<7�a<�a<��a<M�a<��a<��a<Q�a<��a<��a<I�a<�a<��a<0�a<ԣa<m�a<�a<��a<B�a<�a<~�a<�a<��a<B�a<ןa<m�a<��a<��a<.�a<��a<N�a<�a<v�a<�a<��a<8�a<Кa<d�a<�a<��a<)�a<��a<Z�a<��a<��a<1�a<͖a<n�a<
�a<��a<]�a<�a<��a<\�a<�a<��a<f�a<�a<גa<��a<?�a<�a<��a<y�a<P�a<�a<��a<��a<o�a<N�a<$�a<��a<Տa<��a<��a<v�a<Y�a<Q�a<<�a<&�a<�a<�a<�a<��a<�a<�a<�a<�a<%�a</�a<>�a<X�a<w�a<�  �  ��a<��a<��a<��a<�a<F�a<g�a<��a<Аa<�a<7�a<��a<̑a<��a<M�a<��a<�a<�a<n�a<��a<�a<�a<��a<�a<p�a<�a<3�a<��a<�a<K�a<֗a<&�a<��a<��a<Y�a<�a<1�a<Ěa<�a<��a<�a<}�a<��a<I�a<�a<B�a<��a<"�a<��a<�a<{�a<��a<S�a<�a<J�a<��a<#�a<��a<�a<P�a<Ѥa<+�a<��a<�a<M�a<��a<�a<��a<��a<)�a<��a<Ȩa<1�a<[�a<ɩa<�a<U�a<��a<Ъa<(�a<Q�a<��a<īa<�a<:�a<r�a<��a<Ԭa<	�a<%�a<t�a<��a<��a<ԭa<�a<#�a<'�a<O�a<c�a<��a<��a<��a<Ȯa<Ǯa<�a<�a<��a<��a<	�a<#�a<��a<!�a<�a<�a<�a<�a<�a<�a<
�a<Ӯa<�a<ʮa<îa<��a<��a<��a<U�a<c�a<>�a<�a<��a<ԭa<׭a<��a<��a<F�a<0�a<�a<լa<��a<w�a<a�a<�a<�a<��a<�a<g�a<�a<۪a<��a<s�a<%�a<ҩa<��a<K�a<)�a<ɨa<��a<4�a<٧a<��a<7�a<�a<��a<`�a<��a<��a<O�a<դa<��a<+�a<ӣa<e�a<�a<��a<<�a<�a<d�a<�a<��a<@�a<֟a<j�a<�a<��a<0�a<��a<U�a<�a<k�a<�a<��a<K�a<��a<f�a<��a<��a<9�a<��a<h�a<�a<��a<%�a<Ɩa<|�a<�a<ȕa<L�a<�a<��a<Q�a<�a<��a<e�a<�a<�a<��a<@�a<�a<��a<��a<<�a<�a<Ԑa<��a<~�a<7�a<)�a<��a<�a<��a<��a<u�a<`�a<^�a<�a<3�a<�a<�a<�a<��a<�a<��a<%�a<�a<0�a<1�a<L�a<j�a<k�a<�  �  ��a<��a<Əa<��a<"�a<P�a<q�a<��a<Րa<	�a<P�a<��a<��a<��a<N�a<��a<ɒa</�a<s�a<��a<�a<_�a<��a<�a<|�a<a<'�a<��a<��a<U�a<��a<)�a<��a<�a<n�a<�a<C�a<��a<�a<��a<��a<|�a<�a<a�a<ŝa<F�a<��a<1�a<��a<�a<}�a<�a<v�a<ڡa<5�a<��a<$�a<��a<��a<s�a<Ǥa<(�a<��a<�a<[�a<��a<�a<g�a<̧a<&�a<|�a<Ĩa<�a<e�a<��a<�a<X�a<��a<ݪa<�a<V�a<��a<ͫa<�a<E�a<p�a<��a<�a<�a<2�a<W�a<��a<��a<ԭa<�a<
�a<&�a<S�a<b�a<m�a<��a<��a<��a<Ȯa<׮a<�a<��a<�a<�a< �a<�a<�a<�a<�a<�a<
�a<�a<��a<�a<�a<�a<Ǯa<��a<��a<��a<��a<p�a<I�a<5�a<#�a<	�a<ޭa<��a<��a<v�a<^�a<8�a<�a<Ԭa<��a<w�a<F�a<0�a<��a<��a<��a<G�a<�a<�a<��a<S�a<�a<�a<��a<U�a<�a<̨a<~�a<<�a<�a<��a<H�a<��a<��a<S�a<�a<��a<K�a<�a<��a<0�a<ԣa<s�a<�a<��a<>�a<١a<��a<�a<��a<?�a<ןa<]�a<�a<��a<%�a<��a<O�a<ܜa<z�a<�a<��a<+�a<˚a<c�a<��a<��a<'�a<��a<W�a<��a<��a<5�a<Ӗa<h�a<�a<��a<U�a<�a<��a<N�a<��a<��a<i�a<�a<ƒa<��a<;�a<�a<ϑa<x�a<;�a<�a<Ӑa<��a<}�a<V�a<�a<�a<̏a<��a<��a<}�a<\�a<;�a<9�a<0�a<�a<�a<�a<�a<�a<�a<�a<�a<,�a<-�a<J�a<S�a<w�a<�  �  ~�a<ɏa<ɏa<��a<�a<>�a<��a<��a<�a<�a<C�a<u�a<��a<�a<D�a<��a<ǒa<�a<l�a<��a<�a<[�a<єa<
�a<|�a<̕a<?�a<��a<�a<f�a<��a<@�a<��a<��a<b�a<řa<H�a<��a<7�a<��a<�a<{�a<ܜa<~�a<Ɲa<W�a<��a<5�a<��a<�a<��a<�a<e�a<ša<P�a<��a<)�a<��a<�a<^�a<��a<8�a<��a<�a<h�a<��a<&�a<f�a<�a<�a<t�a<Ϩa<�a<��a<��a<
�a<=�a<��a<ܪa<�a<r�a<��a<ܫa< �a<K�a<��a<��a<�a<��a<H�a<S�a<��a<��a<˭a<�a<��a<K�a<P�a<t�a<��a<��a<��a<��a<ڮa<ծa<��a<�a< �a<�a<��a</�a<�a<�a<�a< �a<�a< �a<��a<�a<�a<ٮa<Ӯa<Ѯa<��a<��a<q�a<��a<L�a<B�a< �a<��a<�a<��a<��a<r�a<Q�a<!�a<�a<�a<��a<��a<E�a<�a<�a<��a<��a<C�a<)�a<Ϊa<��a<]�a<1�a<�a<��a<f�a< �a<�a<��a<7�a<�a<��a<N�a<��a<��a<R�a<��a<��a<6�a<	�a<��a<A�a<£a<w�a<�a<��a<P�a<֡a<v�a<��a<��a<H�a<ܟa<z�a<�a<��a< �a<ĝa<V�a<ߜa<��a<��a<��a<*�a<�a<V�a<�a<��a<$�a<Ԙa<T�a<��a<��a<#�a<іa<n�a<(�a<��a<c�a<��a<��a<i�a<��a<��a<R�a<+�a<a<��a<<�a<��a<��a<m�a<`�a<�a<�a<��a<f�a<E�a<�a<�a<ʏa<��a<��a<w�a<m�a<9�a<S�a<�a<$�a<�a<�a<�a<�a<�a<��a<�a<!�a<:�a<Z�a<J�a<��a<�  �  ��a<��a<Ϗa<��a<#�a<H�a<k�a<��a<Ԑa<�a<D�a<��a<֑a<�a<0�a<z�a<�a<%�a<|�a<��a<�a<g�a<��a<�a<y�a<ؕa<1�a<��a<��a<g�a<a<!�a<��a<�a<m�a<��a<G�a<��a<�a<��a<�a<��a<�a<^�a<̝a<K�a<��a<7�a<��a<�a<z�a<�a<^�a<�a<H�a<��a<	�a<��a<�a<X�a<פa<*�a<��a<�a<c�a<��a<�a<l�a<̧a<�a<��a<ըa<�a<X�a<��a<	�a<U�a<��a<ߪa<�a<M�a<��a<ܫa<�a<;�a<v�a<��a<߬a<
�a<6�a<\�a<��a<��a<߭a<�a<)�a<"�a<5�a<K�a<��a<��a<��a<Ʈa<ɮa<�a<�a<��a<�a<�a<
�a<�a<�a<&�a<�a<�a<��a<�a<��a<�a<�a<�a<��a<��a<��a<��a<��a<k�a<R�a<A�a<$�a<�a<حa<ŭa<��a<��a<R�a<<�a<�a<��a<��a<o�a<k�a<&�a<��a<��a<��a<P�a<�a<ݪa<��a<i�a<#�a<ݩa<��a<g�a<�a<Ĩa<~�a<=�a<�a<��a<M�a<��a<��a<O�a<��a<��a<<�a<�a<��a<5�a<ԣa<y�a<�a<��a<;�a<�a<o�a<(�a<��a<(�a<��a<c�a<�a<��a<5�a<��a<U�a<ܜa<��a<�a<��a</�a<ʚa<W�a<�a<��a<%�a<��a<\�a<��a<��a<4�a<Ԗa<n�a<�a<��a<d�a<�a<��a<U�a<�a<��a<e�a<�a<̒a<��a<>�a<�a<��a<��a<7�a<��a<��a<��a<��a<B�a<'�a<�a<؏a<��a<��a<~�a<g�a<E�a<4�a<#�a<,�a<�a<�a<��a<�a<	�a<�a<�a</�a<'�a<G�a<[�a<��a<�  �  �a<�a<�a<7�a<C�a<��a<��a<�a<�a<Q�a<j�a<őa<�a</�a<��a<��a<+�a<X�a<��a<��a<<�a<��a<�a<p�a<��a< �a<r�a<Жa<Q�a<q�a<�a<s�a<Ԙa<-�a<��a<�a<b�a<��a<Y�a<��a<3�a<��a<8�a<��a<�a<q�a<�a<d�a<��a<E�a<��a<0�a<{�a<�a<q�a<�a<g�a<��a<:�a<w�a<��a<L�a<��a<�a<��a<�a<3�a<��a<��a<b�a<��a<�a<{�a<��a<��a<�a<v�a<��a<��a<T�a<��a<�a<�a<V�a<{�a<��a<�a<�a<O�a<Y�a<��a<��a<ԭa<�a<�a<Z�a<D�a<��a<��a<��a<ͮa<��a<�a<�a<�a<��a<=�a<!�a<7�a<L�a<4�a<c�a<0�a<F�a<c�a<:�a<<�a<
�a</�a<��a<�a<��a<�a<�a<��a<Ӯa<��a<��a<m�a<5�a<L�a<��a<�a<��a<��a<j�a<b�a<=�a<��a<�a<��a<��a<L�a<�a<�a<��a<|�a<9�a<(�a<��a<��a<Y�a<�a<�a<f�a<c�a<�a<��a<]�a<��a<̧a<_�a<4�a<Ѧa<��a<�a<ѥa<��a<�a<Ԥa<V�a<��a<��a<*�a<ڢa<a�a<�a<��a<U�a<Ԡa<x�a<�a<��a<D�a<��a<`�a<ݝa<��a<�a<��a<E�a<śa<��a<�a<��a<9�a<��a<��a<��a<��a<�a<ėa<U�a<��a<��a<T�a<�a<u�a<Y�a<�a<��a<Z�a<ғa<��a<J�a<�a<��a<w�a<,�a<�a<בa<h�a<x�a<�a<�a<��a<m�a<c�a<#�a<�a<Տa<�a<��a<��a<��a<h�a<��a<E�a<R�a<l�a<D�a<L�a<$�a<Z�a<3�a<h�a<t�a<��a<��a<��a<�  �  Ǐa<�a< �a<9�a<\�a<��a<��a<��a<�a<[�a<��a<��a<��a<4�a<x�a<��a<�a<]�a<��a<
�a<N�a<��a<��a<P�a<��a<�a<V�a<��a</�a<��a<�a<M�a<Ęa<;�a<��a<!�a<�a<��a<P�a<��a<+�a<��a<�a<��a<��a<��a<�a<a�a<؟a<O�a<��a<8�a<��a<�a<t�a<Ԣa<D�a<��a<*�a<��a<	�a<a�a<˥a<-�a<��a<�a<U�a<��a<�a<C�a<��a<�a<=�a<��a<�a<6�a<��a<̪a<�a<F�a<u�a<��a<��a<=�a<c�a<��a<׬a<�a<5�a<d�a<��a<��a<�a<�a<$�a<E�a<S�a<q�a<��a<��a<®a<�a<��a<��a<�a<�a<%�a<-�a<>�a</�a<9�a<;�a<K�a<1�a<,�a<4�a<A�a<1�a<=�a<�a<�a<��a<׮a<ʮa<ˮa<��a<��a<t�a<o�a<N�a<-�a<�a<�a<έa<��a<��a<[�a<6�a<��a<Ԭa<��a<��a<Q�a<)�a<��a<��a<��a<D�a<�a<֪a<��a<=�a<�a<ͩa<��a<5�a<�a<��a<k�a<!�a<ܧa<|�a<0�a<Ȧa<o�a<�a<եa<k�a<�a<��a<p�a<��a<��a<B�a<�a<u�a< �a<��a<A�a<֠a<`�a<��a<��a<4�a<˞a<l�a<�a<��a<�a<��a<>�a<�a<c�a<�a<��a<0�a<��a<P�a<�a<��a<1�a<ٗa<r�a<�a<��a<8�a<�a<��a<@�a<ؔa<{�a<>�a<��a<��a<U�a<�a<ƒa<��a<H�a<��a<a<w�a<A�a<�a<�a<��a<��a<l�a<7�a<#�a<�a<яa<��a<��a<z�a<m�a<]�a<`�a<=�a<4�a<>�a<Q�a<K�a<g�a<[�a<n�a<k�a<o�a<��a<��a<�  �  ��a<�a< �a</�a<f�a<p�a<Őa<Ґa<�a<9�a<��a<��a<��a<Z�a<t�a<�a<��a<X�a<��a<�a<D�a<��a<
�a<8�a<ŕa<��a<m�a<ۖa<�a<��a<�a<s�a<Θa</�a<��a<��a<}�a<�a<t�a<̛a<G�a<��a<�a<��a<�a<��a<۞a<\�a<֟a<1�a<��a<�a<��a<�a<��a<�a<S�a<Уa<�a<��a<�a<X�a<��a<#�a<��a<Цa<]�a<��a<�a<K�a<��a<	�a<H�a<��a<�a<1�a<m�a<��a< �a<G�a<��a<��a<�a<+�a<y�a<��a<Ƭa<"�a<�a<q�a<��a<��a<֭a<�a<#�a</�a<}�a<p�a<��a<��a<��a<�a<׮a<��a<��a<+�a<�a<.�a<7�a<+�a<f�a<�a<a�a<@�a<F�a<L�a<,�a<0�a<�a<�a<�a<�a<��a<Ԯa<�a<��a<��a<t�a<e�a<Y�a<�a<#�a<߭a<ɭa<��a<��a<N�a<-�a<&�a<Ьa<Ϭa<o�a<L�a<�a<�a<��a<r�a<V�a<�a<�a<��a<T�a<�a<��a<��a<<�a<�a<��a<_�a<�a<��a<z�a<!�a<�a<~�a<1�a<�a<e�a<>�a<��a<q�a<�a<��a<A�a<Ţa<o�a<��a<��a<,�a<�a<x�a<�a<��a<�a<Ӟa<G�a<�a<s�a<�a<��a<*�a<�a<O�a<�a<��a<5�a<ԙa<Z�a<�a<��a<,�a<��a<`�a<�a<��a<_�a<�a<��a<.�a<�a<��a<-�a<�a<��a<b�a< �a<��a<y�a</�a<��a<��a<��a<@�a<+�a<�a<��a<��a<G�a<1�a<��a<�a<Ïa<��a<��a<u�a<��a<A�a<v�a<M�a<O�a<V�a<<�a<K�a<;�a<V�a<[�a<��a<��a<��a<Տa<�  �  ďa<��a<�a<8�a<X�a<��a<a<ϐa<2�a<R�a<~�a<ӑa<��a<>�a<x�a<Ȓa<�a<r�a<��a<
�a<_�a<��a<�a<R�a<��a<�a<t�a<ǖa<*�a<��a<�a<c�a<��a<;�a<��a<�a<��a<�a<L�a<Лa<1�a<��a<�a<��a<�a<~�a<�a<k�a<ٟa<E�a<Ԡa<(�a<��a<�a<o�a<ۢa<F�a<��a<(�a<��a<��a<z�a<ͥa<+�a<��a<�a<F�a<��a<�a<B�a<��a<�a<L�a<��a<ߩa<;�a<��a<ʪa<�a<>�a<��a<��a<��a<5�a<h�a<��a<֬a<�a<5�a<u�a<��a<ĭa<�a<��a<4�a<@�a<^�a<r�a<��a<��a<Үa<֮a<�a<�a<��a<&�a<*�a<.�a<<�a<>�a<E�a<4�a<F�a<5�a<J�a<&�a<3�a<;�a<!�a<$�a<�a<�a<��a<ˮa<Ȯa<��a<��a<��a<m�a<J�a<1�a<!�a<ܭa<�a<��a<~�a<p�a</�a<	�a<Ԭa<��a<~�a<g�a<�a<��a<ƫa<p�a<Z�a<
�a<̪a<��a<Z�a<�a<ɩa<��a<;�a<��a<��a<j�a< �a<Чa<��a<�a<Ħa<��a<�a<ѥa<e�a<#�a<��a<c�a<�a<��a<C�a<ڢa<��a<�a<��a<G�a<Ҡa<g�a<��a<��a<2�a<Ҟa<Y�a<�a<��a<�a<��a<B�a<כa<e�a<�a<��a<.�a<��a<^�a<�a<��a<5�a<ӗa<p�a<�a<��a<H�a<�a<��a<8�a<ޔa<��a<=�a<�a<��a<f�a<�a<Ғa<��a<4�a<�a<��a<��a<B�a<�a<ސa<��a<��a<`�a<S�a<�a<��a<֏a<��a<��a<��a<y�a<V�a<[�a<A�a<S�a<0�a<C�a<U�a<L�a<c�a<f�a<^�a<��a<��a<��a<�  �  �a<؏a<�a<7�a<V�a<��a<��a<�a<�a<P�a<w�a<őa<��a<<�a<��a<a<�a<X�a<��a<��a<F�a<��a<�a<Y�a<��a<�a<k�a<��a<H�a<��a<�a<X�a<˘a<@�a<��a<�a<q�a<�a<L�a<�a<9�a<��a<)�a<��a<�a<m�a<�a<R�a<Οa<C�a<��a<+�a<��a<�a<v�a<�a<Y�a<��a<.�a<~�a<��a<U�a<��a<%�a<z�a<�a<5�a<��a<�a<P�a<��a<��a<a�a<��a<��a<)�a<x�a<��a<�a<O�a<|�a<٫a<�a<S�a<f�a<��a<�a<��a<@�a<Z�a<��a<��a<խa<��a<�a<F�a<Y�a<��a<��a<��a<ʮa<Ȯa<�a<��a<�a<�a< �a<-�a<3�a<H�a<)�a<X�a<E�a<C�a<L�a<-�a<P�a<�a<&�a<�a<%�a<�a<�a<�a<��a<ʮa<��a<��a<m�a<H�a<0�a<�a<��a<ĭa<��a<w�a<b�a<6�a<�a<�a<��a<��a<M�a<�a<�a<��a<��a<=�a<�a<Ūa<��a<Q�a<�a<�a<w�a<U�a<�a<��a<p�a<�a<ȧa<n�a<C�a<Ŧa<��a<#�a<ޥa<}�a<�a<Фa<R�a<�a<��a<8�a<آa<i�a<�a<��a<G�a<ؠa<v�a<�a<��a<8�a<��a<[�a<�a<�a<�a<��a<I�a<ƛa<�a<��a<��a<@�a<��a<s�a<�a<��a<#�a<Ɨa<[�a<	�a<��a<?�a<�a<��a<V�a<ܔa<��a<N�a<�a<��a<K�a<�a<��a<x�a<5�a<�a<Ña<}�a<W�a<�a<�a<��a<v�a<a�a<,�a<�a<�a<̏a<��a<��a<��a<]�a<z�a<Y�a<O�a<U�a<7�a<`�a<:�a<P�a<J�a<}�a<f�a<��a<��a<��a<�  �  ˏa<��a<�a<�a<k�a<��a<��a<�a<�a<N�a<��a<��a< �a<E�a<u�a<ђa<�a<V�a<��a<��a<H�a<��a<�a<Z�a<��a<�a<n�a<Җa<&�a<��a<�a<\�a<Әa<5�a<��a<�a<m�a<��a<Z�a<ʛa<8�a<��a<"�a<��a<�a<l�a<��a<^�a<ӟa<G�a<��a<-�a<��a<�a<{�a<ݢa<I�a<ģa<%�a<��a< �a<Z�a<��a<)�a<��a<��a<:�a<��a<�a<T�a<��a<��a<I�a<��a<�a<$�a<��a<Ūa<�a<N�a<��a<ȫa<��a<0�a<t�a<��a<Ƭa<	�a<@�a<\�a<��a<��a<ݭa<
�a<"�a<D�a<h�a<r�a<��a<��a<��a<�a<�a<�a<�a<�a<'�a<?�a< �a<;�a<L�a<B�a<;�a<>�a<>�a<B�a<7�a<�a<<�a<�a<�a<�a<�a<ݮa<��a<��a<��a<��a<P�a<]�a<5�a<�a<��a<��a<��a<��a<T�a<7�a<�a<Ѭa<��a<��a<J�a<,�a<�a<��a<��a<<�a<�a<תa<y�a<U�a<�a<ũa<~�a<I�a<��a<��a<d�a<�a<٧a<j�a<1�a<Ҧa<}�a<"�a<ȥa<v�a<'�a<��a<Q�a<�a<��a<=�a<ܢa<m�a<�a<��a<=�a<ݠa<i�a<��a<��a</�a<͞a<c�a<�a<��a<�a<��a<N�a<̛a<d�a<
�a<��a<%�a<��a<[�a<�a<��a<�a<֗a<k�a<�a<��a<E�a<�a<��a<3�a<�a<��a<-�a<�a<��a<N�a<�a<��a<��a<G�a<��a<��a<��a<B�a<�a<�a<��a<��a<^�a<'�a<�a<�a<ӏa<ŏa<��a<��a<��a<d�a<P�a<J�a<G�a<L�a<G�a<3�a<f�a<D�a<c�a<|�a<��a<��a<��a<�  �  ʏa<�a<�a<5�a<[�a<��a<��a<��a<)�a<H�a<��a<��a<��a<I�a<��a<͒a<
�a<]�a<��a<��a<\�a<��a<�a<L�a<��a<�a<l�a<ʖa<.�a<��a<�a<a�a<Øa<4�a<��a<�a<��a<�a<^�a<��a<L�a<��a<�a<��a<��a<��a<�a<f�a<Пa<C�a<Πa<�a<��a<��a<{�a<�a<V�a<��a<�a<��a<�a<t�a<ǥa<$�a<��a<�a<Q�a<��a< �a<M�a<��a<�a<<�a<��a<ܩa<6�a<�a<ƪa<�a<?�a<��a<��a<�a<6�a<n�a<��a<Ӭa<�a<.�a<k�a<��a<��a<�a<�a<#�a<7�a<d�a<��a<��a<��a<��a<خa<�a<�a<�a<�a<%�a<-�a<?�a<7�a<F�a<:�a<T�a<E�a<7�a<:�a</�a<2�a<&�a<!�a<�a<��a<�a<ٮa<ڮa<��a<��a<�a<k�a<M�a<.�a<�a<�a<�a<��a<��a<Z�a<0�a<�a<�a<��a<z�a<Q�a<�a<�a<īa<v�a<M�a<�a<٪a<��a<R�a<�a<ͩa<��a<8�a<��a<��a<d�a< �a<Χa<}�a<�a<֦a<p�a<6�a<٥a<l�a<#�a<��a<k�a<��a<��a<:�a<آa<��a<�a<��a<9�a<ݠa<t�a<�a<��a<(�a<ʞa<L�a<�a<��a<�a<��a<:�a<�a<c�a<�a<��a<1�a<ؙa<N�a<��a<��a<0�a<͗a<m�a<	�a<��a<K�a<��a<��a<9�a<�a<��a<:�a<��a<��a<\�a<�a<ϒa<��a<.�a<��a<��a<��a<Q�a<�a<��a<��a<��a<T�a<L�a<�a<�a<Џa<��a<��a<��a<z�a<\�a<i�a<Q�a<@�a<D�a<?�a<M�a<Q�a<`�a<_�a<p�a<�a<��a<Əa<�  �  ۏa<�a<�a<B�a<A�a<��a<��a<ސa<�a<O�a<��a<ɑa<��a</�a<��a<��a<�a<c�a<��a<��a<E�a<��a<�a<P�a<��a<�a<k�a<Ŗa<9�a<��a<��a<p�a<Řa<6�a<��a<�a<��a<�a<^�a<כa<@�a<��a<&�a<��a<�a<y�a<ߞa<f�a<ןa<<�a<��a<)�a<��a<�a<p�a<�a<]�a<��a<2�a<��a<��a<X�a<��a<*�a<��a<ަa<<�a<��a<��a<U�a<��a<��a<S�a<��a<�a<:�a<q�a<��a<�a<C�a<��a<ȫa<��a<>�a<o�a<��a<�a<��a<3�a<o�a<��a<��a<ԭa<��a<"�a<J�a<N�a<��a<��a<��a<ͮa<Ӯa<�a<�a<�a<!�a<(�a<�a<B�a<C�a<6�a<K�a<;�a<D�a<M�a<3�a<8�a<6�a<�a<!�a<�a<��a<��a<ݮa<��a<��a<��a<��a<x�a<3�a<2�a<�a<�a<ía<��a<��a<f�a<4�a<��a<��a<��a<��a<W�a<�a<�a<��a<}�a<P�a<�a<��a<��a<Q�a<	�a<ةa<{�a<D�a<	�a<��a<f�a<�a<��a<��a<)�a<֦a<��a<*�a<ͥa<z�a<�a<Ȥa<^�a<�a<��a<A�a<Ѣa<m�a<�a<��a<I�a<Ҡa<v�a<�a<��a<<�a<a<Z�a<�a<|�a<�a<��a<8�a<Λa<x�a<��a<��a<*�a<Ùa<e�a<��a<��a<4�a<��a<a�a<
�a<��a<U�a<�a<��a<@�a<�a<��a<L�a<ݓa<��a<`�a<	�a<��a<x�a<:�a<��a<Ǒa<r�a<]�a<�a<�a<��a<��a<b�a<*�a<
�a<��a<ӏa<��a<��a<��a<i�a<m�a<P�a<Q�a<V�a<=�a<H�a<Q�a<?�a<_�a<g�a<j�a<��a<��a<��a<�  �  ҏa<�a<�a<-�a<a�a<��a<��a<��a<	�a<V�a<��a<��a<�a<2�a<��a<��a<-�a<O�a<��a<��a<T�a<��a<�a<a�a<��a<�a<c�a<Ėa<2�a<��a<��a<O�a<јa<6�a<��a<�a<x�a<�a<N�a<Ǜa<6�a<��a<%�a<��a<�a<m�a< �a<[�a<˟a<]�a<��a<>�a<��a<�a<u�a<ڢa<M�a<��a<<�a<��a<�a<W�a<ץa<#�a<~�a<��a<5�a<��a<�a<Q�a<��a<�a<H�a<��a<�a<0�a<��a<ƪa<�a<M�a<t�a<ɫa<��a<9�a<j�a<��a<ڬa<��a<H�a<R�a<��a<��a<حa<�a<�a<^�a<T�a<{�a<��a<��a<��a<Үa<��a<�a<$�a<	�a<(�a<5�a<.�a<A�a<9�a<G�a<<�a<B�a<5�a<;�a<7�a<(�a<.�a<�a<�a<�a<�a<ޮa<��a<��a<��a<��a<b�a<S�a<6�a<��a<�a<��a<��a<��a<R�a<L�a<��a<�a<��a<��a<C�a<-�a<�a<��a<��a<0�a<�a<Ǫa<��a<I�a<�a<Щa<��a<H�a<�a<��a<f�a<�a<ԧa<u�a<,�a<Ʀa<y�a< �a<ǥa<y�a<�a<Ȥa<R�a<�a<��a<5�a<�a<j�a<&�a<��a<M�a<ؠa<e�a<�a<��a<F�a<��a<r�a<�a<��a<�a<��a<V�a<Ǜa<u�a<��a<��a<&�a<��a<Z�a<�a<��a<*�a<їa<l�a<�a<��a<7�a<�a<��a<<�a<��a<��a<A�a<�a<��a<C�a<�a<ϒa<{�a<P�a<�a<ۑa<x�a<K�a<
�a<�a<��a<�a<n�a<#�a<)�a<ߏa<ԏa<��a<��a<��a<m�a<h�a<P�a<O�a<>�a<E�a<G�a<B�a<X�a<R�a<e�a<w�a<x�a<��a<��a<�  �  ��a<��a<�a<0�a<_�a<��a<��a<ڐa<�a<?�a<��a<��a<�a<I�a<��a<֒a<�a<H�a<��a<�a<P�a<��a<�a<U�a<��a<�a<q�a<זa<#�a<��a<��a<`�a<՘a</�a<��a<�a<y�a<�a<m�a<śa<T�a<��a<�a<��a<�a<x�a<�a<h�a<ɟa<A�a<��a<$�a<��a< �a<��a<�a<\�a<ƣa< �a<��a<��a<V�a<åa<�a<��a<�a<E�a<��a<�a<S�a<��a<�a<H�a<��a<�a<+�a<p�a<��a<��a<N�a<��a<ūa<�a<6�a<x�a<��a<ڬa<�a<4�a<l�a<}�a<��a<ϭa<�a<�a<:�a<i�a<��a<��a<��a<��a<ݮa<�a<��a<�a<�a<+�a<0�a<3�a<;�a<U�a<1�a<W�a<O�a<5�a<R�a</�a<-�a<�a<�a<�a<�a<�a<�a<�a<��a<��a<��a<e�a<Q�a</�a<�a<�a<ͭa<��a<��a<K�a<8�a<�a<ެa<��a<}�a<<�a<'�a<ݫa<��a<n�a<L�a<�a<ժa<��a<X�a<�a<��a<��a<E�a<��a<��a<_�a<�a<��a<v�a<&�a<�a<x�a<?�a<ݥa<p�a<*�a<��a<]�a<��a<��a<4�a<֢a<n�a<�a<��a<9�a<�a<z�a<�a<��a<*�a<��a<Z�a<�a<��a<�a<��a<;�a<֛a<k�a<�a<��a<:�a<��a<Z�a<�a<��a<%�a<��a<`�a<��a<��a<M�a<�a<��a<8�a<�a<��a<A�a<��a<��a<]�a<��a<Œa<r�a<A�a<�a<��a<��a<O�a<�a<�a<��a<��a<T�a<3�a<�a<�a<׏a<��a<��a<��a<��a<S�a<k�a<[�a<>�a<\�a<?�a<G�a<C�a<W�a<]�a<��a<}�a<��a<͏a<�  �  ��a< �a<��a<C�a<S�a<z�a<Аa<��a<8�a<D�a<��a<̑a<��a<<�a<q�a<̒a<
�a<p�a<��a<��a<h�a<��a<�a<?�a<��a<�a<a�a<ۖa<�a<��a<�a<p�a<��a<9�a<��a<�a<��a<ؚa<`�a<��a<9�a<��a<�a<��a<�a<��a<ٞa<q�a<ڟa<<�a<Ѡa< �a<��a<�a<s�a<ܢa<F�a<��a<"�a<��a<�a<q�a<ƥa<%�a<��a<ͦa<_�a<��a<��a<L�a<��a<�a<8�a<��a<өa<H�a<x�a<˪a<�a<3�a<��a<��a<��a<$�a<w�a<��a<Ȭa<�a<�a<��a<w�a<ɭa<�a<�a<9�a<;�a<b�a<k�a<��a<��a<ˮa<�a<�a<�a<�a<-�a<"�a< �a<K�a<"�a<R�a<5�a<;�a<8�a<>�a<4�a<$�a<M�a<�a<6�a<�a<�a<�a<ˮa<��a<��a<��a<k�a<x�a<E�a<$�a<.�a<̭a<�a<��a<��a<j�a<,�a<�a<ͬa<��a<z�a<e�a<#�a<�a<Ыa<]�a<k�a<��a<Ԫa<��a<G�a<�a<��a<��a<-�a<	�a<��a<i�a<)�a<��a<��a<�a<٦a<p�a<$�a<¥a<m�a<'�a<��a<{�a<�a<��a<D�a<Ѣa<��a<�a<��a<?�a<ՠa<g�a<��a<��a<,�a<�a<U�a<�a<��a<�a<Ɯa<'�a<�a<S�a<�a<��a<�a<��a<J�a<�a<}�a<C�a<Ǘa<q�a<�a<��a<X�a<ڕa<��a<'�a<�a<��a</�a<��a<��a<y�a<��a<גa<��a<=�a<�a<��a<��a<;�a<�a<ܐa<��a<��a<V�a<V�a<�a<�a<Ώa<��a<��a<l�a<��a<W�a<P�a<E�a<F�a<>�a<4�a<g�a<?�a<u�a<Y�a<f�a<��a<��a<��a<�  �  ߏa<�a<�a<5�a<_�a<v�a<��a<ܐa<�a<<�a<m�a<��a<�a<C�a<��a<̒a<�a<U�a<��a<�a<U�a<��a<�a<F�a<��a<	�a<l�a<͖a<>�a<��a<
�a<n�a<ʘa<6�a<��a<�a<r�a<�a<`�a<ٛa<G�a<��a<.�a<��a<�a<��a<�a<L�a<şa<H�a<��a<�a<��a<	�a<y�a<�a<`�a<£a<+�a<��a<�a<Q�a<ƥa<�a<w�a<�a<T�a<��a<��a<Z�a<��a<��a<\�a<��a<�a<-�a<n�a<��a<�a<G�a<��a<֫a< �a<E�a<t�a<��a<Ӭa<�a<+�a<Z�a<��a<��a<ȭa<�a<�a<K�a<c�a<��a<��a<��a<��a<®a<ޮa<��a<	�a<�a<�a</�a<<�a<8�a<=�a<R�a<C�a<R�a<J�a<;�a<6�a<�a<�a<�a<�a<��a<��a<�a<Ǯa<îa<��a<�a<k�a<Q�a<!�a<�a<�a<ϭa<��a<m�a<U�a<>�a<�a<��a<��a<��a<I�a<
�a<ثa<��a<u�a<>�a<��a<תa<��a<R�a<�a<ݩa<��a<R�a<�a<��a<f�a<	�a<��a<o�a<+�a<ئa<��a<2�a<ӥa<��a<�a<��a<j�a<��a<��a</�a<ݢa<l�a<�a<��a<B�a<۠a<|�a<�a<��a<5�a<��a<N�a<�a<��a<
�a<��a<;�a<�a<h�a<�a<��a<4�a<əa<n�a<��a<��a<'�a<��a<V�a<�a<��a<Q�a< �a<��a<G�a<�a<��a<:�a<��a<��a<K�a< �a<ʒa<k�a<+�a<�a<ȑa<��a<a�a<�a<�a<��a<o�a<N�a<0�a<�a<�a<��a<��a<��a<��a<q�a<t�a<W�a<_�a<R�a<E�a<F�a<9�a<C�a<L�a<e�a<s�a<��a<��a<��a<�  �  Џa<؏a<+�a<�a<b�a<��a<��a<�a<��a<a�a<��a<đa< �a<�a<��a<��a<�a<Z�a<ϓa<��a<@�a<��a<�a<e�a<��a<�a<�a<��a<4�a<��a<�a<H�a<טa<8�a<��a<8�a<b�a<�a<L�a<��a<2�a<��a<�a<��a<�a<a�a<
�a<f�a<ߟa<^�a<��a<R�a<��a<�a<g�a<آa<J�a<��a<6�a<��a<(�a<J�a<ԥa<6�a<��a<�a<1�a<��a<��a<H�a<��a<�a<M�a<��a<��a<!�a<��a<Īa<�a<Y�a<j�a<Ыa<�a<;�a<\�a<��a<Ҭa<�a<K�a<\�a<��a<��a<ӭa<*�a< �a<M�a<C�a<��a<w�a<��a<ͮa<�a<
�a<ܮa</�a<�a<+�a<>�a<�a<Y�a<0�a<B�a<0�a<E�a<%�a<:�a<K�a<�a<S�a<�a<�a< �a<Үa<�a<��a<��a<��a<��a<N�a<U�a<9�a<�a<�a<��a<��a<��a<a�a<6�a<�a<�a<��a<��a<O�a<C�a<�a<��a<��a<;�a<�a<Ϫa<��a<e�a<��a<ҩa<v�a<K�a<�a<��a<h�a<�a<�a<_�a<>�a<Ŧa<s�a<�a<ƥa<q�a<�a<Ҥa<F�a<�a<��a<J�a<�a<Y�a<:�a<��a<P�a<ɠa<c�a<��a<��a<@�a<ʞa<��a<۝a<��a<(�a<��a<]�a<a<t�a<��a<��a<)�a<��a<_�a<ޘa<��a<�a<�a<j�a<�a<��a<-�a<��a<��a<>�a<єa<��a<:�a<�a<��a<N�a<#�a<��a<v�a<f�a<��a<ʑa<g�a<Q�a<��a<ݐa<��a<��a<z�a<�a<3�a<�a<׏a<ŏa<�a<��a<d�a<d�a<D�a<Q�a<.�a<D�a<[�a<-�a<}�a<C�a<o�a<v�a<k�a<��a<��a<�  �  ߏa<�a<�a<5�a<_�a<v�a<��a<ܐa<�a<<�a<m�a<��a<�a<C�a<��a<̒a<�a<U�a<��a<�a<U�a<��a<�a<F�a<��a<	�a<l�a<͖a<>�a<��a<
�a<n�a<ʘa<6�a<��a<�a<r�a<�a<`�a<ٛa<G�a<��a<.�a<��a<�a<��a<�a<L�a<şa<H�a<��a<�a<��a<	�a<y�a<�a<`�a<£a<+�a<��a<�a<Q�a<ƥa<�a<w�a<�a<T�a<��a<��a<Z�a<��a<��a<\�a<��a<�a<-�a<n�a<��a<�a<G�a<��a<֫a< �a<E�a<t�a<��a<Ӭa<�a<+�a<Z�a<��a<��a<ȭa<�a<�a<K�a<c�a<��a<��a<��a<��a<®a<ޮa<��a<	�a<�a<�a</�a<<�a<8�a<=�a<R�a<C�a<R�a<J�a<;�a<6�a<�a<�a<�a<�a<��a<��a<�a<Ǯa<îa<��a<�a<k�a<Q�a<!�a<�a<�a<ϭa<��a<m�a<U�a<>�a<�a<��a<��a<��a<I�a<
�a<ثa<��a<u�a<>�a<��a<תa<��a<R�a<�a<ݩa<��a<R�a<�a<��a<f�a<	�a<��a<o�a<+�a<ئa<��a<2�a<ӥa<��a<�a<��a<j�a<��a<��a</�a<ݢa<l�a<�a<��a<B�a<۠a<|�a<�a<��a<5�a<��a<N�a<�a<��a<
�a<��a<;�a<�a<h�a<�a<��a<4�a<əa<n�a<��a<��a<'�a<��a<V�a<�a<��a<Q�a< �a<��a<G�a<�a<��a<:�a<��a<��a<K�a< �a<ʒa<k�a<+�a<�a<ȑa<��a<a�a<�a<�a<��a<o�a<N�a<0�a<�a<�a<��a<��a<��a<��a<q�a<t�a<W�a<_�a<R�a<E�a<F�a<9�a<C�a<L�a<e�a<s�a<��a<��a<��a<�  �  ��a< �a<��a<C�a<S�a<z�a<Аa<��a<8�a<D�a<��a<̑a<��a<<�a<q�a<̒a<
�a<p�a<��a<��a<h�a<��a<�a<?�a<��a<�a<a�a<ۖa<�a<��a<�a<p�a<��a<9�a<��a<�a<��a<ؚa<`�a<��a<9�a<��a<�a<��a<�a<��a<ٞa<q�a<ڟa<<�a<Ѡa< �a<��a<�a<s�a<ܢa<F�a<��a<"�a<��a<�a<q�a<ƥa<%�a<��a<ͦa<_�a<��a<��a<L�a<��a<�a<8�a<��a<өa<H�a<x�a<˪a<�a<3�a<��a<��a<��a<$�a<w�a<��a<Ȭa<�a<�a<��a<w�a<ɭa<�a<�a<9�a<;�a<b�a<k�a<��a<��a<ˮa<�a<�a<�a<�a<-�a<"�a< �a<K�a<"�a<R�a<5�a<;�a<8�a<>�a<4�a<$�a<M�a<�a<6�a<�a<�a<�a<ˮa<��a<��a<��a<k�a<x�a<E�a<$�a<.�a<̭a<�a<��a<��a<j�a<,�a<�a<ͬa<��a<z�a<e�a<#�a<�a<Ыa<]�a<k�a<��a<Ԫa<��a<G�a<�a<��a<��a<-�a<	�a<��a<i�a<)�a<��a<��a<�a<٦a<p�a<$�a<¥a<m�a<'�a<��a<{�a<�a<��a<D�a<Ѣa<��a<�a<��a<?�a<ՠa<g�a<��a<��a<,�a<�a<U�a<�a<��a<�a<Ɯa<'�a<�a<S�a<�a<��a<�a<��a<J�a<�a<}�a<C�a<Ǘa<q�a<�a<��a<X�a<ڕa<��a<'�a<�a<��a</�a<��a<��a<y�a<��a<גa<��a<=�a<�a<��a<��a<;�a<�a<ܐa<��a<��a<V�a<V�a<�a<�a<Ώa<��a<��a<l�a<��a<W�a<P�a<E�a<F�a<>�a<4�a<g�a<?�a<u�a<Y�a<f�a<��a<��a<��a<�  �  ��a<��a<�a<0�a<_�a<��a<��a<ڐa<�a<?�a<��a<��a<�a<I�a<��a<֒a<�a<H�a<��a<�a<P�a<��a<�a<U�a<��a<�a<q�a<זa<#�a<��a<��a<`�a<՘a</�a<��a<�a<y�a<�a<m�a<śa<T�a<��a<�a<��a<�a<x�a<�a<h�a<ɟa<A�a<��a<$�a<��a< �a<��a<�a<\�a<ƣa< �a<��a<��a<V�a<åa<�a<��a<�a<E�a<��a<�a<S�a<��a<�a<H�a<��a<�a<+�a<p�a<��a<��a<N�a<��a<ūa<�a<6�a<x�a<��a<ڬa<�a<4�a<l�a<}�a<��a<ϭa<�a<�a<:�a<i�a<��a<��a<��a<��a<ݮa<�a<��a<�a<�a<+�a<0�a<3�a<;�a<U�a<1�a<W�a<O�a<5�a<R�a</�a<-�a<�a<�a<�a<�a<�a<�a<�a<��a<��a<��a<e�a<Q�a</�a<�a<�a<ͭa<��a<��a<K�a<8�a<�a<ެa<��a<}�a<<�a<'�a<ݫa<��a<n�a<L�a<�a<ժa<��a<X�a<�a<��a<��a<E�a<��a<��a<_�a<�a<��a<v�a<&�a<�a<x�a<?�a<ݥa<p�a<*�a<��a<]�a<��a<��a<4�a<֢a<n�a<�a<��a<9�a<�a<z�a<�a<��a<*�a<��a<Z�a<�a<��a<�a<��a<;�a<֛a<k�a<�a<��a<:�a<��a<Z�a<�a<��a<%�a<��a<`�a<��a<��a<M�a<�a<��a<8�a<�a<��a<A�a<��a<��a<]�a<��a<Œa<r�a<A�a<�a<��a<��a<O�a<�a<�a<��a<��a<T�a<3�a<�a<�a<׏a<��a<��a<��a<��a<S�a<k�a<[�a<>�a<\�a<?�a<G�a<C�a<W�a<]�a<��a<}�a<��a<͏a<�  �  ҏa<�a<�a<-�a<a�a<��a<��a<��a<	�a<V�a<��a<��a<�a<2�a<��a<��a<-�a<O�a<��a<��a<T�a<��a<�a<a�a<��a<�a<c�a<Ėa<2�a<��a<��a<O�a<јa<6�a<��a<�a<x�a<�a<N�a<Ǜa<6�a<��a<%�a<��a<�a<m�a< �a<[�a<˟a<]�a<��a<>�a<��a<�a<u�a<ڢa<M�a<��a<<�a<��a<�a<W�a<ץa<#�a<~�a<��a<5�a<��a<�a<Q�a<��a<�a<H�a<��a<�a<0�a<��a<ƪa<�a<M�a<t�a<ɫa<��a<9�a<j�a<��a<ڬa<��a<H�a<R�a<��a<��a<حa<�a<�a<^�a<T�a<{�a<��a<��a<��a<Үa<��a<�a<$�a<	�a<(�a<5�a<.�a<A�a<9�a<G�a<<�a<B�a<5�a<;�a<7�a<(�a<.�a<�a<�a<�a<�a<ޮa<��a<��a<��a<��a<b�a<S�a<6�a<��a<�a<��a<��a<��a<R�a<L�a<��a<�a<��a<��a<C�a<-�a<�a<��a<��a<0�a<�a<Ǫa<��a<I�a<�a<Щa<��a<H�a<�a<��a<f�a<�a<ԧa<u�a<,�a<Ʀa<y�a< �a<ǥa<y�a<�a<Ȥa<R�a<�a<��a<5�a<�a<j�a<&�a<��a<M�a<ؠa<e�a<�a<��a<F�a<��a<r�a<�a<��a<�a<��a<V�a<Ǜa<u�a<��a<��a<&�a<��a<Z�a<�a<��a<*�a<їa<l�a<�a<��a<7�a<�a<��a<<�a<��a<��a<A�a<�a<��a<C�a<�a<ϒa<{�a<P�a<�a<ۑa<x�a<K�a<
�a<�a<��a<�a<n�a<#�a<)�a<ߏa<ԏa<��a<��a<��a<m�a<h�a<P�a<O�a<>�a<E�a<G�a<B�a<X�a<R�a<e�a<w�a<x�a<��a<��a<�  �  ۏa<�a<�a<B�a<A�a<��a<��a<ސa<�a<O�a<��a<ɑa<��a</�a<��a<��a<�a<c�a<��a<��a<E�a<��a<�a<P�a<��a<�a<k�a<Ŗa<9�a<��a<��a<p�a<Řa<6�a<��a<�a<��a<�a<^�a<כa<@�a<��a<&�a<��a<�a<y�a<ߞa<f�a<ןa<<�a<��a<)�a<��a<�a<p�a<�a<]�a<��a<2�a<��a<��a<X�a<��a<*�a<��a<ަa<<�a<��a<��a<U�a<��a<��a<S�a<��a<�a<:�a<q�a<��a<�a<C�a<��a<ȫa<��a<>�a<o�a<��a<�a<��a<3�a<o�a<��a<��a<ԭa<��a<"�a<J�a<N�a<��a<��a<��a<ͮa<Ӯa<�a<�a<�a<!�a<(�a<�a<B�a<C�a<6�a<K�a<;�a<D�a<M�a<3�a<8�a<6�a<�a<!�a<�a<��a<��a<ݮa<��a<��a<��a<��a<x�a<3�a<2�a<�a<�a<ía<��a<��a<f�a<4�a<��a<��a<��a<��a<W�a<�a<�a<��a<}�a<P�a<�a<��a<��a<Q�a<	�a<ةa<{�a<D�a<	�a<��a<f�a<�a<��a<��a<)�a<֦a<��a<*�a<ͥa<z�a<�a<Ȥa<^�a<�a<��a<A�a<Ѣa<m�a<�a<��a<I�a<Ҡa<v�a<�a<��a<<�a<a<Z�a<�a<|�a<�a<��a<8�a<Λa<x�a<��a<��a<*�a<Ùa<e�a<��a<��a<4�a<��a<a�a<
�a<��a<U�a<�a<��a<@�a<�a<��a<L�a<ݓa<��a<`�a<	�a<��a<x�a<:�a<��a<Ǒa<r�a<]�a<�a<�a<��a<��a<b�a<*�a<
�a<��a<ӏa<��a<��a<��a<i�a<m�a<P�a<Q�a<V�a<=�a<H�a<Q�a<?�a<_�a<g�a<j�a<��a<��a<��a<�  �  ʏa<�a<�a<5�a<[�a<��a<��a<��a<)�a<H�a<��a<��a<��a<I�a<��a<͒a<
�a<]�a<��a<��a<\�a<��a<�a<L�a<��a<�a<l�a<ʖa<.�a<��a<�a<a�a<Øa<4�a<��a<�a<��a<�a<^�a<��a<L�a<��a<�a<��a<��a<��a<�a<f�a<Пa<C�a<Πa<�a<��a<��a<{�a<�a<V�a<��a<�a<��a<�a<t�a<ǥa<$�a<��a<�a<Q�a<��a< �a<M�a<��a<�a<<�a<��a<ܩa<6�a<�a<ƪa<�a<?�a<��a<��a<�a<6�a<n�a<��a<Ӭa<�a<.�a<k�a<��a<��a<�a<�a<#�a<7�a<d�a<��a<��a<��a<��a<خa<�a<�a<�a<�a<%�a<-�a<?�a<7�a<F�a<:�a<T�a<E�a<7�a<:�a</�a<2�a<&�a<!�a<�a<��a<�a<ٮa<ڮa<��a<��a<�a<k�a<M�a<.�a<�a<�a<�a<��a<��a<Z�a<0�a<�a<�a<��a<z�a<Q�a<�a<�a<īa<v�a<M�a<�a<٪a<��a<R�a<�a<ͩa<��a<8�a<��a<��a<d�a< �a<Χa<}�a<�a<֦a<p�a<6�a<٥a<l�a<#�a<��a<k�a<��a<��a<:�a<آa<��a<�a<��a<9�a<ݠa<t�a<�a<��a<(�a<ʞa<L�a<�a<��a<�a<��a<:�a<�a<c�a<�a<��a<1�a<ؙa<N�a<��a<��a<0�a<͗a<m�a<	�a<��a<K�a<��a<��a<9�a<�a<��a<:�a<��a<��a<\�a<�a<ϒa<��a<.�a<��a<��a<��a<Q�a<�a<��a<��a<��a<T�a<L�a<�a<�a<Џa<��a<��a<��a<z�a<\�a<i�a<Q�a<@�a<D�a<?�a<M�a<Q�a<`�a<_�a<p�a<�a<��a<Əa<�  �  ˏa<��a<�a<�a<k�a<��a<��a<�a<�a<N�a<��a<��a< �a<E�a<u�a<ђa<�a<V�a<��a<��a<H�a<��a<�a<Z�a<��a<�a<n�a<Җa<&�a<��a<�a<\�a<Әa<5�a<��a<�a<m�a<��a<Z�a<ʛa<8�a<��a<"�a<��a<�a<l�a<��a<^�a<ӟa<G�a<��a<-�a<��a<�a<{�a<ݢa<I�a<ģa<%�a<��a< �a<Z�a<��a<)�a<��a<��a<:�a<��a<�a<T�a<��a<��a<I�a<��a<�a<$�a<��a<Ūa<�a<N�a<��a<ȫa<��a<0�a<t�a<��a<Ƭa<	�a<@�a<\�a<��a<��a<ݭa<
�a<"�a<D�a<h�a<r�a<��a<��a<��a<�a<�a<�a<�a<�a<'�a<?�a< �a<;�a<L�a<B�a<;�a<>�a<>�a<B�a<7�a<�a<<�a<�a<�a<�a<�a<ݮa<��a<��a<��a<��a<P�a<]�a<5�a<�a<��a<��a<��a<��a<T�a<7�a<�a<Ѭa<��a<��a<J�a<,�a<�a<��a<��a<<�a<�a<תa<y�a<U�a<�a<ũa<~�a<I�a<��a<��a<d�a<�a<٧a<j�a<1�a<Ҧa<}�a<"�a<ȥa<v�a<'�a<��a<Q�a<�a<��a<=�a<ܢa<m�a<�a<��a<=�a<ݠa<i�a<��a<��a</�a<͞a<c�a<�a<��a<�a<��a<N�a<̛a<d�a<
�a<��a<%�a<��a<[�a<�a<��a<�a<֗a<k�a<�a<��a<E�a<�a<��a<3�a<�a<��a<-�a<�a<��a<N�a<�a<��a<��a<G�a<��a<��a<��a<B�a<�a<�a<��a<��a<^�a<'�a<�a<�a<ӏa<ŏa<��a<��a<��a<d�a<P�a<J�a<G�a<L�a<G�a<3�a<f�a<D�a<c�a<|�a<��a<��a<��a<�  �  �a<؏a<�a<7�a<V�a<��a<��a<�a<�a<P�a<w�a<őa<��a<<�a<��a<a<�a<X�a<��a<��a<F�a<��a<�a<Y�a<��a<�a<k�a<��a<H�a<��a<�a<X�a<˘a<@�a<��a<�a<q�a<�a<L�a<�a<9�a<��a<)�a<��a<�a<m�a<�a<R�a<Οa<C�a<��a<+�a<��a<�a<v�a<�a<Y�a<��a<.�a<~�a<��a<U�a<��a<%�a<z�a<�a<5�a<��a<�a<P�a<��a<��a<a�a<��a<��a<)�a<x�a<��a<�a<O�a<|�a<٫a<�a<S�a<f�a<��a<�a<��a<@�a<Z�a<��a<��a<խa<��a<�a<F�a<Y�a<��a<��a<��a<ʮa<Ȯa<�a<��a<�a<�a< �a<-�a<3�a<H�a<)�a<X�a<E�a<C�a<L�a<-�a<P�a<�a<&�a<�a<%�a<�a<�a<�a<��a<ʮa<��a<��a<m�a<H�a<0�a<�a<��a<ĭa<��a<w�a<b�a<6�a<�a<�a<��a<��a<M�a<�a<�a<��a<��a<=�a<�a<Ūa<��a<Q�a<�a<�a<w�a<U�a<�a<��a<p�a<�a<ȧa<n�a<C�a<Ŧa<��a<#�a<ޥa<}�a<�a<Фa<R�a<�a<��a<8�a<آa<i�a<�a<��a<G�a<ؠa<v�a<�a<��a<8�a<��a<[�a<�a<�a<�a<��a<I�a<ƛa<�a<��a<��a<@�a<��a<s�a<�a<��a<#�a<Ɨa<[�a<	�a<��a<?�a<�a<��a<V�a<ܔa<��a<N�a<�a<��a<K�a<�a<��a<x�a<5�a<�a<Ña<}�a<W�a<�a<�a<��a<v�a<a�a<,�a<�a<�a<̏a<��a<��a<��a<]�a<z�a<Y�a<O�a<U�a<7�a<`�a<:�a<P�a<J�a<}�a<f�a<��a<��a<��a<�  �  ďa<��a<�a<8�a<X�a<��a<a<ϐa<2�a<R�a<~�a<ӑa<��a<>�a<x�a<Ȓa<�a<r�a<��a<
�a<_�a<��a<�a<R�a<��a<�a<t�a<ǖa<*�a<��a<�a<c�a<��a<;�a<��a<�a<��a<�a<L�a<Лa<1�a<��a<�a<��a<�a<~�a<�a<k�a<ٟa<E�a<Ԡa<(�a<��a<�a<o�a<ۢa<F�a<��a<(�a<��a<��a<z�a<ͥa<+�a<��a<�a<F�a<��a<�a<B�a<��a<�a<L�a<��a<ߩa<;�a<��a<ʪa<�a<>�a<��a<��a<��a<5�a<h�a<��a<֬a<�a<5�a<u�a<��a<ĭa<�a<��a<4�a<@�a<^�a<r�a<��a<��a<Үa<֮a<�a<�a<��a<&�a<*�a<.�a<<�a<>�a<E�a<4�a<F�a<5�a<J�a<&�a<3�a<;�a<!�a<$�a<�a<�a<��a<ˮa<Ȯa<��a<��a<��a<m�a<J�a<1�a<!�a<ܭa<�a<��a<~�a<p�a</�a<	�a<Ԭa<��a<~�a<g�a<�a<��a<ƫa<p�a<Z�a<
�a<̪a<��a<Z�a<�a<ɩa<��a<;�a<��a<��a<j�a< �a<Чa<��a<�a<Ħa<��a<�a<ѥa<e�a<#�a<��a<c�a<�a<��a<C�a<ڢa<��a<�a<��a<G�a<Ҡa<g�a<��a<��a<2�a<Ҟa<Y�a<�a<��a<�a<��a<B�a<כa<e�a<�a<��a<.�a<��a<^�a<�a<��a<5�a<ӗa<p�a<�a<��a<H�a<�a<��a<8�a<ޔa<��a<=�a<�a<��a<f�a<�a<Ғa<��a<4�a<�a<��a<��a<B�a<�a<ސa<��a<��a<`�a<S�a<�a<��a<֏a<��a<��a<��a<y�a<V�a<[�a<A�a<S�a<0�a<C�a<U�a<L�a<c�a<f�a<^�a<��a<��a<��a<�  �  ��a<�a< �a</�a<f�a<p�a<Őa<Ґa<�a<9�a<��a<��a<��a<Z�a<t�a<�a<��a<X�a<��a<�a<D�a<��a<
�a<8�a<ŕa<��a<m�a<ۖa<�a<��a<�a<s�a<Θa</�a<��a<��a<}�a<�a<t�a<̛a<G�a<��a<�a<��a<�a<��a<۞a<\�a<֟a<1�a<��a<�a<��a<�a<��a<�a<S�a<Уa<�a<��a<�a<X�a<��a<#�a<��a<Цa<]�a<��a<�a<K�a<��a<	�a<H�a<��a<�a<1�a<m�a<��a< �a<G�a<��a<��a<�a<+�a<y�a<��a<Ƭa<"�a<�a<q�a<��a<��a<֭a<�a<#�a</�a<}�a<p�a<��a<��a<��a<�a<׮a<��a<��a<+�a<�a<.�a<7�a<+�a<f�a<�a<a�a<@�a<F�a<L�a<,�a<0�a<�a<�a<�a<�a<��a<Ԯa<�a<��a<��a<t�a<e�a<Y�a<�a<#�a<߭a<ɭa<��a<��a<N�a<-�a<&�a<Ьa<Ϭa<o�a<L�a<�a<�a<��a<r�a<V�a<�a<�a<��a<T�a<�a<��a<��a<<�a<�a<��a<_�a<�a<��a<z�a<!�a<�a<~�a<1�a<�a<e�a<>�a<��a<q�a<�a<��a<A�a<Ţa<o�a<��a<��a<,�a<�a<x�a<�a<��a<�a<Ӟa<G�a<�a<s�a<�a<��a<*�a<�a<O�a<�a<��a<5�a<ԙa<Z�a<�a<��a<,�a<��a<`�a<�a<��a<_�a<�a<��a<.�a<�a<��a<-�a<�a<��a<b�a< �a<��a<y�a</�a<��a<��a<��a<@�a<+�a<�a<��a<��a<G�a<1�a<��a<�a<Ïa<��a<��a<u�a<��a<A�a<v�a<M�a<O�a<V�a<<�a<K�a<;�a<V�a<[�a<��a<��a<��a<Տa<�  �  Ǐa<�a< �a<9�a<\�a<��a<��a<��a<�a<[�a<��a<��a<��a<4�a<x�a<��a<�a<]�a<��a<
�a<N�a<��a<��a<P�a<��a<�a<V�a<��a</�a<��a<�a<M�a<Ęa<;�a<��a<!�a<�a<��a<P�a<��a<+�a<��a<�a<��a<��a<��a<�a<a�a<؟a<O�a<��a<8�a<��a<�a<t�a<Ԣa<D�a<��a<*�a<��a<	�a<a�a<˥a<-�a<��a<�a<U�a<��a<�a<C�a<��a<�a<=�a<��a<�a<6�a<��a<̪a<�a<F�a<u�a<��a<��a<=�a<c�a<��a<׬a<�a<5�a<d�a<��a<��a<�a<�a<$�a<E�a<S�a<q�a<��a<��a<®a<�a<��a<��a<�a<�a<%�a<-�a<>�a</�a<9�a<;�a<K�a<1�a<,�a<4�a<A�a<1�a<=�a<�a<�a<��a<׮a<ʮa<ˮa<��a<��a<t�a<o�a<N�a<-�a<�a<�a<έa<��a<��a<[�a<6�a<��a<Ԭa<��a<��a<Q�a<)�a<��a<��a<��a<D�a<�a<֪a<��a<=�a<�a<ͩa<��a<5�a<�a<��a<k�a<!�a<ܧa<|�a<0�a<Ȧa<o�a<�a<եa<k�a<�a<��a<p�a<��a<��a<B�a<�a<u�a< �a<��a<A�a<֠a<`�a<��a<��a<4�a<˞a<l�a<�a<��a<�a<��a<>�a<�a<c�a<�a<��a<0�a<��a<P�a<�a<��a<1�a<ٗa<r�a<�a<��a<8�a<�a<��a<@�a<ؔa<{�a<>�a<��a<��a<U�a<�a<ƒa<��a<H�a<��a<a<w�a<A�a<�a<�a<��a<��a<l�a<7�a<#�a<�a<яa<��a<��a<z�a<m�a<]�a<`�a<=�a<4�a<>�a<Q�a<K�a<g�a<[�a<n�a<k�a<o�a<��a<��a<�  �  �a<�a<E�a<r�a<n�a<ʐa<ΐa<�a</�a<z�a<��a<��a<?�a<U�a<��a<�a<M�a<��a<˓a<$�a<e�a<Δa<�a<��a<��a<N�a<��a<�a<p�a<��a<7�a<��a<��a<^�a<��a<:�a<��a<"�a<t�a<�a<k�a<ޜa<S�a<��a<<�a<��a<�a<��a<�a<d�a<ʠa<E�a<��a<=�a<��a<��a<i�a<ݣa<[�a<��a<�a<p�a<ޥa<A�a<��a<�a<L�a<ѧa<
�a<y�a<بa<�a<��a<��a<�a<@�a<��a<֪a<�a<r�a<��a<��a<�a<m�a<��a<ìa<�a<�a<p�a<r�a<��a<ŭa<�a<�a<>�a<r�a<t�a<��a<��a<�a<��a<�a<�a<	�a<'�a<*�a<Y�a<=�a<_�a<h�a<L�a<}�a<U�a<y�a<t�a<Q�a<b�a<@�a<O�a<(�a<6�a<�a<�a<�a<Ԯa<�a<��a<��a<��a<V�a<j�a<!�a<�a<ܭa<έa<��a<��a<k�a<�a<�a<Ŭa<��a<y�a<6�a<�a<īa<��a<T�a<I�a<ͪa<˪a<z�a<�a<�a<��a<x�a<�a<٨a<��a<*�a<�a<��a<X�a<�a<��a<Q�a<��a<��a<&�a<�a<p�a<"�a<ȣa<T�a<��a<��a<,�a<��a<v�a<�a<��a<�a<��a<g�a<ݞa<|�a<�a<��a<7�a<Мa<r�a<�a<��a<�a<Śa<e�a<�a<��a<�a<Ęa<C�a<�a<��a<)�a<ۖa<n�a<.�a<��a<y�a<�a<��a<��a<��a<�a<n�a<4�a<ݒa<��a<_�a<#�a<��a<��a<h�a<+�a<!�a<�a<��a<��a<L�a<6�a<�a<�a<Ώa<яa<��a<��a<��a<u�a<��a<��a<f�a<}�a<f�a<��a<r�a<��a<��a<��a<ݏa<ʏa<�  �  ��a<�a<9�a<f�a<��a<��a<ܐa<�a<D�a<w�a<��a<ߑa<�a<u�a<��a<�a<*�a<��a<דa<-�a<��a<ܔa<�a<��a<Օa<6�a<��a<��a<U�a<��a<�a<��a<�a<g�a<ҙa<=�a<��a<�a<{�a<�a<Z�a<Μa<C�a<��a<+�a<��a<�a<��a<��a<z�a<�a<K�a<ša<�a<��a<�a<|�a<�a<9�a<��a<�a<��a<��a<P�a<��a<�a<i�a<��a<�a<m�a<��a<�a<b�a<��a<
�a<T�a<��a<�a<,�a<h�a<��a<ګa<�a<R�a<��a<Ĭa<��a<%�a<W�a<z�a<��a<�a<�a<!�a<C�a<P�a<��a<��a<®a<Ůa<Ԯa<�a<�a<#�a<8�a<;�a<I�a<I�a<`�a<[�a<f�a<_�a<`�a<`�a<V�a<W�a<X�a<L�a<E�a<<�a<2�a<�a<�a<��a<�a<Юa<��a<��a<��a<h�a<T�a</�a<�a<�a<ʭa<��a<r�a<I�a<7�a<�a<�a<��a<r�a<A�a<�a<߫a<��a<]�a</�a<�a<��a<r�a<6�a<�a<��a<[�a<�a<Шa<��a<C�a<�a<��a<K�a<�a<��a<@�a<�a<��a<>�a<ޤa<��a< �a<ģa<e�a<�a<��a<2�a<աa<Q�a<��a<��a<2�a<��a<E�a<�a<��a<#�a<��a<F�a<ќa<e�a< �a<��a<)�a<��a<M�a<�a<{�a<�a<��a<V�a<��a<��a<6�a<іa<k�a<�a<��a<^�a<�a<��a<i�a<�a<˓a<u�a<C�a<��a<��a<h�a<(�a<ؑa<��a<�a<M�a<�a<ΐa<��a<��a<f�a<H�a<�a< �a<ۏa<ҏa<��a<��a<��a<��a<w�a<j�a<l�a<s�a<r�a<{�a<��a<��a<��a<��a<��a<܏a<�  �  ߏa<9�a<.�a<[�a<��a<��a<�a<�a<G�a<[�a<��a<�a<�a<��a<��a<�a<*�a<��a<ϓa<�a<u�a<Ôa<*�a<j�a<�a<'�a<��a<�a<D�a<ڗa<�a<��a<�a<X�a<Ιa<+�a<��a< �a<��a<�a<s�a<�a<?�a<ѝa<�a<��a<�a<��a<�a<X�a<ܠa<-�a<ҡa<�a<��a<�a<m�a<�a<7�a<ɤa< �a<��a<եa<A�a<��a<��a<{�a<��a<1�a<s�a<Ϩa</�a<e�a<ͩa<��a<W�a<��a<�a<#�a<]�a<��a<ګa<9�a<L�a<��a<άa<�a<@�a<C�a<��a<��a<ͭa<�a<�a<T�a<L�a<��a<��a<Ǯa<ɮa<߮a<�a<�a<%�a<�a<=�a<;�a<S�a<\�a<K�a<��a<K�a<��a<f�a<f�a<l�a<D�a<X�a<:�a<C�a<�a<(�a<�a<��a<
�a<��a<ܮa<��a<��a<y�a<B�a<6�a<�a<��a<��a<��a<~�a<J�a<B�a<�a<�a<��a<��a<:�a<��a<ӫa<��a<l�a<�a<�a<��a<s�a<K�a<کa<ȩa<\�a</�a<Ψa<��a<>�a<�a<��a<7�a<�a<��a<X�a< �a<��a<S�a<Ĥa<��a<�a<��a<\�a<�a<��a<�a<�a<U�a<
�a<��a<$�a<џa<C�a<�a<f�a<�a<��a<7�a<Ԝa<U�a<�a<x�a<>�a<��a<\�a<�a<�a<0�a<��a<Y�a<�a<��a<-�a<ǖa<��a<�a<וa<X�a<!�a<Ĕa<V�a<0�a<��a<��a<-�a<�a<��a<X�a<9�a<ԑa<a<]�a<R�a<	�a<ِa<Őa<j�a<h�a<-�a<�a<�a<�a<Ώa<��a<��a<x�a<��a<}�a<z�a<��a<_�a<~�a<o�a<��a<��a<��a<��a<Ïa<�a<�  �  �a<�a<;�a<d�a<}�a<��a<�a<�a<V�a<w�a<��a<�a<(�a<k�a<��a<��a<;�a<��a<ʓa</�a<��a<Ɣa<-�a<x�a<ѕa<;�a<��a<�a<R�a<��a<�a<��a<�a<^�a<͙a<6�a<��a<�a<�a<�a<W�a<؜a<<�a<��a<+�a<��a<�a<��a<��a<c�a<�a<F�a<��a<2�a<��a< �a<k�a<�a<M�a<��a<�a<��a<ߥa<G�a<��a<�a<i�a<��a<�a<g�a<Ǩa<�a<f�a<��a<�a<Y�a<��a<�a<'�a<a�a<��a<۫a<�a<V�a<��a<Ƭa<��a<$�a<S�a<��a<��a<حa<�a<�a<F�a<a�a<��a<��a<��a<Ϯa<�a<�a<
�a<4�a<%�a<B�a<B�a<H�a<\�a<[�a<d�a<[�a<g�a<V�a<g�a<T�a<R�a<X�a<H�a<@�a<'�a<�a<�a<�a<�a<ʮa<��a<��a<��a<e�a<L�a<:�a<�a<�a<˭a<��a<��a<U�a<-�a<�a<֬a<��a<z�a<5�a<�a<�a<��a<p�a<'�a<�a<��a<u�a<*�a<�a<��a<X�a<�a<˨a<��a<=�a<�a<��a<G�a<�a<��a<=�a<��a<��a<=�a<ޤa<��a<�a<ţa<c�a<��a<��a<-�a<ǡa<l�a<�a<��a<"�a<ȟa<Y�a<�a<{�a<#�a<��a<=�a<לa<d�a< �a<��a<*�a<��a<U�a<��a<��a<�a<��a<\�a<�a<��a<1�a<ʖa<v�a<�a<��a<b�a<�a<��a<k�a<�a<Ɠa<��a<2�a<�a<��a<]�a<+�a<�a<��a<c�a<>�a<�a<�a<��a<��a<w�a<4�a<#�a<��a<ُa<͏a<��a<��a<��a<��a<m�a<{�a<i�a<m�a<~�a<}�a<��a<��a<��a<��a<��a<�a<�  �  �a<
�a<?�a<a�a<�a<��a<ڐa<�a<+�a<�a<��a<�a<�a<g�a<ʒa<�a<9�a<|�a<ԓa<'�a<l�a<Дa<�a<��a<͕a<=�a<��a<�a<t�a<��a<1�a<��a<�a<c�a<ęa<7�a<��a<#�a<r�a< �a<W�a<ܜa<R�a<��a<<�a<��a<�a<��a<��a<g�a<ɠa<Z�a<��a<.�a<��a<�a<��a<ңa<N�a<��a<&�a<s�a<�a<H�a<��a<�a<Z�a<ѧa<�a<w�a<Өa<
�a<{�a<��a<�a<F�a<��a<ݪa<&�a<k�a<��a<��a<�a<q�a<��a<��a<�a<�a<g�a<u�a<��a<˭a<��a<#�a<4�a<a�a<y�a<��a<��a<îa<�a<�a<�a<�a<-�a<:�a<I�a<O�a<T�a<f�a<S�a<y�a<a�a<c�a<e�a<M�a<h�a<9�a<E�a<*�a<;�a<�a<�a<�a<�a<�a<��a<��a<��a<g�a<W�a<.�a<�a<حa<ӭa<��a<w�a<L�a<(�a<�a<ͬa<��a<g�a<?�a<�a<˫a<��a<[�a<;�a<�a<��a<s�a<'�a<�a<��a<r�a<�a<Шa<��a<5�a<�a<��a<Z�a<�a<��a<<�a<��a<��a</�a<�a<v�a<-�a<��a<_�a<��a<��a<B�a<��a<g�a<�a<��a<;�a<��a<Z�a<ߞa<��a<�a<��a<?�a<Ȝa<u�a<�a<��a<�a<Úa<`�a<ܙa<��a<�a<Ƙa<H�a<�a<��a<0�a<Ֆa<f�a<'�a<��a<~�a<�a<��a<t�a<
�a<ۓa<p�a<8�a<�a<��a<j�a<�a<�a<��a<��a<B�a<�a<ܐa<��a<��a<H�a<=�a<�a< �a<�a<Əa<��a<��a<��a<��a<z�a<y�a<c�a<��a<_�a<{�a<s�a<��a<��a<��a<͏a<ڏa<�  �  �a<�a<>�a<Y�a<��a<��a<֐a<�a<9�a<z�a<��a<�a<1�a<b�a<��a<�a<B�a<��a<��a<"�a<t�a<ؔa<�a<|�a<��a<,�a<��a<��a<K�a<��a<'�a<��a<��a<T�a<��a<<�a<��a<�a<�a<��a<a�a<͜a<?�a<��a<)�a<��a<�a<��a<��a<o�a<ՠa<N�a<¡a<,�a<��a<��a<h�a<ݣa<K�a<��a<�a<}�a<�a<L�a<��a<�a<c�a<��a<�a<n�a<��a<�a<r�a<��a<
�a<E�a<��a<ܪa<�a<l�a<��a<�a<�a<K�a<��a<ˬa<�a<+�a<V�a<~�a<��a<ӭa<��a<(�a<G�a<d�a<x�a<��a<��a<׮a<�a<�a<�a<�a<5�a<4�a<E�a<X�a<U�a<_�a<e�a<W�a<\�a<h�a<e�a<_�a<\�a<B�a<W�a<-�a<+�a<#�a<�a<�a<ݮa<Ůa<��a<��a<��a<w�a<O�a<)�a<�a<�a<έa<��a<��a<^�a<#�a<�a<ʬa<��a<y�a<K�a<	�a<ҫa<��a<`�a<+�a<��a<��a<|�a<3�a<�a<��a<h�a<!�a<٨a<}�a<1�a<�a<��a<K�a<�a<��a<F�a<�a<��a<<�a<ܤa<�a<(�a<£a<a�a<�a<��a<5�a<ҡa<e�a<��a<��a<�a<��a<X�a<�a<��a<�a<��a<C�a<ќa<k�a<��a<��a<&�a<��a<K�a<�a<��a<�a<��a<G�a<�a<��a<'�a<Ֆa<x�a<�a<��a<X�a<�a<��a<_�a<�a<ʓa<z�a<=�a<�a<��a<o�a<,�a<�a<��a<c�a<8�a<�a<ߐa<��a<��a<X�a<E�a<�a<��a<�a<Əa<��a<��a<��a<|�a<��a<x�a<t�a<w�a<h�a<��a<w�a<��a<��a<��a<͏a<ԏa<�  �  �a<"�a<4�a<a�a<��a<��a<�a<�a<N�a<n�a<��a<�a<*�a<p�a<��a<��a<:�a<��a<̓a<'�a<��a<Ôa<3�a<o�a<�a<.�a<��a<��a<O�a<ϗa<�a<��a<�a<d�a<˙a<3�a<��a<�a<��a<�a<k�a<՜a<>�a<ɝa<�a<��a<�a<��a<��a<b�a<�a<=�a<��a<"�a<��a<�a<s�a<�a<B�a<��a<�a<��a<ߥa<B�a<��a<��a<q�a<��a<'�a<k�a<èa<'�a<_�a<��a<�a<a�a<��a<�a<-�a<_�a<��a<իa<3�a<Q�a<��a<̬a<�a<5�a<H�a<��a<��a<حa< �a<�a<B�a<]�a<��a<��a<��a<ծa<�a<��a< �a</�a<#�a<?�a<J�a<I�a<^�a<Q�a<n�a<Y�a<n�a<b�a<W�a<Z�a<T�a<V�a<B�a<?�a<,�a<�a<�a<��a<�a<Ǯa<Ʈa<��a<��a<m�a<O�a<:�a<�a<��a<­a<��a<{�a<W�a<1�a<��a<ܬa<��a<q�a<6�a<�a<߫a<��a<v�a<�a<��a<��a<y�a<5�a<�a<��a<U�a<�a<Ψa<��a<<�a<�a<��a<C�a<��a<��a<P�a<�a<��a<L�a<Ѥa<��a<�a<ʣa<^�a<��a<��a<$�a<ϡa<\�a<�a<��a<)�a<ϟa<O�a<�a<t�a<%�a<��a<8�a<ޜa<[�a<�a<��a<4�a<��a<P�a<��a<y�a<#�a<��a<d�a<�a<��a<7�a<ɖa<u�a<�a<Еa<^�a<�a<a<]�a<%�a<��a<��a<,�a<�a<��a<\�a<'�a<�a<��a<t�a<F�a<�a<ܐa<��a<{�a<r�a<3�a< �a<�a<ۏa<Ϗa<��a<��a<��a<��a<y�a<k�a<o�a<o�a<|�a<x�a<��a<��a<��a<��a<��a<�a<�  �  �a<�a<8�a<i�a<�a<��a<�a< �a<6�a<~�a<��a<�a<$�a<_�a<��a<�a<C�a<��a<ۓa<)�a<q�a<��a<&�a<~�a<֕a<?�a<��a<�a<_�a<��a<'�a<��a<�a<d�a<��a<#�a<��a<�a<��a<��a<`�a<՜a<N�a<��a<.�a<��a<	�a<��a<��a<]�a<Ѡa<Q�a<��a<0�a<��a<�a<u�a<ԣa<M�a<��a<!�a<x�a<ۥa<E�a<��a<�a<c�a<ŧa<�a<v�a<˨a<�a<o�a<��a<�a<M�a<��a<تa<(�a<g�a<��a<�a<�a<`�a<��a<Ŭa<��a<&�a<T�a<��a<��a<έa<��a<&�a<@�a<f�a<s�a<��a<��a<Ʈa<�a<�a<�a<�a< �a<<�a<O�a<F�a<`�a<[�a<Z�a<q�a<_�a<`�a<k�a<b�a<]�a<G�a<2�a<1�a<3�a< �a<�a<��a<�a<߮a<��a<��a<��a<f�a<V�a<6�a<�a<�a<ҭa<��a<��a<P�a< �a<�a<Ƭa<��a<t�a<F�a<�a<ϫa<��a<i�a<-�a<�a<��a<s�a<.�a<��a<��a<h�a<#�a<Ҩa<��a<0�a<اa<��a<J�a<��a<��a<E�a<�a<��a<7�a<�a<��a<�a<ţa<^�a<�a<��a<8�a<ѡa<i�a<��a<��a<+�a<��a<Y�a<�a<��a<�a<��a<;�a<Ҝa<a�a<��a<��a<$�a<a<X�a<�a<��a<%�a<��a<O�a<�a<��a<2�a<Жa<y�a<�a<��a<l�a<�a<��a<p�a<�a<ȓa<��a<,�a<�a<��a<m�a<%�a<�a<��a<��a<8�a<�a<�a<��a<��a<T�a<0�a<�a<�a<؏a<ҏa<��a<��a<��a<�a<x�a<�a<w�a<x�a<l�a<g�a<{�a<��a<��a<��a<Ǐa<؏a<�  �  ��a<�a<D�a<V�a<��a<��a<Аa<'�a<<�a<��a<��a<�a<5�a<^�a<��a<ޒa<O�a<y�a<ޓa<"�a<w�a<��a<�a<��a<ӕa<9�a<��a<��a<X�a<��a<0�a<�a<�a<P�a<̙a<O�a<��a<�a<s�a<��a<^�a<˜a<I�a<��a<>�a<��a<�a<�a<�a<~�a<͠a<[�a<��a<2�a<��a<�a<s�a<أa<V�a<��a<,�a<p�a<��a<J�a<��a<�a<X�a<Чa<�a<r�a<��a<�a<u�a<��a<
�a<F�a<��a<�a<�a<g�a<��a<��a<�a<X�a<��a<Ĭa<�a<�a<e�a<u�a<��a<٭a<�a<,�a<2�a<s�a<m�a<��a<��a<׮a<�a<�a<�a<�a<I�a</�a<H�a<V�a<M�a<j�a<W�a<g�a<V�a<g�a<]�a<Q�a<P�a<I�a<`�a<6�a<#�a<�a<�a<�a<ծa<֮a<��a<��a<��a<r�a<U�a<$�a<*�a<�a<ԭa<��a<v�a<a�a< �a<�a<��a<��a<c�a<H�a<	�a<իa<��a<Y�a<8�a<�a<��a<t�a<3�a<�a<��a<q�a<�a<Шa<y�a<=�a<�a<��a<I�a<�a<��a<D�a<�a<��a<-�a<�a<s�a<.�a<��a<[�a<�a<��a<B�a<��a<l�a<��a<��a<)�a<��a<b�a<۞a<��a<�a<��a<A�a<ǜa<w�a<�a<��a<�a<��a<N�a<�a<��a<�a<��a<I�a<�a<��a< �a<іa<g�a<(�a<��a<e�a<�a<��a<q�a<�a<ٓa<q�a<B�a<�a<��a<s�a<�a<��a<��a<y�a<<�a<�a<ܐa<��a<��a<Y�a<Y�a<�a<��a<�a<��a<��a<��a<��a<v�a<~�a<q�a<f�a<k�a<o�a<��a<�a<��a<��a<��a<̏a<̏a<�  �  �a<"�a<5�a<V�a<��a<��a<ސa<�a<D�a<g�a<��a<�a<&�a<p�a<��a<��a<9�a<��a<ۓa<�a<{�a<Ĕa<&�a<z�a<ܕa<.�a<��a<��a<Q�a<җa<�a<��a<��a<^�a<řa<#�a<��a<�a<��a<�a<p�a<՜a<E�a<��a<)�a<��a<�a<��a<�a<f�a<Ԡa<C�a<��a<&�a<��a<�a<s�a<�a<F�a<��a<�a<v�a<�a<<�a<��a<�a<g�a<��a< �a<p�a<¨a<'�a<e�a<��a<	�a<Y�a<��a<ڪa<)�a<p�a<��a<߫a<1�a<S�a<��a<Ǭa<�a<,�a<U�a<��a<��a<حa<�a<�a<=�a<`�a<��a<��a<��a<Ϯa<�a<��a< �a<�a<'�a<5�a<H�a<V�a<O�a<X�a<l�a<\�a<q�a<k�a<T�a<d�a<U�a<R�a<+�a<<�a<+�a<%�a<�a<��a<��a<ʮa<Ʈa<��a<��a<t�a<Q�a<2�a<	�a<�a<��a<��a<x�a<R�a<2�a<�a<ݬa<��a<k�a<E�a< �a<٫a<��a<i�a<)�a<��a<��a<p�a<9�a<�a<��a<_�a<�a<ܨa<��a<5�a<اa<��a<I�a<��a<��a<V�a<�a<��a<B�a<ܤa<�a<"�a<ãa<U�a<��a<��a<*�a<ϡa<_�a< �a<��a<*�a<ǟa<R�a<�a<{�a<�a<��a<2�a<՜a<g�a<��a<��a<-�a<��a<O�a<��a<~�a<�a<��a<[�a<�a<��a<3�a<ٖa<m�a<�a<ϕa<`�a<�a<��a<c�a<�a<ɓa<��a<)�a<�a<��a<f�a<"�a<�a<��a<x�a<F�a<�a<ڐa<��a<{�a<b�a<6�a<�a<��a<�a<��a<��a<��a<��a<��a<��a<h�a<y�a<p�a<x�a<a�a<��a<��a<��a<��a<ɏa<�a<�  �  �a<�a<*�a<n�a<��a<��a<��a<�a<d�a<s�a<��a<�a<�a<t�a<��a<��a<*�a<��a<ۓa<,�a<��a<��a<@�a<i�a<�a<4�a<��a<��a<G�a<ėa<�a<��a<�a<\�a<֙a< �a<��a<��a<��a<��a<]�a<˜a<@�a<��a<�a<��a<��a<��a<�a<`�a<�a<A�a<Сa<�a<��a<�a<m�a<�a<;�a<Ǥa<�a<��a<�a<N�a<��a<�a<|�a<��a<�a<j�a<��a<�a<S�a<ϩa<�a<b�a<��a<�a<-�a<X�a<��a<ūa<$�a<G�a<��a<¬a<�a<8�a<=�a<��a<��a<�a<�a<!�a<S�a<O�a<��a<��a<��a<Ȯa<�a<�a<�a<=�a<�a<V�a<C�a<E�a<m�a<K�a<h�a<[�a<e�a<Q�a<_�a<j�a<D�a<i�a<&�a<R�a<�a<"�a<�a<�a<�a<Ǯa<��a<��a<��a<g�a<G�a<Q�a<��a<�a<ǭa<��a<��a<I�a<5�a<��a<ܬa<��a<��a<E�a<�a<�a<��a<��a<�a<��a<��a<k�a<3�a<ީa<��a<D�a</�a<Ȩa<��a<G�a<էa<��a<1�a<�a<��a<C�a<�a<��a<@�a<ˤa<��a<�a<ϣa<n�a<��a<��a<(�a<�a<Y�a<��a<��a<$�a<ğa<G�a<��a<y�a<,�a<��a<D�a<�a<O�a<�a<~�a<*�a<��a<F�a<�a<l�a<3�a<��a<d�a<�a<��a<8�a<a<��a<��a<a<S�a<�a<��a<a�a<(�a<��a<��a<(�a<�a<��a<h�a<8�a<בa<��a<l�a<H�a<�a<ސa<Őa<��a<��a<%�a<7�a<��a<֏a<ޏa<��a<��a<��a<��a<i�a<s�a<�a<_�a<��a<\�a<��a<��a<��a<��a<��a<�a<�  �  �a<�a<>�a<Z�a<��a<��a<�a<�a<?�a<q�a<��a<�a<1�a<p�a<��a<�a<>�a<��a<͓a<!�a<s�a<ɔa<(�a<|�a<�a<.�a<��a<��a<d�a<ėa<"�a<��a<ߘa<T�a<ԙa<>�a<��a<�a<��a<��a<n�a<�a<S�a<��a<+�a<��a<�a<��a<��a<a�a<Ҡa<B�a<��a<,�a<��a<�a<|�a<�a<L�a<��a<�a<x�a<ޥa<D�a<��a<�a<f�a<��a<�a<{�a<֨a<'�a<n�a<��a<��a<T�a<��a<�a<�a<Q�a<��a<�a<-�a<i�a<��a<Ȭa<��a<0�a<U�a<��a<��a<έa<�a<�a<:�a<c�a<}�a<��a<��a<ٮa<�a<�a<�a<�a<+�a<?�a<F�a<S�a<T�a<a�a<Y�a<s�a<l�a<i�a<b�a<Y�a<C�a<\�a<H�a<E�a<�a<�a<�a<��a<�a<�a<��a<��a<��a<t�a<P�a<6�a<�a<�a<ŭa<��a<x�a<^�a<1�a<�a<Ϭa<��a<m�a<7�a<�a<ҫa<��a<k�a<+�a<��a<��a<v�a<3�a<��a<��a<c�a<"�a<��a<}�a<D�a<�a<��a<7�a<��a<��a<T�a<��a<��a<4�a<ޤa<~�a<!�a<��a<]�a<��a<��a<)�a<ġa<f�a<�a<��a<3�a<ğa<X�a<�a<w�a<�a<��a<:�a<Ԝa<e�a<��a<��a<$�a<ǚa<c�a<��a<��a<$�a<��a<V�a<��a<��a<)�a<��a<{�a<�a<˕a<u�a<�a<��a<f�a<!�a<ɓa<��a<1�a<�a<��a<]�a<�a<�a<��a<|�a<J�a<�a<ܐa<��a<��a<_�a<;�a< �a<��a<�a<ŏa<��a<��a<��a<��a<��a<v�a<n�a<^�a<��a<}�a<��a<��a<��a<��a<Ǐa<�a<�  �  ��a<�a<V�a<E�a<��a<��a<Ɛa<-�a<-�a<��a<��a<�a<1�a<X�a<��a<�a<L�a<|�a<�a<;�a<n�a<�a<�a<��a<ڕa<'�a<��a<�a<S�a<��a<!�a<v�a< �a<m�a<��a<&�a<��a<#�a<y�a<�a<X�a<ǜa<D�a<��a<D�a<~�a<'�a<}�a<�a<~�a<Ϡa<c�a<��a<6�a<��a< �a<s�a<ѣa<T�a<��a<1�a<|�a<��a<J�a<��a<�a<H�a<Чa<�a<l�a<��a<
�a<e�a<��a<�a<K�a<��a<Ъa<.�a<w�a<��a<ޫa<�a<U�a<��a<άa<��a<�a<e�a<m�a<��a<حa<�a<5�a<3�a<s�a<l�a<��a<��a<Үa<�a< �a<!�a<�a<I�a<$�a<Q�a<j�a<7�a<{�a<P�a<f�a<R�a<e�a<T�a<e�a<i�a<@�a<5�a<&�a<A�a<'�a<��a<��a<Ԯa<Үa<��a<��a<p�a<��a<[�a<�a<0�a<ۭa<�a<��a<|�a<^�a<�a<�a<Ĭa<��a<f�a<V�a<!�a<ͫa<��a<Q�a<8�a<�a<��a<��a<"�a<�a<��a<b�a<�a<ߨa<��a<%�a<ۧa<��a<Y�a<�a<��a<=�a<�a<��a</�a<��a<`�a<7�a<��a<X�a<�a<��a<J�a<ơa<p�a<��a<��a<*�a<��a<`�a<�a<��a<�a<��a<@�a<Ɯa<x�a<ߛa<��a<"�a<��a<J�a<ܙa<~�a<�a<ʘa<M�a<�a<�a<8�a<�a<b�a<�a<��a<a�a<�a<Ĕa<e�a<�a<ؓa<h�a<D�a<�a<��a<|�a<�a<��a<��a<|�a<0�a<�a<�a<��a<��a<Q�a<X�a<�a<�a<��a<��a<яa<��a<��a<r�a<}�a<h�a<z�a<��a<f�a<k�a<p�a<��a<��a<��a<ɏa<ˏa<�  �  �a<�a<>�a<Z�a<��a<��a<�a<�a<?�a<q�a<��a<�a<1�a<p�a<��a<�a<>�a<��a<͓a<!�a<s�a<ɔa<(�a<|�a<�a<.�a<��a<��a<d�a<ėa<"�a<��a<ߘa<T�a<ԙa<>�a<��a<�a<��a<��a<n�a<�a<S�a<��a<+�a<��a<�a<��a<��a<a�a<Ҡa<B�a<��a<,�a<��a<�a<|�a<�a<L�a<��a<�a<x�a<ޥa<D�a<��a<�a<f�a<��a<�a<{�a<֨a<'�a<n�a<��a<��a<T�a<��a<�a<�a<Q�a<��a<�a<-�a<i�a<��a<Ȭa<��a<0�a<U�a<��a<��a<έa<�a<�a<:�a<c�a<}�a<��a<��a<ٮa<�a<�a<�a<�a<+�a<?�a<F�a<S�a<T�a<a�a<Y�a<s�a<l�a<i�a<b�a<Y�a<C�a<\�a<H�a<E�a<�a<�a<�a<��a<�a<�a<��a<��a<��a<t�a<P�a<6�a<�a<�a<ŭa<��a<x�a<^�a<1�a<�a<Ϭa<��a<m�a<7�a<�a<ҫa<��a<k�a<+�a<��a<��a<v�a<3�a<��a<��a<c�a<"�a<��a<}�a<D�a<�a<��a<7�a<��a<��a<T�a<��a<��a<4�a<ޤa<~�a<!�a<��a<]�a<��a<��a<)�a<ġa<f�a<�a<��a<3�a<ğa<X�a<�a<w�a<�a<��a<:�a<Ԝa<e�a<��a<��a<$�a<ǚa<c�a<��a<��a<$�a<��a<V�a<��a<��a<)�a<��a<{�a<�a<˕a<u�a<�a<��a<f�a<!�a<ɓa<��a<1�a<�a<��a<]�a<�a<�a<��a<|�a<J�a<�a<ܐa<��a<��a<_�a<;�a< �a<��a<�a<ŏa<��a<��a<��a<��a<��a<v�a<n�a<^�a<��a<}�a<��a<��a<��a<��a<Ǐa<�a<�  �  �a<�a<*�a<n�a<��a<��a<��a<�a<d�a<s�a<��a<�a<�a<t�a<��a<��a<*�a<��a<ۓa<,�a<��a<��a<@�a<i�a<�a<4�a<��a<��a<G�a<ėa<�a<��a<�a<\�a<֙a< �a<��a<��a<��a<��a<]�a<˜a<@�a<��a<�a<��a<��a<��a<�a<`�a<�a<A�a<Сa<�a<��a<�a<m�a<�a<;�a<Ǥa<�a<��a<�a<N�a<��a<�a<|�a<��a<�a<j�a<��a<�a<S�a<ϩa<�a<b�a<��a<�a<-�a<X�a<��a<ūa<$�a<G�a<��a<¬a<�a<8�a<=�a<��a<��a<�a<�a<!�a<S�a<O�a<��a<��a<��a<Ȯa<�a<�a<�a<=�a<�a<V�a<C�a<E�a<m�a<K�a<h�a<[�a<e�a<Q�a<_�a<j�a<D�a<i�a<&�a<R�a<�a<"�a<�a<�a<�a<Ǯa<��a<��a<��a<g�a<G�a<Q�a<��a<�a<ǭa<��a<��a<I�a<5�a<��a<ܬa<��a<��a<E�a<�a<�a<��a<��a<�a<��a<��a<k�a<3�a<ީa<��a<D�a</�a<Ȩa<��a<G�a<էa<��a<1�a<�a<��a<C�a<�a<��a<@�a<ˤa<��a<�a<ϣa<n�a<��a<��a<(�a<�a<Y�a<��a<��a<$�a<ğa<G�a<��a<y�a<,�a<��a<D�a<�a<O�a<�a<~�a<*�a<��a<F�a<�a<l�a<3�a<��a<d�a<�a<��a<8�a<a<��a<��a<a<S�a<�a<��a<a�a<(�a<��a<��a<(�a<�a<��a<h�a<8�a<בa<��a<l�a<H�a<�a<ސa<Őa<��a<��a<%�a<7�a<��a<֏a<ޏa<��a<��a<��a<��a<i�a<s�a<�a<_�a<��a<\�a<��a<��a<��a<��a<��a<�a<�  �  �a<"�a<5�a<V�a<��a<��a<ސa<�a<D�a<g�a<��a<�a<&�a<p�a<��a<��a<9�a<��a<ۓa<�a<{�a<Ĕa<&�a<z�a<ܕa<.�a<��a<��a<Q�a<җa<�a<��a<��a<^�a<řa<#�a<��a<�a<��a<�a<p�a<՜a<E�a<��a<)�a<��a<�a<��a<�a<f�a<Ԡa<C�a<��a<&�a<��a<�a<s�a<�a<F�a<��a<�a<v�a<�a<<�a<��a<�a<g�a<��a< �a<p�a<¨a<'�a<e�a<��a<	�a<Y�a<��a<ڪa<)�a<p�a<��a<߫a<1�a<S�a<��a<Ǭa<�a<,�a<U�a<��a<��a<حa<�a<�a<=�a<`�a<��a<��a<��a<Ϯa<�a<��a< �a<�a<'�a<5�a<H�a<V�a<O�a<X�a<l�a<\�a<q�a<k�a<T�a<d�a<U�a<R�a<+�a<<�a<+�a<%�a<�a<��a<��a<ʮa<Ʈa<��a<��a<t�a<Q�a<2�a<	�a<�a<��a<��a<x�a<R�a<2�a<�a<ݬa<��a<k�a<E�a< �a<٫a<��a<i�a<)�a<��a<��a<p�a<9�a<�a<��a<_�a<�a<ܨa<��a<5�a<اa<��a<I�a<��a<��a<V�a<�a<��a<B�a<ܤa<�a<"�a<ãa<U�a<��a<��a<*�a<ϡa<_�a< �a<��a<*�a<ǟa<R�a<�a<{�a<�a<��a<2�a<՜a<g�a<��a<��a<-�a<��a<O�a<��a<~�a<�a<��a<[�a<�a<��a<3�a<ٖa<m�a<�a<ϕa<`�a<�a<��a<c�a<�a<ɓa<��a<)�a<�a<��a<f�a<"�a<�a<��a<x�a<F�a<�a<ڐa<��a<{�a<b�a<6�a<�a<��a<�a<��a<��a<��a<��a<��a<��a<h�a<y�a<p�a<x�a<a�a<��a<��a<��a<��a<ɏa<�a<�  �  ��a<�a<D�a<V�a<��a<��a<Аa<'�a<<�a<��a<��a<�a<5�a<^�a<��a<ޒa<O�a<y�a<ޓa<"�a<w�a<��a<�a<��a<ӕa<9�a<��a<��a<X�a<��a<0�a<�a<�a<P�a<̙a<O�a<��a<�a<s�a<��a<^�a<˜a<I�a<��a<>�a<��a<�a<�a<�a<~�a<͠a<[�a<��a<2�a<��a<�a<s�a<أa<V�a<��a<,�a<p�a<��a<J�a<��a<�a<X�a<Чa<�a<r�a<��a<�a<u�a<��a<
�a<F�a<��a<�a<�a<g�a<��a<��a<�a<X�a<��a<Ĭa<�a<�a<e�a<u�a<��a<٭a<�a<,�a<2�a<s�a<m�a<��a<��a<׮a<�a<�a<�a<�a<I�a</�a<H�a<V�a<M�a<j�a<W�a<g�a<V�a<g�a<]�a<Q�a<P�a<I�a<`�a<6�a<#�a<�a<�a<�a<ծa<֮a<��a<��a<��a<r�a<U�a<$�a<*�a<�a<ԭa<��a<v�a<a�a< �a<�a<��a<��a<c�a<H�a<	�a<իa<��a<Y�a<8�a<�a<��a<t�a<3�a<�a<��a<q�a<�a<Шa<y�a<=�a<�a<��a<I�a<�a<��a<D�a<�a<��a<-�a<�a<s�a<.�a<��a<[�a<�a<��a<B�a<��a<l�a<��a<��a<)�a<��a<b�a<۞a<��a<�a<��a<A�a<ǜa<w�a<�a<��a<�a<��a<N�a<�a<��a<�a<��a<I�a<�a<��a< �a<іa<g�a<(�a<��a<e�a<�a<��a<q�a<�a<ٓa<q�a<B�a<�a<��a<s�a<�a<��a<��a<y�a<<�a<�a<ܐa<��a<��a<Y�a<Y�a<�a<��a<�a<��a<��a<��a<��a<v�a<~�a<q�a<f�a<k�a<o�a<��a<�a<��a<��a<��a<̏a<̏a<�  �  �a<�a<8�a<i�a<�a<��a<�a< �a<6�a<~�a<��a<�a<$�a<_�a<��a<�a<C�a<��a<ۓa<)�a<q�a<��a<&�a<~�a<֕a<?�a<��a<�a<_�a<��a<'�a<��a<�a<d�a<��a<#�a<��a<�a<��a<��a<`�a<՜a<N�a<��a<.�a<��a<	�a<��a<��a<]�a<Ѡa<Q�a<��a<0�a<��a<�a<u�a<ԣa<M�a<��a<!�a<x�a<ۥa<E�a<��a<�a<c�a<ŧa<�a<v�a<˨a<�a<o�a<��a<�a<M�a<��a<تa<(�a<g�a<��a<�a<�a<`�a<��a<Ŭa<��a<&�a<T�a<��a<��a<έa<��a<&�a<@�a<f�a<s�a<��a<��a<Ʈa<�a<�a<�a<�a< �a<<�a<O�a<F�a<`�a<[�a<Z�a<q�a<_�a<`�a<k�a<b�a<]�a<G�a<2�a<1�a<3�a< �a<�a<��a<�a<߮a<��a<��a<��a<f�a<V�a<6�a<�a<�a<ҭa<��a<��a<P�a< �a<�a<Ƭa<��a<t�a<F�a<�a<ϫa<��a<i�a<-�a<�a<��a<s�a<.�a<��a<��a<h�a<#�a<Ҩa<��a<0�a<اa<��a<J�a<��a<��a<E�a<�a<��a<7�a<�a<��a<�a<ţa<^�a<�a<��a<8�a<ѡa<i�a<��a<��a<+�a<��a<Y�a<�a<��a<�a<��a<;�a<Ҝa<a�a<��a<��a<$�a<a<X�a<�a<��a<%�a<��a<O�a<�a<��a<2�a<Жa<y�a<�a<��a<l�a<�a<��a<p�a<�a<ȓa<��a<,�a<�a<��a<m�a<%�a<�a<��a<��a<8�a<�a<�a<��a<��a<T�a<0�a<�a<�a<؏a<ҏa<��a<��a<��a<�a<x�a<�a<w�a<x�a<l�a<g�a<{�a<��a<��a<��a<Ǐa<؏a<�  �  �a<"�a<4�a<a�a<��a<��a<�a<�a<N�a<n�a<��a<�a<*�a<p�a<��a<��a<:�a<��a<̓a<'�a<��a<Ôa<3�a<o�a<�a<.�a<��a<��a<O�a<ϗa<�a<��a<�a<d�a<˙a<3�a<��a<�a<��a<�a<k�a<՜a<>�a<ɝa<�a<��a<�a<��a<��a<b�a<�a<=�a<��a<"�a<��a<�a<s�a<�a<B�a<��a<�a<��a<ߥa<B�a<��a<��a<q�a<��a<'�a<k�a<èa<'�a<_�a<��a<�a<a�a<��a<�a<-�a<_�a<��a<իa<3�a<Q�a<��a<̬a<�a<5�a<H�a<��a<��a<حa< �a<�a<B�a<]�a<��a<��a<��a<ծa<�a<��a< �a</�a<#�a<?�a<J�a<I�a<^�a<Q�a<n�a<Y�a<n�a<b�a<W�a<Z�a<T�a<V�a<B�a<?�a<,�a<�a<�a<��a<�a<Ǯa<Ʈa<��a<��a<m�a<O�a<:�a<�a<��a<­a<��a<{�a<W�a<1�a<��a<ܬa<��a<q�a<6�a<�a<߫a<��a<v�a<�a<��a<��a<y�a<5�a<�a<��a<U�a<�a<Ψa<��a<<�a<�a<��a<C�a<��a<��a<P�a<�a<��a<L�a<Ѥa<��a<�a<ʣa<^�a<��a<��a<$�a<ϡa<\�a<�a<��a<)�a<ϟa<O�a<�a<t�a<%�a<��a<8�a<ޜa<[�a<�a<��a<4�a<��a<P�a<��a<y�a<#�a<��a<d�a<�a<��a<7�a<ɖa<u�a<�a<Еa<^�a<�a<a<]�a<%�a<��a<��a<,�a<�a<��a<\�a<'�a<�a<��a<t�a<F�a<�a<ܐa<��a<{�a<r�a<3�a< �a<�a<ۏa<Ϗa<��a<��a<��a<��a<y�a<k�a<o�a<o�a<|�a<x�a<��a<��a<��a<��a<��a<�a<�  �  �a<�a<>�a<Y�a<��a<��a<֐a<�a<9�a<z�a<��a<�a<1�a<b�a<��a<�a<B�a<��a<��a<"�a<t�a<ؔa<�a<|�a<��a<,�a<��a<��a<K�a<��a<'�a<��a<��a<T�a<��a<<�a<��a<�a<�a<��a<a�a<͜a<?�a<��a<)�a<��a<�a<��a<��a<o�a<ՠa<N�a<¡a<,�a<��a<��a<h�a<ݣa<K�a<��a<�a<}�a<�a<L�a<��a<�a<c�a<��a<�a<n�a<��a<�a<r�a<��a<
�a<E�a<��a<ܪa<�a<l�a<��a<�a<�a<K�a<��a<ˬa<�a<+�a<V�a<~�a<��a<ӭa<��a<(�a<G�a<d�a<x�a<��a<��a<׮a<�a<�a<�a<�a<5�a<4�a<E�a<X�a<U�a<_�a<e�a<W�a<\�a<h�a<e�a<_�a<\�a<B�a<W�a<-�a<+�a<#�a<�a<�a<ݮa<Ůa<��a<��a<��a<w�a<O�a<)�a<�a<�a<έa<��a<��a<^�a<#�a<�a<ʬa<��a<y�a<K�a<	�a<ҫa<��a<`�a<+�a<��a<��a<|�a<3�a<�a<��a<h�a<!�a<٨a<}�a<1�a<�a<��a<K�a<�a<��a<F�a<�a<��a<<�a<ܤa<�a<(�a<£a<a�a<�a<��a<5�a<ҡa<e�a<��a<��a<�a<��a<X�a<�a<��a<�a<��a<C�a<ќa<k�a<��a<��a<&�a<��a<K�a<�a<��a<�a<��a<G�a<�a<��a<'�a<Ֆa<x�a<�a<��a<X�a<�a<��a<_�a<�a<ʓa<z�a<=�a<�a<��a<o�a<,�a<�a<��a<c�a<8�a<�a<ߐa<��a<��a<X�a<E�a<�a<��a<�a<Əa<��a<��a<��a<|�a<��a<x�a<t�a<w�a<h�a<��a<w�a<��a<��a<��a<͏a<ԏa<�  �  �a<
�a<?�a<a�a<�a<��a<ڐa<�a<+�a<�a<��a<�a<�a<g�a<ʒa<�a<9�a<|�a<ԓa<'�a<l�a<Дa<�a<��a<͕a<=�a<��a<�a<t�a<��a<1�a<��a<�a<c�a<ęa<7�a<��a<#�a<r�a< �a<W�a<ܜa<R�a<��a<<�a<��a<�a<��a<��a<g�a<ɠa<Z�a<��a<.�a<��a<�a<��a<ңa<N�a<��a<&�a<s�a<�a<H�a<��a<�a<Z�a<ѧa<�a<w�a<Өa<
�a<{�a<��a<�a<F�a<��a<ݪa<&�a<k�a<��a<��a<�a<q�a<��a<��a<�a<�a<g�a<u�a<��a<˭a<��a<#�a<4�a<a�a<y�a<��a<��a<îa<�a<�a<�a<�a<-�a<:�a<I�a<O�a<T�a<f�a<S�a<y�a<a�a<c�a<e�a<M�a<h�a<9�a<E�a<*�a<;�a<�a<�a<�a<�a<�a<��a<��a<��a<g�a<W�a<.�a<�a<حa<ӭa<��a<w�a<L�a<(�a<�a<ͬa<��a<g�a<?�a<�a<˫a<��a<[�a<;�a<�a<��a<s�a<'�a<�a<��a<r�a<�a<Шa<��a<5�a<�a<��a<Z�a<�a<��a<<�a<��a<��a</�a<�a<v�a<-�a<��a<_�a<��a<��a<B�a<��a<g�a<�a<��a<;�a<��a<Z�a<ߞa<��a<�a<��a<?�a<Ȝa<u�a<�a<��a<�a<Úa<`�a<ܙa<��a<�a<Ƙa<H�a<�a<��a<0�a<Ֆa<f�a<'�a<��a<~�a<�a<��a<t�a<
�a<ۓa<p�a<8�a<�a<��a<j�a<�a<�a<��a<��a<B�a<�a<ܐa<��a<��a<H�a<=�a<�a< �a<�a<Əa<��a<��a<��a<��a<z�a<y�a<c�a<��a<_�a<{�a<s�a<��a<��a<��a<͏a<ڏa<�  �  �a<�a<;�a<d�a<}�a<��a<�a<�a<V�a<w�a<��a<�a<(�a<k�a<��a<��a<;�a<��a<ʓa</�a<��a<Ɣa<-�a<x�a<ѕa<;�a<��a<�a<R�a<��a<�a<��a<�a<^�a<͙a<6�a<��a<�a<�a<�a<W�a<؜a<<�a<��a<+�a<��a<�a<��a<��a<c�a<�a<F�a<��a<2�a<��a< �a<k�a<�a<M�a<��a<�a<��a<ߥa<G�a<��a<�a<i�a<��a<�a<g�a<Ǩa<�a<f�a<��a<�a<Y�a<��a<�a<'�a<a�a<��a<۫a<�a<V�a<��a<Ƭa<��a<$�a<S�a<��a<��a<حa<�a<�a<F�a<a�a<��a<��a<��a<Ϯa<�a<�a<
�a<4�a<%�a<B�a<B�a<H�a<\�a<[�a<d�a<[�a<g�a<V�a<g�a<T�a<R�a<X�a<H�a<@�a<'�a<�a<�a<�a<�a<ʮa<��a<��a<��a<e�a<L�a<:�a<�a<�a<˭a<��a<��a<U�a<-�a<�a<֬a<��a<z�a<5�a<�a<�a<��a<p�a<'�a<�a<��a<u�a<*�a<�a<��a<X�a<�a<˨a<��a<=�a<�a<��a<G�a<�a<��a<=�a<��a<��a<=�a<ޤa<��a<�a<ţa<c�a<��a<��a<-�a<ǡa<l�a<�a<��a<"�a<ȟa<Y�a<�a<{�a<#�a<��a<=�a<לa<d�a< �a<��a<*�a<��a<U�a<��a<��a<�a<��a<\�a<�a<��a<1�a<ʖa<v�a<�a<��a<b�a<�a<��a<k�a<�a<Ɠa<��a<2�a<�a<��a<]�a<+�a<�a<��a<c�a<>�a<�a<�a<��a<��a<w�a<4�a<#�a<��a<ُa<͏a<��a<��a<��a<��a<m�a<{�a<i�a<m�a<~�a<}�a<��a<��a<��a<��a<��a<�a<�  �  ߏa<9�a<.�a<[�a<��a<��a<�a<�a<G�a<[�a<��a<�a<�a<��a<��a<�a<*�a<��a<ϓa<�a<u�a<Ôa<*�a<j�a<�a<'�a<��a<�a<D�a<ڗa<�a<��a<�a<X�a<Ιa<+�a<��a< �a<��a<�a<s�a<�a<?�a<ѝa<�a<��a<�a<��a<�a<X�a<ܠa<-�a<ҡa<�a<��a<�a<m�a<�a<7�a<ɤa< �a<��a<եa<A�a<��a<��a<{�a<��a<1�a<s�a<Ϩa</�a<e�a<ͩa<��a<W�a<��a<�a<#�a<]�a<��a<ګa<9�a<L�a<��a<άa<�a<@�a<C�a<��a<��a<ͭa<�a<�a<T�a<L�a<��a<��a<Ǯa<ɮa<߮a<�a<�a<%�a<�a<=�a<;�a<S�a<\�a<K�a<��a<K�a<��a<f�a<f�a<l�a<D�a<X�a<:�a<C�a<�a<(�a<�a<��a<
�a<��a<ܮa<��a<��a<y�a<B�a<6�a<�a<��a<��a<��a<~�a<J�a<B�a<�a<�a<��a<��a<:�a<��a<ӫa<��a<l�a<�a<�a<��a<s�a<K�a<کa<ȩa<\�a</�a<Ψa<��a<>�a<�a<��a<7�a<�a<��a<X�a< �a<��a<S�a<Ĥa<��a<�a<��a<\�a<�a<��a<�a<�a<U�a<
�a<��a<$�a<џa<C�a<�a<f�a<�a<��a<7�a<Ԝa<U�a<�a<x�a<>�a<��a<\�a<�a<�a<0�a<��a<Y�a<�a<��a<-�a<ǖa<��a<�a<וa<X�a<!�a<Ĕa<V�a<0�a<��a<��a<-�a<�a<��a<X�a<9�a<ԑa<a<]�a<R�a<	�a<ِa<Őa<j�a<h�a<-�a<�a<�a<�a<Ώa<��a<��a<x�a<��a<}�a<z�a<��a<_�a<~�a<o�a<��a<��a<��a<��a<Ïa<�a<�  �  ��a<�a<9�a<f�a<��a<��a<ܐa<�a<D�a<w�a<��a<ߑa<�a<u�a<��a<�a<*�a<��a<דa<-�a<��a<ܔa<�a<��a<Օa<6�a<��a<��a<U�a<��a<�a<��a<�a<g�a<ҙa<=�a<��a<�a<{�a<�a<Z�a<Μa<C�a<��a<+�a<��a<�a<��a<��a<z�a<�a<K�a<ša<�a<��a<�a<|�a<�a<9�a<��a<�a<��a<��a<P�a<��a<�a<i�a<��a<�a<m�a<��a<�a<b�a<��a<
�a<T�a<��a<�a<,�a<h�a<��a<ګa<�a<R�a<��a<Ĭa<��a<%�a<W�a<z�a<��a<�a<�a<!�a<C�a<P�a<��a<��a<®a<Ůa<Ԯa<�a<�a<#�a<8�a<;�a<I�a<I�a<`�a<[�a<f�a<_�a<`�a<`�a<V�a<W�a<X�a<L�a<E�a<<�a<2�a<�a<�a<��a<�a<Юa<��a<��a<��a<h�a<T�a</�a<�a<�a<ʭa<��a<r�a<I�a<7�a<�a<�a<��a<r�a<A�a<�a<߫a<��a<]�a</�a<�a<��a<r�a<6�a<�a<��a<[�a<�a<Шa<��a<C�a<�a<��a<K�a<�a<��a<@�a<�a<��a<>�a<ޤa<��a< �a<ģa<e�a<�a<��a<2�a<աa<Q�a<��a<��a<2�a<��a<E�a<�a<��a<#�a<��a<F�a<ќa<e�a< �a<��a<)�a<��a<M�a<�a<{�a<�a<��a<V�a<��a<��a<6�a<іa<k�a<�a<��a<^�a<�a<��a<i�a<�a<˓a<u�a<C�a<��a<��a<h�a<(�a<ؑa<��a<�a<M�a<�a<ΐa<��a<��a<f�a<H�a<�a< �a<ۏa<ҏa<��a<��a<��a<��a<w�a<j�a<l�a<s�a<r�a<{�a<��a<��a<��a<��a<��a<܏a<�  �  !�a<�a<P�a<o�a<��a<ѐa<�a<>�a<K�a<��a<Ƒa<�a<D�a<��a<��a<�a<X�a<��a<��a<K�a<|�a<��a<'�a<��a<�a<O�a<��a<��a<v�a<ڗa<A�a<��a<�a<w�a<�a<i�a<��a<=�a<��a<��a<��a<�a<d�a<��a<N�a<��a<>�a<��a<�a<t�a<�a<s�a<̡a<R�a<��a<�a<}�a<�a<u�a<��a<@�a<��a<�a<c�a<��a<7�a<g�a<�a<�a<��a<ިa<3�a<w�a<��a<)�a<`�a<êa<��a<8�a<x�a<��a<��a<;�a<t�a<��a<ìa<�a<1�a<��a<��a<խa<֭a<�a<C�a<P�a<��a<��a<��a<��a<�a<
�a<�a<9�a<#�a<Q�a<J�a<Z�a<i�a<\�a<p�a<a�a<��a<w�a<~�a<\�a<d�a<y�a<e�a<r�a<P�a<J�a<+�a<�a<�a<��a<�a<��a<��a<��a<��a<j�a<8�a<;�a<�a<��a<��a<��a<k�a<;�a<�a<�a<��a<��a<^�a<,�a<իa<̫a<e�a<V�a<��a<Ǫa<u�a<3�a<�a<éa<~�a<�a<�a<��a<Q�a<�a<��a<o�a<�a<��a<c�a<�a<��a<;�a<��a<��a<L�a<ˣa<y�a<�a<��a<Y�a<ܡa<��a<�a<��a<4�a<ҟa<��a<��a<��a<!�a<��a<\�a<؜a<��a<�a<��a<'�a<՚a<p�a<	�a<��a<�a<ߘa<h�a<�a<��a<H�a<�a<n�a<4�a<ߕa<��a<�a<��a<��a<'�a<��a<��a<b�a<��a<ʒa<��a<;�a<�a<ȑa<|�a<Q�a<)�a<
�a<Ɛa<��a<l�a<h�a<2�a<�a<�a<ԏa<͏a<��a<��a<��a<��a<w�a<��a<��a<��a<��a<��a<��a<��a<��a<�a<��a<�  �  �a<<�a<Z�a<t�a<��a<ΐa<�a<(�a<]�a<��a<��a<�a<5�a<��a<ϒa<�a<D�a<��a<�a<C�a<��a<�a<5�a<��a<�a<Q�a<��a<�a<d�a<՗a<>�a<��a<�a<s�a<әa<?�a<��a<,�a<��a<�a<�a<ܜa<b�a<ߝa<N�a<��a<+�a<��a<�a<x�a<��a<X�a<ϡa<9�a<��a<(�a<��a<��a<U�a<Ťa<#�a<��a<�a<V�a<��a< �a<m�a<ߧa<:�a<��a<ʨa<3�a<��a<ةa<�a<e�a<��a<�a<9�a<{�a<ȫa<��a<9�a<_�a<��a<�a<�a<3�a<r�a<��a<��a<�a<�a<&�a<V�a<e�a<��a<��a<خa<׮a<��a<�a<!�a<5�a<A�a<H�a<Y�a<a�a<e�a<w�a<�a<w�a<m�a<{�a<~�a<x�a<i�a<a�a<F�a<J�a<>�a<9�a<.�a<�a<�a<�a<ٮa<��a<��a<|�a<g�a<?�a<%�a<�a<�a<��a<��a<[�a<N�a<�a<��a<��a<��a<F�a<$�a<�a<��a<s�a<H�a<��a<Ȫa<��a<Q�a<��a<��a<{�a<?�a<�a<��a<@�a<�a<��a<_�a<�a<��a<b�a<��a<��a<^�a<��a<��a<9�a<Уa<m�a<
�a<��a<?�a<�a<r�a<�a<��a<K�a<֟a<c�a<��a<��a<0�a<��a<O�a<�a<��a<�a<��a<K�a<ښa<[�a<	�a<��a<@�a<՘a<l�a<��a<��a<H�a<�a<��a<7�a<ܕa<q�a<4�a<��a<��a<)�a<�a<��a<N�a<�a<ƒa<t�a<B�a<�a<Ցa<��a<i�a<�a<��a<a<��a<~�a<W�a</�a<�a<��a<ݏa<ӏa<ďa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<؏a<�a<��a<�  �  �a<7�a<C�a<��a<��a<Ӑa<��a<�a<i�a<��a<ϑa<�a<:�a<��a<��a<�a<E�a<��a<�a<B�a<��a<ٔa<K�a<��a<��a<N�a<��a<�a<f�a<�a<�a<��a<��a<x�a<�a<D�a<њa<�a<��a<��a<z�a<�a<X�a<Нa<5�a<��a<&�a<��a<�a<z�a<�a<T�a<�a<:�a<��a<
�a<r�a<��a<R�a<�a<!�a<��a<��a<Y�a<Ѧa<�a<��a<Ƨa<'�a<}�a<Ҩa<4�a<l�a<ԩa<�a<y�a<��a<��a<B�a<h�a<īa<�a<C�a<c�a<��a<̬a<�a<E�a<k�a<��a<��a<�a<�a<*�a<s�a<e�a<��a<��a<Ȯa<ޮa<�a<�a<�a<A�a<4�a<P�a<c�a<h�a<v�a<]�a<w�a<t�a<~�a<h�a<n�a<p�a<_�a<w�a<J�a<`�a<9�a<,�a<!�a<��a<�a<�a<Ԯa<��a<��a<��a<m�a<L�a<�a<�a<ۭa<��a<��a<`�a<A�a<��a<�a<��a<��a<N�a<#�a<�a<��a<��a<C�a<�a<ƪa<w�a<M�a<��a<̩a<\�a<8�a<ըa<��a<V�a<��a<ħa<I�a<�a<��a<]�a<�a<��a<O�a<�a<��a<5�a<�a<s�a<�a<��a<:�a<��a<t�a<�a<��a<)�a<۟a<`�a<�a<��a<;�a<��a<R�a<��a<{�a<�a<��a<8�a<̚a<d�a<�a<��a<<�a<��a<��a<�a<��a<R�a<֖a<��a<�a<�a<u�a<+�a<ǔa<{�a<;�a<�a<��a<E�a<
�a<ɒa<w�a<^�a<�a<ԑa<x�a<Z�a<%�a<�a<֐a<��a<��a<J�a<7�a<!�a<�a<�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ˏa<Ώa<�a<�  �  �a<2�a<R�a<~�a<��a<ΐa<�a<2�a<N�a<��a<ʑa<��a<A�a<��a<̒a<�a<Q�a<��a<�a<?�a<��a<�a</�a<��a<�a<S�a<��a<�a<n�a<Зa<6�a<��a<�a<u�a<יa<H�a<��a</�a<��a<�a<|�a<�a<c�a<ϝa<F�a<��a< �a<��a<�a<��a<�a<e�a<ša<9�a<��a<!�a<��a<��a<Y�a<��a<2�a<��a<��a<_�a<��a<�a<v�a<اa<+�a<��a<֨a<.�a<�a<٩a< �a<a�a<��a<�a<6�a<��a<ëa<��a</�a<j�a<��a<Ѭa<�a<8�a<i�a<��a<̭a<�a<�a<6�a<J�a<q�a<��a<��a<Ѯa<�a<�a<	�a<$�a<&�a<H�a<H�a<X�a<a�a<n�a<n�a<s�a<}�a<s�a<v�a<t�a<��a<p�a<V�a<X�a<B�a<F�a<A�a<#�a<�a<��a<�a<Ϯa<��a<��a<��a<h�a<<�a<.�a<��a<�a<��a<��a<h�a<G�a<�a<�a<��a<z�a<W�a< �a<�a<��a<m�a<B�a<��a<˪a<~�a<H�a< �a<��a<r�a<7�a<�a<��a<C�a<��a<��a<b�a<�a<��a<^�a<�a<��a<O�a<��a<��a<.�a<ͣa<t�a<�a<��a<L�a<աa<s�a<�a<��a<D�a<ڟa<f�a<��a<��a<$�a<��a<X�a<�a<w�a<�a<��a<<�a<֚a<h�a<�a<��a<A�a<טa<h�a<�a<��a<F�a<�a<��a<.�a<ӕa<|�a<+�a<͔a<��a<.�a<�a<��a<Z�a<�a<��a<��a<5�a<��a<ёa<��a<b�a<(�a<�a<Ȑa<��a<p�a<^�a</�a<�a<��a<�a<ʏa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ȏa<͏a<ߏa<��a<�  �   �a<,�a<X�a<q�a<��a<ܐa<�a<?�a<G�a<��a<ˑa<
�a<I�a<w�a<ܒa<��a<f�a<��a<��a<B�a<��a<��a<(�a<��a<�a<P�a<��a<�a<y�a<ʗa<K�a<��a<�a<s�a<�a<g�a<��a<1�a<��a<�a<�a<�a<l�a<ǝa<J�a<��a<5�a<��a<�a<��a<ݠa<t�a<ša<V�a<��a<�a<��a<�a<t�a<��a<B�a<��a<�a<b�a<��a<,�a<f�a<ۧa<&�a<��a<ڨa<-�a<��a<��a<#�a<\�a<êa<��a<3�a<��a<��a<�a<)�a<q�a<��a<Ԭa<�a<-�a<��a<��a<ԭa<�a<�a<B�a<O�a<��a<~�a<��a<®a<�a<�a<
�a<2�a<�a<W�a<C�a<d�a<f�a<_�a<x�a<n�a<��a<m�a<��a<r�a<f�a<r�a<T�a<w�a<C�a<F�a<.�a<�a<�a<�a<�a<ɮa<��a<��a<��a<v�a<4�a<;�a<�a<�a<��a<��a<o�a<2�a<(�a<Ҭa<Ǭa<��a<`�a<#�a<߫a<ɫa<f�a<X�a<��a<Ǫa<��a<B�a<�a<��a<��a< �a<�a<��a<O�a<�a<��a<d�a<��a<��a<a�a< �a<��a<G�a<��a<��a<D�a<ңa<r�a<!�a<��a<Z�a<աa<��a<�a<��a<E�a<a<��a<��a<��a<�a<ʝa<[�a<��a<��a<�a<��a<7�a<��a<k�a<�a<��a< �a<٘a<c�a<�a<��a<B�a<�a<w�a<@�a<͕a<��a<*�a<Дa<��a<#�a<��a<��a<b�a<�a<��a<��a<;�a<�a<��a<��a<S�a<'�a<�a<ɐa<��a<g�a<m�a<*�a<!�a<��a<׏a<ԏa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<Ïa<�a<�a<�  �  �a</�a<S�a<��a<��a<Ða<��a<)�a<e�a<��a<��a<�a<G�a<��a<ђa<�a<X�a<��a<�a<=�a<��a<�a<A�a<��a<�a<\�a<��a<�a<x�a<ޗa<4�a<��a<	�a<t�a<�a<J�a<��a<*�a<��a<�a<{�a<��a<_�a<ɝa<I�a<a<�a<��a<�a<��a<�a<]�a<ǡa<A�a<��a<!�a<��a<��a<]�a<��a<'�a<��a<��a<X�a<��a<�a<��a<ݧa<(�a<��a<�a</�a<��a<ϩa<�a<i�a<��a<�a<7�a<y�a<��a<�a<9�a<u�a<��a<լa<�a<@�a<]�a<��a<��a<�a<�a<*�a<Q�a<v�a<��a<��a<ʮa<�a<��a<�a<"�a<<�a<C�a<M�a<S�a<T�a<y�a<r�a<q�a<v�a<��a<t�a<y�a<j�a<i�a<h�a<P�a<T�a<C�a<.�a<$�a<�a<	�a<�a<̮a<��a<��a<w�a<]�a<H�a<&�a<�a<�a<��a<��a<m�a<;�a<�a<�a<��a<��a<J�a<�a<�a<��a<�a<4�a<�a<Ԫa<��a<@�a<
�a<ǩa<p�a<0�a<�a<��a<P�a<��a<��a<\�a<	�a<��a<]�a<�a<��a<I�a<��a<��a<'�a<ѣa<n�a<�a<��a<C�a<ءa<{�a<�a<��a<D�a<֟a<j�a<��a<��a<+�a<ŝa<Q�a<�a<o�a<�a<��a<8�a<֚a<w�a<�a<��a<7�a<јa<q�a<�a<��a<F�a<�a<��a<*�a<ݕa<��a<'�a<єa<��a<6�a<֓a<��a<N�a<�a<��a<w�a<=�a<�a<Ǒa<��a<[�a</�a<��a<��a<��a<��a<Y�a<5�a<�a<�a<�a<Ϗa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<Ώa<ُa<�a<�  �  �a<I�a<F�a<~�a<��a<��a<�a<�a<i�a<��a<Ցa<�a<;�a<��a<��a<�a<D�a<��a<�a<4�a<��a<Ӕa<S�a<��a<��a<A�a<��a<�a<a�a<��a<)�a<��a<��a<u�a<�a<A�a<͚a<�a<��a<�a<t�a<�a<T�a<�a<,�a<ʞa<�a<��a<�a<t�a<��a<P�a<�a<-�a<��a<�a<��a<�a<I�a<ڤa< �a<��a<�a<V�a<Ǧa<	�a<��a<��a<<�a<}�a<ըa<+�a<r�a<ߩa<�a<t�a<��a<��a<>�a<j�a<ͫa<�a<;�a<a�a<��a<٬a<��a<M�a<R�a<��a<��a<�a<�a<0�a<b�a<c�a<��a<��a<Үa<߮a<�a<�a<�a<>�a</�a<[�a<S�a<Y�a<u�a<^�a<��a<d�a<��a<k�a<z�a<s�a<Y�a<r�a<D�a<Y�a<6�a<1�a<-�a<�a<
�a<Ԯa<�a<��a<��a<��a<X�a<Y�a<�a<�a<έa<ŭa<��a<b�a<J�a<�a<��a<��a<��a<V�a<�a<�a<��a<��a<+�a<�a<��a<��a<N�a<�a<ɩa<f�a<?�a<٨a<��a<T�a<�a<��a<I�a<�a<��a<W�a<�a<��a<c�a<ݤa<��a<'�a<ڣa<t�a<�a<��a<7�a<��a<g�a<�a<��a<9�a<�a<W�a<�a<��a<+�a<��a<N�a<��a<k�a<(�a<��a<L�a<͚a<g�a<�a<��a<H�a<��a<{�a< �a<��a<M�a<ٖa<��a<�a<ޕa<s�a<,�a<Ԕa<r�a<C�a<̓a<��a<A�a<�a<��a<~�a<N�a<�a<ۑa<��a<d�a<&�a<�a<ِa<��a<��a<E�a<B�a<�a<�a<�a<��a<ҏa<��a<��a<��a<��a<��a<{�a<��a<��a<��a<��a<��a<׏a<ҏa<�a<�  �  �a<6�a<K�a<q�a<��a<Ȑa<�a<+�a<g�a<��a<ˑa<�a<F�a<��a<��a<�a<U�a<��a<�a<=�a<��a<�a<8�a<��a<��a<>�a<��a<�a<s�a<ݗa<<�a<��a<
�a<{�a<�a<R�a<��a<*�a<��a< �a<x�a<�a<^�a<ѝa<4�a<��a<6�a<��a<�a<��a<��a<\�a<ӡa<?�a<��a<�a<��a<��a<_�a<ʤa<.�a<��a<�a<\�a<��a<&�a<��a<ŧa<,�a<��a<�a<,�a<u�a<ǩa<�a<d�a<��a<��a<<�a<{�a<��a<��a<7�a<p�a<��a<Ӭa<��a<I�a<o�a<��a<��a<��a<�a<7�a<S�a<u�a<��a<��a<ήa<�a<��a<�a<�a<;�a<G�a<G�a<W�a<s�a<g�a<f�a<z�a<v�a<}�a<w�a<k�a<q�a<l�a<^�a<c�a<I�a<C�a<4�a<�a<�a<�a<�a<Ӯa<��a<��a<��a<a�a<?�a<(�a<�a<֭a<��a<��a<l�a<E�a<�a<�a<��a<��a<X�a<�a<��a<��a<v�a<C�a<�a<��a<�a<B�a<�a<Ʃa<y�a<#�a<�a<��a<O�a<�a<��a<]�a<�a<��a<[�a<�a<��a<Q�a<�a<��a<D�a<ңa<t�a<�a<��a<C�a<�a<x�a<�a<��a<=�a<ڟa<l�a<�a<��a<.�a<ʝa<U�a<�a<��a<�a<��a<=�a<Қa<q�a<�a<��a</�a<Ϙa<k�a<�a<��a<K�a<�a<��a<.�a<ڕa<��a<#�a<Δa<r�a<?�a<�a<��a<N�a<�a<a<��a<?�a<�a<ϑa<��a<_�a<(�a<��a<͐a<��a<��a<]�a<.�a<�a<�a<ߏa<Ïa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<Ïa<�a<�a<�  �  +�a<�a<h�a<t�a<��a<̐a<�a<3�a<P�a<��a<��a<�a<G�a<|�a<�a< �a<^�a<��a<�a<H�a<��a<�a<4�a<��a<�a<S�a<��a<�a<��a<��a<M�a<��a<�a<n�a<ڙa<[�a<��a<?�a<��a<�a<u�a<�a<p�a<��a<X�a<��a<.�a<��a<�a<��a<�a<p�a<��a<G�a<��a<(�a<��a<�a<g�a<��a<>�a<��a<��a<f�a<��a<"�a<g�a<�a<!�a<��a<�a<"�a<��a<ũa<0�a<P�a<��a<�a<*�a<��a<��a<�a<�a<~�a<��a<جa<�a<-�a<r�a<��a<ϭa<�a<�a<9�a<D�a<|�a<��a<̮a<Ǯa<�a<��a< �a<0�a<&�a<K�a<I�a<V�a<b�a<a�a<��a<_�a<��a<j�a<}�a<~�a<m�a<x�a<P�a<o�a<?�a<J�a<5�a<&�a<�a<�a<��a<��a<ˮa<��a<|�a<f�a<?�a<0�a<��a<�a<��a<��a<m�a<8�a<3�a<جa<��a<y�a<T�a<)�a<�a<��a<r�a<H�a<��a<˪a<��a<<�a<�a<��a<��a<*�a<�a<��a<G�a<�a<��a<q�a<�a<Ʀa<W�a<�a<��a<=�a<	�a<��a<<�a<Уa<y�a<�a<��a<W�a<ˡa<��a<�a<��a<R�a<Οa<t�a<�a<��a<(�a<a<^�a<�a<��a<�a<��a<2�a<��a<t�a<��a<��a<-�a<�a<W�a<�a<��a<9�a<��a<��a<C�a<��a<��a<#�a<Ԕa<��a<$�a<�a<��a<]�a< �a<Ȓa<��a</�a<
�a<��a<��a<Y�a<(�a<��a<��a<��a<p�a<a�a<0�a<�a<��a<ُa<�a<��a<��a<��a<��a<��a<��a<��a<|�a<��a<��a<��a<��a<Ϗa<�a<�a<�  �   �a<(�a<X�a<x�a<��a<Ɛa<��a<'�a<W�a<��a<̑a<�a<G�a<y�a<ƒa<�a<^�a<��a<�a<>�a<��a<�a<;�a<��a<�a<K�a<��a<�a<v�a<ʗa<>�a<��a<�a<s�a<�a<S�a<a<&�a<��a<�a<x�a<�a<j�a<Ɲa<A�a<��a</�a<��a<�a<}�a<�a<_�a<ڡa<H�a<��a<�a<��a<�a<e�a<Ѥa<.�a<��a<��a<\�a<��a< �a<u�a<ϧa<%�a<��a<ڨa<(�a<��a<©a<�a<k�a<��a<��a<7�a<s�a<��a<��a<)�a<q�a<��a<Ѭa<�a<;�a<l�a<��a<ƭa<�a<�a<1�a<f�a<|�a<��a<��a<��a<�a<�a<�a<�a<-�a<?�a<Q�a<P�a<g�a<g�a<s�a<h�a<��a<n�a<x�a<x�a<d�a<f�a<i�a<\�a<V�a<?�a<(�a<#�a<�a<�a<�a<Ůa<��a<��a<��a<`�a<F�a<$�a<��a<ܭa<��a<��a<m�a<4�a<�a<۬a<��a<��a<S�a<�a<�a<��a<x�a<=�a<�a<êa<��a<@�a<�a<��a<{�a<)�a<ݨa<��a<T�a<�a<��a<Y�a<��a<��a<[�a<�a<��a<F�a<�a<��a<>�a<Уa<u�a<�a<��a<F�a<�a<��a<�a<��a<9�a<ҟa<r�a<�a<��a<*�a<��a<U�a<�a<��a<�a<��a<6�a<ۚa<k�a<��a<��a<*�a<̘a<r�a<�a<��a<F�a<�a<��a<4�a<̕a<��a<&�a<͔a<z�a<2�a<�a<��a<T�a<�a<Ēa<~�a<R�a<
�a<��a<��a<Q�a<)�a<�a<Ґa<��a<w�a<U�a<8�a<�a< �a<ߏa<Џa<��a<��a<��a<��a<��a<�a<��a<��a<��a<��a<��a<��a<͏a<�a<�a<�  �  �a<<�a<[�a<~�a<��a<��a<��a<�a<e�a<|�a<͑a<��a<>�a<��a<��a<#�a<H�a<��a<�a<3�a<��a<�a<?�a<��a<��a<S�a<��a<�a<e�a<�a<0�a<��a<�a<s�a<ܙa<6�a<ƚa<�a<��a<��a<��a<�a<W�a<�a<C�a<��a<�a<��a<�a<v�a<��a<K�a<ۡa<-�a<��a< �a<��a<�a<K�a<Τa<�a<��a<�a<U�a<��a<�a<��a<ҧa<B�a<��a<ۨa<<�a<r�a<�a<�a<l�a<��a<�a<8�a<x�a<ϫa<�a<E�a<f�a<��a<�a<�a<G�a<[�a<��a<��a<�a<�a<%�a<X�a<c�a<��a<��a<Ԯa<�a<�a<�a<�a<?�a<7�a<V�a<H�a<e�a<q�a<u�a<��a<i�a<��a<y�a<q�a<��a<Z�a<h�a<<�a<Q�a<4�a<H�a<$�a<�a<�a<خa<ٮa<��a<��a<��a<S�a<J�a<�a<�a<ɭa<��a<��a<d�a<O�a<�a<��a<��a<��a<J�a<�a<�a<��a<|�a<-�a<�a<˪a<��a<F�a<��a<ϩa<m�a<=�a<�a<��a<I�a<�a<��a<M�a<&�a<��a<e�a<�a<��a<b�a<�a<��a<-�a<ʣa<s�a<�a<��a<2�a<�a<g�a< �a<��a<?�a<�a<X�a<�a<��a<4�a<��a<M�a<��a<q�a<�a<��a<R�a<Кa<m�a<�a<��a<P�a<Øa<s�a<�a<��a<G�a<�a<��a<$�a<�a<x�a<(�a<�a<��a<=�a<Փa<��a<J�a<�a<��a<s�a<D�a<�a<ߑa<��a<f�a<(�a<�a<Ԑa<��a<��a<M�a<=�a<�a<��a<�a<ҏa<Ǐa<��a<��a<��a<��a<��a<{�a<��a<x�a<��a<��a<Ϗa<Ώa<��a<�a<�  �  �a<,�a<Y�a<q�a<��a<Аa<�a<"�a<S�a<��a<ؑa<�a<@�a<~�a<��a<�a<V�a<��a<��a<A�a<��a<�a<G�a<��a<�a<O�a<��a<�a<o�a<ٗa<9�a<��a<�a<l�a<�a<W�a<Śa<�a<��a<��a<~�a<�a<\�a<ʝa<J�a<��a<0�a<��a<�a<p�a<��a<h�a<ޡa<B�a<��a<�a<z�a<��a<c�a<Ҥa<8�a<��a<�a<c�a<ʦa<%�a<o�a<ڧa<&�a<��a<ըa<3�a<s�a<̩a<�a<h�a<��a<�a<3�a<v�a<��a<�a<8�a<h�a<��a<Ӭa<�a<0�a<t�a<��a<ĭa<٭a<�a<@�a<]�a<x�a<��a<��a<��a<�a<��a<�a<#�a</�a<6�a<Y�a<_�a<b�a<`�a<x�a<n�a<w�a<t�a<{�a<f�a<s�a<W�a<r�a<`�a<\�a<1�a<5�a<�a<�a<��a<�a<ɮa<��a<��a<~�a<j�a<O�a<�a<��a<�a<ȭa<��a<g�a<:�a<�a<�a<��a<��a<^�a<"�a<ݫa<��a<��a<G�a<��a<ƪa<��a<?�a<�a<��a<v�a<)�a<�a<��a<[�a<	�a<��a<O�a<	�a<��a<a�a<�a<��a<I�a<��a<��a<>�a<�a<�a<�a<��a<N�a<�a<|�a<�a<��a<1�a<֟a<p�a<�a<��a<0�a<��a<\�a<��a<��a<	�a<��a<7�a<Кa<g�a<	�a<��a<4�a<ǘa<o�a<�a<��a<B�a<�a<��a<)�a<ەa<z�a<"�a<ϔa<��a<&�a<�a<��a<R�a<��a<ƒa<��a<I�a<�a<ɑa<��a<P�a<'�a<��a<ܐa<��a<y�a<L�a<A�a<�a<��a<؏a<Տa<��a<��a<��a<��a<��a<��a<y�a<��a<��a<��a<��a<��a<��a<�a<��a<�  �  -�a<"�a<]�a<v�a<��a<Ða<�a<3�a<[�a<��a<��a<��a<I�a<��a<�a<�a<g�a<��a<ٓa<E�a<��a<�a<(�a<��a<ߕa<X�a<��a<�a<{�a<Ɨa<S�a<��a<�a<v�a<ՙa<9�a<��a<;�a<��a<�a<�a<ۜa<o�a<��a<_�a<��a<0�a<��a<�a<��a<��a<a�a<��a<B�a<��a<&�a<��a<�a<j�a<��a<*�a<��a<��a<Y�a<��a<'�a<i�a<�a<�a<��a<˨a<)�a<��a<ȩa<2�a<a�a<��a<�a<5�a<��a<��a<�a<$�a<h�a<��a<Ѭa<�a<&�a<s�a<��a<ȭa<�a<�a<%�a<?�a<��a<��a<ήa<ͮa<�a<�a<�a<'�a<4�a<G�a<:�a<J�a<`�a<b�a<��a<`�a<��a<b�a<��a<{�a<o�a<j�a<c�a<H�a<L�a<C�a<8�a<#�a<$�a<�a<��a<��a<��a<��a<z�a<]�a<3�a</�a<�a<�a<��a<��a<p�a<B�a</�a<�a<Ȭa<v�a<>�a<&�a<�a<��a<e�a<B�a<�a<Ъa<��a<D�a<�a<��a<��a<*�a<��a<��a<B�a<�a<��a<m�a<�a<Ŧa<b�a<��a<��a<@�a<�a<��a<>�a<��a<m�a<�a<��a<G�a<ġa<|�a<�a<��a<Q�a<ҟa<w�a<�a<��a<0�a<Ɲa<R�a<Ӝa<��a<�a<ƛa<,�a<ޚa<]�a<��a<��a<0�a<�a<h�a<��a<��a<E�a<��a<��a<C�a<Ǖa<z�a<,�a<̔a<��a<�a<�a<��a<V�a<�a<ʒa<s�a<*�a<�a<Ƒa<��a<^�a<-�a<�a<��a<��a<~�a<]�a<!�a<�a<��a<ڏa<ߏa<��a<ďa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<͏a<��a<�a<�  �  �a<,�a<Y�a<q�a<��a<Аa<�a<"�a<S�a<��a<ؑa<�a<@�a<~�a<��a<�a<V�a<��a<��a<A�a<��a<�a<G�a<��a<�a<O�a<��a<�a<o�a<ٗa<9�a<��a<�a<l�a<�a<W�a<Śa<�a<��a<��a<~�a<�a<\�a<ʝa<J�a<��a<0�a<��a<�a<p�a<��a<h�a<ޡa<B�a<��a<�a<z�a<��a<c�a<Ҥa<8�a<��a<�a<c�a<ʦa<%�a<o�a<ڧa<&�a<��a<ըa<3�a<s�a<̩a<�a<h�a<��a<�a<3�a<v�a<��a<�a<8�a<h�a<��a<Ӭa<�a<0�a<t�a<��a<ĭa<٭a<�a<@�a<]�a<x�a<��a<��a<��a<�a<��a<�a<#�a</�a<6�a<Y�a<_�a<b�a<`�a<x�a<n�a<w�a<t�a<{�a<f�a<s�a<W�a<r�a<`�a<\�a<1�a<5�a<�a<�a<��a<�a<ɮa<��a<��a<~�a<j�a<O�a<�a<��a<�a<ȭa<��a<g�a<:�a<�a<�a<��a<��a<^�a<"�a<ݫa<��a<��a<G�a<��a<ƪa<��a<?�a<�a<��a<v�a<)�a<�a<��a<[�a<	�a<��a<O�a<	�a<��a<a�a<�a<��a<I�a<��a<��a<>�a<�a<�a<�a<��a<N�a<�a<|�a<�a<��a<1�a<֟a<p�a<�a<��a<0�a<��a<\�a<��a<��a<	�a<��a<7�a<Кa<g�a<	�a<��a<4�a<ǘa<o�a<�a<��a<B�a<�a<��a<)�a<ەa<z�a<"�a<ϔa<��a<&�a<�a<��a<R�a<��a<ƒa<��a<I�a<�a<ɑa<��a<P�a<'�a<��a<ܐa<��a<y�a<L�a<A�a<�a<��a<؏a<Տa<��a<��a<��a<��a<��a<��a<y�a<��a<��a<��a<��a<��a<��a<�a<��a<�  �  �a<<�a<[�a<~�a<��a<��a<��a<�a<e�a<|�a<͑a<��a<>�a<��a<��a<#�a<H�a<��a<�a<3�a<��a<�a<?�a<��a<��a<S�a<��a<�a<e�a<�a<0�a<��a<�a<s�a<ܙa<6�a<ƚa<�a<��a<��a<��a<�a<W�a<�a<C�a<��a<�a<��a<�a<v�a<��a<K�a<ۡa<-�a<��a< �a<��a<�a<K�a<Τa<�a<��a<�a<U�a<��a<�a<��a<ҧa<B�a<��a<ۨa<<�a<r�a<�a<�a<l�a<��a<�a<8�a<x�a<ϫa<�a<E�a<f�a<��a<�a<�a<G�a<[�a<��a<��a<�a<�a<%�a<X�a<c�a<��a<��a<Ԯa<�a<�a<�a<�a<?�a<7�a<V�a<H�a<e�a<q�a<u�a<��a<i�a<��a<y�a<q�a<��a<Z�a<h�a<<�a<Q�a<4�a<H�a<$�a<�a<�a<خa<ٮa<��a<��a<��a<S�a<J�a<�a<�a<ɭa<��a<��a<d�a<O�a<�a<��a<��a<��a<J�a<�a<�a<��a<|�a<-�a<�a<˪a<��a<F�a<��a<ϩa<m�a<=�a<�a<��a<I�a<�a<��a<M�a<&�a<��a<e�a<�a<��a<b�a<�a<��a<-�a<ʣa<s�a<�a<��a<2�a<�a<g�a< �a<��a<?�a<�a<X�a<�a<��a<4�a<��a<M�a<��a<q�a<�a<��a<R�a<Кa<m�a<�a<��a<P�a<Øa<s�a<�a<��a<G�a<�a<��a<$�a<�a<x�a<(�a<�a<��a<=�a<Փa<��a<J�a<�a<��a<s�a<D�a<�a<ߑa<��a<f�a<(�a<�a<Ԑa<��a<��a<M�a<=�a<�a<��a<�a<ҏa<Ǐa<��a<��a<��a<��a<��a<{�a<��a<x�a<��a<��a<Ϗa<Ώa<��a<�a<�  �   �a<(�a<X�a<x�a<��a<Ɛa<��a<'�a<W�a<��a<̑a<�a<G�a<y�a<ƒa<�a<^�a<��a<�a<>�a<��a<�a<;�a<��a<�a<K�a<��a<�a<v�a<ʗa<>�a<��a<�a<s�a<�a<S�a<a<&�a<��a<�a<x�a<�a<j�a<Ɲa<A�a<��a</�a<��a<�a<}�a<�a<_�a<ڡa<H�a<��a<�a<��a<�a<e�a<Ѥa<.�a<��a<��a<\�a<��a< �a<u�a<ϧa<%�a<��a<ڨa<(�a<��a<©a<�a<k�a<��a<��a<7�a<s�a<��a<��a<)�a<q�a<��a<Ѭa<�a<;�a<l�a<��a<ƭa<�a<�a<1�a<f�a<|�a<��a<��a<��a<�a<�a<�a<�a<-�a<?�a<Q�a<P�a<g�a<g�a<s�a<h�a<��a<n�a<x�a<x�a<d�a<f�a<i�a<\�a<V�a<?�a<(�a<#�a<�a<�a<�a<Ůa<��a<��a<��a<`�a<F�a<$�a<��a<ܭa<��a<��a<m�a<4�a<�a<۬a<��a<��a<S�a<�a<�a<��a<x�a<=�a<�a<êa<��a<@�a<�a<��a<{�a<)�a<ݨa<��a<T�a<�a<��a<Y�a<��a<��a<[�a<�a<��a<F�a<�a<��a<>�a<Уa<u�a<�a<��a<F�a<�a<��a<�a<��a<9�a<ҟa<r�a<�a<��a<*�a<��a<U�a<�a<��a<�a<��a<6�a<ۚa<k�a<��a<��a<*�a<̘a<r�a<�a<��a<F�a<�a<��a<4�a<̕a<��a<&�a<͔a<z�a<2�a<�a<��a<T�a<�a<Ēa<~�a<R�a<
�a<��a<��a<Q�a<)�a<�a<Ґa<��a<w�a<U�a<8�a<�a< �a<ߏa<Џa<��a<��a<��a<��a<��a<�a<��a<��a<��a<��a<��a<��a<͏a<�a<�a<�  �  +�a<�a<h�a<t�a<��a<̐a<�a<3�a<P�a<��a<��a<�a<G�a<|�a<�a< �a<^�a<��a<�a<H�a<��a<�a<4�a<��a<�a<S�a<��a<�a<��a<��a<M�a<��a<�a<n�a<ڙa<[�a<��a<?�a<��a<�a<u�a<�a<p�a<��a<X�a<��a<.�a<��a<�a<��a<�a<p�a<��a<G�a<��a<(�a<��a<�a<g�a<��a<>�a<��a<��a<f�a<��a<"�a<g�a<�a<!�a<��a<�a<"�a<��a<ũa<0�a<P�a<��a<�a<*�a<��a<��a<�a<�a<~�a<��a<جa<�a<-�a<r�a<��a<ϭa<�a<�a<9�a<D�a<|�a<��a<̮a<Ǯa<�a<��a< �a<0�a<&�a<K�a<I�a<V�a<b�a<a�a<��a<_�a<��a<j�a<}�a<~�a<m�a<x�a<P�a<o�a<?�a<J�a<5�a<&�a<�a<�a<��a<��a<ˮa<��a<|�a<f�a<?�a<0�a<��a<�a<��a<��a<m�a<8�a<3�a<جa<��a<y�a<T�a<)�a<�a<��a<r�a<H�a<��a<˪a<��a<<�a<�a<��a<��a<*�a<�a<��a<G�a<�a<��a<q�a<�a<Ʀa<W�a<�a<��a<=�a<	�a<��a<<�a<Уa<y�a<�a<��a<W�a<ˡa<��a<�a<��a<R�a<Οa<t�a<�a<��a<(�a<a<^�a<�a<��a<�a<��a<2�a<��a<t�a<��a<��a<-�a<�a<W�a<�a<��a<9�a<��a<��a<C�a<��a<��a<#�a<Ԕa<��a<$�a<�a<��a<]�a< �a<Ȓa<��a</�a<
�a<��a<��a<Y�a<(�a<��a<��a<��a<p�a<a�a<0�a<�a<��a<ُa<�a<��a<��a<��a<��a<��a<��a<��a<|�a<��a<��a<��a<��a<Ϗa<�a<�a<�  �  �a<6�a<K�a<q�a<��a<Ȑa<�a<+�a<g�a<��a<ˑa<�a<F�a<��a<��a<�a<U�a<��a<�a<=�a<��a<�a<8�a<��a<��a<>�a<��a<�a<s�a<ݗa<<�a<��a<
�a<{�a<�a<R�a<��a<*�a<��a< �a<x�a<�a<^�a<ѝa<4�a<��a<6�a<��a<�a<��a<��a<\�a<ӡa<?�a<��a<�a<��a<��a<_�a<ʤa<.�a<��a<�a<\�a<��a<&�a<��a<ŧa<,�a<��a<�a<,�a<u�a<ǩa<�a<d�a<��a<��a<<�a<{�a<��a<��a<7�a<p�a<��a<Ӭa<��a<I�a<o�a<��a<��a<��a<�a<7�a<S�a<u�a<��a<��a<ήa<�a<��a<�a<�a<;�a<G�a<G�a<W�a<s�a<g�a<f�a<z�a<v�a<}�a<w�a<k�a<q�a<l�a<^�a<c�a<I�a<C�a<4�a<�a<�a<�a<�a<Ӯa<��a<��a<��a<a�a<?�a<(�a<�a<֭a<��a<��a<l�a<E�a<�a<�a<��a<��a<X�a<�a<��a<��a<v�a<C�a<�a<��a<�a<B�a<�a<Ʃa<y�a<#�a<�a<��a<O�a<�a<��a<]�a<�a<��a<[�a<�a<��a<Q�a<�a<��a<D�a<ңa<t�a<�a<��a<C�a<�a<x�a<�a<��a<=�a<ڟa<l�a<�a<��a<.�a<ʝa<U�a<�a<��a<�a<��a<=�a<Қa<q�a<�a<��a</�a<Ϙa<k�a<�a<��a<K�a<�a<��a<.�a<ڕa<��a<#�a<Δa<r�a<?�a<�a<��a<N�a<�a<a<��a<?�a<�a<ϑa<��a<_�a<(�a<��a<͐a<��a<��a<]�a<.�a<�a<�a<ߏa<Ïa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<Ïa<�a<�a<�  �  �a<I�a<F�a<~�a<��a<��a<�a<�a<i�a<��a<Ցa<�a<;�a<��a<��a<�a<D�a<��a<�a<4�a<��a<Ӕa<S�a<��a<��a<A�a<��a<�a<a�a<��a<)�a<��a<��a<u�a<�a<A�a<͚a<�a<��a<�a<t�a<�a<T�a<�a<,�a<ʞa<�a<��a<�a<t�a<��a<P�a<�a<-�a<��a<�a<��a<�a<I�a<ڤa< �a<��a<�a<V�a<Ǧa<	�a<��a<��a<<�a<}�a<ըa<+�a<r�a<ߩa<�a<t�a<��a<��a<>�a<j�a<ͫa<�a<;�a<a�a<��a<٬a<��a<M�a<R�a<��a<��a<�a<�a<0�a<b�a<c�a<��a<��a<Үa<߮a<�a<�a<�a<>�a</�a<[�a<S�a<Y�a<u�a<^�a<��a<d�a<��a<k�a<z�a<s�a<Y�a<r�a<D�a<Y�a<6�a<1�a<-�a<�a<
�a<Ԯa<�a<��a<��a<��a<X�a<Y�a<�a<�a<έa<ŭa<��a<b�a<J�a<�a<��a<��a<��a<V�a<�a<�a<��a<��a<+�a<�a<��a<��a<N�a<�a<ɩa<f�a<?�a<٨a<��a<T�a<�a<��a<I�a<�a<��a<W�a<�a<��a<c�a<ݤa<��a<'�a<ڣa<t�a<�a<��a<7�a<��a<g�a<�a<��a<9�a<�a<W�a<�a<��a<+�a<��a<N�a<��a<k�a<(�a<��a<L�a<͚a<g�a<�a<��a<H�a<��a<{�a< �a<��a<M�a<ٖa<��a<�a<ޕa<s�a<,�a<Ԕa<r�a<C�a<̓a<��a<A�a<�a<��a<~�a<N�a<�a<ۑa<��a<d�a<&�a<�a<ِa<��a<��a<E�a<B�a<�a<�a<�a<��a<ҏa<��a<��a<��a<��a<��a<{�a<��a<��a<��a<��a<��a<׏a<ҏa<�a<�  �  �a</�a<S�a<��a<��a<Ða<��a<)�a<e�a<��a<��a<�a<G�a<��a<ђa<�a<X�a<��a<�a<=�a<��a<�a<A�a<��a<�a<\�a<��a<�a<x�a<ޗa<4�a<��a<	�a<t�a<�a<J�a<��a<*�a<��a<�a<{�a<��a<_�a<ɝa<I�a<a<�a<��a<�a<��a<�a<]�a<ǡa<A�a<��a<!�a<��a<��a<]�a<��a<'�a<��a<��a<X�a<��a<�a<��a<ݧa<(�a<��a<�a</�a<��a<ϩa<�a<i�a<��a<�a<7�a<y�a<��a<�a<9�a<u�a<��a<լa<�a<@�a<]�a<��a<��a<�a<�a<*�a<Q�a<v�a<��a<��a<ʮa<�a<��a<�a<"�a<<�a<C�a<M�a<S�a<T�a<y�a<r�a<q�a<v�a<��a<t�a<y�a<j�a<i�a<h�a<P�a<T�a<C�a<.�a<$�a<�a<	�a<�a<̮a<��a<��a<w�a<]�a<H�a<&�a<�a<�a<��a<��a<m�a<;�a<�a<�a<��a<��a<J�a<�a<�a<��a<�a<4�a<�a<Ԫa<��a<@�a<
�a<ǩa<p�a<0�a<�a<��a<P�a<��a<��a<\�a<	�a<��a<]�a<�a<��a<I�a<��a<��a<'�a<ѣa<n�a<�a<��a<C�a<ءa<{�a<�a<��a<D�a<֟a<j�a<��a<��a<+�a<ŝa<Q�a<�a<o�a<�a<��a<8�a<֚a<w�a<�a<��a<7�a<јa<q�a<�a<��a<F�a<�a<��a<*�a<ݕa<��a<'�a<єa<��a<6�a<֓a<��a<N�a<�a<��a<w�a<=�a<�a<Ǒa<��a<[�a</�a<��a<��a<��a<��a<Y�a<5�a<�a<�a<�a<Ϗa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<Ώa<ُa<�a<�  �   �a<,�a<X�a<q�a<��a<ܐa<�a<?�a<G�a<��a<ˑa<
�a<I�a<w�a<ܒa<��a<f�a<��a<��a<B�a<��a<��a<(�a<��a<�a<P�a<��a<�a<y�a<ʗa<K�a<��a<�a<s�a<�a<g�a<��a<1�a<��a<�a<�a<�a<l�a<ǝa<J�a<��a<5�a<��a<�a<��a<ݠa<t�a<ša<V�a<��a<�a<��a<�a<t�a<��a<B�a<��a<�a<b�a<��a<,�a<f�a<ۧa<&�a<��a<ڨa<-�a<��a<��a<#�a<\�a<êa<��a<3�a<��a<��a<�a<)�a<q�a<��a<Ԭa<�a<-�a<��a<��a<ԭa<�a<�a<B�a<O�a<��a<~�a<��a<®a<�a<�a<
�a<2�a<�a<W�a<C�a<d�a<f�a<_�a<x�a<n�a<��a<m�a<��a<r�a<f�a<r�a<T�a<w�a<C�a<F�a<.�a<�a<�a<�a<�a<ɮa<��a<��a<��a<v�a<4�a<;�a<�a<�a<��a<��a<o�a<2�a<(�a<Ҭa<Ǭa<��a<`�a<#�a<߫a<ɫa<f�a<X�a<��a<Ǫa<��a<B�a<�a<��a<��a< �a<�a<��a<O�a<�a<��a<d�a<��a<��a<a�a< �a<��a<G�a<��a<��a<D�a<ңa<r�a<!�a<��a<Z�a<աa<��a<�a<��a<E�a<a<��a<��a<��a<�a<ʝa<[�a<��a<��a<�a<��a<7�a<��a<k�a<�a<��a< �a<٘a<c�a<�a<��a<B�a<�a<w�a<@�a<͕a<��a<*�a<Дa<��a<#�a<��a<��a<b�a<�a<��a<��a<;�a<�a<��a<��a<S�a<'�a<�a<ɐa<��a<g�a<m�a<*�a<!�a<��a<׏a<ԏa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<Ïa<�a<�a<�  �  �a<2�a<R�a<~�a<��a<ΐa<�a<2�a<N�a<��a<ʑa<��a<A�a<��a<̒a<�a<Q�a<��a<�a<?�a<��a<�a</�a<��a<�a<S�a<��a<�a<n�a<Зa<6�a<��a<�a<u�a<יa<H�a<��a</�a<��a<�a<|�a<�a<c�a<ϝa<F�a<��a< �a<��a<�a<��a<�a<e�a<ša<9�a<��a<!�a<��a<��a<Y�a<��a<2�a<��a<��a<_�a<��a<�a<v�a<اa<+�a<��a<֨a<.�a<�a<٩a< �a<a�a<��a<�a<6�a<��a<ëa<��a</�a<j�a<��a<Ѭa<�a<8�a<i�a<��a<̭a<�a<�a<6�a<J�a<q�a<��a<��a<Ѯa<�a<�a<	�a<$�a<&�a<H�a<H�a<X�a<a�a<n�a<n�a<s�a<}�a<s�a<v�a<t�a<��a<p�a<V�a<X�a<B�a<F�a<A�a<#�a<�a<��a<�a<Ϯa<��a<��a<��a<h�a<<�a<.�a<��a<�a<��a<��a<h�a<G�a<�a<�a<��a<z�a<W�a< �a<�a<��a<m�a<B�a<��a<˪a<~�a<H�a< �a<��a<r�a<7�a<�a<��a<C�a<��a<��a<b�a<�a<��a<^�a<�a<��a<O�a<��a<��a<.�a<ͣa<t�a<�a<��a<L�a<աa<s�a<�a<��a<D�a<ڟa<f�a<��a<��a<$�a<��a<X�a<�a<w�a<�a<��a<<�a<֚a<h�a<�a<��a<A�a<טa<h�a<�a<��a<F�a<�a<��a<.�a<ӕa<|�a<+�a<͔a<��a<.�a<�a<��a<Z�a<�a<��a<��a<5�a<��a<ёa<��a<b�a<(�a<�a<Ȑa<��a<p�a<^�a</�a<�a<��a<�a<ʏa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ȏa<͏a<ߏa<��a<�  �  �a<7�a<C�a<��a<��a<Ӑa<��a<�a<i�a<��a<ϑa<�a<:�a<��a<��a<�a<E�a<��a<�a<B�a<��a<ٔa<K�a<��a<��a<N�a<��a<�a<f�a<�a<�a<��a<��a<x�a<�a<D�a<њa<�a<��a<��a<z�a<�a<X�a<Нa<5�a<��a<&�a<��a<�a<z�a<�a<T�a<�a<:�a<��a<
�a<r�a<��a<R�a<�a<!�a<��a<��a<Y�a<Ѧa<�a<��a<Ƨa<'�a<}�a<Ҩa<4�a<l�a<ԩa<�a<y�a<��a<��a<B�a<h�a<īa<�a<C�a<c�a<��a<̬a<�a<E�a<k�a<��a<��a<�a<�a<*�a<s�a<e�a<��a<��a<Ȯa<ޮa<�a<�a<�a<A�a<4�a<P�a<c�a<h�a<v�a<]�a<w�a<t�a<~�a<h�a<n�a<p�a<_�a<w�a<J�a<`�a<9�a<,�a<!�a<��a<�a<�a<Ԯa<��a<��a<��a<m�a<L�a<�a<�a<ۭa<��a<��a<`�a<A�a<��a<�a<��a<��a<N�a<#�a<�a<��a<��a<C�a<�a<ƪa<w�a<M�a<��a<̩a<\�a<8�a<ըa<��a<V�a<��a<ħa<I�a<�a<��a<]�a<�a<��a<O�a<�a<��a<5�a<�a<s�a<�a<��a<:�a<��a<t�a<�a<��a<)�a<۟a<`�a<�a<��a<;�a<��a<R�a<��a<{�a<�a<��a<8�a<̚a<d�a<�a<��a<<�a<��a<��a<�a<��a<R�a<֖a<��a<�a<�a<u�a<+�a<ǔa<{�a<;�a<�a<��a<E�a<
�a<ɒa<w�a<^�a<�a<ԑa<x�a<Z�a<%�a<�a<֐a<��a<��a<J�a<7�a<!�a<�a<�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ˏa<Ώa<�a<�  �  �a<<�a<Z�a<t�a<��a<ΐa<�a<(�a<]�a<��a<��a<�a<5�a<��a<ϒa<�a<D�a<��a<�a<C�a<��a<�a<5�a<��a<�a<Q�a<��a<�a<d�a<՗a<>�a<��a<�a<s�a<әa<?�a<��a<,�a<��a<�a<�a<ܜa<b�a<ߝa<N�a<��a<+�a<��a<�a<x�a<��a<X�a<ϡa<9�a<��a<(�a<��a<��a<U�a<Ťa<#�a<��a<�a<V�a<��a< �a<m�a<ߧa<:�a<��a<ʨa<3�a<��a<ةa<�a<e�a<��a<�a<9�a<{�a<ȫa<��a<9�a<_�a<��a<�a<�a<3�a<r�a<��a<��a<�a<�a<&�a<V�a<e�a<��a<��a<خa<׮a<��a<�a<!�a<5�a<A�a<H�a<Y�a<a�a<e�a<w�a<�a<w�a<m�a<{�a<~�a<x�a<i�a<a�a<F�a<J�a<>�a<9�a<.�a<�a<�a<�a<ٮa<��a<��a<|�a<g�a<?�a<%�a<�a<�a<��a<��a<[�a<N�a<�a<��a<��a<��a<F�a<$�a<�a<��a<s�a<H�a<��a<Ȫa<��a<Q�a<��a<��a<{�a<?�a<�a<��a<@�a<�a<��a<_�a<�a<��a<b�a<��a<��a<^�a<��a<��a<9�a<Уa<m�a<
�a<��a<?�a<�a<r�a<�a<��a<K�a<֟a<c�a<��a<��a<0�a<��a<O�a<�a<��a<�a<��a<K�a<ښa<[�a<	�a<��a<@�a<՘a<l�a<��a<��a<H�a<�a<��a<7�a<ܕa<q�a<4�a<��a<��a<)�a<�a<��a<N�a<�a<ƒa<t�a<B�a<�a<Ցa<��a<i�a<�a<��a<a<��a<~�a<W�a</�a<�a<��a<ݏa<ӏa<ďa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<؏a<�a<��a<�  �  "�a<2�a<^�a<y�a<ʐa<ϐa<��a<V�a<@�a<��a<Ցa<�a<=�a<��a<��a<�a<g�a<��a<�a<Z�a<��a<�a<0�a<��a<�a<Y�a<��a<#�a<��a<ٗa<7�a<��a<�a<��a<��a<w�a<��a<5�a<��a<��a<u�a<��a<l�a<��a<T�a<��a<T�a<��a<>�a<��a<��a<��a<ˡa<R�a<��a<�a<��a<�a<q�a<��a<Y�a<��a<�a<��a<��a<>�a<|�a<�a<�a<��a<�a<*�a<o�a<��a<(�a<\�a<֪a<�a<?�a<��a<��a<�a<0�a<z�a<��a<��a<�a<J�a<z�a<��a<��a<�a<"�a<K�a<W�a<��a<��a<��a<ݮa<׮a<�a<�a<D�a<�a<b�a<W�a<V�a<��a<k�a<�a<g�a<��a<��a<u�a<V�a<y�a<k�a<X�a<}�a<O�a<B�a<>�a<��a<�a<�a<�a<ͮa<��a<��a<��a<g�a<F�a<P�a<�a<��a<ía<��a<b�a<N�a<�a<�a<Ƭa<��a<e�a<9�a<ګa<�a<l�a<O�a<�a<Ϫa<w�a<X�a<�a<��a<r�a<�a<�a<��a<`�a<'�a<��a<g�a<��a<��a<W�a<�a<��a<4�a<�a<��a<b�a<ģa<��a<(�a<��a<u�a<ۡa<��a<
�a<��a<?�a<̟a<�a<��a<��a<8�a<ϝa<��a<ٜa<��a<�a<��a<�a<�a<t�a<�a<��a<)�a<��a<e�a<3�a<ėa<O�a<��a<}�a<'�a<Օa<��a<8�a<��a<��a<B�a<��a<��a<��a<�a<ؒa<��a<D�a<�a<ȑa<��a<q�a< �a<
�a<ΐa<Ȑa<g�a<{�a<A�a<�a<)�a<�a<ݏa<��a<��a<��a<��a<s�a<��a<��a<��a<��a<��a<��a<ȏa<��a<�a<
�a<�  �  �a<F�a<n�a<��a<��a<̐a<��a<-�a<U�a<��a<��a<�a<?�a<��a<Вa<�a<[�a<��a<ړa<M�a<��a<�a<>�a<��a<�a<b�a<��a<'�a<l�a<ڗa<I�a<ʘa<�a<z�a<ؙa<C�a<��a<.�a<��a<(�a<��a<�a<r�a<ٝa<V�a<��a<,�a<��a<�a<z�a<�a<X�a<ša<I�a<��a</�a<��a<��a<a�a<��a<#�a<��a<�a<c�a<��a<�a<o�a<�a<7�a<��a<ڨa<9�a<��a<�a<�a<a�a<��a<�a<9�a<��a<�a<�a<7�a<e�a<��a<�a<�a<3�a<h�a<��a<ía<�a<�a<�a<]�a<u�a<��a<��a<߮a<ܮa<	�a<��a<$�a<)�a<@�a<P�a<U�a<f�a<j�a<��a<��a<|�a<y�a<��a<��a<��a<f�a<e�a<P�a<N�a<<�a<M�a<E�a<"�a<��a<�a<�a<Ϯa<��a<��a<d�a<I�a<'�a<��a<�a<��a<��a<d�a<S�a<�a<�a<��a<��a<=�a<,�a<�a<��a<z�a<A�a<��a<تa<��a<]�a<��a<��a<��a<V�a<��a<��a<C�a<�a<��a<`�a<'�a<Ѧa<l�a<�a<��a<X�a<�a<��a<:�a<ǣa<|�a<�a<��a<>�a<աa<��a<�a<��a<U�a<ܟa<o�a<��a<��a<,�a<��a<]�a<ޜa<��a<
�a<��a<I�a<�a<m�a<�a<��a<V�a<֘a<j�a< �a<��a<J�a<��a<��a<=�a<ܕa<y�a<A�a<�a<��a<+�a<�a<��a<S�a<�a<˒a<l�a<K�a<�a<ϑa<��a<r�a<%�a<�a<��a<��a<u�a<X�a<:�a<�a< �a<�a<�a<ɏa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<֏a<�a<��a<��a<�  �  $�a<0�a<Q�a<��a<��a<Րa<�a<&�a<p�a<��a<őa< �a<G�a<��a<��a<�a<W�a<Óa<�a<[�a<��a<�a<Y�a<��a<�a<f�a<��a<
�a<v�a<��a<,�a<��a<��a<��a<�a<]�a<�a<�a<��a<��a<��a<��a<f�a<ŝa<E�a<Şa<'�a<��a<�a<��a<�a<`�a<�a<I�a<��a<�a<��a<�a<c�a<�a<-�a<��a<��a<]�a<Ԧa<�a<��a<اa< �a<��a<�a<7�a<g�a<ѩa<�a<��a<��a<�a<P�a<c�a<��a<�a<K�a<q�a<��a<Ǭa<�a<;�a<l�a<��a<��a<��a<*�a<,�a<w�a<s�a<��a<��a<Ȯa<�a<�a<�a<-�a<E�a<@�a<d�a<i�a<V�a<{�a<q�a<o�a<��a<��a<z�a<n�a<`�a<f�a<��a<\�a<t�a<D�a<�a<�a<
�a<�a<��a<ʮa<��a<��a<v�a<m�a<^�a<!�a<�a<�a<��a<��a<k�a<D�a<	�a<�a<��a<��a<L�a<:�a<��a<��a<��a<D�a<��a<ܪa<v�a<@�a<�a<ܩa<g�a<3�a<Ψa<��a<q�a<�a<էa<N�a<	�a<��a<e�a<�a<��a<D�a<��a<��a<5�a<�a<~�a<�a<��a<G�a<��a<��a< �a<��a<:�a<�a<q�a<"�a<��a<A�a<Ɲa<W�a<�a<~�a<#�a<��a<2�a<ޚa<z�a<�a<��a<:�a<��a<��a<�a<ėa<a�a<Ӗa<��a<�a<�a<��a<'�a<Ĕa<��a<3�a<�a<��a<J�a<�a<ߒa<{�a<e�a<�a<ّa<��a<\�a<1�a<�a<Ԑa<��a<��a<Y�a<N�a<)�a<�a<��a<Џa<��a<��a<��a<��a<��a<~�a<��a<��a<��a<Əa<��a<��a<ˏa<ޏa<�a<�  �  "�a<C�a<g�a<��a<��a<ϐa<�a<J�a<I�a<��a<̑a<��a<J�a<��a<�a< �a<`�a<��a<��a<B�a<��a<�a</�a<��a<�a<f�a<��a<)�a<y�a<�a<T�a<��a<�a<{�a<ۙa<O�a<��a<7�a<��a<�a<��a<�a<p�a<۝a<Z�a<��a<+�a<��a<�a<��a<�a<u�a<ȡa<9�a<��a<9�a<��a<��a<Y�a<��a<>�a<��a<�a<a�a<��a<�a<�a<�a<:�a<��a<�a<@�a<��a<�a<*�a<[�a<��a<�a<8�a<��a<ǫa<	�a<?�a<s�a<��a<�a<%�a<;�a<p�a<��a<ӭa<�a<�a<;�a<A�a<v�a<��a<Ȯa<�a<�a<�a<�a<2�a<�a<X�a<H�a<Z�a<`�a<v�a<��a<�a<��a<{�a<��a<w�a<��a<v�a<Q�a<Z�a<?�a<N�a<@�a<%�a</�a<�a<�a<ޮa<Ȯa<��a<~�a<g�a<;�a<D�a<�a<�a<��a<��a<n�a<Q�a<.�a<��a<��a<s�a<\�a<!�a<߫a<ϫa<k�a<I�a<�a<ܪa<��a<^�a<	�a<˩a<��a<:�a<��a<��a<G�a<��a<��a<i�a<!�a<��a<w�a<�a<��a<[�a<
�a<��a<9�a<Уa<u�a<�a<��a<\�a<ءa<s�a<�a<Ơa<Y�a<ߟa<g�a<��a<��a<!�a<ȝa<Z�a<ߜa<��a<�a<��a<L�a<�a<s�a<�a<��a<N�a<�a<c�a<�a<��a<I�a<��a<��a<D�a<�a<��a<C�a<�a<��a<3�a<�a<��a<c�a<�a<Ēa<��a<.�a<�a<ّa<��a<s�a<2�a<�a<͐a<��a<i�a<q�a<2�a<�a<��a<�a<�a<Ǐa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ʏa<яa<�a< �a<�  �  �a<>�a<e�a<r�a<��a<�a<��a<N�a<R�a<��a<Бa<�a<]�a<k�a<a<�a<��a<��a<�a<J�a<��a<�a<+�a<��a<�a<N�a<��a<�a<h�a<Ɨa<V�a<��a<�a<v�a<��a<k�a<��a<=�a<��a<�a<��a<לa<f�a<ѝa<L�a<��a<K�a<��a<�a<��a<�a<}�a<ȡa<i�a<��a<�a<��a<�a<��a<��a<J�a<��a<�a<]�a<æa<C�a<h�a<٧a<-�a<��a<ƨa<1�a<��a<��a<-�a<\�a<ªa<��a<3�a<��a<��a<�a<*�a<^�a<��a<۬a<	�a<+�a<��a<��a<ҭa<�a<�a<G�a<U�a<��a<s�a<��a<��a<�a<�a<�a<5�a<%�a<`�a<6�a<s�a<v�a<]�a<~�a<x�a<|�a<f�a<��a<r�a<n�a<v�a<\�a<��a<E�a<F�a<3�a<�a<'�a<�a<�a<ٮa<Ʈa<��a<��a<��a<+�a<H�a<��a<�a<��a<��a<��a<%�a<�a<Ĭa<�a<��a<d�a<)�a<�a<Ϋa<g�a<i�a<��a<Īa<��a<Q�a<��a<��a<��a<�a<�a<��a<K�a<�a<��a<o�a<��a<��a<j�a<�a<��a<P�a<��a<��a<Y�a<�a<n�a<&�a<��a<c�a<ءa<��a<
�a<��a<8�a<ȟa<��a<��a<��a<#�a<̝a<V�a<�a<��a<�a<��a<?�a<ښa<Y�a<�a<��a<%�a<�a<d�a<�a<��a<D�a<��a<{�a<K�a<ϕa<r�a<3�a<ٔa<��a<#�a<�a<��a<b�a<�a<ǒa<��a<C�a<.�a<��a<��a<I�a<7�a<�a<ΐa<��a<q�a<y�a<�a<2�a<�a<׏a<ݏa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ɏa<��a<�a<�  �  &�a<4�a<S�a<��a<��a<ېa<�a<�a<l�a<��a<��a<�a<I�a<��a<�a<�a<^�a<��a<�a<T�a<��a<ؔa<Q�a<��a<�a<d�a<��a<�a<��a<�a<6�a<��a<�a<��a<�a<;�a<ɚa<8�a<��a<�a<w�a<��a<d�a<ҝa<P�a<Þa<!�a<��a<�a<��a<�a<h�a<ǡa<E�a<��a<'�a<��a<�a<e�a<��a<4�a<��a<��a<R�a<Цa<�a<��a<�a<,�a<��a<�a<0�a<x�a<ةa<'�a<r�a<��a<��a<G�a<��a<«a<�a<C�a<}�a<��a<Ѭa<�a<>�a<k�a<��a<��a<��a<#�a<-�a<N�a<{�a<��a<̮a<Ѯa<�a<��a<�a<!�a<@�a<8�a<S�a<l�a<`�a<�a<n�a<u�a<��a<��a<e�a<~�a<y�a<t�a<r�a<:�a<]�a<L�a<6�a<.�a<�a<�a<��a<Ϯa<��a<��a<|�a<r�a<Q�a<�a<�a<�a<��a<��a<m�a<G�a<2�a<�a<��a<��a<G�a<4�a<��a<��a<��a<C�a<�a<ڪa<��a<F�a<�a<Щa<q�a<7�a<�a<��a<X�a<�a<��a<j�a<�a<��a<X�a<�a<��a<Q�a< �a<��a</�a<�a<r�a<�a<��a<O�a<סa<�a<�a<��a<Q�a<�a<s�a<��a<��a<>�a<Ýa<L�a<��a<z�a<�a<��a<>�a<ؚa<}�a<�a<��a<B�a<ޘa<z�a< �a<��a<X�a<��a<��a<*�a<�a<��a<*�a<ϔa<��a<6�a<�a<��a<@�a<�a<ْa<|�a<<�a<�a<ؑa<��a<e�a<-�a<�a<Ða<��a<��a<P�a<=�a<+�a<��a<��a<͏a<��a<��a<��a<��a<��a<��a<��a<��a<x�a<��a<��a<��a<ڏa<ԏa<�a<�  �  ��a<Y�a<Q�a<��a<��a<ːa<�a<�a<n�a<��a<��a<�a<<�a<��a<��a<+�a<F�a<��a<
�a<=�a<��a<Քa<d�a<��a<�a<Q�a<��a<,�a<c�a<��a<7�a<Ҙa<�a<u�a<�a<B�a<Кa<�a<��a<�a<��a<��a<S�a<��a<3�a<ƞa<�a<��a<�a<y�a<��a<_�a<��a<1�a<��a<$�a<��a<�a<I�a<�a<1�a<��a<��a<c�a<ۦa<�a<��a<§a<N�a<��a<�a<8�a<��a<�a<�a<u�a<��a<��a<A�a<l�a<�a<��a<=�a<a�a<��a<�a<�a<N�a<Z�a<��a<��a<��a<�a<B�a<s�a<]�a<��a<��a<ܮa<ޮa<��a<=�a<�a<=�a</�a<m�a<`�a<e�a<~�a<f�a<��a<c�a<��a<p�a<��a<��a<[�a<��a<G�a<j�a<5�a<8�a<H�a<�a<�a<Ϯa<��a<��a<��a<��a<c�a<i�a<�a<�a<حa<�a<��a<`�a<Y�a<�a<�a<��a<��a<m�a<�a<��a<��a<��a<4�a<�a<Ǫa<��a<b�a<�a<ǩa<s�a<^�a<�a<��a<\�a<�a<§a<C�a<'�a<��a<d�a<�a<��a<t�a<�a<��a<-�a<�a<��a<�a<��a<E�a<
�a<j�a<�a<��a<>�a<�a<W�a<)�a<��a<7�a<Ýa<\�a<�a<o�a<%�a<��a<`�a<֚a<s�a<�a<��a<\�a<��a<~�a<�a<��a<R�a<ܖa<��a<.�a<�a<u�a<<�a<�a<~�a<F�a<֓a<��a<B�a<�a<ǒa<��a<`�a<�a<��a<��a<p�a<&�a<��a<��a<��a<��a<G�a<W�a< �a< �a<��a<ŏa<�a<��a<��a<��a<��a<��a<�a<��a<��a<��a<��a<a<�a<ڏa<�a<�  �  �a<D�a<b�a<u�a<��a<Ȑa<��a<<�a<s�a<��a<ؑa<	�a<T�a<��a<��a< �a<c�a<��a<��a<1�a<��a<��a<?�a<��a<�a<M�a<Ėa<�a<m�a<�a<>�a<��a<�a<z�a<�a<h�a<̚a<3�a<��a<�a<��a<��a<O�a<�a<D�a<��a<9�a<��a<�a<��a<��a<Y�a<١a<L�a<��a<�a<��a<�a<j�a<Ѥa<'�a<��a<�a<]�a<��a<(�a<��a<Чa<B�a<y�a<ިa<A�a<��a<ǩa<"�a<t�a<��a<��a<<�a<}�a<��a<��a<C�a<k�a<��a<�a<�a<I�a<r�a<��a<ȭa<��a<�a<2�a<a�a<��a<��a<��a<֮a<��a<��a<�a<�a<E�a<T�a<N�a<S�a<x�a<f�a<v�a<��a<g�a<��a<��a<e�a<l�a<p�a<i�a<x�a<T�a<E�a</�a<�a<�a<�a<خa<߮a<îa<��a<��a<`�a<E�a<6�a<�a<ӭa<ƭa<��a<y�a<N�a<��a<��a<¬a<��a<\�a<�a< �a<«a<{�a<@�a<�a<êa<��a<I�a<��a<̩a<z�a<#�a<�a<��a<T�a<�a<��a<e�a<�a<��a<s�a<�a<��a<e�a<��a<��a<F�a<Уa<u�a<!�a<��a<@�a<�a<��a<!�a<��a<:�a<�a<x�a<�a<��a<3�a<Нa<V�a<�a<��a<�a<��a<T�a<ʚa<q�a<�a<��a<0�a<ژa<}�a<�a<��a<M�a<�a<��a<8�a<�a<�a<*�a<�a<|�a<A�a<�a<��a<X�a<�a<��a<��a<N�a<�a<ّa<|�a<j�a<?�a<�a<אa<��a<��a<l�a<8�a<�a<�a<�a<Տa<͏a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<�a<�a<�  �  9�a<�a<{�a<�a<��a<ېa<�a<(�a<H�a<��a<đa<�a<I�a<}�a<�a<
�a<g�a<��a<�a<T�a<��a<�a<>�a<��a<�a<f�a<Ɩa<��a<��a<ʗa<R�a<��a<-�a<~�a<ϙa<I�a<��a<S�a<��a<�a<z�a<�a<m�a<ʝa<q�a<��a<)�a<��a<�a<o�a<�a<y�a<��a<T�a<��a<&�a<��a<�a<r�a<��a<=�a<��a<�a<_�a<��a<�a<i�a<��a</�a<��a<�a<&�a<��a<ũa<C�a<Q�a<��a<�a<4�a<��a<��a<�a<%�a<��a<��a<�a<'�a<+�a<r�a<��a<ȭa<ӭa<�a<7�a<J�a<��a<��a<Ϯa<Ůa<�a<�a<��a<;�a<�a<8�a<[�a<e�a<`�a<e�a<��a<_�a<��a<p�a<��a<��a<y�a<��a<?�a<R�a<-�a<]�a<A�a<(�a<"�a<�a<	�a<��a<ܮa<��a<{�a<r�a<O�a<#�a<�a<��a<��a<��a<n�a<7�a<<�a<�a<Ƭa<��a<T�a<3�a<٫a<��a<z�a<L�a<��a<ܪa<��a<1�a<!�a<��a<��a<,�a<�a<��a<;�a<��a<��a<��a<�a<Ȧa<\�a<�a<��a<J�a<!�a<��a<7�a<֣a<|�a<�a<��a<`�a<ϡa<��a<�a<��a<R�a<Οa<��a<�a<��a<,�a<��a<Y�a<�a<��a<�a<ӛa<A�a<ۚa<s�a<��a<��a<.�a<��a<Z�a<�a<��a<E�a<�a<��a<K�a<ʕa<��a<�a<�a<��a<#�a<�a<��a<X�a<�a<Ԓa<��a<8�a<�a<Ǒa<��a<Y�a<.�a<�a<��a<��a<j�a<Q�a<D�a<%�a<��a<ߏa<��a<��a<̏a<��a<��a<��a<��a<��a<n�a<��a<��a<ɏa<ˏa<ԏa<��a<�a<�  �  8�a<(�a<[�a<x�a<��a<ݐa<�a<4�a<e�a<��a<ёa<�a<S�a<z�a<˒a<��a<c�a<��a<��a<a�a<��a<�a<I�a<��a<��a<O�a<��a<�a<��a<ėa<P�a<��a<��a<��a<��a<f�a<ɚa<)�a<��a<�a<y�a<�a<m�a<Ýa<H�a<��a<D�a<��a<&�a<��a<��a<q�a<�a<R�a<��a<�a<��a<�a<p�a<ݤa<:�a<��a< �a<r�a<˦a<5�a<~�a<اa< �a<��a<ިa<%�a<��a<��a<�a<m�a<Ūa<�a<A�a<p�a<��a<�a<#�a<{�a<��a<լa<�a<D�a<��a<��a<ϭa<�a<+�a<7�a<l�a<��a<��a<��a<îa<�a<�a<�a<=�a<?�a<F�a<f�a<i�a<w�a<i�a<y�a<f�a<��a<i�a<z�a<|�a<\�a<q�a<r�a<s�a<]�a<E�a<�a<$�a<�a<�a<�a<îa<��a<��a<��a<t�a<V�a<.�a<
�a<��a<��a<��a<w�a<3�a<�a<լa<¬a<��a<W�a<@�a<�a<��a<��a<Z�a<�a<Ūa<��a<B�a<�a<��a<��a<+�a<רa<��a<d�a<�a<��a<Z�a<��a<��a<[�a<�a<��a<B�a<��a<��a<R�a<�a<��a<�a<��a<X�a<�a<��a<�a<��a<=�a<Οa<}�a<�a<��a<<�a<ǝa<k�a<��a<��a<�a<��a<2�a<ܚa<q�a<��a<��a<&�a<͘a<v�a<"�a<ėa<R�a<��a<��a<G�a<ȕa<��a<)�a<Ӕa<��a<<�a<��a<��a<_�a<
�a<�a<��a<Y�a<�a<��a<��a<W�a<3�a<	�a<ِa<��a<��a<^�a<O�a<(�a<�a<�a<؏a<��a<̏a<��a<��a<��a<z�a<��a<��a<��a<��a<��a<��a<Џa<�a<�a<�  �  �a<N�a<^�a<o�a<��a<Őa<��a<7�a<s�a<��a<ʑa<�a<O�a<��a<Вa<;�a<P�a<��a<�a<G�a<��a<�a<8�a<��a< �a<D�a<��a<$�a<s�a<�a<F�a<��a<�a<�a<ޙa<?�a<˚a<+�a<��a<�a<��a<��a<Y�a<�a<E�a<��a<3�a<��a<�a<��a<�a<I�a<ԡa<)�a<Ȣa<5�a<��a<�a<J�a<ˤa<�a<��a<�a<c�a<��a<!�a<��a<ԧa<F�a<��a<�a<C�a<|�a<�a<�a<u�a<��a<�a<D�a<��a<˫a<��a<F�a<l�a<��a<�a<�a<J�a<j�a<��a<ƭa<��a<�a<!�a<Q�a<h�a<��a<��a<�a<��a<�a<�a<�a<O�a<D�a<H�a<L�a<{�a<a�a<u�a<��a<p�a<��a<��a<k�a<��a<i�a<j�a<O�a<T�a<A�a<L�a<�a<#�a<�a<�a<�a<��a<��a<��a<\�a<@�a<1�a<�a<խa<��a<}�a<t�a<f�a<�a<�a<��a<{�a<K�a<&�a<��a<��a<t�a<A�a<�a<��a<��a<Z�a<�a<ѩa<��a<9�a<��a<��a<I�a<�a<��a<\�a<,�a<��a<x�a<�a<��a<k�a<��a<��a<@�a<ƣa<u�a<�a<��a<0�a<�a<c�a<,�a< a<V�a<��a<X�a<�a<��a<8�a<̝a<\�a<ۜa<��a<�a<��a<X�a<՚a<u�a<�a<��a<Y�a<՘a<~�a<�a<��a<U�a<��a<��a<4�a<�a<��a<8�a<�a<��a<B�a<�a<��a<V�a<�a<̒a<p�a<>�a<��a<��a<��a<��a<>�a<�a<ѐa<��a<��a<]�a<2�a<�a<�a<ۏa<ԏa<׏a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<Տa<ŏa<��a<�a<�  �  �a<8�a<X�a<{�a<��a<��a<�a<+�a<`�a<��a<�a<!�a<C�a<��a<��a<�a<X�a<��a<�a<T�a<��a<�a<I�a<��a<�a<R�a<��a<�a<q�a<ϗa<<�a<��a<�a<r�a<��a<[�a<��a<*�a<��a<��a<�a<�a<c�a<͝a<C�a<��a<;�a<��a<&�a<z�a<��a<q�a<��a<K�a<��a<�a<~�a<�a<d�a<�a<E�a<��a<��a<v�a<Ȧa</�a<o�a<ԧa<%�a<��a<Ҩa<,�a<p�a<ɩa<�a<j�a<��a<�a<<�a<��a<��a<�a<1�a<g�a<��a<ʬa<�a<5�a<}�a<��a<Эa<�a<�a<R�a<s�a<x�a<��a<��a<��a<�a<�a<3�a<.�a<5�a<;�a<e�a<i�a<t�a<g�a<r�a<w�a<|�a<r�a<��a<]�a<��a<m�a<m�a<_�a<^�a<=�a<D�a<�a<�a<��a<�a<Ӯa<��a<��a<��a<x�a<X�a<&�a<�a<�a<ݭa<��a<h�a<<�a<
�a<�a<��a<��a<w�a<3�a<�a<��a<��a<W�a< �a<Ȫa<~�a<I�a<�a<��a<w�a<�a<��a<��a<`�a<�a<��a<[�a<�a<��a<`�a<��a<��a<L�a<�a<��a<I�a<�a<��a<�a<��a<W�a<�a<��a<�a<��a<6�a<ӟa<r�a<!�a<��a<5�a<��a<p�a<��a<��a<�a<��a<7�a<ݚa<d�a<�a<��a<3�a<јa<r�a<�a<��a<M�a<��a<~�a<*�a<֕a<{�a<1�a<Ȕa<��a<.�a<��a<��a<`�a<�a<Ӓa<��a<a�a<�a<ɑa<��a<T�a<.�a<�a<��a<��a<��a<T�a<O�a<)�a<�a<�a<яa<��a<��a<��a<��a<z�a<��a<��a<��a<��a<��a<��a<Ώa<��a<�a<�a<�  �  F�a<1�a<\�a<��a<��a<ΐa<��a<5�a<k�a<��a<��a<�a<J�a<��a<�a< �a<\�a<��a<Փa<?�a<��a<��a<.�a<��a<��a<|�a<��a<"�a<��a<ȗa<b�a<��a<�a<j�a<�a<Q�a<��a<?�a<��a<)�a<��a<�a<��a<a<V�a<��a<2�a<�a<�a<��a<�a<W�a<¡a<M�a<��a<=�a<��a<�a<l�a<��a<"�a<��a<�a<f�a<��a<)�a<|�a<�a<�a<��a<�a<;�a<��a<ȩa<+�a<[�a<��a<��a</�a<��a<��a<#�a<3�a<��a<ʬa<ʬa<8�a<A�a<{�a<|�a<έa<��a<	�a<�a<N�a<}�a<��a<ٮa<خa<�a<�a<�a< �a<:�a<P�a<^�a<O�a<k�a<��a<|�a<g�a<��a<d�a<��a<��a<x�a<r�a<d�a<N�a<W�a<<�a<<�a<,�a<+�a<�a<�a<̮a<��a<®a<��a<f�a<H�a<0�a<�a<�a<��a<��a<o�a<F�a<9�a<׬a<��a<��a<8�a<�a<��a<��a<j�a<Q�a<�a<�a<��a<W�a< �a<��a<��a<)�a<�a<��a<]�a<�a<��a<q�a<�a<Ҧa<n�a<�a<ߥa<A�a<�a<��a<@�a<��a<~�a<�a<��a<=�a<ҡa<��a<�a<ʠa<h�a<џa<z�a<�a<��a<)�a<ɝa<_�a<ʜa<��a<�a<ƛa</�a<�a<w�a<�a<řa<1�a<�a<d�a<
�a<��a<@�a<��a<��a<]�a<ٕa<��a<Q�a<Ȕa<��a<9�a<��a<�a<^�a<�a<��a<i�a<<�a<�a<��a<��a<l�a<5�a<�a<��a<��a<��a<i�a<G�a<�a<�a<�a<ۏa<��a<�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<Əa<؏a<��a<�a<�  �  �a<8�a<X�a<{�a<��a<��a<�a<+�a<`�a<��a<�a<!�a<C�a<��a<��a<�a<X�a<��a<�a<T�a<��a<�a<I�a<��a<�a<R�a<��a<�a<q�a<ϗa<<�a<��a<�a<r�a<��a<[�a<��a<*�a<��a<��a<�a<�a<c�a<͝a<C�a<��a<;�a<��a<&�a<z�a<��a<q�a<��a<K�a<��a<�a<~�a<�a<d�a<�a<E�a<��a<��a<v�a<Ȧa</�a<o�a<ԧa<%�a<��a<Ҩa<,�a<p�a<ɩa<�a<j�a<��a<�a<<�a<��a<��a<�a<1�a<g�a<��a<ʬa<�a<5�a<}�a<��a<Эa<�a<�a<R�a<s�a<x�a<��a<��a<��a<�a<�a<3�a<.�a<5�a<;�a<e�a<i�a<t�a<g�a<r�a<w�a<|�a<r�a<��a<]�a<��a<m�a<m�a<_�a<^�a<=�a<D�a<�a<�a<��a<�a<Ӯa<��a<��a<��a<x�a<X�a<&�a<�a<�a<ݭa<��a<h�a<<�a<
�a<�a<��a<��a<w�a<3�a<�a<��a<��a<W�a< �a<Ȫa<~�a<I�a<�a<��a<w�a<�a<��a<��a<`�a<�a<��a<[�a<�a<��a<`�a<��a<��a<L�a<�a<��a<I�a<�a<��a<�a<��a<W�a<�a<��a<�a<��a<6�a<ӟa<r�a<!�a<��a<5�a<��a<p�a<��a<��a<�a<��a<7�a<ݚa<d�a<�a<��a<3�a<јa<r�a<�a<��a<M�a<��a<~�a<*�a<֕a<{�a<1�a<Ȕa<��a<.�a<��a<��a<`�a<�a<Ӓa<��a<a�a<�a<ɑa<��a<T�a<.�a<�a<��a<��a<��a<T�a<O�a<)�a<�a<�a<яa<��a<��a<��a<��a<z�a<��a<��a<��a<��a<��a<��a<Ώa<��a<�a<�a<�  �  �a<N�a<^�a<o�a<��a<Őa<��a<7�a<s�a<��a<ʑa<�a<O�a<��a<Вa<;�a<P�a<��a<�a<G�a<��a<�a<8�a<��a< �a<D�a<��a<$�a<s�a<�a<F�a<��a<�a<�a<ޙa<?�a<˚a<+�a<��a<�a<��a<��a<Y�a<�a<E�a<��a<3�a<��a<�a<��a<�a<I�a<ԡa<)�a<Ȣa<5�a<��a<�a<J�a<ˤa<�a<��a<�a<c�a<��a<!�a<��a<ԧa<F�a<��a<�a<C�a<|�a<�a<�a<u�a<��a<�a<D�a<��a<˫a<��a<F�a<l�a<��a<�a<�a<J�a<j�a<��a<ƭa<��a<�a<!�a<Q�a<h�a<��a<��a<�a<��a<�a<�a<�a<O�a<D�a<H�a<L�a<{�a<a�a<u�a<��a<p�a<��a<��a<k�a<��a<i�a<j�a<O�a<T�a<A�a<L�a<�a<#�a<�a<�a<�a<��a<��a<��a<\�a<@�a<1�a<�a<խa<��a<}�a<t�a<f�a<�a<�a<��a<{�a<K�a<&�a<��a<��a<t�a<A�a<�a<��a<��a<Z�a<�a<ѩa<��a<9�a<��a<��a<I�a<�a<��a<\�a<,�a<��a<x�a<�a<��a<k�a<��a<��a<@�a<ƣa<u�a<�a<��a<0�a<�a<c�a<,�a< a<V�a<��a<X�a<�a<��a<8�a<̝a<\�a<ۜa<��a<�a<��a<X�a<՚a<u�a<�a<��a<Y�a<՘a<~�a<�a<��a<U�a<��a<��a<4�a<�a<��a<8�a<�a<��a<B�a<�a<��a<V�a<�a<̒a<p�a<>�a<��a<��a<��a<��a<>�a<�a<ѐa<��a<��a<]�a<2�a<�a<�a<ۏa<ԏa<׏a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<Տa<ŏa<��a<�a<�  �  8�a<(�a<[�a<x�a<��a<ݐa<�a<4�a<e�a<��a<ёa<�a<S�a<z�a<˒a<��a<c�a<��a<��a<a�a<��a<�a<I�a<��a<��a<O�a<��a<�a<��a<ėa<P�a<��a<��a<��a<��a<f�a<ɚa<)�a<��a<�a<y�a<�a<m�a<Ýa<H�a<��a<D�a<��a<&�a<��a<��a<q�a<�a<R�a<��a<�a<��a<�a<p�a<ݤa<:�a<��a< �a<r�a<˦a<5�a<~�a<اa< �a<��a<ިa<%�a<��a<��a<�a<m�a<Ūa<�a<A�a<p�a<��a<�a<#�a<{�a<��a<լa<�a<D�a<��a<��a<ϭa<�a<+�a<7�a<l�a<��a<��a<��a<îa<�a<�a<�a<=�a<?�a<F�a<f�a<i�a<w�a<i�a<y�a<f�a<��a<i�a<z�a<|�a<\�a<q�a<r�a<s�a<]�a<E�a<�a<$�a<�a<�a<�a<îa<��a<��a<��a<t�a<V�a<.�a<
�a<��a<��a<��a<w�a<3�a<�a<լa<¬a<��a<W�a<@�a<�a<��a<��a<Z�a<�a<Ūa<��a<B�a<�a<��a<��a<+�a<רa<��a<d�a<�a<��a<Z�a<��a<��a<[�a<�a<��a<B�a<��a<��a<R�a<�a<��a<�a<��a<X�a<�a<��a<�a<��a<=�a<Οa<}�a<�a<��a<<�a<ǝa<k�a<��a<��a<�a<��a<2�a<ܚa<q�a<��a<��a<&�a<͘a<v�a<"�a<ėa<R�a<��a<��a<G�a<ȕa<��a<)�a<Ӕa<��a<<�a<��a<��a<_�a<
�a<�a<��a<Y�a<�a<��a<��a<W�a<3�a<	�a<ِa<��a<��a<^�a<O�a<(�a<�a<�a<؏a<��a<̏a<��a<��a<��a<z�a<��a<��a<��a<��a<��a<��a<Џa<�a<�a<�  �  9�a<�a<{�a<�a<��a<ېa<�a<(�a<H�a<��a<đa<�a<I�a<}�a<�a<
�a<g�a<��a<�a<T�a<��a<�a<>�a<��a<�a<f�a<Ɩa<��a<��a<ʗa<R�a<��a<-�a<~�a<ϙa<I�a<��a<S�a<��a<�a<z�a<�a<m�a<ʝa<q�a<��a<)�a<��a<�a<o�a<�a<y�a<��a<T�a<��a<&�a<��a<�a<r�a<��a<=�a<��a<�a<_�a<��a<�a<i�a<��a</�a<��a<�a<&�a<��a<ũa<C�a<Q�a<��a<�a<4�a<��a<��a<�a<%�a<��a<��a<�a<'�a<+�a<r�a<��a<ȭa<ӭa<�a<7�a<J�a<��a<��a<Ϯa<Ůa<�a<�a<��a<;�a<�a<8�a<[�a<e�a<`�a<e�a<��a<_�a<��a<p�a<��a<��a<y�a<��a<?�a<R�a<-�a<]�a<A�a<(�a<"�a<�a<	�a<��a<ܮa<��a<{�a<r�a<O�a<#�a<�a<��a<��a<��a<n�a<7�a<<�a<�a<Ƭa<��a<T�a<3�a<٫a<��a<z�a<L�a<��a<ܪa<��a<1�a<!�a<��a<��a<,�a<�a<��a<;�a<��a<��a<��a<�a<Ȧa<\�a<�a<��a<J�a<!�a<��a<7�a<֣a<|�a<�a<��a<`�a<ϡa<��a<�a<��a<R�a<Οa<��a<�a<��a<,�a<��a<Y�a<�a<��a<�a<ӛa<A�a<ۚa<s�a<��a<��a<.�a<��a<Z�a<�a<��a<E�a<�a<��a<K�a<ʕa<��a<�a<�a<��a<#�a<�a<��a<X�a<�a<Ԓa<��a<8�a<�a<Ǒa<��a<Y�a<.�a<�a<��a<��a<j�a<Q�a<D�a<%�a<��a<ߏa<��a<��a<̏a<��a<��a<��a<��a<��a<n�a<��a<��a<ɏa<ˏa<ԏa<��a<�a<�  �  �a<D�a<b�a<u�a<��a<Ȑa<��a<<�a<s�a<��a<ؑa<	�a<T�a<��a<��a< �a<c�a<��a<��a<1�a<��a<��a<?�a<��a<�a<M�a<Ėa<�a<m�a<�a<>�a<��a<�a<z�a<�a<h�a<̚a<3�a<��a<�a<��a<��a<O�a<�a<D�a<��a<9�a<��a<�a<��a<��a<Y�a<١a<L�a<��a<�a<��a<�a<j�a<Ѥa<'�a<��a<�a<]�a<��a<(�a<��a<Чa<B�a<y�a<ިa<A�a<��a<ǩa<"�a<t�a<��a<��a<<�a<}�a<��a<��a<C�a<k�a<��a<�a<�a<I�a<r�a<��a<ȭa<��a<�a<2�a<a�a<��a<��a<��a<֮a<��a<��a<�a<�a<E�a<T�a<N�a<S�a<x�a<f�a<v�a<��a<g�a<��a<��a<e�a<l�a<p�a<i�a<x�a<T�a<E�a</�a<�a<�a<�a<خa<߮a<îa<��a<��a<`�a<E�a<6�a<�a<ӭa<ƭa<��a<y�a<N�a<��a<��a<¬a<��a<\�a<�a< �a<«a<{�a<@�a<�a<êa<��a<I�a<��a<̩a<z�a<#�a<�a<��a<T�a<�a<��a<e�a<�a<��a<s�a<�a<��a<e�a<��a<��a<F�a<Уa<u�a<!�a<��a<@�a<�a<��a<!�a<��a<:�a<�a<x�a<�a<��a<3�a<Нa<V�a<�a<��a<�a<��a<T�a<ʚa<q�a<�a<��a<0�a<ژa<}�a<�a<��a<M�a<�a<��a<8�a<�a<�a<*�a<�a<|�a<A�a<�a<��a<X�a<�a<��a<��a<N�a<�a<ّa<|�a<j�a<?�a<�a<אa<��a<��a<l�a<8�a<�a<�a<�a<Տa<͏a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<�a<�a<�  �  ��a<Y�a<Q�a<��a<��a<ːa<�a<�a<n�a<��a<��a<�a<<�a<��a<��a<+�a<F�a<��a<
�a<=�a<��a<Քa<d�a<��a<�a<Q�a<��a<,�a<c�a<��a<7�a<Ҙa<�a<u�a<�a<B�a<Кa<�a<��a<�a<��a<��a<S�a<��a<3�a<ƞa<�a<��a<�a<y�a<��a<_�a<��a<1�a<��a<$�a<��a<�a<I�a<�a<1�a<��a<��a<c�a<ۦa<�a<��a<§a<N�a<��a<�a<8�a<��a<�a<�a<u�a<��a<��a<A�a<l�a<�a<��a<=�a<a�a<��a<�a<�a<N�a<Z�a<��a<��a<��a<�a<B�a<s�a<]�a<��a<��a<ܮa<ޮa<��a<=�a<�a<=�a</�a<m�a<`�a<e�a<~�a<f�a<��a<c�a<��a<p�a<��a<��a<[�a<��a<G�a<j�a<5�a<8�a<H�a<�a<�a<Ϯa<��a<��a<��a<��a<c�a<i�a<�a<�a<حa<�a<��a<`�a<Y�a<�a<�a<��a<��a<m�a<�a<��a<��a<��a<4�a<�a<Ǫa<��a<b�a<�a<ǩa<s�a<^�a<�a<��a<\�a<�a<§a<C�a<'�a<��a<d�a<�a<��a<t�a<�a<��a<-�a<�a<��a<�a<��a<E�a<
�a<j�a<�a<��a<>�a<�a<W�a<)�a<��a<7�a<Ýa<\�a<�a<o�a<%�a<��a<`�a<֚a<s�a<�a<��a<\�a<��a<~�a<�a<��a<R�a<ܖa<��a<.�a<�a<u�a<<�a<�a<~�a<F�a<֓a<��a<B�a<�a<ǒa<��a<`�a<�a<��a<��a<p�a<&�a<��a<��a<��a<��a<G�a<W�a< �a< �a<��a<ŏa<�a<��a<��a<��a<��a<��a<�a<��a<��a<��a<��a<a<�a<ڏa<�a<�  �  &�a<4�a<S�a<��a<��a<ېa<�a<�a<l�a<��a<��a<�a<I�a<��a<�a<�a<^�a<��a<�a<T�a<��a<ؔa<Q�a<��a<�a<d�a<��a<�a<��a<�a<6�a<��a<�a<��a<�a<;�a<ɚa<8�a<��a<�a<w�a<��a<d�a<ҝa<P�a<Þa<!�a<��a<�a<��a<�a<h�a<ǡa<E�a<��a<'�a<��a<�a<e�a<��a<4�a<��a<��a<R�a<Цa<�a<��a<�a<,�a<��a<�a<0�a<x�a<ةa<'�a<r�a<��a<��a<G�a<��a<«a<�a<C�a<}�a<��a<Ѭa<�a<>�a<k�a<��a<��a<��a<#�a<-�a<N�a<{�a<��a<̮a<Ѯa<�a<��a<�a<!�a<@�a<8�a<S�a<l�a<`�a<�a<n�a<u�a<��a<��a<e�a<~�a<y�a<t�a<r�a<:�a<]�a<L�a<6�a<.�a<�a<�a<��a<Ϯa<��a<��a<|�a<r�a<Q�a<�a<�a<�a<��a<��a<m�a<G�a<2�a<�a<��a<��a<G�a<4�a<��a<��a<��a<C�a<�a<ڪa<��a<F�a<�a<Щa<q�a<7�a<�a<��a<X�a<�a<��a<j�a<�a<��a<X�a<�a<��a<Q�a< �a<��a</�a<�a<r�a<�a<��a<O�a<סa<�a<�a<��a<Q�a<�a<s�a<��a<��a<>�a<Ýa<L�a<��a<z�a<�a<��a<>�a<ؚa<}�a<�a<��a<B�a<ޘa<z�a< �a<��a<X�a<��a<��a<*�a<�a<��a<*�a<ϔa<��a<6�a<�a<��a<@�a<�a<ْa<|�a<<�a<�a<ؑa<��a<e�a<-�a<�a<Ða<��a<��a<P�a<=�a<+�a<��a<��a<͏a<��a<��a<��a<��a<��a<��a<��a<��a<x�a<��a<��a<��a<ڏa<ԏa<�a<�  �  �a<>�a<e�a<r�a<��a<�a<��a<N�a<R�a<��a<Бa<�a<]�a<k�a<a<�a<��a<��a<�a<J�a<��a<�a<+�a<��a<�a<N�a<��a<�a<h�a<Ɨa<V�a<��a<�a<v�a<��a<k�a<��a<=�a<��a<�a<��a<לa<f�a<ѝa<L�a<��a<K�a<��a<�a<��a<�a<}�a<ȡa<i�a<��a<�a<��a<�a<��a<��a<J�a<��a<�a<]�a<æa<C�a<h�a<٧a<-�a<��a<ƨa<1�a<��a<��a<-�a<\�a<ªa<��a<3�a<��a<��a<�a<*�a<^�a<��a<۬a<	�a<+�a<��a<��a<ҭa<�a<�a<G�a<U�a<��a<s�a<��a<��a<�a<�a<�a<5�a<%�a<`�a<6�a<s�a<v�a<]�a<~�a<x�a<|�a<f�a<��a<r�a<n�a<v�a<\�a<��a<E�a<F�a<3�a<�a<'�a<�a<�a<ٮa<Ʈa<��a<��a<��a<+�a<H�a<��a<�a<��a<��a<��a<%�a<�a<Ĭa<�a<��a<d�a<)�a<�a<Ϋa<g�a<i�a<��a<Īa<��a<Q�a<��a<��a<��a<�a<�a<��a<K�a<�a<��a<o�a<��a<��a<j�a<�a<��a<P�a<��a<��a<Y�a<�a<n�a<&�a<��a<c�a<ءa<��a<
�a<��a<8�a<ȟa<��a<��a<��a<#�a<̝a<V�a<�a<��a<�a<��a<?�a<ښa<Y�a<�a<��a<%�a<�a<d�a<�a<��a<D�a<��a<{�a<K�a<ϕa<r�a<3�a<ٔa<��a<#�a<�a<��a<b�a<�a<ǒa<��a<C�a<.�a<��a<��a<I�a<7�a<�a<ΐa<��a<q�a<y�a<�a<2�a<�a<׏a<ݏa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ɏa<��a<�a<�  �  "�a<C�a<g�a<��a<��a<ϐa<�a<J�a<I�a<��a<̑a<��a<J�a<��a<�a< �a<`�a<��a<��a<B�a<��a<�a</�a<��a<�a<f�a<��a<)�a<y�a<�a<T�a<��a<�a<{�a<ۙa<O�a<��a<7�a<��a<�a<��a<�a<p�a<۝a<Z�a<��a<+�a<��a<�a<��a<�a<u�a<ȡa<9�a<��a<9�a<��a<��a<Y�a<��a<>�a<��a<�a<a�a<��a<�a<�a<�a<:�a<��a<�a<@�a<��a<�a<*�a<[�a<��a<�a<8�a<��a<ǫa<	�a<?�a<s�a<��a<�a<%�a<;�a<p�a<��a<ӭa<�a<�a<;�a<A�a<v�a<��a<Ȯa<�a<�a<�a<�a<2�a<�a<X�a<H�a<Z�a<`�a<v�a<��a<�a<��a<{�a<��a<w�a<��a<v�a<Q�a<Z�a<?�a<N�a<@�a<%�a</�a<�a<�a<ޮa<Ȯa<��a<~�a<g�a<;�a<D�a<�a<�a<��a<��a<n�a<Q�a<.�a<��a<��a<s�a<\�a<!�a<߫a<ϫa<k�a<I�a<�a<ܪa<��a<^�a<	�a<˩a<��a<:�a<��a<��a<G�a<��a<��a<i�a<!�a<��a<w�a<�a<��a<[�a<
�a<��a<9�a<Уa<u�a<�a<��a<\�a<ءa<s�a<�a<Ơa<Y�a<ߟa<g�a<��a<��a<!�a<ȝa<Z�a<ߜa<��a<�a<��a<L�a<�a<s�a<�a<��a<N�a<�a<c�a<�a<��a<I�a<��a<��a<D�a<�a<��a<C�a<�a<��a<3�a<�a<��a<c�a<�a<Ēa<��a<.�a<�a<ّa<��a<s�a<2�a<�a<͐a<��a<i�a<q�a<2�a<�a<��a<�a<�a<Ǐa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ʏa<яa<�a< �a<�  �  $�a<0�a<Q�a<��a<��a<Րa<�a<&�a<p�a<��a<őa< �a<G�a<��a<��a<�a<W�a<Óa<�a<[�a<��a<�a<Y�a<��a<�a<f�a<��a<
�a<v�a<��a<,�a<��a<��a<��a<�a<]�a<�a<�a<��a<��a<��a<��a<f�a<ŝa<E�a<Şa<'�a<��a<�a<��a<�a<`�a<�a<I�a<��a<�a<��a<�a<c�a<�a<-�a<��a<��a<]�a<Ԧa<�a<��a<اa< �a<��a<�a<7�a<g�a<ѩa<�a<��a<��a<�a<P�a<c�a<��a<�a<K�a<q�a<��a<Ǭa<�a<;�a<l�a<��a<��a<��a<*�a<,�a<w�a<s�a<��a<��a<Ȯa<�a<�a<�a<-�a<E�a<@�a<d�a<i�a<V�a<{�a<q�a<o�a<��a<��a<z�a<n�a<`�a<f�a<��a<\�a<t�a<D�a<�a<�a<
�a<�a<��a<ʮa<��a<��a<v�a<m�a<^�a<!�a<�a<�a<��a<��a<k�a<D�a<	�a<�a<��a<��a<L�a<:�a<��a<��a<��a<D�a<��a<ܪa<v�a<@�a<�a<ܩa<g�a<3�a<Ψa<��a<q�a<�a<էa<N�a<	�a<��a<e�a<�a<��a<D�a<��a<��a<5�a<�a<~�a<�a<��a<G�a<��a<��a< �a<��a<:�a<�a<q�a<"�a<��a<A�a<Ɲa<W�a<�a<~�a<#�a<��a<2�a<ޚa<z�a<�a<��a<:�a<��a<��a<�a<ėa<a�a<Ӗa<��a<�a<�a<��a<'�a<Ĕa<��a<3�a<�a<��a<J�a<�a<ߒa<{�a<e�a<�a<ّa<��a<\�a<1�a<�a<Ԑa<��a<��a<Y�a<N�a<)�a<�a<��a<Џa<��a<��a<��a<��a<��a<~�a<��a<��a<��a<Əa<��a<��a<ˏa<ޏa<�a<�  �  �a<F�a<n�a<��a<��a<̐a<��a<-�a<U�a<��a<��a<�a<?�a<��a<Вa<�a<[�a<��a<ړa<M�a<��a<�a<>�a<��a<�a<b�a<��a<'�a<l�a<ڗa<I�a<ʘa<�a<z�a<ؙa<C�a<��a<.�a<��a<(�a<��a<�a<r�a<ٝa<V�a<��a<,�a<��a<�a<z�a<�a<X�a<ša<I�a<��a</�a<��a<��a<a�a<��a<#�a<��a<�a<c�a<��a<�a<o�a<�a<7�a<��a<ڨa<9�a<��a<�a<�a<a�a<��a<�a<9�a<��a<�a<�a<7�a<e�a<��a<�a<�a<3�a<h�a<��a<ía<�a<�a<�a<]�a<u�a<��a<��a<߮a<ܮa<	�a<��a<$�a<)�a<@�a<P�a<U�a<f�a<j�a<��a<��a<|�a<y�a<��a<��a<��a<f�a<e�a<P�a<N�a<<�a<M�a<E�a<"�a<��a<�a<�a<Ϯa<��a<��a<d�a<I�a<'�a<��a<�a<��a<��a<d�a<S�a<�a<�a<��a<��a<=�a<,�a<�a<��a<z�a<A�a<��a<تa<��a<]�a<��a<��a<��a<V�a<��a<��a<C�a<�a<��a<`�a<'�a<Ѧa<l�a<�a<��a<X�a<�a<��a<:�a<ǣa<|�a<�a<��a<>�a<աa<��a<�a<��a<U�a<ܟa<o�a<��a<��a<,�a<��a<]�a<ޜa<��a<
�a<��a<I�a<�a<m�a<�a<��a<V�a<֘a<j�a< �a<��a<J�a<��a<��a<=�a<ܕa<y�a<A�a<�a<��a<+�a<�a<��a<S�a<�a<˒a<l�a<K�a<�a<ϑa<��a<r�a<%�a<�a<��a<��a<u�a<X�a<:�a<�a< �a<�a<�a<ɏa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<֏a<�a<��a<��a<�  �  !�a<�a<P�a<o�a<��a<ѐa<�a<>�a<K�a<��a<Ƒa<�a<D�a<��a<��a<�a<X�a<��a<��a<K�a<|�a<��a<'�a<��a<�a<O�a<��a<��a<v�a<ڗa<A�a<��a<�a<w�a<�a<i�a<��a<=�a<��a<��a<��a<�a<d�a<��a<N�a<��a<>�a<��a<�a<t�a<�a<s�a<̡a<R�a<��a<�a<}�a<�a<u�a<��a<@�a<��a<�a<c�a<��a<7�a<g�a<�a<�a<��a<ިa<3�a<w�a<��a<)�a<`�a<êa<��a<8�a<x�a<��a<��a<;�a<t�a<��a<ìa<�a<1�a<��a<��a<խa<֭a<�a<C�a<P�a<��a<��a<��a<��a<�a<
�a<�a<9�a<#�a<Q�a<J�a<Z�a<i�a<\�a<p�a<a�a<��a<w�a<~�a<\�a<d�a<y�a<e�a<r�a<P�a<J�a<+�a<�a<�a<��a<�a<��a<��a<��a<��a<j�a<8�a<;�a<�a<��a<��a<��a<k�a<;�a<�a<�a<��a<��a<^�a<,�a<իa<̫a<e�a<V�a<��a<Ǫa<u�a<3�a<�a<éa<~�a<�a<�a<��a<Q�a<�a<��a<o�a<�a<��a<c�a<�a<��a<;�a<��a<��a<L�a<ˣa<y�a<�a<��a<Y�a<ܡa<��a<�a<��a<4�a<ҟa<��a<��a<��a<!�a<��a<\�a<؜a<��a<�a<��a<'�a<՚a<p�a<	�a<��a<�a<ߘa<h�a<�a<��a<H�a<�a<n�a<4�a<ߕa<��a<�a<��a<��a<'�a<��a<��a<b�a<��a<ʒa<��a<;�a<�a<ȑa<|�a<Q�a<)�a<
�a<Ɛa<��a<l�a<h�a<2�a<�a<�a<ԏa<͏a<��a<��a<��a<��a<w�a<��a<��a<��a<��a<��a<��a<��a<��a<�a<��a<�  �  �a<<�a<Z�a<t�a<��a<ΐa<�a<(�a<]�a<��a<��a<�a<5�a<��a<ϒa<�a<D�a<��a<�a<C�a<��a<�a<5�a<��a<�a<Q�a<��a<�a<d�a<՗a<>�a<��a<�a<s�a<әa<?�a<��a<,�a<��a<�a<�a<ܜa<b�a<ߝa<N�a<��a<+�a<��a<�a<x�a<��a<X�a<ϡa<9�a<��a<(�a<��a<��a<U�a<Ťa<#�a<��a<�a<V�a<��a< �a<m�a<ߧa<:�a<��a<ʨa<3�a<��a<ةa<�a<e�a<��a<�a<9�a<{�a<ȫa<��a<9�a<_�a<��a<�a<�a<3�a<r�a<��a<��a<�a<�a<&�a<V�a<e�a<��a<��a<خa<׮a<��a<�a<!�a<5�a<A�a<H�a<Y�a<a�a<e�a<w�a<�a<w�a<m�a<{�a<~�a<x�a<i�a<a�a<F�a<J�a<>�a<9�a<.�a<�a<�a<�a<ٮa<��a<��a<|�a<g�a<?�a<%�a<�a<�a<��a<��a<[�a<N�a<�a<��a<��a<��a<F�a<$�a<�a<��a<s�a<H�a<��a<Ȫa<��a<Q�a<��a<��a<{�a<?�a<�a<��a<@�a<�a<��a<_�a<�a<��a<b�a<��a<��a<^�a<��a<��a<9�a<Уa<m�a<
�a<��a<?�a<�a<r�a<�a<��a<K�a<֟a<c�a<��a<��a<0�a<��a<O�a<�a<��a<�a<��a<K�a<ښa<[�a<	�a<��a<@�a<՘a<l�a<��a<��a<H�a<�a<��a<7�a<ܕa<q�a<4�a<��a<��a<)�a<�a<��a<N�a<�a<ƒa<t�a<B�a<�a<Ցa<��a<i�a<�a<��a<a<��a<~�a<W�a</�a<�a<��a<ݏa<ӏa<ďa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<؏a<�a<��a<�  �  �a<7�a<C�a<��a<��a<Ӑa<��a<�a<i�a<��a<ϑa<�a<:�a<��a<��a<�a<E�a<��a<�a<B�a<��a<ٔa<K�a<��a<��a<N�a<��a<�a<f�a<�a<�a<��a<��a<x�a<�a<D�a<њa<�a<��a<��a<z�a<�a<X�a<Нa<5�a<��a<&�a<��a<�a<z�a<�a<T�a<�a<:�a<��a<
�a<r�a<��a<R�a<�a<!�a<��a<��a<Y�a<Ѧa<�a<��a<Ƨa<'�a<}�a<Ҩa<4�a<l�a<ԩa<�a<y�a<��a<��a<B�a<h�a<īa<�a<C�a<c�a<��a<̬a<�a<E�a<k�a<��a<��a<�a<�a<*�a<s�a<e�a<��a<��a<Ȯa<ޮa<�a<�a<�a<A�a<4�a<P�a<c�a<h�a<v�a<]�a<w�a<t�a<~�a<h�a<n�a<p�a<_�a<w�a<J�a<`�a<9�a<,�a<!�a<��a<�a<�a<Ԯa<��a<��a<��a<m�a<L�a<�a<�a<ۭa<��a<��a<`�a<A�a<��a<�a<��a<��a<N�a<#�a<�a<��a<��a<C�a<�a<ƪa<w�a<M�a<��a<̩a<\�a<8�a<ըa<��a<V�a<��a<ħa<I�a<�a<��a<]�a<�a<��a<O�a<�a<��a<5�a<�a<s�a<�a<��a<:�a<��a<t�a<�a<��a<)�a<۟a<`�a<�a<��a<;�a<��a<R�a<��a<{�a<�a<��a<8�a<̚a<d�a<�a<��a<<�a<��a<��a<�a<��a<R�a<֖a<��a<�a<�a<u�a<+�a<ǔa<{�a<;�a<�a<��a<E�a<
�a<ɒa<w�a<^�a<�a<ԑa<x�a<Z�a<%�a<�a<֐a<��a<��a<J�a<7�a<!�a<�a<�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ˏa<Ώa<�a<�  �  �a<2�a<R�a<~�a<��a<ΐa<�a<2�a<N�a<��a<ʑa<��a<A�a<��a<̒a<�a<Q�a<��a<�a<?�a<��a<�a</�a<��a<�a<S�a<��a<�a<n�a<Зa<6�a<��a<�a<u�a<יa<H�a<��a</�a<��a<�a<|�a<�a<c�a<ϝa<F�a<��a< �a<��a<�a<��a<�a<e�a<ša<9�a<��a<!�a<��a<��a<Y�a<��a<2�a<��a<��a<_�a<��a<�a<v�a<اa<+�a<��a<֨a<.�a<�a<٩a< �a<a�a<��a<�a<6�a<��a<ëa<��a</�a<j�a<��a<Ѭa<�a<8�a<i�a<��a<̭a<�a<�a<6�a<J�a<q�a<��a<��a<Ѯa<�a<�a<	�a<$�a<&�a<H�a<H�a<X�a<a�a<n�a<n�a<s�a<}�a<s�a<v�a<t�a<��a<p�a<V�a<X�a<B�a<F�a<A�a<#�a<�a<��a<�a<Ϯa<��a<��a<��a<h�a<<�a<.�a<��a<�a<��a<��a<h�a<G�a<�a<�a<��a<z�a<W�a< �a<�a<��a<m�a<B�a<��a<˪a<~�a<H�a< �a<��a<r�a<7�a<�a<��a<C�a<��a<��a<b�a<�a<��a<^�a<�a<��a<O�a<��a<��a<.�a<ͣa<t�a<�a<��a<L�a<աa<s�a<�a<��a<D�a<ڟa<f�a<��a<��a<$�a<��a<X�a<�a<w�a<�a<��a<<�a<֚a<h�a<�a<��a<A�a<טa<h�a<�a<��a<F�a<�a<��a<.�a<ӕa<|�a<+�a<͔a<��a<.�a<�a<��a<Z�a<�a<��a<��a<5�a<��a<ёa<��a<b�a<(�a<�a<Ȑa<��a<p�a<^�a</�a<�a<��a<�a<ʏa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ȏa<͏a<ߏa<��a<�  �   �a<,�a<X�a<q�a<��a<ܐa<�a<?�a<G�a<��a<ˑa<
�a<I�a<w�a<ܒa<��a<f�a<��a<��a<B�a<��a<��a<(�a<��a<�a<P�a<��a<�a<y�a<ʗa<K�a<��a<�a<s�a<�a<g�a<��a<1�a<��a<�a<�a<�a<l�a<ǝa<J�a<��a<5�a<��a<�a<��a<ݠa<t�a<ša<V�a<��a<�a<��a<�a<t�a<��a<B�a<��a<�a<b�a<��a<,�a<f�a<ۧa<&�a<��a<ڨa<-�a<��a<��a<#�a<\�a<êa<��a<3�a<��a<��a<�a<)�a<q�a<��a<Ԭa<�a<-�a<��a<��a<ԭa<�a<�a<B�a<O�a<��a<~�a<��a<®a<�a<�a<
�a<2�a<�a<W�a<C�a<d�a<f�a<_�a<x�a<n�a<��a<m�a<��a<r�a<f�a<r�a<T�a<w�a<C�a<F�a<.�a<�a<�a<�a<�a<ɮa<��a<��a<��a<v�a<4�a<;�a<�a<�a<��a<��a<o�a<2�a<(�a<Ҭa<Ǭa<��a<`�a<#�a<߫a<ɫa<f�a<X�a<��a<Ǫa<��a<B�a<�a<��a<��a< �a<�a<��a<O�a<�a<��a<d�a<��a<��a<a�a< �a<��a<G�a<��a<��a<D�a<ңa<r�a<!�a<��a<Z�a<աa<��a<�a<��a<E�a<a<��a<��a<��a<�a<ʝa<[�a<��a<��a<�a<��a<7�a<��a<k�a<�a<��a< �a<٘a<c�a<�a<��a<B�a<�a<w�a<@�a<͕a<��a<*�a<Дa<��a<#�a<��a<��a<b�a<�a<��a<��a<;�a<�a<��a<��a<S�a<'�a<�a<ɐa<��a<g�a<m�a<*�a<!�a<��a<׏a<ԏa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<Ïa<�a<�a<�  �  �a</�a<S�a<��a<��a<Ða<��a<)�a<e�a<��a<��a<�a<G�a<��a<ђa<�a<X�a<��a<�a<=�a<��a<�a<A�a<��a<�a<\�a<��a<�a<x�a<ޗa<4�a<��a<	�a<t�a<�a<J�a<��a<*�a<��a<�a<{�a<��a<_�a<ɝa<I�a<a<�a<��a<�a<��a<�a<]�a<ǡa<A�a<��a<!�a<��a<��a<]�a<��a<'�a<��a<��a<X�a<��a<�a<��a<ݧa<(�a<��a<�a</�a<��a<ϩa<�a<i�a<��a<�a<7�a<y�a<��a<�a<9�a<u�a<��a<լa<�a<@�a<]�a<��a<��a<�a<�a<*�a<Q�a<v�a<��a<��a<ʮa<�a<��a<�a<"�a<<�a<C�a<M�a<S�a<T�a<y�a<r�a<q�a<v�a<��a<t�a<y�a<j�a<i�a<h�a<P�a<T�a<C�a<.�a<$�a<�a<	�a<�a<̮a<��a<��a<w�a<]�a<H�a<&�a<�a<�a<��a<��a<m�a<;�a<�a<�a<��a<��a<J�a<�a<�a<��a<�a<4�a<�a<Ԫa<��a<@�a<
�a<ǩa<p�a<0�a<�a<��a<P�a<��a<��a<\�a<	�a<��a<]�a<�a<��a<I�a<��a<��a<'�a<ѣa<n�a<�a<��a<C�a<ءa<{�a<�a<��a<D�a<֟a<j�a<��a<��a<+�a<ŝa<Q�a<�a<o�a<�a<��a<8�a<֚a<w�a<�a<��a<7�a<јa<q�a<�a<��a<F�a<�a<��a<*�a<ݕa<��a<'�a<єa<��a<6�a<֓a<��a<N�a<�a<��a<w�a<=�a<�a<Ǒa<��a<[�a</�a<��a<��a<��a<��a<Y�a<5�a<�a<�a<�a<Ϗa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<Ώa<ُa<�a<�  �  �a<I�a<F�a<~�a<��a<��a<�a<�a<i�a<��a<Ցa<�a<;�a<��a<��a<�a<D�a<��a<�a<4�a<��a<Ӕa<S�a<��a<��a<A�a<��a<�a<a�a<��a<)�a<��a<��a<u�a<�a<A�a<͚a<�a<��a<�a<t�a<�a<T�a<�a<,�a<ʞa<�a<��a<�a<t�a<��a<P�a<�a<-�a<��a<�a<��a<�a<I�a<ڤa< �a<��a<�a<V�a<Ǧa<	�a<��a<��a<<�a<}�a<ըa<+�a<r�a<ߩa<�a<t�a<��a<��a<>�a<j�a<ͫa<�a<;�a<a�a<��a<٬a<��a<M�a<R�a<��a<��a<�a<�a<0�a<b�a<c�a<��a<��a<Үa<߮a<�a<�a<�a<>�a</�a<[�a<S�a<Y�a<u�a<^�a<��a<d�a<��a<k�a<z�a<s�a<Y�a<r�a<D�a<Y�a<6�a<1�a<-�a<�a<
�a<Ԯa<�a<��a<��a<��a<X�a<Y�a<�a<�a<έa<ŭa<��a<b�a<J�a<�a<��a<��a<��a<V�a<�a<�a<��a<��a<+�a<�a<��a<��a<N�a<�a<ɩa<f�a<?�a<٨a<��a<T�a<�a<��a<I�a<�a<��a<W�a<�a<��a<c�a<ݤa<��a<'�a<ڣa<t�a<�a<��a<7�a<��a<g�a<�a<��a<9�a<�a<W�a<�a<��a<+�a<��a<N�a<��a<k�a<(�a<��a<L�a<͚a<g�a<�a<��a<H�a<��a<{�a< �a<��a<M�a<ٖa<��a<�a<ޕa<s�a<,�a<Ԕa<r�a<C�a<̓a<��a<A�a<�a<��a<~�a<N�a<�a<ۑa<��a<d�a<&�a<�a<ِa<��a<��a<E�a<B�a<�a<�a<�a<��a<ҏa<��a<��a<��a<��a<��a<{�a<��a<��a<��a<��a<��a<׏a<ҏa<�a<�  �  �a<6�a<K�a<q�a<��a<Ȑa<�a<+�a<g�a<��a<ˑa<�a<F�a<��a<��a<�a<U�a<��a<�a<=�a<��a<�a<8�a<��a<��a<>�a<��a<�a<s�a<ݗa<<�a<��a<
�a<{�a<�a<R�a<��a<*�a<��a< �a<x�a<�a<^�a<ѝa<4�a<��a<6�a<��a<�a<��a<��a<\�a<ӡa<?�a<��a<�a<��a<��a<_�a<ʤa<.�a<��a<�a<\�a<��a<&�a<��a<ŧa<,�a<��a<�a<,�a<u�a<ǩa<�a<d�a<��a<��a<<�a<{�a<��a<��a<7�a<p�a<��a<Ӭa<��a<I�a<o�a<��a<��a<��a<�a<7�a<S�a<u�a<��a<��a<ήa<�a<��a<�a<�a<;�a<G�a<G�a<W�a<s�a<g�a<f�a<z�a<v�a<}�a<w�a<k�a<q�a<l�a<^�a<c�a<I�a<C�a<4�a<�a<�a<�a<�a<Ӯa<��a<��a<��a<a�a<?�a<(�a<�a<֭a<��a<��a<l�a<E�a<�a<�a<��a<��a<X�a<�a<��a<��a<v�a<C�a<�a<��a<�a<B�a<�a<Ʃa<y�a<#�a<�a<��a<O�a<�a<��a<]�a<�a<��a<[�a<�a<��a<Q�a<�a<��a<D�a<ңa<t�a<�a<��a<C�a<�a<x�a<�a<��a<=�a<ڟa<l�a<�a<��a<.�a<ʝa<U�a<�a<��a<�a<��a<=�a<Қa<q�a<�a<��a</�a<Ϙa<k�a<�a<��a<K�a<�a<��a<.�a<ڕa<��a<#�a<Δa<r�a<?�a<�a<��a<N�a<�a<a<��a<?�a<�a<ϑa<��a<_�a<(�a<��a<͐a<��a<��a<]�a<.�a<�a<�a<ߏa<Ïa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<Ïa<�a<�a<�  �  +�a<�a<h�a<t�a<��a<̐a<�a<3�a<P�a<��a<��a<�a<G�a<|�a<�a< �a<^�a<��a<�a<H�a<��a<�a<4�a<��a<�a<S�a<��a<�a<��a<��a<M�a<��a<�a<n�a<ڙa<[�a<��a<?�a<��a<�a<u�a<�a<p�a<��a<X�a<��a<.�a<��a<�a<��a<�a<p�a<��a<G�a<��a<(�a<��a<�a<g�a<��a<>�a<��a<��a<f�a<��a<"�a<g�a<�a<!�a<��a<�a<"�a<��a<ũa<0�a<P�a<��a<�a<*�a<��a<��a<�a<�a<~�a<��a<جa<�a<-�a<r�a<��a<ϭa<�a<�a<9�a<D�a<|�a<��a<̮a<Ǯa<�a<��a< �a<0�a<&�a<K�a<I�a<V�a<b�a<a�a<��a<_�a<��a<j�a<}�a<~�a<m�a<x�a<P�a<o�a<?�a<J�a<5�a<&�a<�a<�a<��a<��a<ˮa<��a<|�a<f�a<?�a<0�a<��a<�a<��a<��a<m�a<8�a<3�a<جa<��a<y�a<T�a<)�a<�a<��a<r�a<H�a<��a<˪a<��a<<�a<�a<��a<��a<*�a<�a<��a<G�a<�a<��a<q�a<�a<Ʀa<W�a<�a<��a<=�a<	�a<��a<<�a<Уa<y�a<�a<��a<W�a<ˡa<��a<�a<��a<R�a<Οa<t�a<�a<��a<(�a<a<^�a<�a<��a<�a<��a<2�a<��a<t�a<��a<��a<-�a<�a<W�a<�a<��a<9�a<��a<��a<C�a<��a<��a<#�a<Ԕa<��a<$�a<�a<��a<]�a< �a<Ȓa<��a</�a<
�a<��a<��a<Y�a<(�a<��a<��a<��a<p�a<a�a<0�a<�a<��a<ُa<�a<��a<��a<��a<��a<��a<��a<��a<|�a<��a<��a<��a<��a<Ϗa<�a<�a<�  �   �a<(�a<X�a<x�a<��a<Ɛa<��a<'�a<W�a<��a<̑a<�a<G�a<y�a<ƒa<�a<^�a<��a<�a<>�a<��a<�a<;�a<��a<�a<K�a<��a<�a<v�a<ʗa<>�a<��a<�a<s�a<�a<S�a<a<&�a<��a<�a<x�a<�a<j�a<Ɲa<A�a<��a</�a<��a<�a<}�a<�a<_�a<ڡa<H�a<��a<�a<��a<�a<e�a<Ѥa<.�a<��a<��a<\�a<��a< �a<u�a<ϧa<%�a<��a<ڨa<(�a<��a<©a<�a<k�a<��a<��a<7�a<s�a<��a<��a<)�a<q�a<��a<Ѭa<�a<;�a<l�a<��a<ƭa<�a<�a<1�a<f�a<|�a<��a<��a<��a<�a<�a<�a<�a<-�a<?�a<Q�a<P�a<g�a<g�a<s�a<h�a<��a<n�a<x�a<x�a<d�a<f�a<i�a<\�a<V�a<?�a<(�a<#�a<�a<�a<�a<Ůa<��a<��a<��a<`�a<F�a<$�a<��a<ܭa<��a<��a<m�a<4�a<�a<۬a<��a<��a<S�a<�a<�a<��a<x�a<=�a<�a<êa<��a<@�a<�a<��a<{�a<)�a<ݨa<��a<T�a<�a<��a<Y�a<��a<��a<[�a<�a<��a<F�a<�a<��a<>�a<Уa<u�a<�a<��a<F�a<�a<��a<�a<��a<9�a<ҟa<r�a<�a<��a<*�a<��a<U�a<�a<��a<�a<��a<6�a<ۚa<k�a<��a<��a<*�a<̘a<r�a<�a<��a<F�a<�a<��a<4�a<̕a<��a<&�a<͔a<z�a<2�a<�a<��a<T�a<�a<Ēa<~�a<R�a<
�a<��a<��a<Q�a<)�a<�a<Ґa<��a<w�a<U�a<8�a<�a< �a<ߏa<Џa<��a<��a<��a<��a<��a<�a<��a<��a<��a<��a<��a<��a<͏a<�a<�a<�  �  �a<<�a<[�a<~�a<��a<��a<��a<�a<e�a<|�a<͑a<��a<>�a<��a<��a<#�a<H�a<��a<�a<3�a<��a<�a<?�a<��a<��a<S�a<��a<�a<e�a<�a<0�a<��a<�a<s�a<ܙa<6�a<ƚa<�a<��a<��a<��a<�a<W�a<�a<C�a<��a<�a<��a<�a<v�a<��a<K�a<ۡa<-�a<��a< �a<��a<�a<K�a<Τa<�a<��a<�a<U�a<��a<�a<��a<ҧa<B�a<��a<ۨa<<�a<r�a<�a<�a<l�a<��a<�a<8�a<x�a<ϫa<�a<E�a<f�a<��a<�a<�a<G�a<[�a<��a<��a<�a<�a<%�a<X�a<c�a<��a<��a<Ԯa<�a<�a<�a<�a<?�a<7�a<V�a<H�a<e�a<q�a<u�a<��a<i�a<��a<y�a<q�a<��a<Z�a<h�a<<�a<Q�a<4�a<H�a<$�a<�a<�a<خa<ٮa<��a<��a<��a<S�a<J�a<�a<�a<ɭa<��a<��a<d�a<O�a<�a<��a<��a<��a<J�a<�a<�a<��a<|�a<-�a<�a<˪a<��a<F�a<��a<ϩa<m�a<=�a<�a<��a<I�a<�a<��a<M�a<&�a<��a<e�a<�a<��a<b�a<�a<��a<-�a<ʣa<s�a<�a<��a<2�a<�a<g�a< �a<��a<?�a<�a<X�a<�a<��a<4�a<��a<M�a<��a<q�a<�a<��a<R�a<Кa<m�a<�a<��a<P�a<Øa<s�a<�a<��a<G�a<�a<��a<$�a<�a<x�a<(�a<�a<��a<=�a<Փa<��a<J�a<�a<��a<s�a<D�a<�a<ߑa<��a<f�a<(�a<�a<Ԑa<��a<��a<M�a<=�a<�a<��a<�a<ҏa<Ǐa<��a<��a<��a<��a<��a<{�a<��a<x�a<��a<��a<Ϗa<Ώa<��a<�a<�  �  �a<,�a<Y�a<q�a<��a<Аa<�a<"�a<S�a<��a<ؑa<�a<@�a<~�a<��a<�a<V�a<��a<��a<A�a<��a<�a<G�a<��a<�a<O�a<��a<�a<o�a<ٗa<9�a<��a<�a<l�a<�a<W�a<Śa<�a<��a<��a<~�a<�a<\�a<ʝa<J�a<��a<0�a<��a<�a<p�a<��a<h�a<ޡa<B�a<��a<�a<z�a<��a<c�a<Ҥa<8�a<��a<�a<c�a<ʦa<%�a<o�a<ڧa<&�a<��a<ըa<3�a<s�a<̩a<�a<h�a<��a<�a<3�a<v�a<��a<�a<8�a<h�a<��a<Ӭa<�a<0�a<t�a<��a<ĭa<٭a<�a<@�a<]�a<x�a<��a<��a<��a<�a<��a<�a<#�a</�a<6�a<Y�a<_�a<b�a<`�a<x�a<n�a<w�a<t�a<{�a<f�a<s�a<W�a<r�a<`�a<\�a<1�a<5�a<�a<�a<��a<�a<ɮa<��a<��a<~�a<j�a<O�a<�a<��a<�a<ȭa<��a<g�a<:�a<�a<�a<��a<��a<^�a<"�a<ݫa<��a<��a<G�a<��a<ƪa<��a<?�a<�a<��a<v�a<)�a<�a<��a<[�a<	�a<��a<O�a<	�a<��a<a�a<�a<��a<I�a<��a<��a<>�a<�a<�a<�a<��a<N�a<�a<|�a<�a<��a<1�a<֟a<p�a<�a<��a<0�a<��a<\�a<��a<��a<	�a<��a<7�a<Кa<g�a<	�a<��a<4�a<ǘa<o�a<�a<��a<B�a<�a<��a<)�a<ەa<z�a<"�a<ϔa<��a<&�a<�a<��a<R�a<��a<ƒa<��a<I�a<�a<ɑa<��a<P�a<'�a<��a<ܐa<��a<y�a<L�a<A�a<�a<��a<؏a<Տa<��a<��a<��a<��a<��a<��a<y�a<��a<��a<��a<��a<��a<��a<�a<��a<�  �  -�a<"�a<]�a<v�a<��a<Ða<�a<3�a<[�a<��a<��a<��a<I�a<��a<�a<�a<g�a<��a<ٓa<E�a<��a<�a<(�a<��a<ߕa<X�a<��a<�a<{�a<Ɨa<S�a<��a<�a<v�a<ՙa<9�a<��a<;�a<��a<�a<�a<ۜa<o�a<��a<_�a<��a<0�a<��a<�a<��a<��a<a�a<��a<B�a<��a<&�a<��a<�a<j�a<��a<*�a<��a<��a<Y�a<��a<'�a<i�a<�a<�a<��a<˨a<)�a<��a<ȩa<2�a<a�a<��a<�a<5�a<��a<��a<�a<$�a<h�a<��a<Ѭa<�a<&�a<s�a<��a<ȭa<�a<�a<%�a<?�a<��a<��a<ήa<ͮa<�a<�a<�a<'�a<4�a<G�a<:�a<J�a<`�a<b�a<��a<`�a<��a<b�a<��a<{�a<o�a<j�a<c�a<H�a<L�a<C�a<8�a<#�a<$�a<�a<��a<��a<��a<��a<z�a<]�a<3�a</�a<�a<�a<��a<��a<p�a<B�a</�a<�a<Ȭa<v�a<>�a<&�a<�a<��a<e�a<B�a<�a<Ъa<��a<D�a<�a<��a<��a<*�a<��a<��a<B�a<�a<��a<m�a<�a<Ŧa<b�a<��a<��a<@�a<�a<��a<>�a<��a<m�a<�a<��a<G�a<ġa<|�a<�a<��a<Q�a<ҟa<w�a<�a<��a<0�a<Ɲa<R�a<Ӝa<��a<�a<ƛa<,�a<ޚa<]�a<��a<��a<0�a<�a<h�a<��a<��a<E�a<��a<��a<C�a<Ǖa<z�a<,�a<̔a<��a<�a<�a<��a<V�a<�a<ʒa<s�a<*�a<�a<Ƒa<��a<^�a<-�a<�a<��a<��a<~�a<]�a<!�a<�a<��a<ڏa<ߏa<��a<ďa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<͏a<��a<�a<�  �  �a<,�a<Y�a<q�a<��a<Аa<�a<"�a<S�a<��a<ؑa<�a<@�a<~�a<��a<�a<V�a<��a<��a<A�a<��a<�a<G�a<��a<�a<O�a<��a<�a<o�a<ٗa<9�a<��a<�a<l�a<�a<W�a<Śa<�a<��a<��a<~�a<�a<\�a<ʝa<J�a<��a<0�a<��a<�a<p�a<��a<h�a<ޡa<B�a<��a<�a<z�a<��a<c�a<Ҥa<8�a<��a<�a<c�a<ʦa<%�a<o�a<ڧa<&�a<��a<ըa<3�a<s�a<̩a<�a<h�a<��a<�a<3�a<v�a<��a<�a<8�a<h�a<��a<Ӭa<�a<0�a<t�a<��a<ĭa<٭a<�a<@�a<]�a<x�a<��a<��a<��a<�a<��a<�a<#�a</�a<6�a<Y�a<_�a<b�a<`�a<x�a<n�a<w�a<t�a<{�a<f�a<s�a<W�a<r�a<`�a<\�a<1�a<5�a<�a<�a<��a<�a<ɮa<��a<��a<~�a<j�a<O�a<�a<��a<�a<ȭa<��a<g�a<:�a<�a<�a<��a<��a<^�a<"�a<ݫa<��a<��a<G�a<��a<ƪa<��a<?�a<�a<��a<v�a<)�a<�a<��a<[�a<	�a<��a<O�a<	�a<��a<a�a<�a<��a<I�a<��a<��a<>�a<�a<�a<�a<��a<N�a<�a<|�a<�a<��a<1�a<֟a<p�a<�a<��a<0�a<��a<\�a<��a<��a<	�a<��a<7�a<Кa<g�a<	�a<��a<4�a<ǘa<o�a<�a<��a<B�a<�a<��a<)�a<ەa<z�a<"�a<ϔa<��a<&�a<�a<��a<R�a<��a<ƒa<��a<I�a<�a<ɑa<��a<P�a<'�a<��a<ܐa<��a<y�a<L�a<A�a<�a<��a<؏a<Տa<��a<��a<��a<��a<��a<��a<y�a<��a<��a<��a<��a<��a<��a<�a<��a<�  �  �a<<�a<[�a<~�a<��a<��a<��a<�a<e�a<|�a<͑a<��a<>�a<��a<��a<#�a<H�a<��a<�a<3�a<��a<�a<?�a<��a<��a<S�a<��a<�a<e�a<�a<0�a<��a<�a<s�a<ܙa<6�a<ƚa<�a<��a<��a<��a<�a<W�a<�a<C�a<��a<�a<��a<�a<v�a<��a<K�a<ۡa<-�a<��a< �a<��a<�a<K�a<Τa<�a<��a<�a<U�a<��a<�a<��a<ҧa<B�a<��a<ۨa<<�a<r�a<�a<�a<l�a<��a<�a<8�a<x�a<ϫa<�a<E�a<f�a<��a<�a<�a<G�a<[�a<��a<��a<�a<�a<%�a<X�a<c�a<��a<��a<Ԯa<�a<�a<�a<�a<?�a<7�a<V�a<H�a<e�a<q�a<u�a<��a<i�a<��a<y�a<q�a<��a<Z�a<h�a<<�a<Q�a<4�a<H�a<$�a<�a<�a<خa<ٮa<��a<��a<��a<S�a<J�a<�a<�a<ɭa<��a<��a<d�a<O�a<�a<��a<��a<��a<J�a<�a<�a<��a<|�a<-�a<�a<˪a<��a<F�a<��a<ϩa<m�a<=�a<�a<��a<I�a<�a<��a<M�a<&�a<��a<e�a<�a<��a<b�a<�a<��a<-�a<ʣa<s�a<�a<��a<2�a<�a<g�a< �a<��a<?�a<�a<X�a<�a<��a<4�a<��a<M�a<��a<q�a<�a<��a<R�a<Кa<m�a<�a<��a<P�a<Øa<s�a<�a<��a<G�a<�a<��a<$�a<�a<x�a<(�a<�a<��a<=�a<Փa<��a<J�a<�a<��a<s�a<D�a<�a<ߑa<��a<f�a<(�a<�a<Ԑa<��a<��a<M�a<=�a<�a<��a<�a<ҏa<Ǐa<��a<��a<��a<��a<��a<{�a<��a<x�a<��a<��a<Ϗa<Ώa<��a<�a<�  �   �a<(�a<X�a<x�a<��a<Ɛa<��a<'�a<W�a<��a<̑a<�a<G�a<y�a<ƒa<�a<^�a<��a<�a<>�a<��a<�a<;�a<��a<�a<K�a<��a<�a<v�a<ʗa<>�a<��a<�a<s�a<�a<S�a<a<&�a<��a<�a<x�a<�a<j�a<Ɲa<A�a<��a</�a<��a<�a<}�a<�a<_�a<ڡa<H�a<��a<�a<��a<�a<e�a<Ѥa<.�a<��a<��a<\�a<��a< �a<u�a<ϧa<%�a<��a<ڨa<(�a<��a<©a<�a<k�a<��a<��a<7�a<s�a<��a<��a<)�a<q�a<��a<Ѭa<�a<;�a<l�a<��a<ƭa<�a<�a<1�a<f�a<|�a<��a<��a<��a<�a<�a<�a<�a<-�a<?�a<Q�a<P�a<g�a<g�a<s�a<h�a<��a<n�a<x�a<x�a<d�a<f�a<i�a<\�a<V�a<?�a<(�a<#�a<�a<�a<�a<Ůa<��a<��a<��a<`�a<F�a<$�a<��a<ܭa<��a<��a<m�a<4�a<�a<۬a<��a<��a<S�a<�a<�a<��a<x�a<=�a<�a<êa<��a<@�a<�a<��a<{�a<)�a<ݨa<��a<T�a<�a<��a<Y�a<��a<��a<[�a<�a<��a<F�a<�a<��a<>�a<Уa<u�a<�a<��a<F�a<�a<��a<�a<��a<9�a<ҟa<r�a<�a<��a<*�a<��a<U�a<�a<��a<�a<��a<6�a<ۚa<k�a<��a<��a<*�a<̘a<r�a<�a<��a<F�a<�a<��a<4�a<̕a<��a<&�a<͔a<z�a<2�a<�a<��a<T�a<�a<Ēa<~�a<R�a<
�a<��a<��a<Q�a<)�a<�a<Ґa<��a<w�a<U�a<8�a<�a< �a<ߏa<Џa<��a<��a<��a<��a<��a<�a<��a<��a<��a<��a<��a<��a<͏a<�a<�a<�  �  +�a<�a<h�a<t�a<��a<̐a<�a<3�a<P�a<��a<��a<�a<G�a<|�a<�a< �a<^�a<��a<�a<H�a<��a<�a<4�a<��a<�a<S�a<��a<�a<��a<��a<M�a<��a<�a<n�a<ڙa<[�a<��a<?�a<��a<�a<u�a<�a<p�a<��a<X�a<��a<.�a<��a<�a<��a<�a<p�a<��a<G�a<��a<(�a<��a<�a<g�a<��a<>�a<��a<��a<f�a<��a<"�a<g�a<�a<!�a<��a<�a<"�a<��a<ũa<0�a<P�a<��a<�a<*�a<��a<��a<�a<�a<~�a<��a<جa<�a<-�a<r�a<��a<ϭa<�a<�a<9�a<D�a<|�a<��a<̮a<Ǯa<�a<��a< �a<0�a<&�a<K�a<I�a<V�a<b�a<a�a<��a<_�a<��a<j�a<}�a<~�a<m�a<x�a<P�a<o�a<?�a<J�a<5�a<&�a<�a<�a<��a<��a<ˮa<��a<|�a<f�a<?�a<0�a<��a<�a<��a<��a<m�a<8�a<3�a<جa<��a<y�a<T�a<)�a<�a<��a<r�a<H�a<��a<˪a<��a<<�a<�a<��a<��a<*�a<�a<��a<G�a<�a<��a<q�a<�a<Ʀa<W�a<�a<��a<=�a<	�a<��a<<�a<Уa<y�a<�a<��a<W�a<ˡa<��a<�a<��a<R�a<Οa<t�a<�a<��a<(�a<a<^�a<�a<��a<�a<��a<2�a<��a<t�a<��a<��a<-�a<�a<W�a<�a<��a<9�a<��a<��a<C�a<��a<��a<#�a<Ԕa<��a<$�a<�a<��a<]�a< �a<Ȓa<��a</�a<
�a<��a<��a<Y�a<(�a<��a<��a<��a<p�a<a�a<0�a<�a<��a<ُa<�a<��a<��a<��a<��a<��a<��a<��a<|�a<��a<��a<��a<��a<Ϗa<�a<�a<�  �  �a<6�a<K�a<q�a<��a<Ȑa<�a<+�a<g�a<��a<ˑa<�a<F�a<��a<��a<�a<U�a<��a<�a<=�a<��a<�a<8�a<��a<��a<>�a<��a<�a<s�a<ݗa<<�a<��a<
�a<{�a<�a<R�a<��a<*�a<��a< �a<x�a<�a<^�a<ѝa<4�a<��a<6�a<��a<�a<��a<��a<\�a<ӡa<?�a<��a<�a<��a<��a<_�a<ʤa<.�a<��a<�a<\�a<��a<&�a<��a<ŧa<,�a<��a<�a<,�a<u�a<ǩa<�a<d�a<��a<��a<<�a<{�a<��a<��a<7�a<p�a<��a<Ӭa<��a<I�a<o�a<��a<��a<��a<�a<7�a<S�a<u�a<��a<��a<ήa<�a<��a<�a<�a<;�a<G�a<G�a<W�a<s�a<g�a<f�a<z�a<v�a<}�a<w�a<k�a<q�a<l�a<^�a<c�a<I�a<C�a<4�a<�a<�a<�a<�a<Ӯa<��a<��a<��a<a�a<?�a<(�a<�a<֭a<��a<��a<l�a<E�a<�a<�a<��a<��a<X�a<�a<��a<��a<v�a<C�a<�a<��a<�a<B�a<�a<Ʃa<y�a<#�a<�a<��a<O�a<�a<��a<]�a<�a<��a<[�a<�a<��a<Q�a<�a<��a<D�a<ңa<t�a<�a<��a<C�a<�a<x�a<�a<��a<=�a<ڟa<l�a<�a<��a<.�a<ʝa<U�a<�a<��a<�a<��a<=�a<Қa<q�a<�a<��a</�a<Ϙa<k�a<�a<��a<K�a<�a<��a<.�a<ڕa<��a<#�a<Δa<r�a<?�a<�a<��a<N�a<�a<a<��a<?�a<�a<ϑa<��a<_�a<(�a<��a<͐a<��a<��a<]�a<.�a<�a<�a<ߏa<Ïa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<Ïa<�a<�a<�  �  �a<I�a<F�a<~�a<��a<��a<�a<�a<i�a<��a<Ցa<�a<;�a<��a<��a<�a<D�a<��a<�a<4�a<��a<Ӕa<S�a<��a<��a<A�a<��a<�a<a�a<��a<)�a<��a<��a<u�a<�a<A�a<͚a<�a<��a<�a<t�a<�a<T�a<�a<,�a<ʞa<�a<��a<�a<t�a<��a<P�a<�a<-�a<��a<�a<��a<�a<I�a<ڤa< �a<��a<�a<V�a<Ǧa<	�a<��a<��a<<�a<}�a<ըa<+�a<r�a<ߩa<�a<t�a<��a<��a<>�a<j�a<ͫa<�a<;�a<a�a<��a<٬a<��a<M�a<R�a<��a<��a<�a<�a<0�a<b�a<c�a<��a<��a<Үa<߮a<�a<�a<�a<>�a</�a<[�a<S�a<Y�a<u�a<^�a<��a<d�a<��a<k�a<z�a<s�a<Y�a<r�a<D�a<Y�a<6�a<1�a<-�a<�a<
�a<Ԯa<�a<��a<��a<��a<X�a<Y�a<�a<�a<έa<ŭa<��a<b�a<J�a<�a<��a<��a<��a<V�a<�a<�a<��a<��a<+�a<�a<��a<��a<N�a<�a<ɩa<f�a<?�a<٨a<��a<T�a<�a<��a<I�a<�a<��a<W�a<�a<��a<c�a<ݤa<��a<'�a<ڣa<t�a<�a<��a<7�a<��a<g�a<�a<��a<9�a<�a<W�a<�a<��a<+�a<��a<N�a<��a<k�a<(�a<��a<L�a<͚a<g�a<�a<��a<H�a<��a<{�a< �a<��a<M�a<ٖa<��a<�a<ޕa<s�a<,�a<Ԕa<r�a<C�a<̓a<��a<A�a<�a<��a<~�a<N�a<�a<ۑa<��a<d�a<&�a<�a<ِa<��a<��a<E�a<B�a<�a<�a<�a<��a<ҏa<��a<��a<��a<��a<��a<{�a<��a<��a<��a<��a<��a<׏a<ҏa<�a<�  �  �a</�a<S�a<��a<��a<Ða<��a<)�a<e�a<��a<��a<�a<G�a<��a<ђa<�a<X�a<��a<�a<=�a<��a<�a<A�a<��a<�a<\�a<��a<�a<x�a<ޗa<4�a<��a<	�a<t�a<�a<J�a<��a<*�a<��a<�a<{�a<��a<_�a<ɝa<I�a<a<�a<��a<�a<��a<�a<]�a<ǡa<A�a<��a<!�a<��a<��a<]�a<��a<'�a<��a<��a<X�a<��a<�a<��a<ݧa<(�a<��a<�a</�a<��a<ϩa<�a<i�a<��a<�a<7�a<y�a<��a<�a<9�a<u�a<��a<լa<�a<@�a<]�a<��a<��a<�a<�a<*�a<Q�a<v�a<��a<��a<ʮa<�a<��a<�a<"�a<<�a<C�a<M�a<S�a<T�a<y�a<r�a<q�a<v�a<��a<t�a<y�a<j�a<i�a<h�a<P�a<T�a<C�a<.�a<$�a<�a<	�a<�a<̮a<��a<��a<w�a<]�a<H�a<&�a<�a<�a<��a<��a<m�a<;�a<�a<�a<��a<��a<J�a<�a<�a<��a<�a<4�a<�a<Ԫa<��a<@�a<
�a<ǩa<p�a<0�a<�a<��a<P�a<��a<��a<\�a<	�a<��a<]�a<�a<��a<I�a<��a<��a<'�a<ѣa<n�a<�a<��a<C�a<ءa<{�a<�a<��a<D�a<֟a<j�a<��a<��a<+�a<ŝa<Q�a<�a<o�a<�a<��a<8�a<֚a<w�a<�a<��a<7�a<јa<q�a<�a<��a<F�a<�a<��a<*�a<ݕa<��a<'�a<єa<��a<6�a<֓a<��a<N�a<�a<��a<w�a<=�a<�a<Ǒa<��a<[�a</�a<��a<��a<��a<��a<Y�a<5�a<�a<�a<�a<Ϗa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<Ώa<ُa<�a<�  �   �a<,�a<X�a<q�a<��a<ܐa<�a<?�a<G�a<��a<ˑa<
�a<I�a<w�a<ܒa<��a<f�a<��a<��a<B�a<��a<��a<(�a<��a<�a<P�a<��a<�a<y�a<ʗa<K�a<��a<�a<s�a<�a<g�a<��a<1�a<��a<�a<�a<�a<l�a<ǝa<J�a<��a<5�a<��a<�a<��a<ݠa<t�a<ša<V�a<��a<�a<��a<�a<t�a<��a<B�a<��a<�a<b�a<��a<,�a<f�a<ۧa<&�a<��a<ڨa<-�a<��a<��a<#�a<\�a<êa<��a<3�a<��a<��a<�a<)�a<q�a<��a<Ԭa<�a<-�a<��a<��a<ԭa<�a<�a<B�a<O�a<��a<~�a<��a<®a<�a<�a<
�a<2�a<�a<W�a<C�a<d�a<f�a<_�a<x�a<n�a<��a<m�a<��a<r�a<f�a<r�a<T�a<w�a<C�a<F�a<.�a<�a<�a<�a<�a<ɮa<��a<��a<��a<v�a<4�a<;�a<�a<�a<��a<��a<o�a<2�a<(�a<Ҭa<Ǭa<��a<`�a<#�a<߫a<ɫa<f�a<X�a<��a<Ǫa<��a<B�a<�a<��a<��a< �a<�a<��a<O�a<�a<��a<d�a<��a<��a<a�a< �a<��a<G�a<��a<��a<D�a<ңa<r�a<!�a<��a<Z�a<աa<��a<�a<��a<E�a<a<��a<��a<��a<�a<ʝa<[�a<��a<��a<�a<��a<7�a<��a<k�a<�a<��a< �a<٘a<c�a<�a<��a<B�a<�a<w�a<@�a<͕a<��a<*�a<Дa<��a<#�a<��a<��a<b�a<�a<��a<��a<;�a<�a<��a<��a<S�a<'�a<�a<ɐa<��a<g�a<m�a<*�a<!�a<��a<׏a<ԏa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<Ïa<�a<�a<�  �  �a<2�a<R�a<~�a<��a<ΐa<�a<2�a<N�a<��a<ʑa<��a<A�a<��a<̒a<�a<Q�a<��a<�a<?�a<��a<�a</�a<��a<�a<S�a<��a<�a<n�a<Зa<6�a<��a<�a<u�a<יa<H�a<��a</�a<��a<�a<|�a<�a<c�a<ϝa<F�a<��a< �a<��a<�a<��a<�a<e�a<ša<9�a<��a<!�a<��a<��a<Y�a<��a<2�a<��a<��a<_�a<��a<�a<v�a<اa<+�a<��a<֨a<.�a<�a<٩a< �a<a�a<��a<�a<6�a<��a<ëa<��a</�a<j�a<��a<Ѭa<�a<8�a<i�a<��a<̭a<�a<�a<6�a<J�a<q�a<��a<��a<Ѯa<�a<�a<	�a<$�a<&�a<H�a<H�a<X�a<a�a<n�a<n�a<s�a<}�a<s�a<v�a<t�a<��a<p�a<V�a<X�a<B�a<F�a<A�a<#�a<�a<��a<�a<Ϯa<��a<��a<��a<h�a<<�a<.�a<��a<�a<��a<��a<h�a<G�a<�a<�a<��a<z�a<W�a< �a<�a<��a<m�a<B�a<��a<˪a<~�a<H�a< �a<��a<r�a<7�a<�a<��a<C�a<��a<��a<b�a<�a<��a<^�a<�a<��a<O�a<��a<��a<.�a<ͣa<t�a<�a<��a<L�a<աa<s�a<�a<��a<D�a<ڟa<f�a<��a<��a<$�a<��a<X�a<�a<w�a<�a<��a<<�a<֚a<h�a<�a<��a<A�a<טa<h�a<�a<��a<F�a<�a<��a<.�a<ӕa<|�a<+�a<͔a<��a<.�a<�a<��a<Z�a<�a<��a<��a<5�a<��a<ёa<��a<b�a<(�a<�a<Ȑa<��a<p�a<^�a</�a<�a<��a<�a<ʏa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ȏa<͏a<ߏa<��a<�  �  �a<7�a<C�a<��a<��a<Ӑa<��a<�a<i�a<��a<ϑa<�a<:�a<��a<��a<�a<E�a<��a<�a<B�a<��a<ٔa<K�a<��a<��a<N�a<��a<�a<f�a<�a<�a<��a<��a<x�a<�a<D�a<њa<�a<��a<��a<z�a<�a<X�a<Нa<5�a<��a<&�a<��a<�a<z�a<�a<T�a<�a<:�a<��a<
�a<r�a<��a<R�a<�a<!�a<��a<��a<Y�a<Ѧa<�a<��a<Ƨa<'�a<}�a<Ҩa<4�a<l�a<ԩa<�a<y�a<��a<��a<B�a<h�a<īa<�a<C�a<c�a<��a<̬a<�a<E�a<k�a<��a<��a<�a<�a<*�a<s�a<e�a<��a<��a<Ȯa<ޮa<�a<�a<�a<A�a<4�a<P�a<c�a<h�a<v�a<]�a<w�a<t�a<~�a<h�a<n�a<p�a<_�a<w�a<J�a<`�a<9�a<,�a<!�a<��a<�a<�a<Ԯa<��a<��a<��a<m�a<L�a<�a<�a<ۭa<��a<��a<`�a<A�a<��a<�a<��a<��a<N�a<#�a<�a<��a<��a<C�a<�a<ƪa<w�a<M�a<��a<̩a<\�a<8�a<ըa<��a<V�a<��a<ħa<I�a<�a<��a<]�a<�a<��a<O�a<�a<��a<5�a<�a<s�a<�a<��a<:�a<��a<t�a<�a<��a<)�a<۟a<`�a<�a<��a<;�a<��a<R�a<��a<{�a<�a<��a<8�a<̚a<d�a<�a<��a<<�a<��a<��a<�a<��a<R�a<֖a<��a<�a<�a<u�a<+�a<ǔa<{�a<;�a<�a<��a<E�a<
�a<ɒa<w�a<^�a<�a<ԑa<x�a<Z�a<%�a<�a<֐a<��a<��a<J�a<7�a<!�a<�a<�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ˏa<Ώa<�a<�  �  �a<<�a<Z�a<t�a<��a<ΐa<�a<(�a<]�a<��a<��a<�a<5�a<��a<ϒa<�a<D�a<��a<�a<C�a<��a<�a<5�a<��a<�a<Q�a<��a<�a<d�a<՗a<>�a<��a<�a<s�a<әa<?�a<��a<,�a<��a<�a<�a<ܜa<b�a<ߝa<N�a<��a<+�a<��a<�a<x�a<��a<X�a<ϡa<9�a<��a<(�a<��a<��a<U�a<Ťa<#�a<��a<�a<V�a<��a< �a<m�a<ߧa<:�a<��a<ʨa<3�a<��a<ةa<�a<e�a<��a<�a<9�a<{�a<ȫa<��a<9�a<_�a<��a<�a<�a<3�a<r�a<��a<��a<�a<�a<&�a<V�a<e�a<��a<��a<خa<׮a<��a<�a<!�a<5�a<A�a<H�a<Y�a<a�a<e�a<w�a<�a<w�a<m�a<{�a<~�a<x�a<i�a<a�a<F�a<J�a<>�a<9�a<.�a<�a<�a<�a<ٮa<��a<��a<|�a<g�a<?�a<%�a<�a<�a<��a<��a<[�a<N�a<�a<��a<��a<��a<F�a<$�a<�a<��a<s�a<H�a<��a<Ȫa<��a<Q�a<��a<��a<{�a<?�a<�a<��a<@�a<�a<��a<_�a<�a<��a<b�a<��a<��a<^�a<��a<��a<9�a<Уa<m�a<
�a<��a<?�a<�a<r�a<�a<��a<K�a<֟a<c�a<��a<��a<0�a<��a<O�a<�a<��a<�a<��a<K�a<ښa<[�a<	�a<��a<@�a<՘a<l�a<��a<��a<H�a<�a<��a<7�a<ܕa<q�a<4�a<��a<��a<)�a<�a<��a<N�a<�a<ƒa<t�a<B�a<�a<Ցa<��a<i�a<�a<��a<a<��a<~�a<W�a</�a<�a<��a<ݏa<ӏa<ďa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<؏a<�a<��a<�  �  �a<�a<E�a<r�a<n�a<ʐa<ΐa<�a</�a<z�a<��a<��a<?�a<U�a<��a<�a<M�a<��a<˓a<$�a<e�a<Δa<�a<��a<��a<N�a<��a<�a<p�a<��a<7�a<��a<��a<^�a<��a<:�a<��a<"�a<t�a<�a<k�a<ޜa<S�a<��a<<�a<��a<�a<��a<�a<d�a<ʠa<E�a<��a<=�a<��a<��a<i�a<ݣa<[�a<��a<�a<p�a<ޥa<A�a<��a<�a<L�a<ѧa<
�a<y�a<بa<�a<��a<��a<�a<@�a<��a<֪a<�a<r�a<��a<��a<�a<m�a<��a<ìa<�a<�a<p�a<r�a<��a<ŭa<�a<�a<>�a<r�a<t�a<��a<��a<�a<��a<�a<�a<	�a<'�a<*�a<Y�a<=�a<_�a<h�a<L�a<}�a<U�a<y�a<t�a<Q�a<b�a<@�a<O�a<(�a<6�a<�a<�a<�a<Ԯa<�a<��a<��a<��a<V�a<j�a<!�a<�a<ܭa<έa<��a<��a<k�a<�a<�a<Ŭa<��a<y�a<6�a<�a<īa<��a<T�a<I�a<ͪa<˪a<z�a<�a<�a<��a<x�a<�a<٨a<��a<*�a<�a<��a<X�a<�a<��a<Q�a<��a<��a<&�a<�a<p�a<"�a<ȣa<T�a<��a<��a<,�a<��a<v�a<�a<��a<�a<��a<g�a<ݞa<|�a<�a<��a<7�a<Мa<r�a<�a<��a<�a<Śa<e�a<�a<��a<�a<Ęa<C�a<�a<��a<)�a<ۖa<n�a<.�a<��a<y�a<�a<��a<��a<��a<�a<n�a<4�a<ݒa<��a<_�a<#�a<��a<��a<h�a<+�a<!�a<�a<��a<��a<L�a<6�a<�a<�a<Ώa<яa<��a<��a<��a<u�a<��a<��a<f�a<}�a<f�a<��a<r�a<��a<��a<��a<ݏa<ʏa<�  �  ��a<�a<9�a<f�a<��a<��a<ܐa<�a<D�a<w�a<��a<ߑa<�a<u�a<��a<�a<*�a<��a<דa<-�a<��a<ܔa<�a<��a<Օa<6�a<��a<��a<U�a<��a<�a<��a<�a<g�a<ҙa<=�a<��a<�a<{�a<�a<Z�a<Μa<C�a<��a<+�a<��a<�a<��a<��a<z�a<�a<K�a<ša<�a<��a<�a<|�a<�a<9�a<��a<�a<��a<��a<P�a<��a<�a<i�a<��a<�a<m�a<��a<�a<b�a<��a<
�a<T�a<��a<�a<,�a<h�a<��a<ګa<�a<R�a<��a<Ĭa<��a<%�a<W�a<z�a<��a<�a<�a<!�a<C�a<P�a<��a<��a<®a<Ůa<Ԯa<�a<�a<#�a<8�a<;�a<I�a<I�a<`�a<[�a<f�a<_�a<`�a<`�a<V�a<W�a<X�a<L�a<E�a<<�a<2�a<�a<�a<��a<�a<Юa<��a<��a<��a<h�a<T�a</�a<�a<�a<ʭa<��a<r�a<I�a<7�a<�a<�a<��a<r�a<A�a<�a<߫a<��a<]�a</�a<�a<��a<r�a<6�a<�a<��a<[�a<�a<Шa<��a<C�a<�a<��a<K�a<�a<��a<@�a<�a<��a<>�a<ޤa<��a< �a<ģa<e�a<�a<��a<2�a<աa<Q�a<��a<��a<2�a<��a<E�a<�a<��a<#�a<��a<F�a<ќa<e�a< �a<��a<)�a<��a<M�a<�a<{�a<�a<��a<V�a<��a<��a<6�a<іa<k�a<�a<��a<^�a<�a<��a<i�a<�a<˓a<u�a<C�a<��a<��a<h�a<(�a<ؑa<��a<�a<M�a<�a<ΐa<��a<��a<f�a<H�a<�a< �a<ۏa<ҏa<��a<��a<��a<��a<w�a<j�a<l�a<s�a<r�a<{�a<��a<��a<��a<��a<��a<܏a<�  �  ߏa<9�a<.�a<[�a<��a<��a<�a<�a<G�a<[�a<��a<�a<�a<��a<��a<�a<*�a<��a<ϓa<�a<u�a<Ôa<*�a<j�a<�a<'�a<��a<�a<D�a<ڗa<�a<��a<�a<X�a<Ιa<+�a<��a< �a<��a<�a<s�a<�a<?�a<ѝa<�a<��a<�a<��a<�a<X�a<ܠa<-�a<ҡa<�a<��a<�a<m�a<�a<7�a<ɤa< �a<��a<եa<A�a<��a<��a<{�a<��a<1�a<s�a<Ϩa</�a<e�a<ͩa<��a<W�a<��a<�a<#�a<]�a<��a<ګa<9�a<L�a<��a<άa<�a<@�a<C�a<��a<��a<ͭa<�a<�a<T�a<L�a<��a<��a<Ǯa<ɮa<߮a<�a<�a<%�a<�a<=�a<;�a<S�a<\�a<K�a<��a<K�a<��a<f�a<f�a<l�a<D�a<X�a<:�a<C�a<�a<(�a<�a<��a<
�a<��a<ܮa<��a<��a<y�a<B�a<6�a<�a<��a<��a<��a<~�a<J�a<B�a<�a<�a<��a<��a<:�a<��a<ӫa<��a<l�a<�a<�a<��a<s�a<K�a<کa<ȩa<\�a</�a<Ψa<��a<>�a<�a<��a<7�a<�a<��a<X�a< �a<��a<S�a<Ĥa<��a<�a<��a<\�a<�a<��a<�a<�a<U�a<
�a<��a<$�a<џa<C�a<�a<f�a<�a<��a<7�a<Ԝa<U�a<�a<x�a<>�a<��a<\�a<�a<�a<0�a<��a<Y�a<�a<��a<-�a<ǖa<��a<�a<וa<X�a<!�a<Ĕa<V�a<0�a<��a<��a<-�a<�a<��a<X�a<9�a<ԑa<a<]�a<R�a<	�a<ِa<Őa<j�a<h�a<-�a<�a<�a<�a<Ώa<��a<��a<x�a<��a<}�a<z�a<��a<_�a<~�a<o�a<��a<��a<��a<��a<Ïa<�a<�  �  �a<�a<;�a<d�a<}�a<��a<�a<�a<V�a<w�a<��a<�a<(�a<k�a<��a<��a<;�a<��a<ʓa</�a<��a<Ɣa<-�a<x�a<ѕa<;�a<��a<�a<R�a<��a<�a<��a<�a<^�a<͙a<6�a<��a<�a<�a<�a<W�a<؜a<<�a<��a<+�a<��a<�a<��a<��a<c�a<�a<F�a<��a<2�a<��a< �a<k�a<�a<M�a<��a<�a<��a<ߥa<G�a<��a<�a<i�a<��a<�a<g�a<Ǩa<�a<f�a<��a<�a<Y�a<��a<�a<'�a<a�a<��a<۫a<�a<V�a<��a<Ƭa<��a<$�a<S�a<��a<��a<حa<�a<�a<F�a<a�a<��a<��a<��a<Ϯa<�a<�a<
�a<4�a<%�a<B�a<B�a<H�a<\�a<[�a<d�a<[�a<g�a<V�a<g�a<T�a<R�a<X�a<H�a<@�a<'�a<�a<�a<�a<�a<ʮa<��a<��a<��a<e�a<L�a<:�a<�a<�a<˭a<��a<��a<U�a<-�a<�a<֬a<��a<z�a<5�a<�a<�a<��a<p�a<'�a<�a<��a<u�a<*�a<�a<��a<X�a<�a<˨a<��a<=�a<�a<��a<G�a<�a<��a<=�a<��a<��a<=�a<ޤa<��a<�a<ţa<c�a<��a<��a<-�a<ǡa<l�a<�a<��a<"�a<ȟa<Y�a<�a<{�a<#�a<��a<=�a<לa<d�a< �a<��a<*�a<��a<U�a<��a<��a<�a<��a<\�a<�a<��a<1�a<ʖa<v�a<�a<��a<b�a<�a<��a<k�a<�a<Ɠa<��a<2�a<�a<��a<]�a<+�a<�a<��a<c�a<>�a<�a<�a<��a<��a<w�a<4�a<#�a<��a<ُa<͏a<��a<��a<��a<��a<m�a<{�a<i�a<m�a<~�a<}�a<��a<��a<��a<��a<��a<�a<�  �  �a<
�a<?�a<a�a<�a<��a<ڐa<�a<+�a<�a<��a<�a<�a<g�a<ʒa<�a<9�a<|�a<ԓa<'�a<l�a<Дa<�a<��a<͕a<=�a<��a<�a<t�a<��a<1�a<��a<�a<c�a<ęa<7�a<��a<#�a<r�a< �a<W�a<ܜa<R�a<��a<<�a<��a<�a<��a<��a<g�a<ɠa<Z�a<��a<.�a<��a<�a<��a<ңa<N�a<��a<&�a<s�a<�a<H�a<��a<�a<Z�a<ѧa<�a<w�a<Өa<
�a<{�a<��a<�a<F�a<��a<ݪa<&�a<k�a<��a<��a<�a<q�a<��a<��a<�a<�a<g�a<u�a<��a<˭a<��a<#�a<4�a<a�a<y�a<��a<��a<îa<�a<�a<�a<�a<-�a<:�a<I�a<O�a<T�a<f�a<S�a<y�a<a�a<c�a<e�a<M�a<h�a<9�a<E�a<*�a<;�a<�a<�a<�a<�a<�a<��a<��a<��a<g�a<W�a<.�a<�a<حa<ӭa<��a<w�a<L�a<(�a<�a<ͬa<��a<g�a<?�a<�a<˫a<��a<[�a<;�a<�a<��a<s�a<'�a<�a<��a<r�a<�a<Шa<��a<5�a<�a<��a<Z�a<�a<��a<<�a<��a<��a</�a<�a<v�a<-�a<��a<_�a<��a<��a<B�a<��a<g�a<�a<��a<;�a<��a<Z�a<ߞa<��a<�a<��a<?�a<Ȝa<u�a<�a<��a<�a<Úa<`�a<ܙa<��a<�a<Ƙa<H�a<�a<��a<0�a<Ֆa<f�a<'�a<��a<~�a<�a<��a<t�a<
�a<ۓa<p�a<8�a<�a<��a<j�a<�a<�a<��a<��a<B�a<�a<ܐa<��a<��a<H�a<=�a<�a< �a<�a<Əa<��a<��a<��a<��a<z�a<y�a<c�a<��a<_�a<{�a<s�a<��a<��a<��a<͏a<ڏa<�  �  �a<�a<>�a<Y�a<��a<��a<֐a<�a<9�a<z�a<��a<�a<1�a<b�a<��a<�a<B�a<��a<��a<"�a<t�a<ؔa<�a<|�a<��a<,�a<��a<��a<K�a<��a<'�a<��a<��a<T�a<��a<<�a<��a<�a<�a<��a<a�a<͜a<?�a<��a<)�a<��a<�a<��a<��a<o�a<ՠa<N�a<¡a<,�a<��a<��a<h�a<ݣa<K�a<��a<�a<}�a<�a<L�a<��a<�a<c�a<��a<�a<n�a<��a<�a<r�a<��a<
�a<E�a<��a<ܪa<�a<l�a<��a<�a<�a<K�a<��a<ˬa<�a<+�a<V�a<~�a<��a<ӭa<��a<(�a<G�a<d�a<x�a<��a<��a<׮a<�a<�a<�a<�a<5�a<4�a<E�a<X�a<U�a<_�a<e�a<W�a<\�a<h�a<e�a<_�a<\�a<B�a<W�a<-�a<+�a<#�a<�a<�a<ݮa<Ůa<��a<��a<��a<w�a<O�a<)�a<�a<�a<έa<��a<��a<^�a<#�a<�a<ʬa<��a<y�a<K�a<	�a<ҫa<��a<`�a<+�a<��a<��a<|�a<3�a<�a<��a<h�a<!�a<٨a<}�a<1�a<�a<��a<K�a<�a<��a<F�a<�a<��a<<�a<ܤa<�a<(�a<£a<a�a<�a<��a<5�a<ҡa<e�a<��a<��a<�a<��a<X�a<�a<��a<�a<��a<C�a<ќa<k�a<��a<��a<&�a<��a<K�a<�a<��a<�a<��a<G�a<�a<��a<'�a<Ֆa<x�a<�a<��a<X�a<�a<��a<_�a<�a<ʓa<z�a<=�a<�a<��a<o�a<,�a<�a<��a<c�a<8�a<�a<ߐa<��a<��a<X�a<E�a<�a<��a<�a<Əa<��a<��a<��a<|�a<��a<x�a<t�a<w�a<h�a<��a<w�a<��a<��a<��a<͏a<ԏa<�  �  �a<"�a<4�a<a�a<��a<��a<�a<�a<N�a<n�a<��a<�a<*�a<p�a<��a<��a<:�a<��a<̓a<'�a<��a<Ôa<3�a<o�a<�a<.�a<��a<��a<O�a<ϗa<�a<��a<�a<d�a<˙a<3�a<��a<�a<��a<�a<k�a<՜a<>�a<ɝa<�a<��a<�a<��a<��a<b�a<�a<=�a<��a<"�a<��a<�a<s�a<�a<B�a<��a<�a<��a<ߥa<B�a<��a<��a<q�a<��a<'�a<k�a<èa<'�a<_�a<��a<�a<a�a<��a<�a<-�a<_�a<��a<իa<3�a<Q�a<��a<̬a<�a<5�a<H�a<��a<��a<حa< �a<�a<B�a<]�a<��a<��a<��a<ծa<�a<��a< �a</�a<#�a<?�a<J�a<I�a<^�a<Q�a<n�a<Y�a<n�a<b�a<W�a<Z�a<T�a<V�a<B�a<?�a<,�a<�a<�a<��a<�a<Ǯa<Ʈa<��a<��a<m�a<O�a<:�a<�a<��a<­a<��a<{�a<W�a<1�a<��a<ܬa<��a<q�a<6�a<�a<߫a<��a<v�a<�a<��a<��a<y�a<5�a<�a<��a<U�a<�a<Ψa<��a<<�a<�a<��a<C�a<��a<��a<P�a<�a<��a<L�a<Ѥa<��a<�a<ʣa<^�a<��a<��a<$�a<ϡa<\�a<�a<��a<)�a<ϟa<O�a<�a<t�a<%�a<��a<8�a<ޜa<[�a<�a<��a<4�a<��a<P�a<��a<y�a<#�a<��a<d�a<�a<��a<7�a<ɖa<u�a<�a<Еa<^�a<�a<a<]�a<%�a<��a<��a<,�a<�a<��a<\�a<'�a<�a<��a<t�a<F�a<�a<ܐa<��a<{�a<r�a<3�a< �a<�a<ۏa<Ϗa<��a<��a<��a<��a<y�a<k�a<o�a<o�a<|�a<x�a<��a<��a<��a<��a<��a<�a<�  �  �a<�a<8�a<i�a<�a<��a<�a< �a<6�a<~�a<��a<�a<$�a<_�a<��a<�a<C�a<��a<ۓa<)�a<q�a<��a<&�a<~�a<֕a<?�a<��a<�a<_�a<��a<'�a<��a<�a<d�a<��a<#�a<��a<�a<��a<��a<`�a<՜a<N�a<��a<.�a<��a<	�a<��a<��a<]�a<Ѡa<Q�a<��a<0�a<��a<�a<u�a<ԣa<M�a<��a<!�a<x�a<ۥa<E�a<��a<�a<c�a<ŧa<�a<v�a<˨a<�a<o�a<��a<�a<M�a<��a<تa<(�a<g�a<��a<�a<�a<`�a<��a<Ŭa<��a<&�a<T�a<��a<��a<έa<��a<&�a<@�a<f�a<s�a<��a<��a<Ʈa<�a<�a<�a<�a< �a<<�a<O�a<F�a<`�a<[�a<Z�a<q�a<_�a<`�a<k�a<b�a<]�a<G�a<2�a<1�a<3�a< �a<�a<��a<�a<߮a<��a<��a<��a<f�a<V�a<6�a<�a<�a<ҭa<��a<��a<P�a< �a<�a<Ƭa<��a<t�a<F�a<�a<ϫa<��a<i�a<-�a<�a<��a<s�a<.�a<��a<��a<h�a<#�a<Ҩa<��a<0�a<اa<��a<J�a<��a<��a<E�a<�a<��a<7�a<�a<��a<�a<ţa<^�a<�a<��a<8�a<ѡa<i�a<��a<��a<+�a<��a<Y�a<�a<��a<�a<��a<;�a<Ҝa<a�a<��a<��a<$�a<a<X�a<�a<��a<%�a<��a<O�a<�a<��a<2�a<Жa<y�a<�a<��a<l�a<�a<��a<p�a<�a<ȓa<��a<,�a<�a<��a<m�a<%�a<�a<��a<��a<8�a<�a<�a<��a<��a<T�a<0�a<�a<�a<؏a<ҏa<��a<��a<��a<�a<x�a<�a<w�a<x�a<l�a<g�a<{�a<��a<��a<��a<Ǐa<؏a<�  �  ��a<�a<D�a<V�a<��a<��a<Аa<'�a<<�a<��a<��a<�a<5�a<^�a<��a<ޒa<O�a<y�a<ޓa<"�a<w�a<��a<�a<��a<ӕa<9�a<��a<��a<X�a<��a<0�a<�a<�a<P�a<̙a<O�a<��a<�a<s�a<��a<^�a<˜a<I�a<��a<>�a<��a<�a<�a<�a<~�a<͠a<[�a<��a<2�a<��a<�a<s�a<أa<V�a<��a<,�a<p�a<��a<J�a<��a<�a<X�a<Чa<�a<r�a<��a<�a<u�a<��a<
�a<F�a<��a<�a<�a<g�a<��a<��a<�a<X�a<��a<Ĭa<�a<�a<e�a<u�a<��a<٭a<�a<,�a<2�a<s�a<m�a<��a<��a<׮a<�a<�a<�a<�a<I�a</�a<H�a<V�a<M�a<j�a<W�a<g�a<V�a<g�a<]�a<Q�a<P�a<I�a<`�a<6�a<#�a<�a<�a<�a<ծa<֮a<��a<��a<��a<r�a<U�a<$�a<*�a<�a<ԭa<��a<v�a<a�a< �a<�a<��a<��a<c�a<H�a<	�a<իa<��a<Y�a<8�a<�a<��a<t�a<3�a<�a<��a<q�a<�a<Шa<y�a<=�a<�a<��a<I�a<�a<��a<D�a<�a<��a<-�a<�a<s�a<.�a<��a<[�a<�a<��a<B�a<��a<l�a<��a<��a<)�a<��a<b�a<۞a<��a<�a<��a<A�a<ǜa<w�a<�a<��a<�a<��a<N�a<�a<��a<�a<��a<I�a<�a<��a< �a<іa<g�a<(�a<��a<e�a<�a<��a<q�a<�a<ٓa<q�a<B�a<�a<��a<s�a<�a<��a<��a<y�a<<�a<�a<ܐa<��a<��a<Y�a<Y�a<�a<��a<�a<��a<��a<��a<��a<v�a<~�a<q�a<f�a<k�a<o�a<��a<�a<��a<��a<��a<̏a<̏a<�  �  �a<"�a<5�a<V�a<��a<��a<ސa<�a<D�a<g�a<��a<�a<&�a<p�a<��a<��a<9�a<��a<ۓa<�a<{�a<Ĕa<&�a<z�a<ܕa<.�a<��a<��a<Q�a<җa<�a<��a<��a<^�a<řa<#�a<��a<�a<��a<�a<p�a<՜a<E�a<��a<)�a<��a<�a<��a<�a<f�a<Ԡa<C�a<��a<&�a<��a<�a<s�a<�a<F�a<��a<�a<v�a<�a<<�a<��a<�a<g�a<��a< �a<p�a<¨a<'�a<e�a<��a<	�a<Y�a<��a<ڪa<)�a<p�a<��a<߫a<1�a<S�a<��a<Ǭa<�a<,�a<U�a<��a<��a<حa<�a<�a<=�a<`�a<��a<��a<��a<Ϯa<�a<��a< �a<�a<'�a<5�a<H�a<V�a<O�a<X�a<l�a<\�a<q�a<k�a<T�a<d�a<U�a<R�a<+�a<<�a<+�a<%�a<�a<��a<��a<ʮa<Ʈa<��a<��a<t�a<Q�a<2�a<	�a<�a<��a<��a<x�a<R�a<2�a<�a<ݬa<��a<k�a<E�a< �a<٫a<��a<i�a<)�a<��a<��a<p�a<9�a<�a<��a<_�a<�a<ܨa<��a<5�a<اa<��a<I�a<��a<��a<V�a<�a<��a<B�a<ܤa<�a<"�a<ãa<U�a<��a<��a<*�a<ϡa<_�a< �a<��a<*�a<ǟa<R�a<�a<{�a<�a<��a<2�a<՜a<g�a<��a<��a<-�a<��a<O�a<��a<~�a<�a<��a<[�a<�a<��a<3�a<ٖa<m�a<�a<ϕa<`�a<�a<��a<c�a<�a<ɓa<��a<)�a<�a<��a<f�a<"�a<�a<��a<x�a<F�a<�a<ڐa<��a<{�a<b�a<6�a<�a<��a<�a<��a<��a<��a<��a<��a<��a<h�a<y�a<p�a<x�a<a�a<��a<��a<��a<��a<ɏa<�a<�  �  �a<�a<*�a<n�a<��a<��a<��a<�a<d�a<s�a<��a<�a<�a<t�a<��a<��a<*�a<��a<ۓa<,�a<��a<��a<@�a<i�a<�a<4�a<��a<��a<G�a<ėa<�a<��a<�a<\�a<֙a< �a<��a<��a<��a<��a<]�a<˜a<@�a<��a<�a<��a<��a<��a<�a<`�a<�a<A�a<Сa<�a<��a<�a<m�a<�a<;�a<Ǥa<�a<��a<�a<N�a<��a<�a<|�a<��a<�a<j�a<��a<�a<S�a<ϩa<�a<b�a<��a<�a<-�a<X�a<��a<ūa<$�a<G�a<��a<¬a<�a<8�a<=�a<��a<��a<�a<�a<!�a<S�a<O�a<��a<��a<��a<Ȯa<�a<�a<�a<=�a<�a<V�a<C�a<E�a<m�a<K�a<h�a<[�a<e�a<Q�a<_�a<j�a<D�a<i�a<&�a<R�a<�a<"�a<�a<�a<�a<Ǯa<��a<��a<��a<g�a<G�a<Q�a<��a<�a<ǭa<��a<��a<I�a<5�a<��a<ܬa<��a<��a<E�a<�a<�a<��a<��a<�a<��a<��a<k�a<3�a<ީa<��a<D�a</�a<Ȩa<��a<G�a<էa<��a<1�a<�a<��a<C�a<�a<��a<@�a<ˤa<��a<�a<ϣa<n�a<��a<��a<(�a<�a<Y�a<��a<��a<$�a<ğa<G�a<��a<y�a<,�a<��a<D�a<�a<O�a<�a<~�a<*�a<��a<F�a<�a<l�a<3�a<��a<d�a<�a<��a<8�a<a<��a<��a<a<S�a<�a<��a<a�a<(�a<��a<��a<(�a<�a<��a<h�a<8�a<בa<��a<l�a<H�a<�a<ސa<Őa<��a<��a<%�a<7�a<��a<֏a<ޏa<��a<��a<��a<��a<i�a<s�a<�a<_�a<��a<\�a<��a<��a<��a<��a<��a<�a<�  �  �a<�a<>�a<Z�a<��a<��a<�a<�a<?�a<q�a<��a<�a<1�a<p�a<��a<�a<>�a<��a<͓a<!�a<s�a<ɔa<(�a<|�a<�a<.�a<��a<��a<d�a<ėa<"�a<��a<ߘa<T�a<ԙa<>�a<��a<�a<��a<��a<n�a<�a<S�a<��a<+�a<��a<�a<��a<��a<a�a<Ҡa<B�a<��a<,�a<��a<�a<|�a<�a<L�a<��a<�a<x�a<ޥa<D�a<��a<�a<f�a<��a<�a<{�a<֨a<'�a<n�a<��a<��a<T�a<��a<�a<�a<Q�a<��a<�a<-�a<i�a<��a<Ȭa<��a<0�a<U�a<��a<��a<έa<�a<�a<:�a<c�a<}�a<��a<��a<ٮa<�a<�a<�a<�a<+�a<?�a<F�a<S�a<T�a<a�a<Y�a<s�a<l�a<i�a<b�a<Y�a<C�a<\�a<H�a<E�a<�a<�a<�a<��a<�a<�a<��a<��a<��a<t�a<P�a<6�a<�a<�a<ŭa<��a<x�a<^�a<1�a<�a<Ϭa<��a<m�a<7�a<�a<ҫa<��a<k�a<+�a<��a<��a<v�a<3�a<��a<��a<c�a<"�a<��a<}�a<D�a<�a<��a<7�a<��a<��a<T�a<��a<��a<4�a<ޤa<~�a<!�a<��a<]�a<��a<��a<)�a<ġa<f�a<�a<��a<3�a<ğa<X�a<�a<w�a<�a<��a<:�a<Ԝa<e�a<��a<��a<$�a<ǚa<c�a<��a<��a<$�a<��a<V�a<��a<��a<)�a<��a<{�a<�a<˕a<u�a<�a<��a<f�a<!�a<ɓa<��a<1�a<�a<��a<]�a<�a<�a<��a<|�a<J�a<�a<ܐa<��a<��a<_�a<;�a< �a<��a<�a<ŏa<��a<��a<��a<��a<��a<v�a<n�a<^�a<��a<}�a<��a<��a<��a<��a<Ǐa<�a<�  �  ��a<�a<V�a<E�a<��a<��a<Ɛa<-�a<-�a<��a<��a<�a<1�a<X�a<��a<�a<L�a<|�a<�a<;�a<n�a<�a<�a<��a<ڕa<'�a<��a<�a<S�a<��a<!�a<v�a< �a<m�a<��a<&�a<��a<#�a<y�a<�a<X�a<ǜa<D�a<��a<D�a<~�a<'�a<}�a<�a<~�a<Ϡa<c�a<��a<6�a<��a< �a<s�a<ѣa<T�a<��a<1�a<|�a<��a<J�a<��a<�a<H�a<Чa<�a<l�a<��a<
�a<e�a<��a<�a<K�a<��a<Ъa<.�a<w�a<��a<ޫa<�a<U�a<��a<άa<��a<�a<e�a<m�a<��a<حa<�a<5�a<3�a<s�a<l�a<��a<��a<Үa<�a< �a<!�a<�a<I�a<$�a<Q�a<j�a<7�a<{�a<P�a<f�a<R�a<e�a<T�a<e�a<i�a<@�a<5�a<&�a<A�a<'�a<��a<��a<Ԯa<Үa<��a<��a<p�a<��a<[�a<�a<0�a<ۭa<�a<��a<|�a<^�a<�a<�a<Ĭa<��a<f�a<V�a<!�a<ͫa<��a<Q�a<8�a<�a<��a<��a<"�a<�a<��a<b�a<�a<ߨa<��a<%�a<ۧa<��a<Y�a<�a<��a<=�a<�a<��a</�a<��a<`�a<7�a<��a<X�a<�a<��a<J�a<ơa<p�a<��a<��a<*�a<��a<`�a<�a<��a<�a<��a<@�a<Ɯa<x�a<ߛa<��a<"�a<��a<J�a<ܙa<~�a<�a<ʘa<M�a<�a<�a<8�a<�a<b�a<�a<��a<a�a<�a<Ĕa<e�a<�a<ؓa<h�a<D�a<�a<��a<|�a<�a<��a<��a<|�a<0�a<�a<�a<��a<��a<Q�a<X�a<�a<�a<��a<��a<яa<��a<��a<r�a<}�a<h�a<z�a<��a<f�a<k�a<p�a<��a<��a<��a<ɏa<ˏa<�  �  �a<�a<>�a<Z�a<��a<��a<�a<�a<?�a<q�a<��a<�a<1�a<p�a<��a<�a<>�a<��a<͓a<!�a<s�a<ɔa<(�a<|�a<�a<.�a<��a<��a<d�a<ėa<"�a<��a<ߘa<T�a<ԙa<>�a<��a<�a<��a<��a<n�a<�a<S�a<��a<+�a<��a<�a<��a<��a<a�a<Ҡa<B�a<��a<,�a<��a<�a<|�a<�a<L�a<��a<�a<x�a<ޥa<D�a<��a<�a<f�a<��a<�a<{�a<֨a<'�a<n�a<��a<��a<T�a<��a<�a<�a<Q�a<��a<�a<-�a<i�a<��a<Ȭa<��a<0�a<U�a<��a<��a<έa<�a<�a<:�a<c�a<}�a<��a<��a<ٮa<�a<�a<�a<�a<+�a<?�a<F�a<S�a<T�a<a�a<Y�a<s�a<l�a<i�a<b�a<Y�a<C�a<\�a<H�a<E�a<�a<�a<�a<��a<�a<�a<��a<��a<��a<t�a<P�a<6�a<�a<�a<ŭa<��a<x�a<^�a<1�a<�a<Ϭa<��a<m�a<7�a<�a<ҫa<��a<k�a<+�a<��a<��a<v�a<3�a<��a<��a<c�a<"�a<��a<}�a<D�a<�a<��a<7�a<��a<��a<T�a<��a<��a<4�a<ޤa<~�a<!�a<��a<]�a<��a<��a<)�a<ġa<f�a<�a<��a<3�a<ğa<X�a<�a<w�a<�a<��a<:�a<Ԝa<e�a<��a<��a<$�a<ǚa<c�a<��a<��a<$�a<��a<V�a<��a<��a<)�a<��a<{�a<�a<˕a<u�a<�a<��a<f�a<!�a<ɓa<��a<1�a<�a<��a<]�a<�a<�a<��a<|�a<J�a<�a<ܐa<��a<��a<_�a<;�a< �a<��a<�a<ŏa<��a<��a<��a<��a<��a<v�a<n�a<^�a<��a<}�a<��a<��a<��a<��a<Ǐa<�a<�  �  �a<�a<*�a<n�a<��a<��a<��a<�a<d�a<s�a<��a<�a<�a<t�a<��a<��a<*�a<��a<ۓa<,�a<��a<��a<@�a<i�a<�a<4�a<��a<��a<G�a<ėa<�a<��a<�a<\�a<֙a< �a<��a<��a<��a<��a<]�a<˜a<@�a<��a<�a<��a<��a<��a<�a<`�a<�a<A�a<Сa<�a<��a<�a<m�a<�a<;�a<Ǥa<�a<��a<�a<N�a<��a<�a<|�a<��a<�a<j�a<��a<�a<S�a<ϩa<�a<b�a<��a<�a<-�a<X�a<��a<ūa<$�a<G�a<��a<¬a<�a<8�a<=�a<��a<��a<�a<�a<!�a<S�a<O�a<��a<��a<��a<Ȯa<�a<�a<�a<=�a<�a<V�a<C�a<E�a<m�a<K�a<h�a<[�a<e�a<Q�a<_�a<j�a<D�a<i�a<&�a<R�a<�a<"�a<�a<�a<�a<Ǯa<��a<��a<��a<g�a<G�a<Q�a<��a<�a<ǭa<��a<��a<I�a<5�a<��a<ܬa<��a<��a<E�a<�a<�a<��a<��a<�a<��a<��a<k�a<3�a<ީa<��a<D�a</�a<Ȩa<��a<G�a<էa<��a<1�a<�a<��a<C�a<�a<��a<@�a<ˤa<��a<�a<ϣa<n�a<��a<��a<(�a<�a<Y�a<��a<��a<$�a<ğa<G�a<��a<y�a<,�a<��a<D�a<�a<O�a<�a<~�a<*�a<��a<F�a<�a<l�a<3�a<��a<d�a<�a<��a<8�a<a<��a<��a<a<S�a<�a<��a<a�a<(�a<��a<��a<(�a<�a<��a<h�a<8�a<בa<��a<l�a<H�a<�a<ސa<Őa<��a<��a<%�a<7�a<��a<֏a<ޏa<��a<��a<��a<��a<i�a<s�a<�a<_�a<��a<\�a<��a<��a<��a<��a<��a<�a<�  �  �a<"�a<5�a<V�a<��a<��a<ސa<�a<D�a<g�a<��a<�a<&�a<p�a<��a<��a<9�a<��a<ۓa<�a<{�a<Ĕa<&�a<z�a<ܕa<.�a<��a<��a<Q�a<җa<�a<��a<��a<^�a<řa<#�a<��a<�a<��a<�a<p�a<՜a<E�a<��a<)�a<��a<�a<��a<�a<f�a<Ԡa<C�a<��a<&�a<��a<�a<s�a<�a<F�a<��a<�a<v�a<�a<<�a<��a<�a<g�a<��a< �a<p�a<¨a<'�a<e�a<��a<	�a<Y�a<��a<ڪa<)�a<p�a<��a<߫a<1�a<S�a<��a<Ǭa<�a<,�a<U�a<��a<��a<حa<�a<�a<=�a<`�a<��a<��a<��a<Ϯa<�a<��a< �a<�a<'�a<5�a<H�a<V�a<O�a<X�a<l�a<\�a<q�a<k�a<T�a<d�a<U�a<R�a<+�a<<�a<+�a<%�a<�a<��a<��a<ʮa<Ʈa<��a<��a<t�a<Q�a<2�a<	�a<�a<��a<��a<x�a<R�a<2�a<�a<ݬa<��a<k�a<E�a< �a<٫a<��a<i�a<)�a<��a<��a<p�a<9�a<�a<��a<_�a<�a<ܨa<��a<5�a<اa<��a<I�a<��a<��a<V�a<�a<��a<B�a<ܤa<�a<"�a<ãa<U�a<��a<��a<*�a<ϡa<_�a< �a<��a<*�a<ǟa<R�a<�a<{�a<�a<��a<2�a<՜a<g�a<��a<��a<-�a<��a<O�a<��a<~�a<�a<��a<[�a<�a<��a<3�a<ٖa<m�a<�a<ϕa<`�a<�a<��a<c�a<�a<ɓa<��a<)�a<�a<��a<f�a<"�a<�a<��a<x�a<F�a<�a<ڐa<��a<{�a<b�a<6�a<�a<��a<�a<��a<��a<��a<��a<��a<��a<h�a<y�a<p�a<x�a<a�a<��a<��a<��a<��a<ɏa<�a<�  �  ��a<�a<D�a<V�a<��a<��a<Аa<'�a<<�a<��a<��a<�a<5�a<^�a<��a<ޒa<O�a<y�a<ޓa<"�a<w�a<��a<�a<��a<ӕa<9�a<��a<��a<X�a<��a<0�a<�a<�a<P�a<̙a<O�a<��a<�a<s�a<��a<^�a<˜a<I�a<��a<>�a<��a<�a<�a<�a<~�a<͠a<[�a<��a<2�a<��a<�a<s�a<أa<V�a<��a<,�a<p�a<��a<J�a<��a<�a<X�a<Чa<�a<r�a<��a<�a<u�a<��a<
�a<F�a<��a<�a<�a<g�a<��a<��a<�a<X�a<��a<Ĭa<�a<�a<e�a<u�a<��a<٭a<�a<,�a<2�a<s�a<m�a<��a<��a<׮a<�a<�a<�a<�a<I�a</�a<H�a<V�a<M�a<j�a<W�a<g�a<V�a<g�a<]�a<Q�a<P�a<I�a<`�a<6�a<#�a<�a<�a<�a<ծa<֮a<��a<��a<��a<r�a<U�a<$�a<*�a<�a<ԭa<��a<v�a<a�a< �a<�a<��a<��a<c�a<H�a<	�a<իa<��a<Y�a<8�a<�a<��a<t�a<3�a<�a<��a<q�a<�a<Шa<y�a<=�a<�a<��a<I�a<�a<��a<D�a<�a<��a<-�a<�a<s�a<.�a<��a<[�a<�a<��a<B�a<��a<l�a<��a<��a<)�a<��a<b�a<۞a<��a<�a<��a<A�a<ǜa<w�a<�a<��a<�a<��a<N�a<�a<��a<�a<��a<I�a<�a<��a< �a<іa<g�a<(�a<��a<e�a<�a<��a<q�a<�a<ٓa<q�a<B�a<�a<��a<s�a<�a<��a<��a<y�a<<�a<�a<ܐa<��a<��a<Y�a<Y�a<�a<��a<�a<��a<��a<��a<��a<v�a<~�a<q�a<f�a<k�a<o�a<��a<�a<��a<��a<��a<̏a<̏a<�  �  �a<�a<8�a<i�a<�a<��a<�a< �a<6�a<~�a<��a<�a<$�a<_�a<��a<�a<C�a<��a<ۓa<)�a<q�a<��a<&�a<~�a<֕a<?�a<��a<�a<_�a<��a<'�a<��a<�a<d�a<��a<#�a<��a<�a<��a<��a<`�a<՜a<N�a<��a<.�a<��a<	�a<��a<��a<]�a<Ѡa<Q�a<��a<0�a<��a<�a<u�a<ԣa<M�a<��a<!�a<x�a<ۥa<E�a<��a<�a<c�a<ŧa<�a<v�a<˨a<�a<o�a<��a<�a<M�a<��a<تa<(�a<g�a<��a<�a<�a<`�a<��a<Ŭa<��a<&�a<T�a<��a<��a<έa<��a<&�a<@�a<f�a<s�a<��a<��a<Ʈa<�a<�a<�a<�a< �a<<�a<O�a<F�a<`�a<[�a<Z�a<q�a<_�a<`�a<k�a<b�a<]�a<G�a<2�a<1�a<3�a< �a<�a<��a<�a<߮a<��a<��a<��a<f�a<V�a<6�a<�a<�a<ҭa<��a<��a<P�a< �a<�a<Ƭa<��a<t�a<F�a<�a<ϫa<��a<i�a<-�a<�a<��a<s�a<.�a<��a<��a<h�a<#�a<Ҩa<��a<0�a<اa<��a<J�a<��a<��a<E�a<�a<��a<7�a<�a<��a<�a<ţa<^�a<�a<��a<8�a<ѡa<i�a<��a<��a<+�a<��a<Y�a<�a<��a<�a<��a<;�a<Ҝa<a�a<��a<��a<$�a<a<X�a<�a<��a<%�a<��a<O�a<�a<��a<2�a<Жa<y�a<�a<��a<l�a<�a<��a<p�a<�a<ȓa<��a<,�a<�a<��a<m�a<%�a<�a<��a<��a<8�a<�a<�a<��a<��a<T�a<0�a<�a<�a<؏a<ҏa<��a<��a<��a<�a<x�a<�a<w�a<x�a<l�a<g�a<{�a<��a<��a<��a<Ǐa<؏a<�  �  �a<"�a<4�a<a�a<��a<��a<�a<�a<N�a<n�a<��a<�a<*�a<p�a<��a<��a<:�a<��a<̓a<'�a<��a<Ôa<3�a<o�a<�a<.�a<��a<��a<O�a<ϗa<�a<��a<�a<d�a<˙a<3�a<��a<�a<��a<�a<k�a<՜a<>�a<ɝa<�a<��a<�a<��a<��a<b�a<�a<=�a<��a<"�a<��a<�a<s�a<�a<B�a<��a<�a<��a<ߥa<B�a<��a<��a<q�a<��a<'�a<k�a<èa<'�a<_�a<��a<�a<a�a<��a<�a<-�a<_�a<��a<իa<3�a<Q�a<��a<̬a<�a<5�a<H�a<��a<��a<حa< �a<�a<B�a<]�a<��a<��a<��a<ծa<�a<��a< �a</�a<#�a<?�a<J�a<I�a<^�a<Q�a<n�a<Y�a<n�a<b�a<W�a<Z�a<T�a<V�a<B�a<?�a<,�a<�a<�a<��a<�a<Ǯa<Ʈa<��a<��a<m�a<O�a<:�a<�a<��a<­a<��a<{�a<W�a<1�a<��a<ܬa<��a<q�a<6�a<�a<߫a<��a<v�a<�a<��a<��a<y�a<5�a<�a<��a<U�a<�a<Ψa<��a<<�a<�a<��a<C�a<��a<��a<P�a<�a<��a<L�a<Ѥa<��a<�a<ʣa<^�a<��a<��a<$�a<ϡa<\�a<�a<��a<)�a<ϟa<O�a<�a<t�a<%�a<��a<8�a<ޜa<[�a<�a<��a<4�a<��a<P�a<��a<y�a<#�a<��a<d�a<�a<��a<7�a<ɖa<u�a<�a<Еa<^�a<�a<a<]�a<%�a<��a<��a<,�a<�a<��a<\�a<'�a<�a<��a<t�a<F�a<�a<ܐa<��a<{�a<r�a<3�a< �a<�a<ۏa<Ϗa<��a<��a<��a<��a<y�a<k�a<o�a<o�a<|�a<x�a<��a<��a<��a<��a<��a<�a<�  �  �a<�a<>�a<Y�a<��a<��a<֐a<�a<9�a<z�a<��a<�a<1�a<b�a<��a<�a<B�a<��a<��a<"�a<t�a<ؔa<�a<|�a<��a<,�a<��a<��a<K�a<��a<'�a<��a<��a<T�a<��a<<�a<��a<�a<�a<��a<a�a<͜a<?�a<��a<)�a<��a<�a<��a<��a<o�a<ՠa<N�a<¡a<,�a<��a<��a<h�a<ݣa<K�a<��a<�a<}�a<�a<L�a<��a<�a<c�a<��a<�a<n�a<��a<�a<r�a<��a<
�a<E�a<��a<ܪa<�a<l�a<��a<�a<�a<K�a<��a<ˬa<�a<+�a<V�a<~�a<��a<ӭa<��a<(�a<G�a<d�a<x�a<��a<��a<׮a<�a<�a<�a<�a<5�a<4�a<E�a<X�a<U�a<_�a<e�a<W�a<\�a<h�a<e�a<_�a<\�a<B�a<W�a<-�a<+�a<#�a<�a<�a<ݮa<Ůa<��a<��a<��a<w�a<O�a<)�a<�a<�a<έa<��a<��a<^�a<#�a<�a<ʬa<��a<y�a<K�a<	�a<ҫa<��a<`�a<+�a<��a<��a<|�a<3�a<�a<��a<h�a<!�a<٨a<}�a<1�a<�a<��a<K�a<�a<��a<F�a<�a<��a<<�a<ܤa<�a<(�a<£a<a�a<�a<��a<5�a<ҡa<e�a<��a<��a<�a<��a<X�a<�a<��a<�a<��a<C�a<ќa<k�a<��a<��a<&�a<��a<K�a<�a<��a<�a<��a<G�a<�a<��a<'�a<Ֆa<x�a<�a<��a<X�a<�a<��a<_�a<�a<ʓa<z�a<=�a<�a<��a<o�a<,�a<�a<��a<c�a<8�a<�a<ߐa<��a<��a<X�a<E�a<�a<��a<�a<Əa<��a<��a<��a<|�a<��a<x�a<t�a<w�a<h�a<��a<w�a<��a<��a<��a<͏a<ԏa<�  �  �a<
�a<?�a<a�a<�a<��a<ڐa<�a<+�a<�a<��a<�a<�a<g�a<ʒa<�a<9�a<|�a<ԓa<'�a<l�a<Дa<�a<��a<͕a<=�a<��a<�a<t�a<��a<1�a<��a<�a<c�a<ęa<7�a<��a<#�a<r�a< �a<W�a<ܜa<R�a<��a<<�a<��a<�a<��a<��a<g�a<ɠa<Z�a<��a<.�a<��a<�a<��a<ңa<N�a<��a<&�a<s�a<�a<H�a<��a<�a<Z�a<ѧa<�a<w�a<Өa<
�a<{�a<��a<�a<F�a<��a<ݪa<&�a<k�a<��a<��a<�a<q�a<��a<��a<�a<�a<g�a<u�a<��a<˭a<��a<#�a<4�a<a�a<y�a<��a<��a<îa<�a<�a<�a<�a<-�a<:�a<I�a<O�a<T�a<f�a<S�a<y�a<a�a<c�a<e�a<M�a<h�a<9�a<E�a<*�a<;�a<�a<�a<�a<�a<�a<��a<��a<��a<g�a<W�a<.�a<�a<حa<ӭa<��a<w�a<L�a<(�a<�a<ͬa<��a<g�a<?�a<�a<˫a<��a<[�a<;�a<�a<��a<s�a<'�a<�a<��a<r�a<�a<Шa<��a<5�a<�a<��a<Z�a<�a<��a<<�a<��a<��a</�a<�a<v�a<-�a<��a<_�a<��a<��a<B�a<��a<g�a<�a<��a<;�a<��a<Z�a<ߞa<��a<�a<��a<?�a<Ȝa<u�a<�a<��a<�a<Úa<`�a<ܙa<��a<�a<Ƙa<H�a<�a<��a<0�a<Ֆa<f�a<'�a<��a<~�a<�a<��a<t�a<
�a<ۓa<p�a<8�a<�a<��a<j�a<�a<�a<��a<��a<B�a<�a<ܐa<��a<��a<H�a<=�a<�a< �a<�a<Əa<��a<��a<��a<��a<z�a<y�a<c�a<��a<_�a<{�a<s�a<��a<��a<��a<͏a<ڏa<�  �  �a<�a<;�a<d�a<}�a<��a<�a<�a<V�a<w�a<��a<�a<(�a<k�a<��a<��a<;�a<��a<ʓa</�a<��a<Ɣa<-�a<x�a<ѕa<;�a<��a<�a<R�a<��a<�a<��a<�a<^�a<͙a<6�a<��a<�a<�a<�a<W�a<؜a<<�a<��a<+�a<��a<�a<��a<��a<c�a<�a<F�a<��a<2�a<��a< �a<k�a<�a<M�a<��a<�a<��a<ߥa<G�a<��a<�a<i�a<��a<�a<g�a<Ǩa<�a<f�a<��a<�a<Y�a<��a<�a<'�a<a�a<��a<۫a<�a<V�a<��a<Ƭa<��a<$�a<S�a<��a<��a<حa<�a<�a<F�a<a�a<��a<��a<��a<Ϯa<�a<�a<
�a<4�a<%�a<B�a<B�a<H�a<\�a<[�a<d�a<[�a<g�a<V�a<g�a<T�a<R�a<X�a<H�a<@�a<'�a<�a<�a<�a<�a<ʮa<��a<��a<��a<e�a<L�a<:�a<�a<�a<˭a<��a<��a<U�a<-�a<�a<֬a<��a<z�a<5�a<�a<�a<��a<p�a<'�a<�a<��a<u�a<*�a<�a<��a<X�a<�a<˨a<��a<=�a<�a<��a<G�a<�a<��a<=�a<��a<��a<=�a<ޤa<��a<�a<ţa<c�a<��a<��a<-�a<ǡa<l�a<�a<��a<"�a<ȟa<Y�a<�a<{�a<#�a<��a<=�a<לa<d�a< �a<��a<*�a<��a<U�a<��a<��a<�a<��a<\�a<�a<��a<1�a<ʖa<v�a<�a<��a<b�a<�a<��a<k�a<�a<Ɠa<��a<2�a<�a<��a<]�a<+�a<�a<��a<c�a<>�a<�a<�a<��a<��a<w�a<4�a<#�a<��a<ُa<͏a<��a<��a<��a<��a<m�a<{�a<i�a<m�a<~�a<}�a<��a<��a<��a<��a<��a<�a<�  �  ߏa<9�a<.�a<[�a<��a<��a<�a<�a<G�a<[�a<��a<�a<�a<��a<��a<�a<*�a<��a<ϓa<�a<u�a<Ôa<*�a<j�a<�a<'�a<��a<�a<D�a<ڗa<�a<��a<�a<X�a<Ιa<+�a<��a< �a<��a<�a<s�a<�a<?�a<ѝa<�a<��a<�a<��a<�a<X�a<ܠa<-�a<ҡa<�a<��a<�a<m�a<�a<7�a<ɤa< �a<��a<եa<A�a<��a<��a<{�a<��a<1�a<s�a<Ϩa</�a<e�a<ͩa<��a<W�a<��a<�a<#�a<]�a<��a<ګa<9�a<L�a<��a<άa<�a<@�a<C�a<��a<��a<ͭa<�a<�a<T�a<L�a<��a<��a<Ǯa<ɮa<߮a<�a<�a<%�a<�a<=�a<;�a<S�a<\�a<K�a<��a<K�a<��a<f�a<f�a<l�a<D�a<X�a<:�a<C�a<�a<(�a<�a<��a<
�a<��a<ܮa<��a<��a<y�a<B�a<6�a<�a<��a<��a<��a<~�a<J�a<B�a<�a<�a<��a<��a<:�a<��a<ӫa<��a<l�a<�a<�a<��a<s�a<K�a<کa<ȩa<\�a</�a<Ψa<��a<>�a<�a<��a<7�a<�a<��a<X�a< �a<��a<S�a<Ĥa<��a<�a<��a<\�a<�a<��a<�a<�a<U�a<
�a<��a<$�a<џa<C�a<�a<f�a<�a<��a<7�a<Ԝa<U�a<�a<x�a<>�a<��a<\�a<�a<�a<0�a<��a<Y�a<�a<��a<-�a<ǖa<��a<�a<וa<X�a<!�a<Ĕa<V�a<0�a<��a<��a<-�a<�a<��a<X�a<9�a<ԑa<a<]�a<R�a<	�a<ِa<Őa<j�a<h�a<-�a<�a<�a<�a<Ώa<��a<��a<x�a<��a<}�a<z�a<��a<_�a<~�a<o�a<��a<��a<��a<��a<Ïa<�a<�  �  ��a<�a<9�a<f�a<��a<��a<ܐa<�a<D�a<w�a<��a<ߑa<�a<u�a<��a<�a<*�a<��a<דa<-�a<��a<ܔa<�a<��a<Օa<6�a<��a<��a<U�a<��a<�a<��a<�a<g�a<ҙa<=�a<��a<�a<{�a<�a<Z�a<Μa<C�a<��a<+�a<��a<�a<��a<��a<z�a<�a<K�a<ša<�a<��a<�a<|�a<�a<9�a<��a<�a<��a<��a<P�a<��a<�a<i�a<��a<�a<m�a<��a<�a<b�a<��a<
�a<T�a<��a<�a<,�a<h�a<��a<ګa<�a<R�a<��a<Ĭa<��a<%�a<W�a<z�a<��a<�a<�a<!�a<C�a<P�a<��a<��a<®a<Ůa<Ԯa<�a<�a<#�a<8�a<;�a<I�a<I�a<`�a<[�a<f�a<_�a<`�a<`�a<V�a<W�a<X�a<L�a<E�a<<�a<2�a<�a<�a<��a<�a<Юa<��a<��a<��a<h�a<T�a</�a<�a<�a<ʭa<��a<r�a<I�a<7�a<�a<�a<��a<r�a<A�a<�a<߫a<��a<]�a</�a<�a<��a<r�a<6�a<�a<��a<[�a<�a<Шa<��a<C�a<�a<��a<K�a<�a<��a<@�a<�a<��a<>�a<ޤa<��a< �a<ģa<e�a<�a<��a<2�a<աa<Q�a<��a<��a<2�a<��a<E�a<�a<��a<#�a<��a<F�a<ќa<e�a< �a<��a<)�a<��a<M�a<�a<{�a<�a<��a<V�a<��a<��a<6�a<іa<k�a<�a<��a<^�a<�a<��a<i�a<�a<˓a<u�a<C�a<��a<��a<h�a<(�a<ؑa<��a<�a<M�a<�a<ΐa<��a<��a<f�a<H�a<�a< �a<ۏa<ҏa<��a<��a<��a<��a<w�a<j�a<l�a<s�a<r�a<{�a<��a<��a<��a<��a<��a<܏a<�  �  �a<�a<�a<7�a<C�a<��a<��a<�a<�a<Q�a<j�a<őa<�a</�a<��a<��a<+�a<X�a<��a<��a<<�a<��a<�a<p�a<��a< �a<r�a<Жa<Q�a<q�a<�a<s�a<Ԙa<-�a<��a<�a<b�a<��a<Y�a<��a<3�a<��a<8�a<��a<�a<q�a<�a<d�a<��a<E�a<��a<0�a<{�a<�a<q�a<�a<g�a<��a<:�a<w�a<��a<L�a<��a<�a<��a<�a<3�a<��a<��a<b�a<��a<�a<{�a<��a<��a<�a<v�a<��a<��a<T�a<��a<�a<�a<V�a<{�a<��a<�a<�a<O�a<Y�a<��a<��a<ԭa<�a<�a<Z�a<D�a<��a<��a<��a<ͮa<��a<�a<�a<�a<��a<=�a<!�a<7�a<L�a<4�a<c�a<0�a<F�a<c�a<:�a<=�a<
�a</�a<��a<�a<��a<�a<�a<��a<Ӯa<��a<��a<m�a<5�a<L�a<��a<�a<��a<��a<j�a<b�a<=�a<��a<�a<��a<��a<L�a<�a<�a<��a<|�a<9�a<(�a<��a<��a<Y�a<�a<�a<f�a<c�a<�a<��a<]�a<��a<̧a<_�a<4�a<Ѧa<��a<�a<ѥa<��a<�a<Ԥa<V�a<��a<��a<*�a<ڢa<a�a<�a<��a<U�a<Ԡa<x�a<�a<��a<D�a<��a<`�a<ݝa<��a<�a<��a<E�a<śa<��a<�a<��a<9�a<��a<��a<��a<��a<�a<ėa<U�a<��a<��a<T�a<�a<u�a<Y�a<�a<��a<Z�a<ғa<��a<J�a<�a<��a<w�a<,�a<�a<בa<h�a<x�a<�a<�a<��a<m�a<c�a<#�a<�a<Տa<�a<��a<��a<��a<h�a<��a<E�a<R�a<l�a<D�a<L�a<$�a<Z�a<3�a<h�a<t�a<��a<��a<��a<�  �  Ǐa<�a< �a<9�a<\�a<��a<��a<��a<�a<[�a<��a<��a<��a<4�a<x�a<��a<�a<]�a<��a<
�a<N�a<��a<��a<P�a<��a<�a<V�a<��a</�a<��a<�a<M�a<Ęa<;�a<��a<!�a<�a<��a<P�a<��a<+�a<��a<�a<��a<��a<��a<�a<a�a<؟a<O�a<��a<8�a<��a<�a<t�a<Ԣa<D�a<��a<*�a<��a<	�a<a�a<˥a<-�a<��a<�a<U�a<��a<�a<C�a<��a<�a<=�a<��a<�a<6�a<��a<̪a<�a<F�a<u�a<��a<��a<=�a<c�a<��a<׬a<�a<5�a<d�a<��a<��a<�a<�a<$�a<E�a<S�a<q�a<��a<��a<®a<�a<��a<��a<�a<�a<%�a<-�a<>�a</�a<9�a<;�a<K�a<1�a<,�a<4�a<A�a<1�a<=�a<�a<�a<��a<׮a<ʮa<ˮa<��a<��a<t�a<o�a<N�a<-�a<�a<�a<έa<��a<��a<[�a<6�a<��a<Ԭa<��a<��a<Q�a<)�a<��a<��a<��a<D�a<�a<֪a<��a<=�a<�a<ͩa<��a<5�a<�a<��a<k�a<!�a<ܧa<|�a<0�a<Ȧa<o�a<�a<եa<k�a<�a<��a<p�a<��a<��a<B�a<�a<u�a< �a<��a<A�a<֠a<`�a<��a<��a<4�a<˞a<l�a<�a<��a<�a<��a<>�a<�a<c�a<�a<��a<0�a<��a<P�a<�a<��a<1�a<ٗa<r�a<�a<��a<8�a<�a<��a<@�a<ؔa<{�a<>�a<��a<��a<U�a<�a<ƒa<��a<H�a<��a<a<w�a<A�a<�a<�a<��a<��a<l�a<7�a<#�a<�a<яa<��a<��a<z�a<m�a<]�a<`�a<=�a<4�a<>�a<Q�a<K�a<g�a<[�a<n�a<k�a<o�a<��a<��a<�  �  ��a<�a< �a</�a<f�a<p�a<Őa<Ґa<�a<9�a<��a<��a<��a<Z�a<t�a<�a<��a<X�a<��a<�a<D�a<��a<
�a<8�a<ŕa<��a<m�a<ۖa<�a<��a<�a<s�a<Θa</�a<��a<��a<}�a<�a<t�a<̛a<G�a<��a<�a<��a<�a<��a<۞a<\�a<֟a<1�a<��a<�a<��a<�a<��a<�a<S�a<Уa<�a<��a<�a<X�a<��a<#�a<��a<Цa<]�a<��a<�a<K�a<��a<	�a<H�a<��a<�a<1�a<m�a<��a< �a<G�a<��a<��a<�a<+�a<y�a<��a<Ƭa<"�a<�a<q�a<��a<��a<֭a<�a<#�a</�a<}�a<p�a<��a<��a<��a<�a<׮a<��a<��a<+�a<�a<.�a<7�a<+�a<f�a<�a<a�a<@�a<F�a<L�a<,�a<0�a<�a<�a<�a<�a<��a<Ԯa<�a<��a<��a<t�a<e�a<Y�a<�a<#�a<߭a<ɭa<��a<��a<N�a<-�a<&�a<Ьa<Ϭa<o�a<L�a<�a<�a<��a<r�a<V�a<�a<�a<��a<T�a<�a<��a<��a<<�a<�a<��a<_�a<�a<��a<z�a<!�a<�a<~�a<1�a<�a<e�a<>�a<��a<q�a<�a<��a<A�a<Ţa<o�a<��a<��a<,�a<�a<x�a<�a<��a<�a<Ӟa<G�a<�a<s�a<�a<��a<*�a<�a<O�a<�a<��a<5�a<ԙa<Z�a<�a<��a<,�a<��a<`�a<�a<��a<_�a<�a<��a<.�a<�a<��a<-�a<�a<��a<b�a< �a<��a<y�a</�a<��a<��a<��a<@�a<+�a<�a<��a<��a<G�a<1�a<��a<�a<Ïa<��a<��a<u�a<��a<A�a<v�a<M�a<O�a<V�a<<�a<K�a<;�a<V�a<[�a<��a<��a<��a<Տa<�  �  ďa<��a<�a<8�a<X�a<��a<a<ϐa<2�a<R�a<~�a<ӑa<��a<>�a<x�a<Ȓa<�a<r�a<��a<
�a<_�a<��a<�a<R�a<��a<�a<t�a<ǖa<*�a<��a<�a<c�a<��a<;�a<��a<�a<��a<�a<L�a<Лa<1�a<��a<�a<��a<�a<~�a<�a<k�a<ٟa<E�a<Ԡa<(�a<��a<�a<o�a<ۢa<F�a<��a<(�a<��a<��a<z�a<ͥa<+�a<��a<�a<F�a<��a<�a<B�a<��a<�a<L�a<��a<ߩa<;�a<��a<ʪa<�a<>�a<��a<��a<��a<5�a<h�a<��a<֬a<�a<5�a<u�a<��a<ĭa<�a<��a<4�a<@�a<^�a<r�a<��a<��a<Үa<֮a<�a<�a<��a<&�a<*�a<.�a<<�a<>�a<E�a<4�a<F�a<5�a<J�a<&�a<3�a<;�a<!�a<$�a<�a<�a<��a<ˮa<Ȯa<��a<��a<��a<m�a<J�a<1�a<!�a<ܭa<�a<��a<~�a<p�a</�a<	�a<Ԭa<��a<~�a<g�a<�a<��a<ƫa<p�a<Z�a<
�a<̪a<��a<Z�a<�a<ɩa<��a<;�a<��a<��a<j�a< �a<Чa<��a<�a<Ħa<��a<�a<ѥa<e�a<#�a<��a<c�a<�a<��a<C�a<ڢa<��a<�a<��a<G�a<Ҡa<g�a<��a<��a<2�a<Ҟa<Y�a<�a<��a<�a<��a<B�a<כa<e�a<�a<��a<.�a<��a<^�a<�a<��a<5�a<ӗa<p�a<�a<��a<H�a<�a<��a<8�a<ޔa<��a<=�a<�a<��a<f�a<�a<Ғa<��a<4�a<�a<��a<��a<B�a<�a<ސa<��a<��a<`�a<S�a<�a<��a<֏a<��a<��a<��a<y�a<V�a<[�a<A�a<S�a<0�a<C�a<U�a<L�a<c�a<f�a<^�a<��a<��a<��a<�  �  �a<؏a<�a<7�a<V�a<��a<��a<�a<�a<P�a<w�a<őa<��a<<�a<��a<a<�a<X�a<��a<��a<F�a<��a<�a<Y�a<��a<�a<k�a<��a<H�a<��a<�a<X�a<˘a<@�a<��a<�a<q�a<�a<L�a<�a<9�a<��a<)�a<��a<�a<m�a<�a<R�a<Οa<C�a<��a<+�a<��a<�a<v�a<�a<Y�a<��a<.�a<~�a<��a<U�a<��a<%�a<z�a<�a<5�a<��a<�a<P�a<��a<��a<a�a<��a<��a<)�a<x�a<��a<�a<O�a<|�a<٫a<�a<S�a<f�a<��a<�a<��a<@�a<Z�a<��a<��a<խa<��a<�a<F�a<Y�a<��a<��a<��a<ʮa<Ȯa<�a<��a<�a<�a< �a<-�a<3�a<H�a<)�a<X�a<E�a<C�a<L�a<-�a<P�a<�a<&�a<�a<%�a<�a<�a<�a<��a<ʮa<��a<��a<m�a<H�a<0�a<�a<��a<ĭa<��a<w�a<b�a<6�a<�a<�a<��a<��a<M�a<�a<�a<��a<��a<=�a<�a<Ūa<��a<Q�a<�a<�a<w�a<U�a<�a<��a<p�a<�a<ȧa<n�a<C�a<Ŧa<��a<#�a<ޥa<}�a<�a<Фa<R�a<�a<��a<8�a<آa<i�a<�a<��a<G�a<ؠa<v�a<�a<��a<8�a<��a<[�a<�a<�a<�a<��a<I�a<ƛa<�a<��a<��a<@�a<��a<s�a<�a<��a<#�a<Ɨa<[�a<	�a<��a<?�a<�a<��a<V�a<ܔa<��a<N�a<�a<��a<K�a<�a<��a<x�a<5�a<�a<Ña<}�a<W�a<�a<�a<��a<v�a<a�a<,�a<�a<�a<̏a<��a<��a<��a<]�a<z�a<Y�a<O�a<U�a<7�a<`�a<:�a<P�a<J�a<}�a<f�a<��a<��a<��a<�  �  ˏa<��a<�a<�a<k�a<��a<��a<�a<�a<N�a<��a<��a< �a<E�a<u�a<ђa<�a<V�a<��a<��a<H�a<��a<�a<Z�a<��a<�a<n�a<Җa<&�a<��a<�a<\�a<Әa<5�a<��a<�a<m�a<��a<Z�a<ʛa<8�a<��a<"�a<��a<�a<l�a<��a<^�a<ӟa<G�a<��a<-�a<��a<�a<{�a<ݢa<I�a<ģa<%�a<��a< �a<Z�a<��a<)�a<��a<��a<:�a<��a<�a<T�a<��a<��a<I�a<��a<�a<$�a<��a<Ūa<�a<N�a<��a<ȫa<��a<0�a<t�a<��a<Ƭa<	�a<@�a<\�a<��a<��a<ݭa<
�a<"�a<D�a<h�a<r�a<��a<��a<��a<�a<�a<�a<�a<�a<'�a<?�a< �a<;�a<L�a<B�a<;�a<>�a<>�a<B�a<7�a<�a<<�a<�a<�a<�a<�a<ݮa<��a<��a<��a<��a<P�a<]�a<5�a<�a<��a<��a<��a<��a<T�a<7�a<�a<Ѭa<��a<��a<J�a<,�a<�a<��a<��a<<�a<�a<תa<y�a<U�a<�a<ũa<~�a<I�a<��a<��a<d�a<�a<٧a<j�a<1�a<Ҧa<}�a<"�a<ȥa<v�a<'�a<��a<Q�a<�a<��a<=�a<ܢa<m�a<�a<��a<=�a<ݠa<i�a<��a<��a</�a<͞a<c�a<�a<��a<�a<��a<N�a<̛a<d�a<
�a<��a<%�a<��a<[�a<�a<��a<�a<֗a<k�a<�a<��a<E�a<�a<��a<3�a<�a<��a<-�a<�a<��a<N�a<�a<��a<��a<G�a<��a<��a<��a<B�a<�a<�a<��a<��a<^�a<'�a<�a<�a<ӏa<ŏa<��a<��a<��a<d�a<P�a<J�a<G�a<L�a<G�a<3�a<f�a<D�a<c�a<|�a<��a<��a<��a<�  �  ʏa<�a<�a<5�a<[�a<��a<��a<��a<)�a<H�a<��a<��a<��a<I�a<��a<͒a<
�a<]�a<��a<��a<\�a<��a<�a<L�a<��a<�a<l�a<ʖa<.�a<��a<�a<a�a<Øa<4�a<��a<�a<��a<�a<^�a<��a<L�a<��a<�a<��a<��a<��a<�a<f�a<Пa<C�a<Πa<�a<��a<��a<{�a<�a<V�a<��a<�a<��a<�a<t�a<ǥa<$�a<��a<�a<Q�a<��a< �a<M�a<��a<�a<<�a<��a<ܩa<6�a<�a<ƪa<�a<?�a<��a<��a<�a<6�a<n�a<��a<Ӭa<�a<.�a<k�a<��a<��a<�a<�a<#�a<7�a<d�a<��a<��a<��a<��a<خa<�a<�a<�a<�a<%�a<-�a<?�a<7�a<F�a<:�a<T�a<E�a<7�a<:�a</�a<2�a<&�a<!�a<�a<��a<�a<ٮa<ڮa<��a<��a<�a<k�a<M�a<.�a<�a<�a<�a<��a<��a<Z�a<0�a<�a<�a<��a<z�a<Q�a<�a<�a<īa<v�a<M�a<�a<٪a<��a<R�a<�a<ͩa<��a<8�a<��a<��a<d�a< �a<Χa<}�a<�a<֦a<p�a<6�a<٥a<l�a<#�a<��a<k�a<��a<��a<:�a<آa<��a<�a<��a<9�a<ݠa<t�a<�a<��a<(�a<ʞa<L�a<�a<��a<�a<��a<:�a<�a<c�a<�a<��a<1�a<ؙa<N�a<��a<��a<0�a<͗a<m�a<	�a<��a<K�a<��a<��a<9�a<�a<��a<:�a<��a<��a<\�a<�a<ϒa<��a<.�a<��a<��a<��a<Q�a<�a<��a<��a<��a<T�a<L�a<�a<�a<Џa<��a<��a<��a<z�a<\�a<i�a<Q�a<@�a<D�a<?�a<M�a<Q�a<`�a<_�a<p�a<�a<��a<Əa<�  �  ۏa<�a<�a<B�a<A�a<��a<��a<ސa<�a<O�a<��a<ɑa<��a</�a<��a<��a<�a<c�a<��a<��a<E�a<��a<�a<P�a<��a<�a<k�a<Ŗa<9�a<��a<��a<p�a<Řa<6�a<��a<�a<��a<�a<^�a<כa<@�a<��a<&�a<��a<�a<y�a<ߞa<f�a<ןa<<�a<��a<)�a<��a<�a<p�a<�a<]�a<��a<2�a<��a<��a<X�a<��a<*�a<��a<ަa<<�a<��a<��a<U�a<��a<��a<S�a<��a<�a<:�a<q�a<��a<�a<C�a<��a<ȫa<��a<>�a<o�a<��a<�a<��a<3�a<o�a<��a<��a<ԭa<��a<"�a<J�a<N�a<��a<��a<��a<ͮa<Ӯa<�a<�a<�a<!�a<(�a<�a<B�a<C�a<6�a<K�a<;�a<D�a<M�a<3�a<8�a<6�a<�a<!�a<�a<��a<��a<ݮa<��a<��a<��a<��a<x�a<3�a<2�a<�a<�a<ía<��a<��a<f�a<4�a<��a<��a<��a<��a<W�a<�a<�a<��a<}�a<P�a<�a<��a<��a<Q�a<	�a<ةa<{�a<D�a<	�a<��a<f�a<�a<��a<��a<)�a<֦a<��a<*�a<ͥa<z�a<�a<Ȥa<^�a<�a<��a<A�a<Ѣa<m�a<�a<��a<I�a<Ҡa<v�a<�a<��a<<�a<a<Z�a<�a<|�a<�a<��a<8�a<Λa<x�a<��a<��a<*�a<Ùa<e�a<��a<��a<4�a<��a<a�a<	�a<��a<U�a<�a<��a<@�a<�a<��a<L�a<ݓa<��a<`�a<	�a<��a<x�a<:�a<��a<Ǒa<r�a<]�a<�a<�a<��a<��a<b�a<*�a<
�a<��a<ӏa<��a<��a<��a<i�a<m�a<P�a<Q�a<V�a<=�a<H�a<Q�a<?�a<_�a<g�a<j�a<��a<��a<��a<�  �  ҏa<�a<�a<-�a<a�a<��a<��a<��a<	�a<V�a<��a<��a<�a<2�a<��a<��a<-�a<O�a<��a<��a<T�a<��a<�a<a�a<��a<�a<c�a<Ėa<2�a<��a<��a<O�a<јa<6�a<��a<�a<x�a<�a<N�a<Ǜa<6�a<��a<%�a<��a<�a<m�a< �a<[�a<˟a<]�a<��a<>�a<��a<�a<u�a<ڢa<M�a<��a<<�a<��a<�a<W�a<ץa<#�a<~�a<��a<5�a<��a<�a<Q�a<��a<�a<H�a<��a<�a<0�a<��a<ƪa<�a<M�a<t�a<ɫa<��a<9�a<j�a<��a<ڬa<��a<H�a<R�a<��a<��a<حa<�a<�a<^�a<T�a<{�a<��a<��a<��a<Үa<��a<�a<$�a<	�a<(�a<5�a<.�a<A�a<9�a<G�a<<�a<B�a<5�a<;�a<7�a<(�a<.�a<�a<�a<�a<�a<ޮa<��a<��a<��a<��a<b�a<S�a<6�a<��a<�a<��a<��a<��a<R�a<L�a<��a<�a<��a<��a<C�a<-�a<�a<��a<��a<0�a<�a<Ǫa<��a<I�a<�a<Щa<��a<H�a<�a<��a<f�a<�a<ԧa<u�a<,�a<Ʀa<y�a< �a<ǥa<y�a<�a<Ȥa<R�a<�a<��a<5�a<�a<j�a<&�a<��a<M�a<ؠa<e�a<�a<��a<F�a<��a<r�a<�a<��a<�a<��a<V�a<Ǜa<u�a<��a<��a<&�a<��a<Z�a<�a<��a<*�a<їa<l�a<�a<��a<7�a<�a<��a<<�a<��a<��a<A�a<�a<��a<C�a<�a<ϒa<{�a<P�a<�a<ۑa<x�a<K�a<
�a<�a<��a<�a<n�a<#�a<)�a<ߏa<ԏa<��a<��a<��a<m�a<h�a<P�a<O�a<>�a<E�a<G�a<B�a<X�a<R�a<e�a<w�a<x�a<��a<��a<�  �  ��a<��a<�a<0�a<_�a<��a<��a<ڐa<�a<?�a<��a<��a<�a<I�a<��a<֒a<�a<H�a<��a<�a<P�a<��a<�a<U�a<��a<�a<q�a<זa<#�a<��a<��a<`�a<՘a</�a<��a<�a<y�a<�a<m�a<śa<T�a<��a<�a<��a<�a<x�a<�a<h�a<ɟa<A�a<��a<$�a<��a< �a<��a<�a<\�a<ƣa< �a<��a<��a<V�a<åa<�a<��a<�a<E�a<��a<�a<S�a<��a<�a<H�a<��a<�a<+�a<p�a<��a<��a<N�a<��a<ūa<�a<6�a<x�a<��a<ڬa<�a<4�a<l�a<}�a<��a<ϭa<�a<�a<:�a<i�a<��a<��a<��a<��a<ݮa<�a<��a<�a<�a<+�a<0�a<3�a<;�a<U�a<1�a<W�a<O�a<5�a<R�a</�a<-�a<�a<�a<�a<�a<�a<�a<�a<��a<��a<��a<e�a<Q�a</�a<�a<�a<ͭa<��a<��a<K�a<8�a<�a<ެa<��a<}�a<<�a<'�a<ݫa<��a<n�a<L�a<�a<ժa<��a<X�a<�a<��a<��a<E�a<��a<��a<_�a<�a<��a<v�a<&�a<�a<x�a<?�a<ݥa<p�a<*�a<��a<]�a<��a<��a<4�a<֢a<n�a<�a<��a<9�a<�a<z�a<�a<��a<*�a<��a<Z�a<�a<��a<�a<��a<;�a<֛a<k�a<�a<��a<:�a<��a<Z�a<�a<��a<%�a<��a<`�a<��a<��a<M�a<�a<��a<8�a<�a<��a<A�a<��a<��a<]�a<��a<Œa<r�a<A�a<�a<��a<��a<O�a<�a<�a<��a<��a<T�a<3�a<�a<�a<׏a<��a<��a<��a<��a<S�a<k�a<[�a<>�a<\�a<?�a<G�a<C�a<W�a<]�a<��a<}�a<��a<͏a<�  �  ��a< �a<��a<C�a<S�a<z�a<Аa<��a<8�a<D�a<��a<̑a<��a<<�a<q�a<̒a<
�a<p�a<��a<��a<h�a<��a<�a<?�a<��a<�a<a�a<ۖa<�a<��a<�a<p�a<��a<9�a<��a<�a<��a<ؚa<`�a<��a<9�a<��a<�a<��a<�a<��a<ٞa<q�a<ڟa<<�a<Ѡa< �a<��a<�a<s�a<ܢa<F�a<��a<"�a<��a<�a<q�a<ƥa<%�a<��a<ͦa<_�a<��a<��a<L�a<��a<�a<8�a<��a<өa<H�a<x�a<˪a<�a<3�a<��a<��a<��a<$�a<w�a<��a<Ȭa<�a<�a<��a<w�a<ɭa<�a<�a<9�a<;�a<b�a<k�a<��a<��a<ˮa<�a<�a<�a<�a<-�a<"�a< �a<K�a<"�a<R�a<5�a<;�a<8�a<>�a<4�a<$�a<M�a<�a<6�a<�a<�a<�a<ˮa<��a<��a<��a<k�a<x�a<E�a<$�a<.�a<̭a<�a<��a<��a<j�a<,�a<�a<ͬa<��a<z�a<e�a<#�a<�a<Ыa<]�a<k�a<��a<Ԫa<��a<G�a<�a<��a<��a<-�a<	�a<��a<i�a<)�a<��a<��a<�a<٦a<p�a<$�a<¥a<m�a<'�a<��a<{�a<�a<��a<D�a<Ѣa<��a<�a<��a<?�a<ՠa<g�a<��a<��a<,�a<�a<U�a<�a<��a<�a<Ɯa<'�a<�a<S�a<�a<��a<�a<��a<J�a<�a<}�a<C�a<Ǘa<q�a<�a<��a<X�a<ڕa<��a<'�a<�a<��a</�a<��a<��a<y�a<��a<גa<��a<=�a<�a<��a<��a<;�a<�a<ܐa<��a<��a<V�a<V�a<�a<�a<Ώa<��a<��a<l�a<��a<W�a<P�a<E�a<F�a<>�a<4�a<g�a<?�a<u�a<Y�a<f�a<��a<��a<��a<�  �  ߏa<�a<�a<5�a<_�a<v�a<��a<ܐa<�a<<�a<m�a<��a<�a<C�a<��a<̒a<�a<U�a<��a<�a<U�a<��a<�a<F�a<��a<	�a<l�a<͖a<>�a<��a<
�a<n�a<ʘa<6�a<��a<�a<r�a<�a<`�a<ٛa<G�a<��a<.�a<��a<�a<��a<�a<L�a<şa<H�a<��a<�a<��a<	�a<y�a<�a<`�a<£a<+�a<��a<�a<Q�a<ƥa<�a<w�a<�a<T�a<��a<��a<Z�a<��a<��a<\�a<��a<�a<-�a<n�a<��a<�a<G�a<��a<֫a< �a<E�a<t�a<��a<Ӭa<�a<+�a<Z�a<��a<��a<ȭa<�a<�a<K�a<c�a<��a<��a<��a<��a<®a<ޮa<��a<	�a<�a<�a</�a<<�a<8�a<=�a<R�a<C�a<R�a<J�a<;�a<6�a<�a<�a<�a<�a<��a<��a<�a<Ǯa<îa<��a<�a<k�a<Q�a<!�a<�a<�a<ϭa<��a<m�a<U�a<>�a<�a<��a<��a<��a<I�a<
�a<ثa<��a<u�a<>�a<��a<תa<��a<R�a<�a<ݩa<��a<R�a<�a<��a<f�a<	�a<��a<o�a<+�a<ئa<��a<2�a<ӥa<��a<�a<��a<j�a<��a<��a</�a<ݢa<l�a<�a<��a<B�a<۠a<|�a<�a<��a<5�a<��a<N�a<�a<��a<
�a<��a<;�a<�a<h�a<�a<��a<4�a<əa<n�a<��a<��a<'�a<��a<V�a<�a<��a<Q�a< �a<��a<G�a<�a<��a<:�a<��a<��a<K�a< �a<ʒa<k�a<+�a<�a<ȑa<��a<a�a<�a<�a<��a<o�a<N�a<0�a<�a<�a<��a<��a<��a<��a<q�a<t�a<W�a<_�a<R�a<E�a<F�a<9�a<C�a<L�a<e�a<s�a<��a<��a<��a<�  �  Џa<؏a<+�a<�a<b�a<��a<��a<�a<��a<a�a<��a<đa< �a<�a<��a<��a<�a<Z�a<ϓa<��a<@�a<��a<�a<e�a<��a<�a<�a<��a<4�a<��a<�a<H�a<טa<8�a<��a<8�a<b�a<�a<L�a<��a<2�a<��a<�a<��a<�a<a�a<
�a<f�a<ߟa<^�a<��a<R�a<��a<�a<g�a<آa<J�a<��a<6�a<��a<(�a<J�a<ԥa<6�a<��a<�a<1�a<��a<��a<H�a<��a<�a<M�a<��a<��a<!�a<��a<Īa<�a<Y�a<j�a<Ыa<�a<;�a<\�a<��a<Ҭa<�a<K�a<\�a<��a<��a<ӭa<*�a< �a<M�a<C�a<��a<w�a<��a<ͮa<�a<
�a<ܮa</�a<�a<+�a<>�a<�a<Y�a<0�a<B�a<0�a<E�a<%�a<:�a<K�a<�a<S�a<�a<�a< �a<Үa<�a<��a<��a<��a<��a<N�a<U�a<9�a<�a<�a<��a<��a<��a<a�a<6�a<�a<�a<��a<��a<O�a<C�a<�a<��a<��a<;�a<�a<Ϫa<��a<e�a<��a<ҩa<v�a<K�a<�a<��a<h�a<�a<�a<_�a<>�a<Ŧa<s�a<�a<ƥa<q�a<�a<Ҥa<F�a<�a<��a<J�a<�a<Y�a<:�a<��a<P�a<ɠa<c�a<��a<��a<@�a<ʞa<��a<۝a<��a<(�a<��a<]�a<a<t�a<��a<��a<)�a<��a<_�a<ޘa<��a<�a<�a<j�a<�a<��a<-�a<��a<��a<>�a<єa<��a<:�a<�a<��a<N�a<#�a<��a<v�a<f�a<��a<ʑa<g�a<Q�a<��a<ݐa<��a<��a<z�a<�a<3�a<�a<׏a<ŏa<�a<��a<d�a<d�a<D�a<Q�a<.�a<D�a<[�a<-�a<}�a<C�a<o�a<v�a<k�a<��a<��a<�  �  ߏa<�a<�a<5�a<_�a<v�a<��a<ܐa<�a<<�a<m�a<��a<�a<C�a<��a<̒a<�a<U�a<��a<�a<U�a<��a<�a<F�a<��a<	�a<l�a<͖a<>�a<��a<
�a<n�a<ʘa<6�a<��a<�a<r�a<�a<`�a<ٛa<G�a<��a<.�a<��a<�a<��a<�a<L�a<şa<H�a<��a<�a<��a<	�a<y�a<�a<`�a<£a<+�a<��a<�a<Q�a<ƥa<�a<w�a<�a<T�a<��a<��a<Z�a<��a<��a<\�a<��a<�a<-�a<n�a<��a<�a<G�a<��a<֫a< �a<E�a<t�a<��a<Ӭa<�a<+�a<Z�a<��a<��a<ȭa<�a<�a<K�a<c�a<��a<��a<��a<��a<®a<ޮa<��a<	�a<�a<�a</�a<<�a<8�a<=�a<R�a<C�a<R�a<J�a<;�a<6�a<�a<�a<�a<�a<��a<��a<�a<Ǯa<îa<��a<�a<k�a<Q�a<!�a<�a<�a<ϭa<��a<m�a<U�a<>�a<�a<��a<��a<��a<I�a<
�a<ثa<��a<u�a<>�a<��a<תa<��a<R�a<�a<ݩa<��a<R�a<�a<��a<f�a<	�a<��a<o�a<+�a<ئa<��a<2�a<ӥa<��a<�a<��a<j�a<��a<��a</�a<ݢa<l�a<�a<��a<B�a<۠a<|�a<�a<��a<5�a<��a<N�a<�a<��a<
�a<��a<;�a<�a<h�a<�a<��a<4�a<əa<n�a<��a<��a<'�a<��a<V�a<�a<��a<Q�a< �a<��a<G�a<�a<��a<:�a<��a<��a<K�a< �a<ʒa<k�a<+�a<�a<ȑa<��a<a�a<�a<�a<��a<o�a<N�a<0�a<�a<�a<��a<��a<��a<��a<q�a<t�a<W�a<_�a<R�a<E�a<F�a<9�a<C�a<L�a<e�a<s�a<��a<��a<��a<�  �  ��a< �a<��a<C�a<S�a<z�a<Аa<��a<8�a<D�a<��a<̑a<��a<<�a<q�a<̒a<
�a<p�a<��a<��a<h�a<��a<�a<?�a<��a<�a<a�a<ۖa<�a<��a<�a<p�a<��a<9�a<��a<�a<��a<ؚa<`�a<��a<9�a<��a<�a<��a<�a<��a<ٞa<q�a<ڟa<<�a<Ѡa< �a<��a<�a<s�a<ܢa<F�a<��a<"�a<��a<�a<q�a<ƥa<%�a<��a<ͦa<_�a<��a<��a<L�a<��a<�a<8�a<��a<өa<H�a<x�a<˪a<�a<3�a<��a<��a<��a<$�a<w�a<��a<Ȭa<�a<�a<��a<w�a<ɭa<�a<�a<9�a<;�a<b�a<k�a<��a<��a<ˮa<�a<�a<�a<�a<-�a<"�a< �a<K�a<"�a<R�a<5�a<;�a<8�a<>�a<4�a<$�a<M�a<�a<6�a<�a<�a<�a<ˮa<��a<��a<��a<k�a<x�a<E�a<$�a<.�a<̭a<�a<��a<��a<j�a<,�a<�a<ͬa<��a<z�a<e�a<#�a<�a<Ыa<]�a<k�a<��a<Ԫa<��a<G�a<�a<��a<��a<-�a<	�a<��a<i�a<)�a<��a<��a<�a<٦a<p�a<$�a<¥a<m�a<'�a<��a<{�a<�a<��a<D�a<Ѣa<��a<�a<��a<?�a<ՠa<g�a<��a<��a<,�a<�a<U�a<�a<��a<�a<Ɯa<'�a<�a<S�a<�a<��a<�a<��a<J�a<�a<}�a<C�a<Ǘa<q�a<�a<��a<X�a<ڕa<��a<'�a<�a<��a</�a<��a<��a<y�a<��a<גa<��a<=�a<�a<��a<��a<;�a<�a<ܐa<��a<��a<V�a<V�a<�a<�a<Ώa<��a<��a<l�a<��a<W�a<P�a<E�a<F�a<>�a<4�a<g�a<?�a<u�a<Y�a<f�a<��a<��a<��a<�  �  ��a<��a<�a<0�a<_�a<��a<��a<ڐa<�a<?�a<��a<��a<�a<I�a<��a<֒a<�a<H�a<��a<�a<P�a<��a<�a<U�a<��a<�a<q�a<זa<#�a<��a<��a<`�a<՘a</�a<��a<�a<y�a<�a<m�a<śa<T�a<��a<�a<��a<�a<x�a<�a<h�a<ɟa<A�a<��a<$�a<��a< �a<��a<�a<\�a<ƣa< �a<��a<��a<V�a<åa<�a<��a<�a<E�a<��a<�a<S�a<��a<�a<H�a<��a<�a<+�a<p�a<��a<��a<N�a<��a<ūa<�a<6�a<x�a<��a<ڬa<�a<4�a<l�a<}�a<��a<ϭa<�a<�a<:�a<i�a<��a<��a<��a<��a<ݮa<�a<��a<�a<�a<+�a<0�a<3�a<;�a<U�a<1�a<W�a<O�a<5�a<R�a</�a<-�a<�a<�a<�a<�a<�a<�a<�a<��a<��a<��a<e�a<Q�a</�a<�a<�a<ͭa<��a<��a<K�a<8�a<�a<ެa<��a<}�a<<�a<'�a<ݫa<��a<n�a<L�a<�a<ժa<��a<X�a<�a<��a<��a<E�a<��a<��a<_�a<�a<��a<v�a<&�a<�a<x�a<?�a<ݥa<p�a<*�a<��a<]�a<��a<��a<4�a<֢a<n�a<�a<��a<9�a<�a<z�a<�a<��a<*�a<��a<Z�a<�a<��a<�a<��a<;�a<֛a<k�a<�a<��a<:�a<��a<Z�a<�a<��a<%�a<��a<`�a<��a<��a<M�a<�a<��a<8�a<�a<��a<A�a<��a<��a<]�a<��a<Œa<r�a<A�a<�a<��a<��a<O�a<�a<�a<��a<��a<T�a<3�a<�a<�a<׏a<��a<��a<��a<��a<S�a<k�a<[�a<>�a<\�a<?�a<G�a<C�a<W�a<]�a<��a<}�a<��a<͏a<�  �  ҏa<�a<�a<-�a<a�a<��a<��a<��a<	�a<V�a<��a<��a<�a<2�a<��a<��a<-�a<O�a<��a<��a<T�a<��a<�a<a�a<��a<�a<c�a<Ėa<2�a<��a<��a<O�a<јa<6�a<��a<�a<x�a<�a<N�a<Ǜa<6�a<��a<%�a<��a<�a<m�a< �a<[�a<˟a<]�a<��a<>�a<��a<�a<u�a<ڢa<M�a<��a<<�a<��a<�a<W�a<ץa<#�a<~�a<��a<5�a<��a<�a<Q�a<��a<�a<H�a<��a<�a<0�a<��a<ƪa<�a<M�a<t�a<ɫa<��a<9�a<j�a<��a<ڬa<��a<H�a<R�a<��a<��a<حa<�a<�a<^�a<T�a<{�a<��a<��a<��a<Үa<��a<�a<$�a<	�a<(�a<5�a<.�a<A�a<9�a<G�a<<�a<B�a<5�a<;�a<7�a<(�a<.�a<�a<�a<�a<�a<ޮa<��a<��a<��a<��a<b�a<S�a<6�a<��a<�a<��a<��a<��a<R�a<L�a<��a<�a<��a<��a<C�a<-�a<�a<��a<��a<0�a<�a<Ǫa<��a<I�a<�a<Щa<��a<H�a<�a<��a<f�a<�a<ԧa<u�a<,�a<Ʀa<y�a< �a<ǥa<y�a<�a<Ȥa<R�a<�a<��a<5�a<�a<j�a<&�a<��a<M�a<ؠa<e�a<�a<��a<F�a<��a<r�a<�a<��a<�a<��a<V�a<Ǜa<u�a<��a<��a<&�a<��a<Z�a<�a<��a<*�a<їa<l�a<�a<��a<7�a<�a<��a<<�a<��a<��a<A�a<�a<��a<C�a<�a<ϒa<{�a<P�a<�a<ۑa<x�a<K�a<
�a<�a<��a<�a<n�a<#�a<)�a<ߏa<ԏa<��a<��a<��a<m�a<h�a<P�a<O�a<>�a<E�a<G�a<B�a<X�a<R�a<e�a<w�a<x�a<��a<��a<�  �  ۏa<�a<�a<B�a<A�a<��a<��a<ސa<�a<O�a<��a<ɑa<��a</�a<��a<��a<�a<c�a<��a<��a<E�a<��a<�a<P�a<��a<�a<k�a<Ŗa<9�a<��a<��a<p�a<Řa<6�a<��a<�a<��a<�a<^�a<כa<@�a<��a<&�a<��a<�a<y�a<ߞa<f�a<ןa<<�a<��a<)�a<��a<�a<p�a<�a<]�a<��a<2�a<��a<��a<X�a<��a<*�a<��a<ަa<<�a<��a<��a<U�a<��a<��a<S�a<��a<�a<:�a<q�a<��a<�a<C�a<��a<ȫa<��a<>�a<o�a<��a<�a<��a<3�a<o�a<��a<��a<ԭa<��a<"�a<J�a<N�a<��a<��a<��a<ͮa<Ӯa<�a<�a<�a<!�a<(�a<�a<B�a<C�a<6�a<K�a<;�a<D�a<M�a<3�a<8�a<6�a<�a<!�a<�a<��a<��a<ݮa<��a<��a<��a<��a<x�a<3�a<2�a<�a<�a<ía<��a<��a<f�a<4�a<��a<��a<��a<��a<W�a<�a<�a<��a<}�a<P�a<�a<��a<��a<Q�a<	�a<ةa<{�a<D�a<	�a<��a<f�a<�a<��a<��a<)�a<֦a<��a<*�a<ͥa<z�a<�a<Ȥa<^�a<�a<��a<A�a<Ѣa<m�a<�a<��a<I�a<Ҡa<v�a<�a<��a<<�a<a<Z�a<�a<|�a<�a<��a<8�a<Λa<x�a<��a<��a<*�a<Ùa<e�a<��a<��a<4�a<��a<a�a<	�a<��a<U�a<�a<��a<@�a<�a<��a<L�a<ݓa<��a<`�a<	�a<��a<x�a<:�a<��a<Ǒa<r�a<]�a<�a<�a<��a<��a<b�a<*�a<
�a<��a<ӏa<��a<��a<��a<i�a<m�a<P�a<Q�a<V�a<=�a<H�a<Q�a<?�a<_�a<g�a<j�a<��a<��a<��a<�  �  ʏa<�a<�a<5�a<[�a<��a<��a<��a<)�a<H�a<��a<��a<��a<I�a<��a<͒a<
�a<]�a<��a<��a<\�a<��a<�a<L�a<��a<�a<l�a<ʖa<.�a<��a<�a<a�a<Øa<4�a<��a<�a<��a<�a<^�a<��a<L�a<��a<�a<��a<��a<��a<�a<f�a<Пa<C�a<Πa<�a<��a<��a<{�a<�a<V�a<��a<�a<��a<�a<t�a<ǥa<$�a<��a<�a<Q�a<��a< �a<M�a<��a<�a<<�a<��a<ܩa<6�a<�a<ƪa<�a<?�a<��a<��a<�a<6�a<n�a<��a<Ӭa<�a<.�a<k�a<��a<��a<�a<�a<#�a<7�a<d�a<��a<��a<��a<��a<خa<�a<�a<�a<�a<%�a<-�a<?�a<7�a<F�a<:�a<T�a<E�a<7�a<:�a</�a<2�a<&�a<!�a<�a<��a<�a<ٮa<ڮa<��a<��a<�a<k�a<M�a<.�a<�a<�a<�a<��a<��a<Z�a<0�a<�a<�a<��a<z�a<Q�a<�a<�a<īa<v�a<M�a<�a<٪a<��a<R�a<�a<ͩa<��a<8�a<��a<��a<d�a< �a<Χa<}�a<�a<֦a<p�a<6�a<٥a<l�a<#�a<��a<k�a<��a<��a<:�a<آa<��a<�a<��a<9�a<ݠa<t�a<�a<��a<(�a<ʞa<L�a<�a<��a<�a<��a<:�a<�a<c�a<�a<��a<1�a<ؙa<N�a<��a<��a<0�a<͗a<m�a<	�a<��a<K�a<��a<��a<9�a<�a<��a<:�a<��a<��a<\�a<�a<ϒa<��a<.�a<��a<��a<��a<Q�a<�a<��a<��a<��a<T�a<L�a<�a<�a<Џa<��a<��a<��a<z�a<\�a<i�a<Q�a<@�a<D�a<?�a<M�a<Q�a<`�a<_�a<p�a<�a<��a<Əa<�  �  ˏa<��a<�a<�a<k�a<��a<��a<�a<�a<N�a<��a<��a< �a<E�a<u�a<ђa<�a<V�a<��a<��a<H�a<��a<�a<Z�a<��a<�a<n�a<Җa<&�a<��a<�a<\�a<Әa<5�a<��a<�a<m�a<��a<Z�a<ʛa<8�a<��a<"�a<��a<�a<l�a<��a<^�a<ӟa<G�a<��a<-�a<��a<�a<{�a<ݢa<I�a<ģa<%�a<��a< �a<Z�a<��a<)�a<��a<��a<:�a<��a<�a<T�a<��a<��a<I�a<��a<�a<$�a<��a<Ūa<�a<N�a<��a<ȫa<��a<0�a<t�a<��a<Ƭa<	�a<@�a<\�a<��a<��a<ݭa<
�a<"�a<D�a<h�a<r�a<��a<��a<��a<�a<�a<�a<�a<�a<'�a<?�a< �a<;�a<L�a<B�a<;�a<>�a<>�a<B�a<7�a<�a<<�a<�a<�a<�a<�a<ݮa<��a<��a<��a<��a<P�a<]�a<5�a<�a<��a<��a<��a<��a<T�a<7�a<�a<Ѭa<��a<��a<J�a<,�a<�a<��a<��a<<�a<�a<תa<y�a<U�a<�a<ũa<~�a<I�a<��a<��a<d�a<�a<٧a<j�a<1�a<Ҧa<}�a<"�a<ȥa<v�a<'�a<��a<Q�a<�a<��a<=�a<ܢa<m�a<�a<��a<=�a<ݠa<i�a<��a<��a</�a<͞a<c�a<�a<��a<�a<��a<N�a<̛a<d�a<
�a<��a<%�a<��a<[�a<�a<��a<�a<֗a<k�a<�a<��a<E�a<�a<��a<3�a<�a<��a<-�a<�a<��a<N�a<�a<��a<��a<G�a<��a<��a<��a<B�a<�a<�a<��a<��a<^�a<'�a<�a<�a<ӏa<ŏa<��a<��a<��a<d�a<P�a<J�a<G�a<L�a<G�a<3�a<f�a<D�a<c�a<|�a<��a<��a<��a<�  �  �a<؏a<�a<7�a<V�a<��a<��a<�a<�a<P�a<w�a<őa<��a<<�a<��a<a<�a<X�a<��a<��a<F�a<��a<�a<Y�a<��a<�a<k�a<��a<H�a<��a<�a<X�a<˘a<@�a<��a<�a<q�a<�a<L�a<�a<9�a<��a<)�a<��a<�a<m�a<�a<R�a<Οa<C�a<��a<+�a<��a<�a<v�a<�a<Y�a<��a<.�a<~�a<��a<U�a<��a<%�a<z�a<�a<5�a<��a<�a<P�a<��a<��a<a�a<��a<��a<)�a<x�a<��a<�a<O�a<|�a<٫a<�a<S�a<f�a<��a<�a<��a<@�a<Z�a<��a<��a<խa<��a<�a<F�a<Y�a<��a<��a<��a<ʮa<Ȯa<�a<��a<�a<�a< �a<-�a<3�a<H�a<)�a<X�a<E�a<C�a<L�a<-�a<P�a<�a<&�a<�a<%�a<�a<�a<�a<��a<ʮa<��a<��a<m�a<H�a<0�a<�a<��a<ĭa<��a<w�a<b�a<6�a<�a<�a<��a<��a<M�a<�a<�a<��a<��a<=�a<�a<Ūa<��a<Q�a<�a<�a<w�a<U�a<�a<��a<p�a<�a<ȧa<n�a<C�a<Ŧa<��a<#�a<ޥa<}�a<�a<Фa<R�a<�a<��a<8�a<آa<i�a<�a<��a<G�a<ؠa<v�a<�a<��a<8�a<��a<[�a<�a<�a<�a<��a<I�a<ƛa<�a<��a<��a<@�a<��a<s�a<�a<��a<#�a<Ɨa<[�a<	�a<��a<?�a<�a<��a<V�a<ܔa<��a<N�a<�a<��a<K�a<�a<��a<x�a<5�a<�a<Ña<}�a<W�a<�a<�a<��a<v�a<a�a<,�a<�a<�a<̏a<��a<��a<��a<]�a<z�a<Y�a<O�a<U�a<7�a<`�a<:�a<P�a<J�a<}�a<f�a<��a<��a<��a<�  �  ďa<��a<�a<8�a<X�a<��a<a<ϐa<2�a<R�a<~�a<ӑa<��a<>�a<x�a<Ȓa<�a<r�a<��a<
�a<_�a<��a<�a<R�a<��a<�a<t�a<ǖa<*�a<��a<�a<c�a<��a<;�a<��a<�a<��a<�a<L�a<Лa<1�a<��a<�a<��a<�a<~�a<�a<k�a<ٟa<E�a<Ԡa<(�a<��a<�a<o�a<ۢa<F�a<��a<(�a<��a<��a<z�a<ͥa<+�a<��a<�a<F�a<��a<�a<B�a<��a<�a<L�a<��a<ߩa<;�a<��a<ʪa<�a<>�a<��a<��a<��a<5�a<h�a<��a<֬a<�a<5�a<u�a<��a<ĭa<�a<��a<4�a<@�a<^�a<r�a<��a<��a<Үa<֮a<�a<�a<��a<&�a<*�a<.�a<<�a<>�a<E�a<4�a<F�a<5�a<J�a<&�a<3�a<;�a<!�a<$�a<�a<�a<��a<ˮa<Ȯa<��a<��a<��a<m�a<J�a<1�a<!�a<ܭa<�a<��a<~�a<p�a</�a<	�a<Ԭa<��a<~�a<g�a<�a<��a<ƫa<p�a<Z�a<
�a<̪a<��a<Z�a<�a<ɩa<��a<;�a<��a<��a<j�a< �a<Чa<��a<�a<Ħa<��a<�a<ѥa<e�a<#�a<��a<c�a<�a<��a<C�a<ڢa<��a<�a<��a<G�a<Ҡa<g�a<��a<��a<2�a<Ҟa<Y�a<�a<��a<�a<��a<B�a<כa<e�a<�a<��a<.�a<��a<^�a<�a<��a<5�a<ӗa<p�a<�a<��a<H�a<�a<��a<8�a<ޔa<��a<=�a<�a<��a<f�a<�a<Ғa<��a<4�a<�a<��a<��a<B�a<�a<ސa<��a<��a<`�a<S�a<�a<��a<֏a<��a<��a<��a<y�a<V�a<[�a<A�a<S�a<0�a<C�a<U�a<L�a<c�a<f�a<^�a<��a<��a<��a<�  �  ��a<�a< �a</�a<f�a<p�a<Őa<Ґa<�a<9�a<��a<��a<��a<Z�a<t�a<�a<��a<X�a<��a<�a<D�a<��a<
�a<8�a<ŕa<��a<m�a<ۖa<�a<��a<�a<s�a<Θa</�a<��a<��a<}�a<�a<t�a<̛a<G�a<��a<�a<��a<�a<��a<۞a<\�a<֟a<1�a<��a<�a<��a<�a<��a<�a<S�a<Уa<�a<��a<�a<X�a<��a<#�a<��a<Цa<]�a<��a<�a<K�a<��a<	�a<H�a<��a<�a<1�a<m�a<��a< �a<G�a<��a<��a<�a<+�a<y�a<��a<Ƭa<"�a<�a<q�a<��a<��a<֭a<�a<#�a</�a<}�a<p�a<��a<��a<��a<�a<׮a<��a<��a<+�a<�a<.�a<7�a<+�a<f�a<�a<a�a<@�a<F�a<L�a<,�a<0�a<�a<�a<�a<�a<��a<Ԯa<�a<��a<��a<t�a<e�a<Y�a<�a<#�a<߭a<ɭa<��a<��a<N�a<-�a<&�a<Ьa<Ϭa<o�a<L�a<�a<�a<��a<r�a<V�a<�a<�a<��a<T�a<�a<��a<��a<<�a<�a<��a<_�a<�a<��a<z�a<!�a<�a<~�a<1�a<�a<e�a<>�a<��a<q�a<�a<��a<A�a<Ţa<o�a<��a<��a<,�a<�a<x�a<�a<��a<�a<Ӟa<G�a<�a<s�a<�a<��a<*�a<�a<O�a<�a<��a<5�a<ԙa<Z�a<�a<��a<,�a<��a<`�a<�a<��a<_�a<�a<��a<.�a<�a<��a<-�a<�a<��a<b�a< �a<��a<y�a</�a<��a<��a<��a<@�a<+�a<�a<��a<��a<G�a<1�a<��a<�a<Ïa<��a<��a<u�a<��a<A�a<v�a<M�a<O�a<V�a<<�a<K�a<;�a<V�a<[�a<��a<��a<��a<Տa<�  �  Ǐa<�a< �a<9�a<\�a<��a<��a<��a<�a<[�a<��a<��a<��a<4�a<x�a<��a<�a<]�a<��a<
�a<N�a<��a<��a<P�a<��a<�a<V�a<��a</�a<��a<�a<M�a<Ęa<;�a<��a<!�a<�a<��a<P�a<��a<+�a<��a<�a<��a<��a<��a<�a<a�a<؟a<O�a<��a<8�a<��a<�a<t�a<Ԣa<D�a<��a<*�a<��a<	�a<a�a<˥a<-�a<��a<�a<U�a<��a<�a<C�a<��a<�a<=�a<��a<�a<6�a<��a<̪a<�a<F�a<u�a<��a<��a<=�a<c�a<��a<׬a<�a<5�a<d�a<��a<��a<�a<�a<$�a<E�a<S�a<q�a<��a<��a<®a<�a<��a<��a<�a<�a<%�a<-�a<>�a</�a<9�a<;�a<K�a<1�a<,�a<4�a<A�a<1�a<=�a<�a<�a<��a<׮a<ʮa<ˮa<��a<��a<t�a<o�a<N�a<-�a<�a<�a<έa<��a<��a<[�a<6�a<��a<Ԭa<��a<��a<Q�a<)�a<��a<��a<��a<D�a<�a<֪a<��a<=�a<�a<ͩa<��a<5�a<�a<��a<k�a<!�a<ܧa<|�a<0�a<Ȧa<o�a<�a<եa<k�a<�a<��a<p�a<��a<��a<B�a<�a<u�a< �a<��a<A�a<֠a<`�a<��a<��a<4�a<˞a<l�a<�a<��a<�a<��a<>�a<�a<c�a<�a<��a<0�a<��a<P�a<�a<��a<1�a<ٗa<r�a<�a<��a<8�a<�a<��a<@�a<ؔa<{�a<>�a<��a<��a<U�a<�a<ƒa<��a<H�a<��a<a<w�a<A�a<�a<�a<��a<��a<l�a<7�a<#�a<�a<яa<��a<��a<z�a<m�a<]�a<`�a<=�a<4�a<>�a<Q�a<K�a<g�a<[�a<n�a<k�a<o�a<��a<��a<�  �  ��a<��a<�a<�a<�a<[�a<_�a<��a<Ɛa<�a<3�a<x�a<��a<��a<��a<u�a<ڒa<�a<p�a<a<�a<v�a<��a<+�a<`�a<ʕa<:�a<��a<��a<H�a<ޗa< �a<��a<�a<b�a<�a<6�a<ʚa<�a<��a<��a<n�a<�a<m�a<��a<*�a<��a<1�a<��a<&�a<m�a<�a<F�a<�a<'�a<עa<R�a<n�a<
�a<C�a<ۤa<�a<��a<�a<T�a<¦a<��a<~�a<ۧa<*�a<q�a<��a<;�a<Y�a<ѩa<��a<O�a<��a<۪a<#�a<H�a<��a<��a<�a<F�a<��a<��a<Ŭa<�a<!�a<h�a<��a<��a<حa<ѭa< �a<�a<��a<k�a<k�a<��a<��a<ˮa<��a<��a<ڮa<�a<��a<�a<"�a<�a<�a<�a<�a<#�a<��a<�a<�a<�a<Ԯa<�a<®a<Ʈa<��a<��a<��a<o�a<f�a<&�a<�a<�a<˭a<٭a<��a<��a<A�a<#�a<��a<Ӭa<��a<k�a<W�a<�a<�a<��a<��a<_�a<�a<�a<��a<[�a<,�a<�a<��a<H�a<1�a<èa<��a<@�a<�a<��a<;�a<�a<��a<n�a<�a<��a<L�a<��a<��a<�a<գa<s�a<��a<��a<-�a<��a<W�a<�a<��a<b�a<�a<K�a<�a<u�a<:�a<��a<`�a<ٜa<r�a<�a<��a<A�a<ښa<f�a<�a<��a<C�a<��a<p�a<�a<��a<,�a<Жa<w�a<��a<ԕa<F�a<��a<��a<b�a<�a<��a<v�a<�a<גa<��a<@�a<�a<��a<��a<,�a<U�a<ܐa<��a<s�a<2�a<,�a<�a<�a<��a<��a<o�a<F�a<]�a<9�a</�a<�a<�a<�a<��a<�a<�a<�a<�a<9�a<(�a<O�a<h�a<f�a<�  �  ��a<��a<Ϗa<��a<#�a<H�a<k�a<��a<Ԑa<�a<D�a<��a<֑a<�a<0�a<z�a<�a<%�a<|�a<��a<�a<g�a<��a<�a<y�a<ؕa<1�a<��a<��a<g�a<a<!�a<��a<�a<m�a<��a<G�a<��a<�a<��a<�a<��a<�a<^�a<̝a<K�a<��a<7�a<��a<�a<z�a<�a<^�a<�a<H�a<��a<	�a<��a<�a<X�a<פa<*�a<��a<�a<c�a<��a<�a<l�a<̧a<�a<��a<ըa<�a<X�a<��a<	�a<U�a<��a<ߪa<�a<M�a<��a<ܫa<�a<;�a<v�a<��a<߬a<
�a<6�a<\�a<��a<��a<߭a<�a<)�a<"�a<5�a<K�a<��a<��a<��a<Ʈa<ɮa<�a<�a<��a<�a<�a<
�a<�a<�a<&�a<�a<�a<��a<�a<��a<�a<�a<�a<��a<��a<��a<��a<��a<k�a<R�a<A�a<$�a<�a<حa<ŭa<��a<��a<R�a<<�a<�a<��a<��a<o�a<k�a<&�a<��a<��a<��a<P�a<�a<ݪa<��a<i�a<#�a<ݩa<��a<g�a<�a<Ĩa<~�a<=�a<�a<��a<M�a<��a<��a<O�a<��a<��a<<�a<�a<��a<5�a<ԣa<y�a<�a<��a<;�a<�a<o�a<(�a<��a<(�a<��a<c�a<�a<��a<5�a<��a<U�a<ܜa<��a<�a<��a</�a<ʚa<W�a<�a<��a<%�a<��a<\�a<��a<��a<4�a<Ԗa<n�a<�a<��a<d�a<�a<��a<U�a<�a<��a<e�a<�a<̒a<��a<>�a<�a<��a<��a<7�a<��a<��a<��a<��a<B�a<'�a<�a<؏a<��a<��a<~�a<g�a<E�a<4�a<#�a<,�a<�a<�a<��a<�a<	�a<�a<�a</�a<'�a<G�a<[�a<��a<�  �  ~�a<ɏa<ɏa<��a<�a<>�a<��a<��a<�a<�a<C�a<u�a<��a<�a<D�a<��a<ǒa<�a<l�a<��a<�a<[�a<єa<
�a<|�a<̕a<?�a<��a<�a<f�a<��a<@�a<��a<��a<b�a<řa<H�a<��a<7�a<��a<�a<{�a<ܜa<~�a<Ɲa<W�a<��a<5�a<��a<�a<��a<�a<e�a<ša<P�a<��a<)�a<��a<�a<^�a<��a<8�a<��a<�a<h�a<��a<&�a<f�a<�a<�a<t�a<Ϩa<�a<��a<��a<
�a<=�a<��a<ܪa<�a<r�a<��a<ܫa< �a<K�a<��a<��a<�a<��a<H�a<S�a<��a<��a<˭a<�a<��a<K�a<P�a<t�a<��a<��a<��a<��a<ڮa<ծa<��a<�a< �a<�a<��a</�a<�a<�a<�a< �a<�a< �a<��a<�a<�a<ٮa<Ӯa<Ѯa<��a<��a<q�a<��a<L�a<B�a< �a<��a<�a<��a<��a<r�a<Q�a<!�a<�a<�a<��a<��a<E�a<�a<�a<��a<��a<C�a<)�a<Ϊa<��a<]�a<1�a<�a<��a<f�a< �a<�a<��a<7�a<�a<��a<N�a<��a<��a<R�a<��a<��a<6�a<	�a<��a<A�a<£a<w�a<�a<��a<P�a<֡a<v�a<��a<��a<H�a<ܟa<z�a<�a<��a< �a<ĝa<V�a<ߜa<��a<��a<��a<*�a<�a<V�a<�a<��a<$�a<Ԙa<T�a<��a<��a<#�a<іa<n�a<(�a<��a<c�a<��a<��a<i�a<��a<��a<R�a<+�a<a<��a<<�a<��a<��a<m�a<`�a<�a<�a<��a<f�a<E�a<�a<�a<ʏa<��a<��a<w�a<m�a<9�a<S�a<�a<$�a<�a<�a<�a<�a<�a<��a<�a<!�a<:�a<Z�a<J�a<��a<�  �  ��a<��a<Əa<��a<"�a<P�a<q�a<��a<Րa<	�a<P�a<��a<��a<��a<N�a<��a<ɒa</�a<s�a<��a<�a<_�a<��a<�a<|�a<a<'�a<��a<��a<U�a<��a<)�a<��a<�a<n�a<�a<C�a<��a<�a<��a<��a<|�a<�a<a�a<ŝa<F�a<��a<1�a<��a<�a<}�a<�a<v�a<ڡa<5�a<��a<$�a<��a<��a<s�a<Ǥa<(�a<��a<�a<[�a<��a<�a<g�a<̧a<&�a<|�a<Ĩa<�a<e�a<��a<�a<X�a<��a<ݪa<�a<V�a<��a<ͫa<�a<E�a<p�a<��a<�a<�a<2�a<W�a<��a<��a<ԭa<�a<
�a<&�a<S�a<b�a<m�a<��a<��a<��a<Ȯa<׮a<�a<��a<�a<�a< �a<�a<�a<�a<�a<�a<
�a<�a<��a<�a<�a<�a<Ǯa<��a<��a<��a<��a<p�a<I�a<5�a<#�a<	�a<ޭa<��a<��a<v�a<^�a<8�a<�a<Ԭa<��a<w�a<F�a<0�a<��a<��a<��a<G�a<�a<�a<��a<S�a<�a<�a<��a<U�a<�a<̨a<~�a<<�a<�a<��a<H�a<��a<��a<S�a<�a<��a<K�a<�a<��a<0�a<ԣa<s�a<�a<��a<>�a<١a<��a<�a<��a<?�a<ןa<]�a<�a<��a<%�a<��a<O�a<ܜa<z�a<�a<��a<+�a<˚a<c�a<��a<��a<'�a<��a<W�a<��a<��a<5�a<Ӗa<h�a<�a<��a<U�a<�a<��a<N�a<��a<��a<i�a<�a<ƒa<��a<;�a<�a<ϑa<x�a<;�a<�a<Ӑa<��a<}�a<V�a<�a<�a<̏a<��a<��a<}�a<\�a<;�a<9�a<0�a<�a<�a<�a<�a<�a<�a<�a<�a<,�a<-�a<J�a<S�a<w�a<�  �  ��a<��a<��a<��a<�a<F�a<g�a<��a<Аa<�a<7�a<��a<̑a<��a<M�a<��a<�a<�a<n�a<��a<�a<�a<��a<�a<p�a<�a<3�a<��a<�a<K�a<֗a<&�a<��a<��a<Y�a<�a<1�a<Ěa<�a<��a<�a<}�a<��a<I�a<�a<B�a<��a<"�a<��a<�a<{�a<��a<S�a<�a<J�a<��a<#�a<��a<�a<P�a<Ѥa<+�a<��a<�a<M�a<��a<�a<��a<��a<)�a<��a<Ȩa<1�a<[�a<ɩa<�a<U�a<��a<Ъa<(�a<Q�a<��a<īa<�a<:�a<r�a<��a<Ԭa<	�a<%�a<t�a<��a<��a<ԭa<�a<#�a<'�a<O�a<c�a<��a<��a<��a<Ȯa<Ǯa<�a<�a<��a<��a<	�a<#�a<��a<!�a<�a<�a<�a<�a<�a<�a<
�a<Ӯa<�a<ʮa<îa<��a<��a<��a<U�a<c�a<>�a<�a<��a<ԭa<׭a<��a<��a<F�a<0�a<�a<լa<��a<w�a<a�a<�a<�a<��a<�a<g�a<�a<۪a<��a<s�a<%�a<ҩa<��a<K�a<)�a<ɨa<��a<4�a<٧a<��a<7�a<�a<��a<`�a<��a<��a<O�a<դa<��a<+�a<ӣa<e�a<�a<��a<<�a<�a<d�a<�a<��a<@�a<֟a<j�a<�a<��a<0�a<��a<U�a<�a<k�a<�a<��a<K�a<��a<f�a<��a<��a<9�a<��a<h�a<�a<��a<%�a<Ɩa<|�a<�a<ȕa<L�a<�a<��a<Q�a<�a<��a<e�a<�a<�a<��a<@�a<�a<��a<��a<<�a<�a<Ԑa<��a<~�a<7�a<)�a<��a<�a<��a<��a<u�a<`�a<^�a<�a<3�a<�a<�a<�a<��a<�a<��a<%�a<�a<0�a<1�a<L�a<j�a<k�a<�  �  ��a<��a<ُa<��a<�a<F�a<|�a<��a<ϐa<�a<L�a<|�a<��a<�a<E�a<��a<͒a<�a<u�a<��a<�a<l�a<Ɣa<�a<q�a<ӕa<;�a<��a<��a<_�a<��a<�a<��a<��a<k�a<�a<H�a<��a< �a<��a<�a<v�a<�a<d�a<֝a<F�a<��a<+�a<��a<�a<��a<��a<m�a<͡a<F�a<��a<$�a<��a<�a<f�a<Ϥa<.�a<��a<�a<W�a<��a<�a<u�a<ѧa<(�a<u�a<ͨa<!�a<j�a<��a<�a<W�a<��a<תa<�a<S�a<��a<֫a<�a<J�a<~�a<��a<ڬa<
�a<8�a<g�a<��a<��a<խa<�a<�a<:�a<N�a<o�a<}�a<��a<��a<îa<Ǯa<�a<��a<��a<��a<�a<�a<�a<�a<�a<�a<�a<�a<�a<��a<�a<�a<ܮa<ɮa<��a<��a<��a<��a<o�a<\�a<5�a<�a< �a<�a<ŭa<��a<~�a<Z�a<'�a<��a<�a<��a<��a<J�a<�a<��a<��a<��a<U�a<�a<ܪa<��a<e�a<-�a<�a<��a<_�a<�a<¨a<��a<7�a<�a<��a<M�a<��a<��a<Q�a<��a<��a<I�a<�a<��a<0�a<ԣa<m�a<�a<��a<B�a<�a<~�a<�a<��a<B�a<ןa<m�a<��a<��a<.�a<��a<N�a<�a<v�a<�a<��a<8�a<Кa<d�a<�a<��a<)�a<��a<Z�a<��a<��a<1�a<͖a<n�a<
�a<��a<]�a<�a<��a<\�a<�a<��a<f�a<�a<גa<��a<?�a<�a<��a<y�a<P�a<�a<��a<��a<o�a<N�a<$�a<��a<Տa<��a<��a<v�a<Y�a<Q�a<<�a<&�a<�a<�a<�a<��a<�a<�a<�a<�a<%�a</�a<>�a<X�a<w�a<�  �  ��a<��a<ŏa<�a<'�a<<�a<w�a<��a<�a< �a<N�a<��a<��a<�a<*�a<��a<Βa<5�a<m�a<��a< �a<W�a<a<	�a<��a<ӕa<'�a<��a<�a<g�a<��a<6�a<��a<��a<h�a<��a<K�a<��a<=�a<��a<�a<��a<�a<_�a<ĝa<[�a<��a<$�a<��a<�a<��a<�a<|�a<ѡa<H�a<��a<�a<��a<�a<x�a<��a<4�a<��a<�a<R�a<��a<-�a<g�a<ǧa<�a<z�a<Ψa<�a<��a<��a<
�a<<�a<��a<٪a<�a<l�a<��a<ޫa<�a<@�a<n�a<��a<�a<��a<6�a<S�a<��a<��a<ɭa<�a<�a<8�a<5�a<i�a<~�a<��a<��a<��a<ݮa<ήa<�a<�a<�a<�a< �a<�a<�a<%�a<	�a<�a<�a< �a<	�a<خa<�a<֮a<ۮa<îa<��a<��a<s�a<p�a<H�a<E�a<(�a<��a<�a<��a<��a<l�a<\�a<8�a< �a<�a<��a<��a<L�a<6�a<�a<��a<��a<?�a<�a<ͪa<��a<d�a<�a<�a<��a<f�a<�a<٨a<��a<5�a<�a<��a<P�a<�a<��a<C�a<��a<��a<<�a<�a<�a<D�a<ˣa<f�a<�a<��a<N�a<ˡa<��a<
�a<��a<6�a<ǟa<n�a<��a<��a<�a<��a<N�a<ޜa<q�a<�a<��a<*�a<Śa<Y�a<��a<��a<�a<טa<L�a<��a<�a<(�a<ϖa<j�a<#�a<��a<e�a<��a<��a<L�a< �a<œa<U�a<�a<a<��a<=�a<��a<בa<v�a<N�a<��a<ڐa<��a<y�a<T�a<�a<�a<Ïa<��a<��a<}�a<m�a<;�a<<�a<�a<*�a<�a<�a<�a<�a<�a<�a< �a<�a<A�a<L�a<N�a<��a<�  �  ��a<��a<Ϗa<�a<�a<O�a<x�a<��a<ܐa<�a<=�a<��a<a<�a<R�a<��a<ђa<�a<n�a<a<�a<h�a<Ŕa< �a<q�a<ҕa<1�a<��a<��a<T�a<Ɨa</�a<��a<��a<p�a<ؙa<L�a<��a<$�a<��a<�a<t�a<��a<_�a<ӝa<E�a<��a<1�a<��a<�a<��a<��a<a�a<סa<F�a<��a<+�a<��a<��a<]�a<̤a<2�a<��a<��a<^�a<��a<�a<u�a<ʧa<.�a<v�a<˨a<"�a<q�a<��a<	�a<P�a<��a<֪a<�a<`�a<��a<ϫa<�a<L�a<w�a<��a<ڬa<�a<:�a<b�a<��a<��a<ҭa<�a<�a<3�a<Z�a<j�a<��a<��a<��a<��a<ծa<�a<�a< �a<�a<�a<�a<�a<�a<�a<�a<�a<�a<��a<�a<�a<�a<Үa<Ʈa<îa<��a<��a<��a<s�a<R�a<8�a<�a<�a<�a<­a<��a<x�a<L�a<+�a<�a<۬a<��a<��a<N�a<�a<�a<��a<��a<Q�a<�a<�a<��a<c�a<#�a<�a<��a<T�a<�a<Ҩa<z�a<3�a<�a<��a<Q�a<�a<��a<S�a<��a<��a<O�a<�a<��a<.�a<ңa<s�a<�a<��a<F�a<�a<r�a<�a<��a<C�a<ޟa<k�a<�a<��a<+�a<��a<L�a<�a<}�a<�a<��a<9�a<ɚa<k�a<��a<��a<+�a<Øa<O�a<��a<��a<4�a<˖a<e�a<�a<��a<W�a<�a<��a<U�a<�a<��a<j�a<�a<ђa<��a<B�a< �a<��a<�a<H�a<�a<ېa<��a<u�a<@�a<�a<��a<Տa<��a<��a<y�a<\�a<G�a<?�a<+�a<�a<�a<�a<��a<��a<�a<�a<�a<�a<,�a<L�a<_�a<j�a<�  �  ��a<��a<Ϗa<��a<$�a<T�a<_�a<��a<͐a<�a<K�a<��a<ʑa<�a<Z�a<z�a<�a<�a<z�a<ȓa<�a<s�a<��a<.�a<s�a<ѕa<.�a<��a<�a<R�a<ʗa<�a<��a<�a<e�a<יa<;�a<Ěa<�a<��a<�a<w�a<��a<N�a<ԝa<>�a<Ξa<$�a<��a<�a<w�a<
�a<[�a<�a<<�a<��a<%�a<~�a<�a<Q�a<ݤa<)�a<��a<��a<M�a<Φa<�a<u�a<��a<2�a<z�a<Ȩa<$�a<]�a<ʩa< �a<N�a<��a<ݪa<'�a<E�a<��a<ɫa<�a<E�a<p�a<��a<جa<�a<�a<i�a<��a<��a<�a<�a<#�a<�a<^�a<U�a<��a<��a<��a<Үa<��a<�a<ٮa<��a<�a<�a<�a<�a<,�a<�a<�a<�a<
�a<�a<��a<��a<�a<�a<Ϯa<��a<��a<��a<��a<^�a<R�a<5�a<%�a<�a<̭a<ҭa<��a<��a<Y�a<.�a<�a<Ŭa<ìa<p�a<b�a<�a<��a<ūa<��a<[�a<��a<�a<��a<b�a< �a<ݩa<��a<R�a<�a<��a<��a<>�a<�a<��a<@�a<�a<��a<T�a<��a<��a<Y�a<ڤa<��a<'�a<�a<f�a<	�a<��a<7�a<�a<l�a< �a<��a<8�a<؟a<Z�a<�a<��a<;�a<��a<Z�a<�a<l�a<"�a<��a<9�a<��a<n�a<��a<��a<,�a<��a<i�a<�a<��a<-�a<Җa<{�a<��a<��a<Q�a<�a<��a<N�a<�a<��a<z�a<�a<ؒa<��a<D�a<�a<��a<��a<4�a<�a<Ɛa<��a<�a<I�a<2�a<�a<�a<��a<��a<��a<[�a<G�a<(�a<?�a<�a<�a<�a<�a<�a< �a<�a<�a<0�a<5�a<9�a<b�a<k�a<�  �  ��a<��a<ُa<��a<�a<>�a<x�a<��a<ؐa<�a<J�a<z�a<ȑa<�a<R�a<��a<ܒa<�a<s�a<��a<�a<q�a<��a<�a<q�a<֕a<6�a<��a<�a<S�a<��a<7�a<��a<�a<f�a<ܙa<8�a<��a<7�a<��a< �a<~�a<�a<^�a<םa<L�a<��a<&�a<��a<�a<�a<��a<a�a<ѡa<K�a<��a<+�a<��a<��a<Z�a<Ȥa<)�a<��a<��a<W�a<��a<�a<v�a<̧a<�a<y�a<Ĩa<�a<�a<��a<��a<Q�a<��a<Ūa<�a<h�a<��a<̫a<	�a<=�a<}�a<��a<ڬa<��a<6�a<f�a<��a<��a<խa<�a<�a<.�a<\�a<m�a<��a<��a<��a<��a<ˮa<�a<�a<�a<��a<�a<�a<�a<�a<�a<�a<�a<�a<��a<��a<��a<�a<̮a<ٮa<Įa<��a<��a<{�a<h�a<\�a<@�a<�a<��a<�a<˭a<��a<r�a<X�a<&�a<�a<ݬa<��a<~�a<Y�a<!�a<��a<��a<��a<Y�a<�a<̪a<��a<g�a<(�a<ݩa<��a<R�a<�a<ڨa<��a<"�a<�a<��a<>�a<�a<��a<Q�a<�a<��a<>�a<�a<��a<5�a<£a<h�a<�a<��a<?�a<ݡa<r�a<
�a<��a<F�a<ޟa<k�a<��a<��a<'�a<��a<S�a<�a<v�a< �a<��a<:�a<˚a<X�a<��a<��a<$�a<јa<W�a<�a<��a<.�a<��a<r�a<�a<��a<S�a<��a<��a<[�a<�a<��a<V�a<�a<Ւa<��a<5�a<�a<��a<��a<C�a<�a<ސa<��a<q�a<K�a<�a<�a<ߏa<��a<��a<k�a<g�a<O�a<1�a<�a<�a<�a<�a<�a<��a< �a<�a<�a<�a<?�a<M�a<W�a<s�a<�  �  ��a<��a<Əa<��a<"�a<E�a<��a<��a<�a<��a<\�a<��a<��a<��a<3�a<��a<Вa<,�a<{�a<��a<�a<Y�a<ݔa<�a<��a<ϕa<-�a<��a<�a<f�a<��a<%�a<��a<�a<v�a<ڙa<]�a<��a<�a<��a<�a<��a<�a<r�a<��a<T�a<��a<@�a<��a<�a<��a<�a<�a<աa<K�a<��a<�a<��a<��a<x�a<Ĥa<5�a<��a<�a<r�a<��a<&�a<`�a<ܧa<�a<�a<Ѩa<�a<h�a<��a<�a<S�a<��a<�a<�a<X�a<��a<߫a<�a<E�a<|�a<��a<�a<��a<T�a<O�a<��a<��a<֭a<�a<�a<3�a<<�a<c�a<�a<��a<®a<��a<ܮa<Үa<��a< �a<��a<�a<�a<$�a<�a<�a<�a<�a<�a<��a<�a<�a<��a<׮a<��a<��a<��a<��a<w�a<}�a<I�a<>�a<#�a<��a<��a<��a<��a<h�a<j�a<4�a<�a<جa<��a<��a<M�a<.�a<��a<��a<��a<A�a<5�a<̪a<��a<`�a<�a<�a<��a<f�a<
�a<Ȩa<o�a<=�a<��a<��a<c�a<�a<��a<G�a<��a<��a<;�a<��a<{�a<=�a<ǣa<��a<�a<��a<M�a<ӡa<��a<�a<��a<2�a<şa<p�a<��a<��a<#�a<��a<H�a<ݜa<��a<�a<��a<#�a<ۚa<Y�a<��a<��a<�a<��a<C�a<�a<��a<:�a<֖a<[�a<�a<��a<g�a<�a<��a<[�a<��a<ēa<W�a<8�a<��a<��a<<�a<�a<ϑa<}�a<H�a<��a<Ԑa<��a<|�a<`�a<�a<�a<Ǐa<ŏa<��a<v�a<g�a<=�a<H�a<�a<$�a<	�a<�a<��a<��a<�a<
�a<'�a<�a<'�a<C�a<T�a<~�a<�  �  ��a<��a<ҏa<��a<$�a<F�a<s�a<��a<�a<�a<F�a<y�a<ʑa<�a<T�a<��a<�a<�a<r�a<��a<$�a<b�a<��a<�a<{�a<ؕa<4�a<��a<��a<S�a<ɗa<�a<��a<
�a<M�a<��a<6�a<ʚa<�a<��a<�a<x�a<�a<b�a<ӝa<I�a<��a<*�a<��a<�a<��a<��a<X�a<ءa<L�a<��a<(�a<��a<��a<N�a<ʤa<:�a<��a<�a<X�a<��a<�a<t�a<ԧa<�a<|�a<Ǩa<*�a<d�a<ѩa<��a<4�a<|�a<ݪa<1�a<Q�a<��a<ȫa<�a<9�a<��a<��a<�a<�a<4�a<V�a<��a<��a<ҭa<ޭa<�a<4�a<X�a<j�a<��a<��a<��a<��a<ݮa<�a<�a<��a<�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<߮a<Ѯa<�a<ٮa<��a<��a<��a<��a<d�a<U�a<@�a<%�a<��a<�a<��a<��a<|�a<T�a<$�a<�a<ܬa<��a<��a<^�a<�a<�a<��a<��a<K�a<�a<תa<��a<i�a<&�a<שa<��a<S�a<�a<¨a<��a<D�a<ͧa<��a<;�a<�a<��a<\�a<��a<��a<B�a<�a<��a<3�a<Σa<m�a<�a<��a<N�a<ߡa<i�a<�a<��a<E�a<۟a<o�a<�a<��a<(�a<Ɲa<^�a<ܜa<w�a<�a<��a<7�a<Қa<X�a<��a<��a<2�a<��a<p�a<�a<w�a<�a<Җa<��a<�a<��a<O�a<�a<��a<_�a<�a<��a<^�a<�a<Œa<��a<G�a< �a<��a<��a<I�a<�a<ېa<��a<r�a<D�a< �a<�a<Տa<��a<��a<�a<d�a<K�a<3�a<)�a<�a<�a<�a<�a<�a<��a<��a< �a<:�a<?�a<G�a<a�a<p�a<�  �  ��a<��a<�a<�a<�a<W�a<y�a<��a<ǐa<�a<K�a<z�a<ӑa<�a<U�a<t�a<�a<�a<��a<��a<�a<o�a<Ĕa<+�a<Y�a<˕a<<�a<��a<�a<B�a<Зa<�a<��a<�a<s�a<�a<(�a<Ěa<�a<��a<�a<��a<�a<N�a<�a</�a<��a<9�a<��a<�a<p�a<�a<S�a<�a<C�a<��a<!�a<��a<�a<N�a<�a<�a<��a<��a<g�a<��a<��a<�a<��a<�a<��a<��a<,�a<N�a<Ωa<�a<��a<��a<��a<�a<;�a<��a<��a<#�a<3�a<�a<��a<��a<�a<A�a<f�a<z�a<��a<�a<�a<(�a< �a<Z�a<_�a<��a<��a<��a<ٮa<��a<�a<�a<�a<��a<��a<!�a<��a<&�a<�a<�a<�a<�a<�a<�a<F�a<ݮa<Үa<��a<��a<��a<��a<��a<W�a<i�a<.�a<�a<�a<�a<ɭa<��a<��a<Y�a<%�a<�a<ˬa<��a<j�a<j�a<�a<�a<��a<y�a<W�a<�a<�a<��a<\�a<.�a<ҩa<��a<B�a<#�a<��a<��a<�a<�a<ܧa<.�a<�a<��a<Z�a<��a<��a<I�a<٤a<��a<�a<ңa<{�a<�a<��a<0�a<��a<d�a<�a<��a<=�a<ԟa<`�a<�a<��a<F�a<��a<J�a<�a<��a<�a<��a<B�a<��a<X�a<�a<�a<4�a<��a<m�a<ԗa<Ǘa<J�a<��a<s�a<�a<ɕa<A�a<�a<��a<]�a<�a<��a<s�a<$�a<Ւa<y�a<<�a<�a<��a<��a<5�a<�a<Аa<��a<v�a<E�a<:�a<�a<׏a<��a<��a<o�a<M�a<\�a<"�a<8�a<�a<�a<�a<�a<�a<��a<a�a<�a<�a<%�a<6�a<b�a<e�a<�  �  ��a<��a<ҏa<��a<$�a<F�a<s�a<��a<�a<�a<F�a<y�a<ʑa<�a<T�a<��a<�a<�a<r�a<��a<$�a<b�a<��a<�a<{�a<ؕa<4�a<��a<��a<S�a<ɗa<�a<��a<
�a<M�a<��a<6�a<ʚa<�a<��a<�a<x�a<�a<b�a<ӝa<I�a<��a<*�a<��a<�a<��a<��a<X�a<ءa<L�a<��a<(�a<��a<��a<N�a<ʤa<:�a<��a<�a<X�a<��a<�a<t�a<ԧa<�a<|�a<Ǩa<*�a<d�a<ѩa<��a<4�a<|�a<ݪa<1�a<Q�a<��a<ȫa<�a<9�a<��a<��a<�a<�a<4�a<V�a<��a<��a<ҭa<ޭa<�a<4�a<X�a<j�a<��a<��a<��a<��a<ݮa<�a<�a<��a<�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<߮a<Ѯa<�a<ٮa<��a<��a<��a<��a<d�a<U�a<@�a<%�a<��a<�a<��a<��a<|�a<T�a<$�a<�a<ܬa<��a<��a<^�a<�a<�a<��a<��a<K�a<�a<תa<��a<i�a<&�a<שa<��a<S�a<�a<¨a<��a<D�a<ͧa<��a<;�a<�a<��a<\�a<��a<��a<B�a<�a<��a<3�a<Σa<m�a<�a<��a<N�a<ߡa<i�a<�a<��a<E�a<۟a<o�a<�a<��a<(�a<Ɲa<^�a<ܜa<w�a<�a<��a<7�a<Қa<X�a<��a<��a<2�a<��a<p�a<�a<w�a<�a<Җa<��a<�a<��a<O�a<�a<��a<_�a<�a<��a<^�a<�a<Œa<��a<G�a< �a<��a<��a<I�a<�a<ېa<��a<r�a<D�a< �a<�a<Տa<��a<��a<�a<d�a<K�a<3�a<)�a<�a<�a<�a<�a<�a<��a<��a< �a<:�a<?�a<G�a<a�a<p�a<�  �  ��a<��a<Əa<��a<"�a<E�a<��a<��a<�a<��a<\�a<��a<��a<��a<3�a<��a<Вa<,�a<{�a<��a<�a<Y�a<ݔa<�a<��a<ϕa<-�a<��a<�a<f�a<��a<%�a<��a<�a<v�a<ڙa<]�a<��a<�a<��a<�a<��a<�a<r�a<��a<T�a<��a<@�a<��a<�a<��a<�a<�a<աa<K�a<��a<�a<��a<��a<x�a<Ĥa<5�a<��a<�a<r�a<��a<&�a<`�a<ܧa<�a<�a<Ѩa<�a<h�a<��a<�a<S�a<��a<�a<�a<X�a<��a<߫a<�a<E�a<|�a<��a<�a<��a<T�a<O�a<��a<��a<֭a<�a<�a<3�a<<�a<c�a<�a<��a<®a<��a<ܮa<Үa<��a< �a<��a<�a<�a<$�a<�a<�a<�a<�a<�a<��a<�a<�a<��a<׮a<��a<��a<��a<��a<w�a<}�a<I�a<>�a<#�a<��a<��a<��a<��a<h�a<j�a<4�a<�a<جa<��a<��a<M�a<.�a<��a<��a<��a<A�a<5�a<̪a<��a<`�a<�a<�a<��a<f�a<
�a<Ȩa<o�a<=�a<��a<��a<c�a<�a<��a<G�a<��a<��a<;�a<��a<{�a<=�a<ǣa<��a<�a<��a<M�a<ӡa<��a<�a<��a<2�a<şa<p�a<��a<��a<#�a<��a<H�a<ݜa<��a<�a<��a<#�a<ۚa<Y�a<��a<��a<�a<��a<C�a<�a<��a<:�a<֖a<[�a<�a<��a<g�a<�a<��a<[�a<��a<ēa<W�a<8�a<��a<��a<<�a<�a<ϑa<}�a<H�a<��a<Ԑa<��a<|�a<`�a<�a<�a<Ǐa<ŏa<��a<v�a<g�a<=�a<H�a<�a<$�a<	�a<�a<��a<��a<�a<
�a<'�a<�a<'�a<C�a<T�a<~�a<�  �  ��a<��a<ُa<��a<�a<>�a<x�a<��a<ؐa<�a<J�a<z�a<ȑa<�a<R�a<��a<ܒa<�a<s�a<��a<�a<q�a<��a<�a<q�a<֕a<6�a<��a<�a<S�a<��a<7�a<��a<�a<f�a<ܙa<8�a<��a<7�a<��a< �a<~�a<�a<^�a<םa<L�a<��a<&�a<��a<�a<�a<��a<a�a<ѡa<K�a<��a<+�a<��a<��a<Z�a<Ȥa<)�a<��a<��a<W�a<��a<�a<v�a<̧a<�a<y�a<Ĩa<�a<�a<��a<��a<Q�a<��a<Ūa<�a<h�a<��a<̫a<	�a<=�a<}�a<��a<ڬa<��a<6�a<f�a<��a<��a<խa<�a<�a<.�a<\�a<m�a<��a<��a<��a<��a<ˮa<�a<�a<�a<��a<�a<�a<�a<�a<�a<�a<�a<�a<��a<��a<��a<�a<̮a<ٮa<Įa<��a<��a<{�a<h�a<\�a<@�a<�a<��a<�a<˭a<��a<r�a<X�a<&�a<�a<ݬa<��a<~�a<Y�a<!�a<��a<��a<��a<Y�a<�a<̪a<��a<g�a<(�a<ݩa<��a<R�a<�a<ڨa<��a<"�a<�a<��a<>�a<�a<��a<Q�a<�a<��a<>�a<�a<��a<5�a<£a<h�a<�a<��a<?�a<ݡa<r�a<
�a<��a<F�a<ޟa<k�a<��a<��a<'�a<��a<S�a<�a<v�a< �a<��a<:�a<˚a<X�a<��a<��a<$�a<јa<W�a<�a<��a<.�a<��a<r�a<�a<��a<S�a<��a<��a<[�a<�a<��a<V�a<�a<Ւa<��a<5�a<�a<��a<��a<C�a<�a<ސa<��a<q�a<K�a<�a<�a<ߏa<��a<��a<k�a<g�a<O�a<1�a<�a<�a<�a<�a<�a<��a< �a<�a<�a<�a<?�a<M�a<W�a<s�a<�  �  ��a<��a<Ϗa<��a<$�a<T�a<_�a<��a<͐a<�a<K�a<��a<ʑa<�a<Z�a<z�a<�a<�a<z�a<ȓa<�a<s�a<��a<.�a<s�a<ѕa<.�a<��a<�a<R�a<ʗa<�a<��a<�a<e�a<יa<;�a<Ěa<�a<��a<�a<w�a<��a<N�a<ԝa<>�a<Ξa<$�a<��a<�a<w�a<
�a<[�a<�a<<�a<��a<%�a<~�a<�a<Q�a<ݤa<)�a<��a<��a<M�a<Φa<�a<u�a<��a<2�a<z�a<Ȩa<$�a<]�a<ʩa< �a<N�a<��a<ݪa<'�a<E�a<��a<ɫa<�a<E�a<p�a<��a<جa<�a<�a<i�a<��a<��a<�a<�a<#�a<�a<^�a<U�a<��a<��a<��a<Үa<��a<�a<ٮa<��a<�a<�a<�a<�a<,�a<�a<�a<�a<
�a<�a<��a<��a<�a<�a<Ϯa<��a<��a<��a<��a<^�a<R�a<5�a<%�a<�a<̭a<ҭa<��a<��a<Y�a<.�a<�a<Ŭa<ìa<p�a<b�a<�a<��a<ūa<��a<[�a<��a<�a<��a<b�a< �a<ݩa<��a<R�a<�a<��a<��a<>�a<�a<��a<@�a<�a<��a<T�a<��a<��a<Y�a<ڤa<��a<'�a<�a<f�a<	�a<��a<7�a<�a<l�a< �a<��a<8�a<؟a<Z�a<�a<��a<;�a<��a<Z�a<�a<l�a<"�a<��a<9�a<��a<n�a<��a<��a<,�a<��a<i�a<�a<��a<-�a<Җa<{�a<��a<��a<Q�a<�a<��a<N�a<�a<��a<z�a<�a<ؒa<��a<D�a<�a<��a<��a<4�a<�a<Ɛa<��a<�a<I�a<2�a<�a<�a<��a<��a<��a<[�a<G�a<(�a<?�a<�a<�a<�a<�a<�a< �a<�a<�a<0�a<5�a<9�a<b�a<k�a<�  �  ��a<��a<Ϗa<�a<�a<O�a<x�a<��a<ܐa<�a<=�a<��a<a<�a<R�a<��a<ђa<�a<n�a<a<�a<h�a<Ŕa< �a<q�a<ҕa<1�a<��a<��a<T�a<Ɨa</�a<��a<��a<p�a<ؙa<L�a<��a<$�a<��a<�a<t�a<��a<_�a<ӝa<E�a<��a<1�a<��a<�a<��a<��a<a�a<סa<F�a<��a<+�a<��a<��a<]�a<̤a<2�a<��a<��a<^�a<��a<�a<u�a<ʧa<.�a<v�a<˨a<"�a<q�a<��a<	�a<P�a<��a<֪a<�a<`�a<��a<ϫa<�a<L�a<w�a<��a<ڬa<�a<:�a<b�a<��a<��a<ҭa<�a<�a<3�a<Z�a<j�a<��a<��a<��a<��a<ծa<�a<�a< �a<�a<�a<�a<�a<�a<�a<�a<�a<�a<��a<�a<�a<�a<Үa<Ʈa<îa<��a<��a<��a<s�a<R�a<8�a<�a<�a<�a<­a<��a<x�a<L�a<+�a<�a<۬a<��a<��a<N�a<�a<�a<��a<��a<Q�a<�a<�a<��a<c�a<#�a<�a<��a<T�a<�a<Ҩa<z�a<3�a<�a<��a<Q�a<�a<��a<S�a<��a<��a<O�a<�a<��a<.�a<ңa<s�a<�a<��a<F�a<�a<r�a<�a<��a<C�a<ޟa<k�a<�a<��a<+�a<��a<L�a<�a<}�a<�a<��a<9�a<ɚa<k�a<��a<��a<+�a<Øa<O�a<��a<��a<4�a<˖a<e�a<�a<��a<W�a<�a<��a<U�a<�a<��a<j�a<�a<ђa<��a<B�a< �a<��a<�a<H�a<�a<ېa<��a<u�a<@�a<�a<��a<Տa<��a<��a<y�a<\�a<G�a<?�a<+�a<�a<�a<�a<��a<��a<�a<�a<�a<�a<,�a<L�a<_�a<j�a<�  �  ��a<��a<ŏa<�a<'�a<<�a<w�a<��a<�a< �a<N�a<��a<��a<�a<*�a<��a<Βa<5�a<m�a<��a< �a<W�a<a<	�a<��a<ӕa<'�a<��a<�a<g�a<��a<6�a<��a<��a<h�a<��a<K�a<��a<=�a<��a<�a<��a<�a<_�a<ĝa<[�a<��a<$�a<��a<�a<��a<�a<|�a<ѡa<H�a<��a<�a<��a<�a<x�a<��a<4�a<��a<�a<R�a<��a<-�a<g�a<ǧa<�a<z�a<Ψa<�a<��a<��a<
�a<<�a<��a<٪a<�a<l�a<��a<ޫa<�a<@�a<n�a<��a<�a<��a<6�a<S�a<��a<��a<ɭa<�a<�a<8�a<5�a<i�a<~�a<��a<��a<��a<ݮa<ήa<�a<�a<�a<�a< �a<�a<�a<%�a<	�a<�a<�a< �a<	�a<خa<�a<֮a<ۮa<îa<��a<��a<s�a<p�a<H�a<E�a<(�a<��a<�a<��a<��a<l�a<\�a<8�a< �a<�a<��a<��a<L�a<6�a<�a<��a<��a<?�a<�a<ͪa<��a<d�a<�a<�a<��a<f�a<�a<٨a<��a<5�a<�a<��a<P�a<�a<��a<C�a<��a<��a<<�a<�a<�a<D�a<ˣa<f�a<�a<��a<N�a<ˡa<��a<
�a<��a<6�a<ǟa<n�a<��a<��a<�a<��a<N�a<ޜa<q�a<�a<��a<*�a<Śa<Y�a<��a<��a<�a<טa<L�a<��a<�a<(�a<ϖa<j�a<#�a<��a<e�a<��a<��a<L�a< �a<œa<U�a<�a<a<��a<=�a<��a<בa<v�a<N�a<��a<ڐa<��a<y�a<T�a<�a<�a<Ïa<��a<��a<}�a<m�a<;�a<<�a<�a<*�a<�a<�a<�a<�a<�a<�a< �a<�a<A�a<L�a<N�a<��a<�  �  ��a<��a<ُa<��a<�a<F�a<|�a<��a<ϐa<�a<L�a<|�a<��a<�a<E�a<��a<͒a<�a<u�a<��a<�a<l�a<Ɣa<�a<q�a<ӕa<;�a<��a<��a<_�a<��a<�a<��a<��a<k�a<�a<H�a<��a< �a<��a<�a<v�a<�a<d�a<֝a<F�a<��a<+�a<��a<�a<��a<��a<m�a<͡a<F�a<��a<$�a<��a<�a<f�a<Ϥa<.�a<��a<�a<W�a<��a<�a<u�a<ѧa<(�a<u�a<ͨa<!�a<j�a<��a<�a<W�a<��a<תa<�a<S�a<��a<֫a<�a<J�a<~�a<��a<ڬa<
�a<8�a<g�a<��a<��a<խa<�a<�a<:�a<N�a<o�a<}�a<��a<��a<îa<Ǯa<�a<��a<��a<��a<�a<�a<�a<�a<�a<�a<�a<�a<�a<��a<�a<�a<ܮa<ɮa<��a<��a<��a<��a<o�a<\�a<5�a<�a< �a<�a<ŭa<��a<~�a<Z�a<'�a<��a<�a<��a<��a<J�a<�a<��a<��a<��a<U�a<�a<ܪa<��a<e�a<-�a<�a<��a<_�a<�a<¨a<��a<7�a<�a<��a<M�a<��a<��a<Q�a<��a<��a<I�a<�a<��a<0�a<ԣa<m�a<�a<��a<B�a<�a<~�a<�a<��a<B�a<ןa<m�a<��a<��a<.�a<��a<N�a<�a<v�a<�a<��a<8�a<Кa<d�a<�a<��a<)�a<��a<Z�a<��a<��a<1�a<͖a<n�a<
�a<��a<]�a<�a<��a<\�a<�a<��a<f�a<�a<גa<��a<?�a<�a<��a<y�a<P�a<�a<��a<��a<o�a<N�a<$�a<��a<Տa<��a<��a<v�a<Y�a<Q�a<<�a<&�a<�a<�a<�a<��a<�a<�a<�a<�a<%�a</�a<>�a<X�a<w�a<�  �  ��a<��a<��a<��a<�a<F�a<g�a<��a<Аa<�a<7�a<��a<̑a<��a<M�a<��a<�a<�a<n�a<��a<�a<�a<��a<�a<p�a<�a<3�a<��a<�a<K�a<֗a<&�a<��a<��a<Y�a<�a<1�a<Ěa<�a<��a<�a<}�a<��a<I�a<�a<B�a<��a<"�a<��a<�a<{�a<��a<S�a<�a<J�a<��a<#�a<��a<�a<P�a<Ѥa<+�a<��a<�a<M�a<��a<�a<��a<��a<)�a<��a<Ȩa<1�a<[�a<ɩa<�a<U�a<��a<Ъa<(�a<Q�a<��a<īa<�a<:�a<r�a<��a<Ԭa<	�a<%�a<t�a<��a<��a<ԭa<�a<#�a<'�a<O�a<c�a<��a<��a<��a<Ȯa<Ǯa<�a<�a<��a<��a<	�a<#�a<��a<!�a<�a<�a<�a<�a<�a<�a<
�a<Ӯa<�a<ʮa<îa<��a<��a<��a<U�a<c�a<>�a<�a<��a<ԭa<׭a<��a<��a<F�a<0�a<�a<լa<��a<w�a<a�a<�a<�a<��a<�a<g�a<�a<۪a<��a<s�a<%�a<ҩa<��a<K�a<)�a<ɨa<��a<4�a<٧a<��a<7�a<�a<��a<`�a<��a<��a<O�a<դa<��a<+�a<ӣa<e�a<�a<��a<<�a<�a<d�a<�a<��a<@�a<֟a<j�a<�a<��a<0�a<��a<U�a<�a<k�a<�a<��a<K�a<��a<f�a<��a<��a<9�a<��a<h�a<�a<��a<%�a<Ɩa<|�a<�a<ȕa<L�a<�a<��a<Q�a<�a<��a<e�a<�a<�a<��a<@�a<�a<��a<��a<<�a<�a<Ԑa<��a<~�a<7�a<)�a<��a<�a<��a<��a<u�a<`�a<^�a<�a<3�a<�a<�a<�a<��a<�a<��a<%�a<�a<0�a<1�a<L�a<j�a<k�a<�  �  ��a<��a<Əa<��a<"�a<P�a<q�a<��a<Րa<	�a<P�a<��a<��a<��a<N�a<��a<ɒa</�a<s�a<��a<�a<_�a<��a<�a<|�a<a<'�a<��a<��a<U�a<��a<)�a<��a<�a<n�a<�a<C�a<��a<�a<��a<��a<|�a<�a<a�a<ŝa<F�a<��a<1�a<��a<�a<}�a<�a<v�a<ڡa<5�a<��a<$�a<��a<��a<s�a<Ǥa<(�a<��a<�a<[�a<��a<�a<g�a<̧a<&�a<|�a<Ĩa<�a<e�a<��a<�a<X�a<��a<ݪa<�a<V�a<��a<ͫa<�a<E�a<p�a<��a<�a<�a<2�a<W�a<��a<��a<ԭa<�a<
�a<&�a<S�a<b�a<m�a<��a<��a<��a<Ȯa<׮a<�a<��a<�a<�a< �a<�a<�a<�a<�a<�a<
�a<�a<��a<�a<�a<�a<Ǯa<��a<��a<��a<��a<p�a<I�a<5�a<#�a<	�a<ޭa<��a<��a<v�a<^�a<8�a<�a<Ԭa<��a<w�a<F�a<0�a<��a<��a<��a<G�a<�a<�a<��a<S�a<�a<�a<��a<U�a<�a<̨a<~�a<<�a<�a<��a<H�a<��a<��a<S�a<�a<��a<K�a<�a<��a<0�a<ԣa<s�a<�a<��a<>�a<١a<��a<�a<��a<?�a<ןa<]�a<�a<��a<%�a<��a<O�a<ܜa<z�a<�a<��a<+�a<˚a<c�a<��a<��a<'�a<��a<W�a<��a<��a<5�a<Ӗa<h�a<�a<��a<U�a<�a<��a<N�a<��a<��a<i�a<�a<ƒa<��a<;�a<�a<ϑa<x�a<;�a<�a<Ӑa<��a<}�a<V�a<�a<�a<̏a<��a<��a<}�a<\�a<;�a<9�a<0�a<�a<�a<�a<�a<�a<�a<�a<�a<,�a<-�a<J�a<S�a<w�a<�  �  ~�a<ɏa<ɏa<��a<�a<>�a<��a<��a<�a<�a<C�a<u�a<��a<�a<D�a<��a<ǒa<�a<l�a<��a<�a<[�a<єa<
�a<|�a<̕a<?�a<��a<�a<f�a<��a<@�a<��a<��a<b�a<řa<H�a<��a<7�a<��a<�a<{�a<ܜa<~�a<Ɲa<W�a<��a<5�a<��a<�a<��a<�a<e�a<ša<P�a<��a<)�a<��a<�a<^�a<��a<8�a<��a<�a<h�a<��a<&�a<f�a<�a<�a<t�a<Ϩa<�a<��a<��a<
�a<=�a<��a<ܪa<�a<r�a<��a<ܫa< �a<K�a<��a<��a<�a<��a<H�a<S�a<��a<��a<˭a<�a<��a<K�a<P�a<t�a<��a<��a<��a<��a<ڮa<ծa<��a<�a< �a<�a<��a</�a<�a<�a<�a< �a<�a< �a<��a<�a<�a<ٮa<Ӯa<Ѯa<��a<��a<q�a<��a<L�a<B�a< �a<��a<�a<��a<��a<r�a<Q�a<!�a<�a<�a<��a<��a<E�a<�a<�a<��a<��a<C�a<)�a<Ϊa<��a<]�a<1�a<�a<��a<f�a< �a<�a<��a<7�a<�a<��a<N�a<��a<��a<R�a<��a<��a<6�a<	�a<��a<A�a<£a<w�a<�a<��a<P�a<֡a<v�a<��a<��a<H�a<ܟa<z�a<�a<��a< �a<ĝa<V�a<ߜa<��a<��a<��a<*�a<�a<V�a<�a<��a<$�a<Ԙa<T�a<��a<��a<#�a<іa<n�a<(�a<��a<c�a<��a<��a<i�a<��a<��a<R�a<+�a<a<��a<<�a<��a<��a<m�a<`�a<�a<�a<��a<f�a<E�a<�a<�a<ʏa<��a<��a<w�a<m�a<9�a<S�a<�a<$�a<�a<�a<�a<�a<�a<��a<�a<!�a<:�a<Z�a<J�a<��a<�  �  ��a<��a<Ϗa<��a<#�a<H�a<k�a<��a<Ԑa<�a<D�a<��a<֑a<�a<0�a<z�a<�a<%�a<|�a<��a<�a<g�a<��a<�a<y�a<ؕa<1�a<��a<��a<g�a<a<!�a<��a<�a<m�a<��a<G�a<��a<�a<��a<�a<��a<�a<^�a<̝a<K�a<��a<7�a<��a<�a<z�a<�a<^�a<�a<H�a<��a<	�a<��a<�a<X�a<פa<*�a<��a<�a<c�a<��a<�a<l�a<̧a<�a<��a<ըa<�a<X�a<��a<	�a<U�a<��a<ߪa<�a<M�a<��a<ܫa<�a<;�a<v�a<��a<߬a<
�a<6�a<\�a<��a<��a<߭a<�a<)�a<"�a<5�a<K�a<��a<��a<��a<Ʈa<ɮa<�a<�a<��a<�a<�a<
�a<�a<�a<&�a<�a<�a<��a<�a<��a<�a<�a<�a<��a<��a<��a<��a<��a<k�a<R�a<A�a<$�a<�a<حa<ŭa<��a<��a<R�a<<�a<�a<��a<��a<o�a<k�a<&�a<��a<��a<��a<P�a<�a<ݪa<��a<i�a<#�a<ݩa<��a<g�a<�a<Ĩa<~�a<=�a<�a<��a<M�a<��a<��a<O�a<��a<��a<<�a<�a<��a<5�a<ԣa<y�a<�a<��a<;�a<�a<o�a<(�a<��a<(�a<��a<c�a<�a<��a<5�a<��a<U�a<ܜa<��a<�a<��a</�a<ʚa<W�a<�a<��a<%�a<��a<\�a<��a<��a<4�a<Ԗa<n�a<�a<��a<d�a<�a<��a<U�a<�a<��a<e�a<�a<̒a<��a<>�a<�a<��a<��a<7�a<��a<��a<��a<��a<B�a<'�a<�a<؏a<��a<��a<~�a<g�a<E�a<4�a<#�a<,�a<�a<�a<��a<�a<	�a<�a<�a</�a<'�a<G�a<[�a<��a<�  �  3�a<\�a<��a<��a<ҏa<��a<!�a<}�a<~�a<Ԑa<�a<&�a<h�a<��a<�a<,�a<��a<��a<?�a<r�a<Гa<7�a<d�a<Ҕa<.�a<��a<�a<H�a<��a<�a<p�a<͗a<W�a<��a<�a<��a<�a<��a<ؚa<O�a<��a<&�a<��a<�a<��a<�a<~�a<�a<d�a<��a<7�a<ՠa<�a<��a<�a<��a<��a<2�a<��a<�a<��a<�a<}�a<ʥa<�a<��a<ݦa<;�a<��a<�a<-�a<{�a<�a<*�a<��a<��a<�a<U�a<��a<��a<�a<^�a<��a<ūa<�a<B�a<l�a<��a<֬a<�a<?�a<^�a<n�a<��a<��a<ܭa<�a<(�a<4�a<3�a<P�a<x�a<��a<��a<Ȯa<��a<��a<ʮa<Ǯa<߮a<ծa<ͮa<ͮa<̮a<Үa<ˮa<�a<��a<Юa<��a<��a<��a<x�a<f�a<O�a<:�a<-�a<$�a<��a<�a<ía<��a<��a<W�a<S�a<,�a<�a<��a<��a<��a<3�a<�a<ʫa<ѫa<��a<U�a<0�a<ͪa<��a<j�a<!�a<�a<��a<T�a<�a<Ѩa<~�a<S�a<��a<��a<h�a<��a<ۦa<b�a<�a<��a<T�a<�a<��a<[�a<�a<��a<(�a<Ԣa<��a<��a<��a<-�a<Ϡa<I�a<�a<��a<�a<��a<?�a<�a<n�a<2�a<��a<*�a<ћa<^�a<��a<��a<�a<��a<0�a<�a<o�a<-�a<��a<P�a<��a<�a<:�a<��a<k�a<��a<��a<[�a<�a<��a<l�a< �a<��a<��a<K�a<�a<ёa<V�a<7�a<�a<֐a<��a<E�a<�a<�a<�a<��a<��a<c�a<?�a<-�a<	�a<�a<�a<ˎa<��a<��a<��a<��a<ӎa<��a<׎a<��a<�a<�a<�a<�a<�a<�  �  I�a<^�a<y�a<��a<ˏa<�a<%�a<E�a<}�a<��a<��a<:�a<��a<��a<�a<<�a<��a<Ԓa<#�a<[�a<ēa<	�a<x�a<ϔa<+�a<��a<�a<H�a<��a<!�a<v�a<�a<G�a<��a<!�a<��a<��a<o�a<�a<Z�a<ța<P�a<��a<�a<��a<�a<r�a<�a<O�a<ɟa<.�a<��a< �a<��a<�a<k�a<բa<T�a<Σa<�a<��a<ܤa<R�a<��a<'�a<y�a<�a<3�a<��a<�a<Y�a<��a<�a<:�a<�a<ĩa<�a<\�a<��a<ުa<-�a<^�a<��a<�a<�a<>�a<r�a<��a<Ϭa<�a<�a<J�a<[�a<��a<��a<�a<��a<�a<*�a<R�a<g�a<j�a<}�a<��a<��a<��a<Ʈa<®a<ծa<̮a<֮a<ޮa<�a<خa<�a<ɮa<ήa<��a<��a<��a<��a<��a<��a<o�a<n�a<P�a</�a<�a<�a<�a<ͭa<��a<s�a<V�a<4�a<�a<��a<٬a<��a<c�a<C�a<+�a<�a<��a<h�a<H�a<�a<�a<��a<g�a<*�a<�a<��a<r�a</�a<֨a<��a<C�a<��a<��a<c�a<�a<��a<j�a<�a<¥a<�a<�a<��a<K�a<��a<��a<:�a<��a<c�a<�a<��a<2�a<�a<o�a<��a<��a<.�a<ўa<M�a<�a<b�a<�a<��a<=�a<ěa<d�a<�a<��a<"�a<˙a<P�a<�a<�a<�a<��a<O�a<�a<��a<#�a<ӕa<j�a<�a<˔a<c�a<�a<��a<n�a<�a<Ԓa<r�a<7�a<ܑa<��a<q�a<I�a<��a<��a<��a<e�a<3�a<�a<ʏa<��a<r�a<_�a<N�a<%�a<�a<�a<�a<܎a<ݎa<��a<̎a<��a<��a<��a<Ďa<a<׎a<ގa<�a<�a<6�a<�  �  2�a<e�a<}�a<��a<��a<��a<2�a<T�a<��a<��a<��a<-�a<k�a<��a<��a<I�a<y�a<Ԓa<"�a<u�a<�a<�a<��a<��a<�a<��a<�a<C�a<��a<�a<h�a<��a<7�a<��a<+�a<��a<�a<`�a<�a<P�a<��a</�a<��a<%�a<��a<�a<^�a<��a<[�a<ߟa<\�a<��a<*�a<��a<�a<}�a<�a<Y�a<��a<*�a<��a<�a<n�a<��a<-�a<f�a<�a<7�a<��a<ߧa<6�a<��a<ܨa<@�a<q�a<ܩa<�a<_�a<��a<ͪa<6�a<N�a<��a<ūa<�a<D�a<t�a<��a<��a<�a<�a<s�a<{�a<��a<��a<ǭa<�a<�a<9�a<?�a<P�a<s�a<��a<��a<��a<��a<��a<��a<�a<Ϯa<�a<Ȯa<׮a<ͮa<�a<ɮa<Ǯa<ծa<��a<��a<��a<��a<��a<`�a<[�a<8�a<6�a<�a<�a<ʭa<ía<��a<��a<��a<=�a<�a<�a<��a<��a<x�a<Q�a<�a<�a<��a<��a<r�a<�a<�a<��a<[�a<.�a<�a<��a<T�a<�a<ɨa<��a<3�a<�a<��a<\�a<!�a<��a<n�a<�a<��a<^�a<��a<��a<N�a<�a<y�a<>�a<ˢa<y�a<�a<��a<<�a<��a<l�a<�a<��a<2�a<��a<W�a<�a<��a<#�a<��a<D�a<��a<i�a<�a<��a<�a<��a<>�a<טa<��a<�a<��a<H�a<�a<��a<�a<ݕa<[�a<�a<��a<Y�a<�a<��a<g�a<�a<�a<w�a<`�a<��a<��a<w�a<"�a<�a<Ða<��a<R�a<�a<��a<Џa<͏a<��a<l�a<G�a<�a<#�a<��a<��a<Ǝa<Ȏa<��a<Ȏa<��a<��a<̎a<��a<َa<׎a<؎a<�a<��a<$�a<�  �  E�a<b�a<��a<��a<Ϗa< �a<�a<k�a<s�a<��a<�a<3�a<w�a<��a<��a<6�a<��a<Вa<*�a<d�a<��a<#�a<g�a<הa<1�a<��a<�a<L�a<��a<!�a<��a<җa<A�a<��a< �a<��a<��a<{�a<ۚa<P�a<ԛa<D�a<��a<�a<��a<�a<{�a<�a<T�a<џa<'�a<��a<0�a<��a<�a<t�a<�a<L�a<��a<)�a<��a<٤a<T�a<��a<�a<��a<�a<4�a<��a<��a<M�a<��a<�a<.�a<��a<ɩa<�a<Z�a<��a<ܪa<�a<i�a<��a<ޫa<�a<=�a<m�a<��a<ܬa<��a<%�a<B�a<_�a<��a<��a<�a<�a<�a<*�a<G�a<_�a<�a<|�a<z�a<��a<��a<��a<Įa<ʮa<Ѯa<خa<�a<�a<�a<ɮa<Ϯa<Ԯa<��a<Юa<��a<��a<��a<s�a<��a<j�a<K�a<2�a<�a<��a<�a<̭a<��a<��a<L�a<5�a<)�a<�a<ͬa<��a<p�a<=�a<!�a<�a<��a<q�a<;�a<�a<Ϫa<��a<m�a<#�a<�a<��a<i�a<.�a<�a<��a<>�a< �a<��a<g�a<�a<ɦa<e�a<�a<Υa<s�a<�a<��a<M�a<�a<��a<3�a<Ģa<k�a<�a<��a<B�a<֠a<f�a<��a<��a<%�a<Þa<W�a<�a<_�a<	�a<��a<3�a<ћa<a�a<�a<��a<)�a<��a<Z�a<�a<s�a<�a<��a<M�a<�a<��a< �a<��a<v�a<#�a<Ôa<i�a<
�a<��a<q�a<%�a<ƒa<��a</�a<�a<��a<p�a<=�a<�a<��a<��a<Y�a<+�a<	�a<ɏa<��a<��a<V�a<I�a<'�a<�a<��a<�a<ގa<؎a<ӎa<��a<��a<��a<��a<׎a<��a<ގa<�a<�a<�a<3�a<�  �  G�a<W�a<��a<��a<Ϗa<�a<�a<m�a<{�a<ېa<�a<,�a<��a<��a<��a<3�a<��a<��a<#�a<��a<��a<1�a<_�a<ݔa<�a<��a<�a<B�a<��a<��a<~�a<ٗa<^�a<��a<�a<��a<�a<��a<ޚa<O�a<��a<!�a<��a<�a<��a<��a<��a<�a<]�a<۟a<F�a<Ҡa<�a<��a<�a<n�a<�a<H�a<̣a<�a<��a<��a<_�a<åa<�a<��a<Цa<K�a<��a<�a</�a<��a<�a<0�a<��a<��a<�a<X�a<��a<��a<�a<e�a<��a<̫a<�a<@�a<{�a<��a<�a<�a<7�a<G�a<��a<��a<��a<��a<�a<�a<$�a<P�a<[�a<[�a<��a<��a<��a<��a<Ǯa<ɮa<Ʈa<�a<̮a<�a<��a<ޮa<Юa<ڮa<׮a<��a<Ȯa<��a<��a<��a<~�a<w�a<D�a<M�a<(�a<'�a<��a<�a<ԭa<��a<��a<T�a<Z�a<
�a<�a<ݬa<��a<z�a<:�a<4�a<Ыa<��a<��a<?�a<)�a<Ǫa<��a<Y�a<,�a<�a<��a<c�a<	�a<ߨa<��a<[�a<��a<��a<h�a<�a<Ӧa<h�a<�a<��a<P�a<�a<��a<i�a<�a<��a<2�a<΢a<u�a<�a<��a<�a<ݠa<d�a<��a<��a<!�a<Ϟa<6�a<��a<��a<�a<��a<.�a<՛a<P�a<�a<z�a<�a<��a<6�a<�a<u�a<*�a<��a<O�a<�a<{�a<=�a<��a<q�a<��a<��a<]�a<�a<Óa<Y�a<)�a<��a<��a<4�a<�a<��a<W�a<Q�a<�a<ɐa<��a<c�a<'�a<�a<�a<��a<��a<Q�a<P�a<,�a<	�a<�a<ݎa<ߎa<��a<Ǝa<��a<��a<Îa<��a<ώa<��a<ێa<�a<�a<�a<�a<�  �  E�a<c�a<|�a<��a<ďa<��a<6�a<D�a<��a<Őa<�a<@�a<f�a<��a<�a<:�a<w�a<ܒa<�a<y�a<Ɠa<�a<��a<ؔa<�a<��a<�a<K�a<��a<�a<x�a<�a<;�a<��a</�a<��a<�a<c�a<ךa<V�a<ϛa<3�a<��a<�a<��a<��a<v�a<��a<`�a<ßa<I�a<��a<%�a<��a<��a<�a<�a<I�a<��a<(�a<��a<��a<M�a<��a<)�a<��a<զa<5�a<��a<�a<>�a<��a<�a<-�a<q�a<۩a<�a<b�a<��a<Ѫa< �a<d�a<��a<Ыa<�a<=�a<p�a<��a<۬a<�a<�a<G�a<{�a<��a<��a<˭a<�a<!�a<0�a<9�a<b�a<j�a<��a<��a<��a<��a<îa<��a<Ѯa<ˮa<خa<�a<ڮa<�a<ۮa<Įa<ʮa<ٮa<��a<Ʈa<��a<��a<��a<v�a<`�a<K�a<4�a<�a<�a<حa<̭a<��a<s�a<f�a<D�a<�a<��a<��a<��a<��a<A�a<�a<�a<��a<��a<K�a<�a<�a<��a<W�a<&�a<�a<��a<c�a<&�a<بa<��a<7�a<��a<��a<Y�a<"�a<��a<a�a<�a<ɥa<b�a<�a<��a<N�a<�a<��a<<�a<Тa<\�a<�a<��a<7�a<Ϡa<^�a<�a<��a<#�a<��a<U�a<�a<��a<�a<��a<?�a<̛a<U�a<�a<��a<�a<��a<S�a<�a<r�a<�a<��a<D�a<�a<��a<�a<ƕa<p�a<�a<��a<c�a<
�a<��a<\�a<%�a<ؒa<x�a<4�a<��a<��a<w�a<&�a<��a<ΐa<��a<K�a<.�a<�a<֏a<��a<s�a<o�a<K�a<!�a<�a<�a<�a<ߎa<ˎa<Ɏa<��a<��a<��a<Ўa<��a<�a<֎a<Ԏa<��a<�a<)�a<�  �  ,�a<u�a<p�a<��a<Տa<�a<<�a<A�a<��a<��a<�a<?�a<m�a<ʑa<֑a<Y�a<{�a<�a<�a<h�a<ٓa<�a<��a<��a<6�a<��a<ޕa<Y�a<��a<#�a<b�a<��a<L�a<��a<(�a<r�a<�a<`�a<��a<C�a<ƛa<@�a<��a<+�a<��a<�a<p�a<�a<g�a<̟a<Q�a<��a<>�a<��a<�a<q�a<Ӣa<i�a<��a<>�a<y�a<��a<[�a<��a<*�a<t�a<�a<,�a<��a<�a<E�a<��a<Ѩa<N�a<s�a<�a<��a<Z�a<��a<ܪa<7�a<G�a<��a<ɫa<�a<?�a<l�a<��a<��a<�a<�a<Z�a<s�a<��a<ҭa<˭a<�a<�a<9�a<H�a<a�a<��a<n�a<��a<��a<Ůa<��a<Ǯa<ڮa<��a<�a<ʮa<�a<ʮa<Ӯa<�a<��a<ݮa<��a<Ůa<��a<��a<��a<_�a<r�a<2�a<F�a<�a<�a<�a<��a<��a<p�a<x�a<-�a<%�a<��a<ìa<��a<Q�a<`�a<	�a<��a<��a<u�a<^�a<�a<�a<��a<r�a<'�a<ߩa<��a<S�a<1�a<èa<��a<I�a<�a<��a<A�a<-�a<��a<��a<�a<��a<n�a<�a<��a<D�a<��a<��a<6�a<עa<e�a<�a<��a<P�a<Ƞa<y�a<��a<��a<B�a<��a<k�a<ҝa<��a<�a<��a<A�a<��a<h�a<�a<��a<�a<��a<Q�a<̘a<��a<�a<ȗa<3�a<�a<��a< �a<ޕa<T�a<�a<��a<l�a<�a<��a<u�a<
�a<ܒa<z�a<G�a<��a<��a<��a<&�a<�a<��a<��a<Z�a<-�a<�a<��a<��a<s�a<w�a<7�a<+�a<�a<�a<��a<Ȏa<��a<��a<��a<̎a<��a<Ԏa<��a<�a<̎a<�a<��a<��a<;�a<�  �  0�a<p�a<��a<��a<ҏa<�a<*�a<X�a<��a<Đa<�a<#�a<r�a<ˑa<�a<U�a<��a<ɒa<'�a<|�a<ēa<#�a<u�a<Ŕa<)�a<��a<�a<Q�a<��a<�a<{�a<ٗa<L�a<��a<&�a<��a<��a<c�a<�a<L�a<˛a<-�a<��a<(�a<��a<��a<v�a<�a<b�a<Пa<N�a<��a<%�a<��a<�a<z�a<�a<^�a<��a< �a<��a<��a<X�a<��a<�a<|�a<Ԧa<>�a<��a<�a<4�a<��a<ߨa<7�a<y�a<ũa<�a<c�a<��a<ߪa<�a<^�a<��a<ëa<�a<H�a<n�a<��a<ʬa<��a<-�a<J�a<�a<��a<��a<ѭa<�a<�a<?�a<F�a<K�a<v�a<��a<��a<��a<��a<��a<Ǯa<��a<ܮa<�a<ɮa<ۮa<߮a<Ϯa<ۮa<��a<��a<ɮa<��a<��a<��a<y�a<v�a<_�a<6�a<A�a<�a<�a<�a<��a<��a<��a<g�a<C�a<!�a<�a<ɬa<��a<i�a<\�a<�a<۫a<��a<��a<I�a<�a<ݪa<��a<e�a<!�a<�a<��a<R�a<$�a<ܨa<��a<I�a<�a<��a<k�a<�a<��a<l�a<�a<ťa<[�a<�a<��a<]�a<�a<��a<2�a<Ңa<i�a<�a<��a<7�a<��a<r�a<�a<��a<7�a<��a<M�a<�a<��a<�a<��a<6�a<ƛa<T�a<��a<��a<�a<��a<N�a<ۘa<|�a<
�a<��a<S�a<�a<z�a<$�a<Õa<k�a<�a<��a<c�a<�a<��a<c�a<�a<ϒa<��a<7�a<�a<��a<j�a<,�a<�a<��a<��a<Y�a<�a< �a<Џa<��a<��a<f�a<@�a<*�a<�a<�a<��a<ǎa<̎a<ǎa<��a<��a<��a<��a<Ўa<Ɏa<Ȏa<�a<�a<�a<(�a<�  �  Y�a<J�a<��a<��a<ʏa<�a<�a<[�a<r�a<ǐa<��a<E�a<u�a<��a<�a<�a<��a<ڒa<�a<v�a<��a<#�a<h�a<�a<!�a<��a<�a<9�a<��a<�a<��a<ȗa<M�a<��a<�a<��a<��a<��a<��a<^�a<՛a<2�a<��a<�a<��a<��a<��a<�a<]�a<ȟa<0�a<��a<!�a<��a<��a<v�a<�a<<�a<ԣa<!�a<��a<�a<L�a<��a<�a<��a<Ϧa<F�a<��a<��a<B�a<��a<��a<�a<��a<éa<�a<R�a<��a<�a<�a<z�a<��a<߫a<�a<B�a<x�a<��a<�a<�a<,�a<7�a<n�a<��a<��a<�a<حa<�a<�a<B�a<o�a<i�a<��a<�a<��a<��a<Ʈa<Ǯa<Įa<�a<®a<�a<̮a<�a<Үa<��a<�a<��a<��a<��a<��a<��a<v�a<��a<N�a<`�a<�a<)�a<��a<ޭa<ӭa<��a<��a<K�a<E�a<�a<�a<ˬa<��a<��a<%�a<&�a<�a<��a<��a<1�a<�a<Ъa<��a<\�a<+�a<�a<��a<t�a<�a<�a<x�a<I�a<�a<��a<e�a<�a<ئa<K�a<!�a<ϥa<`�a<�a<��a<b�a<�a<��a<0�a<͢a<b�a<�a<��a<3�a<�a<\�a<��a<��a<�a<מa<O�a<�a<f�a< �a<��a<+�a<ڛa<O�a< �a<|�a<%�a<��a<T�a<�a<Z�a<%�a<��a<I�a<ݖa<��a</�a<��a<��a<�a<Ĕa<[�a<�a<��a<\�a<0�a<��a<��a<$�a<�a<��a<t�a<H�a<ڐa<ːa<z�a<U�a<;�a<�a<؏a<��a<��a<[�a<N�a<*�a<�a<�a<Ҏa<�a<��a<؎a<��a<��a<Ԏa<��a<Ǝa<��a<�a<َa<�a<(�a<�a<�  �  S�a<O�a<��a<��a<ʏa<��a<'�a<Z�a<��a<ϐa<�a<1�a<{�a<��a<�a<7�a<��a<ђa<�a<��a<ӓa<$�a<s�a<˔a<&�a<��a<�a<<�a<��a<��a<r�a<�a<P�a<��a<�a<��a<��a<v�a<ݚa<S�a<��a<+�a<��a<�a<��a<�a<t�a<�a<i�a<ޟa<W�a<��a<!�a<��a<�a<v�a<�a<O�a<£a< �a<��a<�a<g�a<ɥa<�a<|�a<�a<C�a<��a<�a<8�a<z�a<�a<6�a<��a<ǩa<�a<X�a<��a<�a<+�a<[�a<}�a<֫a<��a<B�a<r�a<��a<ͬa<��a<1�a<\�a<��a<��a<��a<�a<�a<�a<+�a<M�a<T�a<a�a<��a<��a<��a<��a<��a<��a<Ӯa<ݮa<ɮa<�a<Ȯa<̮a<�a<ͮa<Ԯa<��a<��a<��a<��a<��a<��a<f�a<G�a<Y�a< �a<!�a< �a<ޭa<ƭa<��a<��a<p�a<N�a<
�a<�a<Ҭa<��a<��a<>�a<!�a<�a<��a<��a<X�a<�a<۪a<��a<b�a<&�a<�a<��a<p�a<�a<Өa<��a<L�a<��a<��a<[�a<�a<Ŧa<g�a<�a<��a<Z�a<�a<��a<^�a<��a<��a<0�a<٢a<w�a<�a<��a<2�a<Ϡa<h�a<��a<��a<)�a<Şa<M�a<�a<��a<�a<��a<1�a<ƛa<b�a<��a<��a<�a<��a</�a<��a<z�a<�a<��a<F�a<�a<��a<+�a<ҕa<h�a<��a<��a<U�a<�a<��a<f�a<�a<ʒa<��a<I�a<�a<��a<o�a<@�a<��a<̐a<��a<_�a< �a<�a<�a<��a<��a<f�a<F�a<%�a<�a<�a<َa<�a<��a<��a<Ŏa<��a<��a<��a<��a<Îa<ێa<�a<�a<�a<�a<�  �  <�a<m�a<|�a<��a<ݏa<��a<)�a<G�a<��a<��a<	�a<'�a<w�a<Ña<��a<R�a<��a<Βa<,�a<g�a<��a<	�a<|�a<ɔa<<�a<k�a<�a<N�a<��a<3�a<v�a<�a<<�a<��a<,�a<��a<�a<[�a<�a<T�a<Λa<X�a<��a</�a<z�a<�a<y�a<�a<W�a<ğa<=�a<��a<<�a<��a<�a<y�a<�a<a�a<��a<5�a<��a<�a<N�a<��a<'�a<~�a<�a< �a<��a<�a<X�a<��a<�a<:�a<m�a<֩a<�a<b�a<��a<Ϊa<#�a<\�a<��a<ݫa<�a<I�a<X�a<��a<̬a<�a<�a<H�a<g�a<��a<��a<έa<
�a<�a<:�a<L�a<J�a<��a<t�a<��a<��a<��a<��a<ήa<��a<Ǯa<�a<Ϯa< �a<خa<׮a<Ϯa<��a<Ϯa<��a<��a<��a<��a<��a<o�a<��a<B�a<>�a<�a<�a<�a<��a<��a<v�a<a�a</�a<*�a<�a<ͬa<��a<q�a<Y�a<�a<�a<��a<u�a<F�a<�a<�a<��a<x�a<�a<�a<��a<i�a<@�a<רa<��a<9�a<��a<��a<`�a<�a<��a<o�a<�a<ȥa<��a< �a<��a<;�a<��a<��a<:�a<Ȣa<^�a<��a<��a<N�a<��a<v�a<�a<��a<:�a<��a<b�a<ܝa<q�a<�a<��a<>�a<ɛa<f�a<ٚa<��a<�a<ʙa<Y�a<�a<~�a<��a<��a<K�a<�a<��a<�a<ɕa<i�a<,�a<��a<^�a<�a<��a<{�a<�a<֒a<s�a<5�a<�a<��a<t�a<)�a<�a<��a<��a<_�a<�a<�a<��a<��a<s�a<_�a<C�a<1�a<�a<�a<��a<͎a<�a<��a<��a<��a<��a<Ǝa<Ŏa<׎a<͎a<ߎa<��a<�a<K�a<�  �  /�a<`�a<��a<��a<ԏa<��a<$�a<`�a<��a<��a<�a</�a<s�a<��a<��a<8�a<��a<͒a<2�a<s�a<ړa<�a<q�a<ǔa<2�a<��a<�a<B�a<��a<�a<s�a<ڗa<W�a<��a<�a<��a< �a<��a<ޚa<R�a<��a<1�a<��a<$�a<��a<�a<x�a<�a<c�a<�a<P�a<��a<1�a<��a<�a<y�a<�a<I�a<��a<,�a<��a<��a<r�a<ĥa<�a<{�a<�a<4�a<��a<ܧa<8�a<{�a<�a</�a<��a<ϩa<�a<S�a<��a<�a<�a<Z�a<��a<ȫa<��a<H�a<l�a<��a<ɬa<��a<-�a<g�a<x�a<��a<��a<ۭa<�a<�a<+�a<C�a<X�a<��a<��a<��a<��a<��a<��a<ɮa<ͮa<׮a<ٮa<Ʈa<׮a<®a<ծa<Ӯa<ޮa<��a<��a<��a<��a<��a<~�a<b�a<S�a<6�a<1�a<�a<��a<�a<��a<��a<��a<u�a<=�a<,�a<�a<ʬa<��a<v�a<?�a<�a<߫a<īa<��a<_�a<�a<٪a<��a<n�a<#�a<�a<��a<S�a<�a<Өa<��a<T�a<�a<��a<P�a<�a<Ѧa<g�a<�a<��a<`�a<��a<��a<P�a<��a<��a<1�a<Ӣa<��a<�a<��a<C�a<Πa<c�a<�a<��a<#�a<��a<Z�a<�a<��a<&�a<��a<4�a<ƛa<d�a<�a<��a<�a<��a<0�a<�a<s�a<%�a<��a<:�a<ޖa<��a<7�a<��a<g�a<��a<��a<S�a<�a<��a<q�a<�a<Ȓa<��a<T�a<��a<��a<q�a<6�a<�a<Ða<��a<U�a<$�a<�a<Ώa<��a<��a<a�a<=�a<,�a<�a<��a<�a<Ďa<Ȏa<��a<��a<��a<ˎa<��a<��a<Ǝa<�a<�a<�a<��a<�a<�  �  f�a<X�a<��a<��a<ʏa<�a<"�a<G�a<|�a<��a<�a<6�a<��a<��a<
�a<)�a<��a<̒a< �a<d�a<��a<�a<q�a<ڔa<#�a<��a<�a<J�a<Җa<�a<��a<�a<A�a<��a<,�a<��a<�a<p�a<Ěa<n�a<��a<I�a<��a<�a<��a<�a<u�a<�a<V�a<ßa<2�a<��a<�a<��a<��a<u�a<�a<@�a<֣a<�a<��a<ޤa<G�a<��a<�a<�a<ݦa<A�a<��a<��a<]�a<��a<�a<�a<��a<��a<(�a<i�a<��a<ݪa<�a<}�a<��a<��a<�a<6�a<u�a<��a<۬a<��a<�a<>�a<`�a<��a<��a<��a<�a<�a<#�a<O�a<c�a<_�a<z�a<��a<��a<��a<Įa<��a<Ѯa<֮a<ʮa<��a<߮a<ܮa<�a<��a<Ȯa<��a<ˮa<��a<��a<��a<��a<��a<V�a<l�a<(�a<�a<�a<ޭa<Эa<��a<v�a<U�a<4�a<�a<��a<ܬa<��a<��a<0�a<5�a<߫a<��a<q�a<>�a<	�a<٪a<��a<_�a<+�a<�a<��a<��a<�a<��a<��a<=�a<�a<��a<u�a<��a<��a<N�a<1�a<��a<x�a<!�a<��a<Z�a<��a<��a<2�a<Ǣa<\�a<��a<��a<-�a<�a<_�a<��a<��a<�a<ٞa<I�a<�a<d�a<��a<��a<1�a<ʛa<^�a<��a<|�a<-�a<ϙa<=�a<��a<b�a<�a<��a<\�a<��a<h�a<"�a<��a<��a<�a<�a<c�a<�a<��a<e�a<$�a<ɒa<z�a<+�a<�a<��a<l�a<T�a<�a<̐a<��a<b�a</�a<�a<Ǐa<��a<u�a<a�a<M�a<$�a<�a<��a<ڎa<��a<Ўa<Ďa<֎a<��a<��a<��a<Ҏa<��a<Ύa<ӎa<�a<�a<�a<�  �  /�a<`�a<��a<��a<ԏa<��a<$�a<`�a<��a<��a<�a</�a<s�a<��a<��a<8�a<��a<͒a<2�a<s�a<ړa<�a<q�a<ǔa<2�a<��a<�a<B�a<��a<�a<s�a<ڗa<W�a<��a<�a<��a< �a<��a<ޚa<R�a<��a<1�a<��a<$�a<��a<�a<x�a<�a<c�a<�a<P�a<��a<1�a<��a<�a<y�a<�a<I�a<��a<,�a<��a<��a<r�a<ĥa<�a<{�a<�a<4�a<��a<ܧa<8�a<{�a<�a</�a<��a<ϩa<�a<S�a<��a<�a<�a<Z�a<��a<ȫa<��a<H�a<l�a<��a<ɬa<��a<-�a<g�a<x�a<��a<��a<ۭa<�a<�a<+�a<C�a<X�a<��a<��a<��a<��a<��a<��a<ɮa<ͮa<׮a<ٮa<Ʈa<׮a<®a<ծa<Ӯa<ޮa<��a<��a<��a<��a<��a<~�a<b�a<S�a<6�a<1�a<�a<��a<�a<��a<��a<��a<u�a<=�a<,�a<�a<ʬa<��a<v�a<?�a<�a<߫a<īa<��a<_�a<�a<٪a<��a<n�a<#�a<�a<��a<S�a<�a<Өa<��a<T�a<�a<��a<P�a<�a<Ѧa<g�a<�a<��a<`�a<��a<��a<P�a<��a<��a<1�a<Ӣa<��a<�a<��a<C�a<Πa<c�a<�a<��a<#�a<��a<Z�a<�a<��a<&�a<��a<4�a<ƛa<d�a<�a<��a<�a<��a<0�a<�a<s�a<%�a<��a<:�a<ޖa<��a<7�a<��a<g�a<��a<��a<S�a<�a<��a<q�a<�a<Ȓa<��a<T�a<��a<��a<q�a<6�a<�a<Ða<��a<U�a<$�a<�a<Ώa<��a<��a<a�a<=�a<,�a<�a<��a<�a<Ďa<Ȏa<��a<��a<��a<ˎa<��a<��a<Ǝa<�a<�a<�a<��a<�a<�  �  <�a<m�a<|�a<��a<ݏa<��a<)�a<G�a<��a<��a<	�a<'�a<w�a<Ña<��a<R�a<��a<Βa<,�a<g�a<��a<	�a<|�a<ɔa<<�a<k�a<�a<N�a<��a<3�a<v�a<�a<<�a<��a<,�a<��a<�a<[�a<�a<T�a<Λa<X�a<��a</�a<z�a<�a<y�a<�a<W�a<ğa<=�a<��a<<�a<��a<�a<y�a<�a<a�a<��a<5�a<��a<�a<N�a<��a<'�a<~�a<�a< �a<��a<�a<X�a<��a<�a<:�a<m�a<֩a<�a<b�a<��a<Ϊa<#�a<\�a<��a<ݫa<�a<I�a<X�a<��a<̬a<�a<�a<H�a<g�a<��a<��a<έa<
�a<�a<:�a<L�a<J�a<��a<t�a<��a<��a<��a<��a<ήa<��a<Ǯa<�a<Ϯa< �a<خa<׮a<Ϯa<��a<Ϯa<��a<��a<��a<��a<��a<o�a<��a<B�a<>�a<�a<�a<�a<��a<��a<v�a<a�a</�a<*�a<�a<ͬa<��a<q�a<Y�a<�a<�a<��a<u�a<F�a<�a<�a<��a<x�a<�a<�a<��a<i�a<@�a<רa<��a<9�a<��a<��a<`�a<�a<��a<o�a<�a<ȥa<��a< �a<��a<;�a<��a<��a<:�a<Ȣa<^�a<��a<��a<N�a<��a<v�a<�a<��a<:�a<��a<b�a<ܝa<q�a<�a<��a<>�a<ɛa<f�a<ٚa<��a<�a<ʙa<Y�a<�a<~�a<��a<��a<K�a<�a<��a<�a<ɕa<i�a<,�a<��a<^�a<�a<��a<{�a<�a<֒a<s�a<5�a<�a<��a<t�a<)�a<�a<��a<��a<_�a<�a<�a<��a<��a<s�a<_�a<C�a<1�a<�a<�a<��a<͎a<�a<��a<��a<��a<��a<Ǝa<Ŏa<׎a<͎a<ߎa<��a<�a<K�a<�  �  S�a<O�a<��a<��a<ʏa<��a<'�a<Z�a<��a<ϐa<�a<1�a<{�a<��a<�a<7�a<��a<ђa<�a<��a<ӓa<$�a<s�a<˔a<&�a<��a<�a<<�a<��a<��a<r�a<�a<P�a<��a<�a<��a<��a<v�a<ݚa<S�a<��a<+�a<��a<�a<��a<�a<t�a<�a<i�a<ޟa<W�a<��a<!�a<��a<�a<v�a<�a<O�a<£a< �a<��a<�a<g�a<ɥa<�a<|�a<�a<C�a<��a<�a<8�a<z�a<�a<6�a<��a<ǩa<�a<X�a<��a<�a<+�a<[�a<}�a<֫a<��a<B�a<r�a<��a<ͬa<��a<1�a<\�a<��a<��a<��a<�a<�a<�a<+�a<M�a<T�a<a�a<��a<��a<��a<��a<��a<��a<Ӯa<ݮa<ɮa<�a<Ȯa<̮a<�a<ͮa<Ԯa<��a<��a<��a<��a<��a<��a<f�a<G�a<Y�a< �a<!�a< �a<ޭa<ƭa<��a<��a<p�a<N�a<
�a<�a<Ҭa<��a<��a<>�a<!�a<�a<��a<��a<X�a<�a<۪a<��a<b�a<&�a<�a<��a<p�a<�a<Өa<��a<L�a<��a<��a<[�a<�a<Ŧa<g�a<�a<��a<Z�a<�a<��a<^�a<��a<��a<0�a<٢a<w�a<�a<��a<2�a<Ϡa<h�a<��a<��a<)�a<Şa<M�a<�a<��a<�a<��a<1�a<ƛa<b�a<��a<��a<�a<��a</�a<��a<z�a<�a<��a<F�a<�a<��a<+�a<ҕa<h�a<��a<��a<U�a<�a<��a<f�a<�a<ʒa<��a<I�a<�a<��a<o�a<@�a<��a<̐a<��a<_�a< �a<�a<�a<��a<��a<f�a<F�a<%�a<�a<�a<َa<�a<��a<��a<Ŏa<��a<��a<��a<��a<Îa<ێa<�a<�a<�a<�a<�  �  Y�a<J�a<��a<��a<ʏa<�a<�a<[�a<r�a<ǐa<��a<E�a<u�a<��a<�a<�a<��a<ڒa<�a<v�a<��a<#�a<h�a<�a<!�a<��a<�a<9�a<��a<�a<��a<ȗa<M�a<��a<�a<��a<��a<��a<��a<^�a<՛a<2�a<��a<�a<��a<��a<��a<�a<]�a<ȟa<0�a<��a<!�a<��a<��a<v�a<�a<<�a<ԣa<!�a<��a<�a<L�a<��a<�a<��a<Ϧa<F�a<��a<��a<B�a<��a<��a<�a<��a<éa<�a<R�a<��a<�a<�a<z�a<��a<߫a<�a<B�a<x�a<��a<�a<�a<,�a<7�a<n�a<��a<��a<�a<حa<�a<�a<B�a<o�a<i�a<��a<�a<��a<��a<Ʈa<Ǯa<Įa<�a<®a<�a<̮a<�a<Үa<��a<�a<��a<��a<��a<��a<��a<v�a<��a<N�a<`�a<�a<)�a<��a<ޭa<ӭa<��a<��a<K�a<E�a<�a<�a<ˬa<��a<��a<%�a<&�a<�a<��a<��a<1�a<�a<Ъa<��a<\�a<+�a<�a<��a<t�a<�a<�a<x�a<I�a<�a<��a<e�a<�a<ئa<K�a<!�a<ϥa<`�a<�a<��a<b�a<�a<��a<0�a<͢a<b�a<�a<��a<3�a<�a<\�a<��a<��a<�a<מa<O�a<�a<f�a< �a<��a<+�a<ڛa<O�a< �a<|�a<%�a<��a<T�a<�a<Z�a<%�a<��a<I�a<ݖa<��a</�a<��a<��a<�a<Ĕa<[�a<�a<��a<\�a<0�a<��a<��a<$�a<�a<��a<t�a<H�a<ڐa<ːa<z�a<U�a<;�a<�a<؏a<��a<��a<[�a<N�a<*�a<�a<�a<Ҏa<�a<��a<؎a<��a<��a<Ԏa<��a<Ǝa<��a<�a<َa<�a<(�a<�a<�  �  0�a<p�a<��a<��a<ҏa<�a<*�a<X�a<��a<Đa<�a<#�a<r�a<ˑa<�a<U�a<��a<ɒa<'�a<|�a<ēa<#�a<u�a<Ŕa<)�a<��a<�a<Q�a<��a<�a<{�a<ٗa<L�a<��a<&�a<��a<��a<c�a<�a<L�a<˛a<-�a<��a<(�a<��a<��a<v�a<�a<b�a<Пa<N�a<��a<%�a<��a<�a<z�a<�a<^�a<��a< �a<��a<��a<X�a<��a<�a<|�a<Ԧa<>�a<��a<�a<4�a<��a<ߨa<7�a<y�a<ũa<�a<c�a<��a<ߪa<�a<^�a<��a<ëa<�a<H�a<n�a<��a<ʬa<��a<-�a<J�a<�a<��a<��a<ѭa<�a<�a<?�a<F�a<K�a<v�a<��a<��a<��a<��a<��a<Ǯa<��a<ܮa<�a<ɮa<ۮa<߮a<Ϯa<ۮa<��a<��a<ɮa<��a<��a<��a<y�a<v�a<_�a<6�a<A�a<�a<�a<�a<��a<��a<��a<g�a<C�a<!�a<�a<ɬa<��a<i�a<\�a<�a<۫a<��a<��a<I�a<�a<ݪa<��a<e�a<!�a<�a<��a<R�a<$�a<ܨa<��a<I�a<�a<��a<k�a<�a<��a<l�a<�a<ťa<[�a<�a<��a<]�a<�a<��a<2�a<Ңa<i�a<�a<��a<7�a<��a<r�a<�a<��a<7�a<��a<M�a<�a<��a<�a<��a<6�a<ƛa<T�a<��a<��a<�a<��a<N�a<ۘa<|�a<
�a<��a<S�a<�a<z�a<$�a<Õa<k�a<�a<��a<c�a<�a<��a<c�a<�a<ϒa<��a<7�a<�a<��a<j�a<,�a<�a<��a<��a<Y�a<�a< �a<Џa<��a<��a<f�a<@�a<*�a<�a<�a<��a<ǎa<̎a<ǎa<��a<��a<��a<��a<Ўa<Ɏa<Ȏa<�a<�a<�a<(�a<�  �  ,�a<u�a<p�a<��a<Տa<�a<<�a<A�a<��a<��a<�a<?�a<m�a<ʑa<֑a<Y�a<{�a<�a<�a<h�a<ٓa<�a<��a<��a<6�a<��a<ޕa<Y�a<��a<#�a<b�a<��a<L�a<��a<(�a<r�a<�a<`�a<��a<C�a<ƛa<@�a<��a<+�a<��a<�a<p�a<�a<g�a<̟a<Q�a<��a<>�a<��a<�a<q�a<Ӣa<i�a<��a<>�a<y�a<��a<[�a<��a<*�a<t�a<�a<,�a<��a<�a<E�a<��a<Ѩa<N�a<s�a<�a<��a<Z�a<��a<ܪa<7�a<G�a<��a<ɫa<�a<?�a<l�a<��a<��a<�a<�a<Z�a<s�a<��a<ҭa<˭a<�a<�a<9�a<H�a<a�a<��a<n�a<��a<��a<Ůa<��a<Ǯa<ڮa<��a<�a<ʮa<�a<ʮa<Ӯa<�a<��a<ݮa<��a<Ůa<��a<��a<��a<_�a<r�a<2�a<F�a<�a<�a<�a<��a<��a<p�a<x�a<-�a<%�a<��a<ìa<��a<Q�a<`�a<	�a<��a<��a<u�a<^�a<�a<�a<��a<r�a<'�a<ߩa<��a<S�a<1�a<èa<��a<I�a<�a<��a<A�a<-�a<��a<��a<�a<��a<n�a<�a<��a<D�a<��a<��a<6�a<עa<e�a<�a<��a<P�a<Ƞa<y�a<��a<��a<B�a<��a<k�a<ҝa<��a<�a<��a<A�a<��a<h�a<�a<��a<�a<��a<Q�a<̘a<��a<�a<ȗa<3�a<�a<��a< �a<ޕa<T�a<�a<��a<l�a<�a<��a<u�a<
�a<ܒa<z�a<G�a<��a<��a<��a<&�a<�a<��a<��a<Z�a<-�a<�a<��a<��a<s�a<w�a<7�a<+�a<�a<�a<��a<Ȏa<��a<��a<��a<̎a<��a<Ԏa<��a<�a<̎a<�a<��a<��a<;�a<�  �  E�a<c�a<|�a<��a<ďa<��a<6�a<D�a<��a<Őa<�a<@�a<f�a<��a<�a<:�a<w�a<ܒa<�a<y�a<Ɠa<�a<��a<ؔa<�a<��a<�a<K�a<��a<�a<x�a<�a<;�a<��a</�a<��a<�a<c�a<ךa<V�a<ϛa<3�a<��a<�a<��a<��a<v�a<��a<`�a<ßa<I�a<��a<%�a<��a<��a<�a<�a<I�a<��a<(�a<��a<��a<M�a<��a<)�a<��a<զa<5�a<��a<�a<>�a<��a<�a<-�a<q�a<۩a<�a<b�a<��a<Ѫa< �a<d�a<��a<Ыa<�a<=�a<p�a<��a<۬a<�a<�a<G�a<{�a<��a<��a<˭a<�a<!�a<0�a<9�a<b�a<j�a<��a<��a<��a<��a<îa<��a<Ѯa<ˮa<خa<�a<ڮa<�a<ۮa<Įa<ʮa<ٮa<��a<Ʈa<��a<��a<��a<v�a<`�a<K�a<4�a<�a<�a<حa<̭a<��a<s�a<f�a<D�a<�a<��a<��a<��a<��a<A�a<�a<�a<��a<��a<K�a<�a<�a<��a<W�a<&�a<�a<��a<c�a<&�a<بa<��a<7�a<��a<��a<Y�a<"�a<��a<a�a<�a<ɥa<b�a<�a<��a<N�a<�a<��a<<�a<Тa<\�a<�a<��a<7�a<Ϡa<^�a<�a<��a<#�a<��a<U�a<�a<��a<�a<��a<?�a<̛a<U�a<�a<��a<�a<��a<S�a<�a<r�a<�a<��a<D�a<�a<��a<�a<ƕa<p�a<�a<��a<c�a<
�a<��a<\�a<%�a<ؒa<x�a<4�a<��a<��a<w�a<&�a<��a<ΐa<��a<K�a<.�a<�a<֏a<��a<s�a<o�a<K�a<!�a<�a<�a<�a<ߎa<ˎa<Ɏa<��a<��a<��a<Ўa<��a<�a<֎a<Ԏa<��a<�a<)�a<�  �  G�a<W�a<��a<��a<Ϗa<�a<�a<m�a<{�a<ېa<�a<,�a<��a<��a<��a<3�a<��a<��a<#�a<��a<��a<1�a<_�a<ݔa<�a<��a<�a<B�a<��a<��a<~�a<ٗa<^�a<��a<�a<��a<�a<��a<ޚa<O�a<��a<!�a<��a<�a<��a<��a<��a<�a<]�a<۟a<F�a<Ҡa<�a<��a<�a<n�a<�a<H�a<̣a<�a<��a<��a<_�a<åa<�a<��a<Цa<K�a<��a<�a</�a<��a<�a<0�a<��a<��a<�a<X�a<��a<��a<�a<e�a<��a<̫a<�a<@�a<{�a<��a<�a<�a<7�a<G�a<��a<��a<��a<��a<�a<�a<$�a<P�a<[�a<[�a<��a<��a<��a<��a<Ǯa<ɮa<Ʈa<�a<̮a<�a<��a<ޮa<Юa<ڮa<׮a<��a<Ȯa<��a<��a<��a<~�a<w�a<D�a<M�a<(�a<'�a<��a<�a<ԭa<��a<��a<T�a<Z�a<
�a<�a<ݬa<��a<z�a<:�a<4�a<Ыa<��a<��a<?�a<)�a<Ǫa<��a<Y�a<,�a<�a<��a<c�a<	�a<ߨa<��a<[�a<��a<��a<h�a<�a<Ӧa<h�a<�a<��a<P�a<�a<��a<i�a<�a<��a<2�a<΢a<u�a<�a<��a<�a<ݠa<d�a<��a<��a<!�a<Ϟa<6�a<��a<��a<�a<��a<.�a<՛a<P�a<�a<z�a<�a<��a<6�a<�a<u�a<*�a<��a<O�a<�a<{�a<=�a<��a<q�a<��a<��a<]�a<�a<Óa<Y�a<)�a<��a<��a<4�a<�a<��a<W�a<Q�a<�a<ɐa<��a<c�a<'�a<�a<�a<��a<��a<Q�a<P�a<,�a<	�a<�a<ݎa<ߎa<��a<Ǝa<��a<��a<Îa<��a<ώa<��a<ێa<�a<�a<�a<�a<�  �  E�a<b�a<��a<��a<Ϗa< �a<�a<k�a<s�a<��a<�a<3�a<w�a<��a<��a<6�a<��a<Вa<*�a<d�a<��a<#�a<g�a<הa<1�a<��a<�a<L�a<��a<!�a<��a<җa<A�a<��a< �a<��a<��a<{�a<ۚa<P�a<ԛa<D�a<��a<�a<��a<�a<{�a<�a<T�a<џa<'�a<��a<0�a<��a<�a<t�a<�a<L�a<��a<)�a<��a<٤a<T�a<��a<�a<��a<�a<4�a<��a<��a<M�a<��a<�a<.�a<��a<ɩa<�a<Z�a<��a<ܪa<�a<i�a<��a<ޫa<�a<=�a<m�a<��a<ܬa<��a<%�a<B�a<_�a<��a<��a<�a<�a<�a<*�a<G�a<_�a<�a<|�a<z�a<��a<��a<��a<Įa<ʮa<Ѯa<خa<�a<�a<�a<ɮa<Ϯa<Ԯa<��a<Юa<��a<��a<��a<s�a<��a<j�a<K�a<2�a<�a<��a<�a<̭a<��a<��a<L�a<5�a<)�a<�a<ͬa<��a<p�a<=�a<!�a<�a<��a<q�a<;�a<�a<Ϫa<��a<m�a<#�a<�a<��a<i�a<.�a<�a<��a<>�a< �a<��a<g�a<�a<ɦa<e�a<�a<Υa<s�a<�a<��a<M�a<�a<��a<3�a<Ģa<k�a<�a<��a<B�a<֠a<f�a<��a<��a<%�a<Þa<W�a<�a<_�a<	�a<��a<3�a<ћa<a�a<�a<��a<)�a<��a<Z�a<�a<s�a<�a<��a<M�a<�a<��a< �a<��a<v�a<#�a<Ôa<i�a<
�a<��a<q�a<%�a<ƒa<��a</�a<�a<��a<p�a<=�a<�a<��a<��a<Y�a<+�a<	�a<ɏa<��a<��a<V�a<I�a<'�a<�a<��a<�a<ގa<؎a<ӎa<��a<��a<��a<��a<׎a<��a<ގa<�a<�a<�a<3�a<�  �  2�a<e�a<}�a<��a<��a<��a<2�a<T�a<��a<��a<��a<-�a<k�a<��a<��a<I�a<y�a<Ԓa<"�a<u�a<�a<�a<��a<��a<�a<��a<�a<C�a<��a<�a<h�a<��a<7�a<��a<+�a<��a<�a<`�a<�a<P�a<��a</�a<��a<%�a<��a<�a<^�a<��a<[�a<ߟa<\�a<��a<*�a<��a<�a<}�a<�a<Y�a<��a<*�a<��a<�a<n�a<��a<-�a<f�a<�a<7�a<��a<ߧa<6�a<��a<ܨa<@�a<q�a<ܩa<�a<_�a<��a<ͪa<6�a<N�a<��a<ūa<�a<D�a<t�a<��a<��a<�a<�a<s�a<{�a<��a<��a<ǭa<�a<�a<9�a<?�a<P�a<s�a<��a<��a<��a<��a<��a<��a<�a<Ϯa<�a<Ȯa<׮a<ͮa<�a<ɮa<Ǯa<ծa<��a<��a<��a<��a<��a<`�a<[�a<8�a<6�a<�a<�a<ʭa<ía<��a<��a<��a<=�a<�a<�a<��a<��a<x�a<Q�a<�a<�a<��a<��a<r�a<�a<�a<��a<[�a<.�a<�a<��a<T�a<�a<ɨa<��a<3�a<�a<��a<\�a<!�a<��a<n�a<�a<��a<^�a<��a<��a<N�a<�a<y�a<>�a<ˢa<y�a<�a<��a<<�a<��a<l�a<�a<��a<2�a<��a<W�a<�a<��a<#�a<��a<D�a<��a<i�a<�a<��a<�a<��a<>�a<טa<��a<�a<��a<H�a<�a<��a<�a<ݕa<[�a<�a<��a<Y�a<�a<��a<g�a<�a<�a<w�a<`�a<��a<��a<w�a<"�a<�a<Ða<��a<R�a<�a<��a<Џa<͏a<��a<l�a<G�a<�a<#�a<��a<��a<Ǝa<Ȏa<��a<Ȏa<��a<��a<̎a<��a<َa<׎a<؎a<�a<��a<$�a<�  �  I�a<^�a<y�a<��a<ˏa<�a<%�a<E�a<}�a<��a<��a<:�a<��a<��a<�a<<�a<��a<Ԓa<#�a<[�a<ēa<	�a<x�a<ϔa<+�a<��a<�a<H�a<��a<!�a<v�a<�a<G�a<��a<!�a<��a<��a<o�a<�a<Z�a<ța<P�a<��a<�a<��a<�a<r�a<�a<O�a<ɟa<.�a<��a< �a<��a<�a<k�a<բa<T�a<Σa<�a<��a<ܤa<R�a<��a<'�a<y�a<�a<3�a<��a<�a<Y�a<��a<�a<:�a<�a<ĩa<�a<\�a<��a<ުa<-�a<^�a<��a<�a<�a<>�a<r�a<��a<Ϭa<�a<�a<J�a<[�a<��a<��a<�a<��a<�a<*�a<R�a<g�a<j�a<}�a<��a<��a<��a<Ʈa<®a<ծa<̮a<֮a<ޮa<�a<خa<�a<ɮa<ήa<��a<��a<��a<��a<��a<��a<o�a<n�a<P�a</�a<�a<�a<�a<ͭa<��a<s�a<V�a<4�a<�a<��a<٬a<��a<c�a<C�a<+�a<�a<��a<h�a<H�a<�a<�a<��a<g�a<*�a<�a<��a<r�a</�a<֨a<��a<C�a<��a<��a<c�a<�a<��a<j�a<�a<¥a<�a<�a<��a<K�a<��a<��a<:�a<��a<c�a<�a<��a<2�a<�a<o�a<��a<��a<.�a<ўa<M�a<�a<b�a<�a<��a<=�a<ěa<d�a<�a<��a<"�a<˙a<P�a<�a<�a<�a<��a<O�a<�a<��a<#�a<ӕa<j�a<�a<˔a<c�a<�a<��a<n�a<�a<Ԓa<r�a<7�a<ܑa<��a<q�a<I�a<��a<��a<��a<e�a<3�a<�a<ʏa<��a<r�a<_�a<N�a<%�a<�a<�a<�a<܎a<ݎa<��a<̎a<��a<��a<��a<Ďa<a<׎a<ގa<�a<�a<6�a<�  �  Ԏa<�a<+�a<I�a<v�a<��a<��a<�a<1�a<q�a<��a<ʐa<�a<P�a<��a<ܑa<4�a<m�a<ڒa<"�a<p�a<ԓa<�a<b�a<Ӕa</�a<��a<�a<D�a<��a<'�a<��a<��a<d�a<Řa<Q�a<��a<)�a<w�a<��a<o�a<ӛa<M�a<̜a<J�a<��a<+�a<��a<�a<��a<��a<��a<Ѡa<I�a<��a<�a<��a<�a<l�a<ѣa<_�a<��a<$�a<}�a<ɥa<6�a<��a<��a<R�a<��a<�a<I�a<��a<بa<L�a<��a<ީa<�a<]�a<��a<̪a<�a<G�a<�a<��a<�a<1�a<]�a<}�a<��a<�a<�a<9�a<j�a<h�a<��a<��a<��a<ݭa<�a<�a<(�a<P�a<V�a<}�a<\�a<[�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<k�a<��a<U�a<g�a<M�a<2�a<+�a<�a<�a<�a<٭a<��a<��a<d�a<O�a<[�a<!�a<�a<جa<��a<��a<Q�a<�a<��a<ثa<��a<��a<D�a<	�a<�a<��a<I�a<"�a<�a<��a<\�a<�a<̨a<��a<@�a<�a<��a<_�a</�a<��a<��a<�a<˥a<t�a<�a<��a<g�a<�a<��a<L�a<٢a<��a<6�a<��a<m�a<�a<��a<�a<��a<:�a<۞a<k�a<��a<��a<5�a<Мa<Y�a<՛a<u�a<�a<��a<9�a<��a<N�a<�a<��a<�a<̗a<P�a<�a<��a<0�a<ܕa<_�a<�a<��a<O�a<��a<��a<c�a<�a<��a<e�a<5�a<�a<��a<n�a<
�a<ؐa<��a<P�a<#�a<��a<��a<��a<��a<R�a<F�a<��a<ˎa<Վa<��a<��a<��a<l�a<d�a<b�a<U�a<U�a<f�a<J�a<��a<X�a<��a<��a<��a<��a<��a<�  �  ��a<�a<�a<C�a<n�a<��a<Џa<ߏa<$�a<M�a<��a<Ԑa<�a<^�a<��a<�a<'�a<s�a<��a<�a<a�a<��a<*�a<s�a<Ӕa<%�a<��a<��a<f�a<ǖa< �a<��a<�a<[�a<ǘa<?�a<��a<�a<��a<�a<t�a<��a<d�a<ќa<0�a<��a<"�a<��a<
�a<i�a<�a<Z�a<۠a<L�a<áa</�a<��a<�a<q�a<ޣa<5�a<��a<��a<i�a<�a<4�a<��a<�a<O�a<��a<�a<U�a<��a<��a<6�a<��a<ϩa<�a<V�a<��a<�a<�a<b�a<��a<ͫa<�a<#�a<b�a<��a<Ȭa<Ǭa<��a<�a<A�a<p�a<��a<��a<Эa<�a<��a<�a<&�a<'�a<D�a<E�a<n�a<��a<z�a<��a<x�a<��a<��a<��a<��a<��a<��a<�a<s�a<u�a<_�a<V�a<H�a<D�a<#�a<'�a<�a<��a<��a<��a<��a<��a<g�a<$�a<�a<�a<ʬa<��a<{�a<_�a<0�a<�a<˫a<��a<_�a<)�a<��a<��a<��a<[�a<"�a<ةa<��a<h�a</�a<�a<��a<S�a<��a<��a<a�a<�a<Ŧa<p�a<)�a<ԥa<x�a<-�a<Ϥa<l�a<��a<��a<C�a<��a<�a<�a<��a<F�a<�a<��a<#�a<��a<K�a<�a<o�a<�a<��a<�a<��a<D�a<�a<t�a<�a<��a<5�a<әa<q�a<��a<��a<+�a<��a<S�a<�a<��a<)�a<��a<v�a<�a<Ĕa<r�a<�a<��a<U�a<�a<��a<��a<�a<Бa<��a<E�a<�a<Ԑa<��a<f�a<4�a<��a<ˏa<��a<\�a<@�a<�a<�a<�a<Ŏa<��a<��a<��a<��a<��a<[�a<b�a<Z�a<S�a<R�a<c�a<b�a<s�a<��a<��a<��a<؎a<�  �  юa<�a<�a<[�a<e�a<��a<͏a<��a<K�a<]�a<��a<ېa<��a<T�a<��a<ޑa<�a<��a<Ȓa<!�a<��a<��a<)�a<a�a<Дa<6�a<��a<�a<A�a<��a<	�a<��a<�a<o�a<͘a<'�a<��a<�a<��a<��a<[�a<қa<H�a<֜a<6�a<ŝa<�a<��a<�a<��a<�a<c�a<�a<9�a<��a<$�a<��a<��a<\�a<�a<=�a<Ĥa<�a<q�a<�a<&�a<��a<�a<P�a<��a<�a<=�a<��a<��a<,�a<��a<éa<�a<o�a<��a<�a<�a<K�a<z�a<��a<��a<,�a<b�a<u�a<Ǭa<ˬa<�a<=�a<O�a<��a<{�a<��a<ía<�a<�a<�a<7�a<4�a<k�a<J�a<k�a<}�a<n�a<��a<��a<��a<��a<��a<z�a<��a<��a<��a<��a<U�a<s�a<_�a<H�a<B�a<�a<�a<�a<��a<ƭa<ʭa<��a<�a<d�a<&�a<:�a<�a<ܬa<��a<h�a<U�a<$�a<��a<��a<��a<o�a<B�a<�a<��a<��a<H�a<�a<�a<��a<b�a<
�a<Ψa<z�a<V�a<��a<ħa<g�a<�a<ۦa<g�a<,�a<åa<`�a<�a<��a<q�a<��a<��a<7�a<��a<��a<"�a<סa<O�a<��a<r�a<�a<��a<>�a<Ӟa<Z�a<�a<��a<C�a<ɜa<L�a<�a<e�a<�a<��a<7�a<��a<J�a<�a<z�a<0�a<��a<j�a<�a<��a<B�a<��a<~�a<��a<��a<J�a< �a<��a<^�a<�a<��a<��a<�a<��a<��a<S�a<!�a<��a<��a<Y�a<*�a<�a<Ǐa<��a<i�a<g�a<�a<�a<�a<��a<Îa<��a<��a<e�a<f�a<J�a<^�a<[�a<X�a<l�a<C�a<v�a<{�a<��a<��a<��a<��a<�  �  ގa<�a< �a<G�a<s�a<��a<��a<�a<�a<Y�a<��a<ΐa<&�a<U�a<��a<�a<9�a<m�a<˒a<	�a<P�a<͓a<�a<w�a<Δa<.�a<��a<��a<R�a<ʖa<0�a<��a<��a<]�a<��a<8�a<��a<�a<�a<��a<��a<�a<W�a<ɜa<>�a<��a</�a<��a<�a<��a<��a<h�a<Ӡa<N�a<ȡa<(�a<��a<�a<x�a<ԣa<E�a<��a<�a<y�a<֥a<>�a<��a<�a<L�a<��a<��a<k�a<��a<�a<7�a<��a<Ωa<�a<W�a<��a<Ԫa<#�a<i�a<��a<ɫa<��a<-�a<Z�a<��a<��a<�a<��a<�a<U�a<g�a<��a<��a<ȭa<�a<�a<�a<"�a<8�a<1�a<h�a<]�a<{�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<t�a<p�a<\�a<X�a<M�a<3�a<@�a<"�a<��a<�a<έa<��a<��a<��a<R�a<K�a<��a<�a<Ϭa<��a<��a<V�a<'�a<��a<ݫa<��a<r�a<+�a<�a<٪a<��a<^�a<�a<�a<��a<f�a<�a<�a<��a<A�a<�a<��a<Z�a<�a<æa<p�a<�a<Υa<��a<#�a<��a<d�a<�a<��a<Q�a<�a<��a<&�a<��a<S�a<�a<��a<(�a<��a<D�a<�a<v�a<��a<��a<�a<��a<U�a<�a<~�a<�a<��a<2�a<˙a<a�a<�a<��a<�a<��a<R�a<�a<��a<*�a<Еa<g�a<�a<˔a<]�a<�a<��a<_�a<
�a<��a<n�a</�a<ʑa<��a<Y�a<	�a<�a<��a<]�a<,�a<�a<ďa<��a<m�a<-�a<1�a<��a<�a<юa<��a<��a<��a<t�a<v�a<z�a<V�a<T�a<U�a<S�a<^�a<_�a<t�a<��a<��a<Ŏa<ӎa<�  �  �a<��a<)�a<?�a<j�a<��a<��a<�a<�a<��a<��a<ːa<�a<B�a<��a<Αa<<�a<_�a<ǒa<*�a<`�a<ۓa<��a<��a<��a</�a<��a<�a<Z�a<��a<�a<|�a<�a<Y�a<͘a<P�a<��a<-�a<��a<��a<f�a<՛a<b�a<��a<S�a<��a<1�a<��a<�a<��a<�a<��a<��a<V�a<��a<+�a<��a<��a<��a<£a<Z�a<��a<�a<~�a<ɥa<A�a<��a<�a<E�a<��a<�a<A�a<��a<�a<R�a<v�a<�a<�a<M�a<��a<Ѫa<�a<A�a<��a<ǫa<��a<5�a<G�a<��a<��a<��a<�a<8�a<Y�a<Z�a<��a<��a<ܭa<حa<�a<�a<�a<^�a<<�a<x�a<X�a<z�a<~�a<x�a<��a<��a<��a<�a<��a<��a<��a<��a<n�a<��a<_�a<_�a<Z�a<*�a<"�a<��a<�a<�a<׭a<��a<��a<��a<H�a<X�a<�a<�a<Ȭa<��a<��a<C�a<<�a<�a<�a<��a<n�a<L�a<��a<�a<y�a<j�a<�a<�a<��a<_�a<#�a<èa<��a<<�a<�a<��a<g�a<.�a<��a<��a<'�a<ĥa<k�a<�a<ͤa<\�a<�a<��a<R�a<ޢa<��a<2�a<��a<n�a<Ҡa<��a<�a<��a<O�a<ўa<��a<�a<��a<)�a<ǜa<Z�a<՛a<��a<��a<��a<,�a<ϙa<U�a<�a<��a<#�a<җa<F�a<�a<��a< �a<�a<d�a<�a<��a<`�a<�a<��a<g�a<��a<͒a<Y�a<>�a<ۑa<��a<\�a<��a<�a<��a<r�a<�a<��a<Ǐa<��a<��a<9�a<A�a<�a<�a<Ɏa<��a<��a<~�a<��a<W�a<[�a<N�a<f�a<a�a<M�a<|�a<b�a<{�a<��a<��a<��a<��a<�  �  �a<��a<�a<T�a<h�a<��a<Ïa<�a<3�a<W�a<��a<�a<�a<P�a<��a<Ցa<&�a<��a<��a<�a<m�a<��a<�a<w�a<̔a<8�a<��a<�a<S�a<��a<'�a<��a<ߗa<[�a<Ҙa<&�a<��a<�a<��a<��a<{�a<�a<\�a<Üa<<�a<��a<'�a<��a<�a<|�a<��a<Z�a<ߠa<\�a<��a<.�a<��a<��a<z�a<�a<5�a<��a<�a<l�a<ѥa<7�a<��a<�a<E�a<��a<��a<X�a<��a<�a<(�a<��a<��a<�a<Z�a<��a<�a<�a<\�a<��a<ëa<�a<4�a<Z�a<��a<��a<׬a<�a<(�a<B�a<��a<��a<��a<׭a<�a<�a<+�a<#�a<.�a<R�a<T�a<d�a<r�a<x�a<��a<��a<��a<��a<��a<��a<��a<��a<w�a<��a<V�a<s�a<R�a<?�a<G�a<0�a<�a<�a<�a<ƭa<ía<��a<|�a<Y�a<3�a<#�a<�a<Ǭa<��a<u�a<Q�a<:�a<�a<ʫa<��a<_�a<4�a<�a<��a<��a<^�a<�a<�a<��a<]�a<�a<ިa<��a<S�a<�a<��a<l�a<�a<Ҧa<b�a<"�a<ͥa<��a<�a<Ǥa<^�a<�a<��a<H�a<�a<}�a<�a<��a<F�a<�a<��a<�a<��a<L�a<˞a<x�a<�a<��a<&�a<��a<G�a<ݛa<v�a<�a<��a<,�a<ʙa<`�a<��a<��a<$�a<��a<`�a<�a<��a<-�a<��a<t�a<�a<��a<_�a<�a<��a<f�a<�a<��a<g�a<�a<ޑa<��a<F�a<,�a<Ӑa<��a<m�a<)�a<�a<ߏa<��a<c�a<O�a<�a<��a<�a<a<��a<��a<��a<~�a<j�a<l�a<d�a<Q�a<K�a<j�a<E�a<v�a<n�a<y�a<��a<��a<ǎa<�  �  юa<�a<�a<M�a<t�a<��a<܏a<�a<@�a<K�a<��a<ѐa<�a<k�a<��a<��a<�a<~�a<��a<�a<r�a<��a<,�a<d�a<ܔa<.�a<��a< �a<G�a<ϖa<�a<��a<�a<]�a<ژa<%�a<Ǚa<��a<��a<�a<r�a<�a<P�a<؜a</�a<Ɲa<#�a<��a<�a<}�a<�a<T�a<�a<:�a<ǡa<*�a<��a<�a<Z�a<�a<0�a<��a<�a<u�a<�a<,�a<��a<�a<W�a<��a<��a<U�a<��a<��a<"�a<��a<��a<�a<_�a<��a<�a<�a<g�a<��a<Ыa<��a<(�a<m�a<{�a<Ŭa<׬a<�a<-�a<>�a<�a<w�a<Эa<��a<��a<��a<	�a<2�a<$�a<d�a<N�a<|�a<l�a<��a<��a<~�a<��a<��a<��a<��a<��a<��a<h�a<��a<V�a<|�a<E�a<I�a<9�a<�a<'�a<�a<��a<��a<��a<��a<o�a<s�a<-�a<0�a<�a<Ӭa<��a<r�a<l�a<�a<�a<��a<��a<b�a<2�a<�a<��a<��a<L�a<+�a<�a<��a<p�a<�a<�a<y�a<Q�a<�a<��a<t�a<�a<�a<Z�a</�a<��a<w�a<�a<��a<r�a<��a<��a<D�a<�a<��a<�a<ˡa<@�a<��a<s�a<&�a<��a<;�a<�a<X�a<�a<��a<5�a<��a<P�a<�a<l�a<�a<��a<>�a<ęa<[�a<��a<u�a<3�a<��a<n�a<�a<��a<3�a<��a<|�a<��a<ɔa<V�a<�a<��a<Z�a<�a<��a<�a<�a<�a<��a<B�a<!�a<��a<��a<K�a<>�a<�a<��a<��a<Y�a<a�a<�a<�a<܎a<ˎa<��a<��a<��a<i�a<u�a<W�a<S�a<[�a<<�a<u�a<D�a<~�a<a�a<��a<��a<��a<؎a<�  �  ֎a<��a<#�a<A�a<|�a<��a<ďa<��a<.�a<h�a<��a<ɐa<�a<b�a<��a<�a<�a<r�a<Βa<"�a<i�a<Ɠa<�a<m�a<֔a<'�a<��a<�a<L�a<��a<�a<��a<�a<O�a<ɘa<A�a<��a<�a<��a<�a<j�a<��a<N�a<a<A�a<��a<0�a<��a<�a<��a< �a<n�a<�a<9�a<��a<(�a<��a<�a<_�a<ߣa<G�a<��a<�a<w�a<Хa<;�a<��a<�a<E�a<��a<��a<H�a<��a<��a<@�a<t�a<ԩa<�a<J�a<��a<ݪa<
�a<S�a<��a<��a<��a<(�a<a�a<��a<��a<�a<�a<:�a<U�a<s�a<��a<��a<��a<�a<��a<�a<6�a<D�a<T�a<]�a<g�a<i�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<}�a<p�a<��a<^�a<O�a<c�a<.�a<�a<�a<��a<�a<ѭa<��a<��a<r�a<[�a<A�a<�a<��a<ެa<��a<|�a<b�a<�a<�a<��a<��a<t�a<D�a<�a<Ӫa<��a<T�a<%�a<کa<��a<Y�a<�a<ڨa<��a<E�a<�a<��a<d�a<�a<��a<s�a<6�a<��a<n�a<�a<��a<]�a<
�a<��a<Q�a<ޢa<��a<#�a<ġa<Z�a<�a<r�a<�a<��a<=�a<�a<]�a<�a<��a<4�a<a<R�a<ܛa<z�a<�a<��a<,�a<��a<W�a<�a<z�a</�a<��a<D�a<��a<��a<�a<ߕa<p�a<�a<��a<W�a<��a<��a<Z�a<�a<��a<h�a<+�a<ޑa<��a<Y�a<�a<Őa<��a<L�a<5�a<��a<��a<��a<y�a<P�a<&�a<�a<؎a<Վa<��a<��a<��a<l�a<o�a<\�a<M�a<q�a<P�a<O�a<p�a<a�a<k�a<��a<��a<��a<͎a<�  �  ��a<�a<0�a<?�a<i�a<��a<a<�a<�a<[�a<��a<�a<�a<R�a<��a<ґa<7�a<��a<��a<�a<Y�a<ѓa<�a<��a<��a</�a<��a<��a<m�a<��a<A�a<v�a<�a<]�a<��a<H�a<��a<+�a<r�a<�a<v�a<�a<l�a<��a<L�a<��a<6�a<��a<�a<��a<�a<c�a<Ҡa<c�a<��a<5�a<��a<��a<��a<٣a<@�a<��a<�a<{�a<ѥa<K�a<�a<��a<:�a<��a< �a<N�a<��a<Ԩa<L�a<x�a<کa<�a<S�a<��a<êa<5�a<I�a<��a<��a<�a<3�a<J�a<��a<��a<�a<��a<&�a<H�a<|�a<��a<��a<�a<�a<��a<,�a<�a<7�a<9�a<f�a<h�a<v�a<~�a<x�a<��a<t�a<��a<��a<��a<��a<t�a<��a<g�a<��a<Q�a<d�a<;�a<4�a<D�a<�a<�a<Эa<ޭa<��a<��a<��a<Y�a<K�a<�a<�a<��a<��a<��a<S�a<G�a<�a<۫a<��a<a�a<2�a<�a<ݪa<��a<g�a<�a<�a<��a<P�a<6�a<Ǩa<��a<6�a<��a<��a<Z�a<&�a<��a<��a<�a<ץa<{�a<�a<פa<O�a<�a<��a<W�a<�a<��a<!�a<��a<O�a<�a<��a<�a<��a<V�a<̞a<��a<�a<��a<�a<��a<V�a<ޛa<��a<��a<��a<!�a<ՙa<c�a<��a<��a<�a<̗a<H�a<��a<��a<'�a<ӕa<V�a<-�a<��a<r�a< �a<��a<e�a<��a<ϒa<f�a<4�a<Αa<��a<L�a<�a<�a<��a<|�a<-�a<��a<��a<��a<l�a<5�a</�a<�a<�a<Ȏa<��a<��a<l�a<��a<]�a<x�a<Z�a<A�a<f�a<E�a<q�a<T�a<��a<u�a<��a<Ɏa<��a<�  �  �a<��a<(�a<J�a<q�a<��a<ˏa<�a<:�a<y�a<��a<ېa<�a<J�a<��a<ݑa<)�a<q�a<Òa<1�a<u�a<��a<�a<r�a<ϔa<6�a<��a<�a<\�a<��a<�a<~�a<�a<o�a<˘a<5�a<��a<%�a<�a<��a<^�a<ӛa<^�a<Ȝa<B�a<��a<)�a<��a<�a<��a<�a<r�a<Ӡa<N�a<��a<%�a<��a<�a<o�a<Уa<M�a<ɤa<�a<z�a<ץa<8�a<��a<��a<I�a<��a<��a<;�a<��a<�a<C�a<��a<˩a<�a<f�a<��a<Ԫa<�a<<�a<��a<��a<��a<5�a<Z�a<��a<��a<߬a<�a<J�a<R�a<g�a<��a<��a<ʭa<٭a<��a<�a<#�a<P�a<^�a<[�a<q�a<t�a<��a<��a<��a<��a<��a<v�a<��a<��a<��a<��a<{�a<n�a<d�a<i�a<@�a<:�a<�a<��a<�a<߭a<֭a<��a<��a<{�a<a�a<:�a<*�a<�a<ʬa<��a<��a<K�a<)�a<��a<ͫa<��a<i�a<R�a<�a<ɪa<��a<Y�a<�a<�a<��a<U�a<%�a<��a<��a<>�a<��a<ħa<e�a<�a<ɦa<��a<�a<Υa<b�a<�a<ɤa<c�a<�a<��a<K�a<�a<��a<!�a<ӡa<^�a<�a<��a<�a<��a<D�a<؞a<m�a<��a<��a<G�a<��a<U�a<�a<w�a<�a<��a<0�a<̙a<W�a<�a<��a<�a<×a<Z�a<�a<��a<9�a<̕a<f�a<�a<��a<e�a<�a<��a<f�a<�a<��a<p�a<%�a<�a<��a<V�a<	�a<Ӑa<��a<`�a<�a<��a<Џa<��a<��a<[�a<$�a<�a<�a<ˎa<��a<��a<��a<��a<O�a<U�a<`�a<N�a<f�a<Y�a<\�a<g�a<��a<{�a<��a<��a<��a<�  �  Ɏa<�a< �a<@�a<��a<��a<ҏa<�a<%�a<K�a<��a<ѐa<�a<`�a<��a<��a<(�a<�a<ƒa< �a<d�a<��a<$�a<h�a<��a<�a<��a<�a<D�a<Ֆa<�a<��a<�a<H�a<Șa<0�a<��a<�a<��a<��a<��a<��a<F�a<ۜa<+�a<��a<$�a<��a<�a<o�a<�a<U�a<�a<?�a<ӡa<'�a<��a<�a<c�a<�a<3�a<��a<��a<j�a<إa<0�a<��a<�a<Y�a<��a<	�a<c�a<��a<��a<#�a<��a<ũa<�a<J�a<��a<�a<�a<p�a<��a<ƫa<�a<�a<m�a<��a<¬a<Ϭa<��a<�a<M�a<}�a<��a<ŭa<��a<�a<�a<�a<6�a<%�a<F�a<M�a<r�a<l�a<��a<��a<��a<��a<x�a<��a<��a<��a<��a<i�a<w�a<k�a<b�a<?�a<S�a<B�a<&�a<5�a<�a<�a<έa<��a<��a<s�a<i�a<,�a<�a<�a<۬a<��a<��a<a�a<�a<�a<̫a<��a<m�a<"�a<��a<��a<��a<O�a</�a<Ωa<��a<`�a<�a<��a<��a<V�a<��a<��a<c�a<�a<æa<]�a<.�a<ǥa<��a</�a<��a<v�a<��a<��a<E�a<�a<}�a<�a<��a<A�a<��a<x�a<2�a<��a<>�a<�a<a�a<�a<��a<�a<��a<E�a<�a<o�a<�a<��a<@�a<��a<l�a<�a<��a<4�a<��a<O�a<�a<��a<�a<��a<~�a<
�a<Ӕa<Z�a<�a<��a<K�a<�a<��a<}�a<�a<Бa<��a<Q�a<�a<ːa<��a<M�a<0�a<�a<a<��a<Z�a<B�a<�a<�a<܎a<֎a<��a<��a<��a<]�a<��a<g�a<_�a<b�a<<�a<V�a<Y�a<e�a<[�a<��a<��a<��a<�a<�  �  Ȏa<�a<+�a<G�a<j�a<��a<ӏa<�a<<�a<]�a<��a<ѐa<�a<P�a<��a<ڑa<&�a<}�a<͒a<�a<��a<ϓa<!�a<^�a<˔a<(�a<��a<�a<<�a<��a<�a<��a<��a<]�a<Ҙa<=�a<��a<�a<��a<�a<]�a<қa<@�a<ۜa<?�a<��a<�a<��a<�a<��a<�a<m�a<�a<A�a<��a<'�a<��a<�a<k�a<�a<J�a<��a<&�a<��a<إa<.�a<��a<�a<Z�a<��a<�a<;�a<��a<�a<9�a<��a<өa<�a<^�a<��a<۪a<
�a<E�a<s�a<«a<�a<%�a<Z�a<z�a<��a<�a<�a</�a<Y�a<{�a<��a<��a<ԭa<�a<��a<�a<5�a<;�a<^�a<o�a<t�a<h�a<w�a<��a<��a<��a<w�a<��a<��a<��a<��a<~�a<��a<w�a<m�a<R�a<G�a<2�a<�a<�a<�a<��a<ڭa<��a<��a<m�a<j�a<K�a<+�a<�a<ܬa<��a<~�a<Q�a<1�a<��a<ʫa<��a<t�a<4�a<�a<ܪa<��a<E�a<�a<۩a<��a<`�a<�a<̨a<}�a<G�a<�a<��a<l�a<�a<Ӧa<q�a< �a<��a<a�a<�a<��a<v�a<	�a<��a<A�a<�a<��a<6�a<ȡa<X�a<��a<{�a<�a<��a<F�a<؞a<i�a<�a<��a<3�a<Ҝa<[�a<�a<n�a<�a<��a<A�a<��a<E�a<��a<y�a<$�a<��a<d�a<��a<��a<1�a<͕a<m�a<�a<��a<C�a<�a<��a<W�a<�a<��a<x�a<4�a<�a<��a<]�a<�a<ѐa<��a<j�a<'�a<��a<a<��a<o�a<Z�a<7�a<�a<؎a<a<��a<��a<��a<]�a<d�a<Q�a<P�a<S�a<R�a<b�a<e�a<p�a<n�a<��a<��a<��a<��a<�  �  ��a<�a<�a<L�a<p�a<��a<ʏa<�a<&�a<f�a<��a<ܐa<!�a<G�a<��a<ӑa<:�a<q�a<��a<�a<a�a<��a<�a<y�a<Ԕa<8�a<u�a<�a<r�a<��a<4�a<��a<�a<b�a<��a<%�a<��a<�a<��a<�a<|�a<�a<d�a<��a<3�a<��a</�a<��a<�a<u�a<�a<m�a<ɠa<]�a<��a<.�a<��a<�a<��a<ǣa<I�a<��a<�a<n�a<�a<A�a<��a<�a<<�a<��a<
�a<[�a<��a<�a<5�a<��a<��a<�a<\�a<��a<Ѫa<0�a<X�a<��a<ëa<�a<0�a<a�a<��a<��a<լa<��a</�a<N�a<c�a<��a<��a<�a<ۭa<�a< �a<$�a<D�a<E�a<M�a<i�a<��a<�a<��a<z�a<��a<��a<��a<��a<��a<~�a<��a<v�a<a�a<a�a<b�a<=�a<E�a<7�a<�a<�a<ۭa<��a<��a<��a<��a<`�a</�a<�a<��a<ˬa<��a<��a<G�a<N�a<�a<ޫa<��a<g�a<9�a<��a<��a<��a<`�a<#�a<�a<��a<S�a<;�a<ިa<��a<C�a<��a<��a<Z�a<�a<��a<s�a<�a<�a<��a<)�a<Ϥa<X�a<��a<��a<P�a<�a<}�a<�a<��a<Y�a<ܠa<��a<�a<��a<R�a<ٞa<��a<�a<��a<%�a<��a<I�a<�a<��a<�a<��a<#�a<љa<m�a<�a<��a<�a<��a<S�a<�a<��a</�a<ɕa<d�a<(�a<��a<u�a<�a<��a<b�a<�a<ɒa<q�a<�a<ϑa<��a<R�a<�a<�a<��a<~�a<!�a<�a<ԏa<��a<y�a<A�a<�a<�a<�a<Ɏa<��a<��a<~�a<��a<o�a<m�a<m�a<K�a<b�a<T�a<P�a<d�a<~�a<x�a<��a<��a<ʎa<�  �  Ȏa<�a<+�a<G�a<j�a<��a<ӏa<�a<<�a<]�a<��a<ѐa<�a<P�a<��a<ڑa<&�a<}�a<͒a<�a<��a<ϓa<!�a<^�a<˔a<(�a<��a<�a<<�a<��a<�a<��a<��a<]�a<Ҙa<=�a<��a<�a<��a<�a<]�a<қa<@�a<ۜa<?�a<��a<�a<��a<�a<��a<�a<m�a<�a<A�a<��a<'�a<��a<�a<k�a<�a<J�a<��a<&�a<��a<إa<.�a<��a<�a<Z�a<��a<�a<;�a<��a<�a<9�a<��a<өa<�a<^�a<��a<۪a<
�a<E�a<s�a<«a<�a<%�a<Z�a<z�a<��a<�a<�a</�a<Y�a<{�a<��a<��a<ԭa<�a<��a<�a<5�a<;�a<^�a<o�a<t�a<h�a<w�a<��a<��a<��a<w�a<��a<��a<��a<��a<~�a<��a<w�a<m�a<R�a<G�a<2�a<�a<�a<�a<��a<ڭa<��a<��a<m�a<j�a<K�a<+�a<�a<ܬa<��a<~�a<Q�a<1�a<��a<ʫa<��a<t�a<4�a<�a<ܪa<��a<E�a<�a<۩a<��a<`�a<�a<̨a<}�a<G�a<�a<��a<l�a<�a<Ӧa<q�a< �a<��a<a�a<�a<��a<v�a<	�a<��a<A�a<�a<��a<6�a<ȡa<X�a<��a<{�a<�a<��a<F�a<؞a<i�a<�a<��a<3�a<Ҝa<[�a<�a<n�a<�a<��a<A�a<��a<E�a<��a<y�a<$�a<��a<d�a<��a<��a<1�a<͕a<m�a<�a<��a<C�a<�a<��a<W�a<�a<��a<x�a<4�a<�a<��a<]�a<�a<ѐa<��a<j�a<'�a<��a<a<��a<o�a<Z�a<7�a<�a<؎a<a<��a<��a<��a<]�a<d�a<Q�a<P�a<S�a<R�a<b�a<e�a<p�a<n�a<��a<��a<��a<��a<�  �  Ɏa<�a< �a<@�a<��a<��a<ҏa<�a<%�a<K�a<��a<ѐa<�a<`�a<��a<��a<(�a<�a<ƒa< �a<d�a<��a<$�a<h�a<��a<�a<��a<�a<D�a<Ֆa<�a<��a<�a<H�a<Șa<0�a<��a<�a<��a<��a<��a<��a<F�a<ۜa<+�a<��a<$�a<��a<�a<o�a<�a<U�a<�a<?�a<ӡa<'�a<��a<�a<c�a<�a<3�a<��a<��a<j�a<إa<0�a<��a<�a<Y�a<��a<	�a<c�a<��a<��a<#�a<��a<ũa<�a<J�a<��a<�a<�a<p�a<��a<ƫa<�a<�a<m�a<��a<¬a<Ϭa<��a<�a<M�a<}�a<��a<ŭa<��a<�a<�a<�a<6�a<%�a<F�a<M�a<r�a<l�a<��a<��a<��a<��a<x�a<��a<��a<��a<��a<i�a<w�a<k�a<b�a<?�a<S�a<B�a<&�a<5�a<�a<�a<έa<��a<��a<s�a<i�a<,�a<�a<�a<۬a<��a<��a<a�a<�a<�a<̫a<��a<m�a<"�a<��a<��a<��a<O�a</�a<Ωa<��a<`�a<�a<��a<��a<V�a<��a<��a<c�a<�a<æa<]�a<.�a<ǥa<��a</�a<��a<v�a<��a<��a<E�a<�a<}�a<�a<��a<A�a<��a<x�a<2�a<��a<>�a<�a<a�a<�a<��a<�a<��a<E�a<�a<o�a<�a<��a<@�a<��a<l�a<�a<��a<4�a<��a<O�a<�a<��a<�a<��a<~�a<
�a<Ӕa<Z�a<�a<��a<K�a<�a<��a<}�a<�a<Бa<��a<Q�a<�a<ːa<��a<M�a<0�a<�a<a<��a<Z�a<B�a<�a<�a<܎a<֎a<��a<��a<��a<]�a<��a<g�a<_�a<b�a<<�a<V�a<Y�a<e�a<[�a<��a<��a<��a<�a<�  �  �a<��a<(�a<J�a<q�a<��a<ˏa<�a<:�a<y�a<��a<ېa<�a<J�a<��a<ݑa<)�a<q�a<Òa<1�a<u�a<��a<�a<r�a<ϔa<6�a<��a<�a<\�a<��a<�a<~�a<�a<o�a<˘a<5�a<��a<%�a<�a<��a<^�a<ӛa<^�a<Ȝa<B�a<��a<)�a<��a<�a<��a<�a<r�a<Ӡa<N�a<��a<%�a<��a<�a<o�a<Уa<M�a<ɤa<�a<z�a<ץa<8�a<��a<��a<I�a<��a<��a<;�a<��a<�a<C�a<��a<˩a<�a<f�a<��a<Ԫa<�a<<�a<��a<��a<��a<5�a<Z�a<��a<��a<߬a<�a<J�a<R�a<g�a<��a<��a<ʭa<٭a<��a<�a<#�a<P�a<^�a<[�a<q�a<t�a<��a<��a<��a<��a<��a<v�a<��a<��a<��a<��a<{�a<n�a<d�a<i�a<@�a<:�a<�a<��a<�a<߭a<֭a<��a<��a<{�a<a�a<:�a<*�a<�a<ʬa<��a<��a<K�a<)�a<��a<ͫa<��a<i�a<R�a<�a<ɪa<��a<Y�a<�a<�a<��a<U�a<%�a<��a<��a<>�a<��a<ħa<e�a<�a<ɦa<��a<�a<Υa<b�a<�a<ɤa<c�a<�a<��a<K�a<�a<��a<!�a<ӡa<^�a<�a<��a<�a<��a<D�a<؞a<m�a<��a<��a<G�a<��a<U�a<�a<w�a<�a<��a<0�a<̙a<W�a<�a<��a<�a<×a<Z�a<�a<��a<9�a<̕a<f�a<�a<��a<e�a<�a<��a<f�a<�a<��a<p�a<%�a<�a<��a<V�a<	�a<Ӑa<��a<`�a<�a<��a<Џa<��a<��a<[�a<$�a<�a<�a<ˎa<��a<��a<��a<��a<O�a<U�a<`�a<N�a<f�a<Y�a<\�a<g�a<��a<{�a<��a<��a<��a<�  �  ��a<�a<0�a<?�a<i�a<��a<a<�a<�a<[�a<��a<�a<�a<R�a<��a<ґa<7�a<��a<��a<�a<Y�a<ѓa<�a<��a<��a</�a<��a<��a<m�a<��a<A�a<v�a<�a<]�a<��a<H�a<��a<+�a<r�a<�a<v�a<�a<l�a<��a<L�a<��a<6�a<��a<�a<��a<�a<c�a<Ҡa<c�a<��a<5�a<��a<��a<��a<٣a<@�a<��a<�a<{�a<ѥa<K�a<�a<��a<:�a<��a< �a<N�a<��a<Ԩa<L�a<x�a<کa<�a<S�a<��a<êa<5�a<I�a<��a<��a<�a<3�a<J�a<��a<��a<�a<��a<&�a<H�a<|�a<��a<��a<�a<�a<��a<,�a<�a<7�a<9�a<f�a<h�a<v�a<~�a<x�a<��a<t�a<��a<��a<��a<��a<t�a<��a<g�a<��a<Q�a<d�a<;�a<4�a<D�a<�a<�a<Эa<ޭa<��a<��a<��a<Y�a<K�a<�a<�a<��a<��a<��a<S�a<G�a<�a<۫a<��a<a�a<2�a<�a<ݪa<��a<g�a<�a<�a<��a<P�a<6�a<Ǩa<��a<6�a<��a<��a<Z�a<&�a<��a<��a<�a<ץa<{�a<�a<פa<O�a<�a<��a<W�a<�a<��a<!�a<��a<O�a<�a<��a<�a<��a<V�a<̞a<��a<�a<��a<�a<��a<V�a<ޛa<��a<��a<��a<!�a<ՙa<c�a<��a<��a<�a<̗a<H�a<��a<��a<'�a<ӕa<V�a<-�a<��a<r�a< �a<��a<e�a<��a<ϒa<f�a<4�a<Αa<��a<L�a<�a<�a<��a<|�a<-�a<��a<��a<��a<l�a<5�a</�a<�a<�a<Ȏa<��a<��a<l�a<��a<]�a<x�a<Z�a<A�a<f�a<E�a<q�a<T�a<��a<u�a<��a<Ɏa<��a<�  �  ֎a<��a<#�a<A�a<|�a<��a<ďa<��a<.�a<h�a<��a<ɐa<�a<b�a<��a<�a<�a<r�a<Βa<"�a<i�a<Ɠa<�a<m�a<֔a<'�a<��a<�a<L�a<��a<�a<��a<�a<O�a<ɘa<A�a<��a<�a<��a<�a<j�a<��a<N�a<a<A�a<��a<0�a<��a<�a<��a< �a<n�a<�a<9�a<��a<(�a<��a<�a<_�a<ߣa<G�a<��a<�a<w�a<Хa<;�a<��a<�a<E�a<��a<��a<H�a<��a<��a<@�a<t�a<ԩa<�a<J�a<��a<ݪa<
�a<S�a<��a<��a<��a<(�a<a�a<��a<��a<�a<�a<:�a<U�a<s�a<��a<��a<��a<�a<��a<�a<6�a<D�a<T�a<]�a<g�a<i�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<}�a<p�a<��a<^�a<O�a<c�a<.�a<�a<�a<��a<�a<ѭa<��a<��a<r�a<[�a<A�a<�a<��a<ެa<��a<|�a<b�a<�a<�a<��a<��a<t�a<D�a<�a<Ӫa<��a<T�a<%�a<کa<��a<Y�a<�a<ڨa<��a<E�a<�a<��a<d�a<�a<��a<s�a<6�a<��a<n�a<�a<��a<]�a<
�a<��a<Q�a<ޢa<��a<#�a<ġa<Z�a<�a<r�a<�a<��a<=�a<�a<]�a<�a<��a<4�a<a<R�a<ܛa<z�a<�a<��a<,�a<��a<W�a<�a<z�a</�a<��a<D�a<��a<��a<�a<ߕa<p�a<�a<��a<W�a<��a<��a<Z�a<�a<��a<h�a<+�a<ޑa<��a<Y�a<�a<Őa<��a<L�a<5�a<��a<��a<��a<y�a<P�a<&�a<�a<؎a<Վa<��a<��a<��a<l�a<o�a<\�a<M�a<q�a<P�a<O�a<p�a<a�a<k�a<��a<��a<��a<͎a<�  �  юa<�a<�a<M�a<t�a<��a<܏a<�a<@�a<K�a<��a<ѐa<�a<k�a<��a<��a<�a<~�a<��a<�a<r�a<��a<,�a<d�a<ܔa<.�a<��a< �a<G�a<ϖa<�a<��a<�a<]�a<ژa<%�a<Ǚa<��a<��a<�a<r�a<�a<P�a<؜a</�a<Ɲa<#�a<��a<�a<}�a<�a<T�a<�a<:�a<ǡa<*�a<��a<�a<Z�a<�a<0�a<��a<�a<u�a<�a<,�a<��a<�a<W�a<��a<��a<U�a<��a<��a<"�a<��a<��a<�a<_�a<��a<�a<�a<g�a<��a<Ыa<��a<(�a<m�a<{�a<Ŭa<׬a<�a<-�a<>�a<�a<w�a<Эa<��a<��a<��a<	�a<2�a<$�a<d�a<N�a<|�a<l�a<��a<��a<~�a<��a<��a<��a<��a<��a<��a<h�a<��a<V�a<|�a<E�a<I�a<9�a<�a<'�a<�a<��a<��a<��a<��a<o�a<s�a<-�a<0�a<�a<Ӭa<��a<r�a<l�a<�a<�a<��a<��a<b�a<2�a<�a<��a<��a<L�a<+�a<�a<��a<p�a<�a<�a<y�a<Q�a<�a<��a<t�a<�a<�a<Z�a</�a<��a<w�a<�a<��a<r�a<��a<��a<D�a<�a<��a<�a<ˡa<@�a<��a<s�a<&�a<��a<;�a<�a<X�a<�a<��a<5�a<��a<P�a<�a<l�a<�a<��a<>�a<ęa<[�a<��a<u�a<3�a<��a<n�a<�a<��a<3�a<��a<|�a<��a<ɔa<V�a<�a<��a<Z�a<�a<��a<�a<�a<�a<��a<B�a<!�a<��a<��a<K�a<>�a<�a<��a<��a<Y�a<a�a<�a<�a<܎a<ˎa<��a<��a<��a<i�a<u�a<W�a<S�a<[�a<<�a<u�a<D�a<~�a<a�a<��a<��a<��a<؎a<�  �  �a<��a<�a<T�a<h�a<��a<Ïa<�a<3�a<W�a<��a<�a<�a<P�a<��a<Ցa<&�a<��a<��a<�a<m�a<��a<�a<w�a<̔a<8�a<��a<�a<S�a<��a<'�a<��a<ߗa<[�a<Ҙa<&�a<��a<�a<��a<��a<{�a<�a<\�a<Üa<<�a<��a<'�a<��a<�a<|�a<��a<Z�a<ߠa<\�a<��a<.�a<��a<��a<z�a<�a<5�a<��a<�a<l�a<ѥa<7�a<��a<�a<E�a<��a<��a<X�a<��a<�a<(�a<��a<��a<�a<Z�a<��a<�a<�a<\�a<��a<ëa<�a<4�a<Z�a<��a<��a<׬a<�a<(�a<B�a<��a<��a<��a<׭a<�a<�a<+�a<#�a<.�a<R�a<T�a<d�a<r�a<x�a<��a<��a<��a<��a<��a<��a<��a<��a<w�a<��a<V�a<s�a<R�a<?�a<G�a<0�a<�a<�a<�a<ƭa<ía<��a<|�a<Y�a<3�a<#�a<�a<Ǭa<��a<u�a<Q�a<:�a<�a<ʫa<��a<_�a<4�a<�a<��a<��a<^�a<�a<�a<��a<]�a<�a<ިa<��a<S�a<�a<��a<l�a<�a<Ҧa<b�a<"�a<ͥa<��a<�a<Ǥa<^�a<�a<��a<H�a<�a<}�a<�a<��a<F�a<�a<��a<�a<��a<L�a<˞a<x�a<�a<��a<&�a<��a<G�a<ݛa<v�a<�a<��a<,�a<ʙa<`�a<��a<��a<$�a<��a<`�a<�a<��a<-�a<��a<t�a<�a<��a<_�a<�a<��a<f�a<�a<��a<g�a<�a<ޑa<��a<F�a<,�a<Ӑa<��a<m�a<)�a<�a<ߏa<��a<c�a<O�a<�a<��a<�a<a<��a<��a<��a<~�a<j�a<l�a<d�a<Q�a<K�a<j�a<E�a<v�a<n�a<y�a<��a<��a<ǎa<�  �  �a<��a<)�a<?�a<j�a<��a<��a<�a<�a<��a<��a<ːa<�a<B�a<��a<Αa<<�a<_�a<ǒa<*�a<`�a<ۓa<��a<��a<��a</�a<��a<�a<Z�a<��a<�a<|�a<�a<Y�a<͘a<P�a<��a<-�a<��a<��a<f�a<՛a<b�a<��a<S�a<��a<1�a<��a<�a<��a<�a<��a<��a<V�a<��a<+�a<��a<��a<��a<£a<Z�a<��a<�a<~�a<ɥa<A�a<��a<�a<E�a<��a<�a<A�a<��a<�a<R�a<v�a<�a<�a<M�a<��a<Ѫa<�a<A�a<��a<ǫa<��a<5�a<G�a<��a<��a<��a<�a<8�a<Y�a<Z�a<��a<��a<ܭa<حa<�a<�a<�a<^�a<<�a<x�a<X�a<z�a<~�a<x�a<��a<��a<��a<�a<��a<��a<��a<��a<n�a<��a<_�a<_�a<Z�a<*�a<"�a<��a<�a<�a<׭a<��a<��a<��a<H�a<X�a<�a<�a<Ȭa<��a<��a<C�a<<�a<�a<�a<��a<n�a<L�a<��a<�a<y�a<j�a<�a<�a<��a<_�a<#�a<èa<��a<<�a<�a<��a<g�a<.�a<��a<��a<'�a<ĥa<k�a<�a<ͤa<\�a<�a<��a<R�a<ޢa<��a<2�a<��a<n�a<Ҡa<��a<�a<��a<O�a<ўa<��a<�a<��a<)�a<ǜa<Z�a<՛a<��a<��a<��a<,�a<ϙa<U�a<�a<��a<#�a<җa<F�a<�a<��a< �a<�a<d�a<�a<��a<`�a<�a<��a<g�a<��a<͒a<Y�a<>�a<ۑa<��a<\�a<��a<�a<��a<r�a<�a<��a<Ǐa<��a<��a<9�a<A�a<�a<�a<Ɏa<��a<��a<~�a<��a<W�a<[�a<N�a<f�a<a�a<M�a<|�a<b�a<{�a<��a<��a<��a<��a<�  �  ގa<�a< �a<G�a<s�a<��a<��a<�a<�a<Y�a<��a<ΐa<&�a<U�a<��a<�a<9�a<m�a<˒a<	�a<P�a<͓a<�a<w�a<Δa<.�a<��a<��a<R�a<ʖa<0�a<��a<��a<]�a<��a<8�a<��a<�a<�a<��a<��a<�a<W�a<ɜa<>�a<��a</�a<��a<�a<��a<��a<h�a<Ӡa<N�a<ȡa<(�a<��a<�a<x�a<ԣa<E�a<��a<�a<y�a<֥a<>�a<��a<�a<L�a<��a<��a<k�a<��a<�a<7�a<��a<Ωa<�a<W�a<��a<Ԫa<#�a<i�a<��a<ɫa<��a<-�a<Z�a<��a<��a<�a<��a<�a<U�a<g�a<��a<��a<ȭa<�a<�a<�a<"�a<8�a<1�a<h�a<]�a<{�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<t�a<p�a<\�a<X�a<M�a<3�a<@�a<"�a<��a<�a<έa<��a<��a<��a<R�a<K�a<��a<�a<Ϭa<��a<��a<V�a<'�a<��a<ݫa<��a<r�a<+�a<�a<٪a<��a<^�a<�a<�a<��a<f�a<�a<�a<��a<A�a<�a<��a<Z�a<�a<æa<p�a<�a<Υa<��a<#�a<��a<d�a<�a<��a<Q�a<�a<��a<&�a<��a<S�a<�a<��a<(�a<��a<D�a<�a<v�a<��a<��a<�a<��a<U�a<�a<~�a<�a<��a<2�a<˙a<a�a<�a<��a<�a<��a<R�a<�a<��a<*�a<Еa<g�a<�a<˔a<]�a<�a<��a<_�a<
�a<��a<n�a</�a<ʑa<��a<Y�a<	�a<�a<��a<]�a<,�a<�a<ďa<��a<m�a<-�a<1�a<��a<�a<юa<��a<��a<��a<t�a<v�a<z�a<V�a<T�a<U�a<S�a<^�a<_�a<t�a<��a<��a<Ŏa<ӎa<�  �  юa<�a<�a<[�a<e�a<��a<͏a<��a<K�a<]�a<��a<ېa<��a<T�a<��a<ޑa<�a<��a<Ȓa<!�a<��a<��a<)�a<a�a<Дa<6�a<��a<�a<A�a<��a<	�a<��a<�a<o�a<͘a<'�a<��a<�a<��a<��a<[�a<қa<H�a<֜a<6�a<ŝa<�a<��a<�a<��a<�a<c�a<�a<9�a<��a<$�a<��a<��a<\�a<�a<=�a<Ĥa<�a<q�a<�a<&�a<��a<�a<P�a<��a<�a<=�a<��a<��a<,�a<��a<éa<�a<o�a<��a<�a<�a<K�a<z�a<��a<��a<,�a<b�a<u�a<Ǭa<ˬa<�a<=�a<O�a<��a<{�a<��a<ía<�a<�a<�a<7�a<4�a<k�a<J�a<k�a<}�a<n�a<��a<��a<��a<��a<��a<z�a<��a<��a<��a<��a<U�a<s�a<_�a<H�a<B�a<�a<�a<�a<��a<ƭa<ʭa<��a<�a<d�a<&�a<:�a<�a<ܬa<��a<h�a<U�a<$�a<��a<��a<��a<o�a<B�a<�a<��a<��a<H�a<�a<�a<��a<b�a<
�a<Ψa<z�a<V�a<��a<ħa<g�a<�a<ۦa<g�a<,�a<åa<`�a<�a<��a<q�a<��a<��a<7�a<��a<��a<"�a<סa<O�a<��a<r�a<�a<��a<>�a<Ӟa<Z�a<�a<��a<C�a<ɜa<L�a<�a<e�a<�a<��a<7�a<��a<J�a<�a<z�a<0�a<��a<j�a<�a<��a<B�a<��a<~�a<��a<��a<J�a< �a<��a<^�a<�a<��a<��a<�a<��a<��a<S�a<!�a<��a<��a<Y�a<*�a<�a<Ǐa<��a<i�a<g�a<�a<�a<�a<��a<Îa<��a<��a<e�a<f�a<J�a<^�a<[�a<X�a<l�a<C�a<v�a<{�a<��a<��a<��a<��a<�  �  ��a<�a<�a<C�a<n�a<��a<Џa<ߏa<$�a<M�a<��a<Ԑa<�a<^�a<��a<�a<'�a<s�a<��a<�a<a�a<��a<*�a<s�a<Ӕa<%�a<��a<��a<f�a<ǖa< �a<��a<�a<[�a<ǘa<?�a<��a<�a<��a<�a<t�a<��a<d�a<ќa<0�a<��a<"�a<��a<
�a<i�a<�a<Z�a<۠a<L�a<áa</�a<��a<�a<q�a<ޣa<5�a<��a<��a<i�a<�a<4�a<��a<�a<O�a<��a<�a<U�a<��a<��a<6�a<��a<ϩa<�a<V�a<��a<�a<�a<b�a<��a<ͫa<�a<#�a<b�a<��a<Ȭa<Ǭa<��a<�a<A�a<p�a<��a<��a<Эa<�a<��a<�a<&�a<'�a<D�a<E�a<n�a<��a<z�a<��a<x�a<��a<��a<��a<��a<��a<��a<�a<s�a<u�a<_�a<V�a<H�a<D�a<#�a<'�a<�a<��a<��a<��a<��a<��a<g�a<$�a<�a<�a<ʬa<��a<{�a<_�a<0�a<�a<˫a<��a<_�a<)�a<��a<��a<��a<[�a<"�a<ةa<��a<h�a</�a<�a<��a<S�a<��a<��a<a�a<�a<Ŧa<p�a<)�a<ԥa<x�a<-�a<Ϥa<l�a<��a<��a<C�a<��a<�a<�a<��a<F�a<�a<��a<#�a<��a<K�a<�a<o�a<�a<��a<�a<��a<D�a<�a<t�a<�a<��a<5�a<әa<q�a<��a<��a<+�a<��a<S�a<�a<��a<)�a<��a<v�a<�a<Ĕa<r�a<�a<��a<U�a<�a<��a<��a<�a<Бa<��a<E�a<�a<Ԑa<��a<f�a<4�a<��a<ˏa<��a<\�a<@�a<�a<�a<�a<Ŏa<��a<��a<��a<��a<��a<[�a<b�a<Z�a<S�a<R�a<c�a<b�a<s�a<��a<��a<��a<؎a<�  �  m�a<��a<Ďa<ӎa<�a<&�a<=�a<��a<��a<��a<�a<e�a<��a<͐a<$�a<a�a<��a<�a<M�a<��a<�a<_�a<��a<�a<\�a<Ĕa<2�a<t�a<�a<7�a<ǖa<�a<��a<�a<\�a<טa<:�a<̙a<�a<��a<�a<q�a<��a<f�a<�a<E�a<ӝa<,�a<��a<*�a<��a<�a<p�a<�a<b�a<��a<-�a<��a<�a<|�a<�a<\�a<��a<�a<m�a<�a<0�a<��a<��a<N�a<��a<�a<[�a<��a<�a<1�a<~�a<éa<�a<Y�a<x�a<٪a<�a<7�a<h�a<��a<�a<��a<8�a<I�a<��a<��a<�a<��a<�a<C�a<T�a<q�a<y�a<��a<��a<ĭa<��a<�a<
�a< �a<�a</�a<*�a<M�a<3�a<8�a<%�a<J�a<=�a<&�a<F�a<�a<!�a<��a<�a<�a<�a<�a<��a<��a<��a<��a<^�a<L�a<%�a<�a<�a<��a<��a<k�a<S�a<8�a<�a<Ϋa<��a<}�a<G�a<�a<�a<��a<��a<"�a<�a<©a<��a<Z�a<��a<ƨa<j�a<L�a<�a<��a<n�a<�a<Ŧa<g�a<6�a<��a<��a<�a<��a<j�a<�a<ģa<C�a<��a<~�a<$�a<ˡa<c�a<��a<��a<*�a<��a<C�a<מa<z�a<�a<��a<6�a<Ҝa<_�a<�a<m�a<�a<��a<J�a<Йa<b�a<�a<��a<3�a<��a<m�a<�a<��a<%�a<Εa<s�a<�a<��a<7�a<�a<��a<P�a<��a<��a<Q�a<�a<a<l�a<3�a<ߐa<��a<k�a<"�a<�a<��a<��a<W�a<�a<�a<̎a<��a<}�a<n�a<\�a<8�a<>�a<�a< �a<��a<��a<�a<׍a<��a<ٍa<�a<�a<�a<�a<$�a<H�a<?�a<�  �  f�a<��a<��a<Ύa<��a<,�a<g�a<��a<��a<�a<(�a<h�a<��a<�a<4�a<w�a<��a<�a<N�a<��a<��a<W�a<��a<	�a<d�a<��a<$�a<�a<�a<U�a<��a<�a<��a<��a<c�a<՘a<>�a<��a< �a<��a<�a<��a<�a<h�a<לa<N�a<͝a<C�a<��a<#�a<��a<��a<��a<�a<]�a<ܡa<I�a<��a<�a<��a<ޣa<^�a<��a<-�a<��a<�a<<�a<��a<��a<J�a<��a<�a<N�a<��a<�a</�a<|�a<éa<�a<B�a<��a<ͪa<�a<;�a<n�a<��a<Ϋa<
�a<<�a<m�a<��a<��a<ܬa<�a<&�a<2�a<`�a<��a<��a<��a<��a<֭a<ޭa<��a<�a<%�a<&�a<'�a<,�a<4�a<;�a<4�a<E�a<C�a<:�a<.�a<'�a<%�a<$�a<�a< �a<�a<�a<׭a<ȭa<��a<��a<y�a<Y�a<C�a<+�a<�a<�a<ìa<��a<y�a<V�a<&�a<�a<ޫa<��a<m�a<M�a<�a<�a<��a<{�a<J�a<�a<ʩa<~�a<L�a<�a<Ĩa<��a<A�a<�a<��a<\�a<�a<æa<k�a<�a<ťa<t�a<&�a<ͤa<c�a<�a<��a<L�a<��a<��a<:�a<ġa<h�a<�a<��a<!�a<��a<`�a<�a<|�a<�a<��a<(�a<Ӝa<X�a<��a<��a<�a<��a<3�a<Ιa<]�a<��a<��a<&�a<��a<O�a<�a<��a<&�a<��a<\�a< �a<��a<Q�a<�a<��a<F�a<�a<��a<U�a<�a<��a<i�a<,�a<ِa<��a<Z�a<.�a<��a<ďa<��a<V�a<,�a<��a<׎a<��a<��a<y�a<U�a<9�a<%�a<�a<��a<�a<��a<�a<ލa<ލa<�a<��a<��a<��a<�a<%�a<?�a<\�a<�  �  _�a<��a<��a<��a<��a<�a<\�a<w�a<ҏa<�a<,�a<p�a<��a<�a<�a<{�a<��a<�a<K�a<��a<
�a<F�a<��a<�a<s�a<��a<&�a<��a<ܕa<]�a<��a<+�a<��a<��a<p�a<Șa<U�a<��a<?�a<��a<�a<��a<�a<~�a<Ӝa<i�a<��a<0�a<��a<�a<��a<�a<��a<�a<`�a<͡a<7�a<��a<�a<��a<գa<k�a<��a<�a<{�a<եa<V�a<��a<�a<S�a<��a< �a<=�a<��a<�a<E�a<u�a<ũa<�a<I�a<��a<��a<�a<4�a<��a<��a<իa<�a<"�a<e�a<��a<��a<ެa<�a<1�a<1�a<c�a<b�a<��a<��a<ŭa<�a<٭a<�a<��a<�a<�a<'�a<C�a<)�a<R�a<.�a<M�a<-�a<9�a<B�a<$�a<<�a<�a<(�a<��a<��a<�a<��a<ϭa<��a<��a<r�a<k�a<F�a<�a<�a<׬a<ݬa<��a<}�a<^�a<!�a<�a<��a<��a<m�a<Y�a<
�a<ߪa<��a<j�a<B�a<�a<ةa<��a<O�a<�a<��a<��a<'�a<��a<��a<c�a<�a<��a<��a<�a<�a<h�a<�a<Ѥa<c�a<#�a<��a<g�a<�a<��a<+�a<��a<y�a<�a<��a<%�a<��a<Q�a<�a<~�a<�a<��a<�a<��a<W�a<�a<{�a<�a<��a<3�a<�a<f�a<��a<��a<�a<՗a<Q�a< �a<��a<(�a<Εa<c�a<�a<��a<W�a<�a<��a<Q�a<�a<��a<;�a<�a<��a<v�a<.�a<אa<��a<Y�a<1�a<ۏa<��a<��a<]�a<6�a<�a<�a<��a<��a<_�a<U�a<P�a<�a<,�a<��a<	�a<��a<�a<�a<ۍa<��a<ݍa<�a<��a<�a<)�a<(�a<c�a<�  �  l�a<��a<��a<ώa<��a<)�a<Y�a<��a<��a<��a<�a<a�a<��a<�a<0�a<y�a<��a<�a<Q�a<��a<��a<T�a<��a<
�a<_�a<��a<�a<��a<�a<Q�a<��a<$�a<��a<�a<j�a<јa<D�a<��a<$�a<��a<�a<|�a<��a<j�a<ٜa<N�a<ѝa<9�a<��a<�a<��a<�a<y�a<�a<h�a<ϡa<@�a<��a<�a<�a<�a<P�a<��a<�a<}�a<�a<=�a<��a<��a<S�a<��a<��a<Q�a<��a<�a<2�a<{�a<ũa<��a<C�a<��a<˪a<�a<2�a<r�a<��a<ӫa<�a<=�a<_�a<��a<��a<֬a<��a<�a<<�a<e�a<|�a<��a<��a<��a<ǭa<�a<�a<�a<�a<�a<+�a<*�a<*�a<>�a<;�a<:�a<=�a<E�a<0�a<!�a<,�a<�a<�a<��a<�a<�a<׭a<��a<��a<��a<o�a<[�a<D�a<(�a<�a<�a<��a<��a<k�a<O�a<1�a<�a<ګa<��a<w�a<E�a<�a<�a<��a<x�a<;�a<�a<ĩa<��a<<�a<�a<��a<��a<>�a<��a<��a<O�a<�a<��a<r�a<�a<ɥa<|�a<�a<��a<k�a<�a<��a<L�a<��a<��a<*�a<��a<\�a<��a<��a<(�a<ǟa<S�a<�a<��a<�a<��a<8�a<Ŝa<Q�a<�a<~�a<�a<��a<9�a<͙a<f�a<�a<��a<*�a<��a<N�a<�a<��a<(�a<��a<]�a<�a<��a<N�a<�a<��a<<�a<�a<��a<V�a< �a<��a<h�a<&�a<�a<��a<d�a<3�a<��a<��a<��a<T�a<�a<�a<юa<��a<��a<r�a<Y�a<7�a<�a<�a<�a<��a<��a<�a<��a<؍a<�a<ߍa<��a<�a<�a</�a<?�a<Q�a<�  �  ��a<}�a<��a<Վa<��a<1�a<J�a<��a<��a<�a<(�a<b�a<��a<Րa<>�a<Z�a<��a<��a<^�a<��a<�a<e�a<��a<�a<Q�a<ϔa< �a<}�a<��a<D�a<��a<�a<��a<�a<f�a<�a<:�a<��a<�a<��a<�a<��a<�a<W�a<�a<B�a<՝a<9�a<��a<.�a<��a<$�a<t�a<�a<R�a<ѡa<F�a<��a<�a<v�a<�a<E�a<��a<%�a<y�a<��a<.�a<��a<�a<Z�a<��a<�a<O�a<��a<�a<)�a<��a<ȩa<��a<Q�a<z�a<Ҫa<��a<I�a<q�a<��a<�a<��a<M�a<O�a<��a<��a<٬a<	�a<�a<>�a<G�a<��a<��a<��a<��a<ϭa<��a<ݭa<�a<�a<$�a<#�a<*�a<K�a<'�a<P�a<7�a<;�a<0�a<0�a<0�a<"�a<2�a<�a<�a<��a<׭a<حa<��a<��a<��a<��a<`�a<7�a<0�a<��a<��a<��a<��a<y�a<P�a<%�a<�a<�a<��a<t�a<=�a<�a<�a<��a<��a<)�a<�a<��a<��a<I�a<�a<֨a<v�a<C�a<�a<��a<V�a<�a<Ӧa<h�a<&�a<��a<u�a<�a<Ĥa<z�a<��a<ƣa<@�a<��a<��a<.�a<Сa<K�a<�a<��a<*�a<��a<U�a<�a<k�a<�a<��a<N�a<��a<_�a<��a<y�a<)�a<��a<P�a<��a<m�a<��a<��a<'�a<��a<^�a<�a<��a<+�a<��a<k�a<��a<��a<A�a< �a<��a<<�a<�a<��a<g�a<�a<őa<g�a<(�a<�a<��a<f�a<�a<�a<��a<�a<V�a<%�a<�a<��a<ǎa<��a<w�a<Q�a<7�a<=�a<�a<�a<�a<�a<ߍa<�a<�a<�a<�a<��a<�a<�a<�a<@�a<K�a<�  �  k�a<��a<��a<ݎa<��a<-�a<K�a<��a<��a<�a<*�a<l�a<��a<�a<�a<o�a<Ƒa<�a<P�a<��a<��a<b�a<��a<�a<a�a<Δa<�a<��a<�a<J�a<��a<#�a<��a<��a<X�a<Ęa<D�a<��a<4�a<��a<�a<}�a<��a<_�a<�a<[�a<͝a<>�a<��a</�a<��a<
�a<��a<��a<^�a<Ρa<:�a<��a<"�a<��a<�a<X�a<Ǥa<)�a<��a<�a<G�a<��a<�a<Q�a<��a<��a<H�a<��a<�a<6�a<p�a<��a<�a<S�a<��a<Ǫa<��a<8�a<s�a<��a<�a<	�a<8�a<]�a<��a<��a<جa<��a<&�a<I�a<\�a<o�a<��a<��a<ʭa<׭a<߭a<��a<�a<�a<%�a<-�a<7�a<?�a</�a<8�a<;�a<B�a<2�a<A�a<+�a<#�a<�a<�a<�a<�a<�a<حa<��a<��a<��a<~�a<h�a<F�a<,�a<��a<�a<Ĭa<��a<{�a<Z�a</�a<�a<ȫa<��a<��a<P�a<�a<ݪa<��a<��a<5�a<�a<Ʃa<��a<G�a<
�a<¨a<|�a<?�a<��a<��a<d�a<�a<��a<q�a<�a<٥a<p�a< �a<��a<k�a<�a<��a<Y�a<��a<��a<1�a<Сa<b�a<��a<��a<2�a<��a<R�a<�a<{�a<�a<��a<6�a<Μa<i�a<��a<��a<�a<��a<>�a<Ǚa<d�a<��a<��a<!�a<ȗa<V�a<�a<}�a<�a<ʕa<m�a<
�a<��a<F�a<�a<��a<?�a<��a<��a<Q�a<��a<đa<p�a<(�a<��a<��a<q�a<+�a<�a<��a<��a<b�a<,�a<��a<׎a<��a<��a<x�a<Z�a<E�a<1�a<	�a< �a<��a<��a<�a<�a<�a<�a<��a<�a<�a<�a<"�a<@�a<P�a<�  �  _�a<��a<��a<͎a<��a<(�a<g�a<t�a<��a<�a<1�a<_�a<��a<��a<�a<��a<��a<�a<V�a<��a<��a<I�a<��a<��a<Z�a<��a<#�a<��a<ѕa<Y�a<��a<(�a<}�a<��a<n�a<ʘa<Z�a<��a</�a<��a<�a<t�a<�a<~�a<Ϝa<V�a<��a<E�a<��a<�a<��a<�a<��a<ݠa<h�a<֡a<?�a<��a<�a<��a<�a<`�a<��a<"�a<��a<ϥa<J�a<��a<�a<Q�a<��a<�a<G�a<��a<Ҩa<D�a<y�a<ɩa<
�a<7�a<��a<��a<�a<%�a<x�a<��a<ȫa<�a<(�a<x�a<��a<��a<�a<��a<'�a<'�a<u�a<m�a<��a<��a<��a<ݭa<�a<�a<�a<"�a<"�a<�a<(�a<-�a<O�a<1�a<:�a<C�a<9�a<5�a<�a<>�a<�a<&�a<��a<�a<�a<ҭa<­a<��a<��a<w�a<X�a<=�a<'�a<�a<Ԭa<ʬa<��a<��a<M�a<'�a<�a<ǫa<«a<g�a<K�a<�a<�a<��a<m�a<R�a<��a<��a<}�a<L�a<�a<��a<��a<2�a<��a<��a<]�a<�a<��a<��a<�a<ӥa<q�a<*�a<��a<g�a<#�a<��a<T�a<ߢa<��a<1�a<��a<m�a<�a<��a<�a<Ɵa<Z�a<�a<��a<��a<��a<2�a<՜a<M�a<�a<��a<�a<��a<)�a<ߙa<d�a<�a<��a<�a<Ǘa<>�a<��a<��a<,�a<Ǖa<Q�a<�a<��a<W�a<ܓa<��a<J�a<��a<��a<A�a<�a<��a<d�a<4�a<�a<��a<O�a<D�a<�a<ɏa<��a<L�a<2�a<��a<�a<��a<��a<u�a<M�a<5�a<�a<*�a<��a<��a<��a<�a<�a<֍a< �a<ߍa<�a<��a<�a<*�a<:�a<V�a<�  �  y�a<��a<��a<֎a<�a<)�a<N�a<��a<��a<��a<(�a<q�a<��a<ڐa<�a<q�a<��a<�a<Q�a<��a<��a<N�a<��a<�a<i�a<Ɣa<'�a<�a<�a<N�a<��a<!�a<��a<��a<d�a<̘a<D�a<��a<,�a<��a<�a<��a<��a<e�a<�a<T�a<ϝa<7�a<��a<#�a<��a<�a<��a<��a<g�a<ɡa<6�a<��a<�a<��a<�a<T�a<��a< �a<{�a<�a<F�a<��a<��a<Z�a<��a<��a<I�a<��a<�a<1�a<v�a<��a<�a<Q�a<��a<ªa<�a<B�a<s�a<��a<ܫa<�a<?�a<X�a<��a<��a<ݬa<��a<-�a<;�a<]�a<i�a<��a<��a<˭a<حa<�a<��a<�a<�a<�a<5�a</�a<8�a<1�a<K�a<:�a<5�a<2�a<;�a<7�a<$�a<�a<�a<�a<��a<�a<ʭa<��a<��a<��a<�a<a�a<N�a<(�a< �a<�a<��a<��a<z�a<`�a<.�a<��a<ǫa<��a<u�a<U�a<�a<�a<��a<q�a<1�a<�a<Ωa<��a<O�a<�a<ʨa<��a<2�a<��a<��a<^�a<�a<��a<q�a<(�a<Хa<p�a<�a<ɤa<u�a<
�a<��a<R�a<��a<��a<.�a<ša<\�a<��a<��a<2�a<Ɵa<M�a<��a<��a<�a<��a<5�a<ɜa<[�a<�a<|�a<�a<��a<@�a<̙a<m�a<�a<��a<"�a<��a<]�a<�a<��a<#�a<a<k�a<�a<��a<L�a<��a<��a<G�a<��a<��a<X�a<��a<��a<m�a<-�a<��a<��a<c�a<+�a<�a<��a<��a<c�a<-�a<�a<Ԏa<��a<��a<p�a<c�a<<�a<)�a<�a<�a<��a<�a<�a<�a<�a<�a<ߍa<��a<�a<�a<#�a<2�a<S�a<�  �  ��a<��a<��a<Ǝa<�a<4�a<H�a<��a<��a<��a<�a<f�a<��a<�a<A�a<l�a<��a<�a<Q�a<��a<��a<e�a<��a<�a<W�a<��a<$�a<��a<��a<3�a<͖a<�a<��a<�a<Y�a<�a<.�a<��a<�a<��a<�a<{�a<��a<X�a<��a<B�a<ڝa<2�a<��a<2�a<��a<�a<r�a<��a<X�a<ءa<J�a<��a<$�a<x�a<�a<M�a<¤a<(�a<t�a<��a<.�a<��a<�a<W�a<��a<�a<_�a<��a<�a<�a<��a<��a<��a<H�a<~�a<ުa<�a<F�a<r�a<��a<�a<��a<K�a<P�a<��a<��a<Ӭa<��a<�a<F�a<T�a<��a<��a<��a<ía<ĭa<�a<�a<�a<�a<#�a<5�a<�a<H�a<'�a<R�a<,�a<D�a<?�a<+�a<'�a<�a<0�a<��a<��a<�a<�a<�a<��a<��a<��a<��a<Q�a<H�a<3�a<��a<��a<��a<��a<l�a<T�a<'�a< �a<�a<��a<}�a<C�a<�a<ުa<��a<��a<+�a<�a<��a<��a<L�a<�a<רa<e�a<R�a<�a<��a<R�a<�a<Цa<[�a<�a<��a<��a<�a<��a<u�a<��a<ȣa<A�a<�a<��a<0�a<ӡa<W�a<�a<��a<4�a<��a<\�a<��a<s�a<�a<��a<>�a<Üa<d�a<��a<u�a<)�a<��a<Q�a<Ùa<j�a<��a<�a<8�a<��a<W�a<ٖa<��a<!�a<��a<c�a<��a<��a<3�a<��a<��a<C�a<��a<��a<d�a<�a<ʑa<m�a<"�a<�a<��a<n�a<"�a<�a<��a<��a<[�a<�a<�a<̎a<Ǝa<��a<v�a<c�a<-�a<9�a<�a<�a<�a<��a<�a<ۍa<ލa<эa<�a<�a<��a<�a<'�a<I�a<>�a<�  �  o�a<��a<��a<Ԏa<��a<�a<X�a<��a<��a<�a<2�a<b�a<��a<�a<�a<x�a<��a<�a<c�a<��a<��a<P�a<��a<��a<[�a<Ôa<�a<��a<�a<F�a<��a<�a<��a<��a<b�a<֘a<K�a<��a<#�a<��a<
�a<x�a<��a<g�a<�a<R�a<ŝa<7�a<��a<�a<��a<�a<~�a<�a<\�a<ҡa<?�a<��a<�a<��a<�a<W�a<��a<#�a<�a<�a<>�a<��a<��a<O�a<��a<��a<L�a<��a<�a<:�a<~�a<��a<�a<G�a<��a<Ǫa<��a<2�a<q�a<��a<߫a<�a<.�a<c�a<��a<��a<۬a<�a<�a<7�a<^�a<t�a<��a<��a<��a<ۭa<�a<��a<�a<�a<�a<$�a<.�a<:�a<:�a<=�a<9�a<:�a</�a<0�a<.�a<,�a< �a<�a<�a<�a<֭a<֭a<��a<��a<��a<|�a<_�a<?�a<�a<
�a<�a<ìa<��a<��a<P�a<�a<	�a<ʫa<��a<n�a<C�a<"�a<�a<��a<t�a<A�a<��a<��a<��a<F�a<�a<èa<y�a<?�a<�a<��a<e�a<�a<Ħa<x�a<�a<ǥa<v�a<�a<��a<k�a<�a<��a<P�a<�a<��a</�a<��a<c�a< �a<��a<$�a<��a<V�a<�a<|�a<�a<��a<=�a<͜a<S�a<�a<�a<�a<��a<E�a<̙a<b�a<�a<��a<%�a<��a<U�a<��a<��a<$�a<ʕa<a�a<��a<��a<F�a<�a<��a<@�a<��a<��a<G�a<�a<��a<k�a<*�a<�a<��a<_�a<-�a<�a<Ïa<y�a<T�a<1�a<�a<ڎa<��a<��a<e�a<R�a<;�a<+�a<�a<�a<��a<�a<ލa<�a<�a<�a<�a<��a<�a<�a<�a<>�a<P�a<�  �  ^�a<��a<��a<ڎa<�a<!�a<l�a<v�a<ˏa<ݏa</�a<m�a<��a<��a<�a<��a<��a<�a<T�a<��a<�a<E�a<a<��a<w�a<��a<�a<��a<ܕa<i�a<��a<-�a<��a<�a<f�a<��a<G�a<��a<8�a<��a<�a<��a<�a<j�a<ʜa<h�a<ĝa<M�a<��a<"�a<��a<��a<��a<�a<m�a<ѡa<<�a<��a<�a<��a<ޣa<_�a<��a<&�a<��a<ݥa<V�a<��a<��a<L�a<��a<�a<5�a<��a<ܨa<5�a<p�a<��a<�a<G�a<��a<��a<�a<.�a<r�a<��a<ҫa<�a<+�a<y�a<��a<ìa<լa<��a<6�a<:�a<o�a<l�a<��a<��a<ŭa<�a<ԭa<�a<��a<)�a<!�a<+�a<=�a<�a<A�a<.�a<O�a<5�a</�a<D�a<$�a<-�a<��a<�a<��a<�a<�a<ɭa<֭a<��a<��a<a�a<e�a<L�a< �a<�a<׬a<լa<��a<��a<[�a<)�a<�a<ƫa<��a<o�a<Y�a<�a<֪a<��a<h�a<U�a<��a<ܩa<��a<7�a<�a<��a<��a<)�a< �a<��a<W�a<�a<��a<u�a<�a<ܥa<d�a<'�a<Ȥa<d�a<�a<��a<f�a<�a<��a<:�a<áa<m�a<�a<��a<(�a<˟a<U�a<�a<��a<�a<��a<)�a<Ԝa<a�a<��a<��a<�a<��a<+�a<˙a<_�a<��a<��a<�a<ϗa<H�a<�a<}�a<$�a<��a<a�a<�a<��a<d�a<�a<��a<5�a<�a<��a<D�a<�a<��a<~�a<%�a<ܐa<��a<b�a<=�a<�a<̏a<��a<]�a<5�a<�a<�a<��a<��a<t�a<Y�a<J�a<�a<�a<��a<
�a<�a<ލa<�a<ۍa<�a<ύa<��a<��a<�a<$�a<1�a<j�a<�  �  q�a<��a<��a<֎a<��a<'�a<S�a<�a<Ïa<��a<(�a<]�a<��a<�a<2�a<o�a<��a<�a<W�a<��a<�a<J�a<��a<�a<^�a<��a<(�a<��a<�a<O�a<��a<!�a<��a<�a<m�a<ݘa<E�a<��a<.�a<��a<�a<y�a<��a<t�a<�a<S�a<��a<>�a<��a<(�a<��a<�a<}�a<�a<^�a<ӡa<A�a<��a<�a<��a<�a<]�a<��a<�a<��a<ڥa<=�a<��a<�a<[�a<��a<�a<;�a<��a<ݨa<2�a<��a<ͩa<�a<A�a<��a<��a<�a<8�a<�a<��a<ݫa<�a<1�a<c�a<��a<��a<�a<��a<�a<9�a<W�a<|�a<��a<��a<��a<ѭa<�a< �a<�a<�a<"�a<�a<3�a<8�a<H�a<@�a<7�a<;�a<2�a<8�a<#�a<*�a<&�a<�a<��a<��a<�a<ͭa<��a<��a<��a<}�a<a�a<<�a<&�a<�a<߬a<ͬa<��a<z�a<K�a<)�a<�a<ܫa<��a<r�a<B�a<�a<�a<��a<n�a<>�a< �a<éa<��a<P�a<�a<ƨa<��a<0�a<��a<��a<Y�a<�a<˦a<s�a<�a<ҥa<g�a<"�a<��a<r�a<�a<��a<R�a<�a<��a<'�a<ɡa<h�a<�a<��a<#�a<��a<W�a<�a<z�a<�a<��a<<�a<Ҝa<b�a<�a<��a<�a<��a<B�a<ٙa<o�a<�a<��a<�a<Ɨa<I�a<�a<��a<0�a<��a<[�a<�a<��a<P�a<�a<��a<I�a<��a<��a<J�a<�a<��a<w�a<2�a<�a<��a<a�a<&�a<��a<��a<��a<N�a<'�a<�a<��a<��a<��a<u�a<M�a<@�a<)�a<"�a<	�a<�a<�a<�a<�a<ڍa<�a<��a<��a<��a<�a<"�a<5�a<Q�a<�  �  v�a<u�a<��a<ێa<��a<:�a<I�a<��a<��a<��a<$�a<a�a<��a<Րa</�a<e�a<֑a<��a<^�a<��a<�a<N�a<��a<�a<Y�a<Ɣa<�a<r�a<�a<D�a<a<�a<��a< �a<N�a<ʘa<=�a<��a<$�a<��a<�a<~�a<��a<S�a<�a<F�a<ԝa<G�a<��a<"�a<��a<�a<l�a<�a<i�a<ԡa<A�a<��a<0�a<m�a<��a<I�a<��a<�a<��a<�a</�a<��a<�a<S�a<��a<�a<F�a<��a<�a<.�a<m�a<��a<
�a<I�a<y�a<ͪa< �a<@�a<d�a<��a<�a<��a<J�a<]�a<��a<��a<�a<	�a<�a<X�a<Q�a<|�a<��a<��a<ía<ʭa<��a<�a<�a<�a<2�a<+�a</�a<3�a< �a<H�a<2�a<G�a<,�a<2�a<5�a<�a<�a<��a<�a<�a<խa<ݭa<��a<��a<z�a<y�a<f�a<C�a<9�a<��a<�a<��a<��a<v�a<O�a<B�a<�a<٫a<��a<��a<8�a<�a<�a<��a<q�a<7�a<�a<��a<��a<A�a<��a<ɨa<w�a<F�a<�a<��a<g�a<��a<��a<k�a<#�a<ȥa<p�a<)�a<¤a<r�a<��a<��a<D�a<��a<��a<%�a<áa<P�a<�a<��a<<�a<ȟa<X�a<�a<~�a<(�a<��a<H�a<��a<U�a<�a<��a<"�a<��a<E�a<��a<f�a<��a<��a<�a<��a<Y�a<�a<z�a<�a<Ǖa<c�a<��a<��a<I�a<��a<��a<5�a<��a<��a<c�a<��a<��a<\�a<0�a<�a<��a<��a< �a<��a<��a<��a<[�a< �a<�a<a<��a<��a<��a<X�a<<�a<%�a<��a<�a<�a<��a<܍a<�a<�a<Ӎa<�a<ލa<�a<�a<�a<E�a<H�a<�  �  q�a<��a<��a<֎a<��a<'�a<S�a<�a<Ïa<��a<(�a<]�a<��a<�a<2�a<o�a<��a<�a<W�a<��a<�a<J�a<��a<�a<^�a<��a<(�a<��a<�a<O�a<��a<!�a<��a<�a<m�a<ݘa<E�a<��a<.�a<��a<�a<y�a<��a<t�a<�a<S�a<��a<>�a<��a<(�a<��a<�a<}�a<�a<^�a<ӡa<A�a<��a<�a<��a<�a<]�a<��a<�a<��a<ڥa<=�a<��a<�a<[�a<��a<�a<;�a<��a<ݨa<2�a<��a<ͩa<�a<A�a<��a<��a<�a<8�a<�a<��a<ݫa<�a<1�a<c�a<��a<��a<�a<��a<�a<9�a<W�a<|�a<��a<��a<��a<ѭa<�a< �a<�a<�a<"�a<�a<3�a<8�a<H�a<@�a<7�a<;�a<2�a<8�a<#�a<*�a<&�a<�a<��a<��a<�a<ͭa<��a<��a<��a<}�a<a�a<<�a<&�a<�a<߬a<ͬa<��a<z�a<K�a<)�a<�a<ܫa<��a<r�a<B�a<�a<�a<��a<n�a<>�a< �a<éa<��a<P�a<�a<ƨa<��a<0�a<��a<��a<Y�a<�a<˦a<s�a<�a<ҥa<g�a<"�a<��a<r�a<�a<��a<R�a<�a<��a<'�a<ɡa<h�a<�a<��a<#�a<��a<W�a<�a<z�a<�a<��a<<�a<Ҝa<b�a<�a<��a<�a<��a<B�a<ٙa<o�a<�a<��a<�a<Ɨa<I�a<�a<��a<0�a<��a<[�a<�a<��a<P�a<�a<��a<I�a<��a<��a<J�a<�a<��a<w�a<2�a<�a<��a<a�a<&�a<��a<��a<��a<N�a<'�a<�a<��a<��a<��a<u�a<M�a<@�a<)�a<"�a<	�a<�a<�a<�a<�a<ڍa<�a<��a<��a<��a<�a<"�a<5�a<Q�a<�  �  ^�a<��a<��a<ڎa<�a<!�a<l�a<v�a<ˏa<ݏa</�a<m�a<��a<��a<�a<��a<��a<�a<T�a<��a<�a<E�a<a<��a<w�a<��a<�a<��a<ܕa<i�a<��a<-�a<��a<�a<f�a<��a<G�a<��a<8�a<��a<�a<��a<�a<j�a<ʜa<h�a<ĝa<M�a<��a<"�a<��a<��a<��a<�a<m�a<ѡa<<�a<��a<�a<��a<ޣa<_�a<��a<&�a<��a<ݥa<V�a<��a<��a<L�a<��a<�a<5�a<��a<ܨa<5�a<p�a<��a<�a<G�a<��a<��a<�a<.�a<r�a<��a<ҫa<�a<+�a<y�a<��a<ìa<լa<��a<6�a<:�a<o�a<l�a<��a<��a<ŭa<�a<ԭa<�a<��a<)�a<!�a<+�a<=�a<�a<A�a<.�a<O�a<5�a</�a<D�a<$�a<-�a<��a<�a<��a<�a<�a<ɭa<֭a<��a<��a<a�a<e�a<L�a< �a<�a<׬a<լa<��a<��a<[�a<)�a<�a<ƫa<��a<o�a<Y�a<�a<֪a<��a<h�a<U�a<��a<ܩa<��a<7�a<�a<��a<��a<)�a< �a<��a<W�a<�a<��a<u�a<�a<ܥa<d�a<'�a<Ȥa<d�a<�a<��a<f�a<�a<��a<:�a<áa<m�a<�a<��a<(�a<˟a<U�a<�a<��a<�a<��a<)�a<Ԝa<a�a<��a<��a<�a<��a<+�a<˙a<_�a<��a<��a<�a<ϗa<H�a<�a<}�a<$�a<��a<a�a<�a<��a<d�a<�a<��a<5�a<�a<��a<D�a<�a<��a<~�a<%�a<ܐa<��a<b�a<=�a<�a<̏a<��a<]�a<5�a<�a<�a<��a<��a<t�a<Y�a<J�a<�a<�a<��a<
�a<�a<ލa<�a<ۍa<�a<ύa<��a<��a<�a<$�a<1�a<j�a<�  �  o�a<��a<��a<Ԏa<��a<�a<X�a<��a<��a<�a<2�a<b�a<��a<�a<�a<x�a<��a<�a<c�a<��a<��a<P�a<��a<��a<[�a<Ôa<�a<��a<�a<F�a<��a<�a<��a<��a<b�a<֘a<K�a<��a<#�a<��a<
�a<x�a<��a<g�a<�a<R�a<ŝa<7�a<��a<�a<��a<�a<~�a<�a<\�a<ҡa<?�a<��a<�a<��a<�a<W�a<��a<#�a<�a<�a<>�a<��a<��a<O�a<��a<��a<L�a<��a<�a<:�a<~�a<��a<�a<G�a<��a<Ǫa<��a<2�a<q�a<��a<߫a<�a<.�a<c�a<��a<��a<۬a<�a<�a<7�a<^�a<t�a<��a<��a<��a<ۭa<�a<��a<�a<�a<�a<$�a<.�a<:�a<:�a<=�a<9�a<:�a</�a<0�a<.�a<,�a< �a<�a<�a<�a<֭a<֭a<��a<��a<��a<|�a<_�a<?�a<�a<
�a<�a<ìa<��a<��a<P�a<�a<	�a<ʫa<��a<n�a<C�a<"�a<�a<��a<t�a<A�a<��a<��a<��a<F�a<�a<èa<y�a<?�a<�a<��a<e�a<�a<Ħa<x�a<�a<ǥa<v�a<�a<��a<k�a<�a<��a<P�a<�a<��a</�a<��a<c�a< �a<��a<$�a<��a<V�a<�a<|�a<�a<��a<=�a<͜a<S�a<�a<�a<�a<��a<E�a<̙a<b�a<�a<��a<%�a<��a<U�a<��a<��a<$�a<ʕa<a�a<��a<��a<F�a<�a<��a<@�a<��a<��a<G�a<�a<��a<k�a<*�a<�a<��a<_�a<-�a<�a<Ïa<y�a<T�a<1�a<�a<ڎa<��a<��a<e�a<R�a<;�a<+�a<�a<�a<��a<�a<ލa<�a<�a<�a<�a<��a<�a<�a<�a<>�a<P�a<�  �  ��a<��a<��a<Ǝa<�a<4�a<H�a<��a<��a<��a<�a<f�a<��a<�a<A�a<l�a<��a<�a<Q�a<��a<��a<e�a<��a<�a<W�a<��a<$�a<��a<��a<3�a<͖a<�a<��a<�a<Y�a<�a<.�a<��a<�a<��a<�a<{�a<��a<X�a<��a<B�a<ڝa<2�a<��a<2�a<��a<�a<r�a<��a<X�a<ءa<J�a<��a<$�a<x�a<�a<M�a<¤a<(�a<t�a<��a<.�a<��a<�a<W�a<��a<�a<_�a<��a<�a<�a<��a<��a<��a<H�a<~�a<ުa<�a<F�a<r�a<��a<�a<��a<K�a<P�a<��a<��a<Ӭa<��a<�a<F�a<T�a<��a<��a<��a<ía<ĭa<�a<�a<�a<�a<#�a<5�a<�a<H�a<'�a<R�a<,�a<D�a<?�a<+�a<'�a<�a<0�a<��a<��a<�a<�a<�a<��a<��a<��a<��a<Q�a<H�a<3�a<��a<��a<��a<��a<l�a<T�a<'�a< �a<�a<��a<}�a<C�a<�a<ުa<��a<��a<+�a<�a<��a<��a<L�a<�a<רa<e�a<R�a<�a<��a<R�a<�a<Цa<[�a<�a<��a<��a<�a<��a<u�a<��a<ȣa<A�a<�a<��a<0�a<ӡa<W�a<�a<��a<4�a<��a<\�a<��a<s�a<�a<��a<>�a<Üa<d�a<��a<u�a<)�a<��a<Q�a<Ùa<j�a<��a<�a<8�a<��a<W�a<ٖa<��a<!�a<��a<c�a<��a<��a<3�a<��a<��a<C�a<��a<��a<d�a<�a<ʑa<m�a<"�a<�a<��a<n�a<"�a<�a<��a<��a<[�a<�a<�a<̎a<Ǝa<��a<v�a<c�a<-�a<9�a<�a<�a<�a<��a<�a<ۍa<ލa<эa<�a<�a<��a<�a<'�a<I�a<>�a<�  �  y�a<��a<��a<֎a<�a<)�a<N�a<��a<��a<��a<(�a<q�a<��a<ڐa<�a<q�a<��a<�a<Q�a<��a<��a<N�a<��a<�a<i�a<Ɣa<'�a<�a<�a<N�a<��a<!�a<��a<��a<d�a<̘a<D�a<��a<,�a<��a<�a<��a<��a<e�a<�a<T�a<ϝa<7�a<��a<#�a<��a<�a<��a<��a<g�a<ɡa<6�a<��a<�a<��a<�a<T�a<��a< �a<{�a<�a<F�a<��a<��a<Z�a<��a<��a<I�a<��a<�a<1�a<v�a<��a<�a<Q�a<��a<ªa<�a<B�a<s�a<��a<ܫa<�a<?�a<X�a<��a<��a<ݬa<��a<-�a<;�a<]�a<i�a<��a<��a<˭a<حa<�a<��a<�a<�a<�a<5�a</�a<8�a<1�a<K�a<:�a<5�a<2�a<;�a<7�a<$�a<�a<�a<�a<��a<�a<ʭa<��a<��a<��a<�a<a�a<N�a<(�a< �a<�a<��a<��a<z�a<`�a<.�a<��a<ǫa<��a<u�a<U�a<�a<�a<��a<q�a<1�a<�a<Ωa<��a<O�a<�a<ʨa<��a<2�a<��a<��a<^�a<�a<��a<q�a<(�a<Хa<p�a<�a<ɤa<u�a<
�a<��a<R�a<��a<��a<.�a<ša<\�a<��a<��a<2�a<Ɵa<M�a<��a<��a<�a<��a<5�a<ɜa<[�a<�a<|�a<�a<��a<@�a<̙a<m�a<�a<��a<"�a<��a<]�a<�a<��a<#�a<a<k�a<�a<��a<L�a<��a<��a<G�a<��a<��a<X�a<��a<��a<m�a<-�a<��a<��a<c�a<+�a<�a<��a<��a<c�a<-�a<�a<Ԏa<��a<��a<p�a<c�a<<�a<)�a<�a<�a<��a<�a<�a<�a<�a<�a<ߍa<��a<�a<�a<#�a<2�a<S�a<�  �  _�a<��a<��a<͎a<��a<(�a<g�a<t�a<��a<�a<1�a<_�a<��a<��a<�a<��a<��a<�a<V�a<��a<��a<I�a<��a<��a<Z�a<��a<#�a<��a<ѕa<Y�a<��a<(�a<}�a<��a<n�a<ʘa<Z�a<��a</�a<��a<�a<t�a<�a<~�a<Ϝa<V�a<��a<E�a<��a<�a<��a<�a<��a<ݠa<h�a<֡a<?�a<��a<�a<��a<�a<`�a<��a<"�a<��a<ϥa<J�a<��a<�a<Q�a<��a<�a<G�a<��a<Ҩa<D�a<y�a<ɩa<
�a<7�a<��a<��a<�a<%�a<x�a<��a<ȫa<�a<(�a<x�a<��a<��a<�a<��a<'�a<'�a<u�a<m�a<��a<��a<��a<ݭa<�a<�a<�a<"�a<"�a<�a<(�a<-�a<O�a<1�a<:�a<C�a<9�a<5�a<�a<>�a<�a<&�a<��a<�a<�a<ҭa<­a<��a<��a<w�a<X�a<=�a<'�a<�a<Ԭa<ʬa<��a<��a<M�a<'�a<�a<ǫa<«a<g�a<K�a<�a<�a<��a<m�a<R�a<��a<��a<}�a<L�a<�a<��a<��a<2�a<��a<��a<]�a<�a<��a<��a<�a<ӥa<q�a<*�a<��a<g�a<#�a<��a<T�a<ߢa<��a<1�a<��a<m�a<�a<��a<�a<Ɵa<Z�a<�a<��a<��a<��a<2�a<՜a<M�a<�a<��a<�a<��a<)�a<ߙa<d�a<�a<��a<�a<Ǘa<>�a<��a<��a<,�a<Ǖa<Q�a<�a<��a<W�a<ܓa<��a<J�a<��a<��a<A�a<�a<��a<d�a<4�a<�a<��a<O�a<D�a<�a<ɏa<��a<L�a<2�a<��a<�a<��a<��a<u�a<M�a<5�a<�a<*�a<��a<��a<��a<�a<�a<֍a< �a<ߍa<�a<��a<�a<*�a<:�a<V�a<�  �  k�a<��a<��a<ݎa<��a<-�a<K�a<��a<��a<�a<*�a<l�a<��a<�a<�a<o�a<Ƒa<�a<P�a<��a<��a<b�a<��a<�a<a�a<Δa<�a<��a<�a<J�a<��a<#�a<��a<��a<X�a<Ęa<D�a<��a<4�a<��a<�a<}�a<��a<_�a<�a<[�a<͝a<>�a<��a</�a<��a<
�a<��a<��a<^�a<Ρa<:�a<��a<"�a<��a<�a<X�a<Ǥa<)�a<��a<�a<G�a<��a<�a<Q�a<��a<��a<H�a<��a<�a<6�a<p�a<��a<�a<S�a<��a<Ǫa<��a<8�a<s�a<��a<�a<	�a<8�a<]�a<��a<��a<جa<��a<&�a<I�a<\�a<o�a<��a<��a<ʭa<׭a<߭a<��a<�a<�a<%�a<-�a<7�a<?�a</�a<8�a<;�a<B�a<2�a<A�a<+�a<#�a<�a<�a<�a<�a<�a<حa<��a<��a<��a<~�a<h�a<F�a<,�a<��a<�a<Ĭa<��a<{�a<Z�a</�a<�a<ȫa<��a<��a<P�a<�a<ݪa<��a<��a<5�a<�a<Ʃa<��a<G�a<
�a<¨a<|�a<?�a<��a<��a<d�a<�a<��a<q�a<�a<٥a<p�a< �a<��a<k�a<�a<��a<Y�a<��a<��a<1�a<Сa<b�a<��a<��a<2�a<��a<R�a<�a<{�a<�a<��a<6�a<Μa<i�a<��a<��a<�a<��a<>�a<Ǚa<d�a<��a<��a<!�a<ȗa<V�a<�a<}�a<�a<ʕa<m�a<
�a<��a<F�a<�a<��a<?�a<��a<��a<Q�a<��a<đa<p�a<(�a<��a<��a<q�a<+�a<�a<��a<��a<b�a<,�a<��a<׎a<��a<��a<x�a<Z�a<E�a<1�a<	�a< �a<��a<��a<�a<�a<�a<�a<��a<�a<�a<�a<"�a<@�a<P�a<�  �  ��a<}�a<��a<Վa<��a<1�a<J�a<��a<��a<�a<(�a<b�a<��a<Րa<>�a<Z�a<��a<��a<^�a<��a<�a<e�a<��a<�a<Q�a<ϔa< �a<}�a<��a<D�a<��a<�a<��a<�a<f�a<�a<:�a<��a<�a<��a<�a<��a<�a<W�a<�a<B�a<՝a<9�a<��a<.�a<��a<$�a<t�a<�a<R�a<ѡa<F�a<��a<�a<v�a<�a<E�a<��a<%�a<y�a<��a<.�a<��a<�a<Z�a<��a<�a<O�a<��a<�a<)�a<��a<ȩa<��a<Q�a<z�a<Ҫa<��a<I�a<q�a<��a<�a<��a<M�a<O�a<��a<��a<٬a<	�a<�a<>�a<G�a<��a<��a<��a<��a<ϭa<��a<ݭa<�a<�a<$�a<#�a<*�a<K�a<'�a<P�a<7�a<;�a<0�a<0�a<0�a<"�a<2�a<�a<�a<��a<׭a<حa<��a<��a<��a<��a<`�a<7�a<0�a<��a<��a<��a<��a<y�a<P�a<%�a<�a<�a<��a<t�a<=�a<�a<�a<��a<��a<)�a<�a<��a<��a<I�a<�a<֨a<v�a<C�a<�a<��a<V�a<�a<Ӧa<h�a<&�a<��a<u�a<�a<Ĥa<z�a<��a<ƣa<@�a<��a<��a<.�a<Сa<K�a<�a<��a<*�a<��a<U�a<�a<k�a<�a<��a<N�a<��a<_�a<��a<y�a<)�a<��a<P�a<��a<m�a<��a<��a<'�a<��a<^�a<�a<��a<+�a<��a<k�a<��a<��a<A�a< �a<��a<<�a<�a<��a<g�a<�a<őa<g�a<(�a<�a<��a<f�a<�a<�a<��a<�a<V�a<%�a<�a<��a<ǎa<��a<w�a<Q�a<7�a<=�a<�a<�a<�a<�a<ߍa<�a<�a<�a<�a<��a<�a<�a<�a<@�a<K�a<�  �  l�a<��a<��a<ώa<��a<)�a<Y�a<��a<��a<��a<�a<a�a<��a<�a<0�a<y�a<��a<�a<Q�a<��a<��a<T�a<��a<
�a<_�a<��a<�a<��a<�a<Q�a<��a<$�a<��a<�a<j�a<јa<D�a<��a<$�a<��a<�a<|�a<��a<j�a<ٜa<N�a<ѝa<9�a<��a<�a<��a<�a<y�a<�a<h�a<ϡa<@�a<��a<�a<�a<�a<P�a<��a<�a<}�a<�a<=�a<��a<��a<S�a<��a<��a<Q�a<��a<�a<2�a<{�a<ũa<��a<C�a<��a<˪a<�a<2�a<r�a<��a<ӫa<�a<=�a<_�a<��a<��a<֬a<��a<�a<<�a<e�a<|�a<��a<��a<��a<ǭa<�a<�a<�a<�a<�a<+�a<*�a<*�a<>�a<;�a<:�a<=�a<E�a<0�a<!�a<,�a<�a<�a<��a<�a<�a<׭a<��a<��a<��a<o�a<[�a<D�a<(�a<�a<�a<��a<��a<k�a<O�a<1�a<�a<ګa<��a<w�a<E�a<�a<�a<��a<x�a<;�a<�a<ĩa<��a<<�a<�a<��a<��a<>�a<��a<��a<O�a<�a<��a<r�a<�a<ɥa<|�a<�a<��a<k�a<�a<��a<L�a<��a<��a<*�a<��a<\�a<��a<��a<(�a<ǟa<S�a<�a<��a<�a<��a<8�a<Ŝa<Q�a<�a<~�a<�a<��a<9�a<͙a<f�a<�a<��a<*�a<��a<N�a<�a<��a<(�a<��a<]�a<�a<��a<N�a<�a<��a<<�a<�a<��a<V�a< �a<��a<h�a<&�a<�a<��a<d�a<3�a<��a<��a<��a<T�a<�a<�a<юa<��a<��a<r�a<Y�a<7�a<�a<�a<�a<��a<��a<�a<��a<؍a<�a<ߍa<��a<�a<�a</�a<?�a<Q�a<�  �  _�a<��a<��a<��a<��a<�a<\�a<w�a<ҏa<�a<,�a<p�a<��a<�a<�a<{�a<��a<�a<K�a<��a<
�a<F�a<��a<�a<s�a<��a<&�a<��a<ܕa<]�a<��a<+�a<��a<��a<p�a<Șa<U�a<��a<?�a<��a<�a<��a<�a<~�a<Ӝa<i�a<��a<0�a<��a<�a<��a<�a<��a<�a<`�a<͡a<7�a<��a<�a<��a<գa<k�a<��a<�a<{�a<եa<V�a<��a<�a<S�a<��a< �a<=�a<��a<�a<E�a<u�a<ũa<�a<I�a<��a<��a<�a<4�a<��a<��a<իa<�a<"�a<e�a<��a<��a<ެa<�a<1�a<1�a<c�a<b�a<��a<��a<ŭa<�a<٭a<�a<��a<�a<�a<'�a<C�a<)�a<R�a<.�a<M�a<-�a<9�a<B�a<$�a<<�a<�a<(�a<��a<��a<�a<��a<ϭa<��a<��a<r�a<k�a<F�a<�a<�a<׬a<ݬa<��a<}�a<^�a<!�a<�a<��a<��a<m�a<Y�a<
�a<ߪa<��a<j�a<B�a<�a<ةa<��a<O�a<�a<��a<��a<'�a<��a<��a<c�a<�a<��a<��a<�a<�a<h�a<�a<Ѥa<c�a<#�a<��a<g�a<�a<��a<+�a<��a<y�a<�a<��a<%�a<��a<Q�a<�a<~�a<�a<��a<�a<��a<W�a<�a<{�a<�a<��a<3�a<�a<f�a<��a<��a<�a<՗a<Q�a< �a<��a<(�a<Εa<c�a<�a<��a<W�a<�a<��a<Q�a<�a<��a<;�a<�a<��a<v�a<.�a<אa<��a<Y�a<1�a<ۏa<��a<��a<]�a<6�a<�a<�a<��a<��a<_�a<U�a<P�a<�a<,�a<��a<	�a<��a<�a<�a<ۍa<��a<ݍa<�a<��a<�a<)�a<(�a<c�a<�  �  f�a<��a<��a<Ύa<��a<,�a<g�a<��a<��a<�a<(�a<h�a<��a<�a<4�a<w�a<��a<�a<N�a<��a<��a<W�a<��a<	�a<d�a<��a<$�a<�a<�a<U�a<��a<�a<��a<��a<c�a<՘a<>�a<��a< �a<��a<�a<��a<�a<h�a<לa<N�a<͝a<C�a<��a<#�a<��a<��a<��a<�a<]�a<ܡa<I�a<��a<�a<��a<ޣa<^�a<��a<-�a<��a<�a<<�a<��a<��a<J�a<��a<�a<N�a<��a<�a</�a<|�a<éa<�a<B�a<��a<ͪa<�a<;�a<n�a<��a<Ϋa<
�a<<�a<m�a<��a<��a<ܬa<�a<&�a<2�a<`�a<��a<��a<��a<��a<֭a<ޭa<��a<�a<%�a<&�a<'�a<,�a<4�a<;�a<4�a<E�a<C�a<:�a<.�a<'�a<%�a<$�a<�a< �a<�a<�a<׭a<ȭa<��a<��a<y�a<Y�a<C�a<+�a<�a<�a<ìa<��a<y�a<V�a<&�a<�a<ޫa<��a<m�a<M�a<�a<�a<��a<{�a<J�a<�a<ʩa<~�a<L�a<�a<Ĩa<��a<A�a<�a<��a<\�a<�a<æa<k�a<�a<ťa<t�a<&�a<ͤa<c�a<�a<��a<L�a<��a<��a<:�a<ġa<h�a<�a<��a<!�a<��a<`�a<�a<|�a<�a<��a<(�a<Ӝa<X�a<��a<��a<�a<��a<3�a<Ιa<]�a<��a<��a<&�a<��a<O�a<�a<��a<&�a<��a<\�a< �a<��a<Q�a<�a<��a<F�a<�a<��a<U�a<�a<��a<i�a<,�a<ِa<��a<Z�a<.�a<��a<ďa<��a<V�a<,�a<��a<׎a<��a<��a<y�a<U�a<9�a<%�a<�a<��a<�a<��a<�a<ލa<ލa<�a<��a<��a<��a<�a<%�a<?�a<\�a<�  �  2�a<��a<6�a<I�a<u�a<��a<��a<�a<�a<~�a<��a<�a<*�a<H�a<��a<ؐa<I�a<��a<��a<*�a<e�a<ےa<�a<��a<ړa<Q�a<��a<�a<��a<��a<I�a<��a<�a<��a<�a<`�a<a<d�a<��a<:�a<��a<�a<��a<�a<��a<Ϝa<o�a<Ýa<8�a<��a<�a<��a<�a<��a<��a<h�a<ߡa<C�a<ɢa<�a<��a<ڣa<G�a<��a<�a<��a<Хa<[�a<��a<�a<b�a<��a<�a<=�a<��a<ɨa<�a<^�a<��a<��a<�a<z�a<��a<�a<�a<?�a<��a<��a<��a<�a<1�a<9�a<p�a<��a<��a<�a<�a<(�a<�a<L�a<j�a<`�a<��a<y�a<��a<��a<ͭa<ȭa<��a<�a<��a<!�a<έa<ҭa<ܭa<ʭa<�a<��a<��a<��a<��a<��a<��a<n�a<F�a<��a<�a<!�a<��a<ݬa<ڬa<��a<��a<F�a<M�a<�a<��a<ϫa<��a<��a<+�a<#�a<�a<��a<��a<1�a<�a<��a<ũa<Y�a<3�a<�a<��a<��a<�a<�a<��a<R�a<��a<��a<a�a<�a<�a<i�a<&�a<��a<n�a<;�a<��a<i�a<֢a<��a<�a<��a<U�a<ݠa<��a<�a<֟a<R�a<�a<��a<�a<��a<+�a<Ĝa<E�a<ݛa<{�a<��a<a<'�a<�a<I�a<�a<��a<�a<ȗa<G�a<��a<k�a<�a<��a<@�a<��a<��a<?�a<��a<��a<*�a<��a<��a<�a<��a<b�a<>�a<Րa<��a<M�a<�a<��a<��a<��a<$�a<
�a<�a<��a<��a<8�a<0�a<��a<��a<Սa<��a<��a<x�a<ȍa<h�a<c�a<j�a<Y�a<��a<W�a<g�a<j�a<��a<��a<��a<��a<��a<�  �  �a<��a<6�a<N�a<w�a<��a<Ԏa<�a</�a<z�a<��a<؏a<�a<h�a<��a<�a<0�a<��a<�a<9�a<r�a<�a<&�a<��a<ݓa<A�a<��a<��a<d�a<ɕa<D�a<��a<�a<u�a<�a<f�a<ɘa<9�a<��a<%�a<��a< �a<y�a<�a<{�a<ޜa<d�a<ʝa<U�a<��a<4�a<��a<�a<}�a<�a<i�a<סa<>�a<��a<&�a<��a<��a<W�a<Ѥa<�a<��a<٥a<F�a<��a<�a<7�a<��a<�a<8�a<��a<Ψa<'�a<j�a<��a<�a<'�a<j�a<��a<Ϫa<��a<C�a<x�a<��a<�a<��a<@�a<J�a<��a<��a<��a<Ҭa<�a<�a<2�a<>�a<Q�a<x�a<��a<��a<��a<��a<��a<ȭa<˭a<ޭa<ʭa<ԭa<ϭa<ۭa<֭a<ҭa<ȭa<��a<��a<��a<��a<��a<��a<s�a<R�a<@�a< �a< �a<��a<ެa<¬a<��a<��a<Y�a<I�a< �a<�a<��a<��a<s�a<@�a<
�a<�a<��a<��a<?�a<&�a<ԩa<��a<\�a<#�a<�a<��a<Z�a<�a<ߧa<��a<L�a<�a<��a<g�a<	�a<��a<b�a<�a<��a<S�a<��a<��a<X�a<�a<��a<#�a<աa<d�a<��a<��a<2�a<��a<J�a<�a<}�a<	�a<��a<?�a<לa<g�a<�a<��a<�a<��a<0�a<әa<T�a<�a<u�a<�a<��a<B�a<ؖa<p�a<�a<��a<@�a<�a<��a</�a<œa<j�a<
�a<Ēa<s�a<�a<ۑa<{�a<L�a<�a<��a<r�a<'�a<ڏa<��a<n�a<<�a<��a<Ȏa<��a<��a<Q�a<;�a<�a<�a<ԍa<��a<��a<��a<{�a<h�a<l�a<d�a<b�a<]�a<_�a<p�a<m�a<y�a<��a<��a<��a<ōa<�  �  ܍a<�a<%�a<R�a<��a<��a<ێa<�a<3�a<V�a<��a<ُa<�a<}�a<��a<
�a</�a<��a<Αa<�a<u�a<̒a<1�a<u�a<��a<;�a<��a<�a<d�a<��a</�a<��a<�a<u�a<��a<W�a<ژa</�a<��a<�a<��a<$�a<{�a<�a<_�a<�a<T�a<ŝa<N�a<��a<4�a<��a<�a<|�a<�a<d�a<ʡa<[�a<��a<)�a<q�a<��a<?�a<¤a<�a<v�a<�a</�a<��a<�a<U�a<��a<ڧa<K�a<z�a<ۨa<�a<i�a<��a<�a<4�a<U�a<Īa<۪a<�a<M�a<n�a<��a<ūa<�a<(�a<E�a<q�a<��a<��a<Ҭa<�a<��a<?�a<H�a<T�a<v�a<j�a<��a<��a<��a<��a<έa<խa<ǭa<�a<ɭa<��a<ڭa<ɭa<�a<��a<ϭa<��a<��a<��a<��a<y�a<j�a<��a<7�a<C�a<�a<��a<�a<��a<��a<q�a<]�a<%�a<�a<�a<��a<��a<I�a<]�a<�a<�a<��a<r�a<A�a<�a<ߩa<��a<t�a<�a<�a<��a<Y�a<C�a<˧a<��a<J�a<�a<��a<X�a<�a<��a<v�a<�a<ˤa<v�a<��a<��a<<�a<��a<��a<�a<Ρa<G�a< �a<v�a<2�a<��a<d�a<�a<p�a<&�a<��a<B�a<��a<_�a<՛a<��a<�a<��a<D�a<��a<l�a<�a<��a<2�a<��a<U�a<ϖa<~�a<�a<��a<D�a<�a<��a<�a<�a<u�a<#�a<Βa<i�a<1�a<��a<��a<4�a<�a<��a<S�a<'�a<ڏa<��a<O�a<H�a<�a<ʎa<��a<b�a<V�a<�a<�a<ݍa<ۍa<��a<��a<��a<p�a<��a<l�a<V�a<p�a<N�a<p�a<`�a<|�a<m�a<��a<��a<��a<��a<�  �  �a<�a<)�a<Q�a<��a<��a<ߎa<��a<H�a<v�a<��a<�a<�a<d�a<��a<�a<-�a<��a<͑a<6�a<��a<̒a<6�a<��a<�a<I�a<��a<	�a<j�a<ɕa<2�a<��a<�a<��a<��a<K�a<Ԙa<C�a<��a<*�a<��a<�a<��a<��a<p�a<�a<[�a<۝a<U�a<��a<G�a<��a<�a<��a<��a<e�a<աa<D�a<��a<#�a<��a<�a<b�a<̤a<*�a<��a<�a<>�a<��a<�a<<�a<��a<�a<B�a<��a<ڨa<�a<j�a<��a<�a<2�a<`�a<��a<ժa<�a<A�a<{�a<��a<۫a<�a<*�a<b�a<��a<��a<Ƭa<Ѭa<��a<�a<.�a<=�a<f�a<q�a<��a<��a<��a<��a<ŭa<ɭa<έa<ѭa<ۭa<׭a<Эa<˭a<ݭa<ѭa<έa<Эa<��a<��a<��a<��a<��a<`�a<N�a<E�a<0�a<�a<��a<�a<ɬa<��a<w�a<r�a<E�a<�a<��a<��a<��a<j�a<D�a<�a<�a<��a<��a<\�a<�a<�a<��a<d�a<+�a<�a<��a<_�a<�a<ͧa<��a<C�a<��a<��a<M�a<�a<��a<j�a<�a<��a<U�a<�a<��a<M�a<�a<��a<4�a<աa<b�a<�a<��a<,�a<��a<Q�a<�a<{�a<�a<��a<;�a<ɜa<r�a<��a<��a<�a<��a<7�a<˙a<R�a<�a<z�a<�a<��a<L�a<�a<}�a<�a<��a<P�a<�a<��a<%�a<Óa<p�a<�a<a<v�a<�a<֑a<��a<6�a<��a<��a<[�a<,�a<ُa<��a<l�a<7�a<��a<ݎa<��a<��a<g�a<'�a<�a<��a<Սa<��a<��a<��a<~�a<j�a<\�a<j�a<`�a<d�a<q�a<T�a<��a<��a<��a<��a<��a<a<�  �  ��a<��a<A�a<Q�a<q�a<��a<Ďa<�a<$�a<m�a<��a<�a< �a<^�a<��a<�a<A�a<��a<ؑa<'�a<m�a<Вa<!�a<��a<̓a<Q�a<��a<�a<|�a<˕a<[�a<��a<�a<��a<�a<[�a<Ęa<J�a<��a<<�a<��a<�a<��a<�a<��a<Ӝa<_�a<ȝa<:�a<��a<�a<��a<�a<��a<�a<l�a<ޡa<:�a<��a<�a<��a<�a<W�a<��a<�a<��a<ɥa<V�a<��a<��a<L�a<��a<�a<%�a<��a<Ϩa<�a<`�a<��a<�a<�a<��a<��a<�a<�a<J�a<��a<��a<�a<��a<&�a<G�a<r�a<��a<��a<�a<�a<!�a<.�a<E�a<f�a<i�a<��a<��a<��a<��a<��a<ĭa<ɭa<�a<ƭa<�a<ӭa<�a<�a<��a<խa<��a<��a<��a<��a<��a<��a<��a<Q�a<X�a<�a<+�a<��a<جa<ʬa<��a<��a<N�a<<�a<�a<��a<ūa<��a<~�a<:�a<�a<�a<��a<}�a<9�a<�a<Ωa<��a<K�a<3�a<�a<��a<q�a<�a<��a<��a<B�a<�a<��a<\�a<�a<ƥa<M�a<(�a<Ƥa<b�a<�a<��a<f�a<ڢa<��a<!�a<��a<`�a<�a<��a<%�a<ȟa<N�a<�a<��a<�a<��a<2�a<Ҝa<L�a<�a<x�a<�a<��a< �a<�a<R�a<��a<��a<�a<ʗa</�a<�a<r�a<�a<��a<L�a<�a<y�a<J�a<ɓa<��a<�a<˒a<��a<�a<�a<y�a<3�a<�a<��a<h�a<$�a<�a<��a<z�a<8�a<�a<ݎa<��a<~�a<B�a<1�a<��a<�a<Ѝa<��a<��a<�a<��a<m�a<��a<o�a<O�a<k�a<W�a<g�a<j�a<��a<��a<��a<Ѝa<ōa<�  �  �a<�a<&�a<E�a<��a<��a<Ǝa<�a<8�a<o�a<��a<Џa<+�a<k�a<��a<��a<A�a<p�a<Ցa<.�a<{�a<ߒa<!�a<��a<�a<<�a<��a<�a<s�a<ѕa<3�a<��a<!�a<��a<�a<m�a<Řa<M�a<��a<�a<��a<�a<��a<��a<n�a<ޜa<a�a<ϝa<?�a<��a<1�a<��a<	�a<��a<
�a<d�a<ϡa<Y�a<��a<�a<��a<�a<\�a<��a<�a<��a<ܥa<=�a<��a<�a<I�a<��a<ݧa<<�a<��a<ͨa<%�a<_�a<��a<��a<�a<\�a<��a<�a<�a<D�a<t�a<��a<ݫa<��a<2�a<S�a<|�a<��a<��a<�a<
�a<��a<4�a<R�a<O�a<n�a<��a<��a<��a<��a<��a<ԭa<ía<έa<׭a<�a<٭a<ӭa<��a<�a<ҭa<��a<ͭa<��a<��a<��a<g�a<j�a<Y�a<N�a<1�a<�a<�a<�a<Ȭa<��a<��a<b�a<>�a<�a<ܫa<Ыa<��a<W�a<P�a<�a<ͪa<��a<��a<H�a<�a<Ωa<��a<l�a<�a<ߨa<��a<h�a<�a<Χa<�a<U�a<��a<��a<o�a<�a<ɥa<m�a<��a<��a<c�a<�a<��a<K�a<�a<��a<(�a<��a<f�a<��a<��a<�a<��a<g�a<�a<u�a<%�a<��a<(�a<ʜa<]�a<�a<{�a<�a<��a<3�a<ʙa<_�a<�a<��a<�a<��a<F�a<�a<p�a<�a<��a<H�a<��a<�a<!�a<Γa<z�a< �a<Œa<n�a<%�a<ؑa<{�a<?�a<�a<��a<d�a<�a<�a<��a<X�a<=�a<�a<Ǝa<��a<�a<[�a<=�a<�a<�a<��a<��a<��a<��a<��a<s�a<e�a<K�a<r�a<g�a<R�a<}�a<d�a<��a<��a<��a<��a<̍a<�  �  �a<�a<%�a<R�a<w�a<��a<ߎa<��a<<�a<r�a<��a<ۏa<�a<l�a<��a<��a<&�a<��a<ؑa<2�a<|�a<̒a<8�a<��a<�a<>�a<��a<�a<b�a<��a<:�a<��a<�a<r�a<�a<\�a<͘a<)�a<��a<"�a<��a<�a<|�a<�a<c�a<�a<O�a<۝a<F�a<��a<=�a<��a< �a<y�a<��a<n�a<ܡa<F�a<��a<'�a<��a<��a<N�a<��a</�a<u�a<�a<1�a<��a<�a<=�a<��a<�a<B�a<u�a<Ҩa<�a<g�a<��a<۩a<4�a<c�a<��a<Ϊa<�a<M�a<o�a<��a<̫a<�a<$�a<O�a<��a<��a<Ĭa<Ǭa<��a<�a<6�a<:�a<T�a<}�a<��a<��a<��a<��a<��a<­a<խa<ͭa<�a<ҭa<ڭa<�a<׭a<ҭa<��a<ǭa<��a<��a<��a<��a<��a<u�a<^�a<=�a<<�a<�a<��a<ެa<��a<��a<y�a<f�a<A�a<�a<�a<��a<��a<r�a<G�a< �a<�a<��a<��a<H�a<�a<�a<��a<m�a< �a<�a<��a<X�a<*�a<էa<��a<:�a<�a<��a<]�a<�a<��a<m�a<�a<äa<Z�a<��a<��a<@�a<��a<��a<4�a<ǡa<T�a<�a<��a<4�a<��a<R�a<�a<��a<�a<��a<@�a<Ɯa<j�a<�a<~�a<!�a<��a<D�a<��a<k�a<�a<{�a<$�a<��a<L�a<ʖa<u�a<�a<��a<C�a<۔a<��a<(�a<ޓa<i�a<!�a<Βa<i�a<,�a<Ǒa<��a<0�a<�a<��a<d�a<*�a<Ϗa<��a<q�a<?�a<��a<ˎa<��a<|�a<_�a<&�a<�a<�a<΍a<��a<��a<��a<y�a<s�a<r�a<e�a<a�a<K�a<g�a<i�a<y�a<m�a<��a<��a<��a<ҍa<�  �  ��a<��a<3�a<]�a<m�a<��a<Ԏa<
�a<3�a<h�a<��a<�a<'�a<Z�a<��a<�a<E�a<��a<��a<$�a<~�a<ےa<,�a<��a<ۓa<P�a<��a< �a<w�a<ەa<?�a<��a<�a<��a<�a<F�a<ݘa<F�a<��a<%�a<��a<�a<��a<�a<t�a<�a<Y�a<Нa<F�a<��a<.�a<��a<�a<��a<��a<h�a<ޡa<A�a<��a<�a<}�a<�a<\�a<��a<#�a<��a<ޥa<B�a<��a<�a<I�a<��a<�a<)�a<��a<�a<�a<_�a<��a<�a<�a<f�a<��a<�a<�a<E�a<��a<��a<ԫa<�a<.�a<U�a<v�a<��a<Ǭa<�a<�a<+�a<)�a<L�a<o�a<_�a<}�a<��a<��a<��a<��a<��a<حa<ݭa<ʭa<�a<حa<ޭa<ԭa<��a<ѭa<έa<��a<��a<��a<|�a<�a<q�a<[�a<R�a<!�a<�a<�a<Ԭa<��a<��a<��a<]�a<7�a<��a< �a<˫a<��a<��a<4�a<�a<��a<��a<z�a<J�a<�a<کa<��a<Z�a<2�a<�a<��a<m�a<%�a<ڧa<��a<7�a<�a<��a<H�a<�a<¥a<P�a<�a<��a<b�a<	�a<��a<Q�a<�a<��a<*�a<ơa<e�a<��a<��a<!�a<͟a<R�a<�a<��a<�a<��a<6�a<��a<^�a<�a<��a<�a<��a<5�a<Ιa<X�a<�a<��a<�a<��a<3�a<�a<��a<�a<��a<Y�a<�a<�a<+�a<ӓa<}�a<�a<ƒa<|�a<�a<ϑa<��a<;�a<�a<��a<O�a<-�a<�a<��a<��a<2�a<
�a<�a<��a<t�a<Q�a<6�a<�a<�a<ɍa<Ía<��a<��a<��a<r�a<o�a<a�a<I�a<f�a<n�a<M�a<z�a<��a<y�a<��a<��a<΍a<�  �  �a<��a<6�a<D�a<}�a<��a<a<�a<,�a<��a<��a<ޏa<*�a<]�a<��a<�a<H�a<s�a<�a<=�a<x�a<�a<�a<��a<ݓa<C�a<��a<��a<n�a<a<?�a<��a<�a<{�a<�a<d�a<��a<F�a<��a<)�a<��a<�a<|�a<�a<}�a<˜a<n�a<ѝa<F�a<Ğa<+�a<a<�a<��a<��a<h�a<ڡa<E�a<��a<
�a<��a<��a<a�a<Ƥa<�a<��a<ȥa<H�a<��a<�a<C�a<��a<�a<5�a<��a<Ũa<#�a<c�a<��a<�a<"�a<k�a<��a<۪a<�a<@�a<z�a<��a<�a<�a<9�a<R�a<��a<��a<��a<�a<�a<�a<*�a<P�a<[�a<n�a<��a<��a<��a<��a<̭a<Эa<��a<�a<̭a<׭a<ȭa<׭a<խa<ڭa<έa<��a<ƭa<��a<��a<��a<{�a<m�a<I�a<F�a<"�a<!�a<�a<�a<׬a<��a<��a<V�a<Y�a<�a<�a<ϫa<��a<p�a<8�a<"�a<Ъa<��a<��a<D�a<#�a<ʩa<��a<\�a<%�a<�a<��a<c�a<�a<ڧa<��a<L�a<��a<��a<e�a< �a<¥a<c�a<�a<��a<X�a<��a<��a<Z�a<Ӣa<��a<*�a<ơa<j�a<��a<��a<�a<a<W�a<�a<��a<�a<��a<#�a<�a<`�a<��a<��a<�a<��a<�a<ՙa<R�a<�a<��a<
�a<��a<?�a<�a<h�a<�a<��a<E�a<�a<��a<0�a<��a<v�a<�a<��a<u�a<�a<�a<u�a<F�a<�a<��a<z�a<�a<�a<��a<n�a<3�a<�a<юa<��a<��a<L�a<@�a<�a<��a<܍a<��a<��a<��a<~�a<b�a<i�a<c�a<i�a<c�a<Z�a<v�a<i�a<~�a<��a<��a<��a<��a<�  �  ݍa<�a<2�a<W�a<z�a<��a<Ҏa<�a<+�a<_�a<��a<�a<%�a<u�a<��a<��a<@�a<��a<ߑa<�a<t�a<ђa</�a<��a<�a<F�a<��a<�a<f�a<�a<>�a<��a<�a<t�a<�a<X�a<̘a<4�a<��a<�a<��a<�a<��a<�a<s�a<�a<[�a<ȝa<C�a<��a<"�a<��a<�a<��a< �a<m�a<աa<N�a<��a<(�a<��a<�a<P�a<��a<�a<��a<�a<?�a<��a<��a<Q�a<��a<�a<>�a<��a<Ҩa<�a<]�a<��a<�a<*�a<g�a<��a<تa<!�a<Q�a<y�a<��a<٫a<�a<*�a<I�a<g�a<��a<��a<�a<�a<�a<?�a<M�a<]�a<}�a<{�a<��a<��a<��a<��a<ʭa<Эa<ۭa<�a<ϭa<�a<�a<̭a<ڭa<��a<­a<��a<��a<��a<��a<z�a<y�a<l�a<8�a<:�a<�a<�a<�a<��a<��a<��a<U�a<.�a<�a<�a<ɫa<��a<]�a<P�a<�a<�a<��a<q�a<A�a<�a<ݩa<��a<f�a<(�a<�a<��a<[�a<1�a<٧a<��a<I�a<�a<��a<Z�a<�a<��a<l�a<�a<Ȥa<n�a<�a<��a<P�a<�a<��a<!�a<áa<Z�a<�a<��a<3�a<��a<]�a<�a<{�a<�a<��a<A�a<ʜa<M�a<�a<��a<�a<��a<7�a<̙a<f�a<��a<��a<,�a<��a<H�a<Ֆa<u�a<�a<��a<C�a<�a<��a<,�a<�a<s�a<-�a<Ғa<t�a<"�a<ӑa<��a<7�a<�a<��a<l�a<%�a<�a<��a<^�a<H�a<
�a<Ԏa<��a<r�a<J�a<-�a<�a<�a<֍a<��a<��a<��a<v�a<��a<w�a<Z�a<i�a<Q�a<b�a<`�a<p�a<n�a<��a<��a<��a<��a<�  �  ܍a<�a<�a<b�a<v�a<��a<�a<�a<^�a<e�a<��a<��a<�a<o�a<��a< �a<+�a<��a<ɑa<.�a<��a<Ēa<D�a<y�a<�a<H�a<��a<�a<V�a<וa< �a<��a<�a<��a<��a<?�a<�a<4�a<��a<�a<��a<��a<��a<��a<_�a<��a<P�a<ٝa<I�a<��a<N�a<��a<#�a<��a<��a<m�a<ءa<L�a<��a<.�a<v�a<�a<d�a<��a<.�a<u�a<�a</�a<��a<�a</�a<��a<էa<B�a<}�a<�a<�a<a�a<��a<ݩa<0�a<J�a<��a<��a<�a<;�a<u�a<��a<ǫa<�a< �a<m�a<��a<��a<ͬa<ͬa<
�a<�a<:�a<=�a<e�a<v�a<z�a<��a<��a<��a<��a<��a<߭a<��a<ޭa<Эa<ӭa<ʭa<ѭa<̭a<��a<ܭa<��a<ǭa<��a<��a<��a<Y�a<V�a<7�a<8�a<�a<�a<ݬa<��a<��a<t�a<��a<5�a<�a<��a<��a<��a<j�a<S�a<�a<��a<��a<��a<i�a<�a<�a<��a<m�a<*�a<بa<��a<K�a<!�a<��a<��a<9�a<��a<��a<A�a<$�a<��a<l�a<��a<��a<O�a<�a<��a<<�a<��a<��a<3�a<ɡa<e�a<�a<��a<7�a<��a<U�a<�a<~�a<�a<��a<G�a<��a<x�a<��a<��a< �a<��a<E�a<��a<W�a<�a<m�a<�a<��a<L�a<Җa<��a<��a<��a<S�a<ݔa<��a<�a<֓a<[�a<&�a<��a<p�a<,�a<a<��a<-�a<	�a<��a<V�a<3�a<Տa<��a<j�a<C�a<��a<܎a<��a<r�a<{�a<%�a<�a<�a<ʍa<ˍa<��a<��a<w�a<l�a<[�a<_�a<[�a<S�a<|�a<?�a<��a<u�a<��a<��a<��a<ʍa<�  �  ��a<�a<-�a<M�a<v�a<��a<a<��a<.�a<t�a<��a<�a<�a<`�a<��a<�a<9�a<��a<ؑa<)�a<q�a<͒a<�a<��a<��a<G�a<��a<�a<v�a<ҕa<I�a<��a<�a<s�a<�a<Y�a<Øa<3�a<��a<2�a<��a<�a<��a<�a<x�a<ۜa<\�a<˝a<4�a<��a<#�a<��a<�a<��a<�a<s�a<�a<A�a<��a<�a<��a<�a<K�a<��a<�a<��a<إa<F�a<��a<�a<B�a<��a<��a<A�a<{�a<ʨa<�a<b�a<��a<ީa</�a<r�a<��a<�a<�a<A�a<�a<��a<�a<��a<"�a<F�a<t�a<��a<��a<٬a<��a<�a</�a<?�a<e�a<u�a<��a<��a<��a<��a<ía<ía<ȭa<ܭa<ӭa<�a<ϭa<�a<�a<έa<��a<��a<��a<��a<��a<��a<��a<|�a<S�a<W�a<0�a<�a<��a<ެa<ͬa<��a<}�a<W�a<C�a<�a<��a<��a<��a<z�a<A�a<�a<�a<��a<�a<=�a<�a<̩a<��a<_�a<)�a<�a<��a<k�a<�a<�a<��a<9�a<�a<��a<Z�a<�a<��a<k�a<�a<ɤa<Z�a<�a<��a<U�a<�a<��a<%�a<��a<S�a<�a<��a<(�a<şa<N�a<��a<��a<�a<��a<5�a<̜a<S�a<�a<q�a<�a<��a<.�a<әa<S�a<�a<��a<%�a<��a<K�a<Жa<m�a<�a<��a<=�a<ݔa<��a<7�a<ӓa<{�a<*�a<a<z�a<�a<ݑa<w�a<.�a<�a<��a<f�a< �a<�a<��a<y�a<8�a<��a<܎a<��a<��a<J�a<)�a<��a<��a<ύa<��a<��a<��a<��a<i�a<x�a<p�a<]�a<S�a<a�a<k�a<t�a<s�a<��a<��a<Ía<Ǎa<�  �  �a<�a<G�a<J�a<v�a<��a<a<K�a<�a<p�a<��a<�a<7�a<_�a<��a<�a<^�a<��a<�a<�a<y�a<�a<�a<��a<ғa<K�a<��a<��a<k�a<��a<L�a<��a<"�a<�a<ݗa<k�a<��a<O�a<��a<�a<��a<��a<��a<ٛa<��a<؜a<s�a<ŝa<Y�a<�a<�a<��a<�a<��a<�a<e�a<סa<=�a<Ңa<�a<��a<ߣa<|�a<�a<�a<��a<ҥa<]�a<{�a<�a<0�a<��a<�a<.�a<��a<̨a<%�a<\�a<��a<��a<�a<l�a<��a<Ԫa<�a<A�a<��a<��a<�a<�a<h�a<Z�a<h�a<��a<��a<�a<�a<�a<-�a<Q�a<h�a<o�a<��a<|�a<�a<��a<��a<έa<ŭa<��a<��a<�a<ía<߭a<��a<ѭa<׭a<��a<ͭa<��a<��a<��a<i�a<}�a<B�a<I�a<�a<1�a<��a<ݬa<ʬa<��a<ˬa<H�a<?�a<�a<�a<ܫa<��a<r�a<6�a<8�a<ުa<��a<u�a<E�a<Y�a<��a<��a<Q�a<-�a<�a<��a<a�a<�a<�a<�a<V�a<��a<��a<m�a<��a<˥a<Z�a<��a<��a<F�a<	�a<��a<p�a<�a<��a<�a<١a<��a<�a<��a<!�a<ןa<J�a<�a<}�a<�a<ĝa<7�a<�a<J�a<�a<��a<�a<Úa<)�a<�a<@�a<�a<n�a<�a<��a<8�a<�a<o�a<�a<��a<G�a<��a<{�a<1�a<��a<o�a<�a<a<��a<�a<�a<k�a<t�a<��a<��a<x�a<#�a<
�a<��a<s�a<6�a<�a<ߎa<��a<��a<;�a<y�a<	�a<�a<ڍa<��a<ȍa<m�a<��a<]�a<p�a<H�a<`�a<m�a<G�a<}�a<R�a<��a<��a<��a<ča<��a<�  �  ��a<�a<-�a<M�a<v�a<��a<a<��a<.�a<t�a<��a<�a<�a<`�a<��a<�a<9�a<��a<ؑa<)�a<q�a<͒a<�a<��a<��a<G�a<��a<�a<v�a<ҕa<I�a<��a<�a<s�a<�a<Y�a<Øa<3�a<��a<2�a<��a<�a<��a<�a<x�a<ۜa<\�a<˝a<4�a<��a<#�a<��a<�a<��a<�a<s�a<�a<A�a<��a<�a<��a<�a<K�a<��a<�a<��a<إa<F�a<��a<�a<B�a<��a<��a<A�a<{�a<ʨa<�a<b�a<��a<ީa</�a<r�a<��a<�a<�a<A�a<�a<��a<�a<��a<"�a<F�a<t�a<��a<��a<٬a<��a<�a</�a<?�a<e�a<u�a<��a<��a<��a<��a<ía<ía<ȭa<ܭa<ӭa<�a<ϭa<�a<�a<έa<��a<��a<��a<��a<��a<��a<��a<|�a<S�a<W�a<0�a<�a<��a<ެa<ͬa<��a<}�a<W�a<C�a<�a<��a<��a<��a<z�a<A�a<�a<�a<��a<�a<=�a<�a<̩a<��a<_�a<)�a<�a<��a<k�a<�a<�a<��a<9�a<�a<��a<Z�a<�a<��a<k�a<�a<ɤa<Z�a<�a<��a<U�a<�a<��a<%�a<��a<S�a<�a<��a<(�a<şa<N�a<��a<��a<�a<��a<5�a<̜a<S�a<�a<q�a<�a<��a<.�a<әa<S�a<�a<��a<%�a<��a<K�a<Жa<m�a<�a<��a<=�a<ݔa<��a<7�a<ӓa<{�a<*�a<a<z�a<�a<ݑa<w�a<.�a<�a<��a<f�a< �a<�a<��a<y�a<8�a<��a<܎a<��a<��a<J�a<)�a<��a<��a<ύa<��a<��a<��a<��a<i�a<x�a<p�a<]�a<S�a<a�a<k�a<t�a<s�a<��a<��a<Ía<Ǎa<�  �  ܍a<�a<�a<b�a<v�a<��a<�a<�a<^�a<e�a<��a<��a<�a<o�a<��a< �a<+�a<��a<ɑa<.�a<��a<Ēa<D�a<y�a<�a<H�a<��a<�a<V�a<וa< �a<��a<�a<��a<��a<?�a<�a<4�a<��a<�a<��a<��a<��a<��a<_�a<��a<P�a<ٝa<I�a<��a<N�a<��a<#�a<��a<��a<m�a<ءa<L�a<��a<.�a<v�a<�a<d�a<��a<.�a<u�a<�a</�a<��a<�a</�a<��a<էa<B�a<}�a<�a<�a<a�a<��a<ݩa<0�a<J�a<��a<��a<�a<;�a<u�a<��a<ǫa<�a< �a<m�a<��a<��a<ͬa<ͬa<
�a<�a<:�a<=�a<e�a<v�a<z�a<��a<��a<��a<��a<��a<߭a<��a<ޭa<Эa<ӭa<ʭa<ѭa<̭a<��a<ܭa<��a<ǭa<��a<��a<��a<Y�a<V�a<7�a<8�a<�a<�a<ݬa<��a<��a<t�a<��a<5�a<�a<��a<��a<��a<j�a<S�a<�a<��a<��a<��a<i�a<�a<�a<��a<m�a<*�a<بa<��a<K�a<!�a<��a<��a<9�a<��a<��a<A�a<$�a<��a<l�a<��a<��a<O�a<�a<��a<<�a<��a<��a<3�a<ɡa<e�a<�a<��a<7�a<��a<U�a<�a<~�a<�a<��a<G�a<��a<x�a<��a<��a< �a<��a<E�a<��a<W�a<�a<m�a<�a<��a<L�a<Җa<��a<��a<��a<S�a<ݔa<��a<�a<֓a<[�a<&�a<��a<p�a<,�a<a<��a<-�a<	�a<��a<V�a<3�a<Տa<��a<j�a<C�a<��a<܎a<��a<r�a<{�a<%�a<�a<�a<ʍa<ˍa<��a<��a<w�a<l�a<[�a<_�a<[�a<S�a<|�a<?�a<��a<u�a<��a<��a<��a<ʍa<�  �  ݍa<�a<2�a<W�a<z�a<��a<Ҏa<�a<+�a<_�a<��a<�a<%�a<u�a<��a<��a<@�a<��a<ߑa<�a<t�a<ђa</�a<��a<�a<F�a<��a<�a<f�a<�a<>�a<��a<�a<t�a<�a<X�a<̘a<4�a<��a<�a<��a<�a<��a<�a<s�a<�a<[�a<ȝa<C�a<��a<"�a<��a<�a<��a< �a<m�a<աa<N�a<��a<(�a<��a<�a<P�a<��a<�a<��a<�a<?�a<��a<��a<Q�a<��a<�a<>�a<��a<Ҩa<�a<]�a<��a<�a<*�a<g�a<��a<تa<!�a<Q�a<y�a<��a<٫a<�a<*�a<I�a<g�a<��a<��a<�a<�a<�a<?�a<M�a<]�a<}�a<{�a<��a<��a<��a<��a<ʭa<Эa<ۭa<�a<ϭa<�a<�a<̭a<ڭa<��a<­a<��a<��a<��a<��a<z�a<y�a<l�a<8�a<:�a<�a<�a<�a<��a<��a<��a<U�a<.�a<�a<�a<ɫa<��a<]�a<P�a<�a<�a<��a<q�a<A�a<�a<ݩa<��a<f�a<(�a<�a<��a<[�a<1�a<٧a<��a<I�a<�a<��a<Z�a<�a<��a<l�a<�a<Ȥa<n�a<�a<��a<P�a<�a<��a<!�a<áa<Z�a<�a<��a<3�a<��a<]�a<�a<{�a<�a<��a<A�a<ʜa<M�a<�a<��a<�a<��a<7�a<̙a<f�a<��a<��a<,�a<��a<H�a<Ֆa<u�a<�a<��a<C�a<�a<��a<,�a<�a<s�a<-�a<Ғa<t�a<"�a<ӑa<��a<7�a<�a<��a<l�a<%�a<�a<��a<^�a<H�a<
�a<Ԏa<��a<r�a<J�a<-�a<�a<�a<֍a<��a<��a<��a<v�a<��a<w�a<Z�a<i�a<Q�a<b�a<`�a<p�a<n�a<��a<��a<��a<��a<�  �  �a<��a<6�a<D�a<}�a<��a<a<�a<,�a<��a<��a<ޏa<*�a<]�a<��a<�a<H�a<s�a<�a<=�a<x�a<�a<�a<��a<ݓa<C�a<��a<��a<n�a<a<?�a<��a<�a<{�a<�a<d�a<��a<F�a<��a<)�a<��a<�a<|�a<�a<}�a<˜a<n�a<ѝa<F�a<Ğa<+�a<a<�a<��a<��a<h�a<ڡa<E�a<��a<
�a<��a<��a<a�a<Ƥa<�a<��a<ȥa<H�a<��a<�a<C�a<��a<�a<5�a<��a<Ũa<#�a<c�a<��a<�a<"�a<k�a<��a<۪a<�a<@�a<z�a<��a<�a<�a<9�a<R�a<��a<��a<��a<�a<�a<�a<*�a<P�a<[�a<n�a<��a<��a<��a<��a<̭a<Эa<��a<�a<̭a<׭a<ȭa<׭a<խa<ڭa<έa<��a<ƭa<��a<��a<��a<{�a<m�a<I�a<F�a<"�a<!�a<�a<�a<׬a<��a<��a<V�a<Y�a<�a<�a<ϫa<��a<p�a<8�a<"�a<Ъa<��a<��a<D�a<#�a<ʩa<��a<\�a<%�a<�a<��a<c�a<�a<ڧa<��a<L�a<��a<��a<e�a< �a<¥a<c�a<�a<��a<X�a<��a<��a<Z�a<Ӣa<��a<*�a<ơa<j�a<��a<��a<�a<a<W�a<�a<��a<�a<��a<#�a<�a<`�a<��a<��a<�a<��a<�a<ՙa<R�a<�a<��a<
�a<��a<?�a<�a<h�a<�a<��a<E�a<�a<��a<0�a<��a<v�a<�a<��a<u�a<�a<�a<u�a<F�a<�a<��a<z�a<�a<�a<��a<n�a<3�a<�a<юa<��a<��a<L�a<@�a<�a<��a<܍a<��a<��a<��a<~�a<b�a<i�a<c�a<i�a<c�a<Z�a<v�a<i�a<~�a<��a<��a<��a<��a<�  �  ��a<��a<3�a<]�a<m�a<��a<Ԏa<
�a<3�a<h�a<��a<�a<'�a<Z�a<��a<�a<E�a<��a<��a<$�a<~�a<ےa<,�a<��a<ۓa<P�a<��a< �a<w�a<ەa<?�a<��a<�a<��a<�a<F�a<ݘa<F�a<��a<%�a<��a<�a<��a<�a<t�a<�a<Y�a<Нa<F�a<��a<.�a<��a<�a<��a<��a<h�a<ޡa<A�a<��a<�a<}�a<�a<\�a<��a<#�a<��a<ޥa<B�a<��a<�a<I�a<��a<�a<)�a<��a<�a<�a<_�a<��a<�a<�a<f�a<��a<�a<�a<E�a<��a<��a<ԫa<�a<.�a<U�a<v�a<��a<Ǭa<�a<�a<+�a<)�a<L�a<o�a<_�a<}�a<��a<��a<��a<��a<��a<حa<ݭa<ʭa<�a<حa<ޭa<ԭa<��a<ѭa<έa<��a<��a<��a<|�a<�a<q�a<[�a<R�a<!�a<�a<�a<Ԭa<��a<��a<��a<]�a<7�a<��a< �a<˫a<��a<��a<4�a<�a<��a<��a<z�a<J�a<�a<کa<��a<Z�a<2�a<�a<��a<m�a<%�a<ڧa<��a<7�a<�a<��a<H�a<�a<¥a<P�a<�a<��a<b�a<	�a<��a<Q�a<�a<��a<*�a<ơa<e�a<��a<��a<!�a<͟a<R�a<�a<��a<�a<��a<6�a<��a<^�a<�a<��a<�a<��a<5�a<Ιa<X�a<�a<��a<�a<��a<3�a<�a<��a<�a<��a<Y�a<�a<�a<+�a<ӓa<}�a<�a<ƒa<|�a<�a<ϑa<��a<;�a<�a<��a<O�a<-�a<�a<��a<��a<2�a<
�a<�a<��a<t�a<Q�a<6�a<�a<�a<ɍa<Ía<��a<��a<��a<r�a<o�a<a�a<I�a<f�a<n�a<M�a<z�a<��a<y�a<��a<��a<΍a<�  �  �a<�a<%�a<R�a<w�a<��a<ߎa<��a<<�a<r�a<��a<ۏa<�a<l�a<��a<��a<&�a<��a<ؑa<2�a<|�a<̒a<8�a<��a<�a<>�a<��a<�a<b�a<��a<:�a<��a<�a<r�a<�a<\�a<͘a<)�a<��a<"�a<��a<�a<|�a<�a<c�a<�a<O�a<۝a<F�a<��a<=�a<��a< �a<y�a<��a<n�a<ܡa<F�a<��a<'�a<��a<��a<N�a<��a</�a<u�a<�a<1�a<��a<�a<=�a<��a<�a<B�a<u�a<Ҩa<�a<g�a<��a<۩a<4�a<c�a<��a<Ϊa<�a<M�a<o�a<��a<̫a<�a<$�a<O�a<��a<��a<Ĭa<Ǭa<��a<�a<6�a<:�a<T�a<}�a<��a<��a<��a<��a<��a<­a<խa<ͭa<�a<ҭa<ڭa<�a<׭a<ҭa<��a<ǭa<��a<��a<��a<��a<��a<u�a<^�a<=�a<<�a<�a<��a<ެa<��a<��a<y�a<f�a<A�a<�a<�a<��a<��a<r�a<G�a< �a<�a<��a<��a<H�a<�a<�a<��a<m�a< �a<�a<��a<X�a<*�a<էa<��a<:�a<�a<��a<]�a<�a<��a<m�a<�a<äa<Z�a<��a<��a<@�a<��a<��a<4�a<ǡa<T�a<�a<��a<4�a<��a<R�a<�a<��a<�a<��a<@�a<Ɯa<j�a<�a<~�a<!�a<��a<D�a<��a<k�a<�a<{�a<$�a<��a<L�a<ʖa<u�a<�a<��a<C�a<۔a<��a<(�a<ޓa<i�a<!�a<Βa<i�a<,�a<Ǒa<��a<0�a<�a<��a<d�a<*�a<Ϗa<��a<q�a<?�a<��a<ˎa<��a<|�a<_�a<&�a<�a<�a<΍a<��a<��a<��a<y�a<s�a<r�a<e�a<a�a<K�a<g�a<i�a<y�a<m�a<��a<��a<��a<ҍa<�  �  �a<�a<&�a<E�a<��a<��a<Ǝa<�a<8�a<o�a<��a<Џa<+�a<k�a<��a<��a<A�a<p�a<Ցa<.�a<{�a<ߒa<!�a<��a<�a<<�a<��a<�a<s�a<ѕa<3�a<��a<!�a<��a<�a<m�a<Řa<M�a<��a<�a<��a<�a<��a<��a<n�a<ޜa<a�a<ϝa<?�a<��a<1�a<��a<	�a<��a<
�a<d�a<ϡa<Y�a<��a<�a<��a<�a<\�a<��a<�a<��a<ܥa<=�a<��a<�a<I�a<��a<ݧa<<�a<��a<ͨa<%�a<_�a<��a<��a<�a<\�a<��a<�a<�a<D�a<t�a<��a<ݫa<��a<2�a<S�a<|�a<��a<��a<�a<
�a<��a<4�a<R�a<O�a<n�a<��a<��a<��a<��a<��a<ԭa<ía<έa<׭a<�a<٭a<ӭa<��a<�a<ҭa<��a<ͭa<��a<��a<��a<g�a<j�a<Y�a<N�a<1�a<�a<�a<�a<Ȭa<��a<��a<b�a<>�a<�a<ܫa<Ыa<��a<W�a<P�a<�a<ͪa<��a<��a<H�a<�a<Ωa<��a<l�a<�a<ߨa<��a<h�a<�a<Χa<�a<U�a<��a<��a<o�a<�a<ɥa<m�a<��a<��a<c�a<�a<��a<K�a<�a<��a<(�a<��a<f�a<��a<��a<�a<��a<g�a<�a<u�a<%�a<��a<(�a<ʜa<]�a<�a<{�a<�a<��a<3�a<ʙa<_�a<�a<��a<�a<��a<F�a<�a<p�a<�a<��a<H�a<��a<�a<!�a<Γa<z�a< �a<Œa<n�a<%�a<ؑa<{�a<?�a<�a<��a<d�a<�a<�a<��a<X�a<=�a<�a<Ǝa<��a<�a<[�a<=�a<�a<�a<��a<��a<��a<��a<��a<s�a<e�a<K�a<r�a<g�a<R�a<}�a<d�a<��a<��a<��a<��a<̍a<�  �  ��a<��a<A�a<Q�a<q�a<��a<Ďa<�a<$�a<m�a<��a<�a< �a<^�a<��a<�a<A�a<��a<ؑa<'�a<m�a<Вa<!�a<��a<̓a<Q�a<��a<�a<|�a<˕a<[�a<��a<�a<��a<�a<[�a<Ęa<J�a<��a<<�a<��a<�a<��a<�a<��a<Ӝa<_�a<ȝa<:�a<��a<�a<��a<�a<��a<�a<l�a<ޡa<:�a<��a<�a<��a<�a<W�a<��a<�a<��a<ɥa<V�a<��a<��a<L�a<��a<�a<%�a<��a<Ϩa<�a<`�a<��a<�a<�a<��a<��a<�a<�a<J�a<��a<��a<�a<��a<&�a<G�a<r�a<��a<��a<�a<�a<!�a<.�a<E�a<f�a<i�a<��a<��a<��a<��a<��a<ĭa<ɭa<�a<ƭa<�a<ӭa<�a<�a<��a<խa<��a<��a<��a<��a<��a<��a<��a<Q�a<X�a<�a<+�a<��a<جa<ʬa<��a<��a<N�a<<�a<�a<��a<ūa<��a<~�a<:�a<�a<�a<��a<}�a<9�a<�a<Ωa<��a<K�a<3�a<�a<��a<q�a<�a<��a<��a<B�a<�a<��a<\�a<�a<ƥa<M�a<(�a<Ƥa<b�a<�a<��a<f�a<ڢa<��a<!�a<��a<`�a<�a<��a<%�a<ȟa<N�a<�a<��a<�a<��a<2�a<Ҝa<L�a<�a<x�a<�a<��a< �a<�a<R�a<��a<��a<�a<ʗa</�a<�a<r�a<�a<��a<L�a<�a<y�a<J�a<ɓa<��a<�a<˒a<��a<�a<�a<y�a<3�a<�a<��a<h�a<$�a<�a<��a<z�a<8�a<�a<ݎa<��a<~�a<B�a<1�a<��a<�a<Ѝa<��a<��a<�a<��a<m�a<��a<o�a<O�a<k�a<W�a<g�a<j�a<��a<��a<��a<Ѝa<ōa<�  �  �a<�a<)�a<Q�a<��a<��a<ߎa<��a<H�a<v�a<��a<�a<�a<d�a<��a<�a<-�a<��a<͑a<6�a<��a<̒a<6�a<��a<�a<I�a<��a<	�a<j�a<ɕa<2�a<��a<�a<��a<��a<K�a<Ԙa<C�a<��a<*�a<��a<�a<��a<��a<p�a<�a<[�a<۝a<U�a<��a<G�a<��a<�a<��a<��a<e�a<աa<D�a<��a<#�a<��a<�a<b�a<̤a<*�a<��a<�a<>�a<��a<�a<<�a<��a<�a<B�a<��a<ڨa<�a<j�a<��a<�a<2�a<`�a<��a<ժa<�a<A�a<{�a<��a<۫a<�a<*�a<b�a<��a<��a<Ƭa<Ѭa<��a<�a<.�a<=�a<f�a<q�a<��a<��a<��a<��a<ŭa<ɭa<έa<ѭa<ۭa<׭a<Эa<˭a<ݭa<ѭa<έa<Эa<��a<��a<��a<��a<��a<`�a<N�a<E�a<0�a<�a<��a<�a<ɬa<��a<w�a<r�a<E�a<�a<��a<��a<��a<j�a<D�a<�a<�a<��a<��a<\�a<�a<�a<��a<d�a<+�a<�a<��a<_�a<�a<ͧa<��a<C�a<��a<��a<M�a<�a<��a<j�a<�a<��a<U�a<�a<��a<M�a<�a<��a<4�a<աa<b�a<�a<��a<,�a<��a<Q�a<�a<{�a<�a<��a<;�a<ɜa<r�a<��a<��a<�a<��a<7�a<˙a<R�a<�a<z�a<�a<��a<L�a<�a<}�a<�a<��a<P�a<�a<��a<%�a<Óa<p�a<�a<a<v�a<�a<֑a<��a<6�a<��a<��a<[�a<,�a<ُa<��a<l�a<7�a<��a<ݎa<��a<��a<g�a<'�a<�a<��a<Սa<��a<��a<��a<~�a<j�a<\�a<j�a<`�a<d�a<q�a<T�a<��a<��a<��a<��a<��a<a<�  �  ܍a<�a<%�a<R�a<��a<��a<ێa<�a<3�a<V�a<��a<ُa<�a<}�a<��a<
�a</�a<��a<Αa<�a<u�a<̒a<1�a<u�a<��a<;�a<��a<�a<d�a<��a</�a<��a<�a<u�a<��a<W�a<ژa</�a<��a<�a<��a<$�a<{�a<�a<_�a<�a<T�a<ŝa<N�a<��a<4�a<��a<�a<|�a<�a<d�a<ʡa<[�a<��a<)�a<q�a<��a<?�a<¤a<�a<v�a<�a</�a<��a<�a<U�a<��a<ڧa<K�a<z�a<ۨa<�a<i�a<��a<�a<4�a<U�a<Īa<۪a<�a<M�a<n�a<��a<ūa<�a<(�a<E�a<q�a<��a<��a<Ҭa<�a<��a<?�a<H�a<T�a<v�a<j�a<��a<��a<��a<��a<έa<խa<ǭa<�a<ɭa<��a<ڭa<ɭa<�a<��a<ϭa<��a<��a<��a<��a<y�a<j�a<��a<7�a<C�a<�a<��a<�a<��a<��a<q�a<]�a<%�a<�a<�a<��a<��a<I�a<]�a<�a<�a<��a<r�a<A�a<�a<ߩa<��a<t�a<�a<�a<��a<Y�a<C�a<˧a<��a<J�a<�a<��a<X�a<�a<��a<v�a<�a<ˤa<v�a<��a<��a<<�a<��a<��a<�a<Ρa<G�a< �a<v�a<2�a<��a<d�a<�a<p�a<&�a<��a<B�a<��a<_�a<՛a<��a<�a<��a<D�a<��a<l�a<�a<��a<2�a<��a<U�a<ϖa<~�a<�a<��a<D�a<�a<��a<�a<�a<u�a<#�a<Βa<i�a<1�a<��a<��a<4�a<�a<��a<S�a<'�a<ڏa<��a<O�a<H�a<�a<ʎa<��a<b�a<V�a<�a<�a<ݍa<ۍa<��a<��a<��a<p�a<��a<l�a<V�a<p�a<N�a<p�a<`�a<|�a<m�a<��a<��a<��a<��a<�  �  �a<��a<6�a<N�a<w�a<��a<Ԏa<�a</�a<z�a<��a<؏a<�a<h�a<��a<�a<0�a<��a<�a<9�a<r�a<�a<&�a<��a<ݓa<A�a<��a<��a<d�a<ɕa<D�a<��a<�a<u�a<�a<f�a<ɘa<9�a<��a<%�a<��a< �a<y�a<�a<{�a<ޜa<d�a<ʝa<U�a<��a<4�a<��a<�a<}�a<�a<i�a<סa<>�a<��a<&�a<��a<��a<W�a<Ѥa<�a<��a<٥a<F�a<��a<�a<7�a<��a<�a<8�a<��a<Ψa<'�a<j�a<��a<�a<'�a<j�a<��a<Ϫa<��a<C�a<x�a<��a<�a<��a<@�a<J�a<��a<��a<��a<Ҭa<�a<�a<2�a<>�a<Q�a<x�a<��a<��a<��a<��a<��a<ȭa<˭a<ޭa<ʭa<ԭa<ϭa<ۭa<֭a<ҭa<ȭa<��a<��a<��a<��a<��a<��a<s�a<R�a<@�a< �a< �a<��a<ެa<¬a<��a<��a<Y�a<I�a< �a<�a<��a<��a<s�a<@�a<
�a<�a<��a<��a<?�a<&�a<ԩa<��a<\�a<#�a<�a<��a<Z�a<�a<ߧa<��a<L�a<�a<��a<g�a<	�a<��a<b�a<�a<��a<S�a<��a<��a<X�a<�a<��a<#�a<աa<d�a<��a<��a<2�a<��a<J�a<�a<}�a<	�a<��a<?�a<לa<g�a<�a<��a<�a<��a<0�a<әa<T�a<�a<u�a<�a<��a<B�a<ؖa<p�a<�a<��a<@�a<�a<��a</�a<œa<j�a<
�a<Ēa<s�a<�a<ۑa<{�a<L�a<�a<��a<r�a<'�a<ڏa<��a<n�a<<�a<��a<Ȏa<��a<��a<Q�a<;�a<�a<�a<ԍa<��a<��a<��a<{�a<h�a<l�a<d�a<b�a<]�a<_�a<p�a<m�a<y�a<��a<��a<��a<ōa<�  �  ��a<Q�a<��a<��a<؍a<%�a<,�a<��a<��a<Ԏa<�a<`�a<��a<��a<2�a<G�a<ǐa<�a<+�a<��a<ۑa<V�a<��a<�a<:�a<˓a<�a<s�a<�a<@�a<ѕa<�a<��a<�a<l�a<��a<7�a<��a<�a<��a<'�a<��a<,�a<F�a<	�a<K�a<�a<X�a<ǝa<G�a<��a<*�a<v�a<.�a<~�a<��a<m�a<ȡa<]�a<��a<�a<n�a<�a<Q�a<��a<&�a<P�a<�a<��a<��a<��a<9�a<��a<��a< �a<[�a<��a<��a<1�a<��a<��a<�a<.�a<��a<��a<��a<#�a<�a<��a<��a<ͫa<ثa<�a<�a<B�a<��a<w�a<��a<��a<ެa<�a<ܬa<�a<�a<L�a<2�a<Z�a<X�a<X�a<u�a<8�a<��a<n�a<|�a<i�a<P�a<X�a<G�a<_�a<:�a<.�a<�a<�a<�a<�a<�a<��a<��a<��a<c�a<h�a<"�a<'�a<׫a<ƫa<��a<��a<h�a<�a<�a<��a<ªa<o�a<'�a<�a<ǩa<��a<X�a<M�a<רa<ʨa<b�a<+�a<"�a<��a<��a<
�a<Ԧa<�a<B�a<��a<��a<L�a<٤a<��a<X�a<�a<��a<�a<�a<^�a<&�a<��a<N�a<�a<m�a<�a<��a<g�a<ٞa<u�a<�a<��a<G�a<��a<N�a<͛a<p�a<�a<��a<8�a<��a<b�a<��a<��a<�a<��a<6�a<��a<Z�a<�a<��a<)�a<��a<b�a<�a<��a<<�a<�a<��a<�a<��a<s�a<`�a<�a<��a<Q�a<�a<��a<��a<r�a<�a<�a<��a<w�a<Z�a<�a<�a<��a<��a<h�a<f�a<>�a<�a<�a<ˌa<!�a<�a<�a<ьa<��a<Ȍa<��a<�a<ٌa<�a<�a<�a<:�a<4�a<�  �  J�a<u�a<��a<��a<�a<�a<0�a<|�a<��a<�a<�a<K�a<��a<Ǐa<�a<T�a<��a<�a<O�a<��a<�a<R�a<��a<��a<J�a<Ǔa<%�a<�a<̔a<1�a<��a<�a<��a<�a<n�a<חa<R�a<��a<4�a<��a<�a<i�a<�a<�a<�a<^�a<�a<M�a<͝a<M�a<��a<<�a<��a<�a<x�a<�a<\�a<ɡa<5�a<��a<(�a<��a<��a<U�a<��a<�a<d�a<�a<1�a<��a<��a<*�a<��a<ԧa<$�a<v�a<��a<��a<J�a<��a<��a<�a<"�a<T�a<��a<�a<�a<+�a<m�a<��a<ͫa<�a<�a<;�a<G�a<d�a<��a<��a<��a<̬a<�a<�a<$�a<-�a<D�a<9�a<H�a<Z�a<^�a<w�a<i�a<a�a<I�a<p�a<h�a<k�a<^�a<W�a<N�a<?�a<5�a<+�a<�a<�a<ˬa<ʬa<��a<��a<��a<n�a<R�a<%�a<�a<��a<ثa<��a<z�a<J�a<!�a<��a<Ȫa<��a<k�a<J�a<�a<۩a<��a<\�a<2�a<�a<ƨa<��a<8�a<ݧa<��a<q�a<�a<�a<��a<D�a<�a<��a<O�a<��a<��a<J�a<̣a<��a<=�a<�a<q�a<�a<��a<T�a<��a<��a</�a<��a<?�a<Ӟa<k�a<��a<��a<�a<��a<_�a<�a<��a<
�a<��a<+�a<��a<Z�a<�a<n�a<ߗa<��a<-�a<Ŗa<^�a<��a<��a<+�a<ϔa<k�a<��a<��a<0�a<Βa<��a<F�a<��a<��a<F�a<�a<��a<d�a<(�a<��a<��a<H�a<�a<ӎa<��a<e�a<?�a<�a<��a<ƍa<��a<o�a<T�a<A�a<$�a<!�a<��a<�a<��a<یa<Ќa<Ԍa<͌a<ьa<،a<ތa<�a<�a<�a<(�a<�a<�  �  K�a<��a<��a<��a<�a<�a<J�a<\�a<��a<a<�a<L�a<��a<�a<��a<��a<��a<��a<E�a<��a<�a<6�a<��a<�a<g�a<��a<�a<��a<ߔa<m�a<��a<�a<��a<�a<d�a<ȗa<V�a<��a<B�a<��a<2�a<��a<�a<��a<؛a<n�a<��a<W�a<ʝa<&�a<��a<�a<��a<�a<��a<�a<Z�a<�a<0�a<��a<�a<w�a<Уa<G�a<��a<�a<}�a<��a<;�a<��a<�a<O�a<s�a<�a<	�a<t�a<��a<�a<<�a<p�a<ĩa<�a<[�a<o�a<��a<۪a<��a<L�a<g�a<��a<��a<ԫa<��a<$�a<S�a<]�a<��a<��a<Ҭa<ݬa<�a<�a<��a<%�a<�a<N�a<N�a<_�a<Y�a<Q�a<��a<`�a<��a<x�a<Y�a<q�a<I�a<X�a<<�a<A�a<%�a<+�a<�a<	�a<�a<ˬa<Ԭa<��a<��a<|�a<Q�a<@�a<��a<�a<��a<��a<{�a<Q�a<D�a<�a<��a<��a<t�a<@�a<��a<̩a<��a<x�a<)�a<�a<��a<p�a<F�a<�a<ҧa<`�a<�a<Цa<��a<:�a<ߥa<��a<4�a<
�a<��a<c�a<��a<��a<N�a<��a<��a<�a<��a<Q�a<Ҡa<~�a<�a<��a<:�a<��a<q�a<��a<��a<�a<Ȝa<:�a<֛a<Y�a<��a<��a<'�a<��a<3�a<�a<o�a<�a<��a<�a<іa<C�a<��a<{�a<�a<��a<Q�a<�a<��a<i�a<�a<��a<;�a<בa<��a<@�a<�a<��a<M�a<
�a<ɏa<��a<A�a<9�a<Ŏa<��a<v�a<9�a<�a<Ѝa<��a<��a<��a<Z�a<E�a<�a<��a<�a<�a<��a<�a<��a<ڌa<��a<ӌa<ƌa<��a<݌a<�a<�a<+�a<U�a<�  �  ]�a<o�a<��a<��a<ߍa<�a<E�a<k�a<��a<ڎa<�a<V�a<|�a<Џa<�a<Y�a<��a< �a<<�a<��a<��a<@�a<��a<�a<[�a<��a<�a<}�a<�a<?�a<��a<$�a<��a<��a<j�a<ڗa<S�a<��a<5�a<��a<�a<��a<�a<s�a<��a<q�a<֜a<T�a<̝a<B�a<Ȟa<�a<��a<�a<z�a<�a<d�a<ʡa<6�a<��a<�a<��a<�a<L�a<��a<�a<y�a<إa<'�a<��a<ڦa<!�a<v�a<֧a<�a<p�a<��a<��a<A�a<��a<ǩa<�a<)�a<s�a<��a<תa<�a<@�a<^�a<��a<��a<�a<�a<$�a<Z�a<_�a<��a<��a<��a<Ǭa<�a<�a<�a<@�a<3�a<H�a<J�a<Q�a<g�a<k�a<b�a<n�a<j�a<X�a<b�a<g�a<\�a<Z�a<K�a<D�a<2�a<#�a<�a<�a<�a<ݬa<��a<��a<��a<k�a<G�a<:�a<�a<�a<ͫa<��a<��a<B�a<+�a<��a<ͪa<��a<}�a<8�a<�a<�a<��a<s�a<"�a<��a<��a<s�a<6�a<��a<��a<W�a<&�a<٦a<��a<@�a<�a<��a<K�a<��a<��a<8�a<�a<��a<1�a<�a<��a<�a<��a<S�a<�a<��a<�a<��a<A�a<՞a<q�a<�a<��a< �a<Ĝa<E�a<�a<w�a<�a<��a<�a<��a<Q�a<טa<q�a<�a<��a< �a<ǖa<X�a<��a<��a<(�a<Ɣa<e�a<�a<��a<7�a<�a<��a<7�a<�a<��a<6�a<��a<��a<k�a<'�a<ɏa<��a<C�a<�a<؎a<��a<`�a<A�a<�a<�a<ٍa<��a<~�a<U�a<7�a<-�a<�a<��a<�a<݌a<Ìa<ʌa<Ќa<ˌa<Ԍa<Ռa<�a<�a<��a<
�a<�a<4�a<�  �  g�a<b�a<��a<��a<�a<�a<:�a<u�a<��a<؎a<�a<V�a<��a<ˏa<#�a<P�a<��a<��a<;�a<��a<�a<O�a<��a<��a<N�a<��a<�a<r�a<�a<<�a<Еa<�a<��a<��a<Y�a<ߗa<=�a<ǘa<�a<��a<�a<��a<�a<o�a<��a<]�a<�a<Q�a<ǝa<B�a<��a<&�a<��a<�a<y�a<��a<o�a<ơa<P�a<��a<�a<q�a<�a<K�a<��a<�a<f�a<ޥa<$�a<��a<֦a<-�a<��a<��a<%�a<_�a<��a<�a<9�a<��a<��a<�a<,�a<w�a<��a<ݪa<�a<1�a<p�a<��a<ƫa<ܫa< �a<*�a<R�a<x�a<{�a<��a<��a<լa<��a<��a<�a<�a<;�a<=�a<O�a<\�a<X�a<q�a<X�a<z�a<Z�a<|�a<x�a<I�a<e�a<G�a<Q�a</�a<7�a<�a<�a<�a<٬a<�a<��a<��a<��a<p�a<T�a</�a<�a<�a<ʫa<��a<��a<T�a<%�a<�a<Īa<��a<w�a<7�a<�a<ͩa<��a<f�a<4�a<�a<��a<|�a<+�a<��a<��a<��a<�a<Ѧa<��a</�a<��a<��a<V�a<ޤa<��a<P�a<�a<��a<-�a<�a<p�a<%�a<��a<N�a<�a<t�a<�a<��a<W�a<Ԟa<v�a<�a<��a<:�a<��a<N�a<Лa<q�a< �a<��a<1�a<��a<W�a<Ԙa<u�a<��a<��a<H�a<��a<_�a<�a<��a<�a<��a<b�a<��a<��a<:�a<�a<��a<=�a<�a<��a<I�a<�a<��a<U�a<�a<Ϗa<��a<\�a<�a<�a<��a<m�a<L�a<�a<�a<��a<��a<s�a<[�a<C�a<�a<�a<�a<��a<Όa<�a<��a<��a<Ԍa<��a<یa<Όa<�a<�a<�a<9�a<(�a<�  �  W�a<z�a<��a<��a<�a<�a<A�a<v�a<��a<ڎa<�a<H�a<��a<ԏa<
�a<j�a<��a<�a<O�a<��a<�a<O�a<��a<��a<^�a<��a<�a<x�a<�a<M�a<��a<�a<��a<�a<b�a<�a<8�a<Ƙa<,�a<��a<�a<��a< �a<��a<�a<f�a<�a<P�a<ҝa<H�a<��a<0�a<��a<
�a<��a<�a<[�a<סa<<�a<��a<#�a<}�a<�a<V�a<��a<�a<u�a<ɥa<,�a<{�a<ܦa<(�a<s�a<Χa<)�a<]�a<��a<��a<5�a<��a<��a<�a<7�a<s�a<��a<ڪa<�a<E�a<h�a<��a<ɫa<�a<�a<9�a<F�a<m�a<��a<��a<��a<�a<�a<�a<�a<#�a<:�a<J�a<F�a<\�a<V�a<b�a<q�a<m�a<i�a<f�a<Y�a<b�a<c�a<H�a<]�a<6�a<4�a<'�a<�a<��a<�a<׬a<ìa<��a<��a<w�a<J�a<7�a<�a<�a<ͫa<��a<v�a<\�a<.�a<�a<ުa<��a<i�a<J�a<�a<ީa<��a<c�a<+�a<��a<��a<{�a<1�a<��a<��a<_�a<�a<ڦa<��a<8�a<��a<��a<V�a<��a<��a<A�a<�a<��a<@�a<Ӣa<y�a<�a<��a<Y�a<��a<��a<#�a<��a<B�a<�a<h�a<��a<��a<&�a<��a<Z�a<ݛa<y�a<�a<��a<)�a<��a<B�a<ܘa<e�a<�a<��a<�a<��a<c�a<�a<��a<%�a<��a<e�a<��a<��a<E�a<�a<��a<:�a<ܑa<��a<@�a<�a<��a<f�a<�a<ޏa<��a<Q�a< �a<юa<��a<y�a<:�a<�a<�a<��a<��a<��a<R�a<C�a<�a<�a<�a<�a<݌a<ьa<��a<ˌa<Ҍa<Ìa<�a<Ռa<�a<��a<��a<�a<9�a<�  �  B�a<}�a<��a<̍a<�a<�a<F�a<[�a<��a<͎a<#�a<^�a<��a<Ώa<�a<^�a<��a<�a<M�a<��a<��a<2�a<��a<�a<l�a<��a<�a<��a<Ӕa<O�a<��a<4�a<��a<�a<g�a<ӗa<B�a<��a<G�a<��a<�a<��a<��a<��a<�a<��a<לa<Y�a<˝a<=�a<��a< �a<��a<�a<�a<��a<c�a<̡a<9�a<Ǣa<�a<��a<�a<I�a<��a<�a<��a<åa<1�a<|�a<�a</�a<}�a<�a<�a<a�a<��a<��a<7�a<z�a<ةa<�a<:�a<g�a<��a<ުa<	�a<T�a<`�a<��a<��a<�a<�a<1�a<h�a<e�a<��a<��a<¬a<Ҭa<��a<�a<	�a<.�a<$�a<J�a<M�a<_�a<q�a<]�a<p�a<W�a<r�a<^�a<n�a<t�a<M�a<Q�a<@�a<9�a<"�a<1�a<�a<�a<�a<¬a<Ǭa<��a<��a<}�a<K�a<;�a<��a<��a<��a<��a<��a<K�a<(�a<��a<Ҫa<��a<��a<H�a<�a<�a<��a<r�a<(�a<�a<��a<y�a<<�a<�a<��a<Y�a<6�a<٦a<��a<>�a<�a<��a<@�a<�a<��a<C�a<��a<��a<@�a<΢a<��a<�a<��a<R�a<�a<��a<�a<Пa<D�a<ڞa<r�a<�a<��a<#�a<לa<J�a<�a<w�a<��a<��a<�a<Йa<<�a<�a<f�a<	�a<��a<'�a<ٖa<N�a<�a<��a<$�a<��a<[�a<�a<��a<H�a<�a<��a<>�a<�a<��a<8�a<��a<��a<j�a<�a<֏a<��a<H�a<�a<؎a<��a<j�a<I�a<(�a<ۍa<Ǎa<��a<��a<Y�a<E�a<6�a<�a<�a<،a<�a<Ɍa<Ռa<݌a<��a<̌a<ˌa<،a<یa<�a<�a<�a<B�a<�  �  _�a<v�a<��a<Ía<ߍa<�a<@�a<q�a<��a<Ԏa<�a<W�a<��a<̏a<+�a<R�a<��a<��a<:�a<��a<�a<G�a<��a<��a<P�a<��a<�a<��a<�a<D�a<��a<�a<��a<��a<a�a<˗a<O�a<��a<$�a<��a<�a<��a<�a<v�a<�a<p�a<Ԝa<S�a<a<F�a<��a< �a<��a<�a<~�a<��a<o�a<ˡa<N�a<��a<�a<{�a<�a<E�a<��a<�a<w�a<ѥa<*�a<��a<�a<(�a<��a<ǧa<�a<l�a<��a<�a<@�a<u�a<��a<��a<2�a<u�a<��a<Ӫa<�a<8�a<b�a<��a<��a<�a<�a<"�a<N�a<{�a<{�a<��a<��a<֬a<��a<��a<�a<+�a<9�a<A�a<T�a<S�a<e�a<_�a<c�a<u�a<o�a<i�a<m�a<V�a<Y�a<[�a<;�a<@�a<2�a<�a<�a<��a<�a<߬a<��a<��a<��a<k�a<V�a<6�a<�a<�a<ƫa<��a<��a<X�a<&�a<�a<ƪa<��a<s�a<5�a<
�a<٩a<��a<t�a<*�a<�a<��a<n�a<>�a<��a<��a<h�a< �a<Φa<��a<8�a<�a<��a<H�a<�a<��a<A�a<��a<��a<4�a<آa<��a<�a<��a<I�a<�a<��a<�a<��a<S�a<ٞa<w�a<�a<��a<8�a<��a<C�a<ۛa<u�a<��a<��a<�a<��a<J�a<ژa<v�a<�a<��a<5�a<��a<S�a<��a<�a<�a<Ŕa<W�a<��a<��a<@�a<�a<��a<3�a<�a<��a<;�a<��a<��a<a�a<�a<Ǐa<��a<_�a<�a<�a<��a<o�a<F�a<	�a<�a<ča<��a<w�a<_�a<9�a<+�a<	�a<��a<��a<�a<Ԍa<Ԍa<��a<Ȍa<Ռa<Ōa<ߌa<�a<�a<�a<!�a<<�a<�  �  ]�a<q�a<��a<��a<��a<�a<,�a<��a<��a<�a<�a<C�a<��a<Ïa< �a<T�a<��a<ܐa<^�a<��a<ߑa<R�a<��a<�a<Q�a<��a<�a<w�a<�a<<�a<��a<�a<��a<�a<c�a<�a<6�a<Ƙa</�a<��a<�a<��a<	�a<w�a<��a<\�a<�a<W�a<ʝa<G�a<��a<G�a<��a<�a<��a<�a<f�a<͡a<H�a<��a<6�a<~�a<�a<R�a<��a<!�a<f�a<ڥa<(�a<��a<צa<�a<�a<ͧa<+�a<X�a<��a<��a<2�a<��a<��a<��a<&�a<r�a<��a<תa<�a<3�a<w�a<��a<ʫa<ݫa<�a<K�a<6�a<}�a<��a<��a<��a<ެa<�a<�a<3�a<�a<C�a<6�a<V�a<W�a<W�a<g�a<e�a<t�a<^�a<c�a<X�a<e�a<^�a<D�a<U�a<3�a</�a<&�a<�a<��a<ެa<ݬa<��a<��a<��a<l�a<]�a<!�a<$�a<߫a<�a<��a<r�a<]�a<�a<
�a<Ȫa<��a<Z�a<Y�a<�a<ʩa<��a<Y�a<<�a<�a<��a<w�a<0�a<��a<��a<e�a<�a<�a<��a<9�a<��a<��a<V�a<��a<��a<<�a<�a<��a<5�a<�a<o�a<"�a<��a<Q�a<�a<}�a<9�a<��a<N�a<۞a<o�a<�a<��a<2�a<��a<m�a<ݛa<r�a<�a<��a<3�a<��a<S�a<ؘa<l�a<��a<��a<)�a<��a<e�a<ߕa<��a<$�a<��a<k�a<��a<��a<4�a<�a<��a<7�a<�a<��a<O�a<�a<��a<V�a<#�a<�a<x�a<`�a<�a<�a<��a<w�a<:�a<�a<�a<��a<��a<l�a<a�a<=�a<�a<�a<��a<��a<ьa<Όa<��a<Όa<͌a<��a<��a<Ҍa<�a<��a<��a<�a<,�a<�  �  R�a<|�a<��a<��a<�a<�a<:�a<v�a<��a<Ύa<�a<Q�a<��a<؏a<�a<g�a<��a<��a<A�a<��a<�a<H�a<��a< �a<`�a<��a<�a<��a<��a<b�a<��a<�a<��a<�a<e�a<ӗa<=�a<��a<8�a<��a<'�a<��a<�a<�a<�a<m�a<�a<S�a<͝a<D�a<��a<�a<��a<�a<��a<��a<g�a<ۡa<C�a<��a<�a<u�a<�a<Q�a<��a<�a<y�a<ĥa<,�a<��a<�a<=�a<v�a<קa<�a<]�a<��a<��a<0�a<u�a<©a<�a<J�a<p�a<��a<٪a<�a<F�a<p�a<��a<«a<�a<��a<(�a<W�a<q�a<��a<��a<Ƭa<�a<�a<
�a<�a<�a<<�a<B�a<L�a<\�a<b�a<U�a<p�a<f�a<y�a<p�a<[�a<i�a<H�a<M�a<B�a<:�a<�a<(�a<
�a<�a<��a<Ҭa<Ƭa<��a<��a<t�a<V�a</�a<�a<�a<��a<��a<��a<[�a<3�a<�a<۪a<��a<|�a<=�a<��a<کa<��a<b�a<6�a<��a<��a<u�a<8�a<�a<Ƨa<b�a<!�a<Ѧa<y�a<;�a<�a<��a<;�a< �a<��a<X�a<��a<��a<=�a<͢a<��a<"�a<��a<T�a<�a<x�a<�a<��a<O�a<�a<w�a<�a<��a<-�a<Ɯa<E�a<՛a<s�a<�a<��a</�a<��a<=�a<ݘa<k�a<�a<��a< �a<Ȗa<J�a<�a<��a<#�a<��a<V�a<�a<��a<X�a<�a<��a<9�a<ݑa<��a<H�a<�a<��a<`�a<�a<͏a<��a<T�a<!�a<�a<��a<z�a<D�a<�a<؍a<��a<��a<x�a<X�a<C�a<'�a<��a<�a<�a<�a<یa<Ìa<ӌa<��a<Ȍa<̌a<ٌa<Ԍa<��a<�a<$�a<L�a<�  �  E�a<��a<��a<ˍa<؍a<�a<R�a<e�a<��a<ߎa<�a<W�a<��a<Տa<
�a<f�a<��a<	�a<:�a<��a<�a<<�a<��a<�a<T�a<��a<�a<��a<ʔa<G�a<��a<)�a<~�a< �a<r�a<a<h�a<��a<2�a<��a<	�a<y�a<��a<��a<�a<w�a<Μa<Z�a<ԝa<C�a<۞a<!�a<��a<�a<��a<�a<Y�a<ߡa<0�a<��a<�a<��a<�a<R�a<��a<��a<�a<ҥa<3�a<z�a<¦a< �a<l�a<٧a<�a<��a<��a<��a<M�a<o�a<˩a<�a<0�a<V�a<��a<۪a<�a<?�a<O�a<��a<��a<��a<#�a<#�a<d�a<Y�a<��a<��a<��a<լa<�a<�a<�a<I�a<1�a<U�a<F�a<K�a<p�a<^�a<v�a<\�a<a�a<U�a<g�a<`�a<N�a<r�a<*�a<W�a<(�a<�a<�a<�a<�a<Ŭa<̬a<��a<��a<c�a<G�a<G�a<	�a<�a<ѫa<��a<��a<N�a</�a<�a<ڪa<��a<��a<5�a< �a<�a<��a<��a<�a<�a<��a<x�a<>�a<ڧa<��a<O�a<+�a<ʦa<��a<H�a<٥a<��a<7�a<��a<��a<:�a<ۣa<��a<D�a<ۢa<��a<	�a<��a<Z�a<�a<��a<�a<��a<9�a<�a<l�a<��a<��a<�a<Ϝa<C�a<�a<w�a<�a<��a<�a<ęa<K�a<�a<d�a<�a<��a<�a<ɖa<E�a<
�a<z�a<'�a<Ҕa<P�a<�a<��a<>�a<Вa<��a<:�a<�a<��a<'�a<�a<��a<n�a<0�a<ȏa<��a<<�a<#�a<ώa<��a<m�a<@�a<�a<�a<�a<��a<��a<R�a<1�a<5�a<�a<	�a<݌a<Ԍa<��a<όa<Ɍa<��a<�a<��a<��a<��a<��a<�a<	�a<5�a<�  �  b�a<f�a<��a<��a<�a<�a<>�a<a�a<��a<�a<�a<\�a<��a<֏a<�a<d�a<��a< �a<K�a<��a<ˑa<=�a<��a<�a<U�a<��a<�a<v�a<�a<P�a<��a<�a<��a<�a<^�a<̗a<?�a<��a<%�a<��a<(�a<��a<�a<m�a<��a<V�a<�a<`�a<Νa<$�a<��a<2�a<��a<�a<��a<��a<g�a<�a<J�a<��a<�a<z�a<ɣa<P�a<��a<#�a<b�a<֥a<�a<��a<�a<<�a<��a<Ƨa<�a<]�a<��a<�a<0�a<t�a<��a<�a<=�a<|�a<��a<Ӫa<�a<6�a<|�a<��a<��a<ëa<�a<4�a<W�a<r�a<��a<��a<ɬa<�a<��a< �a<!�a<�a<"�a<D�a<[�a<f�a<T�a<e�a<Z�a<x�a<m�a<u�a<l�a<X�a<O�a<G�a<<�a<1�a<$�a<�a<�a<
�a<�a<�a<��a<��a<��a<w�a<a�a<3�a<�a<ҫa<ԫa<��a<��a<\�a<0�a<�a<تa<��a<}�a<G�a<�a<��a<��a<l�a<C�a<�a<��a<o�a<.�a<�a<��a<v�a<�a<Ѧa<}�a<5�a<�a<��a<?�a<�a<��a<Y�a<��a<��a<+�a<ߢa<h�a<)�a<��a<U�a<Ϡa<v�a<%�a<��a<U�a<�a<x�a<	�a<��a<4�a<��a<S�a<ٛa<R�a<�a<��a<5�a<��a<O�a<Ϙa<w�a<�a<��a<9�a<��a<K�a<�a<��a<�a<��a<V�a<��a<��a<K�a<��a<��a<3�a<�a<��a<U�a<��a<��a<;�a<�a<ُa<��a<V�a<�a<ߎa<��a<z�a<P�a<�a<�a<��a<��a<z�a<g�a<L�a<�a<�a<�a<��a<��a<�a<ӌa<��a<��a<a<ƌa<Ќa<܌a<�a<�a<,�a<=�a<�  �  i�a<c�a<��a<��a<�a<�a<!�a<��a<��a<��a<
�a<F�a<��a<ӏa<,�a<P�a<��a<�a<L�a<��a<��a<y�a<k�a<�a<K�a<��a<!�a<o�a<��a<0�a<��a<�a<��a<��a<_�a<�a<4�a<ژa<�a<��a<�a<��a<�a<j�a<�a<F�a<��a<4�a<םa<e�a<��a<B�a<��a<�a<x�a<��a<l�a<ǡa<E�a<��a<)�a<��a<	�a<h�a<��a<-�a<P�a<�a<"�a<��a<Ԧa<�a<|�a<��a<:�a<Y�a<��a<��a<7�a<��a<��a<��a<�a<x�a<��a<�a<�a<&�a<��a<a�a<�a<��a<�a<6�a<6�a<o�a<|�a<��a<Ǭa<Ьa<�a<�a<6�a<�a<g�a<3�a<@�a<i�a<C�a<��a<U�a<|�a<W�a<f�a<G�a<b�a<u�a<<�a<f�a<)�a<D�a<+�a<�a<��a<Ӭa<�a<��a<��a<z�a<x�a<Q�a<�a<I�a<�a<�a<��a<u�a<R�a<.�a<�a<Īa<��a<a�a<G�a<�a<�a<שa<7�a<D�a<�a<��a<�a<(�a<�a<��a<a�a<��a<�a<��a<6�a< �a<��a<i�a<�a<��a<>�a<�a<��a<(�a<��a<Y�a<2�a<��a<^�a<�a<��a<4�a<��a<O�a<Ӟa<x�a<�a<��a</�a<��a<`�a<�a<��a<�a<k�a<?�a<��a<^�a<Ҙa<t�a<��a<��a<&�a<��a<t�a<�a<��a<#�a<��a<{�a<ԓa<��a<*�a<�a<��a<@�a<�a<|�a<Z�a<��a<Րa<q�a<'�a<ۏa<y�a<S�a<�a<�a<��a<h�a<?�a<�a<�a<��a<̍a<i�a<L�a<O�a<	�a<*�a<�a<��a<ˌa<Ҍa<��a<ˌa<�a<��a<��a<Ȍa<��a<�a<�a<�a<"�a<�  �  b�a<f�a<��a<��a<�a<�a<>�a<a�a<��a<�a<�a<\�a<��a<֏a<�a<d�a<��a< �a<K�a<��a<ˑa<=�a<��a<�a<U�a<��a<�a<v�a<�a<P�a<��a<�a<��a<�a<^�a<̗a<?�a<��a<%�a<��a<(�a<��a<�a<m�a<��a<V�a<�a<`�a<Νa<$�a<��a<2�a<��a<�a<��a<��a<g�a<�a<J�a<��a<�a<z�a<ɣa<P�a<��a<#�a<b�a<֥a<�a<��a<�a<<�a<��a<Ƨa<�a<]�a<��a<�a<0�a<t�a<��a<�a<=�a<|�a<��a<Ӫa<�a<6�a<|�a<��a<��a<ëa<�a<4�a<W�a<r�a<��a<��a<ɬa<�a<��a< �a<!�a<�a<"�a<D�a<[�a<f�a<T�a<e�a<Z�a<x�a<m�a<u�a<l�a<X�a<O�a<G�a<<�a<1�a<$�a<�a<�a<
�a<�a<�a<��a<��a<��a<w�a<a�a<3�a<�a<ҫa<ԫa<��a<��a<\�a<0�a<�a<تa<��a<}�a<G�a<�a<��a<��a<l�a<C�a<�a<��a<o�a<.�a<�a<��a<v�a<�a<Ѧa<}�a<5�a<�a<��a<?�a<�a<��a<Y�a<��a<��a<+�a<ߢa<h�a<)�a<��a<U�a<Ϡa<v�a<%�a<��a<U�a<�a<x�a<	�a<��a<4�a<��a<S�a<ٛa<R�a<�a<��a<5�a<��a<O�a<Ϙa<w�a<�a<��a<9�a<��a<K�a<�a<��a<�a<��a<V�a<��a<��a<K�a<��a<��a<3�a<�a<��a<U�a<��a<��a<;�a<�a<ُa<��a<V�a<�a<ߎa<��a<z�a<P�a<�a<�a<��a<��a<z�a<g�a<L�a<�a<�a<�a<��a<��a<�a<ӌa<��a<��a<a<ƌa<Ќa<܌a<�a<�a<,�a<=�a<�  �  E�a<��a<��a<ˍa<؍a<�a<R�a<e�a<��a<ߎa<�a<W�a<��a<Տa<
�a<f�a<��a<	�a<:�a<��a<�a<<�a<��a<�a<T�a<��a<�a<��a<ʔa<G�a<��a<)�a<~�a< �a<r�a<a<h�a<��a<2�a<��a<	�a<y�a<��a<��a<�a<w�a<Μa<Z�a<ԝa<C�a<۞a<!�a<��a<�a<��a<�a<Y�a<ߡa<0�a<��a<�a<��a<�a<R�a<��a<��a<�a<ҥa<3�a<z�a<¦a< �a<l�a<٧a<�a<��a<��a<��a<M�a<o�a<˩a<�a<0�a<V�a<��a<۪a<�a<?�a<O�a<��a<��a<��a<#�a<#�a<d�a<Y�a<��a<��a<��a<լa<�a<�a<�a<I�a<1�a<U�a<F�a<K�a<p�a<^�a<v�a<\�a<a�a<U�a<g�a<`�a<N�a<r�a<*�a<W�a<(�a<�a<�a<�a<�a<Ŭa<̬a<��a<��a<c�a<G�a<G�a<	�a<�a<ѫa<��a<��a<N�a</�a<�a<ڪa<��a<��a<5�a< �a<�a<��a<��a<�a<�a<��a<x�a<>�a<ڧa<��a<O�a<+�a<ʦa<��a<H�a<٥a<��a<7�a<��a<��a<:�a<ۣa<��a<D�a<ۢa<��a<	�a<��a<Z�a<�a<��a<�a<��a<9�a<�a<l�a<��a<��a<�a<Ϝa<C�a<�a<w�a<�a<��a<�a<ęa<K�a<�a<d�a<�a<��a<�a<ɖa<E�a<
�a<z�a<'�a<Ҕa<P�a<�a<��a<>�a<Вa<��a<:�a<�a<��a<'�a<�a<��a<n�a<0�a<ȏa<��a<<�a<#�a<ώa<��a<m�a<@�a<�a<�a<�a<��a<��a<R�a<1�a<5�a<�a<	�a<݌a<Ԍa<��a<όa<Ɍa<��a<�a<��a<��a<��a<��a<�a<	�a<5�a<�  �  R�a<|�a<��a<��a<�a<�a<:�a<v�a<��a<Ύa<�a<Q�a<��a<؏a<�a<g�a<��a<��a<A�a<��a<�a<H�a<��a< �a<`�a<��a<�a<��a<��a<b�a<��a<�a<��a<�a<e�a<ӗa<=�a<��a<8�a<��a<'�a<��a<�a<�a<�a<m�a<�a<S�a<͝a<D�a<��a<�a<��a<�a<��a<��a<g�a<ۡa<C�a<��a<�a<u�a<�a<Q�a<��a<�a<y�a<ĥa<,�a<��a<�a<=�a<v�a<קa<�a<]�a<��a<��a<0�a<u�a<©a<�a<J�a<p�a<��a<٪a<�a<F�a<p�a<��a<«a<�a<��a<(�a<W�a<q�a<��a<��a<Ƭa<�a<�a<
�a<�a<�a<<�a<B�a<L�a<\�a<b�a<U�a<p�a<f�a<y�a<p�a<[�a<i�a<H�a<M�a<B�a<:�a<�a<(�a<
�a<�a<��a<Ҭa<Ƭa<��a<��a<t�a<V�a</�a<�a<�a<��a<��a<��a<[�a<3�a<�a<۪a<��a<|�a<=�a<��a<کa<��a<b�a<6�a<��a<��a<u�a<8�a<�a<Ƨa<b�a<!�a<Ѧa<y�a<;�a<�a<��a<;�a< �a<��a<X�a<��a<��a<=�a<͢a<��a<"�a<��a<T�a<�a<x�a<�a<��a<O�a<�a<w�a<�a<��a<-�a<Ɯa<E�a<՛a<s�a<�a<��a</�a<��a<=�a<ݘa<k�a<�a<��a< �a<Ȗa<J�a<�a<��a<#�a<��a<V�a<�a<��a<X�a<�a<��a<9�a<ݑa<��a<H�a<�a<��a<`�a<�a<͏a<��a<T�a<!�a<�a<��a<z�a<D�a<�a<؍a<��a<��a<x�a<X�a<C�a<'�a<��a<�a<�a<�a<یa<Ìa<ӌa<��a<Ȍa<̌a<ٌa<Ԍa<��a<�a<$�a<L�a<�  �  ]�a<q�a<��a<��a<��a<�a<,�a<��a<��a<�a<�a<C�a<��a<Ïa< �a<T�a<��a<ܐa<^�a<��a<ߑa<R�a<��a<�a<Q�a<��a<�a<w�a<�a<<�a<��a<�a<��a<�a<c�a<�a<6�a<Ƙa</�a<��a<�a<��a<	�a<w�a<��a<\�a<�a<W�a<ʝa<G�a<��a<G�a<��a<�a<��a<�a<f�a<͡a<H�a<��a<6�a<~�a<�a<R�a<��a<!�a<f�a<ڥa<(�a<��a<צa<�a<�a<ͧa<+�a<X�a<��a<��a<2�a<��a<��a<��a<&�a<r�a<��a<תa<�a<3�a<w�a<��a<ʫa<ݫa<�a<K�a<6�a<}�a<��a<��a<��a<ެa<�a<�a<3�a<�a<C�a<6�a<V�a<W�a<W�a<g�a<e�a<t�a<^�a<c�a<X�a<e�a<^�a<D�a<U�a<3�a</�a<&�a<�a<��a<ެa<ݬa<��a<��a<��a<l�a<]�a<!�a<$�a<߫a<�a<��a<r�a<]�a<�a<
�a<Ȫa<��a<Z�a<Y�a<�a<ʩa<��a<Y�a<<�a<�a<��a<w�a<0�a<��a<��a<e�a<�a<�a<��a<9�a<��a<��a<V�a<��a<��a<<�a<�a<��a<5�a<�a<o�a<"�a<��a<Q�a<�a<}�a<9�a<��a<N�a<۞a<o�a<�a<��a<2�a<��a<m�a<ݛa<r�a<�a<��a<3�a<��a<S�a<ؘa<l�a<��a<��a<)�a<��a<e�a<ߕa<��a<$�a<��a<k�a<��a<��a<4�a<�a<��a<7�a<�a<��a<O�a<�a<��a<V�a<#�a<�a<x�a<`�a<�a<�a<��a<w�a<:�a<�a<�a<��a<��a<l�a<a�a<=�a<�a<�a<��a<��a<ьa<Όa<��a<Όa<͌a<��a<��a<Ҍa<�a<��a<��a<�a<,�a<�  �  _�a<v�a<��a<Ía<ߍa<�a<@�a<q�a<��a<Ԏa<�a<W�a<��a<̏a<+�a<R�a<��a<��a<:�a<��a<�a<G�a<��a<��a<P�a<��a<�a<��a<�a<D�a<��a<�a<��a<��a<a�a<˗a<O�a<��a<$�a<��a<�a<��a<�a<v�a<�a<p�a<Ԝa<S�a<a<F�a<��a< �a<��a<�a<~�a<��a<o�a<ˡa<N�a<��a<�a<{�a<�a<E�a<��a<�a<w�a<ѥa<*�a<��a<�a<(�a<��a<ǧa<�a<l�a<��a<�a<@�a<u�a<��a<��a<2�a<u�a<��a<Ӫa<�a<8�a<b�a<��a<��a<�a<�a<"�a<N�a<{�a<{�a<��a<��a<֬a<��a<��a<�a<+�a<9�a<A�a<T�a<S�a<e�a<_�a<c�a<u�a<o�a<i�a<m�a<V�a<Y�a<[�a<;�a<@�a<2�a<�a<�a<��a<�a<߬a<��a<��a<��a<k�a<V�a<6�a<�a<�a<ƫa<��a<��a<X�a<&�a<�a<ƪa<��a<s�a<5�a<
�a<٩a<��a<t�a<*�a<�a<��a<n�a<>�a<��a<��a<h�a< �a<Φa<��a<8�a<�a<��a<H�a<�a<��a<A�a<��a<��a<4�a<آa<��a<�a<��a<I�a<�a<��a<�a<��a<S�a<ٞa<w�a<�a<��a<8�a<��a<C�a<ۛa<u�a<��a<��a<�a<��a<J�a<ژa<v�a<�a<��a<5�a<��a<S�a<��a<�a<�a<Ŕa<W�a<��a<��a<@�a<�a<��a<3�a<�a<��a<;�a<��a<��a<a�a<�a<Ǐa<��a<_�a<�a<�a<��a<o�a<F�a<	�a<�a<ča<��a<w�a<_�a<9�a<+�a<	�a<��a<��a<�a<Ԍa<Ԍa<��a<Ȍa<Ռa<Ōa<ߌa<�a<�a<�a<!�a<<�a<�  �  B�a<}�a<��a<̍a<�a<�a<F�a<[�a<��a<͎a<#�a<^�a<��a<Ώa<�a<^�a<��a<�a<M�a<��a<��a<2�a<��a<�a<l�a<��a<�a<��a<Ӕa<O�a<��a<4�a<��a<�a<g�a<ӗa<B�a<��a<G�a<��a<�a<��a<��a<��a<�a<��a<לa<Y�a<˝a<=�a<��a< �a<��a<�a<�a<��a<c�a<̡a<9�a<Ǣa<�a<��a<�a<I�a<��a<�a<��a<åa<1�a<|�a<�a</�a<}�a<�a<�a<a�a<��a<��a<7�a<z�a<ةa<�a<:�a<g�a<��a<ުa<	�a<T�a<`�a<��a<��a<�a<�a<1�a<h�a<e�a<��a<��a<¬a<Ҭa<��a<�a<	�a<.�a<$�a<J�a<M�a<_�a<q�a<]�a<p�a<W�a<r�a<^�a<n�a<t�a<M�a<Q�a<@�a<9�a<"�a<1�a<�a<�a<�a<¬a<Ǭa<��a<��a<}�a<K�a<;�a<��a<��a<��a<��a<��a<K�a<(�a<��a<Ҫa<��a<��a<H�a<�a<�a<��a<r�a<(�a<�a<��a<y�a<<�a<�a<��a<Y�a<6�a<٦a<��a<>�a<�a<��a<@�a<�a<��a<C�a<��a<��a<@�a<΢a<��a<�a<��a<R�a<�a<��a<�a<Пa<D�a<ڞa<r�a<�a<��a<#�a<לa<J�a<�a<w�a<��a<��a<�a<Йa<<�a<�a<f�a<	�a<��a<'�a<ٖa<N�a<�a<��a<$�a<��a<[�a<�a<��a<H�a<�a<��a<>�a<�a<��a<8�a<��a<��a<j�a<�a<֏a<��a<H�a<�a<؎a<��a<j�a<I�a<(�a<ۍa<Ǎa<��a<��a<Y�a<E�a<6�a<�a<�a<،a<�a<Ɍa<Ռa<݌a<��a<̌a<ˌa<،a<یa<�a<�a<�a<B�a<�  �  W�a<z�a<��a<��a<�a<�a<A�a<v�a<��a<ڎa<�a<H�a<��a<ԏa<
�a<j�a<��a<�a<O�a<��a<�a<O�a<��a<��a<^�a<��a<�a<x�a<�a<M�a<��a<�a<��a<�a<b�a<�a<8�a<Ƙa<,�a<��a<�a<��a< �a<��a<�a<f�a<�a<P�a<ҝa<H�a<��a<0�a<��a<
�a<��a<�a<[�a<סa<<�a<��a<#�a<}�a<�a<V�a<��a<�a<u�a<ɥa<,�a<{�a<ܦa<(�a<s�a<Χa<)�a<]�a<��a<��a<5�a<��a<��a<�a<7�a<s�a<��a<ڪa<�a<E�a<h�a<��a<ɫa<�a<�a<9�a<F�a<m�a<��a<��a<��a<�a<�a<�a<�a<#�a<:�a<J�a<F�a<\�a<V�a<b�a<q�a<m�a<i�a<f�a<Y�a<b�a<c�a<H�a<]�a<6�a<4�a<'�a<�a<��a<�a<׬a<ìa<��a<��a<w�a<J�a<7�a<�a<�a<ͫa<��a<v�a<\�a<.�a<�a<ުa<��a<i�a<J�a<�a<ީa<��a<c�a<+�a<��a<��a<{�a<1�a<��a<��a<_�a<�a<ڦa<��a<8�a<��a<��a<V�a<��a<��a<A�a<�a<��a<@�a<Ӣa<y�a<�a<��a<Y�a<��a<��a<#�a<��a<B�a<�a<h�a<��a<��a<&�a<��a<Z�a<ݛa<y�a<�a<��a<)�a<��a<B�a<ܘa<e�a<�a<��a<�a<��a<c�a<�a<��a<%�a<��a<e�a<��a<��a<E�a<�a<��a<:�a<ܑa<��a<@�a<�a<��a<f�a<�a<ޏa<��a<Q�a< �a<юa<��a<y�a<:�a<�a<�a<��a<��a<��a<R�a<C�a<�a<�a<�a<�a<݌a<ьa<��a<ˌa<Ҍa<Ìa<�a<Ռa<�a<��a<��a<�a<9�a<�  �  g�a<b�a<��a<��a<�a<�a<:�a<u�a<��a<؎a<�a<V�a<��a<ˏa<#�a<P�a<��a<��a<;�a<��a<�a<O�a<��a<��a<N�a<��a<�a<r�a<�a<<�a<Еa<�a<��a<��a<Y�a<ߗa<=�a<ǘa<�a<��a<�a<��a<�a<o�a<��a<]�a<�a<Q�a<ǝa<B�a<��a<&�a<��a<�a<y�a<��a<o�a<ơa<P�a<��a<�a<q�a<�a<K�a<��a<�a<f�a<ޥa<$�a<��a<֦a<-�a<��a<��a<%�a<_�a<��a<�a<9�a<��a<��a<�a<,�a<w�a<��a<ݪa<�a<1�a<p�a<��a<ƫa<ܫa< �a<*�a<R�a<x�a<{�a<��a<��a<լa<��a<��a<�a<�a<;�a<=�a<O�a<\�a<X�a<q�a<X�a<z�a<Z�a<|�a<x�a<I�a<e�a<G�a<Q�a</�a<7�a<�a<�a<�a<٬a<�a<��a<��a<��a<p�a<T�a</�a<�a<�a<ʫa<��a<��a<T�a<%�a<�a<Īa<��a<w�a<7�a<�a<ͩa<��a<f�a<4�a<�a<��a<|�a<+�a<��a<��a<��a<�a<Ѧa<��a</�a<��a<��a<V�a<ޤa<��a<P�a<�a<��a<-�a<�a<p�a<%�a<��a<N�a<�a<t�a<�a<��a<W�a<Ԟa<v�a<�a<��a<:�a<��a<N�a<Лa<q�a< �a<��a<1�a<��a<W�a<Ԙa<u�a<��a<��a<H�a<��a<_�a<�a<��a<�a<��a<b�a<��a<��a<:�a<�a<��a<=�a<�a<��a<I�a<�a<��a<U�a<�a<Ϗa<��a<\�a<�a<�a<��a<m�a<L�a<�a<�a<��a<��a<s�a<[�a<C�a<�a<�a<�a<��a<Όa<�a<��a<��a<Ԍa<��a<یa<Όa<�a<�a<�a<9�a<(�a<�  �  ]�a<o�a<��a<��a<ߍa<�a<E�a<k�a<��a<ڎa<�a<V�a<|�a<Џa<�a<Y�a<��a< �a<<�a<��a<��a<@�a<��a<�a<[�a<��a<�a<}�a<�a<?�a<��a<$�a<��a<��a<j�a<ڗa<S�a<��a<5�a<��a<�a<��a<�a<s�a<��a<q�a<֜a<T�a<̝a<B�a<Ȟa<�a<��a<�a<z�a<�a<d�a<ʡa<6�a<��a<�a<��a<�a<L�a<��a<�a<y�a<إa<'�a<��a<ڦa<!�a<v�a<֧a<�a<p�a<��a<��a<A�a<��a<ǩa<�a<)�a<s�a<��a<תa<�a<@�a<^�a<��a<��a<�a<�a<$�a<Z�a<_�a<��a<��a<��a<Ǭa<�a<�a<�a<@�a<3�a<H�a<J�a<Q�a<g�a<k�a<b�a<n�a<j�a<X�a<b�a<g�a<\�a<Z�a<K�a<D�a<2�a<#�a<�a<�a<�a<ݬa<��a<��a<��a<k�a<G�a<:�a<�a<�a<ͫa<��a<��a<B�a<+�a<��a<ͪa<��a<}�a<8�a<�a<�a<��a<s�a<"�a<��a<��a<s�a<6�a<��a<��a<W�a<&�a<٦a<��a<@�a<�a<��a<K�a<��a<��a<8�a<�a<��a<1�a<�a<��a<�a<��a<S�a<�a<��a<�a<��a<A�a<՞a<q�a<�a<��a< �a<Ĝa<E�a<�a<w�a<�a<��a<�a<��a<Q�a<טa<q�a<�a<��a< �a<ǖa<X�a<��a<��a<(�a<Ɣa<e�a<�a<��a<7�a<�a<��a<7�a<�a<��a<6�a<��a<��a<k�a<'�a<ɏa<��a<C�a<�a<؎a<��a<`�a<A�a<�a<�a<ٍa<��a<~�a<U�a<7�a<-�a<�a<��a<�a<݌a<Ìa<ʌa<Ќa<ˌa<Ԍa<Ռa<�a<�a<��a<
�a<�a<4�a<�  �  K�a<��a<��a<��a<�a<�a<J�a<\�a<��a<a<�a<L�a<��a<�a<��a<��a<��a<��a<E�a<��a<�a<6�a<��a<�a<g�a<��a<�a<��a<ߔa<m�a<��a<�a<��a<�a<d�a<ȗa<V�a<��a<B�a<��a<2�a<��a<�a<��a<؛a<n�a<��a<W�a<ʝa<&�a<��a<�a<��a<�a<��a<�a<Z�a<�a<0�a<��a<�a<w�a<Уa<G�a<��a<�a<}�a<��a<;�a<��a<�a<O�a<s�a<�a<	�a<t�a<��a<�a<<�a<p�a<ĩa<�a<[�a<o�a<��a<۪a<��a<L�a<g�a<��a<��a<ԫa<��a<$�a<S�a<]�a<��a<��a<Ҭa<ݬa<�a<�a<��a<%�a<�a<N�a<N�a<_�a<Y�a<Q�a<��a<`�a<��a<x�a<Y�a<q�a<I�a<X�a<<�a<A�a<%�a<+�a<�a<	�a<�a<ˬa<Ԭa<��a<��a<|�a<Q�a<@�a<��a<�a<��a<��a<{�a<Q�a<D�a<�a<��a<��a<t�a<@�a<��a<̩a<��a<x�a<)�a<�a<��a<p�a<F�a<�a<ҧa<`�a<�a<Цa<��a<:�a<ߥa<��a<4�a<
�a<��a<c�a<��a<��a<N�a<��a<��a<�a<��a<Q�a<Ҡa<~�a<�a<��a<:�a<��a<q�a<��a<��a<�a<Ȝa<:�a<֛a<Y�a<��a<��a<'�a<��a<3�a<�a<o�a<�a<��a<�a<іa<C�a<��a<{�a<�a<��a<Q�a<�a<��a<i�a<�a<��a<;�a<בa<��a<@�a<�a<��a<M�a<
�a<ɏa<��a<A�a<9�a<Ŏa<��a<v�a<9�a<�a<Ѝa<��a<��a<��a<Z�a<E�a<�a<��a<�a<�a<��a<�a<��a<ڌa<��a<ӌa<ƌa<��a<݌a<�a<�a<+�a<U�a<�  �  J�a<u�a<��a<��a<�a<�a<0�a<|�a<��a<�a<�a<K�a<��a<Ǐa<�a<T�a<��a<�a<O�a<��a<�a<R�a<��a<��a<J�a<Ǔa<%�a<�a<̔a<1�a<��a<�a<��a<�a<n�a<חa<R�a<��a<4�a<��a<�a<i�a<�a<�a<�a<^�a<�a<M�a<͝a<M�a<��a<<�a<��a<�a<x�a<�a<\�a<ɡa<5�a<��a<(�a<��a<��a<U�a<��a<�a<d�a<�a<1�a<��a<��a<*�a<��a<ԧa<$�a<v�a<��a<��a<J�a<��a<��a<�a<"�a<T�a<��a<�a<�a<+�a<m�a<��a<ͫa<�a<�a<;�a<G�a<d�a<��a<��a<��a<̬a<�a<�a<$�a<-�a<D�a<9�a<H�a<Z�a<^�a<w�a<i�a<a�a<I�a<p�a<h�a<k�a<^�a<W�a<N�a<?�a<5�a<+�a<�a<�a<ˬa<ʬa<��a<��a<��a<n�a<R�a<%�a<�a<��a<ثa<��a<z�a<J�a<!�a<��a<Ȫa<��a<k�a<J�a<�a<۩a<��a<\�a<2�a<�a<ƨa<��a<8�a<ݧa<��a<q�a<�a<�a<��a<D�a<�a<��a<O�a<��a<��a<J�a<̣a<��a<=�a<�a<q�a<�a<��a<T�a<��a<��a</�a<��a<?�a<Ӟa<k�a<��a<��a<�a<��a<_�a<�a<��a<
�a<��a<+�a<��a<Z�a<�a<n�a<ߗa<��a<-�a<Ŗa<^�a<��a<��a<+�a<ϔa<k�a<��a<��a<0�a<Βa<��a<F�a<��a<��a<F�a<�a<��a<d�a<(�a<��a<��a<H�a<�a<ӎa<��a<e�a<?�a<�a<��a<ƍa<��a<o�a<T�a<A�a<$�a<!�a<��a<�a<��a<یa<Ќa<Ԍa<͌a<ьa<،a<ތa<�a<�a<�a<(�a<�a<�  �  ��a<��a<�a<�a<:�a<{�a<��a<эa<ٍa<?�a<g�a<��a<�a<%�a<��a<��a<�a<N�a<��a<��a<-�a<��a<�a<o�a<��a< �a<d�a<ϓa<E�a<��a<0�a<q�a<��a<F�a<͖a<I�a<��a<#�a<��a<�a<��a<��a<v�a<Śa<y�a<Лa<_�a<֜a<?�a<��a<�a<��a<�a<��a<�a<o�a<�a<<�a<ܡa< �a<��a<�a<]�a<Уa<C�a<��a<�a<l�a<��a<�a<\�a<˦a<�a<I�a<��a<ܧa<E�a<��a<��a<�a<5�a<��a<ϩa<��a<�a<=�a<��a<��a<�a< �a<I�a<S�a<��a<��a<ͫa<�a<��a<3�a<C�a<W�a<|�a<y�a<��a<��a<��a<ˬa<�a<ݬa<֬a<��a<Ȭa<�a<��a<�a<ܬa<�a<Ӭa<Ǭa<Ӭa<��a<��a<��a<��a<��a<{�a<U�a<"�a<*�a<�a<�a<�a<��a<��a<M�a<X�a< �a<�a<تa<��a<��a<@�a<3�a<�a<̩a<��a<;�a<,�a<�a<ƨa<k�a<?�a<�a<��a<t�a<A�a<�a<��a<c�a<��a<��a<y�a<�a<ɤa<p�a<�a<�a<s�a<�a<��a<p�a<�a<��a<A�a<Πa<f�a<�a<��a<�a<ߞa<E�a<�a<}�a<��a<��a<%�a<ԛa<@�a<ךa<u�a<�a<��a<�a<Ϙa< �a<חa<i�a<�a<��a<�a<��a<D�a<��a<��a<�a<ȓa<T�a<�a<��a<M�a<�a<x�a<R�a<�a<��a<X�a<�a<��a<n�a<:�a<�a<a<\�a<?�a<��a<ƍa<��a<_�a<Q�a<��a<��a<׌a<Ča<��a<r�a<u�a<0�a<B�a<A�a<G�a<�a<'�a<�a<�a<2�a<%�a<0�a<[�a<U�a<��a<��a<�  �  ��a<�a<��a<�a<<�a<b�a<��a<Ía<�a<9�a<f�a<��a<ێa<$�a<m�a<��a<��a<L�a<��a<��a<Y�a<��a<�a<W�a<��a<$�a<��a<��a<C�a<��a<�a<��a<��a<j�a<֖a<1�a<Ɨa<5�a<��a<�a<��a<�a<��a<��a<n�a<ߛa<N�a<��a<4�a<��a<,�a<��a<�a<��a<�a<q�a<�a<G�a<��a<'�a<��a<��a<v�a<ţa<&�a<��a<��a<a�a<��a<#�a<P�a<��a<��a<n�a<��a< �a<,�a<|�a<Ϩa<�a<N�a<~�a<��a<�a<J�a<k�a<��a<Ūa<�a<�a<=�a<w�a<��a<��a<Ϋa<�a<�a<'�a<@�a<M�a<n�a<��a<��a<��a<��a<��a<Ȭa<٬a<�a<�a<�a<��a<ܬa<�a<ެa<�a<�a<�a<��a<̬a<��a<��a<��a<}�a<`�a<^�a<[�a<.�a<�a<�a<̫a<��a<��a<y�a<S�a< �a<��a<Ȫa<��a<|�a<J�a<�a<�a<��a<��a<h�a<�a<ިa<��a<x�a<D�a<�a<קa<q�a<+�a<�a<��a<f�a<�a<ƥa<a�a<3�a<ۤa<��a<�a<ˣa<^�a<)�a<̢a<d�a<��a<��a<'�a<àa<q�a< �a<��a<'�a<��a<J�a<�a<�a<�a<��a<,�a<��a<Q�a<�a<i�a<��a<��a<,�a<Řa<X�a<��a<]�a<�a<��a<A�a<͕a<h�a<�a<��a<3�a<ϓa<m�a< �a<��a<E�a<�a<��a<Q�a<��a<��a<D�a<��a<ȏa<o�a<%�a<�a<��a<i�a<2�a<��a<��a<��a<f�a<I�a<�a<�a<ʌa<��a<��a<~�a<o�a<m�a<N�a<%�a<,�a<�a<0�a<0�a<7�a<�a<A�a<L�a<_�a<[�a<u�a<��a<�  �  ��a<ӌa<،a<�a<A�a<n�a<��a<��a<
�a<"�a<p�a<��a<�a<3�a<`�a<ʏa<��a<g�a<��a<�a<\�a<��a<�a<]�a<Œa<�a<m�a<�a<>�a<Ŕa<�a<��a<ܕa<_�a<ۖa<3�a<a<	�a<��a< �a<��a<�a<n�a<�a<F�a<�a<T�a<ۜa<I�a<��a<2�a<��a</�a<��a<�a<j�a<ؠa<]�a<��a<G�a<��a<�a<r�a<ԣa<I�a<��a<	�a<9�a<��a<�a<c�a<ʦa<��a<i�a<��a<��a<1�a<��a<ʨa<�a<U�a<z�a<өa<�a<.�a<U�a<�a<Ѫa<�a<1�a<<�a<v�a<��a<��a<�a<�a< �a<�a<H�a<_�a<r�a<��a<��a<��a<��a<ڬa<٬a<߬a<�a<ͬa<�a<�a<��a<��a<�a<�a<ˬa<�a<��a<Ԭa<��a<��a<��a<��a<y�a<Q�a<F�a<�a<�a<��a<٫a<˫a<��a<~�a<;�a<*�a<�a<Ԫa<��a<n�a<d�a<�a<	�a<��a<��a<k�a<�a<�a<��a<��a<-�a<�a<��a<m�a<G�a<�a<��a<C�a<�a<˥a<c�a<.�a<��a<��a<�a<ߣa<w�a<�a<��a<=�a<�a<��a<F�a<נa<k�a<�a<��a<E�a<��a<`�a<�a<t�a<�a<��a<M�a<��a<W�a<�a<y�a<�a<��a<9�a<��a<G�a<ؗa<p�a<�a<��a<<�a<��a<g�a<�a<��a<-�a<��a<t�a<��a<��a<D�a<��a<��a<2�a<�a<��a<i�a<��a<ȏa<j�a<)�a<�a<��a<��a<%�a<�a<΍a<��a<w�a<0�a<$�a<�a<�a<��a<��a<��a<L�a<[�a<>�a<?�a<:�a<%�a<!�a<�a<9�a<�a<I�a<4�a<H�a<j�a<�a<��a<�  �  ��a<Ȍa<�a< �a<9�a<Z�a<��a<ȍa<��a<5�a<g�a<��a<�a<)�a<p�a<��a< �a<M�a<��a<��a<J�a<��a<��a<G�a<��a< �a<��a<ݓa<D�a<��a<�a<��a<��a<]�a<Ζa<P�a<��a<'�a<��a<�a<��a<�a<q�a<�a<v�a<ߛa<B�a<��a<7�a<��a<4�a<��a<�a<��a<��a<j�a<ܠa<M�a<��a<'�a<��a<
�a<h�a<ɣa</�a<��a<��a<c�a<��a<�a<d�a<��a<��a<d�a<��a<�a<E�a<��a<��a<�a<J�a<~�a<��a<��a<*�a<k�a<��a<Ūa<ܪa<�a<@�a<h�a<��a<��a<ͫa<�a<�a<(�a<A�a<^�a<d�a<��a<��a<��a<��a<��a<ìa<Ьa<�a<��a<�a<�a<�a<�a<�a<��a<ڬa<άa<۬a<��a<��a<��a<��a<|�a<n�a<[�a<;�a<>�a<�a<�a<īa<��a<��a<o�a<N�a<!�a<��a<תa<��a<�a<Q�a< �a<�a<��a<��a<Y�a<!�a<�a<��a<w�a<?�a<	�a<��a<s�a<3�a<�a<��a<^�a<
�a<��a<��a<�a<Τa<��a<�a<ȣa<x�a<�a<��a<l�a<��a<��a<,�a<Ơa<i�a<�a<��a<+�a<��a<T�a<�a<x�a<�a<��a<-�a<a<\�a<�a<n�a< �a<��a<+�a<Ƙa<P�a<֗a<q�a<��a<��a<8�a<ŕa<T�a<��a<��a<#�a<˓a<i�a<�a<��a<J�a<�a<��a<M�a<��a<��a<M�a<�a<��a<}�a<-�a<�a<��a<o�a<3�a<��a<͍a<��a<g�a<?�a<�a<��a<Ȍa<��a<��a<��a<{�a<N�a<G�a<;�a<&�a<&�a<2�a<�a<�a<:�a<.�a<?�a<]�a<e�a<t�a<��a<�  �  Ōa<a<�a<�a<U�a<}�a<��a<эa<�a<C�a<k�a<��a<�a<�a<~�a<��a<�a<G�a<��a<��a<;�a<��a<��a<r�a<͒a<�a<z�a<ޓa<X�a<��a<%�a<t�a<�a<d�a<Ėa<P�a<��a<9�a<��a< �a<}�a<��a<��a<�a<a�a<Λa<j�a<ќa<G�a<��a<!�a<��a<�a<��a<��a<n�a<�a<C�a<֡a<�a<��a<��a<i�a<ףa<7�a<��a<�a<M�a<��a<�a<e�a<��a<�a<E�a<��a<ާa<?�a<z�a<��a<�a<1�a<��a<��a<�a<-�a<]�a<��a<ͪa<�a<�a<M�a<^�a<��a<��a<ëa<�a<��a<9�a<7�a<_�a<w�a<��a<��a<��a<¬a<Ŭa<�a<�a<Ѭa<�a<߬a<�a<�a<�a<�a<٬a<�a<¬a<٬a<��a<��a<��a<��a<��a<_�a<n�a<5�a<*�a<��a<	�a<�a<��a<��a<\�a<\�a<%�a<��a<ުa<��a<��a<=�a<4�a<�a<éa<��a<J�a</�a<�a<ɨa<��a<,�a<��a<��a<��a<#�a<��a<��a<Z�a<�a<��a<�a<
�a<ߤa<h�a<2�a<��a<p�a<$�a<��a<X�a<�a<��a<<�a<֠a<j�a<��a<��a<!�a<՞a<P�a<�a<��a<�a<��a<!�a<ϛa<K�a<�a<|�a<�a<��a<"�a<��a<A�a<�a<r�a<��a<��a<�a<ҕa<F�a<��a<��a<$�a<̓a<P�a<�a<��a<Y�a<��a<��a<<�a<��a<��a<L�a<�a<��a<u�a<2�a<܎a<��a<^�a<E�a<�a<΍a<��a<g�a<R�a<�a<��a<ьa<Ča<��a<l�a<j�a<G�a<Y�a<,�a<+�a<*�a<�a<1�a<�a<9�a<!�a<M�a<I�a<_�a<|�a<��a<�  �  ��a<Όa<��a<�a<4�a<]�a<��a<��a< �a<5�a<m�a<��a<�a<*�a<w�a<��a<��a<O�a<��a<��a<N�a<��a<	�a<P�a<��a<�a<��a<ݓa<J�a<��a<�a<��a<�a<i�a<̖a<9�a<��a<*�a<��a<�a<��a<�a<j�a<��a<f�a<�a<H�a<��a<H�a<��a<2�a<��a<�a<��a<��a<r�a<�a<O�a<��a<!�a<��a<�a<j�a<գa<2�a<��a<��a<V�a<��a<�a<i�a<��a<�a<O�a<��a<�a<3�a<{�a<˨a< �a<H�a<��a<��a<��a<'�a<t�a<��a<��a<�a<"�a<@�a<n�a<��a<��a<˫a<�a<�a<3�a<A�a<[�a<i�a<��a<��a<��a<��a<Ԭa<Ĭa<Ӭa<�a<�a<�a<�a<��a<�a<�a<լa<�a<Ԭa<��a<¬a<��a<��a<��a<��a<v�a<R�a<A�a<6�a<�a<�a<ȫa<ëa<��a<u�a<N�a<'�a<��a<Ӫa<��a<��a<P�a<�a<�a<ɩa<��a<]�a<!�a<��a<��a<p�a<:�a<�a<��a<y�a<6�a<�a<��a<Q�a<�a<��a<i�a<�a<Фa<j�a<.�a<ʣa<y�a<�a<Ƣa<]�a<�a<��a<+�a<נa<d�a<�a<��a<%�a<��a<X�a<�a<��a<�a<��a<&�a<Лa<U�a<�a<y�a<�a<��a<-�a<��a<Z�a<՗a<v�a<�a<��a<"�a<��a<W�a<�a<��a</�a<��a<g�a<�a<��a<P�a<�a<��a<G�a<�a<��a<Z�a<�a<��a<s�a<9�a<�a<��a<n�a<?�a<��a<ʍa<��a<h�a<H�a<�a<�a<ߌa<��a<��a<��a<r�a<W�a<9�a<@�a<2�a<0�a<�a<(�a<$�a<�a<6�a<F�a<B�a<n�a<}�a<��a<�  �  ��a<��a<�a<�a<:�a<d�a<��a<��a<�a<�a<p�a<��a<�a<:�a<b�a<Ώa<��a<U�a<��a<�a<d�a<��a<�a<M�a<��a<�a<~�a<�a<8�a<Ŕa<�a<��a<�a<i�a<Җa<4�a<ȗa<�a<��a<	�a<~�a<�a<^�a<�a<R�a<�a<C�a<؜a<?�a<��a<5�a<��a<!�a<}�a<�a<p�a<ߠa<f�a<��a<6�a<��a<�a<l�a<ǣa<I�a<��a<�a<D�a<ƥa<��a<e�a<��a<��a<\�a<��a<�a<2�a<}�a<Шa<��a<M�a<l�a<ɩa<�a<,�a<k�a<��a<ƪa<�a<6�a<-�a<}�a<��a<��a<֫a<�a<'�a<�a<L�a<e�a<h�a<��a<��a<Ĭa<��a<άa<Ѭa<Ӭa<�a<ܬa<�a<֬a<�a<جa<�a<�a<լa<�a<��a<ͬa<��a<��a<��a<i�a<��a<A�a<S�a<!�a<
�a<�a<ϫa<īa<~�a<��a<5�a<*�a<��a<תa<��a<q�a<g�a<�a<��a<��a<�a<s�a<�a<�a<��a<u�a<.�a<��a<��a<g�a<G�a<զa<��a<K�a<�a<��a<d�a<5�a<Ĥa<z�a<�a<£a<��a<��a<Ӣa<I�a<�a<��a<C�a<͠a<d�a<	�a<��a<8�a<��a<h�a<�a<{�a<$�a<��a<<�a<��a<T�a<�a<k�a<�a<��a<3�a<��a<_�a<̗a<s�a<��a<��a<0�a<��a<k�a<�a<��a<4�a<��a<l�a<�a<��a<B�a<�a<��a<8�a<��a<��a<n�a<�a<Ϗa<j�a<*�a<��a<��a<��a<+�a<�a<ԍa<��a<s�a<,�a<3�a<�a<ڌa<��a<��a<{�a<[�a<k�a<,�a<P�a<�a<"�a<"�a<�a<4�a<�a<B�a<=�a<L�a<c�a<a�a<��a<�  �  ��a<ڌa<�a<�a<A�a<x�a<��a<ōa<�a<8�a<{�a<��a<�a<1�a<j�a<��a<�a<E�a<��a<��a<W�a<��a<�a<d�a<Ēa<�a<n�a<�a<A�a<��a< �a<|�a<�a<[�a<Ȗa<G�a<��a<�a<��a<�a<��a< �a<p�a<�a<X�a<ۛa<S�a<ޜa<=�a<��a</�a<��a<�a<��a<�a<o�a<�a<U�a<��a<)�a<��a<�a<u�a<ͣa<G�a<��a<��a<H�a<��a<
�a<`�a<��a<�a<G�a<��a<�a<=�a<|�a<��a<��a<:�a<��a<��a<�a<6�a<U�a<��a<˪a<��a<&�a<;�a<u�a<��a<��a<ƫa<��a<�a<%�a<E�a<g�a<k�a<��a<��a<��a<��a<Ĭa<�a<ݬa<ڬa<ެa<��a<�a<�a<�a<�a<ެa<֬a<Ѭa<Ϭa<��a<��a<��a<��a<�a<p�a<P�a<M�a<�a<�a<��a<�a<��a<��a<z�a<R�a<5�a<��a<ުa<��a<x�a<T�a<-�a<�a<ϩa<��a<e�a<�a<�a<��a<��a<1�a<�a<ça<p�a<5�a<�a<��a<M�a<�a<��a<v�a<�a<��a<k�a<+�a<ɣa<t�a<�a<��a<O�a<��a<��a<I�a<̠a<p�a<�a<��a<0�a<��a<`�a<�a<|�a<�a<��a</�a<̛a<V�a<�a<q�a<�a<��a<,�a<��a<H�a<ܗa<n�a<��a<��a<�a<��a<R�a<��a<��a<%�a<��a<Y�a<�a<��a<E�a<��a<��a<=�a<��a<��a<^�a<��a<Əa<v�a<>�a<��a<��a<q�a<1�a< �a<֍a<��a<y�a<C�a< �a<��a<όa<Ìa<��a<u�a<]�a<_�a<?�a<8�a<(�a<+�a<�a<�a<!�a<.�a<1�a<;�a<H�a<d�a<x�a<��a<�  �  ��a<Ōa<�a<,�a<-�a<i�a<��a<ލa<�a<;�a<g�a<��a<��a<�a<��a<��a<�a<H�a<��a<��a<E�a<��a<��a<^�a<��a<0�a<��a<��a<M�a<��a<'�a<y�a<��a<]�a<��a<L�a<��a<:�a<��a<�a<��a<�a<z�a<�a<}�a<�a<G�a<Ɯa<D�a<a<%�a<��a<�a<��a<��a<p�a<�a<E�a<ҡa<�a<��a<��a<r�a<أa</�a<��a<��a<o�a<��a<�a<\�a<��a<�a<B�a<��a<ݧa<>�a<v�a<��a<�a<7�a<��a<��a<��a<0�a<j�a<��a<��a<�a<�a<U�a<i�a<��a<��a<ƫa<�a<��a<>�a<:�a<f�a<s�a<|�a<��a<��a<ͬa<¬a<Ьa<ͬa<��a<��a<�a<��a<ڬa<��a<�a<جa<�a<��a<Ԭa<��a<��a<��a<��a<��a<W�a<`�a<8�a<=�a<%�a<�a<ԫa<��a<��a<b�a<U�a<!�a<��a<�a<��a<��a<B�a<7�a<�a<ͩa<��a<T�a<9�a<�a<��a<e�a<O�a<�a<��a<|�a<�a<��a<��a<^�a<�a<��a<|�a<�a<�a<c�a<$�a<ǣa<e�a<�a<��a<t�a< �a<��a<0�a<Ӡa<t�a<��a<��a<�a<Оa<Q�a<�a<��a<�a<��a<"�a<ڛa<M�a<�a<}�a< �a<��a<%�a<Ҙa<H�a<�a<i�a<��a<��a<�a<֕a<F�a<��a<��a< �a<ѓa<V�a<�a<��a<M�a<��a<��a<\�a<�a<��a<I�a<�a<��a<m�a<>�a<ߎa<a<^�a<I�a<��a<Սa<��a<a�a<M�a<�a<�a<Όa<��a<��a<��a<~�a<J�a<L�a<#�a<7�a<%�a<�a</�a<�a<4�a< �a<H�a<I�a<a�a<��a<|�a<�  �  ��a<Ɍa<ߌa<�a<H�a<}�a<��a<ˍa<��a<1�a<r�a<��a<�a<'�a<��a<��a<�a<f�a<��a<�a<S�a<��a<��a<o�a<��a<�a<o�a<Փa<G�a<��a<�a<}�a<�a<_�a<Ȗa<:�a<��a< �a<��a<�a<��a<��a<o�a<�a<O�a<ޛa<Z�a<Ԝa<?�a<��a<.�a<��a<!�a<��a<��a<z�a<�a<P�a<ȡa<:�a<��a<�a<n�a<̣a<>�a<��a<��a<B�a<��a<�a<]�a<��a<�a<N�a<��a<�a<1�a<v�a<��a<��a<?�a<~�a<��a<��a<!�a<W�a<��a<ƪa<�a<�a<B�a<s�a<��a<��a<�a<��a<	�a<>�a<C�a<\�a<{�a<��a<��a<��a<��a<Ĭa<�a<�a<�a<լa<�a<�a<�a<�a<�a<۬a<׬a<Ьa<Ȭa<��a<��a<��a<��a<��a<i�a<W�a<<�a<�a<�a<��a<�a<��a<��a<q�a<J�a<+�a<�a<תa<��a<��a<O�a<#�a<�a<©a<��a<b�a<&�a<�a<ƨa<|�a<+�a<�a<��a<v�a<0�a<�a<��a<H�a<�a<��a<i�a<�a<Ƥa<p�a<�a<ңa<n�a<�a<��a<F�a<��a<��a<?�a<Πa<j�a<�a<��a<8�a<̞a<T�a<��a<��a<�a<��a<@�a<��a<T�a<�a<q�a<�a<��a<*�a<��a<E�a<ԗa<k�a<�a<��a<!�a<��a<R�a<�a<��a<#�a<��a<^�a<�a<��a<K�a<�a<��a<6�a<��a<��a<T�a<�a<ďa<s�a<*�a< �a<��a<j�a<J�a<��a<ˍa<��a<t�a<A�a<�a<�a<όa<Ōa<��a<}�a<U�a<P�a<A�a<3�a<3�a<!�a<�a<�a< �a<(�a</�a<>�a<E�a<\�a<z�a<��a<�  �  ��a<�a<�a<�a<>�a<T�a<��a<Ía<�a<9�a<z�a<��a<�a<A�a<c�a<яa<�a<X�a<��a<�a<U�a<��a<�a<>�a<ɒa<�a<��a<�a<?�a<��a<�a<��a<�a<b�a<̖a<-�a<��a<�a<��a<�a<�a<�a<m�a<�a<`�a<�a<=�a<��a<B�a<��a<D�a<��a<*�a<r�a<
�a<v�a<�a<b�a<��a<@�a<��a<�a<l�a<Уa<1�a<}�a<	�a<R�a<ƥa<�a<g�a<��a<��a<p�a<��a<��a<*�a<w�a<Ȩa<��a<W�a<n�a<��a<��a<6�a<o�a<��a<ժa<Ӫa<!�a<>�a<r�a<��a<��a<�a<ګa<"�a<�a<U�a<[�a<b�a<��a<��a<��a<��a<ʬa<��a<Ӭa<�a<�a<�a<ݬa<��a<۬a<�a<�a<Ѭa<�a<��a<Ȭa<��a<��a<��a<o�a<z�a<F�a<W�a<,�a<�a<�a<��a<��a<��a<��a<R�a<3�a<��a<Ϫa<��a<r�a<j�a<�a<��a<��a<��a<c�a<�a<�a<��a<��a<<�a<�a<ʧa<m�a<7�a<֦a<��a<R�a<�a<��a<]�a<-�a<��a<��a<�a<ãa<y�a<�a<΢a<W�a<	�a<��a<+�a<Ѡa<c�a<�a<��a<A�a<��a<c�a<�a<|�a< �a<��a<F�a<��a<k�a<�a<t�a<�a<}�a<9�a<��a<_�a<ڗa<t�a< �a<��a<C�a<��a<c�a<�a<��a<+�a<��a<v�a<�a<��a<J�a<��a<��a<H�a<�a<��a<Y�a<�a<Ïa<��a<"�a<��a<��a<��a<*�a<�a<ʍa<��a<�a<C�a</�a<�a<֌a<��a<��a<��a<j�a<k�a<3�a<F�a<�a< �a<2�a<�a<2�a<�a<<�a<:�a<W�a<a�a<g�a<��a<�  �  ��a<��a<�a<�a<E�a<o�a<��a<͍a<�a<1�a<h�a<��a<��a<:�a<a�a<яa<�a<c�a<��a<��a<;�a<��a<�a<d�a<��a<�a<q�a<ؓa<E�a<��a<�a<}�a<�a<N�a<˖a<<�a<��a<�a<��a<�a<��a<�a<k�a<ݚa<_�a<ޛa<`�a<֜a<_�a<��a<.�a<��a<'�a<��a<�a<m�a<٠a<b�a<͡a<C�a<��a<�a<]�a<�a<D�a<��a<��a<P�a<��a<��a<j�a<��a<��a<N�a<��a<�a<7�a<|�a<��a< �a<<�a<��a<��a<��a<�a<T�a<��a<ƪa<��a<2�a<V�a<Y�a<��a<��a<�a<�a<'�a<�a<Q�a<j�a<��a<��a<��a<��a<��a<�a<٬a<�a<�a<�a<ݬa<�a<��a<�a<ެa<۬a<Ϭa<ɬa<ìa<��a<��a<��a<��a<��a<v�a<Q�a<2�a<!�a<�a<��a<ګa<Ыa<��a<h�a<J�a<!�a<�a<�a<��a<p�a<j�a<5�a<�a<��a<��a<I�a<1�a<�a<��a<y�a<8�a<�a<��a<s�a<3�a<�a<��a<R�a<��a<��a<k�a<�a<��a<p�a<�a<ģa<{�a<�a<��a<V�a<��a<��a<A�a<�a<a�a<�a<��a<=�a<Ϟa<f�a<�a<u�a< �a<��a<I�a<��a<W�a<ךa<��a<�a<��a<+�a<��a<:�a<Ηa<x�a<��a<��a<"�a<��a<L�a<�a<��a<�a<��a<[�a<�a<��a<Q�a<�a<��a<C�a<��a<��a<i�a<�a<��a<w�a<$�a<�a<��a<��a<(�a<�a<ٍa<��a<l�a<?�a<�a<�a<��a<��a<��a<~�a<c�a<E�a<=�a<B�a<,�a<�a<�a<�a<�a<#�a<)�a<0�a<H�a<Z�a<|�a<��a<�  �  ��a<ӌa<�a<�a<?�a<e�a<�a<ƍa<�a<Q�a<_�a<��a<׎a< �a<z�a<��a< �a<V�a<��a<�a<V�a<��a<ڑa<j�a<��a<�a<��a<�a<E�a<��a<)�a<t�a<��a<U�a<͖a<C�a<��a<:�a<��a<�a<z�a<�a<x�a<�a<y�a<ϛa<b�a<��a<5�a<��a<@�a<��a<
�a<��a<�a<|�a<�a<>�a<¡a<!�a<��a<�a<g�a<ʣa<�a<��a<�a<i�a<��a<
�a<N�a<��a<�a<I�a<��a<֧a<8�a<|�a<��a<�a<3�a<��a<��a<��a<*�a<m�a<��a<��a<�a<��a<E�a<p�a<��a<��a<ѫa<�a<�a<4�a<A�a<F�a<��a<t�a<��a<��a<��a<��a<��a<߬a<٬a<��a<�a<��a<ʬa<�a<�a<ެa<�a<��a<ڬa<��a<��a<��a<��a<��a<I�a<d�a<F�a<:�a<�a<�a<Ыa<��a<��a<��a<k�a<�a<�a<Īa<��a<��a<I�a<�a<��a<��a<��a<d�a<$�a<Ǩa<¨a<g�a<=�a<	�a<��a<t�a<�a<��a<��a<e�a<�a<��a<s�a<�a<�a<n�a<,�a<��a<Z�a<�a<��a<p�a<�a<��a<�a<Ġa<j�a<�a<��a<!�a<Ȟa<B�a<��a<��a<��a<��a<'�a<ƛa<j�a<�a<o�a<ޙa<��a<�a<̘a<V�a<ۗa<[�a<�a<��a<�a<ٕa<>�a<�a<��a<�a<ړa<R�a<�a<��a<K�a<�a<��a<O�a<�a<��a<-�a<�a<a<��a<'�a<�a<��a<f�a<?�a<��a<��a<��a<Z�a<]�a<*�a<�a<��a<��a<��a<t�a<{�a<Y�a<N�a<�a<.�a<+�a<�a<+�a<�a<:�a<)�a<D�a<O�a<`�a<��a<n�a<�  �  ��a<��a<�a<�a<E�a<o�a<��a<͍a<�a<1�a<h�a<��a<��a<:�a<a�a<яa<�a<c�a<��a<��a<;�a<��a<�a<d�a<��a<�a<q�a<ؓa<E�a<��a<�a<}�a<�a<N�a<˖a<<�a<��a<�a<��a<�a<��a<�a<k�a<ݚa<_�a<ޛa<`�a<֜a<_�a<��a<.�a<��a<'�a<��a<�a<m�a<٠a<b�a<͡a<C�a<��a<�a<]�a<�a<D�a<��a<��a<P�a<��a<��a<j�a<��a<��a<N�a<��a<�a<7�a<|�a<��a< �a<<�a<��a<��a<��a<�a<T�a<��a<ƪa<��a<2�a<V�a<Y�a<��a<��a<�a<�a<'�a<�a<Q�a<j�a<��a<��a<��a<��a<��a<�a<٬a<�a<�a<�a<ݬa<�a<��a<�a<ެa<۬a<Ϭa<ɬa<ìa<��a<��a<��a<��a<��a<v�a<Q�a<2�a<!�a<�a<��a<ګa<Ыa<��a<h�a<J�a<!�a<�a<�a<��a<p�a<j�a<5�a<�a<��a<��a<I�a<1�a<�a<��a<y�a<8�a<�a<��a<s�a<3�a<�a<��a<R�a<��a<��a<k�a<�a<��a<p�a<�a<ģa<{�a<�a<��a<V�a<��a<��a<A�a<�a<a�a<�a<��a<=�a<Ϟa<f�a<�a<u�a< �a<��a<I�a<��a<W�a<ךa<��a<�a<��a<+�a<��a<:�a<Ηa<x�a<��a<��a<"�a<��a<L�a<�a<��a<�a<��a<[�a<�a<��a<Q�a<�a<��a<C�a<��a<��a<i�a<�a<��a<w�a<$�a<�a<��a<��a<(�a<�a<ٍa<��a<l�a<?�a<�a<�a<��a<��a<��a<~�a<c�a<E�a<=�a<B�a<,�a<�a<�a<�a<�a<#�a<)�a<0�a<H�a<Z�a<|�a<��a<�  �  ��a<�a<�a<�a<>�a<T�a<��a<Ía<�a<9�a<z�a<��a<�a<A�a<c�a<яa<�a<X�a<��a<�a<U�a<��a<�a<>�a<ɒa<�a<��a<�a<?�a<��a<�a<��a<�a<b�a<̖a<-�a<��a<�a<��a<�a<�a<�a<m�a<�a<`�a<�a<=�a<��a<B�a<��a<D�a<��a<*�a<r�a<
�a<v�a<�a<b�a<��a<@�a<��a<�a<l�a<Уa<1�a<}�a<	�a<R�a<ƥa<�a<g�a<��a<��a<p�a<��a<��a<*�a<w�a<Ȩa<��a<W�a<n�a<��a<��a<6�a<o�a<��a<ժa<Ӫa<!�a<>�a<r�a<��a<��a<�a<ګa<"�a<�a<U�a<[�a<b�a<��a<��a<��a<��a<ʬa<��a<Ӭa<�a<�a<�a<ݬa<��a<۬a<�a<�a<Ѭa<�a<��a<Ȭa<��a<��a<��a<o�a<z�a<F�a<W�a<,�a<�a<�a<��a<��a<��a<��a<R�a<3�a<��a<Ϫa<��a<r�a<j�a<�a<��a<��a<��a<c�a<�a<�a<��a<��a<<�a<�a<ʧa<m�a<7�a<֦a<��a<R�a<�a<��a<]�a<-�a<��a<��a<�a<ãa<y�a<�a<΢a<W�a<	�a<��a<+�a<Ѡa<c�a<�a<��a<A�a<��a<c�a<�a<|�a< �a<��a<F�a<��a<k�a<�a<t�a<�a<}�a<9�a<��a<_�a<ڗa<t�a< �a<��a<C�a<��a<c�a<�a<��a<+�a<��a<v�a<�a<��a<J�a<��a<��a<H�a<�a<��a<Y�a<�a<Ïa<��a<"�a<��a<��a<��a<*�a<�a<ʍa<��a<�a<C�a</�a<�a<֌a<��a<��a<��a<j�a<k�a<3�a<F�a<�a< �a<2�a<�a<2�a<�a<<�a<:�a<W�a<a�a<g�a<��a<�  �  ��a<Ɍa<ߌa<�a<H�a<}�a<��a<ˍa<��a<1�a<r�a<��a<�a<'�a<��a<��a<�a<f�a<��a<�a<S�a<��a<��a<o�a<��a<�a<o�a<Փa<G�a<��a<�a<}�a<�a<_�a<Ȗa<:�a<��a< �a<��a<�a<��a<��a<o�a<�a<O�a<ޛa<Z�a<Ԝa<?�a<��a<.�a<��a<!�a<��a<��a<z�a<�a<P�a<ȡa<:�a<��a<�a<n�a<̣a<>�a<��a<��a<B�a<��a<�a<]�a<��a<�a<N�a<��a<�a<1�a<v�a<��a<��a<?�a<~�a<��a<��a<!�a<W�a<��a<ƪa<�a<�a<B�a<s�a<��a<��a<�a<��a<	�a<>�a<C�a<\�a<{�a<��a<��a<��a<��a<Ĭa<�a<�a<�a<լa<�a<�a<�a<�a<�a<۬a<׬a<Ьa<Ȭa<��a<��a<��a<��a<��a<i�a<W�a<<�a<�a<�a<��a<�a<��a<��a<q�a<J�a<+�a<�a<תa<��a<��a<O�a<#�a<�a<©a<��a<b�a<&�a<�a<ƨa<|�a<+�a<�a<��a<v�a<0�a<�a<��a<H�a<�a<��a<i�a<�a<Ƥa<p�a<�a<ңa<n�a<�a<��a<F�a<��a<��a<?�a<Πa<j�a<�a<��a<8�a<̞a<T�a<��a<��a<�a<��a<@�a<��a<T�a<�a<q�a<�a<��a<*�a<��a<E�a<ԗa<k�a<�a<��a<!�a<��a<R�a<�a<��a<#�a<��a<^�a<�a<��a<K�a<�a<��a<6�a<��a<��a<T�a<�a<ďa<s�a<*�a< �a<��a<j�a<J�a<��a<ˍa<��a<t�a<A�a<�a<�a<όa<Ōa<��a<}�a<U�a<P�a<A�a<3�a<3�a<!�a<�a<�a< �a<(�a</�a<>�a<E�a<\�a<z�a<��a<�  �  ��a<Ōa<�a<,�a<-�a<i�a<��a<ލa<�a<;�a<g�a<��a<��a<�a<��a<��a<�a<H�a<��a<��a<E�a<��a<��a<^�a<��a<0�a<��a<��a<M�a<��a<'�a<y�a<��a<]�a<��a<L�a<��a<:�a<��a<�a<��a<�a<z�a<�a<}�a<�a<G�a<Ɯa<D�a<a<%�a<��a<�a<��a<��a<p�a<�a<E�a<ҡa<�a<��a<��a<r�a<أa</�a<��a<��a<o�a<��a<�a<\�a<��a<�a<B�a<��a<ݧa<>�a<v�a<��a<�a<7�a<��a<��a<��a<0�a<j�a<��a<��a<�a<�a<U�a<i�a<��a<��a<ƫa<�a<��a<>�a<:�a<f�a<s�a<|�a<��a<��a<ͬa<¬a<Ьa<ͬa<��a<��a<�a<��a<ڬa<��a<�a<جa<�a<��a<Ԭa<��a<��a<��a<��a<��a<W�a<`�a<8�a<=�a<%�a<�a<ԫa<��a<��a<b�a<U�a<!�a<��a<�a<��a<��a<B�a<7�a<�a<ͩa<��a<T�a<9�a<�a<��a<e�a<O�a<�a<��a<|�a<�a<��a<��a<^�a<�a<��a<|�a<�a<�a<c�a<$�a<ǣa<e�a<�a<��a<t�a< �a<��a<0�a<Ӡa<t�a<��a<��a<�a<Оa<Q�a<�a<��a<�a<��a<"�a<ڛa<M�a<�a<}�a< �a<��a<%�a<Ҙa<H�a<�a<i�a<��a<��a<�a<֕a<F�a<��a<��a< �a<ѓa<V�a<�a<��a<M�a<��a<��a<\�a<�a<��a<I�a<�a<��a<m�a<>�a<ߎa<a<^�a<I�a<��a<Սa<��a<a�a<M�a<�a<�a<Όa<��a<��a<��a<~�a<J�a<L�a<#�a<7�a<%�a<�a</�a<�a<4�a< �a<H�a<I�a<a�a<��a<|�a<�  �  ��a<ڌa<�a<�a<A�a<x�a<��a<ōa<�a<8�a<{�a<��a<�a<1�a<j�a<��a<�a<E�a<��a<��a<W�a<��a<�a<d�a<Ēa<�a<n�a<�a<A�a<��a< �a<|�a<�a<[�a<Ȗa<G�a<��a<�a<��a<�a<��a< �a<p�a<�a<X�a<ۛa<S�a<ޜa<=�a<��a</�a<��a<�a<��a<�a<o�a<�a<U�a<��a<)�a<��a<�a<u�a<ͣa<G�a<��a<��a<H�a<��a<
�a<`�a<��a<�a<G�a<��a<�a<=�a<|�a<��a<��a<:�a<��a<��a<�a<6�a<U�a<��a<˪a<��a<&�a<;�a<u�a<��a<��a<ƫa<��a<�a<%�a<E�a<g�a<k�a<��a<��a<��a<��a<Ĭa<�a<ݬa<ڬa<ެa<��a<�a<�a<�a<�a<ެa<֬a<Ѭa<Ϭa<��a<��a<��a<��a<�a<p�a<P�a<M�a<�a<�a<��a<�a<��a<��a<z�a<R�a<5�a<��a<ުa<��a<x�a<T�a<-�a<�a<ϩa<��a<e�a<�a<�a<��a<��a<1�a<�a<ça<p�a<5�a<�a<��a<M�a<�a<��a<v�a<�a<��a<k�a<+�a<ɣa<t�a<�a<��a<O�a<��a<��a<I�a<̠a<p�a<�a<��a<0�a<��a<`�a<�a<|�a<�a<��a</�a<̛a<V�a<�a<q�a<�a<��a<,�a<��a<H�a<ܗa<n�a<��a<��a<�a<��a<R�a<��a<��a<%�a<��a<Y�a<�a<��a<E�a<��a<��a<=�a<��a<��a<^�a<��a<Əa<v�a<>�a<��a<��a<q�a<1�a< �a<֍a<��a<y�a<C�a< �a<��a<όa<Ìa<��a<u�a<]�a<_�a<?�a<8�a<(�a<+�a<�a<�a<!�a<.�a<1�a<;�a<H�a<d�a<x�a<��a<�  �  ��a<��a<�a<�a<:�a<d�a<��a<��a<�a<�a<p�a<��a<�a<:�a<b�a<Ώa<��a<U�a<��a<�a<d�a<��a<�a<M�a<��a<�a<~�a<�a<8�a<Ŕa<�a<��a<�a<i�a<Җa<4�a<ȗa<�a<��a<	�a<~�a<�a<^�a<�a<R�a<�a<C�a<؜a<?�a<��a<5�a<��a<!�a<}�a<�a<p�a<ߠa<f�a<��a<6�a<��a<�a<l�a<ǣa<I�a<��a<�a<D�a<ƥa<��a<e�a<��a<��a<\�a<��a<�a<2�a<}�a<Шa<��a<M�a<l�a<ɩa<�a<,�a<k�a<��a<ƪa<�a<6�a<-�a<}�a<��a<��a<֫a<�a<'�a<�a<L�a<e�a<h�a<��a<��a<Ĭa<��a<άa<Ѭa<Ӭa<�a<ܬa<�a<֬a<�a<جa<�a<�a<լa<�a<��a<ͬa<��a<��a<��a<i�a<��a<A�a<S�a<!�a<
�a<�a<ϫa<īa<~�a<��a<5�a<*�a<��a<תa<��a<q�a<g�a<�a<��a<��a<�a<s�a<�a<�a<��a<u�a<.�a<��a<��a<g�a<G�a<զa<��a<K�a<�a<��a<d�a<5�a<Ĥa<z�a<�a<£a<��a<��a<Ӣa<I�a<�a<��a<C�a<͠a<d�a<	�a<��a<8�a<��a<h�a<�a<{�a<$�a<��a<<�a<��a<T�a<�a<k�a<�a<��a<3�a<��a<_�a<̗a<s�a<��a<��a<0�a<��a<k�a<�a<��a<4�a<��a<l�a<�a<��a<B�a<�a<��a<8�a<��a<��a<n�a<�a<Ϗa<j�a<*�a<��a<��a<��a<+�a<�a<ԍa<��a<s�a<,�a<3�a<�a<ڌa<��a<��a<{�a<[�a<k�a<,�a<P�a<�a<"�a<"�a<�a<4�a<�a<B�a<=�a<L�a<c�a<a�a<��a<�  �  ��a<Όa<��a<�a<4�a<]�a<��a<��a< �a<5�a<m�a<��a<�a<*�a<w�a<��a<��a<O�a<��a<��a<N�a<��a<	�a<P�a<��a<�a<��a<ݓa<J�a<��a<�a<��a<�a<i�a<̖a<9�a<��a<*�a<��a<�a<��a<�a<j�a<��a<f�a<�a<H�a<��a<H�a<��a<2�a<��a<�a<��a<��a<r�a<�a<O�a<��a<!�a<��a<�a<j�a<գa<2�a<��a<��a<V�a<��a<�a<i�a<��a<�a<O�a<��a<�a<3�a<{�a<˨a< �a<H�a<��a<��a<��a<'�a<t�a<��a<��a<�a<"�a<@�a<n�a<��a<��a<˫a<�a<�a<3�a<A�a<[�a<i�a<��a<��a<��a<��a<Ԭa<Ĭa<Ӭa<�a<�a<�a<�a<��a<�a<�a<լa<�a<Ԭa<��a<¬a<��a<��a<��a<��a<v�a<R�a<A�a<6�a<�a<�a<ȫa<ëa<��a<u�a<N�a<'�a<��a<Ӫa<��a<��a<P�a<�a<�a<ɩa<��a<]�a<!�a<��a<��a<p�a<:�a<�a<��a<y�a<6�a<�a<��a<Q�a<�a<��a<i�a<�a<Фa<j�a<.�a<ʣa<y�a<�a<Ƣa<]�a<�a<��a<+�a<נa<d�a<�a<��a<%�a<��a<X�a<�a<��a<�a<��a<&�a<Лa<U�a<�a<y�a<�a<��a<-�a<��a<Z�a<՗a<v�a<�a<��a<"�a<��a<W�a<�a<��a</�a<��a<g�a<�a<��a<P�a<�a<��a<G�a<�a<��a<Z�a<�a<��a<s�a<9�a<�a<��a<n�a<?�a<��a<ʍa<��a<h�a<H�a<�a<�a<ߌa<��a<��a<��a<r�a<W�a<9�a<@�a<2�a<0�a<�a<(�a<$�a<�a<6�a<F�a<B�a<n�a<}�a<��a<�  �  Ōa<a<�a<�a<U�a<}�a<��a<эa<�a<C�a<k�a<��a<�a<�a<~�a<��a<�a<G�a<��a<��a<;�a<��a<��a<r�a<͒a<�a<z�a<ޓa<X�a<��a<%�a<t�a<�a<d�a<Ėa<P�a<��a<9�a<��a< �a<}�a<��a<��a<�a<a�a<Λa<j�a<ќa<G�a<��a<!�a<��a<�a<��a<��a<n�a<�a<C�a<֡a<�a<��a<��a<i�a<ףa<7�a<��a<�a<M�a<��a<�a<e�a<��a<�a<E�a<��a<ާa<?�a<z�a<��a<�a<1�a<��a<��a<�a<-�a<]�a<��a<ͪa<�a<�a<M�a<^�a<��a<��a<ëa<�a<��a<9�a<7�a<_�a<w�a<��a<��a<��a<¬a<Ŭa<�a<�a<Ѭa<�a<߬a<�a<�a<�a<�a<٬a<�a<¬a<٬a<��a<��a<��a<��a<��a<_�a<n�a<5�a<*�a<��a<	�a<�a<��a<��a<\�a<\�a<%�a<��a<ުa<��a<��a<=�a<4�a<�a<éa<��a<J�a</�a<�a<ɨa<��a<,�a<��a<��a<��a<#�a<��a<��a<Z�a<�a<��a<�a<
�a<ߤa<h�a<2�a<��a<p�a<$�a<��a<X�a<�a<��a<<�a<֠a<j�a<��a<��a<!�a<՞a<P�a<�a<��a<�a<��a<!�a<ϛa<K�a<�a<|�a<�a<��a<"�a<��a<A�a<�a<r�a<��a<��a<�a<ҕa<F�a<��a<��a<$�a<̓a<P�a<�a<��a<Y�a<��a<��a<<�a<��a<��a<L�a<�a<��a<u�a<2�a<܎a<��a<^�a<E�a<�a<΍a<��a<g�a<R�a<�a<��a<ьa<Ča<��a<l�a<j�a<G�a<Y�a<,�a<+�a<*�a<�a<1�a<�a<9�a<!�a<M�a<I�a<_�a<|�a<��a<�  �  ��a<Ȍa<�a< �a<9�a<Z�a<��a<ȍa<��a<5�a<g�a<��a<�a<)�a<p�a<��a< �a<M�a<��a<��a<J�a<��a<��a<G�a<��a< �a<��a<ݓa<D�a<��a<�a<��a<��a<]�a<Ζa<P�a<��a<'�a<��a<�a<��a<�a<q�a<�a<v�a<ߛa<B�a<��a<7�a<��a<4�a<��a<�a<��a<��a<j�a<ܠa<M�a<��a<'�a<��a<
�a<h�a<ɣa</�a<��a<��a<c�a<��a<�a<d�a<��a<��a<d�a<��a<�a<E�a<��a<��a<�a<J�a<~�a<��a<��a<*�a<k�a<��a<Ūa<ܪa<�a<@�a<h�a<��a<��a<ͫa<�a<�a<(�a<A�a<^�a<d�a<��a<��a<��a<��a<��a<ìa<Ьa<�a<��a<�a<�a<�a<�a<�a<��a<ڬa<άa<۬a<��a<��a<��a<��a<|�a<n�a<[�a<;�a<>�a<�a<�a<īa<��a<��a<o�a<N�a<!�a<��a<תa<��a<�a<Q�a< �a<�a<��a<��a<Y�a<!�a<�a<��a<w�a<?�a<	�a<��a<s�a<3�a<�a<��a<^�a<
�a<��a<��a<�a<Τa<��a<�a<ȣa<x�a<�a<��a<l�a<��a<��a<,�a<Ơa<i�a<�a<��a<+�a<��a<T�a<�a<x�a<�a<��a<-�a<a<\�a<�a<n�a< �a<��a<+�a<Ƙa<P�a<֗a<q�a<��a<��a<8�a<ŕa<T�a<��a<��a<#�a<˓a<i�a<�a<��a<J�a<�a<��a<M�a<��a<��a<M�a<�a<��a<}�a<-�a<�a<��a<o�a<3�a<��a<͍a<��a<g�a<?�a<�a<��a<Ȍa<��a<��a<��a<{�a<N�a<G�a<;�a<&�a<&�a<2�a<�a<�a<:�a<.�a<?�a<]�a<e�a<t�a<��a<�  �  ��a<ӌa<،a<�a<A�a<n�a<��a<��a<
�a<"�a<p�a<��a<�a<3�a<`�a<ʏa<��a<g�a<��a<�a<\�a<��a<�a<]�a<Œa<�a<m�a<�a<>�a<Ŕa<�a<��a<ܕa<_�a<ۖa<3�a<a<	�a<��a< �a<��a<�a<n�a<�a<F�a<�a<T�a<ۜa<I�a<��a<2�a<��a</�a<��a<�a<j�a<ؠa<]�a<��a<G�a<��a<�a<r�a<ԣa<I�a<��a<	�a<9�a<��a<�a<c�a<ʦa<��a<i�a<��a<��a<1�a<��a<ʨa<�a<U�a<z�a<өa<�a<.�a<U�a<�a<Ѫa<�a<1�a<<�a<v�a<��a<��a<�a<�a< �a<�a<H�a<_�a<r�a<��a<��a<��a<��a<ڬa<٬a<߬a<�a<ͬa<�a<�a<��a<��a<�a<�a<ˬa<�a<��a<Ԭa<��a<��a<��a<��a<y�a<Q�a<F�a<�a<�a<��a<٫a<˫a<��a<~�a<;�a<*�a<�a<Ԫa<��a<n�a<d�a<�a<	�a<��a<��a<k�a<�a<�a<��a<��a<-�a<�a<��a<m�a<G�a<�a<��a<C�a<�a<˥a<c�a<.�a<��a<��a<�a<ߣa<w�a<�a<��a<=�a<�a<��a<F�a<נa<k�a<�a<��a<E�a<��a<`�a<�a<t�a<�a<��a<M�a<��a<W�a<�a<y�a<�a<��a<9�a<��a<G�a<ؗa<p�a<�a<��a<<�a<��a<g�a<�a<��a<-�a<��a<t�a<��a<��a<D�a<��a<��a<2�a<�a<��a<i�a<��a<ȏa<j�a<)�a<�a<��a<��a<%�a<�a<΍a<��a<w�a<0�a<$�a<�a<�a<��a<��a<��a<L�a<[�a<>�a<?�a<:�a<%�a<!�a<�a<9�a<�a<I�a<4�a<H�a<j�a<�a<��a<�  �  ��a<�a<��a<�a<<�a<b�a<��a<Ía<�a<9�a<f�a<��a<ێa<$�a<m�a<��a<��a<L�a<��a<��a<Y�a<��a<�a<W�a<��a<$�a<��a<��a<C�a<��a<�a<��a<��a<j�a<֖a<1�a<Ɨa<5�a<��a<�a<��a<�a<��a<��a<n�a<ߛa<N�a<��a<4�a<��a<,�a<��a<�a<��a<�a<q�a<�a<G�a<��a<'�a<��a<��a<v�a<ţa<&�a<��a<��a<a�a<��a<#�a<P�a<��a<��a<n�a<��a< �a<,�a<|�a<Ϩa<�a<N�a<~�a<��a<�a<J�a<k�a<��a<Ūa<�a<�a<=�a<w�a<��a<��a<Ϋa<�a<�a<'�a<@�a<M�a<n�a<��a<��a<��a<��a<��a<Ȭa<٬a<�a<�a<�a<��a<ܬa<�a<ެa<�a<�a<�a<��a<̬a<��a<��a<��a<}�a<`�a<^�a<[�a<.�a<�a<�a<̫a<��a<��a<y�a<S�a< �a<��a<Ȫa<��a<|�a<J�a<�a<�a<��a<��a<h�a<�a<ިa<��a<x�a<D�a<�a<קa<q�a<+�a<�a<��a<f�a<�a<ƥa<a�a<3�a<ۤa<��a<�a<ˣa<^�a<)�a<̢a<d�a<��a<��a<'�a<àa<q�a< �a<��a<'�a<��a<J�a<�a<�a<�a<��a<,�a<��a<Q�a<�a<i�a<��a<��a<,�a<Řa<X�a<��a<]�a<�a<��a<A�a<͕a<h�a<�a<��a<3�a<ϓa<m�a< �a<��a<E�a<�a<��a<Q�a<��a<��a<D�a<��a<ȏa<o�a<%�a<�a<��a<i�a<2�a<��a<��a<��a<f�a<I�a<�a<�a<ʌa<��a<��a<~�a<o�a<m�a<N�a<%�a<,�a<�a<0�a<0�a<7�a<�a<A�a<L�a<_�a<[�a<u�a<��a<�  �  ��a<�a<B�a<Q�a<��a<��a<�a<"�a<-�a<��a<Ǎa<�a<2�a<g�a<��a<��a<T�a<��a<�a<L�a<��a<�a<[�a<��a<�a<g�a<ؒa<*�a<��a<�a<q�a<֔a<_�a<��a<8�a<��a<�a<|�a<�a<s�a<�a<S�a<˙a<G�a<Κa<4�a<͛a<E�a<��a<'�a<��a</�a<~�a<��a<c�a<՟a<E�a<��a<3�a<��a<2�a<w�a<�a<^�a<��a<!�a<d�a<Ԥa<$�a<|�a<Υa<<�a<��a<֦a<%�a<^�a<ӧa<�a<3�a<��a<��a<��a<A�a<`�a<��a<�a<�a<:�a<v�a<��a<Ѫa<Ӫa<�a<N�a<;�a<m�a<}�a<��a<��a<ӫa<�a<�a<+�a<�a<>�a<K�a<U�a<c�a<M�a<h�a<Y�a<S�a<d�a<i�a<Y�a<n�a<F�a<J�a<b�a<;�a<�a<,�a<��a<��a<�a<��a<��a<��a<v�a<t�a<T�a<4�a<�a<ͪa<֪a<��a<g�a<I�a<�a<�a<��a<��a<W�a<T�a<�a<��a<��a<n�a<4�a<�a<��a<x�a<%�a<ڦa<��a<c�a<�a<�a<u�a<D�a<�a<��a<;�a<��a<��a<J�a<ۢa<�a<%�a<ԡa<a�a<�a<��a<T�a<��a<d�a<(�a<��a<1�a<��a<K�a<ۜa<n�a<�a<��a<P�a<��a<K�a<�a<|�a<�a<}�a<�a<��a<3�a<��a<j�a<��a<��a< �a<��a<h�a<��a<r�a<-�a<��a<X�a<�a<��a<;�a<�a<��a<@�a<��a<��a<h�a<��a<ʎa<��a<(�a<��a<��a<n�a<<�a<�a<ތa<��a<��a<O�a<K�a<(�a<�a<��a<��a<��a<��a<z�a<~�a<{�a<h�a<}�a<\�a<k�a<��a<��a<z�a<��a<��a<ŋa<ۋa<�  �  �a<+�a<7�a<e�a<��a<��a<֌a<�a<L�a<j�a<��a<�a<2�a<}�a<��a<�a<O�a<��a<ޏa<:�a<��a<�a<B�a<��a<�a<l�a<Ւa<H�a<��a<�a<a�a<�a<L�a<��a<,�a<��a<�a<z�a<�a<k�a<�a<k�a<�a<\�a<Śa<G�a<��a<"�a<��a<�a<��a<��a<t�a<�a<m�a<�a<V�a<Ġa<)�a<��a<��a<r�a<ߢa<:�a<��a<��a<w�a<Τa<6�a<��a<�a<5�a<z�a<�a<�a<s�a<��a<��a<A�a<��a<ͨa<�a<A�a<�a<��a<�a<�a<C�a<W�a<��a<��a<�a<�a<�a<@�a<e�a<��a<��a<��a<ҫa<�a<�a<��a<'�a<*�a<1�a<4�a<N�a<a�a<[�a<s�a<|�a<q�a<]�a<a�a<f�a<M�a<V�a<*�a<C�a<$�a<#�a<�a<�a<�a<�a<̫a<��a<��a<h�a<6�a<�a<�a<�a<��a<��a<k�a<I�a<'�a<��a<Ωa<��a<_�a<%�a<��a<ڨa<��a<V�a<�a<�a<��a<u�a<C�a<��a<��a<S�a<$�a<ҥa<��a<8�a<֤a<��a<9�a<��a<��a<C�a<�a<��a<:�a<ˡa<s�a<��a<��a<3�a<֟a<n�a<��a<��a<)�a<ĝa<\�a<�a<{�a<�a<��a<�a<��a<I�a<͙a<Y�a<�a<��a<�a<��a<T�a<ٖa<d�a<�a<��a<�a<��a<=�a<ޓa<��a<�a<ƒa<J�a<�a<��a<[�a<��a<��a<I�a<ߏa<��a<G�a<�a<��a<f�a<-�a<�a<a<��a<O�a<�a<یa<��a<v�a<h�a<6�a<�a<�a<ۋa<͋a<��a<��a<��a<��a<o�a<o�a<v�a<c�a<w�a<[�a<��a<��a<��a<��a<��a<�a<�  �  �a<�a<%�a<o�a<��a<��a<��a<��a<S�a<o�a<��a<��a<&�a<p�a<��a<��a<=�a<��a<�a<>�a<��a<ݐa<k�a<��a<�a<m�a<Òa<%�a<��a<	�a<^�a<�a<3�a<��a<=�a<��a<,�a<g�a<��a<l�a<�a<[�a<əa<G�a<��a<V�a<��a<N�a<��a<�a<��a<�a<��a<�a<i�a<ҟa<B�a<��a<"�a<��a<�a<~�a<ݢa<J�a<ˣa<�a<��a<��a<"�a<t�a<إa<3�a<y�a<ئa< �a<��a<��a<�a<J�a<j�a<Өa<�a<>�a<j�a<��a<ѩa<�a<H�a<e�a<��a<��a<�a<	�a<'�a<a�a<X�a<��a<��a<��a<ȫa<�a<
�a< �a</�a<�a<O�a<U�a<O�a<o�a<J�a<X�a<Z�a<d�a<_�a<j�a<Q�a<A�a<g�a<)�a<P�a<�a<�a<�a<�a<�a<īa<��a<��a<��a<g�a<Q�a<B�a<�a<�a<��a<��a<w�a<=�a<�a<�a<��a<��a<y�a<8�a<��a<ܨa<��a<�a<)�a<�a<��a<c�a< �a<�a<��a<P�a<.�a<��a<��a<I�a<ޤa<��a<&�a<�a<��a<D�a<�a<}�a<%�a<��a<��a<�a<àa<I�a<ҟa<}�a<��a<��a<&�a<��a<H�a<ٜa<v�a<��a<��a<!�a<a<G�a<ܙa<��a<�a<��a<	�a<��a<+�a<ɖa<b�a<�a<��a<��a<ʔa<I�a<�a<��a<�a<̒a<I�a<�a<��a<5�a<�a<��a<N�a<�a<��a<E�a<�a<a<x�a<N�a<�a<��a<s�a<A�a<
�a<�a<��a<y�a<p�a<+�a<-�a<�a<܋a<ۋa<��a<��a<��a<~�a<q�a<x�a<a�a<W�a<��a<Z�a<��a<x�a<��a<��a<��a<ߋa<�  �  �a<�a<T�a<Z�a<��a<��a<֌a<�a<8�a<�a<��a<ݍa<:�a<m�a<��a< �a<S�a<��a<�a<>�a<��a<��a<J�a<��a<��a<u�a<�a<:�a<��a<�a<t�a<ؔa<[�a<��a<�a<��a<�a<��a<��a<y�a<�a<]�a<ԙa<e�a<��a<9�a<��a<-�a<��a<!�a<��a<�a<t�a<�a<u�a<�a<V�a<ɠa<,�a<��a<�a<m�a<ܢa<E�a<��a<�a<j�a<�a<E�a<��a<ޥa<9�a<��a<֦a<2�a<a�a<��a<�a<:�a<��a<��a<�a<A�a<u�a<��a<��a<�a<3�a<c�a<��a<êa<تa< �a<.�a<0�a<j�a<��a<��a<��a<ܫa<ثa<��a<�a<�a<8�a<2�a<F�a<N�a<S�a<{�a<o�a<_�a<g�a<o�a<]�a<d�a<\�a<@�a<B�a<)�a</�a<(�a<�a<��a<�a<ɫa<��a<��a<�a<a�a<E�a<�a<�a<تa<Īa<��a<]�a<Q�a<�a<��a<éa<��a<N�a<:�a<��a<èa<��a<]�a<!�a<�a<��a<��a<5�a<�a<��a<f�a<�a<�a<��a<(�a<�a<��a<T�a<��a<��a<L�a<�a<��a<C�a<�a<f�a<�a<��a<8�a<ڟa<g�a<�a<��a<&�a<̝a<Z�a<�a<�a<�a<��a</�a<��a<F�a<יa<f�a<�a<��a</�a<ŗa<:�a<ϖa<g�a<��a<��a<-�a<��a<@�a<דa<y�a<-�a<��a<a�a<�a<��a<I�a<�a<��a<9�a<�a<��a<Z�a<��a<��a<~�a<�a<��a<��a<��a<C�a<�a<Ҍa<��a<��a<T�a<E�a<�a<��a<ۋa<��a<ˋa<��a<��a<��a<��a<k�a<s�a<r�a<a�a<s�a<o�a<��a<��a<��a<ɋa<�a<�  �  �a<�a<5�a<D�a<��a<��a<ʌa</�a<7�a<��a<��a<�a<G�a<]�a<̎a<�a<s�a<��a<��a<F�a<��a<
�a<7�a<a<�a<Y�a<Œa</�a<��a<��a<|�a<Ôa<R�a<��a<#�a<��a<��a<��a<ߗa<o�a<ܘa<c�a<�a<@�a<ǚa<0�a<ԛa<1�a<��a<3�a<��a<�a<p�a<�a<d�a<؟a<O�a<��a<N�a<��a<�a<i�a<�a<P�a<��a<+�a<g�a<Ȥa<�a<��a<�a< �a<��a<��a<7�a<\�a<ħa<��a<:�a<��a<��a<
�a<&�a<~�a<��a<Ωa<��a<:�a<��a<��a<Ѫa<�a<�a<6�a<;�a<��a<m�a<��a<��a<߫a<�a<�a<�a<�a<J�a<-�a<S�a<e�a<>�a<]�a<Z�a<u�a<_�a<d�a<R�a<R�a<e�a<7�a<]�a<&�a<6�a<�a<��a<��a<ګa<ޫa<��a<��a<i�a<v�a<W�a<�a<'�a<תa<Ūa<��a<r�a<^�a<�a<�a<��a<��a<Z�a<=�a<�a<ʨa<��a<J�a<>�a<�a<��a<e�a<*�a<��a<��a<n�a< �a<إa<��a<0�a<��a<��a<\�a<ԣa<��a<5�a<�a<��a<�a<͡a<]�a<%�a<��a<C�a<�a<^�a<�a<��a<E�a<��a<N�a<�a<h�a<&�a<��a<;�a<��a<X�a<�a<a�a<�a<��a<�a<��a<>�a<Ӗa<O�a<��a<g�a<2�a<��a<Z�a<�a<y�a<*�a<��a<f�a<�a<��a<A�a<��a<��a<@�a<�a<��a<g�a<�a<��a<��a<(�a<�a<��a<��a<5�a< �a<�a<��a<��a<O�a<W�a<
�a<�a<�a<��a<��a<��a<��a<y�a<v�a<`�a<b�a<{�a<X�a<��a<l�a<��a<��a<��a<ǋa<ыa<�  �  ��a<�a<:�a<t�a<��a<��a<�a< �a<K�a<{�a<��a<��a<-�a<l�a<Ɏa<�a<P�a<��a<�a<E�a<��a<�a<V�a<��a<�a<}�a<Ғa<.�a<��a<��a<p�a<�a<:�a<��a<'�a<��a<�a<~�a<��a<��a<ޘa<g�a<Ιa<M�a<Κa<V�a<��a</�a<��a<�a<��a<
�a<��a< �a<c�a<�a<X�a<��a<9�a<��a<�a<y�a<ݢa<?�a<��a<�a<~�a<פa<0�a<z�a<�a<)�a<��a<զa<�a<k�a<��a<��a<>�a<t�a<Ѩa<�a<.�a<w�a<��a<�a<�a<A�a<]�a<��a<��a<�a<�a<-�a<P�a<m�a<o�a<��a<��a<ͫa<�a<�a<�a<(�a<!�a<?�a<A�a<J�a<p�a<`�a<]�a<`�a<b�a<Y�a<x�a<V�a<N�a<L�a<9�a<5�a<"�a<�a<#�a<�a<ܫa<̫a<��a<��a<��a<b�a<B�a</�a<��a<�a<��a<��a<u�a<D�a<�a<�a<��a<��a<i�a<9�a<�a<Ҩa<��a<i�a<�a<�a<��a<r�a<(�a<�a<��a<b�a<0�a<��a<��a<3�a<�a<��a<=�a<�a<��a<8�a<�a<��a<+�a<ԡa<��a<��a<��a<=�a<ҟa<t�a<�a<��a<8�a<��a<Y�a<�a<k�a<�a<��a<,�a<��a<G�a<љa<k�a<�a<��a<"�a<��a<0�a<Ԗa<W�a<�a<��a<�a<��a<G�a<ޓa<}�a<�a<ʒa<a�a<�a<��a<=�a<�a<��a<G�a<�a<��a<E�a<�a<��a<}�a<=�a<��a<��a<��a<D�a<�a<�a<��a<��a<h�a<.�a<�a<�a<׋a<݋a<��a<��a<��a<|�a<k�a<��a<e�a<d�a<m�a<j�a<{�a<��a<��a<ŋa<��a<ԋa<�  �  �a<+�a<+�a<h�a<��a<��a<�a<�a<b�a<c�a<��a<�a<4�a<��a<��a<�a<G�a<��a<�a<5�a<��a<�a<j�a<��a<�a<l�a<Ғa<?�a<��a<�a<P�a<�a<8�a<��a<&�a<��a<�a<v�a<��a<a�a<ܘa<m�a<ƙa<l�a<��a<W�a<��a<@�a<��a<$�a<��a<��a<��a<�a<y�a<՟a<C�a<Ҡa<(�a<��a<��a<��a<�a<<�a<ãa<�a<��a<��a<C�a<u�a<�a<1�a<p�a<ۦa<�a<y�a<��a<�a<F�a<q�a<Ψa<�a<N�a<p�a<��a<�a<�a<R�a<T�a<��a<��a<��a<��a<"�a<P�a<`�a<��a<��a<��a<٫a<ݫa<�a<�a<;�a<(�a<L�a<H�a<U�a<h�a<L�a<|�a<T�a<~�a<O�a<_�a<W�a<I�a<[�a<*�a<@�a<"�a<�a<�a<ݫa<��a<��a<̫a<��a<��a<p�a<@�a<=�a<��a<�a<��a<��a<l�a<K�a<,�a<�a<کa<��a<j�a<6�a<��a<�a<��a<}�a<�a<��a<��a<s�a<9�a<�a<��a<B�a<%�a<��a<��a<2�a<Фa<��a<5�a<�a<��a<5�a<��a<z�a<I�a<��a<��a<�a<��a<=�a<ݟa<��a<�a<��a<%�a<Нa<K�a<ٜa<��a< �a<��a<�a<Śa<S�a<ϙa<��a<�a<��a<�a<×a<+�a<Ֆa<`�a<ߕa<��a<�a<��a<6�a<דa<��a<
�a<ǒa<?�a<�a<��a<E�a<��a<��a<X�a<ۏa<��a<E�a<�a<��a<s�a<=�a<�a<΍a<m�a<M�a<�a<׌a<Ìa<m�a<|�a<4�a<)�a<��a<�a<ԋa<��a<��a<|�a<��a<`�a<m�a<f�a<_�a<|�a<[�a<��a<��a<��a<��a<��a<��a<�  �  �a<�a<1�a<Y�a<��a<��a<یa<�a<?�a<y�a<ҍa<�a<1�a<y�a<��a<
�a<O�a<��a<�a<<�a<��a<�a<H�a<��a<#�a<c�a<ɒa<5�a<��a<	�a<j�a<ڔa<L�a<��a<$�a<��a<��a<��a<��a<p�a<�a<`�a<șa<V�a<��a<G�a<ɛa<:�a<��a<)�a<��a<�a<��a<�a<p�a<ޟa<Q�a<Ša<)�a<��a< �a<r�a<�a<>�a<��a<�a<{�a<��a<-�a<x�a<٥a</�a<��a<Ҧa<$�a<W�a<��a<��a<3�a<��a<��a<��a<;�a<e�a<��a<֩a<�a<T�a<o�a<��a<��a<�a<�a<G�a<L�a<h�a<��a<��a<��a<իa<ޫa<�a<�a<�a<1�a<8�a<K�a<d�a<X�a<W�a<i�a<P�a<g�a<`�a<_�a<W�a<N�a<7�a<K�a<%�a<�a<�a<	�a<�a<�a<��a<��a<��a<~�a<{�a<K�a<%�a<	�a<ߪa<��a<��a<j�a<I�a<#�a<�a<̩a<��a<i�a<S�a<��a<Өa<��a<\�a<*�a<�a<��a<j�a</�a<ݦa<��a<\�a<�a<ҥa<{�a<0�a<�a<{�a<D�a<�a<��a<=�a<�a<|�a<3�a<��a<t�a<�a<��a<8�a<�a<j�a<�a<��a<(�a<ǝa<T�a<�a<|�a<�a<��a<>�a<��a<S�a<љa<r�a<�a<��a<	�a<��a</�a<ʖa<]�a<�a<��a<�a<��a<O�a<�a<r�a<�a<��a<S�a<��a<��a<B�a<�a<��a<Z�a<��a<��a<M�a<�a<��a<��a<9�a<��a<��a<�a<K�a<�a<،a<ьa<��a<X�a<>�a<�a<��a<�a<ŋa<��a<��a<w�a<��a<q�a<m�a<f�a<d�a<X�a<|�a<k�a<�a<��a<��a<��a<ދa<�  �  �a<��a<H�a<j�a<o�a<��a<܌a<#�a<>�a<��a<��a<��a<B�a<l�a<َa<�a<h�a<��a<�a<C�a<��a<�a<E�a<��a<�a<��a<גa<'�a<��a<�a<z�a<ʔa<P�a<��a<�a<��a<�a<��a<�a<|�a<ߘa<c�a<�a<>�a<�a<;�a<��a<$�a<��a<.�a<��a<�a<h�a<�a<i�a<�a<c�a<��a<L�a<��a<�a<h�a<�a<J�a<��a<�a<i�a<�a<�a<��a<�a<"�a<��a<��a<=�a<R�a<��a<�a<7�a<��a<��a<�a<#�a<��a<��a<ݩa<&�a<(�a<i�a<��a<˪a<�a<�a<)�a<8�a<��a<t�a<��a<��a<ܫa<�a<�a<�a<�a<@�a<:�a<A�a<>�a<^�a<r�a<I�a<}�a<[�a<c�a<`�a<J�a<o�a<0�a<N�a<�a<=�a<�a<�a<��a<֫a<�a<��a<��a<��a<P�a<F�a<&�a<�a<ުa<̪a<��a<x�a<Y�a<�a<�a<��a<��a<^�a<.�a<�a<Ψa<��a<X�a<&�a<ѧa<ħa<w�a<"�a<�a<��a<l�a<�a<֥a<��a<!�a<�a<y�a<c�a<ۣa<��a<8�a<�a<��a<�a<�a<h�a< �a<��a<>�a<�a<`�a<�a<��a<E�a<��a<`�a<��a<q�a<$�a<�a<5�a<��a<T�a<ܙa<]�a<�a<��a<4�a<��a<D�a<֖a<P�a<��a<q�a<8�a<��a<F�a<Փa<v�a<)�a<��a<d�a<�a<��a<A�a<�a<��a<.�a<��a<��a<b�a<�a<��a<z�a<%�a<�a<��a<��a<C�a<�a<�a<��a<��a<X�a<L�a<�a<�a<ʋa<ʋa<Ëa<��a<��a<u�a<t�a<n�a<Y�a<��a<Q�a<�a<^�a<��a<��a<��a<a<͋a<�  �  ��a<�a<3�a<U�a<��a<όa<�a<�a<P�a<��a<��a<�a<;�a<l�a<��a<��a<^�a<��a<�a<U�a<��a<�a<]�a<Ǒa<�a<h�a<̒a<)�a<��a<��a<t�a<Քa<6�a<��a<#�a<��a<�a<~�a<ۗa<p�a<ژa<S�a<ٙa<L�a<��a<9�a<˛a<S�a<��a<'�a<��a<�a<��a<�a<i�a<ٟa<K�a<��a<G�a<��a<�a<��a<�a<K�a<ʣa<$�a<l�a<Ťa<&�a<��a<ҥa<#�a<��a<��a<�a<m�a<��a<��a<D�a<q�a<��a<�a<,�a<r�a<��a<שa<�a<5�a<��a<��a<��a<�a<�a<4�a<T�a<}�a<��a<��a<��a<ګa<��a<��a<�a<,�a</�a<E�a<k�a<W�a<M�a<X�a<[�a<l�a<V�a<\�a<a�a<=�a<S�a<C�a<@�a<)�a<*�a<��a<
�a<��a<ԫa<իa<��a<��a<z�a<f�a<f�a<2�a<�a<�a<ʪa<��a<��a<R�a<�a<��a<��a<��a<s�a<:�a<�a<Ҩa<��a<q�a<D�a<�a<��a<m�a<#�a<�a<��a<f�a<�a<��a<��a</�a<�a<��a<=�a<Уa<��a<3�a<ڢa<��a<)�a<ǡa<e�a<�a<Ƞa<F�a<��a<|�a<�a<��a<F�a<��a<O�a<�a<s�a<�a<��a<6�a<Śa<Q�a<ݙa<��a<�a<��a<�a<��a<8�a<Öa<Q�a<�a<k�a<�a<��a<J�a<�a<��a<�a<��a<^�a<�a<��a<:�a<�a<��a<;�a<�a<��a<S�a<
�a<юa<��a<B�a<�a<��a<��a<?�a<�a<��a<��a<��a<l�a<<�a<"�a<�a<�a<��a<��a<��a<��a<p�a<n�a<o�a<M�a<i�a<d�a<r�a<o�a<��a<}�a<��a<��a<ˋa<�  �  ߋa<0�a<?�a<]�a<��a<��a<֌a<	�a<L�a<r�a<̍a<�a<*�a<��a<��a<%�a<?�a<��a<��a<E�a<��a<�a<E�a<��a< �a<f�a<ߒa<C�a<��a<�a<[�a<�a<D�a<��a<�a<��a<�a<n�a<�a<g�a<�a<d�a<˙a<m�a<��a<O�a<��a<(�a<��a<�a<��a<�a<��a<�a<�a<�a<X�a<۠a<�a<��a<�a<}�a<ޢa<:�a<��a<�a<��a<Ĥa<I�a<��a<٥a<4�a<w�a<�a<�a<e�a<��a<�a<6�a<v�a<ͨa<�a<D�a<e�a<��a<��a<�a<R�a<W�a<��a<��a<�a<�a<-�a<M�a<S�a<��a<��a<ӫa<ԫa<׫a<�a<�a<'�a<)�a<1�a<;�a<W�a<]�a<b�a<~�a<K�a<q�a<X�a<^�a<e�a<<�a<@�a</�a<,�a<�a<�a<�a<�a<�a<��a<ѫa<��a<��a<u�a<8�a<�a< �a<�a<��a<��a<e�a<A�a<<�a<�a<�a<��a<f�a<A�a<�a<Ψa<��a<X�a<�a<�a<��a<��a<>�a<ۦa<��a<M�a<#�a<ɥa<v�a<*�a<֤a<��a<-�a<�a<��a<@�a<�a<~�a<K�a<ȡa<{�a<�a<��a<2�a<՟a<y�a<��a<��a<�a<֝a<c�a<�a<��a<�a<��a<#�a<��a<H�a<̙a<a�a<�a<��a<�a<ȗa<8�a<ʖa<b�a<�a<��a<�a<��a<7�a<ԓa<u�a<�a<ƒa<I�a<�a<��a<O�a<�a<��a<X�a<ޏa<��a<I�a<�a<Ǝa<~�a<:�a<�a<ݍa<w�a<a�a<�a<ьa<͌a<|�a<h�a<5�a<�a<�a<�a<ɋa<��a<��a<r�a<��a<i�a<l�a<t�a<R�a<a�a<`�a<r�a<u�a<��a<��a<��a<�a<�  �  �a<�a<%�a<_�a<��a<��a<��a<&�a<S�a<t�a<��a<��a<3�a<��a<��a<�a<K�a<��a<�a<C�a<��a<�a<^�a<��a<�a<d�a<��a<&�a<��a<�a<X�a<Ĕa<=�a<��a<,�a<��a<�a<z�a<�a<W�a<ޘa<c�a<șa<A�a<��a<I�a<��a<<�a<a<1�a<��a<�a<��a<��a<t�a<ܟa<J�a<͠a<4�a<��a<�a<��a<�a<b�a<��a<�a<x�a<��a<�a<v�a<ڥa<'�a<k�a<��a<�a<k�a<��a<��a<:�a<v�a<��a<�a<6�a<k�a<��a<˩a<��a<C�a<g�a<��a<تa<�a<�a<+�a<\�a<c�a<��a<��a<ūa<ԫa<�a<�a<�a<-�a<D�a<S�a<N�a<T�a<]�a<K�a<U�a<Z�a<n�a<U�a<K�a<O�a<O�a<P�a<B�a<9�a<#�a<�a<��a<�a<�a<ƫa<��a<��a<��a<m�a<K�a<@�a<�a<��a<��a<��a<}�a<J�a<2�a<�a<թa<��a<y�a<:�a<�a<ݨa<��a<q�a<$�a<�a<��a<\�a<!�a<�a<��a<J�a<�a<åa<}�a<8�a<�a<��a<9�a<�a<��a<7�a<�a<|�a<�a<��a<u�a<�a<��a<Y�a<�a<|�a<��a<��a<4�a<˝a<R�a<��a<��a<�a<��a<%�a<Úa<Y�a<��a<u�a<��a<��a<�a<��a<,�a<˖a<V�a<ڕa<u�a<�a<��a<J�a<�a<y�a<�a<��a<D�a<��a<��a<7�a<ܐa<��a<I�a<�a<��a<o�a<�a<Ďa<{�a<I�a<�a<ɍa<q�a<S�a<�a<�a<Ìa<~�a<m�a<Q�a<0�a<�a<�a<ʋa<��a<��a<��a<��a<g�a<Y�a<^�a<e�a<q�a<s�a<�a<��a<��a<��a<��a<��a<�  �  �a<�a<B�a<i�a<y�a<��a<ڌa<��a<I�a<��a<��a<�a<'�a<��a<�a<�a<E�a<��a<��a<O�a<��a<�a<D�a<��a<��a<�a<ݒa<B�a<��a<�a<��a<ߔa<D�a<��a<�a<��a<�a<��a<�a<��a<�a<P�a<�a<]�a<Ԛa<;�a<��a<3�a<��a<�a<��a<�a<��a<
�a<d�a<��a<q�a<��a<?�a<��a<�a<��a<֢a<A�a<��a<�a<e�a<ޤa<:�a<��a<֥a<0�a<��a<æa<�a<^�a<��a<�a<3�a<~�a<��a<�a<&�a<y�a<��a<�a<!�a<2�a<t�a<��a<��a<ܪa<�a<0�a<[�a<a�a<��a<ƫa<̫a<ȫa<�a<��a<�a<(�a<�a<4�a<Q�a<I�a<b�a<i�a<k�a<w�a<I�a<k�a<v�a<F�a<S�a<;�a<*�a<#�a<%�a<�a<�a<�a<ƫa<ޫa<��a<��a<��a<Z�a<R�a<#�a<�a<�a<ƪa<��a<��a<?�a<,�a<�a<ǩa<��a<�a<7�a<�a<Шa<��a<X�a<3�a<�a<§a<}�a<<�a<��a<��a<y�a<�a<ʥa<}�a<%�a<Фa<��a<B�a<ݣa<��a<E�a<آa<��a<:�a<ۡa<g�a<�a<��a<9�a<̟a<|�a<	�a<��a<A�a<��a<q�a<�a<p�a<�a<��a<.�a<Ța<@�a<ԙa<e�a<��a<�a<)�a<��a<Q�a<ǖa<_�a<�a<v�a<�a<��a<7�a<ԓa<s�a<�a<��a<t�a<�a<��a<V�a<��a<��a<8�a<��a<��a<I�a<�a<͎a<��a<H�a<�a<��a<��a<Y�a<	�a<��a<��a<��a<h�a<*�a<�a<�a<֋a<΋a<��a<��a<��a<c�a<}�a<��a<V�a<i�a<\�a<[�a<i�a<��a<��a<��a<ыa<��a<�  �  �a<�a<%�a<_�a<��a<��a<��a<&�a<S�a<t�a<��a<��a<3�a<��a<��a<�a<K�a<��a<�a<C�a<��a<�a<^�a<��a<�a<d�a<��a<&�a<��a<�a<X�a<Ĕa<=�a<��a<,�a<��a<�a<z�a<�a<W�a<ޘa<c�a<șa<A�a<��a<I�a<��a<<�a<a<1�a<��a<�a<��a<��a<t�a<ܟa<J�a<͠a<4�a<��a<�a<��a<�a<b�a<��a<�a<x�a<��a<�a<v�a<ڥa<'�a<k�a<��a<�a<k�a<��a<��a<:�a<v�a<��a<�a<6�a<k�a<��a<˩a<��a<C�a<g�a<��a<تa<�a<�a<+�a<\�a<c�a<��a<��a<ūa<ԫa<�a<�a<�a<-�a<D�a<S�a<N�a<T�a<]�a<K�a<U�a<Z�a<n�a<U�a<K�a<O�a<O�a<P�a<B�a<9�a<#�a<�a<��a<�a<�a<ƫa<��a<��a<��a<m�a<K�a<@�a<�a<��a<��a<��a<}�a<J�a<2�a<�a<թa<��a<y�a<:�a<�a<ݨa<��a<q�a<$�a<�a<��a<\�a<!�a<�a<��a<J�a<�a<åa<}�a<8�a<�a<��a<9�a<�a<��a<7�a<�a<|�a<�a<��a<u�a<�a<��a<Y�a<�a<|�a<��a<��a<4�a<˝a<R�a<��a<��a<�a<��a<%�a<Úa<Y�a<��a<u�a<��a<��a<�a<��a<,�a<˖a<V�a<ڕa<u�a<�a<��a<J�a<�a<y�a<�a<��a<D�a<��a<��a<7�a<ܐa<��a<I�a<�a<��a<o�a<�a<Ďa<{�a<I�a<�a<ɍa<q�a<S�a<�a<�a<Ìa<~�a<m�a<Q�a<0�a<�a<�a<ʋa<��a<��a<��a<��a<g�a<Y�a<^�a<e�a<q�a<s�a<�a<��a<��a<��a<��a<��a<�  �  ߋa<0�a<?�a<]�a<��a<��a<֌a<	�a<L�a<r�a<̍a<�a<*�a<��a<��a<%�a<?�a<��a<��a<E�a<��a<�a<E�a<��a< �a<f�a<ߒa<C�a<��a<�a<[�a<�a<D�a<��a<�a<��a<�a<n�a<�a<g�a<�a<d�a<˙a<m�a<��a<O�a<��a<(�a<��a<�a<��a<�a<��a<�a<�a<�a<X�a<۠a<�a<��a<�a<}�a<ޢa<:�a<��a<�a<��a<Ĥa<I�a<��a<٥a<4�a<w�a<�a<�a<e�a<��a<�a<6�a<v�a<ͨa<�a<D�a<e�a<��a<��a<�a<R�a<W�a<��a<��a<�a<�a<-�a<M�a<S�a<��a<��a<ӫa<ԫa<׫a<�a<�a<'�a<)�a<1�a<;�a<W�a<]�a<b�a<~�a<K�a<q�a<X�a<^�a<e�a<<�a<@�a</�a<,�a<�a<�a<�a<�a<�a<��a<ѫa<��a<��a<u�a<8�a<�a< �a<�a<��a<��a<e�a<A�a<<�a<�a<�a<��a<f�a<A�a<�a<Ψa<��a<X�a<�a<�a<��a<��a<>�a<ۦa<��a<M�a<#�a<ɥa<v�a<*�a<֤a<��a<-�a<�a<��a<@�a<�a<~�a<K�a<ȡa<{�a<�a<��a<2�a<՟a<y�a<��a<��a<�a<֝a<c�a<�a<��a<�a<��a<#�a<��a<H�a<̙a<a�a<�a<��a<�a<ȗa<8�a<ʖa<b�a<�a<��a<�a<��a<7�a<ԓa<u�a<�a<ƒa<I�a<�a<��a<O�a<�a<��a<X�a<ޏa<��a<I�a<�a<Ǝa<~�a<:�a<�a<ݍa<w�a<a�a<�a<ьa<͌a<|�a<h�a<5�a<�a<�a<�a<ɋa<��a<��a<r�a<��a<i�a<l�a<t�a<R�a<a�a<`�a<r�a<u�a<��a<��a<��a<�a<�  �  ��a<�a<3�a<U�a<��a<όa<�a<�a<P�a<��a<��a<�a<;�a<l�a<��a<��a<^�a<��a<�a<U�a<��a<�a<]�a<Ǒa<�a<h�a<̒a<)�a<��a<��a<t�a<Քa<6�a<��a<#�a<��a<�a<~�a<ۗa<p�a<ژa<S�a<ٙa<L�a<��a<9�a<˛a<S�a<��a<'�a<��a<�a<��a<�a<i�a<ٟa<K�a<��a<G�a<��a<�a<��a<�a<K�a<ʣa<$�a<l�a<Ťa<&�a<��a<ҥa<#�a<��a<��a<�a<m�a<��a<��a<D�a<q�a<��a<�a<,�a<r�a<��a<שa<�a<5�a<��a<��a<��a<�a<�a<4�a<T�a<}�a<��a<��a<��a<ګa<��a<��a<�a<,�a</�a<E�a<k�a<W�a<M�a<X�a<[�a<l�a<V�a<\�a<a�a<=�a<S�a<C�a<@�a<)�a<*�a<��a<
�a<��a<ԫa<իa<��a<��a<z�a<f�a<f�a<2�a<�a<�a<ʪa<��a<��a<R�a<�a<��a<��a<��a<s�a<:�a<�a<Ҩa<��a<q�a<D�a<�a<��a<m�a<#�a<�a<��a<f�a<�a<��a<��a</�a<�a<��a<=�a<Уa<��a<3�a<ڢa<��a<)�a<ǡa<e�a<�a<Ƞa<F�a<��a<|�a<�a<��a<F�a<��a<O�a<�a<s�a<�a<��a<6�a<Śa<Q�a<ݙa<��a<�a<��a<�a<��a<8�a<Öa<Q�a<�a<k�a<�a<��a<J�a<�a<��a<�a<��a<^�a<�a<��a<:�a<�a<��a<;�a<�a<��a<S�a<
�a<юa<��a<B�a<�a<��a<��a<?�a<�a<��a<��a<��a<l�a<<�a<"�a<�a<�a<��a<��a<��a<��a<p�a<n�a<o�a<M�a<i�a<d�a<r�a<o�a<��a<}�a<��a<��a<ˋa<�  �  �a<��a<H�a<j�a<o�a<��a<܌a<#�a<>�a<��a<��a<��a<B�a<l�a<َa<�a<h�a<��a<�a<C�a<��a<�a<E�a<��a<�a<��a<גa<'�a<��a<�a<z�a<ʔa<P�a<��a<�a<��a<�a<��a<�a<|�a<ߘa<c�a<�a<>�a<�a<;�a<��a<$�a<��a<.�a<��a<�a<h�a<�a<i�a<�a<c�a<��a<L�a<��a<�a<h�a<�a<J�a<��a<�a<i�a<�a<�a<��a<�a<"�a<��a<��a<=�a<R�a<��a<�a<7�a<��a<��a<�a<#�a<��a<��a<ݩa<&�a<(�a<i�a<��a<˪a<�a<�a<)�a<8�a<��a<t�a<��a<��a<ܫa<�a<�a<�a<�a<@�a<:�a<A�a<>�a<^�a<r�a<I�a<}�a<[�a<c�a<`�a<J�a<o�a<0�a<N�a<�a<=�a<�a<�a<��a<֫a<�a<��a<��a<��a<P�a<F�a<&�a<�a<ުa<̪a<��a<x�a<Y�a<�a<�a<��a<��a<^�a<.�a<�a<Ψa<��a<X�a<&�a<ѧa<ħa<w�a<"�a<�a<��a<l�a<�a<֥a<��a<!�a<�a<y�a<c�a<ۣa<��a<8�a<�a<��a<�a<�a<h�a< �a<��a<>�a<�a<`�a<�a<��a<E�a<��a<`�a<��a<q�a<$�a<�a<5�a<��a<T�a<ܙa<]�a<�a<��a<4�a<��a<D�a<֖a<P�a<��a<q�a<8�a<��a<F�a<Փa<v�a<)�a<��a<d�a<�a<��a<A�a<�a<��a<.�a<��a<��a<b�a<�a<��a<z�a<%�a<�a<��a<��a<C�a<�a<�a<��a<��a<X�a<L�a<�a<�a<ʋa<ʋa<Ëa<��a<��a<u�a<t�a<n�a<Y�a<��a<Q�a<�a<^�a<��a<��a<��a<a<͋a<�  �  �a<�a<1�a<Y�a<��a<��a<یa<�a<?�a<y�a<ҍa<�a<1�a<y�a<��a<
�a<O�a<��a<�a<<�a<��a<�a<H�a<��a<#�a<c�a<ɒa<5�a<��a<	�a<j�a<ڔa<L�a<��a<$�a<��a<��a<��a<��a<p�a<�a<`�a<șa<V�a<��a<G�a<ɛa<:�a<��a<)�a<��a<�a<��a<�a<p�a<ޟa<Q�a<Ša<)�a<��a< �a<r�a<�a<>�a<��a<�a<{�a<��a<-�a<x�a<٥a</�a<��a<Ҧa<$�a<W�a<��a<��a<3�a<��a<��a<��a<;�a<e�a<��a<֩a<�a<T�a<o�a<��a<��a<�a<�a<G�a<L�a<h�a<��a<��a<��a<իa<ޫa<�a<�a<�a<1�a<8�a<K�a<d�a<X�a<W�a<i�a<P�a<g�a<`�a<_�a<W�a<N�a<7�a<K�a<%�a<�a<�a<	�a<�a<�a<��a<��a<��a<~�a<{�a<K�a<%�a<	�a<ߪa<��a<��a<j�a<I�a<#�a<�a<̩a<��a<i�a<S�a<��a<Өa<��a<\�a<*�a<�a<��a<j�a</�a<ݦa<��a<\�a<�a<ҥa<{�a<0�a<�a<{�a<D�a<�a<��a<=�a<�a<|�a<3�a<��a<t�a<�a<��a<8�a<�a<j�a<�a<��a<(�a<ǝa<T�a<�a<|�a<�a<��a<>�a<��a<S�a<љa<r�a<�a<��a<	�a<��a</�a<ʖa<]�a<�a<��a<�a<��a<O�a<�a<r�a<�a<��a<S�a<��a<��a<B�a<�a<��a<Z�a<��a<��a<M�a<�a<��a<��a<9�a<��a<��a<�a<K�a<�a<،a<ьa<��a<X�a<>�a<�a<��a<�a<ŋa<��a<��a<w�a<��a<q�a<m�a<f�a<d�a<X�a<|�a<k�a<�a<��a<��a<��a<ދa<�  �  �a<+�a<+�a<h�a<��a<��a<�a<�a<b�a<c�a<��a<�a<4�a<��a<��a<�a<G�a<��a<�a<5�a<��a<�a<j�a<��a<�a<l�a<Ғa<?�a<��a<�a<P�a<�a<8�a<��a<&�a<��a<�a<v�a<��a<a�a<ܘa<m�a<ƙa<l�a<��a<W�a<��a<@�a<��a<$�a<��a<��a<��a<�a<y�a<՟a<C�a<Ҡa<(�a<��a<��a<��a<�a<<�a<ãa<�a<��a<��a<C�a<u�a<�a<1�a<p�a<ۦa<�a<y�a<��a<�a<F�a<q�a<Ψa<�a<N�a<p�a<��a<�a<�a<R�a<T�a<��a<��a<��a<��a<"�a<P�a<`�a<��a<��a<��a<٫a<ݫa<�a<�a<;�a<(�a<L�a<H�a<U�a<h�a<L�a<|�a<T�a<~�a<O�a<_�a<W�a<I�a<[�a<*�a<@�a<"�a<�a<�a<ݫa<��a<��a<̫a<��a<��a<p�a<@�a<=�a<��a<�a<��a<��a<l�a<K�a<,�a<�a<کa<��a<j�a<6�a<��a<�a<��a<}�a<�a<��a<��a<s�a<9�a<�a<��a<B�a<%�a<��a<��a<2�a<Фa<��a<5�a<�a<��a<5�a<��a<z�a<I�a<��a<��a<�a<��a<=�a<ݟa<��a<�a<��a<%�a<Нa<K�a<ٜa<��a< �a<��a<�a<Śa<S�a<ϙa<��a<�a<��a<�a<×a<+�a<Ֆa<`�a<ߕa<��a<�a<��a<6�a<דa<��a<
�a<ǒa<?�a<�a<��a<E�a<��a<��a<X�a<ۏa<��a<E�a<�a<��a<s�a<=�a<�a<΍a<m�a<M�a<�a<׌a<Ìa<m�a<|�a<4�a<)�a<��a<�a<ԋa<��a<��a<|�a<��a<`�a<m�a<f�a<_�a<|�a<[�a<��a<��a<��a<��a<��a<��a<�  �  ��a<�a<:�a<t�a<��a<��a<�a< �a<K�a<{�a<��a<��a<-�a<l�a<Ɏa<�a<P�a<��a<�a<E�a<��a<�a<V�a<��a<�a<}�a<Ғa<.�a<��a<��a<p�a<�a<:�a<��a<'�a<��a<�a<~�a<��a<��a<ޘa<g�a<Ιa<M�a<Κa<V�a<��a</�a<��a<�a<��a<
�a<��a< �a<c�a<�a<X�a<��a<9�a<��a<�a<y�a<ݢa<?�a<��a<�a<~�a<פa<0�a<z�a<�a<)�a<��a<զa<�a<k�a<��a<��a<>�a<t�a<Ѩa<�a<.�a<w�a<��a<�a<�a<A�a<]�a<��a<��a<�a<�a<-�a<P�a<m�a<o�a<��a<��a<ͫa<�a<�a<�a<(�a<!�a<?�a<A�a<J�a<p�a<`�a<]�a<`�a<b�a<Y�a<x�a<V�a<N�a<L�a<9�a<5�a<"�a<�a<#�a<�a<ܫa<̫a<��a<��a<��a<b�a<B�a</�a<��a<�a<��a<��a<u�a<D�a<�a<�a<��a<��a<i�a<9�a<�a<Ҩa<��a<i�a<�a<�a<��a<r�a<(�a<�a<��a<b�a<0�a<��a<��a<3�a<�a<��a<=�a<�a<��a<8�a<�a<��a<+�a<ԡa<��a<��a<��a<=�a<ҟa<t�a<�a<��a<8�a<��a<Y�a<�a<k�a<�a<��a<,�a<��a<G�a<љa<k�a<�a<��a<"�a<��a<0�a<Ԗa<W�a<�a<��a<�a<��a<G�a<ޓa<}�a<�a<ʒa<a�a<�a<��a<=�a<�a<��a<G�a<�a<��a<E�a<�a<��a<}�a<=�a<��a<��a<��a<D�a<�a<�a<��a<��a<h�a<.�a<�a<�a<׋a<݋a<��a<��a<��a<|�a<k�a<��a<e�a<d�a<m�a<j�a<{�a<��a<��a<ŋa<��a<ԋa<�  �  �a<�a<5�a<D�a<��a<��a<ʌa</�a<7�a<��a<��a<�a<G�a<]�a<̎a<�a<s�a<��a<��a<F�a<��a<
�a<7�a<a<�a<Y�a<Œa</�a<��a<��a<|�a<Ôa<R�a<��a<#�a<��a<��a<��a<ߗa<o�a<ܘa<c�a<�a<@�a<ǚa<0�a<ԛa<1�a<��a<3�a<��a<�a<p�a<�a<d�a<؟a<O�a<��a<N�a<��a<�a<i�a<�a<P�a<��a<+�a<g�a<Ȥa<�a<��a<�a< �a<��a<��a<7�a<\�a<ħa<��a<:�a<��a<��a<
�a<&�a<~�a<��a<Ωa<��a<:�a<��a<��a<Ѫa<�a<�a<6�a<;�a<��a<m�a<��a<��a<߫a<�a<�a<�a<�a<J�a<-�a<S�a<e�a<>�a<]�a<Z�a<u�a<_�a<d�a<R�a<R�a<e�a<7�a<]�a<&�a<6�a<�a<��a<��a<ګa<ޫa<��a<��a<i�a<v�a<W�a<�a<'�a<תa<Ūa<��a<r�a<^�a<�a<�a<��a<��a<Z�a<=�a<�a<ʨa<��a<J�a<>�a<�a<��a<e�a<*�a<��a<��a<n�a< �a<إa<��a<0�a<��a<��a<\�a<ԣa<��a<5�a<�a<��a<�a<͡a<]�a<%�a<��a<C�a<�a<^�a<�a<��a<E�a<��a<N�a<�a<h�a<&�a<��a<;�a<��a<X�a<�a<a�a<�a<��a<�a<��a<>�a<Ӗa<O�a<��a<g�a<2�a<��a<Z�a<�a<y�a<*�a<��a<f�a<�a<��a<A�a<��a<��a<@�a<�a<��a<g�a<�a<��a<��a<(�a<�a<��a<��a<5�a< �a<�a<��a<��a<O�a<W�a<
�a<�a<�a<��a<��a<��a<��a<y�a<v�a<`�a<b�a<{�a<X�a<��a<l�a<��a<��a<��a<ǋa<ыa<�  �  �a<�a<T�a<Z�a<��a<��a<֌a<�a<8�a<�a<��a<ݍa<:�a<m�a<��a< �a<S�a<��a<�a<>�a<��a<��a<J�a<��a<��a<u�a<�a<:�a<��a<�a<t�a<ؔa<[�a<��a<�a<��a<�a<��a<��a<y�a<�a<]�a<ԙa<e�a<��a<9�a<��a<-�a<��a<!�a<��a<�a<t�a<�a<u�a<�a<V�a<ɠa<,�a<��a<�a<m�a<ܢa<E�a<��a<�a<j�a<�a<E�a<��a<ޥa<9�a<��a<֦a<2�a<a�a<��a<�a<:�a<��a<��a<�a<A�a<u�a<��a<��a<�a<3�a<c�a<��a<êa<تa< �a<.�a<0�a<j�a<��a<��a<��a<ܫa<ثa<��a<�a<�a<8�a<2�a<F�a<N�a<S�a<{�a<o�a<_�a<g�a<o�a<]�a<d�a<\�a<@�a<B�a<)�a</�a<(�a<�a<��a<�a<ɫa<��a<��a<�a<a�a<E�a<�a<�a<تa<Īa<��a<]�a<Q�a<�a<��a<éa<��a<N�a<:�a<��a<èa<��a<]�a<!�a<�a<��a<��a<5�a<�a<��a<f�a<�a<�a<��a<(�a<�a<��a<T�a<��a<��a<L�a<�a<��a<C�a<�a<f�a<�a<��a<8�a<ڟa<g�a<�a<��a<&�a<̝a<Z�a<�a<�a<�a<��a</�a<��a<F�a<יa<f�a<�a<��a</�a<ŗa<:�a<ϖa<g�a<��a<��a<-�a<��a<@�a<דa<y�a<-�a<��a<a�a<�a<��a<I�a<�a<��a<9�a<�a<��a<Z�a<��a<��a<~�a<�a<��a<��a<��a<C�a<�a<Ҍa<��a<��a<T�a<E�a<�a<��a<ۋa<��a<ˋa<��a<��a<��a<��a<k�a<s�a<r�a<a�a<s�a<o�a<��a<��a<��a<ɋa<�a<�  �  �a<�a<%�a<o�a<��a<��a<��a<��a<S�a<o�a<��a<��a<&�a<p�a<��a<��a<=�a<��a<�a<>�a<��a<ݐa<k�a<��a<�a<m�a<Òa<%�a<��a<	�a<^�a<�a<3�a<��a<=�a<��a<,�a<g�a<��a<l�a<�a<[�a<əa<G�a<��a<V�a<��a<N�a<��a<�a<��a<�a<��a<�a<i�a<ҟa<B�a<��a<"�a<��a<�a<~�a<ݢa<J�a<ˣa<�a<��a<��a<"�a<t�a<إa<3�a<y�a<ئa< �a<��a<��a<�a<J�a<j�a<Өa<�a<>�a<j�a<��a<ѩa<�a<H�a<e�a<��a<��a<�a<	�a<'�a<a�a<X�a<��a<��a<��a<ȫa<�a<
�a< �a</�a<�a<O�a<U�a<O�a<o�a<J�a<X�a<Z�a<d�a<_�a<j�a<Q�a<A�a<g�a<)�a<P�a<�a<�a<�a<�a<�a<īa<��a<��a<��a<g�a<Q�a<B�a<�a<�a<��a<��a<w�a<=�a<�a<�a<��a<��a<y�a<8�a<��a<ܨa<��a<�a<)�a<�a<��a<c�a< �a<�a<��a<P�a<.�a<��a<��a<I�a<ޤa<��a<&�a<�a<��a<D�a<�a<}�a<%�a<��a<��a<�a<àa<I�a<ҟa<}�a<��a<��a<&�a<��a<H�a<ٜa<v�a<��a<��a<!�a<a<G�a<ܙa<��a<�a<��a<	�a<��a<+�a<ɖa<b�a<�a<��a<��a<ʔa<I�a<�a<��a<�a<̒a<I�a<�a<��a<5�a<�a<��a<N�a<�a<��a<E�a<�a<a<x�a<N�a<�a<��a<s�a<A�a<
�a<�a<��a<y�a<p�a<+�a<-�a<�a<܋a<ۋa<��a<��a<��a<~�a<q�a<x�a<a�a<W�a<��a<Z�a<��a<x�a<��a<��a<��a<ߋa<�  �  �a<+�a<7�a<e�a<��a<��a<֌a<�a<L�a<j�a<��a<�a<2�a<}�a<��a<�a<O�a<��a<ޏa<:�a<��a<�a<B�a<��a<�a<l�a<Ւa<H�a<��a<�a<a�a<�a<L�a<��a<,�a<��a<�a<z�a<�a<k�a<�a<k�a<�a<\�a<Śa<G�a<��a<"�a<��a<�a<��a<��a<t�a<�a<m�a<�a<V�a<Ġa<)�a<��a<��a<r�a<ߢa<:�a<��a<��a<w�a<Τa<6�a<��a<�a<5�a<z�a<�a<�a<s�a<��a<��a<A�a<��a<ͨa<�a<A�a<�a<��a<�a<�a<C�a<W�a<��a<��a<�a<�a<�a<@�a<e�a<��a<��a<��a<ҫa<�a<�a<��a<'�a<*�a<1�a<4�a<N�a<a�a<[�a<s�a<|�a<q�a<]�a<a�a<f�a<M�a<V�a<*�a<C�a<$�a<#�a<�a<�a<�a<�a<̫a<��a<��a<h�a<6�a<�a<�a<�a<��a<��a<k�a<I�a<'�a<��a<Ωa<��a<_�a<%�a<��a<ڨa<��a<V�a<�a<�a<��a<u�a<C�a<��a<��a<S�a<$�a<ҥa<��a<8�a<֤a<��a<9�a<��a<��a<C�a<�a<��a<:�a<ˡa<s�a<��a<��a<3�a<֟a<n�a<��a<��a<)�a<ĝa<\�a<�a<{�a<�a<��a<�a<��a<I�a<͙a<Y�a<�a<��a<�a<��a<T�a<ٖa<d�a<�a<��a<�a<��a<=�a<ޓa<��a<�a<ƒa<J�a<�a<��a<[�a<��a<��a<I�a<ߏa<��a<G�a<�a<��a<f�a<-�a<�a<a<��a<O�a<�a<یa<��a<v�a<h�a<6�a<�a<�a<ۋa<͋a<��a<��a<��a<��a<o�a<o�a<v�a<c�a<w�a<[�a<��a<��a<��a<��a<��a<�a<�  �  /�a<H�a<��a<��a<ɋa<�a<�a<P�a<i�a<��a<�a<�a<i�a<��a<�a<$�a<��a<Ɏa<6�a<}�a<͏a<<�a<��a<��a<O�a<��a<%�a<k�a<��a<3�a<Ǔa<�a<��a<
�a<|�a<��a<Z�a<�a<4�a<×a<0�a<��a<%�a<��a<$�a<��a<+�a<��a<
�a<��a<�a<z�a<ܝa<N�a<Ğa<*�a<��a<�a<��a<��a<��a<Ρa<I�a<��a<�a<��a<̣a<<�a<��a<�a<A�a<��a<��a<+�a<��a<ئa<7�a<s�a<��a<��a<�a<��a<��a<ܨa<�a<Z�a<r�a<��a<�a<��a<8�a<F�a<i�a<��a<��a<Ϫa<۪a<��a<	�a<7�a<D�a<n�a<��a<t�a<��a<��a<��a<̫a<��a<֫a<ͫa<̫a<��a<ӫa<«a<��a<ɫa<��a<ȫa<��a<��a<y�a<h�a<k�a<6�a<8�a<�a<�a<٪a<۪a<��a<��a<w�a<9�a<1�a<�a<̩a<��a<k�a<H�a<�a<��a<��a<��a<h�a<-�a<�a<��a<��a<Y�a<�a<�a<��a<U�a<��a<ݥa<q�a<9�a<��a<��a<h�a<��a<£a<C�a<�a<��a<A�a<�a<��a<;�a< a<��a<�a<��a<C�a<��a<w�a<��a<��a<�a<��a<0�a<ʛa<^�a<�a<��a<�a<��a<;�a<��a<h�a<̗a<l�a<�a<��a<�a<��a<J�a<��a<x�a<��a<��a<4�a<˒a<h�a<�a<��a<-�a<ސa<~�a<>�a<͏a<~�a<B�a<Վa<��a<<�a<�a<ƍa<d�a<,�a<݌a<��a<e�a<F�a<�a<�a<ʋa<��a<�a<L�a<6�a<%�a<�a<�a<ӊa<��a<��a<��a<��a<��a<��a<��a<Ɗa<��a<Ǌa<Ċa<؊a<�a<��a<�  �  /�a<F�a<v�a<��a<��a<ߋa<�a<G�a<��a<��a<��a<)�a<n�a<��a<��a<@�a<��a<ӎa<�a<s�a<ۏa<.�a<��a<ސa<Q�a<��a<�a<q�a<�a<Q�a<Ɠa<&�a<��a<�a<d�a<ϕa<V�a<Ֆa<I�a<ȗa<@�a<Øa<&�a<��a<&�a<��a<�a<�a<��a<z�a<��a<Z�a<ڝa<T�a<Ӟa<A�a<��a<+�a<��a< �a<`�a<�a<H�a<��a<�a<z�a<�a<A�a<��a<�a<Y�a<��a<��a<A�a<��a<ئa<�a<X�a<��a<�a<3�a<}�a<��a<�a<�a<Q�a<z�a<��a<Ωa<��a<&�a<R�a<j�a<��a<��a<תa<�a<�a<%�a<@�a<O�a<\�a<c�a<��a<��a<��a<��a<��a<ʫa<ѫa<ɫa<Ϋa<۫a<׫a<ѫa<ƫa<��a<��a<��a<��a<��a<��a<z�a<k�a<V�a<9�a<�a<�a<�a<Ъa<��a<��a<o�a<W�a<�a<�a<ةa<��a<��a<]�a</�a<�a<ɨa<��a<^�a<;�a<��a<ʧa<��a<[�a<�a<�a<��a<`�a<�a<ۥa<��a<6�a<�a<��a<8�a<��a<��a<X�a<	�a<��a<`�a<�a<��a<=�a<ܠa<m�a< �a<��a<:�a<ڞa<W�a<��a<��a<'�a<��a<C�a<ڛa<b�a<�a<p�a<�a<��a<,�a<��a<L�a<�a<q�a< �a<��a<*�a<��a<H�a<єa<j�a<��a<}�a<�a<ǒa<]�a<�a<��a<F�a<�a<��a<5�a<֏a<��a<&�a<܎a<��a<G�a<�a<��a<j�a<3�a<�a<��a<��a<O�a<�a<�a<��a<��a<q�a<K�a<*�a<�a<�a<�a<Ίa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ϊa<�a<�a<�a<�  �  $�a<X�a<j�a<��a<��a<�a<(�a<.�a<��a<��a<��a<*�a<Y�a<��a<�a<5�a<}�a<ގa<0�a<��a<܏a<�a<��a<�a<X�a<��a<�a<~�a<ߒa<L�a<��a<-�a<��a<	�a<��a<�a<w�a<Ȗa<T�a<��a<(�a<��a<)�a<��a<�a<��a<�a<��a<�a<i�a<�a<a�a<�a<N�a<��a<2�a<��a<�a<��a<�a<j�a<�a<>�a<��a<.�a<r�a<�a<2�a<��a<�a<J�a<��a<�a<O�a<��a<�a<)�a<x�a<��a<�a<<�a<e�a<��a<�a<�a<K�a<w�a<��a<ͩa<�a<�a<O�a<|�a<��a<��a<Ȫa<�a<��a<�a<+�a<P�a<w�a<o�a<��a<��a<��a<��a<��a<ɫa<īa<ثa<ʫa<իa<��a<ͫa<̫a<��a<Ыa<��a<��a<��a<��a<x�a<M�a<P�a<.�a<+�a<�a<�a<˪a<��a<��a<U�a<_�a<�a<�a<٩a<��a<~�a<J�a<$�a<�a<Өa<��a<o�a<<�a<�a<�a<��a<b�a<�a<֦a<��a<U�a<�a<��a<��a<0�a<��a<��a<R�a<�a<��a<d�a<�a<��a<P�a<�a<��a<-�a<�a<d�a<�a<��a<*�a<�a<^�a<�a<��a<�a<��a<2�a<ʛa<Y�a<�a<y�a<$�a<��a<)�a<՘a<D�a<�a<b�a<�a<��a<�a<��a<>�a<ߔa<_�a<�a<��a<9�a<ђa<S�a<�a<��a<>�a<�a<��a</�a<ҏa<��a<%�a<��a<}�a<E�a<�a<��a<{�a<%�a<�a<��a<x�a<:�a<�a<��a<��a<��a<Y�a<_�a<;�a<	�a<�a<��a<ފa<��a<��a<��a<��a<��a<��a<��a<��a<ʊa<��a<Њa<�a<�a<�a<�  �  /�a<W�a<n�a<��a<a<�a<�a<J�a<s�a<��a<�a<�a<r�a<��a<��a<:�a<��a<Ǝa<3�a<t�a<ԏa<3�a<��a<��a<O�a<��a<�a<~�a<�a<J�a<��a<�a<��a<��a<m�a<��a<P�a<ٖa<?�a<ɗa<;�a<��a<6�a<��a<�a<��a<�a<��a<��a<��a<�a<p�a<ڝa<T�a<Ξa<E�a<��a<'�a<��a<��a<x�a<ѡa<N�a<��a<�a<��a<٣a<7�a<��a<��a<P�a<��a<��a<8�a<��a<Φa<�a<c�a<��a<��a<&�a<w�a<��a<�a<�a<K�a<{�a<��a<ߩa<��a<)�a<M�a<e�a<��a<��a<تa<�a<�a<$�a<?�a<D�a<c�a<|�a<�a<��a<��a<��a<ëa<��a<ȫa<ԫa<ӫa<ϫa<իa<ƫa<ëa<��a<��a<��a<��a<��a<��a<k�a<i�a<N�a<8�a<)�a<�a<�a<Ԫa<��a<��a<q�a<C�a<%�a<�a<ǩa<��a<��a<d�a<)�a<�a<��a<��a<_�a<3�a<�a<��a<��a<X�a<�a<զa<��a<]�a<�a<ӥa<y�a<A�a<�a<��a<I�a<�a<��a<N�a<
�a<��a<Q�a<��a<��a<0�a<Рa<z�a<�a<��a<A�a<a<m�a<��a<��a<"�a<��a<I�a<՛a<b�a<�a<��a<�a<��a<)�a<��a<V�a<ٗa<g�a< �a<��a<"�a<��a<K�a<Ȕa<o�a<�a<��a<$�a<��a<j�a<��a<��a<>�a<�a<��a</�a<׏a<��a<8�a<Ԏa<��a<C�a<�a<��a<_�a<5�a<�a<a<�a<N�a<�a<�a<Ëa<��a<w�a<K�a</�a<�a<��a<�a<ڊa<Ɗa<��a<��a<��a<��a<��a<��a<��a<��a<��a<Њa<ڊa<�a<�a<�  �  2�a<>�a<|�a<��a<��a<�a<�a<i�a<t�a<��a<�a<$�a<t�a<��a<�a<�a<��a<Ɏa<5�a<r�a<ڏa<L�a<x�a<��a<<�a<��a<�a<n�a<�a<=�a<̓a<�a<��a<��a<q�a<��a<H�a<�a<,�a<��a<8�a<��a<-�a<��a<0�a<��a<"�a<��a<��a<��a<�a<�a<ѝa<`�a<��a<5�a<��a<�a<��a<�a<��a<ˡa<^�a<��a<�a<��a<Σa<M�a<��a<�a<N�a<��a<��a<#�a<��a<ɦa<5�a<o�a<��a< �a<�a<��a<��a<�a<�a<E�a<��a<��a<�a<�a<<�a<X�a<c�a<��a<��a<�a<Ҫa<�a<�a<<�a<Q�a<V�a<�a<�a<��a<��a<��a<��a<īa<ثa<��a<ӫa<ƫa<߫a<��a<��a<ǫa<��a<ëa<��a<��a<{�a<c�a<v�a<B�a<;�a<�a<�a<�a<̪a<��a<��a<��a<D�a<%�a<��a<өa<��a<j�a<j�a<
�a<�a<��a<��a<]�a<:�a<�a<��a<��a<E�a<%�a<٦a<��a<]�a<�a<�a<j�a<B�a<�a<��a<f�a<�a<��a<;�a<�a<��a<O�a<��a<��a<H�a<Ǡa<��a< �a<��a<Y�a<a<{�a<�a<��a<�a<��a<?�a<��a<m�a<�a<��a<��a<��a<1�a<��a<a�a<Ηa<}�a<�a<��a< �a<��a<H�a<��a<y�a<�a<��a<0�a<��a<p�a<�a<��a</�a<�a<��a<)�a<�a<s�a<C�a<Ɏa<��a<N�a<�a<ƍa<^�a<?�a<Ԍa<Ìa<i�a<K�a<�a<ۋa<Ƌa<��a<��a<C�a<1�a<�a<��a<��a<��a<Ǌa<��a<��a<��a<��a<��a<��a<��a<��a<��a<Ɗa<ӊa<�a<�a<�  �  5�a<O�a<m�a<��a<��a<��a<#�a<4�a<|�a<��a<�a<'�a<g�a<��a<	�a<3�a<��a<Ԏa<,�a<��a<׏a<#�a<��a<�a<F�a<��a<�a<}�a<�a<C�a<��a<'�a<��a<��a<l�a<�a<S�a<Ɩa<Q�a<ȗa<)�a<��a</�a<��a<�a<��a<�a<��a<�a<s�a<��a<i�a<�a<U�a<a<K�a<a<�a<��a<�a<r�a<ޡa<D�a<��a<0�a<s�a<ޣa<=�a<��a<��a<J�a<��a<��a<K�a<��a<Ӧa<$�a<f�a<��a<�a<4�a<n�a<��a<�a<�a<H�a<��a<��a<֩a<�a<�a<L�a<s�a<��a<��a<תa<�a<!�a<&�a<4�a<R�a<n�a<x�a<��a<��a<��a<ūa<��a<ʫa<ȫa<ҫa<ثa<ƫa<��a<Ыa<īa<��a<��a<��a<��a<��a<��a<w�a<V�a<C�a<?�a<"�a<�a<��a<ªa<��a<��a<[�a<K�a<*�a<�a<֩a<��a<��a<o�a<#�a<�a<ʨa<��a<k�a<6�a<�a<اa<��a<P�a<#�a<֦a<��a<Z�a<
�a<ʥa<��a<2�a<�a<��a<Q�a<��a<��a<`�a<	�a<��a<L�a<��a<��a<6�a<Ԡa<d�a<#�a<��a<4�a<Ӟa<f�a<�a<��a<�a<��a<R�a<̛a<a�a<�a<��a<�a<��a<-�a<טa<F�a<ޗa<m�a<��a<��a<�a<��a<E�a<۔a<^�a<��a<��a<'�a<��a<Y�a<�a<��a<3�a<�a<��a<,�a<ݏa<��a</�a<��a<��a<B�a<��a<��a<l�a<4�a<�a<͌a<��a<C�a<�a<�a<��a<��a<`�a<Y�a<E�a<�a<�a<�a<؊a<ˊa<��a<��a<��a<��a<��a<��a<��a<��a<��a<̊a<�a<�a<�a<�  �  �a<]�a<[�a<��a<��a<ًa<(�a<<�a<��a<��a<�a<,�a<t�a<��a<�a<N�a<��a<�a<)�a<}�a<�a<'�a<��a<Аa<]�a<��a<�a<��a<Ԓa<_�a<��a<-�a<��a<�a<q�a<ԕa<d�a<��a<P�a<��a<=�a<��a<#�a<��a<�a<��a<��a<��a<	�a<z�a<�a<U�a<�a<K�a<۞a<B�a<��a<2�a<��a<�a<_�a<�a<R�a<��a<!�a<`�a<��a<�a<��a<�a<S�a<��a<ۥa<K�a<}�a<�a<�a<f�a<��a<�a<:�a<R�a<��a<بa<�a<K�a<f�a<éa<��a<�a<#�a<_�a<x�a<��a<ªa<˪a< �a<��a<)�a<G�a<O�a<s�a<g�a<��a<��a<��a<��a<��a<ѫa<��a<ޫa<��a<ݫa<īa<ūa<ūa<��a<��a<��a<��a<��a<��a<q�a<Q�a<^�a<(�a</�a<�a<�a<Ъa<��a<��a<d�a<c�a<�a<�a<۩a<��a<��a<H�a<=�a<��a<רa<��a<h�a<H�a<��a<ާa<v�a<f�a<
�a<Ӧa<��a<I�a<&�a<��a<��a<-�a<�a<��a<=�a<�a<��a<_�a<�a<��a<Z�a<�a<��a<�a<�a<W�a<�a<��a<;�a<�a<R�a<�a<��a</�a<��a<>�a<�a<W�a<�a<n�a<!�a<��a<1�a<Șa<2�a<��a<O�a<�a<��a<%�a<��a<(�a<۔a<T�a<�a<��a<'�a<Βa<P�a<	�a<��a<O�a<ڐa<��a</�a<��a<��a<�a<�a<��a<T�a< �a<��a<~�a<(�a<�a<��a<��a<V�a<�a<��a<��a<��a<h�a<_�a<*�a<�a<
�a<͊a<�a<��a<Êa<��a<��a<��a<��a<��a<��a<��a<��a<̊a<��a<�a<"�a<�  �  �a<X�a<z�a<��a<ɋa<�a<�a<R�a<w�a<��a<��a<-�a<j�a<��a<��a<=�a<��a<��a<8�a<x�a<ӏa<=�a<��a<�a<Q�a<��a<%�a<|�a<̒a<G�a<��a<'�a<��a<�a<q�a<��a<P�a<Ζa<=�a<��a<4�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<�a<r�a<�a<U�a<˞a<C�a<��a<%�a<��a<�a<}�a<ӡa<N�a<��a<�a<~�a<ߣa<5�a<��a<�a<A�a<��a<�a<9�a<��a<Φa<.�a<l�a<��a<�a<1�a<f�a<��a<Ҩa<�a<`�a<k�a<��a<کa<	�a<3�a<O�a<h�a<��a<ªa<ͪa<�a<�a<#�a<<�a<Q�a<p�a<{�a<��a<��a<��a<��a<ȫa<��a<ͫa<ثa<��a<˫a<ʫa<ƫa<��a<��a<��a<��a<��a<��a<y�a<q�a<_�a<H�a< �a<*�a<�a<�a<۪a<��a<��a<y�a<G�a<#�a<�a<ܩa<��a<��a<b�a<-�a<��a<ըa<��a<c�a<3�a<�a<ҧa<��a<[�a<�a<�a<��a<B�a<�a<ĥa<��a<3�a<ݤa<��a<_�a<�a<��a<L�a<��a<��a<G�a<�a<��a<3�a<֠a<t�a<
�a<��a<D�a<Ȟa<o�a<�a<��a< �a<��a<I�a<ӛa<c�a<�a<��a<�a<��a<5�a<��a<P�a<ޗa<e�a<�a<��a<�a<��a<8�a<ɔa<_�a<�a<��a<-�a<��a<Y�a< �a<��a<;�a<Ӑa<��a<D�a<Ǐa<��a<2�a<�a<��a<D�a<�a<a<~�a<*�a<��a<��a<~�a<K�a<�a<�a<a<��a<|�a<X�a<0�a<"�a<�a<�a<ފa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<Ŋa<��a<��a<�a<�  �  J�a<9�a<w�a<��a<ŋa<�a<�a<P�a<u�a<Όa<�a<,�a<p�a<��a<�a<0�a<��a<͎a<)�a<��a<ԏa<9�a<~�a<��a<I�a<��a<�a<j�a<��a<8�a<��a<�a<��a<��a<Y�a<�a<9�a<ٖa</�a<Ηa<!�a<��a<7�a<��a<1�a<��a<!�a<��a<�a<��a<�a<��a<̝a<n�a<ƞa<N�a<ǟa<�a<��a<�a<��a<סa<T�a<��a<�a<��a<ͣa<N�a<��a<��a<X�a<��a<�a<)�a<��a<��a<�a<U�a<��a<�a<�a<y�a<��a<��a<�a<?�a<��a<��a<�a<��a<0�a<P�a<}�a<��a<��a<�a<�a<)�a<%�a<;�a<\�a<V�a<��a<��a<��a<��a<��a<ȫa<��a<׫a<��a<�a<ʫa<��a<ɫa<��a<ūa<��a<��a<{�a<��a<t�a<h�a<V�a<B�a<S�a<�a<�a<�a<תa<��a<��a<w�a<D�a<B�a<��a<۩a<��a<��a<y�a< �a<�a<èa<��a<~�a<3�a<	�a<��a<��a<S�a<!�a<Ӧa<��a<s�a<��a<ϥa<m�a<4�a<�a<��a<P�a<ܣa<��a<>�a<�a<��a<W�a<��a<�a<H�a<àa<��a<�a<��a<K�a<ƞa<�a<�a<��a<�a<��a<W�a<ʛa<|�a<ښa<��a<	�a<��a<1�a<��a<_�a<̗a<~�a<�a<��a<*�a<��a<N�a<��a<j�a<ܓa<��a<�a<��a<a�a<�a<��a<+�a<��a<|�a<#�a<�a<x�a<B�a<юa<��a<F�a<�a<��a<_�a<I�a<�a<֌a<��a<K�a<#�a<ۋa<ۋa<��a<|�a<G�a<5�a<"�a<�a<�a<��a<݊a<��a<��a<��a<��a<��a<x�a<��a<��a<Ċa<��a<׊a<�a<�a<�  �  +�a<B�a<s�a<��a<��a<�a<#�a<M�a<��a<��a<�a<4�a<n�a<��a<��a<9�a<��a<܎a<0�a<��a<ۏa<:�a<��a<�a<G�a<��a<�a<p�a<�a<8�a<��a<�a<��a<��a<o�a<�a<V�a<͖a<1�a<ŗa<%�a<��a<%�a<��a<&�a<��a<�a<��a<�a<��a<��a<|�a<ݝa<f�a<Ǟa<>�a<��a<�a<��a< �a<��a<�a<S�a<��a<�a<y�a<ڣa<C�a<��a<�a<K�a<��a<��a</�a<��a<զa<#�a<g�a<��a<�a<#�a<m�a<��a<�a<�a<?�a<��a<��a<ԩa<�a<7�a<T�a<|�a<��a<��a<�a<�a<�a<$�a<<�a<`�a<c�a<��a<��a<��a<��a<��a<��a<ȫa<ϫa<��a<Ϋa<ƫa<��a<˫a<��a<��a<��a<��a<��a<��a<i�a<p�a<W�a<A�a<5�a<�a<
�a<�a<̪a<��a<��a<u�a<S�a<4�a<��a<�a<��a<��a<[�a<(�a<
�a<Ѩa<��a<w�a<;�a<
�a<ѧa<��a<Q�a<!�a<Ҧa<��a<W�a<��a<ɥa<x�a<'�a<�a<��a<R�a<��a<��a<@�a<�a<��a<L�a<�a<��a<=�a<Ѡa<p�a<�a<��a<F�a<֞a<y�a<��a<��a<�a<��a<?�a<͛a<r�a<�a<��a<�a<��a<:�a<Ƙa<K�a<ٗa<s�a<�a<��a<�a<��a<A�a<��a<_�a<��a<��a<(�a<��a<U�a<�a<��a<*�a<�a<�a<#�a<�a<�a<,�a<�a<��a<I�a<�a<��a<o�a<=�a<�a<��a<�a<L�a<'�a<�a<͋a<��a<{�a<Z�a<.�a<�a< �a<�a<Ŋa<a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ߊa<�a<�a<�  �  �a<\�a<k�a<��a<a<�a<$�a<C�a<��a<��a<��a<0�a<q�a<ˍa<��a<`�a<��a<�a<3�a<q�a<��a<2�a<��a<�a<S�a<��a<�a<��a<Òa<\�a<��a</�a<��a<�a<d�a<ϕa<J�a<��a<O�a<��a<@�a<��a<�a<��a<�a<��a<�a<��a<�a<�a<��a<i�a<��a<P�a<�a<R�a<��a<B�a<��a<�a<u�a<ݡa<L�a<��a<"�a<s�a<�a<2�a<��a<�a<?�a<��a<�a<M�a<~�a<ʦa<�a<X�a<��a<�a<<�a<]�a<��a<Ȩa<�a<W�a<n�a<��a<ѩa<�a<,�a<V�a<e�a<��a<Ǫa<Ъa<�a<�a<>�a<H�a<R�a<v�a<s�a<��a<��a<��a<��a<��a<ͫa<��a<�a<��a<ԫa<ȫa<̫a<«a<��a<��a<��a<��a<z�a<�a<z�a<T�a<Y�a<�a</�a<�a<�a<Ԫa<��a<��a<j�a<S�a<�a<�a<ߩa<��a<��a<_�a<O�a<��a<ިa<��a<\�a<@�a<�a<קa<��a<\�a<�a<�a<��a<9�a<#�a<��a<��a<1�a<֤a<��a<8�a<�a<��a<^�a<��a<��a<I�a<ޡa<��a<*�a<�a<j�a<�a<��a<?�a<Ԟa<f�a<�a<��a<5�a<Ĝa<Q�a<�a<b�a<�a<��a<�a<��a<.�a<ɘa<E�a<�a<b�a<�a<~�a<�a<��a<2�a<ޔa<U�a<�a<z�a<�a<��a<T�a<�a<��a<N�a<ʐa<��a<;�a<ʏa<��a<*�a<�a<��a<L�a<�a<��a<��a<-�a<�a<��a<��a<W�a<�a<��a<��a<��a<s�a<Z�a<-�a<�a<�a<܊a<�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ʊa<�a<�a<�a<�  �  +�a<H�a<c�a<��a<��a<�a<�a<P�a<��a<Ōa<��a<0�a<s�a<��a<�a<@�a<��a<�a<7�a<��a<�a<2�a<��a<��a<R�a<��a<	�a<p�a<ܒa<P�a<��a<�a<��a<�a<o�a<�a<W�a<͖a<;�a<��a<.�a<��a<%�a<��a<�a<��a<�a<��a<�a<��a<��a<}�a<�a<Z�a<Ԟa<5�a<��a<)�a<��a<
�a<��a<�a<Z�a<��a< �a<��a<�a<9�a<��a<�a<F�a<��a<إa<7�a<��a<٦a<�a<f�a<��a<�a<#�a<V�a<��a<ڨa<�a<=�a<x�a<��a<�a<�a<*�a<d�a<��a<��a<��a<ܪa<�a<��a<�a<E�a<U�a<p�a<��a<��a<��a<��a<��a<��a<ǫa<��a<˫a<ʫa<Ыa<��a<��a<��a<��a<��a<��a<��a<��a<{�a<^�a<G�a<Q�a<4�a<�a<��a<�a<Ҫa<��a<��a<w�a<Z�a<9�a<�a<ީa<��a<��a<K�a</�a<�a<רa<��a<y�a<G�a<�a<ȧa<��a<\�a<�a<Цa<��a<Q�a<�a<��a<u�a<0�a<�a<��a<L�a<��a<��a<K�a<�a<��a<K�a<�a<��a<.�a<ܠa<r�a<�a<��a<L�a<ݞa<z�a<�a<��a<(�a<��a<6�a<؛a<k�a<��a<��a<�a<��a<,�a<ǘa<R�a<�a<i�a<�a<��a<�a<��a<&�a<ǔa<_�a<��a<��a<'�a<Œa<X�a<�a<��a<D�a<ܐa<}�a<!�a<ԏa<��a<9�a<��a<��a<Y�a<�a<a<z�a<9�a<�a<��a<x�a<T�a<�a<��a<Ջa<��a<�a<K�a<<�a<�a< �a<׊a<ъa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<Ǌa<͊a<ފa<�a<�  �  2�a<A�a<|�a<��a<��a<��a<�a<N�a<k�a<Ča<�a<)�a<y�a<��a<�a<F�a<��a<юa<*�a<��a<ďa</�a<��a<��a<;�a<��a<�a<u�a<�a</�a<��a<#�a<~�a<��a<S�a<ҕa<F�a<ǖa<5�a<̗a<(�a<��a<7�a<��a<3�a<��a<�a<��a<��a<x�a<�a<��a<ӝa<g�a<מa<R�a<˟a<*�a<��a<��a<��a<աa<D�a<��a<#�a<{�a<ͣa<T�a<��a<��a<C�a<��a<��a<2�a<��a<ʦa<
�a<L�a<��a<ߧa<(�a<x�a<��a<�a<�a<D�a<��a<��a<�a<�a<'�a<B�a<s�a<��a<��a<�a<��a<-�a<0�a<J�a<U�a<[�a<��a<x�a<��a<��a<ɫa<��a<ȫa<׫a<«a<իa<��a<ʫa<ͫa<��a<��a<��a<��a<~�a<��a<n�a<s�a<f�a<8�a<;�a<�a<�a<��a<��a<Īa<��a<u�a<;�a<9�a<��a<ةa<��a<��a<}�a<6�a<�a<ƨa<��a<s�a<$�a<��a<̧a<��a<D�a<+�a<ئa<��a<`�a<��a<ѥa<��a<$�a<�a<�a<:�a<�a<��a<D�a<�a<��a<B�a<��a<��a<J�a<ʠa<j�a<�a<��a<9�a<ƞa<�a<�a<��a<+�a<Üa<Z�a<؛a<w�a<�a<��a<�a<��a<*�a<ʘa<M�a<͗a<��a<�a<��a<�a<��a<J�a<a<Z�a<�a<y�a<�a<��a<O�a<��a<��a<(�a<�a<��a<(�a<�a<q�a<9�a<�a<��a<8�a<��a<��a<e�a<L�a<��a<ٌa<��a<Y�a<�a<��a<Ջa<��a<w�a<E�a<H�a<�a<�a<�a<Ǌa<Ɋa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<�a<��a<��a<�  �  +�a<H�a<c�a<��a<��a<�a<�a<P�a<��a<Ōa<��a<0�a<s�a<��a<�a<@�a<��a<�a<7�a<��a<�a<2�a<��a<��a<R�a<��a<	�a<p�a<ܒa<P�a<��a<�a<��a<�a<o�a<�a<W�a<͖a<;�a<��a<.�a<��a<%�a<��a<�a<��a<�a<��a<�a<��a<��a<}�a<�a<Z�a<Ԟa<5�a<��a<)�a<��a<
�a<��a<�a<Z�a<��a< �a<��a<�a<9�a<��a<�a<F�a<��a<إa<7�a<��a<٦a<�a<f�a<��a<�a<#�a<V�a<��a<ڨa<�a<=�a<x�a<��a<�a<�a<*�a<d�a<��a<��a<��a<ܪa<�a<��a<�a<E�a<U�a<p�a<��a<��a<��a<��a<��a<��a<ǫa<��a<˫a<ʫa<Ыa<��a<��a<��a<��a<��a<��a<��a<��a<{�a<^�a<G�a<Q�a<4�a<�a<��a<�a<Ҫa<��a<��a<w�a<Z�a<9�a<�a<ީa<��a<��a<K�a</�a<�a<רa<��a<y�a<G�a<�a<ȧa<��a<\�a<�a<Цa<��a<Q�a<�a<��a<u�a<0�a<�a<��a<L�a<��a<��a<K�a<�a<��a<K�a<�a<��a<.�a<ܠa<r�a<�a<��a<L�a<ݞa<z�a<�a<��a<(�a<��a<6�a<؛a<k�a<��a<��a<�a<��a<,�a<ǘa<R�a<�a<i�a<�a<��a<�a<��a<&�a<ǔa<_�a<��a<��a<'�a<Œa<X�a<�a<��a<D�a<ܐa<}�a<!�a<ԏa<��a<9�a<��a<��a<Y�a<�a<a<z�a<9�a<�a<��a<x�a<T�a<�a<��a<Ջa<��a<�a<K�a<<�a<�a< �a<׊a<ъa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<Ǌa<͊a<ފa<�a<�  �  �a<\�a<k�a<��a<a<�a<$�a<C�a<��a<��a<��a<0�a<q�a<ˍa<��a<`�a<��a<�a<3�a<q�a<��a<2�a<��a<�a<S�a<��a<�a<��a<Òa<\�a<��a</�a<��a<�a<d�a<ϕa<J�a<��a<O�a<��a<@�a<��a<�a<��a<�a<��a<�a<��a<�a<�a<��a<i�a<��a<P�a<�a<R�a<��a<B�a<��a<�a<u�a<ݡa<L�a<��a<"�a<s�a<�a<2�a<��a<�a<?�a<��a<�a<M�a<~�a<ʦa<�a<X�a<��a<�a<<�a<]�a<��a<Ȩa<�a<W�a<n�a<��a<ѩa<�a<,�a<V�a<e�a<��a<Ǫa<Ъa<�a<�a<>�a<H�a<R�a<v�a<s�a<��a<��a<��a<��a<��a<ͫa<��a<�a<��a<ԫa<ȫa<̫a<«a<��a<��a<��a<��a<z�a<�a<z�a<T�a<Y�a<�a</�a<�a<�a<Ԫa<��a<��a<j�a<S�a<�a<�a<ߩa<��a<��a<_�a<O�a<��a<ިa<��a<\�a<@�a<�a<קa<��a<\�a<�a<�a<��a<9�a<#�a<��a<��a<1�a<֤a<��a<8�a<�a<��a<^�a<��a<��a<I�a<ޡa<��a<*�a<�a<j�a<�a<��a<?�a<Ԟa<f�a<�a<��a<5�a<Ĝa<Q�a<�a<b�a<�a<��a<�a<��a<.�a<ɘa<E�a<�a<b�a<�a<~�a<�a<��a<2�a<ޔa<U�a<�a<z�a<�a<��a<T�a<�a<��a<N�a<ʐa<��a<;�a<ʏa<��a<*�a<�a<��a<L�a<�a<��a<��a<-�a<�a<��a<��a<W�a<�a<��a<��a<��a<s�a<Z�a<-�a<�a<�a<܊a<�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ʊa<�a<�a<�a<�  �  +�a<B�a<s�a<��a<��a<�a<#�a<M�a<��a<��a<�a<4�a<n�a<��a<��a<9�a<��a<܎a<0�a<��a<ۏa<:�a<��a<�a<G�a<��a<�a<p�a<�a<8�a<��a<�a<��a<��a<o�a<�a<V�a<͖a<1�a<ŗa<%�a<��a<%�a<��a<&�a<��a<�a<��a<�a<��a<��a<|�a<ݝa<f�a<Ǟa<>�a<��a<�a<��a< �a<��a<�a<S�a<��a<�a<y�a<ڣa<C�a<��a<�a<K�a<��a<��a</�a<��a<զa<#�a<g�a<��a<�a<#�a<m�a<��a<�a<�a<?�a<��a<��a<ԩa<�a<7�a<T�a<|�a<��a<��a<�a<�a<�a<$�a<<�a<`�a<c�a<��a<��a<��a<��a<��a<��a<ȫa<ϫa<��a<Ϋa<ƫa<��a<˫a<��a<��a<��a<��a<��a<��a<i�a<p�a<W�a<A�a<5�a<�a<
�a<�a<̪a<��a<��a<u�a<S�a<4�a<��a<�a<��a<��a<[�a<(�a<
�a<Ѩa<��a<w�a<;�a<
�a<ѧa<��a<Q�a<!�a<Ҧa<��a<W�a<��a<ɥa<x�a<'�a<�a<��a<R�a<��a<��a<@�a<�a<��a<L�a<�a<��a<=�a<Ѡa<p�a<�a<��a<F�a<֞a<y�a<��a<��a<�a<��a<?�a<͛a<r�a<�a<��a<�a<��a<:�a<Ƙa<K�a<ٗa<s�a<�a<��a<�a<��a<A�a<��a<_�a<��a<��a<(�a<��a<U�a<�a<��a<*�a<�a<�a<#�a<�a<�a<,�a<�a<��a<I�a<�a<��a<o�a<=�a<�a<��a<�a<L�a<'�a<�a<͋a<��a<{�a<Z�a<.�a<�a< �a<�a<Ŋa<a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ߊa<�a<�a<�  �  J�a<9�a<w�a<��a<ŋa<�a<�a<P�a<u�a<Όa<�a<,�a<p�a<��a<�a<0�a<��a<͎a<)�a<��a<ԏa<9�a<~�a<��a<I�a<��a<�a<j�a<��a<8�a<��a<�a<��a<��a<Y�a<�a<9�a<ٖa</�a<Ηa<!�a<��a<7�a<��a<1�a<��a<!�a<��a<�a<��a<�a<��a<̝a<n�a<ƞa<N�a<ǟa<�a<��a<�a<��a<סa<T�a<��a<�a<��a<ͣa<N�a<��a<��a<X�a<��a<�a<)�a<��a<��a<�a<U�a<��a<�a<�a<y�a<��a<��a<�a<?�a<��a<��a<�a<��a<0�a<P�a<}�a<��a<��a<�a<�a<)�a<%�a<;�a<\�a<V�a<��a<��a<��a<��a<��a<ȫa<��a<׫a<��a<�a<ʫa<��a<ɫa<��a<ūa<��a<��a<{�a<��a<t�a<h�a<V�a<B�a<S�a<�a<�a<�a<תa<��a<��a<w�a<D�a<B�a<��a<۩a<��a<��a<y�a< �a<�a<èa<��a<~�a<3�a<	�a<��a<��a<S�a<!�a<Ӧa<��a<s�a<��a<ϥa<m�a<4�a<�a<��a<P�a<ܣa<��a<>�a<�a<��a<W�a<��a<�a<H�a<àa<��a<�a<��a<K�a<ƞa<�a<�a<��a<�a<��a<W�a<ʛa<|�a<ښa<��a<	�a<��a<1�a<��a<_�a<̗a<~�a<�a<��a<*�a<��a<N�a<��a<j�a<ܓa<��a<�a<��a<a�a<�a<��a<+�a<��a<|�a<#�a<�a<x�a<B�a<юa<��a<F�a<�a<��a<_�a<I�a<�a<֌a<��a<K�a<#�a<ۋa<ۋa<��a<|�a<G�a<5�a<"�a<�a<�a<��a<݊a<��a<��a<��a<��a<��a<x�a<��a<��a<Ċa<��a<׊a<�a<�a<�  �  �a<X�a<z�a<��a<ɋa<�a<�a<R�a<w�a<��a<��a<-�a<j�a<��a<��a<=�a<��a<��a<8�a<x�a<ӏa<=�a<��a<�a<Q�a<��a<%�a<|�a<̒a<G�a<��a<'�a<��a<�a<q�a<��a<P�a<Ζa<=�a<��a<4�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<�a<r�a<�a<U�a<˞a<C�a<��a<%�a<��a<�a<}�a<ӡa<N�a<��a<�a<~�a<ߣa<5�a<��a<�a<A�a<��a<�a<9�a<��a<Φa<.�a<l�a<��a<�a<1�a<f�a<��a<Ҩa<�a<`�a<k�a<��a<کa<	�a<3�a<O�a<h�a<��a<ªa<ͪa<�a<�a<#�a<<�a<Q�a<p�a<{�a<��a<��a<��a<��a<ȫa<��a<ͫa<ثa<��a<˫a<ʫa<ƫa<��a<��a<��a<��a<��a<��a<y�a<q�a<_�a<H�a< �a<*�a<�a<�a<۪a<��a<��a<y�a<G�a<#�a<�a<ܩa<��a<��a<b�a<-�a<��a<ըa<��a<c�a<3�a<�a<ҧa<��a<[�a<�a<�a<��a<B�a<�a<ĥa<��a<3�a<ݤa<��a<_�a<�a<��a<L�a<��a<��a<G�a<�a<��a<3�a<֠a<t�a<
�a<��a<D�a<Ȟa<o�a<�a<��a< �a<��a<I�a<ӛa<c�a<�a<��a<�a<��a<5�a<��a<P�a<ޗa<e�a<�a<��a<�a<��a<8�a<ɔa<_�a<�a<��a<-�a<��a<Y�a< �a<��a<;�a<Ӑa<��a<D�a<Ǐa<��a<2�a<�a<��a<D�a<�a<a<~�a<*�a<��a<��a<~�a<K�a<�a<�a<a<��a<|�a<X�a<0�a<"�a<�a<�a<ފa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<Ŋa<��a<��a<�a<�  �  �a<]�a<[�a<��a<��a<ًa<(�a<<�a<��a<��a<�a<,�a<t�a<��a<�a<N�a<��a<�a<)�a<}�a<�a<'�a<��a<Аa<]�a<��a<�a<��a<Ԓa<_�a<��a<-�a<��a<�a<q�a<ԕa<d�a<��a<P�a<��a<=�a<��a<#�a<��a<�a<��a<��a<��a<	�a<z�a<�a<U�a<�a<K�a<۞a<B�a<��a<2�a<��a<�a<_�a<�a<R�a<��a<!�a<`�a<��a<�a<��a<�a<S�a<��a<ۥa<K�a<}�a<�a<�a<f�a<��a<�a<:�a<R�a<��a<بa<�a<K�a<f�a<éa<��a<�a<#�a<_�a<x�a<��a<ªa<˪a< �a<��a<)�a<G�a<O�a<s�a<g�a<��a<��a<��a<��a<��a<ѫa<��a<ޫa<��a<ݫa<īa<ūa<ūa<��a<��a<��a<��a<��a<��a<q�a<Q�a<^�a<(�a</�a<�a<�a<Ъa<��a<��a<d�a<c�a<�a<�a<۩a<��a<��a<H�a<=�a<��a<רa<��a<h�a<H�a<��a<ާa<v�a<f�a<
�a<Ӧa<��a<I�a<&�a<��a<��a<-�a<�a<��a<=�a<�a<��a<_�a<�a<��a<Z�a<�a<��a<�a<�a<W�a<�a<��a<;�a<�a<R�a<�a<��a</�a<��a<>�a<�a<W�a<�a<n�a<!�a<��a<1�a<Șa<2�a<��a<O�a<�a<��a<%�a<��a<(�a<۔a<T�a<�a<��a<'�a<Βa<P�a<	�a<��a<O�a<ڐa<��a</�a<��a<��a<�a<�a<��a<T�a< �a<��a<~�a<(�a<�a<��a<��a<V�a<�a<��a<��a<��a<h�a<_�a<*�a<�a<
�a<͊a<�a<��a<Êa<��a<��a<��a<��a<��a<��a<��a<��a<̊a<��a<�a<"�a<�  �  5�a<O�a<m�a<��a<��a<��a<#�a<4�a<|�a<��a<�a<'�a<g�a<��a<	�a<3�a<��a<Ԏa<,�a<��a<׏a<#�a<��a<�a<F�a<��a<�a<}�a<�a<C�a<��a<'�a<��a<��a<l�a<�a<S�a<Ɩa<Q�a<ȗa<)�a<��a</�a<��a<�a<��a<�a<��a<�a<s�a<��a<i�a<�a<U�a<a<K�a<a<�a<��a<�a<r�a<ޡa<D�a<��a<0�a<s�a<ޣa<=�a<��a<��a<J�a<��a<��a<K�a<��a<Ӧa<$�a<f�a<��a<�a<4�a<n�a<��a<�a<�a<H�a<��a<��a<֩a<�a<�a<L�a<s�a<��a<��a<תa<�a<!�a<&�a<4�a<R�a<n�a<x�a<��a<��a<��a<ūa<��a<ʫa<ȫa<ҫa<ثa<ƫa<��a<Ыa<īa<��a<��a<��a<��a<��a<��a<w�a<V�a<C�a<?�a<"�a<�a<��a<ªa<��a<��a<[�a<K�a<*�a<�a<֩a<��a<��a<o�a<#�a<�a<ʨa<��a<k�a<6�a<�a<اa<��a<P�a<#�a<֦a<��a<Z�a<
�a<ʥa<��a<2�a<�a<��a<Q�a<��a<��a<`�a<	�a<��a<L�a<��a<��a<6�a<Ԡa<d�a<#�a<��a<4�a<Ӟa<f�a<�a<��a<�a<��a<R�a<̛a<a�a<�a<��a<�a<��a<-�a<טa<F�a<ޗa<m�a<��a<��a<�a<��a<E�a<۔a<^�a<��a<��a<'�a<��a<Y�a<�a<��a<3�a<�a<��a<,�a<ݏa<��a</�a<��a<��a<B�a<��a<��a<l�a<4�a<�a<͌a<��a<C�a<�a<�a<��a<��a<`�a<Y�a<E�a<�a<�a<�a<؊a<ˊa<��a<��a<��a<��a<��a<��a<��a<��a<��a<̊a<�a<�a<�a<�  �  2�a<>�a<|�a<��a<��a<�a<�a<i�a<t�a<��a<�a<$�a<t�a<��a<�a<�a<��a<Ɏa<5�a<r�a<ڏa<L�a<x�a<��a<<�a<��a<�a<n�a<�a<=�a<̓a<�a<��a<��a<q�a<��a<H�a<�a<,�a<��a<8�a<��a<-�a<��a<0�a<��a<"�a<��a<��a<��a<�a<�a<ѝa<`�a<��a<5�a<��a<�a<��a<�a<��a<ˡa<^�a<��a<�a<��a<Σa<M�a<��a<�a<N�a<��a<��a<#�a<��a<ɦa<5�a<o�a<��a< �a<�a<��a<��a<�a<�a<E�a<��a<��a<�a<�a<<�a<X�a<c�a<��a<��a<�a<Ҫa<�a<�a<<�a<Q�a<V�a<�a<�a<��a<��a<��a<��a<īa<ثa<��a<ӫa<ƫa<߫a<��a<��a<ǫa<��a<ëa<��a<��a<{�a<c�a<v�a<B�a<;�a<�a<�a<�a<̪a<��a<��a<��a<D�a<%�a<��a<өa<��a<j�a<j�a<
�a<�a<��a<��a<]�a<:�a<�a<��a<��a<E�a<%�a<٦a<��a<]�a<�a<�a<j�a<B�a<�a<��a<f�a<�a<��a<;�a<�a<��a<O�a<��a<��a<H�a<Ǡa<��a< �a<��a<Y�a<a<{�a<�a<��a<�a<��a<?�a<��a<m�a<�a<��a<��a<��a<1�a<��a<a�a<Ηa<}�a<�a<��a< �a<��a<H�a<��a<y�a<�a<��a<0�a<��a<p�a<�a<��a</�a<�a<��a<)�a<�a<s�a<C�a<Ɏa<��a<N�a<�a<ƍa<^�a<?�a<Ԍa<Ìa<i�a<K�a<�a<ۋa<Ƌa<��a<��a<C�a<1�a<�a<��a<��a<��a<Ǌa<��a<��a<��a<��a<��a<��a<��a<��a<��a<Ɗa<ӊa<�a<�a<�  �  /�a<W�a<n�a<��a<a<�a<�a<J�a<s�a<��a<�a<�a<r�a<��a<��a<:�a<��a<Ǝa<3�a<t�a<ԏa<3�a<��a<��a<O�a<��a<�a<~�a<�a<J�a<��a<�a<��a<��a<m�a<��a<P�a<ٖa<?�a<ɗa<;�a<��a<6�a<��a<�a<��a<�a<��a<��a<��a<�a<p�a<ڝa<T�a<Ξa<E�a<��a<'�a<��a<��a<x�a<ѡa<N�a<��a<�a<��a<٣a<7�a<��a<��a<P�a<��a<��a<8�a<��a<Φa<�a<c�a<��a<��a<&�a<w�a<��a<�a<�a<K�a<{�a<��a<ߩa<��a<)�a<M�a<e�a<��a<��a<تa<�a<�a<$�a<?�a<D�a<c�a<|�a<�a<��a<��a<��a<ëa<��a<ȫa<ԫa<ӫa<ϫa<իa<ƫa<ëa<��a<��a<��a<��a<��a<��a<k�a<i�a<N�a<8�a<)�a<�a<�a<Ԫa<��a<��a<q�a<C�a<%�a<�a<ǩa<��a<��a<d�a<)�a<�a<��a<��a<_�a<3�a<�a<��a<��a<X�a<�a<զa<��a<]�a<�a<ӥa<y�a<A�a<�a<��a<I�a<�a<��a<N�a<
�a<��a<Q�a<��a<��a<0�a<Рa<z�a<�a<��a<A�a<a<m�a<��a<��a<"�a<��a<I�a<՛a<b�a<�a<��a<�a<��a<)�a<��a<V�a<ٗa<g�a< �a<��a<"�a<��a<K�a<Ȕa<o�a<�a<��a<$�a<��a<j�a<��a<��a<>�a<�a<��a</�a<׏a<��a<8�a<Ԏa<��a<C�a<�a<��a<_�a<5�a<�a<a<�a<N�a<�a<�a<Ëa<��a<w�a<K�a</�a<�a<��a<�a<ڊa<Ɗa<��a<��a<��a<��a<��a<��a<��a<��a<��a<Њa<ڊa<�a<�a<�  �  $�a<X�a<j�a<��a<��a<�a<(�a<.�a<��a<��a<��a<*�a<Y�a<��a<�a<5�a<}�a<ގa<0�a<��a<܏a<�a<��a<�a<X�a<��a<�a<~�a<ߒa<L�a<��a<-�a<��a<	�a<��a<�a<w�a<Ȗa<T�a<��a<(�a<��a<)�a<��a<�a<��a<�a<��a<�a<i�a<�a<a�a<�a<N�a<��a<2�a<��a<�a<��a<�a<j�a<�a<>�a<��a<.�a<r�a<�a<2�a<��a<�a<J�a<��a<�a<O�a<��a<�a<)�a<x�a<��a<�a<<�a<e�a<��a<�a<�a<K�a<w�a<��a<ͩa<�a<�a<O�a<|�a<��a<��a<Ȫa<�a<��a<�a<+�a<P�a<w�a<o�a<��a<��a<��a<��a<��a<ɫa<īa<ثa<ʫa<իa<��a<ͫa<̫a<��a<Ыa<��a<��a<��a<��a<x�a<M�a<P�a<.�a<+�a<�a<�a<˪a<��a<��a<U�a<_�a<�a<�a<٩a<��a<~�a<J�a<$�a<�a<Өa<��a<o�a<<�a<�a<�a<��a<b�a<�a<֦a<��a<U�a<�a<��a<��a<0�a<��a<��a<R�a<�a<��a<d�a<�a<��a<P�a<�a<��a<-�a<�a<d�a<�a<��a<*�a<�a<^�a<�a<��a<�a<��a<2�a<ʛa<Y�a<�a<y�a<$�a<��a<)�a<՘a<D�a<�a<b�a<�a<��a<�a<��a<>�a<ߔa<_�a<�a<��a<9�a<ђa<S�a<�a<��a<>�a<�a<��a</�a<ҏa<��a<%�a<��a<}�a<E�a<�a<��a<{�a<%�a<�a<��a<x�a<:�a<�a<��a<��a<��a<Y�a<_�a<;�a<	�a<�a<��a<ފa<��a<��a<��a<��a<��a<��a<��a<��a<ʊa<��a<Њa<�a<�a<�a<�  �  /�a<F�a<v�a<��a<��a<ߋa<�a<G�a<��a<��a<��a<)�a<n�a<��a<��a<@�a<��a<ӎa<�a<s�a<ۏa<.�a<��a<ސa<Q�a<��a<�a<q�a<�a<Q�a<Ɠa<&�a<��a<�a<d�a<ϕa<V�a<Ֆa<I�a<ȗa<@�a<Øa<&�a<��a<&�a<��a<�a<�a<��a<z�a<��a<Z�a<ڝa<T�a<Ӟa<A�a<��a<+�a<��a< �a<`�a<�a<H�a<��a<�a<z�a<�a<A�a<��a<�a<Y�a<��a<��a<A�a<��a<ئa<�a<X�a<��a<�a<3�a<}�a<��a<�a<�a<Q�a<z�a<��a<Ωa<��a<&�a<R�a<j�a<��a<��a<תa<�a<�a<%�a<@�a<O�a<\�a<c�a<��a<��a<��a<��a<��a<ʫa<ѫa<ɫa<Ϋa<۫a<׫a<ѫa<ƫa<��a<��a<��a<��a<��a<��a<z�a<k�a<V�a<9�a<�a<�a<�a<Ъa<��a<��a<o�a<W�a<�a<�a<ةa<��a<��a<]�a</�a<�a<ɨa<��a<^�a<;�a<��a<ʧa<��a<[�a<�a<�a<��a<`�a<�a<ۥa<��a<6�a<�a<��a<8�a<��a<��a<X�a<	�a<��a<`�a<�a<��a<=�a<ܠa<m�a< �a<��a<:�a<ڞa<W�a<��a<��a<'�a<��a<C�a<ڛa<b�a<�a<p�a<�a<��a<,�a<��a<L�a<�a<q�a< �a<��a<*�a<��a<H�a<єa<j�a<��a<}�a<�a<ǒa<]�a<�a<��a<F�a<�a<��a<5�a<֏a<��a<&�a<܎a<��a<G�a<�a<��a<j�a<3�a<�a<��a<��a<O�a<�a<�a<��a<��a<q�a<K�a<*�a<�a<�a<�a<Ίa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ϊa<�a<�a<�a<�  �  ��a<o�a<��a<��a<݊a<�a<+�a<l�a<��a<�a<�a<?�a<��a<��a<7�a<I�a<��a<��a<S�a<��a<��a<S�a<��a<)�a<r�a<ܐa<P�a<��a<Q�a<X�a<�a<M�a<Гa<@�a<��a<@�a<��a<4�a<j�a<�a<f�a<��a<��a<�a<r�a<˙a<f�a<��a<F�a<��a<'�a<��a<(�a<��a<	�a<��a<	�a<`�a<�a<R�a<Πa<%�a<��a<�a<Y�a<�a<)�a<��a<��a<s�a<��a<�a<s�a<��a<�a<4�a<��a<Цa<�a<a�a<�a<�a<�a<s�a<��a<��a<�a<��a<M�a<@�a<��a<��a<ǩa<��a<�a<2�a<-�a<�a<m�a<��a<��a<��a<�a<̪a<�a<��a<	�a<�a<�a<1�a<,�a<j�a<�a<-�a<,�a<�a<?�a<��a<!�a<�a<�a<֪a<Ϫa<ƪa<��a<ժa<x�a<t�a<>�a<$�a<�a<کa<ȩa<��a<��a<O�a<!�a<�a<ʨa<Ψa<i�a<W�a<�a<��a<ça<��a<Q�a<�a<��a<��a<q�a<A�a<��a<�a<G�a<>�a<Ҥa<��a<N�a<��a<ɣa<K�a<-�a<��a<u�a<�a<��a<y�a<��a<��a<�a<ӟa<K�a<�a<��a<�a<��a<D�a<ڜa<[�a<��a<��a<�a<��a<2�a<͙a<F�a<��a<m�a<�a<��a<�a<��a<C�a<�a<p�a<͔a<��a<��a<��a<,�a<�a<f�a<��a<��a< �a<�a<M�a<E�a<��a<e�a<�a<��a<r�a<�a<��a<m�a<�a<ތa<��a<Y�a<��a<��a<��a<j�a<-�a<�a<��a<��a<��a<g�a<P�a<8�a<�a<�a<��a<&�a<ŉa<҉a<Ήa<��a<�a<��a<�a<ȉa< �a<�a<�a<'�a<�a<�  �  R�a<[�a<��a<��a<�a<�a<G�a<l�a<��a<Ջa<�a<H�a<��a<ǌa<�a<X�a<��a<��a<U�a<��a< �a<_�a<ɏa<�a<��a<ސa<J�a<��a<�a<{�a<��a<Q�a<֓a<>�a<��a<,�a<��a<�a<��a<�a<��a<��a<\�a<ޘa<i�a<�a<h�a<ߚa<\�a<ța<D�a<��a<3�a<��a<�a<��a<�a<t�a<�a<^�a<Ơa<>�a<��a<�a<~�a<�a<?�a<��a<�a<A�a<��a<�a<a�a<��a<��a<.�a<��a<ʦa<�a<_�a<��a<ܧa<�a<L�a<c�a<��a<ߨa<�a<=�a<k�a<��a<��a<ϩa<��a<�a</�a<A�a<h�a<u�a<��a<��a<Īa<Ҫa<�a<��a<�a<�a<%�a<#�a<,�a<�a<#�a<0�a<7�a<%�a<�a<$�a<��a<�a<�a<��a<ߪa<Ȫa<ɪa<��a<��a<d�a<h�a<G�a<5�a<�a<��a<ǩa<��a<}�a<Z�a<*�a<�a<Ѩa<��a<y�a<S�a<$�a<��a<��a<��a<\�a<2�a<�a<��a<s�a<;�a<ޥa<��a<i�a<6�a<פa<��a<L�a<�a<��a<I�a<�a<��a<g�a<�a<��a<:�a<�a<��a<.�a<֟a<m�a<�a<��a<)�a<��a<O�a<ڜa<l�a<��a<��a<�a<��a<>�a<ƙa<_�a<�a<��a<�a<��a<#�a<��a<5�a<��a<i�a<�a<��a<�a<��a<&�a<ђa<_�a<��a<��a<,�a<ݐa<n�a<�a<��a<_�a<	�a<��a<b�a<�a<��a<o�a<"�a<ߌa<��a<V�a<�a<ދa<��a<q�a<6�a<�a<�a<��a<��a<�a<_�a<G�a<#�a<�a<�a<މa<މa<܉a<ǉa<a<Ήa<��a<҉a<ĉa<�a<�a< �a<*�a<6�a<�  �  G�a<��a<��a<��a<�a<��a<H�a<Z�a<��a<ċa<�a<A�a<��a<ӌa<�a<d�a<��a<��a<K�a<��a<
�a<R�a<ˏa<��a<��a<Րa<Z�a<Ǒa<�a<��a<�a<\�a<Гa<8�a<��a<)�a<��a<�a<��a<�a<y�a<�a<i�a<�a<_�a<�a<I�a<Ԛa<R�a<��a<O�a<��a<4�a<��a<�a<��a<��a<w�a<֟a<_�a<��a<B�a<��a<�a<y�a<��a<H�a<��a<�a<X�a<��a<�a<E�a<��a<�a<@�a<��a<Цa<�a<V�a<��a<ça<�a<<�a<��a<ƨa<Өa<�a<�a<o�a<��a<��a<ϩa<�a<�a<�a<L�a<P�a<~�a<��a<��a<êa<��a<��a<�a<�a< �a<�a<"�a<)�a<K�a<�a<?�a<!�a<�a<.�a<�a<�a<�a<�a<�a<�a<ɪa<��a<��a<��a<��a<j�a<E�a<-�a<��a<��a<��a<��a<l�a<X�a<#�a<��a<ݨa<��a<��a<F�a<�a<�a<��a<��a<P�a<4�a<˦a<��a<j�a<K�a<�a<��a<z�a<�a<�a<��a<F�a<�a<��a<`�a<��a<Ģa<O�a<�a<��a<G�a<�a<��a<3�a<��a<a�a<��a<��a<4�a<��a<Q�a<ʜa<h�a<��a<��a<�a<��a<?�a<��a<c�a<ޘa<t�a<�a<x�a<,�a<��a<^�a<Еa<c�a<�a<l�a<�a<��a<8�a<Вa<f�a<��a<��a<<�a<Őa<|�a<�a<͏a<y�a<��a<��a<;�a<�a<��a<p�a<#�a<Ќa<��a<D�a<�a<ǋa<��a<g�a<,�a<�a<͊a<͊a<��a<�a<G�a<8�a<#�a<�a<�a<ډa<�a<ǉa<��a<҉a<��a<щa<҉a<މa<ډa<��a<�a<�a<I�a<�  �  \�a<m�a<{�a<��a<�a<�a<F�a<d�a<��a<Ћa<�a<L�a<��a<Ќa<�a<b�a<��a<��a<P�a<��a<�a<V�a<��a<!�a<��a<ؐa<-�a<��a<�a<y�a<�a<_�a<ēa<0�a<��a<�a<��a<�a<��a<�a<u�a<��a<r�a<ݘa<V�a<�a<g�a<ؚa<\�a<̛a<;�a<��a<*�a<��a<�a<��a<�a<w�a<�a<[�a<Ƞa<2�a<��a<�a<y�a<�a<J�a<��a<�a<T�a<��a<��a<U�a<��a<�a<9�a<��a<Цa<
�a<N�a<��a<ӧa<�a<B�a<x�a<��a<Ҩa<�a<@�a<b�a<��a<��a<ɩa<�a<�a<7�a<L�a<d�a<~�a<��a<��a<��a<ͪa<�a<�a<�a<�a<(�a<(�a<�a<#�a<5�a<'�a<$�a<0�a<�a<�a<�a<��a<��a<�a<۪a<٪a<��a<��a<��a<v�a<H�a<M�a<9�a<�a<��a<��a<��a<w�a<S�a<.�a<�a<٨a<��a<��a<_�a<$�a<�a<��a<��a<T�a<%�a<�a<��a<m�a<�a<��a<��a<h�a<+�a<�a<��a<?�a< �a<��a<U�a<��a<��a<`�a<��a<��a<P�a<�a<��a<8�a<ԟa<e�a<�a<��a< �a<��a<F�a<�a<l�a<��a<��a<�a<��a<;�a<Ǚa<S�a<�a<~�a<	�a<��a<.�a<��a<,�a<̕a<Z�a<�a<|�a<
�a<��a<1�a<˒a<f�a<��a<��a<3�a<Րa<k�a<�a<��a<I�a<��a<��a<e�a<�a<��a<}�a<�a<ڌa<��a<^�a<�a<ۋa<��a<t�a<>�a<	�a<܊a<��a<��a<��a<S�a<I�a<)�a<�a<�a<��a<Չa<ʉa<҉a<a<��a<Éa<��a<։a<؉a<�a<�a<�a<0�a<�  �  `�a<`�a<��a<ʊa<֊a<�a<.�a<r�a<��a<�a<�a<P�a<��a<��a<!�a<L�a<��a<��a<c�a<��a<��a<^�a<��a<(�a<f�a<��a<T�a<��a<�a<p�a<��a<N�a<֓a<;�a<��a<"�a<��a<$�a<��a<�a<��a<�a<r�a<�a<��a<יa<^�a<͚a<F�a<Λa<2�a<͜a<�a<��a<�a<��a<�a<s�a<��a<I�a<ߠa<-�a<��a<	�a<k�a<ߢa<-�a<ģa<��a<U�a<��a<�a<d�a<��a<�a<3�a<��a<ʦa<�a<a�a<��a<�a<�a<K�a<t�a<��a< �a<��a<C�a<U�a<��a<��a<ɩa<�a<�a<4�a<8�a<h�a<n�a<��a<��a<��a<�a<٪a<��a<��a<�a<�a<(�a<@�a<�a<7�a<�a</�a<'�a<�a<+�a<	�a<�a<��a<��a<�a<˪a<ªa<��a<��a<i�a<w�a<V�a<�a<�a<ݩa<Ωa<��a<��a<^�a<1�a<	�a<Ĩa<��a<m�a<[�a<�a<�a<§a<��a<\�a<�a<��a<��a<��a<E�a<�a<��a<_�a<3�a<Ԥa<��a<I�a<��a<��a<S�a<�a<��a<i�a<�a<��a<P�a<�a<��a<$�a<˟a<[�a<�a<��a<�a<Νa<9�a<�a<o�a<��a<��a<�a<��a<*�a<ޙa<M�a<�a<r�a<��a<��a<�a<֖a<:�a<̕a<_�a<�a<��a<�a<��a<*�a<Ȓa<_�a<��a<��a<%�a<�a<j�a<�a<��a<i�a<*�a<��a<i�a< �a<��a<p�a<�a<�a<��a<\�a<�a<ދa<��a<s�a<E�a<�a<��a<��a<��a<j�a<T�a<3�a<)�a<%�a<�a<�a<̉a<Չa<ʉa<a<Չa<��a<̉a<ωa<�a<�a<�a<"�a<&�a<�  �  T�a<{�a<��a<��a<��a<"�a<>�a<q�a<��a<׋a<�a<E�a<��a<ٌa<�a<k�a<��a<��a<X�a<��a<�a<`�a<ŏa<(�a<v�a<Ԑa<D�a<��a<�a<��a<�a<K�a<˓a<7�a<��a<�a<��a<�a<��a<�a<z�a<�a<v�a<��a<c�a<ՙa<a�a<�a<J�a<Ǜa<B�a<��a<0�a<��a<&�a<��a<�a<��a<�a<[�a<Рa<<�a<��a<	�a<��a<�a<3�a<��a<�a<^�a<��a<�a<I�a<��a<�a<8�a<~�a<��a<�a<S�a<��a<̧a<�a<=�a<��a<��a<Ԩa<�a<B�a<p�a<��a<��a<ԩa<��a<
�a<3�a<T�a<c�a<��a<��a<��a<Īa<ժa<�a<��a<�a<'�a<�a<�a<'�a<1�a</�a<+�a<,�a<�a< �a<�a<	�a<�a<�a<�a<ުa<��a<��a<��a<��a<��a<b�a<8�a<'�a<�a<�a<ͩa<��a<~�a<[�a<'�a<�a<�a<��a<��a<]�a<�a<��a<ħa<��a<]�a</�a<��a<��a<i�a<5�a<�a<��a<o�a<$�a<Ѥa<��a<E�a<�a<��a<V�a<��a<��a<L�a<�a<��a<T�a<��a<��a<!�a<Οa<v�a<��a<��a<(�a<��a<L�a<ڜa<x�a<��a<��a<)�a<��a<<�a<ϙa<]�a<�a<q�a<�a<��a<�a<��a<G�a<Օa<R�a<�a<q�a<�a<��a<0�a<Òa<V�a<��a<��a<'�a<ΐa<u�a<�a<Ïa<c�a<��a<��a<g�a<�a<��a<l�a<'�a<�a<��a<Z�a<!�a<ًa<��a<r�a<2�a<�a<�a<��a<��a<u�a<n�a<;�a<�a<�a<��a<�a<ىa<щa<��a<ĉa<��a<��a<ˉa<Ήa<܉a<�a<��a<�a<7�a<�  �  A�a<t�a<��a<ˊa<��a<�a<@�a<`�a<��a<׋a<�a<K�a<��a<݌a<�a<p�a<��a<	�a<O�a<��a<�a<N�a<��a<�a<��a<��a<9�a<��a<�a<��a<ޒa<Z�a<��a<=�a<��a<	�a<��a<��a<��a<�a<��a<�a<b�a<�a<S�a<�a<S�a<Ԛa<O�a<��a<W�a<��a<=�a<��a<-�a<��a<��a<��a<ߟa<j�a<��a<N�a<��a<�a<u�a<͢a<g�a<��a<��a<L�a<��a<�a<C�a<��a<ݥa<F�a<r�a<��a<�a<?�a<��a<��a<�a<4�a<u�a<��a<֨a<1�a<'�a<c�a<|�a<��a<�a<�a<�a<'�a<]�a<U�a<��a<��a<��a<Ȫa<Ъa<��a<�a<�a<�a<�a<;�a<�a<+�a<�a<2�a<)�a<�a<�a<
�a<�a<�a<��a<�a<Ӫa<Ūa<��a<��a<��a<|�a<T�a<X�a<7�a<�a<�a<��a<��a<�a<Z�a<,�a<�a<�a<��a<��a<P�a<.�a<�a<ϧa<��a<L�a<(�a<ݦa<Цa<u�a<+�a<�a<��a<~�a<�a<ߤa<��a<K�a<��a<��a<d�a<��a<��a<L�a<�a<��a<@�a<�a<}�a<U�a<��a<b�a<��a<��a<<�a<��a<Y�a<Ӝa<�a<��a<��a<0�a<��a<J�a<��a<o�a<��a<s�a<�a<��a<K�a<��a<:�a<Õa<Q�a<��a<k�a<�a<��a<>�a<��a<W�a< �a<��a<8�a<a<��a<�a<��a<Y�a< �a<֎a<M�a<�a<��a<t�a<8�a<֌a<��a<N�a<)�a<̋a<��a<w�a<6�a<�a<ߊa<Ҋa<��a<u�a<L�a<?�a<<�a<��a<��a<Ӊa<��a<ωa<��a<��a<��a<ȉa<��a<׉a<Չa<�a<��a<�a<@�a<�  �  Q�a<s�a<��a<��a<֊a<�a<J�a<s�a<��a<�a<�a<X�a<��a<Ռa<#�a<f�a<��a<	�a<L�a<��a<�a<e�a<ŏa<�a<p�a<�a<[�a<��a<�a<{�a<�a<R�a<��a<5�a<��a<�a<��a<	�a<y�a<��a<x�a<�a<j�a<��a<l�a<ؙa<U�a<ߚa<]�a<śa<K�a<��a<.�a<��a<!�a<��a<�a<~�a<�a<\�a<ˠa<B�a<��a<�a<��a<עa<4�a<��a<�a<L�a<��a<��a<Q�a<��a<�a<>�a<x�a<��a<�a<B�a<��a<˧a<�a<>�a<q�a<��a<�a< �a<8�a<n�a<��a<��a<ةa<�a<�a</�a<P�a<m�a<~�a<��a<��a<��a<ڪa<�a<��a<�a<�a<�a<�a<2�a<.�a<*�a<%�a<#�a< �a<�a<�a<�a< �a<��a<�a<̪a<Ȫa<��a<��a<��a<{�a<r�a<C�a<�a<�a<��a<ϩa<��a<��a<S�a<:�a<�a<ߨa<��a<��a<W�a</�a<�a<Χa<��a<c�a</�a<�a<��a<v�a<L�a<�a<��a<j�a<!�a<פa<��a<C�a<�a<��a<Z�a<�a<��a<Y�a<�a<��a<H�a<��a<��a<$�a<a<l�a<�a<��a<0�a<��a<J�a<�a<s�a<��a<��a<#�a<��a<=�a<˙a<b�a<�a<��a<�a<��a<�a<��a<I�a<Õa<Q�a<�a<y�a<�a<��a<5�a<��a<U�a<��a<��a<+�a<͐a<n�a<�a<��a<r�a<	�a<��a<]�a<�a<ƍa<n�a<,�a<Ԍa<��a<V�a<�a<�a<��a<v�a<I�a<	�a<�a<a<��a<��a<W�a</�a<�a<�a<��a<�a<Ӊa<ȉa<a<��a<a<ĉa<ŉa<҉a<މa<��a< �a<�a</�a<�  �  R�a<`�a<��a<��a<��a<#�a<0�a<��a<��a<�a<�a<\�a<��a<׌a<#�a<e�a<͍a<�a<`�a<��a<��a<l�a<��a<:�a<��a<ېa<@�a<��a<�a<m�a<��a<J�a<˓a<6�a<��a<�a<}�a<�a<o�a<	�a<k�a<�a<l�a<ܘa<o�a<͙a<��a<ߚa<O�a<՛a<C�a<Ӝa<+�a<��a<�a<��a<�a<y�a<�a<Y�a<�a<A�a<��a<�a<x�a<�a<+�a<��a<�a<M�a<��a<�a<_�a<��a<�a<*�a<|�a<��a<
�a<U�a<y�a<ܧa<��a<D�a<k�a<��a<ݨa<�a<]�a<W�a<��a<��a<�a<�a<�a<M�a<M�a<p�a<��a<��a<��a<ªa<�a<۪a<�a<��a<!�a<5�a<�a<1�a<�a<(�a<�a<&�a<*�a<�a<�a<�a<�a<֪a<�a<Ӫa<ͪa<��a<��a<��a<i�a<e�a<7�a<>�a< �a<ߩa<۩a<��a<��a<]�a<=�a<�a<�a<��a<��a<r�a<-�a<�a<ҧa<��a<j�a<�a<�a<��a<p�a<1�a<�a<��a<\�a<4�a<Ϥa<��a<D�a<�a<��a<@�a<�a<��a<e�a<��a<��a<J�a<�a<��a<�a<�a<l�a<��a<��a<)�a<ӝa<G�a<��a<q�a<�a<��a<�a<ɚa<:�a<�a<b�a<��a<z�a<�a<��a<�a<��a</�a<ŕa<\�a<ڔa<��a<�a<��a<"�a<��a<Q�a<��a<��a<�a<ސa<^�a<�a<��a<V�a<�a<��a<��a<�a<ča<o�a<4�a<�a<��a<t�a<�a<�a<��a<|�a<Q�a<�a<��a<��a<��a<n�a<i�a<W�a<�a<�a<�a<�a<ˉa<ˉa<͉a<��a<��a<��a<ˉa<��a<ډa<�a<�a<�a<&�a<�  �  E�a<y�a<��a<Ȋa<�a<��a<=�a<y�a<��a<݋a<$�a<T�a<��a<ތa<�a<j�a<��a<�a<d�a<��a<�a<j�a<��a<�a<��a<�a<?�a<��a<�a<u�a<ޒa<J�a<Óa<6�a<��a<�a<��a<�a<�a<��a<l�a<��a<k�a<�a<n�a<�a<O�a<Ěa<P�a<˛a<A�a<a<6�a<��a<"�a<��a<�a<��a<�a<a�a<Ԡa<7�a<��a<�a<e�a<͢a<J�a<��a<��a<V�a<��a<�a<I�a<��a<�a<3�a<x�a<��a<�a<L�a<��a<ŧa<��a<>�a<��a<��a<�a<�a<(�a<X�a<��a<��a<өa<��a<�a<.�a<O�a<e�a<��a<��a<��a<Ѫa<ުa<�a<��a<�a<��a<�a<+�a<+�a<*�a<�a<.�a<�a<�a<�a<�a<�a<��a<�a<�a<Ѫa<��a<��a<��a<��a<��a<c�a<T�a</�a<��a<�a<թa<��a<��a<k�a<5�a<�a<�a<��a<��a<T�a<-�a<�a<ŧa<��a<h�a<�a<צa<��a<��a<0�a<��a<��a<c�a<�a<Фa<��a<D�a<�a<��a<R�a<�a<��a<Q�a<��a<��a<J�a<�a<��a<:�a<��a<Q�a<��a<��a<&�a<Ýa<R�a<�a<t�a<�a<��a<%�a<��a<A�a<ԙa<X�a<�a<y�a<��a<��a<-�a<��a<>�a<Εa<_�a<ݔa<q�a<�a<��a<+�a<��a<V�a<�a<��a<$�a<ǐa<f�a<�a<Ïa<]�a<�a<��a<N�a<�a<ča<u�a<'�a<�a<��a<U�a<�a<ۋa<��a<m�a<A�a<�a<�a<��a<��a<y�a<B�a<8�a<,�a<�a<��a<ىa<܉a<a<��a<��a<a<��a<a<ȉa<��a<�a<��a<�a<4�a<�  �  <�a<}�a<z�a<��a<��a<�a<a�a<e�a<��a<׋a<�a<a�a<��a<�a<+�a<y�a<��a<�a<S�a<��a<�a<U�a<ޏa<�a<�a<ِa<5�a<��a<��a<��a<̒a<T�a<��a<(�a<��a<�a<��a<�a<z�a<�a<u�a<�a<e�a<��a<C�a<�a<R�a<��a<d�a<˛a<P�a<��a<D�a<��a<*�a<��a<�a<��a<�a<r�a<àa<E�a<��a<�a<��a<Ңa<I�a<~�a<��a<L�a<��a<�a<6�a<��a<ӥa<3�a<p�a<��a<��a<6�a<��a<��a<�a</�a<z�a<��a<Ϩa<�a<5�a<��a<��a<éa<թa<�a<+�a<,�a<]�a<w�a<��a<��a<��a<ɪa<Ҫa<��a<�a<%�a<$�a<�a<)�a<�a<7�a<�a</�a<�a<�a<�a<�a<�a<�a<�a<تa<Ǫa<êa<��a<��a<{�a<��a<G�a<L�a<'�a<�a<�a<��a<��a<�a<]�a<C�a<
�a<�a<¨a<��a<R�a<?�a<��a<ŧa<��a<S�a<H�a<�a<��a<n�a<'�a<��a<��a<x�a<�a<٤a<y�a<7�a<�a<��a<S�a<�a<��a<D�a<��a<��a<C�a<��a<l�a<:�a<��a<��a<�a<��a<5�a<��a<`�a<�a<|�a<�a<��a<*�a<��a<R�a<Ùa<f�a<�a<��a<'�a<��a<-�a<��a<@�a<ĕa<M�a<�a<^�a<�a<��a<+�a<��a<T�a<�a<z�a</�a<��a<{�a< �a<��a<W�a<��a<��a<[�a<1�a<��a<��a<(�a<ٌa<��a<S�a<)�a<�a<��a<t�a<N�a<�a<�a<Њa<��a<��a<k�a<3�a<*�a<�a<�a<Չa<݉a<��a<��a<��a<��a<��a<��a<͉a<͉a<ۉa<��a<�a<=�a<�  �  M�a<{�a<��a<Êa<�a<�a<(�a<s�a<��a<�a<�a<\�a<��a<͌a<+�a<[�a<ƍa<�a<^�a<��a<�a<V�a<��a<!�a<~�a<�a<K�a<��a<�a<z�a<�a<S�a<��a<3�a<��a<�a<��a<�a<~�a<��a<t�a<�a<s�a<�a<i�a<�a<`�a<Ԛa<>�a<؛a<D�a<̜a<1�a<��a<"�a<��a<�a<v�a<��a<]�a<ߠa<A�a<��a<��a<q�a<�a<@�a<��a<��a<[�a<��a<�a<I�a<��a<�a<,�a<~�a<��a<�a<E�a<��a<��a<�a<=�a<��a<��a<�a<�a<>�a<W�a<{�a<��a<�a<�a<�a<D�a<B�a<y�a<}�a<��a<��a<��a<�a<�a<��a<�a<�a<�a<+�a<)�a<4�a<&�a<"�a<�a<�a<�a<�a<��a<��a<�a<ުa<Ϫa<Ǫa<��a<��a<��a<��a<f�a<P�a<*�a<�a<שa<ϩa<��a<��a<Z�a<>�a<�a<רa<¨a<{�a<k�a<,�a< �a<٧a<��a<T�a<�a<�a<��a<��a<<�a<��a<��a<i�a<�a<٤a<��a<A�a<�a<��a<H�a<��a<��a<V�a<��a<��a<Q�a<��a<��a<2�a<Οa<a�a<�a<��a<)�a<͝a<M�a<�a<t�a<�a<��a<�a<��a<=�a<ޙa<a�a<��a<g�a< �a<��a<$�a<��a<B�a<ӕa<V�a<�a<q�a<�a<��a<$�a<a<T�a<�a<��a<-�a<a<o�a<�a<��a<f�a<�a<��a<c�a<�a<��a<}�a<6�a<�a<��a<k�a<�a<�a<��a<~�a<R�a<�a<��a<��a<��a<b�a<]�a<9�a<+�a<�a<�a<�a<Љa<a<��a<��a<��a<��a<ĉa<��a<Ӊa<�a<��a<�a<-�a<�  �  J�a<[�a<��a<��a<݊a<$�a<=�a<��a<��a<�a<�a<T�a<��a<Ҍa<>�a<Z�a<�a<��a<e�a<��a<��a<��a<Ïa<%�a<e�a<ސa<7�a<��a<�a<^�a<�a<F�a<��a<*�a<��a<+�a<n�a<�a<s�a<��a<f�a<�a<d�a<Ƙa<y�a<Йa<f�a<ݚa<a�a<��a<%�a<ۜa<#�a<ĝa<"�a<��a<%�a<}�a<�a<N�a<�a<�a<ġa<+�a<}�a<�a<*�a<��a<٣a<I�a<��a<�a<M�a<��a<�a<�a<��a<��a<��a<C�a<��a<ϧa<�a<7�a<m�a<��a<�a<��a<E�a<i�a<��a<��a<˩a<�a<��a<_�a<B�a<��a<��a<��a<��a<��a<�a<Ūa<:�a<�a< �a<�a<�a<2�a<�a<�a< �a<'�a<�a<�a<�a<�a<�a<ܪa<�a<Ȫa<��a<��a<��a<��a<d�a<f�a<>�a<$�a<!�a<�a<�a<��a<��a<_�a<6�a<*�a<ܨa<֨a<z�a<��a<�a<�a<ʧa<��a<��a<,�a<��a<��a<s�a<(�a<�a<��a<M�a<-�a<̤a<}�a<8�a<�a<��a<1�a< �a<��a<W�a<�a<��a<C�a<ˠa<��a<�a<ӟa<j�a<�a<��a<
�a<ܝa<?�a<��a<t�a<�a<��a<"�a<Ӛa<.�a<�a<@�a<�a<��a<�a<��a<�a<��a<�a<��a<M�a<Ӕa<u�a<��a<��a<�a<ɒa<M�a<�a<��a< �a<ѐa<Q�a<	�a<��a<H�a<�a<��a<j�a<�a<�a<r�a<�a<��a<��a<��a<�a<�a<��a<��a<K�a<�a< �a<��a<܊a<z�a<g�a<6�a<�a<�a<ډa<ډa<Ήa<̉a<��a<��a<��a<��a<߉a<��a<׉a<܉a<��a<�a<�a<�  �  M�a<{�a<��a<Êa<�a<�a<(�a<s�a<��a<�a<�a<\�a<��a<͌a<+�a<[�a<ƍa<�a<^�a<��a<�a<V�a<��a<!�a<~�a<�a<K�a<��a<�a<z�a<�a<S�a<��a<3�a<��a<�a<��a<�a<~�a<��a<t�a<�a<s�a<�a<i�a<�a<`�a<Ԛa<>�a<؛a<D�a<̜a<1�a<��a<"�a<��a<�a<v�a<��a<]�a<ߠa<A�a<��a<��a<q�a<�a<@�a<��a<��a<[�a<��a<�a<I�a<��a<�a<,�a<~�a<��a<�a<E�a<��a<��a<�a<=�a<��a<��a<�a<�a<>�a<W�a<{�a<��a<�a<�a<�a<D�a<B�a<y�a<}�a<��a<��a<��a<�a<�a<��a<�a<�a<�a<+�a<)�a<4�a<&�a<"�a<�a<�a<�a<�a<��a<��a<�a<ުa<Ϫa<Ǫa<��a<��a<��a<��a<f�a<P�a<*�a<�a<שa<ϩa<��a<��a<Z�a<>�a<�a<רa<¨a<{�a<k�a<,�a< �a<٧a<��a<T�a<�a<�a<��a<��a<<�a<��a<��a<i�a<�a<٤a<��a<A�a<�a<��a<H�a<��a<��a<V�a<��a<��a<Q�a<��a<��a<2�a<Οa<a�a<�a<��a<)�a<͝a<M�a<�a<t�a<�a<��a<�a<��a<=�a<ޙa<a�a<��a<g�a< �a<��a<$�a<��a<B�a<ӕa<V�a<�a<q�a<�a<��a<$�a<a<T�a<�a<��a<-�a<a<o�a<�a<��a<f�a<�a<��a<c�a<�a<��a<}�a<6�a<�a<��a<k�a<�a<�a<��a<~�a<R�a<�a<��a<��a<��a<b�a<]�a<9�a<+�a<�a<�a<�a<Љa<a<��a<��a<��a<��a<ĉa<��a<Ӊa<�a<��a<�a<-�a<�  �  <�a<}�a<z�a<��a<��a<�a<a�a<e�a<��a<׋a<�a<a�a<��a<�a<+�a<y�a<��a<�a<S�a<��a<�a<U�a<ޏa<�a<�a<ِa<5�a<��a<��a<��a<̒a<T�a<��a<(�a<��a<�a<��a<�a<z�a<�a<u�a<�a<e�a<��a<C�a<�a<R�a<��a<d�a<˛a<P�a<��a<D�a<��a<*�a<��a<�a<��a<�a<r�a<àa<E�a<��a<�a<��a<Ңa<I�a<~�a<��a<L�a<��a<�a<6�a<��a<ӥa<3�a<p�a<��a<��a<6�a<��a<��a<�a</�a<z�a<��a<Ϩa<�a<5�a<��a<��a<éa<թa<�a<+�a<,�a<]�a<w�a<��a<��a<��a<ɪa<Ҫa<��a<�a<%�a<$�a<�a<)�a<�a<7�a<�a</�a<�a<�a<�a<�a<�a<�a<�a<تa<Ǫa<êa<��a<��a<{�a<��a<G�a<L�a<'�a<�a<�a<��a<��a<�a<]�a<C�a<
�a<�a<¨a<��a<R�a<?�a<��a<ŧa<��a<S�a<H�a<�a<��a<n�a<'�a<��a<��a<x�a<�a<٤a<y�a<7�a<�a<��a<S�a<�a<��a<D�a<��a<��a<C�a<��a<l�a<:�a<��a<��a<�a<��a<5�a<��a<`�a<�a<|�a<�a<��a<*�a<��a<R�a<Ùa<f�a<�a<��a<'�a<��a<-�a<��a<@�a<ĕa<M�a<�a<^�a<�a<��a<+�a<��a<T�a<�a<z�a</�a<��a<{�a< �a<��a<W�a<��a<��a<[�a<1�a<��a<��a<(�a<ٌa<��a<S�a<)�a<�a<��a<t�a<N�a<�a<�a<Њa<��a<��a<k�a<3�a<*�a<�a<�a<Չa<݉a<��a<��a<��a<��a<��a<��a<͉a<͉a<ۉa<��a<�a<=�a<�  �  E�a<y�a<��a<Ȋa<�a<��a<=�a<y�a<��a<݋a<$�a<T�a<��a<ތa<�a<j�a<��a<�a<d�a<��a<�a<j�a<��a<�a<��a<�a<?�a<��a<�a<u�a<ޒa<J�a<Óa<6�a<��a<�a<��a<�a<�a<��a<l�a<��a<k�a<�a<n�a<�a<O�a<Ěa<P�a<˛a<A�a<a<6�a<��a<"�a<��a<�a<��a<�a<a�a<Ԡa<7�a<��a<�a<e�a<͢a<J�a<��a<��a<V�a<��a<�a<I�a<��a<�a<3�a<x�a<��a<�a<L�a<��a<ŧa<��a<>�a<��a<��a<�a<�a<(�a<X�a<��a<��a<өa<��a<�a<.�a<O�a<e�a<��a<��a<��a<Ѫa<ުa<�a<��a<�a<��a<�a<+�a<+�a<*�a<�a<.�a<�a<�a<�a<�a<�a<��a<�a<�a<Ѫa<��a<��a<��a<��a<��a<c�a<T�a</�a<��a<�a<թa<��a<��a<k�a<5�a<�a<�a<��a<��a<T�a<-�a<�a<ŧa<��a<h�a<�a<צa<��a<��a<0�a<��a<��a<c�a<�a<Фa<��a<D�a<�a<��a<R�a<�a<��a<Q�a<��a<��a<J�a<�a<��a<:�a<��a<Q�a<��a<��a<&�a<Ýa<R�a<�a<t�a<�a<��a<%�a<��a<A�a<ԙa<X�a<�a<y�a<��a<��a<-�a<��a<>�a<Εa<_�a<ݔa<q�a<�a<��a<+�a<��a<V�a<�a<��a<$�a<ǐa<f�a<�a<Ïa<]�a<�a<��a<N�a<�a<ča<u�a<'�a<�a<��a<U�a<�a<ۋa<��a<m�a<A�a<�a<�a<��a<��a<y�a<B�a<8�a<,�a<�a<��a<ىa<܉a<a<��a<��a<a<��a<a<ȉa<��a<�a<��a<�a<4�a<�  �  R�a<`�a<��a<��a<��a<#�a<0�a<��a<��a<�a<�a<\�a<��a<׌a<#�a<e�a<͍a<�a<`�a<��a<��a<l�a<��a<:�a<��a<ېa<@�a<��a<�a<m�a<��a<J�a<˓a<6�a<��a<�a<}�a<�a<o�a<	�a<k�a<�a<l�a<ܘa<o�a<͙a<��a<ߚa<O�a<՛a<C�a<Ӝa<+�a<��a<�a<��a<�a<y�a<�a<Y�a<�a<A�a<��a<�a<x�a<�a<+�a<��a<�a<M�a<��a<�a<_�a<��a<�a<*�a<|�a<��a<
�a<U�a<y�a<ܧa<��a<D�a<k�a<��a<ݨa<�a<]�a<W�a<��a<��a<�a<�a<�a<M�a<M�a<p�a<��a<��a<��a<ªa<�a<۪a<�a<��a<!�a<5�a<�a<1�a<�a<(�a<�a<&�a<*�a<�a<�a<�a<�a<֪a<�a<Ӫa<ͪa<��a<��a<��a<i�a<e�a<7�a<>�a< �a<ߩa<۩a<��a<��a<]�a<=�a<�a<�a<��a<��a<r�a<-�a<�a<ҧa<��a<j�a<�a<�a<��a<p�a<1�a<�a<��a<\�a<4�a<Ϥa<��a<D�a<�a<��a<@�a<�a<��a<e�a<��a<��a<J�a<�a<��a<�a<�a<l�a<��a<��a<)�a<ӝa<G�a<��a<q�a<�a<��a<�a<ɚa<:�a<�a<b�a<��a<z�a<�a<��a<�a<��a</�a<ŕa<\�a<ڔa<��a<�a<��a<"�a<��a<Q�a<��a<��a<�a<ސa<^�a<�a<��a<V�a<�a<��a<��a<�a<ča<o�a<4�a<�a<��a<t�a<�a<�a<��a<|�a<Q�a<�a<��a<��a<��a<n�a<i�a<W�a<�a<�a<�a<�a<ˉa<ˉa<͉a<��a<��a<��a<ˉa<��a<ډa<�a<�a<�a<&�a<�  �  Q�a<s�a<��a<��a<֊a<�a<J�a<s�a<��a<�a<�a<X�a<��a<Ռa<#�a<f�a<��a<	�a<L�a<��a<�a<e�a<ŏa<�a<p�a<�a<[�a<��a<�a<{�a<�a<R�a<��a<5�a<��a<�a<��a<	�a<y�a<��a<x�a<�a<j�a<��a<l�a<ؙa<U�a<ߚa<]�a<śa<K�a<��a<.�a<��a<!�a<��a<�a<~�a<�a<\�a<ˠa<B�a<��a<�a<��a<עa<4�a<��a<�a<L�a<��a<��a<Q�a<��a<�a<>�a<x�a<��a<�a<B�a<��a<˧a<�a<>�a<q�a<��a<�a< �a<8�a<n�a<��a<��a<ةa<�a<�a</�a<P�a<m�a<~�a<��a<��a<��a<ڪa<�a<��a<�a<�a<�a<�a<2�a<.�a<*�a<%�a<#�a< �a<�a<�a<�a< �a<��a<�a<̪a<Ȫa<��a<��a<��a<{�a<r�a<C�a<�a<�a<��a<ϩa<��a<��a<S�a<:�a<�a<ߨa<��a<��a<W�a</�a<�a<Χa<��a<c�a</�a<�a<��a<v�a<L�a<�a<��a<j�a<!�a<פa<��a<C�a<�a<��a<Z�a<�a<��a<Y�a<�a<��a<H�a<��a<��a<$�a<a<l�a<�a<��a<0�a<��a<J�a<�a<s�a<��a<��a<#�a<��a<=�a<˙a<b�a<�a<��a<�a<��a<�a<��a<I�a<Õa<Q�a<�a<y�a<�a<��a<5�a<��a<U�a<��a<��a<+�a<͐a<n�a<�a<��a<r�a<	�a<��a<]�a<�a<ƍa<n�a<,�a<Ԍa<��a<V�a<�a<�a<��a<v�a<I�a<	�a<�a<a<��a<��a<W�a</�a<�a<�a<��a<�a<Ӊa<ȉa<a<��a<a<ĉa<ŉa<҉a<މa<��a< �a<�a</�a<�  �  A�a<t�a<��a<ˊa<��a<�a<@�a<`�a<��a<׋a<�a<K�a<��a<݌a<�a<p�a<��a<	�a<O�a<��a<�a<N�a<��a<�a<��a<��a<9�a<��a<�a<��a<ޒa<Z�a<��a<=�a<��a<	�a<��a<��a<��a<�a<��a<�a<b�a<�a<S�a<�a<S�a<Ԛa<O�a<��a<W�a<��a<=�a<��a<-�a<��a<��a<��a<ߟa<j�a<��a<N�a<��a<�a<u�a<͢a<g�a<��a<��a<L�a<��a<�a<C�a<��a<ݥa<F�a<r�a<��a<�a<?�a<��a<��a<�a<4�a<u�a<��a<֨a<1�a<'�a<c�a<|�a<��a<�a<�a<�a<'�a<]�a<U�a<��a<��a<��a<Ȫa<Ъa<��a<�a<�a<�a<�a<;�a<�a<+�a<�a<2�a<)�a<�a<�a<
�a<�a<�a<��a<�a<Ӫa<Ūa<��a<��a<��a<|�a<T�a<X�a<7�a<�a<�a<��a<��a<�a<Z�a<,�a<�a<�a<��a<��a<P�a<.�a<�a<ϧa<��a<L�a<(�a<ݦa<Цa<u�a<+�a<�a<��a<~�a<�a<ߤa<��a<K�a<��a<��a<d�a<��a<��a<L�a<�a<��a<@�a<�a<}�a<U�a<��a<b�a<��a<��a<<�a<��a<Y�a<Ӝa<�a<��a<��a<0�a<��a<J�a<��a<o�a<��a<s�a<�a<��a<K�a<��a<:�a<Õa<Q�a<��a<k�a<�a<��a<>�a<��a<W�a< �a<��a<8�a<a<��a<�a<��a<Y�a< �a<֎a<M�a<�a<��a<t�a<8�a<֌a<��a<N�a<)�a<̋a<��a<w�a<6�a<�a<ߊa<Ҋa<��a<u�a<L�a<?�a<<�a<��a<��a<Ӊa<��a<ωa<��a<��a<��a<ȉa<��a<׉a<Չa<�a<��a<�a<@�a<�  �  T�a<{�a<��a<��a<��a<"�a<>�a<q�a<��a<׋a<�a<E�a<��a<ٌa<�a<k�a<��a<��a<X�a<��a<�a<`�a<ŏa<(�a<v�a<Ԑa<D�a<��a<�a<��a<�a<K�a<˓a<7�a<��a<�a<��a<�a<��a<�a<z�a<�a<v�a<��a<c�a<ՙa<a�a<�a<J�a<Ǜa<B�a<��a<0�a<��a<&�a<��a<�a<��a<�a<[�a<Рa<<�a<��a<	�a<��a<�a<3�a<��a<�a<^�a<��a<�a<I�a<��a<�a<8�a<~�a<��a<�a<S�a<��a<̧a<�a<=�a<��a<��a<Ԩa<�a<B�a<p�a<��a<��a<ԩa<��a<
�a<3�a<T�a<c�a<��a<��a<��a<Īa<ժa<�a<��a<�a<'�a<�a<�a<'�a<1�a</�a<+�a<,�a<�a< �a<�a<	�a<�a<�a<�a<ުa<��a<��a<��a<��a<��a<b�a<8�a<'�a<�a<�a<ͩa<��a<~�a<[�a<'�a<�a<�a<��a<��a<]�a<�a<��a<ħa<��a<]�a</�a<��a<��a<i�a<5�a<�a<��a<o�a<$�a<Ѥa<��a<E�a<�a<��a<V�a<��a<��a<L�a<�a<��a<T�a<��a<��a<!�a<Οa<v�a<��a<��a<(�a<��a<L�a<ڜa<x�a<��a<��a<)�a<��a<<�a<ϙa<]�a<�a<q�a<�a<��a<�a<��a<G�a<Օa<R�a<�a<q�a<�a<��a<0�a<Òa<V�a<��a<��a<'�a<ΐa<u�a<�a<Ïa<c�a<��a<��a<g�a<�a<��a<l�a<'�a<�a<��a<Z�a<!�a<ًa<��a<r�a<2�a<�a<�a<��a<��a<u�a<n�a<;�a<�a<�a<��a<�a<ىa<щa<��a<ĉa<��a<��a<ˉa<Ήa<܉a<�a<��a<�a<7�a<�  �  `�a<`�a<��a<ʊa<֊a<�a<.�a<r�a<��a<�a<�a<P�a<��a<��a<!�a<L�a<��a<��a<c�a<��a<��a<^�a<��a<(�a<f�a<��a<T�a<��a<�a<p�a<��a<N�a<֓a<;�a<��a<"�a<��a<$�a<��a<�a<��a<�a<r�a<�a<��a<יa<^�a<͚a<F�a<Λa<2�a<͜a<�a<��a<�a<��a<�a<s�a<��a<I�a<ߠa<-�a<��a<	�a<k�a<ߢa<-�a<ģa<��a<U�a<��a<�a<d�a<��a<�a<3�a<��a<ʦa<�a<a�a<��a<�a<�a<K�a<t�a<��a< �a<��a<C�a<U�a<��a<��a<ɩa<�a<�a<4�a<8�a<h�a<n�a<��a<��a<��a<�a<٪a<��a<��a<�a<�a<(�a<@�a<�a<7�a<�a</�a<'�a<�a<+�a<	�a<�a<��a<��a<�a<˪a<ªa<��a<��a<i�a<w�a<V�a<�a<�a<ݩa<Ωa<��a<��a<^�a<1�a<	�a<Ĩa<��a<m�a<[�a<�a<�a<§a<��a<\�a<�a<��a<��a<��a<E�a<�a<��a<_�a<3�a<Ԥa<��a<I�a<��a<��a<S�a<�a<��a<i�a<�a<��a<P�a<�a<��a<$�a<˟a<[�a<�a<��a<�a<Νa<9�a<�a<o�a<��a<��a<�a<��a<*�a<ޙa<M�a<�a<r�a<��a<��a<�a<֖a<:�a<̕a<_�a<�a<��a<�a<��a<*�a<Ȓa<_�a<��a<��a<%�a<�a<j�a<�a<��a<i�a<*�a<��a<i�a< �a<��a<p�a<�a<�a<��a<\�a<�a<ދa<��a<s�a<E�a<�a<��a<��a<��a<j�a<T�a<3�a<)�a<%�a<�a<�a<̉a<Չa<ʉa<a<Չa<��a<̉a<ωa<�a<�a<�a<"�a<&�a<�  �  \�a<m�a<{�a<��a<�a<�a<F�a<d�a<��a<Ћa<�a<L�a<��a<Ќa<�a<b�a<��a<��a<P�a<��a<�a<V�a<��a<!�a<��a<ؐa<-�a<��a<�a<y�a<�a<_�a<ēa<0�a<��a<�a<��a<�a<��a<�a<u�a<��a<r�a<ݘa<V�a<�a<g�a<ؚa<\�a<̛a<;�a<��a<*�a<��a<�a<��a<�a<w�a<�a<[�a<Ƞa<2�a<��a<�a<y�a<�a<J�a<��a<�a<T�a<��a<��a<U�a<��a<�a<9�a<��a<Цa<
�a<N�a<��a<ӧa<�a<B�a<x�a<��a<Ҩa<�a<@�a<b�a<��a<��a<ɩa<�a<�a<7�a<L�a<d�a<~�a<��a<��a<��a<ͪa<�a<�a<�a<�a<(�a<(�a<�a<#�a<5�a<'�a<$�a<0�a<�a<�a<�a<��a<��a<�a<۪a<٪a<��a<��a<��a<v�a<H�a<M�a<9�a<�a<��a<��a<��a<w�a<S�a<.�a<�a<٨a<��a<��a<_�a<$�a<�a<��a<��a<T�a<%�a<�a<��a<m�a<�a<��a<��a<h�a<+�a<�a<��a<?�a< �a<��a<U�a<��a<��a<`�a<��a<��a<P�a<�a<��a<8�a<ԟa<e�a<�a<��a< �a<��a<F�a<�a<l�a<��a<��a<�a<��a<;�a<Ǚa<S�a<�a<~�a<	�a<��a<.�a<��a<,�a<̕a<Z�a<�a<|�a<
�a<��a<1�a<˒a<f�a<��a<��a<3�a<Րa<k�a<�a<��a<I�a<��a<��a<e�a<�a<��a<}�a<�a<ڌa<��a<^�a<�a<ۋa<��a<t�a<>�a<	�a<܊a<��a<��a<��a<S�a<I�a<)�a<�a<�a<��a<Չa<ʉa<҉a<a<��a<Éa<��a<։a<؉a<�a<�a<�a<0�a<�  �  G�a<��a<��a<��a<�a<��a<H�a<Z�a<��a<ċa<�a<A�a<��a<ӌa<�a<d�a<��a<��a<K�a<��a<
�a<R�a<ˏa<��a<��a<Րa<Z�a<Ǒa<�a<��a<�a<\�a<Гa<8�a<��a<)�a<��a<�a<��a<�a<y�a<�a<i�a<�a<_�a<�a<I�a<Ԛa<R�a<��a<O�a<��a<4�a<��a<�a<��a<��a<w�a<֟a<_�a<��a<B�a<��a<�a<y�a<��a<H�a<��a<�a<X�a<��a<�a<E�a<��a<�a<@�a<��a<Цa<�a<V�a<��a<ça<�a<<�a<��a<ƨa<Өa<�a<�a<o�a<��a<��a<ϩa<�a<�a<�a<L�a<P�a<~�a<��a<��a<êa<��a<��a<�a<�a< �a<�a<"�a<)�a<K�a<�a<?�a<!�a<�a<.�a<�a<�a<�a<�a<�a<�a<ɪa<��a<��a<��a<��a<j�a<E�a<-�a<��a<��a<��a<��a<l�a<X�a<#�a<��a<ݨa<��a<��a<F�a<�a<�a<��a<��a<P�a<4�a<˦a<��a<j�a<K�a<�a<��a<z�a<�a<�a<��a<F�a<�a<��a<`�a<��a<Ģa<O�a<�a<��a<G�a<�a<��a<3�a<��a<a�a<��a<��a<4�a<��a<Q�a<ʜa<h�a<��a<��a<�a<��a<?�a<��a<c�a<ޘa<t�a<�a<x�a<,�a<��a<^�a<Еa<c�a<�a<l�a<�a<��a<8�a<Вa<f�a<��a<��a<<�a<Őa<|�a<�a<͏a<y�a<��a<��a<;�a<�a<��a<p�a<#�a<Ќa<��a<D�a<�a<ǋa<��a<g�a<,�a<�a<͊a<͊a<��a<�a<G�a<8�a<#�a<�a<�a<ډa<�a<ǉa<��a<҉a<��a<щa<҉a<މa<ډa<��a<�a<�a<I�a<�  �  R�a<[�a<��a<��a<�a<�a<G�a<l�a<��a<Ջa<�a<H�a<��a<ǌa<�a<X�a<��a<��a<U�a<��a< �a<_�a<ɏa<�a<��a<ސa<J�a<��a<�a<{�a<��a<Q�a<֓a<>�a<��a<,�a<��a<�a<��a<�a<��a<��a<\�a<ޘa<i�a<�a<h�a<ߚa<\�a<ța<D�a<��a<3�a<��a<�a<��a<�a<t�a<�a<^�a<Ơa<>�a<��a<�a<~�a<�a<?�a<��a<�a<A�a<��a<�a<a�a<��a<��a<.�a<��a<ʦa<�a<_�a<��a<ܧa<�a<L�a<c�a<��a<ߨa<�a<=�a<k�a<��a<��a<ϩa<��a<�a</�a<A�a<h�a<u�a<��a<��a<Īa<Ҫa<�a<��a<�a<�a<%�a<#�a<,�a<�a<#�a<0�a<7�a<%�a<�a<$�a<��a<�a<�a<��a<ߪa<Ȫa<ɪa<��a<��a<d�a<h�a<G�a<5�a<�a<��a<ǩa<��a<}�a<Z�a<*�a<�a<Ѩa<��a<y�a<S�a<$�a<��a<��a<��a<\�a<2�a<�a<��a<s�a<;�a<ޥa<��a<i�a<6�a<פa<��a<L�a<�a<��a<I�a<�a<��a<g�a<�a<��a<:�a<�a<��a<.�a<֟a<m�a<�a<��a<)�a<��a<O�a<ڜa<l�a<��a<��a<�a<��a<>�a<ƙa<_�a<�a<��a<�a<��a<#�a<��a<5�a<��a<i�a<�a<��a<�a<��a<&�a<ђa<_�a<��a<��a<,�a<ݐa<n�a<�a<��a<_�a<	�a<��a<b�a<�a<��a<o�a<"�a<ߌa<��a<V�a<�a<ދa<��a<q�a<6�a<�a<�a<��a<��a<�a<_�a<G�a<#�a<�a<�a<މa<މa<܉a<ǉa<a<Ήa<��a<҉a<ĉa<�a<�a< �a<*�a<6�a<�  �  ��a<x�a<ȉa<׉a<�a<�a<;�a<��a<��a<�a<�a<^�a<��a<ʋa<@�a<V�a<ٌa<��a<W�a<��a<"�a<��a<Îa<1�a<��a<�a<~�a<Аa<c�a<�a<3�a<��a<��a<a�a<Ǔa<P�a<��a<U�a<��a<_�a<��a<(�a<Зa<�a<Ęa<�a<��a<��a<��a<�a<��a<��a<I�a<�a<R�a<ٝa<X�a<��a<C�a<~�a<�a<��a<��a<Z�a<��a<*�a<�a<�a<P�a<ˣa<�a<?�a<դa<�a<c�a<~�a<֥a<�a<]�a<��a<�a<L�a<A�a<��a<ݧa<�a<Q�a<C�a<��a<��a<ިa<�a<�a<3�a<;�a<��a<t�a<ȩa<��a<�a<��a<�a<#�a<3�a<U�a<C�a<N�a<]�a<x�a<��a<i�a<��a<c�a<z�a<��a<d�a<y�a<D�a<h�a<7�a<D�a<(�a<0�a<�a<ԩa<�a<��a<ϩa<��a<i�a<I�a<#�a<)�a<�a<Ǩa<��a<v�a<[�a<
�a<�a<��a<��a<R�a<,�a<�a<�a<��a<]�a<3�a<�a<ܥa<��a<F�a<,�a<��a<��a<2�a<�a<��a<:�a<��a<��a<o�a<�a<١a<@�a<��a<Ơa<4�a<�a<q�a<
�a<��a<;�a<ߝa<l�a<�a<h�a<'�a<��a<A�a<ٚa<D�a<��a<P�a<�a<��a<'�a<��a<&�a<Ɩa<E�a<�a<q�a<�a<��a<�a<ԓa<*�a<�a<I�a<�a<{�a<�a<ΐa<T�a<�a<u�a<X�a<�a<��a<E�a<��a<z�a<�a<ٌa<��a<5�a<�a<��a<��a<�a<�a<��a<��a<R�a<��a<��a<Ήa<��a<y�a<Y�a<B�a<<�a<B�a<��a<+�a<Ԉa<�a<��a<ˈa<�a<��a<�a<Ոa<��a< �a<,�a<>�a<'�a<�  �  a�a<p�a<��a<Ɖa<	�a<.�a<\�a<}�a<��a<�a<-�a<Z�a<��a<ыa<�a<j�a<Ȍa<�a<x�a<��a<�a<x�a<�a<E�a<��a<��a<_�a<��a<7�a<��a<�a<w�a<��a<a�a<�a<f�a<��a<C�a<��a<2�a<��a<'�a<��a<�a<��a<�a<��a<#�a<��a<�a<|�a<��a<o�a<�a<Z�a<��a<4�a<��a<1�a<��a<�a<��a<�a<h�a<ۡa<<�a<��a<�a<>�a<��a<��a<W�a<��a<�a<Q�a<��a<�a<3�a<d�a<��a<ߦa<(�a<c�a<��a<��a<��a<+�a<f�a<��a<Ǩa<ܨa<��a<�a<P�a<V�a<��a<��a<��a<��a<�a<�a<�a<!�a<+�a<A�a<_�a<j�a<y�a<l�a<t�a<f�a<u�a<z�a<z�a<u�a<j�a<j�a<[�a<q�a<K�a<9�a<,�a<�a<�a<��a<ܩa<��a<��a<��a<��a<e�a<D�a<�a<�a<ɨa<��a<s�a<Q�a<�a<�a<��a<��a<f�a<M�a<
�a<զa<��a<��a<F�a<�a<��a<~�a<*�a<�a<��a<z�a<%�a<�a<��a<U�a<�a<��a<]�a<��a<��a<Q�a<��a<��a<-�a<ןa<{�a<$�a<��a<O�a<ԝa<h�a<�a<��a<�a<��a<$�a<��a<S�a<�a<s�a<�a<��a<�a<��a<P�a<ؖa<Y�a<ەa<_�a<�a<��a<�a<��a</�a<Ԓa<[�a<	�a<��a<�a<��a<N�a<��a<��a<4�a<��a<t�a<�a<ԍa<��a<:�a<׌a<��a<8�a<�a<��a<m�a< �a<��a<��a<��a<H�a<&�a<�a<ŉa<��a<��a<u�a<^�a<0�a<�a<��a<�a<�a<�a<ڈa<шa<؈a<Ԉa<��a<�a<�a<�a<�a<3�a<G�a<�  �  N�a<��a<��a<ʉa<�a< �a<R�a<p�a<a<֊a<-�a<Q�a<��a<�a<�a<��a<��a<�a<j�a<��a<"�a<d�a<ێa<�a<��a<��a<��a<�a<(�a<ȑa<�a<��a<��a<`�a<ѓa<:�a<Ҕa<7�a<Еa<$�a<Ŗa<3�a<��a<Q�a<��a<*�a<��a<��a<z�a<��a<��a<�a<|�a<Μa<n�a<՝a<D�a<Ӟa<�a<��a<�a<��a<�a<L�a<��a<�a<��a<�a<z�a<��a<�a<v�a<��a<�a<C�a<��a<ʥa<�a<f�a<��a<��a<�a<��a<��a<ܧa<#�a<&�a<z�a<k�a<��a<Ǩa<��a<�a<:�a<_�a<a�a<��a<��a<թa<�a<�a<�a<
�a<B�a<6�a<P�a<>�a<n�a<q�a<x�a<��a<e�a<��a<�a<o�a<��a<c�a<g�a<=�a<L�a<5�a<:�a<�a<�a<�a<ɩa<�a<��a<��a<��a<7�a<:�a<�a<��a<��a<��a<i�a<L�a<4�a<�a<�a<��a<n�a<@�a<�a<�a<��a<u�a<�a<�a<��a<��a<X�a<�a<�a<f�a<8�a<�a<��a<D�a<�a<��a<P�a<�a<��a<k�a<�a<��a<m�a<ԟa<��a<�a<��a<2�a<ʝa<s�a<�a<��a<�a<��a<=�a<Śa<m�a<͙a<}�a<��a<��a<�a<��a<1�a<��a<l�a<ٕa<��a<��a<��a<8�a<��a<T�a<ǒa<h�a<�a<{�a< �a<��a<g�a<�a<��a<+�a<�a<��a<�a<�a<Y�a<*�a<a<��a<2�a<�a<��a<N�a<A�a<�a<��a<��a<9�a<.�a<މa<݉a<��a<��a<I�a<S�a<5�a< �a<3�a<�a<�a<�a<Ԉa<�a<Јa<߈a<ǈa<�a<�a<�a<�a<-�a<d�a<�  �  f�a<�a<��a<Љa<��a<%�a<k�a<}�a<Êa<�a<#�a<g�a<��a<ۋa<%�a<m�a<��a<!�a<a�a<��a<$�a<w�a<��a<<�a<��a<��a<b�a<ʐa<:�a<��a<�a<��a<�a<k�a<�a<D�a<ߔa<.�a<��a<0�a<��a<#�a<��a<�a<��a<%�a<��a<#�a<��a<�a<��a<��a<x�a<�a<Q�a<˝a<?�a<��a<1�a<��a<�a<��a<�a<f�a<ܡa<1�a<��a<�a<K�a<��a<��a<Y�a<��a<�a<8�a<��a<٥a<&�a<r�a<��a<�a<"�a<e�a<��a<ϧa<��a<+�a<l�a<��a<Шa<بa<�a<#�a<7�a<k�a<t�a<��a<��a<©a<ԩa<��a<�a<�a<F�a<@�a<k�a<i�a<p�a<t�a<p�a<v�a<{�a<y�a<z�a<}�a<e�a<_�a<t�a<K�a<[�a<6�a<�a<&�a<�a<��a<�a<éa<��a<��a<|�a<\�a<S�a<�a< �a<èa<��a<�a<D�a<�a<�a<§a<��a<{�a<6�a<�a<�a<��a<��a<>�a<�a<¥a<��a<@�a<�a<��a<r�a<9�a<գa<��a<U�a<�a<Ģa<H�a<�a<��a<R�a<�a<��a<:�a<՟a<��a<�a<��a<O�a<ӝa<x�a<��a<��a< �a<��a<3�a<��a<N�a<�a<�a<�a<��a<�a<��a<Q�a<͖a<b�a<ܕa<m�a<��a<��a<�a<��a<B�a<��a<t�a<�a<��a<-�a<��a<b�a<�a<��a<6�a<َa<{�a<�a<ۍa<}�a<C�a<ӌa<��a<>�a<�a<��a<a�a< �a<�a<��a<q�a<R�a<#�a<�a<�a<��a<��a<t�a<U�a<8�a<�a<�a<��a<�a<�a<�a<̈a<̈a<�a<Ԉa<��a<�a<��a<"�a<,�a<H�a<�  �  ��a<z�a<��a<̉a<�a<'�a<F�a<�a<��a<��a<�a<\�a<��a<�a<?�a<r�a<ˌa<�a<h�a<͍a<�a<z�a<͎a<<�a<��a<�a<k�a<Đa<O�a<��a<�a<z�a<�a<_�a<ғa<A�a<��a<<�a<��a<1�a<��a<(�a<��a<�a<��a<�a<��a<�a<��a<�a<w�a<�a<\�a<�a<S�a<ޝa<X�a<��a<;�a<��a<�a<��a<�a<]�a<��a<0�a<��a<�a<C�a<��a<�a<N�a<��a<��a<K�a<��a<ҥa<�a<a�a<��a<�a<&�a<T�a<��a<̧a< �a<H�a<Q�a<��a<��a<٨a<��a<(�a<B�a<S�a<��a<��a<ũa<̩a<ݩa<��a<��a<2�a<(�a<@�a<K�a<b�a<`�a<g�a<��a<m�a<��a<s�a<s�a<q�a<g�a<f�a<V�a<L�a<?�a<:�a<(�a<�a<�a<�a<��a<��a<ȩa<��a<o�a<^�a<.�a<�a<�a<بa<��a<u�a<O�a<#�a<�a<ȧa<��a<d�a<=�a<�a<Ҧa<��a<g�a<>�a<�a<ӥa<��a<:�a<�a<��a<x�a<(�a<�a<��a<E�a<�a<��a<V�a<��a<��a<L�a<��a<��a<.�a<��a<k�a<�a<��a<B�a<ӝa<c�a<
�a<z�a<&�a<��a<F�a<ٚa<O�a<�a<a�a<�a<��a<�a<��a<3�a<̖a<F�a<��a<d�a<
�a<��a<�a<��a<6�a<Βa<V�a<�a<��a<�a<��a<Q�a<��a<��a<H�a<׎a<}�a<;�a<��a<}�a<�a<Ԍa<}�a<C�a<�a<��a<r�a<%�a<�a<��a<z�a<N�a<�a<�a<a<��a<��a<m�a<D�a<*�a<;�a<��a<�a<�a<܈a<׈a<Έa<ӈa<ψa<ֈa<ވa<�a< �a<�a<,�a<@�a<�  �  W�a<��a<��a<��a<�a< �a<E�a<��a<��a<ߊa<&�a<h�a<��a<�a<�a<~�a<Ȍa<�a<l�a<��a<$�a<��a<͎a<<�a<��a<�a<e�a<Ӑa<)�a<��a<�a<x�a<�a<Q�a<ٓa<P�a<��a<0�a<��a<"�a<��a<!�a<��a<�a<��a<�a<��a<�a<��a<#�a<z�a<�a<y�a<�a<_�a<ѝa<C�a<��a<4�a<��a<�a<��a<	�a<n�a<��a<C�a<��a<�a<J�a<��a<��a<b�a<��a<�a<>�a<��a<�a<&�a<Z�a<��a<�a<�a<d�a<��a<Чa<��a<#�a<_�a<��a<��a<��a<
�a<�a<A�a<j�a<�a<��a<��a<ѩa<�a<��a<�a<�a</�a<g�a<J�a<Y�a<~�a<[�a<t�a<|�a<r�a<x�a<��a<f�a<r�a<Z�a<[�a<U�a<E�a<*�a<0�a<�a<�a<�a<ҩa<ͩa<��a<��a<��a<W�a<-�a<:�a<�a<��a<��a<��a<X�a<,�a<�a<ӧa<��a<t�a<B�a<�a<�a<Ŧa<g�a<>�a<�a<��a<��a<I�a<�a<��a<x�a<&�a<�a<��a<K�a<��a<��a<J�a<��a<��a<_�a<�a<��a<9�a<ӟa<m�a<)�a<��a<K�a<��a<f�a<��a<��a< �a<��a<9�a<Ěa<X�a<�a<��a<��a<��a<7�a<��a<3�a<ߖa<L�a<וa<k�a<��a<�a<$�a<��a<2�a<��a<Y�a<��a<��a<�a<��a<N�a<�a<��a<(�a<ڎa<z�a<�a<͍a<��a<�a<�a<��a<4�a<�a<��a<l�a<-�a<��a<��a<��a<S�a<$�a<�a<ɉa<͉a<��a<d�a<c�a<�a<�a<�a<��a<�a<�a<ˈa<؈a<ǈa<Ԉa<ވa<�a<�a<�a<
�a<6�a<F�a<�  �  [�a<��a<��a<߉a<�a<�a<[�a<|�a<��a<�a<:�a<q�a<��a<��a<(�a<��a<��a<.�a<s�a<ōa<�a<x�a<�a<4�a<��a<
�a<e�a<אa<0�a<��a<�a<��a<�a<R�a<ٓa<?�a<Ŕa<"�a<ȕa<$�a<��a<�a<��a<&�a<��a<-�a<��a<�a<��a<�a<��a<�a<��a<�a<b�a<ޝa<Q�a<ʞa<(�a<şa<�a<��a<�a<i�a<̡a<.�a<��a<�a<Q�a<��a<��a<Y�a<��a<�a<-�a<��a<ҥa< �a<Z�a<��a<��a<�a<`�a<��a<֧a<��a<8�a<t�a<��a<��a<ݨa<��a<%�a<A�a<|�a<n�a<��a<��a<ީa<ܩa<�a<(�a< �a<7�a<B�a<`�a<`�a<v�a<��a<n�a<��a<r�a<t�a<p�a<u�a<y�a<H�a<b�a<@�a<M�a<�a<2�a<#�a<��a<�a<֩a<Щa<��a<��a<��a<V�a<C�a<�a<�a<ɨa<��a<��a<C�a<8�a<��a<ާa<��a<��a<H�a<�a<ަa<��a<��a<5�a<�a<Υa<��a<M�a<��a<��a<j�a<>�a<ڣa<��a<L�a<�a<��a<;�a<�a<��a<N�a<�a<��a<A�a<ڟa<��a<�a<��a<O�a<؝a<w�a<��a<��a<�a<��a<E�a<Қa<e�a<ݙa<��a<�a<��a<�a<��a<A�a<ʖa<g�a<�a<s�a<�a<��a<�a<��a<M�a<��a<\�a<�a<��a<�a<��a<g�a<�a<��a<-�a<�a<|�a<+�a<�a<x�a<1�a<ٌa<��a<@�a<�a<ɋa<[�a<:�a<�a<Ȋa<z�a<W�a<:�a<�a<щa<��a<��a<k�a<[�a<F�a<�a<�a<�a<�a<؈a<ڈa<��a<��a<ۈa<Ɉa<�a<ֈa<
�a<�a<$�a<B�a<�  �  ��a<v�a<��a<މa<�a<(�a<Y�a<w�a<��a<��a<"�a<p�a<��a<�a<<�a<��a<ǌa<&�a<f�a<ԍa<!�a<z�a<ݎa<7�a<��a<�a<\�a<Ða<S�a<��a<��a<y�a<�a<]�a<̓a<3�a<��a<0�a<��a<%�a<��a<.�a<��a<�a<��a<�a<��a<�a<��a<��a<��a<��a<s�a<�a<c�a<�a<]�a<Ǟa<8�a<��a<�a<��a<�a<c�a<ša<"�a<��a<�a<B�a<��a<�a<I�a<��a<��a<<�a<��a<ĥa<�a<\�a<��a<�a<�a<Q�a<��a<˧a<��a<F�a<S�a<��a<��a<�a< �a<5�a<=�a<k�a<~�a<��a<éa<ةa<ީa<�a<�a<1�a<<�a<<�a<]�a<d�a<U�a<|�a<v�a<k�a<��a<y�a<f�a<k�a<f�a<]�a<W�a<2�a<B�a<5�a<%�a<�a<��a<�a<��a<��a<��a<��a<c�a<_�a<A�a<�a<��a<ۨa<��a<��a<L�a<0�a<	�a<קa<��a<��a<<�a<!�a<�a<��a<w�a<8�a<�a<֥a<{�a<:�a<�a<��a<d�a<'�a<ۣa<��a<?�a<�a<��a<J�a<�a<��a<B�a<��a<��a<1�a<�a<s�a<�a<��a<I�a<ѝa<z�a<��a<��a<*�a<��a<P�a<ޚa<b�a<�a<z�a<�a<��a<�a<��a<:�a<��a<M�a<��a<c�a<�a<��a<�a<��a<7�a<��a<O�a<ۑa<y�a<�a<��a<R�a<�a<��a<M�a<֎a<q�a<9�a<��a<t�a<)�a<݌a<��a<P�a<�a<��a<k�a<4�a<��a<a<{�a<[�a<!�a<�a<։a<��a<��a<o�a<:�a<@�a<�a<��a<�a<�a<ψa<Јa<͈a<ʈa<Јa<��a<��a<�a<��a<�a<�a<C�a<�  �  _�a<v�a<��a<ĉa<��a<8�a<H�a<��a<��a<�a<)�a<j�a<��a<�a<3�a<�a<Ҍa<�a<s�a<ƍa<�a<��a<Ύa<Y�a<��a<��a<d�a<a<,�a<��a<�a<c�a<�a<M�a<˓a<Q�a<��a<8�a<��a<(�a<��a<�a<��a<�a<��a<
�a<��a<�a<��a<�a<{�a<�a<x�a<��a<d�a<ޝa<P�a<Ğa<E�a<��a<�a<��a<�a<l�a<��a<J�a<��a<�a<@�a<��a<�a<M�a<��a<ڤa<C�a<z�a<ݥa<�a<N�a<��a<ʦa<(�a<M�a<��a<ŧa<��a<,�a<S�a<��a<��a<��a<�a<$�a<L�a<f�a<��a<��a<��a<ҩa<�a<�a<�a<.�a<4�a<e�a<K�a<l�a<u�a<d�a<x�a<i�a<w�a<h�a<z�a<e�a<X�a<^�a<L�a<W�a<6�a</�a<�a<�a<�a<�a<کa<��a<��a<��a<{�a<o�a<0�a<7�a<�a<Ҩa<��a<��a<]�a<+�a< �a<ԧa<��a<u�a<I�a<�a<ݦa<Ȧa<i�a<Z�a<��a<��a<��a<8�a<��a<��a<{�a<�a<٣a<��a<=�a<��a<��a<R�a<�a<��a<O�a<�a<��a<.�a<ݟa<i�a<.�a<��a<K�a<�a<g�a<�a<��a<.�a<��a<F�a<њa<_�a<��a<�a<�a<��a<0�a<��a<6�a<�a<F�a<�a<b�a<��a<|�a<�a<��a<�a<ƒa<E�a<��a<��a<�a<��a<8�a<��a<��a<*�a<Ўa<y�a< �a<a<��a<�a<�a<��a<?�a<��a<��a<v�a<2�a<�a<��a<��a<Y�a<%�a<�a<ωa<ʉa<��a<v�a<Z�a<'�a< �a<��a<��a<وa<�a<ʈa<��a<ˈa<ňa<��a<Ոa<�a<��a<�a<1�a<6�a<�  �  \�a<��a<��a<щa<��a< �a<M�a<��a<��a<�a<<�a<`�a<��a<�a<3�a<��a<Ȍa<�a<}�a<͍a<"�a<�a<ڎa<6�a<��a<�a<p�a<��a<+�a<��a<�a<x�a<�a<E�a<��a<4�a<��a<'�a<��a<�a<��a<#�a<��a<7�a<��a<'�a<��a<�a<��a<�a<��a<��a<��a<�a<z�a<�a<W�a<��a</�a<��a<�a<��a<��a<g�a<ǡa<'�a<��a<�a<a�a<��a<��a<T�a<��a<��a<7�a<y�a<åa<
�a<J�a<��a<�a<�a<f�a<��a<٧a<�a<5�a<j�a<��a<��a<�a<�a<*�a<M�a<m�a<|�a<©a<��a<�a<��a<��a<%�a<(�a<@�a<L�a<Q�a<]�a<i�a<u�a<w�a<��a<s�a<}�a<h�a<a�a<n�a<P�a<F�a<?�a</�a<#�a<(�a<�a<��a<��a<שa<�a<��a<��a<y�a<W�a<5�a<�a<��a<Ѩa<��a<x�a<]�a<E�a< �a<�a<��a<v�a<R�a<�a<�a<��a<t�a<7�a<�a<ɥa<��a<V�a<��a<Ťa<h�a<&�a<٣a<z�a<2�a<�a<��a<A�a<�a<��a<M�a<�a<��a<R�a<ݟa<��a<�a<��a<J�a<ߝa<y�a<�a<��a<�a<ʛa<L�a<ؚa<{�a<�a<��a<�a<��a<%�a<��a<<�a<Öa<b�a<�a<��a<��a<��a<�a<��a<8�a<��a<D�a<ّa<q�a<�a<��a<P�a<�a<��a<(�a<�a<��a<(�a<ٍa<u�a<)�a<ތa<��a<E�a<��a<��a<i�a<T�a<�a<Ҋa<��a<M�a<7�a<��a<ډa<��a<��a<h�a<N�a<9�a<�a<#�a<�a<�a<шa<ƈa<Ոa<��a<��a<Ȉa<Έa<ۈa< �a<	�a<�a<N�a<�  �  L�a<��a<��a<܉a<�a<4�a<r�a<p�a<ۊa<�a<2�a<{�a<��a<��a<%�a<��a<Όa<7�a<n�a<֍a<9�a<l�a<�a<9�a<��a<��a<C�a<Đa<$�a<��a<�a<��a<͒a<[�a<ғa<4�a<̔a<�a<��a<�a<��a<�a<��a<�a<}�a<5�a<��a<:�a<��a<�a<��a<�a<��a<�a<o�a<ӝa<H�a<՞a<;�a<˟a<�a<��a<��a<h�a<�a<%�a<��a<Ӣa<D�a<��a<�a<K�a<��a<�a<�a<��a<ťa<�a<g�a<��a<�a<�a<b�a<��a<��a<�a<(�a<l�a<��a<�a<ըa<�a<>�a<A�a<��a<��a<��a<��a<֩a<�a<�a<!�a<�a<a�a<8�a<o�a<x�a<`�a<��a<S�a<y�a<a�a<|�a<_�a<k�a<]�a<I�a<b�a<7�a<J�a<%�a<�a<�a<�a<��a<ǩa<ȩa<��a<��a<r�a<k�a<Z�a<�a<�a<Ψa<��a<��a<X�a<6�a<�a<�a<��a<��a<C�a<"�a<��a<��a<��a<:�a<�a<åa<b�a<:�a<�a<¤a<T�a<1�a<��a<��a<E�a<�a<��a<+�a<��a<��a<B�a<�a<��a<:�a<��a<��a<
�a<՞a<S�a<֝a<��a<��a<��a<)�a<��a<;�a<ɚa<p�a<�a<��a<�a<��a<%�a<��a<h�a<��a<o�a<ƕa<e�a<�a<z�a<�a<��a<2�a<��a<d�a<ܑa<~�a<!�a<��a<W�a<ԏa<��a< �a<Ǝa<c�a<�a<ڍa<t�a<Z�a<Ќa<��a<Y�a<�a<ҋa<r�a<F�a<�a<��a<��a<e�a<3�a<�a<��a<��a<��a<��a<E�a<I�a<��a<
�a<߈a<�a<Ȉa<Јa<Ĉa<��a<ۈa<��a<�a<ވa<�a<�a<�a<M�a<�  �  \�a<��a<��a<��a<�a<!�a<>�a<��a<��a<��a<*�a<p�a<��a<��a<W�a<��a<׌a<�a<w�a<ˍa<"�a<v�a<Ɏa<8�a<��a<�a<o�a<Րa<.�a<��a<�a<x�a<ߒa<U�a<��a<0�a<��a<2�a<��a<4�a<��a<�a<��a<0�a<��a<�a<��a<�a<z�a<
�a<��a<�a<s�a<��a<j�a<��a<o�a<˞a<H�a<��a<"�a<��a<��a<O�a<��a<'�a<��a<��a<^�a<��a<��a<K�a<��a<�a<;�a<}�a<��a<��a<V�a<��a<ݦa<�a<S�a<��a<էa<�a<A�a<a�a<��a<��a<֨a<�a<)�a<N�a<c�a<��a<��a<ܩa<�a<�a<
�a<�a<1�a<@�a<J�a<=�a<[�a<b�a<�a<�a<��a<t�a<j�a<j�a<u�a<X�a<[�a<A�a<5�a<'�a</�a<�a<�a<��a<�a<שa<ѩa<��a<��a<q�a<X�a<&�a<�a<��a<بa<��a<��a<Z�a<8�a<$�a<֧a<��a<w�a<M�a<�a<�a<��a<d�a<:�a<��a<ҥa<��a<K�a<��a<��a<j�a<&�a<ңa<��a<#�a<ݢa<��a<L�a<�a<��a<E�a<�a<��a<L�a<�a<~�a<�a<��a<2�a<ܝa<v�a<
�a<��a<1�a<��a<^�a<�a<f�a<��a<x�a<�a<��a<$�a<��a<.�a<Öa<Z�a<�a<��a< �a<}�a<�a<��a<)�a<��a<H�a<ёa<b�a<�a<��a<L�a<�a<��a<*�a<ߎa<��a<4�a<Ѝa<x�a<�a<ьa<��a<C�a< �a<��a<}�a<5�a<�a<̊a<��a<_�a<$�a<�a<ډa<��a<s�a<f�a<G�a<C�a<'�a<�a<�a<ۈa<ӈa<ۈa<��a<Ɉa<��a<��a<ƈa<�a<��a<�a<#�a<6�a<�  �  r�a<j�a<��a<��a<�a<B�a<J�a<��a<��a<�a<@�a<m�a<��a<�a<M�a<j�a<�a<�a<��a<ƍa<�a<��a<̎a<a�a<��a<�a<T�a<��a<?�a<��a<	�a<P�a<�a<V�a<��a<U�a<��a<E�a<��a<�a<��a<(�a<��a<�a<��a<��a<��a<#�a<��a<*�a<k�a<*�a<t�a<�a<a�a<؝a<Q�a<��a<Y�a<��a<J�a<u�a<�a<��a<Сa<Q�a<{�a<�a<5�a<��a<�a<J�a<��a<Ǥa<L�a<j�a<ߥa<�a<Q�a<��a<��a<!�a<X�a<��a<��a<�a<'�a<_�a<��a<��a<�a<�a<�a<z�a<_�a<��a<��a<ʩa<ʩa<�a<�a<#�a<L�a<�a<w�a<T�a<|�a<~�a<Y�a<i�a<_�a<��a<w�a<g�a<R�a<J�a<l�a<1�a<Y�a<�a<:�a<�a<�a<��a<�a<�a<��a<��a<��a<��a<y�a<2�a<L�a<ըa<�a<��a<��a<b�a<$�a<�a<��a<��a<q�a<q�a<�a<Ѧa<ߦa<f�a<c�a<�a<��a<s�a<2�a<�a<��a<n�a<��a<ߣa<��a<*�a<�a<y�a<_�a<ϡa<��a<B�a<��a<��a<#�a<ܟa<^�a<6�a<��a<^�a<��a<W�a<0�a<��a<A�a<��a<@�a<Қa<U�a<�a<s�a<9�a<��a<9�a<ӗa<E�a<�a<A�a<��a<V�a<��a<��a<�a<��a<�a<Вa<5�a<��a<w�a<�a<��a<&�a<��a<��a<7�a<ʎa<f�a<�a<͍a<��a<�a<�a<��a<6�a<,�a<��a<��a<�a<�a<��a<��a<`�a<5�a< �a<��a<݉a<��a<��a<c�a<�a<�a<�a<�a<�a<Јa<��a<��a<وa<��a<�a<��a<�a<�a<�a<�a<@�a<�  �  \�a<��a<��a<��a<�a<!�a<>�a<��a<��a<��a<*�a<p�a<��a<��a<W�a<��a<׌a<�a<w�a<ˍa<"�a<v�a<Ɏa<8�a<��a<�a<o�a<Րa<.�a<��a<�a<x�a<ߒa<U�a<��a<0�a<��a<2�a<��a<4�a<��a<�a<��a<0�a<��a<�a<��a<�a<z�a<
�a<��a<�a<s�a<��a<j�a<��a<o�a<˞a<H�a<��a<"�a<��a<��a<O�a<��a<'�a<��a<��a<^�a<��a<��a<K�a<��a<�a<;�a<}�a<��a<��a<V�a<��a<ݦa<�a<S�a<��a<էa<�a<A�a<a�a<��a<��a<֨a<�a<)�a<N�a<c�a<��a<��a<ܩa<�a<�a<
�a<�a<1�a<@�a<J�a<=�a<[�a<b�a<�a<�a<��a<t�a<j�a<j�a<u�a<X�a<[�a<A�a<5�a<'�a</�a<�a<�a<��a<�a<שa<ѩa<��a<��a<q�a<X�a<&�a<�a<��a<بa<��a<��a<Z�a<8�a<$�a<֧a<��a<w�a<M�a<�a<�a<��a<d�a<:�a<��a<ҥa<��a<K�a<��a<��a<j�a<&�a<ңa<��a<#�a<ݢa<��a<L�a<�a<��a<E�a<�a<��a<L�a<�a<~�a<�a<��a<2�a<ܝa<v�a<
�a<��a<1�a<��a<^�a<�a<f�a<��a<x�a<�a<��a<$�a<��a<.�a<Öa<Z�a<�a<��a< �a<}�a<�a<��a<)�a<��a<H�a<ёa<b�a<�a<��a<L�a<�a<��a<*�a<ߎa<��a<4�a<Ѝa<x�a<�a<ьa<��a<C�a< �a<��a<}�a<5�a<�a<̊a<��a<_�a<$�a<�a<ډa<��a<s�a<f�a<G�a<C�a<'�a<�a<�a<ۈa<ӈa<ۈa<��a<Ɉa<��a<��a<ƈa<�a<��a<�a<#�a<6�a<�  �  L�a<��a<��a<܉a<�a<4�a<r�a<p�a<ۊa<�a<2�a<{�a<��a<��a<%�a<��a<Όa<7�a<n�a<֍a<9�a<l�a<�a<9�a<��a<��a<C�a<Đa<$�a<��a<�a<��a<͒a<[�a<ғa<4�a<̔a<�a<��a<�a<��a<�a<��a<�a<}�a<5�a<��a<:�a<��a<�a<��a<�a<��a<�a<o�a<ӝa<H�a<՞a<;�a<˟a<�a<��a<��a<h�a<�a<%�a<��a<Ӣa<D�a<��a<�a<K�a<��a<�a<�a<��a<ťa<�a<g�a<��a<�a<�a<b�a<��a<��a<�a<(�a<l�a<��a<�a<ըa<�a<>�a<A�a<��a<��a<��a<��a<֩a<�a<�a<!�a<�a<a�a<8�a<o�a<x�a<`�a<��a<S�a<y�a<a�a<|�a<_�a<k�a<]�a<I�a<b�a<7�a<J�a<%�a<�a<�a<�a<��a<ǩa<ȩa<��a<��a<r�a<k�a<Z�a<�a<�a<Ψa<��a<��a<X�a<6�a<�a<�a<��a<��a<C�a<"�a<��a<��a<��a<:�a<�a<åa<b�a<:�a<�a<¤a<T�a<1�a<��a<��a<E�a<�a<��a<+�a<��a<��a<B�a<�a<��a<:�a<��a<��a<
�a<՞a<S�a<֝a<��a<��a<��a<)�a<��a<;�a<ɚa<p�a<�a<��a<�a<��a<%�a<��a<h�a<��a<o�a<ƕa<e�a<�a<z�a<�a<��a<2�a<��a<d�a<ܑa<~�a<!�a<��a<W�a<ԏa<��a< �a<Ǝa<c�a<�a<ڍa<t�a<Z�a<Ќa<��a<Y�a<�a<ҋa<r�a<F�a<�a<��a<��a<e�a<3�a<�a<��a<��a<��a<��a<E�a<I�a<��a<
�a<߈a<�a<Ȉa<Јa<Ĉa<��a<ۈa<��a<�a<ވa<�a<�a<�a<M�a<�  �  \�a<��a<��a<щa<��a< �a<M�a<��a<��a<�a<<�a<`�a<��a<�a<3�a<��a<Ȍa<�a<}�a<͍a<"�a<�a<ڎa<6�a<��a<�a<p�a<��a<+�a<��a<�a<x�a<�a<E�a<��a<4�a<��a<'�a<��a<�a<��a<#�a<��a<7�a<��a<'�a<��a<�a<��a<�a<��a<��a<��a<�a<z�a<�a<W�a<��a</�a<��a<�a<��a<��a<g�a<ǡa<'�a<��a<�a<a�a<��a<��a<T�a<��a<��a<7�a<y�a<åa<
�a<J�a<��a<�a<�a<f�a<��a<٧a<�a<5�a<j�a<��a<��a<�a<�a<*�a<M�a<m�a<|�a<©a<��a<�a<��a<��a<%�a<(�a<@�a<L�a<Q�a<]�a<i�a<u�a<w�a<��a<s�a<}�a<h�a<a�a<n�a<P�a<F�a<?�a</�a<#�a<(�a<�a<��a<��a<שa<�a<��a<��a<y�a<W�a<5�a<�a<��a<Ѩa<��a<x�a<]�a<E�a< �a<�a<��a<v�a<R�a<�a<�a<��a<t�a<7�a<�a<ɥa<��a<V�a<��a<Ťa<h�a<&�a<٣a<z�a<2�a<�a<��a<A�a<�a<��a<M�a<�a<��a<R�a<ݟa<��a<�a<��a<J�a<ߝa<y�a<�a<��a<�a<ʛa<L�a<ؚa<{�a<�a<��a<�a<��a<%�a<��a<<�a<Öa<b�a<�a<��a<��a<��a<�a<��a<8�a<��a<D�a<ّa<q�a<�a<��a<P�a<�a<��a<(�a<�a<��a<(�a<ٍa<u�a<)�a<ތa<��a<E�a<��a<��a<i�a<T�a<�a<Ҋa<��a<M�a<7�a<��a<ډa<��a<��a<h�a<N�a<9�a<�a<#�a<�a<�a<шa<ƈa<Ոa<��a<��a<Ȉa<Έa<ۈa< �a<	�a<�a<N�a<�  �  _�a<v�a<��a<ĉa<��a<8�a<H�a<��a<��a<�a<)�a<j�a<��a<�a<3�a<�a<Ҍa<�a<s�a<ƍa<�a<��a<Ύa<Y�a<��a<��a<d�a<a<,�a<��a<�a<c�a<�a<M�a<˓a<Q�a<��a<8�a<��a<(�a<��a<�a<��a<�a<��a<
�a<��a<�a<��a<�a<{�a<�a<x�a<��a<d�a<ޝa<P�a<Ğa<E�a<��a<�a<��a<�a<l�a<��a<J�a<��a<�a<@�a<��a<�a<M�a<��a<ڤa<C�a<z�a<ݥa<�a<N�a<��a<ʦa<(�a<M�a<��a<ŧa<��a<,�a<S�a<��a<��a<��a<�a<$�a<L�a<f�a<��a<��a<��a<ҩa<�a<�a<�a<.�a<4�a<e�a<K�a<l�a<u�a<d�a<x�a<i�a<w�a<h�a<z�a<e�a<X�a<^�a<L�a<W�a<6�a</�a<�a<�a<�a<�a<کa<��a<��a<��a<{�a<o�a<0�a<7�a<�a<Ҩa<��a<��a<]�a<+�a< �a<ԧa<��a<u�a<I�a<�a<ݦa<Ȧa<i�a<Z�a<��a<��a<��a<8�a<��a<��a<{�a<�a<٣a<��a<=�a<��a<��a<R�a<�a<��a<O�a<�a<��a<.�a<ݟa<i�a<.�a<��a<K�a<�a<g�a<�a<��a<.�a<��a<F�a<њa<_�a<��a<�a<�a<��a<0�a<��a<6�a<�a<F�a<�a<b�a<��a<|�a<�a<��a<�a<ƒa<E�a<��a<��a<�a<��a<8�a<��a<��a<*�a<Ўa<y�a< �a<a<��a<�a<�a<��a<?�a<��a<��a<v�a<2�a<�a<��a<��a<Y�a<%�a<�a<ωa<ʉa<��a<v�a<Z�a<'�a< �a<��a<��a<وa<�a<ʈa<��a<ˈa<ňa<��a<Ոa<�a<��a<�a<1�a<6�a<�  �  ��a<v�a<��a<މa<�a<(�a<Y�a<w�a<��a<��a<"�a<p�a<��a<�a<<�a<��a<ǌa<&�a<f�a<ԍa<!�a<z�a<ݎa<7�a<��a<�a<\�a<Ða<S�a<��a<��a<y�a<�a<]�a<̓a<3�a<��a<0�a<��a<%�a<��a<.�a<��a<�a<��a<�a<��a<�a<��a<��a<��a<��a<s�a<�a<c�a<�a<]�a<Ǟa<8�a<��a<�a<��a<�a<c�a<ša<"�a<��a<�a<B�a<��a<�a<I�a<��a<��a<<�a<��a<ĥa<�a<\�a<��a<�a<�a<Q�a<��a<˧a<��a<F�a<S�a<��a<��a<�a< �a<5�a<=�a<k�a<~�a<��a<éa<ةa<ީa<�a<�a<1�a<<�a<<�a<]�a<d�a<U�a<|�a<v�a<k�a<��a<y�a<f�a<k�a<f�a<]�a<W�a<2�a<B�a<5�a<%�a<�a<��a<�a<��a<��a<��a<��a<c�a<_�a<A�a<�a<��a<ۨa<��a<��a<L�a<0�a<	�a<קa<��a<��a<<�a<!�a<�a<��a<w�a<8�a<�a<֥a<{�a<:�a<�a<��a<d�a<'�a<ۣa<��a<?�a<�a<��a<J�a<�a<��a<B�a<��a<��a<1�a<�a<s�a<�a<��a<I�a<ѝa<z�a<��a<��a<*�a<��a<P�a<ޚa<b�a<�a<z�a<�a<��a<�a<��a<:�a<��a<M�a<��a<c�a<�a<��a<�a<��a<7�a<��a<O�a<ۑa<y�a<�a<��a<R�a<�a<��a<M�a<֎a<q�a<9�a<��a<t�a<)�a<݌a<��a<P�a<�a<��a<k�a<4�a<��a<a<{�a<[�a<!�a<�a<։a<��a<��a<o�a<:�a<@�a<�a<��a<�a<�a<ψa<Јa<͈a<ʈa<Јa<��a<��a<�a<��a<�a<�a<C�a<�  �  [�a<��a<��a<߉a<�a<�a<[�a<|�a<��a<�a<:�a<q�a<��a<��a<(�a<��a<��a<.�a<s�a<ōa<�a<x�a<�a<4�a<��a<
�a<e�a<אa<0�a<��a<�a<��a<�a<R�a<ٓa<?�a<Ŕa<"�a<ȕa<$�a<��a<�a<��a<&�a<��a<-�a<��a<�a<��a<�a<��a<�a<��a<�a<b�a<ޝa<Q�a<ʞa<(�a<şa<�a<��a<�a<i�a<̡a<.�a<��a<�a<Q�a<��a<��a<Y�a<��a<�a<-�a<��a<ҥa< �a<Z�a<��a<��a<�a<`�a<��a<֧a<��a<8�a<t�a<��a<��a<ݨa<��a<%�a<A�a<|�a<n�a<��a<��a<ީa<ܩa<�a<(�a< �a<7�a<B�a<`�a<`�a<v�a<��a<n�a<��a<r�a<t�a<p�a<u�a<y�a<H�a<b�a<@�a<M�a<�a<2�a<#�a<��a<�a<֩a<Щa<��a<��a<��a<V�a<C�a<�a<�a<ɨa<��a<��a<C�a<8�a<��a<ާa<��a<��a<H�a<�a<ަa<��a<��a<5�a<�a<Υa<��a<M�a<��a<��a<j�a<>�a<ڣa<��a<L�a<�a<��a<;�a<�a<��a<N�a<�a<��a<A�a<ڟa<��a<�a<��a<O�a<؝a<w�a<��a<��a<�a<��a<E�a<Қa<e�a<ݙa<��a<�a<��a<�a<��a<A�a<ʖa<g�a<�a<s�a<�a<��a<�a<��a<M�a<��a<\�a<�a<��a<�a<��a<g�a<�a<��a<-�a<�a<|�a<+�a<�a<x�a<1�a<ٌa<��a<@�a<�a<ɋa<[�a<:�a<�a<Ȋa<z�a<W�a<:�a<�a<щa<��a<��a<k�a<[�a<F�a<�a<�a<�a<�a<؈a<ڈa<��a<��a<ۈa<Ɉa<�a<ֈa<
�a<�a<$�a<B�a<�  �  W�a<��a<��a<��a<�a< �a<E�a<��a<��a<ߊa<&�a<h�a<��a<�a<�a<~�a<Ȍa<�a<l�a<��a<$�a<��a<͎a<<�a<��a<�a<e�a<Ӑa<)�a<��a<�a<x�a<�a<Q�a<ٓa<P�a<��a<0�a<��a<"�a<��a<!�a<��a<�a<��a<�a<��a<�a<��a<#�a<z�a<�a<y�a<�a<_�a<ѝa<C�a<��a<4�a<��a<�a<��a<	�a<n�a<��a<C�a<��a<�a<J�a<��a<��a<b�a<��a<�a<>�a<��a<�a<&�a<Z�a<��a<�a<�a<d�a<��a<Чa<��a<#�a<_�a<��a<��a<��a<
�a<�a<A�a<j�a<�a<��a<��a<ѩa<�a<��a<�a<�a</�a<g�a<J�a<Y�a<~�a<[�a<t�a<|�a<r�a<x�a<��a<f�a<r�a<Z�a<[�a<U�a<E�a<*�a<0�a<�a<�a<�a<ҩa<ͩa<��a<��a<��a<W�a<-�a<:�a<�a<��a<��a<��a<X�a<,�a<�a<ӧa<��a<t�a<B�a<�a<�a<Ŧa<g�a<>�a<�a<��a<��a<I�a<�a<��a<x�a<&�a<�a<��a<K�a<��a<��a<J�a<��a<��a<_�a<�a<��a<9�a<ӟa<m�a<)�a<��a<K�a<��a<f�a<��a<��a< �a<��a<9�a<Ěa<X�a<�a<��a<��a<��a<7�a<��a<3�a<ߖa<L�a<וa<k�a<��a<�a<$�a<��a<2�a<��a<Y�a<��a<��a<�a<��a<N�a<�a<��a<(�a<ڎa<z�a<�a<͍a<��a<�a<�a<��a<4�a<�a<��a<l�a<-�a<��a<��a<��a<S�a<$�a<�a<ɉa<͉a<��a<d�a<c�a<�a<�a<�a<��a<�a<�a<ˈa<؈a<ǈa<Ԉa<ވa<�a<�a<�a<
�a<6�a<F�a<�  �  ��a<z�a<��a<̉a<�a<'�a<F�a<�a<��a<��a<�a<\�a<��a<�a<?�a<r�a<ˌa<�a<h�a<͍a<�a<z�a<͎a<<�a<��a<�a<k�a<Đa<O�a<��a<�a<z�a<�a<_�a<ғa<A�a<��a<<�a<��a<1�a<��a<(�a<��a<�a<��a<�a<��a<�a<��a<�a<w�a<�a<\�a<�a<S�a<ޝa<X�a<��a<;�a<��a<�a<��a<�a<]�a<��a<0�a<��a<�a<C�a<��a<�a<N�a<��a<��a<K�a<��a<ҥa<�a<a�a<��a<�a<&�a<T�a<��a<̧a< �a<H�a<Q�a<��a<��a<٨a<��a<(�a<B�a<S�a<��a<��a<ũa<̩a<ݩa<��a<��a<2�a<(�a<@�a<K�a<b�a<`�a<g�a<��a<m�a<��a<s�a<s�a<q�a<g�a<f�a<V�a<L�a<?�a<:�a<(�a<�a<�a<�a<��a<��a<ȩa<��a<o�a<^�a<.�a<�a<�a<بa<��a<u�a<O�a<#�a<�a<ȧa<��a<d�a<=�a<�a<Ҧa<��a<g�a<>�a<�a<ӥa<��a<:�a<�a<��a<x�a<(�a<�a<��a<E�a<�a<��a<V�a<��a<��a<L�a<��a<��a<.�a<��a<k�a<�a<��a<B�a<ӝa<c�a<
�a<z�a<&�a<��a<F�a<ٚa<O�a<�a<a�a<�a<��a<�a<��a<3�a<̖a<F�a<��a<d�a<
�a<��a<�a<��a<6�a<Βa<V�a<�a<��a<�a<��a<Q�a<��a<��a<H�a<׎a<}�a<;�a<��a<}�a<�a<Ԍa<}�a<C�a<�a<��a<r�a<%�a<�a<��a<z�a<N�a<�a<�a<a<��a<��a<m�a<D�a<*�a<;�a<��a<�a<�a<܈a<׈a<Έa<ӈa<ψa<ֈa<ވa<�a< �a<�a<,�a<@�a<�  �  f�a<�a<��a<Љa<��a<%�a<k�a<}�a<Êa<�a<#�a<g�a<��a<ۋa<%�a<m�a<��a<!�a<a�a<��a<$�a<w�a<��a<<�a<��a<��a<b�a<ʐa<:�a<��a<�a<��a<�a<k�a<�a<D�a<ߔa<.�a<��a<0�a<��a<#�a<��a<�a<��a<%�a<��a<#�a<��a<�a<��a<��a<x�a<�a<Q�a<˝a<?�a<��a<1�a<��a<�a<��a<�a<f�a<ܡa<1�a<��a<�a<K�a<��a<��a<Y�a<��a<�a<8�a<��a<٥a<&�a<r�a<��a<�a<"�a<e�a<��a<ϧa<��a<+�a<l�a<��a<Шa<بa<�a<#�a<7�a<k�a<t�a<��a<��a<©a<ԩa<��a<�a<�a<F�a<@�a<k�a<i�a<p�a<t�a<p�a<v�a<{�a<y�a<z�a<}�a<e�a<_�a<t�a<K�a<[�a<6�a<�a<&�a<�a<��a<�a<éa<��a<��a<|�a<\�a<S�a<�a< �a<èa<��a<�a<D�a<�a<�a<§a<��a<{�a<6�a<�a<�a<��a<��a<>�a<�a<¥a<��a<@�a<�a<��a<r�a<9�a<գa<��a<U�a<�a<Ģa<H�a<�a<��a<R�a<�a<��a<:�a<՟a<��a<�a<��a<O�a<ӝa<x�a<��a<��a< �a<��a<3�a<��a<N�a<�a<�a<�a<��a<�a<��a<Q�a<͖a<b�a<ܕa<m�a<��a<��a<�a<��a<B�a<��a<t�a<�a<��a<-�a<��a<b�a<�a<��a<6�a<َa<{�a<�a<ۍa<}�a<C�a<ӌa<��a<>�a<�a<��a<a�a< �a<�a<��a<q�a<R�a<#�a<�a<�a<��a<��a<t�a<U�a<8�a<�a<�a<��a<�a<�a<�a<̈a<̈a<�a<Ԉa<��a<�a<��a<"�a<,�a<H�a<�  �  N�a<��a<��a<ʉa<�a< �a<R�a<p�a<a<֊a<-�a<Q�a<��a<�a<�a<��a<��a<�a<j�a<��a<"�a<d�a<ێa<�a<��a<��a<��a<�a<(�a<ȑa<�a<��a<��a<`�a<ѓa<:�a<Ҕa<7�a<Еa<$�a<Ŗa<3�a<��a<Q�a<��a<*�a<��a<��a<z�a<��a<��a<�a<|�a<Μa<n�a<՝a<D�a<Ӟa<�a<��a<�a<��a<�a<L�a<��a<�a<��a<�a<z�a<��a<�a<v�a<��a<�a<C�a<��a<ʥa<�a<f�a<��a<��a<�a<��a<��a<ܧa<#�a<&�a<z�a<k�a<��a<Ǩa<��a<�a<:�a<_�a<a�a<��a<��a<թa<�a<�a<�a<
�a<B�a<6�a<P�a<>�a<n�a<q�a<x�a<��a<e�a<��a<�a<o�a<��a<c�a<g�a<=�a<L�a<5�a<:�a<�a<�a<�a<ɩa<�a<��a<��a<��a<7�a<:�a<�a<��a<��a<��a<i�a<L�a<4�a<�a<�a<��a<n�a<@�a<�a<�a<��a<u�a<�a<�a<��a<��a<X�a<�a<�a<f�a<8�a<�a<��a<D�a<�a<��a<P�a<�a<��a<k�a<�a<��a<m�a<ԟa<��a<�a<��a<2�a<ʝa<s�a<�a<��a<�a<��a<=�a<Śa<m�a<͙a<}�a<��a<��a<�a<��a<1�a<��a<l�a<ٕa<��a<��a<��a<8�a<��a<T�a<ǒa<h�a<�a<{�a< �a<��a<g�a<�a<��a<+�a<�a<��a<�a<�a<Y�a<*�a<a<��a<2�a<�a<��a<N�a<A�a<�a<��a<��a<9�a<.�a<މa<݉a<��a<��a<I�a<S�a<5�a< �a<3�a<�a<�a<�a<Ԉa<�a<Јa<߈a<ǈa<�a<�a<�a<�a<-�a<d�a<�  �  a�a<p�a<��a<Ɖa<	�a<.�a<\�a<}�a<��a<�a<-�a<Z�a<��a<ыa<�a<j�a<Ȍa<�a<x�a<��a<�a<x�a<�a<E�a<��a<��a<_�a<��a<7�a<��a<�a<w�a<��a<a�a<�a<f�a<��a<C�a<��a<2�a<��a<'�a<��a<�a<��a<�a<��a<#�a<��a<�a<|�a<��a<o�a<�a<Z�a<��a<4�a<��a<1�a<��a<�a<��a<�a<h�a<ۡa<<�a<��a<�a<>�a<��a<��a<W�a<��a<�a<Q�a<��a<�a<3�a<d�a<��a<ߦa<(�a<c�a<��a<��a<��a<+�a<f�a<��a<Ǩa<ܨa<��a<�a<P�a<V�a<��a<��a<��a<��a<�a<�a<�a<!�a<+�a<A�a<_�a<j�a<y�a<l�a<t�a<f�a<u�a<z�a<z�a<u�a<j�a<j�a<[�a<q�a<K�a<9�a<,�a<�a<�a<��a<ܩa<��a<��a<��a<��a<e�a<D�a<�a<�a<ɨa<��a<s�a<Q�a<�a<�a<��a<��a<f�a<M�a<
�a<զa<��a<��a<F�a<�a<��a<~�a<*�a<�a<��a<z�a<%�a<�a<��a<U�a<�a<��a<]�a<��a<��a<Q�a<��a<��a<-�a<ןa<{�a<$�a<��a<O�a<ԝa<h�a<�a<��a<�a<��a<$�a<��a<S�a<�a<s�a<�a<��a<�a<��a<P�a<ؖa<Y�a<ەa<_�a<�a<��a<�a<��a</�a<Ԓa<[�a<	�a<��a<�a<��a<N�a<��a<��a<4�a<��a<t�a<�a<ԍa<��a<:�a<׌a<��a<8�a<�a<��a<m�a< �a<��a<��a<��a<H�a<&�a<�a<ŉa<��a<��a<u�a<^�a<0�a<�a<��a<�a<�a<�a<ڈa<шa<؈a<Ԉa<��a<�a<�a<�a<�a<3�a<G�a<�  �  m�a<~�a<̈a<ڈa<��a<$�a<8�a<��a<��a<�a<�a<]�a<��a<Պa<P�a<U�a<ۋa<�a<p�a<��a<!�a<��a<ύa<F�a<��a<(�a<��a<�a<J�a<��a<G�a<��a<�a<��a<ݒa<N�a<ߓa<u�a<єa<k�a<ݕa<Q�a<ϖa<@�a<�a<A�a<Řa<2�a<��a<@�a<��a<(�a<}�a</�a<�a<�a<��a<ڝa<��a<��a<U�a<��a<>�a<��a<��a<q�a<Сa<`�a<��a<��a<N�a<��a<�a<;�a<��a<ܤa<�a<W�a<��a<�a<&�a<��a<��a<�a<�a<U�a<��a<��a<ѧa<�a<$�a<E�a<X�a<��a<��a<רa<��a<�a<�a<�a<=�a<6�a<`�a<v�a<��a<z�a<��a<��a<��a<�a<��a<��a<��a<Щa<��a<��a<��a<��a<w�a<t�a<��a<s�a<[�a<g�a<2�a<'�a<�a<�a<ߨa<��a<��a<]�a<]�a<0�a<�a<˧a<��a<��a<O�a<W�a<�a<�a<��a<}�a<C�a<�a<�a<��a<{�a<9�a<�a<ۤa<��a<C�a<��a<ڣa<h�a<4�a<�a<x�a<#�a<�a<��a<?�a<�a<��a<=�a<��a<s�a<E�a<��a<T�a<ܝa<l�a<�a<��a<3�a<��a<e�a<˚a<|�a<�a<j�a<,�a<y�a<1�a<��a<T�a<̖a<O�a<�a<t�a<0�a<��a<&�a<��a<A�a<�a<M�a<��a<v�a<�a<��a<C�a<�a<^�a<)�a<��a<D�a<��a<��a<S�a<Ռa<��a<�a<�a<��a<5�a<��a<��a<��a<�a<�a<��a<u�a<S�a<�a<�a<Јa<��a<o�a<g�a<N�a<9�a<H�a<��a<��a<�a<��a<�a<ԇa<�a<͇a<��a<҇a<�a<�a<�a<K�a<E�a<�  �  y�a<��a<��a<Ĉa< �a<4�a<_�a<u�a<��a<�a<+�a<Q�a<��a<ӊa<�a<d�a<ŋa<�a<{�a<��a<�a<z�a<�a<S�a<��a<�a<r�a<�a<Z�a<Đa<&�a<��a<�a<�a<�a<}�a<��a<Y�a<֔a<I�a<ѕa<Z�a<ܖa<M�a<��a<A�a<ɘa<P�a<��a<-�a<��a<-�a<��a<�a<��a<�a<h�a<�a<h�a<ޞa<Z�a<��a<-�a<��a<�a<~�a<١a<0�a<��a<�a<V�a<��a<�a<D�a<��a<�a<>�a<��a<��a<�a<3�a<m�a<��a<�a<)�a<D�a<m�a<��a<ߧa<�a<�a<>�a<S�a<��a<��a<��a<��a<ިa<��a<�a<(�a<T�a<`�a<e�a<x�a<��a<��a<��a<��a<��a<ȩa<ѩa<Ωa<��a<��a<��a<��a<��a<��a<��a<z�a<o�a<\�a<K�a<G�a<4�a<�a<�a<ɨa<��a<��a<��a<G�a<#�a<�a<�a<��a<��a<L�a<%�a<�a<צa<��a<��a<A�a<�a<ߥa<��a<��a<H�a<��a<¤a<��a<S�a<�a<��a<s�a< �a<ݢa<��a<Q�a<��a<��a<D�a<�a<��a<F�a<�a<��a<�a<��a<Y�a<��a<��a<	�a<��a<7�a<ěa<I�a<Κa<P�a<�a<t�a<�a<��a<6�a<��a<C�a<Ֆa<t�a<��a<~�a<��a<��a<1�a<��a<>�a<��a<V�a<�a<��a<#�a<��a<<�a<ȏa<l�a<�a<��a<S�a<��a<��a<&�a<�a<��a<>�a<؋a<��a<0�a< �a<��a<i�a<�a<ۉa<��a<s�a<=�a<&�a<�a<��a<��a<��a<~�a<V�a<(�a<�a<�a<�a<��a<�a<ڇa<Շa<҇a<��a<��a<��a<�a<�a<�a<0�a<Y�a<�  �  ^�a<��a<��a<وa<�a<�a<W�a<r�a<ɉa<։a<)�a<K�a<��a<�a<!�a<��a<��a<�a<i�a<��a<?�a<q�a<�a<0�a<Îa<�a<�a<��a<C�a<̐a<�a<��a<
�a<~�a<�a<B�a<�a<K�a<��a<I�a<ܕa<M�a<ɖa<`�a<��a<a�a<��a<:�a<��a<B�a<��a<�a<��a<��a<��a<�a<��a<�a<K�a<�a<@�a<ɟa<K�a<��a<	�a<f�a<�a<,�a<��a<��a<F�a<��a<�a<f�a<��a<�a<	�a<e�a<��a<�a<T�a<Y�a<��a<٦a< �a<X�a<r�a<ŧa<��a<��a<�a<^�a<]�a<v�a<��a<��a<�a<�a<�a<'�a<�a<X�a<K�a<��a<{�a<��a<��a<��a<éa<��a<שa<��a<ʩa<��a<��a<ȩa<��a<��a<h�a<��a<w�a<~�a<h�a<=�a<H�a<�a<!�a<�a<ިa<Ȩa<��a<}�a<C�a<B�a<�a<�a<��a<��a<n�a<'�a<�a<Ŧa<��a<u�a<A�a<5�a<եa<��a<e�a<[�a<�a<Ϥa<��a<<�a<�a<��a<��a<(�a<ܢa<��a<�a<�a<��a<e�a<�a<��a<9�a<ڟa<��a<�a<Ӟa<K�a<�a<~�a<�a<��a<�a<̛a<.�a<�a<p�a<��a<��a<�a<��a<�a<a<a�a<Ζa<b�a<�a<��a<��a<��a<!�a<��a<I�a<��a<x�a<בa<��a<�a<��a<>�a<ʏa<��a<�a<��a<>�a<�a<��a<+�a<��a<q�a<1�a<΋a<��a<;�a<�a<��a<Q�a<D�a<�a<a<��a<3�a<*�a<߈a<߈a<��a<��a<[�a<X�a<F�a<�a<'�a<�a<��a<܇a<܇a<�a<̇a<߇a<��a<�a<�a<�a<#�a<"�a<Z�a<�  �  g�a<��a<��a<ψa<��a<+�a<Y�a<w�a<��a<݉a<*�a<o�a<��a<֊a<�a<h�a<��a<)�a<m�a<ǌa<"�a<�a<�a<D�a<��a<�a<~�a<ޏa<I�a<��a<)�a<��a<��a<��a<��a<o�a<��a<H�a<הa<N�a<ݕa<K�a<Ζa<E�a<Ɨa<E�a<Øa<N�a<��a<2�a<��a<�a<��a<�a<��a<��a<p�a<�a<k�a<�a<E�a<ɟa<3�a<��a<�a<r�a<ӡa<6�a<��a<��a<I�a<��a<�a<D�a<|�a<�a<+�a<x�a<¥a<�a<4�a<n�a<��a<ߦa<�a<P�a<w�a<��a<ϧa<�a< �a<?�a<g�a<|�a<��a<��a<ƨa<ܨa<��a<�a<D�a<S�a<P�a<}�a<z�a<��a<��a<��a<��a<��a<��a<��a<��a<ũa<��a<��a<��a<��a<��a<��a<~�a<e�a<X�a<S�a<8�a<!�a<�a<��a<Ԩa<��a<��a<~�a<H�a<3�a<��a<�a<§a<~�a<P�a<!�a<��a<Φa<��a<y�a<K�a<�a<�a<��a<y�a<C�a<�a<Τa<��a<B�a<��a<��a<q�a<�a<�a<��a<C�a<�a<��a<D�a<�a<��a<7�a<ߟa<x�a<�a<��a<R�a<��a<��a<�a<��a<!�a<ɛa<R�a<Қa<]�a<�a<y�a<�a<��a<!�a<��a<I�a<זa<s�a<�a<w�a<�a<��a<!�a<��a<F�a<a<U�a<Бa<��a<�a<��a<H�a<��a<l�a<�a<��a<D�a<�a<��a<0�a<ڌa<��a<B�a<ދa<��a<D�a<��a<��a<b�a<�a<ىa<��a<u�a<Y�a<%�a<�a<ֈa<��a<��a<s�a<P�a<6�a<%�a<�a<��a<�a<�a<Ӈa<ԇa<҇a<�a<�a<��a<��a<��a<�a<8�a<K�a<�  �  ��a<w�a<��a<Јa<��a</�a<P�a<��a<��a<�a<�a<\�a<��a<�a<B�a<u�a<Ӌa<�a<h�a<ߌa<�a<��a<ٍa<Q�a<��a<�a<~�a<ޏa<c�a<��a<2�a<��a<�a<n�a<�a<f�a<˓a<Y�a<ٔa<U�a<ȕa<G�a<�a<:�a<�a<>�a<͘a<<�a<��a</�a<��a<:�a<��a<&�a<��a<�a<��a<�a<z�a<͞a<`�a<˟a<'�a<��a<�a<��a<ϡa<S�a<��a<	�a<L�a<��a<��a<D�a<��a<ɤa<�a<`�a<��a<��a<0�a<{�a<��a<��a<�a<H�a<��a<��a<�a<�a<.�a<0�a<v�a<��a<��a<ɨa<Өa<�a<�a< �a<:�a<9�a<v�a<j�a<��a<��a<��a<��a<��a<ѩa<��a<کa<��a<��a<��a<��a<��a<��a<��a<p�a<u�a<u�a<\�a<V�a<&�a<=�a<��a<�a<ըa<��a<��a<u�a<V�a<�a<�a<ͧa<��a<��a<f�a<H�a<�a<�a<��a<u�a<c�a<	�a<�a<��a<��a<C�a<�a<Τa<��a<\�a<�a<ţa<k�a<.�a<̢a<}�a<:�a<աa<��a<F�a<�a<��a<3�a<��a<n�a<8�a<��a<\�a<�a<��a<�a<��a<D�a<��a<\�a<՚a<w�a<	�a<~�a<"�a<��a<<�a<×a<=�a<��a<Z�a<��a<s�a<"�a<��a<6�a<��a<+�a<̒a<V�a<�a<c�a<�a<��a<%�a<Տa<h�a<�a<��a<Y�a<�a<��a<C�a<ٌa<��a<&�a<�a<|�a<T�a<�a<��a<x�a<&�a<�a<��a<}�a<O�a<�a<
�a<Ĉa<��a<��a<s�a<X�a<4�a<8�a<��a<�a<߇a<�a<݇a<݇a<χa<��a<��a<·a<�a<�a<�a<;�a<9�a<�  �  d�a<��a<��a<҈a<�a<�a<M�a<��a<��a<��a<$�a<k�a<��a<�a<�a<|�a<Ëa<)�a<r�a<Ќa<&�a<��a<ԍa<O�a<��a<�a<��a<܏a<E�a<a<&�a<��a<�a<u�a<�a<W�a<ܓa<^�a<Ӕa<K�a<��a<F�a<Ȗa<C�a<՗a<H�a<ܘa<-�a<��a<<�a<��a</�a<��a< �a<��a<�a<��a<��a<n�a<�a<V�a<Ɵa<8�a<��a<��a<��a<ܡa<G�a<��a<�a<G�a<��a<�a<@�a<��a<פa<�a<h�a<��a<��a<"�a<o�a<��a<ܦa<�a<N�a<��a<��a<�a<�a<-�a<H�a<j�a<��a<��a<��a<ܨa<�a<�a<!�a<E�a<P�a<r�a<s�a<��a<��a<��a<ĩa<��a<��a<��a<��a<��a<ũa<��a<��a<��a<��a<��a<��a<y�a<k�a<D�a<P�a<9�a<�a<�a<��a<רa<Ψa<��a<s�a<_�a<+�a<�a<ާa<��a<��a<]�a<%�a<�a<զa<��a<~�a<S�a<�a<��a<��a<��a<V�a<�a<Фa<��a<>�a<	�a<��a<[�a<+�a<Ӣa<��a<+�a<�a<��a<@�a<�a<��a<2�a<ٟa<w�a<)�a<��a<k�a<םa<��a<�a<��a<:�a<ɛa<V�a<�a<m�a<��a<��a<�a<��a<2�a<��a<N�a<�a<M�a<�a<��a<�a<��a< �a<��a<H�a<��a<R�a<�a<r�a<��a<��a</�a<ҏa<Z�a<�a<��a<A�a<�a<��a<=�a<�a<��a<�a<�a<��a<G�a<��a<��a<g�a</�a<�a<��a<�a<Z�a<"�a<�a<̈a<��a<��a<]�a<h�a<;�a<'�a<�a<��a<�a<�a<Ǉa<҇a<ԇa<ևa<ɇa<�a<�a<�a< �a<5�a<L�a<�  �  Z�a<��a<��a<��a<�a<*�a<n�a<}�a<��a<�a<&�a<j�a<��a<�a<*�a<��a<��a<*�a<p�a<Ќa<*�a<��a<�a<H�a<��a<�a<�a<�a<8�a<��a<�a<��a<��a<g�a<�a<S�a<�a<9�a<֔a<@�a<Εa<A�a<Ɩa<[�a<˗a<.�a<��a<P�a<˙a<(�a<��a<#�a<��a<�a<��a<�a<��a<	�a<`�a<��a<J�a<џa<+�a<��a<�a<u�a<¡a<:�a<��a<�a<:�a<��a<ܣa<G�a<r�a<�a<�a<d�a<��a<ܥa<,�a<]�a<��a<ʦa<"�a<U�a<s�a<��a<اa<�a<!�a<C�a<m�a<��a<��a<��a<��a<�a<�a<�a<>�a<R�a<c�a<��a<}�a<��a<��a<��a<��a<��a<թa<��a<��a<��a<��a<��a<��a<��a<~�a<��a<]�a<g�a<N�a<B�a<7�a<�a<"�a<�a<Ǩa<��a<��a<��a<N�a<:�a<
�a<�a<��a<��a<|�a<0�a<+�a<ʦa<��a<}�a<S�a< �a<�a<Хa<~�a<0�a<��a<Ϥa<��a<1�a<�a<��a<e�a<�a<Ţa<��a<'�a<�a<w�a<C�a<ڠa<��a<-�a<ןa<��a<�a<��a<P�a<��a<��a<�a<��a<.�a<ћa<H�a<�a<v�a<��a<��a<�a<��a<&�a<ɗa<A�a<�a<t�a<�a<f�a<	�a<��a<�a<��a<9�a<��a<X�a<Ǒa<z�a<��a<��a<+�a<��a<d�a<��a<��a</�a<�a<��a<,�a<Ōa<��a<K�a<��a<��a<J�a<��a<��a<[�a<H�a<�a<ɉa<z�a<S�a<#�a<��a<܈a<��a<��a<u�a<C�a<&�a<�a<%�a<�a<�a<ۇa<ˇa<ԇa<��a<�a<Ƈa<�a<Շa<��a<	�a<'�a<J�a<�  �  i�a<{�a<��a<�a<��a</�a<Q�a<��a<ĉa<��a<�a<u�a<��a<��a<-�a<��a<ًa<(�a<p�a<�a<,�a<��a<�a<R�a<��a<(�a<d�a<ڏa<R�a<��a<'�a<��a<�a<j�a<ےa<N�a<ӓa<E�a<͔a<F�a<ȕa<I�a<Жa<,�a<ڗa<Q�a<Иa<C�a<ęa<:�a<ɚa<6�a<��a<-�a<��a<�a<��a<�a<�a<�a<^�a<ߟa<:�a<��a<�a<��a<ޡa<N�a<{�a<��a<E�a<��a<�a<;�a<��a<Фa<�a<Y�a<��a<�a<'�a<k�a<��a<�a<�a<4�a<��a<��a<�a<��a<$�a<G�a<��a<��a<��a<Ѩa<�a<�a<!�a</�a<O�a<H�a<q�a<��a<��a<��a<��a<��a<ȩa<��a<��a<��a<��a<��a<��a<��a<��a<��a<q�a<t�a<d�a<f�a<M�a<K�a<*�a<$�a<��a<�a<�a<��a<��a<v�a<X�a<=�a<�a<֧a<ȧa<��a<u�a<3�a<�a<�a<��a<}�a<e�a<"�a<�a<��a<��a<H�a<�a<��a<��a<K�a<�a<��a<d�a< �a<Ȣa<v�a<"�a<ݡa<��a<:�a<�a<��a<5�a<�a<`�a<.�a<Ğa<_�a<�a<��a<�a<��a<@�a<śa<c�a<�a<x�a<��a<��a<'�a<��a<:�a<חa<P�a<��a<d�a< �a<��a<�a<w�a<$�a<��a</�a<��a<M�a<ԑa<j�a<��a<��a<(�a<ŏa<_�a<�a<��a<G�a<�a<w�a<K�a<ߌa<��a<0�a<�a<��a<^�a<��a<��a<��a<:�a<��a<̉a<��a<d�a<�a<�a<�a<��a<��a<w�a<P�a<K�a<"�a<��a<��a<�a<݇a<̇a<҇a<��a<Ƈa<��a<҇a<܇a<��a<	�a<0�a<<�a<�  �  c�a<~�a<��a<Ԉa<��a<8�a<K�a<��a<��a<�a<3�a<|�a<��a<�a<C�a<r�a<Ջa<1�a<��a<ڌa<#�a<��a<Սa<b�a<��a<�a<y�a<܏a<D�a<��a<+�a<r�a<��a<d�a<�a<h�a<ɓa<W�a<��a<D�a<ҕa<1�a<Жa<:�a<ԗa<@�a<טa<=�a<͙a<M�a<��a<C�a<��a<1�a<��a<�a<��a<��a<��a<�a<j�a<ßa<C�a<��a<�a<��a<Ρa<F�a<��a<��a<1�a<��a<�a<�a<��a<¤a<#�a<b�a<��a<�a<�a<r�a<��a<צa<�a<F�a<��a<��a<�a<�a<B�a<E�a<n�a<��a<��a<̨a<Өa<�a<�a<)�a<T�a<Z�a<|�a<l�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ĩa<��a<��a<��a<��a<��a<{�a<o�a<R�a<?�a<T�a<�a<�a<�a<��a<ڨa<��a<��a<p�a<w�a<'�a<!�a<�a<ϧa<��a<\�a<J�a<�a<�a<¦a<��a<]�a<�a<�a<��a<��a<>�a<�a<ɤa<��a<=�a<�a<��a<L�a<�a<¢a<��a<<�a<ӡa<��a<�a<ޠa<��a<�a<�a<m�a<(�a<��a<f�a<�a<��a<*�a<��a<N�a<ћa<g�a<ޚa<v�a<�a<��a<(�a<��a<F�a<��a<Y�a<�a<_�a<
�a<s�a<�a<��a<#�a<��a<6�a<��a<1�a<�a<]�a<�a<��a<�a<Əa<H�a<�a<��a<;�a<�a<��a<<�a<Ԍa<��a<%�a<�a<��a<K�a<�a<Êa<{�a<'�a<�a<��a<��a<i�a<,�a<�a<ƈa<͈a<��a<y�a<W�a<8�a<(�a<��a<��a<чa<�a<��a<��a<̇a<Ça<݇a<هa<�a<�a<��a<9�a<.�a<�  �  U�a<��a<��a<Ԉa<��a<0�a<U�a<��a<��a<��a<0�a<h�a<��a<�a<H�a<��a<ԋa<+�a<y�a<�a<0�a<��a<��a<L�a<��a<�a<~�a<܏a<9�a<��a<�a<��a< �a<_�a<Вa<A�a<��a<A�a<Ԕa<;�a<Ǖa<@�a<Ėa<V�a<a<C�a<��a<H�a<��a<<�a<��a<7�a<��a<�a<��a<(�a<��a<�a<i�a<�a<^�a<ݟa<<�a<��a<�a<r�a<ӡa<5�a<��a<�a<@�a<��a<أa<=�a<|�a<��a<�a<I�a<��a<�a<(�a<M�a<��a<Ԧa<�a<T�a<y�a<��a<էa<��a<)�a<K�a<~�a<��a<��a<��a<�a<�a<*�a<>�a<=�a<^�a<t�a<}�a<��a<��a<��a<��a<��a<��a<ĩa<��a<��a<��a<��a<��a<��a<|�a<o�a<f�a<\�a<h�a<Q�a<1�a<0�a<�a<�a<�a<ڨa<��a<��a<z�a<\�a<8�a<�a<�a<��a<��a<��a<N�a<,�a<�a<��a<��a<f�a<&�a<�a<��a<��a<C�a<�a<Τa<��a<2�a<��a<��a<f�a<�a<��a<k�a<�a<ɡa<�a<A�a<ՠa<��a<,�a<՟a<��a<�a<��a<Q�a<�a<��a<�a<��a<B�a<՛a<P�a<�a<��a<�a<��a<�a<��a<:�a<՗a<R�a<ޖa<h�a<�a<x�a<�a<��a<�a<��a<2�a<��a<O�a<ёa<V�a<�a<}�a<�a<a<`�a<�a<��a<9�a<�a<��a<2�a<݌a<��a<0�a<�a<��a<[�a<�a<��a<m�a<T�a<�a<Չa<��a<S�a<0�a<�a<׈a<��a<��a<v�a<P�a<9�a<�a<�a<�a<�a<Їa<ʇa<Ӈa<��a<��a<��a<Ça<ԇa< �a<�a<�a<B�a<�  �  N�a<��a<��a<�a<��a<)�a<n�a<��a<҉a<�a<E�a<��a<��a<��a<�a<��a<Ћa<E�a<~�a<Ռa<9�a<��a<�a<?�a<��a<�a<g�a<ޏa<;�a<��a<�a<��a<ّa<s�a<�a<L�a<�a<-�a<͔a<5�a<��a<_�a<��a<D�a<��a<a�a<��a<U�a<șa<7�a<Κa<!�a<ԛa<#�a<��a<�a<|�a<�a<q�a<�a<N�a<�a<7�a<��a<%�a<i�a<�a<(�a<��a<ߢa<[�a<��a<ңa<<�a<`�a<�a<�a<^�a<��a<��a<,�a<J�a<��a<ߦa<�a<>�a<v�a<ça<ȧa<�a<$�a<P�a<z�a<��a<Шa<��a<�a<ۨa<!�a<5�a<P�a<z�a<^�a<��a<��a<��a<��a<��a<ʩa<��a<��a<��a<̩a<��a<��a<��a<��a<��a<u�a<��a<^�a<I�a<M�a<)�a<B�a<�a<
�a<٨a<�a<��a<��a<��a<R�a<K�a<�a<��a<էa<��a<y�a<�a<"�a<�a<צa<��a<Y�a</�a<�a<ӥa<t�a<U�a<	�a<��a<��a<4�a<�a<��a<l�a<��a<Ѣa<��a< �a<�a<j�a<;�a<Ϡa<��a<K�a<Ɵa<x�a<�a<Ԟa<I�a<��a<��a<�a<a<+�a<��a<Y�a<��a<t�a<��a<��a<�a<Ԙa<*�a<ڗa<M�a<�a<~�a<�a<��a<��a<��a<�a<��a<.�a<��a<M�a<��a<|�a<��a<��a<4�a<��a<e�a<�a<��a<D�a<�a<��a</�a<��a<{�a<O�a<�a<��a<W�a<��a<ߊa<n�a<F�a<؉a<̉a<��a<e�a<L�a<�a<�a<��a<��a<t�a<O�a<M�a<�a<	�a<߇a<��a<Ǉa<Ƈa<��a<��a<هa<��a<�a<ևa<�a<	�a<�a<U�a<�  �  S�a<��a<��a<ֈa<�a<%�a<f�a<��a<ωa<��a<4�a<t�a<��a<�a<S�a<��a<؋a<*�a<~�a<׌a<A�a<��a<�a<B�a<��a<�a<��a<�a<6�a<��a<�a<��a<�a<[�a<Œa<>�a<��a<G�a<��a<M�a<��a<>�a<��a<S�a<їa<K�a<��a<?�a<әa<K�a<ƚa<4�a<��a<&�a<��a<9�a<��a<�a<z�a<�a<]�a<ٟa<I�a<��a<�a<k�a<ڡa<C�a<��a<�a<;�a<|�a<�a<.�a<|�a<��a<��a<=�a<��a<եa<%�a<c�a<��a<Цa<�a<Y�a<~�a<��a<ϧa<�a<9�a<[�a<r�a<��a<��a<ͨa< �a<�a<9�a<8�a<F�a<`�a<o�a<��a<��a<��a<��a<��a<��a<ĩa<Ʃa<��a<��a<��a<��a<��a<��a<x�a<s�a<b�a<c�a<K�a<U�a<7�a<!�a<�a<�a<��a<ܨa<��a<��a<��a<m�a<H�a<�a<�a<ȧa<��a<��a<Y�a<4�a<�a<��a<��a<Z�a<7�a<�a<¥a<w�a<4�a<	�a<פa<��a</�a<�a<��a<f�a<�a<��a<`�a<�a<��a<��a<(�a<�a<t�a<*�a<Οa<��a<%�a<��a<G�a<�a<��a<(�a<��a<?�a<՛a<\�a<��a<��a<&�a<��a<"�a<��a<8�a<їa<_�a<�a<i�a<�a<�a<�a<��a<�a<��a<�a<��a<?�a<Бa<P�a<ߐa<p�a<�a<��a<]�a<��a<��a<4�a<�a<��a<7�a<Ԍa<��a<=�a<��a<��a<O�a<��a<��a<|�a<S�a<�a<�a<��a<[�a<1�a<�a<�a<Èa<��a<l�a<D�a<<�a<+�a<�a<�a<ۇa<̇a<Շa<��a<��a<��a<��a<��a<ۇa<�a<�a<�a<4�a<�  �  i�a<j�a<��a<̈a<�a<E�a<P�a<��a<��a<�a</�a<{�a<Ɋa<�a<#�a<��a<�a<(�a<��a<�a<3�a<��a<ٍa<r�a<��a<�a<n�a<��a<L�a<��a<�a<k�a<��a<\�a<��a<w�a<��a<c�a<��a<H�a<��a<H�a<Ɩa</�a<×a<>�a<�a<L�a<əa<=�a<��a<X�a<��a<@�a<��a<�a<y�a<
�a<��a<�a<��a<֟a<@�a<��a<�a<��a<ϡa<5�a<{�a<�a<K�a<��a<�a<	�a<��a<��a</�a<d�a<��a<�a<��a<_�a<��a<�a<��a<<�a<z�a<��a<��a<�a<*�a<Q�a<�a<��a<��a<�a<�a<�a<	�a<K�a<V�a<V�a<��a<u�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<m�a<��a<`�a<k�a<P�a<>�a<7�a<-�a<$�a<�a<�a<Ѩa<ƨa<��a<v�a<`�a<2�a<2�a<�a<ϧa<��a<]�a<*�a<�a<�a<��a<��a<l�a<)�a<�a<��a<��a<C�a<�a<��a<g�a<E�a<�a<��a<E�a<�a<��a<z�a<K�a<��a<��a<�a<�a<{�a<3�a<֟a<c�a<�a<��a<w�a<��a<��a<�a<��a<c�a<Ǜa<w�a<��a<i�a<�a<��a<<�a<��a<]�a<Ηa<V�a<�a<l�a<�a<t�a<�a<x�a<�a<��a< �a<��a<�a<�a<F�a<�a<��a<�a<Ώa<7�a<��a<��a<I�a<͍a<�a<3�a<ٌa<��a<(�a<�a<��a<\�a<�a<��a<��a<;�a<�a<��a<��a<k�a<(�a<#�a<ψa<��a<��a<��a<e�a</�a<�a<�a<��a<އa<̇a<ȇa<��a<χa<��a<�a<��a<�a<�a<��a<�a<@�a<�  �  S�a<��a<��a<ֈa<�a<%�a<f�a<��a<ωa<��a<4�a<t�a<��a<�a<S�a<��a<؋a<*�a<~�a<׌a<A�a<��a<�a<B�a<��a<�a<��a<�a<6�a<��a<�a<��a<�a<[�a<Œa<>�a<��a<G�a<��a<M�a<��a<>�a<��a<S�a<їa<K�a<��a<?�a<әa<K�a<ƚa<4�a<��a<&�a<��a<9�a<��a<�a<z�a<�a<]�a<ٟa<I�a<��a<�a<k�a<ڡa<C�a<��a<�a<;�a<|�a<�a<.�a<|�a<��a<��a<=�a<��a<եa<%�a<c�a<��a<Цa<�a<Y�a<~�a<��a<ϧa<�a<9�a<[�a<r�a<��a<��a<ͨa< �a<�a<9�a<8�a<F�a<`�a<o�a<��a<��a<��a<��a<��a<��a<ĩa<Ʃa<��a<��a<��a<��a<��a<��a<x�a<s�a<b�a<c�a<K�a<U�a<7�a<!�a<�a<�a<��a<ܨa<��a<��a<��a<m�a<H�a<�a<�a<ȧa<��a<��a<Y�a<4�a<�a<��a<��a<Z�a<7�a<�a<¥a<w�a<4�a<	�a<פa<��a</�a<�a<��a<f�a<�a<��a<`�a<�a<��a<��a<(�a<�a<t�a<*�a<Οa<��a<%�a<��a<G�a<�a<��a<(�a<��a<?�a<՛a<\�a<��a<��a<&�a<��a<"�a<��a<8�a<їa<_�a<�a<i�a<�a<�a<�a<��a<�a<��a<�a<��a<?�a<Бa<P�a<ߐa<p�a<�a<��a<]�a<��a<��a<4�a<�a<��a<7�a<Ԍa<��a<=�a<��a<��a<O�a<��a<��a<|�a<S�a<�a<�a<��a<[�a<1�a<�a<�a<Èa<��a<l�a<D�a<<�a<+�a<�a<�a<ۇa<̇a<Շa<��a<��a<��a<��a<��a<ۇa<�a<�a<�a<4�a<�  �  N�a<��a<��a<�a<��a<)�a<n�a<��a<҉a<�a<E�a<��a<��a<��a<�a<��a<Ћa<E�a<~�a<Ռa<9�a<��a<�a<?�a<��a<�a<g�a<ޏa<;�a<��a<�a<��a<ّa<s�a<�a<L�a<�a<-�a<͔a<5�a<��a<_�a<��a<D�a<��a<a�a<��a<U�a<șa<7�a<Κa<!�a<ԛa<#�a<��a<�a<|�a<�a<q�a<�a<N�a<�a<7�a<��a<%�a<i�a<�a<(�a<��a<ߢa<[�a<��a<ңa<<�a<`�a<�a<�a<^�a<��a<��a<,�a<J�a<��a<ߦa<�a<>�a<v�a<ça<ȧa<�a<$�a<P�a<z�a<��a<Шa<��a<�a<ۨa<!�a<5�a<P�a<z�a<^�a<��a<��a<��a<��a<��a<ʩa<��a<��a<��a<̩a<��a<��a<��a<��a<��a<u�a<��a<^�a<I�a<M�a<)�a<B�a<�a<
�a<٨a<�a<��a<��a<��a<R�a<K�a<�a<��a<էa<��a<y�a<�a<"�a<�a<צa<��a<Y�a</�a<�a<ӥa<t�a<U�a<	�a<��a<��a<4�a<�a<��a<l�a<��a<Ѣa<��a< �a<�a<j�a<;�a<Ϡa<��a<K�a<Ɵa<x�a<�a<Ԟa<I�a<��a<��a<�a<a<+�a<��a<Y�a<��a<t�a<��a<��a<�a<Ԙa<*�a<ڗa<M�a<�a<~�a<�a<��a<��a<��a<�a<��a<.�a<��a<M�a<��a<|�a<��a<��a<4�a<��a<e�a<�a<��a<D�a<�a<��a</�a<��a<{�a<O�a<�a<��a<W�a<��a<ߊa<n�a<F�a<؉a<̉a<��a<e�a<L�a<�a<�a<��a<��a<t�a<O�a<M�a<�a<	�a<߇a<��a<Ǉa<Ƈa<��a<��a<هa<��a<�a<ևa<�a<	�a<�a<U�a<�  �  U�a<��a<��a<Ԉa<��a<0�a<U�a<��a<��a<��a<0�a<h�a<��a<�a<H�a<��a<ԋa<+�a<y�a<�a<0�a<��a<��a<L�a<��a<�a<~�a<܏a<9�a<��a<�a<��a< �a<_�a<Вa<A�a<��a<A�a<Ԕa<;�a<Ǖa<@�a<Ėa<V�a<a<C�a<��a<H�a<��a<<�a<��a<7�a<��a<�a<��a<(�a<��a<�a<i�a<�a<^�a<ݟa<<�a<��a<�a<r�a<ӡa<5�a<��a<�a<@�a<��a<أa<=�a<|�a<��a<�a<I�a<��a<�a<(�a<M�a<��a<Ԧa<�a<T�a<y�a<��a<էa<��a<)�a<K�a<~�a<��a<��a<��a<�a<�a<*�a<>�a<=�a<^�a<t�a<}�a<��a<��a<��a<��a<��a<��a<ĩa<��a<��a<��a<��a<��a<��a<|�a<o�a<f�a<\�a<h�a<Q�a<1�a<0�a<�a<�a<�a<ڨa<��a<��a<z�a<\�a<8�a<�a<�a<��a<��a<��a<N�a<,�a<�a<��a<��a<f�a<&�a<�a<��a<��a<C�a<�a<Τa<��a<2�a<��a<��a<f�a<�a<��a<k�a<�a<ɡa<�a<A�a<ՠa<��a<,�a<՟a<��a<�a<��a<Q�a<�a<��a<�a<��a<B�a<՛a<P�a<�a<��a<�a<��a<�a<��a<:�a<՗a<R�a<ޖa<h�a<�a<x�a<�a<��a<�a<��a<2�a<��a<O�a<ёa<V�a<�a<}�a<�a<a<`�a<�a<��a<9�a<�a<��a<2�a<݌a<��a<0�a<�a<��a<[�a<�a<��a<m�a<T�a<�a<Չa<��a<S�a<0�a<�a<׈a<��a<��a<v�a<P�a<9�a<�a<�a<�a<�a<Їa<ʇa<Ӈa<��a<��a<��a<Ça<ԇa< �a<�a<�a<B�a<�  �  c�a<~�a<��a<Ԉa<��a<8�a<K�a<��a<��a<�a<3�a<|�a<��a<�a<C�a<r�a<Ջa<1�a<��a<ڌa<#�a<��a<Սa<b�a<��a<�a<y�a<܏a<D�a<��a<+�a<r�a<��a<d�a<�a<h�a<ɓa<W�a<��a<D�a<ҕa<1�a<Жa<:�a<ԗa<@�a<טa<=�a<͙a<M�a<��a<C�a<��a<1�a<��a<�a<��a<��a<��a<�a<j�a<ßa<C�a<��a<�a<��a<Ρa<F�a<��a<��a<1�a<��a<�a<�a<��a<¤a<#�a<b�a<��a<�a<�a<r�a<��a<צa<�a<F�a<��a<��a<�a<�a<B�a<E�a<n�a<��a<��a<̨a<Өa<�a<�a<)�a<T�a<Z�a<|�a<l�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ĩa<��a<��a<��a<��a<��a<{�a<o�a<R�a<?�a<T�a<�a<�a<�a<��a<ڨa<��a<��a<p�a<w�a<'�a<!�a<�a<ϧa<��a<\�a<J�a<�a<�a<¦a<��a<]�a<�a<�a<��a<��a<>�a<�a<ɤa<��a<=�a<�a<��a<L�a<�a<¢a<��a<<�a<ӡa<��a<�a<ޠa<��a<�a<�a<m�a<(�a<��a<f�a<�a<��a<*�a<��a<N�a<ћa<g�a<ޚa<v�a<�a<��a<(�a<��a<F�a<��a<Y�a<�a<_�a<
�a<s�a<�a<��a<#�a<��a<6�a<��a<1�a<�a<]�a<�a<��a<�a<Əa<H�a<�a<��a<;�a<�a<��a<<�a<Ԍa<��a<%�a<�a<��a<K�a<�a<Êa<{�a<'�a<�a<��a<��a<i�a<,�a<�a<ƈa<͈a<��a<y�a<W�a<8�a<(�a<��a<��a<чa<�a<��a<��a<̇a<Ça<݇a<هa<�a<�a<��a<9�a<.�a<�  �  i�a<{�a<��a<�a<��a</�a<Q�a<��a<ĉa<��a<�a<u�a<��a<��a<-�a<��a<ًa<(�a<p�a<�a<,�a<��a<�a<R�a<��a<(�a<d�a<ڏa<R�a<��a<'�a<��a<�a<j�a<ےa<N�a<ӓa<E�a<͔a<F�a<ȕa<I�a<Жa<,�a<ڗa<Q�a<Иa<C�a<ęa<:�a<ɚa<6�a<��a<-�a<��a<�a<��a<�a<�a<�a<^�a<ߟa<:�a<��a<�a<��a<ޡa<N�a<{�a<��a<E�a<��a<�a<;�a<��a<Фa<�a<Y�a<��a<�a<'�a<k�a<��a<�a<�a<4�a<��a<��a<�a<��a<$�a<G�a<��a<��a<��a<Ѩa<�a<�a<!�a</�a<O�a<H�a<q�a<��a<��a<��a<��a<��a<ȩa<��a<��a<��a<��a<��a<��a<��a<��a<��a<q�a<t�a<d�a<f�a<M�a<K�a<*�a<$�a<��a<�a<�a<��a<��a<v�a<X�a<=�a<�a<֧a<ȧa<��a<u�a<3�a<�a<�a<��a<}�a<e�a<"�a<�a<��a<��a<H�a<�a<��a<��a<K�a<�a<��a<d�a< �a<Ȣa<v�a<"�a<ݡa<��a<:�a<�a<��a<5�a<�a<`�a<.�a<Ğa<_�a<�a<��a<�a<��a<@�a<śa<c�a<�a<x�a<��a<��a<'�a<��a<:�a<חa<P�a<��a<d�a< �a<��a<�a<w�a<$�a<��a</�a<��a<M�a<ԑa<j�a<��a<��a<(�a<ŏa<_�a<�a<��a<G�a<�a<w�a<K�a<ߌa<��a<0�a<�a<��a<^�a<��a<��a<��a<:�a<��a<̉a<��a<d�a<�a<�a<�a<��a<��a<w�a<P�a<K�a<"�a<��a<��a<�a<݇a<̇a<҇a<��a<Ƈa<��a<҇a<܇a<��a<	�a<0�a<<�a<�  �  Z�a<��a<��a<��a<�a<*�a<n�a<}�a<��a<�a<&�a<j�a<��a<�a<*�a<��a<��a<*�a<p�a<Ќa<*�a<��a<�a<H�a<��a<�a<�a<�a<8�a<��a<�a<��a<��a<g�a<�a<S�a<�a<9�a<֔a<@�a<Εa<A�a<Ɩa<[�a<˗a<.�a<��a<P�a<˙a<(�a<��a<#�a<��a<�a<��a<�a<��a<	�a<`�a<��a<J�a<џa<+�a<��a<�a<u�a<¡a<:�a<��a<�a<:�a<��a<ܣa<G�a<r�a<�a<�a<d�a<��a<ܥa<,�a<]�a<��a<ʦa<"�a<U�a<s�a<��a<اa<�a<!�a<C�a<m�a<��a<��a<��a<��a<�a<�a<�a<>�a<R�a<c�a<��a<}�a<��a<��a<��a<��a<��a<թa<��a<��a<��a<��a<��a<��a<��a<~�a<��a<]�a<g�a<N�a<B�a<7�a<�a<"�a<�a<Ǩa<��a<��a<��a<N�a<:�a<
�a<�a<��a<��a<|�a<0�a<+�a<ʦa<��a<}�a<S�a< �a<�a<Хa<~�a<0�a<��a<Ϥa<��a<1�a<�a<��a<e�a<�a<Ţa<��a<'�a<�a<w�a<C�a<ڠa<��a<-�a<ןa<��a<�a<��a<P�a<��a<��a<�a<��a<.�a<ћa<H�a<�a<v�a<��a<��a<�a<��a<&�a<ɗa<A�a<�a<t�a<�a<f�a<	�a<��a<�a<��a<9�a<��a<X�a<Ǒa<z�a<��a<��a<+�a<��a<d�a<��a<��a</�a<�a<��a<,�a<Ōa<��a<K�a<��a<��a<J�a<��a<��a<[�a<H�a<�a<ɉa<z�a<S�a<#�a<��a<܈a<��a<��a<u�a<C�a<&�a<�a<%�a<�a<�a<ۇa<ˇa<ԇa<��a<�a<Ƈa<�a<Շa<��a<	�a<'�a<J�a<�  �  d�a<��a<��a<҈a<�a<�a<M�a<��a<��a<��a<$�a<k�a<��a<�a<�a<|�a<Ëa<)�a<r�a<Ќa<&�a<��a<ԍa<O�a<��a<�a<��a<܏a<E�a<a<&�a<��a<�a<u�a<�a<W�a<ܓa<^�a<Ӕa<K�a<��a<F�a<Ȗa<C�a<՗a<H�a<ܘa<-�a<��a<<�a<��a</�a<��a< �a<��a<�a<��a<��a<n�a<�a<V�a<Ɵa<8�a<��a<��a<��a<ܡa<G�a<��a<�a<G�a<��a<�a<@�a<��a<פa<�a<h�a<��a<��a<"�a<o�a<��a<ܦa<�a<N�a<��a<��a<�a<�a<-�a<H�a<j�a<��a<��a<��a<ܨa<�a<�a<!�a<E�a<P�a<r�a<s�a<��a<��a<��a<ĩa<��a<��a<��a<��a<��a<ũa<��a<��a<��a<��a<��a<��a<y�a<k�a<D�a<P�a<9�a<�a<�a<��a<רa<Ψa<��a<s�a<_�a<+�a<�a<ާa<��a<��a<]�a<%�a<�a<զa<��a<~�a<S�a<�a<��a<��a<��a<V�a<�a<Фa<��a<>�a<	�a<��a<[�a<+�a<Ӣa<��a<+�a<�a<��a<@�a<�a<��a<2�a<ٟa<w�a<)�a<��a<k�a<םa<��a<�a<��a<:�a<ɛa<V�a<�a<m�a<��a<��a<�a<��a<2�a<��a<N�a<�a<M�a<�a<��a<�a<��a< �a<��a<H�a<��a<R�a<�a<r�a<��a<��a</�a<ҏa<Z�a<�a<��a<A�a<�a<��a<=�a<�a<��a<�a<�a<��a<G�a<��a<��a<g�a</�a<�a<��a<�a<Z�a<"�a<�a<̈a<��a<��a<]�a<h�a<;�a<'�a<�a<��a<�a<�a<Ǉa<҇a<ԇa<ևa<ɇa<�a<�a<�a< �a<5�a<L�a<�  �  ��a<w�a<��a<Јa<��a</�a<P�a<��a<��a<�a<�a<\�a<��a<�a<B�a<u�a<Ӌa<�a<h�a<ߌa<�a<��a<ٍa<Q�a<��a<�a<~�a<ޏa<c�a<��a<2�a<��a<�a<n�a<�a<f�a<˓a<Y�a<ٔa<U�a<ȕa<G�a<�a<:�a<�a<>�a<͘a<<�a<��a</�a<��a<:�a<��a<&�a<��a<�a<��a<�a<z�a<͞a<`�a<˟a<'�a<��a<�a<��a<ϡa<S�a<��a<	�a<L�a<��a<��a<D�a<��a<ɤa<�a<`�a<��a<��a<0�a<{�a<��a<��a<�a<H�a<��a<��a<�a<�a<.�a<0�a<v�a<��a<��a<ɨa<Өa<�a<�a< �a<:�a<9�a<v�a<j�a<��a<��a<��a<��a<��a<ѩa<��a<کa<��a<��a<��a<��a<��a<��a<��a<p�a<u�a<u�a<\�a<V�a<&�a<=�a<��a<�a<ըa<��a<��a<u�a<V�a<�a<�a<ͧa<��a<��a<f�a<H�a<�a<�a<��a<u�a<c�a<	�a<�a<��a<��a<C�a<�a<Τa<��a<\�a<�a<ţa<k�a<.�a<̢a<}�a<:�a<աa<��a<F�a<�a<��a<3�a<��a<n�a<8�a<��a<\�a<�a<��a<�a<��a<D�a<��a<\�a<՚a<w�a<	�a<~�a<"�a<��a<<�a<×a<=�a<��a<Z�a<��a<s�a<"�a<��a<6�a<��a<+�a<̒a<V�a<�a<c�a<�a<��a<%�a<Տa<h�a<�a<��a<Y�a<�a<��a<C�a<ٌa<��a<&�a<�a<|�a<T�a<�a<��a<x�a<&�a<�a<��a<}�a<O�a<�a<
�a<Ĉa<��a<��a<s�a<X�a<4�a<8�a<��a<�a<߇a<�a<݇a<݇a<χa<��a<��a<·a<�a<�a<�a<;�a<9�a<�  �  g�a<��a<��a<ψa<��a<+�a<Y�a<w�a<��a<݉a<*�a<o�a<��a<֊a<�a<h�a<��a<)�a<m�a<ǌa<"�a<�a<�a<D�a<��a<�a<~�a<ޏa<I�a<��a<)�a<��a<��a<��a<��a<o�a<��a<H�a<הa<N�a<ݕa<K�a<Ζa<E�a<Ɨa<E�a<Øa<N�a<��a<2�a<��a<�a<��a<�a<��a<��a<p�a<�a<k�a<�a<E�a<ɟa<3�a<��a<�a<r�a<ӡa<6�a<��a<��a<I�a<��a<�a<D�a<|�a<�a<+�a<x�a<¥a<�a<4�a<n�a<��a<ߦa<�a<P�a<w�a<��a<ϧa<�a< �a<?�a<g�a<|�a<��a<��a<ƨa<ܨa<��a<�a<D�a<S�a<P�a<}�a<z�a<��a<��a<��a<��a<��a<��a<��a<��a<ũa<��a<��a<��a<��a<��a<��a<~�a<e�a<X�a<S�a<8�a<!�a<�a<��a<Ԩa<��a<��a<~�a<H�a<3�a<��a<�a<§a<~�a<P�a<!�a<��a<Φa<��a<y�a<K�a<�a<�a<��a<y�a<C�a<�a<Τa<��a<B�a<��a<��a<q�a<�a<�a<��a<C�a<�a<��a<D�a<�a<��a<7�a<ߟa<x�a<�a<��a<R�a<��a<��a<�a<��a<!�a<ɛa<R�a<Қa<]�a<�a<y�a<�a<��a<!�a<��a<I�a<זa<s�a<�a<w�a<�a<��a<!�a<��a<F�a<a<U�a<Бa<��a<�a<��a<H�a<��a<l�a<�a<��a<D�a<�a<��a<0�a<ڌa<��a<B�a<ދa<��a<D�a<��a<��a<b�a<�a<ىa<��a<u�a<Y�a<%�a<�a<ֈa<��a<��a<s�a<P�a<6�a<%�a<�a<��a<�a<�a<Ӈa<ԇa<҇a<�a<�a<��a<��a<��a<�a<8�a<K�a<�  �  ^�a<��a<��a<وa<�a<�a<W�a<r�a<ɉa<։a<)�a<K�a<��a<�a<!�a<��a<��a<�a<i�a<��a<?�a<q�a<�a<0�a<Îa<�a<�a<��a<C�a<̐a<�a<��a<
�a<~�a<�a<B�a<�a<K�a<��a<I�a<ܕa<M�a<ɖa<`�a<��a<a�a<��a<:�a<��a<B�a<��a<�a<��a<��a<��a<�a<��a<�a<K�a<�a<@�a<ɟa<K�a<��a<	�a<f�a<�a<,�a<��a<��a<F�a<��a<�a<f�a<��a<�a<	�a<e�a<��a<�a<T�a<Y�a<��a<٦a< �a<X�a<r�a<ŧa<��a<��a<�a<^�a<]�a<v�a<��a<��a<�a<�a<�a<'�a<�a<X�a<K�a<��a<{�a<��a<��a<��a<éa<��a<שa<��a<ʩa<��a<��a<ȩa<��a<��a<h�a<��a<w�a<~�a<h�a<=�a<H�a<�a<!�a<�a<ިa<Ȩa<��a<}�a<C�a<B�a<�a<�a<��a<��a<n�a<'�a<�a<Ŧa<��a<u�a<A�a<5�a<եa<��a<e�a<[�a<�a<Ϥa<��a<<�a<�a<��a<��a<(�a<ܢa<��a<�a<�a<��a<e�a<�a<��a<9�a<ڟa<��a<�a<Ӟa<K�a<�a<~�a<�a<��a<�a<̛a<.�a<�a<p�a<��a<��a<�a<��a<�a<a<a�a<Ζa<b�a<�a<��a<��a<��a<!�a<��a<I�a<��a<x�a<בa<��a<�a<��a<>�a<ʏa<��a<�a<��a<>�a<�a<��a<+�a<��a<q�a<1�a<΋a<��a<;�a<�a<��a<Q�a<D�a<�a<a<��a<3�a<*�a<߈a<߈a<��a<��a<[�a<X�a<F�a<�a<'�a<�a<��a<܇a<܇a<�a<̇a<߇a<��a<�a<�a<�a<#�a<"�a<Z�a<�  �  y�a<��a<��a<Ĉa< �a<4�a<_�a<u�a<��a<�a<+�a<Q�a<��a<ӊa<�a<d�a<ŋa<�a<{�a<��a<�a<z�a<�a<S�a<��a<�a<r�a<�a<Z�a<Đa<&�a<��a<�a<�a<�a<}�a<��a<Y�a<֔a<I�a<ѕa<Z�a<ܖa<M�a<��a<A�a<ɘa<P�a<��a<-�a<��a<-�a<��a<�a<��a<�a<h�a<�a<h�a<ޞa<Z�a<��a<-�a<��a<�a<~�a<١a<0�a<��a<�a<V�a<��a<�a<D�a<��a<�a<>�a<��a<��a<�a<3�a<m�a<��a<�a<)�a<D�a<m�a<��a<ߧa<�a<�a<>�a<S�a<��a<��a<��a<��a<ިa<��a<�a<(�a<T�a<`�a<e�a<x�a<��a<��a<��a<��a<��a<ȩa<ѩa<Ωa<��a<��a<��a<��a<��a<��a<��a<z�a<o�a<\�a<K�a<G�a<4�a<�a<�a<ɨa<��a<��a<��a<G�a<#�a<�a<�a<��a<��a<L�a<%�a<�a<צa<��a<��a<A�a<�a<ߥa<��a<��a<H�a<��a<¤a<��a<S�a<�a<��a<s�a< �a<ݢa<��a<Q�a<��a<��a<D�a<�a<��a<F�a<�a<��a<�a<��a<Y�a<��a<��a<	�a<��a<7�a<ěa<I�a<Κa<P�a<�a<t�a<�a<��a<6�a<��a<C�a<Ֆa<t�a<��a<~�a<��a<��a<1�a<��a<>�a<��a<V�a<�a<��a<#�a<��a<<�a<ȏa<l�a<�a<��a<S�a<��a<��a<&�a<�a<��a<>�a<؋a<��a<0�a< �a<��a<i�a<�a<ۉa<��a<s�a<=�a<&�a<�a<��a<��a<��a<~�a<V�a<(�a<�a<�a<�a<��a<�a<ڇa<Շa<҇a<��a<��a<��a<�a<�a<�a<0�a<Y�a<�  �  L�a<n�a<��a<ȇa<��a<!�a</�a<��a<��a<׈a<
�a<@�a<��a<��a<<�a<M�a<��a<�a<i�a<��a<"�a<��a<ǌa<T�a<��a<�a<o�a<Ԏa<F�a<Əa<9�a<��a<0�a<��a<�a<o�a<�a<x�a<�a<^�a<��a<Z�a<ѕa<`�a<�a<`�a<�a<\�a<՘a<t�a<͙a<Q�a<��a<B�a<��a</�a<��a<�a<��a<�a<��a<��a<��a<ڟa<>�a<Ơa<�a<��a<ʡa<�a<~�a<�a</�a<��a<�a<�a<a�a<��a<��a<P�a<c�a<��a<�a<�a<A�a<~�a<Ħa<�a<�a<"�a<b�a<��a<��a<ħa<��a<��a<�a<<�a<.�a<D�a<c�a<o�a<��a<��a<Шa<��a<ڨa<��a<�a<��a<�a<�a<�a<�a<٨a<��a<�a<˨a<��a<��a<Ȩa<��a<~�a<��a<h�a<J�a<4�a<*�a<�a<��a<اa<��a<��a<Z�a<3�a<�a<Ӧa<��a<w�a<��a<�a<�a<��a<��a<y�a<Q�a<$�a<Τa<��a<��a<F�a<��a<��a<r�a<@�a<��a<��a<|�a<�a<��a<m�a<�a<ܠa<��a<�a<ڟa<d�a<��a<��a<]�a<�a<��a<�a<��a<[�a<ɛa<a�a<Ța<x�a<�a<��a< �a<��a<<�a<��a<Y�a<Ֆa<��a<��a<x�a<"�a<��a<-�a<��a<�a<��a<R�a<ґa<h�a<�a<��a<�a<��a<F�a<�a<a�a<�a<��a<>�a<֌a<��a<>�a<�a<��a<�a<��a<��a<1�a<��a<�a<g�a< �a<��a<��a<^�a<4�a<��a<�a<��a<��a<h�a<^�a<W�a<)�a<�a<��a<ކa<نa<�a<��a<݆a<نa<��a<��a<φa<��a<�a<��a<3�a<6�a<�  �  j�a<��a<��a<ʇa<݇a<�a<M�a<f�a<��a<шa<�a<H�a<��a<��a<�a<K�a<��a<�a<b�a<��a<�a<p�a<�a<>�a<��a<�a<��a<��a<_�a<Ǐa<,�a<��a<�a<w�a<�a<��a<��a<W�a<��a<m�a<�a<r�a< �a<w�a<�a<_�a<חa<a�a<Әa<F�a<��a<M�a<��a<9�a<��a<�a<��a<�a<��a<�a<��a<�a<Z�a<Οa<M�a<��a<�a<w�a<�a<N�a<��a<�a<9�a<��a<��a<$�a<w�a<��a<�a<+�a<��a<��a<�a<3�a<r�a<��a<��a<ܦa<�a<B�a<L�a<p�a<��a<��a<ǧa<�a<�a<�a<"�a<Q�a<c�a<~�a<��a<��a<��a<Ϩa<Өa<بa<�a<�a<�a<	�a<��a<��a<��a<�a<ɨa<�a<�a<٨a<��a<��a<��a<��a<r�a<i�a<S�a<*�a<�a<ߧa<ŧa<��a<x�a<T�a<-�a<�a<ۦa<��a<q�a<K�a<�a<�a<ϥa<��a<m�a<D�a<�a<�a<��a<l�a<C�a<�a<أa<��a<A�a<�a<��a<Y�a<�a<֡a<��a<0�a<��a<��a<*�a<ןa<}�a<-�a<Şa<R�a<�a<y�a<�a<��a<.�a<��a<]�a<�a<p�a<��a<y�a<�a<��a<,�a<��a<O�a<Öa<W�a<�a<��a< �a<��a< �a<��a<Q�a<Вa<V�a<ܑa<t�a<��a<��a<'�a<��a<4�a<Ўa<~�a<�a<��a<[�a<�a<��a<7�a<Ћa<{�a<8�a<ʊa<{�a<$�a<�a<��a<T�a< �a<ňa<��a<k�a<4�a<�a<߇a<��a<��a<�a<W�a<7�a<+�a<�a<�a<��a<�a<چa<҆a<φa<��a<߆a<�a<�a<Іa<��a<�a<%�a<A�a<�  �  P�a<v�a<��a<߇a<�a<�a<Y�a<j�a<��a<Ɉa<�a<=�a<��a<։a<�a<s�a<��a<�a<S�a<��a<4�a<t�a<��a<8�a<��a<#�a<v�a<��a<E�a<��a< �a<��a<�a<��a<�a<\�a<��a<]�a<�a<d�a<�a<]�a<ߕa<a�a<�a<��a<՗a<i�a<ߘa<[�a<�a<=�a<Śa<!�a<��a<+�a<��a<'�a<z�a<�a<r�a< �a<s�a<ԟa<T�a<��a<-�a<{�a<ҡa<,�a<��a<ޢa<+�a<��a<ƣa<'�a<O�a<��a<�a<0�a<��a<��a<�a<�a<S�a<��a<Ħa<�a<�a<K�a<O�a<��a<��a<��a<Чa<קa<�a<�a<8�a<Q�a<P�a<z�a<��a<èa<��a<ݨa<Ԩa<�a<�a<�a<�a<�a<�a<�a<��a<��a<̨a<�a<��a<˨a<��a<��a<��a<z�a<o�a<N�a<<�a<�a<'�a<�a<ħa<��a<}�a<y�a<%�a<�a<Цa<��a<��a<R�a<>�a<��a<ҥa<��a<r�a<d�a<�a< �a<��a<��a<N�a<��a<��a<p�a<:�a<�a<��a<^�a<�a<ǡa<Z�a</�a<��a<��a<!�a<ɟa<g�a<�a<��a<S�a<
�a<w�a<#�a<��a<B�a<ߛa<M�a<�a<W�a<�a<��a<�a<��a<�a<��a<:�a<�a<p�a<�a<��a<��a<��a<%�a<��a</�a<��a<H�a<ϑa<��a<�a<��a<��a<��a<@�a<Ԏa<��a<��a<��a<B�a<�a<��a<>�a<�a<t�a<A�a<͊a<��a<2�a<Չa<��a<C�a<'�a<шa<��a<k�a<!�a<�a<ԇa<ׇa<��a<��a<Y�a<?�a<I�a<�a<��a<�a<ۆa<Іa<نa<ֆa<��a<׆a<��a<�a<Ԇa<��a<�a<�a<=�a<�  �  j�a<��a<��a<��a<�a<�a<5�a<o�a<��a<Έa<�a<O�a<��a<ʉa<�a<b�a<��a<�a<i�a<��a<�a<y�a<ьa<N�a<��a<�a<��a<�a<_�a<̏a<A�a<��a<�a<��a<��a<��a<�a<p�a<�a<X�a<��a<p�a<�a<l�a<��a<Z�a<�a<\�a<͘a<N�a<řa<A�a<˚a<@�a<��a<$�a<��a<�a<��a<�a<z�a<�a<[�a<̟a<?�a<��a<�a<��a<ۡa<8�a<��a<��a<-�a<x�a<ףa<�a<m�a<��a<�a<2�a<W�a<��a<��a<0�a<Z�a<��a<��a<�a<�a<(�a<U�a<k�a<��a<��a<ԧa<�a<�a<�a</�a<J�a<k�a<��a<��a<��a<��a<��a<٨a<�a<�a<��a<��a<�a<��a<�a<Ԩa<�a<�a<Ѩa<רa<��a<��a<��a<x�a<��a<u�a<h�a<H�a<1�a<�a<�a<ѧa<��a<��a<Y�a<*�a<�a<�a<��a<��a<U�a<.�a<�a<٥a<��a<t�a<@�a<�a<ؤa<��a<{�a<<�a<�a<ãa<��a<E�a<�a<��a<^�a<�a<��a<�a< �a<Ӡa<t�a<�a<�a<z�a<�a<��a<`�a<�a<��a<�a<��a<5�a<��a<Q�a<�a<w�a<��a<��a<�a<��a<3�a<×a<A�a<ʖa<X�a<�a<y�a<�a<��a</�a<��a<;�a<˒a<_�a<Бa<Y�a<��a<��a<�a<��a<;�a<׎a<V�a<�a<��a<X�a<�a<��a<9�a<ڋa<��a<�a<ӊa<v�a<,�a<�a<��a<Y�a<�a<шa<��a<d�a<<�a<�a<ׇa<��a<��a<l�a<]�a<E�a<�a<�a<�a<��a<�a<�a<��a<Æa<Ɔa<a<چa<Іa<�a<�a<�a<4�a<D�a<�  �  n�a<n�a<��a<��a<�a<�a<G�a<��a<��a<�a<�a<L�a<��a<Ήa<'�a<^�a<Ɗa<��a<^�a<͋a<�a<��a<ڌa<T�a<��a<�a<��a<�a<\�a<��a<E�a<��a<$�a<p�a<�a<��a<Вa<w�a<�a<m�a<�a<Q�a<��a<X�a<��a<M�a<�a<Z�a<�a<c�a<Йa<]�a<��a<D�a<��a<2�a<��a<�a<��a<��a<��a<��a<n�a<��a<=�a<��a<��a<��a<ˡa<=�a<z�a<Ңa<A�a<x�a<ߣa< �a<n�a<��a<פa<F�a<`�a<åa<ǥa<"�a<Y�a<��a<��a<Цa<#�a<,�a<��a<q�a<��a<��a<��a<��a<��a<)�a<:�a<X�a<i�a<r�a<��a<��a<بa<Өa<بa<�a<ڨa<��a<�a<�a<Ϩa<��a<�a<�a<ߨa<��a<�a<��a<��a<��a<��a<��a<B�a<m�a<5�a<3�a<�a<�a<Χa<��a<��a<U�a<I�a<�a<ߦa<��a<��a<k�a<)�a<�a<ɥa<��a<��a<A�a<A�a<�a<��a<f�a<9�a<�a<��a<��a<�a<�a<��a<p�a<��a<��a<��a<�a<۠a<v�a<*�a<Ɵa<\�a<!�a<��a<d�a<՝a<��a<�a<Üa<J�a<̛a<m�a<Қa<z�a<��a<��a<�a<��a<;�a<��a<Z�a<ܖa<k�a<�a<w�a<�a<}�a<0�a<��a<@�a<��a<<�a<�a<Y�a<�a<g�a<�a<��a<%�a<�a<^�a< �a<��a<J�a<�a<��a<5�a<ċa<��a<"�a< �a<{�a<@�a<�a<��a<k�a<�a<�a<��a<r�a<:�a<��a<��a<��a<��a<��a<]�a<D�a<�a<�a<�a<�a<��a<چa<ʆa<ˆa<ņa<��a<�a<��a<܆a<��a<�a<.�a<�a<�  �  j�a<j�a<��a<؇a<��a<�a<I�a<i�a<��a<�a<�a<f�a<��a<Չa<!�a<l�a<��a<%�a<b�a<ˋa<�a<z�a<��a<H�a<��a<!�a<t�a<֎a<\�a<��a<(�a<��a<�a<�a<��a<Y�a<�a<g�a<ӓa<X�a<�a<c�a<�a<U�a<�a<o�a<�a<Y�a<�a<O�a<ݙa<P�a<˚a<E�a<��a<*�a<��a<*�a<��a<�a<��a<�a<`�a<�a<>�a<��a<�a<��a<ša<6�a<��a<�a<'�a<o�a<ʣa<�a<Q�a<��a<�a<,�a<_�a<��a<�a<&�a<O�a<}�a<Ǧa<�a<�a<0�a<[�a<v�a<��a<��a<�a<�a<�a<$�a<=�a<U�a<y�a<��a<��a<��a<��a<Ԩa<֨a<�a<��a<�a<�a<�a<�a<�a<�a<ըa<ۨa<Ԩa<��a<��a<��a<��a<��a<~�a<g�a<h�a<0�a<'�a< �a<��a<̧a<��a<|�a<\�a<B�a<�a<��a<��a<��a<e�a<8�a<�a<�a<��a<��a<K�a<�a<�a<��a<��a<M�a<��a<��a<��a<3�a<�a<��a<X�a<
�a<��a<W�a< �a<ʠa<e�a<�a<ɟa<m�a<�a<��a<W�a<��a<��a<�a<��a<6�a<ٛa<`�a<�a<|�a<�a<��a<�a<��a<5�a<ʗa<P�a<�a<]�a<��a<w�a<�a<��a<+�a<��a<9�a<��a<K�a<ˑa<O�a<�a<��a<�a<��a<9�a<юa<]�a<�a<��a<N�a<�a<��a<B�a<�a<��a<'�a<يa<��a<B�a<�a<��a<]�a<�a<݈a<��a<o�a<J�a<�a<�a<��a<��a<��a<[�a<K�a<;�a<�a<�a<��a<نa<цa<��a<��a<��a<Ɔa<��a<׆a<݆a<�a<��a<�a<6�a<�  �  C�a<��a<��a<��a<�a<�a<X�a<h�a<��a<ۈa<�a<]�a<��a<�a<�a<��a<��a<!�a<e�a<ʋa<3�a<w�a<��a<A�a<��a<
�a<�a<�a<:�a<ʏa<�a<��a<��a<q�a<��a<R�a<��a<D�a<�a<N�a<�a<b�a<ߕa<u�a<ݖa<`�a<�a<k�a<�a<R�a<�a<D�a<ߚa<;�a<ɛa<8�a<��a<;�a<��a<'�a<|�a<�a<h�a<�a<U�a<��a<�a<q�a<�a</�a<�a<�a<�a<��a<��a<�a<G�a<��a<�a<�a<q�a<��a<��a<�a<Z�a<��a<��a<�a<�a<M�a<Y�a<��a<��a<��a<�a<�a<,�a<�a<T�a<U�a<q�a<��a<��a<Ĩa<��a<ܨa<�a<ߨa<�a<�a<�a<�a<��a<�a<ۨa<�a<��a<ۨa<��a<Ĩa<��a<��a<��a<q�a<w�a<A�a<N�a<)�a<	�a<�a<֧a<��a<z�a<x�a<7�a<�a<�a<��a<��a<R�a<U�a<��a<�a<��a<��a<b�a<�a<��a<��a<w�a<5�a<�a<ţa<f�a<D�a<٢a<��a<J�a<��a<��a<P�a<(�a<��a<z�a<�a<˟a<l�a<�a<Þa<I�a<�a<��a<%�a<��a<:�a<�a<T�a<�a<q�a<�a<��a<�a<��a<&�a<חa<C�a<�a<d�a<��a<��a<
�a<��a<�a<��a<2�a<��a<Q�a<��a<e�a<ːa<��a<��a<��a<0�a<��a<p�a<��a<��a<5�a<�a<��a<.�a<֋a<~�a<C�a<׊a<��a<E�a<�a<��a<M�a<<�a<шa<��a<o�a<B�a<�a<�a<هa<��a<��a<h�a<>�a<'�a<�a<�a<چa<�a<Ɇa<��a<��a<��a<͆a<��a<܆a<Æa<�a<��a<�a<E�a<�  �  E�a<v�a<��a<͇a<�a<�a<;�a<��a<��a<�a<�a<\�a<��a<�a<�a<��a<ϊa<�a<k�a<ϋa<(�a<��a<׌a<K�a<��a<�a<q�a<�a<8�a<��a<#�a<��a<�a<n�a<�a<Y�a<ڒa<U�a<�a<U�a<��a<R�a<ߕa<W�a<�a<j�a<��a<X�a<�a<g�a<�a<W�a<ɚa<S�a<Λa<C�a<��a<9�a<��a<�a<��a<	�a<w�a<�a<;�a<��a<�a<|�a<ơa<0�a<t�a<ݢa<#�a<|�a<��a<
�a<E�a<��a<ڤa<!�a<]�a<��a<ߥa<
�a<X�a<|�a<æa<��a<�a<+�a<m�a<��a<��a<��a<֧a<�a<#�a<�a<V�a<e�a<{�a<��a<��a<��a<֨a<Ĩa<ڨa<��a<��a<�a<�a<�a<�a<�a<ըa<�a<¨a<��a<��a<��a<��a<��a<z�a<y�a<\�a<C�a<=�a<!�a<�a<�a<Чa<��a<��a<j�a<F�a<�a<�a<ɦa<��a<Y�a<N�a<�a<ߥa<��a<��a<X�a<0�a<ߤa<��a<��a<E�a<��a<��a<d�a<&�a<�a<��a<R�a<��a<��a<W�a<�a<��a<y�a<�a<şa<\�a<�a<��a<U�a<�a<��a<�a<��a<O�a<ߛa<g�a<�a<��a<�a<��a<$�a<��a<C�a<a<V�a<�a<t�a< �a<u�a<�a<��a<%�a<��a<3�a<��a<H�a<Ǒa<]�a<ڐa<p�a<�a<��a<)�a<Ǝa<\�a<��a<��a<2�a<�a<��a<=�a<�a<��a<"�a<�a<��a<E�a<��a<��a<q�a<3�a<؈a<��a<�a<L�a<�a<�a<ʇa<��a<s�a<_�a<U�a<2�a<�a<��a<܆a<φa<͆a<��a<ǆa<��a<��a<��a<��a<Ȇa<��a<�a<�a<+�a<�  �  s�a<t�a<��a<��a<�a<&�a<B�a<��a<��a<��a<!�a<s�a<��a<։a<P�a<d�a<׊a<'�a<y�a<֋a<
�a<��a<܌a<W�a<��a<�a<s�a<�a<[�a<��a<0�a<x�a<��a<p�a<�a<]�a<Ȓa<b�a<��a<Y�a<ܔa<P�a<�a<U�a<��a<K�a<�a<d�a<�a<a�a<ƙa<s�a<ʚa<l�a<��a<F�a<ɜa<!�a<��a<�a<��a<��a<i�a<�a<D�a<��a<��a<��a<ơa<J�a<}�a<Ӣa<+�a<W�a<ãa<��a<K�a<��a<֤a<�a<D�a<��a<ҥa<"�a<]�a<�a<æa<Ϧa<'�a<1�a<v�a<r�a<��a<Чa<�a<�a<�a<P�a<A�a<Z�a<��a<��a<��a<��a<֨a<Ψa<�a<�a<ڨa<��a<�a<�a<ڨa<�a<Ϩa<��a<Ҩa<��a<��a<��a<��a<��a<q�a<�a<S�a<q�a<:�a<%�a< �a<�a<ݧa<��a<��a<B�a<[�a<�a<�a<Ǧa<��a<��a<0�a<&�a<��a<��a<��a<:�a<=�a<�a<Ĥa<d�a<A�a<��a<��a<��a<�a<�a<��a<E�a<��a<��a<[�a<��a<Ša<O�a<�a<��a<Z�a</�a<��a<a�a<ӝa<��a<�a<��a<H�a<a<��a<�a<��a<�a<��a<9�a<��a<[�a<ȗa<p�a<֖a<f�a<�a<~�a<�a<|�a<1�a<��a<M�a<��a<>�a<Αa<8�a<�a<_�a<��a<��a<%�a<��a<C�a<�a<��a<J�a<�a<��a<=�a<Ëa<��a<'�a<�a<|�a<F�a<�a<��a<�a<�a<	�a<��a<s�a<d�a<�a<�a<��a<��a<~�a<k�a<>�a<�a<�a<�a<�a<Ća<цa<��a<��a<��a<��a<��a<��a<ӆa<ֆa<�a<�a<!�a<�  �  I�a<c�a<��a<Ǉa<�a<%�a<R�a<��a<��a<�a<�a<h�a<��a<�a<D�a<�a<Պa<!�a<b�a<�a<4�a<��a<�a<U�a<��a<�a<s�a<̎a<>�a<��a<�a<��a<��a<d�a<Ցa<O�a<͒a<O�a<ғa<O�a<Ȕa<G�a<ԕa<S�a<�a<d�a<�a<p�a<�a<t�a<��a<h�a<Śa<Y�a<ϛa<M�a<ʜa<;�a<��a<�a<��a<�a<��a<�a<Q�a<��a<�a<~�a<ȡa<�a<m�a<��a<�a<o�a<��a<��a<=�a<��a<Ϥa<�a<a�a<��a<ͥa<�a<=�a<��a<��a<ڦa<!�a<D�a<r�a<��a<§a<��a<�a<�a<"�a<J�a<Q�a<m�a<��a<x�a<��a<Ũa<֨a<٨a<�a<�a<�a<��a<ߨa<�a<ڨa<רa<ިa<ͨa<��a<��a<��a<��a<��a<��a<��a<c�a<W�a<H�a<*�a<'�a<�a<�a<ܧa<��a<��a<w�a<]�a<�a<��a<Ԧa<��a<��a<K�a<$�a<�a<��a<��a<d�a<8�a<��a<¤a<n�a<=�a<��a<��a<j�a<�a<Ѣa<��a<G�a<�a<��a<M�a<��a<��a<d�a<�a<��a<R�a<�a<��a<Y�a<�a<��a<*�a<��a<[�a<�a<x�a<�a<��a<�a<��a<:�a<��a<P�a<ȗa<^�a<��a<��a<�a<��a<�a<��a<(�a<��a< �a<��a<*�a<��a<O�a<ِa<^�a<�a<��a<�a<��a<_�a<�a<��a<4�a<ьa<��a<5�a<ϋa<��a<:�a<��a<��a<^�a<�a<��a<y�a<3�a<�a<��a<��a<T�a<�a<�a<ڇa<��a<��a<j�a<@�a<+�a<�a<�a<݆a<Ća<��a<��a<��a<��a<��a<��a<��a<ņa<݆a<��a<�a<%�a<�  �  E�a<��a<��a<Ǉa<�a<�a<G�a<u�a<��a<�a<>�a<m�a<��a<��a<�a<��a<��a<7�a<��a<ϋa<'�a<~�a<�a<E�a<͍a<	�a<s�a<�a<@�a<Əa<	�a<��a<ݐa<k�a<ݑa<R�a<�a<8�a<ϓa<=�a<Ҕa<j�a<Еa<r�a<Ӗa<u�a<�a<e�a<�a<_�a<�a<T�a<��a<T�a<כa<B�a<��a<D�a<��a<D�a<��a<�a<q�a<ޟa<I�a<��a<*�a<b�a<�a<�a<��a<Ԣa<�a<l�a<��a<
�a<E�a<��a<פa<��a<X�a<��a<�a<�a<S�a<��a<��a<�a<�a<8�a<]�a<��a<��a<Χa<�a<��a<3�a<$�a<^�a<g�a<��a<��a<��a<��a<��a<Шa<רa<��a<�a<ߨa<�a<�a<��a<Ѩa<Ȩa<èa<��a<èa<��a<��a<��a<z�a<s�a<^�a<x�a<C�a<P�a<�a<�a<�a<ɧa<��a<��a<q�a<B�a<8�a< �a<Ŧa<��a<_�a<_�a<�a<�a<̥a<��a<V�a<�a<�a<��a<��a<5�a<��a<ãa<k�a<?�a<̢a<��a<)�a<��a<��a<P�a<�a<��a<a�a<��a<��a<t�a<��a<��a<?�a<��a<��a< �a<��a<F�a<ޛa<d�a<�a<��a< �a<��a<!�a<Șa<B�a<��a<V�a<�a<m�a<��a<��a<�a<��a<�a<��a<#�a<��a<>�a<��a<M�a<��a<p�a<�a<��a<%�a<��a<W�a<�a<��a<=�a<�a<��a<%�a<��a<��a</�a<ۊa<��a<G�a< �a<Љa<e�a<C�a<݈a<ňa<��a<U�a<:�a<�a<чa<��a<�a<\�a<W�a<.�a< �a<�a<؆a<�a<��a<��a<��a<��a<��a<��a<��a<Æa<͆a<�a<��a<F�a<�  �  ?�a<}�a<��a<��a<�a<�a<`�a<��a<��a<�a<4�a<e�a<��a<	�a<N�a<��a<��a<0�a<��a<ڋa<2�a<��a<��a<H�a<��a<�a<q�a<ݎa<7�a<��a<�a<��a<�a<i�a<ʑa<E�a<��a<L�a<ēa<S�a<��a<K�a<͕a<k�a<ږa<]�a<�a<s�a<�a<x�a<�a<c�a<�a<O�a<̛a<[�a<՜a<>�a<��a<5�a<��a<�a<��a<��a<Y�a<��a<�a<i�a<ڡa<�a<o�a<��a<"�a<a�a<��a<�a<7�a<{�a<ˤa<�a<W�a<��a<ƥa<�a<G�a<��a<��a<�a<�a<Q�a<|�a<��a<��a<ԧa<��a<��a<5�a<U�a<l�a<\�a<�a<��a<��a<��a<ըa<�a<�a<�a<ިa<�a<��a<ݨa<ݨa<Шa<֨a<Ũa<èa<��a<��a<��a<��a<��a<}�a<a�a<R�a<=�a<C�a<�a<��a<��a<էa<ǧa<��a<t�a<M�a<.�a<��a<��a<��a<��a<d�a<�a<��a<ɥa<��a<b�a<:�a<�a<��a<{�a<1�a<��a<��a<c�a<�a<ۢa<��a<>�a<��a<��a<C�a<�a<��a<V�a<�a<��a<V�a<��a<��a<E�a<�a<��a<-�a<Ӝa<_�a<�a<s�a<�a<��a<�a<��a<E�a<Øa<:�a<�a<d�a<��a<��a<�a<��a<�a<��a<�a<��a<�a<��a<#�a<Ƒa<B�a<Ԑa<R�a<�a<x�a<�a<��a<U�a<��a<��a<+�a<یa<��a<&�a<׋a<��a<G�a<��a<��a<T�a<�a<ǉa<a�a<E�a<�a<ӈa<v�a<P�a<1�a<��a<Շa<��a<��a<h�a<J�a<�a<�a<�a<Ԇa<Ɔa<��a<��a<��a<��a<��a<��a<��a<Ɇa<Ԇa<�a<�a<!�a<�  �  X�a<]�a<��a<҇a<�a<�a<?�a<s�a<��a<��a<�a<��a<��a<�a<*�a<v�a<�a<9�a<g�a<�a<%�a<x�a<�a<S�a<��a<)�a<s�a<ʎa<]�a<��a<�a<s�a<��a<[�a<בa<p�a<��a<_�a<��a<a�a<Δa<e�a<�a<M�a<�a<j�a<�a<Y�a<Ϙa<X�a<�a<d�a<њa<t�a<ٛa<D�a<��a<A�a<ɝa<&�a<��a<�a<j�a<ʟa<=�a<��a<�a<��a<ša<,�a<��a<ʢa</�a<F�a<ţa<�a<U�a<��a<��a<�a<=�a<��a<ҥa</�a<B�a<�a<Ԧa<�a<�a<9�a<P�a<�a<��a<��a<��a<�a<�a<6�a<F�a<{�a<��a<��a<��a<��a<��a<Ũa<ըa<�a<��a<��a<Өa<��a<�a<ۨa<بa<��a<Ȩa<��a<Шa<��a<��a<x�a<x�a<j�a<]�a<W�a<#�a<0�a<�a<��a<ҧa<��a<��a<m�a<[�a<�a<�a<�a<��a<n�a<B�a<2�a<�a<��a<��a<U�a<�a<�a<��a<x�a<T�a<��a<��a<��a<�a<ܢa<|�a<A�a<�a<��a<n�a<�a<àa<@�a<�a<��a<o�a<�a<��a<[�a<�a<��a<�a<��a<@�a<�a<t�a<��a<��a<"�a<��a<0�a<Řa<c�a<֗a<^�a<�a<g�a<�a<w�a<�a<��a<0�a<��a</�a<Ȓa<4�a<ӑa<'�a<�a<H�a<�a<��a<	�a<��a<<�a<��a<��a<X�a<֌a<��a<N�a<׋a<��a</�a<Ίa<��a<Z�a<�a<Éa<��a<+�a<�a<��a<��a<r�a<�a<�a<Ӈa<��a<u�a<Y�a<K�a<5�a<�a<܆a<�a<ӆa<��a<��a<��a<��a<��a<҆a<��a<Ɔa<ˆa<�a<
�a<+�a<�  �  ?�a<}�a<��a<��a<�a<�a<`�a<��a<��a<�a<4�a<e�a<��a<	�a<N�a<��a<��a<0�a<��a<ڋa<2�a<��a<��a<H�a<��a<�a<q�a<ݎa<7�a<��a<�a<��a<�a<i�a<ʑa<E�a<��a<L�a<ēa<S�a<��a<K�a<͕a<k�a<ږa<]�a<�a<s�a<�a<x�a<�a<c�a<�a<O�a<̛a<[�a<՜a<>�a<��a<5�a<��a<�a<��a<��a<Y�a<��a<�a<i�a<ڡa<�a<o�a<��a<"�a<a�a<��a<�a<7�a<{�a<ˤa<�a<W�a<��a<ƥa<�a<G�a<��a<��a<�a<�a<Q�a<|�a<��a<��a<ԧa<��a<��a<5�a<U�a<l�a<\�a<�a<��a<��a<��a<ըa<�a<�a<�a<ިa<�a<��a<ݨa<ݨa<Шa<֨a<Ũa<èa<��a<��a<��a<��a<��a<}�a<a�a<R�a<=�a<C�a<�a<��a<��a<էa<ǧa<��a<t�a<M�a<.�a<��a<��a<��a<��a<d�a<�a<��a<ɥa<��a<b�a<:�a<�a<��a<{�a<1�a<��a<��a<c�a<�a<ۢa<��a<>�a<��a<��a<C�a<�a<��a<V�a<�a<��a<V�a<��a<��a<E�a<�a<��a<-�a<Ӝa<_�a<�a<s�a<�a<��a<�a<��a<E�a<Øa<:�a<�a<d�a<��a<��a<�a<��a<�a<��a<�a<��a<�a<��a<#�a<Ƒa<B�a<Ԑa<R�a<�a<x�a<�a<��a<U�a<��a<��a<+�a<یa<��a<&�a<׋a<��a<G�a<��a<��a<T�a<�a<ǉa<a�a<E�a<�a<ӈa<v�a<P�a<1�a<��a<Շa<��a<��a<h�a<J�a<�a<�a<�a<Ԇa<Ɔa<��a<��a<��a<��a<��a<��a<��a<Ɇa<Ԇa<�a<�a<!�a<�  �  E�a<��a<��a<Ǉa<�a<�a<G�a<u�a<��a<�a<>�a<m�a<��a<��a<�a<��a<��a<7�a<��a<ϋa<'�a<~�a<�a<E�a<͍a<	�a<s�a<�a<@�a<Əa<	�a<��a<ݐa<k�a<ݑa<R�a<�a<8�a<ϓa<=�a<Ҕa<j�a<Еa<r�a<Ӗa<u�a<�a<e�a<�a<_�a<�a<T�a<��a<T�a<כa<B�a<��a<D�a<��a<D�a<��a<�a<q�a<ޟa<I�a<��a<*�a<b�a<�a<�a<��a<Ԣa<�a<l�a<��a<
�a<E�a<��a<פa<��a<X�a<��a<�a<�a<S�a<��a<��a<�a<�a<8�a<]�a<��a<��a<Χa<�a<��a<3�a<$�a<^�a<g�a<��a<��a<��a<��a<��a<Шa<רa<��a<�a<ߨa<�a<�a<��a<Ѩa<Ȩa<èa<��a<èa<��a<��a<��a<z�a<s�a<^�a<x�a<C�a<P�a<�a<�a<�a<ɧa<��a<��a<q�a<B�a<8�a< �a<Ŧa<��a<_�a<_�a<�a<�a<̥a<��a<V�a<�a<�a<��a<��a<5�a<��a<ãa<k�a<?�a<̢a<��a<)�a<��a<��a<P�a<�a<��a<a�a<��a<��a<t�a<��a<��a<?�a<��a<��a< �a<��a<F�a<ޛa<d�a<�a<��a< �a<��a<!�a<Șa<B�a<��a<V�a<�a<m�a<��a<��a<�a<��a<�a<��a<#�a<��a<>�a<��a<M�a<��a<p�a<�a<��a<%�a<��a<W�a<�a<��a<=�a<�a<��a<%�a<��a<��a</�a<ۊa<��a<G�a< �a<Љa<e�a<C�a<݈a<ňa<��a<U�a<:�a<�a<чa<��a<�a<\�a<W�a<.�a< �a<�a<؆a<�a<��a<��a<��a<��a<��a<��a<��a<Æa<͆a<�a<��a<F�a<�  �  I�a<c�a<��a<Ǉa<�a<%�a<R�a<��a<��a<�a<�a<h�a<��a<�a<D�a<�a<Պa<!�a<b�a<�a<4�a<��a<�a<U�a<��a<�a<s�a<̎a<>�a<��a<�a<��a<��a<d�a<Ցa<O�a<͒a<O�a<ғa<O�a<Ȕa<G�a<ԕa<S�a<�a<d�a<�a<p�a<�a<t�a<��a<h�a<Śa<Y�a<ϛa<M�a<ʜa<;�a<��a<�a<��a<�a<��a<�a<Q�a<��a<�a<~�a<ȡa<�a<m�a<��a<�a<o�a<��a<��a<=�a<��a<Ϥa<�a<a�a<��a<ͥa<�a<=�a<��a<��a<ڦa<!�a<D�a<r�a<��a<§a<��a<�a<�a<"�a<J�a<Q�a<m�a<��a<x�a<��a<Ũa<֨a<٨a<�a<�a<�a<��a<ߨa<�a<ڨa<רa<ިa<ͨa<��a<��a<��a<��a<��a<��a<��a<c�a<W�a<H�a<*�a<'�a<�a<�a<ܧa<��a<��a<w�a<]�a<�a<��a<Ԧa<��a<��a<K�a<$�a<�a<��a<��a<d�a<8�a<��a<¤a<n�a<=�a<��a<��a<j�a<�a<Ѣa<��a<G�a<�a<��a<M�a<��a<��a<d�a<�a<��a<R�a<�a<��a<Y�a<�a<��a<*�a<��a<[�a<�a<x�a<�a<��a<�a<��a<:�a<��a<P�a<ȗa<^�a<��a<��a<�a<��a<�a<��a<(�a<��a< �a<��a<*�a<��a<O�a<ِa<^�a<�a<��a<�a<��a<_�a<�a<��a<4�a<ьa<��a<5�a<ϋa<��a<:�a<��a<��a<^�a<�a<��a<y�a<3�a<�a<��a<��a<T�a<�a<�a<ڇa<��a<��a<j�a<@�a<+�a<�a<�a<݆a<Ća<��a<��a<��a<��a<��a<��a<��a<ņa<݆a<��a<�a<%�a<�  �  s�a<t�a<��a<��a<�a<&�a<B�a<��a<��a<��a<!�a<s�a<��a<։a<P�a<d�a<׊a<'�a<y�a<֋a<
�a<��a<܌a<W�a<��a<�a<s�a<�a<[�a<��a<0�a<x�a<��a<p�a<�a<]�a<Ȓa<b�a<��a<Y�a<ܔa<P�a<�a<U�a<��a<K�a<�a<d�a<�a<a�a<ƙa<s�a<ʚa<l�a<��a<F�a<ɜa<!�a<��a<�a<��a<��a<i�a<�a<D�a<��a<��a<��a<ơa<J�a<}�a<Ӣa<+�a<W�a<ãa<��a<K�a<��a<֤a<�a<D�a<��a<ҥa<"�a<]�a<�a<æa<Ϧa<'�a<1�a<v�a<r�a<��a<Чa<�a<�a<�a<P�a<A�a<Z�a<��a<��a<��a<��a<֨a<Ψa<�a<�a<ڨa<��a<�a<�a<ڨa<�a<Ϩa<��a<Ҩa<��a<��a<��a<��a<��a<q�a<�a<S�a<q�a<:�a<%�a< �a<�a<ݧa<��a<��a<B�a<[�a<�a<�a<Ǧa<��a<��a<0�a<&�a<��a<��a<��a<:�a<=�a<�a<Ĥa<d�a<A�a<��a<��a<��a<�a<�a<��a<E�a<��a<��a<[�a<��a<Ša<O�a<�a<��a<Z�a</�a<��a<a�a<ӝa<��a<�a<��a<H�a<a<��a<�a<��a<�a<��a<9�a<��a<[�a<ȗa<p�a<֖a<f�a<�a<~�a<�a<|�a<1�a<��a<M�a<��a<>�a<Αa<8�a<�a<_�a<��a<��a<%�a<��a<C�a<�a<��a<J�a<�a<��a<=�a<Ëa<��a<'�a<�a<|�a<F�a<�a<��a<�a<�a<	�a<��a<s�a<d�a<�a<�a<��a<��a<~�a<k�a<>�a<�a<�a<�a<�a<Ća<цa<��a<��a<��a<��a<��a<��a<ӆa<ֆa<�a<�a<!�a<�  �  E�a<v�a<��a<͇a<�a<�a<;�a<��a<��a<�a<�a<\�a<��a<�a<�a<��a<ϊa<�a<k�a<ϋa<(�a<��a<׌a<K�a<��a<�a<q�a<�a<8�a<��a<#�a<��a<�a<n�a<�a<Y�a<ڒa<U�a<�a<U�a<��a<R�a<ߕa<W�a<�a<j�a<��a<X�a<�a<g�a<�a<W�a<ɚa<S�a<Λa<C�a<��a<9�a<��a<�a<��a<	�a<w�a<�a<;�a<��a<�a<|�a<ơa<0�a<t�a<ݢa<#�a<|�a<��a<
�a<E�a<��a<ڤa<!�a<]�a<��a<ߥa<
�a<X�a<|�a<æa<��a<�a<+�a<m�a<��a<��a<��a<֧a<�a<#�a<�a<V�a<e�a<{�a<��a<��a<��a<֨a<Ĩa<ڨa<��a<��a<�a<�a<�a<�a<�a<ըa<�a<¨a<��a<��a<��a<��a<��a<z�a<y�a<\�a<C�a<=�a<!�a<�a<�a<Чa<��a<��a<j�a<F�a<�a<�a<ɦa<��a<Y�a<N�a<�a<ߥa<��a<��a<X�a<0�a<ߤa<��a<��a<E�a<��a<��a<d�a<&�a<�a<��a<R�a<��a<��a<W�a<�a<��a<y�a<�a<şa<\�a<�a<��a<U�a<�a<��a<�a<��a<O�a<ߛa<g�a<�a<��a<�a<��a<$�a<��a<C�a<a<V�a<�a<t�a< �a<u�a<�a<��a<%�a<��a<3�a<��a<H�a<Ǒa<]�a<ڐa<p�a<�a<��a<)�a<Ǝa<\�a<��a<��a<2�a<�a<��a<=�a<�a<��a<"�a<�a<��a<E�a<��a<��a<q�a<3�a<؈a<��a<�a<L�a<�a<�a<ʇa<��a<s�a<_�a<U�a<2�a<�a<��a<܆a<φa<͆a<��a<ǆa<��a<��a<��a<��a<Ȇa<��a<�a<�a<+�a<�  �  C�a<��a<��a<��a<�a<�a<X�a<h�a<��a<ۈa<�a<]�a<��a<�a<�a<��a<��a<!�a<e�a<ʋa<3�a<w�a<��a<A�a<��a<
�a<�a<�a<:�a<ʏa<�a<��a<��a<q�a<��a<R�a<��a<D�a<�a<N�a<�a<b�a<ߕa<u�a<ݖa<`�a<�a<k�a<�a<R�a<�a<D�a<ߚa<;�a<ɛa<8�a<��a<;�a<��a<'�a<|�a<�a<h�a<�a<U�a<��a<�a<q�a<�a</�a<�a<�a<�a<��a<��a<�a<G�a<��a<�a<�a<q�a<��a<��a<�a<Z�a<��a<��a<�a<�a<M�a<Y�a<��a<��a<��a<�a<�a<,�a<�a<T�a<U�a<q�a<��a<��a<Ĩa<��a<ܨa<�a<ߨa<�a<�a<�a<�a<��a<�a<ۨa<�a<��a<ۨa<��a<Ĩa<��a<��a<��a<q�a<w�a<A�a<N�a<)�a<	�a<�a<֧a<��a<z�a<x�a<7�a<�a<�a<��a<��a<R�a<U�a<��a<�a<��a<��a<b�a<�a<��a<��a<w�a<5�a<�a<ţa<f�a<D�a<٢a<��a<J�a<��a<��a<P�a<(�a<��a<z�a<�a<˟a<l�a<�a<Þa<I�a<�a<��a<%�a<��a<:�a<�a<T�a<�a<q�a<�a<��a<�a<��a<&�a<חa<C�a<�a<d�a<��a<��a<
�a<��a<�a<��a<2�a<��a<Q�a<��a<e�a<ːa<��a<��a<��a<0�a<��a<p�a<��a<��a<5�a<�a<��a<.�a<֋a<~�a<C�a<׊a<��a<E�a<�a<��a<M�a<<�a<шa<��a<o�a<B�a<�a<�a<هa<��a<��a<h�a<>�a<'�a<�a<�a<چa<�a<Ɇa<��a<��a<��a<͆a<��a<܆a<Æa<�a<��a<�a<E�a<�  �  j�a<j�a<��a<؇a<��a<�a<I�a<i�a<��a<�a<�a<f�a<��a<Չa<!�a<l�a<��a<%�a<b�a<ˋa<�a<z�a<��a<H�a<��a<!�a<t�a<֎a<\�a<��a<(�a<��a<�a<�a<��a<Y�a<�a<g�a<ӓa<X�a<�a<c�a<�a<U�a<�a<o�a<�a<Y�a<�a<O�a<ݙa<P�a<˚a<E�a<��a<*�a<��a<*�a<��a<�a<��a<�a<`�a<�a<>�a<��a<�a<��a<ša<6�a<��a<�a<'�a<o�a<ʣa<�a<Q�a<��a<�a<,�a<_�a<��a<�a<&�a<O�a<}�a<Ǧa<�a<�a<0�a<[�a<v�a<��a<��a<�a<�a<�a<$�a<=�a<U�a<y�a<��a<��a<��a<��a<Ԩa<֨a<�a<��a<�a<�a<�a<�a<�a<�a<ըa<ۨa<Ԩa<��a<��a<��a<��a<��a<~�a<g�a<h�a<0�a<'�a< �a<��a<̧a<��a<|�a<\�a<B�a<�a<��a<��a<��a<e�a<8�a<�a<�a<��a<��a<K�a<�a<�a<��a<��a<M�a<��a<��a<��a<3�a<�a<��a<X�a<
�a<��a<W�a< �a<ʠa<e�a<�a<ɟa<m�a<�a<��a<W�a<��a<��a<�a<��a<6�a<ٛa<`�a<�a<|�a<�a<��a<�a<��a<5�a<ʗa<P�a<�a<]�a<��a<w�a<�a<��a<+�a<��a<9�a<��a<K�a<ˑa<O�a<�a<��a<�a<��a<9�a<юa<]�a<�a<��a<N�a<�a<��a<B�a<�a<��a<'�a<يa<��a<B�a<�a<��a<]�a<�a<݈a<��a<o�a<J�a<�a<�a<��a<��a<��a<[�a<K�a<;�a<�a<�a<��a<نa<цa<��a<��a<��a<Ɔa<��a<׆a<݆a<�a<��a<�a<6�a<�  �  n�a<n�a<��a<��a<�a<�a<G�a<��a<��a<�a<�a<L�a<��a<Ήa<'�a<^�a<Ɗa<��a<^�a<͋a<�a<��a<ڌa<T�a<��a<�a<��a<�a<\�a<��a<E�a<��a<$�a<p�a<�a<��a<Вa<w�a<�a<m�a<�a<Q�a<��a<X�a<��a<M�a<�a<Z�a<�a<c�a<Йa<]�a<��a<D�a<��a<2�a<��a<�a<��a<��a<��a<��a<n�a<��a<=�a<��a<��a<��a<ˡa<=�a<z�a<Ңa<A�a<x�a<ߣa< �a<n�a<��a<פa<F�a<`�a<åa<ǥa<"�a<Y�a<��a<��a<Цa<#�a<,�a<��a<q�a<��a<��a<��a<��a<��a<)�a<:�a<X�a<i�a<r�a<��a<��a<بa<Өa<بa<�a<ڨa<��a<�a<�a<Ϩa<��a<�a<�a<ߨa<��a<�a<��a<��a<��a<��a<��a<B�a<m�a<5�a<3�a<�a<�a<Χa<��a<��a<U�a<I�a<�a<ߦa<��a<��a<k�a<)�a<�a<ɥa<��a<��a<A�a<A�a<�a<��a<f�a<9�a<�a<��a<��a<�a<�a<��a<p�a<��a<��a<��a<�a<۠a<v�a<*�a<Ɵa<\�a<!�a<��a<d�a<՝a<��a<�a<Üa<J�a<̛a<m�a<Қa<z�a<��a<��a<�a<��a<;�a<��a<Z�a<ܖa<k�a<�a<w�a<�a<}�a<0�a<��a<@�a<��a<<�a<�a<Y�a<�a<g�a<�a<��a<%�a<�a<^�a< �a<��a<J�a<�a<��a<5�a<ċa<��a<"�a< �a<{�a<@�a<�a<��a<k�a<�a<�a<��a<r�a<:�a<��a<��a<��a<��a<��a<]�a<D�a<�a<�a<�a<�a<��a<چa<ʆa<ˆa<ņa<��a<�a<��a<܆a<��a<�a<.�a<�a<�  �  j�a<��a<��a<��a<�a<�a<5�a<o�a<��a<Έa<�a<O�a<��a<ʉa<�a<b�a<��a<�a<i�a<��a<�a<y�a<ьa<N�a<��a<�a<��a<�a<_�a<̏a<A�a<��a<�a<��a<��a<��a<�a<p�a<�a<X�a<��a<p�a<�a<l�a<��a<Z�a<�a<\�a<͘a<N�a<řa<A�a<˚a<@�a<��a<$�a<��a<�a<��a<�a<z�a<�a<[�a<̟a<?�a<��a<�a<��a<ۡa<8�a<��a<��a<-�a<x�a<ףa<�a<m�a<��a<�a<2�a<W�a<��a<��a<0�a<Z�a<��a<��a<�a<�a<(�a<U�a<k�a<��a<��a<ԧa<�a<�a<�a</�a<J�a<k�a<��a<��a<��a<��a<��a<٨a<�a<�a<��a<��a<�a<��a<�a<Ԩa<�a<�a<Ѩa<רa<��a<��a<��a<x�a<��a<u�a<h�a<H�a<1�a<�a<�a<ѧa<��a<��a<Y�a<*�a<�a<�a<��a<��a<U�a<.�a<�a<٥a<��a<t�a<@�a<�a<ؤa<��a<{�a<<�a<�a<ãa<��a<E�a<�a<��a<^�a<�a<��a<�a< �a<Ӡa<t�a<�a<�a<z�a<�a<��a<`�a<�a<��a<�a<��a<5�a<��a<Q�a<�a<w�a<��a<��a<�a<��a<3�a<×a<A�a<ʖa<X�a<�a<y�a<�a<��a</�a<��a<;�a<˒a<_�a<Бa<Y�a<��a<��a<�a<��a<;�a<׎a<V�a<�a<��a<X�a<�a<��a<9�a<ڋa<��a<�a<ӊa<v�a<,�a<�a<��a<Y�a<�a<шa<��a<d�a<<�a<�a<ׇa<��a<��a<l�a<]�a<E�a<�a<�a<�a<��a<�a<�a<��a<Æa<Ɔa<a<چa<Іa<�a<�a<�a<4�a<D�a<�  �  P�a<v�a<��a<߇a<�a<�a<Y�a<j�a<��a<Ɉa<�a<=�a<��a<։a<�a<s�a<��a<�a<S�a<��a<4�a<t�a<��a<8�a<��a<#�a<v�a<��a<E�a<��a< �a<��a<�a<��a<�a<\�a<��a<]�a<�a<d�a<�a<]�a<ߕa<a�a<�a<��a<՗a<i�a<ߘa<[�a<�a<=�a<Śa<!�a<��a<+�a<��a<'�a<z�a<�a<r�a< �a<s�a<ԟa<T�a<��a<-�a<{�a<ҡa<,�a<��a<ޢa<+�a<��a<ƣa<'�a<O�a<��a<�a<0�a<��a<��a<�a<�a<S�a<��a<Ħa<�a<�a<K�a<O�a<��a<��a<��a<Чa<קa<�a<�a<8�a<Q�a<P�a<z�a<��a<èa<��a<ݨa<Ԩa<�a<�a<�a<�a<�a<�a<�a<��a<��a<̨a<�a<��a<˨a<��a<��a<��a<z�a<o�a<N�a<<�a<�a<'�a<�a<ħa<��a<}�a<y�a<%�a<�a<Цa<��a<��a<R�a<>�a<��a<ҥa<��a<r�a<d�a<�a< �a<��a<��a<N�a<��a<��a<p�a<:�a<�a<��a<^�a<�a<ǡa<Z�a</�a<��a<��a<!�a<ɟa<g�a<�a<��a<S�a<
�a<w�a<#�a<��a<B�a<ߛa<M�a<�a<W�a<�a<��a<�a<��a<�a<��a<:�a<�a<p�a<�a<��a<��a<��a<%�a<��a</�a<��a<H�a<ϑa<��a<�a<��a<��a<��a<@�a<Ԏa<��a<��a<��a<B�a<�a<��a<>�a<�a<t�a<A�a<͊a<��a<2�a<Չa<��a<C�a<'�a<шa<��a<k�a<!�a<�a<ԇa<ׇa<��a<��a<Y�a<?�a<I�a<�a<��a<�a<ۆa<Іa<نa<ֆa<��a<׆a<��a<�a<Ԇa<��a<�a<�a<=�a<�  �  j�a<��a<��a<ʇa<݇a<�a<M�a<f�a<��a<шa<�a<H�a<��a<��a<�a<K�a<��a<�a<b�a<��a<�a<p�a<�a<>�a<��a<�a<��a<��a<_�a<Ǐa<,�a<��a<�a<w�a<�a<��a<��a<W�a<��a<m�a<�a<r�a< �a<w�a<�a<_�a<חa<a�a<Әa<F�a<��a<M�a<��a<9�a<��a<�a<��a<�a<��a<�a<��a<�a<Z�a<Οa<M�a<��a<�a<w�a<�a<N�a<��a<�a<9�a<��a<��a<$�a<w�a<��a<�a<+�a<��a<��a<�a<3�a<r�a<��a<��a<ܦa<�a<B�a<L�a<p�a<��a<��a<ǧa<�a<�a<�a<"�a<Q�a<c�a<~�a<��a<��a<��a<Ϩa<Өa<بa<�a<�a<�a<	�a<��a<��a<��a<�a<ɨa<�a<�a<٨a<��a<��a<��a<��a<r�a<i�a<S�a<*�a<�a<ߧa<ŧa<��a<x�a<T�a<-�a<�a<ۦa<��a<q�a<K�a<�a<�a<ϥa<��a<m�a<D�a<�a<�a<��a<l�a<C�a<�a<أa<��a<A�a<�a<��a<Y�a<�a<֡a<��a<0�a<��a<��a<*�a<ןa<}�a<-�a<Şa<R�a<�a<y�a<�a<��a<.�a<��a<]�a<�a<p�a<��a<y�a<�a<��a<,�a<��a<O�a<Öa<W�a<�a<��a< �a<��a< �a<��a<Q�a<Вa<V�a<ܑa<t�a<��a<��a<'�a<��a<4�a<Ўa<~�a<�a<��a<[�a<�a<��a<7�a<Ћa<{�a<8�a<ʊa<{�a<$�a<�a<��a<T�a< �a<ňa<��a<k�a<4�a<�a<߇a<��a<��a<�a<W�a<7�a<+�a<�a<�a<��a<�a<چa<҆a<φa<��a<߆a<�a<�a<Іa<��a<�a<%�a<A�a<�  �  N�a<Z�a<��a<��a<�a<�a<�a<p�a<z�a<��a<܇a<�a<e�a<��a<�a<,�a<��a<��a<7�a<��a<�a<��a<��a<J�a<��a<��a<n�a<ԍa<T�a<��a</�a<��a<&�a<��a<��a<��a<�a<��a<��a<Z�a<�a<j�a<��a<q�a<��a<s�a<�a<h�a<��a<��a<Әa<d�a<��a<=�a<��a<-�a<��a<%�a<��a<
�a<��a<�a<��a<�a<f�a<��a<F�a<��a<�a<g�a<��a<�a<Z�a<��a<%�a<E�a<��a<�a<$�a<��a<��a<�a<�a<b�a<��a<��a<�a<�a<\�a<S�a<��a<��a<��a<Ӧa<Ϧa<
�a<�a<8�a<;�a<e�a<i�a<��a<��a<��a<��a<��a<�a<&�a<�a<�a<�a<3�a<�a<3�a<�a<+�a<�a<��a<�a<�a<�a<�a<��a<��a<��a<��a<h�a<R�a<*�a<*�a<�a<Ʀa<ɦa<x�a<R�a<�a<إa<ϥa<��a<u�a<8�a<�a<̤a<��a<��a<u�a<_�a<��a<�a<��a<a�a<,�a<�a<��a<b�a<&�a<ˡa<��a<C�a<��a<��a<A�a<�a<��a<<�a<��a<��a<D�a<۝a<{�a<�a<Ɯa<5�a<ڛa<t�a<ؚa<z�a<�a<s�a<��a<��a<�a<��a<4�a<��a<X�a<ѕa<��a<�a<�a<3�a<��a<*�a<��a<=�a<Ƒa<P�a<ʐa<g�a<�a<s�a<�a<��a<7�a<�a<a�a<�a<��a<J�a<֋a<��a<�a<̊a<��a<�a<ԉa<t�a<�a<��a<T�a</�a<ڇa<��a<Z�a<6�a<�a<цa<��a<��a<��a<Y�a<G�a<:�a<�a<�a<݅a<߅a<��a<Ʌa<��a<��a<��a<��a<ƅa<��a<̅a<�a<ޅa<�a<�a<�  �  O�a<m�a<��a<��a<Ɇa<�a<�a<<�a<r�a<��a<�a<"�a<i�a<��a<�a<3�a<��a<�a<A�a<��a<�a<O�a<Ƌa<'�a<��a<�a<��a<�a<R�a<��a<5�a<��a<�a<|�a<��a<n�a<�a<f�a<�a<y�a<��a<z�a<�a<~�a< �a<|�a<�a<l�a<�a<Q�a<֘a<Q�a<Ιa<P�a<͚a<;�a<��a<4�a<��a<"�a<��a<�a<y�a<�a<m�a<џa<K�a<��a<�a<y�a<ˡa<(�a<w�a<��a<��a<Q�a<��a<�a< �a<^�a<��a<�a<)�a<`�a<��a<ҥa<��a<�a<3�a<b�a<o�a<��a<��a<צa<��a<�a<�a<8�a<K�a<u�a<��a<��a<��a<��a<˧a<�a<��a<�a<!�a<,�a</�a<9�a<&�a<-�a<�a<�a<��a<�a<�a<�a<Χa<ϧa<��a<��a<��a<��a<{�a<a�a<?�a<�a<�a<Ʀa<��a<q�a<I�a<'�a<��a<ԥa<��a<p�a<@�a<"�a<��a<Ȥa<��a<\�a<)�a<
�a<ϣa<��a<v�a<>�a<��a<��a<n�a<-�a<ڡa<��a<7�a<�a<��a<Q�a<�a<��a<\�a<�a<��a<S�a<�a<��a<�a<��a<8�a<ěa<D�a<ۚa<g�a<��a<��a<�a<��a<�a<��a<=�a<��a<J�a<֕a<Z�a<�a<��a<
�a<��a<4�a<Œa<O�a<Бa<a�a<�a<d�a<�a<�a<
�a<��a<2�a<ōa<g�a<�a<��a<H�a<�a<��a<0�a<Ɗa<b�a<�a<��a<T�a<�a<Èa<y�a<4�a<�a<��a<i�a<F�a<�a<�a<��a<��a<a�a<N�a<1�a<�a<�a<�a<�a<�a<Ņa<ąa<��a<��a<��a<��a<��a<��a<��a<ׅa<�a<�a<%�a<�  �  3�a<]�a<{�a<��a<͆a<��a<:�a<=�a<��a<��a<�a<�a<T�a<��a<�a<:�a<�a<�a<;�a<��a<�a<V�a<�a<)�a<��a<�a<b�a<؍a<?�a<��a< �a<��a<�a<��a<�a<b�a<�a<k�a<�a<p�a<�a<m�a<�a<k�a<�a<��a<�a<��a<��a<_�a<��a<H�a<ҙa<B�a<��a<1�a<��a<-�a<��a<(�a<��a<1�a<��a<	�a<��a<Пa<S�a<��a<�a<_�a<��a<�a<j�a<��a<�a<k�a<��a<�a<5�a<f�a<��a<�a<�a<K�a<��a<��a<�a<�a<2�a<��a<}�a<��a<ʦa<Ѧa<��a<��a<�a<7�a<N�a<a�a<��a<��a<��a<�a<ϧa<�a<
�a<�a<�a<�a<�a<�a<$�a<�a<�a<�a<�a<�a<اa<�a<�a<ӧa<ħa<��a<��a<z�a<k�a<L�a<<�a<�a<��a<�a<��a<��a<L�a<%�a<��a<��a<��a<r�a<G�a<�a<��a<¤a<��a<y�a<0�a<+�a<ѣa<��a<j�a< �a<�a<��a<i�a<�a<ڡa<��a<H�a<��a<��a<k�a<��a<��a<R�a<�a<��a<:�a<֝a<v�a< �a<��a<T�a<ٛa<R�a< �a<^�a<��a<x�a<�a<��a<�a<��a<,�a<Ŗa<E�a<��a<m�a<�a<��a<	�a<��a<$�a<��a<5�a<��a<K�a<ېa<f�a<�a<��a<�a<��a<G�a<͍a<h�a<��a<��a<2�a<׋a<r�a<!�a<Ίa<a�a<4�a<��a<n�a< �a<��a<}�a< �a<�a<��a<m�a<2�a<�a<�a<��a<��a<e�a<j�a<D�a<�a<�a<�a<݅a<ʅa<Åa<��a<��a<��a<��a<ǅa<��a<хa<Ʌa<܅a<�a<��a<"�a<�  �  H�a<e�a<��a<��a<݆a< �a<�a<M�a<s�a<��a<��a<�a<e�a<��a<��a<:�a<��a<��a<Q�a<��a<��a<f�a<��a<B�a<��a<�a<y�a<��a<Y�a<��a<.�a<~�a<�a<v�a<�a<o�a<בa<x�a<�a<d�a<��a<{�a<��a<�a<��a<k�a<�a<d�a<�a<g�a<ؘa<f�a<ۙa<O�a<Ěa<E�a<��a<4�a<��a<,�a<��a<�a<��a<��a<_�a<�a<@�a<��a<�a<u�a<ѡa<�a<e�a<��a<�a<5�a<��a<أa<�a<u�a<��a<�a<#�a<j�a<��a<ĥa<�a<�a<S�a<H�a<��a<��a<��a<�a<�a<�a<!�a<E�a<Y�a<n�a<��a<��a<��a<��a<�a<�a<�a<%�a<�a<.�a<+�a<.�a<(�a<,�a<�a<�a<�a<�a<�a<ڧa<ۧa<ӧa<��a<��a<��a<��a<t�a<b�a<.�a<&�a<��a<��a<��a<q�a<V�a<3�a<�a<Хa<��a<|�a<G�a<!�a<�a<ؤa<��a<i�a<A�a<�a<�a<��a<i�a<6�a<�a<��a<k�a<&�a<��a<��a<1�a<�a<��a<5�a<�a<��a<F�a<��a<��a<K�a<�a<��a<
�a<Üa<1�a<ʛa<Z�a<ݚa<|�a<�a<��a<
�a<��a<'�a<��a<<�a<ɖa<c�a<ܕa<k�a<��a<w�a<+�a<��a</�a<��a<K�a<בa<V�a<Րa<V�a<��a<d�a<�a<��a<"�a<܍a<O�a<	�a<��a<Q�a<�a<��a<%�a<ϊa<��a<��a<��a<c�a<�a<Ԉa<t�a<2�a<�a<��a<x�a<?�a<�a<�a<��a<��a<u�a<M�a<@�a<8�a< �a<�a<�a<څa<ǅa<a<��a<��a<��a<��a<��a<��a<ąa<ۅa<ԅa<�a<&�a<�  �  B�a<K�a<��a<��a<Ԇa<�a<�a<p�a<r�a<a<�a<�a<p�a<��a<��a<1�a<��a<ۉa<M�a<��a<��a<��a<��a<H�a<��a<�a<z�a<Ǎa<J�a<��a<:�a<{�a<�a<t�a<�a<}�a<͑a<r�a<֒a<w�a<�a<\�a<�a<f�a<�a<a�a<�a<h�a<��a<}�a<٘a<q�a<ʙa<R�a<Śa<H�a<śa<0�a<��a<�a<��a<�a<��a<�a<a�a<��a</�a<��a<�a<d�a<��a<�a<u�a<��a<�a<.�a<��a<ףa<�a<s�a<��a<��a<��a<S�a<�a<åa<��a<�a<X�a<P�a<��a<��a<Ŧa<�a<�a<�a<�a<H�a<O�a<v�a<��a<��a<ɧa<��a<��a<�a<�a<�a<�a<4�a<�a<$�a<�a<(�a<�a<�a<�a<�a<�a<Χa<֧a<ŧa<��a<��a<|�a<��a<Y�a<f�a<0�a<�a< �a<Ħa<Ȧa<q�a<c�a<(�a<��a<ۥa<��a<�a<=�a<2�a<�a<Ԥa<��a<j�a<_�a<��a<�a<��a<p�a<7�a<٢a<��a<B�a<2�a<��a<��a</�a<�a<��a<+�a<��a<��a<Y�a<�a<��a<=�a<ѝa<��a<�a<Ŝa<4�a<ޛa<p�a<ޚa<��a<�a<��a<�a<��a<+�a<��a<A�a<��a<d�a<ݕa<��a<�a<z�a<2�a<��a<9�a<��a<:�a<��a<A�a<�a<J�a<��a<\�a<�a<��a<"�a<ڍa<I�a<�a<��a<;�a<ыa<��a<.�a<��a<��a<�a<ۉa<l�a<�a<ӈa<k�a<B�a<�a<��a<n�a<G�a<�a<ކa<Άa<��a<��a<R�a<>�a<2�a< �a<
�a<ͅa<Ѕa<��a<��a<��a<��a<��a<��a<��a<��a<��a<ͅa<ׅa<�a<�a<�  �  H�a<Y�a<|�a<��a<ʆa<��a<*�a<O�a<��a<��a<�a<7�a<m�a<��a<
�a<J�a<��a<��a<<�a<��a<�a<`�a<؋a<-�a<��a<�a<c�a<׍a<W�a<��a<�a<��a<�a<m�a<�a<V�a<�a<R�a<ڒa<i�a<ݓa<p�a<��a<j�a<��a<{�a<�a<y�a<�a<b�a<�a<P�a<�a<Z�a<Кa<R�a<͛a<@�a<��a<?�a<��a<'�a<��a<�a<|�a<ٟa<L�a<��a<��a<p�a<��a<�a<_�a<��a<�a<H�a<�a<ϣa<�a<C�a<��a<٤a<�a<a�a<��a<��a<��a<�a<:�a<s�a<�a<��a<̦a<̦a<�a<�a<0�a<U�a<e�a<v�a<��a<��a<��a<ߧa<ާa<��a<	�a<�a<�a<�a<�a<.�a<�a<�a<�a<��a<�a<��a<קa<�a<ŧa<��a<��a<��a<��a<��a<g�a<M�a<9�a<�a<��a<צa<��a<��a<S�a<(�a<�a<إa<��a<��a<W�a<'�a<�a<äa<��a<v�a<:�a<�a<գa<��a<q�a< �a<�a<��a<S�a<�a<ˡa<e�a<(�a<�a<��a<K�a<ߟa<��a<K�a<�a<��a<K�a<ԝa<{�a<�a<��a<E�a<қa<U�a<��a<f�a<�a<��a<�a<��a<4�a<��a<A�a<ܖa<E�a<�a<j�a<��a<��a<�a<��a<.�a<��a<F�a<Ǒa<@�a<Аa<S�a<׏a<v�a<��a<��a<$�a<��a<Y�a<��a<��a<H�a<ߋa<u�a<,�a<Ɋa<i�a<%�a<��a<k�a<"�a<��a<��a<6�a<��a<Ƈa<��a<G�a< �a<�a<��a<��a<s�a<^�a<D�a<�a<�a<�a<ۅa<څa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<�a<��a<�a<�  �  "�a<f�a<t�a<��a<цa<��a<8�a<J�a<��a<��a<�a<=�a<f�a<ˈa<�a<b�a<��a<�a<U�a<��a<�a<_�a<�a<'�a<��a< �a<m�a<�a<3�a<��a<��a<��a<��a<a�a<�a<M�a<�a<:�a<��a<Q�a<�a<i�a<ߔa<��a<�a<��a<�a<~�a<��a<n�a< �a<R�a<�a<M�a<ٚa<\�a<Λa<O�a<��a<c�a<��a<6�a<��a<�a<��a<ԟa<c�a<��a<�a<^�a<��a<�a<F�a<̢a<բa<A�a<y�a<Уa<�a<@�a<��a<��a<!�a<E�a<��a<��a<�a<4�a<2�a<~�a<��a<��a<ͦa<�a<'�a<�a<H�a<A�a<y�a<x�a<��a<Чa<��a<�a<ߧa<	�a<�a<�a<)�a<�a</�a<	�a<"�a< �a<�a<�a<ܧa<��a<ħa<ߧa<��a<��a<��a<��a<��a<i�a<u�a<E�a<:�a<�a<�a<�a<��a<��a<O�a<N�a<�a<ѥa<ťa<u�a<o�a<�a<�a<ܤa<��a<��a<9�a<)�a<ϣa<��a<e�a<*�a<�a<��a<j�a<��a<�a<m�a<�a<�a<x�a<C�a<ǟa<��a<4�a<�a<��a<+�a<�a<h�a<3�a<��a<K�a<ߛa<b�a<�a<h�a<4�a<��a<�a<��a<4�a<Ɨa<4�a<�a<P�a<��a<y�a<
�a<��a<�a<��a<�a<��a<4�a<��a<L�a<��a<x�a<��a<o�a<��a<��a<�a<��a<z�a<׌a<��a<,�a<��a<��a<�a<�a<a�a<0�a<��a<{�a<#�a<Јa<��a<(�a<�a<��a<��a<I�a<!�a<�a<��a<��a<u�a<n�a<A�a<#�a<�a<�a<�a<��a<��a<��a<��a<��a<w�a<��a<|�a<��a<��a<Ʌa<�a<��a<#�a<�  �  (�a<X�a<|�a<��a<Ԇa<��a<-�a<q�a<��a<Ǉa<�a<0�a<y�a<͈a< �a<h�a<��a<��a<c�a<��a<�a<��a<ыa<9�a<��a<�a<k�a<эa</�a<��a<��a<|�a<�a<^�a<ېa<\�a<ϑa<G�a<ےa<;�a<ޓa<Y�a<ܔa<w�a<�a<x�a< �a<r�a<�a<��a<�a<r�a<�a<W�a<�a<\�a<ћa<V�a<��a<@�a<��a<'�a<��a<�a<p�a<�a<K�a<��a<�a<T�a<��a<�a<5�a<��a<�a</�a<�a<£a< �a<K�a<��a<��a<�a<;�a<��a<��a<ܥa<�a<D�a<g�a<��a<��a<˦a<��a<�a<�a<P�a<M�a<x�a<��a<��a<��a<ͧa<קa<�a<��a<�a<�a<�a<�a<"�a<�a<�a<�a<�a<��a<�a<ߧa<�a<ɧa<��a<��a<��a<��a<��a<o�a<g�a<N�a<2�a<�a<��a<ڦa<ɦa<��a<h�a<I�a<�a<�a<ȥa<��a<u�a<2�a<�a<�a<��a<��a<^�a<�a<�a<��a<Z�a<(�a<�a<��a<\�a<��a<��a<q�a<�a<Рa<��a<,�a<ԟa<��a<�a<�a<��a<)�a<�a<q�a<�a<��a<>�a<�a<z�a<��a<��a<�a<��a<(�a<��a<8�a<͗a<H�a<ݖa<j�a<�a<��a<�a<��a< �a<��a<"�a<��a<*�a<��a<?�a<��a<T�a<͏a<^�a<��a<��a<�a<��a<P�a<֌a<��a<"�a<Ӌa<|�a<�a<͊a<s�a<�a<݉a<�a<!�a<�a<��a<@�a<�a<��a<��a<U�a<�a<�a<҆a<��a<��a<e�a<;�a<-�a<	�a<�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<Ņa<�a<�a<�  �  I�a<C�a<��a<��a<Άa<�a<�a<i�a<{�a<�a<��a<I�a<��a<��a<,�a<J�a<��a<��a<c�a<Ŋa<��a<v�a<ċa<N�a<��a<�a<b�a<ɍa<O�a<��a<�a<k�a<�a<Z�a<ɐa<R�a<��a<R�a<��a<X�a<Փa<`�a<��a<U�a<
�a<`�a<�a<��a<��a<z�a<�a<��a<ߙa<��a<ښa<h�a<�a<A�a<�a<4�a<ӝa<$�a<��a<�a<y�a<�a</�a<��a<�a<k�a<��a<��a<U�a<��a<�a<�a<w�a<��a<��a<?�a<v�a<٤a<��a<X�a<��a<��a<��a<�a<X�a<_�a<��a<��a<ۦa<�a<�a<9�a</�a<x�a<u�a<��a<��a<��a<�a<ŧa<��a<�a<�a<�a<�a<,�a<�a<0�a<�a<�a<��a<ߧa<�a<ħa<ѧa<��a<��a<��a<��a<��a<r�a<��a<R�a<Z�a<5�a<�a<�a<˦a<¦a<z�a<��a<6�a<�a<�a<��a<��a<W�a<J�a<�a<�a<��a<m�a<P�a<�a<��a<��a<x�a< �a<ۢa<��a<>�a<�a<��a<_�a<�a<��a<}�a<�a<��a<o�a<;�a<ޞa<��a<H�a<��a<��a<��a<��a<M�a<ԛa<m�a<�a<��a<�a<��a< �a<��a<M�a<��a<n�a<іa<��a<�a<|�a<	�a<��a<)�a<��a<A�a<��a<A�a<��a<1�a<Őa</�a<ҏa<M�a<�a<x�a<	�a<��a<6�a<��a<y�a<?�a<؋a<n�a<7�a<��a<��a<�a<Ήa<h�a<0�a<�a<��a<^�a<��a<�a<��a<`�a<;�a<�a<�a<��a<��a<T�a<S�a<*�a<�a<�a<ąa<܅a<��a<��a<��a<t�a<��a<k�a<��a<}�a<��a<��a<Ʌa<�a<��a<�  �  &�a<<�a<��a<��a<ˆa<�a<6�a<q�a<��a<߇a<��a<W�a<��a<ǈa<�a<X�a<��a<�a<V�a<ʊa<!�a<��a<�a<G�a<��a<�a<f�a<Ía<1�a<��a<�a<|�a<��a<S�a<ϐa<N�a<��a<F�a<Òa<Y�a<˓a<S�a<ߔa<M�a<�a<y�a<��a<��a<
�a<��a<�a<��a<�a<��a<ݚa<g�a<�a<H�a<�a<>�a<ĝa<<�a<��a<"�a<��a<�a<C�a<��a<�a<T�a<��a<�a<V�a<��a<ޢa<"�a<r�a<��a<��a<<�a<��a<ˤa<��a<?�a<w�a<��a< �a<�a<P�a<z�a<��a<Ħa<�a<�a<�a<?�a<;�a<f�a<x�a<��a<��a<��a<�a<�a<�a<�a<�a<�a<#�a<&�a<��a<�a<�a<��a<�a<�a<�a<Чa<ͧa<��a<��a<��a<��a<��a<s�a<m�a<K�a<U�a<@�a<�a<�a<�a<ɦa<��a<�a<5�a<.�a<��a<��a<��a<d�a<N�a<�a<ݤa<Ǥa<��a<]�a<$�a<�a<��a<}�a<#�a<բa<��a<:�a<�a<��a<^�a<�a<àa<y�a<�a<ӟa<|�a<;�a<Ԟa<�a<+�a<��a<��a<�a<��a<P�a<�a<��a<�a<��a<�a<��a<#�a<��a<I�a<��a<m�a<ۖa<v�a<�a<��a<�a<��a<�a<��a<9�a<��a<*�a<��a<,�a<ǐa<>�a<ɏa<Q�a<�a<w�a<�a<��a<H�a<�a<u�a<&�a<ɋa<m�a<8�a<��a<�a<,�a<܉a<��a<<�a<݈a<��a<d�a<�a<ׇa<��a<d�a<H�a<�a<�a<��a<��a<m�a<R�a<$�a<�a<��a<��a<��a<��a<��a<��a<y�a<}�a<x�a<��a<��a<��a<��a<хa<�a<��a<�  �  �a<i�a<x�a<��a<׆a<��a<0�a<[�a<��a<̇a<�a<S�a<��a<�a<�a<��a<��a<�a<i�a<��a<�a<s�a<ҋa<2�a<��a<��a<o�a<ۍa<"�a<��a<��a<p�a<ۏa<H�a<Ða<>�a<��a<3�a<ɒa<A�a<��a<\�a<ݔa<��a<��a<|�a<��a<p�a<��a<s�a<��a<}�a<��a<w�a<�a<u�a<�a<z�a<לa<R�a<ŝa<2�a<��a<
�a<s�a<ܟa<R�a<��a<�a<Y�a<��a<�a<:�a<��a<͢a<�a<^�a<��a<�a<1�a<|�a<��a<�a<4�a<��a<ťa<ޥa<"�a<@�a<h�a<��a<��a<ئa< �a<�a<4�a<o�a<U�a<��a<��a<��a<̧a<Чa<�a<�a< �a<�a<�a<�a<�a<1�a< �a<�a< �a<�a<�a<̧a<Χa<§a<��a<��a<��a<��a<��a<��a<]�a<w�a<J�a<4�a<�a<��a<ݦa<��a<��a<m�a<T�a<*�a<�a<�a<��a<��a<J�a< �a<�a<��a<��a<N�a<�a<ڣa<��a<\�a<-�a<�a<��a<_�a<�a<��a<X�a<�a<��a<i�a<�a<��a<��a<#�a<�a<��a<)�a<�a<f�a<�a<��a<<�a<֛a<f�a<�a<��a<#�a<��a<L�a<˘a<M�a<�a<a�a<�a<w�a<��a<|�a<�a<��a<�a<��a<�a<Œa</�a<��a<G�a<��a<>�a<��a<K�a<Ԏa<f�a<��a<��a<=�a<̌a<��a<�a<ًa<��a<�a<ӊa<o�a<�a<ˉa<�a<.�a<�a<��a<Y�a<8�a<Ƈa<��a<u�a<=�a<�a<Նa<��a<��a<f�a<=�a<*�a<�a<�a<��a<��a<��a<��a<��a<~�a<h�a<v�a<{�a<��a<��a<��a<Åa<ޅa<�a<�  �  �a<H�a<n�a<��a<ۆa<�a<A�a<u�a<��a<��a<�a<N�a<��a<ֈa<�a<o�a<��a<�a<g�a<Ίa<�a<��a<�a<E�a<��a<��a<[�a<��a<�a<��a<��a<o�a<�a<]�a<Ða<B�a<��a<G�a<Ēa<G�a<ȓa<F�a<̔a<h�a<�a<t�a<�a<��a<�a<��a<
�a<��a<��a<o�a<�a<n�a<�a<`�a<ќa<O�a<ԝa<F�a<��a<#�a<��a<�a<J�a<��a<��a<D�a<��a<�a<>�a<��a<�a< �a<f�a<��a<��a<@�a<z�a<��a<��a<(�a<r�a<��a<ݥa<�a<P�a<y�a<��a<Ħa<�a<�a<�a<.�a<T�a<d�a<��a<��a<��a<ʧa<�a<�a<�a<�a<�a<�a<�a<�a<�a<��a<��a<��a<��a<�a<�a<Ƨa<��a<��a<��a<��a<��a<��a<q�a<[�a<W�a<@�a</�a<$�a<�a<�a<ͦa<��a<��a<Q�a<%�a<�a<ѥa<��a<|�a<@�a<�a<�a<ʤa<��a<h�a<&�a<�a<��a<Z�a<�a<Ңa<}�a<<�a<�a<��a<c�a<�a<��a<m�a<�a<ԟa<}�a<)�a<Оa<q�a<�a<ҝa<i�a<�a<��a<^�a<�a<|�a<�a<��a< �a<��a<5�a<Ęa<K�a<ؗa<[�a<�a<��a<�a<��a<�a<��a<%�a<��a<�a<��a<�a<��a<&�a<��a<7�a<ˏa<O�a<ݎa<m�a<�a<��a<;�a<Ռa<w�a<�a<ŋa<n�a<�a<Њa<�a<*�a<�a<��a<B�a<�a<��a<S�a<�a<Շa<��a<c�a<6�a<�a<�a<��a<��a<v�a<W�a<3�a<�a<�a<υa<��a<��a<��a<��a<~�a<|�a<m�a<x�a<z�a<��a<��a<Ņa<مa<��a<�  �  H�a<B�a<��a<��a<Ɔa<��a<,�a<u�a<��a<�a<�a<i�a<��a<Јa<9�a<a�a<͉a<$�a<R�a<Њa<�a<��a<ыa<8�a<��a<�a<k�a<΍a<N�a<��a<�a<]�a<ɏa<G�a<��a<?�a<��a<B�a<��a<E�a<��a<g�a<�a<Y�a<�a<x�a<�a<�a<��a<��a<��a<�a<��a<��a<�a<y�a<�a<Y�a<��a<O�a<��a<5�a<��a<�a<�a<ߟa<H�a<��a<�a<`�a<��a<�a<G�a<o�a<٢a<�a<_�a<��a<�a<'�a<h�a<ˤa<�a<Y�a<��a<��a<�a<�a<D�a<k�a<��a<��a<�a<�a<*�a<R�a<E�a<��a<��a<��a<ʧa<��a<�a<�a<�a<��a<�a<
�a< �a<.�a<�a<2�a<�a<��a<�a<ħa<ާa<��a<ȧa<��a<��a<��a<��a<��a<~�a<��a<Q�a<\�a<D�a<�a<��a<٦a<Φa<��a<��a<A�a<@�a<�a<ʥa<��a<m�a<\�a<1�a<٤a<ͤa<�a<`�a<�a<�a<��a<|�a<(�a<�a<��a<;�a<�a<��a<F�a<�a<��a<i�a<�a<ϟa<[�a<'�a<ɞa<��a<>�a<Ýa<��a<�a<��a<K�a<ڛa<}�a< �a<��a<�a<˙a<8�a<Ϙa<Z�a<їa<��a<�a<n�a<��a<��a<�a<��a<�a<��a<A�a<��a<6�a<��a< �a<��a<�a<ďa<@�a<Վa<\�a<��a<��a<(�a<�a<s�a<@�a<ًa<p�a<8�a<Ɗa<s�a<�a<ىa<y�a<9�a<Ոa<��a<w�a<�a<�a<��a<s�a<R�a<��a<�a<��a<��a<c�a<F�a<�a<�a<�a<Ņa<ޅa<��a<��a<}�a<Y�a<z�a<g�a<��a<q�a<��a<��a<��a<ޅa<�a<�  �  �a<H�a<n�a<��a<ۆa<�a<A�a<u�a<��a<��a<�a<N�a<��a<ֈa<�a<o�a<��a<�a<g�a<Ίa<�a<��a<�a<E�a<��a<��a<[�a<��a<�a<��a<��a<o�a<�a<]�a<Ða<B�a<��a<G�a<Ēa<G�a<ȓa<F�a<̔a<h�a<�a<t�a<�a<��a<�a<��a<
�a<��a<��a<o�a<�a<n�a<�a<`�a<ќa<O�a<ԝa<F�a<��a<#�a<��a<�a<J�a<��a<��a<D�a<��a<�a<>�a<��a<�a< �a<f�a<��a<��a<@�a<z�a<��a<��a<(�a<r�a<��a<ݥa<�a<P�a<y�a<��a<Ħa<�a<�a<�a<.�a<T�a<d�a<��a<��a<��a<ʧa<�a<�a<�a<�a<�a<�a<�a<�a<�a<��a<��a<��a<��a<�a<�a<Ƨa<��a<��a<��a<��a<��a<��a<q�a<[�a<W�a<@�a</�a<$�a<�a<�a<ͦa<��a<��a<Q�a<%�a<�a<ѥa<��a<|�a<@�a<�a<�a<ʤa<��a<h�a<&�a<�a<��a<Z�a<�a<Ңa<}�a<<�a<�a<��a<c�a<�a<��a<m�a<�a<ԟa<}�a<)�a<Оa<q�a<�a<ҝa<i�a<�a<��a<^�a<�a<|�a<�a<��a< �a<��a<5�a<Ęa<K�a<ؗa<[�a<�a<��a<�a<��a<�a<��a<%�a<��a<�a<��a<�a<��a<&�a<��a<7�a<ˏa<O�a<ݎa<m�a<�a<��a<;�a<Ռa<w�a<�a<ŋa<n�a<�a<Њa<�a<*�a<�a<��a<B�a<�a<��a<S�a<�a<Շa<��a<c�a<6�a<�a<�a<��a<��a<v�a<W�a<3�a<�a<�a<υa<��a<��a<��a<��a<~�a<|�a<m�a<x�a<z�a<��a<��a<Ņa<مa<��a<�  �  �a<i�a<x�a<��a<׆a<��a<0�a<[�a<��a<̇a<�a<S�a<��a<�a<�a<��a<��a<�a<i�a<��a<�a<s�a<ҋa<2�a<��a<��a<o�a<ۍa<"�a<��a<��a<p�a<ۏa<H�a<Ða<>�a<��a<3�a<ɒa<A�a<��a<\�a<ݔa<��a<��a<|�a<��a<p�a<��a<s�a<��a<}�a<��a<w�a<�a<u�a<�a<z�a<לa<R�a<ŝa<2�a<��a<
�a<s�a<ܟa<R�a<��a<�a<Y�a<��a<�a<:�a<��a<͢a<�a<^�a<��a<�a<1�a<|�a<��a<�a<4�a<��a<ťa<ޥa<"�a<@�a<h�a<��a<��a<ئa< �a<�a<4�a<o�a<U�a<��a<��a<��a<̧a<Чa<�a<�a< �a<�a<�a<�a<�a<1�a< �a<�a< �a<�a<�a<̧a<Χa<§a<��a<��a<��a<��a<��a<��a<]�a<w�a<J�a<4�a<�a<��a<ݦa<��a<��a<m�a<T�a<*�a<�a<�a<��a<��a<J�a< �a<�a<��a<��a<N�a<�a<ڣa<��a<\�a<-�a<�a<��a<_�a<�a<��a<X�a<�a<��a<i�a<�a<��a<��a<#�a<�a<��a<)�a<�a<f�a<�a<��a<<�a<֛a<f�a<�a<��a<#�a<��a<L�a<˘a<M�a<�a<a�a<�a<w�a<��a<|�a<�a<��a<�a<��a<�a<Œa</�a<��a<G�a<��a<>�a<��a<K�a<Ԏa<f�a<��a<��a<=�a<̌a<��a<�a<ًa<��a<�a<ӊa<o�a<�a<ˉa<�a<.�a<�a<��a<Y�a<8�a<Ƈa<��a<u�a<=�a<�a<Նa<��a<��a<f�a<=�a<*�a<�a<�a<��a<��a<��a<��a<��a<~�a<h�a<v�a<{�a<��a<��a<��a<Åa<ޅa<�a<�  �  &�a<<�a<��a<��a<ˆa<�a<6�a<q�a<��a<߇a<��a<W�a<��a<ǈa<�a<X�a<��a<�a<V�a<ʊa<!�a<��a<�a<G�a<��a<�a<f�a<Ía<1�a<��a<�a<|�a<��a<S�a<ϐa<N�a<��a<F�a<Òa<Y�a<˓a<S�a<ߔa<M�a<�a<y�a<��a<��a<
�a<��a<�a<��a<�a<��a<ݚa<g�a<�a<H�a<�a<>�a<ĝa<<�a<��a<"�a<��a<�a<C�a<��a<�a<T�a<��a<�a<V�a<��a<ޢa<"�a<r�a<��a<��a<<�a<��a<ˤa<��a<?�a<w�a<��a< �a<�a<P�a<z�a<��a<Ħa<�a<�a<�a<?�a<;�a<f�a<x�a<��a<��a<��a<�a<�a<�a<�a<�a<�a<#�a<&�a<��a<�a<�a<��a<�a<�a<�a<Чa<ͧa<��a<��a<��a<��a<��a<s�a<m�a<K�a<U�a<@�a<�a<�a<�a<ɦa<��a<�a<5�a<.�a<��a<��a<��a<d�a<N�a<�a<ݤa<Ǥa<��a<]�a<$�a<�a<��a<}�a<#�a<բa<��a<:�a<�a<��a<^�a<�a<àa<y�a<�a<ӟa<|�a<;�a<Ԟa<�a<+�a<��a<��a<�a<��a<P�a<�a<��a<�a<��a<�a<��a<#�a<��a<I�a<��a<m�a<ۖa<v�a<�a<��a<�a<��a<�a<��a<9�a<��a<*�a<��a<,�a<ǐa<>�a<ɏa<Q�a<�a<w�a<�a<��a<H�a<�a<u�a<&�a<ɋa<m�a<8�a<��a<�a<,�a<܉a<��a<<�a<݈a<��a<d�a<�a<ׇa<��a<d�a<H�a<�a<�a<��a<��a<m�a<R�a<$�a<�a<��a<��a<��a<��a<��a<��a<y�a<}�a<x�a<��a<��a<��a<��a<хa<�a<��a<�  �  I�a<C�a<��a<��a<Άa<�a<�a<i�a<{�a<�a<��a<I�a<��a<��a<,�a<J�a<��a<��a<c�a<Ŋa<��a<v�a<ċa<N�a<��a<�a<b�a<ɍa<O�a<��a<�a<k�a<�a<Z�a<ɐa<R�a<��a<R�a<��a<X�a<Փa<`�a<��a<U�a<
�a<`�a<�a<��a<��a<z�a<�a<��a<ߙa<��a<ښa<h�a<�a<A�a<�a<4�a<ӝa<$�a<��a<�a<y�a<�a</�a<��a<�a<k�a<��a<��a<U�a<��a<�a<�a<w�a<��a<��a<?�a<v�a<٤a<��a<X�a<��a<��a<��a<�a<X�a<_�a<��a<��a<ۦa<�a<�a<9�a</�a<x�a<u�a<��a<��a<��a<�a<ŧa<��a<�a<�a<�a<�a<,�a<�a<0�a<�a<�a<��a<ߧa<�a<ħa<ѧa<��a<��a<��a<��a<��a<r�a<��a<R�a<Z�a<5�a<�a<�a<˦a<¦a<z�a<��a<6�a<�a<�a<��a<��a<W�a<J�a<�a<�a<��a<m�a<P�a<�a<��a<��a<x�a< �a<ۢa<��a<>�a<�a<��a<_�a<�a<��a<}�a<�a<��a<o�a<;�a<ޞa<��a<H�a<��a<��a<��a<��a<M�a<ԛa<m�a<�a<��a<�a<��a< �a<��a<M�a<��a<n�a<іa<��a<�a<|�a<	�a<��a<)�a<��a<A�a<��a<A�a<��a<1�a<Őa</�a<ҏa<M�a<�a<x�a<	�a<��a<6�a<��a<y�a<?�a<؋a<n�a<7�a<��a<��a<�a<Ήa<h�a<0�a<�a<��a<^�a<��a<�a<��a<`�a<;�a<�a<�a<��a<��a<T�a<S�a<*�a<�a<�a<ąa<܅a<��a<��a<��a<t�a<��a<k�a<��a<}�a<��a<��a<Ʌa<�a<��a<�  �  (�a<X�a<|�a<��a<Ԇa<��a<-�a<q�a<��a<Ǉa<�a<0�a<y�a<͈a< �a<h�a<��a<��a<c�a<��a<�a<��a<ыa<9�a<��a<�a<k�a<эa</�a<��a<��a<|�a<�a<^�a<ېa<\�a<ϑa<G�a<ےa<;�a<ޓa<Y�a<ܔa<w�a<�a<x�a< �a<r�a<�a<��a<�a<r�a<�a<W�a<�a<\�a<ћa<V�a<��a<@�a<��a<'�a<��a<�a<p�a<�a<K�a<��a<�a<T�a<��a<�a<5�a<��a<�a</�a<�a<£a< �a<K�a<��a<��a<�a<;�a<��a<��a<ܥa<�a<D�a<g�a<��a<��a<˦a<��a<�a<�a<P�a<M�a<x�a<��a<��a<��a<ͧa<קa<�a<��a<�a<�a<�a<�a<"�a<�a<�a<�a<�a<��a<�a<ߧa<�a<ɧa<��a<��a<��a<��a<��a<o�a<g�a<N�a<2�a<�a<��a<ڦa<ɦa<��a<h�a<I�a<�a<�a<ȥa<��a<u�a<2�a<�a<�a<��a<��a<^�a<�a<�a<��a<Z�a<(�a<�a<��a<\�a<��a<��a<q�a<�a<Рa<��a<,�a<ԟa<��a<�a<�a<��a<)�a<�a<q�a<�a<��a<>�a<�a<z�a<��a<��a<�a<��a<(�a<��a<8�a<͗a<H�a<ݖa<j�a<�a<��a<�a<��a< �a<��a<"�a<��a<*�a<��a<?�a<��a<T�a<͏a<^�a<��a<��a<�a<��a<P�a<֌a<��a<"�a<Ӌa<|�a<�a<͊a<s�a<�a<݉a<�a<!�a<�a<��a<@�a<�a<��a<��a<U�a<�a<�a<҆a<��a<��a<e�a<;�a<-�a<	�a<�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<Ņa<�a<�a<�  �  "�a<f�a<t�a<��a<цa<��a<8�a<J�a<��a<��a<�a<=�a<f�a<ˈa<�a<b�a<��a<�a<U�a<��a<�a<_�a<�a<'�a<��a< �a<m�a<�a<3�a<��a<��a<��a<��a<a�a<�a<M�a<�a<:�a<��a<Q�a<�a<i�a<ߔa<��a<�a<��a<�a<~�a<��a<n�a< �a<R�a<�a<M�a<ٚa<\�a<Λa<O�a<��a<c�a<��a<6�a<��a<�a<��a<ԟa<c�a<��a<�a<^�a<��a<�a<F�a<̢a<բa<A�a<y�a<Уa<�a<@�a<��a<��a<!�a<E�a<��a<��a<�a<4�a<2�a<~�a<��a<��a<ͦa<�a<'�a<�a<H�a<A�a<y�a<x�a<��a<Чa<��a<�a<ߧa<	�a<�a<�a<)�a<�a</�a<	�a<"�a< �a<�a<�a<ܧa<��a<ħa<ߧa<��a<��a<��a<��a<��a<i�a<u�a<E�a<:�a<�a<�a<�a<��a<��a<O�a<N�a<�a<ѥa<ťa<u�a<o�a<�a<�a<ܤa<��a<��a<9�a<)�a<ϣa<��a<e�a<*�a<�a<��a<j�a<��a<�a<m�a<�a<�a<x�a<C�a<ǟa<��a<4�a<�a<��a<+�a<�a<h�a<3�a<��a<K�a<ߛa<b�a<�a<h�a<4�a<��a<�a<��a<4�a<Ɨa<4�a<�a<P�a<��a<y�a<
�a<��a<�a<��a<�a<��a<4�a<��a<L�a<��a<x�a<��a<o�a<��a<��a<�a<��a<z�a<׌a<��a<,�a<��a<��a<�a<�a<a�a<0�a<��a<{�a<#�a<Јa<��a<(�a<�a<��a<��a<I�a<!�a<�a<��a<��a<u�a<n�a<A�a<#�a<�a<�a<�a<��a<��a<��a<��a<��a<w�a<��a<|�a<��a<��a<Ʌa<�a<��a<#�a<�  �  H�a<Y�a<|�a<��a<ʆa<��a<*�a<O�a<��a<��a<�a<7�a<m�a<��a<
�a<J�a<��a<��a<<�a<��a<�a<`�a<؋a<-�a<��a<�a<c�a<׍a<W�a<��a<�a<��a<�a<m�a<�a<V�a<�a<R�a<ڒa<i�a<ݓa<p�a<��a<j�a<��a<{�a<�a<y�a<�a<b�a<�a<P�a<�a<Z�a<Кa<R�a<͛a<@�a<��a<?�a<��a<'�a<��a<�a<|�a<ٟa<L�a<��a<��a<p�a<��a<�a<_�a<��a<�a<H�a<�a<ϣa<�a<C�a<��a<٤a<�a<a�a<��a<��a<��a<�a<:�a<s�a<�a<��a<̦a<̦a<�a<�a<0�a<U�a<e�a<v�a<��a<��a<��a<ߧa<ާa<��a<	�a<�a<�a<�a<�a<.�a<�a<�a<�a<��a<�a<��a<קa<�a<ŧa<��a<��a<��a<��a<��a<g�a<M�a<9�a<�a<��a<צa<��a<��a<S�a<(�a<�a<إa<��a<��a<W�a<'�a<�a<äa<��a<v�a<:�a<�a<գa<��a<q�a< �a<�a<��a<S�a<�a<ˡa<e�a<(�a<�a<��a<K�a<ߟa<��a<K�a<�a<��a<K�a<ԝa<{�a<�a<��a<E�a<қa<U�a<��a<f�a<�a<��a<�a<��a<4�a<��a<A�a<ܖa<E�a<�a<j�a<��a<��a<�a<��a<.�a<��a<F�a<Ǒa<@�a<Аa<S�a<׏a<v�a<��a<��a<$�a<��a<Y�a<��a<��a<H�a<ߋa<u�a<,�a<Ɋa<i�a<%�a<��a<k�a<"�a<��a<��a<6�a<��a<Ƈa<��a<G�a< �a<�a<��a<��a<s�a<^�a<D�a<�a<�a<�a<ۅa<څa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<�a<��a<�a<�  �  B�a<K�a<��a<��a<Ԇa<�a<�a<p�a<r�a<a<�a<�a<p�a<��a<��a<1�a<��a<ۉa<M�a<��a<��a<��a<��a<H�a<��a<�a<z�a<Ǎa<J�a<��a<:�a<{�a<�a<t�a<�a<}�a<͑a<r�a<֒a<w�a<�a<\�a<�a<f�a<�a<a�a<�a<h�a<��a<}�a<٘a<q�a<ʙa<R�a<Śa<H�a<śa<0�a<��a<�a<��a<�a<��a<�a<a�a<��a</�a<��a<�a<d�a<��a<�a<u�a<��a<�a<.�a<��a<ףa<�a<s�a<��a<��a<��a<S�a<�a<åa<��a<�a<X�a<P�a<��a<��a<Ŧa<�a<�a<�a<�a<H�a<O�a<v�a<��a<��a<ɧa<��a<��a<�a<�a<�a<�a<4�a<�a<$�a<�a<(�a<�a<�a<�a<�a<�a<Χa<֧a<ŧa<��a<��a<|�a<��a<Y�a<f�a<0�a<�a< �a<Ħa<Ȧa<q�a<c�a<(�a<��a<ۥa<��a<�a<=�a<2�a<�a<Ԥa<��a<j�a<_�a<��a<�a<��a<p�a<7�a<٢a<��a<B�a<2�a<��a<��a</�a<�a<��a<+�a<��a<��a<Y�a<�a<��a<=�a<ѝa<��a<�a<Ŝa<4�a<ޛa<p�a<ޚa<��a<�a<��a<�a<��a<+�a<��a<A�a<��a<d�a<ݕa<��a<�a<z�a<2�a<��a<9�a<��a<:�a<��a<A�a<�a<J�a<��a<\�a<�a<��a<"�a<ڍa<I�a<�a<��a<;�a<ыa<��a<.�a<��a<��a<�a<ۉa<l�a<�a<ӈa<k�a<B�a<�a<��a<n�a<G�a<�a<ކa<Άa<��a<��a<R�a<>�a<2�a< �a<
�a<ͅa<Ѕa<��a<��a<��a<��a<��a<��a<��a<��a<��a<ͅa<ׅa<�a<�a<�  �  H�a<e�a<��a<��a<݆a< �a<�a<M�a<s�a<��a<��a<�a<e�a<��a<��a<:�a<��a<��a<Q�a<��a<��a<f�a<��a<B�a<��a<�a<y�a<��a<Y�a<��a<.�a<~�a<�a<v�a<�a<o�a<בa<x�a<�a<d�a<��a<{�a<��a<�a<��a<k�a<�a<d�a<�a<g�a<ؘa<f�a<ۙa<O�a<Ěa<E�a<��a<4�a<��a<,�a<��a<�a<��a<��a<_�a<�a<@�a<��a<�a<u�a<ѡa<�a<e�a<��a<�a<5�a<��a<أa<�a<u�a<��a<�a<#�a<j�a<��a<ĥa<�a<�a<S�a<H�a<��a<��a<��a<�a<�a<�a<!�a<E�a<Y�a<n�a<��a<��a<��a<��a<�a<�a<�a<%�a<�a<.�a<+�a<.�a<(�a<,�a<�a<�a<�a<�a<�a<ڧa<ۧa<ӧa<��a<��a<��a<��a<t�a<b�a<.�a<&�a<��a<��a<��a<q�a<V�a<3�a<�a<Хa<��a<|�a<G�a<!�a<�a<ؤa<��a<i�a<A�a<�a<�a<��a<i�a<6�a<�a<��a<k�a<&�a<��a<��a<1�a<�a<��a<5�a<�a<��a<F�a<��a<��a<K�a<�a<��a<
�a<Üa<1�a<ʛa<Z�a<ݚa<|�a<�a<��a<
�a<��a<'�a<��a<<�a<ɖa<c�a<ܕa<k�a<��a<w�a<+�a<��a</�a<��a<K�a<בa<V�a<Րa<V�a<��a<d�a<�a<��a<"�a<܍a<O�a<	�a<��a<Q�a<�a<��a<%�a<ϊa<��a<��a<��a<c�a<�a<Ԉa<t�a<2�a<�a<��a<x�a<?�a<�a<�a<��a<��a<u�a<M�a<@�a<8�a< �a<�a<�a<څa<ǅa<a<��a<��a<��a<��a<��a<��a<ąa<ۅa<ԅa<�a<&�a<�  �  3�a<]�a<{�a<��a<͆a<��a<:�a<=�a<��a<��a<�a<�a<T�a<��a<�a<:�a<�a<�a<;�a<��a<�a<V�a<�a<)�a<��a<�a<b�a<؍a<?�a<��a< �a<��a<�a<��a<�a<b�a<�a<k�a<�a<p�a<�a<m�a<�a<k�a<�a<��a<�a<��a<��a<_�a<��a<H�a<ҙa<B�a<��a<1�a<��a<-�a<��a<(�a<��a<1�a<��a<	�a<��a<Пa<S�a<��a<�a<_�a<��a<�a<j�a<��a<�a<k�a<��a<�a<5�a<f�a<��a<�a<�a<K�a<��a<��a<�a<�a<2�a<��a<}�a<��a<ʦa<Ѧa<��a<��a<�a<7�a<N�a<a�a<��a<��a<��a<�a<ϧa<�a<
�a<�a<�a<�a<�a<�a<$�a<�a<�a<�a<�a<�a<اa<�a<�a<ӧa<ħa<��a<��a<z�a<k�a<L�a<<�a<�a<��a<�a<��a<��a<L�a<%�a<��a<��a<��a<r�a<G�a<�a<��a<¤a<��a<y�a<0�a<+�a<ѣa<��a<j�a< �a<�a<��a<i�a<�a<ڡa<��a<H�a<��a<��a<k�a<��a<��a<R�a<�a<��a<:�a<֝a<v�a< �a<��a<T�a<ٛa<R�a< �a<^�a<��a<x�a<�a<��a<�a<��a<,�a<Ŗa<E�a<��a<m�a<�a<��a<	�a<��a<$�a<��a<5�a<��a<K�a<ېa<f�a<�a<��a<�a<��a<G�a<͍a<h�a<��a<��a<2�a<׋a<r�a<!�a<Ίa<a�a<4�a<��a<n�a< �a<��a<}�a< �a<�a<��a<m�a<2�a<�a<�a<��a<��a<e�a<j�a<D�a<�a<�a<�a<݅a<ʅa<Åa<��a<��a<��a<��a<ǅa<��a<хa<Ʌa<܅a<�a<��a<"�a<�  �  O�a<m�a<��a<��a<Ɇa<�a<�a<<�a<r�a<��a<�a<"�a<i�a<��a<�a<3�a<��a<�a<A�a<��a<�a<O�a<Ƌa<'�a<��a<�a<��a<�a<R�a<��a<5�a<��a<�a<|�a<��a<n�a<�a<f�a<�a<y�a<��a<z�a<�a<~�a< �a<|�a<�a<l�a<�a<Q�a<֘a<Q�a<Ιa<P�a<͚a<;�a<��a<4�a<��a<"�a<��a<�a<y�a<�a<m�a<џa<K�a<��a<�a<y�a<ˡa<(�a<w�a<��a<��a<Q�a<��a<�a< �a<^�a<��a<�a<)�a<`�a<��a<ҥa<��a<�a<3�a<b�a<o�a<��a<��a<צa<��a<�a<�a<8�a<K�a<u�a<��a<��a<��a<��a<˧a<�a<��a<�a<!�a<,�a</�a<9�a<&�a<-�a<�a<�a<��a<�a<�a<�a<Χa<ϧa<��a<��a<��a<��a<{�a<a�a<?�a<�a<�a<Ʀa<��a<q�a<I�a<'�a<��a<ԥa<��a<p�a<@�a<"�a<��a<Ȥa<��a<\�a<)�a<
�a<ϣa<��a<v�a<>�a<��a<��a<n�a<-�a<ڡa<��a<7�a<�a<��a<Q�a<�a<��a<\�a<�a<��a<S�a<�a<��a<�a<��a<8�a<ěa<D�a<ۚa<g�a<��a<��a<�a<��a<�a<��a<=�a<��a<J�a<֕a<Z�a<�a<��a<
�a<��a<4�a<Œa<O�a<Бa<a�a<�a<d�a<�a<�a<
�a<��a<2�a<ōa<g�a<�a<��a<H�a<�a<��a<0�a<Ɗa<b�a<�a<��a<T�a<�a<Èa<y�a<4�a<�a<��a<i�a<F�a<�a<�a<��a<��a<a�a<N�a<1�a<�a<�a<�a<�a<�a<Ņa<ąa<��a<��a<��a<��a<��a<��a<��a<ׅa<�a<�a<%�a<�  �  ,�a<�a<j�a<f�a<��a<˅a<�a<,�a<4�a<��a<��a<Ԇa<&�a<R�a<��a<�a<N�a<��a<�a<d�a<��a<S�a<��a<�a<g�a<؋a<c�a<��a<N�a<�a<�a<��a<��a<m�a<��a<��a<ېa<x�a<ޑa<t�a<�a<r�a<	�a<m�a<�a<`�a<��a<l�a<��a<g�a<̗a<f�a<Θa<<�a<��a<)�a<��a<*�a<��a<-�a<��a<�a<��a<,�a<��a<
�a<S�a<ԟa<1�a<��a<��a<<�a<��a<�a<F�a<q�a<�a<�a<G�a<��a<ѣa<�a<,�a<��a<��a<�a<�a<*�a<r�a<w�a<��a<��a<ɥa<�a<��a<�a<�a<6�a<M�a<{�a<��a<��a<զa<Φa<�a<�a< �a<'�a<!�a<R�a<.�a<b�a<.�a<R�a<@�a<1�a<4�a<!�a<H�a<�a<��a<�a<ܦa<ܦa<��a<��a<x�a<��a<A�a<(�a<�a<�a<Υa<|�a<i�a<6�a<�a<פa<��a<h�a<8�a<"�a<�a<ڣa<��a<p�a<n�a<�a<�a<��a<z�a<]�a<�a<�a<g�a<N�a<��a<��a<[�a<�a<�a<g�a<2�a<a<~�a< �a<a<v�a<��a<��a<�a<ʛa<L�a<�a<h�a<ۙa<��a<��a<r�a< �a<x�a<�a<��a<�a<��a<X�a<Ŕa<j�a<�a<~�a<�a<��a<*�a<��a<G�a<̐a<A�a<��a<T�a<��a<c�a<�a<��a<�a<Ìa<P�a<��a<h�a<A�a<Ċa<m�a<��a<��a<Y�a<߈a<��a<2�a<ԇa<��a<3�a<�a<��a<[�a<�a<��a<��a<��a<��a<K�a<I�a<"�a<�a<�a<Ąa<لa<��a<��a<}�a<��a<��a<w�a<��a<y�a<��a<��a<��a<��a<��a<�a<քa<�  �  �a<&�a<d�a<z�a<��a<ƅa<�a<�a<I�a<r�a<��a<�a<�a<o�a<��a<�a<M�a<��a<�a<m�a<Ήa<1�a<��a<�a<��a<�a<\�a<��a<4�a<��a<�a<}�a<��a<w�a<ۏa<M�a<ݐa<d�a<ݑa<l�a<�a<p�a<�a<u�a<�a<��a< �a<r�a<�a<f�a<�a<P�a<ۘa<A�a<��a<G�a<ƚa<5�a<��a<<�a<��a<4�a<��a<�a<��a<�a<x�a<۟a<7�a<��a<�a<D�a<��a<ܡa<4�a<y�a<��a<��a<Q�a<��a<ɣa<�a<K�a<��a<��a<�a<�a<S�a<`�a<y�a<��a<��a<إa<�a<�a<�a<3�a<V�a<j�a<t�a<��a<��a<��a<�a<�a<�a<�a<=�a<>�a<U�a<;�a<J�a<E�a<J�a<6�a<3�a</�a<�a<��a<��a<�a<�a<Ԧa<צa<��a<��a<��a<��a<V�a<D�a<�a<ߥa<��a<��a<[�a<3�a<��a<Ϥa<��a<��a<S�a< �a<��a<ѣa<��a<}�a<M�a<�a<��a<բa<��a<V�a<�a<Сa<��a<M�a<�a<��a<e�a<�a<��a<i�a<�a<��a<w�a<�a<��a<^�a<��a<��a<:�a<͛a<Q�a<ݚa<g�a<��a<l�a<�a<w�a<�a<��a<"�a<��a<$�a<ŕa<D�a<�a<j�a<�a<��a<�a<��a<0�a<��a<3�a<��a<I�a<֏a<O�a<�a<l�a<�a<}�a<$�a<��a<G�a<��a<��a<(�a<��a<j�a<	�a<��a<F�a<�a<��a<5�a<�a<��a<?�a<�a<��a<z�a<<�a<��a<ǅa<��a<v�a<b�a<:�a<�a<
�a<�a<�a<܄a<��a<��a<��a<��a<z�a<y�a<{�a<q�a<`�a<�a<��a<��a<��a<�a<�a<�  �  �a<E�a<N�a<m�a<��a<��a<�a<�a<]�a<h�a<��a<�a<�a<a�a<��a<��a<E�a<��a<��a<i�a<߉a<1�a<��a<��a<��a<׋a<S�a<֌a<+�a<��a<�a<��a<�a<o�a<��a<^�a<��a<O�a<�a<h�a<�a<x�a<�a<��a<�a<}�a<�a<{�a<��a<`�a<��a<?�a<��a<C�a<��a<8�a<��a</�a<��a<=�a<��a<9�a<��a<"�a<��a<��a<y�a<ßa<F�a<��a<�a<B�a<��a<�a<!�a<��a<��a<�a<S�a<��a<֣a<�a<S�a<�a<ɤa<�a<�a<P�a<N�a<��a<��a<åa<إa<֥a<�a<�a<)�a<5�a<Z�a<g�a<��a<��a<��a<��a<�a<�a<�a<5�a<2�a<:�a<V�a<A�a<R�a<5�a<9�a<2�a<�a<7�a<�a<"�a<�a<�a<ܦa<��a<Ȧa<��a<��a<l�a<H�a<<�a<�a<��a<��a<��a<Q�a<0�a<	�a<äa<��a<i�a<J�a<�a<��a<��a<��a<��a<M�a<B�a<�a<Ӣa<y�a<M�a<#�a<ǡa<��a<6�a<��a<��a<]�a< �a<��a<��a<	�a<˞a<s�a<�a<ȝa<_�a<�a<��a<5�a<��a<[�a<�a<a�a<�a<\�a<	�a<y�a<��a<��a<�a<��a<%�a<ƕa<.�a<�a<d�a<��a<��a<	�a<��a<�a<��a<;�a<Őa<F�a<̏a<Z�a<Ҏa<��a<��a<��a<&�a<��a<T�a<�a<��a<!�a<֊a<j�a<��a<��a<5�a<�a<��a<>�a<�a<v�a<A�a<�a<��a<Z�a<,�a<�a<υa<��a<k�a<u�a<5�a<6�a<	�a<��a<Մa<��a<ńa<��a<��a<|�a<|�a<w�a<c�a<��a<p�a<��a<��a<��a<��a<ʄa< �a<�  �  �a<.�a<W�a<z�a<��a<��a<��a<'�a<M�a<z�a<��a<�a<8�a<o�a<��a<�a<d�a<��a<�a<e�a<ډa<E�a<��a<�a<w�a<�a<Z�a<��a<-�a<��a<�a<��a<�a<I�a<��a<\�a<ːa<U�a<�a<l�a<ܒa<n�a<�a<y�a<��a<z�a<��a<b�a<��a<n�a<ޗa<`�a<ʘa<R�a<ՙa<N�a<ƚa<E�a<��a<+�a<��a<%�a<��a<.�a<��a<�a<k�a<ϟa<:�a<��a<�a<0�a<��a<�a<%�a<a�a<��a< �a<,�a<��a<٣a<�a<3�a<�a<��a<�a<�a<9�a<_�a<��a<��a<ĥa<˥a<�a<��a<+�a<7�a<P�a<k�a<��a<��a<��a<Φa<�a< �a<�a<�a</�a<9�a<B�a<D�a<F�a<:�a<1�a<A�a<2�a<�a<�a<�a<��a<٦a<�a<�a<��a<��a<��a<��a<u�a<U�a<2�a<��a<�a<ɥa<��a<d�a<0�a<�a<�a<��a<��a<V�a<8�a<��a<֣a<��a<��a<a�a<'�a<�a<��a<��a<T�a<�a<ʡa<r�a<5�a<�a<��a<7�a<�a<��a<W�a<�a<ʞa<v�a<�a<��a<]�a<�a<��a<2�a<ɛa<B�a<�a<n�a<�a<}�a<��a<��a<�a<��a<"�a<��a<7�a<��a<P�a<Ӕa<m�a<	�a<{�a<�a<��a<$�a<��a<2�a<��a<4�a<Ϗa<Y�a<֎a<T�a<�a<��a<��a<��a<W�a<�a<p�a<"�a<a<j�a<�a<��a<E�a<�a<��a<?�a<ևa<��a<9�a<�a<��a<u�a<=�a<�a<Ӆa<��a<��a<_�a<G�a</�a<��a<�a<݄a<Ʉa<��a<��a<��a<x�a<��a<x�a<\�a<h�a<v�a<{�a<s�a<��a<Ȅa<Ʉa<�a<�  �  �a<�a<_�a<z�a<��a<مa<�a<'�a<<�a<��a<��a<��a<<�a<^�a<ˇa<��a<p�a<��a<(�a<s�a<ωa<C�a<��a<*�a<x�a<�a<Y�a<��a<9�a<��a<�a<d�a<�a<k�a<֏a<[�a<Аa<i�a<đa<b�a<��a<o�a<�a<c�a<�a<u�a<�a<s�a<�a<v�a<ۗa<y�a<Ԙa<f�a<əa<?�a<��a<9�a<қa<7�a<Ҝa<(�a<��a<"�a<��a<�a<f�a<�a<(�a<��a<�a<6�a<��a<¡a<5�a<m�a<��a<��a<F�a<��a<��a<�a<@�a<��a<��a<�a<#�a<8�a<~�a<z�a<��a<��a<֥a<�a<�a<6�a<.�a<]�a<X�a<��a<��a<��a<�a<զa<�a<	�a<)�a<:�a<9�a<O�a<(�a<I�a<D�a<<�a<(�a<�a</�a<�a<	�a<�a<��a<ߦa<Ʀa<ͦa<��a<��a<o�a<|�a<U�a<:�a<!�a<ݥa<ɥa<��a<y�a<E�a<�a<�a<��a<��a<I�a<C�a< �a<�a<��a<~�a<_�a<�a<�a<��a<��a<S�a<�a<֡a<��a<G�a<נa<��a<Y�a<��a<��a<\�a<"�a<��a<l�a<�a<��a<Z�a<�a<��a<-�a<ܛa<S�a<�a<w�a<�a<��a<��a<��a<�a<��a<�a<��a<K�a<��a<l�a<֔a<u�a<��a<��a<.�a<��a<=�a<��a<(�a<a<;�a<Ϗa<6�a<�a<`�a<�a<�a<�a<��a<,�a<�a<|�a<,�a<��a<a�a<�a<��a<e�a<�a<��a<8�a<�a<��a<@�a<�a<��a<��a<*�a<�a<��a<��a<��a<R�a<N�a< �a<�a<��a<܄a<քa<��a<��a<��a<��a<l�a<e�a<|�a<]�a<r�a<l�a<��a<��a<��a<ׄa<�a<�  �  ��a<:�a<U�a<q�a<��a<Ѕa<��a<$�a<f�a<��a<��a<�a<@�a<y�a<ʇa<�a<n�a<��a<�a<��a<�a<?�a<��a<�a<|�a<܋a<T�a<ǌa<"�a<��a< �a<m�a<��a<b�a<ŏa<>�a<Ԑa<F�a<Αa<V�a<Ԓa<g�a<�a<{�a<��a<t�a<�a<��a<�a<w�a<�a<g�a<�a<b�a<ߙa<U�a<њa<R�a<͛a<F�a<��a<P�a<��a<�a<��a<��a<k�a<՟a<8�a<��a<�a<-�a<��a<ϡa<�a<l�a<��a<�a<@�a<u�a<��a< �a<8�a<u�a<��a<�a<�a<?�a<\�a<��a<��a<ӥa<��a<��a<�a<2�a<I�a<a�a<s�a<��a<��a<æa<֦a<�a<�a<�a<2�a<*�a<1�a<@�a<K�a<:�a<>�a<'�a<(�a<�a<�a<�a<��a<�a<�a<Ԧa<Ȧa<��a<��a<��a<��a<s�a<L�a<0�a<�a<��a<ƥa<��a<v�a<G�a<�a<�a<��a<��a<d�a<B�a<�a<�a<ƣa<��a<[�a<=�a<��a<¢a<~�a<M�a<�a<��a<x�a</�a<�a<��a<P�a<�a<��a<`�a< �a<��a<`�a<�a<��a<Y�a<�a<��a<,�a<��a<r�a<��a<w�a<�a<��a<�a<��a<"�a<��a<.�a<��a<F�a<ϕa<V�a<��a<{�a<��a<��a<
�a<��a<*�a<��a<3�a<��a<1�a<��a<B�a<Ŏa<_�a<֍a<d�a<�a<��a<;�a<ۋa<t�a<�a<Êa<c�a<��a<��a<B�a<�a<��a<N�a< �a<��a<K�a<�a<ņa<��a<E�a<�a<߅a<��a<��a<��a<K�a<-�a<�a<�a<Ԅa<Ǆa<��a<��a<��a<n�a<k�a<_�a<[�a<`�a<_�a<k�a<��a<��a<��a<��a<�a<�  �  �a<:�a<>�a<��a<��a<��a<�a<�a<n�a<�a<цa<��a<C�a<��a<��a<,�a<g�a<ψa<"�a<�a<�a<0�a<a<��a<��a<ߋa<J�a<��a<�a<��a<�a<r�a<ˎa<R�a<Ǐa</�a<͐a</�a<Ցa<=�a<ܒa<^�a<ϓa<~�a<ٔa<��a<�a<��a<��a<j�a<�a<`�a<��a<X�a<�a<[�a<њa<e�a<��a<_�a<��a<Q�a<��a<!�a<��a<�a<��a<��a<:�a<v�a<Ԡa<8�a<h�a<աa<��a<e�a<��a<�a<7�a<^�a<��a<ߣa<D�a<Y�a<��a<�a<�a<]�a<N�a<��a<��a<ԥa<�a<��a</�a<)�a<^�a<X�a<��a<��a<��a<Ԧa<̦a<�a<�a<#�a<!�a<3�a<Q�a<&�a<O�a<�a<?�a< �a<�a<�a<��a<�a<ݦa<�a<զa<ɦa<Ȧa<��a<��a<{�a<��a<\�a<f�a<D�a<�a<�a<��a<��a<i�a<W�a<�a<��a<Фa<��a<~�a<;�a< �a<�a<��a<��a<K�a<F�a<�a<ޢa<��a<D�a<�a<��a<��a<�a<�a<~�a<A�a<�a<��a<Y�a<�a<��a<H�a<�a<��a<=�a<�a<{�a<O�a<��a<j�a<�a<j�a<�a<}�a<'�a<��a<5�a<��a<.�a<ϖa<9�a<�a<S�a<��a<r�a<��a<��a< �a<��a<
�a<��a<�a<��a<=�a<��a<H�a<��a<W�a<ʍa<f�a<	�a<��a<>�a<��a<��a<��a<��a<d�a<�a<Ɖa<5�a<	�a<��a<O�a<��a<��a<i�a<�a<ۆa<}�a<X�a< �a<�a<˅a<��a<��a<4�a<9�a<�a<��a<�a<��a<��a<z�a<��a<g�a<b�a<Z�a<K�a<_�a<G�a<k�a<o�a<��a<��a<��a<�a<�  �  ��a<*�a<M�a<r�a<��a<օa<�a<*�a<e�a<��a<φa<�a<U�a<��a<ׇa</�a<x�a<шa<0�a<��a<�a<M�a<��a<�a<u�a<ۋa<[�a<��a<�a<��a<�a<^�a<ˎa<G�a<��a<7�a<��a<9�a<��a<;�a<ޒa<^�a<ۓa<�a<�a<z�a<��a<��a<	�a<��a<��a<��a<��a<o�a<��a<\�a<ٚa<m�a<ڛa<Z�a<՜a<F�a<��a<6�a<��a<
�a<l�a<��a<>�a<y�a<٠a<7�a<j�a<��a<�a<Q�a<��a<٢a<&�a<e�a<��a<�a<C�a<i�a<��a<�a<�a<9�a<q�a<��a<��a<ۥa<�a<�a<(�a<?�a<e�a<j�a<��a<��a<��a<Ϧa<�a<��a<
�a<-�a</�a<)�a<6�a<5�a<C�a<.�a<8�a<)�a<�a<��a<�a<�a<�a<զa<֦a<��a<��a<��a<��a<��a<��a<k�a<M�a</�a<�a<�a<̥a<��a<}�a<U�a<*�a<�a<Ϥa<��a<��a<L�a<"�a<��a<��a<��a<h�a<@�a<�a<��a<}�a<T�a<��a<��a<��a<�a<Рa<}�a<6�a<ݟa<��a<D�a<�a<��a<F�a<�a<��a<I�a<�a<��a<2�a<ƛa<g�a<��a<��a<�a<��a<#�a<��a<=�a<��a<5�a<זa<S�a<�a<p�a<��a<��a<�a<��a<�a<��a<�a<��a<�a<��a<;�a<��a<.�a<��a<D�a<͍a<\�a<��a<��a<&�a<��a<�a<�a<��a<o�a<�a<��a<W�a<�a<��a<V�a<��a<��a<c�a<�a<�a<��a<U�a<2�a<��a<ƅa<��a<x�a<Q�a<D�a<�a<�a<لa<��a<��a<��a<��a<p�a<V�a<B�a<Q�a<F�a<P�a<T�a<p�a<q�a<��a<��a<�a<�  �  ��a<�a<\�a<y�a<��a<݅a<�a<B�a<l�a<��a<̆a<�a<h�a<��a<�a<*�a<��a<҈a<1�a<��a<��a<Z�a<��a<*�a<{�a<��a<J�a<��a<�a<i�a<��a<S�a<Ύa<=�a<��a<0�a<��a<>�a<��a<T�a<��a<L�a<ݓa<Z�a<
�a<s�a<�a<��a<�a<��a<�a<��a<�a<��a< �a<z�a<��a<p�a<��a<M�a<�a<O�a<Нa<%�a<��a<�a<e�a<�a<�a<|�a<Рa<�a<��a<��a<�a<5�a<��a<��a<�a<j�a<��a<��a<�a<l�a<��a<֤a<#�a<<�a<��a<��a<��a<�a<��a<�a<!�a<b�a<`�a<��a<��a<��a<̦a<ʦa< �a<�a<$�a<	�a<5�a<:�a<6�a<N�a<$�a<2�a<�a<�a<�a<��a<�a<Ӧa<�a<��a<Ӧa<��a<��a<��a<��a<��a<i�a<y�a<U�a<:�a<%�a<�a<�a<��a<��a<R�a<7�a<�a<Ԥa<��a<{�a<o�a<#�a<��a<գa<��a<u�a<!�a<�a<¢a<��a<C�a<�a<��a<Q�a<(�a<Ša<��a<,�a<ßa<��a<'�a<��a<��a<^�a<�a<��a<K�a<�a<��a<+�a<ޛa<a�a<�a<��a<�a<��a<�a<��a<B�a<ɗa<U�a<ږa<r�a<֕a<��a<��a<��a< �a<��a<1�a<��a<:�a<��a<!�a<��a<�a<��a<�a<��a<(�a<��a<E�a<�a<��a<�a<ҋa<P�a<�a<��a<R�a<�a<��a<g�a<�a<��a<^�a<�a<��a<[�a<;�a<܆a<��a<b�a<=�a<�a<��a<��a<��a<l�a< �a<!�a<��a<لa<Ԅa<��a<��a<g�a<c�a<c�a<>�a<P�a<+�a<T�a<:�a<m�a<p�a<��a<��a<��a<�  �  ��a<"�a<:�a<s�a<��a<؅a<�a<:�a<a�a<��a<�a<�a<A�a<��a<�a<2�a<�a<�a<F�a<��a<��a<V�a<��a<�a<|�a<�a</�a<��a<�a<u�a<�a<C�a<��a<C�a<��a<(�a<��a<1�a<��a<5�a<��a<P�a<�a<_�a<�a<u�a<��a<��a<	�a<��a<��a<��a<�a<��a<�a<|�a<��a<b�a<�a<q�a<�a<E�a<˝a<4�a<��a<�a<j�a<˟a<�a<��a<ˠa<�a<d�a<��a<��a<A�a<��a<Ӣa<�a<W�a<��a<�a<�a<b�a<��a<��a<�a<>�a<l�a<��a<��a<�a<��a<'�a<A�a<L�a<`�a<��a<��a<��a<˦a<�a<�a<��a<�a<$�a<6�a<0�a<3�a<*�a<2�a<4�a<%�a<�a<�a<�a<��a<�a<ئa<ʦa<̦a<��a<��a<��a<��a<��a<}�a<X�a<N�a<7�a<!�a<��a<ܥa<��a<��a<w�a<>�a<�a<�a<��a<��a<S�a<;�a<�a<ˣa<��a<r�a<<�a<�a<¢a<��a<)�a< �a<��a<]�a<�a<��a<q�a<1�a<ןa<��a<1�a<�a<��a<@�a<�a<��a<R�a<�a<��a<-�a<˛a<m�a<��a<��a<�a<��a<<�a<��a<-�a<̗a<S�a<̖a<d�a<��a<~�a<�a<��a<�a<��a<�a<��a< �a<��a<+�a<��a<�a<��a<�a<��a<4�a<��a<V�a<�a<}�a<�a<��a<V�a<�a<��a<=�a< �a<��a<R�a<�a<��a<[�a< �a<Ǉa<|�a<%�a<܆a<��a<n�a<�a<�a<�a<��a<s�a<`�a<;�a<!�a<��a<ׄa<��a<��a<��a<u�a<R�a<H�a<8�a<E�a<9�a<A�a<I�a<f�a<l�a<��a<��a<Єa<�  �  �a<2�a<;�a<��a<��a<υa<�a<4�a<~�a<��a<�a<�a<\�a<Ƈa<�a<\�a<��a<�a<@�a<��a<�a<S�a<ˊa<�a<x�a<�a<D�a<��a<�a<��a<ɍa<R�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<L�a<ԓa<z�a<ܔa<��a<�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<��a<��a<�a<q�a<�a<]�a<Нa<@�a<��a<��a<|�a<��a<2�a<w�a<Ġa<�a<C�a<��a<�a<0�a<n�a<��a<��a<J�a<��a<��a<4�a<T�a<��a<ڤa<	�a<?�a<d�a<��a<��a<�a<��a<$�a<C�a<H�a<��a<��a<��a<��a<Ʀa<�a<�a<�a<�a<:�a<,�a<$�a<E�a<$�a<J�a<�a<-�a<�a<�a<��a<ئa<զa<��a<��a<��a<��a<��a<��a<��a<x�a<��a<X�a<[�a<*�a<�a<�a<֥a<ƥa<��a<k�a<:�a<�a<�a<��a<��a<U�a<;�a<
�a<ѣa<��a<n�a<N�a<��a<��a<��a<=�a<�a<��a<u�a<��a<Ša<i�a<�a<ğa<f�a<#�a<Ҟa<��a<$�a<�a<��a<B�a<�a<}�a<D�a<��a<p�a<�a<��a<&�a<��a<:�a<��a<T�a<ؗa<[�a<��a<a�a<��a<|�a<
�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<"�a<}�a<#�a<��a<"�a<��a<@�a<Ќa<p�a<"�a<��a<p�a<��a<��a<V�a<��a<��a<J�a<�a<��a<h�a<	�a<Ňa<}�a<!�a<
�a<��a<��a<<�a< �a<�a<��a<��a<[�a<Q�a<�a<�a<�a<��a<��a<y�a<|�a<R�a<7�a<=�a<%�a<.�a<$�a<=�a<A�a<n�a<�a<��a<܄a<�  �  �a<�a<F�a<��a<��a<�a<��a<=�a<s�a<��a<܆a<'�a<q�a<��a<هa<=�a<��a<�a<?�a<��a<��a<[�a<��a</�a<��a<�a<D�a<��a<	�a<z�a<Ӎa<N�a<��a<'�a<��a<+�a<��a<�a<��a<,�a<��a<G�a<͓a<Y�a<�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<
�a<u�a<�a<{�a<��a<f�a<�a<\�a<Νa<2�a<��a<�a<z�a<˟a<�a<o�a<Ƞa<�a<Y�a<��a<�a<6�a<��a<ˢa<�a<F�a<��a<Σa<%�a<Z�a<��a<Ԥa<�a<E�a<�a<��a<��a<�a<
�a<&�a<9�a<^�a<p�a<t�a<��a<Ŧa<Ӧa<�a<�a<�a<�a<�a<7�a<6�a<H�a<3�a<%�a<�a<�a<�a< �a<�a<�a<ަa<ڦa<ʦa<��a<��a<��a<��a<��a<|�a<o�a<c�a<b�a<9�a<*�a<�a<ߥa<��a<��a<b�a<E�a<#�a<�a<��a<��a<l�a<8�a<	�a<�a<��a<w�a<4�a<�a<ɢa<��a<=�a<�a<��a<b�a<�a<��a<b�a<�a<՟a<��a<,�a<՞a<��a<7�a<�a<��a<;�a<�a<��a<D�a<ӛa<m�a<�a<��a<�a<��a</�a<Řa<M�a<ŗa<K�a<�a<u�a<�a<��a<
�a<��a<�a<��a<#�a<��a<!�a<��a<�a<��a<�a<��a<#�a<��a<)�a<a<O�a<ڌa<l�a<�a<��a<a�a<��a<��a<P�a<�a<��a<e�a<��a<��a<^�a<�a<Ǉa<s�a<7�a<�a<��a<k�a<I�a<�a<ׅa<��a<��a<e�a<2�a<"�a<��a<�a<��a<��a<z�a<i�a<X�a<D�a<9�a</�a<7�a<C�a<I�a<M�a<e�a<��a<��a<Ȅa<�  �  �a<�a<M�a<f�a<��a<�a<��a<V�a<T�a<��a<�a<'�a<j�a<��a<(�a<B�a<��a<�a<J�a<��a<�a<t�a<��a<-�a<e�a<ۋa<D�a<��a<�a<c�a<�a<G�a<��a<-�a<��a<�a<��a<�a<��a<;�a<��a<G�a<�a<X�a<��a<d�a<��a<��a<�a<��a<��a<��a<�a<��a<��a<��a<�a<r�a<
�a<l�a<��a<N�a<ݝa<B�a<��a<�a<T�a<՟a<�a<��a<Ǡa<�a<l�a<��a<�a<&�a<n�a<��a<�a<@�a<��a<�a<�a<\�a<��a<Фa<�a<%�a<{�a<��a<֥a<ߥa<�a</�a<9�a<p�a<p�a<��a<��a<��a<٦a<�a<	�a<�a<6�a<�a<A�a<%�a<$�a<A�a<%�a<@�a<
�a<�a<�a<�a<�a<¦a<��a<��a<��a<��a<��a<��a<{�a<��a<q�a<k�a<B�a<&�a<2�a<�a<��a<��a<��a<g�a<E�a<�a<�a<�a<��a<t�a<6�a<�a<�a<��a<��a<&�a<�a<��a<}�a<=�a<��a<��a<K�a<�a<��a<\�a<�a<��a<i�a<�a<Оa<��a<E�a<ݝa<��a<Y�a<�a<��a<�a<Ûa<m�a<��a<��a<�a<��a<8�a<јa<B�a<�a<{�a<ܖa<��a<��a<��a<��a<��a<�a<��a<�a<��a<*�a<��a<-�a<��a<�a<��a<�a<��a<�a<��a<2�a<ڌa<f�a<�a<Ëa<C�a<��a<��a<L�a<��a<��a<b�a<�a<ƈa<Z�a<�a<Їa<s�a<I�a<�a<ކa<��a<A�a<�a<ۅa<��a<h�a<~�a<3�a<-�a<�a<Ȅa<Ȅa<��a<��a<Z�a<S�a<L�a<,�a<2�a<�a<$�a<,�a<T�a<X�a<��a<��a<��a<�  �  �a<�a<F�a<��a<��a<�a<��a<=�a<s�a<��a<܆a<'�a<q�a<��a<هa<=�a<��a<�a<?�a<��a<��a<[�a<��a</�a<��a<�a<D�a<��a<	�a<z�a<Ӎa<N�a<��a<'�a<��a<+�a<��a<�a<��a<,�a<��a<G�a<͓a<Y�a<�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<
�a<u�a<�a<{�a<��a<f�a<�a<\�a<Νa<2�a<��a<�a<z�a<˟a<�a<o�a<Ƞa<�a<Y�a<��a<�a<6�a<��a<ˢa<�a<F�a<��a<Σa<%�a<Z�a<��a<Ԥa<�a<E�a<�a<��a<��a<�a<
�a<&�a<9�a<^�a<p�a<t�a<��a<Ŧa<Ӧa<�a<�a<�a<�a<�a<7�a<6�a<H�a<3�a<%�a<�a<�a<�a< �a<�a<�a<ަa<ڦa<ʦa<��a<��a<��a<��a<��a<|�a<o�a<c�a<b�a<9�a<*�a<�a<ߥa<��a<��a<b�a<E�a<#�a<�a<��a<��a<l�a<8�a<	�a<�a<��a<w�a<4�a<�a<ɢa<��a<=�a<�a<��a<b�a<�a<��a<b�a<�a<՟a<��a<,�a<՞a<��a<7�a<�a<��a<;�a<�a<��a<D�a<ӛa<m�a<�a<��a<�a<��a</�a<Řa<M�a<ŗa<K�a<�a<u�a<�a<��a<
�a<��a<�a<��a<#�a<��a<!�a<��a<�a<��a<�a<��a<#�a<��a<)�a<a<O�a<ڌa<l�a<�a<��a<a�a<��a<��a<P�a<�a<��a<e�a<��a<��a<^�a<�a<Ǉa<s�a<7�a<�a<��a<k�a<I�a<�a<ׅa<��a<��a<e�a<2�a<"�a<��a<�a<��a<��a<z�a<i�a<X�a<D�a<9�a</�a<7�a<C�a<I�a<M�a<e�a<��a<��a<Ȅa<�  �  �a<2�a<;�a<��a<��a<υa<�a<4�a<~�a<��a<�a<�a<\�a<Ƈa<�a<\�a<��a<�a<@�a<��a<�a<S�a<ˊa<�a<x�a<�a<D�a<��a<�a<��a<ɍa<R�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<L�a<ԓa<z�a<ܔa<��a<�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<��a<��a<�a<q�a<�a<]�a<Нa<@�a<��a<��a<|�a<��a<2�a<w�a<Ġa<�a<C�a<��a<�a<0�a<n�a<��a<��a<J�a<��a<��a<4�a<T�a<��a<ڤa<	�a<?�a<d�a<��a<��a<�a<��a<$�a<C�a<H�a<��a<��a<��a<��a<Ʀa<�a<�a<�a<�a<:�a<,�a<$�a<E�a<$�a<J�a<�a<-�a<�a<�a<��a<ئa<զa<��a<��a<��a<��a<��a<��a<��a<x�a<��a<X�a<[�a<*�a<�a<�a<֥a<ƥa<��a<k�a<:�a<�a<�a<��a<��a<U�a<;�a<
�a<ѣa<��a<n�a<N�a<��a<��a<��a<=�a<�a<��a<u�a<��a<Ša<i�a<�a<ğa<f�a<#�a<Ҟa<��a<$�a<�a<��a<B�a<�a<}�a<D�a<��a<p�a<�a<��a<&�a<��a<:�a<��a<T�a<ؗa<[�a<��a<a�a<��a<|�a<
�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<"�a<}�a<#�a<��a<"�a<��a<@�a<Ќa<p�a<"�a<��a<p�a<��a<��a<V�a<��a<��a<J�a<�a<��a<h�a<	�a<Ňa<}�a<!�a<
�a<��a<��a<<�a< �a<�a<��a<��a<[�a<Q�a<�a<�a<�a<��a<��a<y�a<|�a<R�a<7�a<=�a<%�a<.�a<$�a<=�a<A�a<n�a<�a<��a<܄a<�  �  ��a<"�a<:�a<s�a<��a<؅a<�a<:�a<a�a<��a<�a<�a<A�a<��a<�a<2�a<�a<�a<F�a<��a<��a<V�a<��a<�a<|�a<�a</�a<��a<�a<u�a<�a<C�a<��a<C�a<��a<(�a<��a<1�a<��a<5�a<��a<P�a<�a<_�a<�a<u�a<��a<��a<	�a<��a<��a<��a<�a<��a<�a<|�a<��a<b�a<�a<q�a<�a<E�a<˝a<4�a<��a<�a<j�a<˟a<�a<��a<ˠa<�a<d�a<��a<��a<A�a<��a<Ӣa<�a<W�a<��a<�a<�a<b�a<��a<��a<�a<>�a<l�a<��a<��a<�a<��a<'�a<A�a<L�a<`�a<��a<��a<��a<˦a<�a<�a<��a<�a<$�a<6�a<0�a<3�a<*�a<2�a<4�a<%�a<�a<�a<�a<��a<�a<ئa<ʦa<̦a<��a<��a<��a<��a<��a<}�a<X�a<N�a<7�a<!�a<��a<ܥa<��a<��a<w�a<>�a<�a<�a<��a<��a<S�a<;�a<�a<ˣa<��a<r�a<<�a<�a<¢a<��a<)�a< �a<��a<]�a<�a<��a<q�a<1�a<ןa<��a<1�a<�a<��a<@�a<�a<��a<R�a<�a<��a<-�a<˛a<m�a<��a<��a<�a<��a<<�a<��a<-�a<̗a<S�a<̖a<d�a<��a<~�a<�a<��a<�a<��a<�a<��a< �a<��a<+�a<��a<�a<��a<�a<��a<4�a<��a<V�a<�a<}�a<�a<��a<V�a<�a<��a<=�a< �a<��a<R�a<�a<��a<[�a< �a<Ǉa<|�a<%�a<܆a<��a<n�a<�a<�a<�a<��a<s�a<`�a<;�a<!�a<��a<ׄa<��a<��a<��a<u�a<R�a<H�a<8�a<E�a<9�a<A�a<I�a<f�a<l�a<��a<��a<Єa<�  �  ��a<�a<\�a<y�a<��a<݅a<�a<B�a<l�a<��a<̆a<�a<h�a<��a<�a<*�a<��a<҈a<1�a<��a<��a<Z�a<��a<*�a<{�a<��a<J�a<��a<�a<i�a<��a<S�a<Ύa<=�a<��a<0�a<��a<>�a<��a<T�a<��a<L�a<ݓa<Z�a<
�a<s�a<�a<��a<�a<��a<�a<��a<�a<��a< �a<z�a<��a<p�a<��a<M�a<�a<O�a<Нa<%�a<��a<�a<e�a<�a<�a<|�a<Рa<�a<��a<��a<�a<5�a<��a<��a<�a<j�a<��a<��a<�a<l�a<��a<֤a<#�a<<�a<��a<��a<��a<�a<��a<�a<!�a<b�a<`�a<��a<��a<��a<̦a<ʦa< �a<�a<$�a<	�a<5�a<:�a<6�a<N�a<$�a<2�a<�a<�a<�a<��a<�a<Ӧa<�a<��a<Ӧa<��a<��a<��a<��a<��a<i�a<y�a<U�a<:�a<%�a<�a<�a<��a<��a<R�a<7�a<�a<Ԥa<��a<{�a<o�a<#�a<��a<գa<��a<u�a<!�a<�a<¢a<��a<C�a<�a<��a<Q�a<(�a<Ša<��a<,�a<ßa<��a<'�a<��a<��a<^�a<�a<��a<K�a<�a<��a<+�a<ޛa<a�a<�a<��a<�a<��a<�a<��a<B�a<ɗa<U�a<ږa<r�a<֕a<��a<��a<��a< �a<��a<1�a<��a<:�a<��a<!�a<��a<�a<��a<�a<��a<(�a<��a<E�a<�a<��a<�a<ҋa<P�a<�a<��a<R�a<�a<��a<g�a<�a<��a<^�a<�a<��a<[�a<;�a<܆a<��a<b�a<=�a<�a<��a<��a<��a<l�a< �a<!�a<��a<لa<Ԅa<��a<��a<g�a<c�a<c�a<>�a<P�a<+�a<T�a<:�a<m�a<p�a<��a<��a<��a<�  �  ��a<*�a<M�a<r�a<��a<օa<�a<*�a<e�a<��a<φa<�a<U�a<��a<ׇa</�a<x�a<шa<0�a<��a<�a<M�a<��a<�a<u�a<ۋa<[�a<��a<�a<��a<�a<^�a<ˎa<G�a<��a<7�a<��a<9�a<��a<;�a<ޒa<^�a<ۓa<�a<�a<z�a<��a<��a<	�a<��a<��a<��a<��a<o�a<��a<\�a<ٚa<m�a<ڛa<Z�a<՜a<F�a<��a<6�a<��a<
�a<l�a<��a<>�a<y�a<٠a<7�a<j�a<��a<�a<Q�a<��a<٢a<&�a<e�a<��a<�a<C�a<i�a<��a<�a<�a<9�a<q�a<��a<��a<ۥa<�a<�a<(�a<?�a<e�a<j�a<��a<��a<��a<Ϧa<�a<��a<
�a<-�a</�a<)�a<6�a<5�a<C�a<.�a<8�a<)�a<�a<��a<�a<�a<�a<զa<֦a<��a<��a<��a<��a<��a<��a<k�a<M�a</�a<�a<�a<̥a<��a<}�a<U�a<*�a<�a<Ϥa<��a<��a<L�a<"�a<��a<��a<��a<h�a<@�a<�a<��a<}�a<T�a<��a<��a<��a<�a<Рa<}�a<6�a<ݟa<��a<D�a<�a<��a<F�a<�a<��a<I�a<�a<��a<2�a<ƛa<g�a<��a<��a<�a<��a<#�a<��a<=�a<��a<5�a<זa<S�a<�a<p�a<��a<��a<�a<��a<�a<��a<�a<��a<�a<��a<;�a<��a<.�a<��a<D�a<͍a<\�a<��a<��a<&�a<��a<�a<�a<��a<o�a<�a<��a<W�a<�a<��a<V�a<��a<��a<c�a<�a<�a<��a<U�a<2�a<��a<ƅa<��a<x�a<Q�a<D�a<�a<�a<لa<��a<��a<��a<��a<p�a<V�a<B�a<Q�a<F�a<P�a<T�a<p�a<q�a<��a<��a<�a<�  �  �a<:�a<>�a<��a<��a<��a<�a<�a<n�a<�a<цa<��a<C�a<��a<��a<,�a<g�a<ψa<"�a<�a<�a<0�a<a<��a<��a<ߋa<J�a<��a<�a<��a<�a<r�a<ˎa<R�a<Ǐa</�a<͐a</�a<Ցa<=�a<ܒa<^�a<ϓa<~�a<ٔa<��a<�a<��a<��a<j�a<�a<`�a<��a<X�a<�a<[�a<њa<e�a<��a<_�a<��a<Q�a<��a<!�a<��a<�a<��a<��a<:�a<v�a<Ԡa<8�a<h�a<աa<��a<e�a<��a<�a<7�a<^�a<��a<ߣa<D�a<Y�a<��a<�a<�a<]�a<N�a<��a<��a<ԥa<�a<��a</�a<)�a<^�a<X�a<��a<��a<��a<Ԧa<̦a<�a<�a<#�a<!�a<3�a<Q�a<&�a<O�a<�a<?�a< �a<�a<�a<��a<�a<ݦa<�a<զa<ɦa<Ȧa<��a<��a<{�a<��a<\�a<f�a<D�a<�a<�a<��a<��a<i�a<W�a<�a<��a<Фa<��a<~�a<;�a< �a<�a<��a<��a<K�a<F�a<�a<ޢa<��a<D�a<�a<��a<��a<�a<�a<~�a<A�a<�a<��a<Y�a<�a<��a<H�a<�a<��a<=�a<�a<{�a<O�a<��a<j�a<�a<j�a<�a<}�a<'�a<��a<5�a<��a<.�a<ϖa<9�a<�a<S�a<��a<r�a<��a<��a< �a<��a<
�a<��a<�a<��a<=�a<��a<H�a<��a<W�a<ʍa<f�a<	�a<��a<>�a<��a<��a<��a<��a<d�a<�a<Ɖa<5�a<	�a<��a<O�a<��a<��a<i�a<�a<ۆa<}�a<X�a< �a<�a<˅a<��a<��a<4�a<9�a<�a<��a<�a<��a<��a<z�a<��a<g�a<b�a<Z�a<K�a<_�a<G�a<k�a<o�a<��a<��a<��a<�a<�  �  ��a<:�a<U�a<q�a<��a<Ѕa<��a<$�a<f�a<��a<��a<�a<@�a<y�a<ʇa<�a<n�a<��a<�a<��a<�a<?�a<��a<�a<|�a<܋a<T�a<ǌa<"�a<��a< �a<m�a<��a<b�a<ŏa<>�a<Ԑa<F�a<Αa<V�a<Ԓa<g�a<�a<{�a<��a<t�a<�a<��a<�a<w�a<�a<g�a<�a<b�a<ߙa<U�a<њa<R�a<͛a<F�a<��a<P�a<��a<�a<��a<��a<k�a<՟a<8�a<��a<�a<-�a<��a<ϡa<�a<l�a<��a<�a<@�a<u�a<��a< �a<8�a<u�a<��a<�a<�a<?�a<\�a<��a<��a<ӥa<��a<��a<�a<2�a<I�a<a�a<s�a<��a<��a<æa<֦a<�a<�a<�a<2�a<*�a<1�a<@�a<K�a<:�a<>�a<'�a<(�a<�a<�a<�a<��a<�a<�a<Ԧa<Ȧa<��a<��a<��a<��a<s�a<L�a<0�a<�a<��a<ƥa<��a<v�a<G�a<�a<�a<��a<��a<d�a<B�a<�a<�a<ƣa<��a<[�a<=�a<��a<¢a<~�a<M�a<�a<��a<x�a</�a<�a<��a<P�a<�a<��a<`�a< �a<��a<`�a<�a<��a<Y�a<�a<��a<,�a<��a<r�a<��a<w�a<�a<��a<�a<��a<"�a<��a<.�a<��a<F�a<ϕa<V�a<��a<{�a<��a<��a<
�a<��a<*�a<��a<3�a<��a<1�a<��a<B�a<Ŏa<_�a<֍a<d�a<�a<��a<;�a<ۋa<t�a<�a<Êa<c�a<��a<��a<B�a<�a<��a<N�a< �a<��a<K�a<�a<ņa<��a<E�a<�a<߅a<��a<��a<��a<K�a<-�a<�a<�a<Ԅa<Ǆa<��a<��a<��a<n�a<k�a<_�a<[�a<`�a<_�a<k�a<��a<��a<��a<��a<�a<�  �  �a<�a<_�a<z�a<��a<مa<�a<'�a<<�a<��a<��a<��a<<�a<^�a<ˇa<��a<p�a<��a<(�a<s�a<ωa<C�a<��a<*�a<x�a<�a<Y�a<��a<9�a<��a<�a<d�a<�a<k�a<֏a<[�a<Аa<i�a<đa<b�a<��a<o�a<�a<c�a<�a<u�a<�a<s�a<�a<v�a<ۗa<y�a<Ԙa<f�a<əa<?�a<��a<9�a<қa<7�a<Ҝa<(�a<��a<"�a<��a<�a<f�a<�a<(�a<��a<�a<6�a<��a<¡a<5�a<m�a<��a<��a<F�a<��a<��a<�a<@�a<��a<��a<�a<#�a<8�a<~�a<z�a<��a<��a<֥a<�a<�a<6�a<.�a<]�a<X�a<��a<��a<��a<�a<զa<�a<	�a<)�a<:�a<9�a<O�a<(�a<I�a<D�a<<�a<(�a<�a</�a<�a<	�a<�a<��a<ߦa<Ʀa<ͦa<��a<��a<o�a<|�a<U�a<:�a<!�a<ݥa<ɥa<��a<y�a<E�a<�a<�a<��a<��a<I�a<C�a< �a<�a<��a<~�a<_�a<�a<�a<��a<��a<S�a<�a<֡a<��a<G�a<נa<��a<Y�a<��a<��a<\�a<"�a<��a<l�a<�a<��a<Z�a<�a<��a<-�a<ܛa<S�a<�a<w�a<�a<��a<��a<��a<�a<��a<�a<��a<K�a<��a<l�a<֔a<u�a<��a<��a<.�a<��a<=�a<��a<(�a<a<;�a<Ϗa<6�a<�a<`�a<�a<�a<�a<��a<,�a<�a<|�a<,�a<��a<a�a<�a<��a<e�a<�a<��a<8�a<�a<��a<@�a<�a<��a<��a<*�a<�a<��a<��a<��a<R�a<N�a< �a<�a<��a<܄a<քa<��a<��a<��a<��a<l�a<e�a<|�a<]�a<r�a<l�a<��a<��a<��a<ׄa<�a<�  �  �a<.�a<W�a<z�a<��a<��a<��a<'�a<M�a<z�a<��a<�a<8�a<o�a<��a<�a<d�a<��a<�a<e�a<ډa<E�a<��a<�a<w�a<�a<Z�a<��a<-�a<��a<�a<��a<�a<I�a<��a<\�a<ːa<U�a<�a<l�a<ܒa<n�a<�a<y�a<��a<z�a<��a<b�a<��a<n�a<ޗa<`�a<ʘa<R�a<ՙa<N�a<ƚa<E�a<��a<+�a<��a<%�a<��a<.�a<��a<�a<k�a<ϟa<:�a<��a<�a<0�a<��a<�a<%�a<a�a<��a< �a<,�a<��a<٣a<�a<3�a<�a<��a<�a<�a<9�a<_�a<��a<��a<ĥa<˥a<�a<��a<+�a<7�a<P�a<k�a<��a<��a<��a<Φa<�a< �a<�a<�a</�a<9�a<B�a<D�a<F�a<:�a<1�a<A�a<2�a<�a<�a<�a<��a<٦a<�a<�a<��a<��a<��a<��a<u�a<U�a<2�a<��a<�a<ɥa<��a<d�a<0�a<�a<�a<��a<��a<V�a<8�a<��a<֣a<��a<��a<a�a<'�a<�a<��a<��a<T�a<�a<ʡa<r�a<5�a<�a<��a<7�a<�a<��a<W�a<�a<ʞa<v�a<�a<��a<]�a<�a<��a<2�a<ɛa<B�a<�a<n�a<�a<}�a<��a<��a<�a<��a<"�a<��a<7�a<��a<P�a<Ӕa<m�a<	�a<{�a<�a<��a<$�a<��a<2�a<��a<4�a<Ϗa<Y�a<֎a<T�a<�a<��a<��a<��a<W�a<�a<p�a<"�a<a<j�a<�a<��a<E�a<�a<��a<?�a<ևa<��a<9�a<�a<��a<u�a<=�a<�a<Ӆa<��a<��a<_�a<G�a</�a<��a<�a<݄a<Ʉa<��a<��a<��a<x�a<��a<x�a<\�a<h�a<v�a<{�a<s�a<��a<Ȅa<Ʉa<�a<�  �  �a<E�a<N�a<m�a<��a<��a<�a<�a<]�a<h�a<��a<�a<�a<a�a<��a<��a<E�a<��a<��a<i�a<߉a<1�a<��a<��a<��a<׋a<S�a<֌a<+�a<��a<�a<��a<�a<o�a<��a<^�a<��a<O�a<�a<h�a<�a<x�a<�a<��a<�a<}�a<�a<{�a<��a<`�a<��a<?�a<��a<C�a<��a<8�a<��a</�a<��a<=�a<��a<9�a<��a<"�a<��a<��a<y�a<ßa<F�a<��a<�a<B�a<��a<�a<!�a<��a<��a<�a<S�a<��a<֣a<�a<S�a<�a<ɤa<�a<�a<P�a<N�a<��a<��a<åa<إa<֥a<�a<�a<)�a<5�a<Z�a<g�a<��a<��a<��a<��a<�a<�a<�a<5�a<2�a<:�a<V�a<A�a<R�a<5�a<9�a<2�a<�a<7�a<�a<"�a<�a<�a<ܦa<��a<Ȧa<��a<��a<l�a<H�a<<�a<�a<��a<��a<��a<Q�a<0�a<	�a<äa<��a<i�a<J�a<�a<��a<��a<��a<��a<M�a<B�a<�a<Ӣa<y�a<M�a<#�a<ǡa<��a<6�a<��a<��a<]�a< �a<��a<��a<	�a<˞a<s�a<�a<ȝa<_�a<�a<��a<5�a<��a<[�a<�a<a�a<�a<\�a<	�a<y�a<��a<��a<�a<��a<%�a<ƕa<.�a<�a<d�a<��a<��a<	�a<��a<�a<��a<;�a<Őa<F�a<̏a<Z�a<Ҏa<��a<��a<��a<&�a<��a<T�a<�a<��a<!�a<֊a<j�a<��a<��a<5�a<�a<��a<>�a<�a<v�a<A�a<�a<��a<Z�a<,�a<�a<υa<��a<k�a<u�a<5�a<6�a<	�a<��a<Մa<��a<ńa<��a<��a<|�a<|�a<w�a<c�a<��a<p�a<��a<��a<��a<��a<ʄa< �a<�  �  �a<&�a<d�a<z�a<��a<ƅa<�a<�a<I�a<r�a<��a<�a<�a<o�a<��a<�a<M�a<��a<�a<m�a<Ήa<1�a<��a<�a<��a<�a<\�a<��a<4�a<��a<�a<}�a<��a<w�a<ۏa<M�a<ݐa<d�a<ݑa<l�a<�a<p�a<�a<u�a<�a<��a< �a<r�a<�a<f�a<�a<P�a<ۘa<A�a<��a<G�a<ƚa<5�a<��a<<�a<��a<4�a<��a<�a<��a<�a<x�a<۟a<7�a<��a<�a<D�a<��a<ܡa<4�a<y�a<��a<��a<Q�a<��a<ɣa<�a<K�a<��a<��a<�a<�a<S�a<`�a<y�a<��a<��a<إa<�a<�a<�a<3�a<V�a<j�a<t�a<��a<��a<��a<�a<�a<�a<�a<=�a<>�a<U�a<;�a<J�a<E�a<J�a<6�a<3�a</�a<�a<��a<��a<�a<�a<Ԧa<צa<��a<��a<��a<��a<V�a<D�a<�a<ߥa<��a<��a<[�a<3�a<��a<Ϥa<��a<��a<S�a< �a<��a<ѣa<��a<}�a<M�a<�a<��a<բa<��a<V�a<�a<Сa<��a<M�a<�a<��a<e�a<�a<��a<i�a<�a<��a<w�a<�a<��a<^�a<��a<��a<:�a<͛a<Q�a<ݚa<g�a<��a<l�a<�a<w�a<�a<��a<"�a<��a<$�a<ŕa<D�a<�a<j�a<�a<��a<�a<��a<0�a<��a<3�a<��a<I�a<֏a<O�a<�a<l�a<�a<}�a<$�a<��a<G�a<��a<��a<(�a<��a<j�a<	�a<��a<F�a<�a<��a<5�a<�a<��a<?�a<�a<��a<z�a<<�a<��a<ǅa<��a<v�a<b�a<:�a<�a<
�a<�a<�a<܄a<��a<��a<��a<��a<z�a<y�a<{�a<q�a<`�a<�a<��a<��a<��a<�a<�a<�  �  �a<�a<9�a<:�a<R�a<��a<��a<a<لa<+�a<R�a<��a<υa<�a<H�a<��a<�a<]�a<��a<&�a<k�a<��a<d�a<�a</�a<ˊa<C�a<��a<>�a<f�a<�a<_�a<ҍa<?�a<ʎa<j�a<��a<F�a<��a<t�a<ۑa<e�a<
�a<c�a<�a<W�a<��a<j�a<�a<B�a<��a<M�a<��a<K�a<��a<�a<��a<'�a<��a<�a<��a<�a<��a<+�a<��a<"�a<o�a<�a<S�a<ϟa<"�a<\�a<۠a<�a<L�a<��a<�a<0�a<`�a<��a<�a<S�a<X�a<ˣa<أa<�a<K�a<9�a<��a<��a<��a<��a<դa<��a<��a<$�a<�a</�a<<�a<z�a<��a<��a<ͥa<ɥa<�a<�a<,�a<=�a<D�a<{�a<P�a<��a<K�a<a�a<_�a<0�a<6�a<"�a<F�a<�a<�a<�a<��a<��a<��a<��a<��a<��a<f�a<5�a<�a<�a<��a<o�a<a�a<%�a<�a<̣a<~�a<^�a<0�a<(�a<��a<Тa<��a<`�a<V�a<+�a<�a<��a<��a<|�a< �a<�a<��a<x�a<�a<��a<d�a<%�a<��a<q�a</�a<ǝa<��a<2�a<ڜa<��a<�a<Лa<+�a<ښa<^�a<�a<Q�a<٘a<q�a<ܗa<��a<��a<a�a<�a<��a<&�a<��a<5�a<��a<4�a<�a<t�a<�a<v�a<;�a<��a<A�a<��a<(�a<ڎa<%�a<��a<<�a<��a<p�a<�a<��a<�a<�a<L�a<$�a<��a<K�a<�a<U�a<�a<��a<M�a<͆a<��a<E�a<�a<��a<G�a<�a<��a<��a<��a<E�a<1�a<�a<�a<ڃa<ăa<��a<��a<��a<l�a<��a<F�a<T�a<N�a<!�a<.�a<'�a<[�a<@�a<J�a<T�a<��a<��a<��a<�  �  Ӄa<�a< �a<8�a<r�a<}�a<��a<݄a<�a<#�a<K�a<��a<��a<�a<_�a<��a<�a<Q�a<��a<'�a<��a<�a<j�a<؉a<W�a<��a<+�a<��a<�a<z�a<�a<[�a<�a<V�a<��a<;�a<a<Y�a<֐a<L�a<ёa<[�a<ےa<d�a<��a<p�a<��a<d�a<�a<m�a<�a<:�a<��a<&�a<��a<.�a<��a<)�a<��a<%�a<��a<?�a<��a<3�a<��a<%�a<��a<��a<O�a<��a<
�a<Y�a<��a<�a<`�a<��a<ءa<�a<r�a<¢a<�a<-�a<g�a<��a<��a<�a<.�a<a�a<{�a<��a<��a<ؤa<�a<�a<��a<�a<0�a<E�a<]�a<j�a<��a<��a<��a<��a<�a<"�a<&�a<S�a<J�a<`�a<O�a<Y�a<X�a<Y�a<L�a<V�a<K�a<+�a<�a<�a<�a<�a<�a<�a<ɥa<��a<��a<��a<d�a<V�a<�a<��a<ͤa<��a<Y�a<�a<�a<��a<��a<u�a<K�a<�a<�a<��a<��a<��a<h�a<1�a<�a<�a<��a<e�a<�a<�a<��a<W�a<�a<՟a<{�a<�a<ɞa<�a<B�a<�a<��a<(�a<Мa<l�a<�a<��a<D�a<�a<Y�a<�a<|�a<��a<^�a<�a<\�a<�a<v�a< �a<��a<�a<��a<$�a<ѓa<d�a<�a<s�a<�a<��a<�a<��a<�a<��a<%�a<��a<?�a<Ӎa<J�a<Ќa<Z�a< �a<��a<$�a<��a<[�a<��a<��a<3�a<ӈa<~�a<�a<��a<\�a<�a<��a<3�a<��a<��a<\�a<�a<݄a<��a<j�a<F�a<"�a<!�a<�a<�a<��a<ăa<��a<��a<j�a<b�a<S�a<L�a<<�a<H�a<C�a<0�a<,�a<=�a<_�a<x�a<|�a<��a<��a<�  �  ƃa<�a<�a<9�a<s�a<r�a<��a<��a<��a<�a<q�a<��a<˅a<�a<9�a<��a<��a<t�a<̇a<�a<��a<݈a<��a<ĉa<e�a<��a<8�a<��a< �a<��a<یa<a�a<ʍa<G�a<Ύa<C�a<Џa<-�a<ސa<>�a<�a<x�a<ߒa<��a<ߓa<}�a<�a<i�a<ܕa<@�a<Ֆa<=�a<�a<0�a<��a<'�a<��a<8�a<��a<S�a<��a<3�a<��a<�a<��a<�a<��a<��a<s�a<��a<"�a<z�a<��a<�a<7�a<��a<�a<+�a<f�a<��a<��a<�a<��a<��a<�a<�a< �a<r�a<h�a<��a<��a<��a<פa<��a<�a<�a<:�a<'�a<_�a<v�a<��a<̥a<��a<�a<�a<"�a<!�a<O�a<Q�a<O�a<z�a<M�a<x�a<Z�a<E�a<N�a<�a<?�a<!�a<$�a<�a<�a<�a<ߥa<�a<��a<��a<��a<e�a<W�a<	�a<��a<��a<��a<S�a<D�a<�a<ȣa<��a<N�a<S�a<�a<�a<ݢa<��a<��a<=�a<G�a<�a<�a<��a<r�a<:�a<ڠa<àa<F�a<�a<��a<l�a<)�a<Ҟa<��a<�a<�a<t�a<>�a<�a<p�a<6�a<��a<P�a<Қa<^�a<ޙa<O�a<�a<a�a<�a<f�a<��a<o�a<�a<��a<	�a<ǔa<*�a<ēa<@�a<Ԓa<{�a<��a<��a<�a<��a<'�a<��a<F�a<��a<L�a<��a<P�a<،a<l�a<��a<~�a</�a<��a<��a<��a<��a<I�a<Ĉa<��a<�a<ća<5�a<�a<��a<H�a<�a<��a<f�a<��a<߄a<��a<}�a<p�a<�a<�a<Ճa<�a<��a<��a<��a<��a<��a<V�a<s�a<M�a<5�a<@�a<�a<C�a<6�a<P�a<:�a<i�a<w�a<��a<Ӄa<�  �  уa<�a<�a<N�a<_�a<�a<Äa<҄a<�a<4�a<Y�a<��a<ׅa<�a<j�a<��a<�a<Z�a<ˇa<5�a<��a<��a<��a<ωa<P�a<Êa<(�a<��a<�a<p�a<ތa<l�a<Ía<F�a<��a<+�a<��a<0�a<ʐa<K�a<ʑa<P�a<ؒa<l�a<�a<��a<�a<y�a<��a<b�a<�a<Z�a<��a<9�a<��a<7�a<��a<;�a<��a<+�a<��a<G�a<��a<;�a<��a<�a<��a<�a<U�a<��a<��a<S�a<��a<�a<:�a<��a<ȡa<�a<g�a<��a<��a<�a<_�a<��a<ƣa<�a<7�a<]�a<o�a<��a<��a<ݤa<�a<��a<��a< �a<;�a<T�a<c�a<~�a<��a<��a<եa< �a<�a<3�a</�a<=�a<b�a<R�a<]�a<Y�a<K�a<I�a<S�a<<�a<'�a<*�a<
�a<�a<��a<��a<��a<Хa<��a<��a<��a<��a<z�a<C�a<�a<	�a<äa<��a<j�a<,�a<��a<ԣa<��a<��a<T�a<'�a<�a<ܢa<��a<��a<X�a<P�a<��a<١a<��a<b�a<�a<۠a<��a<H�a<�a<��a<k�a<�a<��a<|�a<�a<۝a<��a<!�a<Ɯa<i�a<�a<��a<T�a<˚a<m�a<��a<q�a<�a<~�a<�a<o�a< �a<�a<�a<��a<�a<��a<@�a<ٓa<b�a<�a<��a<��a<��a<�a<��a<�a<��a<�a<��a<=�a<��a<I�a<��a<W�a<��a<z�a<3�a<��a<S�a<�a<��a<6�a<܈a<y�a<	�a<̇a<Q�a<	�a<��a<N�a<�a<��a<f�a<(�a<�a<��a<u�a<M�a<:�a<)�a<��a<��a<ǃa<��a<��a<��a<x�a<b�a<F�a<<�a<C�a<.�a< �a</�a< �a<=�a<C�a<[�a<��a<��a<��a<�  �  �a<�a<�a<9�a<^�a<��a<��a<�a<��a<5�a<j�a<��a<��a<�a<��a<��a<�a<e�a<؇a<%�a<��a<�a<g�a<�a<I�a<��a<$�a<��a<�a<m�a<ތa<9�a<��a<>�a<��a<2�a<��a<B�a<��a<@�a<͑a<`�a<�a<Z�a<�a<f�a<��a<s�a<�a<m�a<ɖa<e�a<ȗa<^�a<��a<D�a<ʙa<)�a<Ϛa<2�a<Λa<'�a<��a<+�a<��a<$�a<��a<��a<G�a<��a<�a<V�a<��a<ؠa<B�a<~�a<ʡa<�a<Z�a<��a<Ǣa<�a<\�a<��a<Σa<��a<3�a<U�a<��a<��a<��a<դa<֤a<�a<�a<2�a<�a<n�a<^�a<��a<��a<��a<ݥa<�a<�a<�a<@�a<@�a<I�a<Y�a<O�a<o�a<O�a<K�a<7�a<�a<:�a<�a<�a<��a<	�a<ڥa<ԥa<եa<��a<ͥa<��a<��a<e�a<B�a<0�a<�a<Ҥa<��a<k�a<=�a<�a<ݣa<��a<��a<9�a<6�a<��a<�a<��a<��a<e�a</�a<�a<ҡa<��a<^�a<�a<��a<��a<H�a<�a<��a<c�a<�a<��a<f�a<+�a<��a<v�a<$�a<՜a<��a<�a<��a<9�a<ښa<h�a<�a<|�a<�a<��a<��a<��a<�a<��a<�a<��a<6�a<��a<O�a<��a<c�a<�a<z�a<�a<��a<�a<��a<*�a<��a<"�a<��a<�a<��a<1�a<��a<L�a<�a<u�a<��a<��a<P�a<
�a<��a</�a<؈a<r�a<#�a<��a<V�a<�a<��a<]�a<�a<��a<J�a<B�a<߄a<��a<��a<`�a<B�a<�a<�a<݃a<؃a<��a<��a<��a<k�a<x�a<J�a<>�a<&�a<�a<3�a<�a<*�a<(�a<P�a<A�a<a�a<��a<��a<�  �  ��a<��a<�a<4�a<`�a<��a<��a<�a<
�a<9�a<��a<��a<��a<*�a<�a<��a<.�a<o�a<�a<0�a<��a<�a<�a<ۉa<P�a<��a<.�a<��a<�a<a�a<ӌa<K�a<a<�a<��a<4�a<��a<"�a<��a<<�a<��a<H�a<Вa<k�a<�a<l�a<�a<~�a<�a<��a<ۖa<l�a<ٗa<S�a<Ҙa<S�a<Йa<J�a<̚a<@�a<כa<<�a<՜a<@�a<��a<�a<��a<�a<W�a<��a<��a<F�a<��a<�a<.�a<^�a<͡a<�a<8�a<��a<ۢa<�a<K�a<��a<ѣa<
�a<"�a<_�a<x�a<��a<ʤa<�a<�a<�a<�a<A�a<E�a<d�a<|�a<��a<��a<ѥa<�a<�a<�a<*�a<9�a<F�a<H�a<T�a<`�a<=�a<B�a<;�a<;�a<.�a<�a<��a<�a<�a<ܥa<�a<ݥa<ťa<��a<��a<��a<��a<`�a<D�a<"�a<�a<ݤa<��a<p�a<T�a<�a<��a<��a<��a<\�a<K�a<�a<��a<��a<��a<u�a<F�a<�a<١a<��a<h�a<%�a<��a<��a<=�a<��a<��a<>�a<��a<a<F�a<�a<Ɲa<r�a<�a<��a<a�a<�a<��a<?�a<ךa<r�a<��a<��a<��a<��a<�a<��a<�a<��a<"�a<��a<3�a<��a<Y�a<͓a<x�a<��a<��a<�a<��a<�a<��a<�a<��a<�a<��a<$�a<��a<�a<Ča<C�a<Ƌa<z�a<�a<��a<>�a<ۉa<��a<<�a<ƈa<|�a<�a<Ƈa<k�a<�a<��a<l�a< �a<ʅa<q�a<8�a<��a<фa<��a<u�a<F�a<�a<�a<�a<уa<��a<��a<��a<{�a<F�a<>�a<.�a<*�a<�a<�a<��a<+�a<�a<#�a<L�a<j�a<|�a<��a<�  �  ��a<�a<��a<M�a<t�a<x�a<Ʉa<܄a<.�a<B�a<��a<��a<�a<B�a<��a<܆a<1�a<��a<�a<D�a<��a<�a<��a<͉a<i�a<��a<�a<��a<�a<o�a<��a<9�a<��a< �a<��a<�a<��a<�a<��a<%�a<��a<M�a<ʒa<j�a<ӓa<��a<�a<v�a<��a<x�a<��a<i�a<�a<\�a<�a<Z�a<ٙa<e�a<Ԛa<U�a<Лa<U�a<Μa<;�a<��a<�a<��a<ܞa<Q�a<��a<��a<C�a<��a<֠a<�a<s�a<��a<�a<B�a<w�a<Ţa<�a<W�a<��a<ãa<��a<&�a<}�a<k�a<��a<��a<�a<��a<�a<(�a<A�a<`�a<n�a<��a<��a<��a<إa<�a<�a<�a<7�a<+�a<M�a<f�a<7�a<\�a<9�a<Q�a</�a<+�a<�a<�a<�a<�a<�a<�a<̥a<ϥa<��a<ƥa<��a<��a<d�a<x�a<X�a<�a<�a<ͤa<Ĥa<x�a<[�a<�a<��a<Σa<��a<x�a<M�a<�a<��a<ɢa<��a<f�a<Q�a<��a<�a<��a<L�a<�a<Ǡa<��a<*�a<�a<��a<E�a<�a<��a<Y�a<��a<��a<[�a<�a<a<[�a<�a<��a<g�a<њa<j�a<��a<��a<�a<��a<�a<��a<'�a<��a<*�a<��a<;�a<ɔa<R�a<�a<r�a<�a<��a<��a<��a<�a<��a<�a<��a<�a<��a<�a<��a<%�a<��a<4�a<Ћa<X�a<��a<��a<K�a<�a<��a<&�a<ˈa<��a<�a<χa<`�a<�a<��a<b�a<�a<ʅa<��a<A�a<�a<؄a<��a<|�a<I�a<B�a<�a<��a<a<��a<��a<j�a<w�a<A�a<L�a<"�a<�a<�a<	�a<�a<�a<�a<)�a<3�a<[�a<k�a<��a<�  �  ��a<�a<	�a<5�a<_�a<��a<̄a<ބa<#�a<U�a<��a<υa<��a<;�a<��a<Άa<2�a<��a<��a<O�a<��a<
�a<��a<�a<I�a<��a< �a<��a<��a<H�a<��a<1�a<��a<�a<��a<�a<��a<�a<��a<1�a<��a<D�a<Ԓa<a�a<ݓa<t�a<�a<��a<�a<q�a<�a<x�a<��a<{�a<ݘa<m�a<��a<R�a<�a<k�a<�a<T�a<˜a<I�a<a<�a<��a<�a<O�a<��a<��a<-�a<��a<��a<�a<Y�a<��a<�a<0�a<l�a<��a<�a<3�a<��a<��a< �a<+�a<U�a<��a<��a<äa<�a<�a<&�a<@�a<J�a<N�a<��a<��a<��a<ӥa<�a<��a<�a<�a<=�a<J�a<?�a<M�a<G�a<P�a<I�a<6�a<�a<)�a<�a<�a<�a<�a<Хa<ݥa<��a<ǥa<��a<��a<��a<��a<x�a<a�a<C�a<0�a<�a<Ϥa<��a<��a<i�a<9�a<��a<ƣa<��a<i�a<N�a<4�a<	�a<Ԣa<��a<j�a<T�a<�a<ѡa<��a<Z�a<�a<Ԡa<l�a<)�a<ݟa<y�a<<�a<�a<��a<@�a<��a<��a<f�a<��a<��a<e�a<�a<��a<H�a<Ϛa<{�a<�a<��a<�a<��a<*�a<��a<�a<��a<G�a<��a<N�a<ޔa<e�a<�a<n�a<�a<��a<�a<��a<	�a<��a<�a<��a<��a<��a<��a<��a<�a<��a<,�a<��a<M�a<�a<��a<'�a<�a<��a<1�a<Јa<r�a<�a<чa<d�a<�a<��a<w�a<+�a<Ӆa<z�a<e�a<�a<фa<��a<��a<^�a<6�a<�a<�a<�a<��a<��a<z�a<k�a<R�a<2�a<�a<�a<�a<�a<�a<��a<��a<%�a<!�a<T�a<_�a<��a<�  �  ��a<΃a<�a<3�a<f�a<��a<��a<�a<(�a<c�a<��a<ƅa<%�a<T�a<��a<�a<[�a<��a<��a<^�a<��a<:�a<|�a<�a<H�a<��a<"�a<u�a<�a<6�a<��a<�a<��a<��a<o�a<�a<Z�a<�a<{�a<#�a<��a<6�a<��a<L�a<�a<i�a<��a<{�a<�a<��a<�a<��a<�a<{�a<��a<t�a<��a<p�a<��a<W�a<�a<c�a<�a<X�a<��a<(�a<��a<�a<<�a<��a<�a<�a<��a<��a<�a<4�a<��a<סa<�a<x�a<��a<��a<!�a<��a<��a<��a<+�a<P�a<��a<��a<�a<��a<�a<)�a<0�a<n�a<m�a<��a<��a<ƥa<ʥa<٥a<�a<�a<E�a<.�a<A�a<J�a<I�a<W�a<9�a<<�a<,�a<�a<�a<��a<��a<ƥa<��a<��a<ťa<��a<��a<��a<��a<��a<{�a<��a<_�a<J�a<.�a<�a<�a<��a<��a<^�a<0�a<"�a<�a<��a<��a<x�a<$�a<�a<�a<��a<��a<D�a<�a<ѡa<��a<\�a<�a<àa<Z�a<$�a<ʟa<��a<�a<˞a<��a<�a<��a<��a<Y�a<�a<��a<P�a<��a<��a<<�a<�a<o�a<	�a<��a<�a<��a<�a<��a<;�a<��a<F�a<̕a<\�a<ʔa<m�a<��a<��a<�a<��a<�a<��a<�a<��a<��a<��a<�a<��a<�a<��a<�a<��a<�a<��a<X�a<ފa<��a<�a<ډa<p�a<)�a<ψa<m�a<&�a<��a<��a<(�a<φa<z�a<�a<��a<��a<d�a<�a<��a<��a<~�a<h�a<@�a<9�a<�a<كa<��a<��a<��a<T�a<E�a<(�a<�a<�a<�a<�a<˂a<�a<݂a<�a< �a<?�a<Z�a<��a<�  �  ��a<�a<��a<7�a<x�a<��a<Ȅa<��a<'�a<`�a<��a<ޅa<�a<h�a<��a<�a<G�a<��a<�a<\�a<��a<#�a<��a<�a<b�a<��a<�a<��a<ًa<W�a<��a<�a<y�a<��a<o�a<��a<u�a<�a<s�a<�a<��a<=�a<��a<f�a<ԓa<r�a< �a<��a<��a<��a<�a<��a<�a<}�a<�a<{�a<��a<��a<�a<��a<�a<b�a<֜a<D�a<��a<+�a<��a<ٞa<M�a<��a<�a<7�a<x�a<��a<��a<J�a<��a<ϡa<�a<T�a<��a<��a<E�a<r�a<ȣa<��a<�a<l�a<��a<��a<Ѥa<�a<�a<7�a<T�a<Y�a<��a<��a<��a<ɥa<إa<
�a<�a<�a<*�a<4�a<C�a<U�a<N�a<;�a<Z�a<,�a<5�a< �a<
�a<�a<�a<ޥa<ӥa<ťa<��a<��a<��a<��a<��a<��a<��a<l�a<b�a<\�a<,�a<�a<�a<��a<��a<��a<H�a<�a<��a<��a<��a<c�a<D�a<�a<�a<��a<��a<R�a<�a<�a<��a<P�a<�a<��a<|�a<�a<��a<d�a<�a<˞a<��a<3�a<ݝa<��a<J�a< �a<��a<O�a<�a<��a<F�a<�a<w�a<��a<��a< �a<��a<K�a<��a<K�a<Öa<F�a<�a<X�a<��a<t�a<�a<z�a<��a<��a<�a<��a<��a<��a<�a<��a<�a<x�a<�a<m�a<��a<��a<�a<��a<5�a<͊a<��a<9�a<ˉa<��a<*�a<Èa<��a< �a<Їa<r�a<�a<̆a<��a<>�a<�a<��a<\�a<1�a<��a<��a<��a<h�a<A�a<�a<��a<ۃa<ƃa<��a<m�a<v�a<5�a<0�a<�a<��a<߂a<�a<�a<�a<�a< �a<�a</�a<]�a<��a<�  �  ��a<�a<��a<L�a<c�a<��a<�a<�a<X�a<k�a<��a<�a<�a<{�a<��a<�a<>�a<��a<�a<q�a<�a<�a<��a<�a<T�a<��a<�a<{�a<��a<A�a<��a<1�a<|�a<�a<h�a<͎a<v�a<��a<��a<
�a<��a<�a<��a<]�a<Гa<��a<�a<��a<�a<��a<3�a<~�a<�a<�a<�a<��a<�a<��a<�a<��a<�a<��a<��a<[�a<۝a<�a<��a<؞a<C�a<w�a<ȟa<#�a<g�a<Ҡa<�a<H�a<o�a<áa<�a<N�a<Ģa<֢a<.�a<P�a<��a<�a<*�a<f�a<{�a<դa<Ѥa<�a<*�a<*�a<h�a<U�a<��a<��a<¥a<ȥa<�a<��a<�a<G�a<&�a<U�a<P�a<B�a<e�a</�a<R�a<�a<�a<�a<�a<�a<٥a<ޥa<��a<ĥa<��a<��a<��a<��a<��a<i�a<��a<^�a<w�a<G�a<2�a<.�a<�a<�a<��a<x�a<S�a<�a<�a<ͣa<��a<Z�a<W�a<�a<��a<ڢa<z�a<p�a<�a<ݡa<��a<B�a<�a<��a<e�a<��a<ݟa<g�a<�a<Þa<[�a<4�a<ɝa<��a<@�a<�a<��a<2�a<�a<��a<Z�a<̚a<��a<�a<��a<L�a<��a<L�a<��a<K�a<ٖa<^�a<�a<U�a<�a<i�a<�a<��a<�a<��a<��a<��a<��a<��a<�a<e�a<�a<f�a<	�a<\�a<��a<g�a<�a<��a<.�a<��a<j�a<!�a<��a<p�a<�a<Έa<��a<�a<��a<s�a<D�a<�a<{�a<S�a<݅a<Åa<t�a<C�a<��a<ʄa<��a<k�a<q�a<�a<�a<�a<��a<��a<a�a<m�a<�a<�a<��a<��a<��a<тa<�a<��a<��a<�a<�a<@�a<F�a<{�a<�  �  ��a<؃a<��a<G�a<d�a<��a<��a<�a<2�a<v�a<��a<��a<4�a<g�a<��a<�a<l�a<Ça<	�a<i�a<ƈa<#�a<~�a<�a<J�a<Ċa<�a<}�a<�a<L�a<��a<�a<l�a<�a<g�a<�a<j�a<܏a<k�a<��a<��a<9�a<Œa<O�a<�a<v�a<��a<�a<��a<��a<�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<��a<h�a<�a<E�a<��a<*�a<��a<�a<8�a<��a<�a<-�a<]�a<��a<�a<:�a<��a<ơa<�a<B�a<��a<Ԣa<<�a<��a<��a<�a<8�a<Y�a<��a<��a<Ӥa<��a<�a<6�a<c�a<��a<��a<��a<��a<ۥa<��a<��a<�a<"�a<2�a<*�a<I�a<I�a<Y�a<A�a<=�a<>�a<7�a<�a<�a<�a<ѥa<ץa<ɥa<��a<��a<��a<��a<��a<��a<��a<��a<l�a<r�a<H�a<6�a<�a<�a<Ȥa<��a<|�a<e�a<1�a<�a<ãa<��a<��a<\�a<�a<�a<��a<��a<F�a<�a<ӡa<��a<B�a<	�a< a<q�a<��a<��a<W�a<
�a<Þa<t�a<(�a<ŝa<|�a<.�a<��a<��a<V�a<��a<��a<J�a<ܚa<s�a<��a<��a<&�a<��a<@�a<ۗa<T�a<˖a<V�a<�a<~�a<��a<w�a<��a<��a<��a<��a<�a<��a<�a<��a<�a<��a<��a<\�a<ݍa<W�a<�a<z�a<�a<��a<"�a<͊a<g�a<0�a<ىa<x�a<�a<݈a<v�a<)�a<ȇa<t�a<'�a<Նa<��a<N�a<�a<��a<l�a<-�a<�a<�a<��a<x�a<L�a<&�a<�a<��a<��a<��a<t�a<Y�a<G�a<2�a<�a<߂a<ւa<ʂa<܂a<߂a<�a<�a<�a<�a<N�a<��a<�  �  ��a<Ѓa<	�a<$�a<j�a<��a<��a<@�a<�a<��a<��a<څa<�a<n�a<݆a<��a<Y�a<��a<!�a<q�a<��a<_�a<~�a<�a<?�a<��a<�a<r�a<ŋa<#�a<��a<�a<��a<��a<J�a<юa<X�a<��a<o�a<�a<��a<�a<��a<M�a<�a<Q�a<�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<(�a<{�a< �a<o�a<"�a<f�a<��a<i�a<Ýa<J�a<o�a<�a<8�a<��a<��a<�a<l�a<��a<�a<3�a<n�a<��a<�a<g�a<��a<�a<�a<X�a<��a<�a<+�a<D�a<��a<��a<�a<��a<"�a<Z�a<B�a<o�a<x�a<ɥa<��a<åa<�a<�a<1�a<�a<j�a<6�a<a�a<V�a<2�a<O�a<5�a<)�a<��a<�a<��a<�a<�a<��a<��a<��a<��a<��a<��a<��a<p�a<�a<}�a<w�a<O�a<N�a<Q�a<�a<0�a<��a<��a<��a<D�a<�a<��a<�a<��a<u�a<7�a<2�a<��a<��a<��a<F�a<9�a<ȡa<��a<H�a<��a<��a<G�a<�a<��a<y�a<�a<��a<`�a<�a<�a<��a<@�a<�a<y�a<J�a<��a<��a<$�a<��a<��a<�a<Ùa<�a<ݘa<2�a<a<C�a<�a<y�a<וa<g�a<�a<��a<��a<��a<!�a<��a<3�a<u�a<�a<��a<��a<S�a<܎a<k�a<֍a<z�a<�a<f�a<�a<��a<H�a<Ŋa<|�a<
�a<��a<p�a<�a<Јa<a�a<E�a<Ƈa<��a<*�a<߆a<��a<,�a<��a<��a<��a<<�a<��a<ʄa<��a<��a<9�a<_�a<��a<��a<ǃa<��a<��a<P�a<2�a<��a<�a<�a<�a<��a<��a<ɂa<ǂa<��a<�a<'�a<U�a<W�a<�  �  ��a<؃a<��a<G�a<d�a<��a<��a<�a<2�a<v�a<��a<��a<4�a<g�a<��a<�a<l�a<Ça<	�a<i�a<ƈa<#�a<~�a<�a<J�a<Ċa<�a<}�a<�a<L�a<��a<�a<l�a<�a<g�a<�a<j�a<܏a<k�a<��a<��a<9�a<Œa<O�a<�a<v�a<��a<�a<��a<��a<�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<��a<h�a<�a<E�a<��a<*�a<��a<�a<8�a<��a<�a<-�a<]�a<��a<�a<:�a<��a<ơa<�a<B�a<��a<Ԣa<<�a<��a<��a<�a<8�a<Y�a<��a<��a<Ӥa<��a<�a<6�a<c�a<��a<��a<��a<��a<ۥa<��a<��a<�a<"�a<2�a<*�a<I�a<I�a<Y�a<A�a<=�a<>�a<7�a<�a<�a<�a<ѥa<ץa<ɥa<��a<��a<��a<��a<��a<��a<��a<��a<l�a<r�a<H�a<6�a<�a<�a<Ȥa<��a<|�a<e�a<1�a<�a<ãa<��a<��a<\�a<�a<�a<��a<��a<F�a<�a<ӡa<��a<B�a<	�a< a<q�a<��a<��a<W�a<
�a<Þa<t�a<(�a<ŝa<|�a<.�a<��a<��a<V�a<��a<��a<J�a<ܚa<s�a<��a<��a<&�a<��a<@�a<ۗa<T�a<˖a<V�a<�a<~�a<��a<w�a<��a<��a<��a<��a<�a<��a<�a<��a<�a<��a<��a<\�a<ݍa<W�a<�a<z�a<�a<��a<"�a<͊a<g�a<0�a<ىa<x�a<�a<݈a<v�a<)�a<ȇa<t�a<'�a<Նa<��a<N�a<�a<��a<l�a<-�a<�a<�a<��a<x�a<L�a<&�a<�a<��a<��a<��a<t�a<Y�a<G�a<2�a<�a<߂a<ւa<ʂa<܂a<߂a<�a<�a<�a<�a<N�a<��a<�  �  ��a<�a<��a<L�a<c�a<��a<�a<�a<X�a<k�a<��a<�a<�a<{�a<��a<�a<>�a<��a<�a<q�a<�a<�a<��a<�a<T�a<��a<�a<{�a<��a<A�a<��a<1�a<|�a<�a<h�a<͎a<v�a<��a<��a<
�a<��a<�a<��a<]�a<Гa<��a<�a<��a<�a<��a<3�a<~�a<�a<�a<�a<��a<�a<��a<�a<��a<�a<��a<��a<[�a<۝a<�a<��a<؞a<C�a<w�a<ȟa<#�a<g�a<Ҡa<�a<H�a<o�a<áa<�a<N�a<Ģa<֢a<.�a<P�a<��a<�a<*�a<f�a<{�a<դa<Ѥa<�a<*�a<*�a<h�a<U�a<��a<��a<¥a<ȥa<�a<��a<�a<G�a<&�a<U�a<P�a<B�a<e�a</�a<R�a<�a<�a<�a<�a<�a<٥a<ޥa<��a<ĥa<��a<��a<��a<��a<��a<i�a<��a<^�a<w�a<G�a<2�a<.�a<�a<�a<��a<x�a<S�a<�a<�a<ͣa<��a<Z�a<W�a<�a<��a<ڢa<z�a<p�a<�a<ݡa<��a<B�a<�a<��a<e�a<��a<ݟa<g�a<�a<Þa<[�a<4�a<ɝa<��a<@�a<�a<��a<2�a<�a<��a<Z�a<̚a<��a<�a<��a<L�a<��a<L�a<��a<K�a<ٖa<^�a<�a<U�a<�a<i�a<�a<��a<�a<��a<��a<��a<��a<��a<�a<e�a<�a<f�a<	�a<\�a<��a<g�a<�a<��a<.�a<��a<j�a<!�a<��a<p�a<�a<Έa<��a<�a<��a<s�a<D�a<�a<{�a<S�a<݅a<Åa<t�a<C�a<��a<ʄa<��a<k�a<q�a<�a<�a<�a<��a<��a<a�a<m�a<�a<�a<��a<��a<��a<тa<�a<��a<��a<�a<�a<@�a<F�a<{�a<�  �  ��a<�a<��a<7�a<x�a<��a<Ȅa<��a<'�a<`�a<��a<ޅa<�a<h�a<��a<�a<G�a<��a<�a<\�a<��a<#�a<��a<�a<b�a<��a<�a<��a<ًa<W�a<��a<�a<y�a<��a<o�a<��a<u�a<�a<s�a<�a<��a<=�a<��a<f�a<ԓa<r�a< �a<��a<��a<��a<�a<��a<�a<}�a<�a<{�a<��a<��a<�a<��a<�a<b�a<֜a<D�a<��a<+�a<��a<ٞa<M�a<��a<�a<7�a<x�a<��a<��a<J�a<��a<ϡa<�a<T�a<��a<��a<E�a<r�a<ȣa<��a<�a<l�a<��a<��a<Ѥa<�a<�a<7�a<T�a<Y�a<��a<��a<��a<ɥa<إa<
�a<�a<�a<*�a<4�a<C�a<U�a<N�a<;�a<Z�a<,�a<5�a< �a<
�a<�a<�a<ޥa<ӥa<ťa<��a<��a<��a<��a<��a<��a<��a<l�a<b�a<\�a<,�a<�a<�a<��a<��a<��a<H�a<�a<��a<��a<��a<c�a<D�a<�a<�a<��a<��a<R�a<�a<�a<��a<P�a<�a<��a<|�a<�a<��a<d�a<�a<˞a<��a<3�a<ݝa<��a<J�a< �a<��a<O�a<�a<��a<F�a<�a<w�a<��a<��a< �a<��a<K�a<��a<K�a<Öa<F�a<�a<X�a<��a<t�a<�a<z�a<��a<��a<�a<��a<��a<��a<�a<��a<�a<x�a<�a<m�a<��a<��a<�a<��a<5�a<͊a<��a<9�a<ˉa<��a<*�a<Èa<��a< �a<Їa<r�a<�a<̆a<��a<>�a<�a<��a<\�a<1�a<��a<��a<��a<h�a<A�a<�a<��a<ۃa<ƃa<��a<m�a<v�a<5�a<0�a<�a<��a<߂a<�a<�a<�a<�a< �a<�a</�a<]�a<��a<�  �  ��a<΃a<�a<3�a<f�a<��a<��a<�a<(�a<c�a<��a<ƅa<%�a<T�a<��a<�a<[�a<��a<��a<^�a<��a<:�a<|�a<�a<H�a<��a<"�a<u�a<�a<6�a<��a<�a<��a<��a<o�a<�a<Z�a<�a<{�a<#�a<��a<6�a<��a<L�a<�a<i�a<��a<{�a<�a<��a<�a<��a<�a<{�a<��a<t�a<��a<p�a<��a<W�a<�a<c�a<�a<X�a<��a<(�a<��a<�a<<�a<��a<�a<�a<��a<��a<�a<4�a<��a<סa<�a<x�a<��a<��a<!�a<��a<��a<��a<+�a<P�a<��a<��a<�a<��a<�a<)�a<0�a<n�a<m�a<��a<��a<ƥa<ʥa<٥a<�a<�a<E�a<.�a<A�a<J�a<I�a<W�a<9�a<<�a<,�a<�a<�a<��a<��a<ƥa<��a<��a<ťa<��a<��a<��a<��a<��a<{�a<��a<_�a<J�a<.�a<�a<�a<��a<��a<^�a<0�a<"�a<�a<��a<��a<x�a<$�a<�a<�a<��a<��a<D�a<�a<ѡa<��a<\�a<�a<àa<Z�a<$�a<ʟa<��a<�a<˞a<��a<�a<��a<��a<Y�a<�a<��a<P�a<��a<��a<<�a<�a<o�a<	�a<��a<�a<��a<�a<��a<;�a<��a<F�a<̕a<\�a<ʔa<m�a<��a<��a<�a<��a<�a<��a<�a<��a<��a<��a<�a<��a<�a<��a<�a<��a<�a<��a<X�a<ފa<��a<�a<ډa<p�a<)�a<ψa<m�a<&�a<��a<��a<(�a<φa<z�a<�a<��a<��a<d�a<�a<��a<��a<~�a<h�a<@�a<9�a<�a<كa<��a<��a<��a<T�a<E�a<(�a<�a<�a<�a<�a<˂a<�a<݂a<�a< �a<?�a<Z�a<��a<�  �  ��a<�a<	�a<5�a<_�a<��a<̄a<ބa<#�a<U�a<��a<υa<��a<;�a<��a<Άa<2�a<��a<��a<O�a<��a<
�a<��a<�a<I�a<��a< �a<��a<��a<H�a<��a<1�a<��a<�a<��a<�a<��a<�a<��a<1�a<��a<D�a<Ԓa<a�a<ݓa<t�a<�a<��a<�a<q�a<�a<x�a<��a<{�a<ݘa<m�a<��a<R�a<�a<k�a<�a<T�a<˜a<I�a<a<�a<��a<�a<O�a<��a<��a<-�a<��a<��a<�a<Y�a<��a<�a<0�a<l�a<��a<�a<3�a<��a<��a< �a<+�a<U�a<��a<��a<äa<�a<�a<&�a<@�a<J�a<N�a<��a<��a<��a<ӥa<�a<��a<�a<�a<=�a<J�a<?�a<M�a<G�a<P�a<I�a<6�a<�a<)�a<�a<�a<�a<�a<Хa<ݥa<��a<ǥa<��a<��a<��a<��a<x�a<a�a<C�a<0�a<�a<Ϥa<��a<��a<i�a<9�a<��a<ƣa<��a<i�a<N�a<4�a<	�a<Ԣa<��a<j�a<T�a<�a<ѡa<��a<Z�a<�a<Ԡa<l�a<)�a<ݟa<y�a<<�a<�a<��a<@�a<��a<��a<f�a<��a<��a<e�a<�a<��a<H�a<Ϛa<{�a<�a<��a<�a<��a<*�a<��a<�a<��a<G�a<��a<N�a<ޔa<e�a<�a<n�a<�a<��a<�a<��a<	�a<��a<�a<��a<��a<��a<��a<��a<�a<��a<,�a<��a<M�a<�a<��a<'�a<�a<��a<1�a<Јa<r�a<�a<чa<d�a<�a<��a<w�a<+�a<Ӆa<z�a<e�a<�a<фa<��a<��a<^�a<6�a<�a<�a<�a<��a<��a<z�a<k�a<R�a<2�a<�a<�a<�a<�a<�a<��a<��a<%�a<!�a<T�a<_�a<��a<�  �  ��a<�a<��a<M�a<t�a<x�a<Ʉa<܄a<.�a<B�a<��a<��a<�a<B�a<��a<܆a<1�a<��a<�a<D�a<��a<�a<��a<͉a<i�a<��a<�a<��a<�a<o�a<��a<9�a<��a< �a<��a<�a<��a<�a<��a<%�a<��a<M�a<ʒa<j�a<ӓa<��a<�a<v�a<��a<x�a<��a<i�a<�a<\�a<�a<Z�a<ٙa<e�a<Ԛa<U�a<Лa<U�a<Μa<;�a<��a<�a<��a<ܞa<Q�a<��a<��a<C�a<��a<֠a<�a<s�a<��a<�a<B�a<w�a<Ţa<�a<W�a<��a<ãa<��a<&�a<}�a<k�a<��a<��a<�a<��a<�a<(�a<A�a<`�a<n�a<��a<��a<��a<إa<�a<�a<�a<7�a<+�a<M�a<f�a<7�a<\�a<9�a<Q�a</�a<+�a<�a<�a<�a<�a<�a<�a<̥a<ϥa<��a<ƥa<��a<��a<d�a<x�a<X�a<�a<�a<ͤa<Ĥa<x�a<[�a<�a<��a<Σa<��a<x�a<M�a<�a<��a<ɢa<��a<f�a<Q�a<��a<�a<��a<L�a<�a<Ǡa<��a<*�a<�a<��a<E�a<�a<��a<Y�a<��a<��a<[�a<�a<a<[�a<�a<��a<g�a<њa<j�a<��a<��a<�a<��a<�a<��a<'�a<��a<*�a<��a<;�a<ɔa<R�a<�a<r�a<�a<��a<��a<��a<�a<��a<�a<��a<�a<��a<�a<��a<%�a<��a<4�a<Ћa<X�a<��a<��a<K�a<�a<��a<&�a<ˈa<��a<�a<χa<`�a<�a<��a<b�a<�a<ʅa<��a<A�a<�a<؄a<��a<|�a<I�a<B�a<�a<��a<a<��a<��a<j�a<w�a<A�a<L�a<"�a<�a<�a<	�a<�a<�a<�a<)�a<3�a<[�a<k�a<��a<�  �  ��a<��a<�a<4�a<`�a<��a<��a<�a<
�a<9�a<��a<��a<��a<*�a<�a<��a<.�a<o�a<�a<0�a<��a<�a<�a<ۉa<P�a<��a<.�a<��a<�a<a�a<ӌa<K�a<a<�a<��a<4�a<��a<"�a<��a<<�a<��a<H�a<Вa<k�a<�a<l�a<�a<~�a<�a<��a<ۖa<l�a<ٗa<S�a<Ҙa<S�a<Йa<J�a<̚a<@�a<כa<<�a<՜a<@�a<��a<�a<��a<�a<W�a<��a<��a<F�a<��a<�a<.�a<^�a<͡a<�a<8�a<��a<ۢa<�a<K�a<��a<ѣa<
�a<"�a<_�a<x�a<��a<ʤa<�a<�a<�a<�a<A�a<E�a<d�a<|�a<��a<��a<ѥa<�a<�a<�a<*�a<9�a<F�a<H�a<T�a<`�a<=�a<B�a<;�a<;�a<.�a<�a<��a<�a<�a<ܥa<�a<ݥa<ťa<��a<��a<��a<��a<`�a<D�a<"�a<�a<ݤa<��a<p�a<T�a<�a<��a<��a<��a<\�a<K�a<�a<��a<��a<��a<u�a<F�a<�a<١a<��a<h�a<%�a<��a<��a<=�a<��a<��a<>�a<��a<a<F�a<�a<Ɲa<r�a<�a<��a<a�a<�a<��a<?�a<ךa<r�a<��a<��a<��a<��a<�a<��a<�a<��a<"�a<��a<3�a<��a<Y�a<͓a<x�a<��a<��a<�a<��a<�a<��a<�a<��a<�a<��a<$�a<��a<�a<Ča<C�a<Ƌa<z�a<�a<��a<>�a<ۉa<��a<<�a<ƈa<|�a<�a<Ƈa<k�a<�a<��a<l�a< �a<ʅa<q�a<8�a<��a<фa<��a<u�a<F�a<�a<�a<�a<уa<��a<��a<��a<{�a<F�a<>�a<.�a<*�a<�a<�a<��a<+�a<�a<#�a<L�a<j�a<|�a<��a<�  �  �a<�a<�a<9�a<^�a<��a<��a<�a<��a<5�a<j�a<��a<��a<�a<��a<��a<�a<e�a<؇a<%�a<��a<�a<g�a<�a<I�a<��a<$�a<��a<�a<m�a<ތa<9�a<��a<>�a<��a<2�a<��a<B�a<��a<@�a<͑a<`�a<�a<Z�a<�a<f�a<��a<s�a<�a<m�a<ɖa<e�a<ȗa<^�a<��a<D�a<ʙa<)�a<Ϛa<2�a<Λa<'�a<��a<+�a<��a<$�a<��a<��a<G�a<��a<�a<V�a<��a<ؠa<B�a<~�a<ʡa<�a<Z�a<��a<Ǣa<�a<\�a<��a<Σa<��a<3�a<U�a<��a<��a<��a<դa<֤a<�a<�a<2�a<�a<n�a<^�a<��a<��a<��a<ݥa<�a<�a<�a<@�a<@�a<I�a<Y�a<O�a<o�a<O�a<K�a<7�a<�a<:�a<�a<�a<��a<	�a<ڥa<ԥa<եa<��a<ͥa<��a<��a<e�a<B�a<0�a<�a<Ҥa<��a<k�a<=�a<�a<ݣa<��a<��a<9�a<6�a<��a<�a<��a<��a<e�a</�a<�a<ҡa<��a<^�a<�a<��a<��a<H�a<�a<��a<c�a<�a<��a<f�a<+�a<��a<v�a<$�a<՜a<��a<�a<��a<9�a<ښa<h�a<�a<|�a<�a<��a<��a<��a<�a<��a<�a<��a<6�a<��a<O�a<��a<c�a<�a<z�a<�a<��a<�a<��a<*�a<��a<"�a<��a<�a<��a<1�a<��a<L�a<�a<u�a<��a<��a<P�a<
�a<��a</�a<؈a<r�a<#�a<��a<V�a<�a<��a<]�a<�a<��a<J�a<B�a<߄a<��a<��a<`�a<B�a<�a<�a<݃a<؃a<��a<��a<��a<k�a<x�a<J�a<>�a<&�a<�a<3�a<�a<*�a<(�a<P�a<A�a<a�a<��a<��a<�  �  уa<�a<�a<N�a<_�a<�a<Äa<҄a<�a<4�a<Y�a<��a<ׅa<�a<j�a<��a<�a<Z�a<ˇa<5�a<��a<��a<��a<ωa<P�a<Êa<(�a<��a<�a<p�a<ތa<l�a<Ía<F�a<��a<+�a<��a<0�a<ʐa<K�a<ʑa<P�a<ؒa<l�a<�a<��a<�a<y�a<��a<b�a<�a<Z�a<��a<9�a<��a<7�a<��a<;�a<��a<+�a<��a<G�a<��a<;�a<��a<�a<��a<�a<U�a<��a<��a<S�a<��a<�a<:�a<��a<ȡa<�a<g�a<��a<��a<�a<_�a<��a<ƣa<�a<7�a<]�a<o�a<��a<��a<ݤa<�a<��a<��a< �a<;�a<T�a<c�a<~�a<��a<��a<եa< �a<�a<3�a</�a<=�a<b�a<R�a<]�a<Y�a<K�a<I�a<S�a<<�a<'�a<*�a<
�a<�a<��a<��a<��a<Хa<��a<��a<��a<��a<z�a<C�a<�a<	�a<äa<��a<j�a<,�a<��a<ԣa<��a<��a<T�a<'�a<�a<ܢa<��a<��a<X�a<P�a<��a<١a<��a<b�a<�a<۠a<��a<H�a<�a<��a<k�a<�a<��a<|�a<�a<۝a<��a<!�a<Ɯa<i�a<�a<��a<T�a<˚a<m�a<��a<q�a<�a<~�a<�a<o�a< �a<�a<�a<��a<�a<��a<@�a<ٓa<b�a<�a<��a<��a<��a<�a<��a<�a<��a<�a<��a<=�a<��a<I�a<��a<W�a<��a<z�a<3�a<��a<S�a<�a<��a<6�a<܈a<y�a<	�a<̇a<Q�a<	�a<��a<N�a<�a<��a<f�a<(�a<�a<��a<u�a<M�a<:�a<)�a<��a<��a<ǃa<��a<��a<��a<x�a<b�a<F�a<<�a<C�a<.�a< �a</�a< �a<=�a<C�a<[�a<��a<��a<��a<�  �  ƃa<�a<�a<9�a<s�a<r�a<��a<��a<��a<�a<q�a<��a<˅a<�a<9�a<��a<��a<t�a<̇a<�a<��a<݈a<��a<ĉa<e�a<��a<8�a<��a< �a<��a<یa<a�a<ʍa<G�a<Ύa<C�a<Џa<-�a<ސa<>�a<�a<x�a<ߒa<��a<ߓa<}�a<�a<i�a<ܕa<@�a<Ֆa<=�a<�a<0�a<��a<'�a<��a<8�a<��a<S�a<��a<3�a<��a<�a<��a<�a<��a<��a<s�a<��a<"�a<z�a<��a<�a<7�a<��a<�a<+�a<f�a<��a<��a<�a<��a<��a<�a<�a< �a<r�a<h�a<��a<��a<��a<פa<��a<�a<�a<:�a<'�a<_�a<v�a<��a<̥a<��a<�a<�a<"�a<!�a<O�a<Q�a<O�a<z�a<M�a<x�a<Z�a<E�a<N�a<�a<?�a<!�a<$�a<�a<�a<�a<ߥa<�a<��a<��a<��a<e�a<W�a<	�a<��a<��a<��a<S�a<D�a<�a<ȣa<��a<N�a<S�a<�a<�a<ݢa<��a<��a<=�a<G�a<�a<�a<��a<r�a<:�a<ڠa<àa<F�a<�a<��a<l�a<)�a<Ҟa<��a<�a<�a<t�a<>�a<�a<p�a<6�a<��a<P�a<Қa<^�a<ޙa<O�a<�a<a�a<�a<f�a<��a<o�a<�a<��a<	�a<ǔa<*�a<ēa<@�a<Ԓa<{�a<��a<��a<�a<��a<'�a<��a<F�a<��a<L�a<��a<P�a<،a<l�a<��a<~�a</�a<��a<��a<��a<��a<I�a<Ĉa<��a<�a<ća<5�a<�a<��a<H�a<�a<��a<f�a<��a<߄a<��a<}�a<p�a<�a<�a<Ճa<�a<��a<��a<��a<��a<��a<V�a<s�a<M�a<5�a<@�a<�a<C�a<6�a<P�a<:�a<i�a<w�a<��a<Ӄa<�  �  Ӄa<�a< �a<8�a<r�a<}�a<��a<݄a<�a<#�a<K�a<��a<��a<�a<_�a<��a<�a<Q�a<��a<'�a<��a<�a<j�a<؉a<W�a<��a<+�a<��a<�a<z�a<�a<[�a<�a<V�a<��a<;�a<a<Y�a<֐a<L�a<ёa<[�a<ےa<d�a<��a<p�a<��a<d�a<�a<m�a<�a<:�a<��a<&�a<��a<.�a<��a<)�a<��a<%�a<��a<?�a<��a<3�a<��a<%�a<��a<��a<O�a<��a<
�a<Y�a<��a<�a<`�a<��a<ءa<�a<r�a<¢a<�a<-�a<g�a<��a<��a<�a<.�a<a�a<{�a<��a<��a<ؤa<�a<�a<��a<�a<0�a<E�a<]�a<j�a<��a<��a<��a<��a<�a<"�a<&�a<S�a<J�a<`�a<O�a<Y�a<X�a<Y�a<L�a<V�a<K�a<+�a<�a<�a<�a<�a<�a<�a<ɥa<��a<��a<��a<d�a<V�a<�a<��a<ͤa<��a<Y�a<�a<�a<��a<��a<u�a<K�a<�a<�a<��a<��a<��a<h�a<1�a<�a<�a<��a<e�a<�a<�a<��a<W�a<�a<՟a<{�a<�a<ɞa<�a<B�a<�a<��a<(�a<Мa<l�a<�a<��a<D�a<�a<Y�a<�a<|�a<��a<^�a<�a<\�a<�a<v�a< �a<��a<�a<��a<$�a<ѓa<d�a<�a<s�a<�a<��a<�a<��a<�a<��a<%�a<��a<?�a<Ӎa<J�a<Ќa<Z�a< �a<��a<$�a<��a<[�a<��a<��a<3�a<ӈa<~�a<�a<��a<\�a<�a<��a<3�a<��a<��a<\�a<�a<݄a<��a<j�a<F�a<"�a<!�a<�a<�a<��a<ăa<��a<��a<j�a<b�a<S�a<L�a<<�a<H�a<C�a<0�a<,�a<=�a<_�a<x�a<|�a<��a<��a<�  �  ��a<��a<ۂa<�a<�a<D�a<L�a<]�a<{�a<كa<�a<9�a<g�a<��a<��a<%�a<��a<��a<c�a<نa<�a<��a<�a<��a<�a<��a<�a<d�a<��a<:�a<��a<�a<��a<�a<��a<�a<��a<&�a<��a<G�a<��a<M�a<��a<>�a<��a<P�a<�a<O�a<Ɣa<�a<��a<C�a<��a<7�a<w�a<�a<��a<�a<��a<�a<��a<�a<��a<&�a<��a<;�a<��a<&�a<]�a<�a<9�a<��a<�a<��a<i�a<��a<��a<<�a<}�a<��a<�a<l�a<x�a<ۢa<��a<�a<e�a<^�a<��a<��a<��a<��a<ۣa<�a<�a<�a<��a<9�a<5�a<V�a<��a<��a<Ҥa<��a<ޤa<�a<A�a<Z�a<X�a<{�a<S�a<��a<d�a<w�a<`�a<:�a<I�a<.�a<3�a<�a<�a<��a<��a<�a<Ѥa<��a<��a<��a<q�a<S�a</�a<�a<��a<c�a<a�a<�a<��a<��a<l�a<`�a<�a<�a<�a<��a<��a<L�a<D�a<)�a<#�a<ՠa<��a<q�a<3�a<�a<��a<��a<��a<��a<{�a<0�a<��a<�a<B�a<Ȝa<��a<D�a<�a<��a<�a<ۚa<A�a<�a<Z�a<ۘa<6�a<��a<o�a<Öa<m�a<��a<H�a<Ҕa<:�a<�a<h�a<�a<��a<�a<��a<J�a<��a<d�a<�a<s�a<'�a<��a<�a<��a<�a<��a<�a<��a<5�a<Êa<P�a<Ӊa<��a<�a<�a<k�a<��a<��a<+�a<�a<[�a<�a<t�a<D�a<�a<��a<R�a<̓a<��a<_�a<2�a<$�a<�a<߂a<��a<{�a<��a<��a<s�a<O�a<U�a<�a<H�a<�a<�a<��a<Ӂa<�a<ځa<��a<�a<�a<�a<)�a<e�a<`�a<�  �  ��a<��a<Ђa<�a<�a<'�a<Z�a<��a<��a<a<��a<�a<T�a<��a<�a<9�a<��a<�a<L�a<Ɇa<Y�a<ȇa<!�a<��a<�a<w�a<�a<i�a<Ίa<7�a<��a<1�a<��a<!�a<��a<�a<��a<4�a<��a<+�a<��a<:�a<Αa<Q�a<ْa<U�a<ۓa<E�a<ݔa<Z�a<��a<!�a<��a<�a<��a<�a<��a<��a<��a< �a<��a<0�a<̛a<F�a<��a<+�a<��a<�a<l�a<͞a<�a<x�a<ȟa<%�a<~�a<��a<�a<=�a<��a<ڡa<�a<A�a<r�a<��a<�a<�a<?�a<e�a<��a<��a<Σa<�a<ԣa<ѣa<�a<�a<
�a<(�a<?�a<P�a<d�a<��a<��a<��a<�a<(�a<'�a<N�a<N�a<e�a<i�a<f�a<[�a<b�a<T�a<^�a<N�a<>�a<+�a<$�a<�a<�a<��a<�a<Ȥa<��a<��a<��a<c�a<N�a<�a<��a<ԣa<��a<J�a<�a<΢a<��a<z�a<N�a<!�a<�a<ˡa<��a<��a<��a<q�a<0�a<�a<٠a<��a<q�a<8�a<�a<��a<`�a<�a<ߞa<��a<2�a<ٝa<��a<P�a<��a<��a<=�a<ٛa<��a<�a<��a<F�a<ڙa<P�a<�a<x�a<�a<M�a<��a<8�a<��a<F�a<̔a<J�a<֓a<\�a<��a<��a<M�a<ّa<J�a<�a<n�a<��a<��a<�a<}�a<�a<��a<�a<��a< �a<��a<6�a<̊a<q�a<��a<��a<�a<��a<e�a<��a<��a<1�a<φa<c�a<�a<��a<=�a<΄a<w�a<&�a<��a<��a<j�a<,�a<��a<ւa<Ȃa<ǂa<��a<��a<f�a<g�a<E�a<?�a<+�a<�a<��a<��a<�a<��a<�a<�a<�a<��a<�a<*�a<*�a<I�a<X�a<�  �  v�a<Ăa<ɂa<�a<�a<+�a<d�a<[�a<��a<��a<�a<+�a<g�a<��a<Ԅa<\�a<��a<�a<w�a<��a<9�a<��a<3�a<��a<�a<n�a<��a<u�a<Ŋa<f�a<��a<,�a<��a<��a<��a<�a<��a<��a<��a<�a<Аa<P�a<đa<l�a<��a<g�a<ѓa<[�a<ʔa<.�a<��a<�a<��a<�a<��a<�a<��a<*�a<��a<:�a<��a<�a<��a<)�a<��a<�a<��a<�a<��a<ɞa<(�a<��a<��a<!�a<=�a<��a<�a<:�a<j�a<��a<	�a<&�a<��a<��a<��a<)�a<2�a<z�a<z�a<��a<��a<��a<��a<�a<�a<�a</�a<�a<O�a<q�a<w�a<��a<��a<٤a<�a<'�a<1�a<L�a<[�a<Y�a<��a<[�a<~�a<a�a<>�a<Q�a< �a<:�a<�a<"�a<��a<�a<�a<�a<�a<��a<Ƥa<��a<h�a<P�a<�a<��a<��a<��a<>�a<:�a<�a<��a<��a<8�a<D�a<�a<�a<ԡa<��a<x�a<=�a<B�a<��a<�a<��a<x�a<D�a<�a<ʟa<L�a<�a<��a<_�a<*�a<ӝa<��a<�a<�a<w�a<S�a<�a<|�a<9�a<��a<X�a<Йa<e�a<ߘa<L�a<Ηa<E�a<�a<>�a<�a<H�a<ǔa<v�a<ԓa<��a<�a<��a<"�a<��a<c�a<ܐa<��a<�a<��a<�a<��a<&�a<o�a<�a<m�a<�a<��a<3�a<��a<9�a<��a<m�a<E�a<��a<m�a<�a<��a<F�a<a<w�a<�a<��a<&�a<�a<��a<&�a<�a<��a<z�a<M�a<	�a<�a<��a<��a<}�a<��a<q�a<d�a<R�a<3�a<K�a<
�a<!�a<��a<Ձa<�a<��a<�a<ہa<��a<�a<�a<�a<B�a<��a<�  �  y�a<��a<ła<��a<�a<A�a<h�a<y�a<��a<Ӄa< �a<$�a<l�a<��a<��a<K�a<��a<�a<e�a<܆a<[�a<��a<@�a<��a<�a<��a<�a<Z�a<Ŋa<9�a<��a<'�a<��a<*�a<}�a<�a<��a<�a<��a<$�a<��a<*�a<Ña<N�a<֒a<k�a<ʓa<n�a<єa<R�a<וa<,�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<I�a<ƛa<5�a<̜a<�a<��a<�a<e�a<Ğa<�a<n�a<��a<�a<T�a<��a<ՠa<�a<��a<��a<�a<6�a<t�a<��a<�a<�a<K�a<s�a<~�a<��a<��a<�a<�a<�a<�a<
�a<�a<8�a<I�a<g�a<}�a<��a<¤a< �a<�a<)�a<K�a<C�a<g�a<]�a<^�a<[�a<V�a<X�a<K�a<I�a<C�a<+�a<��a<�a<�a<��a<�a<�a<̤a<��a<��a<��a<w�a<D�a<,�a<�a<��a<��a<[�a<$�a<ߢa<��a<��a<^�a<4�a<�a<֡a<��a<��a<��a<V�a<O�a<�a<�a<��a<g�a<(�a<��a<��a<V�a<�a<��a<��a<�a<��a<��a<-�a<�a<��a<2�a<ɛa<z�a<�a<��a<\�a<șa<y�a<�a<p�a<��a<X�a<Жa<L�a<ѕa<Q�a<ڔa<b�a<�a<v�a<�a<��a<G�a<Ǒa<r�a<אa<��a<��a<{�a<��a<o�a<��a<��a<�a<��a<"�a<��a<�a<Պa<J�a<�a<}�a<�a<��a<W�a<�a<��a<?�a<Ɔa<��a<�a<��a<R�a<�a<��a<>�a<��a<��a<t�a<C�a<�a<�a<ςa<ӂa<��a<��a<��a<[�a<^�a<7�a< �a<�a<��a<�a<�a<�a<�a<ׁa<��a<�a<�a<�a<!�a<C�a<\�a<�  �  ��a<��a<ςa<�a<�a<D�a<A�a<��a<��a<ڃa<
�a<Q�a<��a<��a<!�a<<�a<Ӆa<�a<v�a<׆a<Z�a<��a<�a<��a<�a<�a<�a<a�a<ۊa<"�a<��a<�a<{�a<�a<n�a< �a<n�a<�a<u�a<#�a<��a<0�a<ڑa<G�a<ݒa<X�a<��a<[�a<��a<]�a<��a<D�a<��a<M�a<��a</�a<��a<�a<ϙa<'�a<��a<-�a<̛a<+�a<��a<3�a<��a<	�a<a�a<؞a<�a<h�a<��a<�a<S�a<��a<֠a<�a<^�a<��a<ޡa<>�a<a�a<��a<�a<�a<D�a<f�a<��a<��a<��a<�a<ޣa<��a<�a<A�a<�a<^�a<R�a<~�a<��a<��a<Ӥa<�a<�a<�a<E�a<M�a<V�a<g�a<X�a<s�a<J�a<\�a<B�a<�a<.�a<
�a<�a<�a<��a<Ӥa<ݤa<�a<��a<̤a<��a<��a<l�a<J�a</�a<ۣa<֣a<��a<b�a<.�a<�a<ڢa<��a<��a<%�a<;�a<��a<ҡa<��a<��a<h�a<*�a<�a<ڠa<��a<k�a</�a<��a<��a<]�a<�a<��a<a�a<�a<ŝa<`�a<)�a<��a<��a<-�a<Λa<��a<�a<��a<H�a<ߙa<f�a<Ҙa<{�a<ߗa<p�a<ݖa<��a<֕a<o�a<��a<_�a<"�a<��a<"�a<��a<M�a<��a<Z�a<�a<r�a<��a<w�a<�a<|�a<��a<��a<ߌa<��a<�a<��a<�a<��a<9�a<ˉa<��a<�a<a<d�a<��a<��a<2�a<݆a<f�a<�a<��a<G�a<��a<��a<v�a<�a<܃a<|�a<Z�a<=�a<��a<��a<Ăa<��a<r�a<��a<f�a<L�a<B�a<�a<#�a<�a<��a<فa<��a<΁a<��a<؁a<ǁa<�a<�a<�a<F�a<H�a<�  �  h�a<��a<͂a<�a<�a<E�a<g�a<��a<��a<�a<+�a<=�a<��a<Ȅa<#�a<e�a<ȅa<�a<��a<�a<O�a<a<5�a<��a<�a<�a<�a<E�a<��a<(�a<��a<�a<��a<ٌa<k�a<��a<L�a<��a<��a<�a<��a<$�a<��a<K�a<֒a<]�a<�a<^�a<ܔa<c�a<��a<f�a<a<8�a<��a<6�a<��a<1�a<��a<8�a<�a<*�a<қa<A�a<��a<6�a<��a<�a<i�a<��a<�a<[�a<��a<��a<H�a<]�a<۠a<�a<5�a<��a<�a< �a<c�a<��a<̢a<�a<B�a<k�a<��a<��a<ģa<ߣa<�a<'�a<�a<1�a<:�a<Y�a<f�a<��a<��a<ˤa<�a<�a<�a<,�a<C�a<V�a<Z�a<e�a<Y�a<J�a<M�a<;�a<9�a</�a<�a<�a<�a<�a<�a<�a<ݤa<��a<��a<��a<��a<��a<p�a<R�a<1�a<�a<գa<��a<u�a<N�a<��a<�a<��a<��a<M�a<1�a<�a< �a<��a<��a<k�a<D�a<�a<ߠa<��a<q�a<�a<͟a<��a<>�a<��a<��a<9�a<��a<ĝa<>�a<�a<ǜa<t�a<�a<Ûa<a�a<�a<��a<N�a<�a<i�a<�a<��a<ԗa<��a<�a<n�a<�a<v�a<��a<}�a<�a<��a<J�a<��a<S�a<ԑa<b�a<�a<v�a<��a<�a<�a<g�a<�a<k�a<�a<x�a<̋a<��a<�a<{�a<:�a<͉a<g�a<	�a<��a<@�a< �a<��a<7�a<߆a<x�a<�a<��a<N�a<$�a<��a<e�a<�a<׃a<��a<k�a<(�a<�a<��a<��a<��a<��a<��a<n�a<Q�a<?�a<�a<��a<��a<Ձa<Ёa<ǁa<��a<��a<сa<��a<ҁa<��a<�a< �a<N�a<�  �  g�a<��a<��a<�a<�a<:�a<y�a<��a<߃a<�a<)�a<V�a<��a<�a<"�a<��a<܅a<#�a<��a<�a<}�a<ʇa<F�a<��a<�a<x�a<݉a<R�a<��a<+�a<�a<�a<e�a<�a<L�a<ƍa<a�a<�a<c�a<��a<��a<6�a<��a<N�a<Òa<b�a<ړa<e�a<�a<s�a<�a<X�a<ϖa<R�a<ԗa<@�a<��a<Q�a<әa<K�a<Қa<U�a<�a<H�a<Ȝa<(�a<��a<��a<c�a<��a<�a<N�a<��a<ٟa<-�a<s�a<��a<�a<F�a<��a<ơa<�a<^�a<��a<Ңa<�a<9�a<s�a<��a<ãa<ͣa<�a<��a<�a<�a<C�a<]�a<\�a<{�a<��a<��a<Фa<�a<�a<&�a<>�a<>�a<M�a<Y�a<N�a<a�a<I�a<[�a<'�a<!�a<�a<�a<��a<ܤa<ݤa<ݤa<��a<¤a<��a<ˤa<��a<��a<z�a<j�a<L�a<%�a<�a<ۣa<ǣa<p�a<M�a<�a<��a<��a<��a<m�a<E�a<�a<�a<��a<��a<s�a<U�a<�a<�a<��a<[�a<!�a<ٟa<��a<(�a<ܞa<��a<D�a<��a<��a<T�a<�a<��a<b�a<�a<ԛa<b�a<�a<��a<S�a<ٙa<p�a<��a<��a<
�a<��a< �a<��a<�a<��a<�a<��a<'�a<��a<9�a<Ȓa<i�a<ۑa<o�a<�a<~�a<�a<y�a<�a<{�a<ލa<Z�a<Ќa<]�a<�a<U�a<�a<��a<�a<��a<U�a<�a<��a<F�a<�a<��a<?�a<φa<��a<�a<݅a<c�a<�a<��a<w�a<4�a<ۃa<��a<��a<E�a<�a<�a<�a<Âa<��a<~�a<f�a<P�a<(�a<$�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<́a<́a<��a<�a<[�a<�  �  a�a<��a<Ƃa<�a<�a<P�a<n�a<��a<Ӄa<��a<D�a<��a<��a<�a<Z�a<x�a<�a<M�a<��a<�a<m�a<ʇa<?�a<��a<�a<�a<މa<C�a<��a<��a<��a<�a<I�a<όa<:�a<��a<>�a<юa<J�a<�a<n�a<�a<��a<:�a<Ӓa<Z�a<�a<x�a<ߔa<a�a<�a<j�a<�a<n�a<��a<l�a<�a<=�a<�a<g�a<�a<a�a<қa<D�a<Ӝa<6�a<��a<�a<S�a<��a< �a<)�a<��a<ğa<�a<R�a<��a<�a<,�a<k�a<��a<�a<%�a<��a<ʢa<�a<C�a<m�a<��a<��a<̣a<�a<�a<,�a<D�a<Y�a<J�a<��a<��a<��a<Ԥa<�a<��a<�a<�a</�a<T�a<S�a<X�a<^�a<P�a<C�a<,�a<�a<0�a<�a<��a<ڤa<ߤa<��a<Ǥa<��a<Ȥa<��a<��a<��a<��a<��a<n�a<R�a<;�a<�a<٣a<��a<��a<h�a<;�a<��a<Ƣa<��a<a�a<U�a<2�a<�a<ҡa<��a<s�a<N�a<"�a<�a<��a<[�a<�a<Οa<[�a<3�a<՞a<o�a<.�a<ϝa<��a<1�a<�a<��a<q�a<�a<��a<Z�a<�a<��a<K�a<�a<��a<��a<�a<�a<��a<�a<��a<��a<��a<7�a<��a<C�a<Óa<K�a<Ԓa<T�a<בa<y�a<�a<u�a<��a<i�a<ߎa<c�a<��a<j�a<��a<E�a<��a<M�a<܊a<r�a<�a<��a<b�a<̈a<��a<>�a<�a<��a<9�a<�a<��a<�a<˅a<t�a<)�a<ڄa<��a< �a<�a<��a<y�a<f�a<7�a<�a<�a<��a<��a<��a<l�a<O�a<8�a<�a<�a<ρa<��a<ǁa<��a<��a<��a<��a<��a<��a<��a<��a<�a<+�a<�  �  c�a<l�a<a<�a<�a<O�a<z�a<��a<ʃa<"�a<B�a<m�a<Ʉa<��a<`�a<��a<��a<8�a<��a<!�a<k�a<�a<<�a<��a<�a<x�a<��a<�a<��a<�a<o�a<ыa<]�a<��a<,�a<Ǎa<�a<�a<C�a<��a<h�a<�a<��a<,�a<Ӓa<U�a<�a<k�a<�a<��a<�a<��a<�a<p�a<�a<g�a<�a<b�a<��a<\�a<��a<k�a<�a<q�a<ɜa<<�a<��a<�a<I�a<��a<��a<(�a<��a<��a<(�a<1�a<��a<٠a<�a<��a<��a<��a<3�a<��a<��a<�a<<�a<h�a<��a<��a<��a<��a<"�a<=�a<2�a<j�a<j�a<��a<��a<��a<Ǥa<�a<�a<
�a<G�a<G�a<Q�a<T�a<R�a<Y�a<2�a<A�a<6�a<�a<�a<��a<��a<��a<ܤa<��a<Ĥa<��a<��a<��a<��a<��a<n�a<��a<h�a<P�a<:�a<�a<�a<��a<��a<e�a<'�a<�a<բa<Ģa<|�a<h�a<�a<�a<�a<��a<��a<K�a<$�a<ݠa<��a<]�a<�a<͟a<i�a<�a<��a<��a<�a<��a<��a<
�a< �a<��a<D�a<�a<��a<R�a<��a<��a<F�a<�a<v�a<�a<��a<�a<��a<�a<��a<#�a<��a<1�a<��a<K�a<��a<c�a<ޒa<m�a<�a<o�a<��a<q�a<��a<_�a<͎a<_�a<��a<A�a<��a<Y�a<��a<S�a<Ҋa<X�a<�a<��a<B�a<ڈa<��a<�a<�a<��a<4�a<�a<��a<J�a<Ӆa<��a<:�a<Ȅa<��a<@�a<�a<Ńa<��a<Y�a<4�a<&�a<܂a<�a<��a<��a<m�a<I�a<3�a<�a<�a<؁a<��a<��a<��a<��a<a�a<��a<v�a<��a<ǁa<ځa<��a<1�a<�  �  I�a<��a<��a<�a< �a<G�a<w�a<��a<�a<�a<S�a<��a<�a<�a<D�a<��a<�a<g�a<��a<�a<t�a<އa<C�a<��a<"�a<k�a<�a<?�a<��a<�a<[�a<ǋa<.�a<��a<�a<��a<"�a<��a<1�a<Ϗa<w�a<�a<��a<J�a<��a<c�a<�a<j�a<��a<p�a<��a<}�a<
�a<}�a<�a<p�a<�a<��a<��a<��a<��a<u�a<ޛa<`�a<˜a<<�a<��a<�a<d�a<��a<��a<A�a<k�a<��a<�a<8�a<}�a<��a<	�a<L�a<��a<�a<O�a<��a<��a<�a<)�a<~�a<��a<��a<�a<��a<&�a<@�a<_�a<r�a<��a<��a<��a<�a<�a< �a<�a<"�a</�a<B�a<K�a<Z�a<W�a<K�a<X�a<,�a<9�a<�a<��a<Ҥa<Τa<Ťa<��a<��a<��a<��a<��a<��a<��a<��a<��a<�a<c�a<X�a<2�a<�a<�a<ʣa<��a<v�a<N�a<5�a<�a<��a<��a<y�a<L�a<�a<�a<��a<��a<R�a<�a<�a<��a<j�a<�a<��a<|�a<�a<��a<T�a<�a<��a<g�a<�a<ɜa<r�a<3�a<��a<��a<L�a<�a<��a<S�a<�a<u�a<�a<��a<$�a<��a<;�a<��a<W�a<��a<4�a<�a<O�a<�a<_�a<�a<_�a<�a<r�a<��a<�a<ۏa<z�a<юa<Y�a<эa<,�a<��a< �a<��a</�a<��a<N�a<�a<��a<+�a<��a<��a<5�a<��a<}�a<J�a<�a<��a<2�a<҅a<��a<=�a<��a<��a<l�a<�a<փa<ăa<y�a<N�a< �a<��a<̂a<��a<��a<s�a<N�a<%�a<�a<ہa<܁a<��a<��a<k�a<m�a<q�a<r�a<��a<��a<��a<΁a<��a<6�a<�  �  -�a<��a<��a<�a<�a<O�a<��a<��a<
�a<�a<O�a<��a<a<(�a<c�a<Åa<��a<r�a<��a<+�a<��a<݇a<l�a<��a<�a<q�a<щa<;�a<v�a<�a<G�a<�a<%�a<��a< �a<��a<2�a<��a<T�a<ҏa<J�a<�a<��a<:�a<��a<i�a<֓a<��a<	�a<|�a<)�a<m�a<�a<i�a<��a<��a<�a<��a<�a<��a<�a<��a<�a<i�a<�a<$�a<��a<�a<U�a<��a<ўa<�a<d�a<ɟa<ٟa<H�a<f�a<��a<�a<A�a<��a<Сa<!�a<]�a<��a<��a</�a<w�a<��a<�a<�a<�a<A�a<.�a<l�a<V�a<��a<��a<��a<��a<�a<�a<	�a<O�a<.�a<_�a<W�a<E�a<`�a<?�a<N�a<�a<�a<�a<
�a<�a<��a<Ѥa<��a<��a<��a<��a<��a<{�a<��a<i�a<��a<l�a<o�a<I�a<:�a<4�a<�a<�a<��a<s�a<S�a<�a<�a<Ǣa<��a<Y�a<W�a<�a<��a<ۡa<��a<{�a<�a<�a<��a<O�a<
�a<��a<S�a<�a<Оa<K�a<�a<��a<G�a<$�a<��a<��a<6�a<͛a<��a<8�a<�a<��a<Z�a<ՙa<��a<�a<��a<N�a<��a<C�a<��a<6�a<͕a<R�a<͔a<9�a<�a<N�a<�a<t�a<��a<��a<�a<��a<ޏa<k�a<Ďa<4�a<��a<%�a<��a<	�a<��a<�a<��a<c�a<؉a<��a<�a<Ȉa<h�a<0�a<އa<��a<C�a<φa<��a<3�a<��a<��a<+�a<�a<��a<k�a< �a<�a<��a<u�a<P�a<�a<"�a<˂a<˂a<��a<^�a<W�a<�a<�a<��a<��a<��a<��a<��a<[�a<}�a<J�a<��a<��a<��a<�a<ہa<�a<�  �  d�a<��a<��a<�a<�a<R�a<��a<��a<݃a<#�a<]�a<��a<�a<+�a<o�a<ƅa<"�a<|�a<Æa<)�a<~�a<�a<M�a<��a<�a<w�a<ĉa<B�a<��a<	�a<U�a<��a<�a<��a<�a<��a<�a<��a<"�a<��a<b�a<�a<��a<&�a<Œa<S�a<�a<v�a<�a<{�a< �a<��a<�a<��a<�a<��a<
�a<��a<&�a<��a<�a<z�a<�a<j�a<Ӝa<8�a<��a<��a<=�a<��a<��a<)�a<Z�a<��a<ܟa<�a<p�a<��a<��a<7�a<��a<ۡa<9�a<��a<ˢa<�a<8�a<f�a<��a<ƣa<�a<�a<0�a<F�a<s�a<��a<��a<��a<ʤa<�a<�a<
�a<�a<�a<8�a<P�a<U�a<K�a<Q�a<F�a<=�a<F�a<5�a<�a<ۤa<Ǥa<��a<��a<��a<��a<��a<�a<y�a<��a<��a<��a<��a<k�a<h�a<G�a<>�a<�a<��a<ģa<��a<��a<m�a<4�a<�a<Ӣa<��a<��a<a�a< �a<��a<��a<��a<\�a<#�a<֠a<��a<B�a<�a<şa<m�a<��a<��a<;�a<�a<��a<Y�a<��a<��a<c�a<�a<�a<��a<e�a<�a<��a<D�a<�a<��a<�a<��a<%�a<��a<I�a<ۖa<P�a<͕a<O�a<ޔa<z�a<�a<i�a<�a<j�a<��a<z�a<��a<m�a<�a<S�a<�a<_�a<��a<�a<��a<�a<��a<"�a<��a<:�a<Ήa<m�a<"�a<��a<��a<?�a<̇a<��a<2�a<�a<��a<>�a<�a<��a<C�a<	�a<Ąa<p�a<(�a<��a<��a<��a<X�a<(�a<�a<Ղa<��a<��a<d�a<H�a<!�a< �a<��a<؁a<��a<r�a<_�a<T�a<\�a<b�a<l�a<w�a<��a<��a<�a<4�a<�  �  1�a<r�a<ǂa<�a<!�a<Z�a<r�a<�a<�a<D�a<U�a<��a<�a<#�a<x�a<��a<�a<T�a<ӆa<;�a<��a<�a<8�a<͈a<�a<��a<݉a<0�a<o�a<؊a<n�a<��a<D�a<��a<�a<��a<��a<Ďa<+�a<ӏa<c�a<ΐa<�a<�a<ܒa<M�a<	�a<n�a<�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<�a<g�a<+�a<��a<�a<��a<Ɯa<Y�a<��a<	�a<9�a<��a<��a<�a<{�a<��a<�a<�a<x�a<��a<�a<j�a<��a<��a<�a<K�a<��a<��a<D�a<e�a<��a<��a<�a<�a<;�a<_�a<H�a<��a<��a<��a<Ǥa<ޤa<�a<��a<C�a<$�a<h�a<E�a<W�a<g�a<M�a<d�a<3�a<�a<�a<�a<�a<ߤa<٤a<��a<��a<��a<��a<��a<��a<��a<b�a<l�a<t�a<��a<k�a<Y�a<E�a<�a<+�a<̣a<̣a<y�a<K�a<1�a<��a<ۢa<��a<��a<9�a</�a<�a<ơa<��a<G�a<>�a<ޠa<��a<Z�a<��a<��a<=�a<�a<��a<k�a<�a<��a<g�a<�a<��a<m�a<7�a<�a<m�a<7�a<�a<��a<=�a<�a<y�a<%�a<Ęa<-�a<ߗa<�a<��a<F�a<̕a<R�a<єa<`�a<Óa<��a<��a<��a<�a<m�a<�a<d�a<��a<N�a<��a<�a<��a<<�a<��a<C�a<}�a<)�a<��a<3�a<�a<v�a<A�a<��a<V�a<*�a<݇a<��a<1�a<�a<y�a<g�a<��a<��a<\�a<ބa<��a<`�a</�a<�a<��a<w�a<B�a<P�a<��a<�a<��a<��a<��a<D�a<?�a<��a<ǁa<��a<��a<��a<x�a<y�a<K�a<v�a<\�a<��a<��a<��a<��a<�a<�  �  d�a<��a<��a<�a<�a<R�a<��a<��a<݃a<#�a<]�a<��a<�a<+�a<o�a<ƅa<"�a<|�a<Æa<)�a<~�a<�a<M�a<��a<�a<w�a<ĉa<B�a<��a<	�a<U�a<��a<�a<��a<�a<��a<�a<��a<"�a<��a<b�a<�a<��a<&�a<Œa<S�a<�a<v�a<�a<{�a< �a<��a<�a<��a<�a<��a<
�a<��a<&�a<��a<�a<z�a<�a<j�a<Ӝa<8�a<��a<��a<=�a<��a<��a<)�a<Z�a<��a<ܟa<�a<p�a<��a<��a<7�a<��a<ۡa<9�a<��a<ˢa<�a<8�a<f�a<��a<ƣa<�a<�a<0�a<F�a<s�a<��a<��a<��a<ʤa<�a<�a<
�a<�a<�a<8�a<P�a<U�a<K�a<Q�a<F�a<=�a<F�a<5�a<�a<ۤa<Ǥa<��a<��a<��a<��a<��a<�a<y�a<��a<��a<��a<��a<k�a<h�a<G�a<>�a<�a<��a<ģa<��a<��a<m�a<4�a<�a<Ӣa<��a<��a<a�a< �a<��a<��a<��a<\�a<#�a<֠a<��a<B�a<�a<şa<m�a<��a<��a<;�a<�a<��a<Y�a<��a<��a<c�a<�a<�a<��a<e�a<�a<��a<D�a<�a<��a<�a<��a<%�a<��a<I�a<ۖa<P�a<͕a<O�a<ޔa<z�a<�a<i�a<�a<j�a<��a<z�a<��a<m�a<�a<S�a<�a<_�a<��a<�a<��a<�a<��a<"�a<��a<:�a<Ήa<m�a<"�a<��a<��a<?�a<̇a<��a<2�a<�a<��a<>�a<�a<��a<C�a<	�a<Ąa<p�a<(�a<��a<��a<��a<X�a<(�a<�a<Ղa<��a<��a<d�a<H�a<!�a< �a<��a<؁a<��a<r�a<_�a<T�a<\�a<b�a<l�a<w�a<��a<��a<�a<4�a<�  �  -�a<��a<��a<�a<�a<O�a<��a<��a<
�a<�a<O�a<��a<a<(�a<c�a<Åa<��a<r�a<��a<+�a<��a<݇a<l�a<��a<�a<q�a<щa<;�a<v�a<�a<G�a<�a<%�a<��a< �a<��a<2�a<��a<T�a<ҏa<J�a<�a<��a<:�a<��a<i�a<֓a<��a<	�a<|�a<)�a<m�a<�a<i�a<��a<��a<�a<��a<�a<��a<�a<��a<�a<i�a<�a<$�a<��a<�a<U�a<��a<ўa<�a<d�a<ɟa<ٟa<H�a<f�a<��a<�a<A�a<��a<Сa<!�a<]�a<��a<��a</�a<w�a<��a<�a<�a<�a<A�a<.�a<l�a<V�a<��a<��a<��a<��a<�a<�a<	�a<O�a<.�a<_�a<W�a<E�a<`�a<?�a<N�a<�a<�a<�a<
�a<�a<��a<Ѥa<��a<��a<��a<��a<��a<{�a<��a<i�a<��a<l�a<o�a<I�a<:�a<4�a<�a<�a<��a<s�a<S�a<�a<�a<Ǣa<��a<Y�a<W�a<�a<��a<ۡa<��a<{�a<�a<�a<��a<O�a<
�a<��a<S�a<�a<Оa<K�a<�a<��a<G�a<$�a<��a<��a<6�a<͛a<��a<8�a<�a<��a<Z�a<ՙa<��a<�a<��a<N�a<��a<C�a<��a<6�a<͕a<R�a<͔a<9�a<�a<N�a<�a<t�a<��a<��a<�a<��a<ޏa<k�a<Ďa<4�a<��a<%�a<��a<	�a<��a<�a<��a<c�a<؉a<��a<�a<Ȉa<h�a<0�a<އa<��a<C�a<φa<��a<3�a<��a<��a<+�a<�a<��a<k�a< �a<�a<��a<u�a<P�a<�a<"�a<˂a<˂a<��a<^�a<W�a<�a<�a<��a<��a<��a<��a<��a<[�a<}�a<J�a<��a<��a<��a<�a<ہa<�a<�  �  I�a<��a<��a<�a< �a<G�a<w�a<��a<�a<�a<S�a<��a<�a<�a<D�a<��a<�a<g�a<��a<�a<t�a<އa<C�a<��a<"�a<k�a<�a<?�a<��a<�a<[�a<ǋa<.�a<��a<�a<��a<"�a<��a<1�a<Ϗa<w�a<�a<��a<J�a<��a<c�a<�a<j�a<��a<p�a<��a<}�a<
�a<}�a<�a<p�a<�a<��a<��a<��a<��a<u�a<ޛa<`�a<˜a<<�a<��a<�a<d�a<��a<��a<A�a<k�a<��a<�a<8�a<}�a<��a<	�a<L�a<��a<�a<O�a<��a<��a<�a<)�a<~�a<��a<��a<�a<��a<&�a<@�a<_�a<r�a<��a<��a<��a<�a<�a< �a<�a<"�a</�a<B�a<K�a<Z�a<W�a<K�a<X�a<,�a<9�a<�a<��a<Ҥa<Τa<Ťa<��a<��a<��a<��a<��a<��a<��a<��a<��a<�a<c�a<X�a<2�a<�a<�a<ʣa<��a<v�a<N�a<5�a<�a<��a<��a<y�a<L�a<�a<�a<��a<��a<R�a<�a<�a<��a<j�a<�a<��a<|�a<�a<��a<T�a<�a<��a<g�a<�a<ɜa<r�a<3�a<��a<��a<L�a<�a<��a<S�a<�a<u�a<�a<��a<$�a<��a<;�a<��a<W�a<��a<4�a<�a<O�a<�a<_�a<�a<_�a<�a<r�a<��a<�a<ۏa<z�a<юa<Y�a<эa<,�a<��a< �a<��a</�a<��a<N�a<�a<��a<+�a<��a<��a<5�a<��a<}�a<J�a<�a<��a<2�a<҅a<��a<=�a<��a<��a<l�a<�a<փa<ăa<y�a<N�a< �a<��a<̂a<��a<��a<s�a<N�a<%�a<�a<ہa<܁a<��a<��a<k�a<m�a<q�a<r�a<��a<��a<��a<΁a<��a<6�a<�  �  c�a<l�a<a<�a<�a<O�a<z�a<��a<ʃa<"�a<B�a<m�a<Ʉa<��a<`�a<��a<��a<8�a<��a<!�a<k�a<�a<<�a<��a<�a<x�a<��a<�a<��a<�a<o�a<ыa<]�a<��a<,�a<Ǎa<�a<�a<C�a<��a<h�a<�a<��a<,�a<Ӓa<U�a<�a<k�a<�a<��a<�a<��a<�a<p�a<�a<g�a<�a<b�a<��a<\�a<��a<k�a<�a<q�a<ɜa<<�a<��a<�a<I�a<��a<��a<(�a<��a<��a<(�a<1�a<��a<٠a<�a<��a<��a<��a<3�a<��a<��a<�a<<�a<h�a<��a<��a<��a<��a<"�a<=�a<2�a<j�a<j�a<��a<��a<��a<Ǥa<�a<�a<
�a<G�a<G�a<Q�a<T�a<R�a<Y�a<2�a<A�a<6�a<�a<�a<��a<��a<��a<ܤa<��a<Ĥa<��a<��a<��a<��a<��a<n�a<��a<h�a<P�a<:�a<�a<�a<��a<��a<e�a<'�a<�a<բa<Ģa<|�a<h�a<�a<�a<�a<��a<��a<K�a<$�a<ݠa<��a<]�a<�a<͟a<i�a<�a<��a<��a<�a<��a<��a<
�a< �a<��a<D�a<�a<��a<R�a<��a<��a<F�a<�a<v�a<�a<��a<�a<��a<�a<��a<#�a<��a<1�a<��a<K�a<��a<c�a<ޒa<m�a<�a<o�a<��a<q�a<��a<_�a<͎a<_�a<��a<A�a<��a<Y�a<��a<S�a<Ҋa<X�a<�a<��a<B�a<ڈa<��a<�a<�a<��a<4�a<�a<��a<J�a<Ӆa<��a<:�a<Ȅa<��a<@�a<�a<Ńa<��a<Y�a<4�a<&�a<܂a<�a<��a<��a<m�a<I�a<3�a<�a<�a<؁a<��a<��a<��a<��a<a�a<��a<v�a<��a<ǁa<ځa<��a<1�a<�  �  a�a<��a<Ƃa<�a<�a<P�a<n�a<��a<Ӄa<��a<D�a<��a<��a<�a<Z�a<x�a<�a<M�a<��a<�a<m�a<ʇa<?�a<��a<�a<�a<މa<C�a<��a<��a<��a<�a<I�a<όa<:�a<��a<>�a<юa<J�a<�a<n�a<�a<��a<:�a<Ӓa<Z�a<�a<x�a<ߔa<a�a<�a<j�a<�a<n�a<��a<l�a<�a<=�a<�a<g�a<�a<a�a<қa<D�a<Ӝa<6�a<��a<�a<S�a<��a< �a<)�a<��a<ğa<�a<R�a<��a<�a<,�a<k�a<��a<�a<%�a<��a<ʢa<�a<C�a<m�a<��a<��a<̣a<�a<�a<,�a<D�a<Y�a<J�a<��a<��a<��a<Ԥa<�a<��a<�a<�a</�a<T�a<S�a<X�a<^�a<P�a<C�a<,�a<�a<0�a<�a<��a<ڤa<ߤa<��a<Ǥa<��a<Ȥa<��a<��a<��a<��a<��a<n�a<R�a<;�a<�a<٣a<��a<��a<h�a<;�a<��a<Ƣa<��a<a�a<U�a<2�a<�a<ҡa<��a<s�a<N�a<"�a<�a<��a<[�a<�a<Οa<[�a<3�a<՞a<o�a<.�a<ϝa<��a<1�a<�a<��a<q�a<�a<��a<Z�a<�a<��a<K�a<�a<��a<��a<�a<�a<��a<�a<��a<��a<��a<7�a<��a<C�a<Óa<K�a<Ԓa<T�a<בa<y�a<�a<u�a<��a<i�a<ߎa<c�a<��a<j�a<��a<E�a<��a<M�a<܊a<r�a<�a<��a<b�a<̈a<��a<>�a<�a<��a<9�a<�a<��a<�a<˅a<t�a<)�a<ڄa<��a< �a<�a<��a<y�a<f�a<7�a<�a<�a<��a<��a<��a<l�a<O�a<8�a<�a<�a<ρa<��a<ǁa<��a<��a<��a<��a<��a<��a<��a<��a<�a<+�a<�  �  g�a<��a<��a<�a<�a<:�a<y�a<��a<߃a<�a<)�a<V�a<��a<�a<"�a<��a<܅a<#�a<��a<�a<}�a<ʇa<F�a<��a<�a<x�a<݉a<R�a<��a<+�a<�a<�a<e�a<�a<L�a<ƍa<a�a<�a<c�a<��a<��a<6�a<��a<N�a<Òa<b�a<ړa<e�a<�a<s�a<�a<X�a<ϖa<R�a<ԗa<@�a<��a<Q�a<әa<K�a<Қa<U�a<�a<H�a<Ȝa<(�a<��a<��a<c�a<��a<�a<N�a<��a<ٟa<-�a<s�a<��a<�a<F�a<��a<ơa<�a<^�a<��a<Ңa<�a<9�a<s�a<��a<ãa<ͣa<�a<��a<�a<�a<C�a<]�a<\�a<{�a<��a<��a<Фa<�a<�a<&�a<>�a<>�a<M�a<Y�a<N�a<a�a<I�a<[�a<'�a<!�a<�a<�a<��a<ܤa<ݤa<ݤa<��a<¤a<��a<ˤa<��a<��a<z�a<j�a<L�a<%�a<�a<ۣa<ǣa<p�a<M�a<�a<��a<��a<��a<m�a<E�a<�a<�a<��a<��a<s�a<U�a<�a<�a<��a<[�a<!�a<ٟa<��a<(�a<ܞa<��a<D�a<��a<��a<T�a<�a<��a<b�a<�a<ԛa<b�a<�a<��a<S�a<ٙa<p�a<��a<��a<
�a<��a< �a<��a<�a<��a<�a<��a<'�a<��a<9�a<Ȓa<i�a<ۑa<o�a<�a<~�a<�a<y�a<�a<{�a<ލa<Z�a<Ќa<]�a<�a<U�a<�a<��a<�a<��a<U�a<�a<��a<F�a<�a<��a<?�a<φa<��a<�a<݅a<c�a<�a<��a<w�a<4�a<ۃa<��a<��a<E�a<�a<�a<�a<Âa<��a<~�a<f�a<P�a<(�a<$�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<́a<́a<��a<�a<[�a<�  �  h�a<��a<͂a<�a<�a<E�a<g�a<��a<��a<�a<+�a<=�a<��a<Ȅa<#�a<e�a<ȅa<�a<��a<�a<O�a<a<5�a<��a<�a<�a<�a<E�a<��a<(�a<��a<�a<��a<ٌa<k�a<��a<L�a<��a<��a<�a<��a<$�a<��a<K�a<֒a<]�a<�a<^�a<ܔa<c�a<��a<f�a<a<8�a<��a<6�a<��a<1�a<��a<8�a<�a<*�a<қa<A�a<��a<6�a<��a<�a<i�a<��a<�a<[�a<��a<��a<H�a<]�a<۠a<�a<5�a<��a<�a< �a<c�a<��a<̢a<�a<B�a<k�a<��a<��a<ģa<ߣa<�a<'�a<�a<1�a<:�a<Y�a<f�a<��a<��a<ˤa<�a<�a<�a<,�a<C�a<V�a<Z�a<e�a<Y�a<J�a<M�a<;�a<9�a</�a<�a<�a<�a<�a<�a<�a<ݤa<��a<��a<��a<��a<��a<p�a<R�a<1�a<�a<գa<��a<u�a<N�a<��a<�a<��a<��a<M�a<1�a<�a< �a<��a<��a<k�a<D�a<�a<ߠa<��a<q�a<�a<͟a<��a<>�a<��a<��a<9�a<��a<ĝa<>�a<�a<ǜa<t�a<�a<Ûa<a�a<�a<��a<N�a<�a<i�a<�a<��a<ԗa<��a<�a<n�a<�a<v�a<��a<}�a<�a<��a<J�a<��a<S�a<ԑa<b�a<�a<v�a<��a<�a<�a<g�a<�a<k�a<�a<x�a<̋a<��a<�a<{�a<:�a<͉a<g�a<	�a<��a<@�a< �a<��a<7�a<߆a<x�a<�a<��a<N�a<$�a<��a<e�a<�a<׃a<��a<k�a<(�a<�a<��a<��a<��a<��a<��a<n�a<Q�a<?�a<�a<��a<��a<Ձa<Ёa<ǁa<��a<��a<сa<��a<ҁa<��a<�a< �a<N�a<�  �  ��a<��a<ςa<�a<�a<D�a<A�a<��a<��a<ڃa<
�a<Q�a<��a<��a<!�a<<�a<Ӆa<�a<v�a<׆a<Z�a<��a<�a<��a<�a<�a<�a<a�a<ۊa<"�a<��a<�a<{�a<�a<n�a< �a<n�a<�a<u�a<#�a<��a<0�a<ڑa<G�a<ݒa<X�a<��a<[�a<��a<]�a<��a<D�a<��a<M�a<��a</�a<��a<�a<ϙa<'�a<��a<-�a<̛a<+�a<��a<3�a<��a<	�a<a�a<؞a<�a<h�a<��a<�a<S�a<��a<֠a<�a<^�a<��a<ޡa<>�a<a�a<��a<�a<�a<D�a<f�a<��a<��a<��a<�a<ޣa<��a<�a<A�a<�a<^�a<R�a<~�a<��a<��a<Ӥa<�a<�a<�a<E�a<M�a<V�a<g�a<X�a<s�a<J�a<\�a<B�a<�a<.�a<
�a<�a<�a<��a<Ӥa<ݤa<�a<��a<̤a<��a<��a<l�a<J�a</�a<ۣa<֣a<��a<b�a<.�a<�a<ڢa<��a<��a<%�a<;�a<��a<ҡa<��a<��a<h�a<*�a<�a<ڠa<��a<k�a</�a<��a<��a<]�a<�a<��a<a�a<�a<ŝa<`�a<)�a<��a<��a<-�a<Λa<��a<�a<��a<H�a<ߙa<f�a<Ҙa<{�a<ߗa<p�a<ݖa<��a<֕a<o�a<��a<_�a<"�a<��a<"�a<��a<M�a<��a<Z�a<�a<r�a<��a<w�a<�a<|�a<��a<��a<ߌa<��a<�a<��a<�a<��a<9�a<ˉa<��a<�a<a<d�a<��a<��a<2�a<݆a<f�a<�a<��a<G�a<��a<��a<v�a<�a<܃a<|�a<Z�a<=�a<��a<��a<Ăa<��a<r�a<��a<f�a<L�a<B�a<�a<#�a<�a<��a<فa<��a<΁a<��a<؁a<ǁa<�a<�a<�a<F�a<H�a<�  �  y�a<��a<ła<��a<�a<A�a<h�a<y�a<��a<Ӄa< �a<$�a<l�a<��a<��a<K�a<��a<�a<e�a<܆a<[�a<��a<@�a<��a<�a<��a<�a<Z�a<Ŋa<9�a<��a<'�a<��a<*�a<}�a<�a<��a<�a<��a<$�a<��a<*�a<Ña<N�a<֒a<k�a<ʓa<n�a<єa<R�a<וa<,�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<I�a<ƛa<5�a<̜a<�a<��a<�a<e�a<Ğa<�a<n�a<��a<�a<T�a<��a<ՠa<�a<��a<��a<�a<6�a<t�a<��a<�a<�a<K�a<s�a<~�a<��a<��a<�a<�a<�a<�a<
�a<�a<8�a<I�a<g�a<}�a<��a<¤a< �a<�a<)�a<K�a<C�a<g�a<]�a<^�a<[�a<V�a<X�a<K�a<I�a<C�a<+�a<��a<�a<�a<��a<�a<�a<̤a<��a<��a<��a<w�a<D�a<,�a<�a<��a<��a<[�a<$�a<ߢa<��a<��a<^�a<4�a<�a<֡a<��a<��a<��a<V�a<O�a<�a<�a<��a<g�a<(�a<��a<��a<V�a<�a<��a<��a<�a<��a<��a<-�a<�a<��a<2�a<ɛa<z�a<�a<��a<\�a<șa<y�a<�a<p�a<��a<X�a<Жa<L�a<ѕa<Q�a<ڔa<b�a<�a<v�a<�a<��a<G�a<Ǒa<r�a<אa<��a<��a<{�a<��a<o�a<��a<��a<�a<��a<"�a<��a<�a<Պa<J�a<�a<}�a<�a<��a<W�a<�a<��a<?�a<Ɔa<��a<�a<��a<R�a<�a<��a<>�a<��a<��a<t�a<C�a<�a<�a<ςa<ӂa<��a<��a<��a<[�a<^�a<7�a< �a<�a<��a<�a<�a<�a<�a<ׁa<��a<�a<�a<�a<!�a<C�a<\�a<�  �  v�a<Ăa<ɂa<�a<�a<+�a<d�a<[�a<��a<��a<�a<+�a<g�a<��a<Ԅa<\�a<��a<�a<w�a<��a<9�a<��a<3�a<��a<�a<n�a<��a<u�a<Ŋa<f�a<��a<,�a<��a<��a<��a<�a<��a<��a<��a<�a<Аa<P�a<đa<l�a<��a<g�a<ѓa<[�a<ʔa<.�a<��a<�a<��a<�a<��a<�a<��a<*�a<��a<:�a<��a<�a<��a<)�a<��a<�a<��a<�a<��a<ɞa<(�a<��a<��a<!�a<=�a<��a<�a<:�a<j�a<��a<	�a<&�a<��a<��a<��a<)�a<2�a<z�a<z�a<��a<��a<��a<��a<�a<�a<�a</�a<�a<O�a<q�a<w�a<��a<��a<٤a<�a<'�a<1�a<L�a<[�a<Y�a<��a<[�a<~�a<a�a<>�a<Q�a< �a<:�a<�a<"�a<��a<�a<�a<�a<�a<��a<Ƥa<��a<h�a<P�a<�a<��a<��a<��a<>�a<:�a<�a<��a<��a<8�a<D�a<�a<�a<ԡa<��a<x�a<=�a<B�a<��a<�a<��a<x�a<D�a<�a<ʟa<L�a<�a<��a<_�a<*�a<ӝa<��a<�a<�a<w�a<S�a<�a<|�a<9�a<��a<X�a<Йa<e�a<ߘa<L�a<Ηa<E�a<�a<>�a<�a<H�a<ǔa<v�a<ԓa<��a<�a<��a<"�a<��a<c�a<ܐa<��a<�a<��a<�a<��a<&�a<o�a<�a<m�a<�a<��a<3�a<��a<9�a<��a<m�a<E�a<��a<m�a<�a<��a<F�a<a<w�a<�a<��a<&�a<�a<��a<&�a<�a<��a<z�a<M�a<	�a<�a<��a<��a<}�a<��a<q�a<d�a<R�a<3�a<K�a<
�a<!�a<��a<Ձa<�a<��a<�a<ہa<��a<�a<�a<�a<B�a<��a<�  �  ��a<��a<Ђa<�a<�a<'�a<Z�a<��a<��a<a<��a<�a<T�a<��a<�a<9�a<��a<�a<L�a<Ɇa<Y�a<ȇa<!�a<��a<�a<w�a<�a<i�a<Ίa<7�a<��a<1�a<��a<!�a<��a<�a<��a<4�a<��a<+�a<��a<:�a<Αa<Q�a<ْa<U�a<ۓa<E�a<ݔa<Z�a<��a<!�a<��a<�a<��a<�a<��a<��a<��a< �a<��a<0�a<̛a<F�a<��a<+�a<��a<�a<l�a<͞a<�a<x�a<ȟa<%�a<~�a<��a<�a<=�a<��a<ڡa<�a<A�a<r�a<��a<�a<�a<?�a<e�a<��a<��a<Σa<�a<ԣa<ѣa<�a<�a<
�a<(�a<?�a<P�a<d�a<��a<��a<��a<�a<(�a<'�a<N�a<N�a<e�a<i�a<f�a<[�a<b�a<T�a<^�a<N�a<>�a<+�a<$�a<�a<�a<��a<�a<Ȥa<��a<��a<��a<c�a<N�a<�a<��a<ԣa<��a<J�a<�a<΢a<��a<z�a<N�a<!�a<�a<ˡa<��a<��a<��a<q�a<0�a<�a<٠a<��a<q�a<8�a<�a<��a<`�a<�a<ߞa<��a<2�a<ٝa<��a<P�a<��a<��a<=�a<ٛa<��a<�a<��a<F�a<ڙa<P�a<�a<x�a<�a<M�a<��a<8�a<��a<F�a<̔a<J�a<֓a<\�a<��a<��a<M�a<ّa<J�a<�a<n�a<��a<��a<�a<}�a<�a<��a<�a<��a< �a<��a<6�a<̊a<q�a<��a<��a<�a<��a<e�a<��a<��a<1�a<φa<c�a<�a<��a<=�a<΄a<w�a<&�a<��a<��a<j�a<,�a<��a<ւa<Ȃa<ǂa<��a<��a<f�a<g�a<E�a<?�a<+�a<�a<��a<��a<�a<��a<�a<�a<�a<��a<�a<*�a<*�a<I�a<X�a<�  �  ;�a<8�a<��a<��a<��a<߁a<�a<�a<�a<Z�a<u�a<��a<܂a<
�a<|�a<��a<$�a<o�a<��a<c�a<��a<Y�a<��a<V�a<��a<B�a<��a<�a<��a<�a<��a<Њa<g�a<ًa<R�a<܌a<_�a<�a<d�a<�a<��a<"�a<��a<�a<ˑa<&�a<ʒa<1�a<��a<�a<f�a<�a<R�a<�a<0�a<֖a<`�a<��a<v�a<ܘa<��a<��a<��a<,�a<��a<H�a<��a<#�a<\�a<�a<=�a<��a<�a<�a<p�a<��a<�a<E�a<��a<Рa<�a<e�a<��a<ϡa<�a<
�a<W�a<`�a<��a<��a<��a<��a<��a<Тa<��a<�a<��a<�a<	�a<&�a<Z�a<n�a<��a<��a<�a<�a<7�a<I�a<O�a<{�a<R�a<�a<n�a<w�a<O�a<J�a<F�a</�a</�a<�a<�a<�a<�a<�a<ߣa<ѣa<��a<��a<j�a<B�a<"�a<עa<��a<A�a<7�a<�a<��a<|�a<7�a<2�a<Πa<ޠa<��a<��a<��a<7�a<O�a<�a<�a<͟a<��a<b�a<*�a<�a<��a<��a<��a<Νa<w�a<"�a<ܜa<��a<>�a<ڛa<��a<I�a<�a<��a<�a<Ιa<5�a<�a<T�a<˗a<5�a<��a<8�a<��a<%�a<h�a<�a<��a<�a<��a< �a<ޑa<J�a<�a<��a<*�a<֏a<6�a<�a<9�a<�a<b�a<݌a<b�a<ċa<Z�a<؊a<l�a<�a<x�a<�a<��a<\�a<�a<��a<�a<��a<W�a<ׅa<��a<�a<��a<�a<̃a<u�a<��a<Ăa<:�a<3�a<فa<��a<��a<`�a<Y�a<�a<'�a<�a<�a<�a<�a<��a<��a<Ҁa<��a<��a<��a<��a<��a<}�a<��a<��a<��a<��a<��a<	�a<�a<�  �  5�a<`�a<��a<��a<��a<ǁa<�a<�a<.�a<D�a<l�a<��a<ׂa<�a<\�a<��a<�a<q�a<ބa<X�a<ۅa<X�a<��a<D�a<��a<E�a<��a<4�a<��a<�a<�a<��a<u�a<ߋa<c�a<ӌa<k�a<�a<��a<�a<��a<�a<��a<?�a<ȑa<9�a<��a<!�a<��a<�a<��a<�a<R�a<֕a<F�a<Öa<I�a<̗a<_�a<ߘa<}�a<�a<��a<)�a<��a<.�a<��a<$�a<��a<�a<-�a<��a<�a<5�a<y�a<��a<��a<H�a<��a<ݠa< �a<U�a<��a<áa<�a<2�a<\�a<m�a<��a<��a<��a<��a<��a<��a<��a<բa<עa<�a<��a<)�a<L�a<k�a<��a<ˣa<�a<�a<#�a<J�a<`�a<w�a<y�a<u�a<`�a<k�a<c�a<Y�a<=�a<:�a<�a<"�a<�a<�a<�a<��a<ԣa<ˣa<��a<��a<t�a<E�a<
�a<Ӣa<��a<l�a<!�a<�a<��a<w�a<5�a<�a<�a<Πa<��a<��a<v�a<g�a<M�a<�a< �a<ٟa<��a<~�a<I�a<��a<��a<l�a<)�a<ܝa<|�a<4�a<Ӝa<��a<>�a<��a<��a<F�a<ٚa<��a<2�a<ʙa<I�a<Ԙa<D�a<Ǘa<L�a<��a<&�a<��a<�a<~�a<��a<��a<�a<��a<"�a<Ǒa<`�a<�a<��a<�a<��a<J�a<�a<g�a<�a<R�a<ߌa<`�a<�a<b�a<�a<`�a<��a<��a<&�a<��a<L�a<�a<|�a<-�a<��a<\�a<�a<{�a<��a<��a<=�a<Ƀa<`�a<��a<��a<T�a<�a<ρa<��a<��a<]�a<F�a<A�a<4�a<�a<�a<�a<��a<�a<ހa<ǀa<��a<��a<��a<��a<�a<��a<z�a<��a<��a<Āa<܀a<��a<�a<�  �  /�a<Z�a<g�a<��a<��a<ԁa<��a<�a<;�a<=�a<��a<��a<�a<)�a<_�a<Ճa<�a<��a<��a<T�a<�a<D�a<چa<I�a<Їa<:�a<��a<#�a<��a<�a<g�a<��a<K�a<��a<`�a<Ȍa<^�a<Ía<u�a<��a<��a<�a<��a<>�a<��a<N�a<��a<<�a<��a<�a<��a<�a<��a<Еa<i�a<Жa<P�a<�a<[�a<�a<��a<�a<��a<$�a<��a<-�a<��a<�a<��a<ޝa<3�a<��a<Ǟa<+�a<M�a<��a<�a<>�a<u�a<��a<�a<>�a<��a<��a<��a<&�a<L�a<�a<��a<��a<��a<��a<��a<ʢa<ߢa<Тa<�a<��a<�a<=�a<L�a<��a<��a<֣a<�a<�a<5�a<O�a<m�a<Z�a<y�a<m�a<v�a<_�a<V�a<G�a<�a<9�a<�a<%�a<�a<��a<��a<�a<�a<ƣa<��a<��a<z�a<O�a<�a<�a<��a<y�a<�a< �a<��a<��a<V�a<�a<�a<͠a<��a<��a<q�a<o�a<:�a<5�a<�a<�a<��a<o�a<8�a<�a<Şa<S�a<"�a<��a<]�a<1�a<Ȝa<��a<�a<�a<��a<E�a<�a<��a<1�a<��a<^�a<јa<_�a<̗a<?�a<��a<'�a<��a<�a<��a<	�a<��a<.�a<��a<S�a<ˑa<c�a<��a<��a<6�a<��a<a�a<ʎa<a�a<ݍa<X�a<�a<E�a<܋a<7�a<׊a<U�a<�a<n�a<��a<��a<5�a<��a<z�a<�a<��a<L�a<��a<}�a<�a<��a<?�a<ȃa<o�a<�a<��a<��a<�a<�a<��a<��a<�a<B�a<L�a<&�a<)�a<�a<�a<�a<׀a<ހa<��a<��a<��a<��a<��a<X�a<��a<p�a<��a<y�a<��a<Հa<�a<�a<�  �  ,�a<K�a<{�a<��a<��a<сa<��a<�a<;�a<W�a<��a<��a<�a<*�a<z�a<ăa<%�a<��a<��a<h�a<��a<[�a<ֆa<@�a<��a<<�a<��a<�a<��a<�a<g�a<؊a<V�a<ʋa<?�a<Ɍa<M�a<ۍa<p�a<��a<z�a<�a<��a<'�a<��a<<�a<��a<3�a<��a<!�a<��a<��a<z�a<�a<]�a<�a<g�a<ߗa<l�a<��a<��a<�a<��a<*�a<��a<!�a<��a<�a<t�a<ޝa<0�a<y�a<ʞa<!�a<b�a<��a<�a<%�a<x�a<��a<��a<=�a<y�a<��a<��a<#�a<T�a<n�a<�a<��a<��a<��a<ɢa<Ѣa<Тa<�a<�a<�a<!�a<=�a<S�a<��a<��a<ӣa<��a<�a<0�a<:�a<\�a<n�a<d�a<k�a<_�a<N�a<G�a<I�a<-�a<�a<�a<�a<��a<��a<�a<գa<ʣa<£a<��a<��a<r�a<<�a<�a<�a<��a<y�a<5�a<��a<��a<��a<W�a<0�a<��a<ߠa<��a<��a<��a<l�a<Q�a<1�a<��a<ןa<��a<u�a<2�a<�a<��a<S�a<�a<��a<h�a<�a<Ȝa<x�a<-�a<�a<��a<,�a<ߚa<��a<�a<��a<L�a<Øa<V�a<˗a<O�a<��a</�a<��a<�a<��a<�a<��a<�a<��a<A�a<ґa<n�a<�a<��a<1�a<��a<J�a<َa<Q�a<ݍa<U�a<Ȍa<H�a<Ӌa<K�a<Ɋa<R�a<Ӊa<q�a<�a<��a<4�a<·a<v�a<�a<��a<U�a<�a<r�a<�a<��a<?�a<ۃa<v�a<�a<��a<k�a<4�a<�a<��a<��a<}�a<Y�a<I�a<<�a<"�a<�a<��a<��a<�a<ɀa<��a<��a<��a<��a<��a<o�a<m�a<w�a<{�a<��a<��a<��a<ڀa<��a<�  �  1�a<?�a<t�a<��a<��a<��a<��a<5�a<1�a<l�a<��a<҂a<�a</�a<��a<Ƀa<_�a<��a<�a<x�a<�a<o�a<͆a<\�a<��a<0�a<��a<�a<��a<܉a<x�a<��a<;�a<��a< �a<��a<"�a<a<3�a<�a<s�a<�a<��a<�a<��a<.�a<Ȓa<A�a<��a<9�a<��a<�a<u�a<�a<u�a<�a<v�a<�a<��a<�a<��a<&�a<��a<?�a<��a<@�a<��a<�a<f�a<ӝa<$�a<k�a<˞a<�a<N�a<~�a<ߟa<�a<X�a<��a<٠a<I�a<c�a<��a<�a<�a<M�a<l�a<��a<��a<Ǣa<âa<Ӣa<�a<�a<#�a<��a</�a<+�a<e�a<��a<��a<��a<Σa<�a<�a<?�a<R�a<N�a<m�a<Y�a<s�a<I�a<P�a<8�a<�a<�a<�a<�a<أa<�a<ңa<ѣa<ޣa<��a<ȣa<��a<��a<c�a<K�a<#�a<�a<΢a<o�a<I�a<�a<�a<��a<]�a<Q�a<�a<�a<ՠa<��a<��a<m�a<d�a<(�a<�a<ٟa<��a<l�a<+�a<��a<��a<d�a<�a<��a<K�a<�a<��a<M�a<�a<��a<��a<$�a<Қa<��a<�a<��a<>�a<�a<d�a<ۗa<g�a<ʖa<O�a<��a<R�a<��a<'�a<��a<-�a<�a<H�a<�a<x�a<�a<��a<8�a<Ώa<@�a<֎a<C�a<Ӎa<I�a<��a<J�a<��a<7�a<��a<G�a<��a<Q�a<��a<w�a<@�a<��a<u�a<�a<��a<M�a<�a<��a<�a<��a<F�a<�a<��a<)�a<��a<s�a<S�a<��a<�a<��a<|�a<q�a<E�a<U�a<#�a<"�a<�a<�a<�a<��a<ŀa<��a<��a<q�a<Q�a<W�a<@�a<r�a<O�a<t�a<��a<��a<�a<�a<�  �  �a<3�a<k�a<��a<��a<��a<�a<%�a<L�a<��a<��a<ɂa<�a<T�a<��a<�a<C�a<��a<)�a<��a<��a<g�a<�a<Y�a<Ça<8�a<��a<��a<}�a<�a<B�a<��a<*�a<��a<�a<��a<�a<��a<3�a<Ɏa<]�a< �a<��a<#�a<��a<=�a<��a<F�a<��a<1�a<��a<=�a<��a<�a<��a<�a<��a<�a<��a<�a<ƙa<8�a<��a<B�a<Ǜa<6�a<��a<�a<s�a<��a<�a<^�a<��a<�a<<�a<w�a<��a<�a<M�a<��a<Ѡa<�a<m�a<��a<Сa<�a<O�a<p�a<��a<��a<��a<ۢa<�a<�a<�a<�a< �a<G�a<K�a<f�a<w�a<��a<�a<�a<�a<1�a<B�a<N�a<]�a<`�a<S�a<R�a<K�a<+�a<$�a<�a<�a<�a<�a<ףa<ݣa<ˣa<��a<��a<��a<��a<��a<��a<q�a<K�a<#�a<��a<��a<��a<k�a<)�a<ءa<��a<��a<g�a<-�a<��a<Ѡa<ՠa<��a<��a<]�a<C�a<�a<ܟa<��a<m�a<�a<ޞa<��a<.�a<۝a<��a<B�a<�a<��a<H�a<
�a<��a<^�a<�a<˚a<d�a<�a<��a<L�a<֘a<i�a<�a<_�a<ߖa<q�a<��a<;�a<Ŕa<D�a<ϓa<S�a<̒a<[�a<�a<��a<�a<��a<B�a<ďa<O�a<Ўa<P�a<��a<A�a<��a<#�a<��a<&�a<��a< �a<��a<F�a<߈a<n�a<�a<a<f�a<�a<��a<O�a<�a<��a<+�a<��a<]�a<��a<��a<,�a<܂a<��a<k�a<�a<�a<��a<��a<��a<`�a<F�a<@�a<%�a<
�a<��a<݀a<��a<��a<��a<g�a<^�a<P�a<Q�a<=�a<A�a<N�a<p�a<�a<��a<��a<�a<�  �  ��a<A�a<`�a<��a<��a<�a<�a<&�a<q�a<{�a<Ăa<�a<3�a<u�a<��a<�a<d�a<ʄa<1�a<��a<�a<h�a<��a<N�a<Ňa<(�a<��a<�a<[�a<ىa<%�a<��a<�a<��a<�a<n�a<�a<��a<)�a<��a<I�a<��a<v�a<+�a<��a<8�a<��a<U�a<Ǔa<D�a<Ĕa<$�a<��a<'�a<��a<�a<��a<@�a<��a<=�a<��a<J�a<ؚa<G�a<ڛa<(�a<��a<��a<w�a<��a<�a<L�a<��a<۞a<�a<s�a<��a<�a<A�a<x�a<Ƞa<��a<[�a<��a<ܡa<�a<:�a<r�a<��a<ɢa<âa<��a<�a<�a<�a<"�a<J�a<<�a<k�a<��a<��a<ţa<ͣa<
�a<	�a<9�a<J�a<J�a<V�a<O�a<^�a<6�a<H�a<�a<�a<��a<�a<�a<��a<ƣa<��a<��a<��a<��a<��a<��a<��a<~�a<f�a<G�a<)�a<
�a<��a<��a<X�a<<�a<��a<ӡa<��a<X�a<U�a<�a<��a<ܠa<��a<��a<^�a<Q�a<
�a<ݟa<��a<h�a<�a<��a<��a<�a<ҝa<u�a</�a<Ҝa<n�a<C�a<ݛa<��a<I�a<��a<Ța<V�a<�a<��a<H�a<Ϙa<x�a<�a<r�a<��a<X�a<�a<]�a<�a<V�a<Փa<|�a<�a<��a< �a<��a<6�a<��a<U�a<��a<I�a<��a<T�a<��a<:�a<��a<	�a<��a<��a<��a<��a<��a<:�a<��a<e�a<�a<��a<L�a<��a<��a<:�a<�a<}�a<<�a<��a<}�a<��a<��a<[�a<��a<ǂa<`�a<;�a<�a<Ձa<��a<~�a<��a<I�a<H�a<-�a<�a<��a<̀a<Àa<��a<��a<P�a<L�a<7�a<*�a<2�a<�a<=�a<N�a<b�a<��a<��a<�a<�  �  �a<1�a<]�a<��a<Áa<�a<�a<H�a<x�a<��a<ςa<�a<S�a<��a<уa<%�a<��a<�a<B�a<��a<�a<��a<�a<a�a<ʇa<.�a<��a<�a<S�a<��a<=�a<��a<�a<h�a<�a<u�a<�a<l�a<��a<��a<?�a<ޏa<q�a<�a<��a<6�a<̒a<T�a<��a<X�a<Քa<C�a<��a<H�a<��a<>�a<��a<E�a<Әa<G�a<әa<\�a<�a<J�a<כa<D�a<��a<�a<d�a<��a<��a<;�a<��a<��a<��a<H�a<��a<Οa<�a<T�a<��a<�a<D�a<��a<֡a<�a<A�a<w�a<��a<��a<עa<��a<�a<�a<*�a<O�a<R�a<d�a<��a<��a<��a<ͣa<�a<�a<-�a<*�a<P�a<Z�a<V�a<V�a<P�a<4�a<&�a<�a<	�a<Уa<ȣa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<z�a<h�a<T�a<2�a<��a<�a<��a<s�a<G�a<�a<�a<��a<��a<`�a<I�a<�a<�a<��a<��a<y�a<G�a<�a<�a<��a<_�a<�a<��a<d�a<*�a<��a<O�a<�a<��a<t�a<�a<��a<t�a<M�a<�a<��a<Q�a<�a<��a<F�a<�a<w�a<�a<��a<�a<w�a<�a<�a<��a<v�a<��a<��a<�a<��a<�a<��a<A�a<��a<R�a<ҏa<L�a<Ďa<B�a<��a<�a<��a<�a<f�a<ߊa<o�a<��a<|�a<�a<��a<>�a<�a<��a<=�a<��a<��a<A�a<�a<��a<4�a<τa<��a<�a<��a<g�a<*�a<ςa<��a<S�a<'�a<�a<��a<��a<��a<n�a<9�a<2�a<�a<��a<Ҁa<��a<��a<k�a<[�a<C�a<�a<
�a<�a< �a<�a<,�a<;�a<|�a<��a<Āa<�  �  �a<�a<^�a<��a<��a<��a<�a<d�a<o�a<ǂa<��a<�a<X�a<��a<��a<'�a<��a<߄a<X�a<ąa<�a<��a<��a<n�a<��a<5�a<��a<�a<b�a<��a<�a<i�a<��a<a�a<ċa<\�a<a<��a<��a<��a<,�a<ʏa<v�a<�a<��a</�a<˒a<I�a<ޓa<d�a<ϔa<r�a<Õa<X�a<̖a<T�a<ߗa<N�a<�a<K�a<��a<b�a<�a<g�a<ɛa<H�a<��a<�a<V�a<��a<�a<+�a<z�a<��a<�a< �a<v�a<��a<�a<h�a<��a<�a<.�a<��a<��a<�a<M�a<h�a<��a<��a<��a<�a<�a<5�a<'�a<X�a<U�a<��a<��a<��a<ɣa<ߣa<!�a<�a<E�a<B�a<R�a<O�a<S�a<Y�a<5�a<>�a<�a<�a<�a<գa<ܣa<��a<��a<}�a<��a<��a<}�a<��a<t�a<��a<r�a<|�a<g�a<H�a<9�a<�a<��a<��a<��a<Y�a<$�a<��a<��a<��a<a�a<O�a<�a<�a<�a<��a<��a<K�a<*�a<ԟa<��a<[�a<��a<Þa<K�a<�a<��a<^�a<��a<��a<[�a<�a<��a<k�a<4�a<ޚa<��a<V�a<��a<��a<?�a<�a<l�a<�a<��a<�a<��a<��a<��a<�a<��a<�a<��a<$�a<��a<F�a<��a<I�a<Ґa<D�a<׏a<?�a<͎a<4�a<��a<�a<{�a<��a<W�a<��a<F�a<މa<_�a<��a<��a<'�a<�a<��a<H�a<�a<��a<M�a<߅a<��a<.�a<��a<��a<.�a<ڃa<e�a<3�a<҂a<��a<W�a<.�a< �a<сa<Ӂa<��a<��a<Q�a<5�a<�a<�a<րa<��a<��a<O�a<>�a<"�a<�a<�a<�a<
�a<�a<4�a<B�a<W�a<��a<��a<�  �  �a<�a<N�a<��a<Ła<��a<%�a<]�a<��a<��a<��a<=�a<n�a<��a<�a<T�a<��a<�a<f�a<Ņa<2�a<��a<��a<m�a<ɇa<�a<��a<�a<I�a<��a<��a<o�a<Ċa<?�a<��a<?�a<��a<N�a<ݍa<��a<#�a<��a<d�a<�a<��a<5�a<ђa<W�a<�a<j�a<�a<h�a<�a<o�a<�a<b�a<�a<p�a<��a<��a<��a<r�a<��a<t�a<؛a<K�a<��a<�a<S�a<��a<ݝa<!�a<[�a<��a<Ԟa<�a<c�a<��a<�a</�a<��a<Ѡa<%�a<w�a<��a<��a<-�a<u�a<��a<Ȣa<��a<�a<!�a<>�a<e�a<q�a<��a<��a<��a<ǣa<�a<��a<�a<"�a<>�a<I�a<[�a<]�a<N�a<B�a<>�a<+�a<�a<�a<أa<��a<��a<��a<��a<x�a<s�a<i�a<s�a<t�a<~�a<��a<y�a<k�a<[�a<V�a<A�a<�a<��a<Ţa<��a<n�a<K�a<�a<�a<��a<��a<g�a<K�a<�a<�a<��a<��a<V�a<)�a<�a<��a<K�a<��a<��a<K�a<�a<��a<+�a<ܜa<��a<?�a<�a<��a<S�a<�a<՚a<��a<D�a<��a<��a<E�a<�a<z�a<�a<��a<�a<��a<#�a<��a<%�a<��a<$�a<��a<7�a<Ēa<A�a<őa<T�a<ߐa<S�a<ُa<H�a<��a<0�a<��a<�a<p�a<ًa<J�a<��a<7�a<ˉa<V�a<�a<x�a<-�a<ȇa<z�a<0�a<Նa<��a<-�a<�a<��a<;�a<�a<��a<2�a<�a<��a<L�a<��a<��a<z�a<H�a< �a<�a<��a<��a<~�a<Y�a<>�a<�a<�a<��a<��a<}�a<T�a<-�a<�a<�a<�a<�a<�a<�a<�a<�a<L�a<x�a<��a<�  �  рa< �a<Q�a<��a<ˁa<�a<3�a<a�a<��a<Âa<�a<5�a<_�a<؃a<�a<l�a<��a<�a<q�a<ׅa<C�a<��a<�a<Z�a<ۇa<-�a<��a<�a<5�a<��a<�a<q�a<��a<A�a<��a<&�a<Ќa<<�a<�a<y�a<�a<��a<R�a<�a<��a<F�a<ǒa<\�a<�a<m�a<�a<g�a<�a<^�a<�a<v�a<�a<z�a<�a<��a<��a<��a<��a<s�a<�a<>�a<��a<��a<W�a<��a<՝a<�a<S�a<��a<Ğa<'�a<K�a<��a<�a<�a<��a<Ša<&�a<f�a<��a<�a<>�a<��a<��a<ߢa<��a<�a<8�a<A�a<g�a<W�a<��a<��a<Σa<��a<ݣa<�a<�a<J�a<B�a<S�a<Q�a<]�a<`�a<H�a<A�a<�a<�a<ڣa<ףa<��a<��a<��a<m�a<|�a<i�a<m�a<w�a<Z�a<~�a<g�a<}�a<o�a<p�a<[�a<0�a<$�a<��a<�a<��a<��a<D�a< �a<�a<��a<��a<O�a<K�a<�a<��a<Рa<��a<k�a<�a<�a<��a<Q�a<��a<��a<N�a<՝a<��a<�a<ޜa<}�a<&�a<��a<��a<c�a<�a<Ěa<��a<2�a<��a<��a<V�a<�a<�a<�a<��a<@�a<��a<<�a<��a<&�a<��a<-�a<��a<$�a<Ԓa<>�a<�a<X�a<ސa<_�a<̏a<_�a<��a<4�a<��a<��a<c�a<ыa<\�a<��a<M�a<��a<C�a<�a<g�a<3�a<��a<{�a<�a<؆a<��a<>�a<��a<��a<R�a<�a<��a<I�a<�a<��a<2�a<�a<��a<��a<;�a<�a<�a<Áa<��a<��a<b�a<3�a<�a<��a<ŀa<��a<c�a<U�a<�a<�a<�a<�a<�a<�a<�a<�a<!�a<Q�a<_�a<��a<�  �  �a<�a<G�a<��a<ȁa<�a<<�a<f�a<��a<ڂa<�a<R�a<��a<Ճa<�a<p�a<��a<&�a<��a<�a</�a<��a<�a<w�a<͇a<+�a<x�a<ֈa<C�a<��a<�a<K�a<��a<*�a<��a<!�a<��a<A�a<ʍa<n�a<�a<��a<a�a<�a<��a<2�a<ےa<g�a<��a<m�a<��a<�a<�a<��a<�a<��a<��a<��a<�a<��a<�a<��a<��a<��a<�a<V�a<��a<��a<8�a<��a<ߝa<�a<L�a<|�a<Ȟa<��a<E�a<��a<ҟa<&�a<h�a<Ǡa< �a<r�a<��a<�a<@�a<t�a<��a<ߢa<�a<�a<=�a<Z�a<t�a<�a<��a<��a<ͣa<ۣa<�a<�a<*�a<1�a<H�a<c�a<c�a<d�a<R�a<B�a<$�a<%�a<�a<�a<��a<��a<��a<q�a<j�a<X�a<`�a<X�a<\�a<a�a<q�a<y�a<d�a<d�a<c�a<Y�a<I�a<-�a< �a<Тa<��a<��a<`�a<$�a<�a<��a<��a<v�a<[�a</�a<��a<��a<��a<j�a<3�a<�a<��a<>�a<�a<��a<E�a<ٝa<v�a<"�a<ǜa<g�a<!�a<Λa<��a<?�a<�a<Ěa<��a<B�a<ޙa<��a<B�a<��a<��a<#�a<��a<*�a<��a<C�a<Õa<9�a<��a<8�a<Ǔa<R�a<ܒa<X�a<ܑa<T�a<�a<g�a<�a<G�a<��a<�a<��a<�a<`�a<ˋa<.�a<��a<#�a<��a<2�a<ˈa<n�a<�a<��a<u�a<+�a<Άa<}�a<@�a<�a<��a<Q�a<��a<��a<N�a<��a<��a<Z�a<�a<Ƃa<��a<\�a<:�a<�a<܁a<��a<��a<r�a<F�a< �a<�a<��a<��a<w�a<L�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<6�a<f�a<��a<�  �  ��a<�a<^�a<��a<��a<��a<�a<m�a<��a<�a<�a<G�a<��a<Ãa<�a<e�a<Ąa<�a<r�a<�a<?�a<��a<�a<{�a<��a<*�a<��a<؈a<1�a<r�a<��a<N�a<ϊa<"�a<��a<=�a<��a<U�a<ča<��a<�a<��a<d�a<�a<��a<&�a<Ւa<;�a<�a<z�a<��a<��a<�a<��a<��a<��a<�a<|�a<	�a<q�a<�a<��a<�a<t�a<��a<S�a<��a<�a<H�a<��a<��a<��a<e�a<y�a<ݞa<��a<_�a<��a<��a<<�a<g�a<٠a<��a<]�a<��a<��a<I�a<a�a<��a<��a<�a<�a<B�a<Q�a<Y�a<��a<��a<��a<��a<ڣa<��a<�a<>�a<:�a<R�a<A�a<N�a<a�a<I�a<U�a<&�a<'�a<٣a<�a<ͣa<��a<��a<a�a<��a<T�a<j�a<[�a<h�a<w�a<G�a<v�a<h�a<{�a<^�a<R�a<C�a<�a<�a<ۢa<ʢa<i�a<V�a<)�a<�a<ԡa<��a<~�a<H�a<�a<�a<ˠa<��a<@�a<7�a<џa<��a<O�a<�a<��a<�a<�a<y�a<5�a<��a<u�a<=�a<��a<��a<:�a<�a<��a<`�a<D�a<�a<��a<6�a<�a<^�a<�a<��a<)�a<��a<�a<��a<+�a<��a<E�a<��a<H�a<��a<]�a<ّa<b�a<ߐa<9�a<�a<5�a<Վa<%�a<��a<��a<O�a<�a<+�a<Ǌa<�a<Ɖa<D�a<��a<��a<�a<Їa<O�a<�a<цa<��a<I�a<؅a<��a<&�a< �a<��a<S�a<��a<��a<]�a<�a<тa<��a<[�a<-�a<�a<��a<��a<��a<P�a<1�a<�a<�a<Ҁa<��a<y�a<�a<+�a<�a<�a<�a<�a<�a<�a<�a<�a<A�a<|�a<{�a<�  �  �a<�a<G�a<��a<ȁa<�a<<�a<f�a<��a<ڂa<�a<R�a<��a<Ճa<�a<p�a<��a<&�a<��a<�a</�a<��a<�a<w�a<͇a<+�a<x�a<ֈa<C�a<��a<�a<K�a<��a<*�a<��a<!�a<��a<A�a<ʍa<n�a<�a<��a<a�a<�a<��a<2�a<ےa<g�a<��a<m�a<��a<�a<�a<��a<�a<��a<��a<��a<�a<��a<�a<��a<��a<��a<�a<V�a<��a<��a<8�a<��a<ߝa<�a<L�a<|�a<Ȟa<��a<E�a<��a<ҟa<&�a<h�a<Ǡa< �a<r�a<��a<�a<@�a<t�a<��a<ߢa<�a<�a<=�a<Z�a<t�a<�a<��a<��a<ͣa<ۣa<�a<�a<*�a<1�a<H�a<c�a<c�a<d�a<R�a<B�a<$�a<%�a<�a<�a<��a<��a<��a<q�a<j�a<X�a<`�a<X�a<\�a<a�a<q�a<y�a<d�a<d�a<c�a<Y�a<I�a<-�a< �a<Тa<��a<��a<`�a<$�a<�a<��a<��a<v�a<[�a</�a<��a<��a<��a<j�a<3�a<�a<��a<>�a<�a<��a<E�a<ٝa<v�a<"�a<ǜa<g�a<!�a<Λa<��a<?�a<�a<Ěa<��a<B�a<ޙa<��a<B�a<��a<��a<#�a<��a<*�a<��a<C�a<Õa<9�a<��a<8�a<Ǔa<R�a<ܒa<X�a<ܑa<T�a<�a<g�a<�a<G�a<��a<�a<��a<�a<`�a<ˋa<.�a<��a<#�a<��a<2�a<ˈa<n�a<�a<��a<u�a<+�a<Άa<}�a<@�a<�a<��a<Q�a<��a<��a<N�a<��a<��a<Z�a<�a<Ƃa<��a<\�a<:�a<�a<܁a<��a<��a<r�a<F�a< �a<�a<��a<��a<w�a<L�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<6�a<f�a<��a<�  �  рa< �a<Q�a<��a<ˁa<�a<3�a<a�a<��a<Âa<�a<5�a<_�a<؃a<�a<l�a<��a<�a<q�a<ׅa<C�a<��a<�a<Z�a<ۇa<-�a<��a<�a<5�a<��a<�a<q�a<��a<A�a<��a<&�a<Ќa<<�a<�a<y�a<�a<��a<R�a<�a<��a<F�a<ǒa<\�a<�a<m�a<�a<g�a<�a<^�a<�a<v�a<�a<z�a<�a<��a<��a<��a<��a<s�a<�a<>�a<��a<��a<W�a<��a<՝a<�a<S�a<��a<Ğa<'�a<K�a<��a<�a<�a<��a<Ša<&�a<f�a<��a<�a<>�a<��a<��a<ߢa<��a<�a<8�a<A�a<g�a<W�a<��a<��a<Σa<��a<ݣa<�a<�a<J�a<B�a<S�a<Q�a<]�a<`�a<H�a<A�a<�a<�a<ڣa<ףa<��a<��a<��a<m�a<|�a<i�a<m�a<w�a<Z�a<~�a<g�a<}�a<o�a<p�a<[�a<0�a<$�a<��a<�a<��a<��a<D�a< �a<�a<��a<��a<O�a<K�a<�a<��a<Рa<��a<k�a<�a<�a<��a<Q�a<��a<��a<N�a<՝a<��a<�a<ޜa<}�a<&�a<��a<��a<c�a<�a<Ěa<��a<2�a<��a<��a<V�a<�a<�a<�a<��a<@�a<��a<<�a<��a<&�a<��a<-�a<��a<$�a<Ԓa<>�a<�a<X�a<ސa<_�a<̏a<_�a<��a<4�a<��a<��a<c�a<ыa<\�a<��a<M�a<��a<C�a<�a<g�a<3�a<��a<{�a<�a<؆a<��a<>�a<��a<��a<R�a<�a<��a<I�a<�a<��a<2�a<�a<��a<��a<;�a<�a<�a<Áa<��a<��a<b�a<3�a<�a<��a<ŀa<��a<c�a<U�a<�a<�a<�a<�a<�a<�a<�a<�a<!�a<Q�a<_�a<��a<�  �  �a<�a<N�a<��a<Ła<��a<%�a<]�a<��a<��a<��a<=�a<n�a<��a<�a<T�a<��a<�a<f�a<Ņa<2�a<��a<��a<m�a<ɇa<�a<��a<�a<I�a<��a<��a<o�a<Ċa<?�a<��a<?�a<��a<N�a<ݍa<��a<#�a<��a<d�a<�a<��a<5�a<ђa<W�a<�a<j�a<�a<h�a<�a<o�a<�a<b�a<�a<p�a<��a<��a<��a<r�a<��a<t�a<؛a<K�a<��a<�a<S�a<��a<ݝa<!�a<[�a<��a<Ԟa<�a<c�a<��a<�a</�a<��a<Ѡa<%�a<w�a<��a<��a<-�a<u�a<��a<Ȣa<��a<�a<!�a<>�a<e�a<q�a<��a<��a<��a<ǣa<�a<��a<�a<"�a<>�a<I�a<[�a<]�a<N�a<B�a<>�a<+�a<�a<�a<أa<��a<��a<��a<��a<x�a<s�a<i�a<s�a<t�a<~�a<��a<y�a<k�a<[�a<V�a<A�a<�a<��a<Ţa<��a<n�a<K�a<�a<�a<��a<��a<g�a<K�a<�a<�a<��a<��a<V�a<)�a<�a<��a<K�a<��a<��a<K�a<�a<��a<+�a<ܜa<��a<?�a<�a<��a<S�a<�a<՚a<��a<D�a<��a<��a<E�a<�a<z�a<�a<��a<�a<��a<#�a<��a<%�a<��a<$�a<��a<7�a<Ēa<A�a<őa<T�a<ߐa<S�a<ُa<H�a<��a<0�a<��a<�a<p�a<ًa<J�a<��a<7�a<ˉa<V�a<�a<x�a<-�a<ȇa<z�a<0�a<Նa<��a<-�a<�a<��a<;�a<�a<��a<2�a<�a<��a<L�a<��a<��a<z�a<H�a< �a<�a<��a<��a<~�a<Y�a<>�a<�a<�a<��a<��a<}�a<T�a<-�a<�a<�a<�a<�a<�a<�a<�a<�a<L�a<x�a<��a<�  �  �a<�a<^�a<��a<��a<��a<�a<d�a<o�a<ǂa<��a<�a<X�a<��a<��a<'�a<��a<߄a<X�a<ąa<�a<��a<��a<n�a<��a<5�a<��a<�a<b�a<��a<�a<i�a<��a<a�a<ċa<\�a<a<��a<��a<��a<,�a<ʏa<v�a<�a<��a</�a<˒a<I�a<ޓa<d�a<ϔa<r�a<Õa<X�a<̖a<T�a<ߗa<N�a<�a<K�a<��a<b�a<�a<g�a<ɛa<H�a<��a<�a<V�a<��a<�a<+�a<z�a<��a<�a< �a<v�a<��a<�a<h�a<��a<�a<.�a<��a<��a<�a<M�a<h�a<��a<��a<��a<�a<�a<5�a<'�a<X�a<U�a<��a<��a<��a<ɣa<ߣa<!�a<�a<E�a<B�a<R�a<O�a<S�a<Y�a<5�a<>�a<�a<�a<�a<գa<ܣa<��a<��a<}�a<��a<��a<}�a<��a<t�a<��a<r�a<|�a<g�a<H�a<9�a<�a<��a<��a<��a<Y�a<$�a<��a<��a<��a<a�a<O�a<�a<�a<�a<��a<��a<K�a<*�a<ԟa<��a<[�a<��a<Þa<K�a<�a<��a<^�a<��a<��a<[�a<�a<��a<k�a<4�a<ޚa<��a<V�a<��a<��a<?�a<�a<l�a<�a<��a<�a<��a<��a<��a<�a<��a<�a<��a<$�a<��a<F�a<��a<I�a<Ґa<D�a<׏a<?�a<͎a<4�a<��a<�a<{�a<��a<W�a<��a<F�a<މa<_�a<��a<��a<'�a<�a<��a<H�a<�a<��a<M�a<߅a<��a<.�a<��a<��a<.�a<ڃa<e�a<3�a<҂a<��a<W�a<.�a< �a<сa<Ӂa<��a<��a<Q�a<5�a<�a<�a<րa<��a<��a<O�a<>�a<"�a<�a<�a<�a<
�a<�a<4�a<B�a<W�a<��a<��a<�  �  �a<1�a<]�a<��a<Áa<�a<�a<H�a<x�a<��a<ςa<�a<S�a<��a<уa<%�a<��a<�a<B�a<��a<�a<��a<�a<a�a<ʇa<.�a<��a<�a<S�a<��a<=�a<��a<�a<h�a<�a<u�a<�a<l�a<��a<��a<?�a<ޏa<q�a<�a<��a<6�a<̒a<T�a<��a<X�a<Քa<C�a<��a<H�a<��a<>�a<��a<E�a<Әa<G�a<әa<\�a<�a<J�a<כa<D�a<��a<�a<d�a<��a<��a<;�a<��a<��a<��a<H�a<��a<Οa<�a<T�a<��a<�a<D�a<��a<֡a<�a<A�a<w�a<��a<��a<עa<��a<�a<�a<*�a<O�a<R�a<d�a<��a<��a<��a<ͣa<�a<�a<-�a<*�a<P�a<Z�a<V�a<V�a<P�a<4�a<&�a<�a<	�a<Уa<ȣa<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<z�a<h�a<T�a<2�a<��a<�a<��a<s�a<G�a<�a<�a<��a<��a<`�a<I�a<�a<�a<��a<��a<y�a<G�a<�a<�a<��a<_�a<�a<��a<d�a<*�a<��a<O�a<�a<��a<t�a<�a<��a<t�a<M�a<�a<��a<Q�a<�a<��a<F�a<�a<w�a<�a<��a<�a<w�a<�a<�a<��a<v�a<��a<��a<�a<��a<�a<��a<A�a<��a<R�a<ҏa<L�a<Ďa<B�a<��a<�a<��a<�a<f�a<ߊa<o�a<��a<|�a<�a<��a<>�a<�a<��a<=�a<��a<��a<A�a<�a<��a<4�a<τa<��a<�a<��a<g�a<*�a<ςa<��a<S�a<'�a<�a<��a<��a<��a<n�a<9�a<2�a<�a<��a<Ҁa<��a<��a<k�a<[�a<C�a<�a<
�a<�a< �a<�a<,�a<;�a<|�a<��a<Āa<�  �  ��a<A�a<`�a<��a<��a<�a<�a<&�a<q�a<{�a<Ăa<�a<3�a<u�a<��a<�a<d�a<ʄa<1�a<��a<�a<h�a<��a<N�a<Ňa<(�a<��a<�a<[�a<ىa<%�a<��a<�a<��a<�a<n�a<�a<��a<)�a<��a<I�a<��a<v�a<+�a<��a<8�a<��a<U�a<Ǔa<D�a<Ĕa<$�a<��a<'�a<��a<�a<��a<@�a<��a<=�a<��a<J�a<ؚa<G�a<ڛa<(�a<��a<��a<w�a<��a<�a<L�a<��a<۞a<�a<s�a<��a<�a<A�a<x�a<Ƞa<��a<[�a<��a<ܡa<�a<:�a<r�a<��a<ɢa<âa<��a<�a<�a<�a<"�a<J�a<<�a<k�a<��a<��a<ţa<ͣa<
�a<	�a<9�a<J�a<J�a<V�a<O�a<^�a<6�a<H�a<�a<�a<��a<�a<�a<��a<ƣa<��a<��a<��a<��a<��a<��a<��a<~�a<f�a<G�a<)�a<
�a<��a<��a<X�a<<�a<��a<ӡa<��a<X�a<U�a<�a<��a<ܠa<��a<��a<^�a<Q�a<
�a<ݟa<��a<h�a<�a<��a<��a<�a<ҝa<u�a</�a<Ҝa<n�a<C�a<ݛa<��a<I�a<��a<Ța<V�a<�a<��a<H�a<Ϙa<x�a<�a<r�a<��a<X�a<�a<]�a<�a<V�a<Փa<|�a<�a<��a< �a<��a<6�a<��a<U�a<��a<I�a<��a<T�a<��a<:�a<��a<	�a<��a<��a<��a<��a<��a<:�a<��a<e�a<�a<��a<L�a<��a<��a<:�a<�a<}�a<<�a<��a<}�a<��a<��a<[�a<��a<ǂa<`�a<;�a<�a<Ձa<��a<~�a<��a<I�a<H�a<-�a<�a<��a<̀a<Àa<��a<��a<P�a<L�a<7�a<*�a<2�a<�a<=�a<N�a<b�a<��a<��a<�a<�  �  �a<3�a<k�a<��a<��a<��a<�a<%�a<L�a<��a<��a<ɂa<�a<T�a<��a<�a<C�a<��a<)�a<��a<��a<g�a<�a<Y�a<Ça<8�a<��a<��a<}�a<�a<B�a<��a<*�a<��a<�a<��a<�a<��a<3�a<Ɏa<]�a< �a<��a<#�a<��a<=�a<��a<F�a<��a<1�a<��a<=�a<��a<�a<��a<�a<��a<�a<��a<�a<ƙa<8�a<��a<B�a<Ǜa<6�a<��a<�a<s�a<��a<�a<^�a<��a<�a<<�a<w�a<��a<�a<M�a<��a<Ѡa<�a<m�a<��a<Сa<�a<O�a<p�a<��a<��a<��a<ۢa<�a<�a<�a<�a< �a<G�a<K�a<f�a<w�a<��a<�a<�a<�a<1�a<B�a<N�a<]�a<`�a<S�a<R�a<K�a<+�a<$�a<�a<�a<�a<�a<ףa<ݣa<ˣa<��a<��a<��a<��a<��a<��a<q�a<K�a<#�a<��a<��a<��a<k�a<)�a<ءa<��a<��a<g�a<-�a<��a<Ѡa<ՠa<��a<��a<]�a<C�a<�a<ܟa<��a<m�a<�a<ޞa<��a<.�a<۝a<��a<B�a<�a<��a<H�a<
�a<��a<^�a<�a<˚a<d�a<�a<��a<L�a<֘a<i�a<�a<_�a<ߖa<q�a<��a<;�a<Ŕa<D�a<ϓa<S�a<̒a<[�a<�a<��a<�a<��a<B�a<ďa<O�a<Ўa<P�a<��a<A�a<��a<#�a<��a<&�a<��a< �a<��a<F�a<߈a<n�a<�a<a<f�a<�a<��a<O�a<�a<��a<+�a<��a<]�a<��a<��a<,�a<܂a<��a<k�a<�a<�a<��a<��a<��a<`�a<F�a<@�a<%�a<
�a<��a<݀a<��a<��a<��a<g�a<^�a<P�a<Q�a<=�a<A�a<N�a<p�a<�a<��a<��a<�a<�  �  1�a<?�a<t�a<��a<��a<��a<��a<5�a<1�a<l�a<��a<҂a<�a</�a<��a<Ƀa<_�a<��a<�a<x�a<�a<o�a<͆a<\�a<��a<0�a<��a<�a<��a<܉a<x�a<��a<;�a<��a< �a<��a<"�a<a<3�a<�a<s�a<�a<��a<�a<��a<.�a<Ȓa<A�a<��a<9�a<��a<�a<u�a<�a<u�a<�a<v�a<�a<��a<�a<��a<&�a<��a<?�a<��a<@�a<��a<�a<f�a<ӝa<$�a<k�a<˞a<�a<N�a<~�a<ߟa<�a<X�a<��a<٠a<I�a<c�a<��a<�a<�a<M�a<l�a<��a<��a<Ǣa<âa<Ӣa<�a<�a<#�a<��a</�a<+�a<e�a<��a<��a<��a<Σa<�a<�a<?�a<R�a<N�a<m�a<Y�a<s�a<I�a<P�a<8�a<�a<�a<�a<�a<أa<�a<ңa<ѣa<ޣa<��a<ȣa<��a<��a<c�a<K�a<#�a<�a<΢a<o�a<I�a<�a<�a<��a<]�a<Q�a<�a<�a<ՠa<��a<��a<m�a<d�a<(�a<�a<ٟa<��a<l�a<+�a<��a<��a<d�a<�a<��a<K�a<�a<��a<M�a<�a<��a<��a<$�a<Қa<��a<�a<��a<>�a<�a<d�a<ۗa<g�a<ʖa<O�a<��a<R�a<��a<'�a<��a<-�a<�a<H�a<�a<x�a<�a<��a<8�a<Ώa<@�a<֎a<C�a<Ӎa<I�a<��a<J�a<��a<7�a<��a<G�a<��a<Q�a<��a<w�a<@�a<��a<u�a<�a<��a<M�a<�a<��a<�a<��a<F�a<�a<��a<)�a<��a<s�a<S�a<��a<�a<��a<|�a<q�a<E�a<U�a<#�a<"�a<�a<�a<�a<��a<ŀa<��a<��a<q�a<Q�a<W�a<@�a<r�a<O�a<t�a<��a<��a<�a<�a<�  �  ,�a<K�a<{�a<��a<��a<сa<��a<�a<;�a<W�a<��a<��a<�a<*�a<z�a<ăa<%�a<��a<��a<h�a<��a<[�a<ֆa<@�a<��a<<�a<��a<�a<��a<�a<g�a<؊a<V�a<ʋa<?�a<Ɍa<M�a<ۍa<p�a<��a<z�a<�a<��a<'�a<��a<<�a<��a<3�a<��a<!�a<��a<��a<z�a<�a<]�a<�a<g�a<ߗa<l�a<��a<��a<�a<��a<*�a<��a<!�a<��a<�a<t�a<ޝa<0�a<y�a<ʞa<!�a<b�a<��a<�a<%�a<x�a<��a<��a<=�a<y�a<��a<��a<#�a<T�a<n�a<�a<��a<��a<��a<ɢa<Ѣa<Тa<�a<�a<�a<!�a<=�a<S�a<��a<��a<ӣa<��a<�a<0�a<:�a<\�a<n�a<d�a<k�a<_�a<N�a<G�a<I�a<-�a<�a<�a<�a<��a<��a<�a<գa<ʣa<£a<��a<��a<r�a<<�a<�a<�a<��a<y�a<5�a<��a<��a<��a<W�a<0�a<��a<ߠa<��a<��a<��a<l�a<Q�a<1�a<��a<ןa<��a<u�a<2�a<�a<��a<S�a<�a<��a<h�a<�a<Ȝa<x�a<-�a<�a<��a<,�a<ߚa<��a<�a<��a<L�a<Øa<V�a<˗a<O�a<��a</�a<��a<�a<��a<�a<��a<�a<��a<A�a<ґa<n�a<�a<��a<1�a<��a<J�a<َa<Q�a<ݍa<U�a<Ȍa<H�a<Ӌa<K�a<Ɋa<R�a<Ӊa<q�a<�a<��a<4�a<·a<v�a<�a<��a<U�a<�a<r�a<�a<��a<?�a<ۃa<v�a<�a<��a<k�a<4�a<�a<��a<��a<}�a<Y�a<I�a<<�a<"�a<�a<��a<��a<�a<ɀa<��a<��a<��a<��a<��a<o�a<m�a<w�a<{�a<��a<��a<��a<ڀa<��a<�  �  /�a<Z�a<g�a<��a<��a<ԁa<��a<�a<;�a<=�a<��a<��a<�a<)�a<_�a<Ճa<�a<��a<��a<T�a<�a<D�a<چa<I�a<Їa<:�a<��a<#�a<��a<�a<g�a<��a<K�a<��a<`�a<Ȍa<^�a<Ía<u�a<��a<��a<�a<��a<>�a<��a<N�a<��a<<�a<��a<�a<��a<�a<��a<Еa<i�a<Жa<P�a<�a<[�a<�a<��a<�a<��a<$�a<��a<-�a<��a<�a<��a<ޝa<3�a<��a<Ǟa<+�a<M�a<��a<�a<>�a<u�a<��a<�a<>�a<��a<��a<��a<&�a<L�a<�a<��a<��a<��a<��a<��a<ʢa<ߢa<Тa<�a<��a<�a<=�a<L�a<��a<��a<֣a<�a<�a<5�a<O�a<m�a<Z�a<y�a<m�a<v�a<_�a<V�a<G�a<�a<9�a<�a<%�a<�a<��a<��a<�a<�a<ƣa<��a<��a<z�a<O�a<�a<�a<��a<y�a<�a< �a<��a<��a<V�a<�a<�a<͠a<��a<��a<q�a<o�a<:�a<5�a<�a<�a<��a<o�a<8�a<�a<Şa<S�a<"�a<��a<]�a<1�a<Ȝa<��a<�a<�a<��a<E�a<�a<��a<1�a<��a<^�a<јa<_�a<̗a<?�a<��a<'�a<��a<�a<��a<	�a<��a<.�a<��a<S�a<ˑa<c�a<��a<��a<6�a<��a<a�a<ʎa<a�a<ݍa<X�a<�a<E�a<܋a<7�a<׊a<U�a<�a<n�a<��a<��a<5�a<��a<z�a<�a<��a<L�a<��a<}�a<�a<��a<?�a<ȃa<o�a<�a<��a<��a<�a<�a<��a<��a<�a<B�a<L�a<&�a<)�a<�a<�a<�a<׀a<ހa<��a<��a<��a<��a<��a<X�a<��a<p�a<��a<y�a<��a<Հa<�a<�a<�  �  5�a<`�a<��a<��a<��a<ǁa<�a<�a<.�a<D�a<l�a<��a<ׂa<�a<\�a<��a<�a<q�a<ބa<X�a<ۅa<X�a<��a<D�a<��a<E�a<��a<4�a<��a<�a<�a<��a<u�a<ߋa<c�a<ӌa<k�a<�a<��a<�a<��a<�a<��a<?�a<ȑa<9�a<��a<!�a<��a<�a<��a<�a<R�a<֕a<F�a<Öa<I�a<̗a<_�a<ߘa<}�a<�a<��a<)�a<��a<.�a<��a<$�a<��a<�a<-�a<��a<�a<5�a<y�a<��a<��a<H�a<��a<ݠa< �a<U�a<��a<áa<�a<2�a<\�a<m�a<��a<��a<��a<��a<��a<��a<��a<բa<עa<�a<��a<)�a<L�a<k�a<��a<ˣa<�a<�a<#�a<J�a<`�a<w�a<y�a<u�a<`�a<k�a<c�a<Y�a<=�a<:�a<�a<"�a<�a<�a<�a<��a<ԣa<ˣa<��a<��a<t�a<E�a<
�a<Ӣa<��a<l�a<!�a<�a<��a<w�a<5�a<�a<�a<Πa<��a<��a<v�a<g�a<M�a<�a< �a<ٟa<��a<~�a<I�a<��a<��a<l�a<)�a<ܝa<|�a<4�a<Ӝa<��a<>�a<��a<��a<F�a<ٚa<��a<2�a<ʙa<I�a<Ԙa<D�a<Ǘa<L�a<��a<&�a<��a<�a<~�a<��a<��a<�a<��a<"�a<Ǒa<`�a<�a<��a<�a<��a<J�a<�a<g�a<�a<R�a<ߌa<`�a<�a<b�a<�a<`�a<��a<��a<&�a<��a<L�a<�a<|�a<-�a<��a<\�a<�a<{�a<��a<��a<=�a<Ƀa<`�a<��a<��a<T�a<�a<ρa<��a<��a<]�a<F�a<A�a<4�a<�a<�a<�a<��a<�a<ހa<ǀa<��a<��a<��a<��a<�a<��a<z�a<��a<��a<Āa<܀a<��a<�a<�  �  �a<�a<�a<!�a<E�a<k�a<u�a<��a<��a<��a<ˀa<�a<:�a<^�a<Ɂa<�a<y�a<��a<S�a<уa<V�a<	�a<]�a<��a<Z�a<�a<`�a<чa<P�a<ƈa<5�a<��a<3�a<��a<�a<��a<�a<��a<H�a<��a<c�a<��a<��a<��a<��a<��a<��a<�a<z�a<��a<0�a<��a<��a<~�a<��a<p�a<��a<�a<�a<��a<K�a<՘a<��a<&�a<��a<:�a<��a<-�a<{�a<�a<P�a<��a<ٝa<=�a<}�a<��a<�a<P�a<}�a<�a<�a<^�a<��a<Ԡa<�a<,�a<Y�a<^�a<��a<��a<��a<��a<��a<��a<p�a<��a<��a<��a<��a<�a<�a<&�a<s�a<��a<��a<��a<)�a<@�a<C�a<o�a<^�a<}�a<n�a<h�a<=�a<T�a</�a<�a<=�a<�a<��a<�a<ޢa<�a<٢a<Ϣa<��a<��a<X�a<3�a<�a<¡a<��a<2�a<��a<��a<N�a<3�a<�a<՟a<��a<��a<J�a<R�a<A�a<3�a<O�a<�a<�a<��a<��a<q�a<1�a<��a<��a<h�a<
�a<ݜa<e�a<"�a<�a<v�a<2�a<��a<��a<G�a<�a<��a<�a<Øa<+�a<җa<>�a<��a<<�a<p�a<�a<8�a<��a<(�a<��a<"�a<��a<>�a<��a<w�a<�a<͏a<f�a<�a<��a<�a<��a<�a<��a<3�a<��a<�a<��a<�a<��a<2�a<��a<$�a<�a<[�a< �a<��a<6�a<˅a<b�a< �a<{�a<,�a<��a<X�a<��a<=�a<ցa<P�a<�a<��a<y�a<+�a<	�a<�a<�a<�a<�a<�a<�a<�a<�a<{a<�a<`a<ma<Qa<Ba<a<,a<a<a<<a<a<,a<^a<Wa<�a<�a<�  �  �a< �a<�a<3�a<C�a<a�a<k�a<v�a<��a<��a<�a<�a<<�a<j�a<��a<�a<y�a<ނa<X�a<ԃa<F�a<Ʉa<X�a<�a<a�a<�a<l�a<�a<O�a<��a<)�a<��a<�a<��a<�a<��a<#�a<��a<B�a<ȍa<d�a<�a<��a<�a<��a<�a<��a<��a<V�a<Ēa<7�a<��a<�a<��a<�a<q�a<��a<��a<�a<��a<C�a<��a<l�a<��a<��a<�a<��a<*�a<��a<��a<I�a<��a<�a<5�a<g�a<a<��a<C�a<��a<ɟa<�a<R�a<��a<ՠa<�a<@�a<d�a<h�a<~�a<��a<~�a<}�a<��a<��a<��a<��a<��a<��a<��a<�a<�a<?�a<i�a<��a<��a<�a<�a<:�a<X�a<m�a<y�a<}�a<d�a<b�a<P�a<I�a<2�a<.�a<�a<�a<�a<��a<�a<�a<Ңa<Тa<��a<��a<k�a<1�a<�a<��a<l�a<0�a<��a<��a<k�a<4�a<�a<˟a<��a<��a<g�a<W�a<E�a<#�a<�a<�a<�a<Ǟa<��a<}�a<F�a<��a<��a<\�a<�a<��a<o�a< �a<a<��a<'�a<�a<��a<G�a<�a<��a</�a<��a<=�a<��a<3�a<��a<�a<w�a<�a<M�a<a<6�a<��a<!�a<��a<D�a<Րa<o�a<�a<��a<<�a<�a<|�a<�a<��a<6�a<��a<-�a<��a<�a<��a<�a<��a<�a<��a<4�a<��a<[�a<�a<��a<7�a<߅a<v�a<�a<��a<�a<��a<�a<��a<B�a<Ձa<k�a<�a<��a<r�a<0�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<|a<ma<Ga<<a<'a<"a<a<a<a<'a<3a<Ma<ga<�a<�a<�  �  �a<�a<�a<1�a<H�a<h�a<��a<��a<��a<��a<��a<�a<<�a<��a<a<�a<v�a<�a<S�a<�a<m�a<ׄa<~�a<�a<h�a<�a<H�a<Ňa<>�a<��a<�a<��a<�a<��a<�a<f�a<,�a<��a<+�a<��a<V�a<�a<o�a<��a<w�a<�a<��a<�a<�a<ْa<_�a<��a<!�a<��a<�a<|�a<��a<��a<�a<��a<B�a<�a<��a<!�a<��a<+�a<��a<�a<u�a<ٜa<:�a<��a<ӝa<%�a<`�a<˞a<�a<?�a<��a<��a<�a<D�a<��a<àa<�a<�a<H�a<q�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<աa<�a<�a<D�a<e�a<��a<¢a<�a<)�a<<�a<Y�a<H�a<_�a<_�a<e�a<U�a<K�a<3�a<&�a<8�a<�a<�a<��a<�a<�a<բa<Ңa<��a<��a<m�a<h�a<6�a<�a<ۡa<u�a<Z�a<��a<��a<u�a<4�a<�a<Οa<��a<��a<x�a<R�a<T�a<K�a<�a<(�a<�a<Ξa<��a<Y�a<%�a<�a<��a<P�a<�a<��a<s�a<�a<��a<��a< �a<ؚa<��a<:�a<�a<|�a<�a<��a<H�a<��a<Q�a<��a<�a<��a<ޔa<\�a<��a<8�a<��a<)�a<��a<@�a<�a<m�a<5�a<��a<a�a<	�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<��a<��a<��a<��a<=�a<��a<\�a<�a<��a<%�a<��a<O�a<�a<��a<�a<��a<-�a<̂a<\�a<сa<��a<�a<ʀa<y�a<G�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<ba<ba<Oa<Ha<.a<"a<a<a<$a<�~a<.a<*a<9a<da<ya<�a<�  �  �a<�a<�a<+�a<M�a<]�a<t�a<��a<��a<��a<��a<�a<O�a<��a<�a<+�a<��a<��a<{�a<�a<^�a<�a<]�a<�a<h�a<�a<m�a<Їa<E�a<��a<�a<{�a<�a<c�a<��a<x�a<�a<��a<�a<��a<C�a<�a<o�a<	�a<��a<�a<��a<�a<z�a<�a<I�a<˓a<6�a<��a<�a<��a<&�a<��a<0�a<̗a<j�a<�a<��a<#�a<��a<8�a<��a<,�a<��a<ݜa<A�a<�a<ǝa<�a<`�a<��a<�a<'�a<Z�a<a<��a<@�a<��a<ʠa<��a<>�a<X�a<k�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<֡a<�a<�a<%�a<_�a<��a<��a<֢a<��a<�a<G�a<Q�a<u�a<i�a<a�a<\�a<F�a<0�a<+�a<�a<��a<��a<�a<ܢa<�a<ʢa<ʢa<Ţa<��a<��a<��a<c�a<;�a<��a<��a<��a<B�a<�a<Рa<��a<G�a<�a<�a<��a<��a<��a<z�a<a�a<;�a<6�a<�a<��a<Ξa<��a<~�a</�a<�a<��a<J�a<�a<��a<C�a<�a<��a<L�a<�a<Ța<u�a<'�a<�a<{�a<%�a<Ƙa<9�a<Ηa</�a<��a<$�a<��a<	�a<p�a<Гa<J�a<Вa<S�a<͑a<Y�a<��a<��a<#�a<��a<c�a<�a<��a<�a<��a<.�a<��a<$�a<��a<��a<z�a<��a<\�a< �a<��a<�a<��a<=�a<�a<��a<,�a<ƅa<s�a<��a<��a<"�a<��a<B�a<a<]�a<��a<��a<*�a<Հa<��a<\�a<&�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<la<Qa<>a< a<a<a<�~a<�~a<�~a<�~a<a<9a<Ca<na<�a<�  �  �a<�a<	�a<�a<`�a<|�a<��a<��a<��a<��a<�a<5�a<q�a<��a< �a<;�a<��a<�a<��a<�a<c�a<�a<j�a<�a<o�a<چa<R�a<��a<0�a<��a<�a<_�a<�a<T�a<ъa<i�a<̋a<��a<��a<��a<-�a<ǎa<_�a<�a<��a<��a<��a<�a<��a<��a<R�a<�a<6�a<Ĕa<0�a<��a<0�a<��a<Y�a<Ηa<��a< �a<��a<=�a<��a<M�a<��a<�a<o�a<̜a<$�a<a�a<ʝa<�a<M�a<n�a<ўa<�a<I�a<��a<ҟa<C�a<^�a<��a<�a<�a<N�a<l�a<��a<��a<áa<��a<��a<áa<��a<ѡa<ǡa<�a<�a<#�a<E�a<^�a<��a<��a<��a<�a<1�a<\�a<@�a<a�a<K�a<W�a<6�a<@�a<#�a<�a<�a<آa<�a<âa<עa<ˢa<��a<ʢa<��a<��a<��a<��a<Q�a<N�a<�a<١a<��a<B�a<1�a<ՠa<��a<i�a<"�a<�a<˟a<��a<��a<��a<v�a<A�a<T�a<�a<�a<֞a<��a<c�a<�a<۝a<q�a<K�a<Мa<��a<3�a<�a<��a<2�a<�a<��a<v�a<�a<��a<k�a<
�a<��a<*�a<�a<D�a<іa<7�a<��a<�a<q�a<��a<d�a<ؒa<]�a<�a<��a<��a<��a<0�a<Ϗa<~�a<�a<��a<�a<��a<�a<��a<�a<l�a<�a<S�a<�a<G�a<�a<i�a<�a<��a<�a<�a<^�a<�a<��a<U�a<��a<��a<<�a<��a<`�a<ɂa<n�a<�a<��a<O�a<�a<��a<b�a<E�a<�a<�a<�a<�a<�a<�a<�a<�a<xa<{a<Na<Ga<a<a<�~a<�~a<�~a<�~a<�~a<�~a<a<a</a<na<va<�  �  �a<�a<�a<.�a<J�a<^�a<��a<��a<�a<��a<�a<_�a<��a<΁a<�a<i�a<Ȃa<=�a<��a<�a<��a<�a<��a<�a<n�a<�a<M�a<��a<,�a<��a<�a<^�a<��a<>�a<��a<*�a<ԋa<J�a<�a<��a< �a<Îa<`�a<��a<|�a<�a<��a<�a<��a<��a<��a<ܓa<c�a<ؔa<L�a<֕a<Z�a<ؖa<h�a<�a<x�a<.�a<��a<6�a<��a<'�a<��a<�a<t�a<Ϝa<�a<V�a<��a<�a<�a<s�a<��a<�a<=�a<o�a<ӟa<�a<X�a<��a<�a<�a<J�a<w�a<��a<��a<��a<͡a<ѡa<��a<�a<�a<�a<	�a<"�a<9�a<h�a<{�a<��a<�a<�a<�a<�a<<�a<Z�a<P�a<V�a<L�a<5�a<'�a<�a<�a<עa<٢a<��a<��a<��a<��a<��a<��a<��a<��a<��a<w�a<f�a<8�a<��a<�a<��a<��a<.�a<�a<Ơa<��a<R�a<#�a<��a<ןa<Ɵa<��a<��a<u�a<N�a<,�a<�a<՞a<��a<^�a<�a<֝a<s�a<�a<Μa<a�a<�a<Ǜa<h�a<:�a<֚a<��a<Z�a<�a<��a<l�a<�a<��a<N�a<��a<E�a<͖a<<�a<̕a<�a<��a<�a<�a<�a<��a<�a<��a<+�a<��a<^�a<ޏa<v�a<�a<��a<&�a<��a<�a<��a<�a<b�a<�a<N�a<��a<M�a<��a<C�a<�a<e�a<�a<��a<X�a<�a<��a<P�a<�a<��a<�a<a<Y�a<�a<��a<�a<Ɓa<c�a<�a<πa<��a<[�a<@�a<�a<�a<�a<�a<�a<�a<�a<�a<ka<Ya<<a<a<a<�~a<�~a<�~a<�~a<�~a<�~a<�~a<�~a<"a<Oa<va<�  �  {a<�a<�a<2�a<Y�a<t�a<��a<��a<��a<�a<X�a<{�a<��a<��a<(�a<��a<̂a<k�a<��a<!�a<��a<��a<��a<�a<��a<Նa<B�a<��a<��a<�a<��a<c�a<��a<�a<��a<�a<��a<�a<��a<b�a<�a<��a<6�a<��a<f�a<5�a<��a<'�a<��a<�a<��a<�a<��a<ޔa<i�a<��a<r�a<��a<o�a<H�a<��a<;�a<��a<>�a<՚a<)�a<ӛa<��a<v�a<��a<��a<H�a<v�a<��a<�a<I�a<��a<Ԟa<
�a<N�a<۟a<�a<Q�a<}�a<ڠa<�a<<�a<��a<��a<ȡa<��a<֡a<ߡa<�a<�a<�a<�a<�a<N�a<H�a<z�a<âa<��a<��a<�a<3�a<6�a<G�a<f�a<@�a<\�a<�a<(�a<��a<��a<�a<��a<��a<��a<��a<u�a<��a<��a<|�a<��a<p�a<��a<j�a<i�a<H�a<�a<�a<��a<��a<9�a<*�a<�a<��a<��a<5�a<(�a<۟a<��a<��a<��a<��a<E�a<M�a<��a<�a<��a<S�a<�a<��a<o�a<�a<Ԝa<K�a<�a<��a<K�a<�a<��a<��a<,�a<�a<��a<B�a<�a<��a<g�a<×a<d�a<ߖa<G�a<וa<+�a<�a<�a<��a<%�a<��a<)�a<��a<r�a<��a<k�a<�a<~�a<"�a<��a<C�a<~�a<�a<k�a<܋a<T�a<��a<]�a<��a<#�a<��a<2�a<��a<D�a<$�a<��a<Q�a<߅a<��a<K�a<�a<��a<�a<��a<S�a<��a<��a<2�a<��a<e�a<=�a<��a<��a<j�a<Q�a<T�a<�a<�a<�a<�a<�a<�a<�a<[a<_a<a<
a<�~a<�~a<�~a<�~a<�~a<�~a<�~a<�~a<�~a<a<!a<la<�  �  �a<�a<�a< �a<[�a<��a<��a<�a<�a<1�a<]�a<{�a<āa<�a<K�a<��a<��a<Z�a<ڃa<H�a<��a<+�a<��a<��a<z�a<ˆa<&�a<��a<�a<p�a<��a<�a<��a<��a<{�a<��a<��a<�a<��a<7�a<��a<��a<:�a<ڏa<f�a<�a<��a<'�a<��a<9�a<��a<$�a<��a<�a<��a<�a<��a<+�a<��a<:�a<ʘa<D�a<�a<^�a<Кa<<�a<��a<��a<X�a<��a<�a<<�a<V�a<��a<�a< �a<m�a<��a<�a<G�a<��a<ԟa<G�a<t�a<Ša<��a<3�a<��a<��a<ša<�a<�a<��a<�a<�a<�a<D�a<:�a<a�a<{�a<��a<��a<ܢa<��a<&�a<7�a<C�a<P�a<M�a<1�a<=�a<'�a<�a<�a<��a<Ƣa<��a<��a<~�a<v�a<m�a<{�a<^�a<q�a<��a<y�a<y�a<V�a<X�a<I�a< �a<��a<סa<��a<i�a</�a<�a<��a<��a<W�a<G�a<
�a<�a<ٟa<��a<��a<q�a<F�a<
�a<�a<��a<7�a<��a<��a<a�a<�a<��a<>�a<؛a<��a<;�a<�a<��a<f�a<�a<ݙa<��a<F�a<��a<��a<F�a<ԗa<d�a<�a<z�a<ޕa<a�a<ܔa<;�a<Γa<5�a<��a<U�a<đa<d�a<��a<u�a<�a<��a<�a<��a<%�a<�a<��a<g�a<΋a<G�a<��a<�a<��a<��a<��a<�a<��a<=�a<܆a<v�a<G�a<օa<��a<-�a<ڄa<��a</�a<݃a<|�a<�a<��a<[�a<�a<��a<c�a< �a<Ӏa<��a<b�a<Q�a<-�a<�a<�a<�a<�a<�a<�a<La<@a<a<�~a<�~a<�~a<�~a<�~a<z~a<|~a<�~a<�~a<�~a<�~a<a<\a<�  �  �a<�a<�a</�a<G�a<��a<��a<�a<��a<T�a<g�a<��a<�a<�a<��a<��a<4�a<��a<��a<]�a<��a<3�a<��a<�a<\�a<�a<6�a<��a<��a<-�a<��a<��a<t�a<�a<I�a<܊a<Y�a<�a<��a<@�a<܍a<w�a<C�a<��a<��a<�a<��a<+�a<��a<>�a<��a<M�a<��a<?�a<��a<2�a<��a<)�a<җa<:�a<�a<O�a<�a<Z�a<Κa<K�a<��a<�a<D�a<��a<՜a<�a<`�a<z�a<ӝa<��a<D�a<��a<؞a<0�a<i�a<؟a<�a<s�a<Ơa<��a<X�a<^�a<��a<��a<�a<�a<�a<.�a<)�a<P�a<<�a<x�a<w�a<��a<Ģa<âa<�a<��a<,�a<*�a<I�a<E�a<S�a<V�a<'�a<+�a<�a<�a<��a<��a<��a<_�a<j�a<F�a<U�a<M�a<Q�a<r�a<J�a<|�a<j�a<x�a<g�a<5�a<,�a<��a<�a<��a<��a<9�a<�a<�a<��a<��a<D�a<C�a<�a<�a<͟a<��a<y�a<;�a<�a<Þa<��a<G�a<��a<��a<�a<�a<j�a<�a<a<Y�a<�a<��a<��a<.�a<
�a<��a<p�a<O�a<ݘa<��a<4�a<ݗa<h�a<�a<�a<�a<��a<ڔa<v�a<֓a<b�a<�a<S�a<��a<d�a<�a<�a<�a<��a<�a<��a<�a<��a<�a<p�a<��a<�a<��a<�a<r�a<׈a<]�a<߇a<�a<&�a<��a<z�a<�a<Յa<��a<3�a<��a<{�a<C�a<ԃa<~�a<�a<Âa<v�a<	�a<́a<[�a<>�a<�a<��a<��a<U�a<X�a<�a<�a<�a<�a<�a<�a<qa<*a<a<�~a<�~a<�~a<k~a<i~a<L~a<i~a<\~a<�~a<�~a<�~a<a<a<�  �  da<�a<�a< �a<Y�a<��a<ƀa<��a<%�a<P�a<~�a<Ёa<��a<@�a<��a<Ղa<7�a<��a<��a<g�a<ۄa<>�a<��a<$�a<n�a<نa<�a<��a<ۇa<*�a<��a<��a<P�a<ŉa<C�a<ʊa<G�a<܋a<~�a<*�a<ˍa<n�a<&�a<��a<r�a<�a<��a<J�a<ƒa<R�a<ʓa<J�a<Ɣa<T�a<��a<L�a<Ԗa<<�a<�a<d�a<�a<n�a<��a<m�a<�a<Y�a<��a<�a<4�a<��a<ɜa<�a<G�a<w�a<��a<�a<7�a<{�a<��a<�a<k�a<ßa< �a<^�a<��a<�a<C�a<p�a<��a<ءa<�a<�a<�a<0�a<I�a<Z�a<Y�a<��a<��a<��a<ޢa<ܢa<�a<!�a<?�a<I�a<d�a<T�a<I�a<6�a<�a<�a<ޢa<Ѣa<��a<��a<e�a<N�a<M�a<7�a<3�a<;�a<K�a<W�a<I�a<Z�a<S�a<X�a<W�a<G�a<E�a<�a<�a<��a<��a<P�a<8�a<�a<Ša<��a<e�a<F�a<)�a<��a<ןa<��a<��a<X�a</�a<Ԟa<��a</�a<�a<��a<�a<Ԝa<l�a<��a<��a<T�a<�a<��a<g�a<*�a<��a<��a<h�a<3�a<Ϙa<��a<7�a<�a<��a<�a<��a<	�a<��a< �a<��a<�a<|�a<�a<g�a<�a<��a<�a<��a<5�a<��a<;�a<��a<�a<��a<֌a<U�a<��a<�a<�a<��a<I�a<Èa<Q�a<هa<d�a<��a<��a<f�a< �a<��a<z�a<�a<�a<��a<S�a<��a<��a<>�a<Ԃa<x�a<)�a<ׁa<x�a<M�a<	�a<ǀa<��a<n�a<U�a<6�a<�a<�a<�a<�a<�a<Qa<a<�~a<�~a<�~a<�~a<_~a<E~a<;~a<L~a<M~a<d~a<�~a<�~a<�~a<a<�  �  Na<�a<�a<�a<\�a<w�a<��a<�a<4�a<\�a<��a<ˁa<�a<l�a<{�a<�a<I�a<��a<�a<x�a<�a<>�a<��a<��a<x�a<͆a<4�a<��a<ɇa<C�a<t�a<�a<B�a<��a<*�a<��a<<�a<a<v�a<�a<эa<v�a<�a<ڏa<l�a<�a<��a<'�a<��a<K�a<ݓa<N�a<�a<N�a<��a<_�a<ؖa<��a<�a<z�a<�a<��a<��a<e�a<њa<7�a<��a<��a<^�a<��a<̜a<�a<!�a<m�a<��a<ڝa<�a<[�a<��a<�a<S�a<��a<�a<O�a<��a<�a<6�a<}�a<��a<ɡa<�a<�a<1�a<A�a<V�a<d�a<��a<p�a<��a<Тa<٢a<�a<�a<3�a<8�a<A�a<=�a<Q�a<H�a<7�a<6�a<��a<�a<��a<��a<x�a<O�a<C�a<*�a<,�a<�a<*�a<+�a<:�a<`�a<D�a<o�a<_�a<T�a<J�a<�a<
�a<�a<͡a<��a<r�a<3�a<�a<�a<��a<��a<X�a<0�a<�a<�a<��a<��a<O�a<�a<ޞa<��a<E�a<�a<s�a<3�a<��a<Q�a<�a<��a<;�a<�a<��a<N�a<#�a<Ιa<��a<p�a<!�a<��a<��a<@�a<ϗa<d�a<��a<��a<�a<��a<�a<��a<'�a<��a<�a<��a<�a<��a<�a<��a<.�a<��a<�a<��a<�a<��a<��a<M�a<��a< �a<Y�a<։a</�a<��a<)�a<��a<S�a<�a<��a<:�a<�a<��a<��a<;�a<ބa<��a<+�a<�a<��a<C�a<�a<��a<6�a<�a<��a<6�a<+�a<�a<��a<��a<]�a<H�a<�a<�a<�a<�a<a<Ra<8a<�~a<�~a<�~a<a~a<Q~a</~a<0~a<)~a<A~a<P~a<|~a<�~a<�~a<5a<�  �  Ca<�a<�a<�a<a�a<��a<݀a<�a<2�a<i�a<��a<߁a<�a<h�a<��a<�a<W�a<��a<�a<��a<�a<]�a<��a<�a<t�a<ˆa<#�a<h�a<��a<�a<w�a<ۈa<A�a<��a<�a<��a<,�a<ċa<^�a<�a<��a<P�a<��a<��a<b�a<�a<��a<N�a<�a<^�a<�a<_�a<�a<\�a<�a<d�a<�a<z�a<�a<��a<�a<��a<	�a<��a<��a<Z�a<��a<�a<9�a<l�a<��a<�a<#�a<W�a<��a<ҝa<�a<L�a<��a<��a<G�a<��a<�a<=�a<��a<�a<2�a<s�a<��a<�a<�a<�a<>�a<M�a<o�a<n�a<��a<��a<��a<Тa<�a<�a<�a<0�a<J�a<a�a<_�a<[�a<A�a<8�a<�a<�a<Ȣa<��a<��a<i�a<R�a<.�a<(�a<�a< �a<�a<-�a<6�a<7�a<9�a<M�a<Z�a<N�a<O�a<:�a<*�a<�a<ˡa<��a<t�a<F�a<�a<�a<��a<��a<f�a<I�a<�a<��a<��a<��a<h�a<'�a<ڞa<��a<5�a<ȝa<f�a<	�a<��a<L�a<�a<��a<&�a<ٚa<��a<P�a<�a<ҙa<��a<J�a<
�a<Иa<��a<5�a<�a<��a<!�a<��a<#�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<1�a<��a<@�a<ʏa<A�a<��a<�a<v�a<یa<,�a<��a<��a<Z�a<��a<3�a<��a< �a<��a<O�a<�a<��a<<�a<�a<��a<X�a<!�a<لa<��a<M�a<��a<��a<D�a<�a<��a<O�a<�a<��a<W�a<+�a<�a<��a<��a<j�a<F�a<)�a<�a<�a<�a<ya<Ra<a<�~a<�~a<�~a<f~a<B~a<2~a<~a<'~a<)~a<R~a<p~a<�~a<�~a<a<�  �  �a<�a<�a<�a<Q�a<��a<Àa<�a<;�a<o�a<��a<��a<�a<_�a<Ղa<��a<W�a<ʃa<�a<��a<�a<[�a<��a< �a<_�a<Նa<.�a<��a<��a<�a<��a<a<"�a<��a<�a<��a<"�a<ȋa<F�a<�a<��a<n�a<9�a<��a<z�a<��a<��a<8�a<͒a<]�a<�a<h�a<�a<|�a<וa<w�a<�a<f�a<�a<��a<�a<��a<�a<w�a<ۚa<Y�a<��a<�a<E�a<��a<ќa<�a<*�a<B�a<��a<ŝa<
�a<L�a<��a<�a<2�a<��a<�a<|�a<��a<��a<E�a<a�a<��a<ȡa<	�a<'�a<@�a<:�a<v�a<v�a<��a<Ţa<��a<Ƣa<�a<��a< �a<:�a<K�a<I�a<U�a<M�a<<�a<E�a<�a<'�a<Ӣa<��a<��a<L�a<Q�a<#�a<3�a<�a< �a<�a<�a<3�a<<�a<x�a<S�a<d�a<N�a<?�a<7�a<�a<�a<ԡa<��a<g�a<^�a<�a<�a<�a<��a<f�a<S�a<�a<��a<˟a<��a<L�a<+�a<ƞa<��a<?�a<�a<��a<�a<��a<3�a<̛a<��a<%�a<ߚa<��a<S�a<�a<ՙa<��a<g�a<E�a<٘a<��a<*�a<�a<u�a<�a<��a<'�a<��a<�a<��a<
�a<��a</�a<��a<1�a<��a<-�a<��a<C�a<��a<(�a<��a<�a<��a<�a<[�a<��a<�a<b�a<��a<1�a<��a<#�a<��a<B�a<ۆa<{�a<H�a<�a<ޅa<z�a<+�a<�a<~�a<O�a<��a<��a<M�a<�a<��a<V�a<�a<��a<��a<)�a<�a<ހa<��a<r�a<P�a<*�a<�a<�a<�a<ta<`a<a<a<�~a<�~a<]~a<%~a<1~a<~a<2~a<~a<Q~a<V~a<�~a<�~a<a<�  �  Ca<�a<�a<�a<a�a<��a<݀a<�a<2�a<i�a<��a<߁a<�a<h�a<��a<�a<W�a<��a<�a<��a<�a<]�a<��a<�a<t�a<ˆa<#�a<h�a<��a<�a<w�a<ۈa<A�a<��a<�a<��a<,�a<ċa<^�a<�a<��a<P�a<��a<��a<b�a<�a<��a<N�a<�a<^�a<�a<_�a<�a<\�a<�a<d�a<�a<z�a<�a<��a<�a<��a<	�a<��a<��a<Z�a<��a<�a<9�a<l�a<��a<�a<#�a<W�a<��a<ҝa<�a<L�a<��a<��a<G�a<��a<�a<=�a<��a<�a<2�a<s�a<��a<�a<�a<�a<>�a<M�a<o�a<n�a<��a<��a<��a<Тa<�a<�a<�a<0�a<J�a<a�a<_�a<[�a<A�a<8�a<�a<�a<Ȣa<��a<��a<i�a<R�a<.�a<(�a<�a< �a<�a<-�a<6�a<7�a<9�a<M�a<Z�a<N�a<O�a<:�a<*�a<�a<ˡa<��a<t�a<F�a<�a<�a<��a<��a<f�a<I�a<�a<��a<��a<��a<h�a<'�a<ڞa<��a<5�a<ȝa<f�a<	�a<��a<L�a<�a<��a<&�a<ٚa<��a<P�a<�a<ҙa<��a<J�a<
�a<Иa<��a<5�a<�a<��a<!�a<��a<#�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<1�a<��a<@�a<ʏa<A�a<��a<�a<v�a<یa<,�a<��a<��a<Z�a<��a<3�a<��a< �a<��a<O�a<�a<��a<<�a<�a<��a<X�a<!�a<لa<��a<M�a<��a<��a<D�a<�a<��a<O�a<�a<��a<W�a<+�a<�a<��a<��a<j�a<F�a<)�a<�a<�a<�a<ya<Ra<a<�~a<�~a<�~a<f~a<B~a<2~a<~a<'~a<)~a<R~a<p~a<�~a<�~a<a<�  �  Na<�a<�a<�a<\�a<w�a<��a<�a<4�a<\�a<��a<ˁa<�a<l�a<{�a<�a<I�a<��a<�a<x�a<�a<>�a<��a<��a<x�a<͆a<4�a<��a<ɇa<C�a<t�a<�a<B�a<��a<*�a<��a<<�a<a<v�a<�a<эa<v�a<�a<ڏa<l�a<�a<��a<'�a<��a<K�a<ݓa<N�a<�a<N�a<��a<_�a<ؖa<��a<�a<z�a<�a<��a<��a<e�a<њa<7�a<��a<��a<^�a<��a<̜a<�a<!�a<m�a<��a<ڝa<�a<[�a<��a<�a<S�a<��a<�a<O�a<��a<�a<6�a<}�a<��a<ɡa<�a<�a<1�a<A�a<V�a<d�a<��a<p�a<��a<Тa<٢a<�a<�a<3�a<8�a<A�a<=�a<Q�a<H�a<7�a<6�a<��a<�a<��a<��a<x�a<O�a<C�a<*�a<,�a<�a<*�a<+�a<:�a<`�a<D�a<o�a<_�a<T�a<J�a<�a<
�a<�a<͡a<��a<r�a<3�a<�a<�a<��a<��a<X�a<0�a<�a<�a<��a<��a<O�a<�a<ޞa<��a<E�a<�a<s�a<3�a<��a<Q�a<�a<��a<;�a<�a<��a<N�a<#�a<Ιa<��a<p�a<!�a<��a<��a<@�a<ϗa<d�a<��a<��a<�a<��a<�a<��a<'�a<��a<�a<��a<�a<��a<�a<��a<.�a<��a<�a<��a<�a<��a<��a<M�a<��a< �a<Y�a<։a</�a<��a<)�a<��a<S�a<�a<��a<:�a<�a<��a<��a<;�a<ބa<��a<+�a<�a<��a<C�a<�a<��a<6�a<�a<��a<6�a<+�a<�a<��a<��a<]�a<H�a<�a<�a<�a<�a<a<Ra<8a<�~a<�~a<�~a<a~a<Q~a</~a<0~a<)~a<A~a<P~a<|~a<�~a<�~a<5a<�  �  da<�a<�a< �a<Y�a<��a<ƀa<��a<%�a<P�a<~�a<Ёa<��a<@�a<��a<Ղa<7�a<��a<��a<g�a<ۄa<>�a<��a<$�a<n�a<نa<�a<��a<ۇa<*�a<��a<��a<P�a<ŉa<C�a<ʊa<G�a<܋a<~�a<*�a<ˍa<n�a<&�a<��a<r�a<�a<��a<J�a<ƒa<R�a<ʓa<J�a<Ɣa<T�a<��a<L�a<Ԗa<<�a<�a<d�a<�a<n�a<��a<m�a<�a<Y�a<��a<�a<4�a<��a<ɜa<�a<G�a<w�a<��a<�a<7�a<{�a<��a<�a<k�a<ßa< �a<^�a<��a<�a<C�a<p�a<��a<ءa<�a<�a<�a<0�a<I�a<Z�a<Y�a<��a<��a<��a<ޢa<ܢa<�a<!�a<?�a<I�a<d�a<T�a<I�a<6�a<�a<�a<ޢa<Ѣa<��a<��a<e�a<N�a<M�a<7�a<3�a<;�a<K�a<W�a<I�a<Z�a<S�a<X�a<W�a<G�a<E�a<�a<�a<��a<��a<P�a<8�a<�a<Ša<��a<e�a<F�a<)�a<��a<ןa<��a<��a<X�a</�a<Ԟa<��a</�a<�a<��a<�a<Ԝa<l�a<��a<��a<T�a<�a<��a<g�a<*�a<��a<��a<h�a<3�a<Ϙa<��a<7�a<�a<��a<�a<��a<	�a<��a< �a<��a<�a<|�a<�a<g�a<�a<��a<�a<��a<5�a<��a<;�a<��a<�a<��a<֌a<U�a<��a<�a<�a<��a<I�a<Èa<Q�a<هa<d�a<��a<��a<f�a< �a<��a<z�a<�a<�a<��a<S�a<��a<��a<>�a<Ԃa<x�a<)�a<ׁa<x�a<M�a<	�a<ǀa<��a<n�a<U�a<6�a<�a<�a<�a<�a<�a<Qa<a<�~a<�~a<�~a<�~a<_~a<E~a<;~a<L~a<M~a<d~a<�~a<�~a<�~a<a<�  �  �a<�a<�a</�a<G�a<��a<��a<�a<��a<T�a<g�a<��a<�a<�a<��a<��a<4�a<��a<��a<]�a<��a<3�a<��a<�a<\�a<�a<6�a<��a<��a<-�a<��a<��a<t�a<�a<I�a<܊a<Y�a<�a<��a<@�a<܍a<w�a<C�a<��a<��a<�a<��a<+�a<��a<>�a<��a<M�a<��a<?�a<��a<2�a<��a<)�a<җa<:�a<�a<O�a<�a<Z�a<Κa<K�a<��a<�a<D�a<��a<՜a<�a<`�a<z�a<ӝa<��a<D�a<��a<؞a<0�a<i�a<؟a<�a<s�a<Ơa<��a<X�a<^�a<��a<��a<�a<�a<�a<.�a<)�a<P�a<<�a<x�a<w�a<��a<Ģa<âa<�a<��a<,�a<*�a<I�a<E�a<S�a<V�a<'�a<+�a<�a<�a<��a<��a<��a<_�a<j�a<F�a<U�a<M�a<Q�a<r�a<J�a<|�a<j�a<x�a<g�a<5�a<,�a<��a<�a<��a<��a<9�a<�a<�a<��a<��a<D�a<C�a<�a<�a<͟a<��a<y�a<;�a<�a<Þa<��a<G�a<��a<��a<�a<�a<j�a<�a<a<Y�a<�a<��a<��a<.�a<
�a<��a<p�a<O�a<ݘa<��a<4�a<ݗa<h�a<�a<�a<�a<��a<ڔa<v�a<֓a<b�a<�a<S�a<��a<d�a<�a<�a<�a<��a<�a<��a<�a<��a<�a<p�a<��a<�a<��a<�a<r�a<׈a<]�a<߇a<�a<&�a<��a<z�a<�a<Յa<��a<3�a<��a<{�a<C�a<ԃa<~�a<�a<Âa<v�a<	�a<́a<[�a<>�a<�a<��a<��a<U�a<X�a<�a<�a<�a<�a<�a<�a<qa<*a<a<�~a<�~a<�~a<k~a<i~a<L~a<i~a<\~a<�~a<�~a<�~a<a<a<�  �  �a<�a<�a< �a<[�a<��a<��a<�a<�a<1�a<]�a<{�a<āa<�a<K�a<��a<��a<Z�a<ڃa<H�a<��a<+�a<��a<��a<z�a<ˆa<&�a<��a<�a<p�a<��a<�a<��a<��a<{�a<��a<��a<�a<��a<7�a<��a<��a<:�a<ڏa<f�a<�a<��a<'�a<��a<9�a<��a<$�a<��a<�a<��a<�a<��a<+�a<��a<:�a<ʘa<D�a<�a<^�a<Кa<<�a<��a<��a<X�a<��a<�a<<�a<V�a<��a<�a< �a<m�a<��a<�a<G�a<��a<ԟa<G�a<t�a<Ša<��a<3�a<��a<��a<ša<�a<�a<��a<�a<�a<�a<D�a<:�a<a�a<{�a<��a<��a<ܢa<��a<&�a<7�a<C�a<P�a<M�a<1�a<=�a<'�a<�a<�a<��a<Ƣa<��a<��a<~�a<v�a<m�a<{�a<^�a<q�a<��a<y�a<y�a<V�a<X�a<I�a< �a<��a<סa<��a<i�a</�a<�a<��a<��a<W�a<G�a<
�a<�a<ٟa<��a<��a<q�a<F�a<
�a<�a<��a<7�a<��a<��a<a�a<�a<��a<>�a<؛a<��a<;�a<�a<��a<f�a<�a<ݙa<��a<F�a<��a<��a<F�a<ԗa<d�a<�a<z�a<ޕa<a�a<ܔa<;�a<Γa<5�a<��a<U�a<đa<d�a<��a<u�a<�a<��a<�a<��a<%�a<�a<��a<g�a<΋a<G�a<��a<�a<��a<��a<��a<�a<��a<=�a<܆a<v�a<G�a<օa<��a<-�a<ڄa<��a</�a<݃a<|�a<�a<��a<[�a<�a<��a<c�a< �a<Ӏa<��a<b�a<Q�a<-�a<�a<�a<�a<�a<�a<�a<La<@a<a<�~a<�~a<�~a<�~a<�~a<z~a<|~a<�~a<�~a<�~a<�~a<a<\a<�  �  {a<�a<�a<2�a<Y�a<t�a<��a<��a<��a<�a<X�a<{�a<��a<��a<(�a<��a<̂a<k�a<��a<!�a<��a<��a<��a<�a<��a<Նa<B�a<��a<��a<�a<��a<c�a<��a<�a<��a<�a<��a<�a<��a<b�a<�a<��a<6�a<��a<f�a<5�a<��a<'�a<��a<�a<��a<�a<��a<ޔa<i�a<��a<r�a<��a<o�a<H�a<��a<;�a<��a<>�a<՚a<)�a<ӛa<��a<v�a<��a<��a<H�a<v�a<��a<�a<I�a<��a<Ԟa<
�a<N�a<۟a<�a<Q�a<}�a<ڠa<�a<<�a<��a<��a<ȡa<��a<֡a<ߡa<�a<�a<�a<�a<�a<N�a<H�a<z�a<âa<��a<��a<�a<3�a<6�a<G�a<f�a<@�a<\�a<�a<(�a<��a<��a<�a<��a<��a<��a<��a<u�a<��a<��a<|�a<��a<p�a<��a<j�a<i�a<H�a<�a<�a<��a<��a<9�a<*�a<�a<��a<��a<5�a<(�a<۟a<��a<��a<��a<��a<E�a<M�a<��a<�a<��a<S�a<�a<��a<o�a<�a<Ԝa<K�a<�a<��a<K�a<�a<��a<��a<,�a<�a<��a<B�a<�a<��a<g�a<×a<d�a<ߖa<G�a<וa<+�a<�a<�a<��a<%�a<��a<)�a<��a<r�a<��a<k�a<�a<~�a<"�a<��a<C�a<~�a<�a<k�a<܋a<T�a<��a<]�a<��a<#�a<��a<2�a<��a<D�a<$�a<��a<Q�a<߅a<��a<K�a<�a<��a<�a<��a<S�a<��a<��a<2�a<��a<e�a<=�a<��a<��a<j�a<Q�a<T�a<�a<�a<�a<�a<�a<�a<�a<[a<_a<a<
a<�~a<�~a<�~a<�~a<�~a<�~a<�~a<�~a<�~a<a<!a<la<�  �  �a<�a<�a<.�a<J�a<^�a<��a<��a<�a<��a<�a<_�a<��a<΁a<�a<i�a<Ȃa<=�a<��a<�a<��a<�a<��a<�a<n�a<�a<M�a<��a<,�a<��a<�a<^�a<��a<>�a<��a<*�a<ԋa<J�a<�a<��a< �a<Îa<`�a<��a<|�a<�a<��a<�a<��a<��a<��a<ܓa<c�a<ؔa<L�a<֕a<Z�a<ؖa<h�a<�a<x�a<.�a<��a<6�a<��a<'�a<��a<�a<t�a<Ϝa<�a<V�a<��a<�a<�a<s�a<��a<�a<=�a<o�a<ӟa<�a<X�a<��a<�a<�a<J�a<w�a<��a<��a<��a<͡a<ѡa<��a<�a<�a<�a<	�a<"�a<9�a<h�a<{�a<��a<�a<�a<�a<�a<<�a<Z�a<P�a<V�a<L�a<5�a<'�a<�a<�a<עa<٢a<��a<��a<��a<��a<��a<��a<��a<��a<��a<w�a<f�a<8�a<��a<�a<��a<��a<.�a<�a<Ơa<��a<R�a<#�a<��a<ןa<Ɵa<��a<��a<u�a<N�a<,�a<�a<՞a<��a<^�a<�a<֝a<s�a<�a<Μa<a�a<�a<Ǜa<h�a<:�a<֚a<��a<Z�a<�a<��a<l�a<�a<��a<N�a<��a<E�a<͖a<<�a<̕a<�a<��a<�a<�a<�a<��a<�a<��a<+�a<��a<^�a<ޏa<v�a<�a<��a<&�a<��a<�a<��a<�a<b�a<�a<N�a<��a<M�a<��a<C�a<�a<e�a<�a<��a<X�a<�a<��a<P�a<�a<��a<�a<a<Y�a<�a<��a<�a<Ɓa<c�a<�a<πa<��a<[�a<@�a<�a<�a<�a<�a<�a<�a<�a<�a<ka<Ya<<a<a<a<�~a<�~a<�~a<�~a<�~a<�~a<�~a<�~a<"a<Oa<va<�  �  �a<�a<	�a<�a<`�a<|�a<��a<��a<��a<��a<�a<5�a<q�a<��a< �a<;�a<��a<�a<��a<�a<c�a<�a<j�a<�a<o�a<چa<R�a<��a<0�a<��a<�a<_�a<�a<T�a<ъa<i�a<̋a<��a<��a<��a<-�a<ǎa<_�a<�a<��a<��a<��a<�a<��a<��a<R�a<�a<6�a<Ĕa<0�a<��a<0�a<��a<Y�a<Ηa<��a< �a<��a<=�a<��a<M�a<��a<�a<o�a<̜a<$�a<a�a<ʝa<�a<M�a<n�a<ўa<�a<I�a<��a<ҟa<C�a<^�a<��a<�a<�a<N�a<l�a<��a<��a<áa<��a<��a<áa<��a<ѡa<ǡa<�a<�a<#�a<E�a<^�a<��a<��a<��a<�a<1�a<\�a<@�a<a�a<K�a<W�a<6�a<@�a<#�a<�a<�a<آa<�a<âa<עa<ˢa<��a<ʢa<��a<��a<��a<��a<Q�a<N�a<�a<١a<��a<B�a<1�a<ՠa<��a<i�a<"�a<�a<˟a<��a<��a<��a<v�a<A�a<T�a<�a<�a<֞a<��a<c�a<�a<۝a<q�a<K�a<Мa<��a<3�a<�a<��a<2�a<�a<��a<v�a<�a<��a<k�a<
�a<��a<*�a<�a<D�a<іa<7�a<��a<�a<q�a<��a<d�a<ؒa<]�a<�a<��a<��a<��a<0�a<Ϗa<~�a<�a<��a<�a<��a<�a<��a<�a<l�a<�a<S�a<�a<G�a<�a<i�a<�a<��a<�a<�a<^�a<�a<��a<U�a<��a<��a<<�a<��a<`�a<ɂa<n�a<�a<��a<O�a<�a<��a<b�a<E�a<�a<�a<�a<�a<�a<�a<�a<�a<xa<{a<Na<Ga<a<a<�~a<�~a<�~a<�~a<�~a<�~a<a<a</a<na<va<�  �  �a<�a<�a<+�a<M�a<]�a<t�a<��a<��a<��a<��a<�a<O�a<��a<�a<+�a<��a<��a<{�a<�a<^�a<�a<]�a<�a<h�a<�a<m�a<Їa<E�a<��a<�a<{�a<�a<c�a<��a<x�a<�a<��a<�a<��a<C�a<�a<o�a<	�a<��a<�a<��a<�a<z�a<�a<I�a<˓a<6�a<��a<�a<��a<&�a<��a<0�a<̗a<j�a<�a<��a<#�a<��a<8�a<��a<,�a<��a<ݜa<A�a<�a<ǝa<�a<`�a<��a<�a<'�a<Z�a<a<��a<@�a<��a<ʠa<��a<>�a<X�a<k�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<֡a<�a<�a<%�a<_�a<��a<��a<֢a<��a<�a<G�a<Q�a<u�a<i�a<a�a<\�a<F�a<0�a<+�a<�a<��a<��a<�a<ܢa<�a<ʢa<ʢa<Ţa<��a<��a<��a<c�a<;�a<��a<��a<��a<B�a<�a<Рa<��a<G�a<�a<�a<��a<��a<��a<z�a<a�a<;�a<6�a<�a<��a<Ξa<��a<~�a</�a<�a<��a<J�a<�a<��a<C�a<�a<��a<L�a<�a<Ța<u�a<'�a<�a<{�a<%�a<Ƙa<9�a<Ηa</�a<��a<$�a<��a<	�a<p�a<Гa<J�a<Вa<S�a<͑a<Y�a<��a<��a<#�a<��a<c�a<�a<��a<�a<��a<.�a<��a<$�a<��a<��a<z�a<��a<\�a< �a<��a<�a<��a<=�a<�a<��a<,�a<ƅa<s�a<��a<��a<"�a<��a<B�a<a<]�a<��a<��a<*�a<Հa<��a<\�a<&�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<la<Qa<>a< a<a<a<�~a<�~a<�~a<�~a<a<9a<Ca<na<�a<�  �  �a<�a<�a<1�a<H�a<h�a<��a<��a<��a<��a<��a<�a<<�a<��a<a<�a<v�a<�a<S�a<�a<m�a<ׄa<~�a<�a<h�a<�a<H�a<Ňa<>�a<��a<�a<��a<�a<��a<�a<f�a<,�a<��a<+�a<��a<V�a<�a<o�a<��a<w�a<�a<��a<�a<�a<ْa<_�a<��a<!�a<��a<�a<|�a<��a<��a<�a<��a<B�a<�a<��a<!�a<��a<+�a<��a<�a<u�a<ٜa<:�a<��a<ӝa<%�a<`�a<˞a<�a<?�a<��a<��a<�a<D�a<��a<àa<�a<�a<H�a<q�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<աa<�a<�a<D�a<e�a<��a<¢a<�a<)�a<<�a<Y�a<H�a<_�a<_�a<e�a<U�a<K�a<3�a<&�a<8�a<�a<�a<��a<�a<�a<բa<Ңa<��a<��a<m�a<h�a<6�a<�a<ۡa<u�a<Z�a<��a<��a<u�a<4�a<�a<Οa<��a<��a<x�a<R�a<T�a<K�a<�a<(�a<�a<Ξa<��a<Y�a<%�a<�a<��a<P�a<�a<��a<s�a<�a<��a<��a< �a<ؚa<��a<:�a<�a<|�a<�a<��a<H�a<��a<Q�a<��a<�a<��a<ޔa<\�a<��a<8�a<��a<)�a<��a<@�a<�a<m�a<5�a<��a<a�a<	�a<��a<�a<��a<�a<��a<�a<��a<�a<��a<��a<��a<��a<��a<=�a<��a<\�a<�a<��a<%�a<��a<O�a<�a<��a<�a<��a<-�a<̂a<\�a<сa<��a<�a<ʀa<y�a<G�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<ba<ba<Oa<Ha<.a<"a<a<a<$a<�~a<.a<*a<9a<da<ya<�a<�  �  �a< �a<�a<3�a<C�a<a�a<k�a<v�a<��a<��a<�a<�a<<�a<j�a<��a<�a<y�a<ނa<X�a<ԃa<F�a<Ʉa<X�a<�a<a�a<�a<l�a<�a<O�a<��a<)�a<��a<�a<��a<�a<��a<#�a<��a<B�a<ȍa<d�a<�a<��a<�a<��a<�a<��a<��a<V�a<Ēa<7�a<��a<�a<��a<�a<q�a<��a<��a<�a<��a<C�a<��a<l�a<��a<��a<�a<��a<*�a<��a<��a<I�a<��a<�a<5�a<g�a<a<��a<C�a<��a<ɟa<�a<R�a<��a<ՠa<�a<@�a<d�a<h�a<~�a<��a<~�a<}�a<��a<��a<��a<��a<��a<��a<��a<�a<�a<?�a<i�a<��a<��a<�a<�a<:�a<X�a<m�a<y�a<}�a<d�a<b�a<P�a<I�a<2�a<.�a<�a<�a<�a<��a<�a<�a<Ңa<Тa<��a<��a<k�a<1�a<�a<��a<l�a<0�a<��a<��a<k�a<4�a<�a<˟a<��a<��a<g�a<W�a<E�a<#�a<�a<�a<�a<Ǟa<��a<}�a<F�a<��a<��a<\�a<�a<��a<o�a< �a<a<��a<'�a<�a<��a<G�a<�a<��a</�a<��a<=�a<��a<3�a<��a<�a<w�a<�a<M�a<a<6�a<��a<!�a<��a<D�a<Րa<o�a<�a<��a<<�a<�a<|�a<�a<��a<6�a<��a<-�a<��a<�a<��a<�a<��a<�a<��a<4�a<��a<[�a<�a<��a<7�a<߅a<v�a<�a<��a<�a<��a<�a<��a<B�a<Ձa<k�a<�a<��a<r�a<0�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<�a<|a<ma<Ga<<a<'a<"a<a<a<a<'a<3a<Ma<ga<�a<�a<�  �  b~a<q~a<�~a<�~a<�~a<�~a<�~a<a<a< a<a<5a<va<�a<�a<;�a<��a<�a<��a<!�a<ւa<h�a<ʃa<��a<�a<��a<�a<v�a<��a<g�a<�a<^�a<�a<A�a<Éa<R�a<��a<|�a<�a<��a<2�a<��a<G�a<ώa<a�a<ڏa<c�a<��a<%�a<��a<ۑa<M�a<��a<��a<��a<�a<o�a<�a<��a<M�a<��a<��a<r�a<��a<{�a<0�a<��a<�a<��a<�a<C�a<��a<�a<<�a<��a<��a<�a<L�a<��a<��a<!�a<c�a<��a<џa<��a<+�a<K�a<k�a<��a<S�a<v�a<z�a<@�a<7�a<'�a<,�a<+�a<2�a<I�a<��a<��a<Рa<�a<R�a<��a<��a<��a<=�a<E�a<^�a<T�a<f�a<U�a<k�a<L�a<I�a</�a<�a<�a<�a<��a< �a<�a<�a<ơa<��a<��a<�a<S�a<1�a<�a<~�a<g�a<��a<��a<A�a<��a<˞a<o�a<J�a<$�a<�a<��a<��a<�a<	�a<�a<ȝa<�a<ŝa<��a<h�a<$�a<�a<��a<d�a<�a<כa<g�a<�a<Қa<b�a<E�a<�a<��a<K�a<Ԙa<��a<�a<��a<0�a<��a<�a<|�a<��a<)�a<��a<ܒa<3�a<��a<�a<��a<.�a<��a<[�a<
�a<��a<�a<
�a<��a<W�a<܌a<g�a<�a<i�a<�a<m�a<҉a<X�a<�a<9�a<·a<U�a<نa<��a<�a<��a<=�a<ׄa<h�a<�a<��a<*�a<��a<�a<��a<@�a<��a<�a<�a<Ga<�~a<�~a<W~a<G~a<~a<�}a<
~a<~a<2~a<~a<~a<0~a<~a<~a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<(~a<6~a<�  �  e~a<�~a<�~a<�~a<�~a<�~a<�~a<�~a<�~a<a<:a<Ga<la<�a<�a<N�a<��a<5�a<��a<2�a<��a<?�a<�a<r�a<�a<��a<�a<��a<��a<o�a<�a<I�a<��a<1�a<��a<6�a<Ċa<E�a<�a<��a<(�a<��a<V�a<�a<e�a<�a<G�a<��a<�a<j�a<��a<P�a<Ēa<�a<��a<�a<��a<�a<��a<n�a<�a<��a<0�a<�a<��a<�a<��a<$�a<��a< �a<L�a<��a<�a<*�a<[�a<��a<�a<8�a<{�a<��a<�a<^�a<��a<ݟa<�a<5�a<S�a<k�a<i�a<r�a<U�a<K�a<L�a<L�a<F�a<)�a<:�a<O�a<j�a<~�a<��a<��a<(�a<P�a<|�a<ʡa<��a<"�a<R�a<g�a<s�a<p�a<b�a<]�a<>�a<)�a<�a<�a<��a<�a<�a<ءa<ڡa<ޡa<Сa<��a<��a<��a<_�a<�a<ܠa<��a</�a<�a<��a<i�a<�a<��a<��a<b�a<8�a<�a<�a<�a<��a<�a<ڝa<�a<ϝa<��a<��a<n�a<>�a<��a<��a<`�a<�a<��a<V�a<
�a<��a<k�a<�a<әa<��a<A�a<�a<��a<(�a<��a<?�a<��a<�a<s�a<��a<.�a<��a<�a<H�a<��a<;�a<��a<7�a<��a<{�a<�a<��a<>�a<��a<��a<>�a<�a<m�a<��a<}�a<�a<g�a<ԉa<E�a<��a<:�a<��a<A�a<̆a<S�a<�a<��a<A�a<�a<��a<�a<��a<*�a<��a<+�a<��a<�a<��a<3�a<�a<Da<�~a<�~a<x~a<<~a<%~a<'~a<~a< ~a<�}a<~a<~a<~a<#~a<~a<~a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<~a<@~a<�  �  H~a<�~a<�~a<�~a<�~a<�~a<a<�~a<$a<a<a<Ka<ma<�a<�a<\�a<��a<8�a<��a<;�a<߂a<_�a<�a<j�a<�a<��a<��a<��a<�a<[�a<҇a<O�a<��a<:�a<��a<�a<ۊa<B�a<�a<��a<�a<��a<=�a<Վa<N�a<�a<C�a<ːa<B�a<��a<�a<0�a<��a<"�a<��a<�a<��a<"�a<��a<f�a<�a<ėa<Q�a<�a<��a<�a<��a<�a<��a<�a<=�a<��a<��a</�a<Y�a<ĝa<۝a<+�a<��a<��a<�a<N�a<��a<ğa<�a<)�a<K�a<u�a<^�a<��a<v�a<q�a<\�a<+�a<J�a<2�a<D�a<D�a<r�a<�a<��a<�a<�a<��a<��a<��a<�a<!�a<P�a<Q�a<n�a<S�a<Z�a<E�a<:�a<,�a<�a<�a<סa<�a<�a<ۡa<סa<ˡa<ơa<��a<��a<w�a<[�a<�a<۠a<��a<P�a<�a<��a<O�a<�a<a<��a<W�a<F�a<�a<�a<�a<�a<�a<��a<
�a<ȝa<ǝa<��a<]�a<4�a<ٜa<��a<P�a<	�a<��a<_�a<��a<��a<��a<�a<ԙa<��a<)�a<Ԙa<x�a<�a<��a<?�a<��a<$�a<��a<ߔa<]�a<w�a<��a<Z�a<��a<9�a<��a<;�a<Ώa<t�a<�a<ώa<_�a<�a<��a<6�a<�a<^�a<�a<i�a<ۊa<Q�a<͉a<J�a<��a<L�a<��a<4�a<چa<U�a<�a<��a<-�a<˄a<v�a<�a<��a<4�a<��a<H�a<��a<7�a<��a<�a<�a<Ma< a<�~a<�~a<=~a</~a<~a<�}a<6~a<~a<=~a<~a<~a<!~a<~a<	~a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<o}a<�}a<�}a<�}a<�}a<
~a<6~a<�  �  T~a<}~a<�~a<�~a<�~a<�~a<�~a<a<a<&a<Da<ya<�a<�a<�a<��a<�a<]�a<ǁa<H�a<؂a<n�a<��a<��a<�a<�a<�a<{�a<�a<T�a<ća<�a<��a<�a<��a<�a<��a<-�a<��a<h�a<
�a<��a<:�a<܎a<b�a<Ϗa<k�a<��a<2�a<��a<�a<m�a<Вa<K�a<��a<*�a<��a<Q�a<�a<��a< �a<��a<_�a<�a<y�a<9�a<��a<#�a<��a<�a<>�a<��a<˜a<��a<M�a<t�a<ҝa<�a<>�a<��a<�a<<�a<��a<ɟa<��a<9�a<J�a<f�a<��a<e�a<��a<o�a<_�a<]�a<j�a<g�a<m�a<j�a<��a<��a<�a<�a<;�a<t�a<��a<סa<��a<<�a<;�a<c�a<d�a<[�a<R�a<?�a<�a<�a<�a<֡a<ޡa<��a<��a<��a<��a<ša<��a<��a<��a<��a<G�a<,�a<�a<��a<d�a<�a<��a<t�a<=�a<��a<��a<}�a<k�a<R�a<>�a<�a<�a<�a<	�a<ߝa<�a<��a<��a<o�a<*�a<�a<��a<A�a<֛a<��a<�a<��a<��a<2�a<��a<��a<j�a<#�a<јa<u�a<#�a<��a<$�a<Öa<�a<��a<�a<Q�a<��a<�a<��a<�a<Q�a<ѐa<i�a<��a<��a<+�a<Ǝa<l�a<�a<��a<`�a<Ќa<m�a<��a<a�a<ۊa<M�a<��a<�a<��a<��a<��a<�a<��a<F�a<҅a<��a<*�a<Єa<j�a<�a<��a<%�a<��a<�a<��a<6�a<��a<D�a<�a<�a<*a<�~a<�~a<s~a<Z~a<2~a<'~a<$~a<'~a<~a<~a<0~a<~a<~a<�}a<�}a<�}a<�}a<�}a<u}a<^}a<\}a<v}a<p}a<w}a<�}a<�}a<~a<-~a<�  �  D~a<L~a<�~a<�~a<�~a<�~a<�~a<,a< a<aa<ca<|a<�a<�a<E�a<��a<�a<\�a<�a<z�a<�a<��a<��a<��a<��a<��a<��a<N�a<نa<(�a<��a<��a<��a<�a<j�a<��a<k�a<2�a<��a<O�a<��a<��a<'�a<��a<c�a<a<x�a<ǐa<R�a<��a<�a<��a<�a<Q�a<Γa<P�a<ڔa<c�a<��a<��a<S�a<җa<t�a<#�a<��a<M�a<��a<&�a<m�a<̛a<�a<]�a<��a<ڜa<L�a<\�a<��a<�a<3�a<��a<��a<.�a<X�a<��a<ԟa<�a<O�a<V�a<��a<z�a<��a<~�a<��a<��a<g�a<q�a<��a<��a<��a<Ša<�a< �a<t�a<��a<̡a<�a<�a<<�a</�a<^�a<2�a<K�a<"�a<!�a<�a<��a<�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<k�a<��a<D�a<)�a<��a<��a<��a<�a<��a<��a<A�a<�a<՞a<��a<��a<[�a<>�a<I�a<A�a<�a<)�a<��a<��a<��a<��a<\�a<��a<Мa<e�a<0�a<��a<��a<�a<��a<w�a<�a<��a<��a<Q�a<��a<��a<b�a<��a<��a<�a<Жa< �a<��a<�a<]�a<�a<!�a<��a<��a<w�a<��a<{�a<�a<��a<^�a<ގa<��a<6�a<��a<t�a<Ča<p�a<ϋa<I�a<��a< �a<��a<��a<��a<�a<z�a<��a<��a<?�a<��a<v�a<��a<��a<A�a<��a<��a<�a<؂a<3�a<ށa<D�a<�a<v�a<�a<�a<?a<�~a<�~a<�~a<_~a<M~a<a~a<0~a<F~a<3~a</~a<0~a< ~a<~a<�}a<�}a<�}a<�}a<q}a<e}a<g}a<:}a<S}a<L}a<{}a<�}a<�}a<�}a<�}a<�  �  5~a<]~a<�~a<�~a<�~a<�~a<a<&a<]a<Xa<ua<�a<�a<$�a<P�a<Ȁa<*�a<��a<�a<��a<�a<��a<�a<��a<�a<~�a<�a<^�a<Æa<�a<��a<�a<H�a<Ոa<?�a<��a<g�a<ڊa<x�a<�a<͌a<v�a<%�a<��a<E�a<ۏa<[�a<�a<Z�a<Ǒa<P�a<��a<�a<��a<��a<v�a<��a<��a<5�a<ʖa<8�a<�a<��a<(�a<��a<&�a<��a<�a<i�a<̛a<�a<K�a<��a<��a<�a<U�a<x�a<ĝa<$�a<P�a<��a<�a<F�a<��a<�a<�a<C�a<e�a<}�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ڠa<��a<1�a<@�a<`�a<��a<̡a<��a<�a<4�a<D�a<C�a<@�a<@�a<�a<�a<ءa<��a<��a<��a<t�a<��a<x�a<p�a<v�a<��a<|�a<��a<|�a<g�a<P�a<'�a<��a<��a<{�a<U�a<�a<��a<��a<6�a<�a<��a<��a<��a<��a<J�a<W�a<D�a< �a<�a<�a<��a<��a<H�a<�a<��a<U�a<�a<��a<:�a<��a<��a<6�a<�a<��a<`�a<!�a<�a<��a<`�a<��a<��a<1�a<��a<<�a<��a<�a<��a<ɓa<Y�a<̒a</�a<��a<�a<��a<G�a<؏a<D�a<�a<��a<;�a<̍a<M�a<܌a<V�a<ˋa<I�a<��a<�a<r�a<Ոa<A�a<݇a<>�a<͆a<u�a<�a<��a<J�a<�a<��a<P�a<�a<��a<$�a<��a<Q�a<؁a<j�a<�a<k�a<0�a<�a<oa<	a<�~a<�~a<�~a<n~a<L~a<o~a<F~a<C~a<:~a<'~a<~a<�}a<�}a<�}a<�}a<u}a<H}a<+}a<}a<)}a<}a<3}a<C}a<]}a<�}a<�}a<�}a<�  �  �}a<^~a<y~a<�~a<�~a<a<9a<,a<va<ya<�a<�a<�a<_�a<��a<�a<*�a<ˁa<!�a<��a<(�a<��a<9�a<��a<�a<r�a<�a<P�a<��a<�a<I�a<Շa<�a<��a<"�a<��a<9�a<��a<u�a<�a<a<N�a<�a<��a</�a<�a<V�a<��a<i�a<ˑa<s�a<��a<N�a<��a<*�a<��a<+�a<a<.�a<��a<^�a<2�a<��a<.�a<Йa<"�a<��a<��a<v�a<��a<�a<J�a<J�a<��a<��a<�a<O�a<��a<�a<�a<��a<Þa<M�a<g�a<˟a<�a<2�a<{�a<{�a<��a<��a<��a<Ѡa<��a<ڠa<��a<�a<ܠa<�a<�a<<�a<}�a<��a<ۡa<ѡa<�a<+�a<5�a<K�a<0�a<G�a<�a<�a<�a<��a<��a<`�a<��a<L�a<h�a<2�a<[�a<Z�a<W�a<t�a<Q�a<|�a<X�a<O�a</�a<�a<�a<��a<n�a<�a<�a<��a<H�a<@�a<�a<�a<��a<��a<x�a<u�a<[�a<)�a<7�a<�a<ѝa<��a<G�a<��a<��a<W�a<Ǜa<��a<�a<��a<v�a<�a<ߙa<d�a<\�a<�a<ۘa<y�a</�a<�a<�a<?�a<��a<T�a<��a<�a<��a<�a<��a<ʒa<Y�a<ґa<J�a<ڐa<@�a<	�a<i�a<=�a<��a<A�a<�a<I�a<�a<>�a<׋a< �a<��a<�a<7�a<ӈa<�a<��a<�a<��a<7�a<��a<��a<�a<�a<n�a<8�a<�a<|�a<;�a<��a<v�a<�a<|�a<%�a<��a<X�a<�a<�a<>a< a<�~a<�~a<�~a<p~a<�~a<K~a<e~a<F~a<(~a<~a<�}a<�}a<�}a<�}a<S}a<'}a< }a<�|a<}a<�|a<}a<�|a<H}a<m}a<�}a<�}a<�  �  �}a<6~a<r~a<�~a<�~a<a<<a<ia<za<�a<�a<�a<8�a<z�a<��a<%�a<n�a<Ձa<H�a<ʂa<A�a<Ƀa<.�a<��a<�a<s�a<؅a<2�a<��a<��a<#�a<��a<�a<v�a<�a<Y�a<�a<��a<K�a<Ƌa<��a<@�a<�a<��a<3�a<ԏa<j�a<��a<��a<��a<j�a<�a<T�a<Ɠa<e�a<Δa<R�a<��a<g�a<��a<��a<-�a<Ęa<S�a<Ùa<:�a<��a<��a<V�a<��a<؛a<*�a<&�a<��a<��a<�a<�a<n�a<��a<�a<g�a<��a<*�a<c�a<��a<�a<6�a<o�a<��a<��a<ڠa<ڠa<�a<ݠa<�a<�a<�a<�a<,�a<U�a<c�a<��a<��a<ۡa<�a<&�a</�a<>�a<:�a<,�a< �a<��a<�a<��a<��a<��a<\�a<H�a<�a<,�a<%�a<?�a<�a<6�a<[�a<K�a<U�a<P�a<D�a<3�a<�a<�a<��a<r�a<B�a<��a<��a<��a<[�a<�a<�a<֞a<��a<��a<��a<t�a<d�a<-�a<��a<ȝa<��a<9�a<�a<|�a<9�a<��a<R�a<�a<��a<B�a<ؙa<��a<m�a<2�a<Șa<��a<k�a<'�a<ߗa<��a<)�a<a<L�a<ܕa<O�a<��a<1�a<��a<��a<��a<��a<q�a<�a<y�a<�a<��a<8�a<юa<f�a<ߍa<a�a<ڌa<B�a<��a<�a<v�a<�a<�a<��a<�a<s�a<��a<w�a<�a<��a<X�a<�a<τa<j�a<%�a<ڃa<�a<.�a<˂a<i�a<�a<��a<5�a<Āa<^�a<�a<�a<fa<9a<a<�~a<�~a<�~a<�~a<�~a<n~a<J~a<2~a<~a<�}a<�}a<�}a<h}a<3}a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<+}a<3}a<v}a<�}a<�  �  �}a<~a<|~a<�~a<�~a<&a<,a<{a<�a<�a<�a<4�a<h�a<��a<��a<3�a<��a<
�a<s�a<�a<K�a<ԃa<$�a<��a<��a<��a<Ʌa<%�a<��a<��a<:�a<r�a<чa<A�a<��a<H�a<Ӊa<e�a< �a<ԋa<x�a<�a<�a<z�a<W�a<��a<z�a<��a<x�a<�a<}�a<�a<k�a<�a<q�a<��a<��a<�a<��a<�a<ϗa<A�a<Ԙa<O�a<ʙa<Q�a<��a< �a<5�a<��a<��a<�a<=�a<D�a<��a<��a<�a<D�a<��a<ڝa<4�a<��a<�a<V�a<��a<�a<M�a<U�a<��a<��a<ߠa<�a<��a<	�a<�a<>�a<�a<H�a<S�a<v�a<��a<��a<�a<�a<!�a<�a<F�a<?�a<4�a<C�a<�a<�a<��a<��a<��a<C�a<*�a<�a<�a<��a<��a<��a<�a<9�a<!�a<P�a<>�a<Z�a<C�a<*�a<'�a<٠a<Рa<~�a<i�a<�a<��a<��a<y�a<\�a<�a<$�a<�a<ʞa<��a<~�a<o�a<"�a<�a<��a<��a<*�a<Ӝa<y�a<��a<��a<,�a<Úa<f�a<�a<Ǚa<y�a<.�a<�a<֘a<��a<H�a<)�a<��a<��a<�a<Җa<V�a<ϕa<d�a<˔a<^�a<��a<S�a<��a<&�a<��a<�a<Ӑa<)�a<ڏa<L�a<�a<a�a<�a<x�a<Ìa<j�a<��a<�a<W�a<��a<*�a<_�a<χa<F�a<ʆa<N�a<ޅa<y�a<%�a<��a<��a<\�a<�a<��a<��a<�a<�a<f�a<�a<��a<I�a<��a<��a<Y�a<�a<�a<aa<4a<a<�~a<�~a<�~a<�~a<^~a<a~a<3~a<~a<�}a<�}a<�}a<7}a<'}a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<%}a<x}a<�}a<�  �  �}a<~a<_~a<�~a<�~a<.a<[a<�a<�a<�a<�a<@�a<f�a<��a<�a<T�a<��a<�a<��a<�a<v�a<�a<U�a<��a<�a<~�a<��a<�a<a�a<��a<�a<X�a<ʇa<0�a<��a<�a<��a<[�a<�a<��a<N�a<�a<̍a<d�a<;�a<яa<t�a<�a<��a<,�a<��a<%�a<��a< �a<�a< �a<��a<�a<a<;�a<ޗa<o�a<��a<k�a<�a<M�a<��a<	�a<�a<y�a<��a<ӛa<	�a<A�a<u�a<��a<ٜa<�a<|�a<ԝa<�a<��a<ߞa<8�a<��a<͟a<E�a<c�a<��a<ܠa<�a<�a<�a<#�a<!�a<6�a<=�a<k�a<v�a<x�a<��a<ɡa< �a<�a<6�a<E�a<U�a<;�a<>�a<&�a<�a<�a<��a<�a<W�a<B�a<�a<��a<ݠa<�a<�a<�a<�a<��a<�a<4�a<-�a<=�a<I�a<+�a</�a<�a<�a<��a<��a<5�a<�a<��a<��a<��a<>�a<�a<��a<�a<͞a<��a<�a<T�a<�a<��a<��a<�a<��a<Y�a<�a<��a<�a<��a<U�a<�a<��a<d�a<$�a<�a<��a<g�a<7�a<�a<��a<��a<&�a<͖a<w�a<��a<�a<��a<l�a<ϓa<W�a<��a<G�a<Ǒa<-�a<Ԑa<I�a<�a<z�a<�a<~�a<�a<t�a<ьa<S�a<�a<��a<E�a<��a<��a<\�a<Ňa<4�a<��a<(�a<ͅa<r�a<�a<̄a<��a<?�a<��a<��a<��a<"�a<�a<��a<,�a<сa<q�a<
�a<��a<Q�a<�a<�a<�a<6a<'a<�~a<�~a<�~a<�~a<�~a<p~a</~a<~a<�}a<�}a<n}a<+}a<�|a<�|a<�|a<�|a<�|a<u|a<�|a<�|a<�|a<}a<>}a<�}a<�  �  �}a<7~a<T~a<�~a<�~a<a<ha<a<�a<�a<-�a<_�a<��a<�a<�a<��a<ցa<H�a<��a<�a<}�a<݃a<[�a<��a<�a<\�a<��a<(�a<O�a<Æa<Ԇa<9�a<��a<��a<��a<��a<��a<'�a<�a<k�a<P�a<�a<Ǎa<��a<�a<�a<r�a<�a<��a<)�a<��a<8�a<ɓa<+�a<̔a<3�a<��a<g�a<̖a<r�a<�a<r�a<�a<u�a<�a<A�a<��a<ޚa<G�a<z�a<��a<ڛa<Λa<$�a<D�a<}�a<��a<�a<I�a<��a<�a<I�a<�a<)�a<��a<�a<�a<|�a<��a<٠a<�a<�a<"�a<?�a<R�a<Q�a<��a<i�a<��a<��a<ˡa<��a<�a< �a<(�a<O�a<C�a<G�a<?�a<�a<�a<ԡa<��a<n�a<,�a<�a<�a<ܠa<��a<Ġa<��a<Ƞa<ʠa<�a<$�a< �a<V�a<2�a<>�a<=�a<�a<�a<Ԡa<��a<��a<\�a<$�a<��a<ǟa<y�a<��a<>�a<*�a< �a<Ҟa<��a<y�a<Z�a<�a<ԝa<k�a<�a<֜a<G�a< �a<Q�a<�a<��a<!�a<ۙa<v�a<8�a<�a<͘a<m�a<i�a<6�a<�a<֗a<c�a<;�a<ʖa<i�a<�a<|�a<��a<�a<�a<c�a<��a<Z�a<ґa<�a<ސa<��a<��a<}�a< �a<��a<�a<h�a<�a<(�a<��a<��a<:�a<��a<��a<@�a<��a<�a<��a<�a<��a<L�a<��a<��a<��a<0�a<�a<��a<f�a<;�a<ӂa<��a<,�a<Ձa<v�a<%�a<рa<k�a<G�a<�a<�a<{a<>a<%a<�~a<�~a<�~a<�~a<^~a<;~a<~a<�}a<�}a<]}a<5}a<�|a<�|a<�|a<a|a<b|a<N|a<s|a<}|a<�|a<�|a<#}a<�}a<�  �  �}a<~a<W~a<�~a<�~a<3a<pa<�a<�a<�a<.�a<[�a<��a<�a<7�a<��a<فa<E�a<��a<$�a<��a<��a<a�a<��a<�a<^�a<��a<��a<1�a<��a<�a<M�a<��a<��a<��a< �a<��a<�a<�a<��a<:�a<�a<��a<u�a<�a<܏a<|�a<�a<��a<>�a<a<G�a<��a<,�a<��a<B�a<ƕa<W�a<Ζa<k�a<��a<��a<�a<��a<�a<O�a<��a<�a<4�a<V�a<y�a<��a<�a<'�a<9�a<z�a<��a<�a<D�a<��a<�a<h�a<��a<�a<}�a<۟a< �a<|�a<��a<�a<	�a<�a<;�a<@�a<Q�a<T�a<u�a<��a<��a<��a<ġa<�a<�a<2�a<F�a<Y�a<V�a<N�a<7�a<�a<��a<��a<��a<k�a<M�a<�a<�a<Πa<��a<��a<��a<Ġa<�a<�a<��a<��a<-�a<6�a<<�a<B�a<4�a<�a<�a<ɠa<��a<^�a<�a<��a<͟a<��a<u�a<A�a<'�a<�a<�a<��a<��a<`�a<�a<ԝa<m�a<�a<��a<)�a<ɛa<l�a<�a<��a<�a<ԙa<�a<2�a<�a<ɘa<��a<S�a<�a<ߗa<��a<n�a<1�a<Ԗa<t�a<�a<��a<�a<��a<��a<d�a<�a<i�a<�a<o�a<��a<y�a<�a<��a<�a<��a<�a<v�a<�a<1�a<��a<ӊa<�a<~�a<ۈa<B�a<��a<�a<��a<�a<��a<;�a<�a<��a<`�a<�a<�a<��a<i�a<;�a<�a<��a<F�a<��a<��a<'�a<πa<o�a<1�a<�a<�a<ta<7a< a<a<�~a<�~a<�~a<q~a<A~a<~a<�}a<�}a<<}a<	}a<�|a<�|a<�|a<]|a<T|a<V|a<d|a<{|a<�|a<�|a<*}a<f}a<�  �  �}a<�}a<a~a<�~a<�~a<'a<Pa<�a<�a<�a<C�a<��a<��a<�a<T�a<}�a<��a<b�a<��a<4�a<y�a<�a<E�a<��a<�a<~�a<��a<��a<n�a<��a<�a<"�a<��a<�a<_�a<��a<�a<�a<Ċa<~�a<1�a<�a<��a<W�a<<�a<׏a<s�a<�a<��a<1�a<��a<K�a<ϓa<o�a<ǔa<Y�a<��a<Y�a<�a<}�a<��a<��a<��a<r�a<�a<F�a<��a<�a<�a<n�a<��a<��a<�a<�a<2�a<o�a<��a<�a<E�a<��a<�a<f�a<��a<E�a<�a<ԟa<?�a<o�a<��a<͠a<��a<�a<I�a<D�a<i�a<��a<h�a<��a<��a<ša<��a<�a<#�a<,�a<A�a<>�a<P�a<F�a<B�a<)�a<ۡa<�a<��a<W�a<.�a<��a<�a<��a<��a<��a<��a<��a<��a<֠a<�a<3�a<�a<@�a<N�a<6�a<(�a<��a<�a< a<��a<r�a<K�a<�a<ʟa<��a<h�a<e�a<C�a<�a<��a<��a<��a<D�a<�a<ɝa<��a<�a<��a<f�a<ɛa<d�a<ܚa<r�a<'�a<��a<_�a<%�a<�a<��a<��a<J�a<F�a<��a<��a<��a<,�a<˖a<g�a<��a<��a<�a<��a<�a<��a<��a<��a<��a<q�a<!�a<��a<�a<��a<�a<��a<��a<m�a<܌a<K�a<{�a<�a<W�a<z�a<Ոa<$�a<��a<��a<]�a<�a<��a<#�a<܄a<��a<\�a<L�a<�a<��a<��a<.�a<�a<��a<7�a<Ӂa<��a<*�a<�a<��a<%�a<�a<�a<�a<qa<8a<a<�~a<�~a<�~a<k~a<9~a<~a<�}a<w}a<j}a<&}a<�|a<�|a<m|a<b|a<>|a<B|a<F|a<�|a<�|a<�|a<}a<x}a<�  �  �}a<~a<W~a<�~a<�~a<3a<pa<�a<�a<�a<.�a<[�a<��a<�a<7�a<��a<فa<E�a<��a<$�a<��a<��a<a�a<��a<�a<^�a<��a<��a<1�a<��a<�a<M�a<��a<��a<��a< �a<��a<�a<�a<��a<:�a<�a<��a<u�a<�a<܏a<|�a<�a<��a<>�a<a<G�a<��a<,�a<��a<B�a<ƕa<W�a<Ζa<k�a<��a<��a<�a<��a<�a<O�a<��a<�a<4�a<V�a<y�a<��a<�a<'�a<9�a<z�a<��a<�a<D�a<��a<�a<h�a<��a<�a<}�a<۟a< �a<|�a<��a<�a<	�a<�a<;�a<@�a<Q�a<T�a<u�a<��a<��a<��a<ġa<�a<�a<2�a<F�a<Y�a<V�a<N�a<7�a<�a<��a<��a<��a<k�a<M�a<�a<�a<Πa<��a<��a<��a<Ġa<�a<�a<��a<��a<-�a<6�a<<�a<B�a<4�a<�a<�a<ɠa<��a<^�a<�a<��a<͟a<��a<u�a<A�a<'�a<�a<�a<��a<��a<`�a<�a<ԝa<m�a<�a<��a<)�a<ɛa<l�a<�a<��a<�a<ԙa<�a<2�a<�a<ɘa<��a<S�a<�a<ߗa<��a<n�a<1�a<Ԗa<t�a<�a<��a<�a<��a<��a<d�a<�a<i�a<�a<o�a<��a<y�a<�a<��a<�a<��a<�a<v�a<�a<1�a<��a<ӊa<�a<~�a<ۈa<B�a<��a<�a<��a<�a<��a<;�a<�a<��a<`�a<�a<�a<��a<i�a<;�a<�a<��a<F�a<��a<��a<'�a<πa<o�a<1�a<�a<�a<ta<7a< a<a<�~a<�~a<�~a<q~a<A~a<~a<�}a<�}a<<}a<	}a<�|a<�|a<�|a<]|a<T|a<V|a<d|a<{|a<�|a<�|a<*}a<f}a<�  �  �}a<7~a<T~a<�~a<�~a<a<ha<a<�a<�a<-�a<_�a<��a<�a<�a<��a<ցa<H�a<��a<�a<}�a<݃a<[�a<��a<�a<\�a<��a<(�a<O�a<Æa<Ԇa<9�a<��a<��a<��a<��a<��a<'�a<�a<k�a<P�a<�a<Ǎa<��a<�a<�a<r�a<�a<��a<)�a<��a<8�a<ɓa<+�a<̔a<3�a<��a<g�a<̖a<r�a<�a<r�a<�a<u�a<�a<A�a<��a<ޚa<G�a<z�a<��a<ڛa<Λa<$�a<D�a<}�a<��a<�a<I�a<��a<�a<I�a<�a<)�a<��a<�a<�a<|�a<��a<٠a<�a<�a<"�a<?�a<R�a<Q�a<��a<i�a<��a<��a<ˡa<��a<�a< �a<(�a<O�a<C�a<G�a<?�a<�a<�a<ԡa<��a<n�a<,�a<�a<�a<ܠa<��a<Ġa<��a<Ƞa<ʠa<�a<$�a< �a<V�a<2�a<>�a<=�a<�a<�a<Ԡa<��a<��a<\�a<$�a<��a<ǟa<y�a<��a<>�a<*�a< �a<Ҟa<��a<y�a<Z�a<�a<ԝa<k�a<�a<֜a<G�a< �a<Q�a<�a<��a<!�a<ۙa<v�a<8�a<�a<͘a<m�a<i�a<6�a<�a<֗a<c�a<;�a<ʖa<i�a<�a<|�a<��a<�a<�a<c�a<��a<Z�a<ґa<�a<ސa<��a<��a<}�a< �a<��a<�a<h�a<�a<(�a<��a<��a<:�a<��a<��a<@�a<��a<�a<��a<�a<��a<L�a<��a<��a<��a<0�a<�a<��a<f�a<;�a<ӂa<��a<,�a<Ձa<v�a<%�a<рa<k�a<G�a<�a<�a<{a<>a<%a<�~a<�~a<�~a<�~a<^~a<;~a<~a<�}a<�}a<]}a<5}a<�|a<�|a<�|a<a|a<b|a<N|a<s|a<}|a<�|a<�|a<#}a<�}a<�  �  �}a<~a<_~a<�~a<�~a<.a<[a<�a<�a<�a<�a<@�a<f�a<��a<�a<T�a<��a<�a<��a<�a<v�a<�a<U�a<��a<�a<~�a<��a<�a<a�a<��a<�a<X�a<ʇa<0�a<��a<�a<��a<[�a<�a<��a<N�a<�a<̍a<d�a<;�a<яa<t�a<�a<��a<,�a<��a<%�a<��a< �a<�a< �a<��a<�a<a<;�a<ޗa<o�a<��a<k�a<�a<M�a<��a<	�a<�a<y�a<��a<ӛa<	�a<A�a<u�a<��a<ٜa<�a<|�a<ԝa<�a<��a<ߞa<8�a<��a<͟a<E�a<c�a<��a<ܠa<�a<�a<�a<#�a<!�a<6�a<=�a<k�a<v�a<x�a<��a<ɡa< �a<�a<6�a<E�a<U�a<;�a<>�a<&�a<�a<�a<��a<�a<W�a<B�a<�a<��a<ݠa<�a<�a<�a<�a<��a<�a<4�a<-�a<=�a<I�a<+�a</�a<�a<�a<��a<��a<5�a<�a<��a<��a<��a<>�a<�a<��a<�a<͞a<��a<�a<T�a<�a<��a<��a<�a<��a<Y�a<�a<��a<�a<��a<U�a<�a<��a<d�a<$�a<�a<��a<g�a<7�a<�a<��a<��a<&�a<͖a<w�a<��a<�a<��a<l�a<ϓa<W�a<��a<G�a<Ǒa<-�a<Ԑa<I�a<�a<z�a<�a<~�a<�a<t�a<ьa<S�a<�a<��a<E�a<��a<��a<\�a<Ňa<4�a<��a<(�a<ͅa<r�a<�a<̄a<��a<?�a<��a<��a<��a<"�a<�a<��a<,�a<сa<q�a<
�a<��a<Q�a<�a<�a<�a<6a<'a<�~a<�~a<�~a<�~a<�~a<p~a</~a<~a<�}a<�}a<n}a<+}a<�|a<�|a<�|a<�|a<�|a<u|a<�|a<�|a<�|a<}a<>}a<�}a<�  �  �}a<~a<|~a<�~a<�~a<&a<,a<{a<�a<�a<�a<4�a<h�a<��a<��a<3�a<��a<
�a<s�a<�a<K�a<ԃa<$�a<��a<��a<��a<Ʌa<%�a<��a<��a<:�a<r�a<чa<A�a<��a<H�a<Ӊa<e�a< �a<ԋa<x�a<�a<�a<z�a<W�a<��a<z�a<��a<x�a<�a<}�a<�a<k�a<�a<q�a<��a<��a<�a<��a<�a<ϗa<A�a<Ԙa<O�a<ʙa<Q�a<��a< �a<5�a<��a<��a<�a<=�a<D�a<��a<��a<�a<D�a<��a<ڝa<4�a<��a<�a<V�a<��a<�a<M�a<U�a<��a<��a<ߠa<�a<��a<	�a<�a<>�a<�a<H�a<S�a<v�a<��a<��a<�a<�a<!�a<�a<F�a<?�a<4�a<C�a<�a<�a<��a<��a<��a<C�a<*�a<�a<�a<��a<��a<��a<�a<9�a<!�a<P�a<>�a<Z�a<C�a<*�a<'�a<٠a<Рa<~�a<i�a<�a<��a<��a<y�a<\�a<�a<$�a<�a<ʞa<��a<~�a<o�a<"�a<�a<��a<��a<*�a<Ӝa<y�a<��a<��a<,�a<Úa<f�a<�a<Ǚa<y�a<.�a<�a<֘a<��a<H�a<)�a<��a<��a<�a<Җa<V�a<ϕa<d�a<˔a<^�a<��a<S�a<��a<&�a<��a<�a<Ӑa<)�a<ڏa<L�a<�a<a�a<�a<x�a<Ìa<j�a<��a<�a<W�a<��a<*�a<_�a<χa<F�a<ʆa<N�a<ޅa<y�a<%�a<��a<��a<\�a<�a<��a<��a<�a<�a<f�a<�a<��a<I�a<��a<��a<Y�a<�a<�a<aa<4a<a<�~a<�~a<�~a<�~a<^~a<a~a<3~a<~a<�}a<�}a<�}a<7}a<'}a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<%}a<x}a<�}a<�  �  �}a<6~a<r~a<�~a<�~a<a<<a<ia<za<�a<�a<�a<8�a<z�a<��a<%�a<n�a<Ձa<H�a<ʂa<A�a<Ƀa<.�a<��a<�a<s�a<؅a<2�a<��a<��a<#�a<��a<�a<v�a<�a<Y�a<�a<��a<K�a<Ƌa<��a<@�a<�a<��a<3�a<ԏa<j�a<��a<��a<��a<j�a<�a<T�a<Ɠa<e�a<Δa<R�a<��a<g�a<��a<��a<-�a<Ęa<S�a<Ùa<:�a<��a<��a<V�a<��a<؛a<*�a<&�a<��a<��a<�a<�a<n�a<��a<�a<g�a<��a<*�a<c�a<��a<�a<6�a<o�a<��a<��a<ڠa<ڠa<�a<ݠa<�a<�a<�a<�a<,�a<U�a<c�a<��a<��a<ۡa<�a<&�a</�a<>�a<:�a<,�a< �a<��a<�a<��a<��a<��a<\�a<H�a<�a<,�a<%�a<?�a<�a<6�a<[�a<K�a<U�a<P�a<D�a<3�a<�a<�a<��a<r�a<B�a<��a<��a<��a<[�a<�a<�a<֞a<��a<��a<��a<t�a<d�a<-�a<��a<ȝa<��a<9�a<�a<|�a<9�a<��a<R�a<�a<��a<B�a<ؙa<��a<m�a<2�a<Șa<��a<k�a<'�a<ߗa<��a<)�a<a<L�a<ܕa<O�a<��a<1�a<��a<��a<��a<��a<q�a<�a<y�a<�a<��a<8�a<юa<f�a<ߍa<a�a<ڌa<B�a<��a<�a<v�a<�a<�a<��a<�a<s�a<��a<w�a<�a<��a<X�a<�a<τa<j�a<%�a<ڃa<�a<.�a<˂a<i�a<�a<��a<5�a<Āa<^�a<�a<�a<fa<9a<a<�~a<�~a<�~a<�~a<�~a<n~a<J~a<2~a<~a<�}a<�}a<�}a<h}a<3}a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<+}a<3}a<v}a<�}a<�  �  �}a<^~a<y~a<�~a<�~a<a<9a<,a<va<ya<�a<�a<�a<_�a<��a<�a<*�a<ˁa<!�a<��a<(�a<��a<9�a<��a<�a<r�a<�a<P�a<��a<�a<I�a<Շa<�a<��a<"�a<��a<9�a<��a<u�a<�a<a<N�a<�a<��a</�a<�a<V�a<��a<i�a<ˑa<s�a<��a<N�a<��a<*�a<��a<+�a<a<.�a<��a<^�a<2�a<��a<.�a<Йa<"�a<��a<��a<v�a<��a<�a<J�a<J�a<��a<��a<�a<O�a<��a<�a<�a<��a<Þa<M�a<g�a<˟a<�a<2�a<{�a<{�a<��a<��a<��a<Ѡa<��a<ڠa<��a<�a<ܠa<�a<�a<<�a<}�a<��a<ۡa<ѡa<�a<+�a<5�a<K�a<0�a<G�a<�a<�a<�a<��a<��a<`�a<��a<L�a<h�a<2�a<[�a<Z�a<W�a<t�a<Q�a<|�a<X�a<O�a</�a<�a<�a<��a<n�a<�a<�a<��a<H�a<@�a<�a<�a<��a<��a<x�a<u�a<[�a<)�a<7�a<�a<ѝa<��a<G�a<��a<��a<W�a<Ǜa<��a<�a<��a<v�a<�a<ߙa<d�a<\�a<�a<ۘa<y�a</�a<�a<�a<?�a<��a<T�a<��a<�a<��a<�a<��a<ʒa<Y�a<ґa<J�a<ڐa<@�a<	�a<i�a<=�a<��a<A�a<�a<I�a<�a<>�a<׋a< �a<��a<�a<7�a<ӈa<�a<��a<�a<��a<7�a<��a<��a<�a<�a<n�a<8�a<�a<|�a<;�a<��a<v�a<�a<|�a<%�a<��a<X�a<�a<�a<>a< a<�~a<�~a<�~a<p~a<�~a<K~a<e~a<F~a<(~a<~a<�}a<�}a<�}a<�}a<S}a<'}a< }a<�|a<}a<�|a<}a<�|a<H}a<m}a<�}a<�}a<�  �  5~a<]~a<�~a<�~a<�~a<�~a<a<&a<]a<Xa<ua<�a<�a<$�a<P�a<Ȁa<*�a<��a<�a<��a<�a<��a<�a<��a<�a<~�a<�a<^�a<Æa<�a<��a<�a<H�a<Ոa<?�a<��a<g�a<ڊa<x�a<�a<͌a<v�a<%�a<��a<E�a<ۏa<[�a<�a<Z�a<Ǒa<P�a<��a<�a<��a<��a<v�a<��a<��a<5�a<ʖa<8�a<�a<��a<(�a<��a<&�a<��a<�a<i�a<̛a<�a<K�a<��a<��a<�a<U�a<x�a<ĝa<$�a<P�a<��a<�a<F�a<��a<�a<�a<C�a<e�a<}�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<ڠa<��a<1�a<@�a<`�a<��a<̡a<��a<�a<4�a<D�a<C�a<@�a<@�a<�a<�a<ءa<��a<��a<��a<t�a<��a<x�a<p�a<v�a<��a<|�a<��a<|�a<g�a<P�a<'�a<��a<��a<{�a<U�a<�a<��a<��a<6�a<�a<��a<��a<��a<��a<J�a<W�a<D�a< �a<�a<�a<��a<��a<H�a<�a<��a<U�a<�a<��a<:�a<��a<��a<6�a<�a<��a<`�a<!�a<�a<��a<`�a<��a<��a<1�a<��a<<�a<��a<�a<��a<ɓa<Y�a<̒a</�a<��a<�a<��a<G�a<؏a<D�a<�a<��a<;�a<̍a<M�a<܌a<V�a<ˋa<I�a<��a<�a<r�a<Ոa<A�a<݇a<>�a<͆a<u�a<�a<��a<J�a<�a<��a<P�a<�a<��a<$�a<��a<Q�a<؁a<j�a<�a<k�a<0�a<�a<oa<	a<�~a<�~a<�~a<n~a<L~a<o~a<F~a<C~a<:~a<'~a<~a<�}a<�}a<�}a<�}a<u}a<H}a<+}a<}a<)}a<}a<3}a<C}a<]}a<�}a<�}a<�}a<�  �  D~a<L~a<�~a<�~a<�~a<�~a<�~a<,a< a<aa<ca<|a<�a<�a<E�a<��a<�a<\�a<�a<z�a<�a<��a<��a<��a<��a<��a<��a<N�a<نa<(�a<��a<��a<��a<�a<j�a<��a<k�a<2�a<��a<O�a<��a<��a<'�a<��a<c�a<a<x�a<ǐa<R�a<��a<�a<��a<�a<Q�a<Γa<P�a<ڔa<c�a<��a<��a<S�a<җa<t�a<#�a<��a<M�a<��a<&�a<m�a<̛a<�a<]�a<��a<ڜa<L�a<\�a<��a<�a<3�a<��a<��a<.�a<X�a<��a<ԟa<�a<O�a<V�a<��a<z�a<��a<~�a<��a<��a<g�a<q�a<��a<��a<��a<Ša<�a< �a<t�a<��a<̡a<�a<�a<<�a</�a<^�a<2�a<K�a<"�a<!�a<�a<��a<�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<k�a<��a<D�a<)�a<��a<��a<��a<�a<��a<��a<A�a<�a<՞a<��a<��a<[�a<>�a<I�a<A�a<�a<)�a<��a<��a<��a<��a<\�a<��a<Мa<e�a<0�a<��a<��a<�a<��a<w�a<�a<��a<��a<Q�a<��a<��a<b�a<��a<��a<�a<Жa< �a<��a<�a<]�a<�a<!�a<��a<��a<w�a<��a<{�a<�a<��a<^�a<ގa<��a<6�a<��a<t�a<Ča<p�a<ϋa<I�a<��a< �a<��a<��a<��a<�a<z�a<��a<��a<?�a<��a<v�a<��a<��a<A�a<��a<��a<�a<؂a<3�a<ށa<D�a<�a<v�a<�a<�a<?a<�~a<�~a<�~a<_~a<M~a<a~a<0~a<F~a<3~a</~a<0~a< ~a<~a<�}a<�}a<�}a<�}a<q}a<e}a<g}a<:}a<S}a<L}a<{}a<�}a<�}a<�}a<�}a<�  �  T~a<}~a<�~a<�~a<�~a<�~a<�~a<a<a<&a<Da<ya<�a<�a<�a<��a<�a<]�a<ǁa<H�a<؂a<n�a<��a<��a<�a<�a<�a<{�a<�a<T�a<ća<�a<��a<�a<��a<�a<��a<-�a<��a<h�a<
�a<��a<:�a<܎a<b�a<Ϗa<k�a<��a<2�a<��a<�a<m�a<Вa<K�a<��a<*�a<��a<Q�a<�a<��a< �a<��a<_�a<�a<y�a<9�a<��a<#�a<��a<�a<>�a<��a<˜a<��a<M�a<t�a<ҝa<�a<>�a<��a<�a<<�a<��a<ɟa<��a<9�a<J�a<f�a<��a<e�a<��a<o�a<_�a<]�a<j�a<g�a<m�a<j�a<��a<��a<�a<�a<;�a<t�a<��a<סa<��a<<�a<;�a<c�a<d�a<[�a<R�a<?�a<�a<�a<�a<֡a<ޡa<��a<��a<��a<��a<ša<��a<��a<��a<��a<G�a<,�a<�a<��a<d�a<�a<��a<t�a<=�a<��a<��a<}�a<k�a<R�a<>�a<�a<�a<�a<	�a<ߝa<�a<��a<��a<o�a<*�a<�a<��a<A�a<֛a<��a<�a<��a<��a<2�a<��a<��a<j�a<#�a<јa<u�a<#�a<��a<$�a<Öa<�a<��a<�a<Q�a<��a<�a<��a<�a<Q�a<ѐa<i�a<��a<��a<+�a<Ǝa<l�a<�a<��a<`�a<Ќa<m�a<��a<a�a<ۊa<M�a<��a<�a<��a<��a<��a<�a<��a<F�a<҅a<��a<*�a<Єa<j�a<�a<��a<%�a<��a<�a<��a<6�a<��a<D�a<�a<�a<*a<�~a<�~a<s~a<Z~a<2~a<'~a<$~a<'~a<~a<~a<0~a<~a<~a<�}a<�}a<�}a<�}a<�}a<u}a<^}a<\}a<v}a<p}a<w}a<�}a<�}a<~a<-~a<�  �  H~a<�~a<�~a<�~a<�~a<�~a<a<�~a<$a<a<a<Ka<ma<�a<�a<\�a<��a<8�a<��a<;�a<߂a<_�a<�a<j�a<�a<��a<��a<��a<�a<[�a<҇a<O�a<��a<:�a<��a<�a<ۊa<B�a<�a<��a<�a<��a<=�a<Վa<N�a<�a<C�a<ːa<B�a<��a<�a<0�a<��a<"�a<��a<�a<��a<"�a<��a<f�a<�a<ėa<Q�a<�a<��a<�a<��a<�a<��a<�a<=�a<��a<��a</�a<Y�a<ĝa<۝a<+�a<��a<��a<�a<N�a<��a<ğa<�a<)�a<K�a<u�a<^�a<��a<v�a<q�a<\�a<+�a<J�a<2�a<D�a<D�a<r�a<�a<��a<�a<�a<��a<��a<��a<�a<!�a<P�a<Q�a<n�a<S�a<Z�a<E�a<:�a<,�a<�a<�a<סa<�a<�a<ۡa<סa<ˡa<ơa<��a<��a<w�a<[�a<�a<۠a<��a<P�a<�a<��a<O�a<�a<a<��a<W�a<F�a<�a<�a<�a<�a<�a<��a<
�a<ȝa<ǝa<��a<]�a<4�a<ٜa<��a<P�a<	�a<��a<_�a<��a<��a<��a<�a<ԙa<��a<)�a<Ԙa<x�a<�a<��a<?�a<��a<$�a<��a<ߔa<]�a<w�a<��a<Z�a<��a<9�a<��a<;�a<Ώa<t�a<�a<ώa<_�a<�a<��a<6�a<�a<^�a<�a<i�a<ۊa<Q�a<͉a<J�a<��a<L�a<��a<4�a<چa<U�a<�a<��a<-�a<˄a<v�a<�a<��a<4�a<��a<H�a<��a<7�a<��a<�a<�a<Ma< a<�~a<�~a<=~a</~a<~a<�}a<6~a<~a<=~a<~a<~a<!~a<~a<	~a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<o}a<�}a<�}a<�}a<�}a<
~a<6~a<�  �  e~a<�~a<�~a<�~a<�~a<�~a<�~a<�~a<�~a<a<:a<Ga<la<�a<�a<N�a<��a<5�a<��a<2�a<��a<?�a<�a<r�a<�a<��a<�a<��a<��a<o�a<�a<I�a<��a<1�a<��a<6�a<Ċa<E�a<�a<��a<(�a<��a<V�a<�a<e�a<�a<G�a<��a<�a<j�a<��a<P�a<Ēa<�a<��a<�a<��a<�a<��a<n�a<�a<��a<0�a<�a<��a<�a<��a<$�a<��a< �a<L�a<��a<�a<*�a<[�a<��a<�a<8�a<{�a<��a<�a<^�a<��a<ݟa<�a<5�a<S�a<k�a<i�a<r�a<U�a<K�a<L�a<L�a<F�a<)�a<:�a<O�a<j�a<~�a<��a<��a<(�a<P�a<|�a<ʡa<��a<"�a<R�a<g�a<s�a<p�a<b�a<]�a<>�a<)�a<�a<�a<��a<�a<�a<ءa<ڡa<ޡa<Сa<��a<��a<��a<_�a<�a<ܠa<��a</�a<�a<��a<i�a<�a<��a<��a<b�a<8�a<�a<�a<�a<��a<�a<ڝa<�a<ϝa<��a<��a<n�a<>�a<��a<��a<`�a<�a<��a<V�a<
�a<��a<k�a<�a<әa<��a<A�a<�a<��a<(�a<��a<?�a<��a<�a<s�a<��a<.�a<��a<�a<H�a<��a<;�a<��a<7�a<��a<{�a<�a<��a<>�a<��a<��a<>�a<�a<m�a<��a<}�a<�a<g�a<ԉa<E�a<��a<:�a<��a<A�a<̆a<S�a<�a<��a<A�a<�a<��a<�a<��a<*�a<��a<+�a<��a<�a<��a<3�a<�a<Da<�~a<�~a<x~a<<~a<%~a<'~a<~a< ~a<�}a<~a<~a<~a<#~a<~a<~a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<~a<@~a<�  �  �|a<}a<>}a<5}a<P}a<U}a<<}a<X}a<B}a<;}a</}a<Y}a<�}a<�}a<�}a<E~a<�~a<5a<�a<f�a< �a<��a<K�a<�a<��a<&�a<��a< �a<��a<��a<��a<�a<w�a<�a<O�a<ֈa<s�a<=�a<��a<Y�a<�a<m�a<$�a<��a<.�a<��a<�a<e�a<��a<0�a<e�a<��a<��a<��a<��a<Y�a<�a<��a<5�a<��a<}�a<;�a<�a<��a<S�a<�a<��a<)�a<��a<
�a<Q�a<��a<�a<�a<��a<��a<�a<1�a<��a<�a<��a<c�a<��a<�a<�a<G�a<V�a<Q�a<b�a<3�a<*�a<�a<�a<a<��a<��a<��a<��a<��a<��a<>�a<Q�a<��a<��a<f�a<��a<٠a<�a<&�a<^�a<\�a<u�a<C�a<G�a<?�a<�a<>�a<�a<ՠa<Рa<�a<Ӡa<Ԡa<ʠa<��a< a<��a<��a<5�a<�a<��a<N�a<�a<��a<4�a<��a<�a<7�a<�a<��a<��a<��a<s�a<t�a<��a<��a<��a<��a<��a<��a<��a<n�a<!�a<�a<��a<O�a<�a<��a<^�a<�a<��a<]�a<G�a<��a<��a<7�a<Ηa<��a<�a<��a<�a<��a<ܔa<,�a<��a<Òa<�a<?�a<̐a<"�a<w�a<��a<��a</�a<��a<f�a<�a<��a<��a<:�a<�a<��a<2�a<��a<@�a<��a<�a<��a<�a<��a<�a<X�a<�a<~�a<%�a<��a<M�a<уa<��a<�a<��a<>�a<��a<8�a<��a<�a<~a<�~a<C~a<�}a<g}a<�|a<�|a<_|a<R|a<H|a<|a<0|a<F|a<u|a<a|a<�|a<�|a<�|a<�|a<�|a<�|a<R|a<N|a<B|a<|a<K|a<
|a< |a<|a<a|a<T|a<}|a<�|a<�|a<�  �  �|a<	}a<)}a<8}a<G}a<S}a<b}a<D}a<@}a<I}a<[}a<b}a<}a<�}a<~a<g~a<�~a<Qa<�a<v�a<�a<��a<y�a<�a<��a<�a<��a<"�a<��a<�a<�a<�a<Q�a<·a<X�a<�a<d�a<�a<��a<:�a<�a<��a<�a<��a<"�a<��a<�a<��a<܏a< �a<|�a<Ԑa<0�a<��a<�a<s�a<��a<��a</�a<�a<��a<U�a<�a<̗a<�a<�a<��a<�a<��a<��a<_�a<��a<�a< �a<Y�a<��a<��a<:�a<p�a<��a<�a<Y�a<��a<�a<�a<3�a<D�a<X�a<R�a<f�a<7�a<�a<��a<�a<Ȟa<��a<��a<��a<�a<��a<7�a<��a<ßa<�a<P�a<��a<�a<
�a<3�a<M�a<Z�a<f�a<g�a<E�a<*�a<�a<�a<�a<�a<Ҡa<��a<��a<àa<Ơa<Πa<��a<��a<o�a<9�a<��a<��a<t�a<��a<��a<B�a<�a<��a<4�a<�a<˜a<��a<��a<��a<��a<��a<��a<��a<Ϝa<��a<��a<�a<]�a<"�a<��a<��a<K�a<�a<��a<=�a<��a<��a<M�a<��a<��a<x�a<3�a<�a<��a<�a<��a<�a<��a<��a<M�a<��a<ڒa<&�a<v�a<��a<�a<��a<�a<��a<)�a<܍a<��a<9�a<�a<��a<e�a<��a<��a<%�a<��a<2�a<��a<�a<��a<�a<T�a<ӆa<k�a<�a<g�a<��a<��a<D�a<�a<��a<�a<��a<,�a<��a<(�a<��a<�a<oa<�~a<k~a<�}a<f}a<}a<�|a<�|a<M|a<A|a<E|a<F|a<L|a<_|a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<v|a<L|a<-|a<
|a<�{a<|a<|a<|a<|a<9|a<m|a<�|a<�|a<�  �  �|a<}a<}a<K}a<]}a<A}a<]}a<D}a<k}a<P}a<i}a<t}a<�}a<�}a<~a<�~a<�~a<`a<�a<��a<2�a<��a<r�a<�a<��a<&�a<��a<'�a<��a<�a<Y�a<�a<Y�a<·a<=�a<��a<_�a<�a<��a<"�a<ċa<r�a<��a<��a<�a<��a<�a<v�a<ڏa<&�a<��a<ʐa<D�a<��a<�a<��a<	�a<��a<7�a<��a<��a<{�a<�a<ȗa<q�a<��a<��a<�a<��a<�a<J�a<��a<ța<?�a<O�a<��a<Ϝa<�a<r�a<��a<�a<5�a<��a<��a<�a<7�a<K�a<y�a<;�a<]�a<2�a<)�a<�a<�a<Ӟa<��a<ڞa<��a<��a<�a<C�a<��a<şa<1�a<O�a<��a<Ѡa<�a<I�a<@�a<d�a<@�a<O�a<'�a<#�a<*�a<�a<ݠa< a< a<��a<֠a< a<��a<��a<��a<��a<c�a<L�a<�a<��a<o�a<��a<ƞa<I�a<��a<��a<B�a<�a<Μa<Мa<��a<��a<��a<��a<��a<��a<ɜa<��a<��a<��a<]�a<(�a<̛a<��a<%�a<�a<��a<=�a<ڙa<��a<H�a<�a<ۘa<`�a<�a<ӗa<l�a<!�a<��a<5�a<�a<�a<J�a<��a<��a<�a<��a<Őa</�a<��a<�a<��a<0�a<�a<��a<_�a<�a<��a<X�a<�a<��a<%�a<��a<%�a<��a<�a<f�a<	�a<J�a<҆a<=�a<ąa<i�a<��a<��a<�a<Ճa<g�a<�a<��a<3�a<ցa<�a<��a<�a<�a<a<f~a<�}a<e}a</}a<�|a<�|a<]|a<M|a<W|a<G|a<w|a<^|a<�|a<�|a<�|a<�|a<�|a<�|a<]|a<]|a<-|a<&|a</|a<�{a<�{a<�{a<|a<|a<X|a<k|a<w|a<�|a<�  �  �|a<�|a<}a<1}a<b}a<h}a<`}a<e}a<j}a<l}a<�}a<�}a<�}a<�}a<0~a<�~a<a<�a<�a<��a<:�a<Ёa<o�a<�a<��a<�a<��a<�a<��a<�a<O�a<��a<!�a<��a<$�a<��a<4�a<ŉa<\�a<�a<��a<V�a<��a<��a<�a<��a<)�a<��a<�a<?�a<��a<�a<]�a<ˑa<4�a<��a<&�a<̓a<r�a<�a<��a<|�a<+�a<ڗa<��a<$�a<��a<�a<x�a<�a<0�a<�a<��a<�a<*�a<q�a<��a<��a<B�a<��a<ϝa<(�a<w�a<��a<�a<�a<7�a<[�a<l�a<_�a<I�a<9�a<$�a<�a<�a<�a<�a<�a<�a<=�a<}�a<��a<�a<+�a<n�a<��a<�a<&�a<)�a<6�a<B�a<J�a<.�a<�a<��a<٠a<Ǡa<��a<��a<��a<��a<��a<��a<��a<��a<��a<{�a<V�a<1�a<�a<ϟa<r�a<�a<Şa<e�a<�a<˝a<u�a<2�a<��a<��a<ɜa<Мa<��a<��a<ǜa<Ĝa<Ɯa<Ȝa<��a<s�a<D�a<	�a<ɛa<v�a<�a<��a<^�a<�a<��a<i�a<�a<Ϙa<��a<L�a<�a<��a<l�a<��a<��a<�a<��a<�a<Y�a<��a<��a<C�a<��a<�a<_�a<��a<7�a<Ўa<k�a<�a<��a<`�a<�a<��a<k�a<�a<��a<�a<��a<�a<��a<��a<V�a<��a<&�a<��a<#�a<��a<8�a<Ǆa<b�a<�a<��a<_�a<��a<��a<�a<��a<C�a<��a<!�a<�a<a<�~a<~a<�}a<D}a<�|a<�|a<�|a<�|a<n|a<e|a<q|a<}|a<�|a<�|a<�|a<�|a<~|a<r|a<f|a<=|a<%|a<|a<�{a<�{a<�{a<�{a<�{a<�{a<|a<@|a<o|a<�|a<�  �  �|a<�|a<5}a<>}a<?}a<i}a<p}a<�}a<t}a<�}a<�}a<�}a<�}a<'~a<z~a<�~a<'a<�a<7�a<ŀa<K�a<�a<v�a<�a<{�a<1�a<��a<�a<|�a<��a<=�a<��a<�a<h�a<�a<|�a<�a<��a<:�a<��a<��a<;�a<��a<g�a<>�a<��a<�a<��a<�a<g�a<��a<5�a<r�a<ڑa<N�a<�a<r�a<�a<��a<+�a<��a<��a<I�a<��a<~�a<%�a<��a<9�a<e�a<ߚa<�a<U�a<��a<ța<�a<,�a<��a<ɜa<�a<u�a<��a<�a<F�a<��a<�a<�a<_�a<?�a<u�a<_�a<y�a<M�a<?�a<9�a<�a<
�a<�a<6�a<H�a<W�a<��a<ȟa<"�a<8�a<��a<àa<�a<	�a<-�a<e�a<�a<G�a<�a<��a<ߠa<��a<��a<y�a<��a<c�a<e�a<n�a<t�a<��a<j�a<��a<X�a<{�a<?�a<��a<ϟa<��a<P�a<Оa<��a<4�a<؝a<��a<g�a<@�a<�a<�a<ܜa<�a<�a<؜a<��a<̜a<Ϝa<��a<��a<R�a<��a<śa<F�a<�a<��a<I�a<יa<��a<A�a<ژa<��a<`�a<5�a<�a<��a<e�a<ܖa<��a<
�a<��a<��a<u�a<ϓa<�a<��a<��a<�a<y�a<�a<��a<�a<��a<�a<�a<r�a<*�a<܌a<e�a<�a<��a<B�a<��a<�a<m�a<ˈa<D�a<��a<�a<_�a<��a<y�a<��a<��a<B�a<�a<��a<W�a<�a<��a<G�a<��a<K�a<��a<R�a<�a<.a<�~a<*~a<�}a<b}a<1}a<�|a<�|a<�|a<�|a<�|a<|a<�|a<�|a<�|a<�|a<�|a<�|a<O|a<d|a<|a<|a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<|a<W|a<q|a<�  �  �|a<�|a<}a<7}a<c}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<~a<a~a<�~a<a<`a<�a<^�a<�a<o�a<�a<��a</�a<��a<�a<t�a<�a<O�a<��a<
�a<]�a<ӆa<B�a<��a<8�a<̈a<l�a<#�a<��a<r�a<�a<ьa<\�a<�a<��a<1�a<��a<�a<v�a<ސa<B�a<��a<#�a<��a<�a<��a<3�a<ϔa<s�a<�a<��a<[�a<�a<��a<1�a<��a<�a<V�a<��a<��a<8�a<i�a<��a<֛a<�a<G�a<��a<ݜa<6�a<��a<��a<+�a<��a<Ҟa<��a<J�a<d�a<��a<t�a<��a<l�a<f�a<T�a<V�a<H�a<S�a<L�a<x�a<��a<ϟa<�a<5�a<k�a<��a<נa<�a<)�a<.�a<7�a<�a<�a<�a<ՠa<��a<��a<m�a<O�a<4�a<2�a<;�a<J�a<;�a<V�a<U�a<n�a<Q�a<K�a<8�a<�a<�a<��a<U�a<��a<��a<n�a<$�a<Нa<��a<W�a<P�a<&�a<�a<�a<�a<��a<��a<�a<�a<��a<��a<)�a<�a<��a<-�a<֚a<c�a<�a<��a<I�a<��a<��a<v�a<I�a<��a<×a<{�a<>�a<іa<��a<�a<��a<�a<��a<ޓa<<�a<��a<��a<[�a<��a<&�a<��a<7�a<Ȏa<c�a<��a<��a<=�a<�a<}�a<�a<��a<%�a<t�a<��a<M�a<��a<�a<s�a<цa<:�a<��a<6�a<Ԅa<x�a<�a<ʃa<q�a<,�a<ނa<q�a<1�a<��a<Z�a<ʀa<[�a<�a<Ua<�~a<n~a<�}a<�}a<G}a<}a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<|a<F|a<;|a<�{a<�{a<�{a<�{a<z{a<i{a<`{a<v{a<�{a<�{a<�{a<+|a<\|a<�  �  u|a<�|a<�|a<,}a<X}a<{}a<�}a<�}a<�}a<�}a<~a<#~a<J~a<�~a<�~a<Oa<�a<�a<��a<�a<��a<�a<��a< �a<��a<�a<p�a<ڄa<�a<��a<مa<9�a<��a<�a<��a<�a<��a<�a<��a<��a<X�a<��a<��a<l�a<�a<��a<&�a<��a<+�a<��a<�a<n�a<�a<D�a<Ӓa<E�a<ѓa<v�a<�a<��a<<�a<��a<v�a<�a<��a<)�a<��a<��a<b�a<��a<˚a<!�a<7�a<|�a<��a<�a<�a<W�a<��a<�a<Y�a<��a< �a<P�a<��a<��a<+�a<Y�a<{�a<��a<��a<��a<��a<�a<��a<i�a<��a<��a<��a<Οa<�a<0�a<c�a<��a<��a<��a<�a<�a<%�a<�a<�a<�a<ՠa<��a<w�a<]�a<�a<0�a<��a<�a<�a<�a<�a</�a<@�a<7�a<S�a<:�a<,�a<�a<�a<��a<e�a<7�a<�a<��a<I�a< �a<�a<��a<��a<L�a<Z�a<9�a<@�a<+�a<�a<	�a<՜a<��a<i�a<$�a<ۛa<d�a<"�a<��a<@�a<ʙa<t�a<!�a<Ƙa<��a<'�a<�a<ŗa<��a<V�a<�a<�a<|�a<�a<��a<+�a<��a<�a<}�a<��a<.�a<|�a<��a<c�a<�a<z�a<�a<��a<%�a<ލa<X�a<�a<��a<�a<��a<�a<��a<Չa<�a<��a<ԇa<E�a<��a<�a<��a<�a<��a<0�a<�a<��a<f�a<��a<a<q�a<�a<��a<Q�a<�a<p�a<�a<�a< a<�~a<~a<�}a<�}a<`}a<$}a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<d|a<M|a<|a<�{a<�{a<{{a<b{a<,{a<J{a<#{a<W{a<O{a<�{a<�{a<|a<G|a<�  �  e|a<�|a< }a<6}a<f}a<�}a<�}a<�}a<�}a<~a<)~a<h~a<�~a<�~a<a<na<�a<Y�a<��a<=�a<��a<I�a<��a<=�a<��a<�a<q�a<��a<	�a<X�a<��a<�a<j�a<ʆa<D�a<��a<a�a<��a<��a<[�a<�a<Ћa<��a<A�a<�a<��a<F�a<��a<L�a<��a<-�a<��a<�a<��a< �a<y�a<�a<��a<7�a<וa<q�a<�a<��a<A�a<��a<G�a<��a<�a<<�a<��a<��a<��a<
�a<@�a<n�a<��a<Λa<�a<n�a<˜a<)�a<}�a<ߝa<>�a<��a<�a<7�a<^�a<��a<��a<��a<��a<��a<��a<ɟa<��a<��a<ɟa<�a<�a<8�a<T�a<��a<��a<�a<�a<�a<2�a<0�a<+�a<��a<ܠa<��a<�a<P�a<'�a<��a<�a<��a<Οa<��a<ܟa<�a<��a<
�a<'�a<1�a<F�a<6�a<�a<�a<��a<��a<J�a<�a<��a<��a<I�a<�a<ӝa<��a<��a<��a<j�a<_�a<C�a<=�a< �a<�a<��a<v�a<%�a<��a<R�a<�a<w�a<�a<��a<9�a<��a<��a<K�a<	�a<ؗa<��a<k�a<1�a<�a<��a<��a<�a<��a<)�a<��a<)�a<��a<��a<W�a<Ƒa<+�a<��a<�a<��a<1�a<Ȏa<Z�a<�a<��a<$�a<��a<5�a<��a<�a<Z�a<��a<�a<V�a<��a<	�a<i�a<Յa<=�a<Ȅa<d�a<�a<��a<g�a<$�a<�a<��a<f�a<�a<��a<o�a<�a<��a<�a<�a<4a<�~a<m~a<~a<�}a<�}a<e}a<B}a<}a<}a<�|a<�|a<�|a<�|a<�|a<�|a<s|a<*|a<�{a<�{a<�{a<T{a<-{a<{a<{a<�za<{a<!{a<^{a<�{a<�{a<|a<�  �  a|a<�|a<�|a<}a<q}a<�}a<�}a<~a<~a<D~a<`~a<�~a<�~a<�~a<]a<�a<
�a<m�a<��a<h�a<сa<q�a<��a<h�a<��a<��a<R�a<��a<�a<%�a<��a<΅a<!�a<��a<�a<��a<�a<��a<m�a<D�a<�a<��a<��a<-�a<��a<�a<\�a<̏a<`�a<�a<G�a<ߑa<<�a<Βa<$�a<��a<G�a<��a<}�a<��a<��a<*�a<ʗa<\�a<��a<b�a<��a<��a<'�a<y�a<��a<��a<��a<��a<'�a<X�a<��a<��a<*�a<��a<�a<r�a<��a<1�a<��a<Оa<!�a<S�a<��a<��a<�a<ԟa<�a<�a<ޟa<��a<�a<�a<�a<8�a<m�a<��a< a<̠a<�a<�a<=�a<B�a<�a<�a<�a<נa<}�a<\�a<$�a<�a<��a<��a<��a<��a<��a<��a<��a<ޟa<ޟa<$�a<�a<,�a<�a<'�a<�a<ǟa<Ɵa<_�a<=�a<�a<��a<s�a<;�a<#�a<ܝa<ϝa<��a<��a<��a<^�a<f�a<
�a<�a<��a<Y�a<�a<��a<J�a<��a<h�a<ՙa<^�a<��a<��a<j�a<�a<Ǘa<��a<��a<C�a<�a<��a<��a<v�a<��a<וa<C�a<Дa<P�a<��a<1�a<��a<�a<O�a<ِa<X�a<��a<w�a<�a<��a<�a<��a<?�a<��a<P�a<~�a<�a<D�a<��a<�a<+�a<��a<Æa<"�a<��a<"�a<��a<!�a<Ńa<{�a<]�a<��a<؂a<��a<G�a<	�a<��a<��a<�a<��a<5�a<�a<oa<�~a<�~a<8~a<~a<�}a<�}a<w}a<K}a<D}a<}a<'}a<�|a<�|a<�|a<m|a<\|a<|a<�{a<�{a<c{a<({a<�za<�za<�za<�za<�za<�za<{a<`{a<�{a<�{a<�  �  /|a<�|a<�|a<5}a<^}a<�}a<�}a<~a<-~a<Z~a<�~a<�~a<�~a<9a<a<�a<0�a<��a<�a<��a<��a<t�a<ւa<6�a<��a<�a<S�a<��a<҄a<�a<X�a<��a<�a<q�a<܆a<W�a< �a<��a<^�a<�a<܊a<��a<c�a<0�a<�a<��a<2�a<Ϗa<k�a<�a<w�a<�a<[�a<ݒa<e�a<�a<v�a<�a<��a<�a<��a<V�a<ݗa<e�a<˘a<5�a<��a<��a<,�a<U�a<�a<��a<��a<�a<�a<=�a<g�a<��a<�a<w�a<Ϝa<,�a<��a<�a<p�a<֞a<1�a<X�a<��a<��a<�a<�a<�a<	�a<�a<�a<$�a<6�a<W�a<g�a<��a<��a<ՠa<��a<�a<%�a<*�a<%�a<)�a<�a<ؠa<��a<n�a<2�a<��a<֟a<��a<y�a<X�a<]�a<g�a<��a<��a<��a<ӟa<�a<
�a<*�a<6�a<�a<��a<�a<ȟa<��a<S�a<�a<՞a<��a<y�a<E�a<�a<��a<ϝa<��a<��a<��a<h�a<,�a<�a<��a<q�a<�a<��a<�a<��a<$�a<��a<V�a<ߘa<x�a<�a<�a<��a<��a<N�a<-�a<�a<Жa<��a<n�a<�a<��a<F�a<۔a<[�a<Փa<@�a<��a<�a<��a<�a<��a<�a<��a<	�a<��a<:�a<��a<H�a<��a<#�a<��a< �a<J�a<��a<҈a<�a<Z�a<��a<	�a<o�a<Մa<b�a<�a<��a<b�a<�a<�a<��a<}�a<M�a<�a<��a<a�a<�a<��a<S�a<�a<�a<a<�~a<y~a<1~a<�}a<�}a<�}a<p}a<W}a<>}a<*}a<}a<�|a<�|a<�|a<W|a<|a<�{a<~{a<8{a<�za<�za<�za<�za<�za<�za<�za<{a<={a<�{a<�{a<�  �  |a<�|a<�|a<5}a<w}a<�}a<�}a<
~a<N~a<b~a<�~a<�~a<a<Ua<�a<�a<Q�a<�a</�a<��a<�a<n�a<��a<A�a<��a<��a<8�a<��a<��a<�a<8�a<��a<܅a<:�a<ǆa<0�a<�a<g�a<2�a<�a<ъa<��a<N�a<)�a<��a<��a<D�a<�a<�a< �a<��a<��a<��a<
�a<��a<�a<��a<0�a<��a<p�a<Ζa<i�a<�a<r�a<�a<E�a<��a<řa<�a<B�a<h�a<��a<��a<Ța<՚a<�a<E�a<��a<ޛa<8�a<��a<�a<��a<�a<e�a<��a<�a<}�a<��a<�a<�a<�a<�a<!�a<Y�a<2�a<M�a<S�a<r�a<��a<��a<�a<ޠa<�a<�a<E�a<@�a<=�a<9�a<�a<ڠa<��a<i�a<�a<��a<��a<c�a<h�a<2�a<J�a<3�a<S�a<z�a<��a<џa<Οa<�a<��a<6�a<-�a<�a<�a<ğa<��a<[�a<E�a<�a<ɞa<��a<_�a<C�a<�a<#�a<�a<��a<��a<b�a<N�a<��a<͜a<]�a<�a<��a<��a<��a<�a<��a<�a<��a<c�a<��a<їa<q�a<X�a<(�a<#�a<�a<��a<��a<:�a<5�a<��a<h�a<�a<h�a<�a<O�a<�a<C�a<��a<"�a<��a<4�a<��a<`�a<��a<M�a<Սa<U�a<،a<4�a<��a<ϊa<:�a<y�a<��a<�a<2�a<��a<Ѕa<O�a<��a<K�a<ԃa<z�a<K�a<��a<�a<��a<r�a<6�a<��a<فa<n�a<6�a<��a<p�a<�a<�a<qa<�~a<�~a<N~a<~a<�}a<�}a<�}a<a}a<]}a<+}a<"}a<�|a<�|a<�|a<)|a<
|a<�{a<x{a<#{a<�za<�za<qza<�za<^za<�za<�za<�za<#{a<h{a<�{a<�  �  |a<�|a<�|a<}a<e}a<�}a<�}a</~a<f~a<�~a<�~a<�~a<a<ha<�a<�a<Y�a<��a<9�a<��a<0�a<��a<�a<L�a<��a<�a<G�a<��a<��a<�a<;�a<��a<҅a<)�a<��a<.�a<ʇa<g�a<'�a<�a<��a<s�a<S�a<4�a<؍a<��a<?�a<�a<~�a< �a<��a<�a<��a<�a<��a<.�a<��a</�a<��a<T�a<�a<��a<
�a<x�a<�a<D�a<��a<ޙa<*�a<H�a<T�a<z�a<��a<��a<Ϛa<�a<=�a<��a<˛a<0�a<��a<�a<}�a<�a<g�a<̞a<�a<e�a<��a<ԟa<�a<'�a<,�a<4�a<2�a<=�a<U�a<��a<��a<��a<��a<ݠa<�a</�a<C�a<=�a<B�a<0�a<�a<�a<ޠa<��a<F�a<�a<۟a<��a<a�a<G�a<-�a<.�a<)�a<A�a<o�a<��a<��a<Пa<�a<�a<�a<�a<�a<��a<�a<a<��a<D�a< �a<Ϟa<��a<��a<N�a<�a<��a<�a<ѝa<��a<��a<E�a<�a<��a<W�a<��a<��a<��a<�a<�a<��a<�a<��a<J�a<�a<��a<q�a<M�a<.�a<�a<Ԗa<��a<��a<R�a<�a<��a<c�a<�a<��a<�a<q�a<ڒa<F�a<��a<L�a<̐a<3�a<��a<D�a<֎a<e�a<�a<Z�a<ьa<2�a<��a<�a<H�a<~�a<��a<��a<;�a<��a<ʅa<5�a<��a<5�a<��a<r�a<7�a<��a<Âa<��a<s�a<D�a<��a<��a<u�a<)�a<܀a<��a<�a<�a<Ja<�~a<�~a<|~a<.~a<�}a<�}a<�}a<�}a<v}a<R}a<}a<�|a<�|a<�|a<8|a<|a<�{a<V{a<{a<�za<�za<nza<aza<Yza<rza<�za<�za<{a<^{a<�{a<�  �  !|a<^|a<�|a<$}a<d}a<�}a<�}a<6~a<B~a<�~a<�~a<�~a<Ta<da<�a<�a<��a<̀a<R�a<��a<�a<��a<�a<Z�a<��a<��a<6�a<c�a<ʄa<�a<#�a<U�a<ޅa<2�a<��a<�a<��a<f�a< �a<ɉa<��a<��a<B�a<�a<�a<��a<S�a<�a<��a< �a<��a<+�a<��a<?�a<��a<$�a<��a<<�a<��a<J�a<�a<z�a<�a<��a<��a<S�a<��a<�a<��a<0�a<e�a<a�a<w�a<��a<њa<��a<'�a<f�a<՛a<?�a<m�a<�a<i�a<��a<B�a<��a<!�a<P�a<��a<՟a<�a<�a<1�a<Q�a<7�a<��a<e�a<h�a<�a<àa<֠a<�a<�a<	�a<D�a<;�a<S�a<6�a<�a<��a<��a<��a<T�a<��a<��a<{�a<e�a<&�a<#�a<�a<+�a<2�a<F�a<{�a<��a<�a<�a<�a<$�a<�a<+�a<��a<�a<��a<��a<Q�a<�a<	�a<��a<s�a<Z�a<o�a<�a<�a<ԝa<��a<��a<G�a<�a<��a<a�a<�a<d�a<�a<t�a<�a<\�a<�a<��a<#�a<ܗa<��a<p�a<&�a<�a<�a<�a<��a<v�a<c�a<�a<͕a<y�a<��a<��a<�a<~�a<Ғa<x�a<ёa<B�a<��a<A�a<��a<;�a<�a<^�a<�a<h�a<ތa<A�a<��a<�a<�a<f�a<��a<ׇa<�a<R�a<̅a<&�a<��a<�a<̃a<��a<�a<܂a<��a<��a<O�a<*�a<	�a<��a<��a<*�a<�a<i�a< �a<�a<Oa<Aa<�~a<b~a<$~a<~a<�}a<�}a<�}a<O}a<S}a<}a<}a<�|a<�|a<F|a<�{a<�{a<c{a<{a<�za<�za<rza<@za<Pza<Sza<�za<�za<�za<Q{a<�{a<�  �  |a<�|a<�|a<}a<e}a<�}a<�}a</~a<f~a<�~a<�~a<�~a<a<ha<�a<�a<Y�a<��a<9�a<��a<0�a<��a<�a<L�a<��a<�a<G�a<��a<��a<�a<;�a<��a<҅a<)�a<��a<.�a<ʇa<g�a<'�a<�a<��a<s�a<S�a<4�a<؍a<��a<?�a<�a<~�a< �a<��a<�a<��a<�a<��a<.�a<��a</�a<��a<T�a<�a<��a<
�a<x�a<�a<D�a<��a<ޙa<*�a<H�a<T�a<z�a<��a<��a<Ϛa<�a<=�a<��a<˛a<0�a<��a<�a<}�a<�a<g�a<̞a<�a<e�a<��a<ԟa<�a<'�a<,�a<4�a<2�a<=�a<U�a<��a<��a<��a<��a<ݠa<�a</�a<C�a<=�a<B�a<0�a<�a<�a<ޠa<��a<F�a<�a<۟a<��a<a�a<G�a<-�a<.�a<)�a<A�a<o�a<��a<��a<Пa<�a<�a<�a<�a<�a<��a<�a<a<��a<D�a< �a<Ϟa<��a<��a<N�a<�a<��a<�a<ѝa<��a<��a<E�a<�a<��a<W�a<��a<��a<��a<�a<�a<��a<�a<��a<J�a<�a<��a<q�a<M�a<.�a<�a<Ԗa<��a<��a<R�a<�a<��a<c�a<�a<��a<�a<q�a<ڒa<F�a<��a<L�a<̐a<3�a<��a<D�a<֎a<e�a<�a<Z�a<ьa<2�a<��a<�a<H�a<~�a<��a<��a<;�a<��a<ʅa<5�a<��a<5�a<��a<r�a<7�a<��a<Âa<��a<s�a<D�a<��a<��a<u�a<)�a<܀a<��a<�a<�a<Ja<�~a<�~a<|~a<.~a<�}a<�}a<�}a<�}a<v}a<R}a<}a<�|a<�|a<�|a<8|a<|a<�{a<V{a<{a<�za<�za<nza<aza<Yza<rza<�za<�za<{a<^{a<�{a<�  �  |a<�|a<�|a<5}a<w}a<�}a<�}a<
~a<N~a<b~a<�~a<�~a<a<Ua<�a<�a<Q�a<�a</�a<��a<�a<n�a<��a<A�a<��a<��a<8�a<��a<��a<�a<8�a<��a<܅a<:�a<ǆa<0�a<�a<g�a<2�a<�a<ъa<��a<N�a<)�a<��a<��a<D�a<�a<�a< �a<��a<��a<��a<
�a<��a<�a<��a<0�a<��a<p�a<Ζa<i�a<�a<r�a<�a<E�a<��a<řa<�a<B�a<h�a<��a<��a<Ța<՚a<�a<E�a<��a<ޛa<8�a<��a<�a<��a<�a<e�a<��a<�a<}�a<��a<�a<�a<�a<�a<!�a<Y�a<2�a<M�a<S�a<r�a<��a<��a<�a<ޠa<�a<�a<E�a<@�a<=�a<9�a<�a<ڠa<��a<i�a<�a<��a<��a<c�a<h�a<2�a<J�a<3�a<S�a<z�a<��a<џa<Οa<�a<��a<6�a<-�a<�a<�a<ğa<��a<[�a<E�a<�a<ɞa<��a<_�a<C�a<�a<#�a<�a<��a<��a<b�a<N�a<��a<͜a<]�a<�a<��a<��a<��a<�a<��a<�a<��a<c�a<��a<їa<q�a<X�a<(�a<#�a<�a<��a<��a<:�a<5�a<��a<h�a<�a<h�a<�a<O�a<�a<C�a<��a<"�a<��a<4�a<��a<`�a<��a<M�a<Սa<U�a<،a<4�a<��a<ϊa<:�a<y�a<��a<�a<2�a<��a<Ѕa<O�a<��a<K�a<ԃa<z�a<K�a<��a<�a<��a<r�a<6�a<��a<فa<n�a<6�a<��a<p�a<�a<�a<qa<�~a<�~a<N~a<~a<�}a<�}a<�}a<a}a<]}a<+}a<"}a<�|a<�|a<�|a<)|a<
|a<�{a<x{a<#{a<�za<�za<qza<�za<^za<�za<�za<�za<#{a<h{a<�{a<�  �  /|a<�|a<�|a<5}a<^}a<�}a<�}a<~a<-~a<Z~a<�~a<�~a<�~a<9a<a<�a<0�a<��a<�a<��a<��a<t�a<ւa<6�a<��a<�a<S�a<��a<҄a<�a<X�a<��a<�a<q�a<܆a<W�a< �a<��a<^�a<�a<܊a<��a<c�a<0�a<�a<��a<2�a<Ϗa<k�a<�a<w�a<�a<[�a<ݒa<e�a<�a<v�a<�a<��a<�a<��a<V�a<ݗa<e�a<˘a<5�a<��a<��a<,�a<U�a<�a<��a<��a<�a<�a<=�a<g�a<��a<�a<w�a<Ϝa<,�a<��a<�a<p�a<֞a<1�a<X�a<��a<��a<�a<�a<�a<	�a<�a<�a<$�a<6�a<W�a<g�a<��a<��a<ՠa<��a<�a<%�a<*�a<%�a<)�a<�a<ؠa<��a<n�a<2�a<��a<֟a<��a<y�a<X�a<]�a<g�a<��a<��a<��a<ӟa<�a<
�a<*�a<6�a<�a<��a<�a<ȟa<��a<S�a<�a<՞a<��a<y�a<E�a<�a<��a<ϝa<��a<��a<��a<h�a<,�a<�a<��a<q�a<�a<��a<�a<��a<$�a<��a<V�a<ߘa<x�a<�a<�a<��a<��a<N�a<-�a<�a<Жa<��a<n�a<�a<��a<F�a<۔a<[�a<Փa<@�a<��a<�a<��a<�a<��a<�a<��a<	�a<��a<:�a<��a<H�a<��a<#�a<��a< �a<J�a<��a<҈a<�a<Z�a<��a<	�a<o�a<Մa<b�a<�a<��a<b�a<�a<�a<��a<}�a<M�a<�a<��a<a�a<�a<��a<S�a<�a<�a<a<�~a<y~a<1~a<�}a<�}a<�}a<p}a<W}a<>}a<*}a<}a<�|a<�|a<�|a<W|a<|a<�{a<~{a<8{a<�za<�za<�za<�za<�za<�za<�za<{a<={a<�{a<�{a<�  �  a|a<�|a<�|a<}a<q}a<�}a<�}a<~a<~a<D~a<`~a<�~a<�~a<�~a<]a<�a<
�a<m�a<��a<h�a<сa<q�a<��a<h�a<��a<��a<R�a<��a<�a<%�a<��a<΅a<!�a<��a<�a<��a<�a<��a<m�a<D�a<�a<��a<��a<-�a<��a<�a<\�a<̏a<`�a<�a<G�a<ߑa<<�a<Βa<$�a<��a<G�a<��a<}�a<��a<��a<*�a<ʗa<\�a<��a<b�a<��a<��a<'�a<y�a<��a<��a<��a<��a<'�a<X�a<��a<��a<*�a<��a<�a<r�a<��a<1�a<��a<Оa<!�a<S�a<��a<��a<�a<ԟa<�a<�a<ޟa<��a<�a<�a<�a<8�a<m�a<��a< a<̠a<�a<�a<=�a<B�a<�a<�a<�a<נa<}�a<\�a<$�a<�a<��a<��a<��a<��a<��a<��a<��a<ޟa<ޟa<$�a<�a<,�a<�a<'�a<�a<ǟa<Ɵa<_�a<=�a<�a<��a<s�a<;�a<#�a<ܝa<ϝa<��a<��a<��a<^�a<f�a<
�a<�a<��a<Y�a<�a<��a<J�a<��a<h�a<ՙa<^�a<��a<��a<j�a<�a<Ǘa<��a<��a<C�a<�a<��a<��a<v�a<��a<וa<C�a<Дa<P�a<��a<1�a<��a<�a<O�a<ِa<X�a<��a<w�a<�a<��a<�a<��a<?�a<��a<P�a<~�a<�a<D�a<��a<�a<+�a<��a<Æa<"�a<��a<"�a<��a<!�a<Ńa<{�a<]�a<��a<؂a<��a<G�a<	�a<��a<��a<�a<��a<5�a<�a<oa<�~a<�~a<8~a<~a<�}a<�}a<w}a<K}a<D}a<}a<'}a<�|a<�|a<�|a<m|a<\|a<|a<�{a<�{a<c{a<({a<�za<�za<�za<�za<�za<�za<{a<`{a<�{a<�{a<�  �  e|a<�|a< }a<6}a<f}a<�}a<�}a<�}a<�}a<~a<)~a<h~a<�~a<�~a<a<na<�a<Y�a<��a<=�a<��a<I�a<��a<=�a<��a<�a<q�a<��a<	�a<X�a<��a<�a<j�a<ʆa<D�a<��a<a�a<��a<��a<[�a<�a<Ћa<��a<A�a<�a<��a<F�a<��a<L�a<��a<-�a<��a<�a<��a< �a<y�a<�a<��a<7�a<וa<q�a<�a<��a<A�a<��a<G�a<��a<�a<<�a<��a<��a<��a<
�a<@�a<n�a<��a<Λa<�a<n�a<˜a<)�a<}�a<ߝa<>�a<��a<�a<7�a<^�a<��a<��a<��a<��a<��a<��a<ɟa<��a<��a<ɟa<�a<�a<8�a<T�a<��a<��a<�a<�a<�a<2�a<0�a<+�a<��a<ܠa<��a<�a<P�a<'�a<��a<�a<��a<Οa<��a<ܟa<�a<��a<
�a<'�a<1�a<F�a<6�a<�a<�a<��a<��a<J�a<�a<��a<��a<I�a<�a<ӝa<��a<��a<��a<j�a<_�a<C�a<=�a< �a<�a<��a<v�a<%�a<��a<R�a<�a<w�a<�a<��a<9�a<��a<��a<K�a<	�a<ؗa<��a<k�a<1�a<�a<��a<��a<�a<��a<)�a<��a<)�a<��a<��a<W�a<Ƒa<+�a<��a<�a<��a<1�a<Ȏa<Z�a<�a<��a<$�a<��a<5�a<��a<�a<Z�a<��a<�a<V�a<��a<	�a<i�a<Յa<=�a<Ȅa<d�a<�a<��a<g�a<$�a<�a<��a<f�a<�a<��a<o�a<�a<��a<�a<�a<4a<�~a<m~a<~a<�}a<�}a<e}a<B}a<}a<}a<�|a<�|a<�|a<�|a<�|a<�|a<s|a<*|a<�{a<�{a<�{a<T{a<-{a<{a<{a<�za<{a<!{a<^{a<�{a<�{a<|a<�  �  u|a<�|a<�|a<,}a<X}a<{}a<�}a<�}a<�}a<�}a<~a<#~a<J~a<�~a<�~a<Oa<�a<�a<��a<�a<��a<�a<��a< �a<��a<�a<p�a<ڄa<�a<��a<مa<9�a<��a<�a<��a<�a<��a<�a<��a<��a<X�a<��a<��a<l�a<�a<��a<&�a<��a<+�a<��a<�a<n�a<�a<D�a<Ӓa<E�a<ѓa<v�a<�a<��a<<�a<��a<v�a<�a<��a<)�a<��a<��a<b�a<��a<˚a<!�a<7�a<|�a<��a<�a<�a<W�a<��a<�a<Y�a<��a< �a<P�a<��a<��a<+�a<Y�a<{�a<��a<��a<��a<��a<�a<��a<i�a<��a<��a<��a<Οa<�a<0�a<c�a<��a<��a<��a<�a<�a<%�a<�a<�a<�a<ՠa<��a<w�a<]�a<�a<0�a<��a<�a<�a<�a<�a</�a<@�a<7�a<S�a<:�a<,�a<�a<�a<��a<e�a<7�a<�a<��a<I�a< �a<�a<��a<��a<L�a<Z�a<9�a<@�a<+�a<�a<	�a<՜a<��a<i�a<$�a<ۛa<d�a<"�a<��a<@�a<ʙa<t�a<!�a<Ƙa<��a<'�a<�a<ŗa<��a<V�a<�a<�a<|�a<�a<��a<+�a<��a<�a<}�a<��a<.�a<|�a<��a<c�a<�a<z�a<�a<��a<%�a<ލa<X�a<�a<��a<�a<��a<�a<��a<Չa<�a<��a<ԇa<E�a<��a<�a<��a<�a<��a<0�a<�a<��a<f�a<��a<a<q�a<�a<��a<Q�a<�a<p�a<�a<�a< a<�~a<~a<�}a<�}a<`}a<$}a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<d|a<M|a<|a<�{a<�{a<{{a<b{a<,{a<J{a<#{a<W{a<O{a<�{a<�{a<|a<G|a<�  �  �|a<�|a<}a<7}a<c}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<~a<a~a<�~a<a<`a<�a<^�a<�a<o�a<�a<��a</�a<��a<�a<t�a<�a<O�a<��a<
�a<]�a<ӆa<B�a<��a<8�a<̈a<l�a<#�a<��a<r�a<�a<ьa<\�a<�a<��a<1�a<��a<�a<v�a<ސa<B�a<��a<#�a<��a<�a<��a<3�a<ϔa<s�a<�a<��a<[�a<�a<��a<1�a<��a<�a<V�a<��a<��a<8�a<i�a<��a<֛a<�a<G�a<��a<ݜa<6�a<��a<��a<+�a<��a<Ҟa<��a<J�a<d�a<��a<t�a<��a<l�a<f�a<T�a<V�a<H�a<S�a<L�a<x�a<��a<ϟa<�a<5�a<k�a<��a<נa<�a<)�a<.�a<7�a<�a<�a<�a<ՠa<��a<��a<m�a<O�a<4�a<2�a<;�a<J�a<;�a<V�a<U�a<n�a<Q�a<K�a<8�a<�a<�a<��a<U�a<��a<��a<n�a<$�a<Нa<��a<W�a<P�a<&�a<�a<�a<�a<��a<��a<�a<�a<��a<��a<)�a<�a<��a<-�a<֚a<c�a<�a<��a<I�a<��a<��a<v�a<I�a<��a<×a<{�a<>�a<іa<��a<�a<��a<�a<��a<ޓa<<�a<��a<��a<[�a<��a<&�a<��a<7�a<Ȏa<c�a<��a<��a<=�a<�a<}�a<�a<��a<%�a<t�a<��a<M�a<��a<�a<s�a<цa<:�a<��a<6�a<Ԅa<x�a<�a<ʃa<q�a<,�a<ނa<q�a<1�a<��a<Z�a<ʀa<[�a<�a<Ua<�~a<n~a<�}a<�}a<G}a<}a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<|a<F|a<;|a<�{a<�{a<�{a<�{a<z{a<i{a<`{a<v{a<�{a<�{a<�{a<+|a<\|a<�  �  �|a<�|a<5}a<>}a<?}a<i}a<p}a<�}a<t}a<�}a<�}a<�}a<�}a<'~a<z~a<�~a<'a<�a<7�a<ŀa<K�a<�a<v�a<�a<{�a<1�a<��a<�a<|�a<��a<=�a<��a<�a<h�a<�a<|�a<�a<��a<:�a<��a<��a<;�a<��a<g�a<>�a<��a<�a<��a<�a<g�a<��a<5�a<r�a<ڑa<N�a<�a<r�a<�a<��a<+�a<��a<��a<I�a<��a<~�a<%�a<��a<9�a<e�a<ߚa<�a<U�a<��a<ța<�a<,�a<��a<ɜa<�a<u�a<��a<�a<F�a<��a<�a<�a<_�a<?�a<u�a<_�a<y�a<M�a<?�a<9�a<�a<
�a<�a<6�a<H�a<W�a<��a<ȟa<"�a<8�a<��a<àa<�a<	�a<-�a<e�a<�a<G�a<�a<��a<ߠa<��a<��a<y�a<��a<c�a<e�a<n�a<t�a<��a<j�a<��a<X�a<{�a<?�a<��a<ϟa<��a<P�a<Оa<��a<4�a<؝a<��a<g�a<@�a<�a<�a<ܜa<�a<�a<؜a<��a<̜a<Ϝa<��a<��a<R�a<��a<śa<F�a<�a<��a<I�a<יa<��a<A�a<ژa<��a<`�a<5�a<�a<��a<e�a<ܖa<��a<
�a<��a<��a<u�a<ϓa<�a<��a<��a<�a<y�a<�a<��a<�a<��a<�a<�a<r�a<*�a<܌a<e�a<�a<��a<B�a<��a<�a<m�a<ˈa<D�a<��a<�a<_�a<��a<y�a<��a<��a<B�a<�a<��a<W�a<�a<��a<G�a<��a<K�a<��a<R�a<�a<.a<�~a<*~a<�}a<b}a<1}a<�|a<�|a<�|a<�|a<�|a<|a<�|a<�|a<�|a<�|a<�|a<�|a<O|a<d|a<|a<|a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<|a<W|a<q|a<�  �  �|a<�|a<}a<1}a<b}a<h}a<`}a<e}a<j}a<l}a<�}a<�}a<�}a<�}a<0~a<�~a<a<�a<�a<��a<:�a<Ёa<o�a<�a<��a<�a<��a<�a<��a<�a<O�a<��a<!�a<��a<$�a<��a<4�a<ŉa<\�a<�a<��a<V�a<��a<��a<�a<��a<)�a<��a<�a<?�a<��a<�a<]�a<ˑa<4�a<��a<&�a<̓a<r�a<�a<��a<|�a<+�a<ڗa<��a<$�a<��a<�a<x�a<�a<0�a<�a<��a<�a<*�a<q�a<��a<��a<B�a<��a<ϝa<(�a<w�a<��a<�a<�a<7�a<[�a<l�a<_�a<I�a<9�a<$�a<�a<�a<�a<�a<�a<�a<=�a<}�a<��a<�a<+�a<n�a<��a<�a<&�a<)�a<6�a<B�a<J�a<.�a<�a<��a<٠a<Ǡa<��a<��a<��a<��a<��a<��a<��a<��a<��a<{�a<V�a<1�a<�a<ϟa<r�a<�a<Şa<e�a<�a<˝a<u�a<2�a<��a<��a<ɜa<Мa<��a<��a<ǜa<Ĝa<Ɯa<Ȝa<��a<s�a<D�a<	�a<ɛa<v�a<�a<��a<^�a<�a<��a<i�a<�a<Ϙa<��a<L�a<�a<��a<l�a<��a<��a<�a<��a<�a<Y�a<��a<��a<C�a<��a<�a<_�a<��a<7�a<Ўa<k�a<�a<��a<`�a<�a<��a<k�a<�a<��a<�a<��a<�a<��a<��a<V�a<��a<&�a<��a<#�a<��a<8�a<Ǆa<b�a<�a<��a<_�a<��a<��a<�a<��a<C�a<��a<!�a<�a<a<�~a<~a<�}a<D}a<�|a<�|a<�|a<�|a<n|a<e|a<q|a<}|a<�|a<�|a<�|a<�|a<~|a<r|a<f|a<=|a<%|a<|a<�{a<�{a<�{a<�{a<�{a<�{a<|a<@|a<o|a<�|a<�  �  �|a<}a<}a<K}a<]}a<A}a<]}a<D}a<k}a<P}a<i}a<t}a<�}a<�}a<~a<�~a<�~a<`a<�a<��a<2�a<��a<r�a<�a<��a<&�a<��a<'�a<��a<�a<Y�a<�a<Y�a<·a<=�a<��a<_�a<�a<��a<"�a<ċa<r�a<��a<��a<�a<��a<�a<v�a<ڏa<&�a<��a<ʐa<D�a<��a<�a<��a<	�a<��a<7�a<��a<��a<{�a<�a<ȗa<q�a<��a<��a<�a<��a<�a<J�a<��a<ța<?�a<O�a<��a<Ϝa<�a<r�a<��a<�a<5�a<��a<��a<�a<7�a<K�a<y�a<;�a<]�a<2�a<)�a<�a<�a<Ӟa<��a<ڞa<��a<��a<�a<C�a<��a<şa<1�a<O�a<��a<Ѡa<�a<I�a<@�a<d�a<@�a<O�a<'�a<#�a<*�a<�a<ݠa< a< a<��a<֠a< a<��a<��a<��a<��a<c�a<L�a<�a<��a<o�a<��a<ƞa<I�a<��a<��a<B�a<�a<Μa<Мa<��a<��a<��a<��a<��a<��a<ɜa<��a<��a<��a<]�a<(�a<̛a<��a<%�a<�a<��a<=�a<ڙa<��a<H�a<�a<ۘa<`�a<�a<ӗa<l�a<!�a<��a<5�a<�a<�a<J�a<��a<��a<�a<��a<Őa</�a<��a<�a<��a<0�a<�a<��a<_�a<�a<��a<X�a<�a<��a<%�a<��a<%�a<��a<�a<f�a<	�a<J�a<҆a<=�a<ąa<i�a<��a<��a<�a<Ճa<g�a<�a<��a<3�a<ցa<�a<��a<�a<�a<a<f~a<�}a<e}a</}a<�|a<�|a<]|a<M|a<W|a<G|a<w|a<^|a<�|a<�|a<�|a<�|a<�|a<�|a<]|a<]|a<-|a<&|a</|a<�{a<�{a<�{a<|a<|a<X|a<k|a<w|a<�|a<�  �  �|a<	}a<)}a<8}a<G}a<S}a<b}a<D}a<@}a<I}a<[}a<b}a<}a<�}a<~a<g~a<�~a<Qa<�a<v�a<�a<��a<y�a<�a<��a<�a<��a<"�a<��a<�a<�a<�a<Q�a<·a<X�a<�a<d�a<�a<��a<:�a<�a<��a<�a<��a<"�a<��a<�a<��a<܏a< �a<|�a<Ԑa<0�a<��a<�a<s�a<��a<��a</�a<�a<��a<U�a<�a<̗a<�a<�a<��a<�a<��a<��a<_�a<��a<�a< �a<Y�a<��a<��a<:�a<p�a<��a<�a<Y�a<��a<�a<�a<3�a<D�a<X�a<R�a<f�a<7�a<�a<��a<�a<Ȟa<��a<��a<��a<�a<��a<7�a<��a<ßa<�a<P�a<��a<�a<
�a<3�a<M�a<Z�a<f�a<g�a<E�a<*�a<�a<�a<�a<�a<Ҡa<��a<��a<àa<Ơa<Πa<��a<��a<o�a<9�a<��a<��a<t�a<��a<��a<B�a<�a<��a<4�a<�a<˜a<��a<��a<��a<��a<��a<��a<��a<Ϝa<��a<��a<�a<]�a<"�a<��a<��a<K�a<�a<��a<=�a<��a<��a<M�a<��a<��a<x�a<3�a<�a<��a<�a<��a<�a<��a<��a<M�a<��a<ڒa<&�a<v�a<��a<�a<��a<�a<��a<)�a<܍a<��a<9�a<�a<��a<e�a<��a<��a<%�a<��a<2�a<��a<�a<��a<�a<T�a<ӆa<k�a<�a<g�a<��a<��a<D�a<�a<��a<�a<��a<,�a<��a<(�a<��a<�a<oa<�~a<k~a<�}a<f}a<}a<�|a<�|a<M|a<A|a<E|a<F|a<L|a<_|a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<v|a<L|a<-|a<
|a<�{a<|a<|a<|a<|a<9|a<m|a<�|a<�|a<�  �  �{a<�{a<�{a<�{a<�{a<�{a<|{a<�{a<b{a<u{a<@{a<T{a<`{a<�{a<|a< |a<�|a<6}a<�}a<�~a<Ja<�a<��a<u�a<�a<͂a<i�a<ڃa<_�a<��a<F�a<��a<�a<��a<�a<m�a<��a<ψa<2�a<#�a<{�a<=�a<��a<p�a<)�a<_�a<͍a<�a<O�a<��a<�a<J�a<^�a<�a<�a<��a<T�a<��a<��a<-�a<'�a<�a<��a<k�a<)�a<��a<��a<`�a<��a<%�a<j�a<��a<"�a<�a<��a<��a<Λa<�a<s�a<Мa<��a<��a<{�a<��a<!�a<K�a<e�a<@�a<6�a<��a<�a<��a<��a<V�a<�a<�a<ڜa<,�a<�a<9�a<��a<˝a<[�a<��a<��a<5�a<��a<�a<'�a<t�a<\�a<s�a<;�a<3�a<@�a<�a<�a<��a<��a<��a<ڟa<��a<ǟa<��a<��a<şa<��a<��a<2�a<ߞa<{�a<��a<��a<&�a<՜a<8�a<ߛa<z�a<+�a<1�a<ʚa<�a<Ԛa<��a<*�a<5�a<O�a<[�a<��a<��a<��a<u�a<1�a<��a<t�a<e�a<ޙa<��a<A�a<˘a<|�a<1�a<�a<��a<��a<�a<ؖa<��a<�a<ѕa<�a<l�a<��a<ڒa<,�a<X�a<��a<��a<�a<=�a<̍a<U�a<��a<��a<��a<�a<��a<e�a<�a<׊a<��a<H�a<%�a<|�a<�a<o�a<��a<j�a<��a<+�a<q�a<߄a<a�a<
�a<��a<1�a<�a<]�a<8�a<ȁa<\�a<�a<5�a<�a<�~a<Q~a<�}a<}a<m|a<�{a<_{a<�za<�za<Qza<"za<2za<!za<oza<nza<�za<�za<�za<{a<{a<K{a<{a<{a<�za<�za<�za<�za<�za<jza<oza<zza<�za<�za<{a<${a</{a<�  �  r{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<i{a<U{a<G{a<U{a<s{a<�{a<�{a<5|a<�|a<G}a<�}a<�~a<Ra<�a<܀a<��a<"�a<��a<?�a<��a<D�a<��a<$�a<��a<��a<e�a<��a<��a<�a<��a<B�a<��a<��a<O�a<Ƌa<Y�a<�a<Y�a<׍a<2�a<~�a<��a<�a<:�a<w�a<֏a<3�a<��a<%�a<Бa<��a<G�a<�a<ޔa<��a<��a<Y�a<�a<��a<�a<��a<�a<m�a<��a<�a<!�a<b�a<��a<��a<0�a<b�a<��a<�a<Y�a<��a<�a<��a<(�a<3�a<G�a<C�a<,�a<��a<��a<y�a<T�a<%�a<�a<�a<�a<�a<T�a<��a<ڝa<=�a<��a<�a<m�a<��a<��a<�a<9�a<B�a<M�a<^�a<6�a<%�a<��a<ݟa<ɟa<��a<��a<��a<��a<��a<��a<��a<��a<u�a<X�a< �a<�a<��a<3�a<��a<,�a<��a<?�a<��a<��a<2�a<��a<ߚa<�a<�a<��a<�a<<�a<e�a<��a<��a<��a<c�a<K�a<	�a<�a<��a<C�a<�a<��a<"�a<��a<��a<3�a<�a<��a<s�a<#�a<�a<i�a< �a<��a<��a<v�a<ɓa<
�a<7�a<S�a<��a<Ïa<�a<Z�a<��a<&�a<��a<t�a<�a<�a<��a<r�a<E�a<�a<��a<D�a<��a<d�a<܈a<r�a<ˇa<7�a<��a<�a<m�a<
�a<��a<��a<��a<7�a<��a<��a<$�a<��a<9�a<��a<<�a<�a<a<j~a<�}a<�|a<k|a<�{a<a{a<�za<za<Pza<=za<.za<0za<Qza<kza<�za<�za< {a<{a<{a<{a<{a<�za<�za<�za<�za<�za<yza<rza<�za<�za<�za<�za<�za<{a<X{a<�  �  S{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<e{a<p{a<d{a<�{a<�{a<�{a<z|a<�|a<e}a<~a<�~a<qa<�a<̀a<_�a<-�a<��a<[�a<σa<%�a<��a<�a<}�a<څa<G�a<��a<B�a<�a<�a<M�a<��a<��a<8�a<��a<��a<�a<w�a<��a<�a<f�a<��a<�a<B�a<��a<Ϗa<n�a<אa<X�a<�a<��a<m�a<#�a<��a<ȕa<|�a<?�a<�a<��a<�a<��a<�a<S�a<��a<��a<,�a<:�a<|�a<��a<�a<F�a<��a<��a<�a<��a<ĝa<�a<N�a<8�a<\�a<"�a<�a<�a<ԝa<��a<f�a<F�a<�a<7�a<�a<Q�a<w�a<��a<�a<I�a<��a<�a<[�a<��a<�a<1�a<C�a<u�a<4�a<K�a<�a<��a<�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<g�a<3�a<ߞa<q�a<%�a<��a<V�a<Ŝa<h�a<�a<��a<o�a<�a<$�a<�a<�a<�a<&�a<\�a<V�a<~�a<n�a<��a<m�a<h�a<'�a<Ěa<��a<
�a<ԙa<g�a<�a<��a<Q�a<�a<Ηa<��a<:�a<�a<Җa<Z�a<3�a<��a<�a<X�a<��a<�a<:�a<w�a<��a<�a<	�a<��a<�a<Z�a<�a<j�a<>�a<�a<��a<{�a<+�a<�a<��a<g�a<߉a<��a<وa<X�a<̇a<��a<��a<܅a<S�a<��a<@�a<܃a<v�a</�a<��a<��a<�a<��a<`�a<��a<R�a<�a<a<T~a<�}a<}a<||a<�{a<\{a<!{a<�za<�za<_za<7za<^za<^za<�za<�za<�za<�za< {a<&{a<{a<4{a<�za<�za<�za<�za<�za<[za<Uza<Aza<bza<xza<�za<�za<�za<L{a<�  �  L{a<}{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<5|a<�|a<�|a<�}a<$~a<�~a<�a</�a<��a<��a<)�a<��a<(�a<��a<�a<��a<�a<L�a<��a<9�a<��a<�a<ׇa<Y�a<��a<��a<k�a<�a<��a<J�a<֌a<j�a<Սa<W�a<��a<��a<*�a<i�a<ȏa<�a<z�a<��a<��a<!�a<Ғa<��a<J�a<�a<�a<��a<��a<	�a<��a<�a<�a<�a<%�a<�a<��a<�a<�a<n�a<��a<ԛa<6�a<]�a<ɜa<�a<s�a<��a<��a<�a<6�a<R�a<R�a<Q�a<�a<�a<��a<��a<w�a<P�a<D�a<T�a<e�a<��a<ٝa<%�a<|�a<֞a<*�a<��a<ڟa<��a<�a<'�a<<�a<4�a<�a<�a<ٟa<��a<��a<��a<L�a<r�a<w�a<U�a<p�a<��a<��a<|�a<q�a<E�a<!�a<�a<��a<O�a<̝a<h�a<��a<��a<(�a<ța<��a<^�a<0�a<&�a<5�a<6�a<[�a<o�a<��a<��a<��a<��a<h�a<4�a<�a<��a<l�a<
�a<��a<+�a<��a<��a<#�a<�a<��a<d�a<,�a<��a<��a<]�a<�a<~�a<�a<u�a<�a< �a<_�a<��a<Ȑa<�a<R�a<��a<
�a<��a<�a<��a<j�a<�a<ڋa<��a<T�a</�a<��a<]�a<׉a<T�a<ֈa<*�a<��a<��a<T�a<��a<E�a<��a<%�a<̃a<>�a<��a<��a<U�a<�a<��a<%�a<��a<H�a<�a<>a<}~a<�}a<D}a<�|a<$|a<�{a<.{a<�za<�za<{za<vza<{za<�za<�za<�za<�za<{a<{a<{a<�za<�za<�za<�za<�za<kza<<za<Dza<;za<za<Eza<gza<hza<�za<�za<{a<�  �  C{a<\{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a< |a<|a<�|a<�|a<\}a<�}a<P~a<
a<�a<_�a<��a<��a<�a<a<,�a<��a<�a<H�a<��a<�a<{�a<ۅa<^�a<��a<x�a< �a<Ĉa<��a<6�a<܊a<��a<4�a<��a<T�a<эa<;�a<��a<	�a<K�a<��a<�a<m�a<��a<?�a<Αa<X�a<,�a<��a<��a<F�a<�a<��a<a�a<�a<��a<6�a<n�a<�a<�a<E�a<��a<��a<ޚa<�a<W�a<��a<֛a<8�a<��a<�a<2�a<��a<�a<�a<S�a<3�a<N�a<4�a<7�a<�a<�a<��a<��a<��a<{�a<��a<��a<�a< �a<@�a<��a<�a<Z�a<��a<̟a<�a<�a<D�a<�a<-�a<�a<ݟa<��a<|�a<[�a<7�a<9�a<�a<#�a<.�a<A�a<Z�a<L�a<s�a<P�a<]�a<'�a<ڞa<��a<A�a<�a<��a<3�a<��a<g�a<�a<��a<��a<h�a<��a<c�a<b�a<��a<��a<��a<��a<��a<v�a<�a<8�a<�a<��a<)�a<ܙa<m�a<�a<��a<F�a<�a<��a<o�a<,�a<�a<Ėa<v�a<[�a<ەa<��a<��a<p�a<ғa<(�a<��a<��a<�a<-�a<��a<�a<S�a<Ѝa<G�a<�a<��a<M�a<�a<ŋa<j�a<�a<��a<>�a<��a<C�a<ψa<�a<j�a<͆a<�a<��a<�a<h�a<�a<m�a<�a<��a<z�a<�a<ׁa<��a<!�a<Ԁa<(�a<�a<!a<�~a<~a<q}a<�|a<J|a<�{a<d{a</{a<�za<�za<�za<�za<�za<�za<�za<�za<{a<	{a<{a<{a<�za<�za<�za<rza<>za<za<�ya<�ya<�ya<�ya<za<@za<{za<�za<�za<�  �  {a<J{a<{a<�{a<�{a<�{a<�{a<|a<�{a<�{a<|a<|a<7|a<j|a<�|a<}a<�}a<~a<�~a<-a<�a<��a<�a<��a</�a<��a<�a<z�a<ʃa<)�a<{�a<τa<?�a<��a<�a<��a<*�a<߇a<��a<3�a<�a<��a<z�a<�a<Ɍa<V�a<�a<M�a<Ǝa<1�a<o�a<�a<2�a<��a<�a<��a<�a<��a<S�a< �a<˔a<j�a<=�a<�a<q�a<7�a<��a<�a<Q�a<��a<ݙa<�a<0�a<r�a<��a<��a<�a<S�a<��a<��a<L�a<��a<�a<`�a<��a<�a<(�a<P�a<v�a<E�a<`�a<8�a<�a<�a<�a<םa<ҝa<֝a<�a<�a<]�a<��a<��a<�a<��a<��a<ڟa<�a<�a<�a<�a<�a<��a<��a<[�a<J�a<�a<��a<�a<۞a<ݞa<��a<�a< �a<$�a<3�a<=�a<2�a<�a<�a<��a<\�a<*�a<��a<X�a<��a<��a<Q�a<�a<ڛa<��a<��a<��a<��a<��a<��a<כa<��a<a<��a<]�a<�a<Қa<h�a<	�a<��a<'�a<̘a<Q�a<�a<��a<\�a<.�a<��a<��a<��a<N�a<�a<ƕa<q�a<��a<��a<�a<R�a<��a<ߑa<B�a<~�a<ӏa<*�a<��a<	�a<��a<2�a<ьa<��a<$�a<��a<��a< �a<�a<K�a<Ɖa<&�a<��a<�a<C�a<y�a<�a<D�a<��a<!�a<��a<'�a<݂a<~�a<1�a<��a<��a<b�a<��a<��a<E�a<�a<2a<�~a<0~a<�}a<"}a<�|a< |a<�{a<e{a<){a<{a<�za<�za<�za<�za<!{a<{a<{a<3{a<{a<�za<�za<�za<^za<?za<�ya<�ya<�ya<�ya<�ya<�ya<�ya<za<-za<�za<�za<�  �  �za<={a<l{a<�{a<�{a<�{a<|a<|a<*|a<4|a<A|a<Y|a<||a<�|a<�|a<n}a<�}a<Q~a<�~a<ra<�a<��a<3�a<��a<*�a<��a<��a<j�a<��a<��a<=�a<��a<�a<Q�a<Ѕa<G�a<�a<��a<L�a< �a<щa<��a<`�a<�a<��a<Y�a<�a<l�a<��a<R�a<��a<�a<��a<Ԑa<V�a<֑a<]�a<��a<��a<R�a<��a<��a<^�a<�a<��a<#�a<��a<��a<G�a<��a<��a<�a<�a<.�a<=�a<��a<��a<�a<P�a<��a<�a<q�a<��a<@�a<��a<�a<)�a<N�a<g�a<{�a<�a<g�a<X�a<5�a</�a<�a<(�a< �a<K�a<h�a<��a<ܞa<�a<`�a<��a<ޟa<�a<�a<�a<�a<��a<ϟa<��a<g�a<"�a<��a<��a<��a<��a<��a<��a<��a<��a<ߞa<��a<�a<0�a<�a<�a<��a<a<��a<?�a<�a<��a<9�a<�a<��a<l�a<"�a<�a<�a<�a<�a<�a<�a<�a<�a<��a<��a<^�a<�a<��a<H�a<ܙa<[�a<�a<s�a<�a<��a<V�a<"�a<Жa<��a<}�a<_�a<-�a<�a<��a<`�a<��a<��a<�a<��a<Вa<&�a<q�a<ΐa<�a<}�a<�a<^�a<�a<l�a<#�a<��a<j�a<�a<Ëa<F�a<Պa<L�a<��a<�a<��a<��a<�a<K�a<��a<��a<[�a<Ńa<T�a<�a<��a<F�a<��a<a<��a<U�a<�a<��a<C�a<�a<ha<�~a<_~a<�}a<L}a<�|a<Y|a<|a<�{a<�{a<P{a<7{a<2{a<,{a<8{a<9{a<L{a<.{a<({a<{a<�za<�za<{za<9za<�ya<�ya<�ya<Yya<_ya<Bya<nya<zya<�ya<�ya<Fza<�za<�  �  �za<�za<g{a<�{a<�{a<|a<-|a<>|a<T|a<t|a<{|a<�|a<�|a<	}a<b}a<�}a<~a<�~a<a<�a<(�a<��a<?�a<��a<&�a<��a<�a<.�a<��a<��a<�a<N�a<��a<�a<t�a<��a<��a<J�a<��a<Ոa<��a<h�a<?�a<ދa<ˌa<[�a<�a<s�a<�a<s�a<�a<H�a<��a<3�a<��a<*�a<��a<:�a<�a<��a<)�a<�a<��a<$�a<��a<(�a<��a<�a<�a<n�a<��a<��a<ԙa<ܙa<�a<,�a<a�a<��a<��a<d�a<Ǜa<@�a<��a<"�a<u�a<Ɲa<9�a<I�a<y�a<��a<��a<��a<��a<j�a<x�a<k�a<b�a<��a<��a<��a<�a<�a<W�a<��a<��a<�a<��a<�a<�a<
�a<��a<��a<d�a<&�a<�a<��a<��a<Z�a<@�a<=�a<H�a<f�a<��a<��a<��a<��a<�a<�a< �a<��a<מa<��a<`�a<�a<ԝa<s�a<>�a<�a<��a<��a<V�a<A�a<=�a<�a<5�a<�a<�a<�a<̛a<��a<h�a<�a<��a<.�a<��a<&�a<��a<7�a<��a<\�a<
�a<̖a<��a<e�a<R�a<�a<�a<�a<��a<s�a< �a<��a<
�a<��a<�a<\�a<��a<�a<m�a<��a<>�a<��a<*�a<ύa<b�a<�a<��a<3�a<Ӌa<N�a<يa<L�a<҉a<�a<X�a<��a<Æa<�a<O�a<��a<�a<r�a<��a<��a<E�a<��a<ǁa<z�a<c�a<�a<׀a<��a<>�a<�a<wa<
a<�~a<~a<�}a<%}a<�|a<K|a<|a<�{a<�{a<�{a<j{a<k{a<c{a<Y{a<]{a<?{a<'{a<{a<�za<}za<bza<za<�ya<�ya<Lya<ya<ya<�xa<ya<8ya<yya<�ya<za<Zza<�  �  �za<�za<O{a<�{a<�{a</|a<@|a<||a<{|a<�|a<�|a<�|a<}a<J}a<�}a<�}a<_~a<�~a<\a<�a<P�a<��a<L�a<�a<1�a<��a<ӂa<�a<h�a<��a<ރa<��a<p�a<ńa<-�a<Ņa<D�a<"�a<��a<��a<d�a<=�a<�a<ϋa<��a<B�a<"�a<��a<4�a<��a<�a<��a<��a<o�a<ݑa<m�a<��a<��a<*�a<ǔa<{�a<�a<��a<Z�a<��a<\�a<��a<٘a<�a<B�a<l�a<y�a<��a<��a<��a<ۙa<*�a<f�a<��a<4�a<t�a<�a<q�a<��a<O�a<��a<�a<M�a<��a<��a<ٞa<��a<a<Þa<��a<��a<��a<ўa<֞a<�a<,�a<^�a<��a<��a<��a<�a<#�a<-�a<��a<�a<��a<��a<6�a<�a<��a<p�a<S�a<�a<�a<�a<�a<!�a<.�a<|�a<��a<Ԟa<؞a<�a<��a<�a<��a<��a<��a<>�a<�a<��a<r�a<+�a<�a<՜a<��a<��a<q�a<n�a<d�a<;�a<N�a<��a<��a<��a<=�a<��a<e�a<�a<h�a<��a<N�a<��a<��a<�a<Ԗa<u�a<q�a<!�a<�a<�a<וa<��a<v�a<G�a<�a<��a</�a<��a<"�a<{�a<�a<D�a<��a<�a<��a<��a<r�a<	�a<��a<@�a<Ɍa<`�a<	�a<n�a<�a<;�a<��a<�a<-�a<q�a<��a<؅a<	�a<��a<��a<;�a<��a<N�a<�a<��a<��a<S�a<=�a<��a<ŀa<��a<B�a<�a<�a<Ia<�~a<F~a<�}a<U}a<�|a<�|a<`|a<|a<�{a<�{a<�{a<�{a<�{a<�{a<u{a<c{a<E{a<�za<�za<gza<<za<�ya<�ya<2ya<ya<�xa<�xa<�xa<�xa<ya<4ya<hya<�ya<-za<�  �  oza<�za<W{a<�{a<�{a<|a<`|a<�|a<�|a<�|a<�|a<}a<i}a<�}a<�}a<M~a<�~a<a<�a<�a<~�a<�a<r�a<́a<7�a<��a<�a<�a<;�a<n�a<��a<܃a<%�a<z�a<�a<w�a<�a<Ća<��a<Q�a<8�a<�a<�a<�a<��a<b�a<�a<��a<C�a<��a<L�a<��a<3�a<��a<>�a<��a<,�a<�a<V�a<�a<��a<J�a<ǖa<d�a<Ηa<:�a<��a<ޘa<.�a<'�a<@�a<O�a<R�a<v�a<��a<��a<ݙa<�a<u�a<�a<[�a<̛a<S�a<ќa<L�a<͝a<�a<]�a<��a<��a<ܞa<۞a<�a<�a<ޞa<�a<�a<�a<!�a<P�a<P�a<��a<şa<�a<�a<"�a<�a<�a<�a<�a<��a<]�a<�a<Оa<w�a<=�a<��a<͝a<ĝa<��a<��a<�a<�a<F�a<w�a<��a<�a<	�a<�a<�a<�a<ܞa<��a<y�a<<�a<�a<��a<��a<A�a<�a<��a<ќa<��a<��a<��a<i�a<S�a<%�a<ܛa<��a<E�a<�a<f�a<ڙa<O�a<��a<4�a<��a<6�a<іa<��a<A�a<�a<��a<Εa<ŕa<��a<��a<��a<J�a<�a<��a<6�a<Γa<9�a<��a<�a<�a<Аa<e�a<��a<.�a<׎a<5�a<Սa<j�a<�a<{�a<�a<|�a<�a<[�a<��a<�a<�a<E�a<s�a<��a<�a<&�a<�a<�a<o�a<�a<Áa<��a<S�a<5�a<�a<�a<ހa<��a<R�a<�a<�a<Ka<�~a<x~a<�}a<�}a<6}a<�|a<{|a<Z|a<9|a<�{a<�{a<�{a<�{a<�{a<�{a<\{a<3{a<{a<�za<za<	za<�ya<fya<
ya<�xa<�xa<vxa<�xa<�xa<�xa<�xa<Gya<�ya<za<�  �  Mza<�za<{a<�{a<�{a<B|a<�|a<�|a<�|a<�|a<"}a<R}a<x}a<�}a<�}a<d~a<�~a<La<�a<$�a<��a<��a<��a<�a<H�a<q�a<��a<��a<�a<R�a<p�a<��a<�a<c�a<Մa<;�a<�a<��a<d�a<0�a<�a<��a<Ŋa<��a<x�a<m�a<�a<ގa<V�a<ڏa<z�a<��a<l�a<ˑa<N�a<Ēa<P�a<��a<��a<H�a<��a<u�a<�a<l�a<�a<?�a<��a<��a<�a<��a<$�a<'�a<+�a<H�a<=�a<��a<��a<�a<f�a<��a<=�a<��a<3�a<��a<�a<��a<�a<l�a<��a<��a<מa<�a<�a<��a<.�a<�a<�a<�a<;�a<^�a<��a<��a<ǟa<�a<�a<F�a<K�a<#�a<�a<��a<��a<6�a<	�a<��a<X�a<	�a<ǝa<��a<��a<��a<��a<��a<�a<�a<h�a<|�a<��a<Ξa<�a<�a<�a<�a<��a<��a<D�a<�a<ޝa<��a<_�a<!�a<�a<�a<�a<��a<��a<��a<P�a<`�a<��a<��a<.�a<��a<8�a<��a<3�a<��a<�a<p�a<�a<��a<J�a<3�a<ѕa<̕a<��a<��a<��a<h�a<Y�a<�a<�a<��a<u�a<�a<X�a<�a<�a<��a<�a<u�a<؏a<Q�a<�a<e�a<�a<j�a</�a<��a<�a<��a<�a<e�a<��a<Èa<�a<)�a<L�a<t�a<��a<��a<q�a<��a<V�a<��a<{�a<n�a<*�a<�a<�a<a<��a<r�a<a�a<�a<�a<Ga<	a<�~a<~a<�}a<X}a<	}a<�|a<t|a<G|a<,|a<|a<�{a<�{a<�{a<�{a<�{a<;{a<{a<�za<Sza<�ya<�ya</ya<�xa<�xa<cxa<ixa<?xa<rxa<�xa<�xa<&ya<wya<za<�  �  Zza<�za<A{a<�{a<�{a</|a<c|a<�|a<�|a<}a<>}a<a}a<�}a<�}a<P~a<~~a<�~a<Ja<�a<<�a<ƀa<�a<y�a<݁a<2�a<��a<ɂa<�a<�a<)�a<d�a<��a<ރa<:�a<��a<�a<��a<��a<C�a<#�a<�a<�a<ߊa<ŋa<��a<S�a< �a<��a<D�a<��a<w�a<��a<o�a<��a<k�a<	�a<��a<�a<��a<@�a<�a<r�a<�a<i�a<ޗa<>�a<��a<ۘa<�a<�a<�a<�a<&�a<%�a<G�a<T�a<}�a<əa<0�a<��a<�a<��a<�a<��a<2�a<��a<�a<Q�a<��a<Þa<�a<'�a<�a<0�a<&�a<1�a<8�a<t�a<p�a<~�a<��a<֟a<��a< �a<1�a<%�a<2�a<�a<	�a<ܟa<��a<D�a<�a<��a<;�a<�a<��a<|�a<^�a<^�a<��a<��a<ŝa<��a<>�a<��a<Ξa<�a<�a<�a< �a<ޞa<Ӟa<��a<r�a<6�a<�a<��a<��a<z�a<(�a<	�a<�a<�a<��a<��a<g�a<,�a<�a<��a<@�a<֚a<L�a<��a<
�a<��a<�a<j�a<��a<��a<%�a<�a<ٕa<��a<��a<��a<��a<��a<l�a<@�a<��a<��a<K�a<Гa<u�a<�a<Z�a<��a<-�a<��a<�a<��a<��a<��a<�a<��a<-�a<��a<�a<��a<��a<C�a<��a<ڈa<�a<�a<3�a<o�a<��a<�a<,�a<��a<�a<Ɓa<~�a<=�a< �a<�a<�a<ـa<��a<��a<F�a<�a<�a<Ya<a<�~a<G~a<�}a<z}a<!}a<}a<�|a<f|a<G|a<,|a<|a<�{a<�{a<�{a<r{a</{a<�za<�za<bza<�ya<�ya<ya<�xa<�xa<]xa<%xa<xa<1xa<uxa<�xa< ya<eya<�ya<�  �  Iza<�za<({a<�{a<�{a<e|a<�|a<�|a<�|a<}a<E}a<i}a<�}a<�}a<#~a<x~a<a<Ca<�a<2�a<��a<=�a<��a<�a<;�a<|�a<��a<��a<�a<-�a<��a<�a<�a<�a<��a<Q�a<��a<��a<'�a<"�a<�a<�a<��a<��a<��a<N�a<9�a<Ԏa<q�a<�a<T�a<+�a<h�a<�a<x�a<�a<q�a<�a<Ӕa<7�a<�a<R�a<�a<��a<��a<��a<��a<Ҙa<Ҙa<�a<�a<�a<*�a<	�a<R�a<>�a<��a<ڙa<�a<��a<��a<��a<�a<��a<�a<��a<�a<V�a<ٞa<ܞa<�a<�a<�a<Z�a<�a<`�a<5�a<I�a<_�a<��a<��a<ҟa<�a<��a<N�a<K�a<`�a<8�a<�a<˟a<m�a<.�a<ݞa<��a<;�a<�a<��a<i�a<��a<S�a<w�a<��a<��a<�a<4�a<x�a<��a<ڞa< �a<�a<5�a<�a<��a<��a<�a<=�a<��a<�a<y�a<M�a<"�a<=�a<�a<�a<��a<��a<��a<D�a<+�a<��a<9�a<��a<�a<��a<�a<��a<חa<r�a<ږa<��a<`�a<֕a<ەa<��a<��a<��a<|�a<d�a<8�a<3�a<�a<ؔa<k�a<��a<��a<Ēa<��a<��a<H�a<��a<��a<r�a<�a<��a<�a<܍a<�a<Ìa<J�a<��a<3�a<E�a<��a<��a<ۇa<�a<<�a<s�a<|�a<��a<�a<a<+�a<��a<��a<%�a<4�a<�a<�a<��a<��a<��a<K�a<G�a<�a<�a<a<�~a<p~a<�}a<�}a<}a<�|a<�|a<�|a<N|a<(|a<,|a<�{a<�{a<�{a<�{a<P{a<�za<�za<,za<�ya<{ya<7ya<�xa<vxa<Vxa<xa<Txa<'xa<gxa<�xa<�xa<�ya<�ya<�  �  Zza<�za<A{a<�{a<�{a</|a<c|a<�|a<�|a<}a<>}a<a}a<�}a<�}a<P~a<~~a<�~a<Ja<�a<<�a<ƀa<�a<y�a<݁a<2�a<��a<ɂa<�a<�a<)�a<d�a<��a<ރa<:�a<��a<�a<��a<��a<C�a<#�a<�a<�a<ߊa<ŋa<��a<S�a< �a<��a<D�a<��a<w�a<��a<o�a<��a<k�a<	�a<��a<�a<��a<@�a<�a<r�a<�a<i�a<ޗa<>�a<��a<ۘa<�a<�a<�a<�a<&�a<%�a<G�a<T�a<}�a<əa<0�a<��a<�a<��a<�a<��a<2�a<��a<�a<Q�a<��a<Þa<�a<'�a<�a<0�a<&�a<1�a<8�a<t�a<p�a<~�a<��a<֟a<��a< �a<1�a<%�a<2�a<�a<	�a<ܟa<��a<D�a<�a<��a<;�a<�a<��a<|�a<^�a<^�a<��a<��a<ŝa<��a<>�a<��a<Ξa<�a<�a<�a< �a<ޞa<Ӟa<��a<r�a<6�a<�a<��a<��a<z�a<(�a<	�a<�a<�a<��a<��a<g�a<,�a<�a<��a<@�a<֚a<L�a<��a<
�a<��a<�a<j�a<��a<��a<%�a<�a<ٕa<��a<��a<��a<��a<��a<l�a<@�a<��a<��a<K�a<Гa<u�a<�a<Z�a<��a<-�a<��a<�a<��a<��a<��a<�a<��a<-�a<��a<�a<��a<��a<C�a<��a<ڈa<�a<�a<3�a<o�a<��a<�a<,�a<��a<�a<Ɓa<~�a<=�a< �a<�a<�a<ـa<��a<��a<F�a<�a<�a<Ya<a<�~a<G~a<�}a<z}a<!}a<}a<�|a<f|a<G|a<,|a<|a<�{a<�{a<�{a<r{a</{a<�za<�za<bza<�ya<�ya<ya<�xa<�xa<]xa<%xa<xa<1xa<uxa<�xa< ya<eya<�ya<�  �  Mza<�za<{a<�{a<�{a<B|a<�|a<�|a<�|a<�|a<"}a<R}a<x}a<�}a<�}a<d~a<�~a<La<�a<$�a<��a<��a<��a<�a<H�a<q�a<��a<��a<�a<R�a<p�a<��a<�a<c�a<Մa<;�a<�a<��a<d�a<0�a<�a<��a<Ŋa<��a<x�a<m�a<�a<ގa<V�a<ڏa<z�a<��a<l�a<ˑa<N�a<Ēa<P�a<��a<��a<H�a<��a<u�a<�a<l�a<�a<?�a<��a<��a<�a<��a<$�a<'�a<+�a<H�a<=�a<��a<��a<�a<f�a<��a<=�a<��a<3�a<��a<�a<��a<�a<l�a<��a<��a<מa<�a<�a<��a<.�a<�a<�a<�a<;�a<^�a<��a<��a<ǟa<�a<�a<F�a<K�a<#�a<�a<��a<��a<6�a<	�a<��a<X�a<	�a<ǝa<��a<��a<��a<��a<��a<�a<�a<h�a<|�a<��a<Ξa<�a<�a<�a<�a<��a<��a<D�a<�a<ޝa<��a<_�a<!�a<�a<�a<�a<��a<��a<��a<P�a<`�a<��a<��a<.�a<��a<8�a<��a<3�a<��a<�a<p�a<�a<��a<J�a<3�a<ѕa<̕a<��a<��a<��a<h�a<Y�a<�a<�a<��a<u�a<�a<X�a<�a<�a<��a<�a<u�a<؏a<Q�a<�a<e�a<�a<j�a</�a<��a<�a<��a<�a<e�a<��a<Èa<�a<)�a<L�a<t�a<��a<��a<q�a<��a<V�a<��a<{�a<n�a<*�a<�a<�a<a<��a<r�a<a�a<�a<�a<Ga<	a<�~a<~a<�}a<X}a<	}a<�|a<t|a<G|a<,|a<|a<�{a<�{a<�{a<�{a<�{a<;{a<{a<�za<Sza<�ya<�ya</ya<�xa<�xa<cxa<ixa<?xa<rxa<�xa<�xa<&ya<wya<za<�  �  oza<�za<W{a<�{a<�{a<|a<`|a<�|a<�|a<�|a<�|a<}a<i}a<�}a<�}a<M~a<�~a<a<�a<�a<~�a<�a<r�a<́a<7�a<��a<�a<�a<;�a<n�a<��a<܃a<%�a<z�a<�a<w�a<�a<Ća<��a<Q�a<8�a<�a<�a<�a<��a<b�a<�a<��a<C�a<��a<L�a<��a<3�a<��a<>�a<��a<,�a<�a<V�a<�a<��a<J�a<ǖa<d�a<Ηa<:�a<��a<ޘa<.�a<'�a<@�a<O�a<R�a<v�a<��a<��a<ݙa<�a<u�a<�a<[�a<̛a<S�a<ќa<L�a<͝a<�a<]�a<��a<��a<ܞa<۞a<�a<�a<ޞa<�a<�a<�a<!�a<P�a<P�a<��a<şa<�a<�a<"�a<�a<�a<�a<�a<��a<]�a<�a<Оa<w�a<=�a<��a<͝a<ĝa<��a<��a<�a<�a<F�a<w�a<��a<�a<	�a<�a<�a<�a<ܞa<��a<y�a<<�a<�a<��a<��a<A�a<�a<��a<ќa<��a<��a<��a<i�a<S�a<%�a<ܛa<��a<E�a<�a<f�a<ڙa<O�a<��a<4�a<��a<6�a<іa<��a<A�a<�a<��a<Εa<ŕa<��a<��a<��a<J�a<�a<��a<6�a<Γa<9�a<��a<�a<�a<Аa<e�a<��a<.�a<׎a<5�a<Սa<j�a<�a<{�a<�a<|�a<�a<[�a<��a<�a<�a<E�a<s�a<��a<�a<&�a<�a<�a<o�a<�a<Áa<��a<S�a<5�a<�a<�a<ހa<��a<R�a<�a<�a<Ka<�~a<x~a<�}a<�}a<6}a<�|a<{|a<Z|a<9|a<�{a<�{a<�{a<�{a<�{a<�{a<\{a<3{a<{a<�za<za<	za<�ya<fya<
ya<�xa<�xa<vxa<�xa<�xa<�xa<�xa<Gya<�ya<za<�  �  �za<�za<O{a<�{a<�{a</|a<@|a<||a<{|a<�|a<�|a<�|a<}a<J}a<�}a<�}a<_~a<�~a<\a<�a<P�a<��a<L�a<�a<1�a<��a<ӂa<�a<h�a<��a<ރa<��a<p�a<ńa<-�a<Ņa<D�a<"�a<��a<��a<d�a<=�a<�a<ϋa<��a<B�a<"�a<��a<4�a<��a<�a<��a<��a<o�a<ݑa<m�a<��a<��a<*�a<ǔa<{�a<�a<��a<Z�a<��a<\�a<��a<٘a<�a<B�a<l�a<y�a<��a<��a<��a<ۙa<*�a<f�a<��a<4�a<t�a<�a<q�a<��a<O�a<��a<�a<M�a<��a<��a<ٞa<��a<a<Þa<��a<��a<��a<ўa<֞a<�a<,�a<^�a<��a<��a<��a<�a<#�a<-�a<��a<�a<��a<��a<6�a<�a<��a<p�a<S�a<�a<�a<�a<�a<!�a<.�a<|�a<��a<Ԟa<؞a<�a<��a<�a<��a<��a<��a<>�a<�a<��a<r�a<+�a<�a<՜a<��a<��a<q�a<n�a<d�a<;�a<N�a<��a<��a<��a<=�a<��a<e�a<�a<h�a<��a<N�a<��a<��a<�a<Ԗa<u�a<q�a<!�a<�a<�a<וa<��a<v�a<G�a<�a<��a</�a<��a<"�a<{�a<�a<D�a<��a<�a<��a<��a<r�a<	�a<��a<@�a<Ɍa<`�a<	�a<n�a<�a<;�a<��a<�a<-�a<q�a<��a<؅a<	�a<��a<��a<;�a<��a<N�a<�a<��a<��a<S�a<=�a<��a<ŀa<��a<B�a<�a<�a<Ia<�~a<F~a<�}a<U}a<�|a<�|a<`|a<|a<�{a<�{a<�{a<�{a<�{a<�{a<u{a<c{a<E{a<�za<�za<gza<<za<�ya<�ya<2ya<ya<�xa<�xa<�xa<�xa<ya<4ya<hya<�ya<-za<�  �  �za<�za<g{a<�{a<�{a<|a<-|a<>|a<T|a<t|a<{|a<�|a<�|a<	}a<b}a<�}a<~a<�~a<a<�a<(�a<��a<?�a<��a<&�a<��a<�a<.�a<��a<��a<�a<N�a<��a<�a<t�a<��a<��a<J�a<��a<Ոa<��a<h�a<?�a<ދa<ˌa<[�a<�a<s�a<�a<s�a<�a<H�a<��a<3�a<��a<*�a<��a<:�a<�a<��a<)�a<�a<��a<$�a<��a<(�a<��a<�a<�a<n�a<��a<��a<ԙa<ܙa<�a<,�a<a�a<��a<��a<d�a<Ǜa<@�a<��a<"�a<u�a<Ɲa<9�a<I�a<y�a<��a<��a<��a<��a<j�a<x�a<k�a<b�a<��a<��a<��a<�a<�a<W�a<��a<��a<�a<��a<�a<�a<
�a<��a<��a<d�a<&�a<�a<��a<��a<Z�a<@�a<=�a<H�a<f�a<��a<��a<��a<��a<�a<�a< �a<��a<מa<��a<`�a<�a<ԝa<s�a<>�a<�a<��a<��a<V�a<A�a<=�a<�a<5�a<�a<�a<�a<̛a<��a<h�a<�a<��a<.�a<��a<&�a<��a<7�a<��a<\�a<
�a<̖a<��a<e�a<R�a<�a<�a<�a<��a<s�a< �a<��a<
�a<��a<�a<\�a<��a<�a<m�a<��a<>�a<��a<*�a<ύa<b�a<�a<��a<3�a<Ӌa<N�a<يa<L�a<҉a<�a<X�a<��a<Æa<�a<O�a<��a<�a<r�a<��a<��a<E�a<��a<ǁa<z�a<c�a<�a<׀a<��a<>�a<�a<wa<
a<�~a<~a<�}a<%}a<�|a<K|a<|a<�{a<�{a<�{a<j{a<k{a<c{a<Y{a<]{a<?{a<'{a<{a<�za<}za<bza<za<�ya<�ya<Lya<ya<ya<�xa<ya<8ya<yya<�ya<za<Zza<�  �  �za<={a<l{a<�{a<�{a<�{a<|a<|a<*|a<4|a<A|a<Y|a<||a<�|a<�|a<n}a<�}a<Q~a<�~a<ra<�a<��a<3�a<��a<*�a<��a<��a<j�a<��a<��a<=�a<��a<�a<Q�a<Ѕa<G�a<�a<��a<L�a< �a<щa<��a<`�a<�a<��a<Y�a<�a<l�a<��a<R�a<��a<�a<��a<Ԑa<V�a<֑a<]�a<��a<��a<R�a<��a<��a<^�a<�a<��a<#�a<��a<��a<G�a<��a<��a<�a<�a<.�a<=�a<��a<��a<�a<P�a<��a<�a<q�a<��a<@�a<��a<�a<)�a<N�a<g�a<{�a<�a<g�a<X�a<5�a</�a<�a<(�a< �a<K�a<h�a<��a<ܞa<�a<`�a<��a<ޟa<�a<�a<�a<�a<��a<ϟa<��a<g�a<"�a<��a<��a<��a<��a<��a<��a<��a<��a<ߞa<��a<�a<0�a<�a<�a<��a<a<��a<?�a<�a<��a<9�a<�a<��a<l�a<"�a<�a<�a<�a<�a<�a<�a<�a<�a<��a<��a<^�a<�a<��a<H�a<ܙa<[�a<�a<s�a<�a<��a<V�a<"�a<Жa<��a<}�a<_�a<-�a<�a<��a<`�a<��a<��a<�a<��a<Вa<&�a<q�a<ΐa<�a<}�a<�a<^�a<�a<l�a<#�a<��a<j�a<�a<Ëa<F�a<Պa<L�a<��a<�a<��a<��a<�a<K�a<��a<��a<[�a<Ńa<T�a<�a<��a<F�a<��a<a<��a<U�a<�a<��a<C�a<�a<ha<�~a<_~a<�}a<L}a<�|a<Y|a<|a<�{a<�{a<P{a<7{a<2{a<,{a<8{a<9{a<L{a<.{a<({a<{a<�za<�za<{za<9za<�ya<�ya<�ya<Yya<_ya<Bya<nya<zya<�ya<�ya<Fza<�za<�  �  {a<J{a<{a<�{a<�{a<�{a<�{a<|a<�{a<�{a<|a<|a<7|a<j|a<�|a<}a<�}a<~a<�~a<-a<�a<��a<�a<��a</�a<��a<�a<z�a<ʃa<)�a<{�a<τa<?�a<��a<�a<��a<*�a<߇a<��a<3�a<�a<��a<z�a<�a<Ɍa<V�a<�a<M�a<Ǝa<1�a<o�a<�a<2�a<��a<�a<��a<�a<��a<S�a< �a<˔a<j�a<=�a<�a<q�a<7�a<��a<�a<Q�a<��a<ݙa<�a<0�a<r�a<��a<��a<�a<S�a<��a<��a<L�a<��a<�a<`�a<��a<�a<(�a<P�a<v�a<E�a<`�a<8�a<�a<�a<�a<םa<ҝa<֝a<�a<�a<]�a<��a<��a<�a<��a<��a<ڟa<�a<�a<�a<�a<�a<��a<��a<[�a<J�a<�a<��a<�a<۞a<ݞa<��a<�a< �a<$�a<3�a<=�a<2�a<�a<�a<��a<\�a<*�a<��a<X�a<��a<��a<Q�a<�a<ڛa<��a<��a<��a<��a<��a<��a<כa<��a<a<��a<]�a<�a<Қa<h�a<	�a<��a<'�a<̘a<Q�a<�a<��a<\�a<.�a<��a<��a<��a<N�a<�a<ƕa<q�a<��a<��a<�a<R�a<��a<ߑa<B�a<~�a<ӏa<*�a<��a<	�a<��a<2�a<ьa<��a<$�a<��a<��a< �a<�a<K�a<Ɖa<&�a<��a<�a<C�a<y�a<�a<D�a<��a<!�a<��a<'�a<݂a<~�a<1�a<��a<��a<b�a<��a<��a<E�a<�a<2a<�~a<0~a<�}a<"}a<�|a< |a<�{a<e{a<){a<{a<�za<�za<�za<�za<!{a<{a<{a<3{a<{a<�za<�za<�za<^za<?za<�ya<�ya<�ya<�ya<�ya<�ya<�ya<za<-za<�za<�za<�  �  C{a<\{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a< |a<|a<�|a<�|a<\}a<�}a<P~a<
a<�a<_�a<��a<��a<�a<a<,�a<��a<�a<H�a<��a<�a<{�a<ۅa<^�a<��a<x�a< �a<Ĉa<��a<6�a<܊a<��a<4�a<��a<T�a<эa<;�a<��a<	�a<K�a<��a<�a<m�a<��a<?�a<Αa<X�a<,�a<��a<��a<F�a<�a<��a<a�a<�a<��a<6�a<n�a<�a<�a<E�a<��a<��a<ޚa<�a<W�a<��a<֛a<8�a<��a<�a<2�a<��a<�a<�a<S�a<3�a<N�a<4�a<7�a<�a<�a<��a<��a<��a<{�a<��a<��a<�a< �a<@�a<��a<�a<Z�a<��a<̟a<�a<�a<D�a<�a<-�a<�a<ݟa<��a<|�a<[�a<7�a<9�a<�a<#�a<.�a<A�a<Z�a<L�a<s�a<P�a<]�a<'�a<ڞa<��a<A�a<�a<��a<3�a<��a<g�a<�a<��a<��a<h�a<��a<c�a<b�a<��a<��a<��a<��a<��a<v�a<�a<8�a<�a<��a<)�a<ܙa<m�a<�a<��a<F�a<�a<��a<o�a<,�a<�a<Ėa<v�a<[�a<ەa<��a<��a<p�a<ғa<(�a<��a<��a<�a<-�a<��a<�a<S�a<Ѝa<G�a<�a<��a<M�a<�a<ŋa<j�a<�a<��a<>�a<��a<C�a<ψa<�a<j�a<͆a<�a<��a<�a<h�a<�a<m�a<�a<��a<z�a<�a<ׁa<��a<!�a<Ԁa<(�a<�a<!a<�~a<~a<q}a<�|a<J|a<�{a<d{a</{a<�za<�za<�za<�za<�za<�za<�za<�za<{a<	{a<{a<{a<�za<�za<�za<rza<>za<za<�ya<�ya<�ya<�ya<za<@za<{za<�za<�za<�  �  L{a<}{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<5|a<�|a<�|a<�}a<$~a<�~a<�a</�a<��a<��a<)�a<��a<(�a<��a<�a<��a<�a<L�a<��a<9�a<��a<�a<ׇa<Y�a<��a<��a<k�a<�a<��a<J�a<֌a<j�a<Սa<W�a<��a<��a<*�a<i�a<ȏa<�a<z�a<��a<��a<!�a<Ғa<��a<J�a<�a<�a<��a<��a<	�a<��a<�a<�a<�a<%�a<�a<��a<�a<�a<n�a<��a<ԛa<6�a<]�a<ɜa<�a<s�a<��a<��a<�a<6�a<R�a<R�a<Q�a<�a<�a<��a<��a<w�a<P�a<D�a<T�a<e�a<��a<ٝa<%�a<|�a<֞a<*�a<��a<ڟa<��a<�a<'�a<<�a<4�a<�a<�a<ٟa<��a<��a<��a<L�a<r�a<w�a<U�a<p�a<��a<��a<|�a<q�a<E�a<!�a<�a<��a<O�a<̝a<h�a<��a<��a<(�a<ța<��a<^�a<0�a<&�a<5�a<6�a<[�a<o�a<��a<��a<��a<��a<h�a<4�a<�a<��a<l�a<
�a<��a<+�a<��a<��a<#�a<�a<��a<d�a<,�a<��a<��a<]�a<�a<~�a<�a<u�a<�a< �a<_�a<��a<Ȑa<�a<R�a<��a<
�a<��a<�a<��a<j�a<�a<ڋa<��a<T�a</�a<��a<]�a<׉a<T�a<ֈa<*�a<��a<��a<T�a<��a<E�a<��a<%�a<̃a<>�a<��a<��a<U�a<�a<��a<%�a<��a<H�a<�a<>a<}~a<�}a<D}a<�|a<$|a<�{a<.{a<�za<�za<{za<vza<{za<�za<�za<�za<�za<{a<{a<{a<�za<�za<�za<�za<�za<kza<<za<Dza<;za<za<Eza<gza<hza<�za<�za<{a<�  �  S{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<e{a<p{a<d{a<�{a<�{a<�{a<z|a<�|a<e}a<~a<�~a<qa<�a<̀a<_�a<-�a<��a<[�a<σa<%�a<��a<�a<}�a<څa<G�a<��a<B�a<�a<�a<M�a<��a<��a<8�a<��a<��a<�a<w�a<��a<�a<f�a<��a<�a<B�a<��a<Ϗa<n�a<אa<X�a<�a<��a<m�a<#�a<��a<ȕa<|�a<?�a<�a<��a<�a<��a<�a<S�a<��a<��a<,�a<:�a<|�a<��a<�a<F�a<��a<��a<�a<��a<ĝa<�a<N�a<8�a<\�a<"�a<�a<�a<ԝa<��a<f�a<F�a<�a<7�a<�a<Q�a<w�a<��a<�a<I�a<��a<�a<[�a<��a<�a<1�a<C�a<u�a<4�a<K�a<�a<��a<�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<g�a<3�a<ߞa<q�a<%�a<��a<V�a<Ŝa<h�a<�a<��a<o�a<�a<$�a<�a<�a<�a<&�a<\�a<V�a<~�a<n�a<��a<m�a<h�a<'�a<Ěa<��a<
�a<ԙa<g�a<�a<��a<Q�a<�a<Ηa<��a<:�a<�a<Җa<Z�a<3�a<��a<�a<X�a<��a<�a<:�a<w�a<��a<�a<	�a<��a<�a<Z�a<�a<j�a<>�a<�a<��a<{�a<+�a<�a<��a<g�a<߉a<��a<وa<X�a<̇a<��a<��a<܅a<S�a<��a<@�a<܃a<v�a</�a<��a<��a<�a<��a<`�a<��a<R�a<�a<a<T~a<�}a<}a<||a<�{a<\{a<!{a<�za<�za<_za<7za<^za<^za<�za<�za<�za<�za< {a<&{a<{a<4{a<�za<�za<�za<�za<�za<[za<Uza<Aza<bza<xza<�za<�za<�za<L{a<�  �  r{a<�{a<�{a<�{a<�{a<�{a<�{a<�{a<i{a<U{a<G{a<U{a<s{a<�{a<�{a<5|a<�|a<G}a<�}a<�~a<Ra<�a<܀a<��a<"�a<��a<?�a<��a<D�a<��a<$�a<��a<��a<e�a<��a<��a<�a<��a<B�a<��a<��a<O�a<Ƌa<Y�a<�a<Y�a<׍a<2�a<~�a<��a<�a<:�a<w�a<֏a<3�a<��a<%�a<Бa<��a<G�a<�a<ޔa<��a<��a<Y�a<�a<��a<�a<��a<�a<m�a<��a<�a<!�a<b�a<��a<��a<0�a<b�a<��a<�a<Y�a<��a<�a<��a<(�a<3�a<G�a<C�a<,�a<��a<��a<y�a<T�a<%�a<�a<�a<�a<�a<T�a<��a<ڝa<=�a<��a<�a<m�a<��a<��a<�a<9�a<B�a<M�a<^�a<6�a<%�a<��a<ݟa<ɟa<��a<��a<��a<��a<��a<��a<��a<��a<u�a<X�a< �a<�a<��a<3�a<��a<,�a<��a<?�a<��a<��a<2�a<��a<ߚa<�a<�a<��a<�a<<�a<e�a<��a<��a<��a<c�a<K�a<	�a<�a<��a<C�a<�a<��a<"�a<��a<��a<3�a<�a<��a<s�a<#�a<�a<i�a< �a<��a<��a<v�a<ɓa<
�a<7�a<S�a<��a<Ïa<�a<Z�a<��a<&�a<��a<t�a<�a<�a<��a<r�a<E�a<�a<��a<D�a<��a<d�a<܈a<r�a<ˇa<7�a<��a<�a<m�a<
�a<��a<��a<��a<7�a<��a<��a<$�a<��a<9�a<��a<<�a<�a<a<j~a<�}a<�|a<k|a<�{a<a{a<�za<za<Pza<=za<.za<0za<Qza<kza<�za<�za< {a<{a<{a<{a<{a<�za<�za<�za<�za<�za<yza<rza<�za<�za<�za<�za<�za<{a<X{a<�  �  za<%za<Nza<Aza<za<�ya<�ya<�ya<_ya<`ya<ya<ya<ya<+ya<�ya<�ya<qza<�za<�{a<�|a<Y}a<O~a<�~a<�a<��a<_�a<�a<|�a<�a<<�a<�a<�a<��a<
�a<u�a<�a<��a<`�a<ׇa<Έa<D�a<�a<a<2�a<�a<�a<o�a<��a<�a< �a<;�a<��a<��a<�a<�a<Վa<q�a<��a<��a<h�a<��a<X�a<H�a<2�a<��a<זa<��a<Y�a<��a<;�a<��a<��a<#�a<
�a<r�a<��a<Қa<�a<d�a<��a<�a<��a<��a<�a<1�a<;�a<_�a<+�a<�a<��a<��a<3�a<��a<��a<E�a<9�a<�a<T�a<1�a<Y�a<��a<�a<��a<��a<��a<�a<a�a<��a<�a<]�a<Z�a<r�a<I�a<3�a<�a<͞a<՞a<��a<��a<v�a<��a<��a<��a<��a<��a<��a<��a<q�a<�a<��a<8�a<��a<J�a<��a<+�a<~�a< �a<��a<7�a<S�a<ۘa<��a<��a<K�a<��a<��a<�a<�a<@�a<Y�a<x�a<[�a</�a<�a<u�a<`�a<��a<r�a<�a<��a<m�a<
�a<��a<��a<��a<�a<�a<��a<�a<��a<�a<6�a<`�a<��a<��a<��a<��a<��a<$�a<7�a<ߋa<b�a<��a<y�a<�a<&�a<�a<ʉa<��a<m�a<H�a<��a<Ոa<-�a<Շa<9�a<j�a<�a<!�a<��a<��a<��a<��a<��a<3�a<��a<��a< �a<��a<n�a<�a<ta<�~a<~a<A}a<�|a<�{a<{a<^za<�ya<ya<kxa<rxa<�wa<�wa<�wa<�wa<Xxa<axa<�xa<�xa<,ya<bya<�ya<�ya<�ya<�ya<qya<Rya<:ya<�xa<�xa<�xa<�xa<�xa<ya<$ya<jya<�ya<�ya<�  �  �ya<za<"za<7za<>za<+za<�ya<�ya<wya<Fya<%ya<ya<)ya<-ya<vya<�ya<~za<{a<�{a<�|a<u}a<Q~a<%a<�a<��a<H�a<؁a<Y�a<�a<N�a<��a< �a<��a<�a<��a<�a<��a<V�a<�a<��a<P�a<	�a<��a<.�a<��a<"�a<��a<،a<�a<*�a<6�a<l�a<��a<��a<H�a<��a<2�a<�a<��a<�a<k�a<K�a<V�a<D�a<%�a<��a<��a<�a<��a<�a<x�a<��a<��a<�a<h�a<��a<ݚa<�a<`�a<��a<��a<Y�a<��a<�a<�a</�a<>�a<E�a<0�a<�a<��a<M�a<�a<��a<[�a<@�a<�a<�a<�a<|�a<˛a<#�a<��a<�a<��a<�a<��a<ߞa<�a<$�a<I�a<L�a<O�a<#�a<�a<�a<מa<��a<��a<��a<��a<��a<��a<��a<��a<��a<x�a<E�a<�a<Νa<j�a<לa<L�a<��a<�a<��a<�a<��a<9�a<�a<�a<
�a<�a<B�a<p�a<��a<�a<7�a<p�a<{�a<a�a<?�a<�a<�a<��a<2�a<͘a<z�a<�a<��a<u�a<�a<�a<��a<n�a<�a<��a<r�a<
�a<w�a<�a<Z�a<��a<��a<��a<��a<׎a<��a<5�a<j�a<��a<#�a<Ċa<��a<.�a<�a<ىa<׉a<��a<��a<k�a<�a<��a<0�a<��a<*�a<��a<�a<5�a<��a<�a<��a<�a<��a<4�a<Ɂa<x�a<�a<ƀa<I�a<�a<Sa<�~a<2~a<g}a<�|a<�{a<�za<Lza<�ya<ya<�xa<$xa<�wa<�wa<�wa<xa<7xa<sxa<�xa<ya<]ya<�ya<�ya<�ya<�ya<�ya<vya<Bya<,ya<ya<�xa<�xa<�xa<�xa<ya<=ya<fya<�ya<�ya<�  �  �ya<:za<6za<Cza<'za<	za<�ya<�ya<�ya<]ya<bya<3ya<Fya<�ya<�ya</za<�za<B{a<�{a<�|a<�}a<R~a<'a<�a<��a<G�a<��a<t�a<ła<K�a<��a<�a<Z�a<Єa<W�a<Ӆa<}�a<�a<Ӈa<q�a<D�a<�a<��a<e�a<��a<:�a<s�a<ƌa<��a<E�a<p�a<��a<�a<�a<��a<�a<u�a<;�a<Đa<őa<��a<~�a<z�a<A�a<�a<֖a<��a<�a<ݘa<	�a<S�a<��a<��a<�a<�a<h�a<��a<�a<-�a<x�a<�a<�a<��a<ɜa<�a<T�a<8�a<A�a<�a<�a<��a<|�a<
�a<ӛa<��a<I�a<a�a<I�a<n�a<��a<ޛa<c�a<��a<I�a<��a<�a<x�a<Ǟa<!�a<4�a<u�a<0�a<;�a<�a<�a<��a<��a<��a<a�a<h�a<V�a<j�a<}�a<x�a<��a<w�a<��a<Y�a<�a<��a<H�a<ڜa<P�a<ޛa<(�a<Ěa<(�a<șa<��a<>�a<@�a<�a<E�a<u�a<��a<�a<�a<9�a<H�a<n�a<`�a<_�a<&�a<��a<��a<��a<��a<:�a<ޗa<��a<0�a<��a<��a<��a<2�a<�a<��a<f�a<A�a<{�a<�a<:�a<�a<��a<ېa<�a<��a<6�a<<�a<��a<�a<f�a<�a<��a<u�a<2�a<�a<��a<��a<��a<H�a<�a<��a<e�a<��a<�a<{�a<��a<%�a<`�a<߃a<F�a<ւa<_�a<�a<��a<=�a<�a<��a<U�a<�a<Na<�~a<
~a<g}a<�|a<|a<!{a<{za<�ya<#ya<�xa<gxa<6xa<xa<xa<Fxa<Rxa<�xa<�xa<ya<Cya<jya<�ya<�ya<�ya<fya<bya<$ya< ya<�xa<�xa<�xa<�xa<�xa<�xa<ya<Cya<lya<�ya<�  �  �ya<�ya<za<?za<5za</za<za<�ya<�ya<�ya<�ya<wya<~ya<�ya<�ya<Hza<�za<v{a<'|a<�|a<�}a<~~a<Ua<�a<��a<H�a<��a<H�a<��a<�a<o�a<փa< �a<��a<�a<��a<M�a<ӆa<��a<W�a<�a<Ɖa<w�a<�a<��a<6�a<�a<��a<%�a<]�a<��a<Ía<�a<F�a<��a<�a<��a<G�a<	�a<�a<ƒa<��a<��a<k�a<N�a<�a<��a<�a<~�a<�a<4�a<t�a<��a<ؙa<�a<?�a<_�a<��a<�a<A�a<��a<�a<b�a<��a<�a<�a<9�a<I�a<"�a<�a<̜a<��a<<�a<��a<ƛa<��a<q�a<��a<��a<̛a<"�a<��a<�a<Y�a<Нa<@�a<��a<Ҟa<�a<�a<&�a<�a<�a<�a<��a<��a<U�a<P�a<.�a<3�a<&�a<-�a<T�a<^�a<n�a<`�a<\�a</�a<�a<ŝa<n�a<�a<{�a<�a<[�a<�a<l�a<�a<��a<��a<X�a<`�a<y�a<��a<ęa<��a</�a<g�a<h�a<w�a<a�a<�a<��a<��a<K�a<�a<��a< �a<��a<W�a<��a<ʖa<k�a<N�a<�a<ߕa<��a<R�a<�a<p�a<�a<F�a<��a<ϑa<��a<�a</�a<_�a<��a<��a<&�a<��a<!�a<͊a<��a<d�a<5�a<�a<�a<��a<T�a<�a<��a<�a<��a<�a<B�a<��a<�a<,�a<��a<�a<��a<9�a<��a<��a<'�a<ۀa<��a<.�a<�a<Na<�~a<$~a<�}a<�|a<|a<S{a<�za<za<hya<�xa<�xa<_xa<Cxa<Lxa<jxa<�xa<�xa<�xa<9ya<kya<uya<�ya<{ya<oya<Pya<4ya<ya<�xa<�xa<{xa<�xa<txa<�xa<�xa<�xa<ya<Rya<�ya<�  �  �ya<�ya<za<3za<@za<Eza<za<za<�ya<�ya<�ya<�ya<�ya<�ya<Xza<�za<D{a<�{a<d|a<;}a<�}a<�~a<Oa<�a<��a<I�a<��a<+�a<��a<Ԃa<&�a<v�a<�a<D�a<��a<E�a<ׅa<��a<R�a<�a<͈a<��a<^�a<�a<��a<�a<��a<��a<8�a<��a<ɍa<�a<0�a<��a<��a<x�a<�a<��a<��a<�a<�a<�a<��a<��a<P�a< �a<��a<&�a<r�a<՘a<�a<3�a<]�a<��a<��a<̙a<�a<D�a<��a<�a<U�a<��a<$�a<��a<֜a<�a<B�a<7�a<B�a<�a<�a<��a<��a<@�a<��a<�a<��a<�a<�a<6�a<��a<��a<F�a<��a<��a<D�a<��a<�a<
�a<!�a<�a<�a<̞a<��a<h�a<L�a<�a<ڝa<۝a<��a<؝a<��a<��a<�a<*�a<Q�a<?�a<3�a<�a<Нa<��a<�a<��a<�a<��a<�a<��a<l�a<��a<�a<��a<Йa<��a<ڙa<�a<#�a<S�a<a�a<��a<n�a<c�a<�a<ݙa<��a<�a<��a<#�a<ȗa<R�a<�a<��a<T�a<-�a<�a<Εa<��a<i�a<:�a<͔a<��a<�a<b�a<��a<�a<�a<K�a<��a<��a<��a< �a<��a<��a<|�a<K�a<Ċa<��a<s�a<7�a<��a<Éa<q�a<�a<��a<��a<p�a<��a< �a<M�a<��a<�a<C�a<��a<2�a<Ёa<��a< �a<߀a<��a<_�a<�a<�a<Wa<�~a<D~a<�}a<�|a<9|a<�{a<�za<2za<�ya<8ya<ya<�xa<�xa<�xa<�xa<�xa<�xa<$ya<=ya<zya<�ya<�ya<�ya<Uya<Bya<�xa<�xa<�xa<jxa<9xa<xa<!xa<xa<Sxa<�xa<�xa<ya<Qya<�  �  cya<�ya<�ya<za<Iza<Xza<Nza<Pza<0za<$za<za<za<'za<_za<�za<{a<z{a<|a<�|a<f}a<~a<�~a<za<4�a<��a<$�a<��a<��a<?�a<��a<�a<+�a<��a<�a<h�a<�a<��a<<�a<��a<��a<��a<]�a<�a<�a<��a<�a<��a<�a<z�a<ɍa<�a<a�a<��a<�a<Y�a<ޏa<n�a<�a<��a<z�a<b�a<�a<��a<��a<f�a<$�a<��a<��a<r�a<��a<Șa<�a<�a<&�a<P�a<|�a<��a<��a<H�a<��a<
�a<w�a<
�a<>�a<��a< �a<�a<8�a<c�a<9�a<)�a<�a<��a<��a<Y�a<:�a<1�a<H�a<Y�a<|�a<a<�a<~�a<Нa<9�a<��a<��a<��a<��a<�a< �a<��a<��a<p�a<�a<�a<��a<��a<w�a<t�a<v�a<��a<��a<��a<�a<�a<)�a<�a<��a<ٝa<��a<7�a<ߜa<_�a<�a<{�a<	�a<��a<k�a<F�a<�a<�a<�a<;�a<J�a<i�a<��a<��a<��a<o�a<>�a<�a<��a<7�a<�a<\�a<ؗa<i�a<��a<��a<F�a<�a<ԕa<��a<o�a<{�a<4�a<��a<͔a<Z�a<�a<~�a<Œa<#�a<`�a<��a<̏a<�a<.�a<{�a<�a<`�a<�a<��a<*�a<��a<��a<y�a<7�a<ىa<��a<�a<y�a<��a</�a<y�a<�a<�a<=�a<��a<�a<\�a<�a<z�a<$�a<Ԁa<��a<��a<�a<�a<�a<-a<�~a<e~a<�}a<+}a<z|a<�{a<J{a<�za<za<�ya<fya<!ya<�xa<�xa<�xa<ya<4ya<eya<{ya<�ya<�ya<wya<dya<Jya<�xa<�xa<�xa<+xa< xa<�wa<�wa<�wa<�wa<�wa<0xa<mxa<�xa<*ya<�  �  2ya<�ya<�ya<&za<Sza<hza<�za<mza<~za<dza<zza<�za<�za<�za<�za<�{a<�{a<|a<}a<�}a<]~a<�~a<�a<0�a<a<,�a<��a<߁a<	�a<^�a<��a<�a< �a<��a<��a<h�a</�a<Ѕa<��a<f�a<B�a<�a<�a<Ǌa<p�a<-�a<��a<2�a<��a<�a<V�a<��a<	�a<R�a<Ϗa<<�a<a<��a<�a<�a<��a<p�a<&�a<�a<��a<�a<��a<�a<F�a<p�a<��a<��a<��a<ܘa<�a< �a<1�a<��a<�a<<�a<Śa<�a<��a<�a<��a<֜a<�a<S�a<U�a<f�a<E�a<.�a<�a<ޜa<ʜa<��a<��a<��a<Ȝa<�a<(�a<��a<��a<�a<T�a<��a<מa<��a<�a<�a<؞a<��a<\�a<�a<͝a<��a<K�a<4�a<�a<�a<�a<:�a<b�a<�a<��a<ԝa<�a<�a<�a<�a<��a<l�a<��a<��a<0�a<ܛa<u�a<�a<��a<��a<��a<s�a<��a<��a<��a<��a<��a<��a<��a<��a<E�a<�a<��a<�a<��a<��a<��a<�a<��a<7�a<ŕa<��a<h�a<S�a<'�a<�a<�a<ʔa<��a<I�a<��a<x�a<�a<L�a<��a<ؐa<��a<]�a<��a<�a<F�a<��a<Z�a<��a<��a<6�a<��a<��a<^�a<�a<��a<�a<k�a<·a<�a<@�a<{�a<��a<�a<*�a<��a<�a<v�a<�a<��a<��a<8�a<!�a<�a<�a<}a</a<�~a<W~a<�}a<G}a<�|a<|a<�{a<{a<~za<%za<�ya<�ya<fya<Rya<cya<Wya<�ya<�ya<�ya<�ya<�ya<�ya<Nya<"ya<�xa<�xa<+xa<�wa<�wa<qwa<hwa<9wa<twa<�wa<�wa<)xa<sxa<�xa<�  �  ya<jya<�ya<za<Hza<�za<�za<�za<�za<�za<�za<�za<�za<4{a<z{a<�{a<O|a<�|a<R}a<~a<�~a<*a<�a<D�a<��a<'�a<l�a<��a<�a<�a<P�a<|�a<��a<�a<��a<#�a<��a<i�a<2�a<,�a<��a<�a<Љa<��a<��a<�a<��a<_�a<��a<$�a<��a<�a<Q�a<��a<.�a<��a<9�a<ݑa<��a<6�a<�a<Քa<\�a<�a<��a<!�a<��a<��a<�a<L�a<[�a<[�a<|�a<k�a<��a<��a<�a<%�a<q�a<ܙa<T�a<�a<Z�a<�a<[�a<��a<�a<=�a<f�a<��a<s�a<o�a<q�a<%�a<�a<�a<�a<�a<0�a<R�a<��a<ŝa<�a<t�a<��a<Ϟa<��a<�a<�a<�a<��a<s�a<�a<Ýa<|�a<"�a<ޜa<��a<��a<��a<��a<͜a<�a<;�a<r�a<��a<ϝa<��a<��a<؝a<ŝa<��a<0�a<��a<��a< �a<ћa<}�a<A�a<�a<�a<ۚa<Қa<Ța<��a<�a<ܚa<�a<��a<v�a<A�a<ԙa<f�a<�a<J�a<Ɨa<)�a<��a<#�a<˕a<��a<2�a<�a<�a<�a<Ôa<��a<��a<x�a<Y�a<�a<z�a<�a<i�a<��a<<�a<Y�a<��a<��a<P�a<��a<+�a<��a<K�a<�a<��a<c�a<݊a<�a<2�a<��a<�a<{�a<��a<�a<�a<)�a<k�a<��a<ɂa<�a<��a<�a<��a<X�a<�a<�a<�a<�a<�a<Za<0a<�~a<h~a<~a<u}a<�|a<�|a<�{a<V{a<�za<za<+za<�ya<�ya<�ya<�ya<�ya<�ya<�ya<�ya<�ya<�ya<qya<Mya<�xa<�xa<>xa<�wa<�wa<Awa<wa<�va<�va<�va<#wa<kwa<�wa</xa<�xa<�  �  �xa<:ya<�ya<za<dza<�za<�za<�za<�za<�za<{a<<{a<X{a<�{a<�{a<&|a<�|a<8}a<�}a<8~a<�~a<ua<�a<e�a<��a<�a<Z�a<s�a<��a<΁a<�a<�a<��a<̂a<%�a<ăa<C�a<5�a<ͅa<̆a<Ǉa<��a<��a<u�a<\�a<�a<ތa<d�a<��a<m�a<Վa<;�a<��a<�a<��a<��a<��a<0�a<�a<��a<@�a<�a<��a<F�a<��a<J�a<��a<ؗa< �a<�a<�a<'�a<$�a<�a<O�a<;�a<��a<��a<�a<��a<�a<��a<�a<��a<�a<��a<�a<F�a<��a<��a<��a<��a<��a<��a<~�a<k�a<S�a<l�a<w�a<��a<�a<�a<S�a<��a<՞a<��a<�a<�a<�a<Ҟa<w�a<8�a<ѝa<��a<�a<Ɯa<��a<E�a<V�a<*�a<j�a<}�a<��a<�a</�a<z�a<��a<�a<�a<��a<֝a<��a<|�a<�a<Ĝa<r�a<1�a<ۛa<��a<p�a<8�a<9�a<;�a<$�a<�a<�a<'�a<�a<Ԛa<��a<-�a<Ùa<%�a<��a<�a<��a<Öa<f�a<ڕa<]�a<!�a<��a<͔a<{�a<��a<��a<w�a<l�a<P�a<5�a<�a<��a<�a<��a<�a<W�a<��a<�a<W�a<��a<�a<��a<	�a<��a<=�a<ދa<��a<!�a<��a<1�a<��a< �a<T�a<��a<��a<̅a<��a<�a<�a<��a<��a<5�a<��a<N�a<$�a<�a<�a<�a<za<Va<Ka<a<�~a<�~a<~a<�}a<+}a<�|a<+|a<�{a<C{a<�za<�za<?za<#za<za<�ya<�ya<�ya<za<�ya<�ya<�ya<oya<4ya<�xa<nxa<�wa<�wa<7wa<�va<�va<yva<�va<�va<�va<wa<jwa< xa<Uxa<�  �  �xa<?ya<�ya<za<mza<�za<�za<�za<.{a<F{a<i{a<t{a<�{a<�{a</|a<�|a<�|a<s}a<~a<�~a<a<�a<�a<[�a<Ҁa<��a<O�a<k�a<��a<��a<��a<�a<�a<a�a<тa<i�a<��a<��a<��a<��a<z�a<w�a<u�a<{�a<>�a<&�a<ьa<e�a<�a<��a<�a<��a<�a<W�a<�a<e�a<�a<��a<�a<�a<��a<3�a<ʕa<`�a<ǖa<6�a<��a<��a<��a<��a<�a<�a<ߗa<ߗa<җa<�a<&�a<d�a<��a<3�a<řa<K�a<�a<z�a<	�a<��a<�a<_�a<~�a<��a<Нa<ڝa<֝a<ѝa<Ýa<��a<ʝa<��a<�a<�a<#�a<p�a<��a<ўa<�a<�a<�a<�a<��a<��a<}�a<�a<��a<:�a<ߜa<��a<9�a<��a<�a<ߛa<��a<.�a<p�a<��a<��a<S�a<��a<ɝa<�a<��a<ԝa<ǝa<��a<]�a<�a<̜a<i�a<2�a<��a<��a<��a<x�a<v�a<z�a<g�a<\�a<7�a<	�a<ʚa<��a<�a<��a<�a<}�a<җa<,�a<��a<��a<p�a<	�a<Ɣa<r�a<T�a<R�a<K�a<H�a<M�a<P�a<V�a<�a<��a<��a<�a<��a<)�a<��a<�a<U�a<��a<�a<o�a<ߍa<y�a<�a<��a<$�a<��a<L�a<يa<:�a<��a<�a<7�a<��a<��a<��a<��a<΃a<��a<�a<\�a<րa<Q�a<�a<�a<�a<ja<Za<Ra<Fa<Ca<�~a<�~a<�~a<(~a<�}a<d}a<�|a<x|a<|a<�{a<B{a<�za<�za<�za<Mza<Sza<@za<5za<za<za<�ya<�ya<tya<ya<�xa<Gxa<�wa<Zwa<�va<�va<_va<.va<7va<=va<zva<�va<6wa<�wa<$xa<�  �  �xa<ya<�ya< za<pza<�za<{a<{a<^{a<^{a<�{a<�{a<�{a<)|a<c|a<�|a< }a<�}a<%~a<�~a<9a<�a<J�a<o�a<؀a<�a<$�a<E�a<e�a<��a<��a<Ɓa<ׁa<@�a<��a<&�a<�a<v�a<v�a<\�a<I�a<o�a<K�a<J�a<(�a<�a<Ҍa<��a<6�a<��a<N�a<��a<;�a<��a<�a<��a<$�a<Œa<U�a<�a<��a<n�a<�a<{�a<#�a<>�a<��a<��a<̗a<̗a<�a<��a<��a<��a<��a<ڗa<�a<1�a<��a<�a<��a<�a<ǚa<`�a<�a<o�a<ݜa<c�a<��a<�a<�a<��a<�a<�a<��a<۝a<��a<��a< �a<7�a<^�a<��a<��a<�a<�a<E�a<@�a<�a<�a<��a<N�a<�a<��a<�a<��a<N�a<��a<��a<��a<a<a<�a<L�a<w�a<��a<&�a<v�a<��a<ܝa< �a<�a<�a<��a<��a<)�a<��a<��a<_�a<5�a<��a<�a<��a<��a<��a<��a<��a<K�a<]�a<ޚa<��a<�a<��a<��a<]�a<��a<��a<s�a<��a<N�a<ܔa<��a<d�a<�a<$�a<�a<�a<E�a<&�a<&�a< �a<�a<��a<q�a<ߒa<H�a<Бa<�a<��a<ȏa<7�a<��a<�a<��a<�a<όa<:�a<��a<j�a<�a<��a<��a<�a<)�a<U�a<g�a<��a<��a<��a<˂a<Ёa<Q�a<��a<�a<�a<ja<ha<5a<@a<8a<a<a<�~a<�~a<�~a<�~a<�}a<�}a<}a<�|a<7|a<�{a<t{a<{a<�za<�za<�za<�za<Uza<jza<4za<>za<za<�ya<iya<�xa<�xa<xa<�wa<%wa<�va<mva<va<va<�ua< va<>va<�va<wa<kwa<xa<�  �  �xa<ya<�ya<za<fza<�za<�za<9{a<h{a<�{a<�{a<�{a<|a<J|a<�|a<�|a<r}a<�}a<V~a<�~a<Qa<�a<�a<c�a<ƀa<�a<<�a<E�a<W�a<J�a<d�a<��a<ȁa<�a<U�a<�a<��a<n�a<4�a<.�a<"�a<A�a<H�a<K�a<O�a<�a<ڌa<��a<1�a<؎a<R�a<׏a<E�a<ϐa<F�a<בa<h�a<�a<��a<,�a<ޔa<t�a<�a<��a<�a<F�a<��a<їa<ӗa<Ηa<��a<��a<��a<n�a<��a<��a<��a<�a<f�a<�a<X�a<��a<��a<I�a<�a<��a<��a<L�a<��a<ҝa<��a<�a<�a<'�a<�a<.�a<�a<?�a<G�a<l�a<��a<��a<�a<�a<.�a<&�a<%�a<�a<��a<��a<M�a<�a<l�a<�a<��a< �a<�a<��a<s�a<n�a<��a<Λa<�a<`�a<��a<$�a<s�a<ɝa<�a<��a<�a<ߝa<ȝa<��a<Y�a<�a<ߜa<��a<W�a<?�a< �a<��a<ۛa<̛a<��a<��a<d�a</�a<Қa<��a<'�a<��a<��a<O�a<��a<ږa<1�a<��a<!�a<��a<>�a<
�a<�a<�a<�a<�a<�a<#�a<'�a<'�a<�a<��a<H�a<ڒa<o�a<ԑa<B�a<��a<
�a<h�a<�a<Z�a<̍a<a�a<یa<|�a<�a<��a<��a<b�a<��a<�a<M�a<\�a<i�a<k�a<W�a<r�a<��a<ˁa<��a<U�a<�a<�a<aa<"a<a<a<!a<$a<)a<a<�~a<�~a<Q~a<�}a<�}a<-}a<�|a<W|a<|a<�{a<\{a<{a<�za<�za<�za<�za<oza<Zza< za<�ya<�ya<zya<ya<�xa<xa<�wa<	wa<�va<?va<
va<�ua<�ua<�ua<$va<mva<�va<Twa<�wa<�  �  �xa<�xa<uya<�ya<sza<�za<{a<^{a<Z{a<�{a<�{a<�{a<|a<:|a<�|a<�|a<q}a<�}a<f~a<�~a<Ra<�a<)�a<��a<ʀa<�a<�a< �a<N�a<=�a<��a<y�a<��a<�a<o�a<-�a<q�a<j�a<�a<D�a<5�a<(�a<@�a<'�a<)�a<�a< �a<��a<V�a<�a<6�a<�a<2�a<ѐa<H�a<ʑa<]�a<�a<��a<�a<�a<V�a<�a<��a<�a<z�a<��a<��a<��a<��a<��a<��a<��a<W�a<��a<Z�a<�a<�a<5�a<՘a<K�a<�a<��a<>�a<Ǜa<Q�a<؜a<L�a<ǝa<ٝa<�a<'�a<�a<C�a<��a<3�a<�a<:�a<:�a<q�a<��a<��a<�a<��a<S�a<F�a<F�a<'�a<֞a<��a<"�a<�a<P�a<��a<��a<�a<қa<|�a<��a<f�a<��a<��a<�a<y�a<��a<"�a<H�a<��a<Νa<�a<�a<��a<�a<��a<{�a<�a<ʜa<��a<F�a<A�a<�a<��a<��a<ݛa<��a<��a<��a<<�a<�a<��a<�a<t�a<Ҙa<G�a<v�a<��a<'�a<��a<��a<��a<��a<�a<�a<Γa<�a<�a<��a<�a<�a<�a<ٓa<Ǔa<M�a<��a<��a<��a<p�a<��a<�a<j�a<Ԏa<N�a<Ǎa<h�a<ǌa<��a<�a<��a<"�a<`�a<�a<��a<*�a<3�a<Z�a<Z�a<g�a<��a<n�a<Ła<рa<��a<�a<ga<Pa<a<>a<a<a<a<�~a<�~a<�~a<�~a<X~a< ~a<�}a<(}a<�|a<<|a<|a<�{a<W{a<{a<�za<�za<�za<�za<`za<za<@za<za<�ya<Vya<�xa<kxa<xa<xwa<wa<�va<-va<�ua<�ua<va<�ua<va<]va<�va<mwa<�wa<�  �  �xa<ya<�ya<za<fza<�za<�za<9{a<h{a<�{a<�{a<�{a<|a<J|a<�|a<�|a<r}a<�}a<V~a<�~a<Qa<�a<�a<c�a<ƀa<�a<<�a<E�a<W�a<J�a<d�a<��a<ȁa<�a<U�a<�a<��a<n�a<4�a<.�a<"�a<A�a<H�a<K�a<O�a<�a<ڌa<��a<1�a<؎a<R�a<׏a<E�a<ϐa<F�a<בa<h�a<�a<��a<,�a<ޔa<t�a<�a<��a<�a<F�a<��a<їa<ӗa<Ηa<��a<��a<��a<n�a<��a<��a<��a<�a<f�a<�a<X�a<��a<��a<I�a<�a<��a<��a<L�a<��a<ҝa<��a<�a<�a<'�a<�a<.�a<�a<?�a<G�a<l�a<��a<��a<�a<�a<.�a<&�a<%�a<�a<��a<��a<M�a<�a<l�a<�a<��a< �a<�a<��a<s�a<n�a<��a<Λa<�a<`�a<��a<$�a<s�a<ɝa<�a<��a<�a<ߝa<ȝa<��a<Y�a<�a<ߜa<��a<W�a<?�a< �a<��a<ۛa<̛a<��a<��a<d�a</�a<Қa<��a<'�a<��a<��a<O�a<��a<ږa<1�a<��a<!�a<��a<>�a<
�a<�a<�a<�a<�a<�a<#�a<'�a<'�a<�a<��a<H�a<ڒa<o�a<ԑa<B�a<��a<
�a<h�a<�a<Z�a<̍a<a�a<یa<|�a<�a<��a<��a<b�a<��a<�a<M�a<\�a<i�a<k�a<W�a<r�a<��a<ˁa<��a<U�a<�a<�a<aa<"a<a<a<!a<$a<)a<a<�~a<�~a<Q~a<�}a<�}a<-}a<�|a<W|a<|a<�{a<\{a<{a<�za<�za<�za<�za<oza<Zza< za<�ya<�ya<zya<ya<�xa<xa<�wa<	wa<�va<?va<
va<�ua<�ua<�ua<$va<mva<�va<Twa<�wa<�  �  �xa<ya<�ya< za<pza<�za<{a<{a<^{a<^{a<�{a<�{a<�{a<)|a<c|a<�|a< }a<�}a<%~a<�~a<9a<�a<J�a<o�a<؀a<�a<$�a<E�a<e�a<��a<��a<Ɓa<ׁa<@�a<��a<&�a<�a<v�a<v�a<\�a<I�a<o�a<K�a<J�a<(�a<�a<Ҍa<��a<6�a<��a<N�a<��a<;�a<��a<�a<��a<$�a<Œa<U�a<�a<��a<n�a<�a<{�a<#�a<>�a<��a<��a<̗a<̗a<�a<��a<��a<��a<��a<ڗa<�a<1�a<��a<�a<��a<�a<ǚa<`�a<�a<o�a<ݜa<c�a<��a<�a<�a<��a<�a<�a<��a<۝a<��a<��a< �a<7�a<^�a<��a<��a<�a<�a<E�a<@�a<�a<�a<��a<N�a<�a<��a<�a<��a<N�a<��a<��a<��a<a<a<�a<L�a<w�a<��a<&�a<v�a<��a<ܝa< �a<�a<�a<��a<��a<)�a<��a<��a<_�a<5�a<��a<�a<��a<��a<��a<��a<��a<K�a<]�a<ޚa<��a<�a<��a<��a<]�a<��a<��a<s�a<��a<N�a<ܔa<��a<d�a<�a<$�a<�a<�a<E�a<&�a<&�a< �a<�a<��a<q�a<ߒa<H�a<Бa<�a<��a<ȏa<7�a<��a<�a<��a<�a<όa<:�a<��a<j�a<�a<��a<��a<�a<)�a<U�a<g�a<��a<��a<��a<˂a<Ёa<Q�a<��a<�a<�a<ja<ha<5a<@a<8a<a<a<�~a<�~a<�~a<�~a<�}a<�}a<}a<�|a<7|a<�{a<t{a<{a<�za<�za<�za<�za<Uza<jza<4za<>za<za<�ya<iya<�xa<�xa<xa<�wa<%wa<�va<mva<va<va<�ua< va<>va<�va<wa<kwa<xa<�  �  �xa<?ya<�ya<za<mza<�za<�za<�za<.{a<F{a<i{a<t{a<�{a<�{a</|a<�|a<�|a<s}a<~a<�~a<a<�a<�a<[�a<Ҁa<��a<O�a<k�a<��a<��a<��a<�a<�a<a�a<тa<i�a<��a<��a<��a<��a<z�a<w�a<u�a<{�a<>�a<&�a<ьa<e�a<�a<��a<�a<��a<�a<W�a<�a<e�a<�a<��a<�a<�a<��a<3�a<ʕa<`�a<ǖa<6�a<��a<��a<��a<��a<�a<�a<ߗa<ߗa<җa<�a<&�a<d�a<��a<3�a<řa<K�a<�a<z�a<	�a<��a<�a<_�a<~�a<��a<Нa<ڝa<֝a<ѝa<Ýa<��a<ʝa<��a<�a<�a<#�a<p�a<��a<ўa<�a<�a<�a<�a<��a<��a<}�a<�a<��a<:�a<ߜa<��a<9�a<��a<�a<ߛa<��a<.�a<p�a<��a<��a<S�a<��a<ɝa<�a<��a<ԝa<ǝa<��a<]�a<�a<̜a<i�a<2�a<��a<��a<��a<x�a<v�a<z�a<g�a<\�a<7�a<	�a<ʚa<��a<�a<��a<�a<}�a<җa<,�a<��a<��a<p�a<	�a<Ɣa<r�a<T�a<R�a<K�a<H�a<M�a<P�a<V�a<�a<��a<��a<�a<��a<)�a<��a<�a<U�a<��a<�a<o�a<ߍa<y�a<�a<��a<$�a<��a<L�a<يa<:�a<��a<�a<7�a<��a<��a<��a<��a<΃a<��a<�a<\�a<րa<Q�a<�a<�a<�a<ja<Za<Ra<Fa<Ca<�~a<�~a<�~a<(~a<�}a<d}a<�|a<x|a<|a<�{a<B{a<�za<�za<�za<Mza<Sza<@za<5za<za<za<�ya<�ya<tya<ya<�xa<Gxa<�wa<Zwa<�va<�va<_va<.va<7va<=va<zva<�va<6wa<�wa<$xa<�  �  �xa<:ya<�ya<za<dza<�za<�za<�za<�za<�za<{a<<{a<X{a<�{a<�{a<&|a<�|a<8}a<�}a<8~a<�~a<ua<�a<e�a<��a<�a<Z�a<s�a<��a<΁a<�a<�a<��a<̂a<%�a<ăa<C�a<5�a<ͅa<̆a<Ǉa<��a<��a<u�a<\�a<�a<ތa<d�a<��a<m�a<Վa<;�a<��a<�a<��a<��a<��a<0�a<�a<��a<@�a<�a<��a<F�a<��a<J�a<��a<ؗa< �a<�a<�a<'�a<$�a<�a<O�a<;�a<��a<��a<�a<��a<�a<��a<�a<��a<�a<��a<�a<F�a<��a<��a<��a<��a<��a<��a<~�a<k�a<S�a<l�a<w�a<��a<�a<�a<S�a<��a<՞a<��a<�a<�a<�a<Ҟa<w�a<8�a<ѝa<��a<�a<Ɯa<��a<E�a<V�a<*�a<j�a<}�a<��a<�a</�a<z�a<��a<�a<�a<��a<֝a<��a<|�a<�a<Ĝa<r�a<1�a<ۛa<��a<p�a<8�a<9�a<;�a<$�a<�a<�a<'�a<�a<Ԛa<��a<-�a<Ùa<%�a<��a<�a<��a<Öa<f�a<ڕa<]�a<!�a<��a<͔a<{�a<��a<��a<w�a<l�a<P�a<5�a<�a<��a<�a<��a<�a<W�a<��a<�a<W�a<��a<�a<��a<	�a<��a<=�a<ދa<��a<!�a<��a<1�a<��a< �a<T�a<��a<��a<̅a<��a<�a<�a<��a<��a<5�a<��a<N�a<$�a<�a<�a<�a<za<Va<Ka<a<�~a<�~a<~a<�}a<+}a<�|a<+|a<�{a<C{a<�za<�za<?za<#za<za<�ya<�ya<�ya<za<�ya<�ya<�ya<oya<4ya<�xa<nxa<�wa<�wa<7wa<�va<�va<yva<�va<�va<�va<wa<jwa< xa<Uxa<�  �  ya<jya<�ya<za<Hza<�za<�za<�za<�za<�za<�za<�za<�za<4{a<z{a<�{a<O|a<�|a<R}a<~a<�~a<*a<�a<D�a<��a<'�a<l�a<��a<�a<�a<P�a<|�a<��a<�a<��a<#�a<��a<i�a<2�a<,�a<��a<�a<Љa<��a<��a<�a<��a<_�a<��a<$�a<��a<�a<Q�a<��a<.�a<��a<9�a<ݑa<��a<6�a<�a<Քa<\�a<�a<��a<!�a<��a<��a<�a<L�a<[�a<[�a<|�a<k�a<��a<��a<�a<%�a<q�a<ܙa<T�a<�a<Z�a<�a<[�a<��a<�a<=�a<f�a<��a<s�a<o�a<q�a<%�a<�a<�a<�a<�a<0�a<R�a<��a<ŝa<�a<t�a<��a<Ϟa<��a<�a<�a<�a<��a<s�a<�a<Ýa<|�a<"�a<ޜa<��a<��a<��a<��a<͜a<�a<;�a<r�a<��a<ϝa<��a<��a<؝a<ŝa<��a<0�a<��a<��a< �a<ћa<}�a<A�a<�a<�a<ۚa<Қa<Ța<��a<�a<ܚa<�a<��a<v�a<A�a<ԙa<f�a<�a<J�a<Ɨa<)�a<��a<#�a<˕a<��a<2�a<�a<�a<�a<Ôa<��a<��a<x�a<Y�a<�a<z�a<�a<i�a<��a<<�a<Y�a<��a<��a<P�a<��a<+�a<��a<K�a<�a<��a<c�a<݊a<�a<2�a<��a<�a<{�a<��a<�a<�a<)�a<k�a<��a<ɂa<�a<��a<�a<��a<X�a<�a<�a<�a<�a<�a<Za<0a<�~a<h~a<~a<u}a<�|a<�|a<�{a<V{a<�za<za<+za<�ya<�ya<�ya<�ya<�ya<�ya<�ya<�ya<�ya<�ya<qya<Mya<�xa<�xa<>xa<�wa<�wa<Awa<wa<�va<�va<�va<#wa<kwa<�wa</xa<�xa<�  �  2ya<�ya<�ya<&za<Sza<hza<�za<mza<~za<dza<zza<�za<�za<�za<�za<�{a<�{a<|a<}a<�}a<]~a<�~a<�a<0�a<a<,�a<��a<߁a<	�a<^�a<��a<�a< �a<��a<��a<h�a</�a<Ѕa<��a<f�a<B�a<�a<�a<Ǌa<p�a<-�a<��a<2�a<��a<�a<V�a<��a<	�a<R�a<Ϗa<<�a<a<��a<�a<�a<��a<p�a<&�a<�a<��a<�a<��a<�a<F�a<p�a<��a<��a<��a<ܘa<�a< �a<1�a<��a<�a<<�a<Śa<�a<��a<�a<��a<֜a<�a<S�a<U�a<f�a<E�a<.�a<�a<ޜa<ʜa<��a<��a<��a<Ȝa<�a<(�a<��a<��a<�a<T�a<��a<מa<��a<�a<�a<؞a<��a<\�a<�a<͝a<��a<K�a<4�a<�a<�a<�a<:�a<b�a<�a<��a<ԝa<�a<�a<�a<�a<��a<l�a<��a<��a<0�a<ܛa<u�a<�a<��a<��a<��a<s�a<��a<��a<��a<��a<��a<��a<��a<��a<E�a<�a<��a<�a<��a<��a<��a<�a<��a<7�a<ŕa<��a<h�a<S�a<'�a<�a<�a<ʔa<��a<I�a<��a<x�a<�a<L�a<��a<ؐa<��a<]�a<��a<�a<F�a<��a<Z�a<��a<��a<6�a<��a<��a<^�a<�a<��a<�a<k�a<·a<�a<@�a<{�a<��a<�a<*�a<��a<�a<v�a<�a<��a<��a<8�a<!�a<�a<�a<}a</a<�~a<W~a<�}a<G}a<�|a<|a<�{a<{a<~za<%za<�ya<�ya<fya<Rya<cya<Wya<�ya<�ya<�ya<�ya<�ya<�ya<Nya<"ya<�xa<�xa<+xa<�wa<�wa<qwa<hwa<9wa<twa<�wa<�wa<)xa<sxa<�xa<�  �  cya<�ya<�ya<za<Iza<Xza<Nza<Pza<0za<$za<za<za<'za<_za<�za<{a<z{a<|a<�|a<f}a<~a<�~a<za<4�a<��a<$�a<��a<��a<?�a<��a<�a<+�a<��a<�a<h�a<�a<��a<<�a<��a<��a<��a<]�a<�a<�a<��a<�a<��a<�a<z�a<ɍa<�a<a�a<��a<�a<Y�a<ޏa<n�a<�a<��a<z�a<b�a<�a<��a<��a<f�a<$�a<��a<��a<r�a<��a<Șa<�a<�a<&�a<P�a<|�a<��a<��a<H�a<��a<
�a<w�a<
�a<>�a<��a< �a<�a<8�a<c�a<9�a<)�a<�a<��a<��a<Y�a<:�a<1�a<H�a<Y�a<|�a<a<�a<~�a<Нa<9�a<��a<��a<��a<��a<�a< �a<��a<��a<p�a<�a<�a<��a<��a<w�a<t�a<v�a<��a<��a<��a<�a<�a<)�a<�a<��a<ٝa<��a<7�a<ߜa<_�a<�a<{�a<	�a<��a<k�a<F�a<�a<�a<�a<;�a<J�a<i�a<��a<��a<��a<o�a<>�a<�a<��a<7�a<�a<\�a<ؗa<i�a<��a<��a<F�a<�a<ԕa<��a<o�a<{�a<4�a<��a<͔a<Z�a<�a<~�a<Œa<#�a<`�a<��a<̏a<�a<.�a<{�a<�a<`�a<�a<��a<*�a<��a<��a<y�a<7�a<ىa<��a<�a<y�a<��a</�a<y�a<�a<�a<=�a<��a<�a<\�a<�a<z�a<$�a<Ԁa<��a<��a<�a<�a<�a<-a<�~a<e~a<�}a<+}a<z|a<�{a<J{a<�za<za<�ya<fya<!ya<�xa<�xa<�xa<ya<4ya<eya<{ya<�ya<�ya<wya<dya<Jya<�xa<�xa<�xa<+xa< xa<�wa<�wa<�wa<�wa<�wa<0xa<mxa<�xa<*ya<�  �  �ya<�ya<za<3za<@za<Eza<za<za<�ya<�ya<�ya<�ya<�ya<�ya<Xza<�za<D{a<�{a<d|a<;}a<�}a<�~a<Oa<�a<��a<I�a<��a<+�a<��a<Ԃa<&�a<v�a<�a<D�a<��a<E�a<ׅa<��a<R�a<�a<͈a<��a<^�a<�a<��a<�a<��a<��a<8�a<��a<ɍa<�a<0�a<��a<��a<x�a<�a<��a<��a<�a<�a<�a<��a<��a<P�a< �a<��a<&�a<r�a<՘a<�a<3�a<]�a<��a<��a<̙a<�a<D�a<��a<�a<U�a<��a<$�a<��a<֜a<�a<B�a<7�a<B�a<�a<�a<��a<��a<@�a<��a<�a<��a<�a<�a<6�a<��a<��a<F�a<��a<��a<D�a<��a<�a<
�a<!�a<�a<�a<̞a<��a<h�a<L�a<�a<ڝa<۝a<��a<؝a<��a<��a<�a<*�a<Q�a<?�a<3�a<�a<Нa<��a<�a<��a<�a<��a<�a<��a<l�a<��a<�a<��a<Йa<��a<ڙa<�a<#�a<S�a<a�a<��a<n�a<c�a<�a<ݙa<��a<�a<��a<#�a<ȗa<R�a<�a<��a<T�a<-�a<�a<Εa<��a<i�a<:�a<͔a<��a<�a<b�a<��a<�a<�a<K�a<��a<��a<��a< �a<��a<��a<|�a<K�a<Ċa<��a<s�a<7�a<��a<Éa<q�a<�a<��a<��a<p�a<��a< �a<M�a<��a<�a<C�a<��a<2�a<Ёa<��a< �a<߀a<��a<_�a<�a<�a<Wa<�~a<D~a<�}a<�|a<9|a<�{a<�za<2za<�ya<8ya<ya<�xa<�xa<�xa<�xa<�xa<�xa<$ya<=ya<zya<�ya<�ya<�ya<Uya<Bya<�xa<�xa<�xa<jxa<9xa<xa<!xa<xa<Sxa<�xa<�xa<ya<Qya<�  �  �ya<�ya<za<?za<5za</za<za<�ya<�ya<�ya<�ya<wya<~ya<�ya<�ya<Hza<�za<v{a<'|a<�|a<�}a<~~a<Ua<�a<��a<H�a<��a<H�a<��a<�a<o�a<փa< �a<��a<�a<��a<M�a<ӆa<��a<W�a<�a<Ɖa<w�a<�a<��a<6�a<�a<��a<%�a<]�a<��a<Ía<�a<F�a<��a<�a<��a<G�a<	�a<�a<ƒa<��a<��a<k�a<N�a<�a<��a<�a<~�a<�a<4�a<t�a<��a<ؙa<�a<?�a<_�a<��a<�a<A�a<��a<�a<b�a<��a<�a<�a<9�a<I�a<"�a<�a<̜a<��a<<�a<��a<ƛa<��a<q�a<��a<��a<̛a<"�a<��a<�a<Y�a<Нa<@�a<��a<Ҟa<�a<�a<&�a<�a<�a<�a<��a<��a<U�a<P�a<.�a<3�a<&�a<-�a<T�a<^�a<n�a<`�a<\�a</�a<�a<ŝa<n�a<�a<{�a<�a<[�a<�a<l�a<�a<��a<��a<X�a<`�a<y�a<��a<ęa<��a</�a<g�a<h�a<w�a<a�a<�a<��a<��a<K�a<�a<��a< �a<��a<W�a<��a<ʖa<k�a<N�a<�a<ߕa<��a<R�a<�a<p�a<�a<F�a<��a<ϑa<��a<�a</�a<_�a<��a<��a<&�a<��a<!�a<͊a<��a<d�a<5�a<�a<�a<��a<T�a<�a<��a<�a<��a<�a<B�a<��a<�a<,�a<��a<�a<��a<9�a<��a<��a<'�a<ۀa<��a<.�a<�a<Na<�~a<$~a<�}a<�|a<|a<S{a<�za<za<hya<�xa<�xa<_xa<Cxa<Lxa<jxa<�xa<�xa<�xa<9ya<kya<uya<�ya<{ya<oya<Pya<4ya<ya<�xa<�xa<{xa<�xa<txa<�xa<�xa<�xa<ya<Rya<�ya<�  �  �ya<:za<6za<Cza<'za<	za<�ya<�ya<�ya<]ya<bya<3ya<Fya<�ya<�ya</za<�za<B{a<�{a<�|a<�}a<R~a<'a<�a<��a<G�a<��a<t�a<ła<K�a<��a<�a<Z�a<Єa<W�a<Ӆa<}�a<�a<Ӈa<q�a<D�a<�a<��a<e�a<��a<:�a<s�a<ƌa<��a<E�a<p�a<��a<�a<�a<��a<�a<u�a<;�a<Đa<őa<��a<~�a<z�a<A�a<�a<֖a<��a<�a<ݘa<	�a<S�a<��a<��a<�a<�a<h�a<��a<�a<-�a<x�a<�a<�a<��a<ɜa<�a<T�a<8�a<A�a<�a<�a<��a<|�a<
�a<ӛa<��a<I�a<a�a<I�a<n�a<��a<ޛa<c�a<��a<I�a<��a<�a<x�a<Ǟa<!�a<4�a<u�a<0�a<;�a<�a<�a<��a<��a<��a<a�a<h�a<V�a<j�a<}�a<x�a<��a<w�a<��a<Y�a<�a<��a<H�a<ڜa<P�a<ޛa<(�a<Ěa<(�a<șa<��a<>�a<@�a<�a<E�a<u�a<��a<�a<�a<9�a<H�a<n�a<`�a<_�a<&�a<��a<��a<��a<��a<:�a<ޗa<��a<0�a<��a<��a<��a<2�a<�a<��a<f�a<A�a<{�a<�a<:�a<�a<��a<ېa<�a<��a<6�a<<�a<��a<�a<f�a<�a<��a<u�a<2�a<�a<��a<��a<��a<H�a<�a<��a<e�a<��a<�a<{�a<��a<%�a<`�a<߃a<F�a<ւa<_�a<�a<��a<=�a<�a<��a<U�a<�a<Na<�~a<
~a<g}a<�|a<|a<!{a<{za<�ya<#ya<�xa<gxa<6xa<xa<xa<Fxa<Rxa<�xa<�xa<ya<Cya<jya<�ya<�ya<�ya<fya<bya<$ya< ya<�xa<�xa<�xa<�xa<�xa<�xa<ya<Cya<lya<�ya<�  �  �ya<za<"za<7za<>za<+za<�ya<�ya<wya<Fya<%ya<ya<)ya<-ya<vya<�ya<~za<{a<�{a<�|a<u}a<Q~a<%a<�a<��a<H�a<؁a<Y�a<�a<N�a<��a< �a<��a<�a<��a<�a<��a<V�a<�a<��a<P�a<	�a<��a<.�a<��a<"�a<��a<،a<�a<*�a<6�a<l�a<��a<��a<H�a<��a<2�a<�a<��a<�a<k�a<K�a<V�a<D�a<%�a<��a<��a<�a<��a<�a<x�a<��a<��a<�a<h�a<��a<ݚa<�a<`�a<��a<��a<Y�a<��a<�a<�a</�a<>�a<E�a<0�a<�a<��a<M�a<�a<��a<[�a<@�a<�a<�a<�a<|�a<˛a<#�a<��a<�a<��a<�a<��a<ߞa<�a<$�a<I�a<L�a<O�a<#�a<�a<�a<מa<��a<��a<��a<��a<��a<��a<��a<��a<��a<x�a<E�a<�a<Νa<j�a<לa<L�a<��a<�a<��a<�a<��a<9�a<�a<�a<
�a<�a<B�a<p�a<��a<�a<7�a<p�a<{�a<a�a<?�a<�a<�a<��a<2�a<͘a<z�a<�a<��a<u�a<�a<�a<��a<n�a<�a<��a<r�a<
�a<w�a<�a<Z�a<��a<��a<��a<��a<׎a<��a<5�a<j�a<��a<#�a<Ċa<��a<.�a<�a<ىa<׉a<��a<��a<k�a<�a<��a<0�a<��a<*�a<��a<�a<5�a<��a<�a<��a<�a<��a<4�a<Ɂa<x�a<�a<ƀa<I�a<�a<Sa<�~a<2~a<g}a<�|a<�{a<�za<Lza<�ya<ya<�xa<$xa<�wa<�wa<�wa<xa<7xa<sxa<�xa<ya<]ya<�ya<�ya<�ya<�ya<�ya<vya<Bya<,ya<ya<�xa<�xa<�xa<�xa<ya<=ya<fya<�ya<�ya<�  �  �xa<�xa<�xa<�xa<�xa<fxa<xa<�wa<Iwa<wa<�va<�va<�va<�va<�va<-wa<�wa<�xa<vya<eza<X{a<�|a<f}a<O~a<a<�a<��a< �a<��a<��a<��a<��a<7�a<��a<�a<τa<4�a<��a<��a<n�a<(�a<ۈa<��a<�a<��a<�a<(�a<^�a<x�a<��a<p�a<��a<��a<ɋa<�a<s�a<�a<��a<��a<|�a<��a<��a<Ւa<�a<�a<ƕa<��a<U�a<ؗa<J�a<��a<ܘa<�a<%�a<n�a<�a<�a<�a<S�a<��a< �a<��a<��a<�a<=�a<Z�a<W�a<�a<�a<��a<G�a<��a<-�a<əa<M�a< �a<Θa<�a<�a<H�a<��a<#�a<њa<Y�a<1�a<��a<D�a<��a<�a<T�a<i�a<m�a<U�a<@�a<�a<ȝa<��a<��a<��a<l�a<|�a<}�a<��a<��a<��a<��a<��a<o�a<�a<��a<�a<s�a<ޚa<�a<G�a<��a<�a<v�a<��a<�a<��a<�a<��a<S�a<��a<�a<��a<ܘa< �a<7�a<h�a<e�a<1�a<��a<��a<R�a<×a<p�a<��a<��a<~�a<�a<ߕa<��a<w�a<;�a<�a<��a<+�a<��a<�a<�a<<�a<A�a<;�a<�a<�a<�a<�a<&�a<r�a<�a<v�a<I�a<�a<�a<�a<"�a</�a<�a<�a<��a<��a<�a<��a<�a<M�a<��a<ڃa<N�a<��a<1�a<��a<�a<Ѐa<^�a<2�a<�a<ua<a<�~a<�}a<)}a<y|a<�{a<�za<�ya<�xa<�wa<wa<�va<�ua<�ua<Cua<Iua<Wua<�ua<�ua<Eva<�va<5wa<�wa<�wa<xa<;xa<7xa<(xa<xa<�wa<�wa<kwa<cwa<<wa<{wa<Owa<}wa<�wa<�wa<7xa<]xa<�  �  �xa<�xa<�xa<�xa<�xa<nxa<xa<�wa<gwa<wa<�va<�va<�va<�va<�va<Swa<�wa<�xa<ya<sza<l{a<_|a<i}a<_~a<.a<�a<��a<�a<��a<�a<`�a<��a<,�a<��a<��a<��a<2�a<�a<��a<[�a<�a<؈a<}�a<�a<��a<��a<1�a<d�a<f�a<z�a<��a<��a<��a<ڋa< �a<z�a<�a<Ӎa<��a<��a<��a<��a<˒a<Փa<�a<ҕa<��a<F�a<ٗa<B�a<��a<ؘa<�a<1�a<e�a<��a<��a<�a<Q�a<��a<�a<b�a<��a<�a<5�a<R�a<V�a<4�a<��a<��a< �a<��a<@�a<șa<`�a<(�a<��a<�a<�a<[�a<��a<9�a<Қa<}�a<�a<��a<H�a<��a<�a<;�a<j�a<c�a<V�a<%�a<��a<ҝa<��a<y�a<]�a<]�a<��a<��a<��a<��a<��a<��a<��a<V�a<�a<��a<!�a<k�a<��a<�a<J�a<��a<��a<��a<�a<ݖa<Ζa<�a<�a<\�a<��a<�a<v�a<��a<0�a<V�a<l�a<X�a<.�a<��a<��a<1�a<×a<e�a<��a<��a<7�a< �a<ڕa<��a<d�a<-�a<�a<��a<.�a<��a<��a<"�a<C�a</�a<+�a<!�a< �a<��a<�a<>�a<y�a<�a<��a<T�a<�a<�a<�a<�a<�a<�a<��a<Շa<t�a<�a<��a<�a<I�a<��a<�a<F�a<��a<��a<s�a<�a<Àa<c�a<�a<�a<qa<a<�~a<�}a<M}a<�|a<�{a<�za<�ya<�xa<�wa<*wa<�va<�ua<�ua<Wua<\ua<lua<�ua<�ua<iva<�va<)wa<�wa<�wa<xa<"xa<8xa<xa<xa<�wa<�wa<uwa<gwa<1wa<(wa<@wa<�wa<�wa<�wa<xa<bxa<�  �  fxa<�xa<�xa<�xa<�xa<uxa<1xa<�wa<�wa<3wa<wa<�va<�va<�va<wa<�wa<xa<�xa<�ya<�za<�{a<r|a<�}a<Z~a<*a<�a<��a<�a<p�a<�a<*�a<��a<�a<Z�a<ڃa<O�a<	�a<��a<r�a<.�a<�a<��a<X�a<�a<p�a<�a<'�a<��a<��a<��a<ċa<��a<�a<��a<H�a<��a<O�a<�a<Ŏa<׏a<ːa<��a<��a<��a<�a<ƕa<��a<0�a<їa<�a<l�a<��a<Ҙa<�a<�a<Z�a<z�a<̙a<�a<h�a<�a<-�a<��a<֛a<�a<F�a<C�a<1�a<�a<a<8�a<�a<n�a<��a<��a<@�a<:�a<#�a<O�a<�a<ޙa<~�a<��a<��a< �a<˜a<W�a<��a<�a<&�a<b�a<8�a<7�a<��a<؝a<��a<g�a<U�a<#�a<8�a<1�a<B�a<l�a<k�a<��a<�a<��a<?�a<�a<��a<'�a<��a<Śa<C�a<n�a<ݘa<%�a<��a<b�a<�a<�a<�a<B�a<��a<�a<S�a<��a<�a<+�a<R�a<]�a<I�a< �a<Ƙa<��a<��a<��a<�a<��a<g�a<��a<֕a<��a<l�a<6�a< �a<Ɣa<p�a<'�a<}�a<�a<�a<^�a<T�a<J�a<Z�a<-�a<>�a<-�a<f�a<��a<0�a<Ȉa<k�a<c�a<>�a<T�a<A�a<4�a<>�a<�a<هa<^�a<�a<b�a<Ņa<�a<b�a<��a<�a<l�a<Áa<Q�a<�a<x�a<@�a<�a<�a<@a<�~a<}~a<�}a<J}a<�|a<�{a<�za<�ya<ya<2xa<fwa<�va<>va<�ua<�ua<�ua<�ua<�ua<"va<�va<�va<Kwa<�wa<�wa<xa<xa<0xa<�wa<�wa<�wa<ywa<>wa<wa<wa<�va<wa<2wa<gwa<�wa<�wa<Fxa<�  �  Ixa<�xa<�xa<�xa<�xa<xa<Jxa<xa<�wa<hwa<Cwa<wa<wa<,wa<lwa<�wa<sxa<!ya<�ya<�za<�{a<�|a<�}a<i~a<4a<�a<`�a<�a<L�a<��a<��a<L�a<��a<��a<�a<�a<��a<]�a<#�a<�a<��a<��a<<�a<݉a<v�a<�a<:�a<��a<��a<ҋa<ыa<�a<�a<T�a<��a<�a<��a<R�a<.�a<�a<
�a<	�a<#�a<"�a<�a<ڕa<��a<5�a<��a<�a<W�a<m�a<��a<��a<Ҙa<��a<9�a<{�a<��a<(�a<��a<��a<\�a<��a<�a<�a<E�a<:�a<�a<ța<x�a<�a<��a<?�a<�a<��a<x�a<q�a<��a<�a<9�a<��a<1�a<Ǜa<m�a<�a<`�a<��a<�a<"�a<-�a<�a<	�a<��a<��a<T�a<�a<��a<�a<֜a<ݜa<�a<$�a<6�a<a�a<b�a<^�a<5�a<�a<��a<1�a<��a<�a<[�a<��a<�a<z�a<	�a<��a<h�a<U�a<h�a<��a<՗a<�a<t�a<Әa<�a<:�a<\�a<^�a<(�a<��a<��a<@�a<ɗa<S�a<ޖa<b�a<�a<ƕa<w�a<C�a<�a<��a<Ɣa<��a<T�a<�a<��a<�a<,�a<e�a<z�a<��a<g�a<l�a<y�a<��a<a<�a<�a<�a<Ԉa<��a<~�a<g�a<o�a<`�a<C�a<�a<Їa<c�a<نa<J�a<��a<߄a<$�a<g�a<��a<	�a<��a< �a<��a<8�a<�a<�a<ga<$a<�~a<W~a<�}a<S}a<�|a<�{a<	{a<za<7ya<txa<�wa<wa<|va<va<�ua<�ua<�ua<$va<Zva<�va< wa<mwa<�wa<�wa<xa<
xa<�wa<�wa<�wa<cwa<3wa<�va<�va<�va<�va<�va<�va<&wa<qwa<�wa<xa<�  �  "xa<Zxa<�xa<�xa<�xa<�xa<kxa<Pxa<�wa<�wa<�wa<xwa<�wa<�wa<�wa<Axa<�xa<}ya<Wza<1{a<|a<�|a<�}a<�~a</a<�a<P�a<��a<!�a<O�a<��a<�a<J�a<��a<�a<��a<&�a<�a<��a<��a<V�a<C�a<�a<��a<x�a<�a<`�a<��a<�a<�a<%�a<i�a<l�a<Ōa<
�a<��a<�a<��a<��a<`�a<�a<a�a<j�a<V�a<-�a<�a<��a<1�a<��a<՗a<�a<�a<>�a<L�a<{�a<{�a<ǘa< �a<Q�a<љa<%�a<��a<��a<��a<՛a<�a<<�a<2�a<,�a<ߛa<��a<P�a<��a<��a<:�a<*�a<�a<��a<�a<L�a<��a<
�a<��a<�a<��a<�a<��a<ϝa<��a<"�a<	�a<��a<��a<k�a<)�a<�a<��a<u�a<x�a<[�a<��a<��a<��a<�a<�a<;�a<5�a<1�a<��a<��a<U�a<Ǜa<P�a<��a<�a<n�a<ܘa<|�a<�a<�a<��a<�a<�a<5�a<|�a<��a<�a<'�a<c�a<X�a<X�a<�a<јa<w�a<�a<y�a<�a<��a<��a<��a<R�a<�a<�a<��a<��a<i�a<[�a<$�a<ѓa<��a<�a<R�a<��a<��a<ɏa<��a<�a<Ȍa<�a<)�a<��a<��a<}�a<G�a<�a<�a<��a<��a<��a<`�a<0�a<a<`�a<��a<�a<e�a<�a<΃a<�a<\�a<��a<�a<��a<�a<�a<�a<\a<	a<�~a<�~a<?~a<�}a<K}a<�|a<�{a<B{a<hza<�ya<�xa<xa<�wa<�va<�va<Sva<Lva<Tva<vva<�va<�va<awa<�wa<�wa<�wa<xa<	xa<�wa<�wa<^wa<wa<�va<�va<kva<-va<Cva<>va<�va<�va<wa<_wa<�wa<�  �  �wa<,xa<uxa<�xa<�xa<�xa<�xa<�xa<Wxa<(xa<xa<�wa<�wa<%xa<rxa<�xa<Mya<�ya<�za<z{a<\|a<*}a<�}a<�~a<0a<�a<<�a<��a<̀a<�a<C�a<��a<��a<�a<��a<�a<Ńa<h�a<H�a<7�a<�a<��a<ňa<��a<L�a<�a<R�a<ʋa<#�a<O�a<��a<��a<��a<-�a<��a<�a<��a<:�a<�a<�a<Ցa<��a<��a<��a<Y�a<��a<��a<
�a<u�a<��a<��a<ӗa<��a<�a<ܗa<�a<F�a<��a<ۘa<1�a<˙a<B�a<Úa<3�a<��a<��a<#�a<3�a<.�a<"�a<�a<��a<A�a< �a<��a<��a<j�a<z�a<��a<��a<�a<��a<�a<o�a<ޜa<]�a<��a<Ɲa<��a<��a<�a<��a<l�a< �a<Ӝa<j�a<+�a<�a<�a<��a<��a<�a<\�a<��a<ǜa<�a<�a<�a<��a<��a<q�a<�a<��a<��a<c�a<�a<T�a<�a<��a<o�a<J�a<C�a<g�a<��a<Ęa<�a<A�a<p�a<o�a<Y�a<D�a<�a<��a<"�a<��a<�a<��a<�a<��a<�a<Δa<��a<N�a<A�a<?�a<(�a<�a<ݓa<��a<X�a<�a<D�a<��a<�a<��a<�a<3�a<Q�a<j�a<��a<�a<�a<��a<��a<z�a<I�a<�a<��a<шa<��a<$�a<Ƈa<9�a<��a<څa<�a<E�a<q�a<��a<��a<#�a<��a<�a<�a<Aa<)a<�~a<�~a<�~a<g~a<4~a<�}a<K}a<�|a<1|a<w{a<�za<�ya<4ya<�xa<�wa<nwa<"wa<�va<�va<�va<�va<wa<[wa<�wa<�wa<�wa<�wa<xa<�wa<�wa<]wa<wa<�va<tva<va<�ua<�ua<�ua<�ua<�ua<2va<�va<wa<vwa<�  �  {wa<�wa<Axa<�xa<�xa<�xa<�xa<�xa<�xa<xxa<�xa<|xa<�xa<�xa<�xa<oya<�ya<�za<-{a<�{a<�|a<Z}a<~a<�~a<ba<�a<�a<P�a<x�a<��a<��a<�a<>�a<��a<��a<p�a<E�a<�a<�a<��a<��a<��a<��a<r�a<�a<�a<f�a<�a<J�a<��a<�a<�a<��a<��a<(�a<��a<�a<ݏa<��a<|�a<&�a<#�a<��a<��a<~�a<�a<Ŗa<��a<9�a<P�a<q�a<m�a<R�a<~�a<]�a<��a<��a<�a<b�a<��a<`�a<��a<m�a<ޚa<[�a<��a<�a<e�a<7�a<K�a<�a<�a<��a<m�a<Q�a<�a<�a<��a<�a<U�a<��a<�a<?�a<ٜa<�a<��a<��a<�a<	�a<Ɲa<��a<W�a<%�a<��a<U�a<�a<��a<��a<?�a<l�a<v�a<��a<�a<�a<y�a<��a<՜a<ٜa<��a<֜a<}�a<9�a<��a<d�a<��a<]�a<ߙa<x�a</�a<Ҙa<�a<˘a<��a<
�a< �a<s�a<q�a<��a<u�a<��a<)�a<ǘa<b�a<Ηa<U�a<��a<#�a<w�a<�a<��a<�a<�a<˓a<�a<��a<��a<Ǔa<��a<��a<(�a<�a<X�a<ɑa<�a<J�a<��a<|�a<ݍa<�a<F�a<��a<�a<��a<(�a<�a<��a<��a<G�a<��a<��a<3�a<�a<�a<p�a<��a<ʄa<ރa<�a<4�a<>�a<��a<�a<qa<)a<�~a<�~a<a~a<x~a<H~a<)~a<�}a<�}a<}}a<�|a<Y|a<�{a<{a<Gza<�ya<ya<gxa<xa<�wa<jwa<Uwa<Mwa<ywa<hwa<�wa<�wa<xa<xa<xa<xa<�wa<}wa<wa<�va<>va<�ua<�ua<Wua<Iua<
ua<Oua<wua<�ua<5va<�va<(wa<�  �  Ewa<�wa<7xa<}xa<�xa<�xa<ya<ya<ya<ya<�xa<�xa<ya<Cya<�ya<�ya<Vza<�za<�{a<X|a<}a<�}a<T~a<�~a<Pa<�a<�a<*�a<5�a<U�a<k�a<��a<��a<�a<w�a<�a<��a<d�a<X�a<I�a<>�a<V�a<S�a<G�a<�a<يa<��a<)�a<��a<�a<I�a<��a<�a<#�a<��a<#�a<��a<X�a<��a<�a<��a<��a<J�a<��a<��a<,�a<��a<Җa<�a<%�a<�a<�a<��a<�a<ܖa<�a</�a<l�a<×a<;�a<Ԙa<h�a<�a<��a<6�a<��a<�a<I�a<i�a<��a<Z�a<E�a<�a<�a<��a<��a<��a<��a<��a<ӛa<�a<z�a<͜a<*�a<r�a<��a<�a<��a<ٝa<��a<��a<&�a<��a<B�a<ߛa<u�a< �a<�a<ޚa<֚a<�a<�a<p�a<��a<�a<^�a<��a<Мa<Μa<ڜa<��a<k�a<�a<��a<A�a<Ϛa<E�a<��a<��a<��a<j�a<M�a<Z�a<��a<��a<��a<��a<˙a<��a<y�a<�a<��a<<�a<��a<�a<<�a<��a<�a<h�a<�a<��a<m�a<J�a<R�a<Q�a<P�a<n�a<k�a<[�a<�a<ڒa<x�a<�a<R�a<��a<ߏa<�a<G�a<a�a<��a<"�a<��a<�a<��a<p�a<*�a<�a<��a<>�a<�a<Z�a<Ça<�a<H�a<j�a<u�a<v�a<��a<��a<��a<�a<wa<�~a<�~a<K~a<3~a<~a<~a< ~a<~a<�}a<�}a<b}a<�|a<�|a<�{a<\{a<�za<'za<zya<�xa<�xa<8xa<�wa<�wa<�wa<�wa<�wa<xa<&xa<7xa<>xa<#xa<�wa<�wa<Zwa<�va<kva<�ua<�ua<ua<�ta<�ta<�ta<�ta<�ta<?ua<�ua<1va<�va<�  �  wa<�wa<xa<�xa<�xa<!ya<Aya<cya<Pya<Zya<Zya<vya<�ya<�ya<za<Qza<�za<h{a<|a<�|a<M}a<�}a<u~a<a<Ma<�a<�a<�a<�a<�a<�a<�a<J�a<��a<�a<��a<�a<�a<̓a<�a<�a<�a<�a<
�a<�a<يa<��a<4�a<ƌa<@�a<��a<��a<G�a<Ďa<�a<��a<6�a<Ɛa<��a<G�a<�a<��a<��a<>�a<ƕa<O�a<��a<ݖa<ߖa<�a<֖a<��a<��a<a�a<��a<p�a<��a<�a<H�a<їa<N�a<�a<��a<c�a<�a<~�a<��a<C�a<��a<��a<��a<��a<`�a<I�a<$�a< �a<�a<�a<�a<W�a<��a<Ԝa<,�a<i�a<ȝa<�a<�a<�a<ٝa<��a<?�a<�a<c�a<��a<z�a<��a<a<b�a<`�a<D�a<�a<��a< �a<l�a<��a<+�a<d�a<��a<ќa<�a<Ӝa<��a<d�a<�a<��a<,�a<ښa<��a<%�a<	�a<͙a<�a<ՙa<�a<�a<�a<
�a<�a<ԙa<v�a<�a<��a<�a<Z�a<��a<�a<�a<��a<�a<w�a<4�a<�a<��a<ƒa<��a<�a<�a<6�a<�a<�a<ڒa<��a<�a<��a<�a<�a<t�a<��a<�a<2�a<��a<�a<��a<D�a<ӊa<��a<�a<�a<|�a<��a<}�a<��a<�a<�a<0�a</�a< �a<3�a<�a<a�a<�a<�~a<h~a<~a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<[}a<'}a<�|a<4|a<�{a<{a<}za<�ya<�ya<�xa<�xa<kxa<Wxa<Sxa<@xa<Uxa<Uxa<{xa<mxa<Wxa<4xa<�wa<�wa<wa<�va<va<�ua<ua<�ta<nta<ta<,ta<(ta<�ta<�ta<Mua<�ua<bva<�  �  �va<jwa<�wa<xa<�xa<&ya<jya<�ya<�ya<�ya<�ya<�ya<�ya<&za<�za<�za<G{a<�{a<j|a<�|a<�}a<~a<�~a<a<[a<�a<�a<�a<�a<�a<�a<�a<�a<%�a<��a<��a<��a<��a<v�a<��a<��a<��a<�a<�a<�a<�a<��a<N�a<�a<y�a<��a<L�a<��a<�a<��a<�a<��a<>�a<�a<��a<i�a<�a<ߔa<n�a<�a<T�a<��a<��a<Ėa<��a<��a<T�a<1�a<�a<	�a<�a<*�a<{�a<��a<b�a<�a<��a<Q�a<�a<Úa<^�a<ڛa<P�a<��a<��a<ќa<�a<��a<��a<��a<y�a<t�a<��a<��a<��a<��a<A�a<}�a<ŝa<�a<�a<�a<�a<ܝa<��a<%�a<��a<$�a<��a<�a<��a<E�a<��a<ٙa<ܙa<	�a<B�a<��a<��a<u�a<�a<D�a<��a<Мa<�a<؜a<Ɯa<��a<L�a<�a<��a<:�a<ݚa<��a<��a<Q�a<>�a<A�a<I�a<B�a<W�a<2�a<�a<әa<��a< �a<r�a<˗a<�a<>�a<w�a<˔a<�a<��a<�a<��a<|�a<u�a<o�a<��a<��a<Ғa<��a<�a<��a<�a<��a<,�a<��a<)�a<v�a<ŏa<�a<V�a<��a<�a<��a<�a<��a<6�a<݊a<}�a<,�a<��a<�a<��a<·a<�a<��a<��a<�a<Ƃa<a<ƀa<�a<a<s~a< ~a<�}a<r}a<_}a<T}a<]}a<�}a<�}a<�}a<~}a<h}a<%}a<�|a<a|a<�{a<`{a<�za<[za<�ya<xya<2ya<�xa<�xa<�xa<�xa<�xa<�xa<�xa<�xa<cxa<<xa<�wa<nwa<�va<rva<�ua</ua<�ta<Ata<�sa<�sa<�sa<�sa<ta<hta<�ta<sua<$va<�  �  �va<Uwa<�wa<sxa<�xa<5ya<�ya<�ya<�ya<�ya<za<za<Bza<�za<�za<3{a<�{a<|a<�|a<.}a<�}a<8~a<�~a< a<ma<wa<�a<�a<xa<�a<la<�a<�a<�a<5�a<��a<p�a<'�a<6�a<D�a<p�a<��a<��a<�a<׉a<݊a<��a<u�a<�a<��a< �a<��a<�a<[�a<�a<e�a<�a<��a<4�a<�a<��a<\�a<��a<��a<�a<Q�a<��a<��a<��a<��a<c�a<;�a<�a<֕a<��a<��a<ܕa<$�a<��a<�a<ŗa<c�a<C�a<ߙa<��a<X�a<ța<d�a<��a<�a<�a<�a<��a<�a<ޜa<��a<Ҝa<��a<�a<�a<;�a<��a<��a<�a<�a<?�a<,�a<�a<ѝa<x�a<�a<k�a<�a<\�a<ߚa<O�a<ݙa<��a<��a<��a<��a<�a<k�a<Ěa<Y�a<��a<0�a<��a<Üa<�a<�a<��a<��a<��a<�a<�a<z�a<3�a< �a<��a<��a<��a<��a<��a<y�a<�a<P�a<E�a<ҙa<��a<�a<k�a<��a<ϖa<-�a<=�a<��a<��a<)�a<��a<b�a<=�a<�a<0�a<L�a<��a<��a<��a< �a<�a<ޒa<��a<T�a<בa<A�a<��a<��a<`�a<��a<�a<c�a<Ќa<d�a<ڋa<��a<�a<��a<B�a<ŉa<E�a<~�a<Їa<Άa<��a<ʄa<��a<��a<��a<��a<�a<�~a<%~a<�}a<I}a<}a<#}a<}a<N}a<H}a<m}a<�}a<m}a<|}a< }a<�|a<�|a<|a<�{a< {a<�za<za<�ya<hya<Dya<ya<�xa<�xa<�xa<�xa<�xa<�xa<xa<<xa<�wa<`wa<�va<&va<�ua<ua<�ta<�sa<�sa<vsa<Psa<�sa<�sa<ta<�ta<@ua<va<�  �  zva<2wa<�wa<sxa<�xa<Lya<�ya<�ya<za<za<1za<Zza<�za<�za<�za<W{a<�{a<P|a<�|a<Z}a<�}a<a~a<�~a<a<ia<{a<�a<ta<ia<aa<Ea<Ba<aa<�a<�a<w�a</�a<�a<��a<�a<?�a<k�a<��a<Ɉa<��a<ߊa<��a<�a<)�a<Ía<I�a<��a<)�a<��a<�a<��a<�a<ʑa<��a<+�a<֓a<��a<%�a<��a<�a<h�a<��a<��a<��a<f�a<8�a<�a<a<��a<��a<��a<��a<ޕa<Z�a<�a<��a<8�a<�a<ƙa<|�a<>�a<ϛa<_�a<��a<��a<�a<*�a< �a<�a<�a<�a<��a<��a<�a<S�a<��a<��a<�a<�a<E�a<K�a<>�a<�a<֝a<|�a<��a<Z�a<Λa<7�a<��a<�a<ƙa<t�a<L�a<S�a<��a<a<*�a<��a<�a<��a<�a<��a<Ĝa<��a<��a<��a<ۜa<��a<N�a<�a<��a<�a<$�a<�a<Ԛa<ݚa<��a<��a<��a<��a<y�a<M�a<�a<��a<��a<X�a<��a<��a<��a<�a<J�a<��a<�a<y�a<&�a<��a<��a<�a<�a<Q�a<��a<��a<ݒa<�a<��a<��a<]�a<�a<t�a<ߐa<.�a<��a<�a<3�a<��a<��a<��a<,�a<��a<J�a<�a<r�a<�a<M�a<��a<χa<چa<ԅa<��a<��a<x�a<T�a<H�a<ia<�~a<�}a<c}a<"}a<�|a<�|a<�|a<}a</}a<I}a<u}a<t}a<x}a<5}a<}a<�|a<A|a<�{a<J{a<�za<xza<�ya<�ya<hya<Sya<7ya<ya<ya<
ya<�xa<�xa<�xa<Ixa<�wa<cwa<�va<va<{ua<�ta<Dta<�sa<rsa<-sa<sa<7sa<�sa<�sa<xta<ua<�ua<�  �  �va<8wa<�wa<\xa<�xa<cya<�ya<�ya<�ya<4za<6za<Yza<�za<�za<A{a<`{a<�{a<E|a<�|a<r}a<�}a<j~a<�~a<.a<Ua<oa<�a<�a<�a<<a<Fa<-a<Ma<�a<�a<w�a<	�a<�a<�a<�a<-�a<c�a<��a<ňa<Љa<��a<ċa<��a<4�a<ōa<B�a<Ўa<#�a<��a<�a<��a<T�a<Ǒa<��a< �a<�a<��a<$�a<��a<�a<r�a<~�a<��a<��a<��a<<�a<�a<˕a<}�a<��a<c�a<��a<ؕa<D�a<Ԗa<i�a<=�a<�a<ٙa<��a<9�a<ƛa<F�a<��a<�a<�a<-�a<2�a<*�a<��a<�a<��a<C�a</�a<Q�a<��a<��a<	�a<�a<I�a<K�a<M�a<�a<��a<n�a<��a<��a<��a<+�a<��a<�a<��a<O�a<R�a<2�a<x�a<��a<�a<��a<�a<��a<�a<y�a<��a<�a<�a<��a<�a<��a<p�a<�a<��a<|�a<6�a<>�a<ݚa<ܚa<��a<Ěa<��a<��a<��a<J�a<�a<~�a<�a<R�a<��a<ؖa<ҕa<�a<5�a<��a<�a<k�a<'�a<֑a<�a<ܑa<�a<?�a<z�a<͒a<ْa<ݒa<��a<��a<e�a<��a<u�a<ؐa<I�a<~�a<�a<3�a<��a<4�a<��a<6�a<��a<`�a<�a<q�a<��a<O�a<��a<��a<͆a<ͅa<˄a<��a<e�a<\�a<3�a<`a<u~a<�}a<]}a<}a<�|a<�|a<�|a<�|a<C}a<X}a<o}a<k}a<^}a<N}a< }a<�|a<D|a<�{a<]{a<�za<|za<za<�ya<�ya<Pya<?ya<ya<2ya<�xa<�xa<�xa<�xa<Cxa<�wa<Vwa<�va<>va<dua<�ta<6ta<�sa<fsa<sa<sa<sa<{sa<�sa<eta<ua<�ua<�  �  zva<2wa<�wa<sxa<�xa<Lya<�ya<�ya<za<za<1za<Zza<�za<�za<�za<W{a<�{a<P|a<�|a<Z}a<�}a<a~a<�~a<a<ia<{a<�a<ta<ia<aa<Ea<Ba<aa<�a<�a<w�a</�a<�a<��a<�a<?�a<k�a<��a<Ɉa<��a<ߊa<��a<�a<)�a<Ía<I�a<��a<)�a<��a<�a<��a<�a<ʑa<��a<+�a<֓a<��a<%�a<��a<�a<h�a<��a<��a<��a<f�a<8�a<�a<a<��a<��a<��a<��a<ޕa<Z�a<�a<��a<8�a<�a<ƙa<|�a<>�a<ϛa<_�a<��a<��a<�a<*�a< �a<�a<�a<�a<��a<��a<�a<S�a<��a<��a<�a<�a<E�a<K�a<>�a<�a<֝a<|�a<��a<Z�a<Λa<7�a<��a<�a<ƙa<t�a<L�a<S�a<��a<a<*�a<��a<�a<��a<�a<��a<Ĝa<��a<��a<��a<ۜa<��a<N�a<�a<��a<�a<$�a<�a<Ԛa<ݚa<��a<��a<��a<��a<y�a<M�a<�a<��a<��a<X�a<��a<��a<��a<�a<J�a<��a<�a<y�a<&�a<��a<��a<�a<�a<Q�a<��a<��a<ݒa<�a<��a<��a<]�a<�a<t�a<ߐa<.�a<��a<�a<3�a<��a<��a<��a<,�a<��a<J�a<�a<r�a<�a<M�a<��a<χa<چa<ԅa<��a<��a<x�a<T�a<H�a<ia<�~a<�}a<c}a<"}a<�|a<�|a<�|a<}a</}a<I}a<u}a<t}a<x}a<5}a<}a<�|a<A|a<�{a<J{a<�za<xza<�ya<�ya<hya<Sya<7ya<ya<ya<
ya<�xa<�xa<�xa<Ixa<�wa<cwa<�va<va<{ua<�ta<Dta<�sa<rsa<-sa<sa<7sa<�sa<�sa<xta<ua<�ua<�  �  �va<Uwa<�wa<sxa<�xa<5ya<�ya<�ya<�ya<�ya<za<za<Bza<�za<�za<3{a<�{a<|a<�|a<.}a<�}a<8~a<�~a< a<ma<wa<�a<�a<xa<�a<la<�a<�a<�a<5�a<��a<p�a<'�a<6�a<D�a<p�a<��a<��a<�a<׉a<݊a<��a<u�a<�a<��a< �a<��a<�a<[�a<�a<e�a<�a<��a<4�a<�a<��a<\�a<��a<��a<�a<Q�a<��a<��a<��a<��a<c�a<;�a<�a<֕a<��a<��a<ܕa<$�a<��a<�a<ŗa<c�a<C�a<ߙa<��a<X�a<ța<d�a<��a<�a<�a<�a<��a<�a<ޜa<��a<Ҝa<��a<�a<�a<;�a<��a<��a<�a<�a<?�a<,�a<�a<ѝa<x�a<�a<k�a<�a<\�a<ߚa<O�a<ݙa<��a<��a<��a<��a<�a<k�a<Ěa<Y�a<��a<0�a<��a<Üa<�a<�a<��a<��a<��a<�a<�a<z�a<3�a< �a<��a<��a<��a<��a<��a<y�a<�a<P�a<E�a<ҙa<��a<�a<k�a<��a<ϖa<-�a<=�a<��a<��a<)�a<��a<b�a<=�a<�a<0�a<L�a<��a<��a<��a< �a<�a<ޒa<��a<T�a<בa<A�a<��a<��a<`�a<��a<�a<c�a<Ќa<d�a<ڋa<��a<�a<��a<B�a<ŉa<E�a<~�a<Їa<Άa<��a<ʄa<��a<��a<��a<��a<�a<�~a<%~a<�}a<I}a<}a<#}a<}a<N}a<H}a<m}a<�}a<m}a<|}a< }a<�|a<�|a<|a<�{a< {a<�za<za<�ya<hya<Dya<ya<�xa<�xa<�xa<�xa<�xa<�xa<xa<<xa<�wa<`wa<�va<&va<�ua<ua<�ta<�sa<�sa<vsa<Psa<�sa<�sa<ta<�ta<@ua<va<�  �  �va<jwa<�wa<xa<�xa<&ya<jya<�ya<�ya<�ya<�ya<�ya<�ya<&za<�za<�za<G{a<�{a<j|a<�|a<�}a<~a<�~a<a<[a<�a<�a<�a<�a<�a<�a<�a<�a<%�a<��a<��a<��a<��a<v�a<��a<��a<��a<�a<�a<�a<�a<��a<N�a<�a<y�a<��a<L�a<��a<�a<��a<�a<��a<>�a<�a<��a<i�a<�a<ߔa<n�a<�a<T�a<��a<��a<Ėa<��a<��a<T�a<1�a<�a<	�a<�a<*�a<{�a<��a<b�a<�a<��a<Q�a<�a<Úa<^�a<ڛa<P�a<��a<��a<ќa<�a<��a<��a<��a<y�a<t�a<��a<��a<��a<��a<A�a<}�a<ŝa<�a<�a<�a<�a<ܝa<��a<%�a<��a<$�a<��a<�a<��a<E�a<��a<ٙa<ܙa<	�a<B�a<��a<��a<u�a<�a<D�a<��a<Мa<�a<؜a<Ɯa<��a<L�a<�a<��a<:�a<ݚa<��a<��a<Q�a<>�a<A�a<I�a<B�a<W�a<2�a<�a<әa<��a< �a<r�a<˗a<�a<>�a<w�a<˔a<�a<��a<�a<��a<|�a<u�a<o�a<��a<��a<Ғa<��a<�a<��a<�a<��a<,�a<��a<)�a<v�a<ŏa<�a<V�a<��a<�a<��a<�a<��a<6�a<݊a<}�a<,�a<��a<�a<��a<·a<�a<��a<��a<�a<Ƃa<a<ƀa<�a<a<s~a< ~a<�}a<r}a<_}a<T}a<]}a<�}a<�}a<�}a<~}a<h}a<%}a<�|a<a|a<�{a<`{a<�za<[za<�ya<xya<2ya<�xa<�xa<�xa<�xa<�xa<�xa<�xa<�xa<cxa<<xa<�wa<nwa<�va<rva<�ua</ua<�ta<Ata<�sa<�sa<�sa<�sa<ta<hta<�ta<sua<$va<�  �  wa<�wa<xa<�xa<�xa<!ya<Aya<cya<Pya<Zya<Zya<vya<�ya<�ya<za<Qza<�za<h{a<|a<�|a<M}a<�}a<u~a<a<Ma<�a<�a<�a<�a<�a<�a<�a<J�a<��a<�a<��a<�a<�a<̓a<�a<�a<�a<�a<
�a<�a<يa<��a<4�a<ƌa<@�a<��a<��a<G�a<Ďa<�a<��a<6�a<Ɛa<��a<G�a<�a<��a<��a<>�a<ƕa<O�a<��a<ݖa<ߖa<�a<֖a<��a<��a<a�a<��a<p�a<��a<�a<H�a<їa<N�a<�a<��a<c�a<�a<~�a<��a<C�a<��a<��a<��a<��a<`�a<I�a<$�a< �a<�a<�a<�a<W�a<��a<Ԝa<,�a<i�a<ȝa<�a<�a<�a<ٝa<��a<?�a<�a<c�a<��a<z�a<��a<a<b�a<`�a<D�a<�a<��a< �a<l�a<��a<+�a<d�a<��a<ќa<�a<Ӝa<��a<d�a<�a<��a<,�a<ښa<��a<%�a<	�a<͙a<�a<ՙa<�a<�a<�a<
�a<�a<ԙa<v�a<�a<��a<�a<Z�a<��a<�a<�a<��a<�a<w�a<4�a<�a<��a<ƒa<��a<�a<�a<6�a<�a<�a<ڒa<��a<�a<��a<�a<�a<t�a<��a<�a<2�a<��a<�a<��a<D�a<ӊa<��a<�a<�a<|�a<��a<}�a<��a<�a<�a<0�a</�a< �a<3�a<�a<a�a<�a<�~a<h~a<~a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<�}a<[}a<'}a<�|a<4|a<�{a<{a<}za<�ya<�ya<�xa<�xa<kxa<Wxa<Sxa<@xa<Uxa<Uxa<{xa<mxa<Wxa<4xa<�wa<�wa<wa<�va<va<�ua<ua<�ta<nta<ta<,ta<(ta<�ta<�ta<Mua<�ua<bva<�  �  Ewa<�wa<7xa<}xa<�xa<�xa<ya<ya<ya<ya<�xa<�xa<ya<Cya<�ya<�ya<Vza<�za<�{a<X|a<}a<�}a<T~a<�~a<Pa<�a<�a<*�a<5�a<U�a<k�a<��a<��a<�a<w�a<�a<��a<d�a<X�a<I�a<>�a<V�a<S�a<G�a<�a<يa<��a<)�a<��a<�a<I�a<��a<�a<#�a<��a<#�a<��a<X�a<��a<�a<��a<��a<J�a<��a<��a<,�a<��a<Җa<�a<%�a<�a<�a<��a<�a<ܖa<�a</�a<l�a<×a<;�a<Ԙa<h�a<�a<��a<6�a<��a<�a<I�a<i�a<��a<Z�a<E�a<�a<�a<��a<��a<��a<��a<��a<ӛa<�a<z�a<͜a<*�a<r�a<��a<�a<��a<ٝa<��a<��a<&�a<��a<B�a<ߛa<u�a< �a<�a<ޚa<֚a<�a<�a<p�a<��a<�a<^�a<��a<Мa<Μa<ڜa<��a<k�a<�a<��a<A�a<Ϛa<E�a<��a<��a<��a<j�a<M�a<Z�a<��a<��a<��a<��a<˙a<��a<y�a<�a<��a<<�a<��a<�a<<�a<��a<�a<h�a<�a<��a<m�a<J�a<R�a<Q�a<P�a<n�a<k�a<[�a<�a<ڒa<x�a<�a<R�a<��a<ߏa<�a<G�a<a�a<��a<"�a<��a<�a<��a<p�a<*�a<�a<��a<>�a<�a<Z�a<Ça<�a<H�a<j�a<u�a<v�a<��a<��a<��a<�a<wa<�~a<�~a<K~a<3~a<~a<~a< ~a<~a<�}a<�}a<b}a<�|a<�|a<�{a<\{a<�za<'za<zya<�xa<�xa<8xa<�wa<�wa<�wa<�wa<�wa<xa<&xa<7xa<>xa<#xa<�wa<�wa<Zwa<�va<kva<�ua<�ua<ua<�ta<�ta<�ta<�ta<�ta<?ua<�ua<1va<�va<�  �  {wa<�wa<Axa<�xa<�xa<�xa<�xa<�xa<�xa<xxa<�xa<|xa<�xa<�xa<�xa<oya<�ya<�za<-{a<�{a<�|a<Z}a<~a<�~a<ba<�a<�a<P�a<x�a<��a<��a<�a<>�a<��a<��a<p�a<E�a<�a<�a<��a<��a<��a<��a<r�a<�a<�a<f�a<�a<J�a<��a<�a<�a<��a<��a<(�a<��a<�a<ݏa<��a<|�a<&�a<#�a<��a<��a<~�a<�a<Ŗa<��a<9�a<P�a<q�a<m�a<R�a<~�a<]�a<��a<��a<�a<b�a<��a<`�a<��a<m�a<ޚa<[�a<��a<�a<e�a<7�a<K�a<�a<�a<��a<m�a<Q�a<�a<�a<��a<�a<U�a<��a<�a<?�a<ٜa<�a<��a<��a<�a<	�a<Ɲa<��a<W�a<%�a<��a<U�a<�a<��a<��a<?�a<l�a<v�a<��a<�a<�a<y�a<��a<՜a<ٜa<��a<֜a<}�a<9�a<��a<d�a<��a<]�a<ߙa<x�a</�a<Ҙa<�a<˘a<��a<
�a< �a<s�a<q�a<��a<u�a<��a<)�a<ǘa<b�a<Ηa<U�a<��a<#�a<w�a<�a<��a<�a<�a<˓a<�a<��a<��a<Ǔa<��a<��a<(�a<�a<X�a<ɑa<�a<J�a<��a<|�a<ݍa<�a<F�a<��a<�a<��a<(�a<�a<��a<��a<G�a<��a<��a<3�a<�a<�a<p�a<��a<ʄa<ރa<�a<4�a<>�a<��a<�a<qa<)a<�~a<�~a<a~a<x~a<H~a<)~a<�}a<�}a<}}a<�|a<Y|a<�{a<{a<Gza<�ya<ya<gxa<xa<�wa<jwa<Uwa<Mwa<ywa<hwa<�wa<�wa<xa<xa<xa<xa<�wa<}wa<wa<�va<>va<�ua<�ua<Wua<Iua<
ua<Oua<wua<�ua<5va<�va<(wa<�  �  �wa<,xa<uxa<�xa<�xa<�xa<�xa<�xa<Wxa<(xa<xa<�wa<�wa<%xa<rxa<�xa<Mya<�ya<�za<z{a<\|a<*}a<�}a<�~a<0a<�a<<�a<��a<̀a<�a<C�a<��a<��a<�a<��a<�a<Ńa<h�a<H�a<7�a<�a<��a<ňa<��a<L�a<�a<R�a<ʋa<#�a<O�a<��a<��a<��a<-�a<��a<�a<��a<:�a<�a<�a<Ցa<��a<��a<��a<Y�a<��a<��a<
�a<u�a<��a<��a<ӗa<��a<�a<ܗa<�a<F�a<��a<ۘa<1�a<˙a<B�a<Úa<3�a<��a<��a<#�a<3�a<.�a<"�a<�a<��a<A�a< �a<��a<��a<j�a<z�a<��a<��a<�a<��a<�a<o�a<ޜa<]�a<��a<Ɲa<��a<��a<�a<��a<l�a< �a<Ӝa<j�a<+�a<�a<�a<��a<��a<�a<\�a<��a<ǜa<�a<�a<�a<��a<��a<q�a<�a<��a<��a<c�a<�a<T�a<�a<��a<o�a<J�a<C�a<g�a<��a<Ęa<�a<A�a<p�a<o�a<Y�a<D�a<�a<��a<"�a<��a<�a<��a<�a<��a<�a<Δa<��a<N�a<A�a<?�a<(�a<�a<ݓa<��a<X�a<�a<D�a<��a<�a<��a<�a<3�a<Q�a<j�a<��a<�a<�a<��a<��a<z�a<I�a<�a<��a<шa<��a<$�a<Ƈa<9�a<��a<څa<�a<E�a<q�a<��a<��a<#�a<��a<�a<�a<Aa<)a<�~a<�~a<�~a<g~a<4~a<�}a<K}a<�|a<1|a<w{a<�za<�ya<4ya<�xa<�wa<nwa<"wa<�va<�va<�va<�va<wa<[wa<�wa<�wa<�wa<�wa<xa<�wa<�wa<]wa<wa<�va<tva<va<�ua<�ua<�ua<�ua<�ua<2va<�va<wa<vwa<�  �  "xa<Zxa<�xa<�xa<�xa<�xa<kxa<Pxa<�wa<�wa<�wa<xwa<�wa<�wa<�wa<Axa<�xa<}ya<Wza<1{a<|a<�|a<�}a<�~a</a<�a<P�a<��a<!�a<O�a<��a<�a<J�a<��a<�a<��a<&�a<�a<��a<��a<V�a<C�a<�a<��a<x�a<�a<`�a<��a<�a<�a<%�a<i�a<l�a<Ōa<
�a<��a<�a<��a<��a<`�a<�a<a�a<j�a<V�a<-�a<�a<��a<1�a<��a<՗a<�a<�a<>�a<L�a<{�a<{�a<ǘa< �a<Q�a<љa<%�a<��a<��a<��a<՛a<�a<<�a<2�a<,�a<ߛa<��a<P�a<��a<��a<:�a<*�a<�a<��a<�a<L�a<��a<
�a<��a<�a<��a<�a<��a<ϝa<��a<"�a<	�a<��a<��a<k�a<)�a<�a<��a<u�a<x�a<[�a<��a<��a<��a<�a<�a<;�a<5�a<1�a<��a<��a<U�a<Ǜa<P�a<��a<�a<n�a<ܘa<|�a<�a<�a<��a<�a<�a<5�a<|�a<��a<�a<'�a<c�a<X�a<X�a<�a<јa<w�a<�a<y�a<�a<��a<��a<��a<R�a<�a<�a<��a<��a<i�a<[�a<$�a<ѓa<��a<�a<R�a<��a<��a<ɏa<��a<�a<Ȍa<�a<)�a<��a<��a<}�a<G�a<�a<�a<��a<��a<��a<`�a<0�a<a<`�a<��a<�a<e�a<�a<΃a<�a<\�a<��a<�a<��a<�a<�a<�a<\a<	a<�~a<�~a<?~a<�}a<K}a<�|a<�{a<B{a<hza<�ya<�xa<xa<�wa<�va<�va<Sva<Lva<Tva<vva<�va<�va<awa<�wa<�wa<�wa<xa<	xa<�wa<�wa<^wa<wa<�va<�va<kva<-va<Cva<>va<�va<�va<wa<_wa<�wa<�  �  Ixa<�xa<�xa<�xa<�xa<xa<Jxa<xa<�wa<hwa<Cwa<wa<wa<,wa<lwa<�wa<sxa<!ya<�ya<�za<�{a<�|a<�}a<i~a<4a<�a<`�a<�a<L�a<��a<��a<L�a<��a<��a<�a<�a<��a<]�a<#�a<�a<��a<��a<<�a<݉a<v�a<�a<:�a<��a<��a<ҋa<ыa<�a<�a<T�a<��a<�a<��a<R�a<.�a<�a<
�a<	�a<#�a<"�a<�a<ڕa<��a<5�a<��a<�a<W�a<m�a<��a<��a<Ҙa<��a<9�a<{�a<��a<(�a<��a<��a<\�a<��a<�a<�a<E�a<:�a<�a<ța<x�a<�a<��a<?�a<�a<��a<x�a<q�a<��a<�a<9�a<��a<1�a<Ǜa<m�a<�a<`�a<��a<�a<"�a<-�a<�a<	�a<��a<��a<T�a<�a<��a<�a<֜a<ݜa<�a<$�a<6�a<a�a<b�a<^�a<5�a<�a<��a<1�a<��a<�a<[�a<��a<�a<z�a<	�a<��a<h�a<U�a<h�a<��a<՗a<�a<t�a<Әa<�a<:�a<\�a<^�a<(�a<��a<��a<@�a<ɗa<S�a<ޖa<b�a<�a<ƕa<w�a<C�a<�a<��a<Ɣa<��a<T�a<�a<��a<�a<,�a<e�a<z�a<��a<g�a<l�a<y�a<��a<a<�a<�a<�a<Ԉa<��a<~�a<g�a<o�a<`�a<C�a<�a<Їa<c�a<نa<J�a<��a<߄a<$�a<g�a<��a<	�a<��a< �a<��a<8�a<�a<�a<ga<$a<�~a<W~a<�}a<S}a<�|a<�{a<	{a<za<7ya<txa<�wa<wa<|va<va<�ua<�ua<�ua<$va<Zva<�va< wa<mwa<�wa<�wa<xa<
xa<�wa<�wa<�wa<cwa<3wa<�va<�va<�va<�va<�va<�va<&wa<qwa<�wa<xa<�  �  fxa<�xa<�xa<�xa<�xa<uxa<1xa<�wa<�wa<3wa<wa<�va<�va<�va<wa<�wa<xa<�xa<�ya<�za<�{a<r|a<�}a<Z~a<*a<�a<��a<�a<p�a<�a<*�a<��a<�a<Z�a<ڃa<O�a<	�a<��a<r�a<.�a<�a<��a<X�a<�a<p�a<�a<'�a<��a<��a<��a<ċa<��a<�a<��a<H�a<��a<O�a<�a<Ŏa<׏a<ːa<��a<��a<��a<�a<ƕa<��a<0�a<їa<�a<l�a<��a<Ҙa<�a<�a<Z�a<z�a<̙a<�a<h�a<�a<-�a<��a<֛a<�a<F�a<C�a<1�a<�a<a<8�a<�a<n�a<��a<��a<@�a<:�a<#�a<O�a<�a<ޙa<~�a<��a<��a< �a<˜a<W�a<��a<�a<&�a<b�a<8�a<7�a<��a<؝a<��a<g�a<U�a<#�a<8�a<1�a<B�a<l�a<k�a<��a<�a<��a<?�a<�a<��a<'�a<��a<Śa<C�a<n�a<ݘa<%�a<��a<b�a<�a<�a<�a<B�a<��a<�a<S�a<��a<�a<+�a<R�a<]�a<I�a< �a<Ƙa<��a<��a<��a<�a<��a<g�a<��a<֕a<��a<l�a<6�a< �a<Ɣa<p�a<'�a<}�a<�a<�a<^�a<T�a<J�a<Z�a<-�a<>�a<-�a<f�a<��a<0�a<Ȉa<k�a<c�a<>�a<T�a<A�a<4�a<>�a<�a<هa<^�a<�a<b�a<Ņa<�a<b�a<��a<�a<l�a<Áa<Q�a<�a<x�a<@�a<�a<�a<@a<�~a<}~a<�}a<J}a<�|a<�{a<�za<�ya<ya<2xa<fwa<�va<>va<�ua<�ua<�ua<�ua<�ua<"va<�va<�va<Kwa<�wa<�wa<xa<xa<0xa<�wa<�wa<�wa<ywa<>wa<wa<wa<�va<wa<2wa<gwa<�wa<�wa<Fxa<�  �  �xa<�xa<�xa<�xa<�xa<nxa<xa<�wa<gwa<wa<�va<�va<�va<�va<�va<Swa<�wa<�xa<ya<sza<l{a<_|a<i}a<_~a<.a<�a<��a<�a<��a<�a<`�a<��a<,�a<��a<��a<��a<2�a<�a<��a<[�a<�a<؈a<}�a<�a<��a<��a<1�a<d�a<f�a<z�a<��a<��a<��a<ڋa< �a<z�a<�a<Ӎa<��a<��a<��a<��a<˒a<Փa<�a<ҕa<��a<F�a<ٗa<B�a<��a<ؘa<�a<1�a<e�a<��a<��a<�a<Q�a<��a<�a<b�a<��a<�a<5�a<R�a<V�a<4�a<��a<��a< �a<��a<@�a<șa<`�a<(�a<��a<�a<�a<[�a<��a<9�a<Қa<}�a<�a<��a<H�a<��a<�a<;�a<j�a<c�a<V�a<%�a<��a<ҝa<��a<y�a<]�a<]�a<��a<��a<��a<��a<��a<��a<��a<V�a<�a<��a<!�a<k�a<��a<�a<J�a<��a<��a<��a<�a<ݖa<Ζa<�a<�a<\�a<��a<�a<v�a<��a<0�a<V�a<l�a<X�a<.�a<��a<��a<1�a<×a<e�a<��a<��a<7�a< �a<ڕa<��a<d�a<-�a<�a<��a<.�a<��a<��a<"�a<C�a</�a<+�a<!�a< �a<��a<�a<>�a<y�a<�a<��a<T�a<�a<�a<�a<�a<�a<�a<��a<Շa<t�a<�a<��a<�a<I�a<��a<�a<F�a<��a<��a<s�a<�a<Àa<c�a<�a<�a<qa<a<�~a<�}a<M}a<�|a<�{a<�za<�ya<�xa<�wa<*wa<�va<�ua<�ua<Wua<\ua<lua<�ua<�ua<iva<�va<)wa<�wa<�wa<xa<"xa<8xa<xa<xa<�wa<�wa<uwa<gwa<1wa<(wa<@wa<�wa<�wa<�wa<xa<bxa<�  �  /wa<Nwa<]wa<<wa<wa<�va<+va<�ua<ua<�ta<#ta<�sa<�sa<�sa<�sa<<ta<�ta<�ua<�va<xa<4ya<�za<�{a<�|a<�}a<�~a<La<�a<Q�a<ŀa<#�a<��a<�a<0�a<��a<d�a<Ѓa<��a<r�a<4�a<�a<��a<[�a<��a<j�a<��a<�a<
�a<�a<Éa<i�a<i�a<I�a<?�a<��a<ˉa<]�a<A�a<&�a<S�a<��a<ďa<9�a<��a<��a<�a<��a<l�a<�a<s�a<��a<�a<3�a<b�a<}�a<��a<�a<&�a<[�a<љa<6�a<��a<�a<&�a<^�a<��a<`�a<5�a<��a<G�a<��a<�a<G�a<��a<�a<��a<\�a<B�a<f�a<Җa<O�a<
�a<טa<��a<��a<D�a<!�a<��a<�a<[�a<w�a<��a<i�a<K�a<"�a<�a<��a<s�a<��a<Y�a<l�a<��a<��a<��a<Ȝa<Ĝa<��a<p�a<�a<��a<��a<��a<.�a<�a<L�a<g�a<��a<��a<q�a<4�a<&�a<Z�a<��a<1�a<��a<P�a< �a<v�a<�a<O�a<e�a<x�a<J�a<	�a<��a<T�a<�a<w�a<�a<��a<k�a<�a<הa<��a<��a<\�a<�a<��a<P�a<��a<�a<*�a<�a<Ўa<��a<�a<�a<��a<~�a<��a<��a<+�a<�a<��a<��a<�a<�a<M�a<��a<��a<Ɇa<��a<I�a<��a<^�a<��a<+�a<`�a<��a<�a<0�a<΀a<=�a<�a<pa<#a<�~a<�~a<~a<�}a<D}a<�|a<�{a<{a<�ya<�xa<�wa<sva<nua<fta<�sa<�ra<qra<>ra<Xra<�ra<�ra<�sa<�sa<�ta<Fua<�ua<\va<�va<�va<�va<�va<�va<nva<Bva<va<�ua<�ua<�ua<�ua<�ua<8va<va<�va<�va<�  �  4wa<cwa<fwa<Zwa< wa<�va<-va<�ua<0ua<�ta<)ta<�sa<�sa<�sa<�sa<nta<ua<�ua<�va<xa<Mya<sza<�{a<�|a<�}a<�~a<Ka<�a<Y�a<��a<�a<f�a<��a<!�a<��a<�a<˃a<|�a<N�a<�a<�a<Ça<q�a<�a<z�a<щa<։a<�a<Ӊa<��a<��a<n�a<f�a<a�a<��a<�a<��a<\�a<C�a<r�a<��a<��a<8�a<o�a<��a<��a<��a<|�a<�a<��a<ݗa<�a<�a<B�a<P�a<��a<��a<�a<N�a<��a<�a<u�a<�a<8�a<v�a<|�a<p�a<<�a<��a<?�a<��a<�a<f�a<��a<8�a<��a<��a<|�a<��a<�a<p�a<�a<֘a<��a<��a<B�a<�a<��a<"�a<g�a<��a<��a<s�a<:�a<�a<��a<��a<`�a<;�a<A�a<N�a<\�a<��a<��a<Μa<ɜa<��a<y�a<$�a<}�a<a<��a<(�a<E�a<L�a<n�a<��a<�a<��a<c�a<X�a<s�a<єa<7�a<ϕa<j�a<�a<q�a<ۗa<G�a<y�a<w�a<`�a<�a<��a<<�a<˖a<A�a<�a<w�a<�a<�a<��a<��a<j�a<K�a< �a<ʓa<W�a<��a<�a<��a<�a<��a<��a<H�a<��a<ˉa<��a<��a<�a<p�a<�a<ʅa<مa<�a<!�a<L�a<o�a<��a<��a<��a<X�a<�a<v�a<ׄa<�a<D�a<��a<ǁa<+�a<��a<�a<�a<=a<a<�~a<~a</~a<�}a<?}a<�|a<�{a<�za<�ya<�xa<�wa<�va<uua<�ta<�sa<sa<�ra<|ra<mra<�ra<sa<�sa<&ta<�ta<Dua<�ua<8va<�va<�va<�va<�va<�va<^va<"va<�ua<�ua<�ua<�ua<�ua<�ua<va<cva<�va< wa<�  �  �va<?wa<@wa<Kwa<wa<�va<�va<�ua<cua<�ta<`ta<ta<�sa<�sa< ta<�ta<Iua<=va<!wa<Gxa<wya<�za<�{a<�|a<�}a<�~a<#a<�a<�a<��a<рa<5�a<m�a<�a<b�a<ނa<��a<3�a<�a<�a<��a<��a<3�a<؈a<S�a<̉a<�a<+�a<�a<Չa<Ӊa<��a<��a<��a<Ήa<D�a<Њa<��a<��a<��a<a<,�a<U�a<��a<�a<��a<��a<Y�a<�a<R�a<��a<ŗa<��a<�a<�a<U�a<o�a<��a<�a<^�a<�a<D�a<��a<��a<H�a<X�a<Y�a<<�a<ښa<��a<יa<8�a<��a<�a<|�a<��a<��a<��a<ۖa<�a<��a<P�a<��a<�a<��a<��a<(�a<��a<�a<<�a<k�a<O�a<D�a<��a<Ӝa<}�a<F�a<5�a<�a<�a<�a<�a<d�a<r�a<��a<��a<��a<S�a<�a<��a<��a<W�a<C�a<x�a<w�a<��a<��a<A�a<��a<��a<��a<��a<�a<j�a<��a<��a<�a<Ǘa< �a<O�a<g�a<O�a<5�a<ԗa<��a<�a<��a<�a<��a<H�a<�a<��a<l�a<_�a<A�a<�a<�a<��a<)�a<��a<��a<�a<2�a<�a<��a<�a<�a<�a<�a<�a<7�a<��a<3�a<�a<�a<
�a<Y�a<i�a<��a<ކa<��a<��a<6�a<Ʌa<=�a<��a<Ճa< �a<Z�a<~�a<��a<K�a<�a<ra<�~a<�~a<�~a<E~a<�}a<�}a<}a<�|a<�{a<�za<*za<�xa<�wa<�va<�ua<�ta<�sa<Ksa<�ra<�ra<�ra<�ra<@sa<�sa<Yta<�ta<�ua<�ua<Hva<�va<�va<�va<�va<qva<#va<�ua<�ua<pua<mua<Qua<|ua<�ua<�ua<3va<pva<�va<�  �  �va<#wa<Owa<2wa<wa<�va<wva<va<�ua<5ua<�ta<�ta<kta<qta<�ta<(ua<�ua<�va<�wa<�xa<�ya<�za<�{a<�|a<�}a<�~a<3a<�a<�a<I�a<��a<��a<�a<^�a<ρa<n�a<��a<�a<��a<��a<p�a<L�a<�a<ވa<b�a<��a<�a<�a<(�a<1�a<�a<
�a<��a<#�a<d�a<��a<J�a<!�a<�a<�a<;�a<d�a<��a<ɒa<֓a<�a<��a<g�a<��a<*�a<j�a<��a<��a<��a<×a<��a<��a<2�a<��a<�a<_�a<��a<n�a<Қa< �a<j�a<[�a<1�a<�a<{�a<�a<��a<�a<U�a<Ηa<{�a<F�a<)�a<S�a<��a<�a<��a<s�a<(�a<�a<��a<+�a<��a<��a<I�a<V�a<,�a<��a<��a<b�a<�a<�a<��a<��a<y�a<��a<Ûa<�a<#�a<W�a<i�a<y�a<a�a<��a<��a<�a<J�a<��a<��a<�a<�a<W�a<͕a<[�a<�a<�a<0�a<l�a<וa<T�a<ݖa<W�a<��a<&�a<N�a<_�a<_�a<�a<��a<@�a<��a<�a<��a<�a<��a<t�a< �a<!�a<��a<�a<˓a<��a<h�a</�a<��a<�a<5�a< �a<�a<��a<��a<��a<]�a<c�a<~�a<��a<�a<ˆa<��a<k�a<��a<��a<��a<Ɇa<Ɔa<ӆa<��a<C�a<؅a<�a<e�a<��a<΂a<ԁa<:�a<Y�a<�a<Ha<�~a<�~a<L~a<;~a<~a<�}a<{}a<-}a<�|a<�{a<{a<za<*ya<$xa<wa<va< ua<gta<�sa<Xsa<*sa<2sa<Rsa<�sa<ta<�ta<&ua<�ua<�ua<eva<�va<�va<�va<fva<)va<�ua<�ua<:ua<ua<�ta<�ta<�ta<,ua<iua<�ua<!va<�va<�  �  �va<�va<wa<"wa</wa<wa<�va<|va<�ua<�ua<Dua<ua<�ta<�ta<Iua<�ua<\va<wa<xa<ya<za<1{a<|a<}a<�}a<e~a<�~a<Da<�a<�a<1�a<1�a<��a<�a<G�a<�a<l�a<t�a< �a<'�a<�a<��a<͇a<��a<;�a<��a<:�a<D�a<k�a<��a<f�a<��a<s�a<��a<܊a<C�a<݋a<��a<��a<��a<a<Đa<�a<�a<�a<�a<��a<C�a<��a<�a<�a<�a<6�a<�a<N�a<(�a<r�a<��a<�a<��a<ؘa<��a<�a<��a<ɚa<�a<>�a<2�a<.�a<��a<f�a<ؙa<H�a<ݘa<O�a<�a<a<ʗa<ԗa<.�a<��a<-�a<�a<z�a<R�a<Ûa<]�a<Ӝa<�a<�a<��a<�a<��a<[�a<�a<|�a<q�a<�a<�a<�a<-�a</�a<r�a<қa<�a<$�a<�a<-�a<�a<��a<6�a<z�a<�a<�a<O�a<��a<ږa<V�a<ڕa<��a<��a<��a<�a<Z�a<��a<+�a<��a<�a<Q�a<N�a<E�a<�a<��a<e�a<a<a�a<��a<'�a<��a<-�a<�a<��a<��a<I�a<{�a<_�a<M�a<&�a<Ւa<��a<ܑa<Y�a<K�a<V�a<b�a<�a<�a<؊a<��a<��a<7�a<��a<C�a<�a<�a<
�a<��a<%�a<�a<�a<��a<|�a< �a<}�a<̄a<�a<"�a<b�a<B�a<ŀa<�a<Ma<�~a<_~a<0~a<�}a<�}a<�}a<z}a<#}a<�|a<o|a<�{a<I{a<Hza<�ya<yxa<twa<�va<�ua<�ta<Lta<�sa<�sa<�sa<�sa<ta<�ta<�ta<�ua<�ua<0va<}va<tva<�va<Hva<va<�ua<ua<ua<�ta<�ta<>ta<Zta<Nta<�ta<�ta<Aua<�ua<va<�  �  ?va<�va<�va<0wa<-wa<.wa< wa<�va<wva<va<�ua<�ua<�ua<�ua<�ua<]va< wa<�wa<�xa<�ya<{za<U{a<f|a<}a<�}a<g~a<�~a<a<Ua<Pa<�a<�a<�a<3�a<��a<,�a<сa<��a<��a<��a<n�a<��a<��a<\�a<�a<��a<"�a<��a<��a<Ŋa<�a<��a<�a<I�a<��a<�a<��a<I�a</�a<+�a<'�a<Q�a<O�a<U�a<d�a<��a<��a<#�a<p�a<��a<��a<��a<��a<�a<r�a<��a<��a<��a<_�a<��a<g�a< �a<o�a<+�a<��a<�a<5�a<F�a<$�a<�a<��a<9�a<ؙa<S�a<��a<��a<u�a<p�a<��a<�a<H�a<Ǚa<V�a<�a<v�a<�a<��a<ǜa<�a<�a<לa<��a<'�a<��a<t�a<�a<��a<k�a<U�a<J�a<h�a<��a<��a<1�a<r�a<ԛa<��a< �a<��a<��a<X�a<Қa<�a<��a<̘a<�a<��a< �a<��a<Y�a<H�a<d�a<��a<ߖa<G�a<��a<֗a<E�a<U�a<]�a<G�a<�a<��a<�a<G�a<��a<&�a<h�a<�a<z�a<3�a<�a<Ӓa<Вa<�a<ɒa<�a<�a<��a<W�a<�a<A�a<��a<��a<��a<��a<y�a<��a<��a<��a<��a<f�a<�a<��a<��a<o�a<}�a<d�a<U�a<T�a<�a<��a< �a<Q�a<��a<��a<��a<ҁa<΀a<�a<1a<�~a<~a<�}a<^}a<T}a<?}a<}a<"}a<�|a<�|a<f|a<�{a<?{a<�za<�ya<�xa<xa<wa<Lva<�ua< ua<�ta<ita<fta<�ta<�ta<ua<qua<�ua<va<gva<qva<�va<Zva<&va<�ua<Tua<�ta<�ta<ta<�sa<�sa<�sa<�sa<�sa<>ta<�ta</ua<�ua<�  �  �ua<qva<�va<"wa<Lwa<Ewa<Swa<wa<wa<�va<rva<Sva<Kva<ova<�va<(wa<�wa<gxa<#ya<za<{a<�{a<�|a<0}a<�}a<C~a<�~a<�~a<�~a<a<�~a<a<1a<�a<�a<c�a</�a<�a<�a<܃a<�a<7�a<�a<?�a<�a<ىa<8�a<Ȋa<�a<K�a<��a<s�a<ŋa<�a<Y�a<��a<H�a<�a<Ύa<ԏa<��a<��a<Ӓa<��a<��a<�a<ؕa<��a<U�a<A�a<Q�a<6�a<�a<�a<Õa<�a<��a<:�a<��a<�a<Ηa<O�a<9�a<��a<N�a<Κa<	�a<i�a<9�a<T�a<�a<Ța<R�a<ߙa<��a<K�a<E�a<#�a<M�a<��a<�a<h�a<њa<��a<�a<l�a<��a<�a<�a<��a<��a<&�a<�a<6�a<��a<W�a<�a<��a<��a<��a<��a<��a<G�a<��a<5�a<b�a<ƛa<ʛa<�a<ɛa<o�a<%�a<��a<�a<C�a<��a<*�a<��a<X�a<
�a<�a<�a<@�a<m�a<��a<+�a<<�a<��a<i�a<��a<$�a<ȗa<K�a<��a<�a<�a<��a<Ǔa<H�a<Œa<j�a<Q�a<�a<7�a<0�a<l�a<��a<t�a<��a<)�a<�a<W�a<ϐa<�a<�a<6�a<��a<*�a<#�a<s�a<��a<�a<��a<U�a<:�a<�a<�a<�a<��a<��a<��a<��a<ԅa<6�a<,�a<L�a<F�a<�a<9�a<:a<�~a<�}a<P}a<}a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<:|a<|a<T{a<�za<za<hya<~xa<�wa<�va<6va<�ua<Qua<$ua<ua<ua<Xua<~ua<va<&va<ova<�va<�va<�va<$va<�ua<aua<ua<Zta<�sa<zsa<sa<�ra<�ra<�ra<2sa<�sa<ta<�ta<gua<�  �  dua< va<�va<wa<_wa<ywa<�wa<�wa<@wa<.wa<#wa<�va<�va< wa<qwa<�wa<Yxa<ya<�ya<|za<V{a<+|a<�|a<c}a<�}a<,~a<|~a<�~a<j~a<�~a<k~a<x~a<�~a<�~a<'a<�a<_�a<E�a<H�a<T�a<��a<��a<��a<��a<Јa<��a<f�a<�a<Y�a<��a<ŋa<)�a<]�a<��a< �a<q�a<
�a<��a<z�a<h�a<g�a<)�a<:�a<�a<��a<E�a<��a<ޕa<�a<�a<̕a<��a<`�a<B�a<"�a<�a<B�a<��a<�a<~�a<%�a<͗a<��a<:�a<��a<��a<��a<U�a<h�a<s�a<]�a<�a<��a<��a<;�a<�a<�a<�a<��a<C�a<��a<�a<v�a<̛a<\�a<��a<ܜa<��a<ߜa<��a<^�a<��a<O�a<Ěa<,�a<��a<E�a<��a<Ϙa<֘a<�a<S�a<��a<)�a<��a<��a<v�a<��a<͛a<ܛa<��a<_�a<��a<V�a<ޙa<h�a<ɘa<a�a<
�a<ޗa<��a<��a<ۗa<)�a<2�a<t�a<��a<��a<��a<z�a<�a<��a<��a<"�a<z�a<��a<ޓa<+�a<��a<�a<��a<��a<}�a<��a<��a<�a<�a<�a<P�a<�a<�a<��a<�a<D�a<��a<q�a<��a<��a<ˋa<�a<e�a<ىa<f�a<�a<ψa<��a<V�a<N�a<�a<��a<*�a<��a<��a< �a<׃a<ǂa<��a<��a<�a<�~a<�}a<}a<�|a<L|a<|a<|a<|a<7|a<1|a<T|a<j|a<&|a<�{a<�{a<{a<wza<�ya<�xa<[xa<�wa<�va<rva<va<�ua<�ua<�ua<va<"va<;va<�va<�va<�va<�va<eva<va<�ua<�ta<|ta<�sa<Msa<�ra<pra<,ra<ra<;ra<�ra<�ra<�sa<(ta<�ta<�  �  <ua<�ua<�va<�va<Twa<�wa<�wa<�wa<�wa<�wa<�wa<�wa<�wa<�wa<*xa<lxa<-ya<�ya<^za<{a<�{a<v|a<�|a<�}a<�}a<<~a<=~a</~a<F~a<�}a<�}a<�}a<�}a<~a<i~a<a<�a<��a<��a<�a< �a<S�a<��a<��a<ވa<��a<t�a<�a<��a<�a<E�a<ƌa<Όa<d�a<��a<(�a<a<Z�a<V�a<ܐa<��a<��a<��a<=�a<ܔa<`�a<��a<�a<��a<��a<��a<�a<��a<��a<��a<k�a<��a<Ȕa<=�a<ԕa<�a<d�a<�a<�a<��a<U�a<�a<=�a<��a<��a<��a<~�a<R�a<$�a<��a<ښa<��a<��a<��a<��a<=�a<��a<�a<G�a<��a<՜a<�a<��a<Ԝa<��a<��a<��a<ܚa<9�a<��a<�a<��a<8�a<+�a<�a<`�a<��a<�a<��a<%�a<Кa<�a<��a<ța<Лa<Лa<��a<J�a<˚a<~�a<ۙa<i�a<#�a<��a<��a<W�a<��a<_�a<��a<Әa<ߘa<��a<٘a<ǘa<d�a<�a<j�a<��a<��a<�a<,�a<@�a<~�a<ۑa<O�a<�a<Ґa<ڐa<�a<9�a<[�a<��a<�a<�a<#�a<ӑa<��a<�a<v�a<ۏa<��a<O�a<2�a<��a<��a<�a<��a<�a<݉a<B�a<F�a<܈a<��a<=�a<̇a<E�a<y�a<Ѕa<��a<��a<��a<.�a<'�a<�~a<�}a<}a<h|a<�{a<�{a<t{a<l{a<�{a<�{a<|a<|a<|a<;|a<�{a<�{a<2{a<�za<za<~ya<�xa<xa<�wa<wa<�va<�va<�va<tva<qva<�va<�va<�va<�va<�va<�va<[va<va<Kua<�ta<	ta<]sa<�ra<*ra<�qa<qqa<wqa<~qa<�qa<Ora<�ra<�sa<Xta<�  �  �ta<�ua<[va<�va<gwa<�wa<	xa<xa<+xa<xa<xa<$xa<<xa<Rxa<�xa<�xa<�ya<!za<�za<v{a<%|a<�|a<X}a<�}a<�}a< ~a<~a<�}a<�}a<�}a<�}a<`}a<f}a<�}a<�}a<f~a<3a<�a<�a<Z�a<��a<��a<@�a<j�a<��a<��a<��a<f�a<�a<`�a<ǌa<(�a<X�a<�a<"�a<��a<F�a<�a<ΐa<l�a<i�a<,�a<�a<��a<6�a<��a<��a<ȕa<��a<e�a< �a<��a<q�a<�a<��a<�a<��a<C�a<a<U�a<�a<�a<��a<��a<o�a<*�a<�a<E�a<��a<��a<�a<ܛa<��a<��a<Q�a<Q�a<�a<1�a<9�a<s�a<ʛa<�a<f�a<a<��a<.�a<E�a<�a<Мa<p�a<̛a<<�a<��a<ҙa<�a<��a<�a<��a<��a<��a<ӗa<%�a<��a<=�a<ՙa<m�a<�a<m�a<��a<�a<�a<ܛa<��a<A�a<Κa<V�a<��a<��a<<�a<�a<�a<�a<��a<�a<-�a<C�a<?�a<7�a<�a<p�a<�a<:�a<m�a<��a<��a<��a<ƒa<��a<]�a<ΐa<l�a<U�a<R�a<e�a<��a<��a<T�a<��a<��a<��a<ґa<��a<l�a<ːa<-�a<s�a<��a<��a<"�a<;�a<��a<�a<��a<U�a<҉a<��a<Y�a< �a<��a<&�a<h�a<|�a<��a<p�a<P�a<�a<̀a<�a<i~a<u}a<�|a<�{a<Z{a<{a<�za<�za<'{a<S{a<�{a<�{a<�{a<|a<�{a<�{a<�{a< {a<|za<�ya<Iya<�xa<<xa<�wa<_wa<wa<�va<wa<�va<wa<1wa<2wa<0wa<wa<�va<Wva<�ua<ua<xta<�sa<�ra<@ra<�qa<<qa<�pa<�pa<�pa<Wqa<�qa<qra<<sa<ta<�  �  �ta<�ua<Dva<�va<|wa<�wa<'xa<<xa<sxa<mxa<�xa<}xa<�xa<�xa<"ya<�ya<�ya<�za<7{a<�{a<n|a<�|a<e}a<�}a<�}a<�}a<~a<�}a<�}a<k}a<}a< }a<�|a<
}a<o}a<�}a<�~a<�a<̀a<�a<Y�a<��a<�a<��a<��a<��a<��a<U�a<�a<��a<�a<q�a<ލa<*�a<��a<4�a<ŏa<��a<�a<�a<��a<g�a<%�a<��a<$�a<w�a<��a<��a<��a<A�a<ϔa<��a<��a<Ɠa<u�a<\�a<w�a<˓a<.�a<ݔa<��a<s�a<��a<N�a<d�a<6�a<��a<e�a<��a<��a<
�a<#�a<��a<�a<ʛa<��a<��a<��a<ϛa<��a<�a<��a<��a<�a<�a<O�a<7�a<�a<̜a<P�a<�a<��a<H�a<v�a<��a<)�a<��a<B�a<�a< �a<J�a<Ǘa<9�a<֘a<��a<&�a<��a<V�a<��a<��a<��a<��a<��a<��a<�a<Ԛa<T�a<�a<ؙa<��a<��a<_�a<g�a<��a<{�a<��a<b�a<E�a<�a<��a<ޗa<;�a<k�a<?�a<b�a<C�a<f�a<��a<ʐa<U�a<�a<ˏa<Ϗa<�a<;�a<��a<�a<h�a<ӑa<ˑa<�a<��a<[�a<��a<^�a<��a<��a<B�a<i�a<ڌa<'�a<��a</�a<��a<X�a<��a<��a<9�a<��a<�a<\�a<��a<v�a<��a<,�a<ʁa<��a<%a<~a<�|a<|a<S{a<�za<�za<|za<�za<�za<{a<E{a<�{a<�{a<�{a<|a<�{a<�{a<#{a<�za<*za<�ya<ya<�xa<?xa<�wa<�wa<ywa<Uwa<rwa<awa<swa<Uwa<Qwa<wa<�va<Sva<�ua<0ua<5ta<usa<�ra<�qa<Mqa<�pa<|pa<Npa<�pa<�pa<nqa<	ra<�ra<�sa<�  �  uta<Lua<va<�va<�wa<�wa<Mxa<xxa<�xa<�xa<�xa<�xa<�xa<ya<Xya<�ya<:za<�za<e{a<|a<�|a<}a<�}a<�}a<~a<�}a<�}a<�}a<q}a<8}a<�|a<�|a<�|a<�|a<:}a<�}a<t~a<Xa<��a<��a<%�a<��a<߅a<0�a<r�a<��a<��a<y�a<9�a<ǌa<C�a<��a<�a<j�a<�a<d�a<��a<��a<W�a<(�a<ےa<��a<X�a<�a<M�a<��a<��a<��a<W�a<�a<��a<K�a<Гa<��a<4�a<.�a<K�a<��a<��a<��a<q�a<N�a<L�a<8�a<�a<�a<��a<j�a<֛a< �a<F�a<V�a<<�a<�a<�a<�a<�a<؛a<��a</�a<Z�a<��a<�a<7�a<\�a<x�a<_�a<-�a<a<'�a<��a<ךa<�a<J�a<�a<�a<R�a<�a<זa<�a<�a<��a<�a<��a<e�a<	�a<��a<&�a<��a<�a<�a< �a<�a<��a<W�a<�a<��a<K�a<�a<řa<��a<��a<��a<��a<��a<��a<��a<i�a<�a<��a<͗a<��a<�a<*�a</�a<�a<.�a<N�a<��a< �a<a<��a<��a<ҏa<�a<��a<�a<8�a<��a<��a<�a<őa<�a<$�a<��a<�a<&�a<x�a<��a<�a<X�a<ȋa<^�a<ފa<��a<#�a<ԉa<m�a<�a<>�a<|�a<��a<g�a<8�a<�a<��a<\�a<�~a<�}a<�|a<�{a<'{a<�za<Vza<:za<^za<�za<�za<.{a<u{a<�{a<�{a<|a<�{a<�{a<_{a<�za<gza<�ya<Rya<�xa<lxa<xa<�wa<�wa<�wa<�wa<�wa<�wa<�wa<{wa<3wa<�va<Iva<�ua<�ta<ta<Gsa<nra<�qa<	qa<~pa<>pa<$pa<Ipa<�pa<*qa<�qa<�ra<�sa<�  �  }ta<Kua<Lva<�va<pwa<�wa<7xa<txa<�xa<�xa<�xa<�xa<ya<4ya<�ya<�ya<_za<�za<�{a<|a<�|a<}a<w}a<�}a<�}a<~a<~a<�}a<x}a<}a<�|a<�|a<�|a<�|a<�|a<}}a<M~a<?a<e�a<��a<��a<~�a<�a<;�a<��a<��a<��a<�a<#�a<��a<P�a<��a<2�a<��a<��a<��a<C�a<��a<��a<I�a<��a<��a<=�a<Ҕa<T�a<��a<��a<��a<j�a<�a<��a<�a<˓a<g�a<�a<�a<�a<T�a<�a<v�a<X�a<G�a<�a<@�a<)�a<�a<��a<H�a<ɛa<�a<4�a<<�a<K�a<<�a<+�a<�a<�a<'�a<#�a<A�a<��a<˜a<�a<7�a<W�a<c�a<_�a<�a<Ϝa<c�a<��a<�a<��a<=�a<y�a<ėa<;�a<Ӗa<��a<��a<��a<d�a<��a<��a<?�a<�a<��a<^�a<��a<�a<�a<
�a<�a<��a<l�a<�a<ƚa<d�a<�a<�a<Ùa<ęa<ҙa<әa<șa<��a<��a<W�a<�a<v�a<��a<0�a<$�a<1�a<��a<�a<�a<,�a<�a<��a<��a<n�a<w�a<��a<�a<Z�a<ڐa<K�a<��a<�a<ԑa<��a<��a<�a<}�a<��a<=�a<��a<ލa<�a<��a<�a<f�a<�a<��a<=�a<�a<R�a<҈a<D�a<j�a<|�a<��a<L�a<	�a<��a<.�a<�~a<�}a<�|a<�{a<�za<kza<;za<za<Dza<�za<�za<6{a<�{a<�{a<|a<�{a<�{a<�{a<N{a<�za<vza<�ya<{ya<�xa<txa<Uxa<�wa<�wa<�wa<�wa<�wa<�wa<�wa<ewa<3wa<�va<Vva<�ua<�ta< ta<*sa<bra<�qa<�pa<gpa<pa<�oa<pa<�pa<qa<�qa<�ra<rsa<�  �  uta<Lua<va<�va<�wa<�wa<Mxa<xxa<�xa<�xa<�xa<�xa<�xa<ya<Xya<�ya<:za<�za<e{a<|a<�|a<}a<�}a<�}a<~a<�}a<�}a<�}a<q}a<8}a<�|a<�|a<�|a<�|a<:}a<�}a<t~a<Xa<��a<��a<%�a<��a<߅a<0�a<r�a<��a<��a<y�a<9�a<ǌa<C�a<��a<�a<j�a<�a<d�a<��a<��a<W�a<(�a<ےa<��a<X�a<�a<M�a<��a<��a<��a<W�a<�a<��a<K�a<Гa<��a<4�a<.�a<K�a<��a<��a<��a<q�a<N�a<L�a<8�a<�a<�a<��a<j�a<֛a< �a<F�a<V�a<<�a<�a<�a<�a<�a<؛a<��a</�a<Z�a<��a<�a<7�a<\�a<x�a<_�a<-�a<a<'�a<��a<ךa<�a<J�a<�a<�a<R�a<�a<זa<�a<�a<��a<�a<��a<e�a<	�a<��a<&�a<��a<�a<�a< �a<�a<��a<W�a<�a<��a<K�a<�a<řa<��a<��a<��a<��a<��a<��a<��a<i�a<�a<��a<͗a<��a<�a<*�a</�a<�a<.�a<N�a<��a< �a<a<��a<��a<ҏa<�a<��a<�a<8�a<��a<��a<�a<őa<�a<$�a<��a<�a<&�a<x�a<��a<�a<X�a<ȋa<^�a<ފa<��a<#�a<ԉa<m�a<�a<>�a<|�a<��a<g�a<8�a<�a<��a<\�a<�~a<�}a<�|a<�{a<'{a<�za<Vza<:za<^za<�za<�za<.{a<u{a<�{a<�{a<|a<�{a<�{a<_{a<�za<gza<�ya<Rya<�xa<lxa<xa<�wa<�wa<�wa<�wa<�wa<�wa<�wa<{wa<3wa<�va<Iva<�ua<�ta<ta<Gsa<nra<�qa<	qa<~pa<>pa<$pa<Ipa<�pa<*qa<�qa<�ra<�sa<�  �  �ta<�ua<Dva<�va<|wa<�wa<'xa<<xa<sxa<mxa<�xa<}xa<�xa<�xa<"ya<�ya<�ya<�za<7{a<�{a<n|a<�|a<e}a<�}a<�}a<�}a<~a<�}a<�}a<k}a<}a< }a<�|a<
}a<o}a<�}a<�~a<�a<̀a<�a<Y�a<��a<�a<��a<��a<��a<��a<U�a<�a<��a<�a<q�a<ލa<*�a<��a<4�a<ŏa<��a<�a<�a<��a<g�a<%�a<��a<$�a<w�a<��a<��a<��a<A�a<ϔa<��a<��a<Ɠa<u�a<\�a<w�a<˓a<.�a<ݔa<��a<s�a<��a<N�a<d�a<6�a<��a<e�a<��a<��a<
�a<#�a<��a<�a<ʛa<��a<��a<��a<ϛa<��a<�a<��a<��a<�a<�a<O�a<7�a<�a<̜a<P�a<�a<��a<H�a<v�a<��a<)�a<��a<B�a<�a< �a<J�a<Ǘa<9�a<֘a<��a<&�a<��a<V�a<��a<��a<��a<��a<��a<��a<�a<Ԛa<T�a<�a<ؙa<��a<��a<_�a<g�a<��a<{�a<��a<b�a<E�a<�a<��a<ޗa<;�a<k�a<?�a<b�a<C�a<f�a<��a<ʐa<U�a<�a<ˏa<Ϗa<�a<;�a<��a<�a<h�a<ӑa<ˑa<�a<��a<[�a<��a<^�a<��a<��a<B�a<i�a<ڌa<'�a<��a</�a<��a<X�a<��a<��a<9�a<��a<�a<\�a<��a<v�a<��a<,�a<ʁa<��a<%a<~a<�|a<|a<S{a<�za<�za<|za<�za<�za<{a<E{a<�{a<�{a<�{a<|a<�{a<�{a<#{a<�za<*za<�ya<ya<�xa<?xa<�wa<�wa<ywa<Uwa<rwa<awa<swa<Uwa<Qwa<wa<�va<Sva<�ua<0ua<5ta<usa<�ra<�qa<Mqa<�pa<|pa<Npa<�pa<�pa<nqa<	ra<�ra<�sa<�  �  �ta<�ua<[va<�va<gwa<�wa<	xa<xa<+xa<xa<xa<$xa<<xa<Rxa<�xa<�xa<�ya<!za<�za<v{a<%|a<�|a<X}a<�}a<�}a< ~a<~a<�}a<�}a<�}a<�}a<`}a<f}a<�}a<�}a<f~a<3a<�a<�a<Z�a<��a<��a<@�a<j�a<��a<��a<��a<f�a<�a<`�a<ǌa<(�a<X�a<�a<"�a<��a<F�a<�a<ΐa<l�a<i�a<,�a<�a<��a<6�a<��a<��a<ȕa<��a<e�a< �a<��a<q�a<�a<��a<�a<��a<C�a<a<U�a<�a<�a<��a<��a<o�a<*�a<�a<E�a<��a<��a<�a<ܛa<��a<��a<Q�a<Q�a<�a<1�a<9�a<s�a<ʛa<�a<f�a<a<��a<.�a<E�a<�a<Мa<p�a<̛a<<�a<��a<ҙa<�a<��a<�a<��a<��a<��a<ӗa<%�a<��a<=�a<ՙa<m�a<�a<m�a<��a<�a<�a<ܛa<��a<A�a<Κa<V�a<��a<��a<<�a<�a<�a<�a<��a<�a<-�a<C�a<?�a<7�a<�a<p�a<�a<:�a<m�a<��a<��a<��a<ƒa<��a<]�a<ΐa<l�a<U�a<R�a<e�a<��a<��a<T�a<��a<��a<��a<ґa<��a<l�a<ːa<-�a<s�a<��a<��a<"�a<;�a<��a<�a<��a<U�a<҉a<��a<Y�a< �a<��a<&�a<h�a<|�a<��a<p�a<P�a<�a<̀a<�a<i~a<u}a<�|a<�{a<Z{a<{a<�za<�za<'{a<S{a<�{a<�{a<�{a<|a<�{a<�{a<�{a< {a<|za<�ya<Iya<�xa<<xa<�wa<_wa<wa<�va<wa<�va<wa<1wa<2wa<0wa<wa<�va<Wva<�ua<ua<xta<�sa<�ra<@ra<�qa<<qa<�pa<�pa<�pa<Wqa<�qa<qra<<sa<ta<�  �  <ua<�ua<�va<�va<Twa<�wa<�wa<�wa<�wa<�wa<�wa<�wa<�wa<�wa<*xa<lxa<-ya<�ya<^za<{a<�{a<v|a<�|a<�}a<�}a<<~a<=~a</~a<F~a<�}a<�}a<�}a<�}a<~a<i~a<a<�a<��a<��a<�a< �a<S�a<��a<��a<ވa<��a<t�a<�a<��a<�a<E�a<ƌa<Όa<d�a<��a<(�a<a<Z�a<V�a<ܐa<��a<��a<��a<=�a<ܔa<`�a<��a<�a<��a<��a<��a<�a<��a<��a<��a<k�a<��a<Ȕa<=�a<ԕa<�a<d�a<�a<�a<��a<U�a<�a<=�a<��a<��a<��a<~�a<R�a<$�a<��a<ښa<��a<��a<��a<��a<=�a<��a<�a<G�a<��a<՜a<�a<��a<Ԝa<��a<��a<��a<ܚa<9�a<��a<�a<��a<8�a<+�a<�a<`�a<��a<�a<��a<%�a<Кa<�a<��a<ța<Лa<Лa<��a<J�a<˚a<~�a<ۙa<i�a<#�a<��a<��a<W�a<��a<_�a<��a<Әa<ߘa<��a<٘a<ǘa<d�a<�a<j�a<��a<��a<�a<,�a<@�a<~�a<ۑa<O�a<�a<Ґa<ڐa<�a<9�a<[�a<��a<�a<�a<#�a<ӑa<��a<�a<v�a<ۏa<��a<O�a<2�a<��a<��a<�a<��a<�a<݉a<B�a<F�a<܈a<��a<=�a<̇a<E�a<y�a<Ѕa<��a<��a<��a<.�a<'�a<�~a<�}a<}a<h|a<�{a<�{a<t{a<l{a<�{a<�{a<|a<|a<|a<;|a<�{a<�{a<2{a<�za<za<~ya<�xa<xa<�wa<wa<�va<�va<�va<tva<qva<�va<�va<�va<�va<�va<�va<[va<va<Kua<�ta<	ta<]sa<�ra<*ra<�qa<qqa<wqa<~qa<�qa<Ora<�ra<�sa<Xta<�  �  dua< va<�va<wa<_wa<ywa<�wa<�wa<@wa<.wa<#wa<�va<�va< wa<qwa<�wa<Yxa<ya<�ya<|za<V{a<+|a<�|a<c}a<�}a<,~a<|~a<�~a<j~a<�~a<k~a<x~a<�~a<�~a<'a<�a<_�a<E�a<H�a<T�a<��a<��a<��a<��a<Јa<��a<f�a<�a<Y�a<��a<ŋa<)�a<]�a<��a< �a<q�a<
�a<��a<z�a<h�a<g�a<)�a<:�a<�a<��a<E�a<��a<ޕa<�a<�a<̕a<��a<`�a<B�a<"�a<�a<B�a<��a<�a<~�a<%�a<͗a<��a<:�a<��a<��a<��a<U�a<h�a<s�a<]�a<�a<��a<��a<;�a<�a<�a<�a<��a<C�a<��a<�a<v�a<̛a<\�a<��a<ܜa<��a<ߜa<��a<^�a<��a<O�a<Ěa<,�a<��a<E�a<��a<Ϙa<֘a<�a<S�a<��a<)�a<��a<��a<v�a<��a<͛a<ܛa<��a<_�a<��a<V�a<ޙa<h�a<ɘa<a�a<
�a<ޗa<��a<��a<ۗa<)�a<2�a<t�a<��a<��a<��a<z�a<�a<��a<��a<"�a<z�a<��a<ޓa<+�a<��a<�a<��a<��a<}�a<��a<��a<�a<�a<�a<P�a<�a<�a<��a<�a<D�a<��a<q�a<��a<��a<ˋa<�a<e�a<ىa<f�a<�a<ψa<��a<V�a<N�a<�a<��a<*�a<��a<��a< �a<׃a<ǂa<��a<��a<�a<�~a<�}a<}a<�|a<L|a<|a<|a<|a<7|a<1|a<T|a<j|a<&|a<�{a<�{a<{a<wza<�ya<�xa<[xa<�wa<�va<rva<va<�ua<�ua<�ua<va<"va<;va<�va<�va<�va<�va<eva<va<�ua<�ta<|ta<�sa<Msa<�ra<pra<,ra<ra<;ra<�ra<�ra<�sa<(ta<�ta<�  �  �ua<qva<�va<"wa<Lwa<Ewa<Swa<wa<wa<�va<rva<Sva<Kva<ova<�va<(wa<�wa<gxa<#ya<za<{a<�{a<�|a<0}a<�}a<C~a<�~a<�~a<�~a<a<�~a<a<1a<�a<�a<c�a</�a<�a<�a<܃a<�a<7�a<�a<?�a<�a<ىa<8�a<Ȋa<�a<K�a<��a<s�a<ŋa<�a<Y�a<��a<H�a<�a<Ύa<ԏa<��a<��a<Ӓa<��a<��a<�a<ؕa<��a<U�a<A�a<Q�a<6�a<�a<�a<Õa<�a<��a<:�a<��a<�a<Ηa<O�a<9�a<��a<N�a<Κa<	�a<i�a<9�a<T�a<�a<Ța<R�a<ߙa<��a<K�a<E�a<#�a<M�a<��a<�a<h�a<њa<��a<�a<l�a<��a<�a<�a<��a<��a<&�a<�a<6�a<��a<W�a<�a<��a<��a<��a<��a<��a<G�a<��a<5�a<b�a<ƛa<ʛa<�a<ɛa<o�a<%�a<��a<�a<C�a<��a<*�a<��a<X�a<
�a<�a<�a<@�a<m�a<��a<+�a<<�a<��a<i�a<��a<$�a<ȗa<K�a<��a<�a<�a<��a<Ǔa<H�a<Œa<j�a<Q�a<�a<7�a<0�a<l�a<��a<t�a<��a<)�a<�a<W�a<ϐa<�a<�a<6�a<��a<*�a<#�a<s�a<��a<�a<��a<U�a<:�a<�a<�a<�a<��a<��a<��a<��a<ԅa<6�a<,�a<L�a<F�a<�a<9�a<:a<�~a<�}a<P}a<}a<�|a<�|a<�|a<�|a<�|a<�|a<�|a<:|a<|a<T{a<�za<za<hya<~xa<�wa<�va<6va<�ua<Qua<$ua<ua<ua<Xua<~ua<va<&va<ova<�va<�va<�va<$va<�ua<aua<ua<Zta<�sa<zsa<sa<�ra<�ra<�ra<2sa<�sa<ta<�ta<gua<�  �  ?va<�va<�va<0wa<-wa<.wa< wa<�va<wva<va<�ua<�ua<�ua<�ua<�ua<]va< wa<�wa<�xa<�ya<{za<U{a<f|a<}a<�}a<g~a<�~a<a<Ua<Pa<�a<�a<�a<3�a<��a<,�a<сa<��a<��a<��a<n�a<��a<��a<\�a<�a<��a<"�a<��a<��a<Ŋa<�a<��a<�a<I�a<��a<�a<��a<I�a</�a<+�a<'�a<Q�a<O�a<U�a<d�a<��a<��a<#�a<p�a<��a<��a<��a<��a<�a<r�a<��a<��a<��a<_�a<��a<g�a< �a<o�a<+�a<��a<�a<5�a<F�a<$�a<�a<��a<9�a<ؙa<S�a<��a<��a<u�a<p�a<��a<�a<H�a<Ǚa<V�a<�a<v�a<�a<��a<ǜa<�a<�a<לa<��a<'�a<��a<t�a<�a<��a<k�a<U�a<J�a<h�a<��a<��a<1�a<r�a<ԛa<��a< �a<��a<��a<X�a<Қa<�a<��a<̘a<�a<��a< �a<��a<Y�a<H�a<d�a<��a<ߖa<G�a<��a<֗a<E�a<U�a<]�a<G�a<�a<��a<�a<G�a<��a<&�a<h�a<�a<z�a<3�a<�a<Ӓa<Вa<�a<ɒa<�a<�a<��a<W�a<�a<A�a<��a<��a<��a<��a<y�a<��a<��a<��a<��a<f�a<�a<��a<��a<o�a<}�a<d�a<U�a<T�a<�a<��a< �a<Q�a<��a<��a<��a<ҁa<΀a<�a<1a<�~a<~a<�}a<^}a<T}a<?}a<}a<"}a<�|a<�|a<f|a<�{a<?{a<�za<�ya<�xa<xa<wa<Lva<�ua< ua<�ta<ita<fta<�ta<�ta<ua<qua<�ua<va<gva<qva<�va<Zva<&va<�ua<Tua<�ta<�ta<ta<�sa<�sa<�sa<�sa<�sa<>ta<�ta</ua<�ua<�  �  �va<�va<wa<"wa</wa<wa<�va<|va<�ua<�ua<Dua<ua<�ta<�ta<Iua<�ua<\va<wa<xa<ya<za<1{a<|a<}a<�}a<e~a<�~a<Da<�a<�a<1�a<1�a<��a<�a<G�a<�a<l�a<t�a< �a<'�a<�a<��a<͇a<��a<;�a<��a<:�a<D�a<k�a<��a<f�a<��a<s�a<��a<܊a<C�a<݋a<��a<��a<��a<a<Đa<�a<�a<�a<�a<��a<C�a<��a<�a<�a<�a<6�a<�a<N�a<(�a<r�a<��a<�a<��a<ؘa<��a<�a<��a<ɚa<�a<>�a<2�a<.�a<��a<f�a<ؙa<H�a<ݘa<O�a<�a<a<ʗa<ԗa<.�a<��a<-�a<�a<z�a<R�a<Ûa<]�a<Ӝa<�a<�a<��a<�a<��a<[�a<�a<|�a<q�a<�a<�a<�a<-�a</�a<r�a<қa<�a<$�a<�a<-�a<�a<��a<6�a<z�a<�a<�a<O�a<��a<ږa<V�a<ڕa<��a<��a<��a<�a<Z�a<��a<+�a<��a<�a<Q�a<N�a<E�a<�a<��a<e�a<a<a�a<��a<'�a<��a<-�a<�a<��a<��a<I�a<{�a<_�a<M�a<&�a<Ւa<��a<ܑa<Y�a<K�a<V�a<b�a<�a<�a<؊a<��a<��a<7�a<��a<C�a<�a<�a<
�a<��a<%�a<�a<�a<��a<|�a< �a<}�a<̄a<�a<"�a<b�a<B�a<ŀa<�a<Ma<�~a<_~a<0~a<�}a<�}a<�}a<z}a<#}a<�|a<o|a<�{a<I{a<Hza<�ya<yxa<twa<�va<�ua<�ta<Lta<�sa<�sa<�sa<�sa<ta<�ta<�ta<�ua<�ua<0va<}va<tva<�va<Hva<va<�ua<ua<ua<�ta<�ta<>ta<Zta<Nta<�ta<�ta<Aua<�ua<va<�  �  �va<#wa<Owa<2wa<wa<�va<wva<va<�ua<5ua<�ta<�ta<kta<qta<�ta<(ua<�ua<�va<�wa<�xa<�ya<�za<�{a<�|a<�}a<�~a<3a<�a<�a<I�a<��a<��a<�a<^�a<ρa<n�a<��a<�a<��a<��a<p�a<L�a<�a<ވa<b�a<��a<�a<�a<(�a<1�a<�a<
�a<��a<#�a<d�a<��a<J�a<!�a<�a<�a<;�a<d�a<��a<ɒa<֓a<�a<��a<g�a<��a<*�a<j�a<��a<��a<��a<×a<��a<��a<2�a<��a<�a<_�a<��a<n�a<Қa< �a<j�a<[�a<1�a<�a<{�a<�a<��a<�a<U�a<Ηa<{�a<F�a<)�a<S�a<��a<�a<��a<s�a<(�a<�a<��a<+�a<��a<��a<I�a<V�a<,�a<��a<��a<b�a<�a<�a<��a<��a<y�a<��a<Ûa<�a<#�a<W�a<i�a<y�a<a�a<��a<��a<�a<J�a<��a<��a<�a<�a<W�a<͕a<[�a<�a<�a<0�a<l�a<וa<T�a<ݖa<W�a<��a<&�a<N�a<_�a<_�a<�a<��a<@�a<��a<�a<��a<�a<��a<t�a< �a<!�a<��a<�a<˓a<��a<h�a</�a<��a<�a<5�a< �a<�a<��a<��a<��a<]�a<c�a<~�a<��a<�a<ˆa<��a<k�a<��a<��a<��a<Ɇa<Ɔa<ӆa<��a<C�a<؅a<�a<e�a<��a<΂a<ԁa<:�a<Y�a<�a<Ha<�~a<�~a<L~a<;~a<~a<�}a<{}a<-}a<�|a<�{a<{a<za<*ya<$xa<wa<va< ua<gta<�sa<Xsa<*sa<2sa<Rsa<�sa<ta<�ta<&ua<�ua<�ua<eva<�va<�va<�va<fva<)va<�ua<�ua<:ua<ua<�ta<�ta<�ta<,ua<iua<�ua<!va<�va<�  �  �va<?wa<@wa<Kwa<wa<�va<�va<�ua<cua<�ta<`ta<ta<�sa<�sa< ta<�ta<Iua<=va<!wa<Gxa<wya<�za<�{a<�|a<�}a<�~a<#a<�a<�a<��a<рa<5�a<m�a<�a<b�a<ނa<��a<3�a<�a<�a<��a<��a<3�a<؈a<S�a<̉a<�a<+�a<�a<Չa<Ӊa<��a<��a<��a<Ήa<D�a<Њa<��a<��a<��a<a<,�a<U�a<��a<�a<��a<��a<Y�a<�a<R�a<��a<ŗa<��a<�a<�a<U�a<o�a<��a<�a<^�a<�a<D�a<��a<��a<H�a<X�a<Y�a<<�a<ښa<��a<יa<8�a<��a<�a<|�a<��a<��a<��a<ۖa<�a<��a<P�a<��a<�a<��a<��a<(�a<��a<�a<<�a<k�a<O�a<D�a<��a<Ӝa<}�a<F�a<5�a<�a<�a<�a<�a<d�a<r�a<��a<��a<��a<S�a<�a<��a<��a<W�a<C�a<x�a<w�a<��a<��a<A�a<��a<��a<��a<��a<�a<j�a<��a<��a<�a<Ǘa< �a<O�a<g�a<O�a<5�a<ԗa<��a<�a<��a<�a<��a<H�a<�a<��a<l�a<_�a<A�a<�a<�a<��a<)�a<��a<��a<�a<2�a<�a<��a<�a<�a<�a<�a<�a<7�a<��a<3�a<�a<�a<
�a<Y�a<i�a<��a<ކa<��a<��a<6�a<Ʌa<=�a<��a<Ճa< �a<Z�a<~�a<��a<K�a<�a<ra<�~a<�~a<�~a<E~a<�}a<�}a<}a<�|a<�{a<�za<*za<�xa<�wa<�va<�ua<�ta<�sa<Ksa<�ra<�ra<�ra<�ra<@sa<�sa<Yta<�ta<�ua<�ua<Hva<�va<�va<�va<�va<qva<#va<�ua<�ua<pua<mua<Qua<|ua<�ua<�ua<3va<pva<�va<�  �  4wa<cwa<fwa<Zwa< wa<�va<-va<�ua<0ua<�ta<)ta<�sa<�sa<�sa<�sa<nta<ua<�ua<�va<xa<Mya<sza<�{a<�|a<�}a<�~a<Ka<�a<Y�a<��a<�a<f�a<��a<!�a<��a<�a<˃a<|�a<N�a<�a<�a<Ça<q�a<�a<z�a<щa<։a<�a<Ӊa<��a<��a<n�a<f�a<a�a<��a<�a<��a<\�a<C�a<r�a<��a<��a<8�a<o�a<��a<��a<��a<|�a<�a<��a<ݗa<�a<�a<B�a<P�a<��a<��a<�a<N�a<��a<�a<u�a<�a<8�a<v�a<|�a<p�a<<�a<��a<?�a<��a<�a<f�a<��a<8�a<��a<��a<|�a<��a<�a<p�a<�a<֘a<��a<��a<B�a<�a<��a<"�a<g�a<��a<��a<s�a<:�a<�a<��a<��a<`�a<;�a<A�a<N�a<\�a<��a<��a<Μa<ɜa<��a<y�a<$�a<}�a<a<��a<(�a<E�a<L�a<n�a<��a<�a<��a<c�a<X�a<s�a<єa<7�a<ϕa<j�a<�a<q�a<ۗa<G�a<y�a<w�a<`�a<�a<��a<<�a<˖a<A�a<�a<w�a<�a<�a<��a<��a<j�a<K�a< �a<ʓa<W�a<��a<�a<��a<�a<��a<��a<H�a<��a<ˉa<��a<��a<�a<p�a<�a<ʅa<مa<�a<!�a<L�a<o�a<��a<��a<��a<X�a<�a<v�a<ׄa<�a<D�a<��a<ǁa<+�a<��a<�a<�a<=a<a<�~a<~a</~a<�}a<?}a<�|a<�{a<�za<�ya<�xa<�wa<�va<uua<�ta<�sa<sa<�ra<|ra<mra<�ra<sa<�sa<&ta<�ta<Dua<�ua<8va<�va<�va<�va<�va<�va<^va<"va<�ua<�ua<�ua<�ua<�ua<�ua<va<cva<�va< wa<�  �  va<va<va<�ua<�ua<(ua<>ta<�sa<�ra<�qa<qa<�pa<7pa<pa<Npa<�pa<�qa<�ra<�sa<`ua<�va<dxa<�ya<X{a<H|a<A}a<~a<�~a<Ia<�a<�a<5�a<��a<�a<P�a<�a<��a<h�a<9�a<�a<��a<��a<��a<��a<m�a<��a<ֈa<��a</�a<͇a<B�a<�a<��a<��a<��a<ӆa<i�a<Z�a<k�a<��a<J�a<��a<j�a< �a<}�a<�a<a<��a<b�a<�a<0�a<v�a<��a<��a<��a<��a<��a<�a<y�a<�a<]�a<ʙa<K�a<��a<��a<ǚa<��a<4�a<�a<��a<�a<�a<&�a<F�a<m�a<ܓa<��a<F�a<r�a<�a<��a<o�a<��a<��a<ǘa<̙a<�a<��a<�a<��a<��a<�a<��a<|�a<,�a<��a<��a<l�a<b�a<P�a<x�a<��a<��a<�a<�a<!�a<�a<��a<�a<��a<Ιa<��a<r�a<�a<�a<Гa<Ւa<�a<|�a<.�a<B�a<��a<��a<��a<��a<O�a<Q�a<�a<��a<@�a<��a<��a<��a<h�a<�a<{�a<��a<��a<�a<��a<J�a<�a<��a<֓a<��a<��a<c�a<#�a<��a<�a<��a<&�a<a<?�a<��a<�a<��a<
�a<Åa<��a<��a<%�a<�a<тa<��a<c�a<��a<C�a<��a<%�a<��a<N�a<@�a<�a<w�a<ǃa<�a<D�a<s�a<��a<�a<Ia<�~a<\~a<~a<�}a<�}a<l}a<}a<�|a<|a<O{a<^za<�ya<xa<�va<6ua<�sa<�ra<Bqa<Kpa<�oa<�na<�na<�na<Ooa<�oa<�pa<oqa<{ra<Ksa<:ta<�ta<ua<yua<�ua<�ua<`ua<ua<�ta<�ta<\ta<ta<(ta</ta<vta<�ta<ua<gua<�ua<�  �  �ua<-va< va<�ua<�ua<�ta<Gta<�sa<�ra<�qa<5qa<�pa<Npa<^pa<�pa<qa<�qa<�ra<ta<�ua<�va<xa<�ya<{a<O|a<[}a<$~a<�~a<5a<�a<�a<�a<P�a<a<%�a<��a<y�a<)�a<�a<�a<܅a<��a<}�a<�a<��a<��a<��a<p�a<B�a<�a<�a<�a<ǆa<��a<��a<�a<��a<��a<��a<�a<W�a<��a<��a<�a<d�a<��a<�a<ѕa<q�a<�a<(�a<Q�a<Z�a<f�a<i�a<��a<��a<�a<_�a<��a<;�a<��a<+�a<��a<Κa<Кa<��a<B�a<��a<�a<4�a<>�a<N�a<[�a<��a<�a<��a<��a<��a<
�a<Ɣa<��a<��a<a<�a<ڙa<��a<��a<6�a<��a<՜a<Ҝa<��a<b�a<�a<Ûa<��a<W�a<&�a<2�a<I�a<e�a<��a<͛a<��a<�a<�a<��a<7�a<|�a<��a<��a<��a<Q�a<�a<�a<�a<%�a<��a<p�a<r�a<��a<+�a<͒a<��a<��a<l�a<�a<��a<G�a<��a<��a<��a<T�a<�a<c�a<�a<G�a<�a<j�a<�a<��a<��a<��a<��a<��a<W�a<�a<��a<�a<�a<�a<��a<R�a<܋a<B�a<��a<6�a<�a<τa<�a<h�a<�a<��a<*�a<p�a<�a<i�a<Єa<�a<M�a<m�a<V�a<��a<z�a<��a<��a<�a<H�a<q�a<�a<a<�~a<B~a<�}a<�}a<v}a<K}a<�|a<�|a<|a<f{a<lza<Aya<xa<�va<dua<�sa<�ra<tqa<^pa<�oa<>oa<oa<oa<~oa<pa<�pa<�qa<�ra<Zsa<ta<�ta<8ua<�ua<�ua<�ua<Mua< ua<�ta<`ta<&ta<	ta<�sa<ta<Gta<�ta<�ta<Hua<�ua<�  �  �ua<�ua<�ua<�ua<�ua<ua<�ta<�sa<�ra<0ra<�qa<qa<�pa<�pa<�pa<dqa<ra<Hsa<Yta<�ua<$wa<�xa<za<5{a<o|a<A}a<�}a<�~a<�~a<Ya<�a<�a<�a<m�a<݀a<c�a<'�a<ɂa<΃a<��a<��a<��a<<�a<߇a<K�a<��a<Èa<��a<��a<�a<��a<G�a< �a<�a<�a<W�a<�a<׈a<�a<I�a<��a<5�a<��a<I�a<��a<Փa<�a<��a<?�a<��a<��a<	�a<�a<.�a<�a<I�a<`�a<��a<�a<]�a<�a<i�a<�a<G�a<��a<��a<��a<a�a<řa<D�a<[�a<f�a<��a<��a<�a<M�a<��a<Ɠa<�a<`�a<*�a<�a<ۖa<��a<��a<%�a<�a<��a<1�a<b�a<��a<��a<t�a<�a<ٛa<��a<#�a<�a<ٚa<�a<�a<"�a<h�a<��a<ɛa<ța<ța<r�a<+�a<��a<��a<�a<��a<��a<X�a<C�a<j�a<��a<�a<��a<��a<��a<��a<�a<�a<��a<��a<i�a<ږa<h�a<��a<y�a<r�a<�a<��a<�a<��a<��a<��a<!�a<Ɠa<��a<X�a<k�a<S�a<<�a<&�a<ےa<q�a<ˑa<�a<�a<�a<��a<�a<��a<�a<��a<H�a<!�a<?�a<��a<g�a<W�a<��a<��a<-�a<��a<�a<Z�a<m�a<�a<%�a<Ąa<;�a<��a<��a<ہa<�a<�a<~a<�~a<L~a<�}a<�}a<|}a<2}a<	}a<�|a<o|a<�{a<E{a<�za<gya<bxa<�va<�ua<?ta<�ra<�qa<�pa<pa<voa<[oa<foa<�oa<^pa<qa<�qa<�ra<�sa<>ta<�ta<3ua<Fua<dua<Aua<ua<�ta<sta< ta<�sa<�sa<�sa<�sa<�sa<Eta<�ta<ua<zua<�  �  ~ua<�ua<�ua<�ua<�ua<,ua<�ta<�sa<Rsa<�ra<ra<�qa<Lqa<Nqa<�qa<	ra<�ra<�sa<�ta<Lva<�wa<�xa<za<W{a<S|a<2}a<�}a<X~a<�~a<�~a<a<Ea<�a<�a<*�a<ˀa<V�a<S�a<0�a</�a<�a<�a< �a<·a<S�a<��a<ވa<��a<��a<d�a<#�a<�a<��a<��a<��a<�a<��a<y�a<q�a<��a<9�a<��a<�a<w�a<��a<��a<єa<��a<6�a<n�a<��a<��a<��a<��a<��a<|�a<Ėa<��a<O�a<�a<b�a<�a<y�a<��a<I�a<��a<��a<C�a<�a<7�a<��a<Ηa<�a<3�a<u�a<�a<��a<��a<��a<�a<��a<h�a<x�a<W�a<G�a</�a<��a<��a<�a<|�a<y�a<V�a<�a<��a<N�a<�a<��a<;�a<J�a<#�a<X�a<��a<֚a<�a<Z�a<��a<��a<��a<�a<��a<ҙa<�a<�a<�a<�a<Ŕa<ޓa<$�a<��a<l�a<f�a<��a<�a<��a<p�a<�a<Ǖa<a�a<��a<M�a<{�a<��a<4�a<Ԗa<E�a<��a<�a<��a<�a<n�a<.�a<Ғa<�a<͒a<Ւa<ƒa<��a<��a<_�a<ӑa<�a<.�a<�a<��a<O�a<�a<��a<�a<Ɇa<Åa<�a<c�a<
�a<؃a<�a<S�a<��a<�a<5�a<X�a<��a<]�a<�a<��a<��a<+�a<@�a<^�a<m�a<�a<�~a<-~a<�}a<2}a<}a<�|a<�|a<�|a<{|a<*|a<�{a<7{a<mza<�ya<Uxa<2wa<�ua<�ta<tsa<Jra<Sqa<�pa<<pa<pa<pa<Zpa<�pa<�qa<Dra<�ra<�sa<Ota<�ta<ua<_ua<Cua<ua<�ta<Cta<�sa<�sa<=sa<�ra<sa<sa<Vsa<�sa<#ta<�ta<ua<�  �  (ua<Tua<�ua<�ua<�ua<wua<�ta<�ta<�sa<6sa<�ra<Nra<
ra<�qa<Vra<�ra<zsa<eta<�ua<�va<�wa<uya<iza<�{a<k|a<}a<�}a<�}a<^~a<f~a<�~a<�~a<�~a<a<la<�a<��a<��a<Z�a<��a<��a<��a<��a<]�a<0�a<��a<�a<�a<�a<�a<��a<x�a<A�a<L�a<c�a<͈a<i�a<$�a<;�a<a�a<ȍa<��a<��a<�a<��a<#�a<Ԕa<��a<ҕa<�a<8�a<�a< �a<��a<��a<ŕa<�a<B�a<��a<3�a<��a<�a<��a<��a<�a<S�a<l�a<P�a<&�a<��a<!�a<>�a<m�a<іa<!�a<��a<E�a<P�a<]�a<a<b�a<�a<��a<��a<�a<��a<H�a<ӛa<�a<F�a<	�a<��a<��a<8�a<��a<�a<�a<�a<��a<e�a<��a<șa<+�a<��a<ޚa<=�a<*�a<M�a<�a<��a<�a<D�a<��a<L�a<_�a<l�a<��a<�a<Y�a<6�a<�a<P�a<��a<C�a<Ԕa<��a<b�a<��a<?�a<d�a<e�a<G�a<ϖa<|�a<a<9�a<L�a<��a<4�a<��a<}�a<�a<B�a<��a<O�a<U�a<[�a<C�a<�a<��a<�a<Q�a<3�a<�a<،a<G�a<�a<��a<��a<y�a<��a<%�a<��a<��a<��a<�a<��a<f�a<��a<��a<��a<`�a<
�a<W�a<��a<ςa<Ɂa<�a<�a<�~a<�}a<x}a<�|a<�|a<]|a<|a<H|a<|a<&|a<�{a<�{a<#{a<zza<�ya<�xa<�wa<cva<ua<ta<�ra<ra<Rqa< qa<�pa<�pa<qa<�qa<"ra<�ra<�sa<ta<�ta<�ta<ua<)ua<�ta<�ta<8ta<�sa<Nsa<�ra<�ra<2ra<bra<Era<�ra<�ra<xsa<"ta<�ta<�  �  �ta<)ua<�ua<�ua<�ua<�ua<Qua<�ta<kta<�sa<ysa< sa<�ra<�ra<9sa<�sa<hta<>ua<Iva<xwa<�xa<�ya<�za<�{a<||a<}a<x}a<�}a<�}a<�}a<�}a<�}a<�}a<0~a<s~a<a<�a<��a<��a<�a<��a<,�a<D�a<1�a<�a<��a<��a<X�a<X�a<J�a<L�a< �a<�a<)�a<S�a<��a<R�a<�a<$�a<9�a<s�a<̏a<��a<)�a<Y�a<�a<�a<l�a<��a<��a<��a<]�a<]�a<�a<�a<�a<�a<A�a<ĕa<X�a<��a<��a<J�a<�a<��a<�a<^�a<g�a<&�a<�a<Z�a<Řa<:�a<��a<��a<��a<D�a<2�a<X�a<��a<3�a<�a<��a<v�a<*�a<�a<~�a<қa<�a<�a<��a<��a<�a<d�a<��a<r�a<�a<��a<��a<w�a<��a<�a<u�a<ҙa<H�a<Ěa<��a<�a<�a<��a<B�a<��a<Řa<��a<�a<6�a<m�a<˔a<Z�a<�a<�a<?�a<��a<�a<��a<�a<��a<�a<H�a<u�a<]�a<�a<��a<��a<�a<k�a<��a<��a<Q�a<��a<r�a<5�a<O�a<W�a<��a<��a<ґa<�a<a<��a<�a<G�a<��a<h�a<5�a<�a<��a<��a<k�a<h�a<��a<�a<��a<��a<w�a<��a<Åa<΅a<�a<�a<��a<v�a<�a<%�a<J�a<F�a<�a< �a<�~a<~a<}a<p|a<�{a<�{a<�{a<q{a<~{a<j{a<�{a<�{a<b{a<{a<�za<�ya<ya<�wa<�va<�ua<�ta<�sa<sa<Qra<�qa<�qa<�qa<�qa<Sra<�ra<csa<�sa<jta<�ta<�ta<ua<�ta<�ta<Cta<�sa<sa<�ra<ra<�qa<Hqa<Lqa<Wqa<�qa<8ra<�ra<Nsa<�sa<�  �  ta<�ta<Dua<�ua<�ua<�ua<�ua<Iua<"ua<�ta<Gta<�sa<�sa<�sa<4ta<�ta<Dua<"va<wa<'xa<=ya<za<6{a<�{a<�|a<�|a<:}a<P}a<4}a<M}a<}a<
}a<�|a<0}a<�}a<~a<�~a<�a<ހa<�a<_�a<��a<��a<��a<��a<��a<�a<��a<��a<ԉa<�a<݉a<��a<��a<I�a<��a<L�a<�a<��a<�a<7�a<��a<��a<��a<��a<8�a<�a<�a<l�a<1�a<�a<�a<��a<D�a<�a<�a<�a<Z�a<Ȕa<X�a<(�a<�a<ٗa<y�a<6�a<ۙa<�a<n�a<R�a<R�a<��a<o�a<�a<K�a<ٗa<q�a<A�a<4�a<Z�a<��a<�a<��a<]�a</�a<��a<R�a<��a<�a<�a<ɛa<��a<�a<��a<ϙa<�a<��a< �a<��a<��a<��a<��a<"�a<��a<.�a<љa<�a<��a<՚a<�a<Ța<v�a<�a<:�a<��a<͗a<�a<K�a<��a<[�a<�a<�a<�a<m�a<Ǖa<M�a<ɖa<��a<��a<t�a<}�a<(�a<Жa<-�a<R�a<��a<��a<Ғa<��a<P�a<ِa<��a<W�a<N�a<{�a<��a<�a<A�a<L�a<��a<>�a<�a<a�a<Ϗa<ˎa<��a<Ča<w�a<f�a<@�a<^�a<��a<�a<��a<^�a<Y�a<P�a<z�a<e�a<L�a<O�a<υa<o�a<��a<�a<��a<��a<��a<Ca<&~a<}a<7|a<�{a<�za<�za<�za<�za<�za<�za<�za<{a<${a<�za<�za<�ya<oya<[xa<�wa<�va<�ua<�ta<�sa<Msa<�ra<�ra<�ra<�ra<&sa<�sa<ta<Wta<�ta<
ua<ua<ua<�ta<jta<�sa<+sa<mra<�qa<%qa<�pa<spa<Ypa<�pa<�pa<Eqa<�qa<�ra<�sa<�  �  �sa<nta<ua<�ua<�ua<va<va<�ua<�ua<Pua<ua<�ta<�ta<�ta<)ua<�ua<Iva<
wa<�wa<�xa<�ya<�za<r{a<|a<�|a<�|a<�|a<�|a<�|a<�|a<]|a<3|a<%|a<?|a<�|a<}a<�}a<�~a<�a<E�a<��a<��a<I�a<��a<��a<��a<[�a<ىa<8�a<w�a<p�a<��a<Ȋa<��a<?�a<��a<:�a< �a<��a<�a<�a<��a<(�a<�a<ݓa<��a<�a<��a<�a<˔a<{�a<2�a<��a<a�a<1�a<�a<�a<b�a<ԓa<��a<L�a<*�a<$�a<��a<Әa<��a<�a<{�a<��a<��a<X�a<��a<n�a<)�a<��a<w�a<�a<(�a<5�a<��a<�a<��a<�a<��a<L�a<��a<��a<�a<��a<��a<5�a<�a<ϙa<�a<R�a<��a<#�a<a<��a<��a<ܖa<B�a<їa<{�a<�a<��a<C�a<��a<ޚa<�a<��a<_�a<�a<&�a<y�a<ܗa<C�a<��a<3�a<
�a<�a< �a<U�a<��a<ۖa<M�a<��a<��a<×a<��a<�a<��a<Ǖa<הa<�a<�a<��a<�a<_�a<ڏa<~�a<X�a<w�a<��a<�a<W�a<��a<�a<4�a<�a<�a<��a<
�a<G�a<b�a<4�a<N�a<6�a<@�a<T�a<��a<��a<��a<^�a<-�a<+�a<�a<�a<ֆa<��a<�a<r�a<~�a<��a<V�a<�a<�a<~~a<D}a<:|a<8{a<�za<za<�ya<�ya<�ya<�ya<Eza<sza<�za<�za<�za<�za<Cza<�ya<�xa<!xa<wa<hva<�ua<�ta<*ta<�sa<�sa<�sa<�sa<�sa<Eta<�ta< ua</ua<Jua<>ua<�ta<�ta<�sa<6sa<wra<�qa<�pa<Bpa<�oa<uoa<]oa<�oa<�oa<fpa<qa<�qa<�ra<�  �  `sa<ta<�ta<�ua<�ua<Gva<>va<mva<1va<$va<�ua<�ua<�ua<�ua<>va<ova<7wa<�wa<�xa<�ya<Mza<{a<�{a<J|a<�|a<�|a<�|a<�|a<k|a<�{a<�{a<d{a<S{a<V{a<�{a<9|a<�|a<�}a<#a<��a<�a<w�a<�a<;�a<��a<��a<l�a<�a<��a<�a<&�a<|�a<b�a<ߋa<�a<��a<C�a<ۍa<�a<��a<Րa<��a<��a<k�a<�a<��a<Дa<�a<��a<��a<�a<c�a<�a<��a<@�a<�a<3�a<q�a<�a<��a<w�a<��a<a�a<��a<��a<I�a<�a<h�a<ƚa<��a<��a<��a<>�a<�a<]�a<h�a<�a<5�a<+�a<��a<Ιa<5�a<�a<B�a<ʛa<�a<1�a<�a<�a<��a<Ӛa<M�a<6�a<X�a<��a<ʖa<5�a<��a<��a<��a<�a<m�a<
�a<��a<r�a<u�a<�a<��a<ؚa<�a<�a<��a<^�a<��a<M�a<��a<��a<��a<$�a<�a<͖a<�a<��a<g�a<��a<ڗa<�a<�a<�a<��a<�a<Q�a<t�a<��a<6�a<B�a<-�a<J�a<v�a<�a<��a<[�a<��a<��a<6�a<��a<�a<��a<̐a<�a<�a<��a<E�a<��a<�a<�a<�a<ыa<!�a</�a<��a<��a<l�a<J�a<ɇa<�a<��a<��a<)�a<��a<3�a<\�a<��a<9�a<�a<��a<a<�}a<j|a<I{a<Aza<�ya<ya<�xa<�xa<�xa<Iya<�ya<za<fza<�za<�za<�za<gza<�ya<\ya<�xa<�wa<.wa<1va<�ua<ua<�ta<�ta<�ta<�ta<�ta<ua</ua<~ua<hua<�ua<Cua<�ta<rta<�sa<sa<�qa<�pa<*pa<hoa<�na<rna<yna<}na<�na<�oa<Wpa<:qa<$ra<�  �  �ra<�sa<�ta<uua<va<�va<�va<�va<�va<�va<�va<yva<rva<�va<�va<)wa<�wa<�xa<Aya<�ya<�za<v{a<	|a<z|a<�|a<�|a<s|a</|a<�{a<s{a<({a<�za<�za<�za<�za<w{a<@|a<0}a<{~a<�a<��a<�a<��a<�a<f�a<|�a<�a<b�a<֊a<X�a<��a<�a<2�a<��a<ʌa<^�a<��a<��a<��a<\�a<J�a<*�a<�a<��a<l�a<��a<̔a<Ӕa<j�a<�a<��a<�a<z�a<ݑa<y�a<d�a<q�a<��a<0�a<�a<ɓa<��a<��a<�a<�a<�a<�a<n�a<�a<!�a<�a<�a<��a<z�a<2�a<�a<��a<�a<�a<.�a<��a<�a<U�a<ěa<#�a<T�a<u�a<1�a<ћa<F�a<}�a<��a<Ęa<�a<�a<�a<w�a<�a<�a<�a<1�a<��a<f�a<Q�a<�a<טa<��a<<�a<��a<��a<-�a<��a<��a<=�a<��a<@�a<ǘa<L�a<�a<̗a<��a<��a<͗a<��a<�a<I�a<e�a<V�a< �a<��a<��a<	�a<�a<�a<ϒa<��a<~�a<��a<��a<,�a<ڍa<��a<��a<�a<��a<,�a<��a<&�a<}�a<�a<�a<ΐa<��a<�a<B�a<d�a<��a<��a<ًa<ߊa<F�a<��a< �a<��a<��a<d�a<"�a<�a<}�a<�a<I�a<X�a<Y�a<��a<��a<)�a<�~a<>}a<�{a<�za<�ya<�xa<Txa<xa<xa<?xa<�xa<ya<�ya<�ya<Lza<�za<�za<�za<>za<�ya<ya<^xa<�wa<wa<rva<�ua<�ua<Aua<2ua<Nua<aua<�ua<�ua<�ua<�ua<�ua<Xua<�ta<*ta<Hsa<era<mqa<�pa<�oa<�na<na<�ma<�ma<�ma<1na<�na<�oa<�pa<�qa<�  �  rra<�sa<�ta<}ua<va<qva<�va<�va<wa<wa<wa< wa<wa<;wa<{wa<�wa<`xa<ya<�ya<nza<({a<�{a<'|a<f|a<�|a<�|a<g|a<!|a<{a<{a<�za<>za<za<�ya<<za<�za<�{a<�|a<~a<Wa<
�a<��a<S�a<��a<>�a<��a<��a<]�a<�a<��a<�a<g�a<،a<�a<��a<�a<��a<Z�a<�a<�a<ȑa<��a<g�a<�a<r�a<��a<�a<��a<p�a<�a<)�a<��a<Ցa<r�a<��a<��a<��a< �a<��a<g�a<S�a<S�a<��a<��a< �a<��a<ՙa<��a<�a<8�a<S�a<V�a<&�a<��a<Кa<��a<��a<z�a<��a<Ԛa<�a<��a<͛a<5�a<`�a<��a<`�a<@�a<�a<(�a<��a<i�a<c�a<e�a<a�a<��a<ٔa<s�a< �a<R�a<��a<C�a<ޕa<��a<��a<��a<��a< �a<Śa<�a<�a</�a<�a<��a<,�a<ՙa<N�a<�a<��a<]�a<V�a<8�a<g�a<��a<��a<��a<��a<s�a<�a<��a<�a<��a<��a<��a<s�a<�a<�a<�a<�a<��a<�a<�a<-�a<��a<��a<��a<A�a<�a<��a<��a<�a<ڐa<��a<-�a<��a<ӎa<�a<F�a<E�a<��a<�a<S�a<�a<g�a<A�a<�a<��a<@�a<ća<�a<Q�a<y�a<3�a<��a<o�a<�a<A~a<�|a<U{a<�ya<�xa<xa<�wa<owa<�wa<�wa<xa<�xa<1ya<�ya<Eza<�za<�za<�za<Uza<�ya<zya<�xa<9xa<�wa<�va<�va<)va<�ua<�ua<�ua<�ua<�ua<"va<va<va<�ua<gua<�ta<ta<Msa< ra<qa<pa<�na<Jna<�ma<(ma<�la<4ma<�ma<gna<,oa<8pa<Vqa<�  �  ara<gsa<dta<^ua<%va<�va<wa<=wa<Uwa<Jwa<Kwa<Ewa<ewa<�wa<�wa<Hxa<�xa<Xya<�ya<�za<Y{a<�{a<_|a<�|a<�|a<�|a<*|a<�{a<m{a<�za<Qza<�ya<�ya<�ya<�ya<xza<G{a<@|a<�}a<a<ˀa<v�a<'�a<��a<�a<�a<��a<��a<_�a<ދa<U�a<��a<�a<S�a<ߍa<H�a<ގa<��a<V�a<:�a<�a<�a<��a<E�a<��a<�a<הa<��a<!�a<��a<�a<Y�a<��a<�a<��a<n�a<t�a<��a<:�a<�a<��a<�a<^�a<��a<��a<��a<��a<��a<�a<l�a<��a<��a<m�a<4�a<	�a<�a<�a<Ěa<�a<*�a<`�a<Ûa<�a<m�a<��a<ǜa<��a<U�a<Ǜa<��a<.�a<S�a<9�a<&�a<�a<C�a<y�a<$�a<�a<�a<3�a<ڔa<��a<�a<w�a<u�a<<�a<��a<��a<�a<V�a<j�a</�a<�a<s�a<	�a<��a<?�a<�a<��a<��a<��a<��a<��a<ۘa<�a<�a<��a<K�a<��a<іa<��a<��a<��a<9�a<�a<��a<��a<��a<:�a<یa<Ìa<όa<C�a<��a<s�a<�a<ŏa<6�a<��a<�a< �a<Ȑa<n�a<ȏa<�a<F�a<|�a<��a<�a<0�a<��a<;�a<��a<x�a<&�a<ۈa<s�a<�a<N�a<~�a<c�a<�a<��a<;�a<�a<~a<]|a<�za<�ya<�xa<�wa<cwa<wa<0wa<qwa<�wa<~xa<ya<�ya< za<mza<�za<�za<�za<3za<�ya<ya<sxa<�wa<Owa<�va<sva<Bva<.va<va<1va<?va<Zva<Tva<Fva<�ua<|ua<�ta<�sa<�ra<	ra<�pa<�oa<�na<�ma<ma<�la<�la<�la<2ma<�ma<�na<�oa<)qa<�  �  Fra<bsa<�ta<gua<va<�va<wa<Uwa<mwa<hwa<jwa<�wa<�wa<�wa<xa<Yxa<�xa<�ya<za<�za<j{a<	|a<G|a<�|a<�|a<�|a<W|a<�{a<O{a<�za<Eza<�ya<�ya<�ya<�ya<0za<{a<+|a<t}a<a<��a<L�a<�a<��a<c�a<l�a<��a<��a<O�a<�a<x�a<Ɍa<2�a<��a<��a<{�a<�a<��a<��a<a�a</�a<�a<��a<=�a<��a<єa<��a<̔a<4�a<��a<�a<!�a<��a<��a<s�a<D�a</�a<y�a<�a<ߑa<Ғa<�a<!�a<��a<��a<ۘa<�a<_�a<�a<U�a<��a<��a<��a<Z�a<<�a<�a<�a<��a<�a<N�a<��a<�a<-�a<��a<��a<��a<��a<;�a<śa<H�a<.�a<9�a<��a<�a<��a<�a<e�a<�a<��a<Ǔa<�a<��a<p�a<h�a<9�a<Z�a<7�a<;�a<��a<��a<J�a<R�a<G�a<��a<��a<(�a<ҙa<j�a<�a<�a<��a<Ϙa<ژa<ؘa<��a<��a<��a<��a<:�a<��a<�a<�a<��a<n�a<��a<ڐa<��a<�a<��a<�a<��a<��a<��a<�a<��a<E�a<�a<��a<A�a<�a<Րa<�a<��a<^�a<؏a<;�a<c�a<��a<܌a<�a<c�a<ъa<N�a<�a<��a<H�a<��a<}�a<��a<A�a<i�a<G�a<R�a<��a<*�a<|a<�}a<N|a<�za<|ya<zxa<�wa<wa<�va<	wa<Gwa<�wa<Axa<�xa<�ya<$za<�za<�za<�za<rza<Aza<�ya<:ya<�xa<xa<�wa<�va<�va<iva<Sva<[va<Ova<Xva<tva<lva<*va<�ua<bua<�ta<,ta<�ra<�qa<�pa<�oa<�na<�ma<ma<�la<rla<�la<ma<�ma<�na<�oa<�pa<�  �  ara<gsa<dta<^ua<%va<�va<wa<=wa<Uwa<Jwa<Kwa<Ewa<ewa<�wa<�wa<Hxa<�xa<Xya<�ya<�za<Y{a<�{a<_|a<�|a<�|a<�|a<*|a<�{a<m{a<�za<Qza<�ya<�ya<�ya<�ya<xza<G{a<@|a<�}a<a<ˀa<v�a<'�a<��a<�a<�a<��a<��a<_�a<ދa<U�a<��a<�a<S�a<ߍa<H�a<ގa<��a<V�a<:�a<�a<�a<��a<E�a<��a<�a<הa<��a<!�a<��a<�a<Y�a<��a<�a<��a<n�a<t�a<��a<:�a<�a<��a<�a<^�a<��a<��a<��a<��a<��a<�a<l�a<��a<��a<m�a<4�a<	�a<�a<�a<Ěa<�a<*�a<`�a<Ûa<�a<m�a<��a<ǜa<��a<U�a<Ǜa<��a<.�a<S�a<9�a<&�a<�a<C�a<y�a<$�a<�a<�a<3�a<ڔa<��a<�a<w�a<u�a<<�a<��a<��a<�a<V�a<j�a</�a<�a<s�a<	�a<��a<?�a<�a<��a<��a<��a<��a<��a<ۘa<�a<�a<��a<K�a<��a<іa<��a<��a<��a<9�a<�a<��a<��a<��a<:�a<یa<Ìa<όa<C�a<��a<s�a<�a<ŏa<6�a<��a<�a< �a<Ȑa<n�a<ȏa<�a<F�a<|�a<��a<�a<0�a<��a<;�a<��a<x�a<&�a<ۈa<s�a<�a<N�a<~�a<c�a<�a<��a<;�a<�a<~a<]|a<�za<�ya<�xa<�wa<cwa<wa<0wa<qwa<�wa<~xa<ya<�ya< za<mza<�za<�za<�za<3za<�ya<ya<sxa<�wa<Owa<�va<sva<Bva<.va<va<1va<?va<Zva<Tva<Fva<�ua<|ua<�ta<�sa<�ra<	ra<�pa<�oa<�na<�ma<ma<�la<�la<�la<2ma<�ma<�na<�oa<)qa<�  �  rra<�sa<�ta<}ua<va<qva<�va<�va<wa<wa<wa< wa<wa<;wa<{wa<�wa<`xa<ya<�ya<nza<({a<�{a<'|a<f|a<�|a<�|a<g|a<!|a<{a<{a<�za<>za<za<�ya<<za<�za<�{a<�|a<~a<Wa<
�a<��a<S�a<��a<>�a<��a<��a<]�a<�a<��a<�a<g�a<،a<�a<��a<�a<��a<Z�a<�a<�a<ȑa<��a<g�a<�a<r�a<��a<�a<��a<p�a<�a<)�a<��a<Ցa<r�a<��a<��a<��a< �a<��a<g�a<S�a<S�a<��a<��a< �a<��a<ՙa<��a<�a<8�a<S�a<V�a<&�a<��a<Кa<��a<��a<z�a<��a<Ԛa<�a<��a<͛a<5�a<`�a<��a<`�a<@�a<�a<(�a<��a<i�a<c�a<e�a<a�a<��a<ٔa<s�a< �a<R�a<��a<C�a<ޕa<��a<��a<��a<��a< �a<Śa<�a<�a</�a<�a<��a<,�a<ՙa<N�a<�a<��a<]�a<V�a<8�a<g�a<��a<��a<��a<��a<s�a<�a<��a<�a<��a<��a<��a<s�a<�a<�a<�a<�a<��a<�a<�a<-�a<��a<��a<��a<A�a<�a<��a<��a<�a<ڐa<��a<-�a<��a<ӎa<�a<F�a<E�a<��a<�a<S�a<�a<g�a<A�a<�a<��a<@�a<ća<�a<Q�a<y�a<3�a<��a<o�a<�a<A~a<�|a<U{a<�ya<�xa<xa<�wa<owa<�wa<�wa<xa<�xa<1ya<�ya<Eza<�za<�za<�za<Uza<�ya<zya<�xa<9xa<�wa<�va<�va<)va<�ua<�ua<�ua<�ua<�ua<"va<va<va<�ua<gua<�ta<ta<Msa< ra<qa<pa<�na<Jna<�ma<(ma<�la<4ma<�ma<gna<,oa<8pa<Vqa<�  �  �ra<�sa<�ta<uua<va<�va<�va<�va<�va<�va<�va<yva<rva<�va<�va<)wa<�wa<�xa<Aya<�ya<�za<v{a<	|a<z|a<�|a<�|a<s|a</|a<�{a<s{a<({a<�za<�za<�za<�za<w{a<@|a<0}a<{~a<�a<��a<�a<��a<�a<f�a<|�a<�a<b�a<֊a<X�a<��a<�a<2�a<��a<ʌa<^�a<��a<��a<��a<\�a<J�a<*�a<�a<��a<l�a<��a<̔a<Ӕa<j�a<�a<��a<�a<z�a<ݑa<y�a<d�a<q�a<��a<0�a<�a<ɓa<��a<��a<�a<�a<�a<�a<n�a<�a<!�a<�a<�a<��a<z�a<2�a<�a<��a<�a<�a<.�a<��a<�a<U�a<ěa<#�a<T�a<u�a<1�a<ћa<F�a<}�a<��a<Ęa<�a<�a<�a<w�a<�a<�a<�a<1�a<��a<f�a<Q�a<�a<טa<��a<<�a<��a<��a<-�a<��a<��a<=�a<��a<@�a<ǘa<L�a<�a<̗a<��a<��a<͗a<��a<�a<I�a<e�a<V�a< �a<��a<��a<	�a<�a<�a<ϒa<��a<~�a<��a<��a<,�a<ڍa<��a<��a<�a<��a<,�a<��a<&�a<}�a<�a<�a<ΐa<��a<�a<B�a<d�a<��a<��a<ًa<ߊa<F�a<��a< �a<��a<��a<d�a<"�a<�a<}�a<�a<I�a<X�a<Y�a<��a<��a<)�a<�~a<>}a<�{a<�za<�ya<�xa<Txa<xa<xa<?xa<�xa<ya<�ya<�ya<Lza<�za<�za<�za<>za<�ya<ya<^xa<�wa<wa<rva<�ua<�ua<Aua<2ua<Nua<aua<�ua<�ua<�ua<�ua<�ua<Xua<�ta<*ta<Hsa<era<mqa<�pa<�oa<�na<na<�ma<�ma<�ma<1na<�na<�oa<�pa<�qa<�  �  `sa<ta<�ta<�ua<�ua<Gva<>va<mva<1va<$va<�ua<�ua<�ua<�ua<>va<ova<7wa<�wa<�xa<�ya<Mza<{a<�{a<J|a<�|a<�|a<�|a<�|a<k|a<�{a<�{a<d{a<S{a<V{a<�{a<9|a<�|a<�}a<#a<��a<�a<w�a<�a<;�a<��a<��a<l�a<�a<��a<�a<&�a<|�a<b�a<ߋa<�a<��a<C�a<ۍa<�a<��a<Րa<��a<��a<k�a<�a<��a<Дa<�a<��a<��a<�a<c�a<�a<��a<@�a<�a<3�a<q�a<�a<��a<w�a<��a<a�a<��a<��a<I�a<�a<h�a<ƚa<��a<��a<��a<>�a<�a<]�a<h�a<�a<5�a<+�a<��a<Ιa<5�a<�a<B�a<ʛa<�a<1�a<�a<�a<��a<Ӛa<M�a<6�a<X�a<��a<ʖa<5�a<��a<��a<��a<�a<m�a<
�a<��a<r�a<u�a<�a<��a<ؚa<�a<�a<��a<^�a<��a<M�a<��a<��a<��a<$�a<�a<͖a<�a<��a<g�a<��a<ڗa<�a<�a<�a<��a<�a<Q�a<t�a<��a<6�a<B�a<-�a<J�a<v�a<�a<��a<[�a<��a<��a<6�a<��a<�a<��a<̐a<�a<�a<��a<E�a<��a<�a<�a<�a<ыa<!�a</�a<��a<��a<l�a<J�a<ɇa<�a<��a<��a<)�a<��a<3�a<\�a<��a<9�a<�a<��a<a<�}a<j|a<I{a<Aza<�ya<ya<�xa<�xa<�xa<Iya<�ya<za<fza<�za<�za<�za<gza<�ya<\ya<�xa<�wa<.wa<1va<�ua<ua<�ta<�ta<�ta<�ta<�ta<ua</ua<~ua<hua<�ua<Cua<�ta<rta<�sa<sa<�qa<�pa<*pa<hoa<�na<rna<yna<}na<�na<�oa<Wpa<:qa<$ra<�  �  �sa<nta<ua<�ua<�ua<va<va<�ua<�ua<Pua<ua<�ta<�ta<�ta<)ua<�ua<Iva<
wa<�wa<�xa<�ya<�za<r{a<|a<�|a<�|a<�|a<�|a<�|a<�|a<]|a<3|a<%|a<?|a<�|a<}a<�}a<�~a<�a<E�a<��a<��a<I�a<��a<��a<��a<[�a<ىa<8�a<w�a<p�a<��a<Ȋa<��a<?�a<��a<:�a< �a<��a<�a<�a<��a<(�a<�a<ݓa<��a<�a<��a<�a<˔a<{�a<2�a<��a<a�a<1�a<�a<�a<b�a<ԓa<��a<L�a<*�a<$�a<��a<Әa<��a<�a<{�a<��a<��a<X�a<��a<n�a<)�a<��a<w�a<�a<(�a<5�a<��a<�a<��a<�a<��a<L�a<��a<��a<�a<��a<��a<5�a<�a<ϙa<�a<R�a<��a<#�a<a<��a<��a<ܖa<B�a<їa<{�a<�a<��a<C�a<��a<ޚa<�a<��a<_�a<�a<&�a<y�a<ܗa<C�a<��a<3�a<
�a<�a< �a<U�a<��a<ۖa<M�a<��a<��a<×a<��a<�a<��a<Ǖa<הa<�a<�a<��a<�a<_�a<ڏa<~�a<X�a<w�a<��a<�a<W�a<��a<�a<4�a<�a<�a<��a<
�a<G�a<b�a<4�a<N�a<6�a<@�a<T�a<��a<��a<��a<^�a<-�a<+�a<�a<�a<ֆa<��a<�a<r�a<~�a<��a<V�a<�a<�a<~~a<D}a<:|a<8{a<�za<za<�ya<�ya<�ya<�ya<Eza<sza<�za<�za<�za<�za<Cza<�ya<�xa<!xa<wa<hva<�ua<�ta<*ta<�sa<�sa<�sa<�sa<�sa<Eta<�ta< ua</ua<Jua<>ua<�ta<�ta<�sa<6sa<wra<�qa<�pa<Bpa<�oa<uoa<]oa<�oa<�oa<fpa<qa<�qa<�ra<�  �  ta<�ta<Dua<�ua<�ua<�ua<�ua<Iua<"ua<�ta<Gta<�sa<�sa<�sa<4ta<�ta<Dua<"va<wa<'xa<=ya<za<6{a<�{a<�|a<�|a<:}a<P}a<4}a<M}a<}a<
}a<�|a<0}a<�}a<~a<�~a<�a<ހa<�a<_�a<��a<��a<��a<��a<��a<�a<��a<��a<ԉa<�a<݉a<��a<��a<I�a<��a<L�a<�a<��a<�a<7�a<��a<��a<��a<��a<8�a<�a<�a<l�a<1�a<�a<�a<��a<D�a<�a<�a<�a<Z�a<Ȕa<X�a<(�a<�a<ٗa<y�a<6�a<ۙa<�a<n�a<R�a<R�a<��a<o�a<�a<K�a<ٗa<q�a<A�a<4�a<Z�a<��a<�a<��a<]�a</�a<��a<R�a<��a<�a<�a<ɛa<��a<�a<��a<ϙa<�a<��a< �a<��a<��a<��a<��a<"�a<��a<.�a<љa<�a<��a<՚a<�a<Ța<v�a<�a<:�a<��a<͗a<�a<K�a<��a<[�a<�a<�a<�a<m�a<Ǖa<M�a<ɖa<��a<��a<t�a<}�a<(�a<Жa<-�a<R�a<��a<��a<Ғa<��a<P�a<ِa<��a<W�a<N�a<{�a<��a<�a<A�a<L�a<��a<>�a<�a<a�a<Ϗa<ˎa<��a<Ča<w�a<f�a<@�a<^�a<��a<�a<��a<^�a<Y�a<P�a<z�a<e�a<L�a<O�a<υa<o�a<��a<�a<��a<��a<��a<Ca<&~a<}a<7|a<�{a<�za<�za<�za<�za<�za<�za<�za<{a<${a<�za<�za<�ya<oya<[xa<�wa<�va<�ua<�ta<�sa<Msa<�ra<�ra<�ra<�ra<&sa<�sa<ta<Wta<�ta<
ua<ua<ua<�ta<jta<�sa<+sa<mra<�qa<%qa<�pa<spa<Ypa<�pa<�pa<Eqa<�qa<�ra<�sa<�  �  �ta<)ua<�ua<�ua<�ua<�ua<Qua<�ta<kta<�sa<ysa< sa<�ra<�ra<9sa<�sa<hta<>ua<Iva<xwa<�xa<�ya<�za<�{a<||a<}a<x}a<�}a<�}a<�}a<�}a<�}a<�}a<0~a<s~a<a<�a<��a<��a<�a<��a<,�a<D�a<1�a<�a<��a<��a<X�a<X�a<J�a<L�a< �a<�a<)�a<S�a<��a<R�a<�a<$�a<9�a<s�a<̏a<��a<)�a<Y�a<�a<�a<l�a<��a<��a<��a<]�a<]�a<�a<�a<�a<�a<A�a<ĕa<X�a<��a<��a<J�a<�a<��a<�a<^�a<g�a<&�a<�a<Z�a<Řa<:�a<��a<��a<��a<D�a<2�a<X�a<��a<3�a<�a<��a<v�a<*�a<�a<~�a<қa<�a<�a<��a<��a<�a<d�a<��a<r�a<�a<��a<��a<w�a<��a<�a<u�a<ҙa<H�a<Ěa<��a<�a<�a<��a<B�a<��a<Řa<��a<�a<6�a<m�a<˔a<Z�a<�a<�a<?�a<��a<�a<��a<�a<��a<�a<H�a<u�a<]�a<�a<��a<��a<�a<k�a<��a<��a<Q�a<��a<r�a<5�a<O�a<W�a<��a<��a<ґa<�a<a<��a<�a<G�a<��a<h�a<5�a<�a<��a<��a<k�a<h�a<��a<�a<��a<��a<w�a<��a<Åa<΅a<�a<�a<��a<v�a<�a<%�a<J�a<F�a<�a< �a<�~a<~a<}a<p|a<�{a<�{a<�{a<q{a<~{a<j{a<�{a<�{a<b{a<{a<�za<�ya<ya<�wa<�va<�ua<�ta<�sa<sa<Qra<�qa<�qa<�qa<�qa<Sra<�ra<csa<�sa<jta<�ta<�ta<ua<�ta<�ta<Cta<�sa<sa<�ra<ra<�qa<Hqa<Lqa<Wqa<�qa<8ra<�ra<Nsa<�sa<�  �  (ua<Tua<�ua<�ua<�ua<wua<�ta<�ta<�sa<6sa<�ra<Nra<
ra<�qa<Vra<�ra<zsa<eta<�ua<�va<�wa<uya<iza<�{a<k|a<}a<�}a<�}a<^~a<f~a<�~a<�~a<�~a<a<la<�a<��a<��a<Z�a<��a<��a<��a<��a<]�a<0�a<��a<�a<�a<�a<�a<��a<x�a<A�a<L�a<c�a<͈a<i�a<$�a<;�a<a�a<ȍa<��a<��a<�a<��a<#�a<Ԕa<��a<ҕa<�a<8�a<�a< �a<��a<��a<ŕa<�a<B�a<��a<3�a<��a<�a<��a<��a<�a<S�a<l�a<P�a<&�a<��a<!�a<>�a<m�a<іa<!�a<��a<E�a<P�a<]�a<a<b�a<�a<��a<��a<�a<��a<H�a<ӛa<�a<F�a<	�a<��a<��a<8�a<��a<�a<�a<�a<��a<e�a<��a<șa<+�a<��a<ޚa<=�a<*�a<M�a<�a<��a<�a<D�a<��a<L�a<_�a<l�a<��a<�a<Y�a<6�a<�a<P�a<��a<C�a<Ԕa<��a<b�a<��a<?�a<d�a<e�a<G�a<ϖa<|�a<a<9�a<L�a<��a<4�a<��a<}�a<�a<B�a<��a<O�a<U�a<[�a<C�a<�a<��a<�a<Q�a<3�a<�a<،a<G�a<�a<��a<��a<y�a<��a<%�a<��a<��a<��a<�a<��a<f�a<��a<��a<��a<`�a<
�a<W�a<��a<ςa<Ɂa<�a<�a<�~a<�}a<x}a<�|a<�|a<]|a<|a<H|a<|a<&|a<�{a<�{a<#{a<zza<�ya<�xa<�wa<cva<ua<ta<�ra<ra<Rqa< qa<�pa<�pa<qa<�qa<"ra<�ra<�sa<ta<�ta<�ta<ua<)ua<�ta<�ta<8ta<�sa<Nsa<�ra<�ra<2ra<bra<Era<�ra<�ra<xsa<"ta<�ta<�  �  ~ua<�ua<�ua<�ua<�ua<,ua<�ta<�sa<Rsa<�ra<ra<�qa<Lqa<Nqa<�qa<	ra<�ra<�sa<�ta<Lva<�wa<�xa<za<W{a<S|a<2}a<�}a<X~a<�~a<�~a<a<Ea<�a<�a<*�a<ˀa<V�a<S�a<0�a</�a<�a<�a< �a<·a<S�a<��a<ވa<��a<��a<d�a<#�a<�a<��a<��a<��a<�a<��a<y�a<q�a<��a<9�a<��a<�a<w�a<��a<��a<єa<��a<6�a<n�a<��a<��a<��a<��a<��a<|�a<Ėa<��a<O�a<�a<b�a<�a<y�a<��a<I�a<��a<��a<C�a<�a<7�a<��a<Ηa<�a<3�a<u�a<�a<��a<��a<��a<�a<��a<h�a<x�a<W�a<G�a</�a<��a<��a<�a<|�a<y�a<V�a<�a<��a<N�a<�a<��a<;�a<J�a<#�a<X�a<��a<֚a<�a<Z�a<��a<��a<��a<�a<��a<ҙa<�a<�a<�a<�a<Ŕa<ޓa<$�a<��a<l�a<f�a<��a<�a<��a<p�a<�a<Ǖa<a�a<��a<M�a<{�a<��a<4�a<Ԗa<E�a<��a<�a<��a<�a<n�a<.�a<Ғa<�a<͒a<Ւa<ƒa<��a<��a<_�a<ӑa<�a<.�a<�a<��a<O�a<�a<��a<�a<Ɇa<Åa<�a<c�a<
�a<؃a<�a<S�a<��a<�a<5�a<X�a<��a<]�a<�a<��a<��a<+�a<@�a<^�a<m�a<�a<�~a<-~a<�}a<2}a<}a<�|a<�|a<�|a<{|a<*|a<�{a<7{a<mza<�ya<Uxa<2wa<�ua<�ta<tsa<Jra<Sqa<�pa<<pa<pa<pa<Zpa<�pa<�qa<Dra<�ra<�sa<Ota<�ta<ua<_ua<Cua<ua<�ta<Cta<�sa<�sa<=sa<�ra<sa<sa<Vsa<�sa<#ta<�ta<ua<�  �  �ua<�ua<�ua<�ua<�ua<ua<�ta<�sa<�ra<0ra<�qa<qa<�pa<�pa<�pa<dqa<ra<Hsa<Yta<�ua<$wa<�xa<za<5{a<o|a<A}a<�}a<�~a<�~a<Ya<�a<�a<�a<m�a<݀a<c�a<'�a<ɂa<΃a<��a<��a<��a<<�a<߇a<K�a<��a<Èa<��a<��a<�a<��a<G�a< �a<�a<�a<W�a<�a<׈a<�a<I�a<��a<5�a<��a<I�a<��a<Փa<�a<��a<?�a<��a<��a<	�a<�a<.�a<�a<I�a<`�a<��a<�a<]�a<�a<i�a<�a<G�a<��a<��a<��a<a�a<řa<D�a<[�a<f�a<��a<��a<�a<M�a<��a<Ɠa<�a<`�a<*�a<�a<ۖa<��a<��a<%�a<�a<��a<1�a<b�a<��a<��a<t�a<�a<ٛa<��a<#�a<�a<ٚa<�a<�a<"�a<h�a<��a<ɛa<ța<ța<r�a<+�a<��a<��a<�a<��a<��a<X�a<C�a<j�a<��a<�a<��a<��a<��a<��a<�a<�a<��a<��a<i�a<ږa<h�a<��a<y�a<r�a<�a<��a<�a<��a<��a<��a<!�a<Ɠa<��a<X�a<k�a<S�a<<�a<&�a<ےa<q�a<ˑa<�a<�a<�a<��a<�a<��a<�a<��a<H�a<!�a<?�a<��a<g�a<W�a<��a<��a<-�a<��a<�a<Z�a<m�a<�a<%�a<Ąa<;�a<��a<��a<ہa<�a<�a<~a<�~a<L~a<�}a<�}a<|}a<2}a<	}a<�|a<o|a<�{a<E{a<�za<gya<bxa<�va<�ua<?ta<�ra<�qa<�pa<pa<voa<[oa<foa<�oa<^pa<qa<�qa<�ra<�sa<>ta<�ta<3ua<Fua<dua<Aua<ua<�ta<sta< ta<�sa<�sa<�sa<�sa<�sa<Eta<�ta<ua<zua<�  �  �ua<-va< va<�ua<�ua<�ta<Gta<�sa<�ra<�qa<5qa<�pa<Npa<^pa<�pa<qa<�qa<�ra<ta<�ua<�va<xa<�ya<{a<O|a<[}a<$~a<�~a<5a<�a<�a<�a<P�a<a<%�a<��a<y�a<)�a<�a<�a<܅a<��a<}�a<�a<��a<��a<��a<p�a<B�a<�a<�a<�a<ǆa<��a<��a<�a<��a<��a<��a<�a<W�a<��a<��a<�a<d�a<��a<�a<ѕa<q�a<�a<(�a<Q�a<Z�a<f�a<i�a<��a<��a<�a<_�a<��a<;�a<��a<+�a<��a<Κa<Кa<��a<B�a<��a<�a<4�a<>�a<N�a<[�a<��a<�a<��a<��a<��a<
�a<Ɣa<��a<��a<a<�a<ڙa<��a<��a<6�a<��a<՜a<Ҝa<��a<b�a<�a<Ûa<��a<W�a<&�a<2�a<I�a<e�a<��a<͛a<��a<�a<�a<��a<7�a<|�a<��a<��a<��a<Q�a<�a<�a<�a<%�a<��a<p�a<r�a<��a<+�a<͒a<��a<��a<l�a<�a<��a<G�a<��a<��a<��a<T�a<�a<c�a<�a<G�a<�a<j�a<�a<��a<��a<��a<��a<��a<W�a<�a<��a<�a<�a<�a<��a<R�a<܋a<B�a<��a<6�a<�a<τa<�a<h�a<�a<��a<*�a<p�a<�a<i�a<Єa<�a<M�a<m�a<V�a<��a<z�a<��a<��a<�a<H�a<q�a<�a<a<�~a<B~a<�}a<�}a<v}a<K}a<�|a<�|a<|a<f{a<lza<Aya<xa<�va<dua<�sa<�ra<tqa<^pa<�oa<>oa<oa<oa<~oa<pa<�pa<�qa<�ra<Zsa<ta<�ta<8ua<�ua<�ua<�ua<Mua< ua<�ta<`ta<&ta<	ta<�sa<ta<Gta<�ta<�ta<Hua<�ua<�  �  ua<�ta<ua<�ta< ta<_sa<@ra<3qa<�oa<�na<�ma<�la<ula<"la<>la<�la<�ma<-oa<�pa<�ra<0ta<6va<�wa<�ya<�za<H|a<}a<�}a<h~a<�~a<�~a<a<Qa<�a<�a<��a<<�a</�a<�a<�a<�a<�a<ֆa<�a<��a<��a<��a<�a<|�a<��a<�a<I�a<��a<a�a<�a<Z�a<�a<��a<`�a<��a<��a<��a<q�a<|�a<>�a<�a<�a<a�a<ٕa<��a<�a<�a<�a<ʖa<�a<іa<�a<P�a<��a<0�a<��a<E�a<��a<2�a<G�a<+�a<�a<Y�a<Әa<��a<z�a<�a<ϓa<��a<o�a<��a<��a<ɏa<�a<��a<��a<��a<�a<N�a<�a<R�a<��a<��a<q�a<�a<�a<e�a<'�a<��a<y�a<�a<��a<x�a<~�a<_�a<z�a<��a<��a<b�a<y�a<��a<F�a<�a<~�a<{�a<��a<�a<��a<ۓa<~�a<ߐa<ŏa<Ǝa<��a<��a<��a<J�a<�a<ُa<�a<-�a<��a<��a<̕a<E�a<��a<�a<�a<�a<k�a<�a<<�a<��a<�a<��a<v�a<�a<�a<��a<�a<�a<��a<��a<�a<��a<F�a<�a<y�a<��a<��a<Ƈa<��a<��a<��a<(�a<6�a<�a<Ua<�a<�a<��a<I�a<
�a<�a<��a<6�a<K�a<��a<��a<ƃa<�a<)�a<E�a<9�a<ya<�~a<~a<y}a<}a<�|a<�|a<�|a<\|a<3|a<�{a<�za<Xza<ya<�wa<:va<�ta<�ra< qa<Coa<�ma<�la<�ka<�ja<�ja<$ka<�ka<mla<�ma<�na<pa<Iqa<pra<;sa<�sa<jta<Xta<�ta<Cta<ta<�sa<sa<�ra<�ra<�ra<�ra<�ra<Nsa<�sa<Wta<�ta<�  �  �ta<ua<ua<�ta<ta<Rsa<Hra<Fqa<pa<�na<�ma<ma<ula<bla<�la< ma<�ma<Poa<�pa<�ra<ota<Iva<�wa<�ya<�za<>|a<$}a<�}a<~a<x~a<�~a<�~a<+a<sa<�a<f�a< �a<��a<�a<�a<�a<��a<��a<A�a<��a<��a<��a< �a<��a<݅a<�a<b�a<��a<Y�a<;�a<��a<!�a<�a<W�a<�a<ǉa<��a<��a<��a<H�a<�a< �a<M�a<��a<p�a<��a<Ȗa<ʖa<��a<��a<��a<ۖa<�a<��a<�a<��a<�a<��a<��a<A�a<F�a<�a<m�a<��a<��a<��a<?�a<��a<��a<��a<��a<7�a<�a<@�a<��a<��a<��a<'�a<��a<�a<X�a<��a<��a<v�a<�a<C�a<.�a<�a<a<Z�a<��a<��a<Z�a<0�a<=�a<^�a<��a<ߚa<+�a<E�a<c�a<h�a<�a<{�a<��a<y�a<�a<��a<�a<��a<�a<ُa<ǎa<9�a<ڍa<��a<D�a<�a<	�a<C�a<l�a<��a<��a<��a<_�a<��a<%�a<�a<��a<>�a<��a<#�a<��a<��a<��a<+�a<��a<�a<�a<�a<�a<��a<��a<�a<o�a<N�a<�a<��a<ˋa<�a<��a<�a<2�a<��a<L�a<i�a<�a<�a<�a<�a<��a<{�a<B�a<�a<��a<*�a<T�a<u�a<�a<��a<��a<�a<�a<*�a<Ia<w~a<�}a<D}a<�|a<�|a<�|a<a|a<1|a<�{a<�{a<{a<Lza<ya<�wa<Ava<�ta<�ra</qa<loa<�ma<�la<�ka<1ka<ka</ka<�ka<�la<�ma<�na<1pa<Pqa<gra<Jsa<�sa<gta<�ta<Yta<ta<�sa<isa<sa<�ra<�ra<kra<�ra<�ra<6sa<�sa<ta<pta<�  �  �ta<�ta<�ta<�ta<7ta<wsa<�ra<qqa<`pa<:oa<Ona<�ma<�la<�la<�la<�ma<una<�oa<7qa<�ra<�ta<rva<=xa<�ya<!{a<|a<�|a<�}a<�}a<a~a<S~a<�~a<�~a<�~a<Xa<�a<��a<p�a<��a<~�a<��a<��a<h�a<�a<k�a<��a<��a<I�a<��a<�a<l�a<��a<G�a<҃a<كa<	�a<��a<��a<φa<z�a<�a<�a<ٍa<��a<{�a<��a<A�a<�a<ٕa<;�a<y�a<��a<V�a<Y�a<#�a<D�a<N�a<��a<�a<m�a< �a<��a<q�a<��a<�a<�a<�a<��a<Иa<�a<��a<w�a<B�a<�a<�a<)�a<Аa<i�a<Đa<;�a<�a<6�a<j�a<��a<4�a<��a<ęa<Ěa<o�a<ƛa<�a<��a<ۛa<j�a<�a<��a<�a<�a<��a<��a<ԙa<�a<l�a<̚a<3�a<.�a<<�a<Ԛa<g�a<��a<��a<_�a<��a<m�a<ߒa<��a<Y�a<N�a<Ďa<?�a<��a<��a<��a<e�a<��a<��a<Гa<��a<ѕa<��a<Жa<�a<�a<{�a<'�a<Q�a<��a<��a<w�a< �a<��a<��a<\�a<��a<z�a<��a<��a<Q�a<�a<+�a<a�a<$�a<��a<��a<�a<I�a<X�a<��a<�a<�a<�a<>�a<"�a<�a<��a<��a<Áa<r�a<3�a<׃a<=�a<u�a<:�a<��a<`�a<��a<܁a<��a<�a<�~a<~a<>}a<�|a<l|a<|a<|a<�{a<|a<�{a<x{a<�za<za<Cya<�wa<�va<�ta<sa<sqa<�oa<ona<ma<Zla<�ka<�ka<�ka<Kla< ma<na<Goa<apa<�qa<�ra<bsa<�sa< ta<Yta<$ta<�sa<}sa<�ra<�ra<)ra<ra<�qa<ra<Hra<�ra<1sa<�sa<]ta<�  �  8ta<�ta<�ta<�ta<,ta<�sa<�ra<�qa<�pa<�oa<�na<=na<�ma<�ma<�ma<nna<Hoa<{pa<�qa<�sa<9ua<�va<~xa<�ya<{a<|a<�|a<>}a<�}a<�}a<�}a<�}a<�}a<1~a<�~a< a<�a<a<߁a<܂a<��a< �a<�a<҆a<l�a<��a<��a<��a<#�a<��a<�a<_�a<��a<��a<��a<�a<v�a<_�a<��a<�a<Ŋa<��a<a�a<"�a<��a<�a<;�a<�a<��a<�a< �a<ݕa<��a<��a<u�a<q�a<��a<Εa<?�a<Ŗa<��a<�a<��a<R�a<��a<�a<�a<��a<�a<(�a<"�a<�a<�a<��a<��a<��a<��a<N�a<��a< �a<ʒa<Γa<�a<p�a<��a<�a<��a<��a<m�a<Ǜa<ěa<��a<@�a<��a<I�a<љa<^�a<�a<�a<�a<�a<k�a<әa<'�a<��a<Ӛa<�a<њa<g�a<��a<Øa<��a<_�a<��a<��a<$�a<�a<�a<��a<'�a<B�a<��a<;�a<�a<4�a<7�a<D�a<9�a<�a<s�a<Жa<ϖa<��a<�a<m�a<��a<�a<O�a<��a<3�a<�a<��a<��a<֑a<ؑa<��a<�a<��a<��a<-�a<]�a<)�a<�a<Z�a<��a<�a<�a<Y�a<׃a<��a<��a<�a<Ԁa<ڀa</�a<��a<f�a<��a<��a<�a<I�a<o�a<8�a<��a<�a<.�a<�a<�a<a<	~a</}a<|a<�{a<�{a<s{a<z{a<R{a<T{a<S{a<{a<�za<za<2ya<xa<�va<Bua<�sa<ra<opa<oa<�ma<ma<{la<`la<�la<�la<�ma<�na<�oa<�pa<�qa<�ra<]sa<�sa< ta<ta<�sa<\sa<�ra<Yra<�qa<xqa<8qa<(qa<Aqa<�qa<ra<�ra<sa<�sa<�  �  �sa< ta<�ta<wta<Mta<�sa</sa<�ra<xqa<�pa<�oa<Hoa<�na<�na<�na<coa<^pa<{qa<�ra<Gta<�ua<vwa<�xa<*za<%{a<�{a<�|a<�|a<}a<�|a<}a<�|a<�|a<'}a<{}a<'~a<�~a<�a<ɀa<"�a<P�a<��a<��a<z�a<A�a<��a<�a<ׇa<��a<#�a<��a<5�a<Ʌa<��a<��a<�a<��a<^�a<��a<�a<��a<;�a<��a<��a<�a<E�a<'�a<�a<@�a<v�a<m�a<3�a<�a<��a<{�a<a�a<��a<Ôa<.�a<Õa<|�a<b�a<�a<̘a<G�a<��a<��a<��a<7�a<l�a<��a<��a<��a<��a<��a<�a<}�a<n�a<��a<�a<ݓa<��a<�a<��a<K�a<J�a<F�a<�a<L�a<��a<]�a<0�a<��a<�a<w�a<Ęa<i�a<��a<�a<ڗa<#�a<d�a<�a<~�a<ݙa<a�a<z�a<��a<B�a<șa<�a<��a<�a<��a<Y�a<�a<�a<,�a<��a<J�a<8�a<��a<:�a<��a<ߒa<ȓa<Քa<}�a<>�a<��a<��a<��a<�a<��a<��a<�a<�a<L�a<��a<#�a<�a<��a<��a<��a<�a<K�a<w�a<��a<Q�a<�a<A�a<f�a<6�a<ˌa</�a<r�a<�a<C�a<��a<��a<Âa<*�a<Ӂa<��a<�a<��a<��a<��a<�a<b�a<��a<[�a<�a<d�a<��a<��a<o�a<Xa<~a<}a< |a<�{a<�za<�za<qza<uza<�za<�za<�za<�za<nza<�ya<<ya<Zxa<wa<�ua<<ta<�ra<Tqa<
pa<oa<na<�ma<`ma<�ma<na<�na<�oa<`pa<xqa<Bra<sa<�sa<�sa<�sa<�sa<\sa<�ra<(ra<�qa<�pa<�pa<&pa<.pa<0pa<�pa<�pa<�qa<sra<sa<�  �  sa<�sa<6ta<ota<jta<ta<�sa<sa<Qra<�qa<�pa<Opa<pa<�oa<pa<�pa<zqa<�ra<�sa<#ua<�va<xa<5ya<Kza<={a<�{a<;|a<`|a<c|a<E|a<|a<�{a<�{a<�{a<D|a<�|a<�}a<�~a<�a<�a<m�a<ڃa<�a<*�a<�a<��a<	�a<�a<�a<�a<��a<,�a<ֆa<��a<Іa<�a<��a<��a<��a<�a<��a<&�a<��a<"�a<V�a<k�a<<�a<��a<�a<�a<��a<T�a<��a<��a<d�a<5�a<M�a<��a<�a<��a<x�a<X�a<D�a<�a<͘a<R�a<��a<��a<U�a<֘a<@�a<g�a<o�a<��a<��a<-�a<ȓa<��a<˓a<>�a<�a<Ǖa<Ζa<ٗa<�a<əa<v�a<�a<P�a<E�a<��a<��a<�a<%�a<m�a<��a<:�a<ʖa<��a<��a<��a<`�a<�a<��a<5�a<��a<�a<K�a<:�a<�a<A�a<~�a<��a<^�a<:�a<�a<�a<W�a<a<l�a<�a<Ǒa<@�a<��a<��a<��a<h�a<�a<_�a<��a<��a<>�a<��a<�a<�a<�a<�a<I�a<��a<�a<��a<u�a<��a<a<�a<h�a<ϐa<�a< �a<Ɛa<P�a<��a<x�a<I�a<�a<_�a<؈a<O�a<��a<�a<��a<[�a<�a<�a<#�a<��a<�a<W�a<��a<��a<��a<q�a<كa<�a<	�a<�a<�a<I~a<}a<�{a<�za<>za<�ya<mya<iya<rya<�ya<�ya<za<0za<za<�ya<Sya<xxa<twa<_va<ua<�sa<Xra<qa<pa<Roa<�na<�na<�na<oa<�oa<spa<@qa<ra<�ra<?sa<�sa<�sa<�sa<<sa<�ra<ra<8qa<}pa<�oa<Toa<�na<�na<�na<loa<�oa<�pa<zqa<`ra<�  �  _ra<Wsa<�sa<`ta<�ta<nta<9ta<�sa</sa<ra<ra<�qa<9qa<Eqa<jqa< ra<�ra<�sa<�ta<va<iwa<�xa<�ya<�za<Q{a<�{a<�{a<�{a<�{a<g{a<{a<�za<�za<�za<{a<�{a<V|a<L}a<�~a<�a<��a<�a<j�a<ǅa<��a<��a<,�a<��a<��a<��a<X�a<�a<�a<�a<�a<�a<�a<�a<�a<A�a<��a<��a<i�a<��a<ʒa<��a<B�a<p�a<��a<S�a<��a<p�a<�a<�a<�a<�a<��a<I�a<��a<m�a<e�a<L�a<f�a<\�a<L�a< �a<p�a<��a<��a<Y�a<��a<(�a<T�a<��a<�a<P�a<�a<�a<#�a<w�a<�a<�a<��a<��a<y�a<T�a<ؚa<+�a<D�a<��a<��a<Йa<$�a<2�a<c�a<��a<�a<��a<F�a<m�a<��a<)�a<��a<��a<e�a<��a<��a<��a<*�a<�a<��a<�a<�a<<�a<$�a<>�a<K�a<��a<�a<Ēa<֒a<�a<t�a<�a<��a<h�a<�a<|�a<��a<��a<m�a<�a</�a<*�a<-�a<�a<�a<�a<5�a<��a<H�a<0�a<8�a<��a<�a<}�a<
�a<R�a<��a<z�a<R�a<��a<�a<؍a<��a<5�a<��a<~�a<)�a<$�a<[�a<��a<Y�a<)�a<V�a<v�a<��a<�a<$�a<&�a<ӄa<w�a<��a<��a<y�a<*�a<�~a<@}a<�{a<�za<�ya<�xa<rxa<%xa<xa<_xa<�xa<	ya<]ya<�ya<�ya<�ya<`ya<�xa<�wa<�va<�ua<�ta<esa<Fra<<qa<�pa<pa<�oa<�oa<Jpa<�pa<[qa<ra<�ra<Lsa<�sa<�sa<�sa<Psa<�ra<�qa<Aqa<Fpa<toa<�na<�ma<�ma<�ma<�ma<na<�na<�oa<�pa<�qa<�  �  �qa<�ra<�sa<@ta<�ta<�ta<�ta<\ta<ta<zsa<sa<�ra<�ra<�ra<�ra<9sa<�sa<�ta<�ua<wa<4xa<1ya<za<�za<[{a<�{a<�{a<[{a<{a<�za<za<�ya<rya<tya<�ya<-za<{a<-|a<r}a<a<��a<Z�a<�a<H�a<��a<��a<T�a<݈a<#�a<@�a<7�a<#�a<�a<8�a<\�a<ĉa<b�a<-�a<@�a<]�a<��a<ݏa<$�a<5�a<#�a<Ǔa<;�a<I�a<�a<Γa<L�a<��a<��a<K�a<�a<��a<��a<�a<z�a<>�a<8�a<d�a<��a<Ŗa<��a<��a<N�a<��a<ՙa<��a<]�a<�a<C�a<��a<�a<��a<R�a<L�a<`�a<Ȗa<Z�a<��a<��a<��a<=�a<ƚa<*�a<C�a<,�a<��a<�a<T�a<Q�a<C�a<K�a<_�a<��a<5�a<�a<�a<n�a<��a<a<��a<��a<x�a<'�a<��a<
�a<�a<�a<m�a<̘a<�a< �a<E�a<��a<ߔa<Y�a<�a<�a<K�a<��a<�a<��a<3�a<��a<ۖa<�a<Ėa<M�a<��a<��a<��a<V�a<�a<�a<Ўa<��a<U�a<�a<�a<�a<h�a<	�a<��a<N�a<֏a<�a<L�a<H�a<؏a<<�a<Z�a<K�a<�a<ϊa<��a<}�a<m�a<��a<
�a<��a<��a<r�a<��a<��a<��a<��a<�a<�a<p�a<r�a<@�a<�a<za<�}a<K|a<�za<yya<hxa<�wa<wa<�va<�va<2wa<�wa<3xa<�xa<"ya<]ya<�ya<aya<�xa<Zxa<|wa<�va<rua<ita<isa<�ra<�qa<xqa<4qa<Hqa<�qa<�qa<]ra<�ra<jsa<�sa<�sa<�sa<�sa<sa<Tra<�qa<npa<Xoa<\na<sma<�la<_la<)la<gla<�la<�ma<�na<�oa<�pa<�  �  Eqa<Mra<isa<$ta<�ta<ua<ua<ua<�ta<xta<ta<�sa<�sa<�sa<ta<kta<*ua<�ua<�va<�wa<�xa<�ya<yza<{a<R{a<r{a<Q{a<�za<eza<�ya</ya<�xa<lxa<@xa<pxa< ya<�ya<{a<n|a<
~a<�a<��a<`�a<�a<m�a<��a<��a<.�a<��a<�a< �a<0�a<�a<C�a<��a<��a<��a<Y�a<S�a<^�a<��a<��a<ؑa<Òa<t�a<��a<$�a<$�a<Ɠa<F�a<��a<��a<��a<F�a<ݏa<d�a<l�a<��a<B�a<7�a<)�a<p�a<��a<�a<D�a<W�a<&�a<��a<�a<�a<��a<��a<'�a<��a<�a<Зa<��a<��a<��a<��a<^�a<�a<��a<=�a<�a<6�a<y�a<_�a<�a<��a<��a<��a<|�a<f�a<L�a<[�a<��a<�a<ϒa<͒a<E�a<�a<��a<��a<��a<ߗa<��a<~�a<�a<(�a<8�a<ڙa<|�a<��a<�a<Q�a<��a<�a<��a<n�a<B�a<x�a<��a< �a<��a<ؖa<:�a<6�a<1�a<��a<+�a<T�a<(�a<�a<s�a<.�a<Ўa<ʍa<ƌa<�a<ċa<��a<�a<e�a<�a<��a<�a<H�a<��a<-�a<0�a<�a<��a<ێa<��a<݌a<܋a<��a<��a<��a<؇a<H�a<φa<��a<r�a<��a<u�a<q�a<;�a<Ѕa<@�a<Y�a<N�a<�a<l�a<�~a<�|a<K{a<�ya<qxa<#wa<]va<�ua<�ua<�ua<"va<�va<Gwa<	xa<�xa<"ya<_ya<Uya<7ya<�xa<xa<;wa<Vva<qua<fta<�sa<sa<�ra<ira<tra<�ra<�ra<asa<�sa<ta<.ta<Ata<�sa<�sa<�ra<�qa<�pa<�oa<{na<^ma<nla<�ka<ka<ka<$ka<�ka<�la<�ma<�na<�oa<�  �  �pa<�qa<sa<ta<�ta<Jua<vua<�ua<Vua<ua<�ta<�ta<�ta<�ta<ua<�ua< va<�va<�wa<�xa<�ya<Iza<�za<R{a<r{a<A{a<�za<~za<�ya<"ya<exa<�wa<Vwa<5wa<nwa<�wa<�xa<�ya<~{a<'}a<#a<�a<؂a<��a<$�a<��a<��a<�a<�a<~�a<��a<ӊa<%�a<B�a<��a<�a<��a<h�a<N�a<k�a<Q�a<a�a<h�a<2�a<ɓa<#�a<1�a<�a<x�a<ǒa<�a<�a<�a<X�a<��a<f�a<\�a<��a<9�a<�a<A�a<��a<�a<t�a<֖a<�a<�a<əa<C�a<i�a<o�a<8�a<әa<s�a<+�a<ɘa<��a<��a<��a<��a<`�a<��a<b�a<�a<b�a<��a<��a<��a<��a<>�a<U�a<.�a<�a<��a<]�a<W�a<�a<��a<��a<Ցa<3�a<�a<ʓa<�a<&�a<M�a<W�a<-�a<Йa<M�a<q�a<D�a<�a<d�a<Řa<9�a<��a<	�a<��a<g�a<W�a<o�a<��a<�a<3�a<��a<��a<��a<g�a<ۖa<��a< �a<Ǔa<Y�a<�a<c�a<�a<��a<��a<�a<��a<��a<�a<t�a<"�a<�a<�a<��a<u�a<�a<.�a<,�a<ޏa<J�a<��a<��a<�a<��a<��a<��a<�a<K�a<݇a<��a<��a<9�a< �a<�a<��a<&�a<h�a<e�a<�a<��a<�a<~a<V|a<lza<�xa<Mwa<%va<Mua<�ta<�ta<�ta<;ua<�ua<�va<uwa<9xa<�xa<&ya<sya<dya<ya<�xa<�wa<wa<1va<}ua<�ta<"ta<�sa<{sa<xsa<�sa<�sa<ta<Qta<�ta<�ta<�ta<%ta<nsa<�ra<�qa<Zpa<oa<�ma<nla<kka<�ja<$ja<�ia<,ja<�ja<�ka<�la<�ma<Roa<�  �  8pa<�qa<�ra<ta<�ta<Rua<�ua<�ua<va<�ua<�ua<sua<nua<�ua<�ua<Uva<�va<�wa<Xxa<Fya<za<�za<0{a<Q{a<s{a<D{a<�za<&za<Pya<�xa<�wa<"wa<�va<tva<�va<�va<xa<,ya<�za<w|a<z~a<j�a<m�a<c�a<�a<��a<��a<��a<o�a<�a<o�a<v�a<ǋa<�a<`�a<Ȍa<c�a<8�a<��a<�a<��a<$�a<ܒa<��a<�a<%�a<9�a<ѓa<<�a<^�a<b�a<r�a<e�a<��a<�a<��a<z�a<ٍa<�a<_�a<��a<�a<��a<��a<v�a<ɗa<�a<ʙa<B�a<��a<Ěa<��a<��a<�a<ݙa<w�a<o�a<G�a<x�a<��a<
�a<��a<�a<��a<śa< �a<̛a<��a<�a<�a<�a<��a<e�a<�a<��a<��a<��a<=�a<��a<�a<d�a<<�a<+�a<N�a<��a<Җa<�a<�a<ޙa<M�a<y�a<��a<N�a<�a<i�a<јa<=�a<a<r�a<�a<,�a<�a<c�a<��a<��a<�a<�a<�a<g�a<ܖa<��a<ʔa<o�a<ۑa<W�a<��a<S�a<��a<��a<K�a<Éa<�a<�a<Ίa<r�a<t�a<^�a<U�a<9�a<ʏa<<�a<0�a<�a<��a<��a<L�a<"�a<@�a<1�a<q�a<��a<�a<��a<>�a<'�a<܇a<�a<u�a<�a<c�a<k�a<m�a<��a<a�a<�a<�}a<�{a<�ya<%xa<�va<rua<jta<ta<�sa<ta<�ta<7ua<#va<�va<�wa<�xa<$ya<tya<cya<Xya<�xa<exa<�wa<�va</va<bua<�ta<sta<Kta<5ta<<ta<xta<�ta<ua<�ta<�ta<�ta<%ta<�sa<zra<Sqa<�oa<�na<ma<�ka<�ja<�ia<hia<�ha<mia<�ia<�ja<�ka<Dma<�na<�  �  pa<jqa<�ra<�sa<�ta<�ua<�ua<va<va<%va<va<�ua<�ua<va<Qva<�va<Zwa<xa<�xa<�ya<#za<�za<V{a<�{a<u{a<.{a<�za<�ya<ya<:xa<mwa<�va<!va<�ua<"va<�va<}wa<�xa<Qza<%|a<5~a<5�a<G�a<�a<�a<n�a<݈a<׉a<��a<
�a<��a<�a<.�a<��a<݌a<S�a<�a<��a<��a<v�a<h�a<I�a<��a<��a<(�a<]�a<�a<��a<�a<:�a<0�a<-�a<�a<)�a<v�a<�a<	�a<[�a<�a<�a<�a<��a<.�a<a<F�a<��a<ۘa<��a<��a<ޚa<��a<Ϛa<˚a<��a<D�a<�a<ݙa<әa<��a<9�a<��a<��a<l�a<��a<�a<-�a<�a<��a<�a<�a<Øa<��a<�a<Ĕa<V�a<,�a<,�a<��a<]�a<��a<ސa<��a<a<�a<O�a<��a<ėa<�a<��a<f�a<��a<ɚa<��a<)�a<˙a<B�a<Ęa<K�a<�a<��a<��a<��a<՗a< �a<3�a<#�a<8�a<�a<��a<ޖa<�a<��a<2�a<��a< �a<k�a<όa<�a<g�a<ɉa<\�a<W�a<��a<G�a< �a</�a<)�a</�a<�a<��a<�a<a�a<6�a<ԏa<�a<j�a<��a<��a<ɋa<�a</�a<��a<&�a<Ԉa<��a<P�a<�a<��a<4�a<��a<��a<H�a<�a<'�a<`a<^}a<j{a<mya<�wa<
va<�ta<�sa<�sa<Msa<�sa<ta<�ta<�ua<�va<�wa<mxa<ya<kya<�ya<{ya<ya<sxa<�wa<Ewa<�va<�ua<eua<�ta<�ta<�ta<�ta<�ta<ua<ua<ua<%ua<�ta<Fta<[sa<]ra<qa<�oa<=na<�la<hka<@ja<Hia<�ha<�ha<�ha<Uia<Xja<�ka<ma<{na<�  �  �oa<cqa<�ra<�sa<�ta<�ua<�ua<Nva<Jva<Zva<$va<va<va<=va<�va<�va<�wa<$xa<�xa<�ya<dza<{a<+{a<�{a<o{a<!{a<�za<�ya<ya<xa<Twa<iva<va<�ua<�ua<cva<Dwa<�xa<(za<|a<~a<�a<3�a<�a<�a<^�a<�a<��a<��a<^�a<��a<�a<A�a<��a<�a<��a<.�a<Ǝa<��a<��a<��a<m�a<M�a<�a<�a<r�a<�a<ϓa<��a<!�a<��a<��a<��a<��a<~�a<�a<ٌa<%�a<ƍa<�a<�a<��a<��a<��a<3�a<��a<Ԙa<��a<��a<��a<5�a<�a<��a<��a<U�a<4�a<��a<�a<(�a<U�a<��a<�a<��a<�a<;�a<�a< �a<��a<ƚa<�a<��a<|�a<ܕa<��a<"�a<�a<2�a<l�a<�a<F�a<�a<��a<��a<�a<	�a<��a<��a<��a<��a<l�a<��a<��a<��a<X�a< �a<^�a<ߘa<f�a<�a<��a<��a<ӗa<�a<"�a<k�a<d�a<p�a<�a<��a<ؖa<ٕa<��a<*�a<��a<ȏa<R�a<��a<|�a<U�a<��a<&�a<�a<��a<�a<��a<��a<�a<�a<�a<Ϗa<�a<q�a<�a<�a<j�a<��a<��a<��a<��a<�a<e�a<։a<;�a<�a<��a<y�a<,�a<�a<[�a<c�a<��a<=�a<��a< �a<Ga<&}a<9{a<Qya<mwa<va<�ta<�sa<Nsa<.sa<�sa<�sa<�ta<�ua<�va<�wa<jxa<ya<dya<�ya<Oya<Sya<�xa<*xa<jwa<�va<va<�ua<Jua<�ta<�ta<�ta<ua<Dua<Kua<gua<ua<�ta<Ota<Asa<rra< qa<�oa<�ma<�la<4ka<"ja<Oia<�ha<Uha<�ha<Yia<Aja<Oka<�la<5na<�  �  pa<jqa<�ra<�sa<�ta<�ua<�ua<va<va<%va<va<�ua<�ua<va<Qva<�va<Zwa<xa<�xa<�ya<#za<�za<V{a<�{a<u{a<.{a<�za<�ya<ya<:xa<mwa<�va<!va<�ua<"va<�va<}wa<�xa<Qza<%|a<5~a<5�a<G�a<�a<�a<n�a<݈a<׉a<��a<
�a<��a<�a<.�a<��a<݌a<S�a<�a<��a<��a<v�a<h�a<I�a<��a<��a<(�a<]�a<�a<��a<�a<:�a<0�a<-�a<�a<)�a<v�a<�a<	�a<[�a<�a<�a<�a<��a<.�a<a<F�a<��a<ۘa<��a<��a<ޚa<��a<Ϛa<˚a<��a<D�a<�a<ݙa<әa<��a<9�a<��a<��a<l�a<��a<�a<-�a<�a<��a<�a<�a<Øa<��a<�a<Ĕa<V�a<,�a<,�a<��a<]�a<��a<ސa<��a<a<�a<O�a<��a<ėa<�a<��a<f�a<��a<ɚa<��a<)�a<˙a<B�a<Ęa<K�a<�a<��a<��a<��a<՗a< �a<3�a<#�a<8�a<�a<��a<ޖa<�a<��a<2�a<��a< �a<k�a<όa<�a<g�a<ɉa<\�a<W�a<��a<G�a< �a</�a<)�a</�a<�a<��a<�a<a�a<6�a<ԏa<�a<j�a<��a<��a<ɋa<�a</�a<��a<&�a<Ԉa<��a<P�a<�a<��a<4�a<��a<��a<H�a<�a<'�a<`a<^}a<j{a<mya<�wa<
va<�ta<�sa<�sa<Msa<�sa<ta<�ta<�ua<�va<�wa<mxa<ya<kya<�ya<{ya<ya<sxa<�wa<Ewa<�va<�ua<eua<�ta<�ta<�ta<�ta<�ta<ua<ua<ua<%ua<�ta<Fta<[sa<]ra<qa<�oa<=na<�la<hka<@ja<Hia<�ha<�ha<�ha<Uia<Xja<�ka<ma<{na<�  �  8pa<�qa<�ra<ta<�ta<Rua<�ua<�ua<va<�ua<�ua<sua<nua<�ua<�ua<Uva<�va<�wa<Xxa<Fya<za<�za<0{a<Q{a<s{a<D{a<�za<&za<Pya<�xa<�wa<"wa<�va<tva<�va<�va<xa<,ya<�za<w|a<z~a<j�a<m�a<c�a<�a<��a<��a<��a<o�a<�a<o�a<v�a<ǋa<�a<`�a<Ȍa<c�a<8�a<��a<�a<��a<$�a<ܒa<��a<�a<%�a<9�a<ѓa<<�a<^�a<b�a<r�a<e�a<��a<�a<��a<z�a<ٍa<�a<_�a<��a<�a<��a<��a<v�a<ɗa<�a<ʙa<B�a<��a<Ěa<��a<��a<�a<ݙa<w�a<o�a<G�a<x�a<��a<
�a<��a<�a<��a<śa< �a<̛a<��a<�a<�a<�a<��a<e�a<�a<��a<��a<��a<=�a<��a<�a<d�a<<�a<+�a<N�a<��a<Җa<�a<�a<ޙa<M�a<y�a<��a<N�a<�a<i�a<јa<=�a<a<r�a<�a<,�a<�a<c�a<��a<��a<�a<�a<�a<g�a<ܖa<��a<ʔa<o�a<ۑa<W�a<��a<S�a<��a<��a<K�a<Éa<�a<�a<Ίa<r�a<t�a<^�a<U�a<9�a<ʏa<<�a<0�a<�a<��a<��a<L�a<"�a<@�a<1�a<q�a<��a<�a<��a<>�a<'�a<܇a<�a<u�a<�a<c�a<k�a<m�a<��a<a�a<�a<�}a<�{a<�ya<%xa<�va<rua<jta<ta<�sa<ta<�ta<7ua<#va<�va<�wa<�xa<$ya<tya<cya<Xya<�xa<exa<�wa<�va</va<bua<�ta<sta<Kta<5ta<<ta<xta<�ta<ua<�ta<�ta<�ta<%ta<�sa<zra<Sqa<�oa<�na<ma<�ka<�ja<�ia<hia<�ha<mia<�ia<�ja<�ka<Dma<�na<�  �  �pa<�qa<sa<ta<�ta<Jua<vua<�ua<Vua<ua<�ta<�ta<�ta<�ta<ua<�ua< va<�va<�wa<�xa<�ya<Iza<�za<R{a<r{a<A{a<�za<~za<�ya<"ya<exa<�wa<Vwa<5wa<nwa<�wa<�xa<�ya<~{a<'}a<#a<�a<؂a<��a<$�a<��a<��a<�a<�a<~�a<��a<ӊa<%�a<B�a<��a<�a<��a<h�a<N�a<k�a<Q�a<a�a<h�a<2�a<ɓa<#�a<1�a<�a<x�a<ǒa<�a<�a<�a<X�a<��a<f�a<\�a<��a<9�a<�a<A�a<��a<�a<t�a<֖a<�a<�a<əa<C�a<i�a<o�a<8�a<әa<s�a<+�a<ɘa<��a<��a<��a<��a<`�a<��a<b�a<�a<b�a<��a<��a<��a<��a<>�a<U�a<.�a<�a<��a<]�a<W�a<�a<��a<��a<Ցa<3�a<�a<ʓa<�a<&�a<M�a<W�a<-�a<Йa<M�a<q�a<D�a<�a<d�a<Řa<9�a<��a<	�a<��a<g�a<W�a<o�a<��a<�a<3�a<��a<��a<��a<g�a<ۖa<��a< �a<Ǔa<Y�a<�a<c�a<�a<��a<��a<�a<��a<��a<�a<t�a<"�a<�a<�a<��a<u�a<�a<.�a<,�a<ޏa<J�a<��a<��a<�a<��a<��a<��a<�a<K�a<݇a<��a<��a<9�a< �a<�a<��a<&�a<h�a<e�a<�a<��a<�a<~a<V|a<lza<�xa<Mwa<%va<Mua<�ta<�ta<�ta<;ua<�ua<�va<uwa<9xa<�xa<&ya<sya<dya<ya<�xa<�wa<wa<1va<}ua<�ta<"ta<�sa<{sa<xsa<�sa<�sa<ta<Qta<�ta<�ta<�ta<%ta<nsa<�ra<�qa<Zpa<oa<�ma<nla<kka<�ja<$ja<�ia<,ja<�ja<�ka<�la<�ma<Roa<�  �  Eqa<Mra<isa<$ta<�ta<ua<ua<ua<�ta<xta<ta<�sa<�sa<�sa<ta<kta<*ua<�ua<�va<�wa<�xa<�ya<yza<{a<R{a<r{a<Q{a<�za<eza<�ya</ya<�xa<lxa<@xa<pxa< ya<�ya<{a<n|a<
~a<�a<��a<`�a<�a<m�a<��a<��a<.�a<��a<�a< �a<0�a<�a<C�a<��a<��a<��a<Y�a<S�a<^�a<��a<��a<ؑa<Òa<t�a<��a<$�a<$�a<Ɠa<F�a<��a<��a<��a<F�a<ݏa<d�a<l�a<��a<B�a<7�a<)�a<p�a<��a<�a<D�a<W�a<&�a<��a<�a<�a<��a<��a<'�a<��a<�a<Зa<��a<��a<��a<��a<^�a<�a<��a<=�a<�a<6�a<y�a<_�a<�a<��a<��a<��a<|�a<f�a<L�a<[�a<��a<�a<ϒa<͒a<E�a<�a<��a<��a<��a<ߗa<��a<~�a<�a<(�a<8�a<ڙa<|�a<��a<�a<Q�a<��a<�a<��a<n�a<B�a<x�a<��a< �a<��a<ؖa<:�a<6�a<1�a<��a<+�a<T�a<(�a<�a<s�a<.�a<Ўa<ʍa<ƌa<�a<ċa<��a<�a<e�a<�a<��a<�a<H�a<��a<-�a<0�a<�a<��a<ێa<��a<݌a<܋a<��a<��a<��a<؇a<H�a<φa<��a<r�a<��a<u�a<q�a<;�a<Ѕa<@�a<Y�a<N�a<�a<l�a<�~a<�|a<K{a<�ya<qxa<#wa<]va<�ua<�ua<�ua<"va<�va<Gwa<	xa<�xa<"ya<_ya<Uya<7ya<�xa<xa<;wa<Vva<qua<fta<�sa<sa<�ra<ira<tra<�ra<�ra<asa<�sa<ta<.ta<Ata<�sa<�sa<�ra<�qa<�pa<�oa<{na<^ma<nla<�ka<ka<ka<$ka<�ka<�la<�ma<�na<�oa<�  �  �qa<�ra<�sa<@ta<�ta<�ta<�ta<\ta<ta<zsa<sa<�ra<�ra<�ra<�ra<9sa<�sa<�ta<�ua<wa<4xa<1ya<za<�za<[{a<�{a<�{a<[{a<{a<�za<za<�ya<rya<tya<�ya<-za<{a<-|a<r}a<a<��a<Z�a<�a<H�a<��a<��a<T�a<݈a<#�a<@�a<7�a<#�a<�a<8�a<\�a<ĉa<b�a<-�a<@�a<]�a<��a<ݏa<$�a<5�a<#�a<Ǔa<;�a<I�a<�a<Γa<L�a<��a<��a<K�a<�a<��a<��a<�a<z�a<>�a<8�a<d�a<��a<Ŗa<��a<��a<N�a<��a<ՙa<��a<]�a<�a<C�a<��a<�a<��a<R�a<L�a<`�a<Ȗa<Z�a<��a<��a<��a<=�a<ƚa<*�a<C�a<,�a<��a<�a<T�a<Q�a<C�a<K�a<_�a<��a<5�a<�a<�a<n�a<��a<a<��a<��a<x�a<'�a<��a<
�a<�a<�a<m�a<̘a<�a< �a<E�a<��a<ߔa<Y�a<�a<�a<K�a<��a<�a<��a<3�a<��a<ۖa<�a<Ėa<M�a<��a<��a<��a<V�a<�a<�a<Ўa<��a<U�a<�a<�a<�a<h�a<	�a<��a<N�a<֏a<�a<L�a<H�a<؏a<<�a<Z�a<K�a<�a<ϊa<��a<}�a<m�a<��a<
�a<��a<��a<r�a<��a<��a<��a<��a<�a<�a<p�a<r�a<@�a<�a<za<�}a<K|a<�za<yya<hxa<�wa<wa<�va<�va<2wa<�wa<3xa<�xa<"ya<]ya<�ya<aya<�xa<Zxa<|wa<�va<rua<ita<isa<�ra<�qa<xqa<4qa<Hqa<�qa<�qa<]ra<�ra<jsa<�sa<�sa<�sa<�sa<sa<Tra<�qa<npa<Xoa<\na<sma<�la<_la<)la<gla<�la<�ma<�na<�oa<�pa<�  �  _ra<Wsa<�sa<`ta<�ta<nta<9ta<�sa</sa<ra<ra<�qa<9qa<Eqa<jqa< ra<�ra<�sa<�ta<va<iwa<�xa<�ya<�za<Q{a<�{a<�{a<�{a<�{a<g{a<{a<�za<�za<�za<{a<�{a<V|a<L}a<�~a<�a<��a<�a<j�a<ǅa<��a<��a<,�a<��a<��a<��a<X�a<�a<�a<�a<�a<�a<�a<�a<�a<A�a<��a<��a<i�a<��a<ʒa<��a<B�a<p�a<��a<S�a<��a<p�a<�a<�a<�a<�a<��a<I�a<��a<m�a<e�a<L�a<f�a<\�a<L�a< �a<p�a<��a<��a<Y�a<��a<(�a<T�a<��a<�a<P�a<�a<�a<#�a<w�a<�a<�a<��a<��a<y�a<T�a<ؚa<+�a<D�a<��a<��a<Йa<$�a<2�a<c�a<��a<�a<��a<F�a<m�a<��a<)�a<��a<��a<e�a<��a<��a<��a<*�a<�a<��a<�a<�a<<�a<$�a<>�a<K�a<��a<�a<Ēa<֒a<�a<t�a<�a<��a<h�a<�a<|�a<��a<��a<m�a<�a</�a<*�a<-�a<�a<�a<�a<5�a<��a<H�a<0�a<8�a<��a<�a<}�a<
�a<R�a<��a<z�a<R�a<��a<�a<؍a<��a<5�a<��a<~�a<)�a<$�a<[�a<��a<Y�a<)�a<V�a<v�a<��a<�a<$�a<&�a<ӄa<w�a<��a<��a<y�a<*�a<�~a<@}a<�{a<�za<�ya<�xa<rxa<%xa<xa<_xa<�xa<	ya<]ya<�ya<�ya<�ya<`ya<�xa<�wa<�va<�ua<�ta<esa<Fra<<qa<�pa<pa<�oa<�oa<Jpa<�pa<[qa<ra<�ra<Lsa<�sa<�sa<�sa<Psa<�ra<�qa<Aqa<Fpa<toa<�na<�ma<�ma<�ma<�ma<na<�na<�oa<�pa<�qa<�  �  sa<�sa<6ta<ota<jta<ta<�sa<sa<Qra<�qa<�pa<Opa<pa<�oa<pa<�pa<zqa<�ra<�sa<#ua<�va<xa<5ya<Kza<={a<�{a<;|a<`|a<c|a<E|a<|a<�{a<�{a<�{a<D|a<�|a<�}a<�~a<�a<�a<m�a<ڃa<�a<*�a<�a<��a<	�a<�a<�a<�a<��a<,�a<ֆa<��a<Іa<�a<��a<��a<��a<�a<��a<&�a<��a<"�a<V�a<k�a<<�a<��a<�a<�a<��a<T�a<��a<��a<d�a<5�a<M�a<��a<�a<��a<x�a<X�a<D�a<�a<͘a<R�a<��a<��a<U�a<֘a<@�a<g�a<o�a<��a<��a<-�a<ȓa<��a<˓a<>�a<�a<Ǖa<Ζa<ٗa<�a<əa<v�a<�a<P�a<E�a<��a<��a<�a<%�a<m�a<��a<:�a<ʖa<��a<��a<��a<`�a<�a<��a<5�a<��a<�a<K�a<:�a<�a<A�a<~�a<��a<^�a<:�a<�a<�a<W�a<a<l�a<�a<Ǒa<@�a<��a<��a<��a<h�a<�a<_�a<��a<��a<>�a<��a<�a<�a<�a<�a<I�a<��a<�a<��a<u�a<��a<a<�a<h�a<ϐa<�a< �a<Ɛa<P�a<��a<x�a<I�a<�a<_�a<؈a<O�a<��a<�a<��a<[�a<�a<�a<#�a<��a<�a<W�a<��a<��a<��a<q�a<كa<�a<	�a<�a<�a<I~a<}a<�{a<�za<>za<�ya<mya<iya<rya<�ya<�ya<za<0za<za<�ya<Sya<xxa<twa<_va<ua<�sa<Xra<qa<pa<Roa<�na<�na<�na<oa<�oa<spa<@qa<ra<�ra<?sa<�sa<�sa<�sa<<sa<�ra<ra<8qa<}pa<�oa<Toa<�na<�na<�na<loa<�oa<�pa<zqa<`ra<�  �  �sa< ta<�ta<wta<Mta<�sa</sa<�ra<xqa<�pa<�oa<Hoa<�na<�na<�na<coa<^pa<{qa<�ra<Gta<�ua<vwa<�xa<*za<%{a<�{a<�|a<�|a<}a<�|a<}a<�|a<�|a<'}a<{}a<'~a<�~a<�a<ɀa<"�a<P�a<��a<��a<z�a<A�a<��a<�a<ׇa<��a<#�a<��a<5�a<Ʌa<��a<��a<�a<��a<^�a<��a<�a<��a<;�a<��a<��a<�a<E�a<'�a<�a<@�a<v�a<m�a<3�a<�a<��a<{�a<a�a<��a<Ôa<.�a<Õa<|�a<b�a<�a<̘a<G�a<��a<��a<��a<7�a<l�a<��a<��a<��a<��a<��a<�a<}�a<n�a<��a<�a<ݓa<��a<�a<��a<K�a<J�a<F�a<�a<L�a<��a<]�a<0�a<��a<�a<w�a<Ęa<i�a<��a<�a<ڗa<#�a<d�a<�a<~�a<ݙa<a�a<z�a<��a<B�a<șa<�a<��a<�a<��a<Y�a<�a<�a<,�a<��a<J�a<8�a<��a<:�a<��a<ߒa<ȓa<Քa<}�a<>�a<��a<��a<��a<�a<��a<��a<�a<�a<L�a<��a<#�a<�a<��a<��a<��a<�a<K�a<w�a<��a<Q�a<�a<A�a<f�a<6�a<ˌa</�a<r�a<�a<C�a<��a<��a<Âa<*�a<Ӂa<��a<�a<��a<��a<��a<�a<b�a<��a<[�a<�a<d�a<��a<��a<o�a<Xa<~a<}a< |a<�{a<�za<�za<qza<uza<�za<�za<�za<�za<nza<�ya<<ya<Zxa<wa<�ua<<ta<�ra<Tqa<
pa<oa<na<�ma<`ma<�ma<na<�na<�oa<`pa<xqa<Bra<sa<�sa<�sa<�sa<�sa<\sa<�ra<(ra<�qa<�pa<�pa<&pa<.pa<0pa<�pa<�pa<�qa<sra<sa<�  �  8ta<�ta<�ta<�ta<,ta<�sa<�ra<�qa<�pa<�oa<�na<=na<�ma<�ma<�ma<nna<Hoa<{pa<�qa<�sa<9ua<�va<~xa<�ya<{a<|a<�|a<>}a<�}a<�}a<�}a<�}a<�}a<1~a<�~a< a<�a<a<߁a<܂a<��a< �a<�a<҆a<l�a<��a<��a<��a<#�a<��a<�a<_�a<��a<��a<��a<�a<v�a<_�a<��a<�a<Ŋa<��a<a�a<"�a<��a<�a<;�a<�a<��a<�a< �a<ݕa<��a<��a<u�a<q�a<��a<Εa<?�a<Ŗa<��a<�a<��a<R�a<��a<�a<�a<��a<�a<(�a<"�a<�a<�a<��a<��a<��a<��a<N�a<��a< �a<ʒa<Γa<�a<p�a<��a<�a<��a<��a<m�a<Ǜa<ěa<��a<@�a<��a<I�a<љa<^�a<�a<�a<�a<�a<k�a<әa<'�a<��a<Ӛa<�a<њa<g�a<��a<Øa<��a<_�a<��a<��a<$�a<�a<�a<��a<'�a<B�a<��a<;�a<�a<4�a<7�a<D�a<9�a<�a<s�a<Жa<ϖa<��a<�a<m�a<��a<�a<O�a<��a<3�a<�a<��a<��a<֑a<ؑa<��a<�a<��a<��a<-�a<]�a<)�a<�a<Z�a<��a<�a<�a<Y�a<׃a<��a<��a<�a<Ԁa<ڀa</�a<��a<f�a<��a<��a<�a<I�a<o�a<8�a<��a<�a<.�a<�a<�a<a<	~a</}a<|a<�{a<�{a<s{a<z{a<R{a<T{a<S{a<{a<�za<za<2ya<xa<�va<Bua<�sa<ra<opa<oa<�ma<ma<{la<`la<�la<�la<�ma<�na<�oa<�pa<�qa<�ra<]sa<�sa< ta<ta<�sa<\sa<�ra<Yra<�qa<xqa<8qa<(qa<Aqa<�qa<ra<�ra<sa<�sa<�  �  �ta<�ta<�ta<�ta<7ta<wsa<�ra<qqa<`pa<:oa<Ona<�ma<�la<�la<�la<�ma<una<�oa<7qa<�ra<�ta<rva<=xa<�ya<!{a<|a<�|a<�}a<�}a<a~a<S~a<�~a<�~a<�~a<Xa<�a<��a<p�a<��a<~�a<��a<��a<h�a<�a<k�a<��a<��a<I�a<��a<�a<l�a<��a<G�a<҃a<كa<	�a<��a<��a<φa<z�a<�a<�a<ٍa<��a<{�a<��a<A�a<�a<ٕa<;�a<y�a<��a<V�a<Y�a<#�a<D�a<N�a<��a<�a<m�a< �a<��a<q�a<��a<�a<�a<�a<��a<Иa<�a<��a<w�a<B�a<�a<�a<)�a<Аa<i�a<Đa<;�a<�a<6�a<j�a<��a<4�a<��a<ęa<Ěa<o�a<ƛa<�a<��a<ۛa<j�a<�a<��a<�a<�a<��a<��a<ԙa<�a<l�a<̚a<3�a<.�a<<�a<Ԛa<g�a<��a<��a<_�a<��a<m�a<ߒa<��a<Y�a<N�a<Ďa<?�a<��a<��a<��a<e�a<��a<��a<Гa<��a<ѕa<��a<Жa<�a<�a<{�a<'�a<Q�a<��a<��a<w�a< �a<��a<��a<\�a<��a<z�a<��a<��a<Q�a<�a<+�a<a�a<$�a<��a<��a<�a<I�a<X�a<��a<�a<�a<�a<>�a<"�a<�a<��a<��a<Áa<r�a<3�a<׃a<=�a<u�a<:�a<��a<`�a<��a<܁a<��a<�a<�~a<~a<>}a<�|a<l|a<|a<|a<�{a<|a<�{a<x{a<�za<za<Cya<�wa<�va<�ta<sa<sqa<�oa<ona<ma<Zla<�ka<�ka<�ka<Kla< ma<na<Goa<apa<�qa<�ra<bsa<�sa< ta<Yta<$ta<�sa<}sa<�ra<�ra<)ra<ra<�qa<ra<Hra<�ra<1sa<�sa<]ta<�  �  �ta<ua<ua<�ta<ta<Rsa<Hra<Fqa<pa<�na<�ma<ma<ula<bla<�la< ma<�ma<Poa<�pa<�ra<ota<Iva<�wa<�ya<�za<>|a<$}a<�}a<~a<x~a<�~a<�~a<+a<sa<�a<f�a< �a<��a<�a<�a<�a<��a<��a<A�a<��a<��a<��a< �a<��a<݅a<�a<b�a<��a<Y�a<;�a<��a<!�a<�a<W�a<�a<ǉa<��a<��a<��a<H�a<�a< �a<M�a<��a<p�a<��a<Ȗa<ʖa<��a<��a<��a<ۖa<�a<��a<�a<��a<�a<��a<��a<A�a<F�a<�a<m�a<��a<��a<��a<?�a<��a<��a<��a<��a<7�a<�a<@�a<��a<��a<��a<'�a<��a<�a<X�a<��a<��a<v�a<�a<C�a<.�a<�a<a<Z�a<��a<��a<Z�a<0�a<=�a<^�a<��a<ߚa<+�a<E�a<c�a<h�a<�a<{�a<��a<y�a<�a<��a<�a<��a<�a<ُa<ǎa<9�a<ڍa<��a<D�a<�a<	�a<C�a<l�a<��a<��a<��a<_�a<��a<%�a<�a<��a<>�a<��a<#�a<��a<��a<��a<+�a<��a<�a<�a<�a<�a<��a<��a<�a<o�a<N�a<�a<��a<ˋa<�a<��a<�a<2�a<��a<L�a<i�a<�a<�a<�a<�a<��a<{�a<B�a<�a<��a<*�a<T�a<u�a<�a<��a<��a<�a<�a<*�a<Ia<w~a<�}a<D}a<�|a<�|a<�|a<a|a<1|a<�{a<�{a<{a<Lza<ya<�wa<Ava<�ta<�ra</qa<loa<�ma<�la<�ka<1ka<ka</ka<�ka<�la<�ma<�na<1pa<Pqa<gra<Jsa<�sa<gta<�ta<Yta<ta<�sa<isa<sa<�ra<�ra<kra<�ra<�ra<6sa<�sa<ta<pta<�  �  ita<%ta<ta<�sa<�ra<�qa<+pa<�na<�la<fka<�ia<�ha<�ga<fga<�ga<#ha<via<ka<�la</oa<_qa<�sa<�ua<(xa<�ya<u{a<>|a<(}a<�}a<�}a<$~a<�}a<)~a<d~a<�~a<wa<�a<!�a<
�a<O�a<e�a<��a<j�a<��a<'�a<�a<u�a<��a<��a<|�a<3�a<�a<�a<�a<�~a<#a<�a<��a<��a<?�a<��a<��a<e�a<�a<��a<�a<��a<&�a<��a<��a<ߖa<��a<��a<G�a<J�a< �a<Y�a<��a<�a<{�a<�a<��a<j�a<'�a<1�a<ߙa<Йa<˘a<ɗa<+�a<Ôa<��a<�a<>�a<ʍa<��a<ǋa<��a<ȋa<�a<Սa<�a<�a<Ւa<��a<��a<q�a<ҙa<�a<��a<ۛa<T�a<�a<��a<�a<a�a<�a<��a<��a<��a<��a<�a<_�a<�a<)�a<��a<	�a<��a<	�a<��a<V�a<|�a<��a<g�a<��a<u�a<�a<��a<��a<��a<r�a<=�a<9�a<{�a<>�a<ҏa<̑a<%�a<��a<��a<��a<��a<�a<��a<�a<��a<��a<�a<S�a<ڒa<��a<U�a<o�a<`�a<��a<��a<ؒa<��a<��a<,�a<͏a<2�a<1�a<�a<��a<-�a<҂a<{�a<�~a<�|a<�{a<Y{a<{a<�{a<&|a<;}a<r~a<�a<�a<�a<�a<��a<�a<d�a<I�a<��a<y�a<��a<=a<a~a<a}a<�|a<5|a<�{a<�{a<{a<�{a<�{a<�{a<{a<)za<�ya<�wa<jva<Gta<_ra<�oa<�ma<yka<�ia<%ha<�fa<Wfa<fa<xfa<ga<zha<#ja<�ka<�ma<)oa<�pa<�qa<�ra<xsa<�sa<�sa<tsa<sa<gra<�qa<�qa<=qa<Jqa<Fqa<�qa<ra<�ra<Ssa<�sa<�  �  �sa<5ta<	ta<�sa<�ra<�qa<Lpa<�na<ma<�ka<�ia<�ha<�ga<�ga<�ga<nha<{ia<*ka<ma<Zoa<�qa<ta<va<Dxa<�ya<A{a<N|a<}a<j}a<�}a<�}a<�}a<-~a<G~a<�~a<8a<�a<��a<�a<'�a<3�a<$�a< �a<��a<��a<׆a<��a<υa<ӄa<��a<f�a<B�a<5�a<na<a<Pa<�a<��a<y�a<z�a<��a<%�a<��a<	�a<.�a<6�a<��a<�a<ҕa<T�a<h�a<|�a<r�a<P�a<,�a<��a<$�a<e�a<˖a<y�a<�a<��a<6�a<��a<�a<��a<��a<͘a<�a<V�a<Ӕa<��a<9�a<y�a<��a<��a<�a<΋a<�a<��a<эa<X�a<0�a<�a<�a<ܖa<��a<�a<�a<��a<��a<�a<��a<E�a<Ԛa<c�a<ܙa<��a<X�a<b�a<��a<�a<U�a<��a<�a<#�a<�a<��a<�a<Θa<y�a<��a<a<��a<��a<��a<�a<��a<��a<��a<��a<B�a<c�a<��a<i�a<�a<בa<J�a<˔a<��a<j�a<��a<Жa<c�a<ݕa<M�a<��a<��a<6�a<��a<c�a</�a<H�a<g�a<�a<��a<m�a<X�a<ޑa<�a<��a<P�a<a�a<6�a<Շa<_�a<�a<��a<�~a<*}a< |a<{a<M{a<�{a<b|a<r}a<�~a<�a<6�a<9�a<#�a<y�a<��a<��a<�a<%�a<E�a<M�a<Ea<D~a<>}a<�|a<|a<�{a<�{a<�{a<|{a<W{a<%{a<�za<Bza<Qya<�wa<�va<rta<pra< pa<�ma<�ka<�ia<&ha<ga<tfa<Nfa<�fa<{ga<�ha<Kja<�ka<�ma<Goa<�pa<�qa<�ra<dsa<�sa<�sa<"sa<�ra<Sra<�qa<eqa<qa<qa<'qa<zqa<ra<�ra<sa<�sa<�  �  �sa<ta<�sa<�sa<�ra<�qa<�pa<oa<�ma<�ka<�ja<�ia<�ha<qha<Zha<Iia<.ja<�ka<�ma<�oa<ra<;ta<Yva<Exa<�ya<*{a<,|a<�|a<}a<�}a<E}a<U}a<^}a<�}a<�}a<{~a<Xa<&�a<Z�a<n�a<�a<�a<҅a<��a<̆a<�a<��a<��a<�a<��a<ׂa<��a<��a<�a<�a<�a<��a<܁a< �a<B�a<<�a<��a<��a<7�a<_�a<4�a<��a<��a<��a<�a<-�a<@�a<��a<��a<T�a<a�a<h�a<��a<�a<��a<g�a<�a<�a<]�a<ԙa<֙a<t�a<�a<�a<��a<�a<j�a<��a<�a<��a<j�a<�a<d�a<̌a<s�a<��a<�a<��a<��a<Z�a<�a<��a<�a<�a<l�a<՛a<��a<q�a<ؚa<%�a<��a<�a<�a<��a<ʘa<јa<=�a<��a</�a<��a<ǚa<�a<��a<�a<ؘa<��a<�a<�a<�a<�a<d�a<Ȍa<~�a<Ɗa<.�a<��a<��a< �a<Z�a<̎a<��a<�a<��a<͔a<ŕa<S�a<��a<��a<�a<��a<��a<�a<'�a<~�a<�a<��a<��a<t�a<��a<Ƒa<9�a<;�a<
�a<��a<ѐa<֏a<S�a<��a<i�a<.�a<хa<p�a<�a<aa<~a<�|a<&|a<4|a<?|a<)}a<�}a<a<P�a<e�a<j�a<"�a<��a<��a<p�a<ǂa<�a<	�a<�a<�~a<l}a<�|a<�{a<Y{a<{a<�za<�za<�za<3{a<�za<�za<za<+ya<xa<�va<�ta<�ra<�pa<Mna<Fla<�ja<�ha<�ga<
ga<ga<lga<*ha<nia<�ja<_la<�ma<�oa<�pa<ra<�ra<7sa<�sa<4sa<�ra<[ra<�qa<%qa<�pa<�pa<Dpa<�pa<�pa<Iqa<�qa<�ra<_sa<�  �  sa<�sa<�sa<�sa<�ra<"ra<qa<�oa<Ena<�la<�ka<sja<�ia<jia<�ia<0ja<0ka<�la<�na<�pa<�ra<�ta<�va<zxa<�ya<7{a<�{a<g|a<�|a<�|a<�|a<�|a<n|a<�|a<�|a<b}a<[~a<9a<��a<��a<	�a<;�a<P�a<�a<��a<�a<��a<Z�a<��a<��a<��a<��a<Ła<#�a<ހa<�a<��a<��a<1�a<�a<�a<l�a<��a<Ȏa<ΐa<H�a<͓a<��a<<�a<��a<��a<Y�a<�a<Ҕa<e�a<q�a<O�a<��a<8�a<��a<��a<W�a<)�a<˘a<X�a<y�a<��a<�a<�a<�a<��a<�a<x�a<ېa<��a<p�a<Ӎa<��a<ˍa<_�a<|�a<�a<q�a<B�a<��a<��a<��a<�a<��a<>�a<Q�a<�a<��a<�a<f�a<Ęa<)�a<ؗa<��a<��a<�a<X�a<�a<h�a<�a<B�a<m�a<C�a<�a<�a<͗a<`�a<��a<Ԓa<�a<9�a<��a<w�a<��a<V�a<��a<��a<��a<'�a<��a<1�a<��a<
�a<�a<ϕa<`�a<K�a< �a<��a<ٔa<��a<)�a<7�a<��a<��a<��a<��a<��a<ܐa<�a<\�a<��a<��a<@�a<��a<�a<e�a<�a<�a<ֈa<��a<C�a<K�a<m�a<�~a<�}a<;}a<}a<P}a<�}a<�~a<�a<��a<��a<قa<6�a<��a<��a<��a<H�a<?�a<"�a<�~a<�}a<}|a<�{a<�za<Fza<za<�ya<za< za<Jza<Iza<9za<�ya<7ya<xa<�va<-ua<Bsa<5qa<$oa<ma<`ka<�ia<�ha<0ha<ha<Wha<&ia<Cja<�ka<ma<�na<pa<9qa<ra<�ra<	sa<sa<�ra<1ra<�qa<�pa<Epa<�oa<poa</oa<yoa<�oa<dpa<qa<�qa<�ra<�  �  �ra<!sa<esa<asa<sa<�ra<cqa<Cpa<oa<�ma<�la<�ka<ka<�ja<ka<�ka<�la<na<�oa<�qa<vsa<Xua<+wa<�xa< za<�za<�{a<�{a<�{a<�{a<�{a<L{a<"{a<={a<r{a<�{a<�|a<�}a<6a<��a<�a<h�a<̈́a<΅a<}�a<ӆa<��a<��a<��a<J�a<��a<��a<�a<��a<A�a<��a<.�a<�a<��a<8�a<A�a<Q�a<J�a<9�a<$�a<��a<��a<��a<�a<�a<��a<k�a<��a<|�a<�a<�a<�a<+�a<��a<j�a<U�a<V�a<5�a<�a<Ԙa<,�a<K�a<�a<r�a<c�a<�a<Ȕa<��a<�a<ΐa<�a<+�a<�a<1�a<ȏa<ؐa<�a<��a<�a<��a<��a<g�a<A�a<��a<�a<�a<��a<a<�a<@�a<p�a<іa<P�a<�a<,�a<��a<�a<��a<r�a<�a<��a<�a<�a<��a<�a<;�a<��a<6�a<��a<�a<`�a<
�a<�a< �a<��a<یa<o�a<=�a<]�a<��a<�a<,�a<[�a<m�a<ەa<%�a< �a<��a<�a<�a<��a<�a<�a<,�a<��a<#�a<�a<5�a<��a<�a<j�a<��a<�a<�a<��a<��a<��a<F�a<^�a<z�a<|�a<}�a<s�a<؁a<N�a<Xa<�~a<m~a<�~a<a<�a<Ԁa<��a<g�a</�a<��a<��a<J�a<��a<��a<x�a<3a<�}a<r|a<-{a</za<Sya<�xa<�xa<�xa<�xa<ya<Vya<�ya<�ya<uya<ya<xa<wa<ua<�sa<�qa<-pa<Lna<�la<Oka<.ja<�ia<}ia<�ia<�ja<gka<�la<�ma<4oa<`pa<�qa<Qra<�ra<�ra<�ra<&ra<Oqa<�pa<�oa<�na<[na<�ma<�ma<�ma<sna<oa<�oa<�pa<�qa<�  �  �qa<�ra<sa<Hsa<Asa<�ra<ra<Hqa<,pa<oa<na<)ma<�la<qla<�la<<ma<*na<loa<qa<�ra<�ta<Jva<�wa<(ya<za<�za<,{a<0{a<�za<�za<Eza<�ya<�ya<�ya<�ya<gza<I{a<t|a<�}a<Da<	�a<��a<�a<I�a<'�a<Ԇa<;�a<	�a<Ɇa<V�a<��a<�a<R�a<�a<��a<�a<��a<҅a<�a<��a<��a<X�a<W�a<�a<��a<�a<��a</�a<w�a<0�a<�a<r�a<��a<�a<��a<X�a<O�a<��a<�a<��a<�a<�a<Q�a<5�a<�a<Øa<�a<�a<��a<�a<�a<��a<��a<f�a<5�a<]�a<�a<��a<Ґa<o�a<=�a<d�a<͔a<+�a<��a<��a<��a<l�a<��a<��a<X�a<��a<�a<�a<ߖa<��a<D�a<̔a<��a<��a<��a<��a<S�a<:�a<)�a<ǘa<c�a<��a<��a<B�a<|�a<m�a<;�a<��a<6�a<��a<p�a<�a<ǎa<q�a<��a<�a<��a<��a<Бa<	�a< �a<��a<��a<��a<�a<��a<�a<��a<�a<��a<~�a<v�a<��a<��a<��a<��a<a<�a<��a<\�a<ُa<#�a<j�a<+�a<��a<��a<��a<+�a<��a<��a<Æa<ׄa<;�a<�a<�a<S�a<*�a<"�a<��a<C�a<ہa<��a<;�a<��a<كa<��a<��a<3�a<�a<�a<;~a<x|a<{a<�ya<�xa<�wa<Dwa<wa<'wa<`wa<�wa<rxa<�xa<�xa<ya<�xa<0xa<[wa<	va<�ta<sa<:qa<�oa<na<�la<�ka<Gka<ka<gka<�ka<�la<�ma<oa<<pa<$qa<�qa<}ra<�ra<vra<ra<=qa<vpa<noa<_na<�ma<�la<ela<?la<mla<�la<�ma<�na<�oa<�pa<�  �  �pa<�qa<�ra<6sa<dsa<3sa<�ra<ra<Cqa<Gpa<�oa<�na<Sna<=na<Sna<oa<�oa<qa<�ra<�sa<�ua<wa<~xa<sya<>za<�za<�za<�za<za<�ya<�xa<�xa<xa<�wa<!xa<�xa<�ya<�za<T|a<�}a<�a<��a<1�a<˄a<�a<܆a<c�a<��a<��a<2�a<Æa<M�a<��a<��a<��a<�a<y�a<��a<��a<V�a<�a<��a<B�a<Ӑa<*�a<�a<Ǔa<��a<��a<��a<ߒa<�a<P�a<��a<��a<��a<��a<ԏa<r�a<M�a<��a<��a<�a<D�a<y�a<T�a<�a<"�a<��a<��a<Ǘa<ߖa<��a<Ӕa<�a<�a<��a<Y�a<��a<�a<�a<�a<�a<N�a<f�a<|�a<&�a<��a<��a<R�a<ԙa<Әa<̗a<��a<��a<|�a<��a<�a<��a<�a<A�a<�a<�a<ڕa<�a<�a<טa<D�a<��a<e�a<ߘa<*�a<�a<ӕa<n�a<U�a<�a<%�a<��a<*�a<Z�a<��a<X�a<3�a<�a<�a<�a<��a<��a<�a<Еa<5�a<X�a<�a<ȑa<_�a<'�a<ԍa<݌a<0�a<��a<ڋa<�a<��a<N�a<��a<Ύa<h�a<�a<�a<��a<�a<5�a<�a<a�a<��a<�a<��a<�a<��a<��a<�a<݁a<Ӂa<=�a<��a<�a<��a<�a<5�a<�a<��a<ła<��a<=�a<�~a<�|a<,{a<�ya<xa<�va<�ua<~ua<Yua<zua<va<~va<&wa<�wa<Zxa<�xa<�xa<Jxa<�wa<�va<bua< ta<ira<qa<�oa<pna<�ma<�la<�la<ma<�ma<fna<(oa<)pa<qa<�qa<ara<�ra<�ra<ra<�qa<ppa<Yoa<na<ma<�ka<ka<�ja<cja<�ja<(ka<la<9ma<Dna<�oa<�  �  	pa<9qa<Mra<sa<xsa<�sa<fsa<�ra<nra<�qa<�pa<dpa<pa<�oa<0pa<�pa<�qa<�ra<�sa<Oua<�va<�wa<�xa<�ya<Cza<~za<Aza<�ya<Jya<ixa<�wa<�va<eva<Eva<Vva<�va<�wa<ya<�za<�|a<v~a<��a<n�a<�a<��a<Ɔa<��a<�a<0�a<(�a<�a<��a<]�a<L�a<N�a<��a<E�a<0�a<j�a<��a<-�a<��a<@�a<y�a<��a<F�a<��a<̓a<Q�a<��a<�a<ِa<��a<�a<=�a<�a<ɍa<�a<Ǝa<��a<�a<l�a<ԓa<m�a<��a<��a<��a<�a<:�a<�a<��a<�a< �a<!�a<c�a<Ȕa<[�a<1�a<b�a<˔a<�a<\�a<c�a<��a<G�a<�a<��a<��a<��a<�a<�a<�a<Ėa<[�a<�a<˒a<�a<J�a<��a< �a<��a<X�a<l�a<��a<�a<-�a<�a<�a<g�a<y�a<F�a<��a<ڗa<��a<˕a<��a<��a<ڒa<Q�a<�a<�a<T�a<ؒa<��a<`�a<%�a<��a<.�a<J�a<�a<��a<��a<��a<C�a<��a<�a<��a<.�a<4�a<f�a<�a<�a<T�a<�a<�a<Ɍa<Ӎa<��a<?�a<��a<��a<I�a<��a<��a<W�a<�a<X�a<�a<��a<Z�a<|�a<كa<��a<��a<��a<��a<r�a<��a<��a<��a<4�a<��a<��a<�a<xa<�}a<�{a<�ya<�wa<Vva<4ua<;ta<�sa<�sa<�sa<[ta<5ua<�ua<�va<�wa<	xa<oxa<Fxa<�wa<7wa<va<ua<�sa<Zra<0qa<-pa<]oa<�na<�na<�na<(oa<�oa<}pa<`qa<�qa<wra<�ra<�ra<qra<�qa<�pa<�oa<Rna<�la<�ka<Nja<ria<�ha<�ha<�ha<�ia<fja<�ka<ma<�na<�  �  oa<�pa<ra<�ra<�sa<�sa<ta<�sa<Jsa<�ra<Qra<�qa<�qa<�qa<�qa<=ra<sa<ta<<ua<rva<�wa<�xa<�ya<za<Nza<Pza<�ya<ya<Axa<Twa<}va<�ua<ua<�ta<�ta<Tua<va<�wa<8ya<?{a<k}a<wa<��a<��a<k�a<��a<Շa<��a<��a<�a<��a<�a<Ɉa<��a<�a<;�a<׉a<͊a<Ջa<$�a<��a<ݏa<�a<L�a<�a<��a<��a<��a<�a<�a<ߐa<Џa<��a<��a<׌a<4�a<9�a<s�a<�a<B�a<��a<-�a<Œa<c�a<�a<p�a<��a<!�a<��a<��a<j�a<Ƙa<5�a<��a<Ԗa<B�a<�a<a<�a<g�a<��a<ėa<��a<c�a<3�a<��a<�a<ۚa<d�a<a<w�a<�a<��a<B�a<��a<c�a<]�a<��a<}�a<u�a<	�a<�a<�a<��a<Ҕa<*�a<k�a<��a<B�a<��a<��a<`�a<ǘa<ڗa<�a<�a<"�a<r�a<ؓa<��a<��a<ۓa<I�a<�a<��a<��a<��a<Öa<��a<*�a<z�a<j�a<ɒa<;�a<��a<�a<$�a<ˊa<��a<ǈa<~�a<Z�a<�a<��a<��a<��a<��a<ōa<��a<o�a<��a<��a<�a<Y�a<7�a<��a<��a<O�a<�a<��a<�a<k�a<%�a<�a<�a<@�a<`�a<q�a<{�a<"�a<��a<z�a<L�a<��a<�~a<�|a<�za<�xa<�va<�ta<vsa<�ra<ra<�qa<ora<�ra<�sa<�ta<�ua<�va<�wa<7xa<Ixa<.xa<�wa<wa<�ua<�ta<�sa<�ra<�qa<�pa<fpa<6pa<^pa<�pa<#qa<�qa<>ra<�ra<,sa<*sa<�ra<Pra<�qa<(pa<�na<2ma<�ka<0ja<�ha<�ga<4ga<+ga<=ga<�ga<ia<Kja<�ka<rma<�  �  zna<4pa<�qa<�ra<�sa<8ta<yta<ita<7ta<�sa<�sa<)sa<sa<sa< sa<�sa<gta<`ua<]va<jwa<gxa<Aya<�ya<Vza<�za<za<�ya<�xa<�wa<�va<Kua<bta<�sa<2sa<Nsa<�sa<�ta<!va<�wa<za<l|a<�~a<�a<K�a< �a<��a<�a<шa<{�a<��a<�a<�a<�a<�a<m�a<��a<F�a<N�a<#�a<z�a<��a<͐a<ܑa<Ғa<d�a<Гa<��a<#�a<��a<q�a<2�a<�a<m�a<Z�a<e�a<׊a<��a<��a<��a<׌a<Y�a<��a<�a<ēa<��a<�a<2�a<T�a<Йa<��a<�a<��a<+�a<��a<$�a<��a<j�a<)�a<i�a<Зa<D�a< �a<��a<U�a<ךa<8�a<7�a<�a<P�a<V�a<%�a<��a<�a<'�a<{�a<�a<�a<>�a<�a<�a<��a<��a<�a<f�a<�a<��a<�a<<�a<�a<ԙa<�a<˙a<\�a<ǘa<��a<>�a<s�a<ԕa<]�a<��a<�a<1�a<��a<�a<|�a<ޖa<�a<!�a<��a<a�a<9�a<�a<o�a<��a<��a<��a<��a<i�a<!�a<^�a<�a<�a<m�a<S�a<_�a<��a<�a<O�a<k�a<�a<��a<Ǐa<a�a<܎a<�a<�a<��a<��a<O�a<y�a<|�a<چa<��a<B�a<a�a<I�a<P�a<3�a< �a<p�a<��a<��a<�a<O�a<+~a<�{a<�ya<Jwa<Qua<}sa<ra<!qa<�pa<�pa<qa<�qa<�ra<ta<Aua<ava<\wa<�wa<{xa<oxa<xa<�wa<�va<�ua<�ta<�sa<�ra<kra<�qa<�qa<�qa<�qa<_ra<�ra<0sa<wsa<�sa<rsa<)sa<<ra<"qa<�oa<4na<xla<�ja<�ha<�ga<ufa<�ea<�ea<�ea<�fa<�ga<ia<�ja<�la<�  �  �ma<�oa<]qa<�ra<�sa<|ta<�ta<�ta<ua<�ta<Lta<ta<�sa<ta<6ta<�ta<Mua<=va<wa<6xa<.ya<�ya<qza<zza<xza<�ya<;ya<4xa<wa<�ua<mta<�sa<�ra<Kra<Kra<�ra<�sa<ua<,wa<8ya<�{a<~a<~�a<Ђa<�a<��a<�a<4�a<��a<V�a<ڊa<��a<ߊa<��a<P�a<��a<^�a<8�a<�a<D�a<H�a<��a<��a<O�a<Փa<͓a<��a<�a<�a<ߐa<��a<�a<��a<��a<V�a<��a<��a<��a<ъa<Ћa<��a<�a<!�a<�a<��a<��a< �a<E�a<�a<~�a<o�a<[�a<�a<T�a<��a<��a<n�a<@�a<}�a<��a<3�a<ʙa<^�a<4�a<\�a<��a<��a<�a<C�a<�a<��a<��a<:�a<M�a<��a<>�a<�a<T�a<��a<"�a<��a<��a<�a<��a<Z�a<��a<��a<��a<�a<˙a<(�a<Q�a<�a<��a<a<�a<]�a<��a<t�a<�a<'�a<�a<y�a<a<I�a<��a<��a<��a<�a<U�a<'�a<��a<�a<��a<��a<ًa<,�a<i�a<;�a<[�a<̅a<&�a<f�a<��a<��a<�a<e�a<��a<��a<�a<��a<��a<ŏa<Y�a<��a<ҍa<h�a<e�a<@�a<]�a<��a<�a<��a<1�a<,�a<��a<9�a<؆a<~�a<�a<��a<��a<ԁa<�a<�}a<I{a<�xa<va<�ta<ora<?qa<pa<�oa<�oa<�oa<qa<�qa<Asa<�ta<�ua<�va<�wa<lxa<�xa<�xa<	xa<{wa<�va<�ua<�ta<�sa<osa<�ra<�ra<�ra<�ra<(sa<xsa<ta<�sa<"ta<�sa<sa</ra<�pa<Voa<�ma<�ka<�ia<1ha<�fa<sea<�da<gda<�da<�ea<�fa<Mha<�ia<�ka<�  �  �ma<poa<Tqa<�ra<�sa<�ta<)ua<Hua<-ua< ua<�ta<�ta<�ta<�ta<�ta<lua<va<�va<�wa<�xa<Vya<za<�za<�za<kza<�ya<#ya<�wa<�va<Nua<	ta<�ra<�qa<pqa<�qa<ra<sa<qta<lva<�xa<*{a<�}a<L�a<��a<�a<��a<,�a<W�a<7�a<��a<�a<T�a<��a<̋a<��a<x�a<�a<؍a<�a<��a<��a<�a<��a<��a<��a<��a<��a<�a<�a<��a<+�a<��a<�a<Ǌa<��a<�a<�a<=�a<�a<&�a<ʌa<��a<��a<ƒa<��a<��a<�a<-�a<�a<��a<Úa<��a<Y�a<�a<��a<R�a<�a< �a< �a<q�a<��a<s�a<��a<U�a<��a<�a<��a<�a</�a<�a<d�a<��a<Óa<�a<�a<��a<-�a<}�a<-�a<R�a<،a<�a<j�a<,�a<�a<��a<S�a<�a<��a<љa<L�a<|�a<<�a<��a<I�a<��a<$�a<y�a<�a<Ζa<��a<�a<6�a<r�a<��a<Ηa<��a<ėa<4�a<H�a<�a<��a<��a<��a<��a<u�a<s�a<��a<_�a<��a<2�a<B�a<��a<��a<�a<|�a<��a<��a<��a<�a<y�a<�a<�a<��a<ʎa<��a<�a<�a<�a<�a<H�a<��a<0�a<
�a<ׇa<��a<m�a<�a<��a< �a<�a<m�a<ׁa<�a<k}a<�za<gxa<�ua<�sa<�qa<Ypa<eoa<�na<�na<Soa<Apa<qa<�ra<Cta<�ua<�va<�wa<Txa<�xa<�xa<\xa<�wa<wa<Cva<�ua<�ta<ta<�sa<jsa<hsa<�sa<�sa<ta</ta<Pta<Tta<�sa<-sa<ra<�pa<oa<Zma<Rka<qia<�ga<fa<�da<da<�ca<da<�da<fa<�ga<�ia<�ka<�  �  �ma<Ooa<4qa<�ra<�sa<�ta<!ua<�ua<pua<aua<�ta<�ta<�ta<�ta<:ua<�ua<Iva<�va<�wa<�xa<�ya<zza<sza<�za<�za<�ya<�xa<�wa<�va<ua<�sa<�ra<�qa<Mqa<Oqa<�qa<�ra<vta<5va<rxa<�za<r}a<6�a<g�a<˄a<��a<b�a<9�a<a�a<�a<6�a<��a<��a<Ջa<�a<��a<I�a<��a<�a<�a<:�a<�a<9�a<ʓa<ϓa<3�a<��a<�a<��a<��a<�a<i�a<�a<��a<ĉa<׈a<Јa<�a<Éa<<�a<��a<��a<{�a<��a<��a<e�a<��a<A�a<?�a<v�a<�a<�a<��a<,�a<��a<|�a<-�a<C�a<B�a<��a<��a<q�a<9�a<��a<*�a<�a<��a<K�a<'�a<��a<@�a<��a<��a<đa<ȏa<]�a<&�a<3�a<�a<�a<Ɍa<�a<'�a<�a<��a<��a<1�a<Зa<�a<��a<K�a<s�a<��a< �a<��a<��a<!�a<��a<-�a<�a<�a<�a<2�a<��a<�a<%�a<R�a<��a<P�a<c�a<�a<n�a<��a<��a<J�a<J�a<4�a<Ƈa<<�a<^�a<�a<��a<a<��a<ȇa<I�a<��a<m�a<��a<Ύa<v�a<�a<ʏa<a<I�a<.�a<X�a<�a<�a<#�a<s�a<݈a<O�a<"�a<Їa<�a<��a<��a<��a<ۅa<!�a<s�a<��a<ta<O}a<�za<3xa<�ua<�sa<�qa<pa<Boa<�na<�na<hoa<pa<Pqa<�ra< ta<�ua<�va<�wa<hxa<�xa<�xa<�xa<
xa<6wa<cva<xua<�ta<.ta<�sa<�sa<�sa<�sa<�sa<Sta<kta<�ta<[ta<�sa<\sa<ra<�pa<�na<Oma<ka<Iia<Jga<�ea<�da<�ca<�ca<�ca<�da<�ea<aga<pia<Cka<�  �  �ma<poa<Tqa<�ra<�sa<�ta<)ua<Hua<-ua< ua<�ta<�ta<�ta<�ta<�ta<lua<va<�va<�wa<�xa<Vya<za<�za<�za<kza<�ya<#ya<�wa<�va<Nua<	ta<�ra<�qa<pqa<�qa<ra<sa<qta<lva<�xa<*{a<�}a<L�a<��a<�a<��a<,�a<W�a<7�a<��a<�a<T�a<��a<̋a<��a<x�a<�a<؍a<�a<��a<��a<�a<��a<��a<��a<��a<��a<�a<�a<��a<+�a<��a<�a<Ǌa<��a<�a<�a<=�a<�a<&�a<ʌa<��a<��a<ƒa<��a<��a<�a<-�a<�a<��a<Úa<��a<Y�a<�a<��a<R�a<�a< �a< �a<q�a<��a<s�a<��a<U�a<��a<�a<��a<�a</�a<�a<d�a<��a<Óa<�a<�a<��a<-�a<}�a<-�a<R�a<،a<�a<j�a<,�a<�a<��a<S�a<�a<��a<љa<L�a<|�a<<�a<��a<I�a<��a<$�a<y�a<�a<Ζa<��a<�a<6�a<r�a<��a<Ηa<��a<ėa<4�a<H�a<�a<��a<��a<��a<��a<u�a<s�a<��a<_�a<��a<2�a<B�a<��a<��a<�a<|�a<��a<��a<��a<�a<y�a<�a<�a<��a<ʎa<��a<�a<�a<�a<�a<H�a<��a<0�a<
�a<ׇa<��a<m�a<�a<��a< �a<�a<m�a<ׁa<�a<k}a<�za<gxa<�ua<�sa<�qa<Ypa<eoa<�na<�na<Soa<Apa<qa<�ra<Cta<�ua<�va<�wa<Txa<�xa<�xa<\xa<�wa<wa<Cva<�ua<�ta<ta<�sa<jsa<hsa<�sa<�sa<ta</ta<Pta<Tta<�sa<-sa<ra<�pa<oa<Zma<Rka<qia<�ga<fa<�da<da<�ca<da<�da<fa<�ga<�ia<�ka<�  �  �ma<�oa<]qa<�ra<�sa<|ta<�ta<�ta<ua<�ta<Lta<ta<�sa<ta<6ta<�ta<Mua<=va<wa<6xa<.ya<�ya<qza<zza<xza<�ya<;ya<4xa<wa<�ua<mta<�sa<�ra<Kra<Kra<�ra<�sa<ua<,wa<8ya<�{a<~a<~�a<Ђa<�a<��a<�a<4�a<��a<V�a<ڊa<��a<ߊa<��a<P�a<��a<^�a<8�a<�a<D�a<H�a<��a<��a<O�a<Փa<͓a<��a<�a<�a<ߐa<��a<�a<��a<��a<V�a<��a<��a<��a<ъa<Ћa<��a<�a<!�a<�a<��a<��a< �a<E�a<�a<~�a<o�a<[�a<�a<T�a<��a<��a<n�a<@�a<}�a<��a<3�a<ʙa<^�a<4�a<\�a<��a<��a<�a<C�a<�a<��a<��a<:�a<M�a<��a<>�a<�a<T�a<��a<"�a<��a<��a<�a<��a<Z�a<��a<��a<��a<�a<˙a<(�a<Q�a<�a<��a<a<�a<]�a<��a<t�a<�a<'�a<�a<y�a<a<I�a<��a<��a<��a<�a<U�a<'�a<��a<�a<��a<��a<ًa<,�a<i�a<;�a<[�a<̅a<&�a<f�a<��a<��a<�a<e�a<��a<��a<�a<��a<��a<ŏa<Y�a<��a<ҍa<h�a<e�a<@�a<]�a<��a<�a<��a<1�a<,�a<��a<9�a<؆a<~�a<�a<��a<��a<ԁa<�a<�}a<I{a<�xa<va<�ta<ora<?qa<pa<�oa<�oa<�oa<qa<�qa<Asa<�ta<�ua<�va<�wa<lxa<�xa<�xa<	xa<{wa<�va<�ua<�ta<�sa<osa<�ra<�ra<�ra<�ra<(sa<xsa<ta<�sa<"ta<�sa<sa</ra<�pa<Voa<�ma<�ka<�ia<1ha<�fa<sea<�da<gda<�da<�ea<�fa<Mha<�ia<�ka<�  �  zna<4pa<�qa<�ra<�sa<8ta<yta<ita<7ta<�sa<�sa<)sa<sa<sa< sa<�sa<gta<`ua<]va<jwa<gxa<Aya<�ya<Vza<�za<za<�ya<�xa<�wa<�va<Kua<bta<�sa<2sa<Nsa<�sa<�ta<!va<�wa<za<l|a<�~a<�a<K�a< �a<��a<�a<шa<{�a<��a<�a<�a<�a<�a<m�a<��a<F�a<N�a<#�a<z�a<��a<͐a<ܑa<Ғa<d�a<Гa<��a<#�a<��a<q�a<2�a<�a<m�a<Z�a<e�a<׊a<��a<��a<��a<׌a<Y�a<��a<�a<ēa<��a<�a<2�a<T�a<Йa<��a<�a<��a<+�a<��a<$�a<��a<j�a<)�a<i�a<Зa<D�a< �a<��a<U�a<ךa<8�a<7�a<�a<P�a<V�a<%�a<��a<�a<'�a<{�a<�a<�a<>�a<�a<�a<��a<��a<�a<f�a<�a<��a<�a<<�a<�a<ԙa<�a<˙a<\�a<ǘa<��a<>�a<s�a<ԕa<]�a<��a<�a<1�a<��a<�a<|�a<ޖa<�a<!�a<��a<a�a<9�a<�a<o�a<��a<��a<��a<��a<i�a<!�a<^�a<�a<�a<m�a<S�a<_�a<��a<�a<O�a<k�a<�a<��a<Ǐa<a�a<܎a<�a<�a<��a<��a<O�a<y�a<|�a<چa<��a<B�a<a�a<I�a<P�a<3�a< �a<p�a<��a<��a<�a<O�a<+~a<�{a<�ya<Jwa<Qua<}sa<ra<!qa<�pa<�pa<qa<�qa<�ra<ta<Aua<ava<\wa<�wa<{xa<oxa<xa<�wa<�va<�ua<�ta<�sa<�ra<kra<�qa<�qa<�qa<�qa<_ra<�ra<0sa<wsa<�sa<rsa<)sa<<ra<"qa<�oa<4na<xla<�ja<�ha<�ga<ufa<�ea<�ea<�ea<�fa<�ga<ia<�ja<�la<�  �  oa<�pa<ra<�ra<�sa<�sa<ta<�sa<Jsa<�ra<Qra<�qa<�qa<�qa<�qa<=ra<sa<ta<<ua<rva<�wa<�xa<�ya<za<Nza<Pza<�ya<ya<Axa<Twa<}va<�ua<ua<�ta<�ta<Tua<va<�wa<8ya<?{a<k}a<wa<��a<��a<k�a<��a<Շa<��a<��a<�a<��a<�a<Ɉa<��a<�a<;�a<׉a<͊a<Ջa<$�a<��a<ݏa<�a<L�a<�a<��a<��a<��a<�a<�a<ߐa<Џa<��a<��a<׌a<4�a<9�a<s�a<�a<B�a<��a<-�a<Œa<c�a<�a<p�a<��a<!�a<��a<��a<j�a<Ƙa<5�a<��a<Ԗa<B�a<�a<a<�a<g�a<��a<ėa<��a<c�a<3�a<��a<�a<ۚa<d�a<a<w�a<�a<��a<B�a<��a<c�a<]�a<��a<}�a<u�a<	�a<�a<�a<��a<Ҕa<*�a<k�a<��a<B�a<��a<��a<`�a<ǘa<ڗa<�a<�a<"�a<r�a<ؓa<��a<��a<ۓa<I�a<�a<��a<��a<��a<Öa<��a<*�a<z�a<j�a<ɒa<;�a<��a<�a<$�a<ˊa<��a<ǈa<~�a<Z�a<�a<��a<��a<��a<��a<ōa<��a<o�a<��a<��a<�a<Y�a<7�a<��a<��a<O�a<�a<��a<�a<k�a<%�a<�a<�a<@�a<`�a<q�a<{�a<"�a<��a<z�a<L�a<��a<�~a<�|a<�za<�xa<�va<�ta<vsa<�ra<ra<�qa<ora<�ra<�sa<�ta<�ua<�va<�wa<7xa<Ixa<.xa<�wa<wa<�ua<�ta<�sa<�ra<�qa<�pa<fpa<6pa<^pa<�pa<#qa<�qa<>ra<�ra<,sa<*sa<�ra<Pra<�qa<(pa<�na<2ma<�ka<0ja<�ha<�ga<4ga<+ga<=ga<�ga<ia<Kja<�ka<rma<�  �  	pa<9qa<Mra<sa<xsa<�sa<fsa<�ra<nra<�qa<�pa<dpa<pa<�oa<0pa<�pa<�qa<�ra<�sa<Oua<�va<�wa<�xa<�ya<Cza<~za<Aza<�ya<Jya<ixa<�wa<�va<eva<Eva<Vva<�va<�wa<ya<�za<�|a<v~a<��a<n�a<�a<��a<Ɔa<��a<�a<0�a<(�a<�a<��a<]�a<L�a<N�a<��a<E�a<0�a<j�a<��a<-�a<��a<@�a<y�a<��a<F�a<��a<̓a<Q�a<��a<�a<ِa<��a<�a<=�a<�a<ɍa<�a<Ǝa<��a<�a<l�a<ԓa<m�a<��a<��a<��a<�a<:�a<�a<��a<�a< �a<!�a<c�a<Ȕa<[�a<1�a<b�a<˔a<�a<\�a<c�a<��a<G�a<�a<��a<��a<��a<�a<�a<�a<Ėa<[�a<�a<˒a<�a<J�a<��a< �a<��a<X�a<l�a<��a<�a<-�a<�a<�a<g�a<y�a<F�a<��a<ڗa<��a<˕a<��a<��a<ڒa<Q�a<�a<�a<T�a<ؒa<��a<`�a<%�a<��a<.�a<J�a<�a<��a<��a<��a<C�a<��a<�a<��a<.�a<4�a<f�a<�a<�a<T�a<�a<�a<Ɍa<Ӎa<��a<?�a<��a<��a<I�a<��a<��a<W�a<�a<X�a<�a<��a<Z�a<|�a<كa<��a<��a<��a<��a<r�a<��a<��a<��a<4�a<��a<��a<�a<xa<�}a<�{a<�ya<�wa<Vva<4ua<;ta<�sa<�sa<�sa<[ta<5ua<�ua<�va<�wa<	xa<oxa<Fxa<�wa<7wa<va<ua<�sa<Zra<0qa<-pa<]oa<�na<�na<�na<(oa<�oa<}pa<`qa<�qa<wra<�ra<�ra<qra<�qa<�pa<�oa<Rna<�la<�ka<Nja<ria<�ha<�ha<�ha<�ia<fja<�ka<ma<�na<�  �  �pa<�qa<�ra<6sa<dsa<3sa<�ra<ra<Cqa<Gpa<�oa<�na<Sna<=na<Sna<oa<�oa<qa<�ra<�sa<�ua<wa<~xa<sya<>za<�za<�za<�za<za<�ya<�xa<�xa<xa<�wa<!xa<�xa<�ya<�za<T|a<�}a<�a<��a<1�a<˄a<�a<܆a<c�a<��a<��a<2�a<Æa<M�a<��a<��a<��a<�a<y�a<��a<��a<V�a<�a<��a<B�a<Ӑa<*�a<�a<Ǔa<��a<��a<��a<ߒa<�a<P�a<��a<��a<��a<��a<ԏa<r�a<M�a<��a<��a<�a<D�a<y�a<T�a<�a<"�a<��a<��a<Ǘa<ߖa<��a<Ӕa<�a<�a<��a<Y�a<��a<�a<�a<�a<�a<N�a<f�a<|�a<&�a<��a<��a<R�a<ԙa<Әa<̗a<��a<��a<|�a<��a<�a<��a<�a<A�a<�a<�a<ڕa<�a<�a<טa<D�a<��a<e�a<ߘa<*�a<�a<ӕa<n�a<U�a<�a<%�a<��a<*�a<Z�a<��a<X�a<3�a<�a<�a<�a<��a<��a<�a<Еa<5�a<X�a<�a<ȑa<_�a<'�a<ԍa<݌a<0�a<��a<ڋa<�a<��a<N�a<��a<Ύa<h�a<�a<�a<��a<�a<5�a<�a<a�a<��a<�a<��a<�a<��a<��a<�a<݁a<Ӂa<=�a<��a<�a<��a<�a<5�a<�a<��a<ła<��a<=�a<�~a<�|a<,{a<�ya<xa<�va<�ua<~ua<Yua<zua<va<~va<&wa<�wa<Zxa<�xa<�xa<Jxa<�wa<�va<bua< ta<ira<qa<�oa<pna<�ma<�la<�la<ma<�ma<fna<(oa<)pa<qa<�qa<ara<�ra<�ra<ra<�qa<ppa<Yoa<na<ma<�ka<ka<�ja<cja<�ja<(ka<la<9ma<Dna<�oa<�  �  �qa<�ra<sa<Hsa<Asa<�ra<ra<Hqa<,pa<oa<na<)ma<�la<qla<�la<<ma<*na<loa<qa<�ra<�ta<Jva<�wa<(ya<za<�za<,{a<0{a<�za<�za<Eza<�ya<�ya<�ya<�ya<gza<I{a<t|a<�}a<Da<	�a<��a<�a<I�a<'�a<Ԇa<;�a<	�a<Ɇa<V�a<��a<�a<R�a<�a<��a<�a<��a<҅a<�a<��a<��a<X�a<W�a<�a<��a<�a<��a</�a<w�a<0�a<�a<r�a<��a<�a<��a<X�a<O�a<��a<�a<��a<�a<�a<Q�a<5�a<�a<Øa<�a<�a<��a<�a<�a<��a<��a<f�a<5�a<]�a<�a<��a<Ґa<o�a<=�a<d�a<͔a<+�a<��a<��a<��a<l�a<��a<��a<X�a<��a<�a<�a<ߖa<��a<D�a<̔a<��a<��a<��a<��a<S�a<:�a<)�a<ǘa<c�a<��a<��a<B�a<|�a<m�a<;�a<��a<6�a<��a<p�a<�a<ǎa<q�a<��a<�a<��a<��a<Бa<	�a< �a<��a<��a<��a<�a<��a<�a<��a<�a<��a<~�a<v�a<��a<��a<��a<��a<a<�a<��a<\�a<ُa<#�a<j�a<+�a<��a<��a<��a<+�a<��a<��a<Æa<ׄa<;�a<�a<�a<S�a<*�a<"�a<��a<C�a<ہa<��a<;�a<��a<كa<��a<��a<3�a<�a<�a<;~a<x|a<{a<�ya<�xa<�wa<Dwa<wa<'wa<`wa<�wa<rxa<�xa<�xa<ya<�xa<0xa<[wa<	va<�ta<sa<:qa<�oa<na<�la<�ka<Gka<ka<gka<�ka<�la<�ma<oa<<pa<$qa<�qa<}ra<�ra<vra<ra<=qa<vpa<noa<_na<�ma<�la<ela<?la<mla<�la<�ma<�na<�oa<�pa<�  �  �ra<!sa<esa<asa<sa<�ra<cqa<Cpa<oa<�ma<�la<�ka<ka<�ja<ka<�ka<�la<na<�oa<�qa<vsa<Xua<+wa<�xa< za<�za<�{a<�{a<�{a<�{a<�{a<L{a<"{a<={a<r{a<�{a<�|a<�}a<6a<��a<�a<h�a<̈́a<΅a<}�a<ӆa<��a<��a<��a<J�a<��a<��a<�a<��a<A�a<��a<.�a<�a<��a<8�a<A�a<Q�a<J�a<9�a<$�a<��a<��a<��a<�a<�a<��a<k�a<��a<|�a<�a<�a<�a<+�a<��a<j�a<U�a<V�a<5�a<�a<Ԙa<,�a<K�a<�a<r�a<c�a<�a<Ȕa<��a<�a<ΐa<�a<+�a<�a<1�a<ȏa<ؐa<�a<��a<�a<��a<��a<g�a<A�a<��a<�a<�a<��a<a<�a<@�a<p�a<іa<P�a<�a<,�a<��a<�a<��a<r�a<�a<��a<�a<�a<��a<�a<;�a<��a<6�a<��a<�a<`�a<
�a<�a< �a<��a<یa<o�a<=�a<]�a<��a<�a<,�a<[�a<m�a<ەa<%�a< �a<��a<�a<�a<��a<�a<�a<,�a<��a<#�a<�a<5�a<��a<�a<j�a<��a<�a<�a<��a<��a<��a<F�a<^�a<z�a<|�a<}�a<s�a<؁a<N�a<Xa<�~a<m~a<�~a<a<�a<Ԁa<��a<g�a</�a<��a<��a<J�a<��a<��a<x�a<3a<�}a<r|a<-{a</za<Sya<�xa<�xa<�xa<�xa<ya<Vya<�ya<�ya<uya<ya<xa<wa<ua<�sa<�qa<-pa<Lna<�la<Oka<.ja<�ia<}ia<�ia<�ja<gka<�la<�ma<4oa<`pa<�qa<Qra<�ra<�ra<�ra<&ra<Oqa<�pa<�oa<�na<[na<�ma<�ma<�ma<sna<oa<�oa<�pa<�qa<�  �  sa<�sa<�sa<�sa<�ra<"ra<qa<�oa<Ena<�la<�ka<sja<�ia<jia<�ia<0ja<0ka<�la<�na<�pa<�ra<�ta<�va<zxa<�ya<7{a<�{a<g|a<�|a<�|a<�|a<�|a<n|a<�|a<�|a<b}a<[~a<9a<��a<��a<	�a<;�a<P�a<�a<��a<�a<��a<Z�a<��a<��a<��a<��a<Ła<#�a<ހa<�a<��a<��a<1�a<�a<�a<l�a<��a<Ȏa<ΐa<H�a<͓a<��a<<�a<��a<��a<Y�a<�a<Ҕa<e�a<q�a<O�a<��a<8�a<��a<��a<W�a<)�a<˘a<X�a<y�a<��a<�a<�a<�a<��a<�a<x�a<ېa<��a<p�a<Ӎa<��a<ˍa<_�a<|�a<�a<q�a<B�a<��a<��a<��a<�a<��a<>�a<Q�a<�a<��a<�a<f�a<Ęa<)�a<ؗa<��a<��a<�a<X�a<�a<h�a<�a<B�a<m�a<C�a<�a<�a<͗a<`�a<��a<Ԓa<�a<9�a<��a<w�a<��a<V�a<��a<��a<��a<'�a<��a<1�a<��a<
�a<�a<ϕa<`�a<K�a< �a<��a<ٔa<��a<)�a<7�a<��a<��a<��a<��a<��a<ܐa<�a<\�a<��a<��a<@�a<��a<�a<e�a<�a<�a<ֈa<��a<C�a<K�a<m�a<�~a<�}a<;}a<}a<P}a<�}a<�~a<�a<��a<��a<قa<6�a<��a<��a<��a<H�a<?�a<"�a<�~a<�}a<}|a<�{a<�za<Fza<za<�ya<za< za<Jza<Iza<9za<�ya<7ya<xa<�va<-ua<Bsa<5qa<$oa<ma<`ka<�ia<�ha<0ha<ha<Wha<&ia<Cja<�ka<ma<�na<pa<9qa<ra<�ra<	sa<sa<�ra<1ra<�qa<�pa<Epa<�oa<poa</oa<yoa<�oa<dpa<qa<�qa<�ra<�  �  �sa<ta<�sa<�sa<�ra<�qa<�pa<oa<�ma<�ka<�ja<�ia<�ha<qha<Zha<Iia<.ja<�ka<�ma<�oa<ra<;ta<Yva<Exa<�ya<*{a<,|a<�|a<}a<�}a<E}a<U}a<^}a<�}a<�}a<{~a<Xa<&�a<Z�a<n�a<�a<�a<҅a<��a<̆a<�a<��a<��a<�a<��a<ׂa<��a<��a<�a<�a<�a<��a<܁a< �a<B�a<<�a<��a<��a<7�a<_�a<4�a<��a<��a<��a<�a<-�a<@�a<��a<��a<T�a<a�a<h�a<��a<�a<��a<g�a<�a<�a<]�a<ԙa<֙a<t�a<�a<�a<��a<�a<j�a<��a<�a<��a<j�a<�a<d�a<̌a<s�a<��a<�a<��a<��a<Z�a<�a<��a<�a<�a<l�a<՛a<��a<q�a<ؚa<%�a<��a<�a<�a<��a<ʘa<јa<=�a<��a</�a<��a<ǚa<�a<��a<�a<ؘa<��a<�a<�a<�a<�a<d�a<Ȍa<~�a<Ɗa<.�a<��a<��a< �a<Z�a<̎a<��a<�a<��a<͔a<ŕa<S�a<��a<��a<�a<��a<��a<�a<'�a<~�a<�a<��a<��a<t�a<��a<Ƒa<9�a<;�a<
�a<��a<ѐa<֏a<S�a<��a<i�a<.�a<хa<p�a<�a<aa<~a<�|a<&|a<4|a<?|a<)}a<�}a<a<P�a<e�a<j�a<"�a<��a<��a<p�a<ǂa<�a<	�a<�a<�~a<l}a<�|a<�{a<Y{a<{a<�za<�za<�za<3{a<�za<�za<za<+ya<xa<�va<�ta<�ra<�pa<Mna<Fla<�ja<�ha<�ga<
ga<ga<lga<*ha<nia<�ja<_la<�ma<�oa<�pa<ra<�ra<7sa<�sa<4sa<�ra<[ra<�qa<%qa<�pa<�pa<Dpa<�pa<�pa<Iqa<�qa<�ra<_sa<�  �  �sa<5ta<	ta<�sa<�ra<�qa<Lpa<�na<ma<�ka<�ia<�ha<�ga<�ga<�ga<nha<{ia<*ka<ma<Zoa<�qa<ta<va<Dxa<�ya<A{a<N|a<}a<j}a<�}a<�}a<�}a<-~a<G~a<�~a<8a<�a<��a<�a<'�a<3�a<$�a< �a<��a<��a<׆a<��a<υa<ӄa<��a<f�a<B�a<5�a<na<a<Pa<�a<��a<y�a<z�a<��a<%�a<��a<	�a<.�a<6�a<��a<�a<ҕa<T�a<h�a<|�a<r�a<P�a<,�a<��a<$�a<e�a<˖a<y�a<�a<��a<6�a<��a<�a<��a<��a<͘a<�a<V�a<Ӕa<��a<9�a<y�a<��a<��a<�a<΋a<�a<��a<эa<X�a<0�a<�a<�a<ܖa<��a<�a<�a<��a<��a<�a<��a<E�a<Ԛa<c�a<ܙa<��a<X�a<b�a<��a<�a<U�a<��a<�a<#�a<�a<��a<�a<Θa<y�a<��a<a<��a<��a<��a<�a<��a<��a<��a<��a<B�a<c�a<��a<i�a<�a<בa<J�a<˔a<��a<j�a<��a<Жa<c�a<ݕa<M�a<��a<��a<6�a<��a<c�a</�a<H�a<g�a<�a<��a<m�a<X�a<ޑa<�a<��a<P�a<a�a<6�a<Շa<_�a<�a<��a<�~a<*}a< |a<{a<M{a<�{a<b|a<r}a<�~a<�a<6�a<9�a<#�a<y�a<��a<��a<�a<%�a<E�a<M�a<Ea<D~a<>}a<�|a<|a<�{a<�{a<�{a<|{a<W{a<%{a<�za<Bza<Qya<�wa<�va<rta<pra< pa<�ma<�ka<�ia<&ha<ga<tfa<Nfa<�fa<{ga<�ha<Kja<�ka<�ma<Goa<�pa<�qa<�ra<dsa<�sa<�sa<"sa<�ra<Sra<�qa<eqa<qa<qa<'qa<zqa<ra<�ra<sa<�sa<�  �  �sa<�sa<�sa<�ra<�qa<pa<na<la<�ia<nga<2ea<�ca<Uba<�aa<�aa<}ba<da<fa<�ha<ska<3na<gqa< ta<�va<�xa<�za<�{a<�|a<c}a<j}a<�}a<M}a<d}a<�}a<�}a<o~a<Fa<U�a<Q�a<Ԃa<�a<:�a<�a<��a<߆a<m�a<��a<J�a<Ȃa<�a<a<V}a<�{a<�za<�ya<�ya<}za<�{a<�}a<	�a<�a<�a<�a<6�a<�a<��a<z�a<)�a<�a<��a<��a<͖a<��a<�a<��a<�a<ӕa<�a<��a<6�a<ۗa<�a<v�a<'�a<E�a<�a<��a<k�a<�a<ٔa<Ӓa<-�a<�a<��a<m�a<�a<��a<m�a<��a<��a<'�a<�a<��a<��a<��a<�a<\�a<N�a<Ěa<Ûa<�a<I�a<�a<o�a<��a<��a<��a<�a<��a<��a<b�a<��a<!�a<ۚa<(�a<}�a<=�a<Ϛa<ƙa<<�a<D�a<ݓa<~�a<��a<�a<p�a<h�a<��a<��a<4�a<M�a<U�a<ņa<��a<��a<!�a<��a<��a<��a<4�a<g�a<ޖa<��a<Жa<�a<w�a<\�a<��a<	�a<M�a<�a<�a<
�a<�a<��a<��a<ܒa<��a<�a<-�a<��a<��a<�a<Y�a<W�a</�a<-a<?|a<�ya<�wa<�va<�ua<�ua<�va<�wa<lya<D{a<$}a<a<��a<�a<�a<��a<^�a<��a<;�a<�a<�a<�~a<�}a<�|a<�{a<1{a<{a<�za<�za<-{a<{a<{a<�za<�ya<�xa<wa<ua<nra<�oa<�la<ja<6ga<�da<�ba<-aa<�`a<X`a<�`a<Cba<�ca<fa<Bha<�ja<�la<oa<�pa<ra<�ra<8sa<Osa<�ra<\ra<�qa<�pa<�pa<pa<pa<'pa<�pa<qa<�qa<�ra<6sa<�  �  ysa<�sa<|sa<�ra<�qa<Epa<Pna<*la<�ia<�ga<pea<�ca<�ba<�aa<ba<�ba<:da<Cfa<�ha<�ka<tna<�qa<Zta<�va<�xa<�za<�{a<�|a<}a<K}a<P}a<D}a<8}a<F}a<�}a<'~a<�~a<�a<R�a<��a<ރa<�a<�a<��a<��a<e�a<��a<~�a<��a<1�a<Va<�}a<�{a<�za<2za< za<�za<|a<�}a<W�a<!�a<1�a<J�a<Z�a<"�a<��a<��a<�a<�a<��a<��a<��a<j�a<�a<a<��a<��a<ѕa<N�a<�a<ٗa<��a<X�a<�a<-�a<�a<��a<r�a<�a<,�a<��a<q�a<�a<��a<��a<�a<�a<��a<�a<ԇa<R�a<M�a<��a<D�a<�a<W�a<��a<V�a<��a<��a<�a<��a<��a<6�a<��a<�a<F�a<טa<��a<��a<��a<~�a<�a<��a<��a<.�a<%�a<��a<��a<G�a<z�a<*�a<��a<ݎa<B�a<��a<��a<�a<Մa<\�a<��a<�a<��a<шa< �a<b�a<܏a<�a<�a<;�a<@�a<Жa<ޖa<��a<�a<.�a<S�a<q�a<��a<�a<��a<��a<ɑa<�a<a�a<��a<��a<x�a<�a< �a<��a<��a<E�a<��a<��a<n�a<ca<�|a<za<;xa<�va<?va<Hva<�va<xa<�ya<s{a<X}a<9a<րa<-�a<�a<`�a<_�a<ւa<�a<�a<�a<�~a<W}a<F|a<y{a<�za<�za<�za<�za<�za<�za<�za<�za<�ya<�xa<wa<5ua<�ra<pa<
ma<5ja<\ga<�da<�ba<�aa<�`a<�`a<@aa<nba<da<Ifa<�ha<�ja<1ma<=oa<�pa< ra<�ra<$sa<sa<�ra<#ra<�qa<�pa<9pa<�oa<�oa<�oa<Npa<�pa<�qa<mra<sa<�  �  
sa<�sa<Msa<�ra<�qa<Zpa<�na<~la<qja<<ha<Pfa<�da<�ca<ca<�ba<�ca<ea<+ga<�ia<:la<oa<�qa<�ta<�va<ya<�za<�{a<o|a<�|a<�|a<}|a<|a<N|a<I|a<�|a<1}a<~a<a<��a<Ɂa<B�a<��a<��a<_�a<��a<��a<��a<��a<I�a<��a<�a<7~a<�|a<�{a<5{a<	{a<�{a<}a<�~a<@�a<փa<Άa<ωa<��a<Z�a<��a<��a<�a<ؕa<9�a<H�a<�a<��a<D�a<Ȕa<��a<��a<�a<V�a<�a<�a<ėa<�a<g�a<�a<�a<t�a<��a<'�a<`�a<:�a<�a<��a<w�a<��a<�a<�a<z�a<�a<ǈa<-�a<.�a<`�a<�a<A�a<��a<��a<j�a<a<k�a<ۛa<��a<Q�a<��a<ƙa<�a<L�a<�a<��a<ۗa<��a<��a<D�a<ҙa<��a<��a<�a<w�a<��a<^�a<��a<n�a<��a<��a<�a<��a<p�a<ֆa<ۅa<9�a<��a<^�a<�a<��a<ŋa<�a<#�a<:�a<��a<]�a<:�a<��a<��a<�a<��a<[�a<��a<��a<��a<5�a<Ȑa<a<͐a<<�a<��a<�a<6�a<�a<Бa<ِa<��a<��a<}�a<وa<��a<�a<�a<r}a<�za<>ya<�wa<#wa<Qwa<�wa<�xa<Qza<|a<�}a<�a<�a<6�a<�a<=�a<&�a<�a<��a<e�a<�~a<�}a<]|a<^{a<�za<za<�ya<�ya<za<za<{za<^za<=za<�ya<�xa<<wa<?ua<�ra<Opa<�ma<�ja<(ha<�ea<�ca<�ba<�aa<�aa<3ba<Ica< ea<�fa<1ia<Qka<yma<]oa<�pa<ra<�ra<�ra<�ra<Gra<lqa<�pa<�oa<?oa<oa<�na<oa<Ooa<pa<�pa<�qa<�ra<�  �  gra<�ra<�ra<�ra<�qa<�pa<1oa<Xma<Nka<Iia<zga<�ea<�da<dda<xda<7ea<|fa<fha<�ja<9ma<�oa<�ra<ua<Hwa<ya<�za<9{a<�{a<�{a<�{a<�{a<E{a<{a<{a<D{a<�{a<�|a<�}a<Ca<ǀa<I�a<��a<�a<̅a<S�a<p�a<�a<-�a<�a<x�a<�a<[a<~a<}a<||a<�|a<.}a<^~a<�a<b�a<��a<Ça<��a<a�a<ُa<ܑa<��a<��a<F�a<��a<o�a<�a<��a<	�a<�a<N�a<1�a<}�a<�a<ɔa<Օa<֖a<ܗa<��a<N�a<a�a<U�a<��a<r�a<�a<�a<�a<��a<��a<ˋa<N�a<l�a<�a<K�a<�a<}�a<T�a<v�a<Ƒa<�a<A�a<�a<��a<��a<�a<E�a<��a<[�a<��a<��a<Зa<�a<��a<J�a<l�a<��a<b�a<�a<ߘa<��a<�a<^�a<�a<��a<v�a<�a<�a<Ӓa<c�a<��a<��a<��a<'�a<;�a<Άa<�a<a<�a<ъa<Ōa<ގa<��a<ǒa<H�a<j�a<�a<"�a<�a<T�a<~�a<k�a<T�a<?�a<c�a<a<^�a<h�a<��a<��a<��a<��a<S�a<�a<<�a<��a<��a<�a<�a<��a<Άa<��a<1�a<�~a<R|a<�za<Nya<�xa<�xa<ya<za<v{a<}a<�~a<@�a<��a<l�a<�a<�a<��a<�a<��a<ga<�}a<|a<{a<za<ya<�xa<lxa<nxa<�xa<ya<uya<�ya<�ya<#ya<�xa<Bwa<�ua<~sa<qa<zna<�ka<Pia<ga<*ea<�ca<%ca<ca<�ca<�da<%fa<ha<ja<-la<na<�oa<qa<ra<Lra<ara<�qa<Rqa<upa<�oa<�na<�ma<�ma<ama<�ma<na<�na<�oa<�pa<�qa<�  �  �qa<Hra<�ra<�ra<ra<9qa<�oa<[na<tla<�ja<ia<�ga<�fa<3fa<qfa<�fa<nha<ja<7la<�na<qa<�sa<�ua<�wa<ya<Xza<�za<4{a<
{a<�za<+za<�ya<Vya<(ya<bya< za<�za<|a<�}a<8a<��a<��a<?�a<E�a<!�a<]�a<B�a<��a<��a<��a<%�a<�a<�a<�~a<N~a<y~a< a<'�a<	�a<
�a<��a<�a<��a<1�a<^�a<>�a<��a<��a<͔a<�a<n�a<ēa<�a<V�a<Ǒa<b�a<f�a<��a<+�a<�a<&�a<l�a<��a<��a<��a< �a<)�a<��a<ߗa<~�a<�a<��a<�a<)�a<{�a<B�a</�a<�a<'�a<��a<T�a<�a<��a<�a<(�a<��a<��a<��a<��a<ښa<��a<,�a<7�a<9�a<�a<�a<A�a<��a<��a<��a<�a<��a<�a<��a<i�a<I�a<��a<Йa<~�a<��a<o�a<��a<Փa<��a<n�a<D�a<��a<�a<
�a<Ȉa<̈a<��a<ъa<[�a<.�a<��a<�a<e�a<��a<l�a<��a<˕a<a�a<w�a<B�a<	�a<��a<��a<��a<�a<��a<z�a<ɍa<H�a<�a<��a<F�a<ːa<��a<o�a<��a<;�a<x�a<K�a<�a<<�a<a<7�a<3~a<W|a<<{a<�za<aza< {a<�{a<}a<S~a<�a<�a<�a<ςa<��a<�a<�a<7�a<�a<~a<l|a<�za<]ya<xa<Rwa<�va<�va<�va<wa<�wa<2xa<�xa<�xa<�xa<Xxa<6wa<�ua<ta<�qa<�oa<1ma<�ja<�ha<ga<�ea<ea<�da<eea<ofa<�ga<�ia<>ka<8ma<�na<Hpa<8qa<�qa<ra<�qa<3qa<.pa<'oa<�ma<ma<5la<�ka<�ka<�ka<Bla<"ma<$na<boa<xpa<�  �  fpa<xqa<6ra<�ra<Gra<�qa<�pa<joa<�ma<Yla<�ja<�ia<�ha<qha<�ha<?ia<wja<la<�ma<.pa<nra<�ta<uva<xa<Nya<'za<bza<Cza<�ya<Mya<rxa<�wa<_wa<wa<Cwa<�wa<�xa<za<�{a<m}a<�a<h�a<�a<��a<ƅa<h�a<��a<C�a<��a<̈́a<��a<��a<��a<Հa<��a<��a<?�a<j�a<��a<�a<3�a<��a<�a<3�a<��a<��a<��a<-�a<0�a<Փa<1�a<g�a<F�a<s�a<��a<<�a<3�a<�a<�a<"�a<T�a<��a<E�a<��a<��a<y�a<�a<��a</�a<,�a<�a<U�a<��a<�a<k�a<@�a<s�a<,�a<\�a< �a<B�a<��a<��a<^�a<C�a<՗a<�a<��a<x�a<n�a<��a<�a<��a<��a<F�a<,�a<0�a<��a<B�a<^�a<ݒa<��a<��a<�a<*�a<�a<�a<`�a<`�a<Әa<��a<��a<�a<��a<�a<�a<w�a<0�a<I�a<��a<�a<��a<��a<�a<��a<^�a<�a<�a<�a<��a<Ǖa<K�a<q�a<@�a<��a<P�a<�a<��a<k�a<��a<Y�a<Q�a<��a<b�a<&�a<=�a<
�a<��a<�a<�a<��a<}�a<
�a<G�a<"�a<��a<^�a<�a<#�a<�~a<a}a<�|a<�|a<�|a<�}a<�~a<�a<�a<�a<��a<�a<	�a<��a<�a<�a<w~a<�|a<�za<�xa<Pwa<�ua< ua<�ta<kta<�ta<Dua<�ua<�va<{wa<�wa<;xa<xa<_wa<Fva<�ta<sa<�pa<�na<�la<�ja<ia<�ga<Dga<ga<�ga<]ha<�ia<ka<�la<Sna<�oa<�pa<vqa<�qa<�qa<�pa<	pa<�na<�ma<0la<ka<%ja<�ia<Zia<�ia<0ja<1ka<Zla<�ma<9oa<�  �  7oa<�pa<�qa<Ira<tra<-ra<�qa<wpa<Xoa<na<�la<�ka<ka<�ja<�ja<�ka<�la</na<�oa<�qa<�sa<�ua<Pwa<�xa<kya<�ya<�ya<iya<�xa<�wa<�va<�ua<!ua<�ta<�ta<Tua<lva<�wa<�ya<�{a<�}a<�a<�a<��a<G�a<R�a<Ɔa<�a<��a<�a<6�a<V�a<��a<��a<҂a<��a<��a<��a<�a<�a<�a</�a<*�a<�a<��a<͒a<��a<��a<��a<ےa<Ցa<��a<��a<|�a<t�a<��a<a<�a<̍a<܎a<k�a<�a<��a<7�a<��a<ܗa<��a<֘a<��a<�a<�a<��a<@�a<ϒa<��a<c�a<ҏa<w�a<ďa<[�a<d�a<ْa<E�a<�a<W�a<��a<��a<0�a<N�a<�a<$�a<��a<��a<�a<u�a<�a<��a<5�a<Ώa<�a<��a<��a<ݒa<0�a<��a<�a<$�a<Θa<&�a< �a<c�a<p�a<�a<o�a<��a<&�a<��a<e�a<��a<9�a<m�a<�a<�a<�a<a�a<��a<�a<��a<��a<��a<i�a<��a<��a< �a<g�a<��a<��a<Z�a<*�a<c�a<�a<�a<p�a<d�a<a�a<��a<��a<��a<`�a<��a<x�a<��a<��a<.�a<>�a<M�a<,�a<;�a<H�a<ڀa<�a<a<�~a<a<�a<��a<r�a<8�a<��a<o�a<^�a<�a<�a<ۀa<"a<}a<{a<�xa<�va<
ua<�sa<�ra<:ra<,ra<�ra<[sa<5ta<Gua<-va<wa<�wa<�wa<vwa<�va<�ua<ta<=ra<apa<~na<�la<=ka<Ija<�ia<�ia<�ia<ja<�ka<�la<5na<goa<�pa<Mqa<�qa<�qa<qa<Apa<�na<yma<�ka<`ja<�ha<�ga<9ga<�fa<@ga<�ga<
ia<�ja<la<�ma<�  �  -na<�oa<(qa<"ra<�ra<�ra<`ra<�qa<�pa<�oa<�na<�ma<\ma<'ma<Rma<�ma<�na<Cpa<�qa<�sa<@ua<�va<xa<ya<�ya<�ya<7ya<�xa<}wa<,va<�ta<�sa<�ra<�ra<|ra<sa<ta<�ua<�wa<�ya<5|a<�~a<!�a<�a<�a<>�a<6�a<��a<��a<=�a<҆a<�a<��a<B�a<�a<i�a<	�a<��a<f�a<�a<ǋa<ҍa<��a<�a<]�a<?�a<��a<f�a<Ēa<�a<��a<�a<��a<X�a<P�a<��a<m�a<��a<��a<��a<F�a<)�a<�a<�a<ٕa<9�a<B�a<�a<�a<��a<��a<�a<�a<��a<��a<��a<�a<�a<�a<��a<��a<��a<�a<t�a<��a<��a<=�a<��a<.�a<q�a<E�a<ۖa<�a<H�a<x�a<�a<��a<؍a<��a<��a<_�a<j�a<Րa<��a<5�a<��a<<�a<R�a<��a<B�a<��a<;�a<&�a<�a<r�a<�a<Ƒa<��a< �a<��a<��a<5�a<��a<�a<�a<1�a<�a<��a<�a<�a<0�a< �a<��a<�a<Վa<ڌa<��a<7�a<�a<��a<��a<��a<L�a<@�a<z�a<�a<_�a<��a<��a<4�a<d�a<.�a<W�a<�a<��a<�a<�a<(�a<��a<�a<,�a<��a<2�a<]�a<��a<B�a<�a<��a<�a<�a<Ѓa< �a<āa<�a<0~a<�{a<gya<wa<�ta<�ra<fqa<Ypa<�oa<�oa<\pa<6qa<jra<�sa<ua<2va<�va<pwa<�wa<-wa<?va<ua<�sa<ra<Fpa<�na<�ma<�la<�ka<�ka<	la<�la<�ma<�na<�oa<�pa<nqa<�qa<ra<�qa<�pa<coa<�ma<la<7ja<dha<�fa<�ea<�da<�da<�da<�ea<�fa<|ha<]ja<Ela<�  �  "ma< oa<�pa<�qa<�ra<5sa<6sa<�ra<ra<hqa<�pa<�oa<ooa<Foa<�oa<pa<�pa<,ra<�sa<ua<~va<�wa<�xa<uya<�ya<Pya<�xa<�wa<[va<�ta<esa<�qa<qa<bpa<Mpa<�pa<�qa<�sa<�ua<xa<�za<m}a<�a<t�a<��a<�a<y�a<�a<��a<z�a<&�a<чa<l�a<>�a<1�a<��a<6�a<�a<l�a<�a<��a<)�a<a<*�a<�a<��a<x�a<!�a<$�a<�a<W�a<��a<�a<o�a<\�a<e�a<M�a<��a<Q�a<Ȋa<i�a<��a<��a<�a<�a<��a<�a<�a<t�a<d�a<�a<K�a<e�a<d�a<{�a<��a<:�a<+�a<<�a<��a<��a<��a<��a<��a<Ǚa<{�a<��a<��a<��a<�a<��a<ԕa<��a<��a<��a<��a<��a<��a<]�a<i�a<D�a<}�a<�a<�a<̒a<Քa<p�a<�a<Øa<e�a<j�a<�a<W�a<5�a<�a<̔a<��a<Œa< �a<��a<ܑa<D�a<�a<��a<��a<o�a<1�a<u�a<v�a<�a<�a<��a<Ǒa<ʏa<i�a<D�a<�a<J�a<��a<˄a<y�a<s�a<R�a<Q�a<Ǉa<c�a<�a<��a<�a<�a<D�a<q�a<��a<!�a<όa<=�a<��a<��a<��a<:�a<T�a<��a<U�a<d�a<��a<�a<l�a<фa<	�a<��a<"�a<�a<�a<sa<,}a<�za<�wa<cua<�ra<�pa<#oa<:na<�ma<�ma<mna<Yoa<�pa<=ra<�sa<<ua<mva<1wa<�wa<�wa<�va<1va<�ta<�sa<ra<�pa<�oa<�na<Bna<�ma<!na<�na<Uoa<?pa<	qa<�qa<Ura<cra<-ra<Nqa<Fpa<�na<�la<�ja<�ha<�fa<�da<�ca<�ba<wba<�ba<�ca<�da<�fa<�ha<�ja<�  �  %la<Zna<?pa<�qa<sa<~sa<�sa<�sa<Ssa<�ra<,ra<�qa<=qa<1qa<[qa<�qa<�ra<�sa<ua<ava<�wa<�xa<aya<�ya<�ya<ya</xa<�va<Kua<�sa<�qa<apa<6oa<�na<mna<�na<pa<�qa<�sa<�va<Tya<R|a<<a<�a<3�a<,�a<��a<��a<;�a<e�a<p�a<C�a<�a<�a<�a<g�a<�a<�a<!�a<��a<
�a<|�a<��a<גa<d�a<��a<��a<��a<��a<�a<=�a<I�a<o�a<ňa<q�a<��a<Y�a<��a<y�a<�a<ϊa<�a<i�a<ԑa<!�a<(�a<��a<�a<��a<�a<יa<]�a<��a<��a<0�a<�a<*�a<�a<#�a<��a<E�a<+�a<�a<��a<��a<"�a<�a<ךa<�a<��a<�a<ޔa<��a<L�a<&�a<@�a<��a<Ήa<d�a<��a<W�a<��a<z�a<{�a<��a<דa<˕a<h�a<��a<��a<��a<��a<+�a<k�a<p�a<l�a<q�a<��a<�a<��a<͓a<�a<��a<F�a<�a<��a<��a<�a<��a<�a<��a<�a<�a<��a<6�a<��a<p�a<p�a<��a<�a<��a<��a<b�a<��a<;�a<�a<�a<ǋa<W�a<��a<Q�a<��a<G�a<ʎa<��a<��a<�a<��a<;�a<�a<*�a<��a<?�a<�a<O�a<��a<��a<ʅa<��a<�a<R�a<��a<�a<�~a<W|a<�ya<�va<�sa<<qa<oa<\ma<Fla<�ka<�ka<�la<�ma<Coa<qa<�ra<zta<�ua<�va<�wa<�wa<�wa<�va<�ua<�ta<�sa<qra<Xqa<�pa<pa<�oa<�oa<^pa<�pa<�qa<Bra<�ra<�ra<�ra<Vra<Eqa<�oa<na<�ka<�ia<=ga<ea</ca<�aa<�`a<~`a<�`a<�aa<0ca<"ea<Uga<�ia<�  �  Lka<�ma<�oa<�qa<sa<�sa<sta<Yta<Pta<�sa<Vsa<�ra<�ra<�ra<�ra<bsa<ta<$ua<6va<Xwa<�xa<?ya<�ya<�ya<�ya<�xa<�wa<=va<qta<�ra<�pa<;oa<�ma<5ma<�la<[ma<�na<Cpa<�ra<\ua<Yxa<|{a<r~a<_�a<�a<)�a<ɇa<
�a<щa<-�a<s�a<1�a<Y�a<;�a<b�a<ڊa<w�a<V�a<n�a<Ԏa<��a<|�a<��a<o�a<�a<�a<��a<|�a<�a<R�a<h�a<P�a<J�a<��a<�a<U�a<̈́a<#�a<2�a<��a<��a<��a<~�a< �a<z�a<��a<��a<�a<�a<��a<r�a<E�a<��a<��a<p�a<ȗa<��a<U�a<��a<ԗa<��a<`�a<�a<��a<T�a<��a<��a<�a<ۙa<@�a<U�a<
�a<��a<F�a<��a<�a<V�a<w�a<͇a<B�a<�a<o�a<O�a<o�a<̐a<��a<1�a<
�a<��a<��a<�a<N�a<ԙa<g�a<`�a<��a<��a<וa<|�a<�a<7�a<P�a<ߕa<]�a<�a<}�a<��a<��a<��a<#�a<��a<��a<l�a<ߍa<U�a<��a<J�a<�a<��a<z�a<�a<^�a<��a<x�a<�a<�a<�a<��a<͌a<7�a<N�a<��a<Џa<a�a<��a<��a<�a<�a<��a<j�a<��a<��a<��a<e�a<��a<y�a<��a<��a<O�a<��a<{�a<�a<ڀa<k~a<�{a<�xa<�ua<�ra<pa<�ma<la<�ja<Fja<�ja<2ka<�la<!na<pa<�qa<�sa<uua<�va<�wa<�wa<xa<�wa<�va<�ua<�ta<�sa<�ra<�qa<kqa<Rqa<=qa<�qa</ra<�ra<Fsa<dsa<�sa<+sa<ora<5qa<yoa<sma<ka<�ha<7fa<�ca<�aa<N`a<}_a<�^a<w_a<W`a<�aa<�ca<Ifa<�ha<�  �  �ja<~ma<�oa<�qa<sa<ta<�ta<�ta<�ta<xta<ta<�sa<sa<zsa<�sa<8ta<�ta<�ua<wa<
xa<�xa<�ya<#za<$za<�ya<�xa<�wa<�ua<ta<ra<!pa<[na<ma<@la<la<~la<�ma<moa<�qa<�ta<�wa<�za<.~a<*�a<�a<�a<އa<@�a<�a<��a<�a<�a<#�a<-�a<U�a<��a<^�a<A�a<d�a<��a<ސa<��a<�a<ēa<,�a<�a<l�a<s�a<�a<�a<ތa<��a<��a<��a<2�a<J�a<�a<7�a<3�a<��a<ňa<:�a<ߍa<��a<'�a<��a<��a<��a<�a<��a<՚a<��a<P�a<ڙa<E�a<Øa<g�a<O�a<p�a<Әa<q�a<&�a<њa<i�a<̛a<��a<��a<�a<��a<3�a<�a<��a<�a<��a<"�a<�a<t�a<h�a<�a<8�a<�a<��a<p�a<ɍa<#�a<��a<�a<��a<z�a<��a<K�a<��a<G�a<ҙa<&�a<_�a<��a<֖a<U�a<�a<�a<H�a<��a<4�a<��a<�a<��a<Зa<&�a<�a<��a<��a<�a<�a<��a< �a<i�a<A�a<��a<��a<�a<R�a<!�a<��a<M�a<l�a<��a<��a<��a</�a<(�a<֏a<�a<��a<��a<�a<�a<��a<|�a<^�a<�a<܇a<{�a<\�a<Y�a<Z�a<A�a<�a<��a<�a<��a<�a<рa<3~a<O{a<&xa<ua<�qa<,oa<�la<	ka<�ia<Zia<�ia<Xja<�ka<{ma<xoa<�qa<�sa<Bua<�va<�wa<&xa<Fxa<�wa<Mwa<pva<�ua<�ta<�sa<�ra<era<-ra<<ra<�ra<�ra<[sa<�sa<�sa<�sa<\sa<qra<qa<loa<8ma<�ja<ha<�ea<ca<aa<k_a<o^a<
^a<m^a<n_a<aa<ca<�ea<4ha<�  �  �ja<0ma<�oa<�qa<-sa<8ta<�ta<ua<�ta<�ta<0ta<�sa<�sa<�sa<	ta<zta<Oua<va<)wa<>xa<%ya<�ya<4za<Oza<�ya<�xa<gwa<�ua<�sa<�qa<�oa<na<�la<�ka<�ka<Hla<Rma<Loa<�qa<ota<�wa<�za<~a<߀a<��a<��a<�a<B�a<6�a<�a<�a<Y�a<"�a<_�a<��a<��a<��a<��a<��a<��a<�a<)�a<A�a<ߓa<+�a<,�a<a�a<T�a<��a<�a<��a<��a<b�a<k�a<�a<�a<��a<�a<�a<��a<x�a< �a<��a<c�a<�a<M�a<w�a<�a<@�a<��a<	�a<�a<��a< �a<H�a<
�a<��a<��a<��a<9�a<��a<2�a<�a<��a<�a<�a<ƛa<�a<��a<��a<��a<��a<Ԑa<��a<�a<�a<F�a<�a<Ɇa<�a<ۇa<b�a<7�a<��a<��a<��a<��a<ǖa<q�a<��a<n�a<��a<��a<��a<o�a<q�a<��a<>�a<��a<c�a<O�a<��a<ǖa<Q�a<Ηa<�a<>�a<��a<R�a<�a<{�a<R�a<ۏa<N�a<f�a<Ǉa<�a<�a<X�a<8�a<�a<�a< �a<E�a<&�a<H�a<G�a<��a<N�a<�a<�a< �a<�a<ŏa<>�a<&�a<.�a<��a<��a<��a<��a<!�a<؇a<��a<R�a<��a<l�a<P�a<��a<�a<��a<ւa<��a<�}a<*{a<�wa<�ta<�qa<�na<�la<�ja<�ia<ia<Dia<6ja<hka<Ama<0oa<Yqa<Jsa<ua<�va<�wa<Uxa<Qxa<xa<}wa<�va<�ua<�ta<�sa<!sa<�ra<hra<�ra<�ra<sa<�sa<�sa<(ta<�sa<psa<�ra<qa<8oa<�la<�ja<�ga<qea<�ba<�`a<>_a<^a<�]a<^a<1_a<�`a<�ba<�ea<�ga<�  �  �ja<~ma<�oa<�qa<sa<ta<�ta<�ta<�ta<xta<ta<�sa<sa<zsa<�sa<8ta<�ta<�ua<wa<
xa<�xa<�ya<#za<$za<�ya<�xa<�wa<�ua<ta<ra<!pa<[na<ma<@la<la<~la<�ma<moa<�qa<�ta<�wa<�za<.~a<*�a<�a<�a<އa<@�a<�a<��a<�a<�a<#�a<-�a<U�a<��a<^�a<A�a<d�a<��a<ސa<��a<�a<ēa<,�a<�a<l�a<s�a<�a<�a<ތa<��a<��a<��a<2�a<J�a<�a<7�a<3�a<��a<ňa<:�a<ߍa<��a<'�a<��a<��a<��a<�a<��a<՚a<��a<P�a<ڙa<E�a<Øa<g�a<O�a<p�a<Әa<q�a<&�a<њa<i�a<̛a<��a<��a<�a<��a<3�a<�a<��a<�a<��a<"�a<�a<t�a<h�a<�a<8�a<�a<��a<p�a<ɍa<#�a<��a<�a<��a<z�a<��a<K�a<��a<G�a<ҙa<&�a<_�a<��a<֖a<U�a<�a<�a<H�a<��a<4�a<��a<�a<��a<Зa<&�a<�a<��a<��a<�a<�a<��a< �a<i�a<A�a<��a<��a<�a<R�a<!�a<��a<M�a<l�a<��a<��a<��a</�a<(�a<֏a<�a<��a<��a<�a<�a<��a<|�a<^�a<�a<܇a<{�a<\�a<Y�a<Z�a<A�a<�a<��a<�a<��a<�a<рa<3~a<O{a<&xa<ua<�qa<,oa<�la<	ka<�ia<Zia<�ia<Xja<�ka<{ma<xoa<�qa<�sa<Bua<�va<�wa<&xa<Fxa<�wa<Mwa<pva<�ua<�ta<�sa<�ra<era<-ra<<ra<�ra<�ra<[sa<�sa<�sa<�sa<\sa<qra<qa<loa<8ma<�ja<ha<�ea<ca<aa<k_a<o^a<
^a<m^a<n_a<aa<ca<�ea<4ha<�  �  Lka<�ma<�oa<�qa<sa<�sa<sta<Yta<Pta<�sa<Vsa<�ra<�ra<�ra<�ra<bsa<ta<$ua<6va<Xwa<�xa<?ya<�ya<�ya<�ya<�xa<�wa<=va<qta<�ra<�pa<;oa<�ma<5ma<�la<[ma<�na<Cpa<�ra<\ua<Yxa<|{a<r~a<_�a<�a<)�a<ɇa<
�a<щa<-�a<s�a<1�a<Y�a<;�a<b�a<ڊa<w�a<V�a<n�a<Ԏa<��a<|�a<��a<o�a<�a<�a<��a<|�a<�a<R�a<h�a<P�a<J�a<��a<�a<U�a<̈́a<#�a<2�a<��a<��a<��a<~�a< �a<z�a<��a<��a<�a<�a<��a<r�a<E�a<��a<��a<p�a<ȗa<��a<U�a<��a<ԗa<��a<`�a<�a<��a<T�a<��a<��a<�a<ۙa<@�a<U�a<
�a<��a<F�a<��a<�a<V�a<w�a<͇a<B�a<�a<o�a<O�a<o�a<̐a<��a<1�a<
�a<��a<��a<�a<N�a<ԙa<g�a<`�a<��a<��a<וa<|�a<�a<7�a<P�a<ߕa<]�a<�a<}�a<��a<��a<��a<#�a<��a<��a<l�a<ߍa<U�a<��a<J�a<�a<��a<z�a<�a<^�a<��a<x�a<�a<�a<�a<��a<͌a<7�a<N�a<��a<Џa<a�a<��a<��a<�a<�a<��a<j�a<��a<��a<��a<e�a<��a<y�a<��a<��a<O�a<��a<{�a<�a<ڀa<k~a<�{a<�xa<�ua<�ra<pa<�ma<la<�ja<Fja<�ja<2ka<�la<!na<pa<�qa<�sa<uua<�va<�wa<�wa<xa<�wa<�va<�ua<�ta<�sa<�ra<�qa<kqa<Rqa<=qa<�qa</ra<�ra<Fsa<dsa<�sa<+sa<ora<5qa<yoa<sma<ka<�ha<7fa<�ca<�aa<N`a<}_a<�^a<w_a<W`a<�aa<�ca<Ifa<�ha<�  �  %la<Zna<?pa<�qa<sa<~sa<�sa<�sa<Ssa<�ra<,ra<�qa<=qa<1qa<[qa<�qa<�ra<�sa<ua<ava<�wa<�xa<aya<�ya<�ya<ya</xa<�va<Kua<�sa<�qa<apa<6oa<�na<mna<�na<pa<�qa<�sa<�va<Tya<R|a<<a<�a<3�a<,�a<��a<��a<;�a<e�a<p�a<C�a<�a<�a<�a<g�a<�a<�a<!�a<��a<
�a<|�a<��a<גa<d�a<��a<��a<��a<��a<�a<=�a<I�a<o�a<ňa<q�a<��a<Y�a<��a<y�a<�a<ϊa<�a<i�a<ԑa<!�a<(�a<��a<�a<��a<�a<יa<]�a<��a<��a<0�a<�a<*�a<�a<#�a<��a<E�a<+�a<�a<��a<��a<"�a<�a<ךa<�a<��a<�a<ޔa<��a<L�a<&�a<@�a<��a<Ήa<d�a<��a<W�a<��a<z�a<{�a<��a<דa<˕a<h�a<��a<��a<��a<��a<+�a<k�a<p�a<l�a<q�a<��a<�a<��a<͓a<�a<��a<F�a<�a<��a<��a<�a<��a<�a<��a<�a<�a<��a<6�a<��a<p�a<p�a<��a<�a<��a<��a<b�a<��a<;�a<�a<�a<ǋa<W�a<��a<Q�a<��a<G�a<ʎa<��a<��a<�a<��a<;�a<�a<*�a<��a<?�a<�a<O�a<��a<��a<ʅa<��a<�a<R�a<��a<�a<�~a<W|a<�ya<�va<�sa<<qa<oa<\ma<Fla<�ka<�ka<�la<�ma<Coa<qa<�ra<zta<�ua<�va<�wa<�wa<�wa<�va<�ua<�ta<�sa<qra<Xqa<�pa<pa<�oa<�oa<^pa<�pa<�qa<Bra<�ra<�ra<�ra<Vra<Eqa<�oa<na<�ka<�ia<=ga<ea</ca<�aa<�`a<~`a<�`a<�aa<0ca<"ea<Uga<�ia<�  �  "ma< oa<�pa<�qa<�ra<5sa<6sa<�ra<ra<hqa<�pa<�oa<ooa<Foa<�oa<pa<�pa<,ra<�sa<ua<~va<�wa<�xa<uya<�ya<Pya<�xa<�wa<[va<�ta<esa<�qa<qa<bpa<Mpa<�pa<�qa<�sa<�ua<xa<�za<m}a<�a<t�a<��a<�a<y�a<�a<��a<z�a<&�a<чa<l�a<>�a<1�a<��a<6�a<�a<l�a<�a<��a<)�a<a<*�a<�a<��a<x�a<!�a<$�a<�a<W�a<��a<�a<o�a<\�a<e�a<M�a<��a<Q�a<Ȋa<i�a<��a<��a<�a<�a<��a<�a<�a<t�a<d�a<�a<K�a<e�a<d�a<{�a<��a<:�a<+�a<<�a<��a<��a<��a<��a<��a<Ǚa<{�a<��a<��a<��a<�a<��a<ԕa<��a<��a<��a<��a<��a<��a<]�a<i�a<D�a<}�a<�a<�a<̒a<Քa<p�a<�a<Øa<e�a<j�a<�a<W�a<5�a<�a<̔a<��a<Œa< �a<��a<ܑa<D�a<�a<��a<��a<o�a<1�a<u�a<v�a<�a<�a<��a<Ǒa<ʏa<i�a<D�a<�a<J�a<��a<˄a<y�a<s�a<R�a<Q�a<Ǉa<c�a<�a<��a<�a<�a<D�a<q�a<��a<!�a<όa<=�a<��a<��a<��a<:�a<T�a<��a<U�a<d�a<��a<�a<l�a<фa<	�a<��a<"�a<�a<�a<sa<,}a<�za<�wa<cua<�ra<�pa<#oa<:na<�ma<�ma<mna<Yoa<�pa<=ra<�sa<<ua<mva<1wa<�wa<�wa<�va<1va<�ta<�sa<ra<�pa<�oa<�na<Bna<�ma<!na<�na<Uoa<?pa<	qa<�qa<Ura<cra<-ra<Nqa<Fpa<�na<�la<�ja<�ha<�fa<�da<�ca<�ba<wba<�ba<�ca<�da<�fa<�ha<�ja<�  �  -na<�oa<(qa<"ra<�ra<�ra<`ra<�qa<�pa<�oa<�na<�ma<\ma<'ma<Rma<�ma<�na<Cpa<�qa<�sa<@ua<�va<xa<ya<�ya<�ya<7ya<�xa<}wa<,va<�ta<�sa<�ra<�ra<|ra<sa<ta<�ua<�wa<�ya<5|a<�~a<!�a<�a<�a<>�a<6�a<��a<��a<=�a<҆a<�a<��a<B�a<�a<i�a<	�a<��a<f�a<�a<ǋa<ҍa<��a<�a<]�a<?�a<��a<f�a<Ēa<�a<��a<�a<��a<X�a<P�a<��a<m�a<��a<��a<��a<F�a<)�a<�a<�a<ٕa<9�a<B�a<�a<�a<��a<��a<�a<�a<��a<��a<��a<�a<�a<�a<��a<��a<��a<�a<t�a<��a<��a<=�a<��a<.�a<q�a<E�a<ۖa<�a<H�a<x�a<�a<��a<؍a<��a<��a<_�a<j�a<Րa<��a<5�a<��a<<�a<R�a<��a<B�a<��a<;�a<&�a<�a<r�a<�a<Ƒa<��a< �a<��a<��a<5�a<��a<�a<�a<1�a<�a<��a<�a<�a<0�a< �a<��a<�a<Վa<ڌa<��a<7�a<�a<��a<��a<��a<L�a<@�a<z�a<�a<_�a<��a<��a<4�a<d�a<.�a<W�a<�a<��a<�a<�a<(�a<��a<�a<,�a<��a<2�a<]�a<��a<B�a<�a<��a<�a<�a<Ѓa< �a<āa<�a<0~a<�{a<gya<wa<�ta<�ra<fqa<Ypa<�oa<�oa<\pa<6qa<jra<�sa<ua<2va<�va<pwa<�wa<-wa<?va<ua<�sa<ra<Fpa<�na<�ma<�la<�ka<�ka<	la<�la<�ma<�na<�oa<�pa<nqa<�qa<ra<�qa<�pa<coa<�ma<la<7ja<dha<�fa<�ea<�da<�da<�da<�ea<�fa<|ha<]ja<Ela<�  �  7oa<�pa<�qa<Ira<tra<-ra<�qa<wpa<Xoa<na<�la<�ka<ka<�ja<�ja<�ka<�la</na<�oa<�qa<�sa<�ua<Pwa<�xa<kya<�ya<�ya<iya<�xa<�wa<�va<�ua<!ua<�ta<�ta<Tua<lva<�wa<�ya<�{a<�}a<�a<�a<��a<G�a<R�a<Ɔa<�a<��a<�a<6�a<V�a<��a<��a<҂a<��a<��a<��a<�a<�a<�a</�a<*�a<�a<��a<͒a<��a<��a<��a<ےa<Ցa<��a<��a<|�a<t�a<��a<a<�a<̍a<܎a<k�a<�a<��a<7�a<��a<ܗa<��a<֘a<��a<�a<�a<��a<@�a<ϒa<��a<c�a<ҏa<w�a<ďa<[�a<d�a<ْa<E�a<�a<W�a<��a<��a<0�a<N�a<�a<$�a<��a<��a<�a<u�a<�a<��a<5�a<Ώa<�a<��a<��a<ݒa<0�a<��a<�a<$�a<Θa<&�a< �a<c�a<p�a<�a<o�a<��a<&�a<��a<e�a<��a<9�a<m�a<�a<�a<�a<a�a<��a<�a<��a<��a<��a<i�a<��a<��a< �a<g�a<��a<��a<Z�a<*�a<c�a<�a<�a<p�a<d�a<a�a<��a<��a<��a<`�a<��a<x�a<��a<��a<.�a<>�a<M�a<,�a<;�a<H�a<ڀa<�a<a<�~a<a<�a<��a<r�a<8�a<��a<o�a<^�a<�a<�a<ۀa<"a<}a<{a<�xa<�va<
ua<�sa<�ra<:ra<,ra<�ra<[sa<5ta<Gua<-va<wa<�wa<�wa<vwa<�va<�ua<ta<=ra<apa<~na<�la<=ka<Ija<�ia<�ia<�ia<ja<�ka<�la<5na<goa<�pa<Mqa<�qa<�qa<qa<Apa<�na<yma<�ka<`ja<�ha<�ga<9ga<�fa<@ga<�ga<
ia<�ja<la<�ma<�  �  fpa<xqa<6ra<�ra<Gra<�qa<�pa<joa<�ma<Yla<�ja<�ia<�ha<qha<�ha<?ia<wja<la<�ma<.pa<nra<�ta<uva<xa<Nya<'za<bza<Cza<�ya<Mya<rxa<�wa<_wa<wa<Cwa<�wa<�xa<za<�{a<m}a<�a<h�a<�a<��a<ƅa<h�a<��a<C�a<��a<̈́a<��a<��a<��a<Հa<��a<��a<?�a<j�a<��a<�a<3�a<��a<�a<3�a<��a<��a<��a<-�a<0�a<Փa<1�a<g�a<F�a<s�a<��a<<�a<3�a<�a<�a<"�a<T�a<��a<E�a<��a<��a<y�a<�a<��a</�a<,�a<�a<U�a<��a<�a<k�a<@�a<s�a<,�a<\�a< �a<B�a<��a<��a<^�a<C�a<՗a<�a<��a<x�a<n�a<��a<�a<��a<��a<F�a<,�a<0�a<��a<B�a<^�a<ݒa<��a<��a<�a<*�a<�a<�a<`�a<`�a<Әa<��a<��a<�a<��a<�a<�a<w�a<0�a<I�a<��a<�a<��a<��a<�a<��a<^�a<�a<�a<�a<��a<Ǖa<K�a<q�a<@�a<��a<P�a<�a<��a<k�a<��a<Y�a<Q�a<��a<b�a<&�a<=�a<
�a<��a<�a<�a<��a<}�a<
�a<G�a<"�a<��a<^�a<�a<#�a<�~a<a}a<�|a<�|a<�|a<�}a<�~a<�a<�a<�a<��a<�a<	�a<��a<�a<�a<w~a<�|a<�za<�xa<Pwa<�ua< ua<�ta<kta<�ta<Dua<�ua<�va<{wa<�wa<;xa<xa<_wa<Fva<�ta<sa<�pa<�na<�la<�ja<ia<�ga<Dga<ga<�ga<]ha<�ia<ka<�la<Sna<�oa<�pa<vqa<�qa<�qa<�pa<	pa<�na<�ma<0la<ka<%ja<�ia<Zia<�ia<0ja<1ka<Zla<�ma<9oa<�  �  �qa<Hra<�ra<�ra<ra<9qa<�oa<[na<tla<�ja<ia<�ga<�fa<3fa<qfa<�fa<nha<ja<7la<�na<qa<�sa<�ua<�wa<ya<Xza<�za<4{a<
{a<�za<+za<�ya<Vya<(ya<bya< za<�za<|a<�}a<8a<��a<��a<?�a<E�a<!�a<]�a<B�a<��a<��a<��a<%�a<�a<�a<�~a<N~a<y~a< a<'�a<	�a<
�a<��a<�a<��a<1�a<^�a<>�a<��a<��a<͔a<�a<n�a<ēa<�a<V�a<Ǒa<b�a<f�a<��a<+�a<�a<&�a<l�a<��a<��a<��a< �a<)�a<��a<ߗa<~�a<�a<��a<�a<)�a<{�a<B�a</�a<�a<'�a<��a<T�a<�a<��a<�a<(�a<��a<��a<��a<��a<ښa<��a<,�a<7�a<9�a<�a<�a<A�a<��a<��a<��a<�a<��a<�a<��a<i�a<I�a<��a<Йa<~�a<��a<o�a<��a<Փa<��a<n�a<D�a<��a<�a<
�a<Ȉa<̈a<��a<ъa<[�a<.�a<��a<�a<e�a<��a<l�a<��a<˕a<a�a<w�a<B�a<	�a<��a<��a<��a<�a<��a<z�a<ɍa<H�a<�a<��a<F�a<ːa<��a<o�a<��a<;�a<x�a<K�a<�a<<�a<a<7�a<3~a<W|a<<{a<�za<aza< {a<�{a<}a<S~a<�a<�a<�a<ςa<��a<�a<�a<7�a<�a<~a<l|a<�za<]ya<xa<Rwa<�va<�va<�va<wa<�wa<2xa<�xa<�xa<�xa<Xxa<6wa<�ua<ta<�qa<�oa<1ma<�ja<�ha<ga<�ea<ea<�da<eea<ofa<�ga<�ia<>ka<8ma<�na<Hpa<8qa<�qa<ra<�qa<3qa<.pa<'oa<�ma<ma<5la<�ka<�ka<�ka<Bla<"ma<$na<boa<xpa<�  �  gra<�ra<�ra<�ra<�qa<�pa<1oa<Xma<Nka<Iia<zga<�ea<�da<dda<xda<7ea<|fa<fha<�ja<9ma<�oa<�ra<ua<Hwa<ya<�za<9{a<�{a<�{a<�{a<�{a<E{a<{a<{a<D{a<�{a<�|a<�}a<Ca<ǀa<I�a<��a<�a<̅a<S�a<p�a<�a<-�a<�a<x�a<�a<[a<~a<}a<||a<�|a<.}a<^~a<�a<b�a<��a<Ça<��a<a�a<ُa<ܑa<��a<��a<F�a<��a<o�a<�a<��a<	�a<�a<N�a<1�a<}�a<�a<ɔa<Օa<֖a<ܗa<��a<N�a<a�a<U�a<��a<r�a<�a<�a<�a<��a<��a<ˋa<N�a<l�a<�a<K�a<�a<}�a<T�a<v�a<Ƒa<�a<A�a<�a<��a<��a<�a<E�a<��a<[�a<��a<��a<Зa<�a<��a<J�a<l�a<��a<b�a<�a<ߘa<��a<�a<^�a<�a<��a<v�a<�a<�a<Ӓa<c�a<��a<��a<��a<'�a<;�a<Άa<�a<a<�a<ъa<Ōa<ގa<��a<ǒa<H�a<j�a<�a<"�a<�a<T�a<~�a<k�a<T�a<?�a<c�a<a<^�a<h�a<��a<��a<��a<��a<S�a<�a<<�a<��a<��a<�a<�a<��a<Άa<��a<1�a<�~a<R|a<�za<Nya<�xa<�xa<ya<za<v{a<}a<�~a<@�a<��a<l�a<�a<�a<��a<�a<��a<ga<�}a<|a<{a<za<ya<�xa<lxa<nxa<�xa<ya<uya<�ya<�ya<#ya<�xa<Bwa<�ua<~sa<qa<zna<�ka<Pia<ga<*ea<�ca<%ca<ca<�ca<�da<%fa<ha<ja<-la<na<�oa<qa<ra<Lra<ara<�qa<Rqa<upa<�oa<�na<�ma<�ma<ama<�ma<na<�na<�oa<�pa<�qa<�  �  
sa<�sa<Msa<�ra<�qa<Zpa<�na<~la<qja<<ha<Pfa<�da<�ca<ca<�ba<�ca<ea<+ga<�ia<:la<oa<�qa<�ta<�va<ya<�za<�{a<o|a<�|a<�|a<}|a<|a<N|a<I|a<�|a<1}a<~a<a<��a<Ɂa<B�a<��a<��a<_�a<��a<��a<��a<��a<I�a<��a<�a<7~a<�|a<�{a<5{a<	{a<�{a<}a<�~a<@�a<փa<Άa<ωa<��a<Z�a<��a<��a<�a<ؕa<9�a<H�a<�a<��a<D�a<Ȕa<��a<��a<�a<V�a<�a<�a<ėa<�a<g�a<�a<�a<t�a<��a<'�a<`�a<:�a<�a<��a<w�a<��a<�a<�a<z�a<�a<ǈa<-�a<.�a<`�a<�a<A�a<��a<��a<j�a<a<k�a<ۛa<��a<Q�a<��a<ƙa<�a<L�a<�a<��a<ۗa<��a<��a<D�a<ҙa<��a<��a<�a<w�a<��a<^�a<��a<n�a<��a<��a<�a<��a<p�a<ֆa<ۅa<9�a<��a<^�a<�a<��a<ŋa<�a<#�a<:�a<��a<]�a<:�a<��a<��a<�a<��a<[�a<��a<��a<��a<5�a<Ȑa<a<͐a<<�a<��a<�a<6�a<�a<Бa<ِa<��a<��a<}�a<وa<��a<�a<�a<r}a<�za<>ya<�wa<#wa<Qwa<�wa<�xa<Qza<|a<�}a<�a<�a<6�a<�a<=�a<&�a<�a<��a<e�a<�~a<�}a<]|a<^{a<�za<za<�ya<�ya<za<za<{za<^za<=za<�ya<�xa<<wa<?ua<�ra<Opa<�ma<�ja<(ha<�ea<�ca<�ba<�aa<�aa<3ba<Ica< ea<�fa<1ia<Qka<yma<]oa<�pa<ra<�ra<�ra<�ra<Gra<lqa<�pa<�oa<?oa<oa<�na<oa<Ooa<pa<�pa<�qa<�ra<�  �  ysa<�sa<|sa<�ra<�qa<Epa<Pna<*la<�ia<�ga<pea<�ca<�ba<�aa<ba<�ba<:da<Cfa<�ha<�ka<tna<�qa<Zta<�va<�xa<�za<�{a<�|a<}a<K}a<P}a<D}a<8}a<F}a<�}a<'~a<�~a<�a<R�a<��a<ރa<�a<�a<��a<��a<e�a<��a<~�a<��a<1�a<Va<�}a<�{a<�za<2za< za<�za<|a<�}a<W�a<!�a<1�a<J�a<Z�a<"�a<��a<��a<�a<�a<��a<��a<��a<j�a<�a<a<��a<��a<ѕa<N�a<�a<ٗa<��a<X�a<�a<-�a<�a<��a<r�a<�a<,�a<��a<q�a<�a<��a<��a<�a<�a<��a<�a<ԇa<R�a<M�a<��a<D�a<�a<W�a<��a<V�a<��a<��a<�a<��a<��a<6�a<��a<�a<F�a<טa<��a<��a<��a<~�a<�a<��a<��a<.�a<%�a<��a<��a<G�a<z�a<*�a<��a<ݎa<B�a<��a<��a<�a<Մa<\�a<��a<�a<��a<шa< �a<b�a<܏a<�a<�a<;�a<@�a<Жa<ޖa<��a<�a<.�a<S�a<q�a<��a<�a<��a<��a<ɑa<�a<a�a<��a<��a<x�a<�a< �a<��a<��a<E�a<��a<��a<n�a<ca<�|a<za<;xa<�va<?va<Hva<�va<xa<�ya<s{a<X}a<9a<րa<-�a<�a<`�a<_�a<ւa<�a<�a<�a<�~a<W}a<F|a<y{a<�za<�za<�za<�za<�za<�za<�za<�za<�ya<�xa<wa<5ua<�ra<pa<
ma<5ja<\ga<�da<�ba<�aa<�`a<�`a<@aa<nba<da<Ifa<�ha<�ja<1ma<=oa<�pa< ra<�ra<$sa<sa<�ra<#ra<�qa<�pa<9pa<�oa<�oa<�oa<Npa<�pa<�qa<mra<sa<�  �  �sa<�sa<�sa<sra<�pa<�na<�ka<	ia<�ea<�ba<�_a<P]a<�[a<�Za<�Za<�[a<`]a<�_a<Dca<�fa<�ja<�na<(ra<�ua<Wxa<vza<)|a<}a<n}a<w}a<q}a<5}a<}a<}a<(}a<�}a<�~a<�a<5�a<Ȃa<*�a<u�a<y�a<$�a<��a<>�a<�a<2�a<؀a<=~a<s{a<�xa<{va<�ta<�sa<Psa<�sa<tua<�wa<�za<�~a<t�a<��a<l�a<	�a<=�a<��a<��a<	�a<��a<��a<i�a<�a<z�a<�a<��a<a<�a<��a<]�a<>�a<?�a<�a<��a<�a<�a<�a<��a<u�a<��a<��a<]�a<�a<�a<��a<ҁa<Z�a<�a<�a<V�a<V�a<�a<_�a<��a<D�a<��a<��a<�a<ۚa<7�a<ٜa<Ӝa<d�a<ћa<�a<�a<��a<͘a<��a<��a<3�a<��a<y�a<)�a<��a<��a<�a<R�a<�a<	�a<��a<U�a<�a<h�a<��a<��a<��a<pa<	~a<�}a<�}a<'a<+�a<�a<��a<.�a<r�a<L�a<!�a<#�a<��a<��a<��a<S�a<��a<ƕa<��a<��a<ܒa<�a<ۑa<��a<�a<\�a<�a<?�a<w�a<`�a<�a<��a<��a<L�a<4�a<��a<��a<�~a<�za<wa<�sa<�qa<pa<Xoa<�oa<�pa<dra<�ta<rwa<Aza<�|a<aa<k�a<��a<��a<�a<R�a<p�a<5�a<�a<h~a<(}a<�{a<!{a<�za<dza<tza<�za<�za<{a<'{a<�za<za<�xa<�va<ta<�pa<9ma<jia<�ea<ba<�^a<\a<CZa<OYa<JYa<0Za<�[a<X^a<Waa<bda<�ga<�ja<�ma<�oa<�qa<�ra<Zsa<>sa<�ra<"ra<Tqa<kpa<�oa<2oa<9oa<8oa<�oa<�pa<�qa<hra<sa<�  �  �sa<�sa<bsa<vra<�pa<�na<Bla<<ia<	fa<�ba<`a<�]a<\a<,[a<[a<\a<�]a<f`a<}ca<)ga<�ja<�na<�ra<�ua<Zxa<rza<�{a<�|a<Y}a<j}a<}a<�|a<z|a<�|a<�|a<^}a<2~a<ea<րa<r�a<��a<o�a<N�a<��a<ۆa<P�a<�a<Q�a<
�a<k~a<�{a<ya<�va<ua<ta<�sa<qta<�ua<Dxa<K{a<�~a<��a<��a<��a<5�a<-�a<a<��a<Ŗa<]�a<��a<A�a<��a<%�a<��a<J�a<L�a<��a<�a<͖a<�a<�a<��a<��a<ޚa<��a<ߙa<�a<n�a<�a<ߐa<��a<G�a<�a<n�a<B�a<׀a<A�a<��a<ˁa<΃a<q�a<��a<�a<t�a<ȓa<��a<	�a<�a<�a<��a<��a<b�a<��a<��a<��a<��a<o�a<J�a<J�a<��a<<�a<�a<ܚa<��a<ޛa<��a<�a<�a<�a<��a<��a<B�a<��a<$�a<ބa<�a<�a<�~a<�}a<d~a<�a<��a< �a<3�a<h�a<��a<��a<"�a<%�a<��a<S�a<|�a<>�a<��a<m�a<X�a<*�a<U�a<��a<h�a<M�a<��a<��a<��a<�a<q�a<5�a<��a<x�a<��a<?�a<S�a<͆a<�a<�~a<	{a<�wa<tta<ra<�pa<�oa<pa<qa<�ra<ua<�wa<qza<#}a<�a<Z�a<˂a<v�a<��a<)�a<g�a<�a<�a<~a<�|a<{{a<�za<za<�ya<�ya<Eza<�za<{a<{a<�za<�ya<�xa<�va<�sa<�pa<gma<�ia<�ea<5ba<$_a<�\a<�Za<�Ya<�Ya<�Za<W\a<�^a<�aa<�da<�ga<ka<�ma<�oa<�qa<�ra<&sa<sa<�ra<�qa<�pa<�oa<Poa<�na<�na<�na<aoa<pa<*qa<ra<sa<�  �  �ra<esa<$sa<wra<qa<oa<�la<�ia<�fa<�ca<!aa<�^a<"]a<[\a<K\a<@]a<�^a<�aa<�da<"ha<�ka<_oa<�ra<�ua<xxa<fza<�{a<u|a<�|a<�|a<|a<�{a<�{a<u{a<�{a<|a<}a<T~a<�a<w�a<�a<��a<��a<��a<��a<d�a<3�a<��a<��a<a<�|a<za<�wa<9va<,ua<�ta<�ua<wa<\ya<\|a<�a<��a<r�a<'�a<��a<]�a<ғa<m�a<v�a<Ԗa<Ӗa<Z�a<��a<+�a<��a<9�a<�a<b�a<�a<ϕa<��a<�a<�a<�a<o�a<d�a<ϙa<��a<��a<\�a<g�a<c�a<C�a<�a<��a<X�a<�a<q�a<́a<�a<�a<{�a<~�a<ލa<	�a<A�a<��a</�a<�a<כa<V�a<�a<��a<��a<��a<��a<�a<Z�a<��a<6�a<��a<B�a<$�a<�a<Кa<3�a<j�a<��a<�a<+�a<Օa<�a<Џa<��a<�a<�a<0�a<��a<�a<%a<�a<��a<��a<#�a<,�a<=�a<*�a<�a<P�a<D�a<~�a<�a<�a<��a<��a<q�a<k�a<0�a<I�a<��a<$�a<8�a<x�a<�a<��a<�a<��a<��a<X�a<T�a<ӏa<n�a<��a<V�a<��a<�a<�{a<�xa<�ua<1sa<�qa<�pa<&qa<*ra<�sa<va<�xa<3{a<�}a<�a<��a<܂a<Z�a<O�a<��a<��a<&�a<�~a<}a<�{a<kza<rya<�xa<�xa<�xa<Yya<�ya<$za<Wza<<za<�ya<sxa<�va<#ta<dqa<�ma<pja<�fa<;ca<?`a<�]a<�[a<�Za<�Za<�[a<r]a<�_a<vba<�ea<�ha<�ka<na<pa<�qa<ura<�ra<zra<�qa<�pa<pa<oa<=na<�ma<qma<�ma<Rna<!oa<0pa< qa<Ira<�  �  ra<�ra<�ra<Cra<Eqa<�oa<Xma<�ja<ha<Vea<�ba<�`a< _a<S^a<U^a<4_a<�`a<-ca<)fa<via<�la<\pa<|sa<kva<�xa<)za<?{a<�{a<�{a<Y{a<�za<.za<�ya<�ya<�ya<1za<{a<�|a<~a<�a<݁a<��a<��a<�a<k�a<<�a<��a<.�a<Z�a<)�a<�}a<�{a<�ya<xa<*wa<�va<�wa<ya<B{a<�}a<j�a<ڄa<{�a<��a<�a<ّa<��a<*�a<��a<�a<a</�a<V�a<`�a<Œa<;�a<#�a<g�a<�a<�a<6�a<��a<�a<�a<��a<�a<��a<��a<*�a<ޔa<X�a<s�a<��a<Éa<*�a<J�a<��a<s�a<ǃa<�a<��a<�a<�a<��a<�a<�a<��a<v�a<��a<y�a<��a<<�a<m�a<^�a<'�a<�a<�a<W�a<�a<0�a<��a<}�a<��a<��a<��a<V�a<a<��a<��a<`�a<i�a<��a<֐a<��a<��a<��a<��a<��a<��a<0�a<��a<��a<f�a<͆a<��a<P�a<'�a<��a<�a<Z�a<B�a<��a<g�a<��a<z�a</�a<��a<u�a<e�a<��a<;�a<8�a<��a<=�a<"�a<�a<��a<�a<͑a<�a<��a<ڍa</�a<�a<��a<
�a<�}a</za<jwa<0ua<�sa<sa<&sa<ta<}ua<�wa<�ya<<|a<�~a<l�a<�a<��a<�a<ӂa<�a<��a<�~a</}a<N{a<�ya<mxa<�wa<�va<�va<,wa<�wa<Uxa<�xa<Yya<�ya<(ya<3xa<�va<�ta<�qa<�na<ka<ha<�da<�aa<�_a<�]a<�\a<�\a<�]a<?_a<Vaa<�ca<�fa<�ia<2la<�na<\pa<yqa<ra<4ra<�qa<�pa<�oa<tna<Ama<gla<�ka<�ka<�ka<wla<\ma<�na<�oa<qa<�  �  �pa<�qa<Xra</ra<eqa<)pa<?na<?la<�ia<>ga<�da<�ba<�aa<�`a<�`a<�aa<Tca<nea<@ha<Ika<ina<�qa<Kta<�va<�xa<za<�za<�za<qza<�ya<ya<xa<�wa<wa<&wa<�wa<�xa<?za<�{a<~a<�a<�a<�a<�a<"�a<1�a<�a<Ԅa<g�a<��a<za<�}a<�{a<|za<�ya<wya<za<s{a<�}a<+�a<f�a<��a<��a<�a<ďa<7�a<��a<�a<�a<�a<b�a<k�a<h�a<?�a<��a<��a<��a<�a<��a<ӑa<�a<ʔa<1�a<��a<��a<B�a<_�a<��a<��a<��a<��a<��a<S�a<Ћa<f�a<��a<c�a<��a<?�a<Y�a<�a<9�a<�a<��a<��a<��a<�a<��a<��a<�a<��a<�a<ݘa<��a<�a<��a<��a<Ԓa<��a<��a<Y�a<F�a<w�a<ޖa<�a<,�a<��a<�a<��a<��a<�a<��a<E�a<6�a<u�a<��a<E�a<u�a<!�a<��a<�a<�a<��a<�a<U�a<׍a<~�a<q�a<a�a<g�a<�a<	�a<]�a<V�a<֒a<[�a<��a<5�a<�a<�a<ًa<��a<c�a<�a<&�a<,�a<�a<͐a<�a<��a<��a<'�a<Ջa<)�a<%�a<��a<�a<Z|a<�ya<�wa<-va<�ua<�ua<}va<�wa<�ya<�{a<�}a<�a<�a<e�a<��a<ւa<�a<Հa<+a<8}a<A{a<-ya<�wa<�ua<ua<�ta<hta<�ta<tua<~va<=wa<xa<xxa<xxa<xa<�va</ua<�ra<'pa<ma<�ia<�fa<da<	ba<J`a<�_a<m_a<1`a<�aa<vca<�ea<Hha<ka<$ma<#oa<�pa<jqa<�qa<9qa<�pa<9oa<�ma<kla<ka<ja<;ia<2ia<Bia<ja<&ka<�la<na<~oa<�  �  �oa<�pa<�qa<ra<�qa<�pa<_oa<�ma<xka<aia<Uga<�ea<ada<�ca<�ca<�da<fa<%ha<�ja<ema<)pa<�ra<_ua<twa<�xa<�ya<�ya<�ya<�xa<�wa<�va<�ua<�ta<Jta<9ta<�ta<�ua<lwa<|ya<�{a<~a<m�a<��a<E�a<��a<?�a<F�a<ƅa<��a<!�a<��a<�a<X~a<5}a<z|a<w|a<}a<d~a<f�a<҂a<��a<��a<��a<H�a<��a<��a<֓a<v�a<F�a<ܓa<��a<n�a<�a<Ԏa<��a<��a<��a<�a<͍a<�a<��a<�a<M�a< �a<��a<y�a<�a<�a<�a<��a<ٔa<��a<n�a<�a<�a<x�a<`�a<�a<8�a<)�a<a<Ía<�a<��a<�a<�a<ݘa<�a<��a<x�a<Йa<a<)�a<w�a<ɓa<,�a<�a<��a<��a<͏a<��a<��a<�a<��a<L�a<ɗa<ɘa<^�a<r�a<ۘa<��a<ƕa<��a<�a<��a<�a<��a<=�a<�a<��a<�a<އa<_�a<=�a<q�a<��a<��a<��a<�a<��a<Օa<C�a<Y�a<ݒa< �a<�a<9�a<��a<�a<+�a<��a<�a<��a<��a<ߋa<*�a<n�a<��a<
�a<;�a<��a<��a<ǌa<O�a<��a<ńa<��a<�~a<�|a<za<-ya<�xa<}xa<4ya<Wza<�{a<�}a<Ha<Ҁa<�a<Âa<��a<d�a< �a<�a<�}a<;{a<�xa<�va<�ta<+sa<
ra<�qa<�qa<+ra<sa<3ta<Yua<�va<ewa<�wa<�wa<�va<�ua<�sa<`qa<�na<la<6ia<�fa<�da<Gca<�ba<fba<ca<Jda< fa<ha<?ja<^la<Dna<�oa<�pa<Sqa<qa<Spa</oa<�ma<�ka<ja<}ha<@ga<efa<fa<efa<Hga<�ha<-ja<�ka<�ma<�  �  �ma<�oa<�pa<�qa<�qa<�qa<�pa<%oa<�ma<�ka<�ia<lha<hga<�fa<�fa<�ga<ia<�ja<#ma<�oa<ra<rta<�va<�wa<	ya<`ya<2ya<�xa<Fwa<va<]ta<sa<�qa<Cqa<+qa<�qa<�ra<Yta<�va<%ya<|a<�~a<8�a<q�a<�a<>�a<��a<��a<��a<߄a<��a<4�a<
�a<�a<�a<�a<D�a<��a<1�a<��a<�a<֊a<K�a<��a<��a<��a<ߓa<�a<��a<u�a<��a<r�a<��a<�a<��a<��a<��a<�a<Ǌa<�a<��a<�a<m�a<j�a<S�a<Ǘa<��a<�a<��a<ʗa<T�a<��a<��a<��a<�a<[�a<��a<�a<o�a<=�a<��a<c�a<f�a<��a<��a<X�a<��a<E�a<j�a<֙a<�a<6�a<X�a<B�a<+�a<O�a<Ѝa<��a<w�a<Ōa<{�a<Ďa<}�a<m�a<v�a<1�a<̗a<��a<:�a<�a<I�a<�a<,�a<1�a<��a<��a<��a<E�a<U�a<ىa<+�a<͊a<#�a<ɍa<��a<��a<@�a<��a<s�a<וa<z�a<��a<)�a<-�a<$�a<��a<��a<��a<�a<�a<��a<�a<|�a<чa<E�a<�a<��a<�a<6�a<��a<��a<ێa<��a<��a<^�a<�a<"�a<��a<Qa<�}a<[|a<�{a<�{a<�{a<}a<A~a<�a<�a<=�a<�a<(�a<�a<сa<\�a<B~a<�{a<?ya<hva<�sa<�qa<)pa<�na<zna<�na<(oa<bpa<�qa<ysa<�ta< va<�va<@wa<wa<va<�ta<�ra<�pa<@na<�ka<�ia<�ga<�fa<�ea<�ea<fa<ga<�ha<]ja<`la<na<�oa<�pa<+qa<*qa<upa<eoa<�ma<�ka<�ia<{ga<�ea<*da<`ca<�ba<^ca<5da<�ea<�ga<�ia<�ka<�  �  Tla<�na<bpa<�qa<6ra<.ra<�qa<�pa<hoa<�ma<�la<Xka<zja< ja<ja<�ja<la<�ma<�oa<�qa<�sa<�ua<vwa<�xa<(ya<ya<xxa<$wa<�ua<�sa<
ra<apa<oa<*na<�ma<{na<�oa<~qa<�sa<�va<�ya<�|a<�a<d�a<��a<)�a<�a<P�a<B�a<��a<��a<��a<��a<�a<��a<��a<Z�a<��a<>�a<O�a<��a<Ȍa<�a<�a<h�a<��a<ғa<z�a<��a<�a<,�a<>�a<�a<M�a<Їa<a<k�a<��a<��a<I�a<R�a<��a<C�a<��a<�a<��a<I�a<�a<0�a<��a<Зa<V�a<ǔa<6�a<��a<q�a<��a<<�a<}�a<H�a<��a<�a<a<��a<2�a<{�a<;�a<��a<>�a<K�a<��a<��a<Y�a<��a<��a<��a<܊a<��a<[�a<��a<y�a<��a<�a<&�a<d�a<��a<��a<�a<�a<R�a<�a<�a<̖a<
�a<,�a<\�a<��a<W�a<`�a<��a<.�a<�a<��a<e�a<�a<^�a<Ŕa<��a<�a<��a<5�a<ܓa<̑a<��a<�a<`�a<�a<��a<��a<�a<��a<��a<��a<�a<Ća<߈a<Ɗa<��a<(�a<.�a<��a<W�a<P�a<�a<�a<ֈa<��a<a�a<X�a<��a<ka<�~a<�~a<a<�a<ʀa<Ɓa<тa<��a<a<��a<܂a<h�a<fa<�|a<�ya<wa<�sa<<qa<�na<�la<�ka<Ika<yka<ala<�ma<_oa<Oqa<sa<�ta<1va<�va< wa<�va<�ua<Uta<_ra<Zpa<Vna<ila<�ja<�ia<�ha<�ha<ia<	ja<Jka<�la<:na<�oa<�pa<Nqa<|qa<�pa<�oa<.na<la<�ia<Rga<�da<�ba<7aa<#`a<�_a<$`a<4aa<�ba<�da<iga<�ia<�  �  ka<ima<�oa<Bqa<lra<�ra<�ra<-ra<&qa<&pa<�na<�ma<Cma<�la<7ma<�ma<�na<Ipa<ra<�sa<�ua<Dwa<Vxa<4ya<7ya<�xa<�wa<va<;ta<�qa<�oa<�ma<Xla<Tka<�ja<zka<�la<�na<3qa<jta<�wa<!{a<�~a<[�a<$�a<�a<s�a<�a<Z�a< �a<��a<��a<"�a<Ʌa<l�a<��a<d�a<\�a<�a<��a<֌a<��a<��a<7�a<8�a<�a<��a<�a<��a<׏a<��a<!�a<�a<��a<�a<̓a<j�a<��a<Äa<��a<��a<��a<5�a<?�a<͓a<�a<�a<	�a<��a<��a<�a<�a<͖a<�a</�a<C�a<k�a<Y�a<f�a<�a</�a<f�a<�a<S�a<��a<z�a<��a<ۚa<�a<��a<��a<l�a<��a<ߎa<:�a<։a<�a<��a<X�a<��a<��a<H�a<v�a<�a<��a<U�a<l�a<n�a<��a<��a<��a<�a<5�a<Ȗa<_�a<��a<N�a<!�a<A�a<�a<�a<��a<��a<��a<��a<�a<�a<�a<��a<�a<ؔa<�a<��a<"�a<�a<;�a<U�a<�a<(�a<�a<�a<�a<�a<X�a<��a<a<!�a<p�a<�a<��a<W�a<��a<�a<�a<��a<��a<�a<Ća<�a<q�a<h�a<ˁa<v�a<ځa<<�a<�a<��a<i�a<a<��a<�a<��a<�a<c~a<�{a<_xa<�ta<�qa<�na<&la< ja<�ha<Kha<�ha<�ia<ka<;ma<Aoa<�qa<�sa<Hua<�va<wa<Gwa<�va<�ua<ta<_ra<�pa<�na<�ma<Pla<�ka<�ka<�ka<�la<�ma<�na<	pa<"qa<�qa<ra<�qa<�pa<Poa<ma<�ja<�ga<4ea<�ba<*`a<u^a<(]a<�\a<(]a<p^a<+`a<�ba<Gea<ha<�  �  �ia<�la<3oa<(qa<�ra<]sa<�sa<Zsa<�ra<�qa<�pa</pa<�oa<eoa<�oa<)pa<=qa<{ra<ta<�ua<*wa<exa<Mya<�ya<Dya<�xa<wa<ua<�ra<Ipa<�ma<�ka<�ia<�ha<�ha<�ha<=ja<Ula<�na<`ra<�ua<�ya<M}a<��a<��a<�a<��a<وa<l�a<s�a<A�a<Ԉa<E�a<�a<�a<)�a<шa<ىa<Q�a<֌a<��a<��a< �a<G�a<�a<+�a<��a<��a<Ԑa<��a<�a<i�a<�a<k�a<��a<e�a<�a<=�a<X�a<.�a<��a<��a<��a<ďa<Ȓa<s�a<��a<�a<	�a<p�a<'�a<��a<��a<��a<]�a<��a<�a<��a<�a<��a<k�a<��a<Ԙa<�a<�a<��a<��a<��a<��a<4�a<��a<�a<�a<�a<!�a<��a<��a<U�a<σa<!�a<9�a<��a<Z�a<�a<��a<�a<��a<�a<��a<��a<!�a<�a<b�a<a�a<0�a<ȕa<��a<��a<ƒa<s�a<��a<�a<��a<��a<��a<��a<5�a<v�a<�a<�a<��a<u�a<��a<��a<j�a<N�a<4�a<��a<�~a<u}a<�|a<U}a<v~a<�a<�a<��a<��a<2�a<`�a<J�a<S�a<�a<ُa<-�a<�a<y�a<a<�a<`�a<�a<ބa<8�a<�a<�a<[�a<��a<��a<a<҅a<j�a<Z�a<��a<��a<�}a<yza<�va<7sa<�oa<Zla<�ia<�ga<Ifa<�ea<+fa<Fga<�ha<Eka<�ma<.pa<�ra<�ta<Lva<'wa<�wa<uwa<�va<�ua<(ta<�ra<qa<�oa<�na<>na<na<bna<�na<�oa<�pa<�qa<Zra<�ra<�ra<�qa<�pa<�na<Cla<}ia<dfa<[ca<s`a<�]a<�[a<�Za<OZa<�Za<�[a<�]a<k`a<cca<xfa<�  �  �ha<�ka<�na<�pa<�ra<�sa<Yta<=ta<�sa</sa<�ra<�qa<�qa<iqa<xqa<*ra<sa<=ta<�ua<�va<Qxa<5ya<�ya<�ya<tya<2xa<�va<Wta<�qa<(oa<gla<ja</ha<�fa<�fa<�fa<Dha<dja<\ma<�pa<�ta<�xa<b|a<�a<�a<�a<�a<N�a<"�a<t�a<s�a<*�a<	�a<ǉa<މa<"�a<Ċa<ԋa<�a<��a<�a<��a<
�a<��a<��a<k�a<��a<,�a<Z�a<͍a<�a<9�a<?�a<ςa<��a<ga<�~a<=a<Y�a<U�a<�a<��a<r�a<��a<�a<�a<F�a<@�a<Z�a<�a<�a<��a<a<��a<#�a<`�a<�a<��a<�a<n�a<*�a<7�a<�a<*�a<Лa<5�a<�a<3�a<a<��a<+�a<�a<�a<��a<y�a<܅a<��a<`�a<Áa<)�a<<�a<=�a<��a<��a<�a<�a<�a<X�a<i�a<әa<��a<a<E�a<��a<h�a<m�a<J�a<l�a<̔a<X�a<��a<ݔa<{�a<E�a<�a<×a<�a<�a<c�a<D�a<O�a<�a< �a<��a<I�a<��a<��a<�~a<�|a<y{a<�za<]{a<�|a<�~a<րa<��a<��a<G�a<�a<��a<W�a<#�a<M�a<�a<�a<��a<�a<��a<�a<�a<؆a<+�a<�a<߅a<%�a<_�a<��a<͆a<��a<�a<��a<Âa<�a<5}a<�ya<�ua<ra<na<�ja<�ga<�ea<Dda<�ca<-da<lea<Uga<�ia<~la<oa<�qa<$ta<�ua<Swa<�wa<xa<uwa<�va<Sua<ta<�ra<�qa<�pa<$pa<pa<Cpa<�pa<rqa<	ra<�ra<Isa<ysa<sa<ra<�pa<>na<�ka<~ha<Rea<ba<�^a<0\a<Za<�Xa<CXa<�Xa<�Ya<!\a<�^a<�aa<cea<�  �  ha<yka<_na<�pa<�ra<ta<�ta<�ta<�ta<*ta<�sa<�ra<�ra<ra<�ra<@sa<"ta<4ua<�va<�wa<ya<�ya<9za<za<hya<
xa<3va<�sa<qa<:na<uka<ia<ga<�ea<Yea<�ea<ga<Nia<Bla<�oa<�sa<�wa<�{a<�a<��a<ׅa<��a<��a<��a<8�a<R�a<(�a<��a<Ŋa<�a<I�a<��a<�a<�a<��a<�a<��a<֓a<��a<֔a<��a<��a<��a<�a<A�a<G�a<@�a<>�a<��a<�a<D~a<�}a<~a<;a<9�a<�a<�a<��a<�a<��a<��a<�a</�a<��a<P�a<��a<i�a<��a<��a<�a<q�a<��a<�a<�a<{�a<#�a<'�a<�a<�a<��a<��a<8�a<<�a<��a<i�a<��a<��a<�a<��a<u�a<a<��a<0�a<��a<��a<&�a<%�a<��a<��a<�a<[�a<{�a<�a<D�a<יa<ǚa<�a<�a<j�a<c�a<d�a<D�a<y�a<�a<��a<��a<�a<s�a<?�a<�a<��a<��a<c�a<��a<8�a<&�a<��a<��a<�a<\�a<˃a<��a<�}a<�{a<Jza<�ya<2za<p{a<f}a<�a<Ăa<ąa<��a<u�a<��a<D�a<5�a<��a<W�a<��a<��a<�a<��a<�a<�a<��a<^�a<��a<�a<�a<^�a<��a<��a<�a<0�a<��a<��a<�a<�|a<ya<ua<qa<ma<�ia<�fa<xda<ca<�ba<ca<Qda<Ifa<�ha<�ka<una<Pqa<�sa<�ua<Awa<xa<Txa<xa<qwa<Eva<ua<�sa<�ra<�qa<oqa<1qa<Qqa<�qa<bra<sa<�sa<�sa<�sa<Ksa<$ra<bpa<
na<@ka<�ga<yda<
aa<�]a<[a<�Xa<�Wa<Wa<�Wa<�Xa<
[a<�]a<aa<�da<�  �  �ga<!ka<Qna<�pa<�ra<8ta<�ta<ua<�ta<xta<�sa<fsa<"sa<�ra<>sa<�sa<�ta<�ua<�va<xa<ya<�ya<rza<>za<^ya<xa<va<�sa<�pa<�ma<Ika<�ha<�fa<Uea<�da<Cea<�fa<�ha<�ka<�oa<vsa<�wa<�{a<ga<�a<ׅa<�a<Չa<��a<H�a<i�a<w�a<R�a<V�a<k�a<��a<k�a<^�a<��a<�a<l�a<��a<�a<��a<�a<��a<��a<�a<��a<�a<�a< �a<�a<N�a<4a<�}a<;}a<�}a<�~a<a<��a<Նa<7�a<ߍa<L�a<z�a<(�a<�a<��a<��a<��a<n�a<�a<P�a<��a<��a<b�a<^�a<f�a<�a<��a<��a<f�a<
�a<��a<��a<o�a<=�a<��a<f�a<b�a<T�a<ڍa<}�a<8�a<O�a< �a<��a<#�a<z�a<��a<��a<e�a<��a<Ìa<&�a<#�a<�a<C�a<ҙa<��a<E�a<�a<k�a<��a<��a<��a<�a<;�a<�a<��a<}�a<��a<��a<+�a<��a<ǘa<��a<��a<.�a<4�a<��a<D�a<Ԋa<�a<��a<4�a<J}a<({a<�ya<Kya<�ya<{a<�|a<�a<��a<��a<��a<*�a<��a<D�a<D�a<Րa<|�a<Əa<��a<e�a<�a<��a<p�a<n�a<҇a<x�a<p�a<r�a<��a<��a<��a<2�a<r�a<Ǆa<��a<�a<�|a<�xa<�ta<�pa<�la<>ia<Bfa<�ca<�ba<%ba<�ba<�ca<�ea<�ha<Bka<Hna<qa<�sa<�ua<0wa<.xa<�xa<1xa<vwa<�va<nua<0ta<Fsa<Era<�qa<�qa<�qa<.ra<�ra<[sa<�sa<ta<ta<�sa<$ra<_pa<na<�ja<�ga<:da<�`a<�]a<�Za<}Xa<Wa<�Va<Wa<nXa<�Za<v]a<�`a<?da<�  �  ha<yka<_na<�pa<�ra<ta<�ta<�ta<�ta<*ta<�sa<�ra<�ra<ra<�ra<@sa<"ta<4ua<�va<�wa<ya<�ya<9za<za<hya<
xa<3va<�sa<qa<:na<uka<ia<ga<�ea<Yea<�ea<ga<Nia<Bla<�oa<�sa<�wa<�{a<�a<��a<ׅa<��a<��a<��a<8�a<R�a<(�a<��a<Ŋa<�a<I�a<��a<�a<�a<��a<�a<��a<֓a<��a<֔a<��a<��a<��a<�a<A�a<G�a<@�a<>�a<��a<�a<D~a<�}a<~a<;a<9�a<�a<�a<��a<�a<��a<��a<�a</�a<��a<P�a<��a<i�a<��a<��a<�a<q�a<��a<�a<�a<{�a<#�a<'�a<�a<�a<��a<��a<8�a<<�a<��a<i�a<��a<��a<�a<��a<u�a<a<��a<0�a<��a<��a<&�a<%�a<��a<��a<�a<[�a<{�a<�a<D�a<יa<ǚa<�a<�a<j�a<c�a<d�a<D�a<y�a<�a<��a<��a<�a<s�a<?�a<�a<��a<��a<c�a<��a<8�a<&�a<��a<��a<�a<\�a<˃a<��a<�}a<�{a<Jza<�ya<2za<p{a<f}a<�a<Ăa<ąa<��a<u�a<��a<D�a<5�a<��a<W�a<��a<��a<�a<��a<�a<�a<��a<^�a<��a<�a<�a<^�a<��a<��a<�a<0�a<��a<��a<�a<�|a<ya<ua<qa<ma<�ia<�fa<xda<ca<�ba<ca<Qda<Ifa<�ha<�ka<una<Pqa<�sa<�ua<Awa<xa<Txa<xa<qwa<Eva<ua<�sa<�ra<�qa<oqa<1qa<Qqa<�qa<bra<sa<�sa<�sa<�sa<Ksa<$ra<bpa<
na<@ka<�ga<yda<
aa<�]a<[a<�Xa<�Wa<Wa<�Wa<�Xa<
[a<�]a<aa<�da<�  �  �ha<�ka<�na<�pa<�ra<�sa<Yta<=ta<�sa</sa<�ra<�qa<�qa<iqa<xqa<*ra<sa<=ta<�ua<�va<Qxa<5ya<�ya<�ya<tya<2xa<�va<Wta<�qa<(oa<gla<ja</ha<�fa<�fa<�fa<Dha<dja<\ma<�pa<�ta<�xa<b|a<�a<�a<�a<�a<N�a<"�a<t�a<s�a<*�a<	�a<ǉa<މa<"�a<Ċa<ԋa<�a<��a<�a<��a<
�a<��a<��a<k�a<��a<,�a<Z�a<͍a<�a<9�a<?�a<ςa<��a<ga<�~a<=a<Y�a<U�a<�a<��a<r�a<��a<�a<�a<F�a<@�a<Z�a<�a<�a<��a<a<��a<#�a<`�a<�a<��a<�a<n�a<*�a<7�a<�a<*�a<Лa<5�a<�a<3�a<a<��a<+�a<�a<�a<��a<y�a<܅a<��a<`�a<Áa<)�a<<�a<=�a<��a<��a<�a<�a<�a<X�a<i�a<әa<��a<a<E�a<��a<h�a<m�a<J�a<l�a<̔a<X�a<��a<ݔa<{�a<E�a<�a<×a<�a<�a<c�a<D�a<O�a<�a< �a<��a<I�a<��a<��a<�~a<�|a<y{a<�za<]{a<�|a<�~a<րa<��a<��a<G�a<�a<��a<W�a<#�a<M�a<�a<�a<��a<�a<��a<�a<�a<؆a<+�a<�a<߅a<%�a<_�a<��a<͆a<��a<�a<��a<Âa<�a<5}a<�ya<�ua<ra<na<�ja<�ga<�ea<Dda<�ca<-da<lea<Uga<�ia<~la<oa<�qa<$ta<�ua<Swa<�wa<xa<uwa<�va<Sua<ta<�ra<�qa<�pa<$pa<pa<Cpa<�pa<rqa<	ra<�ra<Isa<ysa<sa<ra<�pa<>na<�ka<~ha<Rea<ba<�^a<0\a<Za<�Xa<CXa<�Xa<�Ya<!\a<�^a<�aa<cea<�  �  �ia<�la<3oa<(qa<�ra<]sa<�sa<Zsa<�ra<�qa<�pa</pa<�oa<eoa<�oa<)pa<=qa<{ra<ta<�ua<*wa<exa<Mya<�ya<Dya<�xa<wa<ua<�ra<Ipa<�ma<�ka<�ia<�ha<�ha<�ha<=ja<Ula<�na<`ra<�ua<�ya<M}a<��a<��a<�a<��a<وa<l�a<s�a<A�a<Ԉa<E�a<�a<�a<)�a<шa<ىa<Q�a<֌a<��a<��a< �a<G�a<�a<+�a<��a<��a<Ԑa<��a<�a<i�a<�a<k�a<��a<e�a<�a<=�a<X�a<.�a<��a<��a<��a<ďa<Ȓa<s�a<��a<�a<	�a<p�a<'�a<��a<��a<��a<]�a<��a<�a<��a<�a<��a<k�a<��a<Ԙa<�a<�a<��a<��a<��a<��a<4�a<��a<�a<�a<�a<!�a<��a<��a<U�a<σa<!�a<9�a<��a<Z�a<�a<��a<�a<��a<�a<��a<��a<!�a<�a<b�a<a�a<0�a<ȕa<��a<��a<ƒa<s�a<��a<�a<��a<��a<��a<��a<5�a<v�a<�a<�a<��a<u�a<��a<��a<j�a<N�a<4�a<��a<�~a<u}a<�|a<U}a<v~a<�a<�a<��a<��a<2�a<`�a<J�a<S�a<�a<ُa<-�a<�a<y�a<a<�a<`�a<�a<ބa<8�a<�a<�a<[�a<��a<��a<a<҅a<j�a<Z�a<��a<��a<�}a<yza<�va<7sa<�oa<Zla<�ia<�ga<Ifa<�ea<+fa<Fga<�ha<Eka<�ma<.pa<�ra<�ta<Lva<'wa<�wa<uwa<�va<�ua<(ta<�ra<qa<�oa<�na<>na<na<bna<�na<�oa<�pa<�qa<Zra<�ra<�ra<�qa<�pa<�na<Cla<}ia<dfa<[ca<s`a<�]a<�[a<�Za<OZa<�Za<�[a<�]a<k`a<cca<xfa<�  �  ka<ima<�oa<Bqa<lra<�ra<�ra<-ra<&qa<&pa<�na<�ma<Cma<�la<7ma<�ma<�na<Ipa<ra<�sa<�ua<Dwa<Vxa<4ya<7ya<�xa<�wa<va<;ta<�qa<�oa<�ma<Xla<Tka<�ja<zka<�la<�na<3qa<jta<�wa<!{a<�~a<[�a<$�a<�a<s�a<�a<Z�a< �a<��a<��a<"�a<Ʌa<l�a<��a<d�a<\�a<�a<��a<֌a<��a<��a<7�a<8�a<�a<��a<�a<��a<׏a<��a<!�a<�a<��a<�a<̓a<j�a<��a<Äa<��a<��a<��a<5�a<?�a<͓a<�a<�a<	�a<��a<��a<�a<�a<͖a<�a</�a<C�a<k�a<Y�a<f�a<�a</�a<f�a<�a<S�a<��a<z�a<��a<ۚa<�a<��a<��a<l�a<��a<ߎa<:�a<։a<�a<��a<X�a<��a<��a<H�a<v�a<�a<��a<U�a<l�a<n�a<��a<��a<��a<�a<5�a<Ȗa<_�a<��a<N�a<!�a<A�a<�a<�a<��a<��a<��a<��a<�a<�a<�a<��a<�a<ؔa<�a<��a<"�a<�a<;�a<U�a<�a<(�a<�a<�a<�a<�a<X�a<��a<a<!�a<p�a<�a<��a<W�a<��a<�a<�a<��a<��a<�a<Ća<�a<q�a<h�a<ˁa<v�a<ځa<<�a<�a<��a<i�a<a<��a<�a<��a<�a<c~a<�{a<_xa<�ta<�qa<�na<&la< ja<�ha<Kha<�ha<�ia<ka<;ma<Aoa<�qa<�sa<Hua<�va<wa<Gwa<�va<�ua<ta<_ra<�pa<�na<�ma<Pla<�ka<�ka<�ka<�la<�ma<�na<	pa<"qa<�qa<ra<�qa<�pa<Poa<ma<�ja<�ga<4ea<�ba<*`a<u^a<(]a<�\a<(]a<p^a<+`a<�ba<Gea<ha<�  �  Tla<�na<bpa<�qa<6ra<.ra<�qa<�pa<hoa<�ma<�la<Xka<zja< ja<ja<�ja<la<�ma<�oa<�qa<�sa<�ua<vwa<�xa<(ya<ya<xxa<$wa<�ua<�sa<
ra<apa<oa<*na<�ma<{na<�oa<~qa<�sa<�va<�ya<�|a<�a<d�a<��a<)�a<�a<P�a<B�a<��a<��a<��a<��a<�a<��a<��a<Z�a<��a<>�a<O�a<��a<Ȍa<�a<�a<h�a<��a<ғa<z�a<��a<�a<,�a<>�a<�a<M�a<Їa<a<k�a<��a<��a<I�a<R�a<��a<C�a<��a<�a<��a<I�a<�a<0�a<��a<Зa<V�a<ǔa<6�a<��a<q�a<��a<<�a<}�a<H�a<��a<�a<a<��a<2�a<{�a<;�a<��a<>�a<K�a<��a<��a<Y�a<��a<��a<��a<܊a<��a<[�a<��a<y�a<��a<�a<&�a<d�a<��a<��a<�a<�a<R�a<�a<�a<̖a<
�a<,�a<\�a<��a<W�a<`�a<��a<.�a<�a<��a<e�a<�a<^�a<Ŕa<��a<�a<��a<5�a<ܓa<̑a<��a<�a<`�a<�a<��a<��a<�a<��a<��a<��a<�a<Ća<߈a<Ɗa<��a<(�a<.�a<��a<W�a<P�a<�a<�a<ֈa<��a<a�a<X�a<��a<ka<�~a<�~a<a<�a<ʀa<Ɓa<тa<��a<a<��a<܂a<h�a<fa<�|a<�ya<wa<�sa<<qa<�na<�la<�ka<Ika<yka<ala<�ma<_oa<Oqa<sa<�ta<1va<�va< wa<�va<�ua<Uta<_ra<Zpa<Vna<ila<�ja<�ia<�ha<�ha<ia<	ja<Jka<�la<:na<�oa<�pa<Nqa<|qa<�pa<�oa<.na<la<�ia<Rga<�da<�ba<7aa<#`a<�_a<$`a<4aa<�ba<�da<iga<�ia<�  �  �ma<�oa<�pa<�qa<�qa<�qa<�pa<%oa<�ma<�ka<�ia<lha<hga<�fa<�fa<�ga<ia<�ja<#ma<�oa<ra<rta<�va<�wa<	ya<`ya<2ya<�xa<Fwa<va<]ta<sa<�qa<Cqa<+qa<�qa<�ra<Yta<�va<%ya<|a<�~a<8�a<q�a<�a<>�a<��a<��a<��a<߄a<��a<4�a<
�a<�a<�a<�a<D�a<��a<1�a<��a<�a<֊a<K�a<��a<��a<��a<ߓa<�a<��a<u�a<��a<r�a<��a<�a<��a<��a<��a<�a<Ǌa<�a<��a<�a<m�a<j�a<S�a<Ǘa<��a<�a<��a<ʗa<T�a<��a<��a<��a<�a<[�a<��a<�a<o�a<=�a<��a<c�a<f�a<��a<��a<X�a<��a<E�a<j�a<֙a<�a<6�a<X�a<B�a<+�a<O�a<Ѝa<��a<w�a<Ōa<{�a<Ďa<}�a<m�a<v�a<1�a<̗a<��a<:�a<�a<I�a<�a<,�a<1�a<��a<��a<��a<E�a<U�a<ىa<+�a<͊a<#�a<ɍa<��a<��a<@�a<��a<s�a<וa<z�a<��a<)�a<-�a<$�a<��a<��a<��a<�a<�a<��a<�a<|�a<чa<E�a<�a<��a<�a<6�a<��a<��a<ێa<��a<��a<^�a<�a<"�a<��a<Qa<�}a<[|a<�{a<�{a<�{a<}a<A~a<�a<�a<=�a<�a<(�a<�a<сa<\�a<B~a<�{a<?ya<hva<�sa<�qa<)pa<�na<zna<�na<(oa<bpa<�qa<ysa<�ta< va<�va<@wa<wa<va<�ta<�ra<�pa<@na<�ka<�ia<�ga<�fa<�ea<�ea<fa<ga<�ha<]ja<`la<na<�oa<�pa<+qa<*qa<upa<eoa<�ma<�ka<�ia<{ga<�ea<*da<`ca<�ba<^ca<5da<�ea<�ga<�ia<�ka<�  �  �oa<�pa<�qa<ra<�qa<�pa<_oa<�ma<xka<aia<Uga<�ea<ada<�ca<�ca<�da<fa<%ha<�ja<ema<)pa<�ra<_ua<twa<�xa<�ya<�ya<�ya<�xa<�wa<�va<�ua<�ta<Jta<9ta<�ta<�ua<lwa<|ya<�{a<~a<m�a<��a<E�a<��a<?�a<F�a<ƅa<��a<!�a<��a<�a<X~a<5}a<z|a<w|a<}a<d~a<f�a<҂a<��a<��a<��a<H�a<��a<��a<֓a<v�a<F�a<ܓa<��a<n�a<�a<Ԏa<��a<��a<��a<�a<͍a<�a<��a<�a<M�a< �a<��a<y�a<�a<�a<�a<��a<ٔa<��a<n�a<�a<�a<x�a<`�a<�a<8�a<)�a<a<Ía<�a<��a<�a<�a<ݘa<�a<��a<x�a<Йa<a<)�a<w�a<ɓa<,�a<�a<��a<��a<͏a<��a<��a<�a<��a<L�a<ɗa<ɘa<^�a<r�a<ۘa<��a<ƕa<��a<�a<��a<�a<��a<=�a<�a<��a<�a<އa<_�a<=�a<q�a<��a<��a<��a<�a<��a<Օa<C�a<Y�a<ݒa< �a<�a<9�a<��a<�a<+�a<��a<�a<��a<��a<ߋa<*�a<n�a<��a<
�a<;�a<��a<��a<ǌa<O�a<��a<ńa<��a<�~a<�|a<za<-ya<�xa<}xa<4ya<Wza<�{a<�}a<Ha<Ҁa<�a<Âa<��a<d�a< �a<�a<�}a<;{a<�xa<�va<�ta<+sa<
ra<�qa<�qa<+ra<sa<3ta<Yua<�va<ewa<�wa<�wa<�va<�ua<�sa<`qa<�na<la<6ia<�fa<�da<Gca<�ba<fba<ca<Jda< fa<ha<?ja<^la<Dna<�oa<�pa<Sqa<qa<Spa</oa<�ma<�ka<ja<}ha<@ga<efa<fa<efa<Hga<�ha<-ja<�ka<�ma<�  �  �pa<�qa<Xra</ra<eqa<)pa<?na<?la<�ia<>ga<�da<�ba<�aa<�`a<�`a<�aa<Tca<nea<@ha<Ika<ina<�qa<Kta<�va<�xa<za<�za<�za<qza<�ya<ya<xa<�wa<wa<&wa<�wa<�xa<?za<�{a<~a<�a<�a<�a<�a<"�a<1�a<�a<Ԅa<g�a<��a<za<�}a<�{a<|za<�ya<wya<za<s{a<�}a<+�a<f�a<��a<��a<�a<ďa<7�a<��a<�a<�a<�a<b�a<k�a<h�a<?�a<��a<��a<��a<�a<��a<ӑa<�a<ʔa<1�a<��a<��a<B�a<_�a<��a<��a<��a<��a<��a<S�a<Ћa<f�a<��a<c�a<��a<?�a<Y�a<�a<9�a<�a<��a<��a<��a<�a<��a<��a<�a<��a<�a<ݘa<��a<�a<��a<��a<Ԓa<��a<��a<Y�a<F�a<w�a<ޖa<�a<,�a<��a<�a<��a<��a<�a<��a<E�a<6�a<u�a<��a<E�a<u�a<!�a<��a<�a<�a<��a<�a<U�a<׍a<~�a<q�a<a�a<g�a<�a<	�a<]�a<V�a<֒a<[�a<��a<5�a<�a<�a<ًa<��a<c�a<�a<&�a<,�a<�a<͐a<�a<��a<��a<'�a<Ջa<)�a<%�a<��a<�a<Z|a<�ya<�wa<-va<�ua<�ua<}va<�wa<�ya<�{a<�}a<�a<�a<e�a<��a<ւa<�a<Հa<+a<8}a<A{a<-ya<�wa<�ua<ua<�ta<hta<�ta<tua<~va<=wa<xa<xxa<xxa<xa<�va</ua<�ra<'pa<ma<�ia<�fa<da<	ba<J`a<�_a<m_a<1`a<�aa<vca<�ea<Hha<ka<$ma<#oa<�pa<jqa<�qa<9qa<�pa<9oa<�ma<kla<ka<ja<;ia<2ia<Bia<ja<&ka<�la<na<~oa<�  �  ra<�ra<�ra<Cra<Eqa<�oa<Xma<�ja<ha<Vea<�ba<�`a< _a<S^a<U^a<4_a<�`a<-ca<)fa<via<�la<\pa<|sa<kva<�xa<)za<?{a<�{a<�{a<Y{a<�za<.za<�ya<�ya<�ya<1za<{a<�|a<~a<�a<݁a<��a<��a<�a<k�a<<�a<��a<.�a<Z�a<)�a<�}a<�{a<�ya<xa<*wa<�va<�wa<ya<B{a<�}a<j�a<ڄa<{�a<��a<�a<ّa<��a<*�a<��a<�a<a</�a<V�a<`�a<Œa<;�a<#�a<g�a<�a<�a<6�a<��a<�a<�a<��a<�a<��a<��a<*�a<ޔa<X�a<s�a<��a<Éa<*�a<J�a<��a<s�a<ǃa<�a<��a<�a<�a<��a<�a<�a<��a<v�a<��a<y�a<��a<<�a<m�a<^�a<'�a<�a<�a<W�a<�a<0�a<��a<}�a<��a<��a<��a<V�a<a<��a<��a<`�a<i�a<��a<֐a<��a<��a<��a<��a<��a<��a<0�a<��a<��a<f�a<͆a<��a<P�a<'�a<��a<�a<Z�a<B�a<��a<g�a<��a<z�a</�a<��a<u�a<e�a<��a<;�a<8�a<��a<=�a<"�a<�a<��a<�a<͑a<�a<��a<ڍa</�a<�a<��a<
�a<�}a</za<jwa<0ua<�sa<sa<&sa<ta<}ua<�wa<�ya<<|a<�~a<l�a<�a<��a<�a<ӂa<�a<��a<�~a</}a<N{a<�ya<mxa<�wa<�va<�va<,wa<�wa<Uxa<�xa<Yya<�ya<(ya<3xa<�va<�ta<�qa<�na<ka<ha<�da<�aa<�_a<�]a<�\a<�\a<�]a<?_a<Vaa<�ca<�fa<�ia<2la<�na<\pa<yqa<ra<4ra<�qa<�pa<�oa<tna<Ama<gla<�ka<�ka<�ka<wla<\ma<�na<�oa<qa<�  �  �ra<esa<$sa<wra<qa<oa<�la<�ia<�fa<�ca<!aa<�^a<"]a<[\a<K\a<@]a<�^a<�aa<�da<"ha<�ka<_oa<�ra<�ua<xxa<fza<�{a<u|a<�|a<�|a<|a<�{a<�{a<u{a<�{a<|a<}a<T~a<�a<w�a<�a<��a<��a<��a<��a<d�a<3�a<��a<��a<a<�|a<za<�wa<9va<,ua<�ta<�ua<wa<\ya<\|a<�a<��a<r�a<'�a<��a<]�a<ғa<m�a<v�a<Ԗa<Ӗa<Z�a<��a<+�a<��a<9�a<�a<b�a<�a<ϕa<��a<�a<�a<�a<o�a<d�a<ϙa<��a<��a<\�a<g�a<c�a<C�a<�a<��a<X�a<�a<q�a<́a<�a<�a<{�a<~�a<ލa<	�a<A�a<��a</�a<�a<כa<V�a<�a<��a<��a<��a<��a<�a<Z�a<��a<6�a<��a<B�a<$�a<�a<Кa<3�a<j�a<��a<�a<+�a<Օa<�a<Џa<��a<�a<�a<0�a<��a<�a<%a<�a<��a<��a<#�a<,�a<=�a<*�a<�a<P�a<D�a<~�a<�a<�a<��a<��a<q�a<k�a<0�a<I�a<��a<$�a<8�a<x�a<�a<��a<�a<��a<��a<X�a<T�a<ӏa<n�a<��a<V�a<��a<�a<�{a<�xa<�ua<1sa<�qa<�pa<&qa<*ra<�sa<va<�xa<3{a<�}a<�a<��a<܂a<Z�a<O�a<��a<��a<&�a<�~a<}a<�{a<kza<rya<�xa<�xa<�xa<Yya<�ya<$za<Wza<<za<�ya<sxa<�va<#ta<dqa<�ma<pja<�fa<;ca<?`a<�]a<�[a<�Za<�Za<�[a<r]a<�_a<vba<�ea<�ha<�ka<na<pa<�qa<ura<�ra<zra<�qa<�pa<pa<oa<=na<�ma<qma<�ma<Rna<!oa<0pa< qa<Ira<�  �  �sa<�sa<bsa<vra<�pa<�na<Bla<<ia<	fa<�ba<`a<�]a<\a<,[a<[a<\a<�]a<f`a<}ca<)ga<�ja<�na<�ra<�ua<Zxa<rza<�{a<�|a<Y}a<j}a<}a<�|a<z|a<�|a<�|a<^}a<2~a<ea<րa<r�a<��a<o�a<N�a<��a<ۆa<P�a<�a<Q�a<
�a<k~a<�{a<ya<�va<ua<ta<�sa<qta<�ua<Dxa<K{a<�~a<��a<��a<��a<5�a<-�a<a<��a<Ŗa<]�a<��a<A�a<��a<%�a<��a<J�a<L�a<��a<�a<͖a<�a<�a<��a<��a<ޚa<��a<ߙa<�a<n�a<�a<ߐa<��a<G�a<�a<n�a<B�a<׀a<A�a<��a<ˁa<΃a<q�a<��a<�a<t�a<ȓa<��a<	�a<�a<�a<��a<��a<b�a<��a<��a<��a<��a<o�a<J�a<J�a<��a<<�a<�a<ܚa<��a<ޛa<��a<�a<�a<�a<��a<��a<B�a<��a<$�a<ބa<�a<�a<�~a<�}a<d~a<�a<��a< �a<3�a<h�a<��a<��a<"�a<%�a<��a<S�a<|�a<>�a<��a<m�a<X�a<*�a<U�a<��a<h�a<M�a<��a<��a<��a<�a<q�a<5�a<��a<x�a<��a<?�a<S�a<͆a<�a<�~a<	{a<�wa<tta<ra<�pa<�oa<pa<qa<�ra<ua<�wa<qza<#}a<�a<Z�a<˂a<v�a<��a<)�a<g�a<�a<�a<~a<�|a<{{a<�za<za<�ya<�ya<Eza<�za<{a<{a<�za<�ya<�xa<�va<�sa<�pa<gma<�ia<�ea<5ba<$_a<�\a<�Za<�Ya<�Ya<�Za<W\a<�^a<�aa<�da<�ga<ka<�ma<�oa<�qa<�ra<&sa<sa<�ra<�qa<�pa<�oa<Poa<�na<�na<�na<aoa<pa<*qa<ra<sa<�  �  �ta<�ta<ta<�ra<�pa<�ma<�ia<�ea<yaa<]a<Ya<�Ua<LSa<�Qa<�Qa<�Ra<0Ua<�Xa<�\a<�aa<�fa<�ka<npa<�ta</xa<�za<�|a<�}a<O~a<:~a<�}a<�}a<}a<�|a<�|a<�}a<S~a<�a<��a<P�a<�a<i�a<��a<'�a<��a<��a<لa<�a<�~a<4{a<wa<ysa<�oa<Rma<�ka<ka<�ka<�ma<|pa<ita<9ya<"~a<��a<��a</�a<O�a<��a<ɖa<��a<�a<�a<��a<$�a<l�a<Җa<��a<	�a<7�a<Ӗa<�a<%�a<J�a<V�a<!�a<��a<6�a<ךa<�a<;�a<��a<��a<�a<S�a<0�a<;}a<Aza<bxa<�wa<�wa<�ya<:|a<�a<6�a<ֈa<��a<ܑa<�a<1�a<��a<N�a<.�a<=�a<��a<Мa<ޛa<��a<�a<�a<ߘa<��a<��a<J�a<H�a<�a<ޜa<c�a<G�a<b�a<��a<<�a<��a<֐a<p�a<��a<؂a<o~a<�za<�wa<�ua<2ua<�ua<wa<@za<~a<�a<��a<�a<�a<ǒa<y�a<g�a<��a<�a<��a<חa<��a<��a<K�a<�a<G�a<�a<�a<��a<-�a<��a<q�a<єa<ٔa<H�a<��a<u�a<Z�a<[�a<��a<�a<|za<�ua<�pa<�la<�ia<�ga<�fa<�ga<ia<�ka<8oa<�ra<wa<�za<%~a<�a<�a<?�a<܄a<c�a<`�a< �a<p�a<�~a<L}a<�{a<�za<8za<za<�za<�za<l{a<�{a<�{a<�{a<�za<�xa<vva<9sa<oa<{ja<�ea<Y`a<�[a<_Wa<�Sa<�Qa<~Pa<�Pa<�Qa<,Ta<�Wa<�[a<�_a<rda<�ha<fla<zoa<�qa<Msa<ta<ta<dsa<�ra<�qa<npa<�oa<�na<�na<�na<�oa<�pa<�qa<�ra<�sa<�  �  [ta<vta<�sa<�ra<�pa<�ma<ja<�ea<�aa<q]a<�Ya<`Va<�Sa<�Ra<yRa<�Sa<�Ua<;Ya<Y]a<�aa<�fa<�ka<�pa<�ta<Gxa<�za<�|a<�}a<'~a<~a<z}a<�|a<`|a<>|a<J|a<�|a<�}a<>a<܀a<ςa<��a<W�a<b�a<�a<��a<؆a<̈́a<D�a<�~a<Q{a<xwa<�sa<�pa<na<Ola<�ka<^la<7na<-qa<ua<�ya<�~a<��a<��a<b�a<9�a<��a<Ȗa<:�a<�a<�a<y�a<��a<��a< �a<��a<i�a<��a<P�a<=�a<��a<ٙa<�a<��a<I�a<��a<�a<�a<!�a<��a<��a<B�a<a<��a<�}a<�za<ya</xa<�xa<4za<�|a<o�a<��a<�a<��a<�a<��a<8�a<a<0�a<��a<�a<��a<t�a<U�a<�a<.�a<j�a<@�a<?�a<ܘa<��a<��a<��a<ʜa<=�a<�a<?�a<Ța<D�a<��a<�a<��a<�a<4�a<�~a<>{a<Rxa<�va<�ua<vva<+xa<�za<�~a<�a<�a<+�a<E�a<��a<��a<�a<}�a<٘a<��a<��a<K�a<�a<��a<��a<��a<p�a<g�a<בa<u�a<_�a<&�a<��a<��a<�a<��a<��a<O�a<��a<�a<�a<�za<�ua<Dqa<^ma<Qja<fha<�ga<.ha<�ia<Vla<�oa<?sa<.wa<�za<X~a<��a<5�a<>�a<��a<5�a<M�a<��a<�a<~a<z|a<{a<5za<�ya<�ya<�ya<Oza<�za<�{a<�{a<�{a<�za<�xa<�va<sa<8oa<�ja<�ea<�`a<.\a<Xa<�Ta<ZRa<#Qa<6Qa<wRa<�Ta<Xa<�[a<7`a<�da<�ha<nla<�oa<�qa</sa<�sa<�sa<Rsa<#ra< qa<�oa<�na<-na<na<4na<�na<�oa<)qa<^ra<�sa<�  �  bsa<�sa<�sa<�ra<�pa<�ma<�ja<�fa<�ba<�^a<�Za<�Wa<]Ua<0Ta<Ta<Ua<JWa<�Za<�^a<7ca<ha<�la<Yqa< ua<]xa<�za<I|a<!}a<+}a<�|a<V|a<�{a<{a<�za<�za<L{a<q|a<�}a<�a<��a<s�a<F�a<��a<��a<u�a<ņa<�a<ʂa<�a<B|a<�xa<ua<�qa<toa<�ma<]ma<na<�oa<�ra<qva<�za<�a<��a<~�a<��a<z�a<��a<��a<ؗa<9�a< �a<E�a<��a<��a<��a<!�a<ʓa<�a<�a<ڕa<P�a<��a<�a<��a<��a<��a<��a< �a<j�a<r�a<r�a<N�a<	�a<ւa<Za<b|a<�za<�ya<6za<�{a<]~a<Ɓa<Ʌa<N�a<��a<֒a<d�a<\�a<��a<�a<��a<)�a<x�a<I�a<.�a<Ƙa<��a<�a<��a<��a<g�a<G�a<��a<��a<��a<D�a<��a<��a<��a<a�a<S�a<ˑa<w�a<�a<u�a<D�a<�|a<�ya<xa<~wa<�wa<�ya<l|a<�a<ăa<��a<�a<��a<��a<��a<U�a<(�a<D�a<��a<��a<(�a<��a</�a<�a<%�a<Ϗa<�a<n�a<:�a<:�a<�a<��a<�a<��a<h�a<��a<��a<	�a<��a<�a<|a<wa<�ra<�na<�ka<ja<Pia<�ia<Aka<�ma<�pa<�ta<!xa<�{a<�~a<>�a</�a<�a<3�a<��a<A�a<��a<�~a<�|a<{a<�ya<�xa<xa<(xa<]xa<ya<�ya<jza<�za<�za<8za<�xa<�va<gsa<�oa<jka<�fa<ba<h]a<}Ya<Va<�Sa<�Ra<�Ra<�Sa<OVa<lYa<(]a<kaa<}ea<~ia<�la<�oa<�qa<�ra<bsa<�ra<3ra<�pa<�oa<tna<oma<�la<lla<�la<~ma<�na<�oa<6qa<�ra<�  �  Tra<sa<3sa<jra<qa<�na<�ka<8ha<eda<�`a<(]a<CZa<Xa<�Va<�Va<�Wa<�Ya<]a<�`a<ea<�ia<na<ra<�ua<�xa<yza<�{a<1|a<|a<c{a<zza<iya<�xa<)xa<"xa<�xa<�ya<m{a<B}a<�a<ځa<�a<��a<φa<�a<��a<��a<i�a<΀a<�}a<Nza<*wa<3ta<�qa<�pa< pa<�pa<kra<0ua<�xa<�|a<m�a<)�a<��a<��a<&�a<��a<=�a<8�a<4�a<��a<��a<x�a<&�a<9�a<d�a<H�a<u�a<8�a<y�a<�a<Öa<m�a<ۙa<��a<�a<w�a<-�a<&�a<�a<��a<Ōa<Ĉa<
�a<��a<
a<7}a<v|a<�|a<]~a<׀a<�a<ԇa<Ӌa<��a<��a<!�a<Ǚa<v�a<��a<��a<�a<�a<��a<��a<b�a<?�a<I�a<�a<�a<�a<�a<Q�a<ۘa<4�a<5�a<��a<��a<m�a<��a<�a<��a<Ύa<��a<o�a<|�a<#a<{|a<�za< za<�za<G|a<�~a<�a<��a<w�a<S�a<��a<��a<˕a<�a<��a<T�a<w�a<��a<L�a<k�a<ʏa<y�a<��a<N�a<F�a<�a<ڎa<"�a<Z�a<Y�a<ݒa<�a<�a<h�a<�a<��a<ǆa<c�a<�}a<3ya<�ta<Xqa<�na<�la<�ka<bla<�ma< pa<�ra<"va<�ya<�|a<�a<�a< �a<��a<��a<~�a<��a<�~a<�|a<�za<�xa<wa<va<wua<vua<�ua<�va<�wa<�xa<�ya<�ya<�ya<�xa<�va<#ta<�pa<�la<Aha<�ca<�_a<�[a<�Xa<�Va<jUa<uUa<�Va<�Xa<�[a<3_a<�ba<�fa<eja<�ma<pa<�qa<�ra<�ra<�qa<�pa<Poa<�ma<la<�ja<ja<�ia<ja<�ja<#la<�ma<oa<qa<�  �  �pa<�qa<�ra<Ura<Hqa<�oa<�la<ja<�fa<Aca<�_a<']a<G[a<;Za<;Za<-[a<#]a<�_a<�ca<�ga<�ka<�oa<*sa<iva<�xa<Vza<{a<�za<aza<,ya<xa<�va<�ua<ua<�ta<xua<kva<^xa<\za<�|a<�a< �a<�a<��a<Ɔa<��a<�a<X�a<Q�a<�a<�|a<�ya<�va<ua<�sa<ksa<ta<�ua<:xa<�{a<�a<ƃa<(�a<9�a<��a<��a<��a<��a<'�a<��a<Ӕa<k�a<�a<=�a</�a<#�a<��a<5�a<�a<��a<!�a<H�a<.�a<�a<E�a<:�a<J�a<?�a<��a<%�a<a�a<Ўa<:�a<χa<��a<+�a<��a<�a<A�a<��a<ǃa<ʆa<n�a<��a<�a<�a<�a<�a<d�a<�a<v�a<��a<�a<2�a<K�a<{�a<&�a<��a<Őa<ΐa<Ña<��a<��a<h�a<�a<��a<j�a<�a<X�a<��a<ږa<��a<��a<��a<�a<E�a<�a<�a<#~a<�}a<
~a<sa<��a<��a<�a<��a<�a<Бa<d�a<�a<�a<�a<�a<Ĕa<ɒa<Ԑa<��a<݌a<V�a<K�a<��a<��a<��a<�a<��a<�a<h�a<a�a<͑a<��a<b�a<��a<��a<J�a<Z�a<�a<�{a<�wa<]ta<�qa<pa<aoa<�oa<�pa<�ra<�ua<{xa<�{a<i~a<��a<a�a<�a<m�a<��a<�a<a<�|a<5za<�wa<�ua<�sa<�ra<7ra<Jra<	sa<�sa<iua<�va<�wa<�xa<�xa<]xa<�va<�ta<�qa<Xna<Kja<>fa<_ba<�^a<�[a<�Ya<�Xa<�Xa<�Ya<�[a<o^a<�aa<ea<�ha<�ka<dna<]pa<�qa<ra<Zqa<gpa<�na<�la<�ja<)ia<�ga<�fa<�fa<�fa<�ga<;ia<
ka<ma<�na<�  �  �na<�pa<�qa<ra<�qa<qpa<mna<�ka<ia<	fa<Eca<�`a<_a<,^a<*^a<_a<�`a<�ca<�fa<Oja<�ma<rqa<�ta<,wa<�xa<�ya<za<�ya<Txa<�va<ua<rsa<�qa<<qa<�pa<fqa<�ra<�ta<�va<�ya<�|a<�a<��a<��a<�a<��a<��a<��a<΃a<��a<Qa<�|a<�za<�xa<�wa<mwa<xa<�ya<�{a<2a<��a<��a<1�a<��a<�a<!�a<��a<F�a<�a<E�a<��a<��a<�a<�a<X�a<s�a<�a<:�a<L�a<��a<�a<[�a<��a<�a<��a<&�a<��a<t�a<o�a<��a<�a<�a<�a<݊a<F�a<�a<t�a<�a<9�a<i�a<��a<9�a<B�a<��a<��a<��a<��a<x�a<+�a<�a<J�a<ǘa<��a<h�a<3�a<�a<G�a<6�a<��a< �a<�a<_�a<{�a<��a<��a<��a<9�a<�a<	�a<S�a<Ǘa<f�a<y�a<=�a<΋a<��a<Ӆa<|�a<�a<��a<�a<4�a<c�a<އa<ߊa<�a<��a<P�a<'�a<1�a<q�a<�a<��a<��a<K�a<�a<t�a<$�a<��a<d�a<�a<O�a<�a<��a<z�a<O�a<0�a<ҏa<��a<��a<Y�a<�a<ڌa<Ɖa<N�a<��a<�~a<P{a<"xa<�ua<ta<csa<�sa<�ta<�va<�xa<A{a<�}a<�a<ށa<�a<,�a<��a<n�a<�a<�|a<za<4wa<Lta<�qa<pa<�na<<na<�na<Boa<�pa<}ra<ta<�ua<5wa<�wa<�wa<�va<jua<sa<�oa<�la<	ia<lea<gba<�_a<�]a<�\a<�\a<�]a<�_a<�aa<�da<�ga<�ja<Ema<ooa<�pa<Mqa<qa<.pa<�na<fla<ja<�ga<�ea<�ca<�ba<�ba<�ba< da<�ea<�ga<9ja<�la<�  �  �la<(oa<�pa<�qa<�qa<Fqa<pa<�ma<�ka<ia<�fa<�da<.ca<sba<Uba<aca<�da<Xga<ja<Lma<�pa<asa<va<�wa<,ya<wya<ya<�wa<va<0ta<�qa<�oa<+na<&ma<�la<$ma<�na<�pa<isa<cva<	za<t}a<��a<W�a<B�a<��a<��a<��a<��a<��a<�a<�a<4~a<�|a<�{a<�{a<:|a<�}a<�a<ӂa<υa<f�a<��a<��a<	�a<��a<��a<��a<�a<X�a<X�a<�a<j�a<e�a<c�a<V�a<��a<�a<.�a<�a<_�a<��a<�a<��a<A�a<�a<<�a<��a<�a<�a<�a<��a<��a<%�a<�a<މa<ňa<�a<{�a<��a<X�a<��a<[�a<Z�a<ٕa<D�a<�a<ߚa<�a<>�a<�a<��a<J�a<k�a<��a<M�a<A�a<�a<k�a<܈a<܉a<��a<�a<{�a<I�a<��a<×a<�a<ؙa<��a<��a<��a<��a<�a<ގa<�a<��a<��a<^�a<��a<@�a<5�a<�a<;�a<ݍa<��a<��a<��a<ڕa<y�a<�a<�a<�a<}�a<΍a<��a<�a<V�a<t�a<7�a<��a<4�a<�a< �a<�a<��a<ڋa<эa<w�a<3�a<g�a<|�a<�a<��a<��a<z�a<�a<�~a<�{a<�ya<Dxa<�wa<�wa<}xa<"za<�{a<~a<�a<Ła<�a<n�a<M�a<�a<B�a<�}a<�za<Swa<�sa<�pa<�ma<�ka<yja<ja<mja<fka<.ma<oa<�qa<�sa<|ua<�va<Mwa<6wa<va<hta<�qa<oa<�ka<�ha<fa<�ca<ba<�`a<aa<�aa<Hca<^ea<�ga<vja<�la<�na<[pa<)qa<2qa<>pa<�na<xla<ja<ga<Uda<�aa<�_a<�^a<H^a<�^a<�_a<�aa<]da<!ga<*ja<�  �  �ja<�ma<�oa<�qa<;ra<9ra<�qa<pa<*na<;la<Mja<kha<8ga<�fa<�fa<|ga<�ha<�ja<�ma<:pa<�ra<yua<jwa<�xa<<ya<ya<xa<<va<�sa<mqa<�na<_la<eja<�ha<�ha<�ha<Uja<�la<�oa<#sa<wa<�za<�~a<�a<��a<t�a<��a<��a<b�a<@�a<��a<M�a<��a<z�a<�a<�a<o�a<�a<Ƀa<V�a<D�a<�a<�a<t�a<+�a<P�a<��a<�a<��a<z�a<�a<0�a<0�a<Åa<�a<�a<��a<ׁa<�a<�a<Їa<Պa<H�a<z�a<z�a<�a<ǘa<��a<ڙa<5�a<�a<��a<Γa<��a<��a<ߍa<��a<R�a<��a<��a<�a<K�a<��a<ϕa<�a<יa<ޚa<6�a<Śa<��a<t�a<��a<��a<h�a<?�a<��a<8�a<Ǆa<>�a<��a<ǅa<�a<v�a<p�a<��a<��a<6�a<F�a<��a<�a<��a<}�a<��a<\�a<�a<��a<N�a<��a<��a<�a<\�a<;�a<��a<ʎa<͐a<ߒa<ʔa<�a<��a<��a<��a<�a<a�a<V�a<�a<��a<`�a<��a<Fa<�}a<�}a<�}a</a<X�a<��a<��a<W�a<�a<1�a<��a<0�a<�a<��a<Z�a<�a<�a<U�a<n�a<�a<�}a<u|a<�{a<�{a<k|a<�}a<Ea<Àa<\�a<��a<#�a<�a<#�a<|�a<a<�{a<(xa<tta<}pa<#ma<�ia<�ga<Vfa<�ea<3fa<�ga<�ia<�ka<�na<Rqa<�sa<�ua<�va<1wa<�va<�ua<�sa<rqa<�na<?la<�ia<�ga<1fa<Bea<>ea<�ea<
ga<�ha<�ja<�la<�na<�pa<Uqa<�qa<�pa<�oa<Yma<�ja<hga<da<�`a<D^a<�[a<�Za<Za<�Za<�[a<2^a<�`a<da<{ga<�  �  �ha<la<oa<*qa<�ra<0sa<�ra<ra<�pa<oa<oma<la<ka<lja<�ja<7ka<�la<una<�pa<�ra<;ua<=wa<�xa<�ya<iya<�xa<�va<�ta<ra<�na<�ka<�ha<�fa<$ea<�da<ea<rfa<�ha<la<pa<Qta<�xa<}a<��a<�a<I�a<"�a<ֈa<��a<W�a<L�a<?�a<��a<F�a<��a<҃a<��a<��a<��a<��a<A�a<��a<�a<ܒa<B�a<��a<o�a<w�a<T�a<�a<ʋa<e�a<8�a<	�a<�a</~a<�}a<�}a<#a<Q�a<<�a<�a<��a<��a<��a<ޕa<Q�a<a<��a<S�a<��a<:�a<��a<Ŕa<��a<��a<��a<e�a<��a<t�a<Βa<u�a<z�a<G�a<�a<�a<�a<��a<{�a<��a<�a<��a<B�a<��a<�a<ʄa<t�a<��a<N�a<��a<��a<"�a<-�a<��a<�a<Ǒa<��a<f�a<-�a<C�a<��a<��a<��a<ʖa<۔a<ǒa<�a<|�a<X�a<�a<�a<�a<9�a<ߑa<��a<0�a<��a<:�a<��a<��a<7�a<ؒa<ُa<q�a<c�a<��a<�a<�}a<r{a<�ya<�ya<za<p{a<�}a<��a<΃a<�a<Y�a<��a<�a<�a<��a<�a<��a<�a<��a<G�a<��a<��a<��a<z�a<�a<�a<>�a<�a<A�a<f�a<}�a<�a<:�a<��a<
�a<�a<�}a<?za<va<�qa<�ma<jia<:fa<�ca<Uba<�aa<bba<�ca<fa<ia<
la<coa<8ra<�ta<bva<Ewa<�wa<�va<�ua<�sa<�qa<Qoa<ma<pka<�ia<Uia<ia<�ia<�ja<la<�ma<coa<�pa<�qa<Xra<�qa<�pa<�na<�ka<�ha<ea<Xaa<�]a<}Za</Xa<�Va<.Va<�Va<Xa<gZa<�]a<Saa< ea<�  �  ga<�ja<Zna<�pa<�ra<�sa<ta<�sa<�ra<�qa<*pa<�na<0na<�ma< na<�na<�oa<[qa<[sa<eua<Dwa<�xa<�ya<	za<xya<Kxa< va<Qsa<%pa<�la<@ia<fa<�ca<�aa<-aa<�aa<ca<�ea<'ia<_ma<�qa<�va<i{a<�a<q�a<>�a<T�a<��a<+�a<#�a<��a<��a<чa<A�a<��a<�a<ˇa<݈a<��a<��a<Ɏa<��a<�a<U�a<E�a<6�a<o�a<��a<O�a<U�a<ȉa<�a<��a<5a<�|a<�za<za<lza<�{a<O~a<r�a<N�a<U�a<��a<��a<��a<�a<˙a<�a<�a<�a<5�a<�a<b�a<ەa<Δa<ޓa<��a<̓a<��a<��a<:�a<�a<y�a<��a<p�a<��a<śa<N�a<
�a<̔a<7�a<)�a<�a<F�a<�a<Ea<}}a<�|a<;}a<�~a<@�a<d�a<�a<�a<��a<{�a<��a<�a<]�a<&�a<��a<=�a<�a<P�a<��a<ړa<��a<��a<k�a<j�a<1�a< �a<��a<��a<9�a<�a<p�a<�a<ǖa<�a<�a<w�a<��a<5�a<�a<~a<�za<8xa<�va<va<�va<Uxa<�za<�}a<`�a<�a<��a<��a<a�a<��a<Ӑa<��a<"�a<Ύa<�a<Ɗa<��a<��a<�a<��a<�a<Ԃa<E�a<ԃa<Ʉa<��a<[�a<��a<=�a<��a<
�a<p�a<�|a<�xa<ta<Hoa<�ja<�fa<+ca<�`a<�^a<o^a<!_a<�`a<Aca<ofa<�ia<qma<�pa<�sa<va<Mwa<xa<�wa< wa<�ua<�sa<�qa<�oa<�na<,ma<�la<`la<�la<�ma<�na<Mpa<�qa<�ra<sa<sa<ra<rpa<na<�ja<ga<�ba<�^a<�Za<�Wa<Ua<ISa<�Ra<7Sa<�Ta<�Wa<�Za<�^a<�ba<�  �  �ea<ja<�ma<�pa<�ra<Cta<�ta<�ta</ta<Esa<ora<Zqa<�pa<Upa<}pa<3qa<Pra<�sa<�ua<	wa<�xa<�ya<�za<fza<�ya<�wa<kua<ara<�na<ka<-ga<�ca<(aa<0_a<�^a<�^a<k`a<ca<�fa<,ka<1pa<<ua<.za<�~a<��a<<�a<��a<B�a<$�a<N�a<�a<��a<.�a<��a<��a<��a<N�a<��a<��a<�a<Аa<��a<+�a<V�a<ڕa<��a<y�a<G�a<��a<'�a<R�a<`�a<S�a<�|a<za<(xa<swa<�wa< ya<�{a<6a<,�a<Ƈa<+�a<z�a<R�a<c�a<�a<d�a<8�a<�a<��a<��a<��a<>�a<;�a<��a<:�a<f�a<3�a< �a<��a<a<��a<՜a<^�a<�a<
�a< �a<E�a<�a<�a<��a<@�a<�a<�a<�|a<�za<*za<�za<|a<�~a<.�a<(�a<��a<��a<��a<�a<��a<��a<��a<�a<L�a<b�a<�a<ȗa<?�a<(�a<C�a<�a<�a<��a<��a<��a<��a<��a<�a<7�a<f�a<�a<o�a<N�a<��a<'�a<��a< �a<�{a<Sxa<~ua<�sa<msa<�sa<�ua<uxa<�{a<�a<��a<s�a<�a<��a<��a<�a<�a<�a<��a<n�a<��a<��a<��a<��a<G�a<��a<��a<��a<1�a<Іa<8�a<��a<��a<҆a<L�a<�a<�a<|a<twa<�ra<�ma<�ha<Uda<�`a<�]a<A\a<�[a<_\a<L^a<aa<Mda<@ha<la<�oa<�ra<rua<nwa<\xa<�xa<
xa<wa<�ua<ta<[ra<�pa<�oa<)oa<�na<qoa<pa<-qa<ra<sa<�sa<ta<�sa<Ura<Epa<Hma<�ia<�ea<naa<�\a<�Xa<GUa<SRa<�Pa<Pa<�Pa<4Ra<Ua<�Xa<�\a<daa<�  �  �da<[ia<;ma<�pa<sa<�ta<pua<�ua<Wua<mta<�sa<�ra<0ra<�qa<'ra<�ra<�sa<ua<�va<4xa<�ya<�za<�za<�za<�ya<�wa<�ta<�qa<�ma<�ia<�ea<�ba<�_a<�]a<�\a<J]a<�^a<�aa<tea<�ia<�na<8ta<Wya<K~a<r�a<,�a<ʈa<��a<ʋa<R�a<C�a<݋a<_�a<�a<��a<=�a<�a<��a<e�a<�a<��a<��a<3�a<�a<?�a<��a<w�a<�a<�a<W�a<Y�a<�a<a<�{a<�xa<�va<�ua<(va<�wa<Yza<�}a<�a<��a<7�a<��a<ӓa<0�a<�a<��a<��a<�a<��a<��a<��a<{�a<��a< �a<ݗa<�a<��a<z�a<��a<�a<!�a<ϝa<�a<_�a<0�a<	�a<�a<T�a<�a<��a<��a<ρa<~a<'{a<Iya<�xa<ya<�za<`}a<�a<�a<Z�a<��a<��a<��a<��a<��a<�a<j�a<G�a<��a<6�a<��a<��a<��a<Ǖa<��a<��a<�a<ʖa<ݗa<ʘa<��a<��a<��a<��a<
�a<F�a<ېa<��a<3�a<u�a<�~a<�za<�va<ta<Wra<�qa<|ra<Bta<	wa<~za<e~a<��a<��a<h�a<b�a<�a<I�a<�a<��a<��a<��a<�a<�a<]�a<��a<�a<=�a<�a<�a<e�a<��a<l�a<��a<5�a<8�a<�a<�a<za<x{a<�va<�qa<^la<fga<�ba<$_a<Q\a<�Za<+Za<�Za<�\a<�_a<ca<�fa<ka<�na<ura<?ua<�wa<�xa<ya<�xa<xa<�va<2ua<�sa<Zra<Nqa<�pa<�pa<�pa<gqa<Wra<Csa<<ta<�ta<�ta<�sa<{ra<.pa<�la<<ia<�da<R`a<�[a<�Wa<�Sa<�Pa<Oa<jNa<Oa<�Pa<�Sa<XWa<�[a<=`a<�  �  �da<"ia<Ima<�pa<�ra<�ta<�ua<�ua<oua<�ta<*ta<asa<�ra<\ra<�ra<"sa<}ta<�ua<3wa<�xa<�ya<�za<9{a<�za<�ya<�wa<�ta<eqa<�ma<�ia<�ea<�aa<_a<!]a<D\a<�\a<K^a<�`a<�da<�ia<|na<ta<>ya<~a<��a<�a<��a<�a<��a<r�a<�a<O�a<	�a<Ӌa<z�a<Ջa<��a<t�a<8�a<Ɛa<k�a<��a<I�a<2�a<��a<��a<\�a<�a<�a<4�a<6�a<��a<�~a<�za<�wa<va<%ua<}ua<wa<�ya<<}a<��a<5�a<�a<��a<��a<8�a<��a<��a<��a<�a<��a<�a<*�a<1�a<n�a<~�a<��a<�a<7�a<4�a<M�a<O�a<E�a<��a<*�a<��a<�a<��a<�a<!�a<�a<\�a<��a<R�a<c}a<{za<�xa<�wa<_xa<za<�|a<a�a<��a<�a<��a<��a<��a<��a<��a<�a<��a<n�a<��a<��a<��a<G�a<A�a<J�a<2�a<�a<Ֆa<|�a<d�a<$�a<əa<%�a<�a<ɘa<�a<D�a<Ȑa<��a<�a<0�a<r~a<�ya<3va<osa<�qa<&qa<�qa<�sa<]va<za<�}a<w�a<��a<0�a<{�a<ʏa<;�a<)�a<��a<�a<ُa<W�a<��a<-�a<{�a<}�a<ڇa<l�a<ڇa<�a<k�a<��a<��a<c�a<�a<z�a<��a<�a<B{a<�va<{qa<�ka<ga<Gba<q^a<�[a<�Ya<Ya<TZa<-\a<_a<�ba<�fa<�ja<�na<Sra<Hua<awa<�xa<Sya<ya<(xa<�va<�ua<Mta<!sa<�qa<oqa<qa<uqa<"ra<�ra<�sa<`ta<�ta<�ta<ta<`ra<pa<ma<ia<�da<`a<G[a<Wa<Sa<9Pa<lNa<�Ma<\Na<"Pa<�Ra<�Va</[a< `a<�  �  �da<[ia<;ma<�pa<sa<�ta<pua<�ua<Wua<mta<�sa<�ra<0ra<�qa<'ra<�ra<�sa<ua<�va<4xa<�ya<�za<�za<�za<�ya<�wa<�ta<�qa<�ma<�ia<�ea<�ba<�_a<�]a<�\a<J]a<�^a<�aa<tea<�ia<�na<8ta<Wya<K~a<r�a<,�a<ʈa<��a<ʋa<R�a<C�a<݋a<_�a<�a<��a<=�a<�a<��a<e�a<�a<��a<��a<3�a<�a<?�a<��a<w�a<�a<�a<W�a<Y�a<�a<a<�{a<�xa<�va<�ua<(va<�wa<Yza<�}a<�a<��a<7�a<��a<ӓa<0�a<�a<��a<��a<�a<��a<��a<��a<{�a<��a< �a<ݗa<�a<��a<z�a<��a<�a<!�a<ϝa<�a<_�a<0�a<	�a<�a<T�a<�a<��a<��a<ρa<~a<'{a<Iya<�xa<ya<�za<`}a<�a<�a<Z�a<��a<��a<��a<��a<��a<�a<j�a<G�a<��a<6�a<��a<��a<��a<Ǖa<��a<��a<�a<ʖa<ݗa<ʘa<��a<��a<��a<��a<
�a<F�a<ېa<��a<3�a<u�a<�~a<�za<�va<ta<Wra<�qa<|ra<Bta<	wa<~za<e~a<��a<��a<h�a<b�a<�a<I�a<�a<��a<��a<��a<�a<�a<]�a<��a<�a<=�a<�a<�a<e�a<��a<l�a<��a<5�a<8�a<�a<�a<za<x{a<�va<�qa<^la<fga<�ba<$_a<Q\a<�Za<+Za<�Za<�\a<�_a<ca<�fa<ka<�na<ura<?ua<�wa<�xa<ya<�xa<xa<�va<2ua<�sa<Zra<Nqa<�pa<�pa<�pa<gqa<Wra<Csa<<ta<�ta<�ta<�sa<{ra<.pa<�la<<ia<�da<R`a<�[a<�Wa<�Sa<�Pa<Oa<jNa<Oa<�Pa<�Sa<XWa<�[a<=`a<�  �  �ea<ja<�ma<�pa<�ra<Cta<�ta<�ta</ta<Esa<ora<Zqa<�pa<Upa<}pa<3qa<Pra<�sa<�ua<	wa<�xa<�ya<�za<fza<�ya<�wa<kua<ara<�na<ka<-ga<�ca<(aa<0_a<�^a<�^a<k`a<ca<�fa<,ka<1pa<<ua<.za<�~a<��a<<�a<��a<B�a<$�a<N�a<�a<��a<.�a<��a<��a<��a<N�a<��a<��a<�a<Аa<��a<+�a<V�a<ڕa<��a<y�a<G�a<��a<'�a<R�a<`�a<S�a<�|a<za<(xa<swa<�wa< ya<�{a<6a<,�a<Ƈa<+�a<z�a<R�a<c�a<�a<d�a<8�a<�a<��a<��a<��a<>�a<;�a<��a<:�a<f�a<3�a< �a<��a<a<��a<՜a<^�a<�a<
�a< �a<E�a<�a<�a<��a<@�a<�a<�a<�|a<�za<*za<�za<|a<�~a<.�a<(�a<��a<��a<��a<�a<��a<��a<��a<�a<L�a<b�a<�a<ȗa<?�a<(�a<C�a<�a<�a<��a<��a<��a<��a<��a<�a<7�a<f�a<�a<o�a<N�a<��a<'�a<��a< �a<�{a<Sxa<~ua<�sa<msa<�sa<�ua<uxa<�{a<�a<��a<s�a<�a<��a<��a<�a<�a<�a<��a<n�a<��a<��a<��a<��a<G�a<��a<��a<��a<1�a<Іa<8�a<��a<��a<҆a<L�a<�a<�a<|a<twa<�ra<�ma<�ha<Uda<�`a<�]a<A\a<�[a<_\a<L^a<aa<Mda<@ha<la<�oa<�ra<rua<nwa<\xa<�xa<
xa<wa<�ua<ta<[ra<�pa<�oa<)oa<�na<qoa<pa<-qa<ra<sa<�sa<ta<�sa<Ura<Epa<Hma<�ia<�ea<naa<�\a<�Xa<GUa<SRa<�Pa<Pa<�Pa<4Ra<Ua<�Xa<�\a<daa<�  �  ga<�ja<Zna<�pa<�ra<�sa<ta<�sa<�ra<�qa<*pa<�na<0na<�ma< na<�na<�oa<[qa<[sa<eua<Dwa<�xa<�ya<	za<xya<Kxa< va<Qsa<%pa<�la<@ia<fa<�ca<�aa<-aa<�aa<ca<�ea<'ia<_ma<�qa<�va<i{a<�a<q�a<>�a<T�a<��a<+�a<#�a<��a<��a<чa<A�a<��a<�a<ˇa<݈a<��a<��a<Ɏa<��a<�a<U�a<E�a<6�a<o�a<��a<O�a<U�a<ȉa<�a<��a<5a<�|a<�za<za<lza<�{a<O~a<r�a<N�a<U�a<��a<��a<��a<�a<˙a<�a<�a<�a<5�a<�a<b�a<ەa<Δa<ޓa<��a<̓a<��a<��a<:�a<�a<y�a<��a<p�a<��a<śa<N�a<
�a<̔a<7�a<)�a<�a<F�a<�a<Ea<}}a<�|a<;}a<�~a<@�a<d�a<�a<�a<��a<{�a<��a<�a<]�a<&�a<��a<=�a<�a<P�a<��a<ړa<��a<��a<k�a<j�a<1�a< �a<��a<��a<9�a<�a<p�a<�a<ǖa<�a<�a<w�a<��a<5�a<�a<~a<�za<8xa<�va<va<�va<Uxa<�za<�}a<`�a<�a<��a<��a<a�a<��a<Ӑa<��a<"�a<Ύa<�a<Ɗa<��a<��a<�a<��a<�a<Ԃa<E�a<ԃa<Ʉa<��a<[�a<��a<=�a<��a<
�a<p�a<�|a<�xa<ta<Hoa<�ja<�fa<+ca<�`a<�^a<o^a<!_a<�`a<Aca<ofa<�ia<qma<�pa<�sa<va<Mwa<xa<�wa< wa<�ua<�sa<�qa<�oa<�na<,ma<�la<`la<�la<�ma<�na<Mpa<�qa<�ra<sa<sa<ra<rpa<na<�ja<ga<�ba<�^a<�Za<�Wa<Ua<ISa<�Ra<7Sa<�Ta<�Wa<�Za<�^a<�ba<�  �  �ha<la<oa<*qa<�ra<0sa<�ra<ra<�pa<oa<oma<la<ka<lja<�ja<7ka<�la<una<�pa<�ra<;ua<=wa<�xa<�ya<iya<�xa<�va<�ta<ra<�na<�ka<�ha<�fa<$ea<�da<ea<rfa<�ha<la<pa<Qta<�xa<}a<��a<�a<I�a<"�a<ֈa<��a<W�a<L�a<?�a<��a<F�a<��a<҃a<��a<��a<��a<��a<A�a<��a<�a<ܒa<B�a<��a<o�a<w�a<T�a<�a<ʋa<e�a<8�a<	�a<�a</~a<�}a<�}a<#a<Q�a<<�a<�a<��a<��a<��a<ޕa<Q�a<a<��a<S�a<��a<:�a<��a<Ŕa<��a<��a<��a<e�a<��a<t�a<Βa<u�a<z�a<G�a<�a<�a<�a<��a<{�a<��a<�a<��a<B�a<��a<�a<ʄa<t�a<��a<N�a<��a<��a<"�a<-�a<��a<�a<Ǒa<��a<f�a<-�a<C�a<��a<��a<��a<ʖa<۔a<ǒa<�a<|�a<X�a<�a<�a<�a<9�a<ߑa<��a<0�a<��a<:�a<��a<��a<7�a<ؒa<ُa<q�a<c�a<��a<�a<�}a<r{a<�ya<�ya<za<p{a<�}a<��a<΃a<�a<Y�a<��a<�a<�a<��a<�a<��a<�a<��a<G�a<��a<��a<��a<z�a<�a<�a<>�a<�a<A�a<f�a<}�a<�a<:�a<��a<
�a<�a<�}a<?za<va<�qa<�ma<jia<:fa<�ca<Uba<�aa<bba<�ca<fa<ia<
la<coa<8ra<�ta<bva<Ewa<�wa<�va<�ua<�sa<�qa<Qoa<ma<pka<�ia<Uia<ia<�ia<�ja<la<�ma<coa<�pa<�qa<Xra<�qa<�pa<�na<�ka<�ha<ea<Xaa<�]a<}Za</Xa<�Va<.Va<�Va<Xa<gZa<�]a<Saa< ea<�  �  �ja<�ma<�oa<�qa<;ra<9ra<�qa<pa<*na<;la<Mja<kha<8ga<�fa<�fa<|ga<�ha<�ja<�ma<:pa<�ra<yua<jwa<�xa<<ya<ya<xa<<va<�sa<mqa<�na<_la<eja<�ha<�ha<�ha<Uja<�la<�oa<#sa<wa<�za<�~a<�a<��a<t�a<��a<��a<b�a<@�a<��a<M�a<��a<z�a<�a<�a<o�a<�a<Ƀa<V�a<D�a<�a<�a<t�a<+�a<P�a<��a<�a<��a<z�a<�a<0�a<0�a<Åa<�a<�a<��a<ׁa<�a<�a<Їa<Պa<H�a<z�a<z�a<�a<ǘa<��a<ڙa<5�a<�a<��a<Γa<��a<��a<ߍa<��a<R�a<��a<��a<�a<K�a<��a<ϕa<�a<יa<ޚa<6�a<Śa<��a<t�a<��a<��a<h�a<?�a<��a<8�a<Ǆa<>�a<��a<ǅa<�a<v�a<p�a<��a<��a<6�a<F�a<��a<�a<��a<}�a<��a<\�a<�a<��a<N�a<��a<��a<�a<\�a<;�a<��a<ʎa<͐a<ߒa<ʔa<�a<��a<��a<��a<�a<a�a<V�a<�a<��a<`�a<��a<Fa<�}a<�}a<�}a</a<X�a<��a<��a<W�a<�a<1�a<��a<0�a<�a<��a<Z�a<�a<�a<U�a<n�a<�a<�}a<u|a<�{a<�{a<k|a<�}a<Ea<Àa<\�a<��a<#�a<�a<#�a<|�a<a<�{a<(xa<tta<}pa<#ma<�ia<�ga<Vfa<�ea<3fa<�ga<�ia<�ka<�na<Rqa<�sa<�ua<�va<1wa<�va<�ua<�sa<rqa<�na<?la<�ia<�ga<1fa<Bea<>ea<�ea<
ga<�ha<�ja<�la<�na<�pa<Uqa<�qa<�pa<�oa<Yma<�ja<hga<da<�`a<D^a<�[a<�Za<Za<�Za<�[a<2^a<�`a<da<{ga<�  �  �la<(oa<�pa<�qa<�qa<Fqa<pa<�ma<�ka<ia<�fa<�da<.ca<sba<Uba<aca<�da<Xga<ja<Lma<�pa<asa<va<�wa<,ya<wya<ya<�wa<va<0ta<�qa<�oa<+na<&ma<�la<$ma<�na<�pa<isa<cva<	za<t}a<��a<W�a<B�a<��a<��a<��a<��a<��a<�a<�a<4~a<�|a<�{a<�{a<:|a<�}a<�a<ӂa<υa<f�a<��a<��a<	�a<��a<��a<��a<�a<X�a<X�a<�a<j�a<e�a<c�a<V�a<��a<�a<.�a<�a<_�a<��a<�a<��a<A�a<�a<<�a<��a<�a<�a<�a<��a<��a<%�a<�a<މa<ňa<�a<{�a<��a<X�a<��a<[�a<Z�a<ٕa<D�a<�a<ߚa<�a<>�a<�a<��a<J�a<k�a<��a<M�a<A�a<�a<k�a<܈a<܉a<��a<�a<{�a<I�a<��a<×a<�a<ؙa<��a<��a<��a<��a<�a<ގa<�a<��a<��a<^�a<��a<@�a<5�a<�a<;�a<ݍa<��a<��a<��a<ڕa<y�a<�a<�a<�a<}�a<΍a<��a<�a<V�a<t�a<7�a<��a<4�a<�a< �a<�a<��a<ڋa<эa<w�a<3�a<g�a<|�a<�a<��a<��a<z�a<�a<�~a<�{a<�ya<Dxa<�wa<�wa<}xa<"za<�{a<~a<�a<Ła<�a<n�a<M�a<�a<B�a<�}a<�za<Swa<�sa<�pa<�ma<�ka<yja<ja<mja<fka<.ma<oa<�qa<�sa<|ua<�va<Mwa<6wa<va<hta<�qa<oa<�ka<�ha<fa<�ca<ba<�`a<aa<�aa<Hca<^ea<�ga<vja<�la<�na<[pa<)qa<2qa<>pa<�na<xla<ja<ga<Uda<�aa<�_a<�^a<H^a<�^a<�_a<�aa<]da<!ga<*ja<�  �  �na<�pa<�qa<ra<�qa<qpa<mna<�ka<ia<	fa<Eca<�`a<_a<,^a<*^a<_a<�`a<�ca<�fa<Oja<�ma<rqa<�ta<,wa<�xa<�ya<za<�ya<Txa<�va<ua<rsa<�qa<<qa<�pa<fqa<�ra<�ta<�va<�ya<�|a<�a<��a<��a<�a<��a<��a<��a<΃a<��a<Qa<�|a<�za<�xa<�wa<mwa<xa<�ya<�{a<2a<��a<��a<1�a<��a<�a<!�a<��a<F�a<�a<E�a<��a<��a<�a<�a<X�a<s�a<�a<:�a<L�a<��a<�a<[�a<��a<�a<��a<&�a<��a<t�a<o�a<��a<�a<�a<�a<݊a<F�a<�a<t�a<�a<9�a<i�a<��a<9�a<B�a<��a<��a<��a<��a<x�a<+�a<�a<J�a<ǘa<��a<h�a<3�a<�a<G�a<6�a<��a< �a<�a<_�a<{�a<��a<��a<��a<9�a<�a<	�a<S�a<Ǘa<f�a<y�a<=�a<΋a<��a<Ӆa<|�a<�a<��a<�a<4�a<c�a<އa<ߊa<�a<��a<P�a<'�a<1�a<q�a<�a<��a<��a<K�a<�a<t�a<$�a<��a<d�a<�a<O�a<�a<��a<z�a<O�a<0�a<ҏa<��a<��a<Y�a<�a<ڌa<Ɖa<N�a<��a<�~a<P{a<"xa<�ua<ta<csa<�sa<�ta<�va<�xa<A{a<�}a<�a<ށa<�a<,�a<��a<n�a<�a<�|a<za<4wa<Lta<�qa<pa<�na<<na<�na<Boa<�pa<}ra<ta<�ua<5wa<�wa<�wa<�va<jua<sa<�oa<�la<	ia<lea<gba<�_a<�]a<�\a<�\a<�]a<�_a<�aa<�da<�ga<�ja<Ema<ooa<�pa<Mqa<qa<.pa<�na<fla<ja<�ga<�ea<�ca<�ba<�ba<�ba< da<�ea<�ga<9ja<�la<�  �  �pa<�qa<�ra<Ura<Hqa<�oa<�la<ja<�fa<Aca<�_a<']a<G[a<;Za<;Za<-[a<#]a<�_a<�ca<�ga<�ka<�oa<*sa<iva<�xa<Vza<{a<�za<aza<,ya<xa<�va<�ua<ua<�ta<xua<kva<^xa<\za<�|a<�a< �a<�a<��a<Ɔa<��a<�a<X�a<Q�a<�a<�|a<�ya<�va<ua<�sa<ksa<ta<�ua<:xa<�{a<�a<ƃa<(�a<9�a<��a<��a<��a<��a<'�a<��a<Ӕa<k�a<�a<=�a</�a<#�a<��a<5�a<�a<��a<!�a<H�a<.�a<�a<E�a<:�a<J�a<?�a<��a<%�a<a�a<Ўa<:�a<χa<��a<+�a<��a<�a<A�a<��a<ǃa<ʆa<n�a<��a<�a<�a<�a<�a<d�a<�a<v�a<��a<�a<2�a<K�a<{�a<&�a<��a<Őa<ΐa<Ña<��a<��a<h�a<�a<��a<j�a<�a<X�a<��a<ږa<��a<��a<��a<�a<E�a<�a<�a<#~a<�}a<
~a<sa<��a<��a<�a<��a<�a<Бa<d�a<�a<�a<�a<�a<Ĕa<ɒa<Ԑa<��a<݌a<V�a<K�a<��a<��a<��a<�a<��a<�a<h�a<a�a<͑a<��a<b�a<��a<��a<J�a<Z�a<�a<�{a<�wa<]ta<�qa<pa<aoa<�oa<�pa<�ra<�ua<{xa<�{a<i~a<��a<a�a<�a<m�a<��a<�a<a<�|a<5za<�wa<�ua<�sa<�ra<7ra<Jra<	sa<�sa<iua<�va<�wa<�xa<�xa<]xa<�va<�ta<�qa<Xna<Kja<>fa<_ba<�^a<�[a<�Ya<�Xa<�Xa<�Ya<�[a<o^a<�aa<ea<�ha<�ka<dna<]pa<�qa<ra<Zqa<gpa<�na<�la<�ja<)ia<�ga<�fa<�fa<�fa<�ga<;ia<
ka<ma<�na<�  �  Tra<sa<3sa<jra<qa<�na<�ka<8ha<eda<�`a<(]a<CZa<Xa<�Va<�Va<�Wa<�Ya<]a<�`a<ea<�ia<na<ra<�ua<�xa<yza<�{a<1|a<|a<c{a<zza<iya<�xa<)xa<"xa<�xa<�ya<m{a<B}a<�a<ځa<�a<��a<φa<�a<��a<��a<i�a<΀a<�}a<Nza<*wa<3ta<�qa<�pa< pa<�pa<kra<0ua<�xa<�|a<m�a<)�a<��a<��a<&�a<��a<=�a<8�a<4�a<��a<��a<x�a<&�a<9�a<d�a<H�a<u�a<8�a<y�a<�a<Öa<m�a<ۙa<��a<�a<w�a<-�a<&�a<�a<��a<Ōa<Ĉa<
�a<��a<
a<7}a<v|a<�|a<]~a<׀a<�a<ԇa<Ӌa<��a<��a<!�a<Ǚa<v�a<��a<��a<�a<�a<��a<��a<b�a<?�a<I�a<�a<�a<�a<�a<Q�a<ۘa<4�a<5�a<��a<��a<m�a<��a<�a<��a<Ύa<��a<o�a<|�a<#a<{|a<�za< za<�za<G|a<�~a<�a<��a<w�a<S�a<��a<��a<˕a<�a<��a<T�a<w�a<��a<L�a<k�a<ʏa<y�a<��a<N�a<F�a<�a<ڎa<"�a<Z�a<Y�a<ݒa<�a<�a<h�a<�a<��a<ǆa<c�a<�}a<3ya<�ta<Xqa<�na<�la<�ka<bla<�ma< pa<�ra<"va<�ya<�|a<�a<�a< �a<��a<��a<~�a<��a<�~a<�|a<�za<�xa<wa<va<wua<vua<�ua<�va<�wa<�xa<�ya<�ya<�ya<�xa<�va<#ta<�pa<�la<Aha<�ca<�_a<�[a<�Xa<�Va<jUa<uUa<�Va<�Xa<�[a<3_a<�ba<�fa<eja<�ma<pa<�qa<�ra<�ra<�qa<�pa<Poa<�ma<la<�ja<ja<�ia<ja<�ja<#la<�ma<oa<qa<�  �  bsa<�sa<�sa<�ra<�pa<�ma<�ja<�fa<�ba<�^a<�Za<�Wa<]Ua<0Ta<Ta<Ua<JWa<�Za<�^a<7ca<ha<�la<Yqa< ua<]xa<�za<I|a<!}a<+}a<�|a<V|a<�{a<{a<�za<�za<L{a<q|a<�}a<�a<��a<s�a<F�a<��a<��a<u�a<ņa<�a<ʂa<�a<B|a<�xa<ua<�qa<toa<�ma<]ma<na<�oa<�ra<qva<�za<�a<��a<~�a<��a<z�a<��a<��a<ؗa<9�a< �a<E�a<��a<��a<��a<!�a<ʓa<�a<�a<ڕa<P�a<��a<�a<��a<��a<��a<��a< �a<j�a<r�a<r�a<N�a<	�a<ւa<Za<b|a<�za<�ya<6za<�{a<]~a<Ɓa<Ʌa<N�a<��a<֒a<d�a<\�a<��a<�a<��a<)�a<x�a<I�a<.�a<Ƙa<��a<�a<��a<��a<g�a<G�a<��a<��a<��a<D�a<��a<��a<��a<a�a<S�a<ˑa<w�a<�a<u�a<D�a<�|a<�ya<xa<~wa<�wa<�ya<l|a<�a<ăa<��a<�a<��a<��a<��a<U�a<(�a<D�a<��a<��a<(�a<��a</�a<�a<%�a<Ϗa<�a<n�a<:�a<:�a<�a<��a<�a<��a<h�a<��a<��a<	�a<��a<�a<|a<wa<�ra<�na<�ka<ja<Pia<�ia<Aka<�ma<�pa<�ta<!xa<�{a<�~a<>�a</�a<�a<3�a<��a<A�a<��a<�~a<�|a<{a<�ya<�xa<xa<(xa<]xa<ya<�ya<jza<�za<�za<8za<�xa<�va<gsa<�oa<jka<�fa<ba<h]a<}Ya<Va<�Sa<�Ra<�Ra<�Sa<OVa<lYa<(]a<kaa<}ea<~ia<�la<�oa<�qa<�ra<bsa<�ra<3ra<�pa<�oa<tna<oma<�la<lla<�la<~ma<�na<�oa<6qa<�ra<�  �  [ta<vta<�sa<�ra<�pa<�ma<ja<�ea<�aa<q]a<�Ya<`Va<�Sa<�Ra<yRa<�Sa<�Ua<;Ya<Y]a<�aa<�fa<�ka<�pa<�ta<Gxa<�za<�|a<�}a<'~a<~a<z}a<�|a<`|a<>|a<J|a<�|a<�}a<>a<܀a<ςa<��a<W�a<b�a<�a<��a<؆a<̈́a<D�a<�~a<Q{a<xwa<�sa<�pa<na<Ola<�ka<^la<7na<-qa<ua<�ya<�~a<��a<��a<b�a<9�a<��a<Ȗa<:�a<�a<�a<y�a<��a<��a< �a<��a<i�a<��a<P�a<=�a<��a<ٙa<�a<��a<I�a<��a<�a<�a<!�a<��a<��a<B�a<a<��a<�}a<�za<ya</xa<�xa<4za<�|a<o�a<��a<�a<��a<�a<��a<8�a<a<0�a<��a<�a<��a<t�a<U�a<�a<.�a<j�a<@�a<?�a<ܘa<��a<��a<��a<ʜa<=�a<�a<?�a<Ța<D�a<��a<�a<��a<�a<4�a<�~a<>{a<Rxa<�va<�ua<vva<+xa<�za<�~a<�a<�a<+�a<E�a<��a<��a<�a<}�a<٘a<��a<��a<K�a<�a<��a<��a<��a<p�a<g�a<בa<u�a<_�a<&�a<��a<��a<�a<��a<��a<O�a<��a<�a<�a<�za<�ua<Dqa<^ma<Qja<fha<�ga<.ha<�ia<Vla<�oa<?sa<.wa<�za<X~a<��a<5�a<>�a<��a<5�a<M�a<��a<�a<~a<z|a<{a<5za<�ya<�ya<�ya<Oza<�za<�{a<�{a<�{a<�za<�xa<�va<sa<8oa<�ja<�ea<�`a<.\a<Xa<�Ta<ZRa<#Qa<6Qa<wRa<�Ta<Xa<�[a<7`a<�da<�ha<nla<�oa<�qa</sa<�sa<�sa<Rsa<#ra< qa<�oa<�na<-na<na<4na<�na<�oa<)qa<^ra<�sa<�  �  va<Xva<�ua<�sa<�pa<�la<�ga<Mba<?\a<QVa<�Pa<NLa<�Ha<Ga<�Fa<Ha<)Ka<[Oa<�Ta<0[a<�aa<�ha<�na<*ta<|xa<|a<w~a<�a<�a<�a<Ia<g~a<�}a<-}a<)}a<�}a<�~a<��a<S�a<��a<��a<]�a<��a<�a<~�a<��a<	�a<C�a<�|a<�wa<�qa<�la<�ga<,da<�aa<�`a<faa<�ca<Xga<Cla<�ra<�xa<�a<��a<��a<ˑa<ҕa<�a<�a<��a<��a<�a<�a<Řa<�a<��a<�a<�a<ɗa<�a<��a<2�a<�a<}�a<Ԟa<`�a<˜a<�a<L�a<��a<��a<�a<�a<za<�ta<�pa<na<*ma<�ma<�oa<Usa<xa<�}a<�a<m�a<4�a<��a<��a<�a<o�a<v�a<{�a<�a<מa<n�a<֛a<��a<��a<��a<��a<c�a<R�a<��a<�a<�a<��a<��a<��a<A�a<֘a<��a<H�a<w�a<�a<�|a<�va<�qa<�ma<zka<�ja<xka<na<�qa<�va<C|a<h�a<b�a<Ӎa<��a<H�a<7�a<ךa<Z�a<��a<��a<��a<�a<U�a<��a<�a<֒a<ǒa<��a<f�a<��a<��a<3�a<I�a<��a<͔a<͑a<׍a<ǈa<ɂa<l|a<Wua<�na<�ha<�ca<�_a<[]a<�\a<X]a<�_a<Xca<Fha<Zma<)sa<Rxa<%}a<�a<�a<�a<��a<d�a<Q�a<��a<ˁa<�a<�}a< |a<{a<zza<lza<{a<�{a<�|a<a}a<�}a<{}a<q|a<Kza<�va<�ra<fma<aga<�`a<%Za<Ta<MNa<Ja<�Fa<�Ea<�Ea<dGa<�Ja<"Oa<�Ta<�Za<�`a<<fa<]ka<hoa<�ra<�ta<�ua<�ua<�ta<�sa<pra<�pa<�oa<�na<�na<�na<�oa<�pa<�ra<ta<Lua<�  �  �ua<va<\ua<�sa<�pa<�la< ha<qba<�\a<�Va<�Qa<Ma<�Ia<�Ga<oGa<�Ha<�Ka<#Pa<�Ua<�[a<Oba<�ha<�na<Lta<�xa<|a<A~a<�a<�a<�a<�~a<�}a<�|a<�|a<t|a<}a<~a<�a<��a<�a<*�a<�a<Y�a<�a<g�a<�a<-�a<��a<�|a<�wa<cra<Uma<�ha<�da<}ba<caa<ba<]da<ha<ma<%sa<�ya<W�a<ǆa<�a<�a<�a<�a<��a<g�a<\�a<��a<h�a<�a< �a<e�a< �a<]�a<2�a<[�a<ՙa<��a<#�a<?�a<��a<-�a<Ŝa<,�a<h�a<đa<)�a<Z�a<W�a<�za<�ua<�qa<�na<�ma<Rna<�pa<ta<�xa<�~a<{�a<��a<x�a<Õa<��a<>�a<9�a<B�a<A�a<��a<D�a<��a<!�a<��a<�a<Øa<ݘa<��a<��a<�a<~�a<Ȟa<W�a<W�a<I�a<T�a<�a<Ӕa<��a<��a<l�a<I}a<�wa<�ra<�na<8la<_ka<Fla<�na<jra<\wa<�|a<Âa<��a<�a<Ȓa<��a<7�a<��a<+�a<��a<��a<��a<<�a<��a<]�a<a�a<	�a<(�a<Ԓa<��a<��a<�a<�a<
�a<g�a<��a<��a<��a<�a<�a<�|a<�ua<{oa<`ia<Uda<{`a<�]a<7]a<0^a<�`a<&da<�ha<�ma<osa<�xa<u}a<:�a<-�a<߅a<��a<'�a<�a<?�a<�a<�~a< }a<h{a<Pza<�ya<�ya<Cza<
{a<|a<}a<�}a<L}a<>|a<Eza<wa<�ra<�ma<�ga<Baa<�Za<�Ta<Oa<�Ja<�Ga<Fa<QFa<=Ha<sKa<�Oa<BUa<�Za<�`a<�fa<�ka<�oa<�ra<�ta<ua<gua<�ta<Lsa<�qa<%pa<oa<(na<�ma<*na<oa<8pa<�qa<sa<ua<�  �  �ta<�ua<�ta<�sa<qa<ima<�ha<�ca<0^a<�Xa<[Sa<�Na<�Ka<Ja<�Ia<'Ka<�Ma<	Ra<QWa<e]a<�ca<�ia<�oa<�ta<�xa<�{a<�}a<�~a<�~a<!~a<}a<|a<�za<wza<Hza<�za<�{a<�}a<�a<f�a<��a<҆a<g�a<\�a<�a<�a<k�a<:�a<�}a<ya<ta<�na<|ja<�fa<�da<�ca<]da<�fa<�ia<�na<�ta<,{a<��a<҇a<��a<,�a<�a<��a<-�a<��a<�a<�a<ܗa<t�a<�a<M�a<�a<(�a<�a<a�a<@�a<��a<��a<�a<�a<��a<z�a<S�a<ǖa<��a<H�a<��a<�a<P|a<wwa<�sa<0qa<pa<�pa<�ra<�ua<�za<�a<�a<֋a<v�a<K�a<0�a<%�a<Ԟa<��a<6�a<J�a<��a<*�a<d�a<�a<�a<��a<��a<��a<Әa<}�a<�a<l�a<D�a<��a<�a<0�a<J�a<U�a<��a<Ҋa<�a<�~a<@ya<bta<�pa<�na<�ma<�na<�pa<Pta<ya<y~a<8�a<��a<�a<4�a<��a<��a<:�a<r�a<��a<@�a<n�a<��a<��a<H�a<5�a<Ϗa<�a<ɐa<�a<m�a<��a<��a<�a<ߕa<Y�a<��a<9�a<��a<�a<�}a<�wa<qa<Aka<4fa<�ba<V`a<�_a<\`a<qba<fa<qja<�oa<�ta<�ya<(~a<�a<<�a<��a<�a<D�a<̓a<Ɂa<�a<:}a<�za<Pya<xa<�wa<�wa<Ixa<vya<�za<�{a<I|a<�|a<�{a<�ya<Ewa<0sa<na<�ha<�ba<]\a<KVa<Qa<�La<�Ia<uHa<�Ha<JJa<OMa<�Qa<�Va<�\a<ba<~ga<!la<�oa<�ra</ta<�ta<[ta<^sa<�qa<-pa<ina<�la<la<�ka<la<ma<nna<Ipa<�qa<�sa<�  �  Usa<@ta<Uta<jsa<cqa<;na<&ja<rea<C`a<[a<]Va<]Ra<HOa<�Ma<AMa<�Na<\Qa<eUa<IZa<�_a<�ea<�ka<�pa<�ua<'ya<�{a<}a<p}a<"}a<|a<�za<)ya<�wa<wa<�va<�wa<�xa<�za<�|a<�a<`�a<�a<�a<E�a<��a<�a<�a<�a<Oa<�za<8va<�qa<�ma<Jja<ha<.ga<�ga<�ia<zma<-ra<�wa<r}a<��a<X�a<�a<�a<'�a<�a<#�a<#�a<h�a<ؖa<�a<i�a<�a<Ґa<��a<Аa<��a<<�a<E�a<e�a<��a<s�a<��a<ܜa<�a<y�a<��a<��a<�a<��a<X�a<<a<�za<wa<�ta<�sa<ta<va<lya<�}a<��a<(�a<��a<��a<%�a<��a<
�a<C�a<~�a<ʝa<_�a<[�a<B�a<A�a<��a<��a<C�a<P�a<B�a<��a<��a<��a<p�a<՜a<z�a<C�a<�a<��a<(�a<��a<��a<�a<r�a<C|a<�wa<>ta<�qa<3qa<�qa<7ta<�wa<�{a<��a<<�a<a�a<	�a<��a<��a<��a<n�a<�a<�a<'�a<�a<��a<��a<�a<Ռa<��a<��a<��a<�a<��a<R�a<�a<��a<ɔa<ߓa<��a<ގa<��a<��a<�a<�ya<�sa<ena<�ia<fa<�ca<ca<�ca<�ea<Bia<?ma<�qa<�va<({a<a<4�a<I�a<�a<��a<�a<�a<�a<�|a</za<�wa<�ua<�ta<6ta<Pta<%ua<zva<�wa<tya<�za<({a<�za<�ya<kwa<�sa<}oa<Pja<�da<�^a<7Ya<STa<6Pa<XMa<�Ka<La<�Ma<�Pa<�Ta<wYa<�^a<�ca<�ha<�la<Opa<�ra<�sa<�sa<�ra<tqa<doa<Fma<Gka<�ia<�ha<vha<�ha<�ia<Nka<Zma<�oa<�qa<�  �  ?qa<�ra<�sa<:sa<�qa<Toa<�ka<�ga<ca<�^a<Za<cVa<�Sa<"Ra<�Qa<$Sa<�Ua<IYa<�]a<2ca<{ha<�ma<xra<vva<jya<U{a<|a<�{a<�za<!ya<Mwa<sua<�sa<�ra<`ra<�ra<'ta<}va<	ya</|a<Ta<��a<�a<��a<�a<�a<��a<^�a<U�a<m}a<Eya<Fua<eqa<xna<�la<�ka<ula<�na<�qa<�ua<({a<��a<�a<l�a<׏a<��a<-�a<��a<�a<K�a<�a<֓a<��a<��a<�a<u�a<�a<E�a<^�a<Q�a<��a<�a<��a<+�a<��a<Λa<ܛa<��a<r�a<�a<&�a<g�a<��a<�a<�~a<d{a<.ya<>xa<�xa<�za<�}a<r�a<E�a<�a<�a<��a<Q�a<(�a<�a<��a<�a<śa<��a<5�a<��a<g�a<��a<�a<��a<юa<�a<ґa<�a<T�a<��a<��a<ݛa<t�a<֛a<�a<A�a<u�a<��a<މa<��a<�a<�{a<�xa<�va<�ua<�va<�xa<�{a<�a<H�a<�a<��a<��a<��a<8�a<o�a<u�a<c�a<ӕa<?�a<��a<��a<��a<��a<M�a<�a<5�a<��a<�a<4�a<F�a<V�a<͒a<s�a<]�a<�a<~�a<�a<��a<K�a<�|a<kwa<*ra<�ma<�ja<mha<�ga<Sha<+ja<ma<�pa<�ta<2ya<;}a<e�a<�a<N�a<��a<ăa<�a<�a<�|a<rya<[va<�sa<yqa<6pa<�oa<pa<:qa<�ra<�ta<�va<lxa<gya<�ya<Zya<�wa<�ta<�pa<�la<Mga<
ba<�\a<(Xa<�Ta<�Qa<�Pa<�Pa</Ra<�Ta<zXa<]a<�aa<Wfa<�ja<&na<�pa<dra<�ra<1ra<�pa<�na<@la<�ia<nga<�ea<$da<�ca<!da<�ea<pga<�ia<Xla<�na<�  �  �na<qa<�ra<�ra<<ra<�pa<�ma<cja<xfa<\ba<�^a<R[a<�Xa<uWa<>Wa<kXa<�Za<4^a<;ba<�fa<�ka<Cpa<\ta<qwa<�ya<�za<�za<�ya</xa<�ua<�sa<qa<�na<�ma<Bma<�ma<oa<Oqa<eta<xa<�{a<�a<܂a<��a<3�a<؇a<b�a<�a<��a<J�a<�|a<4ya<va<jsa<�qa<%qa<�qa<�sa<�va<�za<'a<)�a<�a<��a<z�a<]�a<5�a<�a<��a<(�a<��a<k�a<��a<��a<̈a<o�a<ˆa<�a<F�a<D�a<�a<=�a<c�a<S�a<��a<��a<;�a<ؚa<X�a<�a<~�a<��a<E�a<�a<��a<`�a<p~a<�}a<~a<�a<p�a<��a<�a<~�a<��a<��a<��a<��a<��a<��a<r�a<L�a<��a<��a<��a<��a<^�a<��a<[�a<a<�a<�a<��a<��a<��a<)�a<O�a<p�a<~�a<��a<o�a<x�a<��a<<�a<��a<r�a<Āa<�}a<�{a<2{a<�{a<�}a<�a<�a<��a<(�a<�a<��a<�a<�a<�a<K�a<��a<�a<�a<ٌa<��a<��a<|�a<.�a<��a<-�a<b�a<v�a<�a<Ƌa<Z�a<��a<	�a<��a<�a<.�a<c�a<��a<'�a<V�a<Z{a<�va<�ra<�oa<�ma<�la<�ma<oa<�qa<�ta<�xa<!|a<ra<�a<��a<W�a<��a<g�a<�a<�|a<ya<pua<�qa<�na<sla<�ja<�ja<�ja<-la<Ana<�pa<Esa<�ua<�wa<�xa<�xa<�wa<�ua<�ra<�na<ija<�ea<aa<]a<Ya<)Wa<�Ua<Va<IWa<�Ya<]a<�`a<�da<�ha<�la<koa<Oqa<+ra<�qa<�pa<tna<�ka<�ha<�ea<�ba<o`a<_a<�^a<_a<d`a<�ba<�ea<�ha<�ka<�  �  �ka<oa<:qa<�ra<�ra<�qa<�oa<ma<ja<tfa<7ca<k`a<1^a< ]a<�\a<^a<`a<@ca<�fa<�ja<#oa<�ra<&va<xa<"za<Uza<sya<�wa<;ua<xra<(oa<dla<�ia<;ha<�ga<�ga<�ia<la<�oa<�sa<xa<p|a<G�a<ƃa<@�a<�a< �a<Y�a<��a<K�a<��a<q}a<�za<�xa<Ewa<�va<rwa<Gya<�{a<�a<t�a<��a<+�a<�a<�a<)�a<h�a<�a<��a<��a<�a<��a<#�a<I�a<��a<�a<�a<o�a<Ђa<-�a<]�a<ʋa<Ϗa<W�a<��a<�a<��a<9�a<R�a<��a<�a<�a<<�a<��a<��a<��a<�a<5�a<��a<�a<��a<��a<5�a<,�a<��a<��a<��a<J�a<��a<f�a<��a<��a<d�a<��a<�a<��a<��a<d�a<��a<'�a<��a<
�a<�a<��a<F�a<[�a<I�a<&�a<F�a<�a<��a<t�a<:�a<ِa<Όa< �a<߅a<*�a<��a<Ӏa<��a<�a<��a<y�a<��a<��a<��a<S�a< �a<�a<q�a<וa<k�a< �a<��a<|�a<�a<��a<
a<�}a<�|a<�}a<a<��a<��a<�a<C�a<��a<G�a<��a< �a<�a<ێa<�a<(�a<�a<�a<�{a<xa<Cua<nsa<�ra<sa<^ta<�va<0ya<b|a<Ea<��a<��a<~�a<��a<�a<��a<q}a<�ya<]ua<�pa<ma<lia<�fa<9ea<�da<tea<ga<�ia<Sla<�oa<�ra<@ua<wa<!xa<)xa<�va<�ta<Hqa<�ma<�ia<�ea<ba<�^a<�\a<�[a<�[a<�\a<�^a<�aa<�da<�ha<�ka<�na<�pa<�qa<ra<�pa<�na<�ka<|ha<�da<�`a<�]a<[a<�Ya<�Xa<zYa<�Za<�]a<�`a<�da<�ha<�  �  ?ia<"ma<pa<ra<sa<sa<�qa<�oa<kma<�ja<�ga<Zea<�ca<�ba<�ba<�ca<kea<ha<gka<�na<Wra<tua<xa<�ya<2za<�ya<xa<�ua<era<�na< ka<�ga<�da<�ba<�aa<Bba<�ca<�fa<�ja<oa<ta<ya<�}a<�a<S�a<��a<ƈa<�a<�a<J�a<4�a<�a<�a<�}a<�|a<�|a<0}a<�~a<$�a<U�a<�a<��a<.�a<R�a<��a<�a<&�a<=�a<L�a<]�a<��a<ψa<Ȅa<Z�a<E~a<K|a<`{a<�{a<C}a<�a<��a<��a<�a<g�a<q�a<��a<�a<0�a<U�a<p�a<��a<�a<�a<-�a<J�a<�a<��a< �a<_�a<��a<��a<h�a<��a<��a<u�a<՚a<J�a<��a<�a<K�a<��a<�a<�a<��a<N�a<��a<��a<�~a<�}a<z~a<�a<�a<e�a<p�a<��a<��a<Y�a<��a<��a<`�a<��a<��a<�a<1�a<�a<ʍa<ϊa<��a<8�a<��a<�a<L�a<^�a<�a<��a<Ғa<K�a<5�a<#�a<�a<Ȗa<��a<W�a<J�a<�a<U�a<�a<s|a<�ya<�wa<Bwa<�wa<�ya<�|a<�a<�a<�a<��a<��a<��a<��a<��a<j�a<4�a<&�a<��a<�a<h�a<+}a<�za<"ya<fxa<�xa<�ya<k{a<�}a<�a<G�a<#�a<6�a<B�a<I�a<7�a<%a< {a<qva<�qa<�la<#ha<'da<Paa<�_a<(_a<�_a<�aa<�da<ha<�ka<�oa<sa<�ua<lwa<xa<�wa<Ova<�sa<�pa<�ma<#ja<�fa<"da<Zba<Vaa<Zaa</ba<�ca<nfa<Eia<la<�na<�pa< ra<\ra<�qa<�oa<�la</ia<�da<�`a<X\a<�Xa<�Ua<�Sa<!Sa<�Sa<�Ua<�Xa<6\a<v`a<�da<�  �  �fa<%ka<�na<�qa<zsa<ta<�sa<�ra<�pa<Zna<&la<Cja<�ha<�ga<�ga<�ha<�ja<�la<�oa<tra<[ua<�wa<�ya<�za<]za< ya<�va<�sa<�oa<Uka<-ga<ca<�_a<�]a<�\a<�\a<�^a<�aa<�ea<�ja<qpa<va<�{a<U�a<w�a<u�a<s�a<.�a<�a<*�a<�a<υa<�a<ڂa<ҁa<��a<c�a<уa<@�a<��a<��a<�a<�a<d�a<��a<��a<�a<q�a<��a<�a<��a<6�a<��a<�|a<Rya<wa<va<kva<#xa<{a<�~a<��a<��a<��a<M�a<0�a<K�a<E�a<:�a<��a<ۚa<�a<��a<M�a<��a<7�a<��a<E�a<y�a<��a<��a<��a<H�a<a<'�a<��a<k�a<+�a<��a<E�a<��a<��a<��a<Їa< �a<�~a<�{a<mya<�xa<*ya<	{a<~a< �a<��a<[�a<2�a<[�a<חa<R�a<��a<�a< �a<��a<M�a<��a<�a<��a<a<J�a<�a<�a<{�a< �a<J�a<��a<ؕa<��a<��a<�a</�a<>�a<2�a<@�a<��a<u�a<��a<�{a<�wa<rta<�ra<�qa<�ra<�ta<�wa<�{a<`�a<�a<F�a<Ռa<Ïa<��a<>�a<��a<$�a<�a<�a<�a<�a<<�a<�a<J~a<�}a<�}a<�~a<�a<��a<w�a<5�a<5�a<��a<�a<8�a<k�a<t}a<�xa<vsa<�ma<vha<Xca<4_a<\a<@Za<�Ya<�Za<�\a<`a<6da<oha<�la<�pa<=ta<�va<2xa<�xa<�wa<9va<�sa<qa<Bna<}ka<Ria<dga<�fa<rfa<Yga<�ha<�ja<ma<>oa<gqa<�ra<Bsa<�ra<Aqa<�na<ka<�fa<�aa<�\a<Xa<�Sa<�Pa<�Na<�Ma<�Na<�Pa<�Sa<�Wa<�\a<�aa<�  �  ada<oia<�ma<[qa<�sa<�ta<2ua<�ta<Tsa<�qa<�oa<"na<�la<Nla<�la<$ma<�na<�pa<sa<�ua<xa<�ya< {a<7{a<zza<�xa<�ua<�qa<:ma<\ha<�ca<H_a<�[a<.Ya<�Wa<KXa<'Za<u]a<�aa<Ega<7ma<msa<jya<�~a<��a<Q�a<��a<E�a<��a<��a<s�a<%�a<�a<ǆa<$�a<?�a<��a<*�a<5�a<��a<X�a<
�a<��a<4�a<&�a<
�a<�a<��a<8�a<�a<+�a<�a<}a<�xa<ua<�ra<iqa<�qa<�sa<�va<{a<�a<��a<�a<Q�a<�a<��a<W�a<ǜa<E�a<˜a<��a<��a<��a<Еa<A�a<�a<�a< �a<�a<u�a<q�a<��a<��a<R�a<4�a<\�a<f�a<t�a<D�a<�a<A�a<�a<n�a<La<�za<:wa<�ta<�sa<�ta<�va<za<G~a<:�a<��a<ݍa<��a<Ŗa<��a<��a<�a<a<Лa<�a<�a<��a<��a<�a<̐a<��a<��a<��a<��a<ǔa<��a<��a<��a<1�a<��a<M�a<��a<��a<\�a<!�a<|�a<�|a<�wa<fsa<�oa<�ma<Kma<3na<�pa<ta<Hxa<&}a<?�a<�a<_�a<�a<_�a<��a<Œa<�a<\�a<�a<I�a<��a<)�a<"�a<قa<+�a<��a<��a<Ƀa<�a<s�a<��a<�a<��a<`�a<(�a<��a<|a<�va<�pa<�ja<�da<�_a<�Za<�Wa<�Ua</Ua<KVa<�Xa<R\a<�`a<hea<Vja<�na<�ra<.va<Dxa<*ya<#ya<(xa<zva<ta<�qa<Uoa<[ma<�ka<6ka<�ja<�ka<�la<vna<Epa<ra<�sa<=ta<2ta<sa<�pa<�ma<^ia<nda< _a<~Ya<XTa<�Oa<PLa<�Ia<&Ia<�Ia<!La<�Oa<Ta<CYa<�^a<�  �  �ba<Lha<ma<qa<�sa<�ua<zva<va<Wua< ta<�ra<Aqa<Fpa<�oa<�oa<�pa<�qa<�sa<�ua<�wa<�ya<C{a<,|a<�{a<�za<xa<�ta<kpa<hka<<fa<�`a<<\a<EXa<�Ua<�Ta<�Ta<�Va<�Ya<�^a<ada<�ja<rqa<�wa<�}a<قa<0�a<!�a<5�a<�a<�a<��a<ȋa<�a<�a<��a<��a<B�a<��a<_�a<��a<�a<E�a<6�a<��a<)�a<|�a<�a<�a<N�a<s�a<8�a<�a<Aza<�ua<�qa<oa<�ma<Vna<6pa<bsa<xa<]}a<Z�a<?�a<�a<�a<�a<`�a<G�a<b�a<0�a<h�a<	�a<��a<�a<y�a<��a<$�a<d�a<P�a<��a<g�a<�a<��a<͞a<��a<�a<��a<3�a<y�a<�a<��a<݇a<��a<O|a<twa<�sa<jqa<vpa<"qa<+sa<�va<E{a<��a<�a<�a<��a<��a<��a<(�a<��a<
�a<C�a<�a<]�a<��a<��a<D�a<4�a<ʓa<�a<Дa<�a<��a<�a<d�a<�a<^�a<H�a<d�a<1�a<"�a<�a<O�a<\�a<Jza<�ta<�oa<�la<tja<�ia<�ja<ma<�pa<cua<�za<D�a<x�a<g�a<#�a<>�a<�a<��a<N�a<��a<#�a<�a<��a<P�a<��a<,�a<x�a<x�a<Ӆa<φa<̇a<��a<Q�a<f�a<��a<҆a<�a<�a<){a<7ua<�na<mha<�aa<N\a<pWa<$Ta<%Ra<�Qa<�Ra<LUa<7Ya<�]a<<ca<ha<�ma< ra<�ua<Lxa<�ya<?za<�ya<Gxa<pva<�ta<tra<�pa<?oa<wna<[na<�na<�oa<kqa<�ra<0ta<ua<�ua<�ta<Tsa<�pa<�la<Pha<�ba<�\a<Wa<\Qa<�La<�Ha<�Fa<�Ea<zFa<�Ha<CLa<Qa<�Va<�\a<�  �  eaa<Uga<�la<�pa<ta<va<wa<.wa<�va<�ua<Nta<sa<^ra<�qa<ra<�ra<�sa<ua<�wa<rya<8{a<I|a<�|a<'|a<�za<�wa<.ta<moa<&ja<�da<\_a<kZa<jVa<�Sa<3Ra<qRa<�Ta<Xa<�\a<�ba<<ia<pa<�va<}a<��a<�a<p�a<��a<�a<W�a<�a<Q�a<{�a<�a<��a<ˋa<|�a<��a<h�a<M�a<��a<��a<s�a<o�a<��a<ϗa<ڕa<��a<��a<c�a<�a<~a<�xa<�sa<�oa<�la<�ka<�ka<na<�qa<%va<�{a<��a<��a<�a<t�a<ޗa<g�a<��a<�a<)�a<��a<��a<"�a<��a<��a<��a<^�a<��a<g�a<x�a<��a<��a<�a<��a<?�a<��a<�a<��a<�a<�a<]�a<d�a<X�a<�za<�ua<�qa<oa<na<�na<-qa<�ta<�ya<a<��a<�a<��a<x�a<i�a<S�a<�a<��a<]�a<�a<�a<;�a<��a<\�a<Y�a<	�a<"�a<��a<җa<>�a<��a<��a<$�a<�a<��a<w�a<��a<��a<�a<�a<�~a<�xa<�ra<na<uja<ha<pga<�ha<!ka<�na<�sa<*ya<�~a<_�a<��a<ˍa<�a<:�a<&�a<�a<2�a<��a<u�a<>�a<P�a<��a<d�a<��a<��a<ۇa<d�a<V�a< �a<��a<A�a<5�a<%�a<��a<�a<mza<'ta<�ma<�fa<j`a<eZa<�Ua<�Qa<�Oa<fOa<�Pa<pSa<ZWa<P\a<�aa<>ga<�la<�qa<Xua<Sxa<za<�za<�za<�ya<�wa<va<ta<�ra<Yqa<�pa<�pa<qa<�qa<sa<Vta<�ua<6va<Hva<Wua<�sa<�pa<gla<bga<�aa<�[a<jUa<�Oa<�Ja<�Fa<EDa<TCa<%Da<�Fa<`Ja<cOa<Ua<@[a<�  �  Faa<ga<[la<�pa<ta<?va<Uwa<lwa<�va<-va<�ta<�sa<sa<�ra<�ra<Qsa<�ta<3va<3xa<�ya<y{a<�|a<�|a<S|a<}za<�wa<�sa<'oa<�ia<*da<�^a<�Ya<�Ua<�Ra<�Qa<�Qa<�Sa<HWa<�[a<%ba<�ha<�oa<�va<�|a<j�a<цa<x�a<׌a<�a<��a<o�a<��a<*�a<��a<?�a<��a<=�a<N�a<1�a<�a<G�a<%�a<��a<��a<֘a<חa<��a<��a<E�a<$�a<��a<}a<xa<�ra<�na<la< ka<Yka<:ma<�pa<Xua<,{a<3�a<Ǉa<��a<)�a<��a<9�a<ŝa<�a<g�a<��a<�a<Μa<N�a<I�a<D�a<.�a<C�a<�a<3�a<��a<6�a<g�a<4�a<r�a<��a<�a<��a<ߖa<֑a<8�a<�a<�a<�ya<�ta< qa<Wna<�ma<
na<bpa<�sa<�xa<t~a<��a<��a<C�a<F�a<+�a<H�a<.�a<�a<��a<ǝa<��a<�a<A�a<�a<
�a<ؖa<Ėa<��a<��a<�a<�a<��a<]�a<�a<ٚa<Q�a<ʔa<S�a<ϊa<߄a<J~a<xa<#ra<Nma<�ia<rga<�fa<�ga<Yja<	na<&sa<�xa<�~a<-�a<V�a<��a<ސa<B�a<W�a<G�a<q�a<�a<"�a<�a<�a<=�a<�a<s�a<"�a<��a<�a<�a<��a<Њa<{�a<g�a<.�a<ăa<�a< za<�sa<Yma<3fa<�_a<�Ya<�Ta<Qa<3Oa<�Na<�Oa<�Ra<�Va<�[a<aa<ga<Jla<5qa<1ua<%xa<'za<�za<�za<�ya<qxa<�va<�ta<asa<�qa<�qa<:qa<�qa<�ra<�sa<�ta<�ua<tva<zva<�ua<�sa<?pa<@la<ga<faa<$[a<�Ta<Oa<�Ia<Fa<~Ca<�Ba<cCa<�Ea<�Ia<�Na<~Ta<�Za<�  �  eaa<Uga<�la<�pa<ta<va<wa<.wa<�va<�ua<Nta<sa<^ra<�qa<ra<�ra<�sa<ua<�wa<rya<8{a<I|a<�|a<'|a<�za<�wa<.ta<moa<&ja<�da<\_a<kZa<jVa<�Sa<3Ra<qRa<�Ta<Xa<�\a<�ba<<ia<pa<�va<}a<��a<�a<p�a<��a<�a<W�a<�a<Q�a<{�a<�a<��a<ˋa<|�a<��a<h�a<M�a<��a<��a<s�a<o�a<��a<ϗa<ڕa<��a<��a<c�a<�a<~a<�xa<�sa<�oa<�la<�ka<�ka<na<�qa<%va<�{a<��a<��a<�a<t�a<ޗa<g�a<��a<�a<)�a<��a<��a<"�a<��a<��a<��a<^�a<��a<g�a<x�a<��a<��a<�a<��a<?�a<��a<�a<��a<�a<�a<]�a<d�a<X�a<�za<�ua<�qa<oa<na<�na<-qa<�ta<�ya<a<��a<�a<��a<x�a<i�a<S�a<�a<��a<]�a<�a<�a<;�a<��a<\�a<Y�a<	�a<"�a<��a<җa<>�a<��a<��a<$�a<�a<��a<w�a<��a<��a<�a<�a<�~a<�xa<�ra<na<uja<ha<pga<�ha<!ka<�na<�sa<*ya<�~a<_�a<��a<ˍa<�a<:�a<&�a<�a<2�a<��a<u�a<>�a<P�a<��a<d�a<��a<��a<ۇa<d�a<V�a< �a<��a<A�a<5�a<%�a<��a<�a<mza<'ta<�ma<�fa<j`a<eZa<�Ua<�Qa<�Oa<fOa<�Pa<pSa<ZWa<P\a<�aa<>ga<�la<�qa<Xua<Sxa<za<�za<�za<�ya<�wa<va<ta<�ra<Yqa<�pa<�pa<qa<�qa<sa<Vta<�ua<6va<Hva<Wua<�sa<�pa<gla<bga<�aa<�[a<jUa<�Oa<�Ja<�Fa<EDa<TCa<%Da<�Fa<`Ja<cOa<Ua<@[a<�  �  �ba<Lha<ma<qa<�sa<�ua<zva<va<Wua< ta<�ra<Aqa<Fpa<�oa<�oa<�pa<�qa<�sa<�ua<�wa<�ya<C{a<,|a<�{a<�za<xa<�ta<kpa<hka<<fa<�`a<<\a<EXa<�Ua<�Ta<�Ta<�Va<�Ya<�^a<ada<�ja<rqa<�wa<�}a<قa<0�a<!�a<5�a<�a<�a<��a<ȋa<�a<�a<��a<��a<B�a<��a<_�a<��a<�a<E�a<6�a<��a<)�a<|�a<�a<�a<N�a<s�a<8�a<�a<Aza<�ua<�qa<oa<�ma<Vna<6pa<bsa<xa<]}a<Z�a<?�a<�a<�a<�a<`�a<G�a<b�a<0�a<h�a<	�a<��a<�a<y�a<��a<$�a<d�a<P�a<��a<g�a<�a<��a<͞a<��a<�a<��a<3�a<y�a<�a<��a<݇a<��a<O|a<twa<�sa<jqa<vpa<"qa<+sa<�va<E{a<��a<�a<�a<��a<��a<��a<(�a<��a<
�a<C�a<�a<]�a<��a<��a<D�a<4�a<ʓa<�a<Дa<�a<��a<�a<d�a<�a<^�a<H�a<d�a<1�a<"�a<�a<O�a<\�a<Jza<�ta<�oa<�la<tja<�ia<�ja<ma<�pa<cua<�za<D�a<x�a<g�a<#�a<>�a<�a<��a<N�a<��a<#�a<�a<��a<P�a<��a<,�a<x�a<x�a<Ӆa<φa<̇a<��a<Q�a<f�a<��a<҆a<�a<�a<){a<7ua<�na<mha<�aa<N\a<pWa<$Ta<%Ra<�Qa<�Ra<LUa<7Ya<�]a<<ca<ha<�ma< ra<�ua<Lxa<�ya<?za<�ya<Gxa<pva<�ta<tra<�pa<?oa<wna<[na<�na<�oa<kqa<�ra<0ta<ua<�ua<�ta<Tsa<�pa<�la<Pha<�ba<�\a<Wa<\Qa<�La<�Ha<�Fa<�Ea<zFa<�Ha<CLa<Qa<�Va<�\a<�  �  ada<oia<�ma<[qa<�sa<�ta<2ua<�ta<Tsa<�qa<�oa<"na<�la<Nla<�la<$ma<�na<�pa<sa<�ua<xa<�ya< {a<7{a<zza<�xa<�ua<�qa<:ma<\ha<�ca<H_a<�[a<.Ya<�Wa<KXa<'Za<u]a<�aa<Ega<7ma<msa<jya<�~a<��a<Q�a<��a<E�a<��a<��a<s�a<%�a<�a<ǆa<$�a<?�a<��a<*�a<5�a<��a<X�a<
�a<��a<4�a<&�a<
�a<�a<��a<8�a<�a<+�a<�a<}a<�xa<ua<�ra<iqa<�qa<�sa<�va<{a<�a<��a<�a<Q�a<�a<��a<W�a<ǜa<E�a<˜a<��a<��a<��a<Еa<A�a<�a<�a< �a<�a<u�a<q�a<��a<��a<R�a<4�a<\�a<f�a<t�a<D�a<�a<A�a<�a<n�a<La<�za<:wa<�ta<�sa<�ta<�va<za<G~a<:�a<��a<ݍa<��a<Ŗa<��a<��a<�a<a<Лa<�a<�a<��a<��a<�a<̐a<��a<��a<��a<��a<ǔa<��a<��a<��a<1�a<��a<M�a<��a<��a<\�a<!�a<|�a<�|a<�wa<fsa<�oa<�ma<Kma<3na<�pa<ta<Hxa<&}a<?�a<�a<_�a<�a<_�a<��a<Œa<�a<\�a<�a<I�a<��a<)�a<"�a<قa<+�a<��a<��a<Ƀa<�a<s�a<��a<�a<��a<`�a<(�a<��a<|a<�va<�pa<�ja<�da<�_a<�Za<�Wa<�Ua</Ua<KVa<�Xa<R\a<�`a<hea<Vja<�na<�ra<.va<Dxa<*ya<#ya<(xa<zva<ta<�qa<Uoa<[ma<�ka<6ka<�ja<�ka<�la<vna<Epa<ra<�sa<=ta<2ta<sa<�pa<�ma<^ia<nda< _a<~Ya<XTa<�Oa<PLa<�Ia<&Ia<�Ia<!La<�Oa<Ta<CYa<�^a<�  �  �fa<%ka<�na<�qa<zsa<ta<�sa<�ra<�pa<Zna<&la<Cja<�ha<�ga<�ga<�ha<�ja<�la<�oa<tra<[ua<�wa<�ya<�za<]za< ya<�va<�sa<�oa<Uka<-ga<ca<�_a<�]a<�\a<�\a<�^a<�aa<�ea<�ja<qpa<va<�{a<U�a<w�a<u�a<s�a<.�a<�a<*�a<�a<υa<�a<ڂa<ҁa<��a<c�a<уa<@�a<��a<��a<�a<�a<d�a<��a<��a<�a<q�a<��a<�a<��a<6�a<��a<�|a<Rya<wa<va<kva<#xa<{a<�~a<��a<��a<��a<M�a<0�a<K�a<E�a<:�a<��a<ۚa<�a<��a<M�a<��a<7�a<��a<E�a<y�a<��a<��a<��a<H�a<a<'�a<��a<k�a<+�a<��a<E�a<��a<��a<��a<Їa< �a<�~a<�{a<mya<�xa<*ya<	{a<~a< �a<��a<[�a<2�a<[�a<חa<R�a<��a<�a< �a<��a<M�a<��a<�a<��a<a<J�a<�a<�a<{�a< �a<J�a<��a<ؕa<��a<��a<�a</�a<>�a<2�a<@�a<��a<u�a<��a<�{a<�wa<rta<�ra<�qa<�ra<�ta<�wa<�{a<`�a<�a<F�a<Ռa<Ïa<��a<>�a<��a<$�a<�a<�a<�a<�a<<�a<�a<J~a<�}a<�}a<�~a<�a<��a<w�a<5�a<5�a<��a<�a<8�a<k�a<t}a<�xa<vsa<�ma<vha<Xca<4_a<\a<@Za<�Ya<�Za<�\a<`a<6da<oha<�la<�pa<=ta<�va<2xa<�xa<�wa<9va<�sa<qa<Bna<}ka<Ria<dga<�fa<rfa<Yga<�ha<�ja<ma<>oa<gqa<�ra<Bsa<�ra<Aqa<�na<ka<�fa<�aa<�\a<Xa<�Sa<�Pa<�Na<�Ma<�Na<�Pa<�Sa<�Wa<�\a<�aa<�  �  ?ia<"ma<pa<ra<sa<sa<�qa<�oa<kma<�ja<�ga<Zea<�ca<�ba<�ba<�ca<kea<ha<gka<�na<Wra<tua<xa<�ya<2za<�ya<xa<�ua<era<�na< ka<�ga<�da<�ba<�aa<Bba<�ca<�fa<�ja<oa<ta<ya<�}a<�a<S�a<��a<ƈa<�a<�a<J�a<4�a<�a<�a<�}a<�|a<�|a<0}a<�~a<$�a<U�a<�a<��a<.�a<R�a<��a<�a<&�a<=�a<L�a<]�a<��a<ψa<Ȅa<Z�a<E~a<K|a<`{a<�{a<C}a<�a<��a<��a<�a<g�a<q�a<��a<�a<0�a<U�a<p�a<��a<�a<�a<-�a<J�a<�a<��a< �a<_�a<��a<��a<h�a<��a<��a<u�a<՚a<J�a<��a<�a<K�a<��a<�a<�a<��a<N�a<��a<��a<�~a<�}a<z~a<�a<�a<e�a<p�a<��a<��a<Y�a<��a<��a<`�a<��a<��a<�a<1�a<�a<ʍa<ϊa<��a<8�a<��a<�a<L�a<^�a<�a<��a<Ғa<K�a<5�a<#�a<�a<Ȗa<��a<W�a<J�a<�a<U�a<�a<s|a<�ya<�wa<Bwa<�wa<�ya<�|a<�a<�a<�a<��a<��a<��a<��a<��a<j�a<4�a<&�a<��a<�a<h�a<+}a<�za<"ya<fxa<�xa<�ya<k{a<�}a<�a<G�a<#�a<6�a<B�a<I�a<7�a<%a< {a<qva<�qa<�la<#ha<'da<Paa<�_a<(_a<�_a<�aa<�da<ha<�ka<�oa<sa<�ua<lwa<xa<�wa<Ova<�sa<�pa<�ma<#ja<�fa<"da<Zba<Vaa<Zaa</ba<�ca<nfa<Eia<la<�na<�pa< ra<\ra<�qa<�oa<�la</ia<�da<�`a<X\a<�Xa<�Ua<�Sa<!Sa<�Sa<�Ua<�Xa<6\a<v`a<�da<�  �  �ka<oa<:qa<�ra<�ra<�qa<�oa<ma<ja<tfa<7ca<k`a<1^a< ]a<�\a<^a<`a<@ca<�fa<�ja<#oa<�ra<&va<xa<"za<Uza<sya<�wa<;ua<xra<(oa<dla<�ia<;ha<�ga<�ga<�ia<la<�oa<�sa<xa<p|a<G�a<ƃa<@�a<�a< �a<Y�a<��a<K�a<��a<q}a<�za<�xa<Ewa<�va<rwa<Gya<�{a<�a<t�a<��a<+�a<�a<�a<)�a<h�a<�a<��a<��a<�a<��a<#�a<I�a<��a<�a<�a<o�a<Ђa<-�a<]�a<ʋa<Ϗa<W�a<��a<�a<��a<9�a<R�a<��a<�a<�a<<�a<��a<��a<��a<�a<5�a<��a<�a<��a<��a<5�a<,�a<��a<��a<��a<J�a<��a<f�a<��a<��a<d�a<��a<�a<��a<��a<d�a<��a<'�a<��a<
�a<�a<��a<F�a<[�a<I�a<&�a<F�a<�a<��a<t�a<:�a<ِa<Όa< �a<߅a<*�a<��a<Ӏa<��a<�a<��a<y�a<��a<��a<��a<S�a< �a<�a<q�a<וa<k�a< �a<��a<|�a<�a<��a<
a<�}a<�|a<�}a<a<��a<��a<�a<C�a<��a<G�a<��a< �a<�a<ێa<�a<(�a<�a<�a<�{a<xa<Cua<nsa<�ra<sa<^ta<�va<0ya<b|a<Ea<��a<��a<~�a<��a<�a<��a<q}a<�ya<]ua<�pa<ma<lia<�fa<9ea<�da<tea<ga<�ia<Sla<�oa<�ra<@ua<wa<!xa<)xa<�va<�ta<Hqa<�ma<�ia<�ea<ba<�^a<�\a<�[a<�[a<�\a<�^a<�aa<�da<�ha<�ka<�na<�pa<�qa<ra<�pa<�na<�ka<|ha<�da<�`a<�]a<[a<�Ya<�Xa<zYa<�Za<�]a<�`a<�da<�ha<�  �  �na<qa<�ra<�ra<<ra<�pa<�ma<cja<xfa<\ba<�^a<R[a<�Xa<uWa<>Wa<kXa<�Za<4^a<;ba<�fa<�ka<Cpa<\ta<qwa<�ya<�za<�za<�ya</xa<�ua<�sa<qa<�na<�ma<Bma<�ma<oa<Oqa<eta<xa<�{a<�a<܂a<��a<3�a<؇a<b�a<�a<��a<J�a<�|a<4ya<va<jsa<�qa<%qa<�qa<�sa<�va<�za<'a<)�a<�a<��a<z�a<]�a<5�a<�a<��a<(�a<��a<k�a<��a<��a<̈a<o�a<ˆa<�a<F�a<D�a<�a<=�a<c�a<S�a<��a<��a<;�a<ؚa<X�a<�a<~�a<��a<E�a<�a<��a<`�a<p~a<�}a<~a<�a<p�a<��a<�a<~�a<��a<��a<��a<��a<��a<��a<r�a<L�a<��a<��a<��a<��a<^�a<��a<[�a<a<�a<�a<��a<��a<��a<)�a<O�a<p�a<~�a<��a<o�a<x�a<��a<<�a<��a<r�a<Āa<�}a<�{a<2{a<�{a<�}a<�a<�a<��a<(�a<�a<��a<�a<�a<�a<K�a<��a<�a<�a<ٌa<��a<��a<|�a<.�a<��a<-�a<b�a<v�a<�a<Ƌa<Z�a<��a<	�a<��a<�a<.�a<c�a<��a<'�a<V�a<Z{a<�va<�ra<�oa<�ma<�la<�ma<oa<�qa<�ta<�xa<!|a<ra<�a<��a<W�a<��a<g�a<�a<�|a<ya<pua<�qa<�na<sla<�ja<�ja<�ja<-la<Ana<�pa<Esa<�ua<�wa<�xa<�xa<�wa<�ua<�ra<�na<ija<�ea<aa<]a<Ya<)Wa<�Ua<Va<IWa<�Ya<]a<�`a<�da<�ha<�la<koa<Oqa<+ra<�qa<�pa<tna<�ka<�ha<�ea<�ba<o`a<_a<�^a<_a<d`a<�ba<�ea<�ha<�ka<�  �  ?qa<�ra<�sa<:sa<�qa<Toa<�ka<�ga<ca<�^a<Za<cVa<�Sa<"Ra<�Qa<$Sa<�Ua<IYa<�]a<2ca<{ha<�ma<xra<vva<jya<U{a<|a<�{a<�za<!ya<Mwa<sua<�sa<�ra<`ra<�ra<'ta<}va<	ya</|a<Ta<��a<�a<��a<�a<�a<��a<^�a<U�a<m}a<Eya<Fua<eqa<xna<�la<�ka<ula<�na<�qa<�ua<({a<��a<�a<l�a<׏a<��a<-�a<��a<�a<K�a<�a<֓a<��a<��a<�a<u�a<�a<E�a<^�a<Q�a<��a<�a<��a<+�a<��a<Λa<ܛa<��a<r�a<�a<&�a<g�a<��a<�a<�~a<d{a<.ya<>xa<�xa<�za<�}a<r�a<E�a<�a<�a<��a<Q�a<(�a<�a<��a<�a<śa<��a<5�a<��a<g�a<��a<�a<��a<юa<�a<ґa<�a<T�a<��a<��a<ݛa<t�a<֛a<�a<A�a<u�a<��a<މa<��a<�a<�{a<�xa<�va<�ua<�va<�xa<�{a<�a<H�a<�a<��a<��a<��a<8�a<o�a<u�a<c�a<ӕa<?�a<��a<��a<��a<��a<M�a<�a<5�a<��a<�a<4�a<F�a<V�a<͒a<s�a<]�a<�a<~�a<�a<��a<K�a<�|a<kwa<*ra<�ma<�ja<mha<�ga<Sha<+ja<ma<�pa<�ta<2ya<;}a<e�a<�a<N�a<��a<ăa<�a<�a<�|a<rya<[va<�sa<yqa<6pa<�oa<pa<:qa<�ra<�ta<�va<lxa<gya<�ya<Zya<�wa<�ta<�pa<�la<Mga<
ba<�\a<(Xa<�Ta<�Qa<�Pa<�Pa</Ra<�Ta<zXa<]a<�aa<Wfa<�ja<&na<�pa<dra<�ra<1ra<�pa<�na<@la<�ia<nga<�ea<$da<�ca<!da<�ea<pga<�ia<Xla<�na<�  �  Usa<@ta<Uta<jsa<cqa<;na<&ja<rea<C`a<[a<]Va<]Ra<HOa<�Ma<AMa<�Na<\Qa<eUa<IZa<�_a<�ea<�ka<�pa<�ua<'ya<�{a<}a<p}a<"}a<|a<�za<)ya<�wa<wa<�va<�wa<�xa<�za<�|a<�a<`�a<�a<�a<E�a<��a<�a<�a<�a<Oa<�za<8va<�qa<�ma<Jja<ha<.ga<�ga<�ia<zma<-ra<�wa<r}a<��a<X�a<�a<�a<'�a<�a<#�a<#�a<h�a<ؖa<�a<i�a<�a<Ґa<��a<Аa<��a<<�a<E�a<e�a<��a<s�a<��a<ܜa<�a<y�a<��a<��a<�a<��a<X�a<<a<�za<wa<�ta<�sa<ta<va<lya<�}a<��a<(�a<��a<��a<%�a<��a<
�a<C�a<~�a<ʝa<_�a<[�a<B�a<A�a<��a<��a<C�a<P�a<B�a<��a<��a<��a<p�a<՜a<z�a<C�a<�a<��a<(�a<��a<��a<�a<r�a<C|a<�wa<>ta<�qa<3qa<�qa<7ta<�wa<�{a<��a<<�a<a�a<	�a<��a<��a<��a<n�a<�a<�a<'�a<�a<��a<��a<�a<Ռa<��a<��a<��a<�a<��a<R�a<�a<��a<ɔa<ߓa<��a<ގa<��a<��a<�a<�ya<�sa<ena<�ia<fa<�ca<ca<�ca<�ea<Bia<?ma<�qa<�va<({a<a<4�a<I�a<�a<��a<�a<�a<�a<�|a</za<�wa<�ua<�ta<6ta<Pta<%ua<zva<�wa<tya<�za<({a<�za<�ya<kwa<�sa<}oa<Pja<�da<�^a<7Ya<STa<6Pa<XMa<�Ka<La<�Ma<�Pa<�Ta<wYa<�^a<�ca<�ha<�la<Opa<�ra<�sa<�sa<�ra<tqa<doa<Fma<Gka<�ia<�ha<vha<�ha<�ia<Nka<Zma<�oa<�qa<�  �  �ta<�ua<�ta<�sa<qa<ima<�ha<�ca<0^a<�Xa<[Sa<�Na<�Ka<Ja<�Ia<'Ka<�Ma<	Ra<QWa<e]a<�ca<�ia<�oa<�ta<�xa<�{a<�}a<�~a<�~a<!~a<}a<|a<�za<wza<Hza<�za<�{a<�}a<�a<f�a<��a<҆a<g�a<\�a<�a<�a<k�a<:�a<�}a<ya<ta<�na<|ja<�fa<�da<�ca<]da<�fa<�ia<�na<�ta<,{a<��a<҇a<��a<,�a<�a<��a<-�a<��a<�a<�a<ܗa<t�a<�a<M�a<�a<(�a<�a<a�a<@�a<��a<��a<�a<�a<��a<z�a<S�a<ǖa<��a<H�a<��a<�a<P|a<wwa<�sa<0qa<pa<�pa<�ra<�ua<�za<�a<�a<֋a<v�a<K�a<0�a<%�a<Ԟa<��a<6�a<J�a<��a<*�a<d�a<�a<�a<��a<��a<��a<Әa<}�a<�a<l�a<D�a<��a<�a<0�a<J�a<U�a<��a<Ҋa<�a<�~a<@ya<bta<�pa<�na<�ma<�na<�pa<Pta<ya<y~a<8�a<��a<�a<4�a<��a<��a<:�a<r�a<��a<@�a<n�a<��a<��a<H�a<5�a<Ϗa<�a<ɐa<�a<m�a<��a<��a<�a<ߕa<Y�a<��a<9�a<��a<�a<�}a<�wa<qa<Aka<4fa<�ba<V`a<�_a<\`a<qba<fa<qja<�oa<�ta<�ya<(~a<�a<<�a<��a<�a<D�a<̓a<Ɂa<�a<:}a<�za<Pya<xa<�wa<�wa<Ixa<vya<�za<�{a<I|a<�|a<�{a<�ya<Ewa<0sa<na<�ha<�ba<]\a<KVa<Qa<�La<�Ia<uHa<�Ha<JJa<OMa<�Qa<�Va<�\a<ba<~ga<!la<�oa<�ra</ta<�ta<[ta<^sa<�qa<-pa<ina<�la<la<�ka<la<ma<nna<Ipa<�qa<�sa<�  �  �ua<va<\ua<�sa<�pa<�la< ha<qba<�\a<�Va<�Qa<Ma<�Ia<�Ga<oGa<�Ha<�Ka<#Pa<�Ua<�[a<Oba<�ha<�na<Lta<�xa<|a<A~a<�a<�a<�a<�~a<�}a<�|a<�|a<t|a<}a<~a<�a<��a<�a<*�a<�a<Y�a<�a<g�a<�a<-�a<��a<�|a<�wa<cra<Uma<�ha<�da<}ba<caa<ba<]da<ha<ma<%sa<�ya<W�a<ǆa<�a<�a<�a<�a<��a<g�a<\�a<��a<h�a<�a< �a<e�a< �a<]�a<2�a<[�a<ՙa<��a<#�a<?�a<��a<-�a<Ŝa<,�a<h�a<đa<)�a<Z�a<W�a<�za<�ua<�qa<�na<�ma<Rna<�pa<ta<�xa<�~a<{�a<��a<x�a<Õa<��a<>�a<9�a<B�a<A�a<��a<D�a<��a<!�a<��a<�a<Øa<ݘa<��a<��a<�a<~�a<Ȟa<W�a<W�a<I�a<T�a<�a<Ӕa<��a<��a<l�a<I}a<�wa<�ra<�na<8la<_ka<Fla<�na<jra<\wa<�|a<Âa<��a<�a<Ȓa<��a<7�a<��a<+�a<��a<��a<��a<<�a<��a<]�a<a�a<	�a<(�a<Ԓa<��a<��a<�a<�a<
�a<g�a<��a<��a<��a<�a<�a<�|a<�ua<{oa<`ia<Uda<{`a<�]a<7]a<0^a<�`a<&da<�ha<�ma<osa<�xa<u}a<:�a<-�a<߅a<��a<'�a<�a<?�a<�a<�~a< }a<h{a<Pza<�ya<�ya<Cza<
{a<|a<}a<�}a<L}a<>|a<Eza<wa<�ra<�ma<�ga<Baa<�Za<�Ta<Oa<�Ja<�Ga<Fa<QFa<=Ha<sKa<�Oa<BUa<�Za<�`a<�fa<�ka<�oa<�ra<�ta<ua<gua<�ta<Lsa<�qa<%pa<oa<(na<�ma<*na<oa<8pa<�qa<sa<ua<�  �  :ya<Uya<>xa<�ua<�qa<Mla<�ea<.^a<�Ua<Na<�Fa<k@a<�;a<9a<9a<):a<;>a<�Ca<)Ka<qSa<*\a<�da<�la<2ta<�ya<�~a<R�a<܂a<A�a<��a<��a<d�a<1a<m~a<&~a<�~a<�a<�a<9�a<�a<X�a<��a<�a<R�a<��a<�a<�a<��a<Eza<*sa<wka<Gda<�]a<�Xa<�Ta<oSa< Ta<rVa<�[a<�aa<ja<�ra<�{a<U�a<=�a<�a<Z�a<m�a<��a<��a<x�a<R�a<*�a<S�a<�a<јa<s�a<��a<��a<+�a<�a<D�a<Ơa<:�a<��a<ۡa<�a<
�a<�a<��a<1�a<�a<�xa<qa<ja<�da<�`a<�_a<I`a<�ba<�ga<Mna<	va<)~a<��a<r�a<��a<R�a<ɟa<��a<�a<L�a<\�a<֡a<�a<�a<�a<@�a<�a<�a<�a<��a<Y�a<�a<t�a<_�a<0�a<̡a<��a<��a<Ԕa<��a<�a<N}a<ua<ma<nfa<Faa<^a<�]a< ^a<�aa<�fa<dma<ua<'}a<Q�a<��a<4�a<8�a<&�a<8�a<�a<��a<>�a<��a<o�a<f�a<ŕa<��a<G�a<|�a<~�a<͖a<��a<řa<�a<'�a<@�a<3�a<Q�a<)�a<��a<��a<=xa<&oa<�fa<a^a<�Wa<�Ra<�Oa<;Oa<Pa<�Sa<�Xa<�_a<�fa<tna<�ua<Z|a<�a<��a<݈a<��a<͉a<��a<e�a<A�a<w�a<$a<0}a<�{a<m{a<�{a<r|a<�}a<.a<�a<�a<��a<Sa<�|a<exa<�ra<�ka<�ca<][a<�Ra<eJa<�Ba<O=a<�8a<�7a<�7a<�9a<�>a<�Da<)La<Ta<W\a<�ca<�ja<Rpa<�ta<fwa<�xa<�xa<�wa<0va<hta<era<�pa<�oa<loa<�oa<�pa<pra<{ta<dva<xa<�  �  �xa<�xa<�wa<�ua<�qa<�la<�ea<�^a<�Va<�Na<�Ga<bAa<�<a<�9a<}9a<-;a<;?a<�Da<La<1Ta<�\a<iea<[ma<rta<za<K~a<��a<��a<ǂa<#�a<݀a<�a<[~a<�}a<T}a<�}a<a<�a<p�a<�a<��a<�a<��a<�a<.�a<��a<<�a<�a<�za<�sa<,la<ea<�^a<cYa<�Ua<Ta<�Ta<�Wa<�\a<�ba<�ja<^sa<H|a<ʄa<��a<E�a<z�a<�a<L�a<*�a<��a<��a<4�a<��a< �a<�a<��a<ӗa<Ęa<^�a<N�a<S�a<K�a<��a<:�a<��a<��a<0�a<O�a<��a<��a<��a<�ya<�qa<ka<�ea<�aa<l`a<aa<da<�ha<Boa<�va<�~a<+�a<�a<ܕa<��a<��a<a�a<ƣa<ɣa<�a<�a<-�a<<�a<��a<v�a<�a<=�a<4�a<��a<{�a<=�a<��a<ޢa<ڢa<y�a<�a<��a<!�a<!�a<a�a<�}a<�ua<na<fga<\ba<�^a<�]a<$_a<�ba<�ga<Ona<�ua<�}a<��a<
�a<u�a<c�a<�a<�a<��a<1�a<ǜa<��a<��a<��a<��a<ɓa<g�a<��a<��a<�a<��a<!�a<g�a<��a<��a<��a<i�a<]�a<�a<*�a<�xa<�oa<bga<e_a<�Xa<�Sa<�Pa<�Oa<EQa<�Ta<�Ya<Y`a<sga<oa<2va<�|a<�a<�a<��a<��a<V�a<�a<υa<K�a<��a<]~a<`|a< {a<�za<�za<�{a<�|a<>~a<�a<d�a<G�a<�~a<|a<�xa<!sa<Dla<wda< \a<dSa<IKa<�Ca<D>a<:a<*8a<u8a<";a<�?a<�Ea<�La<�Ta<�\a<Eda<ka<�pa<�ta<wa<Xxa<Bxa<Hwa<pua<�sa<�qa<�oa<�na<�na<�na<�oa<�qa<�sa<�ua<�wa<�  �  Qwa<2xa<~wa<�ua<ra<?ma<(ga<`a<�Xa<�Pa<Ja<Da<�?a<7=a<�<a<u>a<�Aa<Ga<zNa<HVa<�^a<�fa<sna<�ta<Qza<~a<��a<��a<C�a<{�a<�~a<F}a<�{a<�za<lza<�za<=|a<G~a<�a<܃a<�a<��a<Q�a<m�a<Ћa<�a<��a<�a<�{a<Uua<=na<Gga<+aa<�[a<�Xa<LWa<�Wa<�Za<(_a<�ea<ma<uua<�}a<�a<��a<��a<��a<śa<ȝa<��a<_�a<�a<��a<*�a<Y�a<#�a<��a<�a<�a<��a<�a<!�a<��a<.�a<3�a<�a<_�a<f�a<��a<�a<�a<��a<�{a<>ta<�ma<gha<6ea<�ca<Tda<ga<}ka<�qa<�xa<ڀa<��a<�a<��a<Лa<��a<��a<�a<m�a<H�a<)�a<�a<��a<јa<��a<�a<c�a<i�a<�a<4�a<B�a<^�a<u�a<�a<�a<Ϟa<��a<ƕa<O�a<ۇa<�a<�wa<�pa<ja<;ea<?ba<&aa<mba<bea<Sja<�pa<�wa<�a<$�a<#�a<�a<��a<��a<u�a<��a<��a<�a<��a<Q�a<�a<�a<��a<\�a<Ґa<��a<��a<a�a<T�a<Ϙa<r�a<Z�a<��a<��a<��a<��a<q�a<hza<�qa<�ia<ba<c[a<�Va<�Sa<Sa<vTa<iWa<}\a<�ba<�ia<�pa<�wa<�}a<{�a<?�a<5�a<�a<*�a<y�a<�a<�a<O~a<�{a<�ya<xa<�wa<�wa<�xa<�za<|a<�}a<�~a<?a<�~a<F|a<�xa<�sa<Nma<�ea<�]a<vUa<�Ma<�Fa<�@a<U=a<X;a<�;a<>a<2Ba<7Ha<Oa<�Va<P^a<~ea<�ka<�pa<�ta<�va<�wa<�va<�ua<�sa<Cqa<oa</ma<la<uka<la<.ma<oa<Vqa<�sa<�ua<�  �  Jua<�va<�va<zua<�ra<mna<�ha<�ba<�[a<~Ta<Na<wHa<$Da<�Aa<eAa<�Ba<vFa<�Ka<RRa<�Ya<�aa<ia<pa<�ua<�za<�}a<�a<�a<a<�}a<�{a<kya<�wa<mva<�ua<eva<�wa<�ya<�|a<]�a<ԃa<�a<}�a<�a<L�a<)�a<W�a<d�a<~a<�wa<vqa<�ja<Gea<�`a<?]a<�[a<�\a<,_a<�ca<�ia<�pa<�xa<��a<-�a<�a<|�a<��a<W�a<��a<6�a<�a<�a<��a<�a<�a<ϐa<%�a<r�a<��a<o�a<�a<�a<��a<�a<��a<�a<�a<��a<��a<��a<5�a<C�a<a<xa<�qa<�la<�ia<Wha<�ha<{ka<�oa<�ua<}|a<�a<+�a<��a<ݗa<h�a<��a<E�a<��a<|�a<��a<	�a<I�a<��a<��a<�a<��a<�a<�a<��a<|�a< �a<��a<m�a<��a<D�a<��a<��a<��a<�a<E�a<�a<l{a<�ta<|na<�ia<�fa<�ea<�fa<�ia<�na<�ta<U{a<��a<i�a<̏a<��a<�a<��a<|�a<�a<��a<<�a<c�a<v�a<��a<ōa<g�a<�a<k�a<��a<��a<�a<@�a<L�a<��a< �a<��a<��a<w�a<0�a<v�a<}a<%ua<'ma< fa<�_a<;[a<�Xa<�Wa<�Xa<�[a<�`a<<fa<�la<[sa<�ya</a<V�a<\�a<Ǉa<ʇa<c�a<�a<�a<�}a<?za<Pwa</ua<�sa<4sa<�sa<�ta<�va<�xa<�za<�|a<�}a<{}a<�{a<	ya<�ta<�na<ha<�`a<�Xa<kQa<�Ja<sEa<�Aa<@a<R@a<�Ba<�Fa<6La<�Ra<�Ya<�`a<Zga<ma<hqa<�ta<�ua<"va<�ta<�ra<epa<�ma<�ja<�ha<�ga<	ga<�ga<�ha<�ja<�ma<{pa<-sa<�  �  �ra<�ta<�ua<)ua<Csa<�oa<,ka<�ea<X_a<Ya<�Ra<Na<8Ja<�Ga<�Ga<Ia<vLa<1Qa<9Wa<$^a<ea<�ka<(ra<Uwa<{a<a}a<>~a<�}a<6|a<�ya<<wa<nta<+ra<�pa<�oa<Fpa<�qa<�ta<�wa<�{a<�a<��a<�a<V�a<{�a<�a<O�a<�a<��a<+{a<ua<�oa<bja<Ofa<_ca<?ba<�ba<Oea<�ia<�na<�ua<�|a<�a<Ɗa<ǐa<��a<ɘa<��a<ךa<�a<Ǘa<��a<�a<�a<��a<Ȋa<��a<>�a<��a<�a<��a<��a<ȗa<��a<]�a<��a<��a<��a<��a<��a<�a<Ɖa<a�a<�|a<Awa<�ra<�oa<�na<+oa<�qa<�ua<�za<7�a<Ňa<M�a<F�a<g�a<)�a<o�a<?�a<��a<ݝa<
�a<�a<��a<W�a<ڎa<�a<k�a<��a<Z�a<��a<��a<�a<��a<��a<��a<#�a<c�a<&�a<r�a<U�a<U�a<��a<�a<vya<
ta<�oa<ma<+la<ma<�oa<	ta<xya<�a<�a<X�a<ڑa<Y�a<m�a<�a<%�a<��a<��a<h�a<�a<x�a<`�a<�a<<�a<΅a<b�a<�a<Z�a<P�a<7�a<��a<5�a<C�a<+�a<��a<o�a<،a<�a<>�a<-ya<�qa<;ka<�ea<Zaa<�^a<�]a<�^a<�aa<�ea<ka<�pa<�va</|a<�a<f�a<j�a<�a<!�a<�a<�a<
}a<#ya<'ua<�qa<)oa<�ma<ma<�ma<Xoa<�qa<jta<wa<�ya<i{a<|a<h{a<Vya<�ua<�pa<�ja<da<5]a<PVa<0Pa<kKa<�Ga<SFa<�Fa<�Ha<ULa<4Qa<UWa<�]a<�ca<�ia<�na<*ra<Gta<�ta<4ta<Zra<toa<Fla<�ha<�ea<:ca<taa<�`a<caa<"ca<�ea<�ha<Lla<�oa<�  �  Foa<`ra<<ta<�ta<�sa<�qa<�ma<ia<�ca<H^a<�Xa<`Ta<�Pa<"Oa<�Na<APa<!Sa<�Wa<]a<"ca<Oia<Voa<�ta<�xa<�{a<�|a<�|a<<{a<�xa<�ua<ra<�na<�ka<�ia<�ha<Zia<�ja<�ma<�qa<Ava<${a<�a<�a<k�a<c�a<�a<L�a<�a<��a<a<za<.ua<�pa<�la<[ja<]ia<�ia<Zla<pa<&ua<6{a<��a<�a<�a<˒a<��a<טa<��a<�a<�a<�a<q�a<��a<��a<	�a<�a<�a<l�a<�a<��a<�a<1�a<}�a<Q�a<��a<�a<a<J�a<B�a<՗a<U�a<�a<@�a<��a<�}a<�ya<�va<�ua<Rva<ixa<|a<؀a<y�a<5�a<��a<�a<�a<�a<"�a<��a<{�a<��a<	�a<��a<؎a<�a<*�a<6�a<r�a<�a<��a<g�a<�a<�a<�a<h�a<9�a<ȝa<��a<ʜa<
�a<��a<�a<�a<8�a<sa<gza<�va</ta<Vsa<>ta<�va<`za<Pa<Ƅa<Q�a<��a<@�a<��a<ՙa<\�a<��a<g�a<�a<3�a<܋a<��a<�a<�a<la<�~a<�a<v�a<>�a<ća<��a<�a<*�a<V�a<�a<s�a<j�a<��a<��a<"�a<�}a<rwa<^qa<3la<Wha<�ea<ea<fa<Qha<�ka<�pa<�ua<�za<Ma<�a<|�a<y�a<�a<O�a<"�a<}a<�xa<�sa<oa<Hka<Oha<�fa</fa<�fa<�ha<�ka<oa<�ra<�ua<�xa<iza<�za<�ya<wa<sa<na<4ha<ba<\a<|Va<Ra<Oa<wMa<�Ma<oOa<�Ra<>Wa<�\a<ba<�ga<rla<Mpa<�ra<�sa<�sa<ra<!oa<tka<[ga<1ca<x_a<�\a<�Za<�Ya<�Za<o\a<[_a<	ca<Cga<�ka<�  �  �ka<�oa<�ra<Zta<�ta<#sa<�pa<�la<}ha<�ca<?_a<Y[a<TXa<�Va<dVa<�Wa<aZa<_^a< ca<fha<�ma<�ra<wa<za<�{a<|a<�za<oxa<�ta<�pa<\la<Zha<�da<oba<aaa<�aa<�ca<�fa</ka<Qpa<�ua<�{a<΀a<.�a<8�a<�a<3�a<�a<��a<�a<&a<�za<wa<�sa<�qa<�pa<�qa<�sa<7wa<�{a<��a<��a<�a<�a<�a<��a<�a<��a<�a<ӓa<�a<b�a<��a<��a<�~a<�|a<c{a<�{a<�}a<��a<ʄa<y�a<��a<z�a<��a<�a<��a<��a<��a<J�a<��a<Y�a<y�a<��a<]�a<��a<|~a<[}a<�}a<�a<�a<>�a<�a<�a<ʕa<�a<�a<��a<ܞa<��a<��a<)�a<��a<��a<Ɉa<u�a<�a<�~a<�}a<n~a<U�a<��a<ɇa<i�a<_�a<ѕa<��a<4�a<��a<d�a<��a<��a<��a<ۏa<��a<��a<c�a<�}a<�{a<�za<�{a<�}a<;�a<c�a<�a<��a<3�a<іa<�a<8�a<��a<ӗa<��a<W�a<~�a<7�a<e�a<!}a<�ya<�wa<)wa<+xa<Oza<�}a<Ӂa<d�a<�a<�a<�a<�a<l�a<R�a<ѐa<��a<.�a<Ԃa< }a<�wa<Rsa<�oa<�ma<�la<ma<yoa<�ra<qva<�za<�~a<o�a<!�a<��a<��a<�a<-�a<~a<�xa<xsa<�ma<�ha<1da<�`a<�^a<�^a<�_a<�aa<_ea<cia<�ma<ra<�ua<zxa<�ya<�ya<Yxa<�ua<{qa<�la<Jga<ba<H]a<?Ya<�Va<Ua<MUa<�Va<�Ya<�]a<ba<�fa<gka<Hoa<ra<�sa<�sa<;ra<�oa<�ka<ga<�aa<$]a<�Xa<IUa<1Sa<@Ra<Sa<!Ua<�Xa<�\a<�aa<�fa<�  �  	ha<ma<qa<�sa<�ta<�ta<4sa<tpa<ma<3ia<^ea<#ba<�_a<E^a<^a<A_a<�aa<�da<%ia<�ma<1ra<>va<�ya<{{a<|a<[{a<ya<�ua<qa<�ka<�fa<�aa<�]a<[a<�Ya<Za<\a<�_a<jda<ija<�pa<Fwa<�}a<Ȃa< �a<ȉa<
�a<�a<��a<�a<
�a<��a<d}a<�za<ya<�xa<Qya<&{a<E~a<2�a<҆a<��a<�a<�a<�a<��a<ɘa<z�a<��a<��a<��a<<�a<�a<�{a<�wa<ua<�sa<(ta<!va<�ya<A~a<׃a<��a<|�a<Ôa<�a<$�a<��a<̝a<��a<�a<��a<��a<��a<�a<�a<��a<�a<��a<#�a<�a<i�a<��a<Õa<}�a<��a<��a<,�a<k�a<�a<d�a<��a<	�a<O�a<��a<�}a<�ya<)wa<!va<�va<ya<�|a<��a<�a<��a<)�a<�a<��a<�a<֝a<L�a<^�a<:�a<m�a<%�a<ߋa<.�a<6�a<U�a<��a<B�a<�a<؇a<j�a<`�a<8�a<��a<=�a<��a<m�a<��a<��a<��a<t�a<��a<��a<�za<va<_ra<3pa<�oa<�pa<sa<�va<�{a<2�a<��a<��a<��a<��a<1�a<(�a<Βa<��a<�a<��a<�a<=~a<Lza<wa</ua<lta<�ta<�va<ya<G|a<�a<܂a<��a<8�a<z�a<l�a<�a<�a<�za<�ta<Sna<�ga<�aa<]a<}Ya<NWa<�Va<#Xa<�Za<�^a<�ca<�ha< na<�ra<xva<ya<�ya<�ya<�wa<�ta<�pa<�la<�ga<�ca<m`a<�]a<�\a<�\a<%^a<�`a<�ca<�ga<�ka<oa<ra<�sa<.ta<Dsa<�pa<�la<ha<wba<�\a<Wa<�Qa<Na<�Ka<�Ja<}Ka<�Ma<�Qa<�Va<o\a<Eba<�  �  �da<�ja<�oa<8sa<nua<+va<�ua<�sa<&qa<Gna<&ka<mha<[fa<ea<ea<fa<Iha<-ka<�na<�ra<)va<hya<�{a<�|a<S|a<�za<Iwa<�ra<Qma<nga<�aa<�[a<pWa<,Ta<�Ra<�Ra<�Ta<�Xa<#^a<�da<�ka<.sa<Bza<��a<ƅa<��a<ۋa<��a<L�a<��a<b�a<��a<]�a<_�a<�a<xa<,�a<�a<ӄa<4�a<;�a<�a<�a<��a<ۘa<��a<��a<V�a<��a<x�a<��a<��a<C{a<�ua<:qa<na<�la<	ma</oa<sa<%xa<r~a<�a<��a<ϑa<*�a<7�a<ǝa<�a<��a<�a<�a<n�a<9�a<	�a<��a<��a<�a<W�a<�a<D�a<B�a<��a<�a<��a<!�a< �a<ğa<��a<��a<�a<6�a<ȉa<A�a<�|a<9wa<�ra<�oa<�na<�oa<Bra<Xva<�{a<�a<P�a<��a<W�a<�a<q�a<Q�a<��a<��a<��a<��a<:�a<��a<y�a<�a<$�a<��a<�a<��a<�a<�a<=�a<2�a<˙a<S�a<��a<��a<.�a<4�a<�a<��a<�a<b{a<�ta<�oa<�ka<ia<gha<�ia<�la<�pa<3va<a|a<u�a<_�a<z�a<s�a<��a<��a<t�a<��a<ɏa<�a<:�a<5�a<ɀa<�}a<|a<H{a<�{a<}a<a<��a<5�a<��a<g�a<��a<k�a<P�a<ʂa<�}a<�wa<�pa<�ia<^ba<�[a<|Va<kRa<1Pa<�Oa<1Qa<cTa<�Xa<\^a<\da<Kja<�oa<�ta<xa<za<�za<�ya<�wa<�ta<<qa<�ma<�ia<ga<�da<�ca<�ca<�da<�fa<�ia<�la<�oa<�ra<�ta<Qua<�ta<�ra<_oa<�ja<�da<8^a<�Wa<$Qa<�Ka<QGa<uDa<�Ca<VDa<Ga<RKa<�Pa<OWa<�]a<�  �  �aa<Lha<na<�ra<�ua<Xwa<�wa<�va<�ta<}ra<pa<�ma< la<9ka<-ka<!la<�ma<jpa<�sa<�va<�ya<�{a<}}a<�}a<�|a<�ya<�ua<[pa<)ja<�ca<�\a<�Va<�Qa<Na<`La<�La<�Na<�Ra<�Xa<�_a<�ga<�oa<|wa<�~a<��a<M�a<w�a<1�a<|�a<��a<L�a<`�a<i�a<a<��a<��a<]�a<�a<@�a<H�a<��a<�a<�a<>�a<y�a<;�a<��a<;�a<��a<ϊa<9�a<T}a<cva<ppa<Uka<�ga<^fa<�fa<ia<Xma<sa<�ya<�a<q�a<`�a<��a<M�a<�a<͟a<[�a<��a<ݝa<~�a<טa<;�a<�a<Òa<%�a<��a<��a<��a<9�a<�a<��a<ӟa<9�a<h�a<8�a<�a<C�a<ғa<>�a<%�a<�~a<�wa<�qa<�la<�ia<�ha<~ia<1la<�pa<�va<Y}a<��a<��a<#�a<��a<ݛa<��a<�a<Ɵa<Y�a<1�a<q�a<��a<Ɠa<��a<L�a<��a<&�a<]�a<L�a<ɕa<Y�a<��a<`�a<7�a<��a<�a<a�a<��a<��a<��a<*~a<�va<�oa<�ia<hea<�ba<'ba<`ca<�fa<xka<Nqa<xa<�~a<��a<��a<>�a<��a<��a<��a<�a<ƒa<��a<��a<A�a<,�a<�a<7�a<x�a<��a<��a<"�a<)�a<-�a<��a<��a<��a<�a<1�a<��a<|a< ua<Xma<lea<]a<�Va<�Pa<DLa<�Ia<�Ia<Ka<�Na<�Sa<�Ya<]`a<ga<ima<�ra<.wa<<za<�{a<�{a<Rza<#xa<Jua</ra<"oa<�la<�ja<�ia<�ia<�ja<Mla<�na< qa<�sa<oua<�va<�va<<ua<Zra<�ma<lha<�aa<�Za<*Sa<;La<1Fa<MAa<M>a<>=a<+>a<Aa<�Ea<�Ka<�Ra<3Za<�  �  !_a<�fa<�la<)ra<�ua<+xa<+ya<�xa<�wa<�ua<�sa<�qa<qpa<�oa<�oa<�pa<2ra<�ta<wa<�ya<J|a<�}a<�~a<M~a<�|a<ya<eta<sna<�ga<n`a<6Ya<�Ra<>Ma<�Ia<�Ga<�Ga<eJa<tNa<�Ta<\a<Nda<�la<Tua<}a<��a<�a<ˌa<T�a</�a<�a<H�a<��a<^�a<��a<3�a<�a<Ȋa<P�a<��a<P�a<�a<�a<e�a< �a<��a<��a<e�a<X�a<.�a<��a<��a<za<�ra<<la<�fa<{ca<�aa<ba<�da<�ha<�na<
va<�}a<ޅa<c�a<�a<��a<�a<]�a<��a<l�a<l�a<��a<`�a<R�a<h�a<1�a<��a<��a<�a<əa<�a<1�a<��a<��a<آa<S�a<h�a<�a</�a<!�a<�a<E�a<T{a<�sa<qma<gha<Nea<�ca<�da<�ga<gla<�ra<�ya<��a<?�a<d�a<��a<b�a<͞a<��a<V�a<j�a<�a<��a<L�a<�a<�a<ʔa<'�a<��a<��a<h�a<d�a<u�a<U�a<G�a<��a<Z�a<�a<��a<R�a<��a<�a<{a<sa<�ka<rea<�`a<0^a<n]a<�^a<ba<3ga<�ma<�ta<E|a<o�a<�a<K�a<x�a<�a<�a<��a<�a<��a<�a<6�a<e�a<.�a<��a<�a<��a<Æa<*�a<��a<5�a<#�a<l�a<֋a<~�a<
�a<̀a<|za<�ra<�ja<ba<�Ya<fRa<La<�Ga<8Ea<�Da<�Fa<Ja<�Oa<�Ua</]a<�da<lka<�qa<rva<7za<&|a<}a<-|a<�za<`xa<�ua<8sa<�pa<Eoa<Cna<Rna<
oa<wpa<nra<Kta<mva<�wa<<xa<�wa<lua<�qa<�la<�fa<q_a<�Wa<�Oa<\Ha<�Aa<�<a<�9a<}8a<�9a<�<a<cAa<�Ga<COa<FWa<�  �  �]a<fea<]la<�qa<va<�xa<za<za<Bya<�wa<va<vta<;sa<�ra<�ra<xsa<ua<�va<Vya<�{a<�}a<6a<�a<�~a<�|a<�xa<�sa<6ma<fa<j^a<Wa<:Pa<�Ja<�Fa<�Da<�Da<'Ga<�Ka<�Qa<�Ya<<ba<7ka<�sa<|a<6�a<߈a<�a<ŏa<A�a<��a<��a<�a<��a<��a<�a<�a<ƍa<-�a<F�a<��a<O�a<Ҙa<��a<$�a</�a<�a<;�a<��a<=�a<_�a<�a<�wa<rpa<�ia<7da<F`a<s^a<�^a<�aa<9fa<_la<�sa<�{a<>�a< �a<Q�a<@�a<ȝa<��a<d�a<��a<�a<i�a<��a<a<9�a<�a<��a<��a<ښa<j�a<\�a<M�a<;�a<q�a<��a<Ģa<��a<ќa<��a<�a<��a<^�a<9ya<�qa<�ja<�ea<ba<�`a<�aa<�da<�ia<>pa<�wa<�a<ɇa<<�a<�a<�a<�a<%�a<,�a<١a<��a<��a<��a<��a<Иa<��a<8�a<�a<z�a<�a<��a<Y�a<�a<��a<^�a<ĝa<�a<n�a<��a<f�a<��a<ya<�pa<Eia<�ba<�]a<�Za<<Za<�[a<f_a<�da<=ka<�ra<|za<�a<��a<�a<G�a<&�a<��a<��a<��a<��a<%�a<��a<$�a<�a<��a<�a<ڈa<��a<��a<ŋa<�a<��a<��a<Q�a<͉a<�a<m�a<�ya<�qa<�ha<`a<�Wa<�Oa<yIa<�Da<Ba<�Aa<�Ca<�Ga<�La<�Sa<![a<�ba<(ja<�pa< va<za<�|a<�}a<q}a<H|a<3za<�wa<�ua<�sa<)ra<Qqa<5qa<�qa<sa<�ta<gva<xa<ya<%ya<�wa<�ua<�qa<cla<�ea<
^a<�Ua<�Ma<�Ea</?a<:a<�6a<X5a<S6a<�9a<�>a<lEa<#Ma<VUa<�  �  =]a<�da<la<�qa<+va<�xa<Xza<�za<�ya<yxa<�va<Kua<ta<[sa<�sa<?ta<�ua<�wa<@za<d|a<]~a<�a<�a<a<�|a<�xa<Lsa<�la<�ea<�]a<GVa<EOa<�Ia<�Ea<�Ca<+Da<Fa<�Ja<�Pa<�Xa<aa<�ja<�sa<�{a<��a<��a<Z�a<�a<��a<�a<w�a<אa<}�a<��a<�a<�a<��a<�a<�a<t�a<H�a<a�a<~�a<��a<~�a<C�a<�a<��a<Սa<�a<?a<0wa<�oa<�ha<Mca< _a<�]a<1^a<m`a<Tea<aka<sa<'{a<Ãa<��a<��a<�a<��a<�a<��a<)�a<�a<�a<��a<��a<�a<ۚa<��a<��a<��a<A�a<-�a<(�a<��a<�a<�a<�a<Ƞa<��a<i�a<��a<�a<��a<wxa<�pa<�ia<�da<aa<O`a<�`a<�ca<�ha<Poa<�va<a<Z�a<ˎa<��a<�a<�a<x�a<��a<Z�a<�a<n�a<o�a<[�a<��a<q�a< �a<G�a<W�a<��a<��a<�a<i�a<�a<��a<�a<�a<=�a<9�a<��a<�a<\xa<#pa<Pha<�aa<�\a<0Za<�Ya<�Za<v^a<�ca<Zja<�qa<�ya<��a<��a<��a<�a<v�a<��a< �a<%�a<"�a<�a<U�a<�a<�a<u�a<��a<��a<O�a<N�a<��a<x�a<<�a<�a<��a<"�a<��a</�a<$ya<qa<_ha<I_a<�Va<�Na<�Ha<�Ca<sAa<�@a<pBa<�Fa<�Ka<�Ra<kZa<gba<�ia<jpa<�ua<
za<�|a<�}a<�}a<�|a<�za<�xa<wva<�ta<�ra<5ra<ra<�ra<�sa<�ua<Bwa<�xa<�ya<|ya<Hxa<�ua<�qa<"la<,ea<�]a<'Ua<�La<Ea<2>a<9a<�5a<�4a<o5a<�8a<�=a<~Da<\La<�Ta<�  �  �]a<fea<]la<�qa<va<�xa<za<za<Bya<�wa<va<vta<;sa<�ra<�ra<xsa<ua<�va<Vya<�{a<�}a<6a<�a<�~a<�|a<�xa<�sa<6ma<fa<j^a<Wa<:Pa<�Ja<�Fa<�Da<�Da<'Ga<�Ka<�Qa<�Ya<<ba<7ka<�sa<|a<6�a<߈a<�a<ŏa<A�a<��a<��a<�a<��a<��a<�a<�a<ƍa<-�a<F�a<��a<O�a<Ҙa<��a<$�a</�a<�a<;�a<��a<=�a<_�a<�a<�wa<rpa<�ia<7da<F`a<s^a<�^a<�aa<9fa<_la<�sa<�{a<>�a< �a<Q�a<@�a<ȝa<��a<d�a<��a<�a<i�a<��a<a<9�a<�a<��a<��a<ښa<j�a<\�a<M�a<;�a<q�a<��a<Ģa<��a<ќa<��a<�a<��a<^�a<9ya<�qa<�ja<�ea<ba<�`a<�aa<�da<�ia<>pa<�wa<�a<ɇa<<�a<�a<�a<�a<%�a<,�a<١a<��a<��a<��a<��a<Иa<��a<8�a<�a<z�a<�a<��a<Y�a<�a<��a<^�a<ĝa<�a<n�a<��a<f�a<��a<ya<�pa<Eia<�ba<�]a<�Za<<Za<�[a<f_a<�da<=ka<�ra<|za<�a<��a<�a<G�a<&�a<��a<��a<��a<��a<%�a<��a<$�a<�a<��a<�a<ڈa<��a<��a<ŋa<�a<��a<��a<Q�a<͉a<�a<m�a<�ya<�qa<�ha<`a<�Wa<�Oa<yIa<�Da<Ba<�Aa<�Ca<�Ga<�La<�Sa<![a<�ba<(ja<�pa< va<za<�|a<�}a<q}a<H|a<3za<�wa<�ua<�sa<)ra<Qqa<5qa<�qa<sa<�ta<gva<xa<ya<%ya<�wa<�ua<�qa<cla<�ea<
^a<�Ua<�Ma<�Ea</?a<:a<�6a<X5a<S6a<�9a<�>a<lEa<#Ma<VUa<�  �  !_a<�fa<�la<)ra<�ua<+xa<+ya<�xa<�wa<�ua<�sa<�qa<qpa<�oa<�oa<�pa<2ra<�ta<wa<�ya<J|a<�}a<�~a<M~a<�|a<ya<eta<sna<�ga<n`a<6Ya<�Ra<>Ma<�Ia<�Ga<�Ga<eJa<tNa<�Ta<\a<Nda<�la<Tua<}a<��a<�a<ˌa<T�a</�a<�a<H�a<��a<^�a<��a<3�a<�a<Ȋa<P�a<��a<P�a<�a<�a<e�a< �a<��a<��a<e�a<X�a<.�a<��a<��a<za<�ra<<la<�fa<{ca<�aa<ba<�da<�ha<�na<
va<�}a<ޅa<c�a<�a<��a<�a<]�a<��a<l�a<l�a<��a<`�a<R�a<h�a<1�a<��a<��a<�a<əa<�a<1�a<��a<��a<آa<S�a<h�a<�a</�a<!�a<�a<E�a<T{a<�sa<qma<gha<Nea<�ca<�da<�ga<gla<�ra<�ya<��a<?�a<d�a<��a<b�a<͞a<��a<V�a<j�a<�a<��a<L�a<�a<�a<ʔa<'�a<��a<��a<h�a<d�a<u�a<U�a<G�a<��a<Z�a<�a<��a<R�a<��a<�a<{a<sa<�ka<rea<�`a<0^a<n]a<�^a<ba<3ga<�ma<�ta<E|a<o�a<�a<K�a<x�a<�a<�a<��a<�a<��a<�a<6�a<e�a<.�a<��a<�a<��a<Æa<*�a<��a<5�a<#�a<l�a<֋a<~�a<
�a<̀a<|za<�ra<�ja<ba<�Ya<fRa<La<�Ga<8Ea<�Da<�Fa<Ja<�Oa<�Ua</]a<�da<lka<�qa<rva<7za<&|a<}a<-|a<�za<`xa<�ua<8sa<�pa<Eoa<Cna<Rna<
oa<wpa<nra<Kta<mva<�wa<<xa<�wa<lua<�qa<�la<�fa<q_a<�Wa<�Oa<\Ha<�Aa<�<a<�9a<}8a<�9a<�<a<cAa<�Ga<COa<FWa<�  �  �aa<Lha<na<�ra<�ua<Xwa<�wa<�va<�ta<}ra<pa<�ma< la<9ka<-ka<!la<�ma<jpa<�sa<�va<�ya<�{a<}}a<�}a<�|a<�ya<�ua<[pa<)ja<�ca<�\a<�Va<�Qa<Na<`La<�La<�Na<�Ra<�Xa<�_a<�ga<�oa<|wa<�~a<��a<M�a<w�a<1�a<|�a<��a<L�a<`�a<i�a<a<��a<��a<]�a<�a<@�a<H�a<��a<�a<�a<>�a<y�a<;�a<��a<;�a<��a<ϊa<9�a<T}a<cva<ppa<Uka<�ga<^fa<�fa<ia<Xma<sa<�ya<�a<q�a<`�a<��a<M�a<�a<͟a<[�a<��a<ݝa<~�a<טa<;�a<�a<Òa<%�a<��a<��a<��a<9�a<�a<��a<ӟa<9�a<h�a<8�a<�a<C�a<ғa<>�a<%�a<�~a<�wa<�qa<�la<�ia<�ha<~ia<1la<�pa<�va<Y}a<��a<��a<#�a<��a<ݛa<��a<�a<Ɵa<Y�a<1�a<q�a<��a<Ɠa<��a<L�a<��a<&�a<]�a<L�a<ɕa<Y�a<��a<`�a<7�a<��a<�a<a�a<��a<��a<��a<*~a<�va<�oa<�ia<hea<�ba<'ba<`ca<�fa<xka<Nqa<xa<�~a<��a<��a<>�a<��a<��a<��a<�a<ƒa<��a<��a<A�a<,�a<�a<7�a<x�a<��a<��a<"�a<)�a<-�a<��a<��a<��a<�a<1�a<��a<|a< ua<Xma<lea<]a<�Va<�Pa<DLa<�Ia<�Ia<Ka<�Na<�Sa<�Ya<]`a<ga<ima<�ra<.wa<<za<�{a<�{a<Rza<#xa<Jua</ra<"oa<�la<�ja<�ia<�ia<�ja<Mla<�na< qa<�sa<oua<�va<�va<<ua<Zra<�ma<lha<�aa<�Za<*Sa<;La<1Fa<MAa<M>a<>=a<+>a<Aa<�Ea<�Ka<�Ra<3Za<�  �  �da<�ja<�oa<8sa<nua<+va<�ua<�sa<&qa<Gna<&ka<mha<[fa<ea<ea<fa<Iha<-ka<�na<�ra<)va<hya<�{a<�|a<S|a<�za<Iwa<�ra<Qma<nga<�aa<�[a<pWa<,Ta<�Ra<�Ra<�Ta<�Xa<#^a<�da<�ka<.sa<Bza<��a<ƅa<��a<ۋa<��a<L�a<��a<b�a<��a<]�a<_�a<�a<xa<,�a<�a<ӄa<4�a<;�a<�a<�a<��a<ۘa<��a<��a<V�a<��a<x�a<��a<��a<C{a<�ua<:qa<na<�la<	ma</oa<sa<%xa<r~a<�a<��a<ϑa<*�a<7�a<ǝa<�a<��a<�a<�a<n�a<9�a<	�a<��a<��a<�a<W�a<�a<D�a<B�a<��a<�a<��a<!�a< �a<ğa<��a<��a<�a<6�a<ȉa<A�a<�|a<9wa<�ra<�oa<�na<�oa<Bra<Xva<�{a<�a<P�a<��a<W�a<�a<q�a<Q�a<��a<��a<��a<��a<:�a<��a<y�a<�a<$�a<��a<�a<��a<�a<�a<=�a<2�a<˙a<S�a<��a<��a<.�a<4�a<�a<��a<�a<b{a<�ta<�oa<�ka<ia<gha<�ia<�la<�pa<3va<a|a<u�a<_�a<z�a<s�a<��a<��a<t�a<��a<ɏa<�a<:�a<5�a<ɀa<�}a<|a<H{a<�{a<}a<a<��a<5�a<��a<g�a<��a<k�a<P�a<ʂa<�}a<�wa<�pa<�ia<^ba<�[a<|Va<kRa<1Pa<�Oa<1Qa<cTa<�Xa<\^a<\da<Kja<�oa<�ta<xa<za<�za<�ya<�wa<�ta<<qa<�ma<�ia<ga<�da<�ca<�ca<�da<�fa<�ia<�la<�oa<�ra<�ta<Qua<�ta<�ra<_oa<�ja<�da<8^a<�Wa<$Qa<�Ka<QGa<uDa<�Ca<VDa<Ga<RKa<�Pa<OWa<�]a<�  �  	ha<ma<qa<�sa<�ta<�ta<4sa<tpa<ma<3ia<^ea<#ba<�_a<E^a<^a<A_a<�aa<�da<%ia<�ma<1ra<>va<�ya<{{a<|a<[{a<ya<�ua<qa<�ka<�fa<�aa<�]a<[a<�Ya<Za<\a<�_a<jda<ija<�pa<Fwa<�}a<Ȃa< �a<ȉa<
�a<�a<��a<�a<
�a<��a<d}a<�za<ya<�xa<Qya<&{a<E~a<2�a<҆a<��a<�a<�a<�a<��a<ɘa<z�a<��a<��a<��a<<�a<�a<�{a<�wa<ua<�sa<(ta<!va<�ya<A~a<׃a<��a<|�a<Ôa<�a<$�a<��a<̝a<��a<�a<��a<��a<��a<�a<�a<��a<�a<��a<#�a<�a<i�a<��a<Õa<}�a<��a<��a<,�a<k�a<�a<d�a<��a<	�a<O�a<��a<�}a<�ya<)wa<!va<�va<ya<�|a<��a<�a<��a<)�a<�a<��a<�a<֝a<L�a<^�a<:�a<m�a<%�a<ߋa<.�a<6�a<U�a<��a<B�a<�a<؇a<j�a<`�a<8�a<��a<=�a<��a<m�a<��a<��a<��a<t�a<��a<��a<�za<va<_ra<3pa<�oa<�pa<sa<�va<�{a<2�a<��a<��a<��a<��a<1�a<(�a<Βa<��a<�a<��a<�a<=~a<Lza<wa</ua<lta<�ta<�va<ya<G|a<�a<܂a<��a<8�a<z�a<l�a<�a<�a<�za<�ta<Sna<�ga<�aa<]a<}Ya<NWa<�Va<#Xa<�Za<�^a<�ca<�ha< na<�ra<xva<ya<�ya<�ya<�wa<�ta<�pa<�la<�ga<�ca<m`a<�]a<�\a<�\a<%^a<�`a<�ca<�ga<�ka<oa<ra<�sa<.ta<Dsa<�pa<�la<ha<wba<�\a<Wa<�Qa<Na<�Ka<�Ja<}Ka<�Ma<�Qa<�Va<o\a<Eba<�  �  �ka<�oa<�ra<Zta<�ta<#sa<�pa<�la<}ha<�ca<?_a<Y[a<TXa<�Va<dVa<�Wa<aZa<_^a< ca<fha<�ma<�ra<wa<za<�{a<|a<�za<oxa<�ta<�pa<\la<Zha<�da<oba<aaa<�aa<�ca<�fa</ka<Qpa<�ua<�{a<΀a<.�a<8�a<�a<3�a<�a<��a<�a<&a<�za<wa<�sa<�qa<�pa<�qa<�sa<7wa<�{a<��a<��a<�a<�a<�a<��a<�a<��a<�a<ӓa<�a<b�a<��a<��a<�~a<�|a<c{a<�{a<�}a<��a<ʄa<y�a<��a<z�a<��a<�a<��a<��a<��a<J�a<��a<Y�a<y�a<��a<]�a<��a<|~a<[}a<�}a<�a<�a<>�a<�a<�a<ʕa<�a<�a<��a<ܞa<��a<��a<)�a<��a<��a<Ɉa<u�a<�a<�~a<�}a<n~a<U�a<��a<ɇa<i�a<_�a<ѕa<��a<4�a<��a<d�a<��a<��a<��a<ۏa<��a<��a<c�a<�}a<�{a<�za<�{a<�}a<;�a<c�a<�a<��a<3�a<іa<�a<8�a<��a<ӗa<��a<W�a<~�a<7�a<e�a<!}a<�ya<�wa<)wa<+xa<Oza<�}a<Ӂa<d�a<�a<�a<�a<�a<l�a<R�a<ѐa<��a<.�a<Ԃa< }a<�wa<Rsa<�oa<�ma<�la<ma<yoa<�ra<qva<�za<�~a<o�a<!�a<��a<��a<�a<-�a<~a<�xa<xsa<�ma<�ha<1da<�`a<�^a<�^a<�_a<�aa<_ea<cia<�ma<ra<�ua<zxa<�ya<�ya<Yxa<�ua<{qa<�la<Jga<ba<H]a<?Ya<�Va<Ua<MUa<�Va<�Ya<�]a<ba<�fa<gka<Hoa<ra<�sa<�sa<;ra<�oa<�ka<ga<�aa<$]a<�Xa<IUa<1Sa<@Ra<Sa<!Ua<�Xa<�\a<�aa<�fa<�  �  Foa<`ra<<ta<�ta<�sa<�qa<�ma<ia<�ca<H^a<�Xa<`Ta<�Pa<"Oa<�Na<APa<!Sa<�Wa<]a<"ca<Oia<Voa<�ta<�xa<�{a<�|a<�|a<<{a<�xa<�ua<ra<�na<�ka<�ia<�ha<Zia<�ja<�ma<�qa<Ava<${a<�a<�a<k�a<c�a<�a<L�a<�a<��a<a<za<.ua<�pa<�la<[ja<]ia<�ia<Zla<pa<&ua<6{a<��a<�a<�a<˒a<��a<טa<��a<�a<�a<�a<q�a<��a<��a<	�a<�a<�a<l�a<�a<��a<�a<1�a<}�a<Q�a<��a<�a<a<J�a<B�a<՗a<U�a<�a<@�a<��a<�}a<�ya<�va<�ua<Rva<ixa<|a<؀a<y�a<5�a<��a<�a<�a<�a<"�a<��a<{�a<��a<	�a<��a<؎a<�a<*�a<6�a<r�a<�a<��a<g�a<�a<�a<�a<h�a<9�a<ȝa<��a<ʜa<
�a<��a<�a<�a<8�a<sa<gza<�va</ta<Vsa<>ta<�va<`za<Pa<Ƅa<Q�a<��a<@�a<��a<ՙa<\�a<��a<g�a<�a<3�a<܋a<��a<�a<�a<la<�~a<�a<v�a<>�a<ća<��a<�a<*�a<V�a<�a<s�a<j�a<��a<��a<"�a<�}a<rwa<^qa<3la<Wha<�ea<ea<fa<Qha<�ka<�pa<�ua<�za<Ma<�a<|�a<y�a<�a<O�a<"�a<}a<�xa<�sa<oa<Hka<Oha<�fa</fa<�fa<�ha<�ka<oa<�ra<�ua<�xa<iza<�za<�ya<wa<sa<na<4ha<ba<\a<|Va<Ra<Oa<wMa<�Ma<oOa<�Ra<>Wa<�\a<ba<�ga<rla<Mpa<�ra<�sa<�sa<ra<!oa<tka<[ga<1ca<x_a<�\a<�Za<�Ya<�Za<o\a<[_a<	ca<Cga<�ka<�  �  �ra<�ta<�ua<)ua<Csa<�oa<,ka<�ea<X_a<Ya<�Ra<Na<8Ja<�Ga<�Ga<Ia<vLa<1Qa<9Wa<$^a<ea<�ka<(ra<Uwa<{a<a}a<>~a<�}a<6|a<�ya<<wa<nta<+ra<�pa<�oa<Fpa<�qa<�ta<�wa<�{a<�a<��a<�a<V�a<{�a<�a<O�a<�a<��a<+{a<ua<�oa<bja<Ofa<_ca<?ba<�ba<Oea<�ia<�na<�ua<�|a<�a<Ɗa<ǐa<��a<ɘa<��a<ךa<�a<Ǘa<��a<�a<�a<��a<Ȋa<��a<>�a<��a<�a<��a<��a<ȗa<��a<]�a<��a<��a<��a<��a<��a<�a<Ɖa<a�a<�|a<Awa<�ra<�oa<�na<+oa<�qa<�ua<�za<7�a<Ňa<M�a<F�a<g�a<)�a<o�a<?�a<��a<ݝa<
�a<�a<��a<W�a<ڎa<�a<k�a<��a<Z�a<��a<��a<�a<��a<��a<��a<#�a<c�a<&�a<r�a<U�a<U�a<��a<�a<vya<
ta<�oa<ma<+la<ma<�oa<	ta<xya<�a<�a<X�a<ڑa<Y�a<m�a<�a<%�a<��a<��a<h�a<�a<x�a<`�a<�a<<�a<΅a<b�a<�a<Z�a<P�a<7�a<��a<5�a<C�a<+�a<��a<o�a<،a<�a<>�a<-ya<�qa<;ka<�ea<Zaa<�^a<�]a<�^a<�aa<�ea<ka<�pa<�va</|a<�a<f�a<j�a<�a<!�a<�a<�a<
}a<#ya<'ua<�qa<)oa<�ma<ma<�ma<Xoa<�qa<jta<wa<�ya<i{a<|a<h{a<Vya<�ua<�pa<�ja<da<5]a<PVa<0Pa<kKa<�Ga<SFa<�Fa<�Ha<ULa<4Qa<UWa<�]a<�ca<�ia<�na<*ra<Gta<�ta<4ta<Zra<toa<Fla<�ha<�ea<:ca<taa<�`a<caa<"ca<�ea<�ha<Lla<�oa<�  �  Jua<�va<�va<zua<�ra<mna<�ha<�ba<�[a<~Ta<Na<wHa<$Da<�Aa<eAa<�Ba<vFa<�Ka<RRa<�Ya<�aa<ia<pa<�ua<�za<�}a<�a<�a<a<�}a<�{a<kya<�wa<mva<�ua<eva<�wa<�ya<�|a<]�a<ԃa<�a<}�a<�a<L�a<)�a<W�a<d�a<~a<�wa<vqa<�ja<Gea<�`a<?]a<�[a<�\a<,_a<�ca<�ia<�pa<�xa<��a<-�a<�a<|�a<��a<W�a<��a<6�a<�a<�a<��a<�a<�a<ϐa<%�a<r�a<��a<o�a<�a<�a<��a<�a<��a<�a<�a<��a<��a<��a<5�a<C�a<a<xa<�qa<�la<�ia<Wha<�ha<{ka<�oa<�ua<}|a<�a<+�a<��a<ݗa<h�a<��a<E�a<��a<|�a<��a<	�a<I�a<��a<��a<�a<��a<�a<�a<��a<|�a< �a<��a<m�a<��a<D�a<��a<��a<��a<�a<E�a<�a<l{a<�ta<|na<�ia<�fa<�ea<�fa<�ia<�na<�ta<U{a<��a<i�a<̏a<��a<�a<��a<|�a<�a<��a<<�a<c�a<v�a<��a<ōa<g�a<�a<k�a<��a<��a<�a<@�a<L�a<��a< �a<��a<��a<w�a<0�a<v�a<}a<%ua<'ma< fa<�_a<;[a<�Xa<�Wa<�Xa<�[a<�`a<<fa<�la<[sa<�ya</a<V�a<\�a<Ǉa<ʇa<c�a<�a<�a<�}a<?za<Pwa</ua<�sa<4sa<�sa<�ta<�va<�xa<�za<�|a<�}a<{}a<�{a<	ya<�ta<�na<ha<�`a<�Xa<kQa<�Ja<sEa<�Aa<@a<R@a<�Ba<�Fa<6La<�Ra<�Ya<�`a<Zga<ma<hqa<�ta<�ua<"va<�ta<�ra<epa<�ma<�ja<�ha<�ga<	ga<�ga<�ha<�ja<�ma<{pa<-sa<�  �  Qwa<2xa<~wa<�ua<ra<?ma<(ga<`a<�Xa<�Pa<Ja<Da<�?a<7=a<�<a<u>a<�Aa<Ga<zNa<HVa<�^a<�fa<sna<�ta<Qza<~a<��a<��a<C�a<{�a<�~a<F}a<�{a<�za<lza<�za<=|a<G~a<�a<܃a<�a<��a<Q�a<m�a<Ћa<�a<��a<�a<�{a<Uua<=na<Gga<+aa<�[a<�Xa<LWa<�Wa<�Za<(_a<�ea<ma<uua<�}a<�a<��a<��a<��a<śa<ȝa<��a<_�a<�a<��a<*�a<Y�a<#�a<��a<�a<�a<��a<�a<!�a<��a<.�a<3�a<�a<_�a<f�a<��a<�a<�a<��a<�{a<>ta<�ma<gha<6ea<�ca<Tda<ga<}ka<�qa<�xa<ڀa<��a<�a<��a<Лa<��a<��a<�a<m�a<H�a<)�a<�a<��a<јa<��a<�a<c�a<i�a<�a<4�a<B�a<^�a<u�a<�a<�a<Ϟa<��a<ƕa<O�a<ۇa<�a<�wa<�pa<ja<;ea<?ba<&aa<mba<bea<Sja<�pa<�wa<�a<$�a<#�a<�a<��a<��a<u�a<��a<��a<�a<��a<Q�a<�a<�a<��a<\�a<Ґa<��a<��a<a�a<T�a<Ϙa<r�a<Z�a<��a<��a<��a<��a<q�a<hza<�qa<�ia<ba<c[a<�Va<�Sa<Sa<vTa<iWa<}\a<�ba<�ia<�pa<�wa<�}a<{�a<?�a<5�a<�a<*�a<y�a<�a<�a<O~a<�{a<�ya<xa<�wa<�wa<�xa<�za<|a<�}a<�~a<?a<�~a<F|a<�xa<�sa<Nma<�ea<�]a<vUa<�Ma<�Fa<�@a<U=a<X;a<�;a<>a<2Ba<7Ha<Oa<�Va<P^a<~ea<�ka<�pa<�ta<�va<�wa<�va<�ua<�sa<Cqa<oa</ma<la<uka<la<.ma<oa<Vqa<�sa<�ua<�  �  �xa<�xa<�wa<�ua<�qa<�la<�ea<�^a<�Va<�Na<�Ga<bAa<�<a<�9a<}9a<-;a<;?a<�Da<La<1Ta<�\a<iea<[ma<rta<za<K~a<��a<��a<ǂa<#�a<݀a<�a<[~a<�}a<T}a<�}a<a<�a<p�a<�a<��a<�a<��a<�a<.�a<��a<<�a<�a<�za<�sa<,la<ea<�^a<cYa<�Ua<Ta<�Ta<�Wa<�\a<�ba<�ja<^sa<H|a<ʄa<��a<E�a<z�a<�a<L�a<*�a<��a<��a<4�a<��a< �a<�a<��a<ӗa<Ęa<^�a<N�a<S�a<K�a<��a<:�a<��a<��a<0�a<O�a<��a<��a<��a<�ya<�qa<ka<�ea<�aa<l`a<aa<da<�ha<Boa<�va<�~a<+�a<�a<ܕa<��a<��a<a�a<ƣa<ɣa<�a<�a<-�a<<�a<��a<v�a<�a<=�a<4�a<��a<{�a<=�a<��a<ޢa<ڢa<y�a<�a<��a<!�a<!�a<a�a<�}a<�ua<na<fga<\ba<�^a<�]a<$_a<�ba<�ga<Ona<�ua<�}a<��a<
�a<u�a<c�a<�a<�a<��a<1�a<ǜa<��a<��a<��a<��a<ɓa<g�a<��a<��a<�a<��a<!�a<g�a<��a<��a<��a<i�a<]�a<�a<*�a<�xa<�oa<bga<e_a<�Xa<�Sa<�Pa<�Oa<EQa<�Ta<�Ya<Y`a<sga<oa<2va<�|a<�a<�a<��a<��a<V�a<�a<υa<K�a<��a<]~a<`|a< {a<�za<�za<�{a<�|a<>~a<�a<d�a<G�a<�~a<|a<�xa<!sa<Dla<wda< \a<dSa<IKa<�Ca<D>a<:a<*8a<u8a<";a<�?a<�Ea<�La<�Ta<�\a<Eda<ka<�pa<�ta<wa<Xxa<Bxa<Hwa<pua<�sa<�qa<�oa<�na<�na<�na<�oa<�qa<�sa<�ua<�wa<�  �  �}a<�}a<m|a<$ya<�sa<�la<qca<^Ya<wNa<�Ca<�9a<M1a<�*a<'a<�&a<d(a<�-a<-5a<�>a<�Ia<HUa<�`a<fka<�ta<h|a<7�a<ʅa<��a<��a<�a<��a<��a<��a<�a<Y�a<�a<H�a<��a<Q�a<��a<��a<U�a<�a<%�a<�a<]�a<��a<��a<�wa<�ma<�ca<�Ya<`Pa<OIa<�Ca<�Aa<xBa<�Ea<_La<�Ta<]_a<�ja<�va<	�a<Z�a<?�a<%�a<I�a<��a<2�a<֤a<X�a<��a<�a<M�a<�a<A�a<|�a<̜a<��a<Πa<��a<��a<��a<�a<��a<I�a<B�a<��a<�a<�a<{a<8pa<�ea<4\a<�Ta<�Oa<Na<�Na<�Ra<=Ya<�aa<0la<wa<<�a<��a<>�a<�a<��a<��a<>�a<��a<]�a<m�a<�a<}�a<��a<�a<��a<ϝa<�a<ݠa<-�a<��a<c�a<��a<V�a<��a<�a<=�a<��a<5�a<��a<lva<rka<�`a<�Wa<Qa<�La<�Ka<�La<�Qa<�Xa<�aa<la<�va<ˁa<��a<~�a<B�a<]�a<8�a<Q�a<�a<#�a< �a<$�a<a<ؘa<\�a<��a<l�a<��a<p�a<ʜa<��a< �a<��a<��a<	�a<-�a<y�a<͈a<�~a<Bsa<�ga<\a<PQa<�Ha<�Aa<K>a<x=a<A?a<kDa<XKa<�Ta<�^a<�ha<sa<�{a<��a<;�a<(�a<��a<��a<M�a<Ċa<��a<��a<ށa<�a< ~a<�}a<!~a<-a<��a<�a<Y�a<��a<p�a<Ӄa<��a<{a<�sa<�ja<C`a<�Ta<tIa<Y>a<�4a<�,a<V'a<;%a<�%a<)a<N/a<}7a<�Aa<<La<1Wa<waa<�ja<?ra<�wa<�{a< }a<f}a<|a<za<�wa<ua<2sa<�qa<Rqa<�qa<0sa<ua<�wa<:za<P|a<�  �  #}a<�}a<3|a<ya<�sa<�la<da<7Za<tOa<�Da<�:a<~2a<4,a<c(a<�'a<�)a<�.a<j6a<�?a<�Ja<>Va<�aa<la<@ua<�|a<�a<~�a<'�a<?�a<?�a<��a<��a<݀a<�a<=a<�a<�a<^�a<S�a<��a<ڌa<��a<i�a<ܑa<��a<b�a<<�a<!�a<�xa<�na<�da<�Za<�Qa<dJa<XEa<�Ba<�Ca<&Ga<xMa<Va<``a<�ka<owa<��a<Ռa<��a<:�a<�a<��a<��a<"�a<��a<j�a<(�a<�a<��a<#�a<c�a<v�a<l�a<�a<��a< �a<Ǧa<~�a<��a<�a<k�a<�a<t�a<ʆa<�{a<qa<�fa<q]a<&Va<;Qa</Oa<Pa<�Sa<bZa<�ba<ma<xa<�a<e�a<��a<�a<��a<>�a<�a<�a<��a<��a<��a<n�a<C�a<ݜa<X�a<��a<ѝa<ȟa<1�a<��a<��a<�a<�a<e�a<�a<c�a<�a<یa<��a<iwa<Ola<�aa<Ya<SRa<Na<�La<RNa<�Ra<�Ya<�ba<�la<�wa<��a<=�a<˔a<j�a<+�a<�a<٣a<2�a<n�a<��a<;�a<��a<��a<@�a<וa<9�a<��a<q�a<��a<ʝa<k�a<�a<<�a<��a<2�a<��a<>�a<Ba<ta<sha<]a<�Ra<�Ia<QCa<u?a<�>a<�@a<�Ea<�La<�Ua<u_a<�ia<�sa<z|a<�a<Q�a<Ìa<]�a</�a<��a<��a<׆a<��a<��a<_~a<}a<y|a<�|a<~a<�a<ҁa<��a<̈́a<�a<��a<N�a<+{a<%ta<'ka<�`a<�Ua<NJa<k?a<�5a<.a<�(a<K&a<�&a<_*a<s0a<�8a<�Ba<5Ma<Xa< ba<ka<fra<�wa<A{a<�|a<�|a<\{a<(ya<�va<ta<�qa<�pa<%pa<�pa<�qa<ta<�va<Eya<�{a<�  �  c{a<g|a<�{a<ya<ata<�ma<�ea<\a<�Qa<�Ga<T>a<*6a<0a<�,a<�+a<.a<�2a<:a<FCa<�Ma<�Xa<fca<nma<va<�|a<�a<΄a<�a<i�a< �a<��a<�a<_}a<�{a<P{a<�{a<J}a<�a<�a<��a<v�a<��a<�a<�a<�a<��a<׈a<C�a<"za<�pa<4ga<�]a<EUa<Na<}Ia<(Ga<�Ga<YKa<'Qa<�Ya<�ca<fna<�ya<Y�a<�a<.�a<��a<��a<�a<0�a<3�a<@�a<n�a<��a<|�a<ٖa<�a<l�a<��a<�a<ʜa<��a<Ӣa<�a<1�a<�a<ͣa<ԟa<��a<ˑa<{�a<Y~a<�sa<�ia< aa<�Ya<wUa<CSa<ITa<�Wa<^a<wfa<pa<�za<	�a<�a<��a<��a<ţa<��a<�a<:�a<��a<�a<�a<�a<��a<�a<B�a<Șa<�a<_�a< �a<�a<��a<0�a<�a<ɥa<�a<�a<��a<Z�a<v�a<�ya<2oa<iea<�\a<<Va<?Ra<�Pa<�Ra<�Va<}]a<fa<�oa<3za<J�a<��a<��a<ڛa<	�a<<�a<��a<\�a<O�a<�a<&�a<"�a<��a<T�a<Ƒa<m�a<֓a<6�a<��a<f�a<u�a<|�a<k�a</�a<n�a<Q�a<`�a<ڀa<8va<ka<`a<6Va<�Ma<vGa<�Ca<�Ba<�Da<4Ia<EPa<�Xa<"ba<�ka<Sua<�}a<��a<��a<_�a<��a<��a<��a<��a<ۃa<o�a<}a<�za<�xa<�xa<�xa<�za<�|a<�~a<v�a<�a<��a<˂a<�a<�{a<�ta<~la<�ba<Xa<Ma<�Ba<s9a<�1a<�,a<^*a<+a<[.a<4a<9<a<zEa<�Oa<�Ya<�ca<la<�ra<�wa<�za<�{a<{a<\ya<�va<�sa<�pa<-na<�la<la<�la<na<�pa<�sa<�va<�ya<�  �  �xa<rza<|za<�xa<ua<�oa< ha<a_a<�Ua<qLa<�Ca<�;a<%6a<�2a<.2a</4a<�8a<�?a<]Ha<4Ra<�\a<�fa<�oa<�wa<o}a<��a<y�a<ԃa<��a<N�a<j}a<vza<�wa<va<Aua<�ua<xwa<za<�}a<�a<^�a<S�a<u�a<K�a<c�a<��a<ȉa<D�a<�|a<tta<�ka<�ba<�Za<Ta<�Oa<�Ma<)Na<eQa<8Wa<_a<qha<�ra<=}a<0�a<%�a<?�a<��a<�a<=�a<Ԡa<��a<6�a<��a<��a<�a<�a<�a<R�a<�a<P�a<��a<P�a<�a<�a<�a<}�a<h�a<&�a<��a<�a<��a<"�a<cxa<�na<�fa<`a<�[a<�Ya<�Za<�]a<�ca<�ka<�ta<�~a<j�a<��a<f�a<\�a<��a<��a<
�a<��a<�a<��a<%�a<��a<�a<�a<0�a<˒a<i�a<��a<;�a<��a<��a<��a<�a<��a<��a<��a<��a<�a<��a<�}a<�sa<�ja<�ba<F\a<�Xa<GWa<�Xa<�\a<ca<+ka<cta<~a<i�a<�a<�a<K�a<��a<�a<��a<��a<}�a<їa<�a<��a<�a<D�a<��a<��a<?�a<�a<�a<N�a<�a<�a<��a<~�a<p�a<A�a<`�a<��a<�ya<boa<ea<�[a<�Sa<|Ma<Ja<(Ia<�Ja<DOa<�Ua<�]a<�fa<�oa<+xa<�a<��a<��a<Ћa<�a<d�a<o�a<��a<ma<2{a<vwa<�ta<�ra<ira<Gsa<�ta<�wa<�za<�}a<�a<r�a<W�a<�a<�{a<2va<�na<�ea<�[a<�Qa<�Ga< ?a<�7a<3a<�0a<X1a<a4a<�9a<Aa<LJa<�Sa<^]a<Hfa<�ma<�sa<�wa<�ya<�ya<uxa<�ua<`ra<�na<Uka<�ha<�fa< fa<�fa<|ha<6ka<�na<]ra<�ua<�  �  Bua<�wa<2ya<�xa<�ua<kqa<ka<�ca<[a<�Ra<KJa<�Ca<Q>a<);a<�:a<j<a<�@a<'Ga<Oa<Xa<laa<|ja<yra<5ya<�}a<�a<߁a<�a<�~a<]{a<�wa<�sa<�pa<Dna<;ma<�ma<^oa<�ra<�va<�{a<�a<�a<M�a<�a<{�a<��a<�a<�a<J�a<ya<�pa<�ha<�aa<�[a<�Wa<�Ua<�Va<�Ya<&_a<5fa<�na<Mxa<�a<��a<x�a<��a<Ϝa<�a<'�a<ŝa<Қa<��a<�a<ʎa<j�a<
�a<�a<S�a<�a<��a<�a<��a<ޙa<�a<.�a<��a<¢a<��a<��a<��a<^�a<�a<~a<�ua<na<ha<�ca<@ba<�ba<)fa<�ka<�ra<�za<ڃa<��a<��a<e�a<]�a<r�a<��a<��a<I�a<��a<H�a<��a<��a<=�a<��a<E�a<��a<��a<a<��a<*�a<O�a<�a<w�a<b�a<k�a<h�a<��a<Փa<��a<�a<za<bqa<-ja<uda<�`a<�_a<�`a<�da<�ja<�qa<@za<��a<d�a<��a<Ęa<ۜa<*�a<O�a<͝a<ƚa<��a<!�a<j�a<Q�a<+�a<=�a<��a<��a<��a<�a<�a<��a<֕a<�a<u�a<��a<��a<��a<��a<�a<N~a<�ta<cka<�ba<d[a<�Ua<lRa<�Qa<Sa<2Wa<�\a<da<
la<;ta<�{a<�a<�a<�a<��a<ىa<U�a<L�a<d~a<[ya<Eta<�oa<�la<�ja<jja<\ka<�ma<�pa<�ta<�xa<|a<�~a<�a<a<N|a<�wa<Wqa<�ia<�`a<VWa<TNa<VFa<�?a<K;a<X9a<�9a<�<a<�Aa<NHa<vPa<Ya<�aa<\ia<�oa<�ta<�wa<�xa<�wa<ua<Cqa<�la<dha<1da<�`a<�^a<^a<�^a<�`a<da<7ha<�la<>qa<�  �  �pa<�ta<nwa<&xa<�va<�sa<�na<Pha<�`a<�Ya<YRa<La<~Ga<�Da<6Da<�Ea<�Ia<�Oa<�Va<�^a<ga<�na<�ua<,{a<�~a<C�a<�a<�}a<za<�ua<�pa<la<,ha<;ea<�ca<=da<#fa<�ia<�na<|ta<�za<�a<C�a<x�a<�a<Ǎa<��a<�a<;�a<!~a<wa<apa<�ia<�da<aa<�_a<)`a<ca<�ga<�na<qva<�~a<�a<Ԏa</�a<4�a<�a<�a<��a<ߙa<Еa<�a<��a<ʆa<ςa<�a<�~a<�~a<�a<��a<�a<i�a<�a<D�a<��a<��a<ۡa<'�a<r�a<��a<��a<v�a<��a<T}a<nva<�pa<Uma<�ka<�la<qoa<<ta<�za<'�a<̉a<��a<E�a<��a<��a</�a<�a<��a<��a<3�a<��a<8�a<_�a<d�a<��a<ˀa<h�a<��a<�a<&�a<{�a<ؖa<��a<F�a<��a<�a<g�a<Ŝa<R�a<��a<߈a<�a<rya<�ra<�ma<`ja<Tia<�ja<�ma<sa<�ya<�a<��a<܏a<�a<��a<��a<m�a<P�a<N�a<�a<ܐa<,�a<��a<�a<!}a<�za<Sza<E{a<~a<ځa<��a<͋a<��a<ڔa<՗a<8�a<��a<��a<2�a<�a<m�a<�za<�ra<�ja<da<_a< \a<([a<�\a<�_a<ea<�ka<Tra<xya<�a<քa<��a<$�a<ɉa<p�a<q�a<K~a<Xxa<ra<Fla<bga<�ca<�aa<aa<Eba<%ea< ia<�ma<�ra<Iwa<�za<w}a<$~a<�|a<�ya<Xta<�ma<%fa<�]a<Va<�Na<�Ha<�Da<�Ba<;Ca<�Ea<IJa<nPa<�Wa<�^a<�fa<�la<Ara<�ua<Zwa<�va<�ta<�pa<�ka<mfa<�`a<\a<Xa<pUa<�Ta<ZUa<�Wa<�[a<�`a<-fa<�ka<�  �  #la<}qa<lua<zwa<�wa<�ua<:ra<4ma<(ga<�`a<�Za<TUa<NQa<�Na<tNa<Pa<�Sa<�Xa<�^a<�ea<�la<�sa<ya<	}a<"a<Fa<�}a< za<$ua<Xoa<Wia<�ca<�^a<m[a<�Ya<�Ya<:\a<G`a<�ea<�la<�sa<M{a<�a<��a<��a<��a<��a<ߋa<E�a<p�a<�}a<�wa<�ra<na<ka<�ia<bja<ma<nqa<Twa< ~a<e�a<��a<��a<(�a<��a<��a<u�a<��a<ŕa<O�a<%�a<ރa<~a<Bya<�ua<Qta<�ta<wa<{a<��a<�a<��a<!�a<Ǚa<+�a<��a<i�a<#�a<��a<,�a<@�a<��a<F�a<ka<�za<�wa<va<�va<Qya<�}a<-�a<��a<7�a<��a<�a<(�a<\�a<��a<
�a<|�a<o�a<G�a<��a</�a<Wa<�za<�wa<mva<Swa<za<]~a<�a<D�a<ːa<�a<��a<��a<V�a< �a<�a<�a<��a<"�a<T�a<ׁa<�{a<vwa<�ta<�sa<�ta<�wa<|a<ʁa<�a<��a<|�a<O�a<��a<�a<q�a<�a<��a<�a<��a<��a<I}a<�wa<Ssa<�pa<�oa<Zqa<ita<ya<�~a<�a<�a<��a<��a<��a<]�a<�a<��a<��a<��a<��a<_za<�sa<�ma<ia<7fa<aea<�fa<{ia<�ma<Hsa<#ya<�~a<��a<Їa<�a<�a<W�a<��a<Xa<�xa<�qa<Oja<�ca<�]a<�Ya<4Wa<�Va<mXa<�[a<�`a<+fa<8la<&ra<3wa<{a<�|a<$}a<T{a<�wa<Vra<�ka<�da<^a<�Wa<�Ra<�Na<!Ma<vMa<�Oa<�Sa<�Xa<�^a<iea<�ka<�pa<�ta<�va<�va<ua<dqa<>la<fa<S_a<�Xa< Sa<]Na<jKa<DJa<HKa<Na<�Ra<~Xa<�^a<�ea<�  �  Pga<�ma<Gsa<�va<]xa<�wa<�ua<�qa<Dma<ha<�ba<^a<
[a<Ya<�Xa<Za<@]a<�aa<�fa<�la<�ra<xa<|a<�~a<�a<Y~a<{a<%va<pa<�ha<�aa<*[a<�Ua<�Qa<zOa<�Oa<Ra<�Va<�\a<�da<ma<�ua<�}a<c�a<��a<f�a<��a<e�a<�a<��a<O�a<�a<{a<�wa<�ta<ta<�ta<�va<�za<�a<ƅa<�a<��a<��a<Кa<�a<��a<	�a<�a<��a<Ɋa<H�a< |a<=ua<�oa<�ka<ja<�ja<!ma<�qa<�wa<\a<�a<�a<͕a<}�a<��a<��a<ˡa<�a<{�a<��a<��a</�a<P�a<M�a<r�a<i�a<�a<�a<Ԇa<}�a<�a<x�a<��a<��a<c�a<E�a<3�a<�a<��a<��a<>�a<��a<�|a<2va<�pa<vma<,la<ma<9pa<'ua<�{a<�a<��a<�a<[�a<v�a<��a<�a<�a<`�a<W�a<@�a<��a<�a<%�a<4�a<�~a<�}a<�~a<H�a<�a<ʉa<)�a<e�a<�a<`�a<f�a<o�a<��a<��a<ܒa<�a<�a<Q|a<�ta<Cna<nia<zfa<�ea<8ga<�ja<pa<�va<�}a<a�a<<�a<��a<�a<1�a<V�a<~�a<Ԓa<�a<*�a<�a<|a<�va<�ra<pa<�oa<tpa< sa<�va<�za<�a<S�a<��a<y�a<B�a<�a<�a<��a<{a<Fsa<�ja<�ba<�Za<CTa<�Oa<�La<�La<zNa<LRa<�Wa<�^a<�ea<�la<8sa<Sxa<�{a<j}a<�|a<�za<�va<�qa<�ka<�ea<�`a<)\a<�Xa<{Wa<�Wa<uYa<�\a<9aa<_fa<�ka<pa<Rta<�va<�wa<`va< sa<�ma<�ga<�_a<2Xa<�Pa<�Ia<�Da<9Aa<@a<Aa<VDa<pIa<)Pa<�Wa<�_a<�  �  �ba<uja<%qa<�ua<�xa<�ya<�xa<xva<�ra<�na<�ja<�fa<�ca<`ba<Eba<aca<	fa<�ia<lna<^sa<xa<A|a<
a<h�a<�a<"}a<�xa<mra<ka<�ba<�Za<�Ra<�La<9Ha<�Ea<Fa<�Ha<�Ma<�Ta<]a<|fa<*pa<bya<w�a<.�a<�a<ۏa<��a<ԏa<��a<,�a<��a<��a<�a<~a<_}a<~a<�a<��a<�a<�a<�a<�a<Қa<!�a<�a<��a<j�a<'�a<f�a<y�a<�|a<�ta<�la<�fa<dba<�`a<�`a<�ca<ia<�oa<xa<ڀa<։a<�a<��a<O�a<��a<=�a<��a<��a<$�a<��a<��a<f�a<�a<��a<܉a<@�a<�a<2�a<5�a<Зa<�a</�a<�a<S�a<�a<b�a<�a<��a<5�a<��a<�}a<ua<�ma<�ga<�ca<�ba<�ca<ga<�la<�sa<|a<Ԅa<p�a<�a<S�a<��a<b�a<�a<��a<ܞa<ǚa<]�a<��a<u�a<)�a<�a<k�a<��a<�a<=�a<F�a<��a<��a<2�a<P�a<��a<��a<Q�a<�a<%�a<�a<~a<ua<�la<�ea<`a<�\a</\a<�]a<�aa<�ga<oa<fwa<�a<��a<юa<D�a<��a<P�a<��a<��a<͒a<�a<�a<�a<ya<|a<�ya<ya<�ya<�{a<�~a<9�a<Ѕa<G�a<Ћa<ʌa<c�a<��a<N�a<�~a<�va<�ma<Zda<�Za<fRa<|Ka<Fa<gCa<Ca<Ea<�Ia<�Oa<JWa<{_a<�ga<Yoa<�ua<�za<m}a<k~a<I}a<�za<�va<)ra<Rma<�ha<�da<$ba<�`a<�`a<vba<:ea<�ha<Dma<Lqa<"ua<�wa<�xa<Exa<�ua<qa<�ja<ca<TZa<aQa<�Ha<hAa<�;a<�7a<w6a<�7a<6;a<�@a<(Ha<�Pa<�Ya<�  �  �^a<�ga<Hoa<ua<7ya<!{a<e{a<za<�wa<Zta<qa<na<�ka<lja<.ja<|ka<�ma<�pa<�ta<�xa<�|a<�a<b�a<|�a<�a<|a<�va<Eoa<�fa<�]a<yTa<'La<!Ea<@a<�=a<�=a<c@a<�Ea<XMa<Va<�`a<dka<�ua<�~a<��a<��a<��a<k�a<��a<v�a<I�a<��a<ǉa<g�a<��a<W�a<	�a<�a<�a<ˎa<�a<F�a<��a<ӝa<%�a<͞a<c�a<�a<őa<��a<ǀa<Xwa<na<�ea<�^a<6Za<Xa<�Xa<�[a<2aa<�ha<�qa<�{a<X�a<��a<ɖa<�a<��a<5�a<�a<ӣa<}�a<T�a<ٚa<v�a<��a<ϒa<Αa<K�a<�a<v�a<ҙa<t�a<��a<ڣa<��a<إa<e�a<��a<H�a<�a<+�a<��a<�wa<jna<=fa<�_a<�[a<Za<D[a<�^a<ea<�la<va<�a<G�a<�a<v�a<��a<��a<J�a<.�a<h�a<��a<�a<1�a<��a<�a<�a<W�a<�a<��a<]�a<��a<�a<,�a<��a<��a<�a<��a<=�a<�a<��a<��a<�xa<�na<�ea<�]a<�Wa<�Ta<�Sa<�Ua<�Ya<o`a<�ha<�qa<'{a<.�a<U�a<��a<U�a<�a<��a<n�a<��a<#�a<��a<��a<چa<��a<Ӂa<	�a<��a<�a<d�a<:�a<�a<X�a<юa<ώa<,�a<�a<Ճa<||a<Vsa<Fia<�^a<vTa<@Ka<�Ca<�=a<�:a<�:a<�<a<�Aa<�Ha<�Pa<)Za<[ca<la<�sa<Yya<k}a<ba<�a<�}a<#{a<�wa<�sa<�oa<sla<@ja<�ha<�ha<Hja<}la<�oa<�ra<,va<�xa<hza<_za<�xa<�ta<Toa<�ga<�^a<bUa<yKa<Ba<�9a<w3a<u/a<�-a<A/a<3a<^9a<pAa<�Ja<�Ta<�  �  C[a<ea<�ma<�ta<{ya<L|a<b}a<�|a<;{a<�xa< va<qsa<cqa<npa<@pa<gqa<Esa<>va<�ya<�|a<�a<�a<<�a<a�a<�a<?{a<�ta<�la<Nca<}Ya<�Oa<�Fa<;?a<:a<87a<'7a<J:a<�?a<�Ga<�Qa<R\a<�ga<�ra<�|a<Y�a<J�a<��a<�a<�a<��a<:�a<�a<��a<��a<��a<s�a<$�a<ݍa<��a<�a<s�a<H�a<*�a<#�a< a<N�a<>�a<Ζa<��a<ކa<!}a<�ra<ia<F`a<�Xa<&Ta<�Qa<+Ra<�Ua<6[a<lca<�la<Ewa<ցa<�a<הa<2�a<��a<��a<��a<H�a<�a<u�a<{�a<Üa<3�a<��a<�a<X�a<��a<��a<۞a<��a<Ťa<��a<��a<�a<��a<A�a<��a<��a< �a<�}a<sa<Fia<�`a<�Ya<zUa<�Sa<Ua<�Xa<Q_a<�ga<Tqa<�{a<�a<��a<̗a<]�a<��a<u�a<,�a<�a<9�a<)�a<"�a<�a<��a<�a<j�a<�a<S�a<��a<^�a</�a<��a<�a<��a<��a<ٞa<p�a<6�a<T�a<Ga<�ta<	ja<q`a<�Wa<�Qa<7Na<9Ma<gOa<�Sa<�Za<�ca<:ma<jwa<1�a<�a<n�a<�a<n�a<�a<��a<ʙa<�a<K�a<�a<o�a<��a<�a<#�a<b�a<��a<��a<��a<�a<��a<"�a<l�a<��a<Z�a<��a<Lza<tpa<�ea<\Za<�Oa<�Ea<q=a<�7a<�4a<F4a<�6a<�;a<[Ca<La<�Ua<�_a<Nia<�qa<txa<q}a<#�a<S�a<k�a<�~a<�{a<0xa<ua<	ra<pa<�na<oa<�oa<�qa<�ta<,wa<�ya<�{a<v|a<�{a<ya<qta<�ma<�ea<�[a<yQa<�Fa<�<a<C4a<j-a<C)a<{'a<)a<-a<�3a<@<a<Fa<�Pa<�  �  mYa<�ca<�la<ta<�ya<�|a<�~a<y~a<H}a<P{a<ya<�va<+ua<Qta<Tta<3ua<�va<�ya<�|a<{a<�a<��a<3�a<�a<�a<�za<�sa<ka<Taa<�Va<�La<=Ca<�;a<6a<3a<3a<6a<�;a<#Da<DNa<�Ya<Wea<�pa<i{a<��a<�a<<�a<��a<G�a<a�a<n�a<דa<�a<��a<��a<n�a<)�a<��a<&�a<1�a<l�a<��a<�a<��a<��a<��a<�a<$�a<\�a<;�a<�za<2pa<�ea<�\a<#Ua<�Oa<~Ma<�Ma<sQa<�Wa<�_a<�ia<�ta<�a<R�a<��a<��a<��a<u�a<��a<ۧa<ަa<�a<�a<�a<�a<x�a<�a<A�a<j�a<o�a<�a<��a<ߦa<x�a<�a<˧a<Фa<͟a<�a<$�a<?�a<G{a<Kpa<�ea<�\a<�Ua<;Qa<�Oa<�Pa<�Ta<�[a<Kda<xna<Nya<1�a<�a<�a<��a<�a<�a<M�a<ߦa<G�a<�a<3�a<��a<\�a<�a<�a<әa<�a<�a<j�a<��a<��a<��a<|�a<��a<��a<�a<.�a<ɇa<L}a<ra<ga<�\a<PTa<�Ma< Ja<"Ia<+Ka<	Pa<9Wa<H`a<xja<ua<�a<��a<��a<��a<��a<��a<��a<��a<G�a<<�a<�a<��a<~�a<�a<)�a<6�a<4�a<ʍa<��a<M�a<o�a<��a<*�a<�a<�a<
�a<ya<�na<bca<�Wa<YLa<Ba<�9a<�3a<d0a<0a<�2a<,8a<�?a<
Ia<JSa<�]a<�ga<�pa<�wa<=}a<��a</�a<��a<��a<~a<3{a<Ixa<�ua<�sa<�ra<�ra<�sa<uua<�wa<�ya<|a<k}a<�}a<R|a<*ya<�sa<�la<da<Za<
Oa<Da<�9a<�0a<�)a<%a<i#a<�$a< )a<�/a<�8a<3Ca<GNa<�  �  �Xa<�ba<ola<�sa<�ya<&}a<�~a<5a<�}a<M|a<za<�wa<{va<vua<ua<Yva<Bxa<�za<�}a<`�a<Ăa<o�a<}�a<9�a<�a<�za<Rsa<bja<x`a<�Ua<�Ka<Ba<n:a<�4a<�1a<�1a<�4a<�:a<�Ba<5Ma<�Xa<rda<>pa<�za<Q�a<��a<��a<��a<Ζa<�a<%�a<�a<��a<��a<ڐa<��a<D�a<��a<O�a<�a<��a<N�a<Ǡa<�a<ҡa<�a<ʛa<֕a<܍a<��a<za<Zoa<�da<Y[a<Ta<�Na<eLa<�La<Pa<tVa<�^a<�ha<�sa<�~a<��a<P�a<e�a<��a<ӥa<ԧa<�a<��a<��a<��a<�a<"�a<��a<�a<`�a<��a<��a<ݢa<��a<��a<8�a<]�a<�a<��a<��a<��a<��a<w�a<Lza<moa<�da<�[a<�Ta<�Oa<tNa<kOa<�Sa<mZa<,ca<�ma<Pxa<\�a<t�a<��a<��a<�a<O�a<��a<��a<��a<�a<*�a<��a<��a<'�a<��a<��a<R�a<�a<v�a<��a<a�a<e�a<Ǥa<Ԣa<Ğa<��a<ʐa<�a<q|a<"qa<+fa<�[a</Sa<�La<�Ha<Ha<�Ia<�Na<�Ua<9_a<�ia<4ta<�~a<3�a<f�a<��a< �a<�a<��a<b�a<��a<R�a<�a<"�a<Ҏa<�a<D�a<��a<]�a<��a<��a<�a<"�a<�a<|�a<h�a<�a<��a<�xa<na<�ba<�Va<SKa<�@a<�8a<<2a<K/a<�.a<l1a<7a<~>a<Ha<`Ra<�\a<ga<$pa<�wa<@}a<��a<y�a<��a<7�a<�~a<L|a<Mya<�va<ua<$ta<ta<ua<�va<�xa< {a<�|a<*~a<~a<�|a<Pya<�sa<�la<qca<MYa<Na<$Ca<x8a<Z/a<W(a<�#a<U"a<j#a<�'a<�.a<�7a<UBa<IMa<�  �  mYa<�ca<�la<ta<�ya<�|a<�~a<y~a<H}a<P{a<ya<�va<+ua<Qta<Tta<3ua<�va<�ya<�|a<{a<�a<��a<3�a<�a<�a<�za<�sa<ka<Taa<�Va<�La<=Ca<�;a<6a<3a<3a<6a<�;a<#Da<DNa<�Ya<Wea<�pa<i{a<��a<�a<<�a<��a<G�a<a�a<n�a<דa<�a<��a<��a<n�a<)�a<��a<&�a<1�a<l�a<��a<�a<��a<��a<��a<�a<$�a<\�a<;�a<�za<2pa<�ea<�\a<#Ua<�Oa<~Ma<�Ma<sQa<�Wa<�_a<�ia<�ta<�a<R�a<��a<��a<��a<u�a<��a<ۧa<ަa<�a<�a<�a<�a<x�a<�a<A�a<j�a<o�a<�a<��a<ߦa<x�a<�a<˧a<Фa<͟a<�a<$�a<?�a<G{a<Kpa<�ea<�\a<�Ua<;Qa<�Oa<�Pa<�Ta<�[a<Kda<xna<Nya<1�a<�a<�a<��a<�a<�a<M�a<ߦa<G�a<�a<3�a<��a<\�a<�a<�a<әa<�a<�a<j�a<��a<��a<��a<|�a<��a<��a<�a<.�a<ɇa<L}a<ra<ga<�\a<PTa<�Ma< Ja<"Ia<+Ka<	Pa<9Wa<H`a<xja<ua<�a<��a<��a<��a<��a<��a<��a<��a<G�a<<�a<�a<��a<~�a<�a<)�a<6�a<4�a<ʍa<��a<M�a<o�a<��a<*�a<�a<�a<
�a<ya<�na<bca<�Wa<YLa<Ba<�9a<�3a<d0a<0a<�2a<,8a<�?a<
Ia<JSa<�]a<�ga<�pa<�wa<=}a<��a</�a<��a<��a<~a<3{a<Ixa<�ua<�sa<�ra<�ra<�sa<uua<�wa<�ya<|a<k}a<�}a<R|a<*ya<�sa<�la<da<Za<
Oa<Da<�9a<�0a<�)a<%a<i#a<�$a< )a<�/a<�8a<3Ca<GNa<�  �  C[a<ea<�ma<�ta<{ya<L|a<b}a<�|a<;{a<�xa< va<qsa<cqa<npa<@pa<gqa<Esa<>va<�ya<�|a<�a<�a<<�a<a�a<�a<?{a<�ta<�la<Nca<}Ya<�Oa<�Fa<;?a<:a<87a<'7a<J:a<�?a<�Ga<�Qa<R\a<�ga<�ra<�|a<Y�a<J�a<��a<�a<�a<��a<:�a<�a<��a<��a<��a<s�a<$�a<ݍa<��a<�a<s�a<H�a<*�a<#�a< a<N�a<>�a<Ζa<��a<ކa<!}a<�ra<ia<F`a<�Xa<&Ta<�Qa<+Ra<�Ua<6[a<lca<�la<Ewa<ցa<�a<הa<2�a<��a<��a<��a<H�a<�a<u�a<{�a<Üa<3�a<��a<�a<X�a<��a<��a<۞a<��a<Ťa<��a<��a<�a<��a<A�a<��a<��a< �a<�}a<sa<Fia<�`a<�Ya<zUa<�Sa<Ua<�Xa<Q_a<�ga<Tqa<�{a<�a<��a<̗a<]�a<��a<u�a<,�a<�a<9�a<)�a<"�a<�a<��a<�a<j�a<�a<S�a<��a<^�a</�a<��a<�a<��a<��a<ٞa<p�a<6�a<T�a<Ga<�ta<	ja<q`a<�Wa<�Qa<7Na<9Ma<gOa<�Sa<�Za<�ca<:ma<jwa<1�a<�a<n�a<�a<n�a<�a<��a<ʙa<�a<K�a<�a<o�a<��a<�a<#�a<b�a<��a<��a<��a<�a<��a<"�a<l�a<��a<Z�a<��a<Lza<tpa<�ea<\Za<�Oa<�Ea<q=a<�7a<�4a<F4a<�6a<�;a<[Ca<La<�Ua<�_a<Nia<�qa<txa<q}a<#�a<S�a<k�a<�~a<�{a<0xa<ua<	ra<pa<�na<oa<�oa<�qa<�ta<,wa<�ya<�{a<v|a<�{a<ya<qta<�ma<�ea<�[a<yQa<�Fa<�<a<C4a<j-a<C)a<{'a<)a<-a<�3a<@<a<Fa<�Pa<�  �  �^a<�ga<Hoa<ua<7ya<!{a<e{a<za<�wa<Zta<qa<na<�ka<lja<.ja<|ka<�ma<�pa<�ta<�xa<�|a<�a<b�a<|�a<�a<|a<�va<Eoa<�fa<�]a<yTa<'La<!Ea<@a<�=a<�=a<c@a<�Ea<XMa<Va<�`a<dka<�ua<�~a<��a<��a<��a<k�a<��a<v�a<I�a<��a<ǉa<g�a<��a<W�a<	�a<�a<�a<ˎa<�a<F�a<��a<ӝa<%�a<͞a<c�a<�a<őa<��a<ǀa<Xwa<na<�ea<�^a<6Za<Xa<�Xa<�[a<2aa<�ha<�qa<�{a<X�a<��a<ɖa<�a<��a<5�a<�a<ӣa<}�a<T�a<ٚa<v�a<��a<ϒa<Αa<K�a<�a<v�a<ҙa<t�a<��a<ڣa<��a<إa<e�a<��a<H�a<�a<+�a<��a<�wa<jna<=fa<�_a<�[a<Za<D[a<�^a<ea<�la<va<�a<G�a<�a<v�a<��a<��a<J�a<.�a<h�a<��a<�a<1�a<��a<�a<�a<W�a<�a<��a<]�a<��a<�a<,�a<��a<��a<�a<��a<=�a<�a<��a<��a<�xa<�na<�ea<�]a<�Wa<�Ta<�Sa<�Ua<�Ya<o`a<�ha<�qa<'{a<.�a<U�a<��a<U�a<�a<��a<n�a<��a<#�a<��a<��a<چa<��a<Ӂa<	�a<��a<�a<d�a<:�a<�a<X�a<юa<ώa<,�a<�a<Ճa<||a<Vsa<Fia<�^a<vTa<@Ka<�Ca<�=a<�:a<�:a<�<a<�Aa<�Ha<�Pa<)Za<[ca<la<�sa<Yya<k}a<ba<�a<�}a<#{a<�wa<�sa<�oa<sla<@ja<�ha<�ha<Hja<}la<�oa<�ra<,va<�xa<hza<_za<�xa<�ta<Toa<�ga<�^a<bUa<yKa<Ba<�9a<w3a<u/a<�-a<A/a<3a<^9a<pAa<�Ja<�Ta<�  �  �ba<uja<%qa<�ua<�xa<�ya<�xa<xva<�ra<�na<�ja<�fa<�ca<`ba<Eba<aca<	fa<�ia<lna<^sa<xa<A|a<
a<h�a<�a<"}a<�xa<mra<ka<�ba<�Za<�Ra<�La<9Ha<�Ea<Fa<�Ha<�Ma<�Ta<]a<|fa<*pa<bya<w�a<.�a<�a<ۏa<��a<ԏa<��a<,�a<��a<��a<�a<~a<_}a<~a<�a<��a<�a<�a<�a<�a<Қa<!�a<�a<��a<j�a<'�a<f�a<y�a<�|a<�ta<�la<�fa<dba<�`a<�`a<�ca<ia<�oa<xa<ڀa<։a<�a<��a<O�a<��a<=�a<��a<��a<$�a<��a<��a<f�a<�a<��a<܉a<@�a<�a<2�a<5�a<Зa<�a</�a<�a<S�a<�a<b�a<�a<��a<5�a<��a<�}a<ua<�ma<�ga<�ca<�ba<�ca<ga<�la<�sa<|a<Ԅa<p�a<�a<S�a<��a<b�a<�a<��a<ܞa<ǚa<]�a<��a<u�a<)�a<�a<k�a<��a<�a<=�a<F�a<��a<��a<2�a<P�a<��a<��a<Q�a<�a<%�a<�a<~a<ua<�la<�ea<`a<�\a</\a<�]a<�aa<�ga<oa<fwa<�a<��a<юa<D�a<��a<P�a<��a<��a<͒a<�a<�a<�a<ya<|a<�ya<ya<�ya<�{a<�~a<9�a<Ѕa<G�a<Ћa<ʌa<c�a<��a<N�a<�~a<�va<�ma<Zda<�Za<fRa<|Ka<Fa<gCa<Ca<Ea<�Ia<�Oa<JWa<{_a<�ga<Yoa<�ua<�za<m}a<k~a<I}a<�za<�va<)ra<Rma<�ha<�da<$ba<�`a<�`a<vba<:ea<�ha<Dma<Lqa<"ua<�wa<�xa<Exa<�ua<qa<�ja<ca<TZa<aQa<�Ha<hAa<�;a<�7a<w6a<�7a<6;a<�@a<(Ha<�Pa<�Ya<�  �  Pga<�ma<Gsa<�va<]xa<�wa<�ua<�qa<Dma<ha<�ba<^a<
[a<Ya<�Xa<Za<@]a<�aa<�fa<�la<�ra<xa<|a<�~a<�a<Y~a<{a<%va<pa<�ha<�aa<*[a<�Ua<�Qa<zOa<�Oa<Ra<�Va<�\a<�da<ma<�ua<�}a<c�a<��a<f�a<��a<e�a<�a<��a<O�a<�a<{a<�wa<�ta<ta<�ta<�va<�za<�a<ƅa<�a<��a<��a<Кa<�a<��a<	�a<�a<��a<Ɋa<H�a< |a<=ua<�oa<�ka<ja<�ja<!ma<�qa<�wa<\a<�a<�a<͕a<}�a<��a<��a<ˡa<�a<{�a<��a<��a</�a<P�a<M�a<r�a<i�a<�a<�a<Ԇa<}�a<�a<x�a<��a<��a<c�a<E�a<3�a<�a<��a<��a<>�a<��a<�|a<2va<�pa<vma<,la<ma<9pa<'ua<�{a<�a<��a<�a<[�a<v�a<��a<�a<�a<`�a<W�a<@�a<��a<�a<%�a<4�a<�~a<�}a<�~a<H�a<�a<ʉa<)�a<e�a<�a<`�a<f�a<o�a<��a<��a<ܒa<�a<�a<Q|a<�ta<Cna<nia<zfa<�ea<8ga<�ja<pa<�va<�}a<a�a<<�a<��a<�a<1�a<V�a<~�a<Ԓa<�a<*�a<�a<|a<�va<�ra<pa<�oa<tpa< sa<�va<�za<�a<S�a<��a<y�a<B�a<�a<�a<��a<{a<Fsa<�ja<�ba<�Za<CTa<�Oa<�La<�La<zNa<LRa<�Wa<�^a<�ea<�la<8sa<Sxa<�{a<j}a<�|a<�za<�va<�qa<�ka<�ea<�`a<)\a<�Xa<{Wa<�Wa<uYa<�\a<9aa<_fa<�ka<pa<Rta<�va<�wa<`va< sa<�ma<�ga<�_a<2Xa<�Pa<�Ia<�Da<9Aa<@a<Aa<VDa<pIa<)Pa<�Wa<�_a<�  �  #la<}qa<lua<zwa<�wa<�ua<:ra<4ma<(ga<�`a<�Za<TUa<NQa<�Na<tNa<Pa<�Sa<�Xa<�^a<�ea<�la<�sa<ya<	}a<"a<Fa<�}a< za<$ua<Xoa<Wia<�ca<�^a<m[a<�Ya<�Ya<:\a<G`a<�ea<�la<�sa<M{a<�a<��a<��a<��a<��a<ߋa<E�a<p�a<�}a<�wa<�ra<na<ka<�ia<bja<ma<nqa<Twa< ~a<e�a<��a<��a<(�a<��a<��a<u�a<��a<ŕa<O�a<%�a<ރa<~a<Bya<�ua<Qta<�ta<wa<{a<��a<�a<��a<!�a<Ǚa<+�a<��a<i�a<#�a<��a<,�a<@�a<��a<F�a<ka<�za<�wa<va<�va<Qya<�}a<-�a<��a<7�a<��a<�a<(�a<\�a<��a<
�a<|�a<o�a<G�a<��a</�a<Wa<�za<�wa<mva<Swa<za<]~a<�a<D�a<ːa<�a<��a<��a<V�a< �a<�a<�a<��a<"�a<T�a<ׁa<�{a<vwa<�ta<�sa<�ta<�wa<|a<ʁa<�a<��a<|�a<O�a<��a<�a<q�a<�a<��a<�a<��a<��a<I}a<�wa<Ssa<�pa<�oa<Zqa<ita<ya<�~a<�a<�a<��a<��a<��a<]�a<�a<��a<��a<��a<��a<_za<�sa<�ma<ia<7fa<aea<�fa<{ia<�ma<Hsa<#ya<�~a<��a<Їa<�a<�a<W�a<��a<Xa<�xa<�qa<Oja<�ca<�]a<�Ya<4Wa<�Va<mXa<�[a<�`a<+fa<8la<&ra<3wa<{a<�|a<$}a<T{a<�wa<Vra<�ka<�da<^a<�Wa<�Ra<�Na<!Ma<vMa<�Oa<�Sa<�Xa<�^a<iea<�ka<�pa<�ta<�va<�va<ua<dqa<>la<fa<S_a<�Xa< Sa<]Na<jKa<DJa<HKa<Na<�Ra<~Xa<�^a<�ea<�  �  �pa<�ta<nwa<&xa<�va<�sa<�na<Pha<�`a<�Ya<YRa<La<~Ga<�Da<6Da<�Ea<�Ia<�Oa<�Va<�^a<ga<�na<�ua<,{a<�~a<C�a<�a<�}a<za<�ua<�pa<la<,ha<;ea<�ca<=da<#fa<�ia<�na<|ta<�za<�a<C�a<x�a<�a<Ǎa<��a<�a<;�a<!~a<wa<apa<�ia<�da<aa<�_a<)`a<ca<�ga<�na<qva<�~a<�a<Ԏa</�a<4�a<�a<�a<��a<ߙa<Еa<�a<��a<ʆa<ςa<�a<�~a<�~a<�a<��a<�a<i�a<�a<D�a<��a<��a<ۡa<'�a<r�a<��a<��a<v�a<��a<T}a<nva<�pa<Uma<�ka<�la<qoa<<ta<�za<'�a<̉a<��a<E�a<��a<��a</�a<�a<��a<��a<3�a<��a<8�a<_�a<d�a<��a<ˀa<h�a<��a<�a<&�a<{�a<ؖa<��a<F�a<��a<�a<g�a<Ŝa<R�a<��a<߈a<�a<rya<�ra<�ma<`ja<Tia<�ja<�ma<sa<�ya<�a<��a<܏a<�a<��a<��a<m�a<P�a<N�a<�a<ܐa<,�a<��a<�a<!}a<�za<Sza<E{a<~a<ځa<��a<͋a<��a<ڔa<՗a<8�a<��a<��a<2�a<�a<m�a<�za<�ra<�ja<da<_a< \a<([a<�\a<�_a<ea<�ka<Tra<xya<�a<քa<��a<$�a<ɉa<p�a<q�a<K~a<Xxa<ra<Fla<bga<�ca<�aa<aa<Eba<%ea< ia<�ma<�ra<Iwa<�za<w}a<$~a<�|a<�ya<Xta<�ma<%fa<�]a<Va<�Na<�Ha<�Da<�Ba<;Ca<�Ea<IJa<nPa<�Wa<�^a<�fa<�la<Ara<�ua<Zwa<�va<�ta<�pa<�ka<mfa<�`a<\a<Xa<pUa<�Ta<ZUa<�Wa<�[a<�`a<-fa<�ka<�  �  Bua<�wa<2ya<�xa<�ua<kqa<ka<�ca<[a<�Ra<KJa<�Ca<Q>a<);a<�:a<j<a<�@a<'Ga<Oa<Xa<laa<|ja<yra<5ya<�}a<�a<߁a<�a<�~a<]{a<�wa<�sa<�pa<Dna<;ma<�ma<^oa<�ra<�va<�{a<�a<�a<M�a<�a<{�a<��a<�a<�a<J�a<ya<�pa<�ha<�aa<�[a<�Wa<�Ua<�Va<�Ya<&_a<5fa<�na<Mxa<�a<��a<x�a<��a<Ϝa<�a<'�a<ŝa<Қa<��a<�a<ʎa<j�a<
�a<�a<S�a<�a<��a<�a<��a<ޙa<�a<.�a<��a<¢a<��a<��a<��a<^�a<�a<~a<�ua<na<ha<�ca<@ba<�ba<)fa<�ka<�ra<�za<ڃa<��a<��a<e�a<]�a<r�a<��a<��a<I�a<��a<H�a<��a<��a<=�a<��a<E�a<��a<��a<a<��a<*�a<O�a<�a<w�a<b�a<k�a<h�a<��a<Փa<��a<�a<za<bqa<-ja<uda<�`a<�_a<�`a<�da<�ja<�qa<@za<��a<d�a<��a<Ęa<ۜa<*�a<O�a<͝a<ƚa<��a<!�a<j�a<Q�a<+�a<=�a<��a<��a<��a<�a<�a<��a<֕a<�a<u�a<��a<��a<��a<��a<�a<N~a<�ta<cka<�ba<d[a<�Ua<lRa<�Qa<Sa<2Wa<�\a<da<
la<;ta<�{a<�a<�a<�a<��a<ىa<U�a<L�a<d~a<[ya<Eta<�oa<�la<�ja<jja<\ka<�ma<�pa<�ta<�xa<|a<�~a<�a<a<N|a<�wa<Wqa<�ia<�`a<VWa<TNa<VFa<�?a<K;a<X9a<�9a<�<a<�Aa<NHa<vPa<Ya<�aa<\ia<�oa<�ta<�wa<�xa<�wa<ua<Cqa<�la<dha<1da<�`a<�^a<^a<�^a<�`a<da<7ha<�la<>qa<�  �  �xa<rza<|za<�xa<ua<�oa< ha<a_a<�Ua<qLa<�Ca<�;a<%6a<�2a<.2a</4a<�8a<�?a<]Ha<4Ra<�\a<�fa<�oa<�wa<o}a<��a<y�a<ԃa<��a<N�a<j}a<vza<�wa<va<Aua<�ua<xwa<za<�}a<�a<^�a<S�a<u�a<K�a<c�a<��a<ȉa<D�a<�|a<tta<�ka<�ba<�Za<Ta<�Oa<�Ma<)Na<eQa<8Wa<_a<qha<�ra<=}a<0�a<%�a<?�a<��a<�a<=�a<Ԡa<��a<6�a<��a<��a<�a<�a<�a<R�a<�a<P�a<��a<P�a<�a<�a<�a<}�a<h�a<&�a<��a<�a<��a<"�a<cxa<�na<�fa<`a<�[a<�Ya<�Za<�]a<�ca<�ka<�ta<�~a<j�a<��a<f�a<\�a<��a<��a<
�a<��a<�a<��a<%�a<��a<�a<�a<0�a<˒a<i�a<��a<;�a<��a<��a<��a<�a<��a<��a<��a<��a<�a<��a<�}a<�sa<�ja<�ba<F\a<�Xa<GWa<�Xa<�\a<ca<+ka<cta<~a<i�a<�a<�a<K�a<��a<�a<��a<��a<}�a<їa<�a<��a<�a<D�a<��a<��a<?�a<�a<�a<N�a<�a<�a<��a<~�a<p�a<A�a<`�a<��a<�ya<boa<ea<�[a<�Sa<|Ma<Ja<(Ia<�Ja<DOa<�Ua<�]a<�fa<�oa<+xa<�a<��a<��a<Ћa<�a<d�a<o�a<��a<ma<2{a<vwa<�ta<�ra<ira<Gsa<�ta<�wa<�za<�}a<�a<r�a<W�a<�a<�{a<2va<�na<�ea<�[a<�Qa<�Ga< ?a<�7a<3a<�0a<X1a<a4a<�9a<Aa<LJa<�Sa<^]a<Hfa<�ma<�sa<�wa<�ya<�ya<uxa<�ua<`ra<�na<Uka<�ha<�fa< fa<�fa<|ha<6ka<�na<]ra<�ua<�  �  c{a<g|a<�{a<ya<ata<�ma<�ea<\a<�Qa<�Ga<T>a<*6a<0a<�,a<�+a<.a<�2a<:a<FCa<�Ma<�Xa<fca<nma<va<�|a<�a<΄a<�a<i�a< �a<��a<�a<_}a<�{a<P{a<�{a<J}a<�a<�a<��a<v�a<��a<�a<�a<�a<��a<׈a<C�a<"za<�pa<4ga<�]a<EUa<Na<}Ia<(Ga<�Ga<YKa<'Qa<�Ya<�ca<fna<�ya<Y�a<�a<.�a<��a<��a<�a<0�a<3�a<@�a<n�a<��a<|�a<ٖa<�a<l�a<��a<�a<ʜa<��a<Ӣa<�a<1�a<�a<ͣa<ԟa<��a<ˑa<{�a<Y~a<�sa<�ia< aa<�Ya<wUa<CSa<ITa<�Wa<^a<wfa<pa<�za<	�a<�a<��a<��a<ţa<��a<�a<:�a<��a<�a<�a<�a<��a<�a<B�a<Șa<�a<_�a< �a<�a<��a<0�a<�a<ɥa<�a<�a<��a<Z�a<v�a<�ya<2oa<iea<�\a<<Va<?Ra<�Pa<�Ra<�Va<}]a<fa<�oa<3za<J�a<��a<��a<ڛa<	�a<<�a<��a<\�a<O�a<�a<&�a<"�a<��a<T�a<Ƒa<m�a<֓a<6�a<��a<f�a<u�a<|�a<k�a</�a<n�a<Q�a<`�a<ڀa<8va<ka<`a<6Va<�Ma<vGa<�Ca<�Ba<�Da<4Ia<EPa<�Xa<"ba<�ka<Sua<�}a<��a<��a<_�a<��a<��a<��a<��a<ۃa<o�a<}a<�za<�xa<�xa<�xa<�za<�|a<�~a<v�a<�a<��a<˂a<�a<�{a<�ta<~la<�ba<Xa<Ma<�Ba<s9a<�1a<�,a<^*a<+a<[.a<4a<9<a<zEa<�Oa<�Ya<�ca<la<�ra<�wa<�za<�{a<{a<\ya<�va<�sa<�pa<-na<�la<la<�la<na<�pa<�sa<�va<�ya<�  �  #}a<�}a<3|a<ya<�sa<�la<da<7Za<tOa<�Da<�:a<~2a<4,a<c(a<�'a<�)a<�.a<j6a<�?a<�Ja<>Va<�aa<la<@ua<�|a<�a<~�a<'�a<?�a<?�a<��a<��a<݀a<�a<=a<�a<�a<^�a<S�a<��a<ڌa<��a<i�a<ܑa<��a<b�a<<�a<!�a<�xa<�na<�da<�Za<�Qa<dJa<XEa<�Ba<�Ca<&Ga<xMa<Va<``a<�ka<owa<��a<Ռa<��a<:�a<�a<��a<��a<"�a<��a<j�a<(�a<�a<��a<#�a<c�a<v�a<l�a<�a<��a< �a<Ǧa<~�a<��a<�a<k�a<�a<t�a<ʆa<�{a<qa<�fa<q]a<&Va<;Qa</Oa<Pa<�Sa<bZa<�ba<ma<xa<�a<e�a<��a<�a<��a<>�a<�a<�a<��a<��a<��a<n�a<C�a<ݜa<X�a<��a<ѝa<ȟa<1�a<��a<��a<�a<�a<e�a<�a<c�a<�a<یa<��a<iwa<Ola<�aa<Ya<SRa<Na<�La<RNa<�Ra<�Ya<�ba<�la<�wa<��a<=�a<˔a<j�a<+�a<�a<٣a<2�a<n�a<��a<;�a<��a<��a<@�a<וa<9�a<��a<q�a<��a<ʝa<k�a<�a<<�a<��a<2�a<��a<>�a<Ba<ta<sha<]a<�Ra<�Ia<QCa<u?a<�>a<�@a<�Ea<�La<�Ua<u_a<�ia<�sa<z|a<�a<Q�a<Ìa<]�a</�a<��a<��a<׆a<��a<��a<_~a<}a<y|a<�|a<~a<�a<ҁa<��a<̈́a<�a<��a<N�a<+{a<%ta<'ka<�`a<�Ua<NJa<k?a<�5a<.a<�(a<K&a<�&a<_*a<s0a<�8a<�Ba<5Ma<Xa< ba<ka<fra<�wa<A{a<�|a<�|a<\{a<(ya<�va<ta<�qa<�pa<%pa<�pa<�qa<ta<�va<Eya<�{a<�  �  ��a<��a<ςa<S~a<;wa<�ma<�aa<�Sa<8Ea<�6a<,)a<�a<�a<�a<4a<Sa<+a<H"a</a<�=a<�La<F\a<Oja<�va<m�a<��a<N�a<}�a<�a<x�a<`�a<��a<��a<߄a<�a<��a<4�a<�a<8�a</�a<�a<;�a<A�a<2�a<B�a<s�a<4�a<?�a<Eua<�ga<�Ya<La<w?a<G5a<0.a<�*a<+a<�/a<B8a<�Ca<�Qa<�`a<:pa<ma<�a<��a<��a<�a<��a<�a<o�a<��a<Ƨa<Ϥa<��a<��a<��a<ߟa<[�a<ãa<��a<�a<֬a<�a<{�a<!�a<��a<�a<F�a<��a<s�a<�sa<ea<�Va<GJa<V@a<�9a<}6a<�7a<.=a<�Ea<�Qa<g_a<na<�|a<�a<��a<ԡa<p�a<w�a<��a<%�a<��a<�a<ĩa<��a<J�a<Z�a<��a<�a<��a<�a<ܨa<�a<��a<%�a<ʯa<��a<רa<c�a<b�a<�a<�|a<�ma<_a<�Pa<�Da<�;a<�5a<�3a<v6a<�<a<BFa<iRa<�`a< oa<�}a<�a<Ŗa<ҟa<p�a<H�a<��a<d�a<6�a<W�a<բa<�a<\�a<��a<N�a<�a<ʝa<�a<͢a<��a<��a<]�a<�a<ңa<��a<�a<��a<I|a<8ma<�]a<�Na<�@a<�4a<',a<�&a<�%a<E)a<0a<:a<^Fa<Ta<'ba<�oa<4|a<��a<�a<P�a<��a<�a<9�a<?�a<�a<��a<`�a<��a<́a<@�a<��a<��a<υa<��a<Ҋa<g�a<H�a<\�a<=�a<?a<�ua<�ia<\a<�La<�=a<�.a<�!a<�a<qa<�a<�a<�a<Qa<�&a<54a<�Ba<GQa<,_a<yka<wua<�|a<Ła<ڃa<5�a<��a<�a<�|a<�ya<2wa<Rua<�ta<<ua<wa<�ya<�|a<�a<Âa<�  �  ȃa<E�a<��a<H~a<twa<na<hba<�Ta<�Fa<$8a<�*a<=a<�a<�a<ga<Ga<�a<�#a<t0a<	?a<3Na<E]a<ka<wa<��a<��a<�a<�a<�a<l�a< �a<a�a<�a<)�a<k�a<��a<z�a<L�a<�a<��a<��a<=�a<��a<�a<�a<��a<x�a<�a<2va<�ha<�Za<EMa<Aa<�6a<�/a<�,a<:-a<�1a<�9a<DEa<�Ra<ba<oqa<_�a<��a<�a<��a<�a<X�a<]�a<r�a<o�a<��a<~�a<Ša<Ϟa<�a<9�a<��a<�a<=�a<��a<ƫa<�a<��a<��a<{�a<M�a<��a<w�a<i�a<�ta<Xfa<*Xa<�Ka<�Aa<{;a<�8a<�9a<�>a<{Ga<Sa<�`a<\oa<!~a<�a</�a<�a<k�a<<�a<d�a<O�a<��a<�a<��a<M�a<��a<��a<�a<d�a<	�a<��a<��a<�a<��a<D�a<s�a<l�a<˨a<��a<ߗa<ϋa<�}a<!oa<I`a<^Ra<uFa<J=a<�7a<6a<j8a<E>a<�Ga<�Sa<�aa<Lpa<�~a<݋a<+�a<
�a<c�a<�a<G�a<k�a<+�a<�a<��a<F�a<��a<�a<��a<4�a<�a<��a<��a<u�a<��a<��a<ͦa<��a<��a<S�a<T�a<5}a<mna<_a<�Oa<Ba<[6a<�-a<)a<(a<+a<�1a<�;a<�Ga<dUa<\ca<�pa<�|a<Նa<;�a<(�a<g�a<C�a<<�a<*�a<F�a<@�a<��a<ʁa<�a<�a<D�a<��a<�a<I�a<a<f�a<ɋa<3�a<(�a<oa<=va<�ja<�\a<Na<�>a<O0a<�#a<"a<Ua<a<�a<�a<�a<((a<u5a<�Ca<iRa<`a<la<�ua<�|a<��a<��a<_�a<��a<�~a<m{a</xa<yua<�sa<sa<�sa<`ua<xa<^{a<�~a<��a<�  �  ��a<܂a<��a<V~a<?xa<uoa<tda<�Wa<�Ia<$<a<M/a<J$a<�a<a<�a<�a<�a<�(a<�4a<�Ba<�Qa<�_a< ma<Exa<E�a<�a<!�a<��a<��a<��a<d�a<<�a<P�a<F~a<h}a<�}a<�a<k�a<��a<��a<��a<��a<��a<��a<��a<�a<q�a<��a<rxa<�ka<�^a<{Qa<�Ea<�;a<H5a<2a<�2a<7a<�>a<Ja<'Wa<�ea<�ta<��a<q�a<�a<.�a<k�a<+�a<��a<��a<0�a<��a<3�a<��a<�a<ژa<.�a<��a<j�a<�a<ߤa<Ĩa<��a<a�a<�a<(�a<ڤa<��a<O�a<څa<?xa<4ja<�\a<�Pa<!Ga<�@a<�=a<L?a<(Da<�La<�Wa<�da<�ra<Հa<�a<��a<�a<��a<u�a<�a<<�a<�a<`�a<z�a<Ԡa<��a<��a<њa<l�a<�a<	�a<��a<J�a<ͪa<!�a<	�a<��a<ڨa<g�a<>�a<ڍa<��a<�ra<Ida<�Va<�Ka<�Ba<K=a<f;a<�=a<�Ca<�La<SXa<�ea<�sa<2�a<Ǎa<]�a<��a<1�a<�a<éa<&�a<M�a<\�a<g�a<��a<a<�a<k�a<G�a<&�a<B�a<��a<#�a<�a<��a<��a<�a<!�a<L�a<��a<ua<^qa<�ba<
Ta<�Fa<~;a<?3a<m.a<q-a<o0a<�6a<k@a<�Ka<"Ya<mfa<;sa<�~a<ևa<��a<��a<:�a<g�a<��a<�a<R�a<��a<�a<�|a<{a<�za<d{a<X}a<P�a<{�a<��a<�a<-�a<#�a<ԅa<�a<Zwa<dla<m_a<TQa<�Ba<�4a<}(a<ca<�a<qa<aa<�a<�!a<�,a<�9a<iGa<Ua<+ba<uma<�va<}a<Āa<<�a<L�a<�~a<L{a<]wa<�sa<�pa<�na<�ma<�na<tpa<�sa<Hwa<D{a<
a<�  �  ~a<Q�a<p�a<9~a<6ya<�qa<�ga<\a<MOa<�Ba<X6a<,a<K$a<�a<�a<9!a<J'a<V0a<�;a<Ia<�Va<�ca<
pa<Bza<��a<&�a<��a<��a<هa<��a<��a<�|a<ya<iva<)ua<sua<~wa<�za<�a<ӄa<R�a<p�a<i�a<��a<��a<�a<܍a<�a<|a<pa<Bda<6Xa<�La<Da<�=a<�:a<R;a<�?a<Ga<ZQa<�]a<{ka<Hya<v�a<�a<��a<|�a<��a<�a<y�a<פa<�a<��a<H�a<��a<ݑa<��a<�a<ђa<�a<R�a<��a<��a<ǧa<��a<&�a<��a<o�a<��a<;�a<�a<@}a<8pa<�ca<8Xa<^Oa<mIa<�Fa<�Ga<�La<bTa<�^a<;ka<Lxa<V�a<��a<�a<�a<��a<L�a<��a<Ϊa<V�a<ܢa<%�a<��a<��a<��a<��a<7�a<f�a<ߘa<�a<��a<�a<��a<}�a<J�a<��a<^�a<q�a<"�a<�a<�wa<�ja<^a<<Sa<	Ka<�Ea<5Da<`Fa<�Ka<TTa<Q_a<�ka<�xa<_�a<Ӑa<\�a<c�a<٥a<��a<��a<[�a<U�a<��a<Ėa<c�a<�a<Ìa<"�a<8�a<��a<D�a<o�a<ϛa<��a<��a<h�a<-�a<S�a<��a<��a<�a<va<Qha<�Za<Na<�Ca<�;a<+7a<46a<�8a<�>a<�Ga<�Ra<�^a<6ka<�va<=�a<g�a< �a<�a</�a<a�a<��a<��a<F�a<}a<axa<�ta<�ra<Kra<usa<va<�ya<�}a<��a<(�a<M�a<`�a<_�a<��a<8ya<Ooa<wca<TVa<�Ha<�;a<�/a<�&a<D a<;a<	a<["a<�)a<�3a<@a<�La<�Ya<�ea<�oa<�wa<}a<�a<�a<�}a<Rza<�ua<qa<�la<�ha<�fa<�ea<jfa<�ha<hla<�pa<�ua<Xza<�  �  xya<}a<�~a<�}a<cza<]ta<�ka<�aa<Va<�Ja<�?a<36a</a<�*a<�)a<-,a<�1a<U:a<�Da<�Pa<*]a<;ia<�sa<�|a<ła<��a<��a<$�a<�a</~a< ya<�sa<Woa<la<�ja<�ja<�la<�pa<Hva<�|a<^�a<ǉa<@�a<֒a<w�a<:�a<��a<3�a<��a<�va<vka<�`a<�Va<|Na<�Ha<�Ea<�Fa<pJa<�Qa<[a<�fa<�ra<�a<:�a<a�a<�a<âa<��a<��a<s�a<V�a<�a<��a<�a<��a<K�a<�a<I�a<`�a<J�a<[�a<D�a<*�a<��a<¦a<�a<�a<�a<ߠa<Иa<�a<��a<�wa<zla<ba<�Ya<[Ta<3Ra<Sa<`Wa<�^a<2ha<xsa<;a<&�a<a<Ξa<j�a<e�a<ժa<��a<S�a<]�a<��a<��a<:�a<؋a<݈a<߇a<��a<.�a<J�a<��a<Z�a<��a<�a<=�a<��a<n�a<��a<'�a<0�a<��a<�~a<�ra<Tga<q]a<�Ua<�Pa<�Oa<WQa<�Va<V^a<`ha<�sa<Ja<��a<��a<��a</�a<Q�a<��a<f�a<o�a<�a<��a<�a<��a<��a<�a<��a<��a<��a<��a<K�a<ٔa<�a<Z�a<��a<�a<r�a<k�a<��a<��a<)|a<�oa<Kca<�Wa<�Ma<�Fa<`Ba<Aa<�Ca<rIa<WQa<o[a<2fa<qqa<�{a<��a<P�a<I�a<�a<��a<[�a<#�a<܀a<Iza<�sa<una<Ija<ha<�ga<ia<:la<�pa<�ua<&{a<�a<��a<>�a<��a</�a<u{a<�ra<�ha<�\a<mPa<�Da<�9a<:1a<0+a<�(a<)a<-a<4a<H=a<DHa<�Sa<m_a<�ia<�ra<ya<�|a<&~a<�|a<gya<\ta<�na<�ha<"ca<�^a<�[a<�Za<�[a<�^a<�ba<Gha<Xna<7ta<�  �  �sa<ya<z|a<r}a<�{a<Pwa<wpa<�ga<^a<�Sa<.Ja<�Aa<~;a<�7a<�6a<9a<7>a<�Ea<9Oa<�Ya<�da<(oa<xa<4a<��a<��a<�a<Ła<�|a<�va<�oa<�ia<�ca<�_a<�]a<^a<�`a<2ea<�ka<sa<+{a<�a<�a<o�a<��a<e�a<_�a<a<ޅa<r}a<�sa<pja<�aa<\Za<QUa<�Ra<�Sa<5Wa<�]a<%fa<kpa<k{a<��a<��a<$�a<z�a<'�a<�a<a�a<v�a<˘a<�a<�a<{�a<�~a<	{a<0ya<�ya<3|a<׀a<��a<�a<��a<{�a<0�a</�a<ߧa<ۦa<<�a<��a<Ȕa<�a<��a<�va<wma<.fa<9aa<1_a<
`a<�ca<eja<�ra<�|a<_�a<��a<��a<�a<ݦa<%�a<��a<��a<Ƞa<R�a<�a<ŋa<:�a<�a<d|a< {a<�{a<)a<)�a<z�a<��a<Řa<5�a<:�a<R�a<��a<֥a<�a<��a<�a<��a<|a<�qa<
ia<Bba<�]a<�\a<>^a<�ba<�ia<�ra<�|a<�a<��a<�a<S�a<$�a<b�a<�a<�a<i�a<m�a<�a<��a<Q}a<exa<lua<�ta<Hva<�ya<Aa<��a<��a<^�a<-�a<F�a<@�a<��a<6�a<2�a<ߌa<��a<�wa<�la<�ba<�Ya<GSa<aOa<�Na<�Pa<iUa<w\a<@ea<�na<uxa<�a<K�a<L�a<��a<]�a<s�a<`�a<��a<�xa<�pa<Bia<�ba<^a<][a<�Za<�\a<�`a<;fa<�la<{sa<�ya<�~a<f�a<��a<��a<�}a<wa<Una<+da<NYa<�Na< Ea<i=a<8a<�5a<6a<�9a<�?a<Ha<�Qa<�[a<�ea<�na<�ua<�za<�|a<|a<�xa<�sa<Tma<fa<�^a<%Xa<�Ra<fOa<9Na<7Oa<�Ra<�Wa<=^a<�ea<ma<�  �  uma<�ta<�ya<�|a<�|a<@za<]ua<jna<afa<�]a<aUa<Na<�Ha<wEa<�Da<�Fa<0Ka<�Qa<%Za<bca<�la<Gua<�|a<��a<f�a<_�a<�a<�|a<$va<Tna<fa<2^a<rWa<�Ra<TPa<qPa<?Sa<PXa<�_a<|ha<!ra<�{a<b�a<��a<��a<@�a<�a<b�a<M�a<��a<�|a<�ta<3ma<�fa<�ba<�`a<raa<�da<7ja<�qa<�za<��a<̍a<5�a<��a<G�a<6�a<0�a<Ξa<��a<��a<<�a<��a<�xa<#ra<�ma<�ka<�ka<oa<1ta<�{a<��a<��a<��a<(�a< �a<b�a<Y�a<x�a<I�a<��a<Ȓa<!�a<^�a<}ya<sa<�na<ma<�ma<;qa<�va<I~a<��a<ۏa<J�a<��a<�a<�a<��a<=�a<��a<��a<�a<��a<�a<ya<�ra<oa<pma<�na<$ra<�wa<ua<�a<ʐa<�a<�a<��a<�a<�a<�a<Ǟa<n�a<��a<�a<}a<Qua<roa<�ka<�ja<la<�oa<�ua<�}a<-�a<ˎa<Ėa<k�a<͡a<գa<�a<�a<<�a<��a<�a<��a<\xa<�pa<Lka<�ga<ga<�ha<ma<bsa<{a<��a<�a<y�a<��a<*�a<u�a<לa<Ҙa<M�a<�a<ڀa<>wa<;na<`fa<�`a<6]a<U\a<^a<ba<>ha<�oa<�wa<�a<��a<"�a<�a<��a<x�a<�a<�a<Vya<�oa<\fa<�]a<Va<�Pa<�Ma<cMa<�Oa<"Ta<�Za<�ba<�ja<�ra<�ya<6a<�a<s�a<
�a<U{a<Ita<�ka<�ba<wYa<#Qa<EJa<�Ea<wCa<�Ca<�Fa<La<[Sa<�[a<ada<�la<�sa<�xa<�{a<|a<�ya<�ta<�ma<�ea<�\a<�Sa<La<�Ea<	Ba<�@a<�Aa<�Ea<rKa<;Sa<\a<ea<�  �  ga<�oa<
wa<�{a<�}a<�|a<�ya<�ta<ona<bga<v`a<dZa<�Ua<�Ra<qRa<(Ta<"Xa<�]a<�da<�la<_ta<H{a<��a<�a<�a<�a<�~a<�wa<^oa<�ea<�[a<�Ra<Ka<Ea<�Ba<�Ba<�Ea<�Ka<�Sa<�]a<�ha<ta<�~a<��a<��a<ݒa<��a<��a<q�a<��a<j�a<�~a<�xa<�sa<�oa<Yna<oa<�qa<wa<�}a<*�a<J�a<��a<��a<r�a<�a<�a<I�a<ښa<C�a<'�a<�a<va<�la<pea<,`a<�]a<)^a<�aa<�ga<�oa<�ya<3�a<��a<їa<�a<ڤa<��a<��a<#�a<��a<V�a<D�a<�a<n�a<�a<A|a<�za<[{a<Q~a<7�a<��a<��a<�a<�a<`�a<�a<A�a<��a<��a<��a<v�a<~�a<�a<�ua<�la<�ea<;aa<�_a<�`a< ea<�ka<Qta<A~a<��a<��a<�a<�a<(�a<ԧa<��a<>�a<؝a<�a<��a<3�a<��a<~|a<0ya<2xa<]ya<�|a<��a<\�a<}�a<��a<Ȝa<x�a<+�a<W�a<ʡa<��a<�a<�a<��a<�va<�la<gda<�]a<Za<CYa<M[a<8`a<kga<_pa<Hza<Y�a<��a<X�a<�a<�a<p�a<�a<p�a<�a<w�a<^�a<�ya<sa<�ma<�ja<�ia<Wka<�na<�sa<za<��a<�a<�a<��a<�a<��a<��a<�a<0|a<�qa<�fa<�[a<�Qa<OIa<-Ca<�?a<�?a<IBa<�Ga<6Oa<gXa<-ba<�ka<�ta<�{a<��a<��a<8�a<-a<za<^sa<�ka<da<]a<+Wa<Sa< Qa<fQa<Ta<�Xa<�^a<xea<�la<7sa<mxa<�{a<�|a<:{a<�va<0pa<�ga<�]a<Sa<�Ha<�?a<�8a<D4a<�2a<4a<f8a<6?a<Ha<ERa<�\a<�  �  �`a<Nka<.ta<qza<B~a<Wa<�}a<�za<�ua<6pa<�ja<�ea<�aa<}_a<-_a<�`a<da<�ha<�na<,ua<S{a<��a<Y�a<�a<	�a<��a<^{a<�ra<�ha<�]a<~Ra<�Ga<R?a<�8a<�5a<�5a<�8a<a?a<wHa<�Sa<`a<�la<�xa<r�a<A�a<*�a<ߕa<��a<!�a<ˑa<)�a<'�a<)�a<a<#|a<{a<�{a<8~a<��a<�a<��a<2�a<i�a<u�a<��a<��a<��a<3�a<��a<ˍa<
�a<bwa<2la<�aa<hYa<`Sa<�Pa<'Qa<�Ta<�[a<�da<*pa<�{a<؇a<��a<�a<(�a<��a<��a<��a<եa<%�a<��a<��a<9�a<��a<��a<v�a<�a<q�a<��a<��a<��a<��a<�a<��a<��a<�a<��a<��a<��a<p�a<ɂa<�va<�ka<raa<�Ya<PTa<�Ra<�Sa<�Xa<`a<�ia<ua<��a<Q�a<t�a<�a<�a<k�a<"�a<V�a<��a<P�a<g�a<L�a<܌a<��a<Ʌa<�a<΅a<��a<�a<:�a<��a<��a<<�a</�a<8�a<|�a<C�a<b�a<#�a<V�a<Lya<wma<ba<�Xa<ZQa<Ma<FLa<wNa<Ta<!\a<Yfa<vqa<
}a<��a<E�a<ɘa<]�a<��a<�a<�a<T�a<5�a<��a<0�a<�~a<za<�wa<�va<�wa<jza<s~a<y�a<��a<Z�a<��a<��a<b�a<�a<~�a<�a<�va<�ja<&^a<�Qa<�Fa<I=a<b6a<�2a<�2a<�5a<�;a<?Da<�Na<�Ya<6ea<oa<@xa<�~a<��a<�a<��a<Za<+za<ta<�ma<�ga<�ba<j_a<�]a<^a< `a<�ca<�ha<xna<ta<+ya<�|a<i~a<�}a<2za<Rta<�ka<�aa<�Ua<�Ia<�>a<g4a<�,a<\'a<�%a<'a<�+a<�3a<�=a<Ia<�Ta<�  �  M[a<Yga<�qa<]ya<�~a<�a<B�a<Va<�{a<�wa</sa<.oa<�ka<#ja<�ia<<ka<na<Dra<$wa<O|a<5�a<�a<S�a<r�a< �a<�a<lxa<�na<�ba<�Va</Ja<�>a<�4a<".a<h*a<:*a<�-a<�4a<�>a<�Ja<wXa<_fa<�sa<�a<�a<��a<��a<Әa<�a<�a<ēa<��a<-�a<�a<��a<��a<i�a<Èa<x�a<?�a<��a<�a<Ӡa<i�a<��a<y�a<(�a<3�a<��a<�a<�|a<�oa<vca<�Wa<�Na<�Ha<bEa<�Ea<%Ja<vQa<|[a<�ga<�ta<́a<9�a<��a<��a<��a<��a<v�a<�a<�a<��a<��a<��a<ʕa<A�a<�a<��a<Ŕa<4�a<��a<:�a<�a<��a<+�a<{�a<��a<ҥa<��a<��a<�a<-|a<oa<rba<cWa<�Na<TIa<Ga<�Ha<�Ma<�Ua<�`a<ma<�ya<��a<}�a<c�a<ޣa<ʨa<�a<��a<^�a<��a<ʟa<�a<y�a<͒a<r�a<��a<x�a<Òa<V�a<��a<$�a<d�a<��a<,�a<��a<��a<Ξa<q�a<ҋa<ra<Kra<(ea<�Xa<NNa<�Fa<�Aa<�@a<�Ca<~Ia<GRa<}]a<�ia<�va<�a<Ía<��a<Ԝa<x�a<?�a<�a<��a<Зa<{�a<4�a<e�a<��a<#�a<L�a<�a<N�a<��a<b�a<R�a<Œa<�a<&�a<O�a<��a<�a<�}a<�qa<�da<�Va<8Ia<�<a<�2a<�+a<�'a<c'a<�*a<g1a<�:a<RFa<�Ra<*_a<�ja<,ua<+}a<��a<M�a<|�a<��a<�a<#{a<va</qa<�la<ja<xha<�ha<rja<�ma<�qa< va<eza<~a<7�a<S�a<8~a<Qya<�qa<�ga<&\a<9Oa<Ba<j5a<[*a<�!a<ca<Da<a<A!a<�)a<f4a<Aa<;Na<�  �  �Va<!da<koa<xxa<�~a<p�a<܃a<�a<��a<?}a<�ya<^va<�sa<Yra<ra<^sa<�ua<Yya<g}a<Áa<��a<v�a<��a<��a<�a<�~a<va<ka<`^a<Qa<�Ca<w7a<-a<�%a<�!a<q!a<W%a<�,a<@7a<Da<�Ra<jaa<�oa<}a<I�a<�a<)�a<��a<ۛa<��a<��a<ەa<��a<A�a<��a< �a<��a<ɐa<�a<�a<��a<$�a<ߤa<b�a<�a<"�a<ȡa<��a<�a<�a<�wa<-ja<�\a<�Pa<�Fa<�?a<�<a<C=a<�Aa<{Ia<YTa<aa<"oa<,}a<��a<}�a<2�a<`�a<��a<��a<H�a<@�a<��a<&�a<��a<S�a<V�a<a�a<�a<��a<t�a<�a<��a<˪a<{�a<�a<��a<תa<�a<w�a<��a<Ʉa<wa<�ha<p[a<�Oa<�Fa<�@a<M>a</@a<jEa<ANa<�Ya<�fa<�ta<`�a<E�a<?�a<��a<��a<<�a<H�a<��a<L�a<s�a<p�a<��a<��a<��a<�a<��a<]�a<m�a<ߠa<��a<�a<��a<��a<��a<��a<��a<�a<Y�a<�za<�la<�^a<�Qa<qFa<>a<P9a<8a<;a<JAa<�Ja<�Va<�ca<�qa<�~a<�a<ϔa<P�a<��a<�a<آa<}�a<�a<f�a<��a<��a<��a<l�a<��a<$�a<��a<t�a<b�a<��a<іa<�a<�a<��a<T�a<؅a<�za<na<�_a<�Pa<fBa<~5a<�*a<#a<�a<�a<N"a<m)a<�3a<�?a<Ma<�Za<jga<�ra<�{a<t�a<C�a<��a<Ɇa<B�a<�a<4|a<6xa<�ta<ra<�pa<�pa<Cra<�ta<'xa<�{a<Ma<��a<�a<ׁa<�~a<�xa<�oa<�da<�Wa<Ja<�;a<i.a<�"a<�a<�a<ua<wa<�a<�!a<`-a<�:a<�Ha<�  �  `Ta<ba<na<�wa<�~a<U�a<M�a<�a<e�a<�a<�}a<�za<�xa<Pwa<9wa<Rxa<�za<�}a<s�a<8�a<Q�a<��a<��a<B�a<݄a<�}a<�ta<�ha<�[a<�Ma<�?a<�2a<(a<P a<Ta<a<�a<['a<V2a<�?a<�Na<3^a<rma<I{a<4�a<��a<��a<Ûa<��a<Z�a<��a<��a<.�a<�a<v�a<�a<ȓa<��a<��a<d�a<w�a<V�a<S�a<0�a<�a<��a<M�a<��a<%�a<��a<�ta<gfa<LXa<�Ka<�Aa<�:a<G7a<�7a<N<a<ZDa<�Oa<�\a<ka<Jza<p�a<�a<>�a<
�a<T�a<��a<E�a<ͭa<X�a<,�a<��a<<�a<G�a<��a<�a<�a<�a<=�a<��a<��a<��a<_�a<�a<��a<_�a<:�a<��a<G�a<�sa<�da<�Va<�Ja<8Aa<Y;a<9a<�:a<@a<7Ia<�Ta<�ba<Cqa<�a<@�a<�a<7�a<��a<"�a<��a<&�a<�a<�a<��a<8�a<x�a<��a<�a<��a<M�a<ߡa<�a<�a<��a<	�a<۫a<m�a<U�a<��a<��a<9�a<'xa<Eia<}Za<�La<XAa<�8a<�3a<�2a<�5a<<a<�Ea<-Ra<$`a<{na<�|a<�a<��a<˛a<Z�a<.�a<��a<�a< �a<>�a<4�a<n�a<k�a<x�a<��a<�a<y�a<��a<O�a<��a<E�a<��a<G�a<i�a<ٍa<҄a<>ya<�ka<�\a<-Ma<>a<�0a<g%a<�a<xa<Ja<�a<L$a<�.a<t;a<xIa<�Wa<5ea<qa<�za<�a<ކa<��a<ƈa<Άa<݃a<9�a<�|a<iya<wa<�ua<�ua<*wa<fya<I|a<ta<�a<��a<l�a<ʂa<�~a<�wa<�na<�ba<iUa<�Fa<�7a<�)a<�a<<a<la<+a<a<�a<�a<�(a<�6a<�Ea<�  �  QSa<Eaa<�ma<~wa<�~a<��a<��a<�a<m�a<�a<a<a|a<]za<�xa<�xa<za<\|a<a<��a<c�a<O�a<O�a<E�a<{�a<ބa<�}a<�sa<ha<uZa<)La<D>a<01a<p&a<�a<?a<�a<a<�%a<�0a<?>a<qMa<�\a<|la<�za<��a<q�a<��a<�a<�a<Z�a<�a<�a<~�a<��a<2�a<��a<t�a<f�a<c�a<��a<��a<j�a<Q�a<Ωa<N�a<��a<+�a<=�a<v�a<Ɓa<�sa<ea<�Va<AJa<�?a<�8a<%5a<�5a<�:a<�Ba<Na<�[a<(ja<ya<��a<K�a<��a< �a<��a<6�a<�a<ˮa<z�a<c�a<I�a<��a< �a<I�a<��a<6�a<��a<��a<�a<��a<��a<ΰa<(�a<�a<'�a<Ϛa<ݎa<@�a<Wra<�ca<yUa<>Ia<�?a<_9a<�6a<�8a<�>a<�Ga<zSa<saa<�oa<�~a<h�a<s�a<��a<�a<`�a<�a<�a<�a<S�a<Ǧa<��a<0�a<K�a<Ǟa<E�a<
�a<6�a<'�a<;�a<��a<٬a<"�a<��a<V�a<z�a<�a<P�a<�va<�ga<=Ya<YKa<�?a<7a<�1a<�0a<�3a<�:a<kDa<�Pa<�^a<Ama<�{a<b�a<e�a<��a<s�a<V�a<	�a<�a<�a<u�a<��a<%�a<'�a< �a<W�a<��a<9�a<�a<��a<˘a<D�a<Y�a<z�a<��a<��a<��a<�xa<�ja<h[a<�Ka<�<a</a<�#a<�a<Wa<.a<=a<�"a<I-a<3:a<!Ha<sVa<Hda<|pa<�za<�a<�a<9�a<��a<ˇa<��a<p�a<�}a<){a<�xa<�wa<�wa<�xa<�za<�}a<��a<'�a<�a<ڄa<�a<�~a<�wa<+na<ba<bTa<fEa<�6a<t(a<:a<�a<sa<�	a<
a<�a<Ba<K'a<5a<;Da<�  �  `Ta<ba<na<�wa<�~a<U�a<M�a<�a<e�a<�a<�}a<�za<�xa<Pwa<9wa<Rxa<�za<�}a<s�a<8�a<Q�a<��a<��a<B�a<݄a<�}a<�ta<�ha<�[a<�Ma<�?a<�2a<(a<P a<Ta<a<�a<['a<V2a<�?a<�Na<3^a<rma<I{a<4�a<��a<��a<Ûa<��a<Z�a<��a<��a<.�a<�a<v�a<�a<ȓa<��a<��a<d�a<w�a<V�a<S�a<0�a<�a<��a<M�a<��a<%�a<��a<�ta<gfa<LXa<�Ka<�Aa<�:a<G7a<�7a<N<a<ZDa<�Oa<�\a<ka<Jza<p�a<�a<>�a<
�a<T�a<��a<E�a<ͭa<X�a<,�a<��a<<�a<G�a<��a<�a<�a<�a<=�a<��a<��a<��a<_�a<�a<��a<_�a<:�a<��a<G�a<�sa<�da<�Va<�Ja<8Aa<Y;a<9a<�:a<@a<7Ia<�Ta<�ba<Cqa<�a<@�a<�a<7�a<��a<"�a<��a<&�a<�a<�a<��a<8�a<x�a<��a<�a<��a<M�a<ߡa<�a<�a<��a<	�a<۫a<m�a<U�a<��a<��a<9�a<'xa<Eia<}Za<�La<XAa<�8a<�3a<�2a<�5a<<a<�Ea<-Ra<$`a<{na<�|a<�a<��a<˛a<Z�a<.�a<��a<�a< �a<>�a<4�a<n�a<k�a<x�a<��a<�a<y�a<��a<O�a<��a<E�a<��a<G�a<i�a<ٍa<҄a<>ya<�ka<�\a<-Ma<>a<�0a<g%a<�a<xa<Ja<�a<L$a<�.a<t;a<xIa<�Wa<5ea<qa<�za<�a<ކa<��a<ƈa<Άa<݃a<9�a<�|a<iya<wa<�ua<�ua<*wa<fya<I|a<ta<�a<��a<l�a<ʂa<�~a<�wa<�na<�ba<iUa<�Fa<�7a<�)a<�a<<a<la<+a<a<�a<�a<�(a<�6a<�Ea<�  �  �Va<!da<koa<xxa<�~a<p�a<܃a<�a<��a<?}a<�ya<^va<�sa<Yra<ra<^sa<�ua<Yya<g}a<Áa<��a<v�a<��a<��a<�a<�~a<va<ka<`^a<Qa<�Ca<w7a<-a<�%a<�!a<q!a<W%a<�,a<@7a<Da<�Ra<jaa<�oa<}a<I�a<�a<)�a<��a<ۛa<��a<��a<ەa<��a<A�a<��a< �a<��a<ɐa<�a<�a<��a<$�a<ߤa<b�a<�a<"�a<ȡa<��a<�a<�a<�wa<-ja<�\a<�Pa<�Fa<�?a<�<a<C=a<�Aa<{Ia<YTa<aa<"oa<,}a<��a<}�a<2�a<`�a<��a<��a<H�a<@�a<��a<&�a<��a<S�a<V�a<a�a<�a<��a<t�a<�a<��a<˪a<{�a<�a<��a<תa<�a<w�a<��a<Ʉa<wa<�ha<p[a<�Oa<�Fa<�@a<M>a</@a<jEa<ANa<�Ya<�fa<�ta<`�a<E�a<?�a<��a<��a<<�a<H�a<��a<L�a<s�a<p�a<��a<��a<��a<�a<��a<]�a<m�a<ߠa<��a<�a<��a<��a<��a<��a<��a<�a<Y�a<�za<�la<�^a<�Qa<qFa<>a<P9a<8a<;a<JAa<�Ja<�Va<�ca<�qa<�~a<�a<ϔa<P�a<��a<�a<آa<}�a<�a<f�a<��a<��a<��a<l�a<��a<$�a<��a<t�a<b�a<��a<іa<�a<�a<��a<T�a<؅a<�za<na<�_a<�Pa<fBa<~5a<�*a<#a<�a<�a<N"a<m)a<�3a<�?a<Ma<�Za<jga<�ra<�{a<t�a<C�a<��a<Ɇa<B�a<�a<4|a<6xa<�ta<ra<�pa<�pa<Cra<�ta<'xa<�{a<Ma<��a<�a<ׁa<�~a<�xa<�oa<�da<�Wa<Ja<�;a<i.a<�"a<�a<�a<ua<wa<�a<�!a<`-a<�:a<�Ha<�  �  M[a<Yga<�qa<]ya<�~a<�a<B�a<Va<�{a<�wa</sa<.oa<�ka<#ja<�ia<<ka<na<Dra<$wa<O|a<5�a<�a<S�a<r�a< �a<�a<lxa<�na<�ba<�Va</Ja<�>a<�4a<".a<h*a<:*a<�-a<�4a<�>a<�Ja<wXa<_fa<�sa<�a<�a<��a<��a<Әa<�a<�a<ēa<��a<-�a<�a<��a<��a<i�a<Èa<x�a<?�a<��a<�a<Ӡa<i�a<��a<y�a<(�a<3�a<��a<�a<�|a<�oa<vca<�Wa<�Na<�Ha<bEa<�Ea<%Ja<vQa<|[a<�ga<�ta<́a<9�a<��a<��a<��a<��a<v�a<�a<�a<��a<��a<��a<ʕa<A�a<�a<��a<Ŕa<4�a<��a<:�a<�a<��a<+�a<{�a<��a<ҥa<��a<��a<�a<-|a<oa<rba<cWa<�Na<TIa<Ga<�Ha<�Ma<�Ua<�`a<ma<�ya<��a<}�a<c�a<ޣa<ʨa<�a<��a<^�a<��a<ʟa<�a<y�a<͒a<r�a<��a<x�a<Òa<V�a<��a<$�a<d�a<��a<,�a<��a<��a<Ξa<q�a<ҋa<ra<Kra<(ea<�Xa<NNa<�Fa<�Aa<�@a<�Ca<~Ia<GRa<}]a<�ia<�va<�a<Ía<��a<Ԝa<x�a<?�a<�a<��a<Зa<{�a<4�a<e�a<��a<#�a<L�a<�a<N�a<��a<b�a<R�a<Œa<�a<&�a<O�a<��a<�a<�}a<�qa<�da<�Va<8Ia<�<a<�2a<�+a<�'a<c'a<�*a<g1a<�:a<RFa<�Ra<*_a<�ja<,ua<+}a<��a<M�a<|�a<��a<�a<#{a<va</qa<�la<ja<xha<�ha<rja<�ma<�qa< va<eza<~a<7�a<S�a<8~a<Qya<�qa<�ga<&\a<9Oa<Ba<j5a<[*a<�!a<ca<Da<a<A!a<�)a<f4a<Aa<;Na<�  �  �`a<Nka<.ta<qza<B~a<Wa<�}a<�za<�ua<6pa<�ja<�ea<�aa<}_a<-_a<�`a<da<�ha<�na<,ua<S{a<��a<Y�a<�a<	�a<��a<^{a<�ra<�ha<�]a<~Ra<�Ga<R?a<�8a<�5a<�5a<�8a<a?a<wHa<�Sa<`a<�la<�xa<r�a<A�a<*�a<ߕa<��a<!�a<ˑa<)�a<'�a<)�a<a<#|a<{a<�{a<8~a<��a<�a<��a<2�a<i�a<u�a<��a<��a<��a<3�a<��a<ˍa<
�a<bwa<2la<�aa<hYa<`Sa<�Pa<'Qa<�Ta<�[a<�da<*pa<�{a<؇a<��a<�a<(�a<��a<��a<��a<եa<%�a<��a<��a<9�a<��a<��a<v�a<�a<q�a<��a<��a<��a<��a<�a<��a<��a<�a<��a<��a<��a<p�a<ɂa<�va<�ka<raa<�Ya<PTa<�Ra<�Sa<�Xa<`a<�ia<ua<��a<Q�a<t�a<�a<�a<k�a<"�a<V�a<��a<P�a<g�a<L�a<܌a<��a<Ʌa<�a<΅a<��a<�a<:�a<��a<��a<<�a</�a<8�a<|�a<C�a<b�a<#�a<V�a<Lya<wma<ba<�Xa<ZQa<Ma<FLa<wNa<Ta<!\a<Yfa<vqa<
}a<��a<E�a<ɘa<]�a<��a<�a<�a<T�a<5�a<��a<0�a<�~a<za<�wa<�va<�wa<jza<s~a<y�a<��a<Z�a<��a<��a<b�a<�a<~�a<�a<�va<�ja<&^a<�Qa<�Fa<I=a<b6a<�2a<�2a<�5a<�;a<?Da<�Na<�Ya<6ea<oa<@xa<�~a<��a<�a<��a<Za<+za<ta<�ma<�ga<�ba<j_a<�]a<^a< `a<�ca<�ha<xna<ta<+ya<�|a<i~a<�}a<2za<Rta<�ka<�aa<�Ua<�Ia<�>a<g4a<�,a<\'a<�%a<'a<�+a<�3a<�=a<Ia<�Ta<�  �  ga<�oa<
wa<�{a<�}a<�|a<�ya<�ta<ona<bga<v`a<dZa<�Ua<�Ra<qRa<(Ta<"Xa<�]a<�da<�la<_ta<H{a<��a<�a<�a<�a<�~a<�wa<^oa<�ea<�[a<�Ra<Ka<Ea<�Ba<�Ba<�Ea<�Ka<�Sa<�]a<�ha<ta<�~a<��a<��a<ݒa<��a<��a<q�a<��a<j�a<�~a<�xa<�sa<�oa<Yna<oa<�qa<wa<�}a<*�a<J�a<��a<��a<r�a<�a<�a<I�a<ښa<C�a<'�a<�a<va<�la<pea<,`a<�]a<)^a<�aa<�ga<�oa<�ya<3�a<��a<їa<�a<ڤa<��a<��a<#�a<��a<V�a<D�a<�a<n�a<�a<A|a<�za<[{a<Q~a<7�a<��a<��a<�a<�a<`�a<�a<A�a<��a<��a<��a<v�a<~�a<�a<�ua<�la<�ea<;aa<�_a<�`a< ea<�ka<Qta<A~a<��a<��a<�a<�a<(�a<ԧa<��a<>�a<؝a<�a<��a<3�a<��a<~|a<0ya<2xa<]ya<�|a<��a<\�a<}�a<��a<Ȝa<x�a<+�a<W�a<ʡa<��a<�a<�a<��a<�va<�la<gda<�]a<Za<CYa<M[a<8`a<kga<_pa<Hza<Y�a<��a<X�a<�a<�a<p�a<�a<p�a<�a<w�a<^�a<�ya<sa<�ma<�ja<�ia<Wka<�na<�sa<za<��a<�a<�a<��a<�a<��a<��a<�a<0|a<�qa<�fa<�[a<�Qa<OIa<-Ca<�?a<�?a<IBa<�Ga<6Oa<gXa<-ba<�ka<�ta<�{a<��a<��a<8�a<-a<za<^sa<�ka<da<]a<+Wa<Sa< Qa<fQa<Ta<�Xa<�^a<xea<�la<7sa<mxa<�{a<�|a<:{a<�va<0pa<�ga<�]a<Sa<�Ha<�?a<�8a<D4a<�2a<4a<f8a<6?a<Ha<ERa<�\a<�  �  uma<�ta<�ya<�|a<�|a<@za<]ua<jna<afa<�]a<aUa<Na<�Ha<wEa<�Da<�Fa<0Ka<�Qa<%Za<bca<�la<Gua<�|a<��a<f�a<_�a<�a<�|a<$va<Tna<fa<2^a<rWa<�Ra<TPa<qPa<?Sa<PXa<�_a<|ha<!ra<�{a<b�a<��a<��a<@�a<�a<b�a<M�a<��a<�|a<�ta<3ma<�fa<�ba<�`a<raa<�da<7ja<�qa<�za<��a<̍a<5�a<��a<G�a<6�a<0�a<Ξa<��a<��a<<�a<��a<�xa<#ra<�ma<�ka<�ka<oa<1ta<�{a<��a<��a<��a<(�a< �a<b�a<Y�a<x�a<I�a<��a<Ȓa<!�a<^�a<}ya<sa<�na<ma<�ma<;qa<�va<I~a<��a<ۏa<J�a<��a<�a<�a<��a<=�a<��a<��a<�a<��a<�a<ya<�ra<oa<pma<�na<$ra<�wa<ua<�a<ʐa<�a<�a<��a<�a<�a<�a<Ǟa<n�a<��a<�a<}a<Qua<roa<�ka<�ja<la<�oa<�ua<�}a<-�a<ˎa<Ėa<k�a<͡a<գa<�a<�a<<�a<��a<�a<��a<\xa<�pa<Lka<�ga<ga<�ha<ma<bsa<{a<��a<�a<y�a<��a<*�a<u�a<לa<Ҙa<M�a<�a<ڀa<>wa<;na<`fa<�`a<6]a<U\a<^a<ba<>ha<�oa<�wa<�a<��a<"�a<�a<��a<x�a<�a<�a<Vya<�oa<\fa<�]a<Va<�Pa<�Ma<cMa<�Oa<"Ta<�Za<�ba<�ja<�ra<�ya<6a<�a<s�a<
�a<U{a<Ita<�ka<�ba<wYa<#Qa<EJa<�Ea<wCa<�Ca<�Fa<La<[Sa<�[a<ada<�la<�sa<�xa<�{a<|a<�ya<�ta<�ma<�ea<�\a<�Sa<La<�Ea<	Ba<�@a<�Aa<�Ea<rKa<;Sa<\a<ea<�  �  �sa<ya<z|a<r}a<�{a<Pwa<wpa<�ga<^a<�Sa<.Ja<�Aa<~;a<�7a<�6a<9a<7>a<�Ea<9Oa<�Ya<�da<(oa<xa<4a<��a<��a<�a<Ła<�|a<�va<�oa<�ia<�ca<�_a<�]a<^a<�`a<2ea<�ka<sa<+{a<�a<�a<o�a<��a<e�a<_�a<a<ޅa<r}a<�sa<pja<�aa<\Za<QUa<�Ra<�Sa<5Wa<�]a<%fa<kpa<k{a<��a<��a<$�a<z�a<'�a<�a<a�a<v�a<˘a<�a<�a<{�a<�~a<	{a<0ya<�ya<3|a<׀a<��a<�a<��a<{�a<0�a</�a<ߧa<ۦa<<�a<��a<Ȕa<�a<��a<�va<wma<.fa<9aa<1_a<
`a<�ca<eja<�ra<�|a<_�a<��a<��a<�a<ݦa<%�a<��a<��a<Ƞa<R�a<�a<ŋa<:�a<�a<d|a< {a<�{a<)a<)�a<z�a<��a<Řa<5�a<:�a<R�a<��a<֥a<�a<��a<�a<��a<|a<�qa<
ia<Bba<�]a<�\a<>^a<�ba<�ia<�ra<�|a<�a<��a<�a<S�a<$�a<b�a<�a<�a<i�a<m�a<�a<��a<Q}a<exa<lua<�ta<Hva<�ya<Aa<��a<��a<^�a<-�a<F�a<@�a<��a<6�a<2�a<ߌa<��a<�wa<�la<�ba<�Ya<GSa<aOa<�Na<�Pa<iUa<w\a<@ea<�na<uxa<�a<K�a<L�a<��a<]�a<s�a<`�a<��a<�xa<�pa<Bia<�ba<^a<][a<�Za<�\a<�`a<;fa<�la<{sa<�ya<�~a<f�a<��a<��a<�}a<wa<Una<+da<NYa<�Na< Ea<i=a<8a<�5a<6a<�9a<�?a<Ha<�Qa<�[a<�ea<�na<�ua<�za<�|a<|a<�xa<�sa<Tma<fa<�^a<%Xa<�Ra<fOa<9Na<7Oa<�Ra<�Wa<=^a<�ea<ma<�  �  xya<}a<�~a<�}a<cza<]ta<�ka<�aa<Va<�Ja<�?a<36a</a<�*a<�)a<-,a<�1a<U:a<�Da<�Pa<*]a<;ia<�sa<�|a<ła<��a<��a<$�a<�a</~a< ya<�sa<Woa<la<�ja<�ja<�la<�pa<Hva<�|a<^�a<ǉa<@�a<֒a<w�a<:�a<��a<3�a<��a<�va<vka<�`a<�Va<|Na<�Ha<�Ea<�Fa<pJa<�Qa<[a<�fa<�ra<�a<:�a<a�a<�a<âa<��a<��a<s�a<V�a<�a<��a<�a<��a<K�a<�a<I�a<`�a<J�a<[�a<D�a<*�a<��a<¦a<�a<�a<�a<ߠa<Иa<�a<��a<�wa<zla<ba<�Ya<[Ta<3Ra<Sa<`Wa<�^a<2ha<xsa<;a<&�a<a<Ξa<j�a<e�a<ժa<��a<S�a<]�a<��a<��a<:�a<؋a<݈a<߇a<��a<.�a<J�a<��a<Z�a<��a<�a<=�a<��a<n�a<��a<'�a<0�a<��a<�~a<�ra<Tga<q]a<�Ua<�Pa<�Oa<WQa<�Va<V^a<`ha<�sa<Ja<��a<��a<��a</�a<Q�a<��a<f�a<o�a<�a<��a<�a<��a<��a<�a<��a<��a<��a<��a<K�a<ٔa<�a<Z�a<��a<�a<r�a<k�a<��a<��a<)|a<�oa<Kca<�Wa<�Ma<�Fa<`Ba<Aa<�Ca<rIa<WQa<o[a<2fa<qqa<�{a<��a<P�a<I�a<�a<��a<[�a<#�a<܀a<Iza<�sa<una<Ija<ha<�ga<ia<:la<�pa<�ua<&{a<�a<��a<>�a<��a</�a<u{a<�ra<�ha<�\a<mPa<�Da<�9a<:1a<0+a<�(a<)a<-a<4a<H=a<DHa<�Sa<m_a<�ia<�ra<ya<�|a<&~a<�|a<gya<\ta<�na<�ha<"ca<�^a<�[a<�Za<�[a<�^a<�ba<Gha<Xna<7ta<�  �  ~a<Q�a<p�a<9~a<6ya<�qa<�ga<\a<MOa<�Ba<X6a<,a<K$a<�a<�a<9!a<J'a<V0a<�;a<Ia<�Va<�ca<
pa<Bza<��a<&�a<��a<��a<هa<��a<��a<�|a<ya<iva<)ua<sua<~wa<�za<�a<ӄa<R�a<p�a<i�a<��a<��a<�a<܍a<�a<|a<pa<Bda<6Xa<�La<Da<�=a<�:a<R;a<�?a<Ga<ZQa<�]a<{ka<Hya<v�a<�a<��a<|�a<��a<�a<y�a<פa<�a<��a<H�a<��a<ݑa<��a<�a<ђa<�a<R�a<��a<��a<ǧa<��a<&�a<��a<o�a<��a<;�a<�a<@}a<8pa<�ca<8Xa<^Oa<mIa<�Fa<�Ga<�La<bTa<�^a<;ka<Lxa<V�a<��a<�a<�a<��a<L�a<��a<Ϊa<V�a<ܢa<%�a<��a<��a<��a<��a<7�a<f�a<ߘa<�a<��a<�a<��a<}�a<J�a<��a<^�a<q�a<"�a<�a<�wa<�ja<^a<<Sa<	Ka<�Ea<5Da<`Fa<�Ka<TTa<Q_a<�ka<�xa<_�a<Ӑa<\�a<c�a<٥a<��a<��a<[�a<U�a<��a<Ėa<c�a<�a<Ìa<"�a<8�a<��a<D�a<o�a<ϛa<��a<��a<h�a<-�a<S�a<��a<��a<�a<va<Qha<�Za<Na<�Ca<�;a<+7a<46a<�8a<�>a<�Ga<�Ra<�^a<6ka<�va<=�a<g�a< �a<�a</�a<a�a<��a<��a<F�a<}a<axa<�ta<�ra<Kra<usa<va<�ya<�}a<��a<(�a<M�a<`�a<_�a<��a<8ya<Ooa<wca<TVa<�Ha<�;a<�/a<�&a<D a<;a<	a<["a<�)a<�3a<@a<�La<�Ya<�ea<�oa<�wa<}a<�a<�a<�}a<Rza<�ua<qa<�la<�ha<�fa<�ea<jfa<�ha<hla<�pa<�ua<Xza<�  �  ��a<܂a<��a<V~a<?xa<uoa<tda<�Wa<�Ia<$<a<M/a<J$a<�a<a<�a<�a<�a<�(a<�4a<�Ba<�Qa<�_a< ma<Exa<E�a<�a<!�a<��a<��a<��a<d�a<<�a<P�a<F~a<h}a<�}a<�a<k�a<��a<��a<��a<��a<��a<��a<��a<�a<q�a<��a<rxa<�ka<�^a<{Qa<�Ea<�;a<H5a<2a<�2a<7a<�>a<Ja<'Wa<�ea<�ta<��a<q�a<�a<.�a<k�a<+�a<��a<��a<0�a<��a<3�a<��a<�a<ژa<.�a<��a<j�a<�a<ߤa<Ĩa<��a<a�a<�a<(�a<ڤa<��a<O�a<څa<?xa<4ja<�\a<�Pa<!Ga<�@a<�=a<L?a<(Da<�La<�Wa<�da<�ra<Հa<�a<��a<�a<��a<u�a<�a<<�a<�a<`�a<z�a<Ԡa<��a<��a<њa<l�a<�a<	�a<��a<J�a<ͪa<!�a<	�a<��a<ڨa<g�a<>�a<ڍa<��a<�ra<Ida<�Va<�Ka<�Ba<K=a<f;a<�=a<�Ca<�La<SXa<�ea<�sa<2�a<Ǎa<]�a<��a<1�a<�a<éa<&�a<M�a<\�a<g�a<��a<a<�a<k�a<G�a<&�a<B�a<��a<#�a<�a<��a<��a<�a<!�a<L�a<��a<ua<^qa<�ba<
Ta<�Fa<~;a<?3a<m.a<q-a<o0a<�6a<k@a<�Ka<"Ya<mfa<;sa<�~a<ևa<��a<��a<:�a<g�a<��a<�a<R�a<��a<�a<�|a<{a<�za<d{a<X}a<P�a<{�a<��a<�a<-�a<#�a<ԅa<�a<Zwa<dla<m_a<TQa<�Ba<�4a<}(a<ca<�a<qa<aa<�a<�!a<�,a<�9a<iGa<Ua<+ba<uma<�va<}a<Āa<<�a<L�a<�~a<L{a<]wa<�sa<�pa<�na<�ma<�na<tpa<�sa<Hwa<D{a<
a<�  �  ȃa<E�a<��a<H~a<twa<na<hba<�Ta<�Fa<$8a<�*a<=a<�a<�a<ga<Ga<�a<�#a<t0a<	?a<3Na<E]a<ka<wa<��a<��a<�a<�a<�a<l�a< �a<a�a<�a<)�a<k�a<��a<z�a<L�a<�a<��a<��a<=�a<��a<�a<�a<��a<x�a<�a<2va<�ha<�Za<EMa<Aa<�6a<�/a<�,a<:-a<�1a<�9a<DEa<�Ra<ba<oqa<_�a<��a<�a<��a<�a<X�a<]�a<r�a<o�a<��a<~�a<Ša<Ϟa<�a<9�a<��a<�a<=�a<��a<ƫa<�a<��a<��a<{�a<M�a<��a<w�a<i�a<�ta<Xfa<*Xa<�Ka<�Aa<{;a<�8a<�9a<�>a<{Ga<Sa<�`a<\oa<!~a<�a</�a<�a<k�a<<�a<d�a<O�a<��a<�a<��a<M�a<��a<��a<�a<d�a<	�a<��a<��a<�a<��a<D�a<s�a<l�a<˨a<��a<ߗa<ϋa<�}a<!oa<I`a<^Ra<uFa<J=a<�7a<6a<j8a<E>a<�Ga<�Sa<�aa<Lpa<�~a<݋a<+�a<
�a<c�a<�a<G�a<k�a<+�a<�a<��a<F�a<��a<�a<��a<4�a<�a<��a<��a<u�a<��a<��a<ͦa<��a<��a<S�a<T�a<5}a<mna<_a<�Oa<Ba<[6a<�-a<)a<(a<+a<�1a<�;a<�Ga<dUa<\ca<�pa<�|a<Նa<;�a<(�a<g�a<C�a<<�a<*�a<F�a<@�a<��a<ʁa<�a<�a<D�a<��a<�a<I�a<a<f�a<ɋa<3�a<(�a<oa<=va<�ja<�\a<Na<�>a<O0a<�#a<"a<Ua<a<�a<�a<�a<((a<u5a<�Ca<iRa<`a<la<�ua<�|a<��a<��a<_�a<��a<�~a<m{a</xa<yua<�sa<sa<�sa<`ua<xa<^{a<�~a<��a<�  �  P�a<9�a<ߋa<�a<�|a<�oa<�_a<�Ma<�9a<8&a<�a<a<#�`<��`<��`<��`<��`<�	a<�a<C.a<�Ba<#Wa<�ia<�ya<��a<�a<��a<U�a<��a<��a<��a<C�a<P�a<��a<&�a<��a<*�a<p�a<��a<4�a<�a<۠a<F�a<�a<P�a<��a<J�a<��a<�ra<i`a<Ma<I:a<.)a<a<Pa<a<�a<�a<�a<,-a<�?a<�Sa<�ha<�|a<��a<��a<��a<��a<��a<Ƿa<ٶa<(�a<��a<��a<Ʃa<C�a<~�a<��a<�a<"�a<��a<��a<p�a<D�a<�a<7�a<t�a<3�a<b�a<�a<l~a<�ja<�Va<�Ca<�2a<%a<a<�a<�a<� a<�,a<H<a<�Na<�ba<�va<��a< �a<ϧa<��a<�a<�a<��a<w�a<�a<$�a<N�a<�a<ݨa<F�a<��a<s�a<��a<)�a< �a<U�a<�a<�a<g�a<5�a<��a<>�a<�a<Twa<ca<�Na<<a<�+a<}a<�a<"a<�a<
!a<(.a<�>a<�Qa<xea<$ya<�a<l�a<��a<(�a<;�a<#�a<��a<ܲa<�a<�a<C�a<�a<`�a<��a<��a<ͤa<اa<n�a<�a<��a<�a<o�a<]�a<��a<��a<��a< za<<fa<YQa<=a<T*a<�a<Fa<ya<Ya<a<[a<3#a<4a<�Fa<EZa<�la<)}a<1�a<h�a</�a<\�a<��a<�a<&�a<��a<��a<܌a<}�a<�a<\�a<�a<Y�a<K�a<��a<��a<��a<*�a<ϓa<��a<��a<]ya<|ia<aWa<GCa<�.a<a<�	a<��`<@�`<��`<�`<��`<Ka<�a<�"a<�6a<�Ja<�\a<Ama<�za<f�a<��a<s�a<ߍa<��a<F�a<B�a<i�a<*}a<{a<�za<{a<}a<P�a<'�a<>�a<ًa<�  �  .�a<��a<��a<�a<}a<vpa<�`a<�Na<~;a<(a<�a<aa<e�`<��`<��`<��`<�`<�a<�a<0a<MDa<6Xa<�ja<Oza<�a<�a<j�a<��a<\�a<.�a< �a<v�a<+�a<Èa<��a<�a<�a<9�a<��a<��a<��a<��a<\�a<��a<4�a<�a<��a<��a<�sa<�aa<�Na<<a<g+a<ha<�a<a<�a<Xa< a<f/a<oAa<�Ua<ja<�}a<l�a<H�a<��a<��a<��a<�a<��a<ɲa<	�a<�a<��a<�a<£a<�a<�a<�a<�a<%�a<�a<�a<H�a<�a<x�a<i�a<ןa<��a<~a<Ela<�Xa<�Ea<�4a<H'a<�a<�a<�a<#a<�.a<t>a<�Pa<pda< xa<��a<ؚa<�a<��a<ڷa<��a<w�a<(�a<��a<v�a<\�a<רa<u�a<��a<(�a<?�a<��a<q�a<��a<��a<]�a<��a<�a<;�a<�a<�a<�a<sxa<�da<�Pa<4>a<:.a<�!a<�a<3a<Ra<I#a<l0a<�@a<eSa<�fa<8za<ދa<��a<צa<)�a<�a<z�a<n�a<��a<��a<9�a<�a<ݡa<̟a<;�a<@�a<��a<��a<ީa<��a<��a<�a<�a<A�a<ǥa<ښa<U�a<�za<xga<Sa<�>a<�,a<�a<�a<ta<]
a<�a<�a<m%a<�5a<�Ha<�[a<�ma<~a<��a<��a<!�a<�a<"�a<��a<Ƙa<�a<�a<��a<=�a<+�a<��a<υa<!�a<q�a<�a<d�a<��a<o�a<��a<��a<�a<�ya<rja<rXa<�Da<�0a<a<�a<��`<��`<��`<��`< �`<�a<�a<�$a<H8a<�Ka<�]a<�ma<{a<t�a<n�a<��a<Ɍa<a�a<Άa<��a<x~a<�za<�xa<�wa<�xa<�za<K~a<p�a<��a<��a<�  �  f�a<�a<��a<�a<~a<lra<�ca<�Ra<%@a<j-a<�a<3a<�a<��`<��`<��`<Ka<�a<�"a<J5a<�Ha<�[a<Rma<	|a<��a<��a</�a<��a<i�a<j�a<8�a<�a<��a<S�a<�a<?�a<{�a<�a<֋a<o�a<@�a<Y�a<��a<�a<��a<�a<ԑa<څa<�va<�ea<�Sa<�Aa<�1a<k$a<�a</a<�a<ya<1'a<�5a<Ga<�Za<.na<�a<�a<��a<#�a<�a<4�a<��a<i�a<��a<��a<U�a<;�a<��a<�a<e�a<{�a<��a<<�a<E�a<0�a<��a<�a<��a<$�a< �a<x�a<��a<��a<�pa<�]a<_Ka<�;a<l.a<�%a<�!a<�#a<9*a<�5a<�Da<Va<.ia<�{a<��a<�a<1�a<�a<��a<иa<ȷa<��a<*�a<�a<[�a<r�a<��a<՞a<��a<աa<q�a< �a<�a<p�a<��a<Ʒa<�a<K�a<�a<ܜa<ލa<1|a<]ia<2Va<LDa<5a<�(a<�!a<Oa<x"a<x*a<7a<�Fa<�Xa<hka<�}a<��a<��a<��a<�a<��a<t�a<|�a<��a<Ũa<��a<�a<n�a<+�a<��a<֙a<>�a<'�a<��a<V�a<>�a<��a<~�a<��a<,�a<�a<��a<,~a<}ka<
Xa<fDa<�2a<�#a<�a<�a<wa<�a<�a<�+a<�;a<�Ma<�_a<qa<��a<�a<
�a<��a<��a<��a<{�a<��a<�a<W�a<R�a<ـa<z~a<	~a<da<�a<ʅa<1�a<��a<��a<D�a<5�a<.�a<��a<r{a<%ma<�[a<	Ia<�5a<�"a<�a<a<��`<��`<�`<H�`<}
a<a<<*a<=a<�Oa<aa<pa<|a<��a<��a<@�a<�a<�a<S�a<5}a<yxa<�ta<(ra<!qa<ra<kta<8xa< }a</�a<��a<�  �  ݅a<�a<K�a<3�a<�a<`ua<-ha<�Xa<SGa<�5a<�%a<�a<a<�a<a<�a<�a<�a<	,a<�=a<�Oa<�aa<Gqa<�~a<�a<}�a<��a<S�a<��a<�a<��a<&�a<J{a<�wa<�ua<5va<xxa<�|a<��a<^�a<p�a<Жa<�a<��a<��a<�a<�a<7�a<�{a<&la<G[a<�Ja<;a<#/a<}&a<)"a<�"a</(a<2a<�?a<TPa<Uba<�ta<9�a<d�a<�a<תa<7�a<��a<��a<�a<�a<��a<+�a<@�a<��a<�a<g�a<��a<�a<\�a<��a<ƪa<��a<��a<δa<Ʋa<)�a<
�a<w�a<��a<dwa<�ea<�Ta<�Ea<�9a<�1a< .a<|/a<�5a<?@a<@Na<�^a<{pa<'�a<J�a< �a<ߪa<�a<ӵa<�a<p�a<ծa<�a<Ţa<�a<�a<�a<ɓa<��a<[�a<�a<��a<��a<l�a<	�a<ȴa<Ҵa<a�a<c�a<Пa<9�a<>�a<�pa<�^a<�Ma<f?a<k4a<�-a<^+a<D.a<�5a<9Aa<Pa<�`a<Yra<��a<��a<d�a<٨a<��a<�a<$�a<��a<r�a<D�a<�a<<�a<��a<(�a<��a<юa<%�a<�a<��a<��a<��a<��a<�a<��a<��a</�a<�a<)�a<�qa<�_a<�Ma<�<a<�.a<s$a<�a<ya<[!a<�)a<�5a<�Da<NUa<Afa<Ava<�a<*�a<��a<՚a<`�a<�a<$�a<�a<�a<.�a<Xza<�ua<ysa<sa<�ta<xa<�|a<��a<�a<��a<ɏa<d�a<ύa<��a<~a<�pa<uaa<�Oa<�=a<C,a<�a<)a<�a<�a<�a<�
a<�a<�"a<3a<RDa<�Ua<�ea<"sa<�}a<ބa<j�a<v�a<ąa<�a<;{a<�ta<oa<?ja<$ga<fa<ga<�ia<�na<�ta<�za<�a<�  �  �a<��a<�a<�a<]�a<Iya<�ma<`a<�Pa<�@a<2a<-%a<ka<�a<Xa<Ka<�a<*a<J8a<Ha<�Xa<�ha<}va<1�a<'�a<Ďa<��a<��a<�a<��a<�{a<`ta<bna<�ia<�ga<�ga<~ja<�oa<8va<�~a<E�a<f�a<j�a</�a<�a<^�a<l�a<��a<��a<9ta<ea<LVa<pHa<=a<
5a<F1a<�1a<�6a<@a<�La<\a<Qla<}a<��a<
�a<��a<c�a<�a<��a<m�a<إa<��a<Z�a<�a<�a<��a<��a<)�a<�a<�a<p�a<Q�a</�a<?�a<̮a<�a<رa</�a<?�a<�a<Z�a<�a<1pa<�`a<�Ra<�Ga<F@a<E=a<�>a<?Da<Na<�Za<ja<�ya<ˉa<
�a<�a<�a<��a<ʳa<�a<��a<�a<|�a<��a<H�a<��a<ֆa<t�a<k�a<�a<.�a<$�a<�a<i�a<��a<��a<��a<�a<-�a<��a<͗a<��a<�ya<�ia<qZa<Ma<�Ba<w<a<�:a<=a<Da<�Na<G\a<nka<4{a<��a<ؗa<ܢa< �a<�a<l�a<��a<�a<�a<,�a<#�a<S�a<�a<�a<2a<׀a<�a<��a<őa<W�a<H�a<�a<��a<$�a<	�a<��a<}�a<Q�a<
za<Tia<Ya<�Ia<�<a< 3a<�-a<�,a<�/a<�7a<�Ba<�Pa<J_a<�na<�|a<��a<��a<L�a<��a<�a<��a<�a<��a<V|a<�sa<7ma<�ga<,ea<�da<�fa<'ka<�pa<=xa<~a<��a<��a<��a<��a<��a<5�a<�ua<Hha<�Xa<"Ha<V8a<�)a<aa<pa<
a<�a<Ja<�"a<_/a<">a<�Ma<a]a<cka<=wa<�a<��a<c�a<u�a<�a<Cya<�qa<�ia<lba<�\a<Ya<�Wa<�Xa<}\a<�aa<*ia<5qa<�xa<�  �  �xa<�a<�a<o�a<�a<#}a<ta<Vha<?[a<MMa<,@a<�4a<G,a<'a<�%a<�(a<�/a<{9a<�Ea<'Ta<�ba<Qpa<U|a<u�a<d�a<��a<j�a<+�a<6�a<�xa<�oa<�fa<+_a<�Ya<�Va<�Va<�Ya<�_a<�ga<�qa<5|a<��a<ݏa<֖a<�a<��a<��a<x�a<�a<I}a<zpa< ca<)Wa<HMa<'Fa<�Ba<\Ca<�Ga<iPa<�[a<ia<�wa<f�a<��a<�a<"�a<��a<��a<��a< �a<O�a<�a<��a<΁a<Vza<Cua<�ra<sa<�va<�|a<��a<�a<�a<2�a<	�a<6�a<��a<<�a<@�a<"�a<�a<�a< |a<Lna<#ba<aXa<�Qa<�Na<Pa<1Ua<�]a<Bia<�va<لa<Z�a<��a<E�a<��a<ѱa<�a<?�a<��a<��a<��a<c�a<��a<�za<va<Gta<�ua<�ya<X�a<Ԉa<<�a<�a<��a<��a<��a<��a<խa<��a<�a<��a<|�a<va<�ha<�\a<�Sa<�Ma<-La<~Na<�Ta<^a<�ia<�wa<m�a<^�a<��a<#�a<`�a<��a<��a<��a<L�a<�a<�a<��a<ya<�ra<�na<na<Hpa<ua<1|a<�a<E�a<��a<��a<2�a<��a<a�a<�a<F�a<;�a<�a<�ta<�ea<NXa<�La<Da< ?a< >a<+Aa<Ha<�Qa<�]a<�ja<�wa<Ãa<��a<`�a<�a<��a<�a<W�a<e�a<!za<�oa<�ea<r]a<�Wa<Ta<�Sa<�Va<�[a<=ca<�ka<0ua<�}a<,�a<ɉa<��a<��a<3�a<�{a<�oa<rba<Ta<�Ea<$9a<�.a<�'a<�$a<b%a<8*a<�2a<�=a<�Ja<�Xa<�ea<�qa<h{a<��a<��a<��a<�a<�xa<pa<0fa<�\a<�Sa<�La<SHa<�Fa<Ha<`La<)Sa<�[a<�ea<toa<�  �  pa<�ya<��a<��a<��a<��a<}za<�pa<)fa<fZa<IOa<pEa<�=a<�9a<v8a<;a<�@a<�Ia<�Ta<�`a<!ma<pxa<8�a<��a<��a<:�a<��a<فa<Pxa<�ma<Yba<�Wa<�Na<Ha<�Da<eDa<�Ga<�Na<?Xa<�ca<Tpa<�|a<T�a<�a<:�a<��a<�a<.�a<)�a<��a< |a<�pa<�fa<^a<?Xa<kUa<Va<*Za<Maa<~ka<wa<̃a<�a<5�a<�a<��a<L�a<��a<�a<�a<��a<z�a<�|a<Sra<Gia<Mca<O`a<�`a<�da<�ka<�ua<��a<��a<�a<i�a<"�a<��a<�a<N�a<��a<۞a<:�a<��a<�|a<Nra<�ia<�ca<paa<�ba<
ga<�na<�xa<�a<�a<-�a<F�a<k�a<��a<7�a<�a<��a<V�a<|�a<��a<�{a<�qa<.ia<�ca<�aa<nca<3ha<pa<5za<��a<l�a<<�a<ǥa<)�a<��a<j�a<m�a<��a<��a<h�a<7�a<�wa<Wma<\ea<{`a<�^a<�`a<fa<`na<�xa<,�a<ݏa<��a<��a<q�a<~�a<��a<�a<��a<g�a<�a<�}a<�ra<�ha<"aa<�\a<�[a<C^a<�ca<�la<�va<b�a<��a<��a<J�a<@�a<f�a<D�a<��a<z�a<t�a<e�a<�sa<�ga<�]a<4Va<�Qa<�Pa<WSa<�Xa<�aa<�ka<�va<��a<?�a<��a<�a<8�a<3�a<O�a<�a<�za<na<�aa<[Va<dLa<�Ea<�Aa<�Aa<�Da<�Ja<Ta<�^a<ja<�ta<�~a<��a<��a<��a<>�a<'�a<�wa<�la<s`a<BTa<KIa<@a<:a<.7a<�7a<<a<<Ca<�La<�Wa<�ca<�na<�xa<�a<��a<��a<��a<5za<�pa<�ea<�Ya<#Na<�Ca<b;a<96a<24a<�5a<�:a<�Ba<BMa<�Xa<�da<�  �  �ga<�sa<�|a<�a<��a<��a<i�a<vya<�pa<1ga<�]a<�Ua<�Oa<�Ka<�Ja<+Ma<-Ra<�Ya<�ba<ma<Cwa<q�a<��a<׋a<�a<A�a<?�a<�za<\oa<{ba<�Ta<hHa<�=a< 6a<�1a<�1a<�5a<k=a<*Ha<JUa<da<�ra<��a<�a<O�a<�a<��a<d�a<�a<�a<i�a<y~a<va<�na<ja<�ga<Oha<la<Ira<�za<Єa<N�a<|�a<G�a<��a<�a<ҫa<ާa<��a<J�a<�a<x|a<�na<bba<RXa<Qa<�Ma<8Na<�Ra<�Za<�ea<�ra<0�a<َa<K�a<��a<��a<?�a<)�a<̬a<��a<'�a<��a<�a<�a<�za<
va<�sa<�ta<�xa<a<w�a<��a<Ԛa<��a<t�a<0�a<�a<��a<r�a<��a<�a<�a<�za<#ma<3aa<�Wa<�Qa<-Oa<�Pa<�Va<�_a<1ka<�xa<��a<œa<w�a<t�a<<�a<{�a<��a<z�a<!�a< �a<�a<\�a<�}a<�va<�ra<Eqa<sa<pwa<V~a<��a<u�a<�a<��a<��a<��a<�a<��a<Ңa<֘a<t�a<�~a<ipa<*ca<�Wa<6Oa<'Ja<Ia<�Ka<�Ra<r\a<zha<va<��a<%�a<ךa<S�a<��a<2�a</�a<A�a<��a<��a</�a<5wa<xna<ha<da<ca<Bea<�ia<�pa<Pya<J�a<��a<S�a<4�a<3�a<��a<��a<*�a<�~a<qa<~ba<�Sa<lFa<r;a<W3a</a<�.a<�2a<6:a<�Da<�Pa<~^a<�ka<lwa< �a<��a<��a<�a<2�a<ta<�va<ula<\ba<Ya<[Qa<)La<�Ia<'Ja<�Ma<�Sa<�[a<
ea<�na<�wa<�~a<T�a<��a<a<}a<-ta<yha<9[a<Ma<V?a<e3a<�)a<�#a<�!a<m#a<C)a<w2a<A>a<�Ka<1Za<�  �  z_a<uma<?ya<��a<D�a<��a<��a<�a<_za<�ra<Yka<�da<�_a<�\a<
\a<�]a<6ba<Cha<	pa<jxa<a�a<a�a<6�a<f�a<��a<J�a<�a<_ta<�fa<aWa<IHa<:a<�-a<'%a<s a<@ a<R$a<�,a<�8a<�Ga<8Xa<ia<ya<��a<p�a<�a<t�a<<�a<ٜa<�a<ؑa<ۊa<�a<m~a<pza<�xa<lya<�|a<��a<�a<`�a< �a<�a<q�a<��a<��a<�a<<�a<��a<�a<s�a<�pa<�aa<ZSa<�Ga<�?a<#<a<�<a<�Aa<�Ja<UWa<*fa<�ua<�a<z�a<�a<]�a<
�a<x�a<@�a<C�a<�a<��a<�a<}�a<Ȋa<��a< �a<��a<�a<(�a<��a<��a<��a<��a<ְa<��a<вa<��a<	�a<��a<-�a<�~a<�na<Z_a<�Qa<�Fa<@a<�=a<r?a<�Ea<�Oa<3]a<Dla<|a<��a<I�a<��a<��a<�a<�a<��a<��a<��a<ԛa<��a<��a<�a<��a<s�a<��a<}�a<�a<�a<כa<&�a<z�a<��a<�a<��a<��a<�a<7�a<ƃa<�sa<�ca<�Ta<�Ga<<>a<�8a<�7a<�:a<8Ba<@Ma<+[a<Cja<�ya<��a<S�a<s�a<��a<��a<�a<'�a<ݝa<�a<��a<�a<�}a<dxa<ua<0ta<�ua<�ya<�~a<��a<��a<d�a<}�a<C�a<��a<	�a<�a<�a<Iwa<�ga<�Va<�Fa<e7a<+a<"a<�a<da<�!a<!*a<�5a<Da<+Sa<�ba<�pa<}|a<\�a<~�a<b�a<��a<#�a<fa<�wa<Ooa<rga<Maa<�\a<�Za<[a<�]a<�ba<\ia<qa<�xa<<a<0�a<��a<ąa<k�a<�ya<9na<�`a<�Pa<�@a<�1a<�#a<;a<]a<a<�a<qa<�"a<G0a<�?a<�Oa<�  �   Xa<�ga<qua<�a<��a<��a<؉a<�a<y�a<�|a<�va<jqa<*ma<�ja<Yja<�ka<�oa<�ta<#{a<�a<�a<"�a<�a<L�a<��a<(�a<�{a<�na<�^a<�Ma<=a<>-a<* a<�a<fa< a<�a<�a<�+a<�;a<�Ma<l`a<Yra<�a<_�a<-�a<|�a<6�a<ˡa<�a<��a<7�a<�a<n�a<5�a<��a<��a<_�a<�a<�a<�a<�a< �a<��a<ίa<�a<p�a<k�a<Ėa<��a<xa<�fa<�Ua<=Fa<�9a<01a<�,a<�-a<,3a<�<a<oJa<�Za<3la<�}a<n�a<��a<��a<үa<$�a<�a<ײa<��a<�a<Ңa<�a<�a<��a<S�a<��a<��a<�a<��a<��a<�a<
�a<_�a<�a<l�a<:�a<q�a<g�a<�a<�ua<�ca<�Ra</Da<�8a<;1a<\.a<�0a<j7a<WBa<�Pa<daa<�ra<@�a<ɓa<�a<�a<~�a<m�a<�a<��a<��a<��a<@�a<[�a<��a<��a<Ɛa<ɑa<ؔa<|�a<7�a<S�a<�a<?�a<��a<�a<�a<x�a<P�a<a�a<	|a<?ja<�Xa< Ha<:a<�/a<�)a<F(a<�+a<4a<@a<+Oa<�_a<Eqa<��a<d�a<a�a<Фa<��a<��a<�a<��a<̞a<�a<�a<��a<)�a<[�a<y�a<��a<��a<�a<i�a<��a<��a<��a<q�a<0�a<_�a<�a<0�a<�pa<*_a<�La<�:a<J*a<�a<ta<ba<La<a<6a<�(a<�8a<�Ia<�Za<�ja<xa<��a<C�a<�a<I�a<��a<�a<�a<8za<�sa<�na<�ja<ia<Iia<�ka<�oa<
ua<{a<ـa<��a<��a<9�a<a�a<�a<va<�ha<lYa<�Ga<;6a<9%a<ha<�
a<�a<� a<a<
a<7a<�#a<�4a<}Fa<�  �  (Ra<�ca<�ra<o~a<��a<V�a<�a<��a<��a<�a<[a< {a<�wa<�ua<dua<�va<�ya<6~a<a�a<�a<ߍa<a�a<ʒa<\�a<��a<a�a<�xa<�ia<�Xa<�Fa<34a<�#a<�a<a<�a<�a<�	a<�a<�!a<�2a<�Ea<�Ya<�la<a~a<�a<<�a<�a< �a<[�a<�a<�a<��a<ޘa<A�a<�a<��a<��a<O�a<��a<%�a<ѣa<~�a<?�a<V�a<�a<��a<��a<�a<6�a<I�a<eqa<�^a<vLa<W<a<�.a<u%a<� a<�!a<�'a<O2a<�@a<�Qa<�da<�wa<��a<E�a<�a<`�a<�a<l�a<�a<1�a<�a<�a<=�a<5�a<��a<c�a<��a</�a<��a<Y�a<h�a<A�a<׶a<��a<��a<��a<��a<��a<W�a<7�a<�na<�[a<�Ia<:a<`-a<m%a<M"a<�$a<�+a<8a<*Ga<�Xa<�ka<F~a<��a<�a<��a<x�a<ʵa<��a<Z�a<Աa<��a<ŧa<��a<*�a<��a<ӛa<Ϝa<!�a<�a<w�a<\�a<��a<��a<;�a<�a<��a<��a<)�a<��a<�ua<�ba<�Oa<S>a<�/a<($a<�a<Ca<- a<�(a<	6a<�Ea< Xa<�ja<�|a<��a<�a<ޣa<+�a<�a<��a<ϩa<G�a<��a<��a<͔a<�a<V�a<w�a<}�a<��a<1�a<R�a<|�a<��a<c�a<��a<Ҝa<��a<��a<�|a<�ka<�Xa<�Da<|1a<e a<	a<�a<`a<Ya<ra<�a<Ba<�/a<
Ba<=Ta<�ea<�ta<��a<ωa<��a<ːa<ȏa<��a<Ňa<V�a<,}a<�xa<�ua<ta<Ota<)va<Yya<�}a<{�a<�a<i�a<��a<Ċa<��a<�~a<Psa<�da<�Sa<�@a<�-a<�a<Ba<��`<��`<��`<@�`<��`<�
a<Ca<=,a<b?a<�  �  vNa<�`a<�pa<|}a<��a<f�a<��a<�a<'�a<��a<ӄa<�a<~a<U|a<|a<g}a<4�a<,�a<��a<X�a<I�a<�a<v�a<1�a<p�a<@�a<nva<�fa<�Ta<�Aa<�.a<aa<�a<�a<n�`<��`<�a<�a<;a<�,a<�@a<nUa<yia<�{a<O�a<��a<U�a<��a<��a<�a<��a<�a<��a<��a<y�a<��a<e�a<��a<A�a<ߣa<ըa<��a<h�a<��a<_�a<�a<�a<��a<��a<�a<=ma<�Ya<�Fa<�5a<�'a<Qa<�a<�a<i a<V+a<m:a<.La<�_a<�sa<^�a<�a<Фa<�a<ӵa<	�a<w�a<��a<A�a<7�a<"�a<��a<!�a<�a<��a<��a<۪a<�a<#�a<��a<��a<��a<ʸa<��a<�a<�a<��a<�}a<#ja<dVa<�Ca<J3a<-&a<Ga<1a<�a<�$a<C1a<Aa<�Sa<+ga<�za<��a<'�a<��a<z�a<ڶa<Ըa</�a<o�a<��a<>�a<�a<��a<N�a<��a<J�a<��a<�a<Ьa<Ͱa<�a<$�a<�a<�a<z�a<��a<�a<��a<�qa<^a<MJa<#8a<�(a<a<�a<"a<a<�!a<}/a<@a<�Ra<Efa<ya<�a<N�a<2�a<��a<H�a<�a<�a<:�a<��a<��a<�a<m�a<�a<)�a<�a<ۖa<�a<W�a<��a<�a<��a<�a<W�a<�a<C�a<za<1ha<\Ta<�?a<�+a<�a<�
a<� a<D�`<B�`<Y a<�
a<�a<*a<'=a<DPa<{ba<�ra<�a<v�a<��a<g�a<Q�a<܏a<�a<��a<�a<a<5|a<�za<�za<�|a<�a<=�a<5�a<Ŋa<Q�a<�a<��a<��a<�}a<�qa<ba<Pa<x<a<�(a<�a<�a<s�`<��`<��`<"�`<��`<'a<5a<�&a<�:a<�  �  YMa<�_a<pa<3}a<��a<��a<K�a<��a<~�a<<�a<��a<(�a<Q�a<�~a<�~a<�a<f�a<�a<`�a<Ύa<��a<�a<�a<k�a<`�a<�a<�ua<�ea<�Sa<@a<�,a<.a<aa<�a<��`<��`<3 a<<
a<�a<�*a<?a<Ta<lha<�za<�a<a�a<T�a<ťa<[�a<V�a<U�a<h�a<g�a<��a<��a<Y�a<�a<�a<��a<��a<X�a<�a<��a<}�a<��a<�a<�a<A�a<ďa<�~a<�ka<Xa<�Da<�3a<u%a<�a<�a<�a<	a<�(a<58a<^Ja<^a<Yra<e�a<:�a<��a<�a<��a<o�a<l�a<ĸa<��a<ϱa<��a<ʪa<q�a<˧a<!�a<թa<��a<��a<��a<R�a<�a<1�a<�a<��a<تa<S�a<��a<�|a<�ha<�Ta<�Aa<1a<�#a<�a< a<�a<�"a<�.a< ?a<�Qa<�ea<vya<��a<��a<\�a<w�a<&�a<_�a<U�a<ƶa<�a<��a<�a<̧a<̥a<B�a<��a<��a<˪a<y�a<D�a<`�a<3�a<a�a<+�a<k�a<D�a<I�a<��a<�pa<i\a<vHa<�5a<O&a<�a<�a<a<�a<�a<9-a<>a<Qa<�da<xa<�a<�a<�a<��a<��a<��a< �a<��a<�a<��a<H�a<��a<��a<�a< �a<�a<ța<ٞa<�a<%�a<��a<G�a<]�a<�a<�a<2ya<1ga<
Sa<>a<�)a<�a<�a<�`<:�`<O�`<��`<2a<�a<J(a<k;a<Oa<�aa<�qa<�a<^�a<ޏa<̒a<E�a<�a<��a<1�a<�a<G�a<�~a<z}a<q}a<�~a<��a<�a<��a<!�a<��a<��a<<�a<��a<�}a<�pa<aa<�Na<�:a<�&a<�a<Da<6�`<��`<��`<m�`<@�`<�a<a<%a<-9a<�  �  vNa<�`a<�pa<|}a<��a<f�a<��a<�a<'�a<��a<ӄa<�a<~a<U|a<|a<g}a<4�a<,�a<��a<X�a<I�a<�a<v�a<1�a<p�a<@�a<nva<�fa<�Ta<�Aa<�.a<aa<�a<�a<n�`<��`<�a<�a<;a<�,a<�@a<nUa<yia<�{a<O�a<��a<U�a<��a<��a<�a<��a<�a<��a<��a<y�a<��a<e�a<��a<A�a<ߣa<ըa<��a<h�a<��a<_�a<�a<�a<��a<��a<�a<=ma<�Ya<�Fa<�5a<�'a<Qa<�a<�a<i a<V+a<m:a<.La<�_a<�sa<^�a<�a<Фa<�a<ӵa<	�a<w�a<��a<A�a<7�a<"�a<��a<!�a<�a<��a<��a<۪a<�a<#�a<��a<��a<��a<ʸa<��a<�a<�a<��a<�}a<#ja<dVa<�Ca<J3a<-&a<Ga<1a<�a<�$a<C1a<Aa<�Sa<+ga<�za<��a<'�a<��a<z�a<ڶa<Ըa</�a<o�a<��a<>�a<�a<��a<N�a<��a<J�a<��a<�a<Ьa<Ͱa<�a<$�a<�a<�a<z�a<��a<�a<��a<�qa<^a<MJa<#8a<�(a<a<�a<"a<a<�!a<}/a<@a<�Ra<Efa<ya<�a<N�a<2�a<��a<H�a<�a<�a<:�a<��a<��a<�a<m�a<�a<)�a<�a<ۖa<�a<W�a<��a<�a<��a<�a<W�a<�a<C�a<za<1ha<\Ta<�?a<�+a<�a<�
a<� a<D�`<B�`<Y a<�
a<�a<*a<'=a<DPa<{ba<�ra<�a<v�a<��a<g�a<Q�a<܏a<�a<��a<�a<a<5|a<�za<�za<�|a<�a<=�a<5�a<Ŋa<Q�a<�a<��a<��a<�}a<�qa<ba<Pa<x<a<�(a<�a<�a<s�`<��`<��`<"�`<��`<'a<5a<�&a<�:a<�  �  (Ra<�ca<�ra<o~a<��a<V�a<�a<��a<��a<�a<[a< {a<�wa<�ua<dua<�va<�ya<6~a<a�a<�a<ߍa<a�a<ʒa<\�a<��a<a�a<�xa<�ia<�Xa<�Fa<34a<�#a<�a<a<�a<�a<�	a<�a<�!a<�2a<�Ea<�Ya<�la<a~a<�a<<�a<�a< �a<[�a<�a<�a<��a<ޘa<A�a<�a<��a<��a<O�a<��a<%�a<ѣa<~�a<?�a<V�a<�a<��a<��a<�a<6�a<I�a<eqa<�^a<vLa<W<a<�.a<u%a<� a<�!a<�'a<O2a<�@a<�Qa<�da<�wa<��a<E�a<�a<`�a<�a<l�a<�a<1�a<�a<�a<=�a<5�a<��a<c�a<��a</�a<��a<Y�a<h�a<A�a<׶a<��a<��a<��a<��a<��a<W�a<7�a<�na<�[a<�Ia<:a<`-a<m%a<M"a<�$a<�+a<8a<*Ga<�Xa<�ka<F~a<��a<�a<��a<x�a<ʵa<��a<Z�a<Աa<��a<ŧa<��a<*�a<��a<ӛa<Ϝa<!�a<�a<w�a<\�a<��a<��a<;�a<�a<��a<��a<)�a<��a<�ua<�ba<�Oa<S>a<�/a<($a<�a<Ca<- a<�(a<	6a<�Ea< Xa<�ja<�|a<��a<�a<ޣa<+�a<�a<��a<ϩa<G�a<��a<��a<͔a<�a<V�a<w�a<}�a<��a<1�a<R�a<|�a<��a<c�a<��a<Ҝa<��a<��a<�|a<�ka<�Xa<�Da<|1a<e a<	a<�a<`a<Ya<ra<�a<Ba<�/a<
Ba<=Ta<�ea<�ta<��a<ωa<��a<ːa<ȏa<��a<Ňa<V�a<,}a<�xa<�ua<ta<Ota<)va<Yya<�}a<{�a<�a<i�a<��a<Ċa<��a<�~a<Psa<�da<�Sa<�@a<�-a<�a<Ba<��`<��`<��`<@�`<��`<�
a<Ca<=,a<b?a<�  �   Xa<�ga<qua<�a<��a<��a<؉a<�a<y�a<�|a<�va<jqa<*ma<�ja<Yja<�ka<�oa<�ta<#{a<�a<�a<"�a<�a<L�a<��a<(�a<�{a<�na<�^a<�Ma<=a<>-a<* a<�a<fa< a<�a<�a<�+a<�;a<�Ma<l`a<Yra<�a<_�a<-�a<|�a<6�a<ˡa<�a<��a<7�a<�a<n�a<5�a<��a<��a<_�a<�a<�a<�a<�a< �a<��a<ίa<�a<p�a<k�a<Ėa<��a<xa<�fa<�Ua<=Fa<�9a<01a<�,a<�-a<,3a<�<a<oJa<�Za<3la<�}a<n�a<��a<��a<үa<$�a<�a<ײa<��a<�a<Ңa<�a<�a<��a<S�a<��a<��a<�a<��a<��a<�a<
�a<_�a<�a<l�a<:�a<q�a<g�a<�a<�ua<�ca<�Ra</Da<�8a<;1a<\.a<�0a<j7a<WBa<�Pa<daa<�ra<@�a<ɓa<�a<�a<~�a<m�a<�a<��a<��a<��a<@�a<[�a<��a<��a<Ɛa<ɑa<ؔa<|�a<7�a<S�a<�a<?�a<��a<�a<�a<x�a<P�a<a�a<	|a<?ja<�Xa< Ha<:a<�/a<�)a<F(a<�+a<4a<@a<+Oa<�_a<Eqa<��a<d�a<a�a<Фa<��a<��a<�a<��a<̞a<�a<�a<��a<)�a<[�a<y�a<��a<��a<�a<i�a<��a<��a<��a<q�a<0�a<_�a<�a<0�a<�pa<*_a<�La<�:a<J*a<�a<ta<ba<La<a<6a<�(a<�8a<�Ia<�Za<�ja<xa<��a<C�a<�a<I�a<��a<�a<�a<8za<�sa<�na<�ja<ia<Iia<�ka<�oa<
ua<{a<ـa<��a<��a<9�a<a�a<�a<va<�ha<lYa<�Ga<;6a<9%a<ha<�
a<�a<� a<a<
a<7a<�#a<�4a<}Fa<�  �  z_a<uma<?ya<��a<D�a<��a<��a<�a<_za<�ra<Yka<�da<�_a<�\a<
\a<�]a<6ba<Cha<	pa<jxa<a�a<a�a<6�a<f�a<��a<J�a<�a<_ta<�fa<aWa<IHa<:a<�-a<'%a<s a<@ a<R$a<�,a<�8a<�Ga<8Xa<ia<ya<��a<p�a<�a<t�a<<�a<ٜa<�a<ؑa<ۊa<�a<m~a<pza<�xa<lya<�|a<��a<�a<`�a< �a<�a<q�a<��a<��a<�a<<�a<��a<�a<s�a<�pa<�aa<ZSa<�Ga<�?a<#<a<�<a<�Aa<�Ja<UWa<*fa<�ua<�a<z�a<�a<]�a<
�a<x�a<@�a<C�a<�a<��a<�a<}�a<Ȋa<��a< �a<��a<�a<(�a<��a<��a<��a<��a<ְa<��a<вa<��a<	�a<��a<-�a<�~a<�na<Z_a<�Qa<�Fa<@a<�=a<r?a<�Ea<�Oa<3]a<Dla<|a<��a<I�a<��a<��a<�a<�a<��a<��a<��a<ԛa<��a<��a<�a<��a<s�a<��a<}�a<�a<�a<כa<&�a<z�a<��a<�a<��a<��a<�a<7�a<ƃa<�sa<�ca<�Ta<�Ga<<>a<�8a<�7a<�:a<8Ba<@Ma<+[a<Cja<�ya<��a<S�a<s�a<��a<��a<�a<'�a<ݝa<�a<��a<�a<�}a<dxa<ua<0ta<�ua<�ya<�~a<��a<��a<d�a<}�a<C�a<��a<	�a<�a<�a<Iwa<�ga<�Va<�Fa<e7a<+a<"a<�a<da<�!a<!*a<�5a<Da<+Sa<�ba<�pa<}|a<\�a<~�a<b�a<��a<#�a<fa<�wa<Ooa<rga<Maa<�\a<�Za<[a<�]a<�ba<\ia<qa<�xa<<a<0�a<��a<ąa<k�a<�ya<9na<�`a<�Pa<�@a<�1a<�#a<;a<]a<a<�a<qa<�"a<G0a<�?a<�Oa<�  �  �ga<�sa<�|a<�a<��a<��a<i�a<vya<�pa<1ga<�]a<�Ua<�Oa<�Ka<�Ja<+Ma<-Ra<�Ya<�ba<ma<Cwa<q�a<��a<׋a<�a<A�a<?�a<�za<\oa<{ba<�Ta<hHa<�=a< 6a<�1a<�1a<�5a<k=a<*Ha<JUa<da<�ra<��a<�a<O�a<�a<��a<d�a<�a<�a<i�a<y~a<va<�na<ja<�ga<Oha<la<Ira<�za<Єa<N�a<|�a<G�a<��a<�a<ҫa<ާa<��a<J�a<�a<x|a<�na<bba<RXa<Qa<�Ma<8Na<�Ra<�Za<�ea<�ra<0�a<َa<K�a<��a<��a<?�a<)�a<̬a<��a<'�a<��a<�a<�a<�za<
va<�sa<�ta<�xa<a<w�a<��a<Ԛa<��a<t�a<0�a<�a<��a<r�a<��a<�a<�a<�za<#ma<3aa<�Wa<�Qa<-Oa<�Pa<�Va<�_a<1ka<�xa<��a<œa<w�a<t�a<<�a<{�a<��a<z�a<!�a< �a<�a<\�a<�}a<�va<�ra<Eqa<sa<pwa<V~a<��a<u�a<�a<��a<��a<��a<�a<��a<Ңa<֘a<t�a<�~a<ipa<*ca<�Wa<6Oa<'Ja<Ia<�Ka<�Ra<r\a<zha<va<��a<%�a<ךa<S�a<��a<2�a</�a<A�a<��a<��a</�a<5wa<xna<ha<da<ca<Bea<�ia<�pa<Pya<J�a<��a<S�a<4�a<3�a<��a<��a<*�a<�~a<qa<~ba<�Sa<lFa<r;a<W3a</a<�.a<�2a<6:a<�Da<�Pa<~^a<�ka<lwa< �a<��a<��a<�a<2�a<ta<�va<ula<\ba<Ya<[Qa<)La<�Ia<'Ja<�Ma<�Sa<�[a<
ea<�na<�wa<�~a<T�a<��a<a<}a<-ta<yha<9[a<Ma<V?a<e3a<�)a<�#a<�!a<m#a<C)a<w2a<A>a<�Ka<1Za<�  �  pa<�ya<��a<��a<��a<��a<}za<�pa<)fa<fZa<IOa<pEa<�=a<�9a<v8a<;a<�@a<�Ia<�Ta<�`a<!ma<pxa<8�a<��a<��a<:�a<��a<فa<Pxa<�ma<Yba<�Wa<�Na<Ha<�Da<eDa<�Ga<�Na<?Xa<�ca<Tpa<�|a<T�a<�a<:�a<��a<�a<.�a<)�a<��a< |a<�pa<�fa<^a<?Xa<kUa<Va<*Za<Maa<~ka<wa<̃a<�a<5�a<�a<��a<L�a<��a<�a<�a<��a<z�a<�|a<Sra<Gia<Mca<O`a<�`a<�da<�ka<�ua<��a<��a<�a<i�a<"�a<��a<�a<N�a<��a<۞a<:�a<��a<�|a<Nra<�ia<�ca<paa<�ba<
ga<�na<�xa<�a<�a<-�a<F�a<k�a<��a<7�a<�a<��a<V�a<|�a<��a<�{a<�qa<.ia<�ca<�aa<nca<3ha<pa<5za<��a<l�a<<�a<ǥa<)�a<��a<j�a<m�a<��a<��a<h�a<7�a<�wa<Wma<\ea<{`a<�^a<�`a<fa<`na<�xa<,�a<ݏa<��a<��a<q�a<~�a<��a<�a<��a<g�a<�a<�}a<�ra<�ha<"aa<�\a<�[a<C^a<�ca<�la<�va<b�a<��a<��a<J�a<@�a<f�a<D�a<��a<z�a<t�a<e�a<�sa<�ga<�]a<4Va<�Qa<�Pa<WSa<�Xa<�aa<�ka<�va<��a<?�a<��a<�a<8�a<3�a<O�a<�a<�za<na<�aa<[Va<dLa<�Ea<�Aa<�Aa<�Da<�Ja<Ta<�^a<ja<�ta<�~a<��a<��a<��a<>�a<'�a<�wa<�la<s`a<BTa<KIa<@a<:a<.7a<�7a<<a<<Ca<�La<�Wa<�ca<�na<�xa<�a<��a<��a<��a<5za<�pa<�ea<�Ya<#Na<�Ca<b;a<96a<24a<�5a<�:a<�Ba<BMa<�Xa<�da<�  �  �xa<�a<�a<o�a<�a<#}a<ta<Vha<?[a<MMa<,@a<�4a<G,a<'a<�%a<�(a<�/a<{9a<�Ea<'Ta<�ba<Qpa<U|a<u�a<d�a<��a<j�a<+�a<6�a<�xa<�oa<�fa<+_a<�Ya<�Va<�Va<�Ya<�_a<�ga<�qa<5|a<��a<ݏa<֖a<�a<��a<��a<x�a<�a<I}a<zpa< ca<)Wa<HMa<'Fa<�Ba<\Ca<�Ga<iPa<�[a<ia<�wa<f�a<��a<�a<"�a<��a<��a<��a< �a<O�a<�a<��a<΁a<Vza<Cua<�ra<sa<�va<�|a<��a<�a<�a<2�a<	�a<6�a<��a<<�a<@�a<"�a<�a<�a< |a<Lna<#ba<aXa<�Qa<�Na<Pa<1Ua<�]a<Bia<�va<لa<Z�a<��a<E�a<��a<ѱa<�a<?�a<��a<��a<��a<c�a<��a<�za<va<Gta<�ua<�ya<X�a<Ԉa<<�a<�a<��a<��a<��a<��a<խa<��a<�a<��a<|�a<va<�ha<�\a<�Sa<�Ma<-La<~Na<�Ta<^a<�ia<�wa<m�a<^�a<��a<#�a<`�a<��a<��a<��a<L�a<�a<�a<��a<ya<�ra<�na<na<Hpa<ua<1|a<�a<E�a<��a<��a<2�a<��a<a�a<�a<F�a<;�a<�a<�ta<�ea<NXa<�La<Da< ?a< >a<+Aa<Ha<�Qa<�]a<�ja<�wa<Ãa<��a<`�a<�a<��a<�a<W�a<e�a<!za<�oa<�ea<r]a<�Wa<Ta<�Sa<�Va<�[a<=ca<�ka<0ua<�}a<,�a<ɉa<��a<��a<3�a<�{a<�oa<rba<Ta<�Ea<$9a<�.a<�'a<�$a<b%a<8*a<�2a<�=a<�Ja<�Xa<�ea<�qa<h{a<��a<��a<��a<�a<�xa<pa<0fa<�\a<�Sa<�La<SHa<�Fa<Ha<`La<)Sa<�[a<�ea<toa<�  �  �a<��a<�a<�a<]�a<Iya<�ma<`a<�Pa<�@a<2a<-%a<ka<�a<Xa<Ka<�a<*a<J8a<Ha<�Xa<�ha<}va<1�a<'�a<Ďa<��a<��a<�a<��a<�{a<`ta<bna<�ia<�ga<�ga<~ja<�oa<8va<�~a<E�a<f�a<j�a</�a<�a<^�a<l�a<��a<��a<9ta<ea<LVa<pHa<=a<
5a<F1a<�1a<�6a<@a<�La<\a<Qla<}a<��a<
�a<��a<c�a<�a<��a<m�a<إa<��a<Z�a<�a<�a<��a<��a<)�a<�a<�a<p�a<Q�a</�a<?�a<̮a<�a<رa</�a<?�a<�a<Z�a<�a<1pa<�`a<�Ra<�Ga<F@a<E=a<�>a<?Da<Na<�Za<ja<�ya<ˉa<
�a<�a<�a<��a<ʳa<�a<��a<�a<|�a<��a<H�a<��a<ֆa<t�a<k�a<�a<.�a<$�a<�a<i�a<��a<��a<��a<�a<-�a<��a<͗a<��a<�ya<�ia<qZa<Ma<�Ba<w<a<�:a<=a<Da<�Na<G\a<nka<4{a<��a<ؗa<ܢa< �a<�a<l�a<��a<�a<�a<,�a<#�a<S�a<�a<�a<2a<׀a<�a<��a<őa<W�a<H�a<�a<��a<$�a<	�a<��a<}�a<Q�a<
za<Tia<Ya<�Ia<�<a< 3a<�-a<�,a<�/a<�7a<�Ba<�Pa<J_a<�na<�|a<��a<��a<L�a<��a<�a<��a<�a<��a<V|a<�sa<7ma<�ga<,ea<�da<�fa<'ka<�pa<=xa<~a<��a<��a<��a<��a<��a<5�a<�ua<Hha<�Xa<"Ha<V8a<�)a<aa<pa<
a<�a<Ja<�"a<_/a<">a<�Ma<a]a<cka<=wa<�a<��a<c�a<u�a<�a<Cya<�qa<�ia<lba<�\a<Ya<�Wa<�Xa<}\a<�aa<*ia<5qa<�xa<�  �  ݅a<�a<K�a<3�a<�a<`ua<-ha<�Xa<SGa<�5a<�%a<�a<a<�a<a<�a<�a<�a<	,a<�=a<�Oa<�aa<Gqa<�~a<�a<}�a<��a<S�a<��a<�a<��a<&�a<J{a<�wa<�ua<5va<xxa<�|a<��a<^�a<p�a<Жa<�a<��a<��a<�a<�a<7�a<�{a<&la<G[a<�Ja<;a<#/a<}&a<)"a<�"a</(a<2a<�?a<TPa<Uba<�ta<9�a<d�a<�a<תa<7�a<��a<��a<�a<�a<��a<+�a<@�a<��a<�a<g�a<��a<�a<\�a<��a<ƪa<��a<��a<δa<Ʋa<)�a<
�a<w�a<��a<dwa<�ea<�Ta<�Ea<�9a<�1a< .a<|/a<�5a<?@a<@Na<�^a<{pa<'�a<J�a< �a<ߪa<�a<ӵa<�a<p�a<ծa<�a<Ţa<�a<�a<�a<ɓa<��a<[�a<�a<��a<��a<l�a<	�a<ȴa<Ҵa<a�a<c�a<Пa<9�a<>�a<�pa<�^a<�Ma<f?a<k4a<�-a<^+a<D.a<�5a<9Aa<Pa<�`a<Yra<��a<��a<d�a<٨a<��a<�a<$�a<��a<r�a<D�a<�a<<�a<��a<(�a<��a<юa<%�a<�a<��a<��a<��a<��a<�a<��a<��a</�a<�a<)�a<�qa<�_a<�Ma<�<a<�.a<s$a<�a<ya<[!a<�)a<�5a<�Da<NUa<Afa<Ava<�a<*�a<��a<՚a<`�a<�a<$�a<�a<�a<.�a<Xza<�ua<ysa<sa<�ta<xa<�|a<��a<�a<��a<ɏa<d�a<ύa<��a<~a<�pa<uaa<�Oa<�=a<C,a<�a<)a<�a<�a<�a<�
a<�a<�"a<3a<RDa<�Ua<�ea<"sa<�}a<ބa<j�a<v�a<ąa<�a<;{a<�ta<oa<?ja<$ga<fa<ga<�ia<�na<�ta<�za<�a<�  �  f�a<�a<��a<�a<~a<lra<�ca<�Ra<%@a<j-a<�a<3a<�a<��`<��`<��`<Ka<�a<�"a<J5a<�Ha<�[a<Rma<	|a<��a<��a</�a<��a<i�a<j�a<8�a<�a<��a<S�a<�a<?�a<{�a<�a<֋a<o�a<@�a<Y�a<��a<�a<��a<�a<ԑa<څa<�va<�ea<�Sa<�Aa<�1a<k$a<�a</a<�a<ya<1'a<�5a<Ga<�Za<.na<�a<�a<��a<#�a<�a<4�a<��a<i�a<��a<��a<U�a<;�a<��a<�a<e�a<{�a<��a<<�a<E�a<0�a<��a<�a<��a<$�a< �a<x�a<��a<��a<�pa<�]a<_Ka<�;a<l.a<�%a<�!a<�#a<9*a<�5a<�Da<Va<.ia<�{a<��a<�a<1�a<�a<��a<иa<ȷa<��a<*�a<�a<[�a<r�a<��a<՞a<��a<աa<q�a< �a<�a<p�a<��a<Ʒa<�a<K�a<�a<ܜa<ލa<1|a<]ia<2Va<LDa<5a<�(a<�!a<Oa<x"a<x*a<7a<�Fa<�Xa<hka<�}a<��a<��a<��a<�a<��a<t�a<|�a<��a<Ũa<��a<�a<n�a<+�a<��a<֙a<>�a<'�a<��a<V�a<>�a<��a<~�a<��a<,�a<�a<��a<,~a<}ka<
Xa<fDa<�2a<�#a<�a<�a<wa<�a<�a<�+a<�;a<�Ma<�_a<qa<��a<�a<
�a<��a<��a<��a<{�a<��a<�a<W�a<R�a<ـa<z~a<	~a<da<�a<ʅa<1�a<��a<��a<D�a<5�a<.�a<��a<r{a<%ma<�[a<	Ia<�5a<�"a<�a<a<��`<��`<�`<H�`<}
a<a<<*a<=a<�Oa<aa<pa<|a<��a<��a<@�a<�a<�a<S�a<5}a<yxa<�ta<(ra<!qa<ra<kta<8xa< }a</�a<��a<�  �  .�a<��a<��a<�a<}a<vpa<�`a<�Na<~;a<(a<�a<aa<e�`<��`<��`<��`<�`<�a<�a<0a<MDa<6Xa<�ja<Oza<�a<�a<j�a<��a<\�a<.�a< �a<v�a<+�a<Èa<��a<�a<�a<9�a<��a<��a<��a<��a<\�a<��a<4�a<�a<��a<��a<�sa<�aa<�Na<<a<g+a<ha<�a<a<�a<Xa< a<f/a<oAa<�Ua<ja<�}a<l�a<H�a<��a<��a<��a<�a<��a<ɲa<	�a<�a<��a<�a<£a<�a<�a<�a<�a<%�a<�a<�a<H�a<�a<x�a<i�a<ןa<��a<~a<Ela<�Xa<�Ea<�4a<H'a<�a<�a<�a<#a<�.a<t>a<�Pa<pda< xa<��a<ؚa<�a<��a<ڷa<��a<w�a<(�a<��a<v�a<\�a<רa<u�a<��a<(�a<?�a<��a<q�a<��a<��a<]�a<��a<�a<;�a<�a<�a<�a<sxa<�da<�Pa<4>a<:.a<�!a<�a<3a<Ra<I#a<l0a<�@a<eSa<�fa<8za<ދa<��a<צa<)�a<�a<z�a<n�a<��a<��a<9�a<�a<ݡa<̟a<;�a<@�a<��a<��a<ީa<��a<��a<�a<�a<A�a<ǥa<ښa<U�a<�za<xga<Sa<�>a<�,a<�a<�a<ta<]
a<�a<�a<m%a<�5a<�Ha<�[a<�ma<~a<��a<��a<!�a<�a<"�a<��a<Ƙa<�a<�a<��a<=�a<+�a<��a<υa<!�a<q�a<�a<d�a<��a<o�a<��a<��a<�a<�ya<rja<rXa<�Da<�0a<a<�a<��`<��`<��`<��`< �`<�a<�a<�$a<H8a<�Ka<�]a<�ma<{a<t�a<n�a<��a<Ɍa<a�a<Άa<��a<x~a<�za<�xa<�wa<�xa<�za<K~a<p�a<��a<��a<�  �  l�a<��a<v�a<��a<��a<�sa<^a<Fa<k+a<�a<��`<��`<2�`<Z�`<��`<��`<��`<�`<, a<la<�5a<Qa<�ia<�~a<X�a<@�a<��a<ϥa<��a<'�a<,�a<ƚa<��a<�a<�a<Y�a<C�a<�a<�a<��a<I�a<�a<�a<��a<ݬa<E�a<U�a<c�a<�oa<Wa<�<a<F#a<�a<��`<��`<��`<T�`<a�`<�`<_a<*(a<1Ca<_a<�ya<8�a</�a<!�a<��a<O�a<%�a<��a<r�a<ݼa<)�a<�a<&�a<��a<0�a<�a<f�a<Թa<�a<��a<��a<�a<��a<��a<�a<n�a<8�a<�ya<T_a<PDa<q*a<ja<a<��`<S�`<��`<�`<)a<Y a<z9a<4Ta<Loa<[�a<B�a<��a<ϼa<G�a<�a<r�a<��a<��a<��a<�a<�a<g�a<|�a< �a<H�a< �a<��a<t�a<��a<T�a<(�a<��a<��a<%�a<ܞa<1�a<\pa<GUa<S:a<� a<�
a</�`<��`<��`<0�`<��`<Ca<�$a<S>a<*Ya<�sa<f�a<��a<گa<�a<��a</�a<Q�a<�a<T�a<(�a<��a<٭a<իa<S�a<K�a<��a<�a<n�a<�a<��a<'�a<��a<r�a<p�a<�a<��a<zwa<-]a<[Aa<.&a<a<A�`<��`<.�`<��`<^�`<]�`<a<Ia<�5a<Pa<7ia<?a<ʑa<]�a<��a<��a<��a<�a<��a<�a<[�a<c�a<��a<��a<�a<�a<ݓa<��a<#�a<C�a<�a<��a<�a<�a<a<�~a<ja<Ra<'7a<�a<La<��`<�`<b�`<q�`<T�`<|�`<2�`<�`<�a<Y'a<-Ba<�Za<�pa<-�a<Ўa<�a<a<��a<U�a<	�a<�a<?�a<D�a<Ƀa<��a<��a<�a<��a<̎a<�a<r�a<�  �  1�a<��a<L�a<�a<3�a<�ta<�_a<�Ga<�-a<ra<��`<��`<y�`<��`<b�`<W�`<�`<2�`<�a<�a<�7a<vRa<�ja<�a<Џa<q�a<e�a<�a<^�a<r�a<.�a<��a<9�a<1�a<��a<ӏa<7�a<�a<T�a<Z�a<k�a<��a<�a<B�a<Ҭa<��a<��a<��a<!qa<�Xa<B?a<�%a<�a<��`<H�`<��`<�`<��`<0�`<la<�*a<�Ea<�`a<{a<b�a<ۥa<��a<��a<��a<4�a<X�a<��a<��a<��a<;�a<,�a<w�a<ˬa<�a<��a<��a<ۼa<��a<��a<I�a<��a<ӿa<T�a<!�a<i�a<{a<Saa<�Fa<5-a<�a<Ta<P�`<�`<A�`<k�`<Ia<@#a<<a<�Va<�pa<��a<-�a<��a</�a<*�a<��a<J�a<U�a<��a<r�a<E�a<��a<;�a<�a<ܮa<X�a<Q�a<M�a<��a<�a<�a<��a<��a<�a<��a<��a<u�a<�qa<�Wa<�<a<�#a<a<x�`<o�`<Q�`<��`<��`<`a<�'a<�@a<=[a<	ua<��a<��a<R�a<?�a<}�a<s�a<�a<\�a<V�a<�a<ήa<�a<z�a<ͧa<>�a<�a<O�a<;�a<%�a<
�a<%�a<3�a<f�a<�a<��a<��a<�xa<�^a<�Ca<�(a<a<g�`<>�`<��`<��`<��`<��`<%a<�a<98a<�Qa<�ja<j�a<v�a<Пa<��a<��a<��a<��a<Ȥa<ٞa<ؘa<��a<��a<�a<��a<-�a<�a<S�a<�a<��a<��a<Ƣa<��a<;�a<4�a<za<>ka<fSa<$9a<4a<a<��`<E�`<��`<+�`<��`<��`<R�`<��`<|a<�)a<�Ca<D\a<�qa<��a<0�a<��a<9�a<ՙa<Ɩa<%�a<Ìa<��a<S�a<��a<na<y�a<!�a<N�a<��a<�a<זa<�  �  ��a<��a<%�a<a�a<Ɇa<xwa<�ca<�La<�3a<�a<�a<��`<%�`<��`<U�`<+�`<��`<!�`<�
a<$a<�=a<[Wa<�na<�a<)�a<q�a<��a<}�a<��a<q�a<ݖa<?�a<�a<��a<��a<݆a<o�a<��a<��a<��a<ءa<F�a<ͬa<V�a<�a<|�a<��a<߉a<�ua<E^a<�Ea<{-a<ea<a<�`<��`<��`<~�`<�a<a<u2a<tLa<�fa<�a<ޕa<��a<��a<�a<�a<?�a<@�a<"�a<�a<�a<ڨa<j�a<��a<�a<^�a<r�a<.�a<i�a<��a<��a<��a<�a<��a<��a<��a</�a<�a<8ga<�Ma<5a<da<�a<!a<��`<%�`<%a<xa<�+a<hCa<�\a<va<�a<3�a<>�a<��a<&�a<_�a<��a<��a<�a<y�a<n�a<��a<c�a<��a<��a<ͨa<d�a<9�a<~�a<a�a<��a<G�a<]�a<=�a<E�a<��a<��a<wa<�]a<Da<�+a<4a<%a<U�`<G�`<��`<g	a<Qa<�/a<�Ga<@aa<�ya<��a<I�a<��a<@�a<�a<��a<S�a<[�a<�a<��a<��a<Q�a<��a<מa<u�a<��a<��a<|�a<��a<ʹa<�a<G�a<��a<��a<��a<�a<E}a<cda<oJa<b0a<�a<�a<�`<��`<��`<{�`<��`<�a<�&a< ?a<�Wa<oa<�a<��a<��a<��a<ªa<��a<��a<U�a<3�a<P�a<#�a<׆a<"�a<��a<��a<�a<�a<��a<Y�a<�a<�a<	�a<�a<k�a<�a<oa<*Xa<?a<5%a<�a<��`<��`<��`<�`<��`<��`<��`<T�`<�a<0a<�Ha<�`a<�ta<r�a<��a<��a<�a<}�a<=�a<G�a<ͅa<�a<�za<�wa<uva<�wa<�za<ca<t�a<��a<+�a<�  �  �a<�a<��a<��a<�a<�{a<�ia<�Ta<�=a<4&a<a<��`<s�`<��`<��`<��`<��`<a<�a<"/a<]Ga<_a<ta<��a<�a<E�a<��a<c�a<��a<;�a<�a<��a<Ia<bza<�wa<.xa<�za<6�a<��a<�a<Әa< �a<ȧa<o�a</�a<]�a<Ҝa<i�a<7|a<ga<Pa<�9a<�$a<�a<�a<�a<a<1	a<Ka<�(a<�>a<�Va<loa<��a<��a<�a<��a<O�a<p�a<l�a<P�a<O�a<��a<�a<��a<זa<єa<*�a<�a<u�a<m�a<L�a<Q�a<f�a<A�a<��a<H�a<�a<�a<\�a<M�a<upa<�Xa<�Aa<7-a<�a<�a<=a<a<�a<�%a<�8a< Oa<�fa<n~a<��a<n�a<��a<�a<��a<��a<|�a<2�a<y�a<n�a<��a<ța<��a<B�a<A�a<�a<͠a<�a<�a<��a<�a<��a<��a<u�a<~�a<��a<y�a<a<}ga<�Oa<9a<d%a<va<@a<�
a<]a<�a<F(a<N<a<Sa<�ja<��a<�a<�a<m�a<�a<�a<Ƽa<+�a<&�a<�a<
�a<ݙa<!�a<ڐa<'�a<Αa<;�a<y�a<Уa<��a<��a<�a<^�a<��a<��a<��a<��a<�a<ma<�Ta<�<a<&a<Na<�a<��`<��`<-a<�a<fa<�2a<gIa<n`a<va<��a<��a<١a<;�a<�a<ߤa<��a<��a<��a<G�a<�}a<Exa<pua<ua<)wa<�{a<A�a<��a<�a<q�a<��a<Ҝa<��a<�a<\�a<,ta<�_a<AHa<0a<�a<�a<��`<l�`<V�`<��`<��`<��`<�a<�"a<�9a<OQa<�fa<�xa<�a<�a<��a<��a<�a<��a<܂a<�za<Ksa<"ma<ia<�ga<�ha<�la<�ra<Aza<c�a<`�a<�  �  D�a<��a<�a<��a<��a<a<Yqa<�^a<Ja<�4a<� a<Xa<$a<�`< �`<#�`<8a<.a<(a<G=a<CSa<�ha<{a<n�a<�a<��a<��a<��a<-�a<g�a<�a<%va<na<ha<�da<�da<ha<�na<wa<��a<��a<��a<Πa<��a<k�a<0�a<X�a<t�a<��a<�qa<C]a<Ia<86a<�&a<�a<a<�a<"a<^)a<5:a<mNa<;da<�za<2�a<�a<֮a<��a<ֻa<?�a<��a</�a<��a<��a<ڑa<
�a<:�a<��a<��a<��a<"�a<��a<�a<:�a<ɲa<(�a<S�a<f�a<ιa<w�a<5�a<��a<|a<�fa<�Qa<&?a<80a<&a<�!a<�#a<W+a<g8a<�Ia<^a<psa<��a<כa<�a<��a<S�a<o�a<�a<��a<1�a<�a<��a<,�a<̉a<��a<��a<;�a<Ԉa<׏a<��a<;�a<H�a<&�a<M�a<!�a<n�a<�a<ܫa<�a<(�a<�sa<O^a<�Ia<�7a<,*a<�!a<a<�"a<,a<g:a<�La<;aa<�va<!�a<�a<��a<r�a<x�a<׺a<��a<ׯa<S�a<��a<��a<��a<΁a<�}a<�|a<a<��a<�a<��a<��a<8�a<�a<�a<��a<W�a<�a<��a<G�a<�wa<�aa<�Ka<{7a<8&a<�a<ca<>a<a<� a<�/a<�Ba<�Va<�ka<�~a<�a<u�a<��a<ĥa<�a<1�a<~�a<�a<�a<ua<Vla<�ea<.ba<�aa<�da<�ja<{ra<|a<؅a<Ԏa<��a<A�a<ɘa<��a<ɉa<{a<�ha<�Sa<�=a<�(a<�a<a<}�`<��`<@�`<��`<ia<�a<s1a<�Fa<�[a<zna<U~a<ԉa<Y�a<I�a<��a<��a<��a<{va<la<�ba<+[a<#Va<�Ta<�Ua<�Za<�aa<;ka<�ua<�a<�  �  �a<Z�a<r�a<@�a<�a<��a<�ya<ja<GXa<{Ea<�3a<m$a<�a<�a<�a<�a<�a<�)a<�:a<fMa<�`a<�ra<��a<�a<��a<��a<��a<z�a<�a<U|a<�oa<�ca<�Ya<BRa<3Na<Na<�Qa<YYa<�ca<�pa<�~a<a�a<K�a<��a<�a<ϧa<~�a<ߚa<��a<�}a<{la<[Za<�Ia<N<a<�2a<�-a<[.a<V4a<??a<*Na<`a<�sa<�a<ɘa<��a<L�a<��a<ɹa<�a<��a<'�a<��a<ߊa<�~a<�ta<$na<�ja<Bka<�oa<zwa<F�a<��a<Λa<U�a<��a<۹a<�a<V�a<��a<��a<��a<T�a<�va<da<�Sa<hFa<w=a<�9a<B;a<#Ba<�Ma<]a<�na<�a<;�a<��a<��a</�a<N�a<G�a<ҷa<��a<$�a<�a<3�a<�}a<Tta<Tna<la<�ma<5sa<�{a<G�a<�a<�a<��a<�a<��a<�a<f�a<�a<��a<R�a<,�a<�na<�\a<�La<�@a<J9a<�6a<:a<eBa<Oa<%_a<_qa<(�a<��a<�a<3�a<C�a<�a<��a<�a<��a<A�a<�a<_a<=ta<�ka<ga<�ea<�ha<Zoa<�xa<��a<9�a<ߝa<��a<p�a<��a<��a</�a<�a<��a<�a<�pa<@]a<2Ka<�;a<�0a< *a<�(a<S-a<�6a<�Ca<,Ta<Bfa<xa<L�a<a<�a<�a<��a<ʞa<�a<x�a<�|a<oa<4ba<LWa<�Oa<YKa<"Ka<�Na<�Ua<`a<�ka<lxa<_�a<6�a<Ɣa<w�a<-�a<�a<��a<�ra<aa<�Ma<�:a<�)a<Ka<�a<�a<�a<wa<�!a<�0a<MBa<-Ua<ga<Iwa<�a<f�a<V�a<$�a<��a<T�a<�ta<rga<�Za<�Na<�Ea<�?a<�=a<q?a<Ea<�Ma<�Ya<lfa<�sa<�  �  �ta<��a<��a<
�a<�a<1�a<E�a<lua<�fa<�Va<Ha<�:a<z0a<�*a<)a<a,a<�3a<�?a<2Na<6^a<�na<�}a<��a<m�a<&�a<��a<u�a<5�a<[|a<�ma<a^a<Pa<�Ca<j:a<�5a<;5a<�9a<RBa<Oa<(^a<�na<ma<t�a<#�a<��a<§a<��a<�a<j�a<|�a<�{a<�la<_a<Sa<�Ja<�Fa<sGa<�La<$Va<{ca<�ra<��a<ݓa<��a<S�a<̵a<�a<��a<�a<�a<z�a<�a<�xa<Rja<,^a<�Ua<�Qa<�Ra<�Wa<aa<$na<�|a<�a<Z�a<�a<s�a<��a<g�a<θa< �a<&�a<�a<�a<xwa<\ia<�]a<!Va<�Ra<6Ta<
Za<%da<�qa<��a<��a<�a<g�a<�a<��a<|�a<�a<��a<"�a<��a<��a<va<ha<�\a<�Ua<(Sa<MUa<�[a<@fa<�sa<�a<�a<��a<j�a<-�a<�a<��a<M�a<��a<��a<��a<m�a<qa<;ca<�Xa<2Ra<Pa<�Ra<�Ya<ea<�ra<6�a<�a<e�a<��a<��a<��a<��a<��a<��a<�a<֊a<�za<}ka<^a<%Ta<tNa<.Ma<�Pa<PXa<da< ra<h�a<�a<��a<�a<�a<�a<Y�a<P�a<�a<��a<�a<�oa<G`a<�Ra<�Ha<)Ca<Ba<�Ea<~Ma<7Ya<�fa<va<�a<�a<a�a<n�a<3�a<��a<��a<��a<�}a<Uma<�\a<�Ma<}@a<r7a<�2a<w2a<�6a<�?a<�Ka<"Za<�ia<bxa<��a<\�a<�a<;�a<�a<�a<f}a<�na<P^a<>Na<�?a<�3a<�+a<�'a<�(a<Z.a< 8a<KEa<Ta<da<�ra<	�a<|�a<�a<��a<��a<q�a<�ua<ga<�Va<mGa<|9a<P.a<h'a<�$a<'a<|-a<Q8a<-Fa<�Ua<�ea<�  �  �ia<�ya<��a<	�a<~�a<ԏa<�a<��a<�ta<�ga<�[a<uPa<Ha<Ca<�Aa<�Da<CKa<Ua<8aa<�na<#|a< �a<��a<k�a<Øa<��a<��a<I�a<ipa<�^a<lLa<p;a<-a<r"a<�a<a<!a<)+a<k9a<�Ja<g^a<�qa<6�a<��a<��a<�a<C�a<��a<E�a<��a<�a<�~a<Gsa<�ia<�ba<�_a<4`a<�da<�la<xa<�a<˒a<^�a<Ϋa<4�a<��a<n�a<��a<?�a<1�a<h�a<xa<�ea<�Ta<-Ga<�=a<�8a<�9a<�?a<oJa<2Ya<�ja<�}a<�a<Ѡa<f�a<��a<��a<{�a<��a<0�a<�a<�a<=�a<o~a<�ta<gna<�ka<�la<�qa<2za<b�a<�a<;�a<}�a<x�a<�a<y�a<ٻa<s�a<̨a<6�a<��a<�ta<.ba<Ra<eEa<'=a<�9a<m<a<�Ca<Pa<�_a<�qa<��a<c�a<*�a<&�a<�a<��a<�a<��a<�a<��a<k�a<��a<ya<7pa<�ja<�ha<5ka<+qa<]za<�a<��a<�a<Ϊa<��a<��a<X�a<ܴa<�a<��a<�a<�{a<�ha<�Va<�Ga<,<a<|5a<4a<8a<%Aa<ZNa<�^a<qa<x�a<l�a<ݢa<�a<�a<�a<߯a<�a<��a<i�a<��a<�ta<!ia<�`a<�[a<�Za<�]a<2da<�ma<%ya<\�a<d�a<T�a<C�a<e�a<��a<�a<�a<��a<�pa<[]a<�Ia<8a<�)a<�a<ua<ta<�a<�(a<7a<�Ga<PZa<la<G|a<M�a<�a<w�a<Õa<s�a<l�a<�{a<Nna<�`a<�Ta<�Ja<�Ca<�@a<oAa<!Fa<)Na<Ya<fea<Wra<[~a<�a<o�a<��a<�a<W�a<�za<�ja<	Ya<�Ea<�3a<{#a<�a<�a<�a<(a<�a<'"a<	2a<IDa<}Wa<�  �  �^a<Hqa<�a<܋a<��a<y�a<��a<?�a<_�a<jwa<Qma<zda<�]a<�Ya<�Xa<[a<�`a<�ha<�ra<n}a< �a<*�a<{�a<a�a<��a<H�a<�a<Uwa<�da<Pa<t;a<(a<�a<�a<�a<Ta<�	a<a<%a<�8a<�Na<�da<:za<��a<��a<��a<êa<S�a<ۧa<=�a<��a<�a<Ņa<H~a<�xa<Kva< wa<�za<ˁa<��a<��a<��a<>�a<��a<)�a<��a<^�a<Q�a<>�a<x�a<�}a<�ha<�Sa<�@a<51a<=&a<	!a<�!a<�(a<�4a<�Ea<mYa<�na<�a<��a<0�a<��a<2�a<�a<N�a<�a<��a<��a<Y�a<��a<�a<��a<��a<f�a<��a<~�a<o�a<ԡa<!�a<��a<d�a<��a<H�a<�a<��a<��a<��a<�ya<?da<�Oa<K=a<�.a<�%a<3"a<�$a<f-a<;a<�La<6aa<�va<a�a<̝a<�a<��a<v�a<��a<;�a<��a<N�a<�a<a�a<�a<�a<5�a<�a<��a<��a<؍a<;�a<z�a<a�a<ݳa<}�a<��a<7�a<)�a<�a<a<u�a<ma<�Wa<wCa<+2a<O%a<�a<Ca<� a<+a<:a<�La<Eaa<qva<m�a<��a<�a<��a<n�a<��a<��a<S�a<�a<��a<�a<�}a<�va<�ra<�qa<�sa<&ya<{�a<��a<Q�a<E�a<D�a<9�a<A�a<��a<G�a<�a<�xa<da<�Ma<8a<$a<�a<�a<�a<�a<�a<Qa<n#a<�6a<>Ka<`a<sa<�a<�a<��a<\�a<�a<�a<I�a<�|a<ra<�ga<�_a<Za<�Wa<Xa<�[a<rba<ka<2ua<<a<]�a<�a<m�a<��a<��a<��a<�ra<0`a<DKa<�5a<
!a<�a<o a<�`<��`<��`<P�`<,a<4a<�3a<_Ia<�  �  �Ta<�ia<�{a<i�a<(�a<A�a<�a<*�a<ˋa<)�a<w|a<ua<�oa<�la<la<�ma<�ra<3ya<&�a<��a<֑a<��a<d�a<��a<4�a<3�a<M�a<Zoa<PZa<RCa<j,a<�a<�a<��`<y�`<��`<��`<�a<Ka<�(a<�@a<|Ya<qa<�a<A�a<�a<ʫa<�a<�a<��a<��a<��a<��a<��a<@�a<��a<A�a<f�a<H�a<ۚa<f�a<6�a<9�a<D�a<2�a<�a<�a<S�a<Ǜa<��a<~ra<�Za<Da<%/a<a<Aa<{a<La<�a<�!a<M4a<"Ja<�aa<_ya<Z�a<J�a<X�a<��a<�a<��a<�a<%�a<��a<��a<2�a<ܛa<k�a<ȕa<��a<�a<��a<֦a<Ӯa<Ӷa<��a<�a<�a<ÿa<��a<�a<��a<�a<�ma<�Ua<?a<+a<ha<Ra<�a<ra<�a<�(a<3<a<�Ra<:ja<v�a<Z�a<��a<@�a<��a<^�a<��a<��a<��a<��a<��a<�a<�a<C�a<&�a<o�a<|�a<��a<ݥa<��a<<�a<E�a<j�a<�a<иa<�a<x�a<ɍa<xa<A`a<�Ha<]2a<ya<�a<Q	a<�a<�a<�a<5(a<�<a<�Sa<�ja<P�a<˔a<Ǥa<�a<t�a<;�a<��a<�a<8�a<x�a<�a<F�a<4�a<υa<�a<d�a<��a<��a<��a<Ȟa<A�a<̩a<C�a<��a<[�a<J�a<|�a<#pa<�Xa<B@a<B(a<ga<d a<��`<&�`<3�`<��`<y a<$a<X'a<9>a<dUa<�ja<-}a<��a<P�a<G�a<��a<<�a<֐a<�a<j�a<rxa<�qa<�la<�ja<"ka<(na<�sa<zza</�a<�a<��a<��a<��a< �a<Ήa<�|a<Ska<�Va<>?a<t'a<�a<��`<��`<��`<C�`<7�`<��`<��`<�a<D%a<=a<�  �  �La<da<�wa<O�a<�a<�a<��a<��a<��a<܍a<��a<�a<�}a<Y{a<�za<�|a<)�a<��a<�a< �a<N�a<��a<��a<ҝa<��a<��a< }a<ia<�Qa<b9a<� a<�	a<��`<S�`<|�`<��`<��`<��`<�a<Ra<6a<UPa<�ia<ڀa<�a<��a<C�a<b�a<��a<��a<@�a<˦a<{�a<��a<��a<<�a<��a<�a<x�a<Цa<ǭa<�a<
�a<��a<��a<��a<޴a<(�a<�a<��a<~ia<}Pa<�7a<}!a<:a<�a<Y�`<D�`<#a<va<�&a<>a<�Wa<�pa<܈a<֝a<��a<ºa<�a<��a<(�a<j�a<Ӻa<z�a<w�a<Y�a<�a<{�a<@�a<��a<i�a<T�a<��a<�a<��a<�a<��a<׿a<�a<#�a<�a<!}a<8da<�Ja<A2a<a<6a<{a<[�`<� a<t
a<�a<1/a<;Ga<�`a<}ya<��a<�a<%�a<��a<�a<r�a<N�a<��a<c�a<ذa<��a< �a<��a<ܡa<)�a<!�a<�a<Ӱa<�a<��a<��a<��a<'�a<C�a<��a<,�a<��a<�oa<RVa<�<a<%a<a<
a<S�`<|�`<��`<�a<qa< 0a<�Ha<�aa<�ya<��a<i�a<��a<�a<��a<7�a<��a<��a<��a<��a<S�a<��a<��a<��a<�a<ӗa<��a<�a<��a<�a<��a<ϭa<:�a<(�a<!�a<�a<ia<�Oa<�5a<�a<�a<��`<�`<�`<,�`<R�`<��`<�a<Ta<4a<�La<Nda<�xa<�a<��a<K�a<��a<Y�a<�a<�a<.�a<��a<%a<|{a<uya<�ya<A|a<X�a<��a<�a<�a<��a<��a<m�a<�a<��a<ya<�ea<�Na<�5a<@a<�a<��`<��`<
�`<�`<V�`<f�`<��`<�a<�a<�3a<�  �  �Ga<`a<
ua<Ʌa<ёa<,�a<�a<|�a<r�a<��a<��a<�a<h�a<<�a<��a<m�a<��a<^�a<��a<ɘa<ŝa<'�a<ˡa<a<�a<݊a<�ya<�da<�La<�2a<3a<Na<U�`<��`<��`<��`<�`<^�`<��`<�a<)/a<�Ja<ea<(}a<��a<f�a<��a<��a<T�a<m�a<{�a<K�a<٨a<��a<]�a<%�a<�a<��a<Ϩa<H�a<`�a<O�a<�a<��a<r�a<	�a<ܳa<��a<a�a<�|a<�ca<�Ia<�/a<�a<�a<��`<n�`<^�`<a�`<-
a<fa<�6a<�Pa<Nka<s�a<��a<��a<�a<��a<��a<Q�a<��a<x�a<H�a<)�a<ɱa<�a<t�a<(�a<��a<|�a<��a<��a<��a<`�a<��a<X�a<��a<x�a<y�a<�a<(xa<"^a<�Ca<.*a<a<�a<��`<f�`<��`<� a<ya<�&a<@a<cZa<ita<��a<6�a<��a<M�a<K�a<��a<��a<f�a<�a<��a<��a<��a<�a<תa<��a<��a<��a<��a<�a<1�a<��a<��a<�a<��a<Ūa<�a<?�a<Eja<�Oa<^5a<�a<�a<L�`<p�`<��`<�`<S�`<�a<P(a<�Aa<�[a<Gua<�a<�a<��a<2�a<"�a<��a<��a<��a<+�a<�a<��a<P�a<p�a<��a<��a<*�a<�a<��a<�a<�a<c�a<��a<��a<'�a<�a<|a<|da<$Ja<�.a<+a<�`<.�`<9�`<�`<G�`<��`<��`<=�`<�a<�-a<RGa<�_a<pua<�a<ٓa<�a<��a<�a<j�a<��a<��a<d�a<��a<D�a<l�a<��a<ۄa<j�a<.�a<O�a<��a<;�a<6�a<ǘa<��a<��a<eva<�aa<�Ia<�/a<!a<��`<��`<&�`<2�`<�`<u�`<��`<��`<Z�`<�a<G-a<�  �  Fa<�^a<7ta<C�a<��a<X�a<��a<��a<�a<�a<(�a<̌a<U�a<��a<A�a<��a<��a<�a<<�a<��a<Q�a<E�a<K�a<ٞa<��a<I�a<�xa<�ca<�Ja<�0a<�a<_�`<2�`<D�`<��`<��`<��`<(�`<��`<�a<�,a<�Ha<�ca<�{a<ߐa<��a<y�a<W�a</�a<Ƶa<B�a<f�a<9�a<��a<A�a<��a<Z�a<��a<��a<��a<��a<$�a<t�a<��a<��a<�a<i�a<K�a<5�a<�{a<�aa<Ga<B-a<�a<�a<`�`<��`<��`<�`<a<ga<�3a<�Na<�ia<"�a<{�a<�a<��a<��a<n�a<[�a<D�a<Y�a<~�a<Ÿa<��a<��a<��a<~�a<��a<8�a<ջa<��a<��a<��a<E�a<��a<��a<��a<��a<юa<�va<
\a<Aa<`'a<�a<j�`<�`<��`<�`<��`<\a<$$a<~=a<5Xa<�ra<>�a<d�a<�a<��a<w�a<m�a<�a<	�a<q�a<A�a<o�a<~�a<-�a<`�a<�a<��a<c�a<��a<¾a<��a<�a<X�a<0�a<]�a<1�a<�a<��a<�ha<�Ma<�2a<�a<�a<��`<��`<��`<��`<�`<�a<�%a<??a<�Ya<�sa<يa<b�a<�a< �a<��a<ҽa<ٻa<��a<F�a<x�a<[�a<4�a<ؠa<��a<��a<�a<~�a<��a<��a<~�a<L�a<�a<��a<��a<F�a<�za<"ca<EHa<e,a<�a<��`<��`<��`<b�`<��`<?�`<��`<>�`<.a<+a<�Ea<�^a<\ta<b�a<n�a<'�a<"�a<��a<�a<��a<.�a<��a<��a<X�a<�a<�a<Ƈa<%�a<v�a<G�a<��a<��a<�a<��a<Ña<�a<�ua<�`a<bHa<�-a<�a<��`<r�`<��`<��`<V�`<��`<�`<��`<��`<a<+a<�  �  �Ga<`a<
ua<Ʌa<ёa<,�a<�a<|�a<r�a<��a<��a<�a<h�a<<�a<��a<m�a<��a<^�a<��a<ɘa<ŝa<'�a<ˡa<a<�a<݊a<�ya<�da<�La<�2a<3a<Na<U�`<��`<��`<��`<�`<^�`<��`<�a<)/a<�Ja<ea<(}a<��a<f�a<��a<��a<T�a<m�a<{�a<K�a<٨a<��a<]�a<%�a<�a<��a<Ϩa<H�a<`�a<O�a<�a<��a<r�a<	�a<ܳa<��a<a�a<�|a<�ca<�Ia<�/a<�a<�a<��`<n�`<^�`<a�`<-
a<fa<�6a<�Pa<Nka<s�a<��a<��a<�a<��a<��a<Q�a<��a<x�a<H�a<)�a<ɱa<�a<t�a<(�a<��a<|�a<��a<��a<��a<`�a<��a<X�a<��a<x�a<y�a<�a<(xa<"^a<�Ca<.*a<a<�a<��`<f�`<��`<� a<ya<�&a<@a<cZa<ita<��a<6�a<��a<M�a<K�a<��a<��a<f�a<�a<��a<��a<��a<�a<תa<��a<��a<��a<��a<�a<1�a<��a<��a<�a<��a<Ūa<�a<?�a<Eja<�Oa<^5a<�a<�a<L�`<p�`<��`<�`<S�`<�a<P(a<�Aa<�[a<Gua<�a<�a<��a<2�a<"�a<��a<��a<��a<+�a<�a<��a<P�a<p�a<��a<��a<*�a<�a<��a<�a<�a<c�a<��a<��a<'�a<�a<|a<|da<$Ja<�.a<+a<�`<.�`<9�`<�`<G�`<��`<��`<=�`<�a<�-a<RGa<�_a<pua<�a<ٓa<�a<��a<�a<j�a<��a<��a<d�a<��a<D�a<l�a<��a<ۄa<j�a<.�a<O�a<��a<;�a<6�a<ǘa<��a<��a<eva<�aa<�Ia<�/a<!a<��`<��`<&�`<2�`<�`<u�`<��`<��`<Z�`<�a<G-a<�  �  �La<da<�wa<O�a<�a<�a<��a<��a<��a<܍a<��a<�a<�}a<Y{a<�za<�|a<)�a<��a<�a< �a<N�a<��a<��a<ҝa<��a<��a< }a<ia<�Qa<b9a<� a<�	a<��`<S�`<|�`<��`<��`<��`<�a<Ra<6a<UPa<�ia<ڀa<�a<��a<C�a<b�a<��a<��a<@�a<˦a<{�a<��a<��a<<�a<��a<�a<x�a<Цa<ǭa<�a<
�a<��a<��a<��a<޴a<(�a<�a<��a<~ia<}Pa<�7a<}!a<:a<�a<Y�`<D�`<#a<va<�&a<>a<�Wa<�pa<܈a<֝a<��a<ºa<�a<��a<(�a<j�a<Ӻa<z�a<w�a<Y�a<�a<{�a<@�a<��a<i�a<T�a<��a<�a<��a<�a<��a<׿a<�a<#�a<�a<!}a<8da<�Ja<A2a<a<6a<{a<[�`<� a<t
a<�a<1/a<;Ga<�`a<}ya<��a<�a<%�a<��a<�a<r�a<N�a<��a<c�a<ذa<��a< �a<��a<ܡa<)�a<!�a<�a<Ӱa<�a<��a<��a<��a<'�a<C�a<��a<,�a<��a<�oa<RVa<�<a<%a<a<
a<S�`<|�`<��`<�a<qa< 0a<�Ha<�aa<�ya<��a<i�a<��a<�a<��a<7�a<��a<��a<��a<��a<S�a<��a<��a<��a<�a<ӗa<��a<�a<��a<�a<��a<ϭa<:�a<(�a<!�a<�a<ia<�Oa<�5a<�a<�a<��`<�`<�`<,�`<R�`<��`<�a<Ta<4a<�La<Nda<�xa<�a<��a<K�a<��a<Y�a<�a<�a<.�a<��a<%a<|{a<uya<�ya<A|a<X�a<��a<�a<�a<��a<��a<m�a<�a<��a<ya<�ea<�Na<�5a<@a<�a<��`<��`<
�`<�`<V�`<f�`<��`<�a<�a<�3a<�  �  �Ta<�ia<�{a<i�a<(�a<A�a<�a<*�a<ˋa<)�a<w|a<ua<�oa<�la<la<�ma<�ra<3ya<&�a<��a<֑a<��a<d�a<��a<4�a<3�a<M�a<Zoa<PZa<RCa<j,a<�a<�a<��`<y�`<��`<��`<�a<Ka<�(a<�@a<|Ya<qa<�a<A�a<�a<ʫa<�a<�a<��a<��a<��a<��a<��a<@�a<��a<A�a<f�a<H�a<ۚa<f�a<6�a<9�a<D�a<2�a<�a<�a<S�a<Ǜa<��a<~ra<�Za<Da<%/a<a<Aa<{a<La<�a<�!a<M4a<"Ja<�aa<_ya<Z�a<J�a<X�a<��a<�a<��a<�a<%�a<��a<��a<2�a<ܛa<k�a<ȕa<��a<�a<��a<֦a<Ӯa<Ӷa<��a<�a<�a<ÿa<��a<�a<��a<�a<�ma<�Ua<?a<+a<ha<Ra<�a<ra<�a<�(a<3<a<�Ra<:ja<v�a<Z�a<��a<@�a<��a<^�a<��a<��a<��a<��a<��a<�a<�a<C�a<&�a<o�a<|�a<��a<ݥa<��a<<�a<E�a<j�a<�a<иa<�a<x�a<ɍa<xa<A`a<�Ha<]2a<ya<�a<Q	a<�a<�a<�a<5(a<�<a<�Sa<�ja<P�a<˔a<Ǥa<�a<t�a<;�a<��a<�a<8�a<x�a<�a<F�a<4�a<υa<�a<d�a<��a<��a<��a<Ȟa<A�a<̩a<C�a<��a<[�a<J�a<|�a<#pa<�Xa<B@a<B(a<ga<d a<��`<&�`<3�`<��`<y a<$a<X'a<9>a<dUa<�ja<-}a<��a<P�a<G�a<��a<<�a<֐a<�a<j�a<rxa<�qa<�la<�ja<"ka<(na<�sa<zza</�a<�a<��a<��a<��a< �a<Ήa<�|a<Ska<�Va<>?a<t'a<�a<��`<��`<��`<C�`<7�`<��`<��`<�a<D%a<=a<�  �  �^a<Hqa<�a<܋a<��a<y�a<��a<?�a<_�a<jwa<Qma<zda<�]a<�Ya<�Xa<[a<�`a<�ha<�ra<n}a< �a<*�a<{�a<a�a<��a<H�a<�a<Uwa<�da<Pa<t;a<(a<�a<�a<�a<Ta<�	a<a<%a<�8a<�Na<�da<:za<��a<��a<��a<êa<S�a<ۧa<=�a<��a<�a<Ņa<H~a<�xa<Kva< wa<�za<ˁa<��a<��a<��a<>�a<��a<)�a<��a<^�a<Q�a<>�a<x�a<�}a<�ha<�Sa<�@a<51a<=&a<	!a<�!a<�(a<�4a<�Ea<mYa<�na<�a<��a<0�a<��a<2�a<�a<N�a<�a<��a<��a<Y�a<��a<�a<��a<��a<f�a<��a<~�a<o�a<ԡa<!�a<��a<d�a<��a<H�a<�a<��a<��a<��a<�ya<?da<�Oa<K=a<�.a<�%a<3"a<�$a<f-a<;a<�La<6aa<�va<a�a<̝a<�a<��a<v�a<��a<;�a<��a<N�a<�a<a�a<�a<�a<5�a<�a<��a<��a<؍a<;�a<z�a<a�a<ݳa<}�a<��a<7�a<)�a<�a<a<u�a<ma<�Wa<wCa<+2a<O%a<�a<Ca<� a<+a<:a<�La<Eaa<qva<m�a<��a<�a<��a<n�a<��a<��a<S�a<�a<��a<�a<�}a<�va<�ra<�qa<�sa<&ya<{�a<��a<Q�a<E�a<D�a<9�a<A�a<��a<G�a<�a<�xa<da<�Ma<8a<$a<�a<�a<�a<�a<�a<Qa<n#a<�6a<>Ka<`a<sa<�a<�a<��a<\�a<�a<�a<I�a<�|a<ra<�ga<�_a<Za<�Wa<Xa<�[a<rba<ka<2ua<<a<]�a<�a<m�a<��a<��a<��a<�ra<0`a<DKa<�5a<
!a<�a<o a<�`<��`<��`<P�`<,a<4a<�3a<_Ia<�  �  �ia<�ya<��a<	�a<~�a<ԏa<�a<��a<�ta<�ga<�[a<uPa<Ha<Ca<�Aa<�Da<CKa<Ua<8aa<�na<#|a< �a<��a<k�a<Øa<��a<��a<I�a<ipa<�^a<lLa<p;a<-a<r"a<�a<a<!a<)+a<k9a<�Ja<g^a<�qa<6�a<��a<��a<�a<C�a<��a<E�a<��a<�a<�~a<Gsa<�ia<�ba<�_a<4`a<�da<�la<xa<�a<˒a<^�a<Ϋa<4�a<��a<n�a<��a<?�a<1�a<h�a<xa<�ea<�Ta<-Ga<�=a<�8a<�9a<�?a<oJa<2Ya<�ja<�}a<�a<Ѡa<f�a<��a<��a<{�a<��a<0�a<�a<�a<=�a<o~a<�ta<gna<�ka<�la<�qa<2za<b�a<�a<;�a<}�a<x�a<�a<y�a<ٻa<s�a<̨a<6�a<��a<�ta<.ba<Ra<eEa<'=a<�9a<m<a<�Ca<Pa<�_a<�qa<��a<c�a<*�a<&�a<�a<��a<�a<��a<�a<��a<k�a<��a<ya<7pa<�ja<�ha<5ka<+qa<]za<�a<��a<�a<Ϊa<��a<��a<X�a<ܴa<�a<��a<�a<�{a<�ha<�Va<�Ga<,<a<|5a<4a<8a<%Aa<ZNa<�^a<qa<x�a<l�a<ݢa<�a<�a<�a<߯a<�a<��a<i�a<��a<�ta<!ia<�`a<�[a<�Za<�]a<2da<�ma<%ya<\�a<d�a<T�a<C�a<e�a<��a<�a<�a<��a<�pa<[]a<�Ia<8a<�)a<�a<ua<ta<�a<�(a<7a<�Ga<PZa<la<G|a<M�a<�a<w�a<Õa<s�a<l�a<�{a<Nna<�`a<�Ta<�Ja<�Ca<�@a<oAa<!Fa<)Na<Ya<fea<Wra<[~a<�a<o�a<��a<�a<W�a<�za<�ja<	Ya<�Ea<�3a<{#a<�a<�a<�a<(a<�a<'"a<	2a<IDa<}Wa<�  �  �ta<��a<��a<
�a<�a<1�a<E�a<lua<�fa<�Va<Ha<�:a<z0a<�*a<)a<a,a<�3a<�?a<2Na<6^a<�na<�}a<��a<m�a<&�a<��a<u�a<5�a<[|a<�ma<a^a<Pa<�Ca<j:a<�5a<;5a<�9a<RBa<Oa<(^a<�na<ma<t�a<#�a<��a<§a<��a<�a<j�a<|�a<�{a<�la<_a<Sa<�Ja<�Fa<sGa<�La<$Va<{ca<�ra<��a<ݓa<��a<S�a<̵a<�a<��a<�a<�a<z�a<�a<�xa<Rja<,^a<�Ua<�Qa<�Ra<�Wa<aa<$na<�|a<�a<Z�a<�a<s�a<��a<g�a<θa< �a<&�a<�a<�a<xwa<\ia<�]a<!Va<�Ra<6Ta<
Za<%da<�qa<��a<��a<�a<g�a<�a<��a<|�a<�a<��a<"�a<��a<��a<va<ha<�\a<�Ua<(Sa<MUa<�[a<@fa<�sa<�a<�a<��a<j�a<-�a<�a<��a<M�a<��a<��a<��a<m�a<qa<;ca<�Xa<2Ra<Pa<�Ra<�Ya<ea<�ra<6�a<�a<e�a<��a<��a<��a<��a<��a<��a<�a<֊a<�za<}ka<^a<%Ta<tNa<.Ma<�Pa<PXa<da< ra<h�a<�a<��a<�a<�a<�a<Y�a<P�a<�a<��a<�a<�oa<G`a<�Ra<�Ha<)Ca<Ba<�Ea<~Ma<7Ya<�fa<va<�a<�a<a�a<n�a<3�a<��a<��a<��a<�}a<Uma<�\a<�Ma<}@a<r7a<�2a<w2a<�6a<�?a<�Ka<"Za<�ia<bxa<��a<\�a<�a<;�a<�a<�a<f}a<�na<P^a<>Na<�?a<�3a<�+a<�'a<�(a<Z.a< 8a<KEa<Ta<da<�ra<	�a<|�a<�a<��a<��a<q�a<�ua<ga<�Va<mGa<|9a<P.a<h'a<�$a<'a<|-a<Q8a<-Fa<�Ua<�ea<�  �  �a<Z�a<r�a<@�a<�a<��a<�ya<ja<GXa<{Ea<�3a<m$a<�a<�a<�a<�a<�a<�)a<�:a<fMa<�`a<�ra<��a<�a<��a<��a<��a<z�a<�a<U|a<�oa<�ca<�Ya<BRa<3Na<Na<�Qa<YYa<�ca<�pa<�~a<a�a<K�a<��a<�a<ϧa<~�a<ߚa<��a<�}a<{la<[Za<�Ia<N<a<�2a<�-a<[.a<V4a<??a<*Na<`a<�sa<�a<ɘa<��a<L�a<��a<ɹa<�a<��a<'�a<��a<ߊa<�~a<�ta<$na<�ja<Bka<�oa<zwa<F�a<��a<Λa<U�a<��a<۹a<�a<V�a<��a<��a<��a<T�a<�va<da<�Sa<hFa<w=a<�9a<B;a<#Ba<�Ma<]a<�na<�a<;�a<��a<��a</�a<N�a<G�a<ҷa<��a<$�a<�a<3�a<�}a<Tta<Tna<la<�ma<5sa<�{a<G�a<�a<�a<��a<�a<��a<�a<f�a<�a<��a<R�a<,�a<�na<�\a<�La<�@a<J9a<�6a<:a<eBa<Oa<%_a<_qa<(�a<��a<�a<3�a<C�a<�a<��a<�a<��a<A�a<�a<_a<=ta<�ka<ga<�ea<�ha<Zoa<�xa<��a<9�a<ߝa<��a<p�a<��a<��a</�a<�a<��a<�a<�pa<@]a<2Ka<�;a<�0a< *a<�(a<S-a<�6a<�Ca<,Ta<Bfa<xa<L�a<a<�a<�a<��a<ʞa<�a<x�a<�|a<oa<4ba<LWa<�Oa<YKa<"Ka<�Na<�Ua<`a<�ka<lxa<_�a<6�a<Ɣa<w�a<-�a<�a<��a<�ra<aa<�Ma<�:a<�)a<Ka<�a<�a<�a<wa<�!a<�0a<MBa<-Ua<ga<Iwa<�a<f�a<V�a<$�a<��a<T�a<�ta<rga<�Za<�Na<�Ea<�?a<�=a<q?a<Ea<�Ma<�Ya<lfa<�sa<�  �  D�a<��a<�a<��a<��a<a<Yqa<�^a<Ja<�4a<� a<Xa<$a<�`< �`<#�`<8a<.a<(a<G=a<CSa<�ha<{a<n�a<�a<��a<��a<��a<-�a<g�a<�a<%va<na<ha<�da<�da<ha<�na<wa<��a<��a<��a<Πa<��a<k�a<0�a<X�a<t�a<��a<�qa<C]a<Ia<86a<�&a<�a<a<�a<"a<^)a<5:a<mNa<;da<�za<2�a<�a<֮a<��a<ֻa<?�a<��a</�a<��a<��a<ڑa<
�a<:�a<��a<��a<��a<"�a<��a<�a<:�a<ɲa<(�a<S�a<f�a<ιa<w�a<5�a<��a<|a<�fa<�Qa<&?a<80a<&a<�!a<�#a<W+a<g8a<�Ia<^a<psa<��a<כa<�a<��a<S�a<o�a<�a<��a<1�a<�a<��a<,�a<̉a<��a<��a<;�a<Ԉa<׏a<��a<;�a<H�a<&�a<M�a<!�a<n�a<�a<ܫa<�a<(�a<�sa<O^a<�Ia<�7a<,*a<�!a<a<�"a<,a<g:a<�La<;aa<�va<!�a<�a<��a<r�a<x�a<׺a<��a<ׯa<S�a<��a<��a<��a<΁a<�}a<�|a<a<��a<�a<��a<��a<8�a<�a<�a<��a<W�a<�a<��a<G�a<�wa<�aa<�Ka<{7a<8&a<�a<ca<>a<a<� a<�/a<�Ba<�Va<�ka<�~a<�a<u�a<��a<ĥa<�a<1�a<~�a<�a<�a<ua<Vla<�ea<.ba<�aa<�da<�ja<{ra<|a<؅a<Ԏa<��a<A�a<ɘa<��a<ɉa<{a<�ha<�Sa<�=a<�(a<�a<a<}�`<��`<@�`<��`<ia<�a<s1a<�Fa<�[a<zna<U~a<ԉa<Y�a<I�a<��a<��a<��a<{va<la<�ba<+[a<#Va<�Ta<�Ua<�Za<�aa<;ka<�ua<�a<�  �  �a<�a<��a<��a<�a<�{a<�ia<�Ta<�=a<4&a<a<��`<s�`<��`<��`<��`<��`<a<�a<"/a<]Ga<_a<ta<��a<�a<E�a<��a<c�a<��a<;�a<�a<��a<Ia<bza<�wa<.xa<�za<6�a<��a<�a<Әa< �a<ȧa<o�a</�a<]�a<Ҝa<i�a<7|a<ga<Pa<�9a<�$a<�a<�a<�a<a<1	a<Ka<�(a<�>a<�Va<loa<��a<��a<�a<��a<O�a<p�a<l�a<P�a<O�a<��a<�a<��a<זa<єa<*�a<�a<u�a<m�a<L�a<Q�a<f�a<A�a<��a<H�a<�a<�a<\�a<M�a<upa<�Xa<�Aa<7-a<�a<�a<=a<a<�a<�%a<�8a< Oa<�fa<n~a<��a<n�a<��a<�a<��a<��a<|�a<2�a<y�a<n�a<��a<ța<��a<B�a<A�a<�a<͠a<�a<�a<��a<�a<��a<��a<u�a<~�a<��a<y�a<a<}ga<�Oa<9a<d%a<va<@a<�
a<]a<�a<F(a<N<a<Sa<�ja<��a<�a<�a<m�a<�a<�a<Ƽa<+�a<&�a<�a<
�a<ݙa<!�a<ڐa<'�a<Αa<;�a<y�a<Уa<��a<��a<�a<^�a<��a<��a<��a<��a<�a<ma<�Ta<�<a<&a<Na<�a<��`<��`<-a<�a<fa<�2a<gIa<n`a<va<��a<��a<١a<;�a<�a<ߤa<��a<��a<��a<G�a<�}a<Exa<pua<ua<)wa<�{a<A�a<��a<�a<q�a<��a<Ҝa<��a<�a<\�a<,ta<�_a<AHa<0a<�a<�a<��`<l�`<V�`<��`<��`<��`<�a<�"a<�9a<OQa<�fa<�xa<�a<�a<��a<��a<�a<��a<܂a<�za<Ksa<"ma<ia<�ga<�ha<�la<�ra<Aza<c�a<`�a<�  �  ��a<��a<%�a<a�a<Ɇa<xwa<�ca<�La<�3a<�a<�a<��`<%�`<��`<U�`<+�`<��`<!�`<�
a<$a<�=a<[Wa<�na<�a<)�a<q�a<��a<}�a<��a<q�a<ݖa<?�a<�a<��a<��a<݆a<o�a<��a<��a<��a<ءa<F�a<ͬa<V�a<�a<|�a<��a<߉a<�ua<E^a<�Ea<{-a<ea<a<�`<��`<��`<~�`<�a<a<u2a<tLa<�fa<�a<ޕa<��a<��a<�a<�a<?�a<@�a<"�a<�a<�a<ڨa<j�a<��a<�a<^�a<r�a<.�a<i�a<��a<��a<��a<�a<��a<��a<��a</�a<�a<8ga<�Ma<5a<da<�a<!a<��`<%�`<%a<xa<�+a<hCa<�\a<va<�a<3�a<>�a<��a<&�a<_�a<��a<��a<�a<y�a<n�a<��a<c�a<��a<��a<ͨa<d�a<9�a<~�a<a�a<��a<G�a<]�a<=�a<E�a<��a<��a<wa<�]a<Da<�+a<4a<%a<U�`<G�`<��`<g	a<Qa<�/a<�Ga<@aa<�ya<��a<I�a<��a<@�a<�a<��a<S�a<[�a<�a<��a<��a<Q�a<��a<מa<u�a<��a<��a<|�a<��a<ʹa<�a<G�a<��a<��a<��a<�a<E}a<cda<oJa<b0a<�a<�a<�`<��`<��`<{�`<��`<�a<�&a< ?a<�Wa<oa<�a<��a<��a<��a<ªa<��a<��a<U�a<3�a<P�a<#�a<׆a<"�a<��a<��a<�a<�a<��a<Y�a<�a<�a<	�a<�a<k�a<�a<oa<*Xa<?a<5%a<�a<��`<��`<��`<�`<��`<��`<��`<T�`<�a<0a<�Ha<�`a<�ta<r�a<��a<��a<�a<}�a<=�a<G�a<ͅa<�a<�za<�wa<uva<�wa<�za<ca<t�a<��a<+�a<�  �  1�a<��a<L�a<�a<3�a<�ta<�_a<�Ga<�-a<ra<��`<��`<y�`<��`<b�`<W�`<�`<2�`<�a<�a<�7a<vRa<�ja<�a<Џa<q�a<e�a<�a<^�a<r�a<.�a<��a<9�a<1�a<��a<ӏa<7�a<�a<T�a<Z�a<k�a<��a<�a<B�a<Ҭa<��a<��a<��a<!qa<�Xa<B?a<�%a<�a<��`<H�`<��`<�`<��`<0�`<la<�*a<�Ea<�`a<{a<b�a<ۥa<��a<��a<��a<4�a<X�a<��a<��a<��a<;�a<,�a<w�a<ˬa<�a<��a<��a<ۼa<��a<��a<I�a<��a<ӿa<T�a<!�a<i�a<{a<Saa<�Fa<5-a<�a<Ta<P�`<�`<A�`<k�`<Ia<@#a<<a<�Va<�pa<��a<-�a<��a</�a<*�a<��a<J�a<U�a<��a<r�a<E�a<��a<;�a<�a<ܮa<X�a<Q�a<M�a<��a<�a<�a<��a<��a<�a<��a<��a<u�a<�qa<�Wa<�<a<�#a<a<x�`<o�`<Q�`<��`<��`<`a<�'a<�@a<=[a<	ua<��a<��a<R�a<?�a<}�a<s�a<�a<\�a<V�a<�a<ήa<�a<z�a<ͧa<>�a<�a<O�a<;�a<%�a<
�a<%�a<3�a<f�a<�a<��a<��a<�xa<�^a<�Ca<�(a<a<g�`<>�`<��`<��`<��`<��`<%a<�a<98a<�Qa<�ja<j�a<v�a<Пa<��a<��a<��a<��a<Ȥa<ٞa<ؘa<��a<��a<�a<��a<-�a<�a<S�a<�a<��a<��a<Ƣa<��a<;�a<4�a<za<>ka<fSa<$9a<4a<a<��`<E�`<��`<+�`<��`<��`<R�`<��`<|a<�)a<�Ca<D\a<�qa<��a<0�a<��a<9�a<ՙa<Ɩa<%�a<Ìa<��a<S�a<��a<na<y�a<!�a<N�a<��a<�a<זa<�  �  �a<~�a<��a<�a<�a<�ya<{]a<�<a<�a<<�`<Z�`<;�`<��`<r�`<�`<O�`<ƥ`<]�`<��`<� a<�%a<�Ia<Uja<=�a<Λa<%�a<�a<׷a<Y�a<��a<�a<��a<��a<b�a<��a<�a<E�a<��a<Q�a<��a<�a<��a<�a<��a<�a<Ҳa<��a<�a<�la<FKa<�'a<9a<-�`<��`<ַ`<F�`<��`<ڸ`<��`<�`<g	a<�-a<�Ra<va<��a<��a<��a<0�a<�a</�a<O�a<��a<G�a<��a<��a<�a<_�a<��a<��a<�a<:�a<Z�a<	�a<I�a<��a<!�a<t�a<^�a<'�a<z�a<�sa<�Pa<v,a<�	a<7�`<Z�`<Y�`<q�`<5�`<�`<��`<��`<�a<uAa<�ea<'�a<d�a<��a<k�a<��a<��a<��a<��a<��a<Z�a<��a<	�a<׿a<��a<t�a<K�a<��a<�a<$�a<S�a<��a<��a<q�a<�a<B�a<��a<؈a<�ga<yCa<Pa<��`<_�`<��`<��`<��`<P�`</�`<(�`<�a<X%a<XIa<�la<ʌa< �a<޼a<��a<��a<��a<��a<�a<��a<��a<8�a<лa<4�a<��a<�a<X�a<�a<��a<Q�a<��a<��a<Z�a<�a<��a<جa<��a<�ta<�Qa<�,a<Ta<��`<��`<͵`<��`<#�`<��`<��`<t�`<!�`<�a<:Ca<ea<�a<}�a<n�a<Y�a<��a<Ͽa<üa<K�a<��a<֩a<�a<��a<%�a<��a<P�a<ơa<L�a<իa<�a<��a<��a<l�a<8�a<��a<��a<�ka<�Ka<�'a<$a<��`<�`<��`<.�`<ݍ`<=�`<��`<6�`<��`<>�`<�a<�7a<Ya<va<�a<��a< �a<��a<��a<Z�a<�a<ӝa</�a<��a<_�a<4�a<9�a<>�a<�a<��a<٣a<W�a<�  �  ��a<۬a<X�a<S�a<Ґa< {a<V_a<1?a<a<��`<)�`<[�`<z�`<!�`<��`<�`<8�`<~�`<Q�`<+a<�(a<�Ka<�ka<>�a<t�a<P�a<Գa<�a<˵a<ʱa<C�a<q�a<J�a<z�a<��a<ʛa<W�a<Ţa<�a<	�a<i�a<��a<��a<Z�a<ӽa<e�a<{�a<?�a<�na<�Ma<'+a<�a<(�`<�`<k�`<ٲ`<-�`<|�`<�`< �`<�a<�0a<�Ua<?xa<�a<n�a<��a<$�a<��a<�a<x�a<��a<W�a<<�a<�a<-�a<D�a<��a<	�a<^�a<�a<��a<��a<��a<��a<��a<��a<�a<�a<�a<va<�Sa<�/a<'a<O�`<��`<�`<��`<��`<��`<��`<}�`<� a<�Da<=ha<�a<��a<b�a<��a<��a<!�a<��a<��a<��a<]�a<;�a<#�a<�a<y�a<z�a<h�a<0�a<�a<��a<G�a<J�a<'�a<F�a<��a<��a<Ŧa<��a<$ja<�Fa<�"a<� a<��`< �`<B�`<!�`<�`<��`<K�`<za<�(a<eLa<oa<o�a<�a<��a<��a<}�a< �a<	�a<O�a<�a<x�a<��a<�a<-�a<y�a<�a<��a<��a<��a<��a<��a<��a<��a<��a<�a<��a<�a<�va<nTa<�/a<�a<��`<��`<a�`<�`<��`<F�`<�`<��`<� a<#a<
Fa<-ga<\�a<^�a<�a<M�a<��a<��a<�a<�a<��a<��a<X�a<��a<
�a<��a<`�a<�a<+�a<�a<��a<�a<��a<�a<N�a<A�a<ևa<Dma<�Ma<�*a<ja<X�`<�`<��`<�`<`�`<�`<:�`<R�`<~�`<��`<a<e:a<�Za<Awa<Սa<#�a<�a<�a<X�a<[�a<{�a<ؚa<��a<��a<k�a<�a<@�a<\�a<\�a<��a<:�a<L�a<�  �  R�a</�a<K�a<	�a<1�a< a<�da<Fa<�$a<ua<t�`<��`<��`<�`<Y�`<ʧ`<%�`<��`<?�`<�a<�0a<�Ra<Cqa<�a<��a<��a<|�a<��a<%�a<��a<D�a< �a<h�a<Ǒa<��a<��a<i�a<��a<�a<h�a<q�a<f�a<�a<F�a<U�a<��a<U�a<͏a<�ta<kUa<4a<
a<��`<��`<��`<��`<�`<�`<��`<��`<ma<	:a<%]a<l~a<��a<q�a<�a<��a<��a<u�a<Y�a<��a<��a<Z�a<��a<F�a<�a<{�a<=�a<T�a<�a<X�a<Y�a<��a<��a<X�a<��a<��a<��a<5�a<�|a<�[a<'9a<�a<\�`<��`<��`<��`<��`<��`<k�`<�
a<�*a<SMa<Poa<َa<ɩa<�a<��a<��a<��a<q�a<�a<��a<g�a<ݹa<��a<ݯa<?�a<n�a<زa<��a<�a<��a<f�a<��a<y�a<8�a<��a<[�a<Ūa<N�a<
qa<&Oa<�,a<a<��`<N�`<�`<��`<��`<��`<q�`<ka<;2a<�Ta<�ua<��a<��a<��a<�a<'�a<��a<d�a<�a<�a<�a<��a<5�a<�a<A�a<'�a<?�a<��a<��a<��a<��a< �a<��a<}�a<n�a<��a<t�a<�|a<�[a<�8a<$a<A�`<X�`<��`<�`<��`<��`<��`<V�`<'a<!,a<�Ma<Zma<�a<b�a<��a<	�a<��a<�a<εa<�a<+�a<��a<$�a<ُa<ٌa<��a<��a<�a<��a<Ӡa<B�a</�a<t�a<��a<p�a<*�a<F�a<fra<=Ta<�2a<�a<�`<�`<ѷ`<��`<-�`<��`<��`<��`<��`<��`<�a<xAa<�`a<u{a<c�a<�a<�a<��a<2�a<��a<�a<�a<U�a<%�a<i�a<�~a<7�a<σa<щa<b�a<��a<m�a<�  �  P�a<Υa<��a<ޡa<��a<ׄa<.ma<�Pa<�1a<a<�`<�`<L�`<V�`<=�`<�`<��`<��`<t�`<�a<e=a<�\a<�xa<*�a<I�a<��a<C�a<��a<�a<�a<S�a<��a<Q�a</a<�{a<�{a<Ba<��a<��a<Y�a<��a<}�a<��a<μa<��a<X�a<��a<}�a<�}a<aa<1Ba<R#a<a<��`<��`<S�`<��`<%�`<��`<`
a<�'a<dHa<ia<Ƈa<��a<�a<��a<m�a<��a<��a<��a<U�a<�a<L�a<�a<A�a<y�a<ޙa<��a<�a<�a<'�a<��a<��a<[�a<��a<��a<h�a<��a<��a<��a<�ga<Ha<�(a<;a<��`<�`<��`<3�`<��`<a<�a<�:a<�Za<nza<W�a<�a<��a<��a<��a<��a<��a<r�a<O�a<ϲa<>�a<��a<w�a<��a<��a<��a<ԧa<�a<i�a<��a<��a<�a<��a<j�a<��a<��a<��a<�{a<b\a<*<a<�a<=a<��`<�`<��`<�`<�`<�a<�"a<fAa<Baa<�a<z�a<��a<_�a<Y�a<��a<��a<��a<��a<�a<��a<��a<��a<|�a<��a<��a<u�a<^�a<�a<(�a<��a<��a<Z�a<��a<	�a<��a<!�a<օa<�ga<�Fa<k&a<{a<A�`<��`<��`<A�`<��`<��`<��`<�a<}:a<�Ya<�va<�a<ڣa<z�a<��a<��a<<�a<0�a<��a<e�a<��a<��a<�|a<Bya<�xa<�{a<ȁa<��a<��a<x�a<3�a<,�a<�a<��a<��a<H�a<�ya<6^a<&?a<�a<�`<��`<$�`<Ѽ`<�`<5�`<J�`<O�`<��`<va<=-a<�La<?ia<��a<	�a<�a<��a<u�a<{�a<�a<��a<Q�a<�ya<ra<ma<Qka<�la<�qa<ya<��a<%�a<��a<�  �  ��a<t�a<�a<R�a<k�a<�a<�wa<�^a<�Ba<�%a<�
a<��`<�`<�`<I�`<��`<�`<�`<\a<�/a<iMa<�ia<��a<��a<b�a<��a<��a<�a<�a<��a<'�a<Qya<{na<�fa<ba<ba<�ea<�ma<ya<ʆa<=�a<\�a<h�a<��a<Һa<�a<��a<��a<H�a<�oa<�Sa<8a<ja<<	a<�`<D�`<��`<]�`<�a<�!a<=a<jZa<xa<��a<(�a<Q�a<��a<��a<��a<e�a<��a<&�a<ءa<�a<��a<�a<�a<�a<��a<�a<7�a<��a<�a<�a<��a<��a<�a< �a<��a<�a<$�a<�wa<�Za<�>a<c%a<>a<ya<��`<��`<�
a<2a<�3a<�Na<�ka<w�a<�a<\�a<��a<��a<,�a<��a<X�a<~�a<*�a<��a<�a<c�a<�a<��a<E�a<7�a<p�a<u�a<�a<0�a<+�a<��a<��a<��a<��a<��a<�a<��a<ma<�Oa<-4a<0a<�	a<7�`<��`<��`<�a<�a<�8a<~Ta<Mqa<��a<�a<k�a<}�a<�a<N�a<��a<5�a<|�a<�a<W�a<��a<�a<�{a<�za<�}a<��a<��a<[�a<��a<��a<I�a< �a<��a<��a<��a<L�a<U�a</va<�Xa<5;a<�a<�a<��`<��`<@�`<'�`<�a<ca<�0a<�La<�ha<��a<��a<F�a<j�a<$�a<��a<�a<v�a<��a<-�a<Kwa<la<�ca<`_a<_a<ca<�ja<Jua<�a<�a<L�a<��a<�a<کa<V�a<g�a<�a<�ja<�Na<l1a<�a<�`<u�`<A�`<�`<��`<6�`<}�`<~a<�!a<F>a<�Za<ta<
�a<D�a<�a<B�a<��a<"�a<*�a<�}a<
pa<�ca<�Ya<{Sa<nQa<Sa<:Ya<�ba<�na<�|a<>�a<�  �  O�a<D�a<��a<�a<�a<L�a<ɂa<�ma<UUa<D<a<?$a<Za<��`<��`<��`<\�`<a<�a<v,a<�Ea<g_a<�wa<��a<�a< �a<��a<��a<Ξa<�a<�a<4qa<'aa<kSa<]Ia<�Ca<iCa<Ha<�Qa<�_a<[pa<w�a<��a<p�a<Ӱa<�a<�a<J�a<J�a<̕a<�a<�ga<�Oa<9a<V&a<)a<la<�a<�a<�(a<�<a<Ua<�na<��a<��a<9�a<s�a<H�a<��a<t�a<ݻa<��a<לa<a<�{a<�na<\ea<�`a<�aa<Qga<�qa<�a<D�a<��a<o�a<V�a<M�a<��a<W�a<��a<�a<�a<S�a<pa<eWa<�@a</a<#a<�a< a<P)a<�8a<�Ma<�ea<a<��a<ƭa<#�a<��a<��a<X�a<��a<z�a<Ϊa<v�a<L�a<�xa<�la<�da<�aa<da<qka<�va<�a<іa<�a<�a<��a<��a<��a<�a<�a<,�a<{�a<�a<ffa<�Ma<�8a<C(a</a<.a<va<�*a<�;a<�Qa<&ja<R�a<�a<��a<ܾa< �a<��a<F�a<ʽa<&�a<��a<��a<-}a<�na<�ca<X]a<\a<�_a<�ha<9ua<�a<ٕa<��a<N�a<Y�a<�a<��a<v�a<�a<םa<_�a<�la<�Ra<p:a<&a<a<�a<ra<sa< a<I2a<�Ha<�`a<?ya<~�a<��a<j�a<մa<��a<Y�a<��a<�a<9�a<oa<&^a<%Pa<�Ea<�@a<�@a<�Ea<\Oa<�\a<�la<�}a<ȍa<#�a<��a<J�a<��a<c�a<�a<�xa<m`a<�Fa<�-a<�a<>a<��`<P�`<��`<��`<a<� a<j8a<}Qa<�ia<�a<ѐa<+�a<�a<s�a<˗a<J�a<�{a<ja<�Xa<qIa<`=a<t5a<�2a<�4a<z<a<6Ha<fWa<�ha<'za<�  �  H|a<��a<�a<��a<��a< �a<Ǎa<�|a<�ha<^Sa<?a<R-a<�a<�a<ta<�a<�#a<43a<xFa<�[a<�qa<
�a<�a<�a<Ĩa<�a<�a<*�a<ނa<�na<Za<Fa<�5a<l)a<�"a<�!a<�'a<3a<vCa<�Wa<�ma<ăa<֗a<��a<��a<ĸa<S�a<��a<�a<��a<�|a<	ha<Ua<(Ea<�9a<94a<�4a<�;a<Ha<AYa<�ma<��a<ʙa<D�a<��a<��a<��a<��a<��a<��a<9�a<d�a<\sa<`a<Pa<�Da<w?a<;@a<6Ga<�Sa<�da<�xa<=�a<��a<7�a<N�a<��a<��a<+�a<��a<��a<W�a<��a<qa<�]a<�Na<mDa<�?a<�Aa<�Ia<Wa<�ha<A}a<�a<e�a<1�a<n�a<��a<��a<*�a<��a<�a<#�a<��a<�na<\a<nMa<Da<Z@a<*Ca<�Ka<�Ya<�ka<��a<��a<ީa<ܺa<��a<�a<��a<��a<+�a<��a<O�a<�}a<�ha<�Va<�Ha<�?a<(=a<�@a<gJa<!Ya<�ka<z�a<ӕa<L�a<��a<��a<��a<��a<��a<)�a<#�a<��a<�va<�ba<�Pa<�Ca<$<a<�:a<N?a<�Ia<Ya<la<�a<�a<��a<�a<��a<n�a<}�a<*�a<�a<��a<d�a<ka<sVa<�Da<�7a<t0a<H/a<l4a<"?a<�Na<�aa<va<M�a<8�a<e�a<�a<,�a<�a<z�a<g�a<��a<�la<�Va<hBa<�1a<�%a<Ha<La<�%a<[1a<�Aa<+Ua<$ja<M~a<�a<��a<a�a<ڦa<Сa<��a<8�a<kra<�\a<Ga<�3a<�#a<'a<?a<�a<Sa<X*a<�;a<�Oa<Qea<�ya<�a<�a<K�a<	�a<I�a<��a<�}a<�ia<;Ta<\?a<�,a<a<�a<a<a<�a<&+a<�=a<MRa<ha<�  �  ]ma<Ղa<q�a<�a<G�a<�a<��a<�a<{a<�ia<+Ya<�Ja<q?a<�8a<�6a<:a<Ca<�Oa<�_a<vqa<L�a<]�a<�a<ݧa<��a<��a<�a<��a<�ra<�Za<YBa<+a<Ta<�a<� a< a<ga<�a<�&a<2>a<�Wa<ra<`�a<�a<�a<��a<s�a<Ƕa<r�a<B�a<X�a<�a<Cpa<Nca<Za<�Ua<;Va<�[a<|fa<�ta<�a<$�a<�a<"�a<��a<~�a<�a<��a<��a<��a<�a<sa<_Za<yCa<�0a<�#a<�a<ma<�&a<�4a<�Ha<�`a<�ya<��a<.�a<N�a<��a<�a<��a<*�a<}�a<X�a<+�a<�a<Aza<�ma<	ea<taa<�ba<�ia<�ta<U�a<5�a<��a<,�a<��a<��a<��a<��a<�a<B�a<s�a<f�a<ma<�Ta<�>a<y-a<�"a<]a<�!a<�+a<<a<UQa<�ia<Ăa<�a<�a<T�a<��a<p�a<��a<�a<�a<��a<�a<�a<�sa<:ha<�`a<�^a<�aa<�ia<�ua<�a<�a<G�a<��a<��a<��a<��a<3�a<:�a<��a<A�a<{xa<#_a<Ga<�2a<S#a<[a<�a<a<?*a<;<a<�Ra<9ka<&�a<7�a<��a<��a<T�a<��a<c�a<y�a<��a<�a<�a<�qa<�ba<Xa<�Qa<�Pa<�Ta<�]a<9ja<�ya<A�a<n�a<�a<�a<z�a<��a<1�a<{�a<p�a<rqa<~Wa<�=a<�%a<Sa<�a<k�`<��`<�a<�a<�%a<=a<�Ua<�ma<��a<��a<��a<8�a<K�a<B�a<�a<f�a<�qa<`a<�Oa<�Ba<�9a<�5a<�6a<0=a<�Ga<CVa<�fa<xa<O�a<~�a<h�a<}�a<�a<(�a<?�a<Noa<%Wa<�=a<$%a<+a<�`</�`<&�`<t�`<��`<Qa<�"a<e;a<�Ta<�  �  �^a<�wa<R�a<֚a<̢a<h�a<�a<a�a<Z�a<2~a<�pa<#ea<J\a<�Va<�Ua<zXa<�_a<�ia<�va<�a<��a<��a<��a<q�a<3�a<��a<��a<�|a<|ca<�Ga<V+a<�a<��`<�`<��`<��`<��`<��`<@a<�%a<�Ba<�`a<�|a<N�a<��a<��a<:�a<u�a<A�a<�a<��a<[�a<�a<�~a<�wa<ta<�ta<�ya<:�a<ʍa<֛a<6�a<�a<h�a<��a<��a<d�a<��a<B�a<��a<�za<i^a<,Ba<j(a<ha<�a<]�`<I�`<ya<�a<^.a</Ia<�ea<��a<��a<�a<`�a<D�a<��a<.�a<��a<j�a<4�a<��a<�a<�a<�a<8�a<?�a<��a<��a<Z�a<��a<w�a<�a<n�a<��a<��a<��a<[�a<��a<#�a</ta<9Wa<9;a<�"a<Za<�a<�`<�a<Ra<�a<�7a<[Sa<(pa<<�a<��a<4�a<]�a<��a<3�a<��a<e�a<��a<c�a<��a<n�a<�a<a<�}a<�a<#�a<��a<!�a<��a<¶a<M�a<,�a<X�a<b�a<�a<@�a<��a<Ła<ea< Ha<�,a<�a<|a<F�`<c�`<��`<�a<� a<":a<&Va<�ra<��a<ʤa<Ѷa<R�a<_�a<�a<F�a<g�a<��a<o�a<L�a<y~a<~ua<Npa<Ooa<Rra<Rya<3�a<��a<U�a<��a<`�a<+�a<��a<��a<ئa<0�a<I|a<�`a<�Ba<�%a<�
a<��`<*�`<4�`<_�`<��`<��`<ta<�%a<�Aa<�]a<�wa< �a<�a<h�a<i�a<A�a<>�a<q�a<��a<�va<|ia<_a<�Wa<}Ta<$Ua<:Za<�ba<Dna<�{a<׈a<(�a<V�a<C�a<o�a<7�a<��a<�ya<aa<�Da<�'a<�a<?�`<�`<_�`<��`<��`<r�`<�`<O	a<2%a<JBa<�  �  /Qa<�ma<a�a<+�a<��a<r�a<��a<Y�a<ߘa<ώa<��a<�{a<�ta<pa<�oa<�qa<�wa<�a<�a<�a<y�a<"�a<R�a<ŭa<7�a<6�a<܉a<�qa<IUa<P6a<a<��`<D�`<�`<��`<��`<w�`<��`<?�`<a<G0a<Qa<rpa<I�a<Ǣa<,�a<�a<��a<�a<�a<��a<�a<ŝa<��a<{�a<�a<��a<��a<��a<��a<�a<2�a<��a<j�a<]�a<��a<A�a< �a<��a<��a<�ka<5La<�,a<�a<_�`<=�`<X�`<c�`<d�`<l�`<1a<�4a<bTa<#ta<��a<�a<��a<��a<��a<��a<w�a<��a<�a<i�a<��a<ơa<X�a< �a<	�a<I�a<U�a<��a<��a<a�a<e�a<\�a<�a<�a<��a<��a<ўa<��a<�ca<�Ca<(%a<
a<��`<
�`<
�`<��`<��`<�a<k!a<�?a<�_a<�~a<՚a<A�a<��a<��a<>�a<�a<`�a<�a<�a<o�a<�a<��a<Ҙa<p�a</�a<3�a<ѥa<B�a<��a<��a<x�a<��a<��a<k�a<��a<��a<��a<�sa<�Sa<�3a<�a<|�`<��`<{�`<X�`<!�`<V�`<�a<�$a<�Ca<8ca<C�a<Ûa<۰a<οa<7�a<Q�a<��a<}�a<Y�a<"�a<%�a<��a<o�a<,�a<1�a<n�a<��a<a�a<��a<Q�a< �a<c�a<Ӽa<�a<װa<<�a<��a<Cpa<UQa<�0a<Ta<�`<��`<��`<0�`<{�`<��`<%�`<H�`<a<H0a<wOa<Ula<!�a<;�a<�a<g�a<��a<��a<Şa<b�a<j�a<Ba<�va<�pa<`na<�na<�ra<�ya<k�a<��a<��a<��a<D�a<��a<��a<�a<�a<�oa<�Sa<�4a<�a<��`<��`<r�`<ȷ`<�`<�`<��`<O�`<�`<�a<�1a<�  �  tFa<�ea<�a<�a<ϡa<)�a<+�a<��a<�a<b�a<��a<�a<�a<��a<8�a<I�a<��a<M�a<T�a<�a<�a<��a<@�a<�a<�a<l�a<��a<ia<	Ja<�(a<a<�`<��`<S�`<n�`<�`<O�`<h�`<~�`<;�`<�!a<�Da<�fa<�a<�a<۰a<#�a<j�a<S�a<=�a<��a<e�a<{�a<M�a<C�a<��a<E�a<��a<%�a<�a<��a<u�a<�a<�a<X�a<?�a<;�a<f�a<}�a<�a<�_a<�=a<Ha<�`<=�`<&�`<��`<��`<��`<��`<a<`$a<uFa<�ha<��a<b�a<��a<y�a<��a<>�a<��a<��a<��a<��a<�a<��a<��a<��a<��a<ӱa<[�a<��a<��a<��a<��a<4�a<�a<��a<��a<K�a<�a<�xa<'Wa<�4a<�a<��`<?�`<��`<�`<��`<��`<��`<�a<40a<�Ra<�sa<��a<��a<u�a<��a<��a<��a<��a<��a<��a<h�a<ӵa<�a<S�a<�a<��a<<�a<W�a<��a<��a<��a<�a<��a<��a<;�a<�a<_�a<�a<Uha<9Fa<�#a<a<��`<��`<��`<��`<��`<�`<�`<�a<�4a<�Va<qwa<l�a<��a<{�a<D�a< �a<U�a<��a<I�a<w�a<ۮa<��a<6�a<ǝa<ǜa<\�a<>�a<R�a<C�a<��a<��a<�a<Ͽa<@�a<Ӯa<��a<o�a<�fa<JEa<#"a<��`<��`<��`<ʹ`<o�`<�`<�`<P�`<'�`<� a<["a<�Ca<kca<�~a<+�a<��a<<�a<H�a<G�a<קa<5�a<��a<��a<��a<7�a<�a<w�a<V�a<��a<��a<g�a<�a< �a<�a<��a<�a<��a<w�a<�ga<tIa<�'a<da<��`<��`<�`<y�`<��`<��`< �`<��`<{�`<a<�$a<�  �  �?a<�_a<�{a<��a</�a<I�a<�a<�a<רa<�a<Мa< �a<��a<	�a<o�a<H�a<��a<��a<3�a<B�a<~�a<Ĳa<��a<��a<�a<ʕa<Ma<:ca<�Ba<�a<�`<��`<&�`<�`<��`<�`<��`<��`<��`<��`<.a<�<a<>`a<�a<��a<�a<�a<��a<��a<$�a<�a<��a<(�a<d�a<�a<��a<s�a<r�a<R�a<��a<��a<#�a<�a<��a<�a<f�a<��a<H�a<��a<�ya<Xa<�4a<�a<7�`<��`<��`<��`<�`< �`<�`<h�`<,a<�=a<Gaa<��a<�a<��a<?�a<B�a<q�a<��a<E�a<��a<V�a<1�a<��a<��a<�a<��a<}�a<*�a< �a<��a<��a<p�a<+�a<R�a<�a<��a<��a<��a<�qa<�Na<+a<�a<��`<A�`<��`<P�`<��`<��`<W�`<�a<q&a<Ja<)ma</�a<��a<)�a<Y�a<�a<\�a<��a<{�a<W�a<��a<x�a<��a<d�a<B�a<��a<��a<��a<��a<�a<��a<"�a<N�a<��a<:�a<J�a<�a<D�a<.aa<x=a<�a<��`<\�`<T�`<�`<��`<H�`<J�`<�`<	a<+a<Oa<qa<_�a<��a<��a<9�a<��a<��a<��a<��a<��a<��a<�a<	�a<�a<��a<>�a<k�a<"�a<��a<D�a<��a<��a<��a<h�a<,�a<��a<�a<�`a<�=a<�a<(�`<��`<�`<(�`<��`<
�`<e�`<ǻ`<��`<��`<ua<�<a<t]a< za<d�a<\�a<Ӭa<y�a<*�a<A�a<H�a<Q�a<��a<	�a<+�a<*�a<��a<��a<Y�a<�a<N�a<8�a<��a<�a<�a<��a<ڒa<�}a<�ba<�Ba<�a<��`<��`<e�`<��`<��`<0�`<��`<�`<��`<G�`<S�`<Ca<�  �  ?=a<.^a<�za<�a<ܠa<z�a<��a<[�a<�a<¥a<֟a<��a<��a<�a<��a<;�a<�a<�a</�a<Ϫa<x�a<�a<$�a<ïa<�a<�a<~a<Caa<N@a<�a<��`<��`<
�`<h�`<��`<��`<�`<K�`<j�`<��`<�a<
:a<^a<[~a<��a<b�a<�a<T�a<��a<��a<\�a<��a<P�a<�a<�a<Ʊa<��a<W�a<�a<�a<��a<��a<��a<��a<��a<l�a<��a<a�a<%�a<�wa<8Ua<@1a<(a<!�`<J�`<��`<1�`<W�`<o�`<��`<z�`<�a<T:a<�^a<��a<��a<�a<��a<W�a<��a<��a<9�a<Q�a<Q�a<��a<��a<}�a<�a<��a<`�a<��a<0�a<e�a<�a<��a<��a<��a<��a<��a<��a<�a<�oa<�Ka<�'a<a<��`<��`<3�`<ֹ`<�`<T�`<6�`<� a<#a<�Fa<�ja<b�a<��a<w�a<�a<F�a<
�a<f�a<��a<��a<��a<
�a<`�a<`�a<^�a<�a<��a<�a<��a<��a<��a<g�a<��a<��a<��a<��a<۝a<M�a<�^a<E:a<da<��`<@�`<��`<x�`<+�`<��`<��`<�`<la<=(a< La<�na<эa<��a<�a</�a<��a<��a<9�a<�a<��a<��a<ǵa<��a< �a<�a<#�a<%�a<\�a<��a<��a<j�a<��a<��a<n�a<��a<��a<~a<U^a<�:a<�a<��`<��`<ε`<}�`<�`<r�`<գ`<��`<��`<)�`<9a<�9a<i[a<�xa<��a<Сa<�a<�a<`�a<3�a<ɩa<K�a<�a<�a<�a<K�a<��a<��a<��a<�a<�a<^�a<�a<ҭa<>�a<k�a<5�a<�|a<�`a<t@a<�a<m�`<��`<B�`<}�`<��`<��`<�`<��`<��`<~�`<��`<"a<�  �  �?a<�_a<�{a<��a</�a<I�a<�a<�a<רa<�a<Мa< �a<��a<	�a<o�a<H�a<��a<��a<3�a<B�a<~�a<Ĳa<��a<��a<�a<ʕa<Ma<:ca<�Ba<�a<�`<��`<&�`<�`<��`<�`<��`<��`<��`<��`<.a<�<a<>`a<�a<��a<�a<�a<��a<��a<$�a<�a<��a<(�a<d�a<�a<��a<s�a<r�a<R�a<��a<��a<#�a<�a<��a<�a<f�a<��a<H�a<��a<�ya<Xa<�4a<�a<7�`<��`<��`<��`<�`< �`<�`<h�`<,a<�=a<Gaa<��a<�a<��a<?�a<B�a<q�a<��a<E�a<��a<V�a<1�a<��a<��a<�a<��a<}�a<*�a< �a<��a<��a<p�a<+�a<R�a<�a<��a<��a<��a<�qa<�Na<+a<�a<��`<A�`<��`<P�`<��`<��`<W�`<�a<q&a<Ja<)ma</�a<��a<)�a<Y�a<�a<\�a<��a<{�a<W�a<��a<x�a<��a<d�a<B�a<��a<��a<��a<��a<�a<��a<"�a<N�a<��a<:�a<J�a<�a<D�a<.aa<x=a<�a<��`<\�`<T�`<�`<��`<H�`<J�`<�`<	a<+a<Oa<qa<_�a<��a<��a<9�a<��a<��a<��a<��a<��a<��a<�a<	�a<�a<��a<>�a<k�a<"�a<��a<D�a<��a<��a<��a<h�a<,�a<��a<�a<�`a<�=a<�a<(�`<��`<�`<(�`<��`<
�`<e�`<ǻ`<��`<��`<ua<�<a<t]a< za<d�a<\�a<Ӭa<y�a<*�a<A�a<H�a<Q�a<��a<	�a<+�a<*�a<��a<��a<Y�a<�a<N�a<8�a<��a<�a<�a<��a<ڒa<�}a<�ba<�Ba<�a<��`<��`<e�`<��`<��`<0�`<��`<�`<��`<G�`<S�`<Ca<�  �  tFa<�ea<�a<�a<ϡa<)�a<+�a<��a<�a<b�a<��a<�a<�a<��a<8�a<I�a<��a<M�a<T�a<�a<�a<��a<@�a<�a<�a<l�a<��a<ia<	Ja<�(a<a<�`<��`<S�`<n�`<�`<O�`<h�`<~�`<;�`<�!a<�Da<�fa<�a<�a<۰a<#�a<j�a<S�a<=�a<��a<e�a<{�a<M�a<C�a<��a<E�a<��a<%�a<�a<��a<u�a<�a<�a<X�a<?�a<;�a<f�a<}�a<�a<�_a<�=a<Ha<�`<=�`<&�`<��`<��`<��`<��`<a<`$a<uFa<�ha<��a<b�a<��a<y�a<��a<>�a<��a<��a<��a<��a<�a<��a<��a<��a<��a<ӱa<[�a<��a<��a<��a<��a<4�a<�a<��a<��a<K�a<�a<�xa<'Wa<�4a<�a<��`<?�`<��`<�`<��`<��`<��`<�a<40a<�Ra<�sa<��a<��a<u�a<��a<��a<��a<��a<��a<��a<h�a<ӵa<�a<S�a<�a<��a<<�a<W�a<��a<��a<��a<�a<��a<��a<;�a<�a<_�a<�a<Uha<9Fa<�#a<a<��`<��`<��`<��`<��`<�`<�`<�a<�4a<�Va<qwa<l�a<��a<{�a<D�a< �a<U�a<��a<I�a<w�a<ۮa<��a<6�a<ǝa<ǜa<\�a<>�a<R�a<C�a<��a<��a<�a<Ͽa<@�a<Ӯa<��a<o�a<�fa<JEa<#"a<��`<��`<��`<ʹ`<o�`<�`<�`<P�`<'�`<� a<["a<�Ca<kca<�~a<+�a<��a<<�a<H�a<G�a<קa<5�a<��a<��a<��a<7�a<�a<w�a<V�a<��a<��a<g�a<�a< �a<�a<��a<�a<��a<w�a<�ga<tIa<�'a<da<��`<��`<�`<y�`<��`<��`< �`<��`<{�`<a<�$a<�  �  /Qa<�ma<a�a<+�a<��a<r�a<��a<Y�a<ߘa<ώa<��a<�{a<�ta<pa<�oa<�qa<�wa<�a<�a<�a<y�a<"�a<R�a<ŭa<7�a<6�a<܉a<�qa<IUa<P6a<a<��`<D�`<�`<��`<��`<w�`<��`<?�`<a<G0a<Qa<rpa<I�a<Ǣa<,�a<�a<��a<�a<�a<��a<�a<ŝa<��a<{�a<�a<��a<��a<��a<��a<�a<2�a<��a<j�a<]�a<��a<A�a< �a<��a<��a<�ka<5La<�,a<�a<_�`<=�`<X�`<c�`<d�`<l�`<1a<�4a<bTa<#ta<��a<�a<��a<��a<��a<��a<w�a<��a<�a<i�a<��a<ơa<X�a< �a<	�a<I�a<U�a<��a<��a<a�a<e�a<\�a<�a<�a<��a<��a<ўa<��a<�ca<�Ca<(%a<
a<��`<
�`<
�`<��`<��`<�a<k!a<�?a<�_a<�~a<՚a<A�a<��a<��a<>�a<�a<`�a<�a<�a<o�a<�a<��a<Ҙa<p�a</�a<3�a<ѥa<B�a<��a<��a<x�a<��a<��a<k�a<��a<��a<��a<�sa<�Sa<�3a<�a<|�`<��`<{�`<X�`<!�`<V�`<�a<�$a<�Ca<8ca<C�a<Ûa<۰a<οa<7�a<Q�a<��a<}�a<Y�a<"�a<%�a<��a<o�a<,�a<1�a<n�a<��a<a�a<��a<Q�a< �a<c�a<Ӽa<�a<װa<<�a<��a<Cpa<UQa<�0a<Ta<�`<��`<��`<0�`<{�`<��`<%�`<H�`<a<H0a<wOa<Ula<!�a<;�a<�a<g�a<��a<��a<Şa<b�a<j�a<Ba<�va<�pa<`na<�na<�ra<�ya<k�a<��a<��a<��a<D�a<��a<��a<�a<�a<�oa<�Sa<�4a<�a<��`<��`<r�`<ȷ`<�`<�`<��`<O�`<�`<�a<�1a<�  �  �^a<�wa<R�a<֚a<̢a<h�a<�a<a�a<Z�a<2~a<�pa<#ea<J\a<�Va<�Ua<zXa<�_a<�ia<�va<�a<��a<��a<��a<q�a<3�a<��a<��a<�|a<|ca<�Ga<V+a<�a<��`<�`<��`<��`<��`<��`<@a<�%a<�Ba<�`a<�|a<N�a<��a<��a<:�a<u�a<A�a<�a<��a<[�a<�a<�~a<�wa<ta<�ta<�ya<:�a<ʍa<֛a<6�a<�a<h�a<��a<��a<d�a<��a<B�a<��a<�za<i^a<,Ba<j(a<ha<�a<]�`<I�`<ya<�a<^.a</Ia<�ea<��a<��a<�a<`�a<D�a<��a<.�a<��a<j�a<4�a<��a<�a<�a<�a<8�a<?�a<��a<��a<Z�a<��a<w�a<�a<n�a<��a<��a<��a<[�a<��a<#�a</ta<9Wa<9;a<�"a<Za<�a<�`<�a<Ra<�a<�7a<[Sa<(pa<<�a<��a<4�a<]�a<��a<3�a<��a<e�a<��a<c�a<��a<n�a<�a<a<�}a<�a<#�a<��a<!�a<��a<¶a<M�a<,�a<X�a<b�a<�a<@�a<��a<Ła<ea< Ha<�,a<�a<|a<F�`<c�`<��`<�a<� a<":a<&Va<�ra<��a<ʤa<Ѷa<R�a<_�a<�a<F�a<g�a<��a<o�a<L�a<y~a<~ua<Npa<Ooa<Rra<Rya<3�a<��a<U�a<��a<`�a<+�a<��a<��a<ئa<0�a<I|a<�`a<�Ba<�%a<�
a<��`<*�`<4�`<_�`<��`<��`<ta<�%a<�Aa<�]a<�wa< �a<�a<h�a<i�a<A�a<>�a<q�a<��a<�va<|ia<_a<�Wa<}Ta<$Ua<:Za<�ba<Dna<�{a<׈a<(�a<V�a<C�a<o�a<7�a<��a<�ya<aa<�Da<�'a<�a<?�`<�`<_�`<��`<��`<r�`<�`<O	a<2%a<JBa<�  �  ]ma<Ղa<q�a<�a<G�a<�a<��a<�a<{a<�ia<+Ya<�Ja<q?a<�8a<�6a<:a<Ca<�Oa<�_a<vqa<L�a<]�a<�a<ݧa<��a<��a<�a<��a<�ra<�Za<YBa<+a<Ta<�a<� a< a<ga<�a<�&a<2>a<�Wa<ra<`�a<�a<�a<��a<s�a<Ƕa<r�a<B�a<X�a<�a<Cpa<Nca<Za<�Ua<;Va<�[a<|fa<�ta<�a<$�a<�a<"�a<��a<~�a<�a<��a<��a<��a<�a<sa<_Za<yCa<�0a<�#a<�a<ma<�&a<�4a<�Ha<�`a<�ya<��a<.�a<N�a<��a<�a<��a<*�a<}�a<X�a<+�a<�a<Aza<�ma<	ea<taa<�ba<�ia<�ta<U�a<5�a<��a<,�a<��a<��a<��a<��a<�a<B�a<s�a<f�a<ma<�Ta<�>a<y-a<�"a<]a<�!a<�+a<<a<UQa<�ia<Ăa<�a<�a<T�a<��a<p�a<��a<�a<�a<��a<�a<�a<�sa<:ha<�`a<�^a<�aa<�ia<�ua<�a<�a<G�a<��a<��a<��a<��a<3�a<:�a<��a<A�a<{xa<#_a<Ga<�2a<S#a<[a<�a<a<?*a<;<a<�Ra<9ka<&�a<7�a<��a<��a<T�a<��a<c�a<y�a<��a<�a<�a<�qa<�ba<Xa<�Qa<�Pa<�Ta<�]a<9ja<�ya<A�a<n�a<�a<�a<z�a<��a<1�a<{�a<p�a<rqa<~Wa<�=a<�%a<Sa<�a<k�`<��`<�a<�a<�%a<=a<�Ua<�ma<��a<��a<��a<8�a<K�a<B�a<�a<f�a<�qa<`a<�Oa<�Ba<�9a<�5a<�6a<0=a<�Ga<CVa<�fa<xa<O�a<~�a<h�a<}�a<�a<(�a<?�a<Noa<%Wa<�=a<$%a<+a<�`</�`<&�`<t�`<��`<Qa<�"a<e;a<�Ta<�  �  H|a<��a<�a<��a<��a< �a<Ǎa<�|a<�ha<^Sa<?a<R-a<�a<�a<ta<�a<�#a<43a<xFa<�[a<�qa<
�a<�a<�a<Ĩa<�a<�a<*�a<ނa<�na<Za<Fa<�5a<l)a<�"a<�!a<�'a<3a<vCa<�Wa<�ma<ăa<֗a<��a<��a<ĸa<S�a<��a<�a<��a<�|a<	ha<Ua<(Ea<�9a<94a<�4a<�;a<Ha<AYa<�ma<��a<ʙa<D�a<��a<��a<��a<��a<��a<��a<9�a<d�a<\sa<`a<Pa<�Da<w?a<;@a<6Ga<�Sa<�da<�xa<=�a<��a<7�a<N�a<��a<��a<+�a<��a<��a<W�a<��a<qa<�]a<�Na<mDa<�?a<�Aa<�Ia<Wa<�ha<A}a<�a<e�a<1�a<n�a<��a<��a<*�a<��a<�a<#�a<��a<�na<\a<nMa<Da<Z@a<*Ca<�Ka<�Ya<�ka<��a<��a<ީa<ܺa<��a<�a<��a<��a<+�a<��a<O�a<�}a<�ha<�Va<�Ha<�?a<(=a<�@a<gJa<!Ya<�ka<z�a<ӕa<L�a<��a<��a<��a<��a<��a<)�a<#�a<��a<�va<�ba<�Pa<�Ca<$<a<�:a<N?a<�Ia<Ya<la<�a<�a<��a<�a<��a<n�a<}�a<*�a<�a<��a<d�a<ka<sVa<�Da<�7a<t0a<H/a<l4a<"?a<�Na<�aa<va<M�a<8�a<e�a<�a<,�a<�a<z�a<g�a<��a<�la<�Va<hBa<�1a<�%a<Ha<La<�%a<[1a<�Aa<+Ua<$ja<M~a<�a<��a<a�a<ڦa<Сa<��a<8�a<kra<�\a<Ga<�3a<�#a<'a<?a<�a<Sa<X*a<�;a<�Oa<Qea<�ya<�a<�a<K�a<	�a<I�a<��a<�}a<�ia<;Ta<\?a<�,a<a<�a<a<a<�a<&+a<�=a<MRa<ha<�  �  O�a<D�a<��a<�a<�a<L�a<ɂa<�ma<UUa<D<a<?$a<Za<��`<��`<��`<\�`<a<�a<v,a<�Ea<g_a<�wa<��a<�a< �a<��a<��a<Ξa<�a<�a<4qa<'aa<kSa<]Ia<�Ca<iCa<Ha<�Qa<�_a<[pa<w�a<��a<p�a<Ӱa<�a<�a<J�a<J�a<̕a<�a<�ga<�Oa<9a<V&a<)a<la<�a<�a<�(a<�<a<Ua<�na<��a<��a<9�a<s�a<H�a<��a<t�a<ݻa<��a<לa<a<�{a<�na<\ea<�`a<�aa<Qga<�qa<�a<D�a<��a<o�a<V�a<M�a<��a<W�a<��a<�a<�a<S�a<pa<eWa<�@a</a<#a<�a< a<P)a<�8a<�Ma<�ea<a<��a<ƭa<#�a<��a<��a<X�a<��a<z�a<Ϊa<v�a<L�a<�xa<�la<�da<�aa<da<qka<�va<�a<іa<�a<�a<��a<��a<��a<�a<�a<,�a<{�a<�a<ffa<�Ma<�8a<C(a</a<.a<va<�*a<�;a<�Qa<&ja<R�a<�a<��a<ܾa< �a<��a<F�a<ʽa<&�a<��a<��a<-}a<�na<�ca<X]a<\a<�_a<�ha<9ua<�a<ٕa<��a<N�a<Y�a<�a<��a<v�a<�a<םa<_�a<�la<�Ra<p:a<&a<a<�a<ra<sa< a<I2a<�Ha<�`a<?ya<~�a<��a<j�a<մa<��a<Y�a<��a<�a<9�a<oa<&^a<%Pa<�Ea<�@a<�@a<�Ea<\Oa<�\a<�la<�}a<ȍa<#�a<��a<J�a<��a<c�a<�a<�xa<m`a<�Fa<�-a<�a<>a<��`<P�`<��`<��`<a<� a<j8a<}Qa<�ia<�a<ѐa<+�a<�a<s�a<˗a<J�a<�{a<ja<�Xa<qIa<`=a<t5a<�2a<�4a<z<a<6Ha<fWa<�ha<'za<�  �  ��a<t�a<�a<R�a<k�a<�a<�wa<�^a<�Ba<�%a<�
a<��`<�`<�`<I�`<��`<�`<�`<\a<�/a<iMa<�ia<��a<��a<b�a<��a<��a<�a<�a<��a<'�a<Qya<{na<�fa<ba<ba<�ea<�ma<ya<ʆa<=�a<\�a<h�a<��a<Һa<�a<��a<��a<H�a<�oa<�Sa<8a<ja<<	a<�`<D�`<��`<]�`<�a<�!a<=a<jZa<xa<��a<(�a<Q�a<��a<��a<��a<e�a<��a<&�a<ءa<�a<��a<�a<�a<�a<��a<�a<7�a<��a<�a<�a<��a<��a<�a< �a<��a<�a<$�a<�wa<�Za<�>a<c%a<>a<ya<��`<��`<�
a<2a<�3a<�Na<�ka<w�a<�a<\�a<��a<��a<,�a<��a<X�a<~�a<*�a<��a<�a<c�a<�a<��a<E�a<7�a<p�a<u�a<�a<0�a<+�a<��a<��a<��a<��a<��a<�a<��a<ma<�Oa<-4a<0a<�	a<7�`<��`<��`<�a<�a<�8a<~Ta<Mqa<��a<�a<k�a<}�a<�a<N�a<��a<5�a<|�a<�a<W�a<��a<�a<�{a<�za<�}a<��a<��a<[�a<��a<��a<I�a< �a<��a<��a<��a<L�a<U�a</va<�Xa<5;a<�a<�a<��`<��`<@�`<'�`<�a<ca<�0a<�La<�ha<��a<��a<F�a<j�a<$�a<��a<�a<v�a<��a<-�a<Kwa<la<�ca<`_a<_a<ca<�ja<Jua<�a<�a<L�a<��a<�a<کa<V�a<g�a<�a<�ja<�Na<l1a<�a<�`<u�`<A�`<�`<��`<6�`<}�`<~a<�!a<F>a<�Za<ta<
�a<D�a<�a<B�a<��a<"�a<*�a<�}a<
pa<�ca<�Ya<{Sa<nQa<Sa<:Ya<�ba<�na<�|a<>�a<�  �  P�a<Υa<��a<ޡa<��a<ׄa<.ma<�Pa<�1a<a<�`<�`<L�`<V�`<=�`<�`<��`<��`<t�`<�a<e=a<�\a<�xa<*�a<I�a<��a<C�a<��a<�a<�a<S�a<��a<Q�a</a<�{a<�{a<Ba<��a<��a<Y�a<��a<}�a<��a<μa<��a<X�a<��a<}�a<�}a<aa<1Ba<R#a<a<��`<��`<S�`<��`<%�`<��`<`
a<�'a<dHa<ia<Ƈa<��a<�a<��a<m�a<��a<��a<��a<U�a<�a<L�a<�a<A�a<y�a<ޙa<��a<�a<�a<'�a<��a<��a<[�a<��a<��a<h�a<��a<��a<��a<�ga<Ha<�(a<;a<��`<�`<��`<3�`<��`<a<�a<�:a<�Za<nza<W�a<�a<��a<��a<��a<��a<��a<r�a<O�a<ϲa<>�a<��a<w�a<��a<��a<��a<ԧa<�a<i�a<��a<��a<�a<��a<j�a<��a<��a<��a<�{a<b\a<*<a<�a<=a<��`<�`<��`<�`<�`<�a<�"a<fAa<Baa<�a<z�a<��a<_�a<Y�a<��a<��a<��a<��a<�a<��a<��a<��a<|�a<��a<��a<u�a<^�a<�a<(�a<��a<��a<Z�a<��a<	�a<��a<!�a<օa<�ga<�Fa<k&a<{a<A�`<��`<��`<A�`<��`<��`<��`<�a<}:a<�Ya<�va<�a<ڣa<z�a<��a<��a<<�a<0�a<��a<e�a<��a<��a<�|a<Bya<�xa<�{a<ȁa<��a<��a<x�a<3�a<,�a<�a<��a<��a<H�a<�ya<6^a<&?a<�a<�`<��`<$�`<Ѽ`<�`<5�`<J�`<O�`<��`<va<=-a<�La<?ia<��a<	�a<�a<��a<u�a<{�a<�a<��a<Q�a<�ya<ra<ma<Qka<�la<�qa<ya<��a<%�a<��a<�  �  R�a</�a<K�a<	�a<1�a< a<�da<Fa<�$a<ua<t�`<��`<��`<�`<Y�`<ʧ`<%�`<��`<?�`<�a<�0a<�Ra<Cqa<�a<��a<��a<|�a<��a<%�a<��a<D�a< �a<h�a<Ǒa<��a<��a<i�a<��a<�a<h�a<q�a<f�a<�a<F�a<U�a<��a<U�a<͏a<�ta<kUa<4a<
a<��`<��`<��`<��`<�`<�`<��`<��`<ma<	:a<%]a<l~a<��a<q�a<�a<��a<��a<u�a<Y�a<��a<��a<Z�a<��a<F�a<�a<{�a<=�a<T�a<�a<X�a<Y�a<��a<��a<X�a<��a<��a<��a<5�a<�|a<�[a<'9a<�a<\�`<��`<��`<��`<��`<��`<k�`<�
a<�*a<SMa<Poa<َa<ɩa<�a<��a<��a<��a<q�a<�a<��a<g�a<ݹa<��a<ݯa<?�a<n�a<زa<��a<�a<��a<f�a<��a<y�a<8�a<��a<[�a<Ūa<N�a<
qa<&Oa<�,a<a<��`<N�`<�`<��`<��`<��`<q�`<ka<;2a<�Ta<�ua<��a<��a<��a<�a<'�a<��a<d�a<�a<�a<�a<��a<5�a<�a<A�a<'�a<?�a<��a<��a<��a<��a< �a<��a<}�a<n�a<��a<t�a<�|a<�[a<�8a<$a<A�`<X�`<��`<�`<��`<��`<��`<V�`<'a<!,a<�Ma<Zma<�a<b�a<��a<	�a<��a<�a<εa<�a<+�a<��a<$�a<ُa<ٌa<��a<��a<�a<��a<Ӡa<B�a</�a<t�a<��a<p�a<*�a<F�a<fra<=Ta<�2a<�a<�`<�`<ѷ`<��`<-�`<��`<��`<��`<��`<��`<�a<xAa<�`a<u{a<c�a<�a<�a<��a<2�a<��a<�a<�a<U�a<%�a<i�a<�~a<7�a<σa<щa<b�a<��a<m�a<�  �  ��a<۬a<X�a<S�a<Ґa< {a<V_a<1?a<a<��`<)�`<[�`<z�`<!�`<��`<�`<8�`<~�`<Q�`<+a<�(a<�Ka<�ka<>�a<t�a<P�a<Գa<�a<˵a<ʱa<C�a<q�a<J�a<z�a<��a<ʛa<W�a<Ţa<�a<	�a<i�a<��a<��a<Z�a<ӽa<e�a<{�a<?�a<�na<�Ma<'+a<�a<(�`<�`<k�`<ٲ`<-�`<|�`<�`< �`<�a<�0a<�Ua<?xa<�a<n�a<��a<$�a<��a<�a<x�a<��a<W�a<<�a<�a<-�a<D�a<��a<	�a<^�a<�a<��a<��a<��a<��a<��a<��a<�a<�a<�a<va<�Sa<�/a<'a<O�`<��`<�`<��`<��`<��`<��`<}�`<� a<�Da<=ha<�a<��a<b�a<��a<��a<!�a<��a<��a<��a<]�a<;�a<#�a<�a<y�a<z�a<h�a<0�a<�a<��a<G�a<J�a<'�a<F�a<��a<��a<Ŧa<��a<$ja<�Fa<�"a<� a<��`< �`<B�`<!�`<�`<��`<K�`<za<�(a<eLa<oa<o�a<�a<��a<��a<}�a< �a<	�a<O�a<�a<x�a<��a<�a<-�a<y�a<�a<��a<��a<��a<��a<��a<��a<��a<��a<�a<��a<�a<�va<nTa<�/a<�a<��`<��`<a�`<�`<��`<F�`<�`<��`<� a<#a<
Fa<-ga<\�a<^�a<�a<M�a<��a<��a<�a<�a<��a<��a<X�a<��a<
�a<��a<`�a<�a<+�a<�a<��a<�a<��a<�a<N�a<A�a<ևa<Dma<�Ma<�*a<ja<X�`<�`<��`<�`<`�`<�`<:�`<R�`<~�`<��`<a<e:a<�Za<Awa<Սa<#�a<�a<�a<X�a<[�a<{�a<ؚa<��a<��a<k�a<�a<@�a<\�a<\�a<��a<:�a<L�a<�  �  ��a<8�a<y�a<o�a<ßa<��a<2]a<�1a<�a< �`<��`<F{`<�\`<SJ`<�E`<N`<]d`<��`<�`<��`<�a<�@a<Lla<͐a<��a<h�a<i�a<��a<��a<<�a<D�a<��a<0�a<3�a<U�a<��a<�a<��a<	�a<��a<��a<��a<�a<��a<��a<\�a<��a<��a<Oia<�<a<�a<��`<ñ`<��`<qs`<?f`<f`<�s`<ˎ`<ĳ`<��`<�a<RCa</ra<қa<��a<��a<v�a<��a<�a<~�a<��a<(�a<M�a<��a<��a<��a<:�a<��a<�a<��a<*�a<��a<R�a<K�a</�a<��a<��a<,�a<-�a<ma<>a<Fa<��`<D�`<x�`<>z`<�p`<�t`<�`<��`<��`<��`<r)a<�Ya<o�a<'�a<d�a<;�a<~�a<3�a<G�a<�a<��a<��a<��a<��a<(�a<�a<��a<��a<��a<$�a<A�a<��a<��a<B�a<�a<��a<��a<)�a<:�a<']a<�,a<��`<G�`<�`<@�`<s`<n`<�u`<k�`<�`<��`<�a<f5a<�da<R�a<�a<\�a<T�a<��a<?�a<��a<`�a<��a<_�a< �a<Z�a<��a<�a<��a<5�a<��a<9�a<��a<��a<��a<��a<k�a<��a<w�a<��a<�qa<�Ca<a<��`<Q�`<e�`<iq`<jb`<�``<�l`<��`<Ψ`<�`<Na<C3a<`a<��a<̨a<z�a<��a<��a<��a<�a<F�a<��a<��a<=�a<p�a<�a<d�a<�a<�a<F�a<��a<�a<��a<r�a<��a<ȿa<(�a<D�a<�na<Da<�a<L�`<M�`<O�`<f`<`N`<�D`<�G`<�X`<4v`<�`<��`<"�`<X+a<�Wa<~a<�a<��a<¾a<G�a<1�a<ڿa<q�a<&�a<k�a<,�a<ɢa<͡a<��a<�a<�a<��a<&�a<ſa<�  �  ��a<u�a<7�a<�a<�a<��a<�_a<�4a<�a<��`<M�`<��`<c`<�P`<�K`<hT`<Xj`<?�`<��`<��`<a<FDa<�na<��a<�a<��a<�a<��a<��a<��a<��a<y�a<z�a<�a<�a<N�a<ٯa<Ĵa<��a<��a<��a<f�a<��a<F�a<��a<;�a<0�a<��a<Ola<v@a<,a<O�`<:�`<o�`<�y`<Ol`<�l`<Pz`<��`<D�`<��`<�a<)Ga<Dua<�a<�a<��a<q�a<]�a<��a<4�a<��a<C�a<�a<��a<��a<��a<��a<i�a<C�a<��a<]�a<�a<:�a<-�a<��a<��a<��a<׻a<��a<Mpa<Ba<�a<��`<ڸ`<a�`<��`<�v`<�z`<*�`<S�`<�`<T�`<�-a<w]a<D�a<
�a<��a<��a<D�a<��a<��a<��a<R�a<��a<`�a<��a<��a<��a<��a<��a<2�a<�a<��a<��a<1�a<~�a<��a<1�a<��a<	�a<��a<�`a<�0a<i a<��`<ɪ`<`�`<jy`<�s`<|`<h�`<��`<��`<	a<x9a< ha<ϑa<�a<��a<��a<R�a<@�a<��a<��a<��a<+�a<j�a<:�a<_�a<��a<\�a<J�a<*�a<D�a<��a<S�a<F�a<��a<S�a<��a<�a<��a<�ta<AGa<>a<��`<ȸ`<3�`<�w`<zh`<�f`<�r`<m�`<N�`<��`<�a<7a<�ca<��a<P�a<o�a<��a<a�a<��a<��a<9�a<��a<h�a<]�a<E�a<��a<�a<�a<"�a<�a<�a<2�a<��a<T�a<~�a<�a<J�a<�a<qa<YGa<�a<��`<U�`<�`<�k`<�T`<�J`<N`<_`<�{`<b�`<M�`<N�`<�.a<nZa<�a<k�a<R�a<��a<��a<��a<Z�a<��a<�a<�a<)�a<��a<h�a<t�a<ՠa<��a<��a<��a<5�a<�  �  ��a<��a<��a<��a<��a<5�a<�ga<[>a<Na<�`<��`<ő`<�t`<�c`<�^`<?g`<�{`<ԛ`< �`<��`< a<CMa<va<��a<1�a<��a<�a<c�a<�a<��a<Y�a<E�a<K�a<�a<��a<��a<؟a<ԥa<��a<��a<��a<��a<7�a<X�a<��a<��a<~�a<�a<�ta<~Ja<Ka<c�`<D�`<��`<"�`<H`<s`<ٌ`<�`<s�`<��`<B"a<lQa<�}a<z�a<��a<7�a<��a<��a<��a<��a<=�a<S�a<�a<�a<��a<�a<^�a<��a<��a<Q�a<��a<�a<<�a<��a<��a<��a<��a<��a<��a<ya<�La<Xa<��`<Z�`<�`<l�`<؉`<��`<D�`<>�`<��`<�
a<_9a<ga<#�a<�a<��a<��a<��a<�a<��a<��a<��a<��a<��a<Z�a<��a<׻a<D�a<f�a<b�a<@�a<�a<��a<��a<��a<N�a<��a<��a<��a<��a<�ia<�<a<�a<�`<��`<T�`<^�`<�`<�`<�`<F�`<��`<	a<�Da<qa<�a<�a<��a<��a<T�a<��a<��a<��a<��a<��a<;�a<��a<�a<�a<Z�a<X�a<�a<�a<��a<��a<��a<��a<a�a<��a<8�a<�a<}a<HQa<]"a<��`<��`<\�`<�`<r{`<�y`<m�`<��`<~�`</�`<�a<^Aa<�ka<8�a<Үa<��a<�a<��a<R�a<Y�a<��a<��a<w�a<��a<W�a<ՙa<��a<;�a<��a<��a<��a<3�a<��a<��a<C�a<��a<Q�a<ۘa<xa<%Pa<e#a<Z�`< �`<`�`<s}`<�g`<�]`<a`<3q`<Ռ`<�`<��`<a<y8a<Mba<ͅa<M�a<"�a<0�a< �a<��a<L�a<��a<��a<Z�a<�a<e�a<��a<+�a<~�a<��a<ۡa<��a<�a<�  �  ��a<��a<T�a<n�a<٩a<��a<2sa<(Ma<Y#a<0�`<t�`</�`<,�`<ŀ`<Z|`<8�`<ؗ`<��`<)�`<�a<`1a<W[a<��a<W�a<��a<��a<��a<��a<Ƚa<��a<��a<#�a<��a<�a<��a<c�a<�a<+�a<�a<�a<�a<��a<��a<h�a<��a<~�a<��a<��a<0�a<ZZa<�0a<ma<��`<��`<��`<М`<�`<j�`<;�`<c�`<.
a<�5a<�aa<��a<s�a<%�a<��a<��a<�a<��a<8�a<��a<x�a<�a<��a<��a<ʠa<M�a<�a<߭a<Ӹa<��a<e�a<��a<e�a<��a<��a<��a<�a<7�a<Ԇa<�]a<�2a<�a<��`<��`<G�`<��`<�`<��`<��`<��`<l a<�Ka<2va<�a<��a<�a<��a<�a<P�a<u�a<��a<]�a<ҿa<��a<E�a<�a<��a<{�a<�a<�a<нa<�a<S�a<a�a<��a<��a<��a<��a<	�a<>�a<�xa<�Na<�"a<��`<	�`<��`<��`<��`<�`<�`<(�`<� a<�*a<�Ua<a<�a<��a<9�a<��a<)�a<*�a<��a<��a<�a<Եa<p�a<�a<�a<Лa<��a<��a<��a<ֻa<�a<��a<h�a<��a<G�a<��a<f�a<��a<��a<"aa<�5a<�	a<v�`<x�`<��`<��`<l�`<��`<�`<o�`<~�`<�'a<�Qa<�xa<4�a<`�a<J�a<Y�a<&�a<R�a<��a<>�a<ޤa<Q�a<+�a<0�a<�a<za<q�a<��a<�a<��a<��a<3�a<��a<��a<��a<Z�a<�a<��a<�]a<W4a<�a<��`<�`<(�`<^�`<8{`<_~`<�`<��`<�`<a�`<�a<�Ga<@na<��a<Ȧa<k�a<L�a<l�a<h�a<k�a<�a<v�a<K�a<�ya<�sa<fqa<isa<>ya<f�a<p�a<�a<��a<�  �  �a<2�a<`�a<ùa<��a<e�a<:�a<�_a<�9a<�a<��`<��`<��`<��`<Ţ`<ȩ`<̻`<��`<��`<Ma<�Fa<�la<��a<N�a<T�a<b�a<��a<)�a<��a<�a<C�a<f~a<!pa<�ea<�_a<�_a<rda<�na<�|a<9�a<�a<r�a<r�a<��a<�a<M�a<��a<��a<��a<,na<fHa<q"a<l�`<��`<��`<��`<O�`<��`<f�`<Ka<�&a<8Na<�ua<��a<�a<��a<��a<��a<��a<��a<p�a<@�a<��a<ߙa<H�a<��a<~a<�~a<v�a<!�a<��a<��a<��a<��a<z�a<��a<��a<	�a<��a<��a<�a<sa<�Ka<�%a<�a<_�`<��`<��`<�`<9�`<�`<�a<�;a<�ba<#�a<��a<��a<=�a<��a<��a<Y�a<	�a<�a<[�a<��a<{�a<��a<��a<�~a<��a<��a<q�a<�a<��a<L�a<n�a<4�a<�a<�a<f�a<��a<H�a<E�a<ea<�=a<&a<��`<��`<|�`<�`<��`<��`<5�`<�a<|Da<rka<��a<�a<��a< �a<Z�a<=�a<��a<��a<��a<��a<�a<�a<܀a<Gza<ya<�|a<�a<�a<��a<�a<V�a<�a<��a<��a<��a<}�a<��a<0�a<�ta<tMa<�%a<� a<R�`<��`<�`<��`<&�`<4�`<W�`<�a<�?a<�ea<�a<��a<�a<��a<Y�a<��a<s�a<�a<��a<�a<O{a<�la<Kba<�\a<�\a<�aa<la<�ya<��a<�a<��a<��a<5�a<��a<��a<��a<B�a<�na<yIa<�!a</�`<��`<�`<ϩ`<��`<Q�`<�`<��`<��`<�a<f4a<�Za<�|a<˘a<�a<:�a<Һa<z�a<�a<�a<�a<7va< fa<�Ya<lQa<�Na<�Pa<�Xa<�da<�ta<��a<��a<�  �  ��a<6�a<��a<��a<Ӵa<}�a<$�a<�sa<�Ra<	1a<�a<[�`<��`<��`<b�`<��`<|�`<h�`<�a<8<a<�^a<�a<ƛa<[�a<u�a<h�a<�a<�a<�a<��a<�sa<f^a<La<�>a<7a<p6a<M<a<�Ha<�Za<�pa<��a<i�a<��a<O�a<��a<9�a<��a<+�a<r�a<݃a<ca<@Ba<�#a<�	a<��`<k�`<��`<��`<a<�&a<�Fa<\ia<&�a<��a<�a<-�a<?�a<@�a<�a<��a<�a<��a<��a<^xa<ga<�Za<�Ta<�Ua<]a<�ja<-}a<�a<W�a<��a<��a<*�a<��a<��a<-�a<�a<K�a<h�a<[ha<(Ga<�(a<�a<~ a<��`<_�`<�a<�a<�9a<IZa<M|a<��a<�a<v�a<�a<��a<4�a<��a<&�a<�a<Ԟa<�a<�sa<�ca</Ya<�Ua<PXa<�aa<&qa<�a<��a<��a<��a<4�a<-�a<7�a<��a<��a<4�a<E�a<~a<�[a<�:a<Da<;a<��`<��`<v�`<�a<�"a<�@a<paa<f�a<��a<�a<��a<(�a<e�a<Y�a<x�a<�a<��a<h�a<{a<�ga<�Ya<dQa<�Oa<�Ta<p`a<qa<��a<Ϝa<I�a<O�a<~�a<��a<x�a<l�a<D�a<�a<��a<ha<�Ea<%a<�	a<��`<��`<8�`<y�`<�a<�a<C:a<�Za<|a<R�a<ղa<m�a<
�a<��a<-�a<Y�a<��a<
�a<pa<�Ya<�Ga<Z:a<�3a<�3a<�:a<�Ga<zYa<�na<��a<O�a<��a<úa<�a<+�a<2�a<�a<A�a<�`a<F>a<�a<��`<E�`<��`<<�`<��`<��`<]�`<a<7,a<�Ma<oa<I�a<f�a<Ȳa<�a<��a<�a<&�a<ʅa<�na<�Wa<FCa<U3a<�(a<b%a<P(a<2a<�Aa<�Ua<~la<Ӄa<�  �  ��a<��a<��a<��a<s�a<��a<��a<��a<~la<�Oa<Q4a<�a<o
a<]�`<b�`<�a<xa<�#a<7=a<�Ya<Rwa<�a<�a<,�a<�a<Ϳa<�a<J�a<݌a<�qa<aUa<�:a<J$a<�a<E
a<$	a<na<�a<,5a<�Oa<&ma<��a<��a<��a<��a<}�a<�a<'�a<��a<ҙa<�~a<�ba<�Ha<s3a<&$a<Ma<�a<�%a<	6a<�La<�ga<p�a<��a<ؼa<��a<$�a<�a<��a<�a<�a<�a<��a<?ma<ISa<>a</a<�'a<�(a<�1a<vBa<Ya<�sa<Ȑa<۬a<k�a<i�a<��a<��a<b�a<��a<k�a<C�a<��a<>ia<�Oa<~;a<�-a<�'a<*a<�4a<�Fa< ^a<�ya<��a<c�a<<�a<+�a<?�a<��a<��a<�a<��a<�a<�a<�ea<Ma<�9a<�,a<(a<�+a<�7a<;Ja<^ba<~a<�a<��a<��a<D�a<��a<N�a<�a<��a<T�a<×a<�za<�^a<�Fa<�3a<O(a<�$a<�)a<�6a<MJa<(ca</a<�a<]�a<E�a<��a<��a<��a<:�a<��a<��a<ԏa<�ra<�Wa<4@a<�.a<�$a<�"a<�(a<7a<�Ka<ea<A�a<��a<.�a<��a<|�a<��a<��a<<�a<)�a<��a<��a<�ea<aJa<43a<"a<va<(a<)a<�,a<�Aa<.[a<wa<��a<1�a<m�a<h�a<��a<?�a<$�a<�a<�a<&ma<�Oa<�4a<�a<�a<�a<�a<ha<]a<d5a<�Oa<�ka<�a<��a<��a<�a<-�a<`�a<A�a<Y�a<�xa<v[a<�>a<�$a<�a<�a<:�`<K�`<�a<
a<R0a<~Ka<Dha<ȃa<e�a<�a<��a<$�a<G�a<>�a<ĉa<�na<�Qa<�5a<�a<Y	a<��`<��`<��`<�a<�a<3a<Oa<9la<�  �  �sa<��a<�a<)�a<4�a<¶a<j�a<��a<j�a<uma<Wa<�Ca<�4a<�+a<�)a<.a<J9a<�Ia<�^a<bva<�a<��a<��a<�a<��a<Q�a<�a<�a<�wa<Wa<�5a<Ea<c�`<��`<��`<+�`<r�`<#�`<�a<.a<:Pa<;sa<ޓa</�a<��a<��a<��a<=�a<9�a<�a<h�a<�a</ma<�[a<fOa<]Ia<�Ia<Qa<�^a<pqa<�a<��a<r�a<��a<\�a<:�a<��a<��a<(�a<�a<��a<Cma<	La<6-a<�a<3a<��`<��`<�a<!a< 4a<�Sa<�ua<:�a<t�a<��a<��a<��a<��a<��a<��a<K�a<t�a<q�a<�ua<ea<�Ya<Ua<�Va<�_a< na<r�a<�a<8�a<K�a<��a<��a<��a<��a<��a<d�a<��a<�a<da<Ca<�%a<la<|�`<�`<F�`<a<2"a<�>a<�_a<{�a<4�a<z�a<�a<c�a<�a<:�a<��a<��a<��a<T�a<��a<�ma<b^a<�Ta<5Ra<�Ua<�`a<�pa<�a<��a<��a<x�a<��a<��a<_�a<Z�a<5�a<}�a<��a<7ua<BSa<�2a<Ka<�a<��`<��`<��`<�a<�$a<HCa<Pda<�a<e�a<U�a<��a<��a<B�a<P�a<��a<��a<q�a<d�a<�na<�[a<[Ma<�Ea<TDa<�Ia<�Ua<fa<={a<��a<k�a<Q�a<&�a<��a<��a<��a<?�a<��a<�sa<�Pa<�.a<�a<�`<��`<��`<��`<�`<
�`<Oa<�/a<�Pa<�qa<��a<Q�a<̷a<3�a<��a<6�a<ǣa<��a<Nwa<�_a<uJa<l9a<�-a<�(a<
*a<R2a<�@a<�Sa<�ia<ۀa<��a<��a<�a<M�a<Q�a<$�a<��a<�va<Va<�3a<�a<O�`<4�`<S�`<��`<\�`<L�`<��`<�a<�0a<�Ra<�  �  2`a<�a<�a<(�a<I�a<ٻa<��a<��a<w�a<ۇa<fva<&ga<�[a<�Ta<Sa<�Va<g_a<�la<<}a<��a<ѡa<!�a<��a<$�a<��a<2�a<�a<�a<ca<:=a<�a<��`<��`<�`<0�`<��`<Ҹ`<��`<y�`<�a<34a<!\a<a<<�a<��a<{�a<q�a<��a<j�a<��a</�a<F�a<�a<��a<�va<\ra<sa<�xa<Ճa<��a<��a<[�a<��a<��a<��a<��a<,�a<��a<��a<M�a<mxa<�Qa<d+a<ua<�`<��`<�`<U�`<��`<��`<a<P4a<8[a<Ӂa<�a<g�a<�a<�a<F�a<M�a<��a<��a<�a<K�a<ӗa<Њa<�a<B~a<�a<��a<�a<<�a<�a<��a<��a<�a<��a<8�a<T�a<r�a<K�a<r�a<�ma<�Fa<� a<��`<��`<x�`<d�`<�`<��`<��`<Ja<�Aa<�ha<|�a<دa<��a<a�a<#�a<S�a<��a<e�a<��a<��a<ݠa<)�a<+�a<�}a<�{a<l~a<��a<:�a<C�a<�a<x�a<�a<��a<��a<M�a<@�a<]�a<��a<�a<e[a<P4a<~a<m�`<�`<p�`<��`<=�`<U�`<��`< "a<EHa<�na<D�a<^�a<M�a<��a<�a<�a<��a<>�a<6�a<��a<q�a<?�a<�ta<�na<ima<{qa<�za<��a< �a<��a<��a<�a<r�a<��a< �a<8�a<֡a<$�a<]a<X5a<�a<��`<��`<��`<�`<��`<�`<��`<l�`<a<e6a<t\a<$a<��a< �a<��a<7�a<��a<űa<��a<ݏa<�}a<�la<,_a<�Ua<�Qa<�Ra<\Ya<vda<dsa<Ȅa<y�a<�a<��a<��a<��a<�a<՞a<��a<�ca<�=a<�a<��`<i�`<`�`<Y�`<_�`<?�`<1�`<q�`<�`<�a<:a<�  �  �Ma<ta<w�a<��a</�a<�a<f�a<�a<��a<��a<j�a<�a<Y|a<wa<�ua<�xa<�a<��a<<�a<L�a<�a<F�a<o�a<`�a<y�a<ˮa<��a<Lva<�Oa<&a<{�`<��`<3�`</�`<1�`<-�`<s�`<Q�`<�`<��`<%a<9Ga<�pa<��a<M�a<{�a<��a<��a<��a<k�a<�a<c�a<I�a<d�a<��a<�a<Õa<��a<	�a<z�a<:�a<��a<�a<`�a<��a<`�a<��a<��a<��a<�a<�ca<=9a<�a<W�`<��`<��`<˧`<:�`<��`<?�`<��`<�a<�Ca<=na<ŕa<��a<C�a<��a<�a<~�a<��a<K�a<S�a<��a<z�a<��a<�a<
�a<[�a<��a<6�a<��a<�a<��a<k�a<��a<O�a<��a<Q�a<@�a<�a<��a<Xa<�,a<a<]�`<r�`<̮`<�`<K�`<��`<P�`<�`<0'a<yRa<:|a<�a<�a<��a<	�a<��a<��a<��a<�a<u�a<�a<��a<�a<-�a<J�a<��a<ݦa<>�a<L�a<��a<��a<?�a<��a<��a<F�a<��a<��a<�a<�na<FDa<�a<��`<�`<E�`<n�`<��`<۫`<��`<`�`<a<3/a<Za<v�a<�a<��a<��a<_�a<��a<��a<'�a<�a<��a<Ϊa<"�a<��a<;�a<!�a<J�a<ڙa<��a<��a<K�a<�a<��a<��a<��a<}�a<f�a<�a<�qa<�Ha<�a<?�`<��`<M�`<G�`<ņ`<y�`<1�`<+�`<�`<<�`<�a<�Ha<�oa<!�a<D�a< �a<��a<��a<g�a<��a<�a<!�a<D�a<�~a<�wa<�ta<uua<^za<��a<�a<��a<C�a<ͳa<ݻa<C�a<S�a<�a<��a<Bwa<�Qa<(a<��`<��`<4�`<M�`<�~`<�w`<s}`<�`<ߪ`<��`<I�`<�#a<�  �  U?a<�ha<H�a<åa<n�a<��a<��a<��a<B�a<��a<�a<Z�a<��a<�a<��a<X�a<y�a<p�a<�a<��a<��a<8�a<��a<�a<�a<#�a<��a<+ja<�@a<ra<��`<��`<d�`<�|`<�m`<�k`<�v`<��`<��`<%�`< a<u6a<sca<��a<8�a<��a<��a<~�a<��a<T�a<��a<��a<��a<��a<o�a<&�a<�a<��a<X�a<x�a<��a<��a<k�a<*�a<�a<��a<%�a<4�a<Ҥa<�~a<�Sa<g%a<O�`<>�`<@�`<��`<'�`<��`<3�`<:�`<K�`<�a<�0a<�^a<N�a<2�a<B�a<��a<R�a<��a<)�a<��a<Y�a<L�a<�a<l�a<~�a<C�a<L�a<(�a<��a<��a<��a<��a<��a<K�a<D�a<$�a<��a<m�a<ߛa<bsa<�Fa<�a<��`<W�`<x�`<��`<5�`<�`<r�`< �`<}�`<&a<�@a<�ma<��a<ڸa<��a<H�a<�a<��a<X�a<��a<��a<��a<j�a<F�a<�a<��a<R�a<ھa</�a<*�a<�a<c�a<7�a<6�a<��a<��a<:�a<��a<Ήa<t_a<�1a<Ja<^�`<I�`<�`<	�`<ل`<�`<�`<��`<_�`<a<@Ia<�ta<��a<�a<��a<��a<��a<\�a<�a<��a<��a<y�a<=�a<c�a<O�a<B�a<V�a<)�a<��a<6�a<��a<j�a<��a<��a<;�a<��a<��a<�a<�da<18a<�a<��`<Ű`<ލ`<�u`<$i`<�i`<�w`<'�`<��`<U�`<�a</9a<aca<��a<@�a<4�a<9�a< �a<��a<ռa<�a<��a<��a<��a<\�a<��a<a�a<�a<R�a<١a<p�a<7�a<�a<t�a<9�a<�a<V�a<؍a<#la<�Ca<�a<��`<��`<4�`<Yu`<�a`<?Z`<L``<�r`<��`<S�`<C�`<a<�  �  6a< aa<ƅa</�a<��a<A�a<��a<�a<��a<o�a<�a<@�a<�a<D�a< a<}�a<��a<�a<��a<�a<��a<�a<H�a<K�a<�a<'�a<��a<3ba<�6a<�a<%�`<�`<l�`<�j`<�Z`<�X`<�c`<B|`<5�`<v�`<b�`<�+a<�Za<��a<h�a<��a<L�a<��a<��a<m�a<��a<0�a<��a<��a<.�a<��a<��a<��a<�a<I�a<��a<H�a<��a<4�a<��a<��a<y�a<��a<"�a<Pva<Ia<�a<��`<��`<�`<C�`<9w`<�x`<��`< �`<W�`<��`<�$a<�Ta<)�a<��a<�a<��a<`�a<��a<��a<E�a<U�a<��a<b�a<t�a<��a<�a<��a<��a<��a<��a<��a<I�a<-�a<x�a<(�a<��a<a�a<#�a<��a<Kja<k;a<�
a<��`<��`<`<�~`<Hw`<.}`<��`<=�`<+�`<�a<15a<Pda<
�a<W�a<e�a<��a<��a<��a<��a<�a<a�a<g�a<S�a<��a<]�a<R�a<{�a<�a<��a<��a<Q�a<V�a<�a<��a<��a<��a<@�a<
�a<؁a<�Ua<�%a<��`<��`<O�`<��`<u`<�q`<\|`<��`<��`<��`<ka<�>a<;la<��a<�a<��a<��a<��a< �a<'�a<��a<w�a<�a<��a<!�a<�a<�a<5�a<׿a<[�a<�a<��a<��a<��a<z�a<��a<S�a<�a<D�a</\a<�-a<��`<a�`<��`<�|`<c`<7V`<W`<se`<�`<��`<`�`<��`<D/a<;[a<��a<�a<�a<E�a<�a<��a<��a<�a<׳a<#�a<��a<i�a<w�a<͟a<n�a<h�a<�a<{�a<�a<��a<��a<�a<��a<��a<��a<�da<p:a<ta<��`<}�`<��`<�c`<�N`<VG`<aM`<�``<�`<�`<�`<�a<�  �  �2a<r^a<�a<�a<��a<��a<Y�a<��a<M�a<	�a<�a<߭a<*�a<��a<&�a<��a<��a<Z�a<��a<F�a<�a<��a<��a<}�a<e�a<ȣa<ąa<T_a<?3a<ha<��`<��`<��`<}d`<�T`<�R`<�]`<`v`<��`<x�`<�`<�'a<�Wa<O�a<ƥa<��a<.�a<-�a<��a<��a<��a<�a<��a<��a<X�a<�a<��a<��a<��a<��a<��a<E�a<��a<x�a<�a<��a<z�a<�a<��a<.sa<9Ea<�a<��`<q�`<�`<�|`<9q`<�r`<��`<Z�`<��`<��`<T a<�Pa<3~a<
�a<��a<��a<��a<=�a<?�a<��a<��a<��a<��a<c�a<��a<b�a< �a<��a<��a< �a<V�a<��a<�a<g�a<w�a<��a<$�a<V�a<��a<�fa<Q7a<sa<k�`<�`<��`<~x`<Xq`<�v`<w�`<��`<��`<a a<1a<�`a<[�a<}�a<�a<h�a<�a<w�a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<�a<��a<��a<��a<��a<4�a<�a<:�a<��a<#�a<�~a<)Ra<�!a<��`<7�`<��`<�`<�n`<�k`<�u`<č`<��`<��`<
a<�:a<�ha<i�a<q�a<��a<��a<7�a<J�a<K�a<��a<H�a<F�a<��a<K�a<:�a<D�a<b�a<��a<��a<��a<��a<��a<��a<��a<��a<T�a<��a<�a<Ya<�)a<E�`<{�`<��`<�v`<�\`<8P`<�P`<._`<Hz`<8�`<��`<�`<�+a<EXa<�a<��a<8�a<d�a<��a<�a<��a<V�a<շa<��a<��a<��a<Ԥa<�a<��a<�a<�a<0�a<��a<v�a<��a<m�a<k�a<��a<Ća<Aba<7a<[a<h�`<R�`<�}`<�]`<tH`<hA`<G`<�Z`<'z`<��`<��`<za<�  �  6a< aa<ƅa</�a<��a<A�a<��a<�a<��a<o�a<�a<@�a<�a<D�a< a<}�a<��a<�a<��a<�a<��a<�a<H�a<K�a<�a<'�a<��a<3ba<�6a<�a<%�`<�`<l�`<�j`<�Z`<�X`<�c`<B|`<5�`<v�`<b�`<�+a<�Za<��a<h�a<��a<L�a<��a<��a<m�a<��a<0�a<��a<��a<.�a<��a<��a<��a<�a<I�a<��a<H�a<��a<4�a<��a<��a<y�a<��a<"�a<Pva<Ia<�a<��`<��`<�`<C�`<9w`<�x`<��`< �`<W�`<��`<�$a<�Ta<)�a<��a<�a<��a<`�a<��a<��a<E�a<U�a<��a<b�a<t�a<��a<�a<��a<��a<��a<��a<��a<I�a<-�a<x�a<(�a<��a<a�a<#�a<��a<Kja<k;a<�
a<��`<��`<`<�~`<Hw`<.}`<��`<=�`<+�`<�a<15a<Pda<
�a<W�a<e�a<��a<��a<��a<��a<�a<a�a<g�a<S�a<��a<]�a<R�a<{�a<�a<��a<��a<Q�a<V�a<�a<��a<��a<��a<@�a<
�a<؁a<�Ua<�%a<��`<��`<O�`<��`<u`<�q`<\|`<��`<��`<��`<ka<�>a<;la<��a<�a<��a<��a<��a< �a<'�a<��a<w�a<�a<��a<!�a<�a<�a<5�a<׿a<[�a<�a<��a<��a<��a<z�a<��a<S�a<�a<D�a</\a<�-a<��`<a�`<��`<�|`<c`<7V`<W`<se`<�`<��`<`�`<��`<D/a<;[a<��a<�a<�a<E�a<�a<��a<��a<�a<׳a<#�a<��a<i�a<w�a<͟a<n�a<h�a<�a<{�a<�a<��a<��a<�a<��a<��a<��a<�da<p:a<ta<��`<}�`<��`<�c`<�N`<VG`<aM`<�``<�`<�`<�`<�a<�  �  U?a<�ha<H�a<åa<n�a<��a<��a<��a<B�a<��a<�a<Z�a<��a<�a<��a<X�a<y�a<p�a<�a<��a<��a<8�a<��a<�a<�a<#�a<��a<+ja<�@a<ra<��`<��`<d�`<�|`<�m`<�k`<�v`<��`<��`<%�`< a<u6a<sca<��a<8�a<��a<��a<~�a<��a<T�a<��a<��a<��a<��a<o�a<&�a<�a<��a<X�a<x�a<��a<��a<k�a<*�a<�a<��a<%�a<4�a<Ҥa<�~a<�Sa<g%a<O�`<>�`<@�`<��`<'�`<��`<3�`<:�`<K�`<�a<�0a<�^a<N�a<2�a<B�a<��a<R�a<��a<)�a<��a<Y�a<L�a<�a<l�a<~�a<C�a<L�a<(�a<��a<��a<��a<��a<��a<K�a<D�a<$�a<��a<m�a<ߛa<bsa<�Fa<�a<��`<W�`<x�`<��`<5�`<�`<r�`< �`<}�`<&a<�@a<�ma<��a<ڸa<��a<H�a<�a<��a<X�a<��a<��a<��a<j�a<F�a<�a<��a<R�a<ھa</�a<*�a<�a<c�a<7�a<6�a<��a<��a<:�a<��a<Ήa<t_a<�1a<Ja<^�`<I�`<�`<	�`<ل`<�`<�`<��`<_�`<a<@Ia<�ta<��a<�a<��a<��a<��a<\�a<�a<��a<��a<y�a<=�a<c�a<O�a<B�a<V�a<)�a<��a<6�a<��a<j�a<��a<��a<;�a<��a<��a<�a<�da<18a<�a<��`<Ű`<ލ`<�u`<$i`<�i`<�w`<'�`<��`<U�`<�a</9a<aca<��a<@�a<4�a<9�a< �a<��a<ռa<�a<��a<��a<��a<\�a<��a<a�a<�a<R�a<١a<p�a<7�a<�a<t�a<9�a<�a<V�a<؍a<#la<�Ca<�a<��`<��`<4�`<Yu`<�a`<?Z`<L``<�r`<��`<S�`<C�`<a<�  �  �Ma<ta<w�a<��a</�a<�a<f�a<�a<��a<��a<j�a<�a<Y|a<wa<�ua<�xa<�a<��a<<�a<L�a<�a<F�a<o�a<`�a<y�a<ˮa<��a<Lva<�Oa<&a<{�`<��`<3�`</�`<1�`<-�`<s�`<Q�`<�`<��`<%a<9Ga<�pa<��a<M�a<{�a<��a<��a<��a<k�a<�a<c�a<I�a<d�a<��a<�a<Õa<��a<	�a<z�a<:�a<��a<�a<`�a<��a<`�a<��a<��a<��a<�a<�ca<=9a<�a<W�`<��`<��`<˧`<:�`<��`<?�`<��`<�a<�Ca<=na<ŕa<��a<C�a<��a<�a<~�a<��a<K�a<S�a<��a<z�a<��a<�a<
�a<[�a<��a<6�a<��a<�a<��a<k�a<��a<O�a<��a<Q�a<@�a<�a<��a<Xa<�,a<a<]�`<r�`<̮`<�`<K�`<��`<P�`<�`<0'a<yRa<:|a<�a<�a<��a<	�a<��a<��a<��a<�a<u�a<�a<��a<�a<-�a<J�a<��a<ݦa<>�a<L�a<��a<��a<?�a<��a<��a<F�a<��a<��a<�a<�na<FDa<�a<��`<�`<E�`<n�`<��`<۫`<��`<`�`<a<3/a<Za<v�a<�a<��a<��a<_�a<��a<��a<'�a<�a<��a<Ϊa<"�a<��a<;�a<!�a<J�a<ڙa<��a<��a<K�a<�a<��a<��a<��a<}�a<f�a<�a<�qa<�Ha<�a<?�`<��`<M�`<G�`<ņ`<y�`<1�`<+�`<�`<<�`<�a<�Ha<�oa<!�a<D�a< �a<��a<��a<g�a<��a<�a<!�a<D�a<�~a<�wa<�ta<uua<^za<��a<�a<��a<C�a<ͳa<ݻa<C�a<S�a<�a<��a<Bwa<�Qa<(a<��`<��`<4�`<M�`<�~`<�w`<s}`<�`<ߪ`<��`<I�`<�#a<�  �  2`a<�a<�a<(�a<I�a<ٻa<��a<��a<w�a<ۇa<fva<&ga<�[a<�Ta<Sa<�Va<g_a<�la<<}a<��a<ѡa<!�a<��a<$�a<��a<2�a<�a<�a<ca<:=a<�a<��`<��`<�`<0�`<��`<Ҹ`<��`<y�`<�a<34a<!\a<a<<�a<��a<{�a<q�a<��a<j�a<��a</�a<F�a<�a<��a<�va<\ra<sa<�xa<Ճa<��a<��a<[�a<��a<��a<��a<��a<,�a<��a<��a<M�a<mxa<�Qa<d+a<ua<�`<��`<�`<U�`<��`<��`<a<P4a<8[a<Ӂa<�a<g�a<�a<�a<F�a<M�a<��a<��a<�a<K�a<ӗa<Њa<�a<B~a<�a<��a<�a<<�a<�a<��a<��a<�a<��a<8�a<T�a<r�a<K�a<r�a<�ma<�Fa<� a<��`<��`<x�`<d�`<�`<��`<��`<Ja<�Aa<�ha<|�a<دa<��a<a�a<#�a<S�a<��a<e�a<��a<��a<ݠa<)�a<+�a<�}a<�{a<l~a<��a<:�a<C�a<�a<x�a<�a<��a<��a<M�a<@�a<]�a<��a<�a<e[a<P4a<~a<m�`<�`<p�`<��`<=�`<U�`<��`< "a<EHa<�na<D�a<^�a<M�a<��a<�a<�a<��a<>�a<6�a<��a<q�a<?�a<�ta<�na<ima<{qa<�za<��a< �a<��a<��a<�a<r�a<��a< �a<8�a<֡a<$�a<]a<X5a<�a<��`<��`<��`<�`<��`<�`<��`<l�`<a<e6a<t\a<$a<��a< �a<��a<7�a<��a<űa<��a<ݏa<�}a<�la<,_a<�Ua<�Qa<�Ra<\Ya<vda<dsa<Ȅa<y�a<�a<��a<��a<��a<�a<՞a<��a<�ca<�=a<�a<��`<i�`<`�`<Y�`<_�`<?�`<1�`<q�`<�`<�a<:a<�  �  �sa<��a<�a<)�a<4�a<¶a<j�a<��a<j�a<uma<Wa<�Ca<�4a<�+a<�)a<.a<J9a<�Ia<�^a<bva<�a<��a<��a<�a<��a<Q�a<�a<�a<�wa<Wa<�5a<Ea<c�`<��`<��`<+�`<r�`<#�`<�a<.a<:Pa<;sa<ޓa</�a<��a<��a<��a<=�a<9�a<�a<h�a<�a</ma<�[a<fOa<]Ia<�Ia<Qa<�^a<pqa<�a<��a<r�a<��a<\�a<:�a<��a<��a<(�a<�a<��a<Cma<	La<6-a<�a<3a<��`<��`<�a<!a< 4a<�Sa<�ua<:�a<t�a<��a<��a<��a<��a<��a<��a<K�a<t�a<q�a<�ua<ea<�Ya<Ua<�Va<�_a< na<r�a<�a<8�a<K�a<��a<��a<��a<��a<��a<d�a<��a<�a<da<Ca<�%a<la<|�`<�`<F�`<a<2"a<�>a<�_a<{�a<4�a<z�a<�a<c�a<�a<:�a<��a<��a<��a<T�a<��a<�ma<b^a<�Ta<5Ra<�Ua<�`a<�pa<�a<��a<��a<x�a<��a<��a<_�a<Z�a<5�a<}�a<��a<7ua<BSa<�2a<Ka<�a<��`<��`<��`<�a<�$a<HCa<Pda<�a<e�a<U�a<��a<��a<B�a<P�a<��a<��a<q�a<d�a<�na<�[a<[Ma<�Ea<TDa<�Ia<�Ua<fa<={a<��a<k�a<Q�a<&�a<��a<��a<��a<?�a<��a<�sa<�Pa<�.a<�a<�`<��`<��`<��`<�`<
�`<Oa<�/a<�Pa<�qa<��a<Q�a<̷a<3�a<��a<6�a<ǣa<��a<Nwa<�_a<uJa<l9a<�-a<�(a<
*a<R2a<�@a<�Sa<�ia<ۀa<��a<��a<�a<M�a<Q�a<$�a<��a<�va<Va<�3a<�a<O�`<4�`<S�`<��`<\�`<L�`<��`<�a<�0a<�Ra<�  �  ��a<��a<��a<��a<s�a<��a<��a<��a<~la<�Oa<Q4a<�a<o
a<]�`<b�`<�a<xa<�#a<7=a<�Ya<Rwa<�a<�a<,�a<�a<Ϳa<�a<J�a<݌a<�qa<aUa<�:a<J$a<�a<E
a<$	a<na<�a<,5a<�Oa<&ma<��a<��a<��a<��a<}�a<�a<'�a<��a<ҙa<�~a<�ba<�Ha<s3a<&$a<Ma<�a<�%a<	6a<�La<�ga<p�a<��a<ؼa<��a<$�a<�a<��a<�a<�a<�a<��a<?ma<ISa<>a</a<�'a<�(a<�1a<vBa<Ya<�sa<Ȑa<۬a<k�a<i�a<��a<��a<b�a<��a<k�a<C�a<��a<>ia<�Oa<~;a<�-a<�'a<*a<�4a<�Fa< ^a<�ya<��a<c�a<<�a<+�a<?�a<��a<��a<�a<��a<�a<�a<�ea<Ma<�9a<�,a<(a<�+a<�7a<;Ja<^ba<~a<�a<��a<��a<D�a<��a<N�a<�a<��a<T�a<×a<�za<�^a<�Fa<�3a<O(a<�$a<�)a<�6a<MJa<(ca</a<�a<]�a<E�a<��a<��a<��a<:�a<��a<��a<ԏa<�ra<�Wa<4@a<�.a<�$a<�"a<�(a<7a<�Ka<ea<A�a<��a<.�a<��a<|�a<��a<��a<<�a<)�a<��a<��a<�ea<aJa<43a<"a<va<(a<)a<�,a<�Aa<.[a<wa<��a<1�a<m�a<h�a<��a<?�a<$�a<�a<�a<&ma<�Oa<�4a<�a<�a<�a<�a<ha<]a<d5a<�Oa<�ka<�a<��a<��a<�a<-�a<`�a<A�a<Y�a<�xa<v[a<�>a<�$a<�a<�a<:�`<K�`<�a<
a<R0a<~Ka<Dha<ȃa<e�a<�a<��a<$�a<G�a<>�a<ĉa<�na<�Qa<�5a<�a<Y	a<��`<��`<��`<�a<�a<3a<Oa<9la<�  �  ��a<6�a<��a<��a<Ӵa<}�a<$�a<�sa<�Ra<	1a<�a<[�`<��`<��`<b�`<��`<|�`<h�`<�a<8<a<�^a<�a<ƛa<[�a<u�a<h�a<�a<�a<�a<��a<�sa<f^a<La<�>a<7a<p6a<M<a<�Ha<�Za<�pa<��a<i�a<��a<O�a<��a<9�a<��a<+�a<r�a<݃a<ca<@Ba<�#a<�	a<��`<k�`<��`<��`<a<�&a<�Fa<\ia<&�a<��a<�a<-�a<?�a<@�a<�a<��a<�a<��a<��a<^xa<ga<�Za<�Ta<�Ua<]a<�ja<-}a<�a<W�a<��a<��a<*�a<��a<��a<-�a<�a<K�a<h�a<[ha<(Ga<�(a<�a<~ a<��`<_�`<�a<�a<�9a<IZa<M|a<��a<�a<v�a<�a<��a<4�a<��a<&�a<�a<Ԟa<�a<�sa<�ca</Ya<�Ua<PXa<�aa<&qa<�a<��a<��a<��a<4�a<-�a<7�a<��a<��a<4�a<E�a<~a<�[a<�:a<Da<;a<��`<��`<v�`<�a<�"a<�@a<paa<f�a<��a<�a<��a<(�a<e�a<Y�a<x�a<�a<��a<h�a<{a<�ga<�Ya<dQa<�Oa<�Ta<p`a<qa<��a<Ϝa<I�a<O�a<~�a<��a<x�a<l�a<D�a<�a<��a<ha<�Ea<%a<�	a<��`<��`<8�`<y�`<�a<�a<C:a<�Za<|a<R�a<ղa<m�a<
�a<��a<-�a<Y�a<��a<
�a<pa<�Ya<�Ga<Z:a<�3a<�3a<�:a<�Ga<zYa<�na<��a<O�a<��a<úa<�a<+�a<2�a<�a<A�a<�`a<F>a<�a<��`<E�`<��`<<�`<��`<��`<]�`<a<7,a<�Ma<oa<I�a<f�a<Ȳa<�a<��a<�a<&�a<ʅa<�na<�Wa<FCa<U3a<�(a<b%a<P(a<2a<�Aa<�Ua<~la<Ӄa<�  �  �a<2�a<`�a<ùa<��a<e�a<:�a<�_a<�9a<�a<��`<��`<��`<��`<Ţ`<ȩ`<̻`<��`<��`<Ma<�Fa<�la<��a<N�a<T�a<b�a<��a<)�a<��a<�a<C�a<f~a<!pa<�ea<�_a<�_a<rda<�na<�|a<9�a<�a<r�a<r�a<��a<�a<M�a<��a<��a<��a<,na<fHa<q"a<l�`<��`<��`<��`<O�`<��`<f�`<Ka<�&a<8Na<�ua<��a<�a<��a<��a<��a<��a<��a<p�a<@�a<��a<ߙa<H�a<��a<~a<�~a<v�a<!�a<��a<��a<��a<��a<z�a<��a<��a<	�a<��a<��a<�a<sa<�Ka<�%a<�a<_�`<��`<��`<�`<9�`<�`<�a<�;a<�ba<#�a<��a<��a<=�a<��a<��a<Y�a<	�a<�a<[�a<��a<{�a<��a<��a<�~a<��a<��a<q�a<�a<��a<L�a<n�a<4�a<�a<�a<f�a<��a<H�a<E�a<ea<�=a<&a<��`<��`<|�`<�`<��`<��`<5�`<�a<|Da<rka<��a<�a<��a< �a<Z�a<=�a<��a<��a<��a<��a<�a<�a<܀a<Gza<ya<�|a<�a<�a<��a<�a<V�a<�a<��a<��a<��a<}�a<��a<0�a<�ta<tMa<�%a<� a<R�`<��`<�`<��`<&�`<4�`<W�`<�a<�?a<�ea<�a<��a<�a<��a<Y�a<��a<s�a<�a<��a<�a<O{a<�la<Kba<�\a<�\a<�aa<la<�ya<��a<�a<��a<��a<5�a<��a<��a<��a<B�a<�na<yIa<�!a</�`<��`<�`<ϩ`<��`<Q�`<�`<��`<��`<�a<f4a<�Za<�|a<˘a<�a<:�a<Һa<z�a<�a<�a<�a<7va< fa<�Ya<lQa<�Na<�Pa<�Xa<�da<�ta<��a<��a<�  �  ��a<��a<T�a<n�a<٩a<��a<2sa<(Ma<Y#a<0�`<t�`</�`<,�`<ŀ`<Z|`<8�`<ؗ`<��`<)�`<�a<`1a<W[a<��a<W�a<��a<��a<��a<��a<Ƚa<��a<��a<#�a<��a<�a<��a<c�a<�a<+�a<�a<�a<�a<��a<��a<h�a<��a<~�a<��a<��a<0�a<ZZa<�0a<ma<��`<��`<��`<М`<�`<j�`<;�`<c�`<.
a<�5a<�aa<��a<s�a<%�a<��a<��a<�a<��a<8�a<��a<x�a<�a<��a<��a<ʠa<M�a<�a<߭a<Ӹa<��a<e�a<��a<e�a<��a<��a<��a<�a<7�a<Ԇa<�]a<�2a<�a<��`<��`<G�`<��`<�`<��`<��`<��`<l a<�Ka<2va<�a<��a<�a<��a<�a<P�a<u�a<��a<]�a<ҿa<��a<E�a<�a<��a<{�a<�a<�a<нa<�a<S�a<a�a<��a<��a<��a<��a<	�a<>�a<�xa<�Na<�"a<��`<	�`<��`<��`<��`<�`<�`<(�`<� a<�*a<�Ua<a<�a<��a<9�a<��a<)�a<*�a<��a<��a<�a<Եa<p�a<�a<�a<Лa<��a<��a<��a<ֻa<�a<��a<h�a<��a<G�a<��a<f�a<��a<��a<"aa<�5a<�	a<v�`<x�`<��`<��`<l�`<��`<�`<o�`<~�`<�'a<�Qa<�xa<4�a<`�a<J�a<Y�a<&�a<R�a<��a<>�a<ޤa<Q�a<+�a<0�a<�a<za<q�a<��a<�a<��a<��a<3�a<��a<��a<��a<Z�a<�a<��a<�]a<W4a<�a<��`<�`<(�`<^�`<8{`<_~`<�`<��`<�`<a�`<�a<�Ga<@na<��a<Ȧa<k�a<L�a<l�a<h�a<k�a<�a<v�a<K�a<�ya<�sa<fqa<isa<>ya<f�a<p�a<�a<��a<�  �  ��a<��a<��a<��a<��a<5�a<�ga<[>a<Na<�`<��`<ő`<�t`<�c`<�^`<?g`<�{`<ԛ`< �`<��`< a<CMa<va<��a<1�a<��a<�a<c�a<�a<��a<Y�a<E�a<K�a<�a<��a<��a<؟a<ԥa<��a<��a<��a<��a<7�a<X�a<��a<��a<~�a<�a<�ta<~Ja<Ka<c�`<D�`<��`<"�`<H`<s`<ٌ`<�`<s�`<��`<B"a<lQa<�}a<z�a<��a<7�a<��a<��a<��a<��a<=�a<S�a<�a<�a<��a<�a<^�a<��a<��a<Q�a<��a<�a<<�a<��a<��a<��a<��a<��a<��a<ya<�La<Xa<��`<Z�`<�`<l�`<؉`<��`<D�`<>�`<��`<�
a<_9a<ga<#�a<�a<��a<��a<��a<�a<��a<��a<��a<��a<��a<Z�a<��a<׻a<D�a<f�a<b�a<@�a<�a<��a<��a<��a<N�a<��a<��a<��a<��a<�ia<�<a<�a<�`<��`<T�`<^�`<�`<�`<�`<F�`<��`<	a<�Da<qa<�a<�a<��a<��a<T�a<��a<��a<��a<��a<��a<;�a<��a<�a<�a<Z�a<X�a<�a<�a<��a<��a<��a<��a<a�a<��a<8�a<�a<}a<HQa<]"a<��`<��`<\�`<�`<r{`<�y`<m�`<��`<~�`</�`<�a<^Aa<�ka<8�a<Үa<��a<�a<��a<R�a<Y�a<��a<��a<w�a<��a<W�a<ՙa<��a<;�a<��a<��a<��a<3�a<��a<��a<C�a<��a<Q�a<ۘa<xa<%Pa<e#a<Z�`< �`<`�`<s}`<�g`<�]`<a`<3q`<Ռ`<�`<��`<a<y8a<Mba<ͅa<M�a<"�a<0�a< �a<��a<L�a<��a<��a<Z�a<�a<e�a<��a<+�a<~�a<��a<ۡa<��a<�a<�  �  ��a<u�a<7�a<�a<�a<��a<�_a<�4a<�a<��`<M�`<��`<c`<�P`<�K`<hT`<Xj`<?�`<��`<��`<a<FDa<�na<��a<�a<��a<�a<��a<��a<��a<��a<y�a<z�a<�a<�a<N�a<ٯa<Ĵa<��a<��a<��a<f�a<��a<F�a<��a<;�a<0�a<��a<Ola<v@a<,a<O�`<:�`<o�`<�y`<Ol`<�l`<Pz`<��`<D�`<��`<�a<)Ga<Dua<�a<�a<��a<q�a<]�a<��a<4�a<��a<C�a<�a<��a<��a<��a<��a<i�a<C�a<��a<]�a<�a<:�a<-�a<��a<��a<��a<׻a<��a<Mpa<Ba<�a<��`<ڸ`<a�`<��`<�v`<�z`<*�`<S�`<�`<T�`<�-a<w]a<D�a<
�a<��a<��a<D�a<��a<��a<��a<R�a<��a<`�a<��a<��a<��a<��a<��a<2�a<�a<��a<��a<1�a<~�a<��a<1�a<��a<	�a<��a<�`a<�0a<i a<��`<ɪ`<`�`<jy`<�s`<|`<h�`<��`<��`<	a<x9a< ha<ϑa<�a<��a<��a<R�a<@�a<��a<��a<��a<+�a<j�a<:�a<_�a<��a<\�a<J�a<*�a<D�a<��a<S�a<F�a<��a<S�a<��a<�a<��a<�ta<AGa<>a<��`<ȸ`<3�`<�w`<zh`<�f`<�r`<m�`<N�`<��`<�a<7a<�ca<��a<P�a<o�a<��a<a�a<��a<��a<9�a<��a<h�a<]�a<E�a<��a<�a<�a<"�a<�a<�a<2�a<��a<T�a<~�a<�a<J�a<�a<qa<YGa<�a<��`<U�`<�`<�k`<�T`<�J`<N`<_`<�{`<b�`<M�`<N�`<�.a<nZa<�a<k�a<R�a<��a<��a<��a<Z�a<��a<�a<�a<)�a<��a<h�a<t�a<ՠa<��a<��a<��a<5�a<�  �  V�a<��a<p�a<J�a<�a<i�a<(^a<�#a<l�`<��`<�b`<�,`<`<b�_<��_<O�_<�`<�9`<Ts`<�`<��`<�6a<pa<��a<��a<(�a<��a<1�a<z�a<��a<��a<��a<��a<#�a<3�a<��a<��a<��a<��a<Z�a<��a<�a<��a<��a<7�a<.�a<��a<�a<+fa<**a<��`<�`<Gm`<~;`<|`<�`<�`<P`<�;`<�m`<��`<��`<x/a<na<��a<��a<��a<�b<�b<�b<�b<)b<��a<@�a<��a<��a<��a<��a<[�a<��a<��a<�b<�b<~b<Yb<Cb<rb<��a<��a<��a<!ea<&a<�`<��`<�i`<�;`<�`<�`<�`<�+`<-T`<��`<�`<
a<+Ka<��a<]�a<��a<h�a<b<�b<b<�b<Ib<��a<H�a<E�a<��a<��a<Y�a<x�a<+�a<�a<�b<�b<�b<�b<�b<@�a<��a<��a<݊a<Pa<Ha<�`<��`<W`<-`<�`<�`<�`<T4`< a`<��`<��`<�a<�Za<��a<��a<��a<��a<�
b<Mb<�b<rb< �a<�a<��a<�a<N�a<��a<Q�a<�a<A�a<��a<� b<�b<�b<�
b<�b<�a<2�a<��a<oa<Y1a<��`<��`<�n`<X;`<w`<� `<��_<�`<2`<�b`<��`<��`<�a<�[a<Őa<��a<��a<�a<��a<[�a<v�a<��a<�a<��a<)�a<_�a<��a<=�a<��a<��a<B�a<}�a<e�a<v�a<��a<A�a<��a<��a<'�a<�sa<�;a<�`<w�`<�x`<2>`<s`<V�_<��_<]�_<�_<
&`<1[`<W�`<��`<�a<Wa<��a<��a<�a<y�a<��a<�a<��a<�a<.�a<��a<��a<k�a<_�a<I�a<��a<��a<��a<��a<Q�a<�  �  p�a<��a<e�a<s�a<W�a<^�a<ba<j(a<��`<��`<5j`<z4`<�`<1�_<C�_<�_<�`<�A`<iz`<�`<��`<(;a<�sa<��a<��a<�a<��a<%�a<g�a<��a<K�a<4�a<��a<E�a<�a<H�a<��a<�a<3�a<N�a<B�a<��a<��a<-�a<��a<��a<l�a<R�a<Tja<,/a<`�`<��`<�t`<�C`<1 `<q`<g`< `<�C`<^u`<i�`<��`<�4a<Fra<�a<*�a<{�a<�b<4b<b<�b<�b<��a<��a<�a<��a<��a<��a<t�a<S�a<3�a<��a<�b<Ob<0b<b<4b<��a<k�a<��a<�ia<t+a<6�`<��`<�q`<�C`<�$`<H`<�`<i4`<.\`<�`<��`<�a<�Oa<��a<k�a<��a<��a<b<�b<3b<�
b<,b<6�a<T�a<��a<��a<I�a<9�a<��a<�a<��a<^ b<	b<�b<�b<�b<j�a<��a<�a<��a<�Ta<�a<`�`<-�`<�^`<�5`<�`</`<i`<�<`<�h`<Р`<��`<� a<t_a<`�a<f�a<��a<��a<j
b<Bb<�	b<gb<`�a<��a<]�a<-�a<�a<��a<G�a<h�a<��a<��a<A�a<Vb<[
b<#
b<�b<��a<��a<��a<Csa<Z6a<��`<5�`<lv`<hC`<,`<�	`<�`<j`<%:`<j`<D�`<��`<�#a<�_a<�a<��a<i�a<x�a<M�a<��a<�a<�a<'�a<��a<��a<c�a<�a<
�a<�a<Y�a<��a<��a<-�a<G�a<��a<�a<��a<��a<�a<{wa<�?a<Wa<��`<�`<�E`<�`<�_<C�_<)�_<�`<	.`<�b`<��`<��`<� a<[a<��a<�a<f�a<��a<�a<B�a<��a<��a<��a<��a<%�a<V�a<�a<,�a<ҹa<��a<W�a<l�a<��a<�  �  ��a<��a<��a<��a<��a<X�a<�la<�5a<��`<R�`<`<[K`<�#`<`<C`<�`<�,`<1X`<Ɏ`<��`<Ka<�Ga<�}a<�a<��a<��a<o�a<
�a<��a<��a<@�a<T�a<�a<��a<@�a<=�a<��a<C�a<�a<��a<�a<��a<M�a<��a<��a<��a<��a<8�a<�ua<@=a<, a<��`<^�`<�Z`<,9`<e'`<X'`<;9`<A[`<J�`<��`<�a<Ca<
~a<C�a<��a<��a<vb<'b<�b<�b<��a<��a<��a<��a<��a<��a<��a<��a<a�a<�a<Z�a<��a<fb<�b<�b<Pb<��a<��a<U�a<�ua<�:a<��`<Ͼ`<݇`<�[`<=>`<E1`<�6`<M`<?s`<.�`<(�`< a<Z]a<��a<��a<��a<b<�b<�b<�b<Sb<>�a<>�a<��a<K�a<2�a<*�a<��a<D�a<�a<^�a<�a<# b<�	b<Tb<(b<~b<��a<z�a<i�a<�aa<�$a<��`<�`<�u`<�M`<�5`<4.`<9`<�T`<I`<5�`<��`<R0a<la<z�a<��a<�a<b<<
b<)
b<Db<��a<V�a<��a<��a<l�a<Y�a<|�a<�a<��a<\�a<�a<
�a<_�a<�b<�b<1b<��a<.�a<ܰa<�~a<mDa<�a<v�`<�`<�Z`<&7`<~#`<�!`<�1`<�Q`<�`<Է`<��`<`2a<�ka<J�a<Q�a<��a<��a<C�a<��a<w�a<:�a<�a<"�a<!�a<D�a<��a<1�a<-�a<h�a<}�a<O�a<�a<\�a</�a<��a<��a<��a<�a<D�a<2La<`a<$�`<��`<1\`<�/`<�`<;`<	`<@`<E`<�w`<`�`<��`<.a<�ea<ڔa<˸a<��a<4�a<�a<��a<=�a<�a<�a<?�a<�a<�a<��a<��a<q�a<��a<�a<#�a<��a<�  �  ��a<K�a<A�a<c�a<��a<~�a<�|a<�Ia<xa<�`<��`<uo`<�J`<4`<�-`<|8`<$S`<�{`<l�`<��`<�"a<![a<(�a<)�a<��a<z�a<��a<��a<��a<��a<߸a<0�a<؛a<`�a<o�a<	�a<��a<��a<��a<v�a<q�a<F�a<	�a<�a<��a<��a<2�a<��a<[�a<�Ra<a<��`<�`<�`<M``<�O`<�O`<�``<��`<t�`<Z�`<&a<+Ya<�a<*�a<��a<g�a<	b<�
b<b<�a<��a<��a<�a<Q�a<��a<k�a<��a< �a<ûa<^�a<t�a<��a<��a<�b<xb<�b<1�a<`�a<8�a<��a<�Qa</a<	�`<ݪ`<��`<�e`<�Y`<�^`<�s`<��`<�`<X�`<�8a<!ra<4�a<G�a<S�a<]b<�b< b<\b<��a<�a<��a<��a<��a<��a<�a<�a<��a<��a<:�a<��a<��a<��a<
b<�b<Xb<��a<��a<��a<2va<\=a<�a<��`< �`<�t`<�]`<�V`<�``<�z`<��`<��`<xa<�Ga<za<ɰa<�a<�a<�b<�b<�b<9�a<]�a<��a<��a<�a<E�a<��a<E�a<��a<�a<D�a<��a<i�a<��a<d�a<b<8b<��a<~�a<P�a<G�a<Za<xa<r�`<ԭ`<�`<G^`<�K`<J`<�X`<(w`<�`<7�`<=a<�Ha<�}a<3�a<�a<Y�a<��a<�a<��a<��a<%�a<#�a<��a<٘a<_�a<_�a<=�a<��a<̗a<ڤa<j�a<&�a<��a<s�a<p�a<R�a<%�a<жa< �a< _a<y'a<�`<ղ`<(`<}U`<<9`<�,`<:1`< F`<�i`<��`<��`<�	a<�Ba<�va<q�a<A�a<�a<3�a<H�a<u�a<��a<Q�a<a�a<E�a<��a<z~a<�{a<~a<�a<�a<��a<�a<i�a<�  �  b�a<��a<�a<��a<��a<v�a< �a<�ba<�/a<*�`<��`<L�`<�{`<�g`<6b`<�k`<��`<k�`<��`<�
a<�?a<�ra<0�a<��a<a�a<��a<M�a<6�a<�a<�a<��a<'�a<�sa<=fa<�^a<&^a<da<�pa<��a<��a<�a<�a<��a<��a<��a<�a<��a<e�a<��a<�ma<a:a<�a<��`<M�`<��`<݃`<�`<+�`<P�`<��`<�	a<?a<�ta<ԥa<t�a<��a<b<f	b<Qb<q�a<�a<��a<��a<-�a<��a<k�a<�}a<M~a<��a<%�a<��a<ٻa<��a<F�a<��a<Kb<v
b<b<��a<��a<�a<.na<|9a<�a<A�`<(�`<��`<@�`<��`<��`<�`<��`<#a<�Wa<��a<�a<��a<��a<M	b<)b<Yb<��a<`�a<��a<{�a<�a<�a<��a<�}a<ǀa<D�a<��a<k�a<:�a<��a<��a<�b<i
b<�b<4�a<��a<ܼa<%�a<�[a<�&a<��`<��`<�`<B�`<<�`<.�`<«`<��`<�`<f0a<ea<5�a<��a<��a<��a<1b<"b<\�a<y�a<��a<�a<��a<e�a<�a<�ya<]xa<e}a<�a<˙a<Ѯa<��a<.�a<�a<��a<�b<��a<��a<�a<m�a<�ta<�?a<N
a<��`<&�`<��`<�`<;~`<��`<Ѧ`<d�`<��`<40a<�ca<��a<��a<*�a<�a<��a<u�a<H�a<��a<u�a<�a<��a<?oa<$ba<�[a<�[a<?ba<0oa<+�a<ϖa<�a<:�a<.�a<?�a<��a<�a<	�a<��a<9va<�Ca<�a<z�`<��`<�`<Kl`<&a`<	e`<�w`<ۗ`<d�`<?�`<�(a<V\a<{�a<��a<��a<�a<��a<��a<��a<[�a<{�a<Aa<�ja<�Za<oPa<�La<�Oa<�Ya<ia<8}a<Z�a<`�a<�  �  !�a<6�a<��a<��a<2�a<=�a<R�a<�}a<QQa<H#a<d�`<J�`<-�`<��`<ǝ`<4�`<?�`<R�`<�a<41a<�_a<:�a<�a<i�a<��a<r�a<��a<��a<�a<�a<�xa<�[a<{Ca<�1a<�'a<�&a<,.a<(>a<oUa<ra<Αa<n�a<�a<r�a<v�a<f�a<V�a<G�a<�a<��a<^a<01a<�a<��`<��`</�`<n�`<��`<?�`<�	a<�4a<�ca<?�a<�a<
�a<�a<b<�b<��a<��a<��a<��a<̐a<�ta<�]a<�Ma<Fa<�Fa<�Pa<Nba<�za<��a<��a<��a<�a<b<�	b<�b<o�a<��a<��a<u�a<h_a<M2a<�	a<�`<4�`<��`<��`<D�`<��`<7 a<�Ka<=za<R�a<��a<K�a<�b<2b<�b<X�a<E�a<��a<¦a<W�a<�ma<�Xa<*Ka<SFa<Ja<XVa<vja<��a<��a<`�a<>�a<��a<Ub<�	b<�b<c�a<�a<�a<A}a<�Na<y"a<��`<P�`<7�`<��`<��`< �`<�a<X*a<Wa<�a<��a<��a<f�a<�b<b<��a<��a<��a<׵a<��a<3ya<`a<sMa<�Ba<�@a<sGa<tVa<�la<-�a<��a<�a<W�a<X�a<� b<Eb<��a<��a<̻a<�a<wca<�4a<8	a<��`<��`<H�`<��`<�`<��`<��`<�'a<�Ta<��a<��a<�a<��a<�a<��a<��a<^�a<g�a<�a<?ra<5Ua<U=a<�,a<$a<D$a<@-a<\>a<Va<�ra<�a<��a<��a<�a<��a<��a<��a<��a<ߎa<8ca<�4a<a<��`<̼`<{�`<��`<�`<]�`<V�`<��`<"a<$Ka<�wa<c�a<x�a<��a<��a<C�a<��a<p�a<��a<�ua<)Wa<Z<a<X'a< a<Da<%a<�%a<:a<hTa<�ra<�a<�  �  -�a<��a<t�a<e�a<@�a<�a<*�a<��a<sa<RLa<W'a<ha<�`<j�`<^�`<��`<8�`<7a<32a<�Xa<�a<��a<;�a<��a<%�a<U�a<��a<��a<��a<�va<cPa<�,a<a<��`<,�`<w�`<��`<�a<U#a<�Fa<�ma<[�a<��a<8�a<H�a<!�a<��a<w�a<!�a<V�a<T�a<~\a<�9a<�a< a<��`<��`<?	a<�a<�<a<aa<��a<��a<��a<��a<b<�b<�b<)�a<��a<��a<{�a<!fa<JCa<�&a<�a<�a<5
a<Xa<P,a<�Ja<�na<b�a<$�a<��a<C�a<�b<�	b<� b<Q�a<0�a<��a<(�a<`a<�=a<�"a<ca<ya<�a<�a<[1a<�Pa<�ua<Ȝa<*�a<��a<��a<�b<^
b<��a<��a<�a<֧a<�a<;[a<
:a<�a<=a<�a<�a<Ka<M6a<�Va<�{a<��a<C�a<^�a<��a<Tb<�b<A�a<��a<�a<��a<�wa<wRa<2a<Ba<
a<�a<$a<(a<�7a<�Xa<�~a<1�a<�a<��a<��a<sb<�b<��a<��a<��a<t�a<yna<�Ia<�*a<�a<7a<�a<a<�a<�:a<�\a<˂a<��a<��a<�a<��a<�b<��a<�a<�a<y�a<��a<`a<];a<}a<a<��`<�`<�a<2a<�1a<�Sa<�ya<�a<��a<�a<��a<��a<�a<V�a<��a<2�a<oa<�Ga<�#a<:a<��`<��`<��`<�`<aa<"&a<�Ia<�oa<�a<�a<.�a<�a<c�a<R�a<�a<r�a<n�a<W[a<�4a<$a<I�`<��`<H�`<�`<��`<a<]"a<�Fa<�ma<Βa<�a<�a<��a< �a<�a<�a<N�a<�va<�Oa<*a<�a<��`<"�`<��`<�`<��`<�a<�&a<-La<Bsa<�  �  �~a<5�a<��a<��a<=�a<�a<�a<�a<�a<Hsa<�Ua<�;a<G(a<�a<�a<Ra<�-a<ZCa<�^a<�}a<W�a<P�a<��a<�a<��a<1�a<��a<��a<<�a<�Sa<;&a<~�`<�`<.�`<�`<�`<ߵ`<R�`<c�`<[a<�Ga<�va<`�a<�a<)�a<��a<��a<��a<��a<=�a<�a<��a<ja<�Ra<�Ba<Z:a<�:a<Da<�Ua<�ma<L�a<8�a<|�a<$�a<�a<�b<�b<5�a<��a<l�a<��a<�fa<�9a<a<��`<�`<u�`<��`<]�`<��`<�a<�Ca<�qa<�a<��a<{�a<��a</	b<�b<��a<�a<D�a<��a<�a<|pa<�Za<�Ka<�Ea<1Ha<SSa<pfa<�a<��a<��a<\�a<c�a<�b<Mb<ab<:�a<��a<I�a<\�a<Ya<^,a<�a<��`<��`<G�`<�`<��`<q a<'a<ISa<i�a<��a<��a<K�a<�b<�	b<1b<��a<u�a<�a<ߞa<��a<�fa<�Ra<cFa<�Ba<�Ga<�Ua<�ja<��a<�a<��a<��a<k�a<#b<�b<��a<��a<��a<��a<�ra<RDa<�a<��`<�`<�`<
�`<�`<��`<�a<m/a<u\a<+�a<��a<��a<��a<t�a<b<O�a<i�a<]�a<k�a<|�a<�ka<�Ra<�@a<r6a<5a<k<a<
La<�ba</~a<W�a<�a<��a<�a<��a<��a<��a<��a<S�a<Bxa<�Ia<a<��`<��`<ܴ`<|�`<B�`<
�`<��`<X�`<�a<La<�xa<�a<a�a<;�a<�a<��a<��a<U�a<�a<�a<`a<�Da<#.a<a<�a<�a<Y%a<#8a<FQa<�na<��a<��a<��a<��a<H�a<)�a<��a<<�a<��a<yVa<(a<L�`<��`<��`<��`<V�`<K�`<��`<�`<�`<�#a<�Qa<�  �  da<_�a<��a<�a<[�a<n�a<M�a<��a<�a<S�a<�~a<2ka<]\a<tSa<1Qa<�Ua<�`a<lqa<��a<V�a<��a<M�a<.�a<"�a<N�a<��a<�a<K�a<=da<1a<��`<��`<W�`<l�`<�q`<^o`<�{`<��`<K�`<)�`<"a<�Wa<�a<l�a<��a<{�a<#�a<K�a<4�a<S�a<K�a<��a<k�a<�a<�wa<�qa<Sra<�ya<+�a<��a<��a<8�a<Y�a<��a<Ob<b<Kb<r�a<��a<�a<nva<"Ba<a<x�`<��`<M�`<��`<��`<?�`<x�`<��`<�a<9Na<P�a<��a<��a<��a<Fb<b<�b<P�a<��a<=�a<�a<�a<@�a<��a<N}a<Ga<Շa<r�a<٩a<��a<n�a<��a<f b<�
b<"b<��a<o�a<��a<u�a<�fa<2a<��`<��`<�`<�`<��`<:�`<��`<��`<��`<�+a<6`a<�a<	�a<��a<j�a<�b<�	b< b<(�a<��a<��a<�a<��a<��a<<}a<oza<K~a<ƈa<Ԙa<O�a<^�a<��a<��a< b<>b<�b<D�a<��a<��a<��a<�Oa<a<:�`<�`<@�`<�`<��`<
�`<�`<x�`<5a<�6a<Jka<[�a<B�a<�a<L�a<[b<��a<�a<p�a<��a<�a<�a<܃a<�ua<�ma<�la<�qa<�}a<��a<��a<Y�a<��a<[�a<i�a<��a<Q�a<�a<�a<Ջa<$Za<�$a<��`<�`<X�`<{`<m`<�m`<�}`<��`<�`<��`<�(a<;\a<�a<۱a<��a<�a<N�a<��a<}�a<h�a<T�a<�a<ra<�`a< Ua<Pa<�Qa<�Ya<ha<9{a<��a<J�a<~�a<��a<��a< �a<��a<�a<�a<�ha<6a<a<��`<|�`<}`<
f`<�]`<}d`<z`<Z�`<��`<��`<�0a<�  �  nKa<j~a<ݧa<!�a<E�a<��a<��a<i�a<X�a<2�a<̠a<��a<�a<Ła<!�a<��a<p�a<��a<`�a<Ѹa<��a<��a<w�a<W�a<�a<�a<�a<~a<cJa<�a<��`<ѡ`<�s`<xQ`<>`<;`<�H`<mf`<8�`<��`<  a<~;a<Tsa<E�a<��a<��a<��a<��a<��a<<�a<��a<��a<j�a<�a<g�a<l�a<�a<��a<��a<��a<d�a<��a<��a<� b<�b<Tb<K�a<�a<8�a<��a<�Za<� a<N�`<�`<Ӈ`<�i`<�Z`<�\`<�n`<j�`<��`<�`<I.a<�ga<ߜa<��a<i�a<vb<�b<nb<�b<��a<�a<�a<��a<��a<��a<?�a<ʭa<ѳa<O�a<��a<�a<��a<A�a<�	b<�b<�b<�a<L�a<N�a<n�a<xIa<�a<R�`<b�`<}`<�c`</Z`<�a`<7y`<�`<��`<�a<-Ba<pza<�a<%�a<�a<�b< b<�b<��a<d�a<��a<�a<O�a<B�a<��a<k�a<F�a<��a<"�a<'�a<��a<��a<1�a<Yb<{b<u�a<��a<��a<V�a<�ia<�0a<�`<-�`<^�`<Im`<Y`<'U`<b`<�~`<_�`<��`<�a<Oa<��a<�a<!�a<��a<b<`b<��a<V�a</�a<�a<�a<��a<]�a<��a<V�a<�a<	�a<A�a<J�a<��a<f�a<��a<��a<��a<U�a<��a<s�a<�ua<�>a<ha<��`<|�`<{g`<XH`<�8`< :`<�K`<�l`<��`<�`<�a<�Aa<Bva<o�a<��a<A�a<��a<�a<�a<��a<�a<��a<��a<�a<ςa<�~a<�a<Ņa<�a<�a<3�a<g�a<��a<�a<�a<��a<��a<�a<Ƃa<�Pa<�a<��`<W�`<_s`<L`<�2`<W)`<�0`<�H`<�n`<՟`<�`<�a<�  �  `7a<yna<�a<]�a<��a<��a<k�a<��a<��a<��a<,�a<�a<��a<d�a<^�a<�a<��a<n�a<��a<B�a<��a<��a< �a<�a<��a<V�a<<�a<?ma<b5a<��`<��`<��`<*O`<�*`<�`<|`<V!`<�@`<qn`<Ϧ`<�`<�$a<�`a<��a<M�a<��a<��a<@�a<��a< �a< �a<��a<M�a<��a<��a<q�a<=�a<`�a<��a<��a<�a<V�a<s�a<ab<{b<|b<[�a<�a<�a<�~a<bDa<+a<��`<��`<Ab`<#B`<32`<E4`<�G`<{k`<s�`<B�`<�a<hRa<��a<Y�a<S�a<��a<�
b<ub<�b<�b<��a<��a<�a<_�a<��a<�a<��a<��a<W�a<}�a<:�a<��a<	b<�b<<b<sb<��a<��a<ʣa<�ma<�1a<��`<n�`<̀`<�V`<�;`<�1`<�9`<�R`<{`<��`<"�`<�)a<]fa<�a<7�a<F�a</b<�b<;b<b<��a<h�a<n�a<��a<��a<?�a<��a<��a<��a<��a<y�a<^�a<2�a<Lb<�b<@b<��a<�a<3�a<}�a<�Ta<ba<��`<�`<�k`<nF`<�0`<�,`<�:`<�X`<��`<Ҽ`<��`<.8a<�ra<q�a<��a<O�a<��a<�b<�b<8�a<q�a<0�a<��a<��a<��a<��a<v�a<��a<(�a<��a<��a<z�a<��a<�a<��a<	�a<g�a<��a<M�a<tca< (a<��`<@�`<q`<�A`<� `<F`<�`<�$`<�G`<�w`<:�`<�`<P,a<�da<3�a<��a<G�a<�a< �a<��a<@�a<��a<Z�a<
�a<�a<��a<'�a<֢a<æa<��a<ҷa<N�a<|�a<��a<�a<q�a<w�a<��a<|�a<Gsa<=a<� a<��`<z�`<�O`<�%`<�
`<� `<�`<:"`<�J`<�`<y�`<��`<�  �  X*a<�ca<�a<ڸa<��a<��a<��a<��a<��a<4�a<��a<F�a<�a< �a<t�a<I�a<��a<�a<x�a<��a<?�a<��a<��a<E�a<�a<I�a<͓a<&ba<�'a<)�`<ʧ`<vk`<8`<�`<��_<��_<�`<�(`<3X`<ْ`<��`<�a<~Ta<�a<;�a<��a<��a<��a<z�a<6�a<a�a<D�a<��a<��a<��a<R�a<+�a<o�a<��a<��a<��a<��a<�b<tb<_b<�b<��a<5�a<��a<�ra<�5a<��`<��`<|z`<�J`<�(`<@`<O`</`<-T`<�`<(�`<�a<�Da<8�a<��a<�a<��a<�	b<�b<db<�
b<^b<i�a<]�a<L�a<5�a<��a<K�a<��a<��a<7�a<�a<b<mb<�b<Eb<�b<��a<E�a<��a<aa<"a<��`<�`<,j`<�>`<"`<�`<�`<P:`<@d`<��`<��`<a<RYa<��a<_�a<��a<?�a<�b<�b<b<�b<��a<��a<�a<y�a<��a<��a<�a<��a<��a<N�a<�a<�b<�b<�b<tb<u�a<��a<Ǵa<f�a<QGa<�a<��`<Ј`<�T`<�-`<�`<�`<!`<�@`<To`<ڨ`<b�`<I)a<�fa<Μa<��a<��a<��a<eb<Ob<Nb<��a<��a<O�a<��a<��a<h�a<d�a<��a<��a<J�a<��a< �a<Q�a<3�a<�a<i�a<�a<ӹa<��a<�Wa<�a<��`<��`<[`<9*`<�`<U�_<��_<�`<G0`<tb`< �`<[�`<ga<�Ya<u�a<S�a<z�a<�a<��a<}�a<^�a<^�a<��a<V�a<ʾa<B�a<8�a<��a<k�a<p�a<��a<&�a<��a<
�a<��a<z�a<��a<V�a<�a<ia<c0a<Z�`<�`<�p`<69`<�`<$�_<��_</�_<�	`<	4`<�j`<:�`<��`<�  �  �%a<`a<0�a<��a<��a<��a<��a<��a<��a<��a<�a<a�a<��a<#�a<��a<Z�a<]�a<��a<��a<��a<��a<��a<w�a<'�a<��a<ܷa<��a<!^a<�"a<p�`<V�`<d`<�/`<P	`<�_<��_<!�_<� `<�P`<�`<��`<ua<)Pa<��a<��a<��a<��a<�a<��a<r�a<��a<�a<C�a<"�a<��a<��a<a�a<g�a<y�a<C�a<��a<nb<9	b<�b<�b<Vb<'�a<��a<U�a<Sna<�0a<��`<4�`<�r`<{B`< `<�`<�`<Z&`<L`<|`<��`<�`<�?a<|a<j�a<��a<)�a<�	b<�b<b<Yb<,b<��a<$�a<��a<C�a<��a<y�a<^�a<�a<��a<�b<b<qb<�b<hb<�b<`�a<j�a<̕a<�\a<�a<��`<Ú`<cb`<?6`<B`<�`<`<�1`<b\`<z�`<��`<�a<�Ta<��a<t�a<��a<&�a<�b<�b<b<�	b<Gb<I�a<:�a<M�a<�a<�a<!�a<��a<j�a<��a<"b<M	b<[b<fb<Wb<�a<��a<��a<b~a<�Ba<Aa<n�`<c�`<�L`<%`<`<
`<L`<�8`<�g`<�`<N�`<�#a<\ba<O�a<��a<��a<�a<�b<�b<�b<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<��a<5�a<)�a<��a<JSa<Ya<��`<ŏ`<�S`<)"`<��_<��_<��_<`<7(`<[`<��`<��`<xa<zUa<B�a<бa<��a<��a<0�a<,�a<��a<+�a<��a<�a<o�a<N�a<��a<��a<G�a<��a<	�a<��a<��a<�a<��a<��a<��a<6�a<�a<Nea<�+a<��`<��`<�i`<o1`<N`<`�_<5�_<d�_<�`<-,`<�c`<��`<7�`<�  �  X*a<�ca<�a<ڸa<��a<��a<��a<��a<��a<4�a<��a<F�a<�a< �a<t�a<I�a<��a<�a<x�a<��a<?�a<��a<��a<E�a<�a<I�a<͓a<&ba<�'a<)�`<ʧ`<vk`<8`<�`<��_<��_<�`<�(`<3X`<ْ`<��`<�a<~Ta<�a<;�a<��a<��a<��a<z�a<6�a<a�a<D�a<��a<��a<��a<R�a<+�a<o�a<��a<��a<��a<��a<�b<tb<_b<�b<��a<5�a<��a<�ra<�5a<��`<��`<|z`<�J`<�(`<@`<O`</`<-T`<�`<(�`<�a<�Da<8�a<��a<�a<��a<�	b<�b<db<�
b<^b<i�a<]�a<L�a<5�a<��a<K�a<��a<��a<7�a<�a<b<mb<�b<Eb<�b<��a<E�a<��a<aa<"a<��`<�`<,j`<�>`<"`<�`<�`<P:`<@d`<��`<��`<a<RYa<��a<_�a<��a<?�a<�b<�b<b<�b<��a<��a<�a<y�a<��a<��a<�a<��a<��a<N�a<�a<�b<�b<�b<tb<u�a<��a<Ǵa<f�a<QGa<�a<��`<Ј`<�T`<�-`<�`<�`<!`<�@`<To`<ڨ`<b�`<I)a<�fa<Μa<��a<��a<��a<eb<Ob<Nb<��a<��a<O�a<��a<��a<h�a<d�a<��a<��a<J�a<��a< �a<Q�a<3�a<�a<i�a<�a<ӹa<��a<�Wa<�a<��`<��`<[`<9*`<�`<U�_<��_<�`<G0`<tb`< �`<[�`<ga<�Ya<u�a<S�a<z�a<�a<��a<}�a<^�a<^�a<��a<V�a<ʾa<B�a<8�a<��a<k�a<p�a<��a<&�a<��a<
�a<��a<z�a<��a<V�a<�a<ia<c0a<Z�`<�`<�p`<69`<�`<$�_<��_</�_<�	`<	4`<�j`<:�`<��`<�  �  `7a<yna<�a<]�a<��a<��a<k�a<��a<��a<��a<,�a<�a<��a<d�a<^�a<�a<��a<n�a<��a<B�a<��a<��a< �a<�a<��a<V�a<<�a<?ma<b5a<��`<��`<��`<*O`<�*`<�`<|`<V!`<�@`<qn`<Ϧ`<�`<�$a<�`a<��a<M�a<��a<��a<@�a<��a< �a< �a<��a<M�a<��a<��a<q�a<=�a<`�a<��a<��a<�a<V�a<s�a<ab<{b<|b<[�a<�a<�a<�~a<bDa<+a<��`<��`<Ab`<#B`<32`<E4`<�G`<{k`<s�`<B�`<�a<hRa<��a<Y�a<S�a<��a<�
b<ub<�b<�b<��a<��a<�a<_�a<��a<�a<��a<��a<W�a<}�a<:�a<��a<	b<�b<<b<sb<��a<��a<ʣa<�ma<�1a<��`<n�`<̀`<�V`<�;`<�1`<�9`<�R`<{`<��`<"�`<�)a<]fa<�a<7�a<F�a</b<�b<;b<b<��a<h�a<n�a<��a<��a<?�a<��a<��a<��a<��a<y�a<^�a<2�a<Lb<�b<@b<��a<�a<3�a<}�a<�Ta<ba<��`<�`<�k`<nF`<�0`<�,`<�:`<�X`<��`<Ҽ`<��`<.8a<�ra<q�a<��a<O�a<��a<�b<�b<8�a<q�a<0�a<��a<��a<��a<��a<v�a<��a<(�a<��a<��a<z�a<��a<�a<��a<	�a<g�a<��a<M�a<tca< (a<��`<@�`<q`<�A`<� `<F`<�`<�$`<�G`<�w`<:�`<�`<P,a<�da<3�a<��a<G�a<�a< �a<��a<@�a<��a<Z�a<
�a<�a<��a<'�a<֢a<æa<��a<ҷa<N�a<|�a<��a<�a<q�a<w�a<��a<|�a<Gsa<=a<� a<��`<z�`<�O`<�%`<�
`<� `<�`<:"`<�J`<�`<y�`<��`<�  �  nKa<j~a<ݧa<!�a<E�a<��a<��a<i�a<X�a<2�a<̠a<��a<�a<Ła<!�a<��a<p�a<��a<`�a<Ѹa<��a<��a<w�a<W�a<�a<�a<�a<~a<cJa<�a<��`<ѡ`<�s`<xQ`<>`<;`<�H`<mf`<8�`<��`<  a<~;a<Tsa<E�a<��a<��a<��a<��a<��a<<�a<��a<��a<j�a<�a<g�a<l�a<�a<��a<��a<��a<d�a<��a<��a<� b<�b<Tb<K�a<�a<8�a<��a<�Za<� a<N�`<�`<Ӈ`<�i`<�Z`<�\`<�n`<j�`<��`<�`<I.a<�ga<ߜa<��a<i�a<vb<�b<nb<�b<��a<�a<�a<��a<��a<��a<?�a<ʭa<ѳa<O�a<��a<�a<��a<A�a<�	b<�b<�b<�a<L�a<N�a<n�a<xIa<�a<R�`<b�`<}`<�c`</Z`<�a`<7y`<�`<��`<�a<-Ba<pza<�a<%�a<�a<�b< b<�b<��a<d�a<��a<�a<O�a<B�a<��a<k�a<F�a<��a<"�a<'�a<��a<��a<1�a<Yb<{b<u�a<��a<��a<V�a<�ia<�0a<�`<-�`<^�`<Im`<Y`<'U`<b`<�~`<_�`<��`<�a<Oa<��a<�a<!�a<��a<b<`b<��a<V�a</�a<�a<�a<��a<]�a<��a<V�a<�a<	�a<A�a<J�a<��a<f�a<��a<��a<��a<U�a<��a<s�a<�ua<�>a<ha<��`<|�`<{g`<XH`<�8`< :`<�K`<�l`<��`<�`<�a<�Aa<Bva<o�a<��a<A�a<��a<�a<�a<��a<�a<��a<��a<�a<ςa<�~a<�a<Ņa<�a<�a<3�a<g�a<��a<�a<�a<��a<��a<�a<Ƃa<�Pa<�a<��`<W�`<_s`<L`<�2`<W)`<�0`<�H`<�n`<՟`<�`<�a<�  �  da<_�a<��a<�a<[�a<n�a<M�a<��a<�a<S�a<�~a<2ka<]\a<tSa<1Qa<�Ua<�`a<lqa<��a<V�a<��a<M�a<.�a<"�a<N�a<��a<�a<K�a<=da<1a<��`<��`<W�`<l�`<�q`<^o`<�{`<��`<K�`<)�`<"a<�Wa<�a<l�a<��a<{�a<#�a<K�a<4�a<S�a<K�a<��a<k�a<�a<�wa<�qa<Sra<�ya<+�a<��a<��a<8�a<Y�a<��a<Ob<b<Kb<r�a<��a<�a<nva<"Ba<a<x�`<��`<M�`<��`<��`<?�`<x�`<��`<�a<9Na<P�a<��a<��a<��a<Fb<b<�b<P�a<��a<=�a<�a<�a<@�a<��a<N}a<Ga<Շa<r�a<٩a<��a<n�a<��a<f b<�
b<"b<��a<o�a<��a<u�a<�fa<2a<��`<��`<�`<�`<��`<:�`<��`<��`<��`<�+a<6`a<�a<	�a<��a<j�a<�b<�	b< b<(�a<��a<��a<�a<��a<��a<<}a<oza<K~a<ƈa<Ԙa<O�a<^�a<��a<��a< b<>b<�b<D�a<��a<��a<��a<�Oa<a<:�`<�`<@�`<�`<��`<
�`<�`<x�`<5a<�6a<Jka<[�a<B�a<�a<L�a<[b<��a<�a<p�a<��a<�a<�a<܃a<�ua<�ma<�la<�qa<�}a<��a<��a<Y�a<��a<[�a<i�a<��a<Q�a<�a<�a<Ջa<$Za<�$a<��`<�`<X�`<{`<m`<�m`<�}`<��`<�`<��`<�(a<;\a<�a<۱a<��a<�a<N�a<��a<}�a<h�a<T�a<�a<ra<�`a< Ua<Pa<�Qa<�Ya<ha<9{a<��a<J�a<~�a<��a<��a< �a<��a<�a<�a<�ha<6a<a<��`<|�`<}`<
f`<�]`<}d`<z`<Z�`<��`<��`<�0a<�  �  �~a<5�a<��a<��a<=�a<�a<�a<�a<�a<Hsa<�Ua<�;a<G(a<�a<�a<Ra<�-a<ZCa<�^a<�}a<W�a<P�a<��a<�a<��a<1�a<��a<��a<<�a<�Sa<;&a<~�`<�`<.�`<�`<�`<ߵ`<R�`<c�`<[a<�Ga<�va<`�a<�a<)�a<��a<��a<��a<��a<=�a<�a<��a<ja<�Ra<�Ba<Z:a<�:a<Da<�Ua<�ma<L�a<8�a<|�a<$�a<�a<�b<�b<5�a<��a<l�a<��a<�fa<�9a<a<��`<�`<u�`<��`<]�`<��`<�a<�Ca<�qa<�a<��a<{�a<��a</	b<�b<��a<�a<D�a<��a<�a<|pa<�Za<�Ka<�Ea<1Ha<SSa<pfa<�a<��a<��a<\�a<c�a<�b<Mb<ab<:�a<��a<I�a<\�a<Ya<^,a<�a<��`<��`<G�`<�`<��`<q a<'a<ISa<i�a<��a<��a<K�a<�b<�	b<1b<��a<u�a<�a<ߞa<��a<�fa<�Ra<cFa<�Ba<�Ga<�Ua<�ja<��a<�a<��a<��a<k�a<#b<�b<��a<��a<��a<��a<�ra<RDa<�a<��`<�`<�`<
�`<�`<��`<�a<m/a<u\a<+�a<��a<��a<��a<t�a<b<O�a<i�a<]�a<k�a<|�a<�ka<�Ra<�@a<r6a<5a<k<a<
La<�ba</~a<W�a<�a<��a<�a<��a<��a<��a<��a<S�a<Bxa<�Ia<a<��`<��`<ܴ`<|�`<B�`<
�`<��`<X�`<�a<La<�xa<�a<a�a<;�a<�a<��a<��a<U�a<�a<�a<`a<�Da<#.a<a<�a<�a<Y%a<#8a<FQa<�na<��a<��a<��a<��a<H�a<)�a<��a<<�a<��a<yVa<(a<L�`<��`<��`<��`<V�`<K�`<��`<�`<�`<�#a<�Qa<�  �  -�a<��a<t�a<e�a<@�a<�a<*�a<��a<sa<RLa<W'a<ha<�`<j�`<^�`<��`<8�`<7a<32a<�Xa<�a<��a<;�a<��a<%�a<U�a<��a<��a<��a<�va<cPa<�,a<a<��`<,�`<w�`<��`<�a<U#a<�Fa<�ma<[�a<��a<8�a<H�a<!�a<��a<w�a<!�a<V�a<T�a<~\a<�9a<�a< a<��`<��`<?	a<�a<�<a<aa<��a<��a<��a<��a<b<�b<�b<)�a<��a<��a<{�a<!fa<JCa<�&a<�a<�a<5
a<Xa<P,a<�Ja<�na<b�a<$�a<��a<C�a<�b<�	b<� b<Q�a<0�a<��a<(�a<`a<�=a<�"a<ca<ya<�a<�a<[1a<�Pa<�ua<Ȝa<*�a<��a<��a<�b<^
b<��a<��a<�a<֧a<�a<;[a<
:a<�a<=a<�a<�a<Ka<M6a<�Va<�{a<��a<C�a<^�a<��a<Tb<�b<A�a<��a<�a<��a<�wa<wRa<2a<Ba<
a<�a<$a<(a<�7a<�Xa<�~a<1�a<�a<��a<��a<sb<�b<��a<��a<��a<t�a<yna<�Ia<�*a<�a<7a<�a<a<�a<�:a<�\a<˂a<��a<��a<�a<��a<�b<��a<�a<�a<y�a<��a<`a<];a<}a<a<��`<�`<�a<2a<�1a<�Sa<�ya<�a<��a<�a<��a<��a<�a<V�a<��a<2�a<oa<�Ga<�#a<:a<��`<��`<��`<�`<aa<"&a<�Ia<�oa<�a<�a<.�a<�a<c�a<R�a<�a<r�a<n�a<W[a<�4a<$a<I�`<��`<H�`<�`<��`<a<]"a<�Fa<�ma<Βa<�a<�a<��a< �a<�a<�a<N�a<�va<�Oa<*a<�a<��`<"�`<��`<�`<��`<�a<�&a<-La<Bsa<�  �  !�a<6�a<��a<��a<2�a<=�a<R�a<�}a<QQa<H#a<d�`<J�`<-�`<��`<ǝ`<4�`<?�`<R�`<�a<41a<�_a<:�a<�a<i�a<��a<r�a<��a<��a<�a<�a<�xa<�[a<{Ca<�1a<�'a<�&a<,.a<(>a<oUa<ra<Αa<n�a<�a<r�a<v�a<f�a<V�a<G�a<�a<��a<^a<01a<�a<��`<��`</�`<n�`<��`<?�`<�	a<�4a<�ca<?�a<�a<
�a<�a<b<�b<��a<��a<��a<��a<̐a<�ta<�]a<�Ma<Fa<�Fa<�Pa<Nba<�za<��a<��a<��a<�a<b<�	b<�b<o�a<��a<��a<u�a<h_a<M2a<�	a<�`<4�`<��`<��`<D�`<��`<7 a<�Ka<=za<R�a<��a<K�a<�b<2b<�b<X�a<E�a<��a<¦a<W�a<�ma<�Xa<*Ka<SFa<Ja<XVa<vja<��a<��a<`�a<>�a<��a<Ub<�	b<�b<c�a<�a<�a<A}a<�Na<y"a<��`<P�`<7�`<��`<��`< �`<�a<X*a<Wa<�a<��a<��a<f�a<�b<b<��a<��a<��a<׵a<��a<3ya<`a<sMa<�Ba<�@a<sGa<tVa<�la<-�a<��a<�a<W�a<X�a<� b<Eb<��a<��a<̻a<�a<wca<�4a<8	a<��`<��`<H�`<��`<�`<��`<��`<�'a<�Ta<��a<��a<�a<��a<�a<��a<��a<^�a<g�a<�a<?ra<5Ua<U=a<�,a<$a<D$a<@-a<\>a<Va<�ra<�a<��a<��a<�a<��a<��a<��a<��a<ߎa<8ca<�4a<a<��`<̼`<{�`<��`<�`<]�`<V�`<��`<"a<$Ka<�wa<c�a<x�a<��a<��a<C�a<��a<p�a<��a<�ua<)Wa<Z<a<X'a< a<Da<%a<�%a<:a<hTa<�ra<�a<�  �  b�a<��a<�a<��a<��a<v�a< �a<�ba<�/a<*�`<��`<L�`<�{`<�g`<6b`<�k`<��`<k�`<��`<�
a<�?a<�ra<0�a<��a<a�a<��a<M�a<6�a<�a<�a<��a<'�a<�sa<=fa<�^a<&^a<da<�pa<��a<��a<�a<�a<��a<��a<��a<�a<��a<e�a<��a<�ma<a:a<�a<��`<M�`<��`<݃`<�`<+�`<P�`<��`<�	a<?a<�ta<ԥa<t�a<��a<b<f	b<Qb<q�a<�a<��a<��a<-�a<��a<k�a<�}a<M~a<��a<%�a<��a<ٻa<��a<F�a<��a<Kb<v
b<b<��a<��a<�a<.na<|9a<�a<A�`<(�`<��`<@�`<��`<��`<�`<��`<#a<�Wa<��a<�a<��a<��a<M	b<)b<Yb<��a<`�a<��a<{�a<�a<�a<��a<�}a<ǀa<D�a<��a<k�a<:�a<��a<��a<�b<i
b<�b<4�a<��a<ܼa<%�a<�[a<�&a<��`<��`<�`<B�`<<�`<.�`<«`<��`<�`<f0a<ea<5�a<��a<��a<��a<1b<"b<\�a<y�a<��a<�a<��a<e�a<�a<�ya<]xa<e}a<�a<˙a<Ѯa<��a<.�a<�a<��a<�b<��a<��a<�a<m�a<�ta<�?a<N
a<��`<&�`<��`<�`<;~`<��`<Ѧ`<d�`<��`<40a<�ca<��a<��a<*�a<�a<��a<u�a<H�a<��a<u�a<�a<��a<?oa<$ba<�[a<�[a<?ba<0oa<+�a<ϖa<�a<:�a<.�a<?�a<��a<�a<	�a<��a<9va<�Ca<�a<z�`<��`<�`<Kl`<&a`<	e`<�w`<ۗ`<d�`<?�`<�(a<V\a<{�a<��a<��a<�a<��a<��a<��a<[�a<{�a<Aa<�ja<�Za<oPa<�La<�Oa<�Ya<ia<8}a<Z�a<`�a<�  �  ��a<K�a<A�a<c�a<��a<~�a<�|a<�Ia<xa<�`<��`<uo`<�J`<4`<�-`<|8`<$S`<�{`<l�`<��`<�"a<![a<(�a<)�a<��a<z�a<��a<��a<��a<��a<߸a<0�a<؛a<`�a<o�a<	�a<��a<��a<��a<v�a<q�a<F�a<	�a<�a<��a<��a<2�a<��a<[�a<�Ra<a<��`<�`<�`<M``<�O`<�O`<�``<��`<t�`<Z�`<&a<+Ya<�a<*�a<��a<g�a<	b<�
b<b<�a<��a<��a<�a<Q�a<��a<k�a<��a< �a<ûa<^�a<t�a<��a<��a<�b<xb<�b<1�a<`�a<8�a<��a<�Qa</a<	�`<ݪ`<��`<�e`<�Y`<�^`<�s`<��`<�`<X�`<�8a<!ra<4�a<G�a<S�a<]b<�b< b<\b<��a<�a<��a<��a<��a<��a<�a<�a<��a<��a<:�a<��a<��a<��a<
b<�b<Xb<��a<��a<��a<2va<\=a<�a<��`< �`<�t`<�]`<�V`<�``<�z`<��`<��`<xa<�Ga<za<ɰa<�a<�a<�b<�b<�b<9�a<]�a<��a<��a<�a<E�a<��a<E�a<��a<�a<D�a<��a<i�a<��a<d�a<b<8b<��a<~�a<P�a<G�a<Za<xa<r�`<ԭ`<�`<G^`<�K`<J`<�X`<(w`<�`<7�`<=a<�Ha<�}a<3�a<�a<Y�a<��a<�a<��a<��a<%�a<#�a<��a<٘a<_�a<_�a<=�a<��a<̗a<ڤa<j�a<&�a<��a<s�a<p�a<R�a<%�a<жa< �a< _a<y'a<�`<ղ`<(`<}U`<<9`<�,`<:1`< F`<�i`<��`<��`<�	a<�Ba<�va<q�a<A�a<�a<3�a<H�a<u�a<��a<Q�a<a�a<E�a<��a<z~a<�{a<~a<�a<�a<��a<�a<i�a<�  �  ��a<��a<��a<��a<��a<X�a<�la<�5a<��`<R�`<`<[K`<�#`<`<C`<�`<�,`<1X`<Ɏ`<��`<Ka<�Ga<�}a<�a<��a<��a<o�a<
�a<��a<��a<@�a<T�a<�a<��a<@�a<=�a<��a<C�a<�a<��a<�a<��a<M�a<��a<��a<��a<��a<8�a<�ua<@=a<, a<��`<^�`<�Z`<,9`<e'`<X'`<;9`<A[`<J�`<��`<�a<Ca<
~a<C�a<��a<��a<vb<'b<�b<�b<��a<��a<��a<��a<��a<��a<��a<��a<a�a<�a<Z�a<��a<fb<�b<�b<Pb<��a<��a<U�a<�ua<�:a<��`<Ͼ`<݇`<�[`<=>`<E1`<�6`<M`<?s`<.�`<(�`< a<Z]a<��a<��a<��a<b<�b<�b<�b<Sb<>�a<>�a<��a<K�a<2�a<*�a<��a<D�a<�a<^�a<�a<# b<�	b<Tb<(b<~b<��a<z�a<i�a<�aa<�$a<��`<�`<�u`<�M`<�5`<4.`<9`<�T`<I`<5�`<��`<R0a<la<z�a<��a<�a<b<<
b<)
b<Db<��a<V�a<��a<��a<l�a<Y�a<|�a<�a<��a<\�a<�a<
�a<_�a<�b<�b<1b<��a<.�a<ܰa<�~a<mDa<�a<v�`<�`<�Z`<&7`<~#`<�!`<�1`<�Q`<�`<Է`<��`<`2a<�ka<J�a<Q�a<��a<��a<C�a<��a<w�a<:�a<�a<"�a<!�a<D�a<��a<1�a<-�a<h�a<}�a<O�a<�a<\�a</�a<��a<��a<��a<�a<D�a<2La<`a<$�`<��`<1\`<�/`<�`<;`<	`<@`<E`<�w`<`�`<��`<.a<�ea<ڔa<˸a<��a<4�a<�a<��a<=�a<�a<�a<?�a<�a<�a<��a<��a<q�a<��a<�a<#�a<��a<�  �  p�a<��a<e�a<s�a<W�a<^�a<ba<j(a<��`<��`<5j`<z4`<�`<1�_<C�_<�_<�`<�A`<iz`<�`<��`<(;a<�sa<��a<��a<�a<��a<%�a<g�a<��a<K�a<4�a<��a<E�a<�a<H�a<��a<�a<3�a<N�a<B�a<��a<��a<-�a<��a<��a<l�a<R�a<Tja<,/a<`�`<��`<�t`<�C`<1 `<q`<g`< `<�C`<^u`<i�`<��`<�4a<Fra<�a<*�a<{�a<�b<4b<b<�b<�b<��a<��a<�a<��a<��a<��a<t�a<S�a<3�a<��a<�b<Ob<0b<b<4b<��a<k�a<��a<�ia<t+a<6�`<��`<�q`<�C`<�$`<H`<�`<i4`<.\`<�`<��`<�a<�Oa<��a<k�a<��a<��a<b<�b<3b<�
b<,b<6�a<T�a<��a<��a<I�a<9�a<��a<�a<��a<^ b<	b<�b<�b<�b<j�a<��a<�a<��a<�Ta<�a<`�`<-�`<�^`<�5`<�`</`<i`<�<`<�h`<Р`<��`<� a<t_a<`�a<f�a<��a<��a<j
b<Bb<�	b<gb<`�a<��a<]�a<-�a<�a<��a<G�a<h�a<��a<��a<A�a<Vb<[
b<#
b<�b<��a<��a<��a<Csa<Z6a<��`<5�`<lv`<hC`<,`<�	`<�`<j`<%:`<j`<D�`<��`<�#a<�_a<�a<��a<i�a<x�a<M�a<��a<�a<�a<'�a<��a<��a<c�a<�a<
�a<�a<Y�a<��a<��a<-�a<G�a<��a<�a<��a<��a<�a<{wa<�?a<Wa<��`<�`<�E`<�`<�_<C�_<)�_<�`<	.`<�b`<��`<��`<� a<[a<��a<�a<f�a<��a<�a<B�a<��a<��a<��a<��a<%�a<V�a<�a<,�a<ҹa<��a<W�a<l�a<��a<�  �  �b<H
b<�b<y�a<�a<&�a<�`a<.a<|�`<�b`<�`<��_<_<�f_<�\_<m_<2�_<|�_<�"`<zz`<��`<�*a<Yva<^�a<��a<C b<Mb<�b<�b<�
b<b<n�a<��a<�a<'�a<��a<f�a<��a<�a<�b<�b<�b<�b<� b<�b<Db<?�a<��a<Yca<a<R�`<Ic`<x`<��_<+�_<�_<��_<��_<;�_<`<�b`<u�`<ya<�ia<d�a<��a<b<�+b<�7b<9b<�3b<�+b<4$b<gb<�b<b<b<b<[b<mb<bb<r%b<p-b<R5b<q9b<�6b<�(b<�b<W�a<��a<�[a<�a<�`<qV`<G`<w�_<X�_<�_<'�_<��_<Q�_<�2`<��`<<�`<�8a<�a<[�a<n�a<�b<�3b<�:b<�9b<�2b<Z*b<�"b<hb<�b<$b<�b<�b<�b<`b<N!b<�(b<�0b<�7b<�9b<�3b<&!b<Z b<��a<�a<#@a<�`<�`<@9`<#�_<s�_<֐_<��_<�_<��_<2�_<�I`<ɠ`<W�`<�Oa<x�a<��a<7b<E"b<�1b<b5b<�1b<*b<�!b<�b<$b<�b<b<�b<�b<Bb<Zb<�b<%b<y-b<3b<�2b<)(b<�b<3�a<�a<�la<�a<�`<g`<_`<��_<)�_<}_<�z_<�_<h�_<Z`<+U`<��`</a<�Va<��a< �a<�a<rb<�b<�b<lb<Ob<�b<��a<e�a<��a<��a<P�a<�a<��a<�a<��a<&b<�b<Bb<�b<c b<Y�a<6�a<�{a<�1a<��`<��`<�*`<��_<��_<o_< \_<�b_<p�_<l�_<y`<X`<m�`<�a<�Wa<��a<��a<��a<Cb<U	b<�b<� b<(�a<w�a<�a<3�a<��a<d�a<��a<�a<��a<�a<��a<Y b<�  �  �b<�	b<5b<��a<k�a<��a<-fa<ea<�`<�k`<�`<��_<q�_<�r_<i_</y_<ˡ_<D�_<�,`<��`<��`<�0a<�{a<y�a<��a<*b<�b<�b<�b<!b<��a<h�a<\�a<��a<4�a<��a<��a<�a<��a<� b<Ub<Fb<:b< b<(b<�b<��a<~�a<ia<�a<Y�`<jl`<�`<�_<�_<=�_<ь_<�_<��_<{`<l`<��`<&a<�oa<]�a<7�a<�b<S-b<7b<�7b<i1b<�'b<*b<�b<(b<|b<�
b<b<�b<�b<7b<�b<�)b<3b<J8b<�6b<C*b<�b<P�a<̪a<�aa<�a<g�`<�_`<�`< �_<e�_<�_<P�_<��_<k�_<�<`<s�`<��`<G?a<��a<��a<� b<;"b<�4b<e:b<�7b<�/b<�%b<+b<~b<wb<_b<b<b<�b<Sb<�b<�#b<�-b<�5b<'9b<S4b<]#b<�b<Z�a<��a<[Fa<��`<ԗ`</C`<&�_<$�_<��_<��_<4�_<.�_<�`<�S`<K�`<�a<�Ua<͟a<��a<Eb<,$b<�1b<g4b<�/b<�&b<ub<�b<�b<{b<%b<�b< b<[
b<�b<�b<:!b<�*b<s1b<C2b<c)b<pb<��a<��a<sra<*!a<�`<?p`<�`<��_<�_<E�_<�_<�_<��_<�`<m^`<!�`<�a<u\a<��a<��a<��a<�b<�b<Ob<�b<B	b<x�a<M�a<��a<!�a<��a<G�a<��a<	�a<��a<��a<xb<Gb<b<b<"b<K�a<-�a<"�a<�7a<��`<�`<4`<��_<'�_<{_<@h_<#o_</�_<��_<�`<�``<$�`<1a<8]a<H�a<��a<�a<%b<�b<�b<��a<s�a<��a< �a<�a<	�a<E�a<��a<��a<��a<Z�a<��a<F�a<�  �  ��a<'b<xb<_�a<(�a<f�a<kua<�+a<�`<��`<�3`<[�_<�_<�_<��_<&�_<	�_<�_<>H`<��`<5�`<kBa<,�a<��a<��a<!b<$b<Ub<b<��a<v�a<��a<��a<o�a<?�a<T�a<��a<0�a<L�a<U�a<��a<b<�b<f b<�b<�b<��a<v�a<Uya<9-a<t�`<��`<<9`<G�_<T�_<��_<J�_<f�_<�_<S8`<��`<�`<51a<.�a<��a<M�a<�b<+1b<�7b<�3b<�(b<�b<cb<# b<��a<��a<��a<��a<^�a<�a<@b<b<�b<f+b<[5b<�7b<�.b<�b<#�a<��a<@sa<s#a<��`<V{`<s0`<�_<?�_<��_<��_<��_<!`<�Y`<�`<T�`<&Ra<*�a<�a<�	b<A(b</7b<k9b<2b<�%b<�b<�b<V�a<��a<��a<�a<P�a<��a<��a<�b<kb<#b<�/b<�7b<�6b<)b<eb<6�a<Ϣa<�Xa<�a<�`<�_`<�`<��_<4�_<T�_<3�_<s�_<�%`<Mo`<��`<�a<Mga<S�a<�a<Xb<')b<~3b<2b<�(b<�b<9b<��a<T�a<"�a<.�a<p�a<��a<r�a<��a<lb<zb<�!b<�,b<'2b<�,b<,b<��a<��a<a<�4a<.�`<��`<";`<;�_<S�_<��_<\�_<��_<E�_<�,`<y`<��`<�a<#ma<��a<��a<�b<�b<�b<Mb<Nb<�a<��a<{�a<	�a<-�a<��a<-�a<�a</�a<��a<D�a<U�a<�b<)b<0b<�b<	�a<��a<J�a<Ia<��`<P�`<{O`<`<(�_<�_<Ӌ_<r�_<�_<7�_<P*`<�z`<��`<"a<�la<��a<�a<"�a<�b<�b<A b<��a<��a<��a<��a<��a<��a<ٻa<J�a<�a<9�a<��a<��a<��a<�  �  �a<�b<H	b<�b<��a<1�a<�a<�Ga<D�`<�`<v``<�`<9�_<K�_<��_<�_<`�_<i.`<�s`<2�`<Oa<F]a<��a<j�a<(�a<Ub<�b<�b<$�a<��a<��a<�a<�a<��a<G�a<ڝa<Ӣa<%�a<��a<{�a<��a<��a<Ob<5b<O b<�b<�a<��a<��a<Ka<��`<��`<}g`<+`<b�_<\�_< �_<��_<:*`<g`<T�`<��`<�Oa</�a<��a<Yb<�&b<w5b<I6b<�+b<�b<�b<N�a<�a<
�a<��a<4�a<��a<�a<��a<��a<��a<L	b<?b<
/b<�7b<y4b<�"b<c b<��a<��a<Ca<��`<*�`<U``<(`<`<��_<�_<`<F`<��`<��`<4!a<�na<b�a<`�a<-b<-0b<�9b<�5b<(b<]b<�a<x�a<P�a<��a<v�a<w�a<��a<7�a<�a<��a<K�a<b<�$b<s3b<a8b<g0b<b<�a<s�a<�ta<�'a<(�`<-�`<�I`<�`<��_<b�_<,�_<�`<5V`<��`<��`<�6a<2�a<��a<��a<�b<b/b<�3b<f,b<2b<bb<��a<1�a<z�a<��a<3�a<�a<�a<b�a<��a<��a<��a<b<�$b<�/b<�0b<Q#b<�b<��a<,�a<�Ra<8a<��`<ai`<�*`<`�_<c�_<1�_<��_<i `<`[`<��`<E�`<O>a<&�a<��a<��a<�b<b<lb<�b<��a<)�a<��a<y�a<��a<��a<&�a<�a<1�a<Ȫa<_�a<��a<�a<��a<�b<	b<Pb<��a<5�a<0�a<Aca<6a<R�`<Dz`<�3`<�_<��_<��_<��_<��_<`<mW`<<�`<_�`<�>a<�a<ļa<Q�a<�a<?b<=b<O�a<f�a<a�a<=�a<�a<s�a<4�a<Q�a<��a<w�a<��a<z�a<��a<��a<�  �  ��a<��a<	b<�b<$�a<;�a<��a<�ia<�$a<�`<��`<]`<�/`<�`<N`<@`<�9`<�k`<D�`<��`<�8a<x}a<øa<��a<�b<�b<�b<�b<��a<H�a<��a<M�a<�ya<ia<�_a<�^a<�ea</ua<U�a<_�a<�a< �a<�b<�b<�"b<�b<�b<
�a<��a<Woa<w)a<;�`<ơ`<Ek`<(D`<�/`<{/`<�C`<k`<�`<��`<�,a<�ta<��a<��a<�b<10b<�8b<�1b<�b<hb<��a<(�a<��a<��a<��a<,a<�a<�a<˙a<��a<��a<��a<�
b<$b<�4b<9b<�-b<5b<V�a<�a<�ia<E"a<!�`<М`<j`<�G`<79`<?`<Y`<�`<��`<�a<mKa<v�a<��a<)b<4%b<�7b<F:b<r.b<|b<��a<��a<X�a<]�a<��a<σa<#a<��a<b�a<d�a<��a<I�a<d�a<tb<5+b<48b<A7b<`&b<b<�a<ɖa<8Qa<7	a<W�`<g�`<�Z`<B>`<6`<hB`<jb`<]�`<n�`<a<�^a<r�a<��a<r
b<�'b<�4b<2b<d"b<�	b<��a<w�a<d�a<`�a<��a<�{a<�ya<#�a<e�a<��a<j�a<��a<��a<�b<R*b<�2b<A,b<�b<9�a<$�a<�va<-/a<�`<��`<7k`<%B`<�+`<�)`< <`<Ea`<c�`<�`<a<oca<�a<��a<Lb<Cb<b<�b<�b<��a<L�a<��a<�a<>ta<?da<$\a<^\a<�da<�ta<��a<��a<E�a<�a<��a<,b<�b<b<��a<��a<��a<�>a<��`<-�`<Wp`<=`<�`<W`<�`<t*`<V`<B�`<�`<�a<\aa<g�a<��a<\�a<�b<�b<��a<��a<��a<v�a<+�a< ra<A^a<�Qa<Ma<�Pa<�\a<�oa<~�a<��a<�a<�  �  ��a<w�a<ab<b<{b<h�a<��a<}�a<}Qa<�a<K�`<��`<]|`<yd`<�]`<0i`<^�`<��`<��`<z$a<�ca<J�a<L�a<J�a<�b<pb<%
b<g�a<l�a<Ҩa<�a<�Ya<�9a<H"a<=a<ka<7a<�1a<�Oa<ua<�a<=�a<��a<db<� b<�#b<}b<��a<��a<�a<oYa<�a<[�`<+�`<i�`<ˀ`<ˀ`<��`<��`<��`<Ka<�]a<q�a<��a<Ib<T&b<97b<�7b<H(b<hb<��a<ݾa<�a<�pa<�Ra<9>a<�3a</5a<�Aa<yXa<Jxa<��a<��a<l�a<�b<v-b<�9b<�6b<�"b<�a<��a<��a<BUa<�a<	�`<�`<��`<��`<�`<\�`<��`<F�`<q:a<\ya<+�a<��a<Ab<^1b<<b<p6b<2"b<�b<��a<�a<ωa<�fa<mKa<4:a<�3a<�8a<�Ha<�ba<��a<��a<0�a<k�a<�b<q3b<�:b<�1b<=b<h�a<��a<!~a<?a<a<�`<>�`<׎`<��`<k�`<��`<t�`<4a<�Ja<��a<S�a<��a<�b<v1b<�6b<�+b<&b<��a<>�a<��a<�wa<�Va<�>a<1a<v.a<]7a<�Ja<�ga<�a<��a<��a<b< b<�0b<b2b<`#b<b<#�a<��a<"_a<�a<<�`<�`<e�`<�|`<�z`<��`<�`<��`<�a<Na<0�a<��a<��a<�b<Pb< b<wb<C�a<`�a<Q�a<Uva<bPa<M1a<�a<�a<�a<qa<�3a<�Ra<�xa<��a<��a<��a<�b<�b<�b<o�a<6�a<��a<�ha<�)a<��`<��`< �`<j`<�\`<�a`<�w`<��`<��`<�
a<~Ia<�a<��a<��a<� b<b<)b<��a<��a<˩a<�a<�Wa<�4a<@a<a<�a<�a<a<t1a<�Sa<�{a<�a<�  �  |�a<t�a<r�a<�
b<�
b<��a<h�a<U�a<�}a<8Ia<�a<��`<%�`<��`<�`<��`<��`<��`<(%a<�Xa<}�a<��a<��a<�b<b<Sb<E�a<0�a<�a<a<IKa<a<�`<��`<�`<\�`<��`<��`<�a<�;a<Wpa<a�a<F�a<��a<�b<�%b<X b<,b<E�a<=�a<�a<�Ua<�&a<��`<��`<��`<��`<��`<� a<)a</Ya<'�a<��a<p�a<�b<1b<�9b<h1b<db<��a<�a<z�a<�]a<2/a<�a<?�`<�`<��`<��`<a<�8a<�ha<��a<��a<��a<� b<�5b<$;b<O/b<gb<��a<b�a<G�a<	Ua<�'a<�a<��`<��`<F�`<��`<ma<�@a<ra<��a<�a<vb<�&b<k9b<�;b<e-b<0b<��a<h�a<�a<dNa<�!a<��`<��`<Y�`<�`<��`<a<yHa<rza<Ůa<W�a<�
b<})b<�9b<�8b<�'b<�b<f�a<3�a<ua<wCa<-a<�`<��`<��`<��`<q�`<�a<xLa<-a<W�a<�a<b<^)b<�6b<{3b<�b<��a<2�a<~�a<ja< 9a<ka<��`<��`<`�`<��`<��`<%a<�Ra<�a<۹a<a�a<(b<�)b<4b<6-b<Pb<��a<��a<��a<yYa<�(a<��`<��`<��`<��`<��`<�`<Ya<�Ka<�~a<~�a<r�a<�b<�b<�!b<b<��a<��a<��a<�ra<@>a<�a<5�`<��`<�`<�`<��`<E�`<[a<�Ba<�va<5�a<A�a<��a<�b<`b<b<��a<)�a<h�a<�\a<�(a<��`<��`<�`<�`<�`<�`<\�`<Ta<bBa<�va<��a<�a<��a<�b<�
b<'�a<��a<�a<��a<Oa<Za<��`<��`<ٶ`<h�`<O�`<�`<��`<a<�Ia<�~a<�  �  0�a<��a<��a<.b<Kb<#b<��a<��a<}�a< |a<�Ta<�2a<�a<K
a<a<�a<�a<
<a<�_a<��a<�a<J�a<�a<Lb<�b<�b<��a<5�a<��a<IQa<+a<"�`<ǧ`<?�`<�n`<Dk`<z`<S�`<�`<P�`<�=a<\}a<&�a<��a<�b<�!b<�$b<�b<(�a<B�a<~�a<�a<�fa<rHa<(3a<#(a<�(a<d4a<�Ja<Dja<��a<�a<��a<h
b<�&b<�6b<�6b<-&b<�b<��a<�a<;`a<S"a<-�`<�`<�`< �`<��`<}�`<��`<��`<�/a<na<a�a<��a<�b<�,b<�9b<�6b<�$b<�b<��a<��a<׎a<�ja<Na<S;a<3a<j6a<�Da<�]a<�~a<
�a<��a<��a<b<�1b<<b<�5b<mb<E�a<N�a<
�a<ILa<�a<'�`<)�`<A�`<�`<�`<�`<i�`<�a<�Da<C�a<�a<��a<�b<�2b<�:b<�1b<mb<
�a<4�a<S�a<y�a<_^a<�Da<�4a<0a<�6a<�Ha<!da<Z�a<��a<�a<u�a<�b<�1b<�6b<�*b<b< �a<��a<�pa<�1a<4�`<#�`<ݟ`<c�`<B�`<%�`<q�`<�`<Ba<�Sa<Αa<9�a<O�a<�b<0b<�1b<�#b<�b<��a<*�a<ҏa<�ha<_Ha<"1a<)$a<�"a<�,a<�@a<�^a<�a<w�a<��a<m�a<<b<U b<�b<�b<��a<��a<ŀa<�Aa<�a<��`<��`<�y`<i`<_j`<B}`<2�`<c�`<�	a<�Ga<��a<@�a<%�a<Db<!b<�b<��a<Y�a<ֵa<�a<�ba<->a<� a<�a<a<�a<a<h.a<YOa<`va<ןa<��a<��a<Pb<;b<�b<9�a<��a<��a<LYa<ia<��`<!�`<#~`<Hc`<?Y`<fa`<�z`<0�`<��`<�a<Sa<�  �  �ka<��a<��a<D�a<B	b<T	b<��a<~�a<3�a<"�a<��a<�qa<a_a<`Ta<~Qa<�Va<qda<ya<�a<Ųa<��a<��a<�b<�b<�b<4�a<��a<��a<gha<�"a<��`<��`<�_`<�5`<�`<�`<�*`<�N`<H�`<'�`<�a<Ta<��a<��a<��a<#b<�$b<n b<b</�a<��a<��a<(�a<-�a<�za<sa<�sa<u|a<�a<h�a<P�a<F�a<� b<_b<�/b<!7b<2/b<b<G�a<I�a<�ua<�.a<(�`<>�`<r`<�L`<�:`<�<`<sS`<p|`<��`<X�`<�>a<1�a<��a<}�a<%b<G4b<Y9b<�/b<b<E�a<A�a<��a<��a<-�a<W�a<z~a<��a<f�a<��a<��a<T�a<��a<�b<�(b<�7b<�9b<�+b<�b<;�a<��a<�_a<�a<R�`<��`<Od`<E`<�9`<�B`<�_`<�`<]�`<.a<�Va<��a<�a<�b<�'b<~7b<07b<.)b<�b<��a<��a<��a<l�a<t�a<�~a<�{a<d�a<E�a<E�a<Z�a<��a<��a<�b<D*b<T5b<�1b<qb<{�a<Y�a<��a<JBa<��`<�`<U}`<ZR`<r9`<�4`<�D`<�g`<R�`<�`<=!a<wha<˪a<�a<�b<�'b<_1b<�+b<\b<��a<`�a<U�a<�a<�a<�xa<!oa<�ma<�ta<L�a<��a<��a<��a<��a<h	b<b<� b<Zb<��a<��a<9�a<Xa<Ka<��`<��`<�P`<�*`<�`<;`<=/`<�W`<E�`<��`<La<e^a<��a<��a<��a<ob<�b<�b<��a<-�a<��a<��a<Dza<�da<�Va<^Pa<bRa<�\a<^na<��a<��a<��a<m�a<��a<fb<	b<��a<k�a<߭a<lra<�-a<	�`<j�`<�b`<[2`</`<�`<`<>.`<�\`<��`<��`<�&a<�  �  �Ja<n�a<4�a<Y�a<�b<�	b<]b<{�a<S�a<��a<�a<ݥa<r�a<o�a<��a<\�a<U�a<��a<y�a<)�a<��a<��a<�b<{b<�b<��a<��a<��a<WEa<6�`<��`<�_`<� `<��_<��_<X�_<��_<�`<3G`<��`<g�`<�-a<�xa<w�a<�a<ib<R b<�#b<mb<*b<��a<)�a<U�a<^�a<i�a<ݱa<��a<��a<�a<q�a<��a<��a<�b<�(b<�3b<�3b<'%b<Qb<��a<�a<;Pa<pa<d�`<�k`<�0`<�`<0�_<��_<�`<}<`<�z`<B�`<a<Qaa<l�a<��a<�b<�+b<v7b<�5b<W)b<Wb<� b<e�a<��a<��a<u�a<��a<D�a<�a<H�a<T�a<��a<�b<�"b<o2b<r9b<4b<�b<��a<��a<P�a<�7a<��`<6�`<(W`<!`<��_<��_<�_<]`<�O`<��`<��`<�-a<Gza<ͽa<1�a<�b<�0b<�7b<�1b<�"b<b<�a<�a<s�a<��a<�a<Ժa<�a<:�a<��a< �a<��a<�b<$b<21b<=4b<�)b<
b<S�a<��a<{ea<�a<o�`<�}`<�=`<+`<q�_<I�_<��_<&`<6_`<��`<�`<Ba<ʋa<
�a<*�a<�b<!-b<�.b<�$b<�b<��a<��a<.�a<H�a<b�a<�a<��a<��a<6�a<��a<[�a<3�a<�b<�b<Db<cb<Sb<�a<,�a<	}a<�2a<�`<�`<aK`<�`<U�_<H�_<�_<��_<�`<XU`<q�`<��`<�:a<�a<��a<��a<�b<b<�b<��a<3�a<��a<#�a<�a<=�a<��a<��a<��a<3�a<�a<ݳa<'�a<��a<e�a<b<�b<Ob<��a<��a<e�a<�Qa<�a<:�`<\i`<C%`<��_<��_<+�_<y�_<��_<�`<�a`<�`<��`<�  �  �.a<xa<��a<��a<��a<qb<�b<� b<��a<�a<��a<��a<G�a<�a<A�a<��a<%�a<B�a<��a<�a<b�a<Lb<�b<�b<��a<4�a<F�a<>sa<f(a<�`<��`<Z2`<��_<��_<%�_<d�_<M�_<B�_<�`< d`<��`<pa<�^a<ۤa</�a<�b<b<=$b<"b<�b<�b<�a<9�a<�a<u�a<�a<��a<��a<C�a<�a<�b<b<J$b<0b<5b</b<b<��a<��a<�a<�1a<l�`<t�`<�<`<��_<�_<I�_<�_<��_<�	`<�L`<��`<V�`<�Ca<P�a<��a<�b<�"b<!4b<F8b<+2b<`&b<�b<�	b<��a<��a<o�a<:�a<0�a<e�a<��a<�b<3b<� b<�.b<�7b<�8b<�-b<�b<��a<�a< ha<#a<��`<�o`<�&`<��_<��_<ٹ_<��_<b�_<�`<Ff`<˷`<�a<�^a<r�a<��a<�b<�)b<Q6b<t6b<�-b< b<�b<�b<r�a<s�a<��a<f�a<�a<�a<��a<b<�b<z!b<�-b<z4b<�1b<�!b<b<��a<�a<�Ha<��`<b�`<hP`<�`<��_<�_<Q�_<Q�_<M�_<�/`<�z`<d�`<�"a<�qa<i�a<8�a<6b<�'b<P/b<f+b<< b<Yb<�b<�a<��a<m�a<�a<��a<�a<x�a<c�a<�a<�b<b<b<f b<�b<Kb<��a<�a<�ca<Ia<�`<�i`<S`<0�_<�_<e�_<r�_<��_</�_<]'`<�u`<�`<�a< ia<��a<w�a<��a<�
b<?b<�b<2�a<�a<d�a<��a<��a<��a<�a<��a<{�a<��a<D�a<x�a<�a<X�a<[b<b<��a<��a<t�a<�~a<�6a<��`<<�`<�=`<��_<�_<ڕ_<)�_<E�_<�_<��_<�5`<X�`<��`<�  �  ta<ia<��a<`�a<+�a<`b<�
b<�b<��a<��a<��a<��a<C�a<��a<��a<��a<��a<,�a<x�a<��a<Mb<�b<�b<�
b<��a<��a<ߤa<vca<Ua<}�`<�g`<d`<��_<��_<�{_<�v_<��_<^�_<E�_<�H`<��`<��`<�Ma<�a<��a</�a<�b<X#b<O%b<� b<b<b<eb<b<�a<>�a<,�a<�b<�b<�b<b<"b<�,b<�3b<�4b<�*b<�b<��a<:�a<�na<Ea<��`<�n`<�`<��_<~�_<ė_<��_<Ķ_<��_<Y/`<q�`<m�`<W0a<.�a<��a<A�a<Pb<�0b<�8b<�6b<�/b<�%b<9b<Lb<�b<�b<�
b<b<�b<b<b<4"b<],b<a5b<�9b<�6b<d(b<�b<;�a<9�a<,Va<�a<3�`<�S`<�`<��_<��_<:�_<��_<��_<��_<J`<��`<�`<+La<`�a<��a<�b<h$b<A4b<#8b<&4b<h+b<!b<�b<Ab<ub<�b<�b<�b<�b<zb<b<s!b<k+b<�2b<;5b<�.b<�b<D�a<s�a<R�a<}5a<��`<��`<r3`<
�_<��_<��_<��_<��_<e�_<@`<�_`<]�`<"a<�`a<n�a<��a<�
b<o#b<j.b<�.b<(b<�b<�b<=	b<�b<�a<C�a<>�a<��a<��a<�b<�	b<�b<wb<� b<�b<�b<�a<c�a<��a<�Ra< a<]�`<!O`<N�_<��_<Z�_<�t_<w_<��_<�_<
`<�[`<�`<�	a<�Xa<��a<��a<f�a<db<�b<Wb<�b<�a<��a<s�a<��a<��a<l�a<��a<��a<��a<��a<w�a<g�a<6b<	b<eb<��a<��a< �a<�oa<�$a<�`<�w`<�!`<��_<��_<�r_<�d_<p_<~�_<��_<A`<Gn`<��`<�  �  Ma<�ca<��a<#�a<�a<�b<_b<	b<�b<��a<d�a<��a<|�a<��a<��a<��a<��a<��a<��a<,�a<b<nb<"b<�	b<�a<}�a<B�a<�]a<�a<��`<�^`<G`<��_<:�_<�o_<�j_<�_<�_<��_<�?`<f�`<��`<�Ga<��a<��a<N�a<�b<9#b<�&b<�"b<�b<�b<�b<�
b<�b<Ob<I	b<bb<ab<b<b<�%b</b<25b<�4b<u)b<b<��a<.�a<ia<�a<��`<Ee`<I`<x�_<~�_<��_<g�_<�_<��_< %`<ax`<w�`<�)a<�za<�a<��a<�b<�/b<�8b<�8b<|2b<:*b<�"b<�b<�b<\b<�b<b<�b<eb< b<�'b<�/b<�7b<�:b<�6b<k&b<b<�a<ۛa< Pa<`�`<��`<�I`<��_<�_<~�_<�_<{�_<�_<��_<#@`<�`<��`<Fa<�a<��a<�b<C"b<�3b<�8b<56b<�.b<&&b<ub<ab<�b<jb<�b<Nb<�b<Ob<�b<&b<<.b<�4b<�5b<�-b<.b<��a<��a<�~a</a<(�`<�}`<U)`<��_<ʪ_<f�_<��_<��_<��_<�`<ZV`<
�`<6a<�Za<D�a<��a<�b<�!b<K.b<�/b<s*b<�!b<�b<{b<�
b<�b<Tb<[b<�b<�b<Y	b<xb<�b<�b<B"b<�b<6b<I�a<��a<~�a<Ma<E�`<)�`<�E`<��_<&�_<\�_<�h_<�j_<��_<ҹ_<��_<�R`<'�`<a<7Sa<9�a<Z�a<��a<?b<�b<b<Fb<s�a<9�a<�a<��a<��a<��a<g�a<��a<(�a<��a<��a<��a<bb<g
b<�b<��a<��a<��a<�ja<�a<��`<�n`<`<��_<�_<�f_<sX_<�c_<ֈ_<��_<d`<�e`<��`<�  �  ta<ia<��a<`�a<+�a<`b<�
b<�b<��a<��a<��a<��a<C�a<��a<��a<��a<��a<,�a<x�a<��a<Mb<�b<�b<�
b<��a<��a<ߤa<vca<Ua<}�`<�g`<d`<��_<��_<�{_<�v_<��_<^�_<E�_<�H`<��`<��`<�Ma<�a<��a</�a<�b<X#b<O%b<� b<b<b<eb<b<�a<>�a<,�a<�b<�b<�b<b<"b<�,b<�3b<�4b<�*b<�b<��a<:�a<�na<Ea<��`<�n`<�`<��_<~�_<ė_<��_<Ķ_<��_<Y/`<q�`<m�`<W0a<.�a<��a<A�a<Pb<�0b<�8b<�6b<�/b<�%b<9b<Lb<�b<�b<�
b<b<�b<b<b<4"b<],b<a5b<�9b<�6b<d(b<�b<;�a<9�a<,Va<�a<3�`<�S`<�`<��_<��_<:�_<��_<��_<��_<J`<��`<�`<+La<`�a<��a<�b<h$b<A4b<#8b<&4b<h+b<!b<�b<Ab<ub<�b<�b<�b<�b<zb<b<s!b<k+b<�2b<;5b<�.b<�b<D�a<s�a<R�a<}5a<��`<��`<r3`<
�_<��_<��_<��_<��_<e�_<@`<�_`<]�`<"a<�`a<n�a<��a<�
b<o#b<j.b<�.b<(b<�b<�b<=	b<�b<�a<C�a<>�a<��a<��a<�b<�	b<�b<wb<� b<�b<�b<�a<c�a<��a<�Ra< a<]�`<!O`<N�_<��_<Z�_<�t_<w_<��_<�_<
`<�[`<�`<�	a<�Xa<��a<��a<f�a<db<�b<Wb<�b<�a<��a<s�a<��a<��a<l�a<��a<��a<��a<��a<w�a<g�a<6b<	b<eb<��a<��a< �a<�oa<�$a<�`<�w`<�!`<��_<��_<�r_<�d_<p_<~�_<��_<A`<Gn`<��`<�  �  �.a<xa<��a<��a<��a<qb<�b<� b<��a<�a<��a<��a<G�a<�a<A�a<��a<%�a<B�a<��a<�a<b�a<Lb<�b<�b<��a<4�a<F�a<>sa<f(a<�`<��`<Z2`<��_<��_<%�_<d�_<M�_<B�_<�`< d`<��`<pa<�^a<ۤa</�a<�b<b<=$b<"b<�b<�b<�a<9�a<�a<u�a<�a<��a<��a<C�a<�a<�b<b<J$b<0b<5b</b<b<��a<��a<�a<�1a<l�`<t�`<�<`<��_<�_<I�_<�_<��_<�	`<�L`<��`<V�`<�Ca<P�a<��a<�b<�"b<!4b<F8b<+2b<`&b<�b<�	b<��a<��a<o�a<:�a<0�a<e�a<��a<�b<3b<� b<�.b<�7b<�8b<�-b<�b<��a<�a< ha<#a<��`<�o`<�&`<��_<��_<ٹ_<��_<b�_<�`<Ff`<˷`<�a<�^a<r�a<��a<�b<�)b<Q6b<t6b<�-b< b<�b<�b<r�a<s�a<��a<f�a<�a<�a<��a<b<�b<z!b<�-b<z4b<�1b<�!b<b<��a<�a<�Ha<��`<b�`<hP`<�`<��_<�_<Q�_<Q�_<M�_<�/`<�z`<d�`<�"a<�qa<i�a<8�a<6b<�'b<P/b<f+b<< b<Yb<�b<�a<��a<m�a<�a<��a<�a<x�a<c�a<�a<�b<b<b<f b<�b<Kb<��a<�a<�ca<Ia<�`<�i`<S`<0�_<�_<e�_<r�_<��_</�_<]'`<�u`<�`<�a< ia<��a<w�a<��a<�
b<?b<�b<2�a<�a<d�a<��a<��a<��a<�a<��a<{�a<��a<D�a<x�a<�a<X�a<[b<b<��a<��a<t�a<�~a<�6a<��`<<�`<�=`<��_<�_<ڕ_<)�_<E�_<�_<��_<�5`<X�`<��`<�  �  �Ja<n�a<4�a<Y�a<�b<�	b<]b<{�a<S�a<��a<�a<ݥa<r�a<o�a<��a<\�a<U�a<��a<y�a<)�a<��a<��a<�b<{b<�b<��a<��a<��a<WEa<6�`<��`<�_`<� `<��_<��_<X�_<��_<�`<3G`<��`<g�`<�-a<�xa<w�a<�a<ib<R b<�#b<mb<*b<��a<)�a<U�a<^�a<i�a<ݱa<��a<��a<�a<q�a<��a<��a<�b<�(b<�3b<�3b<'%b<Qb<��a<�a<;Pa<pa<d�`<�k`<�0`<�`<0�_<��_<�`<}<`<�z`<B�`<a<Qaa<l�a<��a<�b<�+b<v7b<�5b<W)b<Wb<� b<e�a<��a<��a<u�a<��a<D�a<�a<H�a<T�a<��a<�b<�"b<o2b<r9b<4b<�b<��a<��a<P�a<�7a<��`<6�`<(W`<!`<��_<��_<�_<]`<�O`<��`<��`<�-a<Gza<ͽa<1�a<�b<�0b<�7b<�1b<�"b<b<�a<�a<s�a<��a<�a<Ժa<�a<:�a<��a< �a<��a<�b<$b<21b<=4b<�)b<
b<S�a<��a<{ea<�a<o�`<�}`<�=`<+`<q�_<I�_<��_<&`<6_`<��`<�`<Ba<ʋa<
�a<*�a<�b<!-b<�.b<�$b<�b<��a<��a<.�a<H�a<b�a<�a<��a<��a<6�a<��a<[�a<3�a<�b<�b<Db<cb<Sb<�a<,�a<	}a<�2a<�`<�`<aK`<�`<U�_<H�_<�_<��_<�`<XU`<q�`<��`<�:a<�a<��a<��a<�b<b<�b<��a<3�a<��a<#�a<�a<=�a<��a<��a<��a<3�a<�a<ݳa<'�a<��a<e�a<b<�b<Ob<��a<��a<e�a<�Qa<�a<:�`<\i`<C%`<��_<��_<+�_<y�_<��_<�`<�a`<�`<��`<�  �  �ka<��a<��a<D�a<B	b<T	b<��a<~�a<3�a<"�a<��a<�qa<a_a<`Ta<~Qa<�Va<qda<ya<�a<Ųa<��a<��a<�b<�b<�b<4�a<��a<��a<gha<�"a<��`<��`<�_`<�5`<�`<�`<�*`<�N`<H�`<'�`<�a<Ta<��a<��a<��a<#b<�$b<n b<b</�a<��a<��a<(�a<-�a<�za<sa<�sa<u|a<�a<h�a<P�a<F�a<� b<_b<�/b<!7b<2/b<b<G�a<I�a<�ua<�.a<(�`<>�`<r`<�L`<�:`<�<`<sS`<p|`<��`<X�`<�>a<1�a<��a<}�a<%b<G4b<Y9b<�/b<b<E�a<A�a<��a<��a<-�a<W�a<z~a<��a<f�a<��a<��a<T�a<��a<�b<�(b<�7b<�9b<�+b<�b<;�a<��a<�_a<�a<R�`<��`<Od`<E`<�9`<�B`<�_`<�`<]�`<.a<�Va<��a<�a<�b<�'b<~7b<07b<.)b<�b<��a<��a<��a<l�a<t�a<�~a<�{a<d�a<E�a<E�a<Z�a<��a<��a<�b<D*b<T5b<�1b<qb<{�a<Y�a<��a<JBa<��`<�`<U}`<ZR`<r9`<�4`<�D`<�g`<R�`<�`<=!a<wha<˪a<�a<�b<�'b<_1b<�+b<\b<��a<`�a<U�a<�a<�a<�xa<!oa<�ma<�ta<L�a<��a<��a<��a<��a<h	b<b<� b<Zb<��a<��a<9�a<Xa<Ka<��`<��`<�P`<�*`<�`<;`<=/`<�W`<E�`<��`<La<e^a<��a<��a<��a<ob<�b<�b<��a<-�a<��a<��a<Dza<�da<�Va<^Pa<bRa<�\a<^na<��a<��a<��a<m�a<��a<fb<	b<��a<k�a<߭a<lra<�-a<	�`<j�`<�b`<[2`</`<�`<`<>.`<�\`<��`<��`<�&a<�  �  0�a<��a<��a<.b<Kb<#b<��a<��a<}�a< |a<�Ta<�2a<�a<K
a<a<�a<�a<
<a<�_a<��a<�a<J�a<�a<Lb<�b<�b<��a<5�a<��a<IQa<+a<"�`<ǧ`<?�`<�n`<Dk`<z`<S�`<�`<P�`<�=a<\}a<&�a<��a<�b<�!b<�$b<�b<(�a<B�a<~�a<�a<�fa<rHa<(3a<#(a<�(a<d4a<�Ja<Dja<��a<�a<��a<h
b<�&b<�6b<�6b<-&b<�b<��a<�a<;`a<S"a<-�`<�`<�`< �`<��`<}�`<��`<��`<�/a<na<a�a<��a<�b<�,b<�9b<�6b<�$b<�b<��a<��a<׎a<�ja<Na<S;a<3a<j6a<�Da<�]a<�~a<
�a<��a<��a<b<�1b<<b<�5b<mb<E�a<N�a<
�a<ILa<�a<'�`<)�`<A�`<�`<�`<�`<i�`<�a<�Da<C�a<�a<��a<�b<�2b<�:b<�1b<mb<
�a<4�a<S�a<y�a<_^a<�Da<�4a<0a<�6a<�Ha<!da<Z�a<��a<�a<u�a<�b<�1b<�6b<�*b<b< �a<��a<�pa<�1a<4�`<#�`<ݟ`<c�`<B�`<%�`<q�`<�`<Ba<�Sa<Αa<9�a<O�a<�b<0b<�1b<�#b<�b<��a<*�a<ҏa<�ha<_Ha<"1a<)$a<�"a<�,a<�@a<�^a<�a<w�a<��a<m�a<<b<U b<�b<�b<��a<��a<ŀa<�Aa<�a<��`<��`<�y`<i`<_j`<B}`<2�`<c�`<�	a<�Ga<��a<@�a<%�a<Db<!b<�b<��a<Y�a<ֵa<�a<�ba<->a<� a<�a<a<�a<a<h.a<YOa<`va<ןa<��a<��a<Pb<;b<�b<9�a<��a<��a<LYa<ia<��`<!�`<#~`<Hc`<?Y`<fa`<�z`<0�`<��`<�a<Sa<�  �  |�a<t�a<r�a<�
b<�
b<��a<h�a<U�a<�}a<8Ia<�a<��`<%�`<��`<�`<��`<��`<��`<(%a<�Xa<}�a<��a<��a<�b<b<Sb<E�a<0�a<�a<a<IKa<a<�`<��`<�`<\�`<��`<��`<�a<�;a<Wpa<a�a<F�a<��a<�b<�%b<X b<,b<E�a<=�a<�a<�Ua<�&a<��`<��`<��`<��`<��`<� a<)a</Ya<'�a<��a<p�a<�b<1b<�9b<h1b<db<��a<�a<z�a<�]a<2/a<�a<?�`<�`<��`<��`<a<�8a<�ha<��a<��a<��a<� b<�5b<$;b<O/b<gb<��a<b�a<G�a<	Ua<�'a<�a<��`<��`<F�`<��`<ma<�@a<ra<��a<�a<vb<�&b<k9b<�;b<e-b<0b<��a<h�a<�a<dNa<�!a<��`<��`<Y�`<�`<��`<a<yHa<rza<Ůa<W�a<�
b<})b<�9b<�8b<�'b<�b<f�a<3�a<ua<wCa<-a<�`<��`<��`<��`<q�`<�a<xLa<-a<W�a<�a<b<^)b<�6b<{3b<�b<��a<2�a<~�a<ja< 9a<ka<��`<��`<`�`<��`<��`<%a<�Ra<�a<۹a<a�a<(b<�)b<4b<6-b<Pb<��a<��a<��a<yYa<�(a<��`<��`<��`<��`<��`<�`<Ya<�Ka<�~a<~�a<r�a<�b<�b<�!b<b<��a<��a<��a<�ra<@>a<�a<5�`<��`<�`<�`<��`<E�`<[a<�Ba<�va<5�a<A�a<��a<�b<`b<b<��a<)�a<h�a<�\a<�(a<��`<��`<�`<�`<�`<�`<\�`<Ta<bBa<�va<��a<�a<��a<�b<�
b<'�a<��a<�a<��a<Oa<Za<��`<��`<ٶ`<h�`<O�`<�`<��`<a<�Ia<�~a<�  �  ��a<w�a<ab<b<{b<h�a<��a<}�a<}Qa<�a<K�`<��`<]|`<yd`<�]`<0i`<^�`<��`<��`<z$a<�ca<J�a<L�a<J�a<�b<pb<%
b<g�a<l�a<Ҩa<�a<�Ya<�9a<H"a<=a<ka<7a<�1a<�Oa<ua<�a<=�a<��a<db<� b<�#b<}b<��a<��a<�a<oYa<�a<[�`<+�`<i�`<ˀ`<ˀ`<��`<��`<��`<Ka<�]a<q�a<��a<Ib<T&b<97b<�7b<H(b<hb<��a<ݾa<�a<�pa<�Ra<9>a<�3a</5a<�Aa<yXa<Jxa<��a<��a<l�a<�b<v-b<�9b<�6b<�"b<�a<��a<��a<BUa<�a<	�`<�`<��`<��`<�`<\�`<��`<F�`<q:a<\ya<+�a<��a<Ab<^1b<<b<p6b<2"b<�b<��a<�a<ωa<�fa<mKa<4:a<�3a<�8a<�Ha<�ba<��a<��a<0�a<k�a<�b<q3b<�:b<�1b<=b<h�a<��a<!~a<?a<a<�`<>�`<׎`<��`<k�`<��`<t�`<4a<�Ja<��a<S�a<��a<�b<v1b<�6b<�+b<&b<��a<>�a<��a<�wa<�Va<�>a<1a<v.a<]7a<�Ja<�ga<�a<��a<��a<b< b<�0b<b2b<`#b<b<#�a<��a<"_a<�a<<�`<�`<e�`<�|`<�z`<��`<�`<��`<�a<Na<0�a<��a<��a<�b<Pb< b<wb<C�a<`�a<Q�a<Uva<bPa<M1a<�a<�a<�a<qa<�3a<�Ra<�xa<��a<��a<��a<�b<�b<�b<o�a<6�a<��a<�ha<�)a<��`<��`< �`<j`<�\`<�a`<�w`<��`<��`<�
a<~Ia<�a<��a<��a<� b<b<)b<��a<��a<˩a<�a<�Wa<�4a<@a<a<�a<�a<a<t1a<�Sa<�{a<�a<�  �  ��a<��a<	b<�b<$�a<;�a<��a<�ia<�$a<�`<��`<]`<�/`<�`<N`<@`<�9`<�k`<D�`<��`<�8a<x}a<øa<��a<�b<�b<�b<�b<��a<H�a<��a<M�a<�ya<ia<�_a<�^a<�ea</ua<U�a<_�a<�a< �a<�b<�b<�"b<�b<�b<
�a<��a<Woa<w)a<;�`<ơ`<Ek`<(D`<�/`<{/`<�C`<k`<�`<��`<�,a<�ta<��a<��a<�b<10b<�8b<�1b<�b<hb<��a<(�a<��a<��a<��a<,a<�a<�a<˙a<��a<��a<��a<�
b<$b<�4b<9b<�-b<5b<V�a<�a<�ia<E"a<!�`<М`<j`<�G`<79`<?`<Y`<�`<��`<�a<mKa<v�a<��a<)b<4%b<�7b<F:b<r.b<|b<��a<��a<X�a<]�a<��a<σa<#a<��a<b�a<d�a<��a<I�a<d�a<tb<5+b<48b<A7b<`&b<b<�a<ɖa<8Qa<7	a<W�`<g�`<�Z`<B>`<6`<hB`<jb`<]�`<n�`<a<�^a<r�a<��a<r
b<�'b<�4b<2b<d"b<�	b<��a<w�a<d�a<`�a<��a<�{a<�ya<#�a<e�a<��a<j�a<��a<��a<�b<R*b<�2b<A,b<�b<9�a<$�a<�va<-/a<�`<��`<7k`<%B`<�+`<�)`< <`<Ea`<c�`<�`<a<oca<�a<��a<Lb<Cb<b<�b<�b<��a<L�a<��a<�a<>ta<?da<$\a<^\a<�da<�ta<��a<��a<E�a<�a<��a<,b<�b<b<��a<��a<��a<�>a<��`<-�`<Wp`<=`<�`<W`<�`<t*`<V`<B�`<�`<�a<\aa<g�a<��a<\�a<�b<�b<��a<��a<��a<v�a<+�a< ra<A^a<�Qa<Ma<�Pa<�\a<�oa<~�a<��a<�a<�  �  �a<�b<H	b<�b<��a<1�a<�a<�Ga<D�`<�`<v``<�`<9�_<K�_<��_<�_<`�_<i.`<�s`<2�`<Oa<F]a<��a<j�a<(�a<Ub<�b<�b<$�a<��a<��a<�a<�a<��a<G�a<ڝa<Ӣa<%�a<��a<{�a<��a<��a<Ob<5b<O b<�b<�a<��a<��a<Ka<��`<��`<}g`<+`<b�_<\�_< �_<��_<:*`<g`<T�`<��`<�Oa</�a<��a<Yb<�&b<w5b<I6b<�+b<�b<�b<N�a<�a<
�a<��a<4�a<��a<�a<��a<��a<��a<L	b<?b<
/b<�7b<y4b<�"b<c b<��a<��a<Ca<��`<*�`<U``<(`<`<��_<�_<`<F`<��`<��`<4!a<�na<b�a<`�a<-b<-0b<�9b<�5b<(b<]b<�a<x�a<P�a<��a<v�a<w�a<��a<7�a<�a<��a<K�a<b<�$b<s3b<a8b<g0b<b<�a<s�a<�ta<�'a<(�`<-�`<�I`<�`<��_<b�_<,�_<�`<5V`<��`<��`<�6a<2�a<��a<��a<�b<b/b<�3b<f,b<2b<bb<��a<1�a<z�a<��a<3�a<�a<�a<b�a<��a<��a<��a<b<�$b<�/b<�0b<Q#b<�b<��a<,�a<�Ra<8a<��`<ai`<�*`<`�_<c�_<1�_<��_<i `<`[`<��`<E�`<O>a<&�a<��a<��a<�b<b<lb<�b<��a<)�a<��a<y�a<��a<��a<&�a<�a<1�a<Ȫa<_�a<��a<�a<��a<�b<	b<Pb<��a<5�a<0�a<Aca<6a<R�`<Dz`<�3`<�_<��_<��_<��_<��_<`<mW`<<�`<_�`<�>a<�a<ļa<Q�a<�a<?b<=b<O�a<f�a<a�a<=�a<�a<s�a<4�a<Q�a<��a<w�a<��a<z�a<��a<��a<�  �  ��a<'b<xb<_�a<(�a<f�a<kua<�+a<�`<��`<�3`<[�_<�_<�_<��_<&�_<	�_<�_<>H`<��`<5�`<kBa<,�a<��a<��a<!b<$b<Ub<b<��a<v�a<��a<��a<o�a<?�a<T�a<��a<0�a<L�a<U�a<��a<b<�b<f b<�b<�b<��a<v�a<Uya<9-a<t�`<��`<<9`<G�_<T�_<��_<J�_<f�_<�_<S8`<��`<�`<51a<.�a<��a<M�a<�b<+1b<�7b<�3b<�(b<�b<cb<# b<��a<��a<��a<��a<^�a<�a<@b<b<�b<f+b<[5b<�7b<�.b<�b<#�a<��a<@sa<s#a<��`<V{`<s0`<�_<?�_<��_<��_<��_<!`<�Y`<�`<T�`<&Ra<*�a<�a<�	b<A(b</7b<k9b<2b<�%b<�b<�b<V�a<��a<��a<�a<P�a<��a<��a<�b<kb<#b<�/b<�7b<�6b<)b<eb<6�a<Ϣa<�Xa<�a<�`<�_`<�`<��_<4�_<T�_<3�_<s�_<�%`<Mo`<��`<�a<Mga<S�a<�a<Xb<')b<~3b<2b<�(b<�b<9b<��a<T�a<"�a<.�a<p�a<��a<r�a<��a<lb<zb<�!b<�,b<'2b<�,b<,b<��a<��a<a<�4a<.�`<��`<";`<;�_<S�_<��_<\�_<��_<E�_<�,`<y`<��`<�a<#ma<��a<��a<�b<�b<�b<Mb<Nb<�a<��a<{�a<	�a<-�a<��a<-�a<�a</�a<��a<D�a<U�a<�b<)b<0b<�b<	�a<��a<J�a<Ia<��`<P�`<{O`<`<(�_<�_<Ӌ_<r�_<�_<7�_<P*`<�z`<��`<"a<�la<��a<�a<"�a<�b<�b<A b<��a<��a<��a<��a<��a<��a<ٻa<J�a<�a<9�a<��a<��a<��a<�  �  �b<�	b<5b<��a<k�a<��a<-fa<ea<�`<�k`<�`<��_<q�_<�r_<i_</y_<ˡ_<D�_<�,`<��`<��`<�0a<�{a<y�a<��a<*b<�b<�b<�b<!b<��a<h�a<\�a<��a<4�a<��a<��a<�a<��a<� b<Ub<Fb<:b< b<(b<�b<��a<~�a<ia<�a<Y�`<jl`<�`<�_<�_<=�_<ь_<�_<��_<{`<l`<��`<&a<�oa<]�a<7�a<�b<S-b<7b<�7b<i1b<�'b<*b<�b<(b<|b<�
b<b<�b<�b<7b<�b<�)b<3b<J8b<�6b<C*b<�b<P�a<̪a<�aa<�a<g�`<�_`<�`< �_<e�_<�_<P�_<��_<k�_<�<`<s�`<��`<G?a<��a<��a<� b<;"b<�4b<e:b<�7b<�/b<�%b<+b<~b<wb<_b<b<b<�b<Sb<�b<�#b<�-b<�5b<'9b<S4b<]#b<�b<Z�a<��a<[Fa<��`<ԗ`</C`<&�_<$�_<��_<��_<4�_<.�_<�`<�S`<K�`<�a<�Ua<͟a<��a<Eb<,$b<�1b<g4b<�/b<�&b<ub<�b<�b<{b<%b<�b< b<[
b<�b<�b<:!b<�*b<s1b<C2b<c)b<pb<��a<��a<sra<*!a<�`<?p`<�`<��_<�_<E�_<�_<�_<��_<�`<m^`<!�`<�a<u\a<��a<��a<��a<�b<�b<Ob<�b<B	b<x�a<M�a<��a<!�a<��a<G�a<��a<	�a<��a<��a<xb<Gb<b<b<"b<K�a<-�a<"�a<�7a<��`<�`<4`<��_<'�_<{_<@h_<#o_</�_<��_<�`<�``<$�`<1a<8]a<H�a<��a<�a<%b<�b<�b<��a<s�a<��a< �a<�a<	�a<E�a<��a<��a<��a<Z�a<��a<F�a<�  �  4b<�8b<�3b<Zb<��a<��a<�ea<q�`<Չ`<!`<D�_<�4_<��^<#�^<_�^<ս^<H�^<�K_<J�_<�.`<�`<a<3�a<��a<a
b<.b<�?b<�Bb<D>b<h6b<k/b<+b<�)b<�*b<$,b<?-b<F-b<�-b<r/b<4b<�;b< Eb<vMb<#Pb<*Gb<�-b<��a<պa<�`a<J�`<�~`<[`<�_< 7_<�^<��^<��^<��^<I3_<��_<�`<�|`<�`<4ea<C�a<�b<�>b<�[b<)hb<�gb<Mab<Yb<sRb<xNb<�Mb<�Mb<�Nb<,Nb<3Mb<�Lb<;Nb<�Rb<�Yb<Hbb<hb<tfb<9Wb<X6b<��a<U�a<�Pa<��`<�f`<��_<U�_<~*_<"�^<:�^<s�^<�_<Y_<ν_<�1`<߫`<�!a<"�a<��a<�"b<Mb<�cb<�jb<?gb<:_b<Wb<$Qb<6Nb<�Mb<JNb<�Nb<5Nb<�Mb<�Mb<�Ob<aUb<B]b<Teb<.ib<�cb<�Nb<�&b<;�a<��a<,a<	�`<�<`<��_<�`_<_<�^<��^<��^<U_<At_<��_<�U`<-�`<kAa<פa<h�a<�-b<�Pb<�ab<7db<�^b<qVb<�Nb<�Ib<'Hb<1Hb<�Hb<PIb<{Hb<Hb<�Hb<2Lb<qRb<�Zb<�ab<�bb<9Xb<+=b<}b<��a<�ja<[�`<Ȅ`<z
`<
�_<17_<��^<��^<��^<��^<)_<��_<��_<�l`<�`<cQa<��a<P�a<�%b<wAb<1Lb<�Jb<�Bb<D9b<�1b<�,b<�*b<H*b<T*b<e)b<�'b<''b< (b<,b<�2b<�:b<B@b<1>b<�.b<&b<��a<�a<&a<~�`<�:`<t�_<JU_<��^<�^<��^<��^<w�^<g)_<Ӎ_<�`<M{`<��`<Za<r�a<6�a<b<[1b<8b<y4b<9,b<�#b<�b<�b<ab<�b<�b<b<�b<b<�b<�#b<�+b<�  �  3b<E9b<�5b<F#b<�a<^�a<�ma<?a<I�`<4`<�_<�C_<��^<��^<n�^<��^<O_<�Z_<��_<:`<�`<�$a<�a<��a<Bb<�1b<qAb<�Bb<]<b<U2b<�(b<G"b<�b< b<�b<�b<c b<"b<�%b<,b<p6b<SBb<�Lb<+Qb<Jb<2b<Pb< �a<�ha<t�`<��`<�`<2�_<�F_<�_<��^<��^<R _<C_<+�_<�`<�`<a�`<gma<��a<8b<@Cb<_b<^ib<]gb<�^b</Tb<Kb<�Db<�Ab<�@b<�@b<�@b<�@b<�Ab<<Eb<Lb<�Ub<7`b<�gb<	hb<�Zb<;b<�b<�a<SYa<��`<r`<��_<�_<y:_<��^<H�^<[�^<_<\h_<��_<$>`<��`<�*a<�a<��a<(b<Qb<fb<+kb<fb<\b<sQb<Ib<�Cb<�Ab<3Ab<\Ab<Ab<JAb<Cb<�Gb<�Ob<�Yb<�cb<�ib<�eb<�Rb<�+b<��a<��a<�4a<�`<�H`<<�_<�o_<I!_<��^<��^<E�^<`/_<(�_<+�_<ia`<+�`<�Ia<��a<��a<v2b<4Tb<Ncb<6db<�\b<^Rb<hHb< Ab<=b<�;b<�;b<�;b<�;b<J<b<�>b<�Db<QMb<�Wb<�`b<�cb<"[b<wAb<�b<��a<�ra<�a<Ϗ`<`<M�_<�F_<� _<��^<��^</�^<�8_<��_<b`<�w`<h�`<�Ya<��a<��a<O*b<�Db<gMb<Jb<7@b<d4b<A*b< #b<6b<yb<�b<�b<Jb<�b<b<]%b<�.b<�8b<@b<�?b<�1b<�b<��a<��a<�.a<9�`<)F`<}�_<	d_<�_<��^<÷^<k�^<��^<�8_<��_<�`<�`<��`<�aa<8�a<h�a<b<�3b<�8b<>3b<)b<Bb<�b<�b<Pb<�b<b<�b<lb<�b<�b<�b<�(b<�  �  .b<>:b<�;b<�-b<Vb<n�a<q�a<F!a<β`<;?`<0�_<4o_<c$_<��^<��^<��^</4_<K�_<��_<�\`<��`<�=a<�a<��a<�b<@;b<]Fb<�Bb<�5b<%b<�b<�b<�a<�a<��a<(�a<��a<��a<�b<�b</&b<�8b<�Ib<�Sb<�Qb<�=b<�b<f�a<;�a<a<ɩ`<Q7`<��_<As_<(2_<�_<_<�/_<�o_<P�_<_4`<��`<pa<�a<c�a<&"b<�Ob<*gb<�lb<eb<Vb<�Db<�4b<�(b<Y b<�b<�b<�b<+b<>!b<5*b<<7b<�Gb<�Xb<gb<plb<�cb<0Hb<wb<��a<�qa<�a<Ǔ`<�!`<5�_<h_<�/_<}_<!_<�K_<$�_<n�_<�a`<��`<FEa<t�a<�a<�6b<�[b<�lb<�lb<�ab<Qb<�?b<�0b<�%b<�b< b<�b<�b<�b<O$b<�.b<�<b<Nb<�^b<�jb<�kb<']b<C:b<� b<��a<�Na<	�`<l`<��_<"�_<�O_<m!_<�_<x(_<J]_<��_<�`<��`<��`<ca<��a<�b<�?b<�]b<?hb<�cb<�Vb< Eb<b4b<�&b<;b<�b<�b<4b<b<=b<�!b<�-b<=b<iNb<�]b<yfb<�bb<JMb<�"b<;�a<3�a<"a<�`<n;`<��_<Qs_<,0_<�_<�_<�'_<�e_<%�_<:&`<w�`<x	a<Pqa<��a<�
b<�6b<�Lb<�Pb<�Gb<�7b<�$b<b<�b<��a<F�a<^�a<��a<��a<u�a<�b<�b<� b<�1b<'?b<(Db<;b<�b<��a<E�a<(Ga<D�`<�g`<c�_<�_<w:_<�_<��^<�^<�_<td_<l�_<V1`<��`<la<Uxa<��a<b<*b<^:b<5:b<�.b<b<zb<h�a<d�a<h�a<��a<b�a<|�a<�a<��a<x�a<;b<�b<�  �  �#b<9b<�Bb<u;b<�b<��a<��a<YHa<��`<�t`<2`<Ͳ_<m_<�B_<7_<�J_<9|_<��_<Y&`<F�`<��`<;ca<��a<� b<�/b<kGb<rKb<�?b<�)b<�b<��a<i�a<��a<��a<��a<2�a<B�a<;�a<	�a<��a<#b<�'b<�Bb<hUb<�Zb<�Mb<D+b<i�a<��a<WCa<��`<zo`<+`<ڸ_<�|_<�\_<6\_<�z_<+�_<T	`<_m`<��`<�Ea<J�a<�a<99b<`b<�pb<ob<_b<QFb<�*b<=b<��a<b�a<��a<��a<�a<'�a<��a<��a< b<0b<�Kb<cb<�pb<5ob<CZb<�.b<��a<Жa<@2a<��`<�\`<��_<��_<n{_<�d_<�m_<��_<w�_<;1`<�`<a<ma<Q�a<�b<�Kb<jjb<tb<^lb<�Xb<�=b<2"b<�b<�a<~�a<��a<��a<��a<��a<��a<Vb<Vb<�9b<�Tb<Sib<{rb<�jb<Nb< b<��a<va<�a<��`<�9`<��_<��_<�m_<�a_<kt_<e�_<��_<N`<J�`<#a<��a<G�a<�$b<�Rb<�ib<Zmb<�`b<7Jb<�.b<`b<?�a<��a<A�a<g�a<8�a<l�a<r�a<8�a<�b<�!b<�=b<�Vb<hb<�kb<(]b<�8b<:�a<��a<cKa<�`<�s`<B`<�_<�z_<�X_<V_<�r_<�_<*�_<<_`<��`<�3a<�a<r�a<�!b<0Gb<�Vb<"Sb<�Ab<�'b<�
b<j�a<�a<��a<2�a<��a<Z�a<ߺa<7�a<Y�a<^�a<�b<$b<%;b<fHb<rFb<1b<b<2�a<�ka<�a<��`<0`<��_<�_<GM_<\6_<�>_<"f_<��_<2`<�g`<��`<A<a<3�a<��a<b<�8b<�Ab<�9b<�%b<b<�a<S�a<��a< �a<F�a<S�a<Ҩa<$�a<;�a<?�a<��a<�b<�  �  9b<�2b<�Fb<dHb<T4b<�	b<��a<�va<�a<�`<�Y`<7`<)�_<�_<��_<�_<��_<	`<�p`<b�`<�2a<��a<��a<	b<�Bb<�Rb<kMb<7b<1b<f�a<s�a<'�a<�a<poa<qda<(ca<_ka<�}a<��a<��a<�a<	b<5b<�Rb<
bb<Q]b<�Bb<�b<��a<�ta<�a<W�`<�[`<�`</�_<�_<q�_<��_<`<�Y`<U�`<>a<xa<t�a<zb<�Qb<{pb<>yb<�mb<�Rb<�-b<b<X�a<��a<��a<A�a<��a<��a<�a<R�a<��a<�a<Lb<�5b<*Yb<�qb<yyb<rlb<*Ib<�b<%�a<&ga<�a<ѥ`<gO`<.
`<~�_<y�_<\�_<��_<�.`<�~`<��`<u=a<��a<��a<�3b<]ab<.xb<@yb<Qgb<-Hb< !b<�a<j�a<	�a<Řa<��a<E�a<c�a<C�a<n�a<��a<��a<ub<�Bb<cb<�vb<�wb<Acb<8b<��a<x�a<Fa<�`<�`<B4`<��_<*�_<�_<��_<� `<�C`<`�`<z�`<Ya<�a<�b<@b<�eb<1ub<[ob<XXb<�5b<tb<��a<��a<O�a<�a<9�a<%a<��a<��a<��a<��a<��a<�#b<"Ib<[eb<sb<�lb<?Pb<�b<��a<�|a<�a<p�`<�]`<`<0�_<�_<Z�_<��_<�`<�M`<5�`</a<*fa<��a<�b<G:b<�Wb<�^b<�Qb<c5b<=b<b�a<��a<��a<}a<�ia<�`a<�`a<�ja<�~a<Úa<l�a<A�a<_b<I1b<:Ib<�Pb<'Cb<Xb<��a<4�a<�;a<��`<'y`<1"`<r�_<F�_<Θ_<I�_<r�_<�_<�N`<K�`<�a<�ka<d�a<Ob<�/b<KFb<Gb<�4b<�b<'�a<�a<=�a<�}a<{ea<[Va<#Qa<pUa<�ca<{a<Úa<.�a<E�a<�  �  �a<f%b<GDb<8Pb<�Eb<E$b<��a<2�a<�Ta<=�`<=�`<Mh`<�2`<�`<�	`<�`<�>`<�x`<^�`<�a<�ka<~�a<xb<�4b<�Qb<,Xb<xHb<�&b<��a<��a<ϊa<?Xa<I.a< a<u�`<��`<	a<�"a<�Ia<cza<��a<��a<Eb<Ib<cb<whb<Wb</b<�a<`�a<�Ua<�a<t�`<\t`<DF`<].`<.`<�E`<~s`<��`<�a<�Wa<��a<��a<�:b<�fb<�|b<a{b<eb<G>b<�b<Y�a<˝a<(ma<Fa<�+a<�a<3 a<�/a<+Ma<�va<̨a<��a<b<�Gb<zkb< ~b<�zb<�`b<�0b<��a<؞a<�Ia<Z�`<�`<�p`<�H`<p7`<Q>`<~\`<'�`<��`<%%a<�za<W�a<~b<�Ob<�sb<�b<�wb<[b<j/b<<�a<C�a<�a<2_a<�;a<�%a<�a<9$a<�8a<4Za<Նa<R�a<�a<�(b<�Ub<tb<�b<�tb<�Rb<�b<��a<݁a<2,a<��`<k�`<�^`<�=`< 4`<�B`<�g`<��`<N�`< =a< �a<!�a<U&b<�Xb<1ub<�zb<qjb<CHb<�b<��a<@�a<wa<uLa<�-a<5a<�a<-$a<
=a<�ba<]�a<p�a<��a<N3b<�[b<�sb<�wb<�db<�:b<�a<d�a<�[a<�a<��`<ht`<ED`<R*`<�'`<p=`<Xi`<Ч`<��`<�Ga<�a< �a<$%b<�Ob<�cb<�`b<%Ib<!b<R�a<��a<}a<pKa<t#a<7a<��`<��`<�
a<o'a<VPa<,�a<�a<��a<�b< Cb<*Ub<lQb<�6b<b<��a<@sa<�a<��`<�~`<�B`<K`<�`<,`<�,`<S``<��`<��`<Ja<u�a<_�a<(b<Bb<<Ob<�Eb<�(b<��a<u�a<O�a<�Ya<,a<�a<��`<��`<]�`<�a<�'a<�Ta<ĉa<��a<�  �  A�a<�b<v9b<Pb<�Ob<;8b<&b<%�a<�a<Ga<Aa<��`<[�`<��`<~`<��`<
�`<��`<Ta<|Za<,�a<��a<Zb<=Fb<�Yb<�Ub<3;b<�b<�a<��a<OFa<7a<5�`<��`<��`<�`<�`<�`<��`<6/a<�ua<s�a< b<�6b<�[b<�kb<Fdb<�Fb<�b<��a<ݓa<FNa<�a<g�`<l�`<M�`<>�`<��`<��`<�a<?Pa<��a<��a<�b<�Sb</ub<�b<;ub<�Sb<� b<@�a<
�a<5Ta<|a<-�`<�`<ȭ`<�`<��`<��`<�!a<�ba</�a<��a<�,b<�\b<[zb<��b<Dqb<)Lb<�b<��a<��a<�Ga<�
a<��`<�`<�`<��`<��`<��`<d,a<�na<׵a<��a<`7b<�db<�~b<�b<'nb<�Eb<b<��a<΂a<�>a<"a<��`<��`<��`<B�`<F�`<��`<�6a<0za<-�a<�b<"?b<8ib<ub<�~b<�fb<J;b<��a<}�a<#ta<�0a<��`<�`<ð`<Ψ`<��`<}�`<�a<^=a<āa<��a<Wb<LCb<kjb<}b<jxb<7]b</b<��a<��a<�ea<$a<[�`<u�`<V�`<ԧ`<��`<��`<�	a<%Ga<f�a<��a<b<*Ib<�lb<{b<�qb<{Rb<� b<��a<�a<YRa<a<q�`<k�`<A�`<'�`<k�`<��`<�a<$Ba<{�a<��a<b<>b<�]b<>hb<�Zb<8b<Mb<��a<gza<3a<��`<��`<��`<��`<F�`<��`<�`<��`<�;a<"�a<0�a<b<�4b<{Qb<&Xb<TGb<�!b<��a<#�a<�`a<a<n�`<�`<��`</}`<�`<^�`<�`<8�`<B>a<,�a<��a<@b<Q3b<'Mb<JPb<<b<�b<��a<;�a<�Oa<�a<�`<��`<��`<�y`<�`<��`<��`<a<�Ha<�a<�  �  �a<�a<&b<�Fb<YPb<�Cb<L$b<��a<��a<�a<�Ta<�(a<a<��`<-�`<��`<�a<4a<�ba<�a<��a<b<�2b<BOb<Xb<Jb<j%b<�a<��a<�Pa<��`<�`<�i`<)8`< `<}`<�*`<U`<��`<��`<j3a<Y�a< �a<�b<�Kb<�eb<�hb<�Ub<.2b<�b<��a<S�a<Rda<a<a<� a<�a<�a<�!a<�=a<�fa<��a<��a<�	b<�<b<db<�zb<|b<Sfb<D:b<��a<��a<OYa<a<ܸ`<bz`<�N`<y9`<<`<2V`<K�`<#�`<�a<�ka<�a<
b<�Eb<�mb<�~b<1yb<F_b<�5b<�b<��a<�a<�da<�?a<�'a<a<e!a<�3a<eSa<�~a<^�a<,�a<� b<�Ob<Qqb<��b<�yb<�[b<P(b<1�a<��a<==a<��`<n�`<�i`<BE`<�7`<yB`<<d`<ƚ`<��`<3a<Q�a<��a<4 b<�Ub<�ub<Eb<1rb<wRb<�$b<7�a<�a<��a<#Ua<�3a<�a<�a<�"a<@9a<�\a<�a<e�a<2�a<�,b<�Wb<�sb<�{b<�lb<yGb<zb<��a<�pa<ma<��`<�`<�U`<�8`<_3`<�E`<o`<��`<n�`<Ja<��a<��a<;.b<�\b<�tb<vb<�ab<<b<�	b<��a<b�a<`fa<i<a<�a<�a<�a<�a<�3a<�Za<܊a<��a<��a<)b<�Nb<|cb<9cb<�Kb<wb<��a<8�a<�9a<[�`<9�`<�W`<f+`<z`<y`<1`<�``<��`<�`<�Da<��a<$�a<�b<�Db<gUb<2Ob<�4b<�
b<�a<��a<ga<?7a<�a<�`<2�`<�`<	a<r#a<sNa<�a<y�a<��a<�b<�?b<Ob<�Gb<�)b<�a<ða<�_a<u
a<׷`<to`<�6`<O`<�`<�`<�1`<�h`<��`<�a<OWa<�  �  <za<��a<�b<�5b<Ib<�Fb<d2b<�b<��a<D�a<��a<�|a<fa<�Xa<�Ua<�[a<�ka<�a<i�a<��a<|�a<b<N>b<Pb<�Nb<;7b< 	b<��a<�qa<�a<ر`<.V`<`<7�_<�_<��_<)�_<4�_<�6`<ˎ`<��`<jRa<ܭa<��a<�4b<�Wb<�db<�\b<aDb<u!b<��a<c�a<��a<'�a<G�a<?xa<�xa<�a<ܖa<i�a<��a<� b<�*b<_Pb<�kb<�wb<Gob<lPb<pb<��a<xa<.a<��`<!^`<w`<��_<��_<��_<s�_<e#`<p`<$�`<_,a<N�a<d�a<|(b<�Yb<Jtb<�xb<�ib<iLb<&b<:�a<��a<n�a<�a<C�a<��a<>�a<��a<��a<��a<>�a<�b<T=b<`_b<�ub<ezb<�ib<�Bb<b<��a<�Xa<�`<�`<�C`<	`<W�_<��_<�_<��_<,;`<��`<��`<1Ma<ƪa<��a<�;b< eb<�wb<[ub<�`b<x?b<_b<f�a<O�a<
�a<�a<a�a<�a<�a<��a<�a<��a<f�a<,b<�Db<gcb<]tb<rb<
Zb<+b<��a<K�a<�2a<I�`<�t`<6&`<��_<��_<~�_<!�_<8	`<�O`<��`<�a<�ga<��a<Db<�Eb<gb<%rb<Jhb<;Nb<j)b<��a<o�a<��a<-�a<Da<1ta<�ra<�za<��a<I�a<��a<��a<�b<�<b<nVb<�`b<�Vb<6b<��a<��a<�Ya<��`<�`<�<`<��_<G�_<ť_<$�_<L�_<��_<�I`<��`<Pa<�da<l�a< b<�0b<�Jb<�Nb<?b</!b<K�a<��a<�a<��a<�la<�[a<�Ta<�Va<�ba<�xa<��a<��a<B�a<fb<@.b<RDb<�Hb<8b<�b<��a<9�a<O&a<[�`<Me`<`<"�_<|�_<�_<��_<o�_<	`<�[`<+�`<>a<�  �  RLa<�a<o�a<}!b<�<b<(Cb<*9b<�#b<�b<z�a<��a<{�a<�a<��a<ƪa<u�a<�a<o�a<��a<7�a<�b<�.b<�Bb<LJb<O@b<,!b<��a<ڞa<�Aa<��`<�m`<8`<O�_<�p_<_K_<;E_<f^_<�_<��_<:F`<��`<"a<�a<��a<b<)Fb<�Zb<X\b<�Nb<�7b<%b<b<��a<S�a<��a<��a<��a<��a<�a<��a<�	b<�%b<iBb<\b<�lb<ob<g^b<�7b<r�a<�a<�Da<��`<$o`<�`<�_<C�_<dg_<�j_<>�_<��_<!`<م`<_�`<N[a<��a<m	b<�Bb<Ceb<rb<�lb<�Zb<�@b<%b<b<��a<+�a<~�a<��a<H�a<��a<��a<|b< b<�5b<Qb<agb<sb<�nb<UVb< 'b<E�a<��a<F"a<J�`<OM`<��_<N�_<�v_<,e_<�r_<]�_<*�_<�A`<��`<~a<�|a<#�a<b<�Pb<}kb<�qb<`gb<�Qb<y6b<�b<�b<��a<�a<�a<��a<��a<��a<{�a<b<�b<e:b<�Tb<�gb<�nb<�cb<Db<�b<I�a<Tba<�`<#�`< '`<i�_<��_< h_<a_<Vy_<	�_<p�_<	^`</�`<j3a<��a<K�a<�+b<WUb<[hb<hb<�Xb<�?b<'#b<b<��a<X�a<��a<��a<��a<��a<��a<��a<��a<�b<�0b<lHb<TWb<�Wb<�Eb<Jb<��a<��a<z&a<i�`<�N`<f�_<��_<	`_<vC_</F_<h_<�_<��_<>_`<P�`<�3a<a<��a<�b<�;b<Hb<EBb<|/b<�b<��a<��a<�a<�a<߭a<��a<۪a<ѱa<��a<-�a<v�a<�b< b<A6b<�Ab<==b<�$b<6�a<'�a<[Va<��`<��`<�`<�_<{s_<�C_<�2_<{@_<m_<.�_<�`<Sx`<��`<�  �  �%a<Q�a<��a<�b<C/b<�<b<�:b<�.b<�b<�b<��a<}�a<j�a<]�a<��a<��a<��a<��a<Mb<b<&&b<?7b<�Bb<cBb<�1b<�b<��a<�}a<[a<��`<�6`<�_<�l_<�&_<��^<��^<�_<�M_<]�_<�`<=`<��`<�^a<M�a<b<|4b<�Ob<�Xb<bSb<�Eb<F5b<�%b<�b< b<�b<zb<mb<�b<�b<. b<�-b<�>b<�Qb<�ab<�ib<�db<jMb< b<v�a<t�a<Za<j�`<�5`<��_<�u_<8_<_<�_<�B_<l�_<�_<N`<��`<[2a<��a<��a<�,b<�Ub<uib<�kb<Ubb<YRb<�@b<k1b<�%b<cb<Wb<�b<ub<�b<�"b<w,b<i:b<hKb<�\b<�ib<�mb<3bb<3Cb<�b<A�a<�ba<��`<�`<e`<<�_<�]_<�*_<�_<�&_<tV_<ڢ_<�`<�t`<�`<Va<c�a<5b<�<b<0^b<qkb<ib<�\b<?Kb<�9b<`+b<� b<tb<�b<�b<b<�b<�!b<�,b<�;b<�Lb<C]b<�gb<�fb<%Ub<�.b<��a<�a<!:a<�`<OV`<��_<Ǌ_<D_<>_<�_<�-_<�g_<G�_<�#`<Ε`<8a<�ra<��a<�b<�Cb<X]b<1db<4]b<�Mb<F;b<�)b<�b<b<�b<kb<Vb<�b<pb<b<�b<�.b<�?b<�Mb<fTb<�Mb<�4b<�b<��a<afa<�`<�`< `<�_<S_<�_<0�^<=�^<�_<�`_<��_<�'`<��`<�
a<�pa<<�a<�b<3,b<R?b<+Ab<�6b<h&b<?b<Kb<>�a<0�a<��a<��a<��a<��a<|�a< �a<�	b<�b<�+b<�8b<M<b<�0b<�b<��a<,�a<i0a<+�`<�O`<��_<|z_<(+_<��^<
�^<5�^<?$_<�p_<Q�_<PC`<>�`<�  �  �a<�qa<��a<��a< %b<#7b<(:b<4b<�)b<�b<�b<�b<�b<�b<ub<�b<�b<rb<Ob<g%b<�0b<:;b<�@b<�;b<P&b<��a<�a<ga<��`<��`<(`<
�_<�@_<��^<��^<��^<�^< _<�y_<T�_<�]`<+�`<SFa<�a<x�a<�'b<Gb<kTb<�Tb<�Mb<�Cb<;b<H5b<�2b<�2b<�3b<�4b<�5b<�7b<)<b<�Cb<Nb<�Yb<}cb<Ffb<�\b<�@b<�b<o�a<|ka<�`<~�`<�`<)�_<hH_<q_<�^<��^<�_<Z_<��_<�)`<ˡ`<a<��a<��a<�b<*Jb<,bb<�ib<�eb<6\b<tQb<�Hb<'Cb<�@b<@b<V@b<F@b<�@b<2Bb<�Fb<Nb<FXb<�bb<�ib<hhb<bXb<z5b<\�a<��a<VIa<��`<�_`<��_<x�_<�/_<>�^<f�^<-�^<(_<�w_<��_<�Q`<��`<I<a<��a<Y�a<�.b<�Sb<�eb<ehb<�ab<ZWb<�Lb<�Db< @b<�=b<�=b<�=b<=b<�=b<�?b<�Db<Mb<�Wb<Gab<�eb<`b<�Ib<�b<�a<�a<\a<ɪ`<�2`<��_<�^_<"_<u�^<{�^<��^<o:_<h�_<�_<`t`<g�`<*Za<C�a<Bb<�6b<Tb<`b<k^b<oUb<�Ib<?b<O7b<�2b<�0b<�/b<�.b<�-b<�-b<0b<�5b<>b<Hb<�Ob<�Pb<cEb<3(b<��a<��a<mNa<��`<h`<�_<��_<&_<A�^<�^<W�^<��^<m4_<��_<[`<�z`<��`<�Ya<�a<��a<� b<8b<�>b<L:b<=0b<�$b<�b<pb<sb<`b<5b<�b<�b<b<&b<�b<�'b<�1b<�8b<7b<�&b<�b<~�a<�za<a<e�`<4-`<�_<�O_< �^<��^<Գ^<��^<��^<�E_<@�_<� `<��`<�  �  a<�ia<&�a<r�a<"!b<�4b<�9b<�5b<b-b<�%b<C b<%b<:b<b< b<�b<�b<� b<9$b<�*b<�3b<X<b<�?b<9b<2"b<��a<�a<_a<��`<�`<�`< �_<^1_<��^<�^<��^<��^<�_<�j_<_�_<bR`<��`<�=a<d�a<��a<�"b<�Cb<�Rb<�Tb<�Ob<'Hb<�Ab<c>b<>b<??b<Ab<JBb<�Bb<hCb<�Eb<�Jb<�Rb<J\b<�cb<�db<FYb<h<b<M
b<�a<:ca<��`<5|`<�`<��_<�8_<��^<��^<��^<Z_<�J_<|�_<y`<ٖ`<�a<�ya<��a<<b<�Eb<d_b<�hb<�fb<_b<�Vb<tPb<Mb<�Lb<Mb<�Mb<�Mb<�Lb<Mb< Ob<gTb<5\b<�db<�ib<|fb<�Tb<�0b<�a<9�a<�@a<��`<�S`<l�_<s_<�_<z�^<R�^<Z�^<�_<�h_<K�_<�E`<s�`<�3a<ؙa<��a<�)b<Pb<�cb<hb<cb<�Zb<�Rb<)Mb<�Jb<OJb<�Jb<!Kb<)Jb<�Ib<�Ib<�Lb<�Rb<�Zb<hbb<=eb<y]b<�Eb<�b<D�a<|�a<^a<
�`<I&`<�_<rO_<�_<��^<o�^<e�^<�*_<��_<!�_<�h`<��`<�Qa<��a<`�a<2b<Qb<�^b<�^b<�Wb<%Nb<�Eb<j@b<>b<:=b<=b<3<b<m:b<H9b<j9b<�<b<�Bb<pJb<QPb<�Ob<*Bb<�#b<�a<Z�a<,Fa<N�`<�\`<4�_<s_<1_<��^<�^<d�^<?�^<�$_<[�_<��_<�o`<m�`<�Qa<��a<1�a<Xb<85b<�=b<0;b<3b<*b<H#b<Ub<Xb<Pb<�b<b<$b<�b<�b<�#b<n+b<�3b<�8b<-5b<+#b<��a<*�a<,sa<ya<I�`<h!`<Ȫ_<�@_<�^<Ѷ^<Ţ^<��^<��^<�6_<��_<�`<��`<�  �  �a<�qa<��a<��a< %b<#7b<(:b<4b<�)b<�b<�b<�b<�b<�b<ub<�b<�b<rb<Ob<g%b<�0b<:;b<�@b<�;b<P&b<��a<�a<ga<��`<��`<(`<
�_<�@_<��^<��^<��^<�^< _<�y_<T�_<�]`<+�`<SFa<�a<x�a<�'b<Gb<kTb<�Tb<�Mb<�Cb<;b<H5b<�2b<�2b<�3b<�4b<�5b<�7b<)<b<�Cb<Nb<�Yb<}cb<Ffb<�\b<�@b<�b<o�a<|ka<�`<~�`<�`<)�_<hH_<q_<�^<��^<�_<Z_<��_<�)`<ˡ`<a<��a<��a<�b<*Jb<,bb<�ib<�eb<6\b<tQb<�Hb<'Cb<�@b<@b<V@b<F@b<�@b<2Bb<�Fb<Nb<FXb<�bb<�ib<hhb<bXb<z5b<\�a<��a<VIa<��`<�_`<��_<x�_<�/_<>�^<f�^<-�^<(_<�w_<��_<�Q`<��`<I<a<��a<Y�a<�.b<�Sb<�eb<ehb<�ab<ZWb<�Lb<�Db< @b<�=b<�=b<�=b<=b<�=b<�?b<�Db<Mb<�Wb<Gab<�eb<`b<�Ib<�b<�a<�a<\a<ɪ`<�2`<��_<�^_<"_<u�^<{�^<��^<o:_<h�_<�_<`t`<g�`<*Za<C�a<Bb<�6b<Tb<`b<k^b<oUb<�Ib<?b<O7b<�2b<�0b<�/b<�.b<�-b<�-b<0b<�5b<>b<Hb<�Ob<�Pb<cEb<3(b<��a<��a<mNa<��`<h`<�_<��_<&_<A�^<�^<W�^<��^<m4_<��_<[`<�z`<��`<�Ya<�a<��a<� b<8b<�>b<L:b<=0b<�$b<�b<pb<sb<`b<5b<�b<�b<b<&b<�b<�'b<�1b<�8b<7b<�&b<�b<~�a<�za<a<e�`<4-`<�_<�O_< �^<��^<Գ^<��^<��^<�E_<@�_<� `<��`<�  �  �%a<Q�a<��a<�b<C/b<�<b<�:b<�.b<�b<�b<��a<}�a<j�a<]�a<��a<��a<��a<��a<Mb<b<&&b<?7b<�Bb<cBb<�1b<�b<��a<�}a<[a<��`<�6`<�_<�l_<�&_<��^<��^<�_<�M_<]�_<�`<=`<��`<�^a<M�a<b<|4b<�Ob<�Xb<bSb<�Eb<F5b<�%b<�b< b<�b<zb<mb<�b<�b<. b<�-b<�>b<�Qb<�ab<�ib<�db<jMb< b<v�a<t�a<Za<j�`<�5`<��_<�u_<8_<_<�_<�B_<l�_<�_<N`<��`<[2a<��a<��a<�,b<�Ub<uib<�kb<Ubb<YRb<�@b<k1b<�%b<cb<Wb<�b<ub<�b<�"b<w,b<i:b<hKb<�\b<�ib<�mb<3bb<3Cb<�b<A�a<�ba<��`<�`<e`<<�_<�]_<�*_<�_<�&_<tV_<ڢ_<�`<�t`<�`<Va<c�a<5b<�<b<0^b<qkb<ib<�\b<?Kb<�9b<`+b<� b<tb<�b<�b<b<�b<�!b<�,b<�;b<�Lb<C]b<�gb<�fb<%Ub<�.b<��a<�a<!:a<�`<OV`<��_<Ǌ_<D_<>_<�_<�-_<�g_<G�_<�#`<Ε`<8a<�ra<��a<�b<�Cb<X]b<1db<4]b<�Mb<F;b<�)b<�b<b<�b<kb<Vb<�b<pb<b<�b<�.b<�?b<�Mb<fTb<�Mb<�4b<�b<��a<afa<�`<�`< `<�_<S_<�_<0�^<=�^<�_<�`_<��_<�'`<��`<�
a<�pa<<�a<�b<3,b<R?b<+Ab<�6b<h&b<?b<Kb<>�a<0�a<��a<��a<��a<��a<|�a< �a<�	b<�b<�+b<�8b<M<b<�0b<�b<��a<,�a<i0a<+�`<�O`<��_<|z_<(+_<��^<
�^<5�^<?$_<�p_<Q�_<PC`<>�`<�  �  RLa<�a<o�a<}!b<�<b<(Cb<*9b<�#b<�b<z�a<��a<{�a<�a<��a<ƪa<u�a<�a<o�a<��a<7�a<�b<�.b<�Bb<LJb<O@b<,!b<��a<ڞa<�Aa<��`<�m`<8`<O�_<�p_<_K_<;E_<f^_<�_<��_<:F`<��`<"a<�a<��a<b<)Fb<�Zb<X\b<�Nb<�7b<%b<b<��a<S�a<��a<��a<��a<��a<�a<��a<�	b<�%b<iBb<\b<�lb<ob<g^b<�7b<r�a<�a<�Da<��`<$o`<�`<�_<C�_<dg_<�j_<>�_<��_<!`<م`<_�`<N[a<��a<m	b<�Bb<Ceb<rb<�lb<�Zb<�@b<%b<b<��a<+�a<~�a<��a<H�a<��a<��a<|b< b<�5b<Qb<agb<sb<�nb<UVb< 'b<E�a<��a<F"a<J�`<OM`<��_<N�_<�v_<,e_<�r_<]�_<*�_<�A`<��`<~a<�|a<#�a<b<�Pb<}kb<�qb<`gb<�Qb<y6b<�b<�b<��a<�a<�a<��a<��a<��a<{�a<b<�b<e:b<�Tb<�gb<�nb<�cb<Db<�b<I�a<Tba<�`<#�`< '`<i�_<��_< h_<a_<Vy_<	�_<p�_<	^`</�`<j3a<��a<K�a<�+b<WUb<[hb<hb<�Xb<�?b<'#b<b<��a<X�a<��a<��a<��a<��a<��a<��a<��a<�b<�0b<lHb<TWb<�Wb<�Eb<Jb<��a<��a<z&a<i�`<�N`<f�_<��_<	`_<vC_</F_<h_<�_<��_<>_`<P�`<�3a<a<��a<�b<�;b<Hb<EBb<|/b<�b<��a<��a<�a<�a<߭a<��a<۪a<ѱa<��a<-�a<v�a<�b< b<A6b<�Ab<==b<�$b<6�a<'�a<[Va<��`<��`<�`<�_<{s_<�C_<�2_<{@_<m_<.�_<�`<Sx`<��`<�  �  <za<��a<�b<�5b<Ib<�Fb<d2b<�b<��a<D�a<��a<�|a<fa<�Xa<�Ua<�[a<�ka<�a<i�a<��a<|�a<b<N>b<Pb<�Nb<;7b< 	b<��a<�qa<�a<ر`<.V`<`<7�_<�_<��_<)�_<4�_<�6`<ˎ`<��`<jRa<ܭa<��a<�4b<�Wb<�db<�\b<aDb<u!b<��a<c�a<��a<'�a<G�a<?xa<�xa<�a<ܖa<i�a<��a<� b<�*b<_Pb<�kb<�wb<Gob<lPb<pb<��a<xa<.a<��`<!^`<w`<��_<��_<��_<s�_<e#`<p`<$�`<_,a<N�a<d�a<|(b<�Yb<Jtb<�xb<�ib<iLb<&b<:�a<��a<n�a<�a<C�a<��a<>�a<��a<��a<��a<>�a<�b<T=b<`_b<�ub<ezb<�ib<�Bb<b<��a<�Xa<�`<�`<�C`<	`<W�_<��_<�_<��_<,;`<��`<��`<1Ma<ƪa<��a<�;b< eb<�wb<[ub<�`b<x?b<_b<f�a<O�a<
�a<�a<a�a<�a<�a<��a<�a<��a<f�a<,b<�Db<gcb<]tb<rb<
Zb<+b<��a<K�a<�2a<I�`<�t`<6&`<��_<��_<~�_<!�_<8	`<�O`<��`<�a<�ga<��a<Db<�Eb<gb<%rb<Jhb<;Nb<j)b<��a<o�a<��a<-�a<Da<1ta<�ra<�za<��a<I�a<��a<��a<�b<�<b<nVb<�`b<�Vb<6b<��a<��a<�Ya<��`<�`<�<`<��_<G�_<ť_<$�_<L�_<��_<�I`<��`<Pa<�da<l�a< b<�0b<�Jb<�Nb<?b</!b<K�a<��a<�a<��a<�la<�[a<�Ta<�Va<�ba<�xa<��a<��a<B�a<fb<@.b<RDb<�Hb<8b<�b<��a<9�a<O&a<[�`<Me`<`<"�_<|�_<�_<��_<o�_<	`<�[`<+�`<>a<�  �  �a<�a<&b<�Fb<YPb<�Cb<L$b<��a<��a<�a<�Ta<�(a<a<��`<-�`<��`<�a<4a<�ba<�a<��a<b<�2b<BOb<Xb<Jb<j%b<�a<��a<�Pa<��`<�`<�i`<)8`< `<}`<�*`<U`<��`<��`<j3a<Y�a< �a<�b<�Kb<�eb<�hb<�Ub<.2b<�b<��a<S�a<Rda<a<a<� a<�a<�a<�!a<�=a<�fa<��a<��a<�	b<�<b<db<�zb<|b<Sfb<D:b<��a<��a<OYa<a<ܸ`<bz`<�N`<y9`<<`<2V`<K�`<#�`<�a<�ka<�a<
b<�Eb<�mb<�~b<1yb<F_b<�5b<�b<��a<�a<�da<�?a<�'a<a<e!a<�3a<eSa<�~a<^�a<,�a<� b<�Ob<Qqb<��b<�yb<�[b<P(b<1�a<��a<==a<��`<n�`<�i`<BE`<�7`<yB`<<d`<ƚ`<��`<3a<Q�a<��a<4 b<�Ub<�ub<Eb<1rb<wRb<�$b<7�a<�a<��a<#Ua<�3a<�a<�a<�"a<@9a<�\a<�a<e�a<2�a<�,b<�Wb<�sb<�{b<�lb<yGb<zb<��a<�pa<ma<��`<�`<�U`<�8`<_3`<�E`<o`<��`<n�`<Ja<��a<��a<;.b<�\b<�tb<vb<�ab<<b<�	b<��a<b�a<`fa<i<a<�a<�a<�a<�a<�3a<�Za<܊a<��a<��a<)b<�Nb<|cb<9cb<�Kb<wb<��a<8�a<�9a<[�`<9�`<�W`<f+`<z`<y`<1`<�``<��`<�`<�Da<��a<$�a<�b<�Db<gUb<2Ob<�4b<�
b<�a<��a<ga<?7a<�a<�`<2�`<�`<	a<r#a<sNa<�a<y�a<��a<�b<�?b<Ob<�Gb<�)b<�a<ða<�_a<u
a<׷`<to`<�6`<O`<�`<�`<�1`<�h`<��`<�a<OWa<�  �  A�a<�b<v9b<Pb<�Ob<;8b<&b<%�a<�a<Ga<Aa<��`<[�`<��`<~`<��`<
�`<��`<Ta<|Za<,�a<��a<Zb<=Fb<�Yb<�Ub<3;b<�b<�a<��a<OFa<7a<5�`<��`<��`<�`<�`<�`<��`<6/a<�ua<s�a< b<�6b<�[b<�kb<Fdb<�Fb<�b<��a<ݓa<FNa<�a<g�`<l�`<M�`<>�`<��`<��`<�a<?Pa<��a<��a<�b<�Sb</ub<�b<;ub<�Sb<� b<@�a<
�a<5Ta<|a<-�`<�`<ȭ`<�`<��`<��`<�!a<�ba</�a<��a<�,b<�\b<[zb<��b<Dqb<)Lb<�b<��a<��a<�Ga<�
a<��`<�`<�`<��`<��`<��`<d,a<�na<׵a<��a<`7b<�db<�~b<�b<'nb<�Eb<b<��a<΂a<�>a<"a<��`<��`<��`<B�`<F�`<��`<�6a<0za<-�a<�b<"?b<8ib<ub<�~b<�fb<J;b<��a<}�a<#ta<�0a<��`<�`<ð`<Ψ`<��`<}�`<�a<^=a<āa<��a<Wb<LCb<kjb<}b<jxb<7]b</b<��a<��a<�ea<$a<[�`<u�`<V�`<ԧ`<��`<��`<�	a<%Ga<f�a<��a<b<*Ib<�lb<{b<�qb<{Rb<� b<��a<�a<YRa<a<q�`<k�`<A�`<'�`<k�`<��`<�a<$Ba<{�a<��a<b<>b<�]b<>hb<�Zb<8b<Mb<��a<gza<3a<��`<��`<��`<��`<F�`<��`<�`<��`<�;a<"�a<0�a<b<�4b<{Qb<&Xb<TGb<�!b<��a<#�a<�`a<a<n�`<�`<��`</}`<�`<^�`<�`<8�`<B>a<,�a<��a<@b<Q3b<'Mb<JPb<<b<�b<��a<;�a<�Oa<�a<�`<��`<��`<�y`<�`<��`<��`<a<�Ha<�a<�  �  �a<f%b<GDb<8Pb<�Eb<E$b<��a<2�a<�Ta<=�`<=�`<Mh`<�2`<�`<�	`<�`<�>`<�x`<^�`<�a<�ka<~�a<xb<�4b<�Qb<,Xb<xHb<�&b<��a<��a<ϊa<?Xa<I.a< a<u�`<��`<	a<�"a<�Ia<cza<��a<��a<Eb<Ib<cb<whb<Wb</b<�a<`�a<�Ua<�a<t�`<\t`<DF`<].`<.`<�E`<~s`<��`<�a<�Wa<��a<��a<�:b<�fb<�|b<a{b<eb<G>b<�b<Y�a<˝a<(ma<Fa<�+a<�a<3 a<�/a<+Ma<�va<̨a<��a<b<�Gb<zkb< ~b<�zb<�`b<�0b<��a<؞a<�Ia<Z�`<�`<�p`<�H`<p7`<Q>`<~\`<'�`<��`<%%a<�za<W�a<~b<�Ob<�sb<�b<�wb<[b<j/b<<�a<C�a<�a<2_a<�;a<�%a<�a<9$a<�8a<4Za<Նa<R�a<�a<�(b<�Ub<tb<�b<�tb<�Rb<�b<��a<݁a<2,a<��`<k�`<�^`<�=`< 4`<�B`<�g`<��`<N�`< =a< �a<!�a<U&b<�Xb<1ub<�zb<qjb<CHb<�b<��a<@�a<wa<uLa<�-a<5a<�a<-$a<
=a<�ba<]�a<p�a<��a<N3b<�[b<�sb<�wb<�db<�:b<�a<d�a<�[a<�a<��`<ht`<ED`<R*`<�'`<p=`<Xi`<Ч`<��`<�Ga<�a< �a<$%b<�Ob<�cb<�`b<%Ib<!b<R�a<��a<}a<pKa<t#a<7a<��`<��`<�
a<o'a<VPa<,�a<�a<��a<�b< Cb<*Ub<lQb<�6b<b<��a<@sa<�a<��`<�~`<�B`<K`<�`<,`<�,`<S``<��`<��`<Ja<u�a<_�a<(b<Bb<<Ob<�Eb<�(b<��a<u�a<O�a<�Ya<,a<�a<��`<��`<]�`<�a<�'a<�Ta<ĉa<��a<�  �  9b<�2b<�Fb<dHb<T4b<�	b<��a<�va<�a<�`<�Y`<7`<)�_<�_<��_<�_<��_<	`<�p`<b�`<�2a<��a<��a<	b<�Bb<�Rb<kMb<7b<1b<f�a<s�a<'�a<�a<poa<qda<(ca<_ka<�}a<��a<��a<�a<	b<5b<�Rb<
bb<Q]b<�Bb<�b<��a<�ta<�a<W�`<�[`<�`</�_<�_<q�_<��_<`<�Y`<U�`<>a<xa<t�a<zb<�Qb<{pb<>yb<�mb<�Rb<�-b<b<X�a<��a<��a<A�a<��a<��a<�a<R�a<��a<�a<Lb<�5b<*Yb<�qb<yyb<rlb<*Ib<�b<%�a<&ga<�a<ѥ`<gO`<.
`<~�_<y�_<\�_<��_<�.`<�~`<��`<u=a<��a<��a<�3b<]ab<.xb<@yb<Qgb<-Hb< !b<�a<j�a<	�a<Řa<��a<E�a<c�a<C�a<n�a<��a<��a<ub<�Bb<cb<�vb<�wb<Acb<8b<��a<x�a<Fa<�`<�`<B4`<��_<*�_<�_<��_<� `<�C`<`�`<z�`<Ya<�a<�b<@b<�eb<1ub<[ob<XXb<�5b<tb<��a<��a<O�a<�a<9�a<%a<��a<��a<��a<��a<��a<�#b<"Ib<[eb<sb<�lb<?Pb<�b<��a<�|a<�a<p�`<�]`<`<0�_<�_<Z�_<��_<�`<�M`<5�`</a<*fa<��a<�b<G:b<�Wb<�^b<�Qb<c5b<=b<b�a<��a<��a<}a<�ia<�`a<�`a<�ja<�~a<Úa<l�a<A�a<_b<I1b<:Ib<�Pb<'Cb<Xb<��a<4�a<�;a<��`<'y`<1"`<r�_<F�_<Θ_<I�_<r�_<�_<�N`<K�`<�a<�ka<d�a<Ob<�/b<KFb<Gb<�4b<�b<'�a<�a<=�a<�}a<{ea<[Va<#Qa<pUa<�ca<{a<Úa<.�a<E�a<�  �  �#b<9b<�Bb<u;b<�b<��a<��a<YHa<��`<�t`<2`<Ͳ_<m_<�B_<7_<�J_<9|_<��_<Y&`<F�`<��`<;ca<��a<� b<�/b<kGb<rKb<�?b<�)b<�b<��a<i�a<��a<��a<��a<2�a<B�a<;�a<	�a<��a<#b<�'b<�Bb<hUb<�Zb<�Mb<D+b<i�a<��a<WCa<��`<zo`<+`<ڸ_<�|_<�\_<6\_<�z_<+�_<T	`<_m`<��`<�Ea<J�a<�a<99b<`b<�pb<ob<_b<QFb<�*b<=b<��a<b�a<��a<��a<�a<'�a<��a<��a< b<0b<�Kb<cb<�pb<5ob<CZb<�.b<��a<Жa<@2a<��`<�\`<��_<��_<n{_<�d_<�m_<��_<w�_<;1`<�`<a<ma<Q�a<�b<�Kb<jjb<tb<^lb<�Xb<�=b<2"b<�b<�a<~�a<��a<��a<��a<��a<��a<Vb<Vb<�9b<�Tb<Sib<{rb<�jb<Nb< b<��a<va<�a<��`<�9`<��_<��_<�m_<�a_<kt_<e�_<��_<N`<J�`<#a<��a<G�a<�$b<�Rb<�ib<Zmb<�`b<7Jb<�.b<`b<?�a<��a<A�a<g�a<8�a<l�a<r�a<8�a<�b<�!b<�=b<�Vb<hb<�kb<(]b<�8b<:�a<��a<cKa<�`<�s`<B`<�_<�z_<�X_<V_<�r_<�_<*�_<<_`<��`<�3a<�a<r�a<�!b<0Gb<�Vb<"Sb<�Ab<�'b<�
b<j�a<�a<��a<2�a<��a<Z�a<ߺa<7�a<Y�a<^�a<�b<$b<%;b<fHb<rFb<1b<b<2�a<�ka<�a<��`<0`<��_<�_<GM_<\6_<�>_<"f_<��_<2`<�g`<��`<A<a<3�a<��a<b<�8b<�Ab<�9b<�%b<b<�a<S�a<��a< �a<F�a<S�a<Ҩa<$�a<;�a<?�a<��a<�b<�  �  .b<>:b<�;b<�-b<Vb<n�a<q�a<F!a<β`<;?`<0�_<4o_<c$_<��^<��^<��^</4_<K�_<��_<�\`<��`<�=a<�a<��a<�b<@;b<]Fb<�Bb<�5b<%b<�b<�b<�a<�a<��a<(�a<��a<��a<�b<�b</&b<�8b<�Ib<�Sb<�Qb<�=b<�b<f�a<;�a<a<ɩ`<Q7`<��_<As_<(2_<�_<_<�/_<�o_<P�_<_4`<��`<pa<�a<c�a<&"b<�Ob<*gb<�lb<eb<Vb<�Db<�4b<�(b<Y b<�b<�b<�b<+b<>!b<5*b<<7b<�Gb<�Xb<gb<plb<�cb<0Hb<wb<��a<�qa<�a<Ǔ`<�!`<5�_<h_<�/_<}_<!_<�K_<$�_<n�_<�a`<��`<FEa<t�a<�a<�6b<�[b<�lb<�lb<�ab<Qb<�?b<�0b<�%b<�b< b<�b<�b<�b<O$b<�.b<�<b<Nb<�^b<�jb<�kb<']b<C:b<� b<��a<�Na<	�`<l`<��_<"�_<�O_<m!_<�_<x(_<J]_<��_<�`<��`<��`<ca<��a<�b<�?b<�]b<?hb<�cb<�Vb< Eb<b4b<�&b<;b<�b<�b<4b<b<=b<�!b<�-b<=b<iNb<�]b<yfb<�bb<JMb<�"b<;�a<3�a<"a<�`<n;`<��_<Qs_<,0_<�_<�_<�'_<�e_<%�_<:&`<w�`<x	a<Pqa<��a<�
b<�6b<�Lb<�Pb<�Gb<�7b<�$b<b<�b<��a<F�a<^�a<��a<��a<u�a<�b<�b<� b<�1b<'?b<(Db<;b<�b<��a<E�a<(Ga<D�`<�g`<c�_<�_<w:_<�_<��^<�^<�_<td_<l�_<V1`<��`<la<Uxa<��a<b<*b<^:b<5:b<�.b<b<zb<h�a<d�a<h�a<��a<b�a<|�a<�a<��a<x�a<;b<�b<�  �  3b<E9b<�5b<F#b<�a<^�a<�ma<?a<I�`<4`<�_<�C_<��^<��^<n�^<��^<O_<�Z_<��_<:`<�`<�$a<�a<��a<Bb<�1b<qAb<�Bb<]<b<U2b<�(b<G"b<�b< b<�b<�b<c b<"b<�%b<,b<p6b<SBb<�Lb<+Qb<Jb<2b<Pb< �a<�ha<t�`<��`<�`<2�_<�F_<�_<��^<��^<R _<C_<+�_<�`<�`<a�`<gma<��a<8b<@Cb<_b<^ib<]gb<�^b</Tb<Kb<�Db<�Ab<�@b<�@b<�@b<�@b<�Ab<<Eb<Lb<�Ub<7`b<�gb<	hb<�Zb<;b<�b<�a<SYa<��`<r`<��_<�_<y:_<��^<H�^<[�^<_<\h_<��_<$>`<��`<�*a<�a<��a<(b<Qb<fb<+kb<fb<\b<sQb<Ib<�Cb<�Ab<3Ab<\Ab<Ab<JAb<Cb<�Gb<�Ob<�Yb<�cb<�ib<�eb<�Rb<�+b<��a<��a<�4a<�`<�H`<<�_<�o_<I!_<��^<��^<E�^<`/_<(�_<+�_<ia`<+�`<�Ia<��a<��a<v2b<4Tb<Ncb<6db<�\b<^Rb<hHb< Ab<=b<�;b<�;b<�;b<�;b<J<b<�>b<�Db<QMb<�Wb<�`b<�cb<"[b<wAb<�b<��a<�ra<�a<Ϗ`<`<M�_<�F_<� _<��^<��^</�^<�8_<��_<b`<�w`<h�`<�Ya<��a<��a<O*b<�Db<gMb<Jb<7@b<d4b<A*b< #b<6b<yb<�b<�b<Jb<�b<b<]%b<�.b<�8b<@b<�?b<�1b<�b<��a<��a<�.a<9�`<)F`<}�_<	d_<�_<��^<÷^<k�^<��^<�8_<��_<�`<�`<��`<�aa<8�a<h�a<b<�3b<�8b<>3b<)b<Bb<�b<�b<Pb<�b<b<�b<lb<�b<�b<�b<�(b<�  �  mgb<�nb<Xlb<�Wb<�(b<-�a<na< �`<�G`<L�_<�_<t^<�^<�]<��]<��]<^<R�^<'_<��_<lp`<�
a<��a<"�a<y=b<�fb<�wb<Ixb<�pb<�hb<�db<�fb<Dnb<�vb<Z}b<.b<;|b<�ub<�nb<�kb<ob<vwb<��b<[�b<��b<�db<�,b<��a<d_a<s�`<�.`<b�_<N�^<l^<�^<A�]<��]<�^<e^<�^<\�_<�(`<s�`<�`a<%�a<9b<vb<��b<�b<��b<
�b<��b<�b<P�b<�b<Q�b<~�b<Ġb<H�b<#�b<��b<{�b<-�b<V�b<��b<�b<��b<�jb<�'b<��a<Da<n�`<`<Gd_<��^<1U^<�^<��]<��]<�+^<c�^<Q _<߿_<�e`<�a<��a<�b<8Sb<��b<D�b<��b<X�b<Q�b<�b<G�b<��b<��b<=�b<�b<��b<�b<ېb<ފb<��b<K�b<�b<�b<�b<��b<dXb<P
b<ǜa<Ga<�u`<��_<�._<��^<�2^<��]<��]<)�]<�F^<X�^<dO_<:�_<�`<�0a<�a<�b<!ab<ډb<-�b<
�b< �b<g�b< �b<p�b<S�b<a�b<*�b<D�b<�b<.�b<H�b<%�b<�b<�b<��b<��b<��b<�tb<`;b<�a<�ia<�`<s5`<Ԏ_<��^<Kl^<�
^<%�]<K�]<V�]<zZ^<c�^<�s_<�`<��`<*La<��a<� b<\b<�zb<b<
b<+ub<zlb<�hb<2kb<�qb<�xb<&|b<�zb<�tb<^lb<�db<bb<deb<9mb<$ub<vb<ygb<1Ab<q�a<ڙa<�a<w�`<��_<7_<�^<�&^<��]<U�]<�]<��]<�d^<��^<ӎ_<�4`<J�`<_a<��a<� b<�Rb<'jb<+nb<�gb<J^b<�Wb<�Vb<�[b<�cb<�jb<amb<Pkb<
eb<6]b<�Wb<�Wb<^b<�  �  Mgb<rqb<=qb<E^b<1b<,�a<�ya<��`<�V`<�_<l_<܈^<�^<s�]<��]<�]<3^<��^<b9_<��_<�~`<Ta<1�a<��a<xEb<Amb<H|b<ozb<pb<�db<\]b<\b<�_b<Ffb<�kb<cmb<kb<Efb<�bb<�bb<dib<$ub<��b<�b<:�b<lb<�5b<�a<hka<��`<J>`<��_<�_<f�^<:#^<��]<@�]<�^<|z^<��^<�_<F8`<%�`<�la<��a<Bb<�}b<X�b<��b<ܞb<�b<@�b<U�b<O�b<��b<Q�b<��b<�b<z�b<v�b<��b<��b<��b<?�b<z�b<(�b<�b<�rb<1b<��a<�Pa<��`<`<Qv_<��^<	k^<�^<i�]<[^<>B^<]�^<Z3_<��_<�t`<�a<��a<�b<�[b<|�b<^�b<��b<��b<C�b<��b<��b<K�b<v�b<��b<�b<+�b<Ĉb<9�b<̀b<�b<�b<��b<��b<֡b<[�b<�`b<Ob<P�a<2 a<��`<\�_<zA_<y�^<I^<^<��]<p^<�\^<��^<�a_<n`<s�`<?=a<T�a<$b<"ib<>�b<��b<2�b<J�b<\�b<�}b<�{b<�~b<��b<��b<w�b<^�b<��b<�|b<,|b<[�b<��b<��b<~�b<0�b<I|b<3Db<��a<�ua<��`<�D`<�_<5_<��^<E!^<��]<��]<3^<�o^<6�^<1�_<�'`<o�`<XXa<k�a<�)b<�cb<��b<��b<N�b<>sb<0gb<0`b<4_b<�bb<�gb<djb<4ib<db<�]b<nYb<&Zb<�`b<"lb<wb<Nzb<�mb<	Ib<�b<�a<(%a<��`<��_<#I_<$�^<�<^<��]<�]<��]<#^<�y^<�_<��_<�C`<\�`<�ja<��a<3)b<�Yb<Cob<'qb<�gb<>[b<UQb<Mb<�Nb<�Sb<DYb<�[b<�Yb<�Tb<�Ob<�Mb<:Qb<�Zb<�  �  Yeb<wb<!~b<�pb<FHb<� b<w�a<�a<.�`<H�_<�J_<��^<�]^<^<�^<)^<�r^<��^<tn_<
`<��`<;a<�a</b<�[b<�~b<ćb<�~b<&lb<MWb<�Eb<�:b<6b<�5b<37b<8b<�8b<$9b<f=b<6Gb<�Wb<mb<`�b<N�b<�b<J�b<VNb<��a<Ќa<�a<�j`<�_<Z;_<&�^<"e^<5^<�3^<�`^<��^<�3_<��_<ne`<xa<�a<:b<[b<R�b<̫b<ܭb<��b<�b<�wb<�gb<$^b<BZb<(Zb<�Zb<>Zb<OYb<�Yb<e^b<
ib<4zb<M�b<�b<�b<��b<��b<-Kb<%�a<�sa<,�`<�F`<��_<>_<V�^<�\^<�:^<5H^<f�^<�^<�j_<�`<�`<�7a<�a<�'b<Nsb<��b<�b<k�b<��b<�b<|qb<�cb<#\b<�Yb<cZb<�Zb<DZb<oYb<[b<�ab<�nb<��b<��b<��b<��b<�b<�wb<�/b<.�a<&Ea<�`<�`<�w_<��^<̉^<�I^<7^<�S^<��^<�_<˖_<�1`<��`<aa<>�a<�>b<qb<��b<$�b<��b<\�b<�wb<fb<�Zb<Ub<,Tb<�Tb<&Ub<�Tb<wTb<�Wb<c`b<�ob<��b<��b<�b< �b<�b<�\b<r	b<a�a<:a<Uq`<u�_<�=_<V�^<-c^<�0^<Q-^<mX^<8�^<M'_<3�_<�T`<��`<Pza<��a<�Bb<Xxb<3�b<��b<�b<Clb<�Vb<~Eb<;b<R6b<z5b<05b<_4b<�2b<�2b<G7b<�Ab<kRb<.gb<�zb<�b<p~b<�^b<� b<N�a<IHa<(�`<�`<}_<q�^<�{^<�-^<�^<s^<BS^<��^<�9_<��_<�n`<�a<�a<��a<�@b<�lb<�|b<xb<�fb<Qb<D=b<//b<�'b<;%b<�%b<$&b<&b<|%b<�'b<�.b<<b<qOb<�  �  �^b<F}b<b�b<��b<�hb<�'b<��a<sMa<��`<-`<͞_<O"_<��^<χ^<8w^<$�^<��^<�=_<,�_<qQ`<C�`<�oa<��a<@b<rzb<��b<ԕb<��b<|bb<?b<b<�b<_�a<��a<��a<��a<��a<j�a<��a<Ob<~8b<#]b<�b<ɜb<`�b<��b<qb<�&b<ؽa<=a<��`<=`<~�_<d_<�^<��^<a�^<f�^<�_<#�_<E`<W�`<�;a<��a<�.b<�~b<o�b<�b<y�b<��b<�}b<Zb<o:b<"b<�b<Gb<Vb<�b<-	b<�b<v%b<|?b<B`b<�b<�b<�b<޽b<�b<Lpb<b<��a<�a<�`<l�_<�w_<[_<O�^<�^<Y�^<-�^<oE_<��_<�L`<��`<oa<=�a<�Ob<o�b<,�b<(�b<j�b<`�b<�qb<�Nb<31b<�b<�b<kb<	b<�b<@b<-b<�-b<WJb<�lb<g�b<Z�b<�b<��b<;�b<Wb<��a<�{a<��`<�Z`<��_<O_<��^<��^<f�^<��^<e _<+g_<��_<y`<a<ؕa<b<~db<1�b<��b<<�b<ƣb<��b<�_b<<>b<2#b<gb<�b<��a<��a<!b<�
b<'b<s1b<ePb<�sb<5�b<X�b<J�b<��b<yb<3b<d�a<�Ea<�`<�`<Δ_<�_<'�^<��^<�^< �^<l_<�_<�`<��`<)a<D�a<b<^fb<z�b<y�b<b�b<2�b<�]b<9b<Yb<�a<��a<��a<�a<��a<��a<��a<[�a<	b<y8b<�[b<a|b<��b<��b<�|b<�Eb<8�a<"|a<t�`<6``<!�_<�I_<��^<_�^<�v^<��^<��^<�_<��_<�`<B�`<s=a<Z�a<�b<�ab<p�b<�b<b<�ab<�=b<�b<��a<%�a<3�a<��a<��a<��a<a�a<��a<��a<�b<�:b<�  �  Ob<@}b<��b<��b<.�b<�Rb<��a<_�a<a<o�`<(`<ɗ_<�B_<G_<��^<|_<bT_<��_<}%`<��`<�.a<3�a<&b<�hb<�b<��b<S�b<�~b<�Nb<
b<��a<c�a<.�a<|a<�oa<Bna<-wa<Ƌa<īa<��a<�	b<~Ab<�vb<p�b<}�b<նb<ɕb<�Tb<7�a<�a<��`<fz`<d�_<Ș_<�N_<w'_<w&_<�K_<��_<{�_<�u`<��`<$�a<v�a<�]b<E�b<��b<e�b<��b</�b<db<�-b<��a<��a<��a<k�a<��a<ޑa<x�a<ϴa<9�a<b<%8b<�nb<�b<��b<��b<��b<�b<iKb<��a<�ga<��`<P_`<��_<B�_<!J_<�._<h9_<j_<U�_<�)`<Ĩ`<�.a<T�a<)"b<�{b< �b<C�b<��b<�b<f�b<�Qb<�b<�a<��a<�a<��a<2�a<��a<8�a<e�a<�a<^b<�Jb<��b<J�b<$�b<��b<ƹb<�b<Q+b<��a<;a<�`<a4`<��_<�n_<:_<+_<(B_<c~_<��_<N`<x�`<�Ua<R�a<y=b<W�b<��b<��b<��b<��b<-pb<�9b<
b<��a<0�a<s�a<g�a<>�a<V�a<�a<��a<��a<�!b<Xb<�b<��b<]�b<��b< �b<�`b<� b<��a<a<�~`<�`<��_<�L_<Z#_<4 _<SC_<��_<��_<Ig`<,�`<wna<��a<#Gb<�b<Ȱb<۶b<��b<�xb<IDb<�b<��a<֬a<��a<�ua<�ka<la<.wa<�a<"�a<��a<[b<rFb<bwb<�b<R�b<�b<�mb<s b<@�a<�;a<�`<�1`<�_<�[_<_<*�^<�	_<�9_<��_<��_<�w`<8�`<�~a<G�a<�Ib<��b<��b<��b<��b<�Sb<b<��a<޶a<L�a<�ra<�aa<�[a<�`a<rpa<��a<}�a<��a<�b<�  �  �2b<1rb<��b<t�b<�b<bxb<f.b<��a<�\a<`�`<�y`<�`<;�_<F�_<�_<�_<}�_<=0`<C�`<�a<�za<l�a<)Gb<��b<;�b<��b<��b<
pb<{.b<��a<ɚa<*Xa<
"a<{�`<6�`<��`<��`<za<�Ca<ׂa< �a<qb<�`b<l�b<�b<b�b< �b<~b<[,b<��a<Ta<L�`<�w`<X `<��_<��_<I�_<��_<�`<�t`<��`<FSa<��a<2b<��b<��b<p�b<I�b<'�b<ۂb<#=b<�a<P�a<�ia<�7a<3a<�a<�a<�a<�@a<�ua<��a<Yb<Lb<p�b<��b<|�b<+�b< �b<$yb<�b<�a<>a<@�`<�f`<$`<�_<��_<�_<�_<�@`<�`<�a<V�a<��a<kUb<��b<��b<A�b<Y�b<��b<mb<S$b<�a<��a<CWa<�*a<�a<na<�a<A&a<Qa<Ίa<�a<�b<9db<.�b<t�b<}�b<{�b<��b<0]b<X�a<�a<a<�`<�G`<��_<;�_<z�_<��_<�`<�Y`<�`<�-a<�a<�b<�lb<��b<�b<��b<5�b<�b<�Ob<Lb<�a<�wa<Aa<�a<�a<��`<	a<�-a<�]a<��a<��a<�.b<�ub<�b<��b<~�b<o�b<��b<�6b<B�a<�Za<��`<
z`<� `<��_<Ӽ_<�_<Z�_<�`<h`<1�`<�Ba<��a<zb<rb<��b<��b<ɿb<%�b<pdb<jb<�a<S�a<�Fa<a<��`<��`<��`<_�`<a<�Na<!�a<��a<�#b<�fb<�b<�b<>�b<��b<Nb<��a<Ӆa<%a<`<�8`<��_<�_<h�_<�_<��_<@`<.m`<��`<�Na<�a<�#b<ypb<��b<��b<m�b<Nwb<�9b<��a<$�a<�^a<#a<B�`<q�`<L�`<��`<��`<�a<�Wa<��a<��a<�  �  Kb<@Yb<Z�b<E�b<��b<l�b<VVb<�b<s�a<�Fa<��`<۟`<Qf`<�C`<<:`<LJ`<�r`<��`<�a<�_a<(�a<�b<�kb<$�b<W�b<۷b<.�b<vSb<��a<סa<2Ba<'�`< `<_k`<|M`<�H`<8]`<�`<��`<� a<�a<�a<I<b<��b<ɺb<0�b<��b<��b<YYb<�b<A�a<�Fa<��`<��`<�y`<-``<�_`<y`<ܩ`<
�`<Fa<��a<�b<�`b<~�b<��b<��b<e�b<��b<p`b<�b<�a<~Ia<��`<��`<{�`<�k`<_n`</�`<��`<^a<�\a<8�a<2b<qb<�b<d�b<�b<��b<k�b<Qb<Z�a<�a<�8a<|�`<�`<�{`<+i`<p`<��`<	�`<.a<�la<$�a<z+b<b<�b<��b<U�b<)�b<8�b<�Db<`�a<��a<�+a<��`<��`< x`<�i`<u`<ݘ`<��`<_!a<E|a<��a<�9b<0�b<��b<J�b<2�b<��b<)�b<O3b<��a<�ta<a<��`<�`<p`<�e`<;u`<�`<%�`<j+a<�a<S�a<�Cb<p�b<��b<N�b<�b<��b<^ub<!b<��a<Tba<�	a<��`<��`<k`<ge`<Ey`<�`<��`<�9a<\�a<s�a<?Qb<�b<��b<B�b<�b<��b<�cb<b<��a<Ka<C�`<�`<�w`<\`<�Y`<�p`<Z�`<r�`<�7a<��a<��a<9Lb<�b<��b<��b<�b<�b<Bb<1�a<0�a<�'a<�`<8�`<�]`<�F`<�H`<�c`<ۖ`<P�`<$5a<l�a<�a<pHb<ߊb<�b<�b<n�b<Iqb<I%b<��a<�ha<�
a<J�`<&w`<CL`<x9`<f@`<$``<J�`<,�`<[;a<��a<��a< Mb<�b<��b<��b<M�b<`b<6b<��a<�Sa<��`<ۧ`<�j`<�C`<�5`<4A`<Te`<|�`<��`<�Ia<ުa<�  �  S�a<2b<	{b<2�b<r�b<��b<)pb<R0b<��a<ܛa<Wa< a<N�`<��`<��`<k�`<��`<�+a<jha<�a<��a< Eb<@�b<��b<��b<0�b<�vb<)b<��a<�Sa<<�`<t`<�`<3�_<�_<��_<Y�_<�_<KN`<��`<�(a<��a<�
b<Ceb<��b<�b<��b<\�b<�xb<�5b<��a<ޢa<cba</a<�a<��`<��`<(a<�/a<�ca<
�a<R�a<�;b<"�b<˹b<��b<��b<��b< �b<�0b<��a<�Sa<��`<�x`<�#`<��_<��_<H�_<��_<�3`<-�`<Q�`<*la<Y�a<�Db<.�b<�b<�b<�b<�b<|vb<�.b<��a<�a<�^a<e/a<�a<�a< 	a< a<gHa<�a<�a<�b<Yb<��b<��b<��b<��b<8�b<�mb<fb<�a<q,a<��`<~Y`<�`<C�_<T�_<��_<^`<OO`<��`<�a<0�a<�b<cb<x�b<2�b<	�b<��b<�b<�^b<�b<��a<��a<=Ka<� a<�a<� a<|a<	(a<bUa<U�a<�a<-#b<ukb<�b<[�b<��b<~�b<��b<�Jb<:�a<�ta<^ a<��`<�7`<~�_<}�_<]�_<Y�_<$`<Vh`<��`<�@a<N�a<�b<�xb<v�b<�b<��b<��b<9�b<>b<�a<;�a<�da<A/a<�	a<��`<��`<�a<P%a<Wa<g�a<��a<
)b<�mb<n�b<��b<��b<F�b<5jb<fb<9�a<�2a<ľ`<�U`<��_<#�_<ʦ_<��_<z�_< `<$f`<��`<^Da<(�a<Ob<!mb<��b<�b<c�b<�b<�Jb<|b<��a<Mna<<0a<� a<w�`<��`<��`<��`<�a<Oa<��a<B�a<k'b<�hb<ʘb<��b<��b<l�b<�:b<�a<dma<��`<�`<�%`<��_<H�_<v�_<ޣ_<��_<:`<�|`<v�`<_aa<�  �  ��a<� b<Vb<�b<T�b< �b<|b<�Mb<�b<L�a<ղa<V�a<�ra<da<o`a<ga<Eya<��a<��a<w�a<;(b<.^b<��b<�b<ߧb<��b<TOb<�a<тa<Ua<T|`<��_<��_<�C_<_<X_<�,_<�o_<M�_<�I`<��`<�Ta<��a<M8b<V�b<z�b<��b<Y�b<6�b<:Yb<�#b<��a<�a<�a<2�a<�a<��a<��a<��a<��a<*�a<�)b<kab<p�b<^�b<6�b<G�b<y�b<w[b<T�a<[a<�`<�v`<R�_<�_<T_<�1_<�5_<!`_<�_<�`<g�`<�a<��a<�b<Rmb<ҭb<$�b<<�b<
�b<b<3Yb<�"b<��a<��a<��a<��a<R�a<9�a<�a<��a<7�a<�b<
Bb<�xb<c�b<��b<.�b<��b<\�b<�=b<D�a<�Sa<D�`<L`<��_<�~_<#D_<�._<�?_<9v_<!�_<�=`<��`<EDa<��a<�1b<k�b<�b<��b<[�b<��b<8|b<�Eb<:b<l�a<��a<��a<b�a<:�a<O�a<Σa<��a<��a<�b<�Ob<��b<u�b<��b<��b<�b<�qb<b<(�a<"a<u�`<`<j�_<b_<�3_<"+_<�H_<��_<I�_<�b`<L�`<�ja<��a<�Kb<	�b<w�b<��b<��b<��b<�ab<�)b<��a<S�a<6�a<5�a<�a<l~a<[�a<�a<��a<��a<b<�Nb<�b<	�b<�b<�b<�b<�>b<�a<�_a<V�`<�T`<��_<Iv_<�/_<�_<S_<�9_<M�_<��_<�j`<��`<Wra<��a<:Db<<�b<�b<��b<��b<�ab<�,b<��a<!�a<{�a<�za<6ga<j_a<�aa<zoa<��a<�a<��a<�b<�Fb<~vb<��b<�b<�b<�\b<�
b<�a<o a<��`<X`<�_<�J_<H_<�^<1_<�B_<(�_<*`<|�`<�a<�  �  OSa<��a<�+b<kb<ϊb<��b<�|b<Y^b<t:b<Db<��a<��a<t�a<`�a<%�a<�a<�a<��a<�b</#b<�Fb<'kb<a�b<ޖb<3�b<�hb<�"b<��a<�@a<��`<�`<�_<�_<��^<؎^<��^<��^<��^<�`_<��_<�y`<6a<r�a<�b<*]b<��b<V�b< �b<�b<�ob<�Lb<-b<Mb<�b<p�a<��a<��a<�a<�b<�b<�3b<Ub<�yb<�b<n�b<.�b<k�b<D|b<�+b<�a<A9a<��`<,`<0�_<�_<H�^<��^<Q�^<��^<4_<��_<4`<h�`<HWa<��a<�?b<��b<v�b<ֿb<:�b< �b<�ub<�Rb<�3b<b<b<�b<	b<:b<
b<b<v)b<Eb<gb<#�b<ڪb<��b<��b<��b<fb<�
b<)�a<w	a<v`<��_<xe_<4 _<h�^<4�^<q�^<��^<BX_<�_<�d`<s�`<��a<��a<\b<�b<g�b<Ͻb<իb<��b<�hb<BFb<�)b<8b<Xb<�b< b<bb<�	b<�b<�-b<�Kb<tnb<ϑb<1�b<ۻb<c�b<��b<�Eb<��a<Cba<Y�`<�?`<m�_<�:_<��^<]�^<��^<u�^<�_<�z_<��_<S�`<v#a<C�a<�b<�nb<��b<��b<P�b<u�b<#xb<+Sb<i1b<�b<�b<q�a<��a<��a<��a<c�a<4b<*%b<eDb<\gb<��b<�b<�b<��b<�`b<�b<ҟa<�a< �`<d�_<rk_<&�^<�^<��^<��^<ڷ^<�_<��_<�`<��`</a<%�a<�b<`b<H�b<�b<وb<�lb<KIb<O%b<�b<��a<�a<c�a<
�a<��a<^�a<�a<E�a<�b<s5b<hYb<�xb<s�b<q�b<ob<S3b<��a<aa<!�`<�B`<H�_<�1_<j�^<��^<�r^<��^<~�^<_%_<��_<�2`<��`<�  �  /a<�a<�b<Kb<rrb<�~b<�wb<�eb<0Pb<r=b<�0b<{*b<)b<*b<�*b<�*b<�*b<�-b<�5b<�Db<YYb<�ob<��b<�b<0tb<�Fb<��a<َa<�a<�q`<
�_<a>_<:�^<u\^<�$^<�^<+@^<-�^<�_<��_<4`<g�`<ba<�a<|8b</ub<��b<��b<�b<�{b<�gb<�Wb<Nb<_Jb<Kb<�Lb<�Mb<zNb<�Ob<	Ub<`b<�qb<��b<7�b<.�b<m�b<֏b<WXb<b<��a<c�`<-c`<,�_<e5_<
�^<bh^<�>^<�C^<Dw^<R�^<�R_<d�_<6�`<Ya<B�a<�b<^gb<��b<�b<e�b<�b<Άb<�rb<�cb<a[b<uXb<�Xb<pYb<lYb<�Xb<Zb<�_b<lb<u~b<�b<�b<�b<8�b<_�b<�?b<��a<�^a<��`<.`<��_<�	_<�^<U^<�:^<�O^<�^<W�^<��_<�`<��`<bNa<��a<5b<{b<
�b<�b<��b<N�b<�~b<}kb<�^b<�Wb<Vb<�Vb<�Vb<Vb<JUb<�Wb<5_b<Mmb<�b<H�b<��b<�b<m�b<qjb<>b<�a<C*a<J�`<*�_<�]_<�^<�z^<B^<�7^<	\^<�^<� _<k�_<�K`<��`<�va<`�a<Jb<�b<סb<�b<M�b<'�b<�mb<�[b<@Pb<Jb<Ib<�Hb<�Gb<Fb<HEb<yHb<lQb<�`b<�tb<��b<�b<_�b<vb<=b<C�a<fma<��`<�B`<m�_<�_<z�^<D^<�^<=^<,Q^<ĭ^<�+_<��_<g]`<�`<�~a<��a<�=b<nnb<?�b<�b<�ob<Zb<IEb<�5b<�,b<S)b<U)b<_)b<�(b<(b<
)b<�.b<�:b<�Lb<Ibb<"ub<�}b<�sb<�Ob<b<ªa<�+a<N�`<��_<`_<��^<]h^<p!^<L^<g^<�^^<��^<1P_<��_<�`<�  �  ��`<Ha<��a<!4b<%`b<Jrb<'rb<hb<�[b<7Sb<[Pb<Sb<�Xb< ^b<�_b<�]b<�Xb<8Tb<[Sb<`Xb<�bb<pb<qyb<,wb<�`b</b<Z�a<<na<�`<�E`<��_<�_<B�^< ^<��]<s�]<~�]<)R^<��^<�b_<�`<&�`<??a<�a<�b<�_b<;�b<D�b<ϋb<6�b<�vb<�pb<�pb<�ub<l|b<��b<�b<d�b<�{b<�xb<.zb<��b<��b<��b<��b<��b<�zb<?b<y�a<Uia<��`<�5`<͒_<��^<~^<�%^<L�]<��]<�5^<Ӗ^<�_<\�_<Y`<��`<#�a<)�a<Ob<��b<��b<e�b<��b<k�b<�b<�b<�b<�b<͋b<юb<ݍb<�b<��b<��b<��b<N�b<y�b<=�b<�b<��b<�kb<%b<v�a<�:a<��`<��_<^_<F�^<\^<�^<R�]<;^<hQ^<w�^<~L_<��_<D�`<�)a<�a<�b<db<��b<��b<�b<Öb<P�b<K�b<~b<k�b<��b<��b<��b<S�b<��b<H~b<�|b<ـb<��b<ܖb<\�b<A�b<
�b<�Rb<b<J�a<pa<�f`<��_<d&_<�^<Q9^<,�]<&�]<W^<m^<��^<a{_<z`<W�`<Ta<@�a<H0b<�ob<]�b<��b<,�b<��b<�|b<�tb<�rb<�ub<lzb<�}b<�|b<xb<Jqb<"lb<�kb<qb<o{b<��b<L�b<��b<ab<�#b<��a<%Ka<C�`<`<q_<L�^<�Z^<�^<T�]<�]<t^<Gp^<��^<��_<21`<��`<s]a<��a<e%b<yZb<�sb<�wb<�ob<�bb<�Wb<Rb<jRb<�Vb<!\b<�^b<c]b<EXb<�Rb<]Ob<�Qb<�Yb<�eb<Vpb<�qb<Ebb<n9b<e�a<��a<�a<�n`<'�_<�*_<��^<e(^</�]<��]<��]<T^<��^<_<��_<�]`<�  �  ��`<�sa<��a<�+b<�Yb<�mb<�ob<`hb<�_b<'Zb<�Zb<�`b<ib<�ob<�qb</ob<�hb<>ab<�\b<�^b<�eb<�ob<Pvb<�qb<�Yb<�&b<�a<vba<��`<�6`<��_<��^<1k^<�^<$�]<��]<l�]<k<^<Ӹ^<�P_<�_<%�`<�2a<��a<`b<�Wb<'}b<,�b<�b<��b<Q{b<�xb<
|b<e�b<I�b<g�b<ǔb<U�b<�b<x�b<��b<��b<��b<��b<��b<��b<'sb<�5b<��a<]a<��`<�%`<#�_<	�^<�h^<^<��]<�]<�^<��^<Z_<2�_<�I`<��`<6za<��a<ZFb<s}b<#�b<�b<�b<�b<�b<?�b<��b<��b<��b<��b<m�b<��b<��b<;�b<Q�b<.�b<	�b<��b<z�b<	�b<�cb<\b<&�a<#.a<��`<E�_<�K_<��^<�E^<v�]<��]<��]<*;^<Ȫ^<�9_<#�_<��`<�a<��a<b<�[b< �b<ǜb<��b<�b<�b<=�b<Z�b<=�b<�b<)�b<؝b<��b<��b<S�b<)�b<�b<��b<q�b<?�b<�b<�}b<Jb<��a<��a<F�`<�W`<ֱ_<8_<�^<�"^<��]<]�]<C^<RW^<��^<zi_<�`<U�`<�Ga<9�a<�&b<�gb<G�b<s�b<u�b<�b<��b<�|b<E~b<��b<I�b<E�b<��b<�b<h�b<�wb<�sb<#vb<%}b<�b<k�b<�{b<qYb<�b<ͻa<�>a<w�`<W`<k__<[�^<dE^<��]<��]<��]<��]<[^<_�^<�|_<�!`<P�`<�Qa<~�a<�b<0Sb<Hnb<�tb<�nb<'eb<�]b<0[b<_b<�fb<Omb<�pb<�nb<�hb<�`b<�Yb<�Xb<�]b<Hfb<nb<kmb<�[b<\1b<��a<T�a<�`<T``<�_<2_<%�^<R^<��]<�]<�]<^<x^<y_<"�_<	O`<�  �  ��`<Ha<��a<!4b<%`b<Jrb<'rb<hb<�[b<7Sb<[Pb<Sb<�Xb< ^b<�_b<�]b<�Xb<8Tb<[Sb<`Xb<�bb<pb<qyb<,wb<�`b</b<Z�a<<na<�`<�E`<��_<�_<B�^< ^<��]<s�]<~�]<)R^<��^<�b_<�`<&�`<??a<�a<�b<�_b<;�b<D�b<ϋb<6�b<�vb<�pb<�pb<�ub<l|b<��b<�b<d�b<�{b<�xb<.zb<��b<��b<��b<��b<��b<�zb<?b<y�a<Uia<��`<�5`<͒_<��^<~^<�%^<L�]<��]<�5^<Ӗ^<�_<\�_<Y`<��`<#�a<)�a<Ob<��b<��b<e�b<��b<k�b<�b<�b<�b<�b<͋b<юb<ݍb<�b<��b<��b<��b<N�b<y�b<=�b<�b<��b<�kb<%b<v�a<�:a<��`<��_<^_<F�^<\^<�^<R�]<;^<hQ^<w�^<~L_<��_<D�`<�)a<�a<�b<db<��b<��b<�b<Öb<P�b<K�b<~b<k�b<��b<��b<��b<S�b<��b<H~b<�|b<ـb<��b<ܖb<\�b<A�b<
�b<�Rb<b<J�a<pa<�f`<��_<d&_<�^<Q9^<,�]<&�]<W^<m^<��^<a{_<z`<W�`<Ta<@�a<H0b<�ob<]�b<��b<,�b<��b<�|b<�tb<�rb<�ub<lzb<�}b<�|b<xb<Jqb<"lb<�kb<qb<o{b<��b<L�b<��b<ab<�#b<��a<%Ka<C�`<`<q_<L�^<�Z^<�^<T�]<�]<t^<Gp^<��^<��_<21`<��`<s]a<��a<e%b<yZb<�sb<�wb<�ob<�bb<�Wb<Rb<jRb<�Vb<!\b<�^b<c]b<EXb<�Rb<]Ob<�Qb<�Yb<�eb<Vpb<�qb<Ebb<n9b<e�a<��a<�a<�n`<'�_<�*_<��^<e(^</�]<��]<��]<T^<��^<_<��_<�]`<�  �  /a<�a<�b<Kb<rrb<�~b<�wb<�eb<0Pb<r=b<�0b<{*b<)b<*b<�*b<�*b<�*b<�-b<�5b<�Db<YYb<�ob<��b<�b<0tb<�Fb<��a<َa<�a<�q`<
�_<a>_<:�^<u\^<�$^<�^<+@^<-�^<�_<��_<4`<g�`<ba<�a<|8b</ub<��b<��b<�b<�{b<�gb<�Wb<Nb<_Jb<Kb<�Lb<�Mb<zNb<�Ob<	Ub<`b<�qb<��b<7�b<.�b<m�b<֏b<WXb<b<��a<c�`<-c`<,�_<e5_<
�^<bh^<�>^<�C^<Dw^<R�^<�R_<d�_<6�`<Ya<B�a<�b<^gb<��b<�b<e�b<�b<Άb<�rb<�cb<a[b<uXb<�Xb<pYb<lYb<�Xb<Zb<�_b<lb<u~b<�b<�b<�b<8�b<_�b<�?b<��a<�^a<��`<.`<��_<�	_<�^<U^<�:^<�O^<�^<W�^<��_<�`<��`<bNa<��a<5b<{b<
�b<�b<��b<N�b<�~b<}kb<�^b<�Wb<Vb<�Vb<�Vb<Vb<JUb<�Wb<5_b<Mmb<�b<H�b<��b<�b<m�b<qjb<>b<�a<C*a<J�`<*�_<�]_<�^<�z^<B^<�7^<	\^<�^<� _<k�_<�K`<��`<�va<`�a<Jb<�b<סb<�b<M�b<'�b<�mb<�[b<@Pb<Jb<Ib<�Hb<�Gb<Fb<HEb<yHb<lQb<�`b<�tb<��b<�b<_�b<vb<=b<C�a<fma<��`<�B`<m�_<�_<z�^<D^<�^<=^<,Q^<ĭ^<�+_<��_<g]`<�`<�~a<��a<�=b<nnb<?�b<�b<�ob<Zb<IEb<�5b<�,b<S)b<U)b<_)b<�(b<(b<
)b<�.b<�:b<�Lb<Ibb<"ub<�}b<�sb<�Ob<b<ªa<�+a<N�`<��_<`_<��^<]h^<p!^<L^<g^<�^^<��^<1P_<��_<�`<�  �  OSa<��a<�+b<kb<ϊb<��b<�|b<Y^b<t:b<Db<��a<��a<t�a<`�a<%�a<�a<�a<��a<�b</#b<�Fb<'kb<a�b<ޖb<3�b<�hb<�"b<��a<�@a<��`<�`<�_<�_<��^<؎^<��^<��^<��^<�`_<��_<�y`<6a<r�a<�b<*]b<��b<V�b< �b<�b<�ob<�Lb<-b<Mb<�b<p�a<��a<��a<�a<�b<�b<�3b<Ub<�yb<�b<n�b<.�b<k�b<D|b<�+b<�a<A9a<��`<,`<0�_<�_<H�^<��^<Q�^<��^<4_<��_<4`<h�`<HWa<��a<�?b<��b<v�b<ֿb<:�b< �b<�ub<�Rb<�3b<b<b<�b<	b<:b<
b<b<v)b<Eb<gb<#�b<ڪb<��b<��b<��b<fb<�
b<)�a<w	a<v`<��_<xe_<4 _<h�^<4�^<q�^<��^<BX_<�_<�d`<s�`<��a<��a<\b<�b<g�b<Ͻb<իb<��b<�hb<BFb<�)b<8b<Xb<�b< b<bb<�	b<�b<�-b<�Kb<tnb<ϑb<1�b<ۻb<c�b<��b<�Eb<��a<Cba<Y�`<�?`<m�_<�:_<��^<]�^<��^<u�^<�_<�z_<��_<S�`<v#a<C�a<�b<�nb<��b<��b<P�b<u�b<#xb<+Sb<i1b<�b<�b<q�a<��a<��a<��a<c�a<4b<*%b<eDb<\gb<��b<�b<�b<��b<�`b<�b<ҟa<�a< �`<d�_<rk_<&�^<�^<��^<��^<ڷ^<�_<��_<�`<��`</a<%�a<�b<`b<H�b<�b<وb<�lb<KIb<O%b<�b<��a<�a<c�a<
�a<��a<^�a<�a<E�a<�b<s5b<hYb<�xb<s�b<q�b<ob<S3b<��a<aa<!�`<�B`<H�_<�1_<j�^<��^<�r^<��^<~�^<_%_<��_<�2`<��`<�  �  ��a<� b<Vb<�b<T�b< �b<|b<�Mb<�b<L�a<ղa<V�a<�ra<da<o`a<ga<Eya<��a<��a<w�a<;(b<.^b<��b<�b<ߧb<��b<TOb<�a<тa<Ua<T|`<��_<��_<�C_<_<X_<�,_<�o_<M�_<�I`<��`<�Ta<��a<M8b<V�b<z�b<��b<Y�b<6�b<:Yb<�#b<��a<�a<�a<2�a<�a<��a<��a<��a<��a<*�a<�)b<kab<p�b<^�b<6�b<G�b<y�b<w[b<T�a<[a<�`<�v`<R�_<�_<T_<�1_<�5_<!`_<�_<�`<g�`<�a<��a<�b<Rmb<ҭb<$�b<<�b<
�b<b<3Yb<�"b<��a<��a<��a<��a<R�a<9�a<�a<��a<7�a<�b<
Bb<�xb<c�b<��b<.�b<��b<\�b<�=b<D�a<�Sa<D�`<L`<��_<�~_<#D_<�._<�?_<9v_<!�_<�=`<��`<EDa<��a<�1b<k�b<�b<��b<[�b<��b<8|b<�Eb<:b<l�a<��a<��a<b�a<:�a<O�a<Σa<��a<��a<�b<�Ob<��b<u�b<��b<��b<�b<�qb<b<(�a<"a<u�`<`<j�_<b_<�3_<"+_<�H_<��_<I�_<�b`<L�`<�ja<��a<�Kb<	�b<w�b<��b<��b<��b<�ab<�)b<��a<S�a<6�a<5�a<�a<l~a<[�a<�a<��a<��a<b<�Nb<�b<	�b<�b<�b<�b<�>b<�a<�_a<V�`<�T`<��_<Iv_<�/_<�_<S_<�9_<M�_<��_<�j`<��`<Wra<��a<:Db<<�b<�b<��b<��b<�ab<�,b<��a<!�a<{�a<�za<6ga<j_a<�aa<zoa<��a<�a<��a<�b<�Fb<~vb<��b<�b<�b<�\b<�
b<�a<o a<��`<X`<�_<�J_<H_<�^<1_<�B_<(�_<*`<|�`<�a<�  �  S�a<2b<	{b<2�b<r�b<��b<)pb<R0b<��a<ܛa<Wa< a<N�`<��`<��`<k�`<��`<�+a<jha<�a<��a< Eb<@�b<��b<��b<0�b<�vb<)b<��a<�Sa<<�`<t`<�`<3�_<�_<��_<Y�_<�_<KN`<��`<�(a<��a<�
b<Ceb<��b<�b<��b<\�b<�xb<�5b<��a<ޢa<cba</a<�a<��`<��`<(a<�/a<�ca<
�a<R�a<�;b<"�b<˹b<��b<��b<��b< �b<�0b<��a<�Sa<��`<�x`<�#`<��_<��_<H�_<��_<�3`<-�`<Q�`<*la<Y�a<�Db<.�b<�b<�b<�b<�b<|vb<�.b<��a<�a<�^a<e/a<�a<�a< 	a< a<gHa<�a<�a<�b<Yb<��b<��b<��b<��b<8�b<�mb<fb<�a<q,a<��`<~Y`<�`<C�_<T�_<��_<^`<OO`<��`<�a<0�a<�b<cb<x�b<2�b<	�b<��b<�b<�^b<�b<��a<��a<=Ka<� a<�a<� a<|a<	(a<bUa<U�a<�a<-#b<ukb<�b<[�b<��b<~�b<��b<�Jb<:�a<�ta<^ a<��`<�7`<~�_<}�_<]�_<Y�_<$`<Vh`<��`<�@a<N�a<�b<�xb<v�b<�b<��b<��b<9�b<>b<�a<;�a<�da<A/a<�	a<��`<��`<�a<P%a<Wa<g�a<��a<
)b<�mb<n�b<��b<��b<F�b<5jb<fb<9�a<�2a<ľ`<�U`<��_<#�_<ʦ_<��_<z�_< `<$f`<��`<^Da<(�a<Ob<!mb<��b<�b<c�b<�b<�Jb<|b<��a<Mna<<0a<� a<w�`<��`<��`<��`<�a<Oa<��a<B�a<k'b<�hb<ʘb<��b<��b<l�b<�:b<�a<dma<��`<�`<�%`<��_<H�_<v�_<ޣ_<��_<:`<�|`<v�`<_aa<�  �  Kb<@Yb<Z�b<E�b<��b<l�b<VVb<�b<s�a<�Fa<��`<۟`<Qf`<�C`<<:`<LJ`<�r`<��`<�a<�_a<(�a<�b<�kb<$�b<W�b<۷b<.�b<vSb<��a<סa<2Ba<'�`< `<_k`<|M`<�H`<8]`<�`<��`<� a<�a<�a<I<b<��b<ɺb<0�b<��b<��b<YYb<�b<A�a<�Fa<��`<��`<�y`<-``<�_`<y`<ܩ`<
�`<Fa<��a<�b<�`b<~�b<��b<��b<e�b<��b<p`b<�b<�a<~Ia<��`<��`<{�`<�k`<_n`</�`<��`<^a<�\a<8�a<2b<qb<�b<d�b<�b<��b<k�b<Qb<Z�a<�a<�8a<|�`<�`<�{`<+i`<p`<��`<	�`<.a<�la<$�a<z+b<b<�b<��b<U�b<)�b<8�b<�Db<`�a<��a<�+a<��`<��`< x`<�i`<u`<ݘ`<��`<_!a<E|a<��a<�9b<0�b<��b<J�b<2�b<��b<)�b<O3b<��a<�ta<a<��`<�`<p`<�e`<;u`<�`<%�`<j+a<�a<S�a<�Cb<p�b<��b<N�b<�b<��b<^ub<!b<��a<Tba<�	a<��`<��`<k`<ge`<Ey`<�`<��`<�9a<\�a<s�a<?Qb<�b<��b<B�b<�b<��b<�cb<b<��a<Ka<C�`<�`<�w`<\`<�Y`<�p`<Z�`<r�`<�7a<��a<��a<9Lb<�b<��b<��b<�b<�b<Bb<1�a<0�a<�'a<�`<8�`<�]`<�F`<�H`<�c`<ۖ`<P�`<$5a<l�a<�a<pHb<ߊb<�b<�b<n�b<Iqb<I%b<��a<�ha<�
a<J�`<&w`<CL`<x9`<f@`<$``<J�`<,�`<[;a<��a<��a< Mb<�b<��b<��b<M�b<`b<6b<��a<�Sa<��`<ۧ`<�j`<�C`<�5`<4A`<Te`<|�`<��`<�Ia<ުa<�  �  �2b<1rb<��b<t�b<�b<bxb<f.b<��a<�\a<`�`<�y`<�`<;�_<F�_<�_<�_<}�_<=0`<C�`<�a<�za<l�a<)Gb<��b<;�b<��b<��b<
pb<{.b<��a<ɚa<*Xa<
"a<{�`<6�`<��`<��`<za<�Ca<ׂa< �a<qb<�`b<l�b<�b<b�b< �b<~b<[,b<��a<Ta<L�`<�w`<X `<��_<��_<I�_<��_<�`<�t`<��`<FSa<��a<2b<��b<��b<p�b<I�b<'�b<ۂb<#=b<�a<P�a<�ia<�7a<3a<�a<�a<�a<�@a<�ua<��a<Yb<Lb<p�b<��b<|�b<+�b< �b<$yb<�b<�a<>a<@�`<�f`<$`<�_<��_<�_<�_<�@`<�`<�a<V�a<��a<kUb<��b<��b<A�b<Y�b<��b<mb<S$b<�a<��a<CWa<�*a<�a<na<�a<A&a<Qa<Ίa<�a<�b<9db<.�b<t�b<}�b<{�b<��b<0]b<X�a<�a<a<�`<�G`<��_<;�_<z�_<��_<�`<�Y`<�`<�-a<�a<�b<�lb<��b<�b<��b<5�b<�b<�Ob<Lb<�a<�wa<Aa<�a<�a<��`<	a<�-a<�]a<��a<��a<�.b<�ub<�b<��b<~�b<o�b<��b<�6b<B�a<�Za<��`<
z`<� `<��_<Ӽ_<�_<Z�_<�`<h`<1�`<�Ba<��a<zb<rb<��b<��b<ɿb<%�b<pdb<jb<�a<S�a<�Fa<a<��`<��`<��`<_�`<a<�Na<!�a<��a<�#b<�fb<�b<�b<>�b<��b<Nb<��a<Ӆa<%a<`<�8`<��_<�_<h�_<�_<��_<@`<.m`<��`<�Na<�a<�#b<ypb<��b<��b<m�b<Nwb<�9b<��a<$�a<�^a<#a<B�`<q�`<L�`<��`<��`<�a<�Wa<��a<��a<�  �  Ob<@}b<��b<��b<.�b<�Rb<��a<_�a<a<o�`<(`<ɗ_<�B_<G_<��^<|_<bT_<��_<}%`<��`<�.a<3�a<&b<�hb<�b<��b<S�b<�~b<�Nb<
b<��a<c�a<.�a<|a<�oa<Bna<-wa<Ƌa<īa<��a<�	b<~Ab<�vb<p�b<}�b<նb<ɕb<�Tb<7�a<�a<��`<fz`<d�_<Ș_<�N_<w'_<w&_<�K_<��_<{�_<�u`<��`<$�a<v�a<�]b<E�b<��b<e�b<��b</�b<db<�-b<��a<��a<��a<k�a<��a<ޑa<x�a<ϴa<9�a<b<%8b<�nb<�b<��b<��b<��b<�b<iKb<��a<�ga<��`<P_`<��_<B�_<!J_<�._<h9_<j_<U�_<�)`<Ĩ`<�.a<T�a<)"b<�{b< �b<C�b<��b<�b<f�b<�Qb<�b<�a<��a<�a<��a<2�a<��a<8�a<e�a<�a<^b<�Jb<��b<J�b<$�b<��b<ƹb<�b<Q+b<��a<;a<�`<a4`<��_<�n_<:_<+_<(B_<c~_<��_<N`<x�`<�Ua<R�a<y=b<W�b<��b<��b<��b<��b<-pb<�9b<
b<��a<0�a<s�a<g�a<>�a<V�a<�a<��a<��a<�!b<Xb<�b<��b<]�b<��b< �b<�`b<� b<��a<a<�~`<�`<��_<�L_<Z#_<4 _<SC_<��_<��_<Ig`<,�`<wna<��a<#Gb<�b<Ȱb<۶b<��b<�xb<IDb<�b<��a<֬a<��a<�ua<�ka<la<.wa<�a<"�a<��a<[b<rFb<bwb<�b<R�b<�b<�mb<s b<@�a<�;a<�`<�1`<�_<�[_<_<*�^<�	_<�9_<��_<��_<�w`<8�`<�~a<G�a<�Ib<��b<��b<��b<��b<�Sb<b<��a<޶a<L�a<�ra<�aa<�[a<�`a<rpa<��a<}�a<��a<�b<�  �  �^b<F}b<b�b<��b<�hb<�'b<��a<sMa<��`<-`<͞_<O"_<��^<χ^<8w^<$�^<��^<�=_<,�_<qQ`<C�`<�oa<��a<@b<rzb<��b<ԕb<��b<|bb<?b<b<�b<_�a<��a<��a<��a<��a<j�a<��a<Ob<~8b<#]b<�b<ɜb<`�b<��b<qb<�&b<ؽa<=a<��`<=`<~�_<d_<�^<��^<a�^<f�^<�_<#�_<E`<W�`<�;a<��a<�.b<�~b<o�b<�b<y�b<��b<�}b<Zb<o:b<"b<�b<Gb<Vb<�b<-	b<�b<v%b<|?b<B`b<�b<�b<�b<޽b<�b<Lpb<b<��a<�a<�`<l�_<�w_<[_<O�^<�^<Y�^<-�^<oE_<��_<�L`<��`<oa<=�a<�Ob<o�b<,�b<(�b<j�b<`�b<�qb<�Nb<31b<�b<�b<kb<	b<�b<@b<-b<�-b<WJb<�lb<g�b<Z�b<�b<��b<;�b<Wb<��a<�{a<��`<�Z`<��_<O_<��^<��^<f�^<��^<e _<+g_<��_<y`<a<ؕa<b<~db<1�b<��b<<�b<ƣb<��b<�_b<<>b<2#b<gb<�b<��a<��a<!b<�
b<'b<s1b<ePb<�sb<5�b<X�b<J�b<��b<yb<3b<d�a<�Ea<�`<�`<Δ_<�_<'�^<��^<�^< �^<l_<�_<�`<��`<)a<D�a<b<^fb<z�b<y�b<b�b<2�b<�]b<9b<Yb<�a<��a<��a<�a<��a<��a<��a<[�a<	b<y8b<�[b<a|b<��b<��b<�|b<�Eb<8�a<"|a<t�`<6``<!�_<�I_<��^<_�^<�v^<��^<��^<�_<��_<�`<B�`<s=a<Z�a<�b<�ab<p�b<�b<b<�ab<�=b<�b<��a<%�a<3�a<��a<��a<��a<a�a<��a<��a<�b<�:b<�  �  Yeb<wb<!~b<�pb<FHb<� b<w�a<�a<.�`<H�_<�J_<��^<�]^<^<�^<)^<�r^<��^<tn_<
`<��`<;a<�a</b<�[b<�~b<ćb<�~b<&lb<MWb<�Eb<�:b<6b<�5b<37b<8b<�8b<$9b<f=b<6Gb<�Wb<mb<`�b<N�b<�b<J�b<VNb<��a<Ќa<�a<�j`<�_<Z;_<&�^<"e^<5^<�3^<�`^<��^<�3_<��_<ne`<xa<�a<:b<[b<R�b<̫b<ܭb<��b<�b<�wb<�gb<$^b<BZb<(Zb<�Zb<>Zb<OYb<�Yb<e^b<
ib<4zb<M�b<�b<�b<��b<��b<-Kb<%�a<�sa<,�`<�F`<��_<>_<V�^<�\^<�:^<5H^<f�^<�^<�j_<�`<�`<�7a<�a<�'b<Nsb<��b<�b<k�b<��b<�b<|qb<�cb<#\b<�Yb<cZb<�Zb<DZb<oYb<[b<�ab<�nb<��b<��b<��b<��b<�b<�wb<�/b<.�a<&Ea<�`<�`<�w_<��^<̉^<�I^<7^<�S^<��^<�_<˖_<�1`<��`<aa<>�a<�>b<qb<��b<$�b<��b<\�b<�wb<fb<�Zb<Ub<,Tb<�Tb<&Ub<�Tb<wTb<�Wb<c`b<�ob<��b<��b<�b< �b<�b<�\b<r	b<a�a<:a<Uq`<u�_<�=_<V�^<-c^<�0^<Q-^<mX^<8�^<M'_<3�_<�T`<��`<Pza<��a<�Bb<Xxb<3�b<��b<�b<Clb<�Vb<~Eb<;b<R6b<z5b<05b<_4b<�2b<�2b<G7b<�Ab<kRb<.gb<�zb<�b<p~b<�^b<� b<N�a<IHa<(�`<�`<}_<q�^<�{^<�-^<�^<s^<BS^<��^<�9_<��_<�n`<�a<�a<��a<�@b<�lb<�|b<xb<�fb<Qb<D=b<//b<�'b<;%b<�%b<$&b<&b<|%b<�'b<�.b<<b<qOb<�  �  Mgb<rqb<=qb<E^b<1b<,�a<�ya<��`<�V`<�_<l_<܈^<�^<s�]<��]<�]<3^<��^<b9_<��_<�~`<Ta<1�a<��a<xEb<Amb<H|b<ozb<pb<�db<\]b<\b<�_b<Ffb<�kb<cmb<kb<Efb<�bb<�bb<dib<$ub<��b<�b<:�b<lb<�5b<�a<hka<��`<J>`<��_<�_<f�^<:#^<��]<@�]<�^<|z^<��^<�_<F8`<%�`<�la<��a<Bb<�}b<X�b<��b<ܞb<�b<@�b<U�b<O�b<��b<Q�b<��b<�b<z�b<v�b<��b<��b<��b<?�b<z�b<(�b<�b<�rb<1b<��a<�Pa<��`<`<Qv_<��^<	k^<�^<i�]<[^<>B^<]�^<Z3_<��_<�t`<�a<��a<�b<�[b<|�b<^�b<��b<��b<C�b<��b<��b<K�b<v�b<��b<�b<+�b<Ĉb<9�b<̀b<�b<�b<��b<��b<֡b<[�b<�`b<Ob<P�a<2 a<��`<\�_<zA_<y�^<I^<^<��]<p^<�\^<��^<�a_<n`<s�`<?=a<T�a<$b<"ib<>�b<��b<2�b<J�b<\�b<�}b<�{b<�~b<��b<��b<w�b<^�b<��b<�|b<,|b<[�b<��b<��b<~�b<0�b<I|b<3Db<��a<�ua<��`<�D`<�_<5_<��^<E!^<��]<��]<3^<�o^<6�^<1�_<�'`<o�`<XXa<k�a<�)b<�cb<��b<��b<N�b<>sb<0gb<0`b<4_b<�bb<�gb<djb<4ib<db<�]b<nYb<&Zb<�`b<"lb<wb<Nzb<�mb<	Ib<�b<�a<(%a<��`<��_<#I_<$�^<�<^<��]<�]<��]<#^<�y^<�_<��_<�C`<\�`<�ja<��a<3)b<�Yb<Cob<'qb<�gb<>[b<UQb<Mb<�Nb<�Sb<DYb<�[b<�Yb<�Tb<�Ob<�Mb<:Qb<�Zb<�  �  �b<[�b<(�b<��b<)hb<�b<X{a<�`<��_<�_<2^<n]<��\<Vw\<�\\<Y�\<l�\<p�]<�d^<�E_<.'`<��`<��a<�(b<)b<t�b<^�b<��b<"�b</�b<��b<)�b<��b<�b<��b<��b<��b<2�b<��b<)�b<]�b<��b<�b<{�b<y�b<��b<=hb<F�a<�_a<��`<��_<��^<_^<W]<O�\<��\<G�\<��\<_K]<L�]<`�^<Z�_<?�`<1]a<s�a<�sb<��b<�b<��b<��b<��b<q�b<)�b<��b<
�b< c<�c<�c<c<D�b<��b<9�b<��b<�b<��b<M�b<��b<�b<]b<��a<�5a<j`<u�_<�^<L�]<�1]<v�\<��\<=�\<��\<ϊ]<K^<'_<!
`<�`<��a<�,b<��b<��b<��b<��b<a�b<Y�b<�b<��b<��b<c<�c<�c<3c<'c<��b<��b<��b<��b<��b<J�b<~�b<��b<i�b<]8b<��a<��`<l `<�=_<�_^<h�]<�]<��\<z�\<{�\<�]<�]<��^<�m_<dN`<�a<�a<zMb<7�b<��b<'�b<��b<��b<x�b<Z�b<��b<��b<�c<fc<�c<[c<��b<�b<��b<��b<V�b<>�b<*�b<q�b<ºb<~wb<�b<�ja<��`<��_<��^<�^<kW]<c�\<΅\<ր\<��\<s@]<+�]<�^<�_<��`<�Ga<��a<-Zb<x�b<-�b<��b<��b<S�b<��b<��b<�b<��b<�b<8�b<��b<��b<y�b<��b<�b<V�b<Y�b<�b<�b<٬b<σb<X2b<Y�a<�	a<�=`<G]_<A{^<۫]<�]<�\<�\\<�o\<��\<�Y]<�^<N�^<�_<��`<�ga<�a<�^b<ߗb<��b<q�b<��b<;�b<��b<ӟb<��b< �b<�b<��b<��b<��b<��b<Y�b<�b<d�b<�  �  ��b< �b<��b<ƨb<�ub<�b<g�a<��`<�`<+'_<�L^<��]<��\<ї\<q}\<��\<�]<�]<�~^<�\_<�;`<�a<"�a<�7b<��b<��b<m�b<��b<��b<֝b<Ȝb<��b<T�b<Q�b<��b<~�b<��b<�b<´b<K�b<��b<ϭb<��b<X�b<��b<5�b<�vb<2
b<nqa<<�`<��_<?�^<�(^<�t]<�\<��\<�\<s�\< i]<�^<4�^<�_</�`<oa<�b<�b<f�b<x�b</�b<[�b<U�b<Q�b<��b<G�b<Z�b<t�b<�c<c<��b<��b<��b<��b<��b<�b<d�b<�b<��b<7�b<�kb<�a<�Ga<�~`<0�_<��^<��]<P]<��\<~�\<��\<�]<�]<�e^<�>_<p`<�`<�a<�<b<�b<��b<J�b<��b<v�b<��b<�b<|�b<��b<2�b<��b<_c<��b<��b<9�b<�b<0�b<C�b<7�b<�b<�b<��b<=�b<�Gb<��a<�a<�5`<QU_<`z^<P�]<�!]</�\<=�\<��\<e=]<��]<k�^<��_<	c`<a/a<��a<\b<��b<�b<8�b<��b<a�b<�b<��b<��b<D�b<��b<��b<��b<j�b<��b<M�b<��b<ѽb<��b<G�b<�b<��b<Z�b<�b<xb<�|a<]�`<��_<
_<J+^<�t]<�\<a�\<z�\<��\<4^]<�^<��^<�_<��`<�Ya<�a<�hb<B�b<��b<��b<y�b<�b<ޡb<?�b<ǯb<�b<n�b<1�b<�b<u�b<��b<��b<��b<i�b<I�b<U�b<��b<ڷb<��b<-Ab<��a<�a<�Q`<�s_<ה^<�]<� ]< �\<i}\<?�\<�\<�v]<^4^<+_<Y�_<��`<Eya<�	b<�lb<��b<L�b<��b<��b<w�b<��b<ӓb<֣b<D�b<��b<��b<0�b<��b<k�b<Еb<q�b<�b<�  �  Φb<��b<l�b<n�b<�b<eBb<�a<�a<�B`<�j_<��^<��]<O]<��\<�\<�]<�k]<^<{�^<Y�_<v`<�<a<f�a< ab<s�b<��b<b�b<��b<�b<��b<;�b<6~b<��b<�b<��b<ܗb<m�b<S�b<�b<�b<��b<S�b<"�b<F�b<��b<��b<�b<#6b<��a<d�`<�`<zB_<{w^<��]<LM]<�	]<q]<;F]<��]<�j^<^5_<�`<�`<�a<�:b<��b<��b<hc<%�b<��b<M�b<�b<"�b<�b<��b<��b<R�b<T�b<²b<d�b<��b<��b<�b<��b<\�b< c<( c<��b<ޔb<�b<�za<�`<�_<�_< H^<e�]<v<]<;]<�]<r]<��]<в^<]�_<(\`<�)a<��a<zgb<i�b<��b<�c<��b<��b<�b<��b<�b<�b<�b<ݷb<��b<w�b<��b<-�b<��b<�b<3�b<N�b<��b<�c<0�b<-�b<,rb<E�a<�<a<kq`<ʘ_<W�^<3^<�{]<�"]<�]<�0]<�]<�0^<u�^<}�_<j�`<!ca<	b<��b<��b<V�b<4�b<�b<��b<ܳb<�b<��b<s�b<��b<u�b<�b<Ұb<קb<��b<l�b<�b<�b<d�b<��b<��b<��b<B�b<eCb<�a<��`<� `<BG_<z^<�]<_K]<�]< ]<�=]<�]<v]^<&_<-�_<��`<e�a<�#b<��b<t�b<��b<��b<��b<�b<��b<��b<��b<g�b<��b<��b<E�b<N�b<��b<�{b<c~b<��b<,�b<J�b<��b<Y�b<M�b<jb<b�a<Oa<}�`<ʹ_<��^<z^<Iy]<�]<�\<1�\<A]<F�]<=�^<�Q_<*`<u�`<Z�a<�4b<(�b<R�b<��b<M�b<1�b<�b<Uxb<Uob<Jqb<0yb<�b<҅b<��b<�zb<orb<�ob<mwb<�b<�  �  �b<X�b<��b<.�b<��b<~b<	 b<R[a<��`<��_<s_<-`^<`�]<�]<�r]<ԗ]<1�]<��^<\9_<�`<6�`<ׇa<�%b<�b<��b<� c< �b<��b<�b<{b<�Sb<s8b</)b<�"b< "b<�"b<T$b<8)b<�5b<�Lb<qb<+�b<��b<��b<8c<jc<��b<�tb<��a<O;a<w`<<�_<�^<9P^<X�]<��]<y�]<�]<�F^<��^<��_<Km`<:5a<��a<^zb<c�b<c<�*c<Dc<+�b<r�b<ܔb<�pb<Yb<`Lb<�Gb<eFb<;Fb<#Gb<�Lb<`[b<�ub<��b<��b<��b<bc<�(c<�c<�b<,^b<,�a<�a<�C`<?{_<+�^<�1^<��]<¢]<̳]<s�]<k^<`(_<�_<�`<fxa<!b< �b<6�b<�%c<�(c<�c<+�b<�b<ˆb<�fb<Sb<nIb<�Fb<Fb<RFb<uHb<Qb<$cb<��b<��b<��b<2c<@%c<�%c<# c<٭b<g/b<M�a<\�`<�_<T:_<��^<h^<s�]<��]<+�]<� ^<��^<qb_<�)`<��`<a�a<dKb<��b<�c<-$c<�c<:�b<��b<Q�b<�tb<�Xb<Ib<?Bb<�@b<�@b<�Ab<�Eb<,Qb<Ugb<#�b<�b<��b<yc<$c<�c<��b<ǁb<��a<hDa<~`<�_<��^<�P^<i�]<z�]<�]<d�]<�;^<��^<i�_<�[`<�!a<r�a<�bb<�b<��b<$c<��b<Z�b<I�b<{rb<.Mb<�4b< 'b<�!b<�b<6b<�b<=%b<Z3b<9Mb<osb<�b<��b<��b<�b<��b<7�b<�2b<!�a<;�`<�`<AM_<��^<k^</�]<�r]<%�]<m�]<N^<��^<2�_<]�`<Fa<a�a<qb<��b<
�b<��b<��b<��b<�|b<�Qb<%1b<pb<�b<�b<jb<�b<eb<ab<�.b<Nb<�xb<�  �  àb<�b<Rc<�c<`c<ֽb<�Jb<��a<Oa<EL`<r�_<�_<��^<�D^<�0^<:Q^<e�^<i#_<�_<�x`<�0a<�a<�mb<u�b<�c<�(c<c<i�b<1�b<�Rb<�b<Z�a<9�a<f�a<��a<.�a<N�a<��a<��a<��a<<b<�b<��b<�c<T3c<�5c<hc<ڷb<�8b<�a<��`<8/`<p�_<��^<��^<�[^<�Y^<y�^<��^<"|_<�%`<�`<��a<�9b<Ծb<Cc<�Jc<yNc<�-c<��b<�b<�bb<�!b<��a<��a<�a<$�a<��a<͵a<c�a<&�a<"-b<apb<-�b<��b<�5c<zOc<Cc<Y
c<<�b<�b<�oa<��`<�`<�`_<d�^<��^<�`^<�o^<$�^<7#_<��_<�h`<!a<}�a<Vmb<��b<�1c<UQc<~Gc<�c<O�b<��b<<Kb<�b<�a<{�a<�a<�a<��a<��a<G�a<Fb<�Bb<Q�b<#�b<�c<�Bc<cPc<�5c<��b<Vzb<��a<�2a<�z`<l�_<�/_<��^<�q^<�\^<�|^<.�^<pM_<G�_<�`<tXa<�b<��b<x�b<!;c<Lc<6c<�c<��b<�sb<l/b<��a<�a<��a<l�a<>�a<��a<��a<�a<Ab<	Ub<��b<��b<"c<.Fc<�Fc<�c<�b< Db<��a<��`<�3`<��_<�^<��^<jW^<nS^<˃^<�^<o_<�`<��`<�a<$b<k�b<�c<|/c<�1c<�c<��b<��b<�@b<g�a<a�a<��a<�a<��a<�a<m�a<��a<&�a<�b<�Gb<_�b<��b<4c<�%c<�c<l�b<�yb<��a<Ca<��`<��_<?2_<�^<�V^<�0^<�>^<�^<��^<�_<�6`<��`<�a<�:b<�b<��b<�c<�c<j�b<ʧb<�]b<b<��a<��a<߉a<Zxa<�ra<Twa<��a<��a<:�a<nb<]Vb<�  �  څb<R�b<# c<�<c</c<��b<Ɏb<	b<�na<u�`<�6`<Ŵ_<�R_<+_<�_<�!_<�f_<T�_<�Y`<P�`<T�a<<.b<^�b<�c<�=c<�Bc<<c<��b<�{b<�b<ױa<�Ya<�a<��`<��`<��`<��`<� a<#>a<�a<!�a<"Yb<�b<�c<EGc<)Wc<;c<��b<�b<��a<�Wa<ݹ`<)`<~�_<�\_<0_<�._<Y_< �_<e"`<;�`<�Ra<��a<��b<g�b<RJc<Wmc<dc<�2c<��b<T�b<�b<7�a<aga<l(a<��`<%�`<E�`<Qa<:3a<eva<��a< 0b<��b<
�b<�>c<Thc<�hc<F<c<&�b<2hb<�a<3a<�`<�`<͞_<�U_<�6_<�B_<z_<��_<�W`<��`<��a<*b<�b<c<�\c<�oc<�Wc<c<�b<__b<�a<כa<IOa<�a<g�`<�`<��`<Qa<�Ga<��a<E�a<�Rb<$�b<c<VQc<�mc<L_c<w#c<:�b<#8b<e�a<��`<�d`<}�_<�_<�C_<�2_<9M_<��_<��_<<�`<�a< �a<	Ub<P�b<�0c<5bc<�fc<7Ac<A�b<c�b<�6b<��a<Vza<�4a<=a<��`<��`<��`<�a<uYa<&�a<
b<�pb<$�b<%c<Zc<)hc<<Jc<�b<1�b<��a<�^a<��`<�+`<˱_<�Z_<�+_<g(_<ZP_<�_<N`<��`<8Aa<S�a</ob<�b<1c<URc<SGc<�c<��b<Iab<?�a<�a<Ca<Na<�`<��`<Z�`<��`<�a<kNa<��a<xb<�mb<��b<ec<[>c<N>c<Ac<��b<�;b<�a<ta<�h`<��_<To_<�%_<%_<�_<�H_<��_<�%`<�`<�[a<��a<M�b<=�b<�)c<�<c<<$c<��b<��b<�*b<!�a<�fa<�a<�`<��`<˳`<��`<��`<#a<�]a<߹a< b<�  �  �Tb<N�b<Kc<�Cc<�Bc<Nc<��b<�Ob<<�a<4Ja<�`<zi`<�`<_�_<��_<j�_<R-`<Z�`<��`<�ja<��a<�ob<��b<�)c<�Nc<�Fc<�c<+�b<�Db<��a<@a<�`< g`<� `<$�_<��_<'`<�G`<��`<a<��a<Wb<>�b<��b<�Dc<fbc<4Sc<�c<l�b<HCb<��a<t?a<��`<rn`<l-`<�`<#`<}+`<~k`<j�`<<a<��a<�Cb<2�b<#c<�cc<�yc<�bc<X!c<Q�b<�Bb<L�a<�=a<U�`<r`<�4`<3`<�`<�>`<l�`<$�`<qWa<��a<�\b<��b<�1c<�jc<Oxc<%Yc<�c<v�b<�)b<l�a<�&a<׸`<Tc`<�+`<�`<,`<CG`<)�`<a�`<�la<��a<sb<�b<w?c<�qc<*xc<�Qc<c<��b<b<��a<�a<t�`<�Y`<�&`<4`<�"`<R`<��`<ga<K�a<ib<�b<��b<sIc<otc<�rc<&Ec<Q�b<�~b<�a<�xa<H�`<V�`<K`<[`<$`<>$`<tX`<��`<5a<`�a<�b<��b<�c<<Oc<+sc<[jc<�5c<��b<�fb<�a<�`a<l�`<͆`<�?`<�`<r`<K*`<�c`<�`<2*a<|�a<�-b<D�b<mc<WWc<Xsc<Ebc<�%c<��b<KLb<k�a<+Da<w�`<�n`<y+`<�`<�`<�"`<�``<V�`<�,a<(�a<�0b<ɩb<�c<�Jc<�^c<KFc<'c<��b<�!b<�a<ya<�`<�L`<`<��_<��_<�`<�Z`<1�`<3/a</�a< 4b<��b<�c<�@c<�Mc<.c<��b<{b<��a<�wa<U�`<͉`<�3`<o�_<#�_<'�_<�`<�^`<��`<�:a<h�a<�@b<`�b<�c<�>c<�Dc<'c<%�b<nab<��a<�\a<��`<Au`<B$`<��_<�_<�_<i`<Tk`<��`<Oa<��a<�  �  �b<A�b<t�b<�0c<�<c<
c<��b<�b<1b<ɶa<�[a<�a<��`<��`<`�`</�`<��`<i#a<�qa<V�a<�7b<��b<3�b<1/c<�Ec<�0c<{�b<�b<k�a<^a<Y�`<�*`<�_<�R_<}_<�_<[8_<��_<=�_<*�`<�a<��a<AVb<��b<�(c<�Sc<�Qc<J'c<��b<y~b<�b<��a<�aa<� a<��`<��`<��`<��`<x a<�aa<��a<�b<�b<�b<p3c<dc<�lc<wHc<��b<��b<��a<�Pa<�`<�$`<0�_<la_<�:_<-?_<�n_<��_<�@`<z�`<xra<�b<��b<�c<VSc<�mc<�\c<?%c<��b<}nb<�b<�a<�Xa<�a<�`<a�`<��`<�
a<�<a<��a<�a<�Ab<h�b<�c<Jc<Cmc<�fc<�2c<��b<�Rb<Ӻa<xa<a�`<��_<��_< O_<�6_<J_<�_<�_<�o`<a<3�a<�Ab<��b<�(c<rac<�lc<�Mc<�c<)�b<!Kb<o�a<?�a<�@a<ma<��`<��`<1�`<Ca<�Ma<e�a<8�a<�_b<��b<lc<�Tc<Fjc<�Tc<�c<��b<Pb<�a<+�`<9K`<��_<�q_<=_<�3_<lU_<��_<g`<4�`<�8a<`�a<5lb<��b<Q;c<�dc<�`c<\4c<��b<t�b<db<@�a<\da<� a<��`<��`<H�`<��`<�a<�Ta<��a<�b<�nb<��b<"c<�Jc<�Qc<�+c<��b<�ab<��a<�.a<�`<� `<8�_<�;_<P_<b_<�G_<*�_<�`<?�`<�Ia<�a<~sb<��b<8)c<CCc<�1c<b�b<3�b<GAb<��a<�ya<�)a<��`<��`<��`<u�`<C�`<�
a<�Qa<��a<�b<�ub<��b<-c<3:c<:3c<��b<
�b<�b<c�a<��`<~K`<��_<x\_<_<�_<X_<tS_<	�_<�;`<��`<�ua<�  �  Y�a<BQb<P�b<�c< c<c<��b<B�b<+Tb<"b<�a<�a<�a<�za<wa<�}a<��a<��a<��a<� b<ib<O�b<��b<�c<K&c<c<��b<�=b<֡a<b�`<�8`<u�_<��^<؉^<K^<&@^<�i^<C�^<K_<��_<e�`<&_a<+b<��b<{�b<�.c<�9c<c<�b<��b<�Zb<�b<F�a<�a<�a<ța<e�a<ça<��a<]�a<{b<y_b<0�b<��b<B-c<�Mc<�Hc<�c<B�b<`5b<e�a<��`<6$`< }_< �^<�^<\e^<�j^<��^<_<��_<<J`<�a<�a<wTb<L�b<c&c<8Mc<�Ic<~#c<��b<�b<�Tb<jb<�a<�a<��a<�a<�a<?�a<��a<j�a<8b<R}b<��b<�c<�=c<Rc<�>c<��b<��b<� b<Ta<K�`<�_<�J_<+�^<~^<�`^<x^<��^<W:_<��_<�`<?a<a�a<˂b<a�b<j8c<PPc<�?c<}c<��b<0�b<�<b<�b<�a<ɷa<!�a<֣a<�a<�a<A�a<�b<�Ib<9�b<��b<�c<?Cc<�Jc< )c<��b<`b<��a<�a<�Y`<��_<m_<��^<�i^<�]^<��^<\�^<)f_<�
`<�`<�va<b<�b<
c<�?c<�Hc<",c<�b<{�b<yab<db<��a<^�a<�a<��a<��a<�a<��a<O�a<Gb<+Nb<Ԗb<w�b<�c<�4c<.c<�b</�b<�b<�oa<��`<`<�X_<�^<wn^<#?^<6D^<p}^<��^<�v_<"`<E�`<<�a<2+b<��b<3�b<}"c<mc<��b<B�b<�ob<�&b<��a<��a<�a<~a<va<�xa<��a<ءa<_�a<�b<�Jb<�b<3�b<c<c<�c<"�b<�^b<��a<�a<�g`<F�_<�_<=�^<.I^<,^<�C^<R�^<h_<��_<T`<za<�  �  �ca<	b<$�b<��b<>�b<��b<3�b<ާb<�wb<eNb<o0b<�b<�b<�b<�b<�b<Vb<�#b<�8b<WZb<��b<Էb<��b<��b<��b<��b<�tb<��a<�Fa<ф`<.�_<F�^<S^<��]<��]<A�]<��]<i^<m�^<#i_<n3`</�`<A�a<JMb<޻b<V�b<c<�c<��b<��b<Їb<�bb< Jb<�<b<A8b<G8b<d9b<�;b<�Ab<Pb<�ib<Ïb<
�b<�b<�c<C)c<�c<�b<vb<��a<!0a<�h`<�_<h�^<�I^<�]<��]<8�]<��]<xg^<1
_<T�_<0�`<vXa<b<��b<0�b<�c<~(c<�c<�b<ѷb<U�b<.ib<�Sb<�Hb<XEb<�Db<!Eb<�Fb<jNb<_b<�{b<4�b<��b<Hc<#c<�)c<c<��b<�Ib<u�a<N�`<�#`<]_<��^<^<�]<��]<[�]<^<p�^<xG_<�`<Y�`<��a<�8b<,�b<~c<|&c<}#c<�c<6�b<��b<:}b<�^b<Mb<�Db<ZBb<�Ab<$Bb<�Db<�Nb<�bb<��b<�b<2�b<?
c<�#c<�c<��b<:�b<b<�ha</�`<��_<�_<�r^<��]<k�]<��]<��]<r5^<r�^<	�_<L`<|a<�a<�ab<q�b<"c<�"c<�c<��b<o�b<��b<Ygb<xLb<0=b<I6b<4b<�2b<�2b<�6b<
Cb<qZb<y~b<��b<��b<s c</c<��b<��b<Xb<y�a<Wa<�F`<�{_<e�^<�$^<��]<��]<��]<��]<�?^<Q�^<�_<�k`<�/a<��a<�eb<��b<��b<�b<��b<R�b<\�b<.]b<Y:b<H$b<�b<�b<�b<�b<7b<}b<�,b<gIb<�qb<p�b<��b<B�b<��b<��b<+�b<�b<�va<�`<��_<~(_<�v^<@�]<W�]<�m]<�]<��]<�e^<_<��_<�`<�  �  �a<c�a<�Gb<T�b<��b<��b<d�b<��b<��b<yb<grb<�ub<�~b<Z�b<@�b<{�b<~b<�vb<�ub<�b<��b<n�b<��b<u�b<��b<��b<8b<�a<��`<�)`<�Q_<��^<��]<�H]<��\<��\<� ]<ݐ]<4^<~�^<x�_<�`<�ka<kb<'�b<h�b<��b<C�b<��b<�b<2�b<.�b<~�b<Q�b<|�b<��b<�b<��b<!�b<��b<��b<��b<��b<��b<��b< c<��b<6�b<)6b<R�a<J�`<]	`<�1_<�i^<\�]<�L]<�]<�]<Qa]<��]<U�^<T__<�7`<(a<��a<�Qb<�b<��b<�c<'�b<��b<A�b<f�b<��b<^�b<�b<�b<�b<f�b<�b<ħb<��b<�b<��b<��b<7�b<�c<;�b<H�b<*�b<�b<�^a<n�`<�_<`�^<;,^<,�]<�1]<�]<'*]<�]<�^<@�^<�_<`<�Ha<��a<�xb<��b<5�b<�c<�b<�b<Һb<�b<
�b<R�b<��b<�b<G�b<�b<©b<��b<ݟb<%�b<�b<��b<(�b<  c<}�b<��b<N[b<��a<�a<(K`<�r_<9�^<3�]<�g]</]<�
]<�=]<٬]<O^<W_<�_<Z�`<s�a<� b<��b<,�b<��b<=�b<��b<��b<��b<әb<�b<��b<��b<]�b<��b<S�b<D�b<�b<��b<b�b<\�b<>�b<��b<�b<��b<Éb<+b<�{a<��`<m�_<�_<�E^<��]<D']<c�\<��\<6:]<�]<yj^< 7_<(`<=�`<A�a<�'b<΍b<��b<V�b<�b<�b<��b<&�b<�tb<�tb<�{b<b�b<��b<�b<�~b<�ub<aqb<�vb<�b<[�b<��b<��b<C�b<�b<�Rb< �a<�*a<Pc`<��_<޶^<��]<}_]<��\<N�\<��\<R]<��]<�^<?t_<�L`<�  �  @�`<#�a<�b<�yb<��b<m�b<i�b<8�b<��b<�b<T�b<��b<d�b<��b<��b<��b<��b<��b<b�b<L�b<9�b<F�b<X�b<��b<��b< rb<�b<�za<��`<��_<�_<�5^<�z]<o�\<��\<9�\<<�\<�8]<'�]<�^<�_<�o`<�8a<�a<Zb<a�b<��b<��b<C�b<��b<�b<I�b<E�b<�b<�b<��b<h�b<l�b<!�b<L�b<��b<�b<��b<y�b<8�b<��b<?�b<~b<i	b<0ia<�`<��_<�^<h^<k]<��\<�\<R�\<U]<ی]<D^<�_<��_<]�`<��a<&b<��b<L�b<�b<��b<G�b<��b<4�b<��b<��b<\�b<��b<�c<�b<?�b<��b<#�b<��b<��b<��b<k�b<*�b<��b<�b<r\b<�a<�*a<�\`<�}_<ڠ^<��]<�:]<C�\< �\<��\< ,]<1�]<��^<d_<�C`<!a<��a<�Nb<:�b<��b<[�b<�b<��b<��b<ۿb<�b<�b<l�b<u�b< c<i�b<W�b<��b<��b<��b<��b<��b<��b<>�b<��b<�b<(0b<F�a<��`<`<�-_<�U^<5�]<~]<�\<�\<�\<�T]<�]<��^<��_<2�`<�Na<N�a<mb<�b<��b<��b<8�b<��b<��b<�b<��b<Q�b<�b<R�b<��b<��b<E�b<C�b<Z�b<��b<��b<.�b<�b<��b<w�b<�ab<p�a<�Ia<;�`<�_<�^<y�]<[F]<<�\<͌\<��\<?�\<^e]<-^<_�^<=�_<p�`<Oea<G�a<�fb<g�b<��b<��b<d�b<�b<�b<��b<1�b<%�b<D�b<��b<��b<n�b<�b<�b<J�b<��b<Z�b<¯b<_�b<��b<�b<)b<��a<��`<�(`<|I_<hl^<��]<]<��\<�x\<?�\<��\<��]<}U^<C1_<8`<�  �  ��`<=�a<ub<�kb<�b<�b<۫b<�b<�b<Ęb<!�b<@�b<��b<K�b<F�b<&�b<0�b<*�b<�b<�b<��b<�b<��b<��b<��b<�cb<+�a<9ia<s�`<>�_<��^<�^<U]]<�\<.{\<zl\<�\<�]<�]<��^<�{_<�[`<�&a<��a<�Kb<S�b<��b< �b<�b<�b<�b<ڻb<��b<�b<P�b<Tc<\c<�c<��b<R�b<��b<��b<��b<��b<��b<(�b<_�b<bob<6�a<*Wa<ܐ`<��_<�^<��]<:M]<��\<5�\<��\<��\<jo]<�(^<C_<�_<�`<}a<=b<��b<��b< �b<$�b<{�b<��b<<�b<��b<��b<��b<c<c<c<�c<��b<w�b<�b<�b< �b<K�b<��b<C�b<��b<WMb<d�a<a<�G`<�f_<Ɇ^<�]<]<ڲ\<_�\<	�\<]<d�]<_n^<�L_<�.`<aa<��a<p?b<��b<C�b<��b<��b<S�b<A�b<��b<��b<��b<�c<�c<dc<�c<�b<?�b<Y�b<Q�b<1�b<v�b<��b<\�b<��b<�b<~ b<ۋa<o�`<��_<�_<�:^<�|]<�\<��\<$�\<�\<�6]<��]<W�^<�_<�r`<�<a<��a<>^b<�b<��b<�b<
�b<��b<�b<|�b<*�b<L�b<U�b<c<�c<H�b<��b<J�b<v�b<��b<��b<{�b<��b< �b<��b<�Rb<@�a<�7a<'p`<��_<�^<��]<y(]<4�\<l\<!s\<��\<�G]<� ^<�^<��_<��`<�Sa<n�a<]Xb<�b<x�b<�b<��b<�b<�b<�b<B�b<l�b<Q�b<��b<��b<�b<�b<@�b<��b<��b<��b<��b<.�b<Q�b<qrb<�b<ѓa<D�`<�`<Y2_<\R^<e�]<y�\<I~\<�W\<�v\< �\<�t]<";^<�_<F�_<�  �  @�`<#�a<�b<�yb<��b<m�b<i�b<8�b<��b<�b<T�b<��b<d�b<��b<��b<��b<��b<��b<b�b<L�b<9�b<F�b<X�b<��b<��b< rb<�b<�za<��`<��_<�_<�5^<�z]<o�\<��\<9�\<<�\<�8]<'�]<�^<�_<�o`<�8a<�a<Zb<a�b<��b<��b<C�b<��b<�b<I�b<E�b<�b<�b<��b<h�b<l�b<!�b<L�b<��b<�b<��b<y�b<8�b<��b<?�b<~b<i	b<0ia<�`<��_<�^<h^<k]<��\<�\<R�\<U]<ی]<D^<�_<��_<]�`<��a<&b<��b<L�b<�b<��b<G�b<��b<4�b<��b<��b<\�b<��b<�c<�b<?�b<��b<#�b<��b<��b<��b<k�b<*�b<��b<�b<r\b<�a<�*a<�\`<�}_<ڠ^<��]<�:]<C�\< �\<��\< ,]<1�]<��^<d_<�C`<!a<��a<�Nb<:�b<��b<[�b<�b<��b<��b<ۿb<�b<�b<l�b<u�b< c<i�b<W�b<��b<��b<��b<��b<��b<��b<>�b<��b<�b<(0b<F�a<��`<`<�-_<�U^<5�]<~]<�\<�\<�\<�T]<�]<��^<��_<2�`<�Na<N�a<mb<�b<��b<��b<8�b<��b<��b<�b<��b<Q�b<�b<R�b<��b<��b<E�b<C�b<Z�b<��b<��b<.�b<�b<��b<w�b<�ab<p�a<�Ia<;�`<�_<�^<y�]<[F]<<�\<͌\<��\<?�\<^e]<-^<_�^<=�_<p�`<Oea<G�a<�fb<g�b<��b<��b<d�b<�b<�b<��b<1�b<%�b<D�b<��b<��b<n�b<�b<�b<J�b<��b<Z�b<¯b<_�b<��b<�b<)b<��a<��`<�(`<|I_<hl^<��]<]<��\<�x\<?�\<��\<��]<}U^<C1_<8`<�  �  �a<c�a<�Gb<T�b<��b<��b<d�b<��b<��b<yb<grb<�ub<�~b<Z�b<@�b<{�b<~b<�vb<�ub<�b<��b<n�b<��b<u�b<��b<��b<8b<�a<��`<�)`<�Q_<��^<��]<�H]<��\<��\<� ]<ݐ]<4^<~�^<x�_<�`<�ka<kb<'�b<h�b<��b<C�b<��b<�b<2�b<.�b<~�b<Q�b<|�b<��b<�b<��b<!�b<��b<��b<��b<��b<��b<��b< c<��b<6�b<)6b<R�a<J�`<]	`<�1_<�i^<\�]<�L]<�]<�]<Qa]<��]<U�^<T__<�7`<(a<��a<�Qb<�b<��b<�c<'�b<��b<A�b<f�b<��b<^�b<�b<�b<�b<f�b<�b<ħb<��b<�b<��b<��b<7�b<�c<;�b<H�b<*�b<�b<�^a<n�`<�_<`�^<;,^<,�]<�1]<�]<'*]<�]<�^<@�^<�_<`<�Ha<��a<�xb<��b<5�b<�c<�b<�b<Һb<�b<
�b<R�b<��b<�b<G�b<�b<©b<��b<ݟb<%�b<�b<��b<(�b<  c<}�b<��b<N[b<��a<�a<(K`<�r_<9�^<3�]<�g]</]<�
]<�=]<٬]<O^<W_<�_<Z�`<s�a<� b<��b<,�b<��b<=�b<��b<��b<��b<әb<�b<��b<��b<]�b<��b<S�b<D�b<�b<��b<b�b<\�b<>�b<��b<�b<��b<Éb<+b<�{a<��`<m�_<�_<�E^<��]<D']<c�\<��\<6:]<�]<yj^< 7_<(`<=�`<A�a<�'b<΍b<��b<V�b<�b<�b<��b<&�b<�tb<�tb<�{b<b�b<��b<�b<�~b<�ub<aqb<�vb<�b<[�b<��b<��b<C�b<�b<�Rb< �a<�*a<Pc`<��_<޶^<��]<}_]<��\<N�\<��\<R]<��]<�^<?t_<�L`<�  �  �ca<	b<$�b<��b<>�b<��b<3�b<ާb<�wb<eNb<o0b<�b<�b<�b<�b<�b<Vb<�#b<�8b<WZb<��b<Էb<��b<��b<��b<��b<�tb<��a<�Fa<ф`<.�_<F�^<S^<��]<��]<A�]<��]<i^<m�^<#i_<n3`</�`<A�a<JMb<޻b<V�b<c<�c<��b<��b<Їb<�bb< Jb<�<b<A8b<G8b<d9b<�;b<�Ab<Pb<�ib<Ïb<
�b<�b<�c<C)c<�c<�b<vb<��a<!0a<�h`<�_<h�^<�I^<�]<��]<8�]<��]<xg^<1
_<T�_<0�`<vXa<b<��b<0�b<�c<~(c<�c<�b<ѷb<U�b<.ib<�Sb<�Hb<XEb<�Db<!Eb<�Fb<jNb<_b<�{b<4�b<��b<Hc<#c<�)c<c<��b<�Ib<u�a<N�`<�#`<]_<��^<^<�]<��]<[�]<^<p�^<xG_<�`<Y�`<��a<�8b<,�b<~c<|&c<}#c<�c<6�b<��b<:}b<�^b<Mb<�Db<ZBb<�Ab<$Bb<�Db<�Nb<�bb<��b<�b<2�b<?
c<�#c<�c<��b<:�b<b<�ha</�`<��_<�_<�r^<��]<k�]<��]<��]<r5^<r�^<	�_<L`<|a<�a<�ab<q�b<"c<�"c<�c<��b<o�b<��b<Ygb<xLb<0=b<I6b<4b<�2b<�2b<�6b<
Cb<qZb<y~b<��b<��b<s c</c<��b<��b<Xb<y�a<Wa<�F`<�{_<e�^<�$^<��]<��]<��]<��]<�?^<Q�^<�_<�k`<�/a<��a<�eb<��b<��b<�b<��b<R�b<\�b<.]b<Y:b<H$b<�b<�b<�b<�b<7b<}b<�,b<gIb<�qb<p�b<��b<B�b<��b<��b<+�b<�b<�va<�`<��_<~(_<�v^<@�]<W�]<�m]<�]<��]<�e^<_<��_<�`<�  �  Y�a<BQb<P�b<�c< c<c<��b<B�b<+Tb<"b<�a<�a<�a<�za<wa<�}a<��a<��a<��a<� b<ib<O�b<��b<�c<K&c<c<��b<�=b<֡a<b�`<�8`<u�_<��^<؉^<K^<&@^<�i^<C�^<K_<��_<e�`<&_a<+b<��b<{�b<�.c<�9c<c<�b<��b<�Zb<�b<F�a<�a<�a<ța<e�a<ça<��a<]�a<{b<y_b<0�b<��b<B-c<�Mc<�Hc<�c<B�b<`5b<e�a<��`<6$`< }_< �^<�^<\e^<�j^<��^<_<��_<<J`<�a<�a<wTb<L�b<c&c<8Mc<�Ic<~#c<��b<�b<�Tb<jb<�a<�a<��a<�a<�a<?�a<��a<j�a<8b<R}b<��b<�c<�=c<Rc<�>c<��b<��b<� b<Ta<K�`<�_<�J_<+�^<~^<�`^<x^<��^<W:_<��_<�`<?a<a�a<˂b<a�b<j8c<PPc<�?c<}c<��b<0�b<�<b<�b<�a<ɷa<!�a<֣a<�a<�a<A�a<�b<�Ib<9�b<��b<�c<?Cc<�Jc< )c<��b<`b<��a<�a<�Y`<��_<m_<��^<�i^<�]^<��^<\�^<)f_<�
`<�`<�va<b<�b<
c<�?c<�Hc<",c<�b<{�b<yab<db<��a<^�a<�a<��a<��a<�a<��a<O�a<Gb<+Nb<Ԗb<w�b<�c<�4c<.c<�b</�b<�b<�oa<��`<`<�X_<�^<wn^<#?^<6D^<p}^<��^<�v_<"`<E�`<<�a<2+b<��b<3�b<}"c<mc<��b<B�b<�ob<�&b<��a<��a<�a<~a<va<�xa<��a<ءa<_�a<�b<�Jb<�b<3�b<c<c<�c<"�b<�^b<��a<�a<�g`<F�_<�_<=�^<.I^<,^<�C^<R�^<h_<��_<T`<za<�  �  �b<A�b<t�b<�0c<�<c<
c<��b<�b<1b<ɶa<�[a<�a<��`<��`<`�`</�`<��`<i#a<�qa<V�a<�7b<��b<3�b<1/c<�Ec<�0c<{�b<�b<k�a<^a<Y�`<�*`<�_<�R_<}_<�_<[8_<��_<=�_<*�`<�a<��a<AVb<��b<�(c<�Sc<�Qc<J'c<��b<y~b<�b<��a<�aa<� a<��`<��`<��`<��`<x a<�aa<��a<�b<�b<�b<p3c<dc<�lc<wHc<��b<��b<��a<�Pa<�`<�$`<0�_<la_<�:_<-?_<�n_<��_<�@`<z�`<xra<�b<��b<�c<VSc<�mc<�\c<?%c<��b<}nb<�b<�a<�Xa<�a<�`<a�`<��`<�
a<�<a<��a<�a<�Ab<h�b<�c<Jc<Cmc<�fc<�2c<��b<�Rb<Ӻa<xa<a�`<��_<��_< O_<�6_<J_<�_<�_<�o`<a<3�a<�Ab<��b<�(c<rac<�lc<�Mc<�c<)�b<!Kb<o�a<?�a<�@a<ma<��`<��`<1�`<Ca<�Ma<e�a<8�a<�_b<��b<lc<�Tc<Fjc<�Tc<�c<��b<Pb<�a<+�`<9K`<��_<�q_<=_<�3_<lU_<��_<g`<4�`<�8a<`�a<5lb<��b<Q;c<�dc<�`c<\4c<��b<t�b<db<@�a<\da<� a<��`<��`<H�`<��`<�a<�Ta<��a<�b<�nb<��b<"c<�Jc<�Qc<�+c<��b<�ab<��a<�.a<�`<� `<8�_<�;_<P_<b_<�G_<*�_<�`<?�`<�Ia<�a<~sb<��b<8)c<CCc<�1c<b�b<3�b<GAb<��a<�ya<�)a<��`<��`<��`<u�`<C�`<�
a<�Qa<��a<�b<�ub<��b<-c<3:c<:3c<��b<
�b<�b<c�a<��`<~K`<��_<x\_<_<�_<X_<tS_<	�_<�;`<��`<�ua<�  �  �Tb<N�b<Kc<�Cc<�Bc<Nc<��b<�Ob<<�a<4Ja<�`<zi`<�`<_�_<��_<j�_<R-`<Z�`<��`<�ja<��a<�ob<��b<�)c<�Nc<�Fc<�c<+�b<�Db<��a<@a<�`< g`<� `<$�_<��_<'`<�G`<��`<a<��a<Wb<>�b<��b<�Dc<fbc<4Sc<�c<l�b<HCb<��a<t?a<��`<rn`<l-`<�`<#`<}+`<~k`<j�`<<a<��a<�Cb<2�b<#c<�cc<�yc<�bc<X!c<Q�b<�Bb<L�a<�=a<U�`<r`<�4`<3`<�`<�>`<l�`<$�`<qWa<��a<�\b<��b<�1c<�jc<Oxc<%Yc<�c<v�b<�)b<l�a<�&a<׸`<Tc`<�+`<�`<,`<CG`<)�`<a�`<�la<��a<sb<�b<w?c<�qc<*xc<�Qc<c<��b<b<��a<�a<t�`<�Y`<�&`<4`<�"`<R`<��`<ga<K�a<ib<�b<��b<sIc<otc<�rc<&Ec<Q�b<�~b<�a<�xa<H�`<V�`<K`<[`<$`<>$`<tX`<��`<5a<`�a<�b<��b<�c<<Oc<+sc<[jc<�5c<��b<�fb<�a<�`a<l�`<͆`<�?`<�`<r`<K*`<�c`<�`<2*a<|�a<�-b<D�b<mc<WWc<Xsc<Ebc<�%c<��b<KLb<k�a<+Da<w�`<�n`<y+`<�`<�`<�"`<�``<V�`<�,a<(�a<�0b<ɩb<�c<�Jc<�^c<KFc<'c<��b<�!b<�a<ya<�`<�L`<`<��_<��_<�`<�Z`<1�`<3/a</�a< 4b<��b<�c<�@c<�Mc<.c<��b<{b<��a<�wa<U�`<͉`<�3`<o�_<#�_<'�_<�`<�^`<��`<�:a<h�a<�@b<`�b<�c<�>c<�Dc<'c<%�b<nab<��a<�\a<��`<Au`<B$`<��_<�_<�_<i`<Tk`<��`<Oa<��a<�  �  څb<R�b<# c<�<c</c<��b<Ɏb<	b<�na<u�`<�6`<Ŵ_<�R_<+_<�_<�!_<�f_<T�_<�Y`<P�`<T�a<<.b<^�b<�c<�=c<�Bc<<c<��b<�{b<�b<ױa<�Ya<�a<��`<��`<��`<��`<� a<#>a<�a<!�a<"Yb<�b<�c<EGc<)Wc<;c<��b<�b<��a<�Wa<ݹ`<)`<~�_<�\_<0_<�._<Y_< �_<e"`<;�`<�Ra<��a<��b<g�b<RJc<Wmc<dc<�2c<��b<T�b<�b<7�a<aga<l(a<��`<%�`<E�`<Qa<:3a<eva<��a< 0b<��b<
�b<�>c<Thc<�hc<F<c<&�b<2hb<�a<3a<�`<�`<͞_<�U_<�6_<�B_<z_<��_<�W`<��`<��a<*b<�b<c<�\c<�oc<�Wc<c<�b<__b<�a<כa<IOa<�a<g�`<�`<��`<Qa<�Ga<��a<E�a<�Rb<$�b<c<VQc<�mc<L_c<w#c<:�b<#8b<e�a<��`<�d`<}�_<�_<�C_<�2_<9M_<��_<��_<<�`<�a< �a<	Ub<P�b<�0c<5bc<�fc<7Ac<A�b<c�b<�6b<��a<Vza<�4a<=a<��`<��`<��`<�a<uYa<&�a<
b<�pb<$�b<%c<Zc<)hc<<Jc<�b<1�b<��a<�^a<��`<�+`<˱_<�Z_<�+_<g(_<ZP_<�_<N`<��`<8Aa<S�a</ob<�b<1c<URc<SGc<�c<��b<Iab<?�a<�a<Ca<Na<�`<��`<Z�`<��`<�a<kNa<��a<xb<�mb<��b<ec<[>c<N>c<Ac<��b<�;b<�a<ta<�h`<��_<To_<�%_<%_<�_<�H_<��_<�%`<�`<�[a<��a<M�b<=�b<�)c<�<c<<$c<��b<��b<�*b<!�a<�fa<�a<�`<��`<˳`<��`<��`<#a<�]a<߹a< b<�  �  àb<�b<Rc<�c<`c<ֽb<�Jb<��a<Oa<EL`<r�_<�_<��^<�D^<�0^<:Q^<e�^<i#_<�_<�x`<�0a<�a<�mb<u�b<�c<�(c<c<i�b<1�b<�Rb<�b<Z�a<9�a<f�a<��a<.�a<N�a<��a<��a<��a<<b<�b<��b<�c<T3c<�5c<hc<ڷb<�8b<�a<��`<8/`<p�_<��^<��^<�[^<�Y^<y�^<��^<"|_<�%`<�`<��a<�9b<Ծb<Cc<�Jc<yNc<�-c<��b<�b<�bb<�!b<��a<��a<�a<$�a<��a<͵a<c�a<&�a<"-b<apb<-�b<��b<�5c<zOc<Cc<Y
c<<�b<�b<�oa<��`<�`<�`_<d�^<��^<�`^<�o^<$�^<7#_<��_<�h`<!a<}�a<Vmb<��b<�1c<UQc<~Gc<�c<O�b<��b<<Kb<�b<�a<{�a<�a<�a<��a<��a<G�a<Fb<�Bb<Q�b<#�b<�c<�Bc<cPc<�5c<��b<Vzb<��a<�2a<�z`<l�_<�/_<��^<�q^<�\^<�|^<.�^<pM_<G�_<�`<tXa<�b<��b<x�b<!;c<Lc<6c<�c<��b<�sb<l/b<��a<�a<��a<l�a<>�a<��a<��a<�a<Ab<	Ub<��b<��b<"c<.Fc<�Fc<�c<�b< Db<��a<��`<�3`<��_<�^<��^<jW^<nS^<˃^<�^<o_<�`<��`<�a<$b<k�b<�c<|/c<�1c<�c<��b<��b<�@b<g�a<a�a<��a<�a<��a<�a<m�a<��a<&�a<�b<�Gb<_�b<��b<4c<�%c<�c<l�b<�yb<��a<Ca<��`<��_<?2_<�^<�V^<�0^<�>^<�^<��^<�_<�6`<��`<�a<�:b<�b<��b<�c<�c<j�b<ʧb<�]b<b<��a<��a<߉a<Zxa<�ra<Twa<��a<��a<:�a<nb<]Vb<�  �  �b<X�b<��b<.�b<��b<~b<	 b<R[a<��`<��_<s_<-`^<`�]<�]<�r]<ԗ]<1�]<��^<\9_<�`<6�`<ׇa<�%b<�b<��b<� c< �b<��b<�b<{b<�Sb<s8b</)b<�"b< "b<�"b<T$b<8)b<�5b<�Lb<qb<+�b<��b<��b<8c<jc<��b<�tb<��a<O;a<w`<<�_<�^<9P^<X�]<��]<y�]<�]<�F^<��^<��_<Km`<:5a<��a<^zb<c�b<c<�*c<Dc<+�b<r�b<ܔb<�pb<Yb<`Lb<�Gb<eFb<;Fb<#Gb<�Lb<`[b<�ub<��b<��b<��b<bc<�(c<�c<�b<,^b<,�a<�a<�C`<?{_<+�^<�1^<��]<¢]<̳]<s�]<k^<`(_<�_<�`<fxa<!b< �b<6�b<�%c<�(c<�c<+�b<�b<ˆb<�fb<Sb<nIb<�Fb<Fb<RFb<uHb<Qb<$cb<��b<��b<��b<2c<@%c<�%c<# c<٭b<g/b<M�a<\�`<�_<T:_<��^<h^<s�]<��]<+�]<� ^<��^<qb_<�)`<��`<a�a<dKb<��b<�c<-$c<�c<:�b<��b<Q�b<�tb<�Xb<Ib<?Bb<�@b<�@b<�Ab<�Eb<,Qb<Ugb<#�b<�b<��b<yc<$c<�c<��b<ǁb<��a<hDa<~`<�_<��^<�P^<i�]<z�]<�]<d�]<�;^<��^<i�_<�[`<�!a<r�a<�bb<�b<��b<$c<��b<Z�b<I�b<{rb<.Mb<�4b< 'b<�!b<�b<6b<�b<=%b<Z3b<9Mb<osb<�b<��b<��b<�b<��b<7�b<�2b<!�a<;�`<�`<AM_<��^<k^</�]<�r]<%�]<m�]<N^<��^<2�_<]�`<Fa<a�a<qb<��b<
�b<��b<��b<��b<�|b<�Qb<%1b<pb<�b<�b<jb<�b<eb<ab<�.b<Nb<�xb<�  �  Φb<��b<l�b<n�b<�b<eBb<�a<�a<�B`<�j_<��^<��]<O]<��\<�\<�]<�k]<^<{�^<Y�_<v`<�<a<f�a< ab<s�b<��b<b�b<��b<�b<��b<;�b<6~b<��b<�b<��b<ܗb<m�b<S�b<�b<�b<��b<S�b<"�b<F�b<��b<��b<�b<#6b<��a<d�`<�`<zB_<{w^<��]<LM]<�	]<q]<;F]<��]<�j^<^5_<�`<�`<�a<�:b<��b<��b<hc<%�b<��b<M�b<�b<"�b<�b<��b<��b<R�b<T�b<²b<d�b<��b<��b<�b<��b<\�b< c<( c<��b<ޔb<�b<�za<�`<�_<�_< H^<e�]<v<]<;]<�]<r]<��]<в^<]�_<(\`<�)a<��a<zgb<i�b<��b<�c<��b<��b<�b<��b<�b<�b<�b<ݷb<��b<w�b<��b<-�b<��b<�b<3�b<N�b<��b<�c<0�b<-�b<,rb<E�a<�<a<kq`<ʘ_<W�^<3^<�{]<�"]<�]<�0]<�]<�0^<u�^<}�_<j�`<!ca<	b<��b<��b<V�b<4�b<�b<��b<ܳb<�b<��b<s�b<��b<u�b<�b<Ұb<קb<��b<l�b<�b<�b<d�b<��b<��b<��b<B�b<eCb<�a<��`<� `<BG_<z^<�]<_K]<�]< ]<�=]<�]<v]^<&_<-�_<��`<e�a<�#b<��b<t�b<��b<��b<��b<�b<��b<��b<��b<g�b<��b<��b<E�b<N�b<��b<�{b<c~b<��b<,�b<J�b<��b<Y�b<M�b<jb<b�a<Oa<}�`<ʹ_<��^<z^<Iy]<�]<�\<1�\<A]<F�]<=�^<�Q_<*`<u�`<Z�a<�4b<(�b<R�b<��b<M�b<1�b<�b<Uxb<Uob<Jqb<0yb<�b<҅b<��b<�zb<orb<�ob<mwb<�b<�  �  ��b< �b<��b<ƨb<�ub<�b<g�a<��`<�`<+'_<�L^<��]<��\<ї\<q}\<��\<�]<�]<�~^<�\_<�;`<�a<"�a<�7b<��b<��b<m�b<��b<��b<֝b<Ȝb<��b<T�b<Q�b<��b<~�b<��b<�b<´b<K�b<��b<ϭb<��b<X�b<��b<5�b<�vb<2
b<nqa<<�`<��_<?�^<�(^<�t]<�\<��\<�\<s�\< i]<�^<4�^<�_</�`<oa<�b<�b<f�b<x�b</�b<[�b<U�b<Q�b<��b<G�b<Z�b<t�b<�c<c<��b<��b<��b<��b<��b<�b<d�b<�b<��b<7�b<�kb<�a<�Ga<�~`<0�_<��^<��]<P]<��\<~�\<��\<�]<�]<�e^<�>_<p`<�`<�a<�<b<�b<��b<J�b<��b<v�b<��b<�b<|�b<��b<2�b<��b<_c<��b<��b<9�b<�b<0�b<C�b<7�b<�b<�b<��b<=�b<�Gb<��a<�a<�5`<QU_<`z^<P�]<�!]</�\<=�\<��\<e=]<��]<k�^<��_<	c`<a/a<��a<\b<��b<�b<8�b<��b<a�b<�b<��b<��b<D�b<��b<��b<��b<j�b<��b<M�b<��b<ѽb<��b<G�b<�b<��b<Z�b<�b<xb<�|a<]�`<��_<
_<J+^<�t]<�\<a�\<z�\<��\<4^]<�^<��^<�_<��`<�Ya<�a<�hb<B�b<��b<��b<y�b<�b<ޡb<?�b<ǯb<�b<n�b<1�b<�b<u�b<��b<��b<��b<i�b<I�b<U�b<��b<ڷb<��b<-Ab<��a<�a<�Q`<�s_<ה^<�]<� ]< �\<i}\<?�\<�\<�v]<^4^<+_<Y�_<��`<Eya<�	b<�lb<��b<L�b<��b<��b<w�b<��b<ӓb<֣b<D�b<��b<��b<0�b<��b<k�b<Еb<q�b<�b<�  �  ͷb<��b<��b<��b<��b<_Cb<�a<^�`<|�_<�K^<�]<\<�2[<R�Z<ʈZ<x�Z<;][<PB\<�]]</�^<��_<��`<��a<�gb<��b<��b<:�b<J�b<l�b<��b<k�b<S
c<>Hc<�c<�c<��c<?�c< gc<x*c<��b<��b<��b<�b<��b<V�b<�b<7�b<],b<�fa<�e`<<_<�^<��\<l�[<�[<,�Z<�Z<�[<��[<��\<b�]< '_<V`<_a<�-b<y�b<�c<�c<�c<g�b<��b<.�b<�c<�Fc<��c<)�c<��c<2�c<��c<(uc<�6c<c<��b<��b<��b<�c<�c<��b<��b<�b<)a<�`<6�^<y�]<�\<��[< [<1�Z<r�Z<&P[<�\<�)]<LZ^<M�_<a�`<�a<�eb<��b<hc<c<�c<��b<��b<C�b<sc<8Zc<ߖc<��c<��c<�c<ڜc<�`c<�$c<��b<#�b<=�b<� c<c<Bc<��b<�sb<��a<��`<��_<�z^<dG]<6\<_`[<m�Z<R�Z<X�Z<`�[<�l\<k�]<ƽ^<Q�_<N	a<��a<�b<)�b<>c<`c<��b<��b<��b<��b<�+c< ic<��c<�c<�c<��c<�c<bGc<]c<?�b<��b<��b<�c<ic<Dc<e�b<v:b<�ra<�o`<�C_<�^<��\<��[<�[<�Z<`�Z<�
[<��[<�\<r�]<�_<�A`<�Ha<cb<��b<��b<��b<��b<�b<�b<0�b<��b<� c<�]c<��c<��c<Ϊc<�c<ILc<�c<��b<{�b<��b<�b<��b<b�b<:�b<zsb<�a<��`<��_<t�^<~]<�]\<�q[<��Z<S�Z<"�Z<u[<��[<R�\<�'^<z`_<K�`<za<2b<Хb<��b<2�b<��b<ȸb<��b<��b<p�b<�"c<}_c<$�c<a�c<�c<=fc<�*c<�b<��b<��b<�  �  �b<�b<��b<R�b<�b<�[b<��a<��`<ȡ_<?m^<C>]<�0\<\^[<�Z<öZ<��Z<�[<%j\<l�]<�^<?�_<��`<&�a<#�b<��b<gc<r�b<H�b<�b<W�b<��b<��b<Q1c<=fc<��c<w�c<�{c<oMc<�c<U�b<��b<��b<f�b<R�b<�c<Cc<��b<Eb<�a<L�`<d[_<�&^<j ]<�\<SL[<�Z<��Z<_@[<��[<^�\<�^<�F_<�r`<aya<�Fb<U�b<fc<�-c<�c<uc<R�b<.�b<Ec<�4c<vkc<כc<n�c<��c<1�c<y]c<l&c<�b<|�b<��b<c<n c</*c<�c<��b<b<�Ca<$4`<�_<��]<��\<�[<?-[<%�Z<>[<(|[<�F\<UO]<S|^<�_<<�`<g�a<)~b<W�b<&c<9+c<�c<��b<�b<b�b<bc<�Ec<�{c<�c<;�c<5�c<&�c<>Kc<�c<��b<p�b<z�b<�c<�'c<�&c<��b<�b<��a<x�`<��_<�^<�l]<�^\<��[<)	[<R�Z<�[<<�[<��\<�]<��^<�`<c$a<b<E�b<Mc<#%c<�c<�c<\�b<9�b<G�b<�c<1Rc<��c<��c<�c<<�c<Pkc<m4c<c<V�b<��b<��b<-c<'c<mc<�b<*Sb<��a<�`<�b_<�+^<A]<m\<rJ[<��Z<<�Z<a7[<d�[<��\<��]<m4_<i^`<�ba<@.b<Ҷb<�b<�c<��b<�b<��b<2�b</�b<�c<�Dc<\tc<p�c<!�c<�hc<�4c<j�b<^�b<<�b<u�b<t�b<��b<��b<(�b<��b<D�a<�a<`<��^<�]<z�\<E�[<��Z<A�Z<��Z<qJ[<�\<]<�I^<_<%�`<�a<wJb<I�b<��b<T�b<M�b<��b<ϲb<��b<g�b<mc<zDc<�oc< �c<<sc<�Jc<(c<�b<��b<M�b<�  �  �b<c<)c<q0c<ac<s�b<z�a<�a<��_<
�^<^�]<��\<�[<6a[<q=[<,v[<�\<�\<��]<_<H;`<AIa<
&b<�b<Sc<	;c<�,c<c<�b<�b<��b<��b<��b<Cc<�)c<|/c<6c<��b<��b<��b<�b<��b<�b<�+c<3Ic<gCc<ic<�b<h�a<��`<`�_<��^<dn]<z}\<��[<(o[<9k[<��[<ll\<�Y]<Ds^<��_<�`<I�a<A�b<$c<Xc<ec<-Lc<�!c<��b<��b<�b<-�b<c<�@c<�Sc<�Pc<�8c<�c<��b<��b<��b<��b<)(c<vPc<cc<�Kc<]�b<ydb<�a<W�`<�__<�6^<i&]<�G\<�[<�n[<�[<��[< �\<ɺ]<^�^<�`<!a<�b<R�b<2c<�ac<k_c<>c<tc<��b<6�b<&�b<�c<$*c<�Hc<�Tc<�Jc<|-c<�	c<��b<��b<��b<~c<�7c<[c<�ac<<8c<��b<i$b<�;a<�%`<��^<��]<��\<�
\<m�[<j[<+�[<#0\<y]<�^<�:_<c`<$pa<Lb<O�b<�Ac<�^c<�Oc<�(c<b�b<��b<�b<��b<uc<�/c<�Ic<�Nc<�=c<ic<|�b<G�b<��b<��b<�c<pAc<<]c<�Uc<�c<.�b<U�a<p�`<׺_<�^<:q]<�}\<��[<�j[<�d[<��[<a\<�K]<Vc^<m�_<��`<Ьa<�sb<��b<�;c<�Fc<f,c<� c<,�b<�b< �b</�b<��b<:c<�+c<n(c<c<��b<��b<}�b<@�b<[�b<��b<�&c<�8c<!c<(�b<�8b<�ba<2Y`<�1_<T^<+�\<\<��[<�=[<zW[<*�[<�\<k�]<��^<�_<��`<`�a<��b<��b<-c<�*c<�c<��b<��b<��b<@�b<��b<��b<Bc<�c<�c<��b<��b<T�b<0�b<ɷb<�  �  M�b<�8c<�nc<y�c<�_c<��b<�Yb<%{a<�s`<sZ_<�I^<1Z]<&�\<�/\<6\<�B\<��\<d�]<�^<z�_<�`<�a<��b<
 c<)tc<�c<�nc<�4c<�b<ƴb<�b<�wb<~wb<��b<d�b<M�b<@�b<�~b<n{b<�b<l�b<�b<#c<�ec<�c<�c<�ac<��b<�2b<Ea<�5`<�_<O^<�7]<�\<�?\<Y<\<�\<l(]<�^<�	_<�#`<�7a<�,b<e�b<nc<��c<=�c<S�c<�Hc<�c<(�b<�b<��b<��b<��b<�b<{�b<ǧb<�b<1�b<$�b<��b<nc<lTc<��c<�c<�c<�Uc<U�b<��a<��`< �_<��^<��]<]<�|\<�@\<TX\<��\<�s]<u^^<�l_<��`<��a<�ub<M!c<�c<ٳc<a�c<�sc<�0c<��b<��b<j�b<�b<��b<�b<�b<ڮb<Z�b<��b<�b<t�b<#�b<�'c<Kkc<��c<۲c<|�c<.c<ŉb<��a<�`<d�_<dx^<p�]<��\<]\<�;\<o\<D�\<��]<ΰ^<Q�_<��`<��a<ïb<TEc<��c<ܭc<ّc<�Wc<Xc<��b<��b<�b<P�b<W�b<M�b<��b<ܦb<��b<9�b<Ţb<��b<�b<�:c<�{c<�c<6�c<�qc<��b<�>b<�Na<F=`<�"_<!^<+8]<�\<�;\<�5\<�\<]<�]<��^<�`<�#a<b<��b<�Sc<E�c<'�c<�hc<�'c<��b<E�b<��b<�xb<�zb<)�b<�b</�b<0b<Lub<9tb<�b<G�b<�b<�*c<�fc<��c<(wc<q*c<p�b<�a<H�`<&�_<I�^<t�]<~�\<CL\<�\<�&\<��\<yA]<,^<1:_<�S`<o^a<�Bb<��b<�Vc<|c<�qc<�>c<��b<��b<'�b<�lb<fb<�lb<�vb<|b<xb<�mb<�fb<�kb<Ʉb<&�b<�  �  �c<�ec<��c<��c<�c<�`c<��b<��a<�a<�`<m_<M:^<͗]<�4]<�]<�E]<'�]<�g^<�F_<A`<�@a<�.b<��b<a�c<��c<T�c<��c<\c<��b<q�b<)@b<��a<�a<�a<D�a<��a<P�a<��a<��a<�'b<vb<U�b<�=c<��c<[�c<��c<!�c<�Pc<��b<��a<��`<�_<�^<	 ^<��]<�G]<�D]<W�]<b^<]�^<i�_<ʿ`<�a</�b<�Tc<s�c<�d<�c<��c<wfc<� c<��b<LQb<�b<�a<	�a<��a<�a<��a<x�a<	 b<*^b<��b<.c<�xc<��c<��c<Q�c<7�c<Q1c<�qb<0�a<��`<��_<��^<��]<j~]<0J]<�^]<\�]<�V^<;'_<T`<4a<Kb<�b<��c<S�c<.d<�c<l�c<�Cc<��b<R�b<&:b<Xb<0�a<��a<��a<��a<��a<�b<�2b<Qxb<��b<7c<-�c<s�c<�d<��c<^�c<��b<�'b<�3a<�3`<+>_<�h^<��]<lb]<�E]<�q]<��]<��^<�p_<j`<�ha<�Ub<c<̦c<5�c<D�c<��c<�~c<$c<Y�b<�ab<� b<��a<k�a<�a<��a<��a<R�a<�b<�Cb<V�b<=�b<�Tc<M�c<G�c<�c<0�c<�^c<��b<��a<C�`<!�_<��^< ^<��]<fC]<9>]<\�]<^<��^<��_<��`<��a<ĉb<S<c<
�c<X�c<��c<ןc<HEc<\�b<�|b<e,b<��a<r�a<��a<ݱa<رa<r�a<��a<�a<5b<B�b<��b<�Nc<��c<z�c<y�c<Ҋc<Mc</Eb<�Za<�[`<�__<"}^<t�]<�M]<�]<-]<[�]<Z$^<��^<��_<C�`<&�a<��b<�Qc<a�c<��c<j�c<Tnc<:c<�b<
Lb<�b<��a<C�a<��a<¡a<�a<^�a<��a<��a<�Cb<�b<�  �  ��b<�yc<A�c<�d<�c<j�c<W%c<�jb<$�a<ϴ`<��_<�0_<��^<�Y^<�B^<kg^<��^<-W_<�`<9�`<��a<M�b<�Nc<D�c<Vd<�d<�c<�ic<q�b<kXb<O�a<:ba<}a<��`<Ǳ`<�`<��`<��`<�=a<�a<,$b<R�b<�=c<�c<�
d<)d<Pd<��c<�c<�Bb<ha<�`<�_<� _<Ĭ^<�o^<�m^<��^<�_<S�_<_�`<�\a<�:b<yc<��c<�d<�@d<g+d<��c<�ic<Y�b<�Sb<��a<Vja<Ja<�`<��`<�`<��`<^)a</}a<��a<eob<��b<�c<��c<�2d<;d<d<�c<�b<�b<�.a<�V`<p�_<C_<��^<=t^<�^<�^<�P_<w�_<]�`<^�a<��b<�Dc<I�c<?,d<�@d<�d<�c<8<c<�b<�%b<\�a<�Ka<Xa<v�`<;�`<^�`<a<?Ba<��a<6b<��b<�+c<��c<d<=d<�/d<��c<gUc<C�b<��a<��`<f`<j__<��^<h�^<p^<��^<[�^<2�_<�<`<sa<��a<��b<Muc<��c<4d<�2d<n�c<��c<�c<Wzb<��a<\�a<7,a<?�`<��`<3�`<_�`<ca<Za<��a<c>b<"�b<�Tc<��c<�d<�:d<Pd<��c<�c<�Lb<ooa<�`<��_<d!_<۪^<lk^<g^<��^<B_<��_<~p`<�Ja<�&b<�b<��c<U�c<�$d<pd<�c<�Hc<ݽb<)0b<��a<�Da<��`<��`<�`<�`<6�`<� a<ITa<��a<%Fb<�b<dYc<��c<Hd<d<}�c<�]c<8�b<"�a<C a<�'`<�h_<��^<�m^<�B^<S^<��^<z_<��_<��`<^ya<�Rb<�c<��c<[�c<Md</�c<�c<�c<�yb<x�a<�ua</a<��`<��`<��`<�`<�`<�a<�ja<��a<�jb<�  �  ��b<Ahc<��c<�d<d<p�c<jac<��b<jb<�Va<�`<�'`<��_<d�_<av_<��_<<�_<JE`<��`<��a<�9b<��b<L�c<�c<�)d<�d<��c<zRc<�b<v�a<�Da<�`<� `<�_<��_<υ_<��_<��_<�j`<@a<&�a<�hb<�c<��c<�d<�>d<A(d<��c<~Lc<T�b<Y�a<7=a<�`< $`<��_</�_<�_<D�_<s`<ߙ`<}5a<g�a<�b<�Lc<�c<�7d<�Wd<�5d<��c<�Hc<'�b<��a<&5a<U�`<$`<@�_<<�_<װ_<��_<�9`<��`<�Wa<�
b<��b<�hc<��c<�@d<�Td<a'd<O�c<�)c<�yb<��a<a<U�`<�`<(�_<��_<<�_<��_<L`<�`< ua<�)b<��b<u�c<�d<�Jd<�Sd<3d<t�c<�c<�]b<�a<��`<�n`<r`<��_<	�_<��_<��_<p``<��`<X�a<KHb<��b<��c<�d<�Nd<�Ld<�
d<��c<��b<�;b<	�a<&�`<]V`<`�_<V�_<ˣ_<r�_<L`<�p`<� a<)�a<bb<Vc<�c<�d<�Nd<Bd<P�c<buc<F�b<db<efa<��`<3A`<H�_<��_<ݤ_<
�_<"`<�`<�a<B�a<��b<�/c<:�c<�'d<�Pd<18d<��c<CXc<�b<��a<JBa<ǣ`<n$`<��_<�_<R�_<K�_<'`<G�`<�%a<S�a<΋b<�6c<��c<�d<�;d<d<	�c<�'c<�yb<6�a<qa<�v`<��_<#�_<��_<ň_<2�_</`<��`<�.a<C�a<~�b<�>c<d�c<d<�)d<��c<��c<��b</Lb<)�a<��`<fR`<"�_<�_<v_<<�_<8�_<u`<D�`<5Ba<��a<e�b<Pc<]�c<�d<�d<��c<�vc<��b<5(b<qa<w�`<k8`<��_<%�_<�q_<��_<��_<+`<Ѷ`<!^a<�b<�  �  Otb<^-c<ʵc<>d<�
d<��c<"tc<}�b<eb<�a<�ga<�a<��`<§`<>�`<<�`<�`<�a<T�a<x�a<Јb<
c<h�c<��c<d<��c<?�c<�c<,Rb<�xa<ԛ`<	�_<y#_<>�^<'_^<�R^<��^<8�^<)�_<�D`<�a<��a<��b<}yc<z�c<�%d<6d<H�c<�hc<�b<�Ub<��a<6ga<�a<D�`<��`<��`<��`<ma<5ea<\�a<�Sb<��b<Zlc<��c<u,d<@d<�d<M�c<� c<�4b<�Wa<t}`<[�_<7_<S�^<�y^<�^<��^<�8_<��_<�`<r�a<�ab<]&c<6�c<} d<�?d<ed<�c<`Pc<��b<t9b<ϼa<�Wa<�a<��`<`�`<t�`<��`<�4a<؍a<� b<��b<5c<3�c<d<�:d<k8d<��c<�rc<��b<��a<�a<7`<=~_<��^<2�^<Ft^<~�^<��^<�k_<D `<��`<��a<,�b<�_c<��c<�2d<�;d< d<P�c<i"c<��b<�b<��a<�:a<~�`<��`<��`<B�`<_a<Ka<�a<''b<��b<�=c<4�c<|d<;d<7#d<��c<�5c<�tb<��a<T�`<�_<D_<c�^<�~^<�q^<ş^<�_<��_<�_`<�8a<Sb<�b<�c<+d<�7d<+d<�c<Ytc<��b<]b<��a<�ia<a<W�`<��`<<�`<��`<$	a<�Wa<��a<�Ab<��b<Vc<n�c<5d<�#d<�c<ۅc<��b<�b<%4a<�X`<Γ_<��^<O�^<�Q^<�W^<��^<_<�_<	�`<1]a<8b<��b<�c<��c<cd<��c<��c<.#c<�b<�
b<]�a<�'a<9�`<n�`<��`<F�`<}�`<a<�Za<��a<gTb<��b<�ec<��c<�d<`d<,�c<>c<��b<%�a<9�`<,`<H_<��^<�^^<'>^<�X^<1�^<y6_<��_<��`<��a<�  �  b<��b<�fc<޼c<P�c<��c<�ac<��b<��b<�Ab<�a<"�a<��a<��a<C�a<�a<˺a<z�a<?b<]Wb<��b<c<6{c<��c<��c<i�c<�Tc<رb<d�a<��`<��_<��^<�'^<x�]<�8]<)]<Qb]<K�]<q�^<�~_<|`<�za<"db<�!c<l�c<��c<:�c<j�c<�_c<��b<q�b<�Hb<�b<��a<�a<v�a<O�a<,�a< �a<�b<�Kb<��b<* c<�fc<W�c<�c<% d<��c<:Oc<�b<A�a<ڸ`<]�_<X�^<R^<�]<NP]<X]<��]<d9^<�_<�_<�`<��a<t�b<Qmc<��c<Pd<��c<(�c<LRc<_�b<,�b<�Bb<b<�a<}�a<F�a<Q�a<��a<4�a<�(b<"kb<�b<�&c<ۉc<��c<fd<�c<�c<�c<�Ob<�`a<�a`<�h_<�^<��]<cr]<�I]<0j]<��]<�v^<	N_<xD`<Da<�5b<�c<��c<�c<(d<x�c<�c<�/c<e�b<Pqb<q,b<@�a<��a<�a<�a<Q�a<S�a<3b<8b<B�b<��b<oCc<.�c<��c<�c<��c<dxc<��b<��a<�a<``<�_<*H^<��]<X]<�G]<s�]<��]<��^<�_<�`<��a<${b<B7c<�c<��c<�c<3�c<�kc<^c<��b<�Mb<bb<X�a<�a<.�a<��a<6�a<��a<Nb<*<b<��b<��b<�Pc<�c<��c<�c<&�c<�/c<8xb<	�a<j�`<ؖ_<�^<�]<�i]<�(]<.0]<o]<�^<�^<�_<��`<m�a<��b<Cc<9�c<�c<��c<��c<�$c<?�b<G_b<�b<��a<�a<��a<K�a<��a<��a<]�a<��a<8b<�b<A�b<vVc<	�c<��c<�c<�rc<�b<�b<�+a<,`<%3_<�V^<��]<]<]<�]<�4]<��]<�A^<�_<�`<�a<�  �  7�a<rcb<>c<�bc<ׁc<�lc<$6c<�b<��b<+�b<�mb<4jb<+rb<�|b<��b<Q{b<]qb<�kb<�sb<�b<�b<[c<7Jc<!|c<�c<u\c< �b<�Ab<�[a<P`<�6_<�*^<WC]<��\<�1\<�\<�a\<��\<;�]<��^<��_<��`<��a<��b<�Dc<-�c< �c<�yc<O=c<2�b<��b<a�b<C�b<��b<9�b<V�b<�b<>�b<��b<W�b<��b<��b<�c<�Gc<݇c<m�c<t�c<�ic<%�b<{$b</a<_`<<_< ^<�(]<��\<pG\<�P\<��\<[R]<�4^<%>_<tW`<7fa<*Rb<�c<|c<(�c<��c<�{c<�9c<y�b<%�b<^�b<�b<?�b<Ūb<g�b<�b<�b<��b<��b<��b<%�b<�c<+ac<z�c<L�c<��c<�Dc<��b<��a<��`<t�_<��^<Ұ]<*�\<�n\<@\<ge\<0�\<ŗ]<��^<n�_<c�`<�a<��b<�5c<�c<��c<q�c<mfc<"c<��b<�b<3�b<y�b<�b<(�b<��b<��b<�b<��b<ݞb<�b<5�b<s.c<Uqc<M�c<3�c<�c<�c<eb<,~a<r`<oX_<�K^<�c]<õ\<JQ\<�>\<�\<�]<m�]<��^<��_<a<�b<��b<Xc<�c<�c<j�c<�Hc<�c<�b<b�b<��b<��b<G�b<�b<|�b<I�b<T�b<Ɇb<��b<ζb<z�b<V1c<�oc<D�c<y�c<5Lc<��b<�b<�a<�_<��^<��]<�]<�j\< \<�(\<Ã\<�)]<�^<$_<1.`<�<a<B(b<K�b<JQc<ăc<}c<�Nc<=c<2�b<�b<�tb<�jb<ob<yb<Db<f|b<Rrb<�ib<�kb<|�b<�b<�b<�-c<�fc<��c<hc<�c<Lwb<�a<��`<�_<r^<{]<R�\<�8\<R
\<�/\<�\< c]<uU^<�g_<,�`<�  �  �a<��a<L�b<�
c<N1c<;(c<�c<b�b<v�b<��b<i�b<�b<v�b<c<"c<�c<O�b<��b<_�b<��b<G�b<��b<7c<Y4c<v5c<+c<��b<E�a<z�`<`�_<|�^<�]<�\<��[<!b[<@N[<��[<�2\<�]<�)^<zT_<c{`<��a<MVb<��b<t8c<�Mc<|:c<bc<9�b<��b<��b<��b<�c<0+c<Cc<�Ec<M2c<�c<��b<�b<��b<�b<Mc<�Jc<wcc<yUc<�c<��b<��a<`�`<�_<tk^<�T]<l\<��[<v[<�[<n�[<�\<��]<��^<��_<��`<}�a<��b<8"c<�[c<k`c<�Bc<Dc<(�b<��b<��b<2�b<"c<�Bc<�Rc<�Lc<.2c<&c<k�b< �b<k�b<Kc<(1c<�Wc<�dc<�Dc<��b<�Gb<hha<Y`<�/_<L	^<C�\<A+\<v�[<n[<)�[<�\<4�\<N�]<�_<8`<HKa<�0b<��b<)<c<'bc<�Xc<4c<�c<m�b<]�b<�b<�c<�+c<�Gc<@Pc<nBc</#c<��b<��b<��b<��b<�c<q:c<�Zc<�Zc<�'c<r�b<f�a<a<]�_<��^<�]<l�\<��[<��[<�l[<~�[<P\<!2]<�D^<>n_<œ`<ٙa<�kb<�b< Jc<�]c<2Hc<�c<��b< �b<��b<��b<c<=)c<�>c<�>c<Y)c<�c<W�b<;�b<��b<��b<	c<k2c<XIc<�9c<��b<Efb<�a<I�`<�r_<G^<�/]<�E\<ՠ[<�N[<PX[<E�[<�p\<�d]<��^<��_<�`<��a<=}b<X�b<v0c<K4c<�c<��b<��b<��b<�b<��b<<�b<�c<� c<c<P�b<�b<B�b<�b<"�b<��b<��b<$c<1c<�c<��b<Eb<�3a<#$`<��^<��]<��\<��[<�k[<�8[<�a[<��[<��\< �]<@�^<�`<�  �  �`<��a<�bb<��b<��b<��b<��b<L�b<-�b<��b<��b<uc<�Pc<�xc<S�c<�rc<�Fc<c<0�b<N�b<I�b<��b<�b<��b<G�b<F�b<?Lb<��a<I�`<�y_<�D^<�]<\<cO[<e�Z<��Z<[<��[<�\<+�]<��^<�)`<58a<$b<3�b<��b<�c<c<(�b<h�b<�b<�b<�c<�Pc<b�c< �c<��c<Ќc<�\c<'c<��b<s�b<a�b<��b<_c<�+c<kc<��b<�?b<hpa<�h`<�<_<^<��\<��[<�D[<��Z<�Z<Uc[<!\<[ ]<�H^<z~_<��`<e�a<�bb<��b<$c<�*c<'c<��b<��b<�b<!	c<e:c<bqc<��c<�c<e�c<l�c<�Sc<&c<��b<��b<A�b<�c<�%c<�*c<c<q�b<t b<Za<�`<
�^<�]<��\<ܭ[<�[<O�Z<[<e�[<�o\<�]<��^<��_<��`<�a<P�b<�b<e'c<&c<�c<w�b<1�b<��b<3c<�Jc<%�c<��c<��c<u�c<�sc<?=c<s
c<��b<��b<�b<Qc<�%c<�c<��b<pb<ҵa<վ`<�_<Yf^<�:]<�5\<Xo[<��Z<^�Z<1[<��[<��\<$�]<�_<B`<Oa<\%b<��b<|c<7%c<�c<��b<��b<G�b<�b<\c<�Pc<n�c<��c<^�c<݃c<wQc<�c<�b<y�b<C�b<��b</c<�c<�b<�b<� b<�Oa<�F`<;_<��]<��\<��[<&[<I�Z<I�Z<2;[<��[<��\<�^<5U_<{`<qwa<m8b<�b<��b<��b<?�b<��b<��b<ȼb<�b<�	c<
@c<�mc<��c<�zc<}Uc<� c<��b<��b<O�b<�b<,�b<\�b<�b<>�b<fpb<%�a<��`<��_<�^<�k]<.V\<?x[<8�Z<ұZ<��Z<nd[<�:\<�K]<%|^<}�_<�  �  ��`<R�a<nJb<��b<1�b<��b<��b<l�b<G�b<��b<��b<91c<�lc<ݘc<��c<	�c<�ac<=%c<��b<��b<��b<r�b<�b<U�b<q�b<��b<�3b<�xa<O�`<*[_<�"^<�\<�[<8#[<��Z<��Z<��Z<X�[<�}\<O�]<��^<�`<�a<��a<(�b<�b<c<b�b<�b<��b<��b<%�b<�)c<�hc<��c<��c<��c<�c<vuc<�8c<�c<��b<}�b<l�b<c<�c<� c<��b<�&b<�Ua<�K`<�_<��]<��\<��[<�[<��Z<5�Z<�6[<��[<�\<,&^<[__<k�`<J�a<4Jb<U�b<	c<Ac<�c<��b<��b<p�b<�c<�Mc<h�c<��c<M�c<��c<�c<`jc<h-c<7�b<��b</�b<G�b<uc<�c<��b<5�b<��a<)a<��_<�^<S|]<�c\<Ђ[<K�Z<L�Z<j�Z<�m[<(G\<�Z]<c�^<i�_<�`<\�a<|b<��b<
c<`c< �b<��b<N�b<��b<�$c<�`c<-�c<��c<��c<��c<��c<nQc<c<��b<�b<��b<f c<�c<�c<[�b<�Wb<ޛa<ܢ`<)}_<!D^<]<�\<+C[<��Z<r�Z<�[<i�[<��\<E�]<��^<�$`<[4a<0b<��b<��b<�c<c<��b<@�b<��b<�b<X,c<�hc<	�c<{�c<W�c<�c<5jc<R+c<
�b<�b<a�b<=�b<��b<��b<��b<��b<�b<=5a<�)`<r�^<V�]<��\<��[<1�Z<h�Z<u�Z<�[<>�[<d�\<0�]<6_<�^`<T]a<�b<g�b<��b<�b<��b<��b<"�b<(�b<��b<c<	Zc<��c<�c<	�c<rc<@7c<.�b<��b<F�b<յb<��b<��b<�b<�b<-Xb<��a<��`<ڲ_<�|^<�F]<1.\<;M[<��Z<փZ<,�Z<9[<�\<�&]<�Z^<Z�_<�  �  �`<��a<�bb<��b<��b<��b<��b<L�b<-�b<��b<��b<uc<�Pc<�xc<S�c<�rc<�Fc<c<0�b<N�b<I�b<��b<�b<��b<G�b<F�b<?Lb<��a<I�`<�y_<�D^<�]<\<cO[<e�Z<��Z<[<��[<�\<+�]<��^<�)`<58a<$b<3�b<��b<�c<c<(�b<h�b<�b<�b<�c<�Pc<b�c< �c<��c<Ќc<�\c<'c<��b<s�b<a�b<��b<_c<�+c<kc<��b<�?b<hpa<�h`<�<_<^<��\<��[<�D[<��Z<�Z<Uc[<!\<[ ]<�H^<z~_<��`<e�a<�bb<��b<$c<�*c<'c<��b<��b<�b<!	c<e:c<bqc<��c<�c<e�c<l�c<�Sc<&c<��b<��b<A�b<�c<�%c<�*c<c<q�b<t b<Za<�`<
�^<�]<��\<ܭ[<�[<O�Z<[<e�[<�o\<�]<��^<��_<��`<�a<P�b<�b<e'c<&c<�c<w�b<1�b<��b<3c<�Jc<%�c<��c<��c<u�c<�sc<?=c<s
c<��b<��b<�b<Qc<�%c<�c<��b<pb<ҵa<վ`<�_<Yf^<�:]<�5\<Xo[<��Z<^�Z<1[<��[<��\<$�]<�_<B`<Oa<\%b<��b<|c<7%c<�c<��b<��b<G�b<�b<\c<�Pc<n�c<��c<^�c<݃c<wQc<�c<�b<y�b<C�b<��b</c<�c<�b<�b<� b<�Oa<�F`<;_<��]<��\<��[<&[<I�Z<I�Z<2;[<��[<��\<�^<5U_<{`<qwa<m8b<�b<��b<��b<?�b<��b<��b<ȼb<�b<�	c<
@c<�mc<��c<�zc<}Uc<� c<��b<��b<O�b<�b<,�b<\�b<�b<>�b<fpb<%�a<��`<��_<�^<�k]<.V\<?x[<8�Z<ұZ<��Z<nd[<�:\<�K]<%|^<}�_<�  �  �a<��a<L�b<�
c<N1c<;(c<�c<b�b<v�b<��b<i�b<�b<v�b<c<"c<�c<O�b<��b<_�b<��b<G�b<��b<7c<Y4c<v5c<+c<��b<E�a<z�`<`�_<|�^<�]<�\<��[<!b[<@N[<��[<�2\<�]<�)^<zT_<c{`<��a<MVb<��b<t8c<�Mc<|:c<bc<9�b<��b<��b<��b<�c<0+c<Cc<�Ec<M2c<�c<��b<�b<��b<�b<Mc<�Jc<wcc<yUc<�c<��b<��a<`�`<�_<tk^<�T]<l\<��[<v[<�[<n�[<�\<��]<��^<��_<��`<}�a<��b<8"c<�[c<k`c<�Bc<Dc<(�b<��b<��b<2�b<"c<�Bc<�Rc<�Lc<.2c<&c<k�b< �b<k�b<Kc<(1c<�Wc<�dc<�Dc<��b<�Gb<hha<Y`<�/_<L	^<C�\<A+\<v�[<n[<)�[<�\<4�\<N�]<�_<8`<HKa<�0b<��b<)<c<'bc<�Xc<4c<�c<m�b<]�b<�b<�c<�+c<�Gc<@Pc<nBc</#c<��b<��b<��b<��b<�c<q:c<�Zc<�Zc<�'c<r�b<f�a<a<]�_<��^<�]<l�\<��[<��[<�l[<~�[<P\<!2]<�D^<>n_<œ`<ٙa<�kb<�b< Jc<�]c<2Hc<�c<��b< �b<��b<��b<c<=)c<�>c<�>c<Y)c<�c<W�b<;�b<��b<��b<	c<k2c<XIc<�9c<��b<Efb<�a<I�`<�r_<G^<�/]<�E\<ՠ[<�N[<PX[<E�[<�p\<�d]<��^<��_<�`<��a<=}b<X�b<v0c<K4c<�c<��b<��b<��b<�b<��b<<�b<�c<� c<c<P�b<�b<B�b<�b<"�b<��b<��b<$c<1c<�c<��b<Eb<�3a<#$`<��^<��]<��\<��[<�k[<�8[<�a[<��[<��\< �]<@�^<�`<�  �  7�a<rcb<>c<�bc<ׁc<�lc<$6c<�b<��b<+�b<�mb<4jb<+rb<�|b<��b<Q{b<]qb<�kb<�sb<�b<�b<[c<7Jc<!|c<�c<u\c< �b<�Ab<�[a<P`<�6_<�*^<WC]<��\<�1\<�\<�a\<��\<;�]<��^<��_<��`<��a<��b<�Dc<-�c< �c<�yc<O=c<2�b<��b<a�b<C�b<��b<9�b<V�b<�b<>�b<��b<W�b<��b<��b<�c<�Gc<݇c<m�c<t�c<�ic<%�b<{$b</a<_`<<_< ^<�(]<��\<pG\<�P\<��\<[R]<�4^<%>_<tW`<7fa<*Rb<�c<|c<(�c<��c<�{c<�9c<y�b<%�b<^�b<�b<?�b<Ūb<g�b<�b<�b<��b<��b<��b<%�b<�c<+ac<z�c<L�c<��c<�Dc<��b<��a<��`<t�_<��^<Ұ]<*�\<�n\<@\<ge\<0�\<ŗ]<��^<n�_<c�`<�a<��b<�5c<�c<��c<q�c<mfc<"c<��b<�b<3�b<y�b<�b<(�b<��b<��b<�b<��b<ݞb<�b<5�b<s.c<Uqc<M�c<3�c<�c<�c<eb<,~a<r`<oX_<�K^<�c]<õ\<JQ\<�>\<�\<�]<m�]<��^<��_<a<�b<��b<Xc<�c<�c<j�c<�Hc<�c<�b<b�b<��b<��b<G�b<�b<|�b<I�b<T�b<Ɇb<��b<ζb<z�b<V1c<�oc<D�c<y�c<5Lc<��b<�b<�a<�_<��^<��]<�]<�j\< \<�(\<Ã\<�)]<�^<$_<1.`<�<a<B(b<K�b<JQc<ăc<}c<�Nc<=c<2�b<�b<�tb<�jb<ob<yb<Db<f|b<Rrb<�ib<�kb<|�b<�b<�b<�-c<�fc<��c<hc<�c<Lwb<�a<��`<�_<r^<{]<R�\<�8\<R
\<�/\<�\< c]<uU^<�g_<,�`<�  �  b<��b<�fc<޼c<P�c<��c<�ac<��b<��b<�Ab<�a<"�a<��a<��a<C�a<�a<˺a<z�a<?b<]Wb<��b<c<6{c<��c<��c<i�c<�Tc<رb<d�a<��`<��_<��^<�'^<x�]<�8]<)]<Qb]<K�]<q�^<�~_<|`<�za<"db<�!c<l�c<��c<:�c<j�c<�_c<��b<q�b<�Hb<�b<��a<�a<v�a<O�a<,�a< �a<�b<�Kb<��b<* c<�fc<W�c<�c<% d<��c<:Oc<�b<A�a<ڸ`<]�_<X�^<R^<�]<NP]<X]<��]<d9^<�_<�_<�`<��a<t�b<Qmc<��c<Pd<��c<(�c<LRc<_�b<,�b<�Bb<b<�a<}�a<F�a<Q�a<��a<4�a<�(b<"kb<�b<�&c<ۉc<��c<fd<�c<�c<�c<�Ob<�`a<�a`<�h_<�^<��]<cr]<�I]<0j]<��]<�v^<	N_<xD`<Da<�5b<�c<��c<�c<(d<x�c<�c<�/c<e�b<Pqb<q,b<@�a<��a<�a<�a<Q�a<S�a<3b<8b<B�b<��b<oCc<.�c<��c<�c<��c<dxc<��b<��a<�a<``<�_<*H^<��]<X]<�G]<s�]<��]<��^<�_<�`<��a<${b<B7c<�c<��c<�c<3�c<�kc<^c<��b<�Mb<bb<X�a<�a<.�a<��a<6�a<��a<Nb<*<b<��b<��b<�Pc<�c<��c<�c<&�c<�/c<8xb<	�a<j�`<ؖ_<�^<�]<�i]<�(]<.0]<o]<�^<�^<�_<��`<m�a<��b<Cc<9�c<�c<��c<��c<�$c<?�b<G_b<�b<��a<�a<��a<K�a<��a<��a<]�a<��a<8b<�b<A�b<vVc<	�c<��c<�c<�rc<�b<�b<�+a<,`<%3_<�V^<��]<]<]<�]<�4]<��]<�A^<�_<�`<�a<�  �  Otb<^-c<ʵc<>d<�
d<��c<"tc<}�b<eb<�a<�ga<�a<��`<§`<>�`<<�`<�`<�a<T�a<x�a<Јb<
c<h�c<��c<d<��c<?�c<�c<,Rb<�xa<ԛ`<	�_<y#_<>�^<'_^<�R^<��^<8�^<)�_<�D`<�a<��a<��b<}yc<z�c<�%d<6d<H�c<�hc<�b<�Ub<��a<6ga<�a<D�`<��`<��`<��`<ma<5ea<\�a<�Sb<��b<Zlc<��c<u,d<@d<�d<M�c<� c<�4b<�Wa<t}`<[�_<7_<S�^<�y^<�^<��^<�8_<��_<�`<r�a<�ab<]&c<6�c<} d<�?d<ed<�c<`Pc<��b<t9b<ϼa<�Wa<�a<��`<`�`<t�`<��`<�4a<؍a<� b<��b<5c<3�c<d<�:d<k8d<��c<�rc<��b<��a<�a<7`<=~_<��^<2�^<Ft^<~�^<��^<�k_<D `<��`<��a<,�b<�_c<��c<�2d<�;d< d<P�c<i"c<��b<�b<��a<�:a<~�`<��`<��`<B�`<_a<Ka<�a<''b<��b<�=c<4�c<|d<;d<7#d<��c<�5c<�tb<��a<T�`<�_<D_<c�^<�~^<�q^<ş^<�_<��_<�_`<�8a<Sb<�b<�c<+d<�7d<+d<�c<Ytc<��b<]b<��a<�ia<a<W�`<��`<<�`<��`<$	a<�Wa<��a<�Ab<��b<Vc<n�c<5d<�#d<�c<ۅc<��b<�b<%4a<�X`<Γ_<��^<O�^<�Q^<�W^<��^<_<�_<	�`<1]a<8b<��b<�c<��c<cd<��c<��c<.#c<�b<�
b<]�a<�'a<9�`<n�`<��`<F�`<}�`<a<�Za<��a<gTb<��b<�ec<��c<�d<`d<,�c<>c<��b<%�a<9�`<,`<H_<��^<�^^<'>^<�X^<1�^<y6_<��_<��`<��a<�  �  ��b<Ahc<��c<�d<d<p�c<jac<��b<jb<�Va<�`<�'`<��_<d�_<av_<��_<<�_<JE`<��`<��a<�9b<��b<L�c<�c<�)d<�d<��c<zRc<�b<v�a<�Da<�`<� `<�_<��_<υ_<��_<��_<�j`<@a<&�a<�hb<�c<��c<�d<�>d<A(d<��c<~Lc<T�b<Y�a<7=a<�`< $`<��_</�_<�_<D�_<s`<ߙ`<}5a<g�a<�b<�Lc<�c<�7d<�Wd<�5d<��c<�Hc<'�b<��a<&5a<U�`<$`<@�_<<�_<װ_<��_<�9`<��`<�Wa<�
b<��b<�hc<��c<�@d<�Td<a'd<O�c<�)c<�yb<��a<a<U�`<�`<(�_<��_<<�_<��_<L`<�`< ua<�)b<��b<u�c<�d<�Jd<�Sd<3d<t�c<�c<�]b<�a<��`<�n`<r`<��_<	�_<��_<��_<p``<��`<X�a<KHb<��b<��c<�d<�Nd<�Ld<�
d<��c<��b<�;b<	�a<&�`<]V`<`�_<V�_<ˣ_<r�_<L`<�p`<� a<)�a<bb<Vc<�c<�d<�Nd<Bd<P�c<buc<F�b<db<efa<��`<3A`<H�_<��_<ݤ_<
�_<"`<�`<�a<B�a<��b<�/c<:�c<�'d<�Pd<18d<��c<CXc<�b<��a<JBa<ǣ`<n$`<��_<�_<R�_<K�_<'`<G�`<�%a<S�a<΋b<�6c<��c<�d<�;d<d<	�c<�'c<�yb<6�a<qa<�v`<��_<#�_<��_<ň_<2�_</`<��`<�.a<C�a<~�b<�>c<d�c<d<�)d<��c<��c<��b</Lb<)�a<��`<fR`<"�_<�_<v_<<�_<8�_<u`<D�`<5Ba<��a<e�b<Pc<]�c<�d<�d<��c<�vc<��b<5(b<qa<w�`<k8`<��_<%�_<�q_<��_<��_<+`<Ѷ`<!^a<�b<�  �  ��b<�yc<A�c<�d<�c<j�c<W%c<�jb<$�a<ϴ`<��_<�0_<��^<�Y^<�B^<kg^<��^<-W_<�`<9�`<��a<M�b<�Nc<D�c<Vd<�d<�c<�ic<q�b<kXb<O�a<:ba<}a<��`<Ǳ`<�`<��`<��`<�=a<�a<,$b<R�b<�=c<�c<�
d<)d<Pd<��c<�c<�Bb<ha<�`<�_<� _<Ĭ^<�o^<�m^<��^<�_<S�_<_�`<�\a<�:b<yc<��c<�d<�@d<g+d<��c<�ic<Y�b<�Sb<��a<Vja<Ja<�`<��`<�`<��`<^)a</}a<��a<eob<��b<�c<��c<�2d<;d<d<�c<�b<�b<�.a<�V`<p�_<C_<��^<=t^<�^<�^<�P_<w�_<]�`<^�a<��b<�Dc<I�c<?,d<�@d<�d<�c<8<c<�b<�%b<\�a<�Ka<Xa<v�`<;�`<^�`<a<?Ba<��a<6b<��b<�+c<��c<d<=d<�/d<��c<gUc<C�b<��a<��`<f`<j__<��^<h�^<p^<��^<[�^<2�_<�<`<sa<��a<��b<Muc<��c<4d<�2d<n�c<��c<�c<Wzb<��a<\�a<7,a<?�`<��`<3�`<_�`<ca<Za<��a<c>b<"�b<�Tc<��c<�d<�:d<Pd<��c<�c<�Lb<ooa<�`<��_<d!_<۪^<lk^<g^<��^<B_<��_<~p`<�Ja<�&b<�b<��c<U�c<�$d<pd<�c<�Hc<ݽb<)0b<��a<�Da<��`<��`<�`<�`<6�`<� a<ITa<��a<%Fb<�b<dYc<��c<Hd<d<}�c<�]c<8�b<"�a<C a<�'`<�h_<��^<�m^<�B^<S^<��^<z_<��_<��`<^ya<�Rb<�c<��c<[�c<Md</�c<�c<�c<�yb<x�a<�ua</a<��`<��`<��`<�`<�`<�a<�ja<��a<�jb<�  �  �c<�ec<��c<��c<�c<�`c<��b<��a<�a<�`<m_<M:^<͗]<�4]<�]<�E]<'�]<�g^<�F_<A`<�@a<�.b<��b<a�c<��c<T�c<��c<\c<��b<q�b<)@b<��a<�a<�a<D�a<��a<P�a<��a<��a<�'b<vb<U�b<�=c<��c<[�c<��c<!�c<�Pc<��b<��a<��`<�_<�^<	 ^<��]<�G]<�D]<W�]<b^<]�^<i�_<ʿ`<�a</�b<�Tc<s�c<�d<�c<��c<wfc<� c<��b<LQb<�b<�a<	�a<��a<�a<��a<x�a<	 b<*^b<��b<.c<�xc<��c<��c<Q�c<7�c<Q1c<�qb<0�a<��`<��_<��^<��]<j~]<0J]<�^]<\�]<�V^<;'_<T`<4a<Kb<�b<��c<S�c<.d<�c<l�c<�Cc<��b<R�b<&:b<Xb<0�a<��a<��a<��a<��a<�b<�2b<Qxb<��b<7c<-�c<s�c<�d<��c<^�c<��b<�'b<�3a<�3`<+>_<�h^<��]<lb]<�E]<�q]<��]<��^<�p_<j`<�ha<�Ub<c<̦c<5�c<D�c<��c<�~c<$c<Y�b<�ab<� b<��a<k�a<�a<��a<��a<R�a<�b<�Cb<V�b<=�b<�Tc<M�c<G�c<�c<0�c<�^c<��b<��a<C�`<!�_<��^< ^<��]<fC]<9>]<\�]<^<��^<��_<��`<��a<ĉb<S<c<
�c<X�c<��c<ןc<HEc<\�b<�|b<e,b<��a<r�a<��a<ݱa<رa<r�a<��a<�a<5b<B�b<��b<�Nc<��c<z�c<y�c<Ҋc<Mc</Eb<�Za<�[`<�__<"}^<t�]<�M]<�]<-]<[�]<Z$^<��^<��_<C�`<&�a<��b<�Qc<a�c<��c<j�c<Tnc<:c<�b<
Lb<�b<��a<C�a<��a<¡a<�a<^�a<��a<��a<�Cb<�b<�  �  M�b<�8c<�nc<y�c<�_c<��b<�Yb<%{a<�s`<sZ_<�I^<1Z]<&�\<�/\<6\<�B\<��\<d�]<�^<z�_<�`<�a<��b<
 c<)tc<�c<�nc<�4c<�b<ƴb<�b<�wb<~wb<��b<d�b<M�b<@�b<�~b<n{b<�b<l�b<�b<#c<�ec<�c<�c<�ac<��b<�2b<Ea<�5`<�_<O^<�7]<�\<�?\<Y<\<�\<l(]<�^<�	_<�#`<�7a<�,b<e�b<nc<��c<=�c<S�c<�Hc<�c<(�b<�b<��b<��b<��b<�b<{�b<ǧb<�b<1�b<$�b<��b<nc<lTc<��c<�c<�c<�Uc<U�b<��a<��`< �_<��^<��]<]<�|\<�@\<TX\<��\<�s]<u^^<�l_<��`<��a<�ub<M!c<�c<ٳc<a�c<�sc<�0c<��b<��b<j�b<�b<��b<�b<�b<ڮb<Z�b<��b<�b<t�b<#�b<�'c<Kkc<��c<۲c<|�c<.c<ŉb<��a<�`<d�_<dx^<p�]<��\<]\<�;\<o\<D�\<��]<ΰ^<Q�_<��`<��a<ïb<TEc<��c<ܭc<ّc<�Wc<Xc<��b<��b<�b<P�b<W�b<M�b<��b<ܦb<��b<9�b<Ţb<��b<�b<�:c<�{c<�c<6�c<�qc<��b<�>b<�Na<F=`<�"_<!^<+8]<�\<�;\<�5\<�\<]<�]<��^<�`<�#a<b<��b<�Sc<E�c<'�c<�hc<�'c<��b<E�b<��b<�xb<�zb<)�b<�b</�b<0b<Lub<9tb<�b<G�b<�b<�*c<�fc<��c<(wc<q*c<p�b<�a<H�`<&�_<I�^<t�]<~�\<CL\<�\<�&\<��\<yA]<,^<1:_<�S`<o^a<�Bb<��b<�Vc<|c<�qc<�>c<��b<��b<'�b<�lb<fb<�lb<�vb<|b<xb<�mb<�fb<�kb<Ʉb<&�b<�  �  �b<c<)c<q0c<ac<s�b<z�a<�a<��_<
�^<^�]<��\<�[<6a[<q=[<,v[<�\<�\<��]<_<H;`<AIa<
&b<�b<Sc<	;c<�,c<c<�b<�b<��b<��b<��b<Cc<�)c<|/c<6c<��b<��b<��b<�b<��b<�b<�+c<3Ic<gCc<ic<�b<h�a<��`<`�_<��^<dn]<z}\<��[<(o[<9k[<��[<ll\<�Y]<Ds^<��_<�`<I�a<A�b<$c<Xc<ec<-Lc<�!c<��b<��b<�b<-�b<c<�@c<�Sc<�Pc<�8c<�c<��b<��b<��b<��b<)(c<vPc<cc<�Kc<]�b<ydb<�a<W�`<�__<�6^<i&]<�G\<�[<�n[<�[<��[< �\<ɺ]<^�^<�`<!a<�b<R�b<2c<�ac<k_c<>c<tc<��b<6�b<&�b<�c<$*c<�Hc<�Tc<�Jc<|-c<�	c<��b<��b<��b<~c<�7c<[c<�ac<<8c<��b<i$b<�;a<�%`<��^<��]<��\<�
\<m�[<j[<+�[<#0\<y]<�^<�:_<c`<$pa<Lb<O�b<�Ac<�^c<�Oc<�(c<b�b<��b<�b<��b<uc<�/c<�Ic<�Nc<�=c<ic<|�b<G�b<��b<��b<�c<pAc<<]c<�Uc<�c<.�b<U�a<p�`<׺_<�^<:q]<�}\<��[<�j[<�d[<��[<a\<�K]<Vc^<m�_<��`<Ьa<�sb<��b<�;c<�Fc<f,c<� c<,�b<�b< �b</�b<��b<:c<�+c<n(c<c<��b<��b<}�b<@�b<[�b<��b<�&c<�8c<!c<(�b<�8b<�ba<2Y`<�1_<T^<+�\<\<��[<�=[<zW[<*�[<�\<k�]<��^<�_<��`<`�a<��b<��b<-c<�*c<�c<��b<��b<��b<@�b<��b<��b<Bc<�c<�c<��b<��b<T�b<0�b<ɷb<�  �  �b<�b<��b<R�b<�b<�[b<��a<��`<ȡ_<?m^<C>]<�0\<\^[<�Z<öZ<��Z<�[<%j\<l�]<�^<?�_<��`<&�a<#�b<��b<gc<r�b<H�b<�b<W�b<��b<��b<Q1c<=fc<��c<w�c<�{c<oMc<�c<U�b<��b<��b<f�b<R�b<�c<Cc<��b<Eb<�a<L�`<d[_<�&^<j ]<�\<SL[<�Z<��Z<_@[<��[<^�\<�^<�F_<�r`<aya<�Fb<U�b<fc<�-c<�c<uc<R�b<.�b<Ec<�4c<vkc<כc<n�c<��c<1�c<y]c<l&c<�b<|�b<��b<c<n c</*c<�c<��b<b<�Ca<$4`<�_<��]<��\<�[<?-[<%�Z<>[<(|[<�F\<UO]<S|^<�_<<�`<g�a<)~b<W�b<&c<9+c<�c<��b<�b<b�b<bc<�Ec<�{c<�c<;�c<5�c<&�c<>Kc<�c<��b<p�b<z�b<�c<�'c<�&c<��b<�b<��a<x�`<��_<�^<�l]<�^\<��[<)	[<R�Z<�[<<�[<��\<�]<��^<�`<c$a<b<E�b<Mc<#%c<�c<�c<\�b<9�b<G�b<�c<1Rc<��c<��c<�c<<�c<Pkc<m4c<c<V�b<��b<��b<-c<'c<mc<�b<*Sb<��a<�`<�b_<�+^<A]<m\<rJ[<��Z<<�Z<a7[<d�[<��\<��]<m4_<i^`<�ba<@.b<Ҷb<�b<�c<��b<�b<��b<2�b</�b<�c<�Dc<\tc<p�c<!�c<�hc<�4c<j�b<^�b<<�b<u�b<t�b<��b<��b<(�b<��b<D�a<�a<`<��^<�]<z�\<E�[<��Z<A�Z<��Z<qJ[<�\<]<�I^<_<%�`<�a<wJb<I�b<��b<T�b<M�b<��b<ϲb<��b<g�b<mc<zDc<�oc< �c<<sc<�Jc<(c<�b<��b<M�b<�  �  CDb<tlb<��b<�b<}�b<�Yb<h�a<�h`<k�^< H]<�[<�Z<	�X<�5X< X<�TX<+Y<�mZ<_�[<*�]<�L_<��`<)�a<
b<��b<��b<-�b<�kb<lLb<�[b<U�b<c<|�c<7d<��d<Z�d<�gd<��c<rcc<��b<~b<Wb<fb<J�b<��b<O�b<o�b<q?b<VWa<6`<!�^<��\<�7[<"�Y<�X<b9X<�2X<��X<��Y<3[<j�\<gd^<��_<mJa<�?b<W�b<mc<��b<��b<ʉb<�wb<s�b<�b<*xc<*
d<H�d<>�d<O�d<�jd<��c<�Tc<��b<'�b<�rb<��b<��b<D�b<��b<��b<�b<�a<�_<^<�X\<{�Z<%yY<�X<3X<�YX<�Y<�'Z<p�[<#J]<[�^<u`<�a<|b<��b<�c<��b<ǧb<�|b<�yb<Y�b<�c<b�c<�5d<\�d<+�d<]�d<RCd<'�c<['c<��b<�{b<�xb<��b<��b<�b<��b<̊b<��a<�`<#_<jw]<7�[<JKZ<fY<dcX<\-X<A�X<�VY<��Z<n&\<?�]<�t_<��`<Z�a<a�b<w�b<�b<��b<Ǝb<ob<.~b<��b<#@c<]�c<�Xd<��d<$�d<��d<>d<�c<G�b<�b<�qb<	b<y�b<�b<��b<��b<qNb<da<�`<&�^<;�\<�:[<��Y<0�X<5X<+,X<B�X<0�Y<�[<ɣ\<jQ^<]�_<�2a<>&b<��b<��b<�b<W�b<�fb<Sb<�sb<@�b<jPc<��c<-Zd<��d<��d<�@d<۽c<�*c<Ǭb<4^b<�Hb<�cb<H�b<��b<
�b<D�b<��a<#�`<nv_<4�]<�)\<��Z<�HY<�dX<_X<�'X<�X< �Y<[n[<�]<��^<;A`<�ta<�Gb<յb<w�b<��b<fqb<�Eb<\Bb<Pwb<2�b<�nc<��c<Vfd<F�d<�nd<0d<�c<��b<��b<QFb<�  �  �[b<��b<��b<��b<��b<�b<6�a<��`<Z_<x]<��[<�UZ<�-Y<kvX<�AX<�X<�gY<E�Z<�/\<{�]<y_</�`<��a<:�b<Z�b<��b<��b<=�b<�ab<@fb<��b<+c<��c<�d<�dd<-ud<:@d<_�c<$Oc<a�b<B�b<�gb<��b<��b<��b<mc<��b<�hb<J�a<�<`<��^<
]<n[<Z<Y<�zX<�tX<��X<_�Y<�K[<S�\<��^<2$`<vta<^ib<��b<�,c<�c<��b<\�b<x�b<�b<��b<)ec<��c<�\d<&�d<��d<pEd<��c<�Dc<��b<f�b<҆b<��b<��b< c<p$c<��b<�9b<C0a<�_<u6^<ԋ\<F�Z<��Y< �X<�tX<ܚX<�DY<�aZ<��[<�z]<�!_<�`<��a<I�b<c<�+c<�c<��b<9�b<;�b<��b<c<\�c<d<�vd<ĝd<0~d<� d<ўc<^c<��b<��b<ߏb<�b<u�b<�'c<Pc<��b<��a<��`<L_<v�]<� \<��Z<J\Y<V�X<oX<��X<ޓY<M�Z<�Y\<�^<%�_<U	a<b<��b<�c<�c<[�b<@�b<M�b<��b<��b<=1c<u�c<=4d<ƅd<�d<a`d<��c<�mc<��b<B�b<m�b<��b<��b<�c<�&c<��b<�wb<�a<�F`<�^<�]</q[<�Z<HY<�vX<�mX<��X<��Y<�=[<��\<�^<�`<�\a<�Ob<��b<�c<F�b<>�b<k�b<eb<Uzb<�b<n=c<?�c<�3d<�od<�fd<}d<��c<�c<��b<sgb<�\b<|�b<o�b<��b<�b<��b<pb<za<��_<"^<�\\<k�Z< �Y<��X<�BX<�hX<bY<	/Z<}�[<KG]<�^<Al`<Ȟa<�pb<>�b<L�b<��b<C�b<K^b<�Pb<�yb<��b<�Wc<�c<�=d<�dd<�Ed<��c<Qgc<��b<��b<mSb<�  �  �b<�b<2c<ec<Zc<�b<�0b<�
a<S�_<^<�h\<��Z<��Y<2Y<��X<+OY<#Z<�H[<��\<�`^<�_<nXa<Skb<c<kc<�fc<�+c<N�b<��b<�b<��b<��b<gCc<5�c<A�c<�c<,�c<�tc<�c<>�b<\�b<&�b<w�b<�c<�ac<��c<]_c<��b<i�a<|�`<C4_<t�]<
\<��Z<n�Y<#8Y</2Y<b�Y<^�Z<��[<Du]<_<ϝ`<��a<��b<Dmc<<�c<��c<�>c<��b<�b<�b<��b<�)c<)�c<u�c<od<ld<��c<�uc<"c<��b<N�b<��b<<�b<�Jc<*�c<ޖc<�Rc< �b<B�a<\K`<��^<]<T�[<�dZ<��Y<�2Y<KWY<��Y<X	[<Go\<^<��_<�a<�Gb<Pc<c�c<��c<^nc<"c<��b<g�b<��b<�b<Ic<N�c<H�c<�d<>d<E�c<�Sc<9�b<R�b<�b<K�b<xc<�dc<�c<|�c<�'c<Xab<�:a<�_<�0^<̗\<|*[<
Z<%`Y<T-Y<�{Y<'DZ<�s[<��\<�^<K`<�a<��b<�Ac<��c<��c<Oc<Y c<��b<��b<3�b<�c<=ec<��c<vd<�d<E�c<�c<*.c<z�b<M�b<��b<W�b<�.c<wc<˗c<�pc<��b<b<ݿ`<C<_<�]<6\<C�Z<��Y<�3Y<[+Y<�Y<��Z<n�[<�d]<_<��`<P�a<��b<�Qc<��c<edc<6c<��b<��b<e�b<�b<c<�fc<m�c<��c<��c<��c< Lc<&�b<˛b<[~b<��b<'�b<� c<�_c<�kc<F'c<ׁb<cya<�`<�^<��\<_n[<�3Z<[^Y<Y<%Y<P�Y<m�Z<<\<��]<m_<��`<�b<��b<�Rc<Nfc<�8c<��b<��b<wb<�|b<³b<nc<zuc<l�c<>�c<��c<I�c<dc<��b<g�b<�ub<�  �  ��b<�[c<��c<+�c<��c<��c<�b<Ȱa<hN`<�^<�K]<��[<
�Z<)VZ<(Z<�pZ<)[<�@\<��]<x$_<r�`<S�a<�	c<ιc<1d<�c<k�c<:Nc<��b<E�b<s|b<)�b<h�b<(�b<c<!c<�c<_�b<��b<\�b<x�b<S�b<+c<��c<r�c<X d<��c<�zc<'�b<f_a<��_<�h^<�\<��[<��Z<�^Z<]YZ<��Z<�[<��\<UI^<��_<-Ia</�b<U{c<�
d<f:d<�d<��c<_Vc<[�b<%�b<#�b<Q�b<��b<�'c<8Fc<�Ac<�c<��b<�b<ʢb<��b<�c<�ic<}�c<�!d<�3d<��c<\Lc<dIb<-�`<�|_<9�]<��\<<s[<�Z<�ZZ<x|Z<�[<�
\<ZU]<��^<�V`<�a<>�b<�c<�$d<56d<��c<�c<�1c<��b<�b<�b<��b<�c<$4c<Hc<�7c<>
c<��b<z�b<��b<��b<%c<3�c<��c<%1d<�(d<��c<� c<��a<K~`<��^<�z]<�(\<�$[<^�Z<�UZ<ٝZ<FU[<2l\<��]<�M_<��`<�#b<E0c<`�c<�,d<9#d<��c<Qqc<H
c<��b<��b</�b<4�b<�c<:9c<�Ac<�&c<��b<Ҿb<��b<T�b<��b<�Cc<��c<�
d<�3d<d<��c<ңb<�ia<��_<=n^<7�\<%�[<��Z<fZZ<�RZ<6�Z<"�[<v�\<�8^<��_<�3a<�sb<�ac<(�c<�d<y�c<��c<�3c<�b<��b<{�b<��b<*�b<��b<�c<�c<��b<��b<*�b<�xb<��b<��b<e?c<)�c< �c<�d<�c< c<bb<e�`<bN_<��]<lc\<iB[<�~Z<�(Z<JZ<��Z<��[<"]<q�^<+#`<�a<+�b<��c<�c<d<6�c<�fc<��b<b�b<Xsb<�pb<m�b< �b<z�b<�c<��b<p�b<��b<�sb<�qb<ܜb<�  �  �>c<m�c<�Pd<әd<��d<2d<�qc<�^b<�a<q�_<!Z^<�1]<`P\<��[<�[<��[<�|\<�o]<�^<�`<�da<ͦb<�c<gWd<>�d<H�d<�Ad<J�c<�)c<ɣb<�?b<+b<��a<��a<�a<��a< �a<,�a<S�a<�'b<K{b<��b<X�c<@d<�d<s�d<W�d<d<�;c<�b<ʽ`<.\_<�^<� ]<2<\<��[<��[<�/\<@�\<��]<CA_<`�`<% b<1c<d<4�d<��d<ծd<�Ed<e�c<&c<_�b<(Rb<~#b<Mb<b<�$b<b#b<�b<"b<�&b<^b<ҽb<Ac<��c<�\d<�d<��d<M�d<(�c<i�b<��a<�W`<Y�^<7�]<v�\<8\<��[<�[<Vn\<G]<�h^<��_<4a<%ob<ˉc<�Td<�d<Z�d<6�d<�d<��c<h�b<m�b<
<b<�b<�b<�b<�$b<t b<�b<�b<}5b<>zb<��b<�rc<�d<>�d<��d<�d<ocd<E�c<3�b<�Ca<5�_<��^<�`]<@\<F�[<��[<\<"�\<��]<��^<h,`<(�a<j�b<��c<$}d<+�d<��d<�ed<q�c<�Lc<B�b<�ab<'&b<pb<Rb<b<�b<b<Gb<zb<�Db<
�b<�c<�c<80d<�d<��d<a�d<�'d<{Hc<Gb<��`<�a_<�^<�]<W:\<��[<��[<L&\<�\<��]<�0_<u�`<��a<�c<s d<��d<&�d<d�d<g$d<��c<�c<�b<�+b<�a<�a<>�a<��a<��a<��a<E�a<�a<4b<�b<
c<Z�c<M2d<_�d<��d<�bd<��c<9�b<��a<�(`<��^<ލ]<k�\<��[<Ѡ[<w�[<h;\<�]<M5^<$�_<��`<G;b<�Uc<u d<Y�d<I�d<�Zd<��c<�Mc<^�b<�Mb<!b<��a<K�a<Q�a<��a<s�a<W�a<��a<%�a<�Db<,�b<�  �  ?gc<�#d<��d<�
e<�e<�d<z�c<��b<��a<Z�`< r_<��^<n�]<c]<4E]<�t]<��]<O�^<��_<��`<�b<�1c<9$d<�d<e<De<[�d<!d< Gc<A�b<�a<[La<^�`<&�`<{�`<�`<��`<_�`<�"a<^�a<{:b<m�b<|�c<�sd<I�d<�.e<Qe<k�d<νc<��b<Ya<�O`<�=_<�`^<��]<�u]<�r]<�]<1R^<+_<�:`<ka<s�b<�c<.�d<4e<Ie<$e<�d<+�c<\0c<�pb<�a<Ra<a<��`<��`<��`<��`<Ja<�fa<��a<i�b<Xc<Wd<�d<|)e<�Ce<�e<ped<E{c<]b<)a<K�_<�^<�2^<��]<�w]<��]<��]<˛^<6�_<}�`<�a<(c<d<��d<�4e<�Be<��d<_kd<M�c<�b<�3b<e�a<<0a<��`<��`<v�`<�`<�`<\&a<m�a<4 b<p�b<#�c<�Vd<2�d<�<e<9e<��d<d<% c<��a<J�`<ء_<�^<��]<ȑ]<`s]<l�]<g^<3�^<��_<oa<�7b<�Yc<Kd<	�d<7=e<�,e<�d<\*d<�ic<��b<8�a<Lna<a<}�`<j�`<Y�`<_�`<X�`<�@a<D�a<Vb<�c<�c<׊d<Je<�Ae<He<8�d<^�c<�b<@�a</U`<�@_<$a^<�]<pq]<�k]<ĳ]<sF^<�_<1*`<"Xa<G�b<��c<�wd<��d<�+e<��d<ցd<��c<Mc<WKb<�a<�*a<��`<�`<��`<�`<��`<�`<�<a<��a<xkb<.c< �c<��d<��d<}e<��d<�8d<�Mc<�.b<�`<u�_<m�^<�^<�}]<�E]<�Z]<Ѽ]<oh^<�S_<�o`<S�a<@�b<
�c<��d<H e<�e<M�d<�5d<�{c<P�b<e�a<�ea<N�`<��`<h�`<w�`<S�`<ɯ`<��`<PXa<��a<ˠb<�  �  Tc<4d<{�d<X4e<�1e<��d<�)d<Hc<dLb<kSa<Nw`<��_<�L_<�_<��^<w_<�d_<s�_<I�`<m�a<�b<j�c<t[d<��d<aBe<�0e<P�d<�d<{)c<�,b<�7a<�b`<�_<�J_<�_<�_<E+_<��_<�`<��`<�a<��b<�c<5�d<9e<�Xe<8e<8�d<d<qc<�b<�&a<xY`<��_<�S_< _<�_<TO_<ٳ_<\N`<a<�	b<	c<;�c<D�d<0Fe<#se<�Be<7�d<��c<�c<�b<Ha<KO`<�_<\X_<l+_<n0_<�g_<g�_<�t`<�Da<�7b<%5c<� d<m�d<�Qe<<ne< .e<�d<^�c<)�b<n�a<g�`<M.`<T�_<J_<,&_<4_<�t_<��_<(�`<�ka<�bb<�_c<�Ed<j�d<1_e<Ile<ue<P~d<��c<[�b<1�a<��`<_`<2�_<RB_<�&_<�<_<|�_<�`<w�`<y�a<�b<c<gd<�e<3fe<Zce<�e<�Zd<�xc<�|b<��a<>�`<��_<|_<�5_<,"_<M@_<_<�`<��`<��a<G�b<��c<��d<�e<�ge<qUe<+�d<M4d<YLc<^Ob<�Ya<��`<��_<�k_<�._<�#_<�J_<w�_<�5`<��`<��a<��b<}�c<��d< 1e<�ke<�He<��d<�d<�c<yb<,a<�\`<N�_<�Q_<�_<�_<F_<�_<7@`<�a<��a<��b<��c<ͩd<�*e<�Ue<�#e<@�d<)�c<��b<��a<��`<(`<�_<�/_<a_<_<9>_<��_<�J`<�a<�b<c<s�c<ٲd<�&e<�Be<�e<6nd<��c<��b<$�a<L�`<m�_<�o_<�_<��^<_<UA_<q�_<y``<8a</b<�+c<�d<%�d<�*e<q7e<;�d<�Hd<�mc<�sb<4xa<��`<��_<iY_<�
_<��^<_<yN_<�_<�`<L^a<�Xb<�  �  ��b<��c<�d<
e<�e<��d<#d<�]c<�b<�a<=Ta<e�`<�`<\�`<	�`<��`<�`<a<Ssa<�b<^�b<��c<�Fd<
�d<�e<ye<5�d<��c<��b<�a<�k`<@R_<�j^<��]<gf]<�U]<��]<�^<��^<��_<la<cRb<�oc<�Wd<��d<s.e<Be<�d<��c<M:c<�xb<��a<�Oa<9�`<�`<�`<B�`<6�`<u�`<�La<��a<�rb<�4c<��c<ŧd<�e<�He<ze<7�d<Ϋc<R�b<�aa<�3`<"(_<�S^<��]<�~]<�]<�]<c{^<�\_<�q`<��a<��b<�c<X�d<@'e<wDe<�e<8�d<8�c<S
c<�Mb<b�a<D=a<��`<��`<<�`<��`<��`<�a<�ya<0b<͵b<�zc<j:d<��d<46e<�Ae<��d<�Ed<Qc<�,b<~�`<�_<^�^<�^<Ϣ]<�w]<	�]<�^<y�^<�_<��`<�	b<S1c<�,d<j�d<�;e<:e<��d<�Kd<c�c<��b<mb<e�a<Ya<��`<��`<ѹ`<��`<O�`<�/a<�a<7b<��b<�c<Ond<e�d<>e<"+e<.�d<E�c<��b<��a<Ս`<t_<B�^<��]<�]<v]<s�]<0:^<;_<�`<�8a<Mlb<@�c<Qnd<ce<OAe<!e<��d<�d<wDc<Ȁb<N�a<�Ra<��`<*�`<��`<o�`<�`<��`<�>a<j�a<�_b<�c<F�c<]�d<�e<�+e<M�d<Yid<d�c<�pb<�<a<�`<_<,^<f�]<�U]<�]]<��]<�Q^<�2_<�G`<�xa<��b<��c<��d<$�d<�e<g�d<,Wd<]�c<��b<db<�a<a<��`</�`<O�`<��`</�`<��`<�Ea<I�a<ہb<�Fc<Sd<f�d<�e<(e<��d<ld<0c<��a<��`<�_<
�^<z�]<Pk]<W@]<�b]<��]<A�^<N~_<ɠ`<��a<�  �  dnb<�}c<�9d<�d<͗d<oKd<��c<�7c<+�b<Bb<H�a<O�a<Y�a<��a<��a<��a<a�a<=�a<hb<�Yb<��b<�]c<��c<�hd<�d<��d<�!d<�Rc<5b<��`<	�_<�0^<[]<@\<�[<��[<] \<Ү\<�]<@�^<�N`<E�a<u�b<�c<@}d<��d<p�d<�Ad<�c<c&c<h�b<hHb< b<�b<zb<�b<�b<Ub<b<�b<Lb<
�b<	'c<Q�c< Id< �d<D�d<?�d<ud<�&c<��a<Q�`<B7_<�]<.�\<x4\<�[<��[<7T\<f]<�4^<��_<��`<�8b<^c<q7d<l�d<��d<<�d<#+d<��c<.
c</�b<Cb<tb<�b<\b<�"b<U b<�b<Tb<c-b<�kb<��b<�Zc<��c<Ard<��d<��d<�|d<��c<`�b<T�a<�`<��^<ő]<Y�\<
\<7�[<��[<��\</s]<Ǟ^<z�_<�Xa<աb<q�c<ld<��d<0�d<�|d<w�c<�hc<��b<�rb<�/b<~b<Fb<�b< b<0b<b<b<A9b<��b<��b<��c<Gd<?�d<��d<V�d<�Ed</vc<	Xb<^a<1�_<uR^<�4]<a\<��[<��[<�\<_�\<��]<�
_<	j`<�a<� c<��c<��d<|�d<,�d<[Pd<P�c<�0c<1�b<�Mb<b<8b<�	b<Zb<�b<b<X b<�b<�;b<@�b<�c<�c<�/d<��d<��d<'�d<��c<;c<F�a<]s`<9_<��]<u�\<#\<C�[<��[<�*\<��\<�
^<-W_<��`<�b<�3c<�d<2�d<æd<�pd<��c<�lc<?�b<dcb<yb<�a<��a<��a<��a<��a<6�a<i�a<e�a<�7b<��b<�&c<��c<>d<s�d<D�d<�Gd<��c<��b<:Ja<C�_<.�^<�Z]<)l\<��[< �[<��[<W\<7=]<bi^<��_<�$a<�  �  1�a<S�b<�c<��c<z�c<��c<�Vc<�b<7�b<sb<xb<��b<�b<bc<�c<N�b<G�b<z�b<1vb<}{b<��b<(c<�tc<]�c<hd<9�c<Ѓc<��b<׃a<�`<&�^<]<�[<��Z<�SZ<�9Z<��Z<�`[<φ\<��]<^v_<X�`<f@b<�?c<��c<�d<�	d<�c<Pc<�b<٨b<5�b<F�b<K�b<�c<�3c<7c<�c<�b<Ĳb<�b<�b<��b<�Vc<��c<cd<�9d<�d<psc<�b<�;a<��_<�<^<��\<��[<�Z<$dZ<qZ<$�Z<��[<T]<��^<;`<��a<�b<>�c<*d<�6d<�	d<<�c<@c<R�b<\�b<%�b<��b<G�b<�+c<�Ec<y;c<�c<��b<e�b<��b<��b<pc<�}c<��c<1,d<�1d<��c<;*c<�b<��`<<>_<�]<:`\<�M[<ڛZ<�YZ<��Z<�4[<W=\<O�]<�_<G�`<��a<c<H�c<�+d<�.d<��c<��c<�c<��b<��b<��b<�b<2	c<-5c<4Cc<-c<9�b<��b<J�b<��b<x�b< 1c<��c<�c<01d<(d< �c<5�b<٦a<`<`<M�^<�<]<~�[<�[<VtZ<�YZ<ܵZ<[<I�\<�^<x�_<a<�Xb<-Vc<h�c<�1d<hd<x�c<w\c<)�b<��b<��b<@�b<��b<�c<X/c<>0c<�c<R�b<��b<|�b<%�b<��b<�?c<��c<�c<ld<��c<�Rc<�]b<�a<��_<	^<%�\<"z[<ȤZ<p;Z<HZ<��Z<s�[<��\<�e^<H�_<W[a<��b<gnc<��c<�
d<��c<�~c<�c<0�b<Z}b<Ksb<��b<��b<��b<7c<�c<�b<��b<Gzb<�pb<z�b<Z�b<{Ic<\�c<��c<*�c<��c<�b<T�a<��`<�_<y�]<j)\<�[<�dZ<�"Z<XZ<[�Z<�\<]]<^�^<Sa`<�  �  �a<^=b<d�b<�\c<�cc<�.c<��b<\�b<3wb<�b<��b<R%c<�c<��c<r�c<��c<�uc<�c<��b<��b<gb<ͬb<o�b<�Dc<^pc<�Xc<,�b<�b<��`<�b_<�]<�3\<X�Z<g�Y<Z.Y<)Y<wY<VSZ<C�[<]<M�^<�E`<ԝa<��b<Bc<-�c<�rc<�2c<��b<�b<��b<Y�b<gc<Ikc<H�c<+d<�	d<��c<}c<c<]�b<��b<�b<I�b<�>c<��c<3�c<ic<��b<��a<X�`<�_<Xg]<_�[<ؖZ<�Y<�<Y<�JY<��Y<`�Z<�/\<ٿ]<�\_<R�`<�b<��b<�yc<U�c<�vc<-c<��b<��b<{�b<^�b<�5c<�c<��c<�d<�	d<+�c<#dc<�c<��b<v�b<{�b<�
c<�Yc<+�c<`�c<�@c<}�b<Xta<.`<y^<h�\<xf[<u;Z<RyY<f1Y<�jY< Z<i@[<��\<#J^<
�_<Oa<pb<�0c<@�c<�c<�_c<�c<=�b<�b<��b<��b<�Uc<T�c<�d<�d<��c<��c<�=c<��b<�b<��b<��b<X c<�kc<D�c<�}c<o
c<^3b<	�`<D�_<4�]<`U\<��Z<U�Y<�NY<2Y<0�Y<�qZ<��[<_3]<Q�^<#_`<�a<�b<�Vc<Ӕc<c�c<Ac<�b<��b<R�b<��b<\c<�kc<^�c<� d<�d<��c<eqc<�
c<�b<�b<�b<�b<�%c<Ric<�c<Jc<�b<Իa<�k`<��^<~A]<��[<PoZ<ˆY<Y<�!Y<_�Y<�Z<+\<�]<3_<#�`<,�a<��b<HNc<Noc<�Ic<z�b<S�b<��b<P}b<X�b<0c<�ic<�c<e�c<�c<�c<�/c<��b<ȉb<Nub<]�b<��b<d%c<�^c<�_c<>c<qVb<�>a<k�_<�B^< �\<�/[<�Z<�BY<��X<�4Y<��Y<�
[<�{\<�^<3�_<�  �  �`<��a<j�b<w�b<��b<	�b<<�b<c[b<�Vb<6�b<!�b<rc<��c<3Md<
id<�>d<��c<�Uc<j�b<�|b<VWb<hb<�b<��b< c<J�b<rb<�a<d`<"�^<�;]<#�[<*Z<�Y<�qX<$TX<�X<+�Y<�Z<��\<�1^<��_<(a<D-b<Y�b<�c<<c<0�b<[�b<psb<��b<*�b<�:c<��c<=;d<Ӄd<�d<�Id<��c<lRc<N�b<��b<��b<g�b< �b<�c<\+c<U�b<,ab<nha<K`<��^<��\<�@[<�Y<��X<�~X<��X<�!Y<�,Z<��[<83]<N�^<�c`<��a<��b<9c<�*c<Gc<��b<N�b<��b<|�b<��b<fwc<i�c<hd<`�d<��d<p2d<��c<N/c<}�b<��b<��b<��b<:�b<�$c<~!c<	�b<�b<��`<��_<�]<�H\< �Z<��Y<��X<sX<�X<�mY<c�Z<|\<��]<�d_<�`<[�a<��b<.c<&c<2�b<>�b<P�b<q�b<�b<�c<��c<#d<J}d<��d<�md<�d<0�c<�c<��b<��b< �b<��b<�c<&c<a
c<h�b<��a<�`<�_<^]<߻[<gKZ<�4Y<�X<�sX<3�X<w�Y<q[<��\<�L^<J�_<@a<�Cb<��b<�"c<�c<��b<��b<w}b<\�b<��b<�=c<H�c<Q9d<td<@�d<�@d<H�c<ZDc<��b<ہb<�mb<A�b<��b<��b<6c<g�b<�@b<PFa<��_<�]^<��\<[<��Y<��X<7VX<�dX<��X<"Z<�j[<u	]<[�^<�9`<'za<�\b<��b<s�b<v�b<�b<�jb<%Ub<6tb<��b<{Ec<��c<�4d<�fd<�Rd<F�c<U�c<�b<>�b<�Xb<oWb<��b<�b<��b<�b<[�b<��a<�`<�[_<�]<~\<|�Z<�SY<�X<�<X<2yX<�7Y<�eZ<��[<k�]<�0_<�  �  'z`<�a<Dab<�b<+�b<��b<�jb<�Db<Jb<݈b<��b<
�c<�d<�vd<\�d<�fd<��c<lc<F�b<�yb<UHb<Ob<�|b<7�b<#�b<�b<�Hb<qa<�8`<��^<2]<�d[<��Y<Q�X<|0X<�X<;~X<iY<��Z<S\<9^<Ξ_<��`<�b<�b<��b<��b<X�b<Axb<�_b<yb<#�b<�Kc<~�c<�`d<��d<�d<5pd<��c<�dc<��b<L�b<pb<J�b<�b<��b<c< �b<�7b<Q>a<��_<:T^<b�\<�	[<i�Y<c�X<9=X<0LX<��X<��Y<�^[<]<��^<}8`<�za<J^b<��b<�c<��b<Ϯb<`b<Utb<�b<'c<k�c<rd<��d<��d<��d<hVd<��c<y=c<��b<��b<�ub<Зb<9�b<��b<�b<ۣb<�a</�`<e_<~�]<	\<e�Z<_MY<~X<c1X<�nX<40Y<>bZ<3�[<�]<�7_<O�`<��a<b�b<��b<��b<��b<��b<�ub<{b<��b<�+c<��c<*Fd<��d<�d<�d<)d<��c<�c<�b<�rb<Bxb<��b<1�b<"�b<��b<.mb<��a< \`<N�^<U-]<n�[<@Z<3�X<�PX<\2X<U�X<R�Y<��Z<Po\<,^<Z�_<�a<b<��b<(�b<�b<ѻb<��b<�ib<b<|�b<�Nc<�c<�^d<6�d<>�d<�fd<!�c<�Vc<K�b<�zb<[b<&ob<��b<S�b<��b<�b<b<6a<%�_<�/^<�\<�Z<�Y<M�X<�X<A#X<��X<l�Y<�4[<D�\<��^<I`<=Pa<V3b<c�b<g�b<��b<(�b<�Pb<�Db<�ob<��b<wZc<��c<r\d<��d<�|d<6"d<��c<+	c<W�b<_Mb<�Ab<�cb<�b<T�b<��b<2ob<+�a<�`<b/_<��]<��[<�SZ<�Y<wGX<��W<m8X<K�X<�,Z<E�[<�]]<�_<�  �  �`<��a<j�b<w�b<��b<	�b<<�b<c[b<�Vb<6�b<!�b<rc<��c<3Md<
id<�>d<��c<�Uc<j�b<�|b<VWb<hb<�b<��b< c<J�b<rb<�a<d`<"�^<�;]<#�[<*Z<�Y<�qX<$TX<�X<+�Y<�Z<��\<�1^<��_<(a<D-b<Y�b<�c<<c<0�b<[�b<psb<��b<*�b<�:c<��c<=;d<Ӄd<�d<�Id<��c<lRc<N�b<��b<��b<g�b< �b<�c<\+c<U�b<,ab<nha<K`<��^<��\<�@[<�Y<��X<�~X<��X<�!Y<�,Z<��[<83]<N�^<�c`<��a<��b<9c<�*c<Gc<��b<N�b<��b<|�b<��b<fwc<i�c<hd<`�d<��d<p2d<��c<N/c<}�b<��b<��b<��b<:�b<�$c<~!c<	�b<�b<��`<��_<�]<�H\< �Z<��Y<��X<sX<�X<�mY<c�Z<|\<��]<�d_<�`<[�a<��b<.c<&c<2�b<>�b<P�b<q�b<�b<�c<��c<#d<J}d<��d<�md<�d<0�c<�c<��b<��b< �b<��b<�c<&c<a
c<h�b<��a<�`<�_<^]<߻[<gKZ<�4Y<�X<�sX<3�X<w�Y<q[<��\<�L^<J�_<@a<�Cb<��b<�"c<�c<��b<��b<w}b<\�b<��b<�=c<H�c<Q9d<td<@�d<�@d<H�c<ZDc<��b<ہb<�mb<A�b<��b<��b<6c<g�b<�@b<PFa<��_<�]^<��\<[<��Y<��X<7VX<�dX<��X<"Z<�j[<u	]<[�^<�9`<'za<�\b<��b<s�b<v�b<�b<�jb<%Ub<6tb<��b<{Ec<��c<�4d<�fd<�Rd<F�c<U�c<�b<>�b<�Xb<oWb<��b<�b<��b<�b<[�b<��a<�`<�[_<�]<~\<|�Z<�SY<�X<�<X<2yX<�7Y<�eZ<��[<k�]<�0_<�  �  �a<^=b<d�b<�\c<�cc<�.c<��b<\�b<3wb<�b<��b<R%c<�c<��c<r�c<��c<�uc<�c<��b<��b<gb<ͬb<o�b<�Dc<^pc<�Xc<,�b<�b<��`<�b_<�]<�3\<X�Z<g�Y<Z.Y<)Y<wY<VSZ<C�[<]<M�^<�E`<ԝa<��b<Bc<-�c<�rc<�2c<��b<�b<��b<Y�b<gc<Ikc<H�c<+d<�	d<��c<}c<c<]�b<��b<�b<I�b<�>c<��c<3�c<ic<��b<��a<X�`<�_<Xg]<_�[<ؖZ<�Y<�<Y<�JY<��Y<`�Z<�/\<ٿ]<�\_<R�`<�b<��b<�yc<U�c<�vc<-c<��b<��b<{�b<^�b<�5c<�c<��c<�d<�	d<+�c<#dc<�c<��b<v�b<{�b<�
c<�Yc<+�c<`�c<�@c<}�b<Xta<.`<y^<h�\<xf[<u;Z<RyY<f1Y<�jY< Z<i@[<��\<#J^<
�_<Oa<pb<�0c<@�c<�c<�_c<�c<=�b<�b<��b<��b<�Uc<T�c<�d<�d<��c<��c<�=c<��b<�b<��b<��b<X c<�kc<D�c<�}c<o
c<^3b<	�`<D�_<4�]<`U\<��Z<U�Y<�NY<2Y<0�Y<�qZ<��[<_3]<Q�^<#_`<�a<�b<�Vc<Ӕc<c�c<Ac<�b<��b<R�b<��b<\c<�kc<^�c<� d<�d<��c<eqc<�
c<�b<�b<�b<�b<�%c<Ric<�c<Jc<�b<Իa<�k`<��^<~A]<��[<PoZ<ˆY<Y<�!Y<_�Y<�Z<+\<�]<3_<#�`<,�a<��b<HNc<Noc<�Ic<z�b<S�b<��b<P}b<X�b<0c<�ic<�c<e�c<�c<�c<�/c<��b<ȉb<Nub<]�b<��b<d%c<�^c<�_c<>c<qVb<�>a<k�_<�B^< �\<�/[<�Z<�BY<��X<�4Y<��Y<�
[<�{\<�^<3�_<�  �  1�a<S�b<�c<��c<z�c<��c<�Vc<�b<7�b<sb<xb<��b<�b<bc<�c<N�b<G�b<z�b<1vb<}{b<��b<(c<�tc<]�c<hd<9�c<Ѓc<��b<׃a<�`<&�^<]<�[<��Z<�SZ<�9Z<��Z<�`[<φ\<��]<^v_<X�`<f@b<�?c<��c<�d<�	d<�c<Pc<�b<٨b<5�b<F�b<K�b<�c<�3c<7c<�c<�b<Ĳb<�b<�b<��b<�Vc<��c<cd<�9d<�d<psc<�b<�;a<��_<�<^<��\<��[<�Z<$dZ<qZ<$�Z<��[<T]<��^<;`<��a<�b<>�c<*d<�6d<�	d<<�c<@c<R�b<\�b<%�b<��b<G�b<�+c<�Ec<y;c<�c<��b<e�b<��b<��b<pc<�}c<��c<1,d<�1d<��c<;*c<�b<��`<<>_<�]<:`\<�M[<ڛZ<�YZ<��Z<�4[<W=\<O�]<�_<G�`<��a<c<H�c<�+d<�.d<��c<��c<�c<��b<��b<��b<�b<2	c<-5c<4Cc<-c<9�b<��b<J�b<��b<x�b< 1c<��c<�c<01d<(d< �c<5�b<٦a<`<`<M�^<�<]<~�[<�[<VtZ<�YZ<ܵZ<[<I�\<�^<x�_<a<�Xb<-Vc<h�c<�1d<hd<x�c<w\c<)�b<��b<��b<@�b<��b<�c<X/c<>0c<�c<R�b<��b<|�b<%�b<��b<�?c<��c<�c<ld<��c<�Rc<�]b<�a<��_<	^<%�\<"z[<ȤZ<p;Z<HZ<��Z<s�[<��\<�e^<H�_<W[a<��b<gnc<��c<�
d<��c<�~c<�c<0�b<Z}b<Ksb<��b<��b<��b<7c<�c<�b<��b<Gzb<�pb<z�b<Z�b<{Ic<\�c<��c<*�c<��c<�b<T�a<��`<�_<y�]<j)\<�[<�dZ<�"Z<XZ<[�Z<�\<]]<^�^<Sa`<�  �  dnb<�}c<�9d<�d<͗d<oKd<��c<�7c<+�b<Bb<H�a<O�a<Y�a<��a<��a<��a<a�a<=�a<hb<�Yb<��b<�]c<��c<�hd<�d<��d<�!d<�Rc<5b<��`<	�_<�0^<[]<@\<�[<��[<] \<Ү\<�]<@�^<�N`<E�a<u�b<�c<@}d<��d<p�d<�Ad<�c<c&c<h�b<hHb< b<�b<zb<�b<�b<Ub<b<�b<Lb<
�b<	'c<Q�c< Id< �d<D�d<?�d<ud<�&c<��a<Q�`<B7_<�]<.�\<x4\<�[<��[<7T\<f]<�4^<��_<��`<�8b<^c<q7d<l�d<��d<<�d<#+d<��c<.
c</�b<Cb<tb<�b<\b<�"b<U b<�b<Tb<c-b<�kb<��b<�Zc<��c<Ard<��d<��d<�|d<��c<`�b<T�a<�`<��^<ő]<Y�\<
\<7�[<��[<��\</s]<Ǟ^<z�_<�Xa<աb<q�c<ld<��d<0�d<�|d<w�c<�hc<��b<�rb<�/b<~b<Fb<�b< b<0b<b<b<A9b<��b<��b<��c<Gd<?�d<��d<V�d<�Ed</vc<	Xb<^a<1�_<uR^<�4]<a\<��[<��[<�\<_�\<��]<�
_<	j`<�a<� c<��c<��d<|�d<,�d<[Pd<P�c<�0c<1�b<�Mb<b<8b<�	b<Zb<�b<b<X b<�b<�;b<@�b<�c<�c<�/d<��d<��d<'�d<��c<;c<F�a<]s`<9_<��]<u�\<#\<C�[<��[<�*\<��\<�
^<-W_<��`<�b<�3c<�d<2�d<æd<�pd<��c<�lc<?�b<dcb<yb<�a<��a<��a<��a<��a<6�a<i�a<e�a<�7b<��b<�&c<��c<>d<s�d<D�d<�Gd<��c<��b<:Ja<C�_<.�^<�Z]<)l\<��[< �[<��[<W\<7=]<bi^<��_<�$a<�  �  ��b<��c<�d<
e<�e<��d<#d<�]c<�b<�a<=Ta<e�`<�`<\�`<	�`<��`<�`<a<Ssa<�b<^�b<��c<�Fd<
�d<�e<ye<5�d<��c<��b<�a<�k`<@R_<�j^<��]<gf]<�U]<��]<�^<��^<��_<la<cRb<�oc<�Wd<��d<s.e<Be<�d<��c<M:c<�xb<��a<�Oa<9�`<�`<�`<B�`<6�`<u�`<�La<��a<�rb<�4c<��c<ŧd<�e<�He<ze<7�d<Ϋc<R�b<�aa<�3`<"(_<�S^<��]<�~]<�]<�]<c{^<�\_<�q`<��a<��b<�c<X�d<@'e<wDe<�e<8�d<8�c<S
c<�Mb<b�a<D=a<��`<��`<<�`<��`<��`<�a<�ya<0b<͵b<�zc<j:d<��d<46e<�Ae<��d<�Ed<Qc<�,b<~�`<�_<^�^<�^<Ϣ]<�w]<	�]<�^<y�^<�_<��`<�	b<S1c<�,d<j�d<�;e<:e<��d<�Kd<c�c<��b<mb<e�a<Ya<��`<��`<ѹ`<��`<O�`<�/a<�a<7b<��b<�c<Ond<e�d<>e<"+e<.�d<E�c<��b<��a<Ս`<t_<B�^<��]<�]<v]<s�]<0:^<;_<�`<�8a<Mlb<@�c<Qnd<ce<OAe<!e<��d<�d<wDc<Ȁb<N�a<�Ra<��`<*�`<��`<o�`<�`<��`<�>a<j�a<�_b<�c<F�c<]�d<�e<�+e<M�d<Yid<d�c<�pb<�<a<�`<_<,^<f�]<�U]<�]]<��]<�Q^<�2_<�G`<�xa<��b<��c<��d<$�d<�e<g�d<,Wd<]�c<��b<db<�a<a<��`</�`<O�`<��`</�`<��`<�Ea<I�a<ہb<�Fc<Sd<f�d<�e<(e<��d<ld<0c<��a<��`<�_<
�^<z�]<Pk]<W@]<�b]<��]<A�^<N~_<ɠ`<��a<�  �  Tc<4d<{�d<X4e<�1e<��d<�)d<Hc<dLb<kSa<Nw`<��_<�L_<�_<��^<w_<�d_<s�_<I�`<m�a<�b<j�c<t[d<��d<aBe<�0e<P�d<�d<{)c<�,b<�7a<�b`<�_<�J_<�_<�_<E+_<��_<�`<��`<�a<��b<�c<5�d<9e<�Xe<8e<8�d<d<qc<�b<�&a<xY`<��_<�S_< _<�_<TO_<ٳ_<\N`<a<�	b<	c<;�c<D�d<0Fe<#se<�Be<7�d<��c<�c<�b<Ha<KO`<�_<\X_<l+_<n0_<�g_<g�_<�t`<�Da<�7b<%5c<� d<m�d<�Qe<<ne< .e<�d<^�c<)�b<n�a<g�`<M.`<T�_<J_<,&_<4_<�t_<��_<(�`<�ka<�bb<�_c<�Ed<j�d<1_e<Ile<ue<P~d<��c<[�b<1�a<��`<_`<2�_<RB_<�&_<�<_<|�_<�`<w�`<y�a<�b<c<gd<�e<3fe<Zce<�e<�Zd<�xc<�|b<��a<>�`<��_<|_<�5_<,"_<M@_<_<�`<��`<��a<G�b<��c<��d<�e<�ge<qUe<+�d<M4d<YLc<^Ob<�Ya<��`<��_<�k_<�._<�#_<�J_<w�_<�5`<��`<��a<��b<}�c<��d< 1e<�ke<�He<��d<�d<�c<yb<,a<�\`<N�_<�Q_<�_<�_<F_<�_<7@`<�a<��a<��b<��c<ͩd<�*e<�Ue<�#e<@�d<)�c<��b<��a<��`<(`<�_<�/_<a_<_<9>_<��_<�J`<�a<�b<c<s�c<ٲd<�&e<�Be<�e<6nd<��c<��b<$�a<L�`<m�_<�o_<�_<��^<_<UA_<q�_<y``<8a</b<�+c<�d<%�d<�*e<q7e<;�d<�Hd<�mc<�sb<4xa<��`<��_<iY_<�
_<��^<_<yN_<�_<�`<L^a<�Xb<�  �  ?gc<�#d<��d<�
e<�e<�d<z�c<��b<��a<Z�`< r_<��^<n�]<c]<4E]<�t]<��]<O�^<��_<��`<�b<�1c<9$d<�d<e<De<[�d<!d< Gc<A�b<�a<[La<^�`<&�`<{�`<�`<��`<_�`<�"a<^�a<{:b<m�b<|�c<�sd<I�d<�.e<Qe<k�d<νc<��b<Ya<�O`<�=_<�`^<��]<�u]<�r]<�]<1R^<+_<�:`<ka<s�b<�c<.�d<4e<Ie<$e<�d<+�c<\0c<�pb<�a<Ra<a<��`<��`<��`<��`<Ja<�fa<��a<i�b<Xc<Wd<�d<|)e<�Ce<�e<ped<E{c<]b<)a<K�_<�^<�2^<��]<�w]<��]<��]<˛^<6�_<}�`<�a<(c<d<��d<�4e<�Be<��d<_kd<M�c<�b<�3b<e�a<<0a<��`<��`<v�`<�`<�`<\&a<m�a<4 b<p�b<#�c<�Vd<2�d<�<e<9e<��d<d<% c<��a<J�`<ء_<�^<��]<ȑ]<`s]<l�]<g^<3�^<��_<oa<�7b<�Yc<Kd<	�d<7=e<�,e<�d<\*d<�ic<��b<8�a<Lna<a<}�`<j�`<Y�`<_�`<X�`<�@a<D�a<Vb<�c<�c<׊d<Je<�Ae<He<8�d<^�c<�b<@�a</U`<�@_<$a^<�]<pq]<�k]<ĳ]<sF^<�_<1*`<"Xa<G�b<��c<�wd<��d<�+e<��d<ցd<��c<Mc<WKb<�a<�*a<��`<�`<��`<�`<��`<�`<�<a<��a<xkb<.c< �c<��d<��d<}e<��d<�8d<�Mc<�.b<�`<u�_<m�^<�^<�}]<�E]<�Z]<Ѽ]<oh^<�S_<�o`<S�a<@�b<
�c<��d<H e<�e<M�d<�5d<�{c<P�b<e�a<�ea<N�`<��`<h�`<w�`<S�`<ɯ`<��`<PXa<��a<ˠb<�  �  �>c<m�c<�Pd<әd<��d<2d<�qc<�^b<�a<q�_<!Z^<�1]<`P\<��[<�[<��[<�|\<�o]<�^<�`<�da<ͦb<�c<gWd<>�d<H�d<�Ad<J�c<�)c<ɣb<�?b<+b<��a<��a<�a<��a< �a<,�a<S�a<�'b<K{b<��b<X�c<@d<�d<s�d<W�d<d<�;c<�b<ʽ`<.\_<�^<� ]<2<\<��[<��[<�/\<@�\<��]<CA_<`�`<% b<1c<d<4�d<��d<ծd<�Ed<e�c<&c<_�b<(Rb<~#b<Mb<b<�$b<b#b<�b<"b<�&b<^b<ҽb<Ac<��c<�\d<�d<��d<M�d<(�c<i�b<��a<�W`<Y�^<7�]<v�\<8\<��[<�[<Vn\<G]<�h^<��_<4a<%ob<ˉc<�Td<�d<Z�d<6�d<�d<��c<h�b<m�b<
<b<�b<�b<�b<�$b<t b<�b<�b<}5b<>zb<��b<�rc<�d<>�d<��d<�d<ocd<E�c<3�b<�Ca<5�_<��^<�`]<@\<F�[<��[<\<"�\<��]<��^<h,`<(�a<j�b<��c<$}d<+�d<��d<�ed<q�c<�Lc<B�b<�ab<'&b<pb<Rb<b<�b<b<Gb<zb<�Db<
�b<�c<�c<80d<�d<��d<a�d<�'d<{Hc<Gb<��`<�a_<�^<�]<W:\<��[<��[<L&\<�\<��]<�0_<u�`<��a<�c<s d<��d<&�d<d�d<g$d<��c<�c<�b<�+b<�a<�a<>�a<��a<��a<��a<E�a<�a<4b<�b<
c<Z�c<M2d<_�d<��d<�bd<��c<9�b<��a<�(`<��^<ލ]<k�\<��[<Ѡ[<w�[<h;\<�]<M5^<$�_<��`<G;b<�Uc<u d<Y�d<I�d<�Zd<��c<�Mc<^�b<�Mb<!b<��a<K�a<Q�a<��a<s�a<W�a<��a<%�a<�Db<,�b<�  �  ��b<�[c<��c<+�c<��c<��c<�b<Ȱa<hN`<�^<�K]<��[<
�Z<)VZ<(Z<�pZ<)[<�@\<��]<x$_<r�`<S�a<�	c<ιc<1d<�c<k�c<:Nc<��b<E�b<s|b<)�b<h�b<(�b<c<!c<�c<_�b<��b<\�b<x�b<S�b<+c<��c<r�c<X d<��c<�zc<'�b<f_a<��_<�h^<�\<��[<��Z<�^Z<]YZ<��Z<�[<��\<UI^<��_<-Ia</�b<U{c<�
d<f:d<�d<��c<_Vc<[�b<%�b<#�b<Q�b<��b<�'c<8Fc<�Ac<�c<��b<�b<ʢb<��b<�c<�ic<}�c<�!d<�3d<��c<\Lc<dIb<-�`<�|_<9�]<��\<<s[<�Z<�ZZ<x|Z<�[<�
\<ZU]<��^<�V`<�a<>�b<�c<�$d<56d<��c<�c<�1c<��b<�b<�b<��b<�c<$4c<Hc<�7c<>
c<��b<z�b<��b<��b<%c<3�c<��c<%1d<�(d<��c<� c<��a<K~`<��^<�z]<�(\<�$[<^�Z<�UZ<ٝZ<FU[<2l\<��]<�M_<��`<�#b<E0c<`�c<�,d<9#d<��c<Qqc<H
c<��b<��b</�b<4�b<�c<:9c<�Ac<�&c<��b<Ҿb<��b<T�b<��b<�Cc<��c<�
d<�3d<d<��c<ңb<�ia<��_<=n^<7�\<%�[<��Z<fZZ<�RZ<6�Z<"�[<v�\<�8^<��_<�3a<�sb<�ac<(�c<�d<y�c<��c<�3c<�b<��b<{�b<��b<*�b<��b<�c<�c<��b<��b<*�b<�xb<��b<��b<e?c<)�c< �c<�d<�c< c<bb<e�`<bN_<��]<lc\<iB[<�~Z<�(Z<JZ<��Z<��[<"]<q�^<+#`<�a<+�b<��c<�c<d<6�c<�fc<��b<b�b<Xsb<�pb<m�b< �b<z�b<�c<��b<p�b<��b<�sb<�qb<ܜb<�  �  �b<�b<2c<ec<Zc<�b<�0b<�
a<S�_<^<�h\<��Z<��Y<2Y<��X<+OY<#Z<�H[<��\<�`^<�_<nXa<Skb<c<kc<�fc<�+c<N�b<��b<�b<��b<��b<gCc<5�c<A�c<�c<,�c<�tc<�c<>�b<\�b<&�b<w�b<�c<�ac<��c<]_c<��b<i�a<|�`<C4_<t�]<
\<��Z<n�Y<#8Y</2Y<b�Y<^�Z<��[<Du]<_<ϝ`<��a<��b<Dmc<<�c<��c<�>c<��b<�b<�b<��b<�)c<)�c<u�c<od<ld<��c<�uc<"c<��b<N�b<��b<<�b<�Jc<*�c<ޖc<�Rc< �b<B�a<\K`<��^<]<T�[<�dZ<��Y<�2Y<KWY<��Y<X	[<Go\<^<��_<�a<�Gb<Pc<c�c<��c<^nc<"c<��b<g�b<��b<�b<Ic<N�c<H�c<�d<>d<E�c<�Sc<9�b<R�b<�b<K�b<xc<�dc<�c<|�c<�'c<Xab<�:a<�_<�0^<̗\<|*[<
Z<%`Y<T-Y<�{Y<'DZ<�s[<��\<�^<K`<�a<��b<�Ac<��c<��c<Oc<Y c<��b<��b<3�b<�c<=ec<��c<vd<�d<E�c<�c<*.c<z�b<M�b<��b<W�b<�.c<wc<˗c<�pc<��b<b<ݿ`<C<_<�]<6\<C�Z<��Y<�3Y<[+Y<�Y<��Z<n�[<�d]<_<��`<P�a<��b<�Qc<��c<edc<6c<��b<��b<e�b<�b<c<�fc<m�c<��c<��c<��c< Lc<&�b<˛b<[~b<��b<'�b<� c<�_c<�kc<F'c<ׁb<cya<�`<�^<��\<_n[<�3Z<[^Y<Y<%Y<P�Y<m�Z<<\<��]<m_<��`<�b<��b<�Rc<Nfc<�8c<��b<��b<wb<�|b<³b<nc<zuc<l�c<>�c<��c<I�c<dc<��b<g�b<�ub<�  �  �[b<��b<��b<��b<��b<�b<6�a<��`<Z_<x]<��[<�UZ<�-Y<kvX<�AX<�X<�gY<E�Z<�/\<{�]<y_</�`<��a<:�b<Z�b<��b<��b<=�b<�ab<@fb<��b<+c<��c<�d<�dd<-ud<:@d<_�c<$Oc<a�b<B�b<�gb<��b<��b<��b<mc<��b<�hb<J�a<�<`<��^<
]<n[<Z<Y<�zX<�tX<��X<_�Y<�K[<S�\<��^<2$`<vta<^ib<��b<�,c<�c<��b<\�b<x�b<�b<��b<)ec<��c<�\d<&�d<��d<pEd<��c<�Dc<��b<f�b<҆b<��b<��b< c<p$c<��b<�9b<C0a<�_<u6^<ԋ\<F�Z<��Y< �X<�tX<ܚX<�DY<�aZ<��[<�z]<�!_<�`<��a<I�b<c<�+c<�c<��b<9�b<;�b<��b<c<\�c<d<�vd<ĝd<0~d<� d<ўc<^c<��b<��b<ߏb<�b<u�b<�'c<Pc<��b<��a<��`<L_<v�]<� \<��Z<J\Y<V�X<oX<��X<ޓY<M�Z<�Y\<�^<%�_<U	a<b<��b<�c<�c<[�b<@�b<M�b<��b<��b<=1c<u�c<=4d<ƅd<�d<a`d<��c<�mc<��b<B�b<m�b<��b<��b<�c<�&c<��b<�wb<�a<�F`<�^<�]</q[<�Z<HY<�vX<�mX<��X<��Y<�=[<��\<�^<�`<�\a<�Ob<��b<�c<F�b<>�b<k�b<eb<Uzb<�b<n=c<?�c<�3d<�od<�fd<}d<��c<�c<��b<sgb<�\b<|�b<o�b<��b<�b<��b<pb<za<��_<"^<�\\<k�Z< �Y<��X<�BX<�hX<bY<	/Z<}�[<KG]<�^<Al`<Ȟa<�pb<>�b<L�b<��b<C�b<K^b<�Pb<�yb<��b<�Wc<�c<�=d<�dd<�Ed<��c<Qgc<��b<��b<mSb<�  �  �`<�`<)Ya<��a<�b<��a<�(a<�_<<�]<��[<��Y<{yW<�U<N�T<�wT<��T<Q"V<��W<�Z<�R\<�o^<@.`<�fa<�b<�b<��a<�Ca<��`<6�`<��`<lla<db<�wc<=id<Ue<x e<Ǽd<��c<1�b<'�a<sa<*�`<��`<*a<��a<�b<~7b<��a<~�`<�__<yh]<1[<�X< W<��U<�T<:�T<�kU<��V<�X<��Z<X:]<>_<#�`<��a<�Lb<�9b<+�a<�Ea<M�`<l�`<!a<3�a<A�b<��c<w�d<�Ce<�4e<̧d<޽c<��b<��a<��`<�`<-�`<�\a<O�a<~Ab<=;b<l�a<�`<��^<Ѿ\<�~Z<=SX<?~V<q:U<��T<��T<8�U<4vW<��Y<a�[<��]<��_<�=a<Sb<LRb<�b<�a<�a<��`<
�`<�Ta<q5b<_Fc<�Id<Je<�Le<Ee<Pbd<Ddc<sQb<0ha<��`<(�`<ca<��a<#b<�Nb<�b<�Ya<�`<z*^<� \<b�Y<��W<?�U<��T<��T<�U<�NV<UX<y;Z<M|\<
�^<�U`</�a<j.b<�Bb<��a<�ga<�`<C�`<��`<a�a<�b<ݚc<�d<�$e<�Be<��d<�d<Yc</�a<(+a<Z�`<�`<�0a<;�a<7*b<�Ib<��a<�`<�j_<q]<(7[<��X<� W<��U<�T<1�T<�aU<K�V<.�X<��Z<}&]<�'_<z�`<��a<�/b<vb<��a<�"a<��`<-�`<��`<|�a<��b<9�c<��d<�e<?	e<o|d<��c<vb<��a<:�`<p�`<ý`</2a<��a<gb<�b<&~a<V`<ܤ^<�\<=OZ<�"X<�LV<U<zT<�T<ߧU<�BW<�OY<Z�[<��]<=�_<�a<<�a<�b<��a<Pga<��`<��`<-�`<Ca<W�a<�c<�d<h�d<e<��d<v(d<"+c<.b<�0a<��`<�  �  �`<�a<=�a<z#b<�bb<T-b<�ga<A`<�:^<F\<�Y<��W<�(V<�!U<��T<=MU<{V<G<X<�ZZ<w�\<U�^<Yl`<<�a<|Kb<�db<�b<��a<		a<�`<��`<mxa<�[b<n]c<�@d<U�d<��d<�d<��c<~�b<�a<�$a< �`<<�`<�[a<��a<�]b<�{b<Kb<�"a<_�_<�]<�w[< FY<�UW<��U<�U<gU<.�U<,W<�Y<?D[<f|]<}_<da<�b<��b<��b<Nb<r�a<na<�`<�:a<Y�a<��b<��c<��d<xe<�e<Q~d<��c<�b<6�a<�a<�`<)%a<��a<�-b<��b<-~b<�a<I�`<;_<]<��Z<��X<r�V<�U<�
U<�AU<v5V<\�W<�Y<�\<�3^<	`<:|a<�Rb<��b<�cb<��a<�[a<Q�`<U�`<�ga<�3b<�1c<M%d<��d<�e<��d<�<d<�Mc<Mb<�xa<�`<D�`<La<��a<
Vb<��b<�^b<��a<�?`<�j^<NE\<�
Z<Q�W<XV<kPU<�U<�zU<��V<�gX<+�Z<�\<��^<��`<��a<�pb<H�b<�6b<N�a<I,a< �`<�
a<a�a<�~b<^�c<�cd<��d<	e<̱d<��c<��b<�a<mBa<J�`<�a<hta<Gb<crb<"�b<F)b<t0a<}�_<��]<�}[<�IY<�VW<��U<�U<_U<��U<�W<(Y<�2[<�h]<�f_<��`<� b<�sb<Vbb<�a<jga<��`<��`<a<��a<�b<��c<�{d<F�d<��d<�Rd<Wvc<�tb<e�a<��`<��`<��`<=xa<�b<�]b<�Rb<Ͻa<5�`<N�^<2�\<�Z<wsX<$�V<�dU<@�T<�U<V<��W<0�Y<��[<}�]<��_<�Ga<�b<bb<�-b<�a<9$a<5�`<��`<'.a<��a<�b<��c<��d<�d<[�d<�d<kc<Eb<�Aa<��`<�  �  KQa<��a<�`b<�b<c<��b<�b<��`<��^<��\<�Z<��X<O'W<�.V<��U<5WV<yuW<!Y<�([<HQ]<]_<Za<Rb<��b<�!c<��b<�Gb<H�a<�La<�<a<i�a<q=b<�
c<3�c<�>d<`Vd<Jd<Fgc<�b<�a<aa<�Da<��a<@b<�b<�c<4c<��b<i�a<�H`<^^<�<\<� Z<GX<��V<�(V< V<��V<�X<�Y<[\<�1^<&(`<��a<`�b<�Gc<�@c<��b<�Bb<��a<�ja<}a<��a<جb<Byc<�!d<�zd<�nd<��c<�Ic<i{b<��a<Fia<
na<U�a<�^b<��b<�Fc<i3c<.�b<aja<�_<$�]<��[<f�Y<��W<��V<�V<�OV<�5W<ӶX<��Z<s�\<��^<��`<�&b<�c<�Qc<�$c<Ȧb<�b<ґa<�aa<*�a<�(b<a�b<�c<�Hd<��d<�Sd<U�c<�c<�;b<�a<�`a<t�a<��a<�b<�c<�Oc<�c<�Cb</�`<�_<]<��Z<K�X<�VW<v]V<V<҄V<C�W<�LY<mS[< {]<��_<�<a<�xb<C%c<�Fc<��b<�kb<��a<�oa<�_a<Y�a<_`b<�-c<��c<ad<�xd<�)d<?�c<�b<�a<�~a<�`a<%�a<�*b<|�b<g2c<YFc<��b<��a<�S`<�f^<�B\<($Z<�GX<��V<y$V<V<�V<`X<F�Y<�[<'^<�`<��a<w�b<�*c<�!c<��b<�b<�a<�Da<�Ua<�a<J�b<�Nc<�c<�Od<QCd<��c<�c<gPb<Ƞa<�>a<�Ca<�a<4b<��b<�c<�c<�jb<0=a<�_<4�]<�c[<�UY<J�W<dmV<�U<�V<mW<�X<�qZ<W�\<��^<5�`<��a<��b<[c<��b<(pb<j�a<�Ya<�(a<�]a<��a<�b<}{c<�d<�Fd<Ud<��c<��b<�b<�ja<q*a<�  �  �b<�b<�bc<>�c<�d<!�c<��b<��a<��_<*�]<��[<�Z<˪X<��W<��W<��W<��X<�sZ<�R\<AW^< J`<��a<�4c<l�c<]d<2�c<�Gc<G�b<6b<��a<��a<�a<cwb<��b<Gc<"Xc<�!c<@�b<�4b<#�a<&�a<��a<^b<�	c</�c<Zd<�'d<*�c<άb</a<cW_<�U]<�`[<��Y<:uX<�W<b�W<�^X<��Y<�5[<�(]<+._<�a<�b<��c<+:d<1@d<_�c<�<c<�b<mb<��a<��a<�Mb<\�b<�?c<�}c<�tc<�'c<$�b<G/b<��a<��a<kb<#�b<�\c<J�c<�Cd<�"d<�zc<�Kb<P�`<�^<z�\<��Z<�EY<�7X<��W<�W<��X<�Z<��[<��]<��_<��a<\c<�c<�Hd<'d<ԩc<@�b<�Zb<��a<��a<�b<<ub<��b<�Yc<��c<yac<�c<�b<�b<d�a<:�a<�Ib<��b<5�c<�d<rHd<~�c<�$c<3�a<Y`<n^<�\<�BZ<R�X<��W<��W<�X<�Y<��Z<�}\<5�^<�r`<�b<�[c<(d<GBd<o�c<�kc<��b<S&b<��a<��a<�b<8�b<dc<�ic<?zc<dCc<�b<�Tb<��a<��a<��a<exb<>"c<��c<�2d</:d<�c<O�b<(:a<�__<�[]<ld[<ɱY<psX<��W<Z�W<UX<��Y<('[<9]<]_<��`<n�b<��c< d<!d<K�c<�c<�lb<\�a<&�a<�a<_$b<1�b<�c<�Rc<�Ic<��b<�b<Sb<׭a<-�a<��a<��b<X2c<h�c<od<��c<Nc<3b<|`<��^<o�\<�Z<SY<YX<ΐW<��W<։X<��Y<ި[<��]<��_<ma<��b<��c<_d<*�c<Tsc<�b<	#b<�a<b�a<��a<';b<��b<�c<�Gc<�'c<H�b<*Jb<�a<k�a<:�a<�  �  ��b<��c<�dd<��d<fe<��d<�c<j|b<��`<�_<3B]<��[<%�Z<6�Y<+�Y<��Y<�Z<�\<j�]<js_<�=a<��b<�d<l�d<	e<��d<hGd<��c<�b<�
b<�a<�a<
�a<��a<n�a<��a<5�a<��a<��a<R�a<8�a<mb<@0c<Cd<!�d<�e<e<��d<��c<�b<Z_`<��^<��\<�f[<_Z<��Y<��Y<UMZ<cJ[<��\<�h^<�:`< �a<]vc<U�d<S#e<�9e<$�d<�6d<�hc<|�b<�b<(�a<��a<��a<w�a<�b<b<�a<��a<)�a<��a<&#b<f�b<�c<�Zd<��d<g:e<�e<Ud<5(c<�a<�_<�^<�`\<r[<p/Z<��Y<��Y<x�Z<�[<�E]<B_<�`<��b<q�c<[�d<�7e<*%e<��d<��c<� c<Ngb<�a<I�a<2�a<��a<>
b<b<�b<�a<�a<U�a<V�a<mTb<�c<��c<ɗd<e<B9e<c�d<�c<6�b<�a<9_<�r]<��[<��Z<��Y<
�Y<0Z<B�Z<
3\<��]<��_<�fa<��b<r5d<`�d<"7e<��d<>kd<�c<-�b<�-b<��a<��a<ɻa<��a<�b<�b<��a<>�a<z�a<��a<��a<�b<pJc<�d<��d<.e<)%e<Λd<��c<�!b<�g`<|�^<��\<rg[<6]Z<R�Y<��Y<�CZ<*>[<̤\<_W^<'`<��a<�]c<�pd<Ze<�e<(�d<�d<%Dc<�}b<��a<ʔa<��a<��a<��a<��a<	�a<��a<��a<Da<ؘa<��a<��b<_fc<B0d<��d<�e<��d<C(d<��b<�la<��_<��]<w/\<}�Z<��Y<}�Y<��Y<�iZ<΋[<Y]<��^<��`<Pb<��c<^�d<Ae<_�d<�ud<��c<��b</b<I�a<�ua<o|a<ɥa<+�a<�a<��a<c�a<��a<�ta<��a<�b<�  �  �Yc<PVd<�%e<֢e<��e<�Ee<�dd<�$c<o�a<5`<�^<oh]<��\<��[<g�[<�\<��\<0�]<��^<]t`<b<:wc<¥d<�ne<z�e<��e<|e<�+d<�+c<�/b<�[a<�`<�k`<�B`<�4`<e3`<<`<�X`<��`<$a<��a<��b<o�c<h�d<&te<��e<,�e<$e<G!d<'�b<�Ca<��_<T^<6]<�q\<�\<�
\<f\<?"]<�9^<Қ_<�%a<��b<�d<�"e<��e<%�e<��e<��d<�d<�c<b<Oa<r�`<o�`<Ge`<�[`<�[`<�g`<2�`<��`<�oa<B=b<56c<�7d<,e<��e<�e<�e<w�d<��c<p\b<��`<wK_<_�]<��\<�R\<�\<)\<r�\<�}]<�^<"!`<��a<b0c<�xd<
fe<��e<��e<#me<��d<��c<��b<x�a<La<��`<�t`<�^`<�Y`<y]`<op`<��`<A	a<B�a<�b<E�c<"�d<�Xe<;�e<q�e<<we<�d<�Uc<;�a<�I`<s�^<՘]<Գ\<�.\<�	\<`C\<o�\< �]<Y_<��`<y-b<��c<��d<�e<��e<�e<u+e<,Od<�Nc<�Rb<�~a<��`<��`<e`<�V`<4U`<A]`<y`<&�`<�6a<��a<7�b<x�c<��d<m�e<�e<0�e<�3e<�.d<�b<La<�_<vW^<�6]<'p\<
\<�\<r\\<]<�*^<��_<8a<��b<�c<e<��e<3�e<�e<��d<��c<��b<��a<�&a<R�`<�Z`<�:`<�0`<�0`<�<`<Eb`<-�`<Ea<�b<�c<`d<\�d<��e<k�e<�{e<o�d<ܚc<�-b<%�`<�_<��]<��\< \<�[<-�[<Ho\<�I]<�z^<��_<){a<��b<DDd<1e<X�e<�e<�6e<�nd<Luc<�rb<��a<L�`<Jr`<�:`< %`<�`<:$`<�7`<uj`<��`<�wa<sXb<�  �  �~c<��d<Oye<��e<��e<lpe<:�d<oc<�*b<��`<�_< _<�w^<r*^<�^<07^<:�^< 0_<�`<�3a<Mwb<�c<n�d<n�e<��e<��e<�Ze<=pd<�Dc<�a<��`<S�_<��^<�s^<71^<"&^<Q^<��^<#a_<5P`<
ya<u�b<T�c<�e<��e<3f<��e<�Me<Vd<�#c<N�a<��`<��_<�^<k|^<�C^<PB^<.w^<#�^<��_<ǘ`<Z�a<Yc<
Jd<�Le<)�e<b0f<_�e<�Ce<0?d<Rc<=�a<��`<E�_<��^<��^<�O^<U^<e�^<c_<W�_<��`<�b<�Hc<Nyd<pme<jf<s)f<�e<�e<d<9�b<�a<m``<tv_<��^<�p^<�I^<�X^<��^<�%_<��_<�`<�9b<�c<5�d<
�e<�f<�&f<�e<��d<9�c<��b<Ta<�7`<�X_<f�^<:h^<XJ^<�a^<D�^<C_<�`<1a<pb<p�c<?�d<B�e<f<kf<�e<x�d<4�c<�[b<}a<�	`<�5_<
�^<�Z^<�E^<.f^<i�^<;]_<�?`<�^a<#�b<��c<��d<��e<"f<h
f<e<ߓd<�gc<"b<j�`<�_<_<U�^<ES^<�G^</r^<I�^<��_<~n`<�a<��b<4d<�#e<$�e<I(f<|�e<`]e<^cd<�.c<��a<�`<��_<��^<�z^<�?^<H;^<�m^<��^<��_<��`<��a<D�b<�1d<�1e<\�e<�f<��e<`!e<d<��b<P�a<}k`<Su_<-�^<NV^<%^<N*^<�f^<��^<��_<�`<��a<c<�Nd<�Be<�e<��e<��e<8�d<��c<�b<�Ta<i/`<�D_<��^<0=^<�^<u$^<k^<�^<A�_<c�`<.b<�Jc<xtd<%[e<]�e<�e< �e<~�d<2�c<�]b<�a<	�_<�_</�^<�.^<2^<)^<�y^<�_<��_<��`<�:b<�  �  �6c<sd<GNe<��e<Ξe<�e<:Jd<�Lc<�Lb<yoa<|�`<�i`<�9`<�'`<�$`<�*`<EB`<�|`<�`<"�a<ևb<f�c<ԃd<�He<V�e<��e<'1e<�>d<��b<�pa<��_<�t^<�H]<[t\<, \<��[<�6\<_�\<�]<OA_<��`<MVb<�c<�d<��e<��e<X�e<��d<�d<c<-b<kTa<��`<_y`<�V`<L`<�L`<eX`<Hz`<a�`<�Ma<�b<�	c<�d<r�d<��e<��e<K�e<�e<�d<d�b<a<��_<a3^<�!]<l\<�\<� \<P�\<IT]<nw^<�_<la<��b<�Ed<�Ce<V�e<_�e<�e<n�d<��c<��b<��a<
/a<`�`<xx`<�^`<�W`<Z`<fj`<\�`<g�`<d�a<�eb<Ecc<cd<e<e<�e<_�e<דe<u�d<4�c<Qb<X�`<{_<��]<��\<�B\<2\<,8\<�\<ث]<�^<�b`<��a<1kc<��d<�e<�e<��e<aNe<�{d<�}c<~b<��a<��`<֚`<�j`<TX`<�T`<Z`<�p`<Q�`<a<��a<�b<g�c<��d<Moe<!�e<��e<nUe<�bd<Rc<�a<a`<��^<Uk]<��\<"\<N\<�W\<�]<D
^<g__<��`<�qb<��c<�d<��e<��e<)�e<y
e<�#d<�c<�&b<FZa<��`<z`<�T`<�G`<�E`<�N`<n`<��`<�<a<��a<��b<0�c<��d<�e<8�e<��e<s�d<��c<�}b<[�`<�g_<�
^<W�\<B\<Z�[<,�[<�_\<�)]<�L^<r�_<�Aa<�b<d<�e<ܥe<S�e<EWe<ۚd<b�c<@�b<�a<��`<�`<qE`<+`<�#`<�%`<�5`<�a`<��`<�Ya<1b<�.c<P.d<�e<�e<�e<^e<<�d<u\c<	�a<�W`<<�^<?�]<"�\<
\<t�[<��[<"�\<ut]<r�^<�,`<r�a<�  �  �b<`�c<ڲd<ye<��d<�[d<��c<.�b<b<z�a<�va<ƅa<��a<��a<q�a<'�a<��a<��a<�}a<.�a<P?b<��b<4�c<*�d<��d<}	e<ߗd<��c<nEb<]�`<��^<�]<��[<+kZ<i�Y<֮Y<Z<1�Z<rV\<�^<�_<��a<�!c<�Id<��d<�#e<��d<v<d<�qc<C�b<�	b<��a<[�a<Q�a<7�a<�b<�b<�a<�a<2�a<)�a<~
b<�b<fnc<c=d<V�d<z;e<�e<X�d<�hc<\�a<R)`<�X^<2�\<�E[<YPZ<��Y<�Y<\zZ<�[<��\<ź^<$�`<p@b<۫c<��d<n,e<�-e<�d<�d<�?c<�b<��a<*�a<0�a<��a<!b<_b<�b<��a<�a<��a<�a<�;b<�b<��c<�{d<�e<�=e<��d<�-d<��b<Ua<9�_<a�]<P$\<�Z<�Z<a�Y<�	Z<��Z<@�[<�]<�U_<�"a<(�b<�d<��d<�:e<�e<_�d<��c<��b<wIb<��a<1�a<"�a<��a<�
b<�b<�b<��a<��a<v�a<��a<�ib<G%c<W�c<1�d<�"e<�.e<L�d<��c<�hb<k�`<{�^<i)]<�[<D�Z<*�Y<#�Y<�6Z<$[<xu\<�^<��_<�a<q;c<�ad<�e<e7e<��d<�Kd<c<�b<b<��a<��a<	�a<\�a<b<�b<y�a<޶a<��a<��a<��a<�b<Vc<�"d<��d<�e<A�d<`d<�Dc<�a<�`<A1^<�\<K[<}&Z<��Y<��Y<�OZ<|^[<�\<3�^<�``<�b<�c<r�d<� e<Te<�d<��c<c<\Pb<��a<sa<�|a<S�a<�a<��a<��a<�a<�a<�ta<'�a<�b<Q�b<:�c<Gd<��d<�e<Z�d<��c<p�b<a<�R_<|�]<�[<��Z<"�Y<�Y<��Y<F�Z<1�[<�W]< _<��`<�  �  �a<;c<9�c<�d<��c<�Zc<F�b<mb<��a<8�a<L�a<�Tb<^�b<0/c<�Kc<= c<@�b<�9b<$�a<n�a<��a<�2b<�b<��c<�c<�d<(�c<��b<gaa<#�_<=�]<֚[<*�Y<шX<��W<��W<� X<8Y<O�Z<��\<ý^<Ψ`<Fb<ioc<1d</,d<��c<z?c<��b<kb<�a< �a<_$b<��b<c<Pgc<�lc<%,c<�b<;b<�a<-�a<�	b<�b<PBc<��c<_Bd<X7d<�c<čb<^�`<�_<h]<�&[<��Y<%_X<��W<<�W<�X<��Y<��[<'�]<��_<Za<u�b<P�c<�@d<�1d<e�c<�c<�pb<r�a<��a<��a<e]b<�b<�Jc<L~c<jc<[c<��b<b<�a<?�a<�3b<��b<�{c<�
d<�Id<�d<MTc<Eb<L_`<k^<�g\<��Z<�Y<}X<��W<�	X<��X<�]Z<�/\<�0^<^)`<��a<{5c<�d<�Hd<�d<,�c<��b<�?b<&�a<��a<�b<:�b<�c<d`c<�|c<_Pc<��b<+hb<n�a<��a<p�a<c\b<kc<۫c<F%d<�@d<��c<��b<ڄa<6�_<�]<]�[<r�Y<ϪX<��W<��W<AX<�WY<.�Z<��\<A�^<��`<_b<�c<�&d<�?d<0�c<�Nc<��b<"b<G�a<��a<�'b<K�b<9c<�bc<�ec<�"c<ʭb<\,b<��a<��a<��a<�{b<�'c<��c<�#d<�d<��c<�ib<)�`<�^<��\<n�Z<�\Y<m5X<��W<�W<qhX<8�Y<b[<�Y]<�Z_<c/a<��b<
�c<�d<7d<:�c<��b<�Ab<l�a<{�a<��a<�*b<p�b<Uc<�Ic<�4c<�b<Abb<��a<�a<I�a<��a<�b<�Fc<��c<�d<,�c<~c<�a<�(`<�3^<>0\<�UZ<��X<W�W<��W<��W<��X<�&Z<|�[<�]<��_<�  �  ��`<� b<��b<Rc<T�b<�Xb<��a<PNa<-a<�sa<�b<x�b<�c<�"d<�Jd<�d<�vc<D�b<��a<�^a<l0a<�fa<��a<�b<�b<T%c<��b<-�a<�|`<��^<�\<caZ<xX<��V<�#V<�U<�V<4�W<~�Y<=�[<޼]<��_<Bea<��b<!!c<�.c<��b<*Bb<�a<�Xa</Za<��a<6ub<Dc<��c<bd<6id<�d<�`c<C�b<�a<�oa<ea<�a<Gb<��b<�Cc<�Ec<�b<&�a<�`<^<�[<��Y<X<��V<�)V<�=V<�W<�nX<�NZ<m\<��^<�t`<�a<Q�b<Lc<�0c<{�b<�#b<R�a<�`a<��a<�b<6�b<�c<h3d<$}d<r`d<$�c<'c<�Zb<��a<�ca<�ya<��a<{b<bc<Oc<�&c<rb<M.a<q_<c]<�;[<Z8Y<
�W<UV<=V<4kV<HmW<�Y<��Z<V%]<�8_<Za<�Sb<}c<}Oc</c<\�b<9�a<�a<�^a<[�a<�Bb<Lc<��c<�Sd<�{d<!=d<J�c<��b<�b<J�a<�[a<��a<`b<��b<}#c<�Jc<d�b<.b<u�`<
�^<٥\<�Z<=�X<p!W<sEV<V<}�V<��W<>�Y<�[<@�]<��_<�~a<B�b<�6c<^Bc<t�b<�Qb<-�a<Vca<mba<��a<sxb<�Dc<��c<�]d</bd<Dd<�Tc<��b<��a<9\a<Oa<�a<�,b<J�b<%c<J%c<��b<v�a<��_<��]<��[<=�Y< �W<��V<��U<bV<��V<�DX<$Z<�B\<
c^<�I`<�a<��b<$ c<Hc<)�b<��a<pa<J0a<BSa<z�a<�b<�`c<��c<)Hd<*+d<��c<��b<T%b<s�a<�.a<Ea<�a<>Fb<��b<c<<�b<r<b<6�`<�:_< ,]<+[<� Y</\W<nGV<r�U<�3V<-6W<�X<�Z<�\<z_<�  �  T$`<�ua<'3b<zab<�b<͙a<*a<]�`<��`<�Ma<�%b<�%c<d<��d<��d<^�d<��c<p�b<��a<,a<!�`<��`<p3a<��a<*<b<�kb<�b<Ba<*�_<�]<e�[<��Y<g�W<9�U<RU<~�T<I�U<1�V<��X<��Z<�]<g_<C�`<U�a<kb<Rpb<�b<�a<�a<;�`<�a<�a<˜b<\�c<�wd<�d<M�d<$�d<=�c<��b<c�a<%*a<��`<�a<��a<b<p�b<��b<�b<�a<Hi_<�e]<�-[<Y<F W<,�U<�U<.U<�V<�~W<1uY<4�[<[�]<T�_<kHa<�7b<M�b<�pb<��a<sna<�a<��`<kKa<
b<�c<��c<��d<�e<��d<.]d< wc<�ub<m�a<�a<��`<9a<$�a<bDb<4�b<�rb<�a<#�`<��^<8�\<lZ<RX<x�V<htU<�U<�^U<�oV<�X<-Z<�g\<��^<X`<��a<�eb<��b<qOb<}�a<�Ca<	�`<� a<�a<�Wb<�Wc<�Cd<-�d<e<��d<_d<>c<s b<�Xa<_�`<��`<(\a<�a<�bb<�b<�Db<fa<��_</^<(�[<�Y<��W< V<�6U<|U<��U<��V</�X<C�Z<!]<H-_<��`<��a<(�b<��b<}#b<m�a<�a<��`<�a<��a<�b<
�c<�ud<��d<G�d<��d<�c<>�b<H�a<�a<��`<��`<?sa<��a<�eb<�nb<��a<R�`<:D_<S?]<M[<��X<H�V<��U<��T<�U<v�U<~TW<�JY<�~[<ů]<��_<ja<b<^gb<�Cb<�a<@a<��`<��`<a<��a<x�b<��c<��d<��d<�d<�'d<tAc<e@b<&aa<��`<ջ`<7a<f�a<�b<>]b<=b<��a<'O`<R�^<`p\<�4Z<�X<�`V<�<U<Z�T<h'U<�8V<x�W<G�Y<w2\<%U^<�  �  /�_<�6a<A�a<vb<��a<Ra<�`<�`<��`<,>a<�*b<�=c<U8d<|�d<�e<��d<d<0c<A�a<a<��`<��`<>�`<�wa<��a<n&b<��a<ua<��_<'�]<�{[<�=Y<�5W<ͣU<��T<:�T<&U<itV<6QX<@�Z<��\<�^<~`<��a<c(b<�(b<��a<nAa<H�`<ݪ`<��`<T�a<s�b<��c<�d<�(e<�1e<R�d<�c<��b<�a<�a<��`<�`<�Ha<��a<�<b<[Kb<��a<��`<2*_<H#]<��Z<��X<J�V<LiU<��T<�T<�U<�)W<�'Y<�b[<��]<��_<�	a<��a<�Nb<6(b<��a<T+a< �`<��`<I5a<Rb<�c<�d<��d<�Ge<1#e<Ԅd<��c<%}b<G�a<��`<�`<"�`<va<G�a<�Kb<g0b<Ԇa<G`<ڂ^<;c\<�!Z< X<Z?V<|U<��T<|U<V<��W<�Y<#\<\I^<�`<�ia<�#b<�Mb<ub<��a<�a<��`<h�`<pa<�\b<�oc<:jd<!e<$Ge<5�d<�6d<1c<!b<�Da<+�`<��`<a<H�a<	b<�Kb<b<�'a<<�_<A�]<��[<M`Y<XW<��U<�T<3�T<fFU<��V<�oX<ϞZ<,�\<��^<_�`<�a<>b<�<b<K�a<�Pa<L�`<��`<�`<�a<��b<-�c< �d<y$e<�*e<��d<��c<��b<��a<�`<�`<��`<[.a<\�a<Eb<+b<±a<�`<)_< �\<��Z<j�X<Q�V<�?U<��T<�T<�}U<2�V<�X<g8[<fn]<�`_<��`<J�a<�"b<��a<#�a<��`<��`<z�`<�a<��a<1�b<}�c<:�d<�e<��d<?Od<[c<�Gb<�Sa<͵`<%�`<X�`<GAa<}�a<�b<3�a<IQa<`<yL^<n,\<��Y<��W<�V<��T<rT<*�T<5�U<��W<F�Y<��[<�^<�  �  T$`<�ua<'3b<zab<�b<͙a<*a<]�`<��`<�Ma<�%b<�%c<d<��d<��d<^�d<��c<p�b<��a<,a<!�`<��`<p3a<��a<*<b<�kb<�b<Ba<*�_<�]<e�[<��Y<g�W<9�U<RU<~�T<I�U<1�V<��X<��Z<�]<g_<C�`<U�a<kb<Rpb<�b<�a<�a<;�`<�a<�a<˜b<\�c<�wd<�d<M�d<$�d<=�c<��b<c�a<%*a<��`<�a<��a<b<p�b<��b<�b<�a<Hi_<�e]<�-[<Y<F W<,�U<�U<.U<�V<�~W<1uY<4�[<[�]<T�_<kHa<�7b<M�b<�pb<��a<sna<�a<��`<kKa<
b<�c<��c<��d<�e<��d<.]d< wc<�ub<m�a<�a<��`<9a<$�a<bDb<4�b<�rb<�a<#�`<��^<8�\<lZ<RX<x�V<htU<�U<�^U<�oV<�X<-Z<�g\<��^<X`<��a<�eb<��b<qOb<}�a<�Ca<	�`<� a<�a<�Wb<�Wc<�Cd<-�d<e<��d<_d<>c<s b<�Xa<_�`<��`<(\a<�a<�bb<�b<�Db<fa<��_</^<(�[<�Y<��W< V<�6U<|U<��U<��V</�X<C�Z<!]<H-_<��`<��a<(�b<��b<}#b<m�a<�a<��`<�a<��a<�b<
�c<�ud<��d<G�d<��d<�c<>�b<H�a<�a<��`<��`<?sa<��a<�eb<�nb<��a<R�`<:D_<S?]<M[<��X<H�V<��U<��T<�U<v�U<~TW<�JY<�~[<ů]<��_<ja<b<^gb<�Cb<�a<@a<��`<��`<a<��a<x�b<��c<��d<��d<�d<�'d<tAc<e@b<&aa<��`<ջ`<7a<f�a<�b<>]b<=b<��a<'O`<R�^<`p\<�4Z<�X<�`V<�<U<Z�T<h'U<�8V<x�W<G�Y<w2\<%U^<�  �  ��`<� b<��b<Rc<T�b<�Xb<��a<PNa<-a<�sa<�b<x�b<�c<�"d<�Jd<�d<�vc<D�b<��a<�^a<l0a<�fa<��a<�b<�b<T%c<��b<-�a<�|`<��^<�\<caZ<xX<��V<�#V<�U<�V<4�W<~�Y<=�[<޼]<��_<Bea<��b<!!c<�.c<��b<*Bb<�a<�Xa</Za<��a<6ub<Dc<��c<bd<6id<�d<�`c<C�b<�a<�oa<ea<�a<Gb<��b<�Cc<�Ec<�b<&�a<�`<^<�[<��Y<X<��V<�)V<�=V<�W<�nX<�NZ<m\<��^<�t`<�a<Q�b<Lc<�0c<{�b<�#b<R�a<�`a<��a<�b<6�b<�c<h3d<$}d<r`d<$�c<'c<�Zb<��a<�ca<�ya<��a<{b<bc<Oc<�&c<rb<M.a<q_<c]<�;[<Z8Y<
�W<UV<=V<4kV<HmW<�Y<��Z<V%]<�8_<Za<�Sb<}c<}Oc</c<\�b<9�a<�a<�^a<[�a<�Bb<Lc<��c<�Sd<�{d<!=d<J�c<��b<�b<J�a<�[a<��a<`b<��b<}#c<�Jc<d�b<.b<u�`<
�^<٥\<�Z<=�X<p!W<sEV<V<}�V<��W<>�Y<�[<@�]<��_<�~a<B�b<�6c<^Bc<t�b<�Qb<-�a<Vca<mba<��a<sxb<�Dc<��c<�]d</bd<Dd<�Tc<��b<��a<9\a<Oa<�a<�,b<J�b<%c<J%c<��b<v�a<��_<��]<��[<=�Y< �W<��V<��U<bV<��V<�DX<$Z<�B\<
c^<�I`<�a<��b<$ c<Hc<)�b<��a<pa<J0a<BSa<z�a<�b<�`c<��c<)Hd<*+d<��c<��b<T%b<s�a<�.a<Ea<�a<>Fb<��b<c<<�b<r<b<6�`<�:_< ,]<+[<� Y</\W<nGV<r�U<�3V<-6W<�X<�Z<�\<z_<�  �  �a<;c<9�c<�d<��c<�Zc<F�b<mb<��a<8�a<L�a<�Tb<^�b<0/c<�Kc<= c<@�b<�9b<$�a<n�a<��a<�2b<�b<��c<�c<�d<(�c<��b<gaa<#�_<=�]<֚[<*�Y<шX<��W<��W<� X<8Y<O�Z<��\<ý^<Ψ`<Fb<ioc<1d</,d<��c<z?c<��b<kb<�a< �a<_$b<��b<c<Pgc<�lc<%,c<�b<;b<�a<-�a<�	b<�b<PBc<��c<_Bd<X7d<�c<čb<^�`<�_<h]<�&[<��Y<%_X<��W<<�W<�X<��Y<��[<'�]<��_<Za<u�b<P�c<�@d<�1d<e�c<�c<�pb<r�a<��a<��a<e]b<�b<�Jc<L~c<jc<[c<��b<b<�a<?�a<�3b<��b<�{c<�
d<�Id<�d<MTc<Eb<L_`<k^<�g\<��Z<�Y<}X<��W<�	X<��X<�]Z<�/\<�0^<^)`<��a<{5c<�d<�Hd<�d<,�c<��b<�?b<&�a<��a<�b<:�b<�c<d`c<�|c<_Pc<��b<+hb<n�a<��a<p�a<c\b<kc<۫c<F%d<�@d<��c<��b<ڄa<6�_<�]<]�[<r�Y<ϪX<��W<��W<AX<�WY<.�Z<��\<A�^<��`<_b<�c<�&d<�?d<0�c<�Nc<��b<"b<G�a<��a<�'b<K�b<9c<�bc<�ec<�"c<ʭb<\,b<��a<��a<��a<�{b<�'c<��c<�#d<�d<��c<�ib<)�`<�^<��\<n�Z<�\Y<m5X<��W<�W<qhX<8�Y<b[<�Y]<�Z_<c/a<��b<
�c<�d<7d<:�c<��b<�Ab<l�a<{�a<��a<�*b<p�b<Uc<�Ic<�4c<�b<Abb<��a<�a<I�a<��a<�b<�Fc<��c<�d<,�c<~c<�a<�(`<�3^<>0\<�UZ<��X<W�W<��W<��W<��X<�&Z<|�[<�]<��_<�  �  �b<`�c<ڲd<ye<��d<�[d<��c<.�b<b<z�a<�va<ƅa<��a<��a<q�a<'�a<��a<��a<�}a<.�a<P?b<��b<4�c<*�d<��d<}	e<ߗd<��c<nEb<]�`<��^<�]<��[<+kZ<i�Y<֮Y<Z<1�Z<rV\<�^<�_<��a<�!c<�Id<��d<�#e<��d<v<d<�qc<C�b<�	b<��a<[�a<Q�a<7�a<�b<�b<�a<�a<2�a<)�a<~
b<�b<fnc<c=d<V�d<z;e<�e<X�d<�hc<\�a<R)`<�X^<2�\<�E[<YPZ<��Y<�Y<\zZ<�[<��\<ź^<$�`<p@b<۫c<��d<n,e<�-e<�d<�d<�?c<�b<��a<*�a<0�a<��a<!b<_b<�b<��a<�a<��a<�a<�;b<�b<��c<�{d<�e<�=e<��d<�-d<��b<Ua<9�_<a�]<P$\<�Z<�Z<a�Y<�	Z<��Z<@�[<�]<�U_<�"a<(�b<�d<��d<�:e<�e<_�d<��c<��b<wIb<��a<1�a<"�a<��a<�
b<�b<�b<��a<��a<v�a<��a<�ib<G%c<W�c<1�d<�"e<�.e<L�d<��c<�hb<k�`<{�^<i)]<�[<D�Z<*�Y<#�Y<�6Z<$[<xu\<�^<��_<�a<q;c<�ad<�e<e7e<��d<�Kd<c<�b<b<��a<��a<	�a<\�a<b<�b<y�a<޶a<��a<��a<��a<�b<Vc<�"d<��d<�e<A�d<`d<�Dc<�a<�`<A1^<�\<K[<}&Z<��Y<��Y<�OZ<|^[<�\<3�^<�``<�b<�c<r�d<� e<Te<�d<��c<c<\Pb<��a<sa<�|a<S�a<�a<��a<��a<�a<�a<�ta<'�a<�b<Q�b<:�c<Gd<��d<�e<Z�d<��c<p�b<a<�R_<|�]<�[<��Z<"�Y<�Y<��Y<F�Z<1�[<�W]< _<��`<�  �  �6c<sd<GNe<��e<Ξe<�e<:Jd<�Lc<�Lb<yoa<|�`<�i`<�9`<�'`<�$`<�*`<EB`<�|`<�`<"�a<ևb<f�c<ԃd<�He<V�e<��e<'1e<�>d<��b<�pa<��_<�t^<�H]<[t\<, \<��[<�6\<_�\<�]<OA_<��`<MVb<�c<�d<��e<��e<X�e<��d<�d<c<-b<kTa<��`<_y`<�V`<L`<�L`<eX`<Hz`<a�`<�Ma<�b<�	c<�d<r�d<��e<��e<K�e<�e<�d<d�b<a<��_<a3^<�!]<l\<�\<� \<P�\<IT]<nw^<�_<la<��b<�Ed<�Ce<V�e<_�e<�e<n�d<��c<��b<��a<
/a<`�`<xx`<�^`<�W`<Z`<fj`<\�`<g�`<d�a<�eb<Ecc<cd<e<e<�e<_�e<דe<u�d<4�c<Qb<X�`<{_<��]<��\<�B\<2\<,8\<�\<ث]<�^<�b`<��a<1kc<��d<�e<�e<��e<aNe<�{d<�}c<~b<��a<��`<֚`<�j`<TX`<�T`<Z`<�p`<Q�`<a<��a<�b<g�c<��d<Moe<!�e<��e<nUe<�bd<Rc<�a<a`<��^<Uk]<��\<"\<N\<�W\<�]<D
^<g__<��`<�qb<��c<�d<��e<��e<)�e<y
e<�#d<�c<�&b<FZa<��`<z`<�T`<�G`<�E`<�N`<n`<��`<�<a<��a<��b<0�c<��d<�e<8�e<��e<s�d<��c<�}b<[�`<�g_<�
^<W�\<B\<Z�[<,�[<�_\<�)]<�L^<r�_<�Aa<�b<d<�e<ܥe<S�e<EWe<ۚd<b�c<@�b<�a<��`<�`<qE`<+`<�#`<�%`<�5`<�a`<��`<�Ya<1b<�.c<P.d<�e<�e<�e<^e<<�d<u\c<	�a<�W`<<�^<?�]<"�\<
\<t�[<��[<"�\<ut]<r�^<�,`<r�a<�  �  �~c<��d<Oye<��e<��e<lpe<:�d<oc<�*b<��`<�_< _<�w^<r*^<�^<07^<:�^< 0_<�`<�3a<Mwb<�c<n�d<n�e<��e<��e<�Ze<=pd<�Dc<�a<��`<S�_<��^<�s^<71^<"&^<Q^<��^<#a_<5P`<
ya<u�b<T�c<�e<��e<3f<��e<�Me<Vd<�#c<N�a<��`<��_<�^<k|^<�C^<PB^<.w^<#�^<��_<ǘ`<Z�a<Yc<
Jd<�Le<)�e<b0f<_�e<�Ce<0?d<Rc<=�a<��`<E�_<��^<��^<�O^<U^<e�^<c_<W�_<��`<�b<�Hc<Nyd<pme<jf<s)f<�e<�e<d<9�b<�a<m``<tv_<��^<�p^<�I^<�X^<��^<�%_<��_<�`<�9b<�c<5�d<
�e<�f<�&f<�e<��d<9�c<��b<Ta<�7`<�X_<f�^<:h^<XJ^<�a^<D�^<C_<�`<1a<pb<p�c<?�d<B�e<f<kf<�e<x�d<4�c<�[b<}a<�	`<�5_<
�^<�Z^<�E^<.f^<i�^<;]_<�?`<�^a<#�b<��c<��d<��e<"f<h
f<e<ߓd<�gc<"b<j�`<�_<_<U�^<ES^<�G^</r^<I�^<��_<~n`<�a<��b<4d<�#e<$�e<I(f<|�e<`]e<^cd<�.c<��a<�`<��_<��^<�z^<�?^<H;^<�m^<��^<��_<��`<��a<D�b<�1d<�1e<\�e<�f<��e<`!e<d<��b<P�a<}k`<Su_<-�^<NV^<%^<N*^<�f^<��^<��_<�`<��a<c<�Nd<�Be<�e<��e<��e<8�d<��c<�b<�Ta<i/`<�D_<��^<0=^<�^<u$^<k^<�^<A�_<c�`<.b<�Jc<xtd<%[e<]�e<�e< �e<~�d<2�c<�]b<�a<	�_<�_</�^<�.^<2^<)^<�y^<�_<��_<��`<�:b<�  �  �Yc<PVd<�%e<֢e<��e<�Ee<�dd<�$c<o�a<5`<�^<oh]<��\<��[<g�[<�\<��\<0�]<��^<]t`<b<:wc<¥d<�ne<z�e<��e<|e<�+d<�+c<�/b<�[a<�`<�k`<�B`<�4`<e3`<<`<�X`<��`<$a<��a<��b<o�c<h�d<&te<��e<,�e<$e<G!d<'�b<�Ca<��_<T^<6]<�q\<�\<�
\<f\<?"]<�9^<Қ_<�%a<��b<�d<�"e<��e<%�e<��e<��d<�d<�c<b<Oa<r�`<o�`<Ge`<�[`<�[`<�g`<2�`<��`<�oa<B=b<56c<�7d<,e<��e<�e<�e<w�d<��c<p\b<��`<wK_<_�]<��\<�R\<�\<)\<r�\<�}]<�^<"!`<��a<b0c<�xd<
fe<��e<��e<#me<��d<��c<��b<x�a<La<��`<�t`<�^`<�Y`<y]`<op`<��`<A	a<B�a<�b<E�c<"�d<�Xe<;�e<q�e<<we<�d<�Uc<;�a<�I`<s�^<՘]<Գ\<�.\<�	\<`C\<o�\< �]<Y_<��`<y-b<��c<��d<�e<��e<�e<u+e<,Od<�Nc<�Rb<�~a<��`<��`<e`<�V`<4U`<A]`<y`<&�`<�6a<��a<7�b<x�c<��d<m�e<�e<0�e<�3e<�.d<�b<La<�_<vW^<�6]<'p\<
\<�\<r\\<]<�*^<��_<8a<��b<�c<e<��e<3�e<�e<��d<��c<��b<��a<�&a<R�`<�Z`<�:`<�0`<�0`<�<`<Eb`<-�`<Ea<�b<�c<`d<\�d<��e<k�e<�{e<o�d<ܚc<�-b<%�`<�_<��]<��\< \<�[<-�[<Ho\<�I]<�z^<��_<){a<��b<DDd<1e<X�e<�e<�6e<�nd<Luc<�rb<��a<L�`<Jr`<�:`< %`<�`<:$`<�7`<uj`<��`<�wa<sXb<�  �  ��b<��c<�dd<��d<fe<��d<�c<j|b<��`<�_<3B]<��[<%�Z<6�Y<+�Y<��Y<�Z<�\<j�]<js_<�=a<��b<�d<l�d<	e<��d<hGd<��c<�b<�
b<�a<�a<
�a<��a<n�a<��a<5�a<��a<��a<R�a<8�a<mb<@0c<Cd<!�d<�e<e<��d<��c<�b<Z_`<��^<��\<�f[<_Z<��Y<��Y<UMZ<cJ[<��\<�h^<�:`< �a<]vc<U�d<S#e<�9e<$�d<�6d<�hc<|�b<�b<(�a<��a<��a<w�a<�b<b<�a<��a<)�a<��a<&#b<f�b<�c<�Zd<��d<g:e<�e<Ud<5(c<�a<�_<�^<�`\<r[<p/Z<��Y<��Y<x�Z<�[<�E]<B_<�`<��b<q�c<[�d<�7e<*%e<��d<��c<� c<Ngb<�a<I�a<2�a<��a<>
b<b<�b<�a<�a<U�a<V�a<mTb<�c<��c<ɗd<e<B9e<c�d<�c<6�b<�a<9_<�r]<��[<��Z<��Y<
�Y<0Z<B�Z<
3\<��]<��_<�fa<��b<r5d<`�d<"7e<��d<>kd<�c<-�b<�-b<��a<��a<ɻa<��a<�b<�b<��a<>�a<z�a<��a<��a<�b<pJc<�d<��d<.e<)%e<Λd<��c<�!b<�g`<|�^<��\<rg[<6]Z<R�Y<��Y<�CZ<*>[<̤\<_W^<'`<��a<�]c<�pd<Ze<�e<(�d<�d<%Dc<�}b<��a<ʔa<��a<��a<��a<��a<	�a<��a<��a<Da<ؘa<��a<��b<_fc<B0d<��d<�e<��d<C(d<��b<�la<��_<��]<w/\<}�Z<��Y<}�Y<��Y<�iZ<΋[<Y]<��^<��`<Pb<��c<^�d<Ae<_�d<�ud<��c<��b</b<I�a<�ua<o|a<ɥa<+�a<�a<��a<c�a<��a<�ta<��a<�b<�  �  �b<�b<�bc<>�c<�d<!�c<��b<��a<��_<*�]<��[<�Z<˪X<��W<��W<��W<��X<�sZ<�R\<AW^< J`<��a<�4c<l�c<]d<2�c<�Gc<G�b<6b<��a<��a<�a<cwb<��b<Gc<"Xc<�!c<@�b<�4b<#�a<&�a<��a<^b<�	c</�c<Zd<�'d<*�c<άb</a<cW_<�U]<�`[<��Y<:uX<�W<b�W<�^X<��Y<�5[<�(]<+._<�a<�b<��c<+:d<1@d<_�c<�<c<�b<mb<��a<��a<�Mb<\�b<�?c<�}c<�tc<�'c<$�b<G/b<��a<��a<kb<#�b<�\c<J�c<�Cd<�"d<�zc<�Kb<P�`<�^<z�\<��Z<�EY<�7X<��W<�W<��X<�Z<��[<��]<��_<��a<\c<�c<�Hd<'d<ԩc<@�b<�Zb<��a<��a<�b<<ub<��b<�Yc<��c<yac<�c<�b<�b<d�a<:�a<�Ib<��b<5�c<�d<rHd<~�c<�$c<3�a<Y`<n^<�\<�BZ<R�X<��W<��W<�X<�Y<��Z<�}\<5�^<�r`<�b<�[c<(d<GBd<o�c<�kc<��b<S&b<��a<��a<�b<8�b<dc<�ic<?zc<dCc<�b<�Tb<��a<��a<��a<exb<>"c<��c<�2d</:d<�c<O�b<(:a<�__<�[]<ld[<ɱY<psX<��W<Z�W<UX<��Y<('[<9]<]_<��`<n�b<��c< d<!d<K�c<�c<�lb<\�a<&�a<�a<_$b<1�b<�c<�Rc<�Ic<��b<�b<Sb<׭a<-�a<��a<��b<X2c<h�c<od<��c<Nc<3b<|`<��^<o�\<�Z<SY<YX<ΐW<��W<։X<��Y<ި[<��]<��_<ma<��b<��c<_d<*�c<Tsc<�b<	#b<�a<b�a<��a<';b<��b<�c<�Gc<�'c<H�b<*Jb<�a<k�a<:�a<�  �  KQa<��a<�`b<�b<c<��b<�b<��`<��^<��\<�Z<��X<O'W<�.V<��U<5WV<yuW<!Y<�([<HQ]<]_<Za<Rb<��b<�!c<��b<�Gb<H�a<�La<�<a<i�a<q=b<�
c<3�c<�>d<`Vd<Jd<Fgc<�b<�a<aa<�Da<��a<@b<�b<�c<4c<��b<i�a<�H`<^^<�<\<� Z<GX<��V<�(V< V<��V<�X<�Y<[\<�1^<&(`<��a<`�b<�Gc<�@c<��b<�Bb<��a<�ja<}a<��a<جb<Byc<�!d<�zd<�nd<��c<�Ic<i{b<��a<Fia<
na<U�a<�^b<��b<�Fc<i3c<.�b<aja<�_<$�]<��[<f�Y<��W<��V<�V<�OV<�5W<ӶX<��Z<s�\<��^<��`<�&b<�c<�Qc<�$c<Ȧb<�b<ґa<�aa<*�a<�(b<a�b<�c<�Hd<��d<�Sd<U�c<�c<�;b<�a<�`a<t�a<��a<�b<�c<�Oc<�c<�Cb</�`<�_<]<��Z<K�X<�VW<v]V<V<҄V<C�W<�LY<mS[< {]<��_<�<a<�xb<C%c<�Fc<��b<�kb<��a<�oa<�_a<Y�a<_`b<�-c<��c<ad<�xd<�)d<?�c<�b<�a<�~a<�`a<%�a<�*b<|�b<g2c<YFc<��b<��a<�S`<�f^<�B\<($Z<�GX<��V<y$V<V<�V<`X<F�Y<�[<'^<�`<��a<w�b<�*c<�!c<��b<�b<�a<�Da<�Ua<�a<J�b<�Nc<�c<�Od<QCd<��c<�c<gPb<Ƞa<�>a<�Ca<�a<4b<��b<�c<�c<�jb<0=a<�_<4�]<�c[<�UY<J�W<dmV<�U<�V<mW<�X<�qZ<W�\<��^<5�`<��a<��b<[c<��b<(pb<j�a<�Ya<�(a<�]a<��a<�b<}{c<�d<�Fd<Ud<��c<��b<�b<�ja<q*a<�  �  �`<�a<=�a<z#b<�bb<T-b<�ga<A`<�:^<F\<�Y<��W<�(V<�!U<��T<=MU<{V<G<X<�ZZ<w�\<U�^<Yl`<<�a<|Kb<�db<�b<��a<		a<�`<��`<mxa<�[b<n]c<�@d<U�d<��d<�d<��c<~�b<�a<�$a< �`<<�`<�[a<��a<�]b<�{b<Kb<�"a<_�_<�]<�w[< FY<�UW<��U<�U<gU<.�U<,W<�Y<?D[<f|]<}_<da<�b<��b<��b<Nb<r�a<na<�`<�:a<Y�a<��b<��c<��d<xe<�e<Q~d<��c<�b<6�a<�a<�`<)%a<��a<�-b<��b<-~b<�a<I�`<;_<]<��Z<��X<r�V<�U<�
U<�AU<v5V<\�W<�Y<�\<�3^<	`<:|a<�Rb<��b<�cb<��a<�[a<Q�`<U�`<�ga<�3b<�1c<M%d<��d<�e<��d<�<d<�Mc<Mb<�xa<�`<D�`<La<��a<
Vb<��b<�^b<��a<�?`<�j^<NE\<�
Z<Q�W<XV<kPU<�U<�zU<��V<�gX<+�Z<�\<��^<��`<��a<�pb<H�b<�6b<N�a<I,a< �`<�
a<a�a<�~b<^�c<�cd<��d<	e<̱d<��c<��b<�a<mBa<J�`<�a<hta<Gb<crb<"�b<F)b<t0a<}�_<��]<�}[<�IY<�VW<��U<�U<_U<��U<�W<(Y<�2[<�h]<�f_<��`<� b<�sb<Vbb<�a<jga<��`<��`<a<��a<�b<��c<�{d<F�d<��d<�Rd<Wvc<�tb<e�a<��`<��`<��`<=xa<�b<�]b<�Rb<Ͻa<5�`<N�^<2�\<�Z<wsX<$�V<�dU<@�T<�U<V<��W<0�Y<��[<}�]<��_<�Ga<�b<bb<�-b<�a<9$a<5�`<��`<'.a<��a<�b<��c<��d<�d<[�d<�d<kc<Eb<�Aa<��`<�  �  �0\<�\<�]<��^<3�_<�!`<��_<
8^<h\<�\Y<�uV<�S<pQ<7�O</�O<8P<L�Q<gIT<�W<� Z<4�\<e�^<��_<�'`<1�_<��^<��]<��\<:9\<�\<��]<�|_<Ia<F�b<��c<��c<sZc<�	b<�P`<�^<� ]<3[\<a\<r]<!>^<�`_<u`<=,`<X]_<x�]<�T[<ĈX<y�U<S<��P<+�O<��O<y�P<z�R<�^U<�BX<�[<\�]<yM_<K8`<)E`<+�_<f^<tZ]<�\<�v\<X(]<��^<SF`<7b<�fc<d<�d<I"c<y�a<S�_<0&^<�\<#c\<9�\<Ս]<��^<��_<M`<7`<��^<J	]<;}Z<h�W<��T<OR<��P<��O<�P<DnQ<2�S<WV<?Y<��[<87^<ݴ_<�R`<�`<�?_<^<�]<Wn\<ϖ\<��]<�_<��`<M�b<ӷc<�,d<��c<��b<}a<-B_<��]<$�\<�f\<�\<�]<�_<r`<�S`<��_<�h^<?\<��Y<�V<;�S<��Q<�)P<�O<�fP<�R<�uT<�GW<�*Z<��\<��^<�_<M`<��_<t�^<�]<�\<�\\<U�\<��]<��_<ma<�b<��c<�d<~c<�,b<s`<�^<�@]<:y\<?}\<�6]<JV^<kv_<�2`<P=`<�k_<c�]<^[<Q�X<J�U<S<:�P<��O<��O<v�P<��R<OU<�0X<[<r]<�3_<�`<�&`<Nx_<p\^<�5]<;j\<�N\<��\<�[^<�`<��a<�9c<�c<y�c<f�b<�va<3�_<��]<ڼ\<D8\<�}\<>c]<��^<��_<{!`<��_<��^<#�\<NZ<=nW<m�T<R<�ZP<L�O<�O<:Q<�iS<w"V<Q
Y<�[<0^<�_<`<��_<�_<d�]<E�\<�4\<{\\<�M]<��^<�`<kKb<�zc< �c<,�c<.ub<��`<N_<�s]<�n\<�  �  ��\<�#]<�,^<�R_<1`<�s`<�_<�~^<�W\<��Y<!�V<$T<+�Q<�~P<�P<�P<[XR<b�T<lvW<POZ<s�\<�^<�`<�{`<�`<w_<�]<]<��\<z�\<� ^<�_<�;a<�b<'�c<��c<#0c<��a<�R`<;�^<i`]<9�\<��\< �]<S�^<��_<\x`<�z`<?�_<t�]<%�[<��X<�V<�sS<l|Q<pcP<�UP<NUQ<�9S<��U<I�X<�d[<��]<��_<��`<ʜ`<\�_<��^<6�]<��\<.�\<'k]<#�^<QK`<��a<>c<m�c<6�c<�b<F�a<�_<�P^<k1]<��\<�]<��]<�$_<�$`<\�`<1^`<�=_<3Q]<�Z<��W<,U<��R<*Q<3KP<��P<��Q<�
T<G�V<�Y<�D\<�}^<��_<o�`<dv`<U�_<m�^<�s]<��\<&�\<q�]<H+_<+�`<Rkb<��c<E�c<(�c<��b<a<3X_<��]<��\<��\<�X]<�`^<Ʌ_<Kc`<m�`<P`<��^<x�\<E�Y<�W<bNT<"R<�P<�BP<H�P<��R<��T<��W<CyZ<(]<�_<0E`<*�`<C6`<l@_<�^<g$]<�\<�]<�$^<��_<�_a<�b<W�c<��c<�Sc<�b<�t`<,�^<�]<8�\<
�\<a�]<v�^<��_<�`<�`<ó_<\^<d�[<z�X<�	V<�tS<�zQ<�^P<NNP<KKQ<-S<-�U<%�X<,P[<F�]<{_<�i`<+~`<��_<��^<R�]<�\<�\<A]<Q^<�`<)�a<'c<]�c<)�c<%�b<�fa<��_<�$^<1]<��\<U�\<��]<��^<n�_<�v`<�1`<o_<�"]<ԛZ<a�W<��T<��R<X�P<�P<dP<��Q<v�S<��V<.\Y<\<�H^<��_<�m`<2@`<o_<�L^<o;]<C�\<�\<Q�]<j�^<��`<�.b<�Mc<z�c<�cc<�Ub<*�`<c_<K�]<��\<�  �  ��]<%R^<!\_<nn`<�.a<Ta<��`<DA_<#]<��Z<��W<+PU<�BS<W�Q<̐Q<&+R<�S<��U<wuX<�,[<�]<�_<�`<;ba<}a<�=`<R&_<,^<��]<�]<{^<��_<�a<dAb<yc<�,c<��b<ڢa<2N`< _<�^<Ф]<X�]<4�^<��_<�`<�ka<�Ra<<k`<.�^<$r\<��Y<.W<(�T<��R<n�Q<��Q<�R<�~T<��V<�Y<y9\<�^<�Y`<$[a<ތa<(a<�`<��^<^<I�]<b^<�_<�O`<��a<�b<�Pc<=c<ևb<�Za<��_<
�^<��]<��]<�=^</_<TH`<�,a<�a<�.a<Q`<^<c�[<��X<�OV<nT<�|R<��Q<�R<�FS<�AU<��W<^xZ<\]<�@_<��`<��a<�pa<پ`<�_<O�^<��]<��]<�W^<$j_<��`<Eb<��b<!\c<c< .b<��`<3�_<o^<Q�]<��]<�^< �_<h�`<&aa<��a<��`<Br_<�S]<3�Z<z
X<��U<�rS<#R<��Q<�YR<��S<MV<נX<�V[<b�]<��_<�a<��a<-;a<�a`<�I_<{O^<��]<x�]<��^<]�_<�/a<�eb<�*c<�Pc<#�b<��a<)p`<� _<u(^<��]<z^<a�^<��_<��`<Ia<�ca<�y`<�^<\{\<C�Y<�W<4�T<(�R<��Q<]�Q<�R<�qT<�V<�xY<�$\<�}^<@`<�>a<Jna<\�`<�_<��^<w�]<�]<��]<�^<6$`<j|a<�b<�#c<c<[b<X.a<��_<i�^<��]<�]<�^<u_<`<�a<X`a<Oa<��_<��]<�u[<*�X<[V<.�S<�IR<F�Q<��Q<&S<UU<�W<�CZ<q�\<�_<H�`<Ka<�:a<�`<�z_<�j^<��]<��]<�^<x._<L�`<��a<C�b<�c<��b<��a< �`<�S_<�6^<
�]<�  �  l_<��_<��`<|�a<��b<6�b<�a<�L`<�@^<8�[<�_Y<BW<RHU<� T<��S<�QT<��U<�W<��Y<�i\<��^<'�`<�b<@�b<�zb<��a<W�`<O�_<�_<��^<_<L�_<U�`<�wa<�b<Ub<j�a<#a<)`<k\_<W�^<�^<n_<u]`<vma<1Nb<��b<�vb<�xa<��_<��]<m'[<��X<�V<m�T<�T<pT<M�T<ddV<X<4�Z<ig]<T�_<@fa<�{b<��b<�}b<�a<��`<�_<�_<H_<jq_<�8`<*a<��a<�Cb<p5b<J�a<�`<�`<�H_<��^<9!_<N�_<��`<��a<A�b<��b<0Ib<�a<�,_<��\<�aZ<�X<�V< �T<� T<�?T<�QU<�W<OY<\�[<�3^<M`<�a<��b<9�b<�>b<oNa<�@`<"d_<��^<�_<�_<x�`<�`a<	b<�Kb<�b<�va<<�`<��_<� _<��^<QP_<x"`<S.a<h%b<��b<�b<b�a<�}`<�q^<\<z�Y<�IW<�xU<�PT<a�S<��T<x�U<��W<LZ<F�\<��^<�`<I+b<��b<ٟb<��a<�`<��_<>*_<E�^<�4_<�_<D�`<��a<�&b<Bb<��a<�-a<�J`<}_<�_<�_<�_<�w`<m�a<�cb<��b<ȇb<*�a<��_<��]<�-[<X�X<�V<��T<	T<0 T<M�T<�WV<pX<�Z<�R]<�_<yLa<y_b<2�b<�\b<D�a<�w`<��_<��^<��^<�F_<`<��`<�a<�b<�b<��a<��`<��_< _<\�^<P�^<��_<�`<��a<�jb<�b<vb<$�`<Y�^<��\<(1Z<F�W<U�U<�lT<��S<NT<>U<��V<)Y<k�[<��]<�`<Ρa<wb<+�b<�b<a<|`<)+_<��^<�^<�m_<�E`<�$a<��a<Ib<��a<~;a<�_`<Q�_<B�^<x�^<�  �  ��`<>�a<�b<�vc<<�c<l�c</�b<\Ra<Ug_<~A]<�[<�2Y<ܰW<�V<7wV<d�V<~�W<ؙY<��[<:�]<=�_<�a<$c<%�c<&�c<Wc<�mb<�]a<i`<g�_<=�_<��_<��_<�C`<&�`<u�`<�h`<�`<D�_<��_<�_<�`<��`<Wb<v	c<#�c<m�c<N�c<{b<��`<v�^<W�\<��Z<5�X<0tW<�V<)�V<c[W<��X<�fZ<�y\<-�^<m�`<hb<`�c<�d<�c<�Ac<!Db<6a<kW`<��_<�_<a�_<�3`<T�`<ټ`<U�`<�v`<`<�_<M�_<7�_<z`<
ha<nxb<�ic<@�c<�c<�Vc<5b<ME`<�,^<j\<�Y<�UX<�/W<�V<#�V<�W<&6Y<�[<�7]< `_<�Ta<��b<P�c<d<��c<��b<1�a<��`<�`<�_<Ѵ_<`�_<�O`<�`<&�`<�`<Y`<)�_<9�_<��_<4
`<L�`<��a<��b<��c<ud<-�c<��b<��a<��_<�r]<�N[<�cY<��W<��V<'�V<�W<�*X<%�Y<��[<�]<�`<6�a<=6c<,�c<E�c<{{c<�b<a�a<~�`<��_<ʦ_<I�_<m`<ug`<�`<�`<�`<G7`<��_<u�_<�_<}<`<qa<@b<K!c<��c<�d<)�c<]�b<^�`<��^<ʰ\<v�Z<6�X<rrW<e�V<�V<eQW<�X<~WZ<�g\<��^<3�`<MNb<Csc<��c<��c<4c<�b<�a<�/`<l�_<��_<�_<�`<�]`<2�`<��`<�I`<��_<#�_<�~_<�_<,O`<8=a<�Mb<h>c<��c<��c<�)c<D�a<V`<��]<X�[< �Y<#X<J�V<�yV<|�V<3�W<Y<��Z<�]<+_<xa<E�b<��c<'�c<,�c<p�b<T�a<=�`<�_<�~_<�y_<�_<�`<�b`<U�`<�i`<5`<'�_<1_<{_<f�_<�  �  ��a<M�b<d�c<q�d<D�d<�ed<Roc<b<LK`<�~^<��\<�R[<�2Z<�Y<�OY<[�Y<�jZ<�[<�)]<Z�^<1�`<�_b<�c<ӏd<N�d<'�d<��c<W�b<�ta<�g`<|�_<e_<��^<ޛ^<j�^<Ґ^<̖^<��^<�^<�Y_<�`<�a<�'b<fQc<�Fd<�d<�d<�@d<.c<\�a<��_<^<�h\<y[<�Z<�Y<��Y<��Y<H�Z<�G\<��]<��_<swa<�c<s>d<�d<�d<{d<7�c<�lb<�Da<�I`<g�_<�_<H�^<��^<��^<�^<�^<��^<�+_<*�_<@u`<a|a<�b<��c<��d<��d<��d<>d<+�b<�a<jI_<;�]<�[<��Z<�Y<��Y<�Y<�MZ<Ib[<��\<р^<lL`<Ib<�c<��d<�d<��d<�2d<�.c<b</�`<��_<a__< �^<��^<
�^<��^<	�^<��^<��^<�P_<��_<<�`<+�a<�c<�d<;�d<{�d<��d<�c<�3b<�|`<>�^<�\<�[<dZ<�Y<
�Y<�Y<ʙZ<��[<OV]<�_<6�`<[�b<��c<0�d<��d<˧d<��c<�b<p�a<'�`<��_< 2_<F�^<��^<�^<+�^<��^<6�^<v_<z_<q*`<�a<�Cb< kc<P^d<��d<B�d<JQd<p-c<�a<��_<t^<Rl\<t[<�Z<`�Y<�|Y<��Y<��Z<h8\<��]<Y�_<I`a<�b<m"d<��d<��d<�Xd<�lc<mFb<9a<� `<:g_<��^<��^<g�^<�^<�^<��^<��^<��^<��_<J`<gQa< }b<��c<Hod<��d<��d<��c<݈b<��`<�_<�W]<��[<A�Z<��Y<�PY<
uY<�Z<�,[<d�\<�K^<*`<
�a<�Jc<+Pd<?�d<p�d<�c<H�b<��a<�`<$�_<�$_< �^<;�^<��^<7}^<�^<��^<L�^<._<�_<��`<�  �  �4b<�c<އd<5e<be<}d<'vc<L"b<��`<�V_<M)^<�8]<��\<�)\<�\<�:\<��\<2j]<�i^<�_<;a<=vb<c�c<&�d<q#e<�e<�ad<MKc<<�a<��`<�,_<5	^<�$]<ۅ\<�.\<�\<9X\<��\<y�]<�^<y�_<qWa<��b<C d<��d<O<e<)	e<UNd<c)c<L�a<�\`<�_<o�]<�]<��\<P@\<�=\<�\<]<��]<�^<%E`<Ʊa<%c<�Id<�e<2Ze<�e<=?d<c<�a<;`</�^<��]<�]<�\<�K\<�R\<��\<V8]< ^<�1_<˂`<~�a<.Oc<pd<�$e</Qe<9�d<�	d<;�b<<_a<[�_<_�^<�]<��\<vw\<D\<�W\<�\<[W]<.@^<fg_<ۿ`<D.b<m�c<B�d<79e<�Me<��d<'�c<Ӓb<y%a<��_<��^<��]<��\<;l\<�D\<�c\<|�\<Rz]<�m^<��_<��`<�ib<M�c<C�d<�De<�@e<��d<اc<�Sb<P�`<��_< [^<�j]<h�\<Z[\<�?\<�j\<�\<��]<ʖ^<��_<�2a<f�b<F�c<��d<)Ie<�,e<��d<$oc<�b<	�`<9P_<�,^<:H]<b�\<�Q\<�B\<�z\<��\<��]<��^<#`<�ta<h�b<�d<S�d<�Qe<2e<�^d<�7c<��a<�e`<�_<�]<�]<��\<�;\<�6\<y\<h]<��]<"�^<�0`<��a<��b<�-d<s�d<�9e<T�d<�d< �b<u}a<1`<>�^<�]<q�\<�_\<\\<b&\<�u\<]]<M�]<V_<�W`<y�a<+$c<�Dd<f�d<%e<m�d<#�c<��b<s/a<u�_<d�^<	�]<Ⱦ\<�B\<\<L"\<@~\<�!]<�
^<�1_<s�`<��a<Rc<�cd<�e<we<�d<�c<�Zb<��`<��_<�S^<2X]<�\<V1\<�	\<�)\<��\<8A]<�5^<�f_<��`<�  �   b<Tc<�nd<�d<Ǒd<�c<�b<��a<��`<3�_<x_<�^<ԑ^<Ѓ^<��^<�^<K�^<��^<E2_<��_<��`<(�a<}c<�d<O�d<��d<�Od<PCc<A�a<�	`<-?^<[�\<�([<�Z<�~Y<kbY<>�Y<v�Z<��[<�]<pE_<�a<�b<j�c<��d<�d<�|d<!�c<�b<�Ya<V`<B�_<�_<��^<5�^<�^<�^<��^<��^<_<��_<WL`<�La<Gwb<�c<�d<��d<\�d<�4d<�b<gfa<d�_<�]<�>\<O�Z<Z<�Y<�Y<],Z<�.[<��\<�5^<_�_<�a<�Ec<ad<W�d<E�d<DSd<.[c<2b<6a<c`<Sr_<�_<N�^<�^<�^<O�^<|�^<��^<�<_<�_<��`<�a<G�b<S�c<�d<< e<M�d<��c<�yb<�`< _<yE]<��[<��Z<��Y<��Y<e�Y<�uZ<��[<`]<r�^<��`<Lb<X�c<�d<��d<��d<�	d<��b<��a<��`<I�_<�F_<Q�^<�^<��^<-�^<��^<A�^<��^<�__</`<��`<�b<�7c< 8d<W�d<��d<td<Jgc<��a<!-`<�b^<Ƕ\<KL[<.>Z<�Y<L�Y<��Y</�Z<\\<��]<�c_<�-a<I�b<�d<��d<G�d<x�d<��c<��b<*ea<�^`<��_<._<��^<i�^<~�^<ԣ^<��^<;�^<�_<�|_<�7`<z5a<�]b<A�c<ed<��d<"�d<vd<F�b<?a<�u_<W�]<\<	�Z<I�Y<dY<�qY<\ Z<�[<&d\<>
^<6�_<�a<�c<�5d<��d<�d<)&d<#-c<�b<��`<	�_<�?_<	�^<��^<�^<�^<l�^<s�^<��^<_<_�_<i`<�ya<�b<�c<a�d<X�d<�~d<�c<Bb<ܓ`<&�^<�]<��[<SWZ<��Y<{JY<�Y<_<Z<�a[<��\<��^<�b`<�  �  ia<��b<�c<�c<Ymc<x�b<�a<w�`<��_<z{_<}�_<L�_<�&`<�p`<}�`<kd`<`<
�_<8~_<)�_<��_<.�`<��a<��b<Ϙc<^�c<#�c<,�b<�a<5_<|�\<
�Z<�X<�W<�V<�V<�W<�HX<K�Y<�\<J.^<�E`<ab<?Lc<]�c<��c<xIc<�Ub<@Fa<~\`<Z�_<�_<��_<�`<j`<̦`<��`<w`<f `<��_< �_<|�_<tY`<>a<�Nb<�Kc<��c<�d<��c<�Xb<E�`<S�^<qe\<WZ<��X<�[W<һV<y�V<ȓW<��X<K�Z<��\<_<�a<�b<^�c<d<��c<�c<�b<a<�2`<�_<Ϭ_<��_<�=`<��`<|�`<��`<|f`<�
`<Z�_<��_<��_<��`< �a<��b<?�c<�	d<��c<n.c<B�a<'�_<��]<��[<��Y<�X<�W<k�V<~�V<�W<��Y<�o[<`�]<0�_<��a<tc<2�c<�d<��c<x�b<�a<~�`< `<ݭ_<�_<��_<xY`<�`<w�`<��`<�D`<u�_<k�_<�_<3`<8�`<q�a<.�b<!�c<�d<˼c<H�b<T5a<�<_<�]<a�Z<]Y<2�W<�V<ǮV<;W<jX<�Z<Y!\<}L^<�b`<g&b<lec<�d<��c<B\c<fb<<Ta<�g`<<�_<_�_<��_<�`<Eh`<E�`<S�`<#m`<�`<>�_<�_<�_<{B`<�$a<3b<�-c<n�c<��c<�bc<�2b<-z`<�h^<�;\<�,Z<�oX<0W<	�V<��V<�gW<5�X<˖Z<��\<��^<��`<�vb<�c<&�c< �c<:�b<^�a<��`<`<W�_<�y_<��_<�`<;\`<��`<hu`<0`<��_<*�_<�w_<̾_<:i`<�aa<=rb<�Wc<5�c<��c<��b<	�a<L�_<z�]<zr[<?zY<��W<��V<�qV<�V<#�W<fHY<D8[<�]]<��_<�  �  [d`<|�a<��b<i�b<��a<�`<��_<i_<O�^<��^<?�_<�o`<Ja<�a</b<��a<ja<�>`<ni_<��^<D�^<Y<_<�`<�.a<b<2�b<�zb<e�a<�`<��]<�{[<dY<��V<uU<"T<��S<�T<	�U<�X<�fZ<�\<�/_<t	a<]=b<�b<hyb<ֵa<�`<Ȱ_<�_<��^<�>_<k�_<E�`<έa<�(b<�0b<z�a<�a<`<�\_<y�^<}_<*�_<ݦ`<:�a<t�b<��b<ktb<�Va<"�_<�M]<��Z<[jX<�VV<P�T<�T<P)T<3U<"�V<:�X<�\[<o�]<��_<}�a<�b<��b<^[b<ywa<�h`<�~_<��^<�_<;�_<RX`<4;a<��a<~Fb<�$b<[�a<9�`<��_<;3_<J�^<%8_<��_<~a<�b<j�b<"�b<�$b<��`<��^<+x\<!�Y<��W<;�U<SyT<��S<�`T<�U<�kW<G�Y<21\<�^<͘`<(b<��b<�b<�b<a<�`<�E_<��^<g#_<�_<ۢ`<}a<�b<�Eb<T�a<VOa<gn`<�_<�
_<�^<�f_<�G`<\Va<�Bb<��b<m�b<��a<�,`<T^<��[<�(Y<�V<�:U<�3T<IT<�T<QV<�"X<ӅZ<�]<�L_<P$a<dVb<��b<T�b<��a<C�`<��_<�_<��^<!E_<��_<%�`<��a<)$b<�)b<��a<��`<�`<�J_<�^<��^<Փ_<3�`<V�a<veb<��b<�Pb<.1a<3h_<�%]<~�Z<+@X<,V<��T<P�S<��S<��T<��V<ϾX<x1[<G�]<j�_<2ta<hb<��b<�.b<�Ia<:`<O_<��^<^�^<�S_<$`<a<غa<&b<O�a<�^a<��`<8�_<�^<t�^<�_<��_<3�`<~�a<�wb<9�b<j�a<��`<h�^<@\<~�Y<~oW<�U<�?T<K�S<�'T<eZU<�3W<<Y<�[<�^^<�  �  Y_<Ӿ`<-Va<U'a<�``<�L_<�F^<�]<a�]<�E^<�h_<��`<�b<\�b<5#c<D�b<L�a<sx`<�"_<�^<�]<��]<��^<%�_<b�`<	Ja<�Pa<��`<�^<��\<�)Z<RtW<��T<�	S<j�Q<n�Q<#kR<#T<dSV<�X<�[<�^<�_<�!a<ua<�a<%`<a_<	 ^<��]<!�]<f�^<�_<\a<`�b<�1c<�<c<�b< �a</`<��^<	^<�]<� ^<~_<i `<)a<O�a<nUa<}J`<�}^<;\<nY<q�V<�mT<��R<>�Q<�Q<
S<��T<�QW<FZ<:�\<��^<i�`<na<�}a<:�`<��_<T�^<��]<��]<�2^<v2_<��`<��a<��b<�Uc<'c<�Zb<(!a<��_<k�^<��]<�]<0b^<�`_<�w`<CKa<2�a<�a<`�_<��]<�7[<�X<0�U<R�S<jPR<�Q<�4R<�S<ۥU<�3X<9�Z<�w]<X�_<`�`<�a<�Ya<Ԓ`<�~_<�x^<[�]<��]<�x^<ڛ_<��`<?9b<zc<�Uc<a�b<��a<��`<�Q_<mE^<-�]<�]<�^<�_<(�`<�oa<�ua<
�`<�_<?�\<�LZ<��W<�U<�,S<R<��Q<��R<C-T<�sV<?Y<��[<�8^<�`<�:a< �a<�"a<�7`<�_<�-^<޼]<��]<��^<�`<�\a<��b<8-c<c5c<��b<�{a<�`<��^<��]<>�]<\^<��^<�`<?�`<ona<�1a<&%`<�V^<%�[<�DY<f�V<�BT<Q�R<ƭQ<��Q<s�R<U�T<0&W<�Y<}\<��^<f`<kBa<_Qa<E�`<��_<p�^<w�]<��]<s ^<��^<%P`<9�a<Y�b<Sc<"�b<�#b<R�`<7�_<$`^<ҫ]<q�]<�,^<�+_<�B`<�a<qXa<P�`<��_<��]< [<�HX<r�U<Q�S<RR<�Q<��Q<�WS<OnU<,�W<F�Z<�B]<�  �  \�^<��_<^t`<�'`<}C_<�^<�]<r�\<��\<_�]<8_<�`<zlb<�qc<��c<�Fc<�b<s�`<��^<�|]<��\<<�\<�P]<-f^<\�_<mQ`<�t`<��_<9^<5�[<c@Y<�eV<��S<Y�Q<�gP<;+P<�P<��R<J2U<jX<r�Z<zV]<K:_<P`<ω`<�`<? _<��]<��\<�\<+]<�R^<j�_<a�a<�b<��c<|�c<�c< �a<�%`<��^<nS]<��\<h�\<��]<J�^<�`<¡`<e�`<�_<��]<EG[<FyX<�U<q&S<@NQ<�]P<�{P<2�Q<ѥS<�>V<XY<r�[<Y)^<��_<�`<��`<��_<v�^<��]<�\<��\<�]<��^<��`<m+b<Bcc<F�c<��c<��b<CMa<��_<�^<3]<��\<06]<0^<�W_<H`<2�`<A`<V�^<�\<�XZ<�W<1�T<]oR<��P<�FP<��P<8R<vT<9.W<�Z<R�\<��^<�&`<C�`<.Z`<�u_<!O^<K]<��\<{�\<\�]<�k_<}a<�b<(�c<��c<)yc<@Qb<ߺ`<
_<��]<�\<�\<z]<F�^<B�_<Kw`<��`<�_<]^<�\<�cY<�V<��S<9�Q<P�P<{MP<� Q<��R<mRU<w X<7�Z<�r]<�T_<�h`<��`<�`<�_<��]<�]<i�\<�3]<Y^<��_<:�a<A�b<U�c<>�c<�c<��a<�`<)w^<?]<ְ\<'�\<H�]<��^<�_<�`<�]`<�`_<��]<D[<1PX<#|U<��R<)#Q<]2P<6PP<�wQ<azS<5V<#�X<K�[<$�]<s�_<Si`<7\`<x�_<}�^<�i]<ݰ\<T�\<T\]<�^</Y`<��a<�,c<x�c<{�c<k�b<La<�f_<*�]<3�\<ߐ\<� ]<��]<�"_<�`<�s`<	`<��^<�\<7!Z<�GW<��T<�6R<�P<P<9�P< R<�>T<��V<+�Y<Wx\<�  �  �O^<��_<�!`<,�_<�^<�]<b�\<j0\<z\<܉]<$_<��`<ʌb<Рc<s�c<Gsc<};b<K�`<��^<=B]<\\<<@\<<�\<�]<&!_<��_<�$`<
{_<j�]<�[<��X<�V<TS<�.Q<U�O<�O<G~P< MR<��T<��W<�Z<�]<H�^<�`<�3`<��_<��^<k]<��\<�R\<K�\<3*^<b�_<��a<G"c<��c<�d<�Gc<j�a<`<�c^<�]<Zj\<��\<d]<,�^<R�_<�J`< 4`<�>_<Bq]<��Z</#X<'BU<O�R<��P<��O<��O<`&Q<�6S<��U<��X<s�[<w�]<��_<�E`</`<�i_<�E^<)]<�w\<�~\<-Q]<K�^<͍`<�Db<`�c<�%d<��c<��b<)Ya<��_<��]<�\<:c\<Y�\<��]<J�^<5�_<�U`<e�_<��^<y�\<�	Z<J%W<bVT<x�Q<�[P<	�O<�<P<��Q<�T<S�V<��Y<=d\<��^<�_<�T`<��_<H_<�]<��\<�b\<8�\<�]<eW_<o$a<S�b<2�c<u&d<��c<mb<ɽ`<��^<p]<��\<+k\<�
]<* ^<H_<�`<�I`<m�_<P^<v�[<GY<	*V<wS<�QQ<�P<�O<��P<�mR<��T<��W<ڥZ<+]<�_<�`<�J`<Z�_<��^<B{]<[�\<�]\<�\<\0^<��_<Ѫa<o c<�c<�d<�=c<��a<�`<�Q^<��\<�S\<�w\<wH]<io^<y�_<�(`<�`<Y_<�J]<��Z<"�W<<U<��R<��P<l�O<9�O<��P<QS<��U<��X<La[<@�]<MW_<4`<�`<q<_<�^<�\<�G\<nM\<]<v�^<�X`<b<�Wc<��c<t�c<вb<&"a<�U_<G�]<�\<�-\<��\<a�]<�^<ܳ_< `<_�_<-^<kr\<�Y<5�V<�T<��Q<�"P<T�O<BP<��Q<f�S<V<��Y<M/\<�  �  \�^<��_<^t`<�'`<}C_<�^<�]<r�\<��\<_�]<8_<�`<zlb<�qc<��c<�Fc<�b<s�`<��^<�|]<��\<<�\<�P]<-f^<\�_<mQ`<�t`<��_<9^<5�[<c@Y<�eV<��S<Y�Q<�gP<;+P<�P<��R<J2U<jX<r�Z<zV]<K:_<P`<ω`<�`<? _<��]<��\<�\<+]<�R^<j�_<a�a<�b<��c<|�c<�c< �a<�%`<��^<nS]<��\<h�\<��]<J�^<�`<¡`<e�`<�_<��]<EG[<FyX<�U<q&S<@NQ<�]P<�{P<2�Q<ѥS<�>V<XY<r�[<Y)^<��_<�`<��`<��_<v�^<��]<�\<��\<�]<��^<��`<m+b<Bcc<F�c<��c<��b<CMa<��_<�^<3]<��\<06]<0^<�W_<H`<2�`<A`<V�^<�\<�XZ<�W<1�T<]oR<��P<�FP<��P<8R<vT<9.W<�Z<R�\<��^<�&`<C�`<.Z`<�u_<!O^<K]<��\<{�\<\�]<�k_<}a<�b<(�c<��c<)yc<@Qb<ߺ`<
_<��]<�\<�\<z]<F�^<B�_<Kw`<��`<�_<]^<�\<�cY<�V<��S<9�Q<P�P<{MP<� Q<��R<mRU<w X<7�Z<�r]<�T_<�h`<��`<�`<�_<��]<�]<i�\<�3]<Y^<��_<:�a<A�b<U�c<>�c<�c<��a<�`<)w^<?]<ְ\<'�\<H�]<��^<�_<�`<�]`<�`_<��]<D[<1PX<#|U<��R<)#Q<]2P<6PP<�wQ<azS<5V<#�X<K�[<$�]<s�_<Si`<7\`<x�_<}�^<�i]<ݰ\<T�\<T\]<�^</Y`<��a<�,c<x�c<{�c<k�b<La<�f_<*�]<3�\<ߐ\<� ]<��]<�"_<�`<�s`<	`<��^<�\<7!Z<�GW<��T<�6R<�P<P<9�P< R<�>T<��V<+�Y<Wx\<�  �  Y_<Ӿ`<-Va<U'a<�``<�L_<�F^<�]<a�]<�E^<�h_<��`<�b<\�b<5#c<D�b<L�a<sx`<�"_<�^<�]<��]<��^<%�_<b�`<	Ja<�Pa<��`<�^<��\<�)Z<RtW<��T<�	S<j�Q<n�Q<#kR<#T<dSV<�X<�[<�^<�_<�!a<ua<�a<%`<a_<	 ^<��]<!�]<f�^<�_<\a<`�b<�1c<�<c<�b< �a</`<��^<	^<�]<� ^<~_<i `<)a<O�a<nUa<}J`<�}^<;\<nY<q�V<�mT<��R<>�Q<�Q<
S<��T<�QW<FZ<:�\<��^<i�`<na<�}a<:�`<��_<T�^<��]<��]<�2^<v2_<��`<��a<��b<�Uc<'c<�Zb<(!a<��_<k�^<��]<�]<0b^<�`_<�w`<CKa<2�a<�a<`�_<��]<�7[<�X<0�U<R�S<jPR<�Q<�4R<�S<ۥU<�3X<9�Z<�w]<X�_<`�`<�a<�Ya<Ԓ`<�~_<�x^<[�]<��]<�x^<ڛ_<��`<?9b<zc<�Uc<a�b<��a<��`<�Q_<mE^<-�]<�]<�^<�_<(�`<�oa<�ua<
�`<�_<?�\<�LZ<��W<�U<�,S<R<��Q<��R<C-T<�sV<?Y<��[<�8^<�`<�:a< �a<�"a<�7`<�_<�-^<޼]<��]<��^<�`<�\a<��b<8-c<c5c<��b<�{a<�`<��^<��]<>�]<\^<��^<�`<?�`<ona<�1a<&%`<�V^<%�[<�DY<f�V<�BT<Q�R<ƭQ<��Q<s�R<U�T<0&W<�Y<}\<��^<f`<kBa<_Qa<E�`<��_<p�^<w�]<��]<s ^<��^<%P`<9�a<Y�b<Sc<"�b<�#b<R�`<7�_<$`^<ҫ]<q�]<�,^<�+_<�B`<�a<qXa<P�`<��_<��]< [<�HX<r�U<Q�S<RR<�Q<��Q<�WS<OnU<,�W<F�Z<�B]<�  �  [d`<|�a<��b<i�b<��a<�`<��_<i_<O�^<��^<?�_<�o`<Ja<�a</b<��a<ja<�>`<ni_<��^<D�^<Y<_<�`<�.a<b<2�b<�zb<e�a<�`<��]<�{[<dY<��V<uU<"T<��S<�T<	�U<�X<�fZ<�\<�/_<t	a<]=b<�b<hyb<ֵa<�`<Ȱ_<�_<��^<�>_<k�_<E�`<έa<�(b<�0b<z�a<�a<`<�\_<y�^<}_<*�_<ݦ`<:�a<t�b<��b<ktb<�Va<"�_<�M]<��Z<[jX<�VV<P�T<�T<P)T<3U<"�V<:�X<�\[<o�]<��_<}�a<�b<��b<^[b<ywa<�h`<�~_<��^<�_<;�_<RX`<4;a<��a<~Fb<�$b<[�a<9�`<��_<;3_<J�^<%8_<��_<~a<�b<j�b<"�b<�$b<��`<��^<+x\<!�Y<��W<;�U<SyT<��S<�`T<�U<�kW<G�Y<21\<�^<͘`<(b<��b<�b<�b<a<�`<�E_<��^<g#_<�_<ۢ`<}a<�b<�Eb<T�a<VOa<gn`<�_<�
_<�^<�f_<�G`<\Va<�Bb<��b<m�b<��a<�,`<T^<��[<�(Y<�V<�:U<�3T<IT<�T<QV<�"X<ӅZ<�]<�L_<P$a<dVb<��b<T�b<��a<C�`<��_<�_<��^<!E_<��_<%�`<��a<)$b<�)b<��a<��`<�`<�J_<�^<��^<Փ_<3�`<V�a<veb<��b<�Pb<.1a<3h_<�%]<~�Z<+@X<,V<��T<P�S<��S<��T<��V<ϾX<x1[<G�]<j�_<2ta<hb<��b<�.b<�Ia<:`<O_<��^<^�^<�S_<$`<a<غa<&b<O�a<�^a<��`<8�_<�^<t�^<�_<��_<3�`<~�a<�wb<9�b<j�a<��`<h�^<@\<~�Y<~oW<�U<�?T<K�S<�'T<eZU<�3W<<Y<�[<�^^<�  �  ia<��b<�c<�c<Ymc<x�b<�a<w�`<��_<z{_<}�_<L�_<�&`<�p`<}�`<kd`<`<
�_<8~_<)�_<��_<.�`<��a<��b<Ϙc<^�c<#�c<,�b<�a<5_<|�\<
�Z<�X<�W<�V<�V<�W<�HX<K�Y<�\<J.^<�E`<ab<?Lc<]�c<��c<xIc<�Ub<@Fa<~\`<Z�_<�_<��_<�`<j`<̦`<��`<w`<f `<��_< �_<|�_<tY`<>a<�Nb<�Kc<��c<�d<��c<�Xb<E�`<S�^<qe\<WZ<��X<�[W<һV<y�V<ȓW<��X<K�Z<��\<_<�a<�b<^�c<d<��c<�c<�b<a<�2`<�_<Ϭ_<��_<�=`<��`<|�`<��`<|f`<�
`<Z�_<��_<��_<��`< �a<��b<?�c<�	d<��c<n.c<B�a<'�_<��]<��[<��Y<�X<�W<k�V<~�V<�W<��Y<�o[<`�]<0�_<��a<tc<2�c<�d<��c<x�b<�a<~�`< `<ݭ_<�_<��_<xY`<�`<w�`<��`<�D`<u�_<k�_<�_<3`<8�`<q�a<.�b<!�c<�d<˼c<H�b<T5a<�<_<�]<a�Z<]Y<2�W<�V<ǮV<;W<jX<�Z<Y!\<}L^<�b`<g&b<lec<�d<��c<B\c<fb<<Ta<�g`<<�_<_�_<��_<�`<Eh`<E�`<S�`<#m`<�`<>�_<�_<�_<{B`<�$a<3b<�-c<n�c<��c<�bc<�2b<-z`<�h^<�;\<�,Z<�oX<0W<	�V<��V<�gW<5�X<˖Z<��\<��^<��`<�vb<�c<&�c< �c<:�b<^�a<��`<`<W�_<�y_<��_<�`<;\`<��`<hu`<0`<��_<*�_<�w_<̾_<:i`<�aa<=rb<�Wc<5�c<��c<��b<	�a<L�_<z�]<zr[<?zY<��W<��V<�qV<�V<#�W<fHY<D8[<�]]<��_<�  �   b<Tc<�nd<�d<Ǒd<�c<�b<��a<��`<3�_<x_<�^<ԑ^<Ѓ^<��^<�^<K�^<��^<E2_<��_<��`<(�a<}c<�d<O�d<��d<�Od<PCc<A�a<�	`<-?^<[�\<�([<�Z<�~Y<kbY<>�Y<v�Z<��[<�]<pE_<�a<�b<j�c<��d<�d<�|d<!�c<�b<�Ya<V`<B�_<�_<��^<5�^<�^<�^<��^<��^<_<��_<WL`<�La<Gwb<�c<�d<��d<\�d<�4d<�b<gfa<d�_<�]<�>\<O�Z<Z<�Y<�Y<],Z<�.[<��\<�5^<_�_<�a<�Ec<ad<W�d<E�d<DSd<.[c<2b<6a<c`<Sr_<�_<N�^<�^<�^<O�^<|�^<��^<�<_<�_<��`<�a<G�b<S�c<�d<< e<M�d<��c<�yb<�`< _<yE]<��[<��Z<��Y<��Y<e�Y<�uZ<��[<`]<r�^<��`<Lb<X�c<�d<��d<��d<�	d<��b<��a<��`<I�_<�F_<Q�^<�^<��^<-�^<��^<A�^<��^<�__</`<��`<�b<�7c< 8d<W�d<��d<td<Jgc<��a<!-`<�b^<Ƕ\<KL[<.>Z<�Y<L�Y<��Y</�Z<\\<��]<�c_<�-a<I�b<�d<��d<G�d<x�d<��c<��b<*ea<�^`<��_<._<��^<i�^<~�^<ԣ^<��^<;�^<�_<�|_<�7`<z5a<�]b<A�c<ed<��d<"�d<vd<F�b<?a<�u_<W�]<\<	�Z<I�Y<dY<�qY<\ Z<�[<&d\<>
^<6�_<�a<�c<�5d<��d<�d<)&d<#-c<�b<��`<	�_<�?_<	�^<��^<�^<�^<l�^<s�^<��^<_<_�_<i`<�ya<�b<�c<a�d<X�d<�~d<�c<Bb<ܓ`<&�^<�]<��[<SWZ<��Y<{JY<�Y<_<Z<�a[<��\<��^<�b`<�  �  �4b<�c<އd<5e<be<}d<'vc<L"b<��`<�V_<M)^<�8]<��\<�)\<�\<�:\<��\<2j]<�i^<�_<;a<=vb<c�c<&�d<q#e<�e<�ad<MKc<<�a<��`<�,_<5	^<�$]<ۅ\<�.\<�\<9X\<��\<y�]<�^<y�_<qWa<��b<C d<��d<O<e<)	e<UNd<c)c<L�a<�\`<�_<o�]<�]<��\<P@\<�=\<�\<]<��]<�^<%E`<Ʊa<%c<�Id<�e<2Ze<�e<=?d<c<�a<;`</�^<��]<�]<�\<�K\<�R\<��\<V8]< ^<�1_<˂`<~�a<.Oc<pd<�$e</Qe<9�d<�	d<;�b<<_a<[�_<_�^<�]<��\<vw\<D\<�W\<�\<[W]<.@^<fg_<ۿ`<D.b<m�c<B�d<79e<�Me<��d<'�c<Ӓb<y%a<��_<��^<��]<��\<;l\<�D\<�c\<|�\<Rz]<�m^<��_<��`<�ib<M�c<C�d<�De<�@e<��d<اc<�Sb<P�`<��_< [^<�j]<h�\<Z[\<�?\<�j\<�\<��]<ʖ^<��_<�2a<f�b<F�c<��d<)Ie<�,e<��d<$oc<�b<	�`<9P_<�,^<:H]<b�\<�Q\<�B\<�z\<��\<��]<��^<#`<�ta<h�b<�d<S�d<�Qe<2e<�^d<�7c<��a<�e`<�_<�]<�]<��\<�;\<�6\<y\<h]<��]<"�^<�0`<��a<��b<�-d<s�d<�9e<T�d<�d< �b<u}a<1`<>�^<�]<q�\<�_\<\\<b&\<�u\<]]<M�]<V_<�W`<y�a<+$c<�Dd<f�d<%e<m�d<#�c<��b<s/a<u�_<d�^<	�]<Ⱦ\<�B\<\<L"\<@~\<�!]<�
^<�1_<s�`<��a<Rc<�cd<�e<we<�d<�c<�Zb<��`<��_<�S^<2X]<�\<V1\<�	\<�)\<��\<8A]<�5^<�f_<��`<�  �  ��a<M�b<d�c<q�d<D�d<�ed<Roc<b<LK`<�~^<��\<�R[<�2Z<�Y<�OY<[�Y<�jZ<�[<�)]<Z�^<1�`<�_b<�c<ӏd<N�d<'�d<��c<W�b<�ta<�g`<|�_<e_<��^<ޛ^<j�^<Ґ^<̖^<��^<�^<�Y_<�`<�a<�'b<fQc<�Fd<�d<�d<�@d<.c<\�a<��_<^<�h\<y[<�Z<�Y<��Y<��Y<H�Z<�G\<��]<��_<swa<�c<s>d<�d<�d<{d<7�c<�lb<�Da<�I`<g�_<�_<H�^<��^<��^<�^<�^<��^<�+_<*�_<@u`<a|a<�b<��c<��d<��d<��d<>d<+�b<�a<jI_<;�]<�[<��Z<�Y<��Y<�Y<�MZ<Ib[<��\<р^<lL`<Ib<�c<��d<�d<��d<�2d<�.c<b</�`<��_<a__< �^<��^<
�^<��^<	�^<��^<��^<�P_<��_<<�`<+�a<�c<�d<;�d<{�d<��d<�c<�3b<�|`<>�^<�\<�[<dZ<�Y<
�Y<�Y<ʙZ<��[<OV]<�_<6�`<[�b<��c<0�d<��d<˧d<��c<�b<p�a<'�`<��_< 2_<F�^<��^<�^<+�^<��^<6�^<v_<z_<q*`<�a<�Cb< kc<P^d<��d<B�d<JQd<p-c<�a<��_<t^<Rl\<t[<�Z<`�Y<�|Y<��Y<��Z<h8\<��]<Y�_<I`a<�b<m"d<��d<��d<�Xd<�lc<mFb<9a<� `<:g_<��^<��^<g�^<�^<�^<��^<��^<��^<��_<J`<gQa< }b<��c<Hod<��d<��d<��c<݈b<��`<�_<�W]<��[<A�Z<��Y<�PY<
uY<�Z<�,[<d�\<�K^<*`<
�a<�Jc<+Pd<?�d<p�d<�c<H�b<��a<�`<$�_<�$_< �^<;�^<��^<7}^<�^<��^<L�^<._<�_<��`<�  �  ��`<>�a<�b<�vc<<�c<l�c</�b<\Ra<Ug_<~A]<�[<�2Y<ܰW<�V<7wV<d�V<~�W<ؙY<��[<:�]<=�_<�a<$c<%�c<&�c<Wc<�mb<�]a<i`<g�_<=�_<��_<��_<�C`<&�`<u�`<�h`<�`<D�_<��_<�_<�`<��`<Wb<v	c<#�c<m�c<N�c<{b<��`<v�^<W�\<��Z<5�X<0tW<�V<)�V<c[W<��X<�fZ<�y\<-�^<m�`<hb<`�c<�d<�c<�Ac<!Db<6a<kW`<��_<�_<a�_<�3`<T�`<ټ`<U�`<�v`<`<�_<M�_<7�_<z`<
ha<nxb<�ic<@�c<�c<�Vc<5b<ME`<�,^<j\<�Y<�UX<�/W<�V<#�V<�W<&6Y<�[<�7]< `_<�Ta<��b<P�c<d<��c<��b<1�a<��`<�`<�_<Ѵ_<`�_<�O`<�`<&�`<�`<Y`<)�_<9�_<��_<4
`<L�`<��a<��b<��c<ud<-�c<��b<��a<��_<�r]<�N[<�cY<��W<��V<'�V<�W<�*X<%�Y<��[<�]<�`<6�a<=6c<,�c<E�c<{{c<�b<a�a<~�`<��_<ʦ_<I�_<m`<ug`<�`<�`<�`<G7`<��_<u�_<�_<}<`<qa<@b<K!c<��c<�d<)�c<]�b<^�`<��^<ʰ\<v�Z<6�X<rrW<e�V<�V<eQW<�X<~WZ<�g\<��^<3�`<MNb<Csc<��c<��c<4c<�b<�a<�/`<l�_<��_<�_<�`<�]`<2�`<��`<�I`<��_<#�_<�~_<�_<,O`<8=a<�Mb<h>c<��c<��c<�)c<D�a<V`<��]<X�[< �Y<#X<J�V<�yV<|�V<3�W<Y<��Z<�]<+_<xa<E�b<��c<'�c<,�c<p�b<T�a<=�`<�_<�~_<�y_<�_<�`<�b`<U�`<�i`<5`<'�_<1_<{_<f�_<�  �  l_<��_<��`<|�a<��b<6�b<�a<�L`<�@^<8�[<�_Y<BW<RHU<� T<��S<�QT<��U<�W<��Y<�i\<��^<'�`<�b<@�b<�zb<��a<W�`<O�_<�_<��^<_<L�_<U�`<�wa<�b<Ub<j�a<#a<)`<k\_<W�^<�^<n_<u]`<vma<1Nb<��b<�vb<�xa<��_<��]<m'[<��X<�V<m�T<�T<pT<M�T<ddV<X<4�Z<ig]<T�_<@fa<�{b<��b<�}b<�a<��`<�_<�_<H_<jq_<�8`<*a<��a<�Cb<p5b<J�a<�`<�`<�H_<��^<9!_<N�_<��`<��a<A�b<��b<0Ib<�a<�,_<��\<�aZ<�X<�V< �T<� T<�?T<�QU<�W<OY<\�[<�3^<M`<�a<��b<9�b<�>b<oNa<�@`<"d_<��^<�_<�_<x�`<�`a<	b<�Kb<�b<�va<<�`<��_<� _<��^<QP_<x"`<S.a<h%b<��b<�b<b�a<�}`<�q^<\<z�Y<�IW<�xU<�PT<a�S<��T<x�U<��W<LZ<F�\<��^<�`<I+b<��b<ٟb<��a<�`<��_<>*_<E�^<�4_<�_<D�`<��a<�&b<Bb<��a<�-a<�J`<}_<�_<�_<�_<�w`<m�a<�cb<��b<ȇb<*�a<��_<��]<�-[<X�X<�V<��T<	T<0 T<M�T<�WV<pX<�Z<�R]<�_<yLa<y_b<2�b<�\b<D�a<�w`<��_<��^<��^<�F_<`<��`<�a<�b<�b<��a<��`<��_< _<\�^<P�^<��_<�`<��a<�jb<�b<vb<$�`<Y�^<��\<(1Z<F�W<U�U<�lT<��S<NT<>U<��V<)Y<k�[<��]<�`<Ρa<wb<+�b<�b<a<|`<)+_<��^<�^<�m_<�E`<�$a<��a<Ib<��a<~;a<�_`<Q�_<B�^<x�^<�  �  ��]<%R^<!\_<nn`<�.a<Ta<��`<DA_<#]<��Z<��W<+PU<�BS<W�Q<̐Q<&+R<�S<��U<wuX<�,[<�]<�_<�`<;ba<}a<�=`<R&_<,^<��]<�]<{^<��_<�a<dAb<yc<�,c<��b<ڢa<2N`< _<�^<Ф]<X�]<4�^<��_<�`<�ka<�Ra<<k`<.�^<$r\<��Y<.W<(�T<��R<n�Q<��Q<�R<�~T<��V<�Y<y9\<�^<�Y`<$[a<ތa<(a<�`<��^<^<I�]<b^<�_<�O`<��a<�b<�Pc<=c<ևb<�Za<��_<
�^<��]<��]<�=^</_<TH`<�,a<�a<�.a<Q`<^<c�[<��X<�OV<nT<�|R<��Q<�R<�FS<�AU<��W<^xZ<\]<�@_<��`<��a<�pa<پ`<�_<O�^<��]<��]<�W^<$j_<��`<Eb<��b<!\c<c< .b<��`<3�_<o^<Q�]<��]<�^< �_<h�`<&aa<��a<��`<Br_<�S]<3�Z<z
X<��U<�rS<#R<��Q<�YR<��S<MV<נX<�V[<b�]<��_<�a<��a<-;a<�a`<�I_<{O^<��]<x�]<��^<]�_<�/a<�eb<�*c<�Pc<#�b<��a<)p`<� _<u(^<��]<z^<a�^<��_<��`<Ia<�ca<�y`<�^<\{\<C�Y<�W<4�T<(�R<��Q<]�Q<�R<�qT<�V<�xY<�$\<�}^<@`<�>a<Jna<\�`<�_<��^<w�]<�]<��]<�^<6$`<j|a<�b<�#c<c<[b<X.a<��_<i�^<��]<�]<�^<u_<`<�a<X`a<Oa<��_<��]<�u[<*�X<[V<.�S<�IR<F�Q<��Q<&S<UU<�W<�CZ<q�\<�_<H�`<Ka<�:a<�`<�z_<�j^<��]<��]<�^<x._<L�`<��a<C�b<�c<��b<��a< �`<�S_<�6^<
�]<�  �  ��\<�#]<�,^<�R_<1`<�s`<�_<�~^<�W\<��Y<!�V<$T<+�Q<�~P<�P<�P<[XR<b�T<lvW<POZ<s�\<�^<�`<�{`<�`<w_<�]<]<��\<z�\<� ^<�_<�;a<�b<'�c<��c<#0c<��a<�R`<;�^<i`]<9�\<��\< �]<S�^<��_<\x`<�z`<?�_<t�]<%�[<��X<�V<�sS<l|Q<pcP<�UP<NUQ<�9S<��U<I�X<�d[<��]<��_<��`<ʜ`<\�_<��^<6�]<��\<.�\<'k]<#�^<QK`<��a<>c<m�c<6�c<�b<F�a<�_<�P^<k1]<��\<�]<��]<�$_<�$`<\�`<1^`<�=_<3Q]<�Z<��W<,U<��R<*Q<3KP<��P<��Q<�
T<G�V<�Y<�D\<�}^<��_<o�`<dv`<U�_<m�^<�s]<��\<&�\<q�]<H+_<+�`<Rkb<��c<E�c<(�c<��b<a<3X_<��]<��\<��\<�X]<�`^<Ʌ_<Kc`<m�`<P`<��^<x�\<E�Y<�W<bNT<"R<�P<�BP<H�P<��R<��T<��W<CyZ<(]<�_<0E`<*�`<C6`<l@_<�^<g$]<�\<�]<�$^<��_<�_a<�b<W�c<��c<�Sc<�b<�t`<,�^<�]<8�\<
�\<a�]<v�^<��_<�`<�`<ó_<\^<d�[<z�X<�	V<�tS<�zQ<�^P<NNP<KKQ<-S<-�U<%�X<,P[<F�]<{_<�i`<+~`<��_<��^<R�]<�\<�\<A]<Q^<�`<)�a<'c<]�c<)�c<%�b<�fa<��_<�$^<1]<��\<U�\<��]<��^<n�_<�v`<�1`<o_<�"]<ԛZ<a�W<��T<��R<X�P<�P<dP<��Q<v�S<��V<.\Y<\<�H^<��_<�m`<2@`<o_<�L^<o;]<C�\<�\<Q�]<j�^<��`<�.b<�Mc<z�c<�cc<�Ub<*�`<c_<K�]<��\<�  �  )lR<�8S<��T<@W<�WY<��Z<)�Z<�Y<�W<#�T<� Q<(�M<�J<XI<��H<gI<DxK<AsN<��Q<�_U<�LX<FZ<�[<��Z<O�X<��V<�T<��R<�tR<=(S<��T<B�W<ˆZ<<]<�^<�_<��]<��[<��X<�V<��S<�R<��R<u�S<��U<DX<�Z<h
[<��Z<�mY<�V<��S<P<#�L<UJ<c�H<`�H<�!J<��L<-�O<�GS<��V<mEY<�Z<�.[<JZ<�wX<�6V<s'T<z�R<�R<��S<+�U<��X<�[<��]<�$_<��^<}]<�[<�X<"jU<�wS<�R<�S<v�T<��V<5�X<n�Z<�0[<��Z<=�X<;�U<�R<PO<��K<��I<�H<�-I<�J<��M<��P<�sT<�W<��Y<�[<��Z<��Y<�W<tU<�S<+�R<c�R<rT<��V<�Y<�{\<^x^<|>_<�^<Ϳ\<�Z<�(W<=�T<DS<T�R<�nS<4U<lsW<D�Y<a�Z<�$[<�Z< �W<!�T<�QQ<	�M<�K<�JI<P�H<�I<J�K<�N<sR<��U<�uX<smZ<�+[<�Z<Y<9�V<-�T< S<L�R<LS<<"U<�W<�Z<�:]<��^<�+_<=^<�[<�Y<�@V<YT<9�R<��R<��S<m�U<�2X<�Z<�[<`�Z<fzY<�V<ϤS<AP<m�L<aSJ<��H<��H<�J<y�L<�O<�4S<�V<�,Y<��Z<[<�)Z<�TX<V<y T<��R<L�R<խS<��U<��X<t[<ɿ]<��^<��^<�N]<�Z<��W<�=U<LS<�uR<��R<�XT<,�V<_�X<`Z<�[<�iZ<�X<ùU<�NR<��N<�K<��I<ڗH<�H<�J<�_M<u�P<~>T<}eW<c�Y<��Z<��Z<ՈY<qW<�;U<m_S<hrR<t�R<5T<�V<>Y<i<\<�8^<2�^<5`^<Ɂ\<��Y<4�V<qT<��R<�  �  �S<!�S<��U<�W<3�Y<�[<�H[<�8Z<"X<��T<��Q<h>N<��K<A�I<�8I<J<qL<�N<�SR<�U<��X<b�Z<k^[<��Z<PqY<�WW<y3U<^�S<�S<W�S<�jU<;�W<w�Z<K]<��^<��^<W�]<m�[<+!Y<zV<aT<\@S<�KS<NwT<�nV<w�X<4vZ<�i[<|0[<F�Y<�4W<
�S<͍P<dM<��J<f�I<ށI<@�J<�M<�8P<&�S<a�V<%�Y<�,[<p�[<0�Z<m�X<H�V<��T<-�S<ZS<�\T<�_V<e�X<}�[<.�]<B_<B�^<p]<%[<�[X<�U<� T<�>S<��S<�$U<|@W<xcY<�Z<��[<��Z<�Y<�>V<=�R<pO<�L<�eJ<ErI<��I<�tK<~N<-`Q<o�T<��W<�;Z<�n[<4c[<�6Z<�BX<�V<�=T<�OS<8�S<��T<�/W<��Y<J|\<�^^<�_<@�^<��\<�2Z<[xW< U<��S<�DS<�T<�U<\X<�Z<�K[<z[<jZ<65X<�*U<��Q<\oN<��K<��I<�hI<27J<�9L<�O<mR<N�U<��X<ԻZ<��[<�[<��Y<:{W<�VU<��S<k7S<'�S<F�U<	X<��Z<�0]<߻^<�_<�^<��[<nEY<@�V<̂T<l`S<�iS<a�T<��V<ݹX<�Z<|[<@[<	�Y<�>W<T<��P<UeM<+�J<׎I<dzI<ݴJ<�M<~(P<-�S<��V<�yY<|[<�n[<�Z<��X<l�V<��T<S\S<�/S<�0T<s2V<E�X<��[<�]<�^<R�^<�A]<:�Z<[.X<��U<2�S<�S<@�S<h�T<�W<�8Y<��Z<�^[<u�Z<4�X<�V<��R<�MO<-SL<�1J<�=I<؜I<�?K<8�M<�*Q<�T<G�W<SZ<9[<-[<��Y<7X<�U<iT<�S<]NS<��T<��V<�Y<!=\<G^<j�^<�D^<�~\<��Y<�<W<��T<iS<�  �  ��T<0�U<]WW<\ZY<z"[<21\<[3\<�[<�X<��U<B�R<&�O<X-M<��K<�K<L�K<�M<J[P<�}S<��V<�rY<�k[<MQ\<�\<�Z<��X<y�V<�oU<o�T<3U<��V<5�X<]�Z<��\<L/^<jp^<ǔ]<��[<T�Y<UmW<��U<�T<NU<�@V<X<�Z<:�[<=p\<�\<^�Z<KX<HU<M�Q<��N<-�L<ChK<XK<�}L<��N<�Q<��T<��W<�fZ<@
\<��\<��[<�nZ<�uX<-�V<�NU<qU<��U<7_W<��Y<�[<��]<Б^<�p^<�<]<+E[<��X<�V<>wU<��T<�xU<I�V<��X<��Z<� \<��\<�[<:�Y<�.W<	T<�P< "N<�+L<YJK<��K<[&M<�O<ߞR<��U<C�X<F[<�U\<�t\<�[<��Y<��W<
V<�U<�U<H0V<!	X<(GZ<�o\<�^<<�^<�%^<~�\<��Z<�DX<�ZV<0U<�U<��U<��W<��Y<�T[<c\<�d\<?[<=Y<�)V<y�R<Q�O<Y^M<��K<AK<� L<K�M<��P<թS<'�V<��Y<��[<�w\<A5\<��Z<_Y<�W<
�U<��T<�VU<<�V<��X<� [<�]<U^<2�^<J�]<��[<u�Y<V�W<3�U<�U<]1U<�\V<�4X<�2Z<�[<m�\<l \<�Z<4#X<VU<y�Q<��N<��L<�cK<�PK<esL<I�N<�{Q<��T<��W<"NZ<!�[<�o\<]�[<hLZ<�PX<QkV<�%U< �T<��U<!2W<�YY<o�[<�i]<�b^<�A^<M]<S[<��X<��V<}KU<��T<�MU<��V<#�X<��Z<I�[<$V\<��[<��Y<&�V<�S<��P<��M<��K<�K<�mK<�L<�bO<diR<��U<ēX<��Z< \<v>\<`J[<D�Y<��W<��U<\�T<�T<��U<x�W<�Z<�0\<��]<Pg^<_�]<�g\<[JZ<o	X<� V<��T<�  �  ZCW<L<X<�Y<܌[<A�\<�]<^p]<q.\<EZ<KjW<��T<��Q<�O<9=N<��M<�yN<�P<zqR<54U<zX<�Z<�\<R�]<m�]<��\<4[<�uY< X<L4W<F>W<�X<�lY<<[<�u\<.f]<ڕ]<��\<4�[<�%Z<E�X<��W<~(W<��W<�X<2~Z<<1\<�l]</�]<�?]<��[<�\Y<ΚV<��S<6Q<�<O<E#N<WN<�O<��P<�S<WV<n"Y<Q�[<;5]<{�]<�]<�z\<P�Z<�Y<��W<sQW<w�W<��X<$#Z<��[< ]<��]<y�]<`�\<t[[<��Y<PYX<�tW<�RW<EX<�mY<�*[<��\<"�]<s�]<��\<�
[<�X<A�U<0�R<��P<��N<�
N<JXN<��O<J�Q<AuT<�NW<� Z<�0\<��]<o�]<FO]<��[<;6Z<0�X<��W<iOW<��W<�Y<B�Z<u0\<$T]<O�]<�j]<�V\<�Z<�AY<��W<CTW<zW<�qX<>Z<�[<�-]<��]<��]<�_\<�CZ<��W<8�T<fR<E�O<JnN<�N<��N<ZHP<#�R<�`U<c6X<w�Z<�\<	�]<��]<]�\<X[<?�Y<|#X<�WW<bW<,3X<g�Y<X)[<��\<͋]<p�]<0]<��[<sIZ<�X<�W<@HW<��W<��X<ǗZ<pH\<��]<I�]<O]<g�[<bfY<ҡV< �S<V7Q<0;O<�N<�N<GO<J�P<drS<DV<�Y<�p[<,]<��]<�]<X\<��Z<&�X<�W<.'W<�uW<�{X<V�Y<'�[<;�\<"�]<�r]<�\<�-[<��Y<�,X<$IW<|'W<l�W<�BY<��Z<��\<F�]<��]<۶\<��Z<�WX<�U<��R<SP<?�N<�M<�"N< uO<��Q<�?T<W<"�Y< �[<�W]<R�]<�]<G�[<�Y<aX<pSW<W<F�W<Q�X<HjZ<�[<�]<҉]<�,]<�\<ȘZ<�Y<=�W<W<�  �  ��Y<��Z<Sq\<v�]<��^<a#_<��^<�9]<�C[<K�X<��V<�aT<P�R<�jQ<�Q<"�Q<k�R<'�T<W<�Y<^�[<z�]<#�^<�+_<G�^<d�]<�%\<��Z<	�Y<�QY<�xY<�Z<}�Z<9�[<{\<4\<��[<�6[<�iZ<��Y<+[Y<I�Y<�HZ<9�[<j
]<�\^<;&_<�)_<�T^<�\<ͦZ<'MX<��U<N�S<�CR<�\Q<�QQ<6$R<ıS<g�U<�X<NvZ<�\<�F^<�5_<�L_<��^<�T]<��[<��Z<}�Y<"�Y<S�Y<;~Z<L[<1�[<_[\<N\<��[<�[<7LZ<ȭY<�wY<j�Y<��Z<�"\<��]<��^<FR_<D_<��]<�(\<��Y<ȐW<�GU<SS<.�Q<eKQ<ۊQ<7�R<�]T<ΈV<k�X<�9[<�<]<�^<�R_<�!_<%5^<�\<FZ[<?0Z<��Y<&�Y<��Y<��Z<މ[<�$\<�b\<�0\<�[<��Z<kZ<��Y<��Y<?Z<2[<g�\<�^<\_<]U_<T�^<8k]<Cu[<(Y<��V<��T<,�R<7�Q<�CQ<�Q<�S<aU<�IW<-�Y<R�[<��]<E�^<rQ_<>�^<��]<iI\<J�Z<��Y<�uY<�Y<2Z<r�Z<z�[<�?\<hY\< \<3[[<��Z<��Y<P|Y<ͤY<<fZ<ק[<�#]<�s^<�:_<�;_<)d^<��\<��Z<TX<��U<��S<�AR<KXQ<9JQ<�R<��S<S�U<�X<�`Z<��\<�+^<_<�,_<Ww^<F0]<Q�[<dZ<p�Y<�UY<��Y<�PZ<�[<��[<�,\<�\<v�[<]�Z<EZ<x�Y<'LY<+�Y<ܘZ<�[<�p]<�^<&_<-�^<��]<b�[<��Y<�^W<�U< S<h�Q<Q<UQ<7jR<v'T<�RV<��X<+[<]<Hv^<�_<^�^<�]<9�\<~![<t�Y<�UY<OMY<��Y<.�Z<�K[<��[<�$\<,�[<+a[<;�Z<��Y<UVY<'OY<�  �  �\< S]<P�^<��_<�*`<��_<�"_<��]<\<�-Z<eX<��V<t�U<k�T<�mT<��T<��U<w"W<n�X<�Z<�m\<-^<^f_<�`<�#`<�_<_d^<X]<<�[< �Z<fZ<='Z<�Z<o'Z<�3Z<�5Z<q/Z<,#Z<�"Z<mHZ<g�Z<�t[<-�\<��]<^_<Z`<\L`<��_<@�^<ZP]<͉[<K�Y<�W<>yV<�SU<�T<��T<�>U<�ZV<F�W<}�Y<f[<T3]<��^<P�_<Ne`<1`<4__<�'^<��\<߶[<��Z<�yZ<�NZ<MZ<aYZ<�`Z<D_Z<�SZ<�FZ<|MZ<��Z<I[<��[<k]<,h^<ҏ_<�B`<TQ`<!�_<�p^<�\< �Z<h,Y<��W<�V<}U<��T<�T<��U<��V<;jX<!/Z<k\<s�]<�5_<C"`<�c`<��_<K�^<�]<~i\<	c[<ݶZ<'`Z<�FZ<�MZ<�ZZ<o_Z<�[Z<�NZ<�EZ<�YZ<<�Z<J[<�F\<�]<:�^<��_<k]`<�/`<�T_<h�]<6\<`Z<p�X<j�V<�U<��T<\�T<�U<��U<ZQW<��X<,�Z<�\<7B^<��_<D`<RI`<��_<b�^<7]<� \<�[<5�Z<�KZ<�@Z<vLZ<�XZ<�ZZ<-TZ<UGZ<�EZ<�jZ<?�Z<�[<��\<�]<�8_<8`<�``<��_<u�^<�\]<��[<3�Y<-�W<nzV<�QU<m�T<�T</4U<�MV<<�W<�|Y<oP[<]<�^<��_<vE`<�`<�:_<J^<��\<�[<��Z<oMZ<p!Z<:Z<'+Z<�2Z<1Z<�%Z<[Z<� Z<JXZ<��Z<��[<Z�\<=^<�d_</`<�$`<��_<"B^</�\<��Z<�X<MW<��U<%�T<�oT<��T<�cU<�V<�3X<��Y<x�[<��]<��^<J�_<A-`<ھ_<��^<�w]<)0\<�([<�{Z<	$Z<
Z<XZ<jZ<*"Z<�Z<|Z<�
Z<�Z<xoZ<�[<�  �  :p]<��^<}�_<�}`<{y`<��_<��^<�]]<w�[<��Z<@�Y<	�X<�X<̩W<�W<��W<�8X<��X<�Y<>�Z<�K\<ű]<._<`<�`<q`<$�_<�^<�,]<�[<�Z<�Y<�X<X<�W<�W<N�W<�cX<w%Y<�Z<�D[<W�\<��]<�L_<LA`<��`<Hp`<O�_<�h^<B]<��[<�xZ<�vY<��X<:X<˽W<��W<�	X<3�X<�gY<�fZ<p�[<��\<�X^<��_<�{`<��`<�t`<.�_<�K^<h�\<��[<AcZ<\hY<�X<X<�W<q�W<W*X<D�X<̕Y<��Z<I�[<�,]<&�^<��_<w�`<\�`<rN`<7U_<�^<c�\<tQ[<(-Z<�;Y<�~X<#�W<N�W<�W<�=X<p�X<��Y<��Z<�
\<�j]<g�^<i�_<d�`<R�`<1`<�%_< �]<�j\<![<�Z<�Y<�gX<��W<��W<�W<�VX<jY<��Y<�Z<|C\<�]<b _<7`<ʰ`<�`<�	`<��^<�]<�-\<�Z<�Y<�X<�IX<��W<v�W<]�W<�iX<� Y<WZ<�*[<�v\<e�]<W/_<�4`<ѵ`<�`<h�_<Ѱ^<ZP]<��[<�Z<H�Y<��X<�2X<��W<��W<� X<��X<rHY<r=Z<e[<G�\<�^<h_<GZ`<��`<��`<�_<�w^<�]<:�[<�Z<�zY<��X<�X<2�W<4�W<g�W<�X<�WY<TZ<�[<��\<�=^<]~_<�[`<��`<�P`<j_<�#^<�\<�e[<47Z<l;Y<�sX<+�W<�W<��W<��W<�X<!iY<�nZ<��[<t]<�c^<��_<�``<6�`<|!`<<'_<��]<�p\<�[<$�Y<Y<gIX<.�W<ʉW<3�W<�X<��X<��Y<��Z<��[<�4]<��^<��_<@m`<��`<��_<��^<H�]<71\<^�Z<y�Y<��X< +X<ӲW<+�W<�W<!X<��X<P�Y<��Z<w\<�  �  b�]<�1_<V`<�'`<#�_<��^<^A]<�\<I	[<�kZ<~ Z<Z<�Z<p#Z<�&Z<�!Z<�Z<Z<&-Z<k�Z<<[<�H\<��]<3�^<k�_<28`<��_<M�^<��]<��[<��Y<h)X<�V<�cU<U�T<��T<��T<�V<9uW<�%Y<V�Z<��\<}k^<�_<R>`<�'`<fm_<3B^<'�\<��[<U�Z<�mZ<:Z<V5Z<�BZ<NNZ<$PZ<�HZ<�=Z<BZ<�qZ<�Z<(�[<��\<�5^<�k_<&8`<�d`<;�_< �^<�"]<�U[<i�Y<I�W<]VV<�AU<��T<��T<rU<�V<D#X<��Y<$�[<�z]<I�^<5`<�a`<�`<!'_<'�]<��\<߄[<��Z< fZ<�DZ<`HZ<VZ<�\Z<[Z<POZ<�DZ<�RZ<�Z<�([<\<�P]<��^<�_<aU`<6F`<چ_<4^<?�\<T�Z<B�X<�BW<��U<��T<4�T<��T<&�U<W<u�X<J}Z<CR\<�^<bf_<�7`<�Z`<��_<��^<�s]<G4\<�;[<��Z<�SZ<�AZ<�JZ<�VZ<�YZ<TZ<jFZ<m@Z<\Z<ҶZ<�g[<�r\<b�]<�_<��_<g]`<c`<d_<�]<��[<�Z<�MX<]�V<L�U<��T<g�T<�#U<E+V<ݗW<9GY<�[<��\<Z�^<��_<W`<>`<{�_<�S^<  ]<��[<��Z<TtZ<>Z<u6Z<#AZ<�IZ<�HZ<{>Z<�0Z<2Z<_Z<��Z<�[<B�\<�^<7L_<U`<�@`<U�_<Q�^<��\<�*[<�UY<��W<!)V<�U<�T<B�T<�DU<qV<��W<�Y<x�[<�O]<��^<��_<6`<?�_<��^<��]<Mi\<�S[<<�Z<^2Z<�Z<�Z<�Z<�%Z<�#Z<�Z<�Z<�Z<�^Z<e�Z<�[<�]<�k^<�_<`<Z`<LO_<��]<M\<ExZ<q�X<W<�U<��T<ShT<g�T<P�U<��V<�zX<�EZ<�\<�  �  �O]<��^<#$_<��^<��]<�\\<F�Z<c�Y<�MY<4]Y<n�Y<�Z<�n[<��[<�(\<1�[<�F[<Z{Z<&�Y<�PY<�aY<[Z<=[<�\<_^<T�^<�#_<�q^<W�\<��Z<]�X<v?V<VT<dR<�ZQ<)Q<�Q<�HS<VEU<=�W<Y�Y<*\<��]<��^<J9_<B�^<�s]<a�[<'�Z<�Y<eY<)�Y<�DZ<l[<��[<@@\<�G\<��[<�1[<(eZ<i�Y<�uY<-�Y<D�Z<��[<of]<y�^<�R_<�1_<[9^<�\<�^Z<��W<_�U<��S<�!R<\Q<�tQ<TgR<�T<�'V<�X<U�Z<��\<�y^<�C_<E5_<�c^<�]<��[<�UZ<��Y<�|Y<��Y<ŘZ<�f[<�\<S]\<U>\<͹[<p�Z<-Z<Q�Y<!~Y<�Y<Z�Z<?f\<q�]<��^<�Y_<��^<P�]<�[<��Y<�/W<0�T< S<N�Q<cHQ<��Q<��R<��T<W�V<�LY<~�[<�]<'�^<�W_<�_<��]<�\<�[<Z<̀Y<��Y<=Z<6�Z<�[<�0\<E\\<H\<�x[<U�Z<��Y<�~Y<�Y<6Z<Nf[<��\<�>^<�"_<�H_<�^<Q]<�[<Q�X<�cV<�=T<ֈR<QQ<=MQ<��Q<lS<�gU<z�W<BZ<mH\<�	^<�_<�Q_<��^<��]<�\<�Z<�Y<�nY<�Y<�HZ<�[<��[<�;\<\@\<��[<q$[<:UZ<��Y<$`Y<(�Y<�zZ<��[<G]<υ^<�._<�_<�^<�_\<�4Z<O�W<�U<�xS<��Q<�.Q<7GQ<-:R<��S<*�U<UX<��Z<�\<N^<�_<+	_<�6^<��\<�b[<�%Z<;kY<
JY<��Y<`cZ<_0[<��[<�%\<k\<߁[<��Z<��Y<VfY<�GY<�Y<}�Z<�0\<��]<��^<K#_<X�^<g|]<P�[<yWY<U�V<d�T<��R<��Q<(Q<�qQ<d�R<M{T<�V<�Y<I`[<�  �  �D\<�y]<9�]<��\<u[<�Y<�*X<=W<J"W<;�W<�Y<ɲZ<N0\<D;]<N�]<K]<M�[<!YZ<�X<ҟW<�W<�dW<
}X<�Z<��[<1]<e�]<�U]<r�[<��Y<z�V<%T<��Q<�jO<�&N<��M<8�N<n�P<U�R<�U<ϑX<W[<6�\<r�]<��]<��\<��Z<%CY<B�W<�<W<�jW<oXX<��Y<y_[<�\<��]<�]<[�\<��[<7�Y<o�X<��W<�IW<��W<�-Y<�Z<>�\<��]<��]<�(]<�r[<�Y<9V<hS<Q�P<�O<]N<i<N<�dO<|hQ<��S<>�V<��Y<��[<ib]<`�]<�u]<:2\<�}Z<G�X<4�W<�FW<Y�W<��X<T`Z<��[<~+]<��]<P�]<�\<�[<�Y<9)X<�bW<�dW<�;X< �Y<�x[<P�\<G�]<��]<ר\<�Z<xX<1?U<'�R<D2P<d�N<�N<=�N<��O<98R<��T<��W<�hZ<�y\<��]<w�]<L]<�[<H�Y<`]X<�oW<�UW<�X<5SY<U�Z<e\<�o]<��]<�A]<\<��Z<D�X<f�W<�EW<�W<��X<�GZ<c\<�V]<\�]<Mz]<�\<��Y<c!W<IT<�Q<�O<�JN<�N<��N<T�P<bS<�U<x�X<y-[<��\<��]<��]<ˮ\<�[<zTY<�W<�HW<tW<_X<��Y<�`[<G�\<�]<i�]<�\<t�[<Q�Y<�vX<;wW<�1W<m�W<�Y<��Z<�l\<�]<	�]<�]<�I[<��X<�V<	<S<��P<��N<%�M<=N<�7O<�;Q<��S<Q�V<�gY<"�[<�6]<��]<�I]<%\<�OZ<�X<�xW<�W<��W<*�X<l*Z<��[<��\<��]<�M]<�T\<x�Z<MIY<�W<�+W<f.W<X<q�Y<�B[<o�\< �]<$�]<Rq\<�tZ<s�W<}U<�FR<��O<�dN<(�M<�FN<��O<N�Q<�T<��W<�2Z<�  �  �#[<�9\<�'\<�[<�=Y<d<W<��U<��T<�U<_:V<(+X<�mZ<�\<��]<cj^<��]<6\<��Y<��W<�U<F�T</�T<D�U<c�W<Q�Y<�g[<�N\<� \<�Z<~yX<N~U<yIR<
IO<�L<
pK<*K<�L<�"N<��P<hT<�<W<d�Y<��[<nm\<��[<�Z<e�X<`�V<�WU<��T<tU<>�V<�Y<"R[<�A]<h^<�y^<�r]<�[<�XY<6W<2�U<
�T<SU<8�V<��X<q�Z<\<,�\<o�[<�NZ<�W<`�T<lQ<o�N<ttL<�_K<��K<��L<�$O<nR<�LU<�SX<ȽZ<�1\<w�\<N�[<�Z<XX<nEV<@&U<�U<I�U<��W<<�Y<�\<�]<ќ^<tL^<��\<��Z<�X<��V<�PU<$�T<�U<E:W<58Y<�[<RH\<�z\<9�[<��Y<@�V<D�S<ZeP<�M<&�K<EK<��K<��M<3P<�'S<YV<I8Y<�X[<�m\<�Z\<3?[<TpY<�nW<G�U<��T<o7U<gnV<�_X<��Z<��\<�.^<�^<��]<fM\<�Z<8�W<V<�U<�U<9V<��W<j�Y<�[< t\<+E\<-�Z<k�X<0�U<emR<mO<M<��K<�MK<�@L<cEN<�Q<.9T<Y\W<XZ<��[<Ç\<\<��Z<�X<��V<ofU<��T<l}U<��V<�Y<,S[<@]<zc^<@r^<�h]<��[<�HY<�#W<�U<"�T<�8U<U�V<�oX<fZ<��[<�k\<R�[<A&Z<�W<WqT<8@Q<�fN<�GL<�2K<�UK<�L<"�N<<�Q<� U<�'X<=�Z<!\<�U\<Њ[<��Y<�W<�V<Y�T<��T<��U<�wW<�Y<X�[<�]<Qd^<�^<�\<>�Z<�hX<IiV<U<��T</uU<�W<�Y<��Z<@\<BD\< O[<�HY<�xV<�IS<�+P<�M<ιK<�
K<��K<BHM<��O<��R<w"V<�Y<�  �  eNZ<M[<�[<շY<{�W<��U<[�S<US<1yS<�U<eW<�Z<�\<�Y^<7�^<7^<� \<��Y<�V<��T<-JS<\"S<�!T<�U<s3X<� Z<B@[<h;[<��Y<��W<�vT<rQ<A�M<;/K<۝I<�RI<BYJ<ۉL<��O<;�R<�NV<�Y<��Z<�s[<�Z<D3Y<�W<��T<ӋS<Z/S<*T<-�U<8pX<L*[<Zy]<a�^<��^<Y�]<l{[<��X<�0V<c;T<�JS<��S<��T<��V<Y<��Z<|�[<�"[<�yY<��V<��S<
P<u M<ʳJ<�I<b�I<�K<F�M<b�P<M?T<�pW<��Y<�O[<}x[<wZ<��X<�hV<6{T<	`S<�gS<�T<�V<�lY<m\<J^<�_<#�^<w]<w�Z<L�W<�vU< �S<�>S<��S<�zU<�W<�Y<�'[<�[<P�Z<��X<��U<�UR<o�N<�L<0)J<�lI<�J<��K<��N<�Q<�\U<T]X<�Z<Ȁ[<�@[<w�Y<��W<�U<�S<s?S<լS<09U<ÙW<�TZ<A�\<�^<4_<�D^<vT\<��Y<\W<�T<�wS<2NS<�KT<�'V<�ZX<�FZ<{e[<�_[<Z<�W<ԚT<R+Q<+�M<&SK<��I<vI<r|J<k�L<��O<�S<,nV<k1Y<��Z<�[<4�Z<>IY<:!W<	U<z�S<b;S<�T<��U<tX<R+[<�w]<��^<c�^<�]<Un[<ɸX<
V<&T<�2S<$nS<��T<��V<��X<Y�Z<,m[<��Z<hQY<�V<�WS<G�O<�L<�J<,\I<{�I<��J<�qM<>�P<sT<�DW<5�Y<)$[<yL[<vJZ<BnX<D:V<}KT<�.S<5S<�eT<��V<k6Y<��[<�]<,�^<9x^<��\<�kZ<7�W<j?U<6�S<KS<��S<=EU<]mW<x�Y<��Z<�S[<FxZ<�oX<��U<{R<ڿN<��K<�I<�2I<D�I<��K<BgN<��Q<F&U<�'X<�  �  � Z<��Z<�Z<?=Y<tW<��T<�&S<WkR<��R<�T<�W<��Y<Ҧ\<4v^<�_<�(^<M\<d[Y<y}V<iT<�R<WR<�|S<jcU<ǨW<�Y<��Z<��Z<�Y<\IW<zT<��P<�AM<ڕJ<��H<��H<�I<��K<UO<��R<E�U<��X<Q�Z<�[<RdZ<�X<�xV<�UT<�R<�R<�zS<WzU<2X<K[<Շ]<b�^<�
_<��]<�l[<��X<��U<�S<��R<��R<�:T<{SV<f�X<�^Z<�5[<��Z<-Y<�zV<2 S<%�O<ZrL<�J<a�H<�	I<��J<lM<�[P<��S<yW<�Y<��Z< [<~Z<\X<��U<�S<[�R<r�R<8T<�eV<�=Y<�\<�3^<k3_<��^<�]<��Z<��W<�U<�@S<ߞR<8S<��T<�W<-;Y<D�Z<2[<4aZ<iYX<�bU<\�Q<qxN<S�K<��I<F�H<VaI<AK<ZN<z�Q<�U<�X<R5Z<y*[<#�Z<�oY<�QW<fU<�YS<~�R<�S<4�T<sLW<(4Z<;�\<��^<7_<E]^<�Q\<ōY<n�V<�NT<��R<B�R<��S<�U<�W<�Y<:[<�[<;�Y<LmW<U>T<��P<�eM<��J<�I<�H<)�I<=L<4O<Q�R<�V<Q�X<j�Z<�2[<z|Z<��X<��V<)gT<"�R<��R<�S<�U<�5X<P[<�]<��^<s_<g�]<�_[<�X<d�U<��S<��R<$�R<�T<U4V<sX<e;Z<s[<ϫZ<�Y<�PV<R�R<mpO<FL<�I<~�H<��H<�UJ<��L<�/P<�S<��V<�qY<��Z<�Z<��Y<��W<N�U<S�S</�R<ѝR<%�S<}0V<>Y<F�[<e�]<��^<��^<��\<�OZ<�gW<N�T<�	S<�hR< S<5�T<T�V<�Y<_�Z<��Z<;*Z<�!X<:*U<c�Q<�>N<|NK<�MI<d�H<�'I<�K<�M<!PQ<]�T<-�W<�  �  eNZ<M[<�[<շY<{�W<��U<[�S<US<1yS<�U<eW<�Z<�\<�Y^<7�^<7^<� \<��Y<�V<��T<-JS<\"S<�!T<�U<s3X<� Z<B@[<h;[<��Y<��W<�vT<rQ<A�M<;/K<۝I<�RI<BYJ<ۉL<��O<;�R<�NV<�Y<��Z<�s[<�Z<D3Y<�W<��T<ӋS<Z/S<*T<-�U<8pX<L*[<Zy]<a�^<��^<Y�]<l{[<��X<�0V<c;T<�JS<��S<��T<��V<Y<��Z<|�[<�"[<�yY<��V<��S<
P<u M<ʳJ<�I<b�I<�K<F�M<b�P<M?T<�pW<��Y<�O[<}x[<wZ<��X<�hV<6{T<	`S<�gS<�T<�V<�lY<m\<J^<�_<#�^<w]<w�Z<L�W<�vU< �S<�>S<��S<�zU<�W<�Y<�'[<�[<P�Z<��X<��U<�UR<o�N<�L<0)J<�lI<�J<��K<��N<�Q<�\U<T]X<�Z<Ȁ[<�@[<w�Y<��W<�U<�S<s?S<լS<09U<ÙW<�TZ<A�\<�^<4_<�D^<vT\<��Y<\W<�T<�wS<2NS<�KT<�'V<�ZX<�FZ<{e[<�_[<Z<�W<ԚT<R+Q<+�M<&SK<��I<vI<r|J<k�L<��O<�S<,nV<k1Y<��Z<�[<4�Z<>IY<:!W<	U<z�S<b;S<�T<��U<tX<R+[<�w]<��^<c�^<�]<Un[<ɸX<
V<&T<�2S<$nS<��T<��V<��X<Y�Z<,m[<��Z<hQY<�V<�WS<G�O<�L<�J<,\I<{�I<��J<�qM<>�P<sT<�DW<5�Y<)$[<yL[<vJZ<BnX<D:V<}KT<�.S<5S<�eT<��V<k6Y<��[<�]<,�^<9x^<��\<�kZ<7�W<j?U<6�S<KS<��S<=EU<]mW<x�Y<��Z<�S[<FxZ<�oX<��U<{R<ڿN<��K<�I<�2I<D�I<��K<BgN<��Q<F&U<�'X<�  �  �#[<�9\<�'\<�[<�=Y<d<W<��U<��T<�U<_:V<(+X<�mZ<�\<��]<cj^<��]<6\<��Y<��W<�U<F�T</�T<D�U<c�W<Q�Y<�g[<�N\<� \<�Z<~yX<N~U<yIR<
IO<�L<
pK<*K<�L<�"N<��P<hT<�<W<d�Y<��[<nm\<��[<�Z<e�X<`�V<�WU<��T<tU<>�V<�Y<"R[<�A]<h^<�y^<�r]<�[<�XY<6W<2�U<
�T<SU<8�V<��X<q�Z<\<,�\<o�[<�NZ<�W<`�T<lQ<o�N<ttL<�_K<��K<��L<�$O<nR<�LU<�SX<ȽZ<�1\<w�\<N�[<�Z<XX<nEV<@&U<�U<I�U<��W<<�Y<�\<�]<ќ^<tL^<��\<��Z<�X<��V<�PU<$�T<�U<E:W<58Y<�[<RH\<�z\<9�[<��Y<@�V<D�S<ZeP<�M<&�K<EK<��K<��M<3P<�'S<YV<I8Y<�X[<�m\<�Z\<3?[<TpY<�nW<G�U<��T<o7U<gnV<�_X<��Z<��\<�.^<�^<��]<fM\<�Z<8�W<V<�U<�U<9V<��W<j�Y<�[< t\<+E\<-�Z<k�X<0�U<emR<mO<M<��K<�MK<�@L<cEN<�Q<.9T<Y\W<XZ<��[<Ç\<\<��Z<�X<��V<ofU<��T<l}U<��V<�Y<,S[<@]<zc^<@r^<�h]<��[<�HY<�#W<�U<"�T<�8U<U�V<�oX<fZ<��[<�k\<R�[<A&Z<�W<WqT<8@Q<�fN<�GL<�2K<�UK<�L<"�N<<�Q<� U<�'X<=�Z<!\<�U\<Њ[<��Y<�W<�V<Y�T<��T<��U<�wW<�Y<X�[<�]<Qd^<�^<�\<>�Z<�hX<IiV<U<��T</uU<�W<�Y<��Z<@\<BD\< O[<�HY<�xV<�IS<�+P<�M<ιK<�
K<��K<BHM<��O<��R<w"V<�Y<�  �  �D\<�y]<9�]<��\<u[<�Y<�*X<=W<J"W<;�W<�Y<ɲZ<N0\<D;]<N�]<K]<M�[<!YZ<�X<ҟW<�W<�dW<
}X<�Z<��[<1]<e�]<�U]<r�[<��Y<z�V<%T<��Q<�jO<�&N<��M<8�N<n�P<U�R<�U<ϑX<W[<6�\<r�]<��]<��\<��Z<%CY<B�W<�<W<�jW<oXX<��Y<y_[<�\<��]<�]<[�\<��[<7�Y<o�X<��W<�IW<��W<�-Y<�Z<>�\<��]<��]<�(]<�r[<�Y<9V<hS<Q�P<�O<]N<i<N<�dO<|hQ<��S<>�V<��Y<��[<ib]<`�]<�u]<:2\<�}Z<G�X<4�W<�FW<Y�W<��X<T`Z<��[<~+]<��]<P�]<�\<�[<�Y<9)X<�bW<�dW<�;X< �Y<�x[<P�\<G�]<��]<ר\<�Z<xX<1?U<'�R<D2P<d�N<�N<=�N<��O<98R<��T<��W<�hZ<�y\<��]<w�]<L]<�[<H�Y<`]X<�oW<�UW<�X<5SY<U�Z<e\<�o]<��]<�A]<\<��Z<D�X<f�W<�EW<�W<��X<�GZ<c\<�V]<\�]<Mz]<�\<��Y<c!W<IT<�Q<�O<�JN<�N<��N<T�P<bS<�U<x�X<y-[<��\<��]<��]<ˮ\<�[<zTY<�W<�HW<tW<_X<��Y<�`[<G�\<�]<i�]<�\<t�[<Q�Y<�vX<;wW<�1W<m�W<�Y<��Z<�l\<�]<	�]<�]<�I[<��X<�V<	<S<��P<��N<%�M<=N<�7O<�;Q<��S<Q�V<�gY<"�[<�6]<��]<�I]<%\<�OZ<�X<�xW<�W<��W<*�X<l*Z<��[<��\<��]<�M]<�T\<x�Z<MIY<�W<�+W<f.W<X<q�Y<�B[<o�\< �]<$�]<Rq\<�tZ<s�W<}U<�FR<��O<�dN<(�M<�FN<��O<N�Q<�T<��W<�2Z<�  �  �O]<��^<#$_<��^<��]<�\\<F�Z<c�Y<�MY<4]Y<n�Y<�Z<�n[<��[<�(\<1�[<�F[<Z{Z<&�Y<�PY<�aY<[Z<=[<�\<_^<T�^<�#_<�q^<W�\<��Z<]�X<v?V<VT<dR<�ZQ<)Q<�Q<�HS<VEU<=�W<Y�Y<*\<��]<��^<J9_<B�^<�s]<a�[<'�Z<�Y<eY<)�Y<�DZ<l[<��[<@@\<�G\<��[<�1[<(eZ<i�Y<�uY<-�Y<D�Z<��[<of]<y�^<�R_<�1_<[9^<�\<�^Z<��W<_�U<��S<�!R<\Q<�tQ<TgR<�T<�'V<�X<U�Z<��\<�y^<�C_<E5_<�c^<�]<��[<�UZ<��Y<�|Y<��Y<ŘZ<�f[<�\<S]\<U>\<͹[<p�Z<-Z<Q�Y<!~Y<�Y<Z�Z<?f\<q�]<��^<�Y_<��^<P�]<�[<��Y<�/W<0�T< S<N�Q<cHQ<��Q<��R<��T<W�V<�LY<~�[<�]<'�^<�W_<�_<��]<�\<�[<Z<̀Y<��Y<=Z<6�Z<�[<�0\<E\\<H\<�x[<U�Z<��Y<�~Y<�Y<6Z<Nf[<��\<�>^<�"_<�H_<�^<Q]<�[<Q�X<�cV<�=T<ֈR<QQ<=MQ<��Q<lS<�gU<z�W<BZ<mH\<�	^<�_<�Q_<��^<��]<�\<�Z<�Y<�nY<�Y<�HZ<�[<��[<�;\<\@\<��[<q$[<:UZ<��Y<$`Y<(�Y<�zZ<��[<G]<υ^<�._<�_<�^<�_\<�4Z<O�W<�U<�xS<��Q<�.Q<7GQ<-:R<��S<*�U<UX<��Z<�\<N^<�_<+	_<�6^<��\<�b[<�%Z<;kY<
JY<��Y<`cZ<_0[<��[<�%\<k\<߁[<��Z<��Y<VfY<�GY<�Y<}�Z<�0\<��]<��^<K#_<X�^<g|]<P�[<yWY<U�V<d�T<��R<��Q<(Q<�qQ<d�R<M{T<�V<�Y<I`[<�  �  b�]<�1_<V`<�'`<#�_<��^<^A]<�\<I	[<�kZ<~ Z<Z<�Z<p#Z<�&Z<�!Z<�Z<Z<&-Z<k�Z<<[<�H\<��]<3�^<k�_<28`<��_<M�^<��]<��[<��Y<h)X<�V<�cU<U�T<��T<��T<�V<9uW<�%Y<V�Z<��\<}k^<�_<R>`<�'`<fm_<3B^<'�\<��[<U�Z<�mZ<:Z<V5Z<�BZ<NNZ<$PZ<�HZ<�=Z<BZ<�qZ<�Z<(�[<��\<�5^<�k_<&8`<�d`<;�_< �^<�"]<�U[<i�Y<I�W<]VV<�AU<��T<��T<rU<�V<D#X<��Y<$�[<�z]<I�^<5`<�a`<�`<!'_<'�]<��\<߄[<��Z< fZ<�DZ<`HZ<VZ<�\Z<[Z<POZ<�DZ<�RZ<�Z<�([<\<�P]<��^<�_<aU`<6F`<چ_<4^<?�\<T�Z<B�X<�BW<��U<��T<4�T<��T<&�U<W<u�X<J}Z<CR\<�^<bf_<�7`<�Z`<��_<��^<�s]<G4\<�;[<��Z<�SZ<�AZ<�JZ<�VZ<�YZ<TZ<jFZ<m@Z<\Z<ҶZ<�g[<�r\<b�]<�_<��_<g]`<c`<d_<�]<��[<�Z<�MX<]�V<L�U<��T<g�T<�#U<E+V<ݗW<9GY<�[<��\<Z�^<��_<W`<>`<{�_<�S^<  ]<��[<��Z<TtZ<>Z<u6Z<#AZ<�IZ<�HZ<{>Z<�0Z<2Z<_Z<��Z<�[<B�\<�^<7L_<U`<�@`<U�_<Q�^<��\<�*[<�UY<��W<!)V<�U<�T<B�T<�DU<qV<��W<�Y<x�[<�O]<��^<��_<6`<?�_<��^<��]<Mi\<�S[<<�Z<^2Z<�Z<�Z<�Z<�%Z<�#Z<�Z<�Z<�Z<�^Z<e�Z<�[<�]<�k^<�_<`<Z`<LO_<��]<M\<ExZ<q�X<W<�U<��T<ShT<g�T<P�U<��V<�zX<�EZ<�\<�  �  :p]<��^<}�_<�}`<{y`<��_<��^<�]]<w�[<��Z<@�Y<	�X<�X<̩W<�W<��W<�8X<��X<�Y<>�Z<�K\<ű]<._<`<�`<q`<$�_<�^<�,]<�[<�Z<�Y<�X<X<�W<�W<N�W<�cX<w%Y<�Z<�D[<W�\<��]<�L_<LA`<��`<Hp`<O�_<�h^<B]<��[<�xZ<�vY<��X<:X<˽W<��W<�	X<3�X<�gY<�fZ<p�[<��\<�X^<��_<�{`<��`<�t`<.�_<�K^<h�\<��[<AcZ<\hY<�X<X<�W<q�W<W*X<D�X<̕Y<��Z<I�[<�,]<&�^<��_<w�`<\�`<rN`<7U_<�^<c�\<tQ[<(-Z<�;Y<�~X<#�W<N�W<�W<�=X<p�X<��Y<��Z<�
\<�j]<g�^<i�_<d�`<R�`<1`<�%_< �]<�j\<![<�Z<�Y<�gX<��W<��W<�W<�VX<jY<��Y<�Z<|C\<�]<b _<7`<ʰ`<�`<�	`<��^<�]<�-\<�Z<�Y<�X<�IX<��W<v�W<]�W<�iX<� Y<WZ<�*[<�v\<e�]<W/_<�4`<ѵ`<�`<h�_<Ѱ^<ZP]<��[<�Z<H�Y<��X<�2X<��W<��W<� X<��X<rHY<r=Z<e[<G�\<�^<h_<GZ`<��`<��`<�_<�w^<�]<:�[<�Z<�zY<��X<�X<2�W<4�W<g�W<�X<�WY<TZ<�[<��\<�=^<]~_<�[`<��`<�P`<j_<�#^<�\<�e[<47Z<l;Y<�sX<+�W<�W<��W<��W<�X<!iY<�nZ<��[<t]<�c^<��_<�``<6�`<|!`<<'_<��]<�p\<�[<$�Y<Y<gIX<.�W<ʉW<3�W<�X<��X<��Y<��Z<��[<�4]<��^<��_<@m`<��`<��_<��^<H�]<71\<^�Z<y�Y<��X< +X<ӲW<+�W<�W<!X<��X<P�Y<��Z<w\<�  �  �\< S]<P�^<��_<�*`<��_<�"_<��]<\<�-Z<eX<��V<t�U<k�T<�mT<��T<��U<w"W<n�X<�Z<�m\<-^<^f_<�`<�#`<�_<_d^<X]<<�[< �Z<fZ<='Z<�Z<o'Z<�3Z<�5Z<q/Z<,#Z<�"Z<mHZ<g�Z<�t[<-�\<��]<^_<Z`<\L`<��_<@�^<ZP]<͉[<K�Y<�W<>yV<�SU<�T<��T<�>U<�ZV<F�W<}�Y<f[<T3]<��^<P�_<Ne`<1`<4__<�'^<��\<߶[<��Z<�yZ<�NZ<MZ<aYZ<�`Z<D_Z<�SZ<�FZ<|MZ<��Z<I[<��[<k]<,h^<ҏ_<�B`<TQ`<!�_<�p^<�\< �Z<h,Y<��W<�V<}U<��T<�T<��U<��V<;jX<!/Z<k\<s�]<�5_<C"`<�c`<��_<K�^<�]<~i\<	c[<ݶZ<'`Z<�FZ<�MZ<�ZZ<o_Z<�[Z<�NZ<�EZ<�YZ<<�Z<J[<�F\<�]<:�^<��_<k]`<�/`<�T_<h�]<6\<`Z<p�X<j�V<�U<��T<\�T<�U<��U<ZQW<��X<,�Z<�\<7B^<��_<D`<RI`<��_<b�^<7]<� \<�[<5�Z<�KZ<�@Z<vLZ<�XZ<�ZZ<-TZ<UGZ<�EZ<�jZ<?�Z<�[<��\<�]<�8_<8`<�``<��_<u�^<�\]<��[<3�Y<-�W<nzV<�QU<m�T<�T</4U<�MV<<�W<�|Y<oP[<]<�^<��_<vE`<�`<�:_<J^<��\<�[<��Z<oMZ<p!Z<:Z<'+Z<�2Z<1Z<�%Z<[Z<� Z<JXZ<��Z<��[<Z�\<=^<�d_</`<�$`<��_<"B^</�\<��Z<�X<MW<��U<%�T<�oT<��T<�cU<�V<�3X<��Y<x�[<��]<��^<J�_<A-`<ھ_<��^<�w]<)0\<�([<�{Z<	$Z<
Z<XZ<jZ<*"Z<�Z<|Z<�
Z<�Z<xoZ<�[<�  �  ��Y<��Z<Sq\<v�]<��^<a#_<��^<�9]<�C[<K�X<��V<�aT<P�R<�jQ<�Q<"�Q<k�R<'�T<W<�Y<^�[<z�]<#�^<�+_<G�^<d�]<�%\<��Z<	�Y<�QY<�xY<�Z<}�Z<9�[<{\<4\<��[<�6[<�iZ<��Y<+[Y<I�Y<�HZ<9�[<j
]<�\^<;&_<�)_<�T^<�\<ͦZ<'MX<��U<N�S<�CR<�\Q<�QQ<6$R<ıS<g�U<�X<NvZ<�\<�F^<�5_<�L_<��^<�T]<��[<��Z<}�Y<"�Y<S�Y<;~Z<L[<1�[<_[\<N\<��[<�[<7LZ<ȭY<�wY<j�Y<��Z<�"\<��]<��^<FR_<D_<��]<�(\<��Y<ȐW<�GU<SS<.�Q<eKQ<ۊQ<7�R<�]T<ΈV<k�X<�9[<�<]<�^<�R_<�!_<%5^<�\<FZ[<?0Z<��Y<&�Y<��Y<��Z<މ[<�$\<�b\<�0\<�[<��Z<kZ<��Y<��Y<?Z<2[<g�\<�^<\_<]U_<T�^<8k]<Cu[<(Y<��V<��T<,�R<7�Q<�CQ<�Q<�S<aU<�IW<-�Y<R�[<��]<E�^<rQ_<>�^<��]<iI\<J�Z<��Y<�uY<�Y<2Z<r�Z<z�[<�?\<hY\< \<3[[<��Z<��Y<P|Y<ͤY<<fZ<ק[<�#]<�s^<�:_<�;_<)d^<��\<��Z<TX<��U<��S<�AR<KXQ<9JQ<�R<��S<S�U<�X<�`Z<��\<�+^<_<�,_<Ww^<F0]<Q�[<dZ<p�Y<�UY<��Y<�PZ<�[<��[<�,\<�\<v�[<]�Z<EZ<x�Y<'LY<+�Y<ܘZ<�[<�p]<�^<&_<-�^<��]<b�[<��Y<�^W<�U< S<h�Q<Q<UQ<7jR<v'T<�RV<��X<+[<]<Hv^<�_<^�^<�]<9�\<~![<t�Y<�UY<OMY<��Y<.�Z<�K[<��[<�$\<,�[<+a[<;�Z<��Y<UVY<'OY<�  �  ZCW<L<X<�Y<܌[<A�\<�]<^p]<q.\<EZ<KjW<��T<��Q<�O<9=N<��M<�yN<�P<zqR<54U<zX<�Z<�\<R�]<m�]<��\<4[<�uY< X<L4W<F>W<�X<�lY<<[<�u\<.f]<ڕ]<��\<4�[<�%Z<E�X<��W<~(W<��W<�X<2~Z<<1\<�l]</�]<�?]<��[<�\Y<ΚV<��S<6Q<�<O<E#N<WN<�O<��P<�S<WV<n"Y<Q�[<;5]<{�]<�]<�z\<P�Z<�Y<��W<sQW<w�W<��X<$#Z<��[< ]<��]<y�]<`�\<t[[<��Y<PYX<�tW<�RW<EX<�mY<�*[<��\<"�]<s�]<��\<�
[<�X<A�U<0�R<��P<��N<�
N<JXN<��O<J�Q<AuT<�NW<� Z<�0\<��]<o�]<FO]<��[<;6Z<0�X<��W<iOW<��W<�Y<B�Z<u0\<$T]<O�]<�j]<�V\<�Z<�AY<��W<CTW<zW<�qX<>Z<�[<�-]<��]<��]<�_\<�CZ<��W<8�T<fR<E�O<JnN<�N<��N<ZHP<#�R<�`U<c6X<w�Z<�\<	�]<��]<]�\<X[<?�Y<|#X<�WW<bW<,3X<g�Y<X)[<��\<͋]<p�]<0]<��[<sIZ<�X<�W<@HW<��W<��X<ǗZ<pH\<��]<I�]<O]<g�[<bfY<ҡV< �S<V7Q<0;O<�N<�N<GO<J�P<drS<DV<�Y<�p[<,]<��]<�]<X\<��Z<&�X<�W<.'W<�uW<�{X<V�Y<'�[<;�\<"�]<�r]<�\<�-[<��Y<�,X<$IW<|'W<l�W<�BY<��Z<��\<F�]<��]<۶\<��Z<�WX<�U<��R<SP<?�N<�M<�"N< uO<��Q<�?T<W<"�Y< �[<�W]<R�]<�]<G�[<�Y<aX<pSW<W<F�W<Q�X<HjZ<�[<�]<҉]<�,]<�\<ȘZ<�Y<=�W<W<�  �  ��T<0�U<]WW<\ZY<z"[<21\<[3\<�[<�X<��U<B�R<&�O<X-M<��K<�K<L�K<�M<J[P<�}S<��V<�rY<�k[<MQ\<�\<�Z<��X<y�V<�oU<o�T<3U<��V<5�X<]�Z<��\<L/^<jp^<ǔ]<��[<T�Y<UmW<��U<�T<NU<�@V<X<�Z<:�[<=p\<�\<^�Z<KX<HU<M�Q<��N<-�L<ChK<XK<�}L<��N<�Q<��T<��W<�fZ<@
\<��\<��[<�nZ<�uX<-�V<�NU<qU<��U<7_W<��Y<�[<��]<Б^<�p^<�<]<+E[<��X<�V<>wU<��T<�xU<I�V<��X<��Z<� \<��\<�[<:�Y<�.W<	T<�P< "N<�+L<YJK<��K<[&M<�O<ߞR<��U<C�X<F[<�U\<�t\<�[<��Y<��W<
V<�U<�U<H0V<!	X<(GZ<�o\<�^<<�^<�%^<~�\<��Z<�DX<�ZV<0U<�U<��U<��W<��Y<�T[<c\<�d\<?[<=Y<�)V<y�R<Q�O<Y^M<��K<AK<� L<K�M<��P<թS<'�V<��Y<��[<�w\<A5\<��Z<_Y<�W<
�U<��T<�VU<<�V<��X<� [<�]<U^<2�^<J�]<��[<u�Y<V�W<3�U<�U<]1U<�\V<�4X<�2Z<�[<m�\<l \<�Z<4#X<VU<y�Q<��N<��L<�cK<�PK<esL<I�N<�{Q<��T<��W<"NZ<!�[<�o\<]�[<hLZ<�PX<QkV<�%U< �T<��U<!2W<�YY<o�[<�i]<�b^<�A^<M]<S[<��X<��V<}KU<��T<�MU<��V<#�X<��Z<I�[<$V\<��[<��Y<&�V<�S<��P<��M<��K<�K<�mK<�L<�bO<diR<��U<ēX<��Z< \<v>\<`J[<D�Y<��W<��U<\�T<�T<��U<x�W<�Z<�0\<��]<Pg^<_�]<�g\<[JZ<o	X<� V<��T<�  �  �S<!�S<��U<�W<3�Y<�[<�H[<�8Z<"X<��T<��Q<h>N<��K<A�I<�8I<J<qL<�N<�SR<�U<��X<b�Z<k^[<��Z<PqY<�WW<y3U<^�S<�S<W�S<�jU<;�W<w�Z<K]<��^<��^<W�]<m�[<+!Y<zV<aT<\@S<�KS<NwT<�nV<w�X<4vZ<�i[<|0[<F�Y<�4W<
�S<͍P<dM<��J<f�I<ށI<@�J<�M<�8P<&�S<a�V<%�Y<�,[<p�[<0�Z<m�X<H�V<��T<-�S<ZS<�\T<�_V<e�X<}�[<.�]<B_<B�^<p]<%[<�[X<�U<� T<�>S<��S<�$U<|@W<xcY<�Z<��[<��Z<�Y<�>V<=�R<pO<�L<�eJ<ErI<��I<�tK<~N<-`Q<o�T<��W<�;Z<�n[<4c[<�6Z<�BX<�V<�=T<�OS<8�S<��T<�/W<��Y<J|\<�^^<�_<@�^<��\<�2Z<[xW< U<��S<�DS<�T<�U<\X<�Z<�K[<z[<jZ<65X<�*U<��Q<\oN<��K<��I<�hI<27J<�9L<�O<mR<N�U<��X<ԻZ<��[<�[<��Y<:{W<�VU<��S<k7S<'�S<F�U<	X<��Z<�0]<߻^<�_<�^<��[<nEY<@�V<̂T<l`S<�iS<a�T<��V<ݹX<�Z<|[<@[<	�Y<�>W<T<��P<UeM<+�J<׎I<dzI<ݴJ<�M<~(P<-�S<��V<�yY<|[<�n[<�Z<��X<l�V<��T<S\S<�/S<�0T<s2V<E�X<��[<�]<�^<R�^<�A]<:�Z<[.X<��U<2�S<�S<@�S<h�T<�W<�8Y<��Z<�^[<u�Z<4�X<�V<��R<�MO<-SL<�1J<�=I<؜I<�?K<8�M<�*Q<�T<G�W<SZ<9[<-[<��Y<7X<�U<iT<�S<]NS<��T<��V<�Y<!=\<G^<j�^<�D^<�~\<��Y<�<W<��T<iS<�  �  kg><�?<�uB<;XF<�fJ<+�M<^�O<��O<D3N<�?K<R�G<Y�C<|@<:k><��=<>�><�A<�D<mbH<GL<H�N<X�O<�[O<zM<��I<�vE<�A<1:?<Zq><%�?<�{B<��F<�:K<QHO<z�Q<_R<}�P<**M<T�H<>D<��@<U�><�><�@<V�C<��G<ҾK<ئN< �O<��O<zM<�1J<\F<�B<��?<I5><� ><[�?<1VB<�E<��I<�:M<t{O< P<Y�N<X?L<�lH<0ZD<N�@<!�><��><�@<��C<f]H<"�L<ȉP<�xR<>7R<��O<��K<�OG<-C<��?<K�><�3?<8�A<�+E<�EI<��L<�YO<CP<�O<m�L<�H<� E<ܥA<�'?<><q{><�e@<u�C<UJG<�K<3#N<��O<x�O<�7N<�K<DG<C<N@<[�><+?<,�A<WE<��I<D;N<�eQ<�R<��Q<&�N<�eJ<��E<J�A<�U?<��><S�?<��B<ŋF<c�J<�M<��O<4�O<�dN<0qK<ԵG<��C<��@<m�><a><�><�LA<e�D<^�H<�+L<��N<sP<{�O<�?M<�I<��E<��A<$]?<��><9�?<��B<��F<^aK<�oO<[R<6�R<��P<�QM<$�H<�cD<��@<��><t�><%�@<	�C<��G<1�K<f�N<�P<l�O<ÄM<�9J<�`F<��B<q�?<�0><)><��?<ZHB<)�E<�I<�#M<�aO<xP<��N<RL<;HH</3D<�@<��><~�><Rd@<��C<�,H<��L<'XP<GR<,R<a�O<W�K<<!G<��B<��?<v><,	?<bA<�E<�I<��L<�-O<F�O<v�N<�ZL<�H<��D<^rA<<�><��=<�E><�/@<tKC<[G<
�J<S�M<��O<L�O<?N<U�J<�F<��B<��?<%p><g�><GA<�E<��I<J�M<�#Q<�_R<bQ<�gN<�&J<5�E<n�A<�?<�  �  �b?<�@<�eC<�.G<�K<0JN<�P<?)P<�N<��K<�H<�KD<#(A<�"?<�><4x?<I�A<�E<��H<�kL<BO<�NP<��O<�M<�KJ<7SF<�B< 8@<xj?< z@<<?C<�9G<��K<�{O<��Q<�kR<d�P<SxM<�2I<��D<3�A<ڲ?<��?<'zA<��D<H�H<�gL<N.O<�kP<@�O<��M<m�J<��F<�LC<�}@<��><��><�D@<8�B<+�F<�NJ<ğM<��O<��P<{�O<9�L<�4I<�?E<�A<��?<�?<oA<�D<E�H<�5M<��P<?�R<HR<*P< DL<��G<%�C<��@<�?<�1@<��B<jF<JJ<'�M<��O<'�P<�uO<��L<Y{I<H�E<FLB<��?<s�><�3?<�A<D<�G<.�K<��N<EP<�`P<5�N<i�K<�G<y D<vA<��?<$@<�VB<��E<�XJ<Y~N<ӀQ<խR<��Q<��N<�J<0sF<��B<)A@<�?<I�@<��C<bG<*NK<|N<EP<�ZP<X�N<��K<09H<?}D<�YA<,T?<�><+�?<+�A<$GE<�I<�L<;O<�uP<��O<}�M<�oJ<GvF<��B<[@<�?<4�@<"dC<^_G<+�K<�O<gR<��R<\�P<ܟM<YYI<GE<[�A<>�?<��?<B�A<S�D<X�H<�}L<�AO<w|P<��O<_�M<�J<G�F<xNC<n|@<��><��>< :@<b�B<MuF<�:J<�M<��O<oP<&bO<9�L<I<�E<��A<��?<�?<b@A<7}D<{�H<2M<�}P<�TR<R<��O<�L<I�G<�C<��@<�m?<@@<�WB<I�E<��I<"_M<٫O<UP<QGO<+�L<2JI<ԀE<�B<+�?<0�><�><��@<��C<�G<9LK<�NN<&P<�*P<��N<#�K<�G< �C<��@<dl?<��?<�B<^�E<�J<<N<�>Q<�kR<>zQ<9�N<�J<�5F<�qB<?@<�  �  �(B<�bC<�F<��I<n	M<C�O<tEQ<N*Q<��O<��L<glI<�E<�C<�/A<ɣ@<�~A<2�C<�F<�5J<��M<ZP<�VQ<�Q<QO<�PL<��H<�`E<BC<p)B<��B<\E<�H<.�L<��O<�R<�}R<$Q<=N<F�J<R�F<
�C<�\B<�{B<�:D<Z;G<��J<�1N<�P<ÈQ<��P<�N<Q�K<WcH<�E<�sB<RA<��@<P?B<�D<�
H<��K<ӪN<U�P<y�Q<V�P<Y�N<�[K<��G<��D<)�B<�tB<��C<�F<JJ<E	N<|Q<��R<�eR<�tP<E7M<�gI<@�E<�WC<�SB<��B<
5E<{H<�L<�1O<�"Q<�Q<pP<GN<,�J<�GG<D D<��A<��@<�CA<0�B<��E<!=I<�L<��O<�CQ<s�Q<~AP<�M<B J<řF<��C<qB<R�B<�D<��G<ÍK<�$O<�Q<��R<"�Q<�}O<E�K<*H<��D<��B<�`B<�C<<;F<�I<�;M<+P<wQ<�[Q<�O<�M<<�I<(F<�?C<LaA<��@<�A<o�C<�F<gbJ<w�M<u6P<(~Q<�>Q<�uO<�tL<��H<��E<S(C<�LB<�!C<�E<��H<��L<	 P<9=R<��R<�BQ<_dN<ٯJ<��F<D<:B<�B<�XD<�VG<��J<�GN<��P<X�Q<��P<��N<��K<�gH<YE<>rB<��@<�@<�4B<�D<��G<�yK<	�N<��P<��Q<�P<k�N<7K<�G<nD<�B<	HB<�C<IpF<bJ<�M<�P<PiR<�4R<`DP<�M<�9I<
�E<�+C<L(B<��B<�
E<�PH<[�K<vO<l�P<�aQ<oAP<6�M<��J<�G<Z�C<�A<f�@<�A<��B<��E<�I<�vL<�OO<�Q<EUQ<�
P<�cM<1�I<�`F<*�C<&5B< xB<:[D<�G<�LK<]�N<.zQ<
{R<�Q<�=O<u�K<��G<�D< �B<�  �  �3F<�qG<��I<M�L<��O<��Q<4�R<^R<)�P<}LN<�QK<CUH<��E<%>D<��C<��D<tTF<��H<5L<I�N< >Q<G�R<-�R<�oQ<yO<�!L<�>I<$G<�(F<��F<-SH<��J<�M<�tP<R<aR<�SQ<gO<�EL<SoI<JBG<>9F<��F<�9H<y�J<��M<|�P<y_R<s�R<eR<�,P<~yM<pqJ<t�G<�XE<mD<�D<�,E<�PG<O&J<[3M<:�O<PR<r�R<f�R<J�P<!ZN<�TK< �H<�F<�ZF<Q@G<1SI<ML<�O<�OQ<<�R<�YR<��P<�^N<pK<e�H<A�F<�KF<G<�I<W�K<�N<xbQ<��R<��R<*�Q<�eO<%�L<I<�F<��D<mD<nWD<T�E<�;H<20K<-1N<S�P<^tR<��R<,R<�(P<.UM<�UJ<��G<�F<�zF< �G<X/J<CM<u�O<^�Q<l�R<��Q<�P<�iM<}J<	H<h�F<�kF<��G<vJ<��L<)�O<��Q<��R<��R<��P<z~N<�K<��H</	F<JpD<[�C<}�D<A�F<(I<*.L<�O<�gQ<=�R<��R<�Q<�<O<IEL<�aI<Y=G<ELF<��F<�wH<5K<nN<��P<�9R<��R<{Q<}FO<�kL<��I<fG<<[F<��F<ZWH<��J<��M<��P<�rR<��R<�$R<V7P<�M<�uJ<�G<+WE<�D<+D<�!E<�BG<}J<�M<~�O<��Q<�R<9zR<y�P<�5N<�-K<wH<,�F</.F<G<�#I<��K<��N<�Q<,QR<;)R<��P<�/N<�AK<A�H<�F<1 F<J�F<=�H<��K<6�N<�6Q<�R<�R<pQ<'5O<2VL<�KI<��F<R�D<h�C<� D<��E<�H<��J<��M<)�P<E>R<��R<��Q<��O<QM<�J<��G<hDF<�=F<�G<��I<��L<��O<-�Q<`ZR<
�Q<C�O<�+M<E@J<��G<UF<�  �  ;�J<p�K<��M<�:P<�AR<�S<��S<�5S<ٳQ<O�O<�6M<��J<WI<��G<�uG<QH<<`I<CeK<��M<bP<#R<�sS<�S<X^S<�Q<��O<~M<էK<b�J<ɎJ<�qK<+M<3�N<��P<;�Q<=�Q<Q<��O<5�M<�L<Z�J<�J<= K<��L<q�N<Q<w�R<o�S<*�S<��R<�/Q<��N<�L<[J<��H<Y�G<�G<��H<�*J<XL<g�N<]Q<��R<��S<]T<�+S<mQ<�0O<�M<�hK<��J<�J<�L<d�M<�O<)+Q<��Q<��Q<!�P<�BO<sdM<��K<��J<��J<d�K<kM<��O<��Q<�hS<>T<��S<�yR<��P<�7N<2�K<g�I<MSH<��G<*�G<�I<f�J<�(M<8�O<��Q<QIS<�T<��S<��R< �P<�gN<�^L<	K<��J<�:K<Y�L<qN<9P<%�Q<	R<��Q<'eP<ťN<��L<rXK<�J<}�J<(,L<&N<)nP<qtR<��S<�T<hgS<��Q<��O<�iM<�K<U4I<�H<Y�G<�2H<ŐI<y�K<��M<bHP<fFR<�S< T< �S<�R<l�O<�M<8�K<�J<�J<N�K<�+M<\	O<D�P<c�Q<��Q<�DQ<��O<$N<�?L<�K<��J<�?K<|�L<��N<�)Q<m�R<��S<��S<.�R<%:Q<z�N<f�L<�\J<��H<��G<g�G<ǁH<�J<IGL<��N<��P<�R<d�S<P�S<A
S<�HQ<
O<��L<@>K<�J<(�J<��K<Z�M<M}O<S�P<��Q<G�Q<d�P<�O<r6M<ԓK<W�J<��J<}{K<[@M<�|O<��Q<�<S<<�S<T�S<�IR<�YP<�N<H�K<W�I<TH<WyG<'�G<��H<P�J<��L<�VO<=}Q<S<y�S<y�S<pR<gxP<&/N<�$L<�J<pgJ<\�J<�_L<1N<��O<�AQ<��Q<�ZQ<A&P<hN<��L<�K< nJ<�  �  �N<�P<�Q<��R<T<dcT<�T<HS<��Q<a3P<��N<E#M<��K<KK<~K<�hK<N7L<rqM<��N<��P<�R<�bS<�2T<�dT<��S<g�R<�7Q<��O<~�N<�N<]	N<�~N<�6O<��O<�`P<�wP<�*P<�O<��N<C7N<�N<�XN<�?O<b�P<t#R<��S<TVT<wT<��S<��R<.fQ<�O< :N<v�L<��K<~TK<�NK<��K<u�L<�N<�O<�JQ<��R<�S<��T<V�T<H�S<8qR<��P<��O<��N<0N<�WN<��N<K�O<�IP<��P<$�P<�'P<�wO<f�N<�:N<	/N<��N<��O<�3Q<��R<��S<�T<�kT<'�S<�sR<z�P<RO<��M<4�L<��K<vPK<�uK<L<5M<$�N<W;P<[�Q<�2S<�-T<�T<JNT<7VS<��Q<{cP<b!O<H[N<�'N<8yN<�"O<�O<�nP<<�P<�yP<��O<t7O<�N<�)N<�LN<�O<79P<�Q<�/S<�8T<��T<�>T<QS<�Q<MfP<��N<�VM<�2L<�~K<�JK<�K<�hL<��M<M!O<O�P<�GR<݋S<HZT<�T<�T<��R<�[Q<��O<<�N<�1N<
.N<�N<�\O<7P<m�P<�P<oQP<δO<p�N<�[N<�%N< zN<Z_O<��P<T>R<�S<lT<"�T<��S<�R<�pQ<��O<p>N<��L<��K<�OK<�FK<�K<��L<
N<m�O<a4Q<F�R<��S<�jT<�^T<S�S<�JR<�P<�^O<�hN<kN<�(N<�N<wO<�P<@qP<eP<f�O<�HO<��N<�N<�N<5�N<��O<	Q<{�R<A�S<r\T<>T<A~S<�CR<��P<�O<)�M<dTL<�xK<#K<>K<Y�K<s�L<�jN<aP<��Q<V�R<��S<�`T<�T<�S<��Q<K*P<�N<�N<�M<O;N<�N<��O<8/P<�gP<�:P<��O<�N<WLN<��M<�N<�  �  ��Q<|�R<|�S<VT<RT<ƽS<��R<x�Q<�P<H�O<�O<ݖN< UN<5N<�,N<B:N<FaN<<�N<�(O<�O<��P<�Q<1	S<k�S<�gT<�JT<��S<+�R<��Q<C{P<��O<3�N<��N<\N<	AN<=N<�NN<X{N<�N<�TO<�P<1Q<�2R<�GS<L T<�T<LT<��S<��R<�nQ<iP<��O<� O<L�N<soN<tYN<�YN<LpN<i�N<��N<ڏO<�_P<�cQ<��R<n�S<<ZT<�T<nTT<��S<�yR<�]Q<�]P<!�O<�O<n�N<,N<�jN<lN<��N<��N<qO<�O<��P<��Q<�R<ܱS<gT<t�T<�-T<3RS<�=R<!$Q<�,P<
mO<��N<8�N<�sN<�dN<�jN<��N<*�N<�.O<��O<��P<%�Q<��R<��S<�|T<C�T<�T<�*S<>R<�P<�P<QWO<0�N<y�N<�rN<�fN<&pN<e�N<��N<PFO<x�O<��P<�Q<�S<j�S<)�T<��T<	�S<��R<�Q<��P<��O<�:O<-�N<��N<{iN<�`N<�mN<��N<6�N<2XO<�P<�Q<R<�1S<AT<�T<^oT<��S<��R<��Q<h�P<+�O<X"O<��N<'�N<|gN<�cN<�tN<5�N<�N<�xO<v<P<7Q<�QR<}dS<�:T<��T<�aT<��S<њR<�{Q<SsP<��O<�O<��N<�mN<�TN<*RN<�eN<��N<��N<:|O<NIP<�JQ<fR<�rS<�8T<4T<f.T<[`S<�OR<�1Q<�0P<�dO<q�N<�N< ON<�:N<V<N<wTN<�N<��N<�O<\P<�dQ<�R<��S<�;T<eiT<� T<$S<R<�P<��O<�8O<%�N<�fN<L<N<�,N<d2N<_ON<��N<��N<]�O<�|P<��Q<��R<T�S<XFT<P[T<I�S<V�R<��Q<.�P<��O<?O<J�N<YN<4N<b(N<2N<TN<Y�N<wO<�O<�P<�  �  �-S<\T<^bT<;�S<7�R<�pQ<�O<ֿN<�N<b�M<xWN<�O<��O<�CP<�kP<.P<"�O<�N<	:N<��M<�-N<��N< GP<%�Q<�9S<c*T<�iT<8�S<��R<r�Q<5�O<�bN<}�L<��K<�GK<+K<��K<huL<��M<WHO<��P<�kR<C�S<{YT<�nT<1�S<R�R<8Q<�O<3�N<�N<�,N<��N<�oO<{P<8�P<w�P<�1P<��O<��N<�DN<(&N<�N<��O<��P<��R<��S<��T<!�T<��S<G�R</?Q<��O<�N<2�L<��K<�\K<SjK<��K<� M<caN<C�O<m�Q<]�R<6
T<ƍT<�cT<�S<H%R<��P<MKO<�mN<S"N<�_N<m�N<��O<�XP<
�P<օP<P<VVO<<�N<�0N<�<N<��N<$�O<QyQ<X�R<ET<H�T<[T<��S<q;R<D�P<XO<,�M<&aL<��K<PK<׊K<�DL<9nM<��N<��P<�R<�cS<IT<�T</.T<�S<	�Q<�#P<��N<KDN<b(N<�N<�=O<��O<*yP<��P<RbP<]�O<O<XjN<RN<�ZN<n(O<pP<��Q<�_S<|OT<�T<DT<�S<��Q<�P<��N<�M<�L<nK<7QK<��K<ԚL<+�M<�kO<�	Q<�R<�S<vT<��T<�S<��R<�Q<�O<O�N<$N<4N<ضN<qO<�P<��P<P<�&P<�~O<3�N<1N<�N<�{N<�vO<[�P<~bR<u�S<�aT<BaT<ʹS<܏R<YQ<�sO<�M<ϒL<'�K< -K< ;K<��K<��L<�3N<��O<UbQ<��R<��S<WbT<�7T<�YS<��Q<�nP<O<<N<��M<�*N< �N<:�O<� P<1iP<�LP<	�O<�O<�gN<�M<�N<M�N<��O<4CQ<�R<��S<^T<�"T<�KS<AR<tP<�N<&XM<�#L<�[K<aK<�MK<�L<�2M<ܪN<�GP<��Q<�  �  jCS<��S<�S<�(R<�P<��M<=�K<�J<�sJ<�0K</�L<�N<�?P<GjQ<�Q<*9Q<:�O<ZN<NL<y�J<8mJ<��J<FL<�WN<�P<�R<ѶS<�S<=S<nQ<NBO<I�L<��J<~�H<�G<��G<�=H<��I<��K<�9N<�P<�tR<�S<�S<�AS<T�Q<asO<�:M<��K<ܞJ<}�J<A�K<lM<�IO<#�P<��Q<��Q<�Q<X�O<��M<�K<��J<,�J<�rK<%M<TNO<~�Q<X@S<T<��S<��R<��P<R�N<jDL<J<�H<i�G<��G<m�H<��J<p�L<�(O<�^Q<�S<�S<��S<p�R<&	Q<�N<;�L<-K<�J<jK<TTL<�N<��O<�TQ<��Q<��Q<ѢP<��N<�M<p�K<ͳJ<��J<h�K<z�M<\P<�)R<��S<�T<�S< 6R<0P<��M<|K<PI<�+H<A�G<�H<�OI<=K<��M<|�O<�R<�xS<OT<e�S<�[R<kMP<XN<�L<O�J<��J<1eK<Z�L<��N<�uP<U�Q<��Q<EnQ<RP<ON<-L<�$K<��J<&K<�oL<�N<��P<n�R<��S<OT<V1S<>�Q<�fO<M<̾J<�H<��G<\�G<cH<��I<�K<!]N<��P<�R<��S<iT<�[S<�Q<��O<mMM<h�K<ګJ<��J<x�K<UpM<5KO<n�P<��Q<?�Q<��P<�vO<�M<��K<~�J<
�J<�VK<��L<^-O<)fQ<�S<��S<-�S<l�R<+�P<�{N<�L<�I<�[H<(�G<��G<�H<�[J<(�L< �N<z2Q<��R<��S<9�S<N�R<=�P<�N<�wL<6�J<�kJ<I�J<�L<��M<x�O<�Q<5�Q<�~Q<.iP<��N<��L<fRK<s|J<��J<"�K<t�M<U�O<V�Q<$dS<�S<j^S<z�Q<��O<\�M<�?K<�BI<��G<ipG<W�G<KI<`K<DVM<T�O<��Q<�  �  1jR<[�R<޳Q<݄O<ҜL<?�I<�XG<�-F<{cF<��G<8kJ<�XM<wP<��Q<]R<D�Q<P|O<��L<5�I<�{G<�;F<�VF<A�G<!NJ<�QM<P<R<A�R<59R<�xP<��M<��J<��G<f�E<�#D<��C<��D<*�F<�I<�L<�mO<�Q<��R<��R<�0Q<��N<!�K<��H<��F<�8F<��F<��H<�K<�sN<��P<qRR<�gR<�#Q<B�N<��K<Z!I<�G<NF<�F<p�H<m{K<[�N<FQ<�R<1�R<��Q<��O<cM<�J<<;G<�$E<D<V8D<��E<��G<x�J<;�M<{`P<~=R<w�R<qbR<��P<�M<y�J<�4H<a�F< ^F<�{G<9�I<L�L<�kO<�Q<��R<.R<-�P<h�M<��J<�^H<�F<�WF<x\G<��I<lyL<RlO<U�Q<��R<иR<�TQ<�N<r
L<I<�jF<ԦD<��C</�D<B,F<9�H<$�K<X�N<�Q<\�R<y�R<(�Q<��O<P�L<��I<��G<caF<��F<�H<�J<ώM<<P<�
R<��R<�Q<(�O<�L<J<��G<�iF<�F<|�G<�vJ<�xM<�DP<9R<��R<g]R<�P<7N<P K< H<��E<ID<(D<��D<��F<�I<жL<�O<˼Q<��R<��R<}JQ<%�N<�K<�H<f�F<�EF<��F<�H<M�K<$uN<��P<�MR<�_R<�Q<��N<
�K<�I<?G<5F<Z�F<�H<�ZK<1_N<��P<�R<��R<$�Q<z�O<�L<x�I<�G<��D<�C<�	D<oUE<֛G<W�J<��M<o4P<�R<��R<�6R<$aP<٤M<�J< H<�mF<+F<GG<�I<�]L<�2O<CZQ<�UR<��Q<FP<��M<лJ<Y&H<�~F<!F<.&G<�YI<�CL<I6O<ـQ<өR<̀R<�Q<3�N<��K<��H<�.F<�jD<��C<wID<@�E<-zH<=zK<�qN<i�P<�  �  �4Q<�9Q<��O<�L<�MI<"�E<
HC<s%B<"�B<�D<'$H<��K<�lO<^�Q<7}R<�cQ<��N<K<WG<)=D<�oB<�EB<x�C<�F<s%J<M<�1P<�fQ<�	Q<:O<sUL<�H<9yE<�B<�A<k�@<�A<�%D<�WG<��J<�N<	oP<&{Q<�P<-�N<��K<�5H<��D<%�B<�DB<]`C<��E<|�I<XM<&�P<�aR<�|R<��P<��M<ZJ<=bF<ܩC<cB<�B<~�D<c�G<��K<S�N<��P<�Q<��P<V�N<<hK<��G<�D<Z3B<��@<�A<�B<JE<�H<� L<�O<�Q<A�Q<Z�P<yN<*�J<�#G<g3D<��B<��B<4+D<�(G<�J<��N</cQ<��R<@-R<^�O<��L<�H<]E<C<pUB<�HC<��E<3I<�L<Q�O<�UQ<R~Q<A"P<��M<F8J<U�F<��C<?�A<1�@<�xA<�gC<2[F<�I<d4M<��O<piQ<�mQ<��O<�M<�I<�F<{C<YB<��B<bE<;ZH<w*L<�O<��Q<=�R<-�Q<��N<PK<��G<�mD<t�B<UrB<�C<��F<�LJ<��M<�VP<��Q<�-Q<8^O<�yL<�I<�E<�B<33A<��@<��A<�ID<q{G<Z�J<5N<��P<��Q<�Q<�O<��K<�JH<0E<��B<�QB<\jC<�E<��I<UYM<h�P<�\R<IuR<;�P<D�M<��I<�NF<��C<"JB<ԮB<@�D<��G<�iK<�N<��P<�}Q<�P<aaN</;K<�G<�tD<�B<��@<.�@<�tB<�E<zH<<�K<��N<��P<mQ<QdP<��M<��J<$�F<7D</ZB<TB<��C<��F<ԭJ<�[N< )Q<�sR<{�Q<��O<�^L<��H<~$E<M�B<�B<mC<��E<}�H<7xL<kO<�Q<�FQ<��O<SM< �I<\F<LuC<�dA<��@<�=A<Q-C<�!F<��I<"�L<ۯO<�  �  �1P<�P<'$N<-�J<7�F<�5C<}@<�`?<v @<p�B<�tF<z�J<a�N<��Q<�mR<�#Q<AN<G�I<ǈE<��A<��?<�{?<��@<hD<��G<�K<��N<@P<OP<Q7N<�'K<qG<��C<��@<K�><��><�?<UB<��E<�I</M<3uO<8lP<�O<8JM<��I<��E<qEB<W@<ƌ?<0�@<��C<FH<�lL<�P<�FR<�fR<3uP<?�L<R�H<hD<�>A<(�?<��?<$B<gqE<'kI<�M<��O<��P<��O<�M<�%J<B]F<��B<m6@<��><�?<~�@<��C<@.G<+�J<6N<9P<+yP<�$O<�LL<t�H<Q�D<qA<��?<��?<Q�A<�KE<��I<�M<�Q< �R<R<�wO< �K<�'G<�9C<�@<��?<*|@<�C<�F<k�J<
N<�P<�wP<6&O<apL<��H<�E<s�A<��?<�><"m?<��A<�D<�rH<�L<'�N<�fP<�7P<5WN<�K<�'G<�hC<7�@<��?<U@<��B<�F<|K<�O<!�Q<�R<lZQ<	BN<�J<��E<�$B<��?<��?<y(A<�+D<
H<2�K<��N<�dP<�0P<�[N<�KK<��G<��C<��@<g"?<��><��?<KyB<&�E<k�I<=#M<��O<�P<��O<�cM<��I<��E<�WB<�@<��?<$�@<��C<oH<�mL<�P<�AR<�^R<�jP<��L<̓H<�TD<�(A<4�?</�?<��A<�PE<2HI<��L<�wO<�iP<W�O<6TM<��I<�/F<��B<�@<��><h�><��@<`C<OG<��J<0�M<m�O<YMP<��N<�L<�RH<bgD<�@A<�?<)�?<ȠA<wE<m_I<\�M<!�P<cR<�Q<�<O<�RK<+�F<� C<9R@<�]?<�E@<�B<y�F<�xJ<u�M<��O<�@P<��N<@7L<	�H<
�D<W�A<_\?<ǅ><I2?<sJA<�zD<�:H<��K<S�N<�  �  ��O<O�O<H�M<k/J<%F<�DB<�?<f><"6?<�A<��E<!kJ<v�N<��Q<�aR<�Q<*�M<sfI<��D<� A<p�><>><�@<"C<zG<K</N<��O<��O<��M<U�J<?�F<J'C< @<�D><m�=<�?<ȯA<�6E< I<��L<\O<�P<�+O<�L<Z�H<��D<�NA<??<ϕ><
@<3C<�}G<1L<��O<�6R<:XR<`MP<�L<�H<�C<a@<Ѻ><��><�A<Z�D<8�H<�oL<O<(P<�lO<M<ìI<��E<�5B<C�?<�'><�R><9�?<��B<�F<�wJ<@�M<c�O<[
P<��N<�K<�G<��C<lv@<y�><��><��@<��D<�I<��M<��P<��R<��Q<BO<i&K<f�F<�sB<��?<ʚ><c~?<�B<��E<��I<�rM<�O<oP<�N<�L<2_H<��D<*A<"�><r><��><X�@<�D<��G<�K<��N<�P<	�O<N�M<bJ<�OF<xwB<�?<�><�j?<�B<]F<=�J<�N<b�Q</�R<�=Q<�M<�I<�E<�QA<z?<;�><�,@<R?C<9G<l6K<nTN<}�O<��O<��M<��J<�G<LC<?@<�i><i><gC?<��A<$ZE<P9I<��L<�4O<8!P<eGO<��L<�I<w�D<aA<�?<��><�@<':C<#�G<fL<��O<�1R<�PR<�BP<y�L<�G<��C<�J@<�><2�><��@<�lD<J�H<�JL<��N<?�O<_BO<W�L<�I<�E<�B<�T?<�=<G$><H�?<V�B<xF<`KJ<;�M<��O<��O<ioN<uK<T�G<�}C<�E@<P�><��><2�@<IfD<��H<�RM<�P<�VR<��Q<+O<	�J<�TF<	;B<�j?<�c><H?<��A<a�E<:�I<�<M<wgO<#�O<ލN<��K<[%H<4JD<�@<�><T�=<{><G�@<��C<��G<nK<�QN<�  �  �1P<�P<'$N<-�J<7�F<�5C<}@<�`?<v @<p�B<�tF<z�J<a�N<��Q<�mR<�#Q<AN<G�I<ǈE<��A<��?<�{?<��@<hD<��G<�K<��N<@P<OP<Q7N<�'K<qG<��C<��@<K�><��><�?<UB<��E<�I</M<3uO<8lP<�O<8JM<��I<��E<qEB<W@<ƌ?<0�@<��C<FH<�lL<�P<�FR<�fR<3uP<?�L<R�H<hD<�>A<(�?<��?<$B<gqE<'kI<�M<��O<��P<��O<�M<�%J<B]F<��B<m6@<��><�?<~�@<��C<@.G<+�J<6N<9P<+yP<�$O<�LL<t�H<Q�D<qA<��?<��?<Q�A<�KE<��I<�M<�Q< �R<R<�wO< �K<�'G<�9C<�@<��?<*|@<�C<�F<k�J<
N<�P<�wP<6&O<apL<��H<�E<s�A<��?<�><"m?<��A<�D<�rH<�L<'�N<�fP<�7P<5WN<�K<�'G<�hC<7�@<��?<U@<��B<�F<|K<�O<!�Q<�R<lZQ<	BN<�J<��E<�$B<��?<��?<y(A<�+D<
H<2�K<��N<�dP<�0P<�[N<�KK<��G<��C<��@<g"?<��><��?<KyB<&�E<k�I<=#M<��O<�P<��O<�cM<��I<��E<�WB<�@<��?<$�@<��C<oH<�mL<�P<�AR<�^R<�jP<��L<̓H<�TD<�(A<4�?</�?<��A<�PE<2HI<��L<�wO<�iP<W�O<6TM<��I<�/F<��B<�@<��><h�><��@<`C<OG<��J<0�M<m�O<YMP<��N<�L<�RH<bgD<�@A<�?<)�?<ȠA<wE<m_I<\�M<!�P<cR<�Q<�<O<�RK<+�F<� C<9R@<�]?<�E@<�B<y�F<�xJ<u�M<��O<�@P<��N<@7L<	�H<
�D<W�A<_\?<ǅ><I2?<sJA<�zD<�:H<��K<S�N<�  �  �4Q<�9Q<��O<�L<�MI<"�E<
HC<s%B<"�B<�D<'$H<��K<�lO<^�Q<7}R<�cQ<��N<K<WG<)=D<�oB<�EB<x�C<�F<s%J<M<�1P<�fQ<�	Q<:O<sUL<�H<9yE<�B<�A<k�@<�A<�%D<�WG<��J<�N<	oP<&{Q<�P<-�N<��K<�5H<��D<%�B<�DB<]`C<��E<|�I<XM<&�P<�aR<�|R<��P<��M<ZJ<=bF<ܩC<cB<�B<~�D<c�G<��K<S�N<��P<�Q<��P<V�N<<hK<��G<�D<Z3B<��@<�A<�B<JE<�H<� L<�O<�Q<A�Q<Z�P<yN<*�J<�#G<g3D<��B<��B<4+D<�(G<�J<��N</cQ<��R<@-R<^�O<��L<�H<]E<C<pUB<�HC<��E<3I<�L<Q�O<�UQ<R~Q<A"P<��M<F8J<U�F<��C<?�A<1�@<�xA<�gC<2[F<�I<d4M<��O<piQ<�mQ<��O<�M<�I<�F<{C<YB<��B<bE<;ZH<w*L<�O<��Q<=�R<-�Q<��N<PK<��G<�mD<t�B<UrB<�C<��F<�LJ<��M<�VP<��Q<�-Q<8^O<�yL<�I<�E<�B<33A<��@<��A<�ID<q{G<Z�J<5N<��P<��Q<�Q<�O<��K<�JH<0E<��B<�QB<\jC<�E<��I<UYM<h�P<�\R<IuR<;�P<D�M<��I<�NF<��C<"JB<ԮB<@�D<��G<�iK<�N<��P<�}Q<�P<aaN</;K<�G<�tD<�B<��@<.�@<�tB<�E<zH<<�K<��N<��P<mQ<QdP<��M<��J<$�F<7D</ZB<TB<��C<��F<ԭJ<�[N< )Q<�sR<{�Q<��O<�^L<��H<~$E<M�B<�B<mC<��E<}�H<7xL<kO<�Q<�FQ<��O<SM< �I<\F<LuC<�dA<��@<�=A<Q-C<�!F<��I<"�L<ۯO<�  �  1jR<[�R<޳Q<݄O<ҜL<?�I<�XG<�-F<{cF<��G<8kJ<�XM<wP<��Q<]R<D�Q<P|O<��L<5�I<�{G<�;F<�VF<A�G<!NJ<�QM<P<R<A�R<59R<�xP<��M<��J<��G<f�E<�#D<��C<��D<*�F<�I<�L<�mO<�Q<��R<��R<�0Q<��N<!�K<��H<��F<�8F<��F<��H<�K<�sN<��P<qRR<�gR<�#Q<B�N<��K<Z!I<�G<NF<�F<p�H<m{K<[�N<FQ<�R<1�R<��Q<��O<cM<�J<<;G<�$E<D<V8D<��E<��G<x�J<;�M<{`P<~=R<w�R<qbR<��P<�M<y�J<�4H<a�F< ^F<�{G<9�I<L�L<�kO<�Q<��R<.R<-�P<h�M<��J<�^H<�F<�WF<x\G<��I<lyL<RlO<U�Q<��R<иR<�TQ<�N<r
L<I<�jF<ԦD<��C</�D<B,F<9�H<$�K<X�N<�Q<\�R<y�R<(�Q<��O<P�L<��I<��G<caF<��F<�H<�J<ώM<<P<�
R<��R<�Q<(�O<�L<J<��G<�iF<�F<|�G<�vJ<�xM<�DP<9R<��R<g]R<�P<7N<P K< H<��E<ID<(D<��D<��F<�I<жL<�O<˼Q<��R<��R<}JQ<%�N<�K<�H<f�F<�EF<��F<�H<M�K<$uN<��P<�MR<�_R<�Q<��N<
�K<�I<?G<5F<Z�F<�H<�ZK<1_N<��P<�R<��R<$�Q<z�O<�L<x�I<�G<��D<�C<�	D<oUE<֛G<W�J<��M<o4P<�R<��R<�6R<$aP<٤M<�J< H<�mF<+F<GG<�I<�]L<�2O<CZQ<�UR<��Q<FP<��M<лJ<Y&H<�~F<!F<.&G<�YI<�CL<I6O<ـQ<өR<̀R<�Q<3�N<��K<��H<�.F<�jD<��C<wID<@�E<-zH<=zK<�qN<i�P<�  �  jCS<��S<�S<�(R<�P<��M<=�K<�J<�sJ<�0K</�L<�N<�?P<GjQ<�Q<*9Q<:�O<ZN<NL<y�J<8mJ<��J<FL<�WN<�P<�R<ѶS<�S<=S<nQ<NBO<I�L<��J<~�H<�G<��G<�=H<��I<��K<�9N<�P<�tR<�S<�S<�AS<T�Q<asO<�:M<��K<ܞJ<}�J<A�K<lM<�IO<#�P<��Q<��Q<�Q<X�O<��M<�K<��J<,�J<�rK<%M<TNO<~�Q<X@S<T<��S<��R<��P<R�N<jDL<J<�H<i�G<��G<m�H<��J<p�L<�(O<�^Q<�S<�S<��S<p�R<&	Q<�N<;�L<-K<�J<jK<TTL<�N<��O<�TQ<��Q<��Q<ѢP<��N<�M<p�K<ͳJ<��J<h�K<z�M<\P<�)R<��S<�T<�S< 6R<0P<��M<|K<PI<�+H<A�G<�H<�OI<=K<��M<|�O<�R<�xS<OT<e�S<�[R<kMP<XN<�L<O�J<��J<1eK<Z�L<��N<�uP<U�Q<��Q<EnQ<RP<ON<-L<�$K<��J<&K<�oL<�N<��P<n�R<��S<OT<V1S<>�Q<�fO<M<̾J<�H<��G<\�G<cH<��I<�K<!]N<��P<�R<��S<iT<�[S<�Q<��O<mMM<h�K<ګJ<��J<x�K<UpM<5KO<n�P<��Q<?�Q<��P<�vO<�M<��K<~�J<
�J<�VK<��L<^-O<)fQ<�S<��S<-�S<l�R<+�P<�{N<�L<�I<�[H<(�G<��G<�H<�[J<(�L< �N<z2Q<��R<��S<9�S<N�R<=�P<�N<�wL<6�J<�kJ<I�J<�L<��M<x�O<�Q<5�Q<�~Q<.iP<��N<��L<fRK<s|J<��J<"�K<t�M<U�O<V�Q<$dS<�S<j^S<z�Q<��O<\�M<�?K<�BI<��G<ipG<W�G<KI<`K<DVM<T�O<��Q<�  �  �-S<\T<^bT<;�S<7�R<�pQ<�O<ֿN<�N<b�M<xWN<�O<��O<�CP<�kP<.P<"�O<�N<	:N<��M<�-N<��N< GP<%�Q<�9S<c*T<�iT<8�S<��R<r�Q<5�O<�bN<}�L<��K<�GK<+K<��K<huL<��M<WHO<��P<�kR<C�S<{YT<�nT<1�S<R�R<8Q<�O<3�N<�N<�,N<��N<�oO<{P<8�P<w�P<�1P<��O<��N<�DN<(&N<�N<��O<��P<��R<��S<��T<!�T<��S<G�R</?Q<��O<�N<2�L<��K<�\K<SjK<��K<� M<caN<C�O<m�Q<]�R<6
T<ƍT<�cT<�S<H%R<��P<MKO<�mN<S"N<�_N<m�N<��O<�XP<
�P<օP<P<VVO<<�N<�0N<�<N<��N<$�O<QyQ<X�R<ET<H�T<[T<��S<q;R<D�P<XO<,�M<&aL<��K<PK<׊K<�DL<9nM<��N<��P<�R<�cS<IT<�T</.T<�S<	�Q<�#P<��N<KDN<b(N<�N<�=O<��O<*yP<��P<RbP<]�O<O<XjN<RN<�ZN<n(O<pP<��Q<�_S<|OT<�T<DT<�S<��Q<�P<��N<�M<�L<nK<7QK<��K<ԚL<+�M<�kO<�	Q<�R<�S<vT<��T<�S<��R<�Q<�O<O�N<$N<4N<ضN<qO<�P<��P<P<�&P<�~O<3�N<1N<�N<�{N<�vO<[�P<~bR<u�S<�aT<BaT<ʹS<܏R<YQ<�sO<�M<ϒL<'�K< -K< ;K<��K<��L<�3N<��O<UbQ<��R<��S<WbT<�7T<�YS<��Q<�nP<O<<N<��M<�*N< �N<:�O<� P<1iP<�LP<	�O<�O<�gN<�M<�N<M�N<��O<4CQ<�R<��S<^T<�"T<�KS<AR<tP<�N<&XM<�#L<�[K<aK<�MK<�L<�2M<ܪN<�GP<��Q<�  �  ��Q<|�R<|�S<VT<RT<ƽS<��R<x�Q<�P<H�O<�O<ݖN< UN<5N<�,N<B:N<FaN<<�N<�(O<�O<��P<�Q<1	S<k�S<�gT<�JT<��S<+�R<��Q<C{P<��O<3�N<��N<\N<	AN<=N<�NN<X{N<�N<�TO<�P<1Q<�2R<�GS<L T<�T<LT<��S<��R<�nQ<iP<��O<� O<L�N<soN<tYN<�YN<LpN<i�N<��N<ڏO<�_P<�cQ<��R<n�S<<ZT<�T<nTT<��S<�yR<�]Q<�]P<!�O<�O<n�N<,N<�jN<lN<��N<��N<qO<�O<��P<��Q<�R<ܱS<gT<t�T<�-T<3RS<�=R<!$Q<�,P<
mO<��N<8�N<�sN<�dN<�jN<��N<*�N<�.O<��O<��P<%�Q<��R<��S<�|T<C�T<�T<�*S<>R<�P<�P<QWO<0�N<y�N<�rN<�fN<&pN<e�N<��N<PFO<x�O<��P<�Q<�S<j�S<)�T<��T<	�S<��R<�Q<��P<��O<�:O<-�N<��N<{iN<�`N<�mN<��N<6�N<2XO<�P<�Q<R<�1S<AT<�T<^oT<��S<��R<��Q<h�P<+�O<X"O<��N<'�N<|gN<�cN<�tN<5�N<�N<�xO<v<P<7Q<�QR<}dS<�:T<��T<�aT<��S<њR<�{Q<SsP<��O<�O<��N<�mN<�TN<*RN<�eN<��N<��N<:|O<NIP<�JQ<fR<�rS<�8T<4T<f.T<[`S<�OR<�1Q<�0P<�dO<q�N<�N< ON<�:N<V<N<wTN<�N<��N<�O<\P<�dQ<�R<��S<�;T<eiT<� T<$S<R<�P<��O<�8O<%�N<�fN<L<N<�,N<d2N<_ON<��N<��N<]�O<�|P<��Q<��R<T�S<XFT<P[T<I�S<V�R<��Q<.�P<��O<?O<J�N<YN<4N<b(N<2N<TN<Y�N<wO<�O<�P<�  �  �N<�P<�Q<��R<T<dcT<�T<HS<��Q<a3P<��N<E#M<��K<KK<~K<�hK<N7L<rqM<��N<��P<�R<�bS<�2T<�dT<��S<g�R<�7Q<��O<~�N<�N<]	N<�~N<�6O<��O<�`P<�wP<�*P<�O<��N<C7N<�N<�XN<�?O<b�P<t#R<��S<TVT<wT<��S<��R<.fQ<�O< :N<v�L<��K<~TK<�NK<��K<u�L<�N<�O<�JQ<��R<�S<��T<V�T<H�S<8qR<��P<��O<��N<0N<�WN<��N<K�O<�IP<��P<$�P<�'P<�wO<f�N<�:N<	/N<��N<��O<�3Q<��R<��S<�T<�kT<'�S<�sR<z�P<RO<��M<4�L<��K<vPK<�uK<L<5M<$�N<W;P<[�Q<�2S<�-T<�T<JNT<7VS<��Q<{cP<b!O<H[N<�'N<8yN<�"O<�O<�nP<<�P<�yP<��O<t7O<�N<�)N<�LN<�O<79P<�Q<�/S<�8T<��T<�>T<QS<�Q<MfP<��N<�VM<�2L<�~K<�JK<�K<�hL<��M<M!O<O�P<�GR<݋S<HZT<�T<�T<��R<�[Q<��O<<�N<�1N<
.N<�N<�\O<7P<m�P<�P<oQP<δO<p�N<�[N<�%N< zN<Z_O<��P<T>R<�S<lT<"�T<��S<�R<�pQ<��O<p>N<��L<��K<�OK<�FK<�K<��L<
N<m�O<a4Q<F�R<��S<�jT<�^T<S�S<�JR<�P<�^O<�hN<kN<�(N<�N<wO<�P<@qP<eP<f�O<�HO<��N<�N<�N<5�N<��O<	Q<{�R<A�S<r\T<>T<A~S<�CR<��P<�O<)�M<dTL<�xK<#K<>K<Y�K<s�L<�jN<aP<��Q<V�R<��S<�`T<�T<�S<��Q<K*P<�N<�N<�M<O;N<�N<��O<8/P<�gP<�:P<��O<�N<WLN<��M<�N<�  �  ;�J<p�K<��M<�:P<�AR<�S<��S<�5S<ٳQ<O�O<�6M<��J<WI<��G<�uG<QH<<`I<CeK<��M<bP<#R<�sS<�S<X^S<�Q<��O<~M<էK<b�J<ɎJ<�qK<+M<3�N<��P<;�Q<=�Q<Q<��O<5�M<�L<Z�J<�J<= K<��L<q�N<Q<w�R<o�S<*�S<��R<�/Q<��N<�L<[J<��H<Y�G<�G<��H<�*J<XL<g�N<]Q<��R<��S<]T<�+S<mQ<�0O<�M<�hK<��J<�J<�L<d�M<�O<)+Q<��Q<��Q<!�P<�BO<sdM<��K<��J<��J<d�K<kM<��O<��Q<�hS<>T<��S<�yR<��P<�7N<2�K<g�I<MSH<��G<*�G<�I<f�J<�(M<8�O<��Q<QIS<�T<��S<��R< �P<�gN<�^L<	K<��J<�:K<Y�L<qN<9P<%�Q<	R<��Q<'eP<ťN<��L<rXK<�J<}�J<(,L<&N<)nP<qtR<��S<�T<hgS<��Q<��O<�iM<�K<U4I<�H<Y�G<�2H<ŐI<y�K<��M<bHP<fFR<�S< T< �S<�R<l�O<�M<8�K<�J<�J<N�K<�+M<\	O<D�P<c�Q<��Q<�DQ<��O<$N<�?L<�K<��J<�?K<|�L<��N<�)Q<m�R<��S<��S<.�R<%:Q<z�N<f�L<�\J<��H<��G<g�G<ǁH<�J<IGL<��N<��P<�R<d�S<P�S<A
S<�HQ<
O<��L<@>K<�J<(�J<��K<Z�M<M}O<S�P<��Q<G�Q<d�P<�O<r6M<ԓK<W�J<��J<}{K<[@M<�|O<��Q<�<S<<�S<T�S<�IR<�YP<�N<H�K<W�I<TH<WyG<'�G<��H<P�J<��L<�VO<=}Q<S<y�S<y�S<pR<gxP<&/N<�$L<�J<pgJ<\�J<�_L<1N<��O<�AQ<��Q<�ZQ<A&P<hN<��L<�K< nJ<�  �  �3F<�qG<��I<M�L<��O<��Q<4�R<^R<)�P<}LN<�QK<CUH<��E<%>D<��C<��D<tTF<��H<5L<I�N< >Q<G�R<-�R<�oQ<yO<�!L<�>I<$G<�(F<��F<-SH<��J<�M<�tP<R<aR<�SQ<gO<�EL<SoI<JBG<>9F<��F<�9H<y�J<��M<|�P<y_R<s�R<eR<�,P<~yM<pqJ<t�G<�XE<mD<�D<�,E<�PG<O&J<[3M<:�O<PR<r�R<f�R<J�P<!ZN<�TK< �H<�F<�ZF<Q@G<1SI<ML<�O<�OQ<<�R<�YR<��P<�^N<pK<e�H<A�F<�KF<G<�I<W�K<�N<xbQ<��R<��R<*�Q<�eO<%�L<I<�F<��D<mD<nWD<T�E<�;H<20K<-1N<S�P<^tR<��R<,R<�(P<.UM<�UJ<��G<�F<�zF< �G<X/J<CM<u�O<^�Q<l�R<��Q<�P<�iM<}J<	H<h�F<�kF<��G<vJ<��L<)�O<��Q<��R<��R<��P<z~N<�K<��H</	F<JpD<[�C<}�D<A�F<(I<*.L<�O<�gQ<=�R<��R<�Q<�<O<IEL<�aI<Y=G<ELF<��F<�wH<5K<nN<��P<�9R<��R<{Q<}FO<�kL<��I<fG<<[F<��F<ZWH<��J<��M<��P<�rR<��R<�$R<V7P<�M<�uJ<�G<+WE<�D<+D<�!E<�BG<}J<�M<~�O<��Q<�R<9zR<y�P<�5N<�-K<wH<,�F</.F<G<�#I<��K<��N<�Q<,QR<;)R<��P<�/N<�AK<A�H<�F<1 F<J�F<=�H<��K<6�N<�6Q<�R<�R<pQ<'5O<2VL<�KI<��F<R�D<h�C<� D<��E<�H<��J<��M<)�P<E>R<��R<��Q<��O<QM<�J<��G<hDF<�=F<�G<��I<��L<��O<-�Q<`ZR<
�Q<C�O<�+M<E@J<��G<UF<�  �  �(B<�bC<�F<��I<n	M<C�O<tEQ<N*Q<��O<��L<glI<�E<�C<�/A<ɣ@<�~A<2�C<�F<�5J<��M<ZP<�VQ<�Q<QO<�PL<��H<�`E<BC<p)B<��B<\E<�H<.�L<��O<�R<�}R<$Q<=N<F�J<R�F<
�C<�\B<�{B<�:D<Z;G<��J<�1N<�P<ÈQ<��P<�N<Q�K<WcH<�E<�sB<RA<��@<P?B<�D<�
H<��K<ӪN<U�P<y�Q<V�P<Y�N<�[K<��G<��D<)�B<�tB<��C<�F<JJ<E	N<|Q<��R<�eR<�tP<E7M<�gI<@�E<�WC<�SB<��B<
5E<{H<�L<�1O<�"Q<�Q<pP<GN<,�J<�GG<D D<��A<��@<�CA<0�B<��E<!=I<�L<��O<�CQ<s�Q<~AP<�M<B J<řF<��C<qB<R�B<�D<��G<ÍK<�$O<�Q<��R<"�Q<�}O<E�K<*H<��D<��B<�`B<�C<<;F<�I<�;M<+P<wQ<�[Q<�O<�M<<�I<(F<�?C<LaA<��@<�A<o�C<�F<gbJ<w�M<u6P<(~Q<�>Q<�uO<�tL<��H<��E<S(C<�LB<�!C<�E<��H<��L<	 P<9=R<��R<�BQ<_dN<ٯJ<��F<D<:B<�B<�XD<�VG<��J<�GN<��P<X�Q<��P<��N<��K<�gH<YE<>rB<��@<�@<�4B<�D<��G<�yK<	�N<��P<��Q<�P<k�N<7K<�G<nD<�B<	HB<�C<IpF<bJ<�M<�P<PiR<�4R<`DP<�M<�9I<
�E<�+C<L(B<��B<�
E<�PH<[�K<vO<l�P<�aQ<oAP<6�M<��J<�G<Z�C<�A<f�@<�A<��B<��E<�I<�vL<�OO<�Q<EUQ<�
P<�cM<1�I<�`F<*�C<&5B< xB<:[D<�G<�LK<]�N<.zQ<
{R<�Q<�=O<u�K<��G<�D< �B<�  �  �b?<�@<�eC<�.G<�K<0JN<�P<?)P<�N<��K<�H<�KD<#(A<�"?<�><4x?<I�A<�E<��H<�kL<BO<�NP<��O<�M<�KJ<7SF<�B< 8@<xj?< z@<<?C<�9G<��K<�{O<��Q<�kR<d�P<SxM<�2I<��D<3�A<ڲ?<��?<'zA<��D<H�H<�gL<N.O<�kP<@�O<��M<m�J<��F<�LC<�}@<��><��><�D@<8�B<+�F<�NJ<ğM<��O<��P<{�O<9�L<�4I<�?E<�A<��?<�?<oA<�D<E�H<�5M<��P<?�R<HR<*P< DL<��G<%�C<��@<�?<�1@<��B<jF<JJ<'�M<��O<'�P<�uO<��L<Y{I<H�E<FLB<��?<s�><�3?<�A<D<�G<.�K<��N<EP<�`P<5�N<i�K<�G<y D<vA<��?<$@<�VB<��E<�XJ<Y~N<ӀQ<խR<��Q<��N<�J<0sF<��B<)A@<�?<I�@<��C<bG<*NK<|N<EP<�ZP<X�N<��K<09H<?}D<�YA<,T?<�><+�?<+�A<$GE<�I<�L<;O<�uP<��O<}�M<�oJ<GvF<��B<[@<�?<4�@<"dC<^_G<+�K<�O<gR<��R<\�P<ܟM<YYI<GE<[�A<>�?<��?<B�A<S�D<X�H<�}L<�AO<w|P<��O<_�M<�J<G�F<xNC<n|@<��><��>< :@<b�B<MuF<�:J<�M<��O<oP<&bO<9�L<I<�E<��A<��?<�?<b@A<7}D<{�H<2M<�}P<�TR<R<��O<�L<I�G<�C<��@<�m?<@@<�WB<I�E<��I<"_M<٫O<UP<QGO<+�L<2JI<ԀE<�B<+�?<0�><�><��@<��C<�G<9LK<�NN<&P<�*P<��N<#�K<�G< �C<��@<dl?<��?<�B<^�E<�J<<N<�>Q<�kR<>zQ<9�N<�J<�5F<�qB<?@<�  �  ��<؝<pn<3%<\�,<��3<�8<�N;<��;< �9<�j6<î2<�T/<�-<Vo,<�w-<� 0<��3<[77<�7:<��;<��:<�7<�+2<+<ɝ#<21<��<��<��<��<Q�%<_@-<ı3<�7<��8<�5<$X0<M")<ܾ!<�<'E<�<
<u� <��'<�;/<��5<��9<7�;<�9;<g�8<�S5<�1<�.<.�,<��,<nW.<�G1<]�4<��8<R;<��;<\:<@Q6<2$0<��(<�!<�<zg<�B<,_<,,!<�|(<�/<��5<I�8<�.8<�w4<�9.<.�&<��<O\<*�<�<��<��"<Z`*<��1<*^7<y�:<��;<��:<��7<�4<��0<��-<u�,<N&-<:/<x|2<w86<=�9<s�;<��;<D9<�o4<��-<�<&<�S<�?<��<j�<K<9}#<��*<(�1<��6<l�8<�I7<�2<��+<�J$<��<}7<��<��<��<�f%<��,<^�3<?�8<�;<�;<��9<��6<�2<'�/<�J-<�,<��-<00<��3<�c7< b:<�;<�;<��7<�O2<�1+<�#<8S<S<��<�<'�<�%<nh-<��3<�7<�8<�6<��0<�K)<[�!<��<9j<�0<}*<9� <��'<�S/<��5<� :<��;<3E;<��8<�X5<��1<s�.<x�,<��,<:L.<B91<��4<�s8<];<��;<>:<006<B 0<8�(<�[!<:�<v9<�<�-<=� <�H(<��/<�\5<-`8<j�7<�E4<�.<��&<�y<�/<��<�<!�<\�"<�6*<Ln1<�27<�:<۲;<3v:<(�7<��3<�Y0<c�-<Zv,<��,<Q/<�E2<�6<�W9<.d;<�q;<�9<�84<؁-<�&<�<�<�<Ū<��<9:#<��*<�1<M�6<�8<>7<�Z2<�+<$<f<�<�  �  nV<K<1  <Ò&<��-<!j4<�D9<��;<��;<:<n�6<;M3<N
0<&�-<�:-<�;.<P�0<�4<�7<Y�:<�<<Ot;<<e8< 3<1=,<�	%<9�<��<�a<uP<E <��&<,.<TO4<48<B�8<f6<<1<�*<f�"<B+<I�<��<�<�$"<�)<+D0<c6<e�:<�9<<��;<
N9<��5<]H2<6S/<��-<��-<�/<��1<�5<49<��;<�Z<<E�:<'7<�$1<#	*<�#<Y<�<��<�<�m"<W~)<��0<\6<�9<��8<5<�	/<Z�'<�� <��<�<Q�<f\< m$<�+<�2<�8<�f;<:S<<�;<6J8<��4<a<1<�.<�w-<�-<�/<�3<u�6<T:<:
<<�!<<��9<�C5<3�.<̕'<�� <�<�<$�<�n<��$<��+<l�2<vk7<�B9< �7<�F3<��,<Vp%<< �<w�<��<E5 <S�&<+.<՛4<-v9<-�;<$<<DN:<�$7<�3<�<0<c.<ll-<dl.<��0<J4<��7<��:<�E<<�;<R�8<�93<�_,<,%<N�<��<��<�t<�D <g '<0?.<tx4<^8<�9<��6<�>1<}F*<�!#<$R<J<��<k�<dB"<�1)<"\0<	x6<;�:<vH<<�;<QV9<��5<)J2<�Q/<��-<ƅ-<�
/<X�1<Et5<f�8<�t;<�?<<2�:<�6<� 1<w�)<Z�"<b-<��<�<}�<�:"<�J)<LZ0<��5<��8<Yp8<��4<��.<٤'<�� <d�<�l<V<�2<�C$<yl+<�_2<K�7<�9;<�$<<��:<�8<��4<�1<zo.<�A-<R�-<*�/<��2<��6<��9<��;<>�;<�9<5<��.<]'<�� <8�<ed<�A<t-<�f$<��+<z\2<'&7<��8<��7<�3<�q,<�0%<��<؎<�  �  �<8�<{X$<JS*<��0<�6<��:<��<<��<<�<;<qL8<N�4<��1<Y
0<�v/</]0<��2<c�5<9<��;<�+=<��<<E:<4}5<k/<V�(<S=#<�]<�<$�<�#<p�)<e0<+�5<�j9<L:<��7<d3<z�,<$m&<�F!<at<�|<L!<�O&<:�,<�3<\c8<��;<dV=<�<<s~:<^U7<
4<�\1<G�/<��/<&1</�3<17<�;:<�<<�r=<+K<</�8<��3<4w-<L'<�!<)�<�}<g!<.�%<�I,<~�2<)�7<):<�9<��6<0C1<��*<�$<�* <A<]<<%�"<ue(<��.<�5<��9<�<<�d=<�,<<��9<�B6<=3<��0<O�/<�0<��1<�4<�$8<�*;<+=<DJ=<.i;<l7<��1< B+<�*%<ݔ <#]<��<0h"<�'<�s.<]{4<��8<h`:<�9</5<D*/<��(<��"<@;<�G<�1 <r�$<̆*<O1<��6<;<q,=<U0=<�n;<�~8<'5<�02<�<0<٨/<�0<�2<�5<�19<��;<�T=<��<<�B:<8�5<	�/<�)<�_#<-�<4<[�<h$<*<��0<!6<��9<�>:<�7<v=3<��,<V�&<�m!</�<"�<Dl!<wm&<�,<�3<4x8<{ <<e=<��<<��:<aZ7<�4<t[1<��/<��/<�1<Ŭ3<��6<�&:<��<<�W=<(-<<:�8<�3<�P-<"�&<t�!<]�<�M<� <��%<V,<ll2< d7<+�9<�9<pt6<X1<_�*<x$<�<�<	<g�"<�;(<��.<4�4<L�9<�<<�5=<��;<�\9<N6<t�2<ċ0<�|/<��/<x�1<�4<��7<�:<��<<�=<�2;<*57<�1<�	+<��$<EY <�<��<J'"<��'<�/.<�64<�y8<�:<��8<Q�4<��.<�f(<��"<= <�  �  O�$<��&<�|*<({/<��4<Jj9<�<<�+><��=<�h<<��9<27<2�4<0&3<��2<�g3<E/5<T�7<f�:<��<<�-><S�=<<<�8</�3<W.<8�)<2&<�$<H&<1])<�=.<Ǝ3<�8< �:<,z;<��9<+�5<��0<�k+<fK'<�&%<�c%<��'<v(,<�^1<�6<<�:<3z=<[k><��=<s�;<z9<�e6<�;4<w3<f�2<%4<'6<A�8<��;<A�=<��><�=<�G;<!67<U2<V�,<4t(<�%<�;%<� '<1+<�;0<�k5<	{9<œ;<�M;<0�8<�L4<� /<�*<�t&<�%<&<v?)<�-<83<�,8<�;<�
><j><�A=<��:<�<8<�5<-�3<��2<hA3<K�4<�	7<#�9<i`<<$><�p><|=<�:<ӎ5<I0<v6+< J'<�C%<��%<D8(<ڰ,<��1<h�6<�k:<��;<v�:<Sh7<M�2<�A-<�(<��%<�+%<!�&<��*<��/<�4<!�9<��<<a]><�0><�<<o:<uR7<��4<}Y3<��2<�3<`5<��7<��:<�	=<TW><'><x=<<h�8<��3<�y.<��)<�T&<i%<�+&<��)<Hd.<v�3<�E8<�;<�;<��9<��5<��0<��+<�q'<"K%<&�%<�(<�E,<@y1<��6<��:<؋=<�y><��=<��;<q#9<�g6<:4<�3<p�2<�4<�6<��8<�};<j�=<f><�=<';<u7<��1<_�,<�H(<Z�%<V%<��&<��*<L0<�75<4G9<=`;<�;<R�8<�4<��.<�)<bH&<\�$<��%<�)<5�-<�3<8<��;<�=<�:><=<6�:<�8<�n5<��3<[�2<�	3<�{4<G�6<ӗ9<t)<<��=<:><�<<��9<nW5<�0<��*<�'<�%<�S%<��'<o,<��1<��6<j':<�|;<$k:< &7<�T2<�-<�e(<�%<�  �  ��,<�A.<o1<��4<Ӄ8<��;<�=<�><�'><N�<<-;<#9<�7<$�6<YG6<e�6<�7<�9<�~;<7<=<�T><�o><pX=<H
;<��7<{�3<�n0<j�-< �,<?F-<̈́/<Z�2<��6<�:<'*<<E�<<84;<p^8<ܫ4<��0<S.<e�,<�+-<�./<kc2<�'6<	�9<��<<�6><5�><��=<�t<<+�:<��8<)M7<��6<V�6<�37<��8<a:<�P<<!�=<M�><�j><`�<<,>:<�6<��2<X�/<[|-<\�,<M.<��0<�n4<O-8<�$;<p�<<5{<<x�:<W[7<ڊ3<�0<5�-<��,<��-<=0<\�3<�|7<�:<�O=<Q�><e�><H�=<��;<a�9<@:8<�7<܁6<��6<'�7<�'9<�;<��<<�C><n�><
><D<<a9<�i5<U�1<f�.<�-<g-<k�.<��1<ӱ5<�E9<�;<��<<Y<<3�9<�6<�L2<�/<�)-<��,<�w.<�S1<��4<?�8<��;<��=<��><Z><O=<�B;<W9<(�7<J�6<{6<U�6<�8<3�9<��;<�h=<4><<�>< =<k/;<��7<�4<ɑ0<c�-<x�,<�j-<�/<�3<.�6<?:<AS<<ɹ<<�];<��8<^�4<C1<:C.<{�,<�M-<EN/<x�2<CB6<��9<w�<<KH><��><�=<�|<<�:<E�8<�K7<2�6<a|6<�(7<P8<�O:<�;<<_�=<�><.M><��<<�:<��6<@�2<Gz/<&O-<D�,<��-<ޓ0<�;4<�7<C�:<Q|<<�H<<�`:<�*7<�[3<��/<�n-<p�,<-�-<�0<!�3<R7<��:<-#=<^><zc><�c=</�;<u�9<8<;�6<�I6<5}6<�f7<[�8<��:<��<<�><ڂ><��=<��;<7�8<�15<&~1<ʁ.<y�,<��,<�.<��1<�o5<%9<�;<ی<<��;<�\9<��5<�2<��.<��,<�  �  �4<�&5<G�6<��8<��:<tP<<�=<a0=<��<<b<<�$;<|]:<}�9<�9<f�9<�9<��9<��:<@W;<�5<<Y�<< :=<��<<�<<�:<�8<Y�6<��4< 4<�4<n/5<W7<�D9<�B;<�<<*�<<��;<9:<�8<P�5<�}4<��3<kn4<��5<��7<��9<��;<0�<<eM=<�:=<ͮ<<P�;<�;<�O:<��9<�9<T�9<��9<�G:<{�:<;�;<�<<�E=<ck=<��<<5�;<:<�8<96<�4<.!4<��4<��5<t�7<�.:<o�;<$�<<��<<*�;<#�9<�w7<e�5<�S4<�4<>�4<_v6<�x8<�|:<�<<N=<�g=<�&=<�}<<�;<C�:<D1:<K�9<G�9<t�9<n:<6�:<XD;<�"<<��<<%`=<�R=<@�<<K;<:i9<lX7<�5<N_4<s4<�4<ތ6<��8<��:<hf<<=<�<<;<��8<Q�6<	5<:'4<3J4<R\5<�7<�,9<�;<��<<�D=<�b=<��<<8<<Y;<O�:<�
:<�9<,�9<	�9<� :<�:<Ά;</c<<�=<�c=<"=<�9<<��:<ů8<��6<�5<�$4<&<4<�T5<57<�k9<�j;<��<<0�<<�<<�a:<�48<,6<,�4<�4<��4<��5<l�7<��9<*�;<��<<�^=<!I=<��<<T�;<�;<:Q:<k�9<L�9<_�9<��9<f9:<�:<��;<m�<<&+=<�M=<\�<<�;<�9<d�7<�5<�4<��3<M_4<1�5<%�7<��9<��;<~�<<Ԝ<<o;<9<�H7<�X5<'4<�3<g�4<�K6<�M8<~Q:<��;<��<<�8=<3�<<�J<<�n;<_�:<�9<�9<j�9<K�9<M�9<aJ:< ;<:�;<��<<g)=<V=<�l<<;<�19<�7<O5<�#4<s�3<��4<�L6<�t8<��:<R$<<��<<�C<<��:<��8<�6<��4<��3<�  �  L�9<�D:<s�:<�;<@;<��:<�=:<��9<7d9<�`9<g�9<�U:<�
;<��;<��;<;<��:<�/:<��9<
[9<Hs9<��9<�a:<��:<,;<�;<Ը:<>0:<Ʊ9<i9<�u9<6�9<Ӂ:<55;<�;<��;<�y;<{�:<�$:<��9<�j9<�9<��9<��:<�;<TD;<5$;<��:<�.:<�9<�{9<T�9<:<ֹ:<Gj;<��;<��;<�;<t�:<�):<�9<'�9<��9<>8:<��:<7:;<&g;<�7;<B�:<y8:<��9<
�9<��9<8B:<��:<�;<l�;<�;<�t;<t�:<G:<��9<��9<E�9<wH:<f�:<�;;<$X;<�;<h�:<�:<
�9<-�9<��9<�R:<4;<��;<��;<��;<�V;<Т:<��9<��9<�9<��9<]c:<��:<�J;< X;<�;<�:<�:<ݤ9<}�9<��9<�s:<=);<��;<�<<��;<r<;<r�:<��9<Q�9<y�9<2�9<�y:<j�:<�Q;<�N;<��:<Tp:<p�9<ė9<�9<��9<t�:<�@;<��;<��;<G�;<�;<Cb:<Z�9<��9<ϟ9<�:<,�:<@
;<UQ;<�>;<��:<�S:<��9<h�9<��9<(:<��:<�\;<6�;<,�;<{�;<��:<\L:<�9<��9<�9<!:<h�:<+%;<^;<+;;<��:<�?:< �9<��9<?�9<�:<p�:<�h;<�;<�;<�t;<+�:<2:<i�9<�t9<<�9<�:<F�:<-;<�A;<�;<�:<:<��9<Nh9<��9<p:<��:<�g;<E�;<m�;<�C;<��:<��9<y9<Nb9<��9<i:<��:<�;<^,;<��:<*o:<��9<Qy9<�W9<X�9<�:<��:<ap;< �;<��;<�;<Ei:<��9<je9<�^9<��9<�,:<3�:<�;<� ;<��:<�Q:<0�9<�h9<�U9<��9<�3:<��:<߀;<��;<��;<.�:<�H:<L�9<�[9<�d9<�  �  �0=<=<�?<<��:<��8<��6<45<�4<��3<�4<U�6<��8<��:<�U<<��<<�<<�}:<�Z8<�66<��4<�3<664<[m5<'E7<�W9<;5;<x�<<L,=<�1=<��<<��;<�;<�O:<O�9<&�9<B�9<B�9<�:<~�:<9�;<�i<<t=<<M=<�<<��;<�M:<�G8<J6<s�4<�4<1L4<��5<Ӄ7<��9<��;<��<<G�<<�;<��9<��7<��5<�u4<54<��4<w26<=+8<O8:<��;<�=<[t=<yI=<��<<J�;<a�:<�P:<e�9<|�9<��9<��9<oj:<� ;<��;<��<<�Q=<c\=<��<<�;<R�9<��7<@�5<}4<�4<߭4<U56<R8<�}:<�.<<��<<_�<<�U;<fQ9<�7<[E5<�:4<�24<� 5<'�6<��8<�:<�S<<�2=<uk=<�=<�_<<��;<��:<�!:<>�9<f�9<)�9<�:<��:<di;<�G<<[=<7g=<�?=<�s<<� ;<�9<L 7<�E5<?4<�)4<5<<�6<>9<�;<�<<��<<�N<<ǲ:<F�8<�h6<I�4<�4<�a4<��5<�l7<�}9<Z;<��<<P=<�U=<�<<�<<~3;<Gv:<��9<��9<=�9<2�9<7::<P�:<��;<M�<<4=<�m=<u=<�<<g:<�^8<�]6<g�4<�4<W4<T�5<��7<�9<�;<�<<S�<<��;<��9<A�7<U�5<G^4<��3<l�4<Y6<n8<�:<��;<��<<YH=<�=<�}<<ߤ;< �:<�:<��9<Ր9<Δ9<��9<;:<��:<��;<��<<�%=< 1=<J�<<�_;<��9<}7<;�5<IL4<N�3<Oy4<��5<8<JD:<��;<˾<<fo<<!;<#9<V�6<�5<4<��3<Q�4<�6<��8<^�:<b<<i�<<�1=<��<<n#<<�D;<�u:<J�9<y�9<�|9<�9<Z�9<�c:<�-;<�<<`�<<�  �  �z><��=<:z;<Q8<�4<��0<^#.<3�,<-<��.<F2<>6<ʋ9<��;<!�<<{;<��8<�>5<�x1<Bm.<��,<
�,<��.<$�1<Aq5<�9<l<<��=<N�><><��<<y�:<��8<3d7<�6<�\6<��6<M+8<��9<��;<�=<>< j><=<?�:<.47<�k3<" 0<��-<c�,<T�-<Q0<B�3<�{7<أ:<v<<�<<��:<,�7<�&4<χ0<�-<��,<s�-<��/<� 3<��6<�l:< =<�}><��><B�=<|C<<T:<��8<y67<��6<��6<Yo7<��8<6�:<��<<�><S�><>:><��<<��9<�6<dH2<�"/<7-<�,<�^.<#K1<N	5<ܶ8<�|;<��<<:C<<�:<�6<��2<6�/<�]-<Y�,<�.<��0<yY4<�8<�`;</�=<��><t~><�[=<ٙ;<d�9<��7<#�6<��6<��6<W�7<�u9<lb;<e/=<~h><y�><�=<��;<��8<��4<#1<LV.<��,<�6-<J4/<�|2<�N6<��9<!<<5�<<|�;<9<�s5<��1<�.<�,<T-<��.<R�1<Η5<(E9<�:<<�><`�><i/><q�<<�:<�
9<�7<]�6<+�6<E7<TR8<<:<3<<�=<+�><6�><<=<�:<PM7<!�3<�0<��-<6�,<!�-<&0<�3<}7<3�:<Jq<<(�<<��:<��7<�4<ss0<��-<��,<Gk-<��/<��2<��6< E:<v�<<R><E�><t�=<�<<T#:<dU8<7<�`6<Dt6<\?7<ү8<�:<�r<<l�=<��><�><<W<<�|9<	�5<@2<6�.<y-<��,<0).<�1<Z�4<�|8<|A;<5�<<g<<&�9< �6<կ2<N/<�%-<�,<M�-<ӑ0<k#4<��7<�);<Lh=<|n><&D><^ =<];<�l9<v�7<r�6<�A6<n�6<�7<�99<�';<p�<<)1><�  �   ><��<<�/9<�~4<�//<�=*<��&<��$<��%<\�(<�O-<Ϣ2<�d7<)�:<J~;<�:<7r6<tv1<-,<��'<&F%<%<dC'<�G+<�e0<��5<�:<�=<�K><��=<3<<�}9<�6<o4<�3<��2<α3<g�5<�B8<Q;<�==<U><�=<í;<��7<��2<�-<$�(<��%<�%<�&<�/*<�9/<�4<��8<QM;<Eq;<,99<25<��/<��*<��&<'%<M�%<u�(<J-<�c2<�y7<1z;<U�=<i�><��=<W{;<x�8<�6<�
4<�3<�#3<�f4<P�6<LX9<j�;<��=<�{><ur=<H�:<�^6<)1<��+<[�'<�m%<hU%<�'<w�+<G1<R,6<��9<ڮ;<";<�8<Ur3<.<pM)<J&<�%<K�&<�)<|�.<�4<��8<�m<<&>><�V><t�<<��:<N�7<H5<�3<��2<Rn3<55<y}7<lE:<_�<<#@><cU><׶<<�b9<��4<*b/<ep*<�&<� %<��%<��(<�-<
�2<��7<P�:<I�;<E@:<}�6<3�1<�`,<p�'<�u%<'I%<9n'<�p+<�0<]�5<h>:<#5=<�o><� ><;<< �9<��6<��4<�33<��2<��3<��5<�h8<*;<aa=<�v><��=<z�;<��7<|�2<R�-<�)<��%<T%<Ò&<�7*<i>/<��4<��8<�H;<Ri;<.9<5<q�/<r�*<��&<�%<A�%<��(<��,<�>2<�R7<�P;<�=<iZ><k=<�K;< �8<��5<��3<��2<��2<O74<xm6<Y*9<U�;<��=<�O><�F=<�:<W26<��0<B�+< �'<{;%<"!%<�f'<O�+<z�0<5�5<ȹ9<Vr;<��:<��7<�63<��-<�)<��%<��$<�I&<�)<��.<��3<R�8<i6<<�><B><��<<W:<{�7<�
5<YQ3<׫2<13<��4<AB7<�:<�<<]	><�  �  ��<<�:<?\6<�w0<��)<�$<0�<N
<�%<M�"<S�(<�G/<5<n�8<�:<HR8<��3<��-<_'<��!<��<N4<K� <HH%<<o+<��1<j�7<g;<3*=<�<<��:<��7<Ow4<?�1<F�/<&�/<�0<�3<uQ6<_�9<�,<<MN=<F�<<�9<�4<�j.<D�'<��"<d
<�7<�H <y�$<�+<M�1<@�6<�9<�:<�K7<p92<��+<}�%<D� <�b<��<�!"<�m'<0�-<R!4<@>9<�o<<�{=<g�<<�:<��6<��3<�1<��/<�/<�1<JH4<��7<�:<��<<�b=<^�;<�58<\�2<T,<�&<�.!<t�<n�<��!<��&<�X-<3<�/8<_K:<�x9<!�5<�80<�)<��#<c�<�;<�<��#<�u)<��/<I�5<q:<��<<U=<��;<�9<q�5<��2<0<h�/<�U0<\Z2<2Z5<�8<��;<�?=<�=<��:<2�6<��0<5**<�@$<� <�><�Z<�/#< �(<��/<�Q5<A09<GV:<`�8<�'4<^.<��'<
"<�<�a<�� <�q%<��+<�2<�7<��;<{N=<o�<<o ;< �7<�4<��1<�0<�/<��0<%D3<�v6<Ͽ9<�O<<�o=<۟<<��9<C�4<;�.<\(<��"<�< E<WS <�$<9+<��1<��6<=�9<��9<�@7<G+2<p�+<=~%<� <�H<�<�"<�K'<q�-<E�3<9<�D<<�N=<G_<<��9<�6<o3<#�0<M�/<��/<�^1<�4<.i7<�:<��<<7=<��;<�	8<��2<g&,<o�%<�� <�S<�u<�n!<ѯ&<M-<�Q3<�7<>:<v;9<g�5<��/<'{)<�#<�q<<vy<�y#<@@)<�/<#�5<�H:<��<<=<��;<��8<N|5<�h2<
B0<jp/<<0<�2<�5<�w8<�\;<?	=<�  �  p�;<J9<�4< j-<|-&<��<^<�S<?�<^<˘%<�,<X3<`�7<E�8<��6<
2<B+<�	$<�<�&<�w<��<�!<��'<�/<ig5<��9<�<<�;<ȳ9<�e6<��2<2�/<9�-<�W-<��.<�F1<�4<�Z8<b;<�;<<40;<O�7<�2<�+<;�#<<kM<�<J<�<!<�((<�V/<XA5<��8<��8<��5<�0<1)<� "<�<��<�(<%�<`[#<�n*<�1<TZ7<�;<�e<<�|;<��8<_5<��1<"/<��-<��-<��/<Ҋ2<s(6<��9<$�;<�C<<�i:<�+6<��/<��(<��!<��<��<q<��<h#<6�*<M�1<��6<�+9<�=8<514<��-<�&<��<L<׉<��<�C<r�%<"�,<p�3<m�8<��;<
G<<<�:<�7<+4<��0<oZ.<�p-<W,.<;j0<&�3<�Z7<v:<�2<<1�;<�@9<�G4<��-<�_&<r�<�O<Y�<��<EQ<��%<4-<��3<��7<j89<h27<�D2<y+<�>$<�<'W<ʥ<Z<C/!<��'<�-/<��5<D
:<.)<<m�;<|�9<��6<w�2<R�/<��-<!~-<�.<�l1<Z�4< 8<E<;<6]<<�O;<��7<�52< 5+<:$<�<�]<��<�<TD!<\-(<!X/<�?5<ץ8<�8<��5<y0<��(<c�!<�u<��<�<�t<.9#<�I*<+]1<L17<��:<9<<�N;<�8<>/5<D�1<��.<Rd-<��-<CX/<M\2<��5<�]9<դ;<�<<�=:<��5<��/<��(<D�!<�^<��<<�<b[<6F#<Yr*< \1<��6<]�8<i 8<'�3<��-<�d&<��<\<KR<3�<�<�b%<��,<�e3<̘8<��;<d<<v�:<�7<u�3<3�0<�.<04-<<�-<�.0<�|3<�!7<�>:<��;<�  �  8;<�h8<�53<�F,<��$<�<in<ɧ<�)<�<�v$<��+<�2<�57<K�8<u6<qY1<UR*<��"<~~<�<��<$C<�z<Aw&<��-<��4<�K9<j�;<J_;<�;9<��5<H 2<,�.<�,<��,<Y�-<��0<�34<u�7<3�:<n�;<5�:<�7<�%1<&�)<�"<d<�<j�<H�<$�<@'<)�.<��4<78<�j8<�:5<�W/<��'<�� <0<�!<7x<|�<h�!<�-)<8�0<��6<~�:<�;<;<gf8<2�4<&1<�F.<�,<�,<A�.<��1<��5<�9<Ta;<N�;<��9<b5<��.<�w'<�] <��<<$�<Q!<tH"<Q�)<��0<�B6<�8<H�7<�3<�-<�%<֞<)�<��<�I<{�<G/$<��+<��2<�$8<�<;<�;<�H:<�97<r�3<v0<�-<1�,<sf-<ϵ/<�3<A�6<T:<��;<�l;</�8<�h3<Iy,<��$<�M<ޡ<E�<i_<�<�$<3,<��2<p7<��8<Ǯ6<�1<o�*<�#<x�<��<�<�n<��<�&<&.<�4<]p9<ư;<��;<�`9<��5<�E2<?/<t-<�,<�.<��0<�X4<��7<�:<��;<��:<&"7<�@1<��)<�"<]w<��<��<ڎ<��<� '<��.<
�4<K28<�b8<�/5<�I/<��'<�� <�<�<X[<��<=�!<?	)<S`0<�t6<�]:<��;<2�:<p78<q�4<��0<T.<ә,<��,<�.<'�1<m5<��8<5;<c�;<Ĩ9<�55<�.<�I'<s. <��<��<�L<��<"<P{)<1�0<�6<G�8<��7<�S3<N�,<�I%<�d<g�<��<<�u<��#<p+<!2<]�7<g;<��;<8:<8�6<�G3<G�/<xY-<�h,<|*-<�z/<��2<s�6<��9<��;<�  �  p�;<J9<�4< j-<|-&<��<^<�S<?�<^<˘%<�,<X3<`�7<E�8<��6<
2<B+<�	$<�<�&<�w<��<�!<��'<�/<ig5<��9<�<<�;<ȳ9<�e6<��2<2�/<9�-<�W-<��.<�F1<�4<�Z8<b;<�;<<40;<O�7<�2<�+<;�#<<kM<�<J<�<!<�((<�V/<XA5<��8<��8<��5<�0<1)<� "<�<��<�(<%�<`[#<�n*<�1<TZ7<�;<�e<<�|;<��8<_5<��1<"/<��-<��-<��/<Ҋ2<s(6<��9<$�;<�C<<�i:<�+6<��/<��(<��!<��<��<q<��<h#<6�*<M�1<��6<�+9<�=8<514<��-<�&<��<L<׉<��<�C<r�%<"�,<p�3<m�8<��;<
G<<<�:<�7<+4<��0<oZ.<�p-<W,.<;j0<&�3<�Z7<v:<�2<<1�;<�@9<�G4<��-<�_&<r�<�O<Y�<��<EQ<��%<4-<��3<��7<j89<h27<�D2<y+<�>$<�<'W<ʥ<Z<C/!<��'<�-/<��5<D
:<.)<<m�;<|�9<��6<w�2<R�/<��-<!~-<�.<�l1<Z�4< 8<E<;<6]<<�O;<��7<�52< 5+<:$<�<�]<��<�<TD!<\-(<!X/<�?5<ץ8<�8<��5<y0<��(<c�!<�u<��<�<�t<.9#<�I*<+]1<L17<��:<9<<�N;<�8<>/5<D�1<��.<Rd-<��-<CX/<M\2<��5<�]9<դ;<�<<�=:<��5<��/<��(<D�!<�^<��<<�<b[<6F#<Yr*< \1<��6<]�8<i 8<'�3<��-<�d&<��<\<KR<3�<�<�b%<��,<�e3<̘8<��;<d<<v�:<�7<u�3<3�0<�.<04-<<�-<�.0<�|3<�!7<�>:<��;<�  �  ��<<�:<?\6<�w0<��)<�$<0�<N
<�%<M�"<S�(<�G/<5<n�8<�:<HR8<��3<��-<_'<��!<��<N4<K� <HH%<<o+<��1<j�7<g;<3*=<�<<��:<��7<Ow4<?�1<F�/<&�/<�0<�3<uQ6<_�9<�,<<MN=<F�<<�9<�4<�j.<D�'<��"<d
<�7<�H <y�$<�+<M�1<@�6<�9<�:<�K7<p92<��+<}�%<D� <�b<��<�!"<�m'<0�-<R!4<@>9<�o<<�{=<g�<<�:<��6<��3<�1<��/<�/<�1<JH4<��7<�:<��<<�b=<^�;<�58<\�2<T,<�&<�.!<t�<n�<��!<��&<�X-<3<�/8<_K:<�x9<!�5<�80<�)<��#<c�<�;<�<��#<�u)<��/<I�5<q:<��<<U=<��;<�9<q�5<��2<0<h�/<�U0<\Z2<2Z5<�8<��;<�?=<�=<��:<2�6<��0<5**<�@$<� <�><�Z<�/#< �(<��/<�Q5<A09<GV:<`�8<�'4<^.<��'<
"<�<�a<�� <�q%<��+<�2<�7<��;<{N=<o�<<o ;< �7<�4<��1<�0<�/<��0<%D3<�v6<Ͽ9<�O<<�o=<۟<<��9<C�4<;�.<\(<��"<�< E<WS <�$<9+<��1<��6<=�9<��9<�@7<G+2<p�+<=~%<� <�H<�<�"<�K'<q�-<E�3<9<�D<<�N=<G_<<��9<�6<o3<#�0<M�/<��/<�^1<�4<.i7<�:<��<<7=<��;<�	8<��2<g&,<o�%<�� <�S<�u<�n!<ѯ&<M-<�Q3<�7<>:<v;9<g�5<��/<'{)<�#<�q<<vy<�y#<@@)<�/<#�5<�H:<��<<=<��;<��8<N|5<�h2<
B0<jp/<<0<�2<�5<�w8<�\;<?	=<�  �   ><��<<�/9<�~4<�//<�=*<��&<��$<��%<\�(<�O-<Ϣ2<�d7<)�:<J~;<�:<7r6<tv1<-,<��'<&F%<%<dC'<�G+<�e0<��5<�:<�=<�K><��=<3<<�}9<�6<o4<�3<��2<α3<g�5<�B8<Q;<�==<U><�=<í;<��7<��2<�-<$�(<��%<�%<�&<�/*<�9/<�4<��8<QM;<Eq;<,99<25<��/<��*<��&<'%<M�%<u�(<J-<�c2<�y7<1z;<U�=<i�><��=<W{;<x�8<�6<�
4<�3<�#3<�f4<P�6<LX9<j�;<��=<�{><ur=<H�:<�^6<)1<��+<[�'<�m%<hU%<�'<w�+<G1<R,6<��9<ڮ;<";<�8<Ur3<.<pM)<J&<�%<K�&<�)<|�.<�4<��8<�m<<&>><�V><t�<<��:<N�7<H5<�3<��2<Rn3<55<y}7<lE:<_�<<#@><cU><׶<<�b9<��4<*b/<ep*<�&<� %<��%<��(<�-<
�2<��7<P�:<I�;<E@:<}�6<3�1<�`,<p�'<�u%<'I%<9n'<�p+<�0<]�5<h>:<#5=<�o><� ><;<< �9<��6<��4<�33<��2<��3<��5<�h8<*;<aa=<�v><��=<z�;<��7<|�2<R�-<�)<��%<T%<Ò&<�7*<i>/<��4<��8<�H;<Ri;<.9<5<q�/<r�*<��&<�%<A�%<��(<��,<�>2<�R7<�P;<�=<iZ><k=<�K;< �8<��5<��3<��2<��2<O74<xm6<Y*9<U�;<��=<�O><�F=<�:<W26<��0<B�+< �'<{;%<"!%<�f'<O�+<z�0<5�5<ȹ9<Vr;<��:<��7<�63<��-<�)<��%<��$<�I&<�)<��.<��3<R�8<i6<<�><B><��<<W:<{�7<�
5<YQ3<׫2<13<��4<AB7<�:<�<<]	><�  �  �z><��=<:z;<Q8<�4<��0<^#.<3�,<-<��.<F2<>6<ʋ9<��;<!�<<{;<��8<�>5<�x1<Bm.<��,<
�,<��.<$�1<Aq5<�9<l<<��=<N�><><��<<y�:<��8<3d7<�6<�\6<��6<M+8<��9<��;<�=<>< j><=<?�:<.47<�k3<" 0<��-<c�,<T�-<Q0<B�3<�{7<أ:<v<<�<<��:<,�7<�&4<χ0<�-<��,<s�-<��/<� 3<��6<�l:< =<�}><��><B�=<|C<<T:<��8<y67<��6<��6<Yo7<��8<6�:<��<<�><S�><>:><��<<��9<�6<dH2<�"/<7-<�,<�^.<#K1<N	5<ܶ8<�|;<��<<:C<<�:<�6<��2<6�/<�]-<Y�,<�.<��0<yY4<�8<�`;</�=<��><t~><�[=<ٙ;<d�9<��7<#�6<��6<��6<W�7<�u9<lb;<e/=<~h><y�><�=<��;<��8<��4<#1<LV.<��,<�6-<J4/<�|2<�N6<��9<!<<5�<<|�;<9<�s5<��1<�.<�,<T-<��.<R�1<Η5<(E9<�:<<�><`�><i/><q�<<�:<�
9<�7<]�6<+�6<E7<TR8<<:<3<<�=<+�><6�><<=<�:<PM7<!�3<�0<��-<6�,<!�-<&0<�3<}7<3�:<Jq<<(�<<��:<��7<�4<ss0<��-<��,<Gk-<��/<��2<��6< E:<v�<<R><E�><t�=<�<<T#:<dU8<7<�`6<Dt6<\?7<ү8<�:<�r<<l�=<��><�><<W<<�|9<	�5<@2<6�.<y-<��,<0).<�1<Z�4<�|8<|A;<5�<<g<<&�9< �6<կ2<N/<�%-<�,<M�-<ӑ0<k#4<��7<�);<Lh=<|n><&D><^ =<];<�l9<v�7<r�6<�A6<n�6<�7<�99<�';<p�<<)1><�  �  �0=<=<�?<<��:<��8<��6<45<�4<��3<�4<U�6<��8<��:<�U<<��<<�<<�}:<�Z8<�66<��4<�3<664<[m5<'E7<�W9<;5;<x�<<L,=<�1=<��<<��;<�;<�O:<O�9<&�9<B�9<B�9<�:<~�:<9�;<�i<<t=<<M=<�<<��;<�M:<�G8<J6<s�4<�4<1L4<��5<Ӄ7<��9<��;<��<<G�<<�;<��9<��7<��5<�u4<54<��4<w26<=+8<O8:<��;<�=<[t=<yI=<��<<J�;<a�:<�P:<e�9<|�9<��9<��9<oj:<� ;<��;<��<<�Q=<c\=<��<<�;<R�9<��7<@�5<}4<�4<߭4<U56<R8<�}:<�.<<��<<_�<<�U;<fQ9<�7<[E5<�:4<�24<� 5<'�6<��8<�:<�S<<�2=<uk=<�=<�_<<��;<��:<�!:<>�9<f�9<)�9<�:<��:<di;<�G<<[=<7g=<�?=<�s<<� ;<�9<L 7<�E5<?4<�)4<5<<�6<>9<�;<�<<��<<�N<<ǲ:<F�8<�h6<I�4<�4<�a4<��5<�l7<�}9<Z;<��<<P=<�U=<�<<�<<~3;<Gv:<��9<��9<=�9<2�9<7::<P�:<��;<M�<<4=<�m=<u=<�<<g:<�^8<�]6<g�4<�4<W4<T�5<��7<�9<�;<�<<S�<<��;<��9<A�7<U�5<G^4<��3<l�4<Y6<n8<�:<��;<��<<YH=<�=<�}<<ߤ;< �:<�:<��9<Ր9<Δ9<��9<;:<��:<��;<��<<�%=< 1=<J�<<�_;<��9<}7<;�5<IL4<N�3<Oy4<��5<8<JD:<��;<˾<<fo<<!;<#9<V�6<�5<4<��3<Q�4<�6<��8<^�:<b<<i�<<�1=<��<<n#<<�D;<�u:<J�9<y�9<�|9<�9<Z�9<�c:<�-;<�<<`�<<�  �  L�9<�D:<s�:<�;<@;<��:<�=:<��9<7d9<�`9<g�9<�U:<�
;<��;<��;<;<��:<�/:<��9<
[9<Hs9<��9<�a:<��:<,;<�;<Ը:<>0:<Ʊ9<i9<�u9<6�9<Ӂ:<55;<�;<��;<�y;<{�:<�$:<��9<�j9<�9<��9<��:<�;<TD;<5$;<��:<�.:<�9<�{9<T�9<:<ֹ:<Gj;<��;<��;<�;<t�:<�):<�9<'�9<��9<>8:<��:<7:;<&g;<�7;<B�:<y8:<��9<
�9<��9<8B:<��:<�;<l�;<�;<�t;<t�:<G:<��9<��9<E�9<wH:<f�:<�;;<$X;<�;<h�:<�:<
�9<-�9<��9<�R:<4;<��;<��;<��;<�V;<Т:<��9<��9<�9<��9<]c:<��:<�J;< X;<�;<�:<�:<ݤ9<}�9<��9<�s:<=);<��;<�<<��;<r<;<r�:<��9<Q�9<y�9<2�9<�y:<j�:<�Q;<�N;<��:<Tp:<p�9<ė9<�9<��9<t�:<�@;<��;<��;<G�;<�;<Cb:<Z�9<��9<ϟ9<�:<,�:<@
;<UQ;<�>;<��:<�S:<��9<h�9<��9<(:<��:<�\;<6�;<,�;<{�;<��:<\L:<�9<��9<�9<!:<h�:<+%;<^;<+;;<��:<�?:< �9<��9<?�9<�:<p�:<�h;<�;<�;<�t;<+�:<2:<i�9<�t9<<�9<�:<F�:<-;<�A;<�;<�:<:<��9<Nh9<��9<p:<��:<�g;<E�;<m�;<�C;<��:<��9<y9<Nb9<��9<i:<��:<�;<^,;<��:<*o:<��9<Qy9<�W9<X�9<�:<��:<ap;< �;<��;<�;<Ei:<��9<je9<�^9<��9<�,:<3�:<�;<� ;<��:<�Q:<0�9<�h9<�U9<��9<�3:<��:<߀;<��;<��;<.�:<�H:<L�9<�[9<�d9<�  �  �4<�&5<G�6<��8<��:<tP<<�=<a0=<��<<b<<�$;<|]:<}�9<�9<f�9<�9<��9<��:<@W;<�5<<Y�<< :=<��<<�<<�:<�8<Y�6<��4< 4<�4<n/5<W7<�D9<�B;<�<<*�<<��;<9:<�8<P�5<�}4<��3<kn4<��5<��7<��9<��;<0�<<eM=<�:=<ͮ<<P�;<�;<�O:<��9<�9<T�9<��9<�G:<{�:<;�;<�<<�E=<ck=<��<<5�;<:<�8<96<�4<.!4<��4<��5<t�7<�.:<o�;<$�<<��<<*�;<#�9<�w7<e�5<�S4<�4<>�4<_v6<�x8<�|:<�<<N=<�g=<�&=<�}<<�;<C�:<D1:<K�9<G�9<t�9<n:<6�:<XD;<�"<<��<<%`=<�R=<@�<<K;<:i9<lX7<�5<N_4<s4<�4<ތ6<��8<��:<hf<<=<�<<;<��8<Q�6<	5<:'4<3J4<R\5<�7<�,9<�;<��<<�D=<�b=<��<<8<<Y;<O�:<�
:<�9<,�9<	�9<� :<�:<Ά;</c<<�=<�c=<"=<�9<<��:<ů8<��6<�5<�$4<&<4<�T5<57<�k9<�j;<��<<0�<<�<<�a:<�48<,6<,�4<�4<��4<��5<l�7<��9<*�;<��<<�^=<!I=<��<<T�;<�;<:Q:<k�9<L�9<_�9<��9<f9:<�:<��;<m�<<&+=<�M=<\�<<�;<�9<d�7<�5<�4<��3<M_4<1�5<%�7<��9<��;<~�<<Ԝ<<o;<9<�H7<�X5<'4<�3<g�4<�K6<�M8<~Q:<��;<��<<�8=<3�<<�J<<�n;<_�:<�9<�9<j�9<K�9<M�9<aJ:< ;<:�;<��<<g)=<V=<�l<<;<�19<�7<O5<�#4<s�3<��4<�L6<�t8<��:<R$<<��<<�C<<��:<��8<�6<��4<��3<�  �  ��,<�A.<o1<��4<Ӄ8<��;<�=<�><�'><N�<<-;<#9<�7<$�6<YG6<e�6<�7<�9<�~;<7<=<�T><�o><pX=<H
;<��7<{�3<�n0<j�-< �,<?F-<̈́/<Z�2<��6<�:<'*<<E�<<84;<p^8<ܫ4<��0<S.<e�,<�+-<�./<kc2<�'6<	�9<��<<�6><5�><��=<�t<<+�:<��8<)M7<��6<V�6<�37<��8<a:<�P<<!�=<M�><�j><`�<<,>:<�6<��2<X�/<[|-<\�,<M.<��0<�n4<O-8<�$;<p�<<5{<<x�:<W[7<ڊ3<�0<5�-<��,<��-<=0<\�3<�|7<�:<�O=<Q�><e�><H�=<��;<a�9<@:8<�7<܁6<��6<'�7<�'9<�;<��<<�C><n�><
><D<<a9<�i5<U�1<f�.<�-<g-<k�.<��1<ӱ5<�E9<�;<��<<Y<<3�9<�6<�L2<�/<�)-<��,<�w.<�S1<��4<?�8<��;<��=<��><Z><O=<�B;<W9<(�7<J�6<{6<U�6<�8<3�9<��;<�h=<4><<�>< =<k/;<��7<�4<ɑ0<c�-<x�,<�j-<�/<�3<.�6<?:<AS<<ɹ<<�];<��8<^�4<C1<:C.<{�,<�M-<EN/<x�2<CB6<��9<w�<<KH><��><�=<�|<<�:<E�8<�K7<2�6<a|6<�(7<P8<�O:<�;<<_�=<�><.M><��<<�:<��6<@�2<Gz/<&O-<D�,<��-<ޓ0<�;4<�7<C�:<Q|<<�H<<�`:<�*7<�[3<��/<�n-<p�,<-�-<�0<!�3<R7<��:<-#=<^><zc><�c=</�;<u�9<8<;�6<�I6<5}6<�f7<[�8<��:<��<<�><ڂ><��=<��;<7�8<�15<&~1<ʁ.<y�,<��,<�.<��1<�o5<%9<�;<ی<<��;<�\9<��5<�2<��.<��,<�  �  O�$<��&<�|*<({/<��4<Jj9<�<<�+><��=<�h<<��9<27<2�4<0&3<��2<�g3<E/5<T�7<f�:<��<<�-><S�=<<<�8</�3<W.<8�)<2&<�$<H&<1])<�=.<Ǝ3<�8< �:<,z;<��9<+�5<��0<�k+<fK'<�&%<�c%<��'<v(,<�^1<�6<<�:<3z=<[k><��=<s�;<z9<�e6<�;4<w3<f�2<%4<'6<A�8<��;<A�=<��><�=<�G;<!67<U2<V�,<4t(<�%<�;%<� '<1+<�;0<�k5<	{9<œ;<�M;<0�8<�L4<� /<�*<�t&<�%<&<v?)<�-<83<�,8<�;<�
><j><�A=<��:<�<8<�5<-�3<��2<hA3<K�4<�	7<#�9<i`<<$><�p><|=<�:<ӎ5<I0<v6+< J'<�C%<��%<D8(<ڰ,<��1<h�6<�k:<��;<v�:<Sh7<M�2<�A-<�(<��%<�+%<!�&<��*<��/<�4<!�9<��<<a]><�0><�<<o:<uR7<��4<}Y3<��2<�3<`5<��7<��:<�	=<TW><'><x=<<h�8<��3<�y.<��)<�T&<i%<�+&<��)<Hd.<v�3<�E8<�;<�;<��9<��5<��0<��+<�q'<"K%<&�%<�(<�E,<@y1<��6<��:<؋=<�y><��=<��;<q#9<�g6<:4<�3<p�2<�4<�6<��8<�};<j�=<f><�=<';<u7<��1<_�,<�H(<Z�%<V%<��&<��*<L0<�75<4G9<=`;<�;<R�8<�4<��.<�)<bH&<\�$<��%<�)<5�-<�3<8<��;<�=<�:><=<6�:<�8<�n5<��3<[�2<�	3<�{4<G�6<ӗ9<t)<<��=<:><�<<��9<nW5<�0<��*<�'<�%<�S%<��'<o,<��1<��6<j':<�|;<$k:< &7<�T2<�-<�e(<�%<�  �  �<8�<{X$<JS*<��0<�6<��:<��<<��<<�<;<qL8<N�4<��1<Y
0<�v/</]0<��2<c�5<9<��;<�+=<��<<E:<4}5<k/<V�(<S=#<�]<�<$�<�#<p�)<e0<+�5<�j9<L:<��7<d3<z�,<$m&<�F!<at<�|<L!<�O&<:�,<�3<\c8<��;<dV=<�<<s~:<^U7<
4<�\1<G�/<��/<&1</�3<17<�;:<�<<�r=<+K<</�8<��3<4w-<L'<�!<)�<�}<g!<.�%<�I,<~�2<)�7<):<�9<��6<0C1<��*<�$<�* <A<]<<%�"<ue(<��.<�5<��9<�<<�d=<�,<<��9<�B6<=3<��0<O�/<�0<��1<�4<�$8<�*;<+=<DJ=<.i;<l7<��1< B+<�*%<ݔ <#]<��<0h"<�'<�s.<]{4<��8<h`:<�9</5<D*/<��(<��"<@;<�G<�1 <r�$<̆*<O1<��6<;<q,=<U0=<�n;<�~8<'5<�02<�<0<٨/<�0<�2<�5<�19<��;<�T=<��<<�B:<8�5<	�/<�)<�_#<-�<4<[�<h$<*<��0<!6<��9<�>:<�7<v=3<��,<V�&<�m!</�<"�<Dl!<wm&<�,<�3<4x8<{ <<e=<��<<��:<aZ7<�4<t[1<��/<��/<�1<Ŭ3<��6<�&:<��<<�W=<(-<<:�8<�3<�P-<"�&<t�!<]�<�M<� <��%<V,<ll2< d7<+�9<�9<pt6<X1<_�*<x$<�<�<	<g�"<�;(<��.<4�4<L�9<�<<�5=<��;<�\9<N6<t�2<ċ0<�|/<��/<x�1<�4<��7<�:<��<<�=<�2;<*57<�1<�	+<��$<EY <�<��<J'"<��'<�/.<�64<�y8<�:<��8<Q�4<��.<�f(<��"<= <�  �  nV<K<1  <Ò&<��-<!j4<�D9<��;<��;<:<n�6<;M3<N
0<&�-<�:-<�;.<P�0<�4<�7<Y�:<�<<Ot;<<e8< 3<1=,<�	%<9�<��<�a<uP<E <��&<,.<TO4<48<B�8<f6<<1<�*<f�"<B+<I�<��<�<�$"<�)<+D0<c6<e�:<�9<<��;<
N9<��5<]H2<6S/<��-<��-<�/<��1<�5<49<��;<�Z<<E�:<'7<�$1<#	*<�#<Y<�<��<�<�m"<W~)<��0<\6<�9<��8<5<�	/<Z�'<�� <��<�<Q�<f\< m$<�+<�2<�8<�f;<:S<<�;<6J8<��4<a<1<�.<�w-<�-<�/<�3<u�6<T:<:
<<�!<<��9<�C5<3�.<̕'<�� <�<�<$�<�n<��$<��+<l�2<vk7<�B9< �7<�F3<��,<Vp%<< �<w�<��<E5 <S�&<+.<՛4<-v9<-�;<$<<DN:<�$7<�3<�<0<c.<ll-<dl.<��0<J4<��7<��:<�E<<�;<R�8<�93<�_,<,%<N�<��<��<�t<�D <g '<0?.<tx4<^8<�9<��6<�>1<}F*<�!#<$R<J<��<k�<dB"<�1)<"\0<	x6<;�:<vH<<�;<QV9<��5<)J2<�Q/<��-<ƅ-<�
/<X�1<Et5<f�8<�t;<�?<<2�:<�6<� 1<w�)<Z�"<b-<��<�<}�<�:"<�J)<LZ0<��5<��8<Yp8<��4<��.<٤'<�� <d�<�l<V<�2<�C$<yl+<�_2<K�7<�9;<�$<<��:<�8<��4<�1<zo.<�A-<R�-<*�/<��2<��6<��9<��;<>�;<�9<5<��.<]'<�� <8�<ed<�A<t-<�f$<��+<z\2<'&7<��8<��7<�3<�q,<�0%<��<؎<�  �  >?�;ا;,��;���;w��;�A<lM<��<��<��<�<!E<�c<�N<�<�<�<��<܍<-�<6_<�< <)u <p��;c��;TB�;:��;Vu�;���;��;��;b��;�<<�<=\	<]�<�;k�;d��;�ѯ;�y�;4_�;բ�;�A�;��;1X�;0a<c<m�<t�<�w<�X<�l<��<m<m�<D�<�!<�<T^<q�<�e<�c<^�<��;6*�;�1�;H��;=V�;�(�;�Y�;Y��;���;���;�E<�W	<گ<�l<%��;�;Sq�;BӪ;��;lʤ;yt�;u�;��;�U�;
 <��<�0<@�<�<8t<��<�<�<�^<�Q<v&<w�<	�<`a<�<��<��<`y�;��;�|�;���;B�;��;�6�;9��;���;�J�;��<j�	<�0<���;�\�;���;b�;��;k��;G�;��;w�;�a�;�r<b~<�'<#<��<8@<	x<��<�<��<��<b-<s<h�<��<G�<Ǽ<D<�� <'�;;�;��;Eť;���;�F�;���;�%�;���;�g<h;<��	<	<m�;���;�A�;�%�;�ɣ;s��;��;ԁ�;�;���;�w<7v<4�<԰<��<2^<�n<;�<�<5�<�t<�<\<�H<J�<iI<�C<v�<
O�;*��;���;(c�;B��;�¢;�;�?�;|��;���;9<� 	<�y<U8<�:�;���;�;�y�;���;Rw�;6#�;�$�;���;��;��
<��<�<��<X�<�@<�K<��<�<h'<�<��<3�<%�<�*<��<�S<��<P	�;��;3�;;�;Dd�;`�;ʮ�;.0�;I��;���;vE<h	<��<�;��;� �;��;O<�;�  �  �#�;\��;���;6�;y��;��<�,<��<�S<I�<l<��<c <a<lk<n]<V�<�a<��<�<��<7<<��<��;���;��;�\�;cQ�;�y�;�y�;3��;h��;�<T1	<�w
<D< �;��;�a�;��;T6�;_G�;	P�;�V�;�;���;1�<6%<�O<��<;�<�<��<b<z�<˽<+<Z�<�<�<�,<��<�<��	<μ�;I�;�0�;�`�;�<�;��;͢�;M:�;���;��;?�<�t
<��	<f�<���;���;,�;�>�;�ާ;���;b��;IG�;��;� <� <�<Ǟ<�?<�O<
�<"<��<*�<�<
�<��<j_<�<��<DU<�_<�<���;E}�;���;wx�;!ʧ;9A�;OF�;�;��;��;�</�
<cY<� <!��; ��;(]�;GN�;�;B�;Fe�;���;���;��<�]<ø<t�<J.<��<��<�3<�:<'�<@�<��<��<�<*=<+�<]<29<�<���;��;��;#��;���;
®;�ſ;�(�;p�;'�<�]	<�
<�G<�Z�;�k�;��;k\�;*��;v��;̕�;���;�I�;���;��<W8<�_<<+�<��<��<�`<��<��<a<O�<�m<�<�<�<%�<�	<�p�;!��;L��;��;ۨ;戨;)9�;���;rA�; ��;�I<�=
<�	<�<�a�;���;���;K�;���;cW�; ��;���;ܴ�;�v <�<�y<�p<�<�<e�<��<m�<�q<��<2�<m<(<��<�<�<%)<��<���;�
�;�C�;=��;iK�;潪;���;]y�;t�;ӄ�;�q<_�
<f<�` <�7�;�2�;޺;�ԫ;�  �  ���;ν;���;���;:�;��<wa<��<�)<�<I<�<��<@�<�m<�9<�<m�<��<��<c�<��<��<�<��;��;���;��;�·;��;��;�4�;���;w+<�H<�u<q	<i<)e�;�;���;�W�;/θ;��;^�;p��;�� <��<�<o<[�<u�<t�<�K<i<s�<L�<��<�<3�<r<��<��<L�<��<�<���;q��;��;���;�(�;���;D�;IC�;�. <-�<�v<��<@<���;b�;v��;���;WA�;#�;�G�;���;t��;��<�<x:<]�<��<�<P�<�<��<�<�	<%�<�<�D<��<L�<w�<�v<�X	<�F�;՞�; 9�;P��;�R�;&�;���;�&�;��;p<��
<*�<��<�s<�Q�;��;bs�;��;h�;�<�;��;�	�;?��;F*<��<�<R[<<�<	|<�)<l�<�$<�<%l<�I<��<��<��<#�<�<&�<߸<�?�;e��;��;w��;=�;7�;Af�;��;�.�;]V<u<��<V�	<�F<��;�]�;�;릹;��;,`�;���;���;,� <��< <�~<��<Y�<�<�M<	<��<�<�<� <�n<P\<��<B�<��<ԑ<��<�0�;��;E��;:[�;ø;i%�;h��;���;��;��<4@<�<�<�<�;E��;Q2�;;/�;R�;���;���;y9�;�O�;W<.�<�<�e<��<7�<+�<>X<b<+s<��<�`<��<H<Ț<�W<�_<�?<�!	<4��;�,�;q��;��;�Է;���;��;%��;XE�;-(<��
<�<=><�-<���;x�;#��;���;�  �  ,��;z	�;$��;��;*<�4<��<��<��<!�<d�<K<h�<n< <t�<��<�<(H<]<+*< <mH<EI
<�� <۹�;�N�;�B�;��;:��;�5�;���;�<�L<Յ<?�<�<L�<�}�;���;,u�;I��;w��;��;��;BS�;�L<G<'�<N0<Q<��<�<B�<hN<�_<ST<i/<�<�u<��<�-<M�<��<�<3x<���;�D�;�Z�;���;���;n��;*$�;���;;<ީ<^�<<f?<U7<�_�;VP�;��;,�;���;��;��;���;�p	<��<z�<?<:<}�<v<*Y<u�< M<S�<��<|P<�<�$<>�<��<��<QZ<�I<�J�;J��;ݍ�;�Y�;�t�;Ԭ�;'�;� <��<�h<��<c�<��	<�<I�;G:�;92�;�$�;Hw�;���;�,�;F5<tf<�<M<ĺ<�.<�+<2<��<��<@E<��<�'<N�<Tv<F7<�S<a'<�m<�l
<N<#��;��;���;��;���;s��;�4�;�,<2w<��<ĳ<rD<�'<���;P�;���;�B�;Z�;���;�O�;H��;(f<s(<�<�?<�<��<N�<E�<M<&[<L<�#<�<pc<��<�<}<Dx<�<�R<�p�;���;���;�>�;�~�;�; ��;�S�;2<s<Y<��<�<<&��;e��;0��;���;�o�;s��;��;"��;�F	<|<P{<$�<�<]j<��<�"<˽<�<}W<�r<�<��<�<:�<QR<s<o#<F<c��;�7�;m�;���;���;�'�;:}�;���;��<D!<t�<ڞ<��	<r� <<��;I��;��;�  �  �;I��;E �;�/<[ 	<t<n�<ZI<�3<��<Ӄ<y�<Z4<��<�<E�<�W<w<؟<e�<�<��<�<�<7�<8� <4��;��;��;$��;�f�;l�<�]
<��<��<ʣ<��<ap<_M<>!�;�{�;4�;���;Q��;{�;��<Y<
|<�6<�:<��<��<�x<��<�-<��<��<N$<��<�r<&�<��<��<��<�4<�5<�r<X��;R��;$��;8�;���;�;G�<��<_�<ܴ<�N<��<,V<}�<w�;���;�|�;�`�;C��;�/ <��<Γ<�L<sw<��<t�<��<�O<��<�<_�<��<�\<=<i�<� <��<��<�d<uP<��	<l$<���;�)�;��;�9�;��;�� <� <`
<%<��<Wg<�<]�<�<�2�;x��;tv�;7]�;_i�;c<u2	<��<�<c{<�f<K�<4�<�<�i<)�<0�<�<ي<�8<,�<m�<�<��<@�<�B<;�<o� <*��;���;[�;��;��;�$<��
<��<�<��<�!<o�<�x<�u�;F��;�R�;�"�;$��;�M�;ק<<r<��<eI<�I<��<c�<�}<��<3,<��<��<�<ͱ<�`<��<��<mp<i�</<9<�J<*d�;��;53�;:��;$v�;��;iw<��<u<<�<]<I$<\�<˹�;���; &�;��;C��;= <�<�h<� <hI<t�<P�<ʩ<�<	i<'�<�<�<#<��<�s<��<=R<��<�-<�<��	<�<C:�;���;�"�;ú�;��;X� <#�<��<߿<��<�!<r<�<�N<P��;$S�;�  �  ҝ<}�<+�<�%	<4�<n<˵<\�<�<%<��<��<.�<a<+<<<jq< �<w�<��<��<xO<*0<�T<,�<�i<Q<�9<o�<3%<5v<�<�<<J<��<+�<5<�W<Zl	<�o<?"<]�<H<�<m
<��<<<;Q<W�<��<�o<�E<��<Y<C`<<Jd<w�<��<��<=�<"�<*�<Hu<h�
<��<��<�<z/<RG<$	<K�<��<��<��<ר<><,�<G�< <��<�<�;<Z,<�0<��<"<�<�H<�<�<�<��<5�<�-<Ft<�Y<'�<�*<�P<�h<�c<�<,<�<G<
�	<�q<��<��<	�<oZ<J�
<��<0[<q�<*<4	<��<�1<+<��<Z�<��<p�<^<uX	<J�<:3<��<��<�?<}J<�3<<��<;M<�r<�6<�<��<&�<�<��<�x<`W<z< <Ќ<�s<�\<��<I<ʛ<�<<D<ɨ<�t<! <�(<n`<<�<�	<��<cH<H�<�i<�#<ֈ
<�<�0<>�<w`<H�<��<�t<�G<@�<GT<X<��<`U<:�<#�<̦<>t<��<�e<P<d�
<�\<ƅ<�<�<8<��<�<F�<�<��<�t<>�<��<n�<��<\i<��<B<q<�<#�<k�<h�<�<�<��<��<<u\<��<�9<�<��<��<*<40<<,<��<n�<yU<<=�	<{8<�<-�<�`<<4`
<`<�<��<g�<%�<�<��<	�
<�<�<�  �  �W<X�<E�<�<z�<��<�<�c<T|<�[<��<��<W-<�<�m<��<ݪ<g
<1G<��<�.<�@<��<��<D�<��<��<�<��<E�<��<}b<*<��<Y%<r<�l<GT<u�<V�<{�<�<c<<��<��<&�<g�<��<2'<��<))<�H<'�<��<�<(f<{<�A<&<�M<��<0o<� <�L<�<�<N<�	<<h[<"<5�<$�<��<F?<�n<3�<<o<% <��<X�<~8<?"<_�<?3<� <��<��<�<�<�^<B;<Q�<�1<U�<��<O�<��<5C<R�<0<_g<L�<!�<�<�)<�<�<S�<��<%<�}<x<L8<�<�n<<
<K�</�<r<CK<�<��<8u<��<B�<�<�<��<��<��<i<�<f�<�< <��<He<R <��<��<��<�><Uy<N<�[<ak<<��<��<B�<��<�%<�<��<�<8�<R<��<lO<(�<m�<�~<g�</<��<2<�_<�<;<��<��<�<t9<��<�4<KQ<T�<f�<?<La<�r<H6<G�<�;<=�<�V<��<�-<��<��<��<|�<N�<s,<@�<�d<l�<mR<N
<�9<�b<�;<��<ur<̭<{
<��<�<�<��<�<��<�<��<o.<�<��<�<ʹ<|e<%r<�f<C<�j<�<<-<.�<�<�x<D�<g�<y�<�<h�<`�<B<�:<5�<+g<�,<?�<�<�j<��<�	<}<�<�9<He<�  �  )�<��<��< }<��<�<�p<I�<s�<�<�4<�:<�<*�<��<Eb<G�<�< "
<��<�N<g�<��<l<q�	<�K<A�<U <i�<�H<�J<v1<k
<5�<�2<�H<��<d<'�<7�<j�<#�<�<q�<��<�i<O�<��<8<��<��<�A<�<.<x3<�<y�<ڗ<��<"�<@�<f<�<�<�<�<.(<$�<�<1
<?�<+�<�<^�<�<D"<�u<�i<E�<�M<�u<�<��<�M<c�<�<1�<PO
<��<�B<��<�T<R�<�	<��<��<KQ<�	<�]<�v<J<��<�h<B/<��<�y<z�<��<�L<߰<I�<b�<�<�%<�<�<��<�C<z<�N<L�<T	<�+<�@<.2<��<��<C<}�<�&	<�<w�<��<8�<0�<l<Gs<?<�!<N<��<�<�S<�U
<�<x}<[�<�<\�< �	<�o<׭<�C<<m<�o<�W<2<��<\<�r<�(<�<^�<Y�<�<�<�7<��<w�<�<r<<?,<��<I�<�I<�	<�<�1<>�<D�<T�<ł<�<�<��<-�<�<Y�<{�<� <;}<ɇ<��<�}<L�<m�<{}<�L<��< B<�6<J�<E<�F<a<d<`"<sZ<��<�<P#
<k�<s<��<!<�<�	<�<�b<�<��<� <:<[�<��</<��<1�<�B<Cm<z�<E<Iy<kK<�`<��<�<B�<c�<v<<-8<X<.�<��<��<�<��<�  �  2 <
r<�<d�<��<f�;��;���;���;z[�;u�<�	<|�<S<ư<-�< q<ox<?$ <���;Z��;1J�;f,�;���;CU<(
<jv<u<��<�l<�<Ty<X�<�)<��<��<w�<,�<�5<$�<f�< �<N/<��<'%<�r<��;�7�;���;�n�;�7�;���;oQ<��<!�<oV<i�<T<3r<�0<�.�;E�;���;&��;g�;b�;�<�<��<��< �<6�<l�<�y<a�<�/<w�<��<>H<'�<��<��<��<�,<�<�?<�<>@<_��;h�;��;�w�;RI�;�.�;��<��<�]<��<z�<a�<�%
<��<H�;5��; g�;�P�;K��;�I<T<�<#<�<�2<�<��<a7<��<�<��<'�<x<e#<��<��<X<V<X�<Q<��<�<���;��;�f�;[�;7��;��<T	<�<܍<��<D�< �<��<6Y <�]�;���;j��;|��;N?�;�{<M
<�<ʘ<��<>�<C�<��<��<R<��<�<�<c�<K^<��<r�<h�<�Q<�<�B<��<*��;�a�;��;H��;�N�;/��;rV<=�<��<�Q<5�<�H<jc<�<)�;=�;���;x�;$�;^�; �<ej<�X<��<6�<�<��<SF<��<��<1�<K�<�<޷<�d<A�<r�<� <}�<�<�
<�<8�;��;i��;��;T��;���;��<8�<�<ş<L�<�k<��	<�<΢�;vW�;���;s��;83�;</�<�m<�<��<��<p�<��<�<�I<��<�<9�<"9<��<�<��<P <�  �  ޯ< d<޹<�y<���;��;���;Ч�;{)�;1��;̠�;we<4
<��<j�<��<xK<ŏ�;���;6s�;f��;��;M��;�+�;���;�<�<��<��<��<_�<��<<m<7]<U(<k�<�K<�<y�<�<��<{L<�*<K�<)��;$��;�0�;	G�;9%�;�q�;��;iJ�;|�<A�<{<z^<�><�<���;��;}��;���;���;���;�0�;���;��<<��<y�<8@<��< m<P�<�/<a<]z<�s<|<7�<�<z<<��<ʳ< �<bn�;�T�;�F�;$��;y�;�n�;���;���;Ş<p�<��<!�<�<�<�2�;���;���;��;��;�p�;@�;g�<�
<��<do<x<�><Ql<��<<M�<�J<��<��<6�<�D<�7<�<2�<ۗ<��<��<� �;��;g��;��;n��;O�;��;�<�B
<y<Q�<�<��<t �;	��;m��;&�;�i�;1�;�}�;�G�;u�<f�<��<�<W�<�<��<�3<F�<��</Q<Y<�t<�3<c�<@<h<?n<:J<Q�<���;K�;NZ�;Qj�;QB�;���;$�;JT�;(�<��<�<GV<}3<��<c�;y��;֖�;�c�;��;��;^��;t��;��<�S<0�<!�<f<��<D:</y<��<H.<JH<�B<��<|�<�<��<K�<[x<K�<�<��;���;���;�b�;��;���;U��;"k�;a<�R<��<F</�
<op<^��;;>�;N�;g��;d��;�;&��;�c<��
<��<�6<�=<?<K/<k�<�<ߎ<�<�u<�<�`<�	<��<�p<�  �  8�<y�<S`<P��;=_�;[��;�9�;:��;��;��;�V�;��;�<��<��<�a
<1�<��;�q�;�1�;6E�;+�;_ǿ;L��;ʈ�;�9�;־	<o�<��<x<b�<f�<#�<<S<5�<4�<�<�<��<�<I�<R<��<W<��<�,�;M6�;$D�;��;�D�;g�;ŀ�;�2�;���;��<�<A<Bn<��;���;h��;k��;Ѹ;���;���;��;���;��<6?<�D<>&<q�<9k<�n<�<��<L�<��<YI<�<��<q�<�<pI<3�<�<� <ew�;Hq�;D��;uθ;(�;���;o��;���;��<��	<��<�@<��<4�;�O�;�l�;_��;,�;ދ�;	 �;\D�;^��;[_<�1<P3<~<�<��<U�<2<`<@�<�;<�<^Q<t�<M�<�B<�<�<ؒ<OK�;:��;\�;���;�	�;n��;Ad�;��;3��;L�<i�<��<��
<6�<%��;��;��;���;�e�;��;�9�;���;Ӆ�;��	<��<��<��<r�<?"<��<�z<L�<��<��< �<u"<!7<c�<|u<�<�><S�<�`�;e�;!m�;��;qa�; +�;���;�<�;Ъ�;�<-�<�8<�b<O��;���;)��;�z�;t��;Y��;z��;���;���;��<�<�<>�<��<�9<P<<W�<ɴ<�<��<�<�P<�<{<��<�<��<��
<���;�;~�;K/�;�f�;���;�p�;T�;Ą�;
�<�	<�w<� <v�<
��;.��;���;�;�;Y��;��;���;���;�<�;�)<2�<W�<�<;�<��<�Y<��<�!<�g<��<�<�<eb< �<v<�  �  P5<��<��<��;���;�ݼ;5�;��;�n�;���;��;m��;�� <�^<Ζ
<!<�i�;)�;9.�;Ƿ;aO�;~�;;ɯ;���;���;h�;v�<�<nr<9�<��<�<wR<j�<��<Շ<v�<K<m�<�J<| <�V<�-<�z<���;�i�;���;�޶;w�;�;	�;n<�;Q;�;���;�<��	<�;
<_�<؈�;Y �;���;Ϧ�;z��;D�;c6�;>p�;9��;(+�;x
<��<<=A<p�<-h<��<&<�<��<��<,-<��<��<��<G"< �<D�<oL�;���;�K�;U��;F�;�ܩ;<C�;���;���;э�;��<ֻ
<�$	<�9<��;6��;/��;%�;���;�>�;:�;j�;��;M�<2�<?�<�!<D<G <�p<x�<}<��<�T<�\<�<��<�9<�h<�i<��<<�y�;|1�;�B�;ij�;ֈ�;Eܬ;�j�;S�;��;9+<��<,�
<�]<���;ޏ�;u��;1�;ͳ�;�ܧ;_"�;���;o��;�X�;��<v�<��<��<�
<�8<y<��<�<
�<��<7=<�<2q<TE<�y< O<��<���;��;	 �;��;O;�;��;���;�L�;E�;���;�<��	<�3
<��<qk�;���;Ϩ�;fv�;�T�;�B�;6��;�(�;_o�;v��;nM
<�_<K�<<y<6<#a<��<�<�<�b<��<K�<��<�<h�<V�<Y�<��;�l�;��;�R�;�ݧ;�n�;�е;p��;�R�;��;�i<^{
<��<D�<.Q�;OY�;�7�;���;�&�;zѫ;ح�;���;��;��<ȗ<��<�<�	<��<4<�g<A<e< <) <��<5�<�<S2<�  �  ��<��<Ў<�s�;D8�;���;�2�;�;�;cݦ;	�;q�;;B�;�)�;�7<�|	<g�<ݕ�;C��;g��;B��;���;��;�;�O�;�*�;;��;+T<��<��<MP<��<��<`�<4<k%<*�<	<ǅ<t|<q�<��<s�<w�<Vt
<���;�s�;���;[S�;C6�;��;�}�;���;[�;���;)�<��<@	<�<�;W�;�9�;�T�;���;���;{��;�{�;���;Z�;'f	<��<�<��<1T<O�<�<�r<<84<��<&�<Ɛ<��<E�<ӡ<J�<��<���;���;\,�;~�;m^�;�%�;P�;���;�1�;��;�v<�	<7<�� <��;���;�ҹ;]��;��;g�;ѭ�;��;W��;�X<��<�#<�<��<�<��<<y�<d�<�<��<A�<�e<��<c<,�<�<"�<O��;:��;��;��;쥡;�J�;-z�;���;���;���;Ju<4�	<f/<{�;^
�;I�;��;u�; ��;�d�;K��;�z�;���;Iy<@<�<�t<��<H�<��<l,<5M<I�<71<��<��<�<B�<�	<��<G�
<��;��;="�;|�;Y�;J5�;a��;Ҝ�;�d�;���;��<��<	<s�<�a�;43�;k�;u$�;R��;)]�;]Z�;24�;�]�;���;$;	<��<+y<��<�"<Q�<x�<O@<�<�<2�<�y<`b</n<�w<�u<��<��<v��;x%�;�̾;���;���;з�;t��;��;k��;�*�;�6<r`	<��<%� <��;�J�;\�;/�;H�;���;|B�;�Q�;8[�;*#<E�<u�<W�<��<�i<3�<��<��<��<�_<6�<:l<,<�<O�<�  �  P5<��<��<��;���;�ݼ;5�;��;�n�;���;��;m��;�� <�^<Ζ
<!<�i�;)�;9.�;Ƿ;aO�;~�;;ɯ;���;���;h�;v�<�<nr<9�<��<�<wR<j�<��<Շ<v�<K<m�<�J<| <�V<�-<�z<���;�i�;���;�޶;w�;�;	�;n<�;Q;�;���;�<��	<�;
<_�<؈�;Y �;���;Ϧ�;z��;D�;c6�;>p�;9��;(+�;x
<��<<=A<p�<-h<��<&<�<��<��<,-<��<��<��<G"< �<D�<oL�;���;�K�;U��;F�;�ܩ;<C�;���;���;э�;��<ֻ
<�$	<�9<��;6��;/��;%�;���;�>�;:�;j�;��;M�<2�<?�<�!<D<G <�p<x�<}<��<�T<�\<�<��<�9<�h<�i<��<<�y�;|1�;�B�;ij�;ֈ�;Eܬ;�j�;S�;��;9+<��<,�
<�]<���;ޏ�;u��;1�;ͳ�;�ܧ;_"�;���;o��;�X�;��<v�<��<��<�
<�8<y<��<�<
�<��<7=<�<2q<TE<�y< O<��<���;��;	 �;��;O;�;��;���;�L�;E�;���;�<��	<�3
<��<qk�;���;Ϩ�;fv�;�T�;�B�;6��;�(�;_o�;v��;nM
<�_<K�<<y<6<#a<��<�<�<�b<��<K�<��<�<h�<V�<Y�<��;�l�;��;�R�;�ݧ;�n�;�е;p��;�R�;��;�i<^{
<��<D�<.Q�;OY�;�7�;���;�&�;zѫ;ح�;���;��;��<ȗ<��<�<�	<��<4<�g<A<e< <) <��<5�<�<S2<�  �  8�<y�<S`<P��;=_�;[��;�9�;:��;��;��;�V�;��;�<��<��<�a
<1�<��;�q�;�1�;6E�;+�;_ǿ;L��;ʈ�;�9�;־	<o�<��<x<b�<f�<#�<<S<5�<4�<�<�<��<�<I�<R<��<W<��<�,�;M6�;$D�;��;�D�;g�;ŀ�;�2�;���;��<�<A<Bn<��;���;h��;k��;Ѹ;���;���;��;���;��<6?<�D<>&<q�<9k<�n<�<��<L�<��<YI<�<��<q�<�<pI<3�<�<� <ew�;Hq�;D��;uθ;(�;���;o��;���;��<��	<��<�@<��<4�;�O�;�l�;_��;,�;ދ�;	 �;\D�;^��;[_<�1<P3<~<�<��<U�<2<`<@�<�;<�<^Q<t�<M�<�B<�<�<ؒ<OK�;:��;\�;���;�	�;n��;Ad�;��;3��;L�<i�<��<��
<6�<%��;��;��;���;�e�;��;�9�;���;Ӆ�;��	<��<��<��<r�<?"<��<�z<L�<��<��< �<u"<!7<c�<|u<�<�><S�<�`�;e�;!m�;��;qa�; +�;���;�<�;Ъ�;�<-�<�8<�b<O��;���;)��;�z�;t��;Y��;z��;���;���;��<�<�<>�<��<�9<P<<W�<ɴ<�<��<�<�P<�<{<��<�<��<��
<���;�;~�;K/�;�f�;���;�p�;T�;Ą�;
�<�	<�w<� <v�<
��;.��;���;�;�;Y��;��;���;���;�<�;�)<2�<W�<�<;�<��<�Y<��<�!<�g<��<�<�<eb< �<v<�  �  ޯ< d<޹<�y<���;��;���;Ч�;{)�;1��;̠�;we<4
<��<j�<��<xK<ŏ�;���;6s�;f��;��;M��;�+�;���;�<�<��<��<��<_�<��<<m<7]<U(<k�<�K<�<y�<�<��<{L<�*<K�<)��;$��;�0�;	G�;9%�;�q�;��;iJ�;|�<A�<{<z^<�><�<���;��;}��;���;���;���;�0�;���;��<<��<y�<8@<��< m<P�<�/<a<]z<�s<|<7�<�<z<<��<ʳ< �<bn�;�T�;�F�;$��;y�;�n�;���;���;Ş<p�<��<!�<�<�<�2�;���;���;��;��;�p�;@�;g�<�
<��<do<x<�><Ql<��<<M�<�J<��<��<6�<�D<�7<�<2�<ۗ<��<��<� �;��;g��;��;n��;O�;��;�<�B
<y<Q�<�<��<t �;	��;m��;&�;�i�;1�;�}�;�G�;u�<f�<��<�<W�<�<��<�3<F�<��</Q<Y<�t<�3<c�<@<h<?n<:J<Q�<���;K�;NZ�;Qj�;QB�;���;$�;JT�;(�<��<�<GV<}3<��<c�;y��;֖�;�c�;��;��;^��;t��;��<�S<0�<!�<f<��<D:</y<��<H.<JH<�B<��<|�<�<��<K�<[x<K�<�<��;���;���;�b�;��;���;U��;"k�;a<�R<��<F</�
<op<^��;;>�;N�;g��;d��;�;&��;�c<��
<��<�6<�=<?<K/<k�<�<ߎ<�<�u<�<�`<�	<��<�p<�  �  2 <
r<�<d�<��<f�;��;���;���;z[�;u�<�	<|�<S<ư<-�< q<ox<?$ <���;Z��;1J�;f,�;���;CU<(
<jv<u<��<�l<�<Ty<X�<�)<��<��<w�<,�<�5<$�<f�< �<N/<��<'%<�r<��;�7�;���;�n�;�7�;���;oQ<��<!�<oV<i�<T<3r<�0<�.�;E�;���;&��;g�;b�;�<�<��<��< �<6�<l�<�y<a�<�/<w�<��<>H<'�<��<��<��<�,<�<�?<�<>@<_��;h�;��;�w�;RI�;�.�;��<��<�]<��<z�<a�<�%
<��<H�;5��; g�;�P�;K��;�I<T<�<#<�<�2<�<��<a7<��<�<��<'�<x<e#<��<��<X<V<X�<Q<��<�<���;��;�f�;[�;7��;��<T	<�<܍<��<D�< �<��<6Y <�]�;���;j��;|��;N?�;�{<M
<�<ʘ<��<>�<C�<��<��<R<��<�<�<c�<K^<��<r�<h�<�Q<�<�B<��<*��;�a�;��;H��;�N�;/��;rV<=�<��<�Q<5�<�H<jc<�<)�;=�;���;x�;$�;^�; �<ej<�X<��<6�<�<��<SF<��<��<1�<K�<�<޷<�d<A�<r�<� <}�<�<�
<�<8�;��;i��;��;T��;���;��<8�<�<ş<L�<�k<��	<�<΢�;vW�;���;s��;83�;</�<�m<�<��<��<p�<��<�<�I<��<�<9�<"9<��<�<��<P <�  �  )�<��<��< }<��<�<�p<I�<s�<�<�4<�:<�<*�<��<Eb<G�<�< "
<��<�N<g�<��<l<q�	<�K<A�<U <i�<�H<�J<v1<k
<5�<�2<�H<��<d<'�<7�<j�<#�<�<q�<��<�i<O�<��<8<��<��<�A<�<.<x3<�<y�<ڗ<��<"�<@�<f<�<�<�<�<.(<$�<�<1
<?�<+�<�<^�<�<D"<�u<�i<E�<�M<�u<�<��<�M<c�<�<1�<PO
<��<�B<��<�T<R�<�	<��<��<KQ<�	<�]<�v<J<��<�h<B/<��<�y<z�<��<�L<߰<I�<b�<�<�%<�<�<��<�C<z<�N<L�<T	<�+<�@<.2<��<��<C<}�<�&	<�<w�<��<8�<0�<l<Gs<?<�!<N<��<�<�S<�U
<�<x}<[�<�<\�< �	<�o<׭<�C<<m<�o<�W<2<��<\<�r<�(<�<^�<Y�<�<�<�7<��<w�<�<r<<?,<��<I�<�I<�	<�<�1<>�<D�<T�<ł<�<�<��<-�<�<Y�<{�<� <;}<ɇ<��<�}<L�<m�<{}<�L<��< B<�6<J�<E<�F<a<d<`"<sZ<��<�<P#
<k�<s<��<!<�<�	<�<�b<�<��<� <:<[�<��</<��<1�<�B<Cm<z�<E<Iy<kK<�`<��<�<B�<c�<v<<-8<X<.�<��<��<�<��<�  �  �W<X�<E�<�<z�<��<�<�c<T|<�[<��<��<W-<�<�m<��<ݪ<g
<1G<��<�.<�@<��<��<D�<��<��<�<��<E�<��<}b<*<��<Y%<r<�l<GT<u�<V�<{�<�<c<<��<��<&�<g�<��<2'<��<))<�H<'�<��<�<(f<{<�A<&<�M<��<0o<� <�L<�<�<N<�	<<h[<"<5�<$�<��<F?<�n<3�<<o<% <��<X�<~8<?"<_�<?3<� <��<��<�<�<�^<B;<Q�<�1<U�<��<O�<��<5C<R�<0<_g<L�<!�<�<�)<�<�<S�<��<%<�}<x<L8<�<�n<<
<K�</�<r<CK<�<��<8u<��<B�<�<�<��<��<��<i<�<f�<�< <��<He<R <��<��<��<�><Uy<N<�[<ak<<��<��<B�<��<�%<�<��<�<8�<R<��<lO<(�<m�<�~<g�</<��<2<�_<�<;<��<��<�<t9<��<�4<KQ<T�<f�<?<La<�r<H6<G�<�;<=�<�V<��<�-<��<��<��<|�<N�<s,<@�<�d<l�<mR<N
<�9<�b<�;<��<ur<̭<{
<��<�<�<��<�<��<�<��<o.<�<��<�<ʹ<|e<%r<�f<C<�j<�<<-<.�<�<�x<D�<g�<y�<�<h�<`�<B<�:<5�<+g<�,<?�<�<�j<��<�	<}<�<�9<He<�  �  ҝ<}�<+�<�%	<4�<n<˵<\�<�<%<��<��<.�<a<+<<<jq< �<w�<��<��<xO<*0<�T<,�<�i<Q<�9<o�<3%<5v<�<�<<J<��<+�<5<�W<Zl	<�o<?"<]�<H<�<m
<��<<<;Q<W�<��<�o<�E<��<Y<C`<<Jd<w�<��<��<=�<"�<*�<Hu<h�
<��<��<�<z/<RG<$	<K�<��<��<��<ר<><,�<G�< <��<�<�;<Z,<�0<��<"<�<�H<�<�<�<��<5�<�-<Ft<�Y<'�<�*<�P<�h<�c<�<,<�<G<
�	<�q<��<��<	�<oZ<J�
<��<0[<q�<*<4	<��<�1<+<��<Z�<��<p�<^<uX	<J�<:3<��<��<�?<}J<�3<<��<;M<�r<�6<�<��<&�<�<��<�x<`W<z< <Ќ<�s<�\<��<I<ʛ<�<<D<ɨ<�t<! <�(<n`<<�<�	<��<cH<H�<�i<�#<ֈ
<�<�0<>�<w`<H�<��<�t<�G<@�<GT<X<��<`U<:�<#�<̦<>t<��<�e<P<d�
<�\<ƅ<�<�<8<��<�<F�<�<��<�t<>�<��<n�<��<\i<��<B<q<�<#�<k�<h�<�<�<��<��<<u\<��<�9<�<��<��<*<40<<,<��<n�<yU<<=�	<{8<�<-�<�`<<4`
<`<�<��<g�<%�<�<��<	�
<�<�<�  �  �;I��;E �;�/<[ 	<t<n�<ZI<�3<��<Ӄ<y�<Z4<��<�<E�<�W<w<؟<e�<�<��<�<�<7�<8� <4��;��;��;$��;�f�;l�<�]
<��<��<ʣ<��<ap<_M<>!�;�{�;4�;���;Q��;{�;��<Y<
|<�6<�:<��<��<�x<��<�-<��<��<N$<��<�r<&�<��<��<��<�4<�5<�r<X��;R��;$��;8�;���;�;G�<��<_�<ܴ<�N<��<,V<}�<w�;���;�|�;�`�;C��;�/ <��<Γ<�L<sw<��<t�<��<�O<��<�<_�<��<�\<=<i�<� <��<��<�d<uP<��	<l$<���;�)�;��;�9�;��;�� <� <`
<%<��<Wg<�<]�<�<�2�;x��;tv�;7]�;_i�;c<u2	<��<�<c{<�f<K�<4�<�<�i<)�<0�<�<ي<�8<,�<m�<�<��<@�<�B<;�<o� <*��;���;[�;��;��;�$<��
<��<�<��<�!<o�<�x<�u�;F��;�R�;�"�;$��;�M�;ק<<r<��<eI<�I<��<c�<�}<��<3,<��<��<�<ͱ<�`<��<��<mp<i�</<9<�J<*d�;��;53�;:��;$v�;��;iw<��<u<<�<]<I$<\�<˹�;���; &�;��;C��;= <�<�h<� <hI<t�<P�<ʩ<�<	i<'�<�<�<#<��<�s<��<=R<��<�-<�<��	<�<C:�;���;�"�;ú�;��;X� <#�<��<߿<��<�!<r<�<�N<P��;$S�;�  �  ,��;z	�;$��;��;*<�4<��<��<��<!�<d�<K<h�<n< <t�<��<�<(H<]<+*< <mH<EI
<�� <۹�;�N�;�B�;��;:��;�5�;���;�<�L<Յ<?�<�<L�<�}�;���;,u�;I��;w��;��;��;BS�;�L<G<'�<N0<Q<��<�<B�<hN<�_<ST<i/<�<�u<��<�-<M�<��<�<3x<���;�D�;�Z�;���;���;n��;*$�;���;;<ީ<^�<<f?<U7<�_�;VP�;��;,�;���;��;��;���;�p	<��<z�<?<:<}�<v<*Y<u�< M<S�<��<|P<�<�$<>�<��<��<QZ<�I<�J�;J��;ݍ�;�Y�;�t�;Ԭ�;'�;� <��<�h<��<c�<��	<�<I�;G:�;92�;�$�;Hw�;���;�,�;F5<tf<�<M<ĺ<�.<�+<2<��<��<@E<��<�'<N�<Tv<F7<�S<a'<�m<�l
<N<#��;��;���;��;���;s��;�4�;�,<2w<��<ĳ<rD<�'<���;P�;���;�B�;Z�;���;�O�;H��;(f<s(<�<�?<�<��<N�<E�<M<&[<L<�#<�<pc<��<�<}<Dx<�<�R<�p�;���;���;�>�;�~�;�; ��;�S�;2<s<Y<��<�<<&��;e��;0��;���;�o�;s��;��;"��;�F	<|<P{<$�<�<]j<��<�"<˽<�<}W<�r<�<��<�<:�<QR<s<o#<F<c��;�7�;m�;���;���;�'�;:}�;���;��<D!<t�<ڞ<��	<r� <<��;I��;��;�  �  ���;ν;���;���;:�;��<wa<��<�)<�<I<�<��<@�<�m<�9<�<m�<��<��<c�<��<��<�<��;��;���;��;�·;��;��;�4�;���;w+<�H<�u<q	<i<)e�;�;���;�W�;/θ;��;^�;p��;�� <��<�<o<[�<u�<t�<�K<i<s�<L�<��<�<3�<r<��<��<L�<��<�<���;q��;��;���;�(�;���;D�;IC�;�. <-�<�v<��<@<���;b�;v��;���;WA�;#�;�G�;���;t��;��<�<x:<]�<��<�<P�<�<��<�<�	<%�<�<�D<��<L�<w�<�v<�X	<�F�;՞�; 9�;P��;�R�;&�;���;�&�;��;p<��
<*�<��<�s<�Q�;��;bs�;��;h�;�<�;��;�	�;?��;F*<��<�<R[<<�<	|<�)<l�<�$<�<%l<�I<��<��<��<#�<�<&�<߸<�?�;e��;��;w��;=�;7�;Af�;��;�.�;]V<u<��<V�	<�F<��;�]�;�;릹;��;,`�;���;���;,� <��< <�~<��<Y�<�<�M<	<��<�<�<� <�n<P\<��<B�<��<ԑ<��<�0�;��;E��;:[�;ø;i%�;h��;���;��;��<4@<�<�<�<�;E��;Q2�;;/�;R�;���;���;y9�;�O�;W<.�<�<�e<��<7�<+�<>X<b<+s<��<�`<��<H<Ț<�W<�_<�?<�!	<4��;�,�;q��;��;�Է;���;��;%��;XE�;-(<��
<�<=><�-<���;x�;#��;���;�  �  �#�;\��;���;6�;y��;��<�,<��<�S<I�<l<��<c <a<lk<n]<V�<�a<��<�<��<7<<��<��;���;��;�\�;cQ�;�y�;�y�;3��;h��;�<T1	<�w
<D< �;��;�a�;��;T6�;_G�;	P�;�V�;�;���;1�<6%<�O<��<;�<�<��<b<z�<˽<+<Z�<�<�<�,<��<�<��	<μ�;I�;�0�;�`�;�<�;��;͢�;M:�;���;��;?�<�t
<��	<f�<���;���;,�;�>�;�ާ;���;b��;IG�;��;� <� <�<Ǟ<�?<�O<
�<"<��<*�<�<
�<��<j_<�<��<DU<�_<�<���;E}�;���;wx�;!ʧ;9A�;OF�;�;��;��;�</�
<cY<� <!��; ��;(]�;GN�;�;B�;Fe�;���;���;��<�]<ø<t�<J.<��<��<�3<�:<'�<@�<��<��<�<*=<+�<]<29<�<���;��;��;#��;���;
®;�ſ;�(�;p�;'�<�]	<�
<�G<�Z�;�k�;��;k\�;*��;v��;̕�;���;�I�;���;��<W8<�_<<+�<��<��<�`<��<��<a<O�<�m<�<�<�<%�<�	<�p�;!��;L��;��;ۨ;戨;)9�;���;rA�; ��;�I<�=
<�	<�<�a�;���;���;K�;���;cW�; ��;���;ܴ�;�v <�<�y<�p<�<�<e�<��<m�<�q<��<2�<m<(<��<�<�<%)<��<���;�
�;�C�;=��;iK�;潪;���;]y�;t�;ӄ�;�q<_�
<f<�` <�7�;�2�;޺;�ԫ;�  �  'R)��-���L8��c�:O�=;�׉;�g�;���;h��;��;��;�;Դ�;O��;� �;7��;�N�;l�;���;�ս;R�;��;��(;"�:WPǹ��к�E�e�(�����͠���T8N�:q�';�qV;�^_;7�@;Ug ;�N-:�3�@�xY!��%���g	{����9���:(�\;�u�;f�;!1�;�+�;e"�;�R�;6��;i��;�y�;qD�;��;�)�;���;���;9�;@��;��f;Gq	;1�:��S��F��92#�W#������T�X�:)�:e�;;��^;<Z;}G/;���:6�_9�}�����P�&�3%��@޺���ѐp:��;Xpy;ȿ�;���;�<�; ��;���;fy�;���;�e�;���;�8�;��;E�;�	�;�;�ޮ;��;��H;^��:R{�8ጟ��l���'��<��κ�ʹ!�:��;|�K;߼a;��O;��;�~�:��y�[����V��e(��M�MC��5O{�$��:o>;�8�;�ȫ;K=�;m9�;�(�;7A�;��;��;qU�;���;c �;֬�;���;KM�;�$�;0�;�H�;�F); �:�lù��Ϻ���(�@A�󛟺[c}8���:�X(;'.W;{ `;^vA;�+;|U0:m�0�7��e� �wW%�&h�u�x���9[��:��\;ў�;���;�K�;A?�;o.�;IW�;��;���;�h�;A,�;?��;J�;ݠ�;���;-��;bJ�;6f;=�;�B:E�V�x���F$���#� J����X�)=:�N�:�:;	�];�XY;l.;t��:�S9m���O��ŗ'�_��x{ߺt^��"n:�;��x;�i�;;��;���;9#�;�z�;��;�[�;���;���;���;��;_��;��;���;�q�;��;*�G;Z��:҇�8Fm��*g�K�(�N�.�кFGӹ�'{:m�;�eJ;և`;��N;��;�=�:�l��'����P��  �  l��^������";&9��:F;���;ܬ;R{�;��;M��;�,�;4��;�w�;���;���;�C�;��;��;Z<�;n��;���;� �;F�1;�,�:��:����D�?@��	����|��g�9pF�:[�1;"__;�h;!!J;f;��b:T��qDǺX����<qߺ�6��s%:��;�c;��;\��;��;�P�;XQ�;��;9(�;�^�;�G�;��;t��;�]�;���;�.�;`B�;ע�;w�m;m�;әQ:���pҺ���J��FҺb�Ͳ?:��;.zE;�g;c;,!9;��:
b�9)Y�&��ح�j

�F︺o̐���:�!(;[�;鑣;�м;+��;��;l"�;��;w��;^7�;���;���;`�;}l�;7�;{��;�6�;��;V�P;�|�:�l�9�x����Ӄ��y�[���k��l��:Yn;z�T;#pj;�Y;$;S��:�iŶ;���O����O��k��J39��:��F;��;i=�;���;m�;RM�;m��;��;b��;�'�;BA�;&��;���;��;��;��;��;?F�;/]2;�*�:A�	�����8��Ÿ�a���=z��~�9q��:�[2;O`;��h;��J;�);��e:*�ํ�ź`��[
�D޺Փ4�f':'�;y0d;!ؘ;&��;���;d�;Z]�;ο�;�%�;�T�;�6�;���;g�;-7�;K��;���;��;
`�;.m;�;#�N:>o���Ӻ���F����ӺO �<:�;O�D;6�f;D5b;F8;�^�:�&�9T\�R��hW�ˬ
�[*�������ސ:��';4;�;�;�u�;�*�;�C�;���; ��;��;���;+K�;Va�;��;���;X��;�8�;�ɯ;���;��O;<��:�2�9�>|�7������ˉ��Ȭ��C.��6�:<;��S;<i;��W;��";uO�:f:�����v���  �  �����9���k��"�O:�;e�[;��;���;EO�;���;d��;d��;���;#N�;���;��;�T�;��;�>�;$�;׿;:b�;|�;��I;C�:�
:S�
�.s��Nf��8G���g��m:7
;c�M;Vx;Y=�;��d;�*;,`�:�օ9 �=�����k��Fmg����7���:� %;�v;$��;;��;_��;���;�@�;�m�;T��;�Q�;�A�;~|�;DQ�;�^�;���;1e�;4�;���;~�;��.;���:p%9O��J���¬��%Q��a9�o�:��#;�N`;,�;�{;��T;�8;���:g;ʸ�{����d��]�!�c�9�h�:�KA;�Ӈ;S��;�E�;҉�;$U�;yL�;c��;s/�;.;�;��;�&�;���;�=�;���;�M�;��;)�;@�e;l;�vw:|Q��慺S´�ȩ��G�	�j�:�-�:	O:;�n;�Z�;�r;rbA;Ő�:}�*:޹)薺�ǵ��|��ʢ�-S:��;��\;�w�;�[�;���; 3�;Y�;� �;T�;ݷ�;�-�;��;���;+2�;��;6z�;�'�;���;�;�rJ;�D�:�	:މ��n��gV���'���u]�"�o:��
;��N;�y;7��;,Te;8M+;�߾:C��9�
;�SĨ�|)��2e�@(8�:�n%;�w;�%�;��;��;��;�L�;�r�;ʟ�;�G�;�0�;Ud�;�1�;V8�;�k�;�0�;l��;�G�;�;Q^.;&�:w�9�"R�3ꭺ�t����T�7�	9���:��";	d_;�;�z;��S;�g;��:B��?m~��Ӵ����.$��)�9�-�:��@;I��;�a�;��;)�;���;���;!��;w��;j��;{,�;���;r�;=��;r��;���;���;�;0�d;	�;>�s:F�_��և��Ƕ��ş�*�	:y��:�9;FYm;���;�Sq;<@;�V�:r]&:��ט��  �  g��"?�8�&G:�g�:�P2;зv;^��;eJ�;�k�;c��;� �;�~�;tl�;~��;���;�;p��;\�;|�;y1�;�{�;���;�k�;kh;T�";߾:�
:�� 8������=9U;f:��:�^<;�"w;M�;ر�;]x�;�sX;6�;�N�:���9R�������f�9<9�:@{;��I;�E�;/��;�·;u|�;��;r �;��;���;�/�;u,�;���;C��;pf�;���;���;�չ;���;���;�<R;��;4��:*��97�b���`�)��92>�:6;��R;���;Ԅ�;2��;	P};�YD;� ;�%�:38�9��͸1��5�c:���:W�;�a;7��;��;�9�;D��;�}�;���;���;1��;�8�;0]�;���;���;N��;Z��;�0�;I߳;�;p�~;-�:;1��:!`b:�'D9�p�ul88,�":�B�:��&;�:f;���;C��;���;H`l;�b.;���:s9:W�8~v�l9�rJ:M��:3;�{w;#�;��;4��;�)�;Q��;���;���;<a�;�/�;Fw�;���;^��;���;���;6ξ;���;x��;q�h;�e#;R�:\:s�!8j��T�F9�h:�W�:	=;.�w;�{�;��;L؅;�3Y;��;5��:S2�90�������9AH�:��;fjJ;eu�;���;=�;���;�;<,�;���;���;&�;�;�~�;��;@�;p�;%��;5��;LC�;���;h�Q;�	;�2�:�q�9%��#B��^��9�u�:8N;r�Q;a4�;C�;TG�;�w|;N�C;& ;�[:G{9�F�r����:߿�:�;�x`;!+�;�9�;�ۼ;�J�;T�;@�;w��;G�;b��;���;�^�;���;�c�;;s�;@��;�q�;;��};i
:;�
�:k�^:��49� ����7:A:~�:P�%;�e;J�;!�; �;>k;�I-;���: 5:<r�8�  �  f�:\��:;��:B");ҲY;@(�;Sښ;+<�;��;h��;~}�;�;N%�;��;���;>`�;5��;/��;�`�;'��;���;�̨;�c�;=�;<�N;;@<�:4��:稯:�:�s;�	@;�v;��;y�;��;��;���;��X;��";���:A�:X�:{��:t<;]9;��j;<�;�j�;6;�;��;�!�;�K�;v��;��;�1�;�C�;�N�;�6�;���;���;!��;��;נ�;.��;3�p;�\?;̃;�1�:�=�:鱷:���:f$;o>S;([�;��;�;�s�;��;$8};=�F;�7;~��:�[�:$ĸ:c�:V�;�I;_${;)c�;pR�;��;r~�;r/�;9��;-��;b��;�o�;(�;c��;BN�;7u�;��;ꁺ;sJ�;�m�;�%�;0`;y,/;��;���:s��:|�:���:��.;<xe;5K�;��;��;��;mǎ;܁k;c�4;a�;�?�:6��:���:1R�:��); yZ;n��;�<�;柬;IU�;v
�;���;���;1��;k	�;�m�;W��;j�;o �;���;.Y�;ֶ;X�;���;�6�;ARO;��;8B�:n�:B��:n.�:;��@;�Lw;�g�;�q�;kY�;?s�;R�;�;Y;��#;��:W��:��:״�:�;��9;k;&4�;���;'\�;���;V4�;QW�;���;��;�'�;�2�;�6�;��;���;���;�u�;���;�^�;�s�;	p;�>; �;@��:0��:��:���:�B;rYR;��;@>�;�y�;J�;�6�;/j|;z
F;~|;]L�:��:�y�:���:m;GBI; }z;�;��;�/�;H�;y��;�O�;Uc�;�;�;���;��;@\�;R��;�;�e�;��;�ܭ;} �;Q��;�)_;tJ.;��;���:��:�p�:���:)�-;hXd;ɸ�;|$�;]N�;��;9�;�mj;�3;ڄ;>]�:�  �  ,}3;��5;�C;Z9X;jq;��;$�;��;�m�;�w�;a0�;>S�;7�;tc�;,��;A��;���;���;�G�;�~�;2[�;:{�;�^�;�;ڼk;,S;�e?;�#4;�5;JrD;�2a;���;h�;�z�;���;���;Hi�;7M�;��;�[q;z�O;�A:;�3;JQ9;��I;��`;��z;*.�;��;�V�;�é;s��;~L�;O�;�#�;���;��;���;���;=Q�;�̳;D�;]��;�a�;R͋;�~;�&d;��L;�m;;?�3;��9; �M;-n;�݊;w��;=}�;�ƶ;;��;Hz�;m�;�6�;+�e;��G;y�6;�+4;F;>;�@Q;kyi;�ǁ;�_�;۩�;���;��;W��;a&�;�y�;m��;d�;�(�;�"�;q��;���;��;��;DL�;���;���;�"u;J�[;��E;�f7;��3;*r>;�W;�z;���;X��;�1�;Zz�;;�;`g�;Eܓ;);*�Z;{}@;>_4;_6;��C; Y;,0r;��;hT�;&�;?զ;��; ��;Z��; ~�;���;H�;��;4'�;i�;���;�ܭ;���;�͚;8��;2�;Hl;�S;6�?;̪4;��5;�E;B�a;=�;�8�;uѩ;Z�;\�;�ů;ͩ�;l�;�r;4�P;)�:;��3;{�9;.ZJ;~9a;}{;l\�;�;cw�;>ݩ;�Ĳ;�W�;��;� �;�z�;��;���;���;)+�;���;T��;�a�;G �;M��;�q};x}c;L;5�:;�3;Ǵ8;"�L;�(m;�l�;�A�;�;W�;�C�;V�;�;EՅ;��d;�F;�6;�3;c�=;ÜP;�h;+r�;g�;�K�;�I�;�|�;VN�;��;��;�@�;���;l��;U��;p(�;!�;ir�;]s�;�ݝ;r3�;�"�;MGt;��Z;R
E;=y6;��2;r=;V;�y;&�;`�;j��;��;ڬ�;5ܥ;AU�;5 ~;e�Y;B�?;�  �  ���;;x;�Ps;&q;�6q;3�s;+�x;F��;cu�;��;��;Sͭ;��;v��;�e�;���;�y�;5ͪ;��;�x�;m��;�e;c>w;��r;q;׌q;YKt;�y;2�;��;#6�;�{�;��;~��;��;HR�;1��;���;⧨;��;��;TO�;� ~;��v;��r;'Yq;V)r;@Wu;j�{;�Z�;8�;B�;}��;Vu�;�z�;���;�.�;R}�;��;���;�;�?�;V�;�};EYv;��r;��q;*s;��v;��};�؄;=�;$�;���;�´;:�;6�;���;-#�;�;^�;��;l��;��;It{;�Yu;wTr;f�q;�/s;�Fw;J�~;���;��;���;���;?��;3V�;?��;�
�;���;ɾ�;L�;�ߔ;��;^�;�?z;m�t;**r;$�q;��s;�^x;�i�;m�;ꑑ;sH�;��;'��;���;~��;:0�;}Ϲ;拭;�ʟ;ޒ;�d�;��;\y;{t;��q;��q;&Lt;miy;�V�;lވ;��; ��;F?�;�Y�;Xr�;Y��;��;��;�9�;Uu�;�ڐ;I��;��;�w;�ss;��q;�r;��t;�z;)U�;�e�;���;�ʢ;Io�;"	�;\H�;R��;�;A�;^�;RN�;<�;���;×~;�&w;�7s;�q;��r;b�u;%�{;�z�;`�;v��;��;�y�;�w�;���;��;[e�;�˳;�y�;C�;,�;��;É|;m�u;yRr;IFq;jgr;@�u;��|;q�;L��;�|�;^�;�R�;î�;"�;�^�;���;��;��;䑖;2,�;�Â;0�z;ȳt;��q;J�p;�r;�v;�6~;���;�4�;b��;F�;1�;�ۿ;HG�;w��;y�;�E�;���;l�;b|�;���;�ey;��s;�Pq;� q;A�r;-vw;��;��;`�;�;ル;��;Y��;Od�;���;�G�;
�;�K�;?d�;,��;�  �  O,�;�I�;��;�o;��V;�B;g5;��3;!�@;i[;O"�;�y�;ɦ;�/�;��;��;��;���;o{w;lT;H�<;N�2;�%7;Z:F;�T\;w�u;��;��;���;e�;�
�;ഹ;���;��;���;��;+�;q��;h�;���;Q%�;��;c��;��;C�;�g;��O;k'=;��3;[7;U�H;Cjg;_2�;�T�;#�;�ӵ;W`�;���;.��;ݑ�; �k;�K;��8;��3;<;��M;��e;��;��;7�;=�;��;�i�;H�;Dx�;��;7��;?��;��;���;���;iY�;�d�;x�;Yv�;̞�;�jy;��_;�I;�9;Ԃ3;D�;;��Q;t;�-�;���;g�;�8�;���;��;D+�;�ւ;�`;2�C;`5;�&5;C�@;�!U;��m;���;�h�;rv�;�M�;&o�;9�;��;^��;�\�;�+�;)��;:8�;T`�;�,�;Gk�;&W�;���;��;�i�;��p;a�W;w�B;[�5;�4;��A;�E\;��;��; @�;��;`�;���;��;�k�;�Qx;�6U;�S=;d�3;#�7;��F;��\;�qv;�1�;N0�;}ʞ;�W�;�U�;0�;* �;i�;�H�;>�;��;K%�;���;O�;�w�;�:�;t*�;͍;�&�;9h;�+P;0�=;64;�@7;��H;�g;]=�;�X�;.�;�ɵ;gO�;���;Ua�;l�;�Wk;XzK;�+8;�N3;W�;;NM;P�d;��~;�)�;��; ס;�!�;���;�|�;&
�;��;���;�(�;G��;�u�;���;���;h�;���;�!�;�J�;��x;+_;�\H;	Q8;ʻ2;X�:;Q;�+s;���;)'�;(�;���;�;9��;¯�;_^�;�_;�C;d�4;QL4;$@;tJT;
m;���;���;� �;�Ӥ;��;ݶ�;���;��;'��;:��;1�;ͳ�;�߿;���;��;��;�  �  :a�;s��;ك;��V;��&;ɥ�:|��:)�:��:�;��6;[}m;Yv�;v<�;rG�;l�;W{�;�ba;�+;��:�p�:���:�y�:�A;�1;.b;��;&�;��;\��;M��;c^�;W"�;��;S��;��;�K�;�c�;Z?�;��;p;;h��;�4�;�;�)x;U�F;�
;�:�ȶ:�в:ۈ�:c�;�I;�;}��;���;�n�;���;�ɂ;w�O;};B�:�ߵ:� �:�.�:z�;B;scs;���;Щ�;��;0A�;�b�;�7�;w��;
��;*r�;�Q�;�&�;���;�3�;���;%�;���;.��;��;/h;�7;�W
;t�:��:��:���:UD&;<\;{Z�;�N�;.��;_�;�N�;�ot;��=;�;Is�:�|�:�8�:�c�:H";e<R;f��;U�;��;ʋ�;���;i�;�d�;�C�; ��;t}�;?	�;���;���;ҫ�;#��;�ø;�̫;_%�;>�;}�W;�V';�4�:G�:��:S��:��;5�7;Uln;a��;;å;o�;��;6Jb;��+;�B�:n��:���:K��:��;��1;Ӣb;�Z�;}l�;�;��;E*�;��;�r�;6��;�1�;�m�;-��;��;H��;���;F�;���;O}�;�N�;G�x;�WG;�o;��:`�:�M�:���:��;��I;��;q~�;���;�]�;�u�;˪�;I�O;��;�u�:b��:� �:��:�0;�fA;��r;���;�H�;6I�;5ٽ;"��;���;��;��;-�;���;[��;p�;C��;���;Ļ;+E�;�2�;���;z�g;pR6;��	;���:}�:�d�:V�:W%;�E[;�ۇ;�͛;0	�;�l�;�Α;zts;9�<;�
;��:ܽ�:���:��:ur!;�eQ;22�;\x�;w��;g�;k^�;_��;���;v��;�f�;D��;k��;9 �;�H�;92�;37�;�S�;�  �  �(�; �;�s;Om.;
!�:^�;:X��8/���G�8��@:}6�:�1;�Jn;j݋;]�;d�;��a;`";���:i�:v�7by�<�T9�fk:T��:�>;�Ӏ;w%�;P��;^�;t��;���;ا�;v�;2�;���;WB�;:��;�V�;��;���;�/�; #�;[��;�];M�;���:���9>o����ŸJ��9��:�E;D�G;��;��;���;J�;[�N;�;�ؔ:3&�9ڐ�|17�}��9�:�~;V;��;��;hѺ;�_�;���;���;�;���;xP�;0[�;3��;��;:,�;���;�	�;��;TP�;̫�;spF;#
;���:��9kļ��~h�ID:曰:q;/\;��;NN�;6ٍ;Qu;`x9;b�:Ծ\:Ϻ+9�Q�G�8؉(:�Q�:�r';�ul;x`�;�D�;�;��;��;���;(��;}��;�=�;)t�;$��;9��;^l�;*��;R!�;ђ�;�|�;9�s;3/;B��:��>:�i�8i��}��8�zD:�:;2;,Do;�[�;���;t�;��b;��";+��:�:2�7�۸@�_9��m:l��:�>;��;�l�;�ܴ;��;7+�;���;���;���;TW�;p=�;Z��;��;��;DZ�;eJ�;�{�;�j�; ��;�]; 
;�g�:���9z)~��轸#2�9WW�:[;ΛG;h�;��;�;I2�;
�N;��;(�:)��9�.���W�%��9�:*�;�eU;�V�;��;�m�; ��;s��;b0�;ϫ�;�J�;���;g��;b�;Ƥ�;H��;t�;���;���;V��;�U�;��E;�U ;�:(؉9T�ָ`eⷙI�9���:Au;c|[;e�;�ɑ;.U�;�t;wy8;��:��X:�@9?,�x�M8�1%:���:7�&;z�k;Q�;)ӭ;�2�;���;L��;�[�;�q�;��;G��;��;vj�;�p�;��;<_�;۲�;�  �  ���;f5�;�wW;uM;�->:-fŹ� ��9���H
����ʹ#�7:��:��C;"8s;���;Ik;V�5;�>�:���9��Ϋ��Oµ�����l"�DR�:�s;
\i;(��;R�;)��;���;���;�z�;���;>=�;0��;���;���;l�;p��;:��;5�;��;���;e<;Ny�:'��90�.�ߓ���Ͳ�J�r�=3��Ǒ:� ;�sW;R�|;��~;g7];�A;�: ~�8�]�������WjD�
�d9�ȼ:@�3;9�;�6�;]�;�;C��;|}�;�[�;���;I_�;���;���;ϩ�;M_�;��;r�;��;k�;��r;ؕ ;N	�:l��N�o��䱺����R�/���9��:/;k�g;��;��w;#oK;c�;o�^: ����.�����u�\d���:n �:q1O;�ʍ;�5�;&�;N�;]��;�7�;��;
��;G:�;��;z�;o�;k�;=��;���;��;Y��;?X;�;�CA:"��B�����'O��ˡùƑ;:�:�D;�8t;V5�;VHl;j�6;�"�:>9�9��9���@��󨁺O�����:�
;��i;��;:�;���;9�;�B�;���;	�;{��;�C�;�L�;I�;�b�;�<�;��;_�;KK�;��;��<;lV�:���9�v-������S���/r��w*���:8;nmW;:�|;ޘ~;�];};�J�:;{�8ݳ^���������5�F�]�[9@��:3;]��;�ע;C��;3��;#��;��;j��;��;���;��;}�;>H�;� �;n~�;�;�\�;��;8�q;$�;S��:�u$���r�Ҍ��vI��uC3�R>�98��:.;�f;N]�;ّv;SgJ;��;I�Z:�F��> ���O���v�����[�:�z�:V\N;^�;�ū;Ȳ�;j��;S�;̺�;�/�;�z�;��;W�;t��;��;ˎ�;�e�;�v�;�  �  S�;}i�;� A;���:[��8ٕ�c��C�����\��1	U8Gܳ:a�&;�Y;6i;G_Q;�\;Qˍ:�$w������)	����U�8k����9#��:|�T;2��;(L�;c%�;:�;�;���;�Z�;�V�; ��;�Q�;>��;���;qA�;4��;���;!��;��z;��";Y�:���	$��c��7@��人vI�aJ:*J�:�;;?�c;�1f;�+B;H4�:��*:,&���غ�2�����3̺����Tf:��;�sr;��;���;+��;*D�;9r�;%��;���;0b�;ϓ�;|p�;��;�w�;�,�;��;<Y�;+�;�Q_;_�;1:�~F�C-�
��h�%|��H+���y:@L;�M;si;��^;��.;��:��]9݄��h��/��}��jV����f�w%�:|�7;���;���;��;M"�;��;l��;c��;@6�;�3�;x�;pF�;_��;�D�;�	�;���;���;�Ί;.�A;i�:�=�8mG���� �6(�� �,���g��8ϵ: �';s�Z;�"j;�aR;�Y;O��:|h��Y��;����A�h�6��9W��:X�U;O��;&��;Dn�;���;�j�;m:�;���;���;�A�;��;')�;�C�;��;
�;�̻;P��;�t{;�*#;
�:����w���y�q��R�k�H���:�X�:��;;�c; f;f�A;��:��):ŋ'��xٺ���3~��Hͺ�/�)�c:?9;Ծq;h!�;l)�;��;���;E	�;��;���;���;n-�;��;\��;��;��;���;��;y��;��^;��;SQ:�I�w��4��cJ��X��(�Ĺ�u:�B;wL;�ch;�~];��-;
��:�DN9"��;��N�����I ��ઍ���:��6;��;�'�;a��;���;ȝ�;�q�;��;c��;״�;׆�;��;B�;%��;c��;���;�  �  �ϩ;���;�v8; ��:�������Tf�ZW)�e!�T���߾;���:q;��P;�h`;LH;��;�g: ����׺���X(�˳������09P�:�*M;�=�;U�;&��;]�;#��;���;ڽ�;���;��;��;�Z�;���;� �;�o�;
��;�̟;�yt;=;9�Y:�;�έ�����x&�j]�^d���f�9��:$02;�%[;Xh];X�8;��:Q��9[h�YP��OX$��8"�+�BNA��t0: �;�k;�{�;#��;8��;J"�;l;�;w�;:E�;Ӓ�;���;G��;���;)K�;'�;���;9*�;{��;]�W;Η�:���9갅�os��H&��Z��;�9m��D:^k;'D;�`;��U;��$;3\�:ra��������:1(�ȴ�Y�Ǻ���{�:�.;��;���;�H�;���;���;h��;�;�x�;Ha�;�B�;G��;�j�;5!�;���;.M�;*8�;��;=9;M��:����b�������(�B��Է�C�,���:q;?�Q;Qna;�!I;ʯ;	�k:���8ֺ-�
�'���
�M���:94��:�M;��;eJ�;��;�Y�;�A�;���;��;>��;7q�;��;F��;2�;$q�;w��;'�;��;|�t;Ņ;�x[:ɳ������;&��-����O�9'�:�)2;�[;�F];�X8;��:���9q�i�E���$��"��?��C� �-:�3;��j;9�;	,�;')�;���;���;#��;*��;�*�;jb�;si�;}<�;���;���;�6�;�Ҳ;�F�;�(W;R3�:f�9�2���>��'��= �溫U"��@:�`;9C;��_;3�T;>�#;�S�:��z���I��w)�َ��ɺZ��,ٗ:��-;k5�;4��;�־;�m�;]|�;
)�;���;M��;���;���;I;�;���;��;wb�;'��;�  �  S�;}i�;� A;���:[��8ٕ�c��C�����\��1	U8Gܳ:a�&;�Y;6i;G_Q;�\;Qˍ:�$w������)	����U�8k����9#��:|�T;2��;(L�;c%�;:�;�;���;�Z�;�V�; ��;�Q�;>��;���;qA�;4��;���;!��;��z;��";Y�:���	$��c��7@��人vI�aJ:*J�:�;;?�c;�1f;�+B;H4�:��*:,&���غ�2�����3̺����Tf:��;�sr;��;���;+��;*D�;9r�;%��;���;0b�;ϓ�;|p�;��;�w�;�,�;��;<Y�;+�;�Q_;_�;1:�~F�C-�
��h�%|��H+���y:@L;�M;si;��^;��.;��:��]9݄��h��/��}��jV����f�w%�:|�7;���;���;��;M"�;��;l��;c��;@6�;�3�;x�;pF�;_��;�D�;�	�;���;���;�Ί;.�A;i�:�=�8mG���� �6(�� �,���g��8ϵ: �';s�Z;�"j;�aR;�Y;O��:|h��Y��;����A�h�6��9W��:X�U;O��;&��;Dn�;���;�j�;m:�;���;���;�A�;��;')�;�C�;��;
�;�̻;P��;�t{;�*#;
�:����w���y�q��R�k�H���:�X�:��;;�c; f;f�A;��:��):ŋ'��xٺ���3~��Hͺ�/�)�c:?9;Ծq;h!�;l)�;��;���;E	�;��;���;���;n-�;��;\��;��;��;���;��;y��;��^;��;SQ:�I�w��4��cJ��X��(�Ĺ�u:�B;wL;�ch;�~];��-;
��:�DN9"��;��N�����I ��ઍ���:��6;��;�'�;a��;���;ȝ�;�q�;��;c��;״�;׆�;��;B�;%��;c��;���;�  �  ���;f5�;�wW;uM;�->:-fŹ� ��9���H
����ʹ#�7:��:��C;"8s;���;Ik;V�5;�>�:���9��Ϋ��Oµ�����l"�DR�:�s;
\i;(��;R�;)��;���;���;�z�;���;>=�;0��;���;���;l�;p��;:��;5�;��;���;e<;Ny�:'��90�.�ߓ���Ͳ�J�r�=3��Ǒ:� ;�sW;R�|;��~;g7];�A;�: ~�8�]�������WjD�
�d9�ȼ:@�3;9�;�6�;]�;�;C��;|}�;�[�;���;I_�;���;���;ϩ�;M_�;��;r�;��;k�;��r;ؕ ;N	�:l��N�o��䱺����R�/���9��:/;k�g;��;��w;#oK;c�;o�^: ����.�����u�\d���:n �:q1O;�ʍ;�5�;&�;N�;]��;�7�;��;
��;G:�;��;z�;o�;k�;=��;���;��;Y��;?X;�;�CA:"��B�����'O��ˡùƑ;:�:�D;�8t;V5�;VHl;j�6;�"�:>9�9��9���@��󨁺O�����:�
;��i;��;:�;���;9�;�B�;���;	�;{��;�C�;�L�;I�;�b�;�<�;��;_�;KK�;��;��<;lV�:���9�v-������S���/r��w*���:8;nmW;:�|;ޘ~;�];};�J�:;{�8ݳ^���������5�F�]�[9@��:3;]��;�ע;C��;3��;#��;��;j��;��;���;��;}�;>H�;� �;n~�;�;�\�;��;8�q;$�;S��:�u$���r�Ҍ��vI��uC3�R>�98��:.;�f;N]�;ّv;SgJ;��;I�Z:�F��> ���O���v�����[�:�z�:V\N;^�;�ū;Ȳ�;j��;S�;̺�;�/�;�z�;��;W�;t��;��;ˎ�;�e�;�v�;�  �  �(�; �;�s;Om.;
!�:^�;:X��8/���G�8��@:}6�:�1;�Jn;j݋;]�;d�;��a;`";���:i�:v�7by�<�T9�fk:T��:�>;�Ӏ;w%�;P��;^�;t��;���;ا�;v�;2�;���;WB�;:��;�V�;��;���;�/�; #�;[��;�];M�;���:���9>o����ŸJ��9��:�E;D�G;��;��;���;J�;[�N;�;�ؔ:3&�9ڐ�|17�}��9�:�~;V;��;��;hѺ;�_�;���;���;�;���;xP�;0[�;3��;��;:,�;���;�	�;��;TP�;̫�;spF;#
;���:��9kļ��~h�ID:曰:q;/\;��;NN�;6ٍ;Qu;`x9;b�:Ծ\:Ϻ+9�Q�G�8؉(:�Q�:�r';�ul;x`�;�D�;�;��;��;���;(��;}��;�=�;)t�;$��;9��;^l�;*��;R!�;ђ�;�|�;9�s;3/;B��:��>:�i�8i��}��8�zD:�:;2;,Do;�[�;���;t�;��b;��";+��:�:2�7�۸@�_9��m:l��:�>;��;�l�;�ܴ;��;7+�;���;���;���;TW�;p=�;Z��;��;��;DZ�;eJ�;�{�;�j�; ��;�]; 
;�g�:���9z)~��轸#2�9WW�:[;ΛG;h�;��;�;I2�;
�N;��;(�:)��9�.���W�%��9�:*�;�eU;�V�;��;�m�; ��;s��;b0�;ϫ�;�J�;���;g��;b�;Ƥ�;H��;t�;���;���;V��;�U�;��E;�U ;�:(؉9T�ָ`eⷙI�9���:Au;c|[;e�;�ɑ;.U�;�t;wy8;��:��X:�@9?,�x�M8�1%:���:7�&;z�k;Q�;)ӭ;�2�;���;L��;�[�;�q�;��;G��;��;vj�;�p�;��;<_�;۲�;�  �  :a�;s��;ك;��V;��&;ɥ�:|��:)�:��:�;��6;[}m;Yv�;v<�;rG�;l�;W{�;�ba;�+;��:�p�:���:�y�:�A;�1;.b;��;&�;��;\��;M��;c^�;W"�;��;S��;��;�K�;�c�;Z?�;��;p;;h��;�4�;�;�)x;U�F;�
;�:�ȶ:�в:ۈ�:c�;�I;�;}��;���;�n�;���;�ɂ;w�O;};B�:�ߵ:� �:�.�:z�;B;scs;���;Щ�;��;0A�;�b�;�7�;w��;
��;*r�;�Q�;�&�;���;�3�;���;%�;���;.��;��;/h;�7;�W
;t�:��:��:���:UD&;<\;{Z�;�N�;.��;_�;�N�;�ot;��=;�;Is�:�|�:�8�:�c�:H";e<R;f��;U�;��;ʋ�;���;i�;�d�;�C�; ��;t}�;?	�;���;���;ҫ�;#��;�ø;�̫;_%�;>�;}�W;�V';�4�:G�:��:S��:��;5�7;Uln;a��;;å;o�;��;6Jb;��+;�B�:n��:���:K��:��;��1;Ӣb;�Z�;}l�;�;��;E*�;��;�r�;6��;�1�;�m�;-��;��;H��;���;F�;���;O}�;�N�;G�x;�WG;�o;��:`�:�M�:���:��;��I;��;q~�;���;�]�;�u�;˪�;I�O;��;�u�:b��:� �:��:�0;�fA;��r;���;�H�;6I�;5ٽ;"��;���;��;��;-�;���;[��;p�;C��;���;Ļ;+E�;�2�;���;z�g;pR6;��	;���:}�:�d�:V�:W%;�E[;�ۇ;�͛;0	�;�l�;�Α;zts;9�<;�
;��:ܽ�:���:��:ur!;�eQ;22�;\x�;w��;g�;k^�;_��;���;v��;�f�;D��;k��;9 �;�H�;92�;37�;�S�;�  �  O,�;�I�;��;�o;��V;�B;g5;��3;!�@;i[;O"�;�y�;ɦ;�/�;��;��;��;���;o{w;lT;H�<;N�2;�%7;Z:F;�T\;w�u;��;��;���;e�;�
�;ഹ;���;��;���;��;+�;q��;h�;���;Q%�;��;c��;��;C�;�g;��O;k'=;��3;[7;U�H;Cjg;_2�;�T�;#�;�ӵ;W`�;���;.��;ݑ�; �k;�K;��8;��3;<;��M;��e;��;��;7�;=�;��;�i�;H�;Dx�;��;7��;?��;��;���;���;iY�;�d�;x�;Yv�;̞�;�jy;��_;�I;�9;Ԃ3;D�;;��Q;t;�-�;���;g�;�8�;���;��;D+�;�ւ;�`;2�C;`5;�&5;C�@;�!U;��m;���;�h�;rv�;�M�;&o�;9�;��;^��;�\�;�+�;)��;:8�;T`�;�,�;Gk�;&W�;���;��;�i�;��p;a�W;w�B;[�5;�4;��A;�E\;��;��; @�;��;`�;���;��;�k�;�Qx;�6U;�S=;d�3;#�7;��F;��\;�qv;�1�;N0�;}ʞ;�W�;�U�;0�;* �;i�;�H�;>�;��;K%�;���;O�;�w�;�:�;t*�;͍;�&�;9h;�+P;0�=;64;�@7;��H;�g;]=�;�X�;.�;�ɵ;gO�;���;Ua�;l�;�Wk;XzK;�+8;�N3;W�;;NM;P�d;��~;�)�;��; ס;�!�;���;�|�;&
�;��;���;�(�;G��;�u�;���;���;h�;���;�!�;�J�;��x;+_;�\H;	Q8;ʻ2;X�:;Q;�+s;���;)'�;(�;���;�;9��;¯�;_^�;�_;�C;d�4;QL4;$@;tJT;
m;���;���;� �;�Ӥ;��;ݶ�;���;��;'��;:��;1�;ͳ�;�߿;���;��;��;�  �  ���;;x;�Ps;&q;�6q;3�s;+�x;F��;cu�;��;��;Sͭ;��;v��;�e�;���;�y�;5ͪ;��;�x�;m��;�e;c>w;��r;q;׌q;YKt;�y;2�;��;#6�;�{�;��;~��;��;HR�;1��;���;⧨;��;��;TO�;� ~;��v;��r;'Yq;V)r;@Wu;j�{;�Z�;8�;B�;}��;Vu�;�z�;���;�.�;R}�;��;���;�;�?�;V�;�};EYv;��r;��q;*s;��v;��};�؄;=�;$�;���;�´;:�;6�;���;-#�;�;^�;��;l��;��;It{;�Yu;wTr;f�q;�/s;�Fw;J�~;���;��;���;���;?��;3V�;?��;�
�;���;ɾ�;L�;�ߔ;��;^�;�?z;m�t;**r;$�q;��s;�^x;�i�;m�;ꑑ;sH�;��;'��;���;~��;:0�;}Ϲ;拭;�ʟ;ޒ;�d�;��;\y;{t;��q;��q;&Lt;miy;�V�;lވ;��; ��;F?�;�Y�;Xr�;Y��;��;��;�9�;Uu�;�ڐ;I��;��;�w;�ss;��q;�r;��t;�z;)U�;�e�;���;�ʢ;Io�;"	�;\H�;R��;�;A�;^�;RN�;<�;���;×~;�&w;�7s;�q;��r;b�u;%�{;�z�;`�;v��;��;�y�;�w�;���;��;[e�;�˳;�y�;C�;,�;��;É|;m�u;yRr;IFq;jgr;@�u;��|;q�;L��;�|�;^�;�R�;î�;"�;�^�;���;��;��;䑖;2,�;�Â;0�z;ȳt;��q;J�p;�r;�v;�6~;���;�4�;b��;F�;1�;�ۿ;HG�;w��;y�;�E�;���;l�;b|�;���;�ey;��s;�Pq;� q;A�r;-vw;��;��;`�;�;ル;��;Y��;Od�;���;�G�;
�;�K�;?d�;,��;�  �  ,}3;��5;�C;Z9X;jq;��;$�;��;�m�;�w�;a0�;>S�;7�;tc�;,��;A��;���;���;�G�;�~�;2[�;:{�;�^�;�;ڼk;,S;�e?;�#4;�5;JrD;�2a;���;h�;�z�;���;���;Hi�;7M�;��;�[q;z�O;�A:;�3;JQ9;��I;��`;��z;*.�;��;�V�;�é;s��;~L�;O�;�#�;���;��;���;���;=Q�;�̳;D�;]��;�a�;R͋;�~;�&d;��L;�m;;?�3;��9; �M;-n;�݊;w��;=}�;�ƶ;;��;Hz�;m�;�6�;+�e;��G;y�6;�+4;F;>;�@Q;kyi;�ǁ;�_�;۩�;���;��;W��;a&�;�y�;m��;d�;�(�;�"�;q��;���;��;��;DL�;���;���;�"u;J�[;��E;�f7;��3;*r>;�W;�z;���;X��;�1�;Zz�;;�;`g�;Eܓ;);*�Z;{}@;>_4;_6;��C; Y;,0r;��;hT�;&�;?զ;��; ��;Z��; ~�;���;H�;��;4'�;i�;���;�ܭ;���;�͚;8��;2�;Hl;�S;6�?;̪4;��5;�E;B�a;=�;�8�;uѩ;Z�;\�;�ů;ͩ�;l�;�r;4�P;)�:;��3;{�9;.ZJ;~9a;}{;l\�;�;cw�;>ݩ;�Ĳ;�W�;��;� �;�z�;��;���;���;)+�;���;T��;�a�;G �;M��;�q};x}c;L;5�:;�3;Ǵ8;"�L;�(m;�l�;�A�;�;W�;�C�;V�;�;EՅ;��d;�F;�6;�3;c�=;ÜP;�h;+r�;g�;�K�;�I�;�|�;VN�;��;��;�@�;���;l��;U��;p(�;!�;ir�;]s�;�ݝ;r3�;�"�;MGt;��Z;R
E;=y6;��2;r=;V;�y;&�;`�;j��;��;ڬ�;5ܥ;AU�;5 ~;e�Y;B�?;�  �  f�:\��:;��:B");ҲY;@(�;Sښ;+<�;��;h��;~}�;�;N%�;��;���;>`�;5��;/��;�`�;'��;���;�̨;�c�;=�;<�N;;@<�:4��:稯:�:�s;�	@;�v;��;y�;��;��;���;��X;��";���:A�:X�:{��:t<;]9;��j;<�;�j�;6;�;��;�!�;�K�;v��;��;�1�;�C�;�N�;�6�;���;���;!��;��;נ�;.��;3�p;�\?;̃;�1�:�=�:鱷:���:f$;o>S;([�;��;�;�s�;��;$8};=�F;�7;~��:�[�:$ĸ:c�:V�;�I;_${;)c�;pR�;��;r~�;r/�;9��;-��;b��;�o�;(�;c��;BN�;7u�;��;ꁺ;sJ�;�m�;�%�;0`;y,/;��;���:s��:|�:���:��.;<xe;5K�;��;��;��;mǎ;܁k;c�4;a�;�?�:6��:���:1R�:��); yZ;n��;�<�;柬;IU�;v
�;���;���;1��;k	�;�m�;W��;j�;o �;���;.Y�;ֶ;X�;���;�6�;ARO;��;8B�:n�:B��:n.�:;��@;�Lw;�g�;�q�;kY�;?s�;R�;�;Y;��#;��:W��:��:״�:�;��9;k;&4�;���;'\�;���;V4�;QW�;���;��;�'�;�2�;�6�;��;���;���;�u�;���;�^�;�s�;	p;�>; �;@��:0��:��:���:�B;rYR;��;@>�;�y�;J�;�6�;/j|;z
F;~|;]L�:��:�y�:���:m;GBI; }z;�;��;�/�;H�;y��;�O�;Uc�;�;�;���;��;@\�;R��;�;�e�;��;�ܭ;} �;Q��;�)_;tJ.;��;���:��:�p�:���:)�-;hXd;ɸ�;|$�;]N�;��;9�;�mj;�3;ڄ;>]�:�  �  g��"?�8�&G:�g�:�P2;зv;^��;eJ�;�k�;c��;� �;�~�;tl�;~��;���;�;p��;\�;|�;y1�;�{�;���;�k�;kh;T�";߾:�
:�� 8������=9U;f:��:�^<;�"w;M�;ر�;]x�;�sX;6�;�N�:���9R�������f�9<9�:@{;��I;�E�;/��;�·;u|�;��;r �;��;���;�/�;u,�;���;C��;pf�;���;���;�չ;���;���;�<R;��;4��:*��97�b���`�)��92>�:6;��R;���;Ԅ�;2��;	P};�YD;� ;�%�:38�9��͸1��5�c:���:W�;�a;7��;��;�9�;D��;�}�;���;���;1��;�8�;0]�;���;���;N��;Z��;�0�;I߳;�;p�~;-�:;1��:!`b:�'D9�p�ul88,�":�B�:��&;�:f;���;C��;���;H`l;�b.;���:s9:W�8~v�l9�rJ:M��:3;�{w;#�;��;4��;�)�;Q��;���;���;<a�;�/�;Fw�;���;^��;���;���;6ξ;���;x��;q�h;�e#;R�:\:s�!8j��T�F9�h:�W�:	=;.�w;�{�;��;L؅;�3Y;��;5��:S2�90�������9AH�:��;fjJ;eu�;���;=�;���;�;<,�;���;���;&�;�;�~�;��;@�;p�;%��;5��;LC�;���;h�Q;�	;�2�:�q�9%��#B��^��9�u�:8N;r�Q;a4�;C�;TG�;�w|;N�C;& ;�[:G{9�F�r����:߿�:�;�x`;!+�;�9�;�ۼ;�J�;T�;@�;w��;G�;b��;���;�^�;���;�c�;;s�;@��;�q�;;��};i
:;�
�:k�^:��49� ����7:A:~�:P�%;�e;J�;!�; �;>k;�I-;���: 5:<r�8�  �  �����9���k��"�O:�;e�[;��;���;EO�;���;d��;d��;���;#N�;���;��;�T�;��;�>�;$�;׿;:b�;|�;��I;C�:�
:S�
�.s��Nf��8G���g��m:7
;c�M;Vx;Y=�;��d;�*;,`�:�օ9 �=�����k��Fmg����7���:� %;�v;$��;;��;_��;���;�@�;�m�;T��;�Q�;�A�;~|�;DQ�;�^�;���;1e�;4�;���;~�;��.;���:p%9O��J���¬��%Q��a9�o�:��#;�N`;,�;�{;��T;�8;���:g;ʸ�{����d��]�!�c�9�h�:�KA;�Ӈ;S��;�E�;҉�;$U�;yL�;c��;s/�;.;�;��;�&�;���;�=�;���;�M�;��;)�;@�e;l;�vw:|Q��慺S´�ȩ��G�	�j�:�-�:	O:;�n;�Z�;�r;rbA;Ő�:}�*:޹)薺�ǵ��|��ʢ�-S:��;��\;�w�;�[�;���; 3�;Y�;� �;T�;ݷ�;�-�;��;���;+2�;��;6z�;�'�;���;�;�rJ;�D�:�	:މ��n��gV���'���u]�"�o:��
;��N;�y;7��;,Te;8M+;�߾:C��9�
;�SĨ�|)��2e�@(8�:�n%;�w;�%�;��;��;��;�L�;�r�;ʟ�;�G�;�0�;Ud�;�1�;V8�;�k�;�0�;l��;�G�;�;Q^.;&�:w�9�"R�3ꭺ�t����T�7�	9���:��";	d_;�;�z;��S;�g;��:B��?m~��Ӵ����.$��)�9�-�:��@;I��;�a�;��;)�;���;���;!��;w��;j��;{,�;���;r�;=��;r��;���;���;�;0�d;	�;>�s:F�_��և��Ƕ��ş�*�	:y��:�9;FYm;���;�Sq;<@;�V�:r]&:��ט��  �  l��^������";&9��:F;���;ܬ;R{�;��;M��;�,�;4��;�w�;���;���;�C�;��;��;Z<�;n��;���;� �;F�1;�,�:��:����D�?@��	����|��g�9pF�:[�1;"__;�h;!!J;f;��b:T��qDǺX����<qߺ�6��s%:��;�c;��;\��;��;�P�;XQ�;��;9(�;�^�;�G�;��;t��;�]�;���;�.�;`B�;ע�;w�m;m�;әQ:���pҺ���J��FҺb�Ͳ?:��;.zE;�g;c;,!9;��:
b�9)Y�&��ح�j

�F︺o̐���:�!(;[�;鑣;�м;+��;��;l"�;��;w��;^7�;���;���;`�;}l�;7�;{��;�6�;��;V�P;�|�:�l�9�x����Ӄ��y�[���k��l��:Yn;z�T;#pj;�Y;$;S��:�iŶ;���O����O��k��J39��:��F;��;i=�;���;m�;RM�;m��;��;b��;�'�;BA�;&��;���;��;��;��;��;?F�;/]2;�*�:A�	�����8��Ÿ�a���=z��~�9q��:�[2;O`;��h;��J;�);��e:*�ํ�ź`��[
�D޺Փ4�f':'�;y0d;!ؘ;&��;���;d�;Z]�;ο�;�%�;�T�;�6�;���;g�;-7�;K��;���;��;
`�;.m;�;#�N:>o���Ӻ���F����ӺO �<:�;O�D;6�f;D5b;F8;�^�:�&�9T\�R��hW�ˬ
�[*�������ސ:��';4;�;�;�u�;�*�;�C�;���; ��;��;���;+K�;Va�;��;���;X��;�8�;�ɯ;���;��O;<��:�2�9�>|�7������ˉ��Ȭ��C.��6�:<;��S;<i;��W;��";uO�:f:�����v���  �  �Iw���m�h�T�VV0����bܴ���L�
����I�9�ģ:,X�:��;�;�;�n;��;56;R;�C�:��:�\�7�H˺xwm���ǻ<W�F+9��[��uq�K�v��-k�a�P�`s,��b�N̻�Z��#����붻U���J�:>A��`���s�� v�"g�8�I��d"�N��P6��3���F�5j0:���:5�:e@
;�;��;1;g;�.;]��:��:�O:1T���s�����u���E��Nd���t���t��}c���D��U�����G������b��ƻ�/�,�'�P�L�h�h�?Sv���r�~�^�_W=����л��}�� 序3��X�:���:iX;�;��;
J;;qV;�;af�:�ί::��9�{�R<�E2���� �Ғ+�-$Q�I�k���v� �p�u�Z��8�͓��*߻�᭻����)��tػ�c��4�QW��o��w���m�J�T��#0��u��|��A�K��4��of�9#U�:���:�|;�;$�;IA;"�;��;��;���:ta�:��7�+ʺ��l�cǻ�9�d9���[�MWq���v��
k��cP��I,��5�i�˻����mT��D���Oh�^�A���`���s���u�A�f��I�NC"����v��e��$�^N1:�O�:di�:0K
;��;��;(�;%�;�
;�:B�:9JM:`D���oZ��;仵��J�E�ƃd�a-u���t�V�c�6E����G���Ż�����ڡ��}ƻf�H0(���L���h��|v���r��^�#|=��/�9.ѻ/i~�ao�'�
����:�j�:L�;|�;�;Ae;v!;p;d�;��:��:��9�t~�-�<�n����� �-�+�!aQ�X�k�zw�q���Z�~/9���� �߻����V����˪��ٻ���P 5�a�W��Go��  �  n�n���e��KM���)�e� �K���=D�#4��wk�9ė�:���:�;E�;�;g�;��;'�
;�m;��:�r�:!%8 ºd�����
�r2���S�:�h�N2n���b�]�H���%��� �{1û�M��┻�`�����zG��!:�/�X�bk�Hm���^�EeB�}s���%O��@$�_
�g0:�4�:���:X�;I�;�;� ;[�;�	;OS�:�:��M:��ѹo��u��^ۻ<��$]>��#\��Cl�R�k�Z[��=�C3���Y�����f��������R�!�.@E�Zm`�d�m�`(j��V��x6�4���ɻ��s���ں�_θT̀:���:T�;j#;p;�];�;R;�;��:6g�:���9y�m�A^4�����\���AO%�T�I��Hc�n�2h�;�R�2�<��:�ջ�����,����ϻ����-��O�c�f��Ln�iKe��M�"�)��� �������C�)���U��9F)�:��:R�;��;�;V;J�;��;�-;m�:�Ì:�:8@�����c��ۿ�6�	�U2�K�S���h��n�W�b���H�)�%��� ��»�電�z��n���Bc�0���9��X���j�.m�I�^�@B��Q�&��i��P������0:���:(�:�;��;��;��;�;vz	;%��:�S�:B$L:�չ���qÊ�R�ۻj����>�fX\�>{l��0l���[���=�7r�����H&���ޙ������'��_�!��oE���`���m��Oj���V��6�@���Qɻ�rt�Z<ܺ;����~:(@�:-� ;�G
;\�;
x;*&;6;`3;5>�:o��:D�9'q�85�������|�%� �I�c�X_n��xh�cS�,P2����+ֻ�5��QГ�ݓ���ϻw	��?.��O�W�f��  �  ��U���M�
8��T�%��HP���1��������99��:J��:9|�:��;�3
;9;G�	;O;.��:���:��:a@�7���/XM�K���.�����[�=���P�J�U��+K��3�Ԉ��%�ra��V~���G}�,���nǻ?�&�zB��R���T�B�G�R@.�LE���ͻzj��NX���� :fð:��:�s;x�;Tr;"�;ac	;��;�N�:�L�:S<:<���F6����x���Ļ(�d�*�WE���S�_S��XD�qL)����9�ͻ����~��Ȃ�=����ۻ=��s+0���H�� U��Q�"q@�K�#�8����t���Z[���ź𨾸�l:՞�:q��:je;
<
;��;�P;�;�n ;���:ڟ:���9�{W�׃"��ꓻ�޻�/�:�4��K��|U��P��y<���������B�����z������=���j�X��!�9���N�:�U���M�C�7�t"����^�<M0��>��Z�9�,�:�*�:�$�:�z;�;*�;.
;[;~�:��:�*�:u�"8&q����L�C���l�������=��P�loU�YK��p3�J_���⻹�����z|��Õ� ǻH�|�%���A���R��T��G�m.�$��Hͻ7��� �.o�Wh!:��:���:�~;��;z^;w;21	;>Y;��:���:+]::b�¹O���y��-Ż3���*���E�9T�I�S���D� �)�v��λ�������?��@*��ܻ��[0�(I�/*U��R��@���#� ������[�i'Ǻ�`ո1i:d�:)�:�;[W	;&;�f
;A3;��:���:��:W �9#�Z��]#��X��،޻�i���4�UL���U��VP��<�G��c����㺻N����S{�+K���ش�o �%���9���N��  �  ��1�y{+�n��� ��*Ļz`��;��XS��~�r8Y/Y:켯:���:SZ�:2� ;��;��:R��:�1�:�G�:��2:��!��ī��6������ѻ�F������-��o1�aE(�����e�q����~�G���;��d�P��C�ջ�.�g ���.��0�n�&�Q��c|�p����g�8(��CN"��l�9*v�:aQ�:'�:�x�:d�;
�;VS�:o�:���:�Ϗ:��99 ��͈Z�uS���������$�K;0� �/�_U"���
��ܻ*����Sk�'�<��B�u;|��Ү��o黲���Z&��0�h�.��� �q+	� Iػ� ���YB�����#���#!:�$�:���:�:1��:�m;_	;�?�:�7�:D�:�n:df39
ze����r���鼻IT����&�)�b|1���,�T��Y���LȻ`ȑ��MV���8��uP�%������~���
��/+�ߓ1�D+��������B�ûE ��z��0̄�dj�8vf\:�c�:���:�:w�;�x;�` ;�l�:��:�¤:�|5:[��f���`o6��S��Άѻ�(�br�F�-��N1��!(�����/��f���t�F�^�:�M�c��蜻(}ջ���}7 �7�.�'�0��|&����:컼5���:g�B{��E1!��,�9�Ǉ:���:�;�:!o�:z{;�;$��:���:T�:��:�c�9��^1�	#[�����V������$�+r0�X�/���"��9�S�ܻg#���Jl���=�M�C�o}�4>��-���)�&��1��.�� �SQ	���ػdO��"�B��e������*:i��:x��:Z@�:W��:��;;e�:�b�:�v�:lk:��%9��h��y�,���?Y������mV��*���1���,�o��V���Ȼ5f��3�W���9�;�Q�� ��;`»���M�jn+��  �  ���x��%��9λ�����xq�D !������}���69��<:V�:Di�:eQ�:���:�:q�:�܊:��:�{87�ZsӺ�2�Q,�������ֻ,�����x���e����ݻ!/��m���,����U޺"���W��q��T_ʻ�8�\m�'L����y组\���;���5U���	���iz���9�9��g:⪦:-;�:�l�:���:���:���:�u:7	�9�:���}��#���K�<��;\�����sU ������a\����λ<k����`��q���ߺ���If$���t��j����ػ0��vZ�}�\����ڻ������r":�l��bL� S�? ::0��:_f�:^u�:s�:���:>)�:S3N:�ǅ9`Eݹ��i���Mg�����GSɻP9�S���Z�JO�` �?���;��,�D����BٺdN �h&<��䉻S{������)�
I���������ͻ3�����p��= �����O�B�C9�"@:��:-�:��:��:���:�"�:�|�:@�":qx;8�e4�|8ҺZv1��聻�U��6�ֻ�\��h���I��#Oݻ.ݯ���~��,�(��]�ܺ!O�W������ɻ���@�"����������u��j�T�ř�`"��*���\{�9N�g:��:>1�:�D�:�N�:��:�>�:E�s:��9�fA�K��� �4L��l������w)�� ��m;������]ϻ$埻��a�-e�#��)�뺟E%�Pmu�qϪ��ٻv��q���+����S(ۻg��������:��j�qcO��+'�x�:���:�'�:��:\��:��:L�:�K�:�J:C}9*C么�����~'h��*��h�ɻ���)�����V�껾L��ҏ�^ F��V���ۺ����P=��t�����.��xg��  �  �������P��u��ݥ���Zr��jC�,����Һ��w����Xݚ9a�O:��:���:�Ë:�6:p�09'0����P溇��ĹM�!�|�����1Ū�κ��g»��� |����O^��[������5-����I�w�JH�G�<������c�������6»WP�������P��¯���$b�!�3��T�������<�4���l��9�-u:a8�:��:Q�:��:�̅��(�?-��y� �A.��c\�<Ʌ����v\��W��»{9��ꥻ�	���D��B��ޥ���M�^���D����
�h3U��Ŏ�����?���P»;ٻ�ו��3◻g����FR�"$�g���]H��%�8(,:���:9�:!�:��_:ڱ�9=ke�U/a��JǺz��-s=�?Jl�����ɣ�W⵻�������p괻!���\v��+�d˺��Q��*�D�B������"��,n�Ug���ϲ��F��HF��q���a��yD��Ƙq�k�B�6���%Ѻtwt�w������9��S:�Ĕ:ݐ�:a��:ӣ9:�X>9��Ṱ���l���%��!M��A|��i������ ����&»�u���4���v����]����X��A*����ot�5��n�;��3�����˧��������@R����?w��W�a�93������I�;����X��9�u:2�:�؝:�:��:f����*�����x�Պ.�[�\����t�$����X���y» ���j]������E�p$��c���W��uM#�����~���U��#������d�����»�(��嬻�2������R��$��0�6���,�����8�b(:\��:'�:��:<\:�9gNt���d��ɺ*���L>��"m����t8��mU�����w���m��RE���xw�}6,�;�ͺ��V���
�ЖG�I��I�#�f9o��晻H���  �  �z�L+�� ����9��0&���@��欇�1yx��%V��(�Up溔�o�à8�坥9n�98"u9,���Oݏ�/��5�3�3�^�r�~�����%���Y���Ґ��`������ds��O�h	 ��`ӺkK�����W��9a�9@y-9�&�骡�yd�WN;���d�]-��5���ڑ��,I��O���K���6��=�m�e�G�%��N쿺Y'��58��9X��9���8
�����R��*WB���i��ɂ��]������q���Ǝ����=��*�g���?����K;��#a���9�v�9C�9ѓ�6'{1�%�źÙ���I�6Yo�0���0���O�� ��*;������=K���b�2)8�&���9��E�ʹmS9]��9�¿9u���T�?#غX."���P�/ct��@���R��瓐���֎�����]3|��[��
0�����|����N�����9���9~9�9�jM�kmw�.��̓*�TzW�[2y�6���P���֐��Đ�xߍ��I���w�=RU�:�'�9��V�k�m�)�+<�9O�9"�9qO�����p��W�2��^���}�c0���ێ�&��֏��/���ͅ���r�0�N��q�Һ*�H�צx����9���9��99�߹�,��ߩ�a�:���c��܀�(H���L���
�����s��X���m��cG�C������Y'���8���9���9᭺8�������(�7�B��9j����̨��T���U��3폻�W���}���h�Ms@�"l�3����\�8
>�9��9|�޶��4�Ǻ�T�tsJ�p�`���	Ќ�����%s������[��=���1�b�\9�>�����M�ҹ\{C9Գ�9f��9D�4�W��ں�#���Q��@u�������������_���������'}���\��1��'������b����9���91�9�_�ް{����~�+��eX��  �  aO��F�|�t�푻 ������r���zJ���%��{*��.
k�]��y���?v@�@�&K^�ywԺ�K0�ir{�}ٞ�+a��0���ɶ��Il������Y����Xj�@�;�!�h�ú�yZ�d�L�o��9k�b:�ʗ:;&�:���:":���8F���蜺xp���
'�U5U��.��b?��縭�%����w»��Xj�����+MQ�[��d������	�����D����H�) ���|������7»{���m���b���u����Y�~Q+�����&ۤ���3��7��:��:J��:ٛ:�&q:���9
Z�q�D�%ٸ�0��]�5���d��ډ�`Z���V��$���f���qܷ�����G����7��ຨ]k�r�	�6�/�������Ϳa�^1��\���꾻V����Ź�m\�����bsy��\J��u��ߺ�p��VιI[b9*�@:�Ï:��:[W�:��M:�X�9�@���}���պ�t�;4E�{6t�����0��+P��F����⿻ι�������j����L���`�<��L��bZ�U�Һ�`/��z��p�������Z��~c����6���!x��e�i��;������ºvX�j�B����9��e:�5�:L��:�q�:�q%:��8������y!�!m&�x�T�l끻I��q����d�� O»g��� P�������5Q�V��o�������扺�����H��N�������X���{»sŽ�Ӿ��ǹ���҄�
tZ�� ,��T������ �!�F7h�:?�:ҝ:c�:�m:q�9�����G��<��;	���6�+)e��-��ɯ��$����￻�3»pG�����A���]�8���⺡zo�7����3�p�����b�����6ϯ��Y���X»T0���Ʃ��|��Pz�AK��c��ấu��ifֹQ9�u<:Ћ�:���:�&�:�{I:��9i3��uŀ�x�׺�  �  �˽�8>%��1v�h��pл7���n�Ak�J��,Z�W���Ƈ��9�Bn��a�ۺ7���`J��x��D�»��������%�����wmǻ*����Xc�h�"�����̹���9g,R:EU�:�T�:�h�:���:��:Z��:1��:�Q
:d����_Z��H���>��1��]���
ݻg���V�D%�"����sֻ�ܧ���o�?'!������⺡$�"�e��R����ѻ�:���m����m��H���������G����;p�q9��#�9Qy|:���:��:��:�t�:�A�:�Ԥ:�1b:,ʸ9<���}Β����Y�Y�����»q�軘A��F�m����^�ǻ�`��bzR�\��|ۺ�+���/����(�� ~߻�9 ����������iԻת�
�~�x�,���ʺY�'�4�8t�*:q��:0z�:�0�:��:�T�:ot�:�2�:�_9:�� 9Y������p$��ju�����л�r�?<��6�c��5���޷�J���8��e���ٺx��dI�����Qg»�5����c��]����h"ǻ�c���b�Z���h��33ȹML�9��T:؟�:a��:���:9�:�0�:��:��:~:����W���J>��`\����ܻ����B���1���,aֻOѧ��o�-!�m����V�f��y���ѻ�o����E��ö��g%�%\��"��w�G�߮����s����� �9��x:6�:U��:<��:���:���:m?�:Y)_:���9{��&��Y�>.Z�,ٗ�.�»O!�Er�zz���5����ǻrᗻ0�S��j�M�ݺIJ���0�����������߻�s ��)�E9�����ԻA��L��y�-��X̺8�+�7Ԏ87�&:=��:DX�:;	�:���:4�:�_�:�.�:�5:��9���  �  ����%�b���F�ǻ�����C%,���1�b�*�r��T�����[�����N��:�H�Z����a$̻��6��[-�V�1��?)�� �[y��Fڹ��{�ν��V���[9y�t:���:߅�:���:��;d�;��:���:�f�:3��:[�:y����ȺR�H�B~����ۻ�
�4�!��E/���0�d|%�����I�?m9x��RA��K>���o��ѥ� �߻ɑ�>q#�-�/��/�c�#�}�:1��줻4BT��ۺh߹�:A�:ˑ�:x�:���:`P;��;n8�:�4�:qW�:S��:�p�9��1�3�H�m�w�����((�i'��1�1>.����w��6һ���E`���9�
�H����N4���K�7��(�g1�q+-��@�;��5λ�搻~X0�B���	"��@:P�:��:_��:�� ;��;�^;�-�:,��:ϊ�:�WS:���7b獺H�$��H��\5ǻ*v�J��P�+�t�1��{*��������,���6	����M�r�8��Y�������˻-Y����s'-��l1��)����,�����j�z�
2��rT���d9�v:��:���:,�:�>;Bc;���:.��:��:$ �:Y: s��Q~Ǻ�%H�0=���ۻ��
��!��1/�<�0��o%�\��Z>�꫻r?x�9gA��n>��o�����߻Ѩ�Ë#�!0�^0���#��������G���U�]ݺ���f�9�W�:���:Q��:y�:t;W�;]��:��:ֽ:ȅ�:q�9��4�����]n��
��a��3W��'�M1��v.� \�O���һL����[a��;�C�I�뛅��������dS��&)���1��a-��u�`���oλ9Q���21�	l���ԸF<:JU�:��:���:��:.�;IU ;<&�:G��:��:��O:��6�  �  �č�Y8��X���"뻬E�֋9�
�N���U�k�M�!S8�C�?B��䱻B����{�hi����!?��� � %>�>Q���U�K�^N3�/d��Eڻ�N���s�4XE����9��:=��:/\ ;i�;ƽ
;�?;�p	;�f;��:f/�:��^:��+�UvҺ�c�8���V���n%�=�A�"�R�H�T�&�G��.���?ػqf�����@C�������<ѻ��	�u+���E�o�S�uS�/D���(���������Lq�K{麻N���I:n��:6��:];�	;Q�;[�;x�;�7;���:} �:��:�K�����(����ѻ6���/���H�p�T�:
R��@��$�7'���û}�����{�iX��C���:`�p<���4���K���U���O��E<����"%���UoE�ח����8�:q��:���:H�;W�
;p;	;xD;m��:A~�:�N�:[�n9�#���B7�%���t��3�VZ9��kN�%�U��M��8������>_��0��zz�bᏻ�n������=q �u�=��P��`U�*�J��#3��<�,�ٻ������� C�z.�9�>�:��:7� ;U[;�j;3�;�"
;�;�W�:��:D1a:��!�EKѺzb��s��)���T%�b�A��}R�&�T�z�G���.�n���:ػ�i��T���T��)����\ѻL�	�g5+��E�>T�7�S�sSD�I
)�%����r�B�"͞�R-F:�߻:
 �:�~;�	;Z;P�
;�#;/p;p�:�:G4:� ��B�c~��.�ѻ�c��0���H��#U�%DR���@�mN$��j��PĻ�B����|�K冻k;��O���|�K;5��-L�
�U��(P�{z<�r����}��SFF��T���8	�:���:���:Ǖ;2�	;[;�
;�E;���:��:���:�
a9�  �  `k���ML�O������,���N�of�v�n�N�e�(N�F1,�e��wj̻�ߠ��> ���ٻq&��K4�ˇT�_5i��-n��ob��H�+H#��E󻇔��n�-��MY�B2:��:'�:��;u�;�q;n�;e�;�?
;�T ;�R�:�Ss:J�:�~��&Z|���ͻ��َ8��-X���j�iYm�?O_�߀C���C������Ө���N���xb�ʹ?��\��}l���k�h�Z��m<�Rp���ֻ92�� \��C��O\:�{�:���:�d
;�Q;�v;LN;q�;��;/�: `�:p_":�)�6"�����~�黯��-D�#�_��ym�Q[j�BW�H 8�_�*�߻ܼ������B����Ż��x�'��J��c�|,n��g�K	R��,0����1��[[��³�J��8+�:v��:%;�;\�;v;��;��;u_;���:���:�ȃ9�͚�'�K������B�+�A�N��;f��Rn���e�:�M�q�+���R�˻V���d��c�����ػ;���4�AMT���h��m�EAb���G�& #�5��L��'�,��W��v:0�:�]�:�;>F;!;Jd;�i;N�
;�;>��:��u:�0�����{�5�ͻ���t8��X�&�j�aIm��B_��wC�p��<�����P���G����g��f���u���?�;�\���l���k���Z�/�<�����׻#����"�����0�X:U��:�
�:�	;:v;t�;�z;��;�;��:�:��:
�,�����ח���黙���]D��+`��m���j�Y�W��A8��G��g��K�����hН�pFƻ���m(��J�'�c��dn�'%h��=R�`0�]��Й���/\�nz����8-	�: �:�;�;��;@r;��;��;�j;s�:&7�:�z9�  �  \Y��9�T�?������2��V�/�n�}Iw�Un�c�U���2����ջ
�����~��":㻐���:;��r\���q���v�r�j�,�O��w)����������4���e�J' :sd�:���:]{;��;�j;\�;q�;G�;S ;�p�:��u:ǞU���N��V�ջH��?��5`��{s�yv���g���J��%��N �	qû�|���������.����!��G�@�d�X.u���t�o�b��C�o"��߻ܡ��1�q���]:�z�:�;�;�n;�f;zC;�;�
;���:q�:�B": �4���$�,�������$���K�CCh��4v�*�r�DD_�9?����v��8��ԛ�TX���λ>6��b.��$R��l���v�H}p���Y���6������»qod�ѓ��qz�8J��:a1�:f�;`;�;�`;��;x�;?�;�>�:��:{9󼢺DT�*'��t���d2�fV���n�vw�-n�[�U���2�
V��?ջ����H7��f���{��	��'�:��7\��q�ӹv���j��TO�_O)��X��V���;\4�0�c�@l:���:���:?	;H{;�;�Q;n;T;��;���:�'x:��K�jl�	��ʈջfb�f?�`��hs�{ v��g���J���%��L �+tû놠�����$������i�!��G��e�
Lu���t��c�)�C��L��l߻� ��c��Pό�Z:	��:/5 ;��
;��;��;3p;�;�X	;��:���:*{:��7�\�%��睻e����$�7�K��vh�lv�4s�Ă_�O?�u;��S껏Ǵ�#d��"祻�wϻz���.��bR��Ol�R$w�b�p�EZ�?7�7���»�Ce��I����8Sϒ:I�:]�;`;_�;D^;��;��;�;Ai�:�C�:��m9�  �  `k���ML�O������,���N�of�v�n�N�e�(N�F1,�e��wj̻�ߠ��> ���ٻq&��K4�ˇT�_5i��-n��ob��H�+H#��E󻇔��n�-��MY�B2:��:'�:��;u�;�q;n�;e�;�?
;�T ;�R�:�Ss:J�:�~��&Z|���ͻ��َ8��-X���j�iYm�?O_�߀C���C������Ө���N���xb�ʹ?��\��}l���k�h�Z��m<�Rp���ֻ92�� \��C��O\:�{�:���:�d
;�Q;�v;LN;q�;��;/�: `�:p_":�)�6"�����~�黯��-D�#�_��ym�Q[j�BW�H 8�_�*�߻ܼ������B����Ż��x�'��J��c�|,n��g�K	R��,0����1��[[��³�J��8+�:v��:%;�;\�;v;��;��;u_;���:���:�ȃ9�͚�'�K������B�+�A�N��;f��Rn���e�:�M�q�+���R�˻V���d��c�����ػ;���4�AMT���h��m�EAb���G�& #�5��L��'�,��W��v:0�:�]�:�;>F;!;Jd;�i;N�
;�;>��:��u:�0�����{�5�ͻ���t8��X�&�j�aIm��B_��wC�p��<�����P���G����g��f���u���?�;�\���l���k���Z�/�<�����׻#����"�����0�X:U��:�
�:�	;:v;t�;�z;��;�;��:�:��:
�,�����ח���黙���]D��+`��m���j�Y�W��A8��G��g��K�����hН�pFƻ���m(��J�'�c��dn�'%h��=R�`0�]��Й���/\�nz����8-	�: �:�;�;��;@r;��;��;�j;s�:&7�:�z9�  �  �č�Y8��X���"뻬E�֋9�
�N���U�k�M�!S8�C�?B��䱻B����{�hi����!?��� � %>�>Q���U�K�^N3�/d��Eڻ�N���s�4XE����9��:=��:/\ ;i�;ƽ
;�?;�p	;�f;��:f/�:��^:��+�UvҺ�c�8���V���n%�=�A�"�R�H�T�&�G��.���?ػqf�����@C�������<ѻ��	�u+���E�o�S�uS�/D���(���������Lq�K{麻N���I:n��:6��:];�	;Q�;[�;x�;�7;���:} �:��:�K�����(����ѻ6���/���H�p�T�:
R��@��$�7'���û}�����{�iX��C���:`�p<���4���K���U���O��E<����"%���UoE�ח����8�:q��:���:H�;W�
;p;	;xD;m��:A~�:�N�:[�n9�#���B7�%���t��3�VZ9��kN�%�U��M��8������>_��0��zz�bᏻ�n������=q �u�=��P��`U�*�J��#3��<�,�ٻ������� C�z.�9�>�:��:7� ;U[;�j;3�;�"
;�;�W�:��:D1a:��!�EKѺzb��s��)���T%�b�A��}R�&�T�z�G���.�n���:ػ�i��T���T��)����\ѻL�	�g5+��E�>T�7�S�sSD�I
)�%����r�B�"͞�R-F:�߻:
 �:�~;�	;Z;P�
;�#;/p;p�:�:G4:� ��B�c~��.�ѻ�c��0���H��#U�%DR���@�mN$��j��PĻ�B����|�K冻k;��O���|�K;5��-L�
�U��(P�{z<�r����}��SFF��T���8	�:���:���:Ǖ;2�	;[;�
;�E;���:��:���:�
a9�  �  ����%�b���F�ǻ�����C%,���1�b�*�r��T�����[�����N��:�H�Z����a$̻��6��[-�V�1��?)�� �[y��Fڹ��{�ν��V���[9y�t:���:߅�:���:��;d�;��:���:�f�:3��:[�:y����ȺR�H�B~����ۻ�
�4�!��E/���0�d|%�����I�?m9x��RA��K>���o��ѥ� �߻ɑ�>q#�-�/��/�c�#�}�:1��줻4BT��ۺh߹�:A�:ˑ�:x�:���:`P;��;n8�:�4�:qW�:S��:�p�9��1�3�H�m�w�����((�i'��1�1>.����w��6һ���E`���9�
�H����N4���K�7��(�g1�q+-��@�;��5λ�搻~X0�B���	"��@:P�:��:_��:�� ;��;�^;�-�:,��:ϊ�:�WS:���7b獺H�$��H��\5ǻ*v�J��P�+�t�1��{*��������,���6	����M�r�8��Y�������˻-Y����s'-��l1��)����,�����j�z�
2��rT���d9�v:��:���:,�:�>;Bc;���:.��:��:$ �:Y: s��Q~Ǻ�%H�0=���ۻ��
��!��1/�<�0��o%�\��Z>�꫻r?x�9gA��n>��o�����߻Ѩ�Ë#�!0�^0���#��������G���U�]ݺ���f�9�W�:���:Q��:y�:t;W�;]��:��:ֽ:ȅ�:q�9��4�����]n��
��a��3W��'�M1��v.� \�O���һL����[a��;�C�I�뛅��������dS��&)���1��a-��u�`���oλ9Q���21�	l���ԸF<:JU�:��:���:��:.�;IU ;<&�:G��:��:��O:��6�  �  �˽�8>%��1v�h��pл7���n�Ak�J��,Z�W���Ƈ��9�Bn��a�ۺ7���`J��x��D�»��������%�����wmǻ*����Xc�h�"�����̹���9g,R:EU�:�T�:�h�:���:��:Z��:1��:�Q
:d����_Z��H���>��1��]���
ݻg���V�D%�"����sֻ�ܧ���o�?'!������⺡$�"�e��R����ѻ�:���m����m��H���������G����;p�q9��#�9Qy|:���:��:��:�t�:�A�:�Ԥ:�1b:,ʸ9<���}Β����Y�Y�����»q�軘A��F�m����^�ǻ�`��bzR�\��|ۺ�+���/����(�� ~߻�9 ����������iԻת�
�~�x�,���ʺY�'�4�8t�*:q��:0z�:�0�:��:�T�:ot�:�2�:�_9:�� 9Y������p$��ju�����л�r�?<��6�c��5���޷�J���8��e���ٺx��dI�����Qg»�5����c��]����h"ǻ�c���b�Z���h��33ȹML�9��T:؟�:a��:���:9�:�0�:��:��:~:����W���J>��`\����ܻ����B���1���,aֻOѧ��o�-!�m����V�f��y���ѻ�o����E��ö��g%�%\��"��w�G�߮����s����� �9��x:6�:U��:<��:���:���:m?�:Y)_:���9{��&��Y�>.Z�,ٗ�.�»O!�Er�zz���5����ǻrᗻ0�S��j�M�ݺIJ���0�����������߻�s ��)�E9�����ԻA��L��y�-��X̺8�+�7Ԏ87�&:=��:DX�:;	�:���:4�:�_�:�.�:�5:��9���  �  aO��F�|�t�푻 ������r���zJ���%��{*��.
k�]��y���?v@�@�&K^�ywԺ�K0�ir{�}ٞ�+a��0���ɶ��Il������Y����Xj�@�;�!�h�ú�yZ�d�L�o��9k�b:�ʗ:;&�:���:":���8F���蜺xp���
'�U5U��.��b?��縭�%����w»��Xj�����+MQ�[��d������	�����D����H�) ���|������7»{���m���b���u����Y�~Q+�����&ۤ���3��7��:��:J��:ٛ:�&q:���9
Z�q�D�%ٸ�0��]�5���d��ډ�`Z���V��$���f���qܷ�����G����7��ຨ]k�r�	�6�/�������Ϳa�^1��\���꾻V����Ź�m\�����bsy��\J��u��ߺ�p��VιI[b9*�@:�Ï:��:[W�:��M:�X�9�@���}���պ�t�;4E�{6t�����0��+P��F����⿻ι�������j����L���`�<��L��bZ�U�Һ�`/��z��p�������Z��~c����6���!x��e�i��;������ºvX�j�B����9��e:�5�:L��:�q�:�q%:��8������y!�!m&�x�T�l끻I��q����d�� O»g��� P�������5Q�V��o�������扺�����H��N�������X���{»sŽ�Ӿ��ǹ���҄�
tZ�� ,��T������ �!�F7h�:?�:ҝ:c�:�m:q�9�����G��<��;	���6�+)e��-��ɯ��$����￻�3»pG�����A���]�8���⺡zo�7����3�p�����b�����6ϯ��Y���X»T0���Ʃ��|��Pz�AK��c��ấu��ifֹQ9�u<:Ћ�:���:�&�:�{I:��9i3��uŀ�x�׺�  �  �z�L+�� ����9��0&���@��欇�1yx��%V��(�Up溔�o�à8�坥9n�98"u9,���Oݏ�/��5�3�3�^�r�~�����%���Y���Ґ��`������ds��O�h	 ��`ӺkK�����W��9a�9@y-9�&�骡�yd�WN;���d�]-��5���ڑ��,I��O���K���6��=�m�e�G�%��N쿺Y'��58��9X��9���8
�����R��*WB���i��ɂ��]������q���Ǝ����=��*�g���?����K;��#a���9�v�9C�9ѓ�6'{1�%�źÙ���I�6Yo�0���0���O�� ��*;������=K���b�2)8�&���9��E�ʹmS9]��9�¿9u���T�?#غX."���P�/ct��@���R��瓐���֎�����]3|��[��
0�����|����N�����9���9~9�9�jM�kmw�.��̓*�TzW�[2y�6���P���֐��Đ�xߍ��I���w�=RU�:�'�9��V�k�m�)�+<�9O�9"�9qO�����p��W�2��^���}�c0���ێ�&��֏��/���ͅ���r�0�N��q�Һ*�H�צx����9���9��99�߹�,��ߩ�a�:���c��܀�(H���L���
�����s��X���m��cG�C������Y'���8���9���9᭺8�������(�7�B��9j����̨��T���U��3폻�W���}���h�Ms@�"l�3����\�8
>�9��9|�޶��4�Ǻ�T�tsJ�p�`���	Ќ�����%s������[��=���1�b�\9�>�����M�ҹ\{C9Գ�9f��9D�4�W��ں�#���Q��@u�������������_���������'}���\��1��'������b����9���91�9�_�ް{����~�+��eX��  �  �������P��u��ݥ���Zr��jC�,����Һ��w����Xݚ9a�O:��:���:�Ë:�6:p�09'0����P溇��ĹM�!�|�����1Ū�κ��g»��� |����O^��[������5-����I�w�JH�G�<������c�������6»WP�������P��¯���$b�!�3��T�������<�4���l��9�-u:a8�:��:Q�:��:�̅��(�?-��y� �A.��c\�<Ʌ����v\��W��»{9��ꥻ�	���D��B��ޥ���M�^���D����
�h3U��Ŏ�����?���P»;ٻ�ו��3◻g����FR�"$�g���]H��%�8(,:���:9�:!�:��_:ڱ�9=ke�U/a��JǺz��-s=�?Jl�����ɣ�W⵻�������p괻!���\v��+�d˺��Q��*�D�B������"��,n�Ug���ϲ��F��HF��q���a��yD��Ƙq�k�B�6���%Ѻtwt�w������9��S:�Ĕ:ݐ�:a��:ӣ9:�X>9��Ṱ���l���%��!M��A|��i������ ����&»�u���4���v����]����X��A*����ot�5��n�;��3�����˧��������@R����?w��W�a�93������I�;����X��9�u:2�:�؝:�:��:f����*�����x�Պ.�[�\����t�$����X���y» ���j]������E�p$��c���W��uM#�����~���U��#������d�����»�(��嬻�2������R��$��0�6���,�����8�b(:\��:'�:��:<\:�9gNt���d��ɺ*���L>��"m����t8��mU�����w���m��RE���xw�}6,�;�ͺ��V���
�ЖG�I��I�#�f9o��晻H���  �  ���x��%��9λ�����xq�D !������}���69��<:V�:Di�:eQ�:���:�:q�:�܊:��:�{87�ZsӺ�2�Q,�������ֻ,�����x���e����ݻ!/��m���,����U޺"���W��q��T_ʻ�8�\m�'L����y组\���;���5U���	���iz���9�9��g:⪦:-;�:�l�:���:���:���:�u:7	�9�:���}��#���K�<��;\�����sU ������a\����λ<k����`��q���ߺ���If$���t��j����ػ0��vZ�}�\����ڻ������r":�l��bL� S�? ::0��:_f�:^u�:s�:���:>)�:S3N:�ǅ9`Eݹ��i���Mg�����GSɻP9�S���Z�JO�` �?���;��,�D����BٺdN �h&<��䉻S{������)�
I���������ͻ3�����p��= �����O�B�C9�"@:��:-�:��:��:���:�"�:�|�:@�":qx;8�e4�|8ҺZv1��聻�U��6�ֻ�\��h���I��#Oݻ.ݯ���~��,�(��]�ܺ!O�W������ɻ���@�"����������u��j�T�ř�`"��*���\{�9N�g:��:>1�:�D�:�N�:��:�>�:E�s:��9�fA�K��� �4L��l������w)�� ��m;������]ϻ$埻��a�-e�#��)�뺟E%�Pmu�qϪ��ٻv��q���+����S(ۻg��������:��j�qcO��+'�x�:���:�'�:��:\��:��:L�:�K�:�J:C}9*C么�����~'h��*��h�ɻ���)�����V�껾L��ҏ�^ F��V���ۺ����P=��t�����.��xg��  �  ��1�y{+�n��� ��*Ļz`��;��XS��~�r8Y/Y:켯:���:SZ�:2� ;��;��:R��:�1�:�G�:��2:��!��ī��6������ѻ�F������-��o1�aE(�����e�q����~�G���;��d�P��C�ջ�.�g ���.��0�n�&�Q��c|�p����g�8(��CN"��l�9*v�:aQ�:'�:�x�:d�;
�;VS�:o�:���:�Ϗ:��99 ��͈Z�uS���������$�K;0� �/�_U"���
��ܻ*����Sk�'�<��B�u;|��Ү��o黲���Z&��0�h�.��� �q+	� Iػ� ���YB�����#���#!:�$�:���:�:1��:�m;_	;�?�:�7�:D�:�n:df39
ze����r���鼻IT����&�)�b|1���,�T��Y���LȻ`ȑ��MV���8��uP�%������~���
��/+�ߓ1�D+��������B�ûE ��z��0̄�dj�8vf\:�c�:���:�:w�;�x;�` ;�l�:��:�¤:�|5:[��f���`o6��S��Άѻ�(�br�F�-��N1��!(�����/��f���t�F�^�:�M�c��蜻(}ջ���}7 �7�.�'�0��|&����:컼5���:g�B{��E1!��,�9�Ǉ:���:�;�:!o�:z{;�;$��:���:T�:��:�c�9��^1�	#[�����V������$�+r0�X�/���"��9�S�ܻg#���Jl���=�M�C�o}�4>��-���)�&��1��.�� �SQ	���ػdO��"�B��e������*:i��:x��:Z@�:W��:��;;e�:�b�:�v�:lk:��%9��h��y�,���?Y������mV��*���1���,�o��V���Ȼ5f��3�W���9�;�Q�� ��;`»���M�jn+��  �  ��U���M�
8��T�%��HP���1��������99��:J��:9|�:��;�3
;9;G�	;O;.��:���:��:a@�7���/XM�K���.�����[�=���P�J�U��+K��3�Ԉ��%�ra��V~���G}�,���nǻ?�&�zB��R���T�B�G�R@.�LE���ͻzj��NX���� :fð:��:�s;x�;Tr;"�;ac	;��;�N�:�L�:S<:<���F6����x���Ļ(�d�*�WE���S�_S��XD�qL)����9�ͻ����~��Ȃ�=����ۻ=��s+0���H�� U��Q�"q@�K�#�8����t���Z[���ź𨾸�l:՞�:q��:je;
<
;��;�P;�;�n ;���:ڟ:���9�{W�׃"��ꓻ�޻�/�:�4��K��|U��P��y<���������B�����z������=���j�X��!�9���N�:�U���M�C�7�t"����^�<M0��>��Z�9�,�:�*�:�$�:�z;�;*�;.
;[;~�:��:�*�:u�"8&q����L�C���l�������=��P�loU�YK��p3�J_���⻹�����z|��Õ� ǻH�|�%���A���R��T��G�m.�$��Hͻ7��� �.o�Wh!:��:���:�~;��;z^;w;21	;>Y;��:���:+]::b�¹O���y��-Ż3���*���E�9T�I�S���D� �)�v��λ�������?��@*��ܻ��[0�(I�/*U��R��@���#� ������[�i'Ǻ�`ո1i:d�:)�:�;[W	;&;�f
;A3;��:���:��:W �9#�Z��]#��X��،޻�i���4�UL���U��VP��<�G��c����㺻N����S{�+K���ش�o �%���9���N��  �  n�n���e��KM���)�e� �K���=D�#4��wk�9ė�:���:�;E�;�;g�;��;'�
;�m;��:�r�:!%8 ºd�����
�r2���S�:�h�N2n���b�]�H���%��� �{1û�M��┻�`�����zG��!:�/�X�bk�Hm���^�EeB�}s���%O��@$�_
�g0:�4�:���:X�;I�;�;� ;[�;�	;OS�:�:��M:��ѹo��u��^ۻ<��$]>��#\��Cl�R�k�Z[��=�C3���Y�����f��������R�!�.@E�Zm`�d�m�`(j��V��x6�4���ɻ��s���ں�_θT̀:���:T�;j#;p;�];�;R;�;��:6g�:���9y�m�A^4�����\���AO%�T�I��Hc�n�2h�;�R�2�<��:�ջ�����,����ϻ����-��O�c�f��Ln�iKe��M�"�)��� �������C�)���U��9F)�:��:R�;��;�;V;J�;��;�-;m�:�Ì:�:8@�����c��ۿ�6�	�U2�K�S���h��n�W�b���H�)�%��� ��»�電�z��n���Bc�0���9��X���j�.m�I�^�@B��Q�&��i��P������0:���:(�:�;��;��;��;�;vz	;%��:�S�:B$L:�չ���qÊ�R�ۻj����>�fX\�>{l��0l���[���=�7r�����H&���ޙ������'��_�!��oE���`���m��Oj���V��6�@���Qɻ�rt�Z<ܺ;����~:(@�:-� ;�G
;\�;
x;*&;6;`3;5>�:o��:D�9'q�85�������|�%� �I�c�X_n��xh�cS�,P2����+ֻ�5��QГ�ݓ���ϻw	��?.��O�W�f��  �  �������F�:)��M��e���R�o� �5����һ&������j�����t���q�ƨv�������� ���?޻����A���~��٢���ȼ+���$��k�N��{��-- �ܛ��.��A���#S������Y���9Ӽ�P��-�9L�
W�
�"����1ټA���D����	[��7%��������T��������4{��3r�b�q��y��ˆ��|��!���� ����HT�򊊼|E��ռ�o��:��������S�o���g�ּ���*O���s�����e�$����ݼx#����
��q����s�ke��̼��ϙG��A��c�\���-��Mރ�#�v��q��+s�7|~�/��S����̻���E�/���h�x�������#ἠ� ���ܶ������LB�§˼x��������W���閼�۪�HȼX�輵��G�W������9�V��5��
�����o��5�i���ѻ&���
���F��N�s���p��u�����Z���&`��L�ݻ۟��vA��f~��ˢ�W�ȼ"��4��d����؍��# �~��m��w��d8���鐼h=��Qֳ���Ҽ�4�m ��?�!K�
�����ټ>���\z��c�Z��$%����ƃ��+����|���8{��Gr���q�E�y��톻צ��K����Z�� ��mT�����\���ռ+���X���������c�����=�ּ�#���p������_<�����aŽ�/�ݼy;��|�
��{��
��|��v���̼������+�G�Bm���以�G|��5M���w���q��t��f�{��Hm���q̻����&0���h�򓖼���[A�� ��R���0��Lk�>�˼�譼����m�����\��T=ȼ<��s,�-X��  �  ��fV	�����߼F9��)㗼��l���4�6V	��tԻL��䎑�;o����y�W@v���{�х����<����V����-*@���z��П��Tļ�����n�
����H �������ۼ�l�������ΐ�T���Ǜ�����f�ͼ�,������������b����<Լ��r7���X���$�9���FĻ`����|��m5����v��Hv���~��������P��ʷ�.��a4R��]��5ʫ�\6мtj�h�M:�L�R��JT�:/Ѽ|���6������A������T����Tؼҷ��� �����T������Nȼ�ã������E��8�WS��p���+��	���n�{�7�u��w�����
��7{λG�X/�k�e�4ߓ�x���ۼ����n�����\
� ��P�ÛƼ\���$┼v�Q������\"ü*�����h�	�K�IH	�o���?�߼f!���˗��l�=�4��%	��Իך���$�����x��gu���z��j��w����R��+�Ⱥ��@���z�y�pGļ{�(��P�
�$���������p�ۼ�U��cw�������}��]��fq���ͼO�H��O�������U����*Լ�௼�)����X�6�$�����Z0ĻB����v��w7����v��lv���~�%߉�����.������J���YR�Nr���ૼ�Nмۄ��v�1I�������u��PѼX���ã��S$��߿��� ������nؼ��������^���԰�Y_ȼ�գ����SF�hd�����ն�e����*����|��lv�9�x��d��B����|��>�λFN��L/��f������'��mܼ� ��L���o
�3��y��Ƽ����������|��dߦ�?Jü��^���״	��  �  ���Ά���!��
ѼO@��-Ɛ� �e�@3�e��2�ݻ�����9���֌�焻�͂�M!�������u��/��K��;�=��Rr�ܗ������׼��� �_n�����c�O�˼��l6���͆�hۃ�����m���⾼|�ۼ��+�*,�w������>�ƼD��xU��Z�S���$��� � hλ󴫻̕�`#��Z>���킻�"��<铻U���Ŧɻ���V ���M��Ⴜk����ü�༾��w��>�������޼V¼�Υ�ɶ���:������ړ�Lī�a�ȼ̓�;���4�<�<S�¹ڼ�
���a���x�3�B�r��_����������h���r��-����+��v������pػ��s.�i_��,��g���s�ͼS_�$���z�r ��sռ�J��.���ъ��=������d���GҼ���������j��e�"�мq(������;�e�a3�X���`ݻ򋵻�͛��h��=x���_��7����!�����������Zq��f=��2r�s͗��q���׼�́ ��f�����SP��˼�֮�w������쿃��ݍ�����ƾ��ۼ���4�i ��r�����\�Ƽ74���G����S���$��� �Rλ����ƕ�w%��rH�������<��B��Uè���ɻ2��T9 ���M�v���㢢�T3ü[�༻���A�����%����޼�&¼�؏�I[��iՅ�����Rૼd�ȼ���-���)>���e�6�ڼ]��t����x���B�'�����`��!������܆��邻�g��������
{��/�ػW��Q.�<�_��G��e�����ͼ�}鼁��K��� ��>�L�ռ�t��쮝����"h��SE�����?��?mҼ���y����  �  h�hἯ�Ҽ����¢��G����_��5�����pͻ7���͟��N���[��U���.���\����Իy��0��H.>���i����������O�ּng㼊���ݼ#�˼,��kΚ�|E����o���j��0|�o|��%���{����ּ�������jݼ��˼�8���͙��w�ˇP��@)�i6
�j[�{�»�Ū�� ��� ��԰��}ҙ�����G���t�໡(��K%�a�K�.�y�r�3E���gɼ%�ۼbY�)O�l�ؼVļk��rؒ��0��0k�z�m�q4��
��_%��}sɼjܼu��V)�Qkؼ	}ļ"����쐼Bo�~B�&����)�ػ;���g���������"��D˝�5��AsɻT|�-X�/1�=EZ�:R��J���lȹ��^м��ZC�=���ҼeU����K����.v��vi�9�s� `��*��_���I~мXc�VJ�bLἶ�Ҽk������n0���V_��\5�9���f�ͻ򯱻�\���ܔ�Oꑻ����l¢������Իû���p��	>���i�{������7���I�ּ�X㼲�弒�ݼ��˼���x����,���o�m[j�f�{��`����������,�ּ�㼯��_Uݼb�˼�&�����v\��pP�~-)�t'
��E廮�»����%#��+����|왻����!ѿ�; �{E�`l%�%�K���y��ؖ�b]����ɼ��ۼ�v��m�'�ؼ�vļ"�������ur��pk�~n��Q���%��6?��X�ɼ`2ܼ¡�W<�{}ؼ�ļ0�������4o�ΨB�<'�}����ػ�)������������������D�������ɻ;��ď��e1�U{Z�im��͟�$幼�|мT8�e������Ҽ�|�����#ɋ�{�v�>�i�Dt�R����P�� �����м`���  �  �üަ���ƶ�y��k9��EY��a��:A�'�%���������H׻ڟ����������o^��*Ļ�ݻ����ѐ��+���G�Z�h�}~���e���3���������ɀ¼mͺ�ɼ��_◼� ���sb��KL�)H�_�V���t�B{��5L���䴼���i(ü�����I����َ��Wx���U�?7������"뻁)λsS�������U��Ņ���X˻[o绡y���5M4�]R��0t�橌��p���[��U��¼����_`��5[��ƴ����x��Y��H�c�J��_������r��џ��b��t���G¼�������g��C���cl��,K��X.�����:�,�໎!ƻOI���g���u���
����ӻ�l�[2��"�o�=�o]�C1��A��Eq���1���ǿ�� ü�,���Y��ö��������l�ޜQ��G�ԋO��0i��h��em��O������z�¼��������`���!���A��c�`��	A�b�%�����P�� �ֻ�+��@��#9���겻�û:ݻSZ��Wb��n+���G�D�h�hn���V��b%��0r�������p¼��������z͗��邼fCb��L�2�G�EeV�b�t�L`���1��+˴�����ü����	���y���ʎ��<x�ѺU��l7�b�������#λ�U�����g�������z˻��b�����m4��?R��Xt���������]u���	����¼�������<{��CՐ�*y�LY�M�H�p�J�.<_�#π�}�������x���¼ZZ¼�ƺ�6���z������w�l�YK��.�^��q����Йƻ�Ĵ��䬻`�$����AԻ���l�""#�2�=�pH]�AL��� ������<O���濼jAü�O��[~��"ݞ�v݉��7m�"�Q��mG���O�ni�����#���祯�
>���  �  Ū��̱��ٝ�s�����ڷ���ip�;D[���E�BT0����q����%ڻDԻR�ݻc(��Б�����#5��J���_�Bu����3���N��4��a桼����ޗ�O���<v�$FU�o9�m(���$�8-0���G��Wg��>�����ޜ�v����ڠ������h��i����U~�"Bi��T���>�� )�
��q�0,�ֻ�ջ��㻠��u��j�&�<���Q���f���{��[��I��%Ě�e_�����t��������ⅼ��j���J��2�#%��&�۲6���Q��Ur�Y[��/���p ��Hڡ������"���7��/��0Gw�9)b���L��W7���!�ru����)߻[�ӻ�1ػ�o��4�����-� PC���X���m��t��5ʋ��_�����Fa���2�������M���/�_�яA��;,�m$�c�*��>�)\�dp}�3��"���.������������Z���錼����9p�g[�ݷE��0�/���6�He�ٻʈӻ�ݻ����Y��}���4���J���_��t�����#���?��!����֡������̗�A��sv��U��?9���'�=�$�~�/�˴G�y#g�%��E���wƜ�W{��GƠ�ʔ���W��Z����;~��+i� �S�A�>�h�(�h��n��.�Rֻ�.ջ`��F@��,���&��:<� �Q��f��|�^q���`��vݚ�Pz��l������������k��"K��G2�a%��	'�%�6���Q�Y�r��r��0������������5��OK��w1��crw��Wb�M�m�7�"��������9�߻�OԻX�ػ���Ms�:����-�ȈC���X��n�l���7勼�{���.�����~�����ݏ�n���`���A�8�,��V$���*�
�>�7r\�׵}��S������  �  �|���숼����4I��/@�� ߋ�����h�� �u��_�0qF�.�,�;���xd��� l�n2�d7L�k�d�Ƽy�m��������N��6[��#��{w���ꇼ*ぼ|1r�'�[��B�	�(�v��%�e��h ����Ւ6� oP���h�Ğ|�k���c#������q\��=猼�����������n��bW���=��$�n�:���;�H_�S"��:���T��0l��B��h����������I�������f�����>H~�%�j�S��-9��� ��s�P��������&�b�>���X���o�#���bO��n��x�Q���k��牼�+��؇{��Hg�t�N���4��v�,3�ZV��g�����)��NC���\�v#s��5�����܄��`���>�����_D������|x� jc��J�V�0��&
���"��o���.��G�"�`�fv�a��T҈��䋼1��n(��Bǋ�=���	���Wu�}_��6F�U�,����Qm��$�l�
��.�32���K���d�H�y��}��߀���<��vJ��0���g���ڇ��ҁ�,r�/v[���A�?�(������~� ��O���_6�==P��|h��p|��w��`��Yy���K��،����|���ۘn�gXW��=�h�$���`���D�+l��c"���:�-�T��Ll��b��z��ת��>ǌ��`��嵌�v����0��e�~�D$k��ES�l9��=!�}����X��%�G&��.?���X���o����Oc���/�����e��%�������D��+�{���g�O�]<5����u�}��n��f�J>*���C�Y]��\s�KQ��l2��b����,���Y���8���a���;��ٽx���c���J�s1��R��r
��[��>	��%��L.�c�G��a���v��  �  �s\�w�q��L��
���2햼�*���š��q������������{��Z���=��)*�hd$�[e-�JXC���a�U�������ړ���6���[��NМ�8����P��3�����l���W��IB�Ю,�����i��g�1�׻mgԻ�~�o��<��'#�r�8��/N�hnc���x�����Ȑ�v����ɟ��ܡ�մ��$��<���Čp��P�@�5��l&���%�*>3�&�L��l��̆�!�������񹡼>.���]��BÑ��Ǉ��z���e�-WP���:��I%����"���F�ӍԻ�UֻK绒M�"!�� *���?��-U�^`j�'r�
��㓼V��������e��o`��'񑼓E���Pe�:&F���.��e$��(�$�:���V�T�w�oҋ�[���ٟ��ȡ�󬞼Aė������\���s�U�^�HI��3��G��C
�� �^ܻ.eӻ3fڻ��ﻃ4�o���L1���F�}=\��cq�[4��x��{Ֆ����ˬ��
X��|v��Hm��|�{�dZ��G=���)��!$�U#-��C��a�#z��w~���z������F��E����攼�?���䀼�l���W�h&B���,��g��>���3�׻pԻ��I�������"��}8�N�lDc��_x����V����������ҡ�����*���)���p�p�m P���5��q&���%�K3�ѱL���l��؆�$�������ˡ��A��s��6ڑ�=�����z�]�e�>�P�w;��%����~���O�⻿ջ��ֻ���-���R��O*���?��WU��j���61������[��|��I���{��l���d��ّe��iF��A/�m�$��(���:��W��&x������w��I���z㡼;Ǟ�mޗ�:���
x��
�s�!�^��I��3����;�
���7�ܻ��ӻ��ڻ�j��x��6���1��G��  �  �B���b�>b��$F��Gl���|��Y���a ü���������g���h����g�t�N�.�G��S�#o���������_���ʾ�%Eü=y�����&���>��Ă~��b[��R<��!��8���� �һ�f���^��-묻j`��T�ǻ��_j��8�)�/���L�kn�C���$v���ۭ��S��p�¼ܿ��-�������VP��~S���]��'J��I���Z��{�Iz��`0�������¼�h�������m������D-r��KP�#�2����R�S����ɻP����嬻�$�����Vhϻ��������9�M�W�tMz��ߏ�i����಼�|���%ü*���E������07��c�r��!U��G�j�L�!�c���P�������Y��N�¼ׂ��#ø�N3���E��7]����f�F��)����<�� �ۻ4z»�2�����"����5���Xػd=��
���'���B�!�b��I��f.���T���d��Y����¼؏������H�� H��;kg���N��:G���R��n��㊼5ޟ�+C������"-ü`c��%t���|������&a~�}A[��0<�]�!������]Uһ���������=����TǻZ#�';�S���/���L��Dn�����Ff��ͭ��G���u¼$���Q�������>M��Q��]��,J��I�b�Z�g{�I���W���I>���(��,�¼�{������>��������`r���P�5�2����,�����OʻA���~Z��ݕ������*�ϻ3�~��>�L+9�k�W�Fvz�W�����l���\���E@ü��������:��Y��bs��hU���G��%M��1d��%���������/w��1�¼����3ݸ�M��|_���w����f�k?F��-*��^������ܻAû>���'���튱�����ػ�������'P'��  �  l�7��b�͸��'>��������Ӽ���|\�6�߼�~ϼ�Q��ힼo����r���i�5�w������ؽ���Ӽ2=��Q��߼"^ϼ}��;L�������W�hO/����s컐Ȼ�`��oj��\,���{���_��eե�t����ڻ&������D���q��k�����z�żUټ���0U�aRۼ�>ȼ7į��Ŗ�Q��]"m�S�k�@����+��嬼�ż͎ټX�优弣�ڼ�2ȼ�կ��G��w�cBI��\#�6��e�޻����k^��_��NW��'4��ˠ�������dĻ�{绯���'+�#�R�L���@��x���zͼ�޼����㼠�ռ*j��&0��k*��cpz�<j�Gop�y.������a���ͼQa޼y�*���ռԐ�����3��� g���;�o��)��̍һ����Ρ�s���Б��0��B���費�λ����yB�5y7���a�̠���&��'彼ŐӼM���A���߼�`ϼ�1���˞�oL����r��i�,�w�7̌�+_��j����Ӽ�!��8�Dy߼ZIϼ�i��C:���냼��W��,/�&���'�3�ǻ�����Iѓ�;��� ��v�����enڻ���v����D�w�q�hZ���󬼓�ż�HټD�优L张Kۼ�9ȼ.����Ė��Q���'m�T�k������3��5לּ�ż��ټ���/��ۼ�GȼT쯼�_���:w�{wI�:�#�)����޻�n��_ԧ�R���ʒ�����6��]��Q�Ļ�������R+��S�.���U������ͼ.1޼��F;��ռx���	S��xN��׹z��Oj�L�p�#R��!0������.ͼ�~޼w-�����ռH���~4��<���Jg�<�������ӻ���V��ג��R[����������|i��Iϻ�T���y��  �  x�5���h�������X�Ҽ�i�8�����f ���o뼲�м�����֙������u���y��y ������*׼�q��d �X{�$5������˼ƫ�t���b�\���+��7�U�ջi����򊻕���ۂ�!����������nlû�񻝼���E���{�5��۽��Nܼ�s��G��������AǼvN��^Ԓ��V�����������R���ü%.༤�����f������hN߼�W��N���4��Y�J����e���!KǻX��4䒻Ņ�������@��L|��ǖ�������лb��d�&��yV�������iȼ9弘c���A�� ����"ڼ_(��������������a=��^E���_��fvͼ��3u���t��3 ������ռɛ�������n�{�:��c�!������=���X��N��+I�����9���㜻:Q����$z��5��h��q��������ҼPQ�6���������P�E�м����+���@u��<Q���U���ܞ�W칼

׼+S��V �xn������:�˼�����t���m\�ø+���>�ջ�c��F���_���ش����������Q���R���ûpn�˒�3bE���{�$���˽�=Aܼ�g���A�t�c�����C�ƼVM��Ւ�<Y��:����ǐ��Z����ü:�g�����������c߼�m���Ӡ�%M���K������
�ǻ�w���X��8���Q��쮃��扻�������	ѻ���.%'���V�����"����ȼQ�w}���O�� �����DڼL������Y!�������b���i��󂰼��ͼk���������@ �B��# ּ񴶼����)o���:���������]���=ގ�#Յ�NЂ��6�������`���ɷ�`��Y���  �  l�7�adp�+ܙ�FB����ă��:�	����O	�~@��CD����󀥼�9*��H㕼�����ȼN,����
�P���	�R���ڼ�������b�.�,��K��#̻����}n��Ɂ��*x��Hv��}�����v����Ը����8��I��₼�ͥ��Tʼ�c���<��i��s��3����ּ=h��䝼[7���h��0����*���Ӽ���&k�;�Q����n�＃=μ.é��}���O�m'�?!��ݼ����Uˈ���}���u�ѻv�E{��p7��H����ƻz���.5'���[�`�����$ּ�\���%���K����i�#�˼������JH��J��=������ݼO;��Yh�����e
��;;�v:¼�����<w�d=��|�8�ܻY>��q������z��=u�V
y�7���?-��mh��J�ֻ�6��[7��3p��ę��*��h��mk��u�	��2A	��!��w#�gl��]��Q�����L�������aȼ,輅��ȳ
�2���������ڼ5�����b�r,��'���˻�a��,��<s��yw�e�u��c|��^���a��{���v��t��H��Ђ�㼥�FEʼOV����#��2��"�K.���ּ!g���䝼�9��Bm�������2���Ӽ�
�r��B���S����＝Sμ�ک������<O��]����O��z���>����~�ܣv���w��䀻����z�� ǻ��`'�
\��,������;ּdu��:�Q��[�!����[	̼<������in���o���ݢ�j$����ݼ[��Hw���s
��%�DT�eS¼
֝�qw��G=����ZQݻ����~�x9���{��Gv�z����r���W߬�_Y׻"l��  �  ?�8�5�s�����i¼����:X�������&r��缎uƼ����T��	���+���xb��֜ͼ�*��A��m����T������@B߼��������[e�X-����y�ɻ򝢻�h���:~���s��q��x�ل�����o���G�综��L�J��ۄ������μ�9�u��J�SQ�A
�����ܼC��dɡ�R����ۑ�x��`����iؼAG�����f��޾�:M�2�����Ҽc+��Y���_ Q� j��r���똻8߅�ڐx��<q�z!r�׵{�X9�����Ļ�\��,�'��Y^�z��y���,,ۼy����
��q������2�� Ѽ�G���@��ﲐ��Ҕ�¦��¼�Q㼈� ��m��E
��h���Y�Ƽ&�����z�f>��P��ڻ�E���[��(遻X1u�?�p��Et�gÀ� ��?e����Ի!�
��}8��\s�l����R¼������qK�0��m���b�����RƼy���/���m���g��>���yͼa	�*2�A_�ŧ�O������.߼IṼ�y���8e��4-�Ɲ�|Qɻ}O�����f�}�>�r��q��ew��|��LG������组��c�J��Ʉ�����i�μG,��kE�M��	
�M����ܼ)��'ʡ�󲒼(���p~�������sؼ'S�����$��y���V������Ӽ�B��/���h4Q���8��V����^��^R��Auy��r���r���|�v����b��4_Ļ����$�'��^�d���b���+Cۼ����1�
���O�������;ѼRm���f��8ِ������榼u�¼�s�p� ���������u����4�ƼY̠���z��>�4��p'ۻO���jۑ��k��:v�"�q�VKu�NC�������۩�Pջ���  �  l�7�adp�+ܙ�FB����ă��:�	����O	�~@��CD����󀥼�9*��H㕼�����ȼN,����
�P���	�R���ڼ�������b�.�,��K��#̻����}n��Ɂ��*x��Hv��}�����v����Ը����8��I��₼�ͥ��Tʼ�c���<��i��s��3����ּ=h��䝼[7���h��0����*���Ӽ���&k�;�Q����n�＃=μ.é��}���O�m'�?!��ݼ����Uˈ���}���u�ѻv�E{��p7��H����ƻz���.5'���[�`�����$ּ�\���%���K����i�#�˼������JH��J��=������ݼO;��Yh�����e
��;;�v:¼�����<w�d=��|�8�ܻY>��q������z��=u�V
y�7���?-��mh��J�ֻ�6��[7��3p��ę��*��h��mk��u�	��2A	��!��w#�gl��]��Q�����L�������aȼ,輅��ȳ
�2���������ڼ5�����b�r,��'���˻�a��,��<s��yw�e�u��c|��^���a��{���v��t��H��Ђ�㼥�FEʼOV����#��2��"�K.���ּ!g���䝼�9��Bm�������2���Ӽ�
�r��B���S����＝Sμ�ک������<O��]����O��z���>����~�ܣv���w��䀻����z�� ǻ��`'�
\��,������;ּdu��:�Q��[�!����[	̼<������in���o���ݢ�j$����ݼ[��Hw���s
��%�DT�eS¼
֝�qw��G=����ZQݻ����~�x9���{��Gv�z����r���W߬�_Y׻"l��  �  x�5���h�������X�Ҽ�i�8�����f ���o뼲�м�����֙������u���y��y ������*׼�q��d �X{�$5������˼ƫ�t���b�\���+��7�U�ջi����򊻕���ۂ�!����������nlû�񻝼���E���{�5��۽��Nܼ�s��G��������AǼvN��^Ԓ��V�����������R���ü%.༤�����f������hN߼�W��N���4��Y�J����e���!KǻX��4䒻Ņ�������@��L|��ǖ�������лb��d�&��yV�������iȼ9弘c���A�� ����"ڼ_(��������������a=��^E���_��fvͼ��3u���t��3 ������ռɛ�������n�{�:��c�!������=���X��N��+I�����9���㜻:Q����$z��5��h��q��������ҼPQ�6���������P�E�м����+���@u��<Q���U���ܞ�W칼

׼+S��V �xn������:�˼�����t���m\�ø+���>�ջ�c��F���_���ش����������Q���R���ûpn�˒�3bE���{�$���˽�=Aܼ�g���A�t�c�����C�ƼVM��Ւ�<Y��:����ǐ��Z����ü:�g�����������c߼�m���Ӡ�%M���K������
�ǻ�w���X��8���Q��쮃��扻�������	ѻ���.%'���V�����"����ȼQ�w}���O�� �����DڼL������Y!�������b���i��󂰼��ͼk���������@ �B��# ּ񴶼����)o���:���������]���=ގ�#Յ�NЂ��6�������`���ɷ�`��Y���  �  l�7��b�͸��'>��������Ӽ���|\�6�߼�~ϼ�Q��ힼo����r���i�5�w������ؽ���Ӽ2=��Q��߼"^ϼ}��;L�������W�hO/����s컐Ȼ�`��oj��\,���{���_��eե�t����ڻ&������D���q��k�����z�żUټ���0U�aRۼ�>ȼ7į��Ŗ�Q��]"m�S�k�@����+��嬼�ż͎ټX�优弣�ڼ�2ȼ�կ��G��w�cBI��\#�6��e�޻����k^��_��NW��'4��ˠ�������dĻ�{绯���'+�#�R�L���@��x���zͼ�޼����㼠�ռ*j��&0��k*��cpz�<j�Gop�y.������a���ͼQa޼y�*���ռԐ�����3��� g���;�o��)��̍һ����Ρ�s���Б��0��B���費�λ����yB�5y7���a�̠���&��'彼ŐӼM���A���߼�`ϼ�1���˞�oL����r��i�,�w�7̌�+_��j����Ӽ�!��8�Dy߼ZIϼ�i��C:���냼��W��,/�&���'�3�ǻ�����Iѓ�;��� ��v�����enڻ���v����D�w�q�hZ���󬼓�ż�HټD�优L张Kۼ�9ȼ.����Ė��Q���'m�T�k������3��5לּ�ż��ټ���/��ۼ�GȼT쯼�_���:w�{wI�:�#�)����޻�n��_ԧ�R���ʒ�����6��]��Q�Ļ�������R+��S�.���U������ͼ.1޼��F;��ռx���	S��xN��׹z��Oj�L�p�#R��!0������.ͼ�~޼w-�����ռH���~4��<���Jg�<�������ӻ���V��ג��R[����������|i��Iϻ�T���y��  �  �B���b�>b��$F��Gl���|��Y���a ü���������g���h����g�t�N�.�G��S�#o���������_���ʾ�%Eü=y�����&���>��Ă~��b[��R<��!��8���� �һ�f���^��-묻j`��T�ǻ��_j��8�)�/���L�kn�C���$v���ۭ��S��p�¼ܿ��-�������VP��~S���]��'J��I���Z��{�Iz��`0�������¼�h�������m������D-r��KP�#�2����R�S����ɻP����嬻�$�����Vhϻ��������9�M�W�tMz��ߏ�i����಼�|���%ü*���E������07��c�r��!U��G�j�L�!�c���P�������Y��N�¼ׂ��#ø�N3���E��7]����f�F��)����<�� �ۻ4z»�2�����"����5���Xػd=��
���'���B�!�b��I��f.���T���d��Y����¼؏������H�� H��;kg���N��:G���R��n��㊼5ޟ�+C������"-ü`c��%t���|������&a~�}A[��0<�]�!������]Uһ���������=����TǻZ#�';�S���/���L��Dn�����Ff��ͭ��G���u¼$���Q�������>M��Q��]��,J��I�b�Z�g{�I���W���I>���(��,�¼�{������>��������`r���P�5�2����,�����OʻA���~Z��ݕ������*�ϻ3�~��>�L+9�k�W�Fvz�W�����l���\���E@ü��������:��Y��bs��hU���G��%M��1d��%���������/w��1�¼����3ݸ�M��|_���w����f�k?F��-*��^������ܻAû>���'���튱�����ػ�������'P'��  �  �s\�w�q��L��
���2햼�*���š��q������������{��Z���=��)*�hd$�[e-�JXC���a�U�������ړ���6���[��NМ�8����P��3�����l���W��IB�Ю,�����i��g�1�׻mgԻ�~�o��<��'#�r�8��/N�hnc���x�����Ȑ�v����ɟ��ܡ�մ��$��<���Čp��P�@�5��l&���%�*>3�&�L��l��̆�!�������񹡼>.���]��BÑ��Ǉ��z���e�-WP���:��I%����"���F�ӍԻ�UֻK绒M�"!�� *���?��-U�^`j�'r�
��㓼V��������e��o`��'񑼓E���Pe�:&F���.��e$��(�$�:���V�T�w�oҋ�[���ٟ��ȡ�󬞼Aė������\���s�U�^�HI��3��G��C
�� �^ܻ.eӻ3fڻ��ﻃ4�o���L1���F�}=\��cq�[4��x��{Ֆ����ˬ��
X��|v��Hm��|�{�dZ��G=���)��!$�U#-��C��a�#z��w~���z������F��E����攼�?���䀼�l���W�h&B���,��g��>���3�׻pԻ��I�������"��}8�N�lDc��_x����V����������ҡ�����*���)���p�p�m P���5��q&���%�K3�ѱL���l��؆�$�������ˡ��A��s��6ڑ�=�����z�]�e�>�P�w;��%����~���O�⻿ջ��ֻ���-���R��O*���?��WU��j���61������[��|��I���{��l���d��ّe��iF��A/�m�$��(���:��W��&x������w��I���z㡼;Ǟ�mޗ�:���
x��
�s�!�^��I��3����;�
���7�ܻ��ӻ��ڻ�j��x��6���1��G��  �  �|���숼����4I��/@�� ߋ�����h�� �u��_�0qF�.�,�;���xd��� l�n2�d7L�k�d�Ƽy�m��������N��6[��#��{w���ꇼ*ぼ|1r�'�[��B�	�(�v��%�e��h ����Ւ6� oP���h�Ğ|�k���c#������q\��=猼�����������n��bW���=��$�n�:���;�H_�S"��:���T��0l��B��h����������I�������f�����>H~�%�j�S��-9��� ��s�P��������&�b�>���X���o�#���bO��n��x�Q���k��牼�+��؇{��Hg�t�N���4��v�,3�ZV��g�����)��NC���\�v#s��5�����܄��`���>�����_D������|x� jc��J�V�0��&
���"��o���.��G�"�`�fv�a��T҈��䋼1��n(��Bǋ�=���	���Wu�}_��6F�U�,����Qm��$�l�
��.�32���K���d�H�y��}��߀���<��vJ��0���g���ڇ��ҁ�,r�/v[���A�?�(������~� ��O���_6�==P��|h��p|��w��`��Yy���K��،����|���ۘn�gXW��=�h�$���`���D�+l��c"���:�-�T��Ll��b��z��ת��>ǌ��`��嵌�v����0��e�~�D$k��ES�l9��=!�}����X��%�G&��.?���X���o����Oc���/�����e��%�������D��+�{���g�O�]<5����u�}��n��f�J>*���C�Y]��\s�KQ��l2��b����,���Y���8���a���;��ٽx���c���J�s1��R��r
��[��>	��%��L.�c�G��a���v��  �  Ū��̱��ٝ�s�����ڷ���ip�;D[���E�BT0����q����%ڻDԻR�ݻc(��Б�����#5��J���_�Bu����3���N��4��a桼����ޗ�O���<v�$FU�o9�m(���$�8-0���G��Wg��>�����ޜ�v����ڠ������h��i����U~�"Bi��T���>�� )�
��q�0,�ֻ�ջ��㻠��u��j�&�<���Q���f���{��[��I��%Ě�e_�����t��������ⅼ��j���J��2�#%��&�۲6���Q��Ur�Y[��/���p ��Hڡ������"���7��/��0Gw�9)b���L��W7���!�ru����)߻[�ӻ�1ػ�o��4�����-� PC���X���m��t��5ʋ��_�����Fa���2�������M���/�_�яA��;,�m$�c�*��>�)\�dp}�3��"���.������������Z���錼����9p�g[�ݷE��0�/���6�He�ٻʈӻ�ݻ����Y��}���4���J���_��t�����#���?��!����֡������̗�A��sv��U��?9���'�=�$�~�/�˴G�y#g�%��E���wƜ�W{��GƠ�ʔ���W��Z����;~��+i� �S�A�>�h�(�h��n��.�Rֻ�.ջ`��F@��,���&��:<� �Q��f��|�^q���`��vݚ�Pz��l������������k��"K��G2�a%��	'�%�6���Q�Y�r��r��0������������5��OK��w1��crw��Wb�M�m�7�"��������9�߻�OԻX�ػ���Ms�:����-�ȈC���X��n�l���7勼�{���.�����~�����ݏ�n���`���A�8�,��V$���*�
�>�7r\�׵}��S������  �  �üަ���ƶ�y��k9��EY��a��:A�'�%���������H׻ڟ����������o^��*Ļ�ݻ����ѐ��+���G�Z�h�}~���e���3���������ɀ¼mͺ�ɼ��_◼� ���sb��KL�)H�_�V���t�B{��5L���䴼���i(ü�����I����َ��Wx���U�?7������"뻁)λsS�������U��Ņ���X˻[o绡y���5M4�]R��0t�橌��p���[��U��¼����_`��5[��ƴ����x��Y��H�c�J��_������r��џ��b��t���G¼�������g��C���cl��,K��X.�����:�,�໎!ƻOI���g���u���
����ӻ�l�[2��"�o�=�o]�C1��A��Eq���1���ǿ�� ü�,���Y��ö��������l�ޜQ��G�ԋO��0i��h��em��O������z�¼��������`���!���A��c�`��	A�b�%�����P�� �ֻ�+��@��#9���겻�û:ݻSZ��Wb��n+���G�D�h�hn���V��b%��0r�������p¼��������z͗��邼fCb��L�2�G�EeV�b�t�L`���1��+˴�����ü����	���y���ʎ��<x�ѺU��l7�b�������#λ�U�����g�������z˻��b�����m4��?R��Xt���������]u���	����¼�������<{��CՐ�*y�LY�M�H�p�J�.<_�#π�}�������x���¼ZZ¼�ƺ�6���z������w�l�YK��.�^��q����Йƻ�Ĵ��䬻`�$����AԻ���l�""#�2�=�pH]�AL��� ������<O���濼jAü�O��[~��"ݞ�v݉��7m�"�Q��mG���O�ni�����#���祯�
>���  �  h�hἯ�Ҽ����¢��G����_��5�����pͻ7���͟��N���[��U���.���\����Իy��0��H.>���i����������O�ּng㼊���ݼ#�˼,��kΚ�|E����o���j��0|�o|��%���{����ּ�������jݼ��˼�8���͙��w�ˇP��@)�i6
�j[�{�»�Ū�� ��� ��԰��}ҙ�����G���t�໡(��K%�a�K�.�y�r�3E���gɼ%�ۼbY�)O�l�ؼVļk��rؒ��0��0k�z�m�q4��
��_%��}sɼjܼu��V)�Qkؼ	}ļ"����쐼Bo�~B�&����)�ػ;���g���������"��D˝�5��AsɻT|�-X�/1�=EZ�:R��J���lȹ��^м��ZC�=���ҼeU����K����.v��vi�9�s� `��*��_���I~мXc�VJ�bLἶ�Ҽk������n0���V_��\5�9���f�ͻ򯱻�\���ܔ�Oꑻ����l¢������Իû���p��	>���i�{������7���I�ּ�X㼲�弒�ݼ��˼���x����,���o�m[j�f�{��`����������,�ּ�㼯��_Uݼb�˼�&�����v\��pP�~-)�t'
��E廮�»����%#��+����|왻����!ѿ�; �{E�`l%�%�K���y��ؖ�b]����ɼ��ۼ�v��m�'�ؼ�vļ"�������ur��pk�~n��Q���%��6?��X�ɼ`2ܼ¡�W<�{}ؼ�ļ0�������4o�ΨB�<'�}����ػ�)������������������D�������ɻ;��ď��e1�U{Z�im��͟�$幼�|мT8�e������Ҽ�|�����#ɋ�{�v�>�i�Dt�R����P�� �����м`���  �  ���Ά���!��
ѼO@��-Ɛ� �e�@3�e��2�ݻ�����9���֌�焻�͂�M!�������u��/��K��;�=��Rr�ܗ������׼��� �_n�����c�O�˼��l6���͆�hۃ�����m���⾼|�ۼ��+�*,�w������>�ƼD��xU��Z�S���$��� � hλ󴫻̕�`#��Z>���킻�"��<铻U���Ŧɻ���V ���M��Ⴜk����ü�༾��w��>�������޼V¼�Υ�ɶ���:������ړ�Lī�a�ȼ̓�;���4�<�<S�¹ڼ�
���a���x�3�B�r��_����������h���r��-����+��v������pػ��s.�i_��,��g���s�ͼS_�$���z�r ��sռ�J��.���ъ��=������d���GҼ���������j��e�"�мq(������;�e�a3�X���`ݻ򋵻�͛��h��=x���_��7����!�����������Zq��f=��2r�s͗��q���׼�́ ��f�����SP��˼�֮�w������쿃��ݍ�����ƾ��ۼ���4�i ��r�����\�Ƽ74���G����S���$��� �Rλ����ƕ�w%��rH�������<��B��Uè���ɻ2��T9 ���M�v���㢢�T3ü[�༻���A�����%����޼�&¼�؏�I[��iՅ�����Rૼd�ȼ���-���)>���e�6�ڼ]��t����x���B�'�����`��!������܆��邻�g��������
{��/�ػW��Q.�<�_��G��e�����ͼ�}鼁��K��� ��>�L�ռ�t��쮝����"h��SE�����?��?mҼ���y����  �  ��fV	�����߼F9��)㗼��l���4�6V	��tԻL��䎑�;o����y�W@v���{�х����<����V����-*@���z��П��Tļ�����n�
����H �������ۼ�l�������ΐ�T���Ǜ�����f�ͼ�,������������b����<Լ��r7���X���$�9���FĻ`����|��m5����v��Hv���~��������P��ʷ�.��a4R��]��5ʫ�\6мtj�h�M:�L�R��JT�:/Ѽ|���6������A������T����Tؼҷ��� �����T������Nȼ�ã������E��8�WS��p���+��	���n�{�7�u��w�����
��7{λG�X/�k�e�4ߓ�x���ۼ����n�����\
� ��P�ÛƼ\���$┼v�Q������\"ü*�����h�	�K�IH	�o���?�߼f!���˗��l�=�4��%	��Իך���$�����x��gu���z��j��w����R��+�Ⱥ��@���z�y�pGļ{�(��P�
�$���������p�ۼ�U��cw�������}��]��fq���ͼO�H��O�������U����*Լ�௼�)����X�6�$�����Z0ĻB����v��w7����v��lv���~�%߉�����.������J���YR�Nr���ૼ�Nмۄ��v�1I�������u��PѼX���ã��S$��߿��� ������nؼ��������^���԰�Y_ȼ�գ����SF�hd�����ն�e����*����|��lv�9�x��d��B����|��>�λFN��L/��f������'��mܼ� ��L���o
�3��y��Ƽ����������|��dߦ�?Jü��^���״	��  �  ~
���Ɔ��{� a���A���!�����ռqխ��v���2x�W�]���M���E��C�� G���P��|b�����&��Lµ��	༑_
���(��H�aog��2������扽����)�w���]�}VB�l�*��d�����,#��"7�:nQ���l�ρ�д��墉�&X��Zps���V�P7�y��3��8#ǼQݢ�������m��W��:J��D��CD��BI�_6U�&�j��M���o��3�¼�c���'b3��dS���p�A_��)Q��$���̂���o�ErT���9�6�$�b�ch�1�(��c?���Z�u�⯄����������P���j�PoL�	K,����U弢׹�����ꁼu�d���Q���G�B�C��?E�?SL�%[��dt�����d���ءм��<D�c(>�ע]���x�V���􉽱�����G�f�=K��1����}���vz/��6H�t�c�)�|������������~{���`�!�A���!�W�q�ռ�����]����w��e]���M�b�E��C���F��OP��Kb����%�������߼�X
���(���H��ig��/�����<㉽]�����w��]�JJB��*��V����+#�]7��^Q���l��ǁ�쭈�s���2R���es���V���6��q��&���Ǽ(բ�������m�*W��;J�8�D�OMD�UPI�!HU�$�j�[���~����¼Kw� �#n3��qS���p��f��$Y������Ղ���o�o�T���9�7�$���/y��(�hr?��Z� u�C���˸������T��͏j�%wL�;S,�Ŗ�6i��칼�+����$e�R���G��D��{E��L��_[�@�t�ˍ����ݼмn��Q�}6>���]�@�x��
������h���r4��f��SK�M2�� ��)�)����/�'LH�`�c���|�S���  �  ᆽ���#v�Ӊ\��o>�c�����ռ�r���ܑ�F�{��'a�g�P���H�òF��J�V�S��f�����j���"���߼����O&��OE�þb���z�$����"���:r�{�X��N>�~�'�Yd�3��f���i3�n�L�N�g�p�}�����~��7g��rRn���R��4�|���v����Ƽ�ʣ�B���_q���Z�(NM�$NG� G��JL�p�X��:n��臼�t���}¼���jX�U�0�riO�}k�'w��50������Ψ�m;j�v�O���5��!���(n� q%�tp;�i�U��o���������n����|��e�S�H�в)�y�F+����D��𗃼"�h��+U��J�<�F��H��}O�̪^���w�
$��󰪼'мY���+���:��JY�q�s����ĕ�2���_y���a��F��U.�b��M(�ߍ���+�QD���^�+w��能Fن����v��}\�d>��������Լ�Z���Ñ�<{���`�L�P��H�U{F�S�I�4�S�p�e�B���sU��J��\�޼����I&��IE��b���z��q����z���0r���X��B>�0�'�V�C��
��Z3�
�L�Fxg���}�9���`x��Ia���Gn�C�R�e 4����i��C�Ƽ�£�<���Wq�d�Z�OM�BSG�c	G�+XL�/�X��Pn����� ���C�¼d��Jc�K�0�xvO�'�k��~��+8�����)��BMj���O��	6��!�0#��~�Ȁ%�;���U��o����Տ��Ms�� }���e�9�H��)�`��>�,��\��;����h��dU���J�"�F��IH���O���^�U'x�+@��n̪�&BмG����8���:�vYY��s�	
��jՆ�ݏ���sy�y�a��G��l.�����?�Ϥ�,�nD���^��#w�B��  �  ��{��v��g��;P�U5���� ��HԼ�3��M���������l�g[�;2R��O��S��|^�0�q�J���훼�:���Mݼ������z;�b�U��Ck�^�x���{��s���b��]K��2�������5W�L��b�(�JW@�!�X�m��zy��]{��`r��`��G��,�{��;��<�Ǽ%g��܉����|�G�e��XW�OP�I$P��6V���c���y�2L���Q��^vü&��)����(�<D���]���p��z�+z�t�n�73[�]C�<++��p���g������40�T�H�/%`�g@r�'O{�X�y��-m�"qX���>���"�pB�X��"ӻ�/����'���t�o�_��<T�آO��_Q��Y�j�i����(��Z���C�ϼ�����k12�TM�X�d��8u�<�{���w��i�~mS�B�:�$$�0�������X�!�!8���P���f�9ev���{�|v��
g��/P��I5����= �~1ԼK������{���Wl��.[�p�Q���O�rhS�@G^��fq��2��K؛��'���<ݼU|�)���s;�z�U�w=k�ңx�A�{��s��b�SK���2�T��t��qH� ���(�H@�I�X��m�omy��P{��Tr��`�s{G� ,�������|Ǽ_��󃏼�|���e��YW�q�P��-P�DV�M�c���y�DY���`����ü��������(�-�D���]���p���z��;z���n��D[�MC�6=+����;����d�C0���H�01`�-Kr��X{�*�y�6m�"yX���>�H�"��K�Q��黼����A���Mt�D/`��xT���O�ޜQ��Z�8j�؁�E���ڭ�V�ϼ�������a?2��bM���d�:Iu��{���w��-i�؂S�|�:��:$�I$�������3
"��-8��P�g��uv��  �  S	b�^�˟Q��?��1)���Z>��w�ּ黸����<Ŏ��	���o�#%d�'a��e���r������l���ӥ�nԾ��F޼f�.���2.�ŖC�M�T��_�V�a�'oZ�(FK��7�}�!�rp��X���U	����~t-���B�A�T�4�_�˰a��Z��K���7�D�!�Da�O�˼���FX��Y���~�z��Sj�4b�ʬa���h��ax�����7���^���rȼ��I�����5���I�xYY��Ja�4.`��V���D���/����Ц
� ��9����_d�
�4��+I��Y�Ea�4P`���V�ǾE���0����W�	⼦����7���;��|	��J;t��f�a�?0c�|+m�VP��ꌼ���q�����ҼT���1-���&�Ӷ<���O���\�]�a�R�]��Q�>�̟(����@��`c���5���D&��;��&O�w�\�F�a�=�]���Q��	?�&)����O'����ּ4�������+����퀼��n���c���`���e�%Tr�d���6T������~����4޼��*��8,.���C��T�M�_��a��fZ��<K��7���!�yc�*������F	�����e-���B�={T��~_�S�a���Z���K�<�7��!�Z��B�˼���qR������H�z��Tj�[!b��a�:i�:sx�����D���m����ȼ
-�	�W�ؓ5�`�I�5hY�'Za��>`��%V�3�D�h�/���P�
�1��I�*���r�9�4��7I�lY��Na�*Y`��V��E��0�Q�a��/�f ¼�P���V���%���vt���f��La��nc��im�,��!���Ȟ�=ϵ��Ӽ&����:�m�&�3�<�2�O��]��b���]��Q��'>�{�(��������y�)����8Y&�B�;��8O���\��  �  �DD�u`B�� :��=-������w���	���ȼĵ��j���kk�����:����|�V��H<��%|���R���$��l�ͼ���̪��C�"X!��d0�:l<�aC��C���<�m�/���PL��[��j�N�开>����	���(�I�7�t�A�eD��=@��96��@(��g�.q��󼳁ؼ�Z���B���������.����}�$M}��X���Ì�/K���*���ڶռ���R��s��I�&�4�4�U?��5D�T'B�o9��*����u��h���C�G�v}���`�j��.'.�y�;��DC���C��s=���1�2#����N���Qgм=P��+��4����F���ہ�T|�HG�����}֐������o���-ƼF޼�d��K��M��e�+��8���A��XD���?���4���$�!�ê�T�P
�6F�Y�����"�s43���>��5D��RB�A:��1-����,��(�����༞�ȼ,����j��UN����������R|� 8��D���`���8����>�ͼ���i��I<�;Q!�,^0��e<�(ZC���C�U�<���/����@��B���N�
��!�A�(��~�(���7�x~A�SYD��2@�a/6�m7(�_�j�{�wؼS���<����:��/���}�uV}��_���̌�V��t7��������ռ��������&���4��c?�ED�d7B�09�,�*�����[���
e�f7�ۛ��o�w�3.�I�;�eNC���C��|=�]�1��#����X����+м1j���F������e��y���	�|���������������򌱼JƼ,޼|�������y�+���8�M�A��iD���?�!�4���$��Q���6��5��p�+�D&�'�"��E3��?��  �  �+'�U9(�O%����o�������4���ϓ��Ѽ¤��򳫼=������e�����a��iw�����)wռ���:�������;���u ��&��_(��F&�]��0�._��u�k�ؼ�ɼ��Ƽ��м��~����?�b����#��(���'�F#��Y�p�������:2�޼	{ʼgS���P��o���T���񑼻R��F���D���Dȼ��ۼ��� �3
�9��~m�d�"��5'��"(�p$����k��׀����pQҼd5Ǽ3�ȼWQּDf���7��uF�g�%�_W(�	~&��-!�������{�����Y�׼��ü�H���n��[R��le���N��)͛�#é��k����μT��S�������`��]��x$��(��v'�Y%"�rB���s���ݣ߼hRͼ^?Ƽy�˼�&ݼ�m��ف	����B!�T'�,(��%�����������i���y�e�мՇ�����������E���t���IZ������%^ռ@�����������о��n ��&�^X(�?&��T�~'��T��^�ؼ��ɼ>�Ƽ��м���T����1���&�#���'���'�<#��P�m������v(��	޼kuʼ�O��fO���o��XW��@���nY������N���Qȼ��ۼ�（� ��
����y�Ȝ"�D'��1(��$�:� ��Ǒ�����rҼVǼ��ȼ'oּ*������MQ�d�%��`(��&��6!�ʲ�?�6����=�꼨�׼4ļ�g�� ����s�����Qp��%4㩼����.�μrp�2o����������7�$� (�ֆ'��6"��T�7)�Ұ��T�߼f|ͼFiƼ�̼�Nݼ���֓	����,R!��  �  �m��>����,��#����������������㼒ͼ ������ʩ�񓯼�ƽ���Ѽ��ԝ������d�����G�>��!���[��6��R��U�߼��ɼ�Z���2�����a������ЎռQg��� �H�	��E�X�P���C����<������F��!��=�ۼ�Ƽ�ᴼ��������_��9�ü�=ټ��ђ�����g��X���:������_��T�
�������׼y�¼>����O���a�������'ǼDݼ���P(��=�����;�����=��j��&����?d	��b ���:Լ����٣���թ�-}�����ʼ��༴p��X���V������e�o-�($�L��S�h��V��':缞�м<����ޮ�E����ԭ�pź��μͬ�0�����_��1�Q��O �:�=�����
����Z����h��̼\߹�x^��9����r��9���$�Ѽ��*������Z���/?�6�����~�kT�"��e-��?����߼�pɼ�B��K�������E��^����sռ�L�� ��	��:�eM��y��:���m���:����������ۼ�Ƽ<ⴼq"��,���Ff����üBHټN#�1��,�7�������%G�B���������
���~�ؼ��¼񻲼�o��R�������7CǼ� ݼ��/3�H�"���D�(��2G��t��1�� ��q	�`q ��-뼛ZԼqƿ��ư��������.<���ʼ7��������Zd�@����r��:�2� �����-z��W_�M�м�ϼ����v���h����뺼@Cμz�伛"���,��  �  ����Z��ǘ�u`��K�,Y%�MH(���&�}� �mN����Y��dܼtq˼�vƼ�9μ
�p?�����o��C�"�H�'���'�:$�����w���u��^���W�2�ͼ�x�������E��^��g����ᖼ�K���Y��nż��ؼ���ǳ��&�����!��!��&�zT(��o%�{����������Tռ�Hȼ��ǼASӼ|�PT��|�Η�	�$��6(�x'�9"�&��}��~	��R ���!�ڼ$Ǽ�6���£�����v����������� ��"P��6�˼߼!7�sg�ڋ�(x�5���#���'���'�y`#�1�o��D��Đ�D�ϼ~�Ƽ� ʼ��ټi��/����Z��5z&�P(���%� 	 ��D���z�#���1��AԼ���b`��e0�����V9���F��ȝ�#������|Ҽ/��|q���u�Ɍ��T�(@�M%�'<(���&��� ��?�$������B�ۼyN˼XSƼ�μ������o��D��\�"���'�}�'��0$�x���o����m��N��"F�O�ͼd���ᨼ�-������}���ǖ�1��9?����ļ��ؼ��{����~�%����F�!�K�&��N(�k%�˺�K������뼨Tռ�Kȼe�Ǽ�YӼ"#鼣Y������T�$�@(��'�=D"�7�����	�>a �8�H�ڼ�CǼ�V��㣼�ߗ��ڑ����)���;��Ui����˼�3߼�K�>q�x����Z��ĝ#�E�'�v�'�vn#�3@�J�g��F�㼑�ϼ�Ƽ�Dʼ��ټ{��o/���������&�R](���%�� ��Q�[��F��0���%���bԼ����j���pV��-.���_���l���일k���b����1ҼP���  �  �|�`��<����5.�ù:���B��)D�?�>�bu2��!�{-��e ����YG��(�=����{�%��5�e@�3qD��gA��>8�9�*�s�������$�ܼ�ż0u�����
8��a�����B�|�K�������ܗ�':��m���x�Ѽ�]�2+����.�#�N�2�1�=��C��
C�O;��H-�S �D{
�A8����缇��Ь��������v+�%�9��yB�)!D���>��4��%�u�����QUԼu���{��Kg��b���肼��|��~�֑��F���d✼�D����¼ �ټr����K	��I�6)�6�6���@�}eD��#A��
7�U�'�X���'�Q�Ho弬��B���1������0�~m=���C��C���;��/��k ��T�� ��P弌{̼趼�<��˒��芈�怼�=|��X���v���
��W�����w�ɼ�b�@G��p�������-��:�b�B�sD�0{>�Kf2���!�v��S �fy�{"��]}���V�%��5�pW@��dD��\A�58�.�*���
�������ܼ>�ļZb������Q"��N}��$�~��|�k1��;܊�R×�!!��Dm��p�ѼMH�!������#�ڝ2���=���C�4C��;�/F-�����z
��8��F��,��q���?�����|+�e�9�6�B�T*D� �>�4�Ȱ%�-����xm�(sԼ�׽��;��ц���3�����5}��S~���֎�U���\��ޜ¼��ټs����U	��S��)���6��@��rD��2A��7�D�'�.�:�2�2��$꼼����B�^ ���0�4|=���C��*C�L�;�k�/�Mx ��a��� ��m�<�̼����^��Q���h������ԇ|�}��b����,��<w��Gϴ��
ʼ�  �  גؼ�t�����?s*��:@�R��v^���a��B\�CN��:�-%�g�V�����x�"���)�sN?���Q�wP^�� b�z\�5�N���;��i%��������;Ѽ�Y��Ť���'��JE~�r�l��c�gWa��[g�wcu�#ׅ��F��⊩���ü�伏��aT���1���F�HHW��`�]a�G`X��"H�'p3��M�A������b�~i��;1���E���V���`��a�B�X�S�H��O4�������
輛�Ƽ>��w(��q8���8w�xIh��ga��Db�Y�j��{�i��3a���v���ͼ�a𼩏���"��,9�~�L�3H[���a�u_�j�S���A�E4,�_�����ϟ�\�A?�?�"��28��;L��[��a�@_�-#T��pB��,��R��� �BܼS,�� ���D_��邼�^q�j$e���`��Gd���o�b���ʋ�������yؼu\��9���g*�4/@�PsR�Zj^�1�a�B4\��3N�`�:�x%��6C�wq��e����?�)��=?���Q�)B^�	�a�un\���N��;��`%�)��_����*Ѽ5H���������~~�/il���b�u&a�*g�F1u�>����.��Ws��|ü�
伶x�UK���1���F��AW���`��
a��\X�* H��n3�GM������e��l�f�
1���E�*�V�%�`��!a�B�X�6�H��[4�1��h��&輥�Ƽ1"��G��\W��Yvw���h�M�a��~b��%k�`�{�Ɂ��sx�������ͼ�u�ϙ�)�"��79�C�L�U[���a��-_��S��A��F,������_��[o��Q�/�"��C8��KL��[���a�1M_��/T��|B�z�,��_��� �^ܼ�I��S���/���\���q��ke�D"a��d��o�F������{;��o;���  �  m�ּ�n��:���6�U�Q�<,h��w��{��u���e�?yO��6�~� ��Z����^���Y%�?<���T�53j� x��{���t���c���K�N�0��@�_G����ͼl2��O��
���+	i�!LY��IQ�k�O���T�y�`���u�[:��}	�����P���	�ZU$��@���Y��n���y�{��xq��^��6G�P�.�����?���N�)o,��pD�){\�[�o�Y�z��z���o�PR\�� C��\'�~v��	�.z��Ϣ�?1��'Fx�A�b�КU��O��P��W���f��~~�\�����ʋɼH�"F�ӏ-�;�H��Ma��s���{��y�Fl�SaW�'�>�֔'���E�?�#���4�׮L��c�0tt�b�{��#x��7j��_T���9��5�Y�F�ڼ�T��m|���8��p�9n]���R��xO��DR���[���m��^���◼	Ѳ�.gּ�b�p/�{�6��Q�e h�w���{�j�u���e�PhO���6��� �G�M��ɷ��F%��,<���T�	#j�Ix���{���t��c�)�K�;�0�8�s6��^�ͼ� ������值��h��Y�CQ�a�O���T�J�`��nu�z"��h����I;�K�	�uL$���?���Y��n�r�y��{�uq���^�`5G���.�;�l������Q�os,�vD�]�\���o�r�z��z���o�]\�|C��h'����O%�ז���좼eO���x�*�b��U�l#P���P��X���f��~���������ɼ�%�wP�x�-�xI��Ya�*s��{�^y�7.l�esW�'�>�~�'��2�M3��R�B��	-4��L�7�c�+�t�T�{��0x�Dj��kT��9��A�@&�wۼ�q��ߚ���X���Pp���]��@S� �O�o�R�b&\��m��|��g����벼�  �  a�׼Ml��<!�H)@�*^�Yw���y߆�I����u��s]��B��*���2M���O�/�цH��Ic�?�z�`ׄ�!ǆ������Xr���W��>9��������ͼ����E����bv�@�]�O�X H���F��K��%V��j�ѳ���ԛ��1����漙���k+��gJ��6g�:~�����n���<��]Rn��vT��:�Vz$�%��b�	�"�
W7�<rQ�2�k��Q��* �� ��n���j���M�R�.���r�EO��=Ԟ�v����l��W�o�K�M�F��dG�3�M�`[���r��j��Js��42ɼ�@���:�#�5��jT�x�o��с�S���IR��צ|��f�nK��2�F��r������(���?�VkZ�5os��ۂ�xǆ�{���q�y�u-a��C�ߒ$�$g��jܼ���pᕼ������d�#�R�#rI�lF�H�H��iQ��b��P}�z��"9��oj׼y`�?1!�	@��^�7Mw�����؆�铃�"�u��b]���B���*����39�'��ɐ/�	tH�8c��z��τ�H��������Mr���W��59�P��y�����ͼ�쨼�⍼);v�;�]���N�G�G��F�V�J� �U���i�=���ڽ����6��	���b+��_J��/g���}�奅��k��2;���On�HuT�N:��z$�}�'e�T�"�M[7�wwQ�b�k�OU��3$���������j�)�M���.����5켰k����V߆�_�l�r�W��K��G�Z�G�w�M�	�[��s����N���cGɼ�U��LE���5�FvT�ȳo�:؁�����FZ���|�$f�_�K��%2��2��������(��?��|Z�os�'ソtΆ����ڱy��9a��C��$��s�K�ܼ�-��V��������d�ZS�X�I�İF��I�s�Q��Xb��}��6���S���  �  E=ؼܧ��#���C�7�b���|����G	��毆��{��`b��F��`.����7��� ��B3���L�?bh��,���􇽪����|�w��\�i<�������9Hμ�7��y��[�r��?Z�@�K��5E��D�x$H���R�aqf��
���������輑0��.��3N��l�|܁��È�e����?��R�s�� Y�9�=���'����U���%��,;�-V���p��M���F��L'��:₽,
o�T�Q���1��l�ό�C���Ý��!���i�%>T�t�H��D��D�;�J��X��To��ቼ9����pɼZ���%���8��X�-�t��Ƅ�����ds��=@��a?k���O���5��G"��^����,���C��A_�ey��ꅽi�q���y/���e��G���&�����Pݼ��������د}���`�l�O���F���C���E��-N��^���y�ȼ������l$ؼ���y#�V�C�Җb���|����v�������{�vOb���F�]M.�����#�ŷ ��.3���L�^Ph�w$��S퇽�牽����X�w���[��_<���b���6μ�%��Of����r��Z�1�K�
E���C�X�G�<�R�mAf�]�헚�m�V�
'�(.��+N��
l�^ف�����1���+>��̻s�mY���=���'��	��W��%��0;�fV��p�\Q���J���+��(炽�o�ܴQ�I�1��y����_��᝼�?���Oi�JzT���H��JD�n�D�\�J��8X�{�o�����@���0�ɼ0,��0���8���X���t�Ÿ́�É�m{���H���Qk�.�O���5�\"�Is�����,�%�C�\S_��y�l�g��������;���e��&G� '�M��kݼ��������G�}��<a�9�O�L�F���C��<F��nN���^�Zz��ؑ�ů��  �  a�׼Ml��<!�H)@�*^�Yw���y߆�I����u��s]��B��*���2M���O�/�цH��Ic�?�z�`ׄ�!ǆ������Xr���W��>9��������ͼ����E����bv�@�]�O�X H���F��K��%V��j�ѳ���ԛ��1����漙���k+��gJ��6g�:~�����n���<��]Rn��vT��:�Vz$�%��b�	�"�
W7�<rQ�2�k��Q��* �� ��n���j���M�R�.���r�EO��=Ԟ�v����l��W�o�K�M�F��dG�3�M�`[���r��j��Js��42ɼ�@���:�#�5��jT�x�o��с�S���IR��צ|��f�nK��2�F��r������(���?�VkZ�5os��ۂ�xǆ�{���q�y�u-a��C�ߒ$�$g��jܼ���pᕼ������d�#�R�#rI�lF�H�H��iQ��b��P}�z��"9��oj׼y`�?1!�	@��^�7Mw�����؆�铃�"�u��b]���B���*����39�'��ɐ/�	tH�8c��z��τ�H��������Mr���W��59�P��y�����ͼ�쨼�⍼);v�;�]���N�G�G��F�V�J� �U���i�=���ڽ����6��	���b+��_J��/g���}�奅��k��2;���On�HuT�N:��z$�}�'e�T�"�M[7�wwQ�b�k�OU��3$���������j�)�M���.����5켰k����V߆�_�l�r�W��K��G�Z�G�w�M�	�[��s����N���cGɼ�U��LE���5�FvT�ȳo�:؁�����FZ���|�$f�_�K��%2��2��������(��?��|Z�os�'ソtΆ����ڱy��9a��C��$��s�K�ܼ�-��V��������d�ZS�X�I�İF��I�s�Q��Xb��}��6���S���  �  m�ּ�n��:���6�U�Q�<,h��w��{��u���e�?yO��6�~� ��Z����^���Y%�?<���T�53j� x��{���t���c���K�N�0��@�_G����ͼl2��O��
���+	i�!LY��IQ�k�O���T�y�`���u�[:��}	�����P���	�ZU$��@���Y��n���y�{��xq��^��6G�P�.�����?���N�)o,��pD�){\�[�o�Y�z��z���o�PR\�� C��\'�~v��	�.z��Ϣ�?1��'Fx�A�b�КU��O��P��W���f��~~�\�����ʋɼH�"F�ӏ-�;�H��Ma��s���{��y�Fl�SaW�'�>�֔'���E�?�#���4�׮L��c�0tt�b�{��#x��7j��_T���9��5�Y�F�ڼ�T��m|���8��p�9n]���R��xO��DR���[���m��^���◼	Ѳ�.gּ�b�p/�{�6��Q�e h�w���{�j�u���e�PhO���6��� �G�M��ɷ��F%��,<���T�	#j�Ix���{���t��c�)�K�;�0�8�s6��^�ͼ� ������值��h��Y�CQ�a�O���T�J�`��nu�z"��h����I;�K�	�uL$���?���Y��n�r�y��{�uq���^�`5G���.�;�l������Q�os,�vD�]�\���o�r�z��z���o�]\�|C��h'����O%�ז���좼eO���x�*�b��U�l#P���P��X���f��~���������ɼ�%�wP�x�-�xI��Ya�*s��{�^y�7.l�esW�'�>�~�'��2�M3��R�B��	-4��L�7�c�+�t�T�{��0x�Dj��kT��9��A�@&�wۼ�q��ߚ���X���Pp���]��@S� �O�o�R�b&\��m��|��g����벼�  �  גؼ�t�����?s*��:@�R��v^���a��B\�CN��:�-%�g�V�����x�"���)�sN?���Q�wP^�� b�z\�5�N���;��i%��������;Ѽ�Y��Ť���'��JE~�r�l��c�gWa��[g�wcu�#ׅ��F��⊩���ü�伏��aT���1���F�HHW��`�]a�G`X��"H�'p3��M�A������b�~i��;1���E���V���`��a�B�X�S�H��O4�������
輛�Ƽ>��w(��q8���8w�xIh��ga��Db�Y�j��{�i��3a���v���ͼ�a𼩏���"��,9�~�L�3H[���a�u_�j�S���A�E4,�_�����ϟ�\�A?�?�"��28��;L��[��a�@_�-#T��pB��,��R��� �BܼS,�� ���D_��邼�^q�j$e���`��Gd���o�b���ʋ�������yؼu\��9���g*�4/@�PsR�Zj^�1�a�B4\��3N�`�:�x%��6C�wq��e����?�)��=?���Q�)B^�	�a�un\���N��;��`%�)��_����*Ѽ5H���������~~�/il���b�u&a�*g�F1u�>����.��Ws��|ü�
伶x�UK���1���F��AW���`��
a��\X�* H��n3�GM������e��l�f�
1���E�*�V�%�`��!a�B�X�6�H��[4�1��h��&輥�Ƽ1"��G��\W��Yvw���h�M�a��~b��%k�`�{�Ɂ��sx�������ͼ�u�ϙ�)�"��79�C�L�U[���a��-_��S��A��F,������_��[o��Q�/�"��C8��KL��[���a�1M_��/T��|B�z�,��_��� �^ܼ�I��S���/���\���q��ke�D"a��d��o�F������{;��o;���  �  �|�`��<����5.�ù:���B��)D�?�>�bu2��!�{-��e ����YG��(�=����{�%��5�e@�3qD��gA��>8�9�*�s�������$�ܼ�ż0u�����
8��a�����B�|�K�������ܗ�':��m���x�Ѽ�]�2+����.�#�N�2�1�=��C��
C�O;��H-�S �D{
�A8����缇��Ь��������v+�%�9��yB�)!D���>��4��%�u�����QUԼu���{��Kg��b���肼��|��~�֑��F���d✼�D����¼ �ټr����K	��I�6)�6�6���@�}eD��#A��
7�U�'�X���'�Q�Ho弬��B���1������0�~m=���C��C���;��/��k ��T�� ��P弌{̼趼�<��˒��芈�怼�=|��X���v���
��W�����w�ɼ�b�@G��p�������-��:�b�B�sD�0{>�Kf2���!�v��S �fy�{"��]}���V�%��5�pW@��dD��\A�58�.�*���
�������ܼ>�ļZb������Q"��N}��$�~��|�k1��;܊�R×�!!��Dm��p�ѼMH�!������#�ڝ2���=���C�4C��;�/F-�����z
��8��F��,��q���?�����|+�e�9�6�B�T*D� �>�4�Ȱ%�-����xm�(sԼ�׽��;��ц���3�����5}��S~���֎�U���\��ޜ¼��ټs����U	��S��)���6��@��rD��2A��7�D�'�.�:�2�2��$꼼����B�^ ���0�4|=���C��*C�L�;�k�/�Mx ��a��� ��m�<�̼����^��Q���h������ԇ|�}��b����,��<w��Gϴ��
ʼ�  �  ����Z��ǘ�u`��K�,Y%�MH(���&�}� �mN����Y��dܼtq˼�vƼ�9μ
�p?�����o��C�"�H�'���'�:$�����w���u��^���W�2�ͼ�x�������E��^��g����ᖼ�K���Y��nż��ؼ���ǳ��&�����!��!��&�zT(��o%�{����������Tռ�Hȼ��ǼASӼ|�PT��|�Η�	�$��6(�x'�9"�&��}��~	��R ���!�ڼ$Ǽ�6���£�����v����������� ��"P��6�˼߼!7�sg�ڋ�(x�5���#���'���'�y`#�1�o��D��Đ�D�ϼ~�Ƽ� ʼ��ټi��/����Z��5z&�P(���%� 	 ��D���z�#���1��AԼ���b`��e0�����V9���F��ȝ�#������|Ҽ/��|q���u�Ɍ��T�(@�M%�'<(���&��� ��?�$������B�ۼyN˼XSƼ�μ������o��D��\�"���'�}�'��0$�x���o����m��N��"F�O�ͼd���ᨼ�-������}���ǖ�1��9?����ļ��ؼ��{����~�%����F�!�K�&��N(�k%�˺�K������뼨Tռ�Kȼe�Ǽ�YӼ"#鼣Y������T�$�@(��'�=D"�7�����	�>a �8�H�ڼ�CǼ�V��㣼�ߗ��ڑ����)���;��Ui����˼�3߼�K�>q�x����Z��ĝ#�E�'�v�'�vn#�3@�J�g��F�㼑�ϼ�Ƽ�Dʼ��ټ{��o/���������&�R](���%�� ��Q�[��F��0���%���bԼ����j���pV��-.���_���l���일k���b����1ҼP���  �  �m��>����,��#����������������㼒ͼ ������ʩ�񓯼�ƽ���Ѽ��ԝ������d�����G�>��!���[��6��R��U�߼��ɼ�Z���2�����a������ЎռQg��� �H�	��E�X�P���C����<������F��!��=�ۼ�Ƽ�ᴼ��������_��9�ü�=ټ��ђ�����g��X���:������_��T�
�������׼y�¼>����O���a�������'ǼDݼ���P(��=�����;�����=��j��&����?d	��b ���:Լ����٣���թ�-}�����ʼ��༴p��X���V������e�o-�($�L��S�h��V��':缞�м<����ޮ�E����ԭ�pź��μͬ�0�����_��1�Q��O �:�=�����
����Z����h��̼\߹�x^��9����r��9���$�Ѽ��*������Z���/?�6�����~�kT�"��e-��?����߼�pɼ�B��K�������E��^����sռ�L�� ��	��:�eM��y��:���m���:����������ۼ�Ƽ<ⴼq"��,���Ff����üBHټN#�1��,�7�������%G�B���������
���~�ؼ��¼񻲼�o��R�������7CǼ� ݼ��/3�H�"���D�(��2G��t��1�� ��q	�`q ��-뼛ZԼqƿ��ư��������.<���ʼ7��������Zd�@����r��:�2� �����-z��W_�M�м�ϼ����v���h����뺼@Cμz�伛"���,��  �  �+'�U9(�O%����o�������4���ϓ��Ѽ¤��򳫼=������e�����a��iw�����)wռ���:�������;���u ��&��_(��F&�]��0�._��u�k�ؼ�ɼ��Ƽ��м��~����?�b����#��(���'�F#��Y�p�������:2�޼	{ʼgS���P��o���T���񑼻R��F���D���Dȼ��ۼ��� �3
�9��~m�d�"��5'��"(�p$����k��׀����pQҼd5Ǽ3�ȼWQּDf���7��uF�g�%�_W(�	~&��-!�������{�����Y�׼��ü�H���n��[R��le���N��)͛�#é��k����μT��S�������`��]��x$��(��v'�Y%"�rB���s���ݣ߼hRͼ^?Ƽy�˼�&ݼ�m��ف	����B!�T'�,(��%�����������i���y�e�мՇ�����������E���t���IZ������%^ռ@�����������о��n ��&�^X(�?&��T�~'��T��^�ؼ��ɼ>�Ƽ��м���T����1���&�#���'���'�<#��P�m������v(��	޼kuʼ�O��fO���o��XW��@���nY������N���Qȼ��ۼ�（� ��
����y�Ȝ"�D'��1(��$�:� ��Ǒ�����rҼVǼ��ȼ'oּ*������MQ�d�%��`(��&��6!�ʲ�?�6����=�꼨�׼4ļ�g�� ����s�����Qp��%4㩼����.�μrp�2o����������7�$� (�ֆ'��6"��T�7)�Ұ��T�߼f|ͼFiƼ�̼�Nݼ���֓	����,R!��  �  �DD�u`B�� :��=-������w���	���ȼĵ��j���kk�����:����|�V��H<��%|���R���$��l�ͼ���̪��C�"X!��d0�:l<�aC��C���<�m�/���PL��[��j�N�开>����	���(�I�7�t�A�eD��=@��96��@(��g�.q��󼳁ؼ�Z���B���������.����}�$M}��X���Ì�/K���*���ڶռ���R��s��I�&�4�4�U?��5D�T'B�o9��*����u��h���C�G�v}���`�j��.'.�y�;��DC���C��s=���1�2#����N���Qgм=P��+��4����F���ہ�T|�HG�����}֐������o���-ƼF޼�d��K��M��e�+��8���A��XD���?���4���$�!�ê�T�P
�6F�Y�����"�s43���>��5D��RB�A:��1-����,��(�����༞�ȼ,����j��UN����������R|� 8��D���`���8����>�ͼ���i��I<�;Q!�,^0��e<�(ZC���C�U�<���/����@��B���N�
��!�A�(��~�(���7�x~A�SYD��2@�a/6�m7(�_�j�{�wؼS���<����:��/���}�uV}��_���̌�V��t7��������ռ��������&���4��c?�ED�d7B�09�,�*�����[���
e�f7�ۛ��o�w�3.�I�;�eNC���C��|=�]�1��#����X����+м1j���F������e��y���	�|���������������򌱼JƼ,޼|�������y�+���8�M�A��iD���?�!�4���$��Q���6��5��p�+�D&�'�"��E3��?��  �  S	b�^�˟Q��?��1)���Z>��w�ּ黸����<Ŏ��	���o�#%d�'a��e���r������l���ӥ�nԾ��F޼f�.���2.�ŖC�M�T��_�V�a�'oZ�(FK��7�}�!�rp��X���U	����~t-���B�A�T�4�_�˰a��Z��K���7�D�!�Da�O�˼���FX��Y���~�z��Sj�4b�ʬa���h��ax�����7���^���rȼ��I�����5���I�xYY��Ja�4.`��V���D���/����Ц
� ��9����_d�
�4��+I��Y�Ea�4P`���V�ǾE���0����W�	⼦����7���;��|	��J;t��f�a�?0c�|+m�VP��ꌼ���q�����ҼT���1-���&�Ӷ<���O���\�]�a�R�]��Q�>�̟(����@��`c���5���D&��;��&O�w�\�F�a�=�]���Q��	?�&)����O'����ּ4�������+����퀼��n���c���`���e�%Tr�d���6T������~����4޼��*��8,.���C��T�M�_��a��fZ��<K��7���!�yc�*������F	�����e-���B�={T��~_�S�a���Z���K�<�7��!�Z��B�˼���qR������H�z��Tj�[!b��a�:i�:sx�����D���m����ȼ
-�	�W�ؓ5�`�I�5hY�'Za��>`��%V�3�D�h�/���P�
�1��I�*���r�9�4��7I�lY��Na�*Y`��V��E��0�Q�a��/�f ¼�P���V���%���vt���f��La��nc��im�,��!���Ȟ�=ϵ��Ӽ&����:�m�&�3�<�2�O��]��b���]��Q��'>�{�(��������y�)����8Y&�B�;��8O���\��  �  ��{��v��g��;P�U5���� ��HԼ�3��M���������l�g[�;2R��O��S��|^�0�q�J���훼�:���Mݼ������z;�b�U��Ck�^�x���{��s���b��]K��2�������5W�L��b�(�JW@�!�X�m��zy��]{��`r��`��G��,�{��;��<�Ǽ%g��܉����|�G�e��XW�OP�I$P��6V���c���y�2L���Q��^vü&��)����(�<D���]���p��z�+z�t�n�73[�]C�<++��p���g������40�T�H�/%`�g@r�'O{�X�y��-m�"qX���>���"�pB�X��"ӻ�/����'���t�o�_��<T�آO��_Q��Y�j�i����(��Z���C�ϼ�����k12�TM�X�d��8u�<�{���w��i�~mS�B�:�$$�0�������X�!�!8���P���f�9ev���{�|v��
g��/P��I5����= �~1ԼK������{���Wl��.[�p�Q���O�rhS�@G^��fq��2��K؛��'���<ݼU|�)���s;�z�U�w=k�ңx�A�{��s��b�SK���2�T��t��qH� ���(�H@�I�X��m�omy��P{��Tr��`�s{G� ,�������|Ǽ_��󃏼�|���e��YW�q�P��-P�DV�M�c���y�DY���`����ü��������(�-�D���]���p���z��;z���n��D[�MC�6=+����;����d�C0���H�01`�-Kr��X{�*�y�6m�"yX���>�H�"��K�Q��黼����A���Mt�D/`��xT���O�ޜQ��Z�8j�؁�E���ڭ�V�ϼ�������a?2��bM���d�:Iu��{���w��-i�؂S�|�:��:$�I$�������3
"��-8��P�g��uv��  �  ᆽ���#v�Ӊ\��o>�c�����ռ�r���ܑ�F�{��'a�g�P���H�òF��J�V�S��f�����j���"���߼����O&��OE�þb���z�$����"���:r�{�X��N>�~�'�Yd�3��f���i3�n�L�N�g�p�}�����~��7g��rRn���R��4�|���v����Ƽ�ʣ�B���_q���Z�(NM�$NG� G��JL�p�X��:n��臼�t���}¼���jX�U�0�riO�}k�'w��50������Ψ�m;j�v�O���5��!���(n� q%�tp;�i�U��o���������n����|��e�S�H�в)�y�F+����D��𗃼"�h��+U��J�<�F��H��}O�̪^���w�
$��󰪼'мY���+���:��JY�q�s����ĕ�2���_y���a��F��U.�b��M(�ߍ���+�QD���^�+w��能Fن����v��}\�d>��������Լ�Z���Ñ�<{���`�L�P��H�U{F�S�I�4�S�p�e�B���sU��J��\�޼����I&��IE��b���z��q����z���0r���X��B>�0�'�V�C��
��Z3�
�L�Fxg���}�9���`x��Ia���Gn�C�R�e 4����i��C�Ƽ�£�<���Wq�d�Z�OM�BSG�c	G�+XL�/�X��Pn����� ���C�¼d��Jc�K�0�xvO�'�k��~��+8�����)��BMj���O��	6��!�0#��~�Ȁ%�;���U��o����Տ��Ms�� }���e�9�H��)�`��>�,��\��;����h��dU���J�"�F��IH���O���^�U'x�+@��n̪�&BмG����8���:�vYY��s�	
��jՆ�ݏ���sy�y�a��G��l.�����?�Ϥ�,�nD���^��#w�B��  �  ht��꽧�۽�iŽ,���Z���o���D���"�	���N�ּG�Ǽ|
��Fｼ�D����ʼ�qۼM���	x�y�)�pM�/�y�N7���(����ʽ�߽��6����`ؽV½C)��ꓗ�wz��-����+����㷽�Ͻ�p�7*�_������Խ�鼽o#������`��u8����9��\��g�м�ļ����V����ü5ϼ���ơ �R���4�44[�B&������#�ҽ�F彯Hｱ���$�2jѽ	v��������������P����ƕ�Ⲩ�o����ֽ�V罃��a����vͽ����*����~��Q�W.-��z}����ݼb�˼5���뽼k��]�Ƽ��Լ4��`����O@���i��o��$��1�½��ٽV���V�bY�1�޽8ʽ8����g���v������zV��v]��$!��yǽR�ܽ�E뽅l� ��8�۽�cŽ~&��mU���o�d�D��"�_v	����5�ּc�Ǽ5ӽ�\)��-�ʼ	Yۼ�����m���)��hM�ُy��4��l&����ʽ��߽��2���5\ؽzP½�"��،���r���$���������z۷�~�ν�h��"�f��d��C�Խw伽�������`�>p8�@|���C�弎�мv�ļ�����Z����üM>ϼ
�⼢� �Q��<�4��>[��~#�������ҽ�N�7Qｪ��+.��sѽ���l��'������9����Ε�����D����"ֽ7\���Z��J��tyͽ�"��X.����~�+�Q��8-�~�������ݼ
̼�����	��������Ƽ��Լ;��v,�s����@�j��v��+����½ �ٽ��?`�c�(�޽�ʽ`���t��s���3͈��b��]i��h,����ǽ��ܽ}N��  �  �$�彌;׽�����V���{���m�4D��r#���
�Y/�G2ڼa	˼��¼>���"/ļ��ͼ&�޼�������j*�ӜL��;w�G"�����O�ƽv/۽h����꽏��:�ӽ�K���ʧ���l��������u��*����'��E�ʽ�uݽ�轴}�b���н�q��֠��N/��J�^�_T8�$R�����S/Լ��Ǽ:{��+����ƼscҼO.����u���4�9�Y��v��"�������UEν^�z��4��X߽��̽x���UР��؏�����7����Hf��۽���}ѽ58�k��5��wݽ\gɽ����`���tb|���P��h-�D�=x��m�!ϼC�ļ����EH¼%�ɼ! ؼ���7h��C �Q@�&h����1j��x��ս;�佫 �罔�ٽ[�ŽN���l���勽W��F͊�.q��
���JHý��׽�
�C���!5׽����Q��v���m��(D��f#���
�/� ڼI�ʼD�¼գ��Zļ�ͼ:�޼����W����)�:�L�E5w��������ƽ -۽��罂�꽓��x�ӽfF��}ħ�ջ������ȸ���m������I���ʽ nݽ����v����M�н�l��@���V+����^��N8��M������}-Լa�Ǽ�}���/����Ƽ�lҼ�9漼��}�ė4���Y��|��v��������Lνf���&�齥&߽#�̽0���ڠ��⏽>!��z@��i
���m���Ļ��ѽq=����4��ݽ�jɽ{�������j|���P�Xs-��#��������=ϼA�ļG���g¼��ɼؼ��Vv��Q ��'@�w3h�ӱ��8q�������ս��
�G!�z�ٽ��Žc$��y��K򋽢c���ي�}��?����RýI�׽���  �  �ܽ�׽ȃʽGA��⭠�6���=nh��C���%��K[���y�%�ԼR̼*�ɼWeͼ"�׼p	�3w�ю���+��:K�\|q�Ʀ��:ԥ��컽�	ν�Tٽ��۽�սtƽ�ٲ�j8������2遽A�����ԕ������#���iϽ��ٽ.�۽�
Խ��Ľ_�D蘽a1���d[�D�8����K���S�fN޼B Ѽyʼ�!ʼ'�ϼrܼM�������z5� /W�ׄ�uM��yj����½��ҽ�)۽{�ڽJ�н�A���׫�З�8��Y(��{1��z ��������foĽ��ӽҁ۽�ڽ)�Ͻ|-��J`��#0��ev�)O���.�'��W'�Q]��
ټ�μJ�ɼ�W˼,OӼ�;⼂$��!����"���?���c�(�����QԴ�ÚȽ8sֽ�ܽTHؽ�̽�����ꤽ�����
�~�⒃�Z��餢��j��8;ʽP׽5ܽ�׽j}ʽa;��G�������-ch���C���%�m���@��^�t�Լ,�˼�ɼ�Hͼ�{׼���nk�F��u�+��2K��uq�ݣ���ѥ�껽ν�Qٽ��۽�սRoƽQԲ�!2�������ၽb���醽}̕�q������#bϽ?�ٽT�۽mԽĝĽ:믽�㘽s-��H^[���8�d}�$���O�L޼� Ѽ�{ʼ�&ʼ(�ϼ8{ܼ���l����܃5�@9W�A���S��Uq���½�ҽ�1۽W�ڽ�нK��"᫽�ٗ��A���1��C:���(��c��߈��euĽ��ӽf�۽�ڽޭϽ1���c��4���v��'O��/���Z4�Ly�S(ټx3μ��ɼ9w˼/nӼ�Y��A��]���#��?��d�������۴���Ƚ�{ֽ�ܽQRؽf̽����m������������������*��揤�t���Dʽ�X׽�  �  ?(ƽX�½ya��iѨ�����Ã�o|d���E��r,�����������m�{�ܼ^�ټ�޼��鼧W��z0�m&���1�(AL�5�k�)���G�������7��.2Ľ��Ž�����ಽ-ա��鏽������n���j�Nw�Z���������x����ĽW�Ž������`䢽n6��l{�=�Y���<�k%�+��t����#?���ڼ�]ڼ���
��Q�K�"�b�9�e5V�ow�����נ��뱽�羽�Ž��ĽK��Mz��ٽ���V��.�y�:sk�hBm�\�~� ���˟����f���.�Ž��Ľ񄼽oj��.Ü��q�o�
O�Q4�B��������A8��޼'�ټq�ۼ��伳+��o_����)�0�B���`������f���٦�#ֶ�����#ƽ��½Ǽ���§�����;��-s�y<j�=jq���������p˥�c+������� ƽu�½/[���˨�|���l���Aqd�
�E��f,����)���o���O�Inܼ'�ټ�޼ ���<��$�M��1��8L���k�݇�w���ޕ��c4��2/Ľ��Ž�����۲��ϡ��㏽����>vn�N�j�>w�@���ﺙ����謺��Ľ��Ž����睳�Sߢ��1��Xd{���Y���<�/%�d(��r����?�h�ڼdbڼ�%��n��X�3�"�k�9��?V�]zw�����ޠ�󱽡ﾽa�Žc�Ľ[������KǛ�`��֗y�V�k��Sm���~�u��Sҟ��#������чŽ��Ľǈ��(n���Ɯ���l�o��O�C\4�lN�f�������V뼼߼W�ټ��ۼ{�伳J��kn�v���)���B���`�/���~m���ঽ�ݶ�=���,ƽ��½1Ƿ��ͧ��ŕ�hG��Es�xTj�q�װ���˓�xե��4������  �  P��m�������ᙽ����j���e�o�N��:�/�'��$���
��� ������[�=�����l��4r���+�l>���S�pdk�B�������w���ی���]��c���z⦽����#�����}�͡d���T��Q��B\�ѻq�C���畽Ȕ���ɪ�n6�������`��н������?�v�:�]��{G��3�3]"�e��.��������6�h���!���� ���1�"E��1[���s�����L���/�������NR��b����n��̰��ݑt� ^��kR���S��Ib��z�~���z��L⥽6A��$���:l���ĝ��p�����3&n�EV��@�7�-������������ e������ ��	�{��%���7�%4L��#c�r|�
����P���	���=-��li��,����䵃�ul���X��iQ�/^W�9~i����w������n���������蚤�(ܙ� ���_�K�e���N�Z:���'�`��
�� ����6<�������1��e��+��a>���S�~\k�ͣ�����������Z��ؙ��cަ�/񛽺���_�}�t�d���T���Q�3\��q�t���ߕ�o����ª��/������?[��ḕ�b�����v���]��vG��3�(Z"�c�.� ���7���
o�������g� ���1� +E��;[��s���pS���6���������Z��B����w�����X�t�;(^�F}R���S��Yb���z�!��π���祽�E��h���:p��sȝ�	u��#���/n��!V��@�R�-��$������������3���� ���	�m���&��7��AL��0c�3|�����������5���r��3������ ���Y5l�*�X�ӀQ��tW��i���,���Þ������  �  ;���c������F���[�������p�y]a��FQ��@�k0�� ��5�pH���	�	������#���3�gdD���T���d��Tt�Դ���爽GB��瓽�ƕ�����&��Ȅ�.br��Z��F�#G:���7�8
@��Q���g����`]��_���Pw���"��˖��Jދ�����{���k��	\���K�2;�Ұ*���f��F�
�{
����d��|�(�m-9��I��:Z�\ j�]Vy�� ��������vڔ�s���}q���V��S���@j��JS��xA��>8��n9��D�X�o�o�L���N@��
��������@��Tݏ�æ��W���s�u���f��V�Q2F��|5���%����E��
�]�� �v��5.���>�fO��_��*o��b~�D����B����������* ������.5���Sz�$Kb�ݖL�!P=��r7�s(<��J��_���w���������ӡ���������wU��'��/�p�XQa�	:Q��@��0�O� �b%��7�+�	���������#�l�3��WD�+�T���d��Kt����L䈽?���㓽�Õ�o����"��SÄ��Wr�=�Z��F�;9:���7�3�?���P���g���EV���ّ��p�����u���~ً�����l{���k�n\���K�8
;��*��������
�w}
�����(�49���I��CZ�L
j�bay��&��%���
��┽m����y���_��4���Rj��\S���A��O8�S9���D��*X���o�6����E��Շ��3ƕ�(E��}ᏽ��������v��f�ĶV�=@F���5��%����+W�c
�ļ�	���UE.�{�>�HtO���_��7o��o~�Б��zI��ޝ��_���x�������>���gz�e`b�¬L�Uf=�
�7�0><��J��_�H�w�����ʏ��  �  G(��?��䓆�e���[���q|��e��Z��x6s�3�b���O���<���,��8"��\�#�� 0�]A��?T��f��\v�{���侄��ӆ�H����s��G/�������}�Ŷp���_���L���9�l�*�R"!�VW�\�%�ی2��)D�oW�W�i�<�x�F���0���������!P��mօ�%߂���{��n��\�xsI�b7�(�S? ����%9'��45��LG���Z��Jl�c�z�.j��A���/0��+���� ���o���-���y��\k��{Y�x5F��C4�/�&�N���z �")� 8�րJ���]�4�n���|���:��Z��,�����F���x����w�F�h��SV��C��1�|�$�A,�}i!��<+�@�:���M��`�؂q��~�����D��#x��$���R���!���󮀽o�u�D�e��S�%�?�/�$m#�@��n�"���-���=�\�P���c��s�T!���8����������ш���v�������)s���b�(�O�`�<�{�,�"'"�O���#���/�'�@��0T�P�f�%Pv�������Qφ�����qp���+��|��Z�}�^�p�Y�_�(�L��9�Ѕ*��!�AI��t%�<~2�D��`W���i�5�x�*���q*�����S����K���҅�܂���{��n�&�\��qI��7�J(��@ �A���<'�95�\RG�4�Z��Rl�$�z�o������!6�������'���v��v5��c�y�ymk��Y��FF�NU4�m�&���� �>1)�*8�čJ���]�� o�[�|��������A_��ʬ����������~��"�w��h��cV��!C�Ҳ1���$��>��{!��N+�J�:���M�X�`�7�q�y�~�����K���~������7���~���඀��u���e�I.S�a@��./�K�#�_�-�"���-���=�?Q�|�c�:t��  �  �>b�d�q�7w��-���?K���K��k���鏔�Uf������Tjv��x^���I��;�Ɣ7��>��M�ׯc���{�ʈ��䐽	)���r���^�����+��d�}�Zn��^��N���=�g]-��W����y��'
����#���h&�nr6�D(G�Q�W�Mtg�t�v��킽I��j+��m�������E���̌�$�jSn���V���C�P9�!�8�}KB�l�T���k�����<׋����⥕�ӷ��绐�����<����|x�? i��QY�~�H�z:8�V(�j�����P
���
��l������+���;�~�L���\�(�l���{�Z���7��ؑ�<<���[��f���JӉ��B~��Cf���O�-F?�X�7���:�F�G���[���s� Z�����})��/���(����뎽���{E���ns���c�R�S�gfC�`�2��#�9���(���	�M��ɹ�%j!���0��A��!R�1b���q�iq�������E��F��{�������n_��9���<Zv��g^���I�e�;��7���=���M���c�]�{���7ސ�#���m��2Z���댽H'���}��Rn��^��~N���=�S-��L��x��l��
�ɫ����Z&��d6�G���W�~hg���v��肽���e'���i������}C���ʌ������Qn�"�V�;�C��9���8��NB��T�+�k�ݳ��ۋ�f�������-�������Ǌ�����x�y/i��aY��I�LK8�Y(�i��ɔ��`
�b
�k{�S��l�+�s<�<�L���\���l�'�{�(_���<��aݑ�B��ab������'ۉ��S~��Uf���O�QY?���7���:���G�I�[�>�s��a��e���N0���ĕ�g���,�f���L���|s� d��T��wC���2�#��"=���	������`|!���0���A��0R��  �  ��O�*Bg�Nq���ʍ�׌��� ���«�j���f>������>��.N��Mh���V��Q�u�Y�F�m�M���}��������ϩ�G=��̶�����Kח��ӊ�F{���a�GK���6��%����?	�<M�����
��s}���f�p�����H�.���A��aW���o�ބ�x+���d���ا� Ϭ����_��_����9���y��8a���S�<�R�Q_�Cv�2����7��dI�������������엟�M���7T���Wr�n�Y�+�C�8�0�������m�s���0��F��[�������#�@#�ڻ4���H��%_��x��R��Ho��K����8��*u��e���B��2���@p��M[���Q��xU���e�YU���������fT�����)�����؛�I>���䁽,�i��PR��C=��*�ċ�����M����,����KZ�Z��4����(��;���O�6g��k��Gō�X���B��߼������K7�����`6��@E��@:h�"�V�A|Q���Y�*{m�(����{������_ȩ��6��2����	���җ�xϊ�� {���a�;K��6�y%������\5���}�����b��Y���f����.�[�A�VW���o�%ل�'���`���է�6̬����^������9��y��8a��S���R��!_��v�񍉽);��)M�����v���������������Z��fr�U�Y��D�E�0���a-�F~����������U���*���0��K#���4��H�c/_�j$x�iW��vt��������m?���|������.���;���Tp��a[��Q�S�U���e��g�)��������[���ì��/�����ޛ�eD��끽�j�M_R�vS=�m�*�J��1���`��?��fS�C���l�њ�����(��#;��  �  8uG�rTf��Ʉ�8����Ʃ�h���.ý�ƽ�<��Me��#פ��В�e낽�p��fj��6t�����Ö�Oƨ�A�����½W#ƽ������5䥽�_�������	_�GGA���(�	����+��n@伣�ۼ(ڼT�߼3�Q �6��;b�8�5��,Q�V�q�J���̝�+Q���&����Ľ�SŽ�����<���˞����)L}�g�l���k���z��@���Ĝ�\j��)���}�ĽahŽ�V������ӟ�����xu��}T�>r8�Ə!�pg�?V�F��p�B'ڼ��ڼ�⼂��'��c>&��A>�As[�f}�>A���⣽�s�������Ž��ý����੪�;�������Z)v�A�j�Z o�hd��7א�"Ϣ����y4��l�Ž�ý.���u���գ���҆��j���J�H0��	�fN
�����_�輼�ݼ7�ټL�ܼ缔���9��{��*�-��hG��Hf�)Ą�ǌ��S������v(ýQƽa5��V]��~Τ�Mǒ��Ⴝ��p�]Rj�v"t����8���M���򀸽&�½�ƽ }������ߥ�@[��}����_�	?A���(���������)�zۼ��ټ)g߼��6 �_���U�e�5��!Q���q������ǝ�WM���#����Ľ�QŽ��*;��˞�2���L}���l��k�>�z��B���ǜ��m��綼���ĽmŽ\��z���ٟ�;����u�%�T�|�8��!�~w�vf������^Fڼ�ۼ���L�34�""�?I&��K>�*}[��o}�UF��%製�y��e���� ƽy�ý���1���Ę��ć�)>v��j��4o�Dn�������ע�5����;��J�Ž{�ý<���[���©���؆��j�[�J��V0���0_
������輛�ݼ�ټ��ܼR2�6�����?�Һ-��  �  x�E���j�Y܊�h���yp��#m˽6ؽGܽ��ֽ1Wɽ(P��	���KH��f'���� ,���풽��L׺�o�̽��ؽ�۽D�ս��ǽ裳�+̜������a�x.>���!�-�������K���Ҽ�.˼��ɼ3�μ��ټ)�켼�|"���0� Q��qx��x�������J���sнqaڽQ۽�ӽFlýS[������b���耽Ad���툽�ܘ����	U��l�ѽU�ڽ��ڽe�ѽNt��?)����� }��U���3�ߑ����K)���ۼ%gϼ��ɼ��ʼ��Ѽ�8߼B�����	������:��]�.g��1���*���Ž�Խ��۽�ٽu�ν����^���ϔ��J���]�#C�������J�������gǽ9�սX�۽�ؽ+ͽW���Æ��]��'o�NAI��O*�
X�� �j��Ŷּ��̼V�ɼ�5̼sHռ�t弳�����qO'�vE�s�j��֊��k��ig˽ؽ�
ܽF�ֽOɽLG������C>�� �����!��7㒽+���ͺ���̽�ؽ	�۽�ս�ǽ����ǜ��ۅ�z�a�&>���!����z���]6�ȱҼ\˼üɼ�μ6�ټ���0�[�m�0�9Q�sgx��s��n����F��spн�^ڽ�N۽�ӽ�jý~Z��b���0b���逽se��b�ޘ����BX��$�ѽ��ڽQ�ڽ��ѽ�y��Q/��c
���-}��,U���3�Z��c��-I�Σۼ��ϼ�ʼ�ʼ�ѼS߼���,�	�����:��]�<l��S6��^0����Ž��Խw�۽+�ٽk�νJ���h��|ڔ��U��&s��M������-T������oǽ��ս:�۽x�ؽ1ͽ!Ǻ�����c���3o��NI��]*�\g�K� �l����ּ�ͼ�ɼ"Y̼�jռw�弁���	#��\'��  �  �DF���o�:㏽1ɩ�z�½MAؽ�l��뽎��X�ֽ>½Jn��i����W��)o��䈌��}���c��{ǽ��ڽ���p���佱Խ��������N��	�e�d(>�����V��s��׼�4ɼ|#¼����LżQ�ϼ�S�"c��n�//��)S� �j���e����ʽ��ݽ��TV�~��bн�{���?���2��臽�X�����������νS�߽���8��ڑ߽ͽ�6���D��g ����W���2����D�伉~Ѽ�	Ƽ^��������ȼ�ռ�d�-$�����9:���`�"�������Һ��ѽ��o��tr�ҍܽ�eɽ�ܲ������������`�����I�������b�Խ�@�.���j�X6ڽ��Žk��������t��mJ�I(��I�]��hݼ��̼{�ü�����ü��˼�(ۼE����q %��8F�T�o��ݏ��é��½�;ؽaf���z��ֽ?
½�d��3|��,M��_d��~��]s��|Y����ƽ��ڽ���?��}�Խ����E����I����e��>�ƾ��M��_�W׼ɼ�¼����2ż��ϼJ:�gJ��!b��#/�(S���~��e��pa����ʽl�ݽ	�T�H|ὓaн{��X?���2��/釽�Y��̟��������.ν�߽�������߽�ͽ�<��NK��8'���W���2�l�)�����Ѽ�(Ƽ���3����ȼ;,ռ_}��/����,D:��`�C������:غ�F�ѽ������z���ܽ`oɽ�沽x���̍�����Ik��O�������������ԽnH���6q�H<ڽR�Ž���w���d�t��zJ�$W(��X�&9��a�ݼͼw�üû��j7ü0�˼�Hۼ������%��  �  ��F�5�q��ϑ�`���8�ƽ�ܽ�뽴q�[��E�۽i:ƽ$讽�k��j݌�و�J��v������Q˽u�߽\��,H�齘{ؽ�6��⨦����4{g�|>������F��Ӽ�+Ƽ�G��c��'Z¼��̼߼p���j��/�G8T�NӀ����������νS���W�i��^��%�Խ�h������8��\��ɉ�Q��G'��Uɻ���ҽ���	'�Xｵr佇Eѽ����+��������X���2���~7���ἻRμrü�*��wž��ļ��Ѽ�0�������k:��{b��'���dW���$ֽ���[������ὧ�ͽ��������_��C����ߋ��w���]��w�ýPsٽ�n齗L𽛘���޽|ɽ���.�����v��-K���'�^$��	��#)ڼ��ɼ����3Ƚ��1���yȼ�׼�𼟩
���$���F�ئq�rʑ������ƽY�ܽ؉��j�Ѱ���۽^1ƽlޮ�ia���Ҍ�3Έ�p���u������BH˽��߽B���@�L��uؽw1��D���z���rg��s>���L���2꼳�Ӽ:Ƽ0������
A¼R�̼��޼qW���^���.��-T�R΀�j���z���b�ν��U��ｎ����Խ�g��:���g񔽝]��Lʉ��R��|)��
̻�Ѣҽ��9+���w�Kѽ��������ꑃ��X�~�2�/��V�����rμg1ü�H���⾼�ż:�Ѽ�I缌����v:�(�b��,��K���!]��+ֽx��
 �t���Ὁ�ͽ}�������~j��2
��Pꋽꁘ�rg����ý�{ٽTv�|S�����޽ʁɽ����������v��:K���'�@3�K)��1Jڼ��ɼ�����꽼T��	�ȼ�
ؼ�𼪷
���$��  �  �DF���o�:㏽1ɩ�z�½MAؽ�l��뽎��X�ֽ>½Jn��i����W��)o��䈌��}���c��{ǽ��ڽ���p���佱Խ��������N��	�e�d(>�����V��s��׼�4ɼ|#¼����LżQ�ϼ�S�"c��n�//��)S� �j���e����ʽ��ݽ��TV�~��bн�{���?���2��臽�X�����������νS�߽���8��ڑ߽ͽ�6���D��g ����W���2����D�伉~Ѽ�	Ƽ^��������ȼ�ռ�d�-$�����9:���`�"�������Һ��ѽ��o��tr�ҍܽ�eɽ�ܲ������������`�����I�������b�Խ�@�.���j�X6ڽ��Žk��������t��mJ�I(��I�]��hݼ��̼{�ü�����ü��˼�(ۼE����q %��8F�T�o��ݏ��é��½�;ؽaf���z��ֽ?
½�d��3|��,M��_d��~��]s��|Y����ƽ��ڽ���?��}�Խ����E����I����e��>�ƾ��M��_�W׼ɼ�¼����2ż��ϼJ:�gJ��!b��#/�(S���~��e��pa����ʽl�ݽ	�T�H|ὓaн{��X?���2��/釽�Y��̟��������.ν�߽�������߽�ͽ�<��NK��8'���W���2�l�)�����Ѽ�(Ƽ���3����ȼ;,ռ_}��/����,D:��`�C������:غ�F�ѽ������z���ܽ`oɽ�沽x���̍�����Ik��O�������������ԽnH���6q�H<ڽR�Ž���w���d�t��zJ�$W(��X�&9��a�ݼͼw�üû��j7ü0�˼�Hۼ������%��  �  x�E���j�Y܊�h���yp��#m˽6ؽGܽ��ֽ1Wɽ(P��	���KH��f'���� ,���풽��L׺�o�̽��ؽ�۽D�ս��ǽ裳�+̜������a�x.>���!�-�������K���Ҽ�.˼��ɼ3�μ��ټ)�켼�|"���0� Q��qx��x�������J���sнqaڽQ۽�ӽFlýS[������b���耽Ad���툽�ܘ����	U��l�ѽU�ڽ��ڽe�ѽNt��?)����� }��U���3�ߑ����K)���ۼ%gϼ��ɼ��ʼ��Ѽ�8߼B�����	������:��]�.g��1���*���Ž�Խ��۽�ٽu�ν����^���ϔ��J���]�#C�������J�������gǽ9�սX�۽�ؽ+ͽW���Æ��]��'o�NAI��O*�
X�� �j��Ŷּ��̼V�ɼ�5̼sHռ�t弳�����qO'�vE�s�j��֊��k��ig˽ؽ�
ܽF�ֽOɽLG������C>�� �����!��7㒽+���ͺ���̽�ؽ	�۽�ս�ǽ����ǜ��ۅ�z�a�&>���!����z���]6�ȱҼ\˼üɼ�μ6�ټ���0�[�m�0�9Q�sgx��s��n����F��spн�^ڽ�N۽�ӽ�jý~Z��b���0b���逽se��b�ޘ����BX��$�ѽ��ڽQ�ڽ��ѽ�y��Q/��c
���-}��,U���3�Z��c��-I�Σۼ��ϼ�ʼ�ʼ�ѼS߼���,�	�����:��]�<l��S6��^0����Ž��Խw�۽+�ٽk�νJ���h��|ڔ��U��&s��M������-T������oǽ��ս:�۽x�ؽ1ͽ!Ǻ�����c���3o��NI��]*�\g�K� �l����ּ�ͼ�ɼ"Y̼�jռw�弁���	#��\'��  �  8uG�rTf��Ʉ�8����Ʃ�h���.ý�ƽ�<��Me��#פ��В�e낽�p��fj��6t�����Ö�Oƨ�A�����½W#ƽ������5䥽�_�������	_�GGA���(�	����+��n@伣�ۼ(ڼT�߼3�Q �6��;b�8�5��,Q�V�q�J���̝�+Q���&����Ľ�SŽ�����<���˞����)L}�g�l���k���z��@���Ĝ�\j��)���}�ĽahŽ�V������ӟ�����xu��}T�>r8�Ə!�pg�?V�F��p�B'ڼ��ڼ�⼂��'��c>&��A>�As[�f}�>A���⣽�s�������Ž��ý����੪�;�������Z)v�A�j�Z o�hd��7א�"Ϣ����y4��l�Ž�ý.���u���գ���҆��j���J�H0��	�fN
�����_�輼�ݼ7�ټL�ܼ缔���9��{��*�-��hG��Hf�)Ą�ǌ��S������v(ýQƽa5��V]��~Τ�Mǒ��Ⴝ��p�]Rj�v"t����8���M���򀸽&�½�ƽ }������ߥ�@[��}����_�	?A���(���������)�zۼ��ټ)g߼��6 �_���U�e�5��!Q���q������ǝ�WM���#����Ľ�QŽ��*;��˞�2���L}���l��k�>�z��B���ǜ��m��綼���ĽmŽ\��z���ٟ�;����u�%�T�|�8��!�~w�vf������^Fڼ�ۼ���L�34�""�?I&��K>�*}[��o}�UF��%製�y��e���� ƽy�ý���1���Ę��ć�)>v��j��4o�Dn�������ע�5����;��J�Ž{�ý<���[���©���؆��j�[�J��V0���0_
������輛�ݼ�ټ��ܼR2�6�����?�Һ-��  �  ��O�*Bg�Nq���ʍ�׌��� ���«�j���f>������>��.N��Mh���V��Q�u�Y�F�m�M���}��������ϩ�G=��̶�����Kח��ӊ�F{���a�GK���6��%����?	�<M�����
��s}���f�p�����H�.���A��aW���o�ބ�x+���d���ا� Ϭ����_��_����9���y��8a���S�<�R�Q_�Cv�2����7��dI�������������엟�M���7T���Wr�n�Y�+�C�8�0�������m�s���0��F��[�������#�@#�ڻ4���H��%_��x��R��Ho��K����8��*u��e���B��2���@p��M[���Q��xU���e�YU���������fT�����)�����؛�I>���䁽,�i��PR��C=��*�ċ�����M����,����KZ�Z��4����(��;���O�6g��k��Gō�X���B��߼������K7�����`6��@E��@:h�"�V�A|Q���Y�*{m�(����{������_ȩ��6��2����	���җ�xϊ�� {���a�;K��6�y%������\5���}�����b��Y���f����.�[�A�VW���o�%ل�'���`���է�6̬����^������9��y��8a��S���R��!_��v�񍉽);��)M�����v���������������Z��fr�U�Y��D�E�0���a-�F~����������U���*���0��K#���4��H�c/_�j$x�iW��vt��������m?���|������.���;���Tp��a[��Q�S�U���e��g�)��������[���ì��/�����ޛ�eD��끽�j�M_R�vS=�m�*�J��1���`��?��fS�C���l�њ�����(��#;��  �  �>b�d�q�7w��-���?K���K��k���鏔�Uf������Tjv��x^���I��;�Ɣ7��>��M�ׯc���{�ʈ��䐽	)���r���^�����+��d�}�Zn��^��N���=�g]-��W����y��'
����#���h&�nr6�D(G�Q�W�Mtg�t�v��킽I��j+��m�������E���̌�$�jSn���V���C�P9�!�8�}KB�l�T���k�����<׋����⥕�ӷ��绐�����<����|x�? i��QY�~�H�z:8�V(�j�����P
���
��l������+���;�~�L���\�(�l���{�Z���7��ؑ�<<���[��f���JӉ��B~��Cf���O�-F?�X�7���:�F�G���[���s� Z�����})��/���(����뎽���{E���ns���c�R�S�gfC�`�2��#�9���(���	�M��ɹ�%j!���0��A��!R�1b���q�iq�������E��F��{�������n_��9���<Zv��g^���I�e�;��7���=���M���c�]�{���7ސ�#���m��2Z���댽H'���}��Rn��^��~N���=�S-��L��x��l��
�ɫ����Z&��d6�G���W�~hg���v��肽���e'���i������}C���ʌ������Qn�"�V�;�C��9���8��NB��T�+�k�ݳ��ۋ�f�������-�������Ǌ�����x�y/i��aY��I�LK8�Y(�i��ɔ��`
�b
�k{�S��l�+�s<�<�L���\���l�'�{�(_���<��aݑ�B��ab������'ۉ��S~��Uf���O�QY?���7���:���G�I�[�>�s��a��e���N0���ĕ�g���,�f���L���|s� d��T��wC���2�#��"=���	������`|!���0���A��0R��  �  G(��?��䓆�e���[���q|��e��Z��x6s�3�b���O���<���,��8"��\�#�� 0�]A��?T��f��\v�{���侄��ӆ�H����s��G/�������}�Ŷp���_���L���9�l�*�R"!�VW�\�%�ی2��)D�oW�W�i�<�x�F���0���������!P��mօ�%߂���{��n��\�xsI�b7�(�S? ����%9'��45��LG���Z��Jl�c�z�.j��A���/0��+���� ���o���-���y��\k��{Y�x5F��C4�/�&�N���z �")� 8�րJ���]�4�n���|���:��Z��,�����F���x����w�F�h��SV��C��1�|�$�A,�}i!��<+�@�:���M��`�؂q��~�����D��#x��$���R���!���󮀽o�u�D�e��S�%�?�/�$m#�@��n�"���-���=�\�P���c��s�T!���8����������ш���v�������)s���b�(�O�`�<�{�,�"'"�O���#���/�'�@��0T�P�f�%Pv�������Qφ�����qp���+��|��Z�}�^�p�Y�_�(�L��9�Ѕ*��!�AI��t%�<~2�D��`W���i�5�x�*���q*�����S����K���҅�܂���{��n�&�\��qI��7�J(��@ �A���<'�95�\RG�4�Z��Rl�$�z�o������!6�������'���v��v5��c�y�ymk��Y��FF�NU4�m�&���� �>1)�*8�čJ���]�� o�[�|��������A_��ʬ����������~��"�w��h��cV��!C�Ҳ1���$��>��{!��N+�J�:���M�X�`�7�q�y�~�����K���~������7���~���඀��u���e�I.S�a@��./�K�#�_�-�"���-���=�?Q�|�c�:t��  �  ;���c������F���[�������p�y]a��FQ��@�k0�� ��5�pH���	�	������#���3�gdD���T���d��Tt�Դ���爽GB��瓽�ƕ�����&��Ȅ�.br��Z��F�#G:���7�8
@��Q���g����`]��_���Pw���"��˖��Jދ�����{���k��	\���K�2;�Ұ*���f��F�
�{
����d��|�(�m-9��I��:Z�\ j�]Vy�� ��������vڔ�s���}q���V��S���@j��JS��xA��>8��n9��D�X�o�o�L���N@��
��������@��Tݏ�æ��W���s�u���f��V�Q2F��|5���%����E��
�]�� �v��5.���>�fO��_��*o��b~�D����B����������* ������.5���Sz�$Kb�ݖL�!P=��r7�s(<��J��_���w���������ӡ���������wU��'��/�p�XQa�	:Q��@��0�O� �b%��7�+�	���������#�l�3��WD�+�T���d��Kt����L䈽?���㓽�Õ�o����"��SÄ��Wr�=�Z��F�;9:���7�3�?���P���g���EV���ّ��p�����u���~ً�����l{���k�n\���K�8
;��*��������
�w}
�����(�49���I��CZ�L
j�bay��&��%���
��┽m����y���_��4���Rj��\S���A��O8�S9���D��*X���o�6����E��Շ��3ƕ�(E��}ᏽ��������v��f�ĶV�=@F���5��%����+W�c
�ļ�	���UE.�{�>�HtO���_��7o��o~�Б��zI��ޝ��_���x�������>���gz�e`b�¬L�Uf=�
�7�0><��J��_�H�w�����ʏ��  �  P��m�������ᙽ����j���e�o�N��:�/�'��$���
��� ������[�=�����l��4r���+�l>���S�pdk�B�������w���ی���]��c���z⦽����#�����}�͡d���T��Q��B\�ѻq�C���畽Ȕ���ɪ�n6�������`��н������?�v�:�]��{G��3�3]"�e��.��������6�h���!���� ���1�"E��1[���s�����L���/�������NR��b����n��̰��ݑt� ^��kR���S��Ib��z�~���z��L⥽6A��$���:l���ĝ��p�����3&n�EV��@�7�-������������ e������ ��	�{��%���7�%4L��#c�r|�
����P���	���=-��li��,����䵃�ul���X��iQ�/^W�9~i����w������n���������蚤�(ܙ� ���_�K�e���N�Z:���'�`��
�� ����6<�������1��e��+��a>���S�~\k�ͣ�����������Z��ؙ��cަ�/񛽺���_�}�t�d���T���Q�3\��q�t���ߕ�o����ª��/������?[��ḕ�b�����v���]��vG��3�(Z"�c�.� ���7���
o�������g� ���1� +E��;[��s���pS���6���������Z��B����w�����X�t�;(^�F}R���S��Yb���z�!��π���祽�E��h���:p��sȝ�	u��#���/n��!V��@�R�-��$������������3���� ���	�m���&��7��AL��0c�3|�����������5���r��3������ ���Y5l�*�X�ӀQ��tW��i���,���Þ������  �  ?(ƽX�½ya��iѨ�����Ã�o|d���E��r,�����������m�{�ܼ^�ټ�޼��鼧W��z0�m&���1�(AL�5�k�)���G�������7��.2Ľ��Ž�����ಽ-ա��鏽������n���j�Nw�Z���������x����ĽW�Ž������`䢽n6��l{�=�Y���<�k%�+��t����#?���ڼ�]ڼ���
��Q�K�"�b�9�e5V�ow�����נ��뱽�羽�Ž��ĽK��Mz��ٽ���V��.�y�:sk�hBm�\�~� ���˟����f���.�Ž��Ľ񄼽oj��.Ü��q�o�
O�Q4�B��������A8��޼'�ټq�ۼ��伳+��o_����)�0�B���`������f���٦�#ֶ�����#ƽ��½Ǽ���§�����;��-s�y<j�=jq���������p˥�c+������� ƽu�½/[���˨�|���l���Aqd�
�E��f,����)���o���O�Inܼ'�ټ�޼ ���<��$�M��1��8L���k�݇�w���ޕ��c4��2/Ľ��Ž�����۲��ϡ��㏽����>vn�N�j�>w�@���ﺙ����謺��Ľ��Ž����睳�Sߢ��1��Xd{���Y���<�/%�d(��r����?�h�ڼdbڼ�%��n��X�3�"�k�9��?V�]zw�����ޠ�󱽡ﾽa�Žc�Ľ[������KǛ�`��֗y�V�k��Sm���~�u��Sҟ��#������чŽ��Ľǈ��(n���Ɯ���l�o��O�C\4�lN�f�������V뼼߼W�ټ��ۼ{�伳J��kn�v���)���B���`�/���~m���ঽ�ݶ�=���,ƽ��½1Ƿ��ͧ��ŕ�hG��Es�xTj�q�װ���˓�xե��4������  �  �ܽ�׽ȃʽGA��⭠�6���=nh��C���%��K[���y�%�ԼR̼*�ɼWeͼ"�׼p	�3w�ю���+��:K�\|q�Ʀ��:ԥ��컽�	ν�Tٽ��۽�սtƽ�ٲ�j8������2遽A�����ԕ������#���iϽ��ٽ.�۽�
Խ��Ľ_�D蘽a1���d[�D�8����K���S�fN޼B Ѽyʼ�!ʼ'�ϼrܼM�������z5� /W�ׄ�uM��yj����½��ҽ�)۽{�ڽJ�н�A���׫�З�8��Y(��{1��z ��������foĽ��ӽҁ۽�ڽ)�Ͻ|-��J`��#0��ev�)O���.�'��W'�Q]��
ټ�μJ�ɼ�W˼,OӼ�;⼂$��!����"���?���c�(�����QԴ�ÚȽ8sֽ�ܽTHؽ�̽�����ꤽ�����
�~�⒃�Z��餢��j��8;ʽP׽5ܽ�׽j}ʽa;��G�������-ch���C���%�m���@��^�t�Լ,�˼�ɼ�Hͼ�{׼���nk�F��u�+��2K��uq�ݣ���ѥ�껽ν�Qٽ��۽�սRoƽQԲ�!2�������ၽb���醽}̕�q������#bϽ?�ٽT�۽mԽĝĽ:믽�㘽s-��H^[���8�d}�$���O�L޼� Ѽ�{ʼ�&ʼ(�ϼ8{ܼ���l����܃5�@9W�A���S��Uq���½�ҽ�1۽W�ڽ�нK��"᫽�ٗ��A���1��C:���(��c��߈��euĽ��ӽf�۽�ڽޭϽ1���c��4���v��'O��/���Z4�Ly�S(ټx3μ��ɼ9w˼/nӼ�Y��A��]���#��?��d�������۴���Ƚ�{ֽ�ܽQRؽf̽����m������������������*��揤�t���Dʽ�X׽�  �  �$�彌;׽�����V���{���m�4D��r#���
�Y/�G2ڼa	˼��¼>���"/ļ��ͼ&�޼�������j*�ӜL��;w�G"�����O�ƽv/۽h����꽏��:�ӽ�K���ʧ���l��������u��*����'��E�ʽ�uݽ�轴}�b���н�q��֠��N/��J�^�_T8�$R�����S/Լ��Ǽ:{��+����ƼscҼO.����u���4�9�Y��v��"�������UEν^�z��4��X߽��̽x���UР��؏�����7����Hf��۽���}ѽ58�k��5��wݽ\gɽ����`���tb|���P��h-�D�=x��m�!ϼC�ļ����EH¼%�ɼ! ؼ���7h��C �Q@�&h����1j��x��ս;�佫 �罔�ٽ[�ŽN���l���勽W��F͊�.q��
���JHý��׽�
�C���!5׽����Q��v���m��(D��f#���
�/� ڼI�ʼD�¼գ��Zļ�ͼ:�޼����W����)�:�L�E5w��������ƽ -۽��罂�꽓��x�ӽfF��}ħ�ջ������ȸ���m������I���ʽ nݽ����v����M�н�l��@���V+����^��N8��M������}-Լa�Ǽ�}���/����Ƽ�lҼ�9漼��}�ė4���Y��|��v��������Lνf���&�齥&߽#�̽0���ڠ��⏽>!��z@��i
���m���Ļ��ѽq=����4��ݽ�jɽ{�������j|���P�Xs-��#��������=ϼA�ļG���g¼��ɼؼ��Vv��Q ��'@�w3h�ӱ��8q�������ս��
�G!�z�ٽ��Žc$��y��K򋽢c���ي�}��?����RýI�׽���  �  �fG�4�B��6��-#�S6������Ľ�+��셆�OWc��rE��(1�fS$�T�ei�nn���&���4�*/K��k���I���ͽٌ���6���'��v9���D��0G���@���2��= �Q��k����X�=|�g������o���*��r;��oE���F�O]?�DB0�x����y�߽���&����}��"X��=��,�d[!�2������ ��*��R;��T���x�H������U�ڽ~-�f��h2.��>��pF�]F���<�-����]���.�<ὸ�'���j�
���n�0�ʟ?�D�F��PE�;���)���Lu���ѽ�������o��0N�*�6�
�'���q�����8#�X/�h�B�l_��ۃ����������,�
�� ��%4�3�A��QG�>�C�:8�V�&�C��4��_���߽/|�~���2����$���6��B��bG���B���5��*#��3�q���Ľ&�� ����Jc�meE�1�.E$��E��Z�S`�3�&��4��#K�{k��
���E��R�ͽ�����5�ٻ'��u9���D�/G��@���2��: ��������P但s�^��@��2k���*�Jn;��kE���F��Y?�!?0��
����:�߽釸�#��
�}�9X���=��,��[!�����+� �՝*��X;�.�T��x��������e�ڽ�0���c6.�>�NuF�)
F���<�6-�3������8�6"�+����^�
�
�l�0�N�?�\�F��RE��;�g�)�����x����ѽ!������o��=N���6���'�P�1��O��yH#�<g/��B�?z_�y⃽H��������
齲�
��� �*4���A��VG���C��?8���&����;�*m�e�߽t��8��1��K�$���6���B��  �  ��B�!v>�r2������
�@��T7ý춡������Pe���G�T�3���&����:��H� ��@)�ɖ7���M��Mm��S��ؕ����˽������\$��s5��,@�]�B�<�+�.�"����	����$Uཙ�ܽ�y齚H��R�F'�{A7��@�-\B�0$;�̓,�������ܽoN��x����~�;WZ��E@�%�.�"�#�����Y�r#�_<-�M�=���V��Mz�;����z���xؽ#����̖*� �9���A�]�A�o�8�u>)��n���n���,ݽ�߽�������b-�O;��cB���@�X�6��}&�8�����Z�Ͻ�!��[��+xq���P��9��w*�f�!����KZ�h�%���1�|<E��za�_���a��-&����!`�*���S0��o=���B��t?�}!4��*#�_�e����5��۽�`�1������!�x2��>���B��r>�K2����
���2ýj����GDe���G��3�|�&�^�����	� �3)�"�7���M��Cm�uO��T���Ƀ˽������[$��r5��+@��B�.}<���.�L����	����L��ܽ�p�D��M��A'�==7��@�oXB�� ;���,�*����w�ܽ�J�������~��SZ�_C@�$�.�L�#�K��\�#�*A-�E�=��V�&Vz����f����~ؽt&�=��Ě*�D�9��A�%�A�k�8��C)�*t�������6ݽ4߽�"���;��`-��Q;��eB���@�� 7�&���G����Ͻ�%��e"����q�q�P�ܟ9�K�*���!�A�j���%�2�4KE��a��e��sh���,��K
潤c����W0�ft=���B��y?�I'4��0#���Ə��NC彊�۽�m㽻=����/!�
}2���>��  �  �(6��O2�dV'��,��V�&t�5L��mC��s���.Ul�kHP��U<��$/�!�'���%���(�6�1��$@��U���s��㍽Kr����ƽ���
��V��M*�y�3���5��=0���#�#Q�v�~��=�Խ�vѽ5Aݽ���V�����lq+��W4�(�5�Q]/��f"�������T?ֽ����S������J�a�l�H��47�i,��j&�S&� +���5��rF�t�^�	��Ż���7���Aҽ�x��\��P� ��2.��b5�	�4�6�,����p��[���d߽4 ҽ3�ӽ�9佲0 ��Z��("�-'/��5�!q4�֭+�F����
���R�ʽ���+m��d�w��X�XB���2���)��%�0/'���-��:��M���h�F����A��>���R޽M-�z'���%��f1�U6���2�h�(�������｡Yٽ��н��׽6������+�V'�`#2�%6�'L2�ES'��)��S��n��F���=�������Hl��:P�qG<�/�(�'���%���(�.1��@� �U�U�s�ߍ��n��~�ƽ$����b��L*�I�3�P�5�<0�m�#�RN�0�!��4�Խ nѽ_8ݽ����}����>m+��S4�x�5��Y/��c"������&;ֽ���m��������a�D�H��37��,�Ol&��!&��#+�Ŭ5��xF���^�Z������`=���Gҽu�����?� �37.�pg5���4�#�,����*u�f��#o߽
ҽ�ӽ�B佚4 �2^��+"��)/�+�5��r4�r�+����,�
�u�@�ʽ����er��9�w�5�X��-B���2�7�)��%�>?'�{.��:�˱M���h�(���EH��ٯ���X޽�0�++���%�Bk1�%6���2��(���W�����fٽ�нv�׽���ҿ��0�D'��'2��  �  i�#�>� ���M�+���.�ؽ�	���%���g��k%{�$�`��FL�L>�Ԣ5��C3���6���@��@P� �e����������R��q½xu߽����0�n���!�c#��A�i|��,�>n콜<ӽ0�ý�����ʽiRཎ���Sg�1�*�!��j#��x����p6�x�νeE��1Û��\���}q�EY���F��:��4���3��9��)E�k�V��nn�uo���d��Lo��݆˽��齟f����R��)#�#^"�z1�R��� ��1��̽N0��+�½��н|D��y�G�M�� #�Ut"�������� ����5ŽJ����ٔ�����)�h�KR��B�۵7��P3�h5�M�<�4WJ�8�]���w��R��F������Wս�%��\f	����U �У#�צ �Ŕ��'
��!��M�ڽ��ǽJ1��	ƽ�ؽQ��K��1C������#��� ��	�y�Ο���ؽ-��$ ���a��p{�Iw`�-8L��=�?�5�L43�;�6�۟@��2P���e����������N��½�r߽=����.��l�>�!��a#��?�z��)��g�h5ӽX�ý9���f�ʽ�I�����c��O�!�2g#�@u���^��1�]�ν�A��W����Z���zq�'Y���F�P�:�C!4���3���9��.E�U�V��un��s��@i���t��Ќ˽&��4j����{��~-#��b"�P6�J��� ��;�	�̽�9��I�½h�н.L�X}�?��O��"#�5v"�V��F��z����89Ž ���ߔ�!ǂ��h�\ZR��B�)�7�Wa3��5���<�gJ�e�]��w��Y������y���]սS,���i	����� �y�#�� �E��^-
��-���ڽu�ǽ>���"ƽ�(ؽ��򽎆��G�����  �  ̛��D�b{����_����ѽ,���I��G|������&{��he���T�y�J�!�G�XLL��X�*�i��K�������KK�����l�ֽ��2� ��	�����9��|	��f �)齵|н3Ȼ��������(�߇ƽ�ݽ�������������%��l%���h�=�ʽ\���Bt��DK�����.[s�8_��P���H�UH�siO�gK]�3�p�Ň��0���s����t��edȽ��ݽ���J��t)�x���+�
���G��Ļ���Ƚ�t�������1��+⹽��ͽaQ潋Y���������>�J�	������ٽ��ý�P��!ڞ�
R�������l���Y��3M�m�G�f�I��QS�;c��sx����絗�>L���㺽1sϽ�J彊���4�����S��	������U��vؽi���-���)��\����ǿ���ս�����K�
���-A�]x�������|�ѽ����C��
v��ō��P{��Ye���T��J���G�<L�"�W�o�i�E���������F��/���N�ֽa���� �z	�R��38��z	�ld ���kvн0���K ��v����괽pƽ��ݽ��������������8��. ��-d�;�ʽ����xq��I����Ys��7_��P�Q�H�~WH�mO�#P]��p�H���G��� ���3z��CjȽ��ݽ������-�˜��0����`Q����ཫ�Ƚ�~������:��r깽-�ͽ X�u_��H�����|@��	����n	��ٽ3�ýV������X��ʱ��T$l���Y��DM���G���I��bS�hKc��x�
��缗��R��G꺽�yϽxQ彂�������˴������ a񽓂ؽ����f9��6��g	��uӿ���ս����w�
��  �  ������T��S�[޽,:ҽ��Ž�k���L��f���������/t��\g�p�c���i��x�m(�� ������ E��sB�� �Ƚ�Խ����6뽣��L���j�5��kڽ�Jǽj���ad���\���u������ݫ�io��^3ҽ������3���H*���"�ʑ�V4ڽa*ν����4��ɧ����\������&#o���d�,dd���m�x��G��g���FC�����nn���̽&�ؽ�W��.�Ȳ���	�����>�'FԽk���1���w1����������;䡽Ū���Žegؽ�a�ߪ�J��Ѩ�=�.���:ֽʽ����6���Q<��ጕ��|��.�z���j���c�bf�C�r��1������"��dǪ�x���M�Ľ��н��ܽE��U������"������/�ͽ�
��a<���ӛ����-嚽����e巽��˽�<޽B��h������o����޽�4ҽ9�Ž�e��AF��d�������y��Pnt�'Kg��rc��ui�rx�� ��������Y?��|=��˸Ƚ��Խ{��4��	��I��Vg�<��[fڽ.EǽH����]��sU���m�������ի�Zg��}+ҽ�㽩��w���$���ｶ���/ڽ{&ν����{���Ƨ�-��[�������c#o�=�d��fd�K�m�-��J��╘�RG�������s����̽�ؽ�^�[6���c������G当OԽ���������:���Ǘ�����L졽)����ŽHmؽg�m��N�����RA�0��_?ֽ�ʽa�������pC������L�����z���j��c�tf�ޠr�:�����*��yΪ�*�����Ľ��н^�ܽ��罀������!��W������ͽ����G���ߛ�d&���𚽏����﷽@�˽�E޽G���  �  үҽ�Cٽ��ܽ�c޽�Y޽Z�ܽ��ؽK8ҽ(�ǽ⍺�n�����%T�������+���"��-�R䞽����Ž�E�ʽԽ�ڽQDݽy{޽d3޽Kܽqؽ��н�Ž����p�����O����Ԅ��`��d������r��#<��3��_̽�>ս��ڽ"�ݽe�޽��ݽ��۽h׽v.Ͻ��ý#����ɥ�S���>Ԋ�������0ˉ�]6������γ�_T½_ν�[ֽ�\۽��ݽN�޽��ݽd'۽S�սsͽƒ���%��{s��XI������sQ��[��р��E���4^����ĽI�Ͻ=k׽=�۽�޽ρ޽kxݽ�ڽ��ԽC�˽2N��/W��=����J��T쇽�A�����r��♽9L���฽՚ƽ�:ѽ�^ؽ�nܽ$<޽Ro޽�ݽX�ٽ��ӽP�ɽ�񼽇������W:��浆�z��K����뎽�U����8V����Ƚ�ҽ�=ٽ(�ܽ�^޽hT޽��ܽ�ؽ*2ҽv�ǽ����������7K��c����"�����-落�۞� ���U����ʽ��ӽ(	ڽI@ݽ�w޽30޽Hܽ8ؽ�н�Ž����k������|���̈́� Y��_\������+k���4�����.X̽8սۺڽ��ݽ|�޽��ݽ"�۽1׽�+Ͻ��ý����ɥ�輖�`Ԋ�������̉��8���
��Hҳ�`X½�ν�`ֽsb۽ �ݽ�޽��ݽ*/۽�ֽ�ͽ��������N.���|��mR��`����Y���b�����Ү��d���Ľ��Ͻ�o׽X�۽�޽.�޽;}ݽx�ڽ��Խ)�˽�U���_��%����S������/K��#������꙽~T��M踽�ƽ�Aѽ�dؽ�tܽUB޽�u޽�&ݽ��ٽ�ӽ�ɽ����������LE������$��/
��v����_�������^��U�Ƚ�  �  -"��֮ƽ]�ҽ��޽-�齤� (��C^��d��#TݽG�ʽ߶�i���8���&0���_���'��p*��U�ν��[��V��׳��xr��V��,ܽ 4н��ý0E��-��Me��t䎽+����q�0f�[�c�.nk�G�{�o3��S��E���w��)\��w�ʽ��ֽ�⽋��;��D���E򽂢��e׽q�ýJ����3��,p�������ٟ���������Tս5��e�"��ev�����u��{3ؽ3̽?���n岽�~��*͗�������}���l��!d��<e���o��T���k��eښ�-����е�6�½��ν��ڽ�'�b�ｺX��n���Po�W���ѽhO��)ꪽi���N��u���� �����S_Ƚ�_۽��꽓��@��ɲ���꽗�58Խ�Ƚ����I���W򠽟K���r��fw�t�h��dc�W�g�adu�����Α��k��U�����ʨƽ��ҽX�޽��8��9"���W��t�뽁Lݽ��ʽ�ֶ�����px��6&���U�����C!����ν��/T��P�������m��R�m)ܽ�0н\�ýwA��	���`��4ߎ�X���_�q���e��c�w_k�d�{�,���K��H���q���U����ʽl�ֽD��T�콏���@��'C�y�罁d׽��ý䬰��3���p��%����۟��������VXս*�Zj�'���{��ٻ��㽛:ؽ�"̽A¿���i���֗�������}�"�l��2d�Me���o��[��Ar��<���s����յ���½��νn�ڽ�,潛�ｗ^������vｉ���$ѽ�X�����;s��Y��m���Y*��=ƴ��gȽ�g۽ʎ�I��eF��и��꽷	཭>Խ�ȽG�������B���$U���|���zw���h��yc���g�Gxu�V)��fב�t������  �  �G��k6���ӽ���"��x���w�\����
�!*��F�tԽ�Ǿ��|���B���ܲ�.ý��ٽ6��`����������*�����6��Hν�ҹ�yX���ݖ��E���2w�W?b�t�R��I���G���M���Z�Lm�{d��a&��Yȟ��Z��H�Ľ0Nڽz9�DF�/
��[�����<�������&�̽� ���ۭ�@�� J��� ʽ�$⽪���NV��c�A����
�XH�$�򽪷ܽT;ǽg��Ϛ�����ʃ���o��U\�l�N�� H�>�H�_CQ��.`���t�����"��g��b����˽��὜M��9<�4����<t��e�]����ܽmTŽ80���k���r�����$�ѽ{�� � �	�}U�
��;���& �d��qսk��"B��c ��L茽�%�D�h��"W���K��G��J�Q�U��lf��m|��T���W��TA���0��P	ӽU���������t�!��$�
�(&�>�?kԽ½���r��8��Ҳ��ý��ٽ���[�,��\����r(�6���P�EνϹ��T���ٖ��@���(w��3b��R�ۋI�'�G���M�d�Z��=m��]����������T����ĽIڽ�4�8D�<-
�;Z�����;�z�����ş̽
��cܭ�SA���K���"ʽ\'����CX��e������
�ZK���򽤾ܽ�Bǽ�n������^ˑ��Ӄ�d�o�Gg\��N�31H�
I�NRQ�i<`�Z�t��Ć�(��l�������˽B�ὮR��?�Y�;��0x�Fj��f����ܽ�^Ž�:���v��W}��ü���ѽ�� ���	��X�&��,���) ��i��wսr��MI��/(�������7�7�h�\6W���K��G��K�>�U��~f��~|�i\���^���  �  -l��0���Eaڽ�a������� !���#���ϙ�g���@��ֽRwŽ�M���\ȽM"ܽ2���]�
��=��!���#�!�������`n�}�ӽ ���tf��lU���:v���\��zI�c2<�+�4�s3��-8�d�B�AiS�&j�\������*T����ƽ���S��%w�6��"��"����
E�����罿�ϽoB½y���<�ͽp��A� �������"�#��T�����t��|�ɽG
��G:���|��u�l�.�U�VD��9���3�L4��;�9�G�29Z��s��T����q���gн������7��M#�e�!�ou�D���"����޽��ɽ���]4ĽhcԽ���] �N0�1���x#���!�����f�����~�ݽ����v����������Hqd�l*O���?��6��*3�J�5���>��-M���a��|� m���e�������[ڽZ\��}��ѧ�!�6�#�m�������7��ֽ�lŽ�B���QȽ�ܽ������
�:9��� �u�#�����l��/j򽏰ӽ@���rb��!Q��y1v�L�\�ZoI�X&<�e�4��e3��8���B��[S��j�ڥ������VN����ƽ�����&u�w���"���"����TD���������Ͻ"C½������ͽ��佪� ���������"��#���K��1��P���ɽ���BB������E�l�&�U�gD�R9���3��[4�\;��G��EZ�js�Z������B����kн���X�������
�#���!�z�:��6-����޽�ʽ���2?Ľ�mԽy���m4���T|#���!�����i�?���]�ݽ����G��핑�� ��l�d�z<O�J�?�"�6��=3�
�5���>��>M���a���|��s���  �  bȢ�!���佇i��*��(�]�2�j$6���1�mL&��:�C����0�ֽ
�н�Mڽ�/񽸜�z�TW)��Z3�&6���0���$��&���Mܽ�湽М�Yz���g�jlL��9�:�-�'���%�]�)�%�3�V5C��"Z��y�n����B��\n̽q�G����?W,���4�r�5���.��L!�b�,������(=ӽ!aҽ_��6���l����`-�Q5�S05�f�-�Q�����V���Jн;����^��<�}�� ]�&OE�M�4�E�*���%���&��w,���7�|�I�(�c��5���뙽_��x>ؽ����I�A#�t�/�$�5��4���*������
��Y���0ܽ6ѽu~ս�:����_F��$���0�s6��x3�7�)�J���*�轇�Ľ�٥�����#�q��LT��?�\�0���(��%���'�?�/�F1=�ƎQ��n��(��]¢��������f�(�(�[�2�!6���1�8H&��5�;�����ֽ��н:Bڽj$�Y��o��R)��V3�u6���0���$�U$����Iܽ~⹽�˜� v����f�9bL�ޤ9�gw-���&���%��)��z3��'C��Z�S�y�a���=��i̽�������U,�/�4�;�5���.�L!��a�ӛ�����=ӽ[bҽ!�����m�ʊ�zb-��5��25��-�?��9��]���QнĐ���f��k�}�;1]��_E���4���*��	&�П&�f�,�=	8�
�I�ǣc�;����d��kCؽ����*D#���/�	�5�K
4�e�*�����
�$e��1<ܽ}Aѽ��սfE�����J��$�B�0��6��{3��)� �ǎ�ӱ轒�Ľ�ॽƣ����q�s]T�*?�c�0��(�T�%�(���/��A=�Z�Q�<)n�/���  �  �f��>DŽ��콧�!��2���>���B�r>�f�1�� �|��~�����7ܽ�?潵D��C'�g9$�"�4�^�?��B���<�m/�}���-���h-���ǜ�!$���_���C�01�_^%��0����!��++���:��%R���s���������ѽU��m4���'���7�*0A�`7B��:��),�����������޽j�ݽf�����;*��^9�4�A�J�A�0(9���)�������\Dֽ�����t��ex��FU�&�<��},��"��5�D��Y^$�?�/��uA��\�ͭ��픙��;���0߽���"B�҈-���;���B��@�E~6��?&�d>��]�|P��Oܽj��hz��b�
�����/�Q
=���B�`�?�V�4�hE#�5i�X���fɽ�Ц�BV3k��L��6�ޔ(�
� �_��n �l'�M�4�9CI��4g�?���`���>Ž[��  �z!�A�2���>�"�B��>� �1�� �[��������⽎�۽�3�?9���!�;4$�`�4��?�D�B�1�<�'j/����+�ֺ�L)���Ü������_�o�C�+%1��R%��$�	���!�>+�W�:��R�A�s��������ѽ���B2���'��7��.A�-6B�)�:�),���q��ڼ｡�޽��ݽ'�B�w��X=*��`9�a�A���A��*9���)�>��C���xKֽ����z|��gx��VU���<��,�B�"��E�U���l$���/��A�/\�:�������@���5߽,���D���-�K�;���B�]�@�&�6��D&��C��c�3\�t[ܽ�	�A���v�
�f��T�/�=���B�k�?�%�4�H#��k�ߩ�lɽ�֦�4���]Bk��'L�ܜ6�y�(��� �[��#" �&}'���4�|RI��Bg��E���  �  �ꣽiǽ�>�w�uU$�y�6�+KC�.dG��~B�'�5�_�#����jb��)�潩�߽q���x+�-�'�9�5VD�CG��3A��63�x��&s	���'���$��-����]��rA�L�.���"�̦�����h��(��	8�]�O�~r��l���׮��+Խ��������+���;�L�E� �F���>�I0����ƭ	�=8���|���b�1�����.�j�=��IF�4F��N=��'-��b����Y�ؽ����k��w�v��R��*:��)�. �I��;���!���,���>���Y�������*���?��3���@�x@1���?��G�EE�p�:�}�)�3S����Q�콎4�i��"������R!���3��hA�FG�m,D���8��&���F��Q˽�s��~����]i���I��3���%���R�����$�H2�|�F��Fe��ه��䣽� ǽ�9�t��R$���6�!HC��`G��zB�ۡ5���#����kW�������߽Re� ��%���'�N9��QD�1?G�<0A��33����p	�ɤ�������ɒ����]��hA�d�.�.�"����܁��[��|(���7���O��q�g��$Ү�Z&Խ������+���;�ڢE�κF��>��0�w����	�l8��X}���#��U�����.�U�=�'LF�y6F�4Q=��*-��e�J��o�ؽ~����s��i�v�V
S�N;:�Z�)�B' ��� J���!�$�,�!�>�Y�Y���Gƙ�1���R������C��C1�F@��G��E�[�:���)��X������H@����-�����xW!�(�3�LlA��IG�w/D�x�8���&��������V˽z��`����li���I���3�H&��"��d������$�u2���F��Te�<����  �  �f��>DŽ��콧�!��2���>���B�r>�f�1�� �|��~�����7ܽ�?潵D��C'�g9$�"�4�^�?��B���<�m/�}���-���h-���ǜ�!$���_���C�01�_^%��0����!��++���:��%R���s���������ѽU��m4���'���7�*0A�`7B��:��),�����������޽j�ݽf�����;*��^9�4�A�J�A�0(9���)�������\Dֽ�����t��ex��FU�&�<��},��"��5�D��Y^$�?�/��uA��\�ͭ��픙��;���0߽���"B�҈-���;���B��@�E~6��?&�d>��]�|P��Oܽj��hz��b�
�����/�Q
=���B�`�?�V�4�hE#�5i�X���fɽ�Ц�BV3k��L��6�ޔ(�
� �_��n �l'�M�4�9CI��4g�?���`���>Ž[��  �z!�A�2���>�"�B��>� �1�� �[��������⽎�۽�3�?9���!�;4$�`�4��?�D�B�1�<�'j/����+�ֺ�L)���Ü������_�o�C�+%1��R%��$�	���!�>+�W�:��R�A�s��������ѽ���B2���'��7��.A�-6B�)�:�),���q��ڼ｡�޽��ݽ'�B�w��X=*��`9�a�A���A��*9���)�>��C���xKֽ����z|��gx��VU���<��,�B�"��E�U���l$���/��A�/\�:�������@���5߽,���D���-�K�;���B�]�@�&�6��D&��C��c�3\�t[ܽ�	�A���v�
�f��T�/�=���B�k�?�%�4�H#��k�ߩ�lɽ�֦�4���]Bk��'L�ܜ6�y�(��� �[��#" �&}'���4�|RI��Bg��E���  �  bȢ�!���佇i��*��(�]�2�j$6���1�mL&��:�C����0�ֽ
�н�Mڽ�/񽸜�z�TW)��Z3�&6���0���$��&���Mܽ�湽М�Yz���g�jlL��9�:�-�'���%�]�)�%�3�V5C��"Z��y�n����B��\n̽q�G����?W,���4�r�5���.��L!�b�,������(=ӽ!aҽ_��6���l����`-�Q5�S05�f�-�Q�����V���Jн;����^��<�}�� ]�&OE�M�4�E�*���%���&��w,���7�|�I�(�c��5���뙽_��x>ؽ����I�A#�t�/�$�5��4���*������
��Y���0ܽ6ѽu~ս�:����_F��$���0�s6��x3�7�)�J���*�轇�Ľ�٥�����#�q��LT��?�\�0���(��%���'�?�/�F1=�ƎQ��n��(��]¢��������f�(�(�[�2�!6���1�8H&��5�;�����ֽ��н:Bڽj$�Y��o��R)��V3�u6���0���$�U$����Iܽ~⹽�˜� v����f�9bL�ޤ9�gw-���&���%��)��z3��'C��Z�S�y�a���=��i̽�������U,�/�4�;�5���.�L!��a�ӛ�����=ӽ[bҽ!�����m�ʊ�zb-��5��25��-�?��9��]���QнĐ���f��k�}�;1]��_E���4���*��	&�П&�f�,�=	8�
�I�ǣc�;����d��kCؽ����*D#���/�	�5�K
4�e�*�����
�$e��1<ܽ}Aѽ��սfE�����J��$�B�0��6��{3��)� �ǎ�ӱ轒�Ľ�ॽƣ����q�s]T�*?�c�0��(�T�%�(���/��A=�Z�Q�<)n�/���  �  -l��0���Eaڽ�a������� !���#���ϙ�g���@��ֽRwŽ�M���\ȽM"ܽ2���]�
��=��!���#�!�������`n�}�ӽ ���tf��lU���:v���\��zI�c2<�+�4�s3��-8�d�B�AiS�&j�\������*T����ƽ���S��%w�6��"��"����
E�����罿�ϽoB½y���<�ͽp��A� �������"�#��T�����t��|�ɽG
��G:���|��u�l�.�U�VD��9���3�L4��;�9�G�29Z��s��T����q���gн������7��M#�e�!�ou�D���"����޽��ɽ���]4ĽhcԽ���] �N0�1���x#���!�����f�����~�ݽ����v����������Hqd�l*O���?��6��*3�J�5���>��-M���a��|� m���e�������[ڽZ\��}��ѧ�!�6�#�m�������7��ֽ�lŽ�B���QȽ�ܽ������
�:9��� �u�#�����l��/j򽏰ӽ@���rb��!Q��y1v�L�\�ZoI�X&<�e�4��e3��8���B��[S��j�ڥ������VN����ƽ�����&u�w���"���"����TD���������Ͻ"C½������ͽ��佪� ���������"��#���K��1��P���ɽ���BB������E�l�&�U�gD�R9���3��[4�\;��G��EZ�js�Z������B����kн���X�������
�#���!�z�:��6-����޽�ʽ���2?Ľ�mԽy���m4���T|#���!�����i�?���]�ݽ����G��핑�� ��l�d�z<O�J�?�"�6��=3�
�5���>��>M���a���|��s���  �  �G��k6���ӽ���"��x���w�\����
�!*��F�tԽ�Ǿ��|���B���ܲ�.ý��ٽ6��`����������*�����6��Hν�ҹ�yX���ݖ��E���2w�W?b�t�R��I���G���M���Z�Lm�{d��a&��Yȟ��Z��H�Ľ0Nڽz9�DF�/
��[�����<�������&�̽� ���ۭ�@�� J��� ʽ�$⽪���NV��c�A����
�XH�$�򽪷ܽT;ǽg��Ϛ�����ʃ���o��U\�l�N�� H�>�H�_CQ��.`���t�����"��g��b����˽��὜M��9<�4����<t��e�]����ܽmTŽ80���k���r�����$�ѽ{�� � �	�}U�
��;���& �d��qսk��"B��c ��L茽�%�D�h��"W���K��G��J�Q�U��lf��m|��T���W��TA���0��P	ӽU���������t�!��$�
�(&�>�?kԽ½���r��8��Ҳ��ý��ٽ���[�,��\����r(�6���P�EνϹ��T���ٖ��@���(w��3b��R�ۋI�'�G���M�d�Z��=m��]����������T����ĽIڽ�4�8D�<-
�;Z�����;�z�����ş̽
��cܭ�SA���K���"ʽ\'����CX��e������
�ZK���򽤾ܽ�Bǽ�n������^ˑ��Ӄ�d�o�Gg\��N�31H�
I�NRQ�i<`�Z�t��Ć�(��l�������˽B�ὮR��?�Y�;��0x�Fj��f����ܽ�^Ž�:���v��W}��ü���ѽ�� ���	��X�&��,���) ��i��wսr��MI��/(�������7�7�h�\6W���K��G��K�>�U��~f��~|�i\���^���  �  -"��֮ƽ]�ҽ��޽-�齤� (��C^��d��#TݽG�ʽ߶�i���8���&0���_���'��p*��U�ν��[��V��׳��xr��V��,ܽ 4н��ý0E��-��Me��t䎽+����q�0f�[�c�.nk�G�{�o3��S��E���w��)\��w�ʽ��ֽ�⽋��;��D���E򽂢��e׽q�ýJ����3��,p�������ٟ���������Tս5��e�"��ev�����u��{3ؽ3̽?���n岽�~��*͗�������}���l��!d��<e���o��T���k��eښ�-����е�6�½��ν��ڽ�'�b�ｺX��n���Po�W���ѽhO��)ꪽi���N��u���� �����S_Ƚ�_۽��꽓��@��ɲ���꽗�58Խ�Ƚ����I���W򠽟K���r��fw�t�h��dc�W�g�adu�����Α��k��U�����ʨƽ��ҽX�޽��8��9"���W��t�뽁Lݽ��ʽ�ֶ�����px��6&���U�����C!����ν��/T��P�������m��R�m)ܽ�0н\�ýwA��	���`��4ߎ�X���_�q���e��c�w_k�d�{�,���K��H���q���U����ʽl�ֽD��T�콏���@��'C�y�罁d׽��ý䬰��3���p��%����۟��������VXս*�Zj�'���{��ٻ��㽛:ؽ�"̽A¿���i���֗�������}�"�l��2d�Me���o��[��Ar��<���s����յ���½��νn�ڽ�,潛�ｗ^������vｉ���$ѽ�X�����;s��Y��m���Y*��=ƴ��gȽ�g۽ʎ�I��eF��и��꽷	཭>Խ�ȽG�������B���$U���|���zw���h��yc���g�Gxu�V)��fב�t������  �  үҽ�Cٽ��ܽ�c޽�Y޽Z�ܽ��ؽK8ҽ(�ǽ⍺�n�����%T�������+���"��-�R䞽����Ž�E�ʽԽ�ڽQDݽy{޽d3޽Kܽqؽ��н�Ž����p�����O����Ԅ��`��d������r��#<��3��_̽�>ս��ڽ"�ݽe�޽��ݽ��۽h׽v.Ͻ��ý#����ɥ�S���>Ԋ�������0ˉ�]6������γ�_T½_ν�[ֽ�\۽��ݽN�޽��ݽd'۽S�սsͽƒ���%��{s��XI������sQ��[��р��E���4^����ĽI�Ͻ=k׽=�۽�޽ρ޽kxݽ�ڽ��ԽC�˽2N��/W��=����J��T쇽�A�����r��♽9L���฽՚ƽ�:ѽ�^ؽ�nܽ$<޽Ro޽�ݽX�ٽ��ӽP�ɽ�񼽇������W:��浆�z��K����뎽�U����8V����Ƚ�ҽ�=ٽ(�ܽ�^޽hT޽��ܽ�ؽ*2ҽv�ǽ����������7K��c����"�����-落�۞� ���U����ʽ��ӽ(	ڽI@ݽ�w޽30޽Hܽ8ؽ�н�Ž����k������|���̈́� Y��_\������+k���4�����.X̽8սۺڽ��ݽ|�޽��ݽ"�۽1׽�+Ͻ��ý����ɥ�輖�`Ԋ�������̉��8���
��Hҳ�`X½�ν�`ֽsb۽ �ݽ�޽��ݽ*/۽�ֽ�ͽ��������N.���|��mR��`����Y���b�����Ү��d���Ľ��Ͻ�o׽X�۽�޽.�޽;}ݽx�ڽ��Խ)�˽�U���_��%����S������/K��#������꙽~T��M踽�ƽ�Aѽ�dؽ�tܽUB޽�u޽�&ݽ��ٽ�ӽ�ɽ����������LE������$��/
��v����_�������^��U�Ƚ�  �  ������T��S�[޽,:ҽ��Ž�k���L��f���������/t��\g�p�c���i��x�m(�� ������ E��sB�� �Ƚ�Խ����6뽣��L���j�5��kڽ�Jǽj���ad���\���u������ݫ�io��^3ҽ������3���H*���"�ʑ�V4ڽa*ν����4��ɧ����\������&#o���d�,dd���m�x��G��g���FC�����nn���̽&�ؽ�W��.�Ȳ���	�����>�'FԽk���1���w1����������;䡽Ū���Žegؽ�a�ߪ�J��Ѩ�=�.���:ֽʽ����6���Q<��ጕ��|��.�z���j���c�bf�C�r��1������"��dǪ�x���M�Ľ��н��ܽE��U������"������/�ͽ�
��a<���ӛ����-嚽����e巽��˽�<޽B��h������o����޽�4ҽ9�Ž�e��AF��d�������y��Pnt�'Kg��rc��ui�rx�� ��������Y?��|=��˸Ƚ��Խ{��4��	��I��Vg�<��[fڽ.EǽH����]��sU���m�������ի�Zg��}+ҽ�㽩��w���$���ｶ���/ڽ{&ν����{���Ƨ�-��[�������c#o�=�d��fd�K�m�-��J��╘�RG�������s����̽�ؽ�^�[6���c������G当OԽ���������:���Ǘ�����L졽)����ŽHmؽg�m��N�����RA�0��_?ֽ�ʽa�������pC������L�����z���j��c�tf�ޠr�:�����*��yΪ�*�����Ľ��н^�ܽ��罀������!��W������ͽ����G���ߛ�d&���𚽏����﷽@�˽�E޽G���  �  ̛��D�b{����_����ѽ,���I��G|������&{��he���T�y�J�!�G�XLL��X�*�i��K�������KK�����l�ֽ��2� ��	�����9��|	��f �)齵|н3Ȼ��������(�߇ƽ�ݽ�������������%��l%���h�=�ʽ\���Bt��DK�����.[s�8_��P���H�UH�siO�gK]�3�p�Ň��0���s����t��edȽ��ݽ���J��t)�x���+�
���G��Ļ���Ƚ�t�������1��+⹽��ͽaQ潋Y���������>�J�	������ٽ��ý�P��!ڞ�
R�������l���Y��3M�m�G�f�I��QS�;c��sx����絗�>L���㺽1sϽ�J彊���4�����S��	������U��vؽi���-���)��\����ǿ���ս�����K�
���-A�]x�������|�ѽ����C��
v��ō��P{��Ye���T��J���G�<L�"�W�o�i�E���������F��/���N�ֽa���� �z	�R��38��z	�ld ���kvн0���K ��v����괽pƽ��ݽ��������������8��. ��-d�;�ʽ����xq��I����Ys��7_��P�Q�H�~WH�mO�#P]��p�H���G��� ���3z��CjȽ��ݽ������-�˜��0����`Q����ཫ�Ƚ�~������:��r깽-�ͽ X�u_��H�����|@��	����n	��ٽ3�ýV������X��ʱ��T$l���Y��DM���G���I��bS�hKc��x�
��缗��R��G꺽�yϽxQ彂�������˴������ a񽓂ؽ����f9��6��g	��uӿ���ս����w�
��  �  i�#�>� ���M�+���.�ؽ�	���%���g��k%{�$�`��FL�L>�Ԣ5��C3���6���@��@P� �e����������R��q½xu߽����0�n���!�c#��A�i|��,�>n콜<ӽ0�ý�����ʽiRཎ���Sg�1�*�!��j#��x����p6�x�νeE��1Û��\���}q�EY���F��:��4���3��9��)E�k�V��nn�uo���d��Lo��݆˽��齟f����R��)#�#^"�z1�R��� ��1��̽N0��+�½��н|D��y�G�M�� #�Ut"�������� ����5ŽJ����ٔ�����)�h�KR��B�۵7��P3�h5�M�<�4WJ�8�]���w��R��F������Wս�%��\f	����U �У#�צ �Ŕ��'
��!��M�ڽ��ǽJ1��	ƽ�ؽQ��K��1C������#��� ��	�y�Ο���ؽ-��$ ���a��p{�Iw`�-8L��=�?�5�L43�;�6�۟@��2P���e����������N��½�r߽=����.��l�>�!��a#��?�z��)��g�h5ӽX�ý9���f�ʽ�I�����c��O�!�2g#�@u���^��1�]�ν�A��W����Z���zq�'Y���F�P�:�C!4���3���9��.E�U�V��un��s��@i���t��Ќ˽&��4j����{��~-#��b"�P6�J��� ��;�	�̽�9��I�½h�н.L�X}�?��O��"#�5v"�V��F��z����89Ž ���ߔ�!ǂ��h�\ZR��B�)�7�Wa3��5���<�gJ�e�]��w��Y������y���]սS,���i	����� �y�#�� �E��^-
��-���ڽu�ǽ>���"ƽ�(ؽ��򽎆��G�����  �  �(6��O2�dV'��,��V�&t�5L��mC��s���.Ul�kHP��U<��$/�!�'���%���(�6�1��$@��U���s��㍽Kr����ƽ���
��V��M*�y�3���5��=0���#�#Q�v�~��=�Խ�vѽ5Aݽ���V�����lq+��W4�(�5�Q]/��f"�������T?ֽ����S������J�a�l�H��47�i,��j&�S&� +���5��rF�t�^�	��Ż���7���Aҽ�x��\��P� ��2.��b5�	�4�6�,����p��[���d߽4 ҽ3�ӽ�9佲0 ��Z��("�-'/��5�!q4�֭+�F����
���R�ʽ���+m��d�w��X�XB���2���)��%�0/'���-��:��M���h�F����A��>���R޽M-�z'���%��f1�U6���2�h�(�������｡Yٽ��н��׽6������+�V'�`#2�%6�'L2�ES'��)��S��n��F���=�������Hl��:P�qG<�/�(�'���%���(�.1��@� �U�U�s�ߍ��n��~�ƽ$����b��L*�I�3�P�5�<0�m�#�RN�0�!��4�Խ nѽ_8ݽ����}����>m+��S4�x�5��Y/��c"������&;ֽ���m��������a�D�H��37��,�Ol&��!&��#+�Ŭ5��xF���^�Z������`=���Gҽu�����?� �37.�pg5���4�#�,����*u�f��#o߽
ҽ�ӽ�B佚4 �2^��+"��)/�+�5��r4�r�+����,�
�u�@�ʽ����er��9�w�5�X��-B���2�7�)��%�>?'�{.��:�˱M���h�(���EH��ٯ���X޽�0�++���%�Bk1�%6���2��(���W�����fٽ�нv�׽���ҿ��0�D'��'2��  �  ��B�!v>�r2������
�@��T7ý춡������Pe���G�T�3���&����:��H� ��@)�ɖ7���M��Mm��S��ؕ����˽������\$��s5��,@�]�B�<�+�.�"����	����$Uཙ�ܽ�y齚H��R�F'�{A7��@�-\B�0$;�̓,�������ܽoN��x����~�;WZ��E@�%�.�"�#�����Y�r#�_<-�M�=���V��Mz�;����z���xؽ#����̖*� �9���A�]�A�o�8�u>)��n���n���,ݽ�߽�������b-�O;��cB���@�X�6��}&�8�����Z�Ͻ�!��[��+xq���P��9��w*�f�!����KZ�h�%���1�|<E��za�_���a��-&����!`�*���S0��o=���B��t?�}!4��*#�_�e����5��۽�`�1������!�x2��>���B��r>�K2����
���2ýj����GDe���G��3�|�&�^�����	� �3)�"�7���M��Cm�uO��T���Ƀ˽������[$��r5��+@��B�.}<���.�L����	����L��ܽ�p�D��M��A'�==7��@�oXB�� ;���,�*����w�ܽ�J�������~��SZ�_C@�$�.�L�#�K��\�#�*A-�E�=��V�&Vz����f����~ؽt&�=��Ě*�D�9��A�%�A�k�8��C)�*t�������6ݽ4߽�"���;��`-��Q;��eB���@�� 7�&���G����Ͻ�%��e"����q�q�P�ܟ9�K�*���!�A�j���%�2�4KE��a��e��sh���,��K
潤c����W0�ft=���B��y?�I'4��0#���Ə��NC彊�۽�m㽻=����/!�
}2���>��  �  Up��)���鳑�{ၾK6_�!�:��8����}uν�w���Ε�>���8�v��nk�D]h�63m�/]z�˪���[����
?׽���V5 ��|B��g��������f���@��EϚ��쎾�U~�;�]��)B�M41���-��9�'lP���o��6��N2����������N���܌�t�w� �R���.�4?���
K½!���h���ח��N�q��{i�Gi�J�p�)b���č��⡽W~��%t���#+�w�N�|�s�*!��z�������@��.s����5s���S��;�f~.�0�R�?�0Z���z��M��8ę����9�������������k��F���#����l�۽rQ��e����E��|V|�c-n�@sh���j���t�B1��邏�c���?ʽ���W��f�6��[�����#������Y`���l��u������9h��ZJ��k5��g-�k�3�+G�J�d��Ԃ��������Kn��c���[�������3_���:�L6�����oν�q��	ȕ�G�����v��_k�rNh��$m�mOz�r���?V��鳽;׽R��.4 �|B��~g�˲��w������U@��jΚ�c뎾�R~�Û]��%B��/1��-��9�3gP�̆o�#4�� 0��U�������s���bڌ�x�w�a�R�U�.�M=��~꽘H½U���=���K���o�q�B}i��i��p��d���Ǎ�_桽����+y����&+� �N�]�s�F#��R|�����$C���u����k;s�R�S�B#;���.�
"0��?�/4Z� �z�O��jř��������6���J�����k�N�F���#����<�۽W���ǜ��L��`e|��<n�-�h���j�L�t��8��X���%j���Fʽk
�����Ŝ6�#[�����%�����b���o��7x��p���Ah�bJ�&s5�5o-���3���G���d��ׂ����k����  �  �����Ә��d��nV~�R-[� �7��������&ϽH���ŗ�巇���z��}o��bl�Gq�\�~������C���V��f�׽�c�f����?��%c��ׂ��4���H��/d�����5�����x�<Y��q>�h.���*���5��AL��gj��������#��"������f�r�:O��,�:�ON�AUýe[���������	
v�.�m�%m�<�t��y��eЏ���������Jk彿&�\)��AK���n�R���锾K͛��k��rߓ�6ˆ�f�m�OO���7�c+���,��<�|�U��"u�u��=��)��eᚾT���z����g�_lC��"�0=��ܽ���꟞�|W���A���Cr�yl�J�n��y��H��c���+��K˽gt��<��j4�-W�J�z��㌾����c���R���y��^����Pc��`F�2�?U*�X�0��C���_����P���!䘾����6Ҙ�Gc���S~��*[���7��������� Ͻ ��+���߰��E�z��no��Sl�a8q�oz~�2����=���Q��N�׽�a�3��ˊ?�;%c��ׂ�F4��4H���c��������۷x��Y��m>��-��*� �5��<L�cj����æ���뚾�!��J���m�r�g7O�ƴ,�-8�6K��Rý�Y��笑�2���+
v���m��m���t�S|��~ӏ�N������Np彖)��)�EK���n�l��씾�ϛ�[n��⓾�͆���m��TO��7�Vh+���,�q
<���U�&u����p���)��'⚾��������g��mC�1"�=?�g!ܽ����R����^��)I��USr��l�e�n�q y�[P��ԩ��M	��&˽{������4��0W��z��匾F�������)�����������Wc�hF�j 2�\*�i�0�֢C�L�_�����s显�  �  gő������C��N�o�TYP��
1���������Mҽ����UX���}��M����
|���x�H�}�#ㅽ腑�����Rv���ڽ e������7��jW�jv�����7ɏ�4���2ǌ�U����h�	L���3�C�$��"�2�+�zu@���[���x�s���V>��'i��J���!���`e��E��'�[����꽑rǽAZ��d���i��}y����y�yy��R.������f˩��Ľ����;	���#��9B�i�a�O�#
�����P���Ӊ���{� _�3<C�<�-���"���#�=�1��I�{�e�	耾^܋��_��wO��ꈾ?5y�m�Z�YG;�ۚ�i��a޽�����������膽��~�3�x��0{����{��C��׳��Ɏν ��j��;�-���L�]-l�H���򹑾8��Q��"�r��qU�1;���(�i�!�A'��8�$GR��ao� 	���b��hÑ��~��+B����o��VP�%1���#���HҽI����Q��pv���3�{�>�x�*�}��ۅ�7������q��[ڽFc�;����7�-jW��
v�?����ȏ�����Rƌ��S����h��L���3���$�"�p�+��p@��[���x�3���6<��-g��z�� ���]e�W�E��'�}�����(pǽ|X���b��ui���y�� �y��{y��À��0������ϩ�FĽ����>	���#�s=B�>�a�BS�a��' ��ճ���Չ�F�{��%_��AC���-�.�"�z�#�ò1��I���e��逾�݋��`��?P���ꈾ}6y���Z��H;�������|#޽ސ��i���7$����
���x�kA{����V���J��
�����ν�&�������-�"�L�1l��������v������#T����r��xU�;";���(���!��G'���8�XMR�fgo�����d���  �  �,��c�	�p��'[�B���(�í�������ڽ�2��)��� ��L͏�����0��,/��C쑽�G��{d��=�Ž�|������M.�O�G�td`�\�t�-��������c{�1ki���Q�h�8�X$�pL�!��~A�B�.��uF��K_�fet�ȹ������a�{�3j�N�R�h�9��� ��
����F;ѽ9����B��Җ�R���函�����8������i��)-���2ν�%��e��(���6��2P���g��z������ ���Iv�l�a��9I��J1����?�tx��:"�hL6���N���f�F�y�����&���v���b��J�?1�u�g���佒bȽF����韽�	��LȊ��?��V����ˎ�i�����p���5|׽}����I�+&��4?��uX���n�L~��*��e�}Ap��Y�c�@��P*�D{��l��I�,'(��3>�+W�@n�U.~��*���{��p�E%[��B�D�(�)��W�����ڽ#,��"�����vŏ�����(��9'���䑽�@��^����Ž;x�0��p���L.�h�G��c`���t��������b{��hi�)�Q��8��$�DH�����<���.��pF�G_�at���������ؐ{��/j�q�R��9��� ��
�����8ѽ|����A���і�g��x懽ʠ���:��f����l���0���6ν�*콜h��+��6��6P���g�Hz�Á� #���Nv���a�?I��O1����-D�B}�?"�bP6�	�N���f���y������&��s�v���b�X�J��1�i��
�7���hȽE���|񟽫���Њ�uH��ۥ��Ԏ�y����#������"�׽!����L�n&��7?�UyX���n�uP~�	-��wj�PGp�C�Y���@��W*�'��rs�FP��-(��9>��0W�<n��2~��  �  ;a�c�^�[U��.F���4���"��B�X��7�G�Խ�)�����,ۡ�?����`������^��uu��,xĽd�ٽ���V�������&���8�d�I���W�-`��`�o�X���I��t6�^J"�ta�G��/����A(��V-�g�A���R�0^��Wa�EU\��P�.�@���.��+���F�����ͽ@��������B��J뗽+���N���X	��W/˽@e������e�zJ��,���>���N�N[�&(a���^���T��C�u�/�m��
�wL��J����_+ ��)4��G���W��*`�v�`�fY�ؑK�k�:�*�(���'����08ܽ��ƽ6@�����l͛��t���$������U@��I��DҽCp�"��6���� �ެ2��ND��S��^��[a��W\���O��4=�M�(�j���	�š�������R�&��:�8�M��G[�B7a��^�kU�1,F�j�4�q�"�Y@�GU�b1콂�Խ�"��9��ҡ�����(X��g���V���m��6qĽ=�ٽs��*�������&���8�i�I���W�`�v�`���X�h�I��q6�G"��]�@���������#�fR-��A���R�,^� Ta��Q\�֑P�g~@�B�.��)�,�W|��b�U�ͽ( ��$��&����B���엽�������d���2˽�iὢ���xh��M�z�,�D�>���N�`R[��,a���^���T��C���/�����hQ�OO�+��D/ �c-4�n�G�1�W��,`�8�`��Y�a�K��:��(�-����	����>ܽq�ƽQH������J֛��}���-��7����H��0���KҽAw�r��i��� �#�2��QD�ʪS�^�,`a��\\���O��:=���(��p�D�	�P�����߭��&�[�:��M��K[��  �  ��?��@�Ҵ<�ru5��y,���"��E��l�W�}����߽�˽̺��g���[����������@Ͻ��㽛����u�`��m�%�q�.�tE7�g�=�<�@�h�>��7���*�G���&�7�����뽢���@����M����#�2�U<�Ҙ@��?�/�:��2�+P)�e�����
����%j�gؽ�Ž/���ƀ������R���3ýI�ս���9] ���
����q���=(��1�e�9��_?���@��<�RX3�4�%����N��,��E(�[������}	��-���(���5�U'>�3�@�Jt>��"8���/��&��}���L��M���l,��aѽ=�������w������H����Ƚ�ܽ{?�q���J�,.��!��j+�5�4�<��`@�@��6:��%/��U ��B��������s=�3� �������-�:9�%�?�Ҙ@���<��r5�rw,�%�"��B��i��h����	߽|˽Aú��^��XR��w���ｽ88ϽI��҄���r���k�u%��.�@D7�9�=���@�ݻ>��7�o�*�����#������n��T8�q������#���1���;�@�@���?�2�:�V�2��M)�X����a	�r��h�Xؽ`ŽK���v�������T��6ýO�ս* �T_ ���
�D��v���@(���1�O�9��c?��@���<�,]3�0�%����(S�v6���1�f��L���_�	�1���(��5�y)>��@�v>��$8�W�/��!&�U������������}4潧jѽd���\��7���j����Q��ɽ9�ܽG����GN�S1�'�!�n+���4��	<��d@�r@��;:�+/�a[ ��H�"�����),轐I�� �������-�>9��  �  ^�#�k�(�}�+�t�,���,�ns+���(���#�Du���~H�����ڽ��̽�Ƚ(Ͻ��޽����,�BL������$��~)�%�+�6�,�t,�Y +�(�5a"�S��3��'�j���׽�i˽)ɽ�ѽg�2��9	��)�p����%�*��,��,��Q,�ܿ*��D'�/'!�("���� ��罧�Խ�Jʽ(�ɽSӽ���c<���L�q��I ���&�5v*�	4,���,��$,��O*�Ho&���U[�D�
�f����P�~�ҽ�sɽ�ʽC�ս�.� � ��[���T�!�B�'���*�d],�2�,�A�+��)�!�%��u�@�����e�������Yн��ȽS�˽ˌؽ�����k`�	_�5�"�F>(��:+��z,��,��+�*K)�&�$�U�����9d����-�ݽ0lν^�ȽvIͽ\۽����`Z������#�Z�(���+�ߑ,��,��p+�Ư(���#��q�b��jD�͗ｮ~ڽ��̽*�Ƚ\
Ͻu�޽������H��}���$�K|)�6�+���,��r,��+��(��_"�_����P$�E���׽�b˽Sɽ�ѽ.����5	��%����;�%���)�,�R�,�xO,��*�C'��%!�!�A��D ������Խ�Kʽm�ɽ�Tӽ��b?��aN����lK �;�&�,y*�K7,�E�,��(,��S*��s&����`��
�"����Z�	�ҽ�|ɽϥʽe�սU6�P� ��^������!�D�'���*�N_,�B�,���+���)�9�%�;y�8��܆�����h���cн��Ƚ<�˽Z�ؽ��L��Pd��b���"�^A(��=+��},�5�,�C�+��N)�<�$������}i��󽱟ݽ�wν�Ƚ�TͽT�۽X��T���^�����  �  \������u#���,���5��=���@�]{?� �8�8�,�?�����������6<��𽬛��(�	=!�B�/���:��9@��B@���;��
4���*��Q!�?��ͽ��Y�5��۽YȽ����PZ��Z���g�������Հҽ<e�*'���0	��J�2�v�&�0�Ǐ8�ϴ>�P�@���=��F5��(��H����f��VD�=��9���k{�^g&��4��%=�~�@��)?��`9�31�J�'����^�R
�Є��$��M�ԽGE½+����ݭ�����5��ƽ�:ٽ��*(�=��2��> ��)��3���:��?�8{@���;�XO1���"����
��K�s�hI�C!��������Q+�ٟ7�f�>���@���=�Q�6��.���$�e��T����M�����o%ν��������G��F°�i���G̽�6��������������r#��,�$�5�=�0�@�Ax?���8�R�,���]��ͱ��_��1�~�𽋖�$��8!�'�/��:��6@�L@@�h�;�	4�C�*�P!����	���W��
񽚉۽_�ǽd���6S��ܓ�������}��yҽ�]����9-	��G�+���&��0���8��>���@�m�=��E5�!(�H�����f��
E꽁���;��A��|�"i&��4�'(=��@��,?�d9��1��'���c�xV
����q�齳�Խ�N½`����歽yƮ��=��Hƽ,Aٽ٣*����S��@ �5�)��3�f�:� �?��~@�l�;��S1�<�"���G�eV�2~��S�M+�����=���U+�y�7��?���@�}�=�.�6��	.�ч$����$�K���V������/νu'�������R��
Ͱ���̽�?��������  �  � ��$���#�_�5��G���U�`1_��a�J�Z�c�L���9��%�h��l'�����
�UX�`�)�hV>��uP�O�\�ha��]���R�`C���1�� ���V����ѽ!
���u��d ��_똽����^=��Bg���3����ǽ��ݽU"�����L��޺)��;��nL���Y�Ѻ`���_���V��F�3��#���+����������0���D�7YU��H_�_
a���Z�N�%�=���+��\�(�
�)��e�8ʽ,���̧�'��^×��p�����֪������ν�a����j����&�/�EvA�!^Q���\�aa���]��'R���@�1,�n/�:0����Q�b(�-X#�#�7���J�ҁY���`���_�(W�1�H���7�!�%�������c�jؽ:Xý|�����������O��� ���l��yǯ�Y1����ս�����!��#��5�G��U��._�Sa���Z�Q�L�%�9�%�%�'���!�"��
��R�"�)��Q>�qP�\�\��da�-�]�i�R��]C��1�6 ����x���Mѽ����o�����䘽�����5���_��I,��T�ǽ�}ݽ������c��5�)���;��lL���Y�;�`�}�_���V�J�F��3��#�������������6�0�c�D�?[U��J_��a���Z�2!N���=���+�v`�=�
����6�;ʽE���է����˗�y��0���ݪ�\��ӵν=g���������o�/��xA��`Q��\��da���]�,R���@�l6,��4��5�N���V��-�]#���7���J�}�Y���`���_��*W���H���7��%�W��/��tk�:sؽ}aýI���ĸ��v����Y���
���v���Я��9����ս����  �  ����x���,*��}C��{\���q�����%��؊}���l�)�U���<�!'�)��^���&�mt+��PB��I[�,Xq�l��O&����}�?�m��W���=�[�$���������սR��F%���阽�Z���o��X���$��h���}ɠ�����ɽ����R�"z2�G L�l.d��w�~S��柁�b�x�1�e��oM�W5��V!���2����W�2�9�J��0c��6w��O������	9y�P�f�(�N��E5�|��	I��N꽞�̽L��������ٔ��Ӌ��~��%��}p��}���1���͹�G�ҽ�����j"���:�~^T�cXk�%L|�
��>}��Lcs���]��E�H�-����� ���%�i2:��S��j� |�s	��(���2�s��_�dTF���,��P��� ���߽S2Ľ�G���o�� V���ډ��!��P���F���ܛ�	*���~���bܽx������Z**�d{C�y\��q�'��"$���}���l�s�U���<��'�d��tz�� ��n+�&KB�QD[�kSq�.��u$����}���m�ZW���=�s�$������F�սdM�� ��?䘽�T��i��Q�����/���M �t���4�ɽ�����O��w2���K�Y,d��w��R��C���`�x�t�e�CoM�&5��V!�B �ԃ�����2���J��2c��8w��P������;y�d�f�|�N�EI5�F��M��V�7�̽������b┽�܋�&���&��x������7��kӹ���ҽ�������"�9�:�(aT�b[k��O|���q��,hs�$�]�kE� �-���Ӵ����N%��7:��S�=�j��#|���������s�m_�	WF�^�,� T��� �j�߽r:ĽXP��y���_���䉽c+���Y���O��_国62��"���Niܽ�  �  �U����x�2�-R��-q��腾'ڎ�����t���b��6�m���P��c7�X�&���!��l)�Bn<�|W��.t���nh�������W��A��ـj�/K�~	,��3����P�̽�Y��WI���b��,�����z���x���`y��k���s(���$���2�n@�Y)��=�G�\�w�z��x��"����<��a���.��Cd���G��0��#��"�w�.���D��`�ug}�s\��Y吾J�s�����}��+`�|z@��K"�����d� \½����o���ϓ���h���?y��2z��ց�G
���R������d.ɽ7�^�Y�(���G��g��؁��x��d���B����#��'Kw�+CZ��?�i+���!�q%�l5�w�M�܉j�L���3��`���B}��w&���mt��U�h6���H  �ؽs븽苡�'����Y��Z}���x��g|�sc�� 1��\_��!����.Խ�O���� �2��R�U+q�3煾�؎�4������i`��Z�m�<�P��]7�Z�&�y�!�jf)�2h<��W�:)t�}���2f�������U���?��^~j��K�z,��1�����̽'U��.D���\�������z�i�x�;��[r��o𓽚!�����f,�y=��&� =��\�p�z��w��`����;���`��p.���d���G��0�J�#���"�_�.�"�D�t�`�/i}�r]��z搾��؉����}�*/`� ~@�mO"�����l�od½�������p���!q��OPy�rBz�Sށ�+��DY�������3ɽ<�a���(�!�G��g�Xځ�cz��o������� &���Pw�IZ��?��+���!��v%�5���M���j�l���5������~���'��pt���U�!6���|# �ؽ6�I������c��m}���x�yz|�ll���9��>g��W���5Խ�  �  "x���}���9��+]�j�����X9��菜��|���፾>~��"^�
KB���/� m*�B�2���G�e�z����������fv������Z ����x��1U�#@2�����2ɽh���e���\����Ox�Hgn�f�l���r�π�"3���ݟ��\��?f޽)��{�#��_E��i�����$��^%����z����A���Xs�9T�3�:���,�Ϲ+��8���P���o�b����v��o���]���CW��>9���m�'II��I'���	����Խ�1\��{玽�⁽�t�`�l��m�u�v��M��`��������6Žk��3����.�
5Q�d�t���������C������"���C���h�\�J�{�4��*�{�.��?�B�Z�C�z�\a��o���Rw���򙾫����g&a�Л=������ �cwս���	���퉽:~}���p��Gl���o�(�{��j��'՘�Ո���4ѽbr��]{�#�9��)]�4��r���7��7����z���ߍ�I~�i^�3EB�u�/��f*���2���G�e�����ﱐ�@��at��󁗾���#�x��/U�>2�������ɽ����B���Ǜ���Cx��Zn��l�&�r�Ȁ�F,��2ן�[V��`޽@��ǿ#�d]E�pi����0#���$��b������*A��jXs�T�J�:��,�q�+��8��P�,�o�=����w�����������X���:���m��LI�;M'�c�	���9ݽ��d��	���*끽�t���l���m��v�ZT����������:<Ž��콪��m�.��7Q�E�t����������E��򥚾����F���h���J�Ƕ4�W�*���.�ò?���Z��z��c��Q����x��������
����(a�f�=�`���� �B~ս����.������C�}��p�=Zl�"�o���{��r���ܘ�⏰�:;ѽ�  �  Q�������<� Ia�ق�u��{����m���7��3B���큾��b�#F��#3�a�-��L6���K��j������,�� ̝��R���-���X���}�K�X�S�4�h(��Y�:Ƚz쨽��������,t�s[j��h��n�Rp}��"��Q��d��]2޽�n�O�%�%�H���m�w�������󞾴ܟ��7���z����x�\�X�+|>�:�/���.��5<��4U�
u�̊�b��{���n���ᗾ�@��`�q�&�L��F)�X}
�������r���ڌ�x��v�o�/�h��i�e�r��5������7��W:Ľ^�����0��T���y�����(������q��釕�8S���m�C�N�w8�v�-� �1��oC�#W_����(���-K���T������꓾�����ke��y@��m���<�ԽQ>��(��Tه�=Ty�6�l��Bh��k�hzw��T���ᖽI��^�н`K����R~<��Fa��ׂ��s���l��6���?��T끾z�b�:F��3�z-�eF6�T�K��
j�����f*���ɝ��P��,��@W��y�}���X�6�4�^&��U�.6Ƚ�稽����&���� t��Nj��h��n��b}�����������5,޽�k���%���H�c�m�v������#�ܟ�d7���z����x�.�X�B|>���/���.��6<��5U�|u��̊�`��0|���o��0㗾B����q���L�~J)�6�
���c���畠��⌽l���o�X�h���i��r�u<��M���
���?Ľx����c�0���T���y�H����)������s������V���m���N��8���-�8�1�kuC�}\_�i��O���M��LV��h���\듾1�ine�2|@�`p��� ս�E��00���ᇽfy�z�l��Th�
�k�ŋw��\��/閽H
����н�  �  "x���}���9��+]�j�����X9��菜��|���፾>~��"^�
KB���/� m*�B�2���G�e�z����������fv������Z ����x��1U�#@2�����2ɽh���e���\����Ox�Hgn�f�l���r�π�"3���ݟ��\��?f޽)��{�#��_E��i�����$��^%����z����A���Xs�9T�3�:���,�Ϲ+��8���P���o�b����v��o���]���CW��>9���m�'II��I'���	����Խ�1\��{玽�⁽�t�`�l��m�u�v��M��`��������6Žk��3����.�
5Q�d�t���������C������"���C���h�\�J�{�4��*�{�.��?�B�Z�C�z�\a��o���Rw���򙾫����g&a�Л=������ �cwս���	���퉽:~}���p��Gl���o�(�{��j��'՘�Ո���4ѽbr��]{�#�9��)]�4��r���7��7����z���ߍ�I~�i^�3EB�u�/��f*���2���G�e�����ﱐ�@��at��󁗾���#�x��/U�>2�������ɽ����B���Ǜ���Cx��Zn��l�&�r�Ȁ�F,��2ן�[V��`޽@��ǿ#�d]E�pi����0#���$��b������*A��jXs�T�J�:��,�q�+��8��P�,�o�=����w�����������X���:���m��LI�;M'�c�	���9ݽ��d��	���*끽�t���l���m��v�ZT����������:<Ž��콪��m�.��7Q�E�t����������E��򥚾����F���h���J�Ƕ4�W�*���.�ò?���Z��z��c��Q����x��������
����(a�f�=�`���� �B~ս����.������C�}��p�=Zl�"�o���{��r���ܘ�⏰�:;ѽ�  �  �U����x�2�-R��-q��腾'ڎ�����t���b��6�m���P��c7�X�&���!��l)�Bn<�|W��.t���nh�������W��A��ـj�/K�~	,��3����P�̽�Y��WI���b��,�����z���x���`y��k���s(���$���2�n@�Y)��=�G�\�w�z��x��"����<��a���.��Cd���G��0��#��"�w�.���D��`�ug}�s\��Y吾J�s�����}��+`�|z@��K"�����d� \½����o���ϓ���h���?y��2z��ց�G
���R������d.ɽ7�^�Y�(���G��g��؁��x��d���B����#��'Kw�+CZ��?�i+���!�q%�l5�w�M�܉j�L���3��`���B}��w&���mt��U�h6���H  �ؽs븽苡�'����Y��Z}���x��g|�sc�� 1��\_��!����.Խ�O���� �2��R�U+q�3煾�؎�4������i`��Z�m�<�P��]7�Z�&�y�!�jf)�2h<��W�:)t�}���2f�������U���?��^~j��K�z,��1�����̽'U��.D���\�������z�i�x�;��[r��o𓽚!�����f,�y=��&� =��\�p�z��w��`����;���`��p.���d���G��0�J�#���"�_�.�"�D�t�`�/i}�r]��z搾��؉����}�*/`� ~@�mO"�����l�od½�������p���!q��OPy�rBz�Sށ�+��DY�������3ɽ<�a���(�!�G��g�Xځ�cz��o������� &���Pw�IZ��?��+���!��v%�5���M���j�l���5������~���'��pt���U�!6���|# �ؽ6�I������c��m}���x�yz|�ll���9��>g��W���5Խ�  �  ����x���,*��}C��{\���q�����%��؊}���l�)�U���<�!'�)��^���&�mt+��PB��I[�,Xq�l��O&����}�?�m��W���=�[�$���������սR��F%���阽�Z���o��X���$��h���}ɠ�����ɽ����R�"z2�G L�l.d��w�~S��柁�b�x�1�e��oM�W5��V!���2����W�2�9�J��0c��6w��O������	9y�P�f�(�N��E5�|��	I��N꽞�̽L��������ٔ��Ӌ��~��%��}p��}���1���͹�G�ҽ�����j"���:�~^T�cXk�%L|�
��>}��Lcs���]��E�H�-����� ���%�i2:��S��j� |�s	��(���2�s��_�dTF���,��P��� ���߽S2Ľ�G���o�� V���ډ��!��P���F���ܛ�	*���~���bܽx������Z**�d{C�y\��q�'��"$���}���l�s�U���<��'�d��tz�� ��n+�&KB�QD[�kSq�.��u$����}���m�ZW���=�s�$������F�սdM�� ��?䘽�T��i��Q�����/���M �t���4�ɽ�����O��w2���K�Y,d��w��R��C���`�x�t�e�CoM�&5��V!�B �ԃ�����2���J��2c��8w��P������;y�d�f�|�N�EI5�F��M��V�7�̽������b┽�܋�&���&��x������7��kӹ���ҽ�������"�9�:�(aT�b[k��O|���q��,hs�$�]�kE� �-���Ӵ����N%��7:��S�=�j��#|���������s�m_�	WF�^�,� T��� �j�߽r:ĽXP��y���_���䉽c+���Y���O��_国62��"���Niܽ�  �  � ��$���#�_�5��G���U�`1_��a�J�Z�c�L���9��%�h��l'�����
�UX�`�)�hV>��uP�O�\�ha��]���R�`C���1�� ���V����ѽ!
���u��d ��_똽����^=��Bg���3����ǽ��ݽU"�����L��޺)��;��nL���Y�Ѻ`���_���V��F�3��#���+����������0���D�7YU��H_�_
a���Z�N�%�=���+��\�(�
�)��e�8ʽ,���̧�'��^×��p�����֪������ν�a����j����&�/�EvA�!^Q���\�aa���]��'R���@�1,�n/�:0����Q�b(�-X#�#�7���J�ҁY���`���_�(W�1�H���7�!�%�������c�jؽ:Xý|�����������O��� ���l��yǯ�Y1����ս�����!��#��5�G��U��._�Sa���Z�Q�L�%�9�%�%�'���!�"��
��R�"�)��Q>�qP�\�\��da�-�]�i�R��]C��1�6 ����x���Mѽ����o�����䘽�����5���_��I,��T�ǽ�}ݽ������c��5�)���;��lL���Y�;�`�}�_���V�J�F��3��#�������������6�0�c�D�?[U��J_��a���Z�2!N���=���+�v`�=�
����6�;ʽE���է����˗�y��0���ݪ�\��ӵν=g���������o�/��xA��`Q��\��da���]�,R���@�l6,��4��5�N���V��-�]#���7���J�}�Y���`���_��*W���H���7��%�W��/��tk�:sؽ}aýI���ĸ��v����Y���
���v���Я��9����ս����  �  \������u#���,���5��=���@�]{?� �8�8�,�?�����������6<��𽬛��(�	=!�B�/���:��9@��B@���;��
4���*��Q!�?��ͽ��Y�5��۽YȽ����PZ��Z���g�������Հҽ<e�*'���0	��J�2�v�&�0�Ǐ8�ϴ>�P�@���=��F5��(��H����f��VD�=��9���k{�^g&��4��%=�~�@��)?��`9�31�J�'����^�R
�Є��$��M�ԽGE½+����ݭ�����5��ƽ�:ٽ��*(�=��2��> ��)��3���:��?�8{@���;�XO1���"����
��K�s�hI�C!��������Q+�ٟ7�f�>���@���=�Q�6��.���$�e��T����M�����o%ν��������G��F°�i���G̽�6��������������r#��,�$�5�=�0�@�Ax?���8�R�,���]��ͱ��_��1�~�𽋖�$��8!�'�/��:��6@�L@@�h�;�	4�C�*�P!����	���W��
񽚉۽_�ǽd���6S��ܓ�������}��yҽ�]����9-	��G�+���&��0���8��>���@�m�=��E5�!(�H�����f��
E꽁���;��A��|�"i&��4�'(=��@��,?�d9��1��'���c�xV
����q�齳�Խ�N½`����歽yƮ��=��Hƽ,Aٽ٣*����S��@ �5�)��3�f�:� �?��~@�l�;��S1�<�"���G�eV�2~��S�M+�����=���U+�y�7��?���@�}�=�.�6��	.�ч$����$�K���V������/νu'�������R��
Ͱ���̽�?��������  �  ^�#�k�(�}�+�t�,���,�ns+���(���#�Du���~H�����ڽ��̽�Ƚ(Ͻ��޽����,�BL������$��~)�%�+�6�,�t,�Y +�(�5a"�S��3��'�j���׽�i˽)ɽ�ѽg�2��9	��)�p����%�*��,��,��Q,�ܿ*��D'�/'!�("���� ��罧�Խ�Jʽ(�ɽSӽ���c<���L�q��I ���&�5v*�	4,���,��$,��O*�Ho&���U[�D�
�f����P�~�ҽ�sɽ�ʽC�ս�.� � ��[���T�!�B�'���*�d],�2�,�A�+��)�!�%��u�@�����e�������Yн��ȽS�˽ˌؽ�����k`�	_�5�"�F>(��:+��z,��,��+�*K)�&�$�U�����9d����-�ݽ0lν^�ȽvIͽ\۽����`Z������#�Z�(���+�ߑ,��,��p+�Ư(���#��q�b��jD�͗ｮ~ڽ��̽*�Ƚ\
Ͻu�޽������H��}���$�K|)�6�+���,��r,��+��(��_"�_����P$�E���׽�b˽Sɽ�ѽ.����5	��%����;�%���)�,�R�,�xO,��*�C'��%!�!�A��D ������Խ�Kʽm�ɽ�Tӽ��b?��aN����lK �;�&�,y*�K7,�E�,��(,��S*��s&����`��
�"����Z�	�ҽ�|ɽϥʽe�սU6�P� ��^������!�D�'���*�N_,�B�,���+���)�9�%�;y�8��܆�����h���cн��Ƚ<�˽Z�ؽ��L��Pd��b���"�^A(��=+��},�5�,�C�+��N)�<�$������}i��󽱟ݽ�wν�Ƚ�TͽT�۽X��T���^�����  �  ��?��@�Ҵ<�ru5��y,���"��E��l�W�}����߽�˽̺��g���[����������@Ͻ��㽛����u�`��m�%�q�.�tE7�g�=�<�@�h�>��7���*�G���&�7�����뽢���@����M����#�2�U<�Ҙ@��?�/�:��2�+P)�e�����
����%j�gؽ�Ž/���ƀ������R���3ýI�ս���9] ���
����q���=(��1�e�9��_?���@��<�RX3�4�%����N��,��E(�[������}	��-���(���5�U'>�3�@�Jt>��"8���/��&��}���L��M���l,��aѽ=�������w������H����Ƚ�ܽ{?�q���J�,.��!��j+�5�4�<��`@�@��6:��%/��U ��B��������s=�3� �������-�:9�%�?�Ҙ@���<��r5�rw,�%�"��B��i��h����	߽|˽Aú��^��XR��w���ｽ88ϽI��҄���r���k�u%��.�@D7�9�=���@�ݻ>��7�o�*�����#������n��T8�q������#���1���;�@�@���?�2�:�V�2��M)�X����a	�r��h�Xؽ`ŽK���v�������T��6ýO�ս* �T_ ���
�D��v���@(���1�O�9��c?��@���<�,]3�0�%����(S�v6���1�f��L���_�	�1���(��5�y)>��@�v>��$8�W�/��!&�U������������}4潧jѽd���\��7���j����Q��ɽ9�ܽG����GN�S1�'�!�n+���4��	<��d@�r@��;:�+/�a[ ��H�"�����),轐I�� �������-�>9��  �  ;a�c�^�[U��.F���4���"��B�X��7�G�Խ�)�����,ۡ�?����`������^��uu��,xĽd�ٽ���V�������&���8�d�I���W�-`��`�o�X���I��t6�^J"�ta�G��/����A(��V-�g�A���R�0^��Wa�EU\��P�.�@���.��+���F�����ͽ@��������B��J뗽+���N���X	��W/˽@e������e�zJ��,���>���N�N[�&(a���^���T��C�u�/�m��
�wL��J����_+ ��)4��G���W��*`�v�`�fY�ؑK�k�:�*�(���'����08ܽ��ƽ6@�����l͛��t���$������U@��I��DҽCp�"��6���� �ެ2��ND��S��^��[a��W\���O��4=�M�(�j���	�š�������R�&��:�8�M��G[�B7a��^�kU�1,F�j�4�q�"�Y@�GU�b1콂�Խ�"��9��ҡ�����(X��g���V���m��6qĽ=�ٽs��*�������&���8�i�I���W�`�v�`���X�h�I��q6�G"��]�@���������#�fR-��A���R�,^� Ta��Q\�֑P�g~@�B�.��)�,�W|��b�U�ͽ( ��$��&����B���엽�������d���2˽�iὢ���xh��M�z�,�D�>���N�`R[��,a���^���T��C���/�����hQ�OO�+��D/ �c-4�n�G�1�W��,`�8�`��Y�a�K��:��(�-����	����>ܽq�ƽQH������J֛��}���-��7����H��0���KҽAw�r��i��� �#�2��QD�ʪS�^�,`a��\\���O��:=���(��p�D�	�P�����߭��&�[�:��M��K[��  �  �,��c�	�p��'[�B���(�í�������ڽ�2��)��� ��L͏�����0��,/��C쑽�G��{d��=�Ž�|������M.�O�G�td`�\�t�-��������c{�1ki���Q�h�8�X$�pL�!��~A�B�.��uF��K_�fet�ȹ������a�{�3j�N�R�h�9��� ��
����F;ѽ9����B��Җ�R���函�����8������i��)-���2ν�%��e��(���6��2P���g��z������ ���Iv�l�a��9I��J1����?�tx��:"�hL6���N���f�F�y�����&���v���b��J�?1�u�g���佒bȽF����韽�	��LȊ��?��V����ˎ�i�����p���5|׽}����I�+&��4?��uX���n�L~��*��e�}Ap��Y�c�@��P*�D{��l��I�,'(��3>�+W�@n�U.~��*���{��p�E%[��B�D�(�)��W�����ڽ#,��"�����vŏ�����(��9'���䑽�@��^����Ž;x�0��p���L.�h�G��c`���t��������b{��hi�)�Q��8��$�DH�����<���.��pF�G_�at���������ؐ{��/j�q�R��9��� ��
�����8ѽ|����A���і�g��x懽ʠ���:��f����l���0���6ν�*콜h��+��6��6P���g�Hz�Á� #���Nv���a�?I��O1����-D�B}�?"�bP6�	�N���f���y������&��s�v���b�X�J��1�i��
�7���hȽE���|񟽫���Њ�uH��ۥ��Ԏ�y����#������"�׽!����L�n&��7?�UyX���n�uP~�	-��wj�PGp�C�Y���@��W*�'��rs�FP��-(��9>��0W�<n��2~��  �  gő������C��N�o�TYP��
1���������Mҽ����UX���}��M����
|���x�H�}�#ㅽ腑�����Rv���ڽ e������7��jW�jv�����7ɏ�4���2ǌ�U����h�	L���3�C�$��"�2�+�zu@���[���x�s���V>��'i��J���!���`e��E��'�[����꽑rǽAZ��d���i��}y����y�yy��R.������f˩��Ľ����;	���#��9B�i�a�O�#
�����P���Ӊ���{� _�3<C�<�-���"���#�=�1��I�{�e�	耾^܋��_��wO��ꈾ?5y�m�Z�YG;�ۚ�i��a޽�����������膽��~�3�x��0{����{��C��׳��Ɏν ��j��;�-���L�]-l�H���򹑾8��Q��"�r��qU�1;���(�i�!�A'��8�$GR��ao� 	���b��hÑ��~��+B����o��VP�%1���#���HҽI����Q��pv���3�{�>�x�*�}��ۅ�7������q��[ڽFc�;����7�-jW��
v�?����ȏ�����Rƌ��S����h��L���3���$�"�p�+��p@��[���x�3���6<��-g��z�� ���]e�W�E��'�}�����(pǽ|X���b��ui���y�� �y��{y��À��0������ϩ�FĽ����>	���#�s=B�>�a�BS�a��' ��ճ���Չ�F�{��%_��AC���-�.�"�z�#�ò1��I���e��逾�݋��`��?P���ꈾ}6y���Z��H;�������|#޽ސ��i���7$����
���x�kA{����V���J��
�����ν�&�������-�"�L�1l��������v������#T����r��xU�;";���(���!��G'���8�XMR�fgo�����d���  �  �����Ә��d��nV~�R-[� �7��������&ϽH���ŗ�巇���z��}o��bl�Gq�\�~������C���V��f�׽�c�f����?��%c��ׂ��4���H��/d�����5�����x�<Y��q>�h.���*���5��AL��gj��������#��"������f�r�:O��,�:�ON�AUýe[���������	
v�.�m�%m�<�t��y��eЏ���������Jk彿&�\)��AK���n�R���锾K͛��k��rߓ�6ˆ�f�m�OO���7�c+���,��<�|�U��"u�u��=��)��eᚾT���z����g�_lC��"�0=��ܽ���꟞�|W���A���Cr�yl�J�n��y��H��c���+��K˽gt��<��j4�-W�J�z��㌾����c���R���y��^����Pc��`F�2�?U*�X�0��C���_����P���!䘾����6Ҙ�Gc���S~��*[���7��������� Ͻ ��+���߰��E�z��no��Sl�a8q�oz~�2����=���Q��N�׽�a�3��ˊ?�;%c��ׂ�F4��4H���c��������۷x��Y��m>��-��*� �5��<L�cj����æ���뚾�!��J���m�r�g7O�ƴ,�-8�6K��Rý�Y��笑�2���+
v���m��m���t�S|��~ӏ�N������Np彖)��)�EK���n�l��씾�ϛ�[n��⓾�͆���m��TO��7�Vh+���,�q
<���U�&u����p���)��'⚾��������g��mC�1"�=?�g!ܽ����R����^��)I��USr��l�e�n�q y�[P��ԩ��M	��&˽{������4��0W��z��匾F�������)�����������Wc�hF�j 2�\*�i�0�֢C�L�_�����s显�  �  ���������^�n�ɾ[:��MD��W"e�,9�L��_���V�ֽ�J8�������j�����
��v�½:yݽC�o��7�A��Ap�$��� ���о�Y�˂���F�����zu߾�ľ�+���O���R��T���/ϊ�'���5��GԾd�뾔����������%ܾ��������烾�SU�)�,��O�(��2ͽɷ����yC��hP���7�$WʽJ��Dc
���(�bJP�=���B���*K���8پ�ﾀ;��Ê�����־IM���Ƞ��}��p���n���?���M��J����ܾu�����l���߫�,-Ӿ~~��������u�O�F��!�8���!��Ž菲�r˧��~���!���鬽x���Gӽ}���~t�Ҷ4�g�_����rΧ� Xƾd���_��Z���{`���8�D�;Q������ˇ�6��!�������� �ʾQ�侟���������?]��ɾ 9��C���e��9�{��<�����ֽ�罽�0�����b����������½�sݽ�@������A��@p�ී�����оkY龏���	F��;��]t߾g�ľ�)���M��LP��Ш���̊�\$��3���Ծ���?���]������#ܾ$�������惾�QU��,�fN�C�1ͽyȷ����'D����@�����]Zʽ+�轋e
�8�(�]MP��ှ���6M�� ;پ|��>��|���{��־EP���ˠ�ŀ��C��Rq��OB���O�����^�ܾ���������R�뾒-Ӿ�~��T ���u�0�F��!� ��G(��Ž����jӧ������)����Iɻ��Nӽ�����w�(�4���_�I��;Ч��Yƾ���cb������c���;���;��x ���χ��9�������������7�ʾ��	���  �  '�����G�޾0ž3ܧ�>��j�b�p]8�L2�����t�ٽ�&��4c��8è�k������;����ŽOf�S���W�@���m��H���n���5˾�~�<󾯝��c���پ���^s���Z��ԁ���~����%͚�r�����ξt��9���1�����k�־p~���������S��I,�l��ｿSн@�������H��󦽌���@(���~ͽ)���<�Y|(���N��\~�Tњ�y>���Ծ���Þ��������� �Ѿ���PX�����8]�����K\��������m5׾����7�����t��	6ξp���Wo���s��yE��>!�U����㽡5Ƚõ��᪽����+��8�����`Wֽ�d��~��64���]�j
��"���d���+ܾ�	� ���{��\�=�ȾG���핾�/����}�%M����!��Eƾ"�޾f�����@��ĵ޾�
ž�ڧ�����b��Z8�w/�����Ìٽ����[������ec��[��s4��	�Ž~`ཡP�����@���m��H���n���5˾�~���5��������پ?���q���X���с���~�0��ʚ�������ξ������x/����뾤�־�|��g������S�@H,�$���ｄRн� �������I��_���|����*��Ɓͽ��?��~(���N�`~�.Ӛ��@���Ծ&��S�����������Ѿ
���I[������b�<����^��*���T���6׾��뾿8��r	����s6ξ䷱��o��]s��{E�A!�(��U��<Ƚ�ʵ��骽ᇦ��3��U������^ֽ�k����$:4�D�]���蔤�R���7-ܾB�������`��ɾ��w��3��\�}���祓��$��V	ƾ��޾˗��  �  gk�J�޾�+Ͼ!���	̞�hc���Q]�:o7��u����t�㽝w˽�\���F��ï�`���P��н&�H'�mw�j)?���f��݊�ʘ��0����aӾ�ι�B�۾�>ʾ&�������R����|u���p�\l��+X��n���O���վ������ھ�6Ⱦ��+%���z���O��,������Ĉڽ�@Ž����8����U��ox���^ý��׽����|��%)�zK���u��H��@���ž��ؾ�M��⾌�־z�¾Rʪ�¤��偾�q���s�/��lw���<����Ǿ _ھ&�㾷��Xվ����4~��्�	�k��*C���"���	�y��քҽ�㿽c����ٯ�A��������Fɽpi�{ ���9�3���X�α���图�µ���̾Ήݾ�X�%�߾��о]���������{��p��Jy�N܊�7��u^��.�ξ��޾`i侎�޾Q*Ͼ͉���ʞ�5b��vO]��l7��r�������Gp˽KU��?��$��������H��1н�꽮$�Pu��'?���f�E݊���������aӾ��<�x�۾�=ʾ��������D���*xu���p��i���U�����M��
վH�������ھ5Ⱦ����#����z� �O�s�,���������ڽ/@Ž����粰�KW��^z��Kaý��׽�����~�P()��|K�H�u��J��B��C�ž��ؾP㾭��V�־Z�¾?ͪ������灾j�q��s�q1���y���>���ǾC`ھ��\�ᾕXվ�����~��������k��,C�|�"���	�2��?�ҽ뿽����⯽����4���Nɽq཰~ �c����3�ڷX�v���i盾ĵ��̾)�ݾ�[��߾��о���Y���b�7�{�np�,Ry��ߊ����ua����ξ�޾�  �  �ɾ��žo���e��uҒ�O�|�:X�o9����q������޽�Rͽ&ý�D����Ľ�н/d㽀a��}���$��?���_��ۂ��u��绫�`Ǽ�:�Ǿ�ɾS�¾����~ݟ�:����#u��I`�~S\���i��^��節��&��۰���Ǿ�ɾ�~¾{峾۪���勾�p��3M�
0��o���n�Y	ؽhɽ�X�������ǽNֽ�6뽙����%-��I�	�k�����`��	챾00��R?ɾ�EȾ�F��O����R��twl�T�\�j�^��r�j��^���%���85��Oɾ�4Ⱦ�U��(ح�gƙ������c���B�ɕ'����Z �I��Eҽ��Ž�_��|n½��˽�Kܽ���t	��:��6��xT�A�x�M���o,�������ľ��ɾZ�žW>���������1?�{we�#�[��c��{��㏾Mo��.i����ľ�ɾ�ž�m��Ld��<ђ���|��7X��9����n�s���^�޽�Jͽ�ý�<����Ľ7�н�\��Z�������$�1�?�1�_�qۂ��u������Ǽ�݃Ǿ��ɾ��¾����ܟ�����u�UE`��N\���i�&\��q���;$��������Ǿښɾ�|¾�㳾X����䋾cp�2M��0��n�*��?��ؽzɽ1Y�����
�ǽ�ֽ�9뽂��2!��'-��I�M�k�˜��b��1�2���AɾHHȾ[I���Q�������T��}l���\�x�^�Fr�!l��!�������`6��Pɾ`5Ⱦ=V���ح� Ǚ������c��B�~�'����] ���iMҽj�Ž{h��@w½M�˽Tܽ���jx	�N>�6��{T�~�x�����B.������H�ľP�ɾ,�žnA��ص��"��qF��~e�p�[�"�c�ھ{��揾3r���k����ľ�  �  +����w��<���ܕ�*���Q�r���X��wA��$-�_:�6��a�����mhܽ��ؽek޽�콽���+��p1�w[F�1^���x�V֊��٘����'����-���楾���։��s���W���F���C���N���e�qt���撾���l9��0���Q���t���6���̂���i�d�P�\d:��&�
������H��?�㽗0ڽӭٽY4�3��T������$�c8���M���f�33���������s��}���Ԫ�Rb������NH��Wi���P��PD���E��PU�v�o�����}���̤�ѫ��ы���M���p���|��a���H�[�3�o� �{���n�����߽��ؽއ۽i��$'��`�	��[�+�w?�b�U�*�o�� ��rS��M��Lѩ�-���캨�TG���Q����}���_�+K�u=C�֚I��]��	z������ʜ�6ݧ�F���1v���:��eە�򜇾��r� �X��tA��!-��6�x��P���b�轖_ܽ��ؽ�b޽j���	�|���
n1�WYF�z/^�s�x��Պ��٘��������-���奾�����ԉ�5s���W���F�$�C���N�)�e�r��X䒾S��O7��8���3O��)s��5���˂�[�i���P��b:���&�&��/��6H��U��I1ڽ!�ٽD6⽼��EV����4�$��8���M���f��4������]u��偬�lת��d��i���K���i�D�P�VD���E�UUU�w�o�?������Τ�ҫ�_﫾|���,N���q���|��a�T�H�U�3��� �U��s����.�߽�ٽ�۽X�潫/��d�	��_��
+��?���U�N�o�}��/U��7��pө���������AJ��U��e�}���_�2K�fDC���I�$]��z�u���͜�eߧ��  �  ���F{��>�����D����ir��wc�?eT�q�D�#(4��r#���Ie�������� �
�	�'3�I'���7�W?H���W���f�R�u��g������������P���M���J����g�u�N��9���,�c5*��2�_tD��P\��u�EF���3��ӫ��赐�V?��J����u|�~im��z^��=O�u=?�k�.����V� %�����A1��*/����TK�5�,�kg=��M�E�\�v�k��z��ل����	[��nÑ�BΎ�TW����x�
#_���F��44�*�*���+��7���K���d�X�}�]���ޏ�iϑ�ꋏ��7��?:���mw�oh��uY�� J��9���(����!�Xt�GG�������<�=[�j�!�hF2�B�B�/�R�>�a�2�p�-���;��.x���C��aK��4̌�s���+Ip�*�V���?��/�5�)�I�.���=���S�Psm��ɂ�`�� ���y���	��� �����wgr�-uc�_bT�;�D��$4��n#�����`����x��� �m�	��.�P'�z�7�V<H��W���f���u�2g��U����� ���/P���L��~I���g�3�N�N�9���,�1*�m�2��oD�L\���u�#D��1��񩑾-����=��㧅�Vs|�Ygm��x^�K<O�I<?���.���V�%������2��0�����L��,��i=��M��\���k���z��ۄ�"���<]���ő��Ў��Y��3�x�Z(_���F�:4�+�*�L�+�f�7���K���d�=�}�P^���ߏ�CБ�����L8��;���ow�sqh��xY��J���9��(����%�By�*Q��{����A��_���!�=J2���B�s�R�U�a�8�p�B��Z=���y���E���M���Ό�1���Op�i�V�>�?���/���)���.���=�|�S��xm��˂�t���  �  ��t��i|�6������8������	|�vtt�d#h��fW�C�C��Q0����h���� ��T#�ă4�VH��q[�zJk��v�A}��<���ƀ����Q��� {�»r�*�e�kFT�"�@�BE-����/�����`���%�׻7�N�K�"\^��~m�v�w���}��a���ˀ�*�����Rz�M�p�q�b��Q��4=�>Q*�p�
�˔�T%�fi(�K�:���N�q*a��o�%;y��~�F��-ˀ�ju��k~�o�x�8�n�,;`��M�W�9��x'�����a��K���G+��N>�%R���c�ށq��hz��4�ș���ɀ��U���}��}w���l��b]�	�J�o�6�(�$��������=��?��B.���A��OU�
wf��Os�!u{��������l��,����|��v��j��mZ��4G��n3�51"��K���g��� ��U1���D��hX���h�j�t��f|����T��������_|�|qt� h�cW��C�aM0���P��������M	#�4��QH��m[�Gk���v��>}��;���ŀ�`������{�:�r�K�e�#DT�i�@�B-�d��P����x\�8�%���7��K�X^�{m���w���}�s`��9ʀ��������z���p�N�b�Q�4=�Q*�"p�\
�r��G&��j(�� ;���N��,a���o��=y���~�����̀�iw��Vo~���x���n�@`��M�r�9��}'����Sf�iP�@��K+�R>��'R� �c���q�jjz�M6������ʀ��V����}�ʀw���l�g]���J�W�6�M�$�9��7��
C��D�gG.��A��SU��zf��Rs�#x{����4����À��.����|��v���j�sZ�:G�yt3�A7"�R�4��
m�W� �;[1���D�;mX���h��  �  ?U�(Ld��?s��(���b���P��g����ߐ�A����.��~l�ϓR�$�<��#.���)�4�0���@��X���q�씄�K-���j��\&��.��nن���~�i�o�6�`�w�Q���A�NZ1�E� �V������*���z��F��o��"��_�)��:���J�>NZ�Di��Dx�J��������Ï��ё�����������|��pc��J�5�6�R|+���*��
5�SH���`�S�y��݇�L���ˑ�)+��p@��Kr���y�x�j�x�[�4�L��z<���+��j�_,�U�������=��ӣ������y/�	&@�mP�AO_��=n�L}����󏌾Oݐ�x���)ލ������~t���Z��@C�z�1�	*�8-�x�:���O��*i�N쀾J���̂����Ԏ�� ������^�t���e���V�	XG���6�|-&��Z��0	�DU ������X��{�� ���W$��5�P�E��;U�IId�5=s��'���a���O�����$ސ������,��l���R��<�-.�.�)���0��@��X�ǲq�����d+��i��%���,���؆���~���o���`���Q���A�X1��� �G��"��&#���r��9��S����^�)��:��J��JZ��@i��Ax�����������'ё�����H���֨|�]pc�עJ�F�6��|+�<�*�}5��H���`�'�y��އ����2͑��,��B��t����y���j���[�ʣL��<���+��o�D1�!��;����F������a��v|/��(@��P�GQ_��?n�N}����:����ސ�7���*���𸅾��t���Z�uFC��1��*�� -���:���O�j/i�R���h���e���"֎�4"�����u�t�"�e���V�U\G�_�6��2&��_�l6	�[ �	���c�����,��z\$�5��E��  �  .�B�/Z��St�Cl��k���4Ң��ª�+����h��Q	��(���;Jx�!�[���H�gUC��	L�qga�mr��;��-���$�������y��@f��#����4��=n��T�l�=�y�)�4t�+'	��������-۽�$ٽm3�F���'��]���!���4�&J�ub���}��=��G�� ��$��њ���9���2��y�� �m�I%T�PvE�H�D�4�Q�q�j��5��G���Q������c�����j���Ԏ��g��{Ue���L�z�6��#�������}�Zsٽ�xڽmr�Mv��������9�'��;���Q�c<k�:���������U���n����੾eg��w������bd��M�4�C�Z�G��Y�H�t�F���mv���j��R���H��'���X��Jhw���\��E�:W0���S���Y ����	�ݽ��ؽ��ܽX������U��&�b1.��B�q�Y�}Qt�k��A����Т�{��������f��:��Ж��Ex���[�#�H�kOC��L��aa��l�/9��� ��}"��˾��Bx���d������3��i;n�=�T���=�r�)��q��$	�����k��&۽7ٽ�+�q��$�Z�2�!��4��J�rb�ԧ}��<��-��
��R��#���9��S2��:����m�\%T��vE��D�$�Q���j��6��.���^������d��� ���k���֎��i���Ye�ʪL���6���#���Κ�M��D��J|ٽ9�ڽUz佊}�����q����'�7�;���Q��>k�W���M ���������V����⩾�i��!��ӊ���gd��M�+�C�%�G�HY�b�t���x���l���S��XJ��y���h�����%kw���\�}E�6[0�B����^ �>����ݽi�ؽ+�ܽv��R���Y��*��4.��  �  ��:�I Z���6���~~��EL���Gƾ��ɾ�Tľ;z��gN��H̎�	z�/�b���[�/�f�ǋ�� B��է��$���\ƾ��ɾ�Dľ������Z��vv�¢R��4�����d�8۽
 ˽�&½����>ƽ�2ӽ�5�F7�����(�c�D���e��6���ᮾ���_�Ⱦ@ɾ���-}���g��Z`���p�kc^�Ye]�_�m�KT�����b�������Ⱦ�ɾ
����밾n:���w����i���G�F�+���������+
ս�Lǽ���c���Ǿɽ�ٽWp���S��y�1���N��7r�F��͡��ڴ��þ�ɾ�4Ǿ�ڻ�3�������f����h�l\�`a�
�v�a�����������&þs�ɾ_ Ǿ����Ҩ��L�������]��=�D�#�\~��������Ͻ�NĽ\2���|ý ν�߽9���p��� �ǯ:��Z�����X}��K��FFƾ$�ɾ�Rľx���K���Ɏ�Hz��b�9�[�Ѓf����� ?��Fҧ�]"��xZƾ��ɾ�Bľ����o���X��Ctv��R��~4����}��^��2۽�˽�½�y���7ƽz+ӽ|.罝3������(�=�D���e�O5���욾�ா�����Ⱦ�ɾ�����|���g��A`��#�p��c^��e]�N�m��T��f��c�����ƔȾ	ɾ���P�(<���y����i���G���+�4 �Z��L��Rս�Uǽ���������ɽ�ٽ�v�ך�����1�0 O��9r�z��YΡ�jܴ��þ �ɾ7Ǿ*ݻ�	�������i����h��\�ra�ǻv����#��Ί��s(þ
�ɾ�!Ǿ�������AM��h���v�]�h�=���#�{��v���])�u�Ͻ�XĽ�<��Ɔý�ν��߽�����s�0!��  �  OT9�n�_�ھ��?���깾Bо�m߾�e�8޾R�;y��О�cމ�}Ex�:)p�%�|���;���b���
Ҿ�eྡྷE�d�ܾl�˾�]���u���^��XsV���1��/�������޽�AȽ�_���f�����e��W�����ӽ*h�&�
��4$�W6E��*n����𨾽���GI־�Q���㾉�پ>�ƾ�ா>���S��hBs�cr�䮂��Ԕ��'���"ľ��׾�⾪� ؾv{ľ�Ы�cݑ�]+s�a[I��w'��4��
�`cֽ�s½;�',��x䰽!��7ƽj�۽�����p��R.�[�Q��w}�����e���kɾBa۾��㾛_��Ծ� ��*����4��m���p��Tv�Lꇾ�:���P��Ii˾ �ܾ}=�#��,\Ҿš���$��{��#ed��.=�&������l�^�ν쁽��J��#���S������K�̽!�չ�@��sQ9��_������=���鹾�@оjl߾ d�H޾�;���J͞�Yۉ�?x��"p�|�|�������_���ҾmcྌC侞�ܾ��˾U\��{t���]��iqV���1��-�������޽<ȽWY��`���2������o�ӽaｺ�
��1$�H3E��'n�M�������]H־�P�X���پߟƾ�ா>���S���Bs�	r�[���UՔ�N(���#ľ��׾3���㾑ؾ	}ľ]ҫ�5ߑ�;/s�t_I�;|'�P9���^lֽ�|½����4���창�(��!>ƽ��۽����:s�U.���Q��y}�򔗾Ί���lɾ!c۾���bᾇԾy��O����7���s�
�p�/[v�C퇾�=��]S��pk˾��ܾ?侁��d]Ҿ좼��%��F|���gd��1=����~��.u�x�νp����T��廯�囲������̽ )�t��z���  �  �z:�y{e�P�������/�ƾ�߾�0�i������c�ݾ��ľ峩�`����]����}�3ᅾ ��h����zʾ��⾘��t���%C���ھdO���񢾵���J[��22�b���1��~�Խ�����z����7����T��˘����ɽ���.�#��G���u�m���Z����Ͼf��g}������Z��N�վ���TS��j��c����������f����z��Ӿ���S���H��7��іҾ靶��5��~{��iL�ʠ&�=�	�ڰ齷̽�B��W6��̦��w��`J���󻽿�ѽ�������9.�zV�񏃾����\��#0ؾ=��i����z���b;�z�����1Q��B.~��K���`��]ئ�X����+۾GY�׿��io�"V�K�ɾJɬ�ɷ��f�j�O�>�������޽��Ľ;t��Ƕ���Z���	��$��n;½b3۽gO��.���w:��xe�-�������ƾ��߾]/��������ݾ	�ľ���C���LZ����}��݅����*����wʾ3����J���LA�T�ھN���𢾪���J[��02�6��4-��H�Խ�񽽐t��	맽Z����M�������zɽ��彴*��#��G�!�u�'��xY���Ͼ�澡|��P��������վ���<S��"j������g��j��� ����{���Ӿ���HT���I�����`�Ҿ�����7��܁{��mL���&���	���齕&̽^K���>��jԦ�����Q������'�ѽb�񽧊�+<.��V�-���O�������1ؾ,��Ak��v��I���e;.~��d����T���4~��N���c��%ۦ�։��.۾$[�l����p�SW�h�ɾiʬ������j�T�>������޽��Ľy}��=���od��������C½,;۽vV��U���  �  35;�*�g�}ݎ�C�A˾���۝��͔��I���r��Zɾ���c����酾'H��&���~Y������g�Ͼr辁���g�����I]��ľ���)���]��2�k�� ��y�ѽ徺��T���褽�����<��kd���Rƽ���7�"�"���H�^�x�����3���ԾA���������o�!J۾����社ZE��5��c��Gd��p$���ݼ�,lؾ�ﾋ���������̼׾@��������~�Z�M���&������潓�ȽW�����2ɣ�,q���'��'���t�ν+@�����.���W�Uo��^����Z���ݾ��a��|#�����$�Ҿ�����ٜ������}��T΄�_��$���1<ƾs��Ǳ���i������\$�vξ�[������lm��?������ �Ө۽gT���D�������Z��s����ۮ�1��3ؽ1��@Z�o2;���g�\܎�,מּ�?˾}��n������G���p�>Xɾ)���?���7慾�D�����V��_���S~Ͼ:o�� ��Qe������[ྸ�ľ������]�	�2�=��a��D�ѽ6����N��V⤽Ē���5��S]���Kƽ��|4���"���H���x�S����1��ܵԾ[����������I۾�����椾eE��d��fc���d��%���޼�mؾ� ﾴ�������y��[�׾�������~�\�M�Ω&�#��M��e�Ƚ���#���ѣ�y��V/��¸�ٯνF�����.�a�W��p������P\����ݾ����
&�����9�Ҿ���Cݜ�5������ф�b��🪾�>ƾ��ྦ����k��7����%�5wξ�\�����Rom��?�3���� ���۽%]��N�����d������䮽����:ؽ0��`]��  �  �z:�y{e�P�������/�ƾ�߾�0�i������c�ݾ��ľ峩�`����]����}�3ᅾ ��h����zʾ��⾘��t���%C���ھdO���񢾵���J[��22�b���1��~�Խ�����z����7����T��˘����ɽ���.�#��G���u�m���Z����Ͼf��g}������Z��N�վ���TS��j��c����������f����z��Ӿ���S���H��7��іҾ靶��5��~{��iL�ʠ&�=�	�ڰ齷̽�B��W6��̦��w��`J���󻽿�ѽ�������9.�zV�񏃾����\��#0ؾ=��i����z���b;�z�����1Q��B.~��K���`��]ئ�X����+۾GY�׿��io�"V�K�ɾJɬ�ɷ��f�j�O�>�������޽��Ľ;t��Ƕ���Z���	��$��n;½b3۽gO��.���w:��xe�-�������ƾ��߾]/��������ݾ	�ľ���C���LZ����}��݅����*����wʾ3����J���LA�T�ھN���𢾪���J[��02�6��4-��H�Խ�񽽐t��	맽Z����M�������zɽ��彴*��#��G�!�u�'��xY���Ͼ�澡|��P��������վ���<S��"j������g��j��� ����{���Ӿ���HT���I�����`�Ҿ�����7��܁{��mL���&���	���齕&̽^K���>��jԦ�����Q������'�ѽb�񽧊�+<.��V�-���O�������1ؾ,��Ak��v��I���e;.~��d����T���4~��N���c��%ۦ�։��.۾$[�l����p�SW�h�ɾiʬ������j�T�>������޽��Ľy}��=���od��������C½,;۽vV��U���  �  OT9�n�_�ھ��?���깾Bо�m߾�e�8޾R�;y��О�cމ�}Ex�:)p�%�|���;���b���
Ҿ�eྡྷE�d�ܾl�˾�]���u���^��XsV���1��/�������޽�AȽ�_���f�����e��W�����ӽ*h�&�
��4$�W6E��*n����𨾽���GI־�Q���㾉�پ>�ƾ�ா>���S��hBs�cr�䮂��Ԕ��'���"ľ��׾�⾪� ؾv{ľ�Ы�cݑ�]+s�a[I��w'��4��
�`cֽ�s½;�',��x䰽!��7ƽj�۽�����p��R.�[�Q��w}�����e���kɾBa۾��㾛_��Ծ� ��*����4��m���p��Tv�Lꇾ�:���P��Ii˾ �ܾ}=�#��,\Ҿš���$��{��#ed��.=�&������l�^�ν쁽��J��#���S������K�̽!�չ�@��sQ9��_������=���鹾�@оjl߾ d�H޾�;���J͞�Yۉ�?x��"p�|�|�������_���ҾmcྌC侞�ܾ��˾U\��{t���]��iqV���1��-�������޽<ȽWY��`���2������o�ӽaｺ�
��1$�H3E��'n�M�������]H־�P�X���پߟƾ�ா>���S���Bs�	r�[���UՔ�N(���#ľ��׾3���㾑ؾ	}ľ]ҫ�5ߑ�;/s�t_I�;|'�P9���^lֽ�|½����4���창�(��!>ƽ��۽����:s�U.���Q��y}�򔗾Ί���lɾ!c۾���bᾇԾy��O����7���s�
�p�/[v�C퇾�=��]S��pk˾��ܾ?侁��d]Ҿ좼��%��F|���gd��1=����~��.u�x�νp����T��廯�囲������̽ )�t��z���  �  ��:�I Z���6���~~��EL���Gƾ��ɾ�Tľ;z��gN��H̎�	z�/�b���[�/�f�ǋ�� B��է��$���\ƾ��ɾ�Dľ������Z��vv�¢R��4�����d�8۽
 ˽�&½����>ƽ�2ӽ�5�F7�����(�c�D���e��6���ᮾ���_�Ⱦ@ɾ���-}���g��Z`���p�kc^�Ye]�_�m�KT�����b�������Ⱦ�ɾ
����밾n:���w����i���G�F�+���������+
ս�Lǽ���c���Ǿɽ�ٽWp���S��y�1���N��7r�F��͡��ڴ��þ�ɾ�4Ǿ�ڻ�3�������f����h�l\�`a�
�v�a�����������&þs�ɾ_ Ǿ����Ҩ��L�������]��=�D�#�\~��������Ͻ�NĽ\2���|ý ν�߽9���p��� �ǯ:��Z�����X}��K��FFƾ$�ɾ�Rľx���K���Ɏ�Hz��b�9�[�Ѓf����� ?��Fҧ�]"��xZƾ��ɾ�Bľ����o���X��Ctv��R��~4����}��^��2۽�˽�½�y���7ƽz+ӽ|.罝3������(�=�D���e�O5���욾�ா�����Ⱦ�ɾ�����|���g��A`��#�p��c^��e]�N�m��T��f��c�����ƔȾ	ɾ���P�(<���y����i���G���+�4 �Z��L��Rս�Uǽ���������ɽ�ٽ�v�ך�����1�0 O��9r�z��YΡ�jܴ��þ �ɾ7Ǿ*ݻ�	�������i����h��\�ra�ǻv����#��Ί��s(þ
�ɾ�!Ǿ�������AM��h���v�]�h�=���#�{��v���])�u�Ͻ�XĽ�<��Ɔý�ν��߽�����s�0!��  �  .�B�/Z��St�Cl��k���4Ң��ª�+����h��Q	��(���;Jx�!�[���H�gUC��	L�qga�mr��;��-���$�������y��@f��#����4��=n��T�l�=�y�)�4t�+'	��������-۽�$ٽm3�F���'��]���!���4�&J�ub���}��=��G�� ��$��њ���9���2��y�� �m�I%T�PvE�H�D�4�Q�q�j��5��G���Q������c�����j���Ԏ��g��{Ue���L�z�6��#�������}�Zsٽ�xڽmr�Mv��������9�'��;���Q�c<k�:���������U���n����੾eg��w������bd��M�4�C�Z�G��Y�H�t�F���mv���j��R���H��'���X��Jhw���\��E�:W0���S���Y ����	�ݽ��ؽ��ܽX������U��&�b1.��B�q�Y�}Qt�k��A����Т�{��������f��:��Ж��Ex���[�#�H�kOC��L��aa��l�/9��� ��}"��˾��Bx���d������3��i;n�=�T���=�r�)��q��$	�����k��&۽7ٽ�+�q��$�Z�2�!��4��J�rb�ԧ}��<��-��
��R��#���9��S2��:����m�\%T��vE��D�$�Q���j��6��.���^������d��� ���k���֎��i���Ye�ʪL���6���#���Κ�M��D��J|ٽ9�ڽUz佊}�����q����'�7�;���Q��>k�W���M ���������V����⩾�i��!��ӊ���gd��M�+�C�%�G�HY�b�t���x���l���S��XJ��y���h�����%kw���\�}E�6[0�B����^ �>����ݽi�ؽ+�ܽv��R���Y��*��4.��  �  ?U�(Ld��?s��(���b���P��g����ߐ�A����.��~l�ϓR�$�<��#.���)�4�0���@��X���q�씄�K-���j��\&��.��nن���~�i�o�6�`�w�Q���A�NZ1�E� �V������*���z��F��o��"��_�)��:���J�>NZ�Di��Dx�J��������Ï��ё�����������|��pc��J�5�6�R|+���*��
5�SH���`�S�y��݇�L���ˑ�)+��p@��Kr���y�x�j�x�[�4�L��z<���+��j�_,�U�������=��ӣ������y/�	&@�mP�AO_��=n�L}����󏌾Oݐ�x���)ލ������~t���Z��@C�z�1�	*�8-�x�:���O��*i�N쀾J���̂����Ԏ�� ������^�t���e���V�	XG���6�|-&��Z��0	�DU ������X��{�� ���W$��5�P�E��;U�IId�5=s��'���a���O�����$ސ������,��l���R��<�-.�.�)���0��@��X�ǲq�����d+��i��%���,���؆���~���o���`���Q���A�X1��� �G��"��&#���r��9��S����^�)��:��J��JZ��@i��Ax�����������'ё�����H���֨|�]pc�עJ�F�6��|+�<�*�}5��H���`�'�y��އ����2͑��,��B��t����y���j���[�ʣL��<���+��o�D1�!��;����F������a��v|/��(@��P�GQ_��?n�N}����:����ސ�7���*���𸅾��t���Z�uFC��1��*�� -���:���O�j/i�R���h���e���"֎�4"�����u�t�"�e���V�U\G�_�6��2&��_�l6	�[ �	���c�����,��z\$�5��E��  �  ��t��i|�6������8������	|�vtt�d#h��fW�C�C��Q0����h���� ��T#�ă4�VH��q[�zJk��v�A}��<���ƀ����Q��� {�»r�*�e�kFT�"�@�BE-����/�����`���%�׻7�N�K�"\^��~m�v�w���}��a���ˀ�*�����Rz�M�p�q�b��Q��4=�>Q*�p�
�˔�T%�fi(�K�:���N�q*a��o�%;y��~�F��-ˀ�ju��k~�o�x�8�n�,;`��M�W�9��x'�����a��K���G+��N>�%R���c�ށq��hz��4�ș���ɀ��U���}��}w���l��b]�	�J�o�6�(�$��������=��?��B.���A��OU�
wf��Os�!u{��������l��,����|��v��j��mZ��4G��n3�51"��K���g��� ��U1���D��hX���h�j�t��f|����T��������_|�|qt� h�cW��C�aM0���P��������M	#�4��QH��m[�Gk���v��>}��;���ŀ�`������{�:�r�K�e�#DT�i�@�B-�d��P����x\�8�%���7��K�X^�{m���w���}�s`��9ʀ��������z���p�N�b�Q�4=�Q*�"p�\
�r��G&��j(�� ;���N��,a���o��=y���~�����̀�iw��Vo~���x���n�@`��M�r�9��}'����Sf�iP�@��K+�R>��'R� �c���q�jjz�M6������ʀ��V����}�ʀw���l�g]���J�W�6�M�$�9��7��
C��D�gG.��A��SU��zf��Rs�#x{����4����À��.����|��v���j�sZ�:G�yt3�A7"�R�4��
m�W� �;[1���D�;mX���h��  �  ���F{��>�����D����ir��wc�?eT�q�D�#(4��r#���Ie�������� �
�	�'3�I'���7�W?H���W���f�R�u��g������������P���M���J����g�u�N��9���,�c5*��2�_tD��P\��u�EF���3��ӫ��赐�V?��J����u|�~im��z^��=O�u=?�k�.����V� %�����A1��*/����TK�5�,�kg=��M�E�\�v�k��z��ل����	[��nÑ�BΎ�TW����x�
#_���F��44�*�*���+��7���K���d�X�}�]���ޏ�iϑ�ꋏ��7��?:���mw�oh��uY�� J��9���(����!�Xt�GG�������<�=[�j�!�hF2�B�B�/�R�>�a�2�p�-���;��.x���C��aK��4̌�s���+Ip�*�V���?��/�5�)�I�.���=���S�Psm��ɂ�`�� ���y���	��� �����wgr�-uc�_bT�;�D��$4��n#�����`����x��� �m�	��.�P'�z�7�V<H��W���f���u�2g��U����� ���/P���L��~I���g�3�N�N�9���,�1*�m�2��oD�L\���u�#D��1��񩑾-����=��㧅�Vs|�Ygm��x^�K<O�I<?���.���V�%������2��0�����L��,��i=��M��\���k���z��ۄ�"���<]���ő��Ў��Y��3�x�Z(_���F�:4�+�*�L�+�f�7���K���d�=�}�P^���ߏ�CБ�����L8��;���ow�sqh��xY��J���9��(����%�By�*Q��{����A��_���!�=J2���B�s�R�U�a�8�p�B��Z=���y���E���M���Ό�1���Op�i�V�>�?���/���)���.���=�|�S��xm��˂�t���  �  +����w��<���ܕ�*���Q�r���X��wA��$-�_:�6��a�����mhܽ��ؽek޽�콽���+��p1�w[F�1^���x�V֊��٘����'����-���楾���։��s���W���F���C���N���e�qt���撾���l9��0���Q���t���6���̂���i�d�P�\d:��&�
������H��?�㽗0ڽӭٽY4�3��T������$�c8���M���f�33���������s��}���Ԫ�Rb������NH��Wi���P��PD���E��PU�v�o�����}���̤�ѫ��ы���M���p���|��a���H�[�3�o� �{���n�����߽��ؽއ۽i��$'��`�	��[�+�w?�b�U�*�o�� ��rS��M��Lѩ�-���캨�TG���Q����}���_�+K�u=C�֚I��]��	z������ʜ�6ݧ�F���1v���:��eە�򜇾��r� �X��tA��!-��6�x��P���b�轖_ܽ��ؽ�b޽j���	�|���
n1�WYF�z/^�s�x��Պ��٘��������-���奾�����ԉ�5s���W���F�$�C���N�)�e�r��X䒾S��O7��8���3O��)s��5���˂�[�i���P��b:���&�&��/��6H��U��I1ڽ!�ٽD6⽼��EV����4�$��8���M���f��4������]u��偬�lת��d��i���K���i�D�P�VD���E�UUU�w�o�?������Τ�ҫ�_﫾|���,N���q���|��a�T�H�U�3��� �U��s����.�߽�ٽ�۽X�潫/��d�	��_��
+��?���U�N�o�}��/U��7��pө���������AJ��U��e�}���_�2K�fDC���I�$]��z�u���͜�eߧ��  �  �ɾ��žo���e��uҒ�O�|�:X�o9����q������޽�Rͽ&ý�D����Ľ�н/d㽀a��}���$��?���_��ۂ��u��绫�`Ǽ�:�Ǿ�ɾS�¾����~ݟ�:����#u��I`�~S\���i��^��節��&��۰���Ǿ�ɾ�~¾{峾۪���勾�p��3M�
0��o���n�Y	ؽhɽ�X�������ǽNֽ�6뽙����%-��I�	�k�����`��	챾00��R?ɾ�EȾ�F��O����R��twl�T�\�j�^��r�j��^���%���85��Oɾ�4Ⱦ�U��(ح�gƙ������c���B�ɕ'����Z �I��Eҽ��Ž�_��|n½��˽�Kܽ���t	��:��6��xT�A�x�M���o,�������ľ��ɾZ�žW>���������1?�{we�#�[��c��{��㏾Mo��.i����ľ�ɾ�ž�m��Ld��<ђ���|��7X��9����n�s���^�޽�Jͽ�ý�<����Ľ7�н�\��Z�������$�1�?�1�_�qۂ��u������Ǽ�݃Ǿ��ɾ��¾����ܟ�����u�UE`��N\���i�&\��q���;$��������Ǿښɾ�|¾�㳾X����䋾cp�2M��0��n�*��?��ؽzɽ1Y�����
�ǽ�ֽ�9뽂��2!��'-��I�M�k�˜��b��1�2���AɾHHȾ[I���Q�������T��}l���\�x�^�Fr�!l��!�������`6��Pɾ`5Ⱦ=V���ح� Ǚ������c��B�~�'����] ���iMҽj�Ž{h��@w½M�˽Tܽ���jx	�N>�6��{T�~�x�����B.������H�ľP�ɾ,�žnA��ص��"��qF��~e�p�[�"�c�ھ{��揾3r���k����ľ�  �  gk�J�޾�+Ͼ!���	̞�hc���Q]�:o7��u����t�㽝w˽�\���F��ï�`���P��н&�H'�mw�j)?���f��݊�ʘ��0����aӾ�ι�B�۾�>ʾ&�������R����|u���p�\l��+X��n���O���վ������ھ�6Ⱦ��+%���z���O��,������Ĉڽ�@Ž����8����U��ox���^ý��׽����|��%)�zK���u��H��@���ž��ؾ�M��⾌�־z�¾Rʪ�¤��偾�q���s�/��lw���<����Ǿ _ھ&�㾷��Xվ����4~��्�	�k��*C���"���	�y��քҽ�㿽c����ٯ�A��������Fɽpi�{ ���9�3���X�α���图�µ���̾Ήݾ�X�%�߾��о]���������{��p��Jy�N܊�7��u^��.�ξ��޾`i侎�޾Q*Ͼ͉���ʞ�5b��vO]��l7��r�������Gp˽KU��?��$��������H��1н�꽮$�Pu��'?���f�E݊���������aӾ��<�x�۾�=ʾ��������D���*xu���p��i���U�����M��
վH�������ھ5Ⱦ����#����z� �O�s�,���������ڽ/@Ž����粰�KW��^z��Kaý��׽�����~�P()��|K�H�u��J��B��C�ž��ؾP㾭��V�־Z�¾?ͪ������灾j�q��s�q1���y���>���ǾC`ھ��\�ᾕXվ�����~��������k��,C�|�"���	�2��?�ҽ뿽����⯽����4���Nɽq཰~ �c����3�ڷX�v���i盾ĵ��̾)�ݾ�[��߾��о���Y���b�7�{�np�,Ry��ߊ����ua����ξ�޾�  �  '�����G�޾0ž3ܧ�>��j�b�p]8�L2�����t�ٽ�&��4c��8è�k������;����ŽOf�S���W�@���m��H���n���5˾�~�<󾯝��c���پ���^s���Z��ԁ���~����%͚�r�����ξt��9���1�����k�־p~���������S��I,�l��ｿSн@�������H��󦽌���@(���~ͽ)���<�Y|(���N��\~�Tњ�y>���Ծ���Þ��������� �Ѿ���PX�����8]�����K\��������m5׾����7�����t��	6ξp���Wo���s��yE��>!�U����㽡5Ƚõ��᪽����+��8�����`Wֽ�d��~��64���]�j
��"���d���+ܾ�	� ���{��\�=�ȾG���핾�/����}�%M����!��Eƾ"�޾f�����@��ĵ޾�
ž�ڧ�����b��Z8�w/�����Ìٽ����[������ec��[��s4��	�Ž~`ཡP�����@���m��H���n���5˾�~���5��������پ?���q���X���с���~�0��ʚ�������ξ������x/����뾤�־�|��g������S�@H,�$���ｄRн� �������I��_���|����*��Ɓͽ��?��~(���N�`~�.Ӛ��@���Ծ&��S�����������Ѿ
���I[������b�<����^��*���T���6׾��뾿8��r	����s6ξ䷱��o��]s��{E�A!�(��U��<Ƚ�ʵ��骽ᇦ��3��U������^ֽ�k����$:4�D�]���蔤�R���7-ܾB�������`��ɾ��w��3��\�}���祓��$��V	ƾ��޾˗��  �  XpF���@�J�0������ ��Mо,���$у�?�S���-�I���� �����޽�2۽�u���H�2����4���]����Ư��Z�ھ�,�ED��4�X�B��&F���=�D@,�yY�WR���^־p��z���
ʾ#�龣�
��m"�7�l�C���E��C<�֌)��~��M��U��k���A�t��qE���#��N�����彁oܽ��۽p0�.��{�	�uw �AA��n�k���c������k��'���:�PAE�b�D��8���$��g��V�k�̾�ӻ�������ҾQ���ѱ���)��Z<�g�E���C���6���!�z	�� ྋ3��7C���7c�7�8�8�����@񽣐�S۽��ݽ��:�����*�N�N���������8˾�k��6�Q.��H?��[F�*�A�"�2�mA�������žd`����¾@�ݾ��!��x�0�h�@�IoF���@���0����$� ��Lо���σ�t�S�{�-����>� �p��.޽�*۽�m���E�L��c�4��]�{���i���<�ھ�,�WD�-�4�R�B��&F�W�=��?,��X�uP���\־�m������ʾJ��9�
�7l"��7�.�C���E��B<��)��}�2L�T��]�����t�0pE���#�j��������1pܽ5�۽p2佴0��&�	�wy ��A�֔n�����#������~��8'��:��BE�ңD���8�-�$�~i�Z�̾�ֻ�� ��W�Ҿ�������p�)�w[<���E�%�C��6���!��	�R�-4��D���9c���8�s����UH�Ϙ�h[۽�ݽ��1������*�ƮN�ŉ�������:˾�m��6�$R.�J?�]F���A���2�YC����J���!ž�d���þ�ݾO������0���@��  �  ��@��;�O�+�,���d��y�̾|��M8���%T��;/���?F������Y�߽�佃�󽝣�C ��h6��^�Rԉ��n��(�־|��#���/�77=�TW@��q8��}'��y�XL���Ѿ�����o����ž��bP�b�0�1�#>��?�|�6�t�$����VZ��S��7���	t�PxF�ys%�e[����>=�>�ཝR���b���J��o"��8B��Dn�w��l���B�b?��"�!E5��|?���>���3�:z ���	���!Ⱦ����5��
sξ������4%���6���?�\>�^�1�������X�۾@İ��F��>Mc��2:����m�����潜�߽��v�������A�+��jO����� ���Ǿ����M��)���9�?�@��:<��-�R�vU��ܾ���_���=��E�ؾn���Ď��+��;��@��;���+�����c��T�̾L��7���"T�m8/�\��B���!��o�߽Y��,��A��O��f6��^��Ӊ��n���־���#���/�/7=�*W@��q8��|'��x�xJ��ҵѾ~���*m����ž2���N����1��!>���?�p�6���$����X뾉R��r6�� t��vF�|r%��Z�p���H=�����S���	����K��q"��:B��Gn��x��*���3�s@�,�"�dF5��}?�!�>�4�3��{ �3�	�C��8�Ⱦ�"���8���uξ)�����5%��6���?��>���1������ʻ۾�İ��G���Oc�t5:�N���q�`�����߽]"�����������+�nO�j�������Ǿ_���N�:�)���9���@�i<<���-�9�wW�$�ܾ�������B���ؾ����a����+��;��  �  �0���+��b��W�0��0þVf���=��,W�[-5�8b�l�
������� ����z.�c*�M5!���;��1`��#���̦���˾Q��������!���-�U0�GP)��C�����i�z�ľ��������I�վ�-�����q#�L].�x0�$(��~��V��޾����씾��s�>�J���+�����B�L���!~�f��a���������l")���F�S�n�����
����~پ%���h�E�&��/��/�j
%�I�����1WپrU��ß��������CH��a�:<�<�'�"0��m.�p�#����p��iо/���t5���d�_?��#�q��FW�����D�)��C���3	�n�Z�1�:�R�[�~��ћ�达�v羐	��{���*�T�0���,�*��q�E�Uξ)����]���Գ��ʾ���1�$�Z�+�ە0��+�9b�W��.쾞/þ#e���<��4)W�.*5��^���
�������a����*��&�02!��;��/`�#��v̦�r�˾D��������!���-��T0��O)�WC�˨��g�P�ľ����g�������վ�*������o#�\.�Y0��"(�	~�V�,޾͏��{딾��s��J���+�@��aB�X����~��_�����d��l$)�O�F��n����ā����پ4��j���&�a�/�	/��%�������HZپ{X����������\���lJ��b��<���'��0�0n.���#���#q���iо꟪�n6����d�b?�~�#�>��Z[�4��jM���ｻ���7	�P�2���R���~�Cӛ��龾gx羈	��|��*���0�,�,�����r�fI�Yξ;����a���س�9�ʾ��G3�w%���+��  �  ���h����n����%ؾ��������N2���3`�B�<�*�}����u��ȗ�^���w�SF�!P/�J&H���g���8�ڒ��=�߾�y �5��`��.��n���R�)�̾O��ʛ�� t���V�����t�޾�Z �����/��"���E�a����̾����~���x��SU�#�9��$����	�T`����"��{��"�A�6�h�Q��Pt� ʏ��L���Tɾ��H���x�&^�����D�K%�����¾�Y����������׮�hTɾJF꾄����@|��v���Q:��n��¾���<���l�k�XMK���1�����ҋ��� *���
�(�5Y(��%?�Ex\��؀�V��3���gԾ~���j
�~������S��X��
�׾gv��f���+霾�2��x�����Ӿ���F�
�������g����*����$ؾ����S����0���0`��B���*������+��s�����s��B��L/�g#H�B�g�7���젾~����߾�y �)��E�������eR�����̾M��t���}q��CT��e�����޾oY ��������$���D�ɰ�\�̾L����}��J�x��RU�/�9�\$����	��`���#��|�~"�<�6���Q��St��ˏ�;N��iVɾ3��i���y�s_����cF��&�����¾�\��j�������ڮ��VɾH�;������|��v�0��:� o㾐¾����T���!�k��PK�:�1�� �j��K��s���.���Z�,](��)?��{\��ڀ�����4��9iԾY���k
������b����F\��Ɖ׾Bz��Nä�
휾�6�������Ӿ �����
�����  �  �n���������ܾ�{ž����ٚ��P��m?t���Y���B�A/�h4 �v�|~�����
#���2��\G��J_�R�z���������ܳ�U�ʾdh� ����\ �������7侟�ʾ�l�������z��U��������������,>پIG����e��3�������Ծ�ѽ������������j���Q���;��)��z�}{����b���'��U9���N�	�g�K��R���Y���9J��^Ҿ�k�h����<�� �od�ܾP���7v���7���`������{ǘ�����՜Ǿ[��FQ���� �� �_�����9;�P���G��$�����}��$b���I�s5���$�n����Px�3��9-�r!@��V��q�����ZĘ�,���[�¾� ھ�����&}�����˶�+tӾ�߸��.���Đ�3�������I)��k�о�K�
J���m�Z������Ȁܾ�zž`��Gؚ�wO��Y<t�4�Y��}B�/� 0 ����y���7#���2��XG�kG_���z�����4��vܳ���ʾ(h�ƿ��b\ �O�����6�2�ʾ�j������Xx�������S��������;پ�D�I���d�2��֧�?�Ծfн�����������j���Q��;�ҁ)��z��{�7��c�?�'�oW9���N�Th��L��м�����L��`Ҿ&n�ƾ���=�'
 �6g��ܾ6���y���:��Bc��B����ɘ�������Ǿɐ�eR��d� �8� ������㾶9;�Q���H��bᎾ��}�}(b���I��5�=�$��r�ƞ�}�����"-��%@���V�q�T����Ř�������¾�ھv������g~�a����뾀wӾM㸾,2��uȐ�ދ�������S��N�оTN�GL���  �  ؆վ�վ�Ͼɫž 	���V��I	���˗�	��9��u�f�TFO�^_<�N0��,�^K2��@�+T��l�b���Î��Q��}����簾���cȾ�sѾ.G־�{ԾC7˾�t���㧾 ���ns�E�o���|��<���螾���:�ľ�FѾDc־GLԾ�̾A������퇪��N��)������@/w�qx^��XH�*z7�Q.�b�-��6��)F���[��bt�Ұ��⫒����WD���ȴ�����=�˾M�Ӿx{־5ҾM�ƾ�-��	!������)�F;p�#%r�G��?��/���Yg���ɾ��Ӿ�n־,AҾKɾI���P1���Ħ�/���������n� �V��B��l3���,�ds/��:�:�L��c��|�G�J����ɡ�5��<���djľf�ξ<Pվ@�վ�Ͼ>I�������~��e����kx��n��v�?톾�U��6a��Be��1�;�վ_�վ��Ͼ��ž���qU����Qʗ�m�����i�f��AO��Z<�"I0��,�_F2�@��&T��l���������TP�������氾�����ȾHsѾ�F־;{Ծl6˾�s��t⧾f������is���o���|�:��W枾�����ľgDѾKa־xJԾI�̾����e��φ���M��b���,��[.w��w^�vXH�6z7��.��-��6�+F�f�[��dt�����.���j���E��pʴ�����a�˾��Ӿ�}־�7Ҿ��ƾz0���#��Z!��D/��@p�*r�\I��>��碥��h���ɾ��Ӿ�o־�AҾ�Kɾ���?2���Ŧ����������[�n�گV��B��q3���,�nx/�ɧ:���L�S�c���|�
Ċ�膖�pˡ��������lľ7�ξJRվ��վ�ϾL��ܟ��D���Σ��qrx���n�ϓv�q����X���c���g��O�;�  �  �V����������ڹ��չ����8l��y𰾹���������M!z���`��AP�w]K� S���e��G��my���������v���4��I��<幾�Ĺ�\�������M���[إ��������uu�wS]��N�L�K��kU�7�i��������R���ƫ�K|��г��:u���깾o����a��e����L���أ��,������p��Z�p;M���L��#X��n��@������_v�� R��g�� ��>���깾��������X��Ь��������vh��g�l��/W��9L���M��%[�jr��ʇ����������Į��<��g�� ����蹾g�������&��#;��V���7)���遾Xmh�ǏT���K�
O�lo^�~�v�sX���j���{��������1θ��ɹ��๾u6��M����� ����S��͜��9�~�k{d��<R�%HK�i�P��a�H�{�茾�ț�1Y���T��=������pٹ��Թ������j��ﰾ	���� ������z���`�W<P�XK���R�S�e�+E��w�����'���u���3��(H���乾�ù�Ե���������uץ�����s~���qu��O]�	�N� �K�xgU���i�o���� ���P���ī�mz������s�� 鹾4����`��}����K��Tأ�*,������p��Z��;M�;�L�}$X��n��A��x���|w��gS���h���!�����칾����������~Ҭ�Lá����� k����l�5W��>L�Q�M�*[��mr�<̇�k���Ά���Ů�_=��4���ӵ���鹾#h������(��=�������+��.쁾�rh�L�T��K�hO��t^�G w��Z���l���}�����v����ϸ�6˹�y⹾ 8��/���������V������S�~���d�CR��NK���P�b�ܷ{��ꌾ˛�0[���  �  �m��p���G���V���Jƾh$оk�վMվiC;�o���D���F�����1�u�Wo�
ty������廯�48¾F�Ͼ+־�վ�8ξ,�þn���m��2,���㕾^���a{��|b���K���9�/��-��4�wC�!�W��7p�{���~����1��e��?ײ�������ɾH�Ҿ�z־!tӾ��Ⱦ]��q����������L�q�R�p�:�����FA���@��_eǾ��Ҿ��־�WӾ�˾�쿾�!��i���o��T��� ����r���Z��E��U5��b-��f.�2:8�tI���_���x�I���Z����퟾P)�����7�¾0;��Ծ"L־��о�ľ\��ʝ�N��
�{��Yo�t�ۃ��7(��z���t����˾I�Ծ�)־EѾZ�Ǿ� ��sA���夾宙����y݁��j���R�W?�B�1�s�,���0�!>=�~uP� �g�qy��Č�l�����	���3����Hƾ:#о�վ�Kվ�A;�m��aB��ND�����r�u�oo�ny����ꖛ�U����5¾C�Ͼy־sվg7ξH�þ���=m��+���╾k��a_{�zb���K��9�./��-��	4�/C���W��3p�z�������%0��uc���ղ�[�����ɾA�Ҿ�y־hsӾ%�Ⱦ]��-���u��������q���p��:��K��B���A��xfǾ��Ҿf�־2YӾ�˾��#������Iq�����2��� s���Z��E��Z5��g-�3k.�`>8�FxI���_���x�����m����=*�����N�¾P1;?�Ծ�M־��оFľ�ﱾm͝��P����{��_o��$t������*������v����˾��Ծb+־�Ѿ��Ǿ2���B��?社ٰ�����߁�i�j�n�R�8?�?�1�l�,�w�0��C=��zP���g��{���Ō��  �  �9���曾�:����ƾ �ݾ(���d���_����M�
Ͼd����ڝ�����K���Pr��[���U����Ծ��쾳Y��#�%.�����ؾ8����|������򡆾y�o�#�U��>�4,�C��4�۵�H��AX%� 6��K��c�Ԑ��ԏ��a������@�ξC�侜[���� �K� ��a���5�T ƾ�^���ٗ�dF��I�����'���t&þ�uݾHk��A �s"�"���I�3ѾH	��ߙ������Mr����f��M��<8�4�&�m��s��H����6b*��<���R�s�l�Z���8��� )�����5־~�������q�����S+���׾�=��к��ے�2̊�����l˱�^̾�徚����3�m' �`��i1��Xɾ���������y���]�F���1�2I"��*�q�Fm�'� ��/���C��[���u��7��W图�9��i�ƾ�ݾ���oc��_�F���)辛
Ͼ�����ם��������o���W���R����Ծ��wW��/~��,�����ھؾS���|��'������y�o�ϒU�k�>�r1,��?�1����F��1T%��6��K��c�8��ӏ�5`�������ξ!�侟Z��$� �� �%a��^5� ƾ�^��ڗ��F������~������<'þ{vݾ\l�`B �$#������J�Ѿ=���������t��j�f��M��A8��&�8����������e*�R�<���R��l�~ᄾF���
*��%���6־��뾖����r�F����-ﾛ�׾�@������Jޒ�Wϊ���⿛�α��̾��h���t4�( ����2�Zɾp����������y��]�"F��1��N"�g0��v��r�`� �� 0�$�C��[�c�u��  �  �c���o���U���ھ����������� �ZT�|�	����Ҿ3@������������򺾽`پ7�����h�=��\���	�kE��o�Ҿi���/����g�g�Z���=�GC'��I�J~
�������l��;h��L3���L��n��ۋ�������þQP�\��������N��"����a��Ǿ��������N���l��QľH����c��"���-����[�����Ǿ�����u�� .r��3P�/�5�P!����Ŵ�$�����}	�Ե�%�+�:�wW�L�z�9ޓ��0����ξ��h�P��������>�X���}ݾ/����_��b>���/��T���܆ξ���%�^X�������,��+��a�ݾ�ϼ�i���І� �e���F�,.��Z���Ȇ�]��]��;��ј�^�+�#�C�+b�kb���n��{T���ھ������������eS�^�	�+���Ҿ=���|������������]پ4��[��0�1��|�B�	�7D��j�Ҿ}���I����e�Q�Z�T�=��@'� G�{
�
��ۿ����Xd�6��3���L�i n�9ڋ������þO���=��9���N��"�����a�̣Ǿū�����N��'m���Qľ��k	�������8.�a��.�����Ǿ´���w���2r�)8P��5�!�P��h�����/����	�t��S%��:�W���z�Zߓ��1��*�ξF��2�=���ܽ�@�a����ݾ����Kc���A���2��T�����ξ3��#&�FY����������,����ݾѼ�pj��s҆���e�ʙF��.��_�?��	��������*��p����+��C��b��  �  ����	8���Zž/��M}�TO�H,�2�0�U+�$3��
���뾬Oɾ�����u��Q����о�}�����{� �.$-��u0�3*�[�����徍̼�i���|���P�*v0�=���s�a$������l����������%��.A�kVg��ƌ�9���өҾ�����2�br$���.�}�/�I'��3��>�	C߾�H���������Z���^J۾� �Y�%�%��R/�_/�z�%��Y��� �-4׾������9El�y�D�Q�'�4���7�i$��'��}���U��H�����>r-���L�ףv����������p�0�����b�(�70�7�-�}�"�O�����X�Ӿw˸��¬��p��>!ƾ�羭��8A���)��p0�9-��!�~���L󾃺ɾ=ꤾ�����]�":����NG��� �\F���e9�_����S��~�6��\Y�����6���Yž'���|��N�mG,�a�0�Z+��1��
����tLɾ|���Jr������nоZz����� ��"-��t0�A*����r���徍˼�r���|���P��s0�����p�����{ｏe������^��>%�V+A�Sg�EŌ�Ď���ҾV���2��q$�o�.�(�/��H'��3��>��B߾�H���������Ԝ���J۾g� �����%�qS/��_/�8�%��Z�x� �6׾����'����Il���D���'����m<�v-�������]�����/��0u-�N�L�O�v���������@r���x��^�(�@80���-���"����|���ִӾ�θ�>Ƭ� t��Z$ƾ������NB���)�hq0��9-�!����M󾭻ɾ�뤾����"�]�	&:����K��� �`P���;C����V��b��#�6��_Y��  �  ք���� %Ͼ���B���,�\�;���@��y:��*��K��d��r�־����Ӷ��3¾�޾����V�Z�.���<��t@��9��n(�
��VU�Siž2��e}�2!M�;3*�١�� ���콱���߽{��9&��U_	��(��'<���e�
�� ���QL޾	/����3�2���>���?�x(6��$�����n��̾���ې���ɾ����3�!��4�7?�Z1?��l4�c!���	��x㾹o��⠒�Atk�<'@��� ��H�{���2��Y�z�k����k�2�&�-�H���v� ��'�������K��%&�Ц7��+@�´=�e�0�6���[��k�ľ�)���^��AhӾ,�������(��%9��u@�;�<�E�.��������Ծ:L���"��]�[��4����h����Y併v߽+]�V~���KQ�T�0�g�V��Ԅ�T���#Ͼ��B�3�,���;���@��x:���*�cJ��a��#�־D��0ж�0¾I�޾:��<U���.�'�<��s@� 9��m(�Z��)T�Ehž0��Y}�M��0*�2��"� ��������߽5������[	�%��$<�Z�e��������K޾r.�b����2�/�>���?�5(6�t$����gn��̾7���1���{�ɾ� �p���!��4��7?�2?��m4��c!���	��z㾲q�������xk��+@�k� ��M�������#ཬ����Tn�''��H�Y�v�X!��e���7L�s&&�է7��,@��=���0��������	�ľH-��Kb��pkӾ���N��ӛ(��&9��v@�۸<���.�%��S��� ԾM��9$����[�Ð4�$��������Xc�s�߽�f㽀���>U���0���V��  �  �~�����g�Ҿ����6���1�;A��kF��@���/�9R����۾�¾�{��EGƾ���P��ڐ�64��jB�9EF��>��'-�K��ɡ��ʸȾ{�����}�0OL��f(�6`��,��)�e]ݽ�w۽23�t���W���:���e����~��T�� m
��8#�s�7��9D�A�E�H�;�4�(�_��1��^ѾJ^��>I���Gξ������4&�[�9�X�D���D���9�9�%��A�p�'��yӓ��k�k�>����5�������y��۽�ܽ�u�h?���"� %�r�G��w�џ����þ�����\�*�=���E�ggC�#6��$!��{	����Y�Ⱦ�Ժ�N;��'ؾ������>i-�]�>��FF��\B�*�3��������ؾGv���눾�,[�23�\���d�R����߽r۽��޽������ ��T/�]
V�J}�����Y�Ҿ��o6�c�1�^:A�"kF��@���/��P������۾�¾	x���Cƾ�㾊��.��� 4�KiB�DF��>��&-����������Ⱦv�����}��LL��d(��]��&���"轰Vݽ�p۽�+��l�-���!�:�x�e�����}���⾊l
�K8#���7�d9D��E��;��(��^��1��^Ѿ{^���I��6HξB��[���4&���9���D�W�D�S�9��%�zB�J�)���Փ�5�k���>�c������������}�۽8�ܽ[}�~F���%�#%�)�G�u�w�����þ���>�*�=���E��hC��	6�^&!��}	�A����Ⱦtغ��>��\"ؾ�������Xj-�H�>�^GF�4]B���3���A��ؾ�w��G툾	0[��3����Vi�����߽)۽7�޽���)��p$�1X/�vV��  �  ք���� %Ͼ���B���,�\�;���@��y:��*��K��d��r�־����Ӷ��3¾�޾����V�Z�.���<��t@��9��n(�
��VU�Siž2��e}�2!M�;3*�١�� ���콱���߽{��9&��U_	��(��'<���e�
�� ���QL޾	/����3�2���>���?�x(6��$�����n��̾���ې���ɾ����3�!��4�7?�Z1?��l4�c!���	��x㾹o��⠒�Atk�<'@��� ��H�{���2��Y�z�k����k�2�&�-�H���v� ��'�������K��%&�Ц7��+@�´=�e�0�6���[��k�ľ�)���^��AhӾ,�������(��%9��u@�;�<�E�.��������Ծ:L���"��]�[��4����h����Y併v߽+]�V~���KQ�T�0�g�V��Ԅ�T���#Ͼ��B�3�,���;���@��x:���*�cJ��a��#�־D��0ж�0¾I�޾:��<U���.�'�<��s@� 9��m(�Z��)T�Ehž0��Y}�M��0*�2��"� ��������߽5������[	�%��$<�Z�e��������K޾r.�b����2�/�>���?�5(6�t$����gn��̾7���1���{�ɾ� �p���!��4��7?�2?��m4��c!���	��z㾲q�������xk��+@�k� ��M�������#ཬ����Tn�''��H�Y�v�X!��e���7L�s&&�է7��,@��=���0��������	�ľH-��Kb��pkӾ���N��ӛ(��&9��v@�۸<���.�%��S��� ԾM��9$����[�Ð4�$��������Xc�s�߽�f㽀���>U���0���V��  �  ����	8���Zž/��M}�TO�H,�2�0�U+�$3��
���뾬Oɾ�����u��Q����о�}�����{� �.$-��u0�3*�[�����徍̼�i���|���P�*v0�=���s�a$������l����������%��.A�kVg��ƌ�9���өҾ�����2�br$���.�}�/�I'��3��>�	C߾�H���������Z���^J۾� �Y�%�%��R/�_/�z�%��Y��� �-4׾������9El�y�D�Q�'�4���7�i$��'��}���U��H�����>r-���L�ףv����������p�0�����b�(�70�7�-�}�"�O�����X�Ӿw˸��¬��p��>!ƾ�羭��8A���)��p0�9-��!�~���L󾃺ɾ=ꤾ�����]�":����NG��� �\F���e9�_����S��~�6��\Y�����6���Yž'���|��N�mG,�a�0�Z+��1��
����tLɾ|���Jr������nоZz����� ��"-��t0�A*����r���徍˼�r���|���P��s0�����p�����{ｏe������^��>%�V+A�Sg�EŌ�Ď���ҾV���2��q$�o�.�(�/��H'��3��>��B߾�H���������Ԝ���J۾g� �����%�qS/��_/�8�%��Z�x� �6׾����'����Il���D���'����m<�v-�������]�����/��0u-�N�L�O�v���������@r���x��^�(�@80���-���"����|���ִӾ�θ�>Ƭ� t��Z$ƾ������NB���)�hq0��9-�!����M󾭻ɾ�뤾����"�]�	&:����K��� �`P���;C����V��b��#�6��_Y��  �  �c���o���U���ھ����������� �ZT�|�	����Ҿ3@������������򺾽`پ7�����h�=��\���	�kE��o�Ҿi���/����g�g�Z���=�GC'��I�J~
�������l��;h��L3���L��n��ۋ�������þQP�\��������N��"����a��Ǿ��������N���l��QľH����c��"���-����[�����Ǿ�����u�� .r��3P�/�5�P!����Ŵ�$�����}	�Ե�%�+�:�wW�L�z�9ޓ��0����ξ��h�P��������>�X���}ݾ/����_��b>���/��T���܆ξ���%�^X�������,��+��a�ݾ�ϼ�i���І� �e���F�,.��Z���Ȇ�]��]��;��ј�^�+�#�C�+b�kb���n��{T���ھ������������eS�^�	�+���Ҿ=���|������������]پ4��[��0�1��|�B�	�7D��j�Ҿ}���I����e�Q�Z�T�=��@'� G�{
�
��ۿ����Xd�6��3���L�i n�9ڋ������þO���=��9���N��"�����a�̣Ǿū�����N��'m���Qľ��k	�������8.�a��.�����Ǿ´���w���2r�)8P��5�!�P��h�����/����	�t��S%��:�W���z�Zߓ��1��*�ξF��2�=���ܽ�@�a����ݾ����Kc���A���2��T�����ξ3��#&�FY����������,����ݾѼ�pj��s҆���e�ʙF��.��_�?��	��������*��p����+��C��b��  �  �9���曾�:����ƾ �ݾ(���d���_����M�
Ͼd����ڝ�����K���Pr��[���U����Ծ��쾳Y��#�%.�����ؾ8����|������򡆾y�o�#�U��>�4,�C��4�۵�H��AX%� 6��K��c�Ԑ��ԏ��a������@�ξC�侜[���� �K� ��a���5�T ƾ�^���ٗ�dF��I�����'���t&þ�uݾHk��A �s"�"���I�3ѾH	��ߙ������Mr����f��M��<8�4�&�m��s��H����6b*��<���R�s�l�Z���8��� )�����5־~�������q�����S+���׾�=��к��ے�2̊�����l˱�^̾�徚����3�m' �`��i1��Xɾ���������y���]�F���1�2I"��*�q�Fm�'� ��/���C��[���u��7��W图�9��i�ƾ�ݾ���oc��_�F���)辛
Ͼ�����ם��������o���W���R����Ծ��wW��/~��,�����ھؾS���|��'������y�o�ϒU�k�>�r1,��?�1����F��1T%��6��K��c�8��ӏ�5`�������ξ!�侟Z��$� �� �%a��^5� ƾ�^��ڗ��F������~������<'þ{vݾ\l�`B �$#������J�Ѿ=���������t��j�f��M��A8��&�8����������e*�R�<���R��l�~ᄾF���
*��%���6־��뾖����r�F����-ﾛ�׾�@������Jޒ�Wϊ���⿛�α��̾��h���t4�( ����2�Zɾp����������y��]�"F��1��N"�g0��v��r�`� �� 0�$�C��[�c�u��  �  �m��p���G���V���Jƾh$оk�վMվiC;�o���D���F�����1�u�Wo�
ty������廯�48¾F�Ͼ+־�վ�8ξ,�þn���m��2,���㕾^���a{��|b���K���9�/��-��4�wC�!�W��7p�{���~����1��e��?ײ�������ɾH�Ҿ�z־!tӾ��Ⱦ]��q����������L�q�R�p�:�����FA���@��_eǾ��Ҿ��־�WӾ�˾�쿾�!��i���o��T��� ����r���Z��E��U5��b-��f.�2:8�tI���_���x�I���Z����퟾P)�����7�¾0;��Ծ"L־��о�ľ\��ʝ�N��
�{��Yo�t�ۃ��7(��z���t����˾I�Ծ�)־EѾZ�Ǿ� ��sA���夾宙����y݁��j���R�W?�B�1�s�,���0�!>=�~uP� �g�qy��Č�l�����	���3����Hƾ:#о�վ�Kվ�A;�m��aB��ND�����r�u�oo�ny����ꖛ�U����5¾C�Ͼy־sվg7ξH�þ���=m��+���╾k��a_{�zb���K��9�./��-��	4�/C���W��3p�z�������%0��uc���ղ�[�����ɾA�Ҿ�y־hsӾ%�Ⱦ]��-���u��������q���p��:��K��B���A��xfǾ��Ҿf�־2YӾ�˾��#������Iq�����2��� s���Z��E��Z5��g-�3k.�`>8�FxI���_���x�����m����=*�����N�¾P1;?�Ծ�M־��оFľ�ﱾm͝��P����{��_o��$t������*������v����˾��Ծb+־�Ѿ��Ǿ2���B��?社ٰ�����߁�i�j�n�R�8?�?�1�l�,�w�0��C=��zP���g��{���Ō��  �  �V����������ڹ��չ����8l��y𰾹���������M!z���`��AP�w]K� S���e��G��my���������v���4��I��<幾�Ĺ�\�������M���[إ��������uu�wS]��N�L�K��kU�7�i��������R���ƫ�K|��г��:u���깾o����a��e����L���أ��,������p��Z�p;M���L��#X��n��@������_v�� R��g�� ��>���깾��������X��Ь��������vh��g�l��/W��9L���M��%[�jr��ʇ����������Į��<��g�� ����蹾g�������&��#;��V���7)���遾Xmh�ǏT���K�
O�lo^�~�v�sX���j���{��������1θ��ɹ��๾u6��M����� ����S��͜��9�~�k{d��<R�%HK�i�P��a�H�{�茾�ț�1Y���T��=������pٹ��Թ������j��ﰾ	���� ������z���`�W<P�XK���R�S�e�+E��w�����'���u���3��(H���乾�ù�Ե���������uץ�����s~���qu��O]�	�N� �K�xgU���i�o���� ���P���ī�mz������s�� 鹾4����`��}����K��Tأ�*,������p��Z��;M�;�L�}$X��n��A��x���|w��gS���h���!�����칾����������~Ҭ�Lá����� k����l�5W��>L�Q�M�*[��mr�<̇�k���Ά���Ů�_=��4���ӵ���鹾#h������(��=�������+��.쁾�rh�L�T��K�hO��t^�G w��Z���l���}�����v����ϸ�6˹�y⹾ 8��/���������V������S�~���d�CR��NK���P�b�ܷ{��ꌾ˛�0[���  �  ؆վ�վ�Ͼɫž 	���V��I	���˗�	��9��u�f�TFO�^_<�N0��,�^K2��@�+T��l�b���Î��Q��}����簾���cȾ�sѾ.G־�{ԾC7˾�t���㧾 ���ns�E�o���|��<���螾���:�ľ�FѾDc־GLԾ�̾A������퇪��N��)������@/w�qx^��XH�*z7�Q.�b�-��6��)F���[��bt�Ұ��⫒����WD���ȴ�����=�˾M�Ӿx{־5ҾM�ƾ�-��	!������)�F;p�#%r�G��?��/���Yg���ɾ��Ӿ�n־,AҾKɾI���P1���Ħ�/���������n� �V��B��l3���,�ds/��:�:�L��c��|�G�J����ɡ�5��<���djľf�ξ<Pվ@�վ�Ͼ>I�������~��e����kx��n��v�?톾�U��6a��Be��1�;�վ_�վ��Ͼ��ž���qU����Qʗ�m�����i�f��AO��Z<�"I0��,�_F2�@��&T��l���������TP�������氾�����ȾHsѾ�F־;{Ծl6˾�s��t⧾f������is���o���|�:��W枾�����ľgDѾKa־xJԾI�̾����e��φ���M��b���,��[.w��w^�vXH�6z7��.��-��6�+F�f�[��dt�����.���j���E��pʴ�����a�˾��Ӿ�}־�7Ҿ��ƾz0���#��Z!��D/��@p�*r�\I��>��碥��h���ɾ��Ӿ�o־�AҾ�Kɾ���?2���Ŧ����������[�n�گV��B��q3���,�nx/�ɧ:���L�S�c���|�
Ċ�膖�pˡ��������lľ7�ξJRվ��վ�ϾL��ܟ��D���Σ��qrx���n�ϓv�q����X���c���g��O�;�  �  �n���������ܾ�{ž����ٚ��P��m?t���Y���B�A/�h4 �v�|~�����
#���2��\G��J_�R�z���������ܳ�U�ʾdh� ����\ �������7侟�ʾ�l�������z��U��������������,>پIG����e��3�������Ծ�ѽ������������j���Q���;��)��z�}{����b���'��U9���N�	�g�K��R���Y���9J��^Ҿ�k�h����<�� �od�ܾP���7v���7���`������{ǘ�����՜Ǿ[��FQ���� �� �_�����9;�P���G��$�����}��$b���I�s5���$�n����Px�3��9-�r!@��V��q�����ZĘ�,���[�¾� ھ�����&}�����˶�+tӾ�߸��.���Đ�3�������I)��k�о�K�
J���m�Z������Ȁܾ�zž`��Gؚ�wO��Y<t�4�Y��}B�/� 0 ����y���7#���2��XG�kG_���z�����4��vܳ���ʾ(h�ƿ��b\ �O�����6�2�ʾ�j������Xx�������S��������;پ�D�I���d�2��֧�?�Ծfн�����������j���Q��;�ҁ)��z��{�7��c�?�'�oW9���N�Th��L��м�����L��`Ҿ&n�ƾ���=�'
 �6g��ܾ6���y���:��Bc��B����ɘ�������Ǿɐ�eR��d� �8� ������㾶9;�Q���H��bᎾ��}�}(b���I��5�=�$��r�ƞ�}�����"-��%@���V�q�T����Ř�������¾�ھv������g~�a����뾀wӾM㸾,2��uȐ�ދ�������S��N�оTN�GL���  �  ���h����n����%ؾ��������N2���3`�B�<�*�}����u��ȗ�^���w�SF�!P/�J&H���g���8�ڒ��=�߾�y �5��`��.��n���R�)�̾O��ʛ�� t���V�����t�޾�Z �����/��"���E�a����̾����~���x��SU�#�9��$����	�T`����"��{��"�A�6�h�Q��Pt� ʏ��L���Tɾ��H���x�&^�����D�K%�����¾�Y����������׮�hTɾJF꾄����@|��v���Q:��n��¾���<���l�k�XMK���1�����ҋ��� *���
�(�5Y(��%?�Ex\��؀�V��3���gԾ~���j
�~������S��X��
�׾gv��f���+霾�2��x�����Ӿ���F�
�������g����*����$ؾ����S����0���0`��B���*������+��s�����s��B��L/�g#H�B�g�7���젾~����߾�y �)��E�������eR�����̾M��t���}q��CT��e�����޾oY ��������$���D�ɰ�\�̾L����}��J�x��RU�/�9�\$����	��`���#��|�~"�<�6���Q��St��ˏ�;N��iVɾ3��i���y�s_����cF��&�����¾�\��j�������ڮ��VɾH�;������|��v�0��:� o㾐¾����T���!�k��PK�:�1�� �j��K��s���.���Z�,](��)?��{\��ڀ�����4��9iԾY���k
������b����F\��Ɖ׾Bz��Nä�
휾�6�������Ӿ �����
�����  �  �0���+��b��W�0��0þVf���=��,W�[-5�8b�l�
������� ����z.�c*�M5!���;��1`��#���̦���˾Q��������!���-�U0�GP)��C�����i�z�ľ��������I�վ�-�����q#�L].�x0�$(��~��V��޾����씾��s�>�J���+�����B�L���!~�f��a���������l")���F�S�n�����
����~پ%���h�E�&��/��/�j
%�I�����1WپrU��ß��������CH��a�:<�<�'�"0��m.�p�#����p��iо/���t5���d�_?��#�q��FW�����D�)��C���3	�n�Z�1�:�R�[�~��ћ�达�v羐	��{���*�T�0���,�*��q�E�Uξ)����]���Գ��ʾ���1�$�Z�+�ە0��+�9b�W��.쾞/þ#e���<��4)W�.*5��^���
�������a����*��&�02!��;��/`�#��v̦�r�˾D��������!���-��T0��O)�WC�˨��g�P�ľ����g�������վ�*������o#�\.�Y0��"(�	~�V�,޾͏��{딾��s��J���+�@��aB�X����~��_�����d��l$)�O�F��n����ā����پ4��j���&�a�/�	/��%�������HZپ{X����������\���lJ��b��<���'��0�0n.���#���#q���iо꟪�n6����d�b?�~�#�>��Z[�4��jM���ｻ���7	�P�2���R���~�Cӛ��龾gx羈	��|��*���0�,�,�����r�fI�Yξ;����a���س�9�ʾ��G3�w%���+��  �  ��@��;�O�+�,���d��y�̾|��M8���%T��;/���?F������Y�߽�佃�󽝣�C ��h6��^�Rԉ��n��(�־|��#���/�77=�TW@��q8��}'��y�XL���Ѿ�����o����ž��bP�b�0�1�#>��?�|�6�t�$����VZ��S��7���	t�PxF�ys%�e[����>=�>�ཝR���b���J��o"��8B��Dn�w��l���B�b?��"�!E5��|?���>���3�:z ���	���!Ⱦ����5��
sξ������4%���6���?�\>�^�1�������X�۾@İ��F��>Mc��2:����m�����潜�߽��v�������A�+��jO����� ���Ǿ����M��)���9�?�@��:<��-�R�vU��ܾ���_���=��E�ؾn���Ď��+��;��@��;���+�����c��T�̾L��7���"T�m8/�\��B���!��o�߽Y��,��A��O��f6��^��Ӊ��n���־���#���/�/7=�*W@��q8��|'��x�xJ��ҵѾ~���*m����ž2���N����1��!>���?�p�6���$����X뾉R��r6�� t��vF�|r%��Z�p���H=�����S���	����K��q"��:B��Gn��x��*���3�s@�,�"�dF5��}?�!�>�4�3��{ �3�	�C��8�Ⱦ�"���8���uξ)�����5%��6���?��>���1������ʻ۾�İ��G���Oc�t5:�N���q�`�����߽]"�����������+�nO�j�������Ǿ_���N�:�)���9���@�i<<���-�9�wW�$�ܾ�������B���ؾ����a����+��;��  �  ����:y���h��*�g�Lw=����龖� g��R�g�ϦA��@(�K;����;�q����+�,�Y�H�JUr��얾y<��~R���]�L�F���p��%���z���`�����ȉ��ԕ_�7�8�J6�����`)�ZK)��M��v�m����S���������M���Y�5�/�s<
�\�־)���M ��n^Y��7�[�!�-��]���#�� ��5���T����F����о�t�RV+�G�T�}P~�C%�������������
fz�fR���,�#j���&d�r�;�4�[�(x��c�����kN��u挿#{u�<{K���"��W��ۤž�䚾��w�ͺL���/����/���S�t��x���
&��B>�ۺb�V׋�����U��
���8�nc��n��OL��̐��b���Nf��Fm���D�)l"�4*��w�q	�N3�{�@��h�������������x��)h����g��v=�w����T쵾�e��7�g�g�A�%=(�j7����7�������,�e�H��Rr��떾�;��8R���]�j�F���p��%���z���`����������_�=�8�5����G��'��I)�l�M�Hv�����4S���
������YM��	�Y�o�/��;
�A�־B������d]Y�U�7��!�1�������)��u �w5���T����:H��q�о�u�VW+�f�T��Q~��%��W���F��|����gz�R�[�,��k�����e�cs�^�4�[��x������B��{N��{挿){u�L{K��"�oX����ž暾��w��L�l�/����_��#X�������&��F>���b�ً����XW�����8�wc�Co���L������?���Bg��S!m���D�an"�q,��y�2s	�V5�^�@�Ġh�ۂ��`����  �  �v������V'���a��8���s��Hٴ�6���)�i���D���+�u�O��8F��
��[��D0�f�K��Lt�����¾�������A���i���u��8��+>��l�~��Y�m�3������pM �@���%�{�G���n��n��D��"甿t䌿�z�5�S���+������Ծn(��s�8�[�%$;��F%����+������e#��98�n�W�����W䢾��ξj"��g'�O�S�v��y���w��C}����r��0L�#�(���� ��������/�g�T���z�팿s锿5?���b�� *n�[F����Q����þ�Κ���y�k�O�F�2�������_���U ��V)�L]A��e�#C��O ��q྾8��R4���\�gE��n���e��ϔ��Y���f�V�?�s�h�dv��1p��Z�܌;���a�%9��Ӓ��Sv��>����&��Ra�[�8�^�I��ش�ͳ���i�O�D� �+�1q�C��'B����W�3A0�b�K�iJt�	���s���3����2�A���i�����u��8��>����~�%Y�t�3�V��9��L ����@%���G�-�n�n��fC���政�㌿�z�T�S���+����Ծ�'������/�[�x#;��F%� ��b+�~����{f#�~;8���W����墾��ξS#��h'�0O���v�mz��mx��F��&�r�=2L�ʈ(�S��� �������/�T�T�P�z�S팿�锿G?���b��	*n�oF����R����þК���y�ĚO��2����9��gc�<��$��Z)�2aA��e��D��"���rྛ9��S4���\��E���n���f������J���f�x�?�:u����z��Qr��\���;�S�a��9��w����  �  _��'��3o���N��,��>���޾uﲾ%����1r���N�#6�r�%�O���������(���:�c�U���{�3��M���`F�1)�T�3���V��Xu�̄��&��7���Kh��.G��#&��x��������1�|8�G	Z��x�Lr��]冿K ��W'e�T[C�� ��Z�P�ξ��������Ve���E�6�/�/�!����Y��� ���-�B�B��`�P���颾��ɾa��Z���q?���a��}�ʅ�����D�z���]�Q�;��G����n���j	���"�D`C���d����ᆿay��r:x��VZ��7���+��T��¦���j���RY��Q=�}:*������Ʈ�n1$�j�3���K�P�m�#��e����tپ���1(��"K���k� 0��FQ�������r�W�R�_�0��U������������-���N���n�����^���&��]2o�B�N�,�7>�\�޾+����R.r�L�N�P6�f�%��J�������ŕ(���:�1�U���{�2�������E�")�a�3�͚V��Xu�̄��&����Kh�.G� #&��w��������{0�	8��Z�;x��q���䆿���_&e�xZC�S� ��Y�;�ξ��������Qe�ގE��/�4�!�q��oZ��� ���-���B�� a�����iꢾ-�ɾ�b��Z���r?�+�a�^�}�|���U����z�M�]���;�'I�t��{�h���	��"�.aC�F�d����&↿wy���:x��VZ��7�P���+��U������+l��nVY�vU=��>*�I����5���5$���3���K�
�m�倎����Tvپ����2(��#K���k��0��R��a����r�O�R�q�0�X� �����7������� -�,�N���n�{���  �  �g���a�k�O��6��c�Ѯ�5Z׾-ѳ�L헾�A���c���I���7�Qz-���*��(/�7L;��N���i�e���ԉ����Zf྇�xm!�g�<�sqT��d��lg��|]��H�[�-�����`����޾��پ�&���
`!� 
=�tMU���d�2g��\���G�B�-������%�ʾ�������^x��Y�cC�H�3���+��9+��\2�	�@�=�V�7�t�����������ƾ�����6�*��&E���Z�M�f���e�W�W�z@�<m$�'�
��W���ھ?Fݾw�������*���E�ݡ[���f�$e��V��?��w$���	���6���ru���ވ�[?m��fQ��=�0�'�*���,�h6��wG���_�2+��3;��\����Ҿ����e���3�c*M��	`���g�3b�H�P�X�6�PY�T/� z�cپ��� ��f�Y�3���M�X�`��g��a���O�{�6�0c�@��Y׾�ϳ��뗾R@���c���I���7��u-�6�*�)$/��G;��N�L�i�Ꙇ�����C���e�d�qm!�o�<�{qT��d��lg��|]���H���-����^��T�޾��پ�#�h��^!��=�'LU�O�d��0g��\���G�m�-�������ʾ����_���]x�_�Y�C�O�3��+��:+��]2�c�@���V�B�t�ě�����L�ƾ~����K�*��'E���Z���f���e�׈W�@��n$���
��Z���ھIݾ�y�������*�A�E�_�[�N�f�\e��V��?��w$���	���K����v������ Cm��jQ��=��#0�ӭ*�\�,��l6�#|G���_�-���<���]��k�Ҿ0���f�u�3�w+M��
`�f�g��4b��P�8�6�J[�_1�?~�x!پ�� � ��h���3�%�M���`��  �  }�>���:�2/�Uj��������s_־k~���u��\��|Ƃ�w�i�,{T��hG���C���I�?�X��eo��>��b��7������`�ܾg�����f"�~\2���<��>���5���%� f�`B��uA׾��¾�Ͼ��3̾4�������/���;�]>���7�1�)�)M�n���7꾓@;_Ŵ�̟�>���ߠ{���a�{"O��E�щD��M��\_��tx�Ŭ�����H��FRʾM�澙��~=��%(��6�>� b<��c1��c�kH
���G�ξhs���d��M7Ծ��� ���#�I�4��=��$=���3�5Z$���& ��ྀ�ľ2p��#o������Tr�+�Z�W�J��C��F���R�?�f����+c���2��r޹�EӾP��	�vc�k�-�-�9�S�>���9�n�+��{�FO�@Sᾃ�Ǿ�%����ž��ݾ�
�"��*���8���>��:�k1/��i�i������:^־}��Lt��ZZ���Ă�6�i��vT��cG��C���I���X�9ao��<��p`�����v�����ܾ�f��y�wf"�q\2�ۂ<��>�_�5��%�Ge��@��]?׾[�¾L;��0̾������z�ɬ/�~�;��[>���7�L�)�\L����P6꾐?;�Ĵ�]˟�Ì��?�{���a��"O�E���D��M�:^_�Pvx�ȭ��0���cI���Sʾ	�澏���>��&(�S�6�j>�cc<�2e1�e��I
���=�ξ>v��-g���9Ծ9������#�ю4�q�=�%=���3�lZ$�# �� �����ľ�q���p����LYr��Z�E�J��C���F�F�R��g���e���4��๾�FӾ�Q�v�	�[d�m�-�S�9���>��9�,��}�"Q�W�f�Ǿ�)��[�ž-�ݾf��#�S*���8��  �  ���;�_������� �:p�*ҾC��P`���.��
7����|��*k�f�Mn�z���ȏ�|/��{k��0ž]�վ��S�����'���z����%��z�������(!ξ{���ԥ�Z󢾺⬾�¾�޾��������d������t���������r�ݾ��̾3e���G��K���(����u��g�`;g�P�s�Đ���_���>���i��z�ʾ47۾~�����������*f���_��)��� �c3⾂�ľ'���cl���ݤ��в�p�ʾ�*����(���L�����*������������羐�׾�Ǿ"l���1��i���������o��;f���i�Hz��z���1��W���P��zSо�ྌ6�jz�C�
��*������Ⱦ�X
����s�׾`��ƛ��[t���1���湾�ԾP��Q�����$���:������������n⾞(Ҿ�A��w^���,���4���|��%k���e�n����hƏ�N-���i���ž�վ�澥���؎�����z�[�������c����oξ}���ҥ���AାE¾��޾w���o���c������s�=��j����q�ݾء̾�d��1G��2K���(����u�h�g�<g�Q�s�o���^`���?���j����ʾ�8۾0�뾿��������[g�@����*�� �H6�e�ľ����o��JाӲ�{�ʾL,龬�����CM����=+�Ԯ�o��n������׾EǾ*n���3������ �����o��@f���i�Mz�}��4��Y��VR��Uо���8�,{��
��+�����%���
������׾􂼾e����w��_5��깾��Ծ!�󾑘�����  �  ����i ����t3��1�C��vG ����Ț�/�ؾ5¾
������u���ֈ��~���~��͇���SǾ�=ݾ<�z,��X� �8���6��+��������3��0���
վ�\��6��9-���7��W$��xK���}���;���"˾��ي񾀙������R8��"�v|�O���>8��g���`Ѿ%���wӤ�^ʓ��8��س��0Q��G�������]�ξ������J����V���7�a��A�jt����l��'�;l���y��������z��������量qͻ�
�Ҿp��������H��$&��7�7��� �4#������v߾��ɾ����w��ۨ��z ��)������r[��Ǣ��"=־I��������������-�F5�0��� �`����@�ܾ�	ƾ�L��ʄ��&Ȉ��ꌾ٦���㬾�zþ��پ��X���Ai �S���2�b1�����F �j����9�ؾ�2¾��������s���ӈ��{���{��'���@QǾ`;ݾ]��*���� ����6��+�k������53��S���	վ}[��n4��S+���5��"��&I���{���9��? ˾��ƈ񾑗�����
��7�/"��{�`���y7�����z`Ѿۇ��VӤ�fʓ�9��/����Q��𤢾U���X�ξ���6������]W���8�t��B��v��+����;/���9���:����}�����������'ϻ�y�Ҿ��������������&�J8���u� ��$�����9y߾�ɾf����y������V��񚋾n���]�����!?־�龐���L���I��P.�6���� �����C��ܾ�ƾ�O�����u�}ˈ��팾򩙾�款N}þO�پ���  �  �Ӿ7X������(<�D^��d��^��S���v��$�ҾJ�������^���qb���ٽ�8�پ����@�
�L0����������7
��� �/E�C�߾^iϾ$X���T���7������y��di��of�9�p��F��D����5���m����Ǿ��ؾC�辦���:�\(��~���u�+�0 �~l羓nɾL����s������鲯��eƾ����{�����m����b��"��������Oھ�ɾ8j��
:��k��kȄ�͇r���f�eh�=�v�v����B��TK��#a���;0�ݾlb���#2	�����1�����*,�W?���	ݾ���m��Q¢��[���8����Ͼ�g�PN��J�E������B9��
�&���'�3�ԾD%ľg���+��"ގ�5e���Dm�#�e�Q�k��~�K��[+���a��9¾6Ӿ�V㾏��I��;��]�Od�^�S������Ҿr�������D���R_���ֽ�J�پ4����
�;/����0��j���7
�x� ��D𾙹߾�hϾ5W���S���6�����}y��`i�tkf�ڡp�sD������3���k����Ǿ��ؾ��� ������'�~�+������8l�tnɾT����s��N���h����fƾ���r|�g��`n�����D��#�����@��VRھ��ɾ�l���<���m��˄��r���f��ih���v�c���nD���L��^b����;�ݾQc�{����2	�����2�����l-�B���ݾ������dŢ��^���;��K�Ͼ4j�UO�cK� �������9�A�����)�2�Ծ�'ľ�i��b.��ᎾCh���Jm�V�e�\�k��~�����-���c���:¾�  �  Gҽ���׾�������k�0�m\;�cr>�g�7��)�������}ܾ�žt>��{�Ⱦ�'㾎v������,�f6:�{�>�\w9�ǧ,��_�}��Q�ﾅ�Ѿ���3��l��B��k�e�W�Q�F���C�/nK�0�[��s�}툾�z��i����
ƾ����S'��P%�
�4��j=��W=���3���"����Q��?�Ҿ[����ܿ�� о���4w�l� ��72���<�"�=�k�5�l6'��5�?��&微�ȾU��В��龊���v��(^�}�L� ND��aE�z�O�gc��;}����]⠾R��2�ξ��뾬���S���*�J^8�Kv>�?*;�G�.����F����/˾�����fþ>�ؾ#m�������&�x�6�l2>�'<���1�hi!��
�.���P ۾����;穾�[��A[����m��yW���H���C�K�G��pU��k�3����X��+����н�`�׾������k��0��[;��q>�y�7��)����I���pܾ{ ž;���ȾZ$��t�<��w�,�45:�w�>��v9��,�_�
����ﾹ�Ѿ$���3���j���@��L�e�ݭQ�DF���C�jK���[���s�t눾�x������<	ƾz��6��&�'P%���4�fj=�PW=���3�x�"����4��H�Ҿ����ݿ� оE�w�� �+82�T�<���=�4�5�I7'��6�A �L���Ⱦ���D���k�����v��-^�l�L��RD�FfE���O�*c�#?}������㠾s��<�ξ���8��;T�E�*�/_8�Zw>�y+;���.�&�����S�澇˾֑��jþ5�ؾ�o��.����&�]�6�,3>��'<���1��i!�#������!۾���L驾�]���]��H�m�{W���H�\�C���G�8vU��k�~����Z�������  �  (�����پ��v��+8��P��3b���g��`��L��[2���� ���K��<پ1��_]����i�8� �Q�s�b�7�g� @_�O�K��)2�t���s����о�����듾�O~��X^��WF�R�5��u,���*���0��	>���R��
o����]������[v�"Q�O�%�j�@�e�W���e��f���Z�6_D��)�ވ�_��S�ܾ�O۾z
������%�zA�i�X���e��Nf�p�Y��C�	)��(��K�W�ľ����Hd��¬r��~U���?���1�+�m�+�UG4�FD��K[��Pz��V���[��֣̾SL�����,!/��=I�ڏ]��gg��d��#T�.�;�������Z��v�پ3�߾dg��0�ZA/�1�I�{\^��g��uc��IS�� ;�������޾"+��m��}��=h���M��h:�ڮ.�|{*���-���8�K�ʴd�vP��@K��������پ
�����*8�u�P�F3b���g��`�ĤL�/Z2�t��Ģ����ᾍ8پ��澕[�-���8���Q�$�b��g�0?_���K�A)2����	s����о�����꓾�M~�V^��TF���5�:r,���*��0��>�ĽR�o������l����t�pP���%���@��W�7�e���f�r�Z�_D�y)�ш�j�󾃎ܾ�O۾�
�@��#�%��zA���X�l�e��Of�5�Y���C��	)��)��M쾌�ľ� ���f����r�w�U���?��1��+���+�bK4��!D��N[��Sz��W���\����̾vM������!/�b>I�Ր]��hg�4d�"%T�͉;����i�����پ��߾�j�����B/�C�I�`]^���g�"vc�dJS�!;���� ��K޾�,��S��3���h���M��m:�E�.��*��-��8��	K��d�dR���L���  �  ��G��t����-���P��p�^���T[�����hNm�8�L��Z+��C������%�]B ����A�2��sT���s��b��A��򬁿Jj�13I��L&��9�U�־������Mrk�3J���2�b�#�1l�S��]��+��>�z2[�����l��e�¾>+�:���9��.\���y�Kƅ�D�����~��c��zA��!�5���&�����]������=��_��|��G���L��VH|���_��}=�) �PE���|Ǿ(���`���_��MA���,�7 �	1����ZK"�Ҵ0��G��$g����i���؊Ѿ�����"�^NE���f�0���@
�����-�v��-X��66���������" �������'�I�l�i�p����>���k����s�y�T�S�1�Ph��`�z�����WNy���S���9�E�'�\�����8I&��27��P��t��8���������.�-�!�P�y�p�
����Z������8Mm���L�#Y+�B����2"�v@ ����n�2��qT�)�s��a���@��q���2Ij��2I�/L&�9�Z�־��������ok�}J���2��#��h�������+��>��.[�O���k��˭¾�)��s�9�R.\�/�y�ƅ����I�~�vc��zA��!�:���&��ߦ���C��t�=���_�"|��G���L��I|���_��~=�!�]G��Ǿh��@c���_�ORA���,�� ��5����SO"�y�0��
G��'g�H������
�Ѿ ����"�OE���f������
��7����v��/X��86���������#��B��"�'�_I���i�✁�X?��	l��6�s��T���1��h��a羊{��̃��\Ry���S�Õ9�J�'�-a�+��(��N&�e77��P���t�C:���  �  &D�����j�B�:��Dc����t��	s�����L��-�_��9����)��֞������ �ޯA�u5h��腿&���R���Վ�gO���\Z��$2��S�hݾ�ԭ�p���y�b�_�?�tK(�������#x��H��� ��4�,�Q��|�ǜ�
�ƾپ���"!��YH��Kp�r0������N���|;��b�x�֟R���-����p��6��A�rQ*�:TN���t��Ɗ��8��5��I����t�*�L��L%��[��̾�Р��/��ْU��6�g|"��2����"\��P��?&�:�<��-^��V���W��s׾˖	��-��U�B�|����U���Ⓙ�����ul�{�E��X#���
�� ��I����H�5��C[�Wf���܎�ZS������م�;�g��a?����J�07������q���I�/����ߥ�.:�G���!�Ī,�iF��wl�?x���B���������:�`Dc�������r������K��ė_�z�9���M���������� ���A��3h�$腿k��R��CՎ��N���[Z��#2�$S��fݾ�ӭ�S����b���?�xH(����1���t��D�+� �/4���Q�z�|��Ŝ�x�ƾe���*"!�YH�pKp�70��y���$���Z;��1�x���R���-������7��A��Q*��TN��t��Ɗ�9��q5������Ղt��L��M%��\��̾�Ҡ�22����U���6��"�W7�(��U`��T�[C&���<��0^�X���X��[t׾m�	���-���U�-�|���������㒿u���^wl�X�E��Z#���
�� �TK�0��ƙ5�<E[��f��Yݎ��S��#���م���g�-b?����2L�8��>��Ȥq���I��/����ڪ�-?�-��3&�(�,�mF�P{l��y���  �  "q��� �V�b�?��j��^���������$P����^f�Χ>���A��������$��#G��^o��R������|��R���ul����`���6���'+�~���l��fS`��<���$��O�}��dl��$�d����0�r�N���z��jȾ�� ��$���M��w�����`���qؙ�)�k���X�q�2�� ����w�ܜ��.�UT���|�Cl���T���P��L^���"|���R�J")�ؙ��ξ,��Ji����R���3�o4�����iK�� ���"��y9�	�[��������"�پ�'�A
2�� \�:[��JV���8���헿1����s��zK�{�'�N����l4�����:���a����^���H}��V��?=���n��pD�tC����=���u���J�o�M�F�,�+�tU�����/�Q������`)�:bC��Hj��9���o��p�����?�/j�x^��T����������<]f�3�>�*��`��������$��!G�]o��Q������{��ȫ��l���`��6�\�*�o���M���P`�L�<���$��L����h�,!��|��0�зN�z�z�=xhȾ� �u�$�d�M�_�w�l���-���Gؙ���j����X�e�2�� ��������Y�.�kUT�(�|��l��U���P���^���#|���R�=#)�ښ��ξb!���k��I�R�U�3�9���&���O��$�5�"��|9��[������c�پz(��
2�]\��[���V���9�������s�e|K�k�'�>����:6�Z����:���a�����ѵ���}�����{=��^�n�8qD��C��󾩘������o��G���+�AZ�y���4�)��z���d)�2fC��Lj�B;���  �  &D�����j�B�:��Dc����t��	s�����L��-�_��9����)��֞������ �ޯA�u5h��腿&���R���Վ�gO���\Z��$2��S�hݾ�ԭ�p���y�b�_�?�tK(�������#x��H��� ��4�,�Q��|�ǜ�
�ƾپ���"!��YH��Kp�r0������N���|;��b�x�֟R���-����p��6��A�rQ*�:TN���t��Ɗ��8��5��I����t�*�L��L%��[��̾�Р��/��ْU��6�g|"��2����"\��P��?&�:�<��-^��V���W��s׾˖	��-��U�B�|����U���Ⓙ�����ul�{�E��X#���
�� ��I����H�5��C[�Wf���܎�ZS������م�;�g��a?����J�07������q���I�/����ߥ�.:�G���!�Ī,�iF��wl�?x���B���������:�`Dc�������r������K��ė_�z�9���M���������� ���A��3h�$腿k��R��CՎ��N���[Z��#2�$S��fݾ�ӭ�S����b���?�xH(����1���t��D�+� �/4���Q�z�|��Ŝ�x�ƾe���*"!�YH�pKp�70��y���$���Z;��1�x���R���-������7��A��Q*��TN��t��Ɗ�9��q5������Ղt��L��M%��\��̾�Ҡ�22����U���6��"�W7�(��U`��T�[C&���<��0^�X���X��[t׾m�	���-���U�-�|���������㒿u���^wl�X�E��Z#���
�� �TK�0��ƙ5�<E[��f��Yݎ��S��#���م���g�-b?����2L�8��>��Ȥq���I��/����ڪ�-?�-��3&�(�,�mF�P{l��y���  �  ��G��t����-���P��p�^���T[�����hNm�8�L��Z+��C������%�]B ����A�2��sT���s��b��A��򬁿Jj�13I��L&��9�U�־������Mrk�3J���2�b�#�1l�S��]��+��>�z2[�����l��e�¾>+�:���9��.\���y�Kƅ�D�����~��c��zA��!�5���&�����]������=��_��|��G���L��VH|���_��}=�) �PE���|Ǿ(���`���_��MA���,�7 �	1����ZK"�Ҵ0��G��$g����i���؊Ѿ�����"�^NE���f�0���@
�����-�v��-X��66���������" �������'�I�l�i�p����>���k����s�y�T�S�1�Ph��`�z�����WNy���S���9�E�'�\�����8I&��27��P��t��8���������.�-�!�P�y�p�
����Z������8Mm���L�#Y+�B����2"�v@ ����n�2��qT�)�s��a���@��q���2Ij��2I�/L&�9�Z�־��������ok�}J���2��#��h�������+��>��.[�O���k��˭¾�)��s�9�R.\�/�y�ƅ����I�~�vc��zA��!�:���&��ߦ���C��t�=���_�"|��G���L��I|���_��~=�!�]G��Ǿh��@c���_�ORA���,�� ��5����SO"�y�0��
G��'g�H������
�Ѿ ����"�OE���f������
��7����v��/X��86���������#��B��"�'�_I���i�✁�X?��	l��6�s��T���1��h��a羊{��̃��\Ry���S�Õ9�J�'�-a�+��(��N&�e77��P���t�C:���  �  (�����پ��v��+8��P��3b���g��`��L��[2���� ���K��<پ1��_]����i�8� �Q�s�b�7�g� @_�O�K��)2�t���s����о�����듾�O~��X^��WF�R�5��u,���*���0��	>���R��
o����]������[v�"Q�O�%�j�@�e�W���e��f���Z�6_D��)�ވ�_��S�ܾ�O۾z
������%�zA�i�X���e��Nf�p�Y��C�	)��(��K�W�ľ����Hd��¬r��~U���?���1�+�m�+�UG4�FD��K[��Pz��V���[��֣̾SL�����,!/��=I�ڏ]��gg��d��#T�.�;�������Z��v�پ3�߾dg��0�ZA/�1�I�{\^��g��uc��IS�� ;�������޾"+��m��}��=h���M��h:�ڮ.�|{*���-���8�K�ʴd�vP��@K��������پ
�����*8�u�P�F3b���g��`�ĤL�/Z2�t��Ģ����ᾍ8پ��澕[�-���8���Q�$�b��g�0?_���K�A)2����	s����о�����꓾�M~�V^��TF���5�:r,���*��0��>�ĽR�o������l����t�pP���%���@��W�7�e���f�r�Z�_D�y)�ш�j�󾃎ܾ�O۾�
�@��#�%��zA���X�l�e��Of�5�Y���C��	)��)��M쾌�ľ� ���f����r�w�U���?��1��+���+�bK4��!D��N[��Sz��W���\����̾vM������!/�b>I�Ր]��hg�4d�"%T�͉;����i�����پ��߾�j�����B/�C�I�`]^���g�"vc�dJS�!;���� ��K޾�,��S��3���h���M��m:�E�.��*��-��8��	K��d�dR���L���  �  Gҽ���׾�������k�0�m\;�cr>�g�7��)�������}ܾ�žt>��{�Ⱦ�'㾎v������,�f6:�{�>�\w9�ǧ,��_�}��Q�ﾅ�Ѿ���3��l��B��k�e�W�Q�F���C�/nK�0�[��s�}툾�z��i����
ƾ����S'��P%�
�4��j=��W=���3���"����Q��?�Ҿ[����ܿ�� о���4w�l� ��72���<�"�=�k�5�l6'��5�?��&微�ȾU��В��龊���v��(^�}�L� ND��aE�z�O�gc��;}����]⠾R��2�ξ��뾬���S���*�J^8�Kv>�?*;�G�.����F����/˾�����fþ>�ؾ#m�������&�x�6�l2>�'<���1�hi!��
�.���P ۾����;穾�[��A[����m��yW���H���C�K�G��pU��k�3����X��+����н�`�׾������k��0��[;��q>�y�7��)����I���pܾ{ ž;���ȾZ$��t�<��w�,�45:�w�>��v9��,�_�
����ﾹ�Ѿ$���3���j���@��L�e�ݭQ�DF���C�jK���[���s�t눾�x������<	ƾz��6��&�'P%���4�fj=�PW=���3�x�"����4��H�Ҿ����ݿ� оE�w�� �+82�T�<���=�4�5�I7'��6�A �L���Ⱦ���D���k�����v��-^�l�L��RD�FfE���O�*c�#?}������㠾s��<�ξ���8��;T�E�*�/_8�Zw>�y+;���.�&�����S�澇˾֑��jþ5�ؾ�o��.����&�]�6�,3>��'<���1��i!�#������!۾���L驾�]���]��H�m�{W���H�\�C���G�8vU��k�~����Z�������  �  �Ӿ7X������(<�D^��d��^��S���v��$�ҾJ�������^���qb���ٽ�8�پ����@�
�L0����������7
��� �/E�C�߾^iϾ$X���T���7������y��di��of�9�p��F��D����5���m����Ǿ��ؾC�辦���:�\(��~���u�+�0 �~l羓nɾL����s������鲯��eƾ����{�����m����b��"��������Oھ�ɾ8j��
:��k��kȄ�͇r���f�eh�=�v�v����B��TK��#a���;0�ݾlb���#2	�����1�����*,�W?���	ݾ���m��Q¢��[���8����Ͼ�g�PN��J�E������B9��
�&���'�3�ԾD%ľg���+��"ގ�5e���Dm�#�e�Q�k��~�K��[+���a��9¾6Ӿ�V㾏��I��;��]�Od�^�S������Ҿr�������D���R_���ֽ�J�پ4����
�;/����0��j���7
�x� ��D𾙹߾�hϾ5W���S���6�����}y��`i�tkf�ڡp�sD������3���k����Ǿ��ؾ��� ������'�~�+������8l�tnɾT����s��N���h����fƾ���r|�g��`n�����D��#�����@��VRھ��ɾ�l���<���m��˄��r���f��ih���v�c���nD���L��^b����;�ݾQc�{����2	�����2�����l-�B���ݾ������dŢ��^���;��K�Ͼ4j�UO�cK� �������9�A�����)�2�Ծ�'ľ�i��b.��ᎾCh���Jm�V�e�\�k��~�����-���c���:¾�  �  ����i ����t3��1�C��vG ����Ț�/�ؾ5¾
������u���ֈ��~���~��͇���SǾ�=ݾ<�z,��X� �8���6��+��������3��0���
վ�\��6��9-���7��W$��xK���}���;���"˾��ي񾀙������R8��"�v|�O���>8��g���`Ѿ%���wӤ�^ʓ��8��س��0Q��G�������]�ξ������J����V���7�a��A�jt����l��'�;l���y��������z��������量qͻ�
�Ҿp��������H��$&��7�7��� �4#������v߾��ɾ����w��ۨ��z ��)������r[��Ǣ��"=־I��������������-�F5�0��� �`����@�ܾ�	ƾ�L��ʄ��&Ȉ��ꌾ٦���㬾�zþ��پ��X���Ai �S���2�b1�����F �j����9�ؾ�2¾��������s���ӈ��{���{��'���@QǾ`;ݾ]��*���� ����6��+�k������53��S���	վ}[��n4��S+���5��"��&I���{���9��? ˾��ƈ񾑗�����
��7�/"��{�`���y7�����z`Ѿۇ��VӤ�fʓ�9��/����Q��𤢾U���X�ξ���6������]W���8�t��B��v��+����;/���9���:����}�����������'ϻ�y�Ҿ��������������&�J8���u� ��$�����9y߾�ɾf����y������V��񚋾n���]�����!?־�龐���L���I��P.�6���� �����C��ܾ�ƾ�O�����u�}ˈ��팾򩙾�款N}þO�پ���  �  ���;�_������� �:p�*ҾC��P`���.��
7����|��*k�f�Mn�z���ȏ�|/��{k��0ž]�վ��S�����'���z����%��z�������(!ξ{���ԥ�Z󢾺⬾�¾�޾��������d������t���������r�ݾ��̾3e���G��K���(����u��g�`;g�P�s�Đ���_���>���i��z�ʾ47۾~�����������*f���_��)��� �c3⾂�ľ'���cl���ݤ��в�p�ʾ�*����(���L�����*������������羐�׾�Ǿ"l���1��i���������o��;f���i�Hz��z���1��W���P��zSо�ྌ6�jz�C�
��*������Ⱦ�X
����s�׾`��ƛ��[t���1���湾�ԾP��Q�����$���:������������n⾞(Ҿ�A��w^���,���4���|��%k���e�n����hƏ�N-���i���ž�վ�澥���؎�����z�[�������c����oξ}���ҥ���AାE¾��޾w���o���c������s�=��j����q�ݾء̾�d��1G��2K���(����u�h�g�<g�Q�s�o���^`���?���j����ʾ�8۾0�뾿��������[g�@����*�� �H6�e�ľ����o��JाӲ�{�ʾL,龬�����CM����=+�Ԯ�o��n������׾EǾ*n���3������ �����o��@f���i�Mz�}��4��Y��VR��Uо���8�,{��
��+�����%���
������׾􂼾e����w��_5��깾��Ծ!�󾑘�����  �  }�>���:�2/�Uj��������s_־k~���u��\��|Ƃ�w�i�,{T��hG���C���I�?�X��eo��>��b��7������`�ܾg�����f"�~\2���<��>���5���%� f�`B��uA׾��¾�Ͼ��3̾4�������/���;�]>���7�1�)�)M�n���7꾓@;_Ŵ�̟�>���ߠ{���a�{"O��E�щD��M��\_��tx�Ŭ�����H��FRʾM�澙��~=��%(��6�>� b<��c1��c�kH
���G�ξhs���d��M7Ծ��� ���#�I�4��=��$=���3�5Z$���& ��ྀ�ľ2p��#o������Tr�+�Z�W�J��C��F���R�?�f����+c���2��r޹�EӾP��	�vc�k�-�-�9�S�>���9�n�+��{�FO�@Sᾃ�Ǿ�%����ž��ݾ�
�"��*���8���>��:�k1/��i�i������:^־}��Lt��ZZ���Ă�6�i��vT��cG��C���I���X�9ao��<��p`�����v�����ܾ�f��y�wf"�q\2�ۂ<��>�_�5��%�Ge��@��]?׾[�¾L;��0̾������z�ɬ/�~�;��[>���7�L�)�\L����P6꾐?;�Ĵ�]˟�Ì��?�{���a��"O�E���D��M�:^_�Pvx�ȭ��0���cI���Sʾ	�澏���>��&(�S�6�j>�cc<�2e1�e��I
���=�ξ>v��-g���9Ծ9������#�ю4�q�=�%=���3�lZ$�# �� �����ľ�q���p����LYr��Z�E�J��C���F�F�R��g���e���4��๾�FӾ�Q�v�	�[d�m�-�S�9���>��9�,��}�"Q�W�f�Ǿ�)��[�ž-�ݾf��#�S*���8��  �  �g���a�k�O��6��c�Ѯ�5Z׾-ѳ�L헾�A���c���I���7�Qz-���*��(/�7L;��N���i�e���ԉ����Zf྇�xm!�g�<�sqT��d��lg��|]��H�[�-�����`����޾��پ�&���
`!� 
=�tMU���d�2g��\���G�B�-������%�ʾ�������^x��Y�cC�H�3���+��9+��\2�	�@�=�V�7�t�����������ƾ�����6�*��&E���Z�M�f���e�W�W�z@�<m$�'�
��W���ھ?Fݾw�������*���E�ݡ[���f�$e��V��?��w$���	���6���ru���ވ�[?m��fQ��=�0�'�*���,�h6��wG���_�2+��3;��\����Ҿ����e���3�c*M��	`���g�3b�H�P�X�6�PY�T/� z�cپ��� ��f�Y�3���M�X�`��g��a���O�{�6�0c�@��Y׾�ϳ��뗾R@���c���I���7��u-�6�*�)$/��G;��N�L�i�Ꙇ�����C���e�d�qm!�o�<�{qT��d��lg��|]���H���-����^��T�޾��پ�#�h��^!��=�'LU�O�d��0g��\���G�m�-�������ʾ����_���]x�_�Y�C�O�3��+��:+��]2�c�@���V�B�t�ě�����L�ƾ~����K�*��'E���Z���f���e�׈W�@��n$���
��Z���ھIݾ�y�������*�A�E�_�[�N�f�\e��V��?��w$���	���K����v������ Cm��jQ��=��#0�ӭ*�\�,��l6�#|G���_�-���<���]��k�Ҿ0���f�u�3�w+M��
`�f�g��4b��P�8�6�J[�_1�?~�x!پ�� � ��h���3�%�M���`��  �  _��'��3o���N��,��>���޾uﲾ%����1r���N�#6�r�%�O���������(���:�c�U���{�3��M���`F�1)�T�3���V��Xu�̄��&��7���Kh��.G��#&��x��������1�|8�G	Z��x�Lr��]冿K ��W'e�T[C�� ��Z�P�ξ��������Ve���E�6�/�/�!����Y��� ���-�B�B��`�P���颾��ɾa��Z���q?���a��}�ʅ�����D�z���]�Q�;��G����n���j	���"�D`C���d����ᆿay��r:x��VZ��7���+��T��¦���j���RY��Q=�}:*������Ʈ�n1$�j�3���K�P�m�#��e����tپ���1(��"K���k� 0��FQ�������r�W�R�_�0��U������������-���N���n�����^���&��]2o�B�N�,�7>�\�޾+����R.r�L�N�P6�f�%��J�������ŕ(���:�1�U���{�2�������E�")�a�3�͚V��Xu�̄��&����Kh�.G� #&��w��������{0�	8��Z�;x��q���䆿���_&e�xZC�S� ��Y�;�ξ��������Qe�ގE��/�4�!�q��oZ��� ���-���B�� a�����iꢾ-�ɾ�b��Z���r?�+�a�^�}�|���U����z�M�]���;�'I�t��{�h���	��"�.aC�F�d����&↿wy���:x��VZ��7�P���+��U������+l��nVY�vU=��>*�I����5���5$���3���K�
�m�倎����Tvپ����2(��#K���k��0��R��a����r�O�R�q�0�X� �����7������� -�,�N���n�{���  �  �v������V'���a��8���s��Hٴ�6���)�i���D���+�u�O��8F��
��[��D0�f�K��Lt�����¾�������A���i���u��8��+>��l�~��Y�m�3������pM �@���%�{�G���n��n��D��"甿t䌿�z�5�S���+������Ծn(��s�8�[�%$;��F%����+������e#��98�n�W�����W䢾��ξj"��g'�O�S�v��y���w��C}����r��0L�#�(���� ��������/�g�T���z�팿s锿5?���b�� *n�[F����Q����þ�Κ���y�k�O�F�2�������_���U ��V)�L]A��e�#C��O ��q྾8��R4���\�gE��n���e��ϔ��Y���f�V�?�s�h�dv��1p��Z�܌;���a�%9��Ӓ��Sv��>����&��Ra�[�8�^�I��ش�ͳ���i�O�D� �+�1q�C��'B����W�3A0�b�K�iJt�	���s���3����2�A���i�����u��8��>����~�%Y�t�3�V��9��L ����@%���G�-�n�n��fC���政�㌿�z�T�S���+����Ծ�'������/�[�x#;��F%� ��b+�~����{f#�~;8���W����墾��ξS#��h'�0O���v�mz��mx��F��&�r�=2L�ʈ(�S��� �������/�T�T�P�z�S팿�锿G?���b��	*n�oF����R����þК���y�ĚO��2����9��gc�<��$��Z)�2aA��e��D��"���rྛ9��S4���\��E���n���f������J���f�x�?�:u����z��Qr��\���;�S�a��9��w����  �  A��]�濞οw��$?��$[S�{L ������7m���gv��S��P>���2�R�/���4�v*B�'FZ�'���˜�˾ƾ-O�]�*�Dm`�搿uN��3�Կ>꿉6�}O�+ǿc1��Hf��&�U���7��L2�'�E���o����j��z�׿�����߿9tÿ�����H|��@���l�޾􈭾�~��,i�7jK� n9��0��I0�G8�[�H��)e�sv��E��huؾ���;�u�ޡ������c@ݿ���}�쿑�ڿ�/���ř�i�u��&I�d83�^�5��9Q����[����ÿB�߿�����׿-��|Ȕ�2/g��/�,K�nk̾ѷ���˂���]�DD�:�5�c�/���1���<�J�P��q�E���I���[�j��M�&}��������ʿW�����!z��aѿ����Ď���d�x+?�F]1�7m<�v[_��:��笿�ο?�濳����@ο�v���>���ZS��K ����a
���k��(dv�S�S��L>���2�2�/��4��&B��BZ�%���ʜ��ƾ�N�B�*�Sm`�#搿�N��U�ԿT꿉6�_O��*ǿ 1���e���U�R�7�OK2���E�L�o���Ji����׿��t���߿�sÿ2���H|�V�@�]�|�޾8���M~��Z+i��iK�n9�C�0��J0�T	8���H�a+e��w������vؾ���;�+u�s���o¿�Aݿz��E��c�ڿ_0���ƙ�%�u��(I�:3���5��:Q�y���[����ÿy�߿�����׿
-��|Ȕ�N/g�R�/��K��l̾@���{͂���]�7HD���5�Ŵ/�,�1��<�p�P��q�(�����e]��j��M��}��K���2�ʿ�俒��{��bѿð�CŎ�
�d��-?��_1�to<��]_��;���笿�ο���  �  �����ݿ��ƿ����kJ��{N�S��)���L���ᖾ�tz��>X�1�B�E�6�L�3�u�8�F�}�^���u��Ȟƾ� �%�'�t�Z�����q2����̿�H�a!�}�ٿ����ş�	����&P�y�3��A.��@�ti�nX�����غϿ8����/�׿����y���tu�/�<�c.�P�ݾ�F��"3��gm��O��=���4��c4�}B<�SDM��oi�Y<��9�����׾���[Q7��n�����'���տ�����㿪}ҿG����䔿��n��(D��#/���1���K�F�z�1��������׿��>��٭Ͽ�ޱ��A��_a�c�,�L��b̾'ۡ������b�$�H��9��3�6�b�@��DU���u�����n����꾥�LwH�����9���Zÿ|�ۿVr�Q�߿��ɿ
Ȫ�Mf��%j^���:��[-�s�7�)jY�m�����ʪƿ��ݿ�濁�ݿ@�ƿ<���#J���zN������`K��_���0qz��:X�-�B��6��3�]�8��|F��^����1��֝ƾ@ ��'��Z�Đ���2����̿�H�_!�^�ٿh��^ş������%P��3�E@.���@��i��W��;���Ͽ���R�応�׿����x��tu���<��-�a�ݾ�E���2��cfm���O��=��4�Pd4��C<��EM�Qqi�j=��|���k�׾���LR7��n��������Gտf�俶��{~ҿ����唿D�n��*D�G%/��1�E�K�o�z����宼���׿;��E��խϿ�ޱ��A��3_a���,�����̾�ܡ�����tb�K�H�d�9�{�3�r6���@�(IU���u�񄓾Pp����꾂�0xH���������Zÿ0�ۿ%s�9�߿��ɿɪ�ng��vl^��:�9^-���7�ClY�f�������ƿA�ݿ�  �  ��ͿS�ƿ,����k��
�u��A�E{��0����_��a��bnf��6P�+�C�DS@�B�E�=DT���l�0ň������Ǿ?����  ���L���}ȝ��㷿�eɿƇͿ,ÿoج��Ȋk���@�Ԗ'���"�,3���V�m������K��L�ʿ�Ϳ������ƍ�Sbc�Ǎ2�B����ܾⱾP���w{���]��K���A�!A�_�I��A[���w�:�����+!׾���6�-���]�)�����������h̿[�˿8���Aأ�������[�$76�2�#��&��=�:f�vō�l穿�
��Ϳ��ʿ^���렿 ,���R��s$��� ���̾ׄ���?��'Bp��uV���F��x@�!�B��YN��kc�^����:���1��b辏g�x�<��eo�6���د��Ŀ�Ϳ�ȿc3���u����|��HM���-�Y"��w+���H���v��I��r���+�ƿH�Ϳ�ƿϞ���k��z�u���A��z��/���s]�����yjf��2P�߽C��N@���E�+@T���l��È������Ǿ�����  ���L�#���ȝ��㷿�eɿ��Ϳÿ.ج�~ˉk���@�~�'�=�"��*3��V�Yl��W���'K����ʿͿv��p��2ƍ��ac��2����ܾ͗f᱾�O��w{�;�]��K���A��!A�k�I�C[�P�w�J�������"׾���$�-��]�����{�������i̿�˿���٣�w�����[��86�ȭ#�F&�=�^f��ō��穿�
��(Ϳ��ʿ^���렿),���R�	t$�� �%�̾d���hA��,Fp�DzV�"�F�\}@���B�a^N�-pc�b⁾�<��h3���ih�W�<��fo��6��ٯ���Ŀ��Ϳ�ȿ[4���v����|��JM���-��"��y+���H���v�{J��3���Їƿ�  �  �g��<ꦿ|̗�\���CZ��I2��.�>���
Ǿ�慨����趀�>i���Z���V�"]�j�m����e���򮾒�ξ����D���:�q�c��퇿�͛�6�����_ţ��V��Ԋx�D#M�]�*���7�����O<���d��̈�뜿ù��ѫ��Ƣ�+I��	iw�XJL�n&����++ྥ����������5x�9c��VX�X�W��a� bu������������۾���֧"�L�G��|r�� ��-��mU��N���Ȟ�>����i�0P@�`�!���������'���H�P�s����Q7��糫���������sR���h�S�>��d��T���Ӿ���혾�߅��p��s^�w�V��Y��g��7~�}ŏ����PFþ���W��*>.�/�U�����߯������Y������阿҃���Z�Q�4������:��,1�	AV�UO��oʖ�:���Zg���馿 ̗���CZ�I2�G.���N	Ǿ�����۴���i���Z�*�V�x]��m����������\�ξ��������:�w�c��͛�;�����9ţ��V���x�O"M�:�*���T6�N��&N<�6�d��ˈ�iꜿ ���qЫ�nƢ��H��+hw��IL�em&���G*�����������I5x�9c�
WX��W��a�ccu�գ����T�����۾�����"�Q�G��}r�����-��!V������Ȟ��>��S�i��Q@���!�R��b����'�ܽH�9�s�����7�������������~R���h���>�.e��U��b	Ӿ����	ⅾ�p��x^�BW���Y��g�T<~��Ǐ����HþO��,��?.��U�/���o�������bZ����꘿|Ӄ���Z�u�4�"!���-<��.1��BV�'P��(˖�ه���  �  ?ɉ������y��N^��6A��r&����Wi���t۾��������������~�>�x��|��Z⊾+���/���}ƾ�����u��,���G�\�d�@�~�v�<n�����jl�K�K�x+�7_���e��������	=��^^�h�{�􈇿撉��g	q�8�T���7�j�&0	�̀�s-Ҿ.ݸ����J���^����z�Z	z��H�������頾FD��X.Ͼ� ��a��;�4�LQ��n��悿�M���&��%�~�P�a���@�d�!���
�'��� � ���a)(�7H��i��恿���m}��������g�o�J���.���� �N5�dVɾ05��i����a���U���y��|�����Mܔ������-��dNؾ����1���#��>�[�`�v��ǅ��ω�q���v�W�:�5������С���*�`��M2�DOS���r�l���ȉ�����H�y�EN^�L6A�Lr&����g��s۾����!�軖�x�� ~�E�x�ez���ߊ��)���_{ƾ5�ᾈ�iu��,�j�G�X�d�@�~�o�'n�����ljl���K�.w+�"^����ɞ�����H���=�i]^� �{�Z���V���Dyq�e�T�"�7�si��/	����,Ҿ�ܸ����lJ���^��J�z�
z�)I��d���l꠾PE���/Ͼ2���E��9�4�+MQ��	n�H炿�N���'����~���a���@���!�x�
����~� ��t*(�H��i�灿����}��ɢ���g���J���.�������6�HXɾT7������ud��vX���y���|�VĆ��ޔ�ٟ��}/��.Pؾ,��������#��>�[�l�v�Aȅ��Љ�8���v��W�-�5������ҥ���,��a��O2��PS��r����  �  ҴW���V���M�5@�r�1��v$��u�	��4�55��yϾ0w��i񣾤���*ߓ��������������#վ���D��˔��
��N'�x�4��]C�6P�a�W�;�V�F-L�d�9��_"��N��$�%�ھ�U־�徿:�����/���D�I-S��VX�V@T�1iI� e;�7-��U �����+	�d)��ڗ�i%ǾQ���垾B�������g��&��rmľ��ݾ�^�����__����ٴ+��9���G�PS��NX�C:T���F�s2�r��d����o	׾�)پ��������7�tJ�&�U���W�u7Q���D��6�_�(�X�w���;�ھ���׾����ũ����F	��Q���
)�������̾�U����~���-�u#��F0�N�>�8L�^�U�{X�n�P��r@��N*�����7��*�6�վJ޾�X���0���'�;4>�LNO��W��V��M�y4@���1�Qv$�5u�Q��3�R3��wϾ�t����}��tܓ�牙����z����!վ���k����
�WN'�B�4��]C�P�<�W���V��,L�ل9�*_"��M�v"�ܒھ�S־]��s9�k��̄/�p�D�&,S��UX�^?T�QhI�8d;�a6-��T �}���+	��(��`��%Ǿ�P���垾3B�����dh�����Knľ��ݾ `��{��&`����е+��9���G�VQS�'PX��;T���F��2��s�`f���:׾P,پc����j��Y7��tJ���U���W��7Q�C�D�_�6���(��X�9���<����]�׾%��Eȩ�ۻ���������+�����۬̾|W澪���M���.�3#�eG0�'�>�9L�x�U��	X�ܶP�Rt@�7P*�̵�];���-��վ�޾\��X2��'��5>�iOO��  �  b�*�.�/��1��1�� 1��0��a/��m*�� ��9��|��Ⱦ�'������5��^Sξ��r��{�Wq#���+���/�Y1�1�2#1�F�0���.�W,)�i���}�.���a߾�+žU_��ie��ꬼ���ҾG��Y<	�_��_.%�I�,��N0�S 1�1�h$1��0�[/.�#�'����L���'��>rھĸ��X򳾏3��0���"D׾q�����<=��&�d�-��0�##1��1�>"1��|0�l-�0C&��x���f���Ĵվ����Ⲿ
`���¾�ܾ$��j��:w�9C(��i.���0�+$1�u1��1�l30���,���$����M���\1Ѿ�û��2���굾`ƾ�ᾟ� �D^������)��/���0��!1�.1��1�$�/�ӌ+�D�"�,��(�����@�̾�G��iⱾѷ�
5ʾ�5�8��D����!��*�n�/��1��1��1�t�0�Fa/��l*�>� �����y�K�Ⱦ%����;��sPξ!���p��z�Zp#���+��/��1��1��"1��0���.�,)����<}�����Y_߾�)ž-]��c�������Ҿ���,;	�>��N-%�K�,��M0��1�U1��#1�Q�0��..���'�C����Q'��rھ˸�����3�������D׾�q��}���=���&�'�-���0�$1��1�X#1�~0�Hm-��D&�z�^�>�����վՖ��2岾�b��L�¾�ܾ���!���w��C(�:j.���0��$1��1�T1�$40���,� �$�!�;O���M4Ѿ�ƻ��5�����bƾN��� �E_����K�)�o/���0�~"1��1��1�#�/���+���"��������龯�̾2K���屾tԷ�>8ʾ�8澓��x��˒!��  �  n��.�+%���2�� A�K4N���V��~W��N��=�IZ&�����|��� ݾ��վ2N��:��'���+���A��_Q�v(X�~U�a�K���=���/�`a"������%O�����=H˾�ҳ��P��cA��-���\���Ҫ�Sm���kپ�)�����z�g ��|)��`7�G�E���Q�PX�{�U��I���5�5f�;��7쾾�ؾ�|׾�-�8������Y3�G�G���T��@X�6�R�2G�T�8���*��Q�?���5�~���Gܾ�þW���`���΃��a�������w����Ⱦ8������	�'F��!�X�-��2<�� J�O�T�NX��R���C��9.����*�~���־]۾S�򾧁�x�#�a�:�3�L���V�|VW�OtO���B��04�N�&��c�]���:�|��Ӿ9����������Г����ڤ�����,�оS��F�����z�s*%�i�2� A��3N���V�~W�7�N�s=�Y&�f���y���ݾx�վ�Jᾘ7�������+�9�A�s^Q��'X�U}U�ǈK�M�=�R�/�a"�6��C�7N������F˾ѳ�$O��Z?���*���Z���Ъ�k���iپ�'�����y�����{)��_7���E�N�Q��X��U�ӍI���5�f�+���7��ؾ�|׾).龍��H��Z3�ۯG�5�T��AX�
�R� 3G�P�8���*�S�t���6�����Iܾ�þ
������X���Đ��ʮ���x��D�Ⱦ��P���g�	��F�l!���-�b3<��!J�%�T�OX��R��C�R;.�x��=,����־`۾3�������#�h�:� M���V�'WW��tO�3�B��14��&��d�c���;��~��Ӿ<���Ħ�R���ԓ�<���ݤ�c�����о���?���  �  pK�������'��B���_���z�"������u���^q��sQ�Œ0��l��G���f��v�w�7��X�_�w��m���ʉ��Y��gu�rY�փ<�_"�Jp�`�����־�ּ��y�����#���8|��;y�!́�#+��Ժ��bv��c�ʾf�������j0�~mL�Hni��9������ 爿�K��zFg��@F�2�&����sX ��8�����_#�*�B�q�c����^m���"���[��X�l���O�%_3�����
�
G��;`���7՟�9Î��Â�(�y�<6{���(��6���,��ȰӾlF�@B
���m9�0V�7�r��l��Q����/��H�z�Q�\�-6;�R�X��?���J�9���%-�w�M�Gn�����>�������ً}��c���E���*��E�� ��Cྛžk���ͥ���$�����a�x�%�~�����ΰ��u ���G¾N
ݾ�I��P���'���B��_�K�z��􆿨��������\q�RrQ�R�0����������Pd��t�ś7�i�X��w��l��ʉ�Y��Nfu�xqY�_�<��^"��o�������־|ռ�cx��H�/"���4|��7y�ˁ��(������Nt��d�ʾ���� ���j0��lL��mi��9��X����房�K��DFg��@F�$�&�����X �&9����e_#���B���c����m��P#��Z\��:�l���O�-`3������xI꾇�;�����ן��Ŏ�5Ƃ��y��:{�򄾳*���7��Z.���Ӿ�G��B
�����m9��0V� �r�Km��᫉��0����z��\��7;��S��eC��-L�����&-���M�Tn�������������f�}�* c�/�E�M�*��F�| ��E��ž
��������'�����R�x��~�i���b����"���I¾ݾ�  �  �����W4���\��K���Ә�t����`���⥿f������+�S��w/�,]�����&���6�MZ]�����򙿗F���E������(���C�~��5S�B,�>b�F4�0q������������|��f��rY�1&W��._��cq�̆�-(������$վ� ��,�A��#k���������M[���u���e��1؎�� q��F�q&��8�fB��O#��_B�Sl�@t�� ����ު��
���V���؍�Xp�ɅE��� �E`�fqپi����������St���`�߃W�~�X�vd�<�y�����衾ؽ��y�FK	�KY(�=�N���y�h��$���� ��F���򛿾����+b��Z:��V�Y�����7(,��_O��{��y��	����6��ܔ���Ԛ����]oa�R�8�/��D��\�̾�f��b[���7���ul��}\��V��W[�0j���������e����Ⱦv�\���V4� �\��K���Ә�!���o`��O⥿г�������S��u/�`[�ץ��$���6�xX]����(��E��*E�����������~�5S��A,��a�O3�p������0�����|�*f�	oY�F"W��*_�z_q�ʆ�2&�����G"վ� �2,�WA�F#k�G�������[���u���e��؎�� q���F�v&��8��B��O#��_B��l�}t��H����ު�F��QW��iٍ�G	p�ʆE�� �fa��sپ����.�������Nt�{�`���W��X��"d��y����� ꡾Xٽ�{��K	��Y(���N���y�rh������(���F��r󛿚����-b��\:�lX�*������),�6aO�A{�z��y���=7��%����Ԛ�X����oa��8��/�;F��L�̾ i���]��n:�� {l�(�\���V�O][�A5j�b�������g��Z�Ⱦ�  �  nN񾰐�mD�q�x�4������Pǿ��Ϳ��ſ�������?t�e�F��h*��4"�v/���O����2�������ȿӰͿ/�ÿ n��㚒�B]l��:��j��)���q���pЀ�j�a��|M���B���@���G��W�
r�D���-T��PMϾے�/�&���T�)Å�xy������˿��̿����i��U2���ec�<;��W%��*$�2�7��+^�=��>a���Ͻ��̿�̿�ܽ�M����􈿕�Z�u[+�H�xԾ	��@(��ڬu�� Z���H���@���A�~�K�#0_��x}�����泾Lf߾X��e5�fZf�ob��̈��'¿�PͿ�ʿ���m/���傿�<T��1���"��u(���B��Sn������I���ÿ�Ϳ(�ȿ ����3����~���I��������%}ž�K��T���u+k�A0S�*-E��C@��0D��)Q���g�7��%�������M����lD���x����l����Oǿ��Ϳ|�ſB�������t���F��f*��2"�u
/���O����G
������\�ȿ-�Ϳ��ÿ�m�������\l��:�!j��(����3���π�U�a�ByM��B���@��|G��W�/r�\���XR���KϾ��o�&���T���2y��Ə���˿��̿�����h��E2���ec�<;��W%��*$�r�7��+^�p��{a��,н��̿̿"ݽ�����D�����Z��\+�b�fzԾn���*����u��Z���H�p�@�G�A���K��3_�&|}����`賾�g߾���5�[f��b��D����¿IQͿ�ʿ���W0��z悿�>T�ټ1�s�"�iw(�B�B�Un�2���@J����ÿu�Ϳl�ȿY����3��l�~��I��������~ž�M������]0k�i5S�q2E��H@��5D��.Q�0�g�'9�����,����  �  �1���" ���Q���m����0ȿ��޿���ݿ�ſJG��b^��2W�X�6��z-��<�
a����{����U˿>���O�y�ڿO���H������E����w���p㑾L�s���S��@�~�5���3��[:��I�4�c����'ӣ���ξD��SA/�g�d��������>ѿnG�:=��]ֿ��M����w���I�)1���/��E�
�q�����n��;�ӿ�`�hZ��ӿJ���ו��Dk�a�4�P�	��Ծ�ާ��̈�S�g�:L�O�;�14�5�Ek>�PQ��ro�湎��~����ྺY�ù?���x�fZ��M��@�ؿ1�忺�=Kο�@��ƕ���Yf�c?���-��4��^R����n���������ڿ�Q�t���F˿�X��9���t�W�_%�Xo��,�þ�1�� Ԁ��\��wE�,8���3��?7�b�C���Y���|�����\̾�{0��m" ��Q����4���W0ȿV�޿���Lݿ6ſ�F���]��aW�f�6��x-�t<�� a���������T˿u��=O���ڿְ�����a���E�{���v����.⑾��s���S��@���5���3��W:�C�I�d�c����]ѣ���ξy���@/���d����I���ѿ:G�=忱]ֿ���L����w���I�B1�ܲ/�M�E�]�q�J���%o����ӿ�`��Z�f�ӿzJ��ؕ��Ek�j�4�f�	�c�Ծ�৾ψ��g��L���;��54�f5�Ho>�Q�8vo�n������.��]Z�k�?�r�x��Z���M��Եؿ��忂�Lο�A��Ö���[f�g?���-�̐4�h`R����������A�ڿ�Q濶��G˿�X��l�����W��%��p����þ�3��Pր���\��|E�(18���3��D7�.�C�L�Y���|�Y����;��  �  �/��R�"�+�V��$��qo��Q�Ͽb����s��fd̿����~����\��,;�F}1�C�@��Lg�
���?���?�ҿ1V鿢h�"n�
�ȿL���֡��w�I���r�辸����L����o��xO�s�;���1�m�/�n(6�PbE���_��+��C���PXϾ�V���2�z�j�n�������ٿ8��E��޿�����r��-�/O��05�}�3��K���x�������ۿJ]�^Y�,�ۿ]⽿W���h�q��68�:���[վn릾�����9c���G��^7�a0�&�0��):��L�	>k���0ԯ�� �2b���C����k���UEſ��?����꿑ֿ=���14����l�(�C��1��8���W�������F�ȿ�t�hi��O���ҿQ[��)����]���'�ۻ����þ2㚾y�}���X�\#A��4��/�3��6?�WcU���x�4������L.����"���V�r$��8o���Ͽ�翧�����c̿���:}����\��*;�9{1�+�@��Jg����G���Z�ҿeU��gￍm㿏�ȿ燦�������I�c�Y�辐����K���o��uO�&�;�<�1���/��$6��^E�ʁ_��)��}����VϾ/V�֞2�Мj�!���W��Yٿ�7쿧E���޿�����r�� �5O��05���3��K��x�!������]�ۿ�]�Y��ۿ�⽿˩��`�q��78�O���]վ����t>c�>�G�,c7��0�j1��-:���L�iAk�����կ��!��b�U�C�w��֑���EſD�����sֿ2���25����l�2�C��1���8�E X�M��F����ȿu㿾i�P��ҿ[��[���r]�P�'�D�����þ!嚾Ⱦ}�P�X�E(A��4��/�3�W;?��gU���x��5������  �  �1���" ���Q���m����0ȿ��޿���ݿ�ſJG��b^��2W�X�6��z-��<�
a����{����U˿>���O�y�ڿO���H������E����w���p㑾L�s���S��@�~�5���3��[:��I�4�c����'ӣ���ξD��SA/�g�d��������>ѿnG�:=��]ֿ��M����w���I�)1���/��E�
�q�����n��;�ӿ�`�hZ��ӿJ���ו��Dk�a�4�P�	��Ծ�ާ��̈�S�g�:L�O�;�14�5�Ek>�PQ��ro�湎��~����ྺY�ù?���x�fZ��M��@�ؿ1�忺�=Kο�@��ƕ���Yf�c?���-��4��^R����n���������ڿ�Q�t���F˿�X��9���t�W�_%�Xo��,�þ�1�� Ԁ��\��wE�,8���3��?7�b�C���Y���|�����\̾�{0��m" ��Q����4���W0ȿV�޿���Lݿ6ſ�F���]��aW�f�6��x-�t<�� a���������T˿u��=O���ڿְ�����a���E�{���v����.⑾��s���S��@���5���3��W:�C�I�d�c����]ѣ���ξy���@/���d����I���ѿ:G�=忱]ֿ���L����w���I�B1�ܲ/�M�E�]�q�J���%o����ӿ�`��Z�f�ӿzJ��ؕ��Ek�j�4�f�	�c�Ծ�৾ψ��g��L���;��54�f5�Ho>�Q�8vo�n������.��]Z�k�?�r�x��Z���M��Եؿ��忂�Lο�A��Ö���[f�g?���-�̐4�h`R����������A�ڿ�Q濶��G˿�X��l�����W��%��p����þ�3��Pր���\��|E�(18���3��D7�.�C�L�Y���|�Y����;��  �  nN񾰐�mD�q�x�4������Pǿ��Ϳ��ſ�������?t�e�F��h*��4"�v/���O����2�������ȿӰͿ/�ÿ n��㚒�B]l��:��j��)���q���pЀ�j�a��|M���B���@���G��W�
r�D���-T��PMϾے�/�&���T�)Å�xy������˿��̿����i��U2���ec�<;��W%��*$�2�7��+^�=��>a���Ͻ��̿�̿�ܽ�M����􈿕�Z�u[+�H�xԾ	��@(��ڬu�� Z���H���@���A�~�K�#0_��x}�����泾Lf߾X��e5�fZf�ob��̈��'¿�PͿ�ʿ���m/���傿�<T��1���"��u(���B��Sn������I���ÿ�Ϳ(�ȿ ����3����~���I��������%}ž�K��T���u+k�A0S�*-E��C@��0D��)Q���g�7��%�������M����lD���x����l����Oǿ��Ϳ|�ſB�������t���F��f*��2"�u
/���O����G
������\�ȿ-�Ϳ��ÿ�m�������\l��:�!j��(����3���π�U�a�ByM��B���@��|G��W�/r�\���XR���KϾ��o�&���T���2y��Ə���˿��̿�����h��E2���ec�<;��W%��*$�r�7��+^�p��{a��,н��̿̿"ݽ�����D�����Z��\+�b�fzԾn���*����u��Z���H�p�@�G�A���K��3_�&|}����`賾�g߾���5�[f��b��D����¿IQͿ�ʿ���W0��z悿�>T�ټ1�s�"�iw(�B�B�Un�2���@J����ÿu�Ϳl�ȿY����3��l�~��I��������~ž�M������]0k�i5S�q2E��H@��5D��.Q�0�g�'9�����,����  �  �����W4���\��K���Ә�t����`���⥿f������+�S��w/�,]�����&���6�MZ]�����򙿗F���E������(���C�~��5S�B,�>b�F4�0q������������|��f��rY�1&W��._��cq�̆�-(������$վ� ��,�A��#k���������M[���u���e��1؎�� q��F�q&��8�fB��O#��_B�Sl�@t�� ����ު��
���V���؍�Xp�ɅE��� �E`�fqپi����������St���`�߃W�~�X�vd�<�y�����衾ؽ��y�FK	�KY(�=�N���y�h��$���� ��F���򛿾����+b��Z:��V�Y�����7(,��_O��{��y��	����6��ܔ���Ԛ����]oa�R�8�/��D��\�̾�f��b[���7���ul��}\��V��W[�0j���������e����Ⱦv�\���V4� �\��K���Ә�!���o`��O⥿г�������S��u/�`[�ץ��$���6�xX]����(��E��*E�����������~�5S��A,��a�O3�p������0�����|�*f�	oY�F"W��*_�z_q�ʆ�2&�����G"վ� �2,�WA�F#k�G�������[���u���e��؎�� q���F�v&��8��B��O#��_B��l�}t��H����ު�F��QW��iٍ�G	p�ʆE�� �fa��sپ����.�������Nt�{�`���W��X��"d��y����� ꡾Xٽ�{��K	��Y(���N���y�rh������(���F��r󛿚����-b��\:�lX�*������),�6aO�A{�z��y���=7��%����Ԛ�X����oa��8��/�;F��L�̾ i���]��n:�� {l�(�\���V�O][�A5j�b�������g��Z�Ⱦ�  �  pK�������'��B���_���z�"������u���^q��sQ�Œ0��l��G���f��v�w�7��X�_�w��m���ʉ��Y��gu�rY�փ<�_"�Jp�`�����־�ּ��y�����#���8|��;y�!́�#+��Ժ��bv��c�ʾf�������j0�~mL�Hni��9������ 爿�K��zFg��@F�2�&����sX ��8�����_#�*�B�q�c����^m���"���[��X�l���O�%_3�����
�
G��;`���7՟�9Î��Â�(�y�<6{���(��6���,��ȰӾlF�@B
���m9�0V�7�r��l��Q����/��H�z�Q�\�-6;�R�X��?���J�9���%-�w�M�Gn�����>�������ً}��c���E���*��E�� ��Cྛžk���ͥ���$�����a�x�%�~�����ΰ��u ���G¾N
ݾ�I��P���'���B��_�K�z��􆿨��������\q�RrQ�R�0����������Pd��t�ś7�i�X��w��l��ʉ�Y��Nfu�xqY�_�<��^"��o�������־|ռ�cx��H�/"���4|��7y�ˁ��(������Nt��d�ʾ���� ���j0��lL��mi��9��X����房�K��DFg��@F�$�&�����X �&9����e_#���B���c����m��P#��Z\��:�l���O�-`3������xI꾇�;�����ן��Ŏ�5Ƃ��y��:{�򄾳*���7��Z.���Ӿ�G��B
�����m9��0V� �r�Km��᫉��0����z��\��7;��S��eC��-L�����&-���M�Tn�������������f�}�* c�/�E�M�*��F�| ��E��ž
��������'�����R�x��~�i���b����"���I¾ݾ�  �  n��.�+%���2�� A�K4N���V��~W��N��=�IZ&�����|��� ݾ��վ2N��:��'���+���A��_Q�v(X�~U�a�K���=���/�`a"������%O�����=H˾�ҳ��P��cA��-���\���Ҫ�Sm���kپ�)�����z�g ��|)��`7�G�E���Q�PX�{�U��I���5�5f�;��7쾾�ؾ�|׾�-�8������Y3�G�G���T��@X�6�R�2G�T�8���*��Q�?���5�~���Gܾ�þW���`���΃��a�������w����Ⱦ8������	�'F��!�X�-��2<�� J�O�T�NX��R���C��9.����*�~���־]۾S�򾧁�x�#�a�:�3�L���V�|VW�OtO���B��04�N�&��c�]���:�|��Ӿ9����������Г����ڤ�����,�оS��F�����z�s*%�i�2� A��3N���V�~W�7�N�s=�Y&�f���y���ݾx�վ�Jᾘ7�������+�9�A�s^Q��'X�U}U�ǈK�M�=�R�/�a"�6��C�7N������F˾ѳ�$O��Z?���*���Z���Ъ�k���iپ�'�����y�����{)��_7���E�N�Q��X��U�ӍI���5�f�+���7��ؾ�|׾).龍��H��Z3�ۯG�5�T��AX�
�R� 3G�P�8���*�S�t���6�����Iܾ�þ
������X���Đ��ʮ���x��D�Ⱦ��P���g�	��F�l!���-�b3<��!J�%�T�OX��R��C�R;.�x��=,����־`۾3�������#�h�:� M���V�'WW��tO�3�B��14��&��d�c���;��~��Ӿ<���Ħ�R���ԓ�<���ݤ�c�����о���?���  �  b�*�.�/��1��1�� 1��0��a/��m*�� ��9��|��Ⱦ�'������5��^Sξ��r��{�Wq#���+���/�Y1�1�2#1�F�0���.�W,)�i���}�.���a߾�+žU_��ie��ꬼ���ҾG��Y<	�_��_.%�I�,��N0�S 1�1�h$1��0�[/.�#�'����L���'��>rھĸ��X򳾏3��0���"D׾q�����<=��&�d�-��0�##1��1�>"1��|0�l-�0C&��x���f���Ĵվ����Ⲿ
`���¾�ܾ$��j��:w�9C(��i.���0�+$1�u1��1�l30���,���$����M���\1Ѿ�û��2���굾`ƾ�ᾟ� �D^������)��/���0��!1�.1��1�$�/�ӌ+�D�"�,��(�����@�̾�G��iⱾѷ�
5ʾ�5�8��D����!��*�n�/��1��1��1�t�0�Fa/��l*�>� �����y�K�Ⱦ%����;��sPξ!���p��z�Zp#���+��/��1��1��"1��0���.�,)����<}�����Y_߾�)ž-]��c�������Ҿ���,;	�>��N-%�K�,��M0��1�U1��#1�Q�0��..���'�C����Q'��rھ˸�����3�������D׾�q��}���=���&�'�-���0�$1��1�X#1�~0�Hm-��D&�z�^�>�����վՖ��2岾�b��L�¾�ܾ���!���w��C(�:j.���0��$1��1�T1�$40���,� �$�!�;O���M4Ѿ�ƻ��5�����bƾN��� �E_����K�)�o/���0�~"1��1��1�#�/���+���"��������龯�̾2K���屾tԷ�>8ʾ�8澓��x��˒!��  �  ҴW���V���M�5@�r�1��v$��u�	��4�55��yϾ0w��i񣾤���*ߓ��������������#վ���D��˔��
��N'�x�4��]C�6P�a�W�;�V�F-L�d�9��_"��N��$�%�ھ�U־�徿:�����/���D�I-S��VX�V@T�1iI� e;�7-��U �����+	�d)��ڗ�i%ǾQ���垾B�������g��&��rmľ��ݾ�^�����__����ٴ+��9���G�PS��NX�C:T���F�s2�r��d����o	׾�)پ��������7�tJ�&�U���W�u7Q���D��6�_�(�X�w���;�ھ���׾����ũ����F	��Q���
)�������̾�U����~���-�u#��F0�N�>�8L�^�U�{X�n�P��r@��N*�����7��*�6�վJ޾�X���0���'�;4>�LNO��W��V��M�y4@���1�Qv$�5u�Q��3�R3��wϾ�t����}��tܓ�牙����z����!վ���k����
�WN'�B�4��]C�P�<�W���V��,L�ل9�*_"��M�v"�ܒھ�S־]��s9�k��̄/�p�D�&,S��UX�^?T�QhI�8d;�a6-��T �}���+	��(��`��%Ǿ�P���垾3B�����dh�����Knľ��ݾ `��{��&`����е+��9���G�VQS�'PX��;T���F��2��s�`f���:׾P,پc����j��Y7��tJ���U���W��7Q�C�D�_�6���(��X�9���<����]�׾%��Eȩ�ۻ���������+�����۬̾|W澪���M���.�3#�eG0�'�>�9L�x�U��	X�ܶP�Rt@�7P*�̵�];���-��վ�޾\��X2��'��5>�iOO��  �  ?ɉ������y��N^��6A��r&����Wi���t۾��������������~�>�x��|��Z⊾+���/���}ƾ�����u��,���G�\�d�@�~�v�<n�����jl�K�K�x+�7_���e��������	=��^^�h�{�􈇿撉��g	q�8�T���7�j�&0	�̀�s-Ҿ.ݸ����J���^����z�Z	z��H�������頾FD��X.Ͼ� ��a��;�4�LQ��n��悿�M���&��%�~�P�a���@�d�!���
�'��� � ���a)(�7H��i��恿���m}��������g�o�J���.���� �N5�dVɾ05��i����a���U���y��|�����Mܔ������-��dNؾ����1���#��>�[�`�v��ǅ��ω�q���v�W�:�5������С���*�`��M2�DOS���r�l���ȉ�����H�y�EN^�L6A�Lr&����g��s۾����!�軖�x�� ~�E�x�ez���ߊ��)���_{ƾ5�ᾈ�iu��,�j�G�X�d�@�~�o�'n�����ljl���K�.w+�"^����ɞ�����H���=�i]^� �{�Z���V���Dyq�e�T�"�7�si��/	����,Ҿ�ܸ����lJ���^��J�z�
z�)I��d���l꠾PE���/Ͼ2���E��9�4�+MQ��	n�H炿�N���'����~���a���@���!�x�
����~� ��t*(�H��i�灿����}��ɢ���g���J���.�������6�HXɾT7������ud��vX���y���|�VĆ��ޔ�ٟ��}/��.Pؾ,��������#��>�[�l�v�Aȅ��Љ�8���v��W�-�5������ҥ���,��a��O2��PS��r����  �  �g��<ꦿ|̗�\���CZ��I2��.�>���
Ǿ�慨����趀�>i���Z���V�"]�j�m����e���򮾒�ξ����D���:�q�c��퇿�͛�6�����_ţ��V��Ԋx�D#M�]�*���7�����O<���d��̈�뜿ù��ѫ��Ƣ�+I��	iw�XJL�n&����++ྥ����������5x�9c��VX�X�W��a� bu������������۾���֧"�L�G��|r�� ��-��mU��N���Ȟ�>����i�0P@�`�!���������'���H�P�s����Q7��糫���������sR���h�S�>��d��T���Ӿ���혾�߅��p��s^�w�V��Y��g��7~�}ŏ����PFþ���W��*>.�/�U�����߯������Y������阿҃���Z�Q�4������:��,1�	AV�UO��oʖ�:���Zg���馿 ̗���CZ�I2�G.���N	Ǿ�����۴���i���Z�*�V�x]��m����������\�ξ��������:�w�c��͛�;�����9ţ��V���x�O"M�:�*���T6�N��&N<�6�d��ˈ�iꜿ ���qЫ�nƢ��H��+hw��IL�em&���G*�����������I5x�9c�
WX��W��a�ccu�գ����T�����۾�����"�Q�G��}r�����-��!V������Ȟ��>��S�i��Q@���!�R��b����'�ܽH�9�s�����7�������������~R���h���>�.e��U��b	Ӿ����	ⅾ�p��x^�BW���Y��g�T<~��Ǐ����HþO��,��?.��U�/���o�������bZ����꘿|Ӄ���Z�u�4�"!���-<��.1��BV�'P��(˖�ه���  �  ��ͿS�ƿ,����k��
�u��A�E{��0����_��a��bnf��6P�+�C�DS@�B�E�=DT���l�0ň������Ǿ?����  ���L���}ȝ��㷿�eɿƇͿ,ÿoج��Ȋk���@�Ԗ'���"�,3���V�m������K��L�ʿ�Ϳ������ƍ�Sbc�Ǎ2�B����ܾⱾP���w{���]��K���A�!A�_�I��A[���w�:�����+!׾���6�-���]�)�����������h̿[�˿8���Aأ�������[�$76�2�#��&��=�:f�vō�l穿�
��Ϳ��ʿ^���렿 ,���R��s$��� ���̾ׄ���?��'Bp��uV���F��x@�!�B��YN��kc�^����:���1��b辏g�x�<��eo�6���د��Ŀ�Ϳ�ȿc3���u����|��HM���-�Y"��w+���H���v��I��r���+�ƿH�Ϳ�ƿϞ���k��z�u���A��z��/���s]�����yjf��2P�߽C��N@���E�+@T���l��È������Ǿ�����  ���L�#���ȝ��㷿�eɿ��Ϳÿ.ج�~ˉk���@�~�'�=�"��*3��V�Yl��W���'K����ʿͿv��p��2ƍ��ac��2����ܾ͗f᱾�O��w{�;�]��K���A��!A�k�I�C[�P�w�J�������"׾���$�-��]�����{�������i̿�˿���٣�w�����[��86�ȭ#�F&�=�^f��ō��穿�
��(Ϳ��ʿ^���렿),���R�	t$�� �%�̾d���hA��,Fp�DzV�"�F�\}@���B�a^N�-pc�b⁾�<��h3���ih�W�<��fo��6��ٯ���Ŀ��Ϳ�ȿ[4���v����|��JM���-��"��y+���H���v�{J��3���Їƿ�  �  �����ݿ��ƿ����kJ��{N�S��)���L���ᖾ�tz��>X�1�B�E�6�L�3�u�8�F�}�^���u��Ȟƾ� �%�'�t�Z�����q2����̿�H�a!�}�ٿ����ş�	����&P�y�3��A.��@�ti�nX�����غϿ8����/�׿����y���tu�/�<�c.�P�ݾ�F��"3��gm��O��=���4��c4�}B<�SDM��oi�Y<��9�����׾���[Q7��n�����'���տ�����㿪}ҿG����䔿��n��(D��#/���1���K�F�z�1��������׿��>��٭Ͽ�ޱ��A��_a�c�,�L��b̾'ۡ������b�$�H��9��3�6�b�@��DU���u�����n����꾥�LwH�����9���Zÿ|�ۿVr�Q�߿��ɿ
Ȫ�Mf��%j^���:��[-�s�7�)jY�m�����ʪƿ��ݿ�濁�ݿ@�ƿ<���#J���zN������`K��_���0qz��:X�-�B��6��3�]�8��|F��^����1��֝ƾ@ ��'��Z�Đ���2����̿�H�_!�^�ٿh��^ş������%P��3�E@.���@��i��W��;���Ͽ���R�応�׿����x��tu���<��-�a�ݾ�E���2��cfm���O��=��4�Pd4��C<��EM�Qqi�j=��|���k�׾���LR7��n��������Gտf�俶��{~ҿ����唿D�n��*D�G%/��1�E�K�o�z����宼���׿;��E��խϿ�ޱ��A��3_a���,�����̾�ܡ�����tb�K�H�d�9�{�3�r6���@�(IU���u�񄓾Pp����꾂�0xH���������Zÿ0�ۿ%s�9�߿��ɿɪ�ng��vl^��:�9^-���7�ClY�f�������ƿA�ݿ�  �  25�`�-��`����!�¿���GjU����o�y+�� o��]݀�P�e�q�V�}�R�JY�J�j�:��D��	ľ�%��ʐ(�b�d�1����ο?�y����0��4�*�V���Pￚڹ�j	��ԉs��k��d��(����ֿz��=!�¸1�o;4�>(���dK�-�������@�-P�7�ھ��l�G�v���_�qT���S���]��s�2#������Ծ�
��R:��?}��Z��`��8����%�ϒ3�l�2�A�#���
�x�ܿ���6���ll��p�7���m�����8��t(��<4���1�C@!�Lk��,տLr��}l�LA.��~�Pɾ;o���F��r�m�*�Z�bS���U�ʝc���}�ce��썵�c�����AN��C������2�������+�s�4�{'/�.�+�Ƨʿ�՜���~��i�d�z�⯘���ĿO���&]�*�-��5�%�-�k`�§��إ¿G���iU�j��2n��)��Zm��rۀ�A�e�?�V�C�R�[FY�[�j�m���𝾞ľ�$����(�L�d�1����ο?������0��4�*�6��+P�ڹ����d�s�M k��c��X���I�ֿ�y�+=!�h�1�;4��(�Ү��J�� ��7���@��O�t�ھ<����v���_�wqT�F�S���]�[�s�$���K�Ծ��
��S:�z@}�E[����ῌ���%�0�3�ӽ2���#��
�[�ܿ�����6��Dnl�x�p�뉍����Y�d���(��<4���1�;@!�Dk��,տWr��M}l��A.�1��Qɾ�p���H����m���Z��S�x�U�-�c��}�jg��ۏ��>������BN�UD������x3����5�+���4��'/����+���ʿ�֜�F�~�}�i���z�������Ŀ:����]���-��  �  ��-�0x&�C?��>�;���=��ksQ��^�����������0���ebk�E\��(X���^��bp�FӇ��n���ž����ۡ&�g�_��і���ǿXi���T�;)�j:-�x!#����*�濶���挿�im�lCe��؀�������ο�H�����e*���,�M2!���
��߿聫�l��e�=�tq�uv۾x���x���d|��	e���Y�tY�p8c��y�����"0��͟վ\*
���7��^w��&��i�ٿ�')��#,�G]+�m��<� �Կ�"��}����f�k�j����Y���������:!���,��^*�����6���Ϳ-Λ�+mg��,�"��ʾ�ڣ�����s�	`��VX�aE[��i�W����	��8������;��_�J�6���.���D �;���$��|-��'�������C�ÿJ"���<x���c�.t�e/���>��J���D���&���-��w&�?��>�:��W=���rQ�@^�.��]���"��@���I^k��@\��$X�ğ^��^p�qч�m����ž������&�K�_��і���ǿi���T�);)�m:-�k!#�|��ƅ�0���o匿8hm��Ae��׀�������ο+H�L���e*�3�,�2!���
���߿~������͵=��p��u۾����x��Od|��	e��Y�+ Y��9c�< y��Ꮎ:1���վ+
�r�7��_w�'���ٿZ��)�%$,��]+���j=���Կ�#��[�����f���j�Ő��򴮿�����:!���,��^*�����6���Ϳ;Λ�omg�,��"���ʾFܣ�����!s�}`�![X��I[�<i�x������'������!��E�J���������� 쿍��e�$�`}-���'�,��)���r�ÿ#��e?x�D�c�`0t�z0���?��2��)E��&��  �  �?��&�`��-ٿ:<���6���G�Wp���`þ��G����|�I�l��kh�|ho����������˾k���o"��T�Xe��<���i�
����R���O��*����ο���:w���Q\�3U���m�׆��Fk���\�6"	�\��������t���ɿ����o�Ս6�+�
�߾x��.����L��}<v��j�:wi��Mt�`�������T��ӓھ~b	��=1��Wh��u�� YĿ?�������[��[l��`���l��$�r��aV���Y��$}�:���.~ɿHX����B��]}�		����|#��񥏿�Z�h0'��@���о�_���H�������p���h���k�x�z��늾 ���྾e �00���A�q�~��h��\�ӿx �&���*�rr����޿𼰿�1���e�D T�r9b�Ǉ����4�ؿB���2��?�O&�1���ٿ�;��~6��{�G��o�,�þ
�Gތ���|���l��gh�do� ��	�������˾U����n"�rT�Ye��P���i�����S���O��*���ο.���v���P\��1U�@�m�����j���[��!	������i��tt����ɿ����o�A�6�+�M�߾���Ӝ���L���<v��j��wi��Nt��������U���ھ=c	��>1�}Xh��v���YĿ�����G�3\�~�4m�a���m��׬r��cV�Q�Y�&}�Ь���~ɿ�X�� ��O��`}�	���迀#�����q�Z��0'�8A�Y�о�a���J��F���i�p�m�h���k���z��튾.��~⾾="�1���A�Y�~�qi����ӿmx ����C+��r�v��2޿����2��q�e��T��;b�'ȇ�����ؿ��� 3��  �  L`��:�,pٿ�����d���n���=��	�L���=�Ӿ�?��혞�Ͳ��3Z������`ۆ�骑�����G��Ϝ۾�L��? ��DG��~z��؜�����f�߿%�������Ul�=-ѿ ѭ�o����sb�H�C��=��Q�d�}��������aL����[���i���ο%;������t\�	10�]�.�-�Ⱦu笾����x؊������U��R���r���>M���žp�辥��� ,�Y�V��-���V���&˿x�� ����_���R忹�ſ���Ӂ�|U���>��A���]�'S��5ө�:pͿ��꿤F���D����ÿ����|���TL��	$���!�߾�n���\���C��]����ӂ�;����S��o���^����Ͼ���w���8���g�ξ������տ�#��D��U����ۿ�ٹ�����q��'K�j�<�$QH�%{l��Ғ��ֵ�T_ؿ����_���9��oٿq���od��� n���=�	�������Ӿ�=��Ԗ�������W��[���ن�����o���E��6�۾.L�J? �IDG�z~z��؜�����z�߿0�������2l��,ѿ�Э�𺋿�rb���C���=�t�Q��~}���������K�h��[���h�o�ο�:�������s\�y00����-��Ⱦ笾c���{؊�˶��)V��ڹ��'���"N���ž���a���,�J�V�t.���W��l'˿%��ڍ���`���S忋�ſb񡿗ԁ��}U�Z�>�d�A���]��S���ө��pͿ.���F���D���%�ÿˤ��*|��UL�8
$�a���߾�p��)_�� F��̻��Cւ������U�������`����Ͼ����V����8�m�g�E������S ֿr$�E��6����ۿ�ڹ�׀��H�q��)K���<�CSH�(}l��Ӓ�o׵�`ؿ���  �  ÿO���y���T��������3[�۬:�g� �F�����%rվ�ۻ�Z���N��;՘��E�����>����۾Ć��c(��&��FA�sc��b������籿�࿿��¿����B��A<���4e��H>��L'��#���1�'9R�d��w���ò��j���x�¿�E��]Ҧ��a��u��O�Oe1��^����U龢P̾#����o��k(��神�2���$Z��fɾ���(�����t.�\�K��~p��ڍ�Om������,¿���h۲�YY��^���ֻV��4�*�#�R�%��:��<`�[^��gա��ض��¿����
峿P����ڈ�Եg�>�D� �(��c�9V��߾�þ��Og�������y��i����[��UҾ�m𾥲	��F��7��7W�"O~��s���s��9L��ÿ�K������ړ���t���I���,��G"�K�*��E��o����F���^㻿�ÿ⟽�������R���O3[�;�:��� �x�����pվ�ٻ��W��CL���Ҙ�jC�������z�۾�����'�Q&�FA��rc��b������籿�࿿��¿�����~���;��4e��G>��K'�P #���1��7R����ȋ�����ˬ���¿TE���Ѧ�%a��Cu�N�O��d1�M^����U�MP̾�����o���(��J��������Z��gɾ���Ȕ����{u.�G�K��p�Hۍ��m��Ǖ���-¿У��,ܲ�#Z��+���o�V���4���#���%�L�:��=`��^���ա��ض�¿����峿d���ۈ�/�g���D���(��d�2X��F!߾��þ����i��" ��E|��ܞ���]��9WҾ�o𾎳	��G���7�a8W�P~�t��.t���L���ÿ�L������ۓ���t���I���,��I"�J�*��E�Ȇo����������㻿�  �  ڲ���C���؊��O����j��nW�ͶF��57�~9'���K{��辺y;i���L���f[����ҾC��[������*��:�rBJ��|[���o�Ă��ߌ�8/������S���z��cX�R�6��p��A��8���Pa)���H�P�k�v���@���_��T�����l9y�5	d���Q��A��1��!�\2����mW޾��ƾ�����׸�o�ľED۾����;����
<0�h�?��O���a���v��\��������1D��b@���o�v�L���,�b��v��r>
��
��3�fyT��&w���\���ޅ���э�������q��]�2L��[<��,�����N
����jվ����"巾2i���˾���5����2_%��z5���D�uU��h��&~�Sŉ�f����哿f���^���"d��ZA��l#�
A����-���� ���=��9`��〿ڦ��]���}C��/؊�8O��=�j�@nW�*�F��47��8'���5z�I�%w;���������X��ȦҾ����Z������*�1�:��AJ�2|[�V�o�Ă��ߌ�(/�����~S����z��bX�k�6��o��@�r7�����_)���H��k�����������T�������8y��d��Q���A���1�à!�2�����GW޾��ƾ(����׸���ľ�D۾g����;�J���<0�5�?� �O���a��v�z]��4������D��A��k�o���L�+�,������?
����3�IzT��'w�J����������э������q���]��L��\<��,����P
�0��Rmվ�����緾�k��X˾O��P����`%�Y{5�g�D��uU�ڈh��'~��ŉ������擿&���2����#d��\A��n#��B����
��p� �7�=�;`��䀿m����  �  ?�b�d�h���i��hi�oi�|�i���h�Ncb��UU��A��y*��,�����/�澔�߾���`��0%�d�/���F��X��Qd�.0i��i��Yi�Մi���i���g���`�{R�|>��z&����W���M��*��y�)�������3��
J��B[�ыe�%�i�x�i�8Pi��i�`�i�K1g�h�^�fsO�tF:��"��������R⾴I�1��4�	�v��Ӱ7�@VM�x]���f�ݶi�άi��Li�ٴi��i��Af���\��@L��b6�E������"������e���=���#�͍;��zP�;{_�Swg���i���i�sRi�T�i��hi��'e��yZ���H�Pr2�w�����\5��߾��%�����b�'��U?��rS�Ja�.h�'�i��|i�Y]i�9�i��i�x�c���W��jE��w.�L�����u���u߾õ�� �e���+�C��=V�V�b���h�(�i�5hi��ni���i��h��bb��TU��A��x*�r+�ː��;�澇�߾p��ܓ��#�
�/�i�F���X�Qd��/i���i�9Yi���i���i���g���`��zR��>�z&�9���U���K�r(�}w��������3��	J��A[�ϊe�7�i���i�xOi�b�i���i��0g��^�sO�8F:���"�������S�Jᾶ���	����V�7��VM��x]�e�f���i�íi��Mi���i�G�i�FCf���\��AL�Dd6����$��m%�S��_�⾶���>���#���;�7{P��{_��wg�F�i�&�i��Ri���i��ii��(e�{Z�:�H��s2�����o8��߾���
�������'��V?��sS��Ja��.h���i�K}i�!^i��i��i���c�;X�GlE�*y.��������ky߾7�羏� ��f��+��C��>V��  �  D8��G��nX���k�2퀿P^��7�������d�����eE^���;�	J���������$��8C�f��c���-��/���x`��9����|�~eg�c|T��D�2�4��q$��$�9��� �D�ɾ=庾���P����־c\��VJ�����-�a7=�9�L�4�^�� s�"����E��	����>��{_���Ou���R��n1�����	�p	�l��".�R�N��q����㝑��ޓ�H#��ƅ�Ҍu�Z�`�K�N���>�3Y/�d��?������پ�þ����󹾁�Ǿ��߾�n���-�
�"���2��]B���R�w%e�tz�R��ȱ��'�����������i�P�F��'�2��l�V��1���N8�YXZ���|�����7�������a��V'��tXn��tZ��\I�\�9�8�)�4 �Ua��>�=OѾ����񘷾�5��Q�ξ���q����#(�j8�S�G�.nX���k��쀿^��䅒��������P��'D^�4�;��H�N� ����`�$�37C��f�c���,������`���8���|�eg�|T�sD�М4�Hq$�$������^�ɾ(㺾��������־Z��7I�����-�o6=�Z�L�j�^�, s�Ҕ��{E��Ψ���>��T_��^Ou�\�R��n1����	��	����g".���N�g�q�`���9���ߓ��#���ƅ�ԍu�p�`�t�N���>�}Z/����s@�� ����پ͢þ����"�����Ǿ��߾ep��T.���"�|�2�^B�6�R��%e��tz����;������D������c�i���F���'�����������P8��YZ��|�}���8�����b���'��"Yn��uZ��]I�m�9�o�)����b��A�~RѾٛ��:����8��\�ξ���Nr����$(��  �  "�K<��:]�:���]A��xî�x=��bÿ%"���^��������l��C���)��`"��.���K���w�J���C��󽿾ÿʖ��8Q��*/�� �{�{CU� �5�����[��]�о�%���ɥ�������6��� ���(ž��
� �w���0*��sF���i��� Ġ��ڴ��1�������䵿<{��;���]��=9��>%��+$��"6�<Y�������
泿�������Ⲷ�+7������	Dn�EJ��-����U��5(�d�Ǿ@���M���r��}q��1���õ�1�;�뾙�����e�2��kQ��Pw��������������¿#��r����!��V}�YP�ؐ0��"��(�D@�L�g������ͥ�󃹿��¿�]���ిǛ�N)���Ya�)�?�f�$�o������5ھ.����������ǘ�w����=�����I׾�������J"�kJ<�-:]�����A��2î�%=���ÿ�!��3^���L�l���C��)��^"�.���K��w�:I��+C��p�(ÿN����P���.����{�CU���5�����$����о5$��ȥ������������y&ž���� �����/*�sF�!�i�����à�Yڴ�}1��y����䵿!{��)���]��=9�?%�,$�;#6��Y����C���U泿��N���L����7��r���En�dJ��-��������*�
�Ǿ�B��_P��u���s��53���ŵ���;>�@������2�lQ�LQw�ޥ��5 ��5���¿�#��8����"��	}�(P���0�м"�;(��@���g�$���8Υ�b���8�¿�]���ిIǛ��)���Za���?�Y�$�������8ھ����������ʘ�o��@��%"���׾����n���  �  ���'�?��q��<���鹿�ۿ#2�W�����/�ֿBճ�1����i�zG�P=�y�L�}�t��^���ڻ��{ݿi����!��8��>Կ���"�le�|�6�q���`����;����~}�������p��P3�����j���x�����ȉ�<�%���N��!��4����ſċ�G���������d�˿Dק�Q����[���@��e?�xW�|i���壿W�ǿ��濬�������h�Hɿwg��ez��U6T���)��z
�>R��[þ����ѕ��0��b,���탾�n��⃙�"<��mNʾ��խ��U2��G_��c��b.��u�п������Z��й�ֿ�i&���z���O�Nz=�ƣD�d�d�x��ѯ��ӿX�����/���Fc޿�ͽ������Ow�w�D��e����A�پ���T᡾x␾`p��֪��ϯ��xf��!���Z�����վ���������?�Dq��<��H鹿�ۿ�1�V���𿖜ֿ�Գ�g���i��G�a�<��L���t��]��ڻ�{ݿ���� !����i>ԿE�����e���6����h_����;(����{�������n��삾B1�����[���w����߈�c�%���N�4!��㍢��ſ����������m��J�˿3ק�J����[��@�f?�]xW��i���壿��ǿ�� �����Di�wHɿ�g���z��k7T��)��{
��T�h^þw
��Yԕ�3���.��<����p��΅���=���OʾR��u��{V2�RH_�d���.���п��쿶����[������ֿ�]'����z���O�-|=���D��d��x���ѯ�rӿǝ�?��u����c޿�ͽ�5����Pw�,�D��f������پ���� 䡾C吾:s����������!i������������վV����  �  ˟���J��7��+�����ۿ������;��������Zֿ|���)#���`��(T�<�g�S���� ��ɭ࿿���!���#����Jѿ���S�z�V�>�� �-<�tܼ�Ϧ�������ky��Rk��h�(�q��C���q����oӾ)��{�)��]�+Б�����<��
�u��S�M������ �ƿ	����cz���X�!W�'u�o�����*����׷���������)8����d�\�.���1ؾ�����Җ��΄��bs��1i�Gvj�!@w��+���훾]3�����G9��5s�TU���̿V���
x�*��9�u���忠�������%�k��T�B�]�����8���0ѿ2���{��=����.��Ɯ��O��>�P�J ����O�ɾ�������Ne��^�n�0Yh�Vlm�:,~�-����n��>1žs,�����J��7��򬭿x�ۿ�����V;�A��[���Yֿ����@"����`��&T�%�g�G������Ϭ�L�T���������rJѿ�����z���>�% �;�,ۼ�b���i���Jhy�=Ok�5�h�3�q��A���o��'���ӾI����)�A�]��ϑ�@������
�Z���R�;��o����ƿ����cz��X�3!W�P'u�Bo��H���h���� ����;��}�����8����d�{�.�F���ؾo���lՖ�ф��gs�S6i��zj�CDw�l-��<�︾���l�dH9�A6s��U��&̿����Vx����������忢�������,�k��T��]������8��q1ѿ������?�]����_������WO����P� �݄��i�ɾV���f����g��Ʒn��^h��qm�I1~��⍾ q��)3ž.���  �  6��h�T���������L�����8'���-�c�%�c��W��Z���8J���Sr��d��qz��/��	|ƿ������(�O`-���#��4�5�}���h���OG�2�_�侞W��P����Ӏ�ch��Z��X���`�g�t�c9��r����W;����.�lPk�]X��S�пk����E�*��~,�7: �ٙ	�B�ݿ&@�����8�i�yxg�?���4w����׿6��o ���+��+���e����ֿ�����Hs��4���{�Ҿ�I��쟍�ۋw��[b��X�dZ�Z�e�B~�)В�6$��\y޾�����@�U��&:���⿹j��)"��-���)�e���� ��̿�l���(��d���n�����N��.�鿓:�>$� b-���(�]�)b����Ŀ�_��D&\���#�s��-þ�Ğ�����+o��]�>X���\�D�l���������|N���������T��������OL��e���7'�X�-�!�%�����￀���HI���Qr��d�coz��.���zƿ���R���(��_-�o�#�V4���$����g���NG�v1�-��QV��☕�Ҁ��h�u�Z��{X��`���t�v7������V;�� �.��Ok�X���пI�� ��+�*�z~,�%: �̙	�2�ݿ@�����R�i��xg�_���^w����׿U��� ��+�1�+�������ֿ
����Is��4�����ҾFL��]�����w��`b���X��Z�qf�	~��ђ��%���z޾<����@�����:������j�	*"��-��)�ܐ�Y� ��̿�m���*��d�j�n������O��ن��:�u$�Ib-���(�t�Tb���Ŀ7`���&\���#�0��/þ�ƞ�h���Bo�Q�]�yX���\�+�l�䫄�����WP��d���  �  �q �Y�摓���ſ�������g.�95�*�,����`����¿X���b�x��i�-��������Ϳ���ok���/���4�+�4����ʳ��^牿��J��Z��6�zU����P|�a�b���U��@S� e[���n��s���?���̾:��z/1�ؒp�����Sؿ���Kw"�?2�|�3�l'��.�3�忹���;ߋ�rso�IQm������򬿑�߿�!�%�$��.3�>-3���$�7���޿������x�Y77�y��N�ѾE���^ߊ���q�_�\�S�S�V�T���`�yx����b��O�ݾA��pD��H���߳���뿸-��)�x}4��$1�6����i�ӿ�q�����Zwj�!u��ݒ�����]y��+���4���/�vn����˿�����`�0�%��W���z��~@��������i�K�X�3�R��xW�Ng�jہ�%�������)���p ��Y�����a�ſ��������f.�5���,�q�������¿f���Z�x���i��������ϓͿv���j�?�/�1�4��+�����o���牿�J�4Z�|5�+T��p1|��b���U��<S�Ja[� �n��q���=���	̾a���.1��p�e���Sؿ���-w"�?2�g�3�['��.�#�忳���>ߋ��so�vQm�������Ů߿�!�I�$�/3�k-3��$�n��޿w�����x�s87������Ѿ�����ኾi�q��\��S���T���`��|x�O�������ݾ��D�$I��೿���-��)��}4�D%1�������w�ӿ�r�����eyj�	#u��ޒ�ď��	z�`�J+��4���/��n�3��I�˿ĝ��}�`���%��Y���|���B��󃾞�i�t�X�_�R��}W�'g��݁�6��̍������  �  6��h�T���������L�����8'���-�c�%�c��W��Z���8J���Sr��d��qz��/��	|ƿ������(�O`-���#��4�5�}���h���OG�2�_�侞W��P����Ӏ�ch��Z��X���`�g�t�c9��r����W;����.�lPk�]X��S�пk����E�*��~,�7: �ٙ	�B�ݿ&@�����8�i�yxg�?���4w����׿6��o ���+��+���e����ֿ�����Hs��4���{�Ҿ�I��쟍�ۋw��[b��X�dZ�Z�e�B~�)В�6$��\y޾�����@�U��&:���⿹j��)"��-���)�e���� ��̿�l���(��d���n�����N��.�鿓:�>$� b-���(�]�)b����Ŀ�_��D&\���#�s��-þ�Ğ�����+o��]�>X���\�D�l���������|N���������T��������OL��e���7'�X�-�!�%�����￀���HI���Qr��d�coz��.���zƿ���R���(��_-�o�#�V4���$����g���NG�v1�-��QV��☕�Ҁ��h�u�Z��{X��`���t�v7������V;�� �.��Ok�X���пI�� ��+�*�z~,�%: �̙	�2�ݿ@�����R�i��xg�_���^w����׿U��� ��+�1�+�������ֿ
����Is��4�����ҾFL��]�����w��`b���X��Z�qf�	~��ђ��%���z޾<����@�����:������j�	*"��-��)�ܐ�Y� ��̿�m���*��d�j�n������O��ن��:�u$�Ib-���(�t�Tb���Ŀ7`���&\���#�0��/þ�ƞ�h���Bo�Q�]�yX���\�+�l�䫄�����WP��d���  �  ˟���J��7��+�����ۿ������;��������Zֿ|���)#���`��(T�<�g�S���� ��ɭ࿿���!���#����Jѿ���S�z�V�>�� �-<�tܼ�Ϧ�������ky��Rk��h�(�q��C���q����oӾ)��{�)��]�+Б�����<��
�u��S�M������ �ƿ	����cz���X�!W�'u�o�����*����׷���������)8����d�\�.���1ؾ�����Җ��΄��bs��1i�Gvj�!@w��+���훾]3�����G9��5s�TU���̿V���
x�*��9�u���忠�������%�k��T�B�]�����8���0ѿ2���{��=����.��Ɯ��O��>�P�J ����O�ɾ�������Ne��^�n�0Yh�Vlm�:,~�-����n��>1žs,�����J��7��򬭿x�ۿ�����V;�A��[���Yֿ����@"����`��&T�%�g�G������Ϭ�L�T���������rJѿ�����z���>�% �;�,ۼ�b���i���Jhy�=Ok�5�h�3�q��A���o��'���ӾI����)�A�]��ϑ�@������
�Z���R�;��o����ƿ����cz��X�3!W�P'u�Bo��H���h���� ����;��}�����8����d�{�.�F���ؾo���lՖ�ф��gs�S6i��zj�CDw�l-��<�︾���l�dH9�A6s��U��&̿����Vx����������忢�������,�k��T��]������8��q1ѿ������?�]����_������WO����P� �݄��i�ɾV���f����g��Ʒn��^h��qm�I1~��⍾ q��)3ž.���  �  ���'�?��q��<���鹿�ۿ#2�W�����/�ֿBճ�1����i�zG�P=�y�L�}�t��^���ڻ��{ݿi����!��8��>Կ���"�le�|�6�q���`����;����~}�������p��P3�����j���x�����ȉ�<�%���N��!��4����ſċ�G���������d�˿Dק�Q����[���@��e?�xW�|i���壿W�ǿ��濬�������h�Hɿwg��ez��U6T���)��z
�>R��[þ����ѕ��0��b,���탾�n��⃙�"<��mNʾ��խ��U2��G_��c��b.��u�п������Z��й�ֿ�i&���z���O�Nz=�ƣD�d�d�x��ѯ��ӿX�����/���Fc޿�ͽ������Ow�w�D��e����A�پ���T᡾x␾`p��֪��ϯ��xf��!���Z�����վ���������?�Dq��<��H鹿�ۿ�1�V���𿖜ֿ�Գ�g���i��G�a�<��L���t��]��ڻ�{ݿ���� !����i>ԿE�����e���6����h_����;(����{�������n��삾B1�����[���w����߈�c�%���N�4!��㍢��ſ����������m��J�˿3ק�J����[��@�f?�]xW��i���壿��ǿ�� �����Di�wHɿ�g���z��k7T��)��{
��T�h^þw
��Yԕ�3���.��<����p��΅���=���OʾR��u��{V2�RH_�d���.���п��쿶����[������ֿ�]'����z���O�-|=���D��d��x���ѯ�rӿǝ�?��u����c޿�ͽ�5����Pw�,�D��f������پ���� 䡾C吾:s����������!i������������վV����  �  "�K<��:]�:���]A��xî�x=��bÿ%"���^��������l��C���)��`"��.���K���w�J���C��󽿾ÿʖ��8Q��*/�� �{�{CU� �5�����[��]�о�%���ɥ�������6��� ���(ž��
� �w���0*��sF���i��� Ġ��ڴ��1�������䵿<{��;���]��=9��>%��+$��"6�<Y�������
泿�������Ⲷ�+7������	Dn�EJ��-����U��5(�d�Ǿ@���M���r��}q��1���õ�1�;�뾙�����e�2��kQ��Pw��������������¿#��r����!��V}�YP�ؐ0��"��(�D@�L�g������ͥ�󃹿��¿�]���ిǛ�N)���Ya�)�?�f�$�o������5ھ.����������ǘ�w����=�����I׾�������J"�kJ<�-:]�����A��2î�%=���ÿ�!��3^���L�l���C��)��^"�.���K��w�:I��+C��p�(ÿN����P���.����{�CU���5�����$����о5$��ȥ������������y&ž���� �����/*�sF�!�i�����à�Yڴ�}1��y����䵿!{��)���]��=9�?%�,$�;#6��Y����C���U泿��N���L����7��r���En�dJ��-��������*�
�Ǿ�B��_P��u���s��53���ŵ���;>�@������2�lQ�LQw�ޥ��5 ��5���¿�#��8����"��	}�(P���0�м"�;(��@���g�$���8Υ�b���8�¿�]���ిIǛ��)���Za���?�Y�$�������8ھ����������ʘ�o��@��%"���׾����n���  �  D8��G��nX���k�2퀿P^��7�������d�����eE^���;�	J���������$��8C�f��c���-��/���x`��9����|�~eg�c|T��D�2�4��q$��$�9��� �D�ɾ=庾���P����־c\��VJ�����-�a7=�9�L�4�^�� s�"����E��	����>��{_���Ou���R��n1�����	�p	�l��".�R�N��q����㝑��ޓ�H#��ƅ�Ҍu�Z�`�K�N���>�3Y/�d��?������پ�þ����󹾁�Ǿ��߾�n���-�
�"���2��]B���R�w%e�tz�R��ȱ��'�����������i�P�F��'�2��l�V��1���N8�YXZ���|�����7�������a��V'��tXn��tZ��\I�\�9�8�)�4 �Ua��>�=OѾ����񘷾�5��Q�ξ���q����#(�j8�S�G�.nX���k��쀿^��䅒��������P��'D^�4�;��H�N� ����`�$�37C��f�c���,������`���8���|�eg�|T�sD�М4�Hq$�$������^�ɾ(㺾��������־Z��7I�����-�o6=�Z�L�j�^�, s�Ҕ��{E��Ψ���>��T_��^Ou�\�R��n1����	��	����g".���N�g�q�`���9���ߓ��#���ƅ�ԍu�p�`�t�N���>�}Z/����s@�� ����پ͢þ����"�����Ǿ��߾ep��T.���"�|�2�^B�6�R��%e��tz����;������D������c�i���F���'�����������P8��YZ��|�}���8�����b���'��"Yn��uZ��]I�m�9�o�)����b��A�~RѾٛ��:����8��\�ξ���Nr����$(��  �  ?�b�d�h���i��hi�oi�|�i���h�Ncb��UU��A��y*��,�����/�澔�߾���`��0%�d�/���F��X��Qd�.0i��i��Yi�Մi���i���g���`�{R�|>��z&����W���M��*��y�)�������3��
J��B[�ыe�%�i�x�i�8Pi��i�`�i�K1g�h�^�fsO�tF:��"��������R⾴I�1��4�	�v��Ӱ7�@VM�x]���f�ݶi�άi��Li�ٴi��i��Af���\��@L��b6�E������"������e���=���#�͍;��zP�;{_�Swg���i���i�sRi�T�i��hi��'e��yZ���H�Pr2�w�����\5��߾��%�����b�'��U?��rS�Ja�.h�'�i��|i�Y]i�9�i��i�x�c���W��jE��w.�L�����u���u߾õ�� �e���+�C��=V�V�b���h�(�i�5hi��ni���i��h��bb��TU��A��x*�r+�ː��;�澇�߾p��ܓ��#�
�/�i�F���X�Qd��/i���i�9Yi���i���i���g���`��zR��>�z&�9���U���K�r(�}w��������3��	J��A[�ϊe�7�i���i�xOi�b�i���i��0g��^�sO�8F:���"�������S�Jᾶ���	����V�7��VM��x]�e�f���i�íi��Mi���i�G�i�FCf���\��AL�Dd6����$��m%�S��_�⾶���>���#���;�7{P��{_��wg�F�i�&�i��Ri���i��ii��(e�{Z�:�H��s2�����o8��߾���
�������'��V?��sS��Ja��.h���i�K}i�!^i��i��i���c�;X�GlE�*y.��������ky߾7�羏� ��f��+��C��>V��  �  ڲ���C���؊��O����j��nW�ͶF��57�~9'���K{��辺y;i���L���f[����ҾC��[������*��:�rBJ��|[���o�Ă��ߌ�8/������S���z��cX�R�6��p��A��8���Pa)���H�P�k�v���@���_��T�����l9y�5	d���Q��A��1��!�\2����mW޾��ƾ�����׸�o�ľED۾����;����
<0�h�?��O���a���v��\��������1D��b@���o�v�L���,�b��v��r>
��
��3�fyT��&w���\���ޅ���э�������q��]�2L��[<��,�����N
����jվ����"巾2i���˾���5����2_%��z5���D�uU��h��&~�Sŉ�f����哿f���^���"d��ZA��l#�
A����-���� ���=��9`��〿ڦ��]���}C��/؊�8O��=�j�@nW�*�F��47��8'���5z�I�%w;���������X��ȦҾ����Z������*�1�:��AJ�2|[�V�o�Ă��ߌ�(/�����~S����z��bX�k�6��o��@�r7�����_)���H��k�����������T�������8y��d��Q���A���1�à!�2�����GW޾��ƾ(����׸���ľ�D۾g����;�J���<0�5�?� �O���a��v�z]��4������D��A��k�o���L�+�,������?
����3�IzT��'w�J����������э������q���]��L��\<��,����P
�0��Rmվ�����緾�k��X˾O��P����`%�Y{5�g�D��uU�ڈh��'~��ŉ������擿&���2����#d��\A��n#��B����
��p� �7�=�;`��䀿m����  �  ÿO���y���T��������3[�۬:�g� �F�����%rվ�ۻ�Z���N��;՘��E�����>����۾Ć��c(��&��FA�sc��b������籿�࿿��¿����B��A<���4e��H>��L'��#���1�'9R�d��w���ò��j���x�¿�E��]Ҧ��a��u��O�Oe1��^����U龢P̾#����o��k(��神�2���$Z��fɾ���(�����t.�\�K��~p��ڍ�Om������,¿���h۲�YY��^���ֻV��4�*�#�R�%��:��<`�[^��gա��ض��¿����
峿P����ڈ�Եg�>�D� �(��c�9V��߾�þ��Og�������y��i����[��UҾ�m𾥲	��F��7��7W�"O~��s���s��9L��ÿ�K������ړ���t���I���,��G"�K�*��E��o����F���^㻿�ÿ⟽�������R���O3[�;�:��� �x�����pվ�ٻ��W��CL���Ҙ�jC�������z�۾�����'�Q&�FA��rc��b������籿�࿿��¿�����~���;��4e��G>��K'�P #���1��7R����ȋ�����ˬ���¿TE���Ѧ�%a��Cu�N�O��d1�M^����U�MP̾�����o���(��J��������Z��gɾ���Ȕ����{u.�G�K��p�Hۍ��m��Ǖ���-¿У��,ܲ�#Z��+���o�V���4���#���%�L�:��=`��^���ա��ض�¿����峿d���ۈ�/�g���D���(��d�2X��F!߾��þ����i��" ��E|��ܞ���]��9WҾ�o𾎳	��G���7�a8W�P~�t��.t���L���ÿ�L������ۓ���t���I���,��I"�J�*��E�Ȇo����������㻿�  �  L`��:�,pٿ�����d���n���=��	�L���=�Ӿ�?��혞�Ͳ��3Z������`ۆ�骑�����G��Ϝ۾�L��? ��DG��~z��؜�����f�߿%�������Ul�=-ѿ ѭ�o����sb�H�C��=��Q�d�}��������aL����[���i���ο%;������t\�	10�]�.�-�Ⱦu笾����x؊������U��R���r���>M���žp�辥��� ,�Y�V��-���V���&˿x�� ����_���R忹�ſ���Ӂ�|U���>��A���]�'S��5ө�:pͿ��꿤F���D����ÿ����|���TL��	$���!�߾�n���\���C��]����ӂ�;����S��o���^����Ͼ���w���8���g�ξ������տ�#��D��U����ۿ�ٹ�����q��'K�j�<�$QH�%{l��Ғ��ֵ�T_ؿ����_���9��oٿq���od��� n���=�	�������Ӿ�=��Ԗ�������W��[���ن�����o���E��6�۾.L�J? �IDG�z~z��؜�����z�߿0�������2l��,ѿ�Э�𺋿�rb���C���=�t�Q��~}���������K�h��[���h�o�ο�:�������s\�y00����-��Ⱦ笾c���{؊�˶��)V��ڹ��'���"N���ž���a���,�J�V�t.���W��l'˿%��ڍ���`���S忋�ſb񡿗ԁ��}U�Z�>�d�A���]��S���ө��pͿ.���F���D���%�ÿˤ��*|��UL�8
$�a���߾�p��)_�� F��̻��Cւ������U�������`����Ͼ����V����8�m�g�E������S ֿr$�E��6����ۿ�ڹ�׀��H�q��)K���<�CSH�(}l��Ӓ�o׵�`ؿ���  �  �?��&�`��-ٿ:<���6���G�Wp���`þ��G����|�I�l��kh�|ho����������˾k���o"��T�Xe��<���i�
����R���O��*����ο���:w���Q\�3U���m�׆��Fk���\�6"	�\��������t���ɿ����o�Ս6�+�
�߾x��.����L��}<v��j�:wi��Mt�`�������T��ӓھ~b	��=1��Wh��u�� YĿ?�������[��[l��`���l��$�r��aV���Y��$}�:���.~ɿHX����B��]}�		����|#��񥏿�Z�h0'��@���о�_���H�������p���h���k�x�z��늾 ���྾e �00���A�q�~��h��\�ӿx �&���*�rr����޿𼰿�1���e�D T�r9b�Ǉ����4�ؿB���2��?�O&�1���ٿ�;��~6��{�G��o�,�þ
�Gތ���|���l��gh�do� ��	�������˾U����n"�rT�Ye��P���i�����S���O��*���ο.���v���P\��1U�@�m�����j���[��!	������i��tt����ɿ����o�A�6�+�M�߾���Ӝ���L���<v��j��wi��Nt��������U���ھ=c	��>1�}Xh��v���YĿ�����G�3\�~�4m�a���m��׬r��cV�Q�Y�&}�Ь���~ɿ�X�� ��O��`}�	���迀#�����q�Z��0'�8A�Y�о�a���J��F���i�p�m�h���k���z��튾.��~⾾="�1���A�Y�~�qi����ӿmx ����C+��r�v��2޿����2��q�e��T��;b�'ȇ�����ؿ��� 3��  �  ��-�0x&�C?��>�;���=��ksQ��^�����������0���ebk�E\��(X���^��bp�FӇ��n���ž����ۡ&�g�_��і���ǿXi���T�;)�j:-�x!#����*�濶���挿�im�lCe��؀�������ο�H�����e*���,�M2!���
��߿聫�l��e�=�tq�uv۾x���x���d|��	e���Y�tY�p8c��y�����"0��͟վ\*
���7��^w��&��i�ٿ�')��#,�G]+�m��<� �Կ�"��}����f�k�j����Y���������:!���,��^*�����6���Ϳ-Λ�+mg��,�"��ʾ�ڣ�����s�	`��VX�aE[��i�W����	��8������;��_�J�6���.���D �;���$��|-��'�������C�ÿJ"���<x���c�.t�e/���>��J���D���&���-��w&�?��>�:��W=���rQ�@^�.��]���"��@���I^k��@\��$X�ğ^��^p�qч�m����ž������&�K�_��і���ǿi���T�);)�m:-�k!#�|��ƅ�0���o匿8hm��Ae��׀�������ο+H�L���e*�3�,�2!���
���߿~������͵=��p��u۾����x��Od|��	e��Y�+ Y��9c�< y��Ꮎ:1���վ+
�r�7��_w�'���ٿZ��)�%$,��]+���j=���Կ�#��[�����f���j�Ő��򴮿�����:!���,��^*�����6���Ϳ;Λ�omg�,��"���ʾFܣ�����!s�}`�![X��I[�<i�x������'������!��E�J���������� 쿍��e�$�`}-���'�,��)���r�ÿ#��e?x�D�c�`0t�z0���?��2��)E��&��  �  �m��.�w�J�Y�Nd0�g������N��ʂE����߾Ż��`z��d5��'z��u���|��D��׫����_��O��A"T���q�Ͽ����:��a�[|�{&��^�r��Q��&��a����������a��U����ݿ�����>� ie�t�}�)̀���o�*�L�j�!��M�@���u���1�����ξ�֨�a���X���v�@Hv��=��M���C����ɾ*� ��+�v�l�ڥ�-�� ��.H��ll��P��e�v�h��tC���3快���n������s>���T��H"��L�ݑo��̀���}�ze�/�>��\�`�׿����[�8� �Y�Z���y����m�~��Vu���x��ф����꯾��پYY���>�A��	���C� �O�+�φU��Ou��[���z���]��<5���
�1Tп�!��S��N����ʿX���o0��Y��w��m����w��Y�%d0��f�V����N���E�J��n�߾󹳾jx��Q3���z�iu���|��B�������﻾��ғ��!T�
��~�Ͽ���:�%�a�o|�~&��R�r��Q���&�!a��g������`������1�ݿa��&�>��he��}��̀���o��L�+�!�9M�?��E�u��1�����ξ�֨�1���X��d�v��Hv�7>�����0���4�ɾ�� ���+�Y�l��ڥ����O��f.H�[ml�Q���e���h�(uC����忎����n��_���,?���U���"�A�L���o��̀���}�ze�%�>��\�l�׿��@�[��� ��Z�\���{�����~�G[u�Q�x� Ԅ����,쯾��پNZ��>��A�������� ���+�'�U�cPu��[��Kz���]�5=5�!�
�qUп#��OT��|����ʿݚ�p0�J�Y�a�w��  �  ��w�a6m�V�P��@)�� �a
���^��NC���c⾻�c����&K����{����(������J���]&��CQ������)ɿ*D	��l2��$X�Pq�?w��@h��eH��7 �BB�b���<w��@u��	����Eֿ�T�J�6��[��s�"�v��^e��+D��g����R���q�O�0��W��Ѿ:2��D#��_���r}���|�����N���ҡ̾��p�*��h��t��:�߿?��;�?��Vb��u��|t��'_��m;����ݿI����t���u��܉��������(D��ke���v�� s�o�[���6�C����пe����X�=$ �f���`Vþ�颾Ib�����'�{� ]�O2������.��/Qܾ�w���<�v���GO�������$��L�z�j��w�po��lT�A�-�<���sɿ�{���s��Zy���ÿ���W)���P�)Em�Q�w�%6m�%�P�~@)�� �
���^��dMC�U�����ﶾg�ꗉ��H����{�轁�����������\�:&��CQ�z����)ɿ9D	� m2�%X�.Pq�?w��@h�beH�s7 ��A󿻉���v��wt��9����Dֿ T���6���[�ts�Ύv�t^e�h+D��g�B��􄧿sq�Њ0��W���Ѿ�1��#��_���lr}�f�|�l���	�����̾���5�*���h�au����߿�����?�Wb�P�u�}t��'_�&n;����ݿ+���}u��iv������/��B���(D��ke���v�� s�g�[���6�A����п����c�X��$ �����5Xþ�뢾xd��M�����{��a��4��F����0��,Sܾ�x���<���O��b�����$�v�L���j�[�w��po�rmT���-����7uɿ}��u���z���ÿr��qX)�I�P��Em��  �  (�Y��XP��7����'��*~���>�6����*¾�g���z�����Bć����"���֟��D�ɾ����k���J��Ї��䷿k�������1>���S��Y��)L�߸0��:� kڿ�(����������U���џ��;�����!��aA�yU��rX���I�P-�Y[
���ѿO]��gf�O.�����p۾ ���u��S���Έ�Hj��� ��]���e��g�־%{�nG)��_��4��,˿v��_)���F�M�W���V��QD��%�d���yǿ. ��h������Aޣ��ӿ�W
��-���I���X��[U��CA���!�����%���o��XQ�C��?��_�;�i��������ㇾډ�5��������k���k�P7��9��u�A9���߿�1�g;4�4FN��bY�p[R�[;�E���+￡�������>���3��R���s�6�q�7�*}P�߂Y�mXP�ܪ7����'�4�)~�J�>�r�߼�G¾�e���x��Ё�������������ם����ɾ^��k�8�J��Ї��䷿��������1>���S��Y��)L���0�z:�xjڿ!(��չ��؊���������q���_�!�oaA��xU�prX�W�I�-�[
�)�ѿ�\��wff��N.����mp۾Ø���t��S��ψ��j��2!���]���f����־�{�1H)�h_�u5���,˿Tv�$`)�!�F���W�!�V�-RD�Y�%�Ԭ��zǿ
!���h��S ���ޣ��ӿ�W
�$-���I��X��[U��CA���!�����%��#p���XQ�������M�;�k�����i���凾u܉�� ��4����m���m�D8��9��u��9����߿2��;4��FN�cY��[R��;�����,�է������k���U��e���r迪�׻7��}P��  �  �0��)�+?�����o�ſ������n��X=�W�������3پn���k������<���$랾�u��%@¾���$���� �w�F�<N|�v����	ѿ���6���+���/��%�R��F�T@���9���u�%�m����y
��՞ӿl���?��,��H/�s�#�x5�-�{�������\�t(0��6����Y�ξ���ꣾ������������ʲ�Hg˾�0�u?��,�C�V�j������<�h�*�!�;�.���-�b�����
mٿs���ч�ko�� s��ߍ��1��iE��;�#��G/���,������ӴֿD;������L�xX$�ٝ�����/žOv������ޙ��<�������.�վ���bt���8��h��;��N���	��٢��~'���/�w*��Y�j���Kȿ΃��^���Kl�w�|����Q�¿�\������)��0��)��>�m���"�ſ\����n��W=���������1پJ���"���&��ѵ���螾@s���=¾���N��R� ���F��M|�i����	ѿ&���6���+���/��%��Q�NF��?��:9����u���m����	���ӿ���?���,�JH/�*�#�65�����A���\��'0�@6������ξ����ꣾ���ၚ�����=˲�0h˾2�@��,��V���� ��U=�gh���!���.�`�-�Ɉ�����mٿL����ч�
o�3"s�����Y2���E�H�X�#��G/���,�������ֿe;��殁��L�=Y$�Ğ���02ž�x��G��ᙾJ?��u��<��Q�վ���Su���8��h�_<��̌�����)���~'�F�/�xw*�nZ�k���Lȿ򄜿<_��9Nl���|����D�¿�]����=)��  �  ���0����K%ɿ�⧿GK��i�i��'G���+���(V����jɾ?����U���?����;��辯m�ڶ�-h1�-N�|�r����������п�c�v���)�Φ���ݿ������np�m	P��J�o�^�Ap��x���JͿ����	���#����߿�ǽ�ޱ��$���*]�d=���#��������ؾ~�¾��c��F�����վC���O.!�J:��;Y�����o�����S�ۿY��]��������!tѿ���������b�$K��N�ǖk�����䳿|�ٿ3������ۤ�-n�}|Կ���&���Vw�I�Q�EM4��(���s�.aоe������������ƾ��޾���Κ��)���C�`e�Y���k��pXſ����) ��}��F����!�Ŀ�y���U�� �W��I�mU���z���������8��: �����/�����$ɿ�⧿�J��Īi��&G���+���U�����ɾ����S��I=��j�;!�辖l���bg1��N��r�������¹п�c�u���)�������ݿ9�����lp�&P�aJ��^��o��Nw��<JͿ�ￇ	���������߿*ǽ�}����#���)]��c=�r�#�������Ѳؾ��¾J��{c������V�վ�C����.!��J:��<Y�����p��>����ۿ�����\��� ��tѿ؏��a���_�b��	K�d
N��k�����e峿֜ٿq��������>n�|Կ9���K&��Ww� �Q�'N4��)�-�����cо���-�������,�ƾ�޾1���Л��)���C��`e����#l���Xſ/��.* ��}�G����!�Ŀ�z���V��$�W��I�wU�q�z�}��������8�-; ��  �  ��ÿ����j���~��4�����ݽy��e���P�5e:��E#�Q��ш��i��G$ܾ�"澦N���7�;_(��?��U��j�j~�Jӊ�����)��트�3�¿^�¿�������D`���g�\A�Z +�L�&��\5�Q�T�mc���J��&
���m��tĿG��X����/ǐ�r��V�r���^��I�I�2�����J�7��%�޾Ѫݾ���G��T�/0�kG�%�\�J�p��؂��<���:���������Q�ÿB����1���������Y��8�Щ'�ѽ)��>�7b�\����a���5��?¿gÿP������5���(C��Mf��4:l���W�B�^�*���ht�'7�&pܾ�ᾠ`���~�1� ��7��bN��Mc�	rw�3�����������ĳ�S��KĿ�ܼ��r������[+v�`eL���0�CE&�ۍ.�އH�q�9������4b��6�ÿ0��@j��`~��蘕����4�y�Q�e��P�9d:��D#���0������n!ܾ ��K���6��](�q~?�'�U�� j��i~�ӊ�����)��ኸ�#�¿B�¿��������_���g��ZA�(+��&�S[5���T��b���I���	��Gm���Ŀ�ｿpX������Ɛ�#����r�z�^�I�
�2�����J�<��V�޾-�ݾ���%H�VU��0�G�ށ\��p�(ق�!=��9;��W���������ÿ�����2��a�����IY�:8�C�'�,�)�>�*8b�Ϙ��%b��66��8?¿�ÿq�����e���jC���f��;l���W�/B���*�F���u�
:�sܾ��Ac��2��Q� �
�7�tcN��Nc��rw�������������_ų�����Ŀ�ݼ�qs������H-v�ZgL���0�9G&���.���H��q���������b���  �  ������&���P���X��J%��	픿=D��&�����v�îV�"�6����
C��o�p���!�K�=���]��/}�/����{���0��K����=��6u���>��w���[0��������q��:Q��2��Y���
�m���g�9&���B��dc�M�y����;��|J��)Ԕ��2��o���tN��'2��:�������FNl�G�K�'o-�?�0H	�(���!��j*��:H���h�2��o���ٓ��Q�����"/��w����P��K���2����t����f��rF��(�w/��L���	��)�P�.�ܛM��n��U���c��%Y���J��݊��G5�������C���������+����a�W-A��$�Î����O�r|�'�3�>
S�y=s��Y����������6���j��	C�����?#��3���k����{��#\��<� � �e>�_����X�g�8��X�Jx��<�������������P���X���$���씿�C������z�v���V���6�k���A�)n����x�!�ʸ=�o�]�s.}�����{���0������=��u���>��X���30��g����q��9Q��2��X���
�;��Df��&�c�B��cc���홌�;��J���Ӕ� 2�����)N���1�����u���
Nl� �K�o-�B�IH	�V��9"�9k*��:H�w�h�h2�����$ړ��Q�������/��
���UQ��񨓿ᘍ��u���f�7tF���(��0��M�د	�+�Z�.���M��n��U���c��XY���J������5������CD������@��h,�� �a��.A���$�U��(�����}�o�3�fS��>s�6Z��{�������O7��3k��qC�����#���3���l��N�{�|%\�\<�Ѥ �:@��`�o�����8��X�YKx��=���  �  �f��z�ٺ��)n��mi��N8��_r����ÿA���)̧�J���+yn�>�F�x�-�|]&��1�gN�c�x��$��P���{��� Ŀ;���"2����&�����_Ov��.b��,M���6�m�?m
����U�t�ܾ�V龲c�����9,� IC��Y�iWm���r��������㫿񶺿�Yÿ6���S?����O6��P�_��z<��#)��(�;z9��C[��u���`��4=��O�����ÿ���{����V���z���9��K�o��Z[�c�E�V�.����K�P�뾷GݾK߾e���Q��D�3���J�J�_�+t����k���pl7��ڃ���Ŀ(־�?쮿D闿~���R��4�	�&�C�+��C�yi��Č�+F��@�-ÿ�3¿qȷ��>�������';}���h�]T��8>�'���.���X&�Xܾ�X�6(����v�$�̫;��Q�)�f�C�z������m��'i��8��	r���ÿȘ���˧������wn���F�Ԝ-��[&�I�1�ZeN���x��#������֍��sĿȘ������}&��m��Ov�N.b�n,M���6��~�dl
� ��|S�5�ܾ�T龅b�h���8,��GC��Y�uVm�� ����������㫿�����Yÿ���,?�����<6��@�_��z<��#)��(�~z9�CD[�v��a���=������X�ÿi��󰭿W��g{��`:����o�>\[���E���.� �GM���VJݾ�߾����R����3�%�J���_��t�D���������7��U���GĿ�־��쮿ꗿ�~�v�R�M4���&���+�fC�azi�DŌ��F����-ÿ�3¿�ȷ��>����y��<}���h�S^T�U:>��'��������)徱ܾ�[�P+�����Ɋ$���;�"�Q��  �  ��H�%�k�����A���q˿��뿗���v�V���Y�N{��R����;x���S��'I�Y�WЁ�s����ƿ�꿊���p��;�����7sÿ����m!���Gc��.B�ȷ'�5u�����6ݾ4�ž�;��h����x��ȴѾ������f���5���S��y�J����v���Zֿ����`����~���*�׿�˱�8Ŏ��Hi��)M�a�K���d��X��������ӿ���������i����ڿ�)���՘��~�DOW���8�A���
�m�jԾ;��Z��Bb��|�þ�,ھ]���/�%���>�d,_�{s���Y�����N�����>����,�1˿*q��y܄�X]�¦I�'Q��r�y�j;��{�߿����5K�ƈ�;����ο2������SYp�>RL���/�)���b���� �̾���E��=P��>5ʾ��W����*-��H�s�k�M�������.˿=��l���v��U��0Y㿡z������2:x��S��%I�ߖY�eρ�r����ƿK��,��`p�\;��V���rÿ����1!��6Gc�.B�?�'��t�{���*5ݾY�ž�9��I���~v����Ѿ`�����e���5���S��y�강�[v��QZֿ����D�����Y����׿�˱�0Ŏ��Hi��)M���K��d�Y��Ѡ���ӿ��������Թ��Kڿ*��^֘��~�wPW�9�8����k�
��o��lԾ���� ���d����þ�.ھ����/��%�G�>��,_��s���Y��h����Nῒ���+?������1˿r��h݄�1]���I��(Q���r�.�	<���߿���cK�������οh2��T���(Zp�:SL� �/�o��.d�����̾/���2H��CS��!8ʾ���QX����+-��  �  ��?�c+r����P�ȿõ�������)�70��8(�xm��V�����|�����z��yl��y�������˿8 �����"+���/��&�N�A��^㽿N"��:ye��6����x����Ӿ�Ǹ�>7��+䛾���"���e����ƾZ�����?:&���N�i~��_����ٿQ���rk-���.���"���I⿃����G��
�q���o�q@���뫿 ]ܿ(	��� �pH.��J.��� ��	�BU߿h���j5���T�E*�i��A
���ɾ�����ס��M���@������M���[о�󾘻�GA2��u_�H��O���O뿯��X�$���/��Y,�G�S9�P�п�բ�؃�6'm��bw������պ�J���Ј&�g�/�x-+�t��K��;ο�<��R�x�|�D�������0�޾����{���e��9���mt��
���.���۾���n�ů?��*r������ȿ����e��W�)�0��8(�*m�
V�����������z�xl��x��ے���˿�7 �2��k"+�z�/���&��M����㽿"���xe�e�6�����w��%�ӾƸ�s5��>⛾������M���βƾU�����V9&�±N�~�������ٿ,�ˮ�Wk-���.���"���I�|����G��$�q��o��@���뫿6]ܿ,(	�¡ ��H.�K.�)� �N�	��U߿삮��5���T�|*������q�ɾO����ڡ�=P���B��1���}O���]о���M���A2��v_��������������$���/�MZ,����9�L�п�֢�ك�)m��dw�����aֺ��J�6���&���/��-+���
L��;ο =���x�\�D��������޾�����}���h�� ���Cw���������(۾���o��  �  ��A�4���ڮ�>��T�HX9�
OQ�'}Y�{O��6�-�Y����?܎�ʅ��
���M�������/�<�t7S��<Y�N+M�Jz2��;�Ibܿ�p��Z�q��B6�VU�Y��_���΢�L���������������n���ݯ�sо|8��t!"�m�T�GЎ��V��7� ��#��B��V��$X�oH�:+�i�:�пPԡ��>����:����~ʿ.��Ay'�^�E��=W��&W��E��'�5����ǿq���,�[���&���hzԾٲ��Z��^���g?��w��-���n���C?��]�ݾ��	��0��*j�����aտ�O���.�K�J�a�X���T��?����(���Ⱦ�V���7��z���Ug����ݿ.�ɂ2��PM��DY�DS���<�!��H8�մ�z���оG�F��$��Ǿ�C���ޖ�����+����݊��>��ڧ����þ�z��ȫA��3��Wڮ���7�'X9��NQ��|Y��zO��6������(��Aێ�
Ʌ��	��tL�����3����<�7S��<Y��*M�z2�];��aܿ�p����q�GB6��T���証�j̢�PJ���������������l���ۯ��о�6��� "���T��ώ�VV��� ���#���B�jV��$X��nH�:+�i�3�пSԡ��>����[����~ʿH��ay'���E� >W��&W��E��'�r��o�ǿ����N�[��&�=���|Ծ�۲�:]��ґ���A���
��G���^���A����ݾI�	���0��+j����bտ�O���.���J���X�=�T���?���3���ɾ�`���8��j���2h����ݿZ.��2�QM�EY�cS��<�9��|8��մ�͑����G�G��&� �Ǿ0F���ᖾm�����~���uA��D����þ�|����  �  [�F��؈�}��n��<�+��~R�YSn���w��l�^�N��'��'�����~��&���p����̿��p/0��PV�Aop�1vw�ʈi��{J��S"�L�����|~�Ԝ9��^��پ�`���g������(�~���{�����G��_��Εž�`����"���\��Ƙ�LRԿ&���39�]p]��s�)v�W�c��B��l�@�翝)��˕��S��F����࿻����=� �`�u�_u�g�`�Y�=�u��2ܿ�����d��(�op���8ʾ�`���!��^
��k|���}�IG��]1���୾q3Ծ�M��3�&uu�X�����|���LF�(�f���v��=r�y�Y���4�5(�1�ҿ{���@�������(��/*��t~"��yJ��i��yw�_`p�mLV��$0�����ſt�>�M�i���,�.꼾	Ş�#ߋ�&X��lu{������S���.���Ḿ������F�H؈��|��R�� �+��~R�1Sn���w��l��N�2'��&������w�����T����̿z���.0�KPV��np��uw�v�i�|{J�WS"��K��o��s{~�:�9��]���پ8_��:f��͈��}�~��{�����E��]���ž�^����"�3�\�BƘ��QԿ����39�>p]���s��(v�F�c��B��l�:�翠)��ؕ��j��g��������ף=�$�`�9u��u���`���=�����ܿ������d� (��r��q;ʾ
c��$������o|�*�}�^I��J3���⭾5Ծ�N�H�3��uu�����쿸��MF�}�f��v�$>r���Y�(�4��(�H�ҿ����H��험�{)���*���~"�zJ�8�i��yw�{`p��LV��$0���Ռſ����M�M���.�y켾�Ǟ��ዾ�Z���z{�[���1V���0���㸾�徯��  �  �I��鋿�Ŀ�����2��[���x�9i����v���W��.�Uu�Sǿ����u��Zڥ�f�ӿ/3��7�6�_��"{�kE����s��_S�
)��Y���I���΁��^;�I+��׾���r,��ZZx�r�u�����֋���>�¾j���~x#��_�m�����ۿ��[1A��Hg�#�~���o n��^J�]��Jh�齶�3������w����������E���j�b�������j���E�܈�5��ར�oQh��	)��/���cǾ%�������1���&�u��dw��삾ȹ��k���ҜѾ�����4��z�0�������^8$�l�N�Aq������}���c�-e<�ݵ��Vڿy�������O᜿
E���? �i:)�AES���s��E��k#{���_�,�7��N�?�˿I��UZP���F?�uι��O���t���"|��
u�O�z�톾+���䳵����6��
I��鋿�Ŀl����2���[���x�i��Y�v�K�W�K.��t�\ǿ����t��;٥�D�ӿ�2�{�7���_�m"{�9E��:�s�N_S��)��Y��NI��΁�B^;��*�w׾G���퓾M*���Vx���u�����ԋ��_�¾�����w#�T�_����T�ۿ۽�91A��Hg�	�~�哀�^ n��^J�U��Ch�콶�@���������:�������E��j�w�������j� �E������g����Rh��
)�2��QfǾ����-���������u�iw������0���r�ѾP��m�4�� z����������8$���N��q����6	}�u�c��e<�i��Xڿ��������I✿�E��@ ��:)��ES���s��E���#{���_�?�7��N�x�˿TI��[P�{�LA龷й� R��Qw���'|��u�y�z��{��������⾒7��  �  [�F��؈�}��n��<�+��~R�YSn���w��l�^�N��'��'�����~��&���p����̿��p/0��PV�Aop�1vw�ʈi��{J��S"�L�����|~�Ԝ9��^��پ�`���g������(�~���{�����G��_��Εž�`����"���\��Ƙ�LRԿ&���39�]p]��s�)v�W�c��B��l�@�翝)��˕��S��F����࿻����=� �`�u�_u�g�`�Y�=�u��2ܿ�����d��(�op���8ʾ�`���!��^
��k|���}�IG��]1���୾q3Ծ�M��3�&uu�X�����|���LF�(�f���v��=r�y�Y���4�5(�1�ҿ{���@�������(��/*��t~"��yJ��i��yw�_`p�mLV��$0�����ſt�>�M�i���,�.꼾	Ş�#ߋ�&X��lu{������S���.���Ḿ������F�H؈��|��R�� �+��~R�1Sn���w��l��N�2'��&������w�����T����̿z���.0�KPV��np��uw�v�i�|{J�WS"��K��o��s{~�:�9��]���پ8_��:f��͈��}�~��{�����E��]���ž�^����"�3�\�BƘ��QԿ����39�>p]���s��(v�F�c��B��l�:�翠)��ؕ��j��g��������ף=�$�`�9u��u���`���=�����ܿ������d� (��r��q;ʾ
c��$������o|�*�}�^I��J3���⭾5Ծ�N�H�3��uu�����쿸��MF�}�f��v�$>r���Y�(�4��(�H�ҿ����H��험�{)���*���~"�zJ�8�i��yw�{`p��LV��$0���Ռſ����M�M���.�y켾�Ǟ��ዾ�Z���z{�[���1V���0���㸾�徯��  �  ��A�4���ڮ�>��T�HX9�
OQ�'}Y�{O��6�-�Y����?܎�ʅ��
���M�������/�<�t7S��<Y�N+M�Jz2��;�Ibܿ�p��Z�q��B6�VU�Y��_���΢�L���������������n���ݯ�sо|8��t!"�m�T�GЎ��V��7� ��#��B��V��$X�oH�:+�i�:�пPԡ��>����:����~ʿ.��Ay'�^�E��=W��&W��E��'�5����ǿq���,�[���&���hzԾٲ��Z��^���g?��w��-���n���C?��]�ݾ��	��0��*j�����aտ�O���.�K�J�a�X���T��?����(���Ⱦ�V���7��z���Ug����ݿ.�ɂ2��PM��DY�DS���<�!��H8�մ�z���оG�F��$��Ǿ�C���ޖ�����+����݊��>��ڧ����þ�z��ȫA��3��Wڮ���7�'X9��NQ��|Y��zO��6������(��Aێ�
Ʌ��	��tL�����3����<�7S��<Y��*M�z2�];��aܿ�p����q�GB6��T���証�j̢�PJ���������������l���ۯ��о�6��� "���T��ώ�VV��� ���#���B�jV��$X��nH�:+�i�3�пSԡ��>����[����~ʿH��ay'���E� >W��&W��E��'�r��o�ǿ����N�[��&�=���|Ծ�۲�:]��ґ���A���
��G���^���A����ݾI�	���0��+j����bտ�O���.���J���X�=�T���?���3���ɾ�`���8��j���2h����ݿZ.��2�QM�EY�cS��<�9��|8��մ�͑����G�G��&� �Ǿ0F���ᖾm�����~���uA��D����þ�|����  �  ��?�c+r����P�ȿõ�������)�70��8(�xm��V�����|�����z��yl��y�������˿8 �����"+���/��&�N�A��^㽿N"��:ye��6����x����Ӿ�Ǹ�>7��+䛾���"���e����ƾZ�����?:&���N�i~��_����ٿQ���rk-���.���"���I⿃����G��
�q���o�q@���뫿 ]ܿ(	��� �pH.��J.��� ��	�BU߿h���j5���T�E*�i��A
���ɾ�����ס��M���@������M���[о�󾘻�GA2��u_�H��O���O뿯��X�$���/��Y,�G�S9�P�п�բ�؃�6'm��bw������պ�J���Ј&�g�/�x-+�t��K��;ο�<��R�x�|�D�������0�޾����{���e��9���mt��
���.���۾���n�ů?��*r������ȿ����e��W�)�0��8(�*m�
V�����������z�xl��x��ے���˿�7 �2��k"+�z�/���&��M����㽿"���xe�e�6�����w��%�ӾƸ�s5��>⛾������M���βƾU�����V9&�±N�~�������ٿ,�ˮ�Wk-���.���"���I�|����G��$�q��o��@���뫿6]ܿ,(	�¡ ��H.�K.�)� �N�	��U߿삮��5���T�|*������q�ɾO����ڡ�=P���B��1���}O���]о���M���A2��v_��������������$���/�MZ,����9�L�п�֢�ك�)m��dw�����aֺ��J�6���&���/��-+���
L��;ο =���x�\�D��������޾�����}���h�� ���Cw���������(۾���o��  �  ��H�%�k�����A���q˿��뿗���v�V���Y�N{��R����;x���S��'I�Y�WЁ�s����ƿ�꿊���p��;�����7sÿ����m!���Gc��.B�ȷ'�5u�����6ݾ4�ž�;��h����x��ȴѾ������f���5���S��y�J����v���Zֿ����`����~���*�׿�˱�8Ŏ��Hi��)M�a�K���d��X��������ӿ���������i����ڿ�)���՘��~�DOW���8�A���
�m�jԾ;��Z��Bb��|�þ�,ھ]���/�%���>�d,_�{s���Y�����N�����>����,�1˿*q��y܄�X]�¦I�'Q��r�y�j;��{�߿����5K�ƈ�;����ο2������SYp�>RL���/�)���b���� �̾���E��=P��>5ʾ��W����*-��H�s�k�M�������.˿=��l���v��U��0Y㿡z������2:x��S��%I�ߖY�eρ�r����ƿK��,��`p�\;��V���rÿ����1!��6Gc�.B�?�'��t�{���*5ݾY�ž�9��I���~v����Ѿ`�����e���5���S��y�강�[v��QZֿ����D�����Y����׿�˱�0Ŏ��Hi��)M���K��d�Y��Ѡ���ӿ��������Թ��Kڿ*��^֘��~�wPW�9�8����k�
��o��lԾ���� ���d����þ�.ھ����/��%�G�>��,_��s���Y��h����Nῒ���+?������1˿r��h݄�1]���I��(Q���r�.�	<���߿���cK�������οh2��T���(Zp�:SL� �/�o��.d�����̾/���2H��CS��!8ʾ���QX����+-��  �  �f��z�ٺ��)n��mi��N8��_r����ÿA���)̧�J���+yn�>�F�x�-�|]&��1�gN�c�x��$��P���{��� Ŀ;���"2����&�����_Ov��.b��,M���6�m�?m
����U�t�ܾ�V龲c�����9,� IC��Y�iWm���r��������㫿񶺿�Yÿ6���S?����O6��P�_��z<��#)��(�;z9��C[��u���`��4=��O�����ÿ���{����V���z���9��K�o��Z[�c�E�V�.����K�P�뾷GݾK߾e���Q��D�3���J�J�_�+t����k���pl7��ڃ���Ŀ(־�?쮿D闿~���R��4�	�&�C�+��C�yi��Č�+F��@�-ÿ�3¿qȷ��>�������';}���h�]T��8>�'���.���X&�Xܾ�X�6(����v�$�̫;��Q�)�f�C�z������m��'i��8��	r���ÿȘ���˧������wn���F�Ԝ-��[&�I�1�ZeN���x��#������֍��sĿȘ������}&��m��Ov�N.b�n,M���6��~�dl
� ��|S�5�ܾ�T龅b�h���8,��GC��Y�uVm�� ����������㫿�����Yÿ���,?�����<6��@�_��z<��#)��(�~z9�CD[�v��a���=������X�ÿi��󰭿W��g{��`:����o�>\[���E���.� �GM���VJݾ�߾����R����3�%�J���_��t�D���������7��U���GĿ�־��쮿ꗿ�~�v�R�M4���&���+�fC�azi�DŌ��F����-ÿ�3¿�ȷ��>����y��<}���h�S^T�U:>��'��������)徱ܾ�[�P+�����Ɋ$���;�"�Q��  �  ������&���P���X��J%��	픿=D��&�����v�îV�"�6����
C��o�p���!�K�=���]��/}�/����{���0��K����=��6u���>��w���[0��������q��:Q��2��Y���
�m���g�9&���B��dc�M�y����;��|J��)Ԕ��2��o���tN��'2��:�������FNl�G�K�'o-�?�0H	�(���!��j*��:H���h�2��o���ٓ��Q�����"/��w����P��K���2����t����f��rF��(�w/��L���	��)�P�.�ܛM��n��U���c��%Y���J��݊��G5�������C���������+����a�W-A��$�Î����O�r|�'�3�>
S�y=s��Y����������6���j��	C�����?#��3���k����{��#\��<� � �e>�_����X�g�8��X�Jx��<�������������P���X���$���씿�C������z�v���V���6�k���A�)n����x�!�ʸ=�o�]�s.}�����{���0������=��u���>��X���30��g����q��9Q��2��X���
�;��Df��&�c�B��cc���홌�;��J���Ӕ� 2�����)N���1�����u���
Nl� �K�o-�B�IH	�V��9"�9k*��:H�w�h�h2�����$ړ��Q�������/��
���UQ��񨓿ᘍ��u���f�7tF���(��0��M�د	�+�Z�.���M��n��U���c��XY���J������5������CD������@��h,�� �a��.A���$�U��(�����}�o�3�fS��>s�6Z��{�������O7��3k��qC�����#���3���l��N�{�|%\�\<�Ѥ �:@��`�o�����8��X�YKx��=���  �  ��ÿ����j���~��4�����ݽy��e���P�5e:��E#�Q��ш��i��G$ܾ�"澦N���7�;_(��?��U��j�j~�Jӊ�����)��트�3�¿^�¿�������D`���g�\A�Z +�L�&��\5�Q�T�mc���J��&
���m��tĿG��X����/ǐ�r��V�r���^��I�I�2�����J�7��%�޾Ѫݾ���G��T�/0�kG�%�\�J�p��؂��<���:���������Q�ÿB����1���������Y��8�Щ'�ѽ)��>�7b�\����a���5��?¿gÿP������5���(C��Mf��4:l���W�B�^�*���ht�'7�&pܾ�ᾠ`���~�1� ��7��bN��Mc�	rw�3�����������ĳ�S��KĿ�ܼ��r������[+v�`eL���0�CE&�ۍ.�އH�q�9������4b��6�ÿ0��@j��`~��蘕����4�y�Q�e��P�9d:��D#���0������n!ܾ ��K���6��](�q~?�'�U�� j��i~�ӊ�����)��ኸ�#�¿B�¿��������_���g��ZA�(+��&�S[5���T��b���I���	��Gm���Ŀ�ｿpX������Ɛ�#����r�z�^�I�
�2�����J�<��V�޾-�ݾ���%H�VU��0�G�ށ\��p�(ق�!=��9;��W���������ÿ�����2��a�����IY�:8�C�'�,�)�>�*8b�Ϙ��%b��66��8?¿�ÿq�����e���jC���f��;l���W�/B���*�F���u�
:�sܾ��Ac��2��Q� �
�7�tcN��Nc��rw�������������_ų�����Ŀ�ݼ�qs������H-v�ZgL���0�9G&���.���H��q���������b���  �  ���0����K%ɿ�⧿GK��i�i��'G���+���(V����jɾ?����U���?����;��辯m�ڶ�-h1�-N�|�r����������п�c�v���)�Φ���ݿ������np�m	P��J�o�^�Ap��x���JͿ����	���#����߿�ǽ�ޱ��$���*]�d=���#��������ؾ~�¾��c��F�����վC���O.!�J:��;Y�����o�����S�ۿY��]��������!tѿ���������b�$K��N�ǖk�����䳿|�ٿ3������ۤ�-n�}|Կ���&���Vw�I�Q�EM4��(���s�.aоe������������ƾ��޾���Κ��)���C�`e�Y���k��pXſ����) ��}��F����!�Ŀ�y���U�� �W��I�mU���z���������8��: �����/�����$ɿ�⧿�J��Īi��&G���+���U�����ɾ����S��I=��j�;!�辖l���bg1��N��r�������¹п�c�u���)�������ݿ9�����lp�&P�aJ��^��o��Nw��<JͿ�ￇ	���������߿*ǽ�}����#���)]��c=�r�#�������Ѳؾ��¾J��{c������V�վ�C����.!��J:��<Y�����p��>����ۿ�����\��� ��tѿ؏��a���_�b��	K�d
N��k�����e峿֜ٿq��������>n�|Կ9���K&��Ww� �Q�'N4��)�-�����cо���-�������,�ƾ�޾1���Л��)���C��`e����#l���Xſ/��.* ��}�G����!�Ŀ�z���V��$�W��I�wU�q�z�}��������8�-; ��  �  �0��)�+?�����o�ſ������n��X=�W�������3پn���k������<���$랾�u��%@¾���$���� �w�F�<N|�v����	ѿ���6���+���/��%�R��F�T@���9���u�%�m����y
��՞ӿl���?��,��H/�s�#�x5�-�{�������\�t(0��6����Y�ξ���ꣾ������������ʲ�Hg˾�0�u?��,�C�V�j������<�h�*�!�;�.���-�b�����
mٿs���ч�ko�� s��ߍ��1��iE��;�#��G/���,������ӴֿD;������L�xX$�ٝ�����/žOv������ޙ��<�������.�վ���bt���8��h��;��N���	��٢��~'���/�w*��Y�j���Kȿ΃��^���Kl�w�|����Q�¿�\������)��0��)��>�m���"�ſ\����n��W=���������1پJ���"���&��ѵ���螾@s���=¾���N��R� ���F��M|�i����	ѿ&���6���+���/��%��Q�NF��?��:9����u���m����	���ӿ���?���,�JH/�*�#�65�����A���\��'0�@6������ξ����ꣾ���ၚ�����=˲�0h˾2�@��,��V���� ��U=�gh���!���.�`�-�Ɉ�����mٿL����ч�
o�3"s�����Y2���E�H�X�#��G/���,�������ֿe;��殁��L�=Y$�Ğ���02ž�x��G��ᙾJ?��u��<��Q�վ���Su���8��h�_<��̌�����)���~'�F�/�xw*�nZ�k���Lȿ򄜿<_��9Nl���|����D�¿�]����=)��  �  (�Y��XP��7����'��*~���>�6����*¾�g���z�����Bć����"���֟��D�ɾ����k���J��Ї��䷿k�������1>���S��Y��)L�߸0��:� kڿ�(����������U���џ��;�����!��aA�yU��rX���I�P-�Y[
���ѿO]��gf�O.�����p۾ ���u��S���Έ�Hj��� ��]���e��g�־%{�nG)��_��4��,˿v��_)���F�M�W���V��QD��%�d���yǿ. ��h������Aޣ��ӿ�W
��-���I���X��[U��CA���!�����%���o��XQ�C��?��_�;�i��������ㇾډ�5��������k���k�P7��9��u�A9���߿�1�g;4�4FN��bY�p[R�[;�E���+￡�������>���3��R���s�6�q�7�*}P�߂Y�mXP�ܪ7����'�4�)~�J�>�r�߼�G¾�e���x��Ё�������������ם����ɾ^��k�8�J��Ї��䷿��������1>���S��Y��)L���0�z:�xjڿ!(��չ��؊���������q���_�!�oaA��xU�prX�W�I�-�[
�)�ѿ�\��wff��N.����mp۾Ø���t��S��ψ��j��2!���]���f����־�{�1H)�h_�u5���,˿Tv�$`)�!�F���W�!�V�-RD�Y�%�Ԭ��zǿ
!���h��S ���ޣ��ӿ�W
�$-���I��X��[U��CA���!�����%��#p���XQ�������M�;�k�����i���凾u܉�� ��4����m���m�D8��9��u��9����߿2��;4��FN�cY��[R��;�����,�է������k���U��e���r迪�׻7��}P��  �  ��w�a6m�V�P��@)�� �a
���^��NC���c⾻�c����&K����{����(������J���]&��CQ������)ɿ*D	��l2��$X�Pq�?w��@h��eH��7 �BB�b���<w��@u��	����Eֿ�T�J�6��[��s�"�v��^e��+D��g����R���q�O�0��W��Ѿ:2��D#��_���r}���|�����N���ҡ̾��p�*��h��t��:�߿?��;�?��Vb��u��|t��'_��m;����ݿI����t���u��܉��������(D��ke���v�� s�o�[���6�C����пe����X�=$ �f���`Vþ�颾Ib�����'�{� ]�O2������.��/Qܾ�w���<�v���GO�������$��L�z�j��w�po��lT�A�-�<���sɿ�{���s��Zy���ÿ���W)���P�)Em�Q�w�%6m�%�P�~@)�� �
���^��dMC�U�����ﶾg�ꗉ��H����{�轁�����������\�:&��CQ�z����)ɿ9D	� m2�%X�.Pq�?w��@h�beH�s7 ��A󿻉���v��wt��9����Dֿ T���6���[�ts�Ύv�t^e�h+D��g�B��􄧿sq�Њ0��W���Ѿ�1��#��_���lr}�f�|�l���	�����̾���5�*���h�au����߿�����?�Wb�P�u�}t��'_�&n;����ݿ+���}u��iv������/��B���(D��ke���v�� s�g�[���6�A����п����c�X��$ �����5Xþ�뢾xd��M�����{��a��4��F����0��,Sܾ�x���<���O��b�����$�v�L���j�[�w��po�rmT���-����7uɿ}��u���z���ÿr��qX)�I�P��Em��  �  mv��'&������bh���-�m��.���_m�*�+������;-������B���\ˉ�j`��W���*��A�׾n	��7�,��g�������::�2�u�wo��v���	��E����:���[�7�"�ؖ�W㾿'��Hտ���6A���{�-ݗ��*����ۯ���\���zT��=�+�ؿ����,T�������+���T壾���㊾z��[����~��XǼ���D����L��:��пgh���M��K��.���P����*��{A����o�G����i�ڿۉ����7�e�׍T��:�����7����+��j����{�k�@��/
�����)E���n>����;�ܾ��������[���쉾T���nܕ�p ���0ɾ@���&�r�d�6����S��L'���a��D��{���^��䤥�᷒���n�}�4�GC�s�ʿ�����?ƿ�����.�;9h������!��Fv��&�����|bh���-����~���^m�e�+�̥���;-����}�����(ɉ�@^��F���(����׾Om	���7��+��X�������::�I�u��o��������?����:��b[���"�+�ￖ⾿Y��tտ���H6A�Z�{��ܗ��*��¡�������\��TzT�L=���ؿ���O,T�#����ɴ��#壾��䊾_z��餑�z��Hȼ�����W�L��:���п�h�,�M��K��]��������*���A��>���G�	��N�ڿ�������7�ee��T�
;�����:����+��e����{�i�@��/
����eE��.o>�i�� ݾȅ������]���� ���ޕ��"���2ɾK���&�m�d�����NT�M'�=�a�E��M{���^��'���*���N�n��4��C���ʿʛ���@ƿ/����.��9h������!���  �  >��d��w����^�'�&����k��Lj��y+����#�Ѿ��|�������\����<���)��GC���K۾^v
�]+7�)]|�?���/ ���2�ik�� ��aϟ��£��Ǚ��d���R�j��a}�RT������xMοf��$s9��*q��i������L���ٗ�����D�K�j��<ҿ����@R�������Ͱľ����3▾v���!A��&���N���0�����뾭=���J�[r��F�ɿ����eE��I}�kӕ�����
��s����:w�]�?��K���ӿ�\�������࿭i���K�ˇ��y��DS��?���e��qAq�6�8�wF��l��4���t=�Ѓ�k��З���+���<��S���-Ώ��ؙ�n=���;V����	&���a�$������ �!QX�_4��[{��X��������]�d��-�"���Ŀ����N��������'�T�^����w ����E��^��ɝ^� �&���쿹j��YKj��x+����B�Ѿ��Y����!����:���'��VA��)J۾�u
��*7��\|�-���/ ���2�k���jϟ��£��Ǚ��d��VR�"���|翓S�������Lο����r9�/*q�|i�������L���ٗ������K��i�|<ҿu��J@R������l�ľe���3▾����A��������� �����Z>���J��r����ɿ��fE�@J}��ӕ�����>������V;w�τ?�cL���ӿ�]��ˊ������i�	�K�⇁����IS��=���e��jAq�6�8��F��l��s��2u=����P��癹��-��6?�������Џ��ڙ��?���;a����
&���a������� �qQX��4���{�����Y��������d���-�S#�� �Ŀꕯ�DO������{�'�͗^���� ���  �  �����]r��MD�&����׿�@����c���,�x���޾Ҽ��,g������T��{t���C����þ�,辤���7��Ys��㦿�1�N���O���z�� ��]���-�����h��y9����]ѿ`���zݢ��㻿w���QH$�PT�,e��9���1���,��`�c��4����;��{�����N�����u��RIҾ\u��y�����������������tξ���*��uH�!ˆ��?���\��.���^�ui��&������������Y��~)����������������Gg˿��U4��c�T���A������FMT�?#$�����h�{�;�<�Z���%�LLǾ�^��l���:z��/͛�����Pպ�wھ
����'�4p\��˕�}пʱ��>��rm��W��sԏ��"��q�v�}�I�Q�a��(���a����wm޿=,�9BD��Pr���������*r��MD������׿n@���c�2�,�����޾�����d��Ɠ��]R��0r���A����þ�*����7�(Ys��㦿�1�W���O���z�� ��_���&�����h��y9����j\ѿ�����ܢ��⻿�����G$��OT��d�p9���1���,���c�N4�g�;��-����N����6u���HҾ-u��y��ܐ����5��?����uξ:���֌��uH��ˆ�|@��]�\�.��^��i��W���%��-����Y��~)�����i������S����g˿���4�G�c�T���A������CMT�B#$�&�������{��<�9���'�}NǾ�`��Ҍ���|���ϛ������׺�Ayھ����'�*q\�6̕��п��c�>��rm��W���ԏ�2#����v��I������^�������B����n޿�,��BD�!Qr�����  �  ��g�37^�#VD��J!�z���8����x���a��q4�������yؾ����,���ᜮ��Ҵ�ž�(߾#��|��|=��Hm��I���4ʿ��>o)�,K���a��dg�U�Y�b�<�A����迯���6I��g���<!����Ϳ�@�ք,�$AN�O�c���f�hW�A9�����N�����9aP�/�(�H�K��cϾ�̺�����������N�̾*꾷t	�%��AK��р��ܧ���ݿp���b5��]T�T�e���d��`Q�ݜ0��G��?Կ�Х�����1p��������~�T�8�dW�z�f�#|c��cN�+w-��	�לпL�����s���A��&��b����lǾq ��ˮ�?���`���Pվ�f��}��7`0��?[��Q���&��dd��3�m�@��	\�`�g�FH`��G��5$�.���z7¿d���,Ӎ�t嘿����0��� �:�C�,M^�F�g��6^��UD��J!�(��������x���a��p4�&�������vؾQ�����k���wд� ž�&߾!������=�_Hm��I���4ʿ��Go)�',K���a��dg�D�Y�?�<���������H������y ���Ϳ]@�x�,��@N���c�o�f�W��@9���j���������`P�ϯ(���cϾ�̺�������s��
�̾�*�Fu	��%��BK�hҀ�ݧ�/�ݿ���c5��]T���e���d�KaQ�H�0�H�[@Կtѥ������p��d��G��I~���8��W���f�)|c��cN�/w-�	���п������s�ΚA��'��c���⾕nǾ�"���ͮ�����ʆ��hRվ�h�����0a0��@[��Q��'���d�64�½@�V
\�Ϲg��H`�j�G�6$�R����8¿����Nԍ��昿¼��1��Y ���C��M^��  �  em-��G'��.������п�Щ��U����l���J�2�.�������p��3�ԾE�Ͼ��׾mK�������4�`�Q�9�u�'$��ʞ��t[ڿ��������)���,�c#�*O��������͑��cx�Hsp���"���jҿ������!*�5�,�
�"�2��-��U�¿�����Q��	�`���@�oi&�-��������߾�Ѿ��о#�ݾ���av�.�#�I�=�(�\�с�Ý���5�����^��� �JH,��+�P����n�׿=d��㯈��q���u��������M(����&!��,��*����(4�:_߿>����1���z��ZU�q�7��m��	�\d�r�پ��Ͼ%�Ӿ6���� ��p�G�+��{G�+�h�����4����˿�Q�������%��c-���'���o���ǿd���w���o��~��嘿���y�������L&�m-��G'�p.�������п�Щ�6U����l���J�=�.��������}羛�Ծ��Ͼ:�׾�H�s��l���4���Q���u��#������e[ڿ��������)���,�N#�O�?�近���_͑�Tbx��qp�I��i����ҿ��A��=!*���,�Ŕ"��������¿e����Q����`�c�@�+i&� ��Յ����߾L�Ѿ>�о��ݾt���v���#���=���\�{с�=����6�����I_��� ��H,��+���2��?�׿e��������q��u�W��������(�0���&!�1�,���*����34�^_߿t����1���z��[U���7�o�	�g�(�پ5�ϾƢӾ����� ��q�N�+��|G��h�󒉿���P�˿;R����R�%�!d-��'�0�v���! ǿz����x���o�&�~��昿����N�������L&��  �  ~9��<����ס̿���Ť�F���.�� Uz��d^�/oA� m&����h��1��+K�����,���G���d�����ƌ��z��td���V��;�ѿ���|���.!�����[�Ϳz<���U��#g�jJ�v�D�ydW��/��~������ݿ��e���D￮�ۿA	ſDE�������L��_ׅ�Bq�]�T�]8��q�\)�H� � �;�	������4�q~Q�W,n��m���萿����7����¿Jbٿ����R�����f�¿n��!����Z�&�E��OH���b��%��U����ɿK1�I���������^QԿ�����G��h����&��쐁�T�g��K�C�.��+����X���%����z�#�)E>�_-[��Uw�A���H��������Kʿ���_g�Gy���&�x�׿�����h��u��5Q�(�C���N��op�f��������VԿ�*��8�����㿁�̿�����Ĥ�틖����<Tz��c^�nA��k&�/�� ��.���I�J��k,�F�G�z�d�+��qƌ�4z��<d��~V��&�ѿ���j���!��\���Ϳ<��mU��
g�4J�+�D�"cW�;/��`}��u��9�ݿ���{d��TD�9�ۿ�ſ�D��g����L��(ׅ��Aq��T�38��q�^)�`� �; ���	�)��W�4��~Q��,n��m��+鐿^��8���¿�bٿ���R��
��n��+�¿5�����@�Z���E��PH��b�L&�����+�ɿ�1�;I��������鿇QԿس���G������'��u�����g�I
K�� /�e-���>����������#�LF>�h.[��Vw��������{������ʿH��h�z���'�[�׿�����i��ńu��7Q�$�C�o�N��qp�A���{³�6WԿq+��  �  v;������L�������ô��d��\�ղ�觿Ԝ���́���Z�`$9��$����[|'�ϥ?��Hc�=���`㚿{��K��M��� ��͐���������-��������i���I����|�xYT��4���!�rk��*���D���i�r���󝿣 ���+��
��b����{���8���߶�L<����������᏿�}u��TN�Ȏ0�H? ��^��.�wJ���p������࠿�ۮ�pݵ������g���u��)���q��֦���B���ꟿ�h���n�m�H���,�P �O� �9�1�{NP���w�A��E���V����d���ζ��"��􀴿�̵�]��洿YV�����䈿Լg��C��{)��1���"�`6��gV���~��g��C������=ö�s����崿������g������F7���ՙ��Y���a�`�=�{�&�=����$���:��\�J���{�������:������PL��6���>ô��d��Aղ��秿K���X́�k�Z��"9�s$�J���z'�7�?�CGc������⚿��cK������ ���������������������si��tI���|��XT��4�x�!�<j���*���D�T�i����^� ��T+���������e{���8��S߶�<��p���񾢿�᏿�}u��TN�̎0�a? ��^�<.�fwJ���p����ᠿ#ܮ��ݵ�����h��v��������~���_C���럿�i��|�n��H�D�,����� �i�1��OP���w�������������d���ζ��"��<���S͵�����洿�V��L򜿍刿d�g��C�f})�=3��"��6�iV��~�h���C��e����ö�Ӓ���崿+�������������8���֙�eZ��la�:�=�W�&�����$�E�:���\����"��������  �  񵊿�E�� ����᷿��Ϳ�5俲`��_��n�-�ҿ1౿fH����m�xUM���C�˧R�H%x��(���g���7ٿ��]�������߿��ȿ�s���.��h������I�u��Y�c�<��Z"�W��$�������G��U��z0�¦L�f�i��I��׎�����>��i澿��տf��;���������,ȿ����I���_�`�ׇG��/F���\�ӌ��z�M�ĿZ,����&���Z��U ؿHS��56���K���7��l�����l�"�O��w3����������3� �����R�9��WV���r��������.���Q���Iƿ�ݿZ�H|��]��Sܿ�%��X�����}���U��bD��K��Ji�����X��v>Ͽe���y���~��p濴yп-,��]w��$���.��~�~��-c��6F�/�*�<��ٮ����r������'��C�G�_���{�|���.E��ɧ��M᷿=�ͿT5�X`������쿝�ҿ�߱��G��@�m��SM�6�C��R��#x��'���f���6ٿ��Ȇ��"�񿉈߿n�ȿas��\.���g��{�����u�w�Y���<��Y"�\���������F�uT��y0���L�Pi�AI���֎�����@>��澿f�տ ���:��������俴,ȿ����@���d�`���G��/F��\� ����򢿐�Ŀ�,�u�������ɒ�� ؿ�S���6��`L��&8������l���O�"y3�y����9���q� �����6�9�aXV�n�r�K�������q���]Q���Iƿ�ݿ���|����TTܿj&��4���?�}�u�U�HdD��K�vLi���������>Ͽ���Lz����jp�
zп�,���w�����������~�:/c�8F�ԥ*�������_�������3�'�C�}�_���{��  �  y�n�⿍�򸫿/�ҿ� ��V���'��a-���%��I�Y��5��<���,}�PJo�U���μ���ɿiq���Q��c(�]O-��%�������~ɿEF��K:����f�b�E�I�*��?�> ����Ӿ о�ھV�&
����+9�.W��l|����ȷ��ῧ������.+�%;,�#- ��/
�SE��O��j���t�ՙr����V�����ڿ=_��!�V�+���+����J�3�
��*���^�����Z��><��]"��W� N��x�ܾՀо9	Ҿ��MR������'�I�B���b�����������Ŀ�l�&��q#��-���)�Ʊ�8���LϿtܢ�>ք�b�o�}�y�!�������������#��*-�l,)�ח��C���׿��������Os�XP�,3��������7׾�yϾ]�վ���y����B@0�C�L���n�����������ҿǟ ��V�\�'��a-�n�%��I�����4��f��+}�qHo�_���ػ���ɿ�p��DQ�Hc(�O-�i%�˛������}ɿF��:��#�f���E���*��>�e ����Ӿ��Ͼ؞ھ��%
����*9� -W��k|�(�}ȷ���῁��u���.+�;,�- ��/
�AE��O��l��6�t��r�������-�ڿ^_��!���+���+�������翕
����������8�Z��?<�_"��X��P���ܾ^�о�Ҿ�OT�������'���B�6�b����	���#�Ŀ-m��&��q#��-��)�3������MϿgݢ�-ׄ�0�o�2�y�ꀓ�������=����#��*-��,)�����C�9�׿񟯿���#Ps��P�Z-3�[��w��%��b׾�|Ͼo�վv�������cA0�A�L��  �  ��c�~���B���ǡ���U#��F�:_�+�g�q;]��'B����Hu�"�������񍿏+���ſ�U�zL&��FI�k1a���g���Z�~�>�)�<���P��<N���sX�/g.��J��G����Ӿ���� 5����7ֶ�9�Ⱦ݃����"����C��'w�^��7�ӿ��
�w/�W�O��+d�"if�K�U���6��l��"޿�꫿����?��cƧ��{׿Q��2�G�R��te��^e���R�Hm3�h����ڿ�P��f~�6�H�vF#��'��=辇C˾�R��P��
r��\���a�о �|���*�S�Oe���ɯ����n��(;��hX��g��b�v�L��s*��B���ʿ�e���f��R����&"쿱���j>�l�Z���g��a�ՂI�h'�&��ǿ���Pj���:��I��� ��mݾ��þ�3��Ս�����"���0ھ� ��"/�ׇ6��c�'�����������pU#�kF��9_���g�/;]��'B����yt�5!�����������*���ſUU��K&�/FI��0a�F�g���Z�;�>��(��ￆP���M��'sX��f.��I�+F���Ӿˊ��3���﮾Զ��Ⱦȁ����+����C��&w��]����ӿ��
��v/�7�O��+d�if�9�U���6��l��"޿뫿����?���Ƨ��{׿*Q�>�2�m�R��te�$_e���R��m3�����ڿeQ���~�o�H��G#��(�o@�F˾1U���R��\t������]�о�!�|}�K�*��S��e��'ʯ�
�迨��(;�#iX�g���b��L�Rt*�<C���ʿ�f���g��S������"����j>���Z�Йg��a��I�/h'�&&�ǿ���8 j�	�:��J�	� ��pݾ��þ�6��Ȑ��v������ھ���10�Ĉ6��  �  G�g����y�ۿ
5�x�F��ct�c��g��_4����o�.�A�P���ۿ�P���ӡ��x��:7�����SL�oy�z�����������k�W6<�X=�p6̿N(��2�X��|%�%:��[ؾ�q���ϥ��u�������"��wz���ɾ��� ��5s?�z��3G��L-����&���V�⏀�Z�������u��tIa��o1������ȿ����Kˤ��3ÿ� �� ,��(\�#����h��
R��&}���\�7,��%���۶�R{��KbE����W���̾<ı��a��百՚�D8��ӿ��CԾ�1 �[� ��R����-�Ŀ�g���6�q0f�*��'i�������T}�`�Q���!��𿆥���j��ZU�� |ԿA���*<�L7k�������甋��x��YL��R����㣿Oo��Y4��'�N�徙W¾�>����G��� ��^P���:�� ᾢ�	�+/���g����4�ۿ�4�Z�F��ct��b��L��=4��k�o�ΏA����ۿ�O���ҡ��w�� 6�T��RSL��y�A�������ۘ���k�6<�'=�6̿�'����X�=|%�u9�PZؾIp��)Υ��s������ ��px���ɾ��3��Ur?����F���,����&���V�ҏ��M�������u��gIa��o1������ȿ����bˤ��3ÿ5� �� ,��(\�6����h��"R��@}���\�t,�(&���ܶ��{��|cE����
����̾�Ʊ�d��p陾Xך�f:�������DԾ�2 �� �:R�[����Ŀ�g�
�6��0f�U��Zi������U}��Q���!��𿓦���k��KV���|Կ���A+<��7k�Կ���������x��YL��R����h㣿�Oo��Z4�)����9Z¾[A�����J������R��8=��`ᾤ�	��+/��  �  �n�2���1���)��a��6��5ҝ� ���X�������w[�%�d��wc��e¯�-�ƿ���@�0���g��č��;�����٠��PӅ�|)U�����;߿�雿Q�]�Ll#��w��)�ʾ�᫾����~��E͍��ɓ�~;��KU���;㾠��b�@������1����p<��Lt�����:o���
��������`�H�E���-ݿ�R��<����ֿ����B��:z�B˔��W��O���Ô��Qz�%CB�[/�3�ſ����$yG�7�����N�n��z����뎾�����@��x�ƾ6����^�tV��앿�|ֿ%9���N�����Ϙ�D����o���9��.n�r6�T4�_�˿Ts��!庿�&�Ds�.6U�1̅�5�������/��#č�; h�̺/��f��J���`�w��"4�����ؾ5����1���������琾�]��ڐ����Ӿo��.J.�e�n�亨�����)�b�a��6��!ҝ����X������Ow[�� %�o��ob��O����ƿ/����0�7�g�sč��;���������+Ӆ�?)U�`��6;߿]雿��]��k#��v����ʾ�߫�>���|��Vˍ��Ǔ��9��WS���9㾸����@�&���g1�����I<��Lt�����-o���
��������X�H�B���-ݿ�R��<���ֿ2����B��:z�T˔�X��O���Ô�Rz�aCB��/���ſ����QzG�n��2���ﾾ�p����o���펾�����B��G�ƾ�����_�3V�8핿$}ֿ]9���N�����Ϙ�y����o���9���n��r6��4�u�˿^t��溿s'뿧s��6U�S̅�O�������/��.č�O h��/��f������%�w�{#4���,�ؾ����D4���ő�_���1ꐾ`��;����Ӿi��K.��  �  ��q�5���0����0�9�k��w��F���p��xP��1����d���+������9Ŀ�ʴ��Ϳ����7��r�J���V��-A��□��ҋ�uq^�?=$��濊x���O`�_N#����D�ƾ�ħ����o�������叾G)��D��w�߾"��Y�A��釿��ÿN��d�C�:)�&%��簨��U��v���/���dKQ�3�� �����7u���޿�T���J�p���g����황�Nv��
�����J�ǋ���˿�c����H��O����.㺾(X��^���L��� ������E%��˾¾^��D��X��(��.Uݿ�4�b�W�}ވ�Ѱ���������Ҟ��V~x�>��B�#>ҿi���A���xs���%�a^�U���u���GA��Y���#��?r�7��-��8���l{�	�4�Ch��վ���g(���荾忉����\Y���t���%о����.��q����������0��k��w��2��qp��VP�������d�3�+�ň���8Ŀ�ɴ��Ϳ���(�7�nr����V���@�������ҋ�7q^�
=$����5x��<O`��M#�������ƾ=ç������������㏾R'��B����߾<����A�W釿&�ÿ$��=�C�)�%��ڰ���U��n���(���\KQ�0��#��)���Nu���޿�T���J������g��������gv��%���׌J���D�˿Rd��*�H��P� �復庾�Z���	��UO���"������;'����¾����X�))���Uݿ15���W��ވ��������ݙ������~x��>�uC�<?ҿv���;���\t�P�%�ta^�w�������ZA��Y���#��?r�.7�.�9��jm{��4�Li�'վ����+��z덾��i���[���v���'оޅ�[�.��  �  �n�2���1���)��a��6��5ҝ� ���X�������w[�%�d��wc��e¯�-�ƿ���@�0���g��č��;�����٠��PӅ�|)U�����;߿�雿Q�]�Ll#��w��)�ʾ�᫾����~��E͍��ɓ�~;��KU���;㾠��b�@������1����p<��Lt�����:o���
��������`�H�E���-ݿ�R��<����ֿ����B��:z�B˔��W��O���Ô��Qz�%CB�[/�3�ſ����$yG�7�����N�n��z����뎾�����@��x�ƾ6����^�tV��앿�|ֿ%9���N�����Ϙ�D����o���9��.n�r6�T4�_�˿Ts��!庿�&�Ds�.6U�1̅�5�������/��#č�; h�̺/��f��J���`�w��"4�����ؾ5����1���������琾�]��ڐ����Ӿo��.J.�e�n�亨�����)�b�a��6��!ҝ����X������Ow[�� %�o��ob��O����ƿ/����0�7�g�sč��;���������+Ӆ�?)U�`��6;߿]雿��]��k#��v����ʾ�߫�>���|��Vˍ��Ǔ��9��WS���9㾸����@�&���g1�����I<��Lt�����-o���
��������X�H�B���-ݿ�R��<���ֿ2����B��:z�T˔�X��O���Ô�Rz�aCB��/���ſ����QzG�n��2���ﾾ�p����o���펾�����B��G�ƾ�����_�3V�8핿$}ֿ]9���N�����Ϙ�y����o���9���n��r6��4�u�˿^t��溿s'뿧s��6U�S̅�O�������/��.č�O h��/��f������%�w�{#4���,�ؾ����D4���ő�_���1ꐾ`��;����Ӿi��K.��  �  G�g����y�ۿ
5�x�F��ct�c��g��_4����o�.�A�P���ۿ�P���ӡ��x��:7�����SL�oy�z�����������k�W6<�X=�p6̿N(��2�X��|%�%:��[ؾ�q���ϥ��u�������"��wz���ɾ��� ��5s?�z��3G��L-����&���V�⏀�Z�������u��tIa��o1������ȿ����Kˤ��3ÿ� �� ,��(\�#����h��
R��&}���\�7,��%���۶�R{��KbE����W���̾<ı��a��百՚�D8��ӿ��CԾ�1 �[� ��R����-�Ŀ�g���6�q0f�*��'i�������T}�`�Q���!��𿆥���j��ZU�� |ԿA���*<�L7k�������甋��x��YL��R����㣿Oo��Y4��'�N�徙W¾�>����G��� ��^P���:�� ᾢ�	�+/���g����4�ۿ�4�Z�F��ct��b��L��=4��k�o�ΏA����ۿ�O���ҡ��w�� 6�T��RSL��y�A�������ۘ���k�6<�'=�6̿�'����X�=|%�u9�PZؾIp��)Υ��s������ ��px���ɾ��3��Ur?����F���,����&���V�ҏ��M�������u��gIa��o1������ȿ����bˤ��3ÿ5� �� ,��(\�6����h��"R��@}���\�t,�(&���ܶ��{��|cE����
����̾�Ʊ�d��p陾Xך�f:�������DԾ�2 �� �:R�[����Ŀ�g�
�6��0f�U��Zi������U}��Q���!��𿓦���k��KV���|Կ���A+<��7k�Կ���������x��YL��R����h㣿�Oo��Z4�)����9Z¾[A�����J������R��8=��`ᾤ�	��+/��  �  ��c�~���B���ǡ���U#��F�:_�+�g�q;]��'B����Hu�"�������񍿏+���ſ�U�zL&��FI�k1a���g���Z�~�>�)�<���P��<N���sX�/g.��J��G����Ӿ���� 5����7ֶ�9�Ⱦ݃����"����C��'w�^��7�ӿ��
�w/�W�O��+d�"if�K�U���6��l��"޿�꫿����?��cƧ��{׿Q��2�G�R��te��^e���R�Hm3�h����ڿ�P��f~�6�H�vF#��'��=辇C˾�R��P��
r��\���a�о �|���*�S�Oe���ɯ����n��(;��hX��g��b�v�L��s*��B���ʿ�e���f��R����&"쿱���j>�l�Z���g��a�ՂI�h'�&��ǿ���Pj���:��I��� ��mݾ��þ�3��Ս�����"���0ھ� ��"/�ׇ6��c�'�����������pU#�kF��9_���g�/;]��'B����yt�5!�����������*���ſUU��K&�/FI��0a�F�g���Z�;�>��(��ￆP���M��'sX��f.��I�+F���Ӿˊ��3���﮾Զ��Ⱦȁ����+����C��&w��]����ӿ��
��v/�7�O��+d�if�9�U���6��l��"޿뫿����?���Ƨ��{׿*Q�>�2�m�R��te�$_e���R��m3�����ڿeQ���~�o�H��G#��(�o@�F˾1U���R��\t������]�о�!�|}�K�*��S��e��'ʯ�
�迨��(;�#iX�g���b��L�Rt*�<C���ʿ�f���g��S������"����j>���Z�Йg��a��I�/h'�&&�ǿ���8 j�	�:��J�	� ��pݾ��þ�6��Ȑ��v������ھ���10�Ĉ6��  �  y�n�⿍�򸫿/�ҿ� ��V���'��a-���%��I�Y��5��<���,}�PJo�U���μ���ɿiq���Q��c(�]O-��%�������~ɿEF��K:����f�b�E�I�*��?�> ����Ӿ о�ھV�&
����+9�.W��l|����ȷ��ῧ������.+�%;,�#- ��/
�SE��O��j���t�ՙr����V�����ڿ=_��!�V�+���+����J�3�
��*���^�����Z��><��]"��W� N��x�ܾՀо9	Ҿ��MR������'�I�B���b�����������Ŀ�l�&��q#��-���)�Ʊ�8���LϿtܢ�>ք�b�o�}�y�!�������������#��*-�l,)�ח��C���׿��������Os�XP�,3��������7׾�yϾ]�վ���y����B@0�C�L���n�����������ҿǟ ��V�\�'��a-�n�%��I�����4��f��+}�qHo�_���ػ���ɿ�p��DQ�Hc(�O-�i%�˛������}ɿF��:��#�f���E���*��>�e ����Ӿ��Ͼ؞ھ��%
����*9� -W��k|�(�}ȷ���῁��u���.+�;,�- ��/
�AE��O��l��6�t��r�������-�ڿ^_��!���+���+�������翕
����������8�Z��?<�_"��X��P���ܾ^�о�Ҿ�OT�������'���B�6�b����	���#�Ŀ-m��&��q#��-��)�3������MϿgݢ�-ׄ�0�o�2�y�ꀓ�������=����#��*-��,)�����C�9�׿񟯿���#Ps��P�Z-3�[��w��%��b׾�|Ͼo�վv�������cA0�A�L��  �  񵊿�E�� ����᷿��Ϳ�5俲`��_��n�-�ҿ1౿fH����m�xUM���C�˧R�H%x��(���g���7ٿ��]�������߿��ȿ�s���.��h������I�u��Y�c�<��Z"�W��$�������G��U��z0�¦L�f�i��I��׎�����>��i澿��տf��;���������,ȿ����I���_�`�ׇG��/F���\�ӌ��z�M�ĿZ,����&���Z��U ؿHS��56���K���7��l�����l�"�O��w3����������3� �����R�9��WV���r��������.���Q���Iƿ�ݿZ�H|��]��Sܿ�%��X�����}���U��bD��K��Ji�����X��v>Ͽe���y���~��p濴yп-,��]w��$���.��~�~��-c��6F�/�*�<��ٮ����r������'��C�G�_���{�|���.E��ɧ��M᷿=�ͿT5�X`������쿝�ҿ�߱��G��@�m��SM�6�C��R��#x��'���f���6ٿ��Ȇ��"�񿉈߿n�ȿas��\.���g��{�����u�w�Y���<��Y"�\���������F�uT��y0���L�Pi�AI���֎�����@>��澿f�տ ���:��������俴,ȿ����@���d�`���G��/F��\� ����򢿐�Ŀ�,�u�������ɒ�� ؿ�S���6��`L��&8������l���O�"y3�y����9���q� �����6�9�aXV�n�r�K�������q���]Q���Iƿ�ݿ���|����TTܿj&��4���?�}�u�U�HdD��K�vLi���������>Ͽ���Lz����jp�
zп�,���w�����������~�:/c�8F�ԥ*�������_�������3�'�C�}�_���{��  �  v;������L�������ô��d��\�ղ�觿Ԝ���́���Z�`$9��$����[|'�ϥ?��Hc�=���`㚿{��K��M��� ��͐���������-��������i���I����|�xYT��4���!�rk��*���D���i�r���󝿣 ���+��
��b����{���8���߶�L<����������᏿�}u��TN�Ȏ0�H? ��^��.�wJ���p������࠿�ۮ�pݵ������g���u��)���q��֦���B���ꟿ�h���n�m�H���,�P �O� �9�1�{NP���w�A��E���V����d���ζ��"��􀴿�̵�]��洿YV�����䈿Լg��C��{)��1���"�`6��gV���~��g��C������=ö�s����崿������g������F7���ՙ��Y���a�`�=�{�&�=����$���:��\�J���{�������:������PL��6���>ô��d��Aղ��秿K���X́�k�Z��"9�s$�J���z'�7�?�CGc������⚿��cK������ ���������������������si��tI���|��XT��4�x�!�<j���*���D�T�i����^� ��T+���������e{���8��S߶�<��p���񾢿�᏿�}u��TN�̎0�a? ��^�<.�fwJ���p����ᠿ#ܮ��ݵ�����h��v��������~���_C���럿�i��|�n��H�D�,����� �i�1��OP���w�������������d���ζ��"��<���S͵�����洿�V��L򜿍刿d�g��C�f})�=3��"��6�iV��~�h���C��e����ö�Ӓ���崿+�������������8���֙�eZ��la�:�=�W�&�����$�E�:���\����"��������  �  ~9��<����ס̿���Ť�F���.�� Uz��d^�/oA� m&����h��1��+K�����,���G���d�����ƌ��z��td���V��;�ѿ���|���.!�����[�Ϳz<���U��#g�jJ�v�D�ydW��/��~������ݿ��e���D￮�ۿA	ſDE�������L��_ׅ�Bq�]�T�]8��q�\)�H� � �;�	������4�q~Q�W,n��m���萿����7����¿Jbٿ����R�����f�¿n��!����Z�&�E��OH���b��%��U����ɿK1�I���������^QԿ�����G��h����&��쐁�T�g��K�C�.��+����X���%����z�#�)E>�_-[��Uw�A���H��������Kʿ���_g�Gy���&�x�׿�����h��u��5Q�(�C���N��op�f��������VԿ�*��8�����㿁�̿�����Ĥ�틖����<Tz��c^�nA��k&�/�� ��.���I�J��k,�F�G�z�d�+��qƌ�4z��<d��~V��&�ѿ���j���!��\���Ϳ<��mU��
g�4J�+�D�"cW�;/��`}��u��9�ݿ���{d��TD�9�ۿ�ſ�D��g����L��(ׅ��Aq��T�38��q�^)�`� �; ���	�)��W�4��~Q��,n��m��+鐿^��8���¿�bٿ���R��
��n��+�¿5�����@�Z���E��PH��b�L&�����+�ɿ�1�;I��������鿇QԿس���G������'��u�����g�I
K�� /�e-���>����������#�LF>�h.[��Vw��������{������ʿH��h�z���'�[�׿�����i��ńu��7Q�$�C�o�N��qp�A���{³�6WԿq+��  �  em-��G'��.������п�Щ��U����l���J�2�.�������p��3�ԾE�Ͼ��׾mK�������4�`�Q�9�u�'$��ʞ��t[ڿ��������)���,�c#�*O��������͑��cx�Hsp���"���jҿ������!*�5�,�
�"�2��-��U�¿�����Q��	�`���@�oi&�-��������߾�Ѿ��о#�ݾ���av�.�#�I�=�(�\�с�Ý���5�����^��� �JH,��+�P����n�׿=d��㯈��q���u��������M(����&!��,��*����(4�:_߿>����1���z��ZU�q�7��m��	�\d�r�پ��Ͼ%�Ӿ6���� ��p�G�+��{G�+�h�����4����˿�Q�������%��c-���'���o���ǿd���w���o��~��嘿���y�������L&�m-��G'�p.�������п�Щ�6U����l���J�=�.��������}羛�Ծ��Ͼ:�׾�H�s��l���4���Q���u��#������e[ڿ��������)���,�N#�O�?�近���_͑�Tbx��qp�I��i����ҿ��A��=!*���,�Ŕ"��������¿e����Q����`�c�@�+i&� ��Յ����߾L�Ѿ>�о��ݾt���v���#���=���\�{с�=����6�����I_��� ��H,��+���2��?�׿e��������q��u�W��������(�0���&!�1�,���*����34�^_߿t����1���z��[U���7�o�	�g�(�پ5�ϾƢӾ����� ��q�N�+��|G��h�󒉿���P�˿;R����R�%�!d-��'�0�v���! ǿz����x���o�&�~��昿����N�������L&��  �  ��g�37^�#VD��J!�z���8����x���a��q4�������yؾ����,���ᜮ��Ҵ�ž�(߾#��|��|=��Hm��I���4ʿ��>o)�,K���a��dg�U�Y�b�<�A����迯���6I��g���<!����Ϳ�@�ք,�$AN�O�c���f�hW�A9�����N�����9aP�/�(�H�K��cϾ�̺�����������N�̾*꾷t	�%��AK��р��ܧ���ݿp���b5��]T�T�e���d��`Q�ݜ0��G��?Կ�Х�����1p��������~�T�8�dW�z�f�#|c��cN�+w-��	�לпL�����s���A��&��b����lǾq ��ˮ�?���`���Pվ�f��}��7`0��?[��Q���&��dd��3�m�@��	\�`�g�FH`��G��5$�.���z7¿d���,Ӎ�t嘿����0��� �:�C�,M^�F�g��6^��UD��J!�(��������x���a��p4�&�������vؾQ�����k���wд� ž�&߾!������=�_Hm��I���4ʿ��Go)�',K���a��dg�D�Y�?�<���������H������y ���Ϳ]@�x�,��@N���c�o�f�W��@9���j���������`P�ϯ(���cϾ�̺�������s��
�̾�*�Fu	��%��BK�hҀ�ݧ�/�ݿ���c5��]T���e���d�KaQ�H�0�H�[@Կtѥ������p��d��G��I~���8��W���f�)|c��cN�/w-�	���п������s�ΚA��'��c���⾕nǾ�"���ͮ�����ʆ��hRվ�h�����0a0��@[��Q��'���d�64�½@�V
\�Ϲg��H`�j�G�6$�R����8¿����Nԍ��昿¼��1��Y ���C��M^��  �  �����]r��MD�&����׿�@����c���,�x���޾Ҽ��,g������T��{t���C����þ�,辤���7��Ys��㦿�1�N���O���z�� ��]���-�����h��y9����]ѿ`���zݢ��㻿w���QH$�PT�,e��9���1���,��`�c��4����;��{�����N�����u��RIҾ\u��y�����������������tξ���*��uH�!ˆ��?���\��.���^�ui��&������������Y��~)����������������Gg˿��U4��c�T���A������FMT�?#$�����h�{�;�<�Z���%�LLǾ�^��l���:z��/͛�����Pպ�wھ
����'�4p\��˕�}пʱ��>��rm��W��sԏ��"��q�v�}�I�Q�a��(���a����wm޿=,�9BD��Pr���������*r��MD������׿n@���c�2�,�����޾�����d��Ɠ��]R��0r���A����þ�*����7�(Ys��㦿�1�W���O���z�� ��_���&�����h��y9����j\ѿ�����ܢ��⻿�����G$��OT��d�p9���1���,���c�N4�g�;��-����N����6u���HҾ-u��y��ܐ����5��?����uξ:���֌��uH��ˆ�|@��]�\�.��^��i��W���%��-����Y��~)�����i������S����g˿���4�G�c�T���A������CMT�B#$�&�������{��<�9���'�}NǾ�`��Ҍ���|���ϛ������׺�Ayھ����'�*q\�6̕��п��c�>��rm��W���ԏ�2#����v��I������^�������B����n޿�,��BD�!Qr�����  �  >��d��w����^�'�&����k��Lj��y+����#�Ѿ��|�������\����<���)��GC���K۾^v
�]+7�)]|�?���/ ���2�ik�� ��aϟ��£��Ǚ��d���R�j��a}�RT������xMοf��$s9��*q��i������L���ٗ�����D�K�j��<ҿ����@R�������Ͱľ����3▾v���!A��&���N���0�����뾭=���J�[r��F�ɿ����eE��I}�kӕ�����
��s����:w�]�?��K���ӿ�\�������࿭i���K�ˇ��y��DS��?���e��qAq�6�8�wF��l��4���t=�Ѓ�k��З���+���<��S���-Ώ��ؙ�n=���;V����	&���a�$������ �!QX�_4��[{��X��������]�d��-�"���Ŀ����N��������'�T�^����w ����E��^��ɝ^� �&���쿹j��YKj��x+����B�Ѿ��Y����!����:���'��VA��)J۾�u
��*7��\|�-���/ ���2�k���jϟ��£��Ǚ��d��VR�"���|翓S�������Lο����r9�/*q�|i�������L���ٗ������K��i�|<ҿu��J@R������l�ľe���3▾����A��������� �����Z>���J��r����ɿ��fE�@J}��ӕ�����>������V;w�τ?�cL���ӿ�]��ˊ������i�	�K�⇁����IS��=���e��jAq�6�8��F��l��s��2u=����P��癹��-��6?�������Џ��ڙ��?���;a����
&���a������� �qQX��4���{�����Y��������d���-�S#�� �Ŀꕯ�DO������{�'�͗^���� ���  �  $b���}��A�� ���R���+�ƿ�0��S�A�UW�N��pt��dF�����uە������\���zþ7Mc��P����p�ؿ���@�b��������8���4����0���������]AE�Iz���޿�Dӿ����Z*�mk�и��܄���^���_�������r��/���#<�-�羮���q�;�.��j��Ծ�J���"����k���c�������W�Ͼ�� ���(���h�ty��=5����4��!{�;���\G�����������n��+���Ds���0��D��&տ^�ڿ��	�)2>�ԓ���6��G����_��a��T���������j���&���"�����W��F�Tl���IǾ����_��� ���R��lm���7��V�ݾ�'�.�:��؂�]h��{��K��މ�j���{v��E���L���>��?đ�~�[�P]�9��Laѿ�	����J�S��������Ju���a��t}��'��
����R������ƿ�0����A�vV�h��gr��?D��Y��:ٕ������Z���xþ~K��b�;P�ؿ��\�ؿ���N�b��������@���6����0�����o���AE��y�0�޿Dӿ(����Y*�k����������^���_������ur������<�������D�q�Ӑ.�Hj�nԾwJ���"��K��ʟ��򬞾����J�Ͼn� �^�(�o�h��y���5���4�"{�g����G���������$o��b����s���0�GE�j'տ/�ڿ-�	�{2>������6��V����_��a��P���������j���&���c���Y�W��G�<n���KǾٞ�����B��=U���o��7:���ݾ�(�3�:�ق��h�����RK��މ������v��YE��M��=?���đ� �[��]�}��bѿ�
�t����S�׼�����xu���  �  �n�����!�����EXJ���������7��,:A�>���E���̩�\i��b��zW����Ⱦ�f����O�Y4��նҿs��QjY�֘��t���l3��3���߻��ġ�T���m=�Pi	�h�׿=Ϳ���#�,za�kE��^���ء��)s��)����V���hx�p�4�'���Ъ��ko���.�)��ؾ*﷾P���AV���ܚ�
�� 4��1Ծ����m)��f��룿`��-�ޘp�4�y��>�������v������fi�$�)������ο�-Կ���϶6�vix�B������|������Ϩ���`��za��V ��ۿ�!��/�V��:��e����˾?4��x���9��䚜�Z짾iཾR�b���:�>!��p��������B�b���:��_���Q������㭫�٪��%�R��z�v濭A˿���s.��fK�"ч��|������n�����������XJ�Բ�����:7��`9A�]���C�����ɩ�g����?U���쭾�Ⱦ&e�6��?O�)4����ҿt��]jY�����~���t3��4���߻��ġ�8��6m=��h	���׿q
Ϳ��0�#��ya�:E��0��������r������V��Chx�8�4������Ϫ�]ko���.��(��ؾ�O���pV���ܚ�����4��$Ծ��sn)��f�:죿�`�7�-�/�p�`����o��������v��! ���i���)������ο�.Կ��!�6��ix��B��#����|������̨���`��{a�W �8�ۿ"���V��;��g����˾�6��oz��6<��B�����⽾|�m��	�:��!��󥹿�����B�����:������Q��Ҵ��-���&���šR�9{����B˿γ�/�0gK�^ч�}������  �  *ۯ�GI��2ٓ��o�c�3�r/ �����큿k?B��z�V��3�о�c�����V��� ���ļ� �׾�� ��� zN�y_���
ÿz�
�j@��e|��G��;5��P��������*����a�.(�{.����Ŀ�㻿��ۿ9'�@G�����i����������H������d�Z�,!�P��<����j��1��������2Ǿ�β�L����4��/3��_ľ����x	��-�6)c�0^��&<ۿ@=��@T��߇�ԋ��8K����[���Ą���M�cU�e��Of������C��gL"���Z�u�����_���i���ӛ��x����F���.�ʿ$s���
U�2�#�]��z۾�'��c[��Ѐ��� ���d���M;�U񾀻���<�K{�8ԭ�����J-��fh�����M�������r���Җ��u�ZK:�o��!ѿw_����̿G���4��o�	��ۄ��ۯ�'I��ٓ��o�8�3�H/ �����=큿�>B��y�T���о�a��k���S��a��[¼��׾�� �"�}yN�@_���
ÿw�
�j@��e|��G��A5��P�������*��d�a��(��-����Ŀ㻿��ۿ�&��G�Ȅ��<��|���{���!�������&�Z��!�����;���j���1�j��*���2Ǿ�β�|���65���3���_ľ��㾆y	�{-� *c��^���<ۿ�=�3AT��߇����iK���������*ń�j�M��U�C��%g��K�����￶L"� �Z�������f���i���ӛ��x����F���c�ʿos���U��#�
^��|۾*���]��C���d#���f���O;�W񾌼���<�I{��ԭ�����;K-�gh�������������'Ӗ���u��K:��o�#ѿ�`��ǒ̿���p4�o�A	��	����  �  푍����o��3C�)���8߿J�������J�&�5�U'ﾯ�ӾZ�þ4k���{ƾ��ؾR���My��0-��U��4���{�����#��kM���w�����K�����+�e��h7��
�=ѿ���q��������󿆷"�КQ�D�{������܌�-+���4a�*�3�X+�Jʿ����7�k��:=��#��������I;�!��"}��4`˾������h�8�p�e�������ÿ���I�.��_\�x���T���ċ��}��V�4�'�ǝ��!����ʤ�hF��W:˿0?��*2���`�5K��Q��E׊���{��wR���$�����D��� ���jZ���0��=�7���^�۾��Ǿ���K�¾1�Ѿ)�뾢����"��3F�`�x�Ⅱ�P�׿VI�U>���j��9��g{������@Ls��0G������F鳿cx���j����ݿ���S�A���n�����Ǒ�����o��3C�����8߿񝦿L���J�&�	4�%�V�Ӿ��þ�h��(yƾK�ؾ���Dx�0-�U�l4��Y{�����"��kM���w�����K������e�Lh7�ٯ
��ѿm�������
�����&�"�s�Q��{������܌�	+��u4a���3�#+��ʿq�����k�):=��#�_������I;""���}���`˾B��^�����8�6�e�%���;�ÿ����.�I`\�2x���T���ċ�~���V���'���������{ˤ�*G��;˿|?��*2��`�EK��Y��I׊� �{��wR� $����RD��� ��kZ���0��>������۾,�Ǿ������¾��Ѿ}�뾼����"��4F�X�x�^�����׿�I��>�݊j��9���{��9���Ls�N1G����'��o곿�y���k����ݿZ����A��n�+����  �  �R��J��5������Gſ}۠�U����Fe��D���(�����= ��뾱��ф���v�ү.��qK��`m��ċ��맿|�ο@�3��%�:�l�M�$R�/�E���+��2�Wؿ��������È��}���Z}����5};���N���Q�n�D���+����;�9����.����~�x�Y��:��� ��<�=���$7�'U澳$��G5	�\��5�7�!V��Gz�.��ˈ����޿x�
�2�(��B�Q��O�,D>��:!��J ��+ƿY1���q��3����ѿ���7P(��`C�P�Q�O�o�=�� "��H�K�ӿq����z����q���N���1�~���`�>���%�8��aa��t�� &�<ZA�"[a�!!�������|��r��;���2���H���R���K���5�`F����E���5��q�������8t����俫��L_2�J�I�ƖR��J��5��������ſ"۠�񘆿�Ee�#�D���(�y���< ������2��vu���.��pK��_m��ċ�I맿T�ο6�1��%�:�j�M�R��E���+��2��ؿb���Q���j�4ģ���|������|;�j�N�`�Q�)�D�q�+�p��;�䲷��.��v�~��Y���:�i� ��<�A���T7羅U�@%���5	������7��V�MHz��.��G���D�޿��
���(�v�B�^Q�|�O��D>�a;!�YK ��,ƿ&2������*	��ڄ����ѿ���eP(��`C�e�Q�+O�{�=�� "��H���ӿ¦��{���q���N���1����Vb����(�ߐ��c�����&�H[A�\a��!�����}����ￄ��2���H�+�R�'�K�:�5��F���G��7����Ñ�4u��~�����_2���I��  �  %|��e����5D�LwԿ	)����Ed��gN��;�}��Q[�8a;��!�g����b��&��B���b�����ƒ�\�������¿Z?ڿ����q	�e�����!�
�N���7ʿj~��
烿�}d�0�]�:�t�?y��"ѷ�^��*�����dw����Ï濵X̿�����-��N����,r�P4P�h�1��F����r9��Z��/�Z�L�Xn�?#���֗�v�������ɿWf��Q �Q�dE�H�����Y�ZU��'��g�x��_�Qb�8B�������ſ�q��a	�W��s���
����&=ݿ��Ŀ?\��Q:��{���r��?�f��E�$f)�����T����6���&8��W���y�����Ĝ��g�������ѿ ���ւ�k�����%E �cVؿ ���Ȍ��"m���\���i�{������ܟӿ�o��|���{��e�x���C��vԿ�(������c���M��3�}��P[��_;���!������(a���&��B���b�����2ƒ�흡�Ǒ��͗¿2?ڿ{���q	�[������
���7ʿ�}��}惿�|d���]��t��x��wз�����)�n�Ł�#w����Z��XX̿�������~��!���o,r�&4P�T�1��F�����9��Z�/�ΕL��Xn��#��Tח��v��<��(�ɿ�f�/R �bQ��E�������Y�!V�������x�<_�wRb��B��-�����ſr�b	�W��s���
����a=ݿF�Ŀ�\���:���{��Ns����f���E��g)�Q��TV������(8�*�W���y�����3Ŝ�fh������ѿ� �<�,��˝�$���E �YWؿ���Ɍ��$m���\���i�f���뺪���ӿlp��̹��  �  �ѿ+�տnԿQ�ѿ�ѿ`>Կ��տ�Kѿ�?Ŀ?)������y�3BQ�I�7�ˬ0�<�Y�q��N���c����ǿ��ҿ`�տ�ӿKdѿ"ҿ��Կ6vտ��Ͽe9�����Be��Rr���K�~x5��I1�s�?��e_�~ ���џ�J"��Peʿ��ӿ+�տ{!ӿ�Dѿ�cҿ�տ1տ��Ϳ����즿{����j���F�"x3�1l2��C�<f�$K����4���`�̿<�Կ/Nտ��ҿ"<ѿ �ҿ�fտ�uԿ��˿Z��������䈿��c�|B���1�t4�o�H�Z$m�����R������ο�7տ��Կ�AҿvLѿ�Iӿv�տ��ӿ �ɿ�涿a��9����=]���>� 1��>6���M�͂t�wԒ��u���A¿�Jп�տb�Կ��ѿxsѿ��ӿK�տk�ҿǿU��v������!W���:���0���8��"S�],|�.(���|���4ſ��ѿ��տԿ��ѿ��ѿ
>ԿK�տ)Kѿ�?Ŀ�(��i�����y��@Q���7�3�0�n<��Y�����~��c���ǿ�ҿ�տ��ӿdѿ�ҿ�ԿvտX�Ͽ*9������d��hr�~�K�Yw5��H1�2�?��d_����!џ��!���dʿG�ӿ��տ!ӿBDѿzcҿKտ�տU�Ϳ�����즿g����j���F�;x3�`l2�c�C��f�]K��J��������̿��Կ�Nտy�ҿ�<ѿ��ҿegտUvԿ��˿���T����刿�c���B��1��4���H�i%m�����RS����Q�ο�7տ��Կ�Aҿ�LѿJӿ�տ��ӿ��ɿ�綿�a���S?]�[�>��1�k@6�)�M��t�Ւ�Bv��B¿lKпq�տƋԿ �ѿ�sѿ�ӿ�տ�ҿ�ǿ'��V��淀��W�i�:�]�0�h�8��$S��-|��(���}��E5ſ�  �  23��=���>����տ����L���Y_�o�W��AEѿf���+��kh��]��n��g��-����ڿ�E�Ї������@H�$a�,Rп���\�������Y�����w�\�U�V�6��f��)��� ��m�*��AG�L�h��`��T��	���E���ƿ�޿6���et� ��
�ߑ�{2�	:ÿx���. ��u^a�ļ_��6{�ܘ�T���ȥ远��+X��Ŷ�l�����A�ȿZ ��:���Y��m8��Wml�U�J�5�-�Ip����iF��H�Kz3��R�1t�`܊��Q��G꨿����ǦͿ;(迭��o�s��c���7�aa߿��������Ħr���]���e�H��L�����̿��ū���ъ����"1��S�ؿu������Ϡ��鑿����`��[@�bx%�i���E[�H�"�/=��2]����-���2���󭿴=��2�տ���L����#_�/�{V���Dѿ����H*��fih�]�:�n��f��9,��ӰڿiE�v��W��v�H��`��Qпg��'����������2�w���U�t�6��e��(���Ӷ�>�*�t@G�*�h�D`���S�����@E��gƿ��޿����Bt����	�ˑ�^2��9ÿo���0 ���^a��_��6{�9ܘ����������XX�8�������.��Ћȿ� ��ܦ����9���nl���J���-��q����G��I�S{3��R��t��܊�R���꨿�����Ϳ�(�����Ŕ����K8�9b߿����������r���]�O�e��H��������̿��� ����������|1����ؿ�u������3Р��ꑿŤ����`�P]@�z%�$�����\���"��=��3]�M��S.���  �  �܇�!���9~ǿ���������6�/�K�ъR���H�&�0�ѻ�B��4$������������Ǹ�q￦�}7��eL�	kR�&�G���0���X�쿪;���㛿�삿�n_���?���$��k��������`德��O�()��+3�)�P�x�s��ޏ�v�����ֿ@����#���>���O�=&Q��(B��&����ο�����Q��S��ힿ�ɿ\��#�-�?�DP��P�MA��'�5#	���ۿ��������x�DT�396�/��H8����徏��P��<G�`�!���<���[�Ϗ��A����ֹ��翚��wx-�d�E�f
R���M��:������������9f���s��Ȗ��?����6ۿ
�*q-���F��IR��"M��l9�Y!����|\̿����q��8Pk���I��6-�	B��������뾒
�����Q*�|TF�tCg�܇������}ǿ����u��^�6� �K���R���H���0�y��}��]#��0����
��%����Ƹ�z�/�7�3eL��jR���G�r�0�����c;���㛿\삿n_���?��$��j�(�������^征��wN�(��*3�$�P���s�9ޏ����%�ֿ����#���>�߯O�%&Q��(B��&����ο�����Q��j��.ힿ�ɿx�#�S�?�DDP�K�P�CMA��'�u#	��ۿ����Q���,x�gET��:6�����9�%��9����羌��@H�H�!�w�<�Z�[�#��������ֹ�G�Ҽ��x-���E��
R��M�Z:�����������*g���t���������W7ۿd
�nq-��F��IR�#M�m9�!����\̿	��0r��mQk��I�8-��C�x��G������������R*��UF�yDg��  �  ��?��u�⿾b�"�E�i4q��3������k����l��M?�����zڿ�Ѯ�����Xϵ��V�y;���I��ru�>���#b�������@h��~;���^Կ&��={u�@�C�� ��|��龏kо6^¾�˿�K�Ⱦ�ݾ��������2��.]�p'���?������l '���T��r}�1D��ϲ���r���C^��/����vȿ�B��Ԅ���7ÿ����o`*�CY����������V���+�Y�*,�@���e���V����b���6����Q� ���wʾO7��ހ���Jξ�i�~�t��/h?�Jo��H��-tͿ�h
�n\6��c�����}��}���6�y�~O��2 �7��!㹿52��/諿bԿO��H	:�^�g�����k��w[��uu�%�J��9���꿨���WN��tR��W+�U����b�׾�žxZ���~ľuվ���]|�k�'�hM�����B?��&�⿚b���E�B4q�q3������I��8�l�UM?�-���yڿ�Ю�����Oε�zU��:�+�I�{ru�����a��r����@h��~;�����]Կ����zu���C�d� ��{�`�龸iо?\¾zɿ�1�Ⱦ�ݾ��������2��-]�'��I?��.���C '�p�T��r}�$D��Ĳ���r���C^��/����vȿ�B��넥�8ÿ����`*�3CY��������%��q���e�Y�F*,����f��gW����b�+�6�C���� ���Szʾ�9��5���Mξ�k�g�G���h?� o�DI���tͿ�h
��\6�[�c�������������y��O�V3 �>��"乿+3��髿5Կ����	:���g�3����k���[��2uu�D�J�:��������N��*uR��X+�������T�׾�žr]��܁ľ?վ`�}���'��hM��  �  74���������6�sr��>��9��@ׯ�4������� �k��1����{ʿ���=�ӿ;�
��t=��!y��-��3���ƞ�� ���I����
e��3*���� �����v�w�9�z��x��ù˾�t�����z���i���i��-tݾ���!&��rX���T�οֲ��DJ����E��c��sî�Y��S����W��|���뿌����X��\忪 ���P�G`��M�����,��{j��5K����P��Z���ֿ剘�b�_��*�Q�� �ᾁþ�p������������>�Ⱦ�@��m���4�S�n��E�����d$�GQ^�`�������f:�����^̚�����C������ؿ�Q��Ѯƿ)��� +��e�����P��@���O���t����y��*=����M��i숿>NK��k��?����վ�������H���|��\l���LҾ����Ji�d1E��3��-��޳�f�6��rr��>��#��$ׯ����W�����k��1�l���zʿ����%�ӿ��
�at=�g!y�r-����������Ӫ��#����
e��3*�%�񿬑��T�v���9��������˾�r��,���~���c���g��,rݾ���4&��qX������ο����DJ�y��5��U��hî�P��L����W�|���뿙���Y��~�� ���P�W`��_���2��D���j��RK��0�P��Z�p�ֿx�����_�>�*�������
þs��9����
��E���=�ȾhB꾴n���4��n�/F���违$��Q^����������:������̚�H����C�H����ؿ�R����ƿ�)��� +�Me�᪏�k��U���^��������y��*=�(��"N���숿>OK��l�tB��b�վc��������J��t��o��OҾ���Qj�K2E��  �  ܈���ſ����N��׉�T�������h������=٦����y�G����=޿�{˿P���:�kLV�p����:��(����.��~��T���&���V?�h��͵��^}�-�7�.����߾�U�����&A��*Z��X���g��:�;������!��oZ��5������#�x�d�`?��P��{-��G$���Z��,y��ʍt�o3�z��A�ҿ��Ͽ���\-��l��ט��̵�2K���=���µ�n����l��K*�=W�"���4�b���&�4� ���Ѿ�䳾c��⨚�T����]���Z��&�ھS��/�1�K�s��b������+8�*Q|����g����������y:���b����]��� �uB�%_̿y�ٿr����@����|�����o3��Fq��@<��<���f�U�}���Jο�Y��+zK��:��ﾭIƾ ֬�kΞ����mם��Ī���¾�������D��ۈ�W�ſ����N�{׉�C�������h������٦�m��
�G�j���<޿�z˿/��8:��KV�(����:�����w.��O��-������V?�8�b͵�^}�~�7�v���߾T��,
��F?��9X��^���e��F�;����ˮ!��nZ��5��C���#�R�d�O?��A��n-��<$���Z��&y��t�o3�|��N�ҿ��Ͽ?���r-�4�l��ט��̵�GK���=��
õ������l�L*��W꿳���a�b���&�r� �@�Ѿ6糾�e��A��������_���\����ھ-����1��s�Zc��0���+8�nQ|�������N��������:���b��M�]�W� ��C�.`̿p�ٿ���@�B���|��(����3��Tq��L<��G����U�����JοZ��{K��;�d��=Lƾ�ج�)ў�?	��ڝ�yǪ�i�¾�龿��ώD��  �  )����0˿g���V�����ű�mn���Z���v���1��ﶋ�%4P���q�֞ѿ��WC!��a_��œ�	޴�r%��c!��
a��V���҇�JG�ս	�[Y��BG��ʷ7��%
�y5۾έ��d���P���n ��y���Rͬ�WGɾ����	� ���[��<������*���n�2�����B�����v����X�����:����")ٿ�TֿsG��4�Tw�k���ս������2���˟��	w�1�I��g����bd��&��9���f;�E������m��qZ���蠾����[־F�h�1�ɫv��������к?�����bI��:��S���Z���� ��׿���+g�3A'�\k���ҿ5��8��~�H�Ĩ��歪�T��m!���)��������3�^�=�c9Կ徐�<NL����X�ڣ��
G���y���Ε����
<��� ��I������E������0˿E���V������ı�Xn���Z���v���1�������3P�s�p忼�ѿ����B!��`_�Pœ��ݴ�4%��-!���`��.���҇��IG���	�Y���F���7��$
��3۾$�������s����������Zˬ�gEɾ���#� ��[�#<����翫*���n�!�����5�����m����X�����:����/)ٿ�Tֿ�G��4�ow�{���!ս������K���˟�,
w�P1��������dd�5&�H<��xi;AH��;���qo���\���꠾����]־ZG�7�1���v�񄲿���?������I��i����������,�����],g��A'�ul���ҿ.�࿩����H�����3T���!���)�������J�^�\��9ԿH���(OL��	�[�a����I��Q|���ѕ������>��K#��|����}E��  �  ܈���ſ����N��׉�T�������h������=٦����y�G����=޿�{˿P���:�kLV�p����:��(����.��~��T���&���V?�h��͵��^}�-�7�.����߾�U�����&A��*Z��X���g��:�;������!��oZ��5������#�x�d�`?��P��{-��G$���Z��,y��ʍt�o3�z��A�ҿ��Ͽ���\-��l��ט��̵�2K���=���µ�n����l��K*�=W�"���4�b���&�4� ���Ѿ�䳾c��⨚�T����]���Z��&�ھS��/�1�K�s��b������+8�*Q|����g����������y:���b����]��� �uB�%_̿y�ٿr����@����|�����o3��Fq��@<��<���f�U�}���Jο�Y��+zK��:��ﾭIƾ ֬�kΞ����mם��Ī���¾�������D��ۈ�W�ſ����N�{׉�C�������h������٦�m��
�G�j���<޿�z˿/��8:��KV�(����:�����w.��O��-������V?�8�b͵�^}�~�7�v���߾T��,
��F?��9X��^���e��F�;����ˮ!��nZ��5��C���#�R�d�O?��A��n-��<$���Z��&y��t�o3�|��N�ҿ��Ͽ?���r-�4�l��ט��̵�GK���=��
õ������l�L*��W꿳���a�b���&�r� �@�Ѿ6糾�e��A��������_���\����ھ-����1��s�Zc��0���+8�nQ|�������N��������:���b��M�]�W� ��C�.`̿p�ٿ���@�B���|��(����3��Tq��L<��G����U�����JοZ��{K��;�d��=Lƾ�ج�)ў�?	��ڝ�yǪ�i�¾�龿��ώD��  �  74���������6�sr��>��9��@ׯ�4������� �k��1����{ʿ���=�ӿ;�
��t=��!y��-��3���ƞ�� ���I����
e��3*���� �����v�w�9�z��x��ù˾�t�����z���i���i��-tݾ���!&��rX���T�οֲ��DJ����E��c��sî�Y��S����W��|���뿌����X��\忪 ���P�G`��M�����,��{j��5K����P��Z���ֿ剘�b�_��*�Q�� �ᾁþ�p������������>�Ⱦ�@��m���4�S�n��E�����d$�GQ^�`�������f:�����^̚�����C������ؿ�Q��Ѯƿ)��� +��e�����P��@���O���t����y��*=����M��i숿>NK��k��?����վ�������H���|��\l���LҾ����Ji�d1E��3��-��޳�f�6��rr��>��#��$ׯ����W�����k��1�l���zʿ����%�ӿ��
�at=�g!y�r-����������Ӫ��#����
e��3*�%�񿬑��T�v���9��������˾�r��,���~���c���g��,rݾ���4&��qX������ο����DJ�y��5��U��hî�P��L����W�|���뿙���Y��~�� ���P�W`��_���2��D���j��RK��0�P��Z�p�ֿx�����_�>�*�������
þs��9����
��E���=�ȾhB꾴n���4��n�/F���违$��Q^����������:������̚�H����C�H����ؿ�R����ƿ�)��� +�Me�᪏�k��U���^��������y��*=�(��"N���숿>OK��l�tB��b�վc��������J��t��o��OҾ���Qj�K2E��  �  ��?��u�⿾b�"�E�i4q��3������k����l��M?�����zڿ�Ѯ�����Xϵ��V�y;���I��ru�>���#b�������@h��~;���^Կ&��={u�@�C�� ��|��龏kо6^¾�˿�K�Ⱦ�ݾ��������2��.]�p'���?������l '���T��r}�1D��ϲ���r���C^��/����vȿ�B��Ԅ���7ÿ����o`*�CY����������V���+�Y�*,�@���e���V����b���6����Q� ���wʾO7��ހ���Jξ�i�~�t��/h?�Jo��H��-tͿ�h
�n\6��c�����}��}���6�y�~O��2 �7��!㹿52��/諿bԿO��H	:�^�g�����k��w[��uu�%�J��9���꿨���WN��tR��W+�U����b�׾�žxZ���~ľuվ���]|�k�'�hM�����B?��&�⿚b���E�B4q�q3������I��8�l�UM?�-���yڿ�Ю�����Oε�zU��:�+�I�{ru�����a��r����@h��~;�����]Կ����zu���C�d� ��{�`�龸iо?\¾zɿ�1�Ⱦ�ݾ��������2��-]�'��I?��.���C '�p�T��r}�$D��Ĳ���r���C^��/����vȿ�B��넥�8ÿ����`*�3CY��������%��q���e�Y�F*,����f��gW����b�+�6�C���� ���Szʾ�9��5���Mξ�k�g�G���h?� o�DI���tͿ�h
��\6�[�c�������������y��O�V3 �>��"乿+3��髿5Կ����	:���g�3����k���[��2uu�D�J�:��������N��*uR��X+�������T�׾�žr]��܁ľ?վ`�}���'��hM��  �  �܇�!���9~ǿ���������6�/�K�ъR���H�&�0�ѻ�B��4$������������Ǹ�q￦�}7��eL�	kR�&�G���0���X�쿪;���㛿�삿�n_���?���$��k��������`德��O�()��+3�)�P�x�s��ޏ�v�����ֿ@����#���>���O�=&Q��(B��&����ο�����Q��S��ힿ�ɿ\��#�-�?�DP��P�MA��'�5#	���ۿ��������x�DT�396�/��H8����徏��P��<G�`�!���<���[�Ϗ��A����ֹ��翚��wx-�d�E�f
R���M��:������������9f���s��Ȗ��?����6ۿ
�*q-���F��IR��"M��l9�Y!����|\̿����q��8Pk���I��6-�	B��������뾒
�����Q*�|TF�tCg�܇������}ǿ����u��^�6� �K���R���H���0�y��}��]#��0����
��%����Ƹ�z�/�7�3eL��jR���G�r�0�����c;���㛿\삿n_���?��$��j�(�������^征��wN�(��*3�$�P���s�9ޏ����%�ֿ����#���>�߯O�%&Q��(B��&����ο�����Q��j��.ힿ�ɿx�#�S�?�DDP�K�P�CMA��'�u#	��ۿ����Q���,x�gET��:6�����9�%��9����羌��@H�H�!�w�<�Z�[�#��������ֹ�G�Ҽ��x-���E��
R��M�Z:�����������*g���t���������W7ۿd
�nq-��F��IR�#M�m9�!����\̿	��0r��mQk��I�8-��C�x��G������������R*��UF�yDg��  �  23��=���>����տ����L���Y_�o�W��AEѿf���+��kh��]��n��g��-����ڿ�E�Ї������@H�$a�,Rп���\�������Y�����w�\�U�V�6��f��)��� ��m�*��AG�L�h��`��T��	���E���ƿ�޿6���et� ��
�ߑ�{2�	:ÿx���. ��u^a�ļ_��6{�ܘ�T���ȥ远��+X��Ŷ�l�����A�ȿZ ��:���Y��m8��Wml�U�J�5�-�Ip����iF��H�Kz3��R�1t�`܊��Q��G꨿����ǦͿ;(迭��o�s��c���7�aa߿��������Ħr���]���e�H��L�����̿��ū���ъ����"1��S�ؿu������Ϡ��鑿����`��[@�bx%�i���E[�H�"�/=��2]����-���2���󭿴=��2�տ���L����#_�/�{V���Dѿ����H*��fih�]�:�n��f��9,��ӰڿiE�v��W��v�H��`��Qпg��'����������2�w���U�t�6��e��(���Ӷ�>�*�t@G�*�h�D`���S�����@E��gƿ��޿����Bt����	�ˑ�^2��9ÿo���0 ���^a��_��6{�9ܘ����������XX�8�������.��Ћȿ� ��ܦ����9���nl���J���-��q����G��I�S{3��R��t��܊�R���꨿�����Ϳ�(�����Ŕ����K8�9b߿����������r���]�O�e��H��������̿��� ����������|1����ؿ�u������3Р��ꑿŤ����`�P]@�z%�$�����\���"��=��3]�M��S.���  �  �ѿ+�տnԿQ�ѿ�ѿ`>Կ��տ�Kѿ�?Ŀ?)������y�3BQ�I�7�ˬ0�<�Y�q��N���c����ǿ��ҿ`�տ�ӿKdѿ"ҿ��Կ6vտ��Ͽe9�����Be��Rr���K�~x5��I1�s�?��e_�~ ���џ�J"��Peʿ��ӿ+�տ{!ӿ�Dѿ�cҿ�տ1տ��Ϳ����즿{����j���F�"x3�1l2��C�<f�$K����4���`�̿<�Կ/Nտ��ҿ"<ѿ �ҿ�fտ�uԿ��˿Z��������䈿��c�|B���1�t4�o�H�Z$m�����R������ο�7տ��Կ�AҿvLѿ�Iӿv�տ��ӿ �ɿ�涿a��9����=]���>� 1��>6���M�͂t�wԒ��u���A¿�Jп�տb�Կ��ѿxsѿ��ӿK�տk�ҿǿU��v������!W���:���0���8��"S�],|�.(���|���4ſ��ѿ��տԿ��ѿ��ѿ
>ԿK�տ)Kѿ�?Ŀ�(��i�����y��@Q���7�3�0�n<��Y�����~��c���ǿ�ҿ�տ��ӿdѿ�ҿ�ԿvտX�Ͽ*9������d��hr�~�K�Yw5��H1�2�?��d_����!џ��!���dʿG�ӿ��տ!ӿBDѿzcҿKտ�տU�Ϳ�����즿g����j���F�;x3�`l2�c�C��f�]K��J��������̿��Կ�Nտy�ҿ�<ѿ��ҿegտUvԿ��˿���T����刿�c���B��1��4���H�i%m�����RS����Q�ο�7տ��Կ�Aҿ�LѿJӿ�տ��ӿ��ɿ�綿�a���S?]�[�>��1�k@6�)�M��t�Ւ�Bv��B¿lKпq�տƋԿ �ѿ�sѿ�ӿ�տ�ҿ�ǿ'��V��淀��W�i�:�]�0�h�8��$S��-|��(���}��E5ſ�  �  %|��e����5D�LwԿ	)����Ed��gN��;�}��Q[�8a;��!�g����b��&��B���b�����ƒ�\�������¿Z?ڿ����q	�e�����!�
�N���7ʿj~��
烿�}d�0�]�:�t�?y��"ѷ�^��*�����dw����Ï濵X̿�����-��N����,r�P4P�h�1��F����r9��Z��/�Z�L�Xn�?#���֗�v�������ɿWf��Q �Q�dE�H�����Y�ZU��'��g�x��_�Qb�8B�������ſ�q��a	�W��s���
����&=ݿ��Ŀ?\��Q:��{���r��?�f��E�$f)�����T����6���&8��W���y�����Ĝ��g�������ѿ ���ւ�k�����%E �cVؿ ���Ȍ��"m���\���i�{������ܟӿ�o��|���{��e�x���C��vԿ�(������c���M��3�}��P[��_;���!������(a���&��B���b�����2ƒ�흡�Ǒ��͗¿2?ڿ{���q	�[������
���7ʿ�}��}惿�|d���]��t��x��wз�����)�n�Ł�#w����Z��XX̿�������~��!���o,r�&4P�T�1��F�����9��Z�/�ΕL��Xn��#��Tח��v��<��(�ɿ�f�/R �bQ��E�������Y�!V�������x�<_�wRb��B��-�����ſr�b	�W��s���
����a=ݿF�Ŀ�\���:���{��Ns����f���E��g)�Q��TV������(8�*�W���y�����3Ŝ�fh������ѿ� �<�,��˝�$���E �YWؿ���Ɍ��$m���\���i�f���뺪���ӿlp��̹��  �  �R��J��5������Gſ}۠�U����Fe��D���(�����= ��뾱��ф���v�ү.��qK��`m��ċ��맿|�ο@�3��%�:�l�M�$R�/�E���+��2�Wؿ��������È��}���Z}����5};���N���Q�n�D���+����;�9����.����~�x�Y��:��� ��<�=���$7�'U澳$��G5	�\��5�7�!V��Gz�.��ˈ����޿x�
�2�(��B�Q��O�,D>��:!��J ��+ƿY1���q��3����ѿ���7P(��`C�P�Q�O�o�=�� "��H�K�ӿq����z����q���N���1�~���`�>���%�8��aa��t�� &�<ZA�"[a�!!�������|��r��;���2���H���R���K���5�`F����E���5��q�������8t����俫��L_2�J�I�ƖR��J��5��������ſ"۠�񘆿�Ee�#�D���(�y���< ������2��vu���.��pK��_m��ċ�I맿T�ο6�1��%�:�j�M�R��E���+��2��ؿb���Q���j�4ģ���|������|;�j�N�`�Q�)�D�q�+�p��;�䲷��.��v�~��Y���:�i� ��<�A���T7羅U�@%���5	������7��V�MHz��.��G���D�޿��
���(�v�B�^Q�|�O��D>�a;!�YK ��,ƿ&2������*	��ڄ����ѿ���eP(��`C�e�Q�+O�{�=�� "��H���ӿ¦��{���q���N���1����Vb����(�ߐ��c�����&�H[A�\a��!�����}����ￄ��2���H�+�R�'�K�:�5��F���G��7����Ñ�4u��~�����_2���I��  �  푍����o��3C�)���8߿J�������J�&�5�U'ﾯ�ӾZ�þ4k���{ƾ��ؾR���My��0-��U��4���{�����#��kM���w�����K�����+�e��h7��
�=ѿ���q��������󿆷"�КQ�D�{������܌�-+���4a�*�3�X+�Jʿ����7�k��:=��#��������I;�!��"}��4`˾������h�8�p�e�������ÿ���I�.��_\�x���T���ċ��}��V�4�'�ǝ��!����ʤ�hF��W:˿0?��*2���`�5K��Q��E׊���{��wR���$�����D��� ���jZ���0��=�7���^�۾��Ǿ���K�¾1�Ѿ)�뾢����"��3F�`�x�Ⅱ�P�׿VI�U>���j��9��g{������@Ls��0G������F鳿cx���j����ݿ���S�A���n�����Ǒ�����o��3C�����8߿񝦿L���J�&�	4�%�V�Ӿ��þ�h��(yƾK�ؾ���Dx�0-�U�l4��Y{�����"��kM���w�����K������e�Lh7�ٯ
��ѿm�������
�����&�"�s�Q��{������܌�	+��u4a���3�#+��ʿq�����k�):=��#�_������I;""���}���`˾B��^�����8�6�e�%���;�ÿ����.�I`\�2x���T���ċ�~���V���'���������{ˤ�*G��;˿|?��*2��`�EK��Y��I׊� �{��wR� $����RD��� ��kZ���0��>������۾,�Ǿ������¾��Ѿ}�뾼����"��4F�X�x�^�����׿�I��>�݊j��9���{��9���Ls�N1G����'��o곿�y���k����ݿZ����A��n�+����  �  *ۯ�GI��2ٓ��o�c�3�r/ �����큿k?B��z�V��3�о�c�����V��� ���ļ� �׾�� ��� zN�y_���
ÿz�
�j@��e|��G��;5��P��������*����a�.(�{.����Ŀ�㻿��ۿ9'�@G�����i����������H������d�Z�,!�P��<����j��1��������2Ǿ�β�L����4��/3��_ľ����x	��-�6)c�0^��&<ۿ@=��@T��߇�ԋ��8K����[���Ą���M�cU�e��Of������C��gL"���Z�u�����_���i���ӛ��x����F���.�ʿ$s���
U�2�#�]��z۾�'��c[��Ѐ��� ���d���M;�U񾀻���<�K{�8ԭ�����J-��fh�����M�������r���Җ��u�ZK:�o��!ѿw_����̿G���4��o�	��ۄ��ۯ�'I��ٓ��o�8�3�H/ �����=큿�>B��y�T���о�a��k���S��a��[¼��׾�� �"�}yN�@_���
ÿw�
�j@��e|��G��A5��P�������*��d�a��(��-����Ŀ㻿��ۿ�&��G�Ȅ��<��|���{���!�������&�Z��!�����;���j���1�j��*���2Ǿ�β�|���65���3���_ľ��㾆y	�{-� *c��^���<ۿ�=�3AT��߇����iK���������*ń�j�M��U�C��%g��K�����￶L"� �Z�������f���i���ӛ��x����F���c�ʿos���U��#�
^��|۾*���]��C���d#���f���O;�W񾌼���<�I{��ԭ�����;K-�gh�������������'Ӗ���u��K:��o�#ѿ�`��ǒ̿���p4�o�A	��	����  �  �n�����!�����EXJ���������7��,:A�>���E���̩�\i��b��zW����Ⱦ�f����O�Y4��նҿs��QjY�֘��t���l3��3���߻��ġ�T���m=�Pi	�h�׿=Ϳ���#�,za�kE��^���ء��)s��)����V���hx�p�4�'���Ъ��ko���.�)��ؾ*﷾P���AV���ܚ�
�� 4��1Ծ����m)��f��룿`��-�ޘp�4�y��>�������v������fi�$�)������ο�-Կ���϶6�vix�B������|������Ϩ���`��za��V ��ۿ�!��/�V��:��e����˾?4��x���9��䚜�Z짾iཾR�b���:�>!��p��������B�b���:��_���Q������㭫�٪��%�R��z�v濭A˿���s.��fK�"ч��|������n�����������XJ�Բ�����:7��`9A�]���C�����ɩ�g����?U���쭾�Ⱦ&e�6��?O�)4����ҿt��]jY�����~���t3��4���߻��ġ�8��6m=��h	���׿q
Ϳ��0�#��ya�:E��0��������r������V��Chx�8�4������Ϫ�]ko���.��(��ؾ�O���pV���ܚ�����4��$Ծ��sn)��f�:죿�`�7�-�/�p�`����o��������v��! ���i���)������ο�.Կ��!�6��ix��B��#����|������̨���`��{a�W �8�ۿ"���V��;��g����˾�6��oz��6<��B�����⽾|�m��	�:��!��󥹿�����B�����:������Q��Ҵ��-���&���šR�9{����B˿γ�/�0gK�^ч�}������  �  � ����������6�� �m��W$���ۿW��VtP�F����)Ǿ`,��G��L���� ��ߒ��/�ξ�/��L	$���`�Tk���g�,3����.������$���~~��C���X��͝��q�]�=�����������
��>��g��H��5���v��]���4z�������=���rS����"�� 1��i^;���P��3F�������]o��4��<X����۾�%	��5�"|��׷��	��K����pT�����"���G����Z��\�������)F�(b����6���<�ƚU�,���7���`��/���!z��l>��ѣ��U]����:�j���р��A<i��h)�����ҾQ���gP���ŝ�+B���/����þ+�W���
I�RO��
ҿ�H�߰d��������e�����������A��Q�� w�>	1��I��������]�*�rn�Wş��@�����f ������������Ոm�VW$�>�ۿ�V���sP�c����'Ǿ6*��������������5�ξ.���$��`�#k���g�,3����.������*���}~��9���X������$�]���������u�
���>��g���G�����v��4���z�������=���rS�����"���0��^;�X��� F��������o������X����۾O&	��5��"|�Wط�_�	�	K�:����T�����S���{����Z��������N*F��b������5=��U�N��8���`��6���#z��k>��ϣ��V]����:���������<i��i)����*�Ҿ����R���ǝ��D��2��?�þ<-�f���I��O���
ҿ�H�-�d������������ ����������ZQ���w��	1�9J����%����*��rn��ş��@��@����  �  ����=��!���ED��x�c��Z�/�տ+	��V�O�|��o����/̾|
�������"���ʧ�#����Ӿ�� �F4%��P_�It���8��e,�@�t�9���������%l������\��KZ����T�����1�[���8�{j7��}�����C��ƛ��/���Y�������
����J���&���¸��"�;�D���徢G¾�l���}�������ҫ��U��P��,�ݞ5�Ƭy��������C����������N��a���,���%f���<���A��b>��a
����)鿘���M�K����i���%��^��������>��r2���}���3�f��W,��ãg��d*���w�׾����XL��'ڤ�5��,�Ⱦ���&���H��M��*�̿���][�-���UF��l������`O������t����l��M*�J����޿ƚ��0$���d��������T�������=�����-D��L�c��Z�֟տ�����O����~���-̾M��{���� ��rȧ��|����Ӿ�� ��3%�9P_�t���8��e,�J�t�A���������$l������\��.Z����T�t���0��࿉8�j7���}����eC���������2�������
����J���ԏ��������;�������pG¾�l���}��I���8ӫ�VV��D������5���y�3������C�����쀮�(O������`���Zf���<���A���b>�Gb
���������M�m��� j���%��f��������>��q2���}���3����,��{�g��e*�����׾7���~���N���ܤ����p�Ⱦ���'��H�AN����̿f��?^[�X����F����������O��9���5u��%�l�BN*�����L�޿����0$��d��������T���  �  i7��٭��୦����ΨI�6��]qƿ������P�b�!����O�ܾ��¾�Y���c��O���Z~Ǿv��u���*� V^�=�����ֿ���%XX��?��Xˬ�����U��� ��dS��D5~�!a<�H	�?�׿TͿ�c��'#��_�	��>��������3���e������X�v��4�����dc����}�e�>����;����Ҿ~���I䱾�S����ƳϾӀ�r��[9�Yu�2���f��i�-��n�.��^���]r�����B�������Xkg�Z!)�xt��bϿE]Կj����5���v�wޜ�\����T���S��K���`��F�_��� ���߿yZ��Ơe��;/�������1ʾ��Б��ve�������YپQ- �ۤ�{~J��������p	��{B�����r��»�����������މ���KQ������ɐ˿е���8*J������������B7������ĭ��鹆���I���qƿ|�����P�x�!����,�ܾ��¾3W��Qa������|ǾV�侀��:�*�wU^� �����ֿ���)XX��?��_ˬ�����T��� ��PS��5~��`<��	���׿=SͿ�b�'#���_�O	�����k����3���e�������v�Ԉ4�B���c�� �}� �>���.;��k�Ҿ~���y䱾�S�������ϾŁ�,s�L\9��Yu��������-�b�n�I.�������r��?���v���ƶ���kg��!)�Uu��8Ͽ^Կƫ���5���v��ޜ�k����T���S��K���b��N�_��� ��߿�Z����e��</�����辔ʾ���H����g�����)\پk. ����J�I��4����	��{B�����r��J»����ĵ����)����LQ�C������˿��࿛���*J�ֽ����������  �  8���1Ә�����d[�;�'�������tU��fZ���1�0Y�9��Mxྑ6Ͼ	Yʾk�Ѿ���`-���8j9��Be�����r¿KF�
�2��g�s��q��~T��,���a��� N�r�����'��%��Nο`H�sf6��l�F�������<ў��֓�Ӓ}��I�����޿�v����~�� K�B�&��v����Yپ\3̾9�˾�G׾*]�P
��p#�YF���w��h���׿�����C��x�	���6��ޞ��\��N�q�X><����#�ӿHe��k����߿,��
 H��A}����k�����������l��d8����tɿF���0k��=����^���辫�ӾM�ʾ6ξ:�ݾ�$������-��T�|��H���x��,"��U����fL�������p���)��/+`�`�*�eR��U�Ŀ4���)���@O���n%��*Z�&���������Ә����d[��'��������U���Z��1�'X�����u�4Ͼ�Vʾ��Ѿh��8,���Ki9��Ae�M����q¿>F��2��g�s��q��{T��!���a��� N�-����u��h��SMο�G�f6�fl��������ў�z֓���}���I����H�޿@v��c�~�B K���&�|v���� Zپ�3̾��˾�H׾�]��
�.q#��YF�Y�w�Si��e׿�����C�x�6���6����������q��><������ӿf���k��C�߿x��I H�(B}����t��
���������l��d8�����ɿ�����0k��=����_���A�Ӿ�ʾ�ξ��ݾ9'�� ���-��T��|���H��@y�+-"�n�U�����L��ֆ��7q��>*���+`���*��S��~�ĿV���@���IP��Vo%�+Z�Y�������  �  �m�Ld��3K���)�c-�wLؿ	��`���0w��`S�x�4�����|�S������[���$�� �SN;� �Z����!e�����vx��Q��1���Q�ؒg���l�Ww^���@��}�@0�ل��J���!��r����5Կ��
���0���R�9�h�Pl��1]�0�@��H����(�ȿ'������Z�j�ղH�#�+�����\d���m���K��I�	)�JBE�s}f��+���ɠ��5Ŀ�����y���<�|�Z�DNk���i��V�T�4����ɓڿ�s�������̗��۳�e�lE�w�<��[�<�k�
i�&�T� c5����(W�R?���j��<]��$�^���>��v#������"#�������e/���1���O�O�r��玿gD��	�ҿ¶���%�Q�G�r�a�!�l�]'e�B	L�Z9(���Fȿ�'�����	Y����¿�����#�NmH�U"c�Wm�d��3K�Y�)�6-�Lؿ�������1/w��_S�a�4�v���{�����[��.Y��#��� �#M;��Z�T���d�����Ix��Q��1���Q�Ԓg�w�l�@w^���@��}��/�A�������o�������4Կ)�
���0���R��h�l�p1]��@��H�K����ȿ�&��¬����j���H���+� �����d��Bn���K�@J�~	)��BE�~f�,���ɠ�G6ĿA���2z�5�<�ӐZ��Nk���i�_V���4�����ڿPt��w���͗�6ܳ��迨E���<�%�[�S�k�-
i�4�T�0c5����hW鿧?���j���]��G�^��>�Jx#�p������%�v���J���0���1���O�N�r�u莿�D����ҿ���%���G���a���l��'e��	L��9(����&Gȿ)��� ��Z����¿o��3�#��mH��"c��  �  -�%�u:"����E��3^���Ͽ����^����כ�������l���I��:-����#b��h���2��P��bu�Z����������������Կ5
���.����#�??%��!�i����߿����/���bv�Io�RV���栿>sʿ���ed�4"�5�%����5,�0L��2�H�ȿ�3�����S땿*0��s�`�r?��&�X�����#���;�c�\�B���擿�F��f��z�ƿ�ݿס���M��s�̠%��#��{�����k�Ͽj�������j@p���s�j/������0ڿ�!�@\�8�$�ѥ$����T�
���g�׿I�¿�Ա������Ώ���y�u�T�c�5�G �՟��J�O�*��E���h�n���㙿`����ݺ��wͿ�)濦����0!��&���������]Z���H������m�	~|�L���6v��\W꿼���P���%�8:"�i�����]鿕�Ͽ<������yכ������l�g�I��9-�4���`�g�+�2���P�jau��������\��<�����Կ
���"��z�#�-?%��!�C��.�߿]�� /���av��o��U��"栿�rʿl���d��"���%�Q���+��K������ȿh3��r��'땿	0��H�`�^?��&�+X�7��6�#�'�;�ם\�����擿�F���f���ƿYݿh���*N�t�$�%��#��{�����2�Ͽ1������Ap� �s�
0������Z1ڿ�!�e\�T�$��$����m�
��󿻉׿��¿sձ�s���.Ϗ��y���T��5�� �L���K���*�W�E���h�o��"䙿ն���ݺ�(xͿ*����_��r0!�V&���+�����^[���I������m��|�8���w��'X���Q��  �  vc翛l�W���忶�忰C�Sj�1��<Tؿ9y��/����y��j�a�d^E�
8=�.�I�}cj��f��.��fƿ3vܿ���2U�p迳��Vd���%B�1���Կ�ܻ�^����6��>�[�3�B��=��N��|q�������ţʿf;߿���E����t�[��d��꿺3�Aѿ�"���噿@~��V��U@��*?�K�R�7y����
ﳿ�ο��R�꿂��`<�+j��l���pG�[���ZͿ�Q�� ���sv�QQ���>�A���W�Tw����������t�ҿ���+	�X8�ʴ濤~�1�I.��k鿧V޿�>ɿBr��]s���o���L���=��nC���]�眄�]��Oi���ֿ����T�u��)?����դ�@a�K��xۿ��Ŀ����c䋿Kh�[�H�,=��kF�(�c��툿YC��j����gٿ�b�'l��鿝��_��VC��i���濿Sؿ�x������y����a��\E�o6=���I��aj��e��J-��^eƿ�uܿ4�迿T��o�o��$d�����A��0忟�Կ]ܻ�����6��1�[��B���=�SN�H{q�G���y��0�ʿ�:߿v������bt��濻c���꿆3��@ѿ�"���噿�?~��V��U@�#+?���R��y�?���Oﳿe�οL�Ώ������<翶j心m翲��H��࿜[Ϳ�R��� ��uv��Q��>�`A���W��w��e������Āҿ��g	뿔8����~忙��.�bl�PW޿c?ɿs��+t���o�#�L�B�=�9pC��]������]���i��bֿ��aU�ݩ鿖?�o��_���a뿸K迒yۿ��Ŀ؊��O勿-h�=�H�=��mF��c��D�����jhٿ�  �  nd��ɰ���ѿ� �#�� o���"�N�%�&��a�ˣ���9����z���m����� ����¿t���^ ��&�� �����������M̿��ѩ�蘿�_��m�f�6D�Wx)����[��� ��#7��V�(�{��֐�����ٸ���ÿ�ؿ�A��Ow�@G�8�$��W$��n������׿�U�����r��q�G��G���>ҿ�;�~�u�#��n%�����\�����j�ۿ�ſ�����Z��Ⓙ?�� �Z��<:�^�"��L�����!'���@���b�)@��w떿������bʿ��� �l�&n��&�5�!�.O�����s�ǿ� 2����n���w������Y��=�J��@���y%�ʒ#������V�:�ӿ����*��p��������Ds�mO�=H1�����P��+�U�.�"YK��o�_���2Ϝ��c��]���^ѿ� �����n���"��%����`�$��f��p��F�z��m�������¿7s�J�w^ �Q&��� �������[�俎M̿���Щ��瘿�_����f�+5D�Xw)����7���� ��"7�ĲV��{�=֐����_���}�ÿ��ؿDA��&w�G��$��W$�un������׿�U�����r��q�i��u��(?ҿ�;�-~���#�o%�Ŀ��\�C�����ۿz�ſV���o[���Ⓙ���k�Z�_>:���"�:N�)���"'���@�w�b��@���떿:��5���ʿև�7 ���pn�&���!��O�����U�ǿg 3��m�n���w�^���MZ���=⿎��{���y%���#��H��%W�ӿ�����+�� ���~���uFs�O��I1�>��eR�--��.��ZK�.o������Ϝ��  �  T��>���5ۿ��	�i�+��L��d�,m��b���F�=�!��A���������>������<(˿6���W*���M�qf��l���`�0F��$�^�kпgp�������p�0�M��_0�Y�����><��dc�L` �����$��7@���`�'��������l���X�h���I7�iRV���i��uk��qZ��:�Q,�0�俙������������p����ݿ����6�܇W��vj���j�l0Y�%;�4���~�i����&�����~d�z�C�~�'�K5������������o�t��gc-�TpJ���l�K􊿊᥿�e˿�W���2 �[nB��q^��gl�q�g��1Q���.����ѿg�������츚�U����������B���_���l�~�f�4(P�b�/�$��ۚ࿂����땿^�}�j�X�h�9�Yx��0�Q��B��Ni���\	�.���6�x5U��_y���������ۿ��	�A�+���L���d��m�Yb�f�F���!�A���������=������A'˿���:W*���M�f���l�S�`��F��$�3��jп!p������0�p���M��^0�z�����0:��<a�1_ �����$��6@���`�����S���Rl��MX�=���I7�HRV���i��uk��qZ��:�H,�(�俜�������ʔ���p����ݿ����6��W��vj�&�j��0Y�a;�t��V�����1'��M�F�d�ҐC�ڞ'��6���f������p�y��Rd-�$qJ�a�l����᥿,f˿�W��3 ��nB��q^�\hl���g�2Q�6�.�~���ѿY���x���Ź�����^��6����B���_�%�l���f�[(P���/�O��A������앿��}���X��9��y�(2�PT��u��ll��^	����V�6��6U��`y��  �  �R�����1,��#V*�:R^�Cއ�ш��=����S���^���(W���"��v����0㰿
ǿR� � �-��(c��a��6��zi���{��ʂ�i�R����rd�O|��7���EUR�},��M��A����ܾ!�;'�ʾ*wԾ�꾦�����2�?��?n��@��:u̿�J��B;�ʧo�YΎ�y������u���tz�#E�e���ܿ?��(<��&�ֿI@��1?���t�!��q���ٝ�>���Ku��	A��%��}ӿ����(�t�;D��!�������wL־�5˾�̾YpھH���+��_�(��eM����t���t⿇C��L�#������t���5��伌��i���3�[���˿����=���꿇\��"Q�ں������w���ך�pG���&d���/���d?��p��bb�Md7�B����.��O9Ѿ+Gʾi�Ͼ ��� �,���v3���\�\R������+���U*�R^�/އ����� ���kS��w^��_(W�H�"��u����/ⰿǿ˽ �z�-�N(c��a�����Hi���{���ɂ�,�R�]��d��{��韄��TR��,�M�=@�� �ܾ(�;�ʾuԾ�}꾜����;�?��>n��@���t̿�J��B;���o�IΎ�k������l���tz��"E�a���ܿ?��?<��H�ֿ_@��1?��t�4�����ڝ�Y���Ku��	A�5&��~ӿ����b�t��D�l�!����C��O־O8˾a�̾�rھN�����5�(�EfM�������Vu⿿C�I�L�7#���������6��"���ui�E�3�����˿����"������\�#Q�����"����w���ך��G���&d���/���?���p��'cb��e7����2�&��R<Ѿ+JʾW�Ͼ���L	 �d��x3���\��  �  ����oʿ8���JM������@��K���r3�����bT���Մ�9�F�o2�gI޿;�˿ ��6����T��m��`���W��5��������ˡ������>�QR�Y��󭅿:wG���9���Q�׾�����������֬���m˾����g���1�ji��T���h��#��c�ȓ�����������Ջ�����L�r�H�2����B�ҿ]/п�5���4,��/k������	���-�����Ӳ���e���'k��y*�*��|����Dq��6�̹�s7ﾆ;ξJ2��>���7��!���WԾݬ��F����A�&��س�u� ���7��fz��i����������������~-���=\�XA ��P�̿8�ٿ0`���?�������������w7���O���a��ТT���.�ҿ�ڔ���Z��>(�
0�Γ�?ƾT����T���۴�|�þ��޾zI���#�T�����.oʿ���JM�{����@��3���U3�����8T���Մ�ͧF��1�hH޿-�˿�迨���T�qm�����������Z���dˡ����Y�>�!R��������vG�I��������׾ǘ���������Ϊ���k˾����f���1�@ii��T��kh���#�ɕc��Ǔ��
����������̋�����D�r�D�2����O�ҿt/п6���4,�0k������	���-��1������e��!(k��y*��������Eq�%�6��� :�>ξ�4������9��K���
YԾ����"����A�����س��� ���7��fz�$j��"�����������Ǐ���-��>\��A �&�Q�̿'�ٿ�`���?��������������7���O���a���T�����ҿ_۔���Z��?(�M1�����Aƾ0���W���޴�)�þ��޾�J���#�T��  �  ���cZڿ�!�)h�Ns��ƿ��A��X����B��~�����@�`�?!�y�����޿ğ ��y-�%-q�����~B��'8���������a��"����7W�m�yȿ�����iE���6�Ǿ����y���n��,���=��I�پ���&-���k���$��P�7����BM�������6���o��|����f��zȉ��PI��B��5���z��V�A��l��P��Y���9{��j��C����t��wi��*(?�Z,����t���2��G	��k޾!콾7���â��ȣ��E��,�þ��Q����>�	C��裿��rO��@������	e�����,���B������V�y��4��D���߿m�����X�f���L��?���P���.!���E���ɟ���p���(�&�79���O[��"��r����Ѿ�P���7��@��#.�������;�f�����H�S�"��Zڿ��!�h�>s��
ƿ��A��<����B��T�����Ѯ`��>!�r�����޿4� �8y-��,q�U���;B���7���������^a�� ����7W��l�ȿ.���5iE��o4�WǾ����w���l��0���;��U�پ���?-��k������#��%�7����1M�������6���o��s����f��vȉ��PI�C��5��俋��l�A��l��P��k���N{��&j��]����t���i��j(?��,�Uﯿ��t��2�1I	�en޾�����Ţ�$ˣ��G��-�þj�/��r�>�oC��P���G��O�A��ҁ��8e��3��i�����������y�Z4�4E���߿b��}��Q�X�����*L��Z���d���>!���E���ɟ���p���(�e&俟9���P[�7�"��t����Ѿ�S��Q:�����0��F��^ ξ�h�����,�S��  �  �z��@��$�'�(r��c���c��[��o��������R��}���/j�'�����Q��3�H`4�"z{���q���;���W����s������k1���R`�'��1eͿ�j��}E��R�mq辋¾�A��'䟾9睾����|G��UվƩ��5,���m�i0��"� ���>�]����ׯ�����P1���r��m������v����Q����ߢ�0V�,���I��.���׳����Pp��q��f��T0��I����F�-��۳��6w�2��D��{پ.񸾊U��9���7���z��;�X/㾸�w�>��ۅ��qĿz)�ĲW�~���՛��
���E5��;���`]��G���*��NF;��������o���!�i�a����]^���a��Q����������W���{��`/�>
����+W\�s!����E�̾h����������ƍ���4����Ⱦ��|��NT�(z���� �'�r��c���c��D��S��������R���|��/j��~'�����9�忡��_4��y{�z���-������� ���{s��Ԩ��I1��_R`�����dͿ�j��P|E��Q��o�����@��G⟾I坾�����E��eվ֨��4,���m�0���� �c�>�J����ׯ�����C1���r��d������r����Q������GV�<��1�I��.���׳�&���ep���q�����p0��2I��'�F�q���۳��7w�;2��E�H~پ���W���;��:���|��Ͼ�61㾘�J�>�2܅�rĿ�)��W���������:���{5��y����]�����++���F;�#������p����!���a�����^���a��f����������b���{��`/��
�6��X\�3t!�h�����̾�j����������s���v7��M�ȾE��}��OT��  �  ���cZڿ�!�)h�Ns��ƿ��A��X����B��~�����@�`�?!�y�����޿ğ ��y-�%-q�����~B��'8���������a��"����7W�m�yȿ�����iE���6�Ǿ����y���n��,���=��I�پ���&-���k���$��P�7����BM�������6���o��|����f��zȉ��PI��B��5���z��V�A��l��P��Y���9{��j��C����t��wi��*(?�Z,����t���2��G	��k޾!콾7���â��ȣ��E��,�þ��Q����>�	C��裿��rO��@������	e�����,���B������V�y��4��D���߿m�����X�f���L��?���P���.!���E���ɟ���p���(�&�79���O[��"��r����Ѿ�P���7��@��#.�������;�f�����H�S�"��Zڿ��!�h�>s��
ƿ��A��<����B��T�����Ѯ`��>!�r�����޿4� �8y-��,q�U���;B���7���������^a�� ����7W��l�ȿ.���5iE��o4�WǾ����w���l��0���;��U�پ���?-��k������#��%�7����1M�������6���o��s����f��vȉ��PI�C��5��俋��l�A��l��P��k���N{��&j��]����t���i��j(?��,�Uﯿ��t��2�1I	�en޾�����Ţ�$ˣ��G��-�þj�/��r�>�oC��P���G��O�A��ҁ��8e��3��i�����������y�Z4�4E���߿b��}��Q�X�����*L��Z���d���>!���E���ɟ���p���(�e&俟9���P[�7�"��t����Ѿ�S��Q:�����0��F��^ ξ�h�����,�S��  �  ����oʿ8���JM������@��K���r3�����bT���Մ�9�F�o2�gI޿;�˿ ��6����T��m��`���W��5��������ˡ������>�QR�Y��󭅿:wG���9���Q�׾�����������֬���m˾����g���1�ji��T���h��#��c�ȓ�����������Ջ�����L�r�H�2����B�ҿ]/п�5���4,��/k������	���-�����Ӳ���e���'k��y*�*��|����Dq��6�̹�s7ﾆ;ξJ2��>���7��!���WԾݬ��F����A�&��س�u� ���7��fz��i����������������~-���=\�XA ��P�̿8�ٿ0`���?�������������w7���O���a��ТT���.�ҿ�ڔ���Z��>(�
0�Γ�?ƾT����T���۴�|�þ��޾zI���#�T�����.oʿ���JM�{����@��3���U3�����8T���Մ�ͧF��1�hH޿-�˿�迨���T�qm�����������Z���dˡ����Y�>�!R��������vG�I��������׾ǘ���������Ϊ���k˾����f���1�@ii��T��kh���#�ɕc��Ǔ��
����������̋�����D�r�D�2����O�ҿt/п6���4,�0k������	���-��1������e��!(k��y*��������Eq�%�6��� :�>ξ�4������9��K���
YԾ����"����A�����س��� ���7��fz�$j��"�����������Ǐ���-��>\��A �&�Q�̿'�ٿ�`���?��������������7���O���a���T�����ҿ_۔���Z��?(�M1�����Aƾ0���W���޴�)�þ��޾�J���#�T��  �  �R�����1,��#V*�:R^�Cއ�ш��=����S���^���(W���"��v����0㰿
ǿR� � �-��(c��a��6��zi���{��ʂ�i�R����rd�O|��7���EUR�},��M��A����ܾ!�;'�ʾ*wԾ�꾦�����2�?��?n��@��:u̿�J��B;�ʧo�YΎ�y������u���tz�#E�e���ܿ?��(<��&�ֿI@��1?���t�!��q���ٝ�>���Ku��	A��%��}ӿ����(�t�;D��!�������wL־�5˾�̾YpھH���+��_�(��eM����t���t⿇C��L�#������t���5��伌��i���3�[���˿����=���꿇\��"Q�ں������w���ך�pG���&d���/���d?��p��bb�Md7�B����.��O9Ѿ+Gʾi�Ͼ ��� �,���v3���\�\R������+���U*�R^�/އ����� ���kS��w^��_(W�H�"��u����/ⰿǿ˽ �z�-�N(c��a�����Hi���{���ɂ�,�R�]��d��{��韄��TR��,�M�=@�� �ܾ(�;�ʾuԾ�}꾜����;�?��>n��@���t̿�J��B;���o�IΎ�k������l���tz��"E�a���ܿ?��?<��H�ֿ_@��1?��t�4�����ڝ�Y���Ku��	A�5&��~ӿ����b�t��D�l�!����C��O־O8˾a�̾�rھN�����5�(�EfM�������Vu⿿C�I�L�7#���������6��"���ui�E�3�����˿����"������\�#Q�����"����w���ך��G���&d���/���?���p��'cb��e7����2�&��R<Ѿ+JʾW�Ͼ���L	 �d��x3���\��  �  T��>���5ۿ��	�i�+��L��d�,m��b���F�=�!��A���������>������<(˿6���W*���M�qf��l���`�0F��$�^�kпgp�������p�0�M��_0�Y�����><��dc�L` �����$��7@���`�'��������l���X�h���I7�iRV���i��uk��qZ��:�Q,�0�俙������������p����ݿ����6�܇W��vj���j�l0Y�%;�4���~�i����&�����~d�z�C�~�'�K5������������o�t��gc-�TpJ���l�K􊿊᥿�e˿�W���2 �[nB��q^��gl�q�g��1Q���.����ѿg�������츚�U����������B���_���l�~�f�4(P�b�/�$��ۚ࿂����땿^�}�j�X�h�9�Yx��0�Q��B��Ni���\	�.���6�x5U��_y���������ۿ��	�A�+���L���d��m�Yb�f�F���!�A���������=������A'˿���:W*���M�f���l�S�`��F��$�3��jп!p������0�p���M��^0�z�����0:��<a�1_ �����$��6@���`�����S���Rl��MX�=���I7�HRV���i��uk��qZ��:�H,�(�俜�������ʔ���p����ݿ����6��W��vj�&�j��0Y�a;�t��V�����1'��M�F�d�ҐC�ڞ'��6���f������p�y��Rd-�$qJ�a�l����᥿,f˿�W��3 ��nB��q^�\hl���g�2Q�6�.�~���ѿY���x���Ź�����^��6����B���_�%�l���f�[(P���/�O��A������앿��}���X��9��y�(2�PT��u��ll��^	����V�6��6U��`y��  �  nd��ɰ���ѿ� �#�� o���"�N�%�&��a�ˣ���9����z���m����� ����¿t���^ ��&�� �����������M̿��ѩ�蘿�_��m�f�6D�Wx)����[��� ��#7��V�(�{��֐�����ٸ���ÿ�ؿ�A��Ow�@G�8�$��W$��n������׿�U�����r��q�G��G���>ҿ�;�~�u�#��n%�����\�����j�ۿ�ſ�����Z��Ⓙ?�� �Z��<:�^�"��L�����!'���@���b�)@��w떿������bʿ��� �l�&n��&�5�!�.O�����s�ǿ� 2����n���w������Y��=�J��@���y%�ʒ#������V�:�ӿ����*��p��������Ds�mO�=H1�����P��+�U�.�"YK��o�_���2Ϝ��c��]���^ѿ� �����n���"��%����`�$��f��p��F�z��m�������¿7s�J�w^ �Q&��� �������[�俎M̿���Щ��瘿�_����f�+5D�Xw)����7���� ��"7�ĲV��{�=֐����_���}�ÿ��ؿDA��&w�G��$��W$�un������׿�U�����r��q�i��u��(?ҿ�;�-~���#�o%�Ŀ��\�C�����ۿz�ſV���o[���Ⓙ���k�Z�_>:���"�:N�)���"'���@�w�b��@���떿:��5���ʿև�7 ���pn�&���!��O�����U�ǿg 3��m�n���w�^���MZ���=⿎��{���y%���#��H��%W�ӿ�����+�� ���~���uFs�O��I1�>��eR�--��.��ZK�.o������Ϝ��  �  vc翛l�W���忶�忰C�Sj�1��<Tؿ9y��/����y��j�a�d^E�
8=�.�I�}cj��f��.��fƿ3vܿ���2U�p迳��Vd���%B�1���Կ�ܻ�^����6��>�[�3�B��=��N��|q�������ţʿf;߿���E����t�[��d��꿺3�Aѿ�"���噿@~��V��U@��*?�K�R�7y����
ﳿ�ο��R�꿂��`<�+j��l���pG�[���ZͿ�Q�� ���sv�QQ���>�A���W�Tw����������t�ҿ���+	�X8�ʴ濤~�1�I.��k鿧V޿�>ɿBr��]s���o���L���=��nC���]�眄�]��Oi���ֿ����T�u��)?����դ�@a�K��xۿ��Ŀ����c䋿Kh�[�H�,=��kF�(�c��툿YC��j����gٿ�b�'l��鿝��_��VC��i���濿Sؿ�x������y����a��\E�o6=���I��aj��e��J-��^eƿ�uܿ4�迿T��o�o��$d�����A��0忟�Կ]ܻ�����6��1�[��B���=�SN�H{q�G���y��0�ʿ�:߿v������bt��濻c���꿆3��@ѿ�"���噿�?~��V��U@�#+?���R��y�?���Oﳿe�οL�Ώ������<翶j心m翲��H��࿜[Ϳ�R��� ��uv��Q��>�`A���W��w��e������Āҿ��g	뿔8����~忙��.�bl�PW޿c?ɿs��+t���o�#�L�B�=�9pC��]������]���i��bֿ��aU�ݩ鿖?�o��_���a뿸K迒yۿ��Ŀ؊��O勿-h�=�H�=��mF��c��D�����jhٿ�  �  -�%�u:"����E��3^���Ͽ����^����כ�������l���I��:-����#b��h���2��P��bu�Z����������������Կ5
���.����#�??%��!�i����߿����/���bv�Io�RV���栿>sʿ���ed�4"�5�%����5,�0L��2�H�ȿ�3�����S땿*0��s�`�r?��&�X�����#���;�c�\�B���擿�F��f��z�ƿ�ݿס���M��s�̠%��#��{�����k�Ͽj�������j@p���s�j/������0ڿ�!�@\�8�$�ѥ$����T�
���g�׿I�¿�Ա������Ώ���y�u�T�c�5�G �՟��J�O�*��E���h�n���㙿`����ݺ��wͿ�)濦����0!��&���������]Z���H������m�	~|�L���6v��\W꿼���P���%�8:"�i�����]鿕�Ͽ<������yכ������l�g�I��9-�4���`�g�+�2���P�jau��������\��<�����Կ
���"��z�#�-?%��!�C��.�߿]�� /���av��o��U��"栿�rʿl���d��"���%�Q���+��K������ȿh3��r��'땿	0��H�`�^?��&�+X�7��6�#�'�;�ם\�����擿�F���f���ƿYݿh���*N�t�$�%��#��{�����2�Ͽ1������Ap� �s�
0������Z1ڿ�!�e\�T�$��$����m�
��󿻉׿��¿sձ�s���.Ϗ��y���T��5�� �L���K���*�W�E���h�o��"䙿ն���ݺ�(xͿ*����_��r0!�V&���+�����^[���I������m��|�8���w��'X���Q��  �  �m�Ld��3K���)�c-�wLؿ	��`���0w��`S�x�4�����|�S������[���$�� �SN;� �Z����!e�����vx��Q��1���Q�ؒg���l�Ww^���@��}�@0�ل��J���!��r����5Կ��
���0���R�9�h�Pl��1]�0�@��H����(�ȿ'������Z�j�ղH�#�+�����\d���m���K��I�	)�JBE�s}f��+���ɠ��5Ŀ�����y���<�|�Z�DNk���i��V�T�4����ɓڿ�s�������̗��۳�e�lE�w�<��[�<�k�
i�&�T� c5����(W�R?���j��<]��$�^���>��v#������"#�������e/���1���O�O�r��玿gD��	�ҿ¶���%�Q�G�r�a�!�l�]'e�B	L�Z9(���Fȿ�'�����	Y����¿�����#�NmH�U"c�Wm�d��3K�Y�)�6-�Lؿ�������1/w��_S�a�4�v���{�����[��.Y��#��� �#M;��Z�T���d�����Ix��Q��1���Q�Ԓg�w�l�@w^���@��}��/�A�������o�������4Կ)�
���0���R��h�l�p1]��@��H�K����ȿ�&��¬����j���H���+� �����d��Bn���K�@J�~	)��BE�~f�,���ɠ�G6ĿA���2z�5�<�ӐZ��Nk���i�_V���4�����ڿPt��w���͗�6ܳ��迨E���<�%�[�S�k�-
i�4�T�0c5����hW鿧?���j���]��G�^��>�Jx#�p������%�v���J���0���1���O�N�r�u莿�D����ҿ���%���G���a���l��'e��	L��9(����&Gȿ)��� ��Z����¿o��3�#��mH��"c��  �  8���1Ә�����d[�;�'�������tU��fZ���1�0Y�9��Mxྑ6Ͼ	Yʾk�Ѿ���`-���8j9��Be�����r¿KF�
�2��g�s��q��~T��,���a��� N�r�����'��%��Nο`H�sf6��l�F�������<ў��֓�Ӓ}��I�����޿�v����~�� K�B�&��v����Yپ\3̾9�˾�G׾*]�P
��p#�YF���w��h���׿�����C��x�	���6��ޞ��\��N�q�X><����#�ӿHe��k����߿,��
 H��A}����k�����������l��d8����tɿF���0k��=����^���辫�ӾM�ʾ6ξ:�ݾ�$������-��T�|��H���x��,"��U����fL�������p���)��/+`�`�*�eR��U�Ŀ4���)���@O���n%��*Z�&���������Ә����d[��'��������U���Z��1�'X�����u�4Ͼ�Vʾ��Ѿh��8,���Ki9��Ae�M����q¿>F��2��g�s��q��{T��!���a��� N�-����u��h��SMο�G�f6�fl��������ў�z֓���}���I����H�޿@v��c�~�B K���&�|v���� Zپ�3̾��˾�H׾�]��
�.q#��YF�Y�w�Si��e׿�����C�x�6���6����������q��><������ӿf���k��C�߿x��I H�(B}����t��
���������l��d8�����ɿ�����0k��=����_���A�Ӿ�ʾ�ξ��ݾ9'�� ���-��T��|���H��@y�+-"�n�U�����L��ֆ��7q��>*���+`���*��S��~�ĿV���@���IP��Vo%�+Z�Y�������  �  i7��٭��୦����ΨI�6��]qƿ������P�b�!����O�ܾ��¾�Y���c��O���Z~Ǿv��u���*� V^�=�����ֿ���%XX��?��Xˬ�����U��� ��dS��D5~�!a<�H	�?�׿TͿ�c��'#��_�	��>��������3���e������X�v��4�����dc����}�e�>����;����Ҿ~���I䱾�S����ƳϾӀ�r��[9�Yu�2���f��i�-��n�.��^���]r�����B�������Xkg�Z!)�xt��bϿE]Կj����5���v�wޜ�\����T���S��K���`��F�_��� ���߿yZ��Ơe��;/�������1ʾ��Б��ve�������YپQ- �ۤ�{~J��������p	��{B�����r��»�����������މ���KQ������ɐ˿е���8*J������������B7������ĭ��鹆���I���qƿ|�����P�x�!����,�ܾ��¾3W��Qa������|ǾV�侀��:�*�wU^� �����ֿ���)XX��?��_ˬ�����T��� ��PS��5~��`<��	���׿=SͿ�b�'#���_�O	�����k����3���e�������v�Ԉ4�B���c�� �}� �>���.;��k�Ҿ~���y䱾�S�������ϾŁ�,s�L\9��Yu��������-�b�n�I.�������r��?���v���ƶ���kg��!)�Uu��8Ͽ^Կƫ���5���v��ޜ�k����T���S��K���b��N�_��� ��߿�Z����e��</�����辔ʾ���H����g�����)\پk. ����J�I��4����	��{B�����r��J»����ĵ����)����LQ�C������˿��࿛���*J�ֽ����������  �  ����=��!���ED��x�c��Z�/�տ+	��V�O�|��o����/̾|
�������"���ʧ�#����Ӿ�� �F4%��P_�It���8��e,�@�t�9���������%l������\��KZ����T�����1�[���8�{j7��}�����C��ƛ��/���Y�������
����J���&���¸��"�;�D���徢G¾�l���}�������ҫ��U��P��,�ݞ5�Ƭy��������C����������N��a���,���%f���<���A��b>��a
����)鿘���M�K����i���%��^��������>��r2���}���3�f��W,��ãg��d*���w�׾����XL��'ڤ�5��,�Ⱦ���&���H��M��*�̿���][�-���UF��l������`O������t����l��M*�J����޿ƚ��0$���d��������T�������=�����-D��L�c��Z�֟տ�����O����~���-̾M��{���� ��rȧ��|����Ӿ�� ��3%�9P_�t���8��e,�J�t�A���������$l������\��.Z����T�t���0��࿉8�j7���}����eC���������2�������
����J���ԏ��������;�������pG¾�l���}��I���8ӫ�VV��D������5���y�3������C�����쀮�(O������`���Zf���<���A���b>�Gb
���������M�m��� j���%��f��������>��q2���}���3����,��{�g��e*�����׾7���~���N���ܤ����p�Ⱦ���'��H�AN����̿f��?^[�X����F����������O��9���5u��%�l�BN*�����L�޿����0$��d��������T���  