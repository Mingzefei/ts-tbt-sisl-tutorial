H   E���}H@                        m��b�@                        �%�J6;@H      �      �         �  f������������<	v�j�)�����h��%Q����������7?��u䚾m[��Q	���嬾��ɾ�����f#��b�,�������%9�fw��{���i���M������O�������6��;~e��#�Y���>���	@E��A��~γ�Z���c������M���`���o���8�Z��L�hĿ{ф���;�����ܾy����c��gi���ޘ�쬡��`��ū׾����5���~�H���C���R��Ԓ��/��s�����������)c���K��Fߍ�?�L��M�P�����\�\�zi���C��3����	��?����c��_���m����A�����j��6�l�1�*��?�jҾT��G���圾ß��J��D�ľ����TM�#���/�ؿA#�*�m�á�u��q���ok���6���)��#�������$�7�V��U�쿬O�=1�:x�HG��!T���*�������@��x���a����dw���*�«��"���V����a����d;���:�����������Թ��	׾Ʉ�k;*��h�ᨧ�4M��6�:�9Y��p��6���U���l�������Œ���I��˲g���%��|��P���szG�H]��T���#��Sz���������A���tǘ�u]�@e�	�ȿ���D�~3��7�$�Ⱦ՝��Ý��t���߱�a�žH��U���D=�px������Z��*2T���� >��8������6����v��n`��������N����t��h�����_��v��`F����������+k���@���:��wH���\C�yQ�W̯���s�=z1����n?߾֢������G訾_|��������Ͼ�q��t�_R������Yۿwi$��o��i��S���U��m��U�������ŏ��u��D�8�T���'�%{��<2��5y��٦���������  �  .���p����������k��D#�a�ڿg���K�P�`��c�u�ƾ~<��C���T���С��񱾕�ξ�����$�P�`����4>￲2���}���>o��He�����P���Y?�������1\��z���򿙽���	�0=�	����F��Y������-j��_���I��lA��<R��+�/���D��� <�%����᾵����H��+������K����~���ܾ��	���5�� |��<��
��ݵI�<����
��O��6u���f��,��Α��,���U�D����翛'�T���
T����w)��)1��ݒ��*��}������D���1":�~��G騿_#k���+��o���׾;#��#�������v��i?����ɾ�X��h���L��ݏ���ҿ�:��d��ۚ�����X�������Q��OT��\ף�w�v�D�0�^<�/�念����]*���m�?[�������/��)+������������1m��$�EMݿ;���=V�� �&�����Ҿ"�����6Y��v��྾,ܾ^���j+���g���������3�������&R��EK������%���FE���Ė�?c^�����[���9�X�	�?�l����`�������3��s��	#���[��vQ��7T�3D��ÿmg���[D���@5�Q�;���vH������-���H�ʾY�쾉����=��+��(]��"�
��K������,��Z���y���%������Q��3�F��D����ˋ����0V��(��e*��%���z���	�������{������;�s���J��Y�q�1x2���
��\侉�žt`��o���z0�����? վ�J������R�F{��k�տ����Re�����jg���M����������Z����n����w�R�1��c����Y�O�+� o�����9�������  �  .��������߬�����P�P�����ʿE����[Q�$� �L�L(ؾJ]��Ĝ�����)���Y¾<:ྖ'�y*��_�`֙�ܿ\Y���_�/����H��xD��:X����X������,�B�e���ܿ��ѿ,���QP(���g�P|��F�����������[U�����������:�P���ҳ��F���B?�Y/�	�.�ξb����լ��8��^���I˾���]Z��o9���w��������l3�y�w�kٞ�>����������j��<����o��i.������ӿ��ؿ_/���;���Iɢ��Ⱦ���������\s������h(h�tD&�m$�2���c�h���0�l_���~�ɾ�g���&���\��':����ھ���j ��uN��\���mĿI����I�J%�������F���	��_n�������'���Y�э�Ë��ѿ���y�#6R��A���̭������Z���y�������O��f�Q��1�;RͿ]��g�V��[&��������-ɾ챺���Ϩ��gFϾ<l���]�0��f�RS���߿i!�ѵa��b���)��-(���B��4 ���Y���˄���D��!�)���տ����r�*��#j�하������������i�������؀��<���������i���}G�`�Ƭ���޾`8Ⱦ�	��Fj��PƾÀ۾6-������A���uװ�9���5��y����μ�B���9"��^~���P��
�q���0�U�� m׿��ܿjW
��=�lɀ��ţ���������q����M��Ag���i�Z�'�x��
���o��g7�'�������?־j�þ�)�������̾M澐��n%�ٿS������ǿ.��IK�/͈�`���f������������w�����Z�T��7��WԿO�V@��[S�ь�iW��7O���  �  ���xt��x���� c�`�,�$�� U���ŋ���Z�q1��9��x�۾�*ʾ5žQ;J�ᾪz���V9���f��s���gƿD��Ə8��Do�A����<���L��{��#���UU�܋��F쿍����'��4�ҿ&��<�L�t��*��e����Ƥ�W��~h��+�P�R�1俪E�������K��s&��\����Xվ��Ǿ~ǾiӾ�������"���F���y�ۢ� ܿ���m�J��{��VE������x���^����z�EB����0ؿ�H��a���	�S#�@O��S��8����������y!��īu��>�n/�A"ο(♿�n�/�?�B,����e龳�Ӿ��ʾ��ξ�O߾����c��1�0�_Y�򠉿,��@���(���]��U���X���������굎�&i�܌1�Y���ʿ�̵�i�ƿ<�����+��c�97���f���:��\%���2��Kad�R3.�?���H��Y���e`��6����-��q�羢@־Q�Ѿ3�پ)����p���*@��m�C񗿙�ɿ��	��N:��q�{s��/��=4��Al��n���cW�M�!�������J���6>׿S[�!�>���v��B��7���ܥ��j��yz��[�R�_n�]3迩o��W����T��.����4�������ؾ�B׾�P㾈��p��!�*���N�l��p���D&���ԢL�6���U���$�����r����|��D����Ʌܿ����^վ��F�7��Q�K��B������f������[w��@�����ѿsD���Bu�-$F�~�$��S�-���ྺ�־�mھ��꾴��;��6��a^��>��+Ʒ�Z����l)��$_�{������-���xP��JV��^j��2�F��EͿ��Aɿ" ���,�v"d�����"���  �  [yu���k�`R�N!/�����ܿ�ϱ��H����x�8T��4�*�������������1�
��  �\;�H�[�62���]��jF�����j�_O7��Y���o��u�gf��zG�_a �A���0���᛿ �� ����>ٿ����6��LZ���p�ԝt�:e�� G�/*#�yW��%Ϳ����wK��Iil��~I�6�+���LW���M��� �uL�Ϸ(�I�E��h����i���ȿӿ����a%C�%b���s��/r�8v]�!�:���a�߿�A��8Ŗ�����5�����C�!�c�Ѭt��q��\�*�;�R��ռ�����dX���x����a���@���$�f�cz ��t��Q���F$�J=���4� �S��x��L��,Ư�Eٿ+(	��,��hO���j�)\v��An�,T�!�.�M��F�ο��������ޢ�+ɿΤ�h*���P��}l���v�|am�QqS�;�0�T4��߿������4x~�A�Y�^:��e ����r� �3��b �<&���&�lB��b�.����ۜ��ǽ�G�|(��9���Z�ޖq�_�v��Bh�=jI��c"�����n��1��R^��T���d�ݿ�(���8��{\��s�F�v��-g��DI�QJ%��s��Vѿ�몿�n���t�4�Q��3�T���s
��'�!� �����g���0�K�M�N4p�����<���(̿���@)!��AE�MDd���u��St�˛_���<��A����싲�m	������^���!�� ��iE�L�e��lv��ps�oO^��g=�aZ�� �k�¿�����ԇ��Wh� GG�C[+�xZ����
< ���o���� ��V:�(Y�)k}�Dꔿ�_��:�ۿ#w
�QY-���P�rl�Q�w�2�o��XU���/����Lѿ���i���*��ML˿Q��0}+��Q�K�m��  �  �+��-'�����5�(��n�ӿ��,E��Y��u��!�n�J���,�r��)�,z��|2���Q�7�w�p��� !��?���1Ŀ Tٿ����R����)��*����-���4��j#��˓x�H�p�iՅ�⫣��&Ͽ�� ����5O'��<+��#��U��o�忑�̿R���h����+�����eb�S�?�_�%�X�����;s#��1<�"^�y��������"�����ʿV���f �M@�C-"���*��4(�����c�'OԿڪ��5&����q�7�u�����X󰿪�߿'	�Kc��B*��6*���Ի�c8����ܿ]ǿ�
���)����~���W���7���!�;�|�I-��zI���m�!���0ԝ�=F��t �� Uӿ$'��*����
'�D;,�I�%� �g	��%xƿ����#e���s������$������������$��,�Đ(��?�N�	��V񿝢ֿ�¿9���Π��獿�nt���O�O�2�� �\U���#��8�y[X�E~��񒿽�������K�ǿi�ܿ9E����&<��*�O,�G�!�����%�Q���EM�����4�y��)�����$�ӿ���b�7{)�@f-���%�ly����uT鿑)ѿ%¾�����H��yڈ��j�[�G���-�ɤ�����+�kLD��:f�`������`��4���h�οL���R\�L$���,��W*���,����ؿv﫿�d���Iz��!~�����(���/ ���+�/�+�>!�Wj�����dK�{ʿ"��~S�����C��pZ^�;#>���'���L�!�H�2�uO��@s��Y��{���㱿��¿P�տ\��Z|��J�_(��-�`�&�qg�\�����ȿP��k���cx��܃��b��U�ÿ
���-����%��  �  b��2��N��� �̎���m�,TݿNwĿ�`��
��}�b�ÛE�^+=�TnJ� l��C��!H��#�ʿƻ�^j�Y�������b�	���(�ٿwӿ��r���Ą�h]�nC�q2>�� O���s��4��Ɖ���LϿ����I���D�%���?���d�����'6ֿ����u��я���`W���@���?�T�S���{�'��抷�dmӿ^6�e?�?��q쿧t���Q�H��<;���ѿ����q:���x���Q�b�>��WA��CY�����]��������׿�-��񿔑��쿉q뿵*�آ�=��0����ο���Ő��Gcs�z�O�$C@��mF�{�a�Y���O���R�¿��ܿ;%� ����1�ē쿴�������ۃ⿈˿����_�����m� oM��}A��BK�^�i����哪�\�ȿ�ῢ�ￖ��G񿦟�2��D����&�Q�XFǿ�>������4�h��K��UC���P��r�����ݛ��q!οD0�p��"����S�C�/��_����i�(�ݿ��ÿ�S����G6e��^K�ĪF�x�W��m|�R����඿ʣӿ�U��#����w���w�C��������
Sڿq������)����|_��H���G���[�$؁�^!������A�׿�P�,_��e��M������)���f$��~�"ֿ�z������Z8Z��G�߅I��Ha������)������E�ۿ���������{ ���9���
�� b������ѿ����\���g�y�\�U��CF�ETL��{g�%u��Qc��h�ſ�p߿F��ei��!�`��@5�*j�6u��'h��!�"�Ϳ���|,����r�+*R��!F���O��En�[$��i���%�ʿ���  �  n ��R����+տ#P�+7	�F����'�]+�ao"�7k�[��Ϳ�������|��{o�7E���{��
ǿi����a�j%�{\+��%�q)�Q�m�鿅dп�U��ϫ��z/��"���şh���D�o1)�������s �Qa7��X�`v~��䒿�.�����rǿ��ݿ�_��c�9 �	4*�	�)��1�v����ܿ!�������?�t�?s�5������/F׿������(���*��{!�I������P��[ɿ����Qئ��Ô�93��:�[�j?:�b-"��P���'�Y�A�e��A��ⴙ�Zz���-����οa]�������3�$���+��'�4����]xͿ"����ƅ���r�b~|����LZ��Ew�Z���!�o�+��)�����.�������ٿb�Ŀ�鳿�cQ��"@y���S��)5��� ����*����2�&�P��u�ǎ�E����Ჿ��ÿ�׿�󿦓
��"��)�,e,���#���f�c���=�� z��]�u�d������DʿI4�����"'��-�%X'����G��D��ӿ<����8��О�X���kHp�}�L�sA1��-!��J���(�
�?��`�]���M7������C���˿���]����~�\"��H,�N�+�E@�1�	�F��J���}���}��{�>������,Uۿ����(���*�H�,�(�#��^�������d�ͿrȻ����=���p���*d�g�B��|*���� �@�.��tI���l��䉿a>��﮿����.ҿT���q��X��n&��b-���(�����h�q�п:ƥ��ш���x��4������w7���D쿎�	�"���,��*���0|��Z���Zܿ��ǿ܎������?撿�P~�L�X�?:��%��)��;$��@7�jU�!z��ѐ������  �  I���\ɳ���߿h��)1���S��m�uu�ej�`M�E�&�}y ���ÿE��O ��=+��L�Ͽe����/�c�T�[On��Vu�2�h���L��%)����/�Կ�)��=����r���N��I0��)���M��%��$�����y$�ض@��b�����M>�����3�cC��]=�d�]�	r��s��>b��MA�S���w����9��s���򖰿[X��d�n=��'_���r��6s���`�F8A��pk����ſFN��,.���e���C���&�1��? �-����[��I�T�-�/#L�Ïo��5���3���_пg�A�%�B^I�R�f�iLu��p��Y��4�-]�׿i穿�֖�@6���������M#��?J�~h�*v��o��5X��)6��a���翪߹�W����Ӂ�?�]��=�m�"����� �����G�����+� �rT;� [��B��fm��0�����}�V�2�.U��an���v��pk�Q�N�2l(�����ƿ�Q�����xE���ҿ1
�v�1�r�V��p�Pw��j�ExN���*�A�lUؿj����Ȓ���y��/V�z�7����^����NC ��E���O-��MI�R�j��>��劢��_ſ�v��<b�-y?�E�_�g-t�v��Ld�<YC����҇���#�� ���Ѣ��@e�Dl�.?��2a�w�t�Fu���b�kMC� .�<���R�ɿ�����j��&n��-L�q_/��H�=�Jg �mg��(�b���c5�.[S�6�v�����/�����ӿ@�5'��K�3`h�j�v�K1r���Z�On6�����*ڿ���ՙ��.��t�¿m���Ÿ$���K�s�i��gw�U#q�4�Y�w7����$&�����?���r��P�b�x�B�#�'���Q�Ff �>_�}���%�v�?�B*_��A���  �  _ƍ��i��r� �1�/��f��͌��4��U���j���(@��_�^���'�^��� �¿ĳ� ˿�5��s3��Ak��~���ܠ�K]��?��䌇�]�Y�v$��@�ۋ������4S�<�+�$1������ؾ�ɾ�Bƾ�@о?��2����@�5p�x����ѿ�T��A�xMx�������?���䠘�Ӂ���K�^��a��9����s��o~ۿs��E�ì}�z�����P����?���~�0�G��N��"ؿ^7���Hv�G1D�h� �&C������Ѿ��ƾȾ׾]�tZ��)� RO����0������l]��)T�����w���5��aH��}5���r��:�`	�=Vѿҵ�8g���:��"��)Y�`������|ڥ��	���ʏ��m��{6��g�e�ĿL��CDg���:��]�gZ��i��Ծ.ξ%�ӾT�����~��68�{�b�b���M-���1��1��mg�?{��2��=��-�������U+`��Q)�H���-�ſLֶ�$ο���5���l��Q�������:������l��C�[��3&����q��s����hZ��3�}��.��x�\6پ'�־��ྚ���7��Ŕ&��H���x��ԟ��Hտv�R�C��hz��%���������֧���؂�I N�D�����`�����*�߿jy�6�G�_������V���ä��H��P����I��h�Zܿ�p���~���L�`O)�E���K���F⾬�־[ؾi��� �ض��H0��VV��j��`���!�,�U��Յ��P�����������s�Ԕ;���
��WԿiи�(cÿ2��	h$�N�Z�����mo��σ�������p���in���7���_tǿ������l�$@�7t ��V	�(��]޾�E׾[ݾLz�1Q�����F<�O�f��  �  �<����ο����QT�̙��8�������T����.������ƭ���dM��T��4�}�Ͽ�^��O��T\�������������p�����ק�ƹ���jE��$
��վ�|8��H�o������kӾ�ƺ�$ۭ�菫�����q�ƾ�;��J���1�.Yk�����<��A)�1�k�K������U��!���x�����U�{��l8�� �V׿��Կx���1��s�N0���ֺ������g���r�����g�s�A�/����cF��s��}6�\Z��1��ɾ�0��$ ��	�������TѾ�������>C�W)�����w��|�>����S���䶿��3�����g���ϕ���d�,�%��7��	ҿq�߿���k�F�����u��.���C������}+������
�\�B�QQٿ����_�3a+��p	�[�Pɾ�Cg��@U���Ⱦ$����~'(�TZ�������ѿd<�f�U�I���2��7i��g^������=���m����N�����G���ҿo�� ���]�2f���߲�����K������������'G����U¿@��@O��5"�,�����>wʾ)߽�&߻��MľZ�׾�)��m���<:�F�s�KV���b+�F�m��X���Ÿ��_��k������u�����}��t:��'�bۿ`�ؿG��c�3��u��4���ۻ�ǣ��o��h{�������u��2����	~���{{�`�>���$���<�پ�pžm���K���ɾ�V�i���%�,?J�̙��@{������4@��ʂ��_���������S��2��q���"f��Z'�K4���տ����u��`H��̆��+��98���������Ҳ�=���>C^��Y�|�ۿ_^��)�d���0�'���Ӿ�o¾N����W���о�d�D���6,��^��  �  `��v}߿o�&��Cp�8�����u���[|��pp���&��I�����h�X*&�Z���������3�>�y�+���P��������>�����DW��� ����^����p�̿!S��F�������]¾@ܪ�l���휾\��[d����վ*s�e-��n�x׫�z ��=��Å���̂��9���o���������ߎ��=P��|�����N����R�H�^Q�� ˲����
������a�������L��	�E�+���4��?w��h2�4����پ�ո����݂�����4���>m����� ���x@�0����Ŀy���V�V���,�������v�������p���V��ɣ���:�m�9�Ո��U� ���`�fN��Κ��%w��x�������\���3���)z�Z%/�#���r��R.`�S�%�D�`�Ծ�����Ʃ��Τ��K���շ���Ҿ~���"���Y��Ǚ��A��9(�_�q�$������_2���.��(��G����B���j�1�'����z��Op�s�4��V{��X��mq��8j���������4�������`�i���п<܎�w5M�T`������Ѿ�}���򮾱,��Lݴ�ǾM������5�ծv����(���?��҆�=���\���	����������e��G���ER�������*Z�×���J��T��5ϳ����� ��=���&������DX��&�G����k��x���:�L���?ɾ��q������E���aϾݒ��m��vG��򉿶�ǿHj�ZX�e���
]���s��4����^��8�����@c��><���	�(�C���m"��hb����S��/)���[����������?ܦ�[|{��x0��R���^le���*��[�&�޾4�¾J��Z���L��:���2۾�e��&�ڬ]��  �  ����$��R-���z��q������ϰ�����]������R���wr���,������?��8:��D���ˬ�h���*�������R����������Vh���s.ҿ�J��#F�HT���k7���꥾�L���I��i����N��.�оFM��,��p�[���gG�!wE���������-���g'��	����?�����"��>�X����Z��!�������P�dO����������l���l���7������l����M��_
��U���iy�}�1�N����Ծ����q蠾i☾b8������M��S�	��M@��2��/�ɿ��_�NP��z���cz��N������������ű��7��NB�M��m����8"'��gj�l������D���4��0��Z:����������	6����Qc��6Ia�gq$�����T�Ͼ�ﳾk��^.��
���7ղ��;m���D� ��oZ�K_��p��e�.��|�%"�����Ka��>���`���v��4��t�U@.�?(�}���
�ļ;�6������MZ��r�������'������lȟ��j�c �A�տӐ��PM�ۤ����}̾k����;��a�������¾���L�
�ר4���x�gӳ��i���G�����D���� ��-1��4���XF��#������Z��$�}f��z��������R��R��ۡ������r��t���@��6��#x����O�]z����bꀿ6#:���a�徙#ľP��'̨�Lթ�o\���=ʾ��ﾌ+��JG�i�����̿���cka��%�������N��S�������L������=���D�C�����j��� �ڤ(���k�����T������� �����������K��y/��0]7��������8�f���)���^�پ���������p���������
־����$��k^��  �  `��v}߿o�&��Cp�8�����u���[|��pp���&��I�����h�X*&�Z���������3�>�y�+���P��������>�����DW��� ����^����p�̿!S��F�������]¾@ܪ�l���휾\��[d����վ*s�e-��n�x׫�z ��=��Å���̂��9���o���������ߎ��=P��|�����N����R�H�^Q�� ˲����
������a�������L��	�E�+���4��?w��h2�4����پ�ո����݂�� ���4���=m����� ���x@�/����Ŀy���V�V���,�������v�������p���V��ɣ���:�m�9�Ո��U� ���`�fN��Κ��%w��x�������\���3���)z�Z%/�#���r��R.`�S�%�D�a�Ծ�����Ʃ��Τ��K���շ���Ҿ~���"���Y��Ǚ��A��9(�_�q�$������_2���.��(��G����B���j�1�'����z��Op�s�4��V{��X��mq��8j���������4�������`�j���п<܎�w5M�U`������Ѿ�}���򮾱,��Lݴ�ǾN������5�ծv����(���?��҆�=���\���	����������e��G���ER�������*Z�×���J��T��5ϳ����� ��=���&������DX��&�G����k��x���:�L���?ɾ��q������E���aϾݒ��m��vG��򉿶�ǿHj�ZX�e���
]���s��4����^��8�����@c��><���	�(�C���m"��hb����S��/)���[����������?ܦ�[|{��x0��R���^le���*��[�&�޾4�¾J��Z���L��:���2۾�e��&�ڬ]��  �  �<����ο����QT�̙��8�������T����.������ƭ���dM��T��4�}�Ͽ�^��O��T\�������������p�����ק�ƹ���jE��$
��վ�|8��H�o������kӾ�ƺ�$ۭ�菫�����q�ƾ�;��J���1�.Yk�����<��A)�1�k�K������U��!���x�����U�{��l8�� �V׿��Կx���1��s�N0���ֺ������g���r�����g�s�A�/����cF��s��}6�\Z��1� �ɾ�0��$ ���������TѾ�������>C�W)�����w��|�>����S���䶿��3�����g���ϕ���d�,�%��7��	ҿq�߿���k�F�����u��.���D������}+�������\�B�RQٿ����_�4a+��p	�\�Pɾ�Cg��@U���Ⱦ#����}'(�SZ�������ѿd<�f�U�I���2��7i��g^������=���m����N�����G���ҿo�� ���]�2f���߲�����K������������'G����U¿A��@O��5"�-�����?wʾ*߽�&߻��Mľ[�׾�)��m���<:�F�s�KV���b+�F�m��X���Ÿ��_��k������u�����}��t:��'�bۿ`�ؿG��c�3��u��4���ۻ�ǣ��o��h{�������u��2����	~���{{�`�>���$���<�پ�pžm���K���ɾ�V�i���%�,?J�̙��@{������4@��ʂ��_���������S��2��q���"f��Z'�K4���տ����u��`H��̆��+��98���������Ҳ�=���>C^��Y�|�ۿ_^��)�d���0�'���Ӿ�o¾N����W���о�d�D���6,��^��  �  _ƍ��i��r� �1�/��f��͌��4��U���j���(@��_�^���'�^��� �¿ĳ� ˿�5��s3��Ak��~���ܠ�K]��?��䌇�]�Y�v$��@�ۋ������4S�<�+�$1������ؾ�ɾ�Bƾ�@о?��2����@�5p�x����ѿ�T��A�xMx�������?���䠘�Ӂ���K�^��a��9����s��o~ۿs��E�ì}�z�����P����?���~�0�G��N��"ؿ^7���Hv�F1D�h� �&C������Ѿ��ƾ��Ⱦ׾]�sZ��)�RO����/������l]��)T�����w���5��aH��}5���r��:�`	�=Vѿҵ�8g���:��"��)Y�`������|ڥ��	���ʏ��m��{6��g�f�ĿM��DDg���:��]�gZ��i��Ծ.ξ%�ӾS�����~��68�z�b�a���L-���1��1��mg�?{��2��=��-�������U+`��Q)�G���-�ſLֶ�$ο���5���l��Q�������:������l��D�[��3&����r��t����hZ��3�~��.��x�]6پ(�־��ྚ���7��Ŕ&��H���x��ԟ��Hտv�R�C��hz��%���������֧���؂�I N�D�����`�����*�߿jy�6�G�_������V���ä��H��P����I��h�Zܿ�p���~���L�`O)�E���K���F⾬�־[ؾi��� �ض��H0��VV��j��`���!�,�U��Յ��P�����������s�Ԕ;���
��WԿiи�(cÿ2��	h$�N�Z�����mo��σ�������p���in���7���_tǿ������l�$@�7t ��V	�(��]޾�E׾[ݾLz�1Q�����F<�O�f��  �  I���\ɳ���߿h��)1���S��m�uu�ej�`M�E�&�}y ���ÿE��O ��=+��L�Ͽe����/�c�T�[On��Vu�2�h���L��%)����/�Կ�)��=����r���N��I0��)���M��%��$�����y$�ض@��b�����M>�����3�cC��]=�d�]�	r��s��>b��MA�S���w����9��s���򖰿[X��d�n=��'_���r��6s���`�F8A��pk����ſFN��,.���e���C���&�1��? �-����[��I�R�-�-#L���o��5���3���_пg�@�%�A^I�R�f�hLu��p��Y��4�-]�׿i穿�֖�@6���������M#��?J�~h�*v��o��5X��)6��a���翫߹�X����Ӂ�A�]��=�n�"����� �����F�����*� �qT;��[��B��em��/�����|�U�2�.U��an���v��pk�Q�N�2l(�����ƿ�Q�����xE���ҿ1
�w�1�r�V��p�Qw��j�FxN���*�A�mUؿk����Ȓ���y��/V�{�7����_����NC ��E���O-��MI�R�j��>��劢��_ſ�v��<b�-y?�E�_�g-t�v��Ld�<YC����҇���#�� ���Ѣ��@e�Dl�.?��2a�w�t�Fu���b�kMC� .�<���R�ɿ�����j��&n��-L�q_/��H�=�Jg �mg��(�b���c5�.[S�6�v�����/�����ӿ@�5'��K�3`h�j�v�K1r���Z�On6�����*ڿ���ՙ��.��t�¿m���Ÿ$���K�s�i��gw�U#q�4�Y�w7����$&�����?���r��P�b�x�B�#�'���Q�Ff �>_�}���%�v�?�B*_��A���  �  n ��R����+տ#P�+7	�F����'�]+�ao"�7k�[��Ϳ�������|��{o�7E���{��
ǿi����a�j%�{\+��%�q)�Q�m�鿅dп�U��ϫ��z/��"���şh���D�o1)�������s �Qa7��X�`v~��䒿�.�����rǿ��ݿ�_��c�9 �	4*�	�)��1�v����ܿ!�������?�t�?s�5������/F׿������(���*��{!�I������P��[ɿ����Qئ��Ô�93��:�[�j?:�b-"��P���'�X�A�e��A��ᴙ�Yz���-����ο`]�������2�$���+��'�4����\xͿ!����ƅ���r�c~|����LZ��Fw�[���!�o�+��)�����.�������ٿc�Ŀ�鳿�dQ��$@y���S��)5��� ����*����2�%�P��u�ǎ�D����Ჿ��ÿ�׿�󿥓
��"��)�,e,���#���f�b���<�� z��]�u�d������DʿJ4�����"'��-�&X'����H��D��ӿ=����8��О�Y���lHp�~�L�tA1��-!��J���(�
�?��`�]���M7������C���˿���]����~�\"��H,�N�+�E@�1�	�F��J���}���}��{�>������,Uۿ����(���*�H�,�(�#��^�������d�ͿrȻ����=���p���*d�g�B��|*���� �@�.��tI���l��䉿a>��﮿����.ҿT���q��X��n&��b-���(�����h�q�п:ƥ��ш���x��4������w7���D쿎�	�"���,��*���0|��Z���Zܿ��ǿ܎������?撿�P~�L�X�?:��%��)��;$��@7�jU�!z��ѐ������  �  b��2��N��� �̎���m�,TݿNwĿ�`��
��}�b�ÛE�^+=�TnJ� l��C��!H��#�ʿƻ�^j�Y�������b�	���(�ٿwӿ��r���Ą�h]�nC�q2>�� O���s��4��Ɖ���LϿ����I���D�%���?���d�����'6ֿ����u��я���`W���@���?�T�S���{�'��抷�dmӿ^6�e?�?��q쿧t���Q�H��<;���ѿ����q:���x���Q�b�>��WA��CY�����]��������׿�-�
�񿒑�	�쿈q뿴*�֢�<��/����ο���Ő��Fcs�z�O�$C@��mF�|�a�Y���P���S�¿��ܿ<%�����1�œ쿵�������܃⿉˿����`�����m� oM��}A��BK�]�i� ���䓪�\�ȿ�ῠ�ￕ��F񿤟�1��D����&�P�WFǿ�>������3�h��K��UC���P��r�����ޛ��r!οE0�q��#����S�C�1��`����i�)�ݿ��ÿ�S����H6e��^K�ĪF�x�W��m|�R����඿ʣӿ�U��#����w���w�C��������
Sڿq������)����|_��H���G���[�$؁�^!������A�׿�P�,_��e��M������)���f$��~�"ֿ�z������Z8Z��G�߅I��Ha������)������E�ۿ���������{ ���9���
�� b������ѿ����\���g�y�\�U��CF�ETL��{g�%u��Qc��h�ſ�p߿F��ei��!�`��@5�*j�6u��'h��!�"�Ϳ���|,����r�+*R��!F���O��En�[$��i���%�ʿ���  �  �+��-'�����5�(��n�ӿ��,E��Y��u��!�n�J���,�r��)�,z��|2���Q�7�w�p��� !��?���1Ŀ Tٿ����R����)��*����-���4��j#��˓x�H�p�iՅ�⫣��&Ͽ�� ����5O'��<+��#��U��o�忑�̿R���h����+�����eb�S�?�_�%�X�����;s#��1<�"^�y��������"�����ʿV���f �M@�C-"���*��4(�����c�'OԿڪ��5&����q�6�u�����X󰿩�߿'	�Kc��B*��6*���ӻ�a8����ܿ\ǿ��	���(����~���W���7���!�;�|�J-��zI���m�"���1ԝ�>F��u ��Uӿ%'��*�����
'�E;,�I�%� �h	��&xƿ����#e���s������$������������$��,�Ð(��?�M�	��V񿜢ֿ�¿8���Π��獿�nt���O�O�2�� �\U���#� �8�z[X��E~��񒿾������L�ǿj�ܿ;E����'<��*�O,�H�!�����%�Q���EM�����4�y��)�����$�ӿ���b�7{)�@f-���%�ly����uT鿑)ѿ%¾�����H��yڈ��j�[�G���-�ɤ�����+�kLD��:f�`������`��4���h�οL���R\�L$���,��W*���,����ؿv﫿�d���Iz��!~�����(���/ ���+�/�+�>!�Wj�����dK�{ʿ"��~S�����C��pZ^�;#>���'���L�!�H�2�uO��@s��Y��{���㱿��¿P�տ\��Z|��J�_(��-�`�&�qg�\�����ȿP��k���cx��܃��b��U�ÿ
���-����%��  �  [yu���k�`R�N!/�����ܿ�ϱ��H����x�8T��4�*�������������1�
��  �\;�H�[�62���]��jF�����j�_O7��Y���o��u�gf��zG�_a �A���0���᛿ �� ����>ٿ����6��LZ���p�ԝt�:e�� G�/*#�yW��%Ϳ����wK��Iil��~I�6�+���LW���M��� �uL�Ϸ(�I�E��h����i���ȿԿ����a%C�%b���s��/r�8v]�!�:���a�߿�A��8Ŗ�����5�����C�!�c�Ѭt��q��\�*�;�Q��Լ�����cX���x����a���@���$�e�cz ��t��Q���F$�K=���4�"�S��x��L��-Ư�Eٿ,(	��,��hO���j�*\v��An�,T�!�.�M��G�ο��������ޢ�+ɿΤ�h*���P��}l���v�{am�QqS�:�0�S4��߿������2x~�?�Y�^:��e ����q� �3��c �<&���&�mB��b�/����ۜ��ǽ�G�}(��9���Z�ޖq�`�v��Bh�>jI��c"�����n��1��S^��T���d�ݿ�(���8��{\��s�F�v��-g��DI�QJ%��s��Vѿ�몿�n���t�4�Q��3�T���s
��'�!� �����g���0�K�M�N4p�����<���(̿���@)!��AE�MDd���u��St�˛_���<��A����싲�m	������^���!�� ��iE�L�e��lv��ps�oO^��g=�aZ�� �k�¿�����ԇ��Wh� GG�C[+�xZ����
< ���o���� ��V:�(Y�)k}�Dꔿ�_��:�ۿ#w
�QY-���P�rl�Q�w�2�o��XU���/����Lѿ���i���*��ML˿Q��0}+��Q�K�m��  �  ���xt��x���� c�`�,�$�� U���ŋ���Z�q1��9��x�۾�*ʾ5žQ;J�ᾪz���V9���f��s���gƿD��Ə8��Do�A����<���L��{��#���UU�܋��F쿍����'��4�ҿ&��<�L�t��*��e����Ƥ�W��~h��+�P�R�1俪E�������K��s&��\����Xվ��Ǿ~ǾiӾ�������"���F���y�ۢ� ܿ���m�J��{��VE������x���^����z�EB����0ؿ�H��a���	�S#�?O��S��8����������x!��īu��>�n/�@"ο'♿�n�.�?�A,����e龲�Ӿ��ʾ��ξ�O߾����d��2�0�`Y�󠉿,��@���(���]��U���X���������굎�&i�܌1�Y���ʿ�̵�i�ƿ<�����+��c�97���f���:��\%���2��Kad�R3.�?���G��X���e`��6����,��p�羡@־Q�Ѿ3�پ*����q���*@��m�D񗿚�ɿ��	��N:��q�{s��0��>4��Al��n���cW�M�!�������J���6>׿S[�!�>���v��B��7���ܥ��j��yz��[�R�_n�]3迩o��W����T��.����4�������ؾ�B׾�P㾈��p��!�*���N�l��p���D&���ԢL�6���U���$�����r����|��D����Ʌܿ����^վ��F�7��Q�K��B������f������[w��@�����ѿsD���Bu�-$F�~�$��S�-���ྺ�־�mھ��꾴��;��6��a^��>��+Ʒ�Z����l)��$_�{������-���xP��JV��^j��2�F��EͿ��Aɿ" ���,�v"d�����"���  �  .��������߬�����P�P�����ʿE����[Q�$� �L�L(ؾJ]��Ĝ�����)���Y¾<:ྖ'�y*��_�`֙�ܿ\Y���_�/����H��xD��:X����X������,�B�e���ܿ��ѿ,���QP(���g�P|��F�����������[U�����������:�P���ҳ��F���B?�Y/�	�.�ξb����լ��8��^���I˾���]Z��o9���w��������l3�y�w�kٞ�>����������j��<����o��i.������ӿ��ؿ_/���;���Iɢ��Ⱦ���������\s������h(h�tD&�l$�1���b�h���0�l_���~�ɾ�g���&���\��(:����ھ���k ��uN��\���mĿI����I�J%�������F���	��_n�������'���Y�ҍ�Ë��ѿ���y�#6R��A���̭������Z���y�������O��f�Q��1�:RͿ]��f�V��[&��������-ɾ챺���Ϩ��hFϾ=l���^�0��f�RS���߿i!�ҵa��b���)��-(���B��4 ���Y���˄���D��!�)���տ����r�*��#j�하������������i�������؀��<���������i���}G�`�Ƭ���޾`8Ⱦ�	��Fj��PƾÀ۾6-������A���uװ�9���5��y����μ�B���9"��^~���P��
�q���0�U�� m׿��ܿjW
��=�lɀ��ţ���������q����M��Ag���i�Z�'�x��
���o��g7�'�������?־j�þ�)�������̾M澐��n%�ٿS������ǿ.��IK�/͈�`���f������������w�����Z�T��7��WԿO�V@��[S�ь�iW��7O���  �  .���p����������k��D#�a�ڿg���K�P�`��c�u�ƾ~<��C���T���С��񱾕�ξ�����$�P�`����4>￲2���}���>o��He�����P���Y?�������1\��z���򿙽���	�0=�	����F��Y������-j��_���I��lA��<R��+�/���D��� <�%����᾵����H��+������K����~���ܾ��	���5�� |��<��
��ݵI�<����
��O��6u���f��,��Α��,���U�D����翛'�T���
T����w)��)1��ݒ��*��|������D���1":�}��G騿^#k���+��o���׾;#��#�������v��i?����ɾ�X��h���L��ݏ���ҿ�:��d��ۚ�����X�������Q��OT��\ף�w�v�D�0�^<�/�念����]*���m�?[�������/��)+������������1m��$�EMݿ;���=V�� �%�����Ҿ"�����6Y��v��྾,ܾ^���j+���g���������3�������&R��EK������%���FE���Ė�?c^�����[���9�X�	�?�l����`�������3��s��	#���[��vQ��7T�3D��ÿmg���[D���@5�Q�;���vH������-���H�ʾY�쾉����=��+��(]��"�
��K������,��Z���y���%������Q��3�F��D����ˋ����0V��(��e*��%���z���	�������{������;�s���J��Y�q�1x2���
��\侉�žt`��o���z0�����? վ�J������R�F{��k�տ����Re�����jg���M����������Z����n����w�R�1��c����Y�O�+� o�����9�������  �  ~i��5_������넟��_l�C/#�r`ٿ6��Z�K���Z�羭��+��"�����|:��d���z�ž�c�����=)\��>��.=�A2��~������H���U����������ѽ�q����\�-��9�򿵰��	���=�����Ĭ���������Y������f�������nR��������(���L7�����ؾ)���r�������,��kƞ�+���iӾ���0�0���w�󩵿����I��	���µ�����e���A��-������3Q����D�-�ω��$�urT��{�����������t��:�������J��h���@:��)���.��V�f���&����seξ�Ѱ��q��N8��Q��|C���
��V�辎v�HH��ݍ��ѿ���}d��f��]�������������������J��w��1��G�l��O�����*��rn�#ɟ��I��y���;�����Ś��t3����m���$��ܿ<Ŕ��aQ�����9�ɾ����6��;
���ߦ�䢶��Ӿp� �{&�c���������3�!��S����+���;�� �������׾��(���^�G��r]��<,�1�:@�	���ޭ�����`
���n������j˒���T���D¿uK���?��+����/[ž�����禾Q]������5¾��G�m�8����ɹ��
�yL�p���ж�a���v��	T������~)��%g��%G��]�h����Z:��V��������������\�����������%���߄��;�����\���d]m�:�-�Z�9۾�b��8����9��󾨾
����8̾������^M��{���8Կa�w�e�����1���:���n��Q���������6;x��-2�(o�.���#�f�+�@�o� [������ۀ���  �  �L��G���?c�������b��2�Rӿ[���Y[K�
��l�3%þ4	�������3��^䞾����I�ʾ6����� �^�Z��G��.翧Q+��s�g��o���s��t����6��ֵ��ӏ���S�����K�޿ 0�Xb6���|�l���f������{D��ב��d��������I��
���`���7���
��_ݾ���:���C������녣������Sؾ��$Y1�k\u�·�����w�A�[����޻��Y���T������@���?���U/=��-	�B`�i�濼��4�K�\m��*��o���m���(������ڥ���|��3��_�Eڣ��e��'�}��	bӾ`ĵ��"����������v��.ƾP���T�G�d܋��̿y�[*[�LƔ�c,��%������L=���w���m��W�l�J*�r���Ǜ޿���H.$���d�1 �������d��R���"V������]��}�c�I��:	ֿ_w����P�ɜ�m����ξRص��Ө�����H�������-ؾ�#�'�W�a��ß�_���-���u�6H��Q���X������Y.��~ڶ�v����U�v���� �5k��8�w�؞��W���X/���Y��E�����^����L���G���8Ӄ���?�~	����\ʾ�r���v���誾@���[2Ǿ��辸�[�9���}�����n	�\D����+���x����i���f�����Ϲ�����N]?��]�F��� ����N��w����� ����S��������)���e�~���4������:����k���.�$9��5�ZU¾�l�������V������$?Ѿ.|���u�'M�	z����ο����w\��m��QԺ�����Q��-���V������!n�r+�4 ���࿉���Y%�(�e�G�������j����  �  Z���a������$��eH����9#Ŀ����6L�/�7�����Ӿ�ù�La��ot������ߠ��½۾sK�Y$&���Y��q��a�ԿK��DW�ȶ���B���o���N���x���̟��(}�AU;�7���տ�@˿�Q��"���^����y�����1���`��i.���u�΄3�_���.[����y���:�3���ʾ׌������@��e����ZǾ�龉6��5��q�B���Y��:�,���m�h���=e����������"��\��k;f�=�'�,��S�̿n ҿق���4��u��b��AN��	��������P��R����$_�  ��~޿>��c��,��m	��5侚�ž���D��0(�����ڶ־����`����I�a���?P����GB�҂��W����������ۡ�����ހ��zAQ����^�心�˿��࿶���/J�#Ć�k���q��N��Uǽ�HȦ�LԆ���I������ƿi��ٶQ���"�V��o߾��ž�u���ϳ�}]���˾�辁��,��`��혿6Qؿ�?��Y�����#���R��N8��m���̠�5?�+|=�m8
��<ڿ�Ͽ�����V$�xa�E�������;$��M�������&@����w�à5��������������B����a��h�ھ@�ľ#ݹ�eA����¾}�׾W��[�B=�	>y��������!�.���o������t�������-��/6���3��fh��*��k���ѿWֿ��ſ6���w�5^��u=��<��������*��u����`��!�e��i����i�3a3�1����uҾ}_��.��R⻾#ɾ��ᾦx���!���N�9��>����(
��C�z��� ���P������LE��.������oR���M�3�Ϳ����bTK�BS������l����  �  (
���<��+��;:Z��m&������ó��	��j�U�� -�l�����w׾U>ƾ�i��ɾ]ݾ
�������5�2�`��d��G��2�̢1���e�`������̞��Y���ڀ�M�����x俘�����t<̿=@��^5��k�]���5���N��T��$�|���H����b�ܿWn��+�z�;�F���"�qb�<��s'Ѿ��þ?þ��ξ������4��B�U�s��:����Կ���/�B�a�v��V��^����	��@z���p�%;�$�
��VѿS�����L�ݿ`��G�DT|�M���9����+���_��7"l�-�7��>�f�ǿ����s�h��;����#�c��O�Ͼ�Ǿ��ʾ5�ھ�}���o�@�,���S��
��{ܯ�Q�!��OU�����+1��om���[������`���*�}@����Ŀ����H����V��xx%��<Z�L��� %��������C�����[���'�E��6{��sÊ��
[��2��{��K �<I�nSҾ�;˶վ��hY��d���;�0�g�lᓿF�ÿ���Ra3�ڷg�Eɋ�Fʛ�����J��^ց��O�������d���a���пnt��7�[6m��t��TL���c���g����~�b�J������࿽���ec��	)O�L�*���������_�,Ծ�nӾ],߾�9��i��Y'�}?J�v�{��Z��uٿd��<�D��y��f��H������I�����r�9=������տ�]���d�����L���I�sA~������m�����8��e�m�Ti9�8�	�˿���XQo�{�A�A@!�K�	�7U�ܾ�Ӿ*�־�u�wY�Z���%2�13Y�N����v�����uF#�ޠV������ڗ����� ��\���'Ma��,����\(ǿ����"ÿ>�����&��U[�]>��U����  �  ��k�[�b�-J���(�����տຬ��Y���r���N��m0�t �'������龑u�����_�Q�6�loV��{��8��@ڴ��Oῢ>��|0�o�P���f� rk��h]�J�?�'q���n���������Ѥ��p%ҿ�	��/���Q�`�g��k��,\���?�^D�8����ƿ��������wf�M�D���'��k��3���*��+�K������$��A�%8b���������¿�i�Y���;��jY�&j���h���T���3����]>ؿj"��7���g���N�����;M��<��[��k��Wh��(T���4��Q�/�翲繿�����k&\��3<��>!�������|��5���O�C���0�ŭN���q��v��%٪���ҿj����%�_�G�&�a�j�l�f�d�'�K�}(�t���-ȿ'������\����¿['��>$���H�;Lc��@m�8d�kK��*�Ab�H�ؿ�q�����x�|gT��6����_�	�˪��L<���� �p&���"���=��A]�<T�������Z��f�俔���82��jR�JCh�*=m��C_�}�A�Vr�K;�9���d䛿�T�����9�ֿ����1��S�Ѯi��=m��S^��A�d�%@��d˿(H��bǋ���n���L���/�2������\��i[���=�#8��,��*I��cj���m���V'ƿ����r���=�t�[�vGl��j���V���5�K��"�ܿ�j��8���zƙ�ֵ���4D���=�8�\�3�l��j���U��f6���a�L��7y���m����b�T�B���'�L����ŗ��p7 ���tv��-6�T�e4w�=���r���/տP��u'�=�H��	c�tn��Ff��)M�I[)�>���ʿ�r��
m�������ſ�/ �&%���I��Od��  �  �$��!��f����a�v�Ϳxo���4��r���nD��qh�yE�E�(������k���E.���L���p��������0⭿
o��q�ҿ���܇����5�"��/$�t�՞�%sݿ���n���9r�)�j��D���֞�?dȿDu��^�[!���$�����'�ZC����ݿ�ƿ{+��U���⓿�&��Q�\� ;���!�};�:{����7�`jX�*�}�đ����n8����Ŀ��ڿ�a��+�_N�`y$���!��Q�Ѐ��jOͿ����N|��C�k���o����䋫��Sؿ�D�.��(�#�<�#�o����	��(�l0ֿx?������$F�������Ew�^�R�c�3��+�K��ئ��.)�-�D���g��↿�f���D���r��4Ϳ�����H���� ���%�
�����P��1.���*�������m���|�cЕ�n���ˋ���||�D$&�cp"����_��.���Bп�%����5O��o��V$n�L�J�(�.�\����? ���4��S���w�$������_�������;ֿI`�1D	�4��D�$���%�������nb�2���@����z��rs�̖��W.��پ̿b������D#��'�����J�7A �q7�_˿�T���4��F���l>����d�U%C�*�)T������'���?�`�`�u���ٕ��8���W�� �ȿ4߿=����F��l���&��$�ku�%� ���ѿ�ꦿ]���c1t���w�S*��;���r.ܿ/!�w\�5�%���%�-��܆�v���:�ٿ�Ŀ�㳿����_ᑿo�}�_�X�r�9��K$�?��1��)�.�1<J�m�Y�������⬿���u�Ͽ�\�Z�����0M"�=2'�� �g��򿆠¿���i^���dr�����,��eʽ�ح���8~��  �  8忺�ѷ�͋���6��/�a�俽
ֿ2��M\��7��� ]�F�@�i�8��E���e�f1�����85ĿzGڿ �濦*鿠G�7v��?�~�翁!�H���ҿ����𣜿����rW�h>���9�Q�I� \m�����G���ȿ�/ݿ,��A�#���k�����[����i+�g8Ͽ����ۗ��)z��R�K9<�O
;���N���t������ѱ�؋̿X�߿�T������*�.(忺�迖��h�޿�˿$��%֒���q�3�L��S:���<���S�}��������6�п?q⿋��?��(^�[&俭��6����ݿWȿ"J��^��P
m�A�J���;���A�@	\�ꃿ!���Xڼ�M�տ�W���*B鿄��D�y6�j��>���ۿ��ĿlH�������g���H��=�0F���c����a}��^E¿��ٿ?�����3|��K�De�+��E��~P���ؿ� ���9��M#��sc���F���>���K� Wl�
s��KN��ҙǿ�ݿ#�^�쿹��k����E2뿇�����4sֿ낽�v������_���F��5B��~R�s�u�)D���[����̿��῀쿕V�i�m��5�Ӌ���M��Tӿ�0����$���Z��QD�z!C�>�V�R�|�|���7㵿=�пR��)t��쿹-鿊[�z^�����9�F�⿁NϿKF��\��/`z��U�t�B�W�D�]�[��s��}~�������Կ�����=��迡���&;�z뿈g࿔Q˿:���d���*Cs���P�6�A�o�G���a�z���Ă��)����>ؿ���k��*��+r�N�翋��Y���꿴�ݿI2ǿ�ͪ�w*��1�l��OM�{�A��
K��_h��A��ș��$SĿ��ۿ�  �  0���V��8�οȫ迺���F���!�f�$�fl��=
��^忇Ͷ��Ǒ��Uv�9|i�ɰ}�$阿Ģ��A�C��wG�S%�������x� �!t�<+ʿYз�A���˖��D����b��@�L%����<�����43��R���w�ʎ��t����������ֿ�8�s
�$C�"�#��S#�7j�-���}տ�J������q�n�+�l����������%п	- �m��{"�RX$���?@�"����iٿhÿ6���������l{��V��5�2�������3#�>=��(_�ל��c��Đ��X���&�ȿs/�w����j�����X%��� �M�������ƿ���B����l�Av�@�������̕�@��f��@@%��]#����fq�9��2,ӿT1���®��Z��4]��P�r��N�7�0��u��G��B���.��K���o�抿�*��Bɭ�3��W�ѿvj�>��#����"�8
&�������A�N���qƔ��h|�ϣo����r��f�ÿ�������� �ڿ&�IM!�9��A�����h�Ϳ�P��?��k������5j�m�G�Y-�����gN%���;�~-[�!��s���Ť������ſ�ۿ�v��v���Z�n&��d%�=x����y�ٿuZ��Ì���v�
�t�3��K��^4Կ�5��w���$��g&�I��bU�����ݿ��ǿs���M���Ք� 󁿈�^�q)>���&��=���B+�7�D���f�%?���똿�������̿��㿌����t �2
'���"��X�������ɿ���^M��`�r�� |�Ⓙ:}���b�7 
�A�Ə&���$�45��������տ!���dg��B������w�m�S���5��3"����[� ��.3�GP���s��,*���  �  ���]�����ؿB�� �*�չK��c�D�k���`�pE�̸ �H���8ѽ��Қ�����t����ȿ���2>)���L��d���k�\�_���D���"����Hο�O��<s���l���I��,,������� ��&�z��I�
�޷ ��<�Qy\�u���왿�b��RO�����E6�MNU���h�vqj�XmY�|�9�S'�"��/����픿�����]���ۿ��$�5�wV�Kci���i�/X���9�Ow�E<�E���Mޜ���� �_��	?�w%#��������Ұ���ə �^���)��7G�K�i�⃉���ʿ���*����A���]�3�k�$g�C�P�.��Q�
(пG	���Ӓ�>���'����$D�|B�[r_�{�l�r�f�#�O��n/�,M��.࿋������}��CX�$9�{
���
�����i��}���\�	�}E��7�F�U��z��p���b��pۿJ$
�K�+�M�R-e��:m�Kb���F�$."�r���G����ޝ��������̿MW���*�V^N���f��m�2{a�)�F�{�$�A��q�ѿ\Ъ�������s��%Q���3������	�+)��*���Ǟ�w�yA)�z�D�Se��̅��8������P��p���`8��eW���j�=�l�.{[���;��0���激�������ԏ��di����߿D����7�j�X��ok���k�')Z��<�ݎ�Kp��<�ÿ����䇿fh�+xG���+��!�8��h������Ae�ɝ��^1�RnN���p�b���G姿JkͿi� �s7!��sC�x_�om���h�;R�O�/���	�&8ӿ����ҕ�`؜����K���Ů���C���`�	�m���g��@Q�Ի0����m��u0���'��n)���o]�~8>�5$�-����]���d�����:�!��2;���Y��~��  �  ������������+)��(]�%J��H���I��.����̄�KV�d�!�6ￄ���`���u�ĿEE��i�,�Qb��Չ�����Sޞ�M���?��+�Q�Pp��A迫[��r���bN�+�'������{eԾ�6ž�t¾�0̾�>⾪b���͙;��(j�%6��7kʿPF
�m>:���n�LL��o���'��N���Apy�D�����ڿ�0��,���}Կ�5�E%>���s�Ӕ���x���N���[���/t���?�7�M9ѿ˱���p���?��R��d����;�þ�ľ'�Ҿ_o�[X
��Q%�&cJ�/�x�������qL�K��Kk��d������s���h��3�����ʿ笰�i���@鿑����P�ב��ܗ���Y��Լ���-����c�w�/�����Ӿ�c����a���6��
�s�������о)7ʾaо�F⾘j ��@��4���]�[����y������*���^�����٢��ں���t��A���\�W�X#��@�˿����o�ǿ<0��D.���c�ݨ��O_��o����Ж�����AS��- �k���ۮ�����NU��+/�ӡ��M��M+�Qվo�Ҿ��ܾ�g�
��#�,D�7�r������ο?g�v\<�O�p��W��U����/�����t{{�@'F��!�á޿�<��;7����ؿ�;�U,@��u�癑���_V���d��_Dv�(B����oտAꟿ�ux�I�G�ķ%���f���o)޾QӾO�Ծ�[����F��c~,��fQ����;��uz�/G���M�ץ���C��9���*����A���#j�b�4��P�Ϳ#��������6�Zn��5R��D���E�����oc���ӊ�@e�[ 1���Hy��e���j�f�y�;�:!����/���cھ{Ӿ�پ�����i�*(8���a��  �  �-���ȿum�' L��	����������~���t}���¤��D���E�F�Xܿk�ɿ��濇���S�����)�����g���0��kA��+{��Q�=�A��㸿.���W=C��u��X��SFϾB�������k��Qf��u,þ���:L	�'�-��Re�#J���^�a�"���b��E�����l���}���	�����S�q��1�~��A�пWο�#��*+��#j�e ��U���f���4s��w&���ז��	j�CY)�����>��k�l�!;2��D��o��žӱ�<����o��2;���H;���F����>��\��v���O �@M7��y���]9���/��p���TI����#�[�$���0�Z�˿e ٿ��
�Y?��Ҁ�G١����]���z���4��G���lT�UR�YHҿNs��kZ�'�������o�žަ��iE��I��~eľ �߾u��`|$��T��B�ʿ��]�M����Z��9���BQ���2��Z}�� ��OG����P߿>�̿������]U�����D�������A��z�����]Y����?�)��Sc�����mJ����G*��޾��ƾ����Ķ��������Ӿ"~���i 6���m��������%�8�d�#S��s���Wv������i�����u�s�h�3�����Կe*ҿ�.��/0-��*l����S���x����z��./��	��� l�Kr+���￺u��Q*u��:�h��8��3־0¾�������o�ž�Gܾ�Q �P��ԞE�J���۵�:��K�8�1k{����:��L���p��T��ϲ��(I]�N!��-���ο��ۿ�p�d�@�%�������$���ۍ��
����۫�z��^�U�����Կ-���N_���,������_Ͼ�)������$���(;�����(���X��  �  G���� ؿJ� ���f��ޚ��1��[���dJ�����������[���_�� �j�� �ܿ���^,��p����H���x������tW��f׷��"��%V��[���ſ�n��0A����J��������n'���"���d������P�Ѿ����(���g�"������{6�����&˧��P����������UE������E��-KH��<��'���J����@�����ȫ�-_������B����N����{ڄ�'>��A���Awp�6.�L��ޮվ(_���������c��f榾+ϼ�c� ����;��Ղ�yC��7n�`^N�4���.��P��'���e����^������G-y���3�����߿h���'��CX�TX��n��Z���{������)�����Gbp���(��㿎њ���Z��"�Q����оL����ަ�Q���i��w�����ξr�����jXT�8i��z�ڿc�!��;h�u���1���]��o����g��z?�����a���!�����7�߿S	�e�-�q��ٟ������������3��#�������S�W�B��zɿ�����]H�K�4����;Z�����B^���᱾\�þg�⾩%
�5�1��np��檿k^��̛8�i���Hب�\��O�������L��3���J���RJ�TC�53���ޓ���B�"��
ͬ�d����������W�������� @�>%� ᱿[�x���6��0��@���ž��������0����˾���]����B�0E��������P�-Î�r��P���Š��wb��'���m���z�5�cR�b����ݨ���Y�����ո�����W,����������LV���q�X�)��_�mu���_�&6'���!�ھ�q���a���H��2k��]���M׾�� �Ǘ"�UX��  �  L��^T޿a�&���p�ϡ������q��{e��C8��&������6i��^&�������h���D3��_z���:I���g��/,��������̧��Z@_�����D˿'L��"CA�b��ྍ���V颾鑗�����W���g��\�̾Z��8(�4�i��%��B4����=�)(���U���b��G�������Go�������;����P������7F������H�è���P���e����������*�������!�����E��j�ꗱ�0�r��-����z�о{h��/	���4��|���P ��fз�\�ܾ���j�;��n��ÿ�}�B
W�M<���I��'���e����f�����gҪ����`�:�/���
���!�^a������/��':�����(�������lҦ���z�q)/���!�����[��� �Z�����˾1ǰ�8��,����ɡ�7���S�ɾ�������U�Hߗ��ῳ,(�58r�:��,���!���������~��3���Z�j���'��������}���4��{��ͦ�m���9�������������\�����`����(�ο�Ԍ�pH� l�T���Ⱦ����C}��pѥ�{(��[�����ݾ�]�0�L:r��k��#����?��6���b��&n����������u������@��1�R����z��.Q�����J�6����T���j������������������fŋ���G���M͵�U{��5�A-��P�����c2��������e����ƾ�%�����B��݇�tuƿB,�r�X�������Q]������3��/�����������S<�R�	�E�q����"�C�b�r��T���K���XB��Q�������{��/!|��|0�D�@��_�`�!�%�R��r�վ����+����æ��ʪ�H{���GҾ)���-!�qY��  �  G���� ؿJ� ���f��ޚ��1��[���dJ�����������[���_�� �j�� �ܿ���^,��p����H���x������tW��f׷��"��%V��[���ſ�n��0A����J��������n'���"���d������P�Ѿ����(���g�"������{6�����&˧��P����������UE������E��-KH��<��'���J����@�����ȫ�-_������B����N����{ڄ�'>��A���Awp�6.�L��ޮվ(_���������c��f榾*ϼ�c� ����;��Ղ�xC��7n�`^N�4���.��P��'���e����^������G-y���3�����߿h���'��CX�TX��n��Z���|������)�����Gbp���(��㿏њ���Z� 	"�Q����оM����ަ�Q���i��w�����ξr�����iXT�7i��y�ڿc�!��;h�u���1���]��o����g��y?�����a���!�����7�߿S	�e�-�q��ٟ������������3��#�������T�W�B��zɿ�����]H�K�5����;Z�����C^���᱾\�þg�⾪%
�5�1��np��檿k^��̛8�i���Hب�\��O�������L��3���J���RJ�TC�53���ޓ���B�"��
ͬ�d����������W�������� @�>%� ᱿[�x���6��0��@���ž��������0����˾���]����B�0E��������P�-Î�r��P���Š��wb��'���m���z�5�cR�b����ݨ���Y�����ո�����W,����������LV���q�X�)��_�mu���_�&6'���!�ھ�q���a���H��2k��]���M׾�� �Ǘ"�UX��  �  �-���ȿum�' L��	����������~���t}���¤��D���E�F�Xܿk�ɿ��濇���S�����)�����g���0��kA��+{��Q�=�A��㸿.���W=C��u��X��SFϾB�������k��Qf��u,þ���:L	�'�-��Re�#J���^�a�"���b��E�����l���}���	�����S�q��1�~��A�пWο�#��*+��#j�e ��U���f���4s��w&���ז��	j�CY)�����>��k�l�!;2��D��o��žӱ�;����o��1;���H;���E���>��\��v���O �@M7��y���]9���/��p���TI����#�[�$���0�Z�˿e ٿ��
�Y?��Ҁ�G١����]���z���4��G���lT�UR�YHҿOs��lZ�Ó'�������p�žަ��iE��H��~eľ��߾u��_|$��T��B�ʿ��]�M����Z��9���BQ���2��Z}�� ��OG����P߿>�̿������]U�����D�������A��z�����]Y����?�)��Tc�����mJ����H*��޾��ƾ����Ķ��������Ӿ#~���i 6���m��������%�8�d�#S��s���Wv������i�����u�s�h�3�����Կe*ҿ�.��/0-��*l����S���x����z��./��	��� l�Kr+���￺u��Q*u��:�h��8��3־0¾�������o�ž�Gܾ�Q �P��ԞE�J���۵�:��K�8�1k{����:��L���p��T��ϲ��(I]�N!��-���ο��ۿ�p�d�@�%�������$���ۍ��
����۫�z��^�U�����Կ-���N_���,������_Ͼ�)������$���(;�����(���X��  �  ������������+)��(]�%J��H���I��.����̄�KV�d�!�6ￄ���`���u�ĿEE��i�,�Qb��Չ�����Sޞ�M���?��+�Q�Pp��A迫[��r���bN�+�'������{eԾ�6ž�t¾�0̾�>⾪b���͙;��(j�%6��7kʿPF
�m>:���n�LL��o���'��N���Apy�D�����ڿ�0��,���}Կ�5�E%>���s�Ӕ���x���N���[���/t���?�7�M9ѿ˱���p���?��R��d����;�þ�ľ&�Ҿ]o�ZX
��Q%�%cJ� /�w�������pL�J��Kk��c������s���h��3�����ʿ笰�i���@鿑����P�ב��ݗ���Y��Լ���-����c�x�/�����Ӿ�d����a���6��
�t�������о)7ʾaо�F⾗j ��@��4���]�Z����y������*���^�����٢��ٺ���t��A���[�W�X#��@�˿����o�ǿ<0��D.���c�ݨ��O_��o����Ж�����AS��- �l���ۮ�����NU��+/�ԡ��M��N+�Qվp�Ҿ��ܾ�h�
��#�,D�7�r������ο?g�v\<�O�p��W��U����/�����t{{�@'F��!�á޿�<��;7����ؿ�;�U,@��u�癑���_V���d��_Dv�(B����oտAꟿ�ux�I�G�ķ%���f���o)޾QӾO�Ծ�[����F��c~,��fQ����;��uz�/G���M�ץ���C��9���*����A���#j�b�4��P�Ϳ#��������6�Zn��5R��D���E�����oc���ӊ�@e�[ 1���Hy��e���j�f�y�;�:!����/���cھ{Ӿ�پ�����i�*(8���a��  �  ���]�����ؿB�� �*�չK��c�D�k���`�pE�̸ �H���8ѽ��Қ�����t����ȿ���2>)���L��d���k�\�_���D���"����Hο�O��<s���l���I��,,������� ��&�z��I�
�޷ ��<�Qy\�u���왿�b��RO�����E6�MNU���h�vqj�XmY�|�9�S'�"��/����픿�����]���ۿ��$�5�wV�Kci���i�/X���9�Ow�E<�E���Mޜ���� �_��	?�w%#��������Ѱ���ə �]���)��7G�I�i�჉���ʿ���*����A���]�2�k�$g�B�P�.��Q�
(пG	���Ӓ�>���'����%D�|B�\r_�{�l�s�f�#�O��n/�,M��.࿍�������}��CX�$9�|
���
�����i��|���[�	�|E��7�D�U��z��p���b��pۿI$
�J�+�M�R-e��:m�Kb���F�$."�r���F����ޝ��������̿MW���*�W^N���f��m�3{a�*�F�{�$�A��r�ѿ^Ъ�������s��%Q���3������	�-)��+���Ȟ�w�zA)�z�D�Se��̅��8������P��o���`8��eW���j�=�l�.{[���;��0���激�������ԏ��di����߿D����7�j�X��ok���k�')Z��<�ݎ�Kp��<�ÿ����䇿fh�+xG���+��!�8��h������Ae�ɝ��^1�RnN���p�b���G姿JkͿi� �s7!��sC�x_�om���h�;R�O�/���	�&8ӿ����ҕ�`؜����K���Ů���C���`�	�m���g��@Q�Ի0����m��u0���'��n)���o]�~8>�5$�-����]���d�����:�!��2;���Y��~��  �  0���V��8�οȫ迺���F���!�f�$�fl��=
��^忇Ͷ��Ǒ��Uv�9|i�ɰ}�$阿Ģ��A�C��wG�S%�������x� �!t�<+ʿYз�A���˖��D����b��@�L%����<�����43��R���w�ʎ��t����������ֿ�8�s
�$C�"�#��S#�7j�-���}տ�J������q�n�+�l����������%п	- �m��{"�RX$���?@�"����iٿhÿ6���������l{��V��5�1�������3#�==��(_�֜��c��Ð��V���$�ȿq/�v����j�����X%��� �M�������ƿ���B����l�Bv�@�������̕�@��f��A@%��]#����gq�:��4,ӿU1���®��Z��5]��Q�r��N�8�0��u��G��B���.��K���o�抿�*��Aɭ�2��U�ѿuj�=��"����"�8
&�������A�N���qƔ��h|�ϣo����r��f�ÿ�������� �ۿ&�JM!�9��A�����j�Ϳ�P��?��k����� 6j�n�G�Y-�����gN%���;�~-[�!��s���Ť������ſ�ۿ�v��v���Z�n&��d%�=x����y�ٿuZ��Ì���v�
�t�3��K��^4Կ�5��w���$��g&�I��bU�����ݿ��ǿs���M���Ք� 󁿈�^�q)>���&��=���B+�7�D���f�%?���똿�������̿��㿌����t �2
'���"��X�������ɿ���^M��`�r�� |�Ⓙ:}���b�7 
�A�Ə&���$�45��������տ!���dg��B������w�m�S���5��3"����[� ��.3�GP���s��,*���  �  8忺�ѷ�͋���6��/�a�俽
ֿ2��M\��7��� ]�F�@�i�8��E���e�f1�����85ĿzGڿ �濦*鿠G�7v��?�~�翁!�H���ҿ����𣜿����rW�h>���9�Q�I� \m�����G���ȿ�/ݿ,��A�#���k�����[����i+�g8Ͽ����ۗ��)z��R�K9<�O
;���N���t������ѱ�؋̿X�߿�T������*�.(忺�迖��h�޿�˿$��%֒���q�2�L��S:���<���S�}��������5�п>q⿊��=��&^�Y&俬��5����ݿVȿ!J��
^��O
m�A�J���;���A�A	\�ꃿ"���Yڼ�N�տ�W���+B鿅��D�z6�k��?���ۿ��ĿmH�������g���H��=�0F���c����`}��]E¿��ٿ>�����1|��K�Be�*��D��}P���ؿ� ���9��M#��sc���F���>���K�!Wl�
s��LN��әǿ�ݿ$�_�쿻��l����F2뿈�����5sֿ삽�v��� ���_���F��5B��~R�t�u�)D���[����̿��῀쿕V�i�m��5�Ӌ���M��Tӿ�0����$���Z��QD�z!C�>�V�R�|�|���7㵿=�пR��)t��쿹-鿊[�z^�����9�F�⿁NϿKF��\��/`z��U�t�B�W�D�]�[��s��}~�������Կ�����=��迡���&;�z뿈g࿔Q˿:���d���*Cs���P�6�A�o�G���a�z���Ă��)����>ؿ���k��*��+r�N�翋��Y���꿴�ݿI2ǿ�ͪ�w*��1�l��OM�{�A��
K��_h��A��ș��$SĿ��ۿ�  �  �$��!��f����a�v�Ϳxo���4��r���nD��qh�yE�E�(������k���E.���L���p��������0⭿
o��q�ҿ���܇����5�"��/$�t�՞�%sݿ���n���9r�)�j��D���֞�?dȿDu��^�[!���$�����'�ZC����ݿ�ƿ{+��U���⓿�&��Q�\� ;���!�};�:{����7�`jX�*�}�đ����n8����Ŀ��ڿ�a��+�_N�`y$���!��Q�Ѐ��jOͿ����N|��B�k���o����㋫��Sؿ�D�-��'�#�;�#�o����	��(�k0ֿw?������#F�������Ew�]�R�b�3��+�K��ئ��.)�.�D���g��↿�f���D���r��5Ϳ�����I���� ���%�
�����Q��1.���*�������m���|�cЕ�n���ʋ���{|�C$&�cp"����^��-���Bп�%����4O��o��U$n�K�J�'�.�[����? ���4��S���w�%������_�������;ֿK`�1D	�4��E�$���%�������nb�3���@����z��rs�͖��W.��پ̿b������D#��'�����J�7A �q7�_˿�T���4��F���l>����d�U%C�*�)T������'���?�`�`�u���ٕ��8���W�� �ȿ4߿=����F��l���&��$�ku�%� ���ѿ�ꦿ]���c1t���w�S*��;���r.ܿ/!�w\�5�%���%�-��܆�v���:�ٿ�Ŀ�㳿����_ᑿo�}�_�X�r�9��K$�?��1��)�.�1<J�m�Y�������⬿���u�Ͽ�\�Z�����0M"�=2'�� �g��򿆠¿���i^���dr�����,��eʽ�ح���8~��  �  ��k�[�b�-J���(�����տຬ��Y���r���N��m0�t �'������龑u�����_�Q�6�loV��{��8��@ڴ��Oῢ>��|0�o�P���f� rk��h]�J�?�'q���n���������Ѥ��p%ҿ�	��/���Q�`�g��k��,\���?�^D�8����ƿ��������wf�M�D���'��k��3���*��+�K������$��A�%8b���������¿�i�Y���;��jY�&j���h���T���3����]>ؿj"��6���g���N�����;M��<��[��k��Wh��(T���4��Q�.�翱繿�����j&\��3<��>!�������|��6���O�D���0�ƭN���q��v��&٪���ҿj����%�`�G�'�a�j�l�f�d�'�K�}(�u���-ȿ'������\����¿['��=$���H�;Lc��@m�8d�kK��*�@b�G�ؿ�q�����x�{gT��6����^�	�˪��L<���� �q&���"���=��A]�=T�������Z��h�俔���82��jR�JCh�*=m��C_�}�A�Vr�L;�9���d䛿�T�����9�ֿ����1��S�Ѯi��=m��S^��A�d�%@��d˿(H��bǋ���n���L���/�2������\��i[���=�#8��,��*I��cj���m���V'ƿ����r���=�t�[�vGl��j���V���5�K��"�ܿ�j��8���zƙ�ֵ���4D���=�8�\�3�l��j���U��f6���a�L��7y���m����b�T�B���'�L����ŗ��p7 ���tv��-6�T�e4w�=���r���/տP��u'�=�H��	c�tn��Ff��)M�I[)�>���ʿ�r��
m�������ſ�/ �&%���I��Od��  �  (
���<��+��;:Z��m&������ó��	��j�U�� -�l�����w׾U>ƾ�i��ɾ]ݾ
�������5�2�`��d��G��2�̢1���e�`������̞��Y���ڀ�M�����x俘�����t<̿=@��^5��k�]���5���N��T��$�|���H����b�ܿWn��+�z�;�F���"�qb�<��s'Ѿ��þ?þ��ξ������4��B�U�s��:����Կ���/�B�a�v��V��^����	��@z���p�%;�$�
��VѿR�����L�ݿ`��G�CT|�M���8����+���_��7"l�,�7��>�e�ǿ����r�h��;����#�b��N�Ͼ�Ǿ��ʾ6�ھ�}���o�A�,���S��
��|ܯ�R�!��OU�����+1��om���[������`���*�}@����Ŀ����H����V��xx%��<Z�K���%��������C�����[���'�E��5{��rÊ��
[��2��{��K �;I�mSҾ�;˶վ��iY��d���;�1�g�mᓿG�ÿ���Sa3�ڷg�Eɋ�Fʛ�����J��^ց��O�������d���a���пnt��7�[6m��t��TL���c���g����~�b�J������࿽���ec��	)O�L�*���������_�,Ծ�nӾ],߾�9��i��Y'�}?J�v�{��Z��uٿd��<�D��y��f��H������I�����r�9=������տ�]���d�����L���I�sA~������m�����8��e�m�Ti9�8�	�˿���XQo�{�A�A@!�K�	�7U�ܾ�Ӿ*�־�u�wY�Z���%2�13Y�N����v�����uF#�ޠV������ڗ����� ��\���'Ma��,����\(ǿ����"ÿ>�����&��U[�]>��U����  �  Z���a������$��eH����9#Ŀ����6L�/�7�����Ӿ�ù�La��ot������ߠ��½۾sK�Y$&���Y��q��a�ԿK��DW�ȶ���B���o���N���x���̟��(}�AU;�7���տ�@˿�Q��"���^����y�����1���`��i.���u�΄3�_���.[����y���:�3���ʾ׌������@��e����ZǾ�龉6��5��q�B���Y��:�,���m�h���=e����������"��\��k;f�<�'�+��S�̿n ҿق���4��u��b��AN��	��������P��R����$_�  ��~޿=��
c��,��m	��5侚�ž���D��0(�����۶־����`����I�b���@P����GB�҂��W����������ۡ�����ހ��zAQ����^�心�˿��࿶���/J�#Ć�k���q��N��Uǽ�HȦ�LԆ���I������ƿi��ضQ���"�V��o߾��ž�u���ϳ�}]���˾�辁��,��`��혿6Qؿ�?��Y�����#���R��N8��m���̠�5?�+|=�m8
��<ڿ�Ͽ�����V$�xa�E�������;$��M�������&@����w�à5��������������B����a��h�ھ@�ľ#ݹ�eA����¾}�׾W��[�B=�	>y��������!�.���o������t�������-��/6���3��fh��*��k���ѿWֿ��ſ6���w�5^��u=��<��������*��u����`��!�e��i����i�3a3�1����uҾ}_��.��R⻾#ɾ��ᾦx���!���N�9��>����(
��C�z��� ���P������LE��.������oR���M�3�Ϳ����bTK�BS������l����  �  �L��G���?c�������b��2�Rӿ[���Y[K�
��l�3%þ4	�������3��^䞾����I�ʾ6����� �^�Z��G��.翧Q+��s�g��o���s��t����6��ֵ��ӏ���S�����K�޿ 0�Xb6���|�l���f������{D��ב��d��������I��
���`���7���
��_ݾ���:���C������녣������Sؾ��$Y1�k\u�·�����w�A�[����޻��Y���T������@���?���U/=��-	�B`�i�濼��4�K�\m��*��n���m���(������ڥ���|��3��_�Eڣ��e��'�}��bӾ`ĵ��"����������v��/ƾQ���T�G�d܋��̿y�[*[�MƔ�c,��&������L=���w���m��W�l�J*�r���Ǜ޿���H.$���d�0 �������d��R���"V������]��}�c�H��9	ֿ_w����P�ɜ�l����ξRص��Ө�����H�������.ؾ�$�'�X�a��ß�`���-���u�6H��Q���X������Y.��~ڶ�v����U�v���� �5k��8�w�؞��W���X/���Y��E�����^����L���G���8Ӄ���?�~	����\ʾ�r���v���誾@���[2Ǿ��辸�[�9���}�����n	�\D����+���x����i���f�����Ϲ�����N]?��]�F��� ����N��w����� ����S��������)���e�~���4������:����k���.�$9��5�ZU¾�l�������V������$?Ѿ.|���u�'M�	z����ο����w\��m��QԺ�����Q��-���V������!n�r+�4 ���࿉���Y%�(�e�G�������j����  �  ������`����]����Q����Ŀ+兿_	=� ����پ#j��3E��k$��P쌾���T��H���V����h�K�q����ֿd��	�a��y�����l���g������[��5���5D�Do�|�ܿ�1ѿt����Q)��j�e5�����������bW��N��)���:�+ �󶬿��m�k�*��X ���˾O���_ގ�M_��4b���<��*Ǿ7���$��yd��L�����?�3�Xz�"��ɴ��������*ٻ�z���q�͉/� �
�ҿ�oؿ
��A=�[��l����V��I�������L��#���M&j�=�%��=����rRU�$������¾�r���>���u�������������2^۾����9�g�����]��T�J��ĉ�_���]��.��:���1�����S~[�5X�[��:[ѿ�� ����S�����>�������w��5����1������S����=ǿ����<�B��[��8��������w6���E�������h����Ǿ��� ���R����9ڿ�y �Imc�|Y��Q��iO���Q������\���'���^F�&��v��U�տ7W���+�pHl��M���������D���j��T��C8���=�d+��ް�v�k�2�Å��+ܾl\��&�������������m��c׾���~�,���l�k���&��7�5�k|��/���ÿ���h�����E���t���1��@�׿�ܿE�
�D0?�6��|���ZG��1��������&���z���k��'�d�俟���\��k"�߾��f�Ͼ�������u���Ϡ��������N�Lw�@A?�����������8L�l��d5����L�������Zϳ�AU����\����Z�®ӿ�Y����yU�CR���~�����  �  �����J��A���R���.I�����O���냿8�<��0�2޾����ʠ�8q��=$��Aq��i��\J����R �r�J����T�п9��WX�����5��G����|���X���=�����a<�K^��տG�ʿ\���"��r`�����:*������������ԝ�1dw�P�3�"��� Ȩ��[k��*���dо�ï�xc�����o����̚��ݬ��˾k���*%�eb�!���k-��,�jyo��0���z��u���5�����Li����g���(�Kh���q̿E�ѿ���S�5�'[w�lƝ��"������5���P��T
���i`�ū��ڿ�ҕ���S�%��8���tǾ{
������Ǯ��{`��� ��`@����߾���Y�9�Я��	:��E����B�4��S ���ս�!:��]�����������R��t��
濣;˿5��U.�	kK�ׇ�$��������������*���"���J�����¿S���(B����a�龴�þo���D����}�����k���lw̾��c��7�Q� ���Q	Կ9���Z���������f��M��b>��l�����>��
��ڿ4gϿf����%��b�Nړ�9A���4�����l�������y�'�5������﬿)�s�3�-D
����� ��V����L��,Ȣ����������۾L���S-�m�j�iݥ�WQ񿇬.��q��>��쉷��.��7G��n��}��j�K�*����j�пu'ֿ,���7�:hy�8�(��������*��{���b�@\!���ݿM0��<�Z�"`#�"\ ��CԾ�����㨾 �������q��Dnƾܱ���$?��M���ӻ����D�Ñ���ȥ��}������ZD��J>���;��X�S�����]� �Ϳe�|W�ڐL��f���������  �  D��в��RC��'�m��f2�l���F���C�w�=�<���B��Ǿ�b������f��}:��=糾k�ξv9��M��J��2��N���@o	��V?��S{������������p��ˣ���`�X'�q��*�¿�й��ٿ$��F����E�������s���1���y���Y� �M��!4��]�f�J�-�Ϋ���߾���������������,騾	���=۾�>�9�(�7�^��1���	ٿ� �p!S�VN��@���q����������.��"xL��&�s�߿�����O�z4!�d�Y�����@���_���U��	}��/#���LF�OC�bpɿ�#���{R�	S!����׾����q��������妾�w����ʾi��-����;�^0z��h��
&��_-�r1h��ߐ��y��Z�������Ö���u�|>:�Kg�0ѿ�Y��q�̿>��$4��(o����P��� ��c������Po���3��c �����D\��(-C�I������Ӿ�0����������ڰ�h����ܾ���f�!��Q�v���.]Ŀ�-��A��}�����������gb��&���Ӫb��#)�on��wHǿ�8��#޿�R�EH����4���s*��I����D��ኋ��\��5"��$濾[����n�96����&"�DϾiѺ�����j ������9̾Sv뾹`���0��g��O��w-ݿ�5��9U��[��G���Ǯ�z��?���B����N��P�����^��-�ÿ+��J#���[�-���"u��я�����0U��������G�O����̿����,Y�h�'�[������Ǿ+Ƕ���������龾��վ9���&���@��k��������d.���i�刑��"���M��<���Ec��
�v��n;�u�	��lӿᬼ�^�οL�<5��Dp�E�������  �  ��������R�m�(	B����z�ܿ*P��v{��bF��s!�T���~�ʾ6�|��l���Xо���]�S�(�r�P���Q��Kq����XL�vtv��Z��Č��]����d��[6�G�	�3�ο����{���F������!���P���z�u��Z������!0`���2�8'�Hȿ���g��)9��.���Ûܾ,žu긾T=��gþ�Dپ ������4���a�T��-^��n���-��=[�������"0��S~�u�U��&�F���g���z��^ ��\ɿQ0�y,1�!�_�_��$����}����z���Q���#��V�� 𵿱Љ���W�?�.����e��Շ׾ľ�������ڕξd��ʃ��!�+=E�n�w�O���׿D�"�=�{Sj����=b��mۈ��*s�rG�÷�)���ܳ��r��hk��v�ݿ���B��n��̇�ѩ��y����;o��iC�4���߿���H����K�='�YW�I�񾑫־�ǾG�¾�2ʾ��ܾ���4���/��W����β�����V �vN��0x�8;��N����L��xxf��b8�Q���;ӿ<ڬ��쥿}c��������#�#�R�\�|�����_n��y���FRb�h�4�B	��>̿i��tp��`A��> ���L�쾋Lվɾ�hȾ�BӾNu�+�����*�<���i�Qr��	�ſ]���/��X]�v��Pь�wA���;��E�W���(�
���u�¿!æ�@��75ͿE=�g)3�-�a�I˃��o�� X����|�*{S��%�T����P��'/��ڋ^��5��f�����來cоcȾ!T˾�ھ�����;�&���J��(}�d���ڿ�b�+?�r�k�YȆ��
������mt��RH�C����L4���Ť�4�����!��C�p��O���  �  �hQ�/�I��3��������¿]����M��̳`��@��[$�>��z���⾌�۾��徬O��n��I*�DG�si�P���	����̿ �����9�"�L��Q���D�U�*�,&
���տ�|������&���eݗ�T���{n�����v:��M�Y�P���C��*�V��3�8����&��пz���U�6�6�*��R'������޾�޾1�쾞
����e�3���Q���u����ZV��3oܿ3�	��'�m[A�#�O���N��=� ��B���ÿ�嚿�P��҉��`����Ͽ���n'���B���P��mN��<�Jw!���K�ҿ�Q��*��yo��tL��O/����P���쾏���M澅k��?-��$��G@��c`�����M��q��"i￿��K�1�ǴH�cSR��fK�c5�}*�g��+���&���ꇿ(Ƒ���������2�L�I��R���J��R5�gP��>����ſ�D��x���4f���E��	*�m	���$"B��6�%��ݜ�
�0���M�;�o�����>���/п���.v�zz;��N���R��{F���,��#�ڿ䯪�܏�` ���4��=�¿m������M�<���O���R���E�-��-�ji濷ٹ��N�����O�]��?���$�\E�����-�h@�����"���!��;���Y��+~����z�������)��xC�R���P��=?�&5"��E��!ȿ�(��[�������%�ӿz���O)��`D�=�R�� P��>� $#�7M��ֿ���Z���H�u��S�L�5�/�ג	�W���i��/�l��u��O`*��E�+�e�]M�����h�¿������83��J��S�7�L�u�6�Lh�D�����퀖��=�����(Ƴ��G�����3���J��  �  N�9��c���}$ҿ�ػ��ʪ�y������y�>�V��6�lM�UF�������qS"���=��|^�Ld������q���g���o���ؿ"����_��������	�6��ȿ�f�� с�	U`�C�Y�-�p�i��Cµ���߿�#����|�xr�<� �!��xPʿ����2��"w���쇿�n�� L���-��.�N�
��
��5�B�*��cH��j����O����I���೿j�ǿB(�9`���,�H��������	�M��Ӿ���ot�r�Z��^�Xa~�Z���:�ÿW��7��Λ����<!
�k�����ۿٔÿ}�� 顿�2���7��`\d��OC��Y'�,��w����D�6��ZV���x����ES��=���'���Eѿ��쿷��L��i�T�� ��ؿ�Ү�������l�m�\�)�i�A���-ު��ӿ����,�������_��4��u�Կ[�������Ҟ��ŏ�H�~�2z\��<�L:#�3Q�����7�N�(�<0D�
)e��Ƀ�y
���좿h汿��ÿx�ۿU)���
����������J���G̿an����N�h�	Wb�� y�}������] 俥N�~6�7��K���	������οS(���7�������Gv� ET���5��G�����.��K���2��P��?r���ə��g����Ż˿�W忑J��I�|>����m��fM迏J��X�����|���b�;Df�	=��������ǿ�p�b
��W�Ou�A���&���E߿��ƿ�h��I��Ë��u�����j��I� �-���9�����#��m<�Y�[��~�������k���G<����ӿt5��(������4��e�'�ڿAF��R����q�fya�݄n�[���>��W�տ|������  �  �dϿL[ӿ�ѿ(EϿ=^Ͽ��ѿ�^ӿ��ο����⬿(r���u���L�73�85,��7�ѣT����UL���2���ſ�п��ӿ|sѿ�=Ͽ��Ͽ&�ҿ�UӿѡͿ��������K����m�u�G��O1��#-�g�;��E[����ĝ�����Yȿ'�ѿS�ӿOѿ<Ͽ�[п�ӿFӿ��˿��
䤿���{�f���B��\/��L.���?��a��2����������vʿ7�ҿLӿ3tп��οd�п�ӿk+ҿ��ɿ <��?c�������R_�>��-���/�G�D��Vi�������������!Ϳ/�ӿ�ӿ��п��Ͽ3�ѿ�HԿnRҿ�Qȿ����5:�������7[�?�<�R@/�]�4�YL�[s��4��t竿9���-�Ͽ�"տ $Կr|ѿbѿAWӿ�Kտ�.ҿ��ƿɲ�ʙ�����Z�V���:���0� 9��TS� |�xb���ǰ�B�ſ/%ҿ�ֿԿҿ�ҿ\�Կ)ֿ4�ѿn�Ŀ#���[N���z�f�R���9��\2���=��[����'���r����.ɿFԿ�	׿��Կ�ҿ�Vӿ
ֿ��ֿO/ѿſ¿*���A'����u���O���9���5�5(D�4�c�T`������g���̿63ֿ��׿�Zտxӿ��Կ�;׿j/׿1п��������%����n���J��r7��a6��G�mj�0@��������s�οɠֿk?׿�ԿH-ӿX�ԿuX׿�gֿ��Ϳ�{��ݡ���ي�۽g��mF�X�5��8��L��q������Q�����пN;׿�ֿ�HԿ`Uӿ�TտB�׿��տҩ˿���� v��6؆��oa��B��?5��}:���Q���x�%��������kĿ0wҿv�׿�ֿ�ԿȨӿ9�տ]�׿��Կ�Iɿ�[��$P������[�$�?��.5���=���W�Oj���~���ղ���ǿ�  �  �֜�]����漿\�ӿ�ￋ$���s9�������d Ͽ�^���ꅿ��c�I�X��qj�80�������~ؿe- �yp�\��x��4��:鿺-ο ḿ�q��֙�y�����s���Q� d2��:�� �[	�����&��#C��d�@T���H��a����;���Ŀ~�ܿ����hp
��������)�h0��͓��_�{�+C]�t�[��w�ǖ�������.��&E�4���6�����߿�Iƿ�ڲ�0^��O���R���q�g��KF��#)���8�	�i3��b���/�"�N�5�p��U������ň�������P̿;�濉��V�(�� ����2@޿텴�����:�p�)�[�
d�6���ˣ�h�˿B{��<k�/���U�o������\ؿ	��sD�� h�������P��kq`���?��.%������zr��6#�L^=�!�]��������b���^��3����KֿVN�(�~�W���N�����o�ѿfN��:爿��i�}�^���p�[���1���ۿ��\'�7I�T��"�����ѿ\[��f��a���(���{��%Y�!8:�#?"�0/���o�%/��K��m�򡇿����2I������#Tȿ��࿅���4��n��8���	�;?�BſS���{ ���Xe��c��'��Қ�X��������1Q���`��A{ ���㿒|ʿ��[�������+���Up���N�r}1��^�L��n9�<> �wr7��V��x��܌��S��������Ͽ81�!������֞�^A�bvῸ����ד�1�v���a�w�i��i��०���ο�5������#�����	�d����ڿ��ÿ걿����(��:僿6�e���D�	*��@�G����ɡ'�R�A�C�a���������  �  H���B9���&ſ����4��Kj5�nJ��dQ�A�G���/�b���g߿�㬿e���υ��Q��7���L��*��5�ANK��TQ���F�w�/������,��4Ù��̀��4[�s�;�� �k<
�����ݾ�Z�C/�i��/��L�b�o�	ԍ�����[�Կ�����"���=��N�<"P��$A���%�?��n�̿�����C�����ۜ���ƿN
���!��>�H1O���O��4@�v�%�F�#�ٿD>���q���s��O���1�~A�G��Jc�X�ݾR�߾lq�ԩ�����K9�3�X�A~��W��?}��_��1���,��7E�~cQ��BM�Su9�	=���������z��x���l���橿oxڿ����$-�X�F�xR���L��99�������S�˿�����
��~�j�;I���,�)��j�:�N����EG��G���*���F�q�g��@��F�����ǿxJ�������6���K�`�R��I�!	1�,��]�寿�n��Wሿk��������r���7�{M�S��H�-A1�^���6����C��uX���jb�<�B��(����׵����6����7�
�d����7�+U��2x�����̯���ؿ-����$�r�?�/�P�02R��1C�/�'�����п�����N�����j堿%�ʿ����#���@�=Q�ܤQ��EB�I(��
���ݿ�s��ѩ��K�{��*X��!:�d� �t$��������ﾨ} �c?�N�%�~~@��_�ґ��켚�ܻ��!���}.���F��S�-�N�n;�(���������������7����Ӭ�>Zݿ���.���G��_S�:N�6�:��:�� ��ο�T��������o��:N���1����{G��������|��������=�.��K�S�k��  �  c�~��妿��)8���D�-p� �������~���vk�C+>�Kx�`:ؿ�����b��ʕ��/�� �0�H��Zt�����֌������,g��k:�����;ҿ��=q���?����I�eo�iȾW�����4���(�Ծ!��������.��Y�����5��`���&�y�S��n|�8��0������y?]�O�.�t��jƿ#5��Su��&�����xT)�45X��$��5���ax��=��-�X�z+��~ � #����Z^��l2�R�(c��o׾�¾.������v�ƾcN߾ƿ�#���h<��(l�蘿8̿ݽ	��5���b�����T���M5��%
y��|N�&��������Q��	��[Fӿ:����9��g������M���@���Au���J�=��=�*C���焿V�Q�.�*����
���־kož(J����ľ��վG��:��D`(��N���������b�1��R�E��fq�tM������0����l���?�����@ۿ򟯿s������;鿍��RJ�� v��̉�;���zՅ���h�*)<����3�տn���Px�t�F��$�W�
����!�׾9ʾ;�ǾѾV��C����v`7� �a�7c���y������8(�V���~��ˋ��8��V����I_��0����vʿ�?��W��<0ſ�� ��Z+��<Z�N)�����m�������Z��"-���&W¿�H����f���:�T{�z��L��FTҾ\Ⱦ�fɾ�5־�Y�m	�N�!�iC�_s��L���yϿ8l��`7���d�%}��=������ĥz�P�o>!���y����O������9ֿ �%;�Hi��0������
��W�v���K�{T�(�쿇簿����i�V���/�F������[�྅�ξZ�Ⱦ8�;X޾�O���(��q,��R��  �  �ׁ�����A���5��Iq�ת������MD����������j���/��� ��=ȿCU���bѿ��	�\Z<�tx�����4�����` ��,�����c��!)���kq����r���5�L����[þe��5l���X��R���)���8վj� ��!��[T�y
���̿B���@I�}���G���jq��tA��Gc��	��K�V�9w�������I����e����O�fم�W"���~���Y���ޞ�׽����O�Q;���Կ�G���Z�n#&��t�2�ؾ!t������퟾ K���B������Ț��H��1���k��墿�(翹s#���]�|/���g����������>�=bC�I/��ؿr��	�ſwQ����*�ߤd�����@ƥ�}����n��>ܗ��x�j�<�=��@㾿օ����J����� ����Ծa����2���8��������Ӿ����
�T�E�4����|��f����6��r��X���.��f���ӧ�����xl��c1��$�KL˿zd���rԿ�6���=���y��q��N
�����J���׏�u�e�v�*�� �L�Ĭy�6�<���m|��c�Ҿn���Z`��򖯾�?��%�Ⱦ��;9	��q*���\�7O����пv��	]K�-���H����z��3I���i��P��ɝX�=~ �����¿uS��������Q�4݆��&�������`�����xǆ�{�Q�9S�~�ؿ�{���ec���.����?Y龯�ʾM���ܯ��
�����оs6�k���8�s�r��I����!%��U_�$���=��*���މ��(Q���e����D�h���
ۿ#o��U�ȿ�J��V,��f��4���t��F6����������1z�<E>���������(��}�O���!�զ���޾i�ľj����{��ѹ��ײ¾a�۾� �p�&�I��  �  ����dÿ��Z�L��B��7���c4������xm��rG��gQ��/�F������ۿ)@ɿ�����1U��������|��������Z��7�������D>�)��&���R!y�l�3� ��6<׾���ͳ��HR��AИ��&����ž�M󾕖��XV�J+��ˋ޿��"�)�c�S���R�������H����ط������s��i2����ːпv�Ϳb��� �+�C�k��P���D�����q���7��&c����k��,)����X���^��O"��#��bHɾtb�����B����퓾b���a���<Ծ����.�7q��������7�Y�{�SƟ�^���p������H����#���B]�y ��b��˿��ؿ�Q��p@��с��P���м����U��i!��z���ffU�Z����Ϳ󍿣�J�ؐ�9afž6���u��r������I����þ����z�FE�@���'ƿo���HN����9�����ކ���"��=�����O<H��
��߿�N̿���f����V��э��|������{��,6���ݣ��d��C�?�P��d+������:�����&�&6þ�G���ԣ�>���@���͹�)y־@��&���^��n��n��k�$�v	f��ɕ�<����������	߸� ���r�u��p4�t��=�ԿO�ѿb����.���m�{T��~I������F���:?���l��I�m�lD+��H�1���ff�U�*������پۼ���?��׉������H��AK����4��"�5�q�w��f��� �:/9��U}������2���B���}��E������e�^�x�!��]�|ο�ۿ@����A������������t�������^ȭ��<���V�2��N�пЕ��\�O���������`Ͼ��������':��x��M���̾�I�݊��CI��  �  훈���ȿ����U��e���0���������S�������%���O����3�cϿ~�' ��F^��8���Q��ƙ��>���j���9Z��AI���7F�����8��Q|�	~3�����Ҿ#O��=8��r����ԍ�bo���������Hf�����W��1��"��A)�w�m�%l��⚺�J�������d���Z֢��~���9�����׿_EԿ�>�l�2��v����+M�����6���Vb��o>����u�)�/��ￌ���#�_��!��e��.�ľ�Ǧ�ѹ��Ir������J��������Ͼi&�Ґ.�7�s�q%���@��?��e��N��������`��\e������Ɓ���f�}�&������ѿ��߿���spH��v��t���,.��S��f���������^��H���ӿVX����K��^��8�|���Φ��� �������Ù�����f뾾��C$���E�>\��,�˿J>��W�{���߱����Ty��2���i[������P�j��D�RqҿM���!�7�_�� �����rl���m�����06���%����G�{h
�����R���ר:�V<����E����ǩ����u���dۤ�8/����Ѿ�) �:%�``�4u��}��#+���o��x��å��{���?������}ۣ�-����;����&ۿ3Oؿ�C���4��	x�W	���Q���������|j���G��xx��2����u륿!Hh�� *�4�*;վ���.إ�N��:@���Ө�Z����Q޾aD
�\�5��z�J������t�@��:��'̧�~���2���2������(E��v7h��M(�̆����Կ����U�I�42���7������r���s������������_���+sֿ���h�P����Qf����ʾ�g��ƣ��z��Ţ�i����pǾ@�4�W�I��  �  ����dÿ��Z�L��B��7���c4������xm��rG��gQ��/�F������ۿ)@ɿ�����1U��������|��������Z��7�������D>�)��&���R!y�l�3� ��6<׾���ͳ��HR��AИ��&����ž�M󾕖��XV�J+��ˋ޿��"�)�c�S���R�������H����ط������s��i2����ːпv�Ϳb��� �+�C�k��P���D�����q���7��&c����k��,)����X���^��O"��#��bHɾtb�����B����퓾a���a���<Ծ����.�6q��������7�Y�{�RƟ�^���p������G����#���B]�y ��b��˿��ؿ�Q��p@��с��P���м����U��i!��z���ffU�Z����Ϳ󍿣�J�ؐ�:afž6���u��r������I���þ����z�FE�@���'ƿo���HN����9�����ކ���"��=�����O<H��
��߿�N̿���f����V��э��|������{��,6���ݣ��d��C�?�P��d+������:�����&�&6þ�G���ԣ�>���@���͹�)y־@��&���^��n��n��k�$�v	f��ɕ�<����������	߸� ���r�u��p4�t��=�ԿO�ѿb����.���m�{T��~I������F���:?���l��I�m�lD+��H�1���ff�U�*������پۼ���?��׉������H��AK����4��"�5�q�w��f��� �:/9��U}������2���B���}��E������e�^�x�!��]�|ο�ۿ@����A������������t�������^ȭ��<���V�2��N�пЕ��\�O���������`Ͼ��������':��x��M���̾�I�݊��CI��  �  �ׁ�����A���5��Iq�ת������MD����������j���/��� ��=ȿCU���bѿ��	�\Z<�tx�����4�����` ��,�����c��!)���kq����r���5�L����[þe��5l���X��R���)���8վj� ��!��[T�y
���̿B���@I�}���G���jq��tA��Gc��	��K�V�9w�������I����e����O�fم�W"���~���Y���ޞ�׽����O�Q;���Կ�G���Z�n#&��t�1�ؾ!t������퟾K���B������ǚ��H��1���k��墿�(翹s#���]�{/���g����������>�=bC�I/��ؿr��	�ſwQ����*�ߤd�����Aƥ�}����n��>ܗ��x�j�<�=��A㾿ׅ����J����� ����Ծb����2���8��������Ӿ����
�S�E�4����|��e����6��r��X���.��e���ӧ�����xl��c1��$�KL˿zd���rԿ�6���=���y��q��N
�����J���׏�v�e�v�*�� �M�Ŭy�8�<���o|��d�Ҿo���[`��󖯾�?��%�Ⱦ��;9	��q*���\�7O����пv��	]K�-���H����z��3I���i��P��ɝX�=~ �����¿uS��������Q�4݆��&�������`�����xǆ�{�Q�9S�~�ؿ�{���ec���.����?Y龯�ʾM���ܯ��
�����оs6�k���8�s�r��I����!%��U_�$���=��*���މ��(Q���e����D�h���
ۿ#o��U�ȿ�J��V,��f��4���t��F6����������1z�<E>���������(��}�O���!�զ���޾i�ľj����{��ѹ��ײ¾a�۾� �p�&�I��  �  c�~��妿��)8���D�-p� �������~���vk�C+>�Kx�`:ؿ�����b��ʕ��/�� �0�H��Zt�����֌������,g��k:�����;ҿ��=q���?����I�eo�iȾW�����4���(�Ծ!��������.��Y�����5��`���&�y�S��n|�8��0������y?]�O�.�t��jƿ#5��Su��&�����xT)�45X��$��5���ax��=��-�X�z+��~ � #����Z^��l2�Q�'c��o׾�¾-������t�ƾaN߾Ŀ�"���h<��(l�蘿7̿ܽ	��5���b�����T���M5��%
y��|N�&��������Q��	��[Fӿ:����9��g������M���@���Au���J�>��=�+C���焿X�Q�0�*�������־kož(J����ľ��վF��9��B`(��N���������b�1��Q�E��fq�tM������0����l���?�����@ۿ򟯿s������;鿍��RJ�� v��̉�;���{Յ���h�+)<����5�տn���Px�u�F��$�X�
����#�׾:ʾ<�ǾѾV��D����w`7� �a�7c���y������8(�V���~��ˋ��8��V����I_��0����vʿ�?��W��<0ſ�� ��Z+��<Z�N)�����m�������Z��"-���&W¿�H����f���:�T{�z��L��FTҾ\Ⱦ�fɾ�5־�Y�m	�N�!�iC�_s��L���yϿ8l��`7���d�%}��=������ĥz�P�o>!���y����O������9ֿ �%;�Hi��0������
��W�v���K�{T�(�쿇簿����i�V���/�F������[�྅�ξZ�Ⱦ8�;X޾�O���(��q,��R��  �  H���B9���&ſ����4��Kj5�nJ��dQ�A�G���/�b���g߿�㬿e���υ��Q��7���L��*��5�ANK��TQ���F�w�/������,��4Ù��̀��4[�s�;�� �k<
�����ݾ�Z�C/�i��/��L�b�o�	ԍ�����[�Կ�����"���=��N�<"P��$A���%�?��n�̿�����C�����ۜ���ƿN
���!��>�H1O���O��4@�v�%�F�#�ٿD>���q���s��O���1�~A�G��Ic�W�ݾP�߾jq�ө�����K9�1�X�A~��W��>}��^��0���,��7E�~cQ��BM�Ru9�=���������z��x���l���橿oxڿ����$-�Y�F�yR���L��99�������T�˿�����
����j�<I���,�*��j�:�N����DG��G���*���F�o�g��@��E�����ǿwJ�������6���K�`�R��I�!	1�+��]�
寿�n��Wሿk��������s���7�|M�S��H�.A1�_���6����C��wX���jb�=�B��(����ص����7����7�
�d����7�+U��2x�����̯���ؿ-����$�r�?�/�P�02R��1C�/�'�����п�����N�����j堿%�ʿ����#���@�=Q�ܤQ��EB�I(��
���ݿ�s��ѩ��K�{��*X��!:�d� �t$��������ﾨ} �c?�N�%�~~@��_�ґ��켚�ܻ��!���}.���F��S�-�N�n;�(���������������7����Ӭ�>Zݿ���.���G��_S�:N�6�:��:�� ��ο�T��������o��:N���1����{G��������|��������=�.��K�S�k��  �  �֜�]����漿\�ӿ�ￋ$���s9�������d Ͽ�^���ꅿ��c�I�X��qj�80�������~ؿe- �yp�\��x��4��:鿺-ο ḿ�q��֙�y�����s���Q� d2��:�� �[	�����&��#C��d�@T���H��a����;���Ŀ~�ܿ����hp
��������)�h0��͓��_�{�+C]�t�[��w�ǖ�������.��&E�4���6�����߿�Iƿ�ڲ�0^��O���R���q�g��KF��#)���7�	�h3��b���/�!�N�3�p��U������Ĉ�������P̿9�濈��V�'�� ����1@޿셴�����:�p�)�[�
d�6���ˣ�i�˿C{��=k�0���U�p������\ؿ	��tD��!h�������P��mq`���?��.%������zr��6#�K^=��]��������a���^��1����KֿUN�'�}�V���N�����n�ѿfN��:爿��i�}�^���p�[���1���ۿ��\'�8I�U��#�����ѿ][��h��a���(���{��%Y�"8:�$?"�1/���p�%/��K��m�򡇿����2I������#Tȿ��࿅���4��n��8���	�;?�BſS���{ ���Xe��c��'��Қ�X��������1Q���`��A{ ���㿒|ʿ��[�������+���Up���N�r}1��^�L��n9�<> �wr7��V��x��܌��S��������Ͽ81�!������֞�^A�bvῸ����ד�1�v���a�w�i��i��०���ο�5������#�����	�d����ڿ��ÿ걿����(��:僿6�e���D�	*��@�G����ɡ'�R�A�C�a���������  �  �dϿL[ӿ�ѿ(EϿ=^Ͽ��ѿ�^ӿ��ο����⬿(r���u���L�73�85,��7�ѣT����UL���2���ſ�п��ӿ|sѿ�=Ͽ��Ͽ&�ҿ�UӿѡͿ��������K����m�u�G��O1��#-�g�;��E[����ĝ�����Yȿ'�ѿS�ӿOѿ<Ͽ�[п�ӿFӿ��˿��
䤿���{�f���B��\/��L.���?��a��2����������vʿ7�ҿLӿ3tп��οd�п�ӿl+ҿ��ɿ <��?c�������R_�>��-���/�F�D��Vi�������������!Ϳ.�ӿ�ӿ��п��Ͽ1�ѿ�HԿlRҿ�Qȿ����4:�������7[�>�<�R@/�]�4�ZL�\s��4��u竿:���.�Ͽ�"տ!$Կs|ѿcѿCWӿ�Kտ�.ҿ��ƿɲ��ʙ�����Z�V���:���0� 9��TS��~|�wb���ǰ�A�ſ-%ҿ�ֿ��Կҿ�ҿZ�Կ(ֿ3�ѿm�Ŀ"���ZN��~�z�e�R���9��\2���=��[����(���s����.ɿFԿ�	׿��Կ	�ҿ�Vӿֿ��ֿP/ѿǿ¿+���B'����u���O���9���5�5(D�5�c�T`������g���̿63ֿ��׿�Zտxӿ��Կ�;׿j/׿1п��������%����n���J��r7��a6��G�mj�0@��������s�οɠֿk?׿�ԿH-ӿX�ԿuX׿�gֿ��Ϳ�{��ݡ���ي�۽g��mF�X�5��8��L��q������Q�����пN;׿�ֿ�HԿ`Uӿ�TտB�׿��տҩ˿���� v��6؆��oa��B��?5��}:���Q���x�%��������kĿ0wҿv�׿�ֿ�ԿȨӿ9�տ]�׿��Կ�Iɿ�[��$P������[�$�?��.5���=���W�Oj���~���ղ���ǿ�  �  N�9��c���}$ҿ�ػ��ʪ�y������y�>�V��6�lM�UF�������qS"���=��|^�Ld������q���g���o���ؿ"����_��������	�6��ȿ�f�� с�	U`�C�Y�-�p�i��Cµ���߿�#����|�xr�<� �!��xPʿ����2��"w���쇿�n�� L���-��.�N�
��
��5�B�*��cH��j����O����I���೿j�ǿB(�9`���,�H��������	�M��Ӿ���ot�q�Z��^�Wa~�Z���9�ÿV��6��͛����;!
�i�����ۿהÿ|���衿�2���7��^\d��OC�Y'�+��w����E�6� [V���x����FS��?���(���Eѿ��쿸��L��i�T�� ��ؿ�Ү�������l�m�\�)�i�@���,ު��ӿ����+�������_��2��s�ԿZ�������Ҟ��ŏ�F�~�0z\��<�L:#�3Q�����7�O�(�=0D�)e��Ƀ�z
���좿j汿��ÿy�ۿV)���
����������K���H̿an����O�h�
Wb�� y�}������] 俥N�~6�7��K���	������οS(���7�������Gv� ET���5��G�����.��K���2��P��?r���ə��g����Ż˿�W忑J��I�|>����m��fM迏J��X�����|���b�;Df�	=��������ǿ�p�b
��W�Ou�A���&���E߿��ƿ�h��I��Ë��u�����j��I� �-���9�����#��m<�Y�[��~�������k���G<����ӿt5��(������4��e�'�ڿAF��R����q�fya�݄n�[���>��W�տ|������  �  �hQ�/�I��3��������¿]����M��̳`��@��[$�>��z���⾌�۾��徬O��n��I*�DG�si�P���	����̿ �����9�"�L��Q���D�U�*�,&
���տ�|������&���eݗ�T���{n�����v:��M�Y�P���C��*�V��3�8����&��пz���U�6�6�*��R'������޾�޾1�쾞
����e�3���Q���u����ZV��3oܿ3�	��'�m[A�#�O���N��=� ��B���ÿ�嚿�P��҉��`����Ͽ���n'���B���P��mN��<�Iw!���I�ҿ�Q��*��wo��tL��O/����P���쾏���M澇k��@-��$��G@��c`�����N��r��$i����L�1�ǴH�dSR��fK�c5�}*�h��+���&���ꇿ(Ƒ���������2�K�I��R���J��R5�gP��>����ſ�D��w���4f���E��	*�l	���#"B��6�&��ޜ��0���M�=�o�����>���/п���/v�zz;��N���R��{F���,��#�ڿ䯪�܏�` ���4��=�¿m������M�<���O���R���E�-��-�ji濷ٹ��N�����O�]��?���$�\E�����-�h@�����"���!��;���Y��+~����z�������)��xC�R���P��=?�&5"��E��!ȿ�(��[�������%�ӿz���O)��`D�=�R�� P��>� $#�7M��ֿ���Z���H�u��S�L�5�/�ג	�W���i��/�l��u��O`*��E�+�e�]M�����h�¿������83��J��S�7�L�u�6�Lh�D�����퀖��=�����(Ƴ��G�����3���J��  �  ��������R�m�(	B����z�ܿ*P��v{��bF��s!�T���~�ʾ6�|��l���Xо���]�S�(�r�P���Q��Kq����XL�vtv��Z��Č��]����d��[6�G�	�3�ο����{���F������!���P���z�u��Z������!0`���2�8'�Hȿ���g��)9��.���Ûܾ,žu긾T=��gþ�Dپ ������4���a�T��-^��n���-��=[�������"0��S~�u�U��&�F���g���z��^ ��\ɿQ0�y,1�!�_�_��$����}����z���Q���#��V��𵿰Љ���W�>�.����e��Ӈ׾ľ�������ەξf��˃��!�,=E�p�w�P���׿E�#�=�|Sj����>b��nۈ��*s�rG�÷�)���ܳ��r��gk��u�ݿ���B��n��̇�ѩ��x����;o��iC�4���߿���H����K�<'�XW�H�񾐫־�ǾG�¾�2ʾ��ܾ���5���/��W����β�����V �wN��0x�8;��N����L��yxf��b8�R���;ӿ<ڬ��쥿}c��������#�#�R�\�|�����_n��y���FRb�h�4�B	��>̿i��tp��`A��> ���L�쾋Lվɾ�hȾ�BӾNu�+�����*�<���i�Qr��	�ſ]���/��X]�v��Pь�wA���;��E�W���(�
���u�¿!æ�@��75ͿE=�g)3�-�a�I˃��o�� X����|�*{S��%�T����P��'/��ڋ^��5��f�����來cоcȾ!T˾�ھ�����;�&���J��(}�d���ڿ�b�+?�r�k�YȆ��
������mt��RH�C����L4���Ť�4�����!��C�p��O���  �  D��в��RC��'�m��f2�l���F���C�w�=�<���B��Ǿ�b������f��}:��=糾k�ξv9��M��J��2��N���@o	��V?��S{������������p��ˣ���`�X'�q��*�¿�й��ٿ$��F����E�������s���1���y���Y� �M��!4��]�f�J�-�Ϋ���߾���������������,騾	���=۾�>�9�(�7�^��1���	ٿ� �p!S�VN��@���q����������.��"xL��&�r�߿�����O�z4!�d�Y�����@���_���U��}��.#���LF�OC�apɿ�#���{R�	S!����׾����q��������妾�w����ʾj��.����;�_0z��h��&��`-�r1h��ߐ��y��Z�������Ö���u�|>:�Kg�0ѿ�Y��q�̿>��$4��(o����P��� ��c������Po���3��c �����C\��'-C�H������Ӿ�0����������ڰ�i����ܾ���g�!��Q�w���.]Ŀ�-��A��}�����������gb��&���Ӫb��#)�on��wHǿ�8��#޿�R�EH����4���s*��I����D��ኋ��\��5"��$濾[����n�96����&"�DϾiѺ�����j ������9̾Sv뾹`���0��g��O��w-ݿ�5��9U��[��G���Ǯ�z��?���B����N��P�����^��-�ÿ+��J#���[�-���"u��я�����0U��������G�O����̿����,Y�h�'�[������Ǿ+Ƕ���������龾��վ9���&���@��k��������d.���i�刑��"���M��<���Ec��
�v��n;�u�	��lӿᬼ�^�οL�<5��Dp�E�������  �  �����J��A���R���.I�����O���냿8�<��0�2޾����ʠ�8q��=$��Aq��i��\J����R �r�J����T�п9��WX�����5��G����|���X���=�����a<�K^��տG�ʿ\���"��r`�����:*������������ԝ�1dw�P�3�"��� Ȩ��[k��*���dо�ï�xc�����o����̚��ݬ��˾k���*%�eb�!���k-��,�jyo��0���z��u���5�����Li����g���(�Kh���q̿E�ѿ���S�5�'[w�lƝ��"������5���P��T
���i`�ū��ڿ�ҕ���S�$��8���tǾ{
������Ǯ��|`��� ��`@����߾���Z�9�Я��	:��E����B�4��S ���ս�!:��]�����������R��t��
濣;˿5��U.�	kK�ׇ�$��������������)���"���J�����¿S���(B����`�龳�þo���C����}�����k���mw̾��d��8�Q� ���R	Կ9���Z���������f��M��b>��l�����>��
��ڿ4gϿf����%��b�Nړ�9A���4�����l�������y�'�5������﬿)�s�3�-D
����� ��V����L��,Ȣ����������۾L���S-�m�j�iݥ�WQ񿇬.��q��>��쉷��.��7G��n��}��j�K�*����j�пu'ֿ,���7�:hy�8�(��������*��{���b�@\!���ݿM0��<�Z�"`#�"\ ��CԾ�����㨾 �������q��Dnƾܱ���$?��M���ӻ����D�Ñ���ȥ��}������ZD��J>���;��X�S�����]� �Ϳe�|W�ڐL��f���������  �  ^ߪ�����ׁ��8g�HY,����1���h�D'��0����ľ��~��G���b܀�az��-A��RV����ξ}�ށ3��{��ʵ�����'9�ot����Ww��b�����,����Z�s�!���ϼ�[ ����ҿ��Z/@��z�Z����U��w-���چ�mvS��9���ֿz���P��w��澧���Ƽ��9Ê������=��v^��e-���h��1�h�RFH� ����Ϳ\M��L�P���{ ��{j������ެ���r���kF���c�ؿV3��ʡ����N���S����8���@���ѧ�[����M{��@�|�	��]��B���Y�;��,�gQؾ�����������8e���ƈ�}�7����ƾ ����%�?�c��P���꿻'�h�a�~*��Ga���F����Ш���n�>�4��:���ʿx���.<ƿ�����.��Gh����s3������P?���1��o�h��-�C���驿�>n�$�,�ǫ��о�}��#J��$ɏ��1��:��E$��
|���@ܾ��	`:�u���C��#w�E�:�+*v�ŕ�QX���w��O
��ɰ��\�k$�����+��lb���U׿���t^B��|��o��/���M2��?�������U��R���ڿ*:���ZX���5�����Ⱦ��[(֒��a�������V��C�ľ�L����sP��+��ҿ�`�L�N��Ǆ�����y��g���Q��������H������ܿ1���C뽿�1�c���U�����%���"��]����q��Q�|���A��4�\����S��f�B����{P�S޽��~���Ɨ�t`���z��va�������Ѿ/Z��Z*���h��ꤿ���cf(���b��ҍ��	������4��GH����o���5��g���̿趿H�ȿ	���/��di�ؑ��^����  �  0����}���P��bs]�%�e�������e���&�|���ρȾ���q�������c����V���L���n��8�Ҿ���2�#x��󰿀7����1�;j�ax��BG��S;���@��ރ��	Q����|g�@���殿<̿i}��k8��#p����Gw��aʢ�EW�����J�*f�>5пA���1N�)��,��M���ן�s���0y�����KJ��E��jn��xU�p����F��G���ǿ����GD�)|��A�����EZ�����tv��X>���&�ѿ����<��;@޿U���J�G���w�������������p��D8�@�����3���#�:�����۾�+����-f���(������'������ʾи��%�� a�����P㿊� �YX����Ya��]���}��+p��߽d��-�V���tĿ����vK������a�'���^�����2���1���-��� ����^���&��]��ե�+k��h,������Ӿ�����K��Ĝ��x���;�V/�� �����߾d��m�9�X�~�cl��� �;o3��k�[V�� (��N"��?1���ل��S������� ����F����п��	���:��Pr��������^ݣ��h��x����L�A��`Կ�%���nV�@ �:����̾ ����������	)��Uo��4n���Ⱦ��W"��N��c��)�˿��#^F�xB~��O��+���j��I/���4x��~@��F���տ7U�������z⿳g�y�L�z���c���ӣ�p������Dr�y�9��K�y�����j�A�Ϩ����r���Ď��]���G$���J���]��˵� �վ����]*�V<f��0��G��[�!��kY�V��	�������!����\�e��.�j� ���ƿ#Ɀ۝¿�!��%�(���_�#y��A����  �  �S���&����p�P#C�����|տ��$_�(�3y�6�վ����!f������e��r����f���"���`߾!�
�n�2�� o�~���0	�!����M���y���������q��;�g�,m8�8�
�+GϿ맿�ʠ�Fҹ�~���@#�IIS�_~�ɶ��f���u����b�f3���?4������f�J�;��IT���$ʾ�L��]K��}\��ݑ��Ǚ�`���,ƾ�Y�L��*D���������A ��-�ӈ]��ׂ�a��Cy������eX�T(������V��z���QX��F1ɿA��3���b����b���Ì��s~��S�T{#��xￄƫ��y�H:�#2�]y�0�¾�;��6����򕾠��������4���ؾ̺���&��[�`��R�Ͽ*}���>��<m�R=�����������v�׌I�T��q�Oz������c��t޿�5�TD��lr����1���։��Rr�}�D���86ؿ����a�d���-��	���@���1������ع��.)��TG��FȾ��쾓[��9�A�u�32�����B����O�ܠ{��x������a��,�i��s:����ӿ=��a$��?/������n%��uU��D��ˍ�d������d��75����_ÿ������R�B�"�����eھ����>w��̂��w���쩾ZϺ��F־$����p�EXL�G����0�� U�}�/�!�_�����"�������+����Z�y*�������¿�����bͿ��5�x�d�ԅ�����֝������PU��'%����"��G��+�@�f��]x���Ͼ��������@�I���(��cþ}㾚	��&,���`�5���A2ҿV���@���n�N���c������8�w�x�J�~>���;ҵ������B�����hV��mE�*}s��x���  �  s�f�E
]�c*C�;  �����ƨ���*��n\���/�������nϾ����2���譥��쫾U(���T־�(�����=�8���h�u��<ȿ��](��J���`��Uf��X��t;����v�ʛ���4�����������˿g9�~+��:M���b���e��V��<8�����⿲���x��RL�t�$������p;Ǿ@����ꧾ�Q��dٰ�pKľ��Ὰ=�� ���F�O}�y�����ۿ���#B4��:S��d���c��8P�.t/��
���ѿ�����f���6����;}߿���K�7��NV��f���b�t�M�X�,�K[��LϿ¦��@4q�a?������G޾xKþ�K��dC���d������-�Ҿ���/���i/�J\Z��勿D����������@�f�[�Z�g��`��gG�$�����¿�����̍�a瘿'ͼ��I��� ��D�Uu^�*h��k^�[�D�܀!��C���b��s㐿��a�4`5�����	���ھz]þ����b ������ɾRt�AC��J�$�?�^�o�������˿����*���K�.�b��h��Z��a=�+��g���Ѵ�{�������e��Bп�e���-�eO�ٷd�g�g��9X��\:�s$�*�=��@����T�X�,��6��7���o׾��¾���Tu������tԾ���5[���(��$O�Â�sͩ�i�߿���M[6�^VU�O�f���e��ZR��1�6B��5ֿ�ǧ�����i��n����㿹|���9�{X�R�g��}d�@fO��z.�H
�Z�ҿ�����w��E��K"������a�Ͼ ���:?������	Ǿ��ݾ����	�.�4���_����WW��u����N�T�A�']���h��ga���H�wW%�<� �#�Ŀh���� ��"5����ل��21!��'E��z_��  �  H?,��&����E��.Aοr���r��;h��DF��A*��T�/���e޾8�˾K�ƾ�ϾCn侀���w��F0�!iM�21q�����jv��5ؿ͂�k��V�(���+��!��A�i�濇�������:t��Ml�� ��)�пC�l���)��+�C�!�������v��� ���MJ���\��<��X"����]򾀺׾=dɾ$�Ⱦ�gվ;��wG	�s}���9�i}X��M��m��? ���_翗>�ǡ��#+�f�)�`������eտ(���l��Rm�Rfq�av��F���BI�r�
�f[ �V�+�i*��&�?��o޿ab��Sᓿ w���R��45� ����H�*�վ�D̾)cоt�ᾶ?���>��*�1�F���g�'��#���j˿�������%��0-���'�E��J��l�ƿ�����f��lo�������������������v&���-��|'�e�D��%�п�9������J�m�b�K���/���*��N���׾L�Ҿy�۾HD��	��#��7��GT��x��s���ﲿx�ۿ�<�Z�\j*��-�<�#��(���h���=ޓ���|�^�t��M���@��oYԿ7�y��wC+�z�-��#�������Ŀ\"���n����d��E���*� ���H����։پc�ؾ��_���:_���'�ݲA�Y�`�-������&���뿀W�@�!�AA-��,��	����u�ٿDZ��������u�r�y�a��������%�a���&"���-���+�D���7��g�ѽ��->���4~�|Y���;�N�"�\?�����O��@ؾ�ܾ}U�;�ƻ��E0���K���l������G���ο�������&��.�,�(�j8�A���Geɿ���q�T�s�*́�w7��I$Ŀ ����&z'��  �  D���`h�d�࿲Lʿ=n���t��+>��h���:�u�Q�Y���<���!��6��$���B��'� �%���'��lC�d`��{�V���P��<��G0��ߝϿDc� ����ʑ�cf˿@#��]>��Y�b���E�ޔ@��AS��?|�`o��������ۿӈ�Z��H;���ٿ� ÿf=�����bE���σ�g2m���P�B�3��]�����������c����C�0�HM��i��H������2替#���R��A"׿};뿸���1���w޿�k���֞��π��rV��DA�1D��^�H7��4����Hȿ������h|��yI�r ӿ�b������#����ٌ��L��~e���H�\�,��!�خ�1	���| �tD��V"��=��Z��\v��0��U�������� �� �ɿ�L����������N׿�F��c9���Au�Q���C���N�<�p��������ŝԿ���ߛ���+��D}�`ͿZ*��-�������s��LD{��l_���B�c�'�� �S���� ������U2.��J�)g��]��E���ʚ�s�����ӿy���[��`���x7�.)Ͽ���L<��k�wEN��I���[��i��G���6E��������9������޿�9ǿCo��*ա��i��
�cu�\�X�
<��w"�
(�������u������8��dU��r�_���ْ����F(��Z~ĿRSۿVq￉��������x�Ŀk������^���I�hBL���f��!���|����˿�1��J��������@Xֿ^���]R����85�������l�{2O��,3��]���
�l���[�J�q�'�j�B��|_���{�mΊ��K���8�������I̿m��x���ʵ���e���ٿqɹ�Ю���z�r�U��lH��+S��u��L��.��H�ֿ���  �  =߰�<���,���d_���p��l��B���≰������U��;��V�ۣ4����bp�V	#�:7;���^�SV�������è�_�����س�sj���Բ���������d���L���.��=Rx�h*P�L0�����E�0l&��@�=�e�����盿W���y!��}������}s��1��ش��4�����H���\ٍ��kq��@J�>x,��%�.A���)�JOF�C�l��w��c���c�������1̴��2���;��A��Vô��`��9��������#���j�b!D�<u(�#��[����-��L�QLt��`��8��������x��г��.���y��kǵ�:���O��Z���򿇿�e��A���'��n�q� ��4�pU���}�ړ�ť������X��!+���}���0��m������������٩�ʄ�����`���=�c&����I�$�]�:�q]��5��#����
��j���lg���������+���˶��V���C��q`���"���b��B�[���:���%�����I)�V�A��\e�᥇����0��ޕ��i��T���㵿pK��L�������ﲿ�Z蔿R��
X��8�M�%���"���.�:KI�/qn��O��K3���?��<i���O���跿����yb������X�����Ϥ��쑿�y�!ZR�B�4��7$�ER#�8�1��bN�F�t��Ӣ�VͰ��η�X츿RX���f��*q����������+5��ޡ��\���vr�SL���0���"��$�}�5�aFT�p�{�������'���h���Ӹ�v)�����׷�&������g��c��������k��NG���-�
l"�+�&�(`:�׮Z����O���m��"%����ø�w��ж��Q��nL��^2��v����1�����e�:�B�!+��m"��o)�0X?�,ea��Q��3�����  �  �Y���딿�P��w�����˿2�ῗ򿙺�����cп\������Ii�{�H�sy?��4N���s����4���׿���Z��0�ￌ`ݿa�ƿAO��'���G��҅�q�$\U���8��+���	�������B%��5��],�ڋH��ge�y>���̌������5�� ޼�܏ӿҙ迋3��w���⿈$ƿ����Q����\�CnC�,B�ȞX�y���۠��p¿@���ƫ��vc���տ���+���,
�����r��h��`K�9/�T�lt��C��a����*�B��$6��S�n�o��������#,������H�Ŀ��ۿ����0�� ��j"ۿ��������{���S�p�B�IsI�]�g�A���x��2�ο]�$������	�пfù����%R��B����~���b��E��9*�������x���������)(��C�.�`�q�|���D������J��OPο2��O����t��Q��3ӿ�y��a�Wro�M�N��E�,nT��
z��,��i~��kaڿ�O�������|�࿂#ʿ`Ǵ����� ƕ�P\����x���\�'@���%�u�����؊�Z�����f�4�Q�J�m�*���c�������r��n����׿��RW�����$���7ʿ)���љ����d�>�K��"J��`������椿t~ƿ�俥���5���"��ڿDÿ/'��=��\)��ߩ���p�"�S��a7��������������#���=�'UZ�V�v�ތ��1��g���X��rRȿO&߿'����,��jf޿�:��Wɝ��ဿ�Y��H��XO�׍m�t�� B��AfѿW�	��������迖�ҿca��ﮩ�����R������!�g���J�0/��e�HD	�"��G/��]��w,���G���d�<C���  �  <j�f��ra���п
���x.�{�&�<,��b$�R&��w����̔�۰x���j��P�������ǿ>��O9�[L'�9,�z�#�Շ������Yǿ�#�����n]b�ڛA�XY&�E�[���2۾̾ʾ۴Ǿ�[Ҿu��d	�
��E5��S�Xx���������߿�}����+*�a7+�>)�z+	�Z<޿ F��=����|p��|n�������5sؿR�L��q*�5�*����m�	�}��͹����:�|��_V���7����'��Z���*ԾCOȾ.%ʾЇپ4)������$�J�?���_�:��\b���ÿ��J}���"�Ca,���(�>���IEο䡿�ꃿj1n��3x�򶒿�]���8��[���#�p�,�^�(��d����x׿�5��o=���r�FO�1�2���D}��-뾄�־�gϾ��վ[[�B�͗��0�o@M���o�(���"���eӿ�� ���/&(�s�-���%�a���Z�a俿	ʗ�O�~���p�oi�����0�ʿ(�������(���-��%�SE����<�ʿ5���W����oi���H��-�6��؉����]�ھ�ؾ���0����v"$��=��[��o���������Y�ߕ	�����<,��E-�5!��4��K�RR��o��Y�x��v�{�����D~ܿ�X���|,�/�,�� ������ ���|雿.�����^��$@��E&�_A��%��My�@aؾ}�پ5��!������+��F�[�f�F���������ƿ�u�,�x$��.��*�>������cѿ����w��,t�C~������;����ߺ���$��@.��C*���1]�ڿױ�������w��T�A�7����v
�&����D�ƭؾ��޾L)򾀋�(����4� AQ��  �  eF_��B�����L��,,"�W�D�^�H�f��\�VA�����2��᷿�c�������¿M; �3%�E.H�`�c{f���Y�M�=������l.���-���6T��-*�����뾟l˾
5���㨾a���Ӑ��Xn��0Iܾ��}���?��s��T��_�ѿ��	�-s.���N��'c�_ee�g�T���5�h��ܿ�ߩ�W���B1������Shտ�E��1��Q�
cd��Jd���Q��S2�l���Wؿ����y�GD�9��8��l�߾�¾���3=������B��#�ɾku龆V
��'��+P�-���r���-��k���:���W��pf��<b��L���)������ɿ|}��1���dz���J��a뿒e��>���Z��^g�,�`��OI�5'���[�ƿ�����Ti��:���,> �&�ܾ�<þ ܳ�}���J��8¾E�ھ*������=7���d�e���^��
����#�	JF��m_�`h�{]��pB�+@��)���⺿�k��*Ď�I���ſ���(�&���I���a�y1h�#�[�r�?������|��������F[��Z1�uf�<���G�ھ��ľ�۸��涾����Ѿ����	��=$�T`H��{�����pֿ���0�.Q�T9e��sg��V���7��o��$��魿���c9��ཀྵ��qٿ2K���3�_�S�bmf�xWf��S��e4������ܿ#B�������L��,'���D��Ӿc.��l0��;W����þ�ؾi��Az�3�.��W��h��ϱ�Ç���.<�BoY�+h���c���M�_~+�MN��Ϳ΀��Z����q���:���E���~?�c\���h��.b��J�u�(��@�2JɿZ>��ȗn�CR?�����R�Z����̾V^�������P����ʾf��,�S���=;��  �  ��b�"����tٿx
��E��;s�~ω�vT�����+�n��m@���y�ؿ���ї��V?�����T��d:K��w��*���/��j����i�*#;�*+�	ʿ�����T�XC!�h����Ͼ���^x���$���N��Hݗ��:������)��{u��\;�:�{��=��t$���%���U����~��������VE`�k0����m�ƿ���ͼ���"������+��[�����ߍ�ȍ����.[���*�{���]����<��$�@���h:�M�þH�����lꑾ(��	㜾�ǯ���;F#�����^EO�����8}ÿ4���)6�m�e�Z������v��)�|��%Q�-8!��������n���y{��r�ӿ���p�;�7�j�Ɯ��^����y��v�x�^&L�����Xz���n���3�����w��6�������%8���9���ѩ�A�����Q
�F�/�BGh��y��6ܿqi��1G�͖t�5}�����U��7Hp�d�A�L���ۿ��������O����F���L�ۗy�# �����\��ߵk���<�"��5�Ϳu���d�[�7m(��P�#�޾cP��c	������x���F��Vط���Ѿ�h��<����C�*9���{���^��c�'���W�/������������Nb��r2����_�ʿ�����Ħ�
+ſ����-�N"]�������KΎ�U����]��-�I �D͸�m��GI��f����xmԾ����==��Pǡ�6����"��}���d8ܾn/��$�_V������ƿRk	�M�7��5g�e�������E��^~��R���"�L�����������t����ֿ��==�3Kl�3J���M��v ��<�y�'sM�am�6����i�s���8��������n˾\_��/���{���=��Ӗ����Ⱦ+p��c���3��  �  ��i�Ua���Y￈�(��`������>��.����ƛ�����FUZ���#�!��y%��������Ŀ� ��i/�N�f��8��J����[��=��8I��OT�f��*ݿ4ə��Y��2��B�¾o���m���K-�����!�����������۾���͠<�0���:(�����M;�Is��
��]������b���!��G�V���"ۿ�E���-��M�Կy��|�A��-y��C��Nϡ�š��8���8y��'A�	�N�ÿ�����C�g����HL��/�������#��]L��gL���S���#�����?i��0S�����'տs���2N�v����~��M=���%�����ٙm�3�5�y��^�ʿ�����	���P�S�"�T�z���d���<ˣ�e�����C�g�6�/�����~+����v��f3�/���׾�ĳ������j��es���!��w���Y����Ծ,\�� /�,mo�;#��+���)�z�a�oP�����#3��Dz��y���.�[�`%�'��0��ƒ����ǿ�'�o�0��hh���߃���3�����J%����U����e��IF��X�`��Z&�i� ��`Ѿ޴���>����Ϟ�������~�þ��b��cE�>���{e������=�y`u�������������g��_���J�I�M��s,߿wN���5��g�ؿ���ŎC�W4{��G��MԢ�Dˢ�@��J{�~;C��'�z�ǿ�����]K�i��e���ƾgE��̜�P��Ж��~��:0��ǩξl���x_"�X	Z�v��ؿ�<�3�O�?����R�������d����$o��}7��@���ͿŐ�����#H�� �
IV�$V���6���t��]���?P���i�O�0����α��&|���8��[��Q���ER��횾E����$��棥��຾�Bݾ�m	���2��  �  V9m�Y�������#}/�ԅj�����X���ݪ����i����c�^�*�zI����������U�ʿvo�/�6���p����B˥����F���H��H^]�+#��q�X���\���/2�]����f�����._������;���g镾_	����׾}��Ŀ=�`߅��������A�B�N%~�C���/���ө���� 2���FP�E���⿄����f�� ܿK���I�������X������|0��.qI��n��ɿ�&��<oD������ܾ}E��뗾)ֈ�Ob�������\��<��1����v��JU�G˗�� ܿ���'W�ی���`��*���gP���Z��U�w�R�=���
�]ѿ馴�B���`�� u%�^�+���Lk��]"��v=���	���
r�U�6�����ϳ�Ԣz�-�3�g����Ӿ����H���u���Ѱ���L���ܘ�K=���-Ѿ�$��S/��r�Of��X�����0�t�k������������(r��V���sJe�x,��R��jſϚ����Ϳ!���B8��~r��M��$���S���s���$���_���$�p���Ԡ�c�0<&������u;����A���.���Ց������w���¿�h达*�t<F�����ſ���E�W��V����7���ڪ�0���6��JNR�9��������n��"�zO���K�5��
��O��-��|��29���K�<���Ϳ�U����L��5�3R�}�¾u/���☾6-�����׊������ʾ�����"��"\�g,���Z߿�8���X�;a��4��If������#���y��?��O��YԿܢ��ĩ¿�����&��s_�H=�����I̫��������`Xs��8��I��r�����(29�3��V$޾���I�����x��N������7Ķ��~پ6�:S3��  �  ��i�Ua���Y￈�(��`������>��.����ƛ�����FUZ���#�!��y%��������Ŀ� ��i/�N�f��8��J����[��=��8I��OT�f��*ݿ4ə��Y��2��B�¾o���m���K-�����!�����������۾���͠<�0���:(�����M;�Is��
��]������b���!��G�V���"ۿ�E���-��M�Կy��|�A��-y��C��Nϡ�š��8���8y��'A�	�N�ÿ�����C�g����GL��/�������#��\L��fL���S���#�����>i��0S�����'տs���2N�v����~��M=���%�����ٙm�3�5�y��^�ʿ�����	���P�S�"�T�z���d���<ˣ�e�����D�g�6�/�����~+����v��f3�0���׾�ĳ������j��es���!��w���Y����Ծ+\� /�,mo�;#��*���)�y�a�nP�����#3��Dz��y���.�[�`%�'��0��ƒ����ǿ�'�o�0��hh��������3�����J%����U����f��IF��Y�`��Z&�j� ��`Ѿߴ���>����О��������þ��b��cE�>���{e������=�y`u�������������g��_���J�I�M��s,߿wN���5��g�ؿ���ŎC�W4{��G��MԢ�Dˢ�@��J{�~;C��'�z�ǿ�����]K�i��e���ƾgE��̜�P��Ж��~��:0��ǩξl���x_"�X	Z�v��ؿ�<�3�O�?����R�������d����$o��}7��@���ͿŐ�����#H�� �
IV�$V���6���t��]���?P���i�O�0����α��&|���8��[��Q���ER��횾E����$��棥��຾�Bݾ�m	���2��  �  ��b�"����tٿx
��E��;s�~ω�vT�����+�n��m@���y�ؿ���ї��V?�����T��d:K��w��*���/��j����i�*#;�*+�	ʿ�����T�XC!�h����Ͼ���^x���$���N��Hݗ��:������)��{u��\;�:�{��=��t$���%���U����~��������VE`�k0����m�ƿ���ͼ���"������+��[�����ߍ�ȍ����.[���*�{���^����<��$�@���h:�M�þH�����kꑾ(��㜾�ǯ���;D#�����]EO�����7}ÿ3���)6�l�e�Y������v��)�|��%Q�-8!��������n���z{��r�ӿ���p�;�7�j�Ɯ��^����y��v�x�_&L�����Yz���n���3�����w��7�������%8���9���ѩ�@�����Q
�E�/�@Gh��y��6ܿpi��1G�̖t�5}�����U��7Hp�d�A�L���ۿ��������O����F���L�ۗy�$ �����\��ߵk���<�#��6�Ϳv���e�[�9m(��P�%�޾dP��d	������x���F��Wط���Ѿ�h��=����C�*9���{���^��c�'���W�/������������Nb��r2����_�ʿ�����Ħ�
+ſ����-�N"]�������KΎ�U����]��-�I �D͸�m��GI��f����xmԾ����==��Pǡ�6����"��}���d8ܾn/��$�_V������ƿRk	�M�7��5g�e�������E��^~��R���"�L�����������t����ֿ��==�3Kl�3J���M��v ��<�y�'sM�am�6����i�s���8��������n˾\_��/���{���=��Ӗ����Ⱦ+p��c���3��  �  eF_��B�����L��,,"�W�D�^�H�f��\�VA�����2��᷿�c�������¿M; �3%�E.H�`�c{f���Y�M�=������l.���-���6T��-*�����뾟l˾
5���㨾a���Ӑ��Xn��0Iܾ��}���?��s��T��_�ѿ��	�-s.���N��'c�_ee�g�T���5�h��ܿ�ߩ�W���B1������Shտ�E��1��Q�
cd��Jd���Q��S2�l���Wؿ����y�GD�9��8��k�߾�¾���2=������B��!�ɾhu龄V
���'��+P�+���r���-��k���:���W��pf��<b��L���)������ɿ|}��1���dz���J��a뿓e��>���Z��^g�,�`��OI�5'���]�ƿ�����Ti��:���-> �(�ܾ�<þ!ܳ�}���J��7¾D�ھ'������=7���d�d���^��
����#�JF��m_�`h�{]��pB�+@��)���⺿�k��*Ď�I���ſ���(�&���I���a�z1h�$�[�r�?������~��������F[��Z1�vf�?���I�ھ��ľ�۸��涾����Ѿ����	��=$�T`H��{�����pֿ���0�.Q�T9e��sg��V���7��o��$��魿���c9��ཀྵ��qٿ2K���3�_�S�bmf�xWf��S��e4������ܿ#B�������L��,'���D��Ӿc.��l0��;W����þ�ؾi��Az�3�.��W��h��ϱ�Ç���.<�BoY�+h���c���M�_~+�MN��Ϳ΀��Z����q���:���E���~?�c\���h��.b��J�u�(��@�2JɿZ>��ȗn�CR?�����R�Z����̾V^�������P����ʾf��,�S���=;��  �  <j�f��ra���п
���x.�{�&�<,��b$�R&��w����̔�۰x���j��P�������ǿ>��O9�[L'�9,�z�#�Շ������Yǿ�#�����n]b�ڛA�XY&�E�[���2۾̾ʾ۴Ǿ�[Ҿu��d	�
��E5��S�Xx���������߿�}����+*�a7+�>)�z+	�Z<޿ F��=����|p��|n�������5sؿR�L��q*�5�*����m�	�}��͹����:�|��_V���7����'��Y���*ԾBOȾ,%ʾ·پ1)������$�H�?���_�:��[b���ÿ��I}���"�Ca,���(�>���IEο
䡿�ꃿj1n��3x�򶒿�]���8��[���#�q�,�_�(��d����x׿�5��q=���r�FO�3�2���F}��-뾅�־�gϾ��վZ[�B�˗��0�m@M���o�
(���"���eӿ�� ���.&(�s�-���%�a���Z�`俿	ʗ�N�~���p�oi�����1�ʿ)�������(���-��%�TE����=�ʿ7���X����oi���H��-�7��ى����_�ھ�ؾ���1����w"$��=��[��o���������Y�ߕ	�����<,��E-�5!��4��K�RR��o��Y�x��v�{�����D~ܿ�X���|,�/�,�� ������ ���|雿.�����^��$@��E&�_A��%��My�@aؾ}�پ5��!������+��F�[�f�F���������ƿ�u�,�x$��.��*�>������cѿ����w��,t�C~������;����ߺ���$��@.��C*���1]�ڿױ�������w��T�A�7����v
�&����D�ƭؾ��޾L)򾀋�(����4� AQ��  �  �Y���딿�P��w�����˿2�ῗ򿙺�����cп\������Ii�{�H�sy?��4N���s����4���׿���Z��0�ￌ`ݿa�ƿAO��'���G��҅�q�$\U���8��+���	�������B%��5��],�ڋH��ge�y>���̌������5�� ޼�܏ӿҙ迋3��w���⿈$ƿ����Q����\�CnC�,B�ȞX�y���۠��p¿@���ƫ��vc���տ���+���,
�����r��h��`K�9/�T�lt��C��_����*�@��$6��S�k�o��������!,������F�Ŀ��ۿ����0�����i"ۿ��������{���S�p�B�JsI�^�g�A���x��3�ο	]�%������	�пhù����'R��D����~���b��E��9*�������x���������)(��C�+�`�n�|���C���}���J��MPο0��N����t��P��3ӿ�y��a�Vro�M�N��E�,nT��
z��,��j~��laڿ�O�������~�࿃#ʿbǴ�򄣿ƕ�Q\����x���\�)@���%�w�����ي�Z�����g�4�Q�J�m�*���c�������r��n����׿��RW�����#���7ʿ)���љ����d�>�K��"J��`������椿t~ƿ�俥���5���"��ڿDÿ/'��=��\)��ߩ���p�"�S��a7��������������#���=�'UZ�V�v�ތ��1��g���X��rRȿO&߿'����,��jf޿�:��Wɝ��ဿ�Y��H��XO�׍m�t�� B��AfѿW�	��������迖�ҿca��ﮩ�����R������!�g���J�0/��e�HD	�"��G/��]��w,���G���d�<C���  �  =߰�<���,���d_���p��l��B���≰������U��;��V�ۣ4����bp�V	#�:7;���^�SV�������è�_�����س�sj���Բ���������d���L���.��=Rx�h*P�L0�����E�0l&��@�=�e�����盿W���y!��}������}s��1��ش��4�����H���\ٍ��kq��@J�>x,��%�.A���)�JOF�C�l��w��c���c�������1̴��2���;��A��Vô��`��9��������#���j�b!D�<u(�"��Z����-�~�L�OLt��`��7��������x��г��.���y��iǵ�9���N��Y���񿇿�e��A���'��n�q� ��4�qU���}�ړ�ť������X��#+���}���0��o������������٩�˄�� ���`���=�c&����H�$�\�:�o]��5��!����
��i���jg���������+���˶��V���C��o`���"���b��A�[���:���%�����I)�W�A��\e�⥇����0������i��T���㵿rK��N�������ﲿ�[蔿T��
X��8�N�%���"���.�:KI�/qn��O��K3���?��<i���O���跿����yb������X�����Ϥ��쑿�y�!ZR�B�4��7$�ER#�8�1��bN�F�t��Ӣ�VͰ��η�X츿RX���f��*q����������+5��ޡ��\���vr�SL���0���"��$�}�5�aFT�p�{�������'���h���Ӹ�v)�����׷�&������g��c��������k��NG���-�
l"�+�&�(`:�׮Z����O���m��"%����ø�w��ж��Q��nL��^2��v����1�����e�:�B�!+��m"��o)�0X?�,ea��Q��3�����  �  D���`h�d�࿲Lʿ=n���t��+>��h���:�u�Q�Y���<���!��6��$���B��'� �%���'��lC�d`��{�V���P��<��G0��ߝϿDc� ����ʑ�cf˿@#��]>��Y�b���E�ޔ@��AS��?|�`o��������ۿӈ�Z��H;���ٿ� ÿf=�����bE���σ�g2m���P�B�3��]�����������c����C�0�HM��i��H������2替#���R��B"׿};뿸���1���w޿�k���֞��π��rV��DA�0D��^�G7��3���Hȿ���	���g|��wI�p ӿ�b������!����ٌ��L��~e���H�[�,��!�خ�1	���| �tD��V"��=��Z��\v��0��W�������� ��!�ɿ�L����!������N׿�F��c9���Au�Q���C���N�;�p��������ÝԿ���ݛ���+��B}�^ͿX*��-�������s��ID{��l_���B�a�'�� �R���� ������W2.��J�)g��]��G���ʚ�t����ӿz���[��b���z7�/)Ͽ���M<��k�xEN��I���[��i��G���6E��������9������޿�9ǿCo��*ա��i��
�cu�\�X�
<��w"�
(�������u������8��dU��r�_���ْ����F(��Z~ĿRSۿVq￉��������x�Ŀk������^���I�hBL���f��!���|����˿�1��J��������@Xֿ^���]R����85�������l�{2O��,3��]���
�l���[�J�q�'�j�B��|_���{�mΊ��K���8�������I̿m��x���ʵ���e���ٿqɹ�Ю���z�r�U��lH��+S��u��L��.��H�ֿ���  �  H?,��&����E��.Aοr���r��;h��DF��A*��T�/���e޾8�˾K�ƾ�ϾCn侀���w��F0�!iM�21q�����jv��5ؿ͂�k��V�(���+��!��A�i�濇�������:t��Ml�� ��)�пC�l���)��+�C�!�������v��� ���MJ���\��<��X"����]򾀺׾=dɾ$�Ⱦ�gվ;��wG	�s}���9�i}X��M��m��? ���_翗>�ǡ��#+�f�)�`������eտ(���l��Rm�Qfq�av��E���BI�q�
�e[ �V�+�i*��&�>��m޿_b��Qᓿ�~w���R��45������	H�)�վ�D̾*cоu�Ᾰ?���>��*�4�F���g�'��%���j˿�������%��0-���'�E��J��m�ƿ�����f��lo�������������������v&���-��|'�e�C��$�п�9������G�m�`�K���/���*��N���׾L�Ҿy�۾JD��	��#��7��GT��x��s���ﲿz�ۿ�<�Z�]j*��-�=�#��(���h���>ޓ���|�^�t��M���@��oYԿ7�y��wC+�z�-��#�������Ŀ\"���n����d��E���*� ���H����։پc�ؾ��_���:_���'�ݲA�Y�`�-������&���뿀W�@�!�AA-��,��	����u�ٿDZ��������u�r�y�a��������%�a���&"���-���+�D���7��g�ѽ��->���4~�|Y���;�N�"�\?�����O��@ؾ�ܾ}U�;�ƻ��E0���K���l������G���ο�������&��.�,�(�j8�A���Geɿ���q�T�s�*́�w7��I$Ŀ ����&z'��  �  s�f�E
]�c*C�;  �����ƨ���*��n\���/�������nϾ����2���譥��쫾U(���T־�(�����=�8���h�u��<ȿ��](��J���`��Uf��X��t;����v�ʛ���4�����������˿g9�~+��:M���b���e��V��<8�����⿲���x��RL�t�$������p;Ǿ@����ꧾ�Q��dٰ�pKľ��Ὰ=�� ���F�O}�y�����ۿ���#B4��:S��d���c��8P�.t/��
���ѿ�����f���6����:}߿���K�7��NV��f���b�s�M�X�,�J[��LϿ����>4q�_?����
��G޾wKþ�K��dC���d������/�Ҿ���1���i/�L\Z��勿F����������@�g�[�[�g��`��gG�$�����¿�����̍�`瘿&ͼ��I��� ��D�Uu^�*h��k^�[�D�ۀ!��C���b��q㐿��a�2`5�����	���ھy]þ����b ������ɾTt�BC��J�%�?�`�o�������˿����*���K�.�b��h��Z��a=�+��g���Ѵ�{�������e��Bп�e���-�eO�ٷd�g�g��9X��\:�s$�*�=��?����T�X�,��6��7���o׾��¾���Tu������tԾ���5[���(��$O�Â�sͩ�i�߿���M[6�^VU�O�f���e��ZR��1�6B��5ֿ�ǧ�����i��n����㿹|���9�{X�R�g��}d�@fO��z.�H
�Z�ҿ�����w��E��K"������a�Ͼ ���:?������	Ǿ��ݾ����	�.�4���_����WW��u����N�T�A�']���h��ga���H�wW%�<� �#�Ŀh���� ��"5����ل��21!��'E��z_��  �  �S���&����p�P#C�����|տ��$_�(�3y�6�վ����!f������e��r����f���"���`߾!�
�n�2�� o�~���0	�!����M���y���������q��;�g�,m8�8�
�+GϿ맿�ʠ�Fҹ�~���@#�IIS�_~�ɶ��f���u����b�f3���?4������f�J�;��IT���$ʾ�L��]K��}\��ݑ��Ǚ�`���,ƾ�Y�L��*D���������A ��-�ӈ]��ׂ�a��Cy������eX�T(������V��y���QX��F1ɿA��3���b����b���Ì��s~��S�S{#��xￄƫ��y�G:�"2�\y�/�¾�;��6����򕾠��������4���ؾͺ���&��[�`��S�Ͽ*}���>��<m�S=�����������v�׌I�T��q�Oz������c��t޿�5�TD��lr����0���։��Rr�|�D���76ؿ����_�d���-��	���@���1������ع��/)��UG��FȾ��쾔[��9�C�u�42�����C����O�ܠ{��x������a��,�i��s:����ӿ=��a$��?/������n%��uU��D��ˍ�d������d��75����_ÿ������R�B�"�����eھ����>w��̂��w���쩾ZϺ��F־$����p�EXL�G����0�� U�}�/�!�_�����"�������+����Z�y*�������¿�����bͿ��5�x�d�ԅ�����֝������PU��'%����"��G��+�@�f��]x���Ͼ��������@�I���(��cþ}㾚	��&,���`�5���A2ҿV���@���n�N���c������8�w�x�J�~>���;ҵ������B�����hV��mE�*}s��x���  �  0����}���P��bs]�%�e�������e���&�|���ρȾ���q�������c����V���L���n��8�Ҿ���2�#x��󰿀7����1�;j�ax��BG��S;���@��ރ��	Q����|g�@���殿<̿i}��k8��#p����Gw��aʢ�EW�����J�*f�>5пA���1N�)��,��M���ן�s���0y�����KJ��E��jn��xU�p����F��G���ǿ����GD�)|��A�����EZ�����tv��X>���&�ѿ����<��;@޿U���J�G���w�������������p��D8�@�����3���"�:�����۾�+����-f���(������(������ʾѸ��%�� a������P㿊� �YX����Ya��]���}��+p��߽d��-�V���tĿ����vK������`�'���^�����2���1���-��� ����^���&��]��ե�+k��h,������Ӿ�����K��Ĝ��x���<�W/��!�����߾d��m�9�X�~�cl��� �<o3��k�[V�� (��O"��?1���ل��S�����������F����п��	���:��Pr��������^ݣ��h��x����L�A��`Կ�%���nV�@ �:����̾�����������	)��Uo��4n���Ⱦ��W"��N��c��)�˿��#^F�xB~��O��+���j��I/���4x��~@��F���տ7U�������z⿳g�y�L�z���c���ӣ�p������Dr�y�9��K�y�����j�A�Ϩ����r���Ď��]���G$���J���]��˵� �վ����]*�V<f��0��G��[�!��kY�V��	�������!����\�e��.�j� ���ƿ#Ɀ۝¿�!��%�(���_�#y��A����  �  �ր�B�v���X��9/��=�6���� ��Q�@�6M���־����ip��iz��"h�BAc�6#k�h���ד�4&�����>7�k�O��㑿-�Ϳ֑�k�8��`�/{�ޞ��}q��P��%�VJ��^m�������N��;v��O�ۿ�����=� cd���|��J��b�n��K��� �IF��8��zq���-��� �B�ƾ��������$]t��f�B�e�\�q��[���6���t��9��� �'�XQh�*���Ʀ����G�Lk��~��@~���g��MB��x�J��t���'���Y������>�$!���K�пn�1n���1}���d�.>�����Iֿ�x���eY��H�(��b�����׆���v��Qn�wr�#끾�v��ݐ����׾ c��=�1Ճ�W��� ��Q+�RU�qu��C��d�y���]�+$5�i�
�6=п!���J�������ʿ��V�0�@�Y�:�w�1����x� �Y�z�0���E�������cF�`��������������������{�a'��hB�����{��jN�R�{�V�bW���ѿ�J���:�lbb�5�|�����Xs���Q���'�fm��~����坿J���Bɭ�$��!�'�?���f����[��J�p���M�h�"��s��_��~�y��6�&	��׾�밾�����O���j�����:��z��b\����ѾA����/�v�p�[ʧ�k��/��a&I��em�À�/����i��nD�{��翘���#f��܏���8���P���#�\�M�ۑp�N����~�x|f�q�?�,a���ٿ�Λ�_`���$�������Ⱦ	ԧ�`U��շ������넾�V�����4������6��PC��o��������,���V�mv����W6{���^��^6����ҿ�l������G���`̿����1�T�Z���x��  �  ��v�u	l��^O�(�]������������>�C@��ؾ�ޭ�l葾.���ɦn���i���q�Dԃ��K���7��-�徬���L�5i��Yǿ1��Z1��W��?p��/v��2g�XG�!+��*�t��#c���b���q���5ԿUM���5��Z�Ur�"�u�.Zd�w'C��c�Q��C~��?m�q},��I�ǀɾ:�������{�m��Kl�ݣx��Љ������;ľ�����&�Md��G��׿ݿU����>��5a�~t�$Xs��^�0G:�9����ڿ;��0���:��_��I��]���BC�w�d�/�u��Or�>[��N6����AϿ�����*V�m��Z ����0����F��n�}�#�t���x�CK����԰�.3ھ�����;��%��:泿?���m$�7SL���j��pw�DFo�gKT�B�-����:\ɿ�l���k���x��S�ÿI��hj)�٦P��jm���w��hm�9�P��u)�� �Ot���ʆ��.D�Y��,��3���s���a���]���%���o�����Sf��.�þ�!�ן�M�S��ܑ��tʿ��	��3�I�X���q���w�Xi�HFI��+!�K��������.����è�ӈؿev��8�l�\� -t���w�zf�~DE��}���0����Iu�F�4�	u	�P�پ�F��d(��7���{����?��jl��*���skԾ(p�C�.�}l�(e��v��n����@�/Oc���v��uu� !`��g<�t��t߿5|���l���n��e���h����(E��kf�\�w�=t�й\�4�7�t����ҿ�	����\��D$��>��C�˾D���Ė�,��:U���*���������Ļ������/A�㿃� ������^�%��M���k�<�x���p���U�;
/�j����˿�ơ�X���ɞ�	�ſ��K�*�S�Q��rn��  �  UX��+O�P6�2�������`�y��#:�d��5������]��z��N����}�2��=ގ��ˢ����(P��ÈF���������.����� =���R��X��K�x�/�'.��Sؿ��q���	y��:����������-� ��[@��sT��mW��H�,�oW	�6�ϿBV��BYb�AA*�����RӾ+x��eP���)��e���m3�������������Zξ�? ��%���Z�����ȿ)Z�bA(��E���V�}�U�v,C�m$�����/ſ	ڙ��(���ˇ�7�����ѿ�a	�M1,���H���W�V�T�Ԛ@��$!�C>���ڼ��%���N��X��D��gSɾ���4e��72���`��0�������X������L㾴@��!8� u�Х��߿���!4�N��1Y��0R���:������Ό��h���������W����*�o!���7���P�M�Y���P�P�7�UT�1�翁X����|�?�H�L��qSľ�騾�B��j����#���ŏ�񵛾�䯾�[ξU������{kM�~��V0���B������>�=�T���Y�[�L�}�1�+��kܿ�A���䍿S��� 뚿=�ÿ ���"��B��V�+�Y��J�,.�Yq��Կ/}����j�	w2��� ��w����y���J��/����L�� ����0���3����޾6^�=)-���b�<%��>Ϳ3n� X*�J�G��X�حW�@KE�׌&�ɦ��oɿ��`�������إ�Q�տ&V�?.���J���Y�E]V�AFB���"�w����/��F|���tU���#��1�\E־&Ķ��⡾Im��TW��ZV��	���s����Ǿ�
�,���]=��Iz��i��!#�~L�KW5�NcO��Z��zS�4<�:��q�S︿�픿�����Z��[߳��f꿄8���8���Q��  �  ��.���'�n��m����ÿ>9���Lj��8��,�_���� оw�����������ɐ�]������l��~ؾˏ ��R���B���w�1a����ο���}%�c�*�d�.�ɔ$��D��-��(��#$��ҳq��i��������q�ѿر��9���+��C.���"�A1�Z�
�������{X��,�W(�=z�t�ƾw���K����˒��J��iC��J���{þs��;	�2�'�r�R�����Qͮ�8��I
��� �އ-�B�,��c�����$׿,O��+���'�j�n�n�$ȋ��2���e���~�"��.��;,�������iտ�勵d��'�I���!�M3�R/�����]��3���[��n��!���i��j4ӾA���M}���7�7�g��Ҕ�#���p�Hm��I'���/�EK*��5�I1���!ȿ)g���L��[=l�|�|�ƚ���¿:���E��3*)��C0�ZH)��t�I.���]ƿ�󙿩�o��8>�0��_� ��v۾*1������>���������rl���ƾhV�R�C)#���I���~�Qգ��Uҿ?i�����z,�Hr0��j&�T+���M5���G��Nz��r�hT��lF����տO���_��.��e0��%�6N�A�v7��p&��%�`�CP4�tS�7���f�־� ��⫾碾
d��_]�����E5Ӿ�����"���/�7�Z�����ﲿ-�b`���"��/��.�܁ �x���aۿ:����ǉ�w�r�-w�Xڏ��-���B�c~�=�$��H0�J�-���j��J�ؿ�E��	����0P�Dy(���� �j�;:ٶ�&m��_R��.�������{�¾Z(޾��;��!=���l��l��P�¿f�������(�(1���+��z�����ʿq̞������p�裀�	ޚ��#ſ������v/*��  �  �R�0 �e��-�ƿ�������De��B��6'��a�+�����ؾ���~Ȱ��f��Z���ľt�߾��U�-�W�I��Pn�Y���wج���ο�A�I����2���yۿ���/���Bl�:�K���E�:�Z��`���i���=˿���]��������|ݿƿ���������Y�;V9����
���оT����ծ��,������Ç;�����`���6�C�T��|��=���Ϸ�R�ٿ����������.ϿVK��pn��a^���F�F�I���g����������׿[b����V����a/ӿU���ْ��t�p%O�t�1���m9�ص�RL̾�㹾���Ty����þ�ܾxN������(���B���d�[������Ŀj"�=����K�����s�ĿL���5��L�W���H�OU�{�P�������{忖d �˰��c�%\꿵�ɿ�L������d�j��H�p�,�����x��x��˾hѼ�c���=忾C�Ѿ��쾜������3�,�P�;u�Tk��qK�� ҿ>��k��\��t0��==߿繿a��Vpt��3T��PN��Bc�M���������Ͽ��'��7�����7��S󿿴ן��C���]a���A�e�'��"����\�ྻ�ʾ�wE����Ⱦ�ݾ���I��P%��+>��]�V����_��������ݿV�� ���������gӿ����O���r�f��N�^�Q���o�́��⵿�ۿ;������s��s��)�ֿ�����0��Uo{��U�.n8��M �4��,k��K�ؾ�ƾ�����.���`Ͼ^P羝��B���b-��(H��i��������ÍǿN���F�ɛ�f�X ��ǿǿ�����ې\�%�M���Y�^���읿=�¿ڐ�fh��  �  �n��Ŭ��!���)��qF�������!u���`�9L��5�g��V+	���ﾨ�پ�5Ӿ/=ݾ�q�������#�4;�/Q�Ĩe�pz����lҖ�����h���h������9�'㡿7G����b��0=�'�&�)�"�s:1��P��|�[=��%����b��u¿"绿yP��B���տ��i����n��Z��rE�9�.�h���8�8n�=f־�tվ��#�*��+���B�?=X�H`l�p��������Y���v��@����=��2�Ù��ـ���T�ۮ3��d#��%��:�to^�oц�����K�������ν������~����e�������4~��i��cU���?�)�(�bb������n���ؾ��ݾ)k�'
�%����6�iM�rib�:�v��K�������?��*Z�����!�ÿʁ��$�����m�u�� L��r0��8&�c�.��H��Nq�,��O�����e+Ŀ~n��zյ�t饿����t��t�z��jf���Q�*m;��j$���9U��b�� {߾���w���O�J�*�$�A��X�m�l�f���!���F���w��cݹ�5�ÿ TĿ*����������N�j� DE�92/�D,+�è9��Y�Ø�������D��*����HƿD%��u���i2���쒿�:��Iw�"�b�T�M���6�M���L����Հ������s1	��;���3�b�J��b`�,�t��Ȅ��,���*��L��������ſes¿�$��\������&�\�M�;���+�&�-��B��.f�~���[`���5���@Ŀ�ſC�����̻���M���r��,Wp��\�/+F��/�c������Y��s~��������U
%�|"<�\�R��g���{��䈿(���ޥ�~���^S¿�Aƿ���᳭�J����z�W�P�]05���*��,3��+M�f�u��K���`��?����  �  �;������Ò�����0���Ԓ����������V��Ur�0%R�&y2�m\�*��Z����
����AP9�,�Y�a�x��ψ�O�����ђ�����P�����}���������Qm�~M�	�-��.��r�J��NE���!���>��J_���}������1��WA���˒��*�����lG��G+��V�������A?h���G�])��
��0�:|���qF&��D�@�d��������%��}��1���*������h��W��v4���b�B��$���������H�8J+��#J��j�QЃ�������E���:;���撿a�������ҷ���֊���}�%Q_��	?���"�������}	�K��\2���Q�$r��ۆ�����O��Zϔ�o��Bړ�ؚ�������Α������z���[�j�;��Z ����S�<���I�u�8���X��x�y���Z����i��D�������=���猕��V��K�������w�+�W�oF8�rE�����	�C���#���?�X*`�J���7��"���[|���G��$���Yŕ���������o���y1����t�*�T��5��)�F��p������b*��LG�8�g��)��mҎ�Br��P~�����D]�������m��XK���
��}���"`p�{�O��p1�~��=�����uT.�W!L���l��#��F��*ʕ��A��B���e�������A������M����g���j�\J�g�,���_<�Ҡ�����2��Q�r��U��`e��p\���O�������=��떿gP�����C%��g>���e��ZE���(��������[��� 8�kUW��w�����.����薿�g������Ax��;<��:]���o������
���`���@��3%����Z������"��M=�z,]���|������  �  ��a�S2v�_c��������糿L$���S���O������K��/�i��+B��")��!�!E-���I�Yat��񒿣p���_�������n���Ű�����v��U郿�r���]���H��T2�TM��>�*��4ؾ.cԾ�ᾏ���˞��(��0?��T�nCi���}����-����ܩ�미�S��Vֿ�>8�����/.��N�[��f8�v%���#�/[5��W��`��1H��� ��ݾ������广
���o!���A������k��V��NA��Z*�ܹ������=�_վW/׾xb�ŷ����0�Q�G�K]��Oq� j���>��g���+鯿8���¿��������m˖�E�{�ԊP��92��$�-B*��A�~h��#��_���Wn��c�¿�����a�� ا�赗�6���;k|��h�@�S���=�q�&�������V�便�۾&�㾻����%��%��C<�Q�R�mg�g�{�'$���֖��Ц�➶�(����Ŀ���~S��0'����o�lH��'/��(�o{3��IP�9�z�9���ǭ��ľ��Xſ�����<�� ���w��F`��ky�;e�%P�p�9�F�"�����T��� ����X����#��0���G��w]���q��3��A-���������ռ��rſ7�ÿ�L������:����c��u@�2-�t
,�g=�m-_�Gi��S���.�� �¿\�ſ)�������F��[k���*��'ss�?_�	�I���2���#7�0��<'徶 �����eI�\� �o�7���N���c��x�Ć�G���)���B��x���V)ƿ�����������l"����V��L8�_�*��#0��VG� �m�Fꎿ�m��&���Yſ�aĿ����_q���R���U��~׀�Y\m���X�5�B�2�+�Λ�?V�&QA�,�쾕��3t�26)�"]@��V��  �  �"D�v)g�a��#O����ȿH鿎� �Q�����ῄ6���n��o�s��)O�z�D��%U�;2� >����Ŀov�E� �zZ����}���L������'����_���=��~#��?��Y��u�Ծnx��믾#j��E4���uɾ��^~��N�ް1��xO���u�ᨓ��n��GSԿ���������m�����տ�ï�?����4e��I�ƎG��`��F������Olѿ@q�>���m������׿.�������.z���R�|L4��u�mW���辍�˾Yŷ�9	�������U��Ӿ�2�r��"�� <��p\�|��	��g[��J�*���v������ʿ]i��{ヿ�3[���G���O�:hq��;��������޿9k���eS��k�pοˬ��9����o��K��@/����������˾�8��T2�������ʾsM�������g�-��I�Ȫl�H!��H���q˿[��������6����������[����y�@0U���J��T[�5����n��ȿ��/[�O�8B �5!���ĿJ��tv��� f���D�ժ*��������+�9!;e㿾6����ƾ�ھ�g������!�',:�C�W�"~�ߗ�����~ؿ7����a��������ٿг��Ő��Cm�1Q��O���h��M�������vտ ����x�������ۿ���Qƚ��B��2[��<���#�_��a?���@ܾ��Ǿ�����F����˾u�ok �6,�O)��B�'3c��x��z`��β��3Y㿶���3F����,�FͿ#��������Aa�8�M��eU��6w����a��;�ῐ��<a�����ѿ8g��sّ��t���P�Pw4�N����O���վ��ľy����þ�{Ӿ�쾻�����1��  �  �:��wm��e��2[ƿ c��S]�x�(�Y�.�'��I���ܽ�Gd���Ov��h�Z�~��\����ȿ7=��N���*���.�ې%��9���!��� ���8a�U2�����ik˾Xj��y���œ��´���U���D��S{����޾���]$"���J�Eu������5�׿��j��h,�j�-�1�!�Z��A࿒����=���m�l�k�1���٩�LHڿ����78-�98-����x���!ݿ$K������ƞO���%�(a�SH�-��?6��F���:T�������Q���T��D�ɾ�����)m/�ɻ\�Ʋ���U��,��<��6$�c�.���+�H�����Ͽ�᡿Egik�ɸu�X0��������h�F&���/���*�X��3���Ϳ ՟�zx��C�.������ݾ.��ު����񙙾V������ƾ�ܾ���	"��s@���r�h%��ɿ���R���*�PG0�Ww(�9��L��������_���W|��n��S���y��̿Ժ ��)�]�+�0��H'����b6��3��w��{1h�Ia9����أ��]Qھ����Kn��8p���ס�����Iַ��3Ͼ�zﾓX��*��S�?���Eͫ���ۿ	1�ʽ�bw.��0�'�#�(��M�󺲿;E��D�u�{�s��6��T୿UP޿+!
�P�!��@/�C/��!� �
�vE��r��F&��u�W�R�-��������Ѿ�������"-���$��{���a<��HPؾu������D6��|c�n��C���"�����%��0�Nb-����C�[�ҿ錄G��aq�~�{�s��0����o������'�k�0��D,���Le��pпt���P}���H�'d#��#����1�ɾ⛴����ߢ������岾VǾ�e侶���$ ��  �  �<���}���� {����08�(P�HWX�fVN�V�4�����T��ڬ�O���e����ё�O��Ǔ�K��ٛ;�0 R��&X�#L�(f1�v(�>ڿ�N����m��2�	� oھ-F���p��L���7@���h�V>���/�������Ǿ}����u�P�$ǌ�EN���R��8�"���A��T��!W��kG�f6*�e�O�οFʟ�3���兿�囿�lȿ��Pm&���D��-V�V���D��h&��l�k�ſ�y��W��h"����O�˾�F������Me���Y��'q������k���~����׾���.�"rg���sԿC���A.�0J��'X��/T�gM?�qI�� ��}ٽ�G)��`Y���ۋ�9����ݿ
���42��M�@	Y�U�R��h<�H�����n���*����F�U��F�� �ƾ�e���A���O���������Q����k����ľ ����oB�����C��8뿀G�1�9�j�Q���Y���O�MM6�si�2I��د�6��������ᔿ�-��$��j��<=���S�o�Y���M�<3������ݿ�Ĥ�}�t��9�;A���辠þ���p������Ï�΋��-���LN��+�ؾ3��n~&��Y����тÿ>��^�$���C�9W��-Y�SuI�>,� k	���ҿ�ѣ�9��뉿�럿Gs̿֌�^r(��F�96X��X���F��w(�M~�`�ɿJ����n_��*�����Hܾ9����0���i������쐾�ݘ�By���3�����ۭ���4��1n�����h׿*T���/���K���Y�?�U���@�� �B3�������*��U���ю�Ԉ����߿�@���3��eN��ZZ�],T�4�=�{�Mm����<ˇ�!7L�2���(��#�о�Z�������є��쐾���N��������H;'�������  �  ��A��~���%��߂��d*��VQ�P,m�ؖv��j��iM�.�%�B����d���ۘ�wY���䞿}Uʿ���/�t8U��Wo��_v��sh��gI�r@!��'�}宿^;z��_5�S%��"Ѿ~���t
���g~�^5n�V`k�P�u����y%��5a���0𾠣�|X�}����Iҿ?��08��l\���r��%u���b���@��h�Y�忘��^���/�����L�޿��ؗ<�?�_�+t��s���_�"�<�n�.�ٿJ��?`�B�#�h���W����֞��ǈ�w�w�Z�l���n�<#~��T���]��Uξ)]���0���r�O������@�E��/f�Rv�-�q�rnY�44�ڬ�Wҿi���D6��,����X��Zf���$"��)J��Qi�~=w�*p��V���/�$���$ſ����7�L���@��fѻ��松�A��t ��_V{�׀��Ԋ����	湾�@澦���qG�3?���徿�����+��R���n���w�AZl��N�Yb'�b����d��᛿�b����iͿ!T�~�0�k�V���p�ox�W'j�BK���"����[�����oi<��H���߾ͷ��)��@���;׆�����Z������Ƭ�"ξ4� �!'���`������}ֿ��E:��~^���t��1w���d��C�tn�����&��P�������������a��Ԝ>���a�qv��	v�w�a�b�>�����ݿ�r��Kdh���+����XҾ�2�������䋾���҆��0��. ��>յ��-ܾHN��7�|y���������!RG���g��w�&Fs��[�*�5��3�hտƻ���1��g���J���M��K�#���K��j�ɏx�uwq��dW�>1�+(���ǿ/,��� R�~9�_0����žܧ�����>���E�ډ�
���:~���:¾�g���  �  9SD�����m(¿���I�1�ۢZ���w�Jր��pu�jV�H�,�T��Ŀ,G��J:��蠣�-`ѿ����6���^��z�Q���f�r�sKR��(��5��^'���\��!7�����ξ���������w���g���d���n����������q��k�b�'�[�J���B�ٿ���-@�fEf���}�:����l�[I�W��d_�峴�ɟ���	��Hﯿu�濬���D�<�i���~���~��i���D��o�]}�(�����c���$��h��ŷ���r���W���:q��Pf��Vh�Zvw�����
���p˾t��*2��hw��6��#N�R�#��WN�|~p�
���2v|��c���;�];�blٿ"������	���t��E�����(���R�߬s�K'����z�!�_� t7��l�˿S␿\�O�X��羟���/q��_ׇ�5s{���t��'{��n��(}������q#侘����I�}P����Ŀ���*3�Q�[�k2y�Յ��i�v���W�\.�+����ǿ�L��rC������VrԿT���8��9`�i�{����[�t�~T���)�m��������)��+>����5ݾ���W����@��Y���y��O���K��;V���/˾?���O�'�Xd�O��� �ݿ����BB�TWh����F���o��bK�=� ��h��������0��������꿊����F���k���������ۺk���F�����念���&4l���,�J��82Ͼ9˫�フ������܂�y���H֊������~��G�پ��
�B�8��&~�b��������<%���O��#r�����7~�u�d��o=�p��0pܿǦ������ ���fÿzQ�@M*�#YT��u��Ё��:|� �`���8�7i��,οĂ����T����C���¾�f��L���Q;��˸�����o3��������IJ�x���  �  ��A��~���%��߂��d*��VQ�P,m�ؖv��j��iM�.�%�B����d���ۘ�wY���䞿}Uʿ���/�t8U��Wo��_v��sh��gI�r@!��'�}宿^;z��_5�S%��"Ѿ~���t
���g~�^5n�V`k�P�u����y%��5a���0𾠣�|X�}����Iҿ?��08��l\���r��%u���b���@��h�Y�忘��^���/�����L�޿��ؗ<�?�_�+t��s���_�"�<�n�.�ٿJ��?`�B�#�h���W����֞��ǈ�v�w�Z�l���n�;#~��T���]��Tξ(]���0���r�~O������@�E��/f�Rv�,�q�rnY�44�ڬ�Wҿi���D6��,����X��Zf���$"��)J��Qi�~=w�*p��V���/�%���$ſ����8�L���B��gѻ��松�A��t ��_V{�׀��Ԋ����湾�@澥���qG�2?���徿�����+��R���n���w�@Zl��N�Yb'�b����d��᛿�b����iͿ!T�~�0�l�V���p�px�W'j�BK���"����[�����pi<��H���߾ͷ��)��A���;׆�����Z������Ƭ�"ξ4� �!'���`������}ֿ��E:��~^���t��1w���d��C�tn�����&��P�������������a��Ԝ>���a�qv��	v�w�a�b�>�����ݿ�r��Kdh���+����XҾ�2�������䋾���҆��0��. ��>յ��-ܾHN��7�|y���������!RG���g��w�&Fs��[�*�5��3�hտƻ���1��g���J���M��K�#���K��j�ɏx�uwq��dW�>1�+(���ǿ/,��� R�~9�_0����žܧ�����>���E�ډ�
���:~���:¾�g���  �  �<���}���� {����08�(P�HWX�fVN�V�4�����T��ڬ�O���e����ё�O��Ǔ�K��ٛ;�0 R��&X�#L�(f1�v(�>ڿ�N����m��2�	� oھ-F���p��L���7@���h�V>���/�������Ǿ}����u�P�$ǌ�EN���R��8�"���A��T��!W��kG�f6*�e�O�οFʟ�3���兿�囿�lȿ��Pm&���D��-V�V���D��h&��l�k�ſ�y��W��h"����O�˾�F������Me���Y��%q������i���|����׾���.� rg�쮜�rԿC���A.� 0J��'X��/T�gM?�qI�� ��|ٽ�G)��`Y���ۋ�9����ݿ
���42��M�A	Y�U�R��h<�I�����n���*����F�V��H��"�ƾ�e���A���O���������P����k����ľ����oB�����C��8�G�0�9�j�Q���Y���O�LM6�si�1I��د�6��������ᔿ�-��$��j��<=���S�o�Y���M�<3������ݿ�Ĥ��t��9�=A���辣þ���p������Ï�ϋ��.���MN��,�ؾ3��n~&��Y����тÿ>��^�$���C�9W��-Y�SuI�>,� k	���ҿ�ѣ�9��뉿�럿Gs̿֌�^r(��F�96X��X���F��w(�M~�`�ɿJ����n_��*�����Hܾ9����0���i������쐾�ݘ�By���3�����ۭ���4��1n�����h׿*T���/���K���Y�?�U���@�� �B3�������*��U���ю�Ԉ����߿�@���3��eN��ZZ�],T�4�=�{�Mm����<ˇ�!7L�2���(��#�о�Z�������є��쐾���N��������H;'�������  �  �:��wm��e��2[ƿ c��S]�x�(�Y�.�'��I���ܽ�Gd���Ov��h�Z�~��\����ȿ7=��N���*���.�ې%��9���!��� ���8a�U2�����ik˾Xj��y���œ��´���U���D��S{����޾���]$"���J�Eu������5�׿��j��h,�j�-�1�!�Z��A࿒����=���m�l�k�1���٩�LHڿ����78-�98-����x���!ݿ$K������ƞO���%�(a�SH�-��?6��F���9T�������Q���T��A�ɾ�����&m/�ƻ\�Ų���U��+��;��6$�b�.���+�G����߽Ͽ�᡿Dgik�ɸu�X0��������h�F&���/���*�Y��4���Ϳ՟�}x��C�.������ݾ1��ު����񙙾V���~���ƾ�ܾ���"��s@���r�g%��ɿ���Q���*�OG0�Vw(�8��K��������_���W|��n��S���y��̿Ժ ��)�]�+�0��H'����d6��3��	w��~1h�Ka9����ۣ��`Qھ����Mn��:p���ס�����Jַ��3Ͼ�zﾓX��*��S�?���Eͫ���ۿ	1�ʽ�bw.��0�'�#�(��M�󺲿;E��D�u�{�s��6��T୿UP޿+!
�P�!��@/�C/��!� �
�vE��r��F&��u�W�R�-��������Ѿ�������"-���$��{���a<��HPؾu������D6��|c�n��C���"�����%��0�Nb-����C�[�ҿ錄G��aq�~�{�s��0����o������'�k�0��D,���Le��pпt���P}���H�'d#��#����1�ɾ⛴����ߢ������岾VǾ�e侶���$ ��  �  �"D�v)g�a��#O����ȿH鿎� �Q�����ῄ6���n��o�s��)O�z�D��%U�;2� >����Ŀov�E� �zZ����}���L������'����_���=��~#��?��Y��u�Ծnx��믾#j��E4���uɾ��^~��N�ް1��xO���u�ᨓ��n��GSԿ���������m�����տ�ï�?����4e��I�ƎG��`��F������Olѿ@q�>���m������׿.�������.z���R�|L4��u�mW���辌�˾Xŷ�7	�������U�� Ӿ}2�p��"�� <��p\�z��	��e[��H�(���u������ʿ\i��{ヿ�3[���G���O�;hq��;��������޿:k���fS��k�pο!ˬ��9����o��K��@/����������˾�8��T2�������ʾpM�������e�-��I�Īl�F!��F���q˿Y��������5����������[����y�?0U���J��T[�5����n��ȿ��0[�P�9B �7!���ĿL��vv��� f���D�ت*��������+�<!;g㿾7����ƾ�ھ h������!�',:�C�W�"~�ߗ�����~ؿ7����a��������ٿг��Ő��Cm�1Q��O���h��M�������vտ ����x�������ۿ���Qƚ��B��2[��<���#�_��a?���@ܾ��Ǿ�����F����˾u�ok �6,�O)��B�'3c��x��z`��β��3Y㿶���3F����,�FͿ#��������Aa�8�M��eU��6w����a��;�ῐ��<a�����ѿ8g��sّ��t���P�Pw4�N����O���վ��ľy����þ�{Ӿ�쾻�����1��  �  ��a�S2v�_c��������糿L$���S���O������K��/�i��+B��")��!�!E-���I�Yat��񒿣p���_�������n���Ű�����v��U郿�r���]���H��T2�TM��>�*��4ؾ.cԾ�ᾏ���˞��(��0?��T�nCi���}����-����ܩ�미�S��Vֿ�>8�����/.��N�[��f8�v%���#�/[5��W��`��1H��� ��ݾ������广
���p!���A������k��V��NA��Z*�ܹ������=�^վU/׾vb�ķ����0�N�G�H]��Oq�j���>��e���(鯿8���¿��������k˖�C�{�ӊP��92��$�-B*��A�h��#��`���Yn��e�¿�����a��#ا�굗�8���?k|��h�C�S���=�s�&�������W�便�۾%�㾹����%��%��C<�N�R�mg�c�{�%$���֖��Ц�����&����Ŀ���}S��/'����o�kH��'/��(�p{3��IP�;�z�9���ǭ��ľ��Xſ�����<��"���w��H`��oy�>e��%P�s�9�H�"�����T��� ����Y����#��0���G��w]���q��3��A-���������ռ��rſ7�ÿ�L������:����c��u@�2-�t
,�g=�m-_�Gi��S���.�� �¿\�ſ)�������F��[k���*��'ss�?_�	�I���2���#7�0��<'徶 �����eI�\� �o�7���N���c��x�Ć�G���)���B��x���V)ƿ�����������l"����V��L8�_�*��#0��VG� �m�Fꎿ�m��&���Yſ�aĿ����_q���R���U��~׀�Y\m���X�5�B�2�+�Λ�?V�&QA�,�쾕��3t�26)�"]@��V��  �  �;������Ò�����0���Ԓ����������V��Ur�0%R�&y2�m\�*��Z����
����AP9�,�Y�a�x��ψ�O�����ђ�����P�����}���������Qm�~M�	�-��.��r�J��NE���!���>��J_���}������1��WA���˒��*�����lG��G+��V�������A?h���G�])��
��0�;|���qF&��D�@�d��������%��}��1���*������h��W��v4���b�B��$���������H�7J+��#J��j�PЃ�������C���8;���撿_�������з���֊���}�#Q_��	?���"�������}	�L��\2���Q�$r��ۆ�����O��\ϔ�q��Dړ�ښ�������Α������z���[�k�;��Z ����S�;���I�t�8���X��x�x���X����i��B�������;���䌕��V��I�������w�)�W�nF8�qE�����	�C���#���?�Z*`�M���7��$���^|���G��'���[ŕ���������q���{1����t�-�T��5��)�G��q������b*��LG�8�g��)��mҎ�Br��P~�����D]�������m��XK���
��}���"`p�{�O��p1�~��=�����uT.�W!L���l��#��F��*ʕ��A��B���e�������A������M����g���j�\J�g�,���_<�Ҡ�����2��Q�r��U��`e��p\���O�������=��떿gP�����C%��g>���e��ZE���(��������[��� 8�kUW��w�����.����薿�g������Ax��;<��:]���o������
���`���@��3%����Z������"��M=�z,]���|������  �  �n��Ŭ��!���)��qF�������!u���`�9L��5�g��V+	���ﾨ�پ�5Ӿ/=ݾ�q�������#�4;�/Q�Ĩe�pz����lҖ�����h���h������9�'㡿7G����b��0=�'�&�)�"�s:1��P��|�[=��%����b��u¿"绿yP��B���տ��i����n��Z��rE�9�.�h���8�8n�=f־�tվ��#�*��+���B�?=X�H`l�p��������Y���v��@����=��2�Ù��ـ���T�ڮ3��d#��%��:�so^�nц�����I�������̽������|����e�������4~��i��cU���?�'�(�ab������n���ؾ��ݾ+k�'
�'����6�iM�uib�>�v��K�������?��-Z�����#�ÿ́��	$�����o�u�� L��r0��8&�c�.��H��Nq�
,��O�����d+Ŀ|n��xյ�q饿����t��p�z��jf��Q�'m;��j$���7U��a�� {߾���x���O�L�*�&�A��X�q�l�h���!���F���w��fݹ�7�ÿ"TĿ,����������P�j�"DE�:2/�E,+�è9��Y�Ø�������D��*����HƿD%��u���i2���쒿�:��Iw�"�b�T�M���6�M���L����Հ������s1	��;���3�b�J��b`�,�t��Ȅ��,���*��L��������ſes¿�$��\������&�\�M�;���+�&�-��B��.f�~���[`���5���@Ŀ�ſC�����̻���M���r��,Wp��\�/+F��/�c������Y��s~��������U
%�|"<�\�R��g���{��䈿(���ޥ�~���^S¿�Aƿ���᳭�J����z�W�P�]05���*��,3��+M�f�u��K���`��?����  �  �R�0 �e��-�ƿ�������De��B��6'��a�+�����ؾ���~Ȱ��f��Z���ľt�߾��U�-�W�I��Pn�Y���wج���ο�A�I����2���yۿ���/���Bl�:�K���E�:�Z��`���i���=˿���]��������|ݿƿ���������Y�;V9����
���оT����ծ��,������Ç;�����`���6�C�T��|��=���Ϸ�R�ٿ����������.ϿVK��pn��a^���F�E�I���g����������׿Zb����U����_/ӿU���ْ�߿t�m%O�r�1���k9�յ�PL̾�㹾���Ty����þ�ܾ{N������(���B���d�]������Ŀl"�?����K�����t�ĿL���5��M�W���H�NU�{�P�������{忕d �ʰ��c�#\꿳�ɿ�L������a�j��H�m�,�����x��x��˾gѼ�c���>忾E�Ѿ��쾞������3�/�P�;u�Vk��sK��ҿ@��l��\��u0��?=߿�繿b��Wpt��3T��PN��Bc�M���������Ͽ��'��7�����7��S󿿴ן��C���]a���A�e�'��"����\�ྺ�ʾ�wE����Ⱦ�ݾ���I��P%��+>��]�V����_��������ݿV�� ���������gӿ����O���r�f��N�^�Q���o�́��⵿�ۿ;������s��s��)�ֿ�����0��Uo{��U�.n8��M �4��,k��K�ؾ�ƾ�����.���`Ͼ^P羝��B���b-��(H��i��������ÍǿN���F�ɛ�f�X ��ǿǿ�����ې\�%�M���Y�^���읿=�¿ڐ�fh��  �  ��.���'�n��m����ÿ>9���Lj��8��,�_���� оw�����������ɐ�]������l��~ؾˏ ��R���B���w�1a����ο���}%�c�*�d�.�ɔ$��D��-��(��#$��ҳq��i��������q�ѿر��9���+��C.���"�A1�Z�
�������{X��,�W(�=z�t�ƾw���K����˒��J��iC��K���{þs��;	�2�'�r�R�����Qͮ�8��I
��� �އ-�B�,��c�����$׿,O��+���&�j�m�n�#ȋ��2���e���~�"��.��;,�������iտ�勵d��%�I���!�K3�P/�����]��3���[��o��#���i��l4ӾD���O}���7�:�g��Ҕ�#���p�Im��I'���/�EK*��5�J1���!ȿ)g���L��\=l�{�|�ƚ���¿9���D��2*)��C0�YH)��t�G.���]ƿ�󙿦�o��8>�.��]� ��v۾(1������=���������tl���ƾkV�R�E)#���I���~�Sգ��Uҿ@i�����z,�Hr0��j&�T+���N5���G��Oz��r�hT��mF����տO���_��.��e0��%�6N�A�v7��p&��%�`�CP4�tS�6���f�־� ��⫾碾
d��_]�����E5Ӿ�����"���/�7�Z�����ﲿ-�b`���"��/��.�܁ �x���aۿ:����ǉ�w�r�-w�Xڏ��-���B�c~�=�$��H0�J�-���j��J�ؿ�E��	����0P�Dy(���� �j�;:ٶ�&m��_R��.�������{�¾Z(޾��;��!=���l��l��P�¿f�������(�(1���+��z�����ʿq̞������p�裀�	ޚ��#ſ������v/*��  �  UX��+O�P6�2�������`�y��#:�d��5������]��z��N����}�2��=ގ��ˢ����(P��ÈF���������.����� =���R��X��K�x�/�'.��Sؿ��q���	y��:����������-� ��[@��sT��mW��H�,�oW	�6�ϿBV��BYb�AA*�����RӾ+x��eP���)��e���m3�������������Zξ�? ��%���Z�����ȿ)Z�bA(��E���V�}�U�v,C�m$�����/ſ	ڙ��(���ˇ�6�����ѿ�a	�L1,���H���W�U�T�Ӛ@��$!�B>���ڼ��%���N��X��D��eSɾ���3e��72���`��0�������X����� M㾵@��!8�"u�Х�!�߿���!4�	N��1Y��0R���:������ό��h���������W����*�n!���7���P�M�Y���P�O�7�UT�0�翀X����z�?�F�I��oSľ�騾�B��i����#���ŏ�򵛾�䯾�[ξW������|kM���W0���B������>�=�T���Y�\�L�}�1�+��kܿ�A���䍿T��� 뚿=�ÿ ���"��B��V�+�Y��J�,.�Yq��Կ/}����j�	w2��� ��w����y���J��/����L�� ����0���3����޾6^�=)-���b�<%��>Ϳ3n� X*�J�G��X�حW�@KE�׌&�ɦ��oɿ��`�������إ�Q�տ&V�?.���J���Y�E]V�AFB���"�w����/��F|���tU���#��1�\E־&Ķ��⡾Im��TW��ZV��	���s����Ǿ�
�,���]=��Iz��i��!#�~L�KW5�NcO��Z��zS�4<�:��q�S︿�픿�����Z��[߳��f꿄8���8���Q��  �  ��v�u	l��^O�(�]������������>�C@��ؾ�ޭ�l葾.���ɦn���i���q�Dԃ��K���7��-�徬���L�5i��Yǿ1��Z1��W��?p��/v��2g�XG�!+��*�t��#c���b���q���5ԿUM���5��Z�Ur�"�u�.Zd�w'C��c�Q��C~��?m�q},��I�ǀɾ:�������{�m��Kl�ݣx��Љ������;ľ�����&�Md��G��׿ݿU����>��5a�~t�$Xs��^�/G:�9����ڿ;��0���:��_��I��]���BC�w�d�/�u��Or�>[��N6����AϿ�����*V�l��X ����/����F��n�}�#�t���x�CK����԰�/3ھ�����;��%��;泿?���m$�7SL���j��pw�DFo�gKT�B�-����:\ɿ�l���k���x��S�ÿH��hj)�٦P��jm���w��hm�9�P��u)�� �Ot���ʆ��.D�X��+��3���s���a���]���%���o�����Sf��/�þ�!�؟�N�S��ܑ��tʿ��	��3�J�X���q���w�Xi�IFI��+!�K��������.����è�Ԉؿev��8�l�\� -t���w�zf�~DE��}���0����Iu�F�4�	u	�P�پ�F��d(��7���z����?��jl��*���skԾ(p�C�.�}l�(e��v��n����@�/Oc���v��uu� !`��g<�t��t߿5|���l���n��e���h����(E��kf�\�w�=t�й\�4�7�t����ҿ�	����\��D$��>��C�˾D���Ė�,��:U���*���������Ļ������/A�㿃� ������^�%��M���k�<�x���p���U�;
/�j����˿�ơ�X���ɞ�	�ſ��K�*�S�Q��rn��  �  �3�wp,��4��R��fS��.Ɏ�7�P��@�1J�P��5\��K�o�.�S��E��A��G�5Y�ix�S'���G��l��18$��1`������̿�,�k���t/���3��)�
���7�÷���.bo�L�f��S��Ȱ��wԿ�s��7 ���0��63��'�(��+D�v���9��?�<��C�E�Ҿyؤ�إ����f��PO��D��|C��\M�.�b�3Ճ������.̾͜��
6��x��,����߿���
�$�cs2���1���"��t	�}Wڿ?�������h��_l��q������h#�@���C'���3�g1�>� ������ӿS,����i��+�Q	 ��ľ�ݜ��*ge��S�L�c�O�G�]���x�����n�������iM��ڋ��?�������Z��+���4���.�]����yʿq�����~�O�i�Y�z�/���ſ�%��7z���-��A5���-�������ÿ�����CV�ú��S�~9��屙��]��yik�y]���Y�ޙ`�}�r��B���m��{�Ⱦ���+��g��w��2пn���b��11�Im5���*����#&�Vλ����]�w�So��������,�ؿ��Y"�u�2��T5��()����mq��!���"����D��p�$��X���̖��_��txo��;d��c�.wm�a����쓾ٲ��.\ܾ���1>�B���?J����;����&�W�4�L�3���$�f���޿'u���,��\p�ܢt�x���������a��W)�B=5�h�2��B"�{n��4׿r|��M�p��]2�����Ѿ���������N~��zk���c���f���t��{��1����,���1�B$�~�R��t�� ۾�?h������-��6�G0��7��L��̿_��}����-n��?����N=ǿ�S�������.��  �  �f,�GK%������I蹿>튿[�L����0j��Ⲿ����Du�CaY�)VJ��KF��L���^�$�}�£���Ҽ����CI"� �[�����ƴſBE��vC�+(�H+,�D"�P��Xm俛����Њ��Ai��a���}�(�����̿,B�߹��`)�Ŀ+��- ���	���ݿ1{����{� �9�Ee
��]Ӿ)��n\��%l���T��bI�ݾH�q�R�-�h�В���Ԣ��4;���R3�is�����ȝ׿h�}�j+��<*���a��~ҿ㢿�M��8b��cf��z��̶��W�޿�)
��n ��,�0�)���0��ԁ̿�����d�7�)�VY����ž�H��`�����j�sX�<]Q�N�T��Qc��C~������a�����9����I�=���$��ӷ�^�.�$�YM-���'�����^��J�ÿ���rx�X�c��/t�o;��(X�����@b���&���-��&�ks�Ȩ��������LR��A�es�����J���,��Z�p��ab�v�^�%�e�sGx�G���餾RHʾ�� ��!)��ab����H"ɿJ������x�)���-���#�7���Y�H���w��q���i�����Ң�I0ѿ:d�����+���-��I"�D�⿔���������A����T���7��+���N.��!�t��i���h���r��]��
���b����aݾ[
��y;��={����ۿ		�d! �L-�'V,�� ��6�h�ֿP����o�j�]�n�Q���鯰�������:"�;�-�`+����9���ϿU؝�o�k��.0�wB��Ҿ�+��ih��񁾅�p�$=i�=l��#z�qK���������S��m���N��֊�)����U����%�>�.��)�b��������ſ�j���|��h���x�r���	�������4q�=�'��  �  ���������ֿ騿e怿C����6��6��ߙ��փ���j�Y�Z�"�V���]�up�D:���P���%þ���j�6�O�7=��%���oE����s�0���A�e����̿�꠿��~�O*X��Q�8�i�ww��>]���O�k���C��a��m���{ǿh����{k���2�R	� �׾0�����_Z~�x�e���Y��Y��c�s�z��M����(Ҿ[$�U�,�<d�_H���&¿7W� ������;�*�	��*�` ���/��]<n��R��U�(y�����ǿ������k�����u�J<�gܸ�}_���X�j�$�������˾�Χ����|��Qi�(�a�vge�۾t��M��۰��:��� 1�K��@���}�� ���zӿ�C �������G����ݿ'������h�e�a�S��=b�)Շ��'��8ٿ����Y�\m��X����RٿY���8����H��R��� ž�5���`��G=��W�r��o��v�g���E��>�����о<T�E�$���V�l���c��۲�T���0���������zlп;��z���}`��xY��Vr�i��������P=
�Ң�H��C��ܟ���˿�%��Ⱦs���:��K����!��-����H�������y��/y������l��ٟ�����U�yB� 5��6l��e���HƿB~�����n���T�Y��_�&U��b��>�v�ZQZ���]�����ǧ��{˿�V��ʮ����~�X 
�	�꿿+�� ���p�^��L+�a���ؾn���e���d劾�ۀ�p�y���|��Ʌ��x������%Ǿ���`���F��y��뛨��ֿ���6��!I������\�5��cz��%Yj��X���f���`���Eۿ���[`��  �  ��G�￹׿��������`i���8�Nr�����ʾ�,��5���=���w�x���s���{�_Έ��3���|����Ҿ����%��%�B�N.v�в������J�ݿ���e����O뿥Ͽ-���T����H^��k?�w�9�Z�M��ay�����Ŀ��@࿍��3R���`��̿�3��X����gX��$,�4����m���ʤ��p�������w��Kv�+����u������ֳ���'ྼ����'�X�R� ���$��%�ȿ��濟O��? ��}�&ÿP����5�?Q�i|:�!w=��Y�=e������˿
V�6����������"M¿�\���i~�e�I���!�����۾B߹�b
���4��H�Э~�7����k���ޙ�� ����;����.��P"8�,g�SV��&���ږտ&�����_���ۿ����R��J�q�k K���<�YH���l�h�0����ؿ�6�{���ݞ�F�ٿ`���Ε� �n�.q>����+�����վ������^w���f��k��G}��B����;��뽿�KMྃ��T�"�R�I��}�r!������I῜&��8N��1����ҿ���<����if���G��B�`V��퀿�C��	Ŀ\��8J��č��\��ѿa���Ì���`�\4��7��Z��%�о(�!����ǒ������1��Ӎ������n����̾�T����/�O�Z�m���F���Ϳ��&~��uQ��?E��ǿ�䣿)Ƀ�iY�-�B�țE��a��N��Ы��nϿ����G���G���忒�ſ
���E���mP�&(�):
�m辇�ƾ�������P$��DG��:3��%ؕ����x���Qlؾq�������W=��_l���[A��j7ؿ�]�e���I��R޿y���Ř�Awv���O�{A�s�L�q�2'��&-��+�ڿ�A���  �  ���}F��V��=����k~�!�V��6�:��=�Z��:_̾Ҳ�}Y��LW���揾�`��;���=���Ӿ�����J�!��<��"_��<���䚿�ů�h���_x��A����d��n#���a��:�O%#���W�-�hN�T�{����,���袽�����8=��ʤ�ZZ����p�F|K�Y-��R�y��o;�@4ľ�|��!L��G���%y��Wƙ����1��U�ݾz�������-*�уG��$l�騋�=7��w[����/e��d������Ox��UR�(S0��y���!���6�:v\�t����,���M�����Pm��퓲�]<��0���&e��'B��H&���̔����ھQv��r
��0��������E��𰣾̶��K�ϾUH��=a�#�6�neV��~}��
���
��l廿��¿���ū������yt�mI��,��8"�<�*�,�E���o�u/���⩿�5���tÿ������{g��n򁿿\���;�β!����� ���׾�]������Y���(���⡾�����>ž,Hྍ ���y�(�%�C�f������S���7��;��uĿH,�����K���~�h��*B��V+��*'�G"6�Y�V����"����岿U�����Ŀ t������1����Fy���S��5��~�Ϋ	�o��YԾ^���_����ń���ҩ�M(��8/Ѿã�+u����S2�I�O��]t�`ʏ�G]�������Ŀ¿�ʹ��L��������Z��8�}�'��)�d�>��3d�@[���ӣ�ظ�DĿ��¿�鵿Ѝ��G㊿d�k���H���,�V������p�V̾�x��oҧ�#q������!������ �ھ6��Z��"�k�;�[�{Z��⨗�D���D����Uſ����LS������ey��AN���1��&�zw/��UJ�v-t��R�����r>���  �  �V��ꏿ�����{�X0f��R��B�M�2�Ħ"�ˆ������߾)yľ񝳾߼���u����ɾ�.�y�������&�NM6��E�J,W�^<k������������䐿D7���v��1T�a2��E�0�(�n���B%���D���g�ߵ���u�������K��8���*u���_���M��t=���-����O%��r�� 8־!z��c������_��:Ӿ2��4
�2����+��;�8kK�4}]�br��'�� T�����\��+��o>k�4MH�|*(��f�H���3�-)�6m/��P��s�)�������(�����𮂿Yo���Z��I���9��8*�/����QEdѾ�1���h���2��Ⱦ��-[��	��d$���4�VD���T�b�g�V}��\���I������V��OC��ՠc���@��%#���E������ �b�=���`�l*�����P��k���wA��0���B�k�qAX���G�w8��*(���Ξ�@���?о,���H�����¾�־%󾊏
�_L��L-��%=���L��^��r�����0��܉��m��9ӌ��}���[��,:��=��7�P������-�q5M��=p�,�r���b5���Ӱ��փ}�`Ih���U�a�E��6���%��>����8R澀�ξgp��:����k̾L��� �����#��4���C���S���e�=�z��L���|���ᕿ�5���2����s�	�P�Po0�G�����,0�����7�,sX�#{��
��Ƈ��숕�u֏����]�u�ʥa��'P�px@���0�u ��w����p�ݾ_ɾ�X����þ��ӾHO�4��-n��)���9�:SI�0�Y���l��H������c꓿="��9�҄�S�h���E���'�����N�9a�_E%��VB�p�d��<������  �  �.^��d��5e���d���d��Ee���c���]���P��@=�:�%��������ݾ'�־��5N��V���g+�~8B�0}T�d�_���d�шe�fe��<e�Ğe���c�ny\�MBN�L�9�%I"��d����۾��׾�6�j�����v�/���E��-W��xa��oe���e��Ae���e���e�%c�O�Z�gK�r96��r�:
�Lb�**ھ�پV������w�3�Q"I��;Y�Qb��ge�tTe���d�-Le�~8e���a��MX�|�G���1��2��w���� �ؾ�ھ�z�R�	�.j ��Y8��wM�1�\��d�3g���f�_�f�-:g���f�0�b�kX���F�C40�p��,���x��iܾ���k���g���&�<=>�EvR�Yc`�'Vg��i�D�h�'�h��i�Ah��c��KW���D���-�my�O�|i��]߾���d� ����A,�F�C�L�V�{�c�[�i���j��:j��?j���j�>ii��Cc��GV���B���+�@q�.����%��<h�2}��/�	�1�Q�H�XB[���f���k�-ll���k� l�)�l���j���c�sU��<A��)�z�� �w쾇6�ؾ����
�>C ��8�lfN���_���i���m�hn�}�m�Y�m��n�[k�w�b�m�S�mR>���&��t���6�%�7a��%����#�E�;�.7Q��Wa��uj���m���m�,m���m�·m��#j�ɣ`�]%P�fI:��x"�H��;������&�������4���'�|�?�]zT� ~c��}k���m���m�jcm�$�m���m��Di��^��M���6������	�����Y�_��F�z�k,�C�C���W�#�e���l�9Fn�@�m���m�JLn�l�m�#Vh�a}\��I���2�Cm�~)�s��M�辕��~V�9�vz0��G���Z��  �  �Y3�h�B��S�\Ug��4}����/8��GD��ъ���{��Y��[7����-���O�ޞ��q ���>���a�"3������ʑ�D6�����\�x�Sc�+8P�q�?��`0��8 ����'���8�ھ����𕲾�˯�)�����ξE$��0�s���})�\$9���H�~�Z�wo�q���p?��񢑿�8��QY���Bq�wxN�F_-�v����������*��~J�	hm�o������B���B�������P-q��Z\�waJ�-~:�\�*��]�n��X��BѾ`Q���y���+��9��$�ؾ|���������	0��?�K�O���b���w�|І�"l��yƒ�Uގ��Ѓ��g�[�D���%�K��1I�2
��.���6��Y�sr{�!p���Ò�ޏ��(�������m���Y�~�H�9�MB)��_�,���i�1�о�A��Z���;b���&Ͼ,|�j����Y�(�=�8��bH��>Y��l��T��Ƌ�c�	 ����������n_�k(=�A� ���uh	������&��9E�Q9h�ㅄ�~^���3�����H������j��!W�z�F�ml7��c'��@�����꾢6Ѿ��¾����A�ɾ2߾,���@��4!�q�1���A�NQ�[�b��hw�?����_������'N���i��[y�,�V��k5���޿���W���2���R�Kvu��ꉿˍ��2Ε���������ky�%�d���R�o�B�`<3�"�"��%�������ᾛy˾Ai�������Ͼ�����J*�͑&���6��cF���V��2i��~��#��:������(%��v��3n��'K��	,���@����� ���<�m�^��o������c���)��D��� Z����r���^���M��A>��t.�f��Z��8V��ppھA�Ǿ���sƾ:�׾��
�����,��  �  �c�s�7�ًX�#g���s��p﻿�����ظ�����G���ah�6F?�e%�d��)�)�AUG��%s�U��`���Ļ�r����l��)��	����w�C�P�ɱ1�����o��8�lȾmɯ� t���͒��֐��]㦾����ؾ���xq��&��bB�+�e����Q���MԲ��+���Ŀ��޳��t��<ꄿW�Y�,5��*!�� ��2���T���V����̱�U�
���h���?���i��m�i�$�E�͘(��i��f���v۾d��Xר�����~���Ȓ��ܜ��ʮ�{0Ǿ�����A��-0�o�N�V�t�W[������θ�����V��m��5��:�z�GN��.��� ��v&���>��Uf�����;��
���P¿��xy��%a��Ä���`���>���#�ZX��^���$پJ⾾X����c������𜾏����׽�x�׾��h��v�"�W=��	^��#��J����*��?����vÿ���樿�#���2n�g/E��d+���#�-�/���M�k�y��U���`�����&EĿGټ�8���jz����~��W�e�8�*�����z���pN׾P�����������FW��tc����;�U�s��\���.���J�1.n�M<���⢿�󶿻Eÿl�ÿ�������q�a�R4=��0)�K(��:�	�\����0���wֵ���¿{�ÿF����&�������#r���M�Y�0����{���!�Ͼ���-'���P���T��e��������վ*�f�
������6�huU�%^{����O
��5���Ŀ�3������6������77T���4�P�&�W,��QD�0l�ю�b���ȭ����Ŀ����(������`^����e��
D��4)�����R��C㾐�Ⱦ�=���妾w������������oƾ�\�4J��]���  �  F��A;��bl��甿ʖ����ؿ��Q��0��$VԿ�������`e���B��8��?H�8Hp��)��9���eKۿ���Z����쿸ҿ��΍�4�`�%{2������h�žJ���!�� Y��Cx��Iu�Q��#݋�MZ��i۷���پ�t�8�!�V�J�������(yÿv��3������n���ɿKХ�������W���<��N;�+]S��Y��Rӡ��ſǮ俫���<����B忱ǿ39���H����O�d�%��:�ݾu���F����|�������v���x�	3��>�������ľ7��=����/���\�[���嬿�dϿh뿿r���,��{�߿�ľ��#����x��)N�ʾ;�O�B�AOc�����*���mҿ2�������*�ݿh�������v�� D�j���8��KؾP������H����
���G䅾{���/g�������־���G��6�@�a�q�;���P����ۿƛ����qW�\'׿�n�������Lk�ˉH�v�>��dN���v�hS��G༿��޿�����V���F𿿄տ�a���?��B�g��o9����:3���Ծ�g��xB���ɓ��݋�����,��QJ��3��Ⱦ�꾅��LN*�=S��G��˰��ѝǿ�������u����뿤�Ϳ�ة�}�����_���D�6SC��a[��\���ץ���ɿ*�迌���, ��=X�i7˿W��@j���X���-��]��(˾�ذ������	��j
��ы�W���q���/���GҾ������K\6��Qc�{j��7���ҿ������k���������Q=���~�2T���A�V�H�%i����������*տ-���B��_)�����P ���+����{��=I�"�"�"k�/�⾔�¾����5�������ދ��쎾��������{���޾���  �  k����E�����X���Yٿ߳�������a�%t ��Կ|��ヿ* \�r�O��<c�0����밿{޿w�����������u���$Ͽ�㡿wv���:�&����߾r���C������>�h�Q�Z��7X��+a�v��9��ޥ��ʾT���x�%���Y�Rȏ�]������	�l��P�=����,�ĿU����Rv��T��	S�Dq�x_���п����g�
����i��K�
�3��𙿿y���o`�hC*��*��NϾ)�	^��ty��Hc��Y�{[�p�h��X��sr��_ǲ��ܾKP�a�6�:�p�
����ʿ���#��}'�v{�ې���信���ܯ���i�lS�k�[��1���}����п���U��}���������q��6��鈿�P�7\�Y���ZȾ�o��������qn�8h���m��%�(����l��qeƾ����_��{K�3���{��7ܿc����#t��������ֿ`i���چ�� b��U��[i��ٍ��������������ܦ�~����ҿIT���^}���A�:��}	�	�¾�	�����������
z�Fx������d��G���ރ��4�۾�I��-��Ib������ξ��+�*&���Z��������u�ȿ���bZ~���\�M[��y�pb��3�ÿN�����ů�������n�1�ÿ(��<�h��2�'o�i�߾�U������U���������x�A<z�Q���H��᣾������� �4N=��?w�\��d"ο����V~�{�����'	���翖������n p���X���a�5���[��cVӿsX �e)�+�R����	��Ѵ�m����[U���$�����Ҿi������䅉�K���\�z�^���\���/���ǭ���ξ�����  �  �#��@P��>���ż����Te� &��i,���$�����G��N��
����m���_���u�����GĿNf�����'�)J,���"�� ���g����E��-C�}���Bܾ>�7����p��_W�x9J�u�G��@P�pd�G��dn���)ž2�����*�.?g��P��!�ο�����<�)��{+�'7����Q�ۿv8��h�Yne��ac��肿�g��g�տ���-���*���*�����B�ԿQT��6�n��?0����jʾ�����2��sg��UR��`I��%K���W��p��\�����B�ؾu���&>�ٳ���﬿v��#��&�!�mj,��F)����F �#˿�}���]}��c��Em�1ڍ�����n��b��L�#�&-��b(����n�����Ŀ�����\[��:#��������<���vⅾT�m��L]���W�j:]��m�'k��ΐ�������\�!����U�I���1���*�������l'�c�-�~�%�Q8�b*��=�������s�o�e��|�R��;gǿ˓����1)� �-�T�$�2���W����!����J�}��m~�?f��*��������v�'{i�E�g�&�p��`��	������Z�վ�_��.3�՞o��}���ҿ	��+����+�i�-��>!�N�
���߿'>��B����sm��ek�놿�j����ٿǬ�����,�ƺ,�P���(�ؿbt��P)w���8������ھ���sp������Vr��h�N�i���u�`����Ú����y澪��h�D�S	���@�����	p�	0#��
.���*�͙�L���4ο����}�����h�4-s��Ő�Wr��˫�nN�(%�x.���)��0�Δ���ǿN�����`�u(�>��̾ҧ��ӏ�����"Np�=~j��Do���B���yꤾ��ǾAg���  �  G���cT�r:���Yÿ������@-�`�3�|�+�=������Lտ�4r���3t��Ke���|��Ɯ��_˿���'S�w�.�j�3���)�#
�k�￴���BŇ�S�F�>��۾몾����~Ok���Q���D���B���J��^��;��r��;�þ;p �w-���l�����Lֿ���&t!�<1�|�2�]�%��+�B��
󯿏։��_k�W:i�?���㪿v�ݿM��#�� 2��2�V�#�~�[�ܿ�c��u�t���2�T�ɾcl��!u��a~a��L�I'D�2�E��QR���j�����稾��׾����OA�����ݕ���>꿌���x(���3���0�Is��d��ҿ����+����h��ws���@ѻ����}��վ*���4�"�/��:�6s�%k˿w7����_�Z%�����J7��-�����Lh��W��R�R�W��h�v�������[���:^�1!���Y�=���ƿ�G��9���.�(H5�w	-��>�p���¿�k���4z�	Yk��k��۟��~ο�=�����j0��t5� �+�b���>�����<8���yM��"����zb��tJ��S����p��*d�irb��k��%�ɸ������C�Ծ����}5���t��D��nuڿ}
�J�#�tH3�I�4��(�M1�h�翵���cڍ��ds�>q�f����宿���g�V�%��&4� %4���%���#��σ���|�;����xwپ�Ȯ�ᯒ��̀���l�,Zc�<�d��Zp�@*����������`���H��M��t浿[��	3��*�΄5�6-2��!����l�տ�����+���n��_y�������������/��,���5���0����p��ο�Ԛ�Ne�_E*��(��~ʾ�M�������{�D�j�#Ae���i��y�+��X��*�ž�h���  �  �#��@P��>���ż����Te� &��i,���$�����G��N��
����m���_���u�����GĿNf�����'�)J,���"�� ���g����E��-C�}���Bܾ>�7����p��_W�x9J�u�G��@P�pd�G��dn���)ž2�����*�.?g��P��!�ο�����<�)��{+�'7����Q�ۿv8��h�Yne��ac��肿�g��g�տ���-���*���*�����B�ԿQT��6�n��?0����jʾ�����2��rg��UR��`I��%K���W� �p��\�����@�ؾt���&>�س���﬿u��#��%�!�mj,��F)����F �#˿�}���]}��c��Em�1ڍ�����o��b��M�#�&-��b(����n�����Ŀ�����\[��:#��������=���vⅾU�m��L]���W�j:]��m�&k��͐�������\� ����U�I���1���*�������l'�b�-�~�%�Q8�b*��=�������s�o�e��|�S��<gǿ̓����1)� �-�T�$�3���W����"����J�~��o~�@f��+��������v�({i�F�g�'�p��`��	������Z�վ�_��.3�՞o��}���ҿ	��+����+�i�-��>!�N�
���߿'>��B����sm��ek�놿�j����ٿǬ�����,�ƺ,�P���(�ؿbt��P)w���8������ھ���sp������Vr��h�N�i���u�`����Ú����y澪��h�D�S	���@�����	p�	0#��
.���*�͙�L���4ο����}�����h�4-s��Ő�Wr��˫�nN�(%�x.���)��0�Δ���ǿN�����`�u(�>��̾ҧ��ӏ�����"Np�=~j��Do���B���yꤾ��ǾAg���  �  k����E�����X���Yٿ߳�������a�%t ��Կ|��ヿ* \�r�O��<c�0����밿{޿w�����������u���$Ͽ�㡿wv���:�&����߾r���C������>�h�Q�Z��7X��+a�v��9��ޥ��ʾT���x�%���Y�Rȏ�]������	�l��P�=����,�ĿU����Rv��T��	S�Dq�x_���п����g�
����i��K�
�3��𙿿y���o`�hC*��*��NϾ)�^��sy��Hc��Y�{[�m�h��X��qr��\ǲ��ܾIP�_�6�8�p�
����ʿ���"��|'�v{�ڐ���信���ܯ���i�lS�l�[��1���}����п���V��~���������q��6��鈿�P�9\�\���ZȾ�o��������sn�8h���m��%�&����l��oeƾ�����_��{K�2���z��5ܿc����"t��������ֿ`i���چ�� b��U��[i��ٍ��������������ݦ������ҿJT���^}���A�<���	��¾�	�����������
z�Hx������d��G���ރ��5�۾�I��-��Ib������ξ��+�*&���Z��������u�ȿ���bZ~���\�M[��y�pb��3�ÿN�����ů�������n�1�ÿ(��<�h��2�'o�i�߾�U������U���������x�A<z�Q���H��᣾������� �4N=��?w�\��d"ο����V~�{�����'	���翖������n p���X���a�5���[��cVӿsX �e)�+�R����	��Ѵ�m����[U���$�����Ҿi������䅉�K���\�z�^���\���/���ǭ���ξ�����  �  F��A;��bl��甿ʖ����ؿ��Q��0��$VԿ�������`e���B��8��?H�8Hp��)��9���eKۿ���Z����쿸ҿ��΍�4�`�%{2������h�žJ���!�� Y��Cx��Iu�Q��#݋�MZ��i۷���پ�t�8�!�V�J�������(yÿv��3������n���ɿKХ�������W���<��N;�+]S��Y��Rӡ��ſǮ俫���<����B忱ǿ39���H����O�d�%��:�ݾt���F����|�������v���x�3��<�������ľ2��:����/���\�Y���嬿�dϿh뿽r���,��z�߿�ľ��#����x��)N�ʾ;�O�B�BOc�����*���mҿ3�������,�ݿ	h�������v�� D�m���8��KؾS������H�� ��
���F䅾y���-g�������־���D��3�@�]�q�9���P����ۿě����oW�Z'׿�n�������Lk�ˉH�v�>��dN���v�iS��H༿��޿�����V���F���տ�a���?��E�g��o9����?3���Ծ�g��{B���ɓ��݋�����,��QJ��4��Ⱦ�꾅��LN*�=S��G��˰��ѝǿ�������u����뿤�Ϳ�ة�}�����_���D�6SC��a[��\���ץ���ɿ*�迌���, ��=X�i7˿W��@j���X���-��]��(˾�ذ������	��j
��ы�W���q���/���GҾ������K\6��Qc�{j��7���ҿ������k���������Q=���~�2T���A�V�H�%i����������*տ-���B��_)�����P ���+����{��=I�"�"�"k�/�⾔�¾����5�������ދ��쎾��������{���޾���  �  �c�s�7�ًX�#g���s��p﻿�����ظ�����G���ah�6F?�e%�d��)�)�AUG��%s�U��`���Ļ�r����l��)��	����w�C�P�ɱ1�����o��8�lȾmɯ� t���͒��֐��]㦾����ؾ���xq��&��bB�+�e����Q���MԲ��+���Ŀ��޳��t��<ꄿW�Y�,5��*!�� ��2���T���V����̱�U�
���h���?���i��m�i�$�E�͘(��i��f���v۾d��Wר�����~���Ȓ��ܜ��ʮ�w0Ǿ�����>�� -0�k�N�R�t�U[������θ�����T��m��4��8�z�FN��.��� ��v&���>��Uf�����;�����P¿��zy��(a��Ä���`���>���#�]X��^���$پM⾾Z����c������𜾍����׽�u�׾���f��r�"�S=��	^��#��H����*��=����vÿ�����樿�#���2n�f/E��d+���#�-�/���M�m�y��U���`�����'EĿIټ�:���lz����~��W�i�8�.��Õ����uN׾S�����������HX��uc����;�U�s��\���.���J�1.n�M<���⢿�󶿻Eÿl�ÿ�������q�a�R4=��0)�K(��:�	�\����0���wֵ���¿{�ÿF����&�������#r���M�Y�0����{���!�Ͼ���-'���P���T��e��������վ*�f�
������6�huU�%^{����O
��5���Ŀ�3������6������77T���4�P�&�W,��QD�0l�ю�b���ȭ����Ŀ����(������`^����e��
D��4)�����R��C㾐�Ⱦ�=���妾w������������oƾ�\�4J��]���  �  �Y3�h�B��S�\Ug��4}����/8��GD��ъ���{��Y��[7����-���O�ޞ��q ���>���a�"3������ʑ�D6�����\�x�Sc�+8P�q�?��`0��8 ����'���8�ھ����𕲾�˯�)�����ξE$��0�s���})�\$9���H�~�Z�wo�q���p?��񢑿�8��QY���Bq�wxN�F_-�v����������*��~J�	hm�o������B���B�������P-q��Z\�waJ�-~:�\�*��]�n��X��BѾ_Q���y���+��9�� �ؾx��������	0��?�G�O���b���w�zІ� l��wƒ�Sގ��Ѓ��g�Y�D���%�K��1I�2
��.���6��Y�vr{�"p���Ò�Ꮢ�*�������Ǌm���Y���H�	9�QB)��_�.���i�3�о�A��Z���:b���&Ͼ)|�h����V�(�9�8��bH��>Y���l��T��Ƌ�a� ������	����n_�i(=�?� ���uh	������&��9E�S9h�兄��^���3�����K������j��!W��F�ql7��c'��@�����꾥6Ѿ��¾����B�ɾ2߾,���@��4!�q�1���A�NQ�Z�b��hw�?����_������'N���i��[y�,�V��k5���޿���W���2���R�Kvu��ꉿˍ��2Ε���������ky�%�d���R�o�B�`<3�"�"��%�������ᾛy˾Ai�������Ͼ�����J*�͑&���6��cF���V��2i��~��#��:������(%��v��3n��'K��	,���@����� ���<�m�^��o������c���)��D��� Z����r���^���M��A>��t.�f��Z��8V��ppھA�Ǿ���sƾ:�׾��
�����,��  �  �.^��d��5e���d���d��Ee���c���]���P��@=�:�%��������ݾ'�־��5N��V���g+�~8B�0}T�d�_���d�шe�fe��<e�Ğe���c�ny\�MBN�L�9�%I"��d����۾��׾�6�j�����v�/���E��-W��xa��oe���e��Ae���e���e�%c�O�Z�gK�r96��r�:
�Lb�**ھ�پV������x�3�Q"I��;Y�Qb��ge�uTe���d�-Le�~8e���a��MX�|�G���1��2��w������ؾ��ھ�z�P�	�+j ��Y8��wM�-�\��d�3g���f�Z�f�(:g���f�,�b�gX���F�A40�n��+���x��iܾ���m���g��&�?=>�IvR�]c`�+Vg��i�I�h�,�h��i�Ah��c��KW���D���-�oy�O�}i��]߾���c� ����A,�C�C�I�V�w�c�V�i���j��:j��?j�}�j�9ii��Cc��GV���B���+�>q�
.����%��>h�3}��/��1�T�H�[B[���f���k�2ll���k� l�.�l���j���c�sU��<A�	�)�|�� �y쾉6�ھ����
�?C ��8�lfN���_���i���m�hn�}�m�Y�m��n�[k�w�b�m�S�mR>���&��t���6�%�6a��%����#�E�;�.7Q��Wa��uj���m���m�,m���m�·m��#j�ɣ`�]%P�fI:��x"�H��;������&�������4���'�|�?�]zT� ~c��}k���m���m�jcm�$�m���m��Di��^��M���6������	�����Y�_��F�z�k,�C�C���W�#�e���l�9Fn�@�m���m�JLn�l�m�#Vh�a}\��I���2�Cm�~)�s��M�辕��~V�9�vz0��G���Z��  �  �V��ꏿ�����{�X0f��R��B�M�2�Ħ"�ˆ������߾)yľ񝳾߼���u����ɾ�.�y�������&�NM6��E�J,W�^<k������������䐿D7���v��1T�a2��E�0�(�n���B%���D���g�ߵ���u�������K��8���*u���_���M��t=���-����O%��r�� 8־!z��c������_��:Ӿ2��4
�2����+��;�9kK�4}]�br��'�� T�����\��+��o>k�4MH�|*(��f�G���3�+)�4m/���P��s�(�������(�������Xo���Z��I���9��8*�,����MEdѾ�1���h���2��Ⱦ��/[��	��d$���4�ZD���T�g�g�V}��\���I������V��QC��נc���@��%#���E������ �`�=���`�j*�����N��i���uA��-���=�k�lAX���G�s8��*(���˞�=���?о+���H�����¾�־�%󾌏
�aL��L-��%=���L��^��r�����0��މ��m��;ӌ� �}���[��,:��=��7�P������-�q5M��=p�,�r���b5���Ӱ��փ}�`Ih���U�a�E��6���%��>����8R澀�ξgp��:����k̾L��� �����#��4���C���S���e�=�z��L���|���ᕿ�5���2����s�	�P�Po0�G�����,0�����7�,sX�#{��
��Ƈ��숕�u֏����]�u�ʥa��'P�px@���0�u ��w����p�ݾ_ɾ�X����þ��ӾHO�4��-n��)���9�:SI�0�Y���l��H������c꓿="��9�҄�S�h���E���'�����N�9a�_E%��VB�p�d��<������  �  ���}F��V��=����k~�!�V��6�:��=�Z��:_̾Ҳ�}Y��LW���揾�`��;���=���Ӿ�����J�!��<��"_��<���䚿�ů�h���_x��A����d��n#���a��:�O%#���W�-�hN�T�{����,���袽�����8=��ʤ�ZZ����p�F|K�Y-��R�y��o;�@4ľ�|��!L��G���%y��Wƙ����1��U�ݾ{�������-*�уG��$l�騋�>7��w[����/e��d������Ox��UR�(S0��y���!���6�8v\�s����,���M�����Nm��ꓲ�[<��.���&e��'B��H&�
��ǔ����ھNv��p
��/��������E��񰣾϶��O�ϾYH��Aa�'�6�seV��~}��
���
��n廿��¿���ū������yt�mI��,��8"�;�*�+�E���o�t/���⩿�5���tÿ������yg��l򁿻\���;�˲!����� ��{�׾�]������Y���(���⡾�����>ž0Hྏ ���}�(�)�C�f������S���7��;��wĿJ,�����L�����h��*B��V+��*'�H"6�Y�V����"����岿U�����Ŀ t������1����Fy���S��5��~�Ϋ	�o��YԾ^���_����ń���ҩ�M(��8/Ѿã�+u����S2�I�O��]t�`ʏ�G]�������Ŀ¿�ʹ��L��������Z��8�}�'��)�d�>��3d�@[���ӣ�ظ�DĿ��¿�鵿Ѝ��G㊿d�k���H���,�V������p�V̾�x��oҧ�#q������!������ �ھ6��Z��"�k�;�[�{Z��⨗�D���D����Uſ����LS������ey��AN���1��&�zw/��UJ�v-t��R�����r>���  �  ��G�￹׿��������`i���8�Nr�����ʾ�,��5���=���w�x���s���{�_Έ��3���|����Ҿ����%��%�B�N.v�в������J�ݿ���e����O뿥Ͽ-���T����H^��k?�w�9�Z�M��ay�����Ŀ��@࿍��3R���`��̿�3��X����gX��$,�4����m���ʤ��p�������w��Kv�+����u������׳���'ྼ����'�X�R� ���$��%�ȿ��濟O��? ��}�&ÿP����5�?Q�i|:� w=��Y�<e������˿V�5���������� M¿�\���i~�a�I���!�����۾?߹�`
���4��G�Э~�8����k���ޙ�� ����;����1��S"8�,g�UV��'���ܖտ(�����a���ۿ����R��K�q�k K���<�YH���l�g�/����ؿ�6�y���ܞ�D�ٿ`���Ε��n�*q>����'�����վ�������]w���f��k��G}��D����;���OM྅��W�"�U�I��}�t!������I῞&��9N��2����ҿ���=����if���G��B�aV��퀿�C��	Ŀ\��8J��č��\��ѿa���Ì���`�\4��7��Z��%�о(�!����ǒ������1��Ӎ������n����̾�T����/�O�Z�m���F���Ϳ��&~��uQ��?E��ǿ�䣿)Ƀ�iY�-�B�țE��a��N��Ы��nϿ����G���G���忒�ſ
���E���mP�&(�):
�m辇�ƾ�������P$��DG��:3��%ؕ����x���Qlؾq�������W=��_l���[A��j7ؿ�]�e���I��R޿y���Ř�Awv���O�{A�s�L�q�2'��&-��+�ڿ�A���  �  ���������ֿ騿e怿C����6��6��ߙ��փ���j�Y�Z�"�V���]�up�D:���P���%þ���j�6�O�7=��%���oE����s�0���A�e����̿�꠿��~�O*X��Q�8�i�ww��>]���O�k���C��a��m���{ǿh����{k���2�R	� �׾0�����_Z~�x�e���Y��Y��c�s�z��M����(Ҿ[$�V�,�<d�_H���&¿7W� ������;�*�	��*�` ���/��]<n��R��U�'y�����ǿ������j�����u�I<�eܸ�|_���X�h�$�������˾�Χ����|��Qi�'�a�wge�ݾt��M��ݰ��<���1�K��@��}�� ���zӿ�C �������G����ݿ'������i�e�a�S��=b�)Շ��'��8ٿ����Y�\m��X����QٿW���7����H��R���ž�5���`��F=��V�r��o��v�h���E��@�����о=T�G�$���V�m���c��ݲ�T���0���������{lп<��z���}`��xY��Vr�i��������P=
�Ң�H��C��ܟ���˿�%��Ⱦs���:��K����!��-����H�������y��/y������l��ٟ�����U�yB� 5��6l��e���HƿB~�����n���T�Y��_�&U��b��>�v�ZQZ���]�����ǧ��{˿�V��ʮ����~�X 
�	�꿿+�� ���p�^��L+�a���ؾn���e���d劾�ۀ�p�y���|��Ʌ��x������%Ǿ���`���F��y��뛨��ֿ���6��!I������\�5��cz��%Yj��X���f���`���Eۿ���[`��  �  �f,�GK%������I蹿>튿[�L����0j��Ⲿ����Du�CaY�)VJ��KF��L���^�$�}�£���Ҽ����CI"� �[�����ƴſBE��vC�+(�H+,�D"�P��Xm俛����Њ��Ai��a���}�(�����̿,B�߹��`)�Ŀ+��- ���	���ݿ1{����{� �9�Ee
��]Ӿ)��n\��%l���T��bI�ݾH�q�R�-�h�В���Ԣ��4;���R3�is�����ȝ׿h�}�j+��<*���a��~ҿ㢿�M��8b��cf��z��̶��V�޿�)
��n ��,�0�)���/��ԁ̿�����d�6�)�TY����ž�H��_�����j�sX�;]Q�O�T��Qc��C~������a�����:����I�=���$��Է�^�.�$�YM-���'�����^��J�ÿ���rx�X�c��/t�n;��(X�����@b���&���-��&�js�Ȩ��������LR��A�cs�����J���,��Y�p��ab�v�^�&�e�tGx�H���餾THʾ�� ��!)��ab����H"ɿK������x�)���-���#�7���Y�H���w��q���i�����Ң�I0ѿ:d�����+���-��I"�D�⿔���������A����T���7��+���N.��!�t��i���h���r��]��
���b����aݾ[
��y;��={����ۿ		�d! �L-�'V,�� ��6�h�ֿP����o�j�]�n�Q���鯰�������:"�;�-�`+����9���ϿU؝�o�k��.0�wB��Ҿ�+��ih��񁾅�p�$=i�=l��#z�qK���������S��m���N��֊�)����U����%�>�.��)�b��������ſ�j���|��h���x�r���	�������4q�=�'��  �  O�=�3�˿"��t솿z�N����xT꾕沾PQ��ZBd�?�A�-P,�\� �6��ֺ"�<r0���H��n�
���������F4&�U\� ����*��KcҿI��~�Q3࿻ſ���xO���Q���3��(.�UjA��k�J����]��b�տ���%�쿟�ݿm��)����<x��<����־ot��]i����X�N6;��2)�x �;���'�vs8��T�a'��%����оAr	�:�6���p�Zu��U����ۿ>��F�꿵MؿJ���ԏ��UQq���D�Y�.�<�1��4M�me~��������^R޿#1� 5��Dֿ�嶿x�����d��b-�����Ǿ���Ĕ|��(U��7<��.�,�(���+���6���K�m��Տ�C��p��?���9L��������1ʿ@$俦/ￄ&迎ѿ!��������Ud��?��J1�q<��w_��V������Pοo�濱����kjοM߬�m���K0T�'!�"L��W�~����z���X���C���8��56�F�;���I���b�$���m��x�˾I��|-���b��*������q�տvw������k�ȿ��DD�� �Y���;�zu6���I��t�h5��ϔ����ٿ���m��[�w�ſ�����>��,E�A?���F�������(y��L[�*:I�v@���?���G��tX���t�w6���Ѱ�1�Y����>�o�x�Ő�����.0߿)�￥�xܿq"��ֹ��k�y�M�'7���9�T-U� ���W����ſ��ῷ��E��t�ٿC3���Ж�'Ck���3�g	���Ծ: �����(jn��U��fF���@���B���M���a�zx������j���������mQ�������?�̿m��G����V�ӿ���_
���&i���C��5��A���c�ڎ���=���mпf���  �  t3�)�ۿ2CĿ~k������j�I�]#��|辘'��ƍ�kOh��+F���0��$�0�!�\�&���4���L�1�r��J���彾x��3#���V��j�����̤ʿ�(߿V�R�׿S���4���s�|���K�}k/��*�J�<���d��J�������Ϳ@����,�տ]����r��iq�3�8��#���վ2������8]�+�?��q-��$��$�8�+���<���X�[큾1���I@Ͼ���	3��Qj������඿��ҿR����Eп{o��D���fj���?�#�*�b�-�R�G�O�v��P��1 ���ֿ$��L῏^οG�������G�^��#*��m��>ǾV)���.��Y�#�@��C2���,���/��;��P�.q�a��K|����辻9�ӤG��O��:����¿B�ۿ	�fi߿�ɿ����{9���)^��o:�oI-���7���Y�:#��I��5�ƿAD޿a�濵O޿� ǿ�(������APO���(t�;4���򘾼�~�_>]��"H��<��J:���?��MN���f�����c���Vk˾���j*�Du]�TՍ��y��ο��⿕��@hۿ���ᆡ�w^���T���7�h2��D��dm�r���h;��!�ѿ��7��ۯٿƶ��#���©y�MA��O�� ��c���?���b}�I�_�(yM���D��D���K�t�\���x�Z��������h߾��~.;�6r�ݥ��n ��a ׿���忧oԿ0����ؖ���r� H�W3���5���O���~���������ٿ4����C�ѿ峿�I��se�Q�0�D��VԾ�#��� ���r��aY���J���D��G�z�Q�p^f�ԇ��O!�����}�8p�v�L�}ꃿ~4��ſ�3޿ڮ�F��I̿�������j�b��.?���1�ۖ<�4^��Z��`s���ɿ�S��  �  ��˿�/Ŀ�G�������p�i'=�O��k��r��-C��|v��[T�26>���1�(w.�(�3��B�2[�w��$A��m(���I�Ԭ��9H�U�}����������Eǿ�i˿������S׎�)]g���<��o#����3/���R��_��Ƴ���@��T�ȿ�˿�����%���zV_�͂.�ە�k�Ծ�ͩ��:��]Ik�ɥM���:�Z1���0�^&9�>�J�gg�|5�����̴ξG���q)��2Y��b���ि�ü��2ʿ_ɿ�s��¡���M��)@W���1��q��!�k9��Hb�c����<���}��7�˿�6ɿ���ѣ���炿(�O���!�����B�ǾHӡ�����7�g�hkN�A`?�R�9�u�<� �H�1^�������>���O�����;�o�n��Γ�>r���yĿ;pͿ�ǿ�괿:���j|��M���-��"�1~+��I�$w��w�������ƿo?ο��ƿl��gԗ��[v�@�B��U�������o��=Z���mk�E�U��I���F�{�L��\�{+u��-��������̾������"�O�%G��>���1��Ǿʿ%�ο �Ŀ�x������:o���D��+�_'��`7���Z�����x颿zv����̿�8Ͽ�9ÿ3���叿�g�θ6�t�����)����\��������m���Z�~WQ���P�� Y���j�G���2D��5�����޾"��U�1�H`a�~��  ������5Yο~�Ϳ1���&˥��u���_�c#:�ؚ'���)�o�@��j��y嫿
ÿ!Ͽo�̿�b�� �74���*V���(����վ^ͮ�����iz���9g�K�W��^Q��S�$b_�u�t��u��١���¾u������@���s�Uk��+��$ǿ�
п�Jʿ�t��M���~�����Q�v_2��&�0��M�N�{�5���Oٴ�M�ȿ�  �  ���r���u��O���C�U���-����b徚彾�ӟ�Q㈾�Zo��W�B�H���D��WK�0�[��v�𾍾W0��q1ƾ;�-��"R6���_�ʅ�ի��A󦿆���4����<���Yt���H�i&������b��18�x�`�3����ߚ�˯��ȩ������A��\s��>H�c"�3���ؾ1��,|��熃��h�!�R�XH�3sG�p#Q��d��`�������I���:Ӿz� ��`��rC��$n�2ь�;���[ ��O�������	���%e���;�x�������b�#�^E��o��_��,����C�������_���	���)f��g<�����a��{0ξ.d���m��1���th�?�V��P�W�S�r9a���x��f���飾YR��H��!�dk-���T�c8��hI��5B��C���hc������X�����Z�&v4����L��{C��Q1���V�.����
���զ�����!L��3���{��~[��3�		�CY�w�Ⱦ�����9��_6��z�n�R�`�o]�|Rd�ju�O>���S���U�Ӿ���sg��)=��df�~6����Wl���~��oF���򓿶�{���P��d.�m�M��#�_�@���h�,􊿉��k㫿����!�
l����{��~P���*�����Y�P3ľ�����������ys�<h��kg�q��x��ef��װ��dc��b����&���K�bZv�,�����E��lv�������0��qom�:D���%�b����j{+�*�L��{w�����6�����L���!����X��1�l�mC��|��F�ZH۾z]��>��\9���n���Ho�t�g�A�j�Hx�Ψ��[��ମ�o�˾�M��Q�G�2���Y��Ԃ�|痿৿�������+��<��	�_�iK9�Ӵ��+�]����5���Z�᥃�D#��U⨿�  �  m��N<��$�t�ŤY�{�<�3�!��0��:�mOҾ�̷�|ᠾ����!#~��l�#�f��/o�=���ԑ�����_����.پ�_���!���'��JC��o`�o�z��х�1P����H6h�1�G�zJ'��4��1���Y��;�������8�$FZ�:�w��~�������灿�l�=�P��3�_��%��l�ʾ�ǰ����0���x��j���i�L3v�`��̧��������ƾ���7����D�0��L���i�������F�6Rz�<�]��W<����ɞ��W�����:5��~$�˦D���e��a��q���?!���~�ILe��CH�m,��[�a� ��^��ľE���n��a��2{�r��ev��ك�9���;�����X־K�����3�"�lB=��BZ�rv��c��	q��ɫ��y~u�S�V��p5�t���q����V7����'�2�϶S�z|s��l��$������rbz� _�_	B�`G'�M���0���Zݾ(�¾p8���=��[Ҋ�s��nc�������KǞ�����˾����}�J��^�.��#J�3Jg������J��%׊�	���O�o��:O�\/�"!�̨�J����� #��JA�U�b�w%��n�������^��YNu�O�X��<���"��P�����Iھ�������:��GD���@���؄����_��謨�����־@��G�
�r��x�8��)U�3�q�aք�Z>��	���N����e���D�:�%����;�+�����,�hL��l�i惿���8���7����k���N��3�4����u�B�Ѿm���	��Ĕ���������s݆�8F��6i��R3����ƾ��྅b������(��wB��{_��?{����O��DA��d�z�l�[�f_:�ޡ�:2
�X�������4�6�F�W�<�w��w���  �  ~�R��Q���H���;�0-�9������q��C��N�Fgƾ�m��+񚾅���񊾏����䞾����XY̾)�f��}<�o����"���0��?�d�K�wOS�%rR���G��P5��.�1!���-GҾQξH�ܾ�9�����tm+�w�@�[O��DT�R0P��ZE�X7�>+)��J�����!�
򾘂ؾn���7��hȖ�; ��!���<9��٥�E,���jվD�ʨ�!"�����f'�&r5�0�C�I�N���S���O��SB�#�-�� ��" ��`߾��ξ5IѾ>��V�LQ��3��qG� $S�M4U�\�N��VB��4��8&�v���_����'��Ӿ�޺�Vɥ�5���T���&q���<��9[��UCʾ�)�C���=�
��S�?"��w/�[�=��kK�hU�!JW��P���?���)��N�����W�߾^�վP3޾����~��(���>���O�nlX�KLW��[N��A�<�2��J%��N�1���'��F뾥�Ѿ
���ر��r���&�����7�������hzپ|�H�	�ŋ���)���7�`�E���R��AZ�w}Y��"O���<��%��������G��J޾�,�e�����3��I�{W�ˣ\��X���M�9�?��j1�x$�:���B�W"�����!ϾA���ʦ��������5���׵��0̾_w���|���<���"��/���=�:�K��/W��/\�aX�L�J��5��Y��N����Y�޾��=�������#��;�:sN���Y�U�[��@U���H�{�:���,�Vp ����\	����uM�ytǾ�'���#���|��/��w�������S@վ����)�z�h��yr'�A�4��C�,�P�7OZ�)�\��2U��D���.�@����+U���޾JQ��� ����X,���B�bT��  �  &���*��W,�vu,�!{,�[^,���*�b�%��Y����Q���r۾�迾�0�����(0��Awž��������W�'���+�k�,�7�,�g�,�u�,��*�B�$���I��`���׾׼�]�����Gk���rʾ���#�2��r!�k�(��>,��-�-��-��,�%*��#�m����	����XҾɛ���Ы�J���i���Ͼ�0����v���"��s)�M,�4�,�4�,���,��,�_
)��!������쾨G;6U���ݪ�����Lg����ԾR����
|��n%���+��$.�6�.���.�2�.���-��*�06"��������;;�������ն��FnþW^޾�2��hE�Q��S�(�G,.��0��S0�P0�-F0��/�F�*�b$"�k
�������(V̾��kɱ�@����ʾ���"�����8"�u�+�,Q0���1�l�1�L�1���1��90�vP+���!��%�o��;���˾�(��7��C���=Ҿ���������%�BX.��w2�t�3�e�3�,�3��3��1�"�+�W�!����D)�M澚o̾���=����ľ4�ھ@S��yz��/�sx)��%1�-�4��b5�'V5��V5��4��N2�<�+��� �V�����a⾂�ɾ�ͻ�7��:eǾ�߾14���������*���1��n4�L 5�?�4�� 5�8\4��L1�?%*�e\����yf��$�ݾlƾQ����A��'�ʾN��<�����ov!��E,��o2���4��05�,5�-25��K4��0�|�(��@��v��v����پ�.ľ�����f����ξ��}�t��+�#�x�-�%c3��L5�Z�5�i�5��5��H4�b0��Q'�h(�9
�y��־�r¾������ |Ӿ%��N�����G&��  �  ���f�6| ���-�:[<���I��6R���R���I���8���!�p
��|�)Ծ��̾%iؾ�^������:'��+=�M�)�S�*Q�s9G��9��9+����K����y���d~ܾ�¾kw������k�b勾X��"����6���:Ѿ�������h�f��bn%��S3�z�A��M��T�n�Q��E�E�1��Z������mkо�UϾ���1g����4/�#�C���P�bT�p�N�j�B�{�4�+�&�"��_�;��dI�W�Ӿ�������f��������]��4���u���}�۾�����6���a�Jd+�O�9�]�G��/R�b�U��7P�/aA��,��v��h��ྕ�Ҿ�%ؾ���}%��v"���9�G�K�nV��{V��N�$�A��d3�Y�%�����2���B�q�Ҿ�f���+��落�z����!��VG���`����Ѿs��K���f�V����%��l3�T�A��O�שW�waX�]�O��>���'�"8�a?��C྆�ؾ���=� �z��Ҽ-�G�C���S���Z�c�W�7N��]@�2�s%�p=�"��{�J뾬�Ѿ�����x������꛾�V�����;�Ⱦ�ᾟ����+
�,���E!�[�-�j�;���I�+�U�.\�ݬY���M�d�9��c"��������g��O߾����e	�a��a97�ǍK�+�X�\�,�V�8K���<�<�.�41"�̝���Ⱦ�� ���ʾ�ȴ�2���w`��p�������c���uо��I��Y���K�H%�D2�}C@�h5N���X��j\���V���G��b2�"��\�� 쾨�޾N��c��J��b�'��?��RQ��R[�ݲ[�3�S��F�"�8�++�Y���i�Ϸ�7�����ܾ}Pľ�⯾�&������3��� ���¾�9ھ���8���  �  ���d>��&#��!>�(F[�/Mv�'���hp��'X���l�L�L�,�������9�������33��{T�;s�K?������{/��q�6&U�<8�@�`0�4h��QξTm����������{��k��h��s�Gt���0E���¾��޾	�����c\,��`H�}be��h~�h���↿d�~��;c��5B��~"�|�	�Ϗ��$����ND��k>�_�_��{��S������:���8h�jZK�Y/�T9����ږ�<ž�n���h�������ku��j��*l��v{�5K����������;���ގ�����6��S��o��.���s������Hx��aZ�)9�Ia�T;�����	� ���S�+�\uL��l�|��/��$5����|��Rb�0E�a�)�c�����`�޾Y�þ�z���ј������y�1�x�;�i/���d�����oþ;_޾���5��ޡ(�g�C�^�`���{�}`��t-��.���kr���R���1��w�� �\���\�tJ�m�9��Z��y�M���P������6�w���[��?���$�c!�q���ܾ��¾$ᬾ�����3��{���C��D���ZC�������׺��@Ӿvg�@F��Z���4��P���m��M���Ɋ�k񊿯Q���Jk�2>J�h�*�����E� �����B'��lF�/�g����)\��~��jJ��p`p�B�S�o=7��r��	��
�1zվ5Ƽ�
���X���c���!����|���֌�N��S(��-%¾R�۾sK��!H�s�#�z=��@Z�ٖv� y������\@��<�~�v�`��c?���!�"F����ǈ����Ll1�lR��er�MÅ�2����Љ�V����g��eJ�g/�_�����=龕ξ�������E��>�����ؓ��K��� ���y���˾v��  �  D��f ���/���W��������y2��2�����lm����{�vlO�a�*�����0�U���$2���X�*Ⴟ��O������Ϣ�1t��oz���N�>�'�T"��޾� ��a?��aT��+�k��_U���H�זF���N���`�f+}���������<�̾������=��g��{������'V���p���`���Ҍ���l�y�B�3"�(�3/�&9�
E>�"�g��a�������Ũ�"6��a���n�k��0A��u������о|^��U'���L��,�c��P��H�s�I���U��l��,��Ǜ������ܾ���$�%��L�=Uw�7'��lM��#̪����vԚ���,&`��o8����?��%���*�-�M�M�y��撿G���⿫��&��l���R��S�`���7�i�����!�˾�*���N���b���Ek��[���V��[�nk�$?�����V���{Lʾ���L���#5��r]�鲄�<���맿xҬ�L^��{<�������9U�Z�0�����>�D��E^8�C_�$��M���i���u��o3���ܕ�C�����U���.�;����7Ǿ�������p��;t��h��Kf�[�n����E ��3~������ݾ���n!�fYE�[o�/���$����i�����[k��ڐ���t���J�>*��%��+��5'�%CF���o�d��7���Yͬ�r���`E���Ǐ���s�dI�1�$��@�85ᾂ���pr���y��1ԁ��_p��<g��mh�L�s����N����੾��ž�~�5Q��b,�R�R���}�_r��~������uV��0��`���hYf�g�>�v�"�v2�H��j0���S��Y�4���Ϊ���b�� ê����눿V�e��<����5��}�վ�j���h���N��ж~���n�_&i��m��|��֊��j��$ȳ�LaҾ�  �  �����G�?�V�s�����Z���ſK�˿�lÿ�׮�o���o�GJB�P�%�����*��!K�Z{��ؙ�T��Րƿ��˿$���	F���t��wh���5��*���ܾn���M��{�p��FQ���<���1�f0�t�6�7(G�W�a�W���'��y%Ǿ���0�"�0�P������s�������ɿ߾ʿ�����c���,��}Y_��-7�!G!�� �;3�RZ�� ��O��������ɿQ�ɿi���-h��b͆��IV�>'������˾�w��8����e�>�I���8��1��#3���=�͵Q�j�p��������e�پ<�
��e2���c����I������O̿�ȿv����"��恿WR�Q�/�h� ���&��.A�8�l��ߑ�n����nÿ09Ϳ�Oȿz3��c͛�~��I�%�6��ľ���l���R�i�� R���D��!@��D�R�Tli�p.���&���0¾���#W�+9E�Foy�Bl���a��A�ǿ�RοK2ƿ;���QK���Ou��/H�.�+���#�Ƿ0�TQ�Ҁ��
��/���D�ɿh�ο?0ſ����ߓ���n���<�p�����ѽ�
��� ��;o�[[��
Q�ߤO�r
W�;�g��.��yՔ������׾Q����*��#Y�@އ����������'Ϳh�ο¿�j���0���\g��-?��D)�(�i�;�0b�� ��Q�����W�Ϳ;�Ϳ/˿��z���㊿�{^��:/���	��;ܾг��������i�~X���P���Q�@�[�	o�����׷���廾vk�P���9��gj��j��0����Ŀ_Ͽs̿^"��D��O����nX���5���&��,�3�F�l�r����Xq���ƿ�ϿG�ʿ|̸�;f��r���0<N�XF"��P �"wξ�O������AY}�8qe�5�W���R���V�O�c���z����s\��Dʾ�  �  *��io���L�Ä��L��D�ſ��ܿL=係�ڿ��¿������R��H2��)� �7���\�鉿�j��H%ɿ�_޿�#�m�ؿW���^���<�{��@A�����޾\���z����b�T%C��[/��%�VX#�M�)�cF9�vkS�B�{�Ѧ��Ϳƾi��T1+��`�f�������ϿJB�;8��XԿ��fG��+�s���E���,���+���A�֙m������\��<�ѿMH�O>���ѿ<&��������f�PB0�<��|̾
R���[��\�V���;���+���$��k&�o[0�"�C���b�?���g����i۾ƪ�y=�Zv�<�����
~׿<�俍���3Ϳ�6��ɘ���wd��D=��2,���2�Y�P�ic���򠿫.��Frڿ������ʿD򫿼U����V��@$����P�¾����J���I[��GD�j�7�]u3�@�7��{D��<[�D�~�ʙ�	%�������� ��VR��������ȿ�B߿/�濿�ݿ*�ſॿ���iX�vA8�/�Y�=�f�b��������a̿G���y�`#ܿD�¿Ca���;���!H��z�����Һ��㗾[$��ra���M�a#D�p�B���I�S�Y�]t�zP���5��C[׾O
��3���h��7��tǵ��&ӿ0U忄F�cؿN���@K��J�{�A�M�R�4��3�:�I���u�Ġ���^��n�տoO��H�r�տ�8��eƗ��"o��v8�����tܾ����`����!w��[�TEK���C��D��8N�:�`�lW�A���Z}���辸_�G�C���|��b��tW����ڿ���A��]п�U������ʋj�qGC��$2�f�8�Y�V�9>������1�ÿ�"ݿr}近��+wͿ*���)���3\��y)�ϯ��̾)5��Qቾ�"o�Q�W��J�|�E�G�I��V�cl�_��������7Ⱦ�  �  ����U�Q��ψ�����_Ϳg>�lX�%S�lʿ*����;��sXX�6�6�?-��6<���b�;\���|����п�'�{<�D��ƿbb���}����E���Fk�!���ㇾL�^�v�>�v+��� �A�*�%���4��O���w�풚�z0ǾE���.�!�f��������$׿�2��@��ܿ����m����z�K�3 1�|�/�t�F���t���������&�ٿE�a=�C�ٿ����]����Am���3��5�/�̾{`���}�o�R�Xy7��'�a� � U"��,�T?��}^�!���)	��X�ܾ����EA��[}��O���Ŀ;�߿/�����*տDy��8���k��
B��:0�l<7�IsV��Z��?u���Vȿ��⿄������ҿ��������bP\�$'��@���¾\�����{�R�V���?�OW3�*`/���3��,@��V�ݹz��a��k���{����#�`]W������֮�Uп���m���̿����%��?^�֩<��3��OB�w
i��|��.���F	Կq꿋��6��\ʿ�ʧ��鄿X�L�v��Dj�sO���K��6|�ã\��I���?�U�>��E�kFU�=�o�aq�� ����׾�����6���n�ט�i.���ۿ�E�O�>��b�ÿ�p���~���S��9�ٶ7���N�A�|�����k���H�ݿL��Gￛ�ݿ�п�����ru��<��i�9ݾj���MɎ���r�PSW��G��?��@�w�I�ʑ\��"{�i���ҷ��%�2h�1�G�t���䙤��Oǿ#㿵 �{��1.ؿ����K���q�<H�U,6��=�6A\��5��$C���˿b��T���}�'!տ�-����a�],�����̾�棾eꇾ4�j�dS�zUF���A�ŒE��Q��h�����M���
Ⱦ�  �  *��io���L�Ä��L��D�ſ��ܿL=係�ڿ��¿������R��H2��)� �7���\�鉿�j��H%ɿ�_޿�#�m�ؿW���^���<�{��@A�����޾\���z����b�T%C��[/��%�VX#�M�)�cF9�vkS�B�{�Ѧ��Ϳƾi��T1+��`�f�������ϿJB�;8��XԿ��fG��+�s���E���,���+���A�֙m������\��<�ѿMH�O>���ѿ<&��������f�PB0�<��|̾
R���[��\�V���;���+���$��k&�n[0� �C��b�=���f����i۾Ū�x=�Zv�;�����
~׿;�俌���3Ϳ�6��ɘ���wd��D=��2,���2�Y�P�ic���򠿬.��Grڿ������ʿD򫿼U����V��@$����R�¾����L���I[��GD�k�7�]u3�?�7��{D��<[�A�~� ʙ�%�������� ��VR��������ȿ�B߿.�濾�ݿ)�ſॿ���iX�vA8�/�Z�=�g�b������� b̿G���y�`#ܿE�¿Da���;���!H��z�����Һ��㗾]$��ta���M�c#D�q�B���I�S�Y�]t�zP���5��C[׾O
��3���h��7��tǵ��&ӿ0U忄F�cؿN���@K��J�{�A�M�R�4��3�:�I���u�Ġ���^��n�տoO��H�r�տ�8��eƗ��"o��v8�����tܾ����`����!w��[�TEK���C��D��8N�:�`�lW�A���Z}���辸_�G�C���|��b��tW����ڿ���A��]п�U������ʋj�qGC��$2�f�8�Y�V�9>������1�ÿ�"ݿr}近��+wͿ*���)���3\��y)�ϯ��̾)5��Qቾ�"o�Q�W��J�|�E�G�I��V�cl�_��������7Ⱦ�  �  �����G�?�V�s�����Z���ſK�˿�lÿ�׮�o���o�GJB�P�%�����*��!K�Z{��ؙ�T��Րƿ��˿$���	F���t��wh���5��*���ܾn���M��{�p��FQ���<���1�f0�t�6�7(G�W�a�W���'��y%Ǿ���0�"�0�P������s�������ɿ߾ʿ�����c���,��}Y_��-7�!G!�� �;3�RZ�� ��O��������ɿQ�ɿi���-h��b͆��IV�>'������˾�w��8����e�=�I���8��1��#3���=�ɵQ�e�p��������a�پ:�
��e2���c����I������N̿�ȿu����"��恿WR�Q�/�h� ���&��.A�9�l��ߑ�o����nÿ19Ϳ�Oȿ|3��e͛�~��I�(�6��ľ���n���V�i�� R���D��!@��D�R�Pli�n.���&���0¾��� W�)9E�Coy�@l���a��@�ǿ�RοJ2ƿ:���QK���Ou��/H�.�+���#�ȷ0�TQ�Ҁ��
��0���E�ɿi�οA0ſ����ߓ���n���<�s�����ѽ���� ���;o�	[[��
Q��O�t
W�<�g��.��yՔ������׾Q����*��#Y�@އ����������'Ϳh�ο¿�j���0���\g��-?��D)�(�i�;�0b�� ��Q�����W�Ϳ;�Ϳ/˿��z���㊿�{^��:/���	��;ܾг��������i�~X���P���Q�@�[�	o�����׷���廾vk�P���9��gj��j��0����Ŀ_Ͽs̿^"��D��O����nX���5���&��,�3�F�l�r����Xq���ƿ�ϿG�ʿ|̸�;f��r���0<N�XF"��P �"wξ�O������AY}�8qe�5�W���R���V�O�c���z����s\��Dʾ�  �  D��f ���/���W��������y2��2�����lm����{�vlO�a�*�����0�U���$2���X�*Ⴟ��O������Ϣ�1t��oz���N�>�'�T"��޾� ��a?��aT��+�k��_U���H�זF���N���`�f+}���������<�̾������=��g��{������'V���p���`���Ҍ���l�y�B�3"�(�3/�&9�
E>�"�g��a�������Ũ�"6��a���n�k��0A��u������о|^��T'���L��+�c���P��H�o�I���U��l��,��Ǜ������ܾ���!�%��L�9Uw�5'��jM��"̪����uԚ���*&`��o8����?��%���*�/�M�O�y��撿H���㿫��&��l���R��V�`���7�
i�����&�˾+���N���b���Ek��[���V��[�kk�"?�����R���vLʾ���I���#5��r]�粄�<���맿vҬ�K^��y<�������9U�Y�0�����>�D��F^8��C_�%��O���i���u��q3���ܕ�E�����U���.�>�$���7Ǿ������s��@t��h��Kf�]�n����E ��4~������ݾ���n!�fYE�[o�/���$����i�����[k��ڐ���t���J�>*��%��+��5'�%CF���o�d��7���Yͬ�r���`E���Ǐ���s�dI�1�$��@�85ᾂ���pr���y��1ԁ��_p��<g��mh�L�s����N����੾��ž�~�5Q��b,�R�R���}�_r��~������uV��0��`���hYf�g�>�v�"�v2�H��j0���S��Y�4���Ϊ���b�� ê����눿V�e��<����5��}�վ�j���h���N��ж~���n�_&i��m��|��֊��j��$ȳ�LaҾ�  �  ���d>��&#��!>�(F[�/Mv�'���hp��'X���l�L�L�,�������9�������33��{T�;s�K?������{/��q�6&U�<8�@�`0�4h��QξTm����������{��k��h��s�Gt���0E���¾��޾	�����c\,��`H�}be��h~�h���↿d�~��;c��5B��~"�|�	�Ϗ��$����ND��k>�_�_��{��S������:���8h�jZK�Y/�T9����ږ�<ž�n���h�������ku��j��*l��v{�1K����������;��ێ�����6���S��o��.���s������Hx��aZ� )9�Ha�S;�����	� � �U�+�^uL�	�l�~��1��&5��ú|��Rb�#0E�e�)�g�����f�޾^�þ�z���ј������y�1�x�9�g/���d�����oþ5_޾���0��ڡ(�b�C�Y�`���{�z`��r-��,���kr���R���1�w�� �\���\�uJ�n�9��Z��y�O���R������:�w���[��?���$�g!�q����ܾ��¾)ᬾ�����3��
{���C��E���[C�������׺��@Ӿvg�@F��Z���4��P���m��M���Ɋ�k񊿯Q���Jk�2>J�h�*�����E� �����B'��lF�/�g����)\��~��jJ��p`p�B�S�o=7��r��	��
�1zվ5Ƽ�
���X���c���!����|���֌�N��S(��-%¾R�۾sK��!H�s�#�z=��@Z�ٖv� y������\@��<�~�v�`��c?���!�"F����ǈ����Ll1�lR��er�MÅ�2����Љ�V����g��eJ�g/�_�����=龕ξ�������E��>�����ؓ��K��� ���y���˾v��  �  ���f�6| ���-�:[<���I��6R���R���I���8���!�p
��|�)Ծ��̾%iؾ�^������:'��+=�M�)�S�*Q�s9G��9��9+����K����y���d~ܾ�¾kw������k�b勾X��"����6���:Ѿ�������h�f��bn%��S3�z�A��M��T�n�Q��E�E�1��Z������mkо�UϾ���1g����4/�$�C���P�bT�p�N�j�B�{�4�+�&�"��_�;��dI�W�Ӿ�������d��������]��0���p���w�۾�����2���a�Ed+�J�9�X�G��/R�^�U��7P�,aA��,��v��h��ྕ�Ҿ�%ؾ���~%��v"���9�K�K�rV��{V��N�*�A��d3�^�%�����2���B�v�Ҿ�f���+��𤘾z����!��TG���`����Ѿn��H���f�R����%��l3�O�A��O�ҩW�raX�Y�O��>���'� 8�_?��B྆�ؾ���?� �|��ռ-�K�C�ŶS�ĕZ�h�W�<N��]@�!2�x%�u=�&���P뾱�Ѿ�����x�������꛾�V�����<�Ⱦ�ᾟ����+
�,���E!�[�-�j�;���I�+�U�.\�ݬY���M�d�9��c"��������g��O߾����e	�a��a97�ǍK�+�X�\�,�V�8K���<�<�.�41"�̝���Ⱦ�� ���ʾ�ȴ�2���w`��p�������c���uо��I��Y���K�H%�D2�}C@�h5N���X��j\���V���G��b2�"��\�� 쾨�޾N��c��J��b�'��?��RQ��R[�ݲ[�3�S��F�"�8�++�Y���i�Ϸ�7�����ܾ}Pľ�⯾�&������3��� ���¾�9ھ���8���  �  &���*��W,�vu,�!{,�[^,���*�b�%��Y����Q���r۾�迾�0�����(0��Awž��������W�'���+�k�,�7�,�g�,�u�,��*�B�$���I��`���׾׼�]�����Gk���rʾ���#�2��r!�k�(��>,��-�-��-��,�%*��#�m����	����XҾɛ���Ы�J���i���Ͼ�0����v���"��s)�M,�4�,�4�,���,��,�_
)��!������쾧G;5U���ݪ�����Ig����ԾR����|��n%���+��$.�1�.���.�-�.���-��*�,6"�����{���;;�������ֶ��HnþZ^޾�2��kE�T��W�(�L,.��0��S0�P0�2F0��/�J�*�f$"�n
�������*V̾��kɱ�?����ʾ��� �����8"�q�+�(Q0���1�g�1�F�1���1��90�rP+���!��%�l��8��
�˾�(��7��D���@ҾŎ�������%�FX.��w2�z�3�j�3�2�3��3�!�1�&�+�[�!����G)�M澞o̾���=����ľ5�ھAS��yz��/�sx)��%1�-�4��b5�'V5��V5��4��N2�<�+��� �V�����a⾂�ɾ�ͻ�7��:eǾ�߾14���������*���1��n4�L 5�?�4�� 5�8\4��L1�?%*�e\����yf��$�ݾlƾQ����A��'�ʾN��<�����ov!��E,��o2���4��05�,5�-25��K4��0�|�(��@��v��v����پ�.ľ�����f����ξ��}�t��+�#�x�-�%c3��L5�Z�5�i�5��5��H4�b0��Q'�h(�9
�y��־�r¾������ |Ӿ%��N�����G&��  �  ~�R��Q���H���;�0-�9������q��C��N�Fgƾ�m��+񚾅���񊾏����䞾����XY̾)�f��}<�o����"���0��?�d�K�wOS�%rR���G��P5��.�1!���-GҾQξH�ܾ�9�����tm+�w�@�[O��DT�R0P��ZE�X7�>+)��J�����!�
򾘂ؾn���7��hȖ�; ��!���<9��٥�E,���jվD�ʨ�!"�����f'�&r5�1�C�I�N���S���O��SB�#�-�� ��" ��`߾��ξ2IѾ>��V�IQ��3��qG��#S�I4U�W�N��VB��4��8&�q���_����!��Ӿ�޺�Sɥ�4���S���'q���<��<[��ZCʾ�)�J���A�
��S�?"��w/�`�=��kK�mU�&JW��P���?���)��N�����X�߾^�վO3޾����~��(���>���O�jlX�FLW��[N��A�7�2��J%��N�-���'��F뾠�Ѿ���ֱ��q���&�����:�������lzپ|�H� 	�ʋ���)��7�e�E���R��AZ�{}Y��"O���<��%��������G��J޾�,�e�����3��I�{W�ˣ\��X���M�9�?��j1�x$�:���B�W"�����!ϾA���ʦ��������5���׵��0̾_w���|���<���"��/���=�:�K��/W��/\�aX�L�J��5��Y��N����Y�޾��=�������#��;�:sN���Y�U�[��@U���H�{�:���,�Vp ����\	����uM�ytǾ�'���#���|��/��w�������S@վ����)�z�h��yr'�A�4��C�,�P�7OZ�)�\��2U��D���.�@����+U���޾JQ��� ����X,���B�bT��  �  m��N<��$�t�ŤY�{�<�3�!��0��:�mOҾ�̷�|ᠾ����!#~��l�#�f��/o�=���ԑ�����_����.پ�_���!���'��JC��o`�o�z��х�1P����H6h�1�G�zJ'��4��1���Y��;�������8�$FZ�:�w��~�������灿�l�=�P��3�_��%��l�ʾ�ǰ����0���x��j���i�L3v�`��̧��������ƾ���7����D�0��L���i�������F�6Rz�;�]��W<����Ȟ��W�����85��~$�ȦD���e��a��o���=!���~�ELe��CH�m,��[�]� ��^��ľ@���n��a��|2{�r��ev��ك�"9���;�����X־R�����7�"�qB=��BZ�wv��c��q��ʫ��|~u�U�V��p5�u���q����V7����%�2�ͶS�w|s��l��$������mbz��_�[	B�[G'�I���0���Zݾ#�¾l8���=��YҊ�r��nc�������NǞ�����˾����}�N��b�.��#J�7Jg������J��'׊����R�o��:O�^/�$!�Ψ�K����� #��JA�U�b�w%��n�������^��YNu�O�X��<���"��P�����Iھ�������:��GD���@���؄����_��謨�����־@��G�
�r��x�8��)U�3�q�aք�Z>��	���N����e���D�:�%����;�+�����,�hL��l�i惿���8���7����k���N��3�4����u�B�Ѿm���	��Ĕ���������s݆�8F��6i��R3����ƾ��྅b������(��wB��{_��?{����O��DA��d�z�l�[�f_:�ޡ�:2
�X�������4�6�F�W�<�w��w���  �  ���r���u��O���C�U���-����b徚彾�ӟ�Q㈾�Zo��W�B�H���D��WK�0�[��v�𾍾W0��q1ƾ;�-��"R6���_�ʅ�ի��A󦿆���4����<���Yt���H�i&������b��18�x�`�3����ߚ�˯��ȩ������A��\s��>H�c"�3���ؾ1��,|��熃��h�!�R�XH�3sG�p#Q��d��`�������I���:Ӿz� ��`��rC��$n�2ь�;���[ ��O�������	���%e���;�x�������a�#�\E���o��_��*����C��ޙ���_���	���)f��g<�����a��v0ξ*d���m��.���ph�=�V��P�X�S�u9a���x��f���飾^R��N��$�gk-���T�e8��jI��7B��E���ic������Y�����Z�'v4����L��{C��Q1���V�-����
���զ�����L��3���{��{[��3�	�=Y�r�Ⱦ�����9��]6��w�n�P�`�o]�~Rd�ju�Q>���W���Z�Ӿ$���vg��)=��df��6����Yl���~��qF���򓿸�{���P��d.�n�M��#�_�@���h�,􊿉��k㫿����!�
l����{��~P���*�����Y�P3ľ�����������ys�<h��kg�q��x��ef��װ��dc��b����&���K�bZv�,�����E��lv�������0��qom�:D���%�b����j{+�*�L��{w�����6�����L���!����X��1�l�mC��|��F�ZH۾z]��>��\9���n���Ho�t�g�A�j�Hx�Ψ��[��ମ�o�˾�M��Q�G�2���Y��Ԃ�|痿৿�������+��<��	�_�iK9�Ӵ��+�]����5���Z�᥃�D#��U⨿�  �  ��˿�/Ŀ�G�������p�i'=�O��k��r��-C��|v��[T�26>���1�(w.�(�3��B�2[�w��$A��m(���I�Ԭ��9H�U�}����������Eǿ�i˿������S׎�)]g���<��o#����3/���R��_��Ƴ���@��T�ȿ�˿�����%���zV_�͂.�ە�k�Ծ�ͩ��:��]Ik�ɥM���:�Z1���0�^&9�>�J�gg�|5�����̴ξG���q)��2Y��b���ि�ü��2ʿ_ɿ�s��¡���M��)@W���1��q��!�j9��Hb�c����<���}��5�˿�6ɿ���ϣ���炿&�O���!�����>�ǾEӡ�����3�g�ekN�@`?�R�9�v�<�"�H�1^�������>���O澂����;�r�n��Γ�?r���yĿ<pͿ	�ǿ�괿:���j|��M���-��"�0~+�I�$w��w�������ƿm?ο��ƿj��eԗ��[v�>�B��U�������o��;Z���mk�C�U��I���F�|�L��\�~+u�.��������̾������"�O�&G��@���1��ɾʿ&�ο�Ŀ�x������:o���D��+�_'��`7���Z�����x颿zv����̿�8Ͽ�9ÿ3���叿�g�θ6�t�����)����\��������m���Z�~WQ���P�� Y���j�G���2D��5�����޾"��U�1�H`a�~��  ������5Yο~�Ϳ1���&˥��u���_�c#:�ؚ'���)�o�@��j��y嫿
ÿ!Ͽo�̿�b�� �74���*V���(����վ^ͮ�����iz���9g�K�W��^Q��S�$b_�u�t��u��١���¾u������@���s�Uk��+��$ǿ�
п�Jʿ�t��M���~�����Q�v_2��&�0��M�N�{�5���Oٴ�M�ȿ�  �  t3�)�ۿ2CĿ~k������j�I�]#��|辘'��ƍ�kOh��+F���0��$�0�!�\�&���4���L�1�r��J���彾x��3#���V��j�����̤ʿ�(߿V�R�׿S���4���s�|���K�}k/��*�J�<���d��J�������Ϳ@����,�տ]����r��iq�3�8��#���վ2������8]�+�?��q-��$��$�8�+���<���X�\큾1���I@Ͼ���	3��Qj������඿��ҿR����Eп{o��D���fj���?�#�*�b�-�Q�G�N�v��P��1 ���ֿ$��L῎^οF�������F�^��#*��m��>ǾU)���.��
Y�!�@��C2���,���/��;��P�.q�a��M|����込9�դG��O��;����¿C�ۿ	�gi߿�ɿ����{9���)^��o:�oI-���7���Y�:#��I��5�ƿAD޿`�濴O޿� ǿ�(������@PO���&t�94���򘾹�~�]>]��"H��<��J:���?��MN���f�����d���Xk˾���k*�Eu]�UՍ��y��ο��⿖��Ahۿ���↡�w^���T���7�h2��D��dm�r���h;��!�ѿ��7��ۯٿƶ��"���©y�MA��O�� ��c���?���b}�I�_�(yM���D��D���K�t�\���x�Z��������h߾��~.;�6r�ݥ��n ��a ׿���忧oԿ0����ؖ���r� H�W3���5���O���~���������ٿ4����C�ѿ峿�I��se�Q�0�D��VԾ�#��� ���r��aY���J���D��G�z�Q�p^f�ԇ��O!�����}�8p�v�L�}ꃿ~4��ſ�3޿ڮ�F��I̿�������j�b��.?���1�ۖ<�4^��Z��`s���ɿ�S��  �  dF��y��&��&c��8�wr���L���3B�� �U�1�/��.��;��H�������F���c	��X��M7��`�H4��������P��|B�O�l����[���B���򐿿o��_e[�GV4����h�b���q	�].%���I�9�q��슿�J��U��Ț��ގ~���U�0�+�t3���ξ�����!z��>I���'�����h��������?����|�$�@vD��Ms�욾n�Ⱦ�8�w'�9�P��y������i���ؖ�.r���v���M�2�(��4�g��%a����V�0��W����%��1�����X���V�r���H�&! �g������ ����n�}�C��'���;H
��u�"��*�k� ���9��o^�����H3�����8��8��Cb� ���듿�5��=�������l�U�D�'("���
��d��v	��S�
�@�d�h�1����ʕ�z����֕��ˇ���h��G>����N��o����R����k��2F��@-�e��M��{������"�175���Q��p{�)���žGA���� ��LI��s�;r���Ҙ��ɛ�Ѝ��"����b�O<����Bt
�d��@��r-���Q��Az�k��rs���*��W����h����]�'�3�[��߾�ϯ��+���Xi�5�G���1�AK$����"]�f#���/��|D��kd�����P�����ؾ�O
��1/�8�X����@��L�����������J~� V���0�iU����tT	�	e��~8��	_��u����������P���ꎿ!�y���O�V�&�|C�	�;a$��B��[]��8@��l-���"�`8�>����'�y#7��lO���s�~��������l��A=��xg�E���Q���=͜�DΘ�����ɦq��I�O�&���_�c�J�#�fE�ALm��ډ��ۗ��  �  ����2���π��c\��4�^s��pݾ����H�����W�"�2��y�eu	�� �����nA����;���<:���b�~A��(����X���R=�Q�e�B����U��S��H"��Z�z�q�T�}{/��o�����T��Q���� �N�C�|j�?d���:���ޒ�+݊��v��O���'����|y̾���f{�}�K��+�� ������ �]� ��h����'�(G���t������lƾh����##�$�J�	Dr��N���J������Dև��in�+�G�C$���	�||�������(,�KQ�$�w�ee���y���⑿h���k���C����`�����
��"�p���F��Y*����Bj�Ҁ	�?��[_�Q$��<�,�`�RL��yN���޾�e���3���[��ဿ�����9B��}�����e��@?��.�����P���v��{�e�;��b��u��ݐ�̕�fꐿ�����a���9�����_��������<"n��@I�'�0��� � �����0�K&�F|8�g�T�Cg}������þf�������"D�
el�����͓�Ƞ������6���}\�O<7��X����WM�5�3)�I&L���r������c�������$�~���W���/�,��7�ܾ�C��΍�,�k�9K�{5��x'�K� ��j �?&���2���G�Og��f��֚��ދ־c���B+��R�(rz��h��bg���ޕ����v�EP�p,������W{����9�3��X��~�V쎿Gꖿ�A���f��6r�*J�e'#��@�(+̾V���)���7`��{C��0�]�%��C!��#�'+�o:�i�R��Vv��锾и��)��@�8�a��|�����e����ӓ��H��]�j��*D�'#�L���U������s5@��mf�����풿�  �  ���G̀�U�j��TJ�b_'�8��ٳվ*���7{��U�_�7�<� $�����a
���������-))��"D�GFj��z��c���ᾦ���r/�YSR�Hq�V���7	����}�}d�c�B��!�^O����� �����O�3���U���s��h��݄��{��a�P?��������ƾ���G�����T�cm5�������
��
��M��p��F2��}P�b�z�������������Q';�3M]�\9y�PY���ك��lv�s]Y��7�d�۞ ����`�F���k�?�S�a�G�|�is��C���u�V�W��5��5�t9뾮u���▾��w��tP���4��H"��3�,��_��n��.�)�F��Vi������謾�׾��nc'�2WJ��*k�Sρ�����n�����q��R�GX0���g���R����e��G_-��&O�go�$e������4�����o���O���,���������e���&Yv�jS��;��+��U"��U �H�$��G0��C��c^��o��BꜾ�����5�q���C6��'Y���w��#�����E���:vk��J���)��1��������,���T��B<��@^��?|�T������N��P\i���G���$��x�L&׾�ծ������u�?oU�m�?��k1�*\*���)��#0��K=��+R�Orp�x��y���o�Ѿv��� ��MC��ze�����qu������~�E�a���?�h0 ����������X���&��XG�
�h��끿�∿�{���B|��b^���;����AZ���ȾD棾}���c�i��N���:�mr/�B�*���,��85��D���\��~��%��$k��|-�B�l�,��O��ap�j������e9��D�v��W��C5����-
��6��̙��9���1��uS�9�s��t���  �  �c�7�\�� K�2�z������"ξ㢪�_Ȏ��Lr���P���7�$�%���u��i_���)��&=�1X���{�Yє�5R���׾���"�Q8�.P�(�_�91c�*EY� dD��)����^�־{�Ѿ�������E���8�q8Q�ۄ`��!c���X���C���)��v��뾭�¾�������?h���I�B�2�@s#��q����"�џ0�9F�?d�vN���3������J��U�ZE&���@��tV��Lb��2a��1S��;��% �NU����ҾEfվ���G�a.'���B�`�X��d��Xb�QT�s�<���!��h��"�๾N����A��8dd�;�H��'5���(���#�Eq&�K�0��8B��"[��|�_B�������CѾ�h��A����2�bL�gG_�{g�s�a�P�O�u}6�X������"�X�ؾZ������wG4��rN��_a�Ʉh�CBb�wP�zz7��4���fپl���<ؙ��U��2�g�;�N�q=�P}3�H1�3D6���B�w�V��jr�=$��%?��zٿ��U�L�	���#�o&?�DW�@�f�;j�s`�h�K�f
1�N0��_ �B����ᾠ<�N"�)�%��>A���Y��h�0nk�^�`��L�D�1���v�����ҾZױ�����+��!�i��R��TC�kJ;���:���A�MzP��cf�����QR��D���<ξ�w��.t�k.�dI�k�^���j�^ki��i[���C��S(��w��-��"�⾱&��\��y��1�.��I�e�_���j�.i�j�Z���C��(�^��D��ƾ����&���}�Vb�*�M���@��;�ݸ=��oG���X�"q�Ɉ��᝾�����۾�h�����8�z�Q�t}d��Bl���f��U��;�z��L�����TR�F���@�k�8�g�R��|e��  �  8�9�V96�Z�*�Q���U�����'; P���P���@��Zhs�X�W�t{B�{5�x�1���7��F��]���z������[���0���Ծ��.��,�%.��C8�<�9���1�z�!��5���k�ξGd��ˉ����þ<�����@��+���7�zL:�-�3�a�%��A�m���%�"0žԵ�������}���~k���Q���>��4�YL4�0G=�gO��
h�cm���X��4奄���SJ޾�n�������#�@:2���9� 8��-�@����X�sƾl��s����̾���!��f� ���1��:��n:��71�S�!����3��-۾"ſ�Į��~Ԕ�i���L�i��R��ZC���<��+@�
�L�8�a�}b}�8��68���	��
�Ѿ����$	������,��69���=��9��j+����S������pǾy����ž�#޾iS�����*�,9�K6?���;�Q�/��7�������&ؾ6J���`���o�����J�n��Y��fM��-J���P�9(`�ڄw����2曾Ư��ƾ=�᾿� ������$�)�4�q2?���@�'�8�{)�Z��a �؈޾�Bʾ,�ƾK8Ծ4����(P!�,�3�
�?���B��<��0.��z�b
�,s�fkվ�߼�Q֧����������q�R�^��T�, T��]���n�����f���[��d���Ҿv����Z�V,��j:�S�A��B@�HF5�H#��.�������־�NǾ�Dɾ�ܾ]������n�'�׌8�ЛA��)A��7�df(��/��-�5��̾���G����U��e���+zk�i�[�H�T�5vW�4�c�4x� ������٬�&�¾��۾���6Y��� �o�1��l>��C�->�΁0�"�S���t���о�ZǾ�Ͼ�������.��E=��  �  ������K��������龊8پ��Ⱦ����D������-��0�j�~=Y��%T�$J\��}p�����e��W����c��s;Kkݾ>^C ��o	��7����������R��I�H�žq�������V���ݢ���ʹ���־��������Q��{���g���������`�F�Ծ%�ľ�U���7���:��,~�.}e���W�o�V�LBc���z�+��@ ��"���l¾E�Ҿ �^c���^��?�h�������K�	�u�����پp���꒦�~���1��[r���þ0���� �>��ty��@���������Q��U�Ҿ}C¾�հ��˞�qn���,}�eZh��]_���c��vt�
ԇ��ɘ�@(���R��-}ξ)�޾юﾫ� ���	�kb�S������x	�v���)׾��3D���W���Q���C��"8վax��7	��o��8�T��������aQ�&���7&�`�Ӿ-.þ=t���t�������#���#q��~l��u��߄��ϓ�ot��K跾u�ɾ�ھ��꾦�����FG�>��w�����9��-��Ծ?���N��`����Ӵ��!ʾ��Z%���8��K��(����~�����P���~/�ܻԾ�nþ�B��:����k����w�X�v�Պ��.Q��'������1!���zҾ���?J�%N�b���i��C�(����	���V ��̾A���qG������Z�����Ҿ��p������N�����3�̺��	��� ���\�߾�AϾ|���D�������=銾H��+!w�6�z� ���[��5ǣ����Z�Ǿ&پ�X�T������u#�ș��O�d@�.<����� �H�Ϡž�Ʋ�Ш���o���-þm�ݾ����H�׆��  �  �$��l��gZ�����N��ja��<W������u⾖�Ͼ�"�������������;���䢓����ω��i|Ծ�c澑|�>���[O�������������7+����Zྼ�̾����7ܟ�/ڍ�;낾Sހ�����C�������¾gؾ�e�wx���������Z���1���������(�:�ݾUQɾew������ϴ���������-���x���ʯ���ƾwy۾�v��x���:��������e������������t�&$ھU&ž�W���S��卉�����D��K��9���9���`̾���iF𾙗������;+��,a���
��z
��K��8쾈�ھ2~ž�Ԯ�W���������=j�����%����4��F	Ծ���p����=���� �_��i��%������4�����F�ھ�ž_�����������������
������Xľ��ھv������*�Ť�� �O�P��
"�������2�ھ;|ľE5���}��Ao����������9��|���]�˾3��>��@���<��v����y��YH����7���	���&۾�ľJ���rC��N����Ȑ��(������[l��3nӾ=��{���͂��J��<��c�,G����ee�EP�����P[پ!v¾��������
���~��2���d�������־Uz�#���v��a1�I����
����T������@y��lվ<����b���r���U��.e��Ft���ڭ�a�þ �ھ�������E�����2��G�4����-�������羇-Ҿ%U��٦�N��us�����兟�%豾8Ⱦ)�޾d��@ ��X�p���d��
]���"��(;��O��Ͼ4d���������Y���8(����4��H�̾�+�"����  �  N�ɾ1�پ?�꾤�����������������QJ�'���ɾn���󗞾�����}�������о
�g������1T�rq�����b��}��n;׾B�ƾ�赾�죾ב��I��	qh��X���U��&`�gv��W������C��iϿ��cо)������d��u�q���������0���[߾�[��詩��Z�����/���6;����۾���˨
�SC�������������7T�⾖�ѾVA��k䯾Sɝ�r��3;y�ޕb��oW��uY��nh��"��tÑ�� �������Ǿ0�ؾ#'龮���ī��f����͝�����	�������ؾS����W���T��D+���F���;��H1��G������J��j�{?�Rs��Ƣ�]qӾ5�¾n5��A(�����f����l�h�e��#l�D�~�^�������{����þ}Ծ��侗��������1�!?�TD��I�����0���{վ3c�����A����ҭ������ݾ������|�FD����>�����~����5�Ծyľ�c��ѕ��VS��h�����w�'�u����nA�����(v��þ�pVоh���6�G&�QE
��K�!������
����Y�9QѾ����	E�������w��&ξ(�뾺X�����H����������^�
�����b�"�J�Ѿ�.������7���������m�v�%x��F���㏾�3��OB��h^ľ��վ���t����YB�����I��"��!��P�KH��c�5�Ⱦl���5��i׮� ����EؾP���Y�
���W�7��~�����t����� ���ݾ�;k��M9��s������l��Sx�K~��R��le��Ʉ��9Ĺ��˾�  �  �a����ξ�n�U�P���b+���6�>�9��c3�$��k�����Ӿ���P���Lھ3 ��C�B�(�(�5��<:��#5�<X(�@�#����澰@ɾ����������D�o���T�DA�8�5��j3�w�:�DgK�apc�y����P��~���齾��پK����F!��0��b9��O9�a�/����b�	�����ʾr���-���J�Ǿ_�� ^�ye�4.��8�ְ9�O�1���"�����o���wܾPN��j������zZ��\f�r�M�f=�E�4���6�M�A�ƐU��_p��b������t���\ɾ0��
c�����g(�g�5��<�9�8��,���r��z�]_Ǿ�!���3��q�վ�����V�_�%��5�3C=�SH;���0�4� ��?�����{�پ��������(���V��8Ol�QV��EH��lC�C;H��NV��tl������v���⨾�=��uپ	^�����; �"�0�M6<��W?�%�8��*�%�/���޾K�Ǿ�j���9̾,���e����/�=|<���@�$�;��"/������������׾���(ר��o��K�����r���_���T��R�&�Z���k�|���"���Ƣ�G����lξ���=�P��r)���8�_}A�6bA���7���&����y���=�ھp�Ⱦ�ǾO�׾����[U�%`$�Q6���@��A�3�9��+��������쾾�о{θ�nW��Y���w>����m��{\��T��!U�5�_�s�r�ˎ���v���ߨ�3����־�	��0�
��c���.�sv<���B��J?���2�c! �@�
�oC�oӾ�Ǿ��˾�W�������M+���:�4�B�M�@���5���%��t�Ű�5�/rɾ_ᲾW_���h����2�i�YE[��U��ZZ�	�g�׷}�x���2�������  �  �#���+о����r:���3�uHL��]��5c�?p[�H�Z�-�ho�$�����ؾ�Nо��ݾ"����o�x4�n^M�6�^�B]c�g�Z�đG�w�-���E��ZȾn5��|���m��M��5�?
%����;�G) �Е-�YB���^��ށ�	ϙ����DY߾XD��!�u�<�{�S�}|a�B�b�6�V��W@�]%��
�J�뾚uԾ>2Ӿy������!��\=��wT���a��b�h�U���?�>�$�9�	����L����z��������a�E���/��"�����B��A&�X�6���N�K,n�ʋ��4Υ�PHǾ��&j��,���F�"[��e���a���Q��i9����������7־g�ܾ�i������-��H�8T]��f��b�nuR�JR:�P����L�ܾ\��������I��� f��K��?9�T.�-V*�p8.��9�UiL��f��q��򗚾� ��۾���Q��C�8�ƻQ��c���h�e�`�)�M�i�3��6��0�p��EbܾD,�o'�D���:�(�S�e�~j�4�a��XN���4�x�jT �l/־A/������!#��M�j�`xS��jC���:�˟9���?���M���b�=b�M��!I��ɾH�ﾕ}��$*��E���[�E�i���j�2�^�[H��-��y�	s��)_侼��������)��VE�v\���i��)j�1�]�,�G���,��� ��UH̾�����(������e�ėO�nA�]�:�%�;��D�@�S�m-k�p��T���_����Ծ+^�����13��QM��a��k�W-h�KHX�
�?�$���
�z��KV�����Z�'�3�GEN��b���k���g���W�?��R$�"-
����x¾e�������%z�x�_���L��A���<��Q@��IK���]�gw�沌������  �  ����@Mؾ�D��F)�WDL�x'l�rK������W����h�[H�(�&���
�֦�T8�%����U��!.��P�*<o�v4��!��+�}�e���D�j"�1���Jξ�8�������Z�`R9�2"�P��_�
�Mk	����¤�A9.�s�J�9s�pG��b���)�qs�Њ5��$X���u�:�p����z��_��r=�������d�����:��k�9��d[�=�w��3��b5��8x�X�[��<9����s�����c�����w�/`N��0�s���}�z�f��^��g#��Y:�m[��=��2%���2̾\\ �����B�Kmd���~��܅������at�QV��74����( ��8� ���Q1�v&���G���h����ņ������s��S��1�ˠ�#��X��D*����v���Q�4�7���&����r����3'��8��bR�]�v�Ɔ��4���9�¼���.�׸Q���q�F��·�g��+^n��N��,�2�������F� ��܇��k4��qV���u��~��hi��1߂��l�i�K���(����`ܾ�/������ \w�[�V���?��11�}�)��(��T.���:�}�N��zk����������˾D��������=�O`�f�}��·�ֹ���R��6g�~pE�n%�h��H����p����	�۽!�"�A��^c�=��5�� :�����ѭc�GYA����L� ��:Ͼ-ͨ�h%��e�n�g�P��}<�i�/�2�)�H�*��2���@�O�V��w�R ��g�����پ{����&��^I�!�j�X���s���-���z��V\�d:�n��c+����/N ����B!,��_M��Kn�#ƃ��j��ә��];x��Y�-76����AG�;j¾�{�������	f���K�:��/��,��/���8�G�I��5c�ۣ��N����  �  �ӭ��lྨY�=E6���^������Î�v'��Ծ�����[��5��]��3�8���D��Ӡ��F=���c�����ޏ��&���DO|�-V�2�-�V	�/�Ծ�]���(��2�Q��/��������;�9������R�A�#�&0A�Cl�,���|��ġ���hND�Bl��+������|����7����t���N���)�@��f���P��P0��<&��;J���p������$����	���5Gp��H��!��-����þ'U��ώq�M�D���&��������v���s
�d �'0��!R�
���"ѣ�0Ҿ����E+�9`S�6;z��\���擿��������`j���C�Ou!��	��������sw�[14�<�Y����V���ٔ�S���o����f�̖>��7�}�ĺ����:o���G�^g-��l����H�4\���.��JH�I�n�0ǒ�y���&Y����P�;�'d�@{��k~��f敿˄��Ղ��`�V�:��<�E&�;^�m�
���!���C�N.j�K��%���x��V�������\��4����4��lR��0K����n��1L�YL5��'�����*��w$�{a0��D�g�a�2���Y����ξ��rM%��L��kt��<��Ѡ������U<����|�v�V�W�1�Ҙ�������#�U1.�H2R�H�x�u���D&��s"������]x�ѵP�))�\9���Ӿ����Z�[#e��hF�2���%��b ��!�G(��6���L��n�T���[���}߾ȟ���1���Y�Na��>���� ���
�����p��J�M�'�g��O�����<���9�ʎ_�捂����9���3���	��il���C��m��1��T'žQ���Ӂ��\�x4A�L�/���%��"��n%��.�	J?�Y�U<��㚾�  �  � ����㾓o�];�bhe�w�������R��襒�jC����a�F#:��&��,��+��=��Ī�u�B���j�_"��qޔ��P��u����D��?k\�LL2����S�׾b+��⮁� �O�.�+�L�ȩ�VQ������)��y�t �m]>���j��ʔ�I������V� ���I���s�5���P����ԗ�le�|���T�W�.�w�W� ��������y�*��<P��sx�K[���@���9��'D��f�w��MN���$�MU ���ž落�gp��?B�(J#�KF�n���D��*����H�۹�p�,�0�O�
��5s��
�ԾV�	�_�/�q�Y�+"��z#�����̖�a����q��I��%��K�!�D���!�L 9��`������.��@�������҉�I�m�˥C��{�k[�$��ä���/m�I�D�{*��-����i�D�L����*��DE�B�l�숒��߹�������@��j� Ȉ��q�����l�������g�u�?���.
���`��s�%���H��Uq�]��I%������;ܔ�����(4c�9�����|�F��;Џ�3l��I���1��#������!O!��-���@���^�⧅��;���о
"�}�(���Q�g�{��ʏ�k����ܛ��󒿦h����\���6������i����2�3X��6��Z��2B��>���K��	��XiV���,�ww���վ&ਾ�-��!fb�k.C��.�)�"��U��
�m�$�|�2�_[I��k�꾎����� ��0��6�`�he��xb��3G��"����,����w�ħO���+�M����r�����>�~"f�����ߕ�'���h3���m��s���H��� �s���Y�ƾ2����΀�]Y�}�=���,�-�"�j���U"�Kr+���;�%V��}�M����  �  �ӭ��lྨY�=E6���^������Î�v'��Ծ�����[��5��]��3�8���D��Ӡ��F=���c�����ޏ��&���DO|�-V�2�-�V	�/�Ծ�]���(��2�Q��/��������;�9������R�A�#�&0A�Cl�,���|��ġ���hND�Bl��+������|����7����t���N���)�@��f���P��P0��<&��;J���p������$����	���5Gp��H��!��-����þ'U��ώq�L�D���&��������t���s
�b �$0��!R���� ѣ�.Ҿ����E+�8`S�4;z��\���擿��������`j���C�Nu!��	��������sw�[14�=�Y����V���ٔ�T���o����f�Ζ>��7��ĺ����:o���G�`g-��l����H�3\���.��JH�F�n�.ǒ�w���$Y����N�;�&d�?{��j~��f敿ʄ��Ղ��`�V�:��<�E&�;^�n�
���!���C�O.j�K��%���x��W�������\��4����6��oR��2K����n��1L�\L5��'�����*��w$�{a0��D�g�a�3���Y����ξ��rM%��L��kt��<��Ѡ������U<����|�v�V�W�1�Ҙ�������#�U1.�H2R�H�x�u���D&��s"������]x�ѵP�))�\9���Ӿ����Z�[#e��hF�2���%��b ��!�G(��6���L��n�T���[���}߾ȟ���1���Y�Na��>���� ���
�����p��J�M�'�g��O�����<���9�ʎ_�捂����9���3���	��il���C��m��1��T'žQ���Ӂ��\�x4A�L�/���%��"��n%��.�	J?�Y�U<��㚾�  �  ����@Mؾ�D��F)�WDL�x'l�rK������W����h�[H�(�&���
�֦�T8�%����U��!.��P�*<o�v4��!��+�}�e���D�j"�1���Jξ�8�������Z�`R9�2"�P��_�
�Mk	����¤�A9.�s�J�9s�pG��b���)�qs�Њ5��$X���u�:�p����z��_��r=�������d�����:��k�9��d[�=�w��3��b5��8x�X�[��<9����s�����c�����w�/`N��0�r���}�x�f��^��g#��Y:�g[��=��.%���2̾Y\ �����B�Hmd���~��܅������at�OV��74����( ��8� ���Q1�v&���G���h����ņ������s��S��1�͠�(��\��H*����v���Q�7�7���&����r����3'��8��bR�W�v���/����8㾿����.�ԸQ���q�D��~·�f��)^n��N��,�1�������F�!��݇��k4��qV���u��~��ii��3߂��l�l�K���(����dܾ�/������&\w�`�V���?��11���)��(��T.���:�~�N��zk����������˾D��������=�O`�f�}��·�ֹ���R��6g�~pE�n%�h��H����p����	�۽!�"�A��^c�=��5�� :�����ѭc�GYA����L� ��:Ͼ-ͨ�h%��e�n�g�P��}<�i�/�2�)�H�*��2���@�O�V��w�R ��g�����پ{����&��^I�!�j�X���s���-���z��V\�d:�n��c+����/N ����B!,��_M��Kn�#ƃ��j��ә��];x��Y�-76����AG�;j¾�{�������	f���K�:��/��,��/���8�G�I��5c�ۣ��N����  �  �#���+о����r:���3�uHL��]��5c�?p[�H�Z�-�ho�$�����ؾ�Nо��ݾ"����o�x4�n^M�6�^�B]c�g�Z�đG�w�-���E��ZȾn5��|���m��M��5�?
%����;�G) �Е-�YB���^��ށ�	ϙ����DY߾XD��!�u�<�{�S�}|a�B�b�6�V��W@�]%��
�J�뾚uԾ>2Ӿy������!��\=��wT���a��b�h�U���?�>�$�9�	����L����z��������a�E���/��"�����B��A&�R�6���N�C,n�ŋ��/Υ�IHǾ��"j���,���F�"[��e���a��Q��i9����������7־h�ܾ�i��	����-��H�;T]��f���b�quR�NR:�T���S�ܾb�������J��� f��K��?9�V.�-V*�n8.��9�PiL��f��q��헚�� ��۾���M��?�8�ûQ��c���h�b�`�'�M�g�3��6��0�o��EbܾE,�o'�E���:�*�S�e��j�8�a��XN���4�x�mT �r/־G/������%#��U�j�fxS��jC���:�Ο9���?���M���b�=b�M��!I��ɾH�ﾔ}��$*��E���[�E�i���j�2�^�[H��-��y�	s��)_侼��������)��VE�v\���i��)j�1�]�,�G���,��� ��UH̾�����(������e�ėO�nA�]�:�%�;��D�@�S�m-k�p��T���_����Ծ+^�����13��QM��a��k�W-h�KHX�
�?�$���
�z��KV�����Z�'�3�GEN��b���k���g���W�?��R$�"-
����x¾e�������%z�x�_���L��A���<��Q@��IK���]�gw�沌������  �  �a����ξ�n�U�P���b+���6�>�9��c3�$��k�����Ӿ���P���Lھ3 ��C�B�(�(�5��<:��#5�<X(�@�#����澰@ɾ����������D�o���T�DA�8�5��j3�w�:�DgK�apc�y����P��~���齾��پK����F!��0��b9��O9�a�/����b�	�����ʾr���-���J�Ǿ_�� ^�ye�4.��8�ְ9�O�1���"�����o���wܾPN��i������yZ��\f�p�M�d=�B�4���6�G�A���U��_p��b������t���\ɾ(��c�����g(�c�5��<�5�8��,���p��w�[_Ǿ�!���3��s�վ�����V�b�%��5�6C=�WH;���0�8� ��?�������پ��������(���V��?Ol�QV��EH��lC�A;H��NV��tl������v���⨾�=���tپ^�����; ��0�I6<��W?�!�8��*�#�	/���޾I�Ǿ�j���9̾.���e����/�A|<���@�(�;��"/������������׾���.ר��o��O�����r���_���T��R�(�Z���k�}���"���Ƣ�G����lξ���=�P��r)���8�_}A�6bA���7���&����y���=�ھp�Ⱦ�ǾO�׾����[U�%`$�Q6���@��A�3�9��+��������쾾�о{θ�nW��Y���w>����m��{\��T��!U�5�_�s�r�ˎ���v���ߨ�3����־�	��0�
��c���.�sv<���B��J?���2�c! �@�
�oC�oӾ�Ǿ��˾�W�������M+���:�4�B�M�@���5���%��t�Ű�5�/rɾ_ᲾW_���h����2�i�YE[��U��ZZ�	�g�׷}�x���2�������  �  N�ɾ1�پ?�꾤�����������������QJ�'���ɾn���󗞾�����}�������о
�g������1T�rq�����b��}��n;׾B�ƾ�赾�죾ב��I��	qh��X���U��&`�gv��W������C��iϿ��cо)������d��u�q���������0���[߾�[��詩��Z�����/���6;����۾���˨
�SC�������������7T�⾖�ѾVA��j䯾Sɝ�q��1;y�ەb��oW��uY��nh��"��oÑ�� ��ل���Ǿ(�ؾ'龤�������f����ɝ�����	�������ؾP����W���T��E+���F���;
��K1��G������!J��j��?�\s��Т�fqӾ<�¾t5��F(�����k����l�i�e��#l�?�~�[�������{����þ}Ծ��侍������	��1�?�PD��I�����0���{վ0c�����A����ҭ������ݾ������|�JD����>���!��"~����=�Ծ�ľ�c��֕��ZS��l�����w�+�u����oA������)v��þ�pVоh���6�G&�QE
��K�!������
����Y�8QѾ����E�������w��&ξ(�뾺X�����H����������^�
�����b�"�J�Ѿ�.������7���������m�v�%x��F���㏾�3��OB��h^ľ��վ���t����YB�����I��"��!��P�KH��c�5�Ⱦl���5��i׮� ����EؾP���Y�
���W�7��~�����t����� ���ݾ�;k��M9��s������l��Sx�K~��R��le��Ʉ��9Ĺ��˾�  �  �$��l��gZ�����N��ja��<W������u⾖�Ͼ�"�������������;���䢓����ω��i|Ծ�c澑|�>���[O�������������7+����Zྼ�̾����7ܟ�/ڍ�;낾Sހ�����C�������¾gؾ�e�wx���������Z���1���������(�:�ݾUQɾew������ϴ���������-���x���ʯ���ƾwy۾�v��x���:��������e������������t�&$ھU&ž�W���S��㍉�����A��K��5���9��z`̾���aF𾏗������1+��"a���
��q
��K��0쾁�ھ-~ž�Ԯ�T���������>j�����(����4��L	Ծ��x���>���� �_��i� &������4�����M�ھ�žc�����������������
������Xľ��ھn������*����� �J�K��"�����م�,�ھ6|ľA5���}��@o����������9������b�˾9��E��I���<��v������^H����@������&۾�ľN���vC��Q����Ȑ��(������[l��3nӾ>��{���͂��J��<��c�,G����ee�EP�����P[پ!v¾��������
���~��2���d�������־Uz�#���v��a1�I����
����T������@y��lվ<����b���r���U��.e��Ft���ڭ�a�þ �ھ�������E�����2��G�4����-�������羇-Ҿ%U��٦�N��us�����兟�%豾8Ⱦ)�޾d��@ ��X�p���d��
]���"��(;��O��Ͼ4d���������Y���8(����4��H�̾�+�"����  �  ������K��������龊8پ��Ⱦ����D������-��0�j�~=Y��%T�$J\��}p�����e��W����c��s;Kkݾ>^C ��o	��7����������R��I�H�žq�������V���ݢ���ʹ���־��������Q��{���g���������`�F�Ծ%�ľ�U���7���:��,~�.}e���W�o�V�MBc���z�+��@ ��"���l¾E�Ҿ �^c���^��?�h�������K�	�u�����پo���蒦�~���1��Xr���þ+�⾽� �:��py��@���������H��M�ҾuC¾�հ��˞�mn���,}�bZh��]_��c��vt�ԇ��ɘ�E(��S��5}ξ2�޾ێﾱ� ���	�pb�W������x	�{��*׾��5D���W���Q���C��8վ\x��4	��o��8�O��������\Q����.&�X�Ӿ%.þ7t���t�������#���#q��~l��u��߄��ϓ�tt��Q跾}�ɾ#�ھ��꾰�����KG�C��w�����<��-��Ծ?���N��b����Ӵ��!ʾ��Z%���8��K��(����~�����O���~/�ܻԾ�nþ�B��:����k����w�X�v�Պ��.Q��'������1!���zҾ���?J�%N�b���i��C�(����	���V ��̾A���qG������Z�����Ҿ��p������N�����3�̺��	��� ���\�߾�AϾ|���D�������=銾H��+!w�6�z� ���[��5ǣ����Z�Ǿ&پ�X�T������u#�ș��O�d@�.<����� �H�Ϡž�Ʋ�Ш���o���-þm�ݾ����H�׆��  �  8�9�V96�Z�*�Q���U�����'; P���P���@��Zhs�X�W�t{B�{5�x�1���7��F��]���z������[���0���Ծ��.��,�%.��C8�<�9���1�z�!��5���k�ξGd��ˉ����þ<�����@��+���7�zL:�-�3�a�%��A�m���%�"0žԵ�������}���~k���Q���>��4�YL4�0G=�gO��
h�cm���X��4奄���SJ޾�n�������#�@:2���9� 8��-�@����X�sƾl��p����̾�����c� ��1��:��n:��71�N�!����3��$۾ſ�����yԔ�d���E�i�
�R��ZC���<��+@��L�>�a��b}�$8��<8���	���Ѿ����$	������,��69��=��9��j+����U������pǾy����ž�#޾hS�����*�,9�G6?���;�L�/��7�������ؾ/J��`���o�����D�n��Y��fM��-J���P�=(`��w����8曾 Ư���ƾE��ĳ ������$�.�4�v2?���@�*�8�~)�\��c �ۈ޾�Bʾ.�ƾM8Ծ5����(P!�,�3�
�?���B��<��0.��z�b
�,s�fkվ�߼�Q֧����������q�R�^��T�, T��]���n�����f���[��d���Ҿv����Z�V,��j:�S�A��B@�HF5�H#��.�������־�NǾ�Dɾ�ܾ]������n�'�׌8�ЛA��)A��7�df(��/��-�5��̾���G����U��e���+zk�i�[�H�T�5vW�4�c�4x� ������٬�&�¾��۾���6Y��� �o�1��l>��C�->�΁0�"�S���t���о�ZǾ�Ͼ�������.��E=��  �  �c�7�\�� K�2�z������"ξ㢪�_Ȏ��Lr���P���7�$�%���u��i_���)��&=�1X���{�Yє�5R���׾���"�Q8�.P�(�_�91c�*EY� dD��)����^�־{�Ѿ�������E���8�q8Q�ۄ`��!c���X���C���)��v��뾭�¾�������?h���I�B�2�@s#��q����"�џ0�9F�@d�vN���3������J��U�ZE&���@��tV��Lb��2a��1S��;��% �MU����ҾCfվ���G�_.'���B�]�X��d��Xb�MT�o�<���!��h�{"�๾H����A��1dd�5�H��'5���(���#�Gq&�N�0��8B��"[��|�dB�������CѾ�h��D����2�"bL�kG_�~g�v�a�S�O�w}6�Y������"�X�ؾY������uG4��rN��_a�Ƅh�@Bb�wP�vz7��4���`پf���7ؙ��U��+�g�6�N�q=�N}3�H1�5D6���B�|�V��jr�A$��*?���ٿ��U�P�	���#�s&?�HW�D�f�;j�
s`�k�K�h
1�P0��_ �D����ᾡ<�N"�)�%��>A���Y��h�0nk�^�`��L�D�1���v�����ҾZױ�����+��!�i��R��TC�kJ;���:���A�MzP��cf�����QR��D���<ξ�w��.t�k.�dI�k�^���j�^ki��i[���C��S(��w��-��"�⾱&��\��y��1�.��I�e�_���j�.i�j�Z���C��(�^��D��ƾ����&���}�Vb�*�M���@��;�ݸ=��oG���X�"q�Ɉ��᝾�����۾�h�����8�z�Q�t}d��Bl���f��U��;�z��L�����TR�F���@�k�8�g�R��|e��  �  ���G̀�U�j��TJ�b_'�8��ٳվ*���7{��U�_�7�<� $�����a
���������-))��"D�GFj��z��c���ᾦ���r/�YSR�Hq�V���7	����}�}d�c�B��!�^O����� �����O�3���U���s��h��݄��{��a�P?��������ƾ���G�����T�cm5�������
��
��M��p��F2��}P�b�z�������������Q';�3M]�\9y�PY���ك��lv�s]Y��7�d�ڞ ����^�F���i�?�Q�a�E�|�gs��A���u�T�W��5��5�o9뾪u���▾z�w��tP���4��H"��3�,��_��n��.�-�F��Vi�����鬾�׾��pc'�5WJ��*k�Uρ�����o�����q��R�HX0���g���R����e��F_-��&O�go�#e������3�����o���O���,���������b��� Yv�jS��;��+��U"��U �J�$��G0��C��c^��o��EꜾ�����5�s���C6��'Y���w��#�����F���<vk��J���)��1��������,���T��B<��@^��?|�T������N��P\i���G���$��x�L&׾�ծ������u�?oU�m�?��k1�*\*���)��#0��K=��+R�Orp�x��y���o�Ѿv��� ��MC��ze�����qu������~�E�a���?�h0 ����������X���&��XG�
�h��끿�∿�{���B|��b^���;����AZ���ȾD棾}���c�i��N���:�mr/�B�*���,��85��D���\��~��%��$k��|-�B�l�,��O��ap�j������e9��D�v��W��C5����-
��6��̙��9���1��uS�9�s��t���  �  ����2���π��c\��4�^s��pݾ����H�����W�"�2��y�eu	�� �����nA����;���<:���b�~A��(����X���R=�Q�e�B����U��S��H"��Z�z�q�T�}{/��o�����T��Q���� �N�C�|j�?d���:���ޒ�+݊��v��O���'����|y̾���f{�}�K��+�� ������ �]� ��h����'�(G���t������lƾh����##�%�J�	Dr��N���J������Dև��in�*�G�C$���	�||�������(,�KQ�#�w�ee���y���⑿g��
�k���C�
���`�� ���
���p���F��Y*����Aj�р	�@��\_�R$��<�/�`�TL��{N���޾�e���3���[��ဿ�����9B��~�����e��@?��.�����P���v��{�e�;��b��u��ݐ�̕�eꐿ~�����a���9�����_��������9"n��@I�&�0��� � �����0�L&�H|8�j�T�Fg}������þi�������"D�el�����͓�Ƞ������6���}\�P<7��X����XM�5�3)�I&L���r������c�������$�~���W���/�,��7�ܾ�C��΍�,�k�9K�{5��x'�K� ��j �?&���2���G�Og��f��֚��ދ־c���B+��R�(rz��h��bg���ޕ����v�EP�p,������W{����9�3��X��~�V쎿Gꖿ�A���f��6r�*J�e'#��@�(+̾V���)���7`��{C��0�]�%��C!��#�'+�o:�i�R��Vv��锾и��)��@�8�a��|�����e����ӓ��H��]�j��*D�'#�L���U������s5@��mf�����풿�  �  $�A��;���+��.�����Ǿ����JFu�	DA�X�m� ��ݽT�ƽ���H~��\弽��˽�I彼l��j#�~bL�����+	��*Ҿ���m��P�0���>���A���9��(��)���kξl%��Zٲ�����U�ᾞ��RW�a�2�+�?���A��68�ʁ%�'u��=�lH��˗���wd�N^5�rx�@���ǮؽwŽ�+��������ý�ս�R����0��^�Ii���%���a⾩o
�s�"��N6�^�@��\@�.�4�e� ��3	�]	�פľٳ�>����˾�d��M�^�&��V9���B��A��B4��]�ʀ�>۾uQ��v����Y��/�v��Ɉ������ҽ��ͽ*'ѽՉݽ�2�����;�%�ɲJ��a}����?�ɾ�����L��-��>��E�$<A��f2����@�����ľ�:��}þ�ݾU���,B1�l<A��G�WRA��W1���T���Ѿ����ġ��mW�_�1� z�/��h���΅꽍B�Z��6���`�y� �&�=�g��r��;���\�߾Ӭ��!�,x7�ŎE�:�H���@��\/�:����h�ݾ�ƾE�¾��Ѿu����f�&�(;��H���I�=j@�į-�x��U}��xɾ\����K�� bU�.c3�������t����U���x��4�
�`d���/�ltP���}�m��q6ľ ��A����*��n>��I���H�G�<���(�HM�I&����Ծ)�þx�ž��ھ�r�����w�-��X@�y�I�Z�G���:��%���8'��a���y����s�!^I��P+����$a	�`��������m���k�H�!��M;��_�7��v����Ӿ��w��2���C�P�J��ZF��v7���!��*
���IIξj�þT<̾
����GO�6}5��bE��  �  ��;�CY6��	'�AI�b�mþ֚��t�m�A������i��˽���ջ��[��^Eн���͍��$�(�L�3%��_ȣ��ξ��������+�_�8�b<��:4�(J#��I���fɾSP���+��ʖ��7bܾ]7�����-��:��;���2�i� ���	�tJ�LF���+���c�e6�[`�����hݽ�ʽd���m���2PȽ�cڽ"���#�M�1�{�]�$���U��_�ݾ���X�=1��6;�n�:�S^/��=����ׇ�KX��(���y����ƾ���i���"�w�3�k%=�Gd;�a/����Q���־!⫾�y����Y��1��
�� ��>�j^׽<ҽ�ս�#�=��� ��'��qK��l|�qE��5'ƾ�f��p����(��
9�t�?���;�I_-������`ܾ���������[
پq$ ����Q,�3�;��BA���;��x,��������Wξǥ����PX�2k3�<��:F����H����j�[o�ѹ�>�"�;Z?��[g�Ԙ��_L��=�۾�������i2���?�H"C�Tb;���*����4��m�ؾ�þ�'����;z���c��*"���5�	JB��"D��	;�I)������uƾXK���
���hV��J5����y��������X�����������1���Q�N�}��'��wf��W��6��s&�D!9�"ZC� �B�߁7�j]$����u��USо����w¾W־����n���/)�a�:���C��B�I�5���!���	���㾉�K}����s���J��e-���*�����+� ��������%�#�/=�n�`�%���h���ɐо������"�-��:>��E�`�@��o2���������5@ʾ\�FȾ⾽���;�:�0���?��  �  ��+�p'�I���������ﹾ�.���r���D���"�\>
�;t��ڽ��̽"lɽ�QϽ��޽c��ע��[*�|�N�O�~�T&��}Sþp������h)�,�(%����y�@ݾL��Uv��⽤�޲��zV;y����p]�L*�y�+�$��s��M ��־���������c��:�������W�'Jؽ�:ν��ͽ.�ֽ[D�6t�A��RP6��A^��E��� ���Ѿ�y��)�w"�V[+���*��� �����K���Ѿ�6��n����ͧ�D���1ھ]����$��--���+��!�����l��v˾����h��x�[��H6�~���]����g�.�߽qR�n�����S��-�{�N�!{�����?��L���=�:��]�)���/��	,�zl�������;�S���9���泾:˾k��_���:,��<1��z,�4$�� ����e�ľ ��s��~[��\9�� �c����p���%(��P} ����J<�F�)���D��ui��猾�����оR����l�>�$��T0��3��>,�%\���	��H쾤�˾)6��2�������F�ݾ�������'�z�2��44��I,�z���t��M澷��� ������Z���;���%���������=�I�
��S��.#���8�)V��/~�I��1���0�����C�d�*��}3���2���(�r�����z&ᾘ)ľ�x��j^��ޑɾ�1龞Y��6��+�94�er2�c�'�H&��G�q�ؾ�Ͳ��k���gu�)�O�	^4�g� �T���
�څ������[K��@+�O9C�)d������ɩǾ�A��p��� �~/���4�#)1��}$�E���]��vw׾�׾�����D��(8Ծ�9�������"��^0��  �  �O�W���;��q��ξ�[�� ����t���M���/�`x�/���5����{὏,����!�
����g�6��V��~��F������[׾�e��fy
����<��O�������epľ����'Q���/����AL��l�־���m�
����1��7���:������ľ��Ks��e�h��@E�)~)�������C��}潨�彣�｝;����&��nA���c�.x��W`���}�Pa��6����^���|���+[ھ�t��SG������ꗾB~���M¾���1{���;��Q��]o�Z��1j޾�+�����ƅ���b�:B�H
)������Lm��2�������=����ّ#�?�:��zX�R�}�>W������N�Ҿ�����	����yP����b���e��f�־�踾g��Nǜ��H��?춾jԾ�]��\��\���������RX���پ�F��e�������d��AF�@+/����ܐ��
�`	�F�����P$���7�
Q��0q�Xь��ɥ�0�þ��R��T������Ⱦ��f
�-�����Ӿ9p��l������,��`�ǾO��s����4�X��7���g�����:.վ����ꑚ��Z���Be�igI�p�3�Y�#��������k����!��m1�UHF�jFa�'ف��z�������Ѿ���{	��T��;���&�j�~�>~ʾ�-���ѥ��k�������=Ѿ�5�B�	���_}�{����E�M��vEʾ�,���ɒ�s|���[��`B��.�c| �D^��������,(���9��`P��m�S����̠�����x2ݾ�������?��3{�Y�����3����¾�ꭾ����p���俾Y2ݾ+����;��~��  �  �l��|�����1.Ӿ�1���ǥ�����"��8�a�'xG��]0�����5��.�B������T��[!�6�5���M��5i��O��^t���>��t¾��ؾa:�h;��>���L���۾-9¾2���j���/��6����a���������Ѿ��������"�|���̾����F�������M�w���Z��A��z+�Mk�j_�JZ�e���/�����)�͓>��W�rt��j��e]���Ჾ��ɾ��߾�;�������� ��©Ӿ�[���I��.5���������*���f���U���L۾�b�����!
���H�d�޾�4Ⱦ�]��gf��Z����t��Y�Q%A���,����A�J���-�B���'��T;���R��m�ͨ��������LL���mؾ�c��J��D� �?h��@��b~Ҿ��������l���h��ڣ��)C������>MѾLJ�x��B��) ��y��޾�Ǿɲ��f���F!��Mx��]��G�:4���%�����3���*���:���O��(h�ak��������̸�q�Ͼ�~澊�����������T�dѾ�-���ˡ�Xє������g���譾��ƾgi�,������;���������(ݾ+�ž�"��[ɜ�����z��ga�[NK��.9��,��	%��$���*��:7�S�H��X^��aw� ����k��Gk��/�¾�ھ�!�A� �����&��0���sɾME������9��
���Q���!���=�Ͼׄ�M����m��y���t��Xվ�w��@v������2����r�xvZ���E�7M5��@*��}%��m'���/�06>��JQ�*(h�,4��3���|���i��9�˾��F���wV�������?���S�ܾ�����O�������uǘ��5���R��Y�پ��7[��  �  o̾Q̾�Pƾ�W����������љ�����n����[m��kT�5=��`*��a����I� ��Y.��B�<}Z��s�V��u����ߜ�TI��;������
�Ⱦ~�;�̾�¾���h����ǋ�L�v���b�_�	El�������iڪ�߻��$ɾKEξu2̾ޒľ�̹�����z��C���싾Q���g��dN�'B8�U_'�����r�N�%�K�5���K�5d�k�|�@h�������蠾�a��"���þu/˾S�;Ҽɾ%���Ҭ�p���=���Ho���`��2c�C/v��3����q3���þO4ξ�
Ѿ;�0ľ���#?��R塾ɖ��h����~�"(f�TlN�^7:��,��&�8&)���4�ܗG��^��]x�����P���!
���c��x����¾�,;��Ӿ5Ծ��;M$��l����������w��n�E�v�fH��B옾/1��.j��YϾ��־g+׾U5Ѿ�@Ǿ"���� ��ä�"����
��|����k�!AT�H�A��;6�<33��;9���G�r\�*ut�w���
Y������^��.ֵ�����2;,�־�۾�ھ��оH���tC���Ϛ�#���9���X�~����!��	��)���;<�پ�޾_�ܾ��Ծ�ʾ�D��򦲾�_��n����������7n��X��G�1�=��=�)�E�A�U� ?k�U䁾5b��t\��]���6����z��*FȾ�EӾSd۾o6޾b�پLTξ��d먾�핾�h�� �������*�����������\����Ѿ9�۾)x޾fQھ�bѾ[ƾ%X����ȣ�7Q��39���p�\g���R��?D��=��h@�©K�e�]���t������h���4��J����е�����>;�׾q7޾�޾qؾ{Mʾ�������������`��U���J���`4���������H�ȾvQ׾�  �  '槾�:������Ȇ������5����4��z§����V瑾�����h��N�0U>�=�9��7A��T�-�n�2���X��0g���ǩ�*���⪰�[O���6���0���?��i6��j���7��a ��m�d���L���=�>;�C�D��^Y�Ru��։�Z+��N���T^�����-_���ױ�����[T���쬾bB���ϛ�M#��4�}���`�J�=�z_<���G� �]�"6z��V���>�����<���Ư��2��P|��.��\���Ȣ���^��\��6^���jx��x\��sG�E�<���>�f�L�v�d��S���ؐ�I����-���ۯ�GH�� ���%派�v��n���7c������}���ڌ���{���`��EM�%�D���H�p�X�T�q��釾3���t���:���7���!��r+���L��z������֯��q=��	-��o����Y}��Zc���Q��K��$Q�=�b���|������Ӝ��������r�������o��@u��B����%�������������rW�����8f��(V���Q�x�Y�I+m�n5��-����w�� ���,�����5���徾{ھ�!罾~���0��X���ܣ���Џ��X��J(k���\�ǨZ�^�d��|y��������؀������������������¾����=��:���N���ͫ�����Ў�	M����i���\�I	\���g��s}�����U7���'�����l���п�I��}���kA������7ջ�8��������s���2��1|�?�f���[��]]�!�j�s��乏�y�v��� Ƕ��E��������+¾	�������^���z��ݧ�by��CB���/y�Ece�'y\��
`��vo��	��U풾5��3"��Yɸ�P�������u�¾��¾�¾V뿾���u����W����������\�v���d�A�]�pXc��t�k)���A���+��Wű��  �  R����A����]��������ƾ �̾̾�ľ�T���2��0>��[<z���c�3]���g�娀��ǒ����w����ƾa;;q̾S�žJ4������L裾�����m�����%�j�ֽQ�;��0)����W���#�ߘ2��G���_�C�x�������IK��5������������ʾ\oξj˾\���GT���w�����"s�Yya��|`�Dp�h���,�����/���dʾ�4ξL ˾�¾偷������/��&���_���'K{��rb��9J��5�T�%�<?�e��Y/*��<���R��cl��삾��&�������W�������CȾ.�Ͼd�Ѿ�&̾Ԍ��㦭�ෙ��r��uRt���h���m�����sx��6����7����ɾ��Ҿ�fԾ�XϾt�ž_l��0����h��%F��!ˌ�5���u�h�NVQ�(�=�h1�B�,�1��
>���Q���i�7�������"˙� ������#G��L�Ǿj�Ѿ��׾�׾�3Ͼ���3���/ę�1ӈ��{��du�I"��L)���{���س���ƾn5Ծ@�ھ��پ\ Ӿ�Ⱦ�$������~���c��Џ�����o���X���G�kV=��;�@C�ÛR���g�,��ʌ���n��'������V�ƾ�Ҿ��ھ�޾�t۾��о�E���_���显�`��������^����ϖ�>���[󽾞Ͼ'VھJ1޾c۾��Ҿ��Ǿ(׻�F[���)��oÙ����C���j�U�T���D�I=��">�cH�6GY�+�o�~?��.���ߝ�������9���׾���ʾ6Wվ��ܾp�޾;پ�I̾�=���#��o����4��d�������������s���?ž?�Ծ�uݾ<�޾��پ�Kо��ľ���g̭�`���	��Hኾ�|�	e��WQ��D�?�=8C���O��c���z�.܉�
0���  �  ɀ�����ݦ��q���tԾJ��[-�������g��޾�ž����-۔����.���E����������q#̾4&�����'O�������E�*о���G���FA��X|���^���D�7<.����D��i���-��k	������%���:�;KS��Ko�Ѷ���G��{w���pƾ|�ܾBNﾮ����@��eX�,ؾ���T��͏��6��͑������c��� ��QIվ6�ID���������޾l�Ⱦ����[*��ST��[r�u�U��1=��
(��Qd�����6��#�I���/���F���`�,�~��^���������j9Ѿ��澃���-��i���g��Z�Ӿ�2���堾�<��qf���Ê��˘������ɾ�@������@ ������%��޾��Ǿ�����������hv�I�[��#D�(e0�;(!�.��vG�}���!�CK1�qE�95]��Nx�X����_���ű��[ȾY^߾��+� �cH��}���*�WѾ`��.���[葾Ͼ���є�F����*��,�ؾj-�;� ����B� �M���ݾ��ƾ�����������z�Dxa��iK��59���+��T$�	X#�|�(�h�4���E��*[�q�s��������A����Ŀ�f�־2�Wu��������T��T���;�3��Ԧ������e���͝�x��T�ʾ6(�u�������jT ����v�ؾ�����Q��y{��R0��
v�n1]���G�x�6�n�*���$�6m%���,��4:���L���b�Qy|��⌾�����9���-ǾBU޾���	�����d�|s��aྺ�žq��FE���>���j���@���W��n�Ծ� �� �Q�����������辐,Ҿ@����즾:����{����o��7X��%D�F�4�
*�\�&���)�>k3��B�:bV���m�YT���  �  ��u����D����о@K�?��2��i����4�˫�ɾ�@���������
�������о�m�p����������W���뾿�ɾ�����,��|n���I�*�,�b��]���󽚾潮v佄��H�����;�"�۝<��]�彃��r���һ��=ݾ��������I�M��� �1X�����K	��^;���T���3��itܾx���X��>��b	���ߛ ���ྦྷ���F�����sa�(�?��.%�m�������轭[� e��,��Q��x�.���K� �o�������9�ɾ'��n�����u��v���R���پ@%���ţ�{ٙ���������˾Et�(�DN����f��R5�����2ܾ�D���띾@g��GYc�fBD��,����Ŵ�1��qf��I�������a�-�q�E��d��Ņ�}Ꝿ&Ế��۾!5���y����Y���M���
�y	����Ծ*����i������慨V���q)ݾT9������=��D�pu����:��g�׾`�������,��Ef�1�I�c�3�5#�o��L���L������S�.��C�1]�mX~� ���í��̾8~�K)����	���M�������>�xϾDx���ަ����C(���̾M�A�����M�������1����\8Ͼuj��p0��Հ�ȶ_�pE�4�0��`!��[�<���F��D�c�$���4�5�J�fg��s���盾pA���־����%'�1��������b����l�VƾHʯ�F�������P��i׾����s�����5����m�����׬ž�O��������w���X�i2@�&�-�� ����P��Ih�3�j8,��p>�$QV���t��  �  :~t�*ї�����Y:�"����g�'�3�+��&������6��@P���	������Fʭ��>Ǿ����+
�B��O�(� ,��%�C4�)���ܾ�F������$k�w�?����Y@�.����ٽXνN\̽��ӽc�~ �ַ�.�0�yW�娄�pv��Гʾ����*��k �#�*�{�+�qD#�Z/�Et��L8׾�;��H榾��˄��_-Ӿ��������!��4+��;+���!�M,�.���ξ������5�[��S4��i�r����9�׽;н�9ҽ��ݽl��L
��x!�A6A�ák��L��!u���d۾�
�`�pl&���-���+��m �~�������ϾU4���^��-A��S(þɿ�Ȉ�����(��z/��T,�!A �����9/Ⱦ�l��Z7���C[���7�E��r��1���~��r�����fe �����V���8���[��������)�ƾm%�;M�g$ �"%-�b{1�[,�B��8��C�`̾:絾񐯾����Ӿ�;��֋���"�^U/�ʽ2�wm,�N��tU
�B)�����w[���|���\��?<��M%��N�b�
�-���,��N	�KK�� �65�wVQ�עw������Ĵ���ھ�~��C�v}(���2���3��A+��&�'-����Ⱦw����ŵ��Wž�c�������)��*3�#73���)��2�.��b�޾g7�������{��aT�uI7��Y"�����
�������q����}�&�L]=���\��T��"���N������	�k��/�,��R4�C2���&����H� �Sܾ�5���5��^칾V�ξa�H�!��
C.�F�4�%�1�z%��'�H ��~�Ҿ�Э�-��� �o��(L��2��t�0���v����c�E�P7�y<0�V�I�=4l��  �  K�v�������ž/���m��Y&(��7��<�v�5�w=&����S\���;�$���歾�O���վ�S��E��"�*��f8�d<���4��$�����꾴㼾�����l��D<��e��� �چ�o{˽(�������(�ŽGֽ�����I�+���U�솾8ު�O6־�%�	����.��z:��;��#2�" ��	��c�j�ľ�����}������%������9f0�&;�};��D0�&6����3۾���F?��'�Z�w�/����s���VGڽ��ɽ��½�Ľ��Ͻ������N6=���k�tє����e�����O�#�;G5��=�4v;���.�T�����޾����"Ƴ�%.���lо����Pz��r'�f8� ?��;�s�-��	��� ���ҾsΨ�߸���X�?92�k���-�T��㽙3߽���B�Co�c ��)3�IY��9��˘��ӱо��������-���<�0�A�Jt;���+�,s������پ� ���빾�~ž��:n�:N��1���>�ʹB��r;���*��p�Q]����ʾlN�������mX���5�8��:�����N���s����:�w�
�V�H.�3IL��Bv��8��#+���}澎D�r�"���6���B���C�� :���'�Ǔ�)B��.�Ծ�a���P��l�Ѿ���f��t�%�X8�1C�l	C�E8��;%�u��.�c'��t[����z�N�O��0�����h�C��0}���E ��J�}O��I�B�6�0�X������)���Ⱦ���[�f9*���;��GD���A��5��� ��:
�p���̾ۜ����ľl�۾� ��	���,�!y=�]�D�HA��33��?��*���ܾ�2������ym�~�F���*����e��N���!�"(���
���T)��C��ei��  �  vx� ����ɾ9���ȑ��-�X�<���A�zv;� #+�B��h�����ҾI������:c����ھD�<,���/��>���A��@:���(�[g��+3���0����l��r;�p���B��Q�۽��ƽ�2��+g���;���ѽ�I�H���*�ʸU�(���1e��R�ھ�c��0���3�4@�B�A���7���$�FZ�Q'�kQɾ�N��Y6��d0ƾ�{�w�
��"��5���@� �@�ʈ5���!��	�I�߾�����r����Z�o.������Q�ս	Ž,E���G��]+˽+�Ǧ ��1��B<���l��Q��v���=�Wn��X(�[�:���C��)A���3���Ё�}	�J$žxq��,
���"վn���Zf��@,�a�=��OE�8wA�3�2������C�־n���ꁇ�b�X�w�0�װ�F�������޽r�ڽ�߽&��;�y���1��X��↾~���klԾq���1�2�HB��UG�~A���0��y����޾��ľ������ɾ9#�A��ǆ ��6�ʖD���H���@�̏/�Y(�֨��E�;����a��=�W�(4�գ�/d�o�6&��/E��������Ũ�k,���J� Cv�6F������c��u��)I'���;��=H��I�d�?��,�M����*پ�#žF	ľ!־DP��P��U*��=�z�H���H��=��)�/���ﾷ���	����#{�wsN��.����
��c��!��V*����.��F�-5�x�W��σ�v�����˾�(�����1�.��'A�|J���G�s,:�AM%�����/��"ѾHþ��ȾX��O��W��+�1���B�;�J���F��68��Q"��+	���ྮ\���ۑ��m��	E�(�(����4	�kF�y�������y�"T���&�dB���h��  �  K�v�������ž/���m��Y&(��7��<�v�5�w=&����S\���;�$���歾�O���վ�S��E��"�*��f8�d<���4��$�����꾴㼾�����l��D<��e��� �چ�o{˽(�������(�ŽGֽ�����I�+���U�솾8ު�O6־�%�	����.��z:��;��#2�" ��	��c�j�ľ�����}������%������9f0�&;�};��D0�&6����3۾���F?��'�Z�w�/����r���TGڽ��ɽ��½ �Ľ��Ͻ�������K6=���k�rє����b�����M�#�:G5��=�3v;���.�S�����޾����"Ƴ�&.���lо����Qz��r'�g8�?��;�t�-��	��� ��ҾvΨ�Ḇ��X�B92�m���-�T��㽙3߽���B�Ao�a ��)3�EY��9��ɘ��ѱо��������-���<�/�A�It;���+�+s������پ� ���빾�~ž��;n�;N��1���>�˹B��r;���*��p�S]����ʾnN�������mX���5�;��<�����Q���u����:�x�
�V�I.�3IL��Bv��8��#+���}澎D�r�"���6���B���C�� :���'�Ǔ�)B��.�Ծ�a���P��l�Ѿ���f��t�%�X8�1C�l	C�E8��;%�u��.�c'��t[����z�N�O��0�����h�C��0}���E ��J�}O��I�B�6�0�X������)���Ⱦ���[�f9*���;��GD���A��5��� ��:
�p���̾ۜ����ľl�۾� ��	���,�!y=�]�D�HA��33��?��*���ܾ�2������ym�~�F���*����e��N���!�"(���
���T)��C��ei��  �  :~t�*ї�����Y:�"����g�'�3�+��&������6��@P���	������Fʭ��>Ǿ����+
�B��O�(� ,��%�C4�)���ܾ�F������$k�w�?����Y@�.����ٽXνN\̽��ӽc�~ �ַ�.�0�yW�娄�pv��Гʾ����*��k �#�*�{�+�qD#�Z/�Et��L8׾�;��H榾��˄��_-Ӿ��������!��4+��;+���!�M,�.���ξ������5�[��S4��i�q����6�׽7н�9ҽ�ݽd��L
��x!�:6A���k��L��u���d۾�
�]�ml&���-���+��m �}��
�����ϾU4���^��.A��T(þʿ�Ɉ�����(��z/��T,�$A �����>/Ⱦ�l��_7���C[���7�J��v��6������r�콾��de �����V���8���[��������$�ƾh%�8M�d$ �%-�_{1�Y,�B��8��C�^̾9絾񐯾����Ӿ�;��׋���"�`U/�ͽ2�ym,�Q��vU
�G)�����{[���|���\�@<��M%��N�e�
�0���,��N	�LK�� �75�xVQ�עw������Ĵ���ھ�~��C�v}(���2���3��A+��&�'-����Ⱦw����ŵ��Wž�c�������)��*3�#73���)��2�.��b�޾g7�������{��aT�uI7��Y"�����
�������q����}�&�L]=���\��T��"���N������	�k��/�,��R4�C2���&����H� �Sܾ�5���5��^칾V�ξa�H�!��
C.�F�4�%�1�z%��'�H ��~�Ҿ�Э�-��� �o��(L��2��t�0���v����c�E�P7�y<0�V�I�=4l��  �  ��u����D����о@K�?��2��i����4�˫�ɾ�@���������
�������о�m�p����������W���뾿�ɾ�����,��|n���I�*�,�b��]���󽚾潮v佄��H�����;�"�۝<��]�彃��r���һ��=ݾ��������I�M��� �1X�����K	��^;���T���3��itܾx���X��>��b	���ߛ ���ྦྷ���F�����sa�(�?��.%�l�������轥[�e��&��J��o�.���K��o�鉎���2�ɾ ��j�����u��v���N���پ>%���ţ�{ٙ����	�����˾Ht�*�GN����i��U5�����!2ܾ�D���띾Fg��RYc�nBD��,����ɴ�3��qf��I�������Z�-�i�E�ۘd��Ņ�vꝾẾ��۾5���y�}��V���M���
�u	����Ծ)����i������慨X���t)ݾX9������=��D�su����:��n�׾g�������,��Of�:�I�k�3�5#�t��P���L������T�.��C�1]�mX~� ���í��̾7~�K)����	���M�������>�xϾDx���ަ����C(���̾M�A�����M�������1����\8Ͼuj��p0��Հ�ȶ_�pE�4�0��`!��[�<���F��D�c�$���4�5�J�fg��s���盾pA���־����%'�1��������b����l�VƾHʯ�F�������P��i׾����s�����5����m�����׬ž�O��������w���X�i2@�&�-�� ����P��Ih�3�j8,��p>�$QV���t��  �  ɀ�����ݦ��q���tԾJ��[-�������g��޾�ž����-۔����.���E����������q#̾4&�����'O�������E�*о���G���FA��X|���^���D�7<.����D��i���-��k	������%���:�;KS��Ko�Ѷ���G��{w���pƾ|�ܾBNﾮ����@��eX�,ؾ���T��͏��6��͑������c��� ��QIվ6�ID���������޾l�Ⱦ����[*��ST��[r�u�U��1=��
(��Nd�����6��#�B���/���F���`��~��^���������a9Ѿ���{��-��b���b��U�Ӿ�2���堾�<��qf���Ê��˘� ���ɾ�@������@ ������%��޾�Ǿ�����������hv�T�[��#D�.e0�?(!�0��vG�{���!�=K1�qE�/5]��Nx�Q����_���ű��[ȾP^߾��&� �_H��}���*��VѾ]��,���Z葾Ͼ���є�H����*��0�ؾp-�?� ����F� �V���ݾ��ƾ�����������z�Oxa��iK��59���+��T$�X#��(�j�4���E��*[�r�s��������A����Ŀ�f�־2�Wu��������T��T���;�3��Ԧ������e���͝�x��T�ʾ6(�u�������jT ����v�ؾ�����Q��y{��R0��
v�n1]���G�x�6�n�*���$�6m%���,��4:���L���b�Qy|��⌾�����9���-ǾBU޾���	�����d�|s��aྺ�žq��FE���>���j���@���W��n�Ծ� �� �Q�����������辐,Ҿ@����즾:����{����o��7X��%D�F�4�
*�\�&���)�>k3��B�:bV���m�YT���  �  R����A����]��������ƾ �̾̾�ľ�T���2��0>��[<z���c�3]���g�娀��ǒ����w����ƾa;;q̾S�žJ4������L裾�����m�����%�j�ֽQ�;��0)����W���#�ߘ2��G���_�C�x�������IK��5������������ʾ\oξj˾\���GT���w�����"s�Yya��|`�Dp�h���,�����/���dʾ�4ξL ˾�¾偷������/��&���_���&K{��rb��9J��5�Q�%�8?�`��R/*��<���R��cl��삾	���������M������}CȾ%�Ͼ\�Ѿ�&̾͌��ަ��ܷ���r��rRt���h���m�����vx��;���8����ɾ��Ҿ�fԾ�XϾ}�žil��:����h��-F��(ˌ�;����h�VVQ�-�=�k1�C�,�
1��
>���Q�~�i�1�������˙� ��󃰾G��B�Ǿ`�Ѿ��׾�׾�3Ͼ���.���+ę�/ӈ��{��du�J"��N)���{���س���ƾv5ԾH�ھ��پe Ӿ"�Ⱦ�$�� ����~���c��Џ������o���X���G�pV=��;�@C�śR���g�,��ʌ���n��'������U�ƾ�Ҿ��ھ�޾�t۾��о�E���_���显�`��������^����ϖ�>���[󽾞Ͼ'VھJ1޾c۾��Ҿ��Ǿ(׻�F[���)��oÙ����C���j�U�T���D�I=��">�cH�6GY�+�o�~?��.���ߝ�������9���׾���ʾ6Wվ��ܾp�޾;پ�I̾�=���#��o����4��d�������������s���?ž?�Ծ�uݾ<�޾��پ�Kо��ľ���g̭�`���	��Hኾ�|�	e��WQ��D�?�=8C���O��c���z�.܉�
0���  �  '槾�:������Ȇ������5����4��z§����V瑾�����h��N�0U>�=�9��7A��T�-�n�2���X��0g���ǩ�*���⪰�[O���6���0���?��i6��j���7��a ��m�d���L���=�>;�C�D��^Y�Ru��։�Z+��N���T^�����-_���ױ�����[T���쬾bB���ϛ�M#��4�}���`�J�=�z_<���G� �]�"6z��V���>�����<���Ư��2��P|��.��\���Ȣ���^��\��6^���jx��x\��sG�@�<���>�_�L�m�d�S���ؐ�B����-���ۯ�=H������派�v��e���.c��햦�w���ڌ���{���`��EM�$�D���H�t�X�[�q��釾$3���t���:���7���!��|+���L���������߯��y=��-��t����Y}��Zc���Q��K��$Q�8�b���|������Ӝ�����򰲾i�������o��6u��8����%����������}��mW�����8f��(V���Q�{�Y�N+m�r5��2����w�����%,�����"5���徾�ھ�+罾����0��`���⣞��Џ�Y��Q(k���\�̨Z�b�d��|y��������ـ������������������¾����=��:���N���ͫ�����Ў�	M����i���\�I	\���g��s}�����U7���'�����l���п�I��}���kA������7ջ�8��������s���2��1|�?�f���[��]]�!�j�s��乏�y�v��� Ƕ��E��������+¾	�������^���z��ݧ�by��CB���/y�Ece�'y\��
`��vo��	��U풾5��3"��Yɸ�P�������u�¾��¾�¾V뿾���u����W����������\�v���d�A�]�pXc��t�k)���A���+��Wű��  �  o̾Q̾�Pƾ�W����������љ�����n����[m��kT�5=��`*��a����I� ��Y.��B�<}Z��s�V��u����ߜ�TI��;������
�Ⱦ~�;�̾�¾���h����ǋ�L�v���b�_�	El�������iڪ�߻��$ɾKEξu2̾ޒľ�̹�����z��C���싾Q���g��dN�'B8�U_'�����r�N�%�L�5���K�5d�k�|�@h�������蠾�a��"���þu/˾S�;Ѽɾ%���Ҭ�o���<���Ho���`��2c�=/v��3����j3���þG4ξ�
Ѿ;�0ľ���?��J塾ɖ��h����~�(f�LlN�Y7:��,��&�:&)���4��G�#�^��]x�����W���)
���c�������¾�,;��Ӿ>Ծ��;T$��q���񸙾�����w��n�C�v�dH��>옾*1��(j��RϾ��־^+׾K5Ѿ~@Ǿ���� ��ä�����
��v����k�AT�C�A��;6�<33��;9���G�y\�3ut�}���Y������^��7ֵ�����2;6�־�۾�ھ��оN���yC���Ϛ�&���;���]�~����!��
��)���;<�پ�޾_�ܾ��Ծ�ʾ�D��򦲾�_��m����������7n��X��G�1�=��=�)�E�A�U� ?k�U䁾5b��t\��]���6����z��*FȾ�EӾSd۾o6޾b�پLTξ��d먾�핾�h�� �������*�����������\����Ѿ9�۾)x޾fQھ�bѾ[ƾ%X����ȣ�7Q��39���p�\g���R��?D��=��h@�©K�e�]���t������h���4��J����е�����>;�׾q7޾�޾qؾ{Mʾ�������������`��U���J���`4���������H�ȾvQ׾�  �  �l��|�����1.Ӿ�1���ǥ�����"��8�a�'xG��]0�����5��.�B������T��[!�6�5���M��5i��O��^t���>��t¾��ؾa:�h;��>���L���۾-9¾2���j���/��6����a���������Ѿ��������"�|���̾����F�������M�w���Z��A��z+�Mk�j_�JZ�e���/�����)�͓>��W�rt��j��e]���Ჾ��ɾ��߾�;�������� ��©Ӿ�[���I��-5���������'���b���P���L۾�b�����
���H�[�޾4Ⱦ�]��_f��S����t��Y�I%A���,����>�J���-�F���'��T;���R��m�Ԩ��������UL���mؾ�c��J��H� �Fh��F��g~Ҿ��������l���h��٣��&C������:MѾFJ�x��>��) ��y��޾�Ǿ����^���?!��Ax��]��G�44��%�����5���*���:���O��(h�gr�������̸�z�Ͼ�~澓����������$T�iѾ�-���ˡ�[є������g���譾��ƾhi�-������;���������(ݾ+�ž�"��[ɜ�����z��ga�[NK��.9��,��	%��$���*��:7�S�H��X^��aw� ����k��Gk��/�¾�ھ�!�A� �����&��0���sɾME������9��
���Q���!���=�Ͼׄ�M����m��y���t��Xվ�w��@v������2����r�xvZ���E�7M5��@*��}%��m'���/�06>��JQ�*(h�,4��3���|���i��9�˾��F���wV�������?���S�ܾ�����O�������uǘ��5���R��Y�پ��7[��  �  �O�W���;��q��ξ�[�� ����t���M���/�`x�/���5����{὏,����!�
����g�6��V��~��F������[׾�e��fy
����<��O�������epľ����'Q���/����AL��l�־���m�
����1��7���:������ľ��Ks��e�h��@E�)~)�������C��}潨�彣�｝;����&��nA���c�.x��W`���}�Pa��6����^���|���*[ھ�t��RG������ꗾ@~���M¾���/{�߻�7��N��Zo�Z��*j޾�+�����ƅ���b��9B�A
)�������Hm��1��������=����ߑ#�G�:��zX�]�}�DW������U�Ҿ#�����	����|P����d���e��i�־�踾g��Nǜ��H��>춾jԾ�]��Z��\���������JX���پ�F��_�������d��AF�9+/����ؐ��
�`	�G�����P$���7�Q��0q�^ь��ɥ�7�þ��U��T������ʾ��f
�1�����Ӿ<p��n������,��a�ǾO��s����4�X��7���g�����:.վ����ꑚ��Z���Be�igI�p�3�Y�#��������k����!��m1�UHF�jFa�'ف��z�������Ѿ���{	��T��;���&�j�~�>~ʾ�-���ѥ��k�������=Ѿ�5�B�	���_}�{����E�M��vEʾ�,���ɒ�s|���[��`B��.�c| �D^��������,(���9��`P��m�S����̠�����x2ݾ�������?��3{�Y�����3����¾�ꭾ����p���俾Y2ݾ+����;��~��  �  ��+�p'�I���������ﹾ�.���r���D���"�\>
�;t��ڽ��̽"lɽ�QϽ��޽c��ע��[*�|�N�O�~�T&��}Sþp������h)�,�(%����y�@ݾL��Uv��⽤�޲��zV;y����p]�L*�y�+�$��s��M ��־���������c��:�������W�'Jؽ�:ν��ͽ.�ֽ[D�6t�A��RP6��A^��E��� ���Ѿ�y��)�w"�V[+���*��� �����K���Ѿ�6��m����ͧ�D���1ھ[����$��--���+��!�����l���u˾����h��q�[��H6�y�	��X����g�.�߽rR�r�����S��-���N�#!{�����?��Q���=�=��`�)���/��	,�|l�������;�S���9���泾:˾k��]���:,��<1��z,�2$�� ����`�ľ ��o��w[��\9�� �`����n���%(��Q} ����M<�J�)���D��ui��猾�����оW����l�A�$��T0��3��>,�'\���	��H쾦�˾*6��3�������G�ݾ�������'�z�2��44��I,�z���t��M澷��� ������Z���;���%���������=�I�
��S��.#���8�)V��/~�I��1���0�����C�d�*��}3���2���(�r�����z&ᾘ)ľ�x��j^��ޑɾ�1龞Y��6��+�94�er2�c�'�H&��G�q�ؾ�Ͳ��k���gu�)�O�	^4�g� �T���
�څ������[K��@+�O9C�)d������ɩǾ�A��p��� �~/���4�#)1��}$�E���]��vw׾�׾�����D��(8Ծ�9�������"��^0��  �  ��;�CY6��	'�AI�b�mþ֚��t�m�A������i��˽���ջ��[��^Eн���͍��$�(�L�3%��_ȣ��ξ��������+�_�8�b<��:4�(J#��I���fɾSP���+��ʖ��7bܾ]7�����-��:��;���2�i� ���	�tJ�LF���+���c�e6�[`�����hݽ�ʽd���m���2PȽ�cڽ"���#�M�1�{�]�$���U��_�ݾ���X�=1��6;�n�:�S^/��=����ׇ�KX��(���y����ƾ��i���"�v�3�j%=�Ed;�`/����Q���־⫾�y����Y��1��
�� ��>�h^׽<ҽ��ս�#�@��� ��'��qK��l|�tE��7'ƾ�f��r����(��
9�u�?���;�J_-������`ܾ���������Z
پp$ �~���Q,�2�;��BA���;��x,��������Wξǥ����LX�/k3�9��9F����G����k�\o�ҹ�A�"�>Z?��[g�֘��aL��@�۾�������i2���?�J"C�Ub;��*�	���4��n�ؾ�þ�'����;z���c��*"���5�	JB��"D��	;�I)������uƾXK���
���hV��J5����y��������X�����������1���Q�N�}��'��wf��W��6��s&�D!9�"ZC� �B�߁7�j]$����u��USо����w¾W־����n���/)�a�:���C��B�I�5���!���	���㾉�K}����s���J��e-���*�����+� ��������%�#�/=�n�`�%���h���ɐо������"�-��:>��E�`�@��o2���������5@ʾ\�FȾ⾽���;�:�0���?��  �  R)����۾�M��D𡾶���R�٨&��k��4ֽQG��Ι��<���߁��p�G}��@����I��>W��d�ὠ���0�^�^����0~��?�Ǿ��c�����3n�B׾Q��ՠ�f ���x���r�������:���˾���B���������oԾ<��������w�OGE�?x�h����ͽH(��̻������'��{ǃ��a��ե�����sȽ&���.���?�6q��V��"���a�оɏ����L-�F�徹�ξ���"���ϒ��W�t���w���__�����l־��4��#*���q� ξ$���Y���Sl�(&=���������Ͻ�������F������1���is���E��˴ɽ5-��n���0��;\�=n��4����ľ�8���K)��C'��$�;~T�������s�����������#����˾�徇������LF�����5*˾�Ҭ��쎾}�h��<������u�߽��ǽ�'��r����Y��^ ��� ���yҽ�C�?�&��XK���y�7���z	��0վ�����Ch����G���˾௾�M��^����#��Gw�������"���ܾ��b��{����E侂�Ǿ���M틾�Ge�=^<����A��s�i�ֽ��ɽ2ýt�½cdȽ��Խ$�������i�7�ڟ_�ߋ��RR��)�þJ��M���z��������S�޾þ]���vO��N��J���!��5���zɾť侮	���n�N����4C۾���%%�� +��A	W��1�rj�.�?a潩Խ�lɽ�BŽ�ǽu�ν}�ݽj����0�p�$��F��,q��ْ�1���3,Ͼ#��UG���8��� �:=�׾O(��5>��$����j��U�������]��V>Ծ��(8 ��  �  �}�P�"Zվ��������Ձ�0kP�&����v�ؽoM�����|g��_섽縂� ���Ґ��}��SD�����B]�ޡ/�R@\�ë�� ڥ�1�¾��ھԅ�()��zѾ驷����Z���s��n�n�����˫�Ŭƾ�ݾ����z��I�ξ�o������t�n�C��@�����ϽII�����񭍽F-��Dˆ���ݘ���� /˽������XT>���m�ނ���篾��˾�q��=�E��E�߾�hɾ.ʮ��H��Fс���o���r�N#��_�>i��y�о���Đ���S��ɾ�������8ei�<�������ҽtӷ�G��"]����������/���P}����̽9��K�0{0��&Z��_�������W���ھ���~��ګ�GྠȾ"O���b���ׄ�M[}�O����链8���H�ƾ��߾8���+�����-�H�ƾ�t��þ���Pf�V<���5�����(˽^Q������QX�����/ý/�ս`.����&�_J�#w��*��me��.CоJ��BV��'��:U�W�߾�kƾ{%��dV�����ȹ�����P���'绾@�־e��r4���S��\���޾�þu������c��&<�-��������j"ڽ��̽i7ƽ�Ž��˽��׽�3�N.�+��&�7� ^��ن�a~��u��۾���4V��������>pپڿ���$������v����ӈ�5>����9�ľI)߾���8��|��-��L־չ�����˳����U�?�1��i��� ���A׽�̽�CȽ�ʽҽ/'�Ч��bl�qW%�ڔE�Io��ː��]����ʾ��4���/���F���Aa꾁Ҿ=#��4��[�����Q,���霾�r��u`Ͼ�W����  �  $�ھ�nվ��ž�7��򁕾�Ex���J��%�-����oH���V��Ga��p������*��r暽jЬ�ǽ�O뽝	���-���U�q@������m��P�ʾ��ؾ7�۾v�Ӿ����X�������[}�n�d��R`��ap��"���蟾�%���̾;�پ��۾ĄҾ�$���������j���?�0����3�ؽq~���3���}��ݖ���.��aA��1���]���qԽJZ������;��,e�����0ꤾ�`���оZ�ھ�=ھ��ξ����𠢾n���/t��6b�ce�g�{���������y����rԾ�޾��ܾ�о����
�������
b��9�N^�k� �mܽ�%½�i��2���W���(��T����ƾ�R�ֽ�0�������/��1U�k���J��5��m˾�ܾ� �]�޾k�Ͼ�������2d����z���o�9qy��&��𛠾����Ͼ�߾S���4ྈ�о��`e��c����`�O;�+^�����콡wս�Gƽ�+��T���.����;ͽ`�߽(���+��g�(��H�fp�M���=����þ��ؾ8Y�X�� ���Oо|U��D����P���������!��� ���OȾsݾK��B��ͼ�sUо76��j4���s��*�_�Xp<�B� �������]a���ֽ[�Ͻ�0Ͻ9Cս��st��5�	����wz8�n�Z���������﴾kn;�����S�}�޾��ʾ���Iq������@����ҁ����_��y*��t�Ͼ]Y����e���fݾ��Ⱦߛ��S˕��|�ߕS��3����j����b��)ֽ�ѽY�ӽ�ܽt��\�����'�AE��$j�,s��_���������վq��I�����پ�ľ�ӫ�����9��{ㅾ�#��
k�������3ؾI��  �  Ɍ��j��������^��� kj���E��&��s�3x򽌰ҽ;w��!W��?O������<���$������?ڽW��3{��+.�6�N�q}t�ᎾY/���B������2�����~'������3����d�u�O�~�K��Y��Rv�}z������v����y��U����h��]ӫ�a����ڃ��`��'=�I ��i��K�Q�ͽ����"���=���Ǡ�٭��˼����ʽ�2罧�����>69��o[�ON����������Ҹ����������\���ϐ���z���\�ìM�B!P���c�Q�������P��^O��:�þ	�¾t�������ɔ�[/���:Z�Za9��]����8��'�ս��½5���ݲ��ﵽ�P����ѽ2@����/��C2�e�P�*>u�<䎾❣��$���\þ��Ⱦ�ľX&��	ť�I`��]'~���d�a[���c��T|�)j��I,���Y����ž@˾�2Ǿ�躾���l�������[���<���#�ͨ�� �Ĕ轁8ؽNϽ-"ͽz�ҽ�k߽/5��	�L���-���H���i�ݼ��l��^ɰ�J���F�̾�+ϾTKȾ����63��,��=|��m�n��!k��(y�� ������Z"���ľ#�Ͼ*�Ѿ7�ʾ���¨�`����� &]�b�?�:5(�]\����)��"�F���߽���C�������.�1t%��y<�X�X�+N{��G�����X���Q�Ⱦ��о� о�ƾ7��u������l|�˥l�Ȭn�&ꀾ�Q��|�� y��y/ɾ�OѾj<оdƾV(䡾�<��;t�'AS��8�X;"����������W�N$��U���My��8�ծ�І.��aG���e�����J��� ��4���:�;��Ҿ��ξ�B¾����W6������c�w�n��v�d#��{4��Rɭ�y���Kξ�  �  �2��!���ޘ����%�|�#J`�u2F�G/�:���	�f�򽙞ؽ4�Ľ�����'���ݺ�Y&ɽ��޽.���؅�� ���4���L�H�g��A��fM��{����	��.���z���E��Dx��rbb��+G��m6��H3��T>�2�U���t�缊�,��������:���b��(��F�u���Y��@��[*���������\<սt�ýT��Շ��#����ҽXJ�߸�&��¹'� �=��FV� �q�fM����������&��˂��c��}o���^x��$Y�|7A��!5�;67�	'G��b�_���1ޑ�7�6��.���XU��=8���t���Jr�}cW�Dh?�@l*��	�X��:���9'߽Uѽ�z˽{Ͻ�g۽����������&��L;��[R�=al��c���Ò�5����_���^���|��d-���b��c|��^�C~J���B���I�<�]��!{�XC��&��������魾�ܫ�����si���9�� v�;\��!E�\1�q���0\���;�X���9��Y������"�F�'�V|:�ïO��g��[���ˏ�睾'����ְ�����������9!��|����e�N?U���R���]�cu��O���ܚ����6O���Ǵ�Yo������bL��Lڊ�)�y�р`�->J�;�6�Um%�st��3
�yY�k��|���* ����خ��L#�94��lG�G]��"v�%����N��"ˤ�*'���6������!���e������x��q`�3�S��U�Ze��t�$鏾V���0Ǭ�	ҳ�h��������c��Ɏ���1��aq�eDY�zD�P~1�J!����
��� ������o���{�p*���%�*�S<�wnP��Tg�ݟ��sˎ�o'���᩾c���쪵�^���}K���_��j懾-r���]��U�d\��o�uU���ږ��-���I���  �  �����������\}�[�n���_��	Q��	B��d2�m�!��O��������ڽ�dֽ�ݽ�F�V��K���b&���6�mF��}U��d���s�G󀾜���ED��X܇�������o�W�U�=���(�s�d���2"��	4���K���e��C|�5��E���ß��;-���5{�\_l��X]�DnN�5?�E7/������ߡ���8�H�۽:۽a*潈������p�b-�5#=�W^L�
<[��2j�;y� A�����wo��灆�1~�%Ih�=O�P7�t�$����B�D�)�\y>�	X�q�q�M���`J���p���W���#���|� �m���^��P���@�	�0�~m ����no�r��o����Zv �=������-���>���N�@^�,]m��|�Ѫ����Oя��a�������gn�w,U���>�o4/��)�^�.�lT>�8U�^o��ă��+��YR���ⒾĈ��!����Z����u�;�f��X��H��^8�i(����!���G��j����0�*�_/��@��?Q��a�%Qp�}��[������$>�����SΕ���8C��?t�o�[�3G���:���8��A���S�X�k��Ⴞ�I��E��ř��ј�Y��k����F���m}��hn��_� O�{:>�Z�-�i��G���d����B�O�+�<�m�L��\�k"l�f{�k������DG�����z��	����������n�tV�|�C�@G:���;�joG��[�¹t��iW���ߗ�Lי�񚗾�M��?X���܃���x���i�}Z�$FJ��9�)�l���E�~�����B�Kr#��2���C�K)T�)d�Z<s�R����������U���*���;��zƕ�l ��A2����h��R�)4B�i.<�t&A��1P���f�e���,���p���  �  Ub�O�i�!dm���n�B�n�W{m�ϭi�"b���U�1E�@�1��A� ����q���@��Y���"��6�7�I���Y�/e���k�?o�{cp��6p�}�n�(j���a���T��{C���/�"������Y��������@��\'��Q;�]N�N@]�^�g���m���p�Bzq��q���n��i���`�\�R�;A�0-��K��g����΂�
�G�	�*���>�y�P�V5_�e�h�A#n��pp�_�p��Gp�=�m��1h�T^��O��=�5�)�¾�S)
�@s�`���5�����1��F��HX��ef���o���t��w���w���v��)t��n�̡c���T��B���.������76�����s���(���<���P��[b��o���w�]N|��~��`~�zQ}��z��Ks���g�i3X��OE�6�1�5!�ƣ������5J!�N�2���F�iZ�2Fk���w� >�����L��lU��ܩ��P���x�.l�(�[��tH��J5��2%����(����V*��B<�K�P�d�"<t�����_�����n���w���턾܂�J�}�� q��%`���L��;:��
+���!�c� ��L'�5�4�OG�.t[�UWn�I�}����|��y���݈�b���փ�������Z��%�r���`�L�L���9���*�{"�� "�)���7�YJ�\@^�Rp�r�~�H������,���y���&��t醾����U~�b�o��V]�sI��7�()�g"��#�D�+��;��)N��b�S�s�����?<��h���M���舾�{������􃾭@}�x�m��&[�SG���5��(� �"�]2%��E/�Z?�T�R�C�f��w��V���r��y���)w��4���9
��Dc��:�6v|�{ul�rOY��E��r4���(��+$���'�D3�Q�C���W��.k�C�{��  �  �^B��~Q�|�`���o��1~�W��JZ�����y���'r�|�Y�k�@�H�*�78�� �T���B/�	vF��&`���w�cv��m�������ߐ��;�|�m�m���^�hP�i�@�1�ߏ ����7� �+��ܽ�rٽE��\���BY	�֐�/_*��:�)J��Y�h h��)w�}��������ˉ�c����݀��l�}lS���:�6�&�_p�#����$���7��fP���i� u��솾����g����eOx��Qi�LZ��bK��<�7,����A{�����[Gݽ=�߽i��7��2Q�zl#�i�4��
E�,�T��c�?/s����䱇����팾HS��zR��3l� �R���;�#�*�dJ#���&���4���J�g@d��W}�����
����菾�!������i���q�wc�0T�X�D�̲4��F$���?�p_��-���������V����%�77�o�G�P�W�b%g�Bv������ �����tO��µ�������J����p���W�]�A�2�3��#0�nK7�.H���_���y�kֈ�W�������ߕ�����ǋ�(���U3z���k�p�\��LM�a(=�g-�w�Q�K�����Ƴ�g��8)�ƣ9���J��Z��pj��ny��6�� ���癒���Aƙ�0���-����*��bs��/Z�/FF�L�:�MJ:��nD�qyW���o�먄�B���l�Lv���֗�7풾� �����*Pz��dk�k\���K�2A;�n�*�v��Z�1�����f����*�.�Ca?��P��`�Z_o�k\~�����-�����j���Ι��������������k�T�ƺB���:�>���K�B�`��Sz�����Xe���1���j��ؕ��*둾CЊ��Q���w�P�h��KY���H�H8�g�(��q����5f��&�Ʉ�AZ'��
7���G��gX��  �  ��/��3G���a�N1~�TT�����������`��rD��v�����9f�E�I���6�O|1��B:���O���m�Os���C���m��[��Ԡ�ɗ�S���Py�B4]��C�^�,��%�ũ�!��x�׽��Ľb�����'E����ν3��U
���~$��9��HR�q�m�k/���������������6��~0���~���]��D��j5�Y�4�P�A��Z��@z��d��⚾��91���Ğ�(�����j:p��T��<�΁&������Kv齱�ҽ3ý����/!ɽ0Fܽ�"���
��v���0�Z>G���`��}�8��@C��h���q���\���
���э��{�Q�\�B�F���<��FA��5S��`o�9F��t1���U��De��9|���>���y��Ls��,\t���Y�|\B���-�a��5�����"X�яܽ�pؽ�vݽ 3�8C ���a7��0��TE���\�fYw����(=���~��b����d���^��a&��8㎾�A}�a���N�b�I���R�h�h�B���W>��
:��늭�CP��Z,��R6���y��/9��/�x��_�"�H�dH5�C3$��g��>	�] �N�������������8���!���1�E�D�8Z�9�r��憾1K��j
�����������������܎��}���c���T��T�Ha�Vz��⌾v+�������Ʋ����Ϫ�����g�������t�{\��jF��_3�b�"�g$�׀�` �q�������.���	��r�=�&��7�.�K���a�[{�����u���B���尾�촾�������R��)����#u���^�xT�x�X�,j�~�T����������� ��/���^栾�ڒ�'�����n�.�V��JB��0�� �W�����>�����_� ��[���� ���.�t	A��  �  8�'��RG�4`l�����g4�����������F0��`_���<��ą�Ch�½P�v�I�N�T��bo��p�����Be��ԥ���@��枻�����z��v͆�Jme���A�ӗ#�
+��j���нr޹�⩽����x���P��}]��8xƽ��὾~�j��SP4�_�U�(I|��ߒ��֦�l��Y|����,���{���e���]����`�1XN��TM��]��|����kG��x궾�j��"���nI����6��� 0��f\Y�0k7��O�a���彏Cʽ"���.������e\������
��z�ֽG\���1��&��bD���g�S��~�������_���ž<�¾6����᥾����Z>}�Z�a�ARU��Z���p��䉾���:?��~����ǾvQžnA��������.8�� [�X#;��!��>������߽�ͽ�ý�忽m(Ľ%�Ͻ�F⽸������Xh#��^=�+]�R��������y����Ⱦ �˾�KƾV���D��� H��}g��qh�S�a��,m����	���̫�EQ��V�ʾvξ��Ⱦd���w���
[��Z���']�9[?�D'��2�Oc�@���u�形�ݽ�ܽ�㽹L�>��B����"��8�n�T��u��E��F���涾�Ǿpsо8�о}`Ⱦ�Q���4���%��j��|�m�_�l��2}�%��Iơ�=���ƾ�=о"�оO-Ⱦg���餾�(��oQy��ZW�6.;�xx$��v�>y��9��M����>὆D����0����'�)�ڃA�C_�8+��"���멾<��PI˾��Ѿ�sϾ�!ľ[���۝��Ǌ���y���l���q�Vރ�T'��\���&����˾fuҾF�Ͼ�ľ�r���������[�o��O���5�� ����=�k.��������Yp�s)�|����I5���3��  �  �s&�	�L�i�z�o떾⠰�oǾ�6־�7۾��Ծw�ľ�����Ǖ�u߀�Zf�"P^�Ek��*���A������Jɾ�׾e�۾�5Ծ<+þ�ȫ�鑾c�q��zE��� �IV��Oݽ�t���禽�!��3D��!���韽����ν����;��I5���]������ᠾ�Ṿ�@ξ�Kھ�۾��Ѿ����ަ��;����x�r7c�@b��Fu�0Ō������:�Ͼf�ھp�ھ5�Ͼ�=��j��������b�i�8�������mӽ�붽���{�������є�� ���Q��[)ý��P��_#��gG��0s�!���͠��q�ľ��־ld߾��ܾ�ϾUݺ��Ȣ�#q���Jx���i�1p�����׀��;α��ɾ��ھK�S�޾��о�������i󇾛wa��l:��b������佛�˽�U��o���j���D�������"Ͻ��C��>X�B<��b��C���ҡ������Ѿn-ᾼ=�P �v�Ͼ-T��L������/	~��Uv���������˧�RQ���-־���;��k�ᾂ�оT?��Vs���z����`�a�<�h ���8�����n�ӽ��̽qN̽�:ҽ�޽5x�2N���+4��DU��D~�������@�ɾ�B޾TA��i�7j�Vtξ%���n����[�������`������#Գ���˾ ~߾����]�߾(̾8��L���`I��!�X���6����{
	����0�ό4սɄϽ(Sн��׽��j����M�le"�U>��b�<ˆ���������{�Ѿ���Z3쾡��@WܾsPǾ�������- ��z���A����m��Ǥ��弾�Ծ<M�n��=�۾�kž����W���1v�vO�:�/���P�X6�f���׽7Խx�׽�!���B��~��-��  �  ��'��R�+B��
-��Q��x�־��羿��|�澈�Ծ y������r�����t���k���y��E�� ���U���T�پ���8�|�徵AҾ����Xe���|�|%J��I!�ˬ��ԽIX��t����<��φ�>����f��MÕ��è��:Ž���u���7���e�`�;L��դǾ�޾hw������6�;�}���P���f���'q���o���������f��M�ʾ���-,�D�o��Zʾ�[�����j��;��D��M���ɽ˶������,N��)Ή��z���^���!������-ڽ�,��K#�Y�K�s�|�ͬ���4���cӾZ�����h&�B���Cɾ3���Eʕ�����tw�E~�km��������ؾ�:쾣���R������	Ⱦ�2���/��'�g�&<���������ڽp���zI��fz����������#�Ľi�޽s��;;�P+=��`h�"%������;Ⱦ�����������F�߾��ƾ0��*7���=�������(������:���cξ/�������8�����[�߾;.ž_����p�e��=�����E�:׽�ɽi@ý"�½�{ȽE�Խ�软�������2�(�W��������c��h�׾���>l��=�������ݾ�Kþq��)��%S��/����J�� W��'���ھ$���������o��sCھrL���栾�r����[��6��V�m]��9뽾q׽�y˽�$ƽ3�ƽ��ͽ�۽�|�}���|�"<>��)f�o����ħ��8ž�V�����ɟ������Ȳվ�Ӻ�-졾纏�l����Ɗ�i䘾rd��ʾ>��e����n��F'��	�^yҾ����������|��P��
.�8��g�k��o�׽[]ν�'˽f�ͽ� ׽z��K ��l��+��  �  �T(��U�X�����������#gܾ�f�#g���$�Xھ[I��މ��u�����y�6�p�k?���>Ȫ��ƾc�߾�L�E���7���׾@��O������: L�
�!��	�BҽCC���d�����Hƃ������N��펒�����d½)�뽏����8�(�h������$����̾�����_�����
HӾ�����䜾�A���v�O�t�Y��,���ɴ��Rо�����󾧳󾫶�~�Ͼ�W��괓�)@n��\=�4K�����ƽX����[���9���҆��{��wC��������׽�t�q�#�MSM��N������u����ؾ~ ��{������c~澿fξK������p���A|�줁��j���ߧ��þ�|޾Y��u��W���k�g�̾4Ů�N���4~j���<�9�]s����׽VK�����j��H��T���4���������۽� ������=���j��c��������̾�U��]���m��B����d�˾I�� H��RɈ��Z��Xɋ�oԝ�PJ���gӾ���O��	� ��/��v���ɾ���آ����g��o=���Ny���齎�ӽF�ƽz1��Cؿ��]Ž^Nѽ��佖�� ���2��Y��|������?;���ܾ\���2~��>�w�������Ǿ���T���Ɗ�Z�����'ө�L�ľ5྿���������B���mi߾�G¾�������@]�h6�fs�@����|;ԽC^Ƚ�!ý��ý]�ʽxXؽl_�Ї����>�t�g��~��U̪�yyɾk�從������N1���4�ھX ��;���i�����;I���⛾>)����ξ�j��W��n��� �A��+@׾;/��O�79�ƋQ���-�) ��������Խ!L˽d'ȽA�ʽ�ӽ�B�9���~E��1+��  �  ��'��R�+B��
-��Q��x�־��羿��|�澈�Ծ y������r�����t���k���y��E�� ���U���T�پ���8�|�徵AҾ����Xe���|�|%J��I!�ˬ��ԽIX��t����<��φ�>����f��MÕ��è��:Ž���u���7���e�`�;L��դǾ�޾hw������6�;�}���P���f���'q���o���������f��M�ʾ���-,�D�o��Zʾ�[�����j��;��D��M���ɽʶ������+N��'Ή��z���^���!������-ڽ�,��K#�T�K�o�|�ˬ���4���cӾW�����f&�@���Cɾ2���Dʕ�����tw�E~�lm��������ؾ�:쾥���T��Ý��	Ⱦ�2���/��+�g�*<���������ڽt���|I��gz����
���	����Ľe�޽p��7;�L+=��`h� %������;Ⱦ����������D�߾��ƾ
0��*7���=�������(������:���cξ1�������8�����]�߾>.žb����t�e��=�����K�:׽ �ɽl@ý%�½�{ȽF�Խ�软�������2�(�W��������c��h�׾���>l��=�������ݾ�Kþq��)��%S��/����J�� W��'���ھ$���������o��sCھrL���栾�r����[��6��V�m]��9뽾q׽�y˽�$ƽ3�ƽ��ͽ�۽�|�}���|�"<>��)f�o����ħ��8ž�V�����ɟ������Ȳվ�Ӻ�-졾纏�l����Ɗ�i䘾rd��ʾ>��e����n��F'��	�^yҾ����������|��P��
.�8��g�k��o�׽[]ν�'˽f�ͽ� ׽z��K ��l��+��  �  �s&�	�L�i�z�o떾⠰�oǾ�6־�7۾��Ծw�ľ�����Ǖ�u߀�Zf�"P^�Ek��*���A������Jɾ�׾e�۾�5Ծ<+þ�ȫ�鑾c�q��zE��� �IV��Oݽ�t���禽�!��3D��!���韽����ν����;��I5���]������ᠾ�Ṿ�@ξ�Kھ�۾��Ѿ����ަ��;����x�r7c�@b��Fu�0Ō������:�Ͼf�ھp�ھ5�Ͼ�=��j��������b�i�8�������lӽ�붽���x�������є�� ���Q��Q)ý��J��_#��gG��0s����ɠ��m�ľ��־hd߾��ܾ�ϾSݺ��Ȣ�"q���Jx���i�2p�����؀��>α�ɾ��ھK�X�޾��о	�����n󇾣wa�m:��b������佢�˽�U��r���j���D�������"Ͻ��=��7X�:<�݋b��C���ҡ������Ѿi-Ᾰ=�L �s�Ͼ*T��	L������-	~��Uv���������˧�TQ���-־���?��o�ᾇ�оY?��[s���z���`�i�<�h ���8�����u�ӽ�̽uN̽�:ҽ�޽7x�2N���+4��DU��D~�������@�ɾ�B޾TA��i�7j�Vtξ%���n����[�������`������#Գ���˾ ~߾����]�߾(̾8��L���`I��!�X���6����{
	����0�ό4սɄϽ(Sн��׽��j����M�le"�U>��b�<ˆ���������{�Ѿ���Z3쾡��@WܾsPǾ�������- ��z���A����m��Ǥ��弾�Ծ<M�n��=�۾�kž����W���1v�vO�:�/���P�X6�f���׽7Խx�׽�!���B��~��-��  �  8�'��RG�4`l�����g4�����������F0��`_���<��ą�Ch�½P�v�I�N�T��bo��p�����Be��ԥ���@��枻�����z��v͆�Jme���A�ӗ#�
+��j���нr޹�⩽����x���P��}]��8xƽ��὾~�j��SP4�_�U�(I|��ߒ��֦�l��Y|����,���{���e���]����`�1XN��TM��]��|����kG��x궾�j��"���nI����6��� 0��f\Y�0k7��O�`��	�彍Cʽ"���.������^\������
��l�ֽ6\���1��&��bD���g�L��w�������_���ž7�¾2����᥾����V>}�X�a�@RU��Z���p��䉾	���>?�������Ǿ}QžuA��%�����48��,[�c#;��!��>������߽�ͽ�ý�忽j(Ľ�Ͻ�F⽬������Oh#��^=�]�K�� ������r����Ⱦ�˾�KƾQ���@����G��yg��qh�S�a��,m�������̫�JQ��[�ʾvξ��Ⱦk���~���[��Z���']�D[?�D'��2�Wc�L����彪�ݽ�ܽ��㽽L�?��C����"��8�n�T��u��E��F���涾�Ǿosо8�о}`Ⱦ�Q���4���%��j��|�m�_�l��2}�%��Iơ�=���ƾ�=о"�оO-Ⱦg���餾�(��oQy��ZW�6.;�xx$��v�>y��9��M����>὆D����0����'�)�ڃA�C_�8+��"���멾<��PI˾��Ѿ�sϾ�!ľ[���۝��Ǌ���y���l���q�Vރ�T'��\���&����˾fuҾF�Ͼ�ľ�r���������[�o��O���5�� ����=�k.��������Yp�s)�|����I5���3��  �  ��/��3G���a�N1~�TT�����������`��rD��v�����9f�E�I���6�O|1��B:���O���m�Os���C���m��[��Ԡ�ɗ�S���Py�B4]��C�^�,��%�ũ�!��x�׽��Ľb�����'E����ν3��U
���~$��9��HR�q�m�k/���������������6��~0���~���]��D��j5�Y�4�P�A��Z��@z��d��⚾��91���Ğ�(�����k:p��T��<�΁&������Hv齭�ҽ�2ý�����#!ɽ!Fܽt"��ڧ
��v���0�L>G���`��}�0��8C��`���j���\���
���э��{�L�\�?�F���<��FA��5S��`o�=F��y1���U��Je��@|���>���y��Us��;\t���Y��\B���-�k��=�����+X�Տܽ�pؽ�vݽ�2�3C ���W7��0��TE���\�WYw�	��� =���~��[����d���^��[&��4㎾�A}�a���N�b�I���R�m�h�E���[>��:��񊭾JP��a,��Z6���y��79��?�x�_�/�H�pH5�N3$��g��>	�] �X�������������:���!���1�E�D�8Z�9�r��憾1K��j
�����������������܎��}���c���T��T�Ha�Vz��⌾v+�������Ʋ����Ϫ�����g�������t�{\��jF��_3�b�"�g$�׀�` �q�������.���	��r�=�&��7�.�K���a�[{�����u���B���尾�촾�������R��)����#u���^�xT�x�X�,j�~�T����������� ��/���^栾�ڒ�'�����n�.�V��JB��0�� �W�����>�����_� ��[���� ���.�t	A��  �  �^B��~Q�|�`���o��1~�W��JZ�����y���'r�|�Y�k�@�H�*�78�� �T���B/�	vF��&`���w�cv��m�������ߐ��;�|�m�m���^�hP�i�@�1�ߏ ����7� �+��ܽ�rٽE��\���BY	�֐�/_*��:�)J��Y�h h��)w�}��������ˉ�c����݀��l�}lS���:�6�&�_p�#����$���7��fP���i� u��솾����g����eOx��Qi�LZ��bK��<�6,����?{������RGݽ3�߽\��/��(Q�nl#�\�4��
E��T��c�-/s����۱�����팾AS��tR��)l���R���;� �*�cJ#���&���4���J�p@d��W}���������菾�!������i���q��c�0T�e�D�ײ4��F$���D�v_��.���������P����%�-7�b�G�A�W�R%g�	Bv������ �����kO�����������J��{�p���W�X�A�0�3��#0�pK7�$.H���_���y�qֈ�^�������ߕ����ȋ�1���g3z���k��\��LM�m(=�q-�w�X�Q�����ɳ�i��8)�ǣ9���J��Z��pj��ny��6�� ���癒���Aƙ�0���-����*��bs��/Z�/FF�L�:�MJ:��nD�qyW���o�먄�B���l�Lv���֗�7풾� �����*Pz��dk�k\���K�2A;�n�*�v��Z�1�����f����*�.�Ca?��P��`�Z_o�k\~�����-�����j���Ι��������������k�T�ƺB���:�>���K�B�`��Sz�����Xe���1���j��ؕ��*둾CЊ��Q���w�P�h��KY���H�H8�g�(��q����5f��&�Ʉ�AZ'��
7���G��gX��  �  Ub�O�i�!dm���n�B�n�W{m�ϭi�"b���U�1E�@�1��A� ����q���@��Y���"��6�7�I���Y�/e���k�?o�{cp��6p�}�n�(j���a���T��{C���/�"������Y��������@��\'��Q;�]N�N@]�^�g���m���p�Bzq��q���n��i���`�\�R�;A�0-��K��g����΂�
�G�	�*���>�z�P�V5_�e�h�A#n��pp�_�p��Gp�>�m��1h�T^��O��=�3�)����P)
�<s�Z���5������1��F��HX��ef���o���t��w���w���v��)t��n���c�t�T��B���.�|����76�����s���(��<���P��[b��o���w�oN|��~��`~��Q}��z��Ks���g�u3X��OE�=�1�;!�ɣ������1J!�G�2��F�iZ�$Fk���w�>�����	L��cU��ө��?���x� l��[��tH��J5��2%����(����V*��B<�U�P�d�0<t����`�����w�������턾!܂�Z�}�� q��%`���L��;:��
+���!�h� ��L'�8�4�OG�/t[�VWn�I�}����|��y���݈�b���փ�������Z��$�r���`�L�L���9���*�{"�� "�)���7�YJ�\@^�Rp�r�~�H������,���y���&��t醾����U~�b�o��V]�sI��7�()�g"��#�D�+��;��)N��b�S�s�����?<��h���M���舾�{������􃾭@}�x�m��&[�SG���5��(� �"�]2%��E/�Z?�T�R�C�f��w��V���r��y���)w��4���9
��Dc��:�6v|�{ul�rOY��E��r4���(��+$���'�D3�Q�C���W��.k�C�{��  �  �����������\}�[�n���_��	Q��	B��d2�m�!��O��������ڽ�dֽ�ݽ�F�V��K���b&���6�mF��}U��d���s�G󀾜���ED��X܇�������o�W�U�=���(�s�d���2"��	4���K���e��C|�5��E���ß��;-���5{�\_l��X]�DnN�5?�E7/������ߡ���8�H�۽:۽a*潈������p�b-�5#=�W^L�
<[��2j�;y� A�����wo��灆�1~�$Ih�;O�M7�q�$�
���B�=�)�Ty>�	X�e�q�G���YJ���p���W���#���|��m���^�}P���@���0�um ����io�r��n���^v �C������-���>���N� @^�=]m��|�ڪ����Wя��h�������'gn�,U���>�q4/��)�\�.�hT>�2U�Uo�ă��+��QR���Ⓘ��������Z���u�+�f��X�r�H��^8�`(������~G��j����0�1�_/��@��?Q��a�5Qp�#}��[�����->�����[Ε����>C��%?t�x�[� 3G���:���8��A���S�Y�k��Ⴞ�I��E��ř��ј�Y��k����F���m}��hn��_� O�{:>�Z�-�i��G���d����B�O�+�<�m�L��\�k"l�f{�k������DG�����z��	����������n�tV�|�C�@G:���;�joG��[�¹t��iW���ߗ�Lי�񚗾�M��?X���܃���x���i�}Z�$FJ��9�)�l���E�~�����B�Kr#��2���C�K)T�)d�Z<s�R����������U���*���;��zƕ�l ��A2����h��R�)4B�i.<�t&A��1P���f�e���,���p���  �  �2��!���ޘ����%�|�#J`�u2F�G/�:���	�f�򽙞ؽ4�Ľ�����'���ݺ�Y&ɽ��޽.���؅�� ���4���L�H�g��A��fM��{����	��.���z���E��Dx��rbb��+G��m6��H3��T>�2�U���t�缊�,��������:���b��(��F�u���Y��@��[*���������\<սt�ýT��Շ��#����ҽXJ�߸�&��¹'� �=��FV�!�q�fM����������&��˂��b��}o���^x��$Y�y7A��!5�667�'G��b�[���+ޑ�1�6��&���PU��58���t���Jr�ocW�6h?�5l*��	�P��.���0'߽Pѽ�z˽}Ͻ�g۽����������&��L;�\R�Mal��c���Ò�=����_���^���|��i-���b��j|��^�E~J�  C���I�8�]��!{�TC��!��������魾�ܫ�����ki��{9���v�-\�s!E�Q1�q���*\����;�X���9��Y������"�O�'�b|:�ЯO�&�g��[���ˏ�睾/����ְ�������ì��=!������e�S?U���R���]�cu��O���ܚ����6O���Ǵ�Yo������bL��Lڊ�)�y�р`�->J�;�6�Um%�st��3
�yY�k��|���* ����خ��L#�94��lG�G]��"v�%����N��"ˤ�*'���6������!���e������x��q`�3�S��U�Ze��t�$鏾V���0Ǭ�	ҳ�h��������c��Ɏ���1��aq�eDY�zD�P~1�J!����
��� ������o���{�p*���%�*�S<�wnP��Tg�ݟ��sˎ�o'���᩾c���쪵�^���}K���_��j懾-r���]��U�d\��o�uU���ږ��-���I���  �  Ɍ��j��������^��� kj���E��&��s�3x򽌰ҽ;w��!W��?O������<���$������?ڽW��3{��+.�6�N�q}t�ᎾY/���B������2�����~'������3����d�u�O�~�K��Y��Rv�}z������v����y��U����h��]ӫ�a����ڃ��`��'=�I ��i��K�R�ͽ����"���=���Ǡ�٭��˼����ʽ�2罧�����>69��o[�ON����������Ҹ����������[���ϐ���z���\���M�>!P���c�M�������P��YO��4�þ�¾n�������ɔ�U/���:Z�Oa9��]����+���ս��½�4���ݲ��ﵽ�P����ѽ>@����/��C2�q�P�6>u�B䎾靣��$���\þ�Ⱦ��ľ]&��ť�L`��a'~���d�a[���c��T|�&j��E,��|Y����ž@˾�2Ǿ�躾�𨾻l�������[���<��#�Ũ�} ����z8ؽJϽ-"ͽ}�ҽ�k߽95��	�L���-���H��i�伇�l��eɰ�Q���L�̾�+ϾYKȾ����:3��,��?|��q�n��!k��(y�� ������Z"���ľ#�Ͼ*�Ѿ7�ʾ���¨�`����� &]�a�?�:5(�]\����)��"�F���߽���C�������.�1t%��y<�X�X�+N{��G�����X���Q�Ⱦ��о� о�ƾ7��u������l|�˥l�Ȭn�&ꀾ�Q��|�� y��y/ɾ�OѾj<оdƾV(䡾�<��;t�'AS��8�X;"����������W�N$��U���My��8�ծ�І.��aG���e�����J��� ��4���:�;��Ҿ��ξ�B¾����W6������c�w�n��v�d#��{4��Rɭ�y���Kξ�  �  $�ھ�nվ��ž�7��򁕾�Ex���J��%�-����oH���V��Ga��p������*��r暽jЬ�ǽ�O뽝	���-���U�q@������m��P�ʾ��ؾ7�۾v�Ӿ����X�������[}�n�d��R`��ap��"���蟾�%���̾;�پ��۾ĄҾ�$���������j���?�0����3�ؽq~���3���}��ݖ���.��aA��1���]���qԽJZ������;��,e�����0ꤾ�`���оZ�ھ�=ھ��ξ�����m���.t��6b�ae�d�{���������u����rԾ�޾��ܾ�о�����������
b���9�H^�f� �mܽ�%½�i��0���W���(��X����ƾ�Z�ֽ�0���� �/��1U�o���J��"5��m˾�ܾ� �`�޾n�Ͼ�������3d����z���o�8qy��&�������Ͼ�߾N���4྄�о��[e��_����`�H;�$^�����콚wս�Gƽ�+��T���0����;ͽf�߽1���1��m�(�
�H�fp�Q���A����þ��ؾ=Y�\�����OоU��F���!�Q���������!��� ���OȾsݾK��B��ͼ�sUо76��j4���s��*�_�Xp<�B� �������]a���ֽ[�Ͻ�0Ͻ9Cս��st��5�	����wz8�n�Z���������﴾kn;�����S�}�޾��ʾ���Iq������@����ҁ����_��y*��t�Ͼ]Y����e���fݾ��Ⱦߛ��S˕��|�ߕS��3����j����b��)ֽ�ѽY�ӽ�ܽt��\�����'�AE��$j�,s��_���������վq��I�����پ�ľ�ӫ�����9��{ㅾ�#��
k�������3ؾI��  �  �}�P�"Zվ��������Ձ�0kP�&����v�ؽoM�����|g��_섽縂� ���Ґ��}��SD�����B]�ޡ/�R@\�ë�� ڥ�1�¾��ھԅ�()��zѾ驷����Z���s��n�n�����˫�Ŭƾ�ݾ����z��I�ξ�o������t�n�C��@�����ϽII�����񭍽F-��Dˆ���ݘ���� /˽������XT>���m�ނ���篾��˾�q��=�E��E�߾�hɾ.ʮ��H��Fс���o���r�M#��^�=i��w�о������Q��ɾ�������3ei�<��������ҽpӷ�G��!]����������1���S}����̽>��N�4{0��&Z��_�������W���ھ���~��ܫ�GྡȾ#O���b���ׄ�N[}�O����链7���F�ƾ��߾7���+�����-�E�ƾ�t�������Pf�R<���2�����(˽\Q������QX�����!/ý2�սd.����&�_J�#w��*��oe��1CоM��EV��'��<U�Y�߾�kƾ|%��eV�����ɹ�����P���'绾@�־e��r4���S��\���޾�þu������c��&<�-��������j"ڽ��̽h7ƽ�Ž��˽��׽�3�N.�+��&�7� ^��ن�a~��u��۾���4V��������>pپڿ���$������v����ӈ�5>����9�ľI)߾���8��|��-��L־չ�����˳����U�?�1��i��� ���A׽�̽�CȽ�ʽҽ/'�Ч��bl�qW%�ڔE�Io��ː��]����ʾ��4���/���F���Aa꾁Ҿ=#��4��[�����Q,���霾�r��u`Ͼ�W����  �  < ���$���V��=q���L��(�I����ս橽���c��C�%�.���#��� �&�ʏ3�o�J�azn���g���8����D1�KXV�}Oz����j����͗�d�������m���L��1�c� �qy���(��@��2_����*�������嗾*���B΄���g���B�q��}��Ɖʽ�Y��˲���y_��\C�2�Ț)��)���0�ߡ@�FD[�3���t.���ŽM������OI>��ac�l肾�@��/l��k��DP���ށ�Ec���C���+�~�,�!�ޜ1�(�L�|�m��%��D哾g���H���Đ��z����a��<��>��)��3�ɽ䶥�*֋��Dt�d�]��wQ�r�M�)�Q��^��[s�P��J���|½r�YE��=3���W���|�����3@������<��Zh��������f��JI�8�4�"-���3��H��e���������T���"���Kݝ�+ ��c��^_b�z�=����� ��Xֽ����������.<�����!���a��eꋽ�O��[ت�u+Ž$�0�q�)��#L�Vq� ���ę�KZ�����҆���唾�i��i�j�o�O�N@?�|r<��G���_���~����P������������[Ԕ��ヾ�b���>�V�������z�ý����qz����My��'2���薽����OV���p��3ݽ��V�o:���]�"����͒��)���U�������.������y_���%c�L�J��&>���?��iO�<�i��;���?��̼��J��|���
	������{�{���V��#4��T�����/fؽ���ݞ������ᴘ������5���}���[��*��̽������@'�H�l�l�ʾ��*������Q��Ng��My�����@iz�c�\���G���?�WSF��Z��Cw�/��ac������  �  t"��xm�������k���H��b%��g��ս"�������Pg�I2G���2���'�\%��0*���7��N��Ir��[��wӴ���)F��S.���Q��t�~����͑�*�k����;���h��aH���-�~v�eb��3%�]�;��Z�b�y�释�/Ғ�����̭����b��-?����r��Vʽd��o���c�݌G��26�;�-��"-�"�4���D�"\_�xt��IS��K Ž0��������:���^�ֱ�ݰ��m���Q=��^����v}�=^�0�?�@(��f�j���-��<H�>h�烾z?��񌖾b}���L����1]�ǰ9��v�����T�ɽ��������ix���a��U�-�Q��U�K*b���w�����D(����½��콯�5�0���S��{w��j��N����5��w��n����ƀ�	�a��PE��l1�*���0�+D�T�`�k����z����ĝ��&��yя�$����V^��2;��P�� ��	׽���x���休�gN��w��������h�������`��������ƽ������(��1I��l��܇��X��8����ࡾU֜�V�������4f���K�<�]X9��{D�g[���y�V쌾z����ڢ�������������f���_�̅<����}���vrŽ���*���6ҙ��}���5����������a���9½�/޽���to��_8���Z��N~�񽏾���������"��ƚ������}}��^�%;G�k;�V�<��K���e��|���������\(���碾ɐ��X����Vw��S�,[2�0�����ҹٽ�ֿ�����3����������L<������Us����6tνb��k����%���E���h��������ݠ�t��á�����F����u�d�X��nD��<�7C��*V�wr��C�������P���  �  NU��/����w���\���=����b3Խ�����!��c(t�ĽT���?��a4�Q\1�#�6���D���\��%�%{���<����P@	���&��CF���d�}~�;N��/$�� \��$�s��5X��o;��G#�Xa�U��o�	0���K�*�h�P����"��UR��'��'r�GMU�q�5���f����˽e���n��+�p��U�RC�C:�E�9�A��;R�1�l�H�������%ƽo������1��Q�V�n�|҂�{鈾̄��}���5�k�]9O�#�3��W�����x�L�#�x�;���X�A�u���7Ƌ�튾����
o��Q�֌1���;����˽�����G����Go�+Hb�G^�WYb�
1o�)���򚒽g֨��bƽ׉�5�jQ*�ĕI�=i�Yt���V��Mk��㍾4C����p�!T��
:�-�'�^Q!��h'�4)9�JES���p�텾�r�������ԏ�~����r�K�S�k[4����$ �1ڽ�
������q���َ�։��$��R���"���} ���#����˽����
�)�#��{A�T@a�a
��X匾���"��z{���I���`u��Y��eA�N�2�Z�0�֮:��O�WFk�8��(����)���\������/��!Iu���U���6�����(�	��}p˽o^���K��EF��<����h���b���ŧ���?YȽ���>������.3��Q�"<q�&T��Ṓ�ј�mh��f�������!�n�5�R��H=�C22��3�`mA���X��u�ڈ��ԓ�%_���U�����������(k��K���-��[�����޽�-ƽ@v���c�����k+���|��X��P6��i����%Խ�$�:m��#�H1?�la^��}�oˌ�E����������9U��fW����g��]M�.�:�"�3���9��$K���d��
���l��6ϗ��  �  �xq�_�l�.^�D�H�p}/�:O�l�����ֽ�2���ț��䆽{n���W�(�J�1G�3HM�!]�
v��E�����	���1!ήF����6��MO�2�c�a�p�ps���j�*�X��@�$=(�q������[�V��у�U6��N� #d��;q���s�pk��Z���B��y)�����P����Ͻ8J��,����Y��k�m��8Z��O�gPO��mX���j�oI������~歽�˽>H����rR&���?�DhW���i��s�e�q�Rf�y�Q��^9�]�!���^_����P���(�1B���Z��#n��Vx���w�P>l���X�T�@��['�����l��%�ҽӶ�˲���Ϗ�uɃ���x�	�s�_x��R�����n��殴�VJϽ��ｚ����"�-�;�G^U���k��|{��ڀ�  }�#n�0X�0y?�@)�J���,�1v���(�9?���X�b�o��*���c����3�s�n0^�9>E�9",��*��~�_��?�Ƚ�\��� ��j����㔽��◽�����ԭ��ɿ�*�ֽO�|���@�7���Q�elj��R��o��kb���Ju�V	^���E�v�1�t<%��:#��,���=��U���n���������鉾h����z���b��aI�r�0��d���	o��׽<Ľ#���oӫ�,���GK���ت�<������ֺԽ9���Y�l���s-���E�{�_��,w�"����s���׈�����cq���X�u�@�g.�B�$��+&���1�pF��^���v�=߄�N���m,���`���s��Z�%]A�dg)��q�����w齩�ҽ�C������g�����􁪽rӰ�sǻ��j˽��^��s)�	� �(�7�2�P�Cj��4�����/��֬���$��sl�5S��<���,��&��+���:���P��i�nj��̃���  �  �ZN�`L��cB�&�3�W"�jd������7�ǽ�P���国S֊�E�{�z�k�"bg��o�3����2��qY��7�����ν�O�[���[�'�˹8�w�F�4O�ۺO�H��#9���%����� ���콸�������	�����O1�|�B�`�M�*Q�1L�`y@��m0�G���%��*��<�ݽ�Ľ.���<��*��
;}��p�y�o��{�#���ꗽ�������[ڽCL��L�
��V�\+.��>���J���P���N��eD���3���������.�����b�� u'���;���K�`	U���U�T�N�YsA��0�	��'���\���ʽEе��.��Yu���y���������)��p����T���Wɽ�5���������op/�24A���P��D[���^���Y��lM�Xe;��^'�tY����f�b��DI���'��n<�*�O�Xv]��c���a�� X��:I���7�w9&����l
�����8ݽ�[ɽ��²���|���������v򲽰���7�Խ=�������W:�mg0�f{B���S��b�Q�j�&�k��8d�A�U�-�B��'/����P���I�~�.)�â<�,!Q���b�`�m�7q��=l�t~`��dP�ɉ>���,�^���h�������ؽ��ȽGS�����������-��E$ǽG�ֽ˼齦���1��<����*�
�;��M��J^�Z�j�p�p��\n��d�(<S�2 ?�%�+� ��}�����ɕ�Q�/�JD���W��xg��)p�A�p��)i���[���J�C9�(�'������
�N�����Y�ս�+ǽ�l��7���	����½�kϽZ�m���>�U%���!��w2�mAD���U�pae���o�v<s�Ln���a��OO�� ;��(�����	����5'�E<9�īM���`�� n��  �  ��,���-���)���"�[��#l�����#��P���Iн�ͺ��}Җ����۫��~����������*���n�ֽ���J ��#
����-f��.&�=�,�C�/�^�-�~;&����LE
�����i�ڽإʽ��ǽ�\ҽ���v������!���+�5k0�ע/��w*�n�"��C�_������l0㽉~ͽ�/���,��-���M������S��	'��������ʽ~t�l�����dV���c6!�f)�� /�9j0��,��7#����T��N���ֽ��˽>ν�޽����r��]��|U*�3�o26��4�	.�o�%�Do�����u	��(��Kw�_cս\��Oo��`Ĥ�Q���1���­�R]����ҽ�G�����Ht
�V���p�#+(��d1��
9�
�=�]g=���7��-�������� �,s��j��,����� �_�/�q;��-B�%TC���?��8���/�VC&������	��1���A�=ս�Žv����������~u̽
�޽����D�L����r�$��.��Y8�gGA��*H�SeK�=�I��^B�M6�bB'�%���B����H���>�^���#�{R3�%�A�X�K�<rP�˪O��xJ�uB�p&9��}/��%�C���'�n=�u��a��W\ս�9ͽ&�̽��ӽ;���b�����O��I,��3$���-�^�7���@�N I���N��$P��3L�}�B�L5�%����C3
��;�P�Á�lH��)�	�8���E�5&N��P���N�6MH��?��h6�P�,��&#���`��q�����o�òԽO:Ͻ��ѽ%Q۽z&�
���X
��9�*����)��Y3�c�<�q)F�U�M�J.R���Q�+L�G-A��p2� q"�z"��3
��w���	��Q'!��B1�Pl@��L��  �  ,�g��������������D��*��-	�����L�܁˽|������W�����GK��j�ѽ�뽬�����d5�����|�x]�/��+{����Y������hʽo��,P�����\0���<���bؽH��|��и������q��X��dE���ND�O+��)��p��/%�RȽ9��)]��~����T���zŽ�!ݽ^l��a�����~��/����-R����L���#�Ơ��G�,i��G�ܽ�Ž8���xG��e_���sϽue�v]�S6����'��B� �[I"���"�eK"��_ �M��w�����& �����ѽ�½����6X����̽�S⽠����
�i6���Ƞ$�V�'��7)��|)���(��s&���!�s���}�������t۽&ͽ�GȽ��ͽ��ܽ!+󽞃��D��6��e&�4�+�#y.�|�/���/�'�.�[4,�<:'��h�����������O�ivؽSսE�ܽ��u�~+�����I&�m .�~�2��a5��j6�&q6��Z5�\�2�<-�%�n�lZ���������a��*�@�����Q����$�:�.�M�5�4�9���;�r�<��$<�I�:�z�6���0���'�5�΀�i������`轻����T����i;&���/�� 6�F�9�˂;��;��};���9�K�5��C/�V�%�/��q��������	꽞N��7b�7���?�c�(�J�1�M�7�e�:��<�	�<��><��0:�-�5�b�.��%��b���-�`����U������L��� �ř �;�+�d4���9���<�->�#D>��q=�L;��q6�	�.�Ы$��~����0���L{�>�)M ������U $�m�.��  �  U6����ͻ��X�X#��*�pD.�� -�qq&�`��-��OA��3�۽6�ɽ��Ľ�ͽ���L������h��G)�y�.���.�yw*���"�T��qK�F�������(�Ͻ���ү��.d��}@�������������vα�W�ƽ��ܽ5��J�������� �t�(��.���0���-��N%�]��T��x��}ؽbWʽ��ɽ�<ֽ�&�]o�yR�|�#�`�,��0�,�.�Y)�� ��`������O��"x߽Lʽ!��������喽�㐽4����/�����W��_�ֽ{r��� ��������s<)��P1�݃6�F7�)�2�̧(����q�
�����?��۽	�߽ ��)��N����&�yp3�v;�=-=��/:���3�M�*���!�B�xi��l����;�޽v8˽����\���묽�N������^ν\㽤���L��������f&��0��#9�^a@�g5D�V1C�ܭ<�c&1�jF"�ӧ��=��1��ŷ��������	�U��49)��E8�7mC�]BI��I��7E�I�=���4�,�+�#"�������/�%��F�c�ҽ)�ʽV�ɽ��нV,޽@��`�O$���}#�^�,�?�6�D�?��^H��vN�&�P��yM���D���7���'���I���}�2�l
��b�a�%���5�dGC�RlL��P��tN���H�rg@��7��u-���#����A8��`����i�m�ӽ�,ͽ�#νɲֽa������3���I��\�&��Y0��:��KC��<K��KP���P��L�5�A�n�3��#�M��f�	�����Y��>��-��<��H��[P��>R�7!O�weH���?�w>6�I�,�o�"�����-��d�Y��%�ὦEֽ�ҽ��ս���oK�S���������  �  �⽜W ��"��#��4�PC���L���N��rH���:���'��x����Uz�е�g�����U�
�,���>�XoK��P��hL���A��82�^� ����a���@�7lƽ臯�-���$#��0�}��o�%&m�%�v�g���c����/��E ���ս���e�a��h�+��b<���I�v�P��O���F���6�@#�R0�<S���j뽘s����ʲ �6�4�<E�� O��P�d�J�3�=�`F-�rc�3
�4���$�ؽ\���y�����f����~�M�u��*y�./�����RA��7����νZ�;X�D����%�4�7�#�G��hS�7X��T�׋I�_=8�-H$�w��9��P�����W�����2�&QF�sKU���\��#\�w�S�
�E���4���"�����I뽕Խ������� ���o������	�����(��(eĽ��ٽ�-�گ�g��j�&���8�UJ�Y-Y�m�b���d�h�^��Q��s>�p~*��/������
����j��v1��@F�y�X�L�e��aj�*�f��h\��M��;�!2*���+��!s��IM�|1սΗŽ?�����������
��t�ý�Yӽ�r潕���^�
�����[(���9��tK�,:\�'ei��jp�i�o��ef�egV�B���.���<^�L��x�Nd,��@��T���d��n��Rp��j��l]�M�L��
;�b�)�����������l�Hֽ��ƽM��"��Jַ�i���lʽ*�ڽx�b���~����]8.��?���Q�.�a�'m���q��<n���b�� Q�p�<��)��ڹ��D�W-#��n4��H�\��j��+r�:q���h�5}Z��PI���7�ǵ&�y���$
��w��݋���սt/ȽgR��8��������ǽս����x����	��  �  !�׽t �s��0���I�Y_���m���q�)Ck��Z��C�h�*�@$�������a	���l�0�(�I���_�t�n��r��cl�b\�i�E�B�,�1��/S����ӽ�<��Ě�Q����.o�fJZ�ūN�ĲL��T��e�"������O���Lƽ��r.
��^"���;�("T��g���r�!Ds�f i���U�|=�%��b�*�C�����P�"�?�:��S�/g��yr�Bs�O�h��\V�.�>���$�J���-�< ʽ�լ�ω�������(m�á\���U���X��{e���{������1�������۽s>������0���J�}�a�1�r�>�z��x�f�j���U�Y.=�p:&�Hi�� ��y��?�w�4��N�b f��w����j\}��]p���[�K+C���)�mr��[����ڽۿ�ϙ������f<��梈��ӆ��ё��H��Ai��Q|Ž��ud�.���$-� �F�*�_�8u��ȁ�N��D���f3q��fZ�9�A�z,�������!�ex2���I�}"c��y�,I������-p���w�
�`���G�9�.�{��ؗ��2��tӽ4���M[��rd���3���ԧ����z׾�Lѽ������ *��LB��[���s����*��o��]D��U>u���\��tD�\�0��z%�#�$���.���A���Y�wr�>�����D���A����u�: ^�1�D�0<,�������̟�B�ӽ����]������Kͦ�^p��;�)����Ž��ٽ������f42��K��d���{�FS��?���������V�n�o�U�%x>�:R-�_�%�ʯ(�6��HK�,d���{�����	����;��R�����p���W��>�p'�@������>轹zҽ����Wֵ������VC���_������ѽ`	�{	��  �  !�ս�9��  �sw?�#�^�rPy�`�����������T�v�$�[�/�>��f%���������*�2pE�Q�b�bh|�r���g������Ju��YY���9�T��{���н����ˎ�Ųs�
 V���B�?�8��7���=�]M�"�f�����#����ÿ��%�-�&�,�ϜL�9�j��u�������>��e��]hp��T���7�K� �`���������4�˺P�]Vm�vO���ӈ�kۈ��l���m���O�q50�4�9l�DĽ�����*����m���T�4F��*@��C�{�N�?�b�Ì�3������lo׽�������=��X]��)z�Ї�����^�������9o��kR�ߚ7�5�#�C4��,��(/�8/H�f�e�򵀾���8���h���Gi��Pq��yR��3��"������(ӽ󒴽�ݝ�gȍ��A����z��x�ٳ}�0���U�������{�����ؽ�A �=���5�o<U�lt�r���+��� �����o����cr�v�U�m�<�_,���'�!�/�MfC��s^�]�{�C
�����&��쑾`����'t���T�,6�˞�C�����7mǽ�E��T��𒜽�N��D���h��Ѥ���Ľ�޽�q������.���L��|l��C���T���`���
���(����~s�iW�g@�N�2��,2���=�I�S��p��V��<���z���K����-��/����~o���O�T�1�8H����G὿�ǽ���j���-���Lq~���S��C������nͽG�ʚ�l�n�8���W�yQw�����ᥔ�鹙�"8���i��o�
�j���O���;�[�2�e6��F�0�^��{�'����ٕ��W���4��'現� ���Kg���G��*���������ܽ��Ž����٩�uS������&��j|��p���Ľ��۽�����  �  ��ֽ����'�9�J�4�m�yޅ�����b���X��QǄ�,�k�yL�EN0�V��I���-!�}!6��wS���s������M��%ɓ�ߎ�G���r�g�RD��9!����нmm��[���df���H���5��3,�$�*�81�W@��Y��~�fؙ����5	�P��jD5�9Y���z�(!��>%��5�������F��Rec�8%D���*�E��g��d�(���@��_�S0�j��7���M���{<���4~���\��9�������½���#���@`�J�G�OS9�t�3�?�6�M�A���U��St��>��٥���
׽]D�U$��AG�k��ȅ�⑾O���>���č��-����`��HC���-�I�#�ON(���9��DU��xu���Vt���|��s���ǎ�9F����]��:����J���c�н�W���e������Py�eTn��k�_(q�7�~��㊽!������G�ս�� �RN���<�wK`����ϐ������m���y������V��pc�X�G�ќ5�y�0�mz9��N��rl�n��
ǔ��D���ᠾ����Ґ��&���_�B_<��\����N߽`�������6������u�����������L#��uW��UCٽ����i�Ɖ3��,U�F�x�$b��T��������У��\��N��bg����c�TCJ���;�_;�J�G�,.`�5	�XC��]���G��Y?������q����X|���X� �6�

�� �ʿܽ�X�����$��\9��񼕽�E���ښ�r⣽�O��ҁǽ���c�����>�<`a�����S������>y���ᢾ�J������
Ky��|[���E��;���?�v�P��k�@ԅ�<��� =���%�����WF��������r�UO�Ф.�4���\���׽�F��G���>�����_�,ݜ��颽`����9�� ֽ�����  �  ��׽�$���)�f�N�}s��4������u@�����'����q���P�W&4��9!����>�$�B':�}oX���y�3n��$��h���*�������ѷl���G�)�#�o2���нƍ��m^��Cdb�bnD�&�1��'(�ݝ&�}�,���;���T���z�����/ý����&x��p8�*�]��p���������ޗ��;��K���u�h�c�H���.������H9,��2E�}	e��Â����j���X��cǏ�)"��j�a��[<�<�1���
�½�㜽�=���/\��fC�8D5�!�/�)�2���=�kzQ��Rp�%���ᬭ��W׽Z�a�&��J�F'p�1�v�������V���I��x>����e��gG��1��'���+�_�=�;�Y�A!{�,c��w'��mY��zۛ��+��#��?b�}p=�[��M����н孽�y��I턽�'u�xCj�ٸg��m�F�z��Έ�/�����'DսB����T}?�id��x���%������K��.5���d��Q:��n�g��wK��8��3���<��R�0gq��m���=���������f����	��������b�?�>�������l޽K�󏪽Wj���퓽���������ꓽ�������ez����׽�g���$��b5�tXX��w}��W���}��9Ȧ�J��������;��\����g�6�M�W?�h+>��K��~d��,���n��#���+�����(����瑾+�����[�c�8����� ��۽����髽�,��P���@���ʘ��ʡ�J��U�ŽE����� ��@�Qe�����ו�\U��bS������UΝ�,���`~���_��H�L�>�E�B�uT��mp����
R����>���l������֊��Vw��2R��90�c_�q���Jֽ�Z��e2���)�������혽 ՚��ՠ�B���F����ԽZD���  �  ��ֽ����'�9�J�4�m�yޅ�����b���X��QǄ�,�k�yL�EN0�V��I���-!�}!6��wS���s������M��%ɓ�ߎ�G���r�g�RD��9!����нmm��[���df���H���5��3,�$�*�81�W@��Y��~�fؙ����5	�P��jD5�9Y���z�(!��>%��5�������F��Rec�8%D���*�E��g��d�(���@��_�S0�j��7���M���{<���4~���\��9�������½���"���@`�H�G�LS9�p�3�9�6�G�A�|�U��St�z>��ӥ���
׽ZD�U$��AG�k��ȅ�⑾M���>���č��-����`��HC���-�I�#�ON(���9��DU��xu���Xt���|��u���ǎ�;F����]�
�:����R���j�н�W���e�����Qy�hTn��k�](q�3�~��㊽!������A�ս�� �NN���<�sK`����ϐ������m���y������V��nc�W�G�М5�y�0�nz9��N��rl�n��ǔ��D���ᠾ����Ґ��&���_�F_<��\����N߽f�������;������x�����������L#��vW��VCٽ����i�Ɖ3��,U�F�x�$b��T��������У��\��N��bg����c�TCJ���;�_;�J�G�,.`�5	�XC��]���G��Y?������q����X|���X� �6�

�� �ʿܽ�X�����$��\9��񼕽�E���ښ�r⣽�O��ҁǽ���c�����>�<`a�����S������>y���ᢾ�J������
Ky��|[���E��;���?�v�P��k�@ԅ�<��� =���%�����WF��������r�UO�Ф.�4���\���׽�F��G���>�����_�,ݜ��颽`����9�� ֽ�����  �  !�ս�9��  �sw?�#�^�rPy�`�����������T�v�$�[�/�>��f%���������*�2pE�Q�b�bh|�r���g������Ju��YY���9�T��{���н����ˎ�Ųs�
 V���B�?�8��7���=�]M�"�f�����#����ÿ��%�-�&�,�ϜL�9�j��u�������>��e��]hp��T���7�K� �`���������4�˺P�]Vm�vO���ӈ�lۈ��l���m���O�q50�4�9l�DĽ�����*����m���T�.F��*@�|C�n�N�0�b�@̀�)��璲�^o׽������ۉ=��X]�y)z�Ї�����[�������4o��kR�ܚ7�3�#�B4��,��(/�;/H�j�e��������<���l���Ki��Xq��yR��3��"�����)ӽ�����ݝ�nȍ��A����z��x�ֳ}�,���O�������q�����ؽ�A �6���5�g<U�lt�n���'��������l����cr�r�U�j�<�~_,���'�"�/�OfC��s^�b�{�F
�����)��쑾e����'t���T�,6�Ҟ�J�����BmǽF��
T�������N��D���h��!Ѥ���Ľ�޽�q������.���L��|l��C���T���`���
���(����~s�iW�g@�N�2��,2���=�I�S��p��V��<���z���K����-��/����~o���O�T�1�8H����G὿�ǽ���j���-���Lq~���S��C������nͽG�ʚ�l�n�8���W�yQw�����ᥔ�鹙�"8���i��o�
�j���O���;�[�2�e6��F�0�^��{�'����ٕ��W���4��'現� ���Kg���G��*���������ܽ��Ž����٩�uS������&��j|��p���Ľ��۽�����  �  !�׽t �s��0���I�Y_���m���q�)Ck��Z��C�h�*�@$�������a	���l�0�(�I���_�t�n��r��cl�b\�i�E�B�,�1��/S����ӽ�<��Ě�Q����.o�fJZ�ūN�ĲL��T��e�"������O���Lƽ��r.
��^"���;�("T��g���r�!Ds�f i���U�|=�%��b�*�C�����P�"�?�:��S�/g��yr�Bs�O�h��\V�.�>���$�J���-�< ʽ�լ�͉�������(m���\���U���X��{e���{������1�������۽h>������0��J�q�a�&�r�4�z��x�^�j���U�T.=�l:&�Fi�� ��y��?�|�4��N�j f��w����u\}��]p���[�W+C���)�xr��[����ڽ#ۿ�ۙ������l<��颈��ӆ��ё��H��6i��C|Ž��ld�#���$-���F��_�8u��ȁ�I��?���^3q��fZ�5�A�z,��������!�hx2���I��"c��y�1I������3p���w��`���G�E�.�������2��tӽ4��&�V[��yd���3���ԧ����|׾�Lѽ������ *��LB��[���s����*��o��]D��U>u���\��tD�\�0��z%�#�$���.���A���Y�wr�>�����D���A����u�: ^�1�D�0<,�������̟�B�ӽ����]������Kͦ�^p��;�)����Ž��ٽ������f42��K��d���{�FS��?���������V�n�o�U�%x>�:R-�_�%�ʯ(�6��HK�,d���{�����	����;��R�����p���W��>�p'�@������>轹zҽ����Wֵ������VC���_������ѽ`	�{	��  �  �⽜W ��"��#��4�PC���L���N��rH���:���'��x����Uz�е�g�����U�
�,���>�XoK��P��hL���A��82�^� ����a���@�7lƽ臯�-���$#��0�}��o�%&m�%�v�g���c����/��E ���ս���e�a��h�+��b<���I�v�P��O���F���6�@#�R0�<S���k뽘s����ʲ �6�4�<E�� O��P�e�J�3�=�`F-�sc�3
�4���#�ؽ[���y�����f����~�?�u��*y�#/�����BA��%�����νB�.X�6����%�%�7��G��hS�7X���T�͋I�V=8�'H$�s��6��P�����W������2�/QF�}KU���\��#\���S��E���4���"�����_뽨Խ����(������o�����������(��eĽt�ٽ�-�ί�Z��\�&���8��TJ�J-Y�_�b���d�]�^��Q��s>�j~*�/������
����j��v1��@F���X�W�e��aj�8�f��h\�M��;�02*���7��8s��]M轍1սܗŽ?�����������
��x�ý�Yӽ�r潖���^�
�����[(���9��tK�,:\�'ei��jp�h�o��ef�egV�B���.���<^�L��x�Nd,��@��T���d��n��Rp��j��l]�M�L��
;�b�)�����������l�Hֽ��ƽM��"��Jַ�i���lʽ*�ڽx�b���~����]8.��?���Q�.�a�'m���q��<n���b�� Q�p�<��)��ڹ��D�W-#��n4��H�\��j��+r�:q���h�5}Z��PI���7�ǵ&�y���$
��w��݋���սt/ȽgR��8��������ǽս����x����	��  �  U6����ͻ��X�X#��*�pD.�� -�qq&�`��-��OA��3�۽6�ɽ��Ľ�ͽ���L������h��G)�y�.���.�yw*���"�T��qK�F�������(�Ͻ���ү��.d��}@�������������vα�W�ƽ��ܽ5��J�������� �t�(��.���0���-��N%�]��T��x��}ؽbWʽ��ɽ�<ֽ�&�]o�yR�|�#�`�,��0�,�.�Y)�� ��`������O��!x߽Jʽ��������喽�㐽*����/�����vW��J�ֽcr�����������c<)��P1�΃6�F7��2���(����j�
�����:��۽�߽��/��U����&��p3��;�L-=�0:���3�]�*���!�Q��i��l����M�޽�8˽����\���묽�N������^ν�[㽐���@��ل����~f&��0��#9�Na@�X5D�H1C�Э<�X&1�bF"�̧��=��1��ŷ��������	�[��<9)��E8�CmC�kBI���I��7E�Y�=���4�<�+�!#"��������/�8��F�p�ҽ4�ʽ^�ɽ��нZ,޽D��a�P$���}#�^�,�?�6�D�?��^H��vN�&�P��yM���D���7���'���I���}�2�l
��b�a�%���5�dGC�RlL��P��tN���H�rg@��7��u-���#����A8��`����i�m�ӽ�,ͽ�#νɲֽa������3���I��\�&��Y0��:��KC��<K��KP���P��L�5�A�n�3��#�M��f�	�����Y��>��-��<��H��[P��>R�7!O�weH���?�w>6�I�,�o�"�����-��d�Y��%�ὦEֽ�ҽ��ս���oK�S���������  �  ,�g��������������D��*��-	�����L�܁˽|������W�����GK��j�ѽ�뽬�����d5�����|�x]�/��+{����Y������hʽo��,P�����\0���<���bؽH��|��и������q��X��dE���ND�O+��)��p��/%�RȽ9��)]��~����T���zŽ�!ݽ^l��a�����~��/����-R����L���#�Ơ��G�*i��D�ܽ�Ž2���pG��Z_��ᗺ�cϽbe�j]�G6������2� �KI"���"�UK"��_ �M��w�����& �����ѽ�½����9X����̽�S⽰����
�u6�$��נ$�f�'��7)��|)���(��s&���!�����}�������t۽&ͽ�GȽ��ͽ��ܽ+󽖃��D��6�ue&�$�+�y.�k�/���/��.�L4,�-:'��h�������ؓ���O�dvؽSսI�ܽ��|��+�����I&�{ .���2��a5��j6�7q6��Z5�l�2�"<-�%�*n�vZ��������� b��*�D�����R����$�:�.�M�5�4�9���;�q�<��$<�I�:�z�6���0���'�5�΀�i������`轻����T����i;&���/�� 6�F�9�˂;��;��};���9�K�5��C/�V�%�/��q��������	꽞N��7b�7���?�c�(�J�1�M�7�e�:��<�	�<��><��0:�-�5�b�.��%��b���-�`����U������L��� �ř �;�+�d4���9���<�->�#D>��q=�L;��q6�	�.�Ы$��~����0���L{�>�)M ������U $�m�.��  �  ��,���-���)���"�[��#l�����#��P���Iн�ͺ��}Җ����۫��~����������*���n�ֽ���J ��#
����-f��.&�=�,�C�/�^�-�~;&����LE
�����i�ڽإʽ��ǽ�\ҽ���v������!���+�5k0�ע/��w*�n�"��C�_������l0㽉~ͽ�/���,��-���M������S��	'��������ʽ~t�l�����eV���c6!�f)�� /�9j0��,��7#����R��I���ֽ��˽u>ν�޽|���h��R��oU*��3�`26��4��.�^�%�4o�z���u	��(��6w�Ncս	\��Fo��[Ĥ�P���1���­�]]����ҽH����Ut
�e���p�3+(��d1��
9��=�kg=���7��-�������� �1s��f��,�|��� �U�/��p;��-B�TC��?�ބ8���/�GC&������	��1���A�0ս��Žq�����������u̽�޽����D�!L������$��.��Y8�xGA��*H�ceK�K�I��^B�&M6�lB'�-���B����M���>�`���#�|R3�&�A�Y�K�<rP�˪O��xJ�~uB�p&9��}/��%�C���'�n=�u��a��W\ս�9ͽ&�̽��ӽ;���b�����O��I,��3$���-�^�7���@�N I���N��$P��3L�}�B�L5�%����C3
��;�P�Á�lH��)�	�8���E�5&N��P���N�6MH��?��h6�P�,��&#���`��q�����o�òԽO:Ͻ��ѽ%Q۽z&�
���X
��9�*����)��Y3�c�<�q)F�U�M�J.R���Q�+L�G-A��p2� q"�z"��3
��w���	��Q'!��B1�Pl@��L��  �  �ZN�`L��cB�&�3�W"�jd������7�ǽ�P���国S֊�E�{�z�k�"bg��o�3����2��qY��7�����ν�O�[���[�'�˹8�w�F�4O�ۺO�H��#9���%����� ���콸�������	�����O1�|�B�`�M�*Q�1L�`y@��m0�G���%��*��<�ݽ�Ľ.���<��*��
;}��p�y�o��{�#���ꗽ�������[ڽCL��L�
��V�\+.��>���J���P���N��eD���3���������&��ｿ�[��u'���;���K�S	U���U�F�N�KsA��0�	�����F��ٲʽ6е�y.��Pu���y�����!����)��z����T���Wɽ	6ὗ������-��}p/�A4A���P��D[�˸^���Y��lM�`e;��^'�yY����f�`��@I���'��n<� �O�Mv]��c���a�� X��:I���7�h9&����`
����z8ݽ�[ɽ�𸽻����|�����ô��~򲽻���E�ԽO��������e:�{g0�t{B���S��b�_�j�3�k��8d�L�U�6�B��'/����U���I�~�.)�Ģ<�-!Q���b�`�m�7q��=l�t~`��dP�ɉ>���,�]���h�������ؽ��ȽGS�����������-��E$ǽG�ֽ˼齦���1��<����*�
�;��M��J^�Z�j�p�p��\n��d�(<S�2 ?�%�+� ��}�����ɕ�Q�/�JD���W��xg��)p�A�p��)i���[���J�C9�(�'������
�N�����Y�ս�+ǽ�l��7���	����½�kϽZ�m���>�U%���!��w2�mAD���U�pae���o�v<s�Ln���a��OO�� ;��(�����	����5'�E<9�īM���`�� n��  �  �xq�_�l�.^�D�H�p}/�:O�l�����ֽ�2���ț��䆽{n���W�(�J�1G�3HM�!]�
v��E�����	���1!ήF����6��MO�2�c�a�p�ps���j�*�X��@�$=(�q������[�V��у�U6��N� #d��;q���s�pk��Z���B��y)�����P����Ͻ8J��,����Y��k�m��8Z��O�gPO��mX���j�oI������~歽�˽?H����rR&���?�DhW���i��s�e�q�Rf�x�Q��^9�[�!���[_�~��P���(�*B���Z��#n��Vx���w�D>l���X�H�@��['�����l���ҽӶ������Ϗ�nɃ���x��s�_x��R�����"n������gJϽ��､��̷"�9�;�S^U��k��|{��ڀ�
 }�#n�7X�5y?�"@)�L���,�/v���(�9?���X�[�o��*���c����(�s�b0^�->E�-",��*��~�N��0�Ƚ�\��� ��d����㔽��◽�����ԭ��ɿ�9�ֽ'O����K�7�	�Q�qlj��W��#o��pb���Ju�^	^���E�{�1�x<%��:#��,���=��U���n���������鉾h����z���b��aI�r�0��d���	o��׽<Ľ#���oӫ�,���GK���ت�<������ֺԽ9���Y�l���s-���E�{�_��,w�"����s���׈�����cq���X�u�@�g.�B�$��+&���1�pF��^���v�=߄�N���m,���`���s��Z�%]A�dg)��q�����w齩�ҽ�C������g�����􁪽rӰ�sǻ��j˽��^��s)�	� �(�7�2�P�Cj��4�����/��֬���$��sl�5S��<���,��&��+���:���P��i�nj��̃���  �  NU��/����w���\���=����b3Խ�����!��c(t�ĽT���?��a4�Q\1�#�6���D���\��%�%{���<����P@	���&��CF���d�}~�;N��/$�� \��$�s��5X��o;��G#�Xa�U��o�	0���K�*�h�P����"��UR��'��'r�GMU�q�5���f����˽e���n��+�p��U�RC�C:�E�9�A��;R�1�l�H�������%ƽo������1��Q�V�n�|҂�{鈾̄��}���5�k�\9O�"�3��W�����x�I�#�t�;���X�;�u���4Ƌ�튾����o��Q�Ό1����:��x�˽�������A����Go�&Hb�E^�ZYb�1o�.�������q֨��bƽ��=�rQ*�͕I�Fi�^t���V��Qk��㍾7C����p�$T��
:�.�'�_Q!��h'�2)9�FES���p�텾�r�������ԏ�z����r�B�S�c[4����$ ��0ڽ�
������k���{َ�}։��$��T���&���� ���#����˽����
�0�#��{A�\@a�f
��]匾���&��~{���I���`u��Y��eA�Q�2�\�0�خ:��O�XFk�8��(����)���\������/��!Iu���U���6�����(�	��}p˽o^���K��EF��<����h���b���ŧ���?YȽ���>������.3��Q�"<q�&T��Ṓ�ј�mh��f�������!�n�5�R��H=�C22��3�`mA���X��u�ڈ��ԓ�%_���U�����������(k��K���-��[�����޽�-ƽ@v���c�����k+���|��X��P6��i����%Խ�$�:m��#�H1?�la^��}�oˌ�E����������9U��fW����g��]M�.�:�"�3���9��$K���d��
���l��6ϗ��  �  t"��xm�������k���H��b%��g��ս"�������Pg�I2G���2���'�\%��0*���7��N��Ir��[��wӴ���)F��S.���Q��t�~����͑�*�k����;���h��aH���-�~v�eb��3%�]�;��Z�b�y�释�/Ғ�����̭����b��-?����r��Vʽd��o���c�݌G��26�;�-��"-�"�4���D�"\_�xt��IS��K Ž0��������:���^�ױ�ݰ��m���Q=��^����v}�<^�/�?�@(��f�j���-��<H�>h�烾x?������`}���L����1]�ð9��v�����N�ɽ��������ix���a��U�,�Q��U�O*b���w�����I(����½��콳�9�0���S��{w��j��P����5��w��o����ƀ��a��PE��l1�*���0�+D�R�`�i����z����ĝ��&��wя�"����V^��2;��P�� �}	׽���t���ἑ�eN��v��������h�������`��������ƽ������(�2I�"�l��܇��X��:����ࡾW֜�W�������7f���K�<�^X9��{D�g[���y�V쌾{����ڢ�������������f���_�̅<����}���vrŽ���*���6ҙ��}���5����������a���9½�/޽���to��_8���Z��N~�񽏾���������"��ƚ������}}��^�%;G�k;�V�<��K���e��|���������\(���碾ɐ��X����Vw��S�,[2�0�����ҹٽ�ֿ�����3����������L<������Us����6tνb��k����%���E���h��������ݠ�t��á�����F����u�d�X��nD��<�7C��*V�wr��C�������P���  �  �4��0�UH#�k���F����Ƚ-����z���C�Ç�������Ѽ2ʸ�<`��
��L���
���=�ܼ���%�%�LvR�c���+���f!ս��֨�Ns(�٣3��M6�0��""�Ɖ��.���s׽~Hý������̽X�轸���X7+��?5��6��A/�0 ����\뽒���e����p�i>�V��UG��(+ټ>�ü�$��V��������ռM)�������8��i�r���������t	�.�H�-��Y6��6��-��D��
�I���Dҽ2�ý0�ƽ@ڽ� ���b���$��4�(�;��:�5�0����H�
�>)齲��	���Rz�%M���,�S'�c�	�e���� �R�"[�)A��I/�6�M�I0w��
��G~���<�z����q>1�3?�9�D�D�A�616��%����, ��9G߽��罬
 ������%��58�DE�V�I��^E�}�8�$&��X�-q��X�˽י��uy���ut���W�A9E��:���4�X�4���9�˥C�	�S�ٍk�ɭ��ˠ��zk���$�7N����~�1��C�YO��R��!L�ѣ>�x,��t�"�	�Ť��E���M���'l&�+:���J�.�T�3mV�x�N���?���+�zK�7�����׽�������)؊�[{�^i�G^��"Y�L�X�&j]�bvg��*x�����3ۚ��i��+
ӽ�r���p�2�(�k�=��WM�\�U�AkU��WL�Dy<�)��D�����. �2�F�
��s���-���@�S�O���V�mZU�))K�:���$������i�ͽ�ޯ����KK����y���j��:b�h�^��`�Bg�P�s�����%���o��?q��m��H�JE�/z2�&�E���S�z2Y�w�U��AJ�{�8��>%��v���IN��9�����#��J7�lJI���U��  �  ��/���+�e��Q�Zu�u�Ž�]���z���D�"��/����(׼	��$x���,��ڳ�(�ļ�0⼝e��^'���R�兽����|�ѽ�����H�Rp$��9/���1�(�+��2�)�����ҽ�D�����E�Ƚ��㽀��-��E'��0��62��+����\	�������Yf��Up�RU?���e� ��s޼ �ȼ�6������|�ƼP(ۼ�\��j��U:���i��Y��JE���⽚��7p�H�)���1�1���(�փ����į�7�ͽ�����½"�ս�����: !�ƶ/��A7�&&6�,�,�d��&��r��漽Ե��xiz���N��F/����3T�]3��i�E��I��,����1�ޕO��4x����m����;߽z(�w���k-�t�:��A@�&=�42��o!�կ��r����㽱f۽ݪ�7J������j"�m+4���@�/E��A���4���"�W��wD�d5ʽ�%��鎽ov�uZ�X�G��<��c7��H7�x-<�f@F��RV���m�����|㝽}����$޽8���[�?R.���?�ƯJ���M���G�r�:�N)�Ѧ�<2�:�������%�� �nM#��v6���F��nP�#�Q���J��5<�Ӻ(�E)����\ֽ����8[��5򋽗�}��l��a���[�.P[���_��j���z�@㉽�����e���ѽp���vf�]&���9��*I�$RQ�=�P�0H���8��%�=����
r��:j��G����*���<��<K��^R�t�P�nG���6��9"�H��*s�/�̽Y���̙��{���<|��gm�+�d�xta��c���i� Mv�&ꄽ\-��0�k������<��6Z/��B�U=O�}�T��hQ�")F��E5��B"����\] ��+����� ���3��>E��iQ��  �  I#��������;��\t���r���y���H���#�C��	9��lμy0��k�����ü'�ռxL󼪎��-�dV������)��#^Ƚ���y
��J���"�%�k�t���̾⽤�Ž�ӳ�����g���Hս�^�� ��66��'$���%��A��T�'���۽xJ�������Nq���D�B]"��7	�s]�Zټ��ͼ�'ͼ]׼��e������?�^k�e��V���8׽����|����O%���$�������E����ڽ�����봽]~����Ƚ�潷��b���#���*�x�)��M!�_���� ���۽	����8��#}��U��Y7��["�:���*�)�'x����a%��/:���V���|�����.u��݆׽J���`�2�"���.��3���0��&��W��;����ؽYн�׽����~����(�`/4��{8���4� *��%��z����Kƽ����N�r}�w�b��`P��D��7?���>��D�oN�@�^��v�Gˊ�=m������xQٽ�����[��
%���4�uT>�$�@���;��/�]������� �𽊁����	��x�/,���:���C�=KE�p�>��2��� ��}�b���ӽAx������u�����yut�F(i��tc�gc�"h��r�����ƍ�I`��.,����ϽE���
�?�E�/��=�|�D��CD��+<��.���T:�����KE����&���-!��2��?�`�E��zD���;�o"-�.��_��M.��n˽Z\���ꜽ%���4e���u���l�G4i���j�r��~�r���˖�n/��=�����޽Y� �]��x�&��w7�14C���G���D��:��.+�b��:
����>������b��'[���)�"�9���D��  �  ���� ��S�=��!ҽc����/���|�3�S��U2�� ����+���ۼ�׼��߼���D�	�ɨ�X<�H�_�ܡ������
��0IܽU8���j	���P���n���h�� $˽���埢�Ɵ��������2ܽ�@����	���GE�]�x���83ͽ�Ү�j]����w��Q�<�1����AO���q7�)|�Q��v��[��,�.���L�i�r��R���X���}ɽ{��!���n����e��X������A�=�Ľ����6������õ��Ͻ������N��p
����o+�����P�ޙϽu^�����������b��dG���2���#��Y����G���%�105��jJ�r�e�����嘽Uұ���ν?���R�-��U�!��T�H��7j�V�\�ؽy@ƽ����mƽ�Fٽ0���A�	�K ��!�)�%��d#����������V߽�ý����7\��!��	s��K`�.�S��M�y�L��R�1�]�1�n�Q	��M֑��)���d����ԽZz�l	�"�U�$�)y,��9.�)��+��U�����x���޽x�ܽJ������[�َ��d)��X1���2�(.�+�#�%��4����ZOҽ)���J7�������7���	����w��(q�׽p��iv����Ɖ�s���ܤ��Է�/�ν1� �N����!�'�,���2���1��*�Xm����;%����2u�O�b�h�M�j�!��:-�/3��}2�ޟ+����|7���D��g�˽ɵ�.ң� ����{��~�����z���v���x��b��T��?@��YV���殽�UýU�۽�Y�����C��}(���1�S�5���2��)�KB��>�c?��62�J�8�9����'5��	)���2��  �  �w��������-�׽T�½ܬ��A������W�i�qYL���2��/�M�����AR �<��@��W#�[a:�Y�U�Qtt��������@���Uʽ�>߽�(�������S��F߽�ǽ�2��Y��������������ȥ�Y��g(ֽ�\���+���V���c�Uֽ�e��ɪ�w���������h�nL�"�3���� #��>	� ��������<&1��?I�xGe�k���U\��A;��g�����ӽ�S罼%��, ��`u��Dڽ����ᝪ��٘��#��	9���ܞ��ݳ�fVͽ7d潃V����̓������`��\۽��Ž����������6'|�
.b�jL��;���0�O1-�a1��^<�PN���d�9��`������������Ƚ�޽��������
���0B	��������ս:´�谽����8_��������׽}k�{��	����#���L
�Ӂ���]�ؽ� Ľ����q���"��І�]fy�.|j���a���`��@g���t��$��YT��!����}���O���Խ ��� ��
�XF��s�y
�1��9��� �L��>�ս(ʽsvȽԌѽ��㽉����z
��6��'��:� \��_�W�
�D�������ս�cýw#���Ť�&]���:��o↽�䂽�����'������ٖ��򢽥��������ҽ����v��+	��1��������K���j���K���ս,?̽��ͽVٽEn�����L�� ��4H����t�����4���@~�Yѽʿ��c��Uޢ��`��gN���5��|��� І����>Ɠ�����r��.J���˽"�ݽ�u�T9��	T������ �������m�
������q�'�ֽ0�н�ս���)���
��}�����  �  ��ν�xн�1̽��ýP���a:��+%��������?�t��Y���@��,�����*��v"���1�`�G���a���}�:q������/���}��/a��!ɽ!ѽgԽ7�ѽk4Ƚf丽�⥽Lq���7����p�=m��Tz����aɝ�����K(ý��Ͻ2�ս7�Խ-�ν�~Ž91���5���<��������t�@�Y���A�b�/�p%���$�K�-�iy?�T�V��Yq��O������Z��㦬����G#Ľ!�ͽ��Խ�ֽ�ѽo�Ž���-䡽��������v���y����iΗ��5�������~ѽ6�ܽ��a߽�&ؽ�Iν�
ý�S��(Y����
��@��Zcq�Ε\��gN��I�a�M���[�:q�;Ʌ�����g��g.��zN����ɽ�HֽS�ὸ�꽚D������A�۽~[ʽ�;��k/���������CR��Χ�K���ӌν�������m���V���P��]�$w���ؽ�ͽ���D���>��~T���|��%	��p�~�	�|�r,�������L��r��>n�����V5ν�4۽8���
����P������ �c��i߽��̽�d��C���1��(����ɽB&ܽ�`���e��l
��%
�.)�la�q\��B���Խ��ƽڸ�Ld��TZ��� ��
��������9��L���ǲ��������Ľ	ҽ�޽G�[c��gt�)f��	�7b
�������5�ŝ߽X�̽N_���������W��A7ѽز佝'�����P	�/���	�KF�+�����	�꽩t޽��ѽ|NĽ6����ө��Þ�������W��8M���Z���屽ڒ���[ͽ!�ڽ�u�������ɘ�U$
�M���l����I����e޽W�̽[|���黽Lڿ���˽~&ݽq�����	��  �  '𬽱���&q������3������"�������m��&��Zֆ���n���T�U�C���>��5G�7[�*Jw�߃��Κ�_���KT������غ�2������D���.�����IJ����������o��V�1�G�,�D�(O���d��̀�p���ӡ��������ω���o��fs������Uϻ��-��R������뻕����r�m��(V�½H���G�[T���j�]0��
쓽�d������M��c@��ݫ��IX��������	���������ۓ�A�����l���W�!N��XQ��Qa���{��������������ù��6½!^ǽ�ʽ��ʽmUʽ��ǽP�½�	��F,��-ޟ�Zѐ�xT��2�s��k�YZq������6��Oq��5ǯ��/��Sgɽ-ѽp�ս��׽.4ؽ�5׽�3Խ�aν�1Ž�ʸ��/��2��/���z�������w��f>��f|���஽������̽m�׽��޽���r���dr㽒	�ɱٽ~�Ͻ�ý�Q��6�������M��:���x��N$��Wﭽgw���\ν1�۽���Ws�$����J��	���� E�6ܽ�.Ͻkt��A���b�����������ä����y���UϽ�޽#��5��\���t���-����!�����V��x�-�⽍EԽ vĽAY��0b��\����:��=�������r½%9ҽi��"��8��������X��'���Y��o�������.J�/o���ѽ(½R����v���ڢ�٬���Ϊ�#��'Nƽeֽ�^�a���~��g"���_��2�������2��������`��ѽ����~ĳ����J��q���o��h���˽Q۽I/齥���;���p��ñ �+� �mI ��_���N��������u�ѽ�\½�����]���秽�󪽚�������Wѽk�བྷN��  �  �b������s��Mv��"sĽ�ͽ_Nѽ��Ͻ�Xǽ]츽3[����Bʁ��`m�kg�A�q��Å�3뗽)⫽u��7�˽�ҽ�%ӽν|ŽC��~-�������dg��\�u���Z��B�f]/���#�i�!�B�)��;:��Q���k�錃����3��u���a¶�u½��̽��ӽ�\ֽqiҽ��ǽ���W.��쐽1t��Saq�'hp�����掽`䡽�t���#ƽlѽ�ֽTaԽL�ͽs�ý���Z��؟��9��# ���q��+X��*B�Aq2�3e+��D.���:�ގO�ɸi�sB���ؑ�����`d���R����ƽv�ҽ�~ܽ"�����1�ݽ��ѽ����Ğ������xM���
���F������b��Nx���9ҽ⽱�뽮�����S�ٽ�Gνso½}T��ǩ�mǜ�]ď������Ss�Vqf�^�b�E�h��"x��T���̔�\#��@`��3���	̽��ؽ}�����ߺ��	:��������彥�ӽ����>{����y���n���}A���ʽ۸޽u�P���3��/�<��C�����ａp�ʺؽF�̽�@���k��sͦ�9k��p��������f��b����Κ������X��m½Y-нPGݽs������� �&���	�m�
�˔��8��!������GϽW�����.n��\K��� ͽ:$����>�����K
��y	����&�������Bt޽�ѽ�ZĽ���r����������T������k��ᠽ�������|cȽ
�ս"���ｲ*��IK�r���)>�W0����[Q�M�޽�d̽r��������"'ƽ��ֽj��o����� :����`�
����(��ת������E߽/fҽ��Ľ�~��ͪ��3�������!ؘ�G̟��_���4����Ľ�ҽ�  �  ���;������4�ý�ؽ%��u��(_��ګ�{�߽�ɽX���К��������qT������w����Ͻ�����������ܝ��a��(W׽}���AB���엽����pj��}M��b4����P�rx������!� ,���C�`_���~����M����)���&н��佟i�����c���'��-Sݽ�*ŽY߬�B�����"������0U��Q½?�ڽ��������
����z��~ҽ*���{B������� ���d���I��2�7� �g�����+L�+y��X-�̸C�{�^��}�Ǟ�������t��,�ͽ���bu��S��X�����L������̽0t��$��2)�����J$���ǽ���-���+��c`
�Z
�U5�����*{Ͻ�ͺ�0��c��@����x�{c�hS��bI���F��L�&aX�6�j�3B�����y����5�� �ýi�ؽ~��F��D���}I����r��~��Qc޽<zɽ����$�������ѽ���,�����o������d��_j�����Ix⽐�ν뾼�����h7���j��(ى������~���~��	���$�����lW��?���vp��O:н#��rc�����
��ڱ�|���5��������D9뽬�׽O\̽��˽
�ս��GG �<���\�����'�1��R���T������ ҽe��؞�������і�>B�������S��؃����K����7��	���n^Ž{�׽��C� �Y������d���*������I��������ս�,ν�VѽԿ޽'��9d�4�s'�ձ��>�$3�]��@X�$����� ѽ���l����ţ�0����������3���}k���ߏ�v������$ఽ����  �  Y}��𗽄%Խ$��*�E���C�OE��e�� �T$ͽ�벽_��������Ԥ�������Խ����������H�-q�����Fн����^����A{�H_S��-3�w��P��i��9[�8�2���[�@���(�
lF�6k�>	�����FpĽʥ㽵u �	�a�������_�y�彁�ǽc��,���Gġ� ��g�Ľ��̠��&�������~�\������ǽ����D��*_q���L��S/���L
	�fT��:���e���z�����)�1<D���e��<������� ��}۽Gv���J���-|����s ��t����8н�@��$ŷ���Ƚ�3�� �ݐ�yi��~�p��X�
�τ����׽u캽����Ό�	�w��\]��I�"�;��14���2��7�k}A���Q���g��0���ޓ�Fc����½�/�q���|��
��$�Y_'���#�X��DM��,��Y����н �̽0sսU꽀G����k^ ��z)��j,���(��s�*�P����O̽����h��������]�z�/Jo���i��j�_Np�b|�k��6쒽K���e����)˽������e�����+�a!2�g2��2,�Ǡ �q��p*��e�X�པ�߽�4����%&������*�$�1��>2�3N,�1!�+��N������ͽW��8X���d��[ɉ�B��5\w�H$r��s���y�	a��A��C��0��Q뼽��Խ���}��Z%��%�=/���3��2���)�2��=��, �	��C�潓j���('��h%���/�P�4�-#3��Y+�����ė ��&���ʽ�s���$��k��Q�u������|�R��~d��֋�G����*���  �  nz�����Z����彧��ޚ��L ���#��n���~���n&ǽ=!��K���Ŷ��ͽ3���}�����!�ȷ$���˺���7G��� ��v� �G���#�Q�	�\7�Sּ��ɼ��Ǽ�м/�W����Z�8���b�����k7��8�н�������]���$�w�%�x���g�� ���޽�<ýX���������6P۽���}���n�]%%�&4%������������Yս>e���̏�Q�i�]s?�������c��⼏�ۼ��%/����j���4�X�Y�mA��h����ý!��j�6����&���,�N+�^Q"�)����Z��U'νI�ý�ɽa�ܽ���ZB�� �&q,��2��/�u&���wb�y���+��m���ڇ��ui�57M�+y9�&�,�41&��%��")��2���A���W���u�ࠎ�Ƨ���ƽZ�5}��d��|+��G6���9�w�5���*�g��;�	����b`�g0ݽcT罧��}��^�!��l1�{�;��>���9�*=.������
�Dg��ν��������V����{���j��w`��[�&C\�t�a���l���}�l犽	���P���˽�a���zV��m-���;��,D���D�4�=���0�Ҵ������ ������� �����_��׽.�4�<��SD��jD���<��.�/2���	���Bν�(�������~������s�|i��d��Ee��]k�iw�Z���7���#��K㹽tsֽzp��/�O"�Έ3�q>@��DF�ED��H;�,�,�G2���
�h�������b��!�=�Am%�u�5��B��aG�?�D�;���+�2���pi�;�ɽl��������X��僽'�y���q��/o�W�q��y��׃�_,��Y���[ٯ��  �  N{����Ƈǽ��
��{ ���,���0���+��m����o���X�Խ'þ�G^��q�½$�۽I��ѫ�qy#�kx.��e1���+�S7��m�4콎����G���v���B�ԡ�|.��7ݼc	Ƽ� ���Y��Y����YӼ��
��2��\`�ħ������ڽ+�<����'��<1�lI2���*��D�k�	�/3���Ͻeɾ�0׽��Uͽ�S�O���O��m)�I�1�}�1�7))���֏�]�߽Rd��8䑽��g���9����dt �i��\0Ҽ��̼R=Ѽ�3༐W����g}-�ڃT���L����ʽ�������R$���2�t�9�L�7�.��(��~����Jڽ�Ͻ6�Խo��Ԃ�����2+��8�W�>�J<��1����T>�^��Y�ýi����*����b��E�.�0�ޏ$�[M��J��I!��g*�ST9��O�|�n�x���@h��]�ʽ����bP$��]6��|B���F��B��5�l�$����������;�<�8��#r���+�-=��IH�`wK�5�E���8�&����V�����ѽt���%��}����Is��Ab�	=X�C�S��kT�u�Y��~d��8u�����i�������̽+��E���"�C7�n9G�;�P���Q��J��;���(��D�.#�������/���C�˷&�Zp9�Y�H���P���P�LfH�N�8�2�$��>������Sн�>���ݚ�s���(�z�K�j�#a�,�\�Yy]��Cc�֚n�\`��kȍ�B���{���<Pٽ�b������y*���=��L�Z�R�WQ��G� �6�*�#����������q������/��A��TN��T��4Q�$F���4�- ��
���콚�ʽ�Ү�⤙��=��=�=�q���i��qg�k�i�n�q��$�p��-%���ﭽ�  �  �U|�8m����ʽ����o���f$�Z�0�f
5��70�Dr#�Ue�C���Ckٽ7�½�@����ƽ���ً��F�j�'�B�2���5���/�� "�ǂ���𽋢Ľe���F�v���A����E��)�׼J�����cK���k��μ�{����1��`�ӌ��������޽h����`�+���5��6��/�& ������zԽ5�½������ѽD����
�1�ѯ-�lT6��96�2P-��&�
b�S��͸��풽�g��E8�"�������ݼ�ͼ~�ǼF>̼ۼ/ ���~��X+��KS�v!��来�Ԝͽt��ƙ�y�'�-�6�a>�vd<��B2��!�ޔ� ����޽�ҽ��ؽ�|�LU��J��(/�<=�	DC��m@��5��D#�������Ž14���څ���`���B��J.���!�������~����'��6�%M�y�l��W��_��}̽���r���'��I:���F��(K�X�F���9�1"(������7��j������s�?�/��A��L��O�C5J��|<��-)��8�/����Eӽ�W��X���^�����p�;�_�&�U�qCQ���Q��IW���a�
�r�����^;��:�����ͽ[����br%��:��QK��U�A'V��^N�y]?�'A,�����`	��} �9���������>�)��:=��L��U�jnU���L�Kj<���'�/=��U��p[ѽ�5��(��5k���.x��h�"p^�q4Z�#�Z�9�`�P�k��.~�����ꟽ������ڽ0�~��x-�O�A��UP��kW���U��3K��:� '������2� �v�R����y2��	E��R�{�X��U�pJ�-.8��"��C�����1˽����������|��n�f\g���d��hg�o�ǀ|��Ȉ�:.��~����  �  N{����Ƈǽ��
��{ ���,���0���+��m����o���X�Խ'þ�G^��q�½$�۽I��ѫ�qy#�kx.��e1���+�S7��m�4콎����G���v���B�ԡ�|.��7ݼc	Ƽ� ���Y��Y����YӼ��
��2��\`�ħ������ڽ+�<����'��<1�lI2���*��D�k�	�/3���Ͻeɾ�0׽��Uͽ�S�O���O��m)�I�1�}�1�7))���֏�]�߽Rd��8䑽��g���9����ct �d��V0Ҽ��̼H=Ѽ}3༂W����]}-�σT���
L����ʽ�������N$���2�q�9�I�7�.��(��~����Jڽ�Ͻ7�Խq��Ղ�����2+�
�8�[�>�N<��1����X>�e��`�ýp����*����b��E�4�0��$�]M��J��I!��g*�NT9���O�s�n�r���:h��V�ʽ����^P$��]6��|B���F��B��5�j�$����������;�<�9��%r��+�0=��IH�cwK�8�E���8�&����]����ѽ{���%�������Is��Ab�=X�H�S��kT�x�Y��~d��8u�����i�������̽+��E���"�C7�n9G�;�P���Q��J��;���(��D�.#�������/���C�˷&�Zp9�Y�H���P���P�LfH�N�8�2�$��>������Sн�>���ݚ�s���(�z�K�j�#a�,�\�Yy]��Cc�֚n�\`��kȍ�B���{���<Pٽ�b������y*���=��L�Z�R�WQ��G� �6�*�#����������q������/��A��TN��T��4Q�$F���4�- ��
���콚�ʽ�Ү�⤙��=��=�=�q���i��qg�k�i�n�q��$�p��-%���ﭽ�  �  nz�����Z����彧��ޚ��L ���#��n���~���n&ǽ=!��K���Ŷ��ͽ3���}�����!�ȷ$���˺���7G��� ��v� �G���#�Q�	�\7�Sּ��ɼ��Ǽ�м/�W����Z�8���b�����k7��8�н�������]���$�w�%�x���g�� ���޽�<ýX���������6P۽���}���n�]%%�&4%������������Yս>e���̏�Q�i�\s?�������[��⼁�ۼϜ�/����j���4�C�Y�aA��h��{�ý��j�/��y�&���,�N+�XQ"�%��
��U��S'νH�ý�ɽe�ܽ���^B�� �+q,��2���/�|&�&��b����	,��y���*ڇ��ui�E7M�7y9�.�,�91&��%��")��2���A���W���u�ՠ���ŧ���ƽ�Y�.}��d��|+��G6���9�q�5���*�c��8�	����``�g0ݽeT罫�����b�!��l1���;��>���9�1=.������
�Sg��ν��������V����{���j��w`���[�.C\�z�a���l��}�m犽
���P���˽�a���zV��m-���;��,D���D�4�=���0�Ҵ������ ������� �����_��׽.�4�<��SD��jD���<��.�/2���	���Bν�(�������~������s�|i��d��Ee��]k�iw�Z���7���#��K㹽tsֽzp��/�O"�Έ3�q>@��DF�ED��H;�,�,�G2���
�h�������b��!�=�Am%�u�5��B��aG�?�D�;���+�2���pi�;�ɽl��������X��僽'�y���q��/o�W�q��y��׃�_,��Y���[ٯ��  �  Y}��𗽄%Խ$��*�E���C�OE��e�� �T$ͽ�벽_��������Ԥ�������Խ����������H�-q�����Fн����^����A{�H_S��-3�w��P��i��9[�8�2���[�@���(�
lF�6k�>	�����FpĽʥ㽵u �	�a�������_�y�彁�ǽc��,���Gġ� ��g�Ľ��̠��'�������~�]������ǽ����D��*_q���L��S/�}�F
	�VT��%���K���z�����)�<D�|�e��<������� ��h۽2v��{J����$|����l ��t����1н���@��&ŷ���Ƚ�3�� ����i��~�y��X�
������׽�캽����"Ό�$�w��\]�'�I�.�;��14���2��7�b}A���Q���g��0���ޓ�5c����½�/�\���r��
��$�P_'���#�Q��>M��,��S����н �̽3sս[꽄G����r^ ��z)��j,���(��s�*�[����O̽(����h��-������q�z�@Jo���i��j�hNp�!b|�n��7쒽K���f����)˽������e�����+�a!2�g2��2,�Ǡ �q��p*��e�X�པ�߽�4����%&������*�$�1��>2�3N,�1!�+��N������ͽW��8X���d��[ɉ�B��5\w�H$r��s���y�	a��A��C��0��Q뼽��Խ���}��Z%��%�=/���3��2���)�2��=��, �	��C�潓j���('��h%���/�P�4�-#3��Y+�����ė ��&���ʽ�s���$��k��Q�u������|�R��~d��֋�G����*���  �  ���;������4�ý�ؽ%��u��(_��ګ�{�߽�ɽX���К��������qT������w����Ͻ�����������ܝ��a��(W׽}���AB���엽����pj��}M��b4����P�rx������!� ,���C�`_���~����M����)���&н��佟i�����c���'��-Sݽ�*ŽY߬�B�����"������0U��Q½?�ڽ������������z��~ҽ*���|B������� ���d���I���2�/� �]��z��L�y��X-���C�Z�^��}����������t���ͽ���Ju��G��M����:������̽(t�� ��1)�����P$���ǽƇ�=���4��n`
�f
�a5�4���'�C{Ͻ�ͺ�F��(c��Q����x��c�wS��bI���F��L�aX�#�j�'B�����f����5���ýP�ؽd��F��D���rI�����r��~��Fc޽5zɽ����#�������ѽŲ�,�����o�ɐ���q��lj����bx⽨�ν�������y7���j��5ى������~���~��	���$�����mW��@���vp��O:н#��rc�����	��ڱ�|���5��������D9뽬�׽O\̽��˽
�ս��GG �<���\�����'�1��R���T������ ҽe��؞�������і�>B�������S��؃����K����7��	���n^Ž{�׽��C� �Y������d���*������I��������ս�,ν�VѽԿ޽'��9d�4�s'�ձ��>�$3�]��@X�$����� ѽ���l����ţ�0����������3���}k���ߏ�v������$ఽ����  �  �b������s��Mv��"sĽ�ͽ_Nѽ��Ͻ�Xǽ]츽3[����Bʁ��`m�kg�A�q��Å�3뗽)⫽u��7�˽�ҽ�%ӽν|ŽC��~-�������dg��\�u���Z��B�f]/���#�i�!�B�)��;:��Q���k�錃����3��u���a¶�u½��̽��ӽ�\ֽqiҽ��ǽ���W.��쐽1t��Saq�'hp�����掽`䡽�t���#ƽlѽ�ֽTaԽM�ͽs�ý���Z��؟��9��" ���q��+X��*B�6q2�$e+��D.�u�:�ÎO���i�_B���ؑ�����Fd���R����ƽY�ҽ�~ܽ�⽨���ݽs�ѽ������������tM���
���F������m��\x���9ҽ����������o�ٽ�Gν�o½�T��ǩ��ǜ�mď������Ss�`qf�`�b�?�h��"x��T���̔�J#��+`�����	̽��ؽ`�����ú���9����������彖�ӽ����6{�� ��y���r����A���ʽ�޽��f���?��<�J��`�����｝p��ؽ_�̽�@���k���ͦ�Hk��|��������f��h����Κ������X��m½Y-нPGݽs������� �&���	�m�
�˔��8��!������GϽW�����.n��\K��� ͽ:$����>�����K
��y	����&�������Bt޽�ѽ�ZĽ���r����������T������k��ᠽ�������|cȽ
�ս"���ｲ*��IK�r���)>�W0����[Q�M�޽�d̽r��������"'ƽ��ֽj��o����� :����`�
����(��ת������E߽/fҽ��Ľ�~��ͪ��3�������!ؘ�G̟��_���4����Ľ�ҽ�  �  '𬽱���&q������3������"�������m��&��Zֆ���n���T�U�C���>��5G�7[�*Jw�߃��Κ�_���KT������غ�2������D���.�����IJ����������o��V�1�G�,�D�(O���d��̀�p���ӡ��������ω���o��fs������Uϻ��-��R������뻕����r�m��(V�½H���G�[T���j�]0��
쓽�d������M��c@��ޫ��JX��������	���������ۓ�>�����l���W�� N��XQ��Qa�~�{��������������ù��6½^ǽ�ʽ��ʽPUʽ��ǽ7�½�	��3,��ޟ�Nѐ�oT��(�s��k�_Zq������6��]q��Gǯ��/��lgɽGѽ��ս�׽L4ؽ�5׽�3Խbν�1Ž�ʸ��/��,2��/���z�������w��_>��[|���஽������̽U�׽�޽ߙ��q����Gr�w	཰�ٽh�Ͻ�ý�Q��*�������M��:���x��V$��cﭽvw���\νG�۽���rs�6$���h��&����E�#6ܽ�.Ͻ}t��P���b����������ä����|���UϽ�޽#��5��\���t���-����!�����V��x�-�⽍EԽ vĽAY��0b��\����:��=�������r½%9ҽi��"��8��������X��'���Y��o�������.J�/o���ѽ(½R����v���ڢ�٬���Ϊ�#��'Nƽeֽ�^�a���~��g"���_��2�������2��������`��ѽ����~ĳ����J��q���o��h���˽Q۽I/齥���;���p��ñ �+� �mI ��_���N��������u�ѽ�\½�����]���秽�󪽚�������Wѽk�བྷN��  �  ��ν�xн�1̽��ýP���a:��+%��������?�t��Y���@��,�����*��v"���1�`�G���a���}�:q������/���}��/a��!ɽ!ѽgԽ7�ѽk4Ƚf丽�⥽Lq���7����p�=m��Tz����aɝ�����K(ý��Ͻ2�ս7�Խ-�ν�~Ž91���5���<��������t�@�Y���A�b�/�p%���$�K�-�iy?�T�V��Yq��O������Z��㦬����G#Ľ"�ͽ��Խ�ֽ�ѽn�Ž���*䡽���������v���y����[Η��5�����o~ѽ�ܽ��F߽�&ؽ�Iν�
ý�S��Y����
��0��Bcq���\��gN��I�f�M��[�Nq�IɅ�����g��.���N���ɽ�Hֽp����꽵D�	����U�۽�[ʽ�;��t/��
�������@R��Χ�@���Ōν�������m���V���P��@�w���ؽmͽ�����C���>��oT��|��	��h�~�	�|�v,�������L�����Pn������n5ν�4۽T����4��^��)���� �x��i߽�̽�d��C���1��.����ɽE&ܽ�`���e��l
��%
�.)�la�q\��B���Խ��ƽڸ�Ld��TZ��� ��
��������9��L���Ʋ��������Ľ	ҽ�޽G�[c��gt�)f��	�7b
�������5�ŝ߽X�̽N_���������W��A7ѽز佝'�����P	�/���	�KF�+�����	�꽩t޽��ѽ|NĽ6����ө��Þ�������W��8M���Z���屽ڒ���[ͽ!�ڽ�u�������ɘ�U$
�M���l����I����e޽W�̽[|���黽Lڿ���˽~&ݽq�����	��  �  �w��������-�׽T�½ܬ��A������W�i�qYL���2��/�M�����AR �<��@��W#�[a:�Y�U�Qtt��������@���Uʽ�>߽�(�������S��F߽�ǽ�2��Y��������������ȥ�Y��g(ֽ�\���+���V���c�Uֽ�e��ɪ�w���������h�nL�"�3���� #��>	� ��������<&1��?I�xGe�k���U\��A;��g�����ӽ�S罼%��, ��_u��Cڽ����ޝ���٘��#�� 9���ܞ��ݳ�WVͽ&d�oV�������j���~`��\۽��Ž����������'|��-b��iL�ӝ;���0�M1-�f1��^<�bN���d�X��#`������آ��ʛȽ!�޽��������
���:B	��������սB´�谽����5_��������׽pk�{��	�������L
�Ɓ���D�ؽ� Ľ����q���"��І�Ify�!|j���a���`��@g���t��$��fT��1����}���O���Խ��� ��
�eF��s��
�;��B��� �Y��I�ս1ʽzvȽٌѽ��㽌����z
��6��'��:� \��_�W�
�D�������ս�cýw#���Ť�&]���:��o↽�䂽�����'������ٖ��򢽥��������ҽ����v��+	��1��������K���j���K���ս,?̽��ͽVٽEn�����L�� ��4H����t�����4���@~�Yѽʿ��c��Uޢ��`��gN���5��|��� І����>Ɠ�����r��.J���˽"�ݽ�u�T9��	T������ �������m�
������q�'�ֽ0�н�ս���)���
��}�����  �  ���� ��S�=��!ҽc����/���|�3�S��U2�� ����+���ۼ�׼��߼���D�	�ɨ�X<�H�_�ܡ������
��0IܽU8���j	���P���n���h�� $˽���埢�Ɵ��������2ܽ�@����	���GE�]�x���83ͽ�Ү�j]����w��Q�<�1����AO���q7�)|�Q��v��\��,�.���L�i�r��R���X���}ɽ{��!���n����e��X������A�:�Ľ����6������õ��Ͻ������E��g
����e+�����P�əϽb^��
���������b�wdG��2���#��Y���H���%�?05��jJ���e�����嘽hұ���νS���R�7��(U�!��T�O��=j�V�c�ؽ|@ƽ����mƽ�Fٽ(���;�	�D ��!� �%��d#����������V߽�ý햪�(\��	!���s��K`�#�S��M�x�L��R�<�]�A�n�\	��Z֑��)���d����Խnz�v	�*"�_�$�3y,��9.�
)��+��U����y���޽}�ܽO������[�ڎ��d)��X1���2�(.�+�#�%��4����ZOҽ)���J7�������7���	����w��(q�׽p��iv����Ɖ�s���ܤ��Է�/�ν1� �N����!�'�,���2���1��*�Xm����;%����2u�O�b�h�M�j�!��:-�/3��}2�ޟ+����|7���D��g�˽ɵ�.ң� ����{��~�����z���v���x��b��T��?@��YV���殽�UýU�۽�Y�����C��}(���1�S�5���2��)�KB��>�c?��62�J�8�9����'5��	)���2��  �  I#��������;��\t���r���y���H���#�C��	9��lμy0��k�����ü'�ռxL󼪎��-�dV������)��#^Ƚ���y
��J���"�%�k�t���̾⽤�Ž�ӳ�����g���Hս�^�� ��66��'$���%��A��T�'���۽xJ�������Nq���D�B]"��7	�s]�Zټ��ͼ�'ͼ]׼��e������?�^k�e��V���8׽����|����O%���$�������D����ڽ�����봽X~����Ƚ�潳��]�z�#���*�q�)��M!�W���� ���۽�����8��}��U��Y7��["�1���*�)�)x����a%� 0:���V���|�����;u���׽Y���g�:�"���.��3���0��&��W��;����ؽYн �׽����{���(�[/4��{8���4��*�~%��z�x��Kƽ겨�C�r}�h�b��`P��D��7?���>��D�wN�K�^��v�Pˊ�Gm�������Qٽ�����[��
%���4�|T>�+�@���;��/�a������� �!𽏁����	��x�/,���:���C�=KE�p�>��2��� ��}�b���ӽAx������u�����yut�F(i��tc�gc�"h��r�����ƍ�I`��.,����ϽE���
�?�E�/��=�|�D��CD��+<��.���T:�����KE����&���-!��2��?�`�E��zD���;�o"-�.��_��M.��n˽Z\���ꜽ%���4e���u���l�G4i���j�r��~�r���˖�n/��=�����޽Y� �]��x�&��w7�14C���G���D��:��.+�b��:
����>������b��'[���)�"�9���D��  �  ��/���+�e��Q�Zu�u�Ž�]���z���D�"��/����(׼	��$x���,��ڳ�(�ļ�0⼝e��^'���R�兽����|�ѽ�����H�Rp$��9/���1�(�+��2�)�����ҽ�D�����E�Ƚ��㽀��-��E'��0��62��+����\	�������Yf��Up�RU?���e� ��s޼ �ȼ�6������|�ƼP(ۼ�\��j��U:���i��Y��JE���⽚��7p�H�)���1�1���(�փ����ï�5�ͽ�����½�ս�����7 !�ö/��A7�"&6�(�,�d��&��r��漽ε��miz���N��F/����/T�[3��i�F��L��1����1��O��4x����s����;߽}(�{���k-�w�:��A@�&=�72��o!�֯��r����㽲f۽ܪ�5J������j"�k+4���@�/E��A���4���"�S��pD�]5ʽ�%��鎽�nv�
uZ�R�G��<��c7��H7�y-<�i@F��RV��m�����㝽�����$޽<���[�CR.���?�ɯJ���M���G�u�:�P)�Ӧ�>2�=�������%�� �oM#��v6���F��nP�#�Q���J��5<�Ӻ(�E)����\ֽ����8[��5򋽗�}��l��a���[�.P[���_��j���z�@㉽�����e���ѽp���vf�]&���9��*I�$RQ�=�P�0H���8��%�=����
r��:j��G����*���<��<K��^R�t�P�nG���6��9"�H��*s�/�̽Y���̙��{���<|��gm�+�d�xta��c���i� Mv�&ꄽ\-��0�k������<��6Z/��B�U=O�}�T��hQ�")F��E5��B"����\] ��+����� ���3��>E��iQ��  �  ��ʽ�dŽ�Z�����`���V��k%����򞳼�n���<�����/7û���-�̻T���q�S��"���ȼ��=�4�2�g�厽)����彽�9˽�wνi*ǽ\ⶽ����5艽k�l���T��P���`�I��K��!���<	½@�ͽ��ϽI�ƽ�紽�뜽=7���O�4s ����20���ˆ��N�� %�_�&� �� ���
���!�%I��Â�����]�W���XJ���~�7��ǲ�ڟŽ��Ͻ*�ϽEŽ���y-���8����j�~6Z��"^��v��莽�ᦽ@���eнX�ٽ:�ؽ�!ͽj_��4���V��w�Y���-�Z�	���ݼq뷼Q�����V����=���A��c���z��=�ļ�꼥��9�0�g[�֘��x������)�ӽ�X�Bc�2��M�ڽr�ƽ�����j��X6��C��x����m������@ʽj�߽t/�N�����ｃ:� @˽/d��Y����#}�ʱS�6�2�w���
����T�4�&�Q���?����� ���/��-L�uq�"������lĽ��޽�'���� ������<}�JRڽ�	Ľ�T��S�������'���k���ս���4 ��4�}����/�󽳜۽���Pk�������u�n�V���?�L�/�.9%�������0���Q��!$�$.�3/=�{%S��2q�/��P��̊��vؽP
���_������x��J�kkٽ�ý&�������A���20���5ȽyQ߽������l��O ��� �\�� �Խ�������ݽ��o��$S�?�ԃ1���(�$�j"�Yq#�EV'���.�Iq:�|�K���d�b���֗��p���J˽������g��~
�6 �Y�9� 
׽'������K����L���y��Zcս%����|��  �  :]Ž�F���ɱ�|Y���1��z�R�zo#����J���#烼�_B�������L�λaȻmػ�} �R�#��0Y��]����ȼ�D��)2�$xc��؋�����=/��TƽhɽP½�2��n윽ȉ��W?g���O���K��O[���{�܎���������ȽDʽ��������7t��Mi���L������`ӵ�����F�T�ކ+�c_�L^�P�����(�m�O�;���MN���\꼀u�zkG�D�y��ږ�d�������|ʽ�1ʽ,��3:��6a�����Yte�'bU��>Y�[�p�����[ܤ��EJ˽�tԽgӽ[Ƚ�Q���c��݃��W�s�,�A
�i�߼:꺼�^���������{��������������Ǽ�켪���0�?�Y��҄�����6Ӹ�*XϽ�E߽D�(���ս0h½�g���o��ॊ��څ��������t����Ž�۽���ܓ�j�꽷�ܽ�{ǽ��������({��)S�)w3����"��4+��b�������S���Ho�3��?�_�0���L��@p�b�}�u_���ڽp�+����0 ��������5Eֽ����Z��������������N��SUѽ�;轆m�����w�rA �iN�D$ؽ�R��	ڤ�mꍽ�uu�`VW��A�$O1�W�&��l ��W��%������%�p�/�?�>��T�1q�,M���١��#���ս{�콅����S�~�������ћսeۿ������P�������k��C�Ľ�Z۽�5��b<��b�g-����齂_ѽ����ٞ��@���=o�1T���@�^#3��x*���%�a�#��$�>�(��J0��<�\CM��ge��Â������Ƚ":�Ǌ��T�f`��z���0��tӽ)ﾽ؎���&��>ï�P���0�ѽV�轋^��A���  �  X���������Ow��9I�0������a���Ry��շV��"(���	��*�.��E���,��58�A"m��P��?�̼���jj,�#�X�k����ʙ�j	���u������v��v���Qz����y��4W�Y�A�)�=��GL��Cj���������������~]��:泽�����4�q�˪D�������2��~���g�i�'�?�fQ%��[�u��Q#�?<��Md�$��x!��}:켪��q@��m�����*΢��������=��'豽v���𛍽�9t�KKV�ܝG��NK���`��M��ȿ������伽�tŽ2�ĽQ�����/ϔ�,|�0�P��*�D��á�	�ļ�Ĭ�Q���V���a����)������ⷼS�Ѽbs��3��U0�aaU�<��:���j���v�½ѽ�׽�ӽVȽJT���9������W���}�wჽ_6��*������{�ͽ�A۽ ���ܽ��Ͻ���Z馽m8���zv���R��5�8A �J���K�l �Ա��P������N�z���.!��4�;VN��n�*��7q�� ��k�ϽG�b(�*R�T�/�ݽS�ʽ����p���q���'����et��v�ƽ1�۽�\�m'��P��t��uJ㽺�ν�����ڠ��O��<v�#�Z�ѫE�y6���+�(%�^�!�|�!�ā$���*�8�4��\C�sW�	r������$�������˽��V=����+C��Һ��!߽��ʽ۶��Y��#a��J������ň��н#'�՜�3q�����.���u޽��Ƚ��������#X���p�H�W��E��Q8�n/�C9*� J(�(h)���-��h5�'%A�b�Q��h������ה�-��.8��� ؽ�콂������"/��e�E�ݽFɽt��>���E������J;����ǽ|�ܽ��ｓ���  �  [i��4���8�����b�1�=�a�� ��!�Ƽ�l����}�5HN��6-���� O�� ��78�U�^�������Jؼ���B�&���J���p��v���6��S�������b���u��pQ]��"?��x,��)�n�5���O�jTr�l$��7M�����������៽����悽��`�5�;���|����T˼q���Sd��@e���G�f�8��28���E��Ea�K���&.����Ƽ������K�7���\�����:��QM������U��f��mێ�F#{��iY���?���2�Z6�IsI�p�h�����`��1���	����|���觽�^���7����m��xJ�&9+���	u��7ؼ<<���ѯ��Ӧ��$��͑��O��.�ʼ���+�����3��*R�ߪu��鍽F����������(���	��hƳ�/g�����P@��g�p��Ri�zr��Ą�0���ao��O���s�Ž�ʽ��ǽ�ڽ�ᰮ��Ŝ��d����r��T�)z<��:)�Ї�������ڏ�q����	��=�1@�=�*�T7=�MT�~�o�IA�����r�.L���nϽI�ؽ�K۽H�ս��ɽ��������LW��պ��+�������1���޶�F2ɽ��ؽ
<�	L�6�޽�Fҽr����㮽�\���u��A�y��b��O�8B@� 35�e�-�W�)���)��-�C�3�v�>���L�N_�r�v��s���������Q���sнݽ�:�5Q㽬�ڽ�Z̽벺�ha���㛽>������؂���h����н�_޽�r�����ܽ�ν+���w��r���ш���&v��[`�&0O��B�\�8�e�2�i^0�`�1��p6�$�>���J�|�Z�Oo�W���A��x���-���&ʽ�Hڽ�����~q�1�۽��˽J��w���?��T홽����$������3˽�۽�_��  �  mW��%�^~��-i���O��m5��4��H��ἊA���I��p{���5d��#M�hG��bS��vp�[T��#���t�˼��D�~R&��@�_v[�Q�t������~���ފ�;D����t�6�X�kL;�g["�����(�	��V0���L��j��-���y���������KP��`�k�SSQ���6�=�o��q�輎ƼgE����h}� �j�\�i��Jz�f����f���¼������/��W4��N��-i�,����o��্����>ʄ���q�1U��{9�|J$����;� ^-�T�G���f��ӂ����O��Pv���ڒ�������{�%b���H���1�\v�Ͳ�����%�߼T̼���������üR:ҼԵ�b�������&���<��tT�q�n�����Y���ĝ�����,���㤽����L��m��;*h�HdV��P�X���k��������������2��������"��Rȟ��R���Z��;�s�Ѭ]��J��$9�T�*�P��Z��A!������2�>�+���:�ٳL���`��
w�@����a���0��o.��ϼ���!��K	½�
��
첽r���&����ދ�1���	)��4��`������i��u��K�ȽƗ˽FȽ����Yf��C?������샍�'I����p�U?_��/P�]�C�;��b6�6��;:�̉B�dgN�/]�;n��ွ��7E��6����Ʋ�f���9�ǽX�˽�ʽ��½�N������~S��,��5n��yF��,����Ӝ�V����2����Ž�0̽��̽��ǽ[��ٱ���������>Ջ��8����o��u_���Q��F�|�?�
�<�%+>��	D���M��[���j�Q}��Ј�pm���9��o���,ͻ��ǽՑν��н�Oͽ3Ľ�޶��������!���������Zڙ��T���o���GĽ�Tν�  �  ��]�6 `��C[�+VQ��lD��6��<'�����/���u#ϼO�������/T���K��8��ɟ�_麼�ۼ�����I�����B/�@�>��GM��@Z���c���g�^wd�kY���F��/�#�}d�4v��,�3������=t&���>�H�S�� c�X{j�d�i��c�i�W�,J�4W;��',�b��@Y�`t���ּ����˓��V[����������-����Ӽ��m�
�����*���9�x�H�S�V�u�b� �j�oll���f��X��#E�R>.��h����|) �p��!�EI%��>���W�[%m��G{����x�&�w��\l��_�E�P�)sB���3�0R$�?��L`������伿`߼y�<"����	��z�|z,�yt>� �O��j`�0�p�l ��J���Ì�������������6���s�L�\�V�H�s�:�Ǣ6� �<���L�۫c�`)}�҇���֓�dX��zĚ������䓽
���Y������cp�UTa��Q�ޚB�_�4�I�)��o#�-�"�{(� �2��A��S��1e�qw����Z���b�����I䢽�����Y���?������쐽�녽t�y���n�Vn��w�����$ϐ�-@���1��t ���ϳ�졳�.��(�������L&���u�������[����w��xg���X���M��fG��G���L�n%W�7ve���u�<��n���X��Q��ɍ��E���J���cq���<���*���"�� 럽�����������v�_x��ρ�А���o���D������r��wε�wk��e&�����������;���@���&��|�w�+h���Z��vQ�!|M�OiO��W��[c���r��́�LE���}���p��#2��~����������'��6���{g���A��2]�����o̊��O����������[������=��ǣ���u���  �  ��4�qM=�\DB�i�D�B�D�6�B��r>��Y6�*����q�����ɼ�4��+����๼��Ҽ=*��.��� �t�0�ǜ<��kD���H���J�?�J�^H�AC�r:�Iz-������	�&���м�,�������ǼCN����o���(�m�7�PC�ZJ���M��\O�T�N�h�K��$F�Ҁ<�]�.�}X�H2
�v����Ҽ <¼�\���7м-)�'�xa�g-��];�8�E��K�UO��P�EO���K���E�ݾ;�L�-���ed
��1�Ղڼ�~ϼ �Լ�p鼒l�%��~�.�N�A��Q���[��b�X�f�yh�( h�#e�T�^���T�
�F���5�p�#�:����J��<��@� �%���9��fN��|`�ڧn���x�`�~�5倽Ce��n߀�?-~��Ew�ihl�:�]�%TL���:��++�!�68�>m#��0���A���V�\�j��7|��ф�f��}(������[፽�,���&��Ve������t�	xb��P�FB�K9���7��]>��L���^��ps�����C(��
����ݖ�}r��8���
���I��a,���H���c��۴����{�e�j�%L]���U��NU���\�&Ak���}����̐���\���	����������AH���@p��zo���������������s�� e�;�\��W\�P�c��q�x遽�����o��@���� �<���8����!��z���H���Ԡ�����z��r������Wr�a�d�2^�_���g��w�݄�����cN��{A��� �����)������0}�������B��PӜ�)[��)Z��Xۂ���t�;h�Y�b�6(e��Bo�5�'��/Β��S��?�������VE��0����檽(+��E'���m�������疽j���QR��x�d�l���h��tl�U�w��3������ m�������  �  ���Ԗ&�6���D�	MR���\�ȸa�3�_�C�U��MD���-�nD�q��-輯��N�����8��5���K��*\���d���e�&�_�~XU��H���9���*�:��J������<ռ����a}��}ے�娐�B<���b���nʼ����Y����'���6�	�E��T�`��"i���k�7g��2Z�*�F��/�|��f�������0�Rc��},��7D�l|X��<f�Fl�g%j�a/b�HV��XH���9���*� E�z���:����ؼ�ᾼӬ�2u�����(�����Լ���B���x1���B�fS���b�m�q��}��͂��j��(!����q�p�]��IG��`2��W#�nc��!�t�0�plF���_��Dx�����g2��K�������P���B����v��qh�P�Y��J�HZ;�Z�+�������
�@+	�3u��P���%�ؙ6�X�H��|Z��k��*|���ƽ��������=Μ�A���q���*��8w��Ucr���^�ȱR�j0P�DX��i�x���\������ǡ�e����~���m���,����ْ�͋�����xz��Yk�^\��,O��E�1�?��?�7�E�k"Q�d`�q��L���Ӊ������ڙ��u��d����î�e��QI��Ǳ��B��]��k����̉��J����u��u���~�������'���\!��v��1�������(��*:���?���Ԛ�+7���a��>D���u���e��W���M��H�k�I�>P��[���j��e{��'���d���Z��c�����Ǡ��a���嵽�&���v���᪽IR��^u���e��l<��R-{�<h~��Ʌ����� ��pȧ�� ��Pල������������˫����9O��Ƕ��ލ�⾅�P{�W�k�,�^�:vV�zS�oiV���^�B�k�	�{�=Q��-Î��  �  �g���/�5�/�P�:�j��"���ꆽ�M�������]s���W�h:��c �/)��;
������&�[�B�X�`���{�����0����-�������&k�rcQ��7���v���>�RAļ����O���u���`���]���l������<���ſۼ�!�Y���H/�f�I�
\d���|�c���s���O������+t��3W��9��"��e����r ���6���S�CKq�k��������d��������h��M���3��v�h	����ifƼrR��QV���ሼ����l������E��{�Ǽ�r鼹���V��95�MhO� 	k����������aW��5���0��H���؁m���R�j?�vm7���<��N�*�i�����;d��L�������m������>5�������w�)�^��$H��4���"����7x�����v|�i��#��=�"������/��C��dY���q�h���Г��젽oܫ�GᲽ}���[L��೦����@���}�ϯm�5j�2�s������8���좽�ܰ����㥾���������Ӫ�QO��ׅ����xu��b�"yR��D�ɱ9�i2�jR.���.���3���<��FI�τX��j���}��ꉽC-���]��W��������gƽ]V˽��ʽC�ýG'�� ����嚽(뎽;��Ҧ��Xэ��L���ͧ�A}��T�½��ɽ�Y˽cǽ������aۤ�X����������4n��f]��O�߀C�~�;��7�q�8�Ɯ=���F��\S�+�b��bt�VB�������8��Q���|ض��x½��ʽ�ν b˽Ný�G�����;����@��皊�o����䔽�ѡ�?ذ�9����ɽ�sϽ�Ͻɽ��������V������d挽����l�r���b�s�U��LK���D��B�8�D�2�K��V�԰c���s��<���  �  �����#��>��d�������V��'k����������K����l]���=��)��#��,-�hoE�^g���������%+��Aw���������f���y{b��p=��K����u�ʼ���Nׅ��M^�Sg?�7�.��,�P�8�d�R�j{�on���'���,꼿���\1��U�7�{�]e��\K��3��ה���B��ۓ��JX~��Z�_&>���-���,�ī;�FiW�@nz�#ڎ����4G���ϥ����\z���G���%[���6�b'�0:����ȼ�'�� ��<~s��^�Z�W��_�F�v��������lɼ�����1�L�T���z�����l���q5���'���d���C��)���"T���r�"OZ�!SP��iV�g�k�����ʘ��g�������⽽�V���r��!����Y���怽��^��c@��'�Z��~��+���� ټ�gؼ>�޼/��s� �<���7 �h/6�LQ���p��v�����',��yݿ��Pʽj�ͽMɽ���������� ���zÃ�kf��G������=T��9��-�Ƚ��ӽ�w׽iӽ�Ƚ�Ҹ�Ϧ�������K�k��lT��GB��4�c�*�YY$�˪!��w"�]�&�^.�f�9��%H�S�Z���q��ǆ�g/���s��1S���ͽu�۽ł�z�㽙fܽ��ν�)���j��&��������2��9���ʁ������̽��ڽ�-�j��k�ܽj|Ͻ�L�������R��x刽��u�&_�D%M��=?�i
5��w.�L�+�x,��:0�g�7��`C���R�#�e��!~��ƍ�Gޞ�=���+LĽJ�Խ"0��潷��A۽��˽����1��خ������p��8h��x����Ž�"ֽ��L�轉�潄�ݽ
�ν��C������k	���x��c���R��.F�pQ=�f8��j6��H8�¹=���F�D}S��d��y��  �  b	��oz�F�J�nZy��K���n��//��w_���E��|�P����z�v�V�t�>���7�SNC��_�z߂�����'���:����M��K`��^C��`���Tu���G���Mc�����󫑼wd���8��w��,�b_���?I.���T��)��=�����߼���(8���d�D����^��I���蔺����}k���ã�����־v�۞U�ĴB���A���R�-�r�[y��kơ�>���@���Y��K\���䡽����E$k�!|>�V��M�B���"@���q�')O�;�<�^�7�V�?�T��:w���������wo伏���3��I^��y����粽\g½l�ɽ�MȽ/뽽����y���(��p�p��e�6�k����}��O墳�����̽)�ӽg[ѽ�ƽ1���8��tm���d��?�!��>
��|�T�ܼ��μG`ȼUȼDiμ��ڼ�8��ib���/��O��;u�R�������پ��0ҽ�,߽L���޽t�ѽ6����{��d왽/���j���=��6���Ԛ���ʽi�ܽ*h�$>����	ڽ?�ƽ�1���͙��j��rh��CM���8�T�*��!�ہ�d\��E�^!�t#%��/��n>�RR�~ql�ú������H밽W(Ƚk�ݽ)��T������������ͽ%L��q����0�����3/������G˽�߽��Q$���F���Q���߽I�ʽՊ��&&���5��G>q��'W�'�C��{5�|�+�3�%�^g#���#�!�'�K�.��9��-I��{^��~z�<͎�����;{��d�ѽ�/�bV������ix��
�ｪ6޽V�ɽsG��f姽rl���#������r���EֽF���;��<�������^+���ݽ��ǽ�Ͱ��*��^���r�[mZ���H�w�<�Y4�]�/�:Y.���/���4��8=��I��+[���r��  �  A���-n$��T� ~���ӝ��B�������fƽ�����q��fӝ�*T���#g�0M�d�E��R��;p�(��*�>Ϸ�(�ĽYGȽ���}����S��ہ�˛P��"�%W��F��v���|�O�9%$� P	��-������)��a�D�?�^�x�v?���ݼӶ�Z�>���p�>h������@
��TLɽX�ʽ'���t���iܚ������@e���P��O�n'b�j��Vd��^���|`���@ʽ�(ʽ� ���������"�w�_�E��a�e�G���Ɖ��"]�Po;�*��6&��$.���A�BCc�/���歼�j޼�.�QA7�Z�f��`������"��=gн��ؽ?=׽4�˽cc������莽޴���r�z��	���%���w���b˽o�۽}��&�߽�ӽ�྽�V��п����i��0@��/��t��ҼA-żh8���t��Tż�&Ѽ
��&���P4�k�-���O�*6z�4����ۯ��cɽ�߽���L����	y߽�R˽?Y��|'��䶕������q���-���ؾ�U9ֽ����4��-�������`��sнm\��56���\��ah��bJ�>s4��o%�������C������i�� ��t*��9���N��j������ԝ�=ٶ���н=*�^h��P��bf����������ؽ��½���0��;���m߮�R5���1ֽ�_��9��R��	�G���|�뽖�ӽ�˹�{����t���&p��S���>�M0���&�MD!�p���m�n�"�ތ)�k4�>�D��i[��z�Q��������[��@<۽�P�Z��������������a1Խp���[���Q���A��C����˽���.*���i�
��"#��6�� ��Z�Ͻh"���睽��p��^V��C��c7�(r/��%+��)�o+���/�N8�u�D�)�V�`cp��  �  ������&�W�X�0a��~����ݷ��ƽ�˽�,ƽ�9������Ί�<�l�|R�1^J��2W��@v�~ǐ��:��-����ʽ�ͽƽc�������-T��#�m���R��������I�Գ�?>����-�� ����Qd9�7�r��8��s�ܼ3���]A��/u�E���\ծ���½j�νr�Ͻq�ƽ�P��Fɞ�t뇽ͽj���U�J{T�čg������=��\���nŽ�Ͻ�oϽ��Ľ纱�����d|�H������鼊=��������V�G35�K$�έ ���(��<�v�\��b���9��'�ܼqe���8���i�q��(��`pýWhս�=޽��ܽ��н�Ž��9��!����y��U�w�G�T������?����н���c4轊�2�׽/�½�T���Ǝ��k�0�@�ѥ�	��d漄[ϼ�¼S��c����t¼yμq��C���-�?�P��K|�م���*6ͽ��Ʒ�����A��yϽ�Ҹ�����:��`���p��(-��lt½Ղڽ�ｦv��� �M������CԽS���럽�6���h���I��3���#�'H�p�nQ��M�E������(��8�r�M���j�gA��#%�����tԽwC�� �}j���]���]�i�ܽD�Ž>��Z������a���hýGڽ���ģ�w�����j����~�ֽ%��,!��o���p���R�Y=��.��;%����t��Q� P!�^�'�3�2�7C�֢Z��Kz�WK��7S��3�ý'�޽�����&�(b��U��H������׽z½B�����������{��W�ν���"���� ���	����� �x����ҽ�)��D	��'T��0�o�?9U�1gB�Z�5���-��)��{(�c�)�n.�Us6��C�.�U�i�o��  �  A���-n$��T� ~���ӝ��B�������fƽ�����q��fӝ�*T���#g�0M�d�E��R��;p�(��*�>Ϸ�(�ĽYGȽ���}����S��ہ�˛P��"�%W��F��v���|�O�9%$� P	��-������)��a�D�?�^�x�v?���ݼӶ�Z�>���p�>h������@
��TLɽX�ʽ'���t���iܚ������@e���P��O�n'b�j��Vd��_���|`���@ʽ�(ʽ� ���������"�w�_�E��a�d�F���Ɖ��"]�Ho;�*��6&��$.���A�(Cc� ���	歼�j޼�.�EA7�N�f��`��������6gн��ؽ:=׽0�˽`c������莽۴���r�z��	���%���w���b˽t�۽���,�߽�ӽ�྽�V��׿����i�1@� �/��t��ҼI-żm8���t��Tż�&Ѽ �����H4�b�-���O�6z�.����ۯ��cɽ�߽���G����y߽�R˽<Y��z'��㶕������q���-���ؾ�X9ֽ����4��-�������`��sнt\��;6���\��#ah��bJ�Gs4��o%� �����H������i�� ��t*��9���N��j������ԝ�=ٶ���н=*�^h��O��bf����������ؽ��½���0��;���m߮�R5���1ֽ�_��9��R��	�G���|�뽖�ӽ�˹�{����t���&p��S���>�M0���&�MD!�p���m�n�"�ތ)�k4�>�D��i[��z�Q��������[��@<۽�P�Z��������������a1Խp���[���Q���A��C����˽���.*���i�
��"#��6�� ��Z�Ͻh"���睽��p��^V��C��c7�(r/��%+��)�o+���/�N8�u�D�)�V�`cp��  �  b	��oz�F�J�nZy��K���n��//��w_���E��|�P����z�v�V�t�>���7�SNC��_�z߂�����'���:����M��K`��^C��`���Tu���G���Mc�����󫑼wd���8��w��,�b_���?I.���T��)��=�����߼���(8���d�D����^��I���蔺����}k���ã�����־v�۞U�ĴB���A���R�-�r�[y��kơ�>���@���Y��K\���䡽����E$k�!|>�V��L�?���@���q�)O�&�<�C�7�4�?���T�T:w�߲������Po�y���3��I^��y��󝽵粽Pg½a�ɽ�MȽ&뽽����t���(��l�p��e�8�k���~��U墳�����̽4�ӽs[ѽ�ƽ>���8���m���d�?�,!��>
��|�i�ܼ��μO`ȼUȼ?iμt�ڼ�8��Yb���/��O�;u�F�������پ�|0ҽ�,߽@����޽l�ѽ/����{��a왽-���j���?��:���ٚ���ʽq�ܽ4h�/>����	ڽL�ƽ2���͙��j��#rh��CM���8�c�*��!���m\��E�d!�x#%��/��n>�RR�~ql�ú������H밽V(Ƚk�ݽ)��T������~������ͽ%L��q����0�����3/������G˽�߽��Q$���F���Q���߽I�ʽՊ��&&���5��G>q��'W�'�C��{5�|�+�3�%�^g#���#�!�'�K�.��9��-I��{^��~z�<͎�����;{��d�ѽ�/�bV������ix��
�ｪ6޽V�ɽsG��f姽rl���#������r���EֽF���;��<�������^+���ݽ��ǽ�Ͱ��*��^���r�[mZ���H�w�<�Y4�]�/�:Y.���/���4��8=��I��+[���r��  �  �����#��>��d�������V��'k����������K����l]���=��)��#��,-�hoE�^g���������%+��Aw���������f���y{b��p=��K����u�ʼ���Nׅ��M^�Sg?�7�.��,�P�8�d�R�j{�on���'���,꼿���\1��U�7�{�]e��\K��3��ה���B��ۓ��JX~��Z�_&>���-���,�ū;�FiW�@nz�#ڎ����4G���ϥ����\z���G���%[���6�b'�.:����ȼ�'�����&~s��^�4�W���_��v��������lɼ���c�1�*�T���z�w���[���`5���'���d���C�����T��|r�OZ� SP��iV�p�k�����ʘ��g�������⽽�V���r��3����Y���怽�^��c@��'�r��~��+���� ټ�gؼ7�޼��f� �*���7 �N/6�.Q���p��v�����,��gݿ��PʽZ�ͽMɽ������������xÃ�jf��I������ET��C��9�Ƚ��ӽ�w׽)iӽ�Ƚ�Ҹ�,Ϧ�#������k�k�mT�HB�1�4�u�*�hY$�ت!��w"�e�&�^.�j�9��%H�U�Z���q��ǆ�g/���s��1S���ͽu�۽ł�z�㽙fܽ��ν�)���j��&��������2��9���ʁ������̽��ڽ�-�j��k�ܽj|Ͻ�L�������R��x刽��u�&_�D%M��=?�i
5��w.�L�+�x,��:0�g�7��`C���R�#�e��!~��ƍ�Gޞ�=���+LĽJ�Խ"0��潷��A۽��˽����1��خ������p��8h��x����Ž�"ֽ��L�轉�潄�ݽ
�ν��C������k	���x��c���R��.F�pQ=�f8��j6��H8�¹=���F�D}S��d��y��  �  �g���/�5�/�P�:�j��"���ꆽ�M�������]s���W�h:��c �/)��;
������&�[�B�X�`���{�����0����-�������&k�rcQ��7���v���>�RAļ����O���u���`���]���l������<���ſۼ�!�Y���H/�f�I�
\d���|�c���s���O������+t��3W��9��"��e����r ���6���S�CKq�k��������d��������h��M���3��v�g	�}��cfƼhR��DV���ሼ����l��귕��E��G�Ǽ�r鼗���V�|95�#hO��k����������NW��$���0��<���ām���R�j?�um7���<�'�N�;�i�����Id��]��������������T5��-���'�w�R�^��$H�4��"����Jx� ����|�l��#��3���Ь���/��C��dY�ѷq�S���Г��젽Yܫ�3Ჽj���JL��ѳ�����@���}�ȯm�5j�8�s������8���좽�ܰ�����������#����Ӫ�gO��텑�-��:xu�7�b�AyR�1�D��9�|2�zR.���.���3���<��FI�҄X��j���}��ꉽC-���]��V��������gƽ]V˽��ʽC�ýG'�� ����嚽(뎽;��Ҧ��Xэ��L���ͧ�A}��T�½��ɽ�Y˽cǽ������aۤ�X����������4n��f]��O�߀C�~�;��7�q�8�Ɯ=���F��\S�+�b��bt�VB�������8��Q���|ض��x½��ʽ�ν b˽Ný�G�����;����@��皊�o����䔽�ѡ�?ذ�9����ɽ�sϽ�Ͻɽ��������V������d挽����l�r���b�s�U��LK���D��B�8�D�2�K��V�԰c���s��<���  �  ���Ԗ&�6���D�	MR���\�ȸa�3�_�C�U��MD���-�nD�q��-輯��N�����8��5���K��*\���d���e�&�_�~XU��H���9���*�:��J������<ռ����a}��}ے�娐�B<���b���nʼ����Y����'���6�	�E��T�`��"i���k�7g��2Z�*�F��/�|��f�������0�Rc��},��7D�l|X��<f�Gl�h%j�b/b�HV��XH���9��*�E�x���:����ؼ�ᾼ�Ҭ�u�����������ԼN���A�����w1�|�B�7S���b�<�q���}�x͂�tj��!��t�q�T�]�zIG��`2��W#�lc��!��0��lF���_�Ex� ��|2��*K��ɯ���P���B����v��qh�{�Y�D�J�iZ;�v�+�.������
�A+	�.u��P�y�%���6�9�H�j|Z�Ũk�Y*|�������� ������&Μ�,���q���*��*w��Acr���^���R�j0P�DX��i�����'\������ǡ�z����~��7�����E����ْ�.͋�����)xz�Zk�}\��,O��E�C�?� �?�A�E�s"Q�i`��q��L���Ӊ������ڙ��u��d����î�e��QI��Ǳ��B��]��k����̉��J����u��u���~�������'���\!��v��1�������(��*:���?���Ԛ�+7���a��>D���u���e��W���M��H�k�I�>P��[���j��e{��'���d���Z��c�����Ǡ��a���嵽�&���v���᪽IR��^u���e��l<��R-{�<h~��Ʌ����� ��pȧ�� ��Pල������������˫����9O��Ƕ��ލ�⾅�P{�W�k�,�^�:vV�zS�oiV���^�B�k�	�{�=Q��-Î��  �  ��4�qM=�\DB�i�D�B�D�6�B��r>��Y6�*����q�����ɼ�4��+����๼��Ҽ=*��.��� �t�0�ǜ<��kD���H���J�?�J�^H�AC�r:�Iz-������	�&���м�,�������ǼCN����o���(�m�7�PC�ZJ���M��\O�T�N�h�K��$F�Ҁ<�]�.�}X�H2
�v����Ҽ<¼�\���7м-)�'�xa�g-��];�8�E��K�UO��P�EO���K���E�ܾ;�J�-���_d
��1󼿂ڼ�~ϼ��Լ�p�wl���[�.�'�A��Q�S�[���b�&�f��xh���g��e�)�^���T���F���5�Y�#�*����H��A��@��%��9��fN��|`��n�΅x���~�N倽]e���߀�o-~�'Fw��hl�]�]�BTL��:��++�!�88�8m#��0���A���V�;�j��7|��ф�f��d(��⋍�B፽�,��h&��@e������at��wb���P��EB�K9���7��]>��L���^��ps�Ѱ��W(������ݖ��r��R���3
���I��y,���H���c�����{���j�;L]���U��NU���\�.Ak���}� ��͐���\���	����������AH���@p��zo���������������s�� e�;�\��W\�P�c��q�x遽�����o��@���� �<���8����!��z���H���Ԡ�����z��r������Wr�a�d�2^�_���g��w�݄�����cN��{A��� �����)������0}�������B��PӜ�)[��)Z��Xۂ���t�;h�Y�b�6(e��Bo�5�'��/Β��S��?�������VE��0����檽(+��E'���m�������疽j���QR��x�d�l���h��tl�U�w��3������ m�������  �  ��]�6 `��C[�+VQ��lD��6��<'�����/���u#ϼO�������/T���K��8��ɟ�_麼�ۼ�����I�����B/�@�>��GM��@Z���c���g�^wd�kY���F��/�#�}d�4v��,�3������=t&���>�H�S�� c�X{j�d�i��c�i�W�,J�4W;��',�b��@Y�`t���ּ����˓��V[����������-����Ӽ��m�
�����*���9�x�H�S�V�u�b�!�j�oll���f��X��#E�M>.��h����o) �_��!�,I%�˲>���W�4%m��G{�����w���w��\l��_��P��rB�Z�3�R$�#��7`�����ފ伻`߼��R"����	��z��z,��t>�(�O�k`�_�p�� ��c���Ì������������6���s�b�\�e�H�|�:�ɢ6��<���L�ȫc�G)}�Ç���֓�PX��dĚ�w���䓽񦍽A������cp�/Ta���Q�ĚB�K�4�;�)��o#�-�"��(��2���A��S��1e��w����!Z���b�����a䢽,�����-Y���?������쐽�녽��y���n�dn��w�����'ϐ�/@���1��t ���ϳ�롳�.��'�������L&���u�������[����w��xg���X���M��fG��G���L�n%W�7ve���u�<��n���X��Q��ɍ��E���J���cq���<���*���"�� 럽�����������v�_x��ρ�А���o���D������r��wε�wk��e&�����������;���@���&��|�w�+h���Z��vQ�!|M�OiO��W��[c���r��́�LE���}���p��#2��~����������'��6���{g���A��2]�����o̊��O����������[������=��ǣ���u���  �  mW��%�^~��-i���O��m5��4��H��ἊA���I��p{���5d��#M�hG��bS��vp�[T��#���t�˼��D�~R&��@�_v[�Q�t������~���ފ�;D����t�6�X�kL;�g["�����(�	��V0���L��j��-���y���������KP��`�k�SSQ���6�=�o��q�輎ƼgE����h}� �j�\�i��Jz�f����f���¼������/��W4��N��-i�,����o��্����=ʄ���q�1U��{9�rJ$����;��]-�=�G���f��ӂ�����O��;v��pڒ�������{��$b���H���1�:v����������߼T̼���������üf:Ҽ��w�������&��<��tT���n�����Y��ŝ�0����,���㤽����L��w��I*h�PdV��P�X���k����������������������"��<ȟ��R��vZ���s���]��J��$9�<�*�>��N��;!������2�O�+���:���L���`��
w�T����a���0���.��强��!��^	½�
��첽����2����ދ�:���)��9��`������i���u��L�ȽƗ˽FȽ����Yf��B?������샍�'I����p�T?_��/P�]�C�;��b6�6��;:�ˉB�dgN�/]�;n��ွ��7E��6����Ʋ�f���9�ǽX�˽�ʽ��½�N������~S��,��5n��yF��,����Ӝ�V����2����Ž�0̽��̽��ǽ[��ٱ���������>Ջ��8����o��u_���Q��F�|�?�
�<�%+>��	D���M��[���j�Q}��Ј�pm���9��o���,ͻ��ǽՑν��н�Oͽ3Ľ�޶��������!���������Zڙ��T���o���GĽ�Tν�  �  [i��4���8�����b�1�=�a�� ��!�Ƽ�l����}�5HN��6-���� O�� ��78�U�^�������Jؼ���B�&���J���p��v���6��S�������b���u��pQ]��"?��x,��)�n�5���O�jTr�l$��7M�����������៽����悽��`�5�;���|����T˼q���Sd��@e���G�f�8��28���E��Ea�L���&.����Ƽ������K�7���\�����:��QM������U��e��lێ�B#{��iY�y�?���2� Z6�9sI�]�h�����`��"��������|���觽�^���7����m��xJ�9+����t��W7ؼ<���ѯ��Ӧ��$��ԑ��_��G�ʼʃ�A�����3�	+R��u��鍽X����������(��
��tƳ�:g�����V@��n�p��Ri�vr��Ą�)���Xo��C���f�Ž �ʽ��ǽ�ڽ�ϰ���Ŝ�~d��ύr���T�z<��:)���������Տ�p����	��=�?@�P�*�k7=�hT���o�YA�������@L��oϽZ�ؽ�K۽V�ս��ɽ��������TW��ܺ��0�������"1���޶�G2ɽ��ؽ
<�	L�6�޽�Fҽq����㮽�\���u��@�y��b��O�8B@� 35�e�-�W�)���)��-�C�3�v�>���L�N_�r�v��s���������Q���sнݽ�:�5Q㽬�ڽ�Z̽벺�ha���㛽>������؂���h����н�_޽�r�����ܽ�ν+���w��r���ш���&v��[`�&0O��B�\�8�e�2�i^0�`�1��p6�$�>���J�|�Z�Oo�W���A��x���-���&ʽ�Hڽ�����~q�1�۽��˽J��w���?��T홽����$������3˽�۽�_��  �  X���������Ow��9I�0������a���Ry��շV��"(���	��*�.��E���,��58�A"m��P��?�̼���jj,�#�X�k����ʙ�j	���u������v��v���Qz����y��4W�Y�A�)�=��GL��Cj���������������~]��:泽�����4�q�˪D�������2��~���g�i�'�?�fQ%��[�u��Q#�?<��Md�$��x!��}:켪��q@��m�����*΢��������=��&豽u�����9t�FKV�՝G��NK���`�M����������伽�tŽ'�ĽE�����"ϔ��+|��P��*�1�������ļ�Ĭ�B���N���_����)������ⷼk�Ѽ�s��3��U0�xaU�<��G���w�����½+ѽ�׽�ӽ_ȽQT���9������W���}�vჽ\6��%������r�ͽ�A۽���ܽ��Ͻ���M馽a8��kzv��R��5�(A �=���K�e �ͱ��O������N�����.!��4�NVN�+�n�6��Dq����w�Ͻ#G�n(�6R�T�8�ݽ\�ʽ����p��r���'����gt��x�ƽ2�۽�\�m'��P��t��uJ㽺�ν�����ڠ��O��<v�#�Z�ѫE�y6���+�(%�^�!�|�!�ā$���*�8�4��\C�sW�	r������$�������˽��V=����+C��Һ��!߽��ʽ۶��Y��#a��J������ň��н#'�՜�3q�����.���u޽��Ƚ��������#X���p�H�W��E��Q8�n/�C9*� J(�(h)���-��h5�'%A�b�Q��h������ה�-��.8��� ؽ�콂������"/��e�E�ݽFɽt��>���E������J;����ǽ|�ܽ��ｓ���  �  :]Ž�F���ɱ�|Y���1��z�R�zo#����J���#烼�_B�������L�λaȻmػ�} �R�#��0Y��]����ȼ�D��)2�$xc��؋�����=/��TƽhɽP½�2��n윽ȉ��W?g���O���K��O[���{�܎���������ȽDʽ��������7t��Mi���L������`ӵ�����F�T�ކ+�c_�L^�P�����(�m�O�;���MN���\꼀u�zkG�D�y��ږ�d�������|ʽ�1ʽ,��3:��5a�����Vte�#bU��>Y�U�p�����Wפ��@J˽�tԽgӽ[Ƚ�Q���c��݃�{W�h�,�7
�X�߼,꺼�^���������z�������������Ǽ�켳���0�K�Y�ӄ�����=Ӹ�1XϽ�E߽J�.���ս4h½�g���o��᥊��څ��������t����Ž�۽���֓�d�꽰�ܽ�{ǽ��������({��)S�w3�}����/+��b�������W���Lo�8���?�g�0�ŀL��@p�h󍽃�|_���ڽ$p�1����0 ��������9Eֽ����]��������������N��SUѽ�;轆m�����w�rA �iN�D$ؽ�R��	ڤ�mꍽ�uu�`VW��A�$O1�W�&��l ��W��%������%�p�/�?�>��T�1q�,M���١��#���ս{�콅����S�~�������ћսeۿ������P�������k��C�Ľ�Z۽�5��b<��b�g-����齂_ѽ����ٞ��@���=o�1T���@�^#3��x*���%�a�#��$�>�(��J0��<�\CM��ge��Â������Ƚ":�Ǌ��T�f`��z���0��tӽ)ﾽ؎���&��>ï�P���0�ѽV�轋^��A���  �  �H��^B��0�5l�9Ｆ���?�i�����v]���9��&;�A�;��;�ٰ;;n�;^ש;i��;�];��:Ұ���[����*�h����ȼ�o�t8#��r<��]L�`P���G��4�$�����;�Ѽ�ݴ�򿯼�SüS���X���+���B��P�9�R���H��y3���T���꯼��n�:�8?��������`:�;�,D;�Z;�rZ;t�E;��;5K:�L��𛈻�u
��5f��ꪼ�����*2���H���T��T�s�H��3�YS��b��Yؼż��ʼ�������)�^F�]�[�1�g�Z�f�ݐY���B��%��l�.SѼ����[�h���+�K����һ�������1���Z�ƻ�6��Z���%��iR��������dw��11��vQ�?�m�[������"F���{w��Z`�F�
.���^$�/���1�!�K���h�7���YǊ�]��	���.���l�S$N��.��-�_���μ_���^��t�	���g��c����������h���f��b׼������}.�;�M���n��@���C�����,2������^���s��[s� S]��NP���N�+�Y�Wo��,���F�����E���m��*N�� ̗����cs�B�S�|7����<���� ��X（��)sݼٔڼvnڼ��ܼ��h�����E�����4�B�P��p����o���&᡽�䧽󼧽����������/�w��c�ZX���Y���g�oT~�v挽�8���z��s��������s������.���mNm���N�m24�϶�����I�2�����|��
�#�#��q�����*�<�-���F��Bd�N9������㟽`���z���V���x���0���
�����z�0Ji���b���h���y�R]���P��&𳬽�  �  �EB��O<��A+����R輰)���e����cab�jB��;�R~;�#�;�-�;��;��;�%�;=�N;�K�: 麺8ݫ�S�(�1凼�ü� �ׇ���6�n6F��J���A�wN/��N����`�ʼrܮ��䩼;����<���W�&�=���J��L�ЬB��[.��������3���dk���P����|º�':��;��7;p�N;O; �9;�	;#�E:�����-l
�_$c�Yr��h��l��)-���B��N���N���B�j>.���������Ѽ�<���żS�u��	(%�1�@���U��Ma�Y�`��S��=�3�!�����Rμwm��Ei�e+.����ڻ[w������$���m̻�����	��;)�
LU�&ψ����%h�[\���-��M��/h��o{���*����q��L[���A��*��z��;�!��.���G�_�c��b}�����5������^d��*h���J��,�!�[#��μK|��E������Y���XΒ����&���.��1v�����ܝؼ��������-��iK��ak�V焽)x���������}���ޏ����	o���Y��HM�QL�0�V��Gk���騐��!��6!���H��d\��u<������hp��R�ǜ6����k3�<d�B"���a�޼�ۼ=�ۼ�u޼i�伧��@5 �Љ������3���N��/m�=���/������ä�����0���s퓽Mچ��s�I�_�]iU��V�Z-d�az�ԋ���}��Pt��}r���s��"������8���F�j�tPM�2�3�����1�k ��v��kV𼣓�%$�q�|��������0h��w��|-�ߢE��)b���������;������!����k�����d��tՇ�Xw�}0f���_�@xe�-v�vD���Ԕ����ߜ���  �  ā0�l[+��6�$���ּ���/�Y�X��gx���%�'�:��P;lN�;�^�;2�;ِ;��q;� ;&U :!���<���b%�����@�����v���P'���4��B8�&�0���������fo�����6��	ժ�9ϼ����,���n,���8�;��>2��& �	����ؼޡ����c����g��k����ǒ�:��;�/*;2�*;�;ķ:��:8�8 �8��g�Y�\�M���]�Լo��F��2�2=�G�<��32��C�/���`⼋_�������7����ϼVw�����P,1��D�h�O�i5O��(D�q�0��������Ƽ7��3�l���6��?� V�k%ջsdʻ Iλ�߻H�������4��>_�nы��@���Jݼ���4%�_!A��dY�o�j��'r�r�n��qa���L��5�)R �������n�$�P�;���U�nWm�)~��W���"��R�q���[�ʴA�R�&��-�ta�+pѼ�Y��_ר�oe���ޘ��u��E��� ���=o��:#����żC
ݼ��������)��D�n�a��|�,���F�������ޏ�3���kz�ȅc��1P�ڬD�`�C�(�M��`�e4y�7=���͓�AI���u���"������恽�dh��6M�4�4�U � �������F;�o 伟�༒]�k��.꼣V�����x���'62�zrJ�.�e����^;���ۖ�����?����*��Bi��*i���#i���V�h	M��|N���Z�%o�A܃�&����꘽����Ɯ�����z���C�z�c���I�{{2����Y�����?�������l�t�����F����j����:���T-�0C���\��{x�����ؕ�84��9�������8���ꍽ����H&m��\]��wW��\�$+l�8N��ȍ�����栽�  �  9��u�������&ֽ�!c��D�O����=U������"�9�F�:�&B;��h;c<p;e�X;�b!;�U�:��C���P�$�λ�T'�%@t����nӼ����U
�,���:��B�Z���較���I}�����.-��%���U��g�ؼ��������Db!�v��`�pa�z�ü�����_�%���Cǻ��a�u{��*wb8�s�:	b�:�i�:��:��9�'��ǺW�΅���o�_�Y��Ŕ�	��R1��!U�o�#�{�"��z����K�鼘A¼n���Õ�����L���ڼ?�N�:�+��5��6��-�|���	�2����V���!�x�VJ�̍'����5���^M�1"��I�Q��+T*�~�J��t�屓�xH��,2ټ�O�����{0�bRD��TR��>X�U�UI���7�*o#����r��� �c���M�)���@�)�U��kd�<�j���g��W\��J���5�{��G������2�ؼW�ü������Ϟ���Z���������!T��뾼��м|��(.�u��&���<��2T���j��
}�Qp��S���(��ϩx�%f�ZIR�ܠA� �7�7���?�ƳP�V@f��d|��}��dL������/H��+
��'At�h�]��G���3��H"��X�l	�D�Я���{�{Y鼑 �(��4���9 �N\�^��� ���1�o�E���[��Ir�9e��p.���8������ŉ�i<��n�m���X���H�@w@���A��sL��T^��s�tD��S�����,-���f���!��kq��[�/�E���2���"�,�,s������������c�����k���f���z,�_����.�NA��+V���l�_���9S�������dȒ�����<���Sq�Z�]�rP���J���O��,]���p��F��2!�����  �  ސ�c�i޼2Tż���5|��}�R����/�ڻO��� ���P��N4�:�k�:��;!�:^�:Ӊ��.H�3���l���8���r�G�����[ؼ���b��~G ��|�ڼ٭��+�����o���J���D��q^�@����諼~�ϼ�=� � �g ��켒�м�����ۑ�V�h���3�>������q�"����Q��D6����@�����Vh�F÷��s�1�qe��A��&��[:м� �2`�Ĝ���<��O�ݼ&J��2���p���4p��z�ݰ���b��ټ����~�����]���� #
�ݵ��ےڼ+��6V��3��9�n��M���2��`������T��v0��L��p�����	���L����ۼ�������sJ��Y-�}7�}�:�M7��-�[��������\��^�5��N����
(��9���F��M�:L���D���8��>*�t�����1��P�pUּ3�Ƽt�����rg��[���7�������zмHK�A���Û�L���%��66��GG�TW�jd�|�l��n�׶h��8]�X�M�@�=�??0��R(�(�'��/�O�=��O�eXb�b.r�\�|�W��g|��Kr��zd���T���D���5���(����y��A:
��9��}��98�����p���#��DZ	�u�����;'��e4�A:C�]7S��Bc�֨q�,X|�R���3t�C�v��#h��V��E��Z8��x1�J�2�~z;�QJ�[ \�/�m��K{�ډ���⁽��}��hr�+�c�	T��D��p6���)��8�K��������̎���������V�����6(�r4��eB���Q� Ab�&r�"��Bp���ꅽ�׃���|�@m�g�[���K�#T@�� <��@��KK�[�8�m�nO~��/���  �  &_��s��Ah�������A��>���Km���I�k�$��+��񻲻U�Z�f_׺�&�����˻q�����a��\mֻIw��V;��b�^��媖�����}��5Cļ_ɼS�ż�a��݉���d��V0W��i(����p��A>���D��{�V���7V����ƼnϼT�μ��Ƽ���4���������Ze�֋?���d��#?����^�ߣ&�N$���W�#k���&໡%�oc=�/�c�㘄�P�������/����ȼܦҼ|>ռ�μ�0���0��l�����h��gC���2���;���]�-g��J騼�Gȼ߫��������g��,��?�ּ��Ƽ�O��4���H���b���7�g��M�P�=��S:��D��\�G8~��œ�������8oռ�꼈&�����������L�s���Q�������"Ｆؼ}�ȼ��ļdpͼλ�|����ڃ��)�{0��&2�R�/���*��e#��f�`)�k�
�p�k���⼎�ӼH/ȼ
¼У¼�	ʼ��׼�7�������
�j��d� �P�*�d�4���>�kQG���M�oQ�T�P��K�5^A�z5��(��9��T��^�����*��8� �G�(&U��^�nc��Wc�\L_���X�VFP��]G��6>���4�K+�aw!�����S�����M��YO��{�9��6b ��<*���3�xM=��F��O��/X��p_��8d�9Ie���a�bqY��SM��J?�9�1��N'�4�!���"�#�)��5�q�C�)R���]���e��ah�/�f��a�nZ�pR�JII��Y@��;7���-�hO$��@�����Q�S"�1^�����'�3D"�1=,��I6�f@�C�I��	S��0\���d�vZk�61o�C�n���i�_Y`��zS��vE��8���/���,�H�/�3�8�p�E��OT��b�f�l��  �  �ⅼ����8��X0��8����З�/����m���zv���P��!%����㨻�xr��}Y��6���Q��

�k�8���e���V-��՚��|��Ä��2���S&��,X���.��`����`�T�4�(T	���˻����l��n��p�����&�KU�P���Ź��"?m����� 쮼0a��W0���v���9��s���i���;�q���ݻ�����ƴ�X<ػ�;�o8���e�i�����7������W���D鱼�������9����m��M|��ѭo�&�E�>��{�����*��6�AG���y�� ������7����ϼ-ټС޼)fἕ��V%߼$�ؼ��ͼ<*������H疼�:���r�q9k��v��=��՟����yҼ��7��������N�	���
�׍
��� *�Q\�����:)ڼ�Ƽ���oL��+���v������.�ռ�S＞/��
��l�b@��� ���"���#�`;#��;!��7�g���J�{Y��������Qiۼ��ڼ��� +��p.���j���)�l�1�͊7�;���<���=��Y=�:T;��=7��0��7(�vo�����t��m	���	�o��%���E#�ɡ/�d1;���D�`�K�<P�d|R�hS�US��aQ���M��"H���?�̓5�&*�T3�2������m�����q�(��J4���>�tmG���M��RQ��SS���S�*}S�=�Q���M�{�G��w?�S5���)��U�Us��}��8�����"�E�-��C9�ǽC�iL�P�Q�$�U�XhW�hX�pW�nU��~Q��1K�uB���7��,�A�"�k{�[���� ���)���4���@�u�J�(�R�{?X���[��M]�U�]�S]�7�Z�e�V���O���F�� <�p�0�eS'�� ��f��� �ז'��1��#=���H�ЃR��  �  �(C��Ni�1o��6���
��C���`7��S1��`����������bTI������n߻Sg ��A'���\�͔��Z9��!�� �ļ�ż�񾼦V��~����E����-[���5�(���{Ի�i���7��2��ẩ����}�k���V��#�.��U�.|��ϐ�f.��妴���üdμ��Ѽ�[̼�2���奼����[}\�Ss/�����]�e,�^�W�t{��\أ�����̼ixӼ�>Ѽ_�Ǽዹ�m����������h���D� � �����i.Ż�x��ᒻah���eͻ�����0�A ^�=Յ��曼4����ż� ڼF�켁<��6�ym�� ���� �ڼc��nB���a���Y�����������ƼW�aL����zb�RE�ѳ�X��o�����AX��&�漕�ռ*�ļޜ������ѧ��3���:ӏ�\��7���?k��Cgɼd�߼�����Z����h���/#���+�B�2���6�J!6��	1���'��[�ps�6l�[6���T��>������c*���8��C�"J�b�K��H��MC��#<�R4�LV,��N$��&�5�����V��Њ��U}�������y��m����k���x&���0�~�:��/D��xM��8V�0�]��b���d���a�O�Y�|0N��@�%2���&�(E ������%���0�v�>���L���X�c)a���d���c�4�^�۽W��]O�/�F��x=�VG4���*��/!�r�����I
�t3�!��"�����M�l!%��$/��8�lrB���K��T���]���d�Y�h�Hmi��.e��C\��O�"�A�+�4��+�̸&���(�>�0��4=�O�K��Y���d���k��n���k�Rf��^��lV�}�M��D��;��52���(�����������5��	�j��� ��*��"4�b*>��  �  r	��P�r��j:��&�Ǽq��(��d�������\Ӽ`�������b�:�8�~X-�EB��Xs��L��=|����߼ɞ���E����������̼ͭ��?���`���+�����Lt���:K�����qg��:G�!:-u�8���j�-��ᙻ�軕�!���U�����짼9Mȼ���������������|ܼ���}9��0?u�yJT�9�R���p�o��RԶ�N�ټŕ����h��� �A����μ�t���Y����g���5�`K���λ͓�leO����<���,���r��n��E���/$��S�6ʃ��;��ģ��z��$�����?��!����a��������Tм�ι�^=��X߸���ϼ�i������,���3�b4���-��F"����ܥ����NrѼ�����M�����*��,	����x�*�y�k4���x��V��Q��jb¼�ڼ���hV	�X����*���:��)H�~�P��YS���N���C�Y�4�r$����ߟ�8�
�`w����v1��KD�aiU��~a�E�f���d���\��TP�4�A��2�ع$�hf�1��L��w��e�Z�輭��y���J���5�Z�}���#���0�2�?���O��_�U�n��*z�����B��Qw��wi��)X���F�=8���/�sz/���6���D�@0V��g��v��~�aJ���n{��p�Yfb���R���B�0N4�Gv'�P�`��`|
�7 ��2��'�������nM������ �;�,�gZ:���I���Y��i���w��a���xy��Ty�j�ĜX�
H�&�;�c)6���8�/�B��xR�>�d���u��F��ǟ���h��(逽��u���f�'5W���G�_":��.�Ɉ#����r��C�h�	�����
�"�������Jq%��\0��  �  H5�/N�R	��˾���뼒��0�����R/�|� P������s����v�&�h�k뀼 l��C�Ƽ-P���ĺ�����r�"
��5�Oe¼/����Z�������Ae>���Y�'Y7:u��:�-;�];x�:Օ|:�,비)�����/�lG�������0�,����H=!���!��;�E	�~���߾�OM���g��"i��e���������o�X`�"���"�6V� �
�8o�ӿ��m���m[�`��b�лxɃ�O������0���
�-�|�0���%Z��Ŭ������X1�2�o��.��RYȼ�%��m��y�'��7���>���<�$�2�D�!�B�����ڼKϼ�׼�k�hB� $�D�9���I�l�Q��P�q�E�:5�Sa �s�
�y�HUȼ�F���ݔ��=���q��gb��P\��Z^�,h�M�y�޿�������ﯼ�lʼ���������W[6� �L���_�K�l��2q�F{l�ۙ_��3M�G9��g'�u�>���A!�Q>1�c�F�&�]��q�G�g������Ks�C
a���K�s�6��#�T���y����ԫ輲�޼cټ�f׼U�ټ�I߼��輤7��������j��5-��A��$W��m�Vw�������g�����5H��C'���o�|pZ��I��?��>�\�G�@DX�w7m�q�����hp��Ǝ�y��� Ă�#q��Z���D��*1� � �-u�1	��d������m��]�q0����5����Y�R��P�՟&�<8���L�Xac���y������H��F���
w���݊�rY�n���Z�6�K�)E�dH��?T�Jg���|�܉�����ܔ���y��b���\��}s��2]�(H�r�5��\&�'T�f��#
��T�������������G����d'��t(��  �  � ��{ Y�}���ݗؼ�]��2�r-�5�2���,��.�\���Lݼ�+��@����`������oA��B�뼒��tU$�f�2�ɉ6�0�/����Ns���ؼZ���Z�a�����f��+CӺ�:��;��=;':Z;�%\;��D;P�;MUk:Ŋ��iu����fG�i��%�ȼ{9 ���Q�.��:���;�T2����bD��-༪���(ơ�����%Z��\�ۼ<����ZJ1�*<��*<���1�����=Ӽ�᝼��]����wE��b+1�����8�B8��:��:�L�8*iF���D�|�ӻ1� ���g������Ӽ}Y���"�3<���N�8WX���V�I+K�L�7�l� ���
�c��4��W�����I�8�r�P�[ c�z~k���h���[���F��X-�mv��e��Ƽg��eԊ��(r�&A[���N��9J�xM��JV�JDf�o~�����v̥�^5ü��}���[&���B��Z^�-�u�ظ��{���Z	��gMw�=b��J��;6�y)�40&�7�.�c�@�3�X���r�߄�l}�������닽����Oq��W��<���$�"���U�*d켍Vݼa�ӼDϼIYμ�м��ռ{޼�뼈k��t�	��t��B-��+E�;`�t�{�슽!���
��P����Җ�1�������nk�B.W���K��K��pU��h�YQ���\��
��}q�����34��j{������<d�xI��1��\��9��o����9�3����\�va��4񼷉��_������$� �9���R��n��߄�s*��3��k����i������݌�^Ā��zj��JY��Q���T��b�%cx�z���(?��vʜ�����w랽���T���=��*e�wEK�(�4���"��Q��}�p��X ������������*�������Z	�2�$��  �  \���d���*뼉���_-�oy>�_D�E#>�!+-�������Ƽrަ�J����S��{�ѼW�w#�~�4�D�	@H�H@�l�-�>���86���Yk�/�|����ҁ�\��:e�/;��f;`;�>�;�k;�<;<_�:����S� ��ZtL�������ּR�
��'���>�}�K��M��UC�LH/�|��Mm��P_˼7���]l����Ǽ/�����-��(B�#�M�*�M�'�A���+�;��⼹�����c�Ј�3������u��k�7:���:��:�S%:Ic%��M��Q�T��1������)g��J����ݼ����G.���J��|_��j�Ηh���[��eF��-��������A�s��j*��FF��`��;t�r@}� z�a]k���S�4�6�������mȼ����5����f���O�Z�C�'�@��D��L�#�[���r�p艼��������m��c,�)L���j��m��5>��=~������4����p�V�� @���1��t.�U7���J�<+e���������;���ɗ�I>��O��w}���_��B�%%'����Pc��7��v׼Bμʼ �ɼ�˼��м��ؼ+�����H�����Q.��I��*g�r+��R���������	���bR��=��UM��4v��`�.T��S��^��s��ц��x��lO���A���C��2\��K?��T�k�o�M�H23�~r����/� ���񼵽缺'⼞�Ϳ�RT伈�뼂����>O� i$��;�t�W�Fv�����|W��Dv���\��w:���]���5�������t��Jb���Y���]���l�����}���#��l��[|��!���oџ�к��S��Urk��N��5���!�)�ڨ�D��~b��{L��ed��72�������L
����#��  �  $���i�vG��o�[��2�T�D���J�LD��2�����7���̼�����ԣ�q���ټUi��;"��{:�0TJ��N�"BF�R�2���bd�vI���oo����|���T���:��=;ngs;�D�;ի�;��w;ȔI;~�:.�$�_�J�""�u�N����Z;ܼBf��j,�t6D��&R���S�{[I�O�4��.� @����Ѽ����6R���hμJ-��oy�)t2��!H�?T���S��zG�4�0�����缒䩼��f�R�?���&��6Ѫ���l:��:��:x P:[�7�9���F�a5��w1�2�g�4)�����^���u2�ɱO��je��Zp�J�n�5�a�C�K�[{1�����������D�����'.�:K��;f�lWz��ȁ�H��X�p��fX�b�:��6������Pɼ����R脼cc�S0L���@�:�=�"iA�YJ�Q�X�M9o��/��I���K"��}�� ��*�.��O�^^o�N(���I��x����Ύ�>x���t��Z��C�ڽ4�\1�`o:�fN�~wi�9��揽`V��.�8��������b��D�f'(����E���I��f�ռ!x̼xpȼ�*ȼ��ʼyaϼD>׼�W�!��H6�����/�e�J���i�K������럽�צ�⫧� U����1���z���c�U%W��sV���a�Uw����Ț��#t���u���`��m'��Hו�#5���xn��mO�k�3��l��T�U- ���	漤�༡�޼�]߼���J�鼀���mM����f�$�E�<�AnY��Oy�ۭ���욽bk�������[���J���̖��:���x�0te��\�ړ`�Rp� ��鑽bힽM{��M������p������"׆�_�m���O�� 6���!��]����s� �n��������
��)���Uy��� �g@	����9#��  �  \���d���*뼉���_-�oy>�_D�E#>�!+-�������Ƽrަ�J����S��{�ѼW�w#�~�4�D�	@H�H@�l�-�>���86���Yk�/�|����ҁ�\��:e�/;��f;`;�>�;�k;�<;<_�:����S� ��ZtL�������ּR�
��'���>�}�K��M��UC�LH/�|��Mm��P_˼7���]l����Ǽ0�����-��(B�#�M�*�M�'�A���+�;��⼹�����c�ψ�/���t�����ސ7:�:��:�T%:�^%�M���T�[1�����p)g��J��u�ݼ���G.��J�w|_��j�ŗh���[��eF��-��������A�v��n*��FF��`��;t�{@}�
z�l]k�	�S�?�6����.���mȼ����5����f���O�h�C�/�@��D��L��[�}�r�e艼��������c��c,�L���j��m��0>��8~������0����p�V�� @���1��t.�U7���J�A+e���������;���ɗ�N>��"O���}���_��B�0%'����ac��7��v׼$Bμʼ(�ɼ
�˼��м��ؼ+�����H�����Q.��I��*g�r+��R���������	���bR��=��UM��4v��`�.T��S��^��s��ц��x��lO���A���C��2\��K?��T�k�o�M�H23�~r����/� ���񼵽缺'⼞�Ϳ�RT伈�뼂����>O� i$��;�t�W�Fv�����|W��Dv���\��w:���]���5�������t��Jb���Y���]���l�����}���#��l��[|��!���oџ�к��S��Urk��N��5���!�)�ڨ�D��~b��{L��ed��72�������L
����#��  �  � ��{ Y�}���ݗؼ�]��2�r-�5�2���,��.�\���Lݼ�+��@����`������oA��B�뼒��tU$�f�2�ɉ6�0�/����Ns���ؼZ���Z�a�����f��+CӺ�:��;��=;':Z;�%\;��D;P�;MUk:Ŋ��iu����fG�i��%�ȼ{9 ���Q�.��:���;�T2����bD��-༪���(ơ�����%Z��\�ۼ<����ZJ1�*<��*<���1�����=Ӽ�᝼��]����oE��G+1�F���)�B8(�:S�:\�8�fF�U�����ӻ� �B�g����y�ӼgY���"�<���N�%WX�o�V�:+K�@�7�b� ���
�\��2��W�����U�8���P�k c��~k���h���[���F��X-��v��e�9�Ƽ>g���Ԋ�*)r�KA[���N��9J�{M��JV�5Df�O~�����[̥�>5ü��j���[&���B��Z^��u�θ��q���Q	��YMw�1b��J��;6�v)�40&�:�.�i�@�<�X���r� ߄�t}�������닽����Oq��W�(�<��$�4���U�Id켨Vݼx�Ӽ'DϼYYμ�м�ռ"{޼�뼋k��u�	��t��B-��+E�:`�t�{�슽!���
��P����Җ�1�������nk�B.W���K��K��pU��h�YQ���\��
��}q�����34��j{������<d�xI��1��\��9��o����9�3����\�va��4񼷉��_������$� �9���R��n��߄�s*��3��k����i������݌�^Ā��zj��JY��Q���T��b�%cx�z���(?��vʜ�����w랽���T���=��*e�wEK�(�4���"��Q��}�p��X ������������*�������Z	�2�$��  �  H5�/N�R	��˾���뼒��0�����R/�|� P������s����v�&�h�k뀼 l��C�Ƽ-P���ĺ�����r�"
��5�Oe¼/����Z�������Ae>���Y�'Y7:u��:�-;�];x�:Օ|:�,비)�����/�lG�������0�,����H=!���!��;�E	�~���߾�OM���g��"i��e���������o�X`�"���"�6V� �
�9o�ӿ��m���m[�]��W�лeɃ��X���</���
�~�|�s.���$Z�0Ŭ�K���wX1�ʂo��.��Yȼ�%��O��[�'��7���>���<��2�3�!�4��ͤ��ڼHϼ�׼�k�sB�# $�X�9���I���Q��P���E�X5�qa ���
���}UȼG���ݔ��=���q��gb��P\��Z^�,h�0�y�ȿ�������ﯼ�lʼ[�꼪��j��8[6��L���_�.�l��2q�.{l�ƙ_��3M�:9��g'�q�>���A!�Y>1�o�F�7�]��q�G�t�����Ls�b
a���K���6��#�o���y� �������޼ټ�f׼g�ټ�I߼�輬7��������j��5-��A��$W��m�Uw�������g�����5H��C'���o�|pZ��I��?��>�\�G�@DX�w7m�q�����hp��Ǝ�y��� Ă�#q��Z���D��*1� � �-u�1	��d������m��]�q0����5����Y�R��P�՟&�<8���L�Xac���y������H��F���
w���݊�rY�n���Z�6�K�)E�dH��?T�Jg���|�܉�����ܔ���y��b���\��}s��2]�(H�r�5��\&�'T�f��#
��T�������������G����d'��t(��  �  r	��P�r��j:��&�Ǽq��(��d�������\Ӽ`�������b�:�8�~X-�EB��Xs��L��=|����߼ɞ���E����������̼ͭ��?���`���+�����Lt���:K�����qg��:G�!:-u�8���j�-��ᙻ�軕�!���U�����짼9Mȼ���������������|ܼ���}9��0?u�yJT�9�R���p�o��RԶ�N�ټŕ����h��� �B����μ�t���Y����g���5�YK�s�λ�̓�eO�0�����,���r�)n�������.$�S��Ƀ�v;��|���0���������>�w!����G��o�����<м�ι�Z=��_߸���ϼj������,���3��4���-��F"���� ����뼏rѼ����	N��:���*��B	����x�.�y�c4���x��:���P��;b¼Oڼ����FV	�4��э*���:�`)H�\�P��YS�|�N�r�C�D�4�c$����ڟ�8�
�ew�����1��KD�ziU��~a�e�f���d��\�#UP�Z�A���2���$��f�P��g��w����{��Ƞ�y�"��J���5�Z����#���0�2�?���O��_�T�n��*z�����B��Qw��wi��)X���F�=8���/�sz/���6���D�@0V��g��v��~�aJ���n{��p�Yfb���R���B�0N4�Gv'�P�`��`|
�7 ��2��'�������nM������ �;�,�gZ:���I���Y��i���w��a���xy��Ty�j�ĜX�
H�&�;�c)6���8�/�B��xR�>�d���u��F��ǟ���h��(逽��u���f�'5W���G�_":��.�Ɉ#����r��C�h�	�����
�"�������Jq%��\0��  �  �(C��Ni�1o��6���
��C���`7��S1��`����������bTI������n߻Sg ��A'���\�͔��Z9��!�� �ļ�ż�񾼦V��~����E����-[���5�(���{Ի�i���7��2��ẩ����}�k���V��#�.��U�.|��ϐ�f.��妴���üdμ��Ѽ�[̼�2���奼����[}\�Ss/�����]�e,�_�W�t{��\أ�����̼ixӼ�>Ѽ`�Ǽ⋹�n����������h���D�� �m���4.ŻZx�������g��	eͻ���^�0��^��ԅ�A曼�3��c�ż� ڼ��0<���5�Um�a �O����ڼ>��TB���a���Y�����ĭ����Ƽ=W�|L���b�xE��������������X��o����ռc�ļ������꧗�A���<ӏ�S��#���k��gɼ/�߼V����Z�t��@��b/#���+��2�ф6�&!6��	1�w�'��[�^s�*l�O6���T��D�
���z*���8�+�C�?"J���K�C�H��MC��#<�:R4�sV,�O$��&�T�����m������t}�������y��m����n���x&���0�~�:��/D��xM��8V�0�]��b���d���a�O�Y�|0N��@�%2���&�(E ������%���0�v�>���L���X�c)a���d���c�4�^�۽W��]O�/�F��x=�VG4���*��/!�r�����I
�t3�!��"�����M�l!%��$/��8�lrB���K��T���]���d�Y�h�Hmi��.e��C\��O�"�A�+�4��+�̸&���(�>�0��4=�O�K��Y���d���k��n���k�Rf��^��lV�}�M��D��;��52���(�����������5��	�j��� ��*��"4�b*>��  �  �ⅼ����8��X0��8����З�/����m���zv���P��!%����㨻�xr��}Y��6���Q��

�k�8���e���V-��՚��|��Ä��2���S&��,X���.��`����`�T�4�(T	���˻����l��n��p�����&�KU�P���Ź��"?m����� 쮼0a��W0���v���9��s���i���;�q���ݻ�����ƴ�X<ػ�;�p8���e�i�����7������W���E鱼�������8����m��I|��ĭo��E�"��U��>��i*�b6��G���y�u ��R���������ϼ�ټz�޼�e�A��%߼��ؼD�ͼ*������!疼�:���r�j9k��v��=��'՟�;���yҼO��������+��y�	���
��
�4��E*��\�����k)ڼ Ƽ��~L��.���v�������ռ�S＂/��
��l�;@��� ��"�q�#�6;#��;!��7�F���J�cY��������Diۼ��ڼ���7+���.�/��j���)���1��7�:;���<���=�Z=�cT;��=7�>�0��7(��o����
u��m	���	�x��-���E#�͡/�f1;���D�`�K�<P�d|R�hS�US��aQ���M��"H���?�̓5�&*�T3�2������m�����q�(��J4���>�tmG���M��RQ��SS���S�*}S�=�Q���M�{�G��w?�S5���)��U�Us��}��8�����"�E�-��C9�ǽC�iL�P�Q�$�U�XhW�hX�pW�nU��~Q��1K�uB���7��,�A�"�k{�[���� ���)���4���@�u�J�(�R�{?X���[��M]�U�]�S]�7�Z�e�V���O���F�� <�p�0�eS'�� ��f��� �ז'��1��#=���H�ЃR��  �  &_��s��Ah�������A��>���Km���I�k�$��+��񻲻U�Z�f_׺�&�����˻q�����a��\mֻIw��V;��b�^��媖�����}��5Cļ_ɼS�ż�a��݉���d��V0W��i(����p��A>���D��{�V���7V����ƼnϼT�μ��Ƽ���4���������Ze�֋?���d��#?����^��&�N$���W�#k���&໢%�pc=�0�c�㘄�P�������/����ȼܦҼ|>ռ�μ�0���0��b�����h��gC���2�t�;���]� g��騼[Gȼ��⼨���T����f�������ּ@�ƼBO��󷥼���3����g���M�3�=��S:��D�\��8~�Ɠ�����@��}oռ���&�����?�����L�����Q�/��ב��"��ؼ��ȼ��ļ[pͼ���\��������|)�X0��&2�)�/�u�*��e#��f�:)�H�
��o�4��[��k�Ӽ0/ȼ�¼ϣ¼�	ʼ��׼�7�!�����
������ �w�*���4�ؠ>��QG���M�.oQ�y�P�!K�T^A��5�0�(��9��T��^�����*���8��G�)&U��^�nc��Wc�[L_���X�VFP��]G��6>���4�K+�aw!�����S�����M��YO��{�9��6b ��<*���3�xM=��F��O��/X��p_��8d�9Ie���a�bqY��SM��J?�9�1��N'�4�!���"�#�)��5�q�C�)R���]���e��ah�/�f��a�nZ�pR�JII��Y@��;7���-�hO$��@�����Q�S"�1^�����'�3D"�1=,��I6�f@�C�I��	S��0\���d�vZk�61o�C�n���i�_Y`��zS��vE��8���/���,�H�/�3�8�p�E��OT��b�f�l��  �  ސ�c�i޼2Tż���5|��}�R����/�ڻO��� ���P��N4�:�k�:��;!�:^�:Ӊ��.H�3���l���8���r�G�����[ؼ���b��~G ��|�ڼ٭��+�����o���J���D��q^�@����諼~�ϼ�=� � �g ��켒�м�����ۑ�V�h���3�>������q�"����Q��D6����@�����Vh�G÷��s�1�qe��A��&��[:м� �2`�Ĝ���<��I�ݼJ��&���p���4p��z������b���ټ���`�����:������"
�������ڼ����U�������n�ˠM���2�s`�������T��v0�U�L��p�Ӻ��@��M��:�ۼ��������J��Y-��7���:�k7��-�)[����&����\��^�-��N�����(���9��F�mM��9L�j�D���8��>*�O�����1���?Uּ�Ƽ�s�����hg��[���A������{мpK�r���ߛ�!L�ؙ%�#76��GG�?TW�'jd���l�n���h�9]�p�M�T�=�Q?0��R(�3�'��/�U�=��O�hXb�d.r�]�|�W��g|��Kr��zd���T���D���5���(����y��@:
��9��}��98�����p���#��DZ	�u�����;'��e4�A:C�]7S��Bc�֨q�,X|�R���3t�C�v��#h��V��E��Z8��x1�J�2�~z;�QJ�[ \�/�m��K{�ډ���⁽��}��hr�+�c�	T��D��p6���)��8�K��������̎���������V�����6(�r4��eB���Q� Ab�&r�"��Bp���ꅽ�׃���|�@m�g�[���K�#T@�� <��@��KK�[�8�m�nO~��/���  �  9��u�������&ֽ�!c��D�O����=U������"�9�F�:�&B;��h;c<p;e�X;�b!;�U�:��C���P�$�λ�T'�%@t����nӼ����U
�,���:��B�Z���較���I}�����.-��%���U��g�ؼ��������Db!�v��`�pa�z�ü�����_�%���Cǻ��a�u{��wb8�s�:b�:�i�:��:��9�'��ȺW�υ���o�_�Y��Ŕ�	��R1��!U�n�#�z�"��z����D�鼎A¼`���Õ�����L���ڼ,�N�"�+�֝5�}6�ˏ-�]����	�������"�����x��UJ���'��������3M�'"�J�m��WT*���J�= t�����H��c2ټ�O�ܚ�|0��RD�UR��>X�)U� UI���7�7o#���r��� �c�{�A�)���@��U��kd�"�j�n�g�pW\���J�ݘ5�^��+�������ؼ/�ü���v�������Z��������1T��뾼Йм���?.���&���<��2T���j��
}�`p��`���(���x�9f�kIR��A�+�7�7���?�˳P�Y@f��d|��}��dL������/H��*
��'At�h�]��G���3��H"��X�l	�D�ϯ���{�{Y鼑 �(��4���9 �N\�^��� ���1�o�E���[��Ir�9e��p.���8������ŉ�i<��n�m���X���H�@w@���A��sL��T^��s�tD��S�����,-���f���!��kq��[�/�E���2���"�,�,s������������c�����k���f���z,�_����.�NA��+V���l�_���9S�������dȒ�����<���Sq�Z�]�rP���J���O��,]���p��F��2!�����  �  ā0�l[+��6�$���ּ���/�Y�X��gx���%�'�:��P;lN�;�^�;2�;ِ;��q;� ;&U :!���<���b%�����@�����v���P'���4��B8�&�0���������fo�����6��	ժ�9ϼ����,���n,���8�;��>2��& �	����ؼޡ����c����g��k����ǒ�:��;�/*;2�*;�;ķ:k�:8�8 �8��g�Z�\�N���]�Լo��F��2�1=�F�<��32��C�-���`⼁_�������7��v�ϼ?w�����A,1���D�V�O�U5O�|(D�\�0�ͭ�����x�Ƽ�6���l���6�X?��U�6%ջUdʻIλ�߻o�������4��>_��ы�A��!Kݼ���4%�u!A��dY���j��'r���n��qa���L��5�0R �������n�$�G�;���U�`Wm�~��W���"��=�q���[���A�=�&��-�Pa�
pѼ�Y��Hר�^e���ޘ��u��E������Ho��K#����ż^
ݼ��������)��D���a��|�7���P�������ޏ�;���kz�ԅc��1P��D�g�C�-�M��`�h4y�8=���͓�BI���u���"������恽�dh��6M�4�4�U � �������F;�n 伟�༒]�k��.꼣V�����x���'62�zrJ�.�e����^;���ۖ�����?����*��Bi��*i���#i���V�h	M��|N���Z�%o�A܃�&����꘽����Ɯ�����z���C�z�c���I�{{2����Y�����?�������l�t�����F����j����:���T-�0C���\��{x�����ؕ�84��9�������8���ꍽ����H&m��\]��wW��\�$+l�8N��ȍ�����栽�  �  �EB��O<��A+����R輰)���e����cab�jB��;�R~;�#�;�-�;��;��;�%�;=�N;�K�: 麺8ݫ�S�(�1凼�ü� �ׇ���6�n6F��J���A�wN/��N����`�ʼrܮ��䩼;����<���W�&�=���J��L�ЬB��[.��������3���dk���P����|º�':��;��7;p�N;O; �9;�	;"�E:����.l
�_$c�Yr��h��l��)-���B��N���N���B�i>.���������Ѽ�<���żS�o��(%�)�@���U��Ma�N�`� �S���=�(�!�����Rμdm��#i�G+.����ڻ@w���󶻋$���m̻�����	��;)�%LU�6ψ����9h�f\���-��M��/h��o{���*����q��L[��A��*��z��;�!��.���G�Y�c��b}�򱇽5������Yd��h���J�տ,��H#�
�μ<|��9������R���TΒ����)���.��:v������ؼ�������-��iK��ak�[焽.x��	�������}���ޏ����	o���Y�IM�TL�3�V��Gk���騐��!��6!���H��d\��u<������hp��R�ǜ6����k3�<d�B"���a�޼�ۼ=�ۼ�u޼i�伧��@5 �Љ������3���N��/m�=���/������ä�����0���s퓽Mچ��s�I�_�]iU��V�Z-d�az�ԋ���}��Pt��}r���s��"������8���F�j�tPM�2�3�����1�k ��v��kV𼣓�%$�q�|��������0h��w��|-�ߢE��)b���������;������!����k�����d��tՇ�Xw�}0f���_�@xe�-v�vD���Ԕ����ߜ���  �  ��������"�]�� ������V���Z;pH�;�B<i�9<��M<]fY<X_<�a<��`<"E^<,FY<tP<"�@<�1(<ei<��;�V�:�{K��^����H�p���������������:Mu���8����5a����!�ۺaGL��Qƻ�("��c��B���坼f^���'����v���3���һ����K;���;$d�;�@<�+<%�5<{;<��<<"�<<�y:<575<� +<��<a��;�b�;h\;=���ϻ[(4���y�*ܗ� Ŧ��V��̙��7��1�E�c�ξ���ړ�q���Y�񻈟4��{��A��Q[���ʼ<�ɼ<]���-��=����7�����g�LP��4�:&?;�3=;�MH;��@;��-;�/;~�:�n:�l;�A��b���e��,-�fNu�^���ȼ��Y���6����G*��C�߼���9]��蓼�������خ���μ[F�1	�c��=>��e�ķ�������ؼ\���,��~.r�#�I���.���(z��r�'k���m&�x0��>�D�R��No�`���N���RdƼ�켢�	�����,�K7���:�)
7�v-�X%��n��������N����4���!�(2��c@��!I�2�J���D��8���'�W,�m��I����ɼ՞��;���񨞼Ll��t���k���i�������-U���_��U��-����4ȼɏ�ɖ����'��i8�ĶE���L���L���E���8���(�9Z��1������v����I.�X�=��J��/P���N�f�F���8�o '��p�?������μ�#���x��Pf����������줼���z����~�����!����̼��⼖���17��C$�%7���G��.S��1X��U��L���>�`�.�%��������	^����͍.�+?�P7N��X��  �  iB����x�\�P��M�.Ȟ�r���%�f;�[�;�<p�8<�UL<��W<�]<j�_<�_<�]<��W<��N<�?<0&'<#N<�ȩ;���:�23����}�=�٨w��G���,��#ʉ�Hh�~�-�G�޻��j��Ѻ!3��6V.�Ľ����XUW�mX��j���w혼%��7sj�2�)�1Ļ.�ٺX�;N��;;��;v�<>C*<�r4<��9<��;<��;<,19<q�3<ϑ)<�y<v�;>
�;J�;��ͺ&»O�*���m�m�]_����;֒��v��P;��'�����D���8��U⻸`+��p�Pߙ� F��I�¼��¼ߞ���l���v�\�1�Il�3@a�M<P�#9�:�Z;��6;��B;�;;6&);��;���:��V:�獹m�}J����޻�\*�2p�����ü�c�x ��;y�����e���ټ���9$���F��M,���q��F���w�ɼjs켣�����������^}	�-�����ԼS9�������'q�!J���/��, �|��5��q�����l�'�K�1���?�T��Lp�g������ļ����R1���)�K�3��7�q3���)�bO�
����S�����;��oR��r��	/���<��mE��F�DA��l5��Z%��Z�)��fp�g�ɼK����L���n��`*���b���;���<��X_��Y��]&����������S	ȼ���$� �PT���$�"g5�>?B�o7I��'I�m%B�c�5��A&���'K��=��?��%��Y��;+���:���F�	uL��NK��IC��5�;�$�D��d�����s�μ�����1���,���]�����W|���V���g��(A���Ѳ��@����̼�T��P�����zL"���4��`D��O�9uT�%R�a6I���;�H ,����$��^������B,��><��J��U��  �  �r\��[P��,�~�ﻧ�e����9=ρ;�^�;Ou<�%4<��F<u�R<DY<��[<�[<��X<1 S<�$I<J�9<��"<��<z�;bv;-�B���N����R�j�s��C|��k��_C��|�(樻����
Ĺ�G��P���xۂ����Y�4���e��������C0s�ȁH����\k��R|w�D�#;S��;*E�;#�<��$<3J/<c=5<D�7<�7<��4<�.<�$<I<���;��;�M&;��l��A���h�J�L�RX{�*���w���G~���R�:.�,�ѻ����>?�Lb�絻�'��JQ�PƇ�5>��紭�J��Iޡ������^��� �S�ͻf�T���f���Q:v�:�� ;R�.;ڿ*;��;�*�:�2�:�2:N��U�	�"�����ܻ]�#���b��n���4����Ҽ��7����9���ȼgF�� (���������D������|�����ۼ����<�������ȉ ����
�ɼ�"�� �� �o�ՊL��d4���%�J�zp�����#���+���6�;DE��GY��qt��O������5��H�����h�B9 �_)�ҁ,�GD)��� ��B��?������<�켕�����}��&M&�3���:��{<�Zy7���,�r��U��EE��D��ɼ�����Ҫ�7.������-���]1��:.������󛜼h桼M���ɶ�0Eȼ#J߼Y���T����]-�D�8�{�>�Ұ>�}B8���,�������L��eY �tJ����2��b]#�z�1��s<�*�A��A�V�9�N�-����X��C���X��Fϼի��cܴ��筼 ֩��ק�"i��#X��h����䮼8���@����"μ������,��]��Z-�`�;�v�E���I���G�$�?��3���$���2���9�0v�ڭ�	%���3��hA���J��  �  ����f��&�����lG�:};�;���;�m<�!)<�;<!�G<ÏO<ƠS<$�S<)pP<-.I<��=<��-<FG<g+�;`��;�9(;/���X~������AL8��>�/�͆��|��I�0���L@�:���:_:0�����a� ���+���E�p(K��:������ӻc$W�03��P0;���;X��;�^<�#<��$<�<,<m�/<�/<��+<�K$<<��<WV�;n��;Sq.;O�:�/�\�o�ٻ�F	D���X���X���C�cz�	��۲����5n���2ں�+h��)Իn�"�9�Y�u�������UO������j�?=��'�亻�bT�B���*9qі:�B�:N\;�];� �::[lD: f �⪫��5��\��Mc���A�R�̏��_��V����%˼-ӼT}м��ü>ʯ���G���m�:f��"v�o����%��ePü��ܼ3��_���z�����e|Ӽ�b��C���`��2r�o�T�	i?�X1��,)� �%�k�&��V+��3��$@�A;P���d�r�~�r����գ��⻼V׼���z�����g~�O�9�F���B�[>����%ݼ�QݼW��.b�����KK���$�Y�+��9-��c)��� �2P�ZA�[����K߼ż˼�E������������������(����������ġ�S����������w�ʼ�<޼-���3���1��e!�L�*���/��L/���)���0_�)E�������>��/> ���
�̣�G$�k�-��2�2��m,�#�"��z�n	�����19��~Ҽo�ļ��������Ԯ�Y��-O��Ye���_��8K��zl��CAż�aҼfa�ځ����-��v#��/��87�ě:�r�8��k1�i�&�+�:����������w��x����'�1[3�j�;��  �  S���V7���$�����1���;B=�;fi�;��;!H<�w&<�5<��?<��E<��F<@B<,�8<L�*<�<��<�+�;�I�;((-;s��9�=������ƻ�r�:�\һ6$���z�`�Y94�;�l;?�y;R<;Ld|:��Ⱥ�'��M/ϻ̈�����w{��L!ʻ":����fY�9�';��;ٻ;��;><�<� <5u"<]s"<�<��<�<y�;c��;l^�;�4;�e$9�\�i����Kػݒ�����(���*����m��S�����9�s:
=�9�6����o�Ϋ׻��U3@��3W��+]�n�R��	<�J:���������w�Jh�%���0k�V�:���:�0�:���:�H:��P�7`��z0'�ޅ���$���/��G(!�T[H���q�I�]j��[ê�����g��i���%��_a�9A^�,�H���C�g+R�ӧq����{J����T̼�4Լ��Ӽ��˼pi���뭼hϜ��ό���}���f�{CT���E��;��5��D4��E8�i�A��SP��	c��Qy�yw��b��"���+ ���eϼZ伄9��tV�,�	��6���(��N+���C�etӼ3C˼w�˼j�ռ3:�GM����	����!��6��W����>��	��.�(�ἣ�Ҽ=�ż�������Ϊ�
���5ܢ��Ţ�_g��4v������(����}ż�^Ҽ?x� ����OG�I��-M��k�u����7)���M�����#��63�{��3g��n�	�d�C4�t� �!���M���j�/:�!���W�輱�ڼ_�μa5żlE���9���Q���籼;��o0���p��l�ż��ϼ֪ۼ���g���X����+K�x!�&'��	)���&�� ��������8��g��q���`���*��h6�����"���)��  �  �b��1�������R[(��p:g�	;�X;;V�;ٟ�;Oi�;=�<�4<�(<�51<Z3<*$-<1 <�
<I��;[�;���;>OT;
��:EJ:}�J����@:��(U��xG��@�o�,��I�:t�P;��;X��;�x�;i�;�Ls;V.�:�!�����\a��������
�`��a!�����\򑸁Ś:#�;s�s;��;S��;�q�;z�<�k<�<q�<���;`��;�ڢ;�Wn;�G;�:�����պs�<��[���h���ڣ��ȗ�<vm��a	�,�����:�*;�6H;{\*;���:AGK�MO����4�����������Ź��%���Z̻���}ш�GWN�~����4��G��O���)���Һi\?�2ב�[ ǻ�����N�n�1��J���b���y��3��~G��]���~ɉ�A���E�g�H�K�{�2��N#��� �p-��\G���j�����j֚����籼������}���ʥ��@��Ő��t򋼒f����u�!�e��bW�wM�[�H��K�ДV��rh��`�ϛ��B
��_\��a���*��-�ͼDڼp/����6�%n�^C��G�M5׼бɼj�����������P¼��м�T⼼���ea�<���
���/����� �����:�����jּ�˼�@������pذ��ܬ������m���f��!���X(˼Mּ��뼜���Z� �S��I
�u�������(L��l ���� "�nռ�ϼwDмu�ؼ�漋L������
��>����(����6������������߼�ռ�˼c�ü7���»�k����¼�˼Sռ}�)��s#��	'���F+�3B��g�x�����lD��������� �������7�^�"�󼰋�t*
��4��e��  �  1�;���:"��:#{:q�h:zԀ::#�:?��:Ӻ:;��;�˶;r�;Ra<�<��<��<s��;�]�;�}�;^xI;��:�y>:i@G8-"�����(�ы�Jz����:���:8-?;p��;i�;���;V <��<��;P��;ϕ�;UJ;>$�:l��9p�'��5���uϺ���6�ߺ~1ƺ���3��	�M:�;��s;ˏ�;�K�;��;;��;���;)P�;�v;��;�
7:�x��c��7���V�����r�#%�ٺ��v��%�8���:o0;
z;��;�i�;�M�;��b;&��:���'@�ϩx��"�� лJ�4\��������6	�ˉ��]��7�ǻVѠ�o�o��'�������x��Ee�n꨻��j���-� �C���S���^��Me�|i��Kj��'h�j�a���U��WE��E1����(v��Q�������� ��<���[�cz��q��:ᔼ1c��\���p���!��	}������w��1?������*z����|�B�l�6d��e�q~r��n��㒼���R���Ǥ��t�ȼX�ϼ��Լk�׼l�ټ�Uڼdټn{ռ�Nϼ��Ƽ輼qE��qͫ��A���ɩ�#����ʻ�D�ɼ��ؼ/<漬������<���#��������� ��������� i���⼯ ּ�ɼ�ٿ��G���
���2��O�ȼpռ�#��!�r���_������2��U3�r����e �6m�����y�6�׼q/̼<Kü�徼�뿼T=Ƽ��м��ݼ���T���x; �������5��n`��.��.�l��� �������m�߼)oԼ?[̼~�ȼf˼YUҼ<ݼ��a������N�	���&��S1�������,�	�k���� �A��;����޼��׼a9ռaFؼ�U༘�.m���M�&	��  �  w�;jjl;τ;bHr:�}��$㣺Z:�7�ۺ�zn���9��;T�;���;f<�;(m�;��;�ٮ;
�^;<<�:B�D���z5�R;�=/�����i����Z:"�;tW;�E�;Fq�;��;��<�;<x�<qX<�b<;�<�X�;���;	�;R�L;��:�$�9ԙd��a��U��Ą�@��<�����A�ύ��$Q :�(;�W�;7�;��;( �;�C/;�.6:�߭�P8G��i��H�����O|��m:��ݺ���`X2:�M�:��C;_��;�-�;���;���;�h�;��;���;˂;:� ;�O:Kj���&�Vg��(@�����/�H�#� �1���6���0�� ��a�}�ػ ����肻�2s�����R㽻��\�'�kM��$k���~��w��	R��bxz��k��Z�O/I�P�7���&�I��S��Pe��ջ��ʻ[�ͻ���0 �\:�0��0K�ɯe���e��˘�	Ԥ��篼"޸��D��Rݾ�����Q��!+���1���l��{�������6��,��z_��ڽ���ϼ�ݼZ"強��8'�Rh߼\�׼4�ϼ�jǼ�D��I-��#��u��ՠ�1-���q���T�������)���*����μ4+ڼ���A�\���r���y<�F[�J�
�ʇ�5���Ar６:߼�Ҽ�ʼ6ʼ� Ѽ,�ݼ�����[�$���Kg��	��o��� ��������t��	ؼ�ͼs�ü�������������q�����"پ�Ʊȼ�Ӽ[�޼��.&��O �M����
� �����
2����� ����+�����,�ݼvټ��ۼ#6������:�
��H��Q�Փ��P��'����s	����<��j/��� �u�߼�ּ�μ�ɼ�	ȼeʼ?]м�ټG����aA���  �  o�;���;��;d��i(��@��鱶��"��'7��_pi�Ƨ����: _;JǞ;�5�;Eϑ;Z�.;�Ee9��ۚ���λ���/ֻ�v����]� ����~�:�~L;F�;�i�;�. <��<� <d<*<�/<�0<��*<�� <��<� <i��;��;#�N;P��:�B����i��ͻ����h��u�B�뻒s���B8�1���{�:��<;��?;w0�:�'��/��J��r��p�������ӻ-L���[�;�+6�~ ;A�m;���;���;�;!��;O>�;^��;O�;���;��;֌;uK7;=8�:�_�Z!G�ꮲ��E���,�G�Q�l�l��nz��w��#e��SF��!��7���cϻ�����sֻ;5��&2�a�a��5���q�����C���K��3�����~�Cs\���;��%��3�e���ɻ#d�����頻RϦ�ͷ��ӻ�����g�)��$F��7f�#-��"���"���N}���CҼu�ݼ)y�G6ݼ]}Ѽ���~=���k��k┼K��s؜�-׭�5ļ��ۼ��� ��y�ӷ�������m޼��ͼ�����n������};������\��y��\���B��������Ȧ�#;���;����ʼ��ڼ�켠#���>	������Ϧ��V�i��������$�����iܼ��ۼ��h�� ���,�`��w��%��E���0����D~�������ӼibǼ���谴��$��ǰ������d���ʫ����U����¼vμ��ۼ�뼴����g���j��z ��#��!�p��[�"0	�������)���������B����#�z�"�g�&��p&��["�6_�'��Z�	��� �(����5ټh�ϼt>ȼ!�¼� ��*6���	��brļ�˼�Ӽ+޼�Y��  �  �w�;7�;�L�:���K֥�R���VE��I'��������<���4�麚�i:�-;��L;x\;SWg8|�=��sƻ~i��K.�E�7��/+�w���|����/���9?Z;M�;���;�-<�[&<_82<��9<Ze=<5N=<r9<0�1<�#&<�<�K�;��;po;�;a:���������z5�L�]�N�w";��x���ɻ9�M�l.�ͪC:+�R:y)���?�`mû{��g�;��WR���S���?�q�LNֻ��\�z���L�;��;���;�;`�<��<�<u�<�<UN�;&��;9`�;��;�i;�K��h�5�û�T�.BS�V���8���6�����<��������U�tT+�7��w�}����0��b��-��Ӈ���]���bż�Sļ���i٥�"'��F�j��F<���2�뻏p��՟��g��@턻l愻.����K���J����ѻ����O���4��7[��ۄ��h��(����׼K��p���p��7 �L��ݼj�Ƽr�����q-��K��4ü�|ݼ����-	���l��@�����J�����fҼ����˪��1��I����Z��}ۉ����]!��q{��ߏ��qR��_���8���d����¼O\ּ���x��K{�<�c�'��-�&.��()�����s�������x��S�F�����O����U�(��s.���.���)�8� ��x�+T��-��̗޼��˼�o�������ͪ�����HS���	��`���j-��៨��9��Sq����ļCռ�h��� ���_��S{'��H0��~4�BS3���,��"�$-��p
��������T���d�H��:��Y+�OL4�
n8�7�+�0�ύ&���� �7� ���켬�ۼ��μ�cżƽ��k����t���o���k������?LɼުӼGn��  �  �C�;貇;���9�}o�y���f�2���W���d�X�9�3�����UR�������PQ:z�:�j�9���������I�ek���t��yd�e=��)��̍�QJ���G;|4�;�4<Et <�2<��<<W�B<;tE<IE<�B<�;<Å1<�M!<�M	<YO�;�Rl;48y9�m��|��8�:�Ƿk�RB��,)���rv�N<K�?u�����Z�/�����:��V#�����_��H�c�v�������Lw�J\I�,Q�7w��o脺�I;L��;��;}�<�<R�<cR<�G<�<H�<R�;���;�!�;ܺ5;�\[9^E�K3߻)4��y�pl�������۾��N��e~��Qj��{���EP�խ,�Փ���,��R��O��1��\ü]ټ�%�O��o+Ӽ���}����|}�`D����	ݻi����N���An��c��h���z�����o��O�����
���,��yY��N���I��j�ʼ9��6&�0������[������;iۼ$Jļ�ڵ�d��������Լ���d	��`�>� ��"$�Z� �����
�������ټ�⾼/���&���U֍��c��t^���΃����r������*�����ϧ��ݭ�[����ּ&��>L	����'H)�=}5�أ<�օ=���7�-�v��� 
�`���������)v�ٷ�;,��7���=�b�=���7��,��9�O�^����g߼3ɼ̃���Ƭ� ���f���𝼃��-������/W��Lh��5����L����Ҽ�3�H:����$�ۖ3��n>���C���B�{];��`/��)!�f���	��1�cP�'���q�E+��&9�ZVC���G��E�Y�=��81���!�D����=K켵:ؼ	�ɼ�����*�������峼������������6��klü�5μ��ݼ�  �  ���;�6q;�������=��.W��"��{}��{���xY�x� �(�Ļg-.�Ճ�e�19�s}���m�S��k�7��p��l��dk�����W`�0r"�$��w����B/;���;� 	<�U%<��7<u1B<?�G<�pI<��H<�ZF<�@<��6<ə&<7J<��;�<^;�м�瘻E1�J�Z�)Έ��꘼�*��TD���co�y�2��c�0 ���W�yH��nz���߻�.��Jl�@*��~����ڜ��Î��Tj�6(�����vںh3;�à;�N�;~�<fc<	�<u<,�<��<�"<� �;���;I��;K�A;��A9�u[�]���OH��]��棬��_Ƽ��ӼS3Ӽ
ż_����̏��	i���A�O	3��@��i��蒼P����ռЫ�L%���"��L���jʼ1���u���ML�!��:&ٻ2%����z�o�X���O��$X���k�y�����������׻���*��Y[� ��S���E�ռ�����6�	��b�\�����q:�|J���ϼ�����:���ȼ��༩� ������ �R$+�o�.��*�X� ���T��B����tC��5���S��Ꮔ�5���!o���䂼`o��t爼
����E��M��Ы�y��zXؼǐ�����g �;N1���>�-�F�^H�w�A�c6�M�&�!K�`�
�D�!��Y�	�����^%�}�4��nA��UH�6?H�h*A��M4�s�#����\ �yzἣ�ȼȣ��+���P��Q����Û��+��I����c��7���ܦ��6;������ӼA��E��p�s�+�)<�-CH��8N��M��E��8�M�(�:�����
��V�IV�AB#�Z3�`pB�+�M��_R�0P�(G���8��'�t�����Pv��F׼ZǼ�μ��v���#���ұ��Ա�=鲼D������ӱ���˼�gܼ�  �  �q�;r�d;��]����� %��:d��^���������f��H,���ػ7O��f��b��X��n���ݜ�8�C���}��Ñ��▼w8����l���,�ӄƻG$̺j�$;�;�;��	<3�&<9<M�C< �H<��J<�J<S�G<OPB<9�8<p(<�7<�T�;�?W;w��糧~c�5�f�;���EI������Z���#|���=�����1����!0���*�ʌ��U�f�8�t�x��0���m��!D��R���VGv�T�1���λ����S�:'�;~��;�@
<��<v�<+�<:�<k�<�^	<3��;n��;�?�;�8D;�9t`e�ս �ƌO�Wk��ݲ��rͼ�Vۼ'�ڼ�˼޲�(����q�EI���9�`�G�9�q�볗�U���=ܼ����YM ��g��b"�r�ϼX|��j��S�O��K�P�ػ[���w�t���R�|JJ��ZS��Bg����Tl�������%Ի+��y*�ك\�A���rz����ټ�( ��z���p  �=������/Լ�üƝ��}̼_7弤&�=���V$��.��J2�|V.�C�#�6�����6�⼍2ü;���ꖼ�����ă��ြ���nH��:؄��@���ی�)y���5��vU������3ټ~����1�a"��74�#YB�}�J���K���E��N9�C�)�ޙ�σ�e �t���z�J%�t(��8�F�D��L���K���D��H7��&��E�.!�.v���ȼ8��x��͉��4%��!��
������p�������᥼�����]��cӼ�#�zv�cK�#O.�PB?�$�K�o�Q���P��H�D;�b!+�E �������n��Z�F�%�36�J�E��Q��V���S�cJ���;��)��6����} 0׼��ƼN��\���Jp���7��dE��xP��q���5ĸ���Y˼�@ܼ�  �  ���;�6q;�������=��.W��"��{}��{���xY�x� �(�Ļg-.�Ճ�e�19�s}���m�S��k�7��p��l��dk�����W`�0r"�$��w����B/;���;� 	<�U%<��7<u1B<?�G<�pI<��H<�ZF<�@<��6<ə&<7J<��;�<^;�м�瘻E1�J�Z�)Έ��꘼�*��TD���co�y�2��c�0 ���W�zH��nz���߻�.��Jl�@*��~����ڜ��Î��Tj�6(�����vںi3;�à;�N�;��<kc<�<
u<7�<��<�"<� �;��;~��;��A;��A9:u[����*H�u]��ԣ���_Ƽ��ӼD3Ӽ
żT����̏��	i���A�M	3��@��i��蒼%P����ռޫ�\%���"��^���jʼ.1���u��NL�A��u&ٻd%��P�z���X���O��$X�ƨk�q�����������׻���*�uY[����A���3�ռ�����6� �xb�T�����k:�tJ���ϼ�����:���ȼ��༬� ������ �Y$+�w�.��*�a� ���^�C�,����C��5���S��폄�?���*o���䂼eo��y爼����E��O��Ы�y��zXؼƐ�����g �;N1���>�-�F�^H�w�A�c6�M�&�!K�`�
�D�!��Y�	�����^%�}�4��nA��UH�6?H�h*A��M4�s�#����\ �yzἣ�ȼȣ��+���P��Q����Û��+��I����c��7���ܦ��6;������ӼA��E��p�s�+�)<�-CH��8N��M��E��8�M�(�:�����
��V�IV�AB#�Z3�`pB�+�M��_R�0P�(G���8��'�t�����Pv��F׼ZǼ�μ��v���#���ұ��Ա�=鲼D������ӱ���˼�gܼ�  �  �C�;貇;���9�}o�y���f�2���W���d�X�9�3�����UR�������PQ:z�:�j�9���������I�ek���t��yd�e=��)��̍�QJ���G;|4�;�4<Et <�2<��<<W�B<;tE<IE<�B<�;<Å1<�M!<�M	<YO�;�Rl;38y9�m��|��8�:�Ƿk�RB��,)���rv�N<K�?u�����[�/�����:��V#�����_��H�d�v�������Lw�J\I�,Q�8w��q脺�I;P��;��;��<�<^�<sR<�G<�<h�<��;��;7"�;��5;Ll[9SE��2߻�(4��y�Ml��c����۾�dN��L~��<j��j��yEP�ǭ,�ғ���,���R��O��1��sü7]ټ�%�p�ἒ+Ӽ �������|}��D�ϯ�zݻ����PO�� Bn��c��h���z�����o������ỵ�
�V�,�yyY��N���I��F�ʼ��%&������r[������,iۼJļ�ڵ�c��������Լ���d	��`�L� ��"$�k� ����!�
�#�����ټ�⾼P���D���p֍��c���^���΃�"���%r�����+�����ҧ��ݭ�\����ּ&��>L	����'H)�=}5�ף<�օ=���7�-�v��� 
�`���������)v�ٷ�;,��7���=�b�=���7��,��9�O�^����g߼3ɼ̃���Ƭ� ���f���𝼃��-������/W��Lh��5����L����Ҽ�3�H:����$�ۖ3��n>���C���B�{];��`/��)!�f���	��1�cP�'���q�E+��&9�ZVC���G��E�Y�=��81���!�D����=K켵:ؼ	�ɼ�����*�������峼������������6��klü�5μ��ݼ�  �  �w�;7�;�L�:���K֥�R���VE��I'��������<���4�麚�i:�-;��L;x\;SWg8|�=��sƻ~i��K.�E�7��/+�w���|����/���9?Z;M�;���;�-<�[&<_82<��9<Ze=<5N=<r9<0�1<�#&<�<�K�;��;po;�;a:���������z5�L�]�N�w";��x���ɻ9�M�l.�˪C:*�R:{)���?�`mû|��g�;��WR���S���?�q�MNֻ��\�����O�;��;���;)�;l�<��<�<��<�<�N�;���;�`�;$�;�j;P����5�KûWT��AS�%���8���6��އ���������k�U�ST+�$��w����ԍ0�b��-��􇧼�]���bż�Sļ����٥�U'����j��F<�r��Ү�q���՟�Oh��~턻�愻4����K���J����ѻ$����N�@�4�T7[��ۄ��h�������׼��A����o��7 ��K���ݼT�Ƽc�����q-��R��Cü}ݼ���.-	�������X��7��K���	gҼ˭��/˪��1��n��� [���ۉ����q!���{��돏�yR��e���<���f����¼O\ּ���w��K{�<�c�'��-�&.��()�����s�������x��S�F�����O����U�(��s.���.���)�8� ��x�+T��-��̗޼��˼�o�������ͪ�����HS���	��`���j-��៨��9��Sq����ļCռ�h��� ���_��S{'��H0��~4�BS3���,��"�$-��p
��������T���d�H��:��Y+�OL4�
n8�7�+�0�ύ&���� �7� ���켬�ۼ��μ�cżƽ��k����t���o���k������?LɼުӼGn��  �  o�;���;��;d��i(��@��鱶��"��'7��_pi�Ƨ����: _;JǞ;�5�;Eϑ;Z�.;�Ee9��ۚ���λ���/ֻ�v����]� ����~�:�~L;F�;�i�;�. <��<� <d<*<�/<�0<��*<�� <��<� <i��;��;#�N;P��:�B����i��ͻ����h��u�B�뻒s���B8�3���{�:��<;��?;v0�:�'��/��J��s��q�������ӻ.L���[�ʇ+6�~ ;M�m;��;���;7�;L��;�>�;���;��;0��;+�;�֌;�L7;V;�:M�_��G�����E�Q�,�͛Q���l�Knz���w�,#e�RSF���!�B7���cϻ�����sֻY5�'2���a��5���q�����|���K��q���Y�~��s\�S�;�8&�a4���|�ɻ�d��Q���A頻YϦ��̷�\ӻ��������)�J$F�E7f��,������䢭�}���CҼ<�ݼ�x�6ݼ3}Ѽ���c=���k��b┼J��|؜�?׭�25ļ��ۼ�� �z���ǫ������m޼��ͼ4����n��Ѻ���;��۶��~��;y��t���B��������Ȧ�(;���;����ʼ��ڼ�켟#���>	������Ϧ��V�i��������$�����iܼ��ۼ��h�� ���,�`��w��%��E���0����D~�������ӼibǼ���谴��$��ǰ������d���ʫ����U����¼vμ��ۼ�뼴����g���j��z ��#��!�p��[�"0	�������)���������B����#�z�"�g�&��p&��["�6_�'��Z�	��� �(����5ټh�ϼt>ȼ!�¼� ��*6���	��brļ�˼�Ӽ+޼�Y��  �  w�;jjl;τ;bHr:�}��$㣺Z:�7�ۺ�zn���9��;T�;���;f<�;(m�;��;�ٮ;
�^;<<�:B�D���z5�R;�=/�����i����Z:"�;tW;�E�;Fq�;��;��<�;<x�<qX<�b<;�<�X�;���;	�;R�L;��:�$�9ԙd��a��U��Ą�@��<�����A�Ѝ��$Q :�(;�W�;7�;��;( �;�C/;�.6:�߭�R8G��i��H�����R|��m:��ݺ���wX2:�M�:��C;v��;�-�;��;̇�;i�;���;=��;�˂;�� ;0�O:Dj���&�Sf��?������.��#�~�1��6���0��� ��a���ػ�����肻�2s������㽻����'��M�]%k��~�x��LR���xz���k���Z��/I���7��&��������e�m�ջ'�ʻd�ͻk�� �&:�y�0�>0K�a�e�����d���ʘ��Ӥ��篼�ݸ�|D��ݾ�J��vQ���*���1���l��q�������6��",���_��@ڽ��ϼݼ�"����|'弘h߼��׼y�ϼ
kǼ�D���-��I#���u��)ՠ�R-���q���T�������2���0����μ5+ڼ���A�\���r���x<�E[�J�
�ʇ�5���Ar５:߼�Ҽ�ʼ6ʼ� Ѽ,�ݼ�����[�$���Kg��	��o��� ��������t��	ؼ�ͼs�ü�������������q�����"پ�Ʊȼ�Ӽ[�޼��.&��O �M����
� �����
2����� ����+�����,�ݼvټ��ۼ#6������:�
��H��Q�Փ��P��'����s	����<��j/��� �u�߼�ּ�μ�ɼ�	ȼeʼ?]м�ټG����aA���  �  1�;���:"��:#{:q�h:zԀ::#�:?��:Ӻ:;��;�˶;r�;Ra<�<��<��<s��;�]�;�}�;^xI;��:�y>:i@G8-"�����(�ы�Jz����:���:8-?;p��;i�;���;V <��<��;P��;ϕ�;UJ;>$�:l��9p�'��5���uϺ���7�ߺ~1ƺ���3���M:�;��s;ʏ�;�K�;��;:��;���;(P�;�v;��;�
7:�x��h��<���Y�����r�"%�ٺ��v��)�8��:�0;mz;��;j�;N�;��b;���:�臸�>��x��!���л3�[�����/����Ј��z��p�ǻ�Р�j�o�]�'�A���u��Sx�)Fe��꨻F�zj�U�-���C�Q�S��^�INe�i�GLj�w(h��a�@�U�XE�@F1�յ�Vv��Q������b� ���<���[��bz��q�������b��:\���p���!���|��}���w���>��Ğ��z��m�|��l�!d��e��~r��n��$㒼F�������������ȼ��ϼ��Լ��׼��ټVڼ�ټ�{ռ'Oϼ��Ƽ@輼�E���ͫ�B���ɩ�4����ʻ�L�ɼ��ؼ2<漮������<���#��������� ��������� i���⼯ ּ�ɼ�ٿ��G���
���2��O�ȼpռ�#��!�r���_������2��U3�r����e �6m�����y�6�׼q/̼<Kü�徼�뿼T=Ƽ��м��ݼ���T���x; �������5��n`��.��.�l��� �������m�߼)oԼ?[̼~�ȼf˼YUҼ<ݼ��a������N�	���&��S1�������,�	�k���� �A��;����޼��׼a9ռaFؼ�U༘�.m���M�&	��  �  �b��1�������R[(��p:g�	;�X;;V�;ٟ�;Oi�;=�<�4<�(<�51<Z3<*$-<1 <�
<I��;[�;���;>OT;
��:EJ:}�J����@:��(U��xG��@�o�,��I�:t�P;��;X��;�x�;i�;�Ls;V.�:�!�����\a��������
�`��a!�����^򑸀Ś:#�;s�s;��;S��;�q�;z�<�k<�<p�<���;`��;�ڢ;�Wn;�G;�:ȑ���պu�<��[���h���ڣ��ȗ�vm��a	�	�����:*;n7H;M]*;���:{BK��KO�L���3��@������;��[%���Y̻'����Ј��UN��|����n���������)���Һ;]?��ב�
!ǻ���� O��1���J�e�b�?�y��3���G�������ɉ�q�����g���K���2��N#��� �p-��\G�\�j�f���=֚�����籼�������}��?ʥ�W@������9�\f����u�ԗe�hbW�OM�F�H��K��V��rh��`�����p
���\���a��+��p�ͼ�ڼ�/��7�dn�C�H�{5׼��ɼ������������P¼��мU�����ga�=���
���/����� �����:�����jּ�˼�@������pذ��ܬ������m���f��!���X(˼Mּ��뼛���Z� �S��I
�u�������(L��l ���� "�nռ�ϼwDмu�ؼ�漋L������
��>����(����6������������߼�ռ�˼c�ü7���»�k����¼�˼Sռ}�)��s#��	'���F+�3B��g�x�����lD��������� �������7�^�"�󼰋�t*
��4��e��  �  S���V7���$�����1���;B=�;fi�;��;!H<�w&<�5<��?<��E<��F<@B<,�8<L�*<�<��<�+�;�I�;((-;s��9�=������ƻ�r�:�\һ6$���z�`�Y94�;�l;?�y;R<;Ld|:��Ⱥ�'��M/ϻ̈�����w{��M!ʻ":����eY�9�';��;ٻ;��;><�<� <5u"<]s"<�<��<�<y�;b��;k^�;�4;�e$9�\�j����Kػݒ������������m�S��K��9M�s:�B�9�4��~�o�.�׻����2@�G3W�+]���R�p	<��9����� ��,�w��f�z���dY���:Ф�:L1�:���:�G:T�P��a��v1'�z����%���0���(!��[H���q��􌼚j���ê��������Fi���%���a�aA^�C�H���C�Y+R���q�쁎�ZJ��� ��%̼X4Լ��Ӽ��˼2i��r뭼+Ϝ�Rό�R�}���f�(CT�r�E�Ҭ;���5��D4��E8�y�A��SP�
c��Qy��w�����W���e ��fϼ]Z��9���V�J�	��6���?��w+���C⼃tӼKC˼��˼y�ռ?:�OM����	����"��7��W����=��	��.�'�ἣ�Ҽ<�ż�������Ϊ�
���5ܢ��Ţ�^g��4v������(����}ż�^Ҽ?x� ����OG�I��-M��k�u����7)���M�����#��63�{��3g��n�	�d�C4�t� �!���M���j�/:�!���W�輱�ڼ_�μa5żlE���9���Q���籼;��o0���p��l�ż��ϼ֪ۼ���g���X����+K�x!�&'��	)���&�� ��������8��g��q���`���*��h6�����"���)��  �  ����f��&�����lG�:};�;���;�m<�!)<�;<!�G<ÏO<ƠS<$�S<)pP<-.I<��=<��-<FG<g+�;`��;�9(;/���X~������AL8��>�/�͆��|��I�0���L@�:���:_:0�����a� ���+���E�p(K��:������ӻc$W�03��P0;���;X��;�^<�#<��$<�<,<m�/<�/<��+<�K$<<��<WV�;n��;Qq.;h�:�0�\�p�ٻ�E	D���X���X���C�Zz��໷������<m���1ں�*h�_)Ի,�"���Y�L�������%O��p����j�?=�2'�Q㺻�aT����*9?Ӗ:D�:�\;,^;� �:���:�jD:�o �y����5�%]���c�p����R�����M_������&˼�-Ӽ|}м��ü[ʯ���G���m�=f��"v�b���z%��JPü��ܼ�2��_��wz��̤�3|Ӽ�b�����1���r�!�T��h?��W1�f,)���%�\�&��V+�+�3��$@�j;P���d���~������գ��⻼�׼3�󼔌���~�f�%9�Y���B�x>�����3%ݼ�Qݼd��7b�����MK���$�Z�+��9-��c)��� �2P�ZA�[����K߼ż˼�E������������������(����������ġ�S����������w�ʼ�<޼-���3���1��e!�L�*���/��L/���)���0_�)E�������>��/> ���
�̣�G$�k�-��2�2��m,�#�"��z�n	�����19��~Ҽo�ļ��������Ԯ�Y��-O��Ye���_��8K��zl��CAż�aҼfa�ځ����-��v#��/��87�ě:�r�8��k1�i�&�+�:����������w��x����'�1[3�j�;��  �  �r\��[P��,�~�ﻧ�e����9=ρ;�^�;Ou<�%4<��F<u�R<DY<��[<�[<��X<1 S<�$I<J�9<��"<��<z�;bv;-�B���N����R�j�s��C|��k��_C��|�(樻����
Ĺ�G��P���xۂ����Y�4���e��������C0s�ȁH����\k��R|w�D�#;S��;*E�;"�<��$<3J/<c=5<D�7<�7<��4<�.<�$<I<���;��;�M&;�l��A���h�J�L�QX{�)���v���G~���R�1.��ѻ����P>?��b��浻�'��JQ�6Ƈ�>��Ǵ��(��&ޡ�}����^�_� ���ͻm�T�v�f���Q:cw�:� ;��.;�*;��;�*�:S2�:81:����	�������ܻ��#�Ȝb��n���4��߸Ҽ��W���(9���ȼwF��,(����������D������m���q�ۼ����/��������� ������ɼ�"�����ío���L��d4�h�%��I�ep������#���+���6�XDE��GY��qt��O��-����5��k�����h�T9 �_)��,�VD)��� ��B��?������<�*켞��������'M&�3���:��{<�Zy7���,�r��U��EE��D��ɼ�����Ҫ�7.������-���]1��:.������󛜼h桼M���ɶ�0Eȼ#J߼Y���T����]-�D�8�{�>�Ұ>�}B8���,�������L��eY �tJ����2��b]#�z�1��s<�*�A��A�V�9�N�-����X��C���X��Fϼի��cܴ��筼 ֩��ק�"i��#X��h����䮼8���@����"μ������,��]��Z-�`�;�v�E���I���G�$�?��3���$���2���9�0v�ڭ�	%���3��hA���J��  �  iB����x�\�P��M�.Ȟ�r���%�f;�[�;�<p�8<�UL<��W<�]<j�_<�_<�]<��W<��N<�?<0&'<#N<�ȩ;���:�23����}�=�٨w��G���,��#ʉ�Hh�~�-�G�޻��j��Ѻ!3��6V.�Ľ����XUW�mX��j���w혼%��7sj�2�)�1Ļ.�ٺX�;N��;;��;v�<>C*<�r4<��9<��;<��;<,19<p�3<ϑ)<�y<v�;>
�;J�;��ͺ&»O�*���m�m�\_����:֒��v��P;��'����{D��{8��2⻣`+���p�Cߙ�F��9�¼��¼̞��}l��Z�v�8�1�l໲?a�}:P��9�:A[;��6;��B;.�;;<&);�;Q��:ԷV:ꍹ�m�J����޻�\*�Vp���
�ü�c伉 ��Cy�����e���ټ���?$���F��M,���q��A���o�ɼ`s켝�����������U}	������ԼA9�������'q�J���/��, �m��+��l�����q�'�U�1���?�*T��Lp�u������ļ��&��[1���)�T�3��7�q3��)�hO�
����S�����=��qR��r��	/���<��mE��F�DA��l5��Z%��Z�)��fp�g�ɼK����L���n��`*���b���;���<��X_��Y��]&����������S	ȼ���$� �PT���$�"g5�>?B�o7I��'I�m%B�c�5��A&���'K��=��?��%��Y��;+���:���F�	uL��NK��IC��5�;�$�D��d�����s�μ�����1���,���]�����W|���V���g��(A���Ѳ��@����̼�T��P�����zL"���4��`D��O�9uT�%R�a6I���;�H ,����$��^������B,��><��J��U��  �  &`Z;Ҵz;;��;���;[#<q\M<;fs<�3�<�}�<���<.��<��<�Q�<1��<�l�<���<�؞<?�<��<f�<.%�<�x{<�bX<��.<�.<�;�N;qd�:��:��;�Aj;rB�;x�<�!<��4<e�7<��)<~^<,�;Y��;�;��P:�:+��:E
S;ݞ�;�<+�/<�9T<�q<w��<2�<�]�<���<4 �<��<���<�^�<��<�<6��<4�<�m<J�P<��+<�� <���;�A-;&;1:a��`��[�9g;V��;�d�;)��;d�<'��;���;wr�;e9�:�R����\�Π��B���rs��� ��`�9� 0;:��;ҍ�;�k<7�<T�<L<��<�<g�
<r�<��;`W�;'V�;���;"J�;��B;�#P:���������77$��wB��Q��wO�d�=�5� �`^���»���.���w�����\��b.G�B�n�޴�������}��~��F]��`6�3��8׻���`yp�-�D�545�;�9��I��1_��v�^��������Y��ͭ����ػ���!�4}G��1t����:���Ee��Z�ɼ��μ�g˼���&t���4��1ܓ������>��v3���"���P��ϼ�e༏�IQ��漺�ؼ:�żOV���|���&��:u���`���S���L�>�I���H���H��*I���I�p�J�>,N�F"U�e�a��sv�ʸ��=+��oe���sǼM�ۼZv뼶���I���
+ݼֹʼ裸�򨪼'����������ʜ����Ѽ�传<�ف��=7�����z߼;V˼���e���3���i����w�f�m��Fi��h�wh��di���j��%l�"�n���s��2}�T��������ע����~�̼���vK��$��.�1��Js���4�)�ڼ7�ɼ ����!Z��·ʼi7ܼ��� �<,��  �  �d};)K�;5J�;zN <CK(<|�P<Xtu<䫉<B��<㓛<Z`�< �<^)�<-ؠ<`O�<z��<1��<�
�<��<L�<�K�<��|<z�Z<E�2<`u<E��;�An;ф;l��:kS%;�@�;zE�;�<G{&<�8<k�;<;.<-a<�2�;庐;m)#;$��:#��:�K;�-p;���;u{
<��2<��U<B�q<ϸ�<��<�&�<ހ�<�ڍ<,ύ<��<n:�<B�<@׊<�\�<��<:n<["R<Ud.<�1<nz�;��I;۾�:�8��V:��;�ґ;k��;,( <+�	<�O<y�;���;4��:�M^�	�;�HE��놻��S���ʺ�!:u�?;��;1�;��<@�<�o<��<k<�l<$�
<-�<	M�;���;D��;�k�;���;��E;0*o:vhҺ�!��dv�l���:���H�=�F���5������/��fΓ��f���K��t޻���v@��!g�#z��o����E���av���V�gu1�Ո��!ӻ�'��;�o�,�E���6�;;�� K��`��mw�I��bQ������f���ٻ[c����GE�fp��L��˙���p���Fż,Yʼ�3Ǽ��.���x�����������B��e�������J���y˼d[ܼ���@��
��ռ��¼)������R��J�t�-�`�e�S��-M�j6J�	EI�'I��fI�m J��[K�h�N��U��b�#�u�"���vŚ�vC����ļ.ؼ�`缢�＀��)���ټ~�Ǽ����}����������[������μ	
Ἑ��$�����e�뼈ܼa�ȼ����Ԡ�d���79���w��(n�;�i��ph���h��i�e�j�>tl��o�2%t��}�����-��j⡼����lʼ��߼u��|������"�����C��:�׼�^Ǽ����K���4L���*ȼ`cټ��X �����  �  ���;X��;���;H�<�5<~�Y<�Pz<��<XT�<�Ú<`i�<0�<*��<]�<��<��<��<�%�<��<��<�?�<��~<�j`<a<<��<[��;���;5�u;D�^;��;w�;��;Q<Jc3<�ZD<��F<�:<E� <wC�;���;$<~;m>8;��,;\�];�`�;���;�<<�:<��Y<��r<<�<F��<�3�<c��<E�<�[�<R'�<��<���<�<�m�<��<"�n<nU<�W5<�f<���;:�;j�';#�:�B�:�8;�q;9C�;��;�B<h�<�n<x�;ۻ�;�p6;���9μ���$��-��X���%ѹ�:ϋh;r��;�*�;��<-O<Px<��<��<|Z<��	<ް<��;3[�;$��;�)�;�Z�;��K;�ԛ:��k�+ǻ���=z"��0�
�.� ��nA��һdԝ��x�1�l��%��o�û���{u-��BQ��k��v��r��3a�?\E��D$�ʼ�Wyɻ�י���q�4[L��>���A���O��c�r�z������ݗ�[g��_����ۻXZ�Sz�AP?��f�#���P��	o���2��L����S��2��ꤼ����p���ń�������v��`���2_����мޏڼ�ܼx׼'�ʼ����h7��D���u����s�s�a���U�bO��K��mJ�J�%GJ��K�e�L�TxP�6XW��'c�EPu�xK��F�����.���xNμ7�ۼ��ӷ�1~ܼ�Tϼ����`ٮ��Y�����&[������j��ѻż�ּ�]㼕�鼒�輢�༒�ҼP@�����ŝ�?���)��:+y��p�f�k�
�i�|�i��|j�E�k���m���p��v��1�r߆�<|������谼5ļ7׼-�F6������B����c�P�'�ϼ��������u��z���y���_Ѽ�㼘����  �  �%�;�-<��<�&*<D�F<ed<٤~<�I�<���<�C�<zܛ<��<Z�<z+�<�Ҟ<Mٝ<�>�<�ߙ<�\�<�*�<���<i<�f<�WH<ţ(<�%
<���;���;H��;c��;�g�;��<xY.<v�F<�9U<FCW<	L<��5<)o<J��;�w�;ۣ;���;��;n�;�u<WF%<�gB<N#\<7�p<C!�<
f�<W��<���<�ϋ<3>�<�<�?�<�ʉ<�w�<0҃<@�|<P�l<�bW<A�<<��<��;�q�;8�;x\t;Vn;�>�;���;�c�;�F<�+<��$<x�<�	<��;N�;'�; ,:g��}Z��RS8���:�T1;�r�;�о;���;��<��<�-<�<oI<u�<N�<Pe<��;��;���;J=�;>�;��H;U�:�t �9:(��ۗ��Ի<n ������<����һz���%�j��'3�+�K�Y�z`��M�ܻ�C���0���G���R���P��$C��5-�;��F�������К���V\`���R��S�̟\���l�~3�������p������ǻ����&������9�X`Z��,}��e������Z���֫�\ʩ��B��&&��1��`���xx���z�����Nؑ������a��W���ȼY�ʼ�nƼü����!���z��'��Yu���e��Z��S�/�O�*SM�UAL��sL���M��P�YLU���\�܉g��Yw�pI���x��f�����~q��ך˼	�ѼӺѼ>|˼�,��2������@��jғ�����朜�O9��R����ƼNҼ��׼�5׼��мreż�c��H���#�����P�����}�m@u�)p��zm��gl��l�(n�!�p�'�t�{��!��fĈ�A쑼�ʝ�o
��O����s˼Fټ�:�Ĭ�/���ݼW�Ѽ7rüDm���`��GF��$ݭ������wż��Լؾ��k��  �  �^%<��'<^2<.C<SW<jlk<T~<�D�<�Ѝ<��<�Ɩ<���<J��<���<R��<�8�<>ɘ<�j�<�'�<�ۋ<�I�<0sz<�>g<�Q<'�:<��$<�<��<bA<�q<�L<�1<)+I<��\<�h<�Yj<E�`<tMN<�'6<�O<�<���;_b�;���;��
<��<`2<�G<�Y<�qi<w"v<�<��<ц<�ڈ<��<��<�`�<���<ڱ�<��|<�=r<F�d<�-T<x�@<w�*<y�<1$�;�C�;���;��;�
�;�3�;�<  %<R3<ܗ7<i�0<�N<�V<���;�y�;�K;"�;���:�.;X�<;�|;�e�;@��;\��;�s�;}�<8�<)�<�	<C<�&<�;[K�;��;8�;�;޾y;�D/;�C�:���?�ֺ�-O��Ǔ�®���Ż�û���]���S�P�3���ĺ���G4
��{\�����]�]�^�M�)�Mu*��"��e���H=⻦���������Ʂ�td{�ͳt�T*v�����㉻ש���«��Z»p#ܻҒ������~!�X8�;�P�J�j�1ၼ�{���ߓ�G���8c����������VM{�l���d�CJg�j�t��c��j���ɠ��K���ĳ�M��yﳼ���k����������Z��H�|���o�ؗe���]�|�W��6S�W�P��Q�ӤS�
OX���^��/g���q�)3��ه������q�����Ӱ���x��툽�����9���^g���袼��������;���E��ꡑ�k������\���:罼�üUü�'��݆��ح����ٟ��I󐼕ω�U1������Hy�ѝt�r�q�*,q���r��w�=}�$�����������0���Q��Tר��4��Gs���Fɼ�=м\Ӽ91Ѽ��ʼ\����,��Ó��4:��2Ơ�Oף����|��/=ļٸϼ^�׼�  �  Q�M<,�K<]zO<H�V<��`<�3k<z�u<��<K�<׻�<�f�<Გ<�.�<oE�<�z�<��<�<��<���<ڣ�<�:y<��l<MR`<nnS<�F<&
;<�1<u-<�-<��4<U�A<̀R<B;d<�Bs<�F|<�9}<"�u<�g<d;T<o�@<p�/<xM$<��<E�<�#%<?.<ݥ8<��C<��N<zqY<��c<n<J�w<�_�<Eσ<���<r��<t�<=i<��u<�
k<��_<DST<�zH<�3<<��/<5#<<:�<!�<K�<��<3!<e0<><��G<�J<q�C<��4<=_<��<W��;�;�;u��;J?�;�;0#�;�#�;�զ;]��;r�;���;Y�;P��;���;2�;���;u��;���; 6�;�;�v�;�q;�2;?-�:�S:�U#�d	���r��D6���Z�U	k���c�$�D������!�4�6?��fP��_m�Y ��Z�q��p�ɻ��f�����Ǡ�+� ������⻜ ӻ�bĻ�ζ��T��y"��������MS�������n���;»��޻U���Y������.���>���N���^�Upm�5�y����}���W���vy��m�X�_�VpU�z�P��T�i�_�B�q��܃�����|��D6��U���z͢��X�����PᖼR��ŋ��V�����ܐw�,|m��`d�gF]�WY�>bY��u]���d�8an��y����ʇ�8���l���'ݙ�m؟�f��wʨ�B$��R���)ˣ��o��i���'Ԋ����ƿ����������َ����
��uǩ������g��BG��	����J��������Ah���W���i��~���D��N>��g+{�[y��{�p����f��ϊ�
���\���پ������v����J��@0��|���+��Rü��S��L������k����#��Gb���㙼�G��n\��"c�������ü�  �  >]o<��h<0d<V�a<�n`<&�`<��b<@g<��n<K�x<�y�<ˈ<t=�<��<�H�<�ҏ<���<��<;mx<>j<`R^<AU<� O<QK<?�H<`H<��H<z:K<�XP<h]X<bc<y�o<�[|<]w�<���<>ʆ<��<M}<M+o<f`<��R<f�G<ff?<��9< �6<�5<��4<�(6<O�9<�?<�H<T<<Pa<cPn<�x<y�~<}�~<�fx<�gm<��_<RUQ<�sD<~:<}2<~-<x*<��(<�K(<#)<=�+<�i0<{�7<�@<�K<�,T<��Y<Z<L�S<��G<�w6<��"<�Q<�%�;�u�;).�;s��;�ʧ;N�;P��;��;�;b��; ��;NY�;���;L��;.��;��;'��;�f�;-��;��S;�;�}�:Z�9L�˹
_�������8�ͺ-VԺ��ɺ8����l��K͹�y9�:.GP:�{,:^9��:��캇C��f�������j���Ի�F�%����sL���T��N����L��߻v�λ+|��U/��"R��.��LŻ!�⻤���2�o)�dI9�0�E���O���V��+\�L,`��b�(�c�iOb�$G^���W�[�O�yG�InA���?�	pC��
M��h[�ޅl�B~�R���4o��ZE������ă��3���������V���=��Ƨ��a�������v��l��f���e�^�k�K�v��?��X�������┼	��������Y���񜼏᜼%
��)%���ꖼ/B��k]��rЅ��$�ƚu��q�Εr�8z�����M������&���C������q���䤼	���٥��ݤ���������J���������{ˈ�����;䂼�P��&���������ݝ��C��0M���欼�A��쩰�Z���Z���{���r��� ���$���/���י�?-��Y���?��x:�����+����G��݉��b����  �  ��<�'{<&1n<�Ba<�8U<�qK<n�E<9E<SK<��V<��f<��x<��<��<%�<���<�
�<�fm<FtY<�G<�:<4<Ye3<�7<R@<J<�T<�^_<��i<�s<s}<�p�<,��<� �<�	�<��<F��<�7�<�M�<F�y<n<�>b<7:V<��I<DX=<B1<� &<�<"j<$�<6%<�Q3<��D<B�V<X�e<��m<�n<[�e<8�V<��C<;�0<�:!<��<�<3O<}x<Xs#<͢-<��7<��A<�sJ<q�R<< Z<��`<e<V�g<�&f<f4`<V<��H<�>9<��(<�<�<�6�;�E�;��;�u�;Nf;I�<;r ';f4);bC;�p;�;��;z��;`f�;��;�֋;��?;9ӽ:[�R8�����s����2���p)ź�D���y
��-��>��9��C:��:U��:Q��:��:T;�:Jw:5�9`%�o�ǺЫ"�ņa�����P���λ	�� J����Y����E?����(Q�@ﻵ�ػ�Uͻ�һ/��$Z�>�i�5��K��\\���f�0�j�C�i� �d�i�]��lV�VHO���H�ԭB�-=��8��4���1�(b2�i�6�`�>���I���V���d��or�������s��n��Vp��������Fܥ�'���UH��e���)�����/�n�v�pv���~�_Ɇ��"�� ���`Q��1q��0t��턧��E��~�����������	��C���K����:� �u��cm��Fg���d���e�sk��ws��}������m���j������@✼3H��2j��w���#B���Y��Uf���^��-ؤ��	��2���~���|���Ό�Y����F��^=������A���{���ѻ�y^���۶�R!���䬼=���;z��с��������������������>��є������f����@���$��*0���  �  �<Ӭ�<��m<#W<��@<�-<[%!<�<�b"<��0<ՕE<��\<�q<__~<���<5�y<h<~=P<?�6<r� <��<�N<�7<�9<m�-<(B<�V<e(i<�y<o߂<�Ӈ<���<rn�<H_�<S�<��<���<<�<�ى<��<�9�<�&s<��b<v|O<��9<�f#<�w<���;֞�;,��;d'�;�<�[%<��<<e�O<�Z<��Z<�OP<k�<<w�$<\�<���;���;��;=o�;�<�t<��(<vN<<�9M<ϽZ<��d<��k<��o<�{q<��p<��m<�5h<��_<]@U<��H<S�:<�V*<�|<��<d&�;�Z�;�hW;*�:2�F:�9�!�8~:�V�:Xp.;�Vu;L/�;���;��;E�=;1�:���$���>h�׌�٦���u���S�������U2�� vL:�:���:��;Sm;��;ݵ;�m�:�q�:�?q:I��9���)������g��V����ϻ9�"���8/�z>�VpE�C���7��&���Z3�S���)�����a��H:���W��r��l������Ն�`z��p�v�łe�fhT��;E�\9��T0���*��w'��T&���&��~)�*&.���4�n=��wG��R���_�F�n�Q^��}������4��cɫ�9!��߸�����R���p���~���i���䄼.����������j���>���I@���ຼ�����������h��Q-�����cw��%�v��vm��Of��a�̒]��@\�P^]���`��kf���m�?w�)R��܅��pJ��ₛ���������	��aü�	Ǽ��ż����h���쪼��ݗ��x�����cޝ�|�������Px��LIʼֹμ
XμЙɼ����oҷ���V����Ĕ��s��f���_��3>����������#��gm�������Ϗ�S���0U���  �  ���<���<Tf<nF<�Z'<��<���;i-�;���;\�
<M�$<��@<=Z< rj<.|n<q(e<�P<�g3<߻<1K�;�Q�;���;�;nB�;{I<�3<"�P<��j<e�<�ɇ<�1�<���<z��<�w�<羓<6h�<�r�<�ې<�v�<�ي<@w�<�{<�f<�M<10/<u�<Ў�;��;w��;Y��;ک;���;"$<�"<�2:<�oG<&�G<��:<t#<�<���;�բ;]��;@N�; R�;6��;�m�;�< �8<DtP<ߋb<m�n<l�u<l�x<|�x<UGv<�9r<��l<ioe<s�\<�IR<�E<`4<\k<k�<R��;��;�l�:�#���Ǻ����"��C���#�p�`:87;�4Q;�&a;)�;;0a�:��ƹ��$�=����,Ż1j߻l�߻d�ǻ�S��#_U���Ӻ?����Ȑ:�;_�%;pe6;�8;&�0;,";n�;���:�(�:[�I:Z"�8�"@����!Q��˟�g�߻��.n3��}P�lMe���n�R�k���]�6�G�/�����`��,��5�c�V�ƻy�y4���㖼 k��ֈ��x!��I놼�s��Z�U�C��2��E&�G���E�?��P� �d$�!Q)��5/�6�	>��H�� U��_f��~|���������謁�ӹ�P�ż��̼��ͼ�_ȼ̗����������I������PV��4���0S���﮼�����)ɼ��ϼ��ϼ��ɼ�'��}=���7��Kԓ��V����z�'|l���b�J�\�֌Y���W�ϢW��X�t�Z�^���c�ySl�Y�x�鄼�:�����{��<��m˼�ּ sۼ�ڼ��Ӽ�Ǽ����(��;������ o���'��g���_�żD$Լ��޼�t�4��G�ڼ��μ���3ﱼzZ������p<��) ���7�������ւ��v��������� !���`���������������  �  ��<^�~<�D[<��4<��<�}�;;�;��;ze�;ZC�;:~<�m)<�jF<QY<#^<ϛS<g�;<3�<�D�;\	�;��;�;};js�;���;�C�;�I#<�.G<p%g<)n�<༉<���<��<���<d �<��<"z�<�Ǔ<���<�ϐ<rr�<KƇ<X~<٭e<NqF<"<�e�;�;{j;�M$;��;��I;���;�!�;H�<؋'<��6<{&7<�(<��<��;|�;��<;� ; R ;_>:;ؑ;�j�;��<g`1<��N<�d<�s<��z<}X}<�%|<3�x<�t<��n<Ah<ǌ`<��V<��I<]�7<0�<X� <1Զ;.�H;�N:���2j��Q��+�~����2���}:Q�	;w;c��:�\�9	��ES��.4ӻ�{�
���w���� �л������I<�HR�:��;�?9;�K;`�J;�d>;��+;�;�s�:<��:�Ά:��9n$�,�Ӻ��P�P���p����#��#L��	o�샼Ԃ��
���~��c���F�|�-������a�-�/�I�Jo�LH����������\D��5M��i����d��񁼄Rc���F���0��2"��`���g���>���!�8�&��Z,��,2�F*9��B��^P���c���}���5����𴼣%Ǽ�ռ�l޼��߼&�ټ
ͼѼ��+������X喼�����֝�N-��������̼@ڼJ�Ἴ���<ڼ��̼L����'��[u��I6��%�x�wh���]�wX���U��,U�9xU��_V�m�W�iwZ�u_�3.g�(�t�+�������\��S6��pȼ��ټ#��^�v켃K伓�ּ�)Ƽ����^ ���4���証�ϲ��¼��Ӽ8�4&�����O�꼸xۼO�ɼE���������𨎼ɱ������ก�� ���7��l����f���z���/���!��������  �  *�<Еy<�0R<I)'<���;���;%J�;YW[;h+y;r��;" �;s�</(9</�M<YS<d�G<u�-<RS
<�	�;D�;4=3;��;�CE;�8�;�{�;��<�?<��b<��<��<y��<��<Sg�<坕<%[�<��<�P�<�k�<պ�<�d�<l�<��}<��b<@<��<.t�;Dڈ;�{;�m�:��Z:
��:�NY;yX�;�k�;��<j|+<��+<B&<)1�;I�;IvV;�j�:<�9���9���:`BU;iW�;��<�*<�DK<��c<%t<V�|<�<�~}<�y<��t<�Ao<�i<��a<��X<�K<>�8<ߏ<�/�;�:�;V;,O�&eG�����Eǻj�ɻ�㬻�	p�}����8d�:��:�$�:�;�@�2�\��� ���"�D,�;`*�����/��V}��T>��%I���|:��;�R?;�R;�Q;��C;{�/;�L;�b;���:��:VH	:{1��M5Ѻ�jX�ܖ�����`1��^��A��ُ��ٕ�9�������v��nV�+�:��*�>�)��A9�S�W�bv�2������j����|��������Vƚ��!��NYk��K���1��X!������c��F���� ���%��)+�R�0�^97�+�@�P�N�l�c��'����������d���м9��ߊ�O��A�1�׼O�ż�����㤼����Z5������{����ļ�׼���������Ǒ���ּ�hüʩ��'ؚ��ɉ�p#y���f�n�[�=V��AT�<T�1�T��wU�e�V�p�X�Z#]�/fe��s�3������3���6����м0��\����u�����B���μP����"��P«�����~R���ɼ��ܼ ������ ��M��B�������мY������o%��ԏ����,���oր��q��궀��<���遼�т�FR���*���T��{����  �  :��<�uw<�N<�#"<0��;=3�;��^;BS8;(PW;�(�;���;�<�y4<"�I<�O<�C<H)<3~<�,�;�j;��;3��:-�#;D�;+�;r<�;<�a<V�~<�<�Ð<C�<���<�ĕ<Kz�<��<�s�<:��<H�<���<?~�<Fv}<�a<I�=<�<�e�;Z�u;L��:"�:�I�9q��:��;;㳦;��;�<��'<;�'<��<���;���;{K9;��}:����AD��Z8{:��8;R�;�Y�;�'<��I<Lrc<�2t<��|<�n<1�}<K�y<t�t<�oo<zXi<yJb<Y<��K<e�8<��<���;_�;w;�Zb��d��^���ػ�/ۻ*���/���&�ǗL�ic�:��:ݧg:�{>��H�s��M��~�%�{�4���2�_ ��8��յ���L��?m��qk:C�;'<@;vT;`=S;E;d�0;/(;�P;( �:P �::��9�Һ�}\��㷻lf��j6���d��������;��Wԗ��ύ��U}��\��?��.�lp-��e=��Y\�˞��q��h���%ٸ��Խ�M��⫮�e؝��t����n���L��2��_!�R/�Ώ�?a����� �K�%���*�U60�[�6�&G@�R�N��:d��΀��X�����q%��%ԼM���i�b�b<ۼ��ȼgA�����܃��/���5�������Ǽ`�ڼ����?��'򼽡�k*ڼ�AƼ���4��y�����y��f�vf[�&�U�"�S���S�,\T�Z:U�'nV�D}X�]�\��e���s� ��zt�������x����Ӽ	�缼���������� ������ѼH���A�����@�������@�̼Y8��� �����������I|ӼjX���ܪ�g���б��dՆ��x��c����G��ѕ��o��gɁ�������a���4��Yٔ��  �  *�<Еy<�0R<I)'<���;���;%J�;YW[;h+y;r��;" �;s�</(9</�M<YS<d�G<u�-<RS
<�	�;D�;4=3;��;�CE;�8�;�{�;��<�?<��b<��<��<y��<��<Sg�<坕<%[�<��<�P�<�k�<պ�<�d�<l�<��}<��b<@<��<.t�;Dڈ;�{;�m�:��Z:
��:�NY;yX�;�k�;��<j|+<��+<B&<)1�;I�;IvV;�j�:�;�9���9���:_BU;iW�;��<�*<�DK<��c<%t<Y�|<�<�~}<�y<�t<�Ao<i<��a<ϴX<#�K<W�8<��<�/�;;�;zV;EM��dG�ֲ���Eǻ9�ɻ�㬻L	p��|���8�d�:��:�$�:�<�p�2�-\��� ���"�)D,�W`*����0���}���>�Q'I�+�|:O�;WR?;��R;�Q;��C;f�/;�L;c;ӡ�:;�:TI	:/���4Ѻ]jX�������� `1��^��A��ُ��ٕ�-����󉼮�v��nV�"�:��*�=�)��A9�\�W�ov�;������v����|�������eƚ�"��lYk�K���1��X!�����t��T���� ���%��)+�W�0�b97�.�@�R�N�m�c��'����������d���м9��ߊ�O��A�1�׼O�ż�����㤼����Z5������{����ļ�׼���������Ǒ���ּ�hüʩ��'ؚ��ɉ�p#y���f�n�[�=V��AT�<T�1�T��wU�e�V�p�X�Z#]�/fe��s�3������3���6����м0��\����u�����B���μP����"��P«�����~R���ɼ��ܼ ������ ��M��B�������мY������o%��ԏ����,���oր��q��궀��<���遼�т�FR���*���T��{����  �  ��<^�~<�D[<��4<��<�}�;;�;��;ze�;ZC�;:~<�m)<�jF<QY<#^<ϛS<g�;<3�<�D�;\	�;��;�;};js�;���;�C�;�I#<�.G<p%g<)n�<༉<���<��<���<d �<��<"z�<�Ǔ<���<�ϐ<rr�<KƇ<X~<٭e<NqF<"<�e�;�;{j;�M$;��;��I;���;�!�;H�<؋'<��6<{&7<�(<��<��;|�;��<;� ;�Q ;^>:;ؑ;�j�;��<g`1<��N<�d<s<��z<�X}<�%|<A�x<�t<��n<]h<�`<��V<	�I<��7<d�<�� <�Զ;�H;�R:��2j�+� ����~����2���}:~�	;!w;2��:�Z�9ÿ麃S��{4ӻ|�<��-x����v�л0�����:C乪P�:	�;�>9;KK;��J;�d>;��+;�;�s�:���:�φ:���9��ʣӺ#�P��O��:p��Z�#��#L��	o��냼����󡇼�~�ɼc���F�j�-������j�-�@�I�co�]H��͡�����vD��QM������e��)񁼿Rc���F���0��2"��`������>���!�K�&��Z,��,2�N*9��B��^P���c���}���5����𴼣%Ǽ�ռ�l޼��߼&�ټ	ͼѼ��+������X喼�����֝�N-��������̼@ڼJ�Ἴ���<ڼ��̼L����'��[u��I6��%�x�wh���]�wX���U��,U�9xU��_V�m�W�iwZ�u_�3.g�(�t�+�������\��S6��pȼ��ټ#��^�v켃K伓�ּ�)Ƽ����^ ���4���証�ϲ��¼��Ӽ8�4&�����O�꼸xۼO�ɼE���������𨎼ɱ������ก�� ���7��l����f���z���/���!��������  �  ���<���<Tf<nF<�Z'<��<���;i-�;���;\�
<M�$<��@<=Z< rj<.|n<q(e<�P<�g3<߻<1K�;�Q�;���;�;nB�;{I<�3<"�P<��j<e�<�ɇ<�1�<���<z��<�w�<羓<6h�<�r�<�ې<�v�<�ي<@w�<�{<�f<�M<10/<u�<Ў�;��;v��;Y��;ک;���;"$<�"<�2:<�oG<&�G<��:<t#<�<���;�բ;]��;?N�;R�;6��;�m�;�< �8<EtP<�b<q�n<s�u<w�x<��x<iGv<:r<��l<�oe<��\<�IR<*E<�4<�k<��<��;%��;-o�:��x�Ǻ����"��A�½#�ޟ`:�7;>5Q;�&a;�;;�`�:��ƹ_�$�����-Ż�j߻�߻�ǻfT��p`U�3�Ӻ�
��]Ɛ:�;w�%;�d6;K�8;��0;�+";c�;@��:�)�:f�I:.8�8_@���� Q�Z˟�Ǌ߻����m3�<}P�Me�f�n��k�Ļ]��G��/������`��,�#�5���V���y��4���㖼Dk�������!��s놼q�s�  Z���C�(2��E&����F�o��x� �0d$�;Q)��5/�6�>��H�� U��_f��~|���������謁�ӹ�P�ż��̼��ͼ�_ȼ̗����������I�����PV��4���0S���﮼�����)ɼ��ϼ��ϼ��ɼ�'��}=���7��Kԓ��V����z�'|l���b�J�\�֌Y���W�ϢW��X�t�Z�^���c�ySl�Y�x�鄼�:�����{��<��m˼�ּ sۼ�ڼ��Ӽ�Ǽ����(��;������ o���'��g���_�żD$Լ��޼�t�4��G�ڼ��μ���3ﱼzZ������p<��) ���7�������ւ��v��������� !���`���������������  �  �<Ӭ�<��m<#W<��@<�-<[%!<�<�b"<��0<ՕE<��\<�q<__~<���<5�y<h<~=P<?�6<r� <��<�N<�7<�9<m�-<(B<�V<e(i<�y<o߂<�Ӈ<���<rn�<H_�<S�<��<���<<�<�ى<��<�9�<�&s<��b<v|O<��9<�f#<�w<���;֞�;,��;d'�;�<�[%<��<<e�O<�Z<��Z<�OP<j�<<w�$<\�<���;���;��;<o�;�<�t<��(<vN<<�9M<ҽZ<��d<��k<��o<�{q<��p<��m<%6h<��_<�@U<1�H<��:<PW*<)}<�<+'�;�[�;kjW;I�:.�F:*9mJ�8��:�X�:q.;.Wu;s/�;��;��;߬=;�/�:��,���?h��׌�����cv����S����� ��zb��apL:��:���:��;�l;g�;��;pm�:Rr�:<Aq:S��9���s'�������g��U��Ūϻ�8����N8/�>��oE�� C���7���&���;3�3���)�������H:��W�r�"m����.ֆ��z��ؔv�,�e��hT�<E��9��T0��*�:x'��T&���&�)�K&.���4��=�xG�%�R���_�I�n�Q^��}������4��bɫ�9!��߸�����R���p���~���i���䄼.����������j���>���I@���ຼ�����������h��Q-�����cw��%�v��vm��Of��a�̒]��@\�P^]���`��kf���m�?w�)R��܅��pJ��ₛ���������	��aü�	Ǽ��ż����h���쪼��ݗ��x�����cޝ�|�������Px��LIʼֹμ
XμЙɼ����oҷ���V����Ĕ��s��f���_��3>����������#��gm�������Ϗ�S���0U���  �  ��<�'{<&1n<�Ba<�8U<�qK<n�E<9E<SK<��V<��f<��x<��<��<%�<���<�
�<�fm<FtY<�G<�:<4<Ye3<�7<R@<J<�T<�^_<��i<�s<s}<�p�<,��<� �<�	�<��<F��<�7�<�M�<F�y<n<�>b<7:V<��I<DX=<B1<� &<�<"j<$�<6%<�Q3<��D<B�V<X�e<��m<�n<[�e<8�V<��C<;�0<�:!<��<�<2O<|x<Xs#<͢-<��7<��A<�sJ<w�R<F Z<��`<ցe<r�g<�&f<�4`<GV<ݤH<?9<��(<$�<"<w7�;�F�;���;dv�;f;��<;"';�5);�C;
p;n�;7�;���;jf�;��;�֋;��?;]ѽ:cR8�����"���������� -źEH����
��_��ْ�9�C:	~�:��:-��:}��:6;�:�Jw:��9�"���Ǻ��"�m�a�����O��4�λ'��I�J��������>�?���P��?�r�ػ�Uͻ�һO��DZ�n���5�X�K��\\��f���j���i���d���]�jmV��HO�\�H�4�B��=�8��4���1�Vb2���6�|�>���I���V���d��or�������s��n��Vp��������Fܥ�'���UH��e���)�����/�m�v�pv���~�_Ɇ��"�� ���`Q��1q��0t��턧��E��~�����������	��C���K����:� �u��cm��Fg���d���e�sk��ws��}������m���j������@✼3H��2j��w���#B���Y��Uf���^��-ؤ��	��2���~���|���Ό�Y����F��^=������A���{���ѻ�y^���۶�R!���䬼=���;z��с��������������������>��є������f����@���$��*0���  �  >]o<��h<0d<V�a<�n`<&�`<��b<@g<��n<K�x<�y�<ˈ<t=�<��<�H�<�ҏ<���<��<;mx<>j<`R^<AU<� O<QK<?�H<`H<��H<z:K<�XP<h]X<bc<y�o<�[|<]w�<���<>ʆ<��<M}<M+o<f`<��R<f�G<ff?<��9< �6<�5<��4<�(6<O�9<�?<�H<T<<Pa<bPn<�x<y�~<}�~<�fx<�gm<��_<QUQ<�sD<~:<}2<~-<x*<��(<�K(<$)<?�+<�i0<��7<�@<�K<-T<��Y<&Z<z�S<.�G<1x6<5�"<$R<�&�;yv�;/�;Y��;�˧;�N�;6;���;«�;��;Ŏ�;�Y�;e��;���;Z��;��;��;�f�;Ҁ�;��S;Q�;�z�:��9Ï˹'	_�H��M����ͺ�YԺ�ɺ-��*�l��T͹�k9��:�EP:D{,:na9��:�r캌C�Sf������i��� Ի�E�<��+��K���S������L��߻��λ�{��/���Q��-��mŻd������2��)��I9���E��O�(�V�j,\��,`���b���c��Ob��G^�'�W���O�HyG��nA�ܡ?�/pC��
M��h[��l�L~�U���6o��[E������ă��2���치�����V���=��Ƨ��`�������v��l��f���e�^�k�J�v��?��X�������┼	��������Y���񜼏᜼%
��)%���ꖼ/B��k]��rЅ��$�ƚu��q�Εr�8z�����M������&���C������q���䤼	���٥��ݤ���������J���������{ˈ�����;䂼�P��&���������ݝ��C��0M���欼�A��쩰�Z���Z���{���r��� ���$���/���י�?-��Y���?��x:�����+����G��݉��b����  �  Q�M<,�K<]zO<H�V<��`<�3k<z�u<��<K�<׻�<�f�<Გ<�.�<oE�<�z�<��<�<��<���<ڣ�<�:y<��l<MR`<nnS<�F<&
;<�1<u-<�-<��4<U�A<̀R<B;d<�Bs<�F|<�9}<"�u<�g<d;T<o�@<p�/<xM$<��<E�<�#%<?.<ݥ8<��C<��N<zqY<��c<n<J�w<�_�<Eσ<���<r��<t�<=i<��u<�
k<��_<DST<�zH<�3<<��/<5#<<;�<$�<O�<��<3!<t0<'><��G<�J<��C<��4<~_<�<���;�<�;?��;!@�;��;$�;�$�;�֦;3��;�r�;���;�Y�;ֿ�;��;_2�;Ȱ�;~��;���;�5�;��;Sv�;��q;v~2;B*�:\S:*q#�����t�|F6���Z��
k��c�f�D���d��q�4��A���P���m�� �0Z��p����ɻ���#��Y���� ��������ӻ�aĻ*ζ�AT���!��I��د��*S�������n��.<»1�޻�������v���.�^�>�N�N���^��pm���y����������wy�!m���_��pU���P��T���_�W�q�݃�����|��F6��V���z͢��X�����PᖼR�� ŋ��V�����ܐw�,|m��`d�gF]�WY�=bY��u]���d�8an��y����ʇ�8���l���'ݙ�m؟�f��wʨ�B$��R���)ˣ��o��i���'Ԋ����ƿ����������َ����
��uǩ������g��BG��	����J��������Ah���W���i��~���D��N>��g+{�[y��{�p����f��ϊ�
���\���پ������v����J��@0��|���+��Rü��S��L������k����#��Gb���㙼�G��n\��"c�������ü�  �  �^%<��'<^2<.C<SW<jlk<T~<�D�<�Ѝ<��<�Ɩ<���<J��<���<R��<�8�<>ɘ<�j�<�'�<�ۋ<�I�<0sz<�>g<�Q<'�:<��$<�<��<bA<�q<�L<�1<)+I<��\<�h<�Yj<E�`<tMN<�'6<�O<�<���;_b�;���;��
<��<`2<�G<�Y<�qi<w"v<�<��<ц<�ڈ<��<��<�`�<���<ڱ�<��|<�=r<F�d<�-T<x�@<v�*<y�<1$�;�C�;���;��;�
�;�3�;�<3 %<k3<��7<��0<�N<�V<:��;�z�;8K;��;���:0;��<;��|;f�; ��;��;Et�;��<t�<X�<�	</C<�&<�;)K�;���;��;��;��y;�C/;�@�:�P��k�ֺ~/O��ȓ�������Ż��û���������P��3�/�ĺ��4
��{\�w��s]�����)��t*���"�Xe�!��<����O��G��a����c{��t��)v�����㉻󩘻2ë�#[»�#ܻ[�����'!��8���P���j�eၼ�{���ߓ�v���dc��̖�������M{�;l���d�eJg���t��c��q���ɠ��K���ĳ�M��yﳼ���k����������Z��H�|���o�ؗe���]�|�W��6S�W�P��Q�ӤS�	OX���^��/g���q�)3��ه������q�����Ӱ���x��툽�����9���^g���袼��������;���E��ꡑ�k������\���:罼�üUü�'��݆��ح����ٟ��I󐼕ω�U1������Hy�ѝt�r�q�*,q���r��w�=}�$�����������0���Q��Tר��4��Gs���Fɼ�=м\Ӽ91Ѽ��ʼ\����,��Ó��4:��2Ơ�Oף����|��/=ļٸϼ^�׼�  �  �%�;�-<��<�&*<D�F<ed<٤~<�I�<���<�C�<zܛ<��<Z�<z+�<�Ҟ<Mٝ<�>�<�ߙ<�\�<�*�<���<i<�f<�WH<ţ(<�%
<���;���;H��;c��;�g�;��<xY.<v�F<�9U<FCW<	L<��5<)o<J��;�w�;ۣ;���;��;n�;�u<WF%<�gB<N#\<7�p<C!�<
f�<W��<���<�ϋ<3>�<�<�?�<�ʉ<�w�<0҃<?�|<P�l<�bW<A�<<��<��;�q�;9�;\t;Vn;�>�;��;�c�;�F<�+<��$<��</�	<r��;�N�;�;F�,:�]���U���S8U��:�U1;gs�;cѾ;r��;
�<�<�-<<�I<��<R�<Ge<���;��;E��;�<�;� �;��H;�|�:�y ��;(��ܗ��Ի�n ��������)�һȇ����j��'3�͕+�$�Y�N`��
�ܻ�C���0���G�`�R�b�P��$C��5-�������`���4К����v[`��R�,S�l�\�o�l�}3��ћ���p�����q�ǻ��9'�'��>�9��`Z��,}��e��ʷ������<֫�ʩ��B��B&��.1��`���xx���z�����Vؑ������a��Y���ȼZ�ʼ�nƼü����!���z��'��Yu���e��Z��S�/�O�*SM�TAL��sL���M��P�YLU���\�܉g��Yw�pI���x��f�����~q��ך˼	�ѼӺѼ>|˼�,��2������@��jғ�����朜�O9��R����ƼNҼ��׼�5׼��мreż�c��H���#�����P�����}�m@u�)p��zm��gl��l�(n�!�p�'�t�{��!��fĈ�A쑼�ʝ�o
��O����s˼Fټ�:�Ĭ�/���ݼW�Ѽ7rüDm���`��GF��$ݭ������wż��Լؾ��k��  �  ���;X��;���;H�<�5<~�Y<�Pz<��<XT�<�Ú<`i�<0�<*��<]�<��<��<��<�%�<��<��<�?�<��~<�j`<a<<��<[��;���;5�u;D�^;��;w�;��;Q<Jc3<�ZD<��F<�:<E� <wC�;���;$<~;m>8;��,;\�];�`�;���;�<<�:<��Y<��r<<�<F��<�3�<c��<E�<�[�<R'�<��<���<�<�m�<��<"�n<nU<�W5<�f<���;:�;l�';#�:�B�:�8;�q;HC�;��;�B<{�<o<Ux�;��;Nq6;7��9�̼��$�-��V��nѹ�	�:��h;���;+�;�<VO<rx<��<��<�Z<��	<ٰ<���;[�;���;�)�;-Z�;��K;/ӛ:��k��ǻ��uz"��0�9�.�I���A�+һ�ԝ�-�x�9�l�s%��P�û���[u-�hBQ��k�Ϸv���r��3a�\E�OD$�����xɻrי�$�q��ZL���>���A�G�O���c�p�z������ݗ��g������[�ۻ�Z��z�xP?�J�f�&#���P��'o���2��g���T���2��ꤼ÷��~���ń�������v��d���5_����мߏڼ�ܼx׼'�ʼ����h7��D���u����s�s�a���U�bO��K��mJ�J�$GJ��K�e�L�TxP�6XW��'c�EPu�xK��F�����.���xNμ7�ۼ��ӷ�1~ܼ�Tϼ����`ٮ��Y�����&[������j��ѻż�ּ�]㼕�鼒�輢�༒�ҼP@�����ŝ�?���)��:+y��p�f�k�
�i�|�i��|j�E�k���m���p��v��1�r߆�<|������谼5ļ7׼-�F6������B����c�P�'�ϼ��������u��z���y���_Ѽ�㼘����  �  �d};)K�;5J�;zN <CK(<|�P<Xtu<䫉<B��<㓛<Z`�< �<^)�<-ؠ<`O�<z��<1��<�
�<��<L�<�K�<��|<z�Z<E�2<`u<E��;�An;ф;l��:kS%;�@�;zE�;�<G{&<�8<k�;<;.<-a<�2�;庐;m)#;$��:#��:�K;�-p;���;u{
<��2<��U<B�q<ϸ�<��<�&�<ހ�<�ڍ<,ύ<��<n:�<B�<@׊<�\�<��<:n<["R<Ud.<�1<nz�;��I;޾�:x�8K��V:��;�ґ;v��;3( <5�	<P</y�;���;���:�L^���;�E���ꆻ3�S���ʺ��!:�?;N��;f�;��<U�<�o<��<k<�l<&�
<*�<�L�;���;%��;ak�;a��;r�E;s(o:aiҺ�!���v黊���:��H�U�F���5�����C��rΓ��f���K���s޻���v@��!g�z��b����E��gav���V�Iu1����Y!ӻ�'����o���E�m�6��:;�] K�u`��mw�Q��rQ������f���ٻrc���cE�4fp�M��ۙ���p��Gż:Yʼ�3Ǽ
�!.���x�����������B��h�������J���y˼d[ܼ���@��
��ռ��¼)������R��J�t�-�`�e�S��-M�j6J�	EI�'I��fI�m J��[K�h�N��U��b�#�u�"���vŚ�vC����ļ.ؼ�`缢�＀��)���ټ~�Ǽ����}����������[������μ	
Ἑ��$�����e�뼈ܼa�ȼ����Ԡ�d���79���w��(n�;�i��ph���h��i�e�j�>tl��o�2%t��}�����-��j⡼����lʼ��߼u��|������"�����C��:�׼�^Ǽ����K���4L���*ȼ`cټ��X �����  �  �<2�<P��<O�<k
�<b��<ַ�<��<���<(��<�E�<�q�<�'�<���<w+�<<��<k��<��<�o�<D~�<�a�<͒�<@�<�N�<y�<1��<��t<�-g<�b<�dh<��v<�I�<���<cΘ<+(�<�Ǟ<wv�<}�<�ن<]�v<чc<��W<4�U<
�]<� n<�ށ<�Ѝ<UC�<���<��<@t�<�_�<V��<�ɯ<�ɮ<��<A��<�ܭ<%H�<��<�ݭ<���<�ͦ<�@�<		�< ��<��w<^�_<1L<�x@<�3><oQE<��S<*'f<�w<(�<��<~�<̿q<��Y<HD><�[#<��<�� <��;��<�?<b&<�:<�M<$[<��c<9�f<"�d<}�_<{Y<�+R<��K<=PF<X�A<�=<��8<Q�1<~'<	=<�<���;�ߜ;��H;���: L�9���q���9ߵ�:F;�I;Gn;��n;ױG;V�:Q��99��;��]��}��9����z��x6��ʺdĝ�neH:���:�'�:��;6��:	d�:���:�m/:G��9�^��B���S�&Gb���������L���%pȻ��5�-u5���F�1�N��L���B���2�l�!�87�Д��6��w�D�0���I��vc���x�&#���ل��n���cs�2+^�[�F���/�8u��� F�/F��� � ����B�����;��@����X��O	����j|!�Ρ5���M���f�Bi~��q������)���y���
����l�7X�x4H�3W@�SB���M�
a�x��&��H���*��t����������]s�2�[��#F���4��(��"�� �(!�NV#�C�%�"�'��}(��(��@(��(�"�+�a42��=�ZZO�Øe���~��F��m���f���D壼]͢���T瓼�\��4y�0Cr���m�d�s�$2��6͋�����&4������  �  �M�<�b�<�ь<�b�<���<۞�<�b�<*ݽ<���< ��<O�<U��<�L�<\&�<�_�<��<��<l�<x�<��<>��<(��<|Ǫ<�q�<�	�<��<ٗy<�-l<]�g<�7m<C {<E�<H`�<��<�E�<`ߟ<T��<US�<x��<q�z<B'h<�\<��Z<��b<�Er<���<�#�<*-�<�<2`�<m��<�h�<���<��<��<�5�<��<��<�c�<���<��<���<��<ş<f�<�$�<R{<q�c<n�P<߁E<�2C<(�I<��W<&�i<v�z<^D�< �<��<�)t<s�\<1�A<'�'<q<��<��<�I	<�@<
�)<+�<<~�N<�\<d<еf<�d<��_<-WY<��R</L<��F<�
B<a�=<Q�8<� 2<��'<��<�<�;�;�ZW;	I�:0�%:�Wh�D�w�D�9�ĩ:�;��S;�-w;��w;��P;wS;�:�͏��i)��7q�y]���F���h�'o'�������6�%�]:���:�� ;4;�K�:
��:�h�:��5:7y�9\857㈹8�
��`�tî��C��I�g����û����:��0�H�A���I�`H�YL>��3/���@��[Q����s�O.���F�Li_��+t�i����M���~�Yo��Z�D�C�j�-�vV�ދ� ��2��� � ��8��p��O�}��~�������	�7��q ���3�K��pc��7z�I���$������"����}��i�NhU�'�E�'&>��@�zK��&^��|t�x���P������𐼮���A�$p�iY�C�D���3�>(��!�V ��� �3#�4s%��9'�X(�4(��(�w�(��y+���1�@Q=�N���c�|�_n���v��ć���Y���T��L˚��������|�p�o���k� Wq����<��׬��n���.���  �  s�<TL�<z�<q��<E|�<�\�<��<���<���<H��<@�<2��<��<��<��<~�<�U�<��<pd�<��<��<��<X��<#t�<K�<�h�<&7�<�0z<�v<��z<,��<TH�<��<���<�d�<Z�<o�<�7�<BE�<��<2u<��j<7(i<�	p<T~<�m�< ��<���<Y֤<��<Q��<.S�<���<M�<�P�<ﱮ<1d�<�i�<��<5��<�ͭ<٭�< ��<��<B�<��<�M�<_o<�1^<�S<�>Q<�W<�`c<ws<,,�<���< �<
�<��z<��d<��K<\i3<��<��<�<_4<�Q"<K2<�6C<8xR<W^<8�d<B�f<�d<��_<��Y<�XS<k0M<��G<ϺB<�><��8<�1<�,(<�b<�<���;l	�;l�;��%;���:Ad:3�O: y�:=� ;�b<;ejq;�f�;�Շ;.�i;N^#;�2�:�L���F:�(�[�ĉY�q17�{����f�5
&9&�:��:�o;G�;�w�:ũ�:㵕:9xE:��9�Ɛ8si����]a��C��Yb��	A��f��{���6��>�*�#���3��E;��e:��2�x�$�I�X�
��������a��$&��<���S�g� s��Ov��p��8c�' Q���<��?)�X��lk�����Y�@� ����u�����Q�p�e��|��B��[	��b��4n/�,D�Z�{�n���~��
��Vn��*����cr���_�jtM��?��8���9�݋D���U�j]j��~�����kj���剼y<����z�Zg�S�l�@�w�1�1�'���!�d. �+� �#�"�P�$�H8&��)'�ʊ'�W�'��(��+�W�1���;�SK�`^��at�9\��{T���Y5���_��Po���y��e8��(\u�K�i���e���j�gyx��˅�K������pE���  �  N�<,K�<]�<͢<0Ī<Ҵ�<���<���<�e�<� �<p��<�Z�<���<��<a�<���<�`�<s��<ϳ�<c̽<��<���<S��<s7�<+�<d�<�c�<�?�<i|�<	h�<	��<��<��<J��<��<yH�<D��<��<�M�<?�<m6�<d�<��}<<9l�<=�<�Q�<kD�<���<y�<��<$��<�
�<��<�<~(�<�ݮ<���<�{�<��<{�<� �<yk�<��<���<��<`��<��<}:q<�'h<s�e<bVj<�Zt<c��<g��<�R�<c�<i_�<k�<�q<֎Z<e�D<�j3<m(<I�$<~�(<��1<
><�K<ȰV<�T_<�d<ye<�c<��^<x�Y<��S<=.N<�H<�C<�=<F�7<�z0<6'<��<<�M�;2t�;�?�;��k;��/;,�;��;�;��A;5-r;���;��;�;�+�;��M;���:�n:��7��'ӺC���

�;M��n����|���:��:���:.�:�S�:�v�:��:I�:b1T:���9> 9K�Y����@�t�����=g���;�&(���I���pӻ�����m��"��G&�$A&�t���M��	�| ����+�����	�ۈ���.���B�x�S�c^�v~a�"]��kR���C��x3�A�#��T��a�K��������R�L���Y�������ɉ��f�	S
��L�c���W*�\;�S\M�f:^�ͥk��ns��$t�7�m��<a��Q���A��Y5��B/��1��m:��I��\[�aXl�Uy�w ���Z���w�J!k�:z[�|+K��@<�tI0�(�i#��!���!�x�"�h�#�L:%�}K&�R5'��G(��*�$-��2�(};��H�X��Aj��|�����Č�=ʏ��(������Y��f�x�`j��7`�]���a��m��o~�mR���r������  �  �ˡ<3~�<��<�:�<o��<�'�<p��<5��<�F�<h��<���<��<�*�<$��<�o�<��<+��<<Y�<�<��<S��<Y��<M`�<�2�<G��<v��<o�<n��<�o�<F��<��<���<_0�<���<�߫<�<^%�<ǐ�<i�<�T�<rb�<	��<Ÿ�<Yy�<`�<[��<�e�<��<Z��<BL�<ǫ<�[�<-U�<��<6,�<�'�<��<sZ�<ω�<�f�<�۪<���<��<6r�<��<���<��<x�<U#�<�g<Bz}<-Z�<"�<#�<铍<c��<��<�(�<��<��~<��k<�NY<z$J<p@<��;<,�<<
B<	hI<�bQ<�xX<y�]<$`<�c`<��^<��[<{X<�S<�GN<yH<*B<�[;<�4<�,<��"<C?<pp<DO�;w?�;��;4ʛ;�p�;�l;Wqd;�xq;~�;�_�;6��;���;��;�w�;̡~;_J7;��:a:C�E��)�CD����j��b�9��`:b�:�A�:��:J��:��:��:7�:4TS:X��9ӈ�8����qF9�)͘�a|ۺ�i�H�B��y�����y��&�ݻ�R��:��2�����
��;�����=�h]�%8��S��2%��>�)/�;?=�F{F�B�I��lG�{k@��v6�&=+��J ���������
��:�����������K�52������s�
�}�����*���t'�j�3��@�J�L�tsV��\��L\�*W��:M���@��,4��T*�
�%��&'�"�.�	X;���I���W��Xb��h�(Gh��]c�k�Z�J�O�l�D��P:���1��+��(���%���$��+$�^$�4 %��f&��6(���*���-�ɪ1���6��G>��G���S��`��cn��jz�W����胼�\��a!���u��Ui���]�_�U�bnS�ЇW��ka��&o�N	~�h���*b���  �  s\�<� �<��<��<W��<�L�<%��<oֹ<I��<�M�<R�<�O�<�d�<?��<��<��<���<�P�<���<�߶<��<��<��<��<{�<�}�<x�<��<��<�z�<���<Kƥ<7U�<�8�<X�<%��<y:�<���<6��<�%�<���<`�<#�<Xj�<P�<틚<�d�<>�<Ӣ<��<��<q��<�Ԫ<Qx�<?��<�:�<���<9�<�4�<���<��< �<�N�<�X�<.��<GH�< p�<^͏<�ǌ<1ӊ<-W�<�v�<��<l�<��<��<�c�<��<,M�<'E�<H�|<��m<��`<m.W<ÇQ<}BO<�pO<�Q<�GS<NCU<*�V<�W<,�V<*mV<��U<Q�S<R�P<�L<��F<��><Z6<��,<�>#<;�<�h<�<q�;��;���;Y�;E��;�0�;��;Qd�;+ͬ; B�;|�;���;x�;^S�;;��;k�r; T5;M��:m�:�E:h%	:e�9��:��9:1~c:��:�Ռ:Ǳ�:4�:@�:k݃:9�h:7�3:�9�Տ��3��L�ֺʏ�E�7�+^�^B��߀��g-��"û�ջ�l仳Q��fﻔ뻪k�ڏػ\ѻYiл�	ػ$��^ ����fZ�6�&���.�z	3�aj3���0�R�,��('���!�O��7 ������������X����������N
�ܑ��L�~:��g�#��k)�hf0��~7���=���B���E���D�m�@�[A9��0���&����b��F�b$�o-��s8�6C���K�k�P�UR�7�P�M�H���B�\S=�s�8�3�4�P1��-��*��Z(���&�;�&�8h(���+�-�/�3#5�w�:�tO@�GF���L�tT���[��@c���i���n�S�p��jo��{j�.�b���Y�_�Q��L�P�J�n�M�P�U��`�|k���u��}��  �  ��<QW�<>�<I;�<꠲<�N�<V�<<�<%(�<�4�<iڸ<m��<��<���<O��<� �<A�<�]�<DX�<D��<>��<�E�< ��<��<Bʦ<J�<��<*?�<��<�s�<���<�~�<c�<�Ʋ<��<��<0E�<�Q�<%��<���<�7�<�k�<�j�<[�<5/�<���<�V�<@]�<,˜<oӝ<���<2�<�?�<�N�<�ª<��<�ث<!�<J0�<3��<�؟<��<���<D�<ʖ<bԕ<�<���<��<M�<~>�<m�<���<��<�\�<���<x��<��<���<��< ǅ<�K<�-t<��j<c<��\<sW<p�R<}�N<��K<	6I<��G<1H<cI<�)K<�XL<��K<�lH<>�A<d�8<IJ-</!<�d<<u<Q<�;�-�;���;f�;�C�;���;f��;�\�;���;���; ��;���;o,�;?��;u�;���;޺�;�u;i5G;+;��:Nh�:�۝:�t:�{6:)�:��9p�g9��C9�s9�v�9�<�9�5:<�9c�9������r��׺q���JJ�K�q��=��$j��}m�����ch��Ժ�����XŻ�ǻj ƻ�
û�׿�䢾�ɏ��U�ɻ��׻^n��L��
��=�����% ���#�H�&��@(��+)�%P)�z�(�kp&�E�"��z��5����;��	� Q	�t���O�Bi�� ��'�:
,�5}/�.�1��-3�~4�\f4��)4�H3�H�0��-�4�'���!�^��C��R�����G.���!��_)�#1��7���<�S�@�	C���D�	 F���F�ײF���E���C���?���:��5���/�I,�Y�*���,���1���8���@���H��JO��gT��
X���Z�Vp\�+�]��o^�v^��]�>O[�NuW�SR�	�L���G��`D�i�C�|F���K�'>S�<V[��c��wi��  �  ���<c��<��<K�<eW�</ �<)�< �<1!�<�ܬ<�ݰ<�Y�<�S�<QԻ<�)�<��<�<_��<;�<��<�~�<���<��<���<t1�<�Ԧ<J��<>��<3�<=�<ϧ�<�L�<�Ǵ<ߵ<fV�<3�<��<��<(ɰ<�8�<��<�Ҩ<��<��<�<l�<�	�<W�<j̓<�ܓ<|��<�>�<�̝<���<h�<k��<�b�<��<4��<vG�<�<f��<��<�<�s�<�#�<wv�<���<1J�<�#�<.y�<�c�<^��<fH�<X �<�I�<_��<��<uP�<:�<@�<T�</d�<��x<ˡn<t�c<��X<�!N< +D<J�;<�6<��3<ߑ4<<8<?=<��A<ٹC<��A<��:< z/<�!<:�<�<�o�;��;
�;��;*��;�Q�;���;n/�;��;^h�;��;q��;�)�;,��;���;S��;�H�;�ж;�1�;C��;�|;z<Z;��4;$�;���:�l:��9拹��8����Y���en�{k'�(©�J���n	��䄹M!I�^�Ⱥx< ���]�a���󄠻fѮ�/ٵ�X+���Ҵ������?����j��ך��o����Q��ĭ�����������$�̻=�ڻ�"껸���R]����r�ű�]�"�z�*�,�1��F7�r:�FO:�ay6�jV/�_&�yu�^����T5������'��D2�d�:�|@�y�A�M@��n<��$7�I1��+���&�:""��8���������������;��7�`��O#���(�co.���4���;�	C�J��2Q�MBV�s�X�t�W�GS�G�K���B��I:�w4�2�1��74�'";��3E���P�t[��Gc��h�5Qi���g��c�S�^�RaY��aT�sP�d]L�I� �E���B�1�@��r?���?�R�A��.E�`�I��#O�
�T��}Z��  �  ��<J��<n��<���<4L�<4x�<�L�<퇝<���<-�<��<��<�<�<���<3�<�߯<�֨<"w�<�<2Ӗ<�A�<�n�<�ޙ<�Ȟ<�Z�<@Щ<��<9%�<���<��<:��<pd�</�<Q�<��<3�<v?�<���<�a�<;�<dC�<�7�<��<]ݝ<P�<w�<-�<!<)�<�]�<[�<�0�<��<��<H�<t�<럠<W�<=ړ<��<�d�<o,�<��<7ȅ<�Љ<K�<_�<�O�<!0�<w��<�<��<Ew�<�;�<h|�<�F�<ۨ�<ӫ�<xS�<��<i��<-�<�r�<��s<I�d<8fT<��C<,@4<�'<$%<�	<	><��$<�-<+�4<��9<��8<�|1<.1$<Ҽ<���;H_�;���;k��;8X�;VL�;.��;P��;��;(��;A��;���;��;���;��;�u�;4T�;���;�[�;Ͻ;C�;!��;;HW~;�\R;��;���:�X:���M\��oU�)��=!�:"��h�KР�_�N����OL��m���w�N�]�ه���嵻��λ
ܻN8޻L׻��ɻ+,��,�������׾��[���e��j1���ע��Ū�����`=���PǻS�ѻd�ܻŢ軙�����T<����w�$�W�2�4�?���I�suP��Q�-M���C��B7�I)*��H���y+�щ���*���8��gF�wFQ��wW��X�M�S���J��@��R4�kX)��3 �i����Z�@m����/d�D��˴�W+��:����8��4`��&��/�/l:��XG�?�T���`�tXj��vo�t,o��ji�|P_�%�R�N�F�>�e�:���=�a}F�G�S���b�h-p�ATz�N^���~�]y��gp��e��Z�ӠP�z�H�=C�I�?�?�=���<�T�<�F)=�o>�&�?�N�A��D��bG�n�K�&FQ��  �  ���<mU�<��<2�<%��<;��<�	�<2��<ؒ<$w�<�x�<m]�<�j�<���<{��<�<��<��<}�<��< �<�e�<�p�<���<×<�ڟ<K��<爮<���<;̶<H]�<Ǹ<υ�<���<�Z�<�ն<�p�<��<Ƅ�<|�<f��<�#�<?�<��<�y�<hf�<���<��<{Xz<Hlx<=�}<���<[��<K��<�Q�<��<V�<��<��<�]�<�ӂ<�x<mp<T�o<�tv<�+�<���<-��<~�<#��<�g�<{�<B"�<��<x��<���<:�<K��<��<�:�<�<�<���<:�<]�<�t<la<O�K<=6<��!< �<�V<�<��<��<J�<g�'<��.<�)/<�x'<G_<�<ǰ�;5`�;Pp�;�+�;10z;Ǉ;̓�;^��;�K�;���;�8�;x<>�<��;��; �;!��;U}�;���;���;�!�;6 �;w�;�:�;�Q[;J;N��:ʝ�E��as%�a�]���|���~���f���<�����Ǻ�?���������΅F�����hG��%H�xO��y�����������]�˻ղ�[�������_Y���������Ꝼ�{��������/�Ż68λ�yֻ��߻ @�8����
������+��[>�CP���^�;�g���i�6d��>X�;�H�|08�3�*��"���"�ɩ*���8�ΰI���Z���g��To�Huo��h��#\�_fL�C�;�M�+�������L�&���:����+��x������Z�' �{w�����m�"�3�.�1>���O�`*b��s�������u����h�r�@#c��S���H�8D�W�G��^R�mb���t�֦��ʈ�]���[ˊ�W�������Np��A`���Q�!�F��-?��5;���9�0>:�,k;���<��7>�NU?�/S@���A���C�iG��M��  �  p��<G��<"��<6��<�k�<?Ȑ<���<6+�<(��<tD�<ړ�<�ܟ<��<fo�<��<)A�<��<]�<���<嫆<f��<%�}<J��<��<ܐ<��<ж�<�&�<�q�<-Z�<� �<]�<���<�Ƿ<;�<�W�<��<_�<��< 5�<�:�<�\�<�+�<=��<�d�<�Z�<Ӏ<&vp<��e<U�c<:j<L�w<��<@��<BN�<ا�<!��<��<C�<��<�Tt<�{d<w�[<*P[<o]c<Mr<�b�<�F�<�c�<:��<�v�<���<�ȣ<�Q�<��<o=�<���<o�<���<#G�<���<�M�<I��<
<�nq<�*[<[ B<;{(<��<�
�;���;���;�7�;�) <��<�r<T%<�q&<�w<��<R��;y�;�M�;��T;�N-;֧);�"G;�@};[K�;/��;��;�B�;��<�-<�� <���;L��;'4�;�[�;{��;2Z�;�;��;�A�;�È;��W;�;3gC:koK�7���Om�"��_��4姻/8��%�{�rh@�_$��j������&�i7r�Yʨ���ڻ�P�O��X��Z�\���p ��C߻�����٣��摻&ى�����M葻Wɜ��꨻I���ѱ��,�ƻ'�ͻԻ��ܻ2黊f���@A��3��^J���_��Iq�*|��F~�O�w��i�bW��QD��4���+���+��4�knD�8X��k�={�m
��2��ٕ{��Sl���X��>D���0�� �e��Q���H�/I����c���������j���]�ڎ�����#�,1���C��?Y�P�o����7É� 썼���Ja��&��q��W_��MR�V�L�w�P���\�{#o����񷋼�Ԓ�����锼#���������{��g���U�ͮG��m>�I�9��8���9�%�;�6�=��8?�L#@���@�3�@��4B��E��4L��  �  ���<L�<<ӭ<�t�<�'�<G��<��<b�</؁<
�<�?�<�x�<dx�<#E�<���<��<p,�<%��<�&�<*E�<ʍs<��o<�u<�܁<�ڋ<#�<+�<U��<>Ȳ<�5�<�3�<!g�<���<�p�<�o�<z׵<���<�۵<V�<}J�<08�<W��<0�<��<=.�<��<�`v<�^c<I�W<�fU<��\<�l<,�<dr�<*ޒ<Q��<2��<��<��<�[~<͞h<U2W<VpM<bM<�V<�f<:�{<�<�-�<�o�<���<a��<�У<�?�<��<�Ɯ<��<fd�<')�<��<��<�Q�<&\�<��<��n<�:V<~�:<��<E�<z��;�&�;2��;W �;W��;PS<|�<8�<Q[ <d6<��<S��;�!�;��k;�;/��:��:�a;PVR;��;g�;���;u��;;A<�B<C� <-��;���;\b�;tB�;���;�	�;���;��;�P�;ɳ�;@�P;@�:iK�9�ۦ��'@��܏�&���s�Ļ]tû�"��\8���fc���*����w��zS@������溻������ �@;(���%��	��X
�"���Ȼ6����`���=���/������o'������F��݁��pȻ:�λtԻ�Hܻo�����c-�JH"�|:��>S�Mk�YX~�+���;��y�����u�rca�K�L�]�;���1��1��A;��wL��b�S�w�ba��`������j��g�w�) b�6�J��85�G#��x��� �{N�K�C.����{��?���!�@Q��e����q9$�!�3�*�H�c�`��Jy�����o�������Ŕ��܏��f���oz��g�D�X�S�F�V�P�c�D�w�S=���ڑ�Q���3���囼����	�}tm�NY��}I���>�/�9��e8�-�9�H<��>�%;@�pA��"A�%!A��B�UiE���L��  �  �`�<\:�<���<:��<U>�<�>�<��<~�z<@�~<iՅ<�]�<C�<�/�<#�<}�<�ۦ<מ<`�<%1�<%|<��n<i�j<��p<�X<5�<r��<�0�<��<�u�<��<)�<�\�<X�<`I�<�=�<X��<���<��<Fܵ<MB�<�#�<���<���<ϝ<���<	A�<�Mr<E�^<ЯR<�XP<V�W<:�g<��|<(��< ��<nv�<�q�<F��<N��<��z<bzd<?|R<�dH<;	H<_PQ<+Yb<�x<��< P�<O�<A��<d��<jã<�,�<���<|��<���<r+�<7��<U�<��<�B�<�8�<�ˀ<�bm<ZST<j8<�<yu <��;��;�y�;���;���;V�<��<�d<�,<��<d<c��;�ɠ;�tZ;%O;;|�:(W�:�';(�B;т�;���;���;�;�� <:$<�� <�G�;��;V��;�i�;
�;p�;@�;�m�;s�;A��;R�M;��:�d�9Q㾺ŁO�O꘻�㼻1�λ�<ͻ���߽��z�o��*5�������qI�!;���K��5M��Kx��%�F-���*��`�r��s���̻����h�������J��L���rt�����������A���ɻ�ϻ$�ԻV\ܻ�\黴���$�-�#�Rl<�?�V��"o�B�����������:��y���d��kO�x�=��%4�
4��=��MO��{e��{�k����������ʆ���{�~e��rM��6�*I$�w���4��-��i�M�w��g6�������JT��g��x��&���$�5��kJ��2c�_�|����"���BD���(���e��ӿ}���i��5[�S2U�!Y�tof���z���������S��� d���c��?䎼�}��5�o�L�Z��NJ��[?���9�@v8�u�9��^<�v�>��@�lA��jA��HA��%B�̄E�i�L��  �  ���<L�<<ӭ<�t�<�'�<G��<��<b�</؁<
�<�?�<�x�<dx�<#E�<���<��<p,�<%��<�&�<*E�<ʍs<��o<�u<�܁<�ڋ<#�<+�<U��<>Ȳ<�5�<�3�<!g�<���<�p�<�o�<z׵<���<�۵<V�<}J�<08�<W��<0�<��<=.�<��<�`v<�^c<I�W<�fU<��\<�l<,�<dr�<*ޒ<Q��<2��<��<��<�[~<͞h<U2W<VpM<bM<�V<�f<:�{<�<�-�<�o�<���<a��<�У<�?�<��<�Ɯ<��<kd�<-)�<��<��<�Q�<0\�<��<�n<;V<��:<ʣ<^�<���;�&�;Z��;z �;u��;\S<��<=�<R[ <a6<��<?��;�!�;��k;̚;���:�:-a;�UR;䤏;6�;x��;J��;'A<xB<4� <��;���;Sb�;sB�;���;�	�;ƚ�; ��;�P�;;��P;�@�:bN�96ۦ�9'@�[܏���H�Ļ6tûo"��@8���fc���*�|��w���S@������溻1��"���� �U;(���%��	��X
�9"�'�Ȼf����`��!>���/�������'�����F�����pȻD�λ
tԻ�Hܻr�����c-�JH"�|:��>S�Mk�YX~�*���;��x�����u�rca�K�L�]�;���1��1��A;��wL��b�S�w�ba��`������j��g�w�) b�6�J��85�G#��x��� �{N�K�C.����{��?���!�@Q��e����q9$�!�3�*�H�c�`��Jy�����o�������Ŕ��܏��f���oz��g�D�X�S�F�V�P�c�D�w�S=���ڑ�Q���3���囼����	�}tm�NY��}I���>�/�9��e8�-�9�H<��>�%;@�pA��"A�%!A��B�UiE���L��  �  p��<G��<"��<6��<�k�<?Ȑ<���<6+�<(��<tD�<ړ�<�ܟ<��<fo�<��<)A�<��<]�<���<嫆<f��<%�}<J��<��<ܐ<��<ж�<�&�<�q�<-Z�<� �<]�<���<�Ƿ<;�<�W�<��<_�<��< 5�<�:�<�\�<�+�<=��<�d�<�Z�<Ӏ<&vp<��e<U�c<:j<L�w<��<@��<BN�<ا�<!��<��<C�<��<�Tt<�{d<w�[<*P[<o]c<Mr<�b�<�F�<�c�<;��<�v�<���<�ȣ<�Q�<��<u=�<���<x�<���<1G�<��<�M�<\��<<�nq<+[<� B<j{(<��<�
�;A��;���;�7�;�) <��<s<T%<�q&<�w<��<+��;F�;DM�;,�T;BN-;'�);"G;�?};�J�;���;'�;�B�;y�<�-<o� <���;.��;4�;�[�;���;JZ�;9�;��;
B�;Ĉ;b�W;��;jC:wlK�z��Om��!�����䧻�7����{�h@�%$�kj�����*�&��7r��ʨ���ڻ�P�t�����Z����+q �QD߻鰾�0ڣ��摻wى�֩���葻�ɜ�먻q���𱾻D�ƻ9�ͻԻ��ܻ2黍f���@A��3��^J���_��Iq�*|��F~�O�w��i�bW��QD��4���+���+��4�knD�8X��k�={�m
��2��ٕ{��Sl���X��>D���0�� �e��Q���H�/I����c���������j���]�ڎ�����#�,1���C��?Y�P�o����7É� 썼���Ja��&��q��W_��MR�V�L�w�P���\�{#o����񷋼�Ԓ�����锼#���������{��g���U�ͮG��m>�I�9��8���9�%�;�6�=��8?�L#@���@�3�@��4B��E��4L��  �  ���<mU�<��<2�<%��<;��<�	�<2��<ؒ<$w�<�x�<m]�<�j�<���<{��<�<��<��<}�<��< �<�e�<�p�<���<×<�ڟ<K��<爮<���<;̶<H]�<Ǹ<υ�<���<�Z�<�ն<�p�<��<Ƅ�<|�<f��<�#�<?�<��<�y�<gf�<���<��<{Xz<Hlx<=�}<���<[��<K��<�Q�<��<V�<��<��<�]�<�ӂ<�x<mp<T�o<�tv<�+�<���<-��<�<$��<�g�<}�<E"�<��<~��<���<E�<X��<��<�:�<�<�<���<V�<|�<$t<�a<��K<�6<��!<@�<W<�<)�<��<j�<~�'<��.<�)/<�x'<5_<�<���;�_�;�o�;�+�;9/z;�Ƈ;F��;ד�;K�;��;X8�;B<�<���;ހ�;��;	��;P}�;���;��;�!�;~ �;pw�;*;�;�R[;B ;V��:[|�,	��Zr%�e�]���|���~���f��<�z��S�Ǻ�?������#���F������G���H��O��Fy�!��!���B����˻�ղ�ݘ��z����Y��[��]���띻|��%�� ��R�ŻP8λ zֻ��߻(@�<����
������+��[>�CP���^�:�g���i�5d��>X�;�H�{08�3�*��"���"�ɩ*���8�ΰI���Z���g��To�Huo��h��#\�_fL�C�;�M�+�������L�&���:����+��x������Z�' �{w�����m�"�3�.�1>���O�`*b��s�������u����h�r�@#c��S���H�8D�W�G��^R�mb���t�֦��ʈ�]���[ˊ�W�������Np��A`���Q�!�F��-?��5;���9�0>:�,k;���<��7>�NU?�/S@���A���C�iG��M��  �  ��<J��<n��<���<4L�<4x�<�L�<퇝<���<-�<��<��<�<�<���<3�<�߯<�֨<"w�<�<2Ӗ<�A�<�n�<�ޙ<�Ȟ<�Z�<@Щ<��<9%�<���<��<:��<pd�</�<Q�<��<3�<v?�<���<�a�<;�<dC�<�7�<��<]ݝ<P�<w�<-�<!<)�<�]�<[�<�0�<��<��<H�<t�<럠<W�<=ړ<��<�d�<o,�<��<7ȅ<�Љ<K�<_�<�O�<"0�<x��<�<��<Kw�<�;�<r|�<�F�<먘<竕<�S�<8��<���<O�<	s�<>�s<��d<�fT<�C<~@4<;�'<m%<�	<D><ҝ$< -<G�4<�9<��8<�|1<1$<��<Y��;�^�;���;߬�;�W�;�K�;���;���;�;���;���;-��;I�;K��;H�;�u�;T�;���;�[�;<Ͻ;VC�;y��;[��;DX~;�]R;��;,��:�]:����Y��:T�	��9!�W!�Ug�'Ϡ�РN�4���OL�&n��)x�ݣ]�6���浻!�λ�ܻ�8޻�׻��ɻ�,������m���o������ f���1���ע��Ū�ڪ���=��Qǻt�ѻ{�ܻԢ転�����U<����w�$�W�2�3�?���I�suP��Q�-M���C��B7�H)*��H���y+�щ���*���8��gF�wFQ��wW��X�M�S���J��@��R4�kX)��3 �i����Z�@m����/d�D��˴�W+��:����8��4`��&��/�/l:��XG�?�T���`�tXj��vo�t,o��ji�|P_�%�R�N�F�>�e�:���=�a}F�G�S���b�h-p�ATz�N^���~�]y��gp��e��Z�ӠP�z�H�=C�I�?�?�=���<�T�<�F)=�o>�&�?�N�A��D��bG�n�K�&FQ��  �  ���<c��<��<K�<eW�</ �<)�< �<1!�<�ܬ<�ݰ<�Y�<�S�<QԻ<�)�<��<�<_��<;�<��<�~�<���<��<���<t1�<�Ԧ<J��<>��<3�<=�<ϧ�<�L�<�Ǵ<ߵ<fV�<3�<��<��<(ɰ<�8�<��<�Ҩ<��<��<�<l�<�	�<W�<j̓<�ܓ<|��<�>�<�̝<���<h�<k��<�b�<��<4��<vG�<�<e��<��<�<�s�<�#�<wv�<���<2J�<�#�</y�<�c�<b��<mH�<a �<J�<n��<��<�P�<U�<'@�<(T�<Vd�<D�x<"�n<��c<�X<1"N<[+D<��;<�6<ߢ3< �4<G<8<>?=<лA<�C<��A<��:<�y/<�!<	�<�<<o�;f��;e	�;A��;r��;Q�;��;�.�;5�;�g�;���;��;�)�;���;���;M��;�H�;�ж;=2�;���;�};�=Z;�4;w�;���:��l:R�9�ڋ���8��z��W���an�3h'����s����_	��䄹!"I�4�Ⱥ= ���]�߻������Ү��ٵ�,���Ӵ�����Ԓ��򢩻sk��u�������VR���ĭ����������U�̻a�ڻ�"�ʤ��W]�Ų�t�Ʊ�]�"�z�*�,�1��F7�r:�FO:�ay6�jV/�_&�yu�^����T5������'��D2�d�:�|@�y�A�M@��n<��$7�I1��+���&�:""��8���������������;��7�`��O#���(�co.���4���;�	C�J��2Q�MBV�s�X�t�W�GS�G�K���B��I:�w4�2�1��74�'";��3E���P�t[��Gc��h�5Qi���g��c�S�^�RaY��aT�sP�d]L�I� �E���B�1�@��r?���?�R�A��.E�`�I��#O�
�T��}Z��  �  ��<QW�<>�<I;�<꠲<�N�<V�<<�<%(�<�4�<iڸ<m��<��<���<O��<� �<A�<�]�<DX�<D��<>��<�E�< ��<��<Bʦ<J�<��<*?�<��<�s�<���<�~�<c�<�Ʋ<��<��<0E�<�Q�<%��<���<�7�<�k�<�j�<[�<5/�<���<�V�<@]�<,˜<oӝ<���<2�<�?�<�N�<�ª<��<�ث<!�<J0�<3��<�؟<��<���<D�<ʖ<bԕ< �<���<��<N�<>�<p�<���<��<�\�<
��<���<��<���<��< ǅ<FL<�-t<�j<cc<+�\<osW<��R<��N<�K<]6I<��G<tH<>cI<�)K<�XL<�K<�lH<4�A<L�8<#J-<�!<�d<�<�t<�;�;�,�;	��;��;�B�;��;���;�[�;��;��;ǰ�;i��;L,�;9��;��;.��;+��;�u;d6G;1,;���:k�:�ޝ:�t:��6:��:*ɭ91 h9n�C9's9�}�9�A�9�7:��9��9S�����r�2�׺G���KJ�v�q�*>���j��9n������&i���Ժ�n��XYŻ6ǻ� ƻxû/ؿ�E��������ɻ��׻�n��L��#
��=����% ���#�I�&��@(��+)�%P)�y�(�kp&�D�"��z��5����;��	� Q	�t���O�Bi�� ��'�:
,�5}/�.�1��-3�~4�\f4��)4�H3�H�0��-�4�'���!�^��C��R�����G.���!��_)�#1��7���<�S�@�	C���D�	 F���F�ײF���E���C���?���:��5���/�I,�Y�*���,���1���8���@���H��JO��gT��
X���Z�Vp\�+�]��o^�v^��]�>O[�NuW�SR�	�L���G��`D�i�C�|F���K�'>S�<V[��c��wi��  �  s\�<� �<��<��<W��<�L�<%��<oֹ<I��<�M�<R�<�O�<�d�<?��<��<��<���<�P�<���<�߶<��<��<��<��<{�<�}�<x�<��<��<�z�<���<Kƥ<7U�<�8�<X�<%��<y:�<���<6��<�%�<���<`�<#�<Xj�<P�<틚<�d�<>�<Ӣ<��<��<q��<�Ԫ<Qx�<?��<�:�<���<9�<�4�<���<��< �<�N�<�X�<.��<GH�< p�<_͏<�ǌ<2ӊ</W�<�v�<�<r�<��<*��<�c�<��<CM�<BE�<��|<ʜm<D�`<�.W<�Q<�BO<�pO<@Q<HS<�CU<{�V<W<m�V<amV<ʂU<o�S<c�P<�L<��F<��><66<Q�,<r>#<��<Ch<��<��;��;@��;��;���;0�;y��;�c�;�̬;�A�;?�;���;x�;tS�;l��;�r;�T5;3��:5o�:��E:�*	:��9��:`�9:Ѓc:���:،:
��:+�:��:�ރ:�h:�3:+�9�t5�>���ֺĐ�e�7�M,^�C������".���û��ջZm�]R�~g�$�*l�I�ػ�\ѻ�iл�	ػU��p ����oZ�<�&���.�|	3�bj3���0�R�,��('���!�O��6 ������������W����������N
�ܑ��L�~:��g�#��k)�hf0��~7���=���B���E���D�m�@�[A9��0���&����b��F�b$�o-��s8�6C���K�k�P�UR�7�P�M�H���B�\S=�s�8�3�4�P1��-��*��Z(���&�;�&�8h(���+�-�/�3#5�w�:�tO@�GF���L�tT���[��@c���i���n�S�p��jo��{j�.�b���Y�_�Q��L�P�J�n�M�P�U��`�|k���u��}��  �  �ˡ<3~�<��<�:�<o��<�'�<p��<5��<�F�<h��<���<��<�*�<$��<�o�<��<+��<<Y�<�<��<S��<Y��<M`�<�2�<G��<v��<o�<n��<�o�<F��<��<���<_0�<���<�߫<�<^%�<ǐ�<i�<�T�<rb�<	��<Ÿ�<Yy�<`�<[��<�e�<��<Z��<BL�<ǫ<�[�<-U�<��<6,�<�'�<��<sZ�<Ή�<�f�<�۪<���<��<6r�<��<���<��<x�<V#�<�g<Fz}<0Z�<&�<)�<�<m��<��<�(�<��<�~<�k<OY<�$J<�@<�;<~�<<q
B<\hI<�bQ< yX<]<D$`<d`<��^<��[<�X<��S<�GN<wyH<�)B<�[;<�4<�,<��"<�><$p<�N�;�>�;�;�ɛ;&p�;kl;Lpd;�wq;�;b_�;���;���;��;�w�;$�~;�J7;k��:�d:q�E�7)�]>D���uV��l�9��`:��:	D�:��:��:*�:�:��:�TS:f��9���8�����H9��Θ� ~ۺ�j�g�B�K�y�%��� ��ϒݻ�S�����2���#�
��;�G���>軮]�]8� T��B%��>�%)/�A?=�J{F�D�I��lG�|k@��v6�&=+��J ���������
��:�����������K�52������s�
�}�����*���t'�j�3��@�J�L�tsV��\��L\�*W��:M���@��,4��T*�
�%��&'�"�.�	X;���I���W��Xb��h�(Gh��]c�k�Z�J�O�l�D��P:���1��+��(���%���$��+$�^$�4 %��f&��6(���*���-�ɪ1���6��G>��G���S��`��cn��jz�W����胼�\��a!���u��Ui���]�_�U�bnS�ЇW��ka��&o�N	~�h���*b���  �  N�<,K�<]�<͢<0Ī<Ҵ�<���<���<�e�<� �<p��<�Z�<���<��<a�<���<�`�<s��<ϳ�<c̽<��<���<S��<s7�<+�<d�<�c�<�?�<i|�<	h�<	��<��<��<J��<��<yH�<D��<��<�M�<?�<m6�<d�<��}<<9l�<=�<�Q�<kD�<���<y�<��<$��<�
�<��<�<~(�<�ݮ<���<�{�<��<{�<� �<yk�<��<���<��<`��<��<~:q<�'h<v�e<gVj<�Zt<h��<m��<�R�<)c�<w_�<0k�<$q<�Z<��D<�j3<Em(<��$<��(<��1<P
><K<�V<�T_<d<�e<�c<��^<��Y<��S<?.N<�H<�C<ǜ=<#�7<�z0<�5'<x�<�<cM�;�s�;W?�;��k;��/;<�;��;V�;��A;�,r;���;��; �;�+�;>�M;���:q:	�7��%Ӻ]���	
�1KẴl���|��:���:|��:�/�:GU�:�w�:���:�I�:2T:���9� 9�Y�����t�-���h���;��(��J��sqӻU����m�#��G&�^A&�����M��	�� �;���Y���̦	�����.���B�|�S�!c^�x~a�#]��kR���C��x3�A�#��T��a�J��������R�K���Y�������ɉ��f�	S
��L�c���W*�\;�S\M�f:^�ͥk��ns��$t�7�m��<a��Q���A��Y5��B/��1��m:��I��\[�aXl�Uy�w ���Z���w�J!k�:z[�|+K��@<�tI0�(�i#��!���!�x�"�h�#�L:%�}K&�R5'��G(��*�$-��2�(};��H�X��Aj��|�����Č�=ʏ��(������Y��f�x�`j��7`�]���a��m��o~�mR���r������  �  s�<TL�<z�<q��<E|�<�\�<��<���<���<H��<@�<2��<��<��<��<~�<�U�<��<pd�<��<��<��<X��<#t�<K�<�h�<&7�<�0z<�v<��z<,��<TH�<��<���<�d�<Z�<o�<�7�<BE�<��<2u<��j<7(i<�	p<T~<�m�< ��<���<Y֤<��<Q��<.S�<���<M�<�P�<ﱮ<1d�<�i�<��<5��<�ͭ<٭�< ��<��<B�<��<�M�<_o<�1^<	�S<�>Q<�W<�`c<~s<1,�<���<(�<"
�<��z<��d<�K<�i3<��<�<2�<�4<�Q"<2K2<7C<exR<�^<^�d<c�f<"�d<��_<
�Y<�XS<m0M<��G<ĺB<�><��8<��1<�,(<�b<�<3��;	�;�;�%;{��:j>d:ɑO:�w�:�� ;?b<;%jq;�f�;�Շ;E�i;�^#;J3�:�I���rE:���[��Y��07�����f��&9��:^��:Up;ɿ;�x�:j��:S��:�xE:�9QÐ8vvi����&_a��D���b��
A�g��٠�����F>�Z�#��3��E;��e:��2���$�8I�q�
�������a��$&��<���S�
g�"s��Ov��p��8c�' Q���<��?)�X��kk�����Y�?� ����u�����Q�p�e��|��B��[	��b��4n/�,D�Z�{�n���~��
��Vn��*����cr���_�jtM��?��8���9�݋D���U�j]j��~�����kj���剼y<����z�Zg�S�l�@�w�1�1�'���!�d. �+� �#�"�P�$�H8&��)'�ʊ'�W�'��(��+�W�1���;�SK�`^��at�9\��{T���Y5���_��Po���y��e8��(\u�K�i���e���j�gyx��˅�K������pE���  �  �M�<�b�<�ь<�b�<���<۞�<�b�<*ݽ<���< ��<O�<U��<�L�<\&�<�_�<��<��<l�<x�<��<>��<(��<|Ǫ<�q�<�	�<��<ٗy<�-l<]�g<�7m<C {<E�<H`�<��<�E�<`ߟ<T��<US�<x��<q�z<B'h<�\<��Z<��b<�Er<���<�#�<*-�<�<2`�<m��<�h�<���<��<��<�5�<��<��<�c�<���<��<���<��<ş<f�<�$�<R{<r�c<o�P<��E<�2C<)�I<��W<)�i<{�z<aD�<	 �<��<�)t<��\<B�A<:�'<*q<ɩ<��<J	<A<#�)<C�<<��N<�\<3d<�f<#�d<��_<5WY<��R</L<��F<�
B<W�=<D�8<� 2<��'<��<�<��;���;�ZW;FH�:��%:.�i�@x��A�9�ĩ:�;��S;�-w;��w;��P;�S;��:�͏�i)�V7q�O]��zF����h��n'�������6���]:���:�� ;X4;=L�:_��:�h�:��5:;y�9�*57�㈹ߘ
�˩`��î�3D��I������û8����:��0�`�A���I�uH�lL>��3/���L��eQ����z�T.���F�Ni_��+t�j����M���~�Yo��Z�D�C�j�-�vV�ދ� ��2��� � ��8��p��O�}��~�������	�7��q ���3�K��pc��7z�I���$������"����}��i�NhU�'�E�'&>��@�zK��&^��|t�x���P������𐼮���A�$p�iY�C�D���3�>(��!�V ��� �3#�4s%��9'�X(�4(��(�w�(��y+���1�@Q=�N���c�|�_n���v��ć���Y���T��L˚��������|�p�o���k� Wq����<��׬��n���.���  �  g8�<
A�<��<�;�<]r�<�v�<�_�<��<`��<��<P�<�P�<eE�<���<��<���<H-�<��<-��<>��<���<���<,��<QU�<��<���<�z�<�<�<J��<��<��<�h�<[O�<?F�<g,�<�Q�<���<�k�<Ƹ<#�<�/�<4��<�<��<Ɇ�<��<	��<���<���<J^�<ig�<
��<h��<���<��<���<�s�<���<}��<}��<^��<�~�<e��<�Y�<��<�,�<���<_\�<VX�<hq�<�0�<���<K�<v��<��<�Ī<@�<�D�<Y��<䱚<é�<�݈<[��<��y<�.v<�Ax<.�~<ƿ�<�X�<�<<S�<y��<�%�<:�<�n�<�U�<�|<�8v<�.q<�m<�k<u�h<�ie<�(`<�W<jGL<�V=<�(,<�s<�1
<_��;q��;P��;6��;���;�<��<��<< <C8<�D�;���;��;��;��a;|�E;�QA;�R;R�q;R�;TA�;��;�ɲ;ٱ;��;]�;?\�;o?z;�r\;�D;�32;��%;�3;n�;[�;Xx�:�:1��9�@�ﺨ�>���}�����̣�縥�W����b�����f���^���k�����U|����»]��1������
�����i��5��k�ϻb���x��D�����Ϙ��J��.M��.ϫ�41��Bo��s}��CO��5~�����J���X��I����˻}Y廓�������q% �� ��.�P��K�?���-��0eܻ�{߻{��Wp�*'�Uj���'��-�O�,�K�&��������P�����ڻ:Iٻ�hݻ�们����󻺒����� Y��8 �����e��������A���/!��0�ޘ=���G�<�L�2L��F�!<�wj0���%���@��xf ��)��[6��D�WJQ��XZ��  �  ���<��<?,�<�]�<^W�<��<���<���<�*�<���<C�<��<ȓ�<2��<��<���<�w�<H�<6��<{��<^��<��<�7�<��<���<�<�׵<���<M$�<Uc�<��<�i�<�<~��<���<���<�1�<'�<\��<�
�<�}�<S�<f�<x�<̯<���<�ǻ<s~�<���<���<t��<N�<|��<���<}W�<�6�<��<�/�<��<��<���<��<W�<u��<���<��<w��<��<���<K�<���<��<>�<홤<<(^�<��<6Ш<A:�<�v�<韒<��<��<h�|<\y<��z<�<ݶ�<a�<֜�<��<Vَ<�N�<�d�<c��<p��<�}<��v<g�q<cIn<��k<�i<$�e<׋`<"�X<� M<��><.�-<��<��<Z0 <�|�;x�;ͫ�;=�;5Y<8�<6<<�\<@��;$(�;U�;��;�l;�YQ;V�L;K�\;ۄz;Uv�;Ԡ;�­;5�;���;���;
̝;�T�;¾|;e_;�.G;5;7(;�;um;� ;B�:�+�:�2�9��)��ߺ�)5��r�N����䝻01���ޘ��R����x��ya�Z�*Vg��#��փ������d{޻\���0�3�����fN�����J�̻JH��M�LF���e���#���|��@��V��L����ﯻq'��^;��a����c��/���ki���%����Ȼ�7� �� B�k��2�����>��O"���T�[+ڻ�;ݻ5A��� �?1�����$��%*�F�)�f$��z���2��P�sn��ٻs�ػ+�ܻ���α�O�����{��Q�����h��[��k��@���'�m���s�P�-��:��D���I�V_I���C���9��.�^$�oh�I{��=��)(�8�4�gB���N���W��  �  ���<���<4��<�x�<���<r��<���<���<W��<�<�<���<4)�<�a�<"��<��<���<%;�<V��<�[�<wM�<.�<Κ�<qq�<���<j��<p%�<���<gɵ<�@�<�@�<���<d@�<�c�<���<_I�<�^�<���<�3�<E�<L4�<-,�<��<ɇ�<�j�<�M�<q�<3��<��<���<y,�<���<6z�<�5�<���<C4�<�2�<���<��<��<מ�<�3�<��<���<v��<���<E�<Iq�<t�<���< �<M��<r��<ml�<.3�<�Ǫ<��<��<�I�<��<��<X�<QS�<���<�[�<ƚ�<�G�<G̃<�T�<���<qߍ<4h�<|M�<s��<�Ê<,�<X�<p]<�x<��s<��o<��l<�j<A�f<ea<%�Y<8CO<n�A<��2<��"<�<@<Ɗ <�i�;D�;��<*A<��<�I<�<~	<�u�;x��;�Һ;��;z�;�#r;9�l;��y;��;^
�;/��; �;���;VD�;�
�;؋�;�͐;ǩ�;+=g;FuO;z�<;'�.;y�";s;�+;���:���:e(�9��ٹU���f��i(T��*���O��ė�����£��f��R��]M��[���|�?2��������ѻ������I3��o����4���ػe�ûNE���(�������ݔ�ͩ��(���������� �����������Jq������栻�!���H��>����:ûi�ٻ��
^����������|
�p����B뻱�ۻ�&Ի]׻h)以���ߤ�.[��U���!��!��s�a���X	��m���'�yF޻��׻23׻'ۻ��6�����G󻨛��������ﻋT5������g`����P�'�?�3�Y�<���A�~lA��n<�&�3�o�)�Wx ��.�����6\$�S�/��v<�(�G��O��  �  "��<d��<�<���<���<{��<�<��<���<�b�<kE�<���<Jb�<�0�<�h�<��<�)�<*o�<S��<�o�<�i�<�@�<Z��<^?�<���<���<���<��<-?�<��<ň�<�l�<���<EN�<�g�<Rg�<.0�<�$�<0�<�ݺ<Ș�<��<��<��<u:�<�_�<3��<L��<���<݌�<��<��<���<wm�<�L�<�{�<}�<�/�<h��<��<mg�<%�<]��<�j�<G��<i��<"8�<*ή<�)�<��<���<��<a�<	 �<G��<Q�<���<�J�<�Z�<���<�T�<4.�<�B�<�C�<4u�<Z��<�Z�<�؊<(c�<L�<M�<?��<:��<���<#��<R8�<�ـ<N�{<�gv<r<�Xn<��j<�f<C�a<X�Z<�Q<��E<��8<i2+<�g<^�<�<�f	<�
<�<h<�b<~�<<��<�<�X�;;�;�}�;<�;��;4��;���;��;k��;l��;E̶;ܗ�;S��;g��;��;���;�ǅ;�}q;cdZ;��F;��6;�<(;=�;v�;%��: 5�:g�&:�Y���{�P��j�(��P�A8j�nJs�C�m���]��DK���=�e�;�(iJ��i��<���>���羻�@ԻJ-�+�TB��cػ�ɻ
g�����\���o���@���ە�����c��Ꞣ�;���𽦻���!'��W���R��ѕ��o𤻊.������ϻ@��6o����� 	�� 
���� �2�r)߻oһ��˻�λ*ڻ-�n ��z
�s�������,����
��4�<��%D��kۻ��ֻc�ֻ�ڻdl߻W&廔2�D������.�����)��;�������^
�����z�'�)��F1��5�l�5��1���*�U�"������4w�h��q����(�O�3�]=��D��  �  ٩�<�<���<.(�<-��<��<���<j��<w�<��<"�<��<�-�<�V�<r��<�.�<���<ۚ�<+P�<Z��<���<��<���<*�<K�<�Y�<w��<�F�<*�<�x�<�T�<�1�<�[�<��<1��<�u�<2��<3_�<aR�<�:�<pڼ<�Ǻ<�J�<PN�<z�<�P�<AN�<��<���<��<�h�<*�<��<l��<M;�<��<RV�<)(�<��<��< ��<eq�<v\�<9v�< ��<0	�<S��<�ݳ<�@�<h��<|<�<�I�<��<YN�<���<̶�<D�<�N�<K�<�-�<�ݝ<�×<R��<���<�<[��<��<G>�<Ub�<e�<T�<dގ<��<���<Ň<�Ԅ<��<,~<m�x<��s<�o<ݏj<��e<ݍ`<�.Z<�_R<�I<��><�3<�~)<̴ <�M<q�<>I<L�<�w<Vg<9G<�<m8<�M<��;���;c3�;2[�;���;�(�;ͧ;p��;���;#Q�;>��;#C�;�F�;k;�;��;eɔ;:�;�{;�d;8P;~�<;�X*;\;Er;�k�:��:��?:�� 9^"�ze����d�3�2�a>���>��7�yA-��*'��*�1h9�ĩU��"|��㓻�8�� ��>�ƻ\�˻Nʻ�=û;7���/��h#�������I���񖻥җ����@}��Sڞ�����̡��-���
�����v塻'Q������㭻$9���ŻggԻ���.ﻌ��2������'C��޻��ѻL�ǻ��û�;ƻ݆ϻ��ݻGg��.��7#�gW��d�æ��� �Ȇ���I��Ở�ۻ�ٻ�Sٻ��ۻ �޻�����廸�軺�껨F�H�K����"@�Z���"�Gh��������~��w$��'��`(���%�� ���������d�O-��!�y�)�`1�w�6��  �  �7�<��< ��<���<���<���<"��<k��<��<���<��<��<._�<��<~�<���<q��<���<z��<m��<ٹ�<Hh�<8��< ��<��<&.�<��<Zy�<+��<~��<e��<��<���<�g�<�I�<�<��<�A�<tW�<�h�<C��<�W�<ʼ�<��<���<%A�<k��<V��<B��<��<*[�<�z�<��<Ġ�<N��<v�<V�<��<���< �<*J�< d�<�W�<��<F�<G�<,��<#�<�ʵ<*�<4��<�]�<.��<�X�<س<K��<�l�<.گ<�<qJ�<�&�<�)�<�Ҙ<y�<7/�<�ˑ<��<m��<V�<[�<�>�<)��<���<�<q��<4Ƅ<m�<R�<x<z<�at<wXn<�Mh<`b<Ӈ\<I�V<bGP<�jI<�B<�~:<�23<��,<1m'<��#<�,"<8�!<��!<�!< �<�<��<6J<�~< ��;Z8�;<��;���;B��;�W�;2��;լ�;@�;$u�;��;S�;�Ӣ;��;�ؒ;�;�~�;�*l;��U;�>;��%;0�;���:jI�:��:�f+:�j[9�㊹�RC�����;Һ	$����
�)�����E��X������+���D��td�!���.<���^��rm���ұ������`J��~֨��Ƥ�)Ρ�I����-�����������F��;��������b�������{��y^���o��  ����������N_ɻƢѻX�ػmvݻ?�޻r$ܻ�ֻ��ͻ/�Żc����1��I����zƻ�л"�ܻ��Z�sQ��h�������������.軂q仙.��E��8����	�Ȳ�G��0��G軫;����.�)��$���aG �l[��,�-��ba�}��"��1���]�������ǉ��X�A=���6�����e �ȵ%��)��  �  ���<1��<.�<�s�<���<`<�<ǯ�<�N�<�>�<���<9�<�<B��<���<Ֆ�<Օ�<*�<S�<�#�<�Z�<?��<���<z�<���<��<a�<��<�]�<8�<*�<���<vd�<�A�<���<�7�<���<���<Q�<�}�<��<#
�<���<?��<�\�<}��<�{�<�<��<�i�<�Z�<(��<�Y�<�Q�<�W�<5&�<{�<�*�<2�<���<��<;�<=��<���<���<���<;Y�<�<�Һ<B�<��<��<Tk�<S�<��<3�<�ִ<�<��<bW�<��<$��<m��<���<�˚<�<ʙ�<(N�<��<C�<��<$��<ވ<^X�<��<���<���<u'�<��<�,z<�3s<�sk<�c<s�[<X%U<!YO<XhJ<YF</�A<��=<,�9<�5<�$2<��.<p,<��)<2�'<�X%<�"<֓<V�<~�<��<O<J�;-�;��;6q�;9��;��;���;զ�;X��;C�;���;�[�;2�;둌;�f�;�c�;V�m;2�T;d�7;#>;�)�:$�:��:'	):1��9��8�?P����]�?��r���Ԣ��ξ�.rպ���N7��
���|���$��y:�oNS�l8m���������;V��u���	w���"���1��w˪��������������̭�k󪻥馻�������u���b��#롻�u��|��`���������O����~»��ûd>Ż�ƻ�ǻw�Ȼ��ȻP�ǻ7�Ļ�������s��gṻM�������m6ǻa�λ��ջ��ۻ����㻘0�R軖k�Â��� |��r�y��ع黺������&�V0�g������	����(�HK����]	���
�����#��T��q�LE����������:�E���-�ǩ�t|�T��H�zJ�6����  �  �2�<���<���<�N�<A��<w��<���<���<���<A��<�c�<�K�<��<���<m��<+x�<`�<&�<O�<�`�<\|�<?��<��<�P�<j�<���<J��<�l�<���<9��<���<���<��<��<->�<��<�#�<�X�<�w�<���<���<���<g^�<���<=��<X��<��<㵿<�b�<u�<{h�<pտ<��<���<��<���<�Q�<3��<uy�<���<�ͼ<��<��<ډ�<�Ӹ<��<x��<<��<�"�<�6�<�Ȼ<��<]ѹ<�v�<a�<�<��<�q�<��<���<?��<���<L��<�i�<��<�~�<��<h��<�ǋ<,C�<_�<�T�<�7�<ځ<7ف<5��<��<�Q~<kMx<�p<R\f<�/\<��R<��J<��D<0�@<��><��=< I=<0�<<k;<�V9<�z6<�3<�J/<�G+<�&<p["<#K<��<J<.<<�F <0 �;;'�;>x�;B��;տ;�Ű;[�;��;���;� �;! �;���;�ց;XӀ;�Ny;B�g;��L;m�);�;��:��P:Jj�9T�i7`�H�B根�¹�ݹ0w�4  �#�K�:W���ꟺ~���c��������$�1}7�$cJ�y�\�Jn��;~�Pކ��̎�'q������b������˼�J�»��Ļ�»��T���k�ɷ���렻+���;���_��"_��!'ƻ|�λ��ӻ�+ջ�ӻ�λ��ȻBaûͷ������Ĺ�����������a���p���"��X��x��������pŻk&ɻ�ͻ*�ѻ!׻%*޻��V������
 ��}��%����{���C�����}�黳Z���뻎��FO��F���������{������#�Z������
�h&	�����	��Z	���	��*
�^�
�{���A����w�����5�q}��  �  ���<
��<�<�<�_�<�[�<���<���<d\�<�j�<���<t��<v��<Tx�<#�<\8�<��<Lg�<VS�<^�<bh�<~��<�<<��<o��<4�<7�<^��<��<��<M��<̥�<���<i�<�<�<A��<y��<��<	i�<~F�<v�<��<���<���<,[�<e�<�C�<���<2H�<��<�N�<� �<]�<��<��<8��<{��<��<'��<g�<Sc�<n�<�D�<|o�<}#�<p<�<NU�<T�<�t�<�w�<���<>��<�ݼ<PL�<Q>�<��<�t�<8��<@��< 4�<_�<l��<P5�<}�<J;�<$A�<l��<�$�<��<��<�d�<��}<pgy<�-x<)Xy<�{<��}<��}<�#{<�t<nRk<��_<S<�_G<��=<��7<y�4<��4<�l6<�(9<��;<i=<��<<o�:<��6<c2<�,<�&<]!<��<�d<�<5<_�<K�<8��;t��;���;���;G޷;�K�;z�;H[z;U�b;Q�V;��U;�^];�gg;��m;�yk;7�[;�?>;
�;t��:w,H:֝�8��!�H���j��Dd�B�D����q���Q�����=��(��E���ٺ�����n�*��;��?I�z�U��]a���m��|��X�����73������j�Ļ|aһ��ۻ��޻h�ۻ��һ6ƻ|������?����:��򾯻�����;̻ �ۻ���zI�Ӣ6���߻Ԣӻ��ǻ�������g����氻�Q�� ���#��zﺻ\V���
����������4�� L»(�Ļ��ɻ�
һŴݻ&������q�4���m��?�w���	���B���jn���D��P�����+���������!_�bh�1��p����%f�ؼ����}8����o��V
�v����	���P�<��Zx��v��V��  �  �@�<��<z��<�L�<+��<� �<4\�<���<���<=	�<l��<���<1��<���<..�<c8�<xT�<;�<o��<�F�<�?�<�C�<�Z�<�%�<��<(K�<<�<�F�<��<֩�<�3�<u�<D��<�^�<|S�<з�<���<���<v1�<�y�<�H�<G7�<$��<y�<���<���<��<UF�<2g�<=|�<뮱<���<&�<HL�<���<Y��<���<�*�<P �<��<��<��<���<d�<��<\>�<b(�<�<�c�<h}�<�)�<�u�<�<-�<FA�<Y�<R��<�:�<V,�<�[�<Ҙ�<���<�<���<r�<V$�<nt�<�l�<���<�x<I�o<t�k<8�k<x�n<,s<Lw<1y<c	w<�p<a�e<F,X<�|I<��;<��0<�*<��'<)<zF-<��2<8<��;<L=<��;<�;8<��2<�$,<U%<h�<�<�<��<Cb<K�<n�<;_�;���;r��;a��;�`�;}8�;�ln;�F;9�+;f|!;�b&;V�5;Z�H;�EW;�Z;(L;�0,;���:�҇:��9;�*��{��)�Ϻ�ٺҬǺWƣ��}s��d*����$���zW%��p�����+�ݺv	�� �n�3���B���M�5�U�\�]���g�H�w�[击|Y��D���=�»�@ػ�K껍@���-���x��G黤aػ��ƻw�����w����幻�*ʻ�޻'��e� �6������� ����w�ҳл���nǵ�p����-��l�����(?��(J»��ûa�ûAl»�����6��»R Ȼ2�һ1��1������q��+��������_����$a��T����+���ղ��,n�������"�'�)��Q-���,�}�'�3� ���A]���	��P�M���������������K�	�w����ld�|���<���  �  3��<B��<�]�<
�<ϊ�<��<���<˄�<t�<���<�^�<�q�<���<R��<t(�<���<T��<���<�\�<���<5f�<�B�<���<N�<���<�G�<�I�<8�<A��<��<��<g��<���<�Q�<{�<�g�<�h�<d��<��<�:�<�&�<|��<�:�<G��<�\�<H�<v�< ˮ<Jw�<���<F�<�ӯ<��<�#�<`j�<E��<Ǉ�<���<.�<!��<O�<V�<ͤ�<?h�<ل�<�o�<^�<�h�<N��<]��<>Ƚ<B�<�Z�<挸<V�<��<�;�<H۬<^ �<���<�<cZ�<أ<��<��<�<�<��<�^�<#_y<�l<z�c<��_<:�`<MOe<��k<�rq<�st<f�r<X?l<p�`<�Q<�A<Ƕ1<"�%<n%<��<�<�p$<�,<f�3<L9<s<<,�;<��7< 2<:�*<�i#<�W<'H<C�<��<� <�0<B�<:f�;�l�;�|�;��;�/�;�s};h<D;�8;n��:���:�I�:�R;~u-;M'B;5	I;xg<;\�;���::��й�*��g����5�l����rr��=�f�}d�&�	���(��s�'������,���9*���=�%�K�b+T���Y�7>_���h���y������F�����g$ѻO��g �������6��c����q��8ӻ�����D��HƸ��û�mֻ���&r���{��������Wj��x��HۻҞǻp��Ѱ�^���pp�����К���}û�ǻgɻ�Ȼ�yŻ�»�����»��ɻ��ֻ &���z������#���(���)��&%���T���!	���3��x��	����*.!���,��T5��Q9��A8���2�i�)�II�v��V���,���8����
��������cQ������	������j��  �  ?�<I��<f��<���<af�<b�<
z�<qd�<G�<1c�<�n�<H�<�
�<�(�<`��<�W�<$��<)�<�K�<�[�<�h�< �<q��<�{�<��<I��<d��<�3�<)	�<��<��<�<�<�U�<�{�<T�<�g�<���<�1�<� �<���<���<�q�<�j�<��<�b�<�d�<5��<��<L[�<am�<EJ�<L��<�$�<��<⨼<�6�<v�<�<�ʶ<aL�< ϩ<���<���<�E�<u��<� �<&��<eS�<SJ�<���<!9�<�ټ<��<���<!��<U.�</�<�ѫ<D�<�ɨ<<��<�i�<f}�<W�<	��<T>�<}h�<�7r<�d<)w[<c�W<_Y<	�^<e�f<�^m<? q<h�o<�%i<��\<h�L<Qh;<��*<~�<�<��<;
<s<�'<e�/<<�6<\�:<A�:<�I7<�F1<G�)<~�!<#r<G=<&�<�?<"�	<I<�<��;���;���;��;fG�;�'d;�s&;�]�:�ȴ:tѧ:z_�:��:�;H3;��<;W�0;��;gŮ:�N�9�H�����Z�P�7�ӫ9��1(���	�lͺ�\����>�>R�b4�<�}����N-�`���1���E���R���Y�0�]�8b��1k��^}�׍��t�� ^��<�ۻA(�� ���(��'�{�L�d���ۻ��Ȼ�Y���ξ�cʻ��޻x��u���� ��0������=
�����X���+ͻ<~���ⲻC*��z�P��3o���ǻ�~˻@�̻'{˻ ȻYoĻ�c»�4Ļ�˻;�ڻA�|����!��t+�9B1�l�1��v,��5#�`���-�#m��~��:�L�gF���&�=�3�Q=���A�h@�+:�j40��Z$�<��u�����>��=���i�3��8������"8��i�y��8w�:��D��  �  ��<�,�<���<��<A�<��<��<��<䷻<�&�<|e�<�>�<^�<f��<K�<<��<3��<�<�<�6�<x�<���<��<�/�<�.�<"Խ<�!�<>�<���<���<��<��<|�<��<�*�<���<8�<�(�<���<���<��<���<�9�<��<��<⤽<g�<�]�<���<��<���<p�<LV�<�,�<�,�<��<@��<qu�<�h�<��<�Y�<&��<_=�<��<5˟<�4�<���<���<鋲<,��<�X�<���<r��<���<"ķ<�I�<�Ӱ<Sʭ<n�<���<&��<�W�<N¥<�7�<'9�<(~�<��<�g�<0S�<@�o<��a<�|X<��T<��V<U�\<p�d<C�k<n�o<@�n<6h<��[<�[K<�d9<�y(<�<=<F�<�X<K�<�/%<��.<6<�:<�L:<��6<5�0<P)<)B!<U�<y<^�<p�<E	<�<Yz<F��;�b�;��;�S�;���;w�Z;�;��:�.�:j��:y��:j-�:��;��-;�8;�s,;�a	;I��:�R9i�j�
���*�ދC��E��x2��~�spں�ꕺ�dK�k^$���9��W��ӓ��D���b����4��H�CU�S�[��T_��]c��sl�
��%��5x���M��E�߻. ��k�
���V�Z+�^��B��r߻�e˻����,	����̻����@��A����?�������
��N ���YPϻ"轻.ͳ�ٰ�ʝ��������fȻ��̻�iλ��̻(ɻ.9Ż?ûq�Ļ�̻�0ܻݗ��"������#�gN.�g64� k4�g/��k%�������i��ܙ��^�5��	����(�6���?��|D��SC���<�r�2�:&����������<�a@����������M�q�i�����X�`��э�����  �  ?�<I��<f��<���<af�<b�<
z�<qd�<G�<1c�<�n�<H�<�
�<�(�<`��<�W�<$��<)�<�K�<�[�<�h�< �<q��<�{�<��<I��<d��<�3�<)	�<��<��<�<�<�U�<�{�<T�<�g�<���<�1�<� �<���<���<�q�<�j�<��<�b�<�d�<5��<��<L[�<am�<EJ�<L��<�$�<��<⨼<�6�<v�<�<�ʶ<aL�< ϩ<���<���<�E�<u��<� �<&��<eS�<SJ�<���<!9�<�ټ<��<���<#��<W.�</�<�ѫ<I�<�ɨ<�<��<�i�<o}�<a�<��<^>�<�h�<�7r<�d<;w[<s�W<_Y<�^<n�f<�^m<C q<i�o<�%i<��\<`�L<Gh;<��*<o�<��<��<(
<`<�'<R�/<*�6<J�:<2�:<�I7<�F1<>�)<x�!<r<G=<(�<�?<*�	<I<�<��;��;���;�;�G�;�'d;�s&;�^�:�ɴ:�ѧ:�_�:C��:*�;H3;��<;X�0;��;7Ů:�M�9��H�^��[���7��9��1(���	�ͺ@]����>�cS�s4�5�}�}����-��`�Ҷ1�ưE��R���Y�<�]�@b��1k��^}�׍��t�� ^��<�ۻA(�� ���(��'�{�L�d���ۻ��Ȼ�Y���ξ�cʻ��޻x��u���� ��0������=
�����X���+ͻ<~���ⲻC*��z�P��3o���ǻ�~˻@�̻'{˻ ȻYoĻ�c»�4Ļ�˻;�ڻA�|����!��t+�9B1�l�1��v,��5#�`���-�#m��~��:�L�gF���&�=�3�Q=���A�h@�+:�j40��Z$�<��u�����>��=���i�3��8������"8��i�y��8w�:��D��  �  3��<B��<�]�<
�<ϊ�<��<���<˄�<t�<���<�^�<�q�<���<R��<t(�<���<T��<���<�\�<���<5f�<�B�<���<N�<���<�G�<�I�<8�<A��<��<��<g��<���<�Q�<{�<�g�<�h�<d��<��<�:�<�&�<|��<�:�<G��<�\�<H�<v�< ˮ<Jw�<���<F�<�ӯ<��<�#�<`j�<E��<Ǉ�<���<.�<!��<N�<V�<ͤ�<?h�<ل�<�o�<^�<�h�<N��<]��<?Ƚ<B�<�Z�<錸<V�<��<�;�<P۬<h �<���<�<qZ�<أ<��<��<�<�<��<�^�<H_y<*�l<��c<�_<U�`<dOe<��k<�rq<�st<h�r<T?l<f�`<ٌQ<�A<��1<�%<N%<��<��<�p$<�,<A�3<[L9<Q<<�;<��7<�2<(�*<�i#<�W<&H<H�<��<� <�0<[�<tf�;�l�;}�;��;�/�;6t};�<D;9;y��:���:tJ�:S;�u-;|'B;M	I;yg<;E�;8��:�:��йz+��Y���t6�������s�O򨺤�f��f�\�	�ɡ(�Ȟs�����=��{��:*���=�N�K��+T���Y�F>_���h���y������F�����g$ѻO��g �������6��c����q��8ӻ�����D��HƸ��û�mֻ���%r���{��������Wj��x��HۻҞǻp��Ѱ�^���pp�����К���}û�ǻgɻ�Ȼ�yŻ�»�����»��ɻ��ֻ &���z������#���(���)��&%���T���!	���3��x��	����*.!���,��T5��Q9��A8���2�i�)�II�v��V���,���8����
��������cQ������	������j��  �  �@�<��<z��<�L�<+��<� �<4\�<���<���<=	�<l��<���<1��<���<..�<c8�<xT�<;�<o��<�F�<�?�<�C�<�Z�<�%�<��<(K�<<�<�F�<��<֩�<�3�<u�<D��<�^�<|S�<з�<���<���<v1�<�y�<�H�<G7�<$��<y�<���<���<��<UF�<2g�<=|�<뮱<���<&�<HL�<���<Y��<���<�*�<P �<��<��<��<���<d�<��<\>�<b(�<�<�c�<i}�<�)�<�u�<���<1�<KA�<"Y�<[��<�:�<c,�<�[�<䘨<���<�<���<��<q$�<�t�<m�<���<x<y�o<��k<^�k<��n<3,s<'Lw<<y<f	w<�p<S�e<0,X<�|I<��;<a�0<�*<��'<�)<DF-<L�2<�8<{�;<�K=<l�;<�;8<f�2<�$,<U%<^�<�<�<��<Yb<h�<��<�_�;D��;֗�;���;a�;�8�;�mn;PF;��+;}!;Jc&;��5;��H;�EW;�Z;(L;�0,;%��:�ч:8�9�+�<}����Ϻ��ٺ~�Ǻȣ��s�h*�����f���dZ%�=p�篨�3�ݺ�	�E� ���3�׿B�'�M�U�U�q�]���g�P�w�^击~Y��D���=�»�@ػ�K껌@���-���x��G黤aػ��ƻw�����v����幻�*ʻ�޻'��d� �6������� ����w�ҳл���nǵ�p����-��l�����(?��'J»��ûa�ûAl»�����6��»R Ȼ2�һ1��1������q��+��������_����$a��T����+���ղ��,n�������"�'�)��Q-���,�}�'�3� ���A]���	��P�M���������������K�	�w����ld�|���<���  �  ���<
��<�<�<�_�<�[�<���<���<d\�<�j�<���<t��<v��<Tx�<#�<\8�<��<Lg�<VS�<^�<bh�<~��<�<<��<o��<4�<7�<^��<��<��<M��<̥�<���<i�<�<�<A��<y��<��<	i�<~F�<v�<��<���<���<,[�<e�<�C�<���<2H�<��<�N�<� �<]�<��<��<8��<{��<��<'��<g�<Sc�<n�<�D�<|o�<}#�<p<�<NU�<T�<�t�<�w�<���<?��<�ݼ<SL�<V>�<��<�t�<D��<N��<04�<s�<���<i5�<'}�<h;�<DA�<���<�$�<$��<��<�d�<��}<�gy<�-x<QXy<<�{<ɵ}<��}<�#{<�t<]Rk<��_<�S<�_G<��=<L�7<<�4<V�4<ul6<P(9<h�;<*=<��<<:�:<e�6<<2<Ì,<�&<Q!<��<�d<&�<P<��<v�<���;���;P��; ��;�޷;L�;��;@\z;<�b;#�V;Q�U;_];(hg;�m;�yk;9�[;�?>;��;���:*H:&��8#���H���j�Id�x�D�&��͏��h����u�=�7*���F��ٺ���a��ʋ*�E;�@I���U��]a���m�'�|��X�����83������j�Ļ{aһ��ۻ��޻h�ۻ��һ6ƻ|������?����:��򾯻�����;̻ �ۻ���zI�Ӣ6���߻Ԣӻ��ǻ�������g����氻�Q�� ���#��zﺻ\V���
����������4�� L»(�Ļ��ɻ�
һŴݻ&������q�4���m��?�w���	���B���jn���D��P�����+���������!_�bh�1��p����%f�ؼ����}8����o��V
�v����	���P�<��Zx��v��V��  �  �2�<���<���<�N�<A��<w��<���<���<���<A��<�c�<�K�<��<���<m��<+x�<`�<&�<O�<�`�<\|�<?��<��<�P�<j�<���<J��<�l�<���<9��<���<���<��<��<->�<��<�#�<�X�<�w�<���<���<���<g^�<���<=��<X��<��<㵿<�b�<u�<{h�<pտ<��<���<��<���<�Q�<3��<uy�<���<�ͼ<��<��<ډ�<�Ӹ<��<x��<<��<�"�<�6�<�Ȼ<��<aѹ<w�<h�<�<��<�q�<0��<���<X��<���<k��<�i�<�<�<2��<���<ȋ<OC�<1_�<U�<�7�<5ځ<Hف<B��<�<�Q~<cMx<qp<4\f<�/\<\�R<y�J<��D<��@<��><��=<�H=<�<<�j;<�V9<]z6<�3<�J/<aG+<�&<c["< K<��<^<L<E<�F <� �;�'�;�x�;Ѣ�;�տ;[ư;�[�;���; ��;!�;� �;�;2ׁ;�Ӏ;�Ny;C�g;��L;�);q�;|�:��P:c�9��h7��H�jM�¹�ݹ�{�� �l�K�8Y���쟺���ͬ�l�s���$��}7�acJ���\�in��;~�Vކ��̎�)q������b������˼�I�»��Ļ�»��S���k�ɷ���렻+���;���_��"_��!'ƻ|�λ��ӻ�+ջ�ӻ�λ��ȻBaûͷ������Ĺ�����������a���p���"��X��x��������pŻk&ɻ�ͻ*�ѻ!׻%*޻��V������
 ��}��%����{���C�����}�黳Z���뻎��FO��F���������{������#�Z������
�h&	�����	��Z	���	��*
�^�
�{���A����w�����5�q}��  �  ���<1��<.�<�s�<���<`<�<ǯ�<�N�<�>�<���<9�<�<B��<���<Ֆ�<Օ�<*�<S�<�#�<�Z�<?��<���<z�<���<��<a�<��<�]�<8�<*�<���<vd�<�A�<���<�7�<���<���<Q�<�}�<��<#
�<���<?��<�\�<}��<�{�<�<��<�i�<�Z�<(��<�Y�<�Q�<�W�<5&�<{�<�*�<2�<���<��<;�<=��<���<���<���<;Y�<�<�Һ<C�<	��<��<Wk�<W�<���<;�<�ִ<"�<'��<uW�<3��<>��<���<���<�˚<:�<<ON�<�<h�<<��<E��<#ވ<yX�<��<���<���<}'�<��<�,z<�3s<�sk<�c<A�[<%U<�XO<hJ<F<��A<m�=<��9<��5<u$2<G�.<:,<��)<�'<�X%<�"<ԓ<_�<��<��<y<lJ�;�-�;7�;�q�;���;���;.��;j��;罨;�C�;���;e\�;��;.��;$g�;d�;X�m;�T;�7;�=;a(�:��:�}�:�):-�9�8�RP�R��4�?�/u��ע��о�tպ����8�����P}�\�$��y:��NS��8m���������BV��y���w���"���1��w˪��������������̭�k󪻥馻������u���b��#롻�u��|��`���������O����~»��ûd>Ż�ƻ�ǻw�Ȼ��ȻP�ǻ7�Ļ�������s��gṻM�������m6ǻa�λ��ջ��ۻ����㻘0�R軖k�Â��� |��r�y��ع黺������&�V0�g������	����(�HK����]	���
�����#��T��q�LE����������:�E���-�ǩ�t|�T��H�zJ�6����  �  �7�<��< ��<���<���<���<"��<k��<��<���<��<��<._�<��<~�<���<q��<���<z��<m��<ٹ�<Hh�<8��< ��<��<&.�<��<Zy�<+��<~��<e��<��<���<�g�<�I�<�<��<�A�<tW�<�h�<C��<�W�<ʼ�<��<���<%A�<k��<V��<B��<��<*[�<�z�<��<Ġ�<N��<v�<V�<��<���< �<*J�< d�<�W�<��<F�<G�<,��<#�<�ʵ<+�<6��<�]�<2��<�X�<�س<U��<�l�<>گ<#�<�J�<�&�<�)�<Ә<%y�<Z/�<�ˑ<��<���<{�<5[�<?�<G��<���<%�<���<@Ƅ<"m�<V�<p<z<�at<ZXn<tMh<�_b<��\<
�V<GP<VjI<�B<9~:<n23<:�,<�l'<��#<�,"<�!<��!<��!<��<�<�<JJ<<O��;�8�;���;G��;���;X�;Ũ�;h��;�@�;�u�;e�;��;�Ӣ;��;#ْ;L�;�~�;�*l;r�U;�>;�%;��;���:�G�:��:9b+:aX[9>특�WC�󡝺Y=Һ/&����
�����������|��}�+�D�D�ud�8���><���^��ym���ұ������aJ��~֨��Ƥ�)Ρ�I����,�����������F��;��������b�������{��y^���o��  ����������N_ɻƢѻX�ػmvݻ?�޻r$ܻ�ֻ��ͻ/�Żc����1��I����zƻ�л"�ܻ��Z�sQ��h�������������.軂q仙.��E��8����	�Ȳ�G��0��G軫;����.�)��$���aG �l[��,�-��ba�}��"��1���]�������ǉ��X�A=���6�����e �ȵ%��)��  �  ٩�<�<���<.(�<-��<��<���<j��<w�<��<"�<��<�-�<�V�<r��<�.�<���<ۚ�<+P�<Z��<���<��<���<*�<K�<�Y�<w��<�F�<*�<�x�<�T�<�1�<�[�<��<1��<�u�<2��<3_�<aR�<�:�<pڼ<�Ǻ<�J�<PN�<z�<�P�<AN�<��<���<��<�h�<*�<��<l��<M;�<��<RV�<)(�<��<��< ��<eq�<v\�<9v�<��<0	�<S��<�ݳ<�@�<i��<~<�<�I�<��<^N�<���<Զ�<O�<�N�<\�<�-�<�ݝ<ė<n��<���<=�<|��<��<i>�<vb�<��<q�<ގ<��<���< Ň<�Ԅ<��</~<f�x<��s<�o<��j<a�e<��`<�.Z<i_R<�I<��><��3<F~)<�� <�M<;�<I<$�<�w<@g<-G<�<t8<�M<J��;���;�3�;�[�;F��;r)�;�ͧ;���;	��;�Q�;���;�C�;	G�;�;�;C�;�ɔ;a�;#{;�d;�7P;1�<;SX*;�;�q;�i�:��:��?:3� 9�&��g��&��e�*�2��a>�y�>��7�B-��+'�G*��h9��U��"|��㓻�8��
��D�ƻ`�˻Pʻ�=û<7���/��h#�������I���񖻤җ����@}��Rڞ�����̡��-���
�����v塻'Q������㭻$9���ŻggԻ���.ﻌ��2������'C��޻��ѻL�ǻ��û�;ƻ݆ϻ��ݻGg��.��7#�gW��d�æ��� �Ȇ���I��Ở�ۻ�ٻ�Sٻ��ۻ �޻�����廸�軺�껨F�H�K����"@�Z���"�Gh��������~��w$��'��`(���%�� ���������d�O-��!�y�)�`1�w�6��  �  "��<d��<�<���<���<{��<�<��<���<�b�<kE�<���<Jb�<�0�<�h�<��<�)�<*o�<S��<�o�<�i�<�@�<Z��<^?�<���<���<���<��<-?�<��<ň�<�l�<���<EN�<�g�<Rg�<.0�<�$�<0�<�ݺ<Ș�<��<��<��<u:�<�_�<3��<L��<���<݌�<��<��<���<wm�<�L�<�{�<}�<�/�<h��<��<mg�<%�<]��<�j�<G��<i��<#8�<*ή<�)�<��<���<��<d�< �<L��<Q�<���<�J�<[�<ѻ�<�T�<I.�<�B�<�C�<Nu�<u��<[�<�؊<Bc�<&L�<e�<U��<M��<���</��<[8�<�ـ<Q�{<�gv<r<�Xn<��j<��f<�a<*�Z<ډQ<L�E<��8<32+<�g<+�<�<Yf	<�
<�<�g<}b<t�< <��< �<�X�;v�;<~�;��;�;���;&��;x��;ֵ�;���;�̶;9��;���;���;8�;���;�ǅ;!~q;ddZ;o�F;^�6;p<(;��;��;���:�3�:;�&:Qt��a�{���E�(���P�9j�*Ks��m�,�]�JEK�o�=���;�tiJ�M�i�=���>���羻�@ԻO-�.�VB��cػ�ɻ
g�����\���o���@���ە�����c��Ꞣ�;���𽦻���!'��W���R��ѕ��o𤻊.������ϻ@��6o����� 	�� 
���� �2�r)߻oһ��˻�λ*ڻ-�n ��z
�s�������,����
��4�<��%D��kۻ��ֻc�ֻ�ڻdl߻W&廔2�D������.�����)��;�������^
�����z�'�)��F1��5�l�5��1���*�U�"������4w�h��q����(�O�3�]=��D��  �  ���<���<4��<�x�<���<r��<���<���<W��<�<�<���<4)�<�a�<"��<��<���<%;�<V��<�[�<wM�<.�<Κ�<qq�<���<j��<p%�<���<gɵ<�@�<�@�<���<d@�<�c�<���<_I�<�^�<���<�3�<E�<L4�<-,�<��<ɇ�<�j�<�M�<q�<3��<��<���<y,�<���<6z�<�5�<���<C4�<�2�<���<��<��<מ�<�3�<��<���<v��<���<E�<Iq�<t�<���< �<N��<s��<ol�<13�<�Ǫ<��<��<�I�<��<&��<X�<`S�<���< \�<ٚ�<�G�<[̃<U�<���<�ߍ<Eh�<�M�<���<�Ê<,�<X�<w]<
�x<��s<��o<��l<�j<(�f<�da<�Y<CO<I�A<��2<_�"<�<�?<�� <�i�;�;��<A<��<�I<�<!~	<�u�;���;�Һ;��;��;$r;��l;c�y;]��;�
�;y��;J �;щ�;�D�;�
�;��;�͐;ݩ�;C=g;GuO;d�<;��.;7�";;�+;���:���:�#�9��ٹ������)T�H+���O�����)��/��f�1�R��]M��[�Ҭ|�O2��ʆ���ѻ������L3��p����4���ػe�ûNE���(������ݔ�ͩ��(���������� �����������Iq������栻�!���H��>����:ûi�ٻ��
^����������|
�p����B뻱�ۻ�&Ի]׻h)以���ߤ�.[��U���!��!��s�a���X	��m���'�yF޻��׻23׻'ۻ��6�����G󻨛��������ﻋT5������g`����P�'�?�3�Y�<���A�~lA��n<�&�3�o�)�Wx ��.�����6\$�S�/��v<�(�G��O��  �  ���<��<?,�<�]�<^W�<��<���<���<�*�<���<C�<��<ȓ�<2��<��<���<�w�<H�<6��<{��<^��<��<�7�<��<���<�<�׵<���<M$�<Uc�<��<�i�<�<~��<���<���<�1�<'�<\��<�
�<�}�<S�<f�<x�<̯<���<�ǻ<s~�<���<���<t��<N�<|��<���<}W�<�6�<��<�/�<��<��<���<��<V�<u��<���<��<w��<��<���<K�<���<��<>�<<�<+^�<��<:Ш<G:�<�v�<�<��<��<z�|<oy<��z<���<綄<j�<ߜ�<��<^َ<�N�<�d�<g��<t��<�}<��v<e�q<^In<}�k<�i<�e<ȋ`<�X<� M<��><�-<��<��<G0 <�|�;�w�;���;�<�;,Y<1�<2<<�\<K��;4(�;k�;��;D�l;(ZQ;��L;��\;)�z;}v�;:Ԡ;�­;X�;ʜ�;͢�; ̝;U�;پ|;&e_;�.G;5;�6(;�;Hm;� ;� �:+�:0�9��)���ߺ)*5�B�r�t����䝻R1���ޘ�
S��"�x�za�4Z�FVg��#��߃�����h{޻_���1�3�����fN�����K�̻JH��M�LF���e���#���|��@��V��L����ﯻq'��^;��a����c��/���ki���%����Ȼ�7� �� B�k��2�����>��O"���T�[+ڻ�;ݻ5A��� �?1�����$��%*�F�)�f$��z���2��P�sn��ٻs�ػ+�ܻ���α�O�����{��Q�����h��[��k��@���'�m���s�P�-��:��D���I�V_I���C���9��.�^$�oh�I{��=��)(�8�4�gB���N���W��  �  ��<��<���<!��<H��<'��<���<T:�<-��<�,�<1��<x�<�/�<^v�<��<Aq�<"�<QD�<���<?o�<���<ڟ�<�m�<��<?��<���<Q��<]2�<��<Y�<�t�<Wf�<#��<M�<��<���<���<���<Dw�<H�<f��<�<\�<�
�<Tb�<l��<���<���</L�<��<a�<
��<�Z�<Y�<P/�<���<�v�<���<���<aG�<1��<�g�<6F�<���<�I�<'��<H�<ȏ�<���<��<瘻<M��<~�<g�<���<U��<���<�m�<3,�<$��<�Z�<}J�<�'�<3�<���<�*�<���<tt�<�נ<4��<=�<�<�<�G�<�p�<� �<j̏<Z݋<���<�6�<���<Ҥ�<7��<6)�<�ˀ<�	}<d4v<ym<�-b<�V<(�K<�_B<w�;<S�8</=8<�":<��<<�?<?<w<<�j5<9�+<��<�|<	<���;)�;�@�;�J�;~e�;,�;�b�;/� <Z��;36�;�C�;h=�;9��;��;9�;�i�;���;a��;�E�;���;7ǃ;�Lz;o�d;�E;�;�[�:y�:;��9�M��O�T�7��-2����x
¹t���h�����&s�E&ź����8�CJ]���u�#E��@$}�Cn��(X�7)@��+��������!�'t.���?��CQ�Y9`�*�i�r�l�� i���_� �S��$H��|@��@���H���[��~w�c��������!��ZP��H6��1���ĵ���ʗ�ꊻ]&���y���k؈��8��{��6;����Ļ!�˻��˻�ƻ۽������¢�a����������ro���f��Q���)f��I�������»�F��V����������찻V2���]��Smƻ�Bֻ���K���/A�o��*
�%)�����Tﻄ�㻅gܻ+ۻޔ��b컖v��������I���  �  i��<k��<ŧ�<�R�<�S�<��<���<Wx�<%��<Wg�<�5�<M��<B��<���<���<��<}t�<���<���<���<0��<��<��<ӈ�<V��<�]�<U��<+
�<-��<"D�<}�<��<��<��<�<��<��<���<���<H��<���<�d�<Z��<��<�#�<+�<�Q�<���<��<��<HU�<K��<U��<|n�<V��<�N�<���<�5�<'6�<���<���<��<��<5�<p��<%�<ڭ�<�L�<�}�<f��<g�<�y�<Z��<J�<�"�<@��<�"�<K��<|t�<L��<K߮<X�<w�<gO�<�^�<~��<P��<��<KN�<�١<IF�<�s�<�~�<���<�j�<�"�<�=�<N�<	��<n��<���<�=�<Af�<*�<s�}<P�v<+�m<Hc<'�W<1"M<�D<ړ=<�&:<�9<P;<��=<S�?<W�?<�k<<��5<�[,<J� <�<�f	<� <&z�;Ԓ�;Wf�;��;�?�;a� <=(<��;�;�.�;�M�;O&�;�|�;q̨;��;Ԇ�;��;���;���;�;�*|;�g;нH;a�!;{��:���:;o�9<�����蹝��ӄ���q����Rh� ׈��2���Fj�f'���
�C4�SkW�=vo��y�}v��+h���R�� <�T�(�0��)����o�,�Q=���N�kF]�еf���i�}&f��O]�i�Q�c2F�B�>�34>��F���X�|s��m��5����٥��ﭻ��G����2��>Ǖ��d��h	���x��G}����󘕻糧A�������AUȻ�ȻK�»_ٸ�2����ߠ�T������jۓ�I���xe��ѩ��	�����;)��f����־��Ժ��㵻�����K?���$����Ļ�Իz�������� �*�Qs����ԁ���|����cۻ�+ڻH�߻p����`��-y�����  �  ���<�C�<���<63�<
��<T!�<���<d�<*u�<���<���<ך�<��<)��<�
�<���<Sf�<�[�<am�<�4�<~R�<���<���<l��<D �<�P�<b��<�f�<�1�<�o�<� �<�w�<z.�<Mo�<���<�s�<|��<*��<�O�<$��<T��<Z��<�9�<�+�<�9�<���<ް�<���<L�<��<���<QW�<t[�<O�<ґ�<�h�<���<�<�<l�<:L�<�r�<�$�<=	�<���<���<`Q�<_`�<�T�<���<�<���<w��<�m�<I��<m"�<���<���<P1�<�4�<��<�O�<���<8�<S��<���<�,�<���<��<���<ķ�<��<��<��<TM�<�-�<��<�J�<�"�<Գ�<h��<�ф<��<g��<Ꮑ<�~<gx<Op<�=f<��[<xtQ<�H<UUB<o�><�=<Q�><Zd@<O�A<f�@<��=<�%7<.<5#<��<�A<��<J��;���;� �;���;�<.�<��<�� <�)�;6p�;��;�}�;'r�;S6�;j��;R�;E�;ӎ;de�;��;�V�;�Ol;��O;v�+;U�;d?�:�G9:�zQ9-J"�����Ᾱx���?6�>D����@�v�׹,�R��Ԯ�����&���F��]�
�f���c�aW���D�O�0��� �b���Q��{�o�'��~7���G��U�X�]�v�`���]��#V���K��VA��|:���9�g2A��5Q���h�U����Ɛ�b���tr��㿦�(W��*#���/���@���.z��s���x��z���%����C>��'/��g��3��鹻�谻����曻Rh���鐻����xb���ݝ������R���I��ز���-��Nົ�t������n��w��������ot��r<λ}�ݻ�:�W�����������r���-��Kd���޻`�ػ��׻Aݻ5�˾��_�� �	�*~��  �  �]�<6��<��<%��<���<���<���<���</��<i��<u��<I��<���<}�<?��<@i�<x��<�`�<�,�<Y��<���<�&�<���<�>�<U>�<6�<��<���<Ξ�<���<s��<��<V��<���<f�<�&�<c��<F�<�7�<k�<���<v�<8��<:x�<�%�<�N�<�v�<=&�<��<O�<f^�<���<�?�<�|�<� �<���<Џ�<J��<�N�<�6�<��<���<܌�<��<{��<���<7��<+�<���<݁�<P �<T��<���<��<8y�<�s�<�O�<�ݿ<�*�<&�<fY�<=Y�<b�<y��<�<R�<`�<+ʣ<P�<'��<7��<�p�<���<���<�$�<�O�<&Ɏ<���<RG�<�`�<��<(΄<r��<�<[�<�+z<��r<fj<G�`<��W<�O<�EI<&EE<tyC<�[C<X�C<�D<Z�B<}�><��8<�a0<��&<�N<�<T<9<֛<�<��<u<x<C|<y�<2$�;��;�C�;��;o��;%��;�6�;f+�;�O�; �;���;T��;���;?�q;;X;118;:J;v9�:��:+#:��9�?m8�ʷC=[����7���7�)���H����4��՘��ߺ9��d�.�xB�L�J�mTI�w�?�$�1��"���������S�z�"��M0�!>�T�I�2Q���S�N2R�qL��<D�?�;��U6�c�5��M;��H��4[��r��K��v���`����B��a��s搻�K��S��r���m�l�r��\���������W�������H^��^�����*ॻ~a��P���A���9�������9��j���`Ģ�X<���G���?��o絻V��#����˯�����󫻡������%-����ƻ�ӻ�"�7l�]������Gq黣J�Y�ٻLaջ�-ջ�ٻ���y������Q���  �  {D�<�f�<d7�<Rm�<���<N��<3�<���<�	�<>��<HD�<>��<K�<�1�<s�<��<]	�<uI�<��<}��<��<�^�<>�<���<�I�<m��<.�<���<ā�<?�<@��<���<�^�<��<�<���<���<���<<�<z��<���<N��<��<��<'C�<d��<��<��<�o�<�:�<�y�<�Q�<���<7��<���<��<T�<A�<8��<���<�w�<r��<p��<���<��<�{�<��<�*�<��<�T�<���<���<���<��<��<+4�<��<X^�<��<��<��<rD�<֔�<]��<Uا<4��<4�<�ܥ<�W�<\Y�<û�<�x�<(��<Wh�<���< ��<�g�<$��<r�< ۈ<T
�<8v�<��<�8�<�&�<{-{<��t<%�m<��e<�^<oW<�Q<��L<iJ<�H<�G<�VF<��C<�?<�9<|�2<D�)<�@!<(7<�<^�<R<�	<h	<ت<�<�w<��<�m�;R��;E��;��;���;���;���;�	�;��;��;��;���;�3�;�Et;��];�B;,$;�;	��:7��:@�D:��:L�9���9�o9��9�I���5��$��*��"��ݟ������=#�^+���+���&��0��������������^�K��1�*���4�/G=���B��E��E�Q�B��>�g�8��W5��4��8�+�A�O�T%`��?r�g?���$���쉻�=��X�������Jt���k�Wji�^�m�iCy�j�,���݀���M��ࡻ����$��QN���ؔ�96�������7��o^������x0��>S������©�v��� ������î��M��~񫻎������Ѱ����-|���Lɻ�ӻM�ۻ+P������߻{�ٻV3ջ@�һ�ӻ}׻^޻�经��-����� ��  �  ���<0��<P�<h��<���<
��<���<+�<�X�<H[�<O�<nO�<�o�<��<�<R��<��<���<r��<1n�<b1�<���<-�<��<5��<��<��<?)�<�)�<ԧ�<���<��<[��<��<�3�<��<��<���<r��<,d�<�+�<m�<p2�<�h�<���<���<���<�!�<���<���<���<%�<�0�< p�<���<jR�<��<3��<�Z�<8@�<"6�<"�<V��<�b�<݃�<z>�<y��<x��<<��<���<BR�<C�<t9�<��<��<l��<g��<ln�<ro�<���<�d�<S�<�د<SO�<�Q�<>ǩ<��<�I�<`�<�*�<��<���<��<�:�<�\�<щ�<D͑<�$�<@��<s�<ܿ�<֚�<|��<◁<;<=�z<
�u<
p<�j<5�c< �]<u|X<+�S<�4P<�>M<�J<��G<trD<)�?<�f:<p�3<'�,<9�%<�<[�<� <��<�N<0<�
<N><+�<� <i��;Z��;G��;���;ky�;��;[F�;��;Tc�;�X�;@�;�߈;*��;&p;`
];�G;�/;ۇ;ȱ�:u�:��:��s:D�::v�:���9	m9d6�7��m�����f�e&���ͺ���������5��!�r��Y7����8 ��j�jV�K"�K�(��^.���2��_6�+	9�:�:��;���;�b�:�5:���:�D�<�VRA��H��R���]��h�1eq�O�v��|x�=Kv�͋q��Cl�w�h��eh��l�u�0L������|��1ݐ��H��t�6����Đ�&ڎ�ƍ�<���}����8���ŕ�a���k����%�����m���t਻�������;㬻?���rO���¯�o@��T��a��DM����ǻ��ͻb�һ��ջ�ֻ��ջ��ӻ�һ{gѻU�һJֻb�ۻ�%�������!��  �  W��<+h�<��<��<���<0�<3O�<�o�<��<o	�<��<�K�<b
�<���<�1�<�t�<ʍ�<ܚ�<%��<� �<Yv�<��<���<�o�<� �<	f�<!��<��<'�<qP�<���<Gs�<�<�<��<	��<�Q�<���<���<���<�7�<5��<<�<&��<���<���<bA�<!��<��<Vk�<I��<�<�<���<H��<^��<@��<g�<��<]c�<ܟ�<4��<' �<Y��<��<���</c�<F��<z0�<4�<N��<��<��<���<O�<p��<���<�<�<�9�<��<�=�<Bm�<ޘ�<��<�\�<��<��<߫<vϩ<|��<�O�<�ܢ<^�<��<��<)@�<Q�<��<`��<�D�<D��<���<�ׇ<��<�^�<��<��{<`�w<@�s<:p<�l<1�g<"�b< 0^<XxY<�T<}�P<�aL<<.H<g�C<��><~�9<��3<�/.<ʢ(<�}#<��<��<��<*<2<<<b�<V�<�F�;���;P��;��;T��;�
�;���;�;�,�;���;��;��;d��;}jt;Jbc;eS;8�C;�-3;�d!;FF;c��:���:���:0��:.�<:5��9ϣr9,���񑹜���[��p��i���V�ɺQ|޺���I����m�3	�h������M��U#��(�;+��\,��,�F�,��-��-0�cd4���9��>��yC�ȱF�,�H��vI�iJ�&K��\M�Q�kV��T[�9S`�xXd�g�|vh��4i��j�g6l�zp�ķu��I|�_g��H<���f���釻n�������\?��h$���ŏ��蒻U,���2������$t��s����{��L���@(������f��'Ы��m��ދ������ὶ�i��^t������n���r��,�û�fǻO�ʻ0ͻvϻ�\лWhѻa�һ��Ի��׻|ۻ��޻_�����63��  �  �|�<l��<���<sp�<���<�4�<ֹ�<ʘ�<���<��<��<���<o��<��<���<���<�Z�<G��<H�<!��<���<�A�<�H�<e��<��<Ms�<s��<
N�<��<���<��<�<�#�<Y^�<���<�2�<2��<�n�<EA�<�/�<�!�<���<���<���<+	�<���<�R�<��<u��<���<֤�<���<p�<�#�<��<D��<px�<h��<�1�<��<�)�<`��<�B�<���< �<yT�<ٌ�<!��<2	�<��<f��<��<���<��<֎�<�J�<=�<b��<'c�<%�<��<��<��<E��<�]�<�ì<��<���<i��<�_�<%��<G	�<~�<�j�<�	�<]��<��<�<�<�Ɗ<:7�<���<r>�<:�z<�v<T�r<��o<�m<<�k<��h<�e<��a<��\<��W<<R<�L<� G<��A<N�<<Ά7<ȯ2<{-.<�*<L&<� "<o�<�y<�m<a�<��<Ǘ<7g�;���;R��;ѿ�;T��;��;{��;	��;�Q�;���; 4�;aÕ;�{�;�t;�_;a�M;9T@;z�5;��,;�s";�;��;���:O.�:ʞ�:{1R:z6�9��#9J���aչ��+�O9e�.ꊺ�0���ذ�ߤ��VdӺÐ�o��������a(���2�h�9�>�<�=;��l6��0���+���)�Nd,�h3�#�<��^H��
S�l[��2_�bf_��[\�*YW�)R��GN���L�fcN��FR��X�/�^���e�j�k�E�p�u��x���{���}� �~������)〻�ւ�G��y���._��/���s���[���d��9i��瘤������w���.��=�����lt���4��_=�������»y�»����I���}���㽻���̕��˴û,�ǻ��˻=�ϻuӻ-�ֻ�-ٻMۻ$iݻt�޻��߻�g�d��  �  �!�<��<�d�<2�<Z��<F�<�A�<��<�v�<h��<���<O,�< K�<���<��<�r�<5��<["�<8��<��<�"�<`��</��<���<]#�<�h�<�R�<K��<�p�<j��<�c�<g��<1n�<J&�<�0�<ȗ�<�\�<{�<{��<�X�<J��<w��<0�<,�<>a�<9�<���<]��<c"�<zH�<O�<�$�<���<��<$0�<ΰ�<cT�<d�<m$�<���<���<���<2��<B\�<~��<l��<���<���<��<>��<�b�<���<��<�d�<(��<���<LP�<��<p�<�D�<�<�)�<�m�<R�<C��<9��<�ۨ<8Ӥ<���<��</͙<�e�<�Е<4�<O[�<ܶ�<���<��<�Ӎ<3.�<��<���<�z<�s<q�n<%�k<{j<�]i<M�h<�h<�*f<��b<�h^<>�X<WR<�K<_�D<3�><vK9<�v4<C[0<�,<g�)<z�&<�f#<�+<!�<h�<@><Nd<�R�;m�;0 �;r��;���;�9�;\G�;�Y�;���;�%�;���;4C�;��;��|;�];-cC;�01;�&;�W ;��;I�;��;V�
;��:���:���:UP:�.�9��7Gʥ�M���EV��߀�k7��곛��񦺍c��ϵɺ���h����� .���@��9O�9�V��1W�3�P��E�T~9�3�/�'0+��p-�S�6�OE���V�dh�B@u��1|�x1|�"v� �k�"K_��ET�F�L�n<J�u�L�r?S�Y]��*h���r��{��쀻����䂻�ꁻ���ڑ|��z��3|����b���2g��Ǘ��j��|੻�读`���u	��7o��u5��r ��ޠ�֟��<죻򎪻r���������ƻ�iͻ��л��л�ͻ��Ȼr�û�ȿ�J���%������L�ŻA�˻��ѻ��׻<_ܻt�߻vộ�ỉ�;�߻{�޻{�޻�  �  9��<F��<}?�<I�<��<���<6{�<[	�<���<E��<}d�<r�<�7�<1�<��<C��<�T�<7>�<X�<�8�<�_�<��<�3�<ʡ�<���<���<�T�<L@�<O�<2��<��<�C�<`Y�<���<qt�<���<s��<6�<p�<��<���<y��<��<�[�<P��<��</��<�:�<�G�<�j�< ��<6-�<J�<`��<DG�<l�<5��<�:�<��<���<���<�.�<��<bw�<�9�<]��<��<�-�<�&�<s2�<�:�<OR�<���<K��<"D�<�,�<4s�<�0�<ji�<��<��<dµ<c>�<s �<�>�<،�<%�<�R�<ɉ�<nA�<�ٕ<�<2c�<�#�<sY�<-k�<�ˑ<��<�5�<�.�<:V�<^~<��t<|�l<�)g<" d<�Ec<j�c<ye<V�e<�e<=�b<[J^<$dX<dSQ<x�I<,=B<�q;<��5<�1<z-<L�*<��(<-M&<K%#<�<b�<�-<�W<���;���;�:�;^w�;2�;�9�;�V�;s�;�+�;�~�;|;�;�;���;]��;~;h;�$C;��%;Ѥ;�	;�/;��	;�g;ۀ;�;���:w�:9�:XN=:hɋ9M�%���LS����IV���Ŝ��ġ����s���vRͺ�`�	@�.*��=E���\���m�`�u�K}s��\h��pW��^E� �6���/�p�1��l=���P�rh��,�����y��!���2L���Ɓ��eq��`��"S��L��KM��LT�) `�`wn�Ѧ|�1+�����o�����Zo���セ����{�t}������J�������������舸��|�����_���7Z��4��87��~��Ǣ��m���5��22ǻ�.ӻ%�ۻ�R໤�߻�^ۻEԻ=�˻��Ļ����[/���dƻF�ͻ�ջW$ݻo㻺��#=�-z�=����;{߻�޻�  �  �X�<V��<���<XE�<�g�<���<��<��<���<���<��<���<%�<4e�<�]�<s��<��<oo�<^��<�I�<1�<A�<��<���<Z"�<���<l
�<rk�<\��<i	�<�}�<k�<�7�<�E�<#��<�2�<�A�<U��<��<6�<�<�<&;�<�K�<b�<��<�,�<N�<f��<��<8��<*��<7�<�<�D�<�_�<�<�B�<I�<M��<t�<U�<?Z�<=�<���<��<�<�<Rx�<A��<an�<��<I��<W��<B��<-��<~��<Cǻ<؈�<H�<2Ѷ<���<��<)��<|��<ce�<�C�<~H�<�ڟ<!��<��<Z�<G,�<�]�<g��<'s�<��<��<Hi�<&r�<E�<Ѿ�<kz<�3o<�`f<�\`<�`]<[]<"�^<��`<h�b<0#c<}Xa<`O]<IW<��O<2�G<_�?<�Z8<�a2<��-<�*<��(<'<[%<�"<�n<v�<9I<A<�V�;�X�;��;?��;>3�;r�;�G�;S��;���;	q�;��;Q�;��;���;k�U;]3,;/;%�:Ë�:�P�:��:5��:ܕ;
A;�d�:q'�:�:��#:�9n`��Z�9�����L��ʧ�ݬ���r���������E�׺�s �����;��_[���v�W���ri���3���}���g�h;Q�~�>���5���7�gE�%\��x��񉻙딻@��Z��|M��:%��-Ձ��pm�\��pR�jyQ��{X���e�$�u�;�����
s������r������Tf��W�� �������Յ�Q6��7��S0��tй���ŻTLͻ6:ϻW~˻27û�����u��	{��ď�����p��8����л�B޻X�軪�0��=���޻�4Ի�ʻ��û�s���1û��Ȼ��лj�ٻ�g�,黓F��l�컔Q�Q����O���  �  ��<���<��<���<X��</��<j��<�<�<�R�<F��<��<6��<'1�<-��<���<�1�<�!�<$�<���<oH�<��<���<���<���<-Q�<x\�<k��<���<�+�<g��<���<��<S]�<HF�<���<5�<�4�<��<�J�<ە�<dy�<ې�<��<�b�<i�<-�<!,�<���<�y�<ư�<ހ�< ��<���<���< }�<���<�v�<ʁ�<#:�<�7�<�9�<���<��<:��<ة�<���<��<�#�<��<0��<��<�,�<�D�<���<��<K��<���<�c�<�ܶ<d�<�8�<um�<��<�<��<�5�<�ڣ<g�<oh�<_��<��<?ߍ<�M�<A�<��<��<1�<َ<�Ջ<?D�<_��<��v<wqk<�b<��[<˳X<r�X<N�Z<��]<dx`<�ya<� `<AE\<%1V<؁N<�	F<	�=<%26<�0<+�+<?�(<��&<+�%<�#<l� <�.<�*<?�< *<���;Ë�;�)�;00�;+X�;W-�;���;^��;�9�;���;���;uP�;PP�;OOy;A�H;%;æ�:��:9��:�ӽ:!��:�#�:���:t��:>��:�=�:!�:[9:��8j�[�[�����������8������������ź���ܑ��%�D�H��Ik��C����ڬ��0��������s�,�Y��*E�cJ:��5<��K�Fsd� �������Q���<��_֤��g���I��
�����w��c��W���U�ٽ\��{j���{��؆��3���䒻�^��𲒻����3C��Cs���ၻP�������[J���ʡ��K���6»+	ϻ��ֻ�Rػ�ӻh
ʻw�aa���E���ϧ�7����d���YŻ�1ֻr��6��2q������V�����Q{ڻGQϻIXǻ/�ûMŻ�ʻ8Iӻ�ܻ97滀t��������컍��A�.��  �  3��<1z�<�B�<-�<���<6��<p��<�f�<���<�6�<��<��<��<ׄ�<��<���<���<(��<�W�<���<��<P�<s��<B��<]��<���<	��<�]�<w��<�K�<ĭ�<zr�<�<���<�d�<���<6��<1��<���<!V�<�@�<�W�<O�<s�<ţ�<a��<�q�<��<���<���<ѿ�<A�<�:�<���<22�<��<#>�<"9�<���<���<	��<�<�<�6�<��<X��<��<���<���<��<�p�< ��<���<�<�p�<	��<,�<7�<Z��<�{�<��<+�<�,�<1�<���<mT�<�ͨ<�Q�<&a�<���<���<?�<��<ג�<�L�<қ�<��<u�<���<}��<��<{*�<��u<�j<L�`<Z<9W<�W<ecY<V�\<��_<��`<͡_<��[<��U<1�M<�nE<9�<<?l5<QQ/<��*<�(<�U&<�%<no#<H� <��<;�<�<� <��;�^�;���;յ;�5�;�n�;b��;�<�;H�;��;��;@T�;��;�u;��C;�;��:T��:�ث:��:�:���:wa�:�K�:[�:��:މ�:$�:+���������g�=M��u���A]����O湺���A4ɺ�溣]
��)�?�M��q��~���p��~������k�����w�,#]�xG�%<���=�;^M��g��ƃ�T����J��9���7������?��\����{��f�@Z���W��^�nql��E~�]-��n����y��-�j)���ۏ��^���f��:���0샻�牻ޔ��⣻_鴻mBŻ�Yһ�'ڻ��ۻ�ֻ�x̻�߿�?ӳ��U������������ǻ�gػ�� ������� S�����S�_�ܻ
ѻ(�ȻP�Ļ�.ƻ��˻QԻB4޻��/���U�bJ���"�7����}�����  �  ��<���<��<���<X��</��<j��<�<�<�R�<F��<��<6��<'1�<-��<���<�1�<�!�<$�<���<oH�<��<���<���<���<-Q�<x\�<k��<���<�+�<g��<���<��<S]�<HF�<���<5�<�4�<��<�J�<ە�<dy�<ې�<��<�b�<i�<-�<!,�<���<�y�<ư�<ހ�< ��<���<���< }�<���<�v�<ʁ�<#:�<�7�<�9�<���<��<:��<ة�<���<��<�#�<��<1��<��<�,�<�D�<���<��<M��<���<�c�<ݶ<h�<�8�<{m�<��<�<&��<�5�<�ڣ<o�<wh�<g��<��<Eߍ<�M�<F�<��<��<1�<َ<�Ջ<=D�<\��<��v<mqk<�b<��[<��X<b�X<?�Z<��]<Tx`<�ya<� `<5E\<1V<ρN<�	F<�=<"26<�0<-�+<C�(<��&<3�%<!�#<x� <�.<�*<N�<*<ǰ�;��;�)�;L0�;DX�;m-�;���;l��;�9�;���;���;pP�;FP�;3Oy;�H;�~;_��:���:���:1ӽ:���:f#�:y��:���:ɰ�:=�:� �:�8:��8!k�˴[���������K������ǳ����ź���ݑ��%�D�H��Ik��C����ڬ��0������ߟs�,�Y��*E�cJ:��5<��K�Fsd� �������Q���<��_֤��g���I��
�����w��c��W���U�ٽ\��{j���{��؆��3���䒻�^��𲒻����3C��Cs���ၻP�������[J���ʡ��K���6»+	ϻ��ֻ�Rػ�ӻh
ʻw�aa���E���ϧ�7����d���YŻ�1ֻr��6��2q������V�����Q{ڻGQϻIXǻ/�ûMŻ�ʻ8Iӻ�ܻ97滀t��������컍��A�.��  �  �X�<V��<���<XE�<�g�<���<��<��<���<���<��<���<%�<4e�<�]�<s��<��<oo�<^��<�I�<1�<A�<��<���<Z"�<���<l
�<rk�<\��<i	�<�}�<k�<�7�<�E�<#��<�2�<�A�<U��<��<6�<�<�<&;�<�K�<b�<��<�,�<N�<f��<��<8��<*��<7�<�<�D�<�_�<�<�B�<I�<M��<t�<U�<?Z�<=�<���<��<�<�<Sx�<B��<bn�<��<J��<Y��<D��<1��<���<Hǻ<ވ�<P�<;Ѷ<���<��<6��<���<re�<�C�<�H�<�ڟ<0��<��< Z�<S,�<�]�<p��<.s�<��<��<Hi�<%r�<A�<˾�<[z<�3o<�`f<�\`<m`]<>]<�^<|�`<J�b<#c<bXa<HO]<�HW<��O<$�G<U�?<�Z8<�a2<��-<��*<Ȥ(<,'<o%<�"<�n<��<VI<4A<�V�;�X�;D��;t��;n3�;��;�G�;n��;���;q�;��;H�;��;���;%�U;
3,;�;P�:ފ�:P�:��:=��:b�;�@;�c�:�&�:@�:R�#:S�9ub��2�9�g���M��9ʧ�����r��'�������M�׺�s �����;��_[���v�W���ri���3���}���g�h;Q�~�>���5���7�gE�%\��x��񉻙딻@��Z��|M��:%��-Ձ��pm�\��pR�jyQ��{X���e�$�u�;�����
s������r������Tf��W�� �������Յ�Q6��7��S0��tй���ŻTLͻ6:ϻW~˻27û�����u��	{��ď�����p��8����л�B޻X�軪�0��=���޻�4Ի�ʻ��û�s���1û��Ȼ��лj�ٻ�g�,黓F��l�컔Q�Q����O���  �  9��<F��<}?�<I�<��<���<6{�<[	�<���<E��<}d�<r�<�7�<1�<��<C��<�T�<7>�<X�<�8�<�_�<��<�3�<ʡ�<���<���<�T�<L@�<O�<2��<��<�C�<`Y�<���<qt�<���<s��<6�<p�<��<���<y��<��<�[�<P��<��</��<�:�<�G�<�j�< ��<6-�<J�<`��<DG�<l�<5��<�:�<��<���<���<�.�<��<bw�<�9�<]��<��<�-�<�&�<t2�<�:�<QR�<���<O��<&D�<�,�<<s�<�0�<ui�<��<��<tµ<v>�<� �<�>�<팫<!%�<�R�<މ�<�A�<�ٕ<Ԍ�<Bc�<$�<~Y�<5k�<�ˑ<��<�5�<�.�<2V�<�]~<��t<\�l<e)g<�d<bEc<@�c<Oe<+�e<�e<�b<8J^<dX<KSQ<d�I<=B<~q;<��5<�1<%z-<^�*<�(<IM&<k%#<&�<��<�-<(X< ��;���;3;�;�w�;I2�;�9�;�V�;*s�;�+�;�~�;|;�;��;���;8��;;h;8$C;)�%;:�;	;#/;��	;g;.�;e�;���:�u�:( �:oL=:Ƌ9�%�O���LS�)���V���Ŝ��ġ�9��������Rͺ�`�@�/*��=E���\���m�_�u�K}s��\h��pW��^E��6���/�p�1��l=���P�rh��,�����y��!���2L���Ɓ��eq��`��"S��L��KM��LT�) `�`wn�Ѧ|�1+�����o�����Zo���セ����{�t}������J�������������舸��|�����_���7Z��4��87��~��Ǣ��m���5��22ǻ�.ӻ%�ۻ�R໤�߻�^ۻEԻ=�˻��Ļ����[/���dƻF�ͻ�ջW$ݻo㻺��#=�-z�=����;{߻�޻�  �  �!�<��<�d�<2�<Z��<F�<�A�<��<�v�<h��<���<O,�< K�<���<��<�r�<5��<["�<8��<��<�"�<`��</��<���<]#�<�h�<�R�<K��<�p�<j��<�c�<g��<1n�<J&�<�0�<ȗ�<�\�<{�<{��<�X�<J��<w��<0�<,�<>a�<9�<���<]��<c"�<zH�<O�<�$�<���<��<$0�<ΰ�<cT�<d�<m$�<���<���<���<2��<B\�<~��<l��<���<���<��<?��<�b�<��<��<�d�<.��<���<UP�<��<}�<E�<��<�)�<�m�<4R�<\��<S��<ܨ<SӤ<���<(��<F͙<�e�<�Е<D�<[[�<嶓<���<��<�Ӎ<,.�<��<狁<��z<��s<E�n<��k<Hj<O]i<�h<�h<�*f<��b<�h^<�X<�VR<�K<N�D<)�><tK9<�v4<Q[0<1�,<��)<��&<g#<�+<Q�<��<t><�d<BS�;qm�;� �;���; ��;:�;�G�;Z�;���;�%�;��;C�;��;/�|;4];�bC;A01;�&;�V ;!�;q�;!�;��
;���:?��:6��:�P:�*�9�ـ74ͥ�|���FV��߀��7������񦺣c��ݵɺ���h����� .���@��9O�9�V��1W�2�P��E�S~9�3�/�&0+��p-�S�6�OE���V�dh�B@u��1|�x1|�"v� �k�"K_��ET�F�L�n<J�u�L�r?S�Y]��*h���r��{��쀻����䂻�ꁻ���ڑ|��z��3|����b���2g��Ǘ��j��|੻�读`���u	��7o��u5��r ��ޠ�֟��<죻򎪻r���������ƻ�iͻ��л��л�ͻ��Ȼr�û�ȿ�J���%������L�ŻA�˻��ѻ��׻<_ܻt�߻vộ�ỉ�;�߻{�޻{�޻�  �  �|�<l��<���<sp�<���<�4�<ֹ�<ʘ�<���<��<��<���<o��<��<���<���<�Z�<G��<H�<!��<���<�A�<�H�<e��<��<Ms�<s��<
N�<��<���<��<�<�#�<Y^�<���<�2�<2��<�n�<EA�<�/�<�!�<���<���<���<+	�<���<�R�<��<u��<���<֤�<���<p�<�#�<��<D��<px�<h��<�1�<��<�)�<`��<�B�<���< �<yT�<ڌ�<"��<3	�<��<h��<��<���<��<܎�<�J�<H�<n��<6c�<0%�<��<��<��<`��<�]�<�ì<��<���<���<�_�<?��<^	�<��<�j�<�	�<g��<��<�<�<�Ɗ</7�<���<_>�<�z<�v<�r<O�o<��m<�k<k�h<��e<{�a<��\<w�W<�;R<֡L<� G<��A<L�<<Ն7<ׯ2<�-.<*<s&<� "<��<�y<.n<��<�< �<�g�;��;���;"��;���;#��;���;��;�Q�;���;�3�;.Õ;_{�;s�t;_;��M;\S@;��5;��,;�r";�;��;���:�,�:U��:�.R:�1�9�#9Ў�odչ��+�:e�{ꊺ�0���ذ�����fdӺ͐�u��������a(���2�g�9�>�<�=;��l6��0���+���)�Md,�h3�#�<��^H��
S�k[��2_�bf_��[\�*YW�)R��GN���L�fcN��FR��X�/�^���e�j�k�E�p�u��x���{���}� �~������)〻�ւ�G��y���._��/���s���[���d��9i��瘤������w���.��=�����lt���4��_=�������»y�»����I���}���㽻���̕��˴û,�ǻ��˻=�ϻuӻ-�ֻ�-ٻMۻ$iݻt�޻��߻�g�d��  �  W��<+h�<��<��<���<0�<3O�<�o�<��<o	�<��<�K�<b
�<���<�1�<�t�<ʍ�<ܚ�<%��<� �<Yv�<��<���<�o�<� �<	f�<!��<��<'�<qP�<���<Gs�<�<�<��<	��<�Q�<���<���<���<�7�<5��<<�<&��<���<���<bA�<!��<��<Vk�<I��<�<�<���<H��<^��<@��<g�<��<]c�<ܟ�<4��<' �<Y��<��<���</c�<G��<z0�<4�<O��<���<��<���<S�<u��<���<�<�<:�<��<�=�<Tm�<�<��<�\�<��<��<%߫<�ϩ<���<�O�<ݢ<7^�<��<#��<;@�<_�<��<f��<�D�<A��<���<�ׇ<��<�^�<��<i�{<(�w<�s<�p<Rl<��g<��b<�/^<'xY<��T<Y�P<�aL<(.H<\�C<��><��9<��3<�/.<�(<~#<��<��<(�<d<o<<J<��<��<G�;B��;���;��;���;�
�;���;�;�,�;`��;g�;��;��;�it;vac;0dS;G�C;�,3;�c!;PE;���:9��:9��:���:z�<:z��9��r97G����������[�q������~�ɺl|޺���T����m�3	�h������M��U#��(�:+��\,��,�F�,��-��-0�cd4���9��>��yC�ȱF�,�H��vI�iJ�&K��\M�Q�jV��T[�9S`�xXd�g�|vh��4i��j�g6l�zp�ķu��I|�_g��H<���f���釻n�������\?��h$���ŏ��蒻U,���2������$t��s����{��L���@(������f��'Ы��m��ދ������ὶ�i��^t������n���r��,�û�fǻO�ʻ0ͻvϻ�\лWhѻa�һ��Ի��׻|ۻ��޻_�����63��  �  ���<0��<P�<h��<���<
��<���<+�<�X�<H[�<O�<nO�<�o�<��<�<R��<��<���<r��<1n�<b1�<���<-�<��<5��<��<��<?)�<�)�<ԧ�<���<��<[��<��<�3�<��<��<���<r��<,d�<�+�<m�<p2�<�h�<���<���<���<�!�<���<���<���<%�<�0�< p�<���<jR�<��<2��<�Z�<8@�<"6�<"�<V��<�b�<݃�<z>�<y��<y��<<��<���<CR�<F�<w9�<��<��<u��<q��<yn�<�o�<���<�d�<j�<ٯ<nO�<�Q�<[ǩ<#��<J�<}�<�*�<��<��<��<;�<�\�<ۉ�<J͑<�$�<=��<k�<ѿ�<ƚ�<i��<̗�<
<�z<ёu<�p<�j<��c<��]<A|X<��S<�4P<�>M<��J<��G<irD<'�?<�f:<��3<?�,<Y�%<�<��<� <*�<�N<J0<;�
<�><b�<$� <Š�;���;���;ǈ�;�y�;���;\F�;��;1c�;jX�;��;P߈;κ�;8%p;�	];/�G;+�/;�;��:��:;�:f�s:Y�::٥:��95m9#�7.�m�����f��&��E�ͺ�� ����6��!�t��Z7����7 ��j�jV�K"�K�(��^.���2��_6�*	9�:�:� �;���;�a�:�5:���:�D�<�URA��H��R���]��h�1eq�O�v��|x�=Kv�͋q��Cl�w�h��eh��l�u�0L������|��1ݐ��H��t�6����Đ�&ڎ�ƍ�<���}����8���ŕ�a���k����%�����m���t਻�������;㬻?���rO���¯�o@��T��a��DM����ǻ��ͻb�һ��ջ�ֻ��ջ��ӻ�һ{gѻU�һJֻb�ۻ�%�������!��  �  {D�<�f�<d7�<Rm�<���<N��<3�<���<�	�<>��<HD�<>��<K�<�1�<s�<��<]	�<uI�<��<}��<��<�^�<>�<���<�I�<m��<.�<���<ā�<?�<@��<���<�^�<��<�<���<���<���<<�<z��<���<N��<��<��<'C�<d��<��<��<�o�<�:�<�y�<�Q�<���<7��<���<��<T�<A�<8��<���<�w�<r��<p��<���<��<�{�<��<�*�<��<�T�<���<���<���<��<���<34�<%��<d^�<��<��<-��<�D�<씬<u��<nا<O��<"4�<�ܥ<�W�<uY�<ڻ�<y�<;��<gh�<���<	��<�g�<%��<o�<ۈ<J
�<*v�<��<�8�<�&�<K-{<y�t<��m<��e<g^<=W<YQ<��L<DJ<єH<�G<�VF<��C<�?<�9<��2<Z�)<�@!<K7<.�<��<�<�	<�	<�<$�<�w<��<�m�;���;���;:��;���;��;���;�	�;h�;s�;r�;���;�3�;Et;��];C�B;E+$;E�;]��:���:+�D:�:��9܄�9W o9��9f��Z8����c*��g�����	���=#�!^+���+���&��0��������������^�J��1�*���4�.G=���B��E��E�Q�B��>�g�8��W5��4��8�+�A�O�T%`��?r�g?���$���쉻�=��X�������Jt���k�Wji�^�m�iCy�j�,���݀���M��ࡻ����$��QN���ؔ�96�������7��o^������x0��>S������©�v��� ������î��M��~񫻎������Ѱ����-|���Lɻ�ӻM�ۻ+P������߻{�ٻV3ջ@�һ�ӻ}׻^޻�经��-����� ��  �  �]�<6��<��<%��<���<���<���<���</��<i��<u��<I��<���<}�<?��<@i�<x��<�`�<�,�<Y��<���<�&�<���<�>�<U>�<6�<��<���<Ξ�<���<s��<��<V��<���<f�<�&�<c��<F�<�7�<k�<���<v�<8��<:x�<�%�<�N�<�v�<=&�<��<O�<f^�<���<�?�<�|�<� �<���<Џ�<J��<�N�<�6�<��<���<܌�<��<{��<���<8��<+�<���<ށ�<R �<V��<���<��<<y�<�s�<�O�<�ݿ<�*�<3�<tY�<NY�<t�<���<-�<R�<2`�<@ʣ<e�<;��<J��<�p�<Ɔ�<���<�$�<�O�<*Ɏ<���<PG�<�`�<��<΄<d��<�<7�<`+z<��r<;j<�`<q�W<�O<�EI<EE<UyC<�[C<D�C<�D<R�B<{�><µ8<�a0<��&<�N<7�<)T<29<��<'<��<�<=x<k|<��<u$�;L��;D�;@��;���;2��;�6�;Y+�;�O�;��;Y��;��;O��;��q;u:X;�08;�I;8�:t�:�#:��9�m8tGʷN�[�њ�7�[�7w3���J��|�4�&֘�ߺN��s�.��B�R�J�qTI�z�?�%�1��"���������S�z�"��M0�!>�T�I�2Q���S�M2R�qL��<D�?�;��U6�c�5��M;��H��4[��r��K��v���`����B��a��s搻�K��S��r���m�l�r��\���������W�������H^��^�����*ॻ~a��P���A���9�������9��j���`Ģ�X<���G���?��o絻V��#����˯�����󫻡������%-����ƻ�ӻ�"�7l�]������Gq黣J�Y�ٻLaջ�-ջ�ٻ���y������Q���  �  ���<�C�<���<63�<
��<T!�<���<d�<*u�<���<���<ך�<��<)��<�
�<���<Sf�<�[�<am�<�4�<~R�<���<���<l��<D �<�P�<b��<�f�<�1�<�o�<� �<�w�<z.�<Mo�<���<�s�<|��<*��<�O�<$��<T��<Z��<�9�<�+�<�9�<���<ް�<���<L�<��<���<QW�<t[�<O�<ґ�<�h�<���<�<�<l�<:L�<�r�<�$�<=	�<���<���<`Q�<_`�<�T�<���<�<���<x��<�m�<K��<p"�<���<���<V1�<�4�< �<�O�<���<E�<a��<���<�,�<���<��<���<ҷ�<��<��<��<]M�<�-�<�<�J�<�"�<ҳ�<d��<�ф<��<]��<֏�<��~<�fx<2p<�=f<��[<ZtQ<�H<:UB<W�><ӣ=<?�><Ld@<E�A<`�@<��=<�%7<.<5#<	�<�A<�<~��;7��;� �;;��;�<K�<��<�� <*�;_p�;��;�}�;:r�;\6�;j��;I�;3�;�Ҏ;Ae�;��;�V�;WOl;Y�O;��+;��;k>�:�E9:fsQ9NQ"�.���侹2���6�cL���@�ׅ׹��R� ծ�����&���F��]��f���c�aW���D�O�0��� �b���Q��{�n�'��~7���G��U�X�]�u�`���]��#V���K��VA��|:���9�g2A��5Q���h�U����Ɛ�b���tr��㿦�(W��*#���/���@���.z��s���x��z���%����C>��'/��g��3��鹻�谻����曻Rh���鐻����xb���ݝ������R���I��ز���-��Nົ�t������n��w��������ot��r<λ}�ݻ�:�W�����������r���-��Kd���޻`�ػ��׻Aݻ5�˾��_�� �	�*~��  �  i��<k��<ŧ�<�R�<�S�<��<���<Wx�<%��<Wg�<�5�<M��<B��<���<���<��<}t�<���<���<���<0��<��<��<ӈ�<V��<�]�<U��<+
�<-��<"D�<}�<��<��<��<�<��<��<���<���<H��<���<�d�<Z��<��<�#�<+�<�Q�<���<��<��<HU�<K��<U��<|n�<V��<�N�<���<�5�<'6�<���<���<��<��<5�<p��<%�<ڭ�<�L�<�}�<f��<g�<�y�<[��<K�<�"�<B��<�"�<N��<�t�<Q��<Q߮<^�<~�<nO�<�^�<���<X��<��<SN�<�١<PF�<�s�<�~�<���<�j�<�"�<�=�<N�<��<l��<���<�=�<<f�<$�<e�}<A�v<�m<oHc<�W<""M<�D<̓=<�&:<٦9<�O;<��=<N�?<T�?<�k<<��5<�[,<P� <��<�f	<� <Az�;��;vf�;	�;@�;q� <L(<,��;&�;�.�;�M�;]&�;�|�;v̨;��;І�;���;���;w��;ݸ�;q*|;vg;��H;#�!;���:��:=m�9�������z�������������Th��׈�[3��CGj��'���
�K4�XkW�Avo��y�}v��+h���R�� <�T�(�0��(����n�,�Q=���N�kF]�еf���i�}&f��O]�h�Q�c2F�B�>�34>��F���X�|s��m��5����٥��ﭻ��G����2��>Ǖ��d��h	���x��G}����󘕻糧A�������AUȻ�ȻK�»_ٸ�2����ߠ�T������jۓ�I���xe��ѩ��	�����;)��f����־��Ժ��㵻�����K?���$����Ļ�Իz�������� �*�Qs����ԁ���|����cۻ�+ڻH�߻p����`��-y�����  �  T�<��<z��<�.�<U��<a��<��<�k�<V�<���<�q�<���<��<{�<�&�<�</��<���<��<d<�<���<f �<�#�<�m�<��<`r�<��<</�<�9�<�;�<� �<'��<�f�<��<Ƥ�<$]�<Z��<3��<���<�;�<���<�}�<���<�d�<���<��<���<���<��<�$�<���<}��<�4�<���<�<��<�G�<���<�l�<z��<T#�<E�<���<x�<�2�<��<�L�<�S�<H��<�p�<��<K��<~��<�*�<k��<n�<�L�<���<*�<�.�<���<���<��<��<~��<�֮<�c�<l4�<�έ<^ˬ<��<Y#�<���<[e�<��<�З<��<5�<���<y�<�<lw�<��<~�<���<�|�<Nu�<�x<Aw<so<��g<fCb<�k^<�V\<Ǜ[<ـ[<z[<7mY<��U<��O< �G<
�><u5<g�,<\�%<Vc <+<Z�<�I<�<�(<��<��<�<�<k�;���;�z�;�Q�;���;鶷;�R�;�"�;	�;֪�;���;��;;Е;�y�;=Kq;��O;�;/;|�;��:��:_'�:�D�:��:�:�:��:'�o:���9�Y��Vz�/ej��̚�����]����𲕺�"��5�n�Z�m�����Wٜ�N���?���]�����| �������
�g*��A��ٺ�ںV%��)����;$)��:�)OE��NI�*�E�Y�;���-�0��>��>���i"�I6�{UL��Ta�y�q��.{��	}�h�w�]�m��za�15W���Q��LS�O�[�m�j�25}�K����ߑ��*��/����(��ӫ��)Ι����*k����������Kތ���������q���SL��-���S���{��l=��o��,t��S?��$d��we��-ܫ�]L���I���ʻ�Dջ��ܻ�  �  ��<	��<rT�<���<���<c��<�0�<H��<�4�<M$�<z��<w8�< 
�<Lk�</��<_�<Z��<���<E�<�q�<�,�<|3�<a�<V��<�p�<���<�}�<4��<���<���<���<v��<��<���<R��<�c�<M�<G��<�7�<��<c�<��<Hx�<	��<��<���<��<���<��<U�<~��<,��<�y�<�:�<p`�<�$�<|��<���<���<��<�^�<%w�<��<$��<�s�<`�<R��<���<�<���<��<B��<�<Ck�<���<Z~�<�P�<B��<���<�Z�<Jǽ<mX�<W|�< |�<s�<kO�<FѮ<w��<d�<v�<�<�Q�<Խ�<N��<�P�<'#�<�f�<OP�<3��<\�<�[�<U��<�(�<�N�<"�<���<㽃<2�<~x<:p<��h<AAc<H[_<~(]<�B\<��[<Z[<�Y<��U<��O<�5H<�D?<�6<[�-<{�&<K[!<�$<C�<W<�<��<i6<��<9�<�f<N�;���;���;l��;=y�;�*�;-��;jU�;��;���;�q�;7��;�ϖ;*��;�Nt;S;�3;S�;9�;�?�:�b�:��:K�:���:&��:V�::�q:��9�+7����\��$��-���z��񝠺*H����{�ef��f���� ���1N��`���8����S.�ڔ�e��� �����k����⺽�ֺe�׺��� ����I�%�h$6��WA��|E��HB�T�8�ы+��������Z��1�!�@�4�HJ��X^�8%n�Pw�xy�xt��j��y^�M�T��O�`�Q��TZ���h�zD{��y����������<��[���$P��3�������͈���劻�ɉ�M���ט�����P��Iq���ƶ��	��U���	���3Ƕ�A���긪��-���M������ѳ��k��&�ɻʫӻ��ڻ�  �  ��<���<դ�<}��<���<m��<���<��<��<���<�e�<��<���<�q�<��<Bb�<N��<���<���<��<K��<���<�<m��<}s�<��<Y��<��< �<a��< ��<4��<��<N;�<M��<pl�<�4�<�@�<J��<h��<o��<+L�<u��<]B�<�H�<���<��<���<=��<9��<
]�<�g�<�7�<x�<[�<.�<���<>��<��<���<���<2��<#v�<k6�<��<<�<=��<f�<�j�<O�<e��<#�<2��<��<��<o��<S�<��<N��< ��<|��<�W�<y��<�ѳ<�ұ<��<��<���<L�<Z��<W��<Jʨ<�C�<�E�<)�<�<g�<�[�<� �<}S�<7�<�t�<���<�Ҋ<bg�<�P�<��<�
�<fz<2�r<��k<�f<D�a<On_<�
^<�*]<��[<�Y<w�U<> P<x�H<�_@<�7< �/<�)<j$<S� <B3<eh<ұ<�8<�c<��<U�<|�<���;EV�;��;���;��;�N�;�y�;v��;Uٰ;�٭;���;��;kp�;�	�;ŗ|;t�\;�>;�#;��;*��:T��:�+�:w��:���:�*�:�ަ:�^w:��:���8e���>�6�o1{��r���@��� ���{���^�dXO�Z�T�Baq�{h�����O�Ժ,h��p��&��5=�
�o�����r�y}ں�*Ϻ��κ�ۺ�9��	���2+�3"6�A�:���8�1�&�%����$C�ܵ�6R�����0� �C�XV��<d��el���m��6i��\`��7V��"N���J�U{M�ilV���d�kv��Q���댻ݺ��J��m���fy���3������i3��s㈻�̇�X���0���s[�����Z>���7��Rx��if�����9�����.k��붦�X/��F��M���n"���9ƻ�=ϻ �ջ�  �  ���<e��<��<�f�<89�<.��<���<���<�O�<Fs�<�X�<M=�<wa�<���<|!�<���<o2�<���<2��<e��<�B�<�U�<���<���<:��<���<l��<6�<��<Ͼ�<��<���<���<"y�<���<^�<�P�<ϱ�<u��<e��<�=�<E:�<���<�A�<��<)%�<��<u�<�A�<�h�<� �<�4�<�>�<�\�<���<���<�<�<�R�<���<;��<���<	��<�	�<q��<��<�a�<�8�<���<�^�<�Q�<]��<N��<�G�<���<���<E��<y:�<��<���<{R�<Iy�<c��<�k�<���<�ҳ<'��<���<���<f��<"o�<�9�<kZ�<��<��<b/�<�\�<��<��<�<���<Dq�<>s�<E��<5w�<�<*�<B{�<X�<i�}<�uv<��o<�$j<N�e<}�b<�w`<��^<۲\<��Y<�U<�%P<�ZI<�A<�:<��2<�,<�(<f�$<��"<��!<H <1+<j�<�<�<[	<�Z<� �;FR�;z%�;!�;:y�;��;^�;`��;+ְ;��;���;v��;�r�;o�;I�j;]�M;��3;�/;;;��;���:JF�:�W�:���:�q�:��{:�:��T9��3��& ���<�~�^�f�g��]��}I���7��L2���>��@^����i���2;ĺ�*����Dj�����M�!��ø�/@�	к'�ź�IĺAͺd�������8�@S�]�%�#+��+�+9&������i$�a�����G��&,���;�y�J�,V�.�\�N�]���Y���R�`�J�&aE��ED� rH��Q��_�xo����(���X�Eʑ��r���Ӓ�[��hΌ��+��k��fk��IɆ�͊��?���U���š�B#���Y���ڰ������a����������|���p��%$��
[��@�������Ȼbλ�  �  ;;�<�;�<b��< �<݄�<C��<��<i#�<���<��<+K�<��<���<Z��<"��<���<S��<� �<���<�I�<���<���<0j�<
��<<�<՗�<���<f�<�O�<��<ě�<���<5;�<#��<���<��<�5�<���<;��</*�<��<^�<�0�<�x�<�<ź�<N.�<s7�<)��<I��<��<2��<}M�<���<<v�<��<��<��<S�<��<z��<�#�<p�<�Q�<���<�u�<���<��<C��<D��<���<��<���<���<���<G��<���<���<~��<$��<Sb�<�+�<�K�<'�<1�<c��<`��<�\�<h�<��<{��<뽩<bv�<��<V�<�֛<���<�Õ<�Y�<�_�<�ȏ<�u�<m>�<���<�x�<���<�Y�<О�<Ӈ�<d�z<St<R�n<��i<f</�b</`<�]<�xY<6U<P�O<��I<��B<�@<<�6<��0<]�,<`W)<9�&<o%<��"<��<$�<H�<��<�R
<kD<gT�;ѿ�;�g�;>��;e��;�X�;�o�;�\�;zv�;m�;ǎ�;y�;L��;b͉;�y;�-_;@F;�^0;UA;��;�	;� �:���:f�:-j�:��y:��%:(v�9񥗶򀊹�s�/���( �Q����-Y��x��m.��P���}�)����,����˺��ߺ���3����E�캗$���ӺƙǺ���O���������κ`8������	�Ʉ����o-�����������W�n���<�ɕ(�� 4�,�>��F���J�@K�3`H�+�C��F?�uJ=��	?�^�D��JN�R�Z�PYh�fv�����Sֆ�hn��DB���a��q��'ވ�t��ވ������🄻s��#C������=���p&��~H�������Щ�����nV��@���'�������꫻ϰ�0Ƕ�V�T»�/ƻ�  �  �E�<yB�<�d�<��<�f�<���<-�<M�<���<�f�<}��<N��<~u�<`�<���<?W�<�#�<�&�<�M�<���<��<���<��<7�<�:�<>�<���<�r�<S�<sx�<���<��<�d�<A4�<���<�i�<i��<U��<�<T8�<���<�I�<f@�<}q�<s��<h��<��<���<'��<��<ۜ�<a]�<"�<:�<��<�T�<���<��<���<��<��<4B�<Mc�<�L�<u��<A�<���<'@�<:n�<s��<u��<z+�<k��<$>�<���<N�<�&�<��<Lj�<`��<���<tU�<��<�Թ<�	�<�x�<n��<w[�<�q�<�+�<t��<ٯ�<���<}t�<cI�<�3�<�G�<S��<J�<��<���<�9�<���<d�<�v�<+��<<B{�<�<�"~<�dx<�r<�m<[
i<X�d<�`<$�\<�\X<I�S<��N<
I<bhC<~�=<a�8<�M4<��0<XO-<�*<_�'<�$<g� <�<��<K
<��
<L�<���;���;���;��;��;�E�;���;��;V��;7Z�;���;cP�;T֗;�;���;�n;�W;��@;ߦ,;Џ;DS
;�j�:���:�l�:��:��k:$%:���9�i9�����@b�]ǣ������ι�ܹ�I�����NC-��~Q�s�y�����ڼ��e����Lƺ�к�a׺J�ٺ[�׺�Ӻ:o̺pźH�����������pBĺE�к^���T��'�X9
�3@��$�4m�Q�9�������!�
�'��.���4���8��:�X�:�\=9�j7�2�6��8�.�=��E��cN��X�$�c���n�J7x�Z���.���8���B��*j��!셻|���M��C�_������􈻣R��_�����������c���P˥�_񦻏��L���U���*������Y����z��7����⾻�  �  ���<Ϋ�<х�<�-�<��</��< ��<�^�<�7�<,&�<�2�<^�<���<d��<�T�<��<�8�<5��<�h�<M-�<�<>�<9��<���<�~�<d��<]��<9��<��<,��<ű�<B��<
�<�l�<��<L�<b��<�_�<��<��<C��<���<���<���<̺�<�r�<���<��<��<��<��<�A�<Ȅ�<z��<
V�<��<+_�<-��<l��<P5�<���<���<���<m��<yb�<��<UC�<�&�<,��<���<�!�<2�<�8�<M:�<�2�<��<���<S��<���<�D�<��<|��<��<0�<rl�<]��<*��<���<'5�<���<h˫<���<P2�<�x�<;Ѡ<�7�<�<��<���<�%�<�Ƒ<W��<r�<���<>ȉ<��<�m�<���<���<O/�<R9{<��u<*_p<|�j<��e<�x`<�a[<�WV<!YQ<�iL<��G<��B<}�><�|:<j�6<IW3<b0<[�,<��(<��$<U�<��<V<��<n
<<;��;��;c��;|y�;ʎ�;���;'��;꾻;��;��;��;G�;2�;NY�;�a�;�x;?c;Z�L;��6;Q!;��;�I�:��:�C�:zy�:�O:Tq:o�9&gT9`o�8��6�����P��>��#������!^��B�-�g�����D���f��?Y������bø�����;]ĺD�ȺA�˺Kͺ�̺�ʺ �ǺOwźpź߂ɺ�jҺ�Yߺ}�`'������4�������b��o �4$���'��*�!+-��.�uy/�s/��&/��F/�t�0��C4��8:�V
B���J���S��\���c��j�v�o��0u��z���~��l��K��Ԅ��ꅻ͉���І�����do�������ي��F�������1��ԛ�U*��p���v�����#C���ԯ�<��Ws���f��������������  �  O; =_% =���<K �<��<�}�<l�<���<%��<8G�<i��<���<�V�<���<�s�<��<F��<���<���<%4�<���<
��< ��<���<���<<��<�X�<?��<�|�<C:�<��<��<XF�<G2�<~Y�<��<fp�<�\�<�}�<���<.�<NS�<�p�<lQ�<���<
�<��<b��<w��<H��<	��<��<B]�<I�<6,�<j��<�w�< ��<���<��<�J�<���<vA�<��<��<�	�<���<=5�<�$�<���<���<��<E.�<B��<�(�<���<�Z�<<+�<�(�<�R�<���<n	�<�u�<Tһ<��<��<���<R�<�!�<(�<�D�<"��<�!�<Z�<\Ӡ<�<N��<�:�<��<��<N�<�G�<橌<'X�<x^�<���<�F�<��<�U�<�w�<�v|<.Sw<��q<h�k<�ce<�-_<&Y<�uS<w5N<$tI<6E<�sA<
><)�:<c�7<˲4<�21<\2-<\�(<�I#<�<C�<�b<O<��<�u<k <T��;>��;c+�;��;��;�;�;�/�;K�;��;`��;�;�6�;�A�;�a�;�<|;��h;�S;=�;;)5#;��
;0=�:��:mQ�:�u_:�t%:�:�9(�9�'W98��8wF48� �^a����Ϲ�t�)E��p��I���閺�a��鴡��٢�!��3K��|N���G���q���Gͺ9�׺�޺Q��@ߺ�/ں�!Ժ{кg�к�Q׺\+㺴7� �1�����6��z'�ަ,�h90���1��1��
0�L�-�b+���)��)�=�+�k�0�$�8��]B�*�L�l�V��^��/d�i�g���i��kk���m�fq�!6v�l�|��)����//���w��V�������1�����1ˋ�yC��r*��ZK���S���㞻����	���ꮻ�󲻩 �����{
���1������ ��Y���  �  �@ =� =b�<�<^q�<���<��<���<�$�<_��<D�<�U�<ܕ�<��<( �<|?�<���<D|�<���<}��<9��<}�<���<��<v��<���<{��<)��<��<�(�<"��<K��<b�<��<��<���<���<\ �<��<�9�<:��<�W�<�u�<0 �<wK�<��<Jt�<��<��<_��<�F�<>W�<���<5�<���<��<��<9�<���<҆�<�!�<� �<G�<8 �<��<0g�<��<��<M��<&��<=��<�[�<H��<Դ�<2��<���<�y�<(O�<��<4�<���<���<�J�<�ʻ<��<���<3�<���<�b�<"�<�(�<`��<ь�<O١<�Z�<�՞<1�<��<9E�<;;�<��<Պ�<_�<���<�b�<���<�w�<qv�<f�<��<�@|<�ow<%�q<�"k<I(d<.]<~?V<��O<ކJ<�E<7/B<{.?<B�<<�I:<ż7<�4<�0<4=,<�&<k <��<��<�J<1�	<��<��<���;��;�@�;��;��;q�;���;���;�[�;��;���;R�;���;hP�;�l�;M�y;��h;��S;ux;;� ;	;�:�!�:�m:':GK�9��9-T9�39I��8�hR8���.�b���v	�>�F�Ľ���#��B˩�<���厱��ȫ����������ܢ�v���x���kֺ��麽���P: �U ��"��#��H�vۺ!�ں�㺽��0�y��2���5*�Q04�/;�my>��r>�w;���6�h�0��!,��r)�/�)��L.�Ķ6�BxB�^�O�ٺ\��g���m�R�p���o��_m���j�l�i�Y�k�;mq��qz�������r|��s�������ꔻ"����r��ө��A7��%����%��u]���ߟ�7���9������u͹��D�����򾻘����f��!���t���  �  [
 =���<�{�<��<Q��<k��<>��<���<q�<�A�<I��<��<�x�<���<�l�<�f�<]��<e��<2��<���<f��<�7�<A[�<��<���<���<!.�<���<��<���<d��<u��<���<�<H��<f�<g�<���<�b�<�f�<S�<���<� �<it�<�B�<��<���<ٷ�<�G�<x�<c[�<���<���<���<ُ�<���<Wb�<@E�< ��<á�<���<P�<��<̲�<q��<w�<��<wi�<J�<��<�A�<H��<��<t��<�B�<8�<���<m�<���<���<ʣ�<�Ľ<g��<_Q�<�^�<�Ͷ<���<��<�Y�<�٨<�֥<�u�<���<��<��<��<�-�<�0�<y��<x-�<jg�<��<�Љ<���<t.�<�v�<�b�<���<z�<�,~<o{<ǚv<��p<��i<�_b<]�Z<)'S<�sL<n�F<�RB<%�><`�<<�:<[�8<��6<K�3<�/<�^*<��#<x�<��<�6<�	<L�<ب<9� <H��;�Z�;�5�;�j�;��;��;�h�;{�;z��;�;㿎;���;Ƶ�;��;7~};x�s;�e;�P;S8;h�;��: [�:Ո:�Q5:AI�9�o9��8�*�8��R8 o"8�N6j���/m�t��7��逺���o���̺�2к�ɺպ�����i����ɘ��d�������tǺg���V �`����c����.�:���K캅>溼�꺑l��:{��*��&��5���A�P�I���L���K�!vF���>���6��0�ڿ,�5�-�T�4�m@��UO���_��n��Iy���~��~��ez�݀s��l��h��ji�!�o�~�z����$J���Ԕ�<�������������$����#���������ᕻ���)O������8$��Ժ�����ĻKƻ9Ż��»���V���NA���  �  �y�<i��<py�<�o�<�
�<]��<���<c��<EC�<���<���<��<t,�<��<�|�<�T�<|e�<��< ��<UZ�<���</�<\W�<�+�<�]�<l��<�<�<�E�<��<��<��<���<4��<M��<w<�<���<��<�4�<wJ�<���<#��<�T�<�]�<���<�%�<��<T��<���<<�<~�<���<�q�<���<�;�<_�<���<=l�<[�<��<��< R�<�`�<"�<��<"��<d��<���<x<�<C=�<�b�<Ơ�</�<Z��<�i�<6��<���<���<���<�I�<sD�<���<��<N�<��<���<Vٵ<&b�<.y�<�{�<�Ϧ<�ã<G��<�
�<�4�<"��<��<8�<N?�<P��<��<�Ő</n�<�U�<�ل<�3�<Gs�<�~<~<�i}<� |<�y<gu<¡o<��h<,�`<�OX<jP<�gI<�C<?<?<�+<<.:<��8<�l7<�}5<��2<�!.<3M(<�?!<p�<��<N<�<��<�$�;���;$��;�<�;9�;M��;��;�~�;�l�;�)�;�a�;2_�;fІ;컀;��z;�}w;�s;��l;r�_;�}L;�R3;��;���:OT�:�Je:�
:�qr9"zV81J)�݄��jU�8�'�T9���T"�ȩ�Ǧ�I<e�훜�N@º��ݺ�B�\=�a�ߺ��ʺ�U�������D��毝�����Ϻ���jQ�1�bO!��"����b�F	�b���c�����j����]��Eu/��@�O�M�}7V��dY��*W�ssP���F�t=��+5��w1�px3�O�;���I���[�Bhn���~�x̄�����	��S���?z�zp��}i���h�7�o�X}����]���Cؚ��Ρ�񪥻*������Q\�����S)���2��8U���j%���E������PG���ƻ2�ʻ�$̻��ʻTǻQ�»w���i����  �  ���<�B�<���<�u�<���<<`�<ke�< 9�<���<@��<��<i~�<���<���<�t�<�4�<V�<;]�<���<�5�<{��<%��<g��<��<E<�<���<��<(��<m�<2��<�v�<3�<���<A��<"4�<Q��<���<�L�<e��<���<P�<��<N��<��<{O�<p�<G��<g�<��<�!�<�]�<:m�<��<���<�)�<���<�`�<[��<��<~��<�S�<y)�<���<�:�<7��<�i�<��<�[�<��<��<t�<���<�=�<���<5��<��<���<��<�G�<�]�<�ͼ<�J�<X��<�(�<��<,�<5s�<�V�<N.�<4h�<bX�<�)�<f۞<�A�<��<���<��<�6�<�o�<ﭔ<�B�<ա�<�G�<Й�<7׀<."~<aV|<��{<dq{<��z<pYx<�et<(�n<�lg<�6_<�V<��N<�[G<��A<E*=<%A:<w~8<�a7<�A6<�v4<xt1<��,<�&<�C<B&<�;<�O<]�<
��;���;�C�;?��;�%�;���;q��;3N�;:?�;��; ��;Q�;@�;�\�;��v;��p;5�n;;�l;��f;�Q[;��H;pw/;�,;�x�:��:;G:�\�9w��81��������#��9���׸� �*�c���ҹ`	0����C��]�׺�F���� ��������׈ֺ����M飺r��k]��
��kֺ���9�5�"�e,���-�h�(�gU���	6�}�������=Q����"���5��GG�]U��^���a�I�^�'eW��L�k�A��B9�,e5��7�fA�2 Q�*�d�H�x��˄��c���^��*������uy�hs�s�j��5i�
=p��"�����n唻U���ަ��,��*ë���X ������V��Z����a��zz��]������W���;Ļ��ʻ�ϻ�;л��λ��ʻ�Żp���z����  �  ���<7�<�i�<c�<{r�<���<���<���<Ņ�<9�<���<=H�<J��<4��<�n�<[&�<J��<P!�<fD�<7��<��<�K�<�v�<�j�<���<?�<�;�<�y�<���<M\�<�=�<���<;]�<�K�<���<>$�<b6�<���<�9�<��<���<��<���<^��<���<X��<�*�<���<
V�<Z��</��<��<z��<֗�<Q�<���<(Y�<9��<�{�<ű�<B��<	��<vF�<���<5	�<���<��<��< I�<ڛ�<@��<,M�<���<T�<��<�O�<���<�a�<w�<G�<(��<��<M�<d��<�ѷ<մ<f�<��<F��<��<�ס<��<n�<t�<�ȝ<��<yܜ<a0�<�e�<���<0�<OV�<��<q'�<�[�<1'}<�e{<�z<J�z<*�y<��w<�t< Jn<g<Z�^<�V<��M</�F<��@<�p<<M�9<Y�7<H�6<��5<�4<C1<i,<6"&<e�<�K<�H<Q<q�<U��;/�;#�;"��;���;���;���;l�;��;,�;�f�;YV�;�l�;��~;��r;G9m;gzk;��i;
�d;)�Y;�CG;� .;�s;�a�:$?�:�n<:]��9���8e_�PCD��3G�i#��������^}�BK�6�9�� ����rߺ�-��{���j�\�����ں[~���G������_Ξ�G��5ٺ��D�(S&�r�/���1�Ǧ,�d�!�u������X��~ ������_�$�b�7��I��KX�lva�.�d�5�a��Y�,�N�߮C�w�:���6�[�9��C���S���g� F|�]���8^���A��Va��j�������=t��%k�hi�c�p��������?��,���筨�c ������J򪻈֥���Ѕ��Z���V,���:���3��9���%���SŻi_̻Îл-�ѻ�ϻ	�˻,�ƻ����oh���  �  ���<�B�<���<�u�<���<<`�<ke�< 9�<���<@��<��<i~�<���<���<�t�<�4�<V�<;]�<���<�5�<{��<%��<g��<��<E<�<���<��<(��<m�<2��<�v�<3�<���<A��<"4�<Q��<���<�L�<e��<���<P�<��<N��<��<{O�<p�<G��<g�<��<�!�<�]�<:m�<��<���<�)�<���<�`�<[��<��<~��<�S�<y)�<���<�:�<7��<�i�<��<�[�<��<��<u�<���<�=�< ��<7��<��<���<��<�G�<�]�<�ͼ<�J�<]��<�(�<��<2�<<s�<�V�<T.�<:h�<hX�<�)�<k۞<�A�<��<���<��<�6�<�o�<�<�B�<ѡ�<�G�<̙�<2׀<#"~<UV|<��{<Xq{<��z<eYx<�et<�n<�lg<�6_<�V<��N<�[G<��A<G*=<(A:<|~8<�a7<�A6<�v4<�t1<��,<�&<�C<N&<�;<�O<h�<��;���;�C�;I��;�%�;���;q��;/N�;3?�;��;�;@�;@�;�\�;X�v;��p;�n;�l;_�f;�Q[;e�H;Ew/;�,;�x�:e�:�G:6\�9*��8������v�#��9� �׸2� �K�c���ҹd	0����D��]�׺�F���� ��������׈ֺ����L飺r��k]��
��kֺ���9�5�"�e,���-�h�(�gU���	6�}�������=Q����"���5��GG�\U��^���a�I�^�'eW��L�k�A��B9�,e5��7�fA�2 Q�*�d�H�x��˄��c���^��*������uy�hs�s�j��5i�
=p��"�����n唻U���ަ��,��*ë���X ������V��Z����a��zz��]������W���;Ļ��ʻ�ϻ�;л��λ��ʻ�Żp���z����  �  �y�<i��<py�<�o�<�
�<]��<���<c��<EC�<���<���<��<t,�<��<�|�<�T�<|e�<��< ��<UZ�<���</�<\W�<�+�<�]�<l��<�<�<�E�<��<��<��<���<4��<M��<w<�<���<��<�4�<wJ�<���<#��<�T�<�]�<���<�%�<��<T��<���<<�<~�<���<�q�<���<�;�<_�<���<=l�<[�<��<��< R�<�`�<"�<��<"��<d��<���<x<�<C=�<�b�<Ǡ�<0�<\��<�i�<8��<���<���<���<�I�<zD�<���<��<X�<��<���<aٵ<2b�<:y�<�{�<�Ϧ<�ã<P��<�
�<�4�<(��<��<:�<N?�<O��<��<�Ő<(n�<�U�<�ل<�3�<<s�<�~<�~<�i}<� |<ˑy<jgu<��o<��h<�`<�OX<jP<�gI<�C<B<?<�+<<
.:<��8<�l7<�}5<��2<�!.<JM(<�?!<��<��<d<�<��<%�;���;9��;�<�;$9�;M��;���;�~�;�l�;�)�;�a�;_�;<І;���;i�z;P}w;��s;W�l;�_;�}L;@R3;E�;"��:�S�:-Je:�	:�or9sV8�O)�߄��mU�X�'�:��U"�ȩ�ͦ�M<e��O@º��ݺ�B�\=�a�ߺ��ʺ�U�������D��毝�����Ϻ���jQ�1�bO!��"����b�F	�b���c�����j����]��Eu/��@�O�M�}7V��dY��*W�ssP���F�t=��+5��w1�px3�O�;���I���[�Bhn���~�x̄�����	��S���?z�zp��}i���h�7�o�X}����]���Cؚ��Ρ�񪥻*������Q\�����S)���2��8U���j%���E������PG���ƻ2�ʻ�$̻��ʻTǻQ�»w���i����  �  [
 =���<�{�<��<Q��<k��<>��<���<q�<�A�<I��<��<�x�<���<�l�<�f�<]��<e��<2��<���<f��<�7�<A[�<��<���<���<!.�<���<��<���<d��<u��<���<�<H��<f�<g�<���<�b�<�f�<S�<���<� �<it�<�B�<��<���<ٷ�<�G�<x�<c[�<���<���<���<ُ�<���<Wb�<@E�< ��<á�<���<P�<��<̲�<q��<w�<��<xi�<J�<��<�A�<J��<��<w��<�B�<8�<���<#m�<���<ȑ�<֣�<Ž<v��<nQ�<�^�<�Ͷ<ɥ�<��<Z�<�٨<�֥<�u�<���<��<��<��<�-�<�0�<w��<t-�<dg�<��<�Љ<���<e.�<�v�<�b�<���<i�<�,~<O{<��v<��p<��i<�_b<M�Z<'S<�sL<l�F<�RB<.�><n�<<'�:<q�8<��6<g�3<�/<�^*<��#<��<ݼ<�6< �	<g�<�<L� <f��;�Z�;�5�;�j�;��; ��;�h�;U�;L��;�;���;p��;���;q�;�}};��s;Te;��P;�8;��;O��:UZ�:�Ԉ:Q5:�G�9��o9���8�'�8C�R8l"8��M6$���C/m�3t��7��逺���o���̺�2к�ɺպ�����i����ɘ��d�������tǺg���V �`����c����.�:���K캅>溼�꺑l��:{��*��&��5���A�P�I���L���K�!vF���>���6��0�ڿ,�5�-�T�4�m@��UO���_��n��Iy���~��~��ez�݀s��l��h��ji�!�o�~�z����$J���Ԕ�<�������������$����#���������ᕻ���)O������8$��Ժ�����ĻKƻ9Ż��»���V���NA���  �  �@ =� =b�<�<^q�<���<��<���<�$�<_��<D�<�U�<ܕ�<��<( �<|?�<���<D|�<���<}��<9��<}�<���<��<v��<���<{��<)��<��<�(�<"��<K��<b�<��<��<���<���<\ �<��<�9�<:��<�W�<�u�<0 �<wK�<��<Jt�<��<��<_��<�F�<>W�<���<5�<���<��<��<9�<���<҆�<�!�<� �<G�<8 �<��<0g�<��<��<M��<'��<>��<�[�<J��<״�<7��<���<�y�<1O�<��<A�<���<���<�J�<�ʻ<��<Σ�<H�<¹�<�b�<5�<�(�<p��<ߌ�<[١<�Z�<�՞<5�<��<7E�<6;�<��<ʊ�<_�<���<�b�<{��<�w�<]v�<�e�<��<�@|<�ow<�q<�"k<1(d<]<p?V<��O<܆J<�E<B/B<�.?<X�<<�I:<�7<�4<+�0<\=,<F�&<Hk <��<��<�J<Q�	<�<��<���;��;�@�;��;��;�p�;���;T��;i[�;��;���;�Q�;H��;P�;4l�;��y;�h;�S;�w;;�� ;�;L�:� �:ߧm:�':�I�9x�9C+T9�29d��8�eR8����.�z���v	�B�F�Ž���#��B˩�;���厱��ȫ����������ܢ�v���x���kֺ��麽���P: �U ��"��#��H�vۺ!�ں�㺽��0�y��2���5*�Q04�/;�my>��r>�w;���6�h�0��!,��r)�/�)��L.�Ķ6�BxB�^�O�ٺ\��g���m�R�p���o��_m���j�l�i�Y�k�;mq��qz�������r|��s�������ꔻ"����r��ө��A7��%����%��u]���ߟ�7���9������u͹��D�����򾻘����f��!���t���  �  O; =_% =���<K �<��<�}�<l�<���<%��<8G�<i��<���<�V�<���<�s�<��<F��<���<���<%4�<���<
��< ��<���<���<<��<�X�<?��<�|�<C:�<��<��<XF�<G2�<~Y�<��<fp�<�\�<�}�<���<.�<NS�<�p�<lQ�<���<
�<��<b��<w��<H��<	��<��<B]�<I�<6,�<j��<�w�< ��<���<��<�J�<���<vA�<��<��<�	�<���<>5�<�$�<���<���<��<H.�<F��<�(�<���<�Z�<F+�<�(�<S�<���<�	�<�u�<iһ<��<��<خ�<i�<�!�<(�<�D�<5��<"�<h�<gӠ<�<R��<�:�< ��<��<E�<�G�<ש�<X�<e^�<���<xF�<��<�U�<�w�<xv|<Sw<��q<H�k<�ce<~-_< &Y<�uS<u5N<*tI<6E<�sA<#><H�:<��7<�4<�21<�2-<��(<�I#<�<n�< c<*O<��<�u<k <p��;L��;c+�;���;Ԙ�;�;�;�/�;�;j�;��;��;96�;4A�;�a�;/<|;��h;S;��;;�4#;+�
;G<�:��:�P�:vt_:t%:89�9'�9v&W9��8tC48#�h �za����Ϲ�t�+E��p��I���閺�a��贡��٢�!��3K��{N���G���q���Gͺ9�׺�޺Q��@ߺ�/ں�!Ժ{кg�к�Q׺\+㺴7� �1�����6��z'�ަ,�h90���1��1��
0�L�-�b+���)��)�=�+�k�0�$�8��]B�*�L�l�V��^��/d�i�g���i��kk���m�fq�!6v�l�|��)����//���w��V�������1�����1ˋ�yC��r*��ZK���S���㞻����	���ꮻ�󲻩 �����{
���1������ ��Y���  �  ���<Ϋ�<х�<�-�<��</��< ��<�^�<�7�<,&�<�2�<^�<���<d��<�T�<��<�8�<5��<�h�<M-�<�<>�<9��<���<�~�<d��<]��<9��<��<,��<ű�<B��<
�<�l�<��<L�<b��<�_�<��<��<C��<���<���<���<̺�<�r�<���<��<��<��<��<�A�<Ȅ�<z��<
V�<��<+_�<-��<l��<P5�<���<���<���<n��<zb�<��<UC�<�&�<,��<���<�!�<2�<�8�<Q:�<�2�<��<���<]��<���<�D�<��<���<��<+0�<�l�<u��<B��<��<>5�<ʐ�<}˫<���<a2�<�x�<FѠ<�7�<���<��<���<�%�<�Ƒ<J��<r�<퉋<*ȉ<t�<nm�<���<���<8/�<%9{<��u<_p<Z�j<��e<�x`<va[<�WV<YQ<�iL<��G<��B<��><}:<��6<rW3<�0<��,<*�(<�$<��<��<8V<��<;n
<3<d��;��;r��;}y�;���;���;���;���;ٚ�;9�;{�;�F�;�1�;�X�;�a�;)�x;�c;��L;W�6;�P!;�;�H�:?��:C�:�x�:)�O:�p:a�9�eT9m�8֭6�P��LP��>��5�����$^��B�-�g�����D���f��?Y������bø�����;]ĺD�ȺA�˺Kͺ�̺�ʺ �ǺOwźpź߂ɺ�jҺ�Yߺ}�`'������4�������b��o �4$���'��*�!+-��.�uy/�s/��&/��F/�t�0��C4��8:�V
B���J���S��\���c��j�v�o��0u��z���~��l��K��Ԅ��ꅻ͉���І�����do�������ي��F�������1��ԛ�U*��p���v�����#C���ԯ�<��Ws���f��������������  �  �E�<yB�<�d�<��<�f�<���<-�<M�<���<�f�<}��<N��<~u�<`�<���<?W�<�#�<�&�<�M�<���<��<���<��<7�<�:�<>�<���<�r�<S�<sx�<���<��<�d�<A4�<���<�i�<i��<U��<�<T8�<���<�I�<f@�<}q�<s��<h��<��<���<'��<��<ۜ�<a]�<"�<:�<��<�T�<���<��<���<��<��<4B�<Mc�<�L�<u��<A�<���<'@�<:n�<t��<v��<}+�<n��<)>�<���<T�<�&�<��<Xj�<n��<��<�U�< �<�Թ<�	�<�x�<���<�[�<�q�<�+�<���<쯩<���<�t�<mI�<�3�<�G�<T��<H�<��<~��<x9�<���<S�<�v�<��<���<,{�<��<�"~<fdx<��r<�m<;
i<<�d<ν`<�\<�\X<H�S<��N<�
I<uhC<��=<�8<�M4<��0<�O-<�*<��'<K�$<�� < <��<o
<�
<f�<���;��;���;��;���;�E�;���;��;��;�Y�;N��;P�;�՗;��;g��;Pn;@W;,�@;>�,;=�;�R
;�i�:��:�k�:���:��k:`#%:���96h9�����Ab��ǣ����ι�ܹ�I�����OC-��~Q�r�y�����ڼ��e����Lƺ�к�a׺I�ٺ[�׺�Ӻ:o̺pźH�����������pBĺE�к^���T��'�X9
�3@��$�4m�Q�9�������!�
�'��.���4���8��:�X�:�\=9�j7�2�6��8�.�=��E��cN��X�$�c���n�J7x�Z���.���8���B��*j��!셻|���M��C�_������􈻣R��_�����������c���P˥�_񦻏��L���U���*������Y����z��7����⾻�  �  ;;�<�;�<b��< �<݄�<C��<��<i#�<���<��<+K�<��<���<Z��<"��<���<S��<� �<���<�I�<���<���<0j�<
��<<�<՗�<���<f�<�O�<��<ě�<���<5;�<#��<���<��<�5�<���<;��</*�<��<^�<�0�<�x�<�<ź�<N.�<s7�<)��<I��<��<2��<}M�<���<<v�<��<��<��<S�<��<z��<�#�<p�<�Q�<���<�u�<���<��<D��<E��<���<��<���<���<���<M��<���<���<���<1��<bb�<�+�<�K�<:�<E�<w��<u��<�\�<}�<��<���<���<pv�<��<
V�<�֛<���<�Õ<�Y�<�_�<�ȏ<�u�<_>�<���<�x�<���<�Y�<���<���<<�z<�Rt<.�n<v�i<�f<�b<`<�]<�xY<5U<U�O<��I<��B<�@<<6<��0<��,<�W)<a�&<�%<��"<�<J�<l�<��<�R
<�D<�T�;��;�g�;>��;Y��;�X�;go�;h\�;Bv�;,�;���;�x�;���;͉;6�y;�,_;`?F;^0;�@;I�;
	;���:%��:oe�:�i�:ĕy:��%:<u�9�ї�q���t�N���( �_���2Y��x��m.��P���}�)����,����˺��ߺ���3����E�캗$���ӺƙǺ���O���������κ_8������	�Ʉ����o-�����������W�n���<�ɕ(�� 4�,�>��F���J�@K�3`H�+�C��F?�uJ=��	?�^�D��JN�R�Z�PYh�fv�����Sֆ�hn��DB���a��q��'ވ�t��ވ������🄻s��#C������=���p&��~H�������Щ�����nV��@���'�������꫻ϰ�0Ƕ�V�T»�/ƻ�  �  ���<e��<��<�f�<89�<.��<���<���<�O�<Fs�<�X�<M=�<wa�<���<|!�<���<o2�<���<2��<e��<�B�<�U�<���<���<:��<���<l��<6�<��<Ͼ�<��<���<���<"y�<���<^�<�P�<ϱ�<u��<e��<�=�<E:�<���<�A�<��<)%�<��<u�<�A�<�h�<� �<�4�<�>�<�\�<���<���<�<�<�R�<���<;��<���<	��<�	�<q��<��<�a�<�8�<���<�^�<�Q�<^��<P��<�G�<���<���<J��<:�<��<���<�R�<Uy�<p��<�k�<���<�ҳ<8��<��<���<w��<2o�<�9�<xZ�<��<��<j/�<�\�<��<��<�<���<>q�<6s�<:��<(w�<�<�<2{�<�W�<G�}<suv<��o<�$j<2�e<e�b<�w`<�^<в\<��Y<�U<�%P<�ZI<#�A<�:<��2<�,<�(<��$<�"<ɢ!<>H <R+<��<�<�<r	<�Z<� �;ZR�;�%�;!�;0y�;��;�]�;:��;�հ;K�;d��;7��;rr�;*�;��j;��M;,�3;B/;�;v�;3��:�E�:W�:��:�q�:�{:k�:y�T9��3��& ��<���^�w�g�#�]��}I���7��L2���>��@^����i���2;ĺ�*����Cj�����M�!��ø�/@�	к'�ź�IĺAͺd�������8�@S�]�%�#+��+�+9&������i$�a�����G��&,���;�y�J�,V�.�\�N�]���Y���R�`�J�&aE��ED� rH��Q��_�xo����(���X�Eʑ��r���Ӓ�[��hΌ��+��k��fk��IɆ�͊��?���U���š�B#���Y���ڰ������a����������|���p��%$��
[��@�������Ȼbλ�  �  ��<���<դ�<}��<���<m��<���<��<��<���<�e�<��<���<�q�<��<Bb�<N��<���<���<��<K��<���<�<m��<}s�<��<Y��<��< �<a��< ��<4��<��<N;�<M��<pl�<�4�<�@�<J��<h��<o��<+L�<u��<]B�<�H�<���<��<���<=��<9��<
]�<�g�<�7�<x�<[�<.�<���<>��<��<���<���<2��<#v�<k6�<��<<�<=��<g�<�j�<O�<f��<#�<4��<��<��<r��<#S�<��<T��<'��<���<�W�<���<�ѳ<�ұ<(��<��<���<X�<e��<a��<Tʨ<�C�<�E�</�<�<g�<�[�<� �<zS�<7�<�t�<���<�Ҋ<Xg�<�P�<��<�
�<�ez<�r<޶k<�f<1�a<>n_<y
^<�*]<��[<ܾY<v�U<A P<~�H<�_@<��7<�/<)<~$<i� <Y3<}h<�<�8<�c<��<g�<��<���;ZV�;��;���;��;�N�;�y�;a��;:ٰ;`٭;k��;��;?p�;�	�;d�|;�\;B>;L#;~�;���:���:K+�:���:��:U*�:Pަ:^w:M�:���8����c�6��1{��r���@��� ���{���^�fXO�Z�T�Baq�{h�����O�Ժ,h��p��&��5=�
�o�����r�y}ں�*Ϻ��κ�ۺ�9��	���2+�3"6�A�:���8�1�&�%����$C�ܵ�6R�����0� �C�XV��<d��el���m��6i��\`��7V��"N���J�U{M�ilV���d�kv��Q���댻ݺ��J��m���fy���3������i3��s㈻�̇�X���0���s[�����Z>���7��Rx��if�����9�����.k��붦�X/��F��M���n"���9ƻ�=ϻ �ջ�  �  ��<	��<rT�<���<���<c��<�0�<H��<�4�<M$�<z��<w8�< 
�<Lk�</��<_�<Z��<���<E�<�q�<�,�<|3�<a�<V��<�p�<���<�}�<4��<���<���<���<v��<��<���<R��<�c�<M�<G��<�7�<��<c�<��<Hx�<	��<��<���<��<���<��<U�<~��<,��<�y�<�:�<p`�<�$�<|��<���<���<��<�^�<%w�<��<$��<�s�<`�<R��<���<�<���<��<B��<�<Dk�<»�<[~�<�P�<E��<���<�Z�<Nǽ<rX�<]|�<|�<s�<qO�<LѮ<}��<j�<|�<�<�Q�<ٽ�<R��<�P�<)#�<�f�<OP�<2��<\�<�[�<R��<�(�<�N�<�<���<ݽ�<,�<rx<-p<��h<6Ac<>[_<u(]<�B\<��[<Z[<�Y<��U<��O<�5H<�D?< 6<c�-<��&<U[!<�$<O�<c<�<��<t6<��<C�<�f<\�;���;���;p��;=y�;�*�;%��;_U�;��;~��;�q�;"��;�ϖ;��;vNt;�S;�3;"�;
�;|?�:�b�:��:�J�:o��:���:1�:��q:���9�+77��Դ\��$��1���z��󝠺+H��{�ff��f��������0N��`���8����S.�ڔ�e��� �����k����⺽�ֺe�׺��� ����I�%�h$6��WA��|E��HB�T�8�ы+��������Z��1�!�@�4�HJ��X^�8%n�Pw�xy�xt��j��y^�M�T��O�`�Q��TZ���h�zD{��y����������<��[���$P��3�������͈���劻�ɉ�M���ט�����P��Iq���ƶ��	��U���	���3Ƕ�A���긪��-���M������ѳ��k��&�ɻʫӻ��ڻ�  �  z =q��<� =�M =� =_� =`K =�s�<���<���<�2�<=��<���<ZV�<�u�<hC�<��<��<���<��<.��<��<c��<r�<��<+��<�H�<���<��<��<�3�<���<P��<Ē�<��<s�<Z`�<$��<h��<7��<;�<��<��<���<�-�<`��<�G�<�M�<v��<ۆ�<���<N��<�h�<�K�<���<"W�<���<���<,��<���<���<���<�w�<֋�<���<K��<���<յ�<��<���<}b�<n��<��<,��<O\�<���<�,�<���<3�<��<��<N.�<��<{/�<��<���<�o�<QR�<�<��<�~�<�N�<ۖ�<���<Lj�<x�<�<���<⭓<�<���<�7�<���<�׎<���<��<,؉<g�<��<#��<]1{<��u<u�q<)�n<��l<k<'i<yef<�bb<�\<�HV<��N<�0G<�	@<#�9<Q�4<yI1<��.<'�,<�l*<�{'<e#<��<�L<Ӫ<��<q��;�;L+�;vI�;6�;�o�;��;��;R��;��;��;���;��;-�;�ލ;�Ԁ;' j;2V;c�G;˶=;��6;�1;=N*;�( ;'N;#�:#�:�ٙ:Q�R:[8�9I�}9�^�8U��7��7'8��Y8��7|f��z���U���lB��������@bú�պ�sݺK#ں��ͺ�������ې��6��nCx�b7�����,x��B^��9�Ӻ��3>�ƪ�\����ҺR�ú�縺f��~�Ӻ��ﺧ���Z�jE"��)�\q,�E�*�4m&��!�����!�Pn(��N4�^1D��jV���h���y�*����ㇻjy���x���e��Y����x� 
q�X�l�C�l���q��{�tp���j��䖑�y敻S͗�aP�����𯑻���d4���$��������������B�������l���  �  �0 = =5 =Gq =E� =�� =�` =x��<=��<|��<�h�<]#�<�&�<Χ�<���<��<���<���<���<_��<��<�:�<��<=7�<���<&@�<��<o<�<b�<# �<Zj�<��<&��<̍�<���<�a�<�U�<l��<6��<c�<�z�<�f�<���<���<z�<��<̀�<u}�<D��<'��<���<���<��<���<���<���<o�<45�<v��<$��<��<���<���<���<��<��<]�<g �<o��<��<��<?��<�4�<���<�`�<5��<��<.��<��<o��<J��<�`�<A)�<K|�<�k�<��<���<�<J#�<�4�<⤯<Zt�<`��<���<"��<-��<�<�<�J�<���<�X�<�8�<�o�<HǏ<� �<9�<�@�<�
�<�L�<�0�<2��<��{<o�v<=xr<Mgo<�%m<�?k<)'i<�Jf<c=b<��\<NCV<��N<�}G<|@<�g:<D�5<M�1<@N/<�,-<&�*<��'<^�#<KF<b�<�<G�< ��;ƺ�;Yu�;&��;Fc�;���;��;p��;Y7�;��;���;�B�;���;W�;Y	�;V�;�l;�Y;�J;�v?;(�7;��1;01*;߶;�;؋�:[y�:w�:��X:T3:�,�9�+9oz8I,^8lٗ8eԦ8��2849r��m��n<�?���V��s����кhFغ�7պ]ɺѶ�l衺�E����I9s��z�ʖ��qQ�������κ��ߺyl�@���޺jHѺDEú~}�����q��GGԺ�ﺕ~�۶��  �qW'���)��<(�9$�8��+�G$ ��2'��3���B�I�T�og��w�nZ��o����1���G���X���0���kw���o��Wk��ak��kp���y��X���1���L��L�������@_��NP��2`�������g���l�����!�����������Ю��I���  �  �� =Q� =w� =\� =�� =�� =l� =| =0O�<�<�<��<=��<'��<-��<Ĵ�<�x�<]��<!��<�|�<�x�<C�<���<��<���<K��<(�<�y�<#�<�=�<���<X��<�o�<��<�x�<7��<g(�<u0�<{��<I$�<���<(�<8�<���<G��<FP�<���<E�<� �<mT�<�<�`�<�^�<I�<�U�<���<���<�<��<���<~�<Q�<�j�<Y�<� �<D��<;w�<���<���<���<~��<�}�<�n�<{��<2�<f�<�d�<a��<���<{��<��<
>�<Y��<L޾<�O�<aL�<�¸<}��<�>�<���<�<}�<�۬<X5�<�K�<�V�<���<�<�6�<'�<�2�<���<��<&L�<s�<zO�<p��<���< ��<n��<Yԁ<%�}<ax<^t<خp<  n<��k<,i<@�e<�a<�t\<�%V<�?O<�BH<,�A<��;<�A7</�3<R1<@�.<0,<��(<��$<�<+v<�<�-	<
c<��;B�;�Z�;Z�;V��;�;+K�;�7�;)��;�b�;�>�;'�;���;-M�;>��;��s;�`;4P;F(D;.�:;u�2;��);?:;�;�m�:���:&��:�Hh:I8:7�9pmy9H29��#9�@+9(�#9�?�8�Uq�� 8�%<ѹMQ+�lSo���a���_º�ɺ�?Ǻ����2���2������Vr�]e���j��›.����f��y���ѺR(ۺXsܺ��ֺ��̺��ºr���L����\ĺg�պ����\V��G��� ���"�b/!�V���W��]��F��#�ȿ/��?�&FP��a��q�Ϝ}��炻�����䃻�_���f{��Ys��Pl�#h���g��%l���t��L���Ɔ�U������0z��Yӓ�����꜐�7Ȏ�����T��_Ғ��O��v	��b
���Z���,���  �  F>=�,= A=�`=�l=~J=�� =�J =N��<���<���<���<m;�<���<J�<���<� �<9��<�W�<)�<4��<:8�<�%�<,��<��<h.�</��<Fk�<Br�<��<U��<0��<�<�B�<�.�<��<���<M��<`h�<r!�<"�<�Z�<r�<�)�<ȁ�<D��<��<y��<���<���<8�<q%�<�>�<ny�<��<���<f�<_�<���<�w�<nI�<��<]��<B��<�G�<K�<	��<w��<�<�1�<m��<�W�<VL�<�Z�<�V�<:�<�e�<0<�<���<���<P��<���<�ӿ<2w�<�<+��<ӟ�<�2�<Wz�< M�<㙰<j�<�ܩ<��<�Y�<���<�o�<���<�D�<�v�<�<, �<��<9�<b�<X�<�V�<���<�<M�<_�<.�z<2Dv<�cr<�o<�l<��h<O9e<��`<Ʊ[<��U<�O<X4I<EC<�><��9<#86<�m3<]�0<� .<zk*<F�%<6 <�<�u<�
<�<D%�;���;���;Vt�;���;���;@��;��;���;ͼ;0��;5�;j��;1��;Eъ;�v~;c�i;��X;n]J;�b>;Rr3;_+(;�E;x�;���:�]�:K�:�Q|:M�::��:^}�9�Ы9�7�9�'�9��9��I9��8~ݸ�r��<P��vP�������#��{����z��B���{��t��vay��&`�Y�R���T��f�^��V����!��CX����Ⱥ kͺA�̺�Ⱥ�úG,��Bºa�ʺ��ٺ���x� �[�
�1Q����n�T��v��x����N�9��"+���9���I��PY�l�g�Ms�c�z��K~���}�,�y�Qt��om�psg��c�3�b��Jf���m���w��偻����i$������m��H{���ُ��E��:{������G��옻�l��L�����㬻�  �  !�=��=��=��=��=�=�3=l� =���<���<��<�4�<#��<~~�<���<�]�<l�<��<&L�<5��<�i�<���<���<�V�<��<�a�<)�<���< ��<���<<q�<�+�<'�<A��<̈�<8
�<	V�<�x�<���<˪�<���<-��<Sh�<ވ�<���< ��<���<"]�<!v�<�/�<"��<T��<)V�<���<��<���<S�<,��<��<2��<*'�<��<+�<`8�<���<U�<���<f4�<^]�<m��<���<�=�<=��<:}�<b�<S��<��<���<��<�{�<���<�0�<���<*��<�ݼ<�L�<�͹<T,�<�;�<�<Y�<��<��<��<d��<��<0��<�6�<�ޗ<��<�a�<Z�<ߑ<x��<rp�<q�<��<�ω<26�<�b�<���<x�}<}�x<�t</�o<+l<�-h<kd<s_<DmZ<SU< uO<��I<��D<q*@<�8<<��8<�6< 3<��/<M�+<�&<=!<��<< <�<�;`
�;3��;���;���;p��;*��;y5�;�u�;��;J��;�r�;VЦ;��;WW�;�݄;�Qt;j+a;�IP; *A;73;@�$;�U;��;G��:H��:秦:�&�:��X:	/:��:�v:���9���9���9R4�9�9\�%��S}�����N-���^�wɃ�IJ��ٱ��p���
R��*���\�|�Nd���N���A�S�?�3�K��d��j��@������8d��|k���>ú�Dź-\ƺ�xȺI5ͺlmպẳ���u��-K�"E
�	�.}��E���
�`_
�j���"���լ&��4��*B�+�O�\\���f���m��q�)�q���o�C�k��g�L�b�vT_� m^�'�`��Of�d�n��Zy����bކ��������ꯎ������ؑ�ړ�Ǻ��]���k���q���糧�}���  �  �q=Mr=�u=jh=�8=��=OW=)� =7��<�W�<���<#j�<�'�<d�<c�<#��<���<���<T"�<�o�<w��<P��<��<���<;<�<cU�<�1�<���<���<��<���<q8�<ޣ�<��<O��<�<�}�<���<�f�<~��<t��<��<���<��<@��<���<�k�<~��<+��<�w�<^�<��<�W�<�<?�<^4�<���<q�<�r�<$��<$��<�)�<�c�<!t�<e<�<���<k��<�1�<�{�<	��<���<#��<�<yX�<b��<ѡ�<E��<'�<hH�<�<i��<{��<~��<���<��<c�<��<�޸<=��<�'�<VN�<�;�<J	�<Nͧ<ș�<M�<�<<�<A��<ws�<-��<*�<Ɉ�<�!�<���<9�<�<)w�<�<�{�<�<C�<�bz<?u<�Zp<M�k<��f<�3b<�f]<V�X<٪S<8�N<�,J<��E<R�A<�Y><�0;<�$8<��4<m1<>�,<,}'<�!<��<P<<:�<K�<�<h��;q�;�q�;���;ɪ�;�i�;X��;#�;eF�;f�;ˉ�;ک;3�;�;a��;G!};Dh;OT;��A;�a0;5�;�;���:ȕ�:��:�:O/�:
�n:f�N:�<8:�j(:�:$�
:���9���9��19��gC�,i��!��<�4��pV�9fo� ~��"��s~��s�Ne��U�AyE�`�9��4��l:��JK��)f��ǃ�kS���~����x����ƺ�Pκ��պ�ݺ���$�����j�����k���53��1�����r����Ü����$���/�R�;�lG��DQ���Y��g`�\dd���e�J�e��<d���a�b_�d:]�G\��n]�_Ha�E�g�n�p�|�z��j������JÊ��덻F���6	��lk��ߗ�gc��t�������Zݡ����������  �  ~�=q�=�=9�=WL=�=C==�� =���<K��<�s�<.e�<�q�<��<���<.n�<V�<���<���<v��<���<���<��<���<Gr�<���<j��<���<cn�<-�<���<L��<m��<*�<R�<���<1T�<�<M��<��<���<��<�C�<i�<&c�<h�<o}�<���<��<OR�<y)�<s�<��<1�<�f�<Z��<�5�<9��<���<�d�<4J�<@�< ?�<V8�<�<F��<;��<��<F&�<N�<�H�<�,�<J�< ��<���<co�<�B�<(�<T#�<_1�<XR�<���<���<�;�<J��<q�<�-�<�<*��<l�<�<	�<=+�<�F�<�q�<í�<���<p�<�<GȘ<���<h��<�ݒ<I+�<w��<�
�<�m�<���<8��<��<�r�<휀<Sp{<Ҭu<� p<�qj<�e<w�_<ܽZ<
V<�Q<�M<��I<�F<��B<X�?<%�<<=W9<�5<�\1<�u,<�'<MX!<n�<��<�<5�
<�!<���;"��;�x�;���;��;��;n��;��;!��;�h�;-��;m�;���;9ؗ;iҌ;�[�;r�k;�TU;��?;+;�l;�9;���:���:�M�:a��:�S�:�*y:c4b:`6P:],@:��-:�:@r�9�,�90'9����o9�mr�����>��b*�{K>���L�~U��Y�0�Z��W���Q��I��a@���9�X9�Q�A���T�Iq�T�������]뭺���d�ͺ'�ۺl��	��tN���m��h� �k��ޖ�S� ��?���������������Ԭ�D�|����$���.�˽7��@� �G��cN�v�S�~RX�2s[�T�]���^��}_�gM_�[�^���]��1^�cH`���d���k�;�t�r=��߄��퉻����:�Ӗ��@����8M��+頻}
������������  �  ��=�=��=��=�=a�=�� =�? =�c�<Sv�<p��<+�<�q�<���<�?�<���<_��<�`�<0��<h�<�'�<�<�!�<�.�<s�<t��<G��<���<��<�&�<ʪ�<�9�<���< ��<5��<'1�<���<��<+�<b�<���<�+�<�y�<%��<�a�<��<���<���<���<̱�<��<x�<w�<���<m~�<��<<�<Y��<�`�<���<
M�<���<c��<�x�<�X�<��<��<.��<�C�<�y�<�Z�<@�<���<���<Eo�<%��<���<��<ζ�<��<��<�<ɺ�<<T�<5Ѿ<��<\�<h��<��<S-�<�M�<^��<�ު<�[�<i�<v��<Q*�<ӽ�<�J�<*ԙ<Bb�<��<�Ȓ<F��<��<XU�<5͋<�0�<)Y�<�-�<J��<bӀ<h�{<�Au<X�n<�h<��b<��\<k�W<ZS<�O<�K<cH<�E<v�B<��?<u�<<ch9<�A5<<v0<%+<�%<��<��<j}<��<��<�.<%n<�3�;�r�;Z��;���;��;���;�;e�;T��;�r�;ڟ�;���;�s�;�ٍ;�3�;��k;�S;Ғ:;�	#;;��:*d�:�F�:��:��:.5�:|�u:�hf:L�W:�rF:T�.:{�:KR�9��l9�-p8�;ǸH8h�*R��>�й���S2��$��4#�y1���?���L�W�@�\���\���W�3�O���I��J�
�U�l�HD�����ο���ź<�ںS�LF���9�C���
�Pf	��\�R}��K�����}1��D����:���B��K�]��Oo ��B)�}�0���6���;�I�@�0�D�W�I�qHN��.S�\X�?�\��X`�c�b���c���c�tpc�9�c�pbf�	�k�Kns���}�+����Ɋ�ߐ�7���Λ�I"���R��P@�����㥻/(������䢻�  �  g�=��=��=�1=��=d� =gI =@h�<��<$��<h��<8X�<��<���<�@�<u��<I��<)��<0��<���<�:�<g��<��<��<m6�<�<@��<,��<�T�<X��<�<�D�<���<_:�<)�<���<�Q�<���<5��<ט�<�D�<p��<`:�<{A�<��<��<���<���<��<2��<.�<p��<�{�<ke�<�C�<���<z�<���<��<F��<^��<U(�<C��<�M�<�,�<�<r��<��<���<�/�<��<�z�<���<v��<��<�X�<L��<E��<"�<[��<�{�<I]�< >�<���<��<証<�h�<�ʷ<��<��<�"�<W��<�0�<n�<��<��<��<~��<�=�<U��<]��<2��<�R�<��<��<�1�<Q��<mF�<W��<6��<Na�<G��<��z<�#t<�-m<<Cf<¢_<��Y<n2T<��O<�L<I<�F<@D<�A<�d?<�L<<zy8<��3<:�.<��(<�/#<��<��<�p<�e<(�<C�<�V<^�;�&�;�;�;��;�;&��;e��;ٸ;�D�;�`�;�]�;�q�;��;���;M�;�h;&N;6;3;/N;�f;A�:�1�:C��:E��:jh:Zp:�\f:qY]:��P:��<:+�:9,�9mB�9��86��� �e��i��?��	Ϲ�kչ��ܹ��빜������h0�^�J��Ob�t�k}��|���t�Kj�+�c��f�c�v�?���枺�r����Ѻ���<��+����j�A�L��?K���	���`� �;P��͌��3Q����� �~~)�r�0�E�5���8�\�:�<��!>��A���F���M��OU��5]�j:d���i�a}l�L0m��]l��nk���k�E6o��u����������>I���C��E���R���	�������Ы�����f���`q��n[���  �  �~=�{=�8=j�=<=�K =�2�<��<Qp�<�*�<�1�<�]�<�~�<�f�<���<�<���<��<�$�<?��<-�<"��<���<���<��<�,�<	��<2�<S��<��<�3�<T7�<`W�<~��<��<��< ��<Y�<���<���<��<N�<t��<���<��<��<���<2i�<�=�<�l�<��<I�<�<�<���<ü�<K��<#'�<�?�<�<��<AT�<B1�<�`�<:��<���<&��<���<\7�<�8�<n��<�m�</��<���<֮�<���<���<�A�<1�<|��<�V�<mZ�<�z�<���<l�<��<��<S~�<���<-��<���<�í<�T�<�G�<È�<��<�Z�<���<�n�<��<���<�ӗ<�<W��<��<���<�׊<�e�<��<��<A �<7΂<��<��y<�r<%>k<��c<��\<�]V<�P<_�L<N I<ȋF<�D<t�B<��@<K><P;<��6<��1<�6,<9&<zi <�*<Э<��<�<��<�]	<ʢ<h$<���;ɠ�;2��;U�;Q��;tB�;k��;N��;�]�;��;��;�p�;��;��~;�Nd;��G;b+;P9;���:@��:���:�M�:��k:�4[:�T:Q:�L:?�@:�):�:���9�9����߁�����2�J�p޹1�˹����p�����۹�}��K*���P�x�u�G����������,��2��g�������Ξ�����䕧�I:º'�ߺ������������K�"�wK"�[;���������	�%��$��'��O���X��+�24��>:�� =��=�*�;���9��9��<�u�A�;J���T�Q�_��j���q�I�v�1.x�w��t���s�qCu��z��聻�X�������(��� ���:��ݬ����F����������8���,}�������  �  h6=�+=��=�@=q} =�Z�<���<���<#a�<�]�<ŷ�<;�<m��<��<}a�<�m�<�<wO�<n��<��<U��<�c�<O�<&��<e�<PH�<�&�<�{�<!>�<���< t�<�I�<i:�<�y�<�3�<0��<�t�<z��<v��<f��<���<��<2 �<2��<,A�<�<���<�%�<���<^>�<@�<xO�<���<���<5��<x�<[��<��<G	�<V�<&��<;�<$4�<��<���<
��<���<�\�<p��<��<���<��<���<x��<�i�<{k�<N��<��<�A�<f*�<]�<(��<��<&Ҿ<AI�<�3�<���<|��<Y_�<�B�<�{�<Q.�<]�<W�<���<�k�<��<bܠ<�F�<�,�<н�<�8�<gސ<��<5u�<b��<+�< �<�ǅ<=�<|.�<�<A�x<\Iq<�i<E�a<�NZ<V�S<N!N<9�I<Z�F<�[D<��B<�2A<|?<�=<��9<f5<�0<��)<�#<q�<R�<0�<zO<��<�V<�	<�k<U<:�;�0�;:?�;>G�;�D�;���;��;+��;5��;�;ґ�;���;���;kz;l�_;!-B;��#;�;���:��:� �:cZa:��F:l�;:qf::�}<:��::�/:>:���9�"^9�W�?�o���ҹC[����,�(L��͹Rխ�񀦹�����T����)��B[�eW��K���k����Q��w��Iݛ�A璺����pp���
��B���C�̺��캦��:	�[T"���*��-�m�,�(J'���\�����\	�����
��J��$���)��G5�?>��?C�O*D���A��=�:W9��7�X�8�B�>���H���U��hc��.p��7z��4���8��������}��f{�tz{�t��J-��	���Gɒ�����gW��"���2������q��莶��곻|=���W������  �  	=��= �=�� =� =�|�<X�<9�<ś�<	��<�T�<�<q��<���<g��<���<h�<V�<\'�<5p�<�.�<��<7i�<}��<�C�<ä�<x��<��<	��<��<T��<���<�z�<���<tJ�<f��<���<"�<��<MK�<�q�<$P�<��<O|�<ê�<�\�<���<qC�<��<f�<4S�<K��<Ӑ�<�o�<��<AC�<|��<?��<���<�</%�<k��<�\�<Ͼ�<.��<���<���<��<-�<��<�d�<���<�_�<���<��<��<���<���<U_�<�`�<��<*�<m�<b�<lҼ<���<�<+ϴ< ��<�X�<��<�Z�<���<�s�<ps�<�g�<��<��<�y�<A�</��<�ޓ<RL�<+(�<���<���<WN�<Q8�<��<]��<5��<c9~<��w<�Sp<�Uh<�I`<��X<��Q<EL<��G<��D<��B<}sA<W/@<�><�A<<��8<3E4<�.<*c(<)�!<�<��<�<o<��<�<��	<��<G�<l��;[T�;���;��;���;��;�w�;�z�;�W�;f��;��;Ȣ�;��;\@w;�D\;�3>;��;� ;�T�:�^�:rIs:h�E:#�-:I6&:��(:�.:��-:��!:4�:��99j�����E��<!���'�"3�Gi��ѹ�Ǧ�j���@˲�bS��ޭ+��?d�>���̣��ﱺꤶ�s���E��Ha�������d�����Y��|�Ӻ'���a?��T��V)���1�F/5�1f3�gc-��$�+��a�Ԭ��O�5��L�#��I0�=q<��XE�?�I���I�f{E�-b?�i9�6�5���6�c�<��H�ؚV��Kf��t��!��ۧ���ӄ�p���#��fj����������څ��b��d��������.���d��ȵ��������`⹻�϶�󥲻P��C̪��  �  ��=8�=fw=� =���<o-�<���<���<�S�<���<.�<��<��<H�<B��<B��<�<.�<Y��<3�<A��<e0�<��<�r�<���<�i�<Sn�<8��<���<���<��<.p�<�6�<S�<g��<iF�<C�<���<���<�<EG�<�)�<v��<�N�<ht�<�<V��<u��<��<��<`�<Ԓ�<�q�<=f�<��<�S�<]��<���<-��<E��<���<�B�<��<�k�<K�<�y�<��<Ն�<u��<|f�<�<�<n�<�,�<x��<�P�<�3�<���<���<��<��<(v�<��<fB�<�9�<M��<�w�<b��<9��<{4�<.�<�@�<��<�n�<�E�<[�<�c�<��<]'�<)��<�E�<���<g��<��<t�<�L�<_�<\��<���<_߄<�{�<��<��}<�vw<��o<��g<��_<�X<>Q<d�K<�UG<�VD<�]B<�A<��?<�H><��;<-�8<��3<N-.<]�'< Y!<{\<BS<r<�<ƣ<Q�<m�	<��<İ<+�;wV�;:�;���;�ۿ;pĳ;f:�;A9�;0(�;��;L4�;2�;�B�;6v;}[;�<;�C;�.�:���:QT�:i:��;:��$:G�:v�":��(:E):�:ko :?��9�T�8";��Ĺ�T�-�*��;0�k�"��D��<Թ[ �������)#�W�,���g�Ø��狀Nȶ��̻��������O~��$���J���n��Z����ֺ����"�܌�C�+�ts4�7�7�C�5���/�}x&��|�V��~��٘��u�m��7%���2��?���G�L��wK�e�F��@���9���5�,<6�;}<�,�G��
W�ng���v��<��o焻����E��	F��-d���΀�X^���v������f��"͞��0���������
���Q��h���շ��|������i���  �  	=��= �=�� =� =�|�<X�<9�<ś�<	��<�T�<�<q��<���<g��<���<h�<V�<\'�<5p�<�.�<��<7i�<}��<�C�<ä�<x��<��<	��<��<T��<���<�z�<���<tJ�<f��<���<"�<��<MK�<�q�<$P�<��<O|�<ê�<�\�<���<qC�<��<f�<4S�<K��<Ӑ�<�o�<��<AC�<|��<?��<���<�</%�<k��<�\�<Ͼ�<.��<���<���<��<-�<��<�d�<���<�_�<���<��<��<���<���<W_�<�`�<��<.�<m�<b�<pҼ<���<�<0ϴ<%��<�X�<��<�Z�<���<�s�<rs�<�g�<��<��<�y�<A�<-��<�ޓ<OL�<'(�<���<���<RN�<L8�<��<X��<0��<Z9~<��w<�Sp<�Uh<�I`<��X<��Q<EL<��G<��D<��B<�sA<]/@<�><�A<<��8<<E4<��.<3c(<2�!<<�<�<v<��<�<��	<��<G�<i��;UT�;}��;���;~��;��;�w�;|z�;�W�;S��;��;���;��;8@w;yD\;�3>;��;�� ;�T�:�^�:7Is:9�E:��-:,6&:x�(:�.:��-:��!:.�:��9�9v�����E��<!���'�!3�Gi��ѹ�Ǧ�j���@˲�bS��ޭ+��?d�>���̣��ﱺꤶ�s���E��Ha�������d�����Y��|�Ӻ'���a?��T��V)���1�F/5�1f3�gc-��$�+��a�Ԭ��O�5��L�#��I0�=q<��XE�?�I���I�f{E�-b?�i9�6�5���6�c�<��H�ؚV��Kf��t��!��ۧ���ӄ�p���#��fj����������څ��b��d��������.���d��ȵ��������`⹻�϶�󥲻P��C̪��  �  h6=�+=��=�@=q} =�Z�<���<���<#a�<�]�<ŷ�<;�<m��<��<}a�<�m�<�<wO�<n��<��<U��<�c�<O�<&��<e�<PH�<�&�<�{�<!>�<���< t�<�I�<i:�<�y�<�3�<0��<�t�<z��<v��<f��<���<��<2 �<2��<,A�<�<���<�%�<���<^>�<@�<xO�<���<���<5��<x�<[��<��<G	�<V�<&��<;�<$4�<��<���<
��<���<�\�<p��<��<���<��<���<z��<�i�<~k�<R��<��<�A�<l*�<]�<0��<��</Ҿ<II�<�3�<���<���<b_�<�B�<�{�<X.�<
]�<\�<���<�k�<��<cܠ<�F�<�,�<̽�<�8�<aސ<��<-u�<Z��<�*�< �<�ǅ<=�<t.�<�<2�x<OIq<�i<=�a<�NZ<R�S<M!N<<�I<_�F<�[D<��B<�2A<+|?<�=<��9<f5<�0<��)<.�#<��<b�<?�<�O<�<�V<	�	<�k<U<4�;�0�;*?�;)G�;�D�;���;��;��;��;��;���;���;���;�jz;*�_;�,B;��#;�;O��:ڮ�:� �:Za:c�F:4�;:Hf::�}<:��::�/:
>:���9�"^9UW�F�o���ҹD[����,�(L��͹Qխ�񀦹�����T����)��B[�eW��K���k����Q��w��Iݛ�A璺����pp���
��B���C�̺��캦��:	�[T"���*��-�m�,�(J'���\�����\	�����
��J��$���)��G5�?>��?C�O*D���A��=�:W9��7�X�8�B�>���H���U��hc��.p��7z��4���8��������}��f{�tz{�t��J-��	���Gɒ�����gW��"���2������q��莶��곻|=���W������  �  �~=�{=�8=j�=<=�K =�2�<��<Qp�<�*�<�1�<�]�<�~�<�f�<���<�<���<��<�$�<?��<-�<"��<���<���<��<�,�<	��<2�<S��<��<�3�<T7�<`W�<~��<��<��< ��<Y�<���<���<��<N�<t��<���<��<��<���<2i�<�=�<�l�<��<I�<�<�<���<ü�<K��<#'�<�?�<�<��<AT�<B1�<�`�<:��<���<'��<���<]7�<�8�<o��<�m�<0��<���<خ�<���<���<�A�<1�<���<�V�<vZ�<�z�<���<l�<��<��<`~�<���<:��<Ð�<�í<�T�<�G�<ˈ�<��<�Z�<���<�n�<��<���<�ӗ<ꤔ<O��<��<���<�׊<�e�<��<���<4 �<+΂<��<��y<�r<>k<��c<��\<�]V<�P<b�L<U I<ӋF<�D<��B<Ϸ@<%K><g;<��6<��1<�6,</9&<�i <�*<�<��<�<��<�]	<΢<h$<���;���;��;�T�;.��;KB�;>��;��;�]�;��;��;�p�;n�;&�~;@Nd;|�G;+;9;5��:���:1��:�M�:D�k:74[:nT:�Q:ӍL:)�@:�):�:{��9�9����߁�����2�I�p޹0�˹����o�����۹�}��K*���P�x�u�G����������,��2��g�������Ξ�����䕧�I:º'�ߺ������������K�"�wK"�[;���������	�%��$��'��O���X��+�24��>:�� =��=�*�;���9��9��<�u�A�;J���T�Q�_��j���q�I�v�1.x�w��t���s�qCu��z��聻�X�������(��� ���:��ݬ����F����������8���,}�������  �  g�=��=��=�1=��=d� =gI =@h�<��<$��<h��<8X�<��<���<�@�<u��<I��<)��<0��<���<�:�<g��<��<��<m6�<�<@��<,��<�T�<X��<�<�D�<���<_:�<)�<���<�Q�<���<5��<ט�<�D�<p��<`:�<{A�<��<��<���<���<��<2��<.�<p��<�{�<ke�<�C�<���<z�<���<��<F��<^��<V(�<C��<�M�<�,�<�<r��<��<���<�/�<��<�z�<���<y��<��<�X�<R��<L��<#"�<e��<�{�<U]�<>�<���<��<���<�h�<�ʷ<��<*��<�"�<d��<�0�<x�<��<��<��<��<�=�<Q��<W��<)��<�R�<��<��<�1�<A��<]F�<G��<&��<?a�<8��<��z<#t<�-m<.Cf<��_<��Y<m2T<��O<�L<&I<��F<@D<'�A<�d?<�L<<�y8<��3<Z�.<
�(<0#<�<��<�p<�e<5�<L�<�V<^�;�&�;q;�;��;��;���;2��;�ظ;oD�;|`�;~]�;Yq�;G�;���;�L�;��h;�%N;�:3;�M;Ff;��:�1�:�:��:	h:�Yp:�\f:JY]:��P:o�<:�:(,�9cB�9��8D����e��i��?��	Ϲ�kչ��ܹ��빜������h0�^�J��Ob�t�k}��|���t�Kj�+�c��f�c�v�?���枺�r����Ѻ���<��+����j�A�L��?K���	���`� �;P��͌��3Q����� �~~)�r�0�E�5���8�\�:�<��!>��A���F���M��OU��5]�j:d���i�a}l�L0m��]l��nk���k�E6o��u����������>I���C��E���R���	�������Ы�����f���`q��n[���  �  ��=�=��=��=�=a�=�� =�? =�c�<Sv�<p��<+�<�q�<���<�?�<���<_��<�`�<0��<h�<�'�<�<�!�<�.�<s�<t��<G��<���<��<�&�<ʪ�<�9�<���< ��<5��<'1�<���<��<+�<b�<���<�+�<�y�<%��<�a�<��<���<���<���<̱�<��<x�<w�<���<m~�<��<<�<Y��<�`�<���<
M�<���<c��<�x�<�X�<��<��</��<�C�<�y�<�Z�<A�<���<���<Jo�<*��<���<��<ض�<��<��<�<غ�<MT�<FѾ<��<o�<z��<��<d-�<N�<m��<�ު<�[�<r�<|��<T*�<ӽ�<�J�<%ԙ<;b�<��<�Ȓ<9��<��<HU�<$͋<�0�<Y�<�-�<9��<RӀ<L�{<�Au<C�n<�h<��b<��\<i�W<^S<�O<�K<cH<�E<��B<��?<��<<�h9<B5<`v0<A%+<	�%<��<ܗ<�}<�<�<�.<*n<�3�;�r�;E��;���;ݧ�;}��;G�;&�;��;hr�;���;M��;�s�;Tٍ;m3�;v�k;2S;j�:;_	#;�;���:�c�:0F�:��:٤�:5�:?�u:ahf:-�W:�rF:F�.:q�:?R�9��l9�-p8�;ǸI8h�*R��=�й���R2��$��4#�y1���?���L�W�?�\���\���W�3�O���I��J�
�U�l�HD�����ο���ź<�ںS�LF���9�C���
�Pf	��\�R}��K�����}1��D����:���B��K�]��Oo ��B)�}�0���6���;�I�@�0�D�W�I�qHN��.S�\X�?�\��X`�c�b���c���c�tpc�9�c�pbf�	�k�Kns���}�+����Ɋ�ߐ�7���Λ�I"���R��P@�����㥻/(������䢻�  �  ~�=q�=�=9�=WL=�=C==�� =���<K��<�s�<.e�<�q�<��<���<.n�<V�<���<���<v��<���<���<��<���<Gr�<���<j��<���<cn�<-�<���<L��<m��<*�<R�<���<1T�<�<M��<��<���<��<�C�<i�<&c�<h�<o}�<���<��<OR�<y)�<s�<��<1�<�f�<Z��<�5�<9��<���<�d�<4J�<@�< ?�<V8�<�<F��<;��<��<F&�<N�<�H�<�,�<L�<$��<���<ho�<�B�<(�<^#�<k1�<eR�<Ȉ�<���<�;�<\��<��<�-�<'�<<��<}�</�<�<J+�<�F�<�q�<ʭ�<���<p�<�<CȘ<���<_��<�ݒ<;+�<h��<�
�<�m�<睊<&��<��<�r�<ݜ�<5p{<��u<� p<�qj<�e<p�_<۽Z<
V<�Q<+�M<ШI<�F<��B<w�?<G�<<`W9<�5<�\1<v,<�'<lX!<��<��<�<E�
<�!<	��;"��;�x�;޷�;��;���;<��;���;᱿;�h�;㠲;"�;���;�ח; Ҍ;�[�;��k;]TU;P�?;�+;zl;_9;<��:$��:�M�:)��:�S�:�*y:54b:?6P:G,@:��-:�:3r�9�,�9('9���o9�mr�����=��b*�zK>���L�~U��Y�0�Z��W���Q��I��a@���9�X9�Q�A���T�Iq�T�������]뭺���d�ͺ'�ۺl��	��tN���m��h� �k��ޖ�S� ��?���������������Ԭ�D�|����$���.�˽7��@� �G��cN�v�S�~RX�2s[�T�]���^��}_�gM_�[�^���]��1^�cH`���d���k�;�t�r=��߄��퉻����:�Ӗ��@����8M��+頻}
������������  �  �q=Mr=�u=jh=�8=��=OW=)� =7��<�W�<���<#j�<�'�<d�<c�<#��<���<���<T"�<�o�<w��<P��<��<���<;<�<cU�<�1�<���<���<��<���<q8�<ޣ�<��<O��<�<�}�<���<�f�<~��<t��<��<���<��<@��<���<�k�<~��<+��<�w�<^�<��<�W�<�<?�<^4�<���<q�<�r�<$��<$��<�)�<�c�<!t�<e<�<���<k��<�1�<�{�<
��<���<%��<�<}X�<g��<ס�<L��</�<rH�<�<v��<���<���<ħ�<��<c�<-��<�޸<O��<�'�<fN�<�;�<W	�<Xͧ<Й�<S�<Ő�<=�<?��<ss�<&��< �<���<�!�<|��<9�<�~�<w�<m�<�{�<Ⲃ<$�<ebz<�>u<�Zp<=�k<��f<�3b<�f]<Z�X<�S<F�N<�,J<�E<m�A<�Y><�0;<�$8<��4<�1<`�,<M}'<��!<��<h<<N�<[�<��<s��;q�;�q�;���;���;�i�;(��;��;'F�;#�;���;�٩;��;� �;��;� };�h;�NT;��A;pa0;�;�;���:n��:���:��:&/�:��n:9�N:�<8:�j(:�:�
:y��9���9��19���gC�,i�� ��;�4��pV�9fo� ~��"��r~��s�Ne��U�AyE�`�9��4��l:��JK��)f��ǃ�kS���~����x����ƺ�Pκ��պ�ݺ���$�����j�����k���53��1�����r����Ü����$���/�R�;�lG��DQ���Y��g`�\dd���e�J�e��<d���a�b_�d:]�G\��n]�_Ha�E�g�n�p�|�z��j������JÊ��덻F���6	��lk��ߗ�gc��t�������Zݡ����������  �  !�=��=��=��=��=�=�3=l� =���<���<��<�4�<#��<~~�<���<�]�<l�<��<&L�<5��<�i�<���<���<�V�<��<�a�<)�<���< ��<���<<q�<�+�<'�<A��<̈�<8
�<	V�<�x�<���<˪�<���<-��<Sh�<ވ�<���< ��<���<"]�<!v�<�/�<"��<T��<)V�<���<��<���<S�<,��<��<2��<*'�<��<+�<`8�<���<U�<���<g4�<_]�<n��<���<�=�<?��<=}�<f�<W��<!��<���<��<|�< ��<�0�<���<8��<�ݼ<M�<ι<e,�<�;�<#�<h�<��< ��<��<k��<��<3��<�6�<�ޗ<��<�a�<R�<�ޑ<l��<dp�<c�<��<�ω<"6�<�b�<q��<\�}<d�x<�t<�o<l<�-h<fd<s_<HmZ<[U<,uO<��I<��D<�*@<9<<��8<�6<< 3<�/<l�+<$�&<=!<��<1<<�</�;j
�;3��;���;���;T��;��;M5�;zu�;��;��;�r�;Ц;j�;W�;I݄;7Qt;�*a;GIP;�)A;�3;��$;�U;f�;���:	��:���:z&�:W�X:�/:��:�v:���9���9���9L4�9�9j�%��S}�����N-���^�wɃ�HJ��ٱ��p���
R��*���\�|�Nd���N���A�S�?�3�K��d��j��@������8d��|k���>ú�Dź-\ƺ�xȺI5ͺlmպẳ���u��-K�"E
�	�.}��E���
�`_
�j���"���լ&��4��*B�+�O�\\���f���m��q�)�q���o�C�k��g�L�b�vT_� m^�'�`��Of�d�n��Zy����bކ��������ꯎ������ؑ�ړ�Ǻ��]���k���q���糧�}���  �  F>=�,= A=�`=�l=~J=�� =�J =N��<���<���<���<m;�<���<J�<���<� �<9��<�W�<)�<4��<:8�<�%�<,��<��<h.�</��<Fk�<Br�<��<U��<0��<�<�B�<�.�<��<���<M��<`h�<q!�<"�<�Z�<r�<�)�<ȁ�<D��<��<y��<���<���<8�<q%�<�>�<ny�<��<���<f�<_�<���<�w�<nI�<��<]��<B��<�G�<K�<
��<w��<�<�1�<n��<�W�<XL�<�Z�<�V�<>�<�e�<6<�<���<���<Y��<���<�ӿ<>w�< ��<8��<៸<�2�<dz�<M�<<j�<�ܩ<��<�Y�<���<�o�<���<�D�<�v�<	�<% �<�</�<W�<X�<�V�<���<�<A�<R�<�z<Dv<�cr<�o<�l<��h<K9e<��`<ɱ[<��U< �O<f4I<-EC<�><��9<;86<�m3<w�0<� .<�k*<^�%<"6 <��<
v<�
<�<S%�;���;���;Nt�;���;���;#��;��;k��;�̼;��;�4�;4��;���;ъ;�v~; �i;a�X;]J;eb>;r3;%+(;�E;O�;G��:�]�:#�:�Q|: �::��:/}�9�Ы9�7�9s'�9��9��I9
��8�ݸ�r��<P��vP�������#��z����z��B���{��t��vay��&`�Y�R���T��f�^��V����!��CX����Ⱥ kͺA�̺�Ⱥ�úG,��Bºa�ʺ��ٺ���x� �[�
�1Q����n�T��v��x����N�9��"+���9���I��PY�l�g�Ms�c�z��K~���}�,�y�Qt��om�psg��c�3�b��Jf���m���w��偻����i$������m��H{���ُ��E��:{������G��옻�l��L�����㬻�  �  �� =Q� =w� =\� =�� =�� =l� =| =0O�<�<�<��<=��<'��<-��<Ĵ�<�x�<]��<!��<�|�<�x�<C�<���<��<���<K��<(�<�y�<#�<�=�<���<X��<�o�<��<�x�<7��<g(�<u0�<{��<I$�<���<(�<8�<���<G��<FP�<���<E�<� �<mT�<�<�`�<�^�<I�<�U�<���<���<�<��<���<~�<Q�<�j�<Y�<� �<E��<;w�<���<���<���<��<�}�<�n�<}��<3�<f�<�d�<d��<���<���<	��<>�<`��<T޾<�O�<jL�<�¸<���<�>�<���<���<��<ܬ<^5�<�K�<�V�<���<�<�6�<&�<�2�<���<��< L�< s�<sO�<h��<���<��<d��<Pԁ<�}<ax<Pt<ˮp<��m<�k<&i<=�e<�a<�t\<&V<�?O<�BH<8�A<��;<�A7<@�3<d1<R�.<'0,<��(<��$<�<9v<�<�-	<c<�;H�;�Z�;T�;K��;���;K�;�7�;��;`b�;�>�;�;���;M�;��;_�s;w`;�3P;
(D;��:;F�2;˦);:;�;rm�:{��:
��:uHh:(8:�6�9,my9�G29��#9�@+9�#9�?�8�Vq�� 8�%<ѹLQ+�kSo���a���_º�ɺ�?Ǻ����2���2������Vr�]e���j��›.����f��y���ѺR(ۺXsܺ��ֺ��̺��ºr���L����\ĺg�պ����\V��G��� ���"�b/!�V���W��]��F��#�ȿ/��?�&FP��a��q�Ϝ}��炻�����䃻�_���f{��Ys��Pl�#h���g��%l���t��L���Ɔ�U������0z��Yӓ�����꜐�7Ȏ�����T��_Ғ��O��v	��b
���Z���,���  �  �0 = =5 =Gq =E� =�� =�` =x��<=��<|��<�h�<]#�<�&�<Χ�<���<��<���<���<���<_��<��<�:�<��<=7�<���<&@�<��<o<�<b�<# �<Zj�<��<&��<̍�<���<�a�<�U�<l��<6��<c�<�z�<�f�<���<���<z�<��<̀�<u}�<D��<'��<���<���<��<���<���<���<o�<45�<v��<$��<��<���<���<���<��<��<]�<g �<o��<��<��<?��<�4�<���<�`�<6��<��<0��<��<r��<M��<�`�<E)�<O|�<�k�<��<���<ǐ�<O#�<�4�<椯<^t�<d��<���<$��</��<�<�<�J�<���<�X�<�8�<�o�<EǏ<� �<5�<�@�<�
�<�L�<�0�<-��<��{<f�v<6xr<Fgo<�%m<�?k<&'i<�Jf<b=b<��\<PCV<��N<�}G<|@<�g:<M�5<V�1<IN/<--<0�*<��'<f�#<SF<i�<�<L�<(��;̺�;\u�;&��;Dc�;���;ߴ�;e��;L7�;���;x��;�B�;���;D�;F	�;C�;�l;�Y;|J;xv?;�7;i�1;1*;Ͷ;��;���:Hy�:�v�:��X:D3:�,�9�+9�nz8,^8Vٗ8WԦ8��28>9r��m��n<�?���V��s����кhFغ�7պ]ɺѶ�l衺�E����I9s��z�ʖ��qQ�������κ��ߺyl�@���޺jHѺDEú~}�����q��GGԺ�ﺕ~�۶��  �qW'���)��<(�9$�8��+�G$ ��2'��3���B�I�T�og��w�nZ��o����1���G���X���0���kw���o��Wk��ak��kp���y��X���1���L��L�������@_��NP��2`�������g���l�����!�����������Ю��I���  �  (w=�G=�9=�4=�=*�=�p=�� =y��<#��<��<���<s�<��<���<|��<&��<�f�<_4�<�
�<���<�#�<W$�<��<���<���<a��<��<~��<�l�<o�<B��<��<P:�<$&�<b��<���<���<�3�<��<Z��<͛�<��<���<���<M�<���<�`�<Au�<��<Ah�<}�<ф�<���<� �<��<�l�<�\�<���<rh�<�3�<���<�l�<~��<W)�<#K�<W��<Yf�<[��<��<���<қ�<;��<*��<��<���<�M�<�7�<ɪ�<���<��<���<ؽ�<�?�<�'�<�b�<qù<��<c%�<ҳ<�
�</ԭ<SG�<��<�Ţ<D,�<K�<�<�ז<��<9Г<!Β<��<c��<׏<�[�<�x�<1�<雇<�<;1�<!v<={<ܾw<��t< r<�o<e�k<HUg<�?b<	l\<�V<ѤO<�tI<��C<�'?<�=;<��7<*�4<pO1<_H-<Ci(<��"<�<�<O<��<���;km�;��;d��;Y��;8��;^)�;��;���;R��;c�;<M�;���;�"�;9�;�ɋ;Ǌ�;��u;�ii;8)_;�U;�\K;+?;Z0;��;yL;���:c%�:���:忆:le:�UK:�;:�-:�}:P�:0)�9z.9��v��	�� ��e�L�?�}�s���d���Ǘ� ���VT����d�,�E��;-��N�O����,�d�E��	f�h���_?������X���ZD�������ˋ�����㊺_���8ꢺ#����ͺ���m��ZZ����5U���@K�H��?�?��z?"��1�� A�,)Q���_��ek�	Es���v��v��r��l�68e��_�[���Y��X\��b�Qwj�It��C}�SI��lt�����wy���`��ˊ��h���8A���}��9������������O���  �  ��=�c=�U=�N=6=��=Z�=4� =%��<�
�<Y��<C�<�J�<;��<�#�<���<-�<��<)a�<�1�<���<�F�<�I�<��<m�<���<)��<���<���<��<��<��<���<�(�<��<ו�<ͻ�<��<�4�<1��<��<���<�K�<�%�</�<�6�<a�<6��</��<?�<��<&��<y��<���<u_�<�F�<��<��<6��<���<*^�<��<%��<ë�<�O�<Jv�<,/�<���<D��<	H�<���<���<���<I��<|�<���<�2�<<�<���<׸�<��<��<���<5n�<�\�<G��<���<�C�<�N�<���<�,�<-��<dm�<~��<s��<*f�<�'�<�]�<��<�Z�<��<���<;�<"�<��<耎<���<�_�<�χ<��<Pi�<D�<�{<��w<L�t<��q<b�n<|ek<� g<6b<4K\<`V<��O<��I<t3D<��?<�;<�R8<| 5<�1<�-<��(<��"<�J<�<(�<�Q<���;Ty�;�;���;���;���;L��;+S�;U]�;�e�;��;��;	�;���;'�;E��;(T�;��v;u*j;�n_;�sU;H�J;q>;)�/;~8;��
;c��:F3�:��:
��:��k:�eR:��A:��3:�":*�:�=�9
a@9�+�pv����
�*�E�ev��狺�-��;Г�o"��v~�!�_��)A���(����o ��'���?�oA_�	��N荺̪���{���'���֑��x��)x���;��;������fOͺ�P⺺�����������g\�V��bF������� !���/���?���O���]�!`i�('q���t�[.t�mp��j���c���]���Y���X��[��`�/�h��Rr��{��z���Ƀ�2����F���i���Ă����D����ڇ�|w���
���ꗻ=W��P����  �  !�=3�=d�=��=�u=�.=��=�	=j2 =g|�<<��<G��<���<���<N��<ϑ�<��</�<���<w��<�D�<{��<��<KR�<ԓ�<���<�l�<aY�<��<M��<%��<���<���<���<���<�G�<z�<gh�<\2�<� �<`��<�@�<��<��<0��<���<��<
��<��<ڠ�<���<o�<�?�<Ʉ�<r�<^�<8m�<dO�<��<&�<���<�}�<1��<��<���<b��<T��<9-�<�<
��<DW�<��<2��<���<R��<܌�<���<���<W�<�<��<���<o=�<��<��<�-�<q��<ĸ<��<�[�<���<�W�<"ت<�/�<���<��<ޜ<��<[֗<'
�<���<y��<Ŋ�<֊�<�^�<|�<��<�ފ<+^�<y��<��<�{�<�v|<��x<� u<��q<�n<��j<~�f<G}a<�[<��U<x�O<v/J<$E<�@<��<<}9<�76<�2<$v.<�y)<��#<t<:<�<��<]� <�l�;��;���;�2�;d�;5��;��;���;��;���;rط;e��;�M�;��;&�;cq�;<z;},l;E`;~�T;�0I;#5<;,<-;�?;�	;��:���:�n�:<�:f�}:Y�e:��T:=?E:�1:59:3B�9x�q9J�!7��n�)��E�1�j�_����WQ�����
���Z�l�`P�j�3��|�x��(����`�.�Z�L��l�9Մ�%������A��N�������l捺�L����������X����̺��޺7��8���p}������@���`O��ן�������I�&g,���;�uK�A�X�0�c�!5k�)�n���n���k�*^f�HS`�'�Z�@�V�ƦU���W���\��yd���m���v�n�~���o��{ȃ�v���K~�����ⅻN���;>��:I��I����<��S����  �  �1==�=��=;�=�z=��=�L=�y =� �<D�<ҁ�<���<b��<���<5��<ǰ�<E�<?��<?�<f��<.�<�<�<���<F�<�U�<L=�<}$�<N1�<�}�<�<x��<���<���<�A�<���<o�<��<��<�.�<h�<���<f��<8��<��<{�<�*�<��<ǂ�<(�<X��<��<��<�s�<��<s�<��<�[�<��<���<|��<M�<gw�<���<!F�<���<�i�<���<K�<���<���<"~�<\)�<h��<>��<��<�R�<�A�<*��<�U�<��<��<���<y��<J��<I��<�F�<�r�<dY�<��<��<�ݮ<vp�<��<�_�<��<��<,8�<5�<�<؍�<�N�<5�<��<)�<-s�<嫍<ь�<
!�<Z��<{Ӄ<|9�<�}<&Py<'`u<ʥq<��m<F�i<ke<�{`<�$[<|�U<^P<�J<� F<� B<!g><�;<ϴ7<��3<e�/<ψ*<�$<$2<�J<�=<%T	<��<9��;`��;�!�;[=�;k��; ��;��;I�;�.�;2��;Td�;(z�;�|�;��;xO�;/M�;��~;��n;�`;jQS;o/F;J8;�$);`�;��;��:��:�t�:Jw�:PZ�:��:�n:\]:��F:z�':�`�9�9E0�8�t�<#������H>���\��(m��oo�9�e�2�R�06:��� �	u��w��z���ɩ���rj3��R��q�ު��t���됺Ej������������Q0��sP��m���%g̺ՎںZ��M�캌��I��!���� S���*������?�'��6��5D���P�'[��Rb��f�0�f��Od�)`��[��;V�>�R��dQ���R� qW�uz^�n)g��Rp���x��[������I�����؄�������%m����咻���Oٚ�y����  �  e�=y~=�q=�W=)!=��=<=&�=x� =e��<-#�<���<�.�<�<�U�<n��<?��<&�<Aq�<P��<�^�<c��<
��<���<���<B�<��<<��<g��<|��<5G�<���<�T�<���<��<=��<X�<]��<���<	F�<���<�}�<�a�<�a�<^�<y5�<>��<��<��<J��<�'�<K��</��<���<=Z�<�p�<&��<���<���<5��<K�<��<���<��<���<I'�<�<˺�<��<mV�<���<���<�@�<I��<�<:b�<Ņ�<�w�<�<�<(��<���<�B�<�"�<�4�<ar�<�ý<��<��<��<�c�<���<zd�<	�<��<�Z�<5*�<N5�<���<�@�<�J�<��<6�<��<鸒<Cp�<���<@�<�7�<p�<]V�<=��<E��<��~<��y<�lu<�q<��l<�oh<��c<k_<��Y<�T<��O<$_K<�*G<�hC<�?<��<<=09<�E5<r�0<g�+<��%<X<k�<��<s<}A<!&�;��;f�;@�;3��;�p�;j��;��;�W�;.�;��;�X�;���;�Q�;⢕;-�;LZ�;��p;�`;�P;E�A;ۋ2;�/#;k~;6�;F��:U��:;з:Α�:�:���:]m�:u�t:K[:ȇ9:��:[)�9*#$9�0X�@6��)��S��:2��|B�!G�p�A��4�f!�V��w���6۹�ӹV�߹ � �'��l8��$X�P
u��;���펺$B���\��臟�X饺�/��kE��Uú�-κ��׺E޺h��D*��W���交�躖�����i�	��R��L"� �/��F<���G�X�P��W��[�\�\�~�[�TY��VU��Q��N��RM��qN�09R�{}X��`�V�i�h�r�G�z������1��H1�����%ۈ�����΍��搻���)��ʳ�������  �  ��=��=u�=2�=k\=*�=he=�=v� =�9 =���<u��<�o�<�x�<���<�K�<w�<��<�:�<�}�<��<@�<�<��<<r�<L��<��<��<Vh�<!M�<�Q�<z�<���<�<��<���<o�<q��<H��<y-�<���<���<H��<�<���<��<�9�<�j�<�U�<|�<j��<\=�<���<˯�<��<���<�D�<��<���<��<���<�2�<[�<�]�<��<���<��<0Q�<g��<���< �<�<�'�<iC�<�^�< s�<jy�<�n�<mW�<e>�<c0�<�9�<fb�<P��<&�<`�<��<���<dI�<L��<PԲ<=ů<���<�o�<iT�<�Y�<N��<���<���<���<���<��<���<�3�<
ϑ<Q�<���<.��<�v�<��<�P�<��<K�<>z<�u<6 p<�Jk<��f<��a<d]<�cX<�S<�O<�K<�G<NyD<;A<��=<�G:<*6< v1<n*,<s^&<M; <a�<|�<�<��<�b<���;p��;��;�	�;��;���;�y�;���;}��;���;lp�;�2�;:	�;K�;�d�;"��;/<q;�'^;�/L;�*;;��*;1S;�j;���:���:���:�k�:��:�ơ:�@�:c��:t'�:�?i:�E:<4:�Q�96�d9ճ8����z����ع�#��<����E��<��Ό
�������ܹ��ƹ@����Ĺ��߹wB��#���D�g.f�偂��珺0M��i���˭���������ź�ͺ�ӺEb׺��ٺ��ٺ ,ٺ"�غ�ۺ���V^�A�������@���z)��\4��>��F�oBL��lP��R�.S�% R�v3P�D�M���K�`�J�H�K�ΜN�hT���[���d�f;n�c�w�����ۃ���*���ڟ���&��ܡ��<���,������E������  �  *�=/�=S�=��=sm=��=g=!�=�=�o =��<���<D��<���<<!�<���<S6�<S��<���<5��<"��<��<��<���<M��<���<y
�<���<���<�Z�<��<k��<V��<�<�W�<_��<�O�<N�<s��<���<��<��<�G�<_�<�H�<���<lS�<|q�<�Z�<�%�<J��<ɾ�<ɫ�<���<T��<@2�<���<�.�<���<H��<���<{�<u�<
`�<I!�<C��<<��<B��<��<J1�<�&�<���<��<��<]o�<hL�<�5�<�.�<L:�<�\�<���<:��<m]�<���<�P�<_��<GҼ<m��<�R�<*��<ֲ<��<|�<�<�-�<�r�<�ա<�X�<���<�ǚ<���<�і<��<�r�<\�<.Z�<ܰ�<^Ԍ<���</P�<ë�<�؂<��<}z<�Ft<�n<LUi<C2d<+O_<ůZ<[ZV<SR<��N<�/K<'H<��D<��A<N�><%�:<"e6<ׅ1<�+,<~{&<� <Q�<�<��<�1
<�<�> <�S�;��;���;�l�;M��;nO�;�.�;���;���;%9�;c�;���;�;!~�;��;�o;�SZ;kF;�3;�!;��; �;��:l��: �:Y�:�:G��:{�:���:���:c�l:,UF:3:cK�9��9�M�8C|3�6B*�1_���F���ӹ5鹋[���P������I8չG�Ĺ�������'iӹ�	�����n�:��)`��􂺉ה�:���U��w���oɺ�AѺ�ֺmhں��ۺEۺ30ٺ�Rֺ��ӺY�Ӻ�ֺ#3޺ ?�sX��W��9��L��$��r-��'5���;�6JA���E�(I�<@K��gL���L�"L�+K���J��=K���M�N<R�`Y���a���k���v�����+~���򉻙ߍ�a>������N��% ���"�����Gܙ�ߠ���  �  ��=�=�=ܬ=LN=��=�;=y�==`� =B =9S�<T��<���<�Z�<2��<�+�<���<?�<��<r��<��<7��<���<�a�<��<s�<���<���<�<,��<~<�<p��<���<���<�b�<��<���<��<qA�<���<|��<K?�<[�<q5�<;��<�<C�<��<;��<���<� �<�:�<��<���<Vf�<Q��<�E�<��<�:�<&��<|�<W?�<_�< ��<YQ�<���<�w�<���<�!�<J��<���<Y6�<ɾ�<Q�<���<���<���<'��<MK�<���<e�<}�<���<dA�<s��<}��<pw�<���<\M�<��<���<���<�Y�<�ҧ<�^�<���<���<�.�<(қ<���<XT�<3H�<g�<+��<
�<Db�<`��<���<�E�<���<5ς<��<�By<��r<��l<�g<p�a<��\<� X<��S<5gP<Z7M<�PJ<f�G<��D<��A<�[><�e:<��5<��0<�y+<��%</t <X!<?<�<�?<g~<<�<��;���;k��;5+�;&:�;���;�5�;/��;��;��;V�;���;�֙;O�;~G�;�Zl;"�T;�S>;�);�;=;OI�:1��:=��:Pǿ:1�:�D�:�Ӧ:��:[ʒ:B+�:�d:^�;:�7:��9�Ń9ݲ9l��7��t�=��a�K��C���֢�n&��3ҹv�߹S�����,ٹ$Oѹ+Eѹ�L߹�l���Y��;��d��ׇ�}���Z1���xĺz�ӺJߺZ��E�꺌������%�ySݺ��׺=ԺԺ\jغ����o����	�	0�����!��*(��-��2�w�7�,7<�]�@��D��uH��K���L�(M�%PM�6�M�F�O��pS��Y���a�^l�Rx����u�������r���{��B����������F᜻1j���~��g���  �  B�=�= �=�p=1=�}=��=,Z=� =�x =C+ =���<�i�<M��<&^�<r��<��<?�<e�<H��<�g�<2�<Z�<��<���<�d�<���<��<�6�<��<���<U\�<���<���<X��<���<#��<1��<��<g��<��<���<���<f�<J��<D�<ds�<�t�<�h�<{o�<���<��<΍�<�/�<���<d�<���<C&�<M`�<*��<R��<-:�<���<@k�<A�<Ȱ�<��<��<�<��<���<��<{r�<o��<n�<+��<eV�<U�<6��<� �<���<~��<��<�N�<;�<�5�<�4�<��<�T�<$��<��<�?�<Ĭ<�q�<�<�<:�<\ߣ< ��<s)�<7��<��<p��<�=�<��<*�<�l�<w<`�<	�<}�<|[�<E|�<��~<x<qeq<��j<?�d<��^<P�Y< 6U<�qQ<BN<��K<�I<��F<gD<A<ݐ=<�k9<��4<5�/<�,*<��$<��<4�<Nw<�'<7�<Uw	<��<���;l��;5��;6��;���;�|�;�;�A�;���;as�;�o�;T6�;���;��;{��;5^g;��M;B�5;d�;}*;��:>�:�:2s�:S1�:D��:�M�:4��:��:-��:(�x:`�Q:"�':�g�9��9ge9��9�΋8��7��ϷrT���
���T�M������ݹn���� �/% �����i,��$' � ���4$�'�E��\p�`>��dA��Ol���׺���@���X���U�������`�������^�ݺ]ٺ1�ٺ�]ߺ+꺑��K����£��	��� ���$�I�'��`+�6l/�;k4��@:��t@�mF�K�K��:O��iQ��dR�S��RT�TIW�I�\�r�d�8
o��m{��s��v@�������Y�����=�����!���l��޶�� '���  �  �=I�=|l=0=��=�=́=i� =6� =V =�. =� =r��<���<#�<�a�<5n�<a�<�Z�<y�<���<�r�<�I�<8�<��<Q��<��<�<H��<-�<bC�<�u�<r��<�[�<�H�<b��<�i�<��<{�<���<�h�<�<�j�<�}�<�3�<A��<���<��<���<X��<)-�<!��<5��<Z��<-t�<X$�<���<��<���<���<v��<��<\�<Ο�<�C�<���<�M�<�d�<t�<;?�<W�<�m�<��<���<���<�O�<��<���<�S�<���<���<���<���<���<[�<���<��<?!�<�~�</ų<��<ӟ�<�a�<]Z�<;s�<X��<W��<�X�<��<s>�<�u�<���<��<��<E{�<���<��<�F�<�r�<5U�<�ل<���<Ԗ}<B�v<m�o<.�h<�/b<0\<|�V< �R<O<�#L<F�I<՞G<�uE<	C<�@<�`<<�8<�$3<��-</�(<d#<f�<�j<t�<��<y	<"�
</n<�k<O�;-��;S��;0��;�Q�;9�;|�;�s�;���;���;$�;�Ɩ;��;��|;��a;��F;'[-;�;��;'��:�9�:7�:��:I��:���::�:37�:��:8�:��b:9:dv:YN�9]�9+M,9G<�8έ�8��8�f]8��7�"�~���m�Ӯ��g湺������.����Ј����&� ��T5��V�ཀ�YY���̵�|�к8麦.������C	���	�d�8���������e��gr�W�⺛��z������j�����kt������!���"��
$��%��E)���.���5�t�=���E�mM�DS�yW���X�*�Y��Z���\��Ha���h�ps�$���(��o���ĕ����>!������DR���n���=���(��ɳ��3o���  �  AA=_J=�=��=B=�=3=Ѣ =;R =N+ =S$ =�+ =�, =T =���<���<&��<s~�<d7�<�<;�<մ�<�z�<�j�<�W�<��<��<2��<�+�<�|�<`��<���<h��<�T�<0�<1��<>Y�<���<�4�<���<���<D|�<3��<��<���<i��<��<��<}��<��<���<���<ή�<n��<��<g��<��<�:�<�<���<x�<AT�<:r�<9��<Hp�<��<���<6��<.y�<ճ�<�s�<���<=��<���<���<�9�<���<+��<�B�<��<��<�/�<�H�<�1�<0;<	�<�ܺ<�^�<���<�<�T�<���<w��<l,�<���<	ۦ<��<1�<sh�<���<���<ϡ�<o��<2�<>ˏ<=ڍ<'�<5��<�Ĉ<���<�P�<0y�<��|<��u<�;n<�g<�0`<�Z<^�T<BaP<��L<�VJ<27H<�PF<�QD<v�A<)�><4';< �6<!�1<#=,<w�&<��!<ێ<��<�a<�*<��<��<�<j<�w�;�w�;�z�;�*�;`�;]_�;Y��;XX�;���;�l�;Iޞ;u��;v�;�%x;��\;M�@;�2&;��;�`�:�h�:H~�:?ܩ:1�:���:gY�:N��:��:B�:��r:
RL:M :oB�9
��9�79ą�8p�8�h�8$ �8#��8PG�8$��7�{��*�K�����K�����)�c�1�p2��.��-���4�1BG���f��G��0ܣ������޺y����	�~�F����C������W����Kj�����A���� ��^	�3�����a�S="���"�K:"��!�4"��%�R�*��q2��<��\F���O���W�	�\��8_�T`���`��Bb�$f�hm��Cw��%��Ȩ��𓑻*@�� ��ir��������s���Ȩ�-��H?��Ǧ���  �  �=�=s�=�=��=�`=�� =�^ =� =+	 =D =�4 =SF =s8 =���<��<���<s��<a�<���<[��<�(�<���<D��<C��<n��<��<3%�<n��<a�<�%�<�%�<�A�<R��<%t�<��<1��<<��<O��<(��<ta�<9�<O��<>��<��<tU�<�N�<?7�<�A�<��<}Q�<�_�<O��<k��<��<)��<hi�<ex�<�3�<���<cF�<e��<I��<�C�<���<>~�<��<CD�<%�<2N�<��<�_�<�h�<S�<�L�<x��<�<��<N��<�d�<_�<ô�<���<�˿<�e�<L��<(^�<�з<O�<GT�<oï<���<ٟ�<D�<`��<�<�D�<*.�<���<�ٝ<��<g��<�{�<��<9H�<�F�<Ր�<W��<(E�<�K�<��<��<��{<��t<�:m<Q�e<��^<��X<:5S<��N<��K<D"I<�,G<]iE<��C<x%A<�><�@:<&�5<ax0<m
+<��%<�� <ٷ<�8<�2<+Q<�5<�<+<��<;�;���;7�;g�;�U�;�@�;i��;��;G��;���;�5�;T=�;Ӕ�;[u;�Y;��<;4g!;��;+��: ��:bN�:3��:Z�:��:[��:���:y!�:@؁:(bd:��;:�0:�c�9If9{O�8��~8��c8n��8���8�i9+��8�k�8��'��:������= ��"�@%9�5D��E�V3A�4�>���C�/�T��s�Lo�������Ⱥ���&]�����k�w���k�|��>�H���������W�y�z���*(�=�/��]��#���$��$�""��K �� �W�"��2(�|�0��m;�R�F���Q��Z�P�`���c���d��'e�?Of���i��Hp�IOz�����ef��]�����������2U��������A#���'��38��|���;���  �  ��==��=�l=��=(E=,� =�E =B =���<) =�6 =gN =1D =�	 =�5�<���<߈�<��<R��<��<���<��</��<(��<l�<���<� �<��<:��<���<<��<�<�g�<x1�<k��<�b�<g��<�q�<nU�<�:�<_��<�_�<a�<���<�$�<��<^��<��</j�<�-�<kK�<>��<&��<�-�<��<u��<6��<}=�<���<x3�<���<3��<k�<:��<~G�<���<��<{��<^)�<���<U8�<<�<��<��<?�<���<���<;L�<�+�<iM�<V��<���<���<�?�<Mm�<0�<��<Q۴<Q�<���<<W�<��<H�<���<T�<�Y�<�G�<�ʠ<W�<�ƚ<���<�d�<�<Y�<]�<�Y�<UÉ<e�<�"�<�ƃ<��<�q{<�St<U�l<Sqe<$d^<X<s�R<�dN<�$K<Y�H<��F<\E<�6C<�@<�=<��9<)F5<�0<W�*<xK%<H} <gf<z<�<�Z<�W<��<�`<�)<x�;f��;\��;��;(��;\w�;�ո;�9�;�֫;gۤ;ܚ�;��;T�;��s;�W;�H;;��;��; ��:,��:Y�:�$�:V��:\W�:�d�:Ac�:���:�:�_:�5:p�:Љ�9b9K9��8c78�;83͡8ڗ�809��	9쮛8����#�5�/������O&���>���J�iL���G�Q�D�I5I�UY��w������qO˺�꺋%������i��^�P8����Y�\q ������Y�����q��G��N����� �Jv$�&�%���$�""�����q�]�!�s'��50�E>;�X:G�a�R���[��Xb��e�s�f���f���g��k�/sq��i{��H�����K��=g��'���Z[������������n����層٣���͢��  �  �=�=s�=�=��=�`=�� =�^ =� =+	 =D =�4 =SF =s8 =���<��<���<s��<a�<���<[��<�(�<���<D��<C��<n��<��<3%�<n��<a�<�%�<�%�<�A�<R��<%t�<��<1��<<��<O��<(��<ta�<9�<O��<>��<��<tU�<�N�<?7�<�A�<��<}Q�<�_�<O��<k��<��<)��<hi�<ex�<�3�<���<cF�<e��<I��<�C�<���<>~�<��<CD�<&�<2N�<��<�_�<�h�<S�<�L�<y��<�<��<P��<�d�<b�<ƴ�<���<�˿<�e�<P��<,^�<�з<S�<KT�<rï<���<۟�<F�<b��<�<�D�<*.�<���<�ٝ<��<e��<�{�<��<6H�<~F�<Ґ�<S��<$E�<�K�<��<��<��{<��t<�:m<N�e<��^<�X<:5S<��N<��K<G"I<�,G<aiE<āC<%A<�><�@:<.�5<hx0<t
+<��%<�� <߷<�8<�2</Q<�5<�<+<��<;�;���;/�;]�;�U�;�@�;[��;��;8��;u��;�5�;E=�;Ŕ�;Au;{Y;x�<;!g!;x�;��:��:ON�:$��:N�:��:T��:���:u!�:>؁:%bd:��;:�0:�c�9Ff9xO�8��~8��c8n��8���8�i9,��8�k�8��'��:������= ��"�?%9�5D��E�V3A�4�>���C�/�T��s�Lo�������Ⱥ���&]�����k�w���k�|��>�H���������W�y�z���*(�=�/��]��#���$��$�""��K �� �W�"��2(�|�0��m;�R�F���Q��Z�P�`���c���d��'e�?Of���i��Hp�IOz�����ef��]�����������2U��������A#���'��38��|���;���  �  AA=_J=�=��=B=�=3=Ѣ =;R =N+ =S$ =�+ =�, =T =���<���<&��<s~�<d7�<�<;�<մ�<�z�<�j�<�W�<��<��<2��<�+�<�|�<`��<���<h��<�T�<0�<1��<>Y�<���<�4�<���<���<D|�<3��<��<���<i��<��<��<}��<��<���<���<ή�<n��<��<g��<��<�:�<�<���<x�<AT�<:r�<9��<Hp�<��<���<6��<.y�<ֳ�<�s�<���<>��<���<���<�9�<���</��<�B�<��<��<0�<�H�<�1�<6;<�<�ܺ<�^�<���<�<�T�<���<|��<p,�<���<ۦ<��<1�<rh�<���<���<ˡ�<j��<,�<8ˏ<7ڍ<'�<.��<�Ĉ<���<�P�<)y�<��|<��u<�;n<�g<�0`<�Z<]�T<DaP<��L<�VJ<:7H<�PF<�QD<��A<6�><B';<�6</�1<0=,<��&<��!<�<��<�a<+<��<��<�<j<�w�;�w�;�z�;w*�;J�;D_�;>��;<X�;i��;�l�;,ޞ;Y��;[�;p%x;[�\;#�@;�2&;��;�`�:�h�:"~�:!ܩ:�:䙜:ZY�:D��:��:B�:��r:RL:M :jB�9��9�79���8o�8�h�8% �8$��8QG�8)��7�{��)�K�����K�����)�c�1�p2��.��-���4�1BG���f��G��0ܣ������޺y����	�~�F����C������W����Kj�����A���� ��^	�3�����a�S="���"�K:"��!�4"��%�R�*��q2��<��\F���O���W�	�\��8_�T`���`��Bb�$f�hm��Cw��%��Ȩ��𓑻*@�� ��ir��������s���Ȩ�-��H?��Ǧ���  �  �=I�=|l=0=��=�=́=i� =6� =V =�. =� =r��<���<#�<�a�<5n�<a�<�Z�<y�<���<�r�<�I�<8�<��<Q��<��<�<H��<-�<bC�<�u�<r��<�[�<�H�<b��<�i�<��<{�<���<�h�<�<�j�<�}�<�3�<A��<���<��<���<X��<)-�<!��<5��<Z��<-t�<X$�<���<��<���<���<v��<��<\�<Ο�<�C�<���<�M�<�d�<u�<<?�<X�<�m�<��<���<���<�O�<��<���<�S�<��<���<���<���<��<#[�<���<(��<I!�<�~�<9ų<��<۟�<�a�<cZ�<?s�<[��<Y��<�X�<��<p>�<�u�<���<��<��<={�<���<��<�F�<�r�<+U�<�ل<���<Ė}<4�v<a�o<$�h<�/b<0\<{�V<"�R<!O<�#L<Q�I<�G<�uE<C<�@<�`<<�8<�$3<��-<A�(<d#<u�<�j<�<��<~	<%�
</n<�k<D�;��;<��;��;�Q�;�8�;V�;�s�;y��;���;��;rƖ;l�;x�|;[�a;u�F;�Z-;�;��;���:n9�:�:��:0��:u��:+�:)7�:��:8�:��b:9:av:UN�9[�9)M,9E<�8έ�8��8�f]8��7�"�}���m�Ӯ��g湺������.����Ј����&� ��T5��V�ཀ�YY���̵�|�к8麦.������C	���	�d�8���������e��gr�W�⺛��z������j�����kt������!���"��
$��%��E)���.���5�t�=���E�mM�DS�yW���X�*�Y��Z���\��Ha���h�ps�$���(��o���ĕ����>!������DR���n���=���(��ɳ��3o���  �  B�=�= �=�p=1=�}=��=,Z=� =�x =C+ =���<�i�<M��<&^�<r��<��<?�<e�<H��<�g�<2�<Z�<��<���<�d�<���<��<�6�<��<���<U\�<���<���<X��<���<#��<1��<��<g��<��<���<���<f�<J��<D�<ds�<�t�<�h�<{o�<���<��<΍�<�/�<���<d�<���<C&�<M`�<*��<R��<-:�<���<@k�<A�<Ȱ�<��<��<Ü�<��<���<��<}r�<r��<q�</��<jV�<U�<=��<� �<���<���<��<�N�<G�<�5�<5�<��<�T�<0��<��<�?�<Ĭ<�q�<�<�<>�<^ߣ< ��<q)�<4��<��<j��<�=�<��<
*�<�l�<k<T�<��<q�<q[�<:|�<�~<x<beq<��j<7�d<��^<O�Y<#6U<�qQ<BN<̄K<�I<äF<{D<"A<��=<�k9<ղ4<M�/<�,*<��$<��<D�<[w<�'<>�<Yw	<��<���;^��; ��;��;���;c|�;��;hA�;Ɛ�;/s�;�o�;!6�;Q��;R�;P��;�]g;[�M;�5;,�;N*;���:�=�:��:
s�:31�:,��:�M�:(��:��:'��:�x:Z�Q:�':�g�9��9de9�9�΋8��7��ϷpT���
���T�M������ݹm���� �/% �����i,��$' � ���4$�'�E��\p�`>��dA��Ol���׺���@���X���U�������`�������^�ݺ]ٺ1�ٺ�]ߺ+꺑��K����£��	��� ���$�I�'��`+�6l/�;k4��@:��t@�mF�K�K��:O��iQ��dR�S��RT�TIW�I�\�r�d�8
o��m{��s��v@�������Y�����=�����!���l��޶�� '���  �  ��=�=�=ܬ=LN=��=�;=y�==`� =B =9S�<T��<���<�Z�<2��<�+�<���<?�<��<r��<��<7��<���<�a�<��<s�<���<���<�<,��<~<�<p��<���<���<�b�<��<���<��<qA�<���<|��<K?�<[�<q5�<;��<�<C�<��<;��<���<� �<�:�<��<���<Vf�<Q��<�E�<��<�:�<&��<|�<W?�<_�< ��<YQ�<���<�w�<���<�!�<K��<���<[6�<̾�<�Q�<���<���<���<.��<VK�<���<e�<��<���<qA�<���<���<}w�<���<iM�<*��<���<���<�Y�<�ҧ<�^�<���<���<�.�<%қ<���<QT�<*H�<g�< ��<
�<7b�<S��<���<�E�<���<)ς<��<�By<��r<��l<�g<k�a<��\<� X<��S<@gP<h7M<�PJ<{�G<��D<��A<�[><�e:<��5<��0<�y+<��%<Dt <j!<N<�<�?<k~<<�<��;���;S��;+�;:�;���;�5�;���;��;��;�;���;�֙;�N�;NG�;�Zl;ѼT;�S>;�);l;;I�:���:��:-ǿ:�:�D�:�Ӧ:��:Tʒ:=+�:x�d:Y�;:�7:��9�Ń9ܲ9l��7��t�<��_�K��C���֢�m&��3ҹu�߹S�����,ٹ$Oѹ+Eѹ�L߹�l���Y��;��d��ׇ�}���Z1���xĺz�ӺJߺZ��E�꺌������%�ySݺ��׺=ԺԺ\jغ����o����	�	0�����!��*(��-��2�w�7�,7<�]�@��D��uH��K���L�(M�%PM�6�M�F�O��pS��Y���a�^l�Rx����u�������r���{��B����������F᜻1j���~��g���  �  *�=/�=S�=��=sm=��=g=!�=�=�o =��<���<D��<���<<!�<���<S6�<S��<���<5��<"��<��<��<���<M��<���<y
�<���<���<�Z�<��<k��<V��<�<�W�<_��<�O�<N�<s��<���<��<��<�G�<_�<�H�<���<lS�<|q�<�Z�<�%�<J��<ɾ�<ɫ�<���<T��<@2�<���<�.�<���<H��<���<{�<u�<`�<I!�<C��<=��<B��<��<K1�<�&�<���<��<��<`o�<mL�<�5�<�.�<T:�<�\�<Ș�<E��<y]�<���<�P�<m��<VҼ<{��<�R�<8��<ֲ<��<��<�<�-�<�r�<�ա<�X�<���<�ǚ<���<�і<��<{r�<Q�<!Z�<ΰ�<PԌ<���<!P�<���<�؂<��<iz<�Ft<s�n<CUi<>2d<*O_<ȯZ<cZV<"SR<ЛN<�/K<<H<��D<�A<i�><A�:<>e6<�1<,,<�{&<�� <d�<�<��<�1
<�<�> <�S�;ܾ�;���;nl�;&��;BO�;k.�;���;���;�8�;�b�;^��;�;�}�;P�;��o;`SZ;"F;�3;͝!;��;۩;ұ�:<��:���:=�:��:8��:q�:���:���:\�l:(UF:3:`K�9��9�M�8C|3�6B*�0_���F���ӹ4鹊[���P������I8չG�Ĺ�������'iӹ�	�����n�:��)`��􂺉ה�:���U��w���oɺ�AѺ�ֺmhں��ۺEۺ30ٺ�Rֺ��ӺY�Ӻ�ֺ#3޺ ?�sX��W��9��L��$��r-��'5���;�6JA���E�(I�<@K��gL���L�"L�+K���J��=K���M�N<R�`Y���a���k���v�����+~���򉻙ߍ�a>������N��% ���"�����Gܙ�ߠ���  �  ��=��=u�=2�=k\=*�=he=�=v� =�9 =���<u��<�o�<�x�<���<�K�<w�<��<�:�<�}�<��<@�<�<��<<r�<L��<��<��<Vh�<!M�<�Q�<z�<���<�<��<���<o�<q��<H��<y-�<���<���<H��<�<���<��<�9�<�j�<�U�<|�<j��<\=�<���<˯�<��<���<�D�<��<���<��<���<�2�<[�<�]�<��<���<��<1Q�<g��<���< �<�<�'�<lC�<�^�<s�<py�<�n�<uW�<m>�<l0�<�9�<rb�<\��<3�<`�<"��<���<rI�<Y��<\Բ<Hů<Û�<�o�<oT�<�Y�<Q��<���<���<���<���<��<���<�3�<�Α<�P�<���< ��<�v�<���<�P�<��<5�<�=z<�u<* p<xJk<��f<��a<g]<dX<�S<��O<��K<�G<dyD<;A<��=<H:<2*6<v1<�*,<�^&<b; <s�<��<��<��<�b<���;h��;��;}	�;��;[��;�y�;W��;J��;Ǖ�;4p�;u2�;	�;�J�;�d�;�;�;q;�'^;p/L;�*;;��*;S;�j;���:[��:���:sk�:��:xơ:�@�:\��:o'�:�?i:�E:94:�Q�92�d9г8����z����ع�#��<����D��<��͌
�������ܹ��ƹ?����Ĺ��߹wB��#���D�g.f�偂��珺0M��i���˭���������ź�ͺ�ӺEb׺��ٺ��ٺ ,ٺ"�غ�ۺ���V^�A�������@���z)��\4��>��F�oBL��lP��R�.S�% R�v3P�D�M���K�`�J�H�K�ΜN�hT���[���d�f;n�c�w�����ۃ���*���ڟ���&��ܡ��<���,������E������  �  e�=y~=�q=�W=)!=��=<=&�=x� =e��<-#�<���<�.�<�<�U�<n��<?��<&�<Aq�<P��<�^�<c��<
��<���<���<B�<��<<��<g��<|��<5G�<���<�T�<���<��<=��<X�<]��<���<	F�<���<�}�<�a�<�a�<^�<y5�<>��<��<��<J��<�'�<K��</��<���<=Z�<�p�<&��<���<���<5��<K�<��<���<��<���<I'�<�<˺�<��<nV�<���<���<�@�<L��<�<>b�<ʅ�<�w�<�<�</��<���<�B�<�"�<�4�<mr�<�ý<��<��<��<�c�<���<�d�<�<#��<�Z�<9*�<Q5�<���<�@�<�J�<��<�5�<��<ฒ<9p�<���<@�<�7�<d�<QV�<1��<:��<��~<��y<�lu<�q<��l<�oh<��c<n_<��Y<&�T<��O<4_K<�*G<iC<*�?<��<<V09<�E5<��0<}�+<ұ%</X<|�<��<�s<�A<(&�;��;xf�;2�;��;�p�;I��;ǥ�;pW�;�-�;f�;sX�;q��;xQ�;���;�,�; Z�;��p;\`;��P;�A;��2;\/#;J~;�;��:5��:#з:���:��:���:Wm�:l�t:E[:ć9:��:X)�9'#$9�0X�@6��)��S��:2��|B�!G�p�A��4�f!�V��w���6۹�ӹV�߹ � �'��l8��$X�P
u��;���펺$B���\��臟�X饺�/��kE��Uú�-κ��׺E޺h��D*��W���交�躖�����i�	��R��L"� �/��F<���G�X�P��W��[�\�\�~�[�TY��VU��Q��N��RM��qN�09R�{}X��`�V�i�h�r�G�z������1��H1�����%ۈ�����΍��搻���)��ʳ�������  �  �1==�=��=;�=�z=��=�L=�y =� �<D�<ҁ�<���<b��<���<5��<ǰ�<E�<?��<?�<f��<.�<�<�<���<F�<�U�<L=�<}$�<N1�<�}�<�<x��<���<���<�A�<���<o�<��<��<�.�<h�<���<f��<8��<��<{�<�*�<��<ǂ�<(�<X��<��<��<�s�<��<s�<��<�[�<��<���<|��<M�<gw�<���<!F�<���<�i�<���<K�<���<���<#~�<])�<j��<@��<��<�R�<�A�<0��<�U�<��<��<���<���<T��<S��<�F�<�r�<nY�<��<��<�ݮ<}p�<��<�_�<��<��<-8�<4�<	�<ԍ�<�N�<5�<��<!�<$s�<ܫ�<ǌ�< !�<P��<qӃ<s9�<�}<Py<`u<��q<��m<B�i<ke<�{`<�$[<��U<hP<�J<� F<B<3g><�;<�7<��3<x�/<�*<��$<42<�J<�=<.T	<��<?��;`��;�!�;O=�;Z��;	��;Ѵ�;�H�;n.�;��;,d�;�y�;�|�;��;QO�;	M�;T�~;C�n;��`;6QS;B/F;�I8;�$);E�;��;���:��:�t�:;w�:FZ�:��:�n:T]:��F:w�':�`�9�9@0�8�t�<#������H>���\��(m��oo�9�e�2�R�06:��� �	u�w��z���ɩ���rj3��R��q�ު��t���됺Ej������������Q0��sP��m���%g̺ՎںZ��M�캌��I��!���� S���*������?�'��6��5D���P�'[��Rb��f�0�f��Od�)`��[��;V�>�R��dQ���R� qW�uz^�n)g��Rp���x��[������I�����؄�������%m����咻���Oٚ�y����  �  !�=3�=d�=��=�u=�.=��=�	=j2 =g|�<<��<G��<���<���<N��<ϑ�<��</�<���<w��<�D�<{��<��<KR�<ԓ�<���<�l�<aY�<��<M��<%��<���<���<���<���<�G�<z�<gh�<\2�<� �<`��<�@�<��<��<0��<���<��<
��<��<ڠ�<���<o�<�?�<Ʉ�<r�<^�<8m�<dO�<��<&�<���<�}�<1��<��<���<b��<T��<9-�<�<
��<EW�< �<3��<���<T��<ތ�<���<���<W�<Ǘ�<��<���<u=�<��<��<�-�<y��<ĸ< ��<�[�<���<�W�<'ت<�/�<�<��<ޜ<��<Z֗<%
�<���<u��<���<ъ�<�^�<u�<��<�ފ<$^�<r��<}�<{{�<xv|<z�x<� u<}�q<�n<��j<~�f<H}a<�[<��U<�O</J</E<��@<��<<#}9<�76<��2<2v.<�y)<��#<<C<��<��<a� <�l�;��;���;�2�;X�;&��;��;���; ��;���;Vط;H��;eM�;�;
�;Hq�;�;z;O,l;`;Z�T;�0I;5<;<-;?;�	;���:���:�n�:<�:W�}:N�e:��T:8?E:�1:39:0B�9t�q9-�!7��n�)��E�1�j�_����WQ�����
���Z�l�`P�j�3��|�x��(����`�.�Z�L��l�9Մ�%������A��N�������l捺�L����������X����̺��޺7��8���p}������@���`O��ן�������I�&g,���;�uK�A�X�0�c�!5k�)�n���n���k�*^f�HS`�'�Z�@�V�ƦU���W���\��yd���m���v�n�~���o��{ȃ�v���K~�����ⅻN���;>��:I��I����<��S����  �  ��=�c=�U=�N=6=��=Z�=4� =%��<�
�<Y��<C�<�J�<;��<�#�<���<-�<��<)a�<�1�<���<�F�<�I�<��<m�<���<)��<���<���<��<��<��<���<�(�<��<ו�<ͻ�<��<�4�<1��<��<���<�K�<�%�</�<�6�<a�<6��</��<?�<��<&��<y��<���<u_�<�F�<��<��<6��<���<*^�<��<%��<ë�<�O�<Jv�<,/�<���<D��<	H�<���< ��<���<I��<}�<���<�2�<>�<���<ٸ�< ��<��<���<8n�<�\�<K��<���<�C�<�N�<���<�,�<0��<gm�<���<u��<+f�<�'�<�]�<��<�Z�<��<���<8�<"�<��<䀎<���<�_�<�χ<��<Li�<>�<�{<��w<H�t<��q<`�n<{ek<� g<6b<6K\<cV<��O<�I<y3D<��?<�;<�R8<� 5<��1<�-< �(<��"<�J<�<,�<�Q<���;Vy�;�;���;��;���;D��;!S�;I]�;�e�;��;��;�~�;���;�;7��;T�;��v;]*j;�n_;�sU;7�J;q>;�/;t8;��
;W��:=3�:��:��:z�k:�eR:��A:��3:�":)�:�=�9a@9�+�pv����
�*�E�ev��狺�-��;Г�o"��v~�!�_��)A���(����o ��'���?�oA_�	��N荺̪���{���'���֑��x��)x���;��;������fOͺ�P⺺�����������g\�V��bF������� !���/���?���O���]�!`i�('q���t�[.t�mp��j���c���]���Y���X��[��`�/�h��Rr��{��z���Ƀ�2����F���i���Ă����D����ڇ�|w���
���ꗻ=W��P����  �  ��=�M=I=��=׬=�O=��=2(=b =��<�M�<���<u-�<r�<�B�<W��<���<� �<��<��<v��<���<&��<��<��<1�<U�<��<P��<�O�<��<���<��<���<3��<��<�>�<G�<�1�<��<))�<�h�<��<s��<)@�<���<�s�<��<F��<�d�<*��<m2�<T��<���<c��<ɪ�<�
�<	��<}��<�"�<���<^��<w&�<��<���<P�<n��<_��<IB�<���<�j�<x'�<1 �<x��< ��<�H�<���<���<J�<Ҿ�<�<�n�<���<A��<���<ꑼ< ��<���<tv�<���<�3�<;!�<$ת<�p�<��<�Р<�ם<Z6�<p��<C�<���<�?�<0�<H�<&��<��<H�<�:�<��<���<� �<Gʁ<	><	Q{<շw<�Bt<�p<k�l<�}h<��c<�L^<j�X<sS<�M<ŀH</�C<��?<��;<8<�4<x/<�X*<Ϝ$<hW<�<R�<@
<��<��;���;Q1�;�A�;���;6��;��;T�;$��;��;�<�;�ѳ;���;�"�;×;0�;��;�;`s;�tg;�I[;@N;�|?;�^/;�4;��;�#�:'�:���:��:���:�V�:|��:��h:�F:�4:P��9YQX9�~;�vk��p۹R���R6��H��%M���F���7��$�L������	깇�繝M�������"���:���P��b��/l��o�sho���n�;rq�U�z��"��Jᒺo�������.ĺ�LҺ��ܺi�ܛ�QG��W��Ĕ��C�����G,��'�A�4��)B�s4N� X�]�^���b���c�'5b���^���Z���V��$T��kS��U���X� �^�.�e��l���r��w�B�z��?|�Z�|��}��������>󄻕ֈ�7V��y����U������  �  ��=�]=N/=)�=I�=S`=b�=�7=(r =1�<�s�<3��<WZ�<$7�<�q�<��<�<�I�<��<�;�<Q��<���<���<[��<i�<�U�<fx�<��<���<�_�<��<���<���<���<�l�<���<O(�<q6�<�)�<N�<�4�<�}�<m��<@��<�d�<��<��<\��<r��<��<���<�U�<S��<�#�<���<���<�9�<���<��<KJ�<O��<�<�E�<[<�<l��<�(�<��<C��<�c�<���<��<;3�<��<��<1��<�1�<F��<��<4�<k��<z�<�r�<p��<���<��<߳�<�˺<E˸<���<��<�Q�<C@�<��<���<�5�<���<��<te�<Z%�<�D�<��<wf�<N5�<%�<ڴ�<q0�<Ii�<^�<��<���<�A�<b�<�d<#d{<3�w<�-t<=�p<�l<�Ih<oc<&&^<b�X<"S< �M<��H<�$D<@<�7<<�^8<\F4<�/<*�*<��$<��<��<56<�
<�Q<3G�;4X�;1��;L��;�4�;�@�;r��;��;�s�;%�;�ż;ec�;�;�;!��;!C�;hX�;IA�;[�;Es;�g;�Z;1`M;��>;?�.;s�;T�;�E�:2��:�C�:G��:�:���:�ׄ:�&m:�J:$!:���9��h9_�6��W�n�й��go0��5B��iG��fA��2�H��z��,��~@��߹���^9�XH���6�VM�8G_�	�j�J�o��Sp�9�p��-t�J�}������,���|�����S�ú{^Ѻ�ۺ?��lk���뺧�}�����b��}.�V&��3���@���L�o�V�e�]��ka�hb���`���]�-�Y���U��+S��pR�<T���W�5�]���d�P�k��r��)w��tz�8F|�ZR}��~�Cf���`��ER���!������L��Z4�������  �  ʼ=��='_=�/=�=�=	=b=$� =Y��<��<!A�<���<���<���<���<B��<��<�!�<��<'�<B�<�D�<v �<w�<���<��<'��<')�<���<��<���<}��<<z�<L#�<��<p��<J�<R�<O �<�R�<��<�L�<x�<K��<�r�<8��<1�<)'�<7��<�V�<��<}�<��<�W�<qa�<���<"x�<�{�<J��<1�<g�<4��<ԏ�<W5�<���<�|�<3�<���<�7�<��<�Q�<��<���<i�<���<j1�<�1�<0��<��<���<�y�<F�<C��<a�<��<�)�<r'�<��<�o�<0��<���<�R�<��<���<�w�<���<F�<���<Tŗ<.�<SҔ<떓<,^�<+�<(��<oÍ<���<�{�<��<̛�<|0�<_�<g�{<1�w<5�s<�p<kl<'�g<�b<��]<�LX<��R<!�M<� I<�D<��@<v�<<19<��4<�h0<w@+<�%<XG< �<�
<%�<�R<yh�;,��;E�;.��;l
�;���;$�;g@�;���;>��;�:�;��;,ˬ;�9�;2��;Ip�;��;W�;��r;�e;��X;k&K;k<;��,;,;ǽ;�s�:���:'��:{��:Y��:4Ǘ:��:��x:q�U:3�+:�F�9��9�^8n� �t�����h�.$1�P7��)2��%��)��Q �q���͹��ɹ��ع���.�:+��PC���W�of���n�W]s���v�{|�N���NR�����%;���)��86ú�κ�u׺Hݺ�������.�P������w1��{�Q/#�x0��]=�>�H�ylR�b9Y��3]��f^�,3]��LZ���V�S��P���O�6<Q���T�z�Z�υa���h�l�o�Ջu��y�\r|�|Z~�!"��������Rp��%�����O*���ᕻh蘻�  �  ��=3�=��=Zp=C+=��=iA=Ϛ=}� =} =Vv�<0��<L��<-��<}��<a�<�A�<Re�<��<	�<�x�<ֲ�</��<Sw�<���<�8�<�V�<�g�<P��<q��<3+�<M��<�f�<��<���<��<2q�<E��<D��<��<}w�<��<Ѷ�<3��<gG�<���<l�<0��<G��<8L�<a��<uD�<l��<�P�<��<3�<��<z@�<[2�<�Y�<���<���<y�<8��<إ�<q��<���<!��</7�<j��<.�<]v�<���<���<N�<u�<$��<1��<J�<4,�<���<z�<wJ�<�D�<�_�<ވ�<6��<t��<hb�<Uݴ<&�<��<lѫ<���<OK�<M2�<�T�<���<�}�<���<�ߖ<�o�<�!�<[ڒ<��<���<c:�<�:�<���<\��<<�<W��<,�<��{<g�w<\ps<1^o<!&k<�f<��a<��\<9�W<_�R< �M<{I<�mE<8�A<"�=<N:<%�5<P1<,<{d&<l8 </�<j?<��<>�<eY<���;�Q�;���;6��;�Q�;�D�;*/�;Z��;Gc�;�)�;��;�;�J�;��;8�;��;��;T�q;��c;=�U;OdG;�8;�");s};6
;��:pa�:��:`W�:���:k�:z�:W#�:Lwd:d
::\�	:�{�9�r�8�%������ѹ����]���<����Q�e��ù��?��뛺���ع����i���5��M�KEa��jo��Ky�v���N������k ��4���-��$�����º�˺��Ѻ�1ֺ��ٺ��ݺ�G��Y�!���f��p�� %�v�+�/%8�C��L�-�R�?�V��HX��W��oU��QR��6O�s�L�\DL�ƗM�Q���V�y]��e���l��gs���x��}�	!��ɡ���\�������S��񔋻(�����������旻�  �  h=� ='�=4�=wg=��=�w=�=C=ZU ='�<���<y��<��<��<�^�<v)�<�.�<�`�<��<���<�!�<�"�<S��< o�<���<���<���<���<��<�&�<���<���<�z�<=��<=l�<c��<�'�<&��<c��<���<IK�<��<���<���<rp�<���<��<�<��<1W�<��<ou�<@+�< �<�6�<���<
7�<��<{�<^=�<�h�<��<i�<��<�j�<�r�<\/�<s��<�<�K�<��<��<�3�<���<���<���<���<���<e��<���<�h�<nm�<��<�ɿ<k�<-"�<��<�Ϸ<eE�<�z�<{�<LY�<:-�<��<L�<�O�<�ǝ<[��<{�<���</&�<�<�\�<��<�i�<2��<<���<��<��<���<�k�<��{<r2w<^�r<�En<��i<YBe<ь`<��[<��V<�MR<��M<��I<�$F<r�B<��><@;<q�6<o,2<��,<�C'<33!<��<У<4�<ֻ<�b<��;W]�;V��;��;��;��;�1�;���;�0�;@�;���;� �;�`�;lc�;d�;}��;���;6p;fU`;�Q;EB; $3;/$;4�;ص;u��:^/�:>��:4 �:;��:,T�:�:���:��r:t�G:UX:c��9[6M9^lX7R�F1��v�ȹ!"�c���c�����ŒڹBt��bu��[��������p��>Z���i�W���=(��;D�Fm]�eNr�g���Q���N������t��}���Y�������uú�ɺ �̺*$Ϻ<�Ѻ�պ��ܺ�+纘����;��������&���1�p�;��.D�pkJ�S�N��P�>Q��O�:�M�3:K��iI�
�H�1J��ZM�%�R��oY��Ua�ېi��sq�)tx�CU~�y����̓�\����X������Ѝ�C���mH��El��
 ���  �  �>=N-=u= �=�=q&=��=!�=�M=�� =���<��<���<ʥ�<6��<yr�<[!�<���<t�<�*�<�U�<s�<�n�<8�<Y��<��<�6�<V0�<v�<��<P�<N"�<�`�<p��<Q�<o��<G��<�{�<��<ȼ�<0��<�v�<�k�<�X�<L)�<s��<�3�<z^�<HQ�<s�< ��<�u�<d3�<��<�<�R�<%��<B�<l��<4��<���<&��<��<Y��<tY�<*��<���<���<�<�O�<�t�<���<���<޹�<R��<\��<,�<��<��<N�<��<6�<r�<���<z�<�Y�<�z�<yh�<�<��<�Ų<�֯<�Ѭ<�˩<�ئ<z�<``�<g�<���<c�<���<�ݖ<lJ�<̓<�M�<���<���<m�<���<o}�<�<�B�<ӎ�<��{<��v<��q<��l<v#h<_yc<��^<�BZ<��U<k�Q<,�M<�J<�F<�3C<k�?<�;<N�7</�2<:�-<��'<W"< <�<c?<��
<��<�� <���;���;�d�;���;���;K��;���;I~�;d�;to�;(��;z��;ZӞ;�k�;��;!�;kpm;m�[;!5K;�i;;VG,;��;�S;
;���:{3�:���:9#�:'��:ғ�:��:��:@V|:��Q:'�#:��9Y�9[g�8M ��F#�߹����������1�ùH���]?�����Tx���!��ڒ}��#���̢�EV˹o �Jd��E>�37]��-y������(��9����䬺ݴ�(��>º�ƺ�HȺ�4ɺ�ɺn�˺ҿϺ�׺]4�;,�ƺ�)	������!�Q�+��Q4�ޡ;�QuA���E�6�H��J��(J�R9I�0�G���F��}F�E�G���J��O�ujV���^��_g��dp�n�x��U��Ĳ��A���rQ��ߋ��Z��#����ג������Ǖ�d����  �  6H=�?=S%=y�=�=1=;�=�=%n=V� =>9 =^h�<���<���<��<���<��<_��<w��<J��<M��<��<p��<TN�<a��<?�<�`�<�R�<%�<-��<���<s��<ԥ�<��<��<̄�<��<��<Wp�<�X�<�^�<qt�<Z��<���<+R�<���<�L�<.s�<�k�<,F�<B�<���<���<*��<� �<�l�<<��<J�<,��<;��<R�<�+�<g�< ��<�j�<r��<��<��<�*�<�e�<�o�<-Z�<�8�<T�<��<���<���<��<3�<�@�<��<���<�K�<h��<�-�<"{�<K��<^��<*)�<2��<�޲<��<>(�<UR�<���<�<�m�<��<��<�~�<�l�<ǁ�<���<��<y�<�Ր<��<(+�<�<��<��<YZ�<���<W{<O�u<WPp<�k<�(f<bda<R�\<`|X<�kT<I�P<�0M<��I<a�F<utC<�?<
<<��7<{�2<ǳ-< 2(<$�"<�<�A<��<j�<�<�<�%�;���;i��;�.�;�Z�;���;n��;'��;���;��;YP�;@��;6x�;޸�;Љ;~;��i;�$V;�)D;m�3;�?$;�W;�	;ɱ�:�	�:��:F��:��:NV�:�^�:�Q�:鱒:�C:�cU:ݢ):�x�9�ժ9�+D9��8�؄��;���p�����?*��q������y���Pv�us����8~���5����������>�1b�*q�����:����B������)���ú�*Ⱥէʺ�#˺�ʺ7�Ⱥ?�ǺDɺGKͺ2պ�����ﺑ� �SW
�9��I�r�%���,�I-3���8�g=��@�X{C�bE�b�E��E�F~E��E�G���I�n�N��U�;N]��f�.�p�߽z�m��(X������=�������P���3������j�������ǖ��  �  36=z4=�=:�=R�=4=��==�v=� =\v =Y =�b�<1��<D�<k}�<���<�i�<��<���<���<}�<�]�<�$�<���<�$�<�K�<:�<2��<��<G�<B��<~��<L��<�<�g�<���<���<K��<V��<I�<�?�<)h�<�k�<�:�<���<�$�<�I�<�K�<�>�<�5�<�B�<�l�<d��<]�<=p�<���<�9�<
��<��<ê�<�N�<
 �<b��<F>�<"��<���<���<��<�B�<�6�<q��<���<V\�<]�<���<0��<��<(�<�[�<���<�[�<���<C��<��<[^�<y�<�V�<>��<)l�<���<��<�S�<���<�0�<3å<�c�<a
�<���<�e�<\'�<m�<��<�.�<�n�<���<���<��<	�<��<L�<t:�<�K�<�z<P�t<I�n<�5i<��c<x"_<z�Z<�V<��R<�mO<�XL<|eI<gjF<q=C<Z�?<Q�;<;b7<��2<g-<�(<3�"<�Y<�9<KL<m�<_�	<|2<,� </�;oL�;��;�T�;�+�;S�;�}�;�X�;�;n�;���;�1�;n0�;�͈;��z;��d;c�O;�Z<;��*;Z�;�;�;LX�:���:[w�:���:�w�:�E�:�'�:f��:jh�:qkz:��Q:��(:Zo:#=�9q��9D�)9+U�8f�I7%�`�t���31��B^��{��5��\c�����^Ń����줢��1ǹ���I^��3D�دl�����Js�����建��ƺ-�κ��Ӻ��պxFպȐҺ!�κY˺\~ɺ*fʺ4�κpH׺�W��P򺬌��6
������:� ��R&��u+��R0�[5���9�e�=�4A���C��E���E���F�YH��K��{O��U�?�]���g���r��}�d���p���ڍ�}���t������=���Ø��̘�.^��eė��  �  }=�=��=i�=U^=��=�j=y�=�i=� =�� =XT =[ =*��<���<�Q�<˝�<���<hL�<���<Ns�<b5�<S�<2��<jd�<���<���<���<j��<�6�<���<4C�<U��<���<���<#I�<D��<���<���<�1�<Z��<���<��< �<���<u�</��<X��<7��<��<�+�<�o�<��<�Q�<���<�M�<z��<�<KG�<'��<���<4H�<���<�Y�<y��</<�<�a�<�:�<���< ��<4��<��<��<���<� �<$��<���<i��<P��<xm�<"	�<���<�~�<�-�<߶�<�
�<m�<@��<E��<�	�<qo�<�د<�V�<��<ʩ�<�o�<4�<H�<B��<{'�<b��<uc�<Z+�<��<5�<�c�<<��<���<���<�K�<��<M�<��<l�y<]Cs<�m<?g<��a<Q�\<�mX<_�T<Q<�	N<�BK<��H<a�E<�B<�?<�;<+�6<��1<ײ,<(�'<'s"<"�<��<�m<�<��<� <�I<m��;=s�;E�;���;���;U�;�0�;���;@D�;�ұ;Rq�;��;��;51�;�v;	_;��H;�b4;�M";��;e�;7��:P�::;�:*�:�::��:U˷:c�:.6�:D��:��n:J�G:]q":{Y:G��9S�9o�y9��:9,�8N5_8�v��A����&��a� N��W͐������_��w�����s[۹?�f/(��O���{��B��D˩��$�̺v�غ�w�AF�R;�:Ẻ�ۺ��պ��кOκ�)Ϻ�Ժn ݺ�`�����F~��P�g	�W��� ���$��I)�J6.���3�V9��?>�Q�B�+�E���G���I�r[K�=	N�61R�AX��\`��Rj�{�u�$񀻆��*�������nە���m������$��т��bw���a���  �  |�=I�=M�=�{=W=��=�/=��=�M=�� =P� =� =�W =� =��<2��<�&�<DH�<:s�<��<p2�<���<���<�B�<���<Z�<���<��<g3�<3��<p �<3��<��<���<���<�B�<���<���<�&�<���<0�<i�<���<β�<�w�<\��<�C�<�k�<v��<��<�<}�<H�<F��<�o�<���<Fc�<ޡ�<���<d��<R��<�$�<�{�<���<\�<���<>��<c��<L�<;{�<jW�<���<9c�<��<�9�<��<g��<ޱ�<� �<���<H�<��<���<c��<tC�<���<J��<[p�<Q�<m��<�<�<�<�<-�<:��<h�<%פ<�<^=�<g��<�+�<k��<�/�<��<ޑ<�<f�<+0�<�#�<q܇<iO�<�|�<z�~<�rx<��q<ׁk<~je<��_<�Z<�gV<�R<emO<-�L<J<]�G<��D<~�A<X.><�:<�5<B�0<��+<��&<k"<(�<P<A<�.<7�<�n<ס<�7�;b �;r��;��;k��;D��;/f�;�
�;c�;��;�˦;2~�;r<�;�C�;R�q;C�Y;p@B;8 -;^;^�
;l%�:��:��:92�:i��:���:H �:�-�:�_�:ͧ�:���::H_:��9:wV:,2�9���9���9~��9#��9��S9�<9�t8����� �/{W������U��,ͱ�6����gŹ�+عZd�������5�`�^�RF���]���Ե��ʺ�IܺM��\����h��Q��po��޺�غ�պ�ֺ�mۺU���w�A���-���4���
�������L�#�\�(���.�r�5�t<�:xB��?G��J�X+M�\O�8R�+ V���[�:�c���m���y��.������돻�e��ՙ����[���/����^���>��y����S���  �  ۛ=�=w�=�==s�=*k=��=��=�.=� =:� =ũ =-� =�[ =@ =rn�<ބ�<��<%��<���<���<�j�<�<'��<�d�<���<f�<��</��<�;�<ۖ�<z��<g�<��<��<�o�<C%�<11�<���<���<���<���<6:�<�@�<���<�z�<���<��<�<�_�<{��<�x�<B�<��<���<�y�<��<�<��<� �<9��<���<�'�< z�<P��<�2�<�^�<BF�<���<��<���<*n�<d��<�<�{�<��<���<4��<�4�<���<P��<���<Ss�<C;�<ξ<�<:$�<`�<��<\
�<��<A�<��<��<�2�<�K�<�J�< �<�<@&�<+u�<��<�#�<���<���<,��<���<��<M��<�g�<��<�<*�}<�kw<ȿp<�+j<�c</1^<(!Y<A�T<�Q<
N<�mK<�I<��F<�C<W�@<�==<� 9<\�4</�/<��*<M
&<��!<{a<�<��<U�<��<hu	<��<���;& �;�Q�;�(�;���;K]�;`��;��;;s�;x6�;+�;�Κ;���;�i�;��m;��T;V�<;�&;��;�3;��:��:���:!M�:���:�Ż:H�:\:�:��:ތ:Ou: �O: ,:M�:Z�9���9*�9�ʮ9���9�o�9_�O9�&�8�g7�aԸ��V�Ԓ���޸��E͹�ڹ(��l��(K��#���C��m�4���W�����/uֺ@��{(��P���������D���R(����aCߺ$ܺ�Mݺ�����w�������e
�����L��WX�v��}&������$�~�+�6y3�~;�#�B��I���M�+�P��^S��V���Y���_�jJg��Sq��E}�g>��'�������`�����Z���;��'���V������>מ�V4���  �  �q=u=�S=�=�=q;=��=d=3=�� =h� =b� =u� =� =>< =B��<S��<���<��<p��<���<h�<q��<�`�<0�<���<��<���<Hl�<���<6�<��<>��<9��<���<���<b��<���<{�<{��<�$�<ҝ�<���<9��<���<]�<�`�<x��<M��<0 �<���<�o�<(V�<�D�<��<���<�+�<aR�<�C�<��<���</��<���<�'�<;~�<$��<���<���<�|�<���<��<��<�f�<\��<���<�|�<o>�<�N�<U��<EW�<3�<?'�<6�<��<�u�<¼<�ĺ<V��<�!�<��<�F�<�<(��<��<�M�<0�<���<�g�<6�<`c�<��<�Θ<j�<#��<�@�<�,�<G<�<Q�<TK�<L�<��<]��<D}<u�v<k�o<�Di<o�b<�$]<�X<2�S<�P<�!M<]�J<CH<��E<=C<y&@<��<<�a8<�3<B�.<�$*<�{%<5)!<-<<�<1<�u<�~<
<(<��;���;Wo�;���;G�;�=�;k<�;̤�;��;Ϭ;G��;���;�;�;��;	�j;#sQ;,/9;�#;#�;  ;��:v��:��:��:4E�:���:T�:��:q�:� �:nVi:kD:Q�!:�:��9,��9��9�-�9��97�9%u9W�9#!8xu����Y��A��''ȹ���0I�0��;�����-��uN���w�e瓺ܙ��Ǻ�޺��x����&�X ��E��V���F��
`�=���k�p�������̠��]�� ��������q���r�JB�*�Bb�ܱ"���)��92��;�UgC��mJ���O�~S�VV��%Y���\�tPb��i��s����絆�ɬ��$b���W��^"��Q~��+T������㣻GC���R������  �  b=_e=OC=(�=Ě=�)=�=0W=k=�� =�� =N� =� =ċ =�H =`��<��<w��<I��<t|�<��<6�<X��<w<�<���<t_�<i��<<��<M�<4��<1�<�^�<���<i�<�_�<ҷ�<Cs�<ʉ�<T��<Cq�<:�<'~�<���<R��<)��<���<�;�<�l�<!��<��</��<yk�<�[�<@S�<�1�<���<�D�<�g�<�R�<��<V��<���<���<
�<P[�<��<��<S��<�[�<���<�e�<���<B�<z��<,��<�M�<�<x�<���<\+�<�
�<��<U��<M¿<�U�<���<���<2c�<a��<���<*�<��<l�<9�<lV�<ߏ�<.��<<��<��<gw�<4��<�Ҙ<Q�<0|�<r(�<�<D�<-�<�(�<��<�k�<���<�}<�lv<Q�o<��h<�b<�\<��W<XS<P�O<��L<LJ<G�G<S�E<��B<B�?<�D<<�8<6�3<ʹ.<�)<�G%<!<�,<��<�0<�<�<�F
<1X<��;���;u�;׭�;���;��;���;��;.q�;I�;�8�;0�;�;b��;j�i;�FP;��7;��!;�[;��:���:�?�:��:�:�9�:ْ�:6�:\��:�`�:�̈́:��d:)�?:B$:�:��9W��9ڑ�9�ڽ9�S�9�`�9K�9Q� 9�"8 ���/T[�����޹͹�������Ъ�Jl�H����1�YR���{�����Wׯ�g|ɺ��ມ��#� �����k�Ț�����y��k�T��[_�������w.��O� � ������a��P�����+�o��"M����F�!�\3)�d�1���:��C���J�O�P��yT��rW�JZ���]��Yc��j�|�t��~���=���@��/���	��ܟ��:�����i��S���J٢��۠�S���  �  �q=u=�S=�=�=q;=��=d=3=�� =h� =b� =u� =� =>< =B��<S��<���<��<p��<���<h�<q��<�`�<0�<���<��<���<Hl�<���<6�<��<>��<9��<���<���<b��<���<{�<{��<�$�<ҝ�<���<9��<���<]�<�`�<x��<M��<0 �<���<�o�<(V�<�D�<��<���<�+�<aR�<�C�<��<���</��<���<�'�<;~�<$��<���<���<�|�<���<��<��<�f�<]��<���<�|�<p>�<�N�<V��<GW�<3�<A'�<8�<��<�u�<	¼<�ĺ<Y��<�!�<��<�F�<�<*��<��<�M�<1�<���<�g�<6�<_c�<��<�Θ<h�<!��<�@�<�,�<D<�<Q�<QK�<J�<��<[��<D}<q�v<h�o<�Di<m�b<�$]<�X<2�S<�P<�!M<`�J<CH<��E<	=C<~&@<��<<b8<�3<H�.<�$*<�{%<:)!<1<<
�<4<�u<�~<
<(<��;���;Qo�;���;>�;�=�;a<�;���;��;Ϭ;<��;���;�;�;��;��j;sQ;/9;�#;�;���:Ғ�:j��:��:��:.E�:���:P�:��:q�:� �:lVi:iD:Q�!:�:��9+��9��9�-�9��97�9%u9W�9$!8xu����Y��A��''ȹ���0I�0��;�����-��uN���w�e瓺ܙ��Ǻ�޺��x����&�X ��E��V���F��
`�=���k�p�������̠��]�� ��������q���r�JB�*�Bb�ܱ"���)��92��;�UgC��mJ���O�~S�VV��%Y���\�tPb��i��s����絆�ɬ��$b���W��^"��Q~��+T������㣻GC���R������  �  ۛ=�=w�=�==s�=*k=��=��=�.=� =:� =ũ =-� =�[ =@ =rn�<ބ�<��<%��<���<���<�j�<�<'��<�d�<���<f�<��</��<�;�<ۖ�<z��<g�<��<��<�o�<C%�<11�<���<���<���<���<6:�<�@�<���<�z�<���<��<�<�_�<{��<�x�<B�<��<���<�y�<��<�<��<� �<9��<���<�'�< z�<P��<�2�<�^�<BF�<���<��<���<+n�<e��<�<�{�<��<���<7��<�4�<���<T��<���<Xs�<H;�<ξ<�<@$�<e�<��<a
�<���<	A�<��<��<�2�<�K�<�J�< �<�<>&�<)u�<��<�#�<���<���<'��<���<z��<H��<�g�<��<�<"�}<�kw<¿p<�+j<�c<-1^<(!Y<C�T<�Q<N<�mK<�I<�F<�C<a�@<�==<� 9<f�4<9�/<��*<V
&<��!<�a<��<��<X�<��<hu	<��<���; �;�Q�;r(�;���;8]�;L��;��;%s�;b6�;�;}Κ;z��;�i�;k�m;s�T;9�<;��&;��;�3;ʫ�:ӄ�:���:M�:���:�Ż:H�:W:�:��:�݌:Ou:�O:,:L�: Z�9���9*�9�ʮ9���9�o�9`�O9�&�8�g7�aԸ��V�Ԓ���޸��E͹�ڹ(��l��(K��#���C��m�4���W�����/uֺ@��{(��P���������D���R(����aCߺ$ܺ�Mݺ�����w�������e
�����L��WX�v��}&������$�~�+�6y3�~;�#�B��I���M�+�P��^S��V���Y���_�jJg��Sq��E}�g>��'�������`�����Z���;��'���V������>מ�V4���  �  |�=I�=M�=�{=W=��=�/=��=�M=�� =P� =� =�W =� =��<2��<�&�<DH�<:s�<��<p2�<���<���<�B�<���<Z�<���<��<g3�<3��<p �<3��<��<���<���<�B�<���<���<�&�<���<0�<i�<���<β�<�w�<\��<�C�<�k�<v��<��<�<}�<H�<F��<�o�<���<Fc�<ޡ�<���<d��<R��<�$�<�{�<���<\�<���<>��<c��<L�<<{�<kW�<���<;c�<��<�9�<"��<k��<��<� �<���<H�<��<���<j��<{C�<���<R��<bp�<X�<t��<�<���<�<�<1�<=��<j�<'פ<�<]=�<e��<�+�<g��<�/�<��<�ݑ<
�<_�<$0�<#�<j܇<bO�<�|�<n�~<�rx<��q<Ёk<yje<��_<�Z<�gV<�R<kmO<5�L<J<h�G<��D<��A<g.><�:<�5<P�0<��+<��&<w"<2�<P<#A<�.<:�<�n<ԡ<�7�;U �;b��;��;S��;)��;f�;�
�;�b�;��;x˦;~�;T<�;�C�; �q;�Y;G@B; -;�];E�
;B%�:���:��:#2�:X��:���:> �:�-�:�_�:ʧ�:���:7H_:��9:vV:*2�9���9���9~��9#��9��S9�<9�t8����� �/{W������U��+ͱ�6����gŹ�+عZd�������5�`�^�RF���]���Ե��ʺ�IܺM��\����h��Q��po��޺�غ�պ�ֺ�mۺU���w�A���-���4���
�������L�#�\�(���.�r�5�t<�:xB��?G��J�X+M�\O�8R�+ V���[�:�c���m���y��.������돻�e��ՙ����[���/����^���>��y����S���  �  }=�=��=i�=U^=��=�j=y�=�i=� =�� =XT =[ =*��<���<�Q�<˝�<���<hL�<���<Ns�<b5�<S�<2��<jd�<���<���<���<j��<�6�<���<4C�<U��<���<���<#I�<D��<���<���<�1�<Z��<���<��< �<���<u�</��<X��<7��<��<�+�<�o�<��<�Q�<���<�M�<z��<�<KG�<'��<���<4H�<���<�Y�<y��</<�<�a�<�:�<���<��<5��<��<��<���<� �<'��<���<n��<U��<~m�<)	�<���<�~�<�-�<趿<�
�<w�<I��<N��<�	�<yo�<�د<�V�<��<ϩ�<�o�<4�<H�<A��<x'�<_��<pc�<U+�<��<�4�<�c�<3��<���<���<�K�<���<E�<��<_�y<RCs<zm<?g<��a<P�\<�mX<c�T<Q<�	N<�BK<��H<q�E<'�B<�?<�;<=�6<��1<�,<8�'<5s"<.�<��<�m<�<��<� <�I<b��;-s�;�D�;���;ػ�;�T�;�0�;���;D�;�ұ;,q�;��;s�;1�;��v;�_;y�H;�b4;�M";��;K�;��:.�: ;�:�:�:.��:M˷:c�:*6�:A��:|�n:G�G:\q":zY:F��9S�9n�y9��:9-�8P5_8�v��@����&��a� N��W͐������_��w�����s[۹?�f/(��O���{��B��D˩��$�̺v�غ�w�AF�R;�:Ẻ�ۺ��պ��кOκ�)Ϻ�Ժn ݺ�`�����F~��P�g	�W��� ���$��I)�J6.���3�V9��?>�Q�B�+�E���G���I�r[K�=	N�61R�AX��\`��Rj�{�u�$񀻆��*�������nە���m������$��т��bw���a���  �  36=z4=�=:�=R�=4=��==�v=� =\v =Y =�b�<1��<D�<k}�<���<�i�<��<���<���<}�<�]�<�$�<���<�$�<�K�<:�<2��<��<G�<B��<~��<L��<�<�g�<���<���<K��<V��<I�<�?�<)h�<�k�<�:�<���<�$�<�I�<�K�<�>�<�5�<�B�<�l�<d��<]�<=p�<���<�9�<
��<��<ê�<�N�<
 �<b��<F>�<"��<���<���<��<�B�<�6�<s��<���<Y\�<`�<���<4��<��<.�<�[�<���<�[�<���<M��<��<f^�<y�<�V�<I��<3l�<���<��<�S�<���<�0�<6å<�c�<a
�<���<�e�<X'�<h�<��<{.�<�n�<���<���<��<��<��<B�<k:�<�K�<��z<D�t<@�n<�5i<��c<w"_<|�Z<�V<��R<nO<�XL<�eI<xjF<�=C<n�?<e�;<Pb7<��2<g-<�(<B�"<�Y<�9<TL<s�<b�	<|2<)� <#�;^L�;��;oT�;�+�;�R�;�}�;�X�;ȗ�;C�;f��;q1�;F0�;�͈;��z;��d;+�O;�Z<;��*;7�;�;�;&X�:q��:Dw�:o��:�w�:�E�:�'�:a��:gh�:lkz:��Q:��(:Yo:!=�9p��9D�)9,U�8n�I7#�`�r���31��B^��{��5��\c�����^Ń����줢��1ǹ���I^��3D�دl�����Js�����建��ƺ-�κ��Ӻ��պxFպȐҺ!�κY˺\~ɺ*fʺ4�κpH׺�W��P򺬌��6
������:� ��R&��u+��R0�[5���9�e�=�4A���C��E���E���F�YH��K��{O��U�?�]���g���r��}�d���p���ڍ�}���t������=���Ø��̘�.^��eė��  �  6H=�?=S%=y�=�=1=;�=�=%n=V� =>9 =^h�<���<���<��<���<��<_��<w��<J��<M��<��<p��<TN�<a��<?�<�`�<�R�<%�<-��<���<s��<ԥ�<��<��<̄�<��<��<Wp�<�X�<�^�<qt�<Z��<���<+R�<���<�L�<.s�<�k�<,F�<B�<���<���<*��<� �<�l�<<��<J�<,��<;��<R�<�+�<g�< ��<�j�<r��<��<��<�*�<�e�<�o�</Z�<�8�<W�<��<���<���<��<9�<�@�<��<���<�K�<s��<�-�<-{�<V��<i��<5)�<<��<�޲<��<E(�<[R�<���<�<�m�<��<��<�~�<�l�<���<���<��<y�<�Ր<��<+�<�<���<��<PZ�<���<W{<B�u<NPp<�k<�(f<ada<U�\<f|X<�kT<T�P<1M<��I<s�F<�tC<+�?<&
<<��7<��2<۳-<22(<4�"<�<�A<��<p�<�<�<�%�;���;W��;�.�;�Z�;l��;I��;���;���;��;-P�;��;x�;���;�ω;�~;��i;I$V;�)D;B�3;v?$;�W;�	;���:�	�:ˮ�:4��:��:DV�:�^�:�Q�:汒:�C:�cU:ۢ):�x�9�ժ9�+D9��8�ׄ��;���p�����>*��q������y���Pv�us����8~���5����������>�1b�*q�����:����B������)���ú�*Ⱥէʺ�#˺�ʺ7�Ⱥ?�ǺDɺGKͺ2պ�����ﺑ� �SW
�9��I�r�%���,�I-3���8�g=��@�X{C�bE�b�E��E�F~E��E�G���I�n�N��U�;N]��f�.�p�߽z�m��(X������=�������P���3������j�������ǖ��  �  �>=N-=u= �=�=q&=��=!�=�M=�� =���<��<���<ʥ�<6��<yr�<[!�<���<t�<�*�<�U�<s�<�n�<8�<Y��<��<�6�<V0�<v�<��<P�<N"�<�`�<p��<Q�<o��<G��<�{�<��<ȼ�<0��<�v�<�k�<�X�<L)�<s��<�3�<z^�<HQ�<s�< ��<�u�<d3�<��<�<�R�<%��<B�<l��<4��<���<&��<��<Y��<uY�<+��<���<���<�<�O�<�t�<���<���<��<U��<`��<0�<��<��<T�<��<6�<#r�<���<��<�Y�<�z�<�h�<�<'��<�Ų<�֯<�Ѭ<�˩<�ئ<}�<b`�<h�<���<`�<���<�ݖ<fJ�<̓<�M�<���<���<c�<���<e}�<�<�B�<ˎ�<��{<��v<��q<��l<r#h<^yc<��^<�BZ<��U<v�Q<9�M<J<#�F<�3C<�?<�;<c�7<C�2<M�-< �'<g"< <�<l?<��
<��<�� <���;���;�d�;���;j��;+��;���;"~�;�c�;Jo�;���;P��;1Ӟ;�k�;v�;� �;-pm;6�[;�4K;i;;3G,;��;�S;�;c��:d3�:���:,#�:��:˓�:��:��:;V|:��Q:%�#:��9X�9Yg�8N ��F#�޹����������1�ùH���\?�����Tx���!��ڒ}��#���̢�EV˹o �Jd��E>�37]��-y������(��9����䬺ݴ�(��>º�ƺ�HȺ�4ɺ�ɺn�˺ҿϺ�׺]4�;,�ƺ�)	������!�Q�+��Q4�ޡ;�QuA���E�6�H��J��(J�R9I�0�G���F��}F�E�G���J��O�ujV���^��_g��dp�n�x��U��Ĳ��A���rQ��ߋ��Z��#����ג������Ǖ�d����  �  h=� ='�=4�=wg=��=�w=�=C=ZU ='�<���<y��<��<��<�^�<v)�<�.�<�`�<��<���<�!�<�"�<S��< o�<���<���<���<���<��<�&�<���<���<�z�<=��<=l�<c��<�'�<&��<c��<���<IK�<��<���<���<rp�<���<��<�<��<1W�<��<ou�<@+�< �<�6�<���<
7�<��<{�<^=�<�h�<��<i�<��<�j�<�r�<]/�<t��<�<�K�<��<��<�3�<���<���<���<���<���<k��<���<�h�<vm�<��<�ɿ<u�<7"�<��<�Ϸ<nE�<�z�<!{�<RY�<?-�<��<O�<�O�<�ǝ<Z��<{�<���<*&�<纔<�\�<	��<�i�<)��<䴌<���<��<��<���<�k�<��{<h2w<V�r<�En<��i<XBe<ӌ`<��[<��V<�MR<��M<�I<�$F<��B<��><R;<��6<�,2<
�,<�C'<A3!<��<ڣ<<�<ۻ<�b<��;Q]�;L��;��;��;ɗ�;�1�;���;�0�;�;���;o �;�`�;Gc�;�c�;\��;c��;�5p;5U`;nQ;B;�#3;�.$;�;ǵ;Z��:I/�:.��:( �:3��:&T�:�:���:��r:q�G:SX:a��9Y6M9LlX7R�F1��v�ȹ!"�c���c�����ŒڹBt��bu��[��������p��>Z���i�W���=(��;D�Fm]�eNr�g���Q���N������t��}���Y�������uú�ɺ �̺*$Ϻ<�Ѻ�պ��ܺ�+纘����;��������&���1�p�;��.D�pkJ�S�N��P�>Q��O�:�M�3:K��iI�
�H�1J��ZM�%�R��oY��Ua�ېi��sq�)tx�CU~�y����̓�\����X������Ѝ�C���mH��El��
 ���  �  ��=3�=��=Zp=C+=��=iA=Ϛ=}� =} =Vv�<0��<L��<-��<}��<a�<�A�<Re�<��<	�<�x�<ֲ�</��<Sw�<���<�8�<�V�<�g�<P��<q��<3+�<M��<�f�<��<���<��<2q�<E��<D��<��<}w�<��<Ѷ�<3��<gG�<���<l�<0��<G��<8L�<a��<uD�<l��<�P�<��<3�<��<z@�<[2�<�Y�<���<���<y�<8��<إ�<q��<���<!��<07�<j��</�<^v�<���<���<P�<u�<'��<5��<O�<9,�<���<�z�<~J�<�D�<�_�<戽<>��<|��<ob�<\ݴ<-�<�<qѫ<���<RK�<P2�<�T�<���<�}�<���<�ߖ<�o�<�!�<Uڒ<|�<���<\:�<}:�<���<U��<5�<Q��<,�<��{<^�w<Vps<-^o<&k<�f<��a<��\<?�W<g�R<)�M<!{I<�mE<E�A<0�=<]:<4�5<P1<&,<�d&<x8 <9�<r?<��<B�<gY<���;�Q�;���;)��;sQ�;zD�;/�;@��;+c�;�)�;��;��;�J�;瀛;�;f�;���;'�q;Z�c;�U;0dG;��8;�");b};6
;j�:_a�:���:VW�:���:f�:w�:U#�:Iwd:b
::[�	:�{�9�r�8�%������ѹ����]���<����Q�e��ù��?��뛺���ع����i���5��M�KEa��jo��Ky�v���N������k ��4���-��$�����º�˺��Ѻ�1ֺ��ٺ��ݺ�G��Y�!���f��p�� %�v�+�/%8�C��L�-�R�?�V��HX��W��oU��QR��6O�s�L�\DL�ƗM�Q���V�y]��e���l��gs���x��}�	!��ɡ���\�������S��񔋻(�����������旻�  �  ʼ=��='_=�/=�=�=	=b=$� =Y��<��<!A�<���<���<���<���<B��<��<�!�<��<'�<B�<�D�<v �<w�<���<��<'��<')�<���<��<���<}��<<z�<L#�<��<p��<J�<R�<O �<�R�<��<�L�<x�<K��<�r�<8��<1�<)'�<7��<�V�<��<}�<��<�W�<qa�<���<"x�<�{�<J��<1�<g�<4��<ԏ�<X5�<���<�|�<3�<���<�7�<��<�Q�<��<���<i�<���<l1�<�1�<3��<��<���<�y�<K�<H��<f�<��<�)�<x'�<��<�o�<4��<���<�R�<��<���< x�<���<F�<���<Sŗ<.�<PҔ<薓<(^�<'�<$��<jÍ<���<�{�<��<Ǜ�<w0�<V�<_�{<+�w<0�s<�p<il<'�g<�b<��]<�LX<��R<(�M<� I<�D<�@<��<<;9<��4<�h0<�@+<�%<`G<�<�
<)�<S<|h�;,��;A�;'��;c
�;���;�#�;W@�;���;*��;�:�;��;ˬ;u9�;��;5p�;��;�V�;��r;��e;��X;V&K;�j<;��,;,;��;{s�:���:��:t��:T��:0Ǘ:��:��x:n�U:2�+:�F�9��9�^8n� �t�����h�.$1�P7��)2��%��)��Q �p���͹��ɹ��ع���.�:+��PC���W�of���n�V]s���v�{|�N���NR�����%;���)��86ú�κ�u׺Hݺ�������.�P������w1��{�Q/#�x0��]=�>�H�ylR�b9Y��3]��f^�,3]��LZ���V�S��P���O�6<Q���T�z�Z�υa���h�l�o�Ջu��y�\r|�|Z~�!"��������Rp��%�����O*���ᕻh蘻�  �  ��=�]=N/=)�=I�=S`=b�=�7=(r =1�<�s�<3��<WZ�<$7�<�q�<��<�<�I�<��<�;�<Q��<���<���<[��<i�<�U�<fx�<��<���<�_�<��<���<���<���<�l�<���<O(�<q6�<�)�<N�<�4�<�}�<m��<@��<�d�<��<��<\��<r��<��<���<�U�<S��<�#�<���<���<�9�<���<��<KJ�<O��<�<�E�<[<�<l��<�(�<��<C��<�c�<���<��<<3�<��<��<2��<�1�<G��<��<4�<m��<|�<�r�<r��<���<��<⳼<�˺<H˸<��<��<�Q�<E@�<��<���<�5�<���<��<te�<Z%�<�D�<��<vf�<L5�<"�<״�<o0�<Gi�<^�<��<���<�A�<_�<�d<d{<0�w<�-t<;�p<�l<�Ih<oc<(&^<d�X<%S<#�M<��H<�$D<#@<�7<<�^8<bF4<��/</�*<��$<��<��<86<!�
<�Q<5G�;4X�;/��;H��;�4�;�@�;k��;���;�s�;�$�;�ż;Zc�;�;�;��;C�;]X�;@A�;R�;�Ds;�g;�Z;&`M;��>;7�.;m�;N�;�E�:,��:�C�:D��:�:���:�ׄ:�&m:�J:$!:���9��h9H�6��W�n�й��go0��5B��iG��fA��2�H��z��,��~@��߹���^9�XH���6�VM�8G_�	�j�J�o��Sp�9�p��-t�J�}������,���|�����S�ú{^Ѻ�ۺ?��lk���뺧�}�����b��}.�V&��3���@���L�o�V�e�]��ka�hb���`���]�-�Y���U��+S��pR�<T���W�5�]���d�P�k��r��)w��tz�8F|�ZR}��~�Cf���`��ER���!������L��Z4�������  �  ��=ӯ=m=�%=��=�f=��=_H=� =ͼ�<�E�<K��<���<��<���<�}�<I�<�J�<�r�<���<���<���<���<ߞ�<[*�<I��<@��<�&�<�|�<��<_v�<��<x��<�x�<-�<B��<���<a�<=%�<N�<:��<<��<�[�<���<>m�<:��<QB�<yn�<wg�<�0�<���<�h�<���<��<܎�<��<���<��<Ka�<�Y�<�i�<Dx�<�n�<�7�<���<:�<��<*��<ӭ�<(O�<t��<ҋ�<�1�<��<Sm�<���<�(�<9�<��<���<.u�<e�< ��<���<-��<㏼<j��<�]�<��<풳<%ް<���<��<�ۧ<|Τ<�<�"�<���<df�<�m�<#��<�#�<���<2G�<E̐<)0�<h�<bq�<�Q�<��<�̈́<k��<�W�<L{|<urx<�t<y�p<�kl<nh<RQc<�[^<�@Y<^(T<W7O<ƂJ<mF<��A<��=<�u9<�5<�Q0<m.+<ԣ%<��<�<u�<K<��<"|<ie�;i��;+q�;���;���;�d�;���;���;If�;8�;Z�;d�;":�;�|�;���;��;�^�;�~;5q;ɬc;�U;�zG;wc8;��(;�;�&;���:���:2m�:O��:�B�:�$�:�:F}t:YVJ:�:Ԥ�9��c9F8�e	�����@�Ź����������G���6�ۖҹ:��r���삹���ǹ'��U�m��$^)��:��*I��T�UZ\�8�c��&m��y�(Ʌ�nߐ�I����ܪ�!���d�ºXY̺KmԺ��ۺ>�<-����������S��-!���,�9�7�؆A���I�3P��iT���V�*�V�x�U�T��UR�n=Q��[Q��S��<V�d�Z�nZ`��<f��k�H�p��*u���x�H\{�@.~��ɀ�3���hƅ�T������|[��j������  �  ��=ط={v=�/=��=�p=1�=S=S� =���<#`�<� �<���<b��<}�<��<�g�<g�<���<C��<,��<�
�<���<w��<?�<^��<���<6�<���<F��<uu�<{�<��<�f�<��<�k�<��<���<�<MJ�<ӎ�<���<�h�<���<���<���<�V�<#��<m|�<;F�<k��<`��<��<T��<Y��<���<��<���<�~�<)u�<J��<"��<&��<�L�<��<z&�<�3�<?�<���<L\�<���<[��<�-�<���<>]�<b��<]�<�"�<'�<��<l�<��<���<���<��<%��<���<�q�<�%�<��<��<|�<��<���<�<��<�B�<nÜ<��<���<NΖ<�>�<6˓<,^�<)�<xE�<}�<t��<lf�<)�<Eބ<Ζ�<J_�<�}|<�gx<�lt<�kp<�Bl<r�g<m'c<&8^<�'Y<cT<T7O<ӎJ<�&F<��A<��=<��9<u65< z0<�W+<n�%<��<6�<]�<>�<1<�<���;�i�;���;>T�;b�;���;�*�;N<�;���;���;��;�D�;���;���;�*�;?�;�]�;Tb~;y�p; c;�CU;`�F;��7;�v(;�Y;g;�"�:�7�:H�:㴿:��:s�:�i�:�w:��L:�:�k�9aBp9ƇF8�7��@Ņ�8���Ȱ�i���ّ���l���|�̹ޠ��P[��kT��c�¹(�ܹQ���ص���'�c�9���H�GuT��]���e���o�G�|�������_v��$_��$���i�ºR�˺��Ӻ}�ںT�ẓ���8��\O�u��C�u[ ��+�1�6�]�@���H��,O�eS�a�U���U��U�2VS���Q�X�P�]�P��\R�$�U�2Z���_�/�e���k���p�!u���x�5�{�`�~�����R�����fZ��L医fs��S���ħ���  �  �=��=�=�K=��=�=\=�p=�� =� =���<�S�<?%�<<-�<�s�<��<���<d��<���<`�<22�<�E�<�1�<b��<px�<O��<q!�<�_�<���<���<�p�<���<��<�/�<s��<�+�<��<���<i��<:=�<^��<D�<D��<�"�<���<P5�<���<,��<��<���<�,�<���<�h�<u#�<V	�<
%�<|�<�<|��<���<6��<���<.��<b��<%�<_�<Vk�<<@�<k��<(��<�	�<���<p �<���<e,�<���<���<���<q��<?��<�O�<>�<���<���<�̾<�ϼ<�ɺ<���<�]�<q߳< ,�<�J�<�I�<�<�<�9�<�T�<鞟<j"�<a�<\�<�"�<ߋ�<[�<���<�<�<:��</��<e��<�]�<��<��<�r�<%�|<�Dx<%t<p<��k<�Vg<`�b<=�]<��X<]�S<3O<R�J<)dF<�DB<�2><�
:<��5<��0<]�+<�D&<�l <�b<fP<�`<"�<�|<n�;���;�V�;s��;���;��;�,�;�2�;���;�~�;���;>)�;@V�;�j�;}��;�@�;R�;|�};�ro; xa;W\S;��D;B�5;�';�h;��
;A��:v��:o��:��:0�:��:u�:�v~:�dT:n_&:o��9��9���8D���/�]�6	��(�˹��แ
�2�޹�Ϲ|���i�������ʥ��P��%�ι�]������"���6�k�G���U��@a�	�k���v�sU�����D��� $��'�����&���S�ɺT�к%�׺^�޺�N�ښ��} ��@	�$W��G��t)�`04���=���E�A4L��sP���R��ZS�i�R��,Q���O�ǲN�X�N�y�P���S�rX��"^��Rd�{j��'p�Uu�I?y���|�d%��X��BT��U�� +��%{��~������b���  �  "=��=˳=0r='=^�=%3=Y�=�� =�> =�< ��<���<A��<��<݋�<H�<h4�<E�<Bh�<c��<��<7��<A<�<��<�&�<�f�<��<}��<H�<nb�<y��<�O�<���<�R�<���<:�<�q�<���<G"�<��<� �<��<�b�<���<-��<��<��<>�<���<	��<s0�<���<���<�<��<E�<)��<�X�<S:�<_2�<�,�<��<���<V`�<��<7��<E��<d+�<��<�$�<���<��<�s�<��<-�<�a�<t�<g�<E�<��<o��<���<���<���<^�<��<��<z��<�+�<�z�<���<J��<��<沥<Iۢ<�.�<E��<0x�<�s�<D��< �<�x�<c��<gt�<�ҏ<��<��<N�<^��<bJ�<��<���<hx|<x<<�s<Zo<��j<Zf<��a<\]<�TX<�S<�O<T�J<W�F<�B<F�><�:<�A6<��1<�h,<��&<� !<�,<%5<�a<L�	</�<7��;�5�;��;	��;%\�;5t�;8��;��;���;/��;Y�;Eh�;qy�;�Y�;6K�;!��;�$�;�o|;sYm;�^;35P;<�A;03;?�$;ݾ;��	;?��:^��:n��:���:f��:{�:��:�<�:r�^:1:F�:�;�9^9��]����� ����������Ĺ���������㤹3���)|��v������b��b�߹������2��<G���X��g��Su�jn���ٕ��V�����⯺�+��>$����Ǻa�ͺ�?Ӻ�ٺmg����	��д�y��uB��&�-\0���9��sA���G���K�adN��UO�	O���M�B�L��L��bL��N��SQ�V��[�1gb�'i�-vo��:u��Jz���~�Yx��;�������ݤ��҆���|���T���ᓻ����  �  �5=R	=��=ژ=tF=��=�[=��="=�x =`��<�n�<*]�<�w�<���<XB�<���<���<���<g��<���<'��<V��<��<��<'s�<���<���<���<
�<D�<���<��<�V�<���<�0�<���<�<�q�<���<ϊ�<5�<���<3��<�I�</��<!.�<[�<�Y�<�1�<|��<��<�l�<�H�<H�<2r�<���<�N�<	��<���<1��<���<�n�<�&�<}��<��<��<���<�i�<���<q8�<���<���<m �<�g�<���<���<G��<���<��<e��<m��<���<��<0�<P�<nY�<>�<��<�w�<�˱<���<��<R&�<_F�<��<Q�<r�<�1�<o#�<�C�<_��<��<�a�<�Α<&�<Z�<cb�<�=�<��<숅<A�<\��<�S|<�w<O�r<Rkn<��i<�Xe<�`<$\<�W<5(S<;�N<c�J<��F<�(C<�G?<�6;<�6<="2<*-<ߖ'<��!<<
F<�<q3<�<�c<��;?�;4�;�z�;HE�;0�;���;�P�;�;n4�;㬳;*��;�H�;T��;��;;#zz; Xj;��Z;�K;27=;m�.;�,!;|G;"�;�M�:��:���:��:�d�:n�:w �:HJ�:Si:��<:�:���9e�[9}�8��v�4�$��.p��5��޲��Ƙ��P���A�������pu��d|��錹������̹����wo���/�$'H�|^�8�q�����������������r]���!���J��kQ���!����ź�9ʺ��κպ%�ݺ��躎��t�M������"�b�+��_4��;�G�A��F�I�H�-eJ���J��RJ��I�AUI���I�P�K���N��S���Y��~`���g�>o�M�u���{�)ƀ��Q���ǅ��C��ӊ�k������A>��2<��Fꕻ�  �  �?=�=��=!�=.c=��=�z=�=�N=�� =0 =X�<��<�E�<A��<��<۫�<�m�<�M�<�B�<?�<�2�<j�<���<�N�<$��<���<u��<7��<���<��<2�<gk�<Ÿ�<��<	~�<@��<r�<��<B��<cj�<Z7�<��<���<��<9
�<�g�<2��<^��<�~�<R�<�#�<��<��<��<�B�<՚�<��<���<ya�<�(�<���<ǻ�<{f�<���<�.�<S8�<��<
��<���<�8�<�f�<w��<���<���<��<��<*(�<�9�<�L�<�i�<A��<���</�<�L�<x{�<���<Xr�<�(�<���<��<�I�<>x�<���<�<78�<���<=D�<l�<'�<k�<��<f�<��<a�<�g�<3��<b��<y�<�(�<���<�)�<9��< |<{�v<�	r<h>m<c�h<�c<�a_<z�Z<k�V<bzR<4�N<��J<}G<[sC<}�?<��;<\I7<�2<`�-<Z&(<��"<H�<�`<)�<"�<�<4<�`�;�;�;b��;���;�
�;ޜ�;"�;�\�;p�;o0�;F��;��;f�;�-�;�s�;���;1�w;@uf;�V;��F;n�7;�);m�;��;�x;Q�:[_�:���:��:��:Ľ�:�ڟ:��:�`q:�eF:=�:���9i�9G�9B38zp�|5���<�v^�6�l�=�l�xFc�N~X�bT�P�^��}��8��K��4���!H/��K��df�k�~�;��e��y��T����d��h��FM��.뾺9eºz.ź�Ⱥ9�˺�Ѻ��ٺ6%��C���������*��(�&���.��w5�n";�U�?���B��E�$CF��F���F�\G�V�G��I��M���Q�!�W�,_��g�w.o�bw�Mw~�����妅�`s�����L���"̏��ԑ�싓��	���  �  �:=�!=k�=|�=�m=a=��=- =Vp=A� ={Y =��<U��<��<�m�<���<�e�<4
�<r��<=��<8|�<�Z�<*�<��<d�<y��<���<b��<t��<���<���<I��<C��<{�<�M�<Բ�<�1�<���<j�<~M�</0�<��<��<���<̒�<,�<�|�<���<ڻ�<���<��<ʎ�<v��<T��<��<2�<p�<���<n]�<���<Y��<YD�<	��<,��<���<�@�<�I�<�<���<���<��<�*�<�+�<�)�<�*�<r2�<A�<�W�<Uy�<ʨ�<h��<;:�<F��<��<�I�<{��<ڙ�<<�9�<�Ŵ<�-�<i��<�ʬ<��<�y�<��<�x�<�<�ԝ<���<��<���<�̕<��<�L�<ω�<`��<O��<W��<�<�<d��<�#�<it�<�{< &v<��p<��k<�g<�Qb<��]<ƅY<�rU<A�Q<�M<�vJ<�G<�|C<��?<;�;<�n7<��2<�-<@}(<h#<ʹ<�h<�;<�;<Jj	<��<#X <�:�;�9�;���;ӊ�;ݫ�;#��;���;8��;
��;�
�;�ի;��;_�;�ڍ;CЃ;>t;a�a;��P;�l@;�1;�#;6�;��;��;��:q��:���:2��:�O�:�7�:ZV�:(Î:[�u:��L:��$:ؼ�9��9�s9��96B;8�5��B���t���#���4���;���=�}�B���Q�H<r���lp��գ�׵��22�zR���q�Ko��z{��0柺����j����6�������ĺXRź�Fƺ��Ǻ%�ʺ^к��غ�㺋��`� �3?	�m���:�'�!�V�(��/��j4��9���<���?� B���C���D�
�E���F��I�oiL�w-Q�idW���^��Kg��4p�('y�$܀��τ��]��)����>�����������X=�����~����  �  Q%="=�=�=pc=��=�=�=A�=n=�� =�& =p��<[��<+9�<6��<��<~��<w.�<J��<Y��<a�<��<���<:O�<>��<C��<���<��<*��<Z�<5�<�)�<�>�<z�<��<je�<*�<7��<��<���<���<]��<N��<�|�<
�<�h�<���<���<h��<���<���<=
�<�C�<���<%��<�9�<{��<���<�o�<Q��<w�<��<u��<D��<"*�<�0�<M��<�~�<���<���<���<B��<���<�q�<2a�<�c�<�{�<1��<���<7V�<���<�E�<���<p"�<Df�<�~�<ng�<�!�<#��<O-�<_��<z�<�y�<���<��<�8�<C�<���<�^�<�0�<��<��<�4�<�\�<���<棎<���<�}�<�(�<"��<	��<�6�<�z<E,u<ïo<#gj<_e<��`<�)\<�X<'(T<��P<1M<��I<(�F<8;C<�?<-�;<�@7<�2<��-<��(<j#<�K<�H<g<ץ<��
<i<��<��;��;[`�;u��;	C�;��;���;{X�;�a�;=ʹ;�;찡;�^�;nь;L�;!"p;v�\;��J;��9;�*;Ƕ;�0;�\;E ;��:���:h��:Z��:}!�:��:�=�:���:��u:"�O:��*:�&	:Q�9�d�9�=f9��9���8���6͚P��ȸ]�v9!���2���B�l�X���{��3��oտ����c1��9��\����V�����������%��bg��Pź��Ⱥ�ʺ��ʺ��ɺnaɺ�ɺ�s̺�Ѻ�ٺ����P�� ��_�l��+�h��{�#��	)�N.���2�,/7�>!;��z>�9.A��QC��'E�2G���I�M���Q�RX���_��h�)r�� |�ς�:I��eK���������ޓ�ꇕ�k����?��烗�*����  �  z=�=��=-�=9G=
�=
r=%�=��=�=z� =d =� =���< ��<MI�<���<��<�{�<��<���<�H�<���<���<^�<�p�<���<>��<?q�</�<���<5��<�}�<4}�<Q��<�	�<��<�^�<�J�<)W�<�t�<���<���<���<9C�<���<e1�<o�<���<Q��<���<@�<=l�<���<.�<z��<���<�;�<���<_��<-�<���< ��<�b�<J��<)��<>��<غ�<k>�<���<P��<�i�<0�<;��<M��<��<��<���<���<N@�<���<�J�<���<k�<�۾<�%�<�?�<9)�<�<�<F�<k��<�"�<���<�k�<&$�<�ߣ<ʘ�<�K�<"��<M��<�u�<SQ�<�E�<�O�<�c�<�s�<
o�<�F�<���<j�<��<��<b�y<2t<)hn<~�h<C�c<$�^<щZ<2�V<��R<�uO<�JL<�4I<�F<��B<�?<�;<L�6<I,2<�W-<sj(<*#<N�<��<2a< �<d_<��<|E<=f�;&c�;Ĭ�;Y�;7i�;���;�A�;���;U��;[��;R��;�Ơ;�F�;�o�;>��;��k;$wW;أD;�3;ۉ$;`�;��;�;�N�:���:���:+��:��:���:d��:O�:��:��q:
sN:��-:��:���9>"�9ӳ�9ˀl9�b"9��8�7+�B���ϸ��2"6��R��pp���������7ιy �*���C�N.i�����JK���ު����Bĺ�o̺�ѺG�Ӻ��Ӻ�8ҺW�Ϻ)κ��ͺs#кtJպhwݺ�N����s�a�o�����A�%���#��y(��T-�K2�+7�O�;���?���B��E�iEH��'K�R�N�-�S���Y���a�	�j���t��f��섻�Չ�8��{�~攻0���}���9���i��	B������  �  .�=��=��=�p=� =[�=�T=i�=
�=,)=�� =q� =�P =o =�}�<���<��<8`�<��<��<��<��<���<�J�<���<"�<�M�<�H�<��<��<En�<p�<���<���<���<N�<9��<���<ٶ�<���<C�<:4�<�H�<E6�<s��<&��<|��<+�<c�<���<*��<wC�<���<&2�<G��<��<}z�<ܾ�<���<� �<VT�<���<���<x.�<yu�<I��< ��<�h�<8��<5)�<�)�<o��<ڭ�<+X�<��<���<���<e��<�*�<F��<�(�<}��<�s�<�<ф�<Ѽ<d�<�ָ<혶<w@�<4ݱ< ~�<�,�<��<׽�<蔦<�f�<�)�<�ٟ<�y�<��<ʷ�<�o�<yB�<I/�<�-�<�/�<$�<+��<<��<�b�<�<�y<Ms<�5m<&�g<sRb<Oy]<�Y<�$U<��Q<�cN<�`K<4kH<�[E<�B<�t><G|:<#-6<��1<��,<f(<6m#<p�<�q<C"<��<~<�	<x`<�L�;���;_��;߱�;?@�;�1�;R_�;��;3r�;�ղ;���;_��;k��;N�;�~};��g;��R;�E?;��-;��;;)�;d�:��:wH�:��:��:'�:Y�:eި:1K�:��:�]k:PK:%.:�j:>� :%�9�:�9/<�9��j9k}9k �8�}%��;��Z;�;�B� �k�j؈�����������Ag
���)�ЊN��xv�豏�Pf��w1���=ĺB�Ϻ�غٝܺQ�ݺ��ܺ��ٺ�^ֺ[�Ӻ�Ӻ�պT5ں�V���캤��A��J������b������������#���(��c.��4�Ȩ9�V�>�C���F��	J��ZM��4Q��V�g]\��-d�ptm���w�t��7���{8���␻f̔��֗����.��Ĥ��T����
�������  �  Ӭ=�=%�=�I=2�=ۛ=L7=��=	{=�-=�� =X� =�| =�> =���<m6�<In�<C��<���<��<]w�<'��<�x�<��<{�<\��<���<���<���<~n�<��<���<b]�<bA�<�]�< ��<mW�<1�<=�<�k�<8��<N��<B��<3��<���<�3�<���<`��<X-�<a{�<���<fV�<y��<�{�<��<���<g��<��<�>�<=S�<�i�<���<+��<5��<P1�<iU�<�R�<`�<h��<&��<#��<ܗ�<"?�<���<݂�<&F�<�1�<�L�<��<�<��<>`�<��<\��<�0�<�~�<���<���<6L�<���<���<Za�<�*�<8�<��<7�<�Ȥ<ړ�<)A�<�ԝ<�Z�<��<�}�<"5�< 
�<;��<��<�ً<#��<zV�<�̈́<T�<�S~<IMx<�6r<\;l<��f<�-a<ON\<��W<UT<��P<~M<}�J<��G<#�D<�nA<F�=<i�9<n�5<4
1<�h,<��'<0I#<+�<��<��<i�<O<�	<�.<�T <W��;�"�;���;���;���;�v�;�x�;�K�;���;{a�;/`�;Բ�;���;cz;�d;�N;k�:;�i);@;�;�b;Ѩ�:���:�o�:���:���:�V�:%�:��:���:�ł:��d:��F:l-:S�:�: �9f��9d��9���9b]J9 ��8�t7�䐸�>�7�R�9Ȃ�{p��<��Ȝι;����D�x4�hMY��)��$^���ꪺ�����-ͺ�4ٺ�F�yq庋��些Aມ(ܺ�ٺغ�ں�!ߺ3���b��]�C�	�����~������v��� �ï%���+���1��Z8�?L>���C���G�d�K���O���S���X�]�^�v�f��p�
�z�*���)����+�������C'���:���W��M���KE�����8��  �  �=�='f=�,=s�=q�=�!= �=�r=�.=0� =�� =)� =c] = =�r�<]��<��<��<Y�<Uc�<���<?K�<���<�B�<���<���<Z��<���<�.�<&��<�X�<?	�<��<���<[�<���<���<���<�"�<
f�<��<]��< ��<�k�<���<�c�<���<��<�`�<a��<7^�<��<���<#E�<��<�"�<W�<�k�<{o�<s�<^��<@��<���<T �<Y�<-�<���<r]�<d��<���<�S�<���<��<�)�<h��<���<Z��<(;�<M��<�^�<4�<���<�t�<��<tB�<�]�<�J�<e�<�ͳ<(��<�I�<�$�<*�<9�<*�<��<�Ӣ<��<@�<a��<b��<���<�'�<R�<N͏<Ϻ�<���<�t�<m�<��<�ց<$�}<��w<�q<~�k<��e<�q`<T�[<V1W<�WS<7�O<-�L<c	J<:3G<8D<p�@<�\=</f9<�5<�0<�,<b�'<�(#<�<��<9�<|�<��<C`
<_�<z� <�i�;cn�;���;p��;��;#��;��;�t�;̰;I��;�;7˒;���;Fx;�a;�L;�68;��&;BV;E�
;� ;���:���:
f�:M�:��:)ȼ:���:"��:�U�:T�:��_:j�C:��+:a�:(
: !�9?��9�b�9E��9F6g9�#9��7׆��y��_�Ta���g��̭��b�ܹ����v`;�8�`��B��ܚ��ޯ���º�Һ�"ߺ�/纀��j�a�躈��.ຏ�ܺE�ۺ��ݺ����S���~���{�wy
�$�������(~�������#���)�Y�0�ϥ7�h.>���C���H�>%M��Q��QU�WZ��`��zh���q��|����-≻Xr���h��]�����������ໞ�$螻�q������'휻�  �  k�=s|=�[=h"=P�=y=�=P�=�o=�.=[� =�� =� =�g =� =׆�<��<
��<���<��<�[�<N��<�:�<u��<{.�<��<��<l��<,s�<�<˩�<;>�<,��<���<	��<S:�<��<��<>��<�	�<�N�<��<<��<5��<W�<���<�O�<���<��<�V�<��<,`�<��<ص�<�W�<]��<<8�<%j�<�z�<{x�<�u�<�<���<x��<Z��<9
�<�<���<H�<���<cz�<�;�<���<}m�<�<���<1��<���<��<���<�B�<���<.��<�]�<�ݽ<�,�<|H�<�5�<O�<��<�w�<RA�<�!�<��<f�<�$�<��<��<���<`�<���<��<���<�"�<��<E��<���<�<[`�<'	�<r�<���<߫}<`�w<]nq<�^k<T�e<1`<L[<��V<}S<8�O<��L<��I<rG<�D<��@<�2=<<9<p�4<}0<��+<rt'<#<��<��<�<R<�<ό
<�<� <���;���;���;��;���;9��;�h�;&�;y|�;�2�;W.�;�w�;�;�;|�w;Z�`;d3K;�A7;��%;�T;��	;f��:(�:���:���:��:\��:���:.N�:cL�:�:�Z}:�!^:ckB:Y+:�2:+*: ��9���9ǿ�9��9��p9X�9r+	8���-I���c��㏹�ͩ�ܙù��ṙ��� ��>���c�v���1m��������ĺ��Ժm/Ắ:���@�m��0�����,޺�
ݺ1�޺��L�o��|� ����c�
�!��
����(��������#�S)�YJ0�6m7�*>�o#D�k;I���M�ܯQ���U���Z��Ha��!i�/�r�/F}��j���I��{㏻�┻C���&��3��7��\Z��ڞ�S
���F���  �  �=�='f=�,=s�=q�=�!= �=�r=�.=0� =�� =)� =c] = =�r�<]��<��<��<Y�<Uc�<���<?K�<���<�B�<���<���<Z��<���<�.�<&��<�X�<?	�<��<���<[�<���<���<���<�"�<
f�<��<]��< ��<�k�<���<�c�<���<��<�`�<a��<7^�<��<���<#E�<��<�"�<W�<�k�<{o�<s�<^��<@��<���<T �<Y�<-�<���<r]�<d��<���<�S�<���<��<�)�<h��<���<[��<);�<O��<�^�<6�<���<�t�<��<vB�<�]�<�J�<g�<�ͳ<*��<�I�<�$�<+�<:�<+�<��<�Ӣ<��<@�<`��<a��<���<�'�<Q�<L͏<ͺ�<���<�t�<k�<��<�ց<!�}<��w<�q<|�k<��e<�q`<T�[<W1W<�WS<8�O</�L<f	J<=3G<�8D<s�@<�\=<3f9<�5<�0<�,<f�'<�(#<�<��<;�<}�<��<C`
<_�<y� <�i�;^n�;|��;i��;��;��;��;�t�;̰;@��;�;/˒;���;�Ex;ݫa;�L;�68;��&;:V;?�
;� ;���:��:f�:I�:��:'ȼ:���: ��:�U�:S�:��_:j�C:��+:a�:'
: !�9?��9�b�9E��9F6g9�#9��7׆��y��_�Ta���g��̭��a�ܹ����v`;�8�`��B��ܚ��ޯ���º�Һ�"ߺ�/纀��j�a�躈��.ຏ�ܺE�ۺ��ݺ����S���~���{�wy
�$�������(~�������#���)�Y�0�ϥ7�h.>���C���H�>%M��Q��QU�WZ��`��zh���q��|����-≻Xr���h��]�����������ໞ�$螻�q������'휻�  �  Ӭ=�=%�=�I=2�=ۛ=L7=��=	{=�-=�� =X� =�| =�> =���<m6�<In�<C��<���<��<]w�<'��<�x�<��<{�<\��<���<���<���<~n�<��<���<b]�<bA�<�]�< ��<mW�<1�<=�<�k�<8��<N��<B��<3��<���<�3�<���<`��<X-�<a{�<���<fV�<y��<�{�<��<���<g��<��<�>�<=S�<�i�<���<+��<5��<Q1�<iU�<�R�<`�<h��<'��<$��<ݗ�<"?�<���<ނ�<(F�<�1�<�L�<��<�<��<A`�<��<`��<�0�<�~�<��<���<:L�<���<���<^a�<�*�<:�<���<8�<�Ȥ<ړ�<(A�<�ԝ<�Z�<��<�}�<5�<
�<8��<��<�ً<��<vV�<�̈́<Q�<�S~<CMx<�6r<Y;l<��f<�-a<ON\<��W<WT<��P<~M<��J<��G<*�D<�nA<M�=<q�9<v�5<<
1<�h,<��'<6I#<1�<��<��<l�<O<�	<�.<�T <P��;�"�;���;���;���;�v�;�x�;tK�;���;ja�;`�;Ų�;���;�bz;�d;�N;X�:;�i);@;��;�b;¨�:{��:�o�:���:���:�V�:"�:��:�:�ł:��d:��F:k-:R�:�: �9e��9d��9���9b]J9 ��8�t7�䐸�>�7�R�9Ȃ�{p��<��Ȝι;����D�x4�hMY��)��$^���ꪺ�����-ͺ�4ٺ�F�yq庋��些Aມ(ܺ�ٺغ�ں�!ߺ3���b��]�C�	�����~������v��� �ï%���+���1��Z8�?L>���C���G�d�K���O���S���X�]�^�v�f��p�
�z�*���)����+�������C'���:���W��M���KE�����8��  �  .�=��=��=�p=� =[�=�T=i�=
�=,)=�� =q� =�P =o =�}�<���<��<8`�<��<��<��<��<���<�J�<���<"�<�M�<�H�<��<��<En�<p�<���<���<���<N�<9��<���<ٶ�<���<C�<:4�<�H�<E6�<s��<&��<|��<+�<c�<���<*��<wC�<���<&2�<G��<��<}z�<ܾ�<���<� �<VT�<���<���<x.�<yu�<I��< ��<�h�<8��<5)�<�)�<p��<ۭ�<,X�<��<���<���<h��<�*�<J��<�(�<���<�s�<�<ׄ�<�Ѽ<j�<�ָ<�<|@�<9ݱ<%~�<�,�<��<ٽ�<ꔦ<�f�<�)�<�ٟ<�y�<��<ȷ�<�o�<uB�<D/�<�-�<�/�<z$�<%��<飇<��<�b�<�<�y<Fs<�5m<#�g<qRb<Oy]<�Y<�$U<��Q<�cN<�`K<=kH<\E<�B<�t><R|:<.-6<��1<��,<o(<?m#<x�<�q<H"<��<~<�	<w`<�L�;���;S��;б�;.@�;�1�;<_�;i��;r�;�ղ;}��;H��;U��;9�;�~};q�g;m�R;gE?;��-;�;�;�;M�:��:iH�:��:��:'�:U�:aި:.K�:��:�]k:NK:%.:�j:>� :$�9�:�9/<�9��j9l}9l �8�}%��;��Z;�:�B� �k�j؈�����������Ag
���)�ЊN��xv�豏�Pf��w1���=ĺB�Ϻ�غٝܺQ�ݺ��ܺ��ٺ�^ֺ[�Ӻ�Ӻ�պT5ں�V���캤��A��J������b������������#���(��c.��4�Ȩ9�V�>�C���F��	J��ZM��4Q��V�g]\��-d�ptm���w�t��7���{8���␻f̔��֗����.��Ĥ��T����
�������  �  z=�=��=-�=9G=
�=
r=%�=��=�=z� =d =� =���< ��<MI�<���<��<�{�<��<���<�H�<���<���<^�<�p�<���<>��<?q�</�<���<5��<�}�<4}�<Q��<�	�<��<�^�<�J�<)W�<�t�<���<���<���<9C�<���<e1�<o�<���<Q��<���<@�<=l�<���<.�<z��<���<�;�<���<_��<-�<���< ��<�b�<J��<)��<>��<ٺ�<l>�<���<Q��<�i�<0�<=��<O��<���<��<���<���<R@�<���<�J�<���<k�<ܾ<�%�<�?�<@)�<�<���<M�<p��<�"�<���<�k�<)$�<�ߣ<ʘ�<�K�< ��<J��<�u�<NQ�<�E�<�O�<�c�<�s�<o�<�F�<���<yj�<��<��<X�y<*t<#hn<z�h<@�c<$�^<ӉZ<6�V<��R<�uO<KL<�4I<F<��B<�?<
;<Z�6<W,2<�W-<j(<5#<W�<��<8a<�<f_<��<zE<5f�;c�;���;Y�;!i�;o��;�A�;l��;9��;>��;5��;�Ơ;�F�;�o�;'��;z�k;�vW;��D;��3;$;K�;��;�;�N�:���:���:!��:��:�:`��:M�:��:��q:sN:��-:��:���9>"�9ӳ�9ˀl9�b"9��8�7)�B���ϸ��2"6��R��pp���������7ιy �*���C�N.i�����JK���ު����Bĺ�o̺�ѺG�Ӻ��Ӻ�8ҺW�Ϻ)κ��ͺs#кtJպhwݺ�N����s�a�o�����A�%���#��y(��T-�K2�+7�O�;���?���B��E�iEH��'K�R�N�-�S���Y���a�	�j���t��f��섻�Չ�8��{�~攻0���}���9���i��	B������  �  Q%="=�=�=pc=��=�=�=A�=n=�� =�& =p��<[��<+9�<6��<��<~��<w.�<J��<Y��<a�<��<���<:O�<>��<C��<���<��<*��<Z�<5�<�)�<�>�<z�<��<je�<*�<7��<��<���<���<]��<N��<�|�<
�<�h�<���<���<h��<���<���<=
�<�C�<���<%��<�9�<{��<���<�o�<Q��<w�<��<u��<D��<#*�<�0�<N��<�~�<���<���<���<D��<���<�q�<5a�<�c�<�{�<6��<���<=V�<���<�E�<½�<x"�<Lf�<�~�<vg�<�!�<*��<V-�<e��<�<�y�<���< ��<�8�<C�<���<�^�<�0�<��<��<�4�<�\�<�<ޣ�<���<�}�<�(�<��<��<�6�<�z<<,u<��o<gj<_e<��`<�)\<�X<-(T<��P<1M<��I<5�F<F;C<��?<=�;<�@7<�2<��-<��(< j#<�K<�H<g<ۥ<��
<i<��<��;��;J`�;`��;�B�;��;���;\X�;�a�;ʹ;ԍ�;Ͱ�;~^�;Qь;�K�;�!p;L�\;x�J;w�9;��*;��;�0;�\;9 ;��:���:]��:Q��:v!�:��:�=�:���:��u:�O:��*:�&	:P�9�d�9�=f9��9���8���6˚P��ȸ]�u9!���2���B�l�X���{��3��oտ����c1��9��\����V�����������%��bg��Pź��Ⱥ�ʺ��ʺ��ɺnaɺ�ɺ�s̺�Ѻ�ٺ����P�� ��_�l��+�h��{�#��	)�N.���2�,/7�>!;��z>�9.A��QC��'E�2G���I�M���Q�RX���_��h�)r�� |�ς�:I��eK���������ޓ�ꇕ�k����?��烗�*����  �  �:=�!=k�=|�=�m=a=��=- =Vp=A� ={Y =��<U��<��<�m�<���<�e�<4
�<r��<=��<8|�<�Z�<*�<��<d�<y��<���<b��<t��<���<���<I��<C��<{�<�M�<Բ�<�1�<���<j�<~M�</0�<��<��<���<̒�<,�<�|�<���<ڻ�<���<��<ʎ�<v��<T��<��<2�<p�<���<n]�<���<Y��<YD�<	��<,��<���<�@�<�I�<�<���<���<��<�*�<�+�<�)�<�*�<u2�<A�<�W�<Zy�<Ϩ�<n��<A:�<M��<��<�I�<���<♻<���<�9�<�Ŵ<�-�<o��<�ʬ<��<�y�<��<�x�<�<�ԝ<���<��<���<�̕<��<�L�<ǉ�<Y��<G��<O��<�<�<\��<�#�<ct�<�{<�%v<��p<��k<�g<�Qb<��]<˅Y<�rU<J�Q<�M<�vJ<�G<�|C<��?<K�;<�n7<�2<'�-<N}(<u#<չ<�h<�;<�;<Lj	<��<!X <y:�;�9�;|��;���;ë�;��;���;��;霽;�
�;�ի;m�;@�;�ڍ;'Ѓ;�=t;5�a;��P;�l@;Ό1;�#;"�;��;��;��:b��:���:)��:�O�:�7�:VV�:&Î:X�u:��L:��$:ּ�9��9�s9��96B;8�5��B���t���#���4���;���=�}�B���Q�H<r���lp��գ�׵��22�zR���q�Ko��z{��0柺����j����6�������ĺXRź�Fƺ��Ǻ%�ʺ^к��غ�㺋��`� �3?	�m���:�'�!�V�(��/��j4��9���<���?� B���C���D�
�E���F��I�oiL�w-Q�idW���^��Kg��4p�('y�$܀��τ��]��)����>�����������X=�����~����  �  �?=�=��=!�=.c=��=�z=�=�N=�� =0 =X�<��<�E�<A��<��<۫�<�m�<�M�<�B�<?�<�2�<j�<���<�N�<$��<���<u��<7��<���<��<2�<gk�<Ÿ�<��<	~�<@��<r�<��<B��<cj�<Z7�<��<���<��<9
�<�g�<2��<^��<�~�<R�<�#�<��<��<��<�B�<՚�<��<���<ya�<�(�<���<ǻ�<{f�<���<�.�<S8�<��<��<���<�8�<�f�<y��<���<���<
��<��<.(�<�9�<�L�<�i�<G��<���<6�<�L�<�{�<���<`r�<)�<���<��<�I�<Dx�<���<�<:8�<���<=D�<k�<%�<h�<|�<f�<��<[�<�g�<,��<[��<�x�<�(�<�<�)�<3��<�|<r�v<�	r<c>m<`�h<�c<�a_<~�Z<q�V<jzR<>�N<��J<�G<isC<��?<��;<lI7<*�2<n�-<h&(<��"<S�<�`<0�<&�< �<4<�`�;�;�;T��;��;�
�;Ŝ�;�!�;�\�;P�;O0�;&��;e�;G�;�-�;~s�;���;�w;uf;[V;߇F;R�7;��);Z�;��;�x;=�:L_�:���:x�:��:���:�ڟ:��:�`q:�eF:;�:���9i�9F�9@38zp�|5���<�u^�6�l�=�l�xFc�N~X�bT�P�^��}��8��K��4���!H/��K��df�k�~�;��e��y��T����d��h��FM��.뾺9eºz.ź�Ⱥ9�˺�Ѻ��ٺ6%��C���������*��(�&���.��w5�n";�U�?���B��E�$CF��F���F�\G�V�G��I��M���Q�!�W�,_��g�w.o�bw�Mw~�����妅�`s�����L���"̏��ԑ�싓��	���  �  �5=R	=��=ژ=tF=��=�[=��="=�x =`��<�n�<*]�<�w�<���<XB�<���<���<���<g��<���<'��<V��<��<��<'s�<���<���<���<
�<D�<���<��<�V�<���<�0�<���<�<�q�<���<ϊ�<5�<���<3��<�I�</��<!.�<[�<�Y�<�1�<|��<��<�l�<�H�<H�<2r�<���<�N�<	��<���<1��<���<�n�<�&�<~��<��<��<���<�i�<���<r8�<���<���<o �<�g�<���<���<J��<���< ��<j��<r��<���<��<	0�<P�<vY�<>�<��<�w�<�˱<���<��<V&�<bF�<��<R�<r�<�1�<m#�<�C�<[��<��<�a�<�Α<&�<�Y�<\b�<�=�<��<戅<;�<V��<�S|<�w<I�r<Nkn<��i<�Xe<�`<$\< �W<<(S<D�N<m�J<��F<�(C<�G?<7;<#�6<K"2<7-<�'<��!<<F<�<u3<�<�c<��;�>�;)�;�z�;5E�;�/�;���;�P�;��;R4�;Ƭ�;��;�H�;9��;���;ֺ�;�yz;�Wj;��Z;��K;7=;X�.;�,!;nG;�;sM�:��:���:��:�d�:j�:t �:FJ�:Pi:��<: �:���9c�[9{�8��v�4�$��.p��5��޲��Ƙ��P���A�������pu��d|��錹������̹����wo���/�$'H�|^�8�q�����������������r]���!���J��kQ���!����ź�9ʺ��κպ%�ݺ��躎��t�M������"�b�+��_4��;�G�A��F�I�H�-eJ���J��RJ��I�AUI���I�P�K���N��S���Y��~`���g�>o�M�u���{�)ƀ��Q���ǅ��C��ӊ�k������A>��2<��Fꕻ�  �  "=��=˳=0r='=^�=%3=Y�=�� =�> =�< ��<���<A��<��<݋�<H�<h4�<E�<Bh�<c��<��<7��<A<�<��<�&�<�f�<��<}��<H�<nb�<y��<�O�<���<�R�<���<:�<�q�<���<G"�<��<� �<��<�b�<���<-��<��<��<>�<���<	��<s0�<���<���<�<��<E�<)��<�X�<S:�<_2�<�,�<��<���<W`�<��<7��<E��<e+�<��<�$�<���<��<�s�<���<-�<�a�<"t�<g�<E�<��<t��<���< ��<���<c�<�<��<���<�+�<�z�<���<N��<!��<鲥<Kۢ<�.�<E��</x�<�s�<B��< �<�x�<_��<bt�<�ҏ<��<��<H�<Y��<]J�<��<���<`x|<�x<7�s<Zo<��j<Zf<��a<_]<�TX<�S<�O<\�J<a�F<��B<Q�>< �:<�A6<��1<�h,<��&<� !<�,<+5<�a<O�	<1�<7��;�5�; ��;���;\�;&t�;&��;��;���;��;A�;-h�;Zy�;�Y�; K�;��;�$�;�o|;TYm;׵^;5P;'�A;3;1�$;Ҿ;��	;1��:S��:e��:���:b��:x�:��:�<�:p�^:1:E�:�;�9]9��]����� ����������Ĺ���������㤹3���)|��v������b��b�߹������2��<G���X��g��Su�jn���ٕ��V�����⯺�+��>$����Ǻa�ͺ�?Ӻ�ٺmg����	��д�y��uB��&�-\0���9��sA���G���K�adN��UO�	O���M�B�L��L��bL��N��SQ�V��[�1gb�'i�-vo��:u��Jz���~�Yx��;�������ݤ��҆���|���T���ᓻ����  �  �=��=�=�K=��=�=\=�p=�� =� =���<�S�<?%�<<-�<�s�<��<���<d��<���<`�<22�<�E�<�1�<b��<px�<O��<q!�<�_�<���<���<�p�<���<��<�/�<s��<�+�<��<���<i��<:=�<^��<D�<D��<�"�<���<P5�<���<,��<��<���<�,�<���<�h�<u#�<V	�<
%�<|�<�<|��<���<6��<���<.��<b��<%�<_�<Vk�<<@�<k��<)��<�	�<���<p �<���<f,�<���<���<���<t��<A��<�O�<A�<���<���<�̾<�ϼ<�ɺ<��<�]�<u߳<,�<�J�<�I�<�<�<�9�<�T�<ꞟ<j"�<`�<[�<�"�<݋�<X�<���<�<�<6��<+��<a��<�]�<��<
��<�r�< �|<�Dx<%t<	p<��k<�Vg<a�b<?�]<��X<a�S<3O<X�J</dF<�DB<�2><�
:<��5<��0<e�+<�D&<�l <�b<jP<�`<$�<�|<n�;���;�V�;l��;���;��;�,�;�2�;���;�~�;���;-)�;/V�;�j�;n��;@�;R�;c�};�ro;xa;F\S;��D;6�5;�';}h;��
;7��:o��:i��:��:-�:��:s�:�v~:�dT:l_&:m��9��9���8E���/�]�6	��(�˹��แ
�2�޹�Ϲ|���i�������ʥ��P��%�ι�]������"���6�j�G���U��@a�	�k���v�sU�����D��� $��'�����&���S�ɺT�к%�׺^�޺�N�ښ��} ��@	�$W��G��t)�`04���=���E�A4L��sP���R��ZS�i�R��,Q���O�ǲN�X�N�y�P���S�rX��"^��Rd�{j��'p�Uu�I?y���|�d%��X��BT��U�� +��%{��~������b���  �  ��=ط={v=�/=��=�p=1�=S=S� =���<#`�<� �<���<b��<}�<��<�g�<g�<���<C��<,��<�
�<���<w��<?�<^��<���<6�<���<F��<uu�<{�<��<�f�<��<�k�<��<���<�<MJ�<ӎ�<���<�h�<���<���<���<�V�<#��<m|�<;F�<k��<`��<��<T��<Y��<���<��<���<�~�<)u�<J��<"��<&��<�L�<��<z&�<�3�<?�<���<L\�<���<[��<�-�<���<>]�<c��<^�<�"�<)�<��<l�<��<���<���<��<'��<���<�q�<�%�<��<��<}�<��<���<�<��<�B�<nÜ<��<���<NΖ<�>�<5˓<+^�<'�<vE�<}�<r��<jf�<)�<Cބ<̖�<H_�<�}|<�gx<�lt<�kp<�Bl<q�g<m'c<'8^<�'Y<eT<W7O<֎J<�&F<�A<��=<��9<y65<$z0<�W+<q�%<��<9�<_�<@�<2<�<���;�i�;���;;T�; b�;���;�*�;G<�;���;���;��;�D�;���;���;�*�;7�;�]�;Gb~;m�p;�c;�CU;X�F;��7;�v(;�Y;d;�"�:�7�:H�:ി:��:s�:�i�:�w:��L:�:�k�9`Bp9ćF8�7��@Ņ�8���Ȱ�i���ّ���l���|�̹ޠ��P[��kT��c�¹(�ܹQ���ص���'�c�9���H�GuT��]���e���o�G�|�������_v��$_��$���i�ºR�˺��Ӻ}�ںT�ẓ���8��\O�u��C�u[ ��+�1�6�]�@���H��,O�eS�a�U���U��U�2VS���Q�X�P�]�P��\R�$�U�2Z���_�/�e���k���p�!u���x�5�{�`�~�����R�����fZ��L医fs��S���ħ���  �  /=�=�x=_&=��=\=u�=Q=�� =b =���<���<��<���<G$�<���<�K�<D�<i
�<��<s �<���<,��<uq�<z�<dw�<=��<;0�<<��<���<_�<m��<�`�<��<r^�<���<$�<%r�<ѻ�<��<�_�<��<�3�<��<��<�z�<R��<g��<���<��<^��<xb�<�,�<_	�<=�<�&�<�t�<���<��<�G�<0�<z��<���<'.�<۞�<���<���<��<]��<�E�<���<�t�<�<���<���<�R�<��<���<H��<қ�<7z�<gV�<�7�<�!�<��<��<��<Y��<�h�<���<^�<$��<�۪<	�<{>�<<9��<<��<�X�<Q�<t�<r��<_�<t�<>ϐ<'�<pC�<@P�<�?�<��<��<1��<=w�<n�|<pVx<.t<��o<גk<$g<%�b<�]<z$Y<ulT<Y�O<MGK<��F<&�B<P><��9<�l5<ɩ0<��+<�T&<8� <�3<j�<�<��
<��<�<���;!��;o��;c�;s��;m�;���;�2�;���;�W�;}Q�;|
�;\��;l�;�`�;���;�)�;��w;��i;t~[;�CM;��>;)�0;�#;��;l�	;�#�:���:���:;��:�+�:nϟ:.k�:՛o:�LD:o�:\��9�
�9���8���+7 ���P��b��#L�����������ܒ����s���w*����T�ùt�F�R��ħ'��@8�DEG��U��nb�Bep�����ڈ�ɒ� j���=���ò������źeEκR�ֺ��ߺB������*��.
�g0�|��Y\&��/�8�5x?��fE�d�I�g�L�XwN�60O�-YO��dO�K�O�g�P�d�R�!+V�hQZ��5_���d�q�i��o�b�s�*Mx�r|�gH��Br���Մ��~���c���f��hi��9L��d����  �  =��=y}=�+=��=/b=��=�W=D� =�  =t�</��<���<���<C;�<I��<a�<.1�<��<�<A�<O��<���<�}�<
�<ԁ�<Y��<:7�<��<��<9[�<���<QU�<���<8N�<��<��<Le�<X��<�<Y^�<h��<�9�<S��<�#�<���<-��<���<���<5��<���<�s�<�?�<�<��<�=�<���<�<���<�Z�<�"�<��<ơ�<;�< ��<`��<���<���<p��<0K�<��<is�<M��<�y�<M��<C�<���<��<ܡ�<@��<5q�<bQ�<�6�<�$�<��<<
�<>�<A·<<t�<��<k�<a��<o�<��<R�< ��<��<-��<�o�<g�<���<}˕<�#�<���<qݐ<c$�<�O�<@\�<K�<{"�<��<O��<�x�<��|<`Ix<�	t<K�o<sk<Bg<�pb<��]<kY<�]T<��O<�HK<K�F<��B<4b><�:<��5<��0<(�+<5p&<�� <AU<�<�5<��
<1�<�E<��;�9�;t�;�c�;c��;Ѫ�;}2�;3h�;�1�;���;�}�;,1�;�͢;�}�;�c�;1��;��;��w;25i;= [;��L;�>;�f0;��";��;Ӳ	;�O�:'%�:�v�:
��:��:��:34�:�Dq:�F:(�:!6�9eވ9��8���Yt�ZAE��{����!ݒ��G��9莹�o���N��I������ ���u���4�2��1O'��`8�4�G�S0V� d�Jr�����߉�����f'��$¨����������ź��ͺ$ֺ�ߺ�3�C1��6����	�]��X8��%��/�@u7�V�>�
�D�KI�wL���M�t�N� �N� �N��WO��}P���R�A�U���Y�c�^��Id���i�Uo���s�Q�x�G�|�l~��)���k��u���ޚ��<���C����W�������  �  �=��=G�=�:=��= s=��=>k=�� =v8 =�<�<��<>�<F2�<�~�<n��<���<�j�<kP�<&D�<�8�<& �<Q��<	��<�-�<���<���<�I�<��<���<"O�<���<v2�<+��<��<q��<���<]>�<c��<���<�X�<��<wH�<u��<�>�<(��<���<=�<l�<��<���<���<�v�<?Z�<[�<���<���<�D�<D��<��<	T�<�<L��<S_�<���<S�<o�<���<��<zY�<4��<�m�<c��<B\�<X��<h�<=M�<�l�<vs�<-i�<�U�<�A�<d3�<z+�<�'�<k �<��<�<���<�#�<A��<Jݭ<��<)M�<6��<vܢ<YO�<n�<���<B��<Dė<��<JT�<b��<#�<aI�<�r�<_}�<�i�<;=�<� �<���<�|�<Є|<%!x<J�s<�so<�k<��f<�b<Co]<0�X<�0T<��O<KK<'G<x�B<�><B:<��5<Q1<1,<ϼ&<qF!<x�<�"<V�<sj<�q<�<;�;:�;��;":�;8��;pX�;b��;g��;��;~�;���;���;a�;���; i�;�h�;@��;�wv;�g;��Y;�@K;�=;9/;��!;�=;w�	;l��:�"�:���:[_�:
״:ا�:Zf�:g�u:dK:�l:���9Y��9�9�[�7�5���#�K�Z���{��|ͅ��ă��c����B]�������5����ٹ����/���u&�p�8��I� �Y�ʾh�&�w�J���팺�w��If���U���߳�d���`�ĺ��̺r�ԺBݺ�<纁󺓎 �R���r����3$�&>-���5�q�<���B�G��J���K���L�QM�l�M�� N�b\O��Q�y�T�*Y�m^�ͣc��Zi���n�+7t��!y�w�}��!��n��
߅�8}��B������ڐ�l}�����  �  O =��=��=�N=��=��=/=	�=�� =\ =6��<s�<Bt�<���<}��<�_�< �<���<���<Z��<�u�<xV�<!�<���<*Y�<#��<��<�`�<���<U��<�7�<:��<g��<c�<���<�6�<��<��<Id�<m��<�K�<���<uZ�<���<�c�<���<��<fF�<xP�<x>�<�<&��<o��<,��<���<���<�6�<?��<�;�<���<���<aW�<��<Ȓ�<"��<A7�<�A�<��<���<�j�<��<}_�<=��<�)�<O�<���<���<|�<�'�<*�<'�<R%�<�(�<-1�<�:�<�=�<0�<��<���<�R�<�°<��<�Z�<S��<U�<p;�<ƴ�<'S�<g�<u
�<2 �<zT�<���<��<�>�<�}�<���<��<���<�a�<��<p͂<}�<�b|<j�w<`s<t�n<�wj<��e<\qa<K�\<�ZX<��S<ĄO<�CK<�G<��B<��><m�:<�6<�`1<De,<T+'<��!<�C<��<�b<K1<�C<��<���;J��;�i�;��;���;�W�;���;q��;P��;`Ǽ;p��;�(�;��;Yߚ;4\�;��;��;��t;�e;vW;��H;	�:;�E-;*c ;�R; 4	;��:�[�:���:H��:w��:���:ay�:W�|:�jR:��':�O�9˫9��F9���8jo��Nf޸�x(���L��M_���e��jf���g���o�&5���[������3йs.��3���%�O:���M�P�_�<�p��������x瑺�����!������s��+5��hĺ�_˺#�Һ��ںϋ�<:���x��������E�!��*�^�2�9��M?���C��G�� I�g]J�VK�%�K��^L�t�M�P��fS�8�W�H�\�8�b���h���n��t�N<z��e�A.������F"������T���펻9p��;ʓ�����  �  5$=	�=&�=�b=[=��=�+=9�=�=�� =	��<��<���<�<Gl�<*��<(y�<0�<���<���<���<��<�V�<+��<^��<���<�9�<�t�<p��<���<p�<#W�<���<�<�c�<���<�4�<c��<��<֢�<j2�<F��<�g�<���<W��<���<�I�<~y�<q��<��<of�<�H�<�1�<+�<�<�<!l�<���<�'�<���<�N�<���<:��<�C�<��<.�<wd�<5j�<z@�<���<Rv�<b��<E�<a��<���<c$�<\�<���<`��<���<���<(��<��<u�<�.�<�H�<�W�<mR�<�0�<��<���<���<�Y�<S��<���<�J�<y��<�4�<�מ<���<m��<���<��<���<C;�<��<��<c׍<dڋ<�<�<�5�<�ׂ<�t�<'|<%qw<��r<�2n<�i<�e<�`<�#\<��W<pS<+?O<,)K<�%G<v%C<�?<�:<p6<��1<f�,<C�'<^T"<��<H�<�E<�+<NM<�<���;W��;]-�;?�;�7�;t�;C��;&��; V�;߆�;@I�;>��;��;���;�)�;��;1�;#Jr;��b;��S;�zE;D�7;N�*;�H;i�;�|;���:�P�:M��:��:DA�:e��:q��:��:Y�Z:�S1:��:v��99)[9tX8c�3���Ѹ?��3�*�_28��b?��<F���R���j�f�������ǹE�T���&��'=�;7S��g��r{�����Z珺&����$���N������.�UU��@Jĺ�>ʺ/�к�tغH��47�!������l��#����K&'���.��5�?(;�ձ?��"C�f�E��:G��YH�nII��cJ��L�N���Q��}V��[��b���h�Y6o���u���{��ۀ�ڞ��(E���ֈ��Z��Bˍ����vL��;L��?$���  �  e!=�=ն=Wq=�=^�=C=��=�;=�� =	- =U^�<y�<���<Y�<r�<���<���<�d�<�/�<f��<���<���<�$�<���<u�<#M�<z{�<���<'��<��<_�<eB�<��<���<6F�<��<v7�<P��<fa�<y	�<���<�g�<�<���<��<�m�<G��<`��<6��<��<���<h��<H��<���<���<�N�<l��<�1�<���<�W�<^��<l��<���<�V�<Ć�<-��<�V�<���<|t�<7��<��<:U�<@��<���<���< �<�!�<�B�<f�<���<Һ�<���<d�<�I�<pe�<&i�<�M�<��<v��<6.�<=��<��<�W�<��<�6�<Yġ<l�<1�<��<��<y'�<PQ�<%��<J��<��<��<>��<Z݉<ל�<,B�<6Ղ<@^�<
�{<Y�v<Wr<4Mm<��h<Bd<��_<8[<��V<�R<��N<��J<�G<m4C<-:?<!;<��6<}2<\--<�(<��"<�<�c<�?<�B<nw	<]�<Ό <���;��;��;M��;B��;���;�|�;��;��;�ȵ;�;��;��;[��;|��;��;�:o;�,_;��O;5vA;n�3;>';ɖ;��;7K;+��:�w�:ȝ�:��:�O�:��:%v�:��:J�b:;:�:���94ݠ9')O9�8���7*�1#���g�% ����&��29�K1U�}�~��������4a칍y�A(��A�\[��r��v�����*���ɠ�e����Ư������5f��{ź��ɺp�Ϻ��ֺ#�ߺ��꺚����`�[�B��Դ��w#���*���0���6��;���>��A�/�C��E�G�i�H���J��;M���P��U��9[�u�a��h���o��#w�~��T��f��
A��"犻�Z��ٙ�����=r��"��y����  �  r=��=ķ=�u=�#=��=R=s�=�Y=!� =o` =���<-�<]E�<��<-�<���<��<���<�{�<�7�<j��<r��< 8�<��<�<	M�<�o�<���<,��<̔�<3��<���<�<]P�<���<F+�<b��<�[�<w�<r��<w��<<U�<e�<��<�!�<~�<ٺ�<"��<���<���<w��< �<�,�<�Y�<��<"��<�F�<���<�.�<E��<a5�<c��<��<m�<g��<ҏ�<�X�<���<�_�<��<���<&�<C�<f2�<�J�<Mg�<��<��<���<W&�<�k�<δ�<��<]7�<�_�<�k�<"V�<v�<cĳ<Q�<�̮<t@�<2��<02�<���<�W�<��<�ȝ<V��<^��<4��<m��<�Ɠ<S�<U
�<��<l�<��<?��<J<�<5��<(6�<5M{<�4v<�/q<�Gl<=�g<��b<Ts^<',Z<�V<�R<�NN<ӔJ</�F<�C<9?<� ;<��6<�52<�g-<Gn(<Q\#<C<u3<�9<�_<�
<�<ɾ<T�;Z�;�R�;��;V��;�X�;��;cb�;�e�;���;��;��;҄�;�;ӱ�;�+};�k;�[;NxK;��<;<�/;�g#;�d;�};��;���:�{�:|z�:�,�:��:��:j
�:ZR�:�h:$�C:��:��9h�9�֋9�%:9si�85	8?�k���e�������긋S�j�'��H��v�[0���p��c;���VZ,���H���d�C���7���f��sQ���ꩺz6���B���'���$��A�ú=�ƺپʺ�Ϻ�WֺZ�޺��麓J��?/��	��B����7���e&��^,��1��\6�\_:���=�j�@�E�B��
E��&G���I� �L��gP��BU��#[�]�a�lbi��5q��y��h��'��om��A|��7��ܙ��9���Pe���ٔ�����6���  �  O =��=w�=�n=�=,�=�V=��=p=�� =� =�% =���<���</�<w��<�	�<��<��<ٹ�<�_�<��< ��<�4�<��<� �<�6�<�O�<S�<SJ�<D@�<�>�<bN�<�u�<s��<�<���<'3�<��<1��<���<�^�<�/�<C��<ȑ�<9�<�w�<z��<��<x�<l)�<�I�<�q�<��<���<�)�<�y�<���<�.�<���<��<1j�<���<�+�<�m�<$��< ��<D�<,��<8�<t�<���<���<���<���<��<y��<��<s�<�b�<��<0�<�m�<�ƿ<D�<�C�<�V�<EG�<e�<�ų<�`�<�<y�<A�<+��<T:�<L�<���<NZ�<@(�<��<��<�<���<7�<Z�<i�<v
�<݉<��<]!�<���<��<��z<nu<>p<P2k<WUf<Ѯa<CB]<�Y<U<NQ<h�M<J<)�F<��B<?<' ;<�6<02<Ox-<�(<�#<��<B�<Y!<hm<�<ZM<)�<2,�;t��;���;���;	J�;?��;)-�;�h�;VP�;!͵;7ج;�~�;�ݙ;e�;�n�;G�y;��g;ֺV;�F;�C8;�+;2P;|�;��;(d;���:�O�:l �:$-�:�x�:�ī:�?�:"J�:Y�l:A%J:2w):)O:���9\I�9uȁ9��39��8�;8гж��N��Y������J���gG���x�"����ùZ�j
���2�~�Q�op��}�����P檺{r���3��NK��e�ºl�źͭǺ��ɺ��̺�(ѺZ׺��ߺ���%���ٔ��{�Sh����{�tm"��'��-���1�E.6�W:���=�f�@�ߔC��PF��6I�b�L�s�P���U��[���b��j��s�ֈ{�����A����Ҍ�����󑻜Փ��N��1p���V��S%���  �  ��=��=ę=�]='=��=)R=-�=w}=�=m� =�V =)��<V�<��<��<zz�<���<b�<���<�u�<E	�<��<��<��<U��<��<��<��<d �<J��<���<p��<B��<"%�<5��<�<���<?s�<-N�<Y5�<��<���<n��<8l�<���<�\�<���<���<G�<�K�<��<|��<g�<�[�<J��<?��<�J�<ʘ�<��<F:�<؍�<P��<8'�<m[�<q�<�^�<!�<Ӧ�<� �<T0�<�?�<�:�<-�<� �<V�<�.�<�R�<���<���<�?�</��<��<��<3۽<��<�.�<�$�<���<���<�^�<���<䠬<�F�<��<��<�`�<4�<�۞<8��<j�<s@�<�$�<��<��<��<�	�<T��<-��<�i�<#��<Gb�<�r<c	z<؟t<Lo<�!j<=0e<f�`<V\<��W<�T<wP<3�L<�I<�F<&|B<�><۷:<Yy6<�2< d-<d�(<��#<g0<�<5�<�Z<|�<�[<Q�<���;�W�;
��;��;��;��;o�;��;��;Q�;�E�;�̢;I��;f�;n�;��v;� d;�zR;�TB;�3;�&;eE;�Q;�;�� ;���:)�:�h�:���: ��:O8�:"A�:n�:�n:;�N:A�0:&�:��9��9��9\�u9F�*9x��8l�8����F��)[��� ��vO�₹3���	͹�=�������:�ʚ[���|�5�������w��V/��C���}�ºSEǺ�ɺ�b˺�h̺��ͺZ�Ϻ��Ӻ��ٺ��zn�;���Ӎ����/��������
$���(��-�[|2�Z�6�6;��?�ުB�qF�tI�p.M���Q���V��\��:d�bl�g'u�\1~�,��� ч�ⱋ�������;������8��P�������>���  �  	�=}�=�="G=I�=}�=EG=��=��=�&=�� =�} =b. =���<# �<|�<���<2�<]��<��<0}�<���<g��<���<
c�<[��<���<���<���<���<Ӎ�<�l�<P^�<cm�<ɡ�<���<���<L7�<"�<���<2��<X��<���<ȍ�<><�<<��<[7�<���<D��<Y�<�^�<��<�<�`�<���<��<5h�<���<���<�)�<e�<O��<=��<��<m=�<DJ�<`1�<��<�o�<<��<���<���<��<U��<���<d��<��<���<T�<�e�<���<�O�<���<!@�<���<߻<���<���<]ӵ<(��<�O�<��<&��<�u�<9�<� �<fǣ<
��<�F�< �<���<�|�<�J�<�&�<��<��<��<�ʋ<5��<I:�<]��<1&�<��~<�cy<��s<@on<�,i<�*d<	u_<v[<�W<�:S<��O<�HL<�H<��E<�
B<ZQ><�Z:<'6<��1<7-<��(<1$<�t<��<!�<�<�<�;	<�<s= <0��;���;�4�;��;7��;���;��;U�;姴;D��;���; �;��;���;�s;_�`;ߪN;Q>;w�/;_�";�;;,�;��:��:���:�>�:��:��:<��:*��:<�:(�n:�Q:\#6:��:��:���9��9a �90�\9�i9��8U�}5�+s�1��(�#�]����kͮ���ع�����"��%C��pe�����������p���u��@�ĺ��ʺ9}κ�Nк��к�%ѺۺѺtӺ��ֺe~ܺ�&�ȡ��j�����ײ��B�(���p��)�s� ��%�Qt*��z/��4�y_9�+�=��6B�z2F��J��*N��R�� X�l^���e�vIn��[w��d��^��܈������������E���㗻��������x��^���  �  h�=D�=�i=(1='�=R�=�:=X�=�=�0=�� =<� =�P = =�p�<���<<�<�e�<���<��<E|�<���<�e�<���<�9�<���<��<8��<B��<!v�<E�<B�<��<N
�<�9�<ʖ�<&"�< ��<���<���<���<���<<��<�\�<@�<X��<��<�m�<���<I�<g�<$��<J0�<U��<Y�<lg�<��<R��<�+�<>W�<���<٫�<���<� �<t�<�"�< �<k��<�<�<��<_��<��</��<�f�<�D�<3�<�9�<_�< ��<��<~�<��<���<��<�g�<.��<͹<>˷<F��<Jy�<<�<D��<�Ŭ<Ԕ�<oj�<�@�<��<�ڡ<���<G�<���<ܥ�<�a�<�,�<��<p�<�ˍ<s��<�g�<��<4��<5��<�l~<��x<?@s<0�m<�ih<�[c<$�^<�AZ<^;V<,�R<�
O<�K<prH<�E<��A<��=< :<_�5<=z1<w-<ł(<�$<��<�D<=�<�<"P<t�	<L\<�� <9f�;=X�;4��;��;}��;\�;�"�;軼;� �;�֪;�7�;�4�;��;���;�q;�];)�K;�#;;�s,;�;V�;xi;ut;-��:X�:U]�:�D�: L�:PZ�:��:֖�:�ͅ:�m:�5R:�|9:�d#:S3:���9T��9��9�9�.9NI�8r�r7�6^��:���2��l�:����i���M� ���e)�!�J���m�Dň������������ ú'n˺�Ѻ�GԺ��պ��պ�1պ�Oպ��ֺ�ٺ�Mߺa��d�ﺵ3���z�������_�����g!�s��	#���'��F-�g�2�u8��D=��B���F���J��6O��S��}Y�t�_��yg���o�Fy��{���O���늻F�����a���Tᗻ�j��p\��Aݚ�M��xV���  �  =�=^=�X="!=v�=��=�0=��=�=�5=�� =ҩ =f = =���<���<�@�<���<
��<D�<Fx�<f��<�P�<G��<��<Cb�<���<��<)x�<�J�<��<:��<(��<5��<��<~S�<r��<W��<�x�<�p�<Ft�<�t�<�d�<�9�<	��<�<|��<'V�<���<��<&i�<,��<J�<���<�3�<>��<��<Q%�<�P�<�q�<���<���<���<���<z�<��<���<&��<��<De�<S��<�y�<X�<�,�<��<���<r��<��<ia�<���<8E�<���<[�<5ھ<<A�<���<���<)��<׏�<b�<\,�<���<�ʬ<��<N��<�g�<A�<�<hƟ<ir�<w�<Ͻ�<�m�<-�<
��<֏<���<>��<�H�<��</l�<�ʁ<�~<L|x<�r<RIm<��g<F�b<!^<S�Y<Q�U<�R<q�N<�WK<�H<�D<cYA<"�=<[�9<C�5<vF1<��,<Vk(<�$<��<�q<�:<q�<?�<kG
<P�<�<���;���;���; ��;�d�;��;���;�J�;��;�T�;p��;Ӟ�;GL�;e�;�to;��[;��I;�9;d*;�;��;b�	;�;�(�:��: �:Q#�:DG�:Pr�:�:�%�:ń:b�l:n�R:�K;:��&:��:��:���9bt�9!\�9%RA9�u�8?M�7S<W�����:��_x�����)��u�����.���O��\s��狺֎���ƭ�ֻ��3ǺR�ϺPպnغ0�غL�غ��׺��׺��غ�ܺ2X���4�񺐐�������,�������-�����B}!�{&�D�+� �1��a7�8�<�?B���F�4mK�$�O��T�-|Z�a�Q�h��.q��z�5�� ���ҋ�����ƶ��F똻"g���E��/����ۛ�a����  �  `�=�x=�R=L= �=��=%-=[�=��=s7=b� =B� =m =' =8��<]�<�M�<���<V��<p�<}v�<>��<�H�<���<��<V�<�}�<��<,j�<�;�<��<I��<���< ��<)��<�<�<���<2��<Ne�<�^�<6d�<Of�<W�<�,�<��<�s�<@��<MM�<��<��<xi�<���<�R�<���<�B�<���<���<E4�<�\�<�z�<o��<V��<���<B��<���<���<T��<�<��<�W�<Zs�<�h�<�E�<��<���<b��<���<G�<lJ�<<��<_1�<ý�<�J�<k˾<�3�< {�<C��<���<���<TY�<g&�<X��<̬<���<���<�t�<gP�<��<�֟<Ӏ�<�"�<�Ř<�q�<�,�<I��<�Ϗ<ɪ�<�}�<S=�<�߆<�_�<.��<M�}<r[x<H�r<3!m<��g<m�b<��]<"�Y<P�U<��Q<�yN<�5K<�G<�D<?A<:�=<w�9<s�5<f31<s�,<Zb(<�$<�<t�<2Q<<�<�i
<��<�7<{�;c��;��;���;�R�;Z��;Ȝ�;�!�;yY�;&�;�{�;i�;��;��;��n;�K[;�I;�d8;9�);A�;.;�	;�[;V.�:���:pH�:e_�:ϋ�:B��:oH�:���:�_�:.Kl:ƖR:��;:��':4M:�q:x�9���9@!�9ԅG9wa�8{G�7&�U��t����=�J�|����S�ù������/��XQ�gYu���nƞ�����=����Ⱥ�ѺF�ֺRٺ!"ں*�ٺ��غz�غu�ٺ��ܺ�iX�F5�������������2~���J� ���%��{+��I1��$7�_�<�aB�"G�i�K��FP�H:U��Z� ba�@�h�5�q�){��v��~i���"���l��������F��𽚻Q���g���1���;���  �  =�=^=�X="!=v�=��=�0=��=�=�5=�� =ҩ =f = =���<���<�@�<���<
��<D�<Fx�<f��<�P�<G��<��<Cb�<���<��<)x�<�J�<��<:��<(��<5��<��<~S�<r��<W��<�x�<�p�<Ft�<�t�<�d�<�9�<	��<�<|��<'V�<���<��<&i�<,��<J�<���<�3�<>��<��<Q%�<�P�<�q�<���<���<���<���<z�<��<���<&��<��<De�<S��<�y�<X�<�,�<��<���<s��<��<ja�<���<9E�<���<[�<6ھ<>A�<�<���<+��<ُ�<b�<^,�<���<�ʬ<��<O��<�g�<A�<�<hƟ<ir�<v�<ν�<�m�<-�<	��<~֏<���<<��<�H�<��<-l�<�ʁ<�~<J|x<��r<QIm<��g<F�b<!^<S�Y<R�U<�R<s�N<�WK<�H<�D<fYA<%�=<^�9<F�5<yF1<��,<Yk(<�$<��<�q<�:<r�<@�<kG
<P�<�<���;���;���;��;�d�;��;���;�J�;��;�T�;j��;͞�;AL�;_�;wto;��[;��I;�9;d*;�;��;^�	;�;�(�:��:�:O#�:CG�:Or�:�:�%�:ń:b�l:n�R:�K;:��&:��:��:���9bt�9!\�9%RA9�u�8?M�7S<W�����:��_x�����)��u�����.���O��\s��狺֎���ƭ�ֻ��3ǺR�ϺPպnغ0�غL�غ��׺��׺��غ�ܺ2X���4�񺐐�������,�������-�����B}!�{&�D�+� �1��a7�8�<�?B���F�4mK�$�O��T�-|Z�a�Q�h��.q��z�5�� ���ҋ�����ƶ��F똻"g���E��/����ۛ�a����  �  h�=D�=�i=(1='�=R�=�:=X�=�=�0=�� =<� =�P = =�p�<���<<�<�e�<���<��<E|�<���<�e�<���<�9�<���<��<8��<B��<!v�<E�<B�<��<N
�<�9�<ʖ�<&"�< ��<���<���<���<���<<��<�\�<@�<X��<��<�m�<���<I�<g�<$��<J0�<U��<Y�<lg�<��<R��<�+�<>W�<���<٫�<���<� �<t�<�"�< �<k��<�<�<��<_��<��</��<�f�<�D�<3�<�9�< _�<!��<��<~�<��<��<��<�g�<1��<͹<A˷<I��<My�<<�<F��<�Ŭ<֔�<pj�<�@�<��<�ڡ<���<G�<���<ڥ�<�a�<�,�<��<n�<�ˍ<p��<�g�<��<1��<2��<�l~<��x<;@s<-�m<�ih<�[c<$�^<�AZ<`;V<.�R<�
O<�K<urH<�E<��A<��=< :<e�5<Cz1<}-<˂(<�$<�<�D<?�<�<#P<t�	<K\<�� <4f�;6X�;,��;��;r��;\�;t"�;ܻ�;� �;u֪;�7�;�4�;��;���;�q;ٻ];�K;�#;;{s,;�;N�;qi;ot;$��:Q�:P]�:�D�:L�:NZ�:��:Ֆ�:�ͅ:�m:�5R:�|9:�d#:R3:���9T��9��9�9�.9NI�8t�r7�6^��:���2��l�:����i���M� ���e)�!�J���m�Dň������������ ú'n˺�Ѻ�GԺ��պ��պ�1պ�Oպ��ֺ�ٺ�Mߺa��d�ﺵ3���z�������_�����g!�s��	#���'��F-�g�2�u8��D=��B���F���J��6O��S��}Y�t�_��yg���o�Fy��{���O���늻F�����a���Tᗻ�j��p\��Aݚ�M��xV���  �  	�=}�=�="G=I�=}�=EG=��=��=�&=�� =�} =b. =���<# �<|�<���<2�<]��<��<0}�<���<g��<���<
c�<[��<���<���<���<���<Ӎ�<�l�<P^�<cm�<ɡ�<���<���<L7�<"�<���<2��<X��<���<ȍ�<><�<<��<[7�<���<D��<Y�<�^�<��<�<�`�<���<��<5h�<���<���<�)�<e�<P��<=��<��<m=�<DJ�<`1�<��<�o�<<��<���<���<��<V��<���<f��<��<���<W�<�e�<���<�O�<���<&@�<���<#߻<���<���<aӵ<,��<�O�<��<)��< v�<�9�<� �<gǣ<
��<�F�< �<���<�|�<J�<�&�<��<��<��<�ʋ<1��<E:�<Y��<-&�<��~<�cy<��s<<on<�,i<�*d<	u_<w[<�W<�:S<��O<�HL<�H<��E<B<bQ><�Z:<'6<��1<7-<�(<8$<�t<��<%�<�<�<�;	<�<q= <)��;���;�4�;��;(��;���;ҥ�;�T�;ӧ�;2��;���;��;v�;濃;��s;G�`;ɪN;�P>;g�/;Q�";�;;%�;��:֢�:���:�>�:��:��::��:(��:;�:'�n:�Q:[#6:��:��:���9��9a �90�\9�i9��8~�}5�+s�0�
�(�#�]����kͮ���ع�����"��%C��pe�����������p���u��@�ĺ��ʺ9}κ�Nк��к�%ѺۺѺtӺ��ֺe~ܺ�&�ȡ��j�����ײ��B�(���p��)�s� ��%�Qt*��z/��4�y_9�+�=��6B�z2F��J��*N��R�� X�l^���e�vIn��[w��d��^��܈������������E���㗻��������x��^���  �  ��=��=ę=�]='=��=)R=-�=w}=�=m� =�V =)��<V�<��<��<zz�<���<b�<���<�u�<E	�<��<��<��<U��<��<��<��<d �<J��<���<p��<B��<"%�<5��<�<���<?s�<-N�<Y5�<��<���<n��<8l�<���<�\�<���<���<G�<�K�<��<|��<g�<�[�<J��<?��<�J�<ʘ�<��<F:�<؍�<P��<8'�<m[�<q�<�^�<!�<Ӧ�<� �<U0�<�?�<�:�<-�<� �<X�<�.�<S�<���<���<�?�<4��<��< ��<8۽<��<�.�<�$�<���<���<�^�<���<蠬<�F�<��<��<�`�<4�<�۞<7��<j�<p@�<�$�<��<��<��<�	�<O��<'��<�i�<��<Bb�<�r<[	z<ҟt<Lo<�!j<;0e<e�`<W\<��W<�T<
wP<:�L<�I<�F</|B<�><�:<cy6<�2<*d-<m�(<��#<n0<�<:�<�Z<~�<�[<O�<���;�W�;���;��;ִ�;��;[�;l�;��;�P�;vE�;�̢;4��;S�;\�;��v;� d;}zR;�TB;��3;�&;WE;�Q;�;�� ;���:)�:�h�:���:���:L8�: A�:m�:�n::�N:@�0:%�:��9��9��9\�u9F�*9y��8m�8����F��)[��� ��vO�₹3���	͹�=�������:�ʚ[���|�5�������w��V/��C���}�ºSEǺ�ɺ�b˺�h̺��ͺZ�Ϻ��Ӻ��ٺ��zn�;���Ӎ����/��������
$���(��-�[|2�Z�6�6;��?�ުB�qF�tI�p.M���Q���V��\��:d�bl�g'u�\1~�,��� ч�ⱋ�������;������8��P�������>���  �  O =��=w�=�n=�=,�=�V=��=p=�� =� =�% =���<���</�<w��<�	�<��<��<ٹ�<�_�<��< ��<�4�<��<� �<�6�<�O�<S�<SJ�<D@�<�>�<bN�<�u�<s��<�<���<'3�<��<1��<���<�^�<�/�<C��<ȑ�<9�<�w�<z��<��<x�<l)�<�I�<�q�<��<���<�)�<�y�<���<�.�<���<��<1j�<���<�+�<�m�<%��<!��<D�<-��<8�<t�<���<���<ä�<���<��<|��<��<w�<�b�<��<5�<�m�<�ƿ<J�<�C�<�V�<KG�<k�<�ų<�`�<�<y�<D�<.��<V:�<M�<���<NZ�<>(�<��<��<�<���<2�<U�<c�<q
�<݉<��<X!�<���<��<�z<nu<>p<L2k<UUf<Ѯa<DB]<�Y<U<$NQ<o�M<J<3�F<��B<%?<2 ;<#�6<'02<Zx-<�(<�#<��<H�<^!<km<�<ZM<'�<,,�;j��;��;z��;�I�;+��;-�;�h�;>P�;͵;ج;�~�;�ݙ;P�;�n�;"�y;��g;��V;��F;�C8;�+;#P;o�;��; d;���:�O�:d �:-�:�x�:�ī:�?�:!J�:W�l:?%J:1w):(O:���9[I�9uȁ9��39��8�;8ʳж��N��Y������J���gG���x�"����ùZ�j
���2�~�Q�op��}�����P檺{r���3��NK��e�ºl�źͭǺ��ɺ��̺�(ѺZ׺��ߺ���%���ٔ��{�Sh����{�tm"��'��-���1�E.6�W:���=�f�@�ߔC��PF��6I�b�L�s�P���U��[���b��j��s�ֈ{�����A����Ҍ�����󑻜Փ��N��1p���V��S%���  �  r=��=ķ=�u=�#=��=R=s�=�Y=!� =o` =���<-�<]E�<��<-�<���<��<���<�{�<�7�<j��<r��< 8�<��<�<	M�<�o�<���<,��<̔�<3��<���<�<]P�<���<F+�<b��<�[�<w�<r��<w��<<U�<e�<��<�!�<~�<ٺ�<"��<���<���<w��< �<�,�<�Y�<��<"��<�F�<���<�.�<E��<a5�<c��<��<m�<g��<ҏ�<�X�<���<�_�<��<���<'�<D�<g2�<�J�<Pg�<��<��<���<[&�<�k�<Ӵ�<���<c7�<�_�<�k�<(V�<|�<iĳ<Q�<�̮<x@�<6��<22�<���<�W�<��<�ȝ<U��<[��<1��<i��<�Ɠ<N�<P
�<��<f�<��<9��<D<�<0��<#6�<-M{<�4v<{/q<�Gl<;�g<��b<Vs^<*,Z<�V<�R<�NN<ܔJ<9�F<�C<"9?<� ;<�6<�52<�g-<Rn(<Z\#<C<|3<�9<�_<�
<�<Ⱦ<M�;O�;�R�;���;C��;�X�;��;Kb�;ke�;���;��;��;���;��;���;�+};«k;r[;3xK;s�<;)�/;zg#;xd;�};��;���:�{�:tz�:�,�:��:��:h
�:XR�:�h:#�C:��:��9h�9�֋9�%:9si�85	8=�k���e�������긋S�j�'��H��v�[0���p��c;���VZ,���H���d�C���7���f��sQ���ꩺz6���B���'���$��A�ú=�ƺپʺ�Ϻ�WֺZ�޺��麓J��?/��	��B����7���e&��^,��1��\6�\_:���=�j�@�E�B��
E��&G���I� �L��gP��BU��#[�]�a�lbi��5q��y��h��'��om��A|��7��ܙ��9���Pe���ٔ�����6���  �  e!=�=ն=Wq=�=^�=C=��=�;=�� =	- =U^�<y�<���<Y�<r�<���<���<�d�<�/�<f��<���<���<�$�<���<u�<#M�<z{�<���<'��<��<_�<eB�<��<���<6F�<��<v7�<P��<fa�<y	�<���<�g�<�<���<��<�m�<G��<`��<6��<��<���<h��<H��<���<���<�N�<l��<�1�<���<�W�<^��<l��<���<�V�<Ć�<-��<�V�<���<}t�<8��<��<;U�<B��<���<���< �<�!�<�B�<f�<���<׺�<���<j�<�I�<ve�<,i�<�M�<��<{��<;.�<A��<#��<�W�<��<�6�<Zġ<l�<1�<��<��<v'�<LQ�< ��<E��<��<��<8��<T݉<ќ�<&B�<0Ղ<;^�<�{<R�v<Rr<0Mm<��h<Bd<��_<8[<��V<�R<��N<��J<�G<w4C<8:?<,;<��6<�2<g--<�(<��"<��<�c<�?<�B<pw	<]�<̌ <���;��;��;=��;/��;���;}|�;��;��;lȵ;��;��;��;F��;h��;��;�:o;�,_;��O;vA;\�3;�=';��;��;/K;��:�w�:���:��:�O�:��:#v�:��:G�b:~;:~�:���93ݠ9&)O9�8���7*�1#���g�% ����&��29�K1U�}�~��������4a칍y�A(��A�\[��r��v�����*���ɠ�e����Ư������5f��{ź��ɺp�Ϻ��ֺ#�ߺ��꺚����`�[�B��Դ��w#���*���0���6��;���>��A�/�C��E�G�i�H���J��;M���P��U��9[�u�a��h���o��#w�~��T��f��
A��"犻�Z��ٙ�����=r��"��y����  �  5$=	�=&�=�b=[=��=�+=9�=�=�� =	��<��<���<�<Gl�<*��<(y�<0�<���<���<���<��<�V�<+��<^��<���<�9�<�t�<p��<���<p�<#W�<���<�<�c�<���<�4�<c��<��<֢�<j2�<F��<�g�<���<W��<���<�I�<~y�<q��<��<of�<�H�<�1�<+�<�<�<!l�<���<�'�<���<�N�<���<:��<�C�<��<.�<xd�<5j�<{@�<���<Sv�<c��<E�<b��<���<e$�<\�<���<c��<���<���<,��<��<z�<�.�<�H�<�W�<rR�<�0�<��<���<���<�Y�<W��<���<�J�<z��<�4�<�מ<���<l��<���< ��<���<?;�<��<��<^׍<_ڋ<轉<섇<�5�<�ׂ<�t�<'|<qw<��r<�2n<�i<�e<�`<�#\<��W<pS<1?O<3)K<�%G<%C<?<�:<p6<��1<o�,<L�'<fT"<��<N�<�E<�+<OM<�<���;P��;T-�;3�;�7�;d�;1��;��;V�;ʆ�;*I�;(��;��;���;�)�;	��;1�;Jr;��b;��S;�zE;4�7;@�*;�H;`�;�|;���:�P�:F��:��:@A�:b��:o��:��:W�Z:�S1:��:u��99([9rX8c�3���Ѹ?��3�*�^28��b?��<F���R���j�f�������~ǹE�T���&��'=�;7S��g��r{�����Z珺&����$���N������.�UU��@Jĺ�>ʺ/�к�tغH��47�!������l��#����K&'���.��5�?(;�ձ?��"C�f�E��:G��YH�nII��cJ��L�N���Q��}V��[��b���h�Y6o���u���{��ۀ�ڞ��(E���ֈ��Z��Bˍ����vL��;L��?$���  �  O =��=��=�N=��=��=/=	�=�� =\ =6��<s�<Bt�<���<}��<�_�< �<���<���<Z��<�u�<xV�<!�<���<*Y�<#��<��<�`�<���<U��<�7�<:��<g��<c�<���<�6�<��<��<Id�<m��<�K�<���<uZ�<���<�c�<���<��<fF�<xP�<x>�<�<&��<o��<,��<���<���<�6�<?��<�;�<���<���<aW�<��<Ȓ�<"��<A7�<�A�<��<���<�j�<��<}_�<>��<�)�<P�<���<���<~�<�'�<*�<!'�<V%�<�(�<11�<�:�<�=�<0�<��<���<�R�<�°<��<�Z�<U��<W�<q;�<Ǵ�<'S�<f�<t
�<0 �<xT�<���<��<�>�<�}�<���<��<���<�a�<��<l͂<}�<�b|<e�w<`s<q�n<�wj<��e<]qa<M�\<�ZX<��S<ʄO<�CK<�G<��B<��><u�:<�6<�`1<Le,<[+'<��!<�C<��<�b<M1<�C<��<���;E��;�i�;��;���;�W�;���;`��;?��;NǼ;_��;q(�;�;Hߚ;%\�;��;��;�t;һe;cW;{�H;��:;�E-;!c ;�R;�3	;��:�[�:���:D��:s��:���:_y�:U�|:�jR:��':�O�9~˫9��F9���8lo��Nf޸�x(���L��M_���e��jf���g���o�&5���[������3йs.��3���%�O:���M�P�_�<�p��������x瑺�����!������s��+5��hĺ�_˺#�Һ��ںϋ�<:���x��������E�!��*�^�2�9��M?���C��G�� I�g]J�VK�%�K��^L�t�M�P��fS�8�W�H�\�8�b���h���n��t�N<z��e�A.������F"������T���펻9p��;ʓ�����  �  �=��=G�=�:=��= s=��=>k=�� =v8 =�<�<��<>�<F2�<�~�<n��<���<�j�<kP�<&D�<�8�<& �<Q��<	��<�-�<���<���<�I�<��<���<"O�<���<v2�<+��<��<q��<���<]>�<c��<���<�X�<��<wH�<u��<�>�<(��<���<=�<l�<��<���<���<�v�<?Z�<[�<���<���<�D�<D��<��<	T�<�<L��<S_�<���<S�<o�<���<��<{Y�<5��<�m�<d��<C\�<Y��<i�<>M�<�l�<xs�</i�<�U�<�A�<g3�<}+�<�'�<n �<��<�<��<�#�<D��<Mݭ<��<*M�<8��<wܢ<ZO�<n�<���<B��<Cė<��<HT�<_��<!�<^I�<�r�<\}�<�i�<8=�<� �<���<�|�<̄|<!!x<H�s<�so<�k<��f<�b<Do]<2�X<�0T<��O<KK<,G<~�B<��>< B:<��5<V1<6,<Լ&<vF!<|�<�"<Y�<tj<�q<�<9�;:�;��;:�;0��;gX�;W��;\��;ݾ�;q�;���;;T�;���;�h�;�h�;6��;�wv;��g;��Y;�@K;�=;�8/;��!;�=;s�	;f��:�"�:���:X_�:״:֧�:Yf�:e�u:cK:�l:���9Y��9�9�[�7�5���#�K�Z���{��|ͅ��ă��c����B]�������5����ٹ����/���u&�p�8��I� �Y�ʾh�&�w�J���팺�w��If���U���߳�d���`�ĺ��̺r�ԺBݺ�<纁󺓎 �R���r����3$�&>-���5�q�<���B�G��J���K���L�QM�l�M�� N�b\O��Q�y�T�*Y�m^�ͣc��Zi���n�+7t��!y�w�}��!��n��
߅�8}��B������ڐ�l}�����  �  =��=y}=�+=��=/b=��=�W=D� =�  =t�</��<���<���<C;�<I��<a�<.1�<��<�<A�<O��<���<�}�<
�<ԁ�<Y��<:7�<��<��<9[�<���<QU�<���<8N�<��<��<Le�<X��<�<Y^�<h��<�9�<S��<�#�<���<-��<���<���<5��<���<�s�<�?�<�<��<�=�<���<�<���<�Z�<�"�<��<ơ�<;�< ��<`��<���<���<p��<0K�<��<is�<M��<�y�<M��<C�<���<���<ݡ�<A��<6q�<dQ�<�6�<�$�<��<=
�<?�<B·<=t�<��<k�<b��<p�<��<R�<��<��<.��<�o�<g�<���<|˕<�#�<���<pݐ<a$�<�O�<?\�<�J�<y"�<��<M��<�x�<��|<^Ix<~	t<J�o<sk<Bg<�pb<��]<mY<�]T<��O<�HK<M�F<��B<7b><�:<��5<��0<+�+<8p&<�� <CU<�<�5<��
<2�<�E<��;�9�;q�;�c�;^��;̪�;w2�;-h�;�1�;���;�}�;%1�;|͢;�}�;�c�;,��;��;��w;*5i;6 [;��L;�>;�f0;��";��;в	;�O�:$%�:�v�:��:��:��:34�:�Dq:�F:'�:!6�9eވ9��8���Zt�ZAE��{����!ݒ��G��9莹�o���N��I������ ���u���4�2��1O'��`8�4�G�S0V� d�Jr�����߉�����f'��$¨����������ź��ͺ$ֺ�ߺ�3�C1��6����	�]��X8��%��/�@u7�V�>�
�D�KI�wL���M�t�N� �N� �N��WO��}P���R�A�U���Y�c�^��Id���i�Uo���s�Q�x�G�|�l~��)���k��u���ޚ��<���C����W�������  �  N=R�=5h=�=U�=eH=�=�S=�� =FB =r�<�l�<�|�<{��<��<�l�<q �<��<�s�<�B�<��<��<��<m/�<K��<�0�<���<���<�P�<���<��<�|�<���<XY�<���<*�<ވ�<���<�;�<a��<���<�\�<���<�/�<���<
��<�'�<�Q�<�c�<Ua�<9P�<�8�<�$�<�<?*�<^R�<��<>��<v�<��<��<d.�<���<t%�<�v�<���<c��<g��<�Z�<
�<Z��<%4�<���<d*�<��<���<M#�<xM�<[d�<l�<�i�<�b�<�Z�<\S�<EJ�<6;�<Y �<��<
��<O�<0ׯ<5J�<8��<i�<+u�<��</x�<u$�<A�<��<��<4�<jL�<���<���<��<u
�<a�<��<��<E��<͇�<1U�<9J|<��w<��s<pDo<��j<Xwf<��a<�r]<y�X<5aT<b�O<_�K< (G<E�B<s�><�:<��5<!�0<��+<��&<��!<��<�C<�<5<�K<��<��;��;E��;Bm�;ل�;1��;���;۲�;t]�;E��;��;�٭;���;���;˶�;��;�a�;c~;�o;r^a;�\S;P�E;@8;z+;;�;R ;o;��:�'�:�c�:���:{�:�:O�:pzi:Z�@:Y:X8�9ek�98E9�%�8<�6��h���ҸzZ
��0!�ZA3���E�y`]��s}�^��I����ι���
���r/��?@��P��"a���q��d��]m���哺�����w������p��ntúyV̺hպߺ̴麙������������}1���!���)��1�\�7��i=�B�?�E��/H�$ J�*�K��M�ձN�t�P���S��V�[���_���d��j��So�Pht��Oy�~��e���̃�GJ���䈻�����S�����j����G���  �  �=�=�j=�=ʵ=>L=R�=sX=� =)H =Z�<�z�<d��<���<w
�<�|�<��<G��<��<N�<�<J��<X��<�6�<���<�6�<;��<}��<�Q�<��<P�<�u�<���<uN�<۸�<�<g}�<���<�3�<��<���<K\�<���<�3�<���<V��<./�<�Y�<~l�<#k�<"[�<E�<(2�<�+�<:�<�b�<$��<$
�<τ�<N�<_��<Q9�<Q��<7.�<�~�<���<}��<O��<�^�<��<ѥ�<"1�<���<="�<�<��<��<A�<�X�<b�<b�<�]�<ZX�<PS�<{L�< ?�<e%�<��<��<�V�<�߯<T�<Q��<��<"��<���<;��<�4�<��<��<���<�#�<�X�<���<fː<���<r�<��<�	�<��<���<t��<_T�<NC|<��w<��s<a/o<)�j<�^f<��a<*]]<��X< TT<A�O<�}K<	*G<��B<��><N&:<+�5<<�0<�,<�'<��!<��<w^<6<�5<�l<_�<�G�;aM�;��;��;´�;h��;S��;���;^}�;�ܽ;8��;��;x˥;Q��;���;��;(H�;L�};�>o;�a;��R;@:E;��7;��*;,�;��;�;x��:wj�:��:�6�:�|�:�D�:���:��j:�@B:�:���9&!�9��L9l{�8ot7��H���ø�n�#���-���@��X��ly��.�����{�̹���9l
�?�AY/�<�@���Q�\]b�!s��$��1+�� ���n<���觺�e��`����lú+̺�!պ�޺eK��3���I����=������!!��')��0�h?7���<� �A�PE�y�G��I��EK�\�L��eN�7�P��DS��V���Z���_��d�nj��Zo�5�t��y�vU~�����Y����z���������zv��'���œ�8L���  �  ;
=&�=q=�=F�=�V=4�=�e=�� =Y =P��<��<���<��<M:�<���<6<�<`��<��<�n�<.9�<"��<z��<�K�<p��<$F�<6��<���<�R�<p��<	�<%a�<D��<�-�<6��<���<[�<��<��<O��<���<�Z�<E��<�=�<���<���<�B�<�o�<��<���<?z�<h�<vY�<�V�<h�<$��<���<R8�<���<�8�<���<rX�<���<�F�<��<þ�<:��<֥�<�g�<��<���<�'�<���<�	�<�f�<���<���<��<6�<bD�<�J�<�M�<YP�<=R�<Q�<9I�<P3�<�	�<Tȴ<�l�<���<�o�<�٪<�?�<R��<�%�<޶�<�d�<2�<G�<?)�<�J�<.{�<p��<��<.�<�(�<\,�<!�<i��<7Ƅ<���<UQ�<-.|<'�w<�Ws<��n<��j<�f<V�a<�]< �X<g,T<��O<�sK<�-G<��B<У><�E:<�5<�1<�>,<]:'<�"<o�<�<�<c�<��< G<E <U�;�s�;`<�;�=�;�T�;~\�;<8�;���;*,�;�?�;�"�;��;���;͟�;��;���;��|;vBn;��_;t�Q;�/D;��6;�%*;?
;	�;I;��:S�:���:ZU�:p��:⫞:@�:7n:0F:t:��9c�95$d9tM�8y�8�׷�w���޸'	����>�2��lL��Ln��0�������"ɹ�<�U�	�:�m\0�#�B�ǪT�3f�kKw�th��i��S���`���p@���G��h����eúx�˺�iԺ�ݺ�(躨��t� �n����i�����,�'��:/���5��g;�6@�%�C�iF���H�Q4J���K���M���O��R�\"V�@`Z�i7_�yd���i�sto�_�t��z����������d������@?��tގ�Is����C\���  �  �
=�=iy=�'=C�=�e=;�=y=6� =�r =D��<���<���<�3�<��<���<S��<�&�<S��<���<:d�<� �<���<�h�<���<	[�<���<��<�Q�<���<���<D>�<��<���<u[�<"��<�#�<؉�<��<�c�<���<�T�<|��<!J�<]��<��<^�<���<���<��<Ũ�<`��<���<a��<k��<H��<�!�<��<���<cu�<.��<��<�<�i�<ò�<E��<���<���<es�<S�</��<��<G��<���<U4�< {�<߳�<���<���<��<9$�<�2�<�@�<�M�<VV�<�U�<�E�<� �<�<���<��<���<�	�<�v�<�<�i�<:��<5��</|�<Af�<'k�< ��<ͯ�<x��<�<�3�<�G�<�G�<R2�<�	�<ф<���<�I�<�|<ׁw<�s<W�n<Cj<�e<\'a<=�\<�GX<!�S<��O<�^K<<-G<��B<�><vo:<V�5<,S1<ʁ,<T�'<�n"</F< <�<�<�b	<��<� <� �;y�;�&�;;�;/
�;��;���;�R�;a��;���;sh�;�;N��;x�;4\�;Zu�;�{;ݦl;�,^;�P;�B;�i5;��(;u1;!/;�;j�:H��:r��:l��:Ԃ�:}��:?V�:�Xs:�L:��%:�]:*��9��9�r!9�"�8Z�7F�)�mҡ��ܸR3��5��c:��m^�A��j���yPĹ��鹍	����O2��EF��{Y��l��+~�����	�����pࢺ����Fѳ�(Ȼ��ú�P˺�Ӻ={ܺ�溣#�������$\��L��?���%�-�+�3�<9�h�=��oA��]D���F���H�M`J�^TL�ưN��Q�
OU�_�Y���^��#d��i���o��tu�H
{��7���ւ�i��4�����������������@F��U����  �  �=A�=��=D2=��=�u=�='�=Z=p� =b =r6�<VX�<F��<'��<~Q�<m��<�u�<�#�<��<���<UK�<���<N��<&�<�n�<���<��<�J�<t��<6��<7�<[�<���<��<]p�<���<G�<��<�:�<]��<TH�<��<tS�<d��<-�<xz�<D��<��<���< ��<=��<'��<���<�	�<t:�<M��<���<G�<}��<�@�<���<�1�<���<���<���<���<e��<�{�<��<n��<K��<�V�<%��<j��<m-�<�a�<c��<���<���<?��<;�<�'�<KB�<pV�<�^�<
V�<7�<���<Ϭ�<�C�<�ȭ<�B�<���<�5�<"��<[�<�<5ڜ<���<���<mϖ<��<��<Q=�<[�<ni�<)d�<LI�<�<�ل<Z��<n:�<��{<%)w<�r<]�m<zi<��d<@�`<�$\<��W<�S<�YO<9K<�!G<XC<��><`�:<�*6<C�1<��,<(�'<.�"<n�<��<ѱ<��<|!
<�<�W</��;���;�G�;]�;���;���;Ib�;��;�;���;��;K0�;۪�;�0�;bی;U��;&�y;�zj;F�[;E�M;+8@;c3;�J';T�;Ei;��;}�:���:^�:�_�:Y[�:֢:�ݏ:�Jy:S:��-:
�
:	��99^�P9��84[8�u��q�+�Mޙ���Ӹ/W��3&�eHM�5~�<͜��ۿ�7b繵	��+��l5�72K��.`��Bt�C���
���땺Q����Ԧ�%������$��;ĺ�˺��ҺSGۺ���A�7���.e�����x���#��c*�/�0�66�x�:���>��A��fD��F��H��J��M���P��tT�7�X�0^���c�#�i�<1p�Ibv�kl|�N��wꃻ����2��D���%���w��=����Ô��Ŗ��  �  �=O�=s�=�9=�=(�=�=}�=�+=�� =9: =ݏ�<^��<e��<	O�<���<�9�<z��<�n�<f�<I��<�s�<��<��<��<"|�<#��<��<�:�<�h�<֘�<	��<��<�Y�<ׯ�<0�<�}�<���<Ex�<?�<��<�1�<���<�T�<T��<�=�<F��<B��<���<��<��<h#�<�1�<�I�<o�<X��<]��<o@�<s��<��<U��<���<�_�<��<���<Y
�<���<���<|{�<��<�w�<`��<��<ha�<��<���<��<+�<UU�<X�<s��<2��<��<�,�<lM�<`�<7_�<�F�<��<�ɲ<�h�<���<�}�<v�<e��<h�<*¡<�x�<�C�<e$�<�<z�<]3�<�N�<|j�<N�<u��<{�<�Y�<j#�<�ل<���<P!�<�z{<��v<��q<;Vm<˿h<�<d<��_<;w[<�7W<�S< O<��J<�G<��B<�><��:<�Q6<!�1<-<�3(<�A#<�E<�M<)g<<�<��
<z|<�-<��;5(�;ۀ�;��;���;�b�;$��;
M�;Vf�;B8�;�ɮ;H+�;?u�;K;�,�;Ỹ;�ew;;�g;=�X;��J;!u=;��0;7%;�];�N;z�;u�:\��:���:��:*޶:���:8�:�&:cLZ:��6:�:I�9�>�9-�9�l19O�8<8<���&������yݸZd��Z>�_7r��o��d'��׽�)
���!�!�9�V�Q�(�h�ZH~�Z��p蒺ZЛ����ޭ����������'���(ź�v˺3tҺ�ں���P�������(��D�ː����a� �tb'�8d-���2�+y7�*�;�8�>���A��D��G��I�iL�?�O���S�Z�X���]���c��Yj���p�,�w�]4~��>��:���
��r���*��My�����(����n��m2���  �  ��=ο=}�=J;=��=��=m$=�=�C=�� =�` =7��<� �< g�<���<%�<��<�#�<���<U�<��<���<*�<��<"�<~�<`��<I��<)�<?�<�_�<���<���<���<�F�<��<��<��<")�<L��<�i�<~�<@��<K�<���<EC�<C��<���<��<�2�<!M�<
f�<��<ϧ�< ��<��<X�<��<��<e�<���<�,�<��<���<i�<,�<	�<���< p�<���<tT�<S��<���<�<O<�<tf�<ܐ�<���<���<�"�<\�<c��<���<�<9�<�U�<�\�<=K�< �<�ܲ<셰<
!�<´�<�G�<'ߦ<��<`,�<�<:��<s��<�u�<�n�<,t�<g��<���<随<���<��<f_�<�!�<�΄<�k�<x�<�{<
0v<Yq<��l<L�g<fec<��^<��Z<�V<��R<�N<:�J<��F<�B<��><W�:<�b6<��1<�>-<�y(<]�#<;�<��<�<�k<f�<�^<h
<ܱ�;��;���;?�;{�;!��;z\�;���;j��;�M�;8��;���;b�;�(�;)U�;#��;��t;��d;��U;t�G;r[:;_.;��";-q;��;��;���:�O�:/��:"��:���:G�:��:��:W�`:&!?:FQ:��:�s�9��9Z�h9t�9N �81!8�1綐�F��ȴ�����&4���k�Pؖ�kF����蹴f���%�ѳ?�}pY�mBr��ք����i����d��pD���3���K��i��� ���+�ƺ�̺��Һ�oں<e�/��s���9,�j�	�������� ��P$�**��O/�]4�R8�<�q|?�ÎB�xE��iH�ʘK��8O�tS�_bX�^��Md��k�a"r��Gy��'��懃����������Y���Ɏ������쒻p���dD��˗��  �  p�=��=Hz=�6=v�=��=7+=��=RW=� =� =q =y��<"��<�'�<���<4��<�u�<y��<��<��<��<`5�<���<��<s�<B��<���<���<f�<��<7�<�[�<���<���<�8�<���<w7�<���<T~�<L1�<���<<��<h5�<���<�;�<���<���<�!�<@P�<�x�<m��<���<� �<x:�<�z�<e��<"�<]]�<���<9�<NY�<���<���<��<K�<��<%��<pX�<���<�'�<g�<��<`��<���<���<]�<�K�<���<���<4�<BR�<���<��<��<?�<�M�<�B�<��<R�<e��<�@�<��<���<�-�<�ۤ<���<#Q�<�<��<�̙<���<���<z��<���<=��<���<K��<�W�<+�<f��<K�<R�<d�z<o�u<ȧp<��k<�g<��b<, ^<�Y<��U<��Q<�N<�KJ<q�F<�B<6�><>�:<2Z6<m�1<�X-<y�(<y�#<�/<\v<��<�0<�<�8<�<8�;#��;���;���;�;"^�;
��;ݱ�;ᒿ;�/�;J��;���;7��;�l�;�_�;l��;��q;��a;oR;Q7D;(7;"+;�: ;�L;b.;m�;h�:��:q�:���:z��:댦:�1�:���:K�f:�F:��(:\:2y�9-�9Oَ9�5Q9�Y9Y�8>�7G�ַ����k����0�
�k�1���@�����!��*���F�^b���|��܊�5D���k��@���ð�����V�����%ź�^ɺ�9κ�Ժ*ۺ$�������������� ?�D��\��2h!���&���+�%�0��D5��j9��?=���@� 3D���G��"K�~O�/�S���X���^�)
e�`l��s��#{�rP���脻EE���V��3��={��w���?S���ڕ��8��T����  �  ^�=ˢ=�l=L,=O�=E�=s,=��=Qe=�=K� =vD =��<:,�<F��<���<�N�<���<�2�< ��<�2�<s��<�5�<���<��<=]�<M��<z��<���<W��<a��<���<W �<4,�<�o�<���<=F�<���<�~�<�5�< ��<ݴ�<,m�<d�<U��<W)�<z��<���<�'�<�b�<��<Z��<J�<�N�<ݒ�<��<��<1f�<F��<���<68�<{�<���<���<-�<>�<=��<��<�7�<��<��<�(�<J�<�`�<�u�<'��<ү�<w��<w�<H`�<&��<�	�<�`�<���<��<�<�3�<D/�<R�<��<���<�U�<N�<���<r�<-�<��<9��<�w�<�D�<��<���<0ܕ<}ʓ<Ľ�<_��<�<z�<nE�<d��<���<�"�<�:<�z<	u<��o<)	k<Cf<n�a<�K]<�Y<�U<"IQ<	�M<��I<b,F<�fB<ɀ><Ts:<&;6<��1<0\-<8�(<�'$<�<I�<Aa<+�<ih<-�<G�<�H <l�;��;8��;���;��;���;��;�a�;��;,"�;��;��;қ�;^�;aQ�;�3o;�^;�5O;_�@;@�3;88(;ۤ;_;^];�4;y��:�?�:f��:ۉ�:��:n^�:���:�6�:9�j:"�L:w�0:0�:��9Q��9%��9�~9�549��8�	D8����u��%n��1�\Iq�񜹯�ƹʦ�����C�0�Z�M��k�x����Ő�W������U᯺��+ּ�Yh���*źf�ȺE5̺(|к��պA�ܺW���I�����u3�f�f�,��8u�q���$��)��-��2��7�U;��b?��EC��G��K��>O���S�FGY�(R_�\f�9fm�g)u��}��~��'G���ˉ�k���ؿ���������������F:��~Y���  �  z�==�=4]==��=$�=�)=2�=?n=�=�� =tb =� =Ey�<0��<�3�<��<���<^�<���<~A�<���<�-�<��<���<�A�<�u�<���<2��<���<��<���< ��<���<��<�n�<;��<��<b1�<���<��<߃�<�C�<1��<���<��<�}�<���<4%�<�k�<h��<5��<}A�<_��<���<'�<�m�<���<���<�&�<	^�<R��<���<���<��<y��<^��<���<��<�{�<]��<��<e�<��<<�<U/�<�M�<�{�<���<�	�<�d�<���<�&�<�<�Ǽ<���<�<��<,��<�ղ<<ga�<�!�<��<ʨ�<�o�<�7�<���<�Ş<���<�V�<
'�<���<ߓ<,ő<ܬ�<ˏ�<g�<�,�<a܆<u�<C��<��~<ڧy<xt<iXo<Yj<��e<+�`<m�\<�jX<�{T<�P<UM<tI<��E<=B<�>><�;:<>6<z�1<dO-<V�(<wK$<#�<N<l�<�n<<4�	<�7<�� <��;�u�;�;���;���;���;ji�;��;Ă�;���;���;H;�;�Α;5j�;�l~;S�l;��[;WL;">;/'1;f�%;eJ; 
;n�	;�;�A�:�%�:'��:t�:0��:���:#��:'Ӆ:��m:S�Q:�g7:� :o:m�9�P�9Ӕ�9��T9�k
9���8��/6��m����z�6��Zz�b���͹aI��Y��I�6�yU��Ys��^������e������Ƶ������
º�
ƺ2ɺn̺�Ϻ��Һx�׺OT޺�,溳Tﺟ���3+�����1����������Ѩ!�N�&�r+��T0�;$5���9��T>���B���F��+K�*�O���T�>Z�J`��2g�A�n�
�v���~�q��������)��l��C<������x������*��/���(���  �  E�=T=dN=/=�=�z=�$=��=1s=�=� =<x =�( =}��<��<l�<<��<-�<|�<���<�H�<��<�"�<N��<��<'�<W�<4q�<�x�<
s�<�h�<�c�<@l�<���<���<1$�<���<�=�<7��<x��<���<�Y�<��<���<q�<!��<ii�<���<w�<9n�<��<Z�<f�<��<��<�`�<��<��<%�<<L�<x�<���<���<T��<v��<���<���<,f�<4��<�U�<��<3��<���<���<��<���<n �<�.�<�p�<���<&�<q��<��<{T�<��<�ٺ<���<���<��<�ǲ<���<#f�<:2�< �<:Ч<���<�n�<m9�<J��<���<��<�I�<g�<!�<�Ƒ<N��<��<�R�<*�<ￆ<OT�<�ҁ<�~<-Dy<\t<��n<f�i<��d<V`<v�[<��W<��S<jBP<b�L<bI<N�E<A�A<i><:<`�5<c�1<�;-<��(<\_$<a�<>�<?4<��<?{<�
<P�<{?<ү�;��;�e�;���;S��;�q�;�+�;#þ;� �;{8�;�
�;ܤ�;- �;���;�|;��j;��Y;�J;�;;J�.;�#;�e;�[;$;}u ;u	�:�1�:��:ܛ�:�Ǵ:�ܤ:@*�:�:wyo:p�T:�<:F�$:��:��9 ��9�L�95�l9Rq9WZ�8�0$7�!f��p����=�������Թ�"�,���<���Z��+z�J5���Q���禺㪱�_k���/��R1ƺk�ɺ�̺M�κ8�Ѻ�#պ��ٺkພ�红z��A���H�9�� ��H���t��0�a��_�$�E�)���.��3���8��=�aQB��F�pK�
(P��=U��Z��3a��=h��o�5x�*F���y��5���<?������lg��P���E���c����������ٚ��  �  �=�s=�C=�=��=�t=� =��=gu=�"=�� =i� =�8 =���<>5�<֎�<���<8�<V��<���<�K�<n��<r�<�z�<6��<��<pA�<Y�<�]�<{T�<^F�<�<�<�A�<�]�<:��<\��<�r�<��<���<1��<Uj�<>=�<��<��<�\�<��<TZ�<U��<E�<n�<���<��<�{�<1��<�2�<̄�<���<��<�8�<�b�<
��<ק�<��<6��<	��<>��<^��<Q�<���<y;�<y�<��<F��<&��<��<���<���<v��<A�<���<L��<�i�<�տ<�7�<.��<Hº<��<H�<�۴<��<U��<Vg�<�:�<|�<��<\��<7��<�]�<�"�<>�<~��<�^�<�#�<��<�ő<���<nu�<�C�<�<���<f=�<+��<EE~<=y<Իs<��n<ysi<�d<_�_<��[<1�W<�S<m�O<�cL<Q�H<LE<��A<��=<��9<�5<R�1<D+-<�(<Bh$<� <�<j<<{�<�a
<�<�<��;�E�;l��;S�;��;WS�;���;���;2ٵ;y�;��;�=�;Ȫ�;��;�u{;�hi;aX;=�H;�P:;��-;R,";�);�@;�);�/�:���:,��:���:���:�߳:�0�:�Δ:��:_p:!�V:�>:�s(:�:��9��9���9�M{9��(9Ͳ8t�a7v�d�������B�6���V`��c�ٹ�����!���?���^�u�~�𵎺S��Щ�����oe���ĺ3�Ⱥ�;̺��κ��к�SӺ?�ֺ=ۺ{>��躤X������j�Wq�[�	�Q��/?������#��(��-���2��8�99=��'B�
�F�E�K���P�;�U��u[�O�a�E�h�2�p�y�aʀ����q(����oM���&��ow��dD��B����������P���  �  i�=Jo=@=T=�=?r=/=4�=
v=�$=� =͉ =�= =u��<bA�<t��<S��<e@�<1��<6��<|L�<���<��<�u�<��<��<�9�<PP�<�S�<�I�<]:�<a/�<(3�<ON�<���<���<�b�<��<���<|��<	_�<3�<m��<��<eU�<���<�T�<��<��<�m�<���<�#�<��<���<�=�<���<���<��<�B�<j�<���<��<���<���<���<���<���<wI�<L��<2�<o�<t��<D��<���<e��<��<��<���<�0�<���<#��<B]�<$ʿ<M-�<�~�<Ṻ<V۸<��<[ִ<Ḳ<��<�g�<�=�<��<��<`ȥ<���<�i�<�.�<�<���<|e�<%(�<��<ő<���<
q�<'>�<���<-��<.5�<��<�0~<(�x<��s<in<�Ti<>td<O�_<�x[<�aW<ʆS<��O<�KL<��H<�8E<&�A<,�=<~�9<�5<�w1<�$-<��(<�j$<� <��<�{<�/<��<�z
<<�<<�;_�;���;b�;k��;�F�;���;�n�;Ծ�;�ɬ;���;��;���;`�;A{;��h;��W;!H;��9;�-;��!;ͻ;��;�;��:���:]T�:Nm�:� �:닳:J�:���:�	�:�p:HAW:��?:̥):Cn::	�9��9���9��9$�,9�߷8jau7#�d��H��pE����������۹�����"���@��Z`����^���]���SЪ�
����i��xź��ɺyͺirϺF�Ѻ�ӺK8׺�ۺ���麗��{��/z�km��B�p��s����z��4#��*(�rU-���2�}�7�=�?B�'�F���K�x�P���U�ī[��b�;i�:q�Yy������B���a��C/��5���5h��_�������٘�mܙ������y���  �  �=�s=�C=�=��=�t=� =��=gu=�"=�� =i� =�8 =���<>5�<֎�<���<8�<V��<���<�K�<n��<r�<�z�<6��<��<pA�<Y�<�]�<{T�<^F�<�<�<�A�<�]�<:��<\��<�r�<��<���<1��<Uj�<>=�<��<��<�\�<��<TZ�<U��<E�<n�<���<��<�{�<1��<�2�<̄�<���<��<�8�<�b�<
��<ק�<��<6��<	��<>��<^��<Q�<���<y;�<�y�<��<F��<&��<��<���<���<v��<A�<���<M��<�i�<�տ<�7�</��<Iº<��<I�<�۴<��<V��<Vg�<�:�<|�<��<]��<8��<�]�<�"�<>�<}��<�^�<�#�<��<�ő<���<mu�<�C�<�<���<e=�<*��<CE~<;y<ӻs<��n<ysi<�d<_�_<��[<1�W<�S<n�O<�cL<S�H<LE<��A<��=<��9<�5<T�1<F+-<�(<Dh$<� <�<j<<{�<�a
<�<�<��;�E�;h��;O�;��;RS�;���;|��;-ٵ;t�;��;�=�;Ī�;��;�u{;�hi;	aX;8�H;�P:;��-;O,";�);�@;�);�/�:���:*��:���:���:�߳:�0�:�Δ:��:_p:!�V:�>:�s(:�:��9��9���9�M{9��(9Ͳ8u�a7v�d�������B�6���V`��c�ٹ�����!���?���^�u�~�𵎺S��Щ�����oe���ĺ3�Ⱥ�;̺��κ��к�SӺ?�ֺ=ۺ{>��躤X������j�Wq�[�	�Q��/?������#��(��-���2��8�99=��'B�
�F�E�K���P�;�U��u[�O�a�E�h�2�p�y�aʀ����q(����oM���&��ow��dD��B����������P���  �  E�=T=dN=/=�=�z=�$=��=1s=�=� =<x =�( =}��<��<l�<<��<-�<|�<���<�H�<��<�"�<N��<��<'�<W�<4q�<�x�<
s�<�h�<�c�<@l�<���<���<1$�<���<�=�<7��<x��<���<�Y�<��<���<q�<!��<ii�<���<w�<9n�<��<Z�<f�<��<��<�`�<��<��<%�<<L�<x�<���<���<U��<v��<���<���<,f�<4��<�U�<��<4��<���<���<��<���<o �<�.�<�p�<���<&�<s��<��<~T�<"��<�ٺ<���<���<��<�ǲ<���<$f�<<2�< �<;Ч<���<�n�<m9�<I��<���<��<�I�<f�<�<�Ƒ<L��<��<�R�<(�<�<MT�<�ҁ<�~<*Dy<Yt<��n<d�i<��d<V`<w�[<��W<��S<mBP<e�L<eI<Q�E<E�A<m><�:<e�5<g�1<�;-<��(<__$<d�<A�<A4<��<@{<�
<O�<z?<ί�;z��;�e�;���;K��;�q�;�+�;þ;� �;r8�;�
�;Ӥ�;% �;���;�|;v�j;��Y;�J;��;;C�.;��#;�e;�[;$;zu ;p	�:�1�:��:ڛ�:�Ǵ:�ܤ:@*�:�:vyo:o�T:�<:F�$:��:��9 ��9�L�95�l9Rq9XZ�8�0$7�!f��p����=�������Թ�"�,���<���Z��+z�J5���Q���禺㪱�_k���/��R1ƺk�ɺ�̺M�κ8�Ѻ�#պ��ٺkພ�红z��A���H�9�� ��H���t��0�a��_�$�E�)���.��3���8��=�aQB��F�pK�
(P��=U��Z��3a��=h��o�5x�*F���y��5���<?������lg��P���E���c����������ٚ��  �  z�==�=4]==��=$�=�)=2�=?n=�=�� =tb =� =Ey�<0��<�3�<��<���<^�<���<~A�<���<�-�<��<���<�A�<�u�<���<2��<���<��<���< ��<���<��<�n�<;��<��<b1�<���<��<߃�<�C�<1��<���<��<�}�<���<4%�<�k�<h��<5��<}A�<_��<���<'�<�m�<���<���<�&�<	^�<S��<���<���<��<y��<^��<���<��<�{�<]��<��<f�<��<=�<V/�<�M�<�{�<���<�	�<�d�<��<�&�<�<�Ǽ<���<�<��</��<�ղ<�<ja�< "�< �<̨�<�o�<�7�<���<�Ş<���<�V�<'�<���<ߓ<)ő<٬�<ȏ�<g�<�,�<^܆<u�<@��<��~<էy<xt<gXo<Yj<��e<+�`<n�\<�jX<�{T<�P<YM<tI<��E<CB<�>><�;:<D6<��1<jO-<[�(<|K$<(�<"N<n�<�n<<4�	<�7<�� <��;�u�;�;���;}��;���;]i�;s�;���;驭;u��;;;�;�Α;*j�;�l~;A�l;��[;�VL;>;$'1;]�%;]J;
;i�	;�;�A�:�%�:#��:q�:.��:�:"��:&Ӆ:��m:S�Q:�g7:� :o:m�9�P�9Ӕ�9��T9�k
9���8��/6��m����z�6��Zz�b���͹aI��Y��I�6�yU��Ys��^������e������Ƶ������
º�
ƺ2ɺn̺�Ϻ��Һx�׺OT޺�,溳Tﺟ���3+�����1����������Ѩ!�N�&�r+��T0�;$5���9��T>���B���F��+K�*�O���T�>Z�J`��2g�A�n�
�v���~�q��������)��l��C<������x������*��/���(���  �  ^�=ˢ=�l=L,=O�=E�=s,=��=Qe=�=K� =vD =��<:,�<F��<���<�N�<���<�2�< ��<�2�<s��<�5�<���<��<=]�<M��<z��<���<W��<a��<���<W �<4,�<�o�<���<=F�<���<�~�<�5�< ��<ݴ�<,m�<d�<U��<W)�<z��<���<�'�<�b�<��<Z��<J�<�N�<ݒ�<��<��<1f�<F��<���<68�<{�<���<���<-�<>�<=��<��<�7�<��<��<�(�<J�<�`�<�u�<)��<ԯ�<y��<y�<K`�<)��<�	�<�`�<���<��<�<�3�<H/�<U�<��<��<�U�<Q�<���<r�<-�<��<9��<�w�<�D�<��<���<.ܕ<zʓ<���<\��<<z�<jE�<`��<���<�"�<�:<�z<u<��o<'	k<Cf<n�a<�K]<�Y<�U<&IQ<�M<�I<i,F<�fB<Ѐ><[s:<.;6<��1<7\-<>�(<�'$<�<M�<Ea<-�<jh<-�<F�<�H <f�;ٻ�;.��;��;��;��;��;�a�;��;"�;��;��;ě�;^�;TQ�;�3o;��^;�5O;P�@;3�3;-8(;Ҥ;W;X];�4;q��:�?�:b��:؉�:��:l^�:���:�6�:8�j:!�L:v�0:0�: ��9Q��9%��9�~9�549��8�	D8����u��$n��1�\Iq�񜹯�ƹʦ�����C�0�Z�M��k�x����Ő�W������U᯺��+ּ�Yh���*źf�ȺE5̺(|к��պA�ܺW���I�����u3�f�f�,��8u�q���$��)��-��2��7�U;��b?��EC��G��K��>O���S�FGY�(R_�\f�9fm�g)u��}��~��'G���ˉ�k���ؿ���������������F:��~Y���  �  p�=��=Hz=�6=v�=��=7+=��=RW=� =� =q =y��<"��<�'�<���<4��<�u�<y��<��<��<��<`5�<���<��<s�<B��<���<���<f�<��<7�<�[�<���<���<�8�<���<w7�<���<T~�<L1�<���<<��<h5�<���<�;�<���<���<�!�<@P�<�x�<m��<���<� �<x:�<�z�<e��<"�<]]�<���<9�<NY�<���<���<��<K�<��<&��<pX�<���<�'�<g�<��<a��<���<���<_�<�K�<���<���<7�<FR�<���<��<��<?�<�M�<�B�<��<V�<h��<�@�<��<���<�-�<�ۤ< ��<#Q�<�<��<�̙<���<}��<w��<���<9��<���<G��<�W�<&�<b��<K�<K�<^�z<j�u<ħp<��k<�g<��b<- ^<!�Y<��U<��Q<�N<�KJ<x�F<!�B<?�><F�:<;Z6<u�1<�X-<��(<��#<�/<av<��<�0<�<�8<�<8�;��;���;���;r�;^�;���;˱�;ϒ�;�/�;8��;���;&��;}l�;�_�;^��;��q;�a;�nR;@7D;7;�!+;�: ;�L;[.;h�;`�:��:m�:���:w��:錦:�1�:���:I�f:�F:��(:[:1y�9-�9Oَ9�5Q9�Y9Y�8?�7F�ַ����k����0�
�k�1���@�����!��*���F�^b���|��܊�5D���k��@���ð�����V�����%ź�^ɺ�9κ�Ժ*ۺ$�������������� ?�D��\��2h!���&���+�%�0��D5��j9��?=���@� 3D���G��"K�~O�/�S���X���^�)
e�`l��s��#{�rP���脻EE���V��3��={��w���?S���ڕ��8��T����  �  ��=ο=}�=J;=��=��=m$=�=�C=�� =�` =7��<� �< g�<���<%�<��<�#�<���<U�<��<���<*�<��<"�<~�<`��<I��<)�<?�<�_�<���<���<���<�F�<��<��<��<")�<L��<�i�<~�<@��<K�<���<EC�<C��<���<��<�2�<!M�<
f�<��<ϧ�< ��<��<X�<��<��<e�<���<�,�<��<���<j�<,�<	�<���< p�<���<tT�<T��<���<�<P<�<vf�<ސ�<���<���<�"�< \�<g��<���<�<9�<�U�<�\�<BK�< �<�ܲ<���<!�<Ŵ�<�G�<*ߦ<��<a,�<�<:��<q��<�u�<�n�<)t�<d��<���<嚏<���<��<a_�<�!�<�΄<�k�<q�<�{<0v<
Yq<�l<K�g<fec<��^<��Z<�V<��R<�N<A�J<��F<�B<��><`�:<�b6<��1<�>-<�y(<d�#<A�<��<�<�k<h�<�^<f
<ױ�;��;��;3�;{�;��;i\�;���;W��;�M�;%��;���;P�;�(�;U�;��;��t;��d;��U;b�G;c[:;R.;��";%q;��;��;���:�O�:*��:��:���:E�:��:��:V�`:%!?:EQ:�:�s�9��9Z�h9t�9N �82!8�1綏�F��ȴ�����&4���k�Pؖ�jF����蹴f���%�ѳ?�}pY�mBr��ք����i����d��pD���3���K��i��� ���+�ƺ�̺��Һ�oں<e�/��s���9,�j�	�������� ��P$�**��O/�]4�R8�<�q|?�ÎB�xE��iH�ʘK��8O�tS�_bX�^��Md��k�a"r��Gy��'��懃����������Y���Ɏ������쒻p���dD��˗��  �  �=O�=s�=�9=�=(�=�=}�=�+=�� =9: =ݏ�<^��<e��<	O�<���<�9�<z��<�n�<f�<I��<�s�<��<��<��<"|�<#��<��<�:�<�h�<֘�<	��<��<�Y�<ׯ�<0�<�}�<���<Ex�<?�<��<�1�<���<�T�<T��<�=�<F��<B��<���<��<��<h#�<�1�<�I�<o�<X��<]��<o@�<s��<��<U��<���<�_�<��<���<Y
�<���<���<|{�<��<�w�<a��<��<ia�<���<���<��<+�<XU�<[�<w��<6��<��<�,�<pM�<`�<<_�<�F�<��<�ɲ<�h�<���<�}�<y�<g��<j�<+¡<�x�<�C�<d$�<
�<x�<Z3�<�N�<xj�<K�<q��<{�<�Y�<f#�<�ل<���<M!�<�z{<�v<��q<8Vm<ʿh<�<d<��_<=w[<�7W<�S< O<��J<�G<��B<�><ű:<�Q6<*�1<-<�3(<�A#<�E<�M<-g<?�<��
<z|<�-<��;.(�;Ҁ�;�;~��;�b�;��;�L�;Df�;/8�;�ɮ;6+�;.u�;:;�,�;K̃;ew;$�g;)�X;t�J;u=;��0;�6%;�];�N;u�;m�:V��:���:��:(޶:���:8�:�&:bLZ:��6:�:H�9�>�9,�9�l19O�8<85���&������yݸZd��Z>�_7r��o��d'��׽�)
���!�!�9�V�Q�(�h�ZH~�Z��p蒺ZЛ����ޭ����������'���(ź�v˺3tҺ�ں���P�������(��D�ː����a� �tb'�8d-���2�+y7�*�;�8�>���A��D��G��I�iL�?�O���S�Z�X���]���c��Yj���p�,�w�]4~��>��:���
��r���*��My�����(����n��m2���  �  �=A�=��=D2=��=�u=�='�=Z=p� =b =r6�<VX�<F��<'��<~Q�<m��<�u�<�#�<��<���<UK�<���<N��<&�<�n�<���<��<�J�<t��<6��<7�<[�<���<��<]p�<���<G�<��<�:�<]��<TH�<��<tS�<d��<-�<xz�<D��<��<���< ��<=��<'��<���<�	�<t:�<M��<���<G�<}��<�@�<���<�1�<���<���<���<���<e��<�{�<��<o��<L��<�V�<&��<k��<o-�<�a�<e��<���<���<B��<?�<�'�<OB�<tV�<�^�<V�<7�<���<Ӭ�<�C�<�ȭ<�B�<���<�5�<#��<[�<�<5ڜ<���<���<kϖ<��<��<N=�<	[�<ji�<%d�<HI�< �<�ل<W��<k:�<��{< )w<��r<Z�m<zi<��d<A�`<�$\<��W<�S<�YO<9K<�!G<_C<��><h�:<�*6<J�1<��,</�'<4�"<s�<��<Ա<��<}!
<�<�W<*��;���;�G�;R�;���;z��;:b�;��;�;���; ��;;0�;˪�;�0�;Tی;H��;�y;ozj;4�[;5�M;8@;�b3;�J';L�;?i;��;}�:���:Z�:�_�:W[�: ֢:�ݏ:�Jy:S:��-:	�
:��99]�P9��84[8v��q�+�Lޙ���Ӹ/W��3&�eHM�4~�<͜��ۿ�7b繵	��+��l5�72K��.`��Bt�C���
���땺Q����Ԧ�%������$��;ĺ�˺��ҺSGۺ���A�7���.e�����x���#��c*�/�0�66�x�:���>��A��fD��F��H��J��M���P��tT�7�X�0^���c�#�i�<1p�Ibv�kl|�N��wꃻ����2��D���%���w��=����Ô��Ŗ��  �  �
=�=iy=�'=C�=�e=;�=y=6� =�r =D��<���<���<�3�<��<���<S��<�&�<S��<���<:d�<� �<���<�h�<���<	[�<���<��<�Q�<���<���<D>�<��<���<u[�<"��<�#�<؉�<��<�c�<���<�T�<|��<!J�<]��<��<^�<���<���<��<Ũ�<`��<���<a��<k��<H��<�!�<��<���<cu�<.��<��<�<�i�<ò�<E��<���<���<fs�<S�<0��< �<H��<���<V4�<{�<��<���<���<��<;$�<�2�<�@�<�M�<ZV�<�U�<�E�<� �<�<���<�<���<�	�<�v�<�<�i�<;��<5��<.|�<@f�<%k�<���<˯�<u��<�<�3�<�G�<�G�<O2�<�	�<|ф<���<�I�<�|<Ӂw<~s<U�n<Bj<�e<]'a<?�\<�GX<%�S<��O<�^K<A-G<��B<#�><|o:<]�5<2S1<Ё,<Y�'<�n"<3F< <�<�< c	<��<� <� �;y�;�&�;3�;%
�;���;���;�R�;S��;曶;eh�;��;A��;x�;(\�;Pu�;��{;̦l;�,^;�P;�B;�i5;��(;o1;/;�;j�:C��:n��:i��:҂�:{��:>V�:�Xs:�L:��%:�]:)��9��9�r!9�"�8Y�7F�)�mҡ��ܸQ3��5��c:��m^�A��j���yPĹ��鹍	����O2��EF��{Y��l��+~�����	�����pࢺ����Fѳ�(Ȼ��ú�P˺�Ӻ={ܺ�溣#�������$\��L��?���%�-�+�3�<9�h�=��oA��]D���F���H�M`J�^TL�ưN��Q�
OU�_�Y���^��#d��i���o��tu�H
{��7���ւ�i��4�����������������@F��U����  �  ;
=&�=q=�=F�=�V=4�=�e=�� =Y =P��<��<���<��<M:�<���<6<�<`��<��<�n�<.9�<"��<z��<�K�<p��<$F�<6��<���<�R�<p��<	�<%a�<D��<�-�<6��<���<[�<��<��<O��<���<�Z�<E��<�=�<���<���<�B�<�o�<��<���<?z�<h�<vY�<�V�<h�<$��<���<R8�<���<�8�<���<rX�<���<�F�<��<þ�<:��<֥�< h�<��<���<�'�<���<�	�<�f�<���<���<��<	6�<dD�<�J�<�M�<[P�<?R�<�Q�<;I�<R3�<�	�<Wȴ<�l�<���<p�<�٪<�?�<S��<�%�<߶�<�d�<2�<G�<>)�<�J�<-{�<n��<��<,�<~(�<Y,�<�<g��<5Ƅ<���<TQ�<*.|<$�w<�Ws<��n<��j<�f<V�a<�]<"�X<i,T<��O<�sK<�-G<��B<ԣ><�E:<�5<�1<�>,<a:'<�"<r�<�<�<e�<��< G<D <R�;�s�;[<�;�=�;�T�;v\�;48�;���; ,�;�?�;�"�;��;���;ş�;��;���;��|;jBn;��_;k�Q;�/D;��6;�%*;;
;�;F;��:O�:���:XU�:n��:᫞:?�:7n: 0F:s:��9c�95$d9sM�8y�8�׷�w���޸'	����>�2��lL��Ln��0�������"ɹ�<�U�	�:�m\0�#�B�ǪT�3f�kKw�th��i��S���`���p@���G��h����eúx�˺�iԺ�ݺ�(躨��t� �n����i�����,�'��:/���5��g;�6@�%�C�iF���H�Q4J���K���M���O��R�\"V�@`Z�i7_�yd���i�sto�_�t��z����������d������@?��tގ�Is����C\���  �  �=�=�j=�=ʵ=>L=R�=sX=� =)H =Z�<�z�<d��<���<w
�<�|�<��<G��<��<N�<�<J��<X��<�6�<���<�6�<;��<}��<�Q�<��<P�<�u�<���<uN�<۸�<�<g}�<���<�3�<��<���<K\�<���<�3�<���<V��<./�<�Y�<~l�<#k�<"[�<E�<(2�<�+�<:�<�b�<$��<$
�<τ�<N�<_��<Q9�<Q��<7.�<�~�<���<}��<O��<�^�<��<ѥ�<"1�<���<>"�<�<��<��<A�<�X�<b�<b�<�]�<[X�<QS�<|L�<!?�<g%�<��<��<�V�<�߯<T�<R��<��<#��<���<;��<�4�<��<��<���<�#�<�X�<���<eː<���<q�<��<�	�<��<���<s��<^T�<LC|<��w<��s<a/o<)�j<�^f<��a<*]]<��X<!TT<C�O<�}K<*G<��B<��><P&:<-�5<>�0<�,<�'<��!<��<x^<6<�5<�l<_�<�G�;`M�;��;��;���;d��;O��;���;Y}�;�ܽ;3��;��;s˥;L��;���;��;$H�;E�};�>o;�a;��R;=:E;��7;��*;*�;��;�;v��:uj�:߸�:�6�:�|�:�D�:���:��j:�@B:�:���9&!�9��L9l{�8ot7��H���ø�n�#���-���@��X��ly��.�����{�̹���9l
�?�AY/�<�@���Q�\]b�!s��$��1+�� ���n<���觺�e��`����lú+̺�!պ�޺eK��3���I����=������!!��')��0�h?7���<� �A�PE�y�G��I��EK�\�L��eN�7�P��DS��V���Z���_��d�nj��Zo�5�t��y�vU~�����Y����z���������zv��'���œ�8L���  �  ��=��=�S=�=��=�7=!�=ZU=�� =�_ =W��<���<{�<(=�<&��<s��<�}�<��<��<Yi�<��<��<Nb�<N��<�t�<;��<�M�<~��<g�<Cb�<s��<��<��<��<0J�<��<�	�<�f�<!��<�!�<т�<h��<pJ�<«�<!�<�T�<ٔ�<���<Y��<^��<���<���<���<� �<��<�B�<-��<���<v1�<8��<��<_z�<��<$+�<�a�<�|�<(z�<�Z�<
!�<���<Rm�<���<Zx�<R��<gL�<��<���<k�<�<�<�U�<f�<�p�<fw�<nz�<�x�<�n�<VY�<m4�<7��<���<aU�< �<�r�<���<Â�<��<ؽ�<My�<�L�<8�<�8�<gK�<�i�<���</��<Ȏ<�Ռ<xՊ<'ƈ<���<6��<mV�<�&�<��{<U�w<"3s<+�n<uj<f<k�a<�0]<N�X<�TT<5�O<��K<BHG<��B<q�><A>:<��5<%%1<�i,<��'<A�"<ئ<��<��<��<-]
<o�<Ʊ<dQ�;v��;�&�;t��;���;���;[3�;��;��;�U�;@p�;�~�;���;S��;��;؄�;�)�;[�u;1�g;Z;P�L;��?;��2;K�&;�f;�;5;ܢ�:t�:-��:u��:3��:_��:xV�:,�f:v{A:�:y��9��99ފ9�<9���8��V8��60�E=����޸����C�8�w��}���r��'޹=���m��0'��9���K�W�]�5eo����������\���ݜ��`��4¯�����Gº4D˺�ԺG�޺P麵����� �����lH�ȵ���$���+���1��l7��$<��@�\oC��>F�;�H��(K�^�M���P�$�S� �W���[�Ԑ`���e���j�[ p��3u��Rz�}[�&-�������:��OЉ��n�����Ʈ��QA���Ȗ��  �  ��=��=U=��=�=n:=�=�X=F� =�c =���<4��<��<�H�<��<�<���<�<(��<qq�< �<P��<�g�<��<�x�<l��<P�<���<�<=`�<���<a�<�{�<���<cA�<1��<�<�^�<��<�<��<>��<�J�<���<��<�X�<B��<���<X��<��<���<���<] �<u�<D$�<N�<���<+��<!<�<��<5�<��<���<1�<-g�<-��<�}�<f]�<�"�<���<l�<���<�s�<���<_D�<��<Q��<(�<�3�<1N�<`�<_l�<�t�<|y�<y�<�p�<\�<8�<��<ķ�<X[�<��<]z�<��<���<�"�<\ɠ<-��<yX�<MC�<�C�<U�<r�<L��<޴�<Ύ<1ی<�ي<�Ɉ<g��<̄�<�V�<[%�<I�{<��w<�%s<��n<�cj<�e<��a<@ ]<M�X<#JT<�O<��K<�GG<E�B<��><�D:<��5<�.1<�t,<Y�'< �"<��<��<�<I<u
<�<��<�~�;���;�L�;M�;���;l��;RK�;���;�/�;�c�;�z�;��;Ԓ�;z��;���;op�;X�;�u;��g;�Y;�VL;MK?;ͻ2;S�&;�Q;]�;{:;��:N��:���:l��:�
�:\�:�Æ:όg:��B:7X:2�9���9�ԍ9�}B9�=�8�xl8��7��!o��N�׸���+,A�quu�����A����ݹ�~����R�'�J,:��uL�}|^�up��L��!���1㓺LS�����-��} ��%º>5˺-�Ժ�i޺W麤���4� �"w����j��m���$�:c+�D�1�\7���;���?�~C���E��{H���J�}M��YP�U�S�JuW���[�d|`�	�e���j��p��Mu��yz�[��;M��^҄��^��+�K���,�����N���ϖ��  �  �=&�=IX=n=��=JA=��=�a=�� =�o =���<C�<�.�<�j�<H��<�'�<n��<{<�<���<���<�4�</��<[w�<T�<ă�< ��<�U�<¯�<�<�Y�<���<�	�<�f�<��<'�<���<���<2H�<[��<+�<w�<8��<UK�<���<N�<�b�<���<<��<��<n
�<��<��<��<@*�<E�<|p�<���<��<[�<X��<k/�<I��<��<�A�<Pu�<��<j��<dd�<o&�<���<�g�<���<Be�<���<�,�<�|�<y��<{��<�<�7�<�M�<�^�<Ll�<�u�<�y�<�t�<qc�<�A�<��<Ʊ<'l�<q�<��<W�<���< B�<��<W��<mz�<d�<b�<�p�<���<P��<Ȑ<�ގ<��<�<�ӈ<���<���<WV�<g �<T�{<�gw<|�r<��n<�/j<��e<�Za<��\<�X<�)T<��O<=�K<�DG</ C<ҳ><OV:<@�5<�I1<`�,<�'<��"<7�<��<�<�U<�
<�K<j<��;{<�;)��;�g�;�)�;Q��;x��;��;�`�;犸;{��;���;���;W��;�Ӑ;�1�;ὁ;m�t;0�f;�X;��K;��>;-2;�P&;�;Df;�B;Y�:#"�:u�:���:���:���:���:l]j:5�E:��":pz:�:�9c�9�S9��9�o�8*ֻ7 ���m�V*ĸ~]��9��0o��򕹓ʷ�$cܹ�a�%���(�D�;�ݷN��Ba�K�s������+��dl������F˧��Ű�y����Lº�˺85Ժ��ݺ�b�"��/ ����U��N�A��e�#�2f*���0���5���:�w�>��(B�;E���G�@J���L�x�O��7S��W�/u[�.F`��le���j�>5p���u�r�z�b��h���>9��Rɇ��Z���팻-|��� ��Dy���喻�  �  {�=��=Y\=�=խ=K=��=wo=�� =l� =t =�5�<~a�<���<���<&\�<G��<%j�<��<���<VS�<���<���<>�<��<���<�\�<V��<> �<iM�<��<*��<�D�<��<p��<f\�<���<T#�<���<���<�g�<:��</J�<r��<��<]p�<ݶ�<���<~�<'�<4�<$=�< H�<>Z�<ux�<���<*��<�0�<S��<��<%V�<���<��<�Y�<���<��<k��<Wm�<t*�<��<�^�<>��<�L�<��<��<�Q�<l��<���< ��<��<S/�<!H�<j]�<`n�<�x�<�y�<�l�<UO�<��<�ڱ<ބ�<� �<4��<�B�<֥<
s�<��<�ܞ<���<��<���<ޛ�<���<5˒<��<��<Q��<R��< �<���<|��<T�<��<�{<35w<��r<DJn<��i<-ne<	a<5�\<xEX<�S<X�O<frK< <G<)C<m�><�m:<c�5<"p1<"�,<j�'<#<n2<\M<�w<��<�%<P�<z<��;~��;Ge�;���;/��;�W�;���;�_�;��;o��;�;9��;W��;�u�;���;�Ȉ;�9�;B�s;}e;�W;�QJ;B=;&@1;�%;��;n.;0A;Uh�:���:6[�:y��:N�:ǐ�:Sщ:�n:ݝJ:�a(:�:�'�9���9�en9��"9$�8�M68lI ���)�t�-���r;/�(Lf�Cm���@���۹p�A��9f*�z�>�1xR��e�´x�����َ�>헺٠�������d��~�ºI
˺��Ӻ�2ݺ"t續��, ��;�%��5��Y�K"�h�(���.��N4�<9��(=���@�B�C�$�F��=I��L��O�\�R��V��[�� `�[Pe��j�6�p�"(v���{�K���xB��ᅻAv�������������h����������  �  ��=��=�_=�=8�=�U=��=r=�=� =�& =�p�<s��<���<)7�<ў�<8�<{��<6:�<X��<"x�<@�<��<�,�<ܢ�<�	�<b�<���<w��<j:�<x�<��<��<�i�<X��<�"�<"��<���<�a�<���<;P�<d��<	E�<���<{"�<�}�<+��<��<�,�<�H�<�\�<�l�<P~�<Ɩ�<���<<��<�&�<�q�<,��<�%�<��<C��<d4�<�u�<��<���<-��<�t�<�+�<��<P�<���<�*�<r��<W��<��<-U�<���<���<��<��<�'�<�F�<5a�<t�<�{�< u�<�\�<�0�<��<Z��<5C�<�ܪ<�s�<��<ణ<�`�<� �<�<�ך<z͘<qі<�ߔ<�<�<��<#�<{	�<}�<�Ć<ٍ�<�M�<h�<`~{<�v<Her<��m<ii<��d<(�`<'7\<w�W<��S<�vO<NK<�)G<�C<��><ʃ:<Z6<��1<�,<�7(<�f#<s�<ٶ<��<�><׮<�D<�<���;%��;�8�;,��;�G�;���;�[�;��;���;��;?հ;���;b�;11�;��;F7�;���;�$r;��c;��U;��H;�;;��/;a�$;��;`�;";��:�c�:�D�:�:iʰ:�^�:���:(�s:%�P:�</:w':N��9�ɴ9�B�9��C9��9�p�8jŽ7�έ�+5��j��s#���\��ᎹQ�9GڹS��&{�|,-�^�B��W���k����RB��0n���J��У�e���쳺󤻺Rú;2˺�Ӻ|�ܺ����w�Vv���*�d��������� �+�&���,�--2�W�6�-%;�.�>��B�E�"H��K��CN��Q��V�H�Z���_�Je��k�4q�@�v���|��F����������]���勻�W��H�������+��dS���  �  w�=ӧ=}`=�=�=<_=6�=U�=� =B� =2C =��<E��<�.�<S��<"��<�_�<E��<�q�<��<%��<\2�<g��<9>�<��<"�<Mb�<^��<=��<2 �<iZ�<q��<���<_)�<�~�<���<�D�<ڴ�<l-�<���<>1�<ڶ�<�9�<���<9&�<���<K��<��<�G�<Bk�<*��<��<V��<\��<��<�5�<ys�<���<,�<>b�<���<$�<�V�<`��<F��<ٽ�<��<�w�<�'�<���<K:�<���<���<�N�<���<���<��<�A�<�s�<m��<���<���<�(�<M�<i�<�x�<�x�<�e�<�?�<m�<Լ�<�f�<	�<��<�K�<��</��<�m�<�?�<� �<H�<o�<�<��<�'�<�-�<�)�<t�<���<�ǆ<܉�<A�<��<�;{<��v<k�q<mem<��h<jkd<�`<ٶ[<�xW<LS<�.O<aK<�
G<�B<_�><^�:<;76<��1<�&-<w(<��#<�<�*<ys<��<�I<��<��<���;��;f �;�y�;U��;_�;���;�
�;�'�;�;�߰;͊�;A*�;*ї;�;9��;�T;�2p;v�a;��S;��F;]&:;�h.;>a#;�;�2;��;���:	��:���::�:�%�:�:�+�:�#y:�W:"�6:��:�9�
�9���9�h9	$9O��8� H8B�/4��A�XŸ�����T��G��Ա�!�ڹb;����}�0�^�G�l�]�nfs�%ꃺŚ��þ��Y��Lp�����HQ��Z[���fĺ$�˺��Ӻ�.ܺ���h�'	��:@���
��q�6�����$�Xz*�2�/���4���8�%�<�|H@�i�C�_�F���I��vM�LLQ��U� fZ���_�koe��{k��q�_�w��3~����Z��Ї�u�������S��Ï��G������鲗��  �  ��=��=�]=	=S�=�e=2=P�={3=�� =�_ =���<P3�<�}�<h��<:8�<Z��<�#�<Ȩ�<�3�<H��<sL�<���<�I�<���<��<�[�<��<���<���<.�<oa�<I��<P��<>2�<���<%��<�p�<���<�{�<
�<$��<�'�<ѫ�<#�<���<��<�&�<^�<��<���<~��<���<v�<�N�<���<���<��<�Q�<E��<���<�5�<�u�<���<���<���<ū�<Gs�<p�<4��<+�<�|�<���<V�<)N�<��<U��<���<�'�<�^�<q��<���<��<�1�<�V�<\n�<�t�<(h�<"H�<��<ԯ<���<l3�<�ݨ<���<3=�<k��<̽�<͎�<�k�<dT�<�G�<mC�<ED�<�E�<�C�<�8�<!�<���<2Ć<�~�<]-�<ۦ<��z<s/v<�|q<��l<oHh<��c<Qn_<�&[<o�V<��R<��N<&�J<B�F<8�B< �><ې:< C6<��1<�M-<��(<[$<zN<�<��<�g<��<��<W><� <2��;(�;o9�;y��;��;��;�D�;�H�;0!�;ϰ;�[�;�֟;+U�;
�;9��;}a};bn;eY_;�rQ;�ZD;�8;��,;�!;p�;:b;�O;���:���:�5�:��:�)�:��:1'�:�K~:g�]:�t>:Od!:��:x�9��9ꎇ9^IG9�9��8}�7\������ۨ��0P�b`���m��ݹ�`��;��5�[�M��Fe���{�d����k��i���I䣺񉫺咲�0)��f�����źɩ̺�Ժ�?ܺy�ѹﺦ����v��	����f� ���y"�(��C-��2���6���:��t>�B�L�E�RI�v�L�,�P��[U��YZ�=�_�E�e�4l���r�OCy�������������G����$��+n��B���񀔻�]��"/���  �  �=Η=�W=�=	�=�h=�
=.�=KC=!� =�z =� =Nz�<}��<�!�<I��<���< a�<���<�[�<���<&`�<���< N�<���<��<fM�<܄�<t��<���<"��<g&�<OX�<:��<���<�?�<���<#)�<Ų�<UF�<���<�y�<��<���<��<��<l��<�.�<�m�< ��<���<q �<P/�<Sa�<Y��<{��<��<�P�<B��<q��<9�<fY�<���<��<5��<M��<��<�g�<�	�<��<)��<P�<���<*��<u�<e6�<9i�<ߞ�<���<e�<W�<���<�׿<2�<�=�<�\�<�i�<c�<@I�<��<��<x��<�X�<?�<�Ŧ<,��<�B�<�
�< ۝<³�<"��<�~�<p�<f�<�]�<R�<@�<6"�<���<$��<�l�<]�<4`<��z<ɿu<��p<�El<M�g<�,c<��^<��Z<TqV<�jR<nwN<��J<B�F<7�B<-�><v�:<�?6<Z�1<�f-<��(<�@$</�<�
<{<~�<	�<�%	<��<נ <���;���;���;��;�-�;�Q�;�`�;kL�;��;��;�;�j�;Ö;o0�;+˅;nS{;�k;��\;+O;��A;$�5;A�*;�I ;ő;Gc;��; �:��: �:E��:���:���:MÑ:8c�:�\c:�E:	�):�:yK�9I��9[ �9��h9ܹ#9#V�8�$8�˚�gМ�jM�`!O�Y��*ᴹ�.��Z��J!�[�:��AT��m��S��V���i������+����ׯ�AT��K���º��Ǻ�
κ��Ժ]�ܺ���)���J��3����@����4���S �0�%�$�*�"�/�AN4�פ8��<���@���D��`H��aL�	�P�c[U���Z��7`�pbf���l���s�
�z��ƀ�����C��U6���ꌻ2_��씑�ƒ��ld��c�� ��  �  n�=��=BN==	=B�=�g=�=��=�O=�� =v� =�5 =���<��<�g�<���<�+�<���<>�<�|�<���<�l�<0��<CK�<ө�<���<�9�<�j�<h��<���<.��<���<��<�M�<���<���<b�<���<Dt�<d�<���<�T�<��<��<��<�z�<���<�/�<Vv�<���<���<0'�<`�<���<P��<^�<�T�<3��<"��<N
�<�B�<�u�<���<���<���<	��<ș�<�U�<��<�p�<��<W!�<�]�<̏�<���<)��<6�<+O�<6��<���<_�<�b�<���<w�<| �<�E�<IX�<AW�<�C�<Y�<|�<ⴭ<�v�<w7�<F��<���<��<yP�<��<��<FΙ<���<_��<���<on�<oZ�<�@�<V�<�<��<�U�<\��<�<12z<�Ou<�xp<ζk<�g<��b<�4^<��Y<��U<�Q<�N<�;J<�aF<mzB<�}><5e:<�.6<Y�1<�q-<��(<�q$<`�<h<K�<�y<�<ϴ	<�c<!<P��;s��;�r�;+g�;�j�;�m�;�`�;3�;�ݸ;�[�;���;��;�&�;Sq�;��;�Ny;��i;r�Z;��L;�?;��3;��(;�;�5;�J; �;p��:��:/^�:���:�ֳ:25�:��:;-�:�Ih:��K:
1:8�:=T :GG�9��9�P�9�=9��8y�W8Y������`�ЄQ�(��[帹&�������%�Q@���Z� �t�.���0���99���K��4��P�����Vz���ĺO�ɺ�Ϻ�;ֺ(�ݺx9������y��v,�������<��k�4�#�.�(���-��N2�,�6��H;��?���C�:�G��*L���P���U�?�Z���`�J!g���m���t�R(|�h���f��5_��Ud��g����������ꖔ��G��Vؗ��_���  �  ��=~~=�C=� =a�=�d=�=��=;X=;� =�� =^L =���<WF�<]��<���<�^�<��<�)�<���<-�<9s�<��<�C�<���<��<n#�<�O�<ro�<2��<Ĝ�<P��<���<��<�R�<t��<��<t��<�;�<���<��</1�<A��<�k�<.��<�k�<���<i+�<5y�<��<�<OE�<���<L��<;�<�O�<���<}��<\��<e2�<Ia�<���<���<m��<+��<H��<���<�@�<���<�Q�<��<���<�*�<�U�<�|�<ä�<��<��<�H�<��<���<�0�<��<gǽ<E�<�,�<D�<�G�<~9�<��<w�<���<h��<�W�<�"�<%�<I��<*��<�X�<P)�<���<�ԗ<0��<��<�x�<�\�<�;�<��<�ڈ< ��<�<�<�ց<.�~<[�y<��t<�p<�7k<�f<vb<׬]<~Y<�uU<��Q<��M<��I<	 F<DB<RQ><VB:<�6<��1<�q-<�)<ה$<�! <^�<�H<j�<��<�+
<V�<ي<���;I*�;l��;��;@��;Vr�;nK�;*	�;L��;��;�M�;�s�;���;/��;��;w;u�g;U�X;ЕJ;��=;J�1;�';�';��;�7;?�;?�:��:�~�:q
�:���:Vo�:ǩ�:h�:8 l:��P:7:5�:g�:3��9�3�9���9�aQ9Ru9ʘ�8�m�@��[��@V��������W��I��"*�%�E�Q�`�U�{�4z������z������E���Է��p��Kmº�*Ǻ�̺tѺ7�׺~�޺W纫<�&3���W�ƹ�=!�Pz�������!���&���+��0��n5� :���>�5%C��G�$!L�c�P�S�U�Pl[�$la��g���n�� v���}��r��(��
\���o��y0������ױ��{����������T����  �  �= s=�9=��=I�=�`=�=��=�]=�=�� =] =Y
 =�p�<���<h(�<N��<���<sB�<k��<a�<mu�<.��<�:�<���<H��<3�<�7�<pS�<�f�<w�<���<���<���<��<�x�<���<-t�<�<Ҷ�<;e�<E�<���<�U�<���<�\�<���<0%�<�x�<���<k�<rZ�<���<x��<[6�<Az�<���<���<�"�<�O�<�v�<o��<)��<���<���<���<�z�<�-�<���<7�<��<���<��<�'�<�I�<�n�<
��<w��<"�< _�<c��<��<�\�<��<1�<W�<;1�<�8�<�.�<��<��<ɭ<q��<�n�<A�<��<}�<=��<���<�P�<F�<��<;ƕ<i��<�}�<g[�<N5�<��<�ˈ<���<�&�<���<͌~<��y<O�t<��o<��j<� f<�a<�A]<�Y<�U<N7Q<qmM<ԬI<�E<SB<�(><� :<j�5< �1<l-<)<��$<�G <�<n�<�3<`�<��
<�-<\�<��;��;�)�;��;T��;9j�;�.�;��;�c�;"��;���;
�;��;.�;0u�;�v;f;��V;��H;)<;�e0;)�%;��;��;�P
;�;���:��:���:\h�:fG�:�n�:��:a\�:��n:/zT:�;:7�#:1�:���9j�9��9>`9ʎ9+�8���?��K���l[��,��s%¹��񹷩�<�-���I���e�-��������V��,ң��ܬ��z���Һ��%��T�ĺ�<ɺ�ͺ��Һ��غj�ߺ$��E��?z���K��v�U��@�����հ��� �W�%�gu*�fl/��^4�%B9��>���B�auG�n0L��Q�1JV���[��b���h���o�Lw���~���ֹ��$$��B����!n��L{��-:���������u���  �  �=k=$3=?�=��=�]=&= �=�`=�=׸ =$g =@ =���<D��<B�<l��<C��<%Q�<*��<3�<�u�<���<�3�<F��<Z��<�<w'�<�@�<�P�<V^�<�o�<��</��<���<�V�<D��<�T�<��<М�<)N�<#��<"��<�F�<���<&R�<���<��<w�<���<��<�f�<���<��<�N�<���<��<�	�<�8�<6a�<���<'��<���<5��<a��<r��<do�<` �<>��<�$�<A{�<͹�<���<�	�<q)�<oL�<�w�<!��<���<�>�<��<t��<�E�<���<~ֻ<��<$�<�-�<r&�<��<��<�̭<��<�|�<�S�<R*�<���<�Ϡ<���<$i�<=4�<E�<ҕ<=��<��<uY�<�/�<���<��<�t�<�<���<�c~<5cy<�at<mo<m�j<�e<�Ta<{�\<J�X<�T< Q<0<M<n�I<L�E<��A<�><!	:<a�5<�1<f-<K)<��$<�] <<<ȵ<nd<�<|�
<�b<�	<�i�;=��;lU�;���;���;;`�;��;���;p8�;;���;>;b��;�΋;�	�;�!u;se;��U;��G;�;;p/;/�$;�&;�,;�	;B�;�	�:��:7��:���:���:r[�:B�:�؅:}kp:��V:X@>:R�&:�>: 0�9h��9��9	/i9u9]�8�<�5�3���D�r^_��͘��NŹޛ�����2I0���L�i�Di���{���i���������H���z��������bƺ+�ʺ�Ϻ�Ժ��ٺ٫�ͅ�iG񺈺��~M�]T��W�J�}(���������$�Σ)�l�.�#�3���8�M�=�1�B��gG��CL�NFQ��V��B\��ob�i��Bp��w�Sf�����J0������ȍ����� ���,���ֱ���)��~���ɚ��  �  ��=;h=�0=2�=�=�\=�
=2�=~a=�=f� =�j =X =s��<0��<�J�<b��<���<�U�<J��<��<yu�<���<61�<���<��<���<�!�<�9�<[I�<�U�<7f�<~��<��<��<�J�<���<�I�<��<ݓ�<6F�<"��<��<dA�<@��<CN�<���<��<$v�<3��<<�<�j�<���<_�<^W�<i��<���< �<A@�<g�<ԇ�<���<���<X��<B��<O��<[k�<��<���<��<t�<���<���<i��<@�<�@�<Lk�<��<;��<�3�<��<t��<�=�<���<%л<V�<S�<�)�<i#�<�<�<�ͭ<���<��<Z�<2�<@�<�ؠ<���<wq�<h;�<��<�Օ<P��<[��<xX�<�-�<m��<6��<�o�<��<w��<3U~<�Ry<jOt<{Xo<7|j<��e<�<a<��\<��X<�T<�P<N+M<erI<�E<��A<]><� :<��5<�1<bc-<�)<�$<�d <�<��<*u<�#<��
<�t<<r��;���;pc�;A��;���;�[�;��;��;�(�;�y�;[��;6��;���;?��;��;�t;��d;��U;��G;��:;8/;��$;��;>�;�~	;p[;��:���:���:T��:ܲ:�O�:&N�:���:��p:�bW:@/?:��':L[:Zi�9@��9��9X#l9�99ߒ�8���5�搸�;���`�����rƹ��������%1�Z�M��6j����/(��� ��󲦺i����=��Uh��Z�º��ƺ1˺sϺaԺ�)ں�����s�����P�WJ�h@�}%����!��Ј��g$��])�5i.�r�3�X�8��=���B�feG��LL��XQ�ݪV�c\�u�b�RKi��up�2�w�l������LY��:Њ�+��������#���(��-ۖ� O��
����暻�  �  �=k=$3=?�=��=�]=&= �=�`=�=׸ =$g =@ =���<D��<B�<l��<C��<%Q�<*��<3�<�u�<���<�3�<F��<Z��<�<w'�<�@�<�P�<V^�<�o�<��</��<���<�V�<D��<�T�<��<М�<)N�<#��<"��<�F�<���<&R�<���<��<w�<���<��<�f�<���<��<�N�<���<��<�	�<�8�<6a�<���<'��<���<5��<a��<r��<do�<` �<>��<�$�<A{�<͹�<���<�	�<r)�<pL�<�w�<"��< ��<�>�<��<u��<�E�<���<ֻ<��<$�<�-�<s&�<��<��<�̭<��<�|�<�S�<S*�<���<�Ϡ<���<#i�<=4�<E�<ҕ<<��<��<tY�<�/�<���<��<�t�<~�<���<�c~<4cy<�at<mo<l�j<�e<�Ta<{�\<J�X<�T< Q<1<M<p�I<M�E<��A<�><#	:<c�5<�1<f-<M)<��$<�] <=<ȵ<od<�<|�
<�b<�	<�i�;;��;iU�;���;���;7`�;��;���;l8�;댯;���;:;_��;�΋;�	�;�!u;ne;��U;��G;�;;p/;-�$;�&;�,;�	;A�;�	�:��:6��:���:���:r[�:B�:�؅:}kp:��V:X@>:R�&:�>: 0�9h��9��9	/i9u9]�8�<�5�3���D�r^_��͘��NŹޛ�����2I0���L�i�Di���{���i���������H���z��������bƺ+�ʺ�Ϻ�Ժ��ٺ٫�ͅ�iG񺈺��~M�]T��W�J�}(���������$�Σ)�l�.�#�3���8�M�=�1�B��gG��CL�NFQ��V��B\��ob�i��Bp��w�Sf�����J0������ȍ����� ���,���ֱ���)��~���ɚ��  �  �= s=�9=��=I�=�`=�=��=�]=�=�� =] =Y
 =�p�<���<h(�<N��<���<sB�<k��<a�<mu�<.��<�:�<���<H��<3�<�7�<pS�<�f�<w�<���<���<���<��<�x�<���<-t�<�<Ҷ�<;e�<E�<���<�U�<���<�\�<���<0%�<�x�<���<k�<rZ�<���<x��<[6�<Az�<���<���<�"�<�O�<�v�<o��<)��<���<���<���<�z�<�-�<���<7�<��<���<��<�'�<�I�<�n�<��<x��<#�<_�<d��<��<�\�<��<2�<Y�<=1�<�8�<�.�<��<��<ɭ<r��<�n�<A�<��<~�<=��<���<�P�<E�<��<:ƕ<g��<�}�<e[�<M5�<��<�ˈ<���<�&�<���<ʌ~<��y<M�t<��o<��j<� f<�a<�A]<�Y< U<O7Q<smM<֬I<�E<VB<�(><� :<m�5<�1<l-<)<��$<�G < �<o�<�3<a�<��
<�-<[�<��;��;�)�;��;N��;3j�;�.�;��;�c�;��;���;
�;��;.�;*u�;�v;�f;��V;��H;#<;�e0;%�%;��;��;�P
;�;���:��:���:[h�:eG�:�n�:��:a\�:��n:/zT:�;:7�#:1�:���9j�9��9>`9ʎ9+�8���?��K���l[��,��s%¹��񹷩�<�-���I���e�-��������V��,ң��ܬ��z���Һ��%��T�ĺ�<ɺ�ͺ��Һ��غj�ߺ$��E��?z���K��v�U��@�����հ��� �W�%�gu*�fl/��^4�%B9��>���B�auG�n0L��Q�1JV���[��b���h���o�Lw���~���ֹ��$$��B����!n��L{��-:���������u���  �  ��=~~=�C=� =a�=�d=�=��=;X=;� =�� =^L =���<WF�<]��<���<�^�<��<�)�<���<-�<9s�<��<�C�<���<��<n#�<�O�<ro�<2��<Ĝ�<P��<���<��<�R�<t��<��<t��<�;�<���<��</1�<A��<�k�<.��<�k�<���<i+�<5y�<��<�<OE�<���<L��<;�<�O�<���<}��<\��<e2�<Ia�<���<���<m��<+��<H��<���<�@�<���<�Q�<��<���<�*�<�U�<�|�<Ĥ�<���<��<�H�<��<���<�0�<��<iǽ<G�<�,�<D�<�G�<�9�<��<y�<���<i��<�W�<�"�<&�<J��<*��<�X�<O)�<���<�ԗ</��<
��<�x�<�\�<�;�<��<�ڈ<��<�<�<�ց<+�~<W�y<��t<�p<�7k<
�f<vb<׬]<~Y<�uU<��Q<��M<��I< F<DB<VQ><[B:<�6<��1<�q-<�)<۔$< " <a�<�H<k�<��<�+
<V�<؊<���;D*�;f��;���;8��;Mr�;dK�; 	�;B��;|�;�M�;�s�;쐕;&��;��;�~w;h�g;I�X;ƕJ;��=;C�1;�';�';��;�7;=�;?�:��:�~�:o
�:���:Uo�:ǩ�:g�:7 l:��P:7:5�:g�:3��9�3�9���9�aQ9Ru9ʘ�8�m�@��[��@V��������W��H��"*�%�E�Q�`�U�{�4z������z������E���Է��p��Kmº�*Ǻ�̺tѺ7�׺~�޺W纫<�&3���W�ƹ�=!�Pz�������!���&���+��0��n5� :���>�5%C��G�$!L�c�P�S�U�Pl[�$la��g���n�� v���}��r��(��
\���o��y0������ױ��{����������T����  �  n�=��=BN==	=B�=�g=�=��=�O=�� =v� =�5 =���<��<�g�<���<�+�<���<>�<�|�<���<�l�<0��<CK�<ө�<���<�9�<�j�<h��<���<.��<���<��<�M�<���<���<b�<���<Dt�<d�<���<�T�<��<��<��<�z�<���<�/�<Vv�<���<���<0'�<`�<���<P��<^�<�T�<3��<"��<N
�<�B�<�u�<���<���<���<	��<ș�<�U�<��<�p�<��<W!�<�]�<͏�<���<+��<7�<,O�<8��<���<b�<�b�<���<z�< �<�E�<LX�<DW�<�C�<\�<~�<崭<�v�<y7�<H��<���<��<yP�<��<��<EΙ<���<]��<���<ln�<mZ�<�@�<T�<�<��<�U�<Y��<�<-2z<�Ou<�xp<̶k<�g<��b<�4^<��Y<��U<��Q<�N<�;J<�aF<szB<�}><;e:</6<_�1<�q-<��(<�q$<c�<h<N�<�y<�<ϴ	<�c<!<K��;m��;�r�;"g�;�j�;�m�;�`�;s3�;�ݸ;�[�;���;��;�&�;Hq�;��;�Ny;��i;d�Z;�L;�?;��3;��(;�;�5;�J;��;k��:��:,^�:���:�ֳ:15�:��::-�:�Ih:��K:	1:7�:=T :GG�9��9�P�9�=9��8y�W8X������`�ЄQ�(��[帹&�������%�Q@���Z� �t�.���0���99���K��4��P�����Vz���ĺO�ɺ�Ϻ�;ֺ(�ݺx9������y��v,�������<��k�4�#�.�(���-��N2�,�6��H;��?���C�:�G��*L���P���U�?�Z���`�J!g���m���t�R(|�h���f��5_��Ud��g����������ꖔ��G��Vؗ��_���  �  �=Η=�W=�=	�=�h=�
=.�=KC=!� =�z =� =Nz�<}��<�!�<I��<���< a�<���<�[�<���<&`�<���< N�<���<��<fM�<܄�<t��<���<"��<g&�<OX�<:��<���<�?�<���<#)�<Ų�<UF�<���<�y�<��<���<��<��<l��<�.�<�m�< ��<���<q �<P/�<Sa�<Y��<{��<��<�P�<B��<q��<9�<fY�<���<��<5��<M��<��<�g�<�	�<	��<*��<P�<���<+��<v�<f6�<:i�<��<���<h�<W�<���<�׿<5�<�=�<�\�<�i�<c�<CI�<��<��<{��<�X�<A�<�Ŧ<-��<�B�<�
�<۝<���< ��<�~�<
p�<f�<�]�<|R�<@�<3"�<���<!��<�l�<[�</`<��z<ſu<��p<�El<L�g<�,c<��^<��Z<VqV<�jR<rwN<��J<H�F<=�B<3�><}�:<�?6<`�1<�f-<��(<�@$<3�<<"{<��<
�<�%	<��<ՠ <���;���;���;��;�-�;�Q�;�`�;]L�;��;��;�;�j�;�;c0�; ˅;[S{;��k;��\;O;��A;�5;9�*;�I ;��;Cc;��;�:��: �:B��:���:���:LÑ:8c�:�\c:�E:	�):�:yK�9I��9[ �9��h9ܹ#9#V�8�$8�˚�fМ�jM�_!O�Y��*ᴹ�.��Z��J!�[�:��AT��m��S��V���i������+����ׯ�AT��K���º��Ǻ�
κ��Ժ]�ܺ���)���J��3����@����4���S �0�%�$�*�"�/�AN4�פ8��<���@���D��`H��aL�	�P�c[U���Z��7`�pbf���l���s�
�z��ƀ�����C��U6���ꌻ2_��씑�ƒ��ld��c�� ��  �  ��=��=�]=	=S�=�e=2=P�={3=�� =�_ =���<P3�<�}�<h��<:8�<Z��<�#�<Ȩ�<�3�<H��<sL�<���<�I�<���<��<�[�<��<���<���<.�<oa�<I��<P��<>2�<���<%��<�p�<���<�{�<
�<$��<�'�<ѫ�<#�<���<��<�&�<^�<��<���<~��<���<v�<�N�<���<���<��<�Q�<E��<���<�5�<�u�<���<���<���<ū�<Gs�<p�<4��<+�<�|�<���<W�<*N�<���<V��<���<�'�<�^�<t��<���<��<�1�<�V�<`n�<�t�<,h�<%H�<��<ԯ<���<n3�<�ݨ<���<4=�<l��<̽�<͎�<�k�<cT�<�G�<kC�<BD�<�E�<�C�<�8�<!�<|��</Ć<�~�<Z-�<զ<��z<o/v<�|q<��l<nHh<��c<Rn_<�&[<r�V<��R<��N<+�J<H�F<>�B<&�><�:<C6<��1<�M-<��(<`$<~N<�<��<�g<��<��<V><� <,��;!�;f9�;n��;��;��;�D�;�H�;!!�;ϰ;�[�;�֟;U�;��;.��;ha};Pn;UY_;�rQ;�ZD;�8;��,;�!;j�;5b;�O;���:���:�5�:��:�)�:��:0'�:�K~:f�]:�t>:Nd!:��:w�9��9ꎇ9]IG9�9��8}�7\������ۨ��0P�b`���m��ݹ�`��;��5�[�M��Fe���{�d����k��i���I䣺񉫺咲�0)��f�����źɩ̺�Ժ�?ܺy�ѹﺦ����v��	����f� ���y"�(��C-��2���6���:��t>�B�L�E�RI�v�L�,�P��[U��YZ�=�_�E�e�4l���r�OCy�������������G����$��+n��B���񀔻�]��"/���  �  w�=ӧ=}`=�=�=<_=6�=U�=� =B� =2C =��<E��<�.�<S��<"��<�_�<E��<�q�<��<%��<\2�<g��<9>�<��<"�<Mb�<^��<=��<2 �<iZ�<q��<���<_)�<�~�<���<�D�<ڴ�<l-�<���<>1�<ڶ�<�9�<���<9&�<���<K��<��<�G�<Bk�<*��<��<V��<\��<��<�5�<ys�<���<,�<>b�<���<$�<�V�<`��<G��<ڽ�<��<�w�<�'�<���<K:�<���<���<�N�<���<���<��<�A�<�s�<p��<���<���<�(�< M�<i�<�x�<�x�<�e�<�?�<p�<׼�<�f�<	�<��<�K�<��<0��<�m�<�?�<� �<F�<n�<�<��<�'�<�-�<�)�<q�<���<�ǆ<ى�<A�<��<�;{<��v<h�q<jem<��h<ikd<�`<۶[<�xW<LS<�.O<fK<�
G<�B<e�><d�:<A76<��1<�&-<!w(<��#<#�<�*<{s<��<�I<��<��<���;���;_ �;�y�;K��;_�;t��;�
�;}'�;��;�߰;���;3*�;ї;蒏;.��;�T;�2p;f�a;t�S;��F;S&:;�h.;7a#;�;~2;��;���:��:���:7�:�%�:�:�+�:�#y:�W:!�6:��:�9�
�9���9�h9$9O��8� H8o�/4��A�XŸ�����T��G��Ա�!�ڹb;����}�0�^�G�l�]�nfs�%ꃺŚ��þ��Y��Lp�����HQ��Z[���fĺ$�˺��Ӻ�.ܺ���h�'	��:@���
��q�6�����$�Xz*�2�/���4���8�%�<�|H@�i�C�_�F���I��vM�LLQ��U� fZ���_�koe��{k��q�_�w��3~����Z��Ї�u�������S��Ï��G������鲗��  �  ��=��=�_=�=8�=�U=��=r=�=� =�& =�p�<s��<���<)7�<ў�<8�<{��<6:�<X��<"x�<@�<��<�,�<ܢ�<�	�<b�<���<w��<j:�<x�<��<��<�i�<X��<�"�<"��<���<�a�<���<;P�<d��<	E�<���<{"�<�}�<+��<��<�,�<�H�<�\�<�l�<P~�<Ɩ�<���<<��<�&�<�q�<,��<�%�<��<C��<d4�<�u�<��<���<-��<�t�<�+�<��<P�<���<�*�<s��<X��<��<.U�<���<���<���<��<�'�<�F�<7a�<t�<�{�<#u�<�\�<�0�<��<\��<8C�<�ܪ<�s�<��<ᰣ<�`�<� �<�<�ך<y͘<oі<�ߔ<�<�<��<!�<x	�<z�<�Ć<֍�<�M�<f�<\~{<�v<Eer<��m<ii<��d<)�`<(7\<y�W<��S<�vO<NK<�)G<�C<��><Ѓ:<_6<��1<�,<�7(<�f#<w�<ܶ<��<�><خ<�D<�<���; ��;�8�;$��;�G�;���;�[�;��;���;��;3հ;���;�a�;&1�;��;=7�;���;�$r;��c;��U;��H;�;;��/;[�$;��;\�;
";	��:�c�:�D�:�:gʰ:�^�:���:'�s:$�P:�</:v':M��9�ɴ9�B�9��C9��9�p�8jŽ7�έ�+5��i��s#���\��ᎹQ�9GڹS��&{�|,-�^�B��W���k����RB��0n���J��У�e���쳺󤻺Rú;2˺�Ӻ|�ܺ����w�Vv���*�d��������� �+�&���,�--2�W�6�-%;�.�>��B�E�"H��K��CN��Q��V�H�Z���_�Je��k�4q�@�v���|��F����������]���勻�W��H�������+��dS���  �  {�=��=Y\=�=խ=K=��=wo=�� =l� =t =�5�<~a�<���<���<&\�<G��<%j�<��<���<VS�<���<���<>�<��<���<�\�<V��<> �<iM�<��<*��<�D�<��<p��<f\�<���<T#�<���<���<�g�<:��</J�<r��<��<]p�<ݶ�<���<~�<'�<4�<$=�< H�<>Z�<ux�<���<*��<�0�<S��<��<%V�<���<��<�Y�<���<��<k��<Xm�<t*�<��<�^�<?��<�L�<��<��<�Q�<n��<���<��<��<U/�<#H�<l]�<bn�<�x�<�y�<�l�<WO�<��<�ڱ<���<� �<6��<�B�<֥<s�<��<�ܞ<���<��<���<ݛ�<���<3˒<��<���<O��<O��<�<���<z��<T�<��<�{<15w<��r<BJn<��i<-ne<	a<6�\<zEX<�S<[�O<jrK<$<G<.C<q�><�m:<h�5<'p1<&�,<n�'<#<q2<_M<�w<��<�%<P�<z<��;z��;Ae�;���;'��;�W�;���;{_�;ؤ�;e��;鷰;/��;M��;�u�;���;}Ȉ;�9�;5�s;}e;�W;�QJ;;=; @1;�%;ܛ;j.;.A;Qh�:���:4[�:w��:N�:Ɛ�:Sщ:�n:ܝJ:�a(:~�:�'�9���9�en9��"9$�8�M68kI ���)�t�-���r;/�(Lf�Cm���@���۹p�A��9f*�z�>�1xR��e�´x�����َ�>헺٠�������d��~�ºI
˺��Ӻ�2ݺ"t續��, ��;�%��5��Y�K"�h�(���.��N4�<9��(=���@�B�C�$�F��=I��L��O�\�R��V��[�� `�[Pe��j�6�p�"(v���{�K���xB��ᅻAv�������������h����������  �  �=&�=IX=n=��=JA=��=�a=�� =�o =���<C�<�.�<�j�<H��<�'�<n��<{<�<���<���<�4�</��<[w�<T�<ă�< ��<�U�<¯�<�<�Y�<���<�	�<�f�<��<'�<���<���<2H�<[��<+�<w�<8��<UK�<���<N�<�b�<���<<��<��<n
�<��<��<��<@*�<E�<|p�<���<��<[�<X��<k/�<I��<��<�A�<Pu�<��<j��<dd�<o&�<���<�g�<���<Be�<���<�,�<�|�<z��<|��<�<�7�<�M�<�^�<Ml�<�u�<�y�<�t�<sc�<�A�<��<Ʊ<(l�<r�<��<X�<���< B�<��<W��<mz�<d�<b�<�p�<���<O��<Ȑ<�ގ<��<�<�ӈ<���<���<VV�<f �<Q�{<�gw<z�r<��n<�/j<��e<�Za<��\<�X<�)T<��O<@�K<�DG<2 C<ճ><RV:<C�5<�I1<d�,<�'<��"<9�<��<�<�U<�
<�K<i<��;x<�;%��;�g�;�)�;K��;q��;��;�`�;���;t��;���;���;Q��;�Ӑ;�1�;۽�;d�t;(�f;�X;��K;��>;-2;�P&;�;Af;�B;V�:!"�:u�:���:���:���:���:k]j:4�E:��":pz:�:�9c�9�S9��9�o�8*ֻ7 ���m�V*ĸ~]��9��0o��򕹓ʷ�$cܹ�a�%���(�D�;�ݷN��Ba�K�s������+��dl������F˧��Ű�y����Lº�˺85Ժ��ݺ�b�"��/ ����U��N�A��e�#�2f*���0���5���:�w�>��(B�;E���G�@J���L�x�O��7S��W�/u[�.F`��le���j�>5p���u�r�z�b��h���>9��Rɇ��Z���팻-|��� ��Dy���喻�  �  ��=��=U=��=�=n:=�=�X=F� =�c =���<4��<��<�H�<��<�<���<�<(��<qq�< �<P��<�g�<��<�x�<l��<P�<���<�<=`�<���<a�<�{�<���<cA�<1��<�<�^�<��<�<��<>��<�J�<���<��<�X�<B��<���<X��<��<���<���<] �<u�<D$�<N�<���<+��<!<�<��<5�<��<���<1�<-g�<-��<�}�<g]�<�"�<���<l�<���<�s�<���<_D�<��<Q��<(�<�3�<2N�<`�<`l�<�t�<}y�<y�<�p�<\�<8�<��<ŷ�<Y[�<��<^z�<��<���<�"�<\ɠ<-��<yX�<MC�<�C�<U�<r�<K��<ݴ�<Ύ<0ی<�ي<�Ɉ<g��<˄�<�V�<Z%�<H�{<��w<�%s<��n<�cj< �e<��a<A ]<N�X<$JT<�O<��K<�GG<F�B<��><�D:<��5<�.1<�t,<Z�'<�"<��<��<	�<I<u
<�<��<�~�;���;�L�;J�;���;h��;OK�;���;�/�;�c�;�z�;��;В�;w��;���;lp�;U�;�u;��g;�Y;�VL;KK?;ʻ2;Q�&;�Q;\�;z:;��:L��:���:k��:�
�:\�:�Æ:όg:��B:7X:~2�9���9�ԍ9�}B9�=�8�xl8��7��!o��N�׸���+,A�quu�����A����ݹ�~����R�'�J,:��uL�}|^�up��L��!���1㓺LS�����-��} ��%º>5˺-�Ժ�i޺W麤���4� �"w����j��m���$�:c+�D�1�\7���;���?�~C���E��{H���J�}M��YP�U�S�JuW���[�d|`�	�e���j��p��Mu��yz�[��;M��^҄��^��+�K���,�����N���ϖ��  �  �=;�=�A=��=��=d*=U�=U=R� =�s =� =-.�<�`�<͢�<?��<�[�<���< X�<���<I�<v�<+��<�9�<I��<�5�<���<U�< f�<��<}�<}q�<���<�'�<��<t��<�?�<0��<���<�U�<��<�<�r�<6��<,�<��<���<�	�<�;�<�a�<R|�<��<@��< ��<'��<!��<t
�<\@�<R��<���<��<s�<���<��<W<�<�]�< i�<�[�<�6�<���<���<�F�<u��<�Q�<|��<�%�<�{�<���<� �<�0�<�V�<�t�<���<;��<��<K��<�<m��<��<�V�<��<�֮<��<�)�<Cͧ<�r�<; �<k٠<���<kz�<3d�<Z]�<c�<\q�<���<��<j��<���<���<Î�<%t�<TQ�<�(�<��<g�{<jAw<u�r<q�n<,j<��e<Cma<Y]<��X<VT<tP<u�K<�iG<�C<k�><zm:<�5<�v1<��,<�*(<l#<	�<^�<�0<�<�<��<�<_��;��;k�;m��;���;e�;L��;)%�;���;k˺;��;�3�;�k�;���;��;���;2_�;�y|;Ӌn;�`;A�S;��F;��:;�.;�m#;|�;(6;+5;���:���:,��:N1�:��:z��:���:0(f:�lD:��$:��:_��9i�9���9�-@9��9�8ǯ7��F������D�����ߌ��b?ʹ�M���h��.2��AE�!X�6�j���}��J�����8��������N�����z�ɺ �ӺͿݺrp� ������c��������ZD!�)�'�ay-�	�2�U�7�K�;�j�?��:C�LrF�L�I�(�L�
6P���S��W�.n\��-a��-f�Yk��p�7�u��{�#������8I���ۇ��q����6���.��/����?���  �  ��=W�=�B=��=?�=,=N�=�W=�� =�v = =�5�<�h�<9��<���<Dd�<���<�_�<8��<"��<s�<t��<y=�<e��<U8�<_��<;	�<f�<��<s�<Cn�<���<x"�<�~�<���<�8�<���<���<�P�<%��<��<aq�<���<�,�<���<���<��<t?�<�e�<��<���<���<<��<���<E��<��<�H�<}��<���<'�<iy�<{��<{�<Q@�<wa�<�k�<�]�<�7�<���<6��<"E�<���<�M�<o��<��<'u�<���<|��<*�<�P�<�o�<��<���<ç�<孻<q��<❷<#��<�Y�<,!�<�ڮ<ˈ�<�/�<�ӧ<7z�<$(�<��<��<���<Zl�<e�<j�<�w�<��<���<���<��<\��<␈<xu�<�Q�<(�<��<ݗ{<a9w<(�r<E}n<�j<�e<�_a<� ]<��X<�MT<L�O<��K<5hG<�C<r�><+q:<�6<.}1<P�,<T3(<�v#<1�< �<"@<��<%<"�<�<d
�;^-�;���;��;ՙ�;�0�;��;�2�;b��;�Ӻ;��;�4�;�h�;Y��;��;��;
J�;�I|;Xn;l�`;R�S;(�F;�v:;�.;xZ#;�;@4;t:;t�:&�:�*�:Il�:O©:B�:N�:h�f:�RE:��%:h�:Z�9ъ�9�9�D9��9v�8�5�70oԷ|*����� C�P.���(��sʹ�`�f��]8�1�2���E�s�X�'�k���~�����o'�����8��rq��z����ɺe�Ӻ,�ݺ�J�*��F����A����Ҫ��n�_	!�KV'��6-�ە2��i7�Y�;�D�?�mC�bAF��jI�c�L�P���S�E�W��]\��#a�Y+f��]k���p��u��5{��7���΂�`c�����%���� ��6����>���Ĕ��F���  �  �=��=D=v�=ӑ=�0=��=4^=�� =� =� =pK�<1��<|��<`�<X|�<���<�t�<h�<-��<7+�<���<�G�<���<?�<(��<��< f�<ֻ�<��<@d�<U��<��<�l�<Q��<%�<���<���<tB�<���<g�<�l�<T��<�-�<N��<���<_�<"I�<6q�<���<���<���<���< ��<� �<H+�<8a�<��<��<m;�<���<���<2�<�K�<�j�<Es�<�c�<d;�<���<d��<@�<2��<�A�<k��<%�<�a�<��<���<��<�?�<:a�<�|�<ђ�<@��<���<Ϭ�<���<���<Pa�<�*�<S�<̖�<�?�<;�<���<�>�<���<�<?��<ڃ�<{�<5~�<���<Ԙ�<4��<��<���<��<���<�x�<�R�<&�<��<&�{<� w<ռr<Zn<G�i<��e<�8a<��\<(�X<�3T<��O<�K<QbG<�C<��><�z:<�6<ю1<��,<=M(<�#<u�<�<l<��<�V<x�<��<�h�;n��;{��;kM�;?��;<f�;K��;zX�;���;�;��;I7�;�^�;���;z�;h�;��;��{;s�m;/)`;��R;�CF;�:;�O.;�#;/l;,;�H;tQ�:�g�:y��:7�:���:,"�:A�:'?i:��G:��(:�:�>�9߰�9��9�`O9��9��8��8'7���H��1��O!?�դ��W%���ɹ���5��0 � 4��G�?�Z�Mn�r���!�J������0ȥ� ߮��᷺P���LʺEtӺq[ݺ���!���`���p�B$�&��	a ��&�w,�)�1���6�#�:�7�>�@dB�t�E���H�H=L���O���S�g�W�&2\��	a�)%f�Cok�p�p��8v�`�{��s���������\F���؊�"g����p���锻�]���  �  ��=G�=�E=��=�=7=��=�g=�� =� =,  ==m�<���<���<>�<J��<��<��<$ �<��<WA�<���<KW�<~��<vH�<>��<;�<yd�<���<��<�S�<���<Y��<O�<���<�<-d�<��<�*�<ȑ�<���<3d�<���<�.�<ԉ�<���<��<W�<`��<C��<���<���<��<��<&�<�Q�<���<^��<��<[�<���<���<�-�<�\�<�x�<~�<k�<b?�<2��<K��<�6�< ��<R.�<���<:��<�A�<}��<���<L��<}#�<aI�<j�<���<��<2��<���<��<Ɛ�<el�<�8�<���<���<�X�<��<@��<b�<"�</�<���<Ҩ�<~��<o��<*��<���<���<���<���<��<P��<!}�<�R�<�!�<�<�h{<��v<��r<@ n<:�i<�Ve<�`<��\<EQX<�T<��O<p�K<�VG<>C<#�><��:<#6<U�1<�-<t(<��#<N<�X<��<3<��<�K<|<���;��;|R�;��;6�;���;�,�;ŏ�;\��;��;�#�;�5�;�J�;do�;߯�;`�;`��;\�z;S�l;1_;R;�kE;�O9;h�-;�";�.;�;TT;:��:��:h�:��:���:�r�:��:��l:��K:��,:�i:���9�_�9v�9��`9?�9_{�8��48���3����c���X9�� }��颹�_ɹ-h�1�l�!�dP6�݉J�4c^���q�<���<닺�*��v@��>-����
����M��c%ʺSRӺH ݺ�Q�^�'*��HL����Y�}���Z�4�%��H+�y�0�rt5���9��=�)mA���D�4H���K�L9O��S�p[W�a�[���`�P&f�x�k��q�,�v��7|�׀� ���^,��{ƈ�PV��ۍ��T��#Ò�'��b����  �  ��=��=�F=�=�=V>=�=�s=	=�� =D3 =��<��<I�<Zo�<���<HC�<���<<E�<��<P\�<���<�h�<��<�Q�<ҵ�<8�<)`�<~��<���<�<�<��<��<k'�<�~�<���<:;�<���<Q
�<�w�<S��<6W�<���<O-�<u��<|��<5+�<�f�<i��<���<^��<���<��<�/�<U�<y��<���<���<;�<��<���<b�<bF�<�p�< ��<D��<r�<TB�<#��<���<-)�<���<'�<9t�<~��<��<
[�<r��<?��<���<)�<-P�<Hr�<_��<x��<M��<���<M��<x�<�H�<7�<Ŭ<-w�<�&�<�ץ<쎣<�N�<M�<n�<�ך<�Ș<�Ė<~ǔ<�͒<�Ӑ<�Վ<Ќ<t��<̥�<C��<�P�<��<��<?{<��v<�Gr<��m<aei<S e<E�`<wR\<]X<��S<~�O<?nK<KCG<WC<��><%�:<�66<W�1<5<-<O�(<G�#<8O<̥<\<�{<�<��<�w<�\ <
��;��;%A�;��;v�;�z�;���;'�;y$�;.�; +�;8(�;�2�;�X�;v��;� �;�y;�k;�];t�P;�JD;BW8;8�,;0$";6�;�;�P;���:Ex�:4.�:��:��:��:5��:<4q:��P:�2:aX:�7�9o��9���9AEw9u49R�8j�q88Tl6kX����?3�3y�]ߡ�D�ɹ���p���'$��}9�C}N�P�b��v��)������C����}�����gp��߳������?tʺ�KӺo�ܺl��*�����0��]�
�J]�����$���)��/�G�3�`_8��q<�{7@���C�'OG�&�J���N���R��W�3�[���`�Q:f���k�5�q�FVw�}� ]��i ��5҆��p�����9v��,ݐ�4��~��×��  �   �=`�=F=�=h�=E=Q�=o=�=�� =oH =���<u�<�Q�<T��<H	�<�v�<���<&n�<���<�x�<g��<@z�<W��<�Y�<���<��<X�<ߜ�<*��</�<|b�<(��<���<L�<q��<
�<\s�<���<W�<!��<uE�<��<m(�<��<��<Y5�<�u�<���<���<I��<~�<�<�<Fa�<i��<���<	��<,�<�l�<���<���<j-�<`�<���<���<ђ�<�v�<B�<X��<ҏ�<j�<G��<_��<bK�<���<���<�%�<lb�<֚�<���<��<�/�<bY�<�|�<���<>��<䩷<���<"��<�W�<� �<�߬<'��<N�<��<���<��< R�<�)�<��<��<'�<��<#�<!�<}�<�ތ<_ʊ<�<*��<1K�<��<n�<m	{<!}v<R�q<{um<� i<��d<�>`<�[<:�W<��S<�aO<�CK< 'G<�C<[�><^�:<�F6<�1<a`-<u�(</7$<�<��<�h<8�<�x<O#	<A�<�� <�;��;
��;(#�;�x�;���;4�;�+�;g7�;�+�;�;���;h�;�;0�;z{�;6x;X�i;�Y\;�RO;j�B;�&7;8�+;�d!;�J;֘;r2;K�:���:���:T��:h1�:۫�:/��:{v:AyV:��8:H:8�:���9�x�9�7�9{�J98�	9<��8ޏ�7�.��wո��-���u�������ʹ�}�����!3'��u=�TS�*�h��}��Y��๑�&����6��Le��bR��~��8�º1 ˺�|Ӻ��ܺ>N�F���
��F���
��L�E��D��"��(�R-��22�6�6���:�1�>�ǥB�gZF�#J��N�%7R���V�q�[�?�`�kf��7l��+r�K-x�U%~�� ���ل�?����=��;Ō�u1��v���ݿ���앻����  �  �==eC=�=�=J=4�=l�=c&=�� =�] =<��<�=�<���<���<=B�<��<��<���<!�<��<��<���<'��<�]�<b��<�<vK�<r��<���<���<�8�<z�<���</�<�n�<��<�@�<N��<x1�<��<�.�<l��<6�<C��<���<�;�<���<=��<���<Y�<�A�<j�<��<���<���<�)�<�c�<���<���<��<�L�<%x�<��<��<Ę�<�w�<q=�<(��<'�<���<l�<k��<I�<:g�<:��<���<�'�<�b�<���<���<7
�<�;�<If�<��<՝�< ��<��<���<�c�<3�<���<���<�u�<4�<���<a��<<��<�c�<�C�<G,�<z�<G�<x�<��<���<1�<�Њ<5��< |�</A�<2��<�e<?�z<�.v<ߘq<{m<L�h<�%d<��_<�[<�VW<�4S<�O<�K<� G<L�B<��><��:<8O6<��1<;-<�(<�p$<r�<�R<	�<�T<�<ܚ	<�]<�5<�F�;1G�;f�;��;���;�
�;-2�;�C�;�:�;@�;g�;ˮ�;��;Uh�;,z�;1;�v;Lh;ƢZ;��M;ucA;��5;��*;� ;��;w%;��;���:n	�:�U�:I��:%Y�:<8�:3��:��z:�-\:,?:�$:��
:ED�9��9|&�9ѥa9#�9��8�p�7Bw	��ȸK*���t�[��t�̹�4��
���*�mB��X�J�n��끺<����;������A��
�������Լ�35ĺ�˺��Ӻ�ܺm�DL�s.��gQ�V=	��@��@��#��� �)O&�,�+�pe0��5��]9��=��A��mE��gI��M�~�Q�I�V�:�[��a�h�f���l���r��*y��^�p���&����u������������9>���_��o��[w���  �  >�=	�=�>=��=�=�L=��=��=3=� =r =" =r�<���<&�<Ey�<_��<4L�<i��<d4�<���<�!�<��<���<�\�<���<7��<�:�<br�<���<���<��<�G�<Ƌ�<o��<�4�<���<h�<T��<!	�<���<��<��<��<D��<���<>�<)��<���<<�<5�<,e�<���<���<?��<�+�<�a�<l��<(��<��<E;�<�h�<���<���<%��<M��<�s�<~4�<���<�j�<|��<�I�<���<���<�0�<�p�<5��<_��<�(�<Ig�<c��<���<p�<)L�<Pt�<'��<���<���<���<�k�<�A�<R�<�ժ<ؚ�<3`�<�'�<��<�ğ<���<�x�<i\�<)F�<�4�<c&�<��<��<[�<nҊ<���<�s�<�2�<��<�.<��z<��u<�7q<��l<�h<�c<�Y_<�[<��V<�R<%�N<~�J<w�F<F�B<D�><a�:<{N6<G�1<��-<d!)<ģ$<�" <i�<�,<��<�_<�
<��<��<Q�;���;���;� �;��;8<�;�L�;NI�;�+�;���;1��;8Z�;.�;�ڑ;�Љ;y �;�t;H�f;��X;�K;*�?;�a4;~�);J�;��; �;f�;�j�:|��:��:�E�:@�:&��:�N�:_:x�a:tVE:��*:�:�f�9�9'��9Jmw9.�/9�p�8)� 8��ط����(�\v��5���Ϲ��������.�x G�&�^�-Pu�kn��]���#ژ��y��Km��.ذ��㷺�����źc�̺
�Ժ�ݺj.�X����]��ۅ� M������1C�;�$�!�)��.�]3�@�7�"8<�4q@���D�;�H��"M�گQ�҇V�ƺ[�~Ka��5g��gm���s��@z��V���y��~��NZ��%	��U����ِ����$
��.����蘻�  �  ��=�z= 8=y�=B�=�M=��=K�=U==,� =Ã =) =��<���<^M�<��<x�<�t�<,��<�N�<���<�-�<���<��<�W�<%��<��<f'�<�Y�<���<���<s��<�<�V�<��<���<�d�<��<SY�<?��<<m�<Z��<P��<B�<�v�<���<<�<w��<���<��<L�<���<��<���<N'�<'^�<���<���<?��<�-�<Z�<��<~��<���<��<ʗ�<Pl�<%(�<=��<�S�<���<�&�<xw�<:��<S��<F8�<t�<[��<:��<3�<w�<���<���<�0�<[^�<a�<���<���<ψ�<ko�<XK�<4�<L�<亨<L��<�T�<�$�<���<�͝<h��<e��<�j�<UR�<<�<�'�<g�<P�<Њ<���<�g�<�!�<Jҁ<��~<	?z<�u<��p<i9l<�g<�>c<��^<ѰZ<;�V<�R<��N<H�J<��F<�B<A�><�y:<�E6<m�1< �-<<)<	�$<�[ <�<�<�<w�<"x
<V5<��<خ�;�y�;�]�;�T�;�W�;�[�;�V�;U>�;�;�Ĳ;rf�;���;Y��;oM�;�)�;OC�;�Us;^�d;�*W;�KJ;U@>;��2; p(;�};};��;';���:҇�:�s�:.��:�۰:��:7Ȑ:㞁:BOf:��J:k�0:O:�:�C�9_��9�S�9��?9�s�8��A8�V��F���9�)�m<y�H𦹁�ӹܓ���3� �K�	Bd��{�Sψ������T��:Ϥ�M�������t?��[���OHǺ!+κ;�պ��ݺ>�溂�@C��Ew����=����~�����#��"(��-�b�1���6�|;�ډ?�y�C�^]H��L�y�Q�r�V�!�[��a�>�g�	n���t�Y{�����m6��M���5��錻�d��z������������_���  �  �=�q=�0=d�="�=�L=5�=��=E=:� =� =J: =��<��<�w�<8��<�3�<��<]��<~c�<���<�5�<ߚ�<.��<�P�<��<���<�<�A�<�i�<���<x��<���<�'�<r�<���<�4�<k��<F0�<���<N�<3��<�k�<E��<�i�<���<$7�<M��<(��<�<�]�<؛�<���<��<XO�<B��<���<���<!�<�L�<�r�<ȑ�<���<���<���<j��<�b�<��<l��<�=�<���<j�<�Q�<Ғ�<���<��<�@�<[~�<��<��<�M�<$��< پ<8�<�H�<n�<���<���<���<�o�<FQ�<v+�<D�<�Ԩ<>��<z�<�M�<"�<��<Л<���<���<�i�<`M�<2�<�<��<�ʊ<c��<SZ�<f�<.��<��~<~�y<?=u<��p<�k<�Mg<��b<M�^<�RZ<�:V<b9R<�GN<�]J<�rF<�~B<B{><Dd:<C86<��1<Y�-<0N)<=�$<�� <1&<$�<>o<<��
<��<�N<�9�;��;I��;��;P~�;�k�;OR�;�(�;��;ˎ�;u�;¤�;�,�;�ʐ;���;J��;S�q;,_c;H�U;��H;��<;�1;W';��;�?;�L;��;0�:b�:�0�:)��:�8�:7L�:��:D*�:@-j:chO:~�5:�:rj:*n�9��9x+�9�L9�y 9��Y8����7����+�7p}�G	��zع�.��C�-�6�]P�Ti�ę��6ɋ�p��dd�������A������i��W�ºb�ȺnhϺ�ֺ�c޺����F�)��>�������4�wy�ũ�5�!�Y�&��+��0��s5�>-:���>�WoC��H��L���Q���V��G\�Eb�aQh���n���u��[|�_���oބ�j��8�������&��&c���j���I�����bΙ��  �  e�=�i=j*=l�=Κ=,K=��=��=IJ=� =�� =
G =4��<�=�<���<M��<P�<��<�<�q�<��<�9�<Ț�<9��<uI�<p��<X��<o�<�-�<CR�<5u�<d��<Z��<�<�K�<��<��<׈�<��<ҟ�<�4�<���<�Y�<v��<�]�<���<�1�<]��<`��<$�<�i�<0��<��<W/�<\m�<��<c��<"�<|<�<lc�<B��<���<Ю�<ʳ�<���<���<wY�<��<��<�*�<O��<c��<�3�<7q�<��<���<��<UV�<`��<t��<�,�<�w�<ſ�<N �<U6�<�^�<Zx�<���<~�<n�<T�<V3�<Z�<,�<⾦<ؕ�<=l�<B�<��<��<�ę<T��<[z�<�X�<e8�<��<~�<(Ŋ<J��<N�<>�<u��<^�~<|�y<Nu<�Ap<H�k<� g<��b<�9^<�Z<�U<d�Q<vN</J<�JF<�]B<-`><]O:<*6<��1<��-<�X)<%<� <�P<&�<֪<�\<�<��<�<H��;UA�;C��;���;��;�p�;�G�;��;1ú;�]�;��;Y�;LӘ;�a�;��;Q�;&�p;`4b;�}T;ڰG;��;;��0;u&;P�;n�;�
;�";L�:w��:`��:]x�:�c�:x¡:���:rE�:�m:��R:ŵ9:ŝ!:�j
:N�9¼9+��9c%U9u�9�i8����`���L.�ր�w�����۹�g�����9���S�%Zm�΂�W"���|���ˡ�����k�����'��tĺʺ�xк�k׺]ߺx�V��Y2�� �BD�yr���������� �]�%�{�*��/��4�q�9�fQ>��C���G���L���Q�W�U�\�n�b�M�h�Hio�#=v�o,}�	���c�����H���I����������h� Ö��y��)���  �  �=od=�%=��==�=�I=u�=�=NM=�� =٢ =�N =���<0Q�<ʫ�<N�<[a�<g��<�<�z�<O��<�;�<ܙ�<���<�C�<���<���<&��</ �<�B�<Zc�<`��<^��<���<K3�<X��<��<"r�<���<���<'$�<4��<�M�<A��<�U�<r��<0-�<J��<���<�'�<�p�<���<���<�?�<��<c��<���<"�<�L�<6q�<���<K��<���<^��<Y��<��<�R�<7�<D��<��<e��<!��<~ �<�[�<���<���<5��<�<�<ʀ�<M��<S�<�d�<﮾<��<�)�<�T�<�o�<	|�<$z�<Al�<'U�<�7�<6�<p�<.ͦ<¦�<�~�<�U�<+�<���<�ԙ<���<s��<�_�<�;�</�<7�<���<���<�E�<���<���<�u~<<�y<��t<�p<�ek<�f<�Zb<�^<��Y<�U<y�Q<��M<�J<10F<GB<�M><�@:<K6<��1<��-<�])<@%<M� <�j<�<(�<�<f:<O�<(�<��;�t�;q�;=��;\��;�p�;�=�;|��;���;J;�;ͷ�;�&�;���;7�;P·;!�;�p;lva;)�S;a�F;�;;0;��%;�H;I*;2c
;��;C��:N!�:��:D\�:�q�:
�:}'�:s�:��n:��T:/<:$:u�:���9���9xy�9ТZ9)�
9fhq8�����j��}`0��d��$����%޹����!�[�;�2EV� �o��6��i���.��S��,����β��K���H��ź]�ʺ�0Ѻغ)�ߺ������|E�������/�\>��C�@�28 �0%�V,*�e*/��%4�Z9��>���B�"�G��L�]�Q�P(W�-�\�&�b�B"i���o�:�v���}�OV����� ��x���g ���Q���G��!��b����e���  �  ě=yb=Q$=��=F�=2I=_�=H�=5N=?� =� =uQ =��<�W�<���<��<[g�<v��<�<Q}�<���<T<�<���<���<�A�<X��<���<$��<��<>=�<2]�<l��<���<s��<�*�<҃�<���<,j�<o��<���<n�<e��<SI�<~��<�R�<��<}+�<���<��<�(�<!s�<#��<B�<ME�<��<��<���<�(�<�R�<�u�<x��<���<���<~��<���<$��<BP�<.�<\��<��<q��<7��<��<T�<R��<J��<_��<4�<Ox�<7��<��<-^�<%��<��<�%�<�P�<�l�<�y�<�x�<�k�<fU�<�8�<��<(��<Ҧ<���<`��<�\�<�1�<�<eڙ<�<���<�a�<�<�<>�<]�<Ͼ�<V��<�B�<�<���<�k~<w�y<N�t<�p<�Uk<3�f<�Ib<��]<f�Y<��U<��Q<}�M<>J<*'F<�>B<�F><P;:<>6<��1<<�-<�_)<�%<c� <s<�&<��<��<dH<��<��<R��;���;�(�;{��;ȣ�;Xp�;�9�;c��;7��;�.�;Ҩ�;��;��;��;n��;�F;l�o;�4a;�{S;��F;��:;��/;��%;�;6;�B
;�;x��:��:߆�:R�:�u�:��:gL�:c)�:�Uo:�U:��<:�$:(�:dM�9�a�92��9�o\9O�9�s8������5.1���y����߹�j�DF"�˰<�GW���p�Q���2#��R����ڣ�����J����������gźE;˺vqѺ�=غK�ߺ���#���L��>�������0���r ���$��)���.��3���8���=���B���G�~�L��Q�97W��\�v�b�NAi�	�o���v���}��p���օ�C��I���͎�B���q���e��-,��dט�Vz���  �  �=od=�%=��==�=�I=u�=�=NM=�� =٢ =�N =���<0Q�<ʫ�<N�<[a�<g��<�<�z�<O��<�;�<ܙ�<���<�C�<���<���<&��</ �<�B�<Zc�<`��<^��<���<K3�<X��<��<"r�<���<���<'$�<4��<�M�<A��<�U�<r��<0-�<J��<���<�'�<�p�<���<���<�?�<��<c��<���<"�<�L�<6q�<���<K��<���<^��<Y��<��<�R�<7�<E��<��<e��<!��< �<�[�<���<���<6��<�<�<ˀ�<N��<T�<�d�<﮾<��<�)�<�T�<�o�<
|�<%z�<Bl�<(U�<�7�<7�<p�<.ͦ<¦�<�~�<�U�<+�<���<�ԙ<���<s��<�_�<�;�<.�<6�<���<���<�E�<���<���<�u~<;�y<��t<�p<�ek<�f<�Zb<�^<��Y<�U<z�Q<��M<�J<20F<GB<�M><�@:<M6<��1<��-<�])<A%<M� <�j<�<)�<�<f:<O�<(�<��;�t�;o�;;��;Y��;�p�;�=�;y��;���;G;�;ʷ�;�&�;���;4�;N·;�;�p;iva;&�S;^�F;�;;0;��%;�H;H*;1c
;��;B��:M!�:��:D\�:�q�:	�:}'�:s�:��n:��T:/<:$:u�:���9���9xy�9ТZ9)�
9fhq8�����j��}`0��d��$����%޹����!�[�;�2EV� �o��6��i���.��S��,����β��K���H��ź]�ʺ�0Ѻغ)�ߺ������|E�������/�\>��C�@�28 �0%�V,*�e*/��%4�Z9��>���B�"�G��L�]�Q�P(W�-�\�&�b�B"i���o�:�v���}�OV����� ��x���g ���Q���G��!��b����e���  �  e�=�i=j*=l�=Κ=,K=��=��=IJ=� =�� =
G =4��<�=�<���<M��<P�<��<�<�q�<��<�9�<Ț�<9��<uI�<p��<X��<o�<�-�<CR�<5u�<d��<Z��<�<�K�<��<��<׈�<��<ҟ�<�4�<���<�Y�<v��<�]�<���<�1�<]��<`��<$�<�i�<0��<��<W/�<\m�<��<c��<"�<|<�<lc�<B��<���<Ю�<ʳ�<���<���<wY�<��<��<�*�<P��<c��<�3�<7q�<��<���<��<VV�<`��<u��<�,�<�w�<ƿ�<P �<W6�<�^�<[x�<���<�~�<n�<T�<W3�<[�<-�<⾦<ؕ�<=l�<B�<��<��<�ę<S��<[z�<�X�<d8�<��<|�<'Ŋ<H��<N�<<�<t��<\�~<z�y<Lu<�Ap<G�k<� g<��b<�9^<�Z<�U<f�Q<xN</J<�JF<�]B</`><_O:<*6<��1<��-<�X)<%<!� <�P<'�<֪<�\<�<��<�<F��;SA�;@��;���;��;�p�;�G�;�;,ú;�]�;��;Y�;GӘ;�a�;��;M�;�p;Y4b;�}T;հG;��;;��0;u&;N�;l�;�
;�";L�:u��:_��:\x�:�c�:w¡:���:rE�:�m:��R:ŵ9:ŝ!:�j
:N�9¼9+��9c%U9u�9�i8����`���L.�ր�w�����۹�g�����9���S�%Zm�΂�W"���|���ˡ�����k�����'��tĺʺ�xк�k׺]ߺx�V��Y2�� �BD�yr���������� �]�%�{�*��/��4�q�9�fQ>��C���G���L���Q�W�U�\�n�b�M�h�Hio�#=v�o,}�	���c�����H���I����������h� Ö��y��)���  �  �=�q=�0=d�="�=�L=5�=��=E=:� =� =J: =��<��<�w�<8��<�3�<��<]��<~c�<���<�5�<ߚ�<.��<�P�<��<���<�<�A�<�i�<���<x��<���<�'�<r�<���<�4�<k��<F0�<���<N�<3��<�k�<E��<�i�<���<$7�<M��<(��<�<�]�<؛�<���<��<XO�<B��<���<���<!�<�L�<�r�<ȑ�<���<���<���<j��<�b�<��<m��<�=�<���<j�<�Q�<Ӓ�<���<��<�@�<\~�<��<��<�M�<&��<"پ<:�<�H�<n�<���<���<���<�o�<HQ�<x+�<E�<�Ԩ<?��<z�<�M�<"�<��<Л<���<���<�i�<_M�< 2�<�<��<�ʊ<a��<QZ�<e�<,��<��~<|�y<==u<��p<�k<�Mg<��b<N�^<�RZ<�:V<d9R<�GN<�]J<�rF<�~B<E{><Gd:<F86<��1<\�-<3N)<@�$<�� <3&<&�<?o<<��
<��<�N<�9�;��;D��;��;I~�;�k�;GR�;�(�;��;Î�;m�;���;�,�;�ʐ;���;D��;I�q;#_c;@�U;��H;��<;�1;W';��;�?;�L;��;-�:`�:�0�:(��:�8�:7L�:��:D*�:@-j:chO:~�5:�:rj:*n�9��9x+�9�L9�y 9��Y8����7����+�7p}�G	��zع�.��C�-�6�]P�Ti�ę��6ɋ�p��dd�������A������i��W�ºb�ȺnhϺ�ֺ�c޺����F�)��>�������4�wy�ũ�5�!�Y�&��+��0��s5�>-:���>�WoC��H��L���Q���V��G\�Eb�aQh���n���u��[|�_���oބ�j��8�������&��&c���j���I�����bΙ��  �  ��=�z= 8=y�=B�=�M=��=K�=U==,� =Ã =) =��<���<^M�<��<x�<�t�<,��<�N�<���<�-�<���<��<�W�<%��<��<f'�<�Y�<���<���<s��<�<�V�<��<���<�d�<��<SY�<?��<<m�<Z��<P��<B�<�v�<���<<�<w��<���<��<L�<���<��<���<N'�<'^�<���<���<?��<�-�<Z�<��<~��<���<��<ʗ�<Pl�<%(�<>��<�S�<���<�&�<yw�<;��<T��<G8�<	t�<\��<<��<�3�<w�<ù�<���<�0�<]^�<d�<Ñ�<���<ш�<mo�<ZK�<6�<M�<庨<M��<�T�<�$�<���<�͝<g��<d��<�j�<TR�<}<�<'�<e�<M�<Њ<���<�g�<�!�<Hҁ<��~<?z<�u<��p<g9l<�g<�>c<��^<ҰZ<=�V<�R<��N<K�J<��F<
�B<E�><�y:<�E6<q�1<$�-<<)<�$<�[ < �<�<�<x�<"x
<U5<��<ծ�;�y�;�]�;�T�;�W�;�[�;�V�;L>�;	�;�Ĳ;if�;���;Q��;gM�;�)�;HC�;�Us;S�d;�*W;�KJ;N@>;��2;p(;�};y;��;%;���:χ�:�s�:,��:�۰:��:6Ȑ:㞁:AOf:��J:k�0:O:�:�C�9^��9�S�9��?9�s�8��A8�V��F���9�)�m<y�H𦹁�ӹܓ���3� �K�	Bd��{�Sψ������T��:Ϥ�M�������t?��[���OHǺ!+κ;�պ��ݺ>�溂�@C��Ew����=����~�����#��"(��-�b�1���6�|;�ډ?�y�C�^]H��L�y�Q�r�V�!�[��a�>�g�	n���t�Y{�����m6��M���5��錻�d��z������������_���  �  >�=	�=�>=��=�=�L=��=��=3=� =r =" =r�<���<&�<Ey�<_��<4L�<i��<d4�<���<�!�<��<���<�\�<���<7��<�:�<br�<���<���<��<�G�<Ƌ�<o��<�4�<���<h�<T��<!	�<���<��<��<��<D��<���<>�<)��<���<<�<5�<,e�<���<���<?��<�+�<�a�<l��<(��<��<E;�<�h�<���<���<%��<M��<�s�<~4�<���<�j�<|��<�I�<���<���<�0�<�p�<6��<`��<�(�<Kg�<e��<���<s�<,L�<Rt�<*��<���<ě�<���<�k�<�A�<T�<�ժ<ٚ�<5`�<�'�<��<�ğ<���<�x�<h\�<'F�<�4�<a&�<�<��<Y�<lҊ<���<�s�<�2�<��<�.<�z<��u<�7q<��l<�h<�c<�Y_<�[<��V<�R<(�N<��J<{�F<J�B<I�><f�:<�N6<L�1<��-<i!)<ȣ$<# <l�<�,<��<�_<�
<��<��<M�;���;���;� �;��;/<�;�L�;DI�;�+�;���;'��;.Z�;%�;�ڑ;�Љ;r �;�t;<�f;��X;�K;"�?;�a4;y�);F�;��;�;c�;�j�:y��: ��:�E�:@�:%��:�N�:_:w�a:sVE:��*:�:�f�9�9'��9Jmw9.�/9�p�8)� 8��ط����(�\v��5���Ϲ��������.�x G�&�^�-Pu�kn��]���#ژ��y��Km��.ذ��㷺�����źc�̺
�Ժ�ݺj.�X����]��ۅ� M������1C�;�$�!�)��.�]3�@�7�"8<�4q@���D�;�H��"M�گQ�҇V�ƺ[�~Ka��5g��gm���s��@z��V���y��~��NZ��%	��U����ِ����$
��.����蘻�  �  �==eC=�=�=J=4�=l�=c&=�� =�] =<��<�=�<���<���<=B�<��<��<���<!�<��<��<���<'��<�]�<b��<�<vK�<r��<���<���<�8�<z�<���</�<�n�<��<�@�<N��<x1�<��<�.�<l��<6�<C��<���<�;�<���<=��<���<Y�<�A�<j�<��<���<���<�)�<�c�<���<���<��<�L�<%x�<��<��<Ę�<�w�<q=�<(��<'�<���<l�<l��<J�<;g�<;��<���<�'�<�b�<���<���<9
�<�;�<Lf�<��<ם�<��<��<���<�c�<3�<���<���<�u�<4�<���<a��<<��<�c�<�C�<F,�<y�<E�<v�<��<���</�<�Њ<2��<�{�<-A�<0��<�e<<�z<�.v<ܘq<ym<K�h<�%d<��_<�[<�VW<�4S<�O<�K<� G<P�B<��><��:<=O6<��1<?-<#�(<�p$<u�<�R<�<�T<�<ܚ	<�]<�5<�F�;+G�;�e�;ܘ�;���;�
�;#2�;�C�;�:�;5�;\�;���;��;Kh�;$z�;);��v;Lh;��Z;��M;mcA;��5;��*; ;��;t%;��;���:k	�:�U�:G��:#Y�:;8�:3��:��z:�-\:,?:�$:��
:DD�9��9|&�9ѥa9#�9��8�p�7Bw	��ȸK*���t�[��t�̹�4��
���*�mB��X�J�n��끺<����;������A��
�������Լ�35ĺ�˺��Ӻ�ܺm�DL�s.��gQ�V=	��@��@��#��� �)O&�,�+�pe0��5��]9��=��A��mE��gI��M�~�Q�I�V�:�[��a�h�f���l���r��*y��^�p���&����u������������9>���_��o��[w���  �   �=`�=F=�=h�=E=Q�=o=�=�� =oH =���<u�<�Q�<T��<H	�<�v�<���<&n�<���<�x�<g��<@z�<W��<�Y�<���<��<X�<ߜ�<*��</�<|b�<(��<���<L�<q��<
�<\s�<���<W�<!��<uE�<��<m(�<��<��<Y5�<�u�<���<���<I��<~�<�<�<Fa�<i��<���<	��<,�<�l�<���<���<j-�<`�<���<���<ђ�<�v�<B�<X��<ӏ�<k�<G��<`��<cK�<���<���<�%�<mb�<ؚ�<���<��<�/�<eY�<�|�<���<A��<穷<���<$��<�W�<� �<�߬<)��<N�<��<���<��< R�<�)�<��<��<%�<��<!�<�<{�<�ތ<\ʊ<�<'��</K�<��<j�<j	{<}v<P�q<yum<� i<��d<�>`<�[<<�W<��S<�aO<�CK<'G<�C<`�><c�:<�F6<�1<f`-<y�(<37$<�<��<�h<:�<�x<O#	<@�<�� <�~�;��;��; #�;�x�;���;*�;�+�;\7�;�+�;�;���;_�;�;(�;r{�;6x;L�i;�Y\;�RO;b�B;&7;2�+;�d!;�J;Ә;p2;H�:���:���:S��:g1�:ګ�:.��:zv:AyV:��8:H:7�:���9�x�9�7�9{�J98�	9<��8ޏ�7�.��wո��-���u�������ʹ�}�����!3'��u=�TS�*�h��}��Y��๑�&����6��Le��bR��~��8�º1 ˺�|Ӻ��ܺ>N�F���
��F���
��L�E��D��"��(�R-��22�6�6���:�1�>�ǥB�gZF�#J��N�%7R���V�q�[�?�`�kf��7l��+r�K-x�U%~�� ���ل�?����=��;Ō�u1��v���ݿ���앻����  �  ��=��=�F=�=�=V>=�=�s=	=�� =D3 =��<��<I�<Zo�<���<HC�<���<<E�<��<P\�<���<�h�<��<�Q�<ҵ�<8�<)`�<~��<���<�<�<��<��<k'�<�~�<���<:;�<���<Q
�<�w�<S��<6W�<���<O-�<u��<|��<5+�<�f�<i��<���<^��<���<��<�/�<U�<y��<���<���<;�<��<���<b�<bF�<�p�< ��<D��<r�<TB�<$��<���<-)�<���<(�<:t�<��<��<[�<s��<@��<���<)�</P�<Jr�<a��<z��<O��<���<P��<x�<�H�<9�<Ŭ<.w�<�&�<�ץ<펣<�N�<M�<m�<�ך<�Ș<�Ė<|ǔ<�͒<�Ӑ<�Վ<Ќ<r��<ɥ�<@��<�P�<��<��<�>{<��v<�Gr<��m<aei<S e<F�`<xR\<_X<��S<��O<BnK<NCG<[C<��><*�:<�66<[�1<9<-<S�(<J�#<;O<Υ<^<�{<�<��<�w<�\ <��;z��;A�;���;n�;�z�;���;�;p$�;.�;�*�;/(�;�2�;�X�;o��;� �;צy;�k;�];l�P;�JD;<W8;3�,;,$";3�;�;�P;���:Bx�:2.�:��:��:��:4��:;4q:��P:�2:aX:�7�9n��9���9AEw9u49R�8j�q89Tl6kX����?3�3y�]ߡ�D�ɹ���p���'$��}9�C}N�P�b��v��)������C����}�����gp��߳������?tʺ�KӺo�ܺl��*�����0��]�
�J]�����$���)��/�G�3�`_8��q<�{7@���C�'OG�&�J���N���R��W�3�[���`�Q:f���k�5�q�FVw�}� ]��i ��5҆��p�����9v��,ݐ�4��~��×��  �  ��=G�=�E=��=�=7=��=�g=�� =� =,  ==m�<���<���<>�<J��<��<��<$ �<��<WA�<���<KW�<~��<vH�<>��<;�<yd�<���<��<�S�<���<Y��<O�<���<�<-d�<��<�*�<ȑ�<���<3d�<���<�.�<ԉ�<���<��<W�<`��<C��<���<���<��<��<&�<�Q�<���<^��<��<[�<���<���<�-�<�\�<�x�<~�<k�<b?�<2��<K��<�6�<��<S.�<���<;��<�A�<~��<���<M��<#�<cI�<j�<���<��<3��<���<��<Ȑ�<fl�<�8�<���<���<�X�<��<A��<b�<"�</�<���<Ѩ�<}��<n��<)��<���<���<���<���< ��<N��<}�<�R�<�!�<�<�h{<��v<ފr<? n<9�i<�Ve<�`<��\<FQX<�T<��O<s�K<�VG<AC<&�><��:<#6<Y�1<�-<"t(<��#<P<�X<��<4<��<�K<|<���;��;xR�;
��;6�;���;�,�;���;U��;~�;�#�;�5�;�J�;]o�;ٯ�;Z�;Z��;R�z;J�l;1_;R;�kE;�O9;d�-;�";�.;�;ST;7��:��:h�:��:���:�r�:��:��l:��K:��,:�i:���9�_�9v�9��`9?�9_{�8��48���3����c���X9�� }��颹�_ɹ-h�1�l�!�dP6�݉J�4c^���q�<���<닺�*��v@��>-����
����M��c%ʺSRӺH ݺ�Q�^�'*��HL����Y�}���Z�4�%��H+�y�0�rt5���9��=�)mA���D�4H���K�L9O��S�p[W�a�[���`�P&f�x�k��q�,�v��7|�׀� ���^,��{ƈ�PV��ۍ��T��#Ò�'��b����  �  �=��=D=v�=ӑ=�0=��=4^=�� =� =� =pK�<1��<|��<`�<X|�<���<�t�<h�<-��<7+�<���<�G�<���<?�<(��<��< f�<ֻ�<��<@d�<U��<��<�l�<Q��<%�<���<���<tB�<���<g�<�l�<T��<�-�<N��<���<_�<"I�<6q�<���<���<���<���< ��<� �<H+�<8a�<��<��<m;�<���<���<2�<�K�<�j�<Es�<�c�<d;�<���<d��<	@�<2��<�A�<l��<%�<�a�<��<���<��<�?�<;a�<�|�<Ғ�<A��<���<Ь�<���<�<Ra�<�*�<T�<͖�<�?�<<�<���<�>�<���<�<?��<ك�<{�<4~�<���<Ә�<3��<��<���<��<���<�x�<�R�<&�<��<%�{<� w<Լr<
Zn<F�i<��e<�8a<��\<)�X<�3T<��O<�K<SbG<�C<��><�z:<�6<ӎ1<��,<?M(<!�#<w�<�<l<��<�V<x�<��<�h�;k��;x��;hM�;;��;7f�;F��;uX�;���;�;��;D7�;�^�;���;v�;h�;��;��{;l�m;*)`;��R;�CF;�:;�O.;�#;-l;,;�H;rQ�:�g�:x��:6�:���:+"�:A�:&?i:��G:��(:�:�>�9ް�9��9�`O9��9��8��8'7���H��1��O!?�դ��W%���ɹ���5��0 � 4��G�?�Z�Mn�r���!�J������0ȥ� ߮��᷺P���LʺEtӺq[ݺ���!���`���p�B$�&��	a ��&�w,�)�1���6�#�:�7�>�@dB�t�E���H�H=L���O���S�g�W�&2\��	a�)%f�Cok�p�p��8v�`�{��s���������\F���؊�"g����p���锻�]���  �  ��=W�=�B=��=?�=,=N�=�W=�� =�v = =�5�<�h�<9��<���<Dd�<���<�_�<8��<"��<s�<t��<y=�<e��<U8�<_��<;	�<f�<��<s�<Cn�<���<x"�<�~�<���<�8�<���<���<�P�<%��<��<aq�<���<�,�<���<���<��<t?�<�e�<��<���<���<<��<���<E��<��<�H�<}��<���<'�<iy�<{��<{�<Q@�<wa�<�k�<�]�<�7�<���<6��<"E�<���<�M�<p��<��<'u�<���<|��<*�<�P�<�o�<��<���<ħ�<死<r��<㝷<$��<�Y�<-!�<�ڮ<ˈ�<�/�<�ӧ<7z�<$(�<��<��<���<Zl�<e�<j�<�w�<��<���<���<��<[��<␈<wu�<�Q�<(�<��<ܗ{<`9w<(�r<D}n<�j<߿e<�_a<� ]<��X<�MT<M�O<��K<6hG<�C<t�><,q:<�6<0}1<Q�,<U3(<�v#<2�<!�<"@<��<%<"�<�<c
�;]-�;���;��;ә�;�0�;��;�2�;_��;�Ӻ;��;�4�;�h�;V��;��;��;J�;�I|;Xn;i�`;O�S;&�F;�v:;�.;vZ#;�;?4;t:;s�:%�:�*�:Hl�:N©:B�:N�:h�f:�RE:��%:h�:Z�9ъ�9�9�D9��9v�8�5�70oԷ|*����� C�P.���(��sʹ�`�f��]8�1�2���E�s�X�'�k���~�����o'�����8��rq��z����ɺe�Ӻ,�ݺ�J�*��F����A����Ҫ��n�_	!�KV'��6-�ە2��i7�Y�;�D�?�mC�bAF��jI�c�L�P���S�E�W��]\��#a�Y+f��]k���p��u��5{��7���΂�`c�����%���� ��6����>���Ĕ��F���  �  !�=L�=c2=b�=�~=�=T�=cT=&� =6� =M =.d�<���<���<<�<8��<�
�<4��<��<Ĉ�<L�<���<�<���<���< e�<���<#�<u{�<���<�'�<d~�<���<0.�<>��<���<�:�<K��<1��<�K�<���<��<�[�<���< �<gG�<���<���<!��<`�<F"�<�:�<eS�<�n�<��<9��<��<��<V�<ٓ�<���<k�<7�<3X�<�h�<�f�<(P�<%�<0��<���<�1�<B��<�>�<'��<��<�p�<���<��<E:�<j�<ő�<���<�̾<I�<`�<��<�<-״<-��<2��<�Z�<��<)٩<-��<jN�<��<�֠<ҩ�<'��<br�<rg�<�e�<�i�<�p�<�w�<�z�<9x�<�n�<�\�<{C�<�#�<���<��<�W{<�w<��r<Tn<5�i<Y�e<�Qa<��\<�X<�aT<�P<�K<F�G<�HC<��><��:<�C6<�1<~O-<��(<�($<E�<v�<4h<��<'�<�>	<�<�<T�;�V�;���;�(�;d��;��;���;���;GA�;���;߭;�6�;ܟ�;L$�;$ɏ;���;���;vKu;&�g;l�Z;8GN;�B;�c6;�+;HK ;}�;�;t�;c��:���:�0�:�̸:T��:��:�:�g:"H:�J+:s�:��9�3�9���9C�r9Y�/9�Q�8n�H8��D����w�˴U�땏�����*�ܹKD��;�u*���=��Q���d��Xx�Oх��l��$����������f��\޾�(yȺ�QҺʈܺ2�b�\��#�3g�*��f��R��P$�"�)�xM/��74�;�8�r�<��@�H�D��BH���K�N�O�+�S�a:X�2�\�͢a�/�f�9�k��q��`v�~�{�Jw��[��B����I��mኻ�u�����%��� ��Щ���  �  ��= �=�2=��=�= =��=�U=� =e� =� =�i�<[��<���<(B�<B��<��<���<w�<��<��<���<��<ʍ�<��<f�<!��<�"�<Xz�< ��<-%�<�z�<���<�)�<D��<���<�5�<א�<j��<�H�<_��<]�<[�<հ�<� �<�H�<J��<��<���<�	�<G&�<�?�<�X�<#t�<ה�<M��< ��<� �<�[�<���<A��<k�<D:�<�Z�<+k�<gh�<\Q�<�%�<���<���<10�<��<�;�<6��<\�<�k�<M��<?��<O5�<�e�<��<|��<�ʾ<�޼<��<��<��<tش<���<���<P]�<8 �<:ݩ<ӗ�<�S�<`�<�ܠ<ޯ�<<��<Hx�<m�<�j�<'n�<�t�<�z�<�}�<�z�<Mp�<�]�<�C�<i#�<���<��<;S{<*�v<��r<�Jn<T�i<�e<�Ga<[�\<¥X<�ZT<xP<��K<�G<HC<p�><��:<�F6<_�1<�T-<	�(<>0$<�<��<^s<��<��<:K	<f<�<�-�;�j�;k��;�7�;K��;�&�;���;���;�E�;��;�ݭ;03�;���;=�;ӻ�;���;�t�;�$u;��g;'�Z;�$N;��A;�K6;�+;�A ;��;��;7�;\��:���:�X�:t��:��:�G�:�3�:/�g:��H:8
,:��:b��9 ��9��9�Su9X29"g�83O8�-�s�������U��h��î��~�ܹ�k�}|� �*��^>��R�ݖe�_�x��!��+���Y@��f���y!��*�����e�Ⱥ�OҺ�zܺx�GB����^�3K����o��Y(��"$���)��/� 4�<�8��<��@��qD��#H�@�K�
�O���S��,X���\�C�a�b�f���k�r"q��sv���{�����'���ą�^����������������)�������  �  �=Ć=!3=\�=Ɂ=#=��=�Z=�� =�� =�! =by�<0��<���<�S�<���<L!�<���<T�<K��<��<���<�<]��<�<�h�<���<R!�<�v�<1��<�<�p�<j��<��<�s�<(��<�'�<��<G��<�?�<���<���<�X�<ư�<h�<
L�<'��<g��<��<r�<�1�<�L�<7g�<5��<��<���<���<�1�<�k�<���<g��<��<D�<c�<�q�<m�<~T�<'�<���<
��<M+�<ѵ�<(2�<���<��<�\�<��<���<�&�<UX�<���<e��<�þ<eڼ<o�<��<h�<�۴<ؿ�<9��<�e�<B*�<��<:��<�b�<�$�<J�<���<柜<G��<�|�<$y�<#{�<��<t��<���<뀌<u�<.a�<�E�<#�<1��<��<D{<��v<b�r<0n<}�i<=e<�*a<��\<��X<<FT<�P<{�K<L�G<FC<$�><�:<*O6<��1<�c-<v�(<MF$<�<C<=�<�<z�<�o	<WB<!0<�m�;���;��;e�;^��;F�;���;[�;QR�;{��;lۭ;?'�;���;���;ڔ�;�T�;H@�;�t;LMg;QOZ;��M;��A;6;��*;T  ;��;1�;�;�
�:�F�:��:K��:���:�:��:��i:;�J:11.:¹:�
�9,�9��9��|9h�89�)�83Nc8�.ֶ/돸P�BS��쎹����jzݹ���O�0�+�ػ?���S�Vg��z�d
������&��`��P���B嵺�-���Ⱥ;GҺVܺ������S~�������
��@���]��؞#��C)���.��y3��8�HB<��;@�hD�z�G�ƕK���O� �S�bX���\���a�;�f��k�$Kq��v��|�Z����\������ꘈ�h.��Ͻ���F���ɒ��H��Gŗ��  �  k�=��=�3=3�=��=�'=*�=�a=�� =w� =- =��<���<>�<�o�<4��<x;�<*��<,�<��<�-�<��<�'�<�<��<�k�<��<��<�p�<l��<��<�_�<~��<��<N\�<k��<��<�n�<���<�0�<&��<���<�T�<���<;�<�P�<^��<��<F��<Q"�<GC�<a�<E~�<~��<���<���<��<�L�<&��<��<���<m)�<�R�<o�<�z�<t�<�X�<�(�<��<Y��<�"�<��<�"�<���<��<�D�<��<4��<)�<�B�<Gp�<{��<x��<�Ҽ<5�<��<;�<O�<ǲ<㡰<�q�<e9�<���<*��<>z�<l>�<~	�<�ݞ<���<��<��<�<K��<V��<$��<���<m��<|�<{e�<G�<�!�<f��<��<H,{<k�v<-er<�n<��i<	Oe<b�`<p�\<�eX<�$T<_�O<o�K<�zG<�@C< ?<~�:<3[6<7�1<Az-<_�(<�g$<��<MI<U�<�P<��<�	<�z<-f<���;)��;aJ�;`��;7�;.u�;9��;s �;�b�;L��;�ӭ;-�;a�;�ɖ;�T�;D�;��;h�s;t�f;�Y;bM;�A;�5;F�*;��;��;��;: ;P[�:&��:�c�:�I�:9�:��:)T�:0l:xN:��1:�8:��9���9o�9OD�9�+C9�9q��8�jڴ� ��==�X�P�b���ӵ��o޹���ʭ�m-���A�@V��.j�l�}�p�������]J��5t��n���ۇ�������ȺvHҺ])ܺ��j�#����\��y
�ج�������"��h(�î-��2��17��z;�M�?��lC�CG�4#K��%O�]S�M�W���\�ފa���f��l�ޏq�w�e�|�P��ٲ��rZ�������������7���b
���z��;闻�  �  K�=��=�3=��=H�=�,=��=	j=.=�� =; =A��<}��<�>�<�<J��<�\�<���<WG�<���<`A�<��<P4�<��<��<Zn�<$��<}�<^g�<���<-��<�H�<��<(��<=�<ٕ�<���<�R�<I��<$�<4��<���<�M�<۬�<^�<U�<"��<"��<�	�<j4�<2Y�<�z�<R��<���<��<�<<�<;o�<L��<��<��<e?�<�d�<_}�<���<o{�<�\�<$)�<���<Մ�<
�<1��<4�<�t�<���<9%�<p�<S��<���<}&�<cW�<���<���<�Ǽ<\޺<��<H�<��<�β<��<���<�K�<��<�ԧ<���<_�<7,�<4�<ߜ<9ƚ<ٵ�<���<���<⦒<�<͟�<O��<���<�i�<�G�<,�<��<mv<w
{<@�v<�1r<��m<Xii<�e<o�`<~r\<1X<��S<�O<v�K<�hG<P7C<��><U�:<�g6<�2<p�-<)<�$<C <�<�<��<)9<x�	<�<�<�P�;�q�;^��;���; V�;ɬ�;���;K=�;�r�;i��;�ĭ;��;K.�;V��;p��;Y��;�x�;�s;Ӡe;.�X;�EL;�\@;j�4;`*;��;�{;մ;�.;l��:]F�:G�:�8�:���:���:��:�+p:TR:��5:��:�:N��9���9���9OIP9�A9t{�8=1�6=�t�x%�cdN�����i���๟:�n����/�.E�G�Y���m��ڀ��x���֓������饺 ����m���2���#ɺY_Һhܺ?,���� ��J����	����(�L���!�.Q'���,�y�1�&"6��~:���>�0�B�0�F���J�N�N��	S�#�W��p\��a���f�Xl��q���w��:}�g��>%���Ն��v��\������o���Yb������j���  �  ��=X�=[2=��=�=O1=��=�r=f=+� =�J =���<��<�f�<z��<B�<w��<8��<�e�<���<�V�<��<A�<���<��<6o�<���<��<�Z�<٠�<C��<�,�<�v�<���<��<2p�<(��<
1�<|��<��<!o�<���<�C�<���<g�<X�<��<
��<��<�G�<q�<��< ��<���<

�<�5�<od�<R��<���<���<-�<ZW�<&x�<'��<Y��<��<<_�<�'�<���<Dz�<W�<:��<��<�U�<î�<U��<�H�<��<o��<	�<@9�<�i�<���<���<�Ժ<��<;�<��<�ղ<0��<��<�_�<$*�<��<���< ��<�S�<�)�<��<��<�٘<�̖<pĔ<Z��<ط�<}��<ퟌ<.��<_l�<FF�<o�<)�<�V<2�z<�hv<�q<D�m< i<r�d<Uq`<�+\<�W<��S<ٗO<�sK<PG<�(C<��><��:<r6<2<M�-<�:)<�$<�> <��<�L<��<z�<F
<T< �<���;���;E�;�Y�;��;'��;�$�;�V�;|�;0��;ܫ�;ť;��;�-�;!��;t&�;X�;��q;�|d;*�W;�?K;�v?;W54;�s);G#;�3;l�;
-;���:1��:e��:�0�:��:�
�:Ŀ�:�Nt:űV:��::�� :љ:�a�9>˺9.��9��^9�9�h�8B�l7$^��u �0�L���������Y�0��
��3��H�3�]��yr�?4���ό�|��\�������+�����������ɺ˚Һ��ۺ���9X��N���[�17	��&�x����w� ��&��J+�J=0�J�4�!a9�5�=�"�A���E��J�^GN�z�R�gjW�(_\�4�a��g���l�Grr�KAx��~�7⁻@����h��a��)������|x��}͓�����^���  �  H�=�{=�/=�=�=$5=��=m{=h=ĺ =�Z =��<�A�<ܐ�<��<�D�<���<��<Ȅ�<���<�k�<���<AL�<n��<@�<�m�<��<?�<K�<���<���<��<�R�<���<���<�F�<���<��<w�<b��<�W�<���<�6�<ğ�<� �<�X�<��<��<c&�<=Z�<ƈ�<ϳ�<���<g�<�2�<�_�<���<��<���<��<J�<o�<���<���<%��<Q��<_�<X#�<,��<�l�<|��<�k�<U��<[3�<��<}��<M�<�`�<��<���<��<�L�<D}�<���<�Ǻ<l޸<��<s�<�ڲ<���<B��<.s�<�B�<{�<"ܥ<���<�|�<BT�<�1�<a�<��<��<���<�Ւ<�ɐ<׻�<���<̎�<�l�<>B�<��<�ց<�0<Y�z<3-v<�q<I8m<��h<&nd<r`<�[<ѩW<g�S<�cO<�JK<c1G<C<A�><6�:<'x6<�&2<=�-<C\)<P�$<ou <�<Ė<.5<w�<j�
<Bk<1J<(u�;�s�;��;
��;��;��;.F�;%h�;:|�;���;���;P��;��;]ʕ;��;М�;��~;�p;�:c;L`V;�J;�t>;IY3;��(;ś;��;�Y;;3�:��:r�:��:��:G��:̓�:`�x:�q[:{�?:Z&:�:���9�X�9��9�m9�$9F��8���7~�J�5����K��ގ�[k���i�z/	�K��Ƃ6���L���b��xw�_˅�Uc������fF��L����ٱ�t깺V	º)Yʺ�Ӻ�ܺ��庨��<���4��Д�%[�!����d���$�e�)��.���3��98���<���@��-E�zI�{�M�fxR�JW��_\�;�a��Sg�Gm�s�6y���~��k���G��(��ͳ��]>��έ�����WF��|��z����  �  ��=�u=),=��=Q�=�7=��=Ԃ=f%=v� =j = =bh�<���<��<vm�<���<�6�</��<�<u~�<���<�T�<���<�<di�<���<B��<V9�<u�<��<���<�-�<@u�<o��<�<�|�<���<T�<��<�>�<ڴ�<�'�<W��<���<�V�<.��<���<�1�<�j�<z��<���<���<�+�<Z�<ň�<̷�<���<�<�>�<Je�<��<��<��<{��<)��<�\�<��<���<�\�<���<�Q�<��<�<�_�<t��<���<�4�<vv�<p��<#��<n.�<�c�<���<w��<�Ӹ<T�<W�<ݲ<�Ȱ<1��<]��<hY�<�+�<,��<�ϣ<��<�}�<�Z�<�<�<�"�<g�<0��<��<�ِ<�Ǝ<���<���<pj�<�;�<��<�Ɓ<�<�zz<Z�u<�fq<��l<zxh<�d<A�_<'�[<�_W<�@S<i,O<mK<lG<��B<��><6�:<�x6<502<H�-<�y)<o%<�� <�@<$�<%�</5<��
<־<��<��;���;f��;��;�#�;OC�;�]�;!n�;�q�;�i�;�Y�;FK�;EI�;�_�;1��;��;y};|fo;�a;�U;�H;$f=;�o2;� (;�;�c;�;&�;���:GH�:���:gս:o%�:��:�L�:��|:�`:��D:�L+: :��9���9���9�j{9R�/9ľ�8g��7G<� ���ҵL�D��!仹��/��w�"�#::�\Q�VMg���|�`s������������
ī������a��=.ú.1˺��Ӻ�iܺ������ ��tx�����:�����7�u�#��(���-��s2��7���;��@�%�D��H��M��JR��?W�>w\���a��g�0�m�D�s���y�������y养J���^��/捻�L������Ŕ��疻g���  �  &�=�n=z'=�=��=
9=�=��=�-=� =�w =� =R��<���<Z6�<"��< ��<�U�<&��<�$�<2��<8��<�Z�<[��<��<c�<H��<���<�&�<�]�<H��<���<�	�<�N�<���<g��<�T�<���<>2�<���<l%�<0��<��<<��<���<�R�<���<���<*:�<x�<��<���<�<gL�<�}�<��<"��<`
�<�4�<�[�<&}�<���<}��<9��<��<���<#X�<��<)��<�K�<��<�7�<H��<��<9�<:��<o��<L
�<�M�<]��<���<��<�J�<�}�<��<�Ǹ<#۶<�<ݲ<�̰<;��<���<�l�<SD�<��<U�<:ɡ<D��<��<�_�<"C�<_)�<G�<���<��<�Ύ<���<*��<�e�<J3�<)��<ѵ�<��~<�Fz<	�u<!q<��l<�'h<t�c<�w_<q>[<�W<1S<}�N<u�J<��F<&�B<��>< �:<�t6<�42<��-<�)<K4%<V� <�w<K<��<�<e@<�
<M�<b��;R]�;2L�;8K�;�T�;a�;�j�;�j�;�^�;QF�;&�;x�;��;���;�!�;��;�L|;[,n;ų`;W�S;��G;�_<;R�1;�>';�e;5�;k�
;5�;��:LO�:�.�:pd�:�:� �:$Ύ:��:P+d:oI:A0:*�:�� :���9R�9΃9�99w��8��8�k3�qh���N�'��Y˾����S!��
&�'�=��FU���k��ƀ� ���Ǒ�����@㥺�̭�%e��{ݼ��_ĺ�̺";Ժ-�ܺS����T���r'��������n�����'��`"��|'�z,��Y1��6���:��f?���C�O�H��SM��2R�>HW���\�/:b�h�b)n��at�q�z��t��􅃻}��{R����񆎻o吻�!��SB��jR��&]���  �  ˪=Vh=�"=��=�=19=?�=��=\4=^� =�� =�* =[��<���<�U�<ذ�<r�<�n�<q��<�5�<7��<���<E^�<ʹ�<��<�[�<���<��<5�<�H�<({�<��<G��<k,�<zx�<���<2�<Ğ�<2�<���<Y�<���<2�<3}�<��<KM�<Ѧ�<K��<�?�<��<���<���<�1�<bg�<e��<F��<f��<6(�<P�<Ms�<���<L��<y��<̲�<���<	��<FR�<�
�<r��<s;�<
��<��<�{�<���<�<
]�<2��<-��<�)�<�n�<K��<���<G3�<oj�<g��<T��<FҶ<�ܴ<�ڲ<�ΰ<b��<?��<e|�<�X�<3�< �<��<�<>��<f}�<�]�<]@�<�$�<�
�<>�<Ԏ<ҳ�<���<?`�<7*�<��<���<4�~<�z<�yu<c�p<LYl<��g<�|c<0_<�Z<��V<�R<��N<1�J<��F<��B<�><5�:<jm6<�42<��-<�)<�N%<=� <��<FS<�<��<u�<J<t<<��;���;H��;���;Bx�;Kt�;n�;*`�;�F�;!�;~�;#Ť;5��;���;��;��;�D{;�m;��_;B�R;�F;�v;;H�0;�&;��;Vs;�X
;�r;�i�:#6�:AQ�:�ƾ:���:�:��:���:S�g:�/M:r�3:=�:��:/��9��92ƈ9�-A9^�8�^8�/�h��\Q�<��U���6���y���(��'A�~�X�,�o�v�q9���ʖ������⧺Z��������9���~ź:ͺ��Ժ�Nݺ>>�m���������-�-z�P�����F�_l!��&���+�+o0��J5��:���>���C�nTH��-M��,R�X_W�=�\�ʅb��|h�˫n��u��h{��※� �����߉�G���	���k������᱕����������  �  ۣ=�b=,=��=*�=�8=c�=��=�8=�� =֊ =�4 =F��<(�<�m�<���<�#�<���<���<�A�<���<��<�_�<l��<�
�<U�<p��<F��<��<u7�<!g�<X��<:��<��<�\�<���<��<��<f��<{z�<��<]}�<:��<�r�<	��<�G�<)��<���<C�<ƈ�<���<��<�B�<�{�<б�<���<��<�>�<�d�<ބ�<���<���<C��< ��<���<!��<�L�<9�<���<�-�<ɥ�<��<�e�<N��<I��<�@�<��<+��<��<bT�<��<�<� �<�Z�<G��<ϰ�<8ʶ<C״<dز<"ϰ<��<���<c��<0g�<,E�<"�<W��<oڟ<���<���<�q�<PQ�<d2�<��<���<׎<ʳ�<ۊ�<�Z�<�!�<�<Z��<�~<��y<,Nu<��p<b$l<	�g<IDc<"�^<8�Z<��V<ٚR<śN<-�J<�F<d�B<��><�:<�e6<�22<�-<��)<a%<!<��<�z<�3<��<b�<�y<H<H<�;���;&��;x��;���;�~�;�l�;�S�;�/�;���;CȬ;�;x`�;�I�;�\�;٧�;�tz;�@l;�^;�R; F;�:;�0;o�%;�Z;J;�

;7;��:��:[�:?�:D�:��:u�:5��:�%j:�P:��6:��:�z:��9���9�^�9q�F9���8�8�-�nj��ʒS�T&���7Ĺ���;d��+�i�C�N�[�p4s�ۤ��|�������V��w��1��QC���O��&kƺ)�ͺ��պ!�ݺ��P�ﺦ�����������MO��z�V���� ���%��*��/���4���9��k>�cDC��$H�|M��/R�_yW���\�	�b���h�ho�U�u�� |�<:���a���k��'M��K ��r����Ց�����V
��	�����  �  F�=�^=A=��=ʇ=M8=��=V�=�;=�� =͏ =�: =���<�#�<q|�<%��<1�<��<q��<�H�<���<1�<B`�<���<��<xP�<<��<b��<4��<-,�<>Z�<݊�<N��<� �<K�<��<O�<st�<:��<�l�<���<s�<���<�k�<���<'D�<��<��<�D�<���<��<"�<wM�<��<���<A��<r"�<�L�<q�<���<,��<��<2��<���< ��<��<�H�<���<V��<�$�<��<3 �<}W�<���<B��<�.�<�q�<���<���<�C�<���<:ҿ<��<%P�<���<ǩ�<�Ķ<fӴ<6ֲ<�ΰ< ��<ꨬ<
��<'p�</P�<�.�<X�<�<*ŝ<S��<�}�<�[�<�:�<p�<@��<W؎<0��<���<�V�<�<�ك<���<�~~<>�y<<2u<x�p<�l<��g<F c<z�^<�Z<��V<�}R<�N<��J<(�F<��B<o�><��:<�_6<S02<��-<@�)<�k%<�"!<�<D�<LO<<��<:�<~c<tl�;"�;���;��;ڜ�;��;�i�;�I�;��;��;��;!k�;�5�;��;�$�;>j�;��y;��k;�9^;�Q;�E;8H:;[�/;��%;1;K�;��	;;���:���:�W�:\�:C]�:��:�t�:�_�:��k:E�Q:ſ8:� :�9	:--�9�?�9���9��I9��8��8dh.��k��zaU��n����Ź<��S���,��sE���]��>u�E������)���2h��x������N������ǺNDκ��պ�޺��溑��N���z�������C�� �5��C �GL%��Q*�,Q/��K4��>9��+>��C�)	H��M��6R��W�{ ]�X�b��i�#`o�'�u��c|�r��럄�V���8���|G���ȏ����]>���B��,3������  �  ��=�]=-=��=@�=&8=��=ّ=x<=�� =�� =�< =`��<r(�<���<��<�5�<���<���<K�<���<�<`�<���<L�<�N�<��<���<��<G(�<�U�<΅�<���<���<�D�<Л�<L��<�n�<���<*h�<���<�o�<���<Oi�<���<�B�<��<���<UE�<ڍ�<���<��<Q�<b��<G��<B��<x'�<CQ�<iu�<"��<��<ظ�<S��<5��<��<�~�<G�<���<���<�!�<���<���<�R�<)��<R��<m(�<:k�<^��<���<�=�<]��<rͿ<`�<�L�<}�<0��<�¶<�Ѵ<uղ<�ΰ<���<��<��<7s�<�S�<L3�<%�<!�<ʝ<���<��<(_�<J=�<6�<j��<�؎<��<���<HU�<y�<E׃<���<�w~<��y<�(u<��p<�k<zyg<c<2�^<B�Z<�{V<�sR<'yN<�J<ɐF<�B<�><�~:<�]6<�/2<N�-<G�)</o%<�'!<�<��<�X<0<�<M�<�l<�|�;�/�;���;p��;h��;���;�h�;�E�;��;)�;���;#_�;�&�;��;P�;�T�;.�y;:�k;|
^;�PQ;d[E;:;͉/;|�%;��;ŷ;��	;U ;S��:���:X�:�)�:
q�:�>�:,��:(��:dDl:sZR:�a9:�;!:.�	:�E�9�+�9�O�9Q�J9��8C�8'W.��+���V�+痹�ƹ=���P�0-��F��t^�
�u�1��6v������Ƣ��Ѫ�kH���\���F���:Ǻtqκ�ֺ)޺��溴�ﺛ������Z��R�����N�4� ��#%��)*�,/��*4��"9�t>�P	C�} H�KM�I8R�ՕW��,]�c�+$i�Pxo�=�u�م|�p��������Ň�a����_��ᏻ@0��HT���V���D��f+���  �  F�=�^=A=��=ʇ=M8=��=V�=�;=�� =͏ =�: =���<�#�<q|�<%��<1�<��<q��<�H�<���<1�<B`�<���<��<xP�<<��<b��<4��<-,�<>Z�<݊�<N��<� �<K�<��<O�<st�<:��<�l�<���<s�<���<�k�<���<'D�<��<��<�D�<���<��<"�<wM�<��<���<A��<r"�<�L�<q�<���<,��<��<2��<���< ��<��<�H�<���<V��<�$�<��<3 �<}W�<���<C��<�.�<�q�<���<���<�C�<���<:ҿ<��<&P�<���<ǩ�<�Ķ<gӴ<7ֲ<�ΰ<��<ꨬ<��<(p�</P�<�.�<X�<�<*ŝ<S��<�}�<�[�<�:�<p�<@��<V؎<0��<���<�V�<�<�ك<��<�~~<=�y<<2u<x�p<�l<��g<F c<z�^<�Z<��V<�}R<�N<��J<)�F<��B<p�><��:<�_6<T02<��-<A�)<�k%<�"!<�<E�<MO<<��<:�<~c<sl�;"�;���;��;ٜ�;��;�i�;�I�;��;��;��;k�;�5�;��;�$�;=j�;��y;��k;�9^;�Q;�E;6H:;Z�/;��%;1;J�;��	;;���:���:�W�:\�:C]�:��:�t�:�_�:��k:E�Q:ſ8:� :�9	:--�9�?�9���9��I9��8��8dh.��k��zaU��n����Ź<��S���,��sE���]��>u�E������)���2h��x������N������ǺNDκ��պ�޺��溑��N���z�������C�� �5��C �GL%��Q*�,Q/��K4��>9��+>��C�)	H��M��6R��W�{ ]�X�b��i�#`o�'�u��c|�r��럄�V���8���|G���ȏ����]>���B��,3������  �  ۣ=�b=,=��=*�=�8=c�=��=�8=�� =֊ =�4 =F��<(�<�m�<���<�#�<���<���<�A�<���<��<�_�<l��<�
�<U�<p��<F��<��<u7�<!g�<X��<:��<��<�\�<���<��<��<f��<{z�<��<]}�<:��<�r�<	��<�G�<)��<���<C�<ƈ�<���<��<�B�<�{�<б�<���<��<�>�<�d�<ބ�<���<���<C��< ��<���<!��<�L�<:�<���<�-�<ɥ�<��<�e�<O��<J��<�@�<��<+��<��<cT�< ��<�<� �<�Z�<H��<а�<9ʶ<D״<eز<#ϰ<��<���<c��<1g�<,E�<"�<W��<oڟ<���<���<�q�<PQ�<c2�<��<���<׎<ɳ�<ڊ�<�Z�<�!�<�<Y��<
�~<��y<+Nu<��p<a$l<	�g<IDc<"�^<9�Z<��V<ښR<ƛN</�J<�F<f�B<��><	�:<�e6<�22<�-<��)<a%<!<��< {<�3<��<b�<�y< H<F<�;���;#��;u��;���;�~�;�l�;�S�;�/�;���;?Ȭ;펤;t`�;�I�;�\�;֧�;�tz;�@l;�^;�R;�F;�:;�0;m�%;�Z;I;�

;7;��:��:[�:>�:D�:��:u�:4��:�%j:�P:��6:��:�z:��9���9�^�9q�F9���8�8�-�nj��ʒS�T&���7Ĺ���;d��+�i�C�N�[�p4s�ۤ��|�������V��w��1��QC���O��&kƺ)�ͺ��պ!�ݺ��P�ﺦ�����������MO��z�V���� ���%��*��/���4���9��k>�cDC��$H�|M��/R�_yW���\�	�b���h�ho�U�u�� |�<:���a���k��'M��K ��r����Ց�����V
��	�����  �  ˪=Vh=�"=��=�=19=?�=��=\4=^� =�� =�* =[��<���<�U�<ذ�<r�<�n�<q��<�5�<7��<���<E^�<ʹ�<��<�[�<���<��<5�<�H�<({�<��<G��<k,�<zx�<���<2�<Ğ�<2�<���<Y�<���<2�<3}�<��<KM�<Ѧ�<K��<�?�<��<���<���<�1�<bg�<e��<F��<f��<6(�<P�<Ms�<���<L��<y��<̲�<���<	��<FR�<�
�<r��<s;�<��<��<�{�<���<�<]�<3��<.��<�)�<�n�<L��<���<H3�<pj�<h��<V��<HҶ<�ܴ<�ڲ<�ΰ<d��<@��<f|�<�X�<3�<!�<��<�<>��<f}�<�]�<\@�<�$�<�
�<=�<Ԏ<ѳ�<���<>`�<6*�<��<���<2�~<�z<�yu<b�p<KYl<��g<�|c<0_<�Z<��V<�R<��N<3�J<��F<��B<�><8�:<lm6<�42<��-<�)<�N%<?� <��<GS<�<��<u�<J<s<:��;���;D��;���;=x�;Ft�;n�;$`�;�F�;� �;x�;Ť;0��;���;���;��;�D{;�m;��_;=�R;�F;�v;;E�0;�&;��;Ts;�X
;�r;�i�:"6�:@Q�:�ƾ:���:�:��:���:R�g:�/M:r�3:=�:��:/��9��92ƈ9�-A9^�8�^8�/�h��\Q�<��U���6���y���(��'A�~�X�,�o�v�q9���ʖ������⧺Z��������9���~ź:ͺ��Ժ�Nݺ>>�m���������-�-z�P�����F�_l!��&���+�+o0��J5��:���>���C�nTH��-M��,R�X_W�=�\�ʅb��|h�˫n��u��h{��※� �����߉�G���	���k������᱕����������  �  &�=�n=z'=�=��=
9=�=��=�-=� =�w =� =R��<���<Z6�<"��< ��<�U�<&��<�$�<2��<8��<�Z�<[��<��<c�<H��<���<�&�<�]�<H��<���<�	�<�N�<���<g��<�T�<���<>2�<���<l%�<0��<��<<��<���<�R�<���<���<*:�<x�<��<���<�<gL�<�}�<��<"��<`
�<�4�<�[�<&}�<���<}��<:��<��<���<#X�<��<)��<�K�<��<�7�<H��<��<9�<;��<p��<M
�<�M�<^��<���<��<�J�<�}�<��<�Ǹ<%۶<�<ݲ<�̰<<��<���<�l�<TD�<��<V�<;ɡ<E��<��<�_�<!C�<^)�<F�<���<��<�Ύ<���<)��<�e�<H3�<'��<ϵ�<��~<�Fz<�u<!q<��l<�'h<t�c<�w_<r>[<�W<3S<�N<w�J<��F<)�B<��><#�:<�t6<�42<��-<�)<M4%<Y� <�w<L<��<�<e@<�
<L�<_��;N]�;.L�;3K�;�T�;a�;�j�;�j�;{^�;IF�;&�;q�;��;���;�!�;��;�L|;S,n;��`;P�S;z�G;�_<;N�1;�>';�e;3�;j�
;3�;��:JO�:�.�:od�:�:� �:$Ύ:��:O+d:oI:A0:*�:�� :���9R�9΃9�99w��8��8�k3�qh���N�'��Y˾����S!��
&�'�=��FU���k��ƀ� ���Ǒ�����@㥺�̭�%e��{ݼ��_ĺ�̺";Ժ-�ܺS����T���r'��������n�����'��`"��|'�z,��Y1��6���:��f?���C�O�H��SM��2R�>HW���\�/:b�h�b)n��at�q�z��t��􅃻}��{R����񆎻o吻�!��SB��jR��&]���  �  ��=�u=),=��=Q�=�7=��=Ԃ=f%=v� =j = =bh�<���<��<vm�<���<�6�</��<�<u~�<���<�T�<���<�<di�<���<B��<V9�<u�<��<���<�-�<@u�<o��<�<�|�<���<T�<��<�>�<ڴ�<�'�<W��<���<�V�<.��<���<�1�<�j�<z��<���<���<�+�<Z�<ň�<̷�<���<�<�>�<Je�<��<��<��<{��<)��<�\�<��<���<�\�<���<�Q�<��<�<�_�<u��<���<�4�<wv�<q��<$��<p.�<�c�<���<y��<�Ӹ<V�<Y�<!ݲ<�Ȱ<2��<^��<jY�<�+�<-��<�ϣ<��<�}�<�Z�<�<�<�"�<f�</��<��<�ِ<�Ǝ<���<���<nj�<�;�<��<�Ɓ<�<�zz<X�u<�fq<��l<zxh<�d<B�_<(�[<�_W<�@S<k,O<oK<oG<��B<��><9�:<�x6<902<L�-<�y)<r%<�� <�@<%�<&�<05<��
<վ<��<��;���;a��;��;~#�;HC�;�]�;n�;�q�;�i�;�Y�;?K�;>I�;�_�;+��;��;y};rfo;�a;�U;�H;f=;�o2;� (;�;�c;�;$�;���:EH�:���:fս:o%�:��:�L�:��|:�`:��D:�L+: :��9���9���9�j{9R�/9þ�8g��7G<� ���ҵL�D��!仹��/��w�"�#::�\Q�VMg���|�`s������������
ī������a��=.ú.1˺��Ӻ�iܺ������ ��tx�����:�����7�u�#��(���-��s2��7���;��@�%�D��H��M��JR��?W�>w\���a��g�0�m�D�s���y�������y养J���^��/捻�L������Ŕ��疻g���  �  H�=�{=�/=�=�=$5=��=m{=h=ĺ =�Z =��<�A�<ܐ�<��<�D�<���<��<Ȅ�<���<�k�<���<AL�<n��<@�<�m�<��<?�<K�<���<���<��<�R�<���<���<�F�<���<��<w�<b��<�W�<���<�6�<ğ�<� �<�X�<��<��<c&�<=Z�<ƈ�<ϳ�<���<g�<�2�<�_�<���<��<���<��<J�<o�<���<���<%��<Q��<_�<X#�<-��<�l�<|��<�k�<V��<\3�<��<~��<N�<�`�<��<���<��<�L�<F}�<���<�Ǻ<n޸<��<u�<�ڲ<���<D��</s�<�B�<|�<"ܥ<���<�|�<BT�<�1�<a�<��<��<���<Ւ<�ɐ<ջ�<���<ʎ�<�l�<<B�<��<�ց<�0<V�z<1-v<�q<H8m<��h<%nd<s`<�[<ҩW<i�S<�cO<�JK<f1G<C<E�><:�:<*x6<�&2<@�-<F\)<S�$<ru <�<Ŗ<05<x�<j�
<Bk<0J<%u�;�s�;	��;��;��;��;'F�;h�;2|�;���;���;H��; ��;Vʕ;�;ʜ�;��~;�p;|:c;E`V;�J;�t>;EY3;��(;;��;�Y;;0�:��:r�:��:��:F��:˓�:_�x:�q[:z�?:Z&:�:���9�X�9��9�m9�$9F��8���7~�J�5����K��ގ�[k���i�z/	�K��Ƃ6���L���b��xw�_˅�Uc������fF��L����ٱ�t깺V	º)Yʺ�Ӻ�ܺ��庨��<���4��Д�%[�!����d���$�e�)��.���3��98���<���@��-E�zI�{�M�fxR�JW��_\�;�a��Sg�Gm�s�6y���~��k���G��(��ͳ��]>��έ�����WF��|��z����  �  ��=X�=[2=��=�=O1=��=�r=f=+� =�J =���<��<�f�<z��<B�<w��<8��<�e�<���<�V�<��<A�<���<��<6o�<���<��<�Z�<٠�<C��<�,�<�v�<���<��<2p�<(��<
1�<|��<��<!o�<���<�C�<���<g�<X�<��<
��<��<�G�<q�<��< ��<���<

�<�5�<od�<R��<���<���<-�<ZW�<&x�<'��<Y��<��<<_�<�'�<���<Dz�<W�<:��<��<�U�<Į�<V��<�H�<��<p��<
�<B9�<�i�<���<���<�Ժ<��<=�<��<�ղ<2��<��<�_�<%*�<��<���<!��<�S�<�)�<��<��<�٘<�̖<oĔ<Y��<׷�<|��<럌<,��<^l�<EF�<m�<(�<�V<0�z<�hv<�q<B�m< i<r�d<Vq`<�+\<�W<��S<ܗO<�sK<PG<�(C<��><��:<r6<2<P�-<�:)<"�$<�> <��<�L<��<{�<F
<S<��<���;���;@�;�Y�;��; ��;�$�;�V�;�{�;)��;ԫ�;�ĥ;��;�-�;��;n&�;N�;��q;�|d;#�W;�?K;�v?;S54;�s);D#;�3;j�;-;���:/��:d��:�0�:��:�
�:Ŀ�:�Nt:űV:��::�� :љ:�a�9>˺9.��9��^9�9�h�8B�l7$^��u �0�L���������Y�0��
��3��H�3�]��yr�?4���ό�|��\�������+�����������ɺ˚Һ��ۺ���9X��N���[�17	��&�x����w� ��&��J+�J=0�J�4�!a9�5�=�"�A���E��J�^GN�z�R�gjW�(_\�4�a��g���l�Grr�KAx��~�7⁻@����h��a��)������|x��}͓�����^���  �  K�=��=�3=��=H�=�,=��=	j=.=�� =; =A��<}��<�>�<�<J��<�\�<���<WG�<���<`A�<��<P4�<��<��<Zn�<$��<}�<^g�<���<-��<�H�<��<(��<=�<ٕ�<���<�R�<I��<$�<4��<���<�M�<۬�<^�<U�<"��<"��<�	�<j4�<2Y�<�z�<R��<���<��<�<<�<;o�<L��<��<��<e?�<�d�<_}�<���<o{�<�\�<$)�<���<ք�<
�<2��<5�<�t�<���<:%�<p�<T��<���<~&�<dW�<��<���<�Ǽ<^޺<��<J�<��<�β<��<���<�K�<��<�ԧ<���<_�<8,�<4�<ߜ<9ƚ<ص�<���<���<঒<�<̟�<M��<���<�i�<�G�<+�<��<kv<u
{<>�v<�1r<��m<Wii<�e<p�`<r\<1X<��S<�O<x�K<�hG<S7C<��><Y�:<�g6<�2<s�-<)<�$<E <�<�<��<*9<x�	<�<�<�P�;�q�;Z��;���;�U�;ì�;���;D=�;�r�;b��;�ĭ;��;E.�;P��;j��;S��;�x�;�s;̠e;'�X;�EL;�\@;f�4;]*;��;�{;Ӵ;�.;j��:[F�:E�:�8�:���:���:��:�+p:TR:��5:��:�:N��9���9���9OIP9�A9s{�8=1�6=�t�x%�cdN�����i���๟:�n����/�.E�G�Y���m��ڀ��x���֓������饺 ����m���2���#ɺY_Һhܺ?,���� ��J����	����(�L���!�.Q'���,�y�1�&"6��~:���>�0�B�0�F���J�N�N��	S�#�W��p\��a���f�Xl��q���w��:}�g��>%���Ն��v��\������o���Yb������j���  �  k�=��=�3=3�=��=�'=*�=�a=�� =w� =- =��<���<>�<�o�<4��<x;�<*��<,�<��<�-�<��<�'�<�<��<�k�<��<��<�p�<l��<��<�_�<~��<��<N\�<k��<��<�n�<���<�0�<&��<���<�T�<���<;�<�P�<^��<��<F��<Q"�<GC�<a�<E~�<~��<���<���<��<�L�<&��<��<���<m)�<�R�<o�<�z�<t�<�X�<�(�<��<Z��<�"�<��<�"�<���<��<�D�<��<5��<*�<�B�<Hp�<|��<y��<�Ҽ<7�<��<=�<P�<ǲ<塰<�q�<f9�<���<+��<>z�<l>�<~	�<�ݞ<���<��<��<���<J��<U��<#��<���<l��<|�<ze�<�F�<�!�<e��<��<F,{<i�v<,er<�n<��i<	Oe<c�`<q�\<�eX<�$T<`�O<q�K<�zG<�@C< ?<��:<5[6<9�1<Cz-<a�(<�g$<��<OI<V�<�P<��<�	<�z<,f<���;&��;]J�;\��;3�;)u�;3��;m �;�b�;F��;�ӭ;(�;a�;�ɖ;�T�;@�;�;b�s;n�f;�Y;^M;�A;�5;C�*;��;��;��;9 ;N[�:%��:�c�:�I�:8�:��:)T�:/l:wN:��1:�8:��9���9o�9ND�9�+C9�9q��8�jڴ� ��==�X�P�b���ӵ��o޹���ʭ�m-���A�@V��.j�l�}�p�������]J��5t��n���ۇ�������ȺvHҺ])ܺ��j�#����\��y
�ج�������"��h(�î-��2��17��z;�M�?��lC�CG�4#K��%O�]S�M�W���\�ފa���f��l�ޏq�w�e�|�P��ٲ��rZ�������������7���b
���z��;闻�  �  �=Ć=!3=\�=Ɂ=#=��=�Z=�� =�� =�! =by�<0��<���<�S�<���<L!�<���<T�<K��<��<���<�<]��<�<�h�<���<R!�<�v�<1��<�<�p�<j��<��<�s�<(��<�'�<��<G��<�?�<���<���<�X�<ư�<h�<
L�<'��<g��<��<r�<�1�<�L�<7g�<5��<��<���<���<�1�<�k�<���<g��<��<D�<c�<�q�<m�<~T�<'�<���<
��<M+�<ѵ�<)2�<���<��<�\�<��<���<�&�<VX�<���<f��<�þ<fڼ<p�<��<i�<�۴<ٿ�<:��<�e�<B*�<��<:��<�b�<�$�<J�<���<柜<F��<�|�<#y�<"{�<��<t��<���<ꀌ<u�<-a�<E�<#�<0��<��<}D{<��v<b�r<0n<|�i<=e<�*a<��\<��X<=FT<�P<|�K<N�G<FC<&�><�:<,O6<��1<�c-<x�(<NF$<��<D<>�<�<{�<�o	<WB< 0<�m�;���;	��;e�;Z��;F�;���;W�;MR�;w��;hۭ;;'�;���;���;ה�;�T�;F@�;�t;HMg;MOZ;��M;��A;6;��*;S  ;��;0�;�;�
�:�F�:��:K��:���:�:��:�i::�J:11.:¹:�
�9,�9��9��|9h�89�)�83Nc8�.ֶ/돸O�BS��쎹����jzݹ���O�0�+�ػ?���S�Vg��z�d
������&��`��P���B嵺�-���Ⱥ;GҺVܺ������S~�������
��@���]��؞#��C)���.��y3��8�HB<��;@�hD�z�G�ƕK���O� �S�bX���\���a�;�f��k�$Kq��v��|�Z����\������ꘈ�h.��Ͻ���F���ɒ��H��Gŗ��  �  ��= �=�2=��=�= =��=�U=� =e� =� =�i�<[��<���<(B�<B��<��<���<w�<��<��<���<��<ʍ�<��<f�<!��<�"�<Xz�< ��<-%�<�z�<���<�)�<D��<���<�5�<א�<j��<�H�<_��<]�<[�<հ�<� �<�H�<J��<��<���<�	�<G&�<�?�<�X�<#t�<ה�<M��< ��<� �<�[�<���<A��<k�<D:�<�Z�<+k�<gh�<\Q�<�%�<���<���<10�<��<�;�<6��<]�<�k�<M��<?��<O5�<�e�<��<}��<�ʾ<�޼<��<��<��<uش<���<���<P]�<9 �<:ݩ<ԗ�<�S�<a�<�ܠ<ޯ�<<��<Gx�<m�<�j�<'n�<�t�<�z�<�}�<�z�<Mp�<�]�<�C�<i#�<���<��<:S{<*�v<��r<�Jn<T�i<�e<�Ga<[�\<¥X<�ZT<yP<��K<�G<HC<q�><��:<�F6<`�1<�T-<
�(<?0$<�<��<^s<��<��<:K	<f<�<�-�;�j�;i��;�7�;J��;�&�;���;���;�E�;��;�ݭ;.3�;���;;�;ѻ�;���;�t�;�$u;��g;%�Z;�$N;��A;�K6;�+;�A ;��;��;7�;[��:���:�X�:s��:��:�G�:�3�:/�g:��H:8
,:��:b��9��9��9�Su9X29"g�83O8�-�s�������U��h��î��~�ܹ�k�}|� �*��^>��R�ݖe�_�x��!��+���Y@��f���y!��*�����e�Ⱥ�OҺ�zܺx�GB����^�3K����o��Y(��"$���)��/� 4�<�8��<��@��qD��#H�@�K�
�O���S��,X���\�C�a�b�f���k�r"q��sv���{�����'���ą�^����������������)�������  �  ��=Tz=%=J�=�r=B=ߴ=/R=�� =i� =�% =���<���<z�<�i�<O��<'.�<���<��<��<��<�y�<3��<�]�<i��<X+�<ω�<���<G:�<Ύ�<���<G6�<P��<%��<�4�<ۊ�<���<A9�<���<$��<�@�<��<���<;�<��<��<��<�;�<�h�<��<��<1��<B��<W
�<�*�<&O�<hw�<��<���<���<.*�<�O�<�l�<�}�<���<�s�<U�<�$�<���</��<�-�<���<>�<���<��<Jy�<R��<l�<ZU�<Ì�<n��< �<@�<� �<G3�<�=�<�>�<�5�<*#�<��<�<e��<̂�<�N�<5�<��<h��<]��<�<"k�<�^�<hX�<�V�<�V�<�V�<T�<mM�<6A�<J/�<��<k��<-ف<ti<�{<�v<!~r<�.n<��i<��e<Ga<I�\<�X<VuT<M5P<��K<P�G<HyC<�4?<,�:<!�6<�12<��-<S)<��$<a_ <K�<9z<<4�<��
<�m<*`< ��;x��;$I�;���;��;�}�;���;P�;���;��;���;<��;�|�;��;Cܒ;���;�Ȅ;�{;�n;0�a;pU;bI;��=;*�2;Z�';�9;&;n5	;��:8�:���:3w�:)��:K�:}��:�e�:�*h:�JK:�N0:�=:� :W��9A̬9��9�E9��8%]]8̀�_n���M$�}oq�J��_�ȹ�M��a�!�9�5��J��^���q�xЂ�����)Q�����g����<��鼺d�ƺڶкۺ���˫������+�	�$����F����!��9'��~,��|1��06���:���>��C�L!G��<K�tpO�b�S�FRX��
]���a�Mg�B2l�vvq���v��|�+���8V������Q���q/��Lō�qX���璻�u�����  �  i�=z=%=��=Is=�=׵=WS=_� =�� =h' =���<���<��<n�<���<E2�<a��<s�<���<��<�{�<
��<"_�<s��<�+�<���<��<=9�<I��<j��<�3�<7��<���<1�<8��<6��<�5�< ��<���<�>�<���<��<�:�<��<���<�<_=�<�j�<���<ҳ�<z��<���<[�<9/�<�S�<�{�<_��<���<��<{-�<�R�<Ao�<��<���<�t�<�U�<�$�<���<S��<W,�<���<v;�<���<;�<�u�<���<��<�Q�<j��<r��<l�<t�<W�<�2�<c=�<�>�<�6�<d$�<5�<&�<���<�<>R�<��<��<�à<���<o��<io�<�b�<#\�<�Y�<�Y�<Y�<V�<O�<sB�< 0�<��<��<K؁<�f<�{<��v<%xr<(n<��i<9�e<�?a<X�\<˱X<�oT<�0P<��K<@�G<HxC<�4?<5�:<G�6<�42<��-<�W)<c�$<�e <��<?�<�"<4�<~�
<�v<�h<6��;D�;V�;��;`�;���;2��;�T�;(��;L�;��;��;Zw�;	�;�ђ;Ȳ�;���;U�{;�n;�a;�VU;LI;B�=;-x2;G�';J4;�;P7	;-�:xM�:���:]��:�ε:�z�:Ϸ�:ա�:��h:��K:��0:��:n� :��9���9���93�F9��8��a8k4t�!��i�#��Rq��U��=�ȹ��{S���!�O76�pJ��}^��^r�
���ό������'������FV��������ƺl�к�ںɖ���,���/����	�����������!��'�`\,��Y1��6���:�a�>���B��
G��)K��`O�+�S��HX��]���a�Dg��9l�2�q�f�v��)|�����c��
��룈��=���ҍ��d��{�[~���
���  �  ��=�y=&%=Z�=�t=�=��=�V=^� =�� =�, =��<��<�&�<{�<���<S>�<���<��<��<U�<H��<��<�b�<���<-�<���<���<�5�<t��<���<�+�<�}�<V��< &�<2|�<���<,�<���<k��<&9�<���<���<:�<���<���<C�<�A�<�p�<��<1��<��<���<�<�;�<j`�<���<ݳ�<���<V�<7�<[�<Dv�<���<��<�w�<�W�<b%�<���<ƌ�<(�<Ǵ�<�3�<æ�<��<j�<���<"�<�F�<_�<Ȱ�<)ۿ<���<Y�<E0�<�<�<�?�<�8�<�'�<��<��<+��<H��<\�<�)�<���<qР<���<e��<�{�<Gn�<�f�<Kc�<�a�<�_�<�[�<SS�<�E�<�1�< �<7��<�Ձ<M^<�{<ιv<Rfr<�n<�i<�te<�)a<��\<U�X<`T<
$P<��K<�G<uC<�4?<��:<��6<p<2<�-<�d)<o�$<=x <�<}�<�;<��<&�
<�<��<��;�6�;�{�;���;�5�;ƛ�; �;a�;���;��;�{�;O�;�e�;���;���;��;ϓ�;N�{;�Nn;�wa;4
U;
I;Dv=;�M2;Ί';�#;�;>	;HP�:N��:��:��:�A�:�:�S�:�P�:�%j:�hM:�|2:mj:�#:���9!{�9�0�9��J9��9pjm8�gO�\���I�"���p��v���Gɹ~��� ���"�xD7��K�|�_��s�Ҹ��w����.����*�������1����ƺ3�кG�ںLp�i\��������	�n�����Mq�)-!���&�}�+���0�L�5�x*:��w>�\�B���F���J��4O��S�"1X��\���a�g�UOl���q�
w��e|�}ျ����0��Ј��h�������������얕�����  �  z�=9x=%=Q�=�v==��=�[=~� =Ė =�4 =$��<_��<�:�<^��<e��<jQ�<Q��<u.�<Т�<�<���<���<sh�<���<�.�<ӈ�<j��<l0�<B��<4��<��<�n�<���<��<�j�<���<@�<�w�<���<�/�<��<���<18�<3��<n��<��<�H�<wy�<ԣ�<��<��<��<{,�<#O�<�t�<���<\��<.��<7�<F�<�g�<��<O��<v��<c|�<Z�<�%�<w��<=��< !�<���<�'�<"��<s��<�X�<}��<���<5�<(o�<���<SϿ<���<��<,�<�:�<@�<Y;�<I,�<��<��<<ɫ<���<Rk�<-;�<l�<�<���<z��<8��<���<pw�<r�<�n�<�j�<\d�<�Y�<J�<94�<U�< ��<с<�O<@�z</�v<,Ir<�m<<�i<Qe<�a<S�\<5�X<+FT<�P<��K<C�G<�oC<Q3?<4�:<(�6<;H2<�-<y)<%<>� <�%<,�<�b<�<��
<��<�<~U�;y�;j��;��;y_�;���;��;Qr�;�ƿ;��;&r�;Ԩ;�G�;�ԙ;���;6U�; T�;�{;��m;?�`;?�T;�H;�=;I2; Y';C;�;EE	;��:���:��:Y��:-�:�ե:iF�:%a�:{l:��O:�5:��:U�:���9�ô9f��9�oQ9�{9�q8T���ب��^!�ōp��ݠ�y?ʹ�%��#"��#$�,�8�{�M���a�t�u�pЄ�f������D~���٪�z.������oǺ\�к�ںl;庀��0��aY�R7	�%���p��g� �4&�LR+�=Q0�H5���9�A�=��2B��eF���J�3�N��iS�MX���\��a�2!g��tl���q��Rw���|�o���̃��u�����歋��<��]Ð�/C��q����:���  �  ��=%v=x$=(�=�x=�=]�=�a==ɟ =? =��<�<�T�<���<�<�i�<���<�B�<A��<�&�<ӗ�<��<�n�<E��<�/�<��<���<�(�<u�<���<��<�Z�<���<p��<%S�<ɫ�<7�<�d�<���< #�<���<z��<5�<��<���<!�<XP�<��<*��<3��<���<� �<D�<:h�<h��<���<~��<�
�<�3�<�X�<x�<H��<���<��<T��<4\�<%�<���<���<�<���<�<���<���<�@�<��<;��<��<�Y�<���<\��<��<U�<�%�<�7�<�?�<�=�<�1�<|�<���<�֫< ��<�~�<�P�<`%�<w��<�ڞ<d��<4��<���<���<���<a~�<�w�<�n�<�a�<O�<�6�<��<j�<wʁ<�;<|�z<�v<k"r<��m<�qi<w!e<��`<�\<2YX<e#T<p�O<��K<�G<GfC<C0?<��:<5�6<�U2<�-<�)<k&%<�� <|O<��<F�<YL<�<��<��<ܲ�;;��;* �;7D�;���;���;U7�;P��;JϿ;a�;�b�;5��;c�;@��;V?�;X�;���;�Pz;1m;D`;��S;�H;Ţ<;Ħ1;�';��; �;VH	;��:�.�:��:7�:η:>ܦ:
y�:���:6uo:�	S:`K8:";:��:���9"0�9�ђ9��Y9V9ߩ�8�p���J�����sp����{�˹f����~&�]L;�6P�V�d���x��E��f揺�T�������ƫ�贺����cǺ��кY�ںW庸�ﺃ������C�����^q�4�����E%�Ӏ*� �/�$J4�f�8� M=��A���E��:J���N�~/S� �W��\�$�a��?g�4�l�%/r�<�w�NL}�|h���"���ц�t��^
������}������~����d���  �  �=4s=3#=w�=�z=�!=i�=�h=t	=ѩ =�J =��<0#�<r�<[��<A#�<w��<3��<$Y�<���<�6�<���<�<u�<Z��<}/�<փ�<���<�<�f�<��<���<�B�<]��<���<h7�<Ґ�<���<;N�<y��<��<�u�<��<V0�<���<���<��<AX�<)��<���<��<�<9�<�^�<���<��<2��<��<}%�<�K�<5n�<��<���<ģ�<Ü�<ԅ�<s]�<#�<���<�x�<]
�<Q��<��<%m�<G��<�$�<�t�<3��<��<�?�<�x�<꫿<ٽ<5��<��<�2�<P>�<�?�<q6�<�#�<2�<��<m��<l��<�i�<~@�<\�<���<�ۜ<�Ě<c��<w��<��<叒<텐<�y�<-i�<�S�<�7�<��<1�<u��<]"<��z<�Wv<��q<��m<�:i<0�d<.�`<3`\<)X<m�S<��O<ݨK<��G<gYC<3*?<0�:<�6<�b2<�.<��)<H%<$� <�~<�!<��<��<�Q<+<�<��;,�;R�;���;���;�;�T�;`��;~ӿ;��;UL�;���;r�;�[�;��;���;l��;�{y;x:l;Rs_;�*S;`G;�<;�/1;,�&;)�;��;�@	;���:���:��:g��:���:���:�З:VC�:��r:��V:D<:��":�d:-c�9�\�9�:�9/�b9��9�A�8���������q�ȣ���͹AN��_���q(��>��TS�eh�U|�# ��]���qۚ����[謺�ε�v�����Ǻh(Ѻ�ںy�亁F�R��f��SH�s�9���j�,��:]$���)���.��g3�y8��<�U�@��`E��I�ON���R�7�W�c�\��b��kg���l�Εr��Ax���}�FŁ�R����>���㉻�w��?����o��Yؓ��9��♘��  �  Y�=Po=!=�=|=�$=�=*o=�=� =�V =��<�@�<���<���<�A�<s��<��<Xp�<K��<�F�<���<��<7z�<'��<�-�<�~�<Q��<��<�V�<���<0��<�'�<rs�<���<��<*s�</��<,5�<�<��<�g�<���<�)�<h��<���<��<P_�<���<���<��<�(�<R�<vz�<���<���<7��<�<lA�<�d�<݃�<��<��<-��<���<��<Y]�<n�<i��<�m�<���<�z�<b��<S�<T��<��<�T�<X��< ��<d#�</_�<<�ƽ<�<2�<1,�<-;�<�?�<!:�<�*�<�<���<ѩ<���<l��<�\�<�8�<��<���<d�<�͘<��<���<���<Ǔ�<ʃ�<�o�<�V�<�7�<l�<�<���<�<#�z<�*v<��q<�Zm<�h<�d<c`<&\<��W<Z�S<̧O<�K<WjG<�HC<� ?<��:<Q�6<En2<_.<��)<�i%<�!<T�<�X<�
<��<��<Vj<�P<D��;Í�;���;'��;� �;�7�;�n�;���;Aҿ;���;�.�;f�;*��;��;c��; E�;�)�;i�x;RMk;��^;�SR;��F;�g;;��0;�M&;P;�;�,	;���:���:��:���:���:&�:�/�:�؉:*Xv:�kZ:��?:\�&:0:[w�9���9���9�!l9I095J�8d�!6H��o���ar�R1��8#йS�������+��)A��V��k�+�� 扺F`��F����s���0��ٶ�"����eȺnѺ��ں���o�����<�}���i������6��h#�M�(���-�kz2�z27�=�;�0U@���D��`I�� N��R�#�W���\��%b���g�`Mm��s�H�x��~�:,��q���r���2^���>m���ב�4��؆��&ט��  �  ��=�j=3=��=�|=*'=�=u=�=ѽ ==b =� =>]�<��<O�<�_�<���<7!�<���<���<[U�<���<��<�}�<[��<�*�<Ex�<L��<'�<QE�<��<���<d�<�U�<���<���<�T�<���<2�<��<a��<X�<?��<�!�<�}�<���<��<�d�<��<���<��<A=�<(j�<}��<���<(��<��<<8�<�\�<2}�<���<߬�<Ƿ�<4��<��<Ҋ�<�[�<X�<���<sa�<|��<�f�<���<8�<���<��<4�<�}�<���<�<�D�<�<���<��<s�<$�<�6�<�>�<Y<�<�0�<��<�<��<��<2��<~x�<8V�<Q6�<1�<R��<��<�Ԗ< Ô<�<N��<���<<u�<�X�<<6�<m�<�ރ<m��<��~<_pz<��u<��q<> m<��h<�kd<j$`<_�[<ȼW<��S<�}O<lfK<�OG<5C<?<	�:<��6<�v2<�-.<��)< �%<�2!<3�<�<#E<�<�< �<f�<��;���;~��; �;(1�;�Y�;���;���;�ʿ;{�;c�;84�;�l�;���;�6�;0ۉ;���;��w;�Zj;�];�uQ;��E;D�:;�0;��%;�;�c;�	;��:*��:�f�:;�:�{�:\9�:D��:a_�:��y:�^:�C:е*:��:oX�9���9�9��t9��$9y�8�Ʊ6K�������ut����-�ҹ�8 �q�_�-�R]D�RQZ���o�-��(؋��?��HH��A��&���d���Km��(ɺ��Ѻ�&ۺ\�����-$�����sY�4��IY�����2��z"�E�'�ݫ,��1�F^6��;��?��VD���H�w�M�>�R�/�W�y�\��Pb�a�g�u�m���s��wy�"\������n��x1��dۊ�lk���⏻iC��(���"ؖ�����  �  Q�=�e=�=�=J|=�(=(�=�y=\ =S� =�l =� =Hw�<���<!�<�z�<4��<@8�<���<!��<�a�<���<<$�<��<;��<�&�<�p�<���<(��<�3�<?q�<ׯ�<��<G9�<���<���<�7�<=��<%�<n�<���<�H�<��<��<x�<��<> �<�h�</��<���<h�<|O�<��<��</��<��<-�<�R�<u�<��<���<u��<���<h��<x��<&��<�X�< �<W��<�T�<Y��<S�<��<�</v�<���<��<�^�<���<��<K+�<�h�<���<һ<3��<�<�0�<�;�<=�<�4�<d$�<��<��<�ҧ<y��<���<q�<�Q�<�4�<��<� �<�<�Ԕ<%��<���<���<�x�<�X�<X3�<]�<=Ճ<���<��~<tIz<�u<Wq<E�l<Ƅh<M/d<��_<g�[<�W<%jS<�TO<DK<�3G<% C<�?<��:<��6<�{2<�9.<e�)<#�%<bU!<<[�<]z<�=<%
< �<��<�V�;�?�;;�;RE�;�Y�;�s�;���;Ѩ�;|��;eѷ;J�;� �;�+�;4q�;Hې;�u�;	I�;ӻv;�si;�\;+�P;E;�:;��/;Cc%;w�;J";i�;���:��::��:���:B2�:(�:v��:O��:��|:�pa:�<G:�0.:�;:���9l�9���9�V|9��*9��8��6��� ��#w�9��W�չ��h�Z�0��uG��]��1s��⃺;�������񟺠����ذ�V���R��H�ɺ�iҺqۺ��争������������Y�I��	�h���!�S�&���+��0�a�5��i:�U*?�#�C��H�l�M�ӃR�ϧW���\���b��9h��n�Lt��z�)	������݅������R��
፻�R��窒���'��\���  �  )�= a=k= �=�{=$)=P�=�}=�%=K� =u =V =��<���<�8�<��<���<aK�<��<^�<�k�<3��<�'�<���<��<�!�<pi�<���<;��<[$�<�^�<њ�<���<M �<m�<���<)�<��<��<SZ�<���<�:�<���<1�<r�<���<��<�j�<t��<-��<#(�<g^�<���<D��<i��<��<HD�<i�<���<���<���<@��<$��<���<���<5��<�T�<��<?��<�H�<���<lA�<x��<?�<"]�<P��<���<�C�<c��<d��<��<�T�<���<�û<��<V�<�*�<�8�<|<�</7�<�)�<u�<��<��<�ĥ<e��<���<Wi�<�K�<�/�<��<���<Y�<�˒< ��<���<�z�<X�<�/�<�<L̃<瑁<N�~<W&z<��u<�)q<�l<�Ph<=�c<g�_<>[<iYW<9@S<)0O<%K<8G<BC<�><��:<D�6<�}2<-B.<��)<��%<�q!<�*<r�<�<Vm<w:<�<��<���;V��; t�;Jq�;�x�;���;"��;i��;L��;���;���;�Ч;��;�*�;���;��;e�;��u;��h;/�[;�O;liD;�v9;K/;Z�$;�F;�;��;E��:
��:���:�:^��:��:㜜:��:o:�@d:,J:� 1:W:p�:Q�9Ș�9�7�9�/9_d�8f7[Ӗ�8�!�U�y�|K����ع\���|�|3�.J���`��]v�����+R��暘�3j���ة�"�����~&º�bʺ[�Һ��ۺ��������q��������<�$������ ��	&��+�40��4���9��>���C�fpH�[dM�wR���W��]��b�7�h��wn��t�i�z��Y��=W���?��Z��b���'H��������A��+o������  �  %�=]=p=�=�z=X)=��="�=�)=n� =f{ =�$ =k��<���<'J�<��<���<�Y�<��<�<s�<���<%*�<i��<���<o�<c�<"��<���<��<P�<C��<p��<��<�X�<M��<d
�<2o�<���<�J�<��<"/�<X��<��<�l�<���<h�<l�<��<��<�0�<mi�<��<���<�<M-�<�U�<�y�<���<q��<��<���<��<���<���<Ո�<�Q�<%�<���<�>�<���<Z3�<a��<;��<~I�<���<���<p.�<�v�<��<,�<�D�<ׁ�<��<B�<�
�<c%�<v5�<p;�<�8�<�-�<��<�<�<�ҥ<��<���<�z�<Z]�<L@�<$�<��<�<�Ӓ<���<Λ�<�{�<�V�<],�<���<�ă<8��<��~<U
z<��u<�q<[�l<�(h<3�c<�_<X[<�4W<.S<�O<K<jG<��B<��><��:<,�6<	~2<wG.<
*<2�%<`�!<sD<�<`�<��<�^<'3<g<��;��;���;��;��;Ȓ�;Θ�;|��;��;��;�;m��;��;��;K�;5Ո;5��;�Vu;Uh;�`[;=TO;��C;�8;Ҙ.;��$;��;ժ;ޑ;�[�:���:���:M�:5!�:7v�:�P�:��:
��:C]f:w_L:�U3:K.:A�:^r�9�p�9Wt�9C429�(�8�k7/���#�lx|����~�ڹe:��&���4��SL��
c���x��Ȇ����/ә�����7媺d�fߺ�6�º?�ʺBOӺxܺ^*�V������eO�2t���������?�Hc ��|%�ˊ*�@�/���4�gw9��c>�YOC�ZEH�kLM��qR�v�W��8]���b�6�h��n��t��{�����Y���s����\��x��������M�����?����ș��  �  �=cZ=z=��=�y=H)=Q�=��=�+=�� =? =F) =���<���<2U�<˭�<��<�b�<{��<��<Ow�<\��<	+�<��<��<h�<�^�<���<���<��<�F�<��<߼�<� �<�K�<R��<���<Bc�<���<�@�<[��<�'�<F��<�<Pi�<7��<n�<`l�<���<���<�5�<0p�<3��<��<��<,8�<�`�<D��<���<���<���<	��<���<���<Я�<���<�N�<`�<���<�8�<���<J*�<��<���<=�<���<��<� �<�i�<ʱ�<���<�:�<�x�<���<�<�<�!�<3�<~:�<�8�<�/�<� �<��<$��<Pۥ<俣<7��<⅟<7h�<�J�<l-�<��<���<�ؒ<��<o��<�{�<�U�<�)�<���<���<<C�~<a�y<#qu<E�p<�wl<�h<�c<�q_<S?[<�W<�	S< O<��J<��F<��B<K�><��:<�6<�}2<�I.<*<_�%<�!<T<*<P�<�<�u<JI<W#<� <`��;g��;��;���;a��;/��;u��;ٖ�;��;���;��;��;�Η;7"�;���;Wm�;	�t;��g;��Z;��N;r�C;Ա8;�U.;�f$;x�;l�;�w;:�:���:x��:%m�:?\�:Rʬ:d��:Y?�:J�:��g:}�M:2�4:��:):���9�/�9ʄ949�6�87ᇘ�<$$�"-~��9���eܹ�#�^9��+6���M���d��gz�M����d��R���L��^���4����d���Aú>H˺1�Ӻ>ܺ�H�ܴ�)u���;��S��y�������3�� ��$%��3*��;/�=4��89�G0>�|)C��+H��@M��qR��W��M]�c��h��n�*#u��X{����˃�ؼ��n���z@���ˎ��2���{�������̗�7虻�  �  ��=mY=�=!�=�y=M)=��= �=�,=�� =�� =�* =��<[�<�X�<T��<�<|e�<��<��<�x�<A��<`+�<��<d��<2�<D]�<���<���<��<nC�<�{�<۸�<8��<�G�<��<H��<5_�<���<a=�<Q��<%�<��<M�<�g�<@��<�<zl�<Y��<���<y7�<�r�<���<@��<��<�;�</d�<���<���<p��<L��<���<���<^��<��<a��<�M�<��<���<W6�<7��<!'�<w��<���<�8�<���<x��<N�<ee�<���<���<X7�<�u�<���<�ݹ<M�<X �<02�<<:�<9�<�0�<�!�<Z�<���<#ޥ<,ã<���<���<�k�<N�<�0�<��< ��<=ڒ<��<���<�{�<0U�<�(�<���<⽃<��<�z~<8�y< ju<u�p<�ol<�h<2�c<�h_<�6[<�W<�S<��N<�J<*�F<��B<=�><X�:<��6<�}2<�J.<�*<=�%<r�!<�Y<f<L�<d�<}<�P<W*</
 <u��;��;۩�;Ԟ�;m��;���;Y��;���;��;2��;��;3��;z;��;��;�\�;��t;�g;��Z;$�N;�nC;�8;*>.;4R$;��;,y;Tm;�+�:F��:,��:�w�:�n�:n�:��:�l�:c}�::h:E3N:!*5:��:Dt:�?�9�Ͱ9D9�9�496�8�N 7ɘ�-�$�v�~�$���[�ܹ�v�J��p�6�h,N��e���z��݇�ت���ߚ������̫�����S����hú.i˺ĮӺRܺ;U�ö�|p��15��I�Rj�Q�����������b%�=*�. /�h$4��"9�>��C��#H��<M�qR���W�CV]�|c��h�o��8u�Mq{��Ѐ�ۃ�f͆������Q��<ݎ��C��?������5ٗ�;��  �  �=cZ=z=��=�y=H)=Q�=��=�+=�� =? =F) =���<���<2U�<˭�<��<�b�<{��<��<Ow�<\��<	+�<��<��<h�<�^�<���<���<��<�F�<��<߼�<� �<�K�<R��<���<Bc�<���<�@�<[��<�'�<F��<�<Pi�<7��<n�<`l�<���<���<�5�<0p�<3��<��<��<,8�<�`�<D��<���<���<���<	��<���<���<Я�<���<�N�<`�<���<�8�<���<J*�<��<���<=�<���<��<� �<�i�<ʱ�<���<�:�<�x�<���<�<�<�!�<3�<~:�<�8�<�/�<� �<��<$��<Pۥ<忣<7��<⅟<7h�<�J�<l-�<��<���<�ؒ<��<o��<�{�<�U�<�)�<���<���<<B�~<`�y<#qu<E�p<�wl<�h<�c<�q_<S?[<�W<�	S< O<��J<��F<��B<L�><��:<�6<�}2<�I.<*<`�%<�!<T<*<Q�<�<�u<JI<W#<� <_��;f��;��;���;_��;.��;s��;ז�;��;���;��;��;�Η;6"�;���;Vm�;�t;~�g;��Z;��N;p�C;ӱ8;�U.;�f$;w�;l�;�w;:�:���:w��:%m�:?\�:Rʬ:d��:Y?�:J�:��g:}�M:2�4:��:):���9�/�9ʄ949�6�87ᇘ�<$$�"-~��9���eܹ�#�^9��+6���M���d��gz�M����d��R���L��^���4����d���Aú>H˺1�Ӻ>ܺ�H�ܴ�)u���;��S��y�������3�� ��$%��3*��;/�=4��89�G0>�|)C��+H��@M��qR��W��M]�c��h��n�*#u��X{����˃�ؼ��n���z@���ˎ��2���{�������̗�7虻�  �  %�=]=p=�=�z=X)=��="�=�)=n� =f{ =�$ =k��<���<'J�<��<���<�Y�<��<�<s�<���<%*�<i��<���<o�<c�<"��<���<��<P�<C��<p��<��<�X�<M��<d
�<2o�<���<�J�<��<"/�<X��<��<�l�<���<h�<l�<��<��<�0�<mi�<��<���<�<M-�<�U�<�y�<���<q��<��<���<��<���<���<Ո�<�Q�<%�<���<�>�<���<Z3�<a��<;��<I�<���<���<p.�<�v�<��<,�<�D�<؁�<��<B�<�
�<c%�<w5�<q;�<�8�<�-�<��<�<�<�ҥ<��<���<�z�<Z]�<L@�<$�<��<�<�Ӓ<���<Λ�<�{�<�V�<\,�<���<�ă<8��<��~<T
z<��u<�q<Z�l<�(h<3�c<�_<X[<�4W</S<�O<K<kG<��B<��><��:<-�6<~2<xG.<
*<3�%<a�!<tD<�<`�<��<�^<'3<g<��;��;���;��;��;ƒ�;˘�;y��;��;��;�;j��;��;��;	K�;3Ո;3��;�Vu;Rh;�`[;:TO;��C;�8;И.;��$;��;Ԫ;ݑ;�[�:���:���:
M�:4!�:7v�:�P�:��:
��:C]f:w_L:�U3:K.:A�:^r�9�p�9Wt�9C429�(�8�k7/���#�lx|����~�ڹe:��&���4��SL��
c���x��Ȇ����/ә�����7媺d�fߺ�6�º?�ʺBOӺxܺ^*�V������eO�2t���������?�Hc ��|%�ˊ*�@�/���4�gw9��c>�YOC�ZEH�kLM��qR�v�W��8]���b�6�h��n��t��{�����Y���s����\��x��������M�����?����ș��  �  )�= a=k= �=�{=$)=P�=�}=�%=K� =u =V =��<���<�8�<��<���<aK�<��<^�<�k�<3��<�'�<���<��<�!�<pi�<���<;��<[$�<�^�<њ�<���<M �<m�<���<)�<��<��<SZ�<���<�:�<���<1�<r�<���<��<�j�<t��<-��<#(�<g^�<���<D��<i��<��<HD�<i�<���<���<���<@��<$��<���<���<5��<�T�<��<?��<�H�<���<lA�<x��<@�<"]�<Q��<���<�C�<c��<e��<��<�T�<���<�û<��<W�<�*�<�8�<}<�<07�<�)�<u�<��<��<�ĥ<e��<���<Wi�<�K�<�/�<��<���<X�<�˒<���<���<�z�<X�<�/�<�<K̃<摁<M�~<V&z<��u<�)q<�l<�Ph<=�c<g�_<?[<iYW<:@S<+0O<%K<:G<DC<�><��:<E�6<�}2</B.<��)<��%<�q!<�*<s�<�<Vm<w:<�<��<���;T��;�s�;Gq�;�x�;~��;��;d��;H��;���;���;�Ч;��;�*�;���;��;b�;��u;��h;+�[;�O;hiD;�v9;I/;X�$;�F;�;��;D��:	��:���:�:^��:��:✜:��:o:�@d:,J:� 1:W:p�:Q�9Ș�9�7�9�/9_d�8f7[Ӗ�8�!�U�y�|K����ع\���|�|3�.J���`��]v�����+R��暘�3j���ة�"�����~&º�bʺ[�Һ��ۺ��������q��������<�$������ ��	&��+�40��4���9��>���C�fpH�[dM�wR���W��]��b�7�h��wn��t�i�z��Y��=W���?��Z��b���'H��������A��+o������  �  Q�=�e=�=�=J|=�(=(�=�y=\ =S� =�l =� =Hw�<���<!�<�z�<4��<@8�<���<!��<�a�<���<<$�<��<;��<�&�<�p�<���<(��<�3�<?q�<ׯ�<��<G9�<���<���<�7�<=��<%�<n�<���<�H�<��<��<x�<��<> �<�h�</��<���<h�<|O�<��<��</��<��<-�<�R�<u�<��<���<u��<���<h��<x��<&��<�X�< �<W��<�T�<Y��<S�<��<�<0v�<���<��<�^�<���<��<L+�<�h�<���<һ<5��<�<�0�<�;�<=�<�4�<e$�<��<��<�ҧ<z��<���<q�<�Q�<�4�<��<� �<�<�Ԕ<$��<���<���<�x�<�X�<V3�<\�<<Ճ<���<�~<sIz<�u<Wq<E�l<ńh<M/d<��_<g�[<�W<'jS<�TO<DK<�3G<' C<�?<��:<��6<�{2<�9.<g�)<%�%<cU!<<\�<^z<�=<%
<�<��<�V�;�?�; ;�;NE�;�Y�;�s�;���;˨�;v��;`ѷ;E�;� �;�+�;/q�;Dې;�u�;I�;̻v;�si;�\;'�P;E;�:;ރ/;Ac%;u�;I";h�;���:��:9��:���:A2�:(�:u��:N��:��|:�pa:�<G:�0.:�;:���9l�9���9�V|9��*9��8��6��� ��#w�9��W�չ��h�Z�0��uG��]��1s��⃺;�������񟺠����ذ�V���R��H�ɺ�iҺqۺ��争������������Y�I��	�h���!�S�&���+��0�a�5��i:�U*?�#�C��H�l�M�ӃR�ϧW���\���b��9h��n�Lt��z�)	������݅������R��
፻�R��窒���'��\���  �  ��=�j=3=��=�|=*'=�=u=�=ѽ ==b =� =>]�<��<O�<�_�<���<7!�<���<���<[U�<���<��<�}�<[��<�*�<Ex�<L��<'�<QE�<��<���<d�<�U�<���<���<�T�<���<2�<��<a��<X�<?��<�!�<�}�<���<��<�d�<��<���<��<A=�<(j�<}��<���<(��<��<<8�<�\�<2}�<���<߬�<Ƿ�<4��<��<Ҋ�<�[�<X�<���<sa�<|��<�f�<���<8�<���<��<4�<�}�<���<�<�D�<�<���<��<u�<$�<�6�<�>�<[<�<�0�<��<�<��<��<2��<~x�<8V�<Q6�<1�<Q��<��<�Ԗ<�<ﱒ<M��<���<;u�<�X�<;6�<l�<�ރ<l��<��~<]pz<��u<��q<= m<��h<�kd<j$`<`�[<ɼW<��S<�}O<nfK<�OG<5C<?<�:<��6<�v2<�-.<��)<"�%<�2!<4�<�<$E<�<�< �<e�<��;���;z��;��;#1�;�Y�;���;���;�ʿ;u�;]�;24�;�l�;���;�6�;,ۉ;���;�w;�Zj;�];�uQ;��E;A�:;�0;��%;�;�c;~	;��:(��:�f�:;�:�{�:[9�:D��:a_�:��y:�^:�C:е*:��:oX�9���9�9��t9��$9y�8�Ʊ6K�������ut����-�ҹ�8 �q�_�-�R]D�RQZ���o�-��(؋��?��HH��A��&���d���Km��(ɺ��Ѻ�&ۺ\�����-$�����sY�4��IY�����2��z"�E�'�ݫ,��1�F^6��;��?��VD���H�w�M�>�R�/�W�y�\��Pb�a�g�u�m���s��wy�"\������n��x1��dۊ�lk���⏻iC��(���"ؖ�����  �  Y�=Po=!=�=|=�$=�=*o=�=� =�V =��<�@�<���<���<�A�<s��<��<Xp�<K��<�F�<���<��<7z�<'��<�-�<�~�<Q��<��<�V�<���<0��<�'�<rs�<���<��<*s�</��<,5�<�<��<�g�<���<�)�<h��<���<��<P_�<���<���<��<�(�<R�<vz�<���<���<7��<�<lA�<�d�<݃�<��<��<-��<���<��<Y]�<n�<i��<�m�<���<�z�<b��<S�<U��<��<�T�<X��<!��<e#�<0_�<�<�ƽ<�<4�<3,�<.;�<�?�<#:�<�*�<�<���<ѩ<���<m��<�\�<�8�<��<���<c�<�͘<��<���<���<Ɠ�<Ƀ�<�o�<�V�<�7�<k�<�<���<�<!�z<�*v<��q<�Zm<�h<�d<c`< &\<��W<\�S<ͧO<��K<YjG<�HC<� ?<��:<T�6<Hn2<b.<��)<�i%<�!<V�<�X<�
<��<��<Uj<�P<B��;���;��;"��;� �;�7�;�n�;���;;ҿ;���;�.�;f�;$��;��;^��;E�;�)�;a�x;KMk;��^;�SR;��F;�g;;��0;�M&;P;�;�,	;���:���:��:���:���:&�:�/�:�؉:*Xv:�kZ:��?:\�&:0:[w�9���9���9�!l9I095J�8d�!6H��o���ar�R1��8#йS�������+��)A��V��k�+�� 扺F`��F����s���0��ٶ�"����eȺnѺ��ں���o�����<�}���i������6��h#�M�(���-�kz2�z27�=�;�0U@���D��`I�� N��R�#�W���\��%b���g�`Mm��s�H�x��~�:,��q���r���2^���>m���ב�4��؆��&ט��  �  �=4s=3#=w�=�z=�!=i�=�h=t	=ѩ =�J =��<0#�<r�<[��<A#�<w��<3��<$Y�<���<�6�<���<�<u�<Z��<}/�<փ�<���<�<�f�<��<���<�B�<]��<���<h7�<Ґ�<���<;N�<y��<��<�u�<��<V0�<���<���<��<AX�<)��<���<��<�<9�<�^�<���<��<2��<��<}%�<�K�<5n�<��<���<ģ�<Ü�<ԅ�<s]�<	#�<���<�x�<]
�<R��<��<&m�<G��<�$�<�t�<4��<��<�?�<�x�<뫿<ٽ<6��<��<�2�<R>�<�?�<r6�<�#�<3�<��<n��<m��<�i�<@�<\�<���<�ۜ<�Ě<b��<v��<~��<䏒<셐<�y�<+i�<�S�<�7�<��<0�<t��<Z"<��z<�Wv<��q<��m<�:i<0�d</�`<4`\<)X<n�S<��O<ߨK<��G<jYC<6*?<3�:<
�6<�b2<�.<��)<H%<&� <�~<�!<��<��<�Q<+<�<��;,�;R�;���;���;�;�T�;Z��;xӿ;��;OL�;���;m�;�[�;��;���;h��;�{y;q:l;Ls_;�*S;�_G;�<;�/1;)�&;'�;��;�@	;���:���:��:f��:���:���:�З:VC�:��r:��V:C<:��":�d:-c�9�\�9�:�9/�b9��9�A�8���������q�ȣ���͹AN��_���q(��>��TS�eh�U|�# ��]���qۚ����[謺�ε�v�����Ǻh(Ѻ�ںy�亁F�R��f��SH�s�9���j�,��:]$���)���.��g3�y8��<�U�@��`E��I�ON���R�7�W�c�\��b��kg���l�Εr��Ax���}�FŁ�R����>���㉻�w��?����o��Yؓ��9��♘��  �  ��=%v=x$=(�=�x=�=]�=�a==ɟ =? =��<�<�T�<���<�<�i�<���<�B�<A��<�&�<ӗ�<��<�n�<E��<�/�<��<���<�(�<u�<���<��<�Z�<���<p��<%S�<ɫ�<7�<�d�<���< #�<���<z��<5�<��<���<!�<XP�<��<*��<3��<���<� �<D�<:h�<h��<���<~��<�
�<�3�<�X�<x�<H��<���<��<T��<4\�<%�<���<���<�<���<�<���<���<�@�<��<<��<��<�Y�<���<^��<��<W�<�%�<�7�<�?�<�=�<�1�<}�<���<�֫<!��<�~�<�P�<`%�<w��<�ڞ<d��<3��<�<���<���<`~�<�w�<�n�<�a�<O�<�6�<��<i�<vʁ<�;<{�z<�v<i"r<��m<�qi<w!e<��`<�\<3YX<g#T<r�O<��K<��G<IfC<E0?<��:<8�6<�U2<�-<�)<m&%<�� <~O<��<G�<YL<�<��<��<ڲ�;8��;' �;3D�;���;���;P7�;K��;DϿ;\�;�b�;0��;^�;<��;Q?�;T�;���;�Pz;+m;D`;��S;�H;¢<;��1;�';��;�;UH	;��:�.�:��:7�:η:>ܦ:
y�:���:6uo:�	S:_K8:!;:��:���9!0�9�ђ9��Y9V9ީ�8�p���J�����sp����{�˹f����~&�]L;�6P�V�d���x��E��f揺�T�������ƫ�贺����cǺ��кY�ںW庸�ﺃ������C�����^q�4�����E%�Ӏ*� �/�$J4�f�8� M=��A���E��:J���N�~/S� �W��\�$�a��?g�4�l�%/r�<�w�NL}�|h���"���ц�t��^
������}������~����d���  �  z�=9x=%=Q�=�v==��=�[=~� =Ė =�4 =$��<_��<�:�<^��<e��<jQ�<Q��<u.�<Т�<�<���<���<sh�<���<�.�<ӈ�<j��<l0�<B��<4��<��<�n�<���<��<�j�<���<@�<�w�<���<�/�<��<���<18�<3��<n��<��<�H�<wy�<ԣ�<��<��<��<{,�<#O�<�t�<���<\��<.��<7�<F�<�g�<��<O��<v��<c|�<Z�<�%�<w��<>��< !�<���<�'�<"��<s��<�X�<~��<���<5�<)o�<���<TϿ<���<��<,�<�:�<@�<Z;�<J,�<��<��<=ɫ<���<Rk�<-;�<l�<�<���<z��<7��<���<pw�<r�<�n�<�j�<[d�<�Y�<J�<84�<T�<���<с<�O<?�z<.�v<+Ir<�m<<�i<Qe<�a<S�\<6�X<,FT<�P<��K<E�G<�oC<S3?<6�:<*�6<=H2<�-<y)<%<?� <�%<-�<�b<�<��
<��<�<|U�;y�;g��;��;u_�;}��;��;Mr�;�ƿ;��;"r�;Ԩ;�G�;�ԙ;���;2U�;�S�;�{;��m;:�`;;�T;�H;�=;G2;�X';A;�;DE	;��:���: ��:X��:-�:�ե:iF�:$a�:~{l:��O:�5:��:U�:���9�ô9f��9�oQ9�{9�q8T���ب��^!�ōp��ݠ�y?ʹ�%��#"��#$�,�8�{�M���a�t�u�pЄ�f������D~���٪�z.������oǺ\�к�ںl;庀��0��aY�R7	�%���p��g� �4&�LR+�=Q0�H5���9�A�=��2B��eF���J�3�N��iS�MX���\��a�2!g��tl���q��Rw���|�o���̃��u�����歋��<��]Ð�/C��q����:���  �  ��=�y=&%=Z�=�t=�=��=�V=^� =�� =�, =��<��<�&�<{�<���<S>�<���<��<��<U�<H��<��<�b�<���<-�<���<���<�5�<t��<���<�+�<�}�<V��< &�<2|�<���<,�<���<k��<&9�<���<���<:�<���<���<C�<�A�<�p�<��<1��<��<���<�<�;�<j`�<���<ݳ�<���<V�<7�<[�<Dv�<���<��<�w�<�W�<b%�<���<ƌ�<(�<Ǵ�<�3�<Ħ�<��<j�<���<"�<�F�<`�<ɰ�<)ۿ<���<Z�<F0�<�<�<�?�<�8�<�'�<��<��<,��<H��<\�<�)�<���<qР<���<e��<�{�<Gn�<�f�<Kc�<�a�<�_�<�[�<RS�<�E�<�1�<�<6��<�Ձ<L^<�{<ιv<Rfr<�n<�i<�te<�)a<��\<U�X<`T<$P<��K<�G<�uC<�4?<��:<��6<r<2<�-<�d)<p�$<>x <�<~�<�;<��<&�
<�<��<��;�6�;�{�;���;�5�;Û�; �;a�;���;��;�{�;L�;�e�;���;���;��;͓�;J�{;�Nn;�wa;2
U;
I;Cv=;�M2;̊';�#;�;>	;FP�:M��:��:��:�A�:�:�S�:�P�:�%j:�hM:�|2:mj:�#:���9!{�9�0�9��J9��9pjm8�gO�\���I�"���p��v���Gɹ~��� ���"�xD7��K�|�_��s�Ҹ��w����.����*�������1����ƺ3�кG�ںLp�i\��������	�n�����Mq�)-!���&�}�+���0�L�5�x*:��w>�\�B���F���J��4O��S�"1X��\���a�g�UOl���q�
w��e|�}ျ����0��Ј��h�������������얕�����  �  i�=z=%=��=Is=�=׵=WS=_� =�� =h' =���<���<��<n�<���<E2�<a��<s�<���<��<�{�<
��<"_�<s��<�+�<���<��<=9�<I��<j��<�3�<7��<���<1�<8��<6��<�5�< ��<���<�>�<���<��<�:�<��<���<�<_=�<�j�<���<ҳ�<z��<���<[�<9/�<�S�<�{�<_��<���<��<{-�<�R�<Ao�<��<���<�t�<�U�<�$�<���<S��<X,�<���<v;�<���<;�<�u�<���<��<�Q�<j��<r��<m�<t�<W�<�2�<c=�<�>�<�6�<d$�<5�<&�<���<�<>R�<��<��<�à<���<o��<io�<�b�<#\�<�Y�<�Y�<Y�<V�<O�<sB�<�/�<��<��<J؁<�f<�{<��v<$xr<(n<��i<9�e<�?a<X�\<˱X<�oT<�0P< �K<@�G<IxC<�4?<6�:<H�6<�42<��-<�W)<d�$<�e <��<?�<�"<4�<~�
<�v<�h<5��;C�;V�;��;_�;���;1��;�T�;&��;J�;��;��;Yw�;�;�ђ;ǲ�;���;S�{;�n;�a;�VU;LI;A�=;,x2;F�';I4;�;P7	;-�:wM�:���:]��:�ε:�z�:Ϸ�:ա�:��h:��K:��0:��:n� :��9���9���93�F9��8��a8k4t�!��i�#��Rq��U��=�ȹ��{S���!�O76�pJ��}^��^r�
���ό������'������FV��������ƺl�к�ںɖ���,���/����	�����������!��'�`\,��Y1��6���:�a�>���B��
G��)K��`O�+�S��HX��]���a�Dg��9l�2�q�f�v��)|�����c��
��룈��=���ҍ��d��{�[~���
���  �  ��=Xo=�=?�=�h=�=î=8O=�� =�� =- =���<���<2�<��<���<�A�<Ȩ�<�<��<���<�^�<`��<w2�<.��<���<�P�<*��<���<�O�<[��<���<�C�<���<1��<>;�<���<���<�6�<���<#��<�/�<�~�<<��<3�<\R�<e��<���<��<��<�<�<�]�<}�<ܛ�<"��<���<��<� �<�C�<�d�<v��<ޙ�<��<E��<7��<���<gi�<y4�<���<��<�9�<���<oM�<���<1�<Β�<���<=9�<�<��<��<"�<�I�<fj�<V��<J��<��<ʜ�<��<���<pj�<�K�<�(�<��<�ݤ<׹�<ۘ�<�|�<�e�<wT�<AH�<2@�<7;�<f7�<k3�<v-�<�$�<v�<��<��<�Ճ<���<%/<��z<�v<�\r<Mn<��i<��e<�Ga<�]<�X<ۏT<�WP<< L< �G<��C<�r?<0;<�6<��2<�>.<��)<��%<�!!<��<�o<�%<��<n�<U�<�<C�;�n�;��;!�;�h�;V��;@�;���;)#�;К�;��;��;M�;6�;W��;ێ;���;|E�;�vu;��h;Ye\;�nP;��D;@�9;��.;
R$;�;~5;y�;2$�:ɢ�:l��:��:U��:y�:��:�ǂ:}h:%	M:�)3: �:��:�J�9�ֲ9l̊9LMG9M��8��08��JE��WB��0�������Yݹ������N-���A�XrV�Z�j���~��m��cV���1��*���ְ�õ���ĺ��κY5ٺ&�������w��c|�lQ�:#����с�P�$�9*�+H/��!4���8�OS=�`�A��$F�|�J�O���S��JX��#]� b�q<g��pl�ѷq��w�\^|��ـ�Ձ���&���ǈ��e��l��������)������oQ���  �  �=(o=�=_�=�h=5=r�=P=�� =� =�. ={��<���<'5�<��<���<�D�<���<��<?��<���<q`�<���<W3�<ǖ�<���<P�<���<���<9N�<{��<o��<�A�<1��<���<�8�<+��<R��<�4�<��<���<�.�<#~�< ��<'�<�R�<��<���<���<��<?�<W`�<��<���<E��<���<	�<�#�<�F�<�g�<ׄ�<��<ê�<���<1��<���<�i�<_4�<h��<H��<�8�<T��<[K�<���<�.�<��<���<n6�<\|�<`��<���< �<:H�<7i�<���<���<���<>��<ϔ�<��<�k�<�M�<+�<�<��<���<��<��<�h�<�W�<"K�<�B�<�=�<�9�<;5�<�.�<�%�<,�<N�<��<LՃ<-��<�,<\�z<�v<Xr<>n<��i<�e<{Ba<�]<��X<��T<�SP<�L<#�G<ͮC<|r?<�0;<Q�6<�2<�A.<n�)<Յ%<1&!<M�<�u<,<+�<��<�<��<�N�;gy�;X��;��;p�;���;D�;���;3$�;���;l�;���;�G�;'�;]ؕ;Ҏ;��;S;�;�au;��h;kR\;^P;]�D;*�9;!�.;�L$;y;�5;k�;�0�:}��: ��:���:�Ѳ:�6�:�<�:���:w�h:�jM:s�3:)1:`=:��9>r�9�T�9�CH9��8�38���⸣XB��<���Ƴ��ݹ���-����-��CB��V�k��6�����t|��8S��� ��{��ƺ��ĺ��κ4ٺ�㺳��8���Y��Nl�@�����4j���$�!*�C//�	4���8��==��A��F�Q}J���N�*�S��EX�!]�� b�/?g�wwl���q�aw��n|��※ڋ��V1���҈�$p���	��۞���1���Õ��V���  �  ��=xn=�=��=�i=�=\�=lR=~� =:� =�2 =��<���<�>�<���< ��<�M�<��<%�<���<Z��<�d�<;��<�5�<h��<K��<�O�< ��<��<UJ�<f��<U��<�:�<f��<Q��<30�<*��<���<-.�<i��<!��<G+�<�{�<��<-�<�S�<C��<%��<���<��<#E�<[g�<�<K��<k��<e��<r
�</-�<JO�<�o�<��<���<���<ǲ�<F��<���<�j�<>4�<D��<���<5�<���<�E�<���<�&�<���<��<�-�<t�<���<%��<i�<�C�<�e�<o��< ��<���<k��<���<F��<p�<�R�<?1�<K�<��<hŢ<Y��<N��<mr�<�`�<�S�<�J�<oD�<�?�<&:�<�2�<�(�<;�<R�<��<$ԃ<���<�%<�z<j�v<bJr<� n<V�i<�se<�1a<��\<��X<�T<�IP<�L<��G<��C<�q?<52;<��6<�2<.I.<��)<g�%<�3!<��<Æ<j><�<��<I�<�<Sq�;Ә�;���;S'�;���;���;�O�;���;�'�;��;/�;v��;�9�;$�;<��;���;�Ӈ;��;K!u;�kh;�\;}+P;��D;�z9;��.;�<$;[;_7;��;�U�:x��:��:�M�:F4�:먢:l��:䀃:�
j:ΛN:�4:�Z:�R:��9�=�9�ߌ9x�J9�M�8�98�~�I���EB��r��IL���o޹�U�m��b.��/C���W� l������yڶ���s��w-��s�����ĺ]�κ�-ٺط�J�� ���)��'A�6�������1$���$���)�`�.���3�r8�C�<��wA���E��VJ�P�N��vS�6X��]�a"b�Ig�j�l��q��;w��|�����G����Q��K􈻶���5(��t���cI���֕�-e���  �  ��=3m=2=?�=k=�=C�=V=� =�� =�8 =��<��<:M�<_��<���<�[�<���<�)�<��< �<�k�<���<�9�<���<���<�N�<��<b��<�C�<��<D��</�<�<T��<#�<}w�<��<r#�<Kz�<���<�%�<4x�<��<�<gU�<W��<���<��<�'�<�N�<Ur�<	��<ʴ�<���<��<&�<Y;�<�\�<�{�<ٖ�<���<���<���<��<���<l�<�3�<��<ݔ�<</�<��<�;�<s��<Y�<pz�<U��<��<�f�<���<4��<1�<T<�<O`�<�|�<��<蜵<埳<��<!��<�v�<[�<;�<v�<A��<Ӣ<���<��<��<�n�<a�<�V�<UO�<�H�<�A�<'9�<:-�<)�<��<o�<�у<İ�<�<�z<R�v<04r<��m<j�i<lYe<�a<1�\<͠X<�kT<Z9P<�L<j�G<�C<�o?<�3;<��6<�2<�T.<��)<��%<
I!<��<��<)[<p!<p�<(�<��<&��;b��;5�;PL�;,��;  �;�a�;���;�,�;��;��;��;�!�;�Μ; ��;]��;���;��;,�t;
h;��[;��O;�[D;�B9;a�.;�!$;(;^9;�;#��:�8�:uK�:���:�г:~[�:���:�[�:��k:�vP:��6:�%:�	:S#�9�	�9�V�9|�N9o��8�C8q���D�߸�3B�u㊹�+����߹V<�h����/���D�;VY�W�m�1���hڊ�~����Z��g���h���D��[	ź��κ7&ٺ���6S�S��]I�_����qx�~$�]��U $��^)�n.�xO3�\8��<��!A��E�mJ���N��SS�/ X��]��%b��[g���l��r�zw��|��)��dڃ������(��;ċ��X��琻8p�������}���  �  ��=Wk=u=��=�l=)=ŷ=�Z=�� =6� =3@ =���<9�<'`�<���<e�<�m�<T��<�8�<��<��<�t�<6��<8>�<���<#��<�L�<��<���<�:�<چ�<���<��<�n�<��<��<vf�<1��<;�<'n�<���<�<s�<��<]�<�V�<ߖ�<l��<��<~1�<�Z�<J��<���<$��<���<	
�<%,�<�M�<8n�<���<Ϥ�<r��<h��<���<F��<ԗ�<5m�<�2�<���<D��<$'�<a��<J/�<���<�	�<�h�<��<��<WU�<C��<���<��<+2�<�X�<qw�<��<"��<R��<���<Ǒ�<�~�<#e�<OG�<�&�<I�<��<=Ơ<;��<��<1��<Br�<|f�<!]�<�T�<�K�<�@�<�2�< �<�	�<f�<�΃<0��<�	<��z<hv<�r<�m<�|i<26e<��`<��\<��X<QT<$#P<5�K<��G<��C<7l?<~4;<��6<��2<wb.<�*<�%<d!<�<��<K�<0H<�<�<	�<���;k�;�8�;�z�;^��;S�;�v�;p��;�0�;2��;���;�u�;G �;Ǥ�;.h�;1Q�;�d�;���;�5t;��g;~C[;�kO;��C;v�8;�M.;�#;��;�6;�;#��:��:���:�q�: ��:�>�:4��:�t�:�(n:d�R:��8:�z :A>	:�#�9���9�b�9W�S9��9#O8ˠ�D1޸,rB�#���fg��řṭt��u1�/�F��t[���o����拺\����3��u����.�������Pź�Ϻ�&ٺ�u������5�ڨ��V������~&���#�$�(�H�-��2��~7�%$<���@�~?E���I�\oN��*S��X�u	]��/b��wg���l�qOr���w�N}�=d������Ɇ�)n��0	��ՙ��:"�������!��ҟ���  �  Ը=�h=@=��=�m=�=��=�_=�=�� =�H =,��<�%�<�u�<c��<�#�<��</��<sI�<^��<��</~�<��<�B�<
��<���<�I�<A��<���<�/�<6y�<���<��<�Z�<���< ��<cR�<i��<?�<]_�<���<��<&l�<���<��<�W�<R��<5��<�<L<�<�g�<!��<���<���<���<��<�A�<�b�<ہ�<���<���<���<'��<���<ݸ�<��<�m�<�0�<5��<��<�<���<��<��<9��<�S�<u��<4��<�@�<���<m��<���<�%�<O�<�p�<�<|��<I��<5��<���<��<Cp�<�T�<�6�<��<���<o۠<���<���<	��<���<Kx�<�l�<�a�<2V�<�H�<38�<�#�<p
�<|�<ʃ<棁<��~< �z<XIv<��q<q�m<�Si<Ze<a�`<��\<s^X<1T<+P<��K<v�G<.�C<�f?<4;<��6<C�2<%q.<�#*</�%<p�!<
4<�<j�<ht<�J<'.<9<M <�N�;2v�;��;���;�<�;o��;U��;'2�;㊺;��;�W�;�ף;bq�;F+�;�;J�;�W�;��s;T�f;��Z;��N;��C;�8;
.;a�#;��;-;�;��:g��:�V�:�#�:�k�:l@�: ��:���:��p:��U:��;:�"#:��:Z��9v��9Tʕ9�Y9�D9�S[81�ٷC�ܸ�C�Q���:
�����8�������3��H���]��r�UM���!�������7��p����Ⲻ-;��ЯźYQϺ!3ٺ	Y㺍�� ������^K����!~�������"��(�')-��2���6�2�;�_:@�B�D�s|I�`1N�l S�0�W�B]�Ab�8�g�m��r��3x�w�}�𩁻�g���������lZ��玻�h���ᓻ�U��Tɘ��  �  S�=�e=�=D�=�n=�=!�=�d=J	=j� =�Q =I��<�;�<���<c��<x:�<���<���<�Z�<7��<�#�<���<���<�F�<R��<X��<�E�<t��<���<O#�<�i�<��<���<zE�<'��<y��<s<�<���<z��<�N�<̬�<�	�<d�<���<4�<�W�<���<���<,�<;G�<�u�<@��<H��<f��<
�<q6�<�X�<�x�<���<Z��<���<`��<	��<���<#��<p��<�m�<�-�<l��<c�<��<G��<��<W|�<���<�<�<���<���<�)�<�m�<A��<-�<
�<D�<mh�<���<���<i��<���<R��<p��<�{�<c�<�G�<�*�<��<��<�מ<���<��<;��<���<�|�<o�<�`�<�P�<a=�<&�<H
�<��<dă<\��<��~<g�z<P'v<"�q<wm<�&i<Z�d<4�`<�f\<�6X<�T<��O<�K<��G<ۅC<�^?<�1;<��6<��2<l.<�7*<��%<~�!<GX<<��<�<	z<�\<�K<UF <{��;h��;���;I�;I[�;��;_��;�0�;`~�;KӲ;	5�;a��;�7�;y�;ÿ�;�Ɔ;6�;��r;�Af;�Z;XN;/C;�08;�-;g�#;��;�;��;U8�:*V�:1��:9��:L�:G�:�Ֆ:�:Ӛs:�yX:�>:}�%:L]:�v�9H��9�O�9�:_9��9��f8M�ͷ~�ܸ25D������������U�	������5��~K�W�`�hSu�?����z������X��苪�Y����ټ�c!ƺ��Ϻ�Lٺ�H�����Zs����p����dq�M��k+"��^'�\r,�(g1�9A6�
;�C�?�pD��)I���M���R�h�W��	]�Zb���g��Zm���r�
�x�FP~�����z���-s�����W����;�������&�����������  �  e�=,b=V=m�=+o=�=Q�=Ri=E=ִ =�Z =�  =�P�<̢�<��<�P�<i��<�
�<�k�<s��<J/�<��<���<�I�<���<��<�@�<���<l��<��<"Z�<Ԟ�<���<r/�<G}�<|��<�%�<}��<1��<>�<U��<���<0[�<e��<��<�V�<���<.��<c�<=Q�<t��<��<_��<��<�(�<�L�<�n�<t��<Ū�<~��<���<L��<���<���<{��<��<il�<*�<���<�u�<U�<&��<��<Fh�<���<3%�<�y�<���<��<�W�<���<Ծ<X	�</8�<j_�<D~�<}��<���<ѥ�<��<���<�<qp�<�W�<4=�<@"�<��<r�<�֜<���<)��<��<���<�{�<�j�<�W�<�A�<�'�<(	�<��<ƽ�<���<B�~<�ez<\v<c�q<�Km<&�h<��d<�o`<<:\<�X<J�S<i�O<��K<�G<�vC<oU?<�-;<��6<��2<�.<J*<&<��!<�{<�;<\<��<��<��<Cw<Hn <���;'��;	�;dA�;Xv�;ݯ�;|��;�+�;n�;-��;��;�w�;���;���;4q�;�q�;�Q;�5r;��e;snY;N�M;c�B;8�7;�Z-;�J#;х;[;t�;�Z�:Ȥ�:�W�:�}�:Z�:�F�:���:,G�:�Sv:�N[:ArA:J�(:��:��9���9���9`nd9IL9G�p8�Fŷ�ݸ'�E��=�����ue� c���!�r>8�� N�zc��2x��#��9ݏ�"M��*��������������1�ƺ��Ϻ5uٺ�H㺙f�d����1���f�Jq�`��O4�{!�p�&�e�+�+�0���5��x:�D?��D��H���M�=�R��W�]��zb�,h�Ϧm��^s��y���~��E������͇��w��U����������m���͖�L+���  �  x�=�^=�=-�=1o==��=Am=�=p� =Yb =�	 =Cd�<#��<��<�d�<w��<@�<�z�<
��<99�<_��<��<�K�<��<
��<v;�<ق�< ��<	�<�J�<��<��<��<�g�<���<��<`l�<���<u-�<P��<f��< R�<��<��<NU�<���<���<s!�<�Y�<ˍ�<��<���<��<;<�<4a�<a��<0��<��<���<���<���<���<���<���<���<pj�<�%�<���<gl�<<��<�x�<���<�T�<���<��<�b�<���<}��<EC�<���<7þ<&��<~,�<AV�<�w�<I��<石<Ѧ�<���<U��<��<;|�<6f�<�M�<�4�<��<��<R�<՚<9��<���<���<���<s�<a]�<�D�<6(�<6�<`�<�<���<=�~<WHz<$�u<Iq<q"m<��h<��d<8D`<a\<��W<��S<��O<�K<WG<WgC<�J?<A(;<a�6<j�2<��.<�Y*<6&<6�!<b�<`<�)<��<5�<M�<�<�� <��;(�;k?�;9b�;@��;���;���;#�;�[�;��;M�;EG�;3��;�]�;�&�;H!�;��~;Ɍq;v�d;��X;�3M;�B;�V7;�-;�#;�U;��;��;�o�:!��:��:��:uٷ:]+�:��:�n�:7�x:��]:�D:C++:�>:W@�9#j�9/��9'�h9-�9'x8�\���i޸ڳG�:ʐ�O��36�����#�!�:���P�� f���z�[���,������?���ۈ���[�� 2��x$Ǻ�Gк��ٺ�U�fJ�p����� ��F�(�����Q�O���� ��&�'+� 0��5���9��>�0�C���H��M���R�n�W��&]�͟b�x;h�x�m���s���y�Ud�����lc���#���Ί��d���䏻�R��򲔻%	���\���  �  �=[=z=Ͽ=�n=�=��=Np=�=�� =�h =: =�t�<g��<�<�u�<���<�*�<C��<h��<RA�<��<q��<�L�<��<���<A6�<t{�<k��<���<�<�<�}�<���<<�<�T�<|��<���<�Z�<d��<��<ǃ�<���<�I�<ŧ�<o �<JS�<���<���< &�<�`�<)��<s��<H��<$�<�L�<sr�<���<��<{��<���<2��<��<���<Y��<���<{��<*h�<!�<L��<�c�<I��<�k�<���<D�<��<u��<�N�<ǝ�<��<1�<u�<j��<{�<�!�<�M�<yq�<��<읳<��<��<��<_��<<r�<�[�<�D�<,�<H�<���<��<nϘ<���<��<Ꮢ<�y�<�a�<�F�<#(�<��<�܅<v��<��<��~<Y.z<T�u<�]q<�l<��h<�\d<�`<u�[<}�W<��S<o�O<~K<_lG<�XC<�@?<<";<��6<J�2<}�.<�e*<�+&<*�!<Ե<a~<rK<�<�<��<J�<� <�S�;�T�;�b�;�{�;Ԝ�;I��; ��;S�;J�;f��;�Ī;��;%��;�"�;v�;_څ;�~;�p;�]d;�HX;h�L;�A;��6;��,;��";G(;��;�;(w�:
�:��:��:ns�:8�:�:!h�:��z:M`:'5F:�J-:/4:k��9_�9���9Ϡl9��9�?}8�ʾ��'�ئI�&A���W��������%���<���R�pth��P}����LT���������\g������ξ�͞Ǻi�кu�ٺ\j㺐<�R��!� �U�,N���#���R ��y%���*���/�К4���9�i>�
pC��iH�sM���R��W��:]���b��ph�~:n��t���y�T��Ԃ�����o�����&���`-��$���A;>��8����  �  A�=5X=o=��=zn=5= �=|r=�=�� =�m =� =ʀ�<O��<.+�<���<���<�5�<���<��<'G�<��<���<M�<ѝ�<��<�1�<du�<õ�<2��<%2�<�q�<���<��<�E�<���<���<�L�<���<��<�y�<���<�B�<���<���<ZQ�<R��<<��<*)�<�e�<��<
��<��<�/�<LY�<g�<���<W��<���<���<���<���<���<v��<"��<��<f�<M�<���<\�<���<a�<���<�6�<���<w��<:?�<U��<2��<�"�<h�<Ȩ�<H�<\�<�F�<,l�<���<���<���<���<x��<���<��<{�<�f�<IP�<9�<U!�<�	�<��<�ژ<Ė<f��<���<w~�<�d�<H�<�'�<��<<م<��<�x�<;�~<�z<��u<�Cq<��l<^�h<�>d<B `<��[<��W<ˎS<�zO<�kK</]G<�LC<�7?<�;<��6<��2<��.<�n*<08&<z "<��<C�<^d<w8<<;�<?�<�� <�{�;�u�;�|�;
��;I��;��;~��;c�;o:�;ik�;t��;���; d�;W��;ذ�;���;3�};�p;2�c;��W;-TL;;FA;�6;�r,;��";� ;ϯ;I�;�t�:�$�:�A�:"��:��:�s�:d��:�"�:e|:�a:X�G:'�.:��:�_�9ו�9-ȣ9�8o9$�9�N�8F������)UK���������������b*'�>�ɊT�m>j��*�����7��2t���^��������#L���Ⱥ��к�ں���Q:�1��ϰ �f��+�5N������]���%�**��9/�@4��?9�}=>�:<C�AEH��\M��R���W�M]���b��h��sn��\t��Nz�I����yㅻ)����V��uꍻ�e���ʒ�r��Fh��묙��  �  �=RV==��=n=`=��=�s=�=U� =�p =O =~��<z��<�3�<���<��<p<�<n��<���<�J�<W��<���<6M�<ٜ�<��<�.�<hq�<��<E��<J+�<�i�<��<���<l<�<3��<5��<D�<{��<=�<ds�<6��<�>�<��<x��<�O�<���<���<	+�<�h�<��<I��<��<�6�<a�<���<թ�<3��<?��<1��<��<���<���<M��<���<{��<pd�<��<��<�W�<���<rZ�<P��<W.�<���<���<T5�<h��<���<��<�_�<_��<�ݼ<��<uB�<�h�<��<���<]��<h��<~��<���<d��<���<m�<�W�<A�<�)�<��<���<��<7ʖ<���<|��<j��<uf�<�H�<)'�<E�<�օ<r��<Dt�<(|~<�z<ԝu<3q<�l<Nwh<q+d<�_<��[<��W<"S<:mO<�_K<�SG<EC<.2?<;<�6<�2<`�.<�s*<�?&<b
"<��<q�<$t<<I<P#<�	<�<� <��;���;��;H��;���;��;'��;�	�;�/�;�\�;t��;X�;�I�;"֓;)��;���;�[};�;p;��c;g�W;�L;�A;�x6;J,;�r";��;�;
�;Kr�:�1�:b�:��:C'�:Tɩ:@�:���:%}}:�b:,�H:A�/:}�:���9���9P֤9��p9f�9L�8c��C8�U{L�-[���ù}�l��U(�8!?���U�!hk��,���3��7ʓ�����Oޥ�4���[��z����CȺHѺ*3ں#���9� ���� ����H�
�!��S���)����$�W�)���.��4��9�Q>��C��.H��OM���R�W�W�|Z]���b�M�h�ݗn�k�t��z��:��Y)������Έ��|��K��K���6쒻=��Â���Ù��  �  �=�U=�
=]�=n=r=�=It=~=;� =�q =w =��<��<E6�<V��<���<�>�<r��<e��<�K�<$��<.��<OM�<���<U��<�-�<�o�<��<,��<�(�<�f�<2��<���<S9�<5��<��<A�<���<�	�<<q�<9��<�<�<��<���<WO�<��<��<�+�<�i�<���</��<�
�</9�<�c�<K��<}��<���<���<J��< ��<l �<���<���<���<d��<�c�<��<��<?V�<���<0X�<���<q+�<���<e��</2�<4��<O��<��<�\�<ើ<�ۼ<��<�@�<�g�<<��<	��<R��<���<&��<ٟ�<�<y��<7o�<Z�<�C�<V,�<m�<W��<Q�<U̖<h��<ߛ�<i��<�f�<�H�<
'�<� �<�Յ<1��<�r�<x~<2z<��u<^-q<�l<�ph<n%d<��_<~�[<ɒW<�yS<�hO<�[K<PG<;BC<:0?<�;<��6<T�2<*�.<�u*<MB&<"<	�<*�<Uy<�N<�(<S	<6�<�� <w��;��;���;��;M��;��;K��;��;�,�;�W�;���;lڢ;A�;�˓;"��;�t�;�C};�$p;��c;��W;�K;>�@;�g6;�:,;=f";U�;�;#�;-r�:@5�:l�:��:�>�:]�:v�:J��:k�}:�c:=;I:q/0:U�:^B :m�9K6�9�^q9��9H�8,k��3��&�L������pùƚ����_(��y?���U�X�k��\���d��b���++���	������3��$���o[Ⱥ�*Ѻ�>ں����8�k���� �
��D�
��/B�Lo����W�$�D�)�N�.��3���8�{>��C�'H�BLM�P�R���W�j_]� c���h�S�n�ϙt���z��D���4������ۈ��������~��������G��ǋ��̙��  �  �=RV==��=n=`=��=�s=�=U� =�p =O =~��<z��<�3�<���<��<p<�<n��<���<�J�<W��<���<6M�<ٜ�<��<�.�<hq�<��<E��<J+�<�i�<��<���<l<�<3��<5��<D�<{��<=�<ds�<6��<�>�<��<x��<�O�<���<���<	+�<�h�<��<I��<��<�6�<a�<���<թ�<3��<?��<1��<��<���<���<M��<���<{��<pd�<��<��<�W�<���<rZ�<P��<W.�<���<���<T5�<h��<���<��<�_�<_��<�ݼ<��<uB�<�h�<��<���<^��<i��<~��<���<d��<���<m�<�W�<A�<�)�<��<���<��<7ʖ<���<{��<j��<tf�<�H�<('�<E�<�օ<r��<Dt�<'|~<�z<ԝu<3q<�l<Nwh<q+d<�_<��[<��W<"S<:mO<�_K<�SG<EC<.2?<;<�6<�2<a�.<�s*<�?&<b
"<��<r�<%t<=I<P#<�	<�<� <��;���;��;G��;���;��;%��;�	�;�/�;�\�;s��;W�;�I�;!֓;(��;���;�[};�;p;��c;f�W;�L;�A;�x6;J,;�r";��;�;
�;Jr�:�1�:b�:��:C'�:Tɩ:@�:���:%}}:�b:,�H:A�/:}�:���9���9P֤9��p9f�9L�8c��C8�U{L�-[���ù}�l��U(�8!?���U�!hk��,���3��7ʓ�����Oޥ�4���[��z����CȺHѺ*3ں#���9� ���� ����H�
�!��S���)����$�W�)���.��4��9�Q>��C��.H��OM���R�W�W�|Z]���b�M�h�ݗn�k�t��z��:��Y)������Έ��|��K��K���6쒻=��Â���Ù��  �  A�=5X=o=��=zn=5= �=|r=�=�� =�m =� =ʀ�<O��<.+�<���<���<�5�<���<��<'G�<��<���<M�<ѝ�<��<�1�<du�<õ�<2��<%2�<�q�<���<��<�E�<���<���<�L�<���<��<�y�<���<�B�<���<���<ZQ�<R��<<��<*)�<�e�<��<
��<��<�/�<LY�<g�<���<W��<���<���<���<���<���<v��<"��<��<f�<M�<���<\�<���<a�<���<�6�<���<x��<;?�<U��<3��<�"�<h�<Ȩ�<H�<\�<�F�<,l�<���<���<���<���<y��<���<��<{�<�f�<JP�<9�<U!�<�	�<��<�ژ<Ė<f��<���<w~�<�d�<H�<�'�<��<<م<��<�x�<:�~<�z<��u<�Cq<��l<^�h<�>d<B `<��[<��W<̎S<�zO<�kK<0]G<�LC<�7?<�;<��6<��2<��.<�n*<08&<{ "<��<C�<^d<w8<<;�<?�<�� <{�;�u�;�|�;��;G��;��;{��;a�;m:�;gk�;q��;���;�c�;U��;ְ�;���;0�};�p;/�c;��W;+TL;:FA;�6;�r,;��";� ;ί;H�;�t�:�$�:�A�:"��:��:�s�:d��:�"�:e|:�a:X�G:'�.:��:�_�9ו�9-ȣ9�8o9$�9�N�8F������)UK���������������b*'�>�ɊT�m>j��*�����7��2t���^��������#L���Ⱥ��к�ں���Q:�1��ϰ �f��+�5N������]���%�**��9/�@4��?9�}=>�:<C�AEH��\M��R���W�M]���b��h��sn��\t��Nz�I����yㅻ)����V��uꍻ�e���ʒ�r��Fh��묙��  �  �=[=z=Ͽ=�n=�=��=Np=�=�� =�h =: =�t�<g��<�<�u�<���<�*�<C��<h��<RA�<��<q��<�L�<��<���<A6�<t{�<k��<���<�<�<�}�<���<<�<�T�<|��<���<�Z�<d��<��<ǃ�<���<�I�<ŧ�<o �<JS�<���<���< &�<�`�<)��<s��<H��<$�<�L�<sr�<���<��<{��<���<2��<��<���<Y��<���<{��<*h�<!�<L��<�c�<J��<�k�<���<D�<��<v��<�N�<ȝ�<��<1�<u�<k��<|�<�!�<�M�<zq�<��<읳<��<��<��<`��<<r�<�[�<�D�<,�<H�<���<��<nϘ<���<��<���<�y�<�a�<�F�<"(�<��<�܅<u��<��<��~<W.z<S�u<�]q<�l<��h<�\d<�`<u�[<}�W<��S<p�O<~K<`lG<�XC<�@?<=";<��6<K�2<~�.<�e*<�+&<+�!<յ<a~<sK<�<�<��<J�<� <�S�;�T�;�b�;�{�;ќ�;F��;���;O�;J�;b��;�Ī;��;"��;�"�;t�;\څ;�~;�p;�]d;�HX;e�L;�A;��6;��,;��";F(;��;~�;'w�:
�:��:��:ms�:8�:�:!h�:��z:M`:'5F:�J-:.4:k��9_�9���9Ϡl9��9�?}8�ʾ��'�ئI�&A���W��������%���<���R�pth��P}����LT���������\g������ξ�͞Ǻi�кu�ٺ\j㺐<�R��!� �U�,N���#���R ��y%���*���/�К4���9�i>�
pC��iH�sM���R��W��:]���b��ph�~:n��t���y�T��Ԃ�����o�����&���`-��$���A;>��8����  �  x�=�^=�=-�=1o==��=Am=�=p� =Yb =�	 =Cd�<#��<��<�d�<w��<@�<�z�<
��<99�<_��<��<�K�<��<
��<v;�<ق�< ��<	�<�J�<��<��<��<�g�<���<��<`l�<���<u-�<P��<f��< R�<��<��<NU�<���<���<s!�<�Y�<ˍ�<��<���<��<;<�<4a�<a��<0��<��<���<���<���<���<���<���<���<pj�<�%�<���<gl�<<��<�x�<���<�T�<���<��<�b�<���<~��<FC�<���<8þ<'��<,�<BV�<�w�<J��<蟳<Ҧ�<���<U��<��<<|�<7f�<�M�<�4�<��<��<R�<՚<8��<���<���<���<s�<`]�<�D�<5(�<5�<_�<�<���<;�~<VHz<#�u<Hq<q"m<��h<��d<8D`<b\<��W<��S<��O<�K<YG<YgC<�J?<C(;<c�6<l�2<�.<�Y*<7&<8�!<c�<`<�)<��<5�<M�<�<�� <��;(�;h?�;6b�;<��;���;���;#�;�[�;���;I�;AG�;/��;�]�;~&�;F!�;��~;Ōq;r�d;��X;�3M;�B;�V7;�-;�#;�U;��;��;�o�: ��:��:��:uٷ:]+�:��:�n�:7�x:��]:�D:C++:�>:V@�9#j�9/��9'�h9-�9'x8�\���i޸ڳG�:ʐ�O��36�����#�!�:���P�� f���z�[���,������?���ۈ���[�� 2��x$Ǻ�Gк��ٺ�U�fJ�p����� ��F�(�����Q�O���� ��&�'+� 0��5���9��>�0�C���H��M���R�n�W��&]�͟b�x;h�x�m���s���y�Ud�����lc���#���Ί��d���䏻�R��򲔻%	���\���  �  e�=,b=V=m�=+o=�=Q�=Ri=E=ִ =�Z =�  =�P�<̢�<��<�P�<i��<�
�<�k�<s��<J/�<��<���<�I�<���<��<�@�<���<l��<��<"Z�<Ԟ�<���<r/�<G}�<|��<�%�<}��<1��<>�<U��<���<0[�<e��<��<�V�<���<.��<c�<=Q�<t��<��<_��<��<�(�<�L�<�n�<t��<Ū�<~��<���<L��<���<���<{��<��<il�<*�<���<�u�<U�<&��<��<Fh�<���<4%�<�y�<���<��<�W�<���<Ծ<Y	�<08�<k_�<E~�<~��<���<ҥ�<��<���<���<rp�<�W�<5=�<A"�<��<r�<�֜<���<(��<~��<���<�{�<�j�<�W�<�A�<�'�<'	�<��<Ž�<���<@�~<~ez<[v<c�q<�Km<&�h<��d<�o`<<:\<�X<K�S<j�O<��K<�G<�vC<qU?<�-;<��6<��2<�.<J*<&<��!<�{<�;<]<��<��<��<Bw<Gn <���;$��;�;`A�;Tv�;ٯ�;x��;�+�;n�;(��;��;�w�;���;���;0q�;�q�;�Q;�5r;��e;pnY;J�M;a�B;5�7;�Z-;�J#;υ;Z;s�;�Z�:Ǥ�:�W�:�}�:Y�:�F�:���:+G�:�Sv:�N[:ArA:J�(:��:��9���9���9`nd9IL9G�p8�Fŷ�ݸ'�E��=�����ue� c���!�r>8�� N�zc��2x��#��9ݏ�"M��*��������������1�ƺ��Ϻ5uٺ�H㺙f�d����1���f�Jq�`��O4�{!�p�&�e�+�+�0���5��x:�D?��D��H���M�=�R��W�]��zb�,h�Ϧm��^s��y���~��E������͇��w��U����������m���͖�L+���  �  S�=�e=�=D�=�n=�=!�=�d=J	=j� =�Q =I��<�;�<���<c��<x:�<���<���<�Z�<7��<�#�<���<���<�F�<R��<X��<�E�<t��<���<O#�<�i�<��<���<zE�<'��<y��<s<�<���<z��<�N�<̬�<�	�<d�<���<4�<�W�<���<���<,�<;G�<�u�<@��<H��<f��<
�<q6�<�X�<�x�<���<Z��<���<`��<	��<���<#��<p��<�m�<�-�<l��<c�<��<H��<��<W|�<���<�<�<���<���<�)�<�m�<B��<.�<�<D�<nh�<���<���<j��<���<S��<q��<�{�<c�<�G�<�*�<��<��<�מ<���<��<;��<���<�|�<o�<�`�<�P�<`=�<&�<G
�<��<că<[��<��~<f�z<N'v<!�q<wm<�&i<Z�d<4�`<�f\<�6X<�T<��O<�K<��G<݅C<�^?<�1;<��6<��2<n.<�7*<�%<��!<HX<<��<�<	z<�\<�K<TF <x��;e��;���;E�;E[�;��;Z��;�0�;\~�;FӲ;5�;\��;�7�;u�;���;�Ɔ;3�;}�r;�Af;�Z;XN;,C;�08;�-;e�#;��;�;��;T8�:)V�:0��:8��:L�:G�:�Ֆ:�:Ӛs:�yX:�>:}�%:K]:�v�9H��9�O�9�:_9��9��f8M�ͷ~�ܸ25D������������U�	������5��~K�W�`�hSu�?����z������X��苪�Y����ټ�c!ƺ��Ϻ�Lٺ�H�����Zs����p����dq�M��k+"��^'�\r,�(g1�9A6�
;�C�?�pD��)I���M���R�h�W��	]�Zb���g��Zm���r�
�x�FP~�����z���-s�����W����;�������&�����������  �  Ը=�h=@=��=�m=�=��=�_=�=�� =�H =,��<�%�<�u�<c��<�#�<��</��<sI�<^��<��</~�<��<�B�<
��<���<�I�<A��<���<�/�<6y�<���<��<�Z�<���< ��<cR�<i��<?�<]_�<���<��<&l�<���<��<�W�<R��<5��<�<L<�<�g�<!��<���<���<���<��<�A�<�b�<ہ�<���<���<���<'��<���<ݸ�<��<�m�<�0�<5��<��<�<���<��<��<:��<�S�<v��<5��<�@�<���<n��<���<�%�<O�<�p�<���<}��<J��<6��<���<��<Cp�<�T�<�6�<��<���<o۠<���<���<	��<���<Jx�<�l�<�a�<2V�<�H�<28�<�#�<o
�<{�<ʃ<壁<��~<�z<WIv<��q<p�m<�Si<Ze<a�`<��\<t^X<1T<,P<��K<x�G<0�C<�f?<4;<��6<E�2<'q.<�#*<0�%<r�!<4<�<j�<it<�J<&.<8<L <�N�;/v�;��;���;�<�;k��;Q��;#2�;ފ�;��;�W�;�ף;^q�;B+�;�;G�;�W�;��s;O�f;�Z;��N;��C;�8;.;_�#;��;-;�;��:f��:�V�:�#�:�k�:k@�: ��:���:��p:��U:��;:�"#:��:Z��9v��9Tʕ9�Y9�D9�S[81�ٷC�ܸ�C�Q���:
�����8�������3��H���]��r�UM���!�������7��p����Ⲻ-;��ЯźYQϺ!3ٺ	Y㺍�� ������^K����!~�������"��(�')-��2���6�2�;�_:@�B�D�s|I�`1N�l S�0�W�B]�Ab�8�g�m��r��3x�w�}�𩁻�g���������lZ��玻�h���ᓻ�U��Tɘ��  �  ��=Wk=u=��=�l=)=ŷ=�Z=�� =6� =3@ =���<9�<'`�<���<e�<�m�<T��<�8�<��<��<�t�<6��<8>�<���<#��<�L�<��<���<�:�<چ�<���<��<�n�<��<��<vf�<1��<;�<'n�<���<�<s�<��<]�<�V�<ߖ�<l��<��<~1�<�Z�<J��<���<$��<���<	
�<%,�<�M�<8n�<���<Ϥ�<r��<h��<���<F��<ԗ�<5m�<�2�<���<D��<$'�<b��<J/�<���<�	�<�h�<��<��<WU�<D��<���<��<,2�<�X�<rw�<��<#��<S��<���<ȑ�<�~�<$e�<OG�<�&�<J�<��<=Ơ<;��<��<1��<Ar�<{f�< ]�<�T�<�K�<�@�<�2�<~ �<�	�<e�<�΃<0��<�	<��z<hv<�r<�m<�|i<26e<��`<��\<��X<QT<%#P<6�K<��G<��C<9l?<�4;<��6<��2<xb.<�*<�%<d!<�<��<L�<0H<�<�<	�<���;i�;�8�;�z�;[��;O�;�v�;l��;�0�;.��;���;�u�;C �;ä�;+h�;-Q�;�d�;���;�5t;}�g;zC[;�kO;��C;t�8;�M.;�#;��;�6;�;"��:��:���:�q�:���:�>�:4��:�t�:�(n:d�R:��8:�z :A>	:�#�9���9�b�9W�S9��9#O8ˠ�D1޸,rB�#���fg��řṭt��u1�/�F��t[���o����拺\����3��u����.�������Pź�Ϻ�&ٺ�u������5�ڨ��V������~&���#�$�(�H�-��2��~7�%$<���@�~?E���I�\oN��*S��X�u	]��/b��wg���l�qOr���w�N}�=d������Ɇ�)n��0	��ՙ��:"�������!��ҟ���  �  ��=3m=2=?�=k=�=C�=V=� =�� =�8 =��<��<:M�<_��<���<�[�<���<�)�<��< �<�k�<���<�9�<���<���<�N�<��<b��<�C�<��<D��</�<�<T��<#�<}w�<��<r#�<Kz�<���<�%�<4x�<��<�<gU�<W��<���<��<�'�<�N�<Ur�<	��<ʴ�<���<��<&�<Y;�<�\�<�{�<ٖ�<���<���<���<��<���<l�<�3�<��<ݔ�<</�<��<�;�<s��<Z�<pz�<V��<  �<�f�<���<5��<2�<U<�<P`�<�|�<��<霵<柳<��<"��<�v�<[�<;�<v�<A��<Ӣ<���<��<��<�n�<a�<�V�<TO�<�H�<�A�<'9�<9-�<)�<��<n�<�у<ð�<�<~�z<Q�v<04r<��m<j�i<lYe<�a<1�\<͠X<�kT<[9P<�L<k�G<�C<�o?<�3;<��6<�2<�T.<��)<��%<I!<��<��<)[<p!<p�<(�<��<%��;`��;3�;ML�;)��; �;�a�;���;�,�;��;��;��;�!�;�Μ;���;[��;��;��;)�t;
h;��[;��O;�[D;�B9;`�.;�!$;';]9;�;"��:�8�:tK�:���:�г:}[�:���:�[�:��k:�vP:��6:�%:�	:S#�9�	�9�V�9|�N9o��8�C8q���D�߸�3B�u㊹�+����߹V<�h����/���D�;VY�W�m�1���hڊ�~����Z��g���h���D��[	ź��κ7&ٺ���6S�S��]I�_����qx�~$�]��U $��^)�n.�xO3�\8��<��!A��E�mJ���N��SS�/ X��]��%b��[g���l��r�zw��|��)��dڃ������(��;ċ��X��琻8p�������}���  �  ��=xn=�=��=�i=�=\�=lR=~� =:� =�2 =��<���<�>�<���< ��<�M�<��<%�<���<Z��<�d�<;��<�5�<h��<K��<�O�< ��<��<UJ�<f��<U��<�:�<f��<Q��<30�<*��<���<-.�<i��<!��<G+�<�{�<��<-�<�S�<C��<%��<���<��<#E�<[g�<�<K��<k��<e��<r
�</-�<JO�<�o�<��<���<���<ǲ�<F��<���<�j�<>4�<D��<���<5�<���<�E�<���<�&�<���<��<�-�<t�<���<%��<i�<�C�<�e�<p��<��<���<l��<���<F��<p�<�R�<@1�<L�<��<hŢ<Y��<N��<mr�<�`�<�S�<�J�<oD�<�?�<%:�<�2�<�(�<;�<R�<��<$ԃ<���<�%<�z<i�v<bJr<� n<V�i<�se<�1a<��\<��X<�T<�IP<�L<��G<��C<�q?<62;<��6<��2</I.<��)<h�%<�3!<��<Ć<j><�<��<I�<�<Rq�;Ҙ�;���;Q'�;���;���;�O�;���;�'�;��;-�;t��;�9�;"�;:��;���;�Ӈ;��;H!u;�kh;�\;{+P;��D;�z9;��.;�<$;Z;_7;��;�U�:x��:��:�M�:E4�:먢:l��:䀃:�
j:ΛN:�4:�Z:�R:��9�=�9�ߌ9x�J9�M�8�98�~�I���EB��r��IL���o޹�U�m��b.��/C���W� l������yڶ���s��w-��s�����ĺ]�κ�-ٺط�J�� ���)��'A�6�������1$���$���)�`�.���3�r8�C�<��wA���E��VJ�P�N��vS�6X��]�a"b�Ig�j�l��q��;w��|�����G����Q��K􈻶���5(��t���cI���֕�-e���  �  �=(o=�=_�=�h=5=r�=P=�� =� =�. ={��<���<'5�<��<���<�D�<���<��<?��<���<q`�<���<W3�<ǖ�<���<P�<���<���<9N�<{��<o��<�A�<1��<���<�8�<+��<R��<�4�<��<���<�.�<#~�< ��<'�<�R�<��<���<���<��<?�<W`�<��<���<E��<���<	�<�#�<�F�<�g�<ׄ�<��<ê�<���<1��<���<�i�<_4�<h��<H��<�8�<T��<\K�<���<�.�<��<���<n6�<\|�<`��<���< �<:H�<7i�<���<���<���<?��<ϔ�<��<�k�<�M�<+�<�<��<���<��<��<�h�<�W�<"K�<�B�<�=�<�9�<;5�<�.�<�%�<+�<M�<��<LՃ<-��<�,<\�z<
�v<Xr<>n<��i<�e<{Ba<�]<��X<��T<�SP<�L<#�G<ήC<|r?<�0;<Q�6<��2<�A.<o�)<օ%<2&!<M�<�u<,<+�<��<�<��<�N�;gy�;W��;��;p�;���;
D�;���;2$�;���;j�;���;�G�;&�;\ؕ;Ҏ;��;R;�;�au;��h;jR\;^P;\�D;)�9; �.;�L$;x;�5;k�;�0�:|��: ��:���:�Ѳ:�6�:�<�:���:w�h:�jM:s�3:)1:`=:��9>r�9�T�9�CH9��8�38���⸣XB��<���Ƴ��ݹ���-����-��CB��V�k��6�����t|��8S��� ��{��ƺ��ĺ��κ4ٺ�㺳��8���Y��Nl�@�����4j���$�!*�C//�	4���8��==��A��F�Q}J���N�*�S��EX�!]�� b�/?g�wwl���q�aw��n|��※ڋ��V1���҈�$p���	��۞���1���Õ��V���  �  ɺ=	f= =ĸ=�_='=�=�K=i� =8� =p1 =���<���<B�<^��<j��<{J�<���<��<�u�<���<�B�<k��<V	�<�g�<-��<�<p�<���<��<Mc�<h��<��<�P�<,��<��<V@�<̐�<��<�0�<��<���<+�<D^�<]��<x��<n�<�K�<�y�<��<���<���<��<'�<D�<�`�<J}�<���<���<?��<���<��<h��<���<^��<���<N��<QR�<8�<���<�T�<���<ck�<���<(U�<���<��<bj�<���<���<�4�<2i�<���<伺<�۸<3�<��<�
�<�<�<���<��<!ͨ<泦<���<��<�g�<�R�<A�<�2�<1(�< �<��<D�<��<�<X��<Z��<�߇<�˅<���<l��<�~<�z<�v<,Cr<|n<��i<`�e<DPa<�]<�X<��T<^~P<�ML<!H<��C<;�?<�};<V@7</�2<B�.<Nm*<�!&<A�!<L�<�O<l<U�<��<�<9�<�� <޴�;N��;�J�;ά�;��;���;��; ��;��;b��;�R�;�;�;�Ҙ;��;��;�w�;y�{;co;!#c;s>W;��K;)�@;Ǯ5;(+;�� ;��;�B;��;��:� �:Rf�:J�:��:B��:"h�:^��:�ug:B�L:�3:sd:�N:q<�9�'�9M�9��:9�'�8�Q�7Ey��W�g�$����ȹ��*��e$�6y9�dN��c���w�Q���!���2���8��8@��4R���yº��̺y4׺���j�캧����|�](�������%�Z���#��Y(�)w-�n2�TB7���;��@��DE���I���N��SS�{-X�m"]��1b�!Zg���l�#�q�4w��|���@����E��wꈻ����c)��kĐ�^�����������  �  n�=�e==ܸ=�_=o=e�=0L=3� =� =d2 =���<���<`D�<���<���<�L�<���<��<�w�<&��<D�<=��<�	�<<h�<C��<��<�o�<���<w�<�a�<ݰ�<���<�N�<)��<��<_>�<��<f��<d/�<o~�<���<��<^�<R��<���<��<rL�<�z�<=��<t��<l��<�
�<)�<aF�<4c�<��<���<���<@��<X��<��<���<���<��<��<���<9R�<�
�<��<�S�<���<�i�<���<,S�<���<��<<h�<q��<���<�2�<�g�<b��<���<C۸<��<��<�<��<��<���<?�<�Ψ<���<���<��<@j�<,U�<oC�<55�<B*�< "�<��<��<��<�<���<���<��<�˅<F��<Ǚ�<�~<y�z<�~v<�?r<� n<��i<7�e<9La<�]<v�X<��T<�{P<�KL<�H<F�C<��?<�};<A7<G�2<�.<�o*<�$&<��!<(�<T<
<!�< �<��<ս<�� <���;U��;XQ�;̱�;8�;���;��;ډ�;��;+��;�O�;
�;�ܟ;�̘;�ݑ;�;�o�;��{;�So;hc;�1W;=�K;�}@;��5;�#+;�� ;��;pE;r�;��:��:�|�:�d�:�ׯ:oߟ:���:D݁:+�g:QM:<�3:��:�:���9���9}_�9�g;9c��8`�7ϣx�hZ��2g��G��oɹk��Y��$�E�9�}�N��`c���w��$���?���K��8O��LR��\_��<�º!�̺�3׺��ẳ�������s������mw�r�כ��#��G(��d-��[2��17�4�;�:�@��7E���I�ʋN��NS�f*X�� ]�j2b�F\g�ۚl�!�q�Y>w���|��������lM���򈻕���&1��~ː�d�����ϕ���  �  Y�=5e=�=	�=�`=o=̪=�M=T� =�� =75 =ұ�<���<DK�<���<���<+S�<���<�<U|�<:��<gG�<��<��<Di�<m��<;�< n�<���<W�<�]�<$��<B��<�H�<��<���<h8�<?��<c��<+�<�z�<��<��< ]�<��<j��<C�<�N�<�}�<��<���<���<��<^/�<M�<j�<m��<���<��<��<x��<���<r��<���<@��<X��<!��<�Q�<�	�<ٳ�<�P�<��<Je�<���<AM�<b��<[�<�a�<5��<��<�-�<?c�<ؑ�<<��<Yٸ<��<��<��<��<$�<���<�<BӨ<뺦<���<n��<q�<\�<WJ�<�;�<�0�<�'�<� �<O�<l�<�<* �<"�<���<w˅<��<���<m�~<�z<�uv<=5r<��m<}�i<�ye<�?a<�]<��X<5�T<�sP<~EL<	H<Y�C<��?<r~;<9C7<)3<��.<�v*<H-&<��!<��<�`<{*<?�<N�<�<;�<�� <���;��;�b�;*��;�'�;k��;��;���;O�;*��;�G�;���;�͟; ��;ɑ;���;�X�;}�{;�%o;�b;
W;E�K;Yc@;��5;�+;u� ;��;�K;��;C�:�C�:e��:��:+�:�=�:$�:fJ�:R�h:U�M:�4:bs:�M:���9��9QS�9B�<9�A�8�$�7|w��j�w�g�庞���ɹ����5��&8%�vh:��`O��#d�ŭx�)���񗐺j��������������º�̺�2׺?��2�����Z����>��XL�K���h�'�"�_(�<--��&2�: 7�Z�;�Wn@�5E�F�I��tN�>S�/ X��]��5b�8fg�s�l���q�\w�ȼ|�<������qe��������AH������Uv��U�������  �  ��=d=o=?�=fa=�=۬=�P=�� =m� =�9 =���<��<�U�<s��<K�<c]�<+��<��<��<���<�L�<���<L�<�j�<���<�<�k�<���<
�<uW�<w��<���<�?�<Q��< ��<�.�<[��<C��<$�<u�<���<��<C[�<���<6��<Z�<R�<R��<���<���<���<��<G9�<�W�<�t�<2��<(��<���<*��<���<���<5��<���<{��<M��<Ì�<RQ�<��<���<L�<���<�]�<	��<�C�<\��<	�<~W�<P��<���<i%�< \�<���<���<9ָ<.�<L�<��<�<�
�<l��<��<vڨ<5æ<ɪ�<w��<�{�<�f�<U�<IF�<Z:�<�0�<�(�</!�<�<r�<^�<�<R�<�ʅ<#��<u��<��~<�z<Lgv<�$r<��m<�i<�ee<2,a<�\<{�X<��T<�fP<5;L<�H<��C<Ͳ?<�~;<XF7<�3<��.<s�*<�:&<_�!<~�<Wt<�?<2<��<�<k�<i� <���;�2�;�}�;���;I9�;٣�;P�;��;��;蜵;:�;N�;���;᝘;_��;�؊; 3�;s{;	�n;��b;��V;�SK;�6@;Pr5;|�*;�� ;��;�S;1�;P{�:̎�:��:� �:��:_Ѡ:ˏ�:�:�i:GZO:+�5:��:�u:�9灴9�щ9�L?9���8��7�0u����qh��u����ʹ�;��~���8&��;���P��\e�y�y�����!��*��,���ܮ��Ÿ�A�ºf�̺92׺���%h�9P��$2�����j�a�ߙ�A�_x"��'�K�,���1��6�x;�/@�:�D�ӒI��RN��%S��X��]��:b��vg�O�l�(%r�Čw��|�n/��-���4���?2���ҋ��l��&������6$��D����  �  (�=�b=�=\�=\b=�	=r�=T=�� =`� =:? =���<>�<�c�<y��<�<�j�<]��<�*�<p��<���<S�<���<��<3l�<s��<K�<h�<y��<�<�N�<L��<K��<;3�<j��</��<,"�<|t�<q��<��<Wm�<���<P�<�X�<˟�<���<��<V�<��<��<���< �<|%�<F�<e�<���<��<���<���<���<���<T��<t��<���<h��<���<U��<(P�<��<��<�E�<���<6T�<���<�7�<��<g��<�I�</��<���<_�<�R�<��<���<�Ѹ<��<f�<Y�<��<��<J�<r��<~�<�ͦ<���<v��<,��<�t�<�b�<�S�<G�<B<�<�2�<�)�<Q �<�<J�<d��<��<�Ʌ<G��<ߏ�<�~<ϙz<�Sv<@r<`�m<
�i<�Ke<a<Q�\<��X<�T<�UP<Q-L<NH<��C<|�?<;<�I7<�3<��.<�*<WK&<_"<?�<��<�Z<�1<�<�	<��<�<�%�;[�;d��;���;�N�;+��;��;��;�
�;���;2'�;IѦ;~��;Gw�;�|�;���;K�;5{;czn;Ib;qyV;|K;��?;�D5;�*;F� ;��;`\;O;^��:!��:V��:���:�W�:��:�^�:�̓:ʻk:}Q:��7:�U:�:���9�Ķ9���9�EB9p�8G�7�:s���6�i��{��zM̹0!�����F�'�|�<��#R��f�%�{��߇�Tڑ�����l����O������ ú�ͺk7׺ݜ�.7캄���� �N����Ʊ�V9�����
"��H'�Eh,��g1�9M6�6;�s�?��D��ZI��'N��S�� X�f]��Db�_�g���l��Xr�D�w�5D}��[��m��M���f�����k����.��<���E���Ϙ��  �  �=z`=�=H�=;c=�=B�=�W=�� =�� =�E =+��<v#�<�s�<���<��<�y�<@��<07�<@��<���<Z�<���<��<�m�<���<��<�c�<��<���<fD�<7��<���<�$�<Ar�<���<@�<of�<���<��<�c�<��<��<@U�<V��<w��<2!�<fZ�<F��<��<���<��<�2�<�T�<~t�<���<��<%��< ��<��<� �<L�<�<���<���<̾�<���<nN�<5�<��<�=�<���<wH�<i��<�(�<u��<J��<�9�<���<#��<R�<3G�<�z�< ��<X̸<�<���<��<�<�<��<���<��<�٦< Ĥ<)��<ۘ�<�<�r�</c�<mU�<mI�<|>�<�3�<*(�<�<f�<���<)�<ȅ<���<��<��~<*�z<�<v<��q<��m<�ji<�,e<y�`<�\<��X<�gT<AP<�L<l�G<��C<��?<>~;<�L7<�3<�.<�*<=^&<"<\�<��<z<QR<�4<M"	<<�<|Z�;��;&��;��;�f�;���;�%�;i��;P�;x��;��;�;n�;[I�;�H�;�q�;�ƃ;��z;=n;��a;lV;��J;s�?;�5;\�*;6� ;.�;c;�;�	�:V�:[�:.T�:'�:~e�:�I�:kȄ:[�m:;"S:��9:�,!:�	:P��9�U�9�ˍ9˄E9���8�]�7��q�8|�i;k��ˡ��ιyj��B�� )�C�>���S���h��k}�Xʈ�2����~��=1���گ�����Mú�1ͺ�C׺G��N�۶���� ��E�����N�a���6�#�!���&�#�+�$�0���5���:�2�?�:ND��I��M���R��W��]�-Tb�1�g�m���r��x��}�����I��[�������&B���֎��c��MꓻQm����  �  ��=^=A=�=�c=7=�=�[=[=�� =`L ='��<�3�<���<���<�/�<���<���<1D�<f��<��<'a�<н�<��<dn�<���<��<6^�<o��<��<�8�<��<���<��<�a�<��<��<�V�<���<$�<{Y�<���<��<Q�<4��<a��<1#�<�^�<`��<`��<��<��<�@�<�c�<ʄ�<y��<ڿ�<y��<~��<�<��<��<��<���<���<���<?��<�K�<���<\��<�4�<��<�;�<���<��<mz�<���<N(�<�u�<B��<���<�:�<�o�<���<�Ÿ<��<���<��<*�<`�<��<Y�<G��<F�<^Ҥ<���<[��<ו�<҃�<os�<�d�<2W�<jJ�<�=�<80�<!�<I�<X��<��<�Ņ<��<b��<�~<[pz<*#v<
�q<��m<�Ii<�
e<�`<՟\<�sX<
MT<*P<�	L<��G<��C<��?<C|;<;O7<I3<��.<�*<�q&<_6"<��<"�<��<�t<�W<�D	<<<�=<I��;���;��;F1�;�}�;���;�,�;{��;&��;
o�;j��;���;fB�;��;�;4�;ކ�;cz;��m;�ea;7�U;_WJ;�d?;g�4;h�*;C� ;9�;?e;J*;^P�:[��:Ҟ�:��:�ܲ:(H�:�B�:�Ѕ:t�o:xBU:��;:D #:�h:���9��9(�9��H9���8�h�7kq��m��1m�(O��Y$й���
��L�*���@��V�x�j� ��ˉ�8����V�����v�������ú�iͺ1[׺������>i��� ����Js�r��DW����!�@&�)a+��k0��a5��G:�3%?���C� �H�X�M�z�R���W��]��hb���g�NQm��r�Xsx��~��Ɂ�6����<���扻������띑���噖�K���  �  ܪ=_[=�
=M�=Sd=�={�= _=�=a� =�R =���<jC�<��<S��<@�<$��<8��<�P�<4��<��<�g�<L��<&�<�n�<���<��<eX�<|��<	��<�,�<+s�<���<p�<�P�<��<d��<DG�<5��<s��<�N�<ץ�<���<WL�<���<���<�$�<b�<
��<2��<���<�&�<7N�<�r�<ǔ�<��<r��<v��<���<��<��<_�<s�<U�<���<���<s��<I�<���<<��<�+�<���<A.�<���<D�<i�<���<��<�d�<��<(�<�-�<�d�<���</��<�<*��<P�<��<�<��<^�<t�<l�<:�<͢<���<���<_��<j��<�s�<�d�<V�<gG�<�7�<u&�<��<���<�<�<��<G|�<}�~<�Yz<�v<X�q<�mm<�'i<�d<�`<\<UUX<�1T<}P<��K<�G<8�C<W�?<Qy;<�P7<�"3<��.<M�*<-�&<$M"<<��<b�<��<Ez<�f	<�\<o[<���;���;��;�N�;ܒ�;���;"1�;Ê�;��;�Z�;k׭;8i�;��;W�;�Ր;���;�E�;Y�y;i	m;%�`;�;U;��I;�?;�4;V*;�m ;p�;�c;T9;ю�:��:@ �:��:ޝ�:O$�:�5�:�ӆ:�q:�\W:��=:]	%:g#:P��9;��9C��9��K9f��8b��7	�q����lpo�}��Lҹ����W�٤,�:�B�HX�9m��΀��Њ�����K5��ɮ�����ㇺ��ĺ��ͺ�y׺�}���%���^ � �������1���<��� ��%���*��/���4� �9�o�>���C��H�šM�Q�R���W�� ]�Z�b�d�g��m��(s�b�x��o~����Ȅ�����*��/ǌ�RV���ّ�US���ǖ��:���  �  0�=�X=�=}�=ud=�=��=<b=
=u� =�X =�  =�Q�<5��<���< O�<\��<6�<Y\�<��<>�<�m�<��<��<�n�<��<�	�<sR�<���<T��<v!�<f�<V��<��<�@�<���<���<o8�<���<)��<D�<#��<���<uG�<���<���<�%�<�d�<��<	��<��<i1�<{Z�<���<h��</��<���<��<<�<��<d#�<%$�<=�<"
�<���<���<-��<�E�<a��<��<y"�<���<s!�<i��<���<�X�<���<��<5T�<���<�<&!�<4Z�<Ռ�<K��</ܶ<<��<G�<��<�<��<u�<��<i��<��<�ڢ<TȠ<ӵ�<���<���<��<�p�<�`�<�O�<x>�<+�<P�<[��<�߇<���<ꛃ<<u�<l�~<Dz<��u<E�q<nOm<�i<u�d<~�`<9`\<�8X<�T<��O<��K<��G<��C<��?<�u;<�P7<'3<��.<��*<��&<�a"<.0<<��<��<��<��	<z<�v<N��;D�;�6�;i�;���;���;23�;V��;�߼;�E�;��;�D�;�;R��;���;4��;��;�y;i�l;�y`;��T;h�I; �>;�G4;#*;�I ;,�;E^;�B;���:�m�:���:7.�:�L�:��:��:��:t�s:FHY:��?:+�&:��:���9���9ü�9�FN97��8�7N�s����2�q�����PjԹ�k��|U.��kD�]Z��o��ρ��ȋ�����F	���i��6������hiĺ�ͺ��׺G�������2 ��}���
�*������# �?%��c*��w/��4�~9�rv>��pC��pH�e~M��R� �W�:,]��b��%h�.�m��qs��$y���~�g<��?������k�����������z�������_���  �  ѣ=V==��=cd=�=9�=�d=d=�� =�] =' =^�<��<��<�[�<a��<:�<�e�<��<��<2r�<���<�<n�<���<��<�L�<���<���<N�<�Z�<���<���<�2�<���<���<Q+�<���<f��<�:�<`��<���<�B�<���<���<&�<g�<���<���<��<8:�<�d�<��<ͯ�<��<q��<��<��<O%�<7,�<j+�<�!�<��<���<���<���<�B�<���<���<U�<ܝ�<:�<��<��<BJ�<H��<��<�E�<B��<�տ<$�<�P�<턺<��<�׶<?��<�<>�<@ �<� �<?�<�<��<w��<��<�Ԡ<�<a��<P��<���<�z�<?i�<W�<�C�<�.�<:�<���<^އ<���<%��<�n�<W�~<�0z<t�u<��q<�4m<��h<�d<hs`<E\<3X<� T<s�O<��K<żG<�C<H�?<�q;<P7<�)3<F�.<��*<-�&<�r"<PD<�<��<�<��<�	<�<��<��;�2�;pR�;�}�;���;���;�3�;�~�;�Ҽ;�1�;ᠭ;�$�;�Þ;���;	n�;6��;"҂;S�x;{%l;+`;�uT;�DI;z>;�4;G�);#( ;ɟ;wV;>H;`��:p��:]��:ѥ�:�ܴ:Ŕ�:)ϖ:)��:�u:��Z:7,A:B?(:�:v��9_��9�.�9JP9<�8��7�u�RU���s�_���Oֹ�=��-�V�/�PF�ʿ[���p����w����N��������E���{����ĺ-κa�׺	��(������  ��L���
�"���(�el������$�x�)��/�%4��-9��2>�29C�GH��bM�$�R���W�d9]�a�b�Mh���m�y�s��qy�-�om��^9���������P>��lȏ��C�����\��ۀ���  �  "�=
T=�=õ=5d=�=Z�=�f=�=�� =�a =_
 =8g�<ͺ�<q�<ge�<b��<{�<m�<���<N�<|u�<���<��<�m�<й�<��<�H�<��<���<U�<�Q�<ڕ�<#��<(�<w�<W��<.!�<&{�<���<r3�<8��<���<D?�<C��<^��<&�<Zh�<h��<���<T�<�@�<�l�<���<"��<���<'��<��<o �<&-�<�2�<�0�<�%�<{�<���<���<d��<@�<���<c��<��<)��<n�<#{�<���<2?�<���<���<�:�<ͅ�<7̿<��<II�<�~�<��<�Ӷ<��<�	�<E�<�!�<�#�< �<��<f�<w��<��<mޠ<r̞<&��<���<��<���<�o�<_\�<�G�<R1�<e�<}��<݇<鹅<N��<�i�<�{~<�!z<�u<^qq<�m<�h<��d<�]`<0\<wX<��S<��O<�K<��G<h�C<9�?<�m;<O7<W+3<�/<��*<C�&<B"<�S<5*<�<�<��<�	<�<�<]>�;oL�;g�;Ì�;X��;���;3�;y�;ȼ;k"�;��;�;[��;ib�;FH�;%^�;���;�Vx;��k;��_;r-T;�I;fA>;��3;'�);� ;$�;�N;J;���:j��:�0�:d��:aI�:�:[�:�!�:��v:�#\:�\B:�X):�:1��9U�9�>�9L�Q9���8U�7��w��z���u�=B����׹�%�*8���0�>NG�]��9r��[���H���햺�S��P���ﴲ��׻�BźMaκ��׺ԚẀ��֤������:(��d
�X��0���$��Z�M�$�A�)�y�.���3���8�>�=��C�%)H�MOM���R���W� E]��b�~lh�m"n���s���y�Fr�����]b��R!���Ί�i����Cj��"֔�W:������  �  n�=�R=�=0�=d=A=�=�g=b=�� =�c = =m�<���<��<gk�<��<��<�q�<���<!�<�w�<��<�<m�<���<� �<�E�<p��<���<O
�<�K�<���<r��<&!�<(p�<��<��<&u�<���<�.�<G��<���<�<�<���<r��< &�<!i�<��<	��<��<�D�<|q�<-��<��<���<1��<��<�%�<�1�<�6�<4�<*(�<�<���<���<_��<=>�<���<��<��<J��<��<�t�<���<8�<���<i��<�3�<2�<ƿ<�<�D�<�z�<ǩ�<SѶ<�<		�<R�<�"�<�%�<#�<"�<��<i�<��<Z�<�Ҟ<0��<s��<���<W��<�s�<�_�<J�<�2�< �<]��<܇<��<���<Rf�<js~<
z<�u<eq<�m<6�h<�d<�O`<�"\<��W<?�S<��O<_�K<��G<��C<�?<�k;<XN7<Z,3<g/<)�*<B�&<�"<�\<5<�<v�<r�<��	<Ʊ<ש<0Q�;/\�;ys�;��;S��;���;@2�;�t�;���;��;�~�;���;H��;WL�;S0�;XD�;͍�;e!x;��k;k�_;�S;a�H;�>;ʿ3;�);��;�;�H;�J;�:��:|Y�:�4�:���:mb�:���:뀉:V�w:��\:�C:]*:��:4��9��9���9v�R97��8ª�7Qy�*A�z�v�
����عĸ����!�1��H�_�]��s��ʃ������Q��ܰ���᩺�������:ź�κ�׺���ǃ�P���������`H
����ž�����*�jX$��})�֜.�ǵ3�$�8���=�M�B��H�rCM�ڃR�6�W��M]��b��h�=n��t�&�y�X�����T|���<���ꊻ�������ł���씻�M��⫙��  �  ՞=5R=j=�=�c=M=7�=�g=�=Y� =�d =� =�n�<���<��<`m�<
��<Y�<s�<���<"�<&x�<R��<�<�l�<��< �<�D�<'��<���<��<�I�<���<-��<��<�m�<"��<��<s�<���<&-�<ԉ�<���<�;�< ��< ��<�%�<Li�<���<���<��<bF�<s�<��<���<���<9��<��<�'�<�3�<i8�<A5�<)�<��<���<���<���<�=�<.��<׀�<F�<���<��<�r�<���<�5�<<��< ��<�1�<}�<�ÿ<=�<�B�<<y�<���<�ж<��<��<H�<�"�<&�<�#�<U�<�<�<���<M�<�Ԟ<1<f��<[��<䈖<)u�<�`�<�J�<M3�<C�<I��<�ۇ<���<܏�<+e�<Vp~<�z<V�u<�`q<em<m�h<_�d<�J`<"\<��W<_�S<�O<(�K<�G<��C<�?<�j;<�M7<�,3</<��*<Z�&<Ɖ"<�_<�8<�<��<��<��	<Ե<|�<�W�;�a�;�w�;���;���;��;�1�;�s�;���;I�;z�;���;ŋ�;�D�;p(�;�;�;ل�;�x;S�k;��_;R�S;~�H;>;��3;��);�;�~;vF;K;{�:� �:�g�:�G�:ң�:|�:�җ:���:��w:�)]:7ZC:AH*:u�:� �9F6�9b�9K�R9v��8!��7��y��z��Ew��O��H!ٹ����p�1�E]H�6^�`s�Lٍ��r��JР���������'��QKźi�κ�غ
����ŏ�������
�[>
��w�"��I��2��G$��m)�O�.�3�3��8���=���B��H�v@M���R��W�CP]��b���h�lFn�t���y�<��a���I���MF��s��������������T��#����  �  n�=�R=�=0�=d=A=�=�g=b=�� =�c = =m�<���<��<gk�<��<��<�q�<���<!�<�w�<��<�<m�<���<� �<�E�<p��<���<O
�<�K�<���<r��<&!�<(p�<��<��<&u�<���<�.�<G��<���<�<�<���<r��< &�<!i�<��<	��<��<�D�<|q�<-��<��<���<1��<��<�%�<�1�<�6�<4�<*(�<�<���<���<_��<=>�<���<��<��<J��<��<�t�<���<8�<���<i��<�3�<2�<ƿ<�<�D�<�z�<ǩ�<TѶ<�<
	�<R�<�"�<�%�<#�<"�<��<i�<��<Z�<�Ҟ<0��<s��<���<W��<�s�<�_�<J�<�2�<�<]��<܇<��<���<Rf�<js~<
z<�u<eq<�m<6�h<�d<�O`<�"\<��W<?�S<��O<_�K<��G<��C<�?<�k;<XN7<Z,3<g/<)�*<B�&<�"<�\<5<�<v�<r�<��	<Ʊ<ש<0Q�;.\�;ys�;��;R��;���;?2�;�t�;���;��;�~�;���;G��;VL�;S0�;WD�;̍�;d!x;��k;j�_;�S;a�H;�>;ʿ3;�);��;�;�H;�J;�:��:|Y�:�4�:���:mb�:���:뀉:V�w:��\:�C:]*:��:4��9��9���9v�R97��8ª�7Qy�*A�z�v�
����عĸ����!�1��H�_�]��s��ʃ������Q��ܰ���᩺�������:ź�κ�׺���ǃ�P���������`H
����ž�����*�jX$��})�֜.�ǵ3�$�8���=�M�B��H�rCM�ڃR�6�W��M]��b��h�=n��t�&�y�X�����T|���<���ꊻ�������ł���씻�M��⫙��  �  "�=
T=�=õ=5d=�=Z�=�f=�=�� =�a =_
 =8g�<ͺ�<q�<ge�<b��<{�<m�<���<N�<|u�<���<��<�m�<й�<��<�H�<��<���<U�<�Q�<ڕ�<#��<(�<w�<W��<.!�<&{�<���<r3�<8��<���<D?�<C��<^��<&�<Zh�<h��<���<T�<�@�<�l�<���<"��<���<'��<��<o �<&-�<�2�<�0�<�%�<{�<���<���<d��<@�<���<c��<��<)��<o�<#{�<���<2?�<���<���<�:�<΅�<8̿<��<II�<�~�<��<�Ӷ<��<�	�<E�<�!�<�#�< �<��<f�<w��<��<mޠ<r̞<&��<���<��<���<�o�<_\�<�G�<R1�<d�<|��<݇<鹅<M��<�i�<�{~<�!z<�u<]qq<�m<�h<��d<�]`<0\<xX<��S<��O<�K<��G<h�C<:�?<�m;< O7<X+3<�/<��*<D�&<C"<�S<5*<�<�<��<�	<�<�<\>�;nL�;g�;�;W��;���;3�;y�;ȼ;i"�;��;�;Y��;gb�;DH�;$^�;���;�Vx;��k;��_;q-T;�I;eA>;��3;'�);� ;#�;�N;J;���:i��:�0�:d��:aI�:�:[�:�!�:��v:�#\:�\B:�X):�:1��9U�9�>�9L�Q9���8U�7��w��z���u�=B����׹�%�*8���0�>NG�]��9r��[���H���햺�S��P���ﴲ��׻�BźMaκ��׺ԚẀ��֤������:(��d
�X��0���$��Z�M�$�A�)�y�.���3���8�>�=��C�%)H�MOM���R���W� E]��b�~lh�m"n���s���y�Fr�����]b��R!���Ί�i����Cj��"֔�W:������  �  ѣ=V==��=cd=�=9�=�d=d=�� =�] =' =^�<��<��<�[�<a��<:�<�e�<��<��<2r�<���<�<n�<���<��<�L�<���<���<N�<�Z�<���<���<�2�<���<���<Q+�<���<f��<�:�<`��<���<�B�<���<���<&�<g�<���<���<��<8:�<�d�<��<ͯ�<��<q��<��<��<O%�<8,�<j+�<�!�<��<���<���<���<�B�<���<���<U�<ݝ�<:�<��<��<BJ�<I��<��<�E�<B��<�տ<%�<�P�<턺<��<�׶<@��<�<>�<@ �<� �<?�<�<��<w��<��<�Ԡ<�<a��<O��<���<�z�<>i�<W�<�C�<�.�<9�<���<^އ<���<%��<�n�<V�~<�0z<s�u<��q<�4m<��h<�d<hs`<E\<3X<� T<t�O<��K<ƼG<�C<I�?<�q;<P7<�)3<H�.<��*<.�&<�r"<QD<�<��<�<��<�	<�<��<��;�2�;nR�;�}�;���;���;�3�;�~�;�Ҽ;�1�;ޠ�;�$�;�Þ;���;n�;4��;!҂;P�x;y%l;)`;�uT;�DI;z>;�4;F�);"( ;ȟ;vV;=H;_��:o��:]��:Х�:�ܴ:Ŕ�:)ϖ:)��:�u:��Z:7,A:B?(:�:v��9_��9�.�9JP9<�8��7�u�RU���s�_���Oֹ�=��-�V�/�PF�ʿ[���p����w����N��������E���{����ĺ-κa�׺	��(������  ��L���
�"���(�el������$�x�)��/�%4��-9��2>�29C�GH��bM�$�R���W�d9]�a�b�Mh���m�y�s��qy�-�om��^9���������P>��lȏ��C�����\��ۀ���  �  0�=�X=�=}�=ud=�=��=<b=
=u� =�X =�  =�Q�<5��<���< O�<\��<6�<Y\�<��<>�<�m�<��<��<�n�<��<�	�<sR�<���<T��<v!�<f�<V��<��<�@�<���<���<o8�<���<)��<D�<#��<���<uG�<���<���<�%�<�d�<��<	��<��<i1�<{Z�<���<h��</��<���<��<<�<��<d#�<%$�<=�<"
�<���<���<-��<�E�<a��<��<y"�<���<s!�<i��<���<�X�<���<��<6T�<���<�<&!�<4Z�<֌�<L��<0ܶ<=��<H�<��<�<��<v�<��<j��<��<�ڢ<TȠ<ӵ�<���<���<��<�p�<�`�<�O�<w>�<+�<P�<Z��<�߇<���<ꛃ<<u�<k�~<Dz<��u<D�q<mOm<�i<u�d<~�`<9`\<�8X<�T<��O<��K<��G<��C<��?<�u;<�P7<'3<��.<��*<��&<�a"<.0<<��<��<��<��	<z<�v<L��;B�;�6�;i�;���;���;/3�;S��;�߼;�E�;��;�D�;�;O��;���;1��;��;�y;f�l;�y`;�T;f�I;�>;�G4;#*;�I ;+�;D^;�B;���:�m�:���:7.�:�L�:��:��:��:t�s:FHY:��?:+�&:��:���9���9ü�9�FN97��8�7N�s����2�q�����PjԹ�k��|U.��kD�]Z��o��ρ��ȋ�����F	���i��6������hiĺ�ͺ��׺G�������2 ��}���
�*������# �?%��c*��w/��4�~9�rv>��pC��pH�e~M��R� �W�:,]��b��%h�.�m��qs��$y���~�g<��?������k�����������z�������_���  �  ܪ=_[=�
=M�=Sd=�={�= _=�=a� =�R =���<jC�<��<S��<@�<$��<8��<�P�<4��<��<�g�<L��<&�<�n�<���<��<eX�<|��<	��<�,�<+s�<���<p�<�P�<��<d��<DG�<5��<s��<�N�<ץ�<���<WL�<���<���<�$�<b�<
��<2��<���<�&�<7N�<�r�<ǔ�<��<r��<v��<���<��<��<_�<s�<U�<���<���<s��<I�<���<=��<�+�<���<B.�<���<D�<i�<���<��<�d�<��<(�<�-�<�d�<���<0��<�<+��<Q�<��<�<��<_�<u�<l�<;�<͢<���<���<_��<j��<�s�<�d�<V�<fG�<�7�<t&�<��<���<�<�<��<G|�<{�~<�Yz<�v<W�q<�mm<�'i<�d<�`<\<UUX<�1T<~P<��K< �G<:�C<X�?<Sy;<�P7<�"3<��.<N�*</�&<%M"<<��<c�<��<Ez<�f	<\<n[<���;���;��;�N�;ْ�;���;1�;���;��;�Z�;h׭;5i�;��;T�;�Ր;���;�E�;U�y;f	m;"�`;�;U;��I;�?;�4;V*;�m ;o�;�c;T9;Ў�:��:? �:��:ޝ�:O$�:�5�:�ӆ:�q:�\W:��=:]	%:g#:P��9;��9C��9��K9f��8b��7	�q����lpo�}��Lҹ����W�٤,�:�B�HX�9m��΀��Њ�����K5��ɮ�����ㇺ��ĺ��ͺ�y׺�}���%���^ � �������1���<��� ��%���*��/���4� �9�o�>���C��H�šM�Q�R���W�� ]�Z�b�d�g��m��(s�b�x��o~����Ȅ�����*��/ǌ�RV���ّ�US���ǖ��:���  �  ��=^=A=�=�c=7=�=�[=[=�� =`L ='��<�3�<���<���<�/�<���<���<1D�<f��<��<'a�<н�<��<dn�<���<��<6^�<o��<��<�8�<��<���<��<�a�<��<��<�V�<���<$�<{Y�<���<��<Q�<4��<a��<1#�<�^�<`��<`��<��<��<�@�<�c�<ʄ�<y��<ڿ�<y��<~��<�<��<��<��<���<���<���<?��<�K�<���<\��<�4�<��<�;�<���<��<nz�<���<N(�<�u�<C��<���<�:�<�o�<���<�Ÿ<��<���<��<+�<a�< �<Y�<H��<G�<^Ҥ<���<\��<ו�<҃�<os�<�d�<1W�<iJ�<�=�<70�<!�<H�<X��<��<�Ņ<��<a��<�~<Zpz<)#v<	�q<��m<�Ii<�
e<�`<֟\<�sX<MT<*P<�	L<��G<��C<��?<E|;<=O7<K3<��.<�*<�q&<`6"<��<#�<��<�t<�W<�D	<<<�=<G��;���;��;C1�;�}�;���;|,�;w��;"��;o�;g��;���;cB�;��;��;4�;܆�;_z;��m;�ea;4�U;\WJ;�d?;e�4;f�*;A� ;9�;>e;I*;]P�:[��:Ҟ�:��:�ܲ:'H�:�B�:�Ѕ:t�o:xBU:��;:C #:�h:���9��9(�9��H9���8�h�7kq��m��1m�(O��Y$й���
��L�*���@��V�x�j� ��ˉ�8����V�����v�������ú�iͺ1[׺������>i��� ����Js�r��DW����!�@&�)a+��k0��a5��G:�3%?���C� �H�X�M�z�R���W��]��hb���g�NQm��r�Xsx��~��Ɂ�6����<���扻������띑���噖�K���  �  �=z`=�=H�=;c=�=B�=�W=�� =�� =�E =+��<v#�<�s�<���<��<�y�<@��<07�<@��<���<Z�<���<��<�m�<���<��<�c�<��<���<fD�<7��<���<�$�<Ar�<���<@�<of�<���<��<�c�<��<��<@U�<V��<w��<2!�<fZ�<F��<��<���<��<�2�<�T�<~t�<���<��<%��< ��<��<� �<L�<��<���<���<̾�<���<nN�<5�<��<�=�<���<wH�<j��<�(�<u��<J��<�9�<���<$��<R�<4G�<�z�<!��<Y̸<�<���<��<�<�<��<���<��<�٦<!Ĥ<)��<ۘ�<�<�r�</c�<mU�<lI�<{>�<�3�<)(�<�<e�<���<)�<ȅ<���<��<��~<)�z<�<v<��q<��m<�ji<�,e<y�`<�\<��X<�gT<AP<�L<n�G<��C<��?<?~;<�L7<�3<�.<�*<>^&<"<]�<��<z<QR<�4<M"	<<�<{Z�;��;$��;��;�f�;���;�%�;f��;L�;u��;��;�;n�;XI�;�H�;�q�;�ƃ;��z;:n;��a;jV;�J;q�?;�5;[�*;5� ;-�;c;�;�	�:V�:Z�:.T�:'�:}e�:�I�:kȄ:[�m:;"S:��9:�,!:�	:P��9�U�9�ˍ9˄E9���8�]�7��q�8|�i;k��ˡ��ιyj��B�� )�C�>���S���h��k}�Xʈ�2����~��=1���گ�����Mú�1ͺ�C׺G��N�۶���� ��E�����N�a���6�#�!���&�#�+�$�0���5���:�2�?�:ND��I��M���R��W��]�-Tb�1�g�m���r��x��}�����I��[�������&B���֎��c��MꓻQm����  �  (�=�b=�=\�=\b=�	=r�=T=�� =`� =:? =���<>�<�c�<y��<�<�j�<]��<�*�<p��<���<S�<���<��<3l�<s��<K�<h�<y��<�<�N�<L��<K��<;3�<j��</��<,"�<|t�<q��<��<Wm�<���<P�<�X�<˟�<���<��<V�<��<��<���< �<|%�<F�<e�<���<��<���<���<���<���<T��<t��<���<h��<���<U��<(P�<��<��<�E�<���<7T�<���<�7�<��<g��<�I�</��<���<`�<�R�<��<���<�Ѹ<��<g�<Z�<��<��<K�<s��<�<�ͦ<���<v��<,��<�t�<�b�<�S�<G�<B<�<�2�<�)�<P �<�<I�<d��<��<�Ʌ<G��<ޏ�<�~<Ιz<�Sv<?r<`�m<
�i<�Ke<a<R�\<��X<�T<�UP<R-L<OH<��C<}�?<;<�I7<�3<��.<�*<XK&<`"<@�<��<�Z<�1<�<�	<��<�<�%�;[�;b��;���;�N�;(��;��;��;�
�;�;/'�;FѦ;|��;Ew�;�|�;���;I�;2{;`zn;Ib;oyV;zK;��?;�D5;�*;E� ;��;_\;O;]��: ��:V��:���:�W�:��:�^�:�̓:ʻk:}Q:��7:�U:�:���9�Ķ9���9�EB9p�8G�7�:s���6�i��{��zM̹0!�����F�'�|�<��#R��f�%�{��߇�Tڑ�����l����O������ ú�ͺk7׺ݜ�.7캄���� �N����Ʊ�V9�����
"��H'�Eh,��g1�9M6�6;�s�?��D��ZI��'N��S�� X�f]��Db�_�g���l��Xr�D�w�5D}��[��m��M���f�����k����.��<���E���Ϙ��  �  ��=d=o=?�=fa=�=۬=�P=�� =m� =�9 =���<��<�U�<s��<K�<c]�<+��<��<��<���<�L�<���<L�<�j�<���<�<�k�<���<
�<uW�<w��<���<�?�<Q��< ��<�.�<[��<C��<$�<u�<���<��<C[�<���<6��<Z�<R�<R��<���<���<���<��<G9�<�W�<�t�<2��<(��<���<*��<���<���<5��<���<{��<M��<Č�<SQ�<��<���<L�<���<�]�<	��<�C�<\��<	�<W�<P��<���<i%�< \�<���<���<:ָ</�<M�<��<�<�
�<m��<��<vڨ<6æ<ɪ�<w��<�{�<�f�<U�<IF�<Z:�<�0�<�(�<.!�<�<r�<]�<�<Q�<�ʅ<#��<t��<��~<�z<Lgv<�$r<��m<�i<�ee<2,a<�\<{�X<��T<�fP<6;L<�H<��C<β?<�~;<YF7<�3<��.<s�*<�:&<`�!<�<Xt<�?<2<��<�<k�<i� <���;�2�;�}�;���;G9�;ף�;N�;��;��;朵;:�;L�;���;ޝ�;]��;�؊;�2�;s{;�n;��b;��V;~SK;�6@;Nr5;{�*;�� ;��;�S;1�;O{�:ˎ�:��:� �:��:_Ѡ:ˏ�:�:�i:GZO:+�5:��:�u:�9灴9�щ9�L?9���8��7�0u����qh��u����ʹ�;��~���8&��;���P��\e�y�y�����!��*��,���ܮ��Ÿ�A�ºf�̺92׺���%h�9P��$2�����j�a�ޙ�A�_x"��'�K�,���1��6�x;�/@�:�D�ӒI��RN��%S��X��]��:b��vg�O�l�(%r�Čw��|�n/��-���4���?2���ҋ��l��&������6$��D����  �  Y�=5e=�=	�=�`=o=̪=�M=T� =�� =75 =ұ�<���<DK�<���<���<+S�<���<�<U|�<:��<gG�<��<��<Di�<m��<;�< n�<���<W�<�]�<$��<B��<�H�<��<���<h8�<?��<c��<+�<�z�<��<��< ]�<��<j��<C�<�N�<�}�<��<���<���<��<^/�<M�<j�<m��<���<��<��<x��<���<r��<���<@��<X��<!��<�Q�<�	�<ٳ�<�P�<��<Je�<���<AM�<b��<\�<�a�<5��<��<�-�<?c�<ّ�<=��<Yٸ<��<��<��< �<$�<���<�<CӨ<캦<���<n��<q�<\�<WJ�<�;�<�0�<�'�<� �<N�<l�<�<* �<!�<���<v˅<��<���<l�~<�z<�uv<<5r<��m<}�i<�ye<�?a<�]<��X<5�T<�sP<EL<
H<Z�C<��?<s~;<9C7<)3<��.<�v*<I-&<��!<��<�`<{*<?�<N�<�<;�<�� <���;��;�b�;)��;�'�;j��;��;���;N�;(��;�G�;���;�͟;���;�ȑ;���;�X�;{�{;�%o; �b;	W;D�K;Xc@;��5;�+;t� ;��;�K;��;C�:�C�:e��:��:+�:�=�:#�:fJ�:R�h:U�M:�4:bs:�M:���9��9QS�9B�<9�A�8�$�7|w��j�w�g�庞���ɹ����5��&8%�vh:��`O��#d�ŭx�)���񗐺j��������������º�̺�2׺?��2�����Z����>��XL�K���h�'�"�_(�<--��&2�: 7�Z�;�Wn@�5E�F�I��tN�>S�/ X��]��5b�8fg�s�l���q�\w�ȼ|�<������qe��������AH������Uv��U�������  �  n�=�e==ܸ=�_=o=e�=0L=3� =� =d2 =���<���<`D�<���<���<�L�<���<��<�w�<&��<D�<=��<�	�<<h�<C��<��<�o�<���<w�<�a�<ݰ�<���<�N�<)��<��<_>�<��<f��<d/�<o~�<���<��<^�<R��<���<��<rL�<�z�<=��<t��<l��<�
�<)�<aF�<4c�<��<���<���<@��<X��<��<���<���<��<��<���<9R�<�
�<��<�S�<���<�i�<���<,S�<���<��<<h�<q��<���<�2�<�g�<c��<���<D۸<��<��<�<��<��<���<@�<�Ψ<���<���<��<@j�<,U�<oC�<55�<B*�< "�<��<��<��<�<���<���<��<�˅<E��<Ǚ�<�~<y�z<�~v<�?r<� n<��i<7�e<9La<�]<w�X<��T<�{P<�KL<�H<F�C<��?<�};<A7<G�2<�.<�o*<�$&<��!<(�<T<
<!�< �<��<ս<�� <���;T��;XQ�;˱�;8�;���;��;ى�;��;*��;�O�;
�;�ܟ;�̘;�ݑ;�;�o�;��{;�So;hc;�1W;<�K;�}@;��5;�#+;�� ;��;pE;r�;��:��:�|�:�d�:�ׯ:nߟ:���:D݁:+�g:QM:<�3:��:�:���9���9}_�9�g;9c��8`�7ϣx�hZ��2g��G��oɹk��Y��$�E�9�}�N��`c���w��$���?���K��8O��LR��\_��<�º!�̺�3׺��ẳ�������s������mw�r�כ��#��G(��d-��[2��17�4�;�:�@��7E���I�ʋN��NS�f*X�� ]�j2b�F\g�ۚl�!�q�Y>w���|��������lM���򈻕���&1��~ː�d�����ϕ���  �  v�=*^=�=��=
X=:�=C�=rG=� =�� =c2 =0��<���<�H�<?��<c��<�J�<0��<��<�e�<^��<x&�<��<���<�;�<u��<p��<�:�<}��<l��<.(�<=u�<��<��<�[�<���<a��<5B�<���<[��<�$�<~m�<���<���<�5�<�p�<d��<���<��<V.�<�R�<�s�<Q��<���<���<���<���<��<��<�-�<7�<�9�<�4�<f&�<��<���<���<2}�<4�<���<�|�<I�<���<H�<���<*��<�O�<H��<���<?�<��<���<<�<��<j<�<�Y�<p�<H�<���<���<υ�<}�<~p�<fa�<�P�<@�<�/�<!�<c�<�	�<=�<7��<X��<��<��<���<l׋<eˉ<���<��<���<-��<N�~<��z<�ev<�/r<��m<P�i<v�e<>^a<�-]<��X<��T<�P<%L<PUH<X*D<��?<^�;<@�7<�f3<�./<D�*<�&<��"<�M<�<Y�<V�<��<f�	<U�<��<d��;��;�v�;?��;O�;F��;
S�;���;{��;�.�;]�;��;��;N��;ؔ;;"�;Ƒ�;�(�;4�u;Τi;s�];�OR;�$G;K<;I�1;[|';�~;�;SB
;�� ;���:KQ�:5�:1��:���:�"�:�F�:��:ֳd:q�J:Fa1:�):��::��9�B�9��z9}6#9���8x+���ø�9�DI���	��z�߹���@��0�*F�-[� "p��w��"Ɍ�v���G������õ�����~ʺ 	պ[�ߺΊ�ӄ��M �����}���V����{!�C�&���+���0���5�J�:�h�?�kyD�FHI�� N��S��W�3]�,b��_g���l�L�q��Iw���|�� ��ŭ��hX��S ������pH���萻����a&��ǘ��  �  (�=^=�=��=-X=p�=��=�G=�� =/� =3 =���<���<�J�<��<%��<mL�<���<9�<'g�<g��</'�<���<%��<(<�<���<O��<�:�<׊�<���</'�<t�<���<H�<�Y�<Ħ�<���<�@�<a��<B��<�#�<�l�<.��<r��<�5�<q�<���<y��<��<//�<�S�<Iu�<ѓ�<"��<���<��<���<U�<C!�<X/�<P8�<�:�<z5�<	'�</�<	��<ȹ�<"}�<�3�<���<�{�<H�<h��<��<u��<���<�M�<��<f��<�=�<�~�<o��<E�<�<�;�<�Y�<p�<o�<���<��<r��<�}�<�q�<�b�<_R�<�A�<�1�<�"�<7�<v�<��<���<���<��<S�<��<�׋<�ˉ<���<���<v��<��<��~<��z<�cv<-r<��m<�i<�e<�Za<�*]< �X<T�T<�P<w}L<TH<�)D<��?<��;<��7<�g3<"0/<��*<I�&<M�"<�P<�!<��<�<��<�	<��<��<A��;$�;{�;k��;�Q�;��;IT�;@��;D��;w-�;�;廩;]��;��;MӔ;��;N��;�!�;v�u;��i;��];[GR;�G;hE<;��1;�z';;�;,E
;S;���:S_�:�H�:���:��:9<�:ga�:�!�:��d: �J:9�1:�Z:?�:3�9�|�9�z9p�#9��8P�)��øK99�Tg��l7����߹˿��h���0��=F��d[�cXp�����ߌ� ��dX������ε�[����ʺպ˳ߺ?��Q{���G ����Zs���ے�*��m!�]�&�I�+���0�1�5���:��?�2pD�BI�zN� S���W��
]��,b��ag�A�l���q�bQw���|��������^��e��+���ON���퐻���;*��=ʘ��  �  J�=r]=�=��=�X='�=��=I=#� =�� =*5 =K��<x �<�O�<��<��<1Q�<5��<8�<�j�<h��<�)�<���<n��<�<�<���<���<O9�<���<��<$�<zp�<���<��<|U�<H��<w��<�<�<���<���<#!�<�j�<���<|��<�5�<q�<���<$��<��<�1�<JW�<y�<��<ô�<w��<i��<r��<-�<�%�<�3�<<�<*>�<38�<3)�<��<���<��<�|�<�2�<O��<�y�<X�<ܑ�<��<��<���<�H�<ɠ�<���<A9�<�z�<���<q�<��<W:�<�X�<�o�<��<���<ǋ�<���<ŀ�<u�<�f�<�V�<LF�<{6�<�'�<'�<U�<m�<���<_��<�<�<��<|ً<�̉< ��<���<k��<�}�<B�~<ȓz<�\v<0%r<�m<*�i<ǃe<�Qa<9"]<�X<�T<ʠP<�xL<[PH<:'D<C�?<��;<8�7<�j3<=4/<��*<��&<��"<Y<7+<�<,�<�<0�	<��<:�<��;3�; ��;��;�Z�;��;�W�;"��;O��;&)�;~�;���;���;I��;�Ô;&�;9z�;��;��u;0yi;>�];�-R;�G;�5<;O�1;4t';"};
�;�M
;o;��:��:�:�:t��:]��: ��:Aq�:�e:CYK:�*2:��:�c:��92�9|9ba$9���8:�%���øȪ9��ň�,���0��*�R���p1���F���[���p��ӂ�� ���Z��񋡺Ӹ��~쵺�0���ʺ�	պ�ߺ�q�3]���4 �/��VW�)��{o�>���F!���&���+���0�w�5�=�:���?�~VD�-I�q
N��R���W��]��0b��jg���l��
r��hw�d�|�����ă�jp��W��꽋�__������<���I6���Ә��  �  ް=�\=B=Ͱ=!Y=, =�=!K=�� =ߓ =o8 =a��<�<�W�<5��<���<�X�<-��<��<<p�<��<v-�<M��<B��<�=�<w��<���<B7�<��<���<�<�j�<6��<��< N�<��<$��<�5�<w��<���<��<
g�<��<��<#5�<�q�<��<f��<�<E6�<]\�<�<ƞ�<��<;��<`��<m�<��<,-�<M:�<B�<:C�<�<�<{,�<��<E��<h��<|�<1�<���<�u�<��<C��<��<y�<G��<5A�<��<8��<Y2�<`t�<���<��<V�<�7�<%W�<@o�<H��<m��<��<&��<*��<Yz�<�l�<~]�<�M�<N>�<�/�< #�<�<��<��<O��<��<F��<��<�ۋ<�͉<R��<�<Ɠ�<L{�<��~<`�z<�Qv<�r<1�m<F�i<�te<�Ba<]<&�X<��T<ݖP<zpL<^JH<E#D<j�?<��;<B�7<}n3<:/<�+<Z�&<C�"<Wf<�9<7<z�<��<��	<D�<��<��;�J�;#��;���;�f�;���;�\�;2��;�}�;L"�;~ذ;���;���;W��;`��;���;�]�;>�;<ju;�Ei;|y];�R;I�F;�<;ڝ1;j';�z;��;�Z
;�#;�Q�:%��:@��:hU�:Qa�:8��:.�:i�:�f:�UL:�3:�:�):�Z�9;P�9�}99�%9���8$m!��7ĸ�T:��_��ŗ��0�ṟ��ܡ��D2��G��\�M�q��F�����������ܡ���� ���S����ʺ�պ��ߺ3V��3��� �G���+����:8�/��_!��L&��x+��0�H�5�at:��S?�/D��I� �M��R�(�W�%]��5b�Zxg�f�l� )r���w���|��.��
���܍���6��Uۋ�{���������~I��+㘻�  �  �=5[=�=̰=�Y=z=��=�M=�� =�� =�< =���<��<�a�<|��<
�<b�<;��<��<Nw�<
��<62�<֍�<���<�>�<'��<���<Z4�<���<���<~�<�b�<���<���<�D�<O��<���<�,�<A{�<r��<��<Tb�<���<���<?4�<Tr�<ݫ�<g��<A�<�;�<�b�<���<j��<n��<��<���<��<�%�<�6�<�B�<�I�<�I�<�A�<�0�<��<���<���<�z�<�.�<���<�p�<X �<Ԅ�<���<�o�<u��<7�<��<z��<&)�<�k�<G��<�ݻ<��<D4�<�T�<^n�<���<A��<'��<r��<���<	��<�t�<Hf�<AW�<@H�<1:�<R-�<�!�<��<&�<��<���<���<
�<�ދ<�ω<���<ݨ�<V��<�w�<ҷ~<~z<�Bv<�r<�m<"�i<Xae<�/a<�]<��X<�T<ЉP<�eL</BH<�D<n�?<~�;<��7<�s3<�A/<+<��&<�"<Zw<wL<Y(<S<��<[�	<~�<��<Q+�;�h�;���;��;�v�; ��;�b�;���;�x�;o�;�ɰ;���;Ko�;�k�;���;�͍;9�;)π;&"u;�i;l:];��Q;2�F;D�;;�1;=Z';�u;��;.j
;N=;���:9-�:{=�:�ҽ:��:���:`Ώ:˗�:��g:H�M:J4:��:%:a�9���9��9u''9�q�8���a�ĸ�_;��4��\���G*�Q��'���]3���H�0^�ws��ك�.���6���G���T���d��w����ʺ�պ/�ߺ�2�,��������p�t�
�(v�����\�� �|�%�>'+��<0��>5�j0:�2?���C�y�H���M�%�R�x�W�]�X?b���g�s�l��Pr��w��1}�3P���������>]��W��@����8���Γ��b�������  �  ��=�Y=�=��=[Z=�=�=nP=9� =�� =]A ='��<I�<�m�<_��<��<�m�<���< #�<]�<���<t7�<ő�<���<�?�<���<���<�0�<�|�<��<��<�Y�<g��<���<<9�<݅�<���<g"�<�q�<���<w�<�\�<]��<��<3�<�r�<l��<���<��<�A�<|j�<`��<:��<8��<���<\�<d�<N1�<eA�<�L�<eR�<EQ�<�G�< 5�<��<M��<���<�y�<�+�<V��<�j�<���<�{�<���<�d�<���<+�<��<���<2�<%b�<���<xֻ<��<�/�<R�<1m�<��<⍰<��<%��<���<���<p}�<Kp�<0b�<�S�<F�<(9�<b-�<�"�<��<j�<��<t��<��<��<�Љ<���<j��<j��<s�<�~< oz<e1v<�q<m�m<�i<Je<�a<��\<{�X<��T<�yP<�XL<-8H<�D<��?<��;<��7<�x3<�I/<&+<+�&<�"<��<�a<~?<�$<Y<�	
<�
<D<*R�;���;
��;�'�;���;U��;gh�;���;�r�;L�;<��;mw�;QQ�;{I�;�c�; ��;��;��;��t;�h;�\;��Q;<�F;��;;�d1;�F';-n;`�;�x
;�X;~��:��:���:e_�:���:3E�:I��:�V�:�Zi:PO:��5:P:@:T��9�E�9C,�9w�(9�0�8\ ���Ÿ��<��8��������������,�4��=J�r�_��pt����e����ɘ��ɢ�;�������ؿ����ʺ:պ�ߺ�����l����;�δ
�j-�ߞ��XY �i�%�v�*���/���4���9���>��C���H�f�M���R�/�W�]��Kb���g�Fm��r�-�w�Fw}�dw���.��k������<.��tʎ��`��	�l���~���  �  ͩ=�W=�=i�=�Z==4�=HS=�� =� =nF =E��<#)�<z�<���<*"�<[y�<���<�,�<Ň�<���<�<�<���<��<S@�<���<W��<�,�<�v�<Ϳ�<��<�O�<S��<���<�,�<vy�<���<��<?g�<���<��<,V�<o��<���<D1�<�r�<���<���<��<�G�<3r�<���<���<���<���<��<�)�<`=�<�L�<>W�<�[�<�X�<	N�<�9�<��<���<���<�w�<.(�<��<d�<y��<&r�<��<�X�<��<��<�u�<?��<V�<iW�<��<sλ< �<+�<�N�<pk�<��<z��<���<�<f��<���<݆�<�z�<�m�<`�<�R�<�E�<Z9�<�-�<9#�<q�<��<��<'�<�<f҉<v��<y��<���<�m�<t�~<�^z<1v<��q<Ѡm<�fi<�0e<��`<��\<S�X<�T<�hP<�JL<�,H<�D<��?<>�;<��7<�}3<2R/<�$+<��&<��"<4�<�x<�W<(><@,<>#
<#<2,<�{�;Ү�;'��;�?�;~��;���;�m�;9��;�j�;���;��;�\�;o0�;�#�;,9�;7v�;5ކ;As�;Wot;QWh;��\;2FQ;�EF;��;;�?1;�/';�b;R�;C�
;ss;I4�:���:V8�:E��:18�:���:�K�:� �:��j:��P:�7:�p:Xm:o��9,�9�e�9Q�*9Y��8V��^�Ǹ�(>�Bg������\�湒�	�/ �
6��K��a�?�u��H��Xk���j���W��,6��~�� ��?˺}1պ�{ߺL�����$?�����r
�����G�������6%��d*�M�/���4�d�9���>���C���H�c�M���R�(�W�\	]��\b��g��7m�%�r�->x���}�C����]��*��˼��_����������������",���  �  ��=�U=[=�=?[=>=�=V=\� =N� =NK =+��<�4�<G��<[��<U.�<��<,��<Y6�<���<z��<B�<��<��<�@�<S��<}��<5(�<�p�<E��<���<�E�<��<���<s �<�l�<H��<N�<i\�<��<e��<tO�<N��<B��<D/�<%r�<E��<v��<�<�M�<�y�<z��<���<���<��<�<6�<LI�<�W�<Va�<~d�<``�<	T�<>�<��<���<��<Ou�<Q$�<���<�\�<���<h�<���<tL�<5��<��<�h�<��<U�<FL�<7��< ƻ<Q��<�%�<9K�<di�<���<Ӑ�<���<���<���<P��<���<F��<y�<l�<�^�<�Q�<FE�<9�<3-�<9!�<��<i�<\��<$�<vӉ<̼�<H��<"��<|h�<v�~<�Mz<P
v<^�q<"�m<�Mi<me<��`<��\<��X<ltT<�VP<�;L<� H<D<8�?<��;<��7<��3<�Y/<�/+<�'<��"<�<ێ<�o<HW<�E<o<
<F;<�B<Σ�;���;.�;�V�;���;��;%q�;.��;�a�;V�;[��;�@�;��;d��; �;.H�;%��;�B�;wt;�g;IM\;j�P;�F;�h;;�1;�';�T;
�;��
;��;h~�:\�:D��:��:Eܯ:v��:R�:u�:�|l:R:��8:��:��:t��9�t�9䏃9,9t�8̪�@Xɸ+�?�X���bR��@���@t!���7�SGM���b�f�w��	��� ��d��꣺����z��SO���;˺qIպ�yߺ��麩Q������2���2
�������J������$�~*�-#/��74�bB9�hH>�rMC��WH�lM���R���W��]�"ob���g�>cm�{�r��x�.~�E΁������B��ϐ���(��F���A���Ŗ��H���  �  >�=�S==^�=_[='=ï=}X= =-� =�O =-��<�?�<���<���<}9�<���<���<?�<a��<h��<�F�<��<���<�@�<���<���<�#�<
k�<��<Q��<�;�<^��<z��<��<a�<���<@ �<@R�<��<}��<�H�<N��<���<C-�<sq�<��<���<�!�<>S�<c��<���<���<��<p�<T*�<gA�<2T�<>b�<�j�<�l�<%g�<=Y�<�A�<��<n��<���<s�<c �<T��<,V�<���<�^�<��<�@�<���<>�<;\�<_��<���<�A�<���<���<��<� �<�G�<ag�<��<���<�<���<��<Q��<F��<���<���<w�<Fj�<)]�<.P�<CC�<Q6�<>)�<m�<��<���<M�<ԉ<���<��<8��<<c�<ǂ~<X=z<��u<�q<�rm<6i<X�d<��`<��\<?�X<aT<�EP<-L<�H<N�C<��?<Z�;<ڧ7<m�3<2`/<V9+<�'<m�"< �<H�<�<dn<z]<�S
<�Q<�V<k��;���;(�;�j�;���;�;s�;���;X�;}޷;w�;%�;��;�ך;"�;?�;z��;��;/�s;˨g;�[;"�P;J�E;@7;;�0;��&;)G;��;{�
;��;��:���:�!�:��:r�:-Z�:E��:���:��m:AyS:W�9:�� :��:ߠ�9�Ҳ9,��9�A-9�e�8����&˸ٙA��ڎ�*缹���A,���"��8���N��d�y�����u͐�/����s���)���ڷ�/���|m˺gaպr}ߺ-���$��e���(����	��P�Ħ�����<��w$��)�%�.���3�8�8�8	>��C��/H�mPM��R���W��]��b�� h�׍m��&s��x�o]~�����p����q���������U��:⑻�f���斻,e���  �  ġ=�Q=� =��=j[=�=�=wZ==\� =�S =���<�H�<��<s��<�B�<���<>��<PF�<���<S��<;J�<|��<���<Z@�<n��<���<��<�e�<���<���<X3�<y�<���<^
�<�V�<���<���<XI�<���<���</C�<���<7��<+�<�p�<���<���<�$�<�W�<���<S��<���<���<��<�3�<�J�<^]�<�j�<xr�<Zs�<�l�<�]�<�D�<�!�<���<	��<�p�<��<���<!P�<g��<QV�<���<�6�<u��<p��<oQ�<��<���<�8�<�z�<���<��<�<(D�<>e�<#�<?��<瞮<å�<��<��<;��<Ŗ�<G��<e��<�s�<�f�<VY�<�K�<>�<�/�<� �<��<���<��<fԉ<��<���<��<{^�<�v~</z<1�u<1�q<�^m<�!i<��d<�`<��\<|mX<PT<�6P<_ L<6H<}�C<V�?<��;<˧7<
�3<�e/<=A+<'<V�"<��<��<��<��<Wq<g
<*d<gh<Y��;��;�=�;�{�;J��;W�;t�;���;�N�;Mз;�c�;I�;#ҡ;���;R��;)��;Y�;��;�hs;\^g;l�[;�yP;��E;�;;��0;��&;�7;��;.�
;�;���:���:T}�:�y�:��:��:
S�:\9�:�!o:��T:{�::��!:Rz	:E�9n�9La�9�E.9��8x�"��"͸X6C��􏹌N���}칈(�V�#�j:�!�O�yce�aOz��`��-d���9�� ȑ��k0�� �����˺}|պ�ߺڮ����tp���|���	�<��d��������*$��[)��.��3���8�D�=��B��H��9M�fsR�ǿW�; ]�M�b��h�`�m��Vs�'�x�M�~�/������?����G���茻<}������������}���  �  Ɵ=KP=��=;�=c[=F=�=�[==ɭ =]V = ��<�O�<f��<���<HJ�<w��<p��<�K�<*��<��<�L�<"��<N��<@�<%��<���<��<�a�<���<���<�,�<�q�<ظ�<_�<�N�<���< ��<vB�<���<>��<�>�<��<���<m)�<�o�<���<���<'�<�Z�<4��<f��<���<& �<��<+;�<:R�<�d�<`q�<Xx�<lx�<�p�<�`�<�F�<�"�<���<2��<�n�<�<���<OK�<���<�O�<���</�<2��<���<I�<���<E��<�1�<it�<���</�<h�<�A�<�c�<n~�<u��<$��<��<說<o��<t��<Ĝ�<뒢<���<({�<n�<g`�<NR�<�C�<�4�<%�<��<�<�<�ԉ</��<�<}�<�Z�<pm~<�#z<R�u<�q<�Om<�i<�d<��`<	�\<_X<�BT<'+P<sL<�H<v�C<�?<I�;<��7<��3<<i/<G+<�#'<)#<�<��<��<�<��<Uv
<_r<iu<���;��;�M�;���;R��;@�;\t�;���;nG�;0ŷ;dT�;���;Ȼ�;���;ͥ�;k،;5:�;�;�+s;�$g;f�[;NIP;�mE;��:;&�0;�&;�+;��;H�
;��;x�:M2�:��:���:�R�:5P�:XǓ:�:?p:1�U:{�;:̪":!
:�)�9�δ9���9T�.9qg�8��'���θ�kD�{֐�n����������$�b	;���P��ef��O{�U݇�Pؑ�����:N���⮺�u��º`�˺��պ�ߺ������G���_�$�	�,���3��x� ��4�#�� )��J.�o3���8�í=���B���G��)M��kR�s�W��']�G�b��3h�i�m�s|s��(y���~�38������幇�;h��r��ě��8#��	������ꐙ��  �  ��=EO= �=٭=T[=�=��=�\=D=P� =%X =�  =T�<ئ�<H��<�N�<���<T��<=O�<��<K��<�N�<0��<���<�?�<C��<��<w�<�^�<J��<1��<�(�<;m�<���<n��<�I�<ʘ�<f��<>�<ϒ�<���<�;�<���<���<?(�<[o�<ݱ�<���<x(�<�\�<Ό�<���<m��<@�<$�<�?�<�V�<�h�<}u�<|�<�{�<�s�<�b�<RH�<\#�<��<���<�m�<"�<3��<@H�<+��<�K�<���<*�<��<���<�C�<���<^��<-�<fp�<���<:�<��<�?�<\b�<�}�<���<���<~��<<"��<���<���<��<��<��<r�<�d�<^V�<�G�<8�<�'�<��<b�<��<�ԉ<���<���<{�<3X�<fg~<�z<<�u<�q<�Em<�i<��d<�`<:w\<�UX<Y:T<�#P<L<��G</�C<$�?<��;<*�7<��3<�k/<�J+<�('<Y#<D�<��<��<7�<ŉ<y
<4{<�}<-�;>,�;�W�;��;q��;�;7t�;4��;B�;k��;�J�;��;ǭ�;���;��;�Ō;)'�;�u;s; g;rc[;G+P;�RE;y�:;b�0;4�&;h#;��;&�
;��;�/�:_R�:���:��:[��:뒢:v�:���:�p:�V:�J<:�"#:�
:w��9�O�9sU�9�X/9���8˛+�k�ϸlNE�Ai���$������i�	5%���;�F�Q�g��{�_+���"���蛺L���x������f2º��˺١պ��ߺe�����Y.���N���	�������V����X�#�6�(�E(.��N3��q8�Ŕ=��B��G��M�^fR�˿W�G-]��b��Ch�B�m���s�qEy���~�&J�� ���͇�"|��4��
���U5��p����(��\����  �  !�=�N=��=��=@[=�=ϲ=]=�=̯ =�X =� =�U�<}��<��<AP�<,��<���<[P�<���<��<O�<p��<���<�?�<���<���<��<%^�<��<���<	'�<�k�<P��<���<�G�<��<���<�<�<q��<{��<�:�<��<=��<�'�<"o�<Ա�<���<�(�<s]�<���<���<���<��<�%�<GA�<^X�<Sj�<�v�<;}�<�|�<jt�<\c�<�H�<�#�<���<D��<Fm�<|�<u��<>G�<���<EJ�<[��<b(�<I��<���<�A�<Д�<���<w+�<�n�<���<P�<:�<?�<�a�<�}�<���<"��<���<���<��<Ѩ�<Ρ�<���<���<_��<)t�<.f�<�W�<�H�<	9�<m(�<w�<��<��<wԉ<P��<M��<yz�<|W�<Qe~<@z<m�u<��q<�Bm<i<5�d<M�`<�s\<�RX<r7T<(!P<�L<�G<��C<C�?<�;<Ц7<�3<'l/<�K+<l*'<P	#<��<r�<��<��<f�<��
<E~<\�<��;L0�;[�;���;���;��;�s�;Y��;q@�;$��;�G�;(�;ب�;��;��;K��; �;3g;��r;��f;tW[;� P;IE;�:;B�0;Ѽ&;� ;u�;%�
;G�;7�:�]�:~��:��:���:^��:�$�:$�:��p:�HV:2x<:�J#:��
:n�9�|�9�r�9�r/9K��8�c-�g"иN�E�v���y`��M���!f%���;���Q��?g��)|��E���;��� ��m����*��N����<ºA�˺ݦպ��ߺ۟�2��&���H��	�*���
�9K����=�#���(��.��C3��h8��=�8�B���G��M�}eR���W�9/]��b�tHh��m�"�s��Oy�#�~�XP��s���ԇ�����^#�������;�����	.�������  �  ��=EO= �=٭=T[=�=��=�\=D=P� =%X =�  =T�<ئ�<H��<�N�<���<T��<=O�<��<K��<�N�<0��<���<�?�<C��<��<w�<�^�<J��<1��<�(�<;m�<���<n��<�I�<ʘ�<f��<>�<ϒ�<���<�;�<���<���<?(�<[o�<ݱ�<���<x(�<�\�<Ό�<���<m��<@�<$�<�?�<�V�<�h�<}u�<|�<�{�<�s�<�b�<RH�<\#�<��<���<�m�<"�<3��<@H�<+��<�K�<���<*�<��<���<�C�<���<^��<-�<gp�<���<:�<��<�?�<\b�<�}�<���<���<~��<<"��<���<���<��<��<��<r�<�d�<^V�<�G�<8�<�'�<��<a�<��<�ԉ<���<���<{�<3X�<fg~<�z<<�u<�q<�Em<�i<��d<�`<:w\<�UX<Z:T<�#P<L<��G<0�C<$�?<��;<*�7<��3<�k/<�J+<�('<Y#<D�<��<��<7�<ŉ<y
<4{<�}<-�;=,�;�W�;��;p��;�;6t�;3��;B�;k��;�J�;��;ǭ�;���;��;�Ō;)'�;�u;s; g;qc[;F+P;�RE;y�:;a�0;4�&;h#;��;&�
;��;�/�:_R�:���:��:[��:뒢:v�:���:�p:�V:�J<:�"#:�
:w��9�O�9sU�9�X/9���8˛+�k�ϸlNE�Ai���$������i�	5%���;�F�Q�g��{�_+���"���蛺L���x������f2º��˺١պ��ߺe�����Y.���N���	�������V����X�#�6�(�E(.��N3��q8�Ŕ=��B��G��M�^fR�˿W�G-]��b��Ch�B�m���s�qEy���~�&J�� ���͇�"|��4��
���U5��p����(��\����  �  Ɵ=KP=��=;�=c[=F=�=�[==ɭ =]V = ��<�O�<f��<���<HJ�<w��<p��<�K�<*��<��<�L�<"��<N��<@�<%��<���<��<�a�<���<���<�,�<�q�<ظ�<_�<�N�<���< ��<vB�<���<>��<�>�<��<���<m)�<�o�<���<���<'�<�Z�<4��<f��<���<& �<��<+;�<:R�<�d�<`q�<Xx�<lx�<�p�<�`�<�F�<�"�<���<2��<�n�<�<���<OK�<���<�O�<���</�<2��<���<I�<���<E��<�1�<it�<���<0�<h�<�A�<�c�<n~�<u��<%��<��<說<o��<t��<Ĝ�<뒢<���<({�<n�<g`�<NR�<�C�<�4�<%�<��<�<�<�ԉ</��<�<}�<�Z�<pm~<�#z<R�u<�q<�Om<�i<�d<��`<	�\<_X<�BT<(+P<sL<�H<v�C<�?<J�;<��7<��3<=i/<G+<�#'<*#<�<��<��<�<��<Uv
<_r<hu<���;��;�M�;���;Q��;>�;Zt�;���;lG�;/ŷ;bT�;���;ǻ�;���;̥�;j،;4:�;�;�+s;�$g;e�[;NIP;�mE;��:;%�0;�&;�+;��;G�
;��;w�:M2�:��:���:�R�:5P�:XǓ:�:?p:1�U:{�;:̪":!
:�)�9�δ9���9T�.9qg�8��'���θ�kD�{֐�n����������$�b	;���P��ef��O{�U݇�Pؑ�����:N���⮺�u��º`�˺��պ�ߺ������G���_�$�	�,���3��x� ��4�#�� )��J.�o3���8�í=���B���G��)M��kR�s�W��']�G�b��3h�i�m�s|s��(y���~�38������幇�;h��r��ě��8#��	������ꐙ��  �  ġ=�Q=� =��=j[=�=�=wZ==\� =�S =���<�H�<��<s��<�B�<���<>��<PF�<���<S��<;J�<|��<���<Z@�<n��<���<��<�e�<���<���<X3�<y�<���<^
�<�V�<���<���<XI�<���<���</C�<���<7��<+�<�p�<���<���<�$�<�W�<���<S��<���<���<��<�3�<�J�<^]�<�j�<xr�<Zs�<�l�<�]�<�D�<�!�<���<	��<�p�<��<���<!P�<h��<QV�<���<�6�<u��<q��<oQ�<��<���<�8�<�z�<���<��<�<)D�<?e�<#�<?��<螮<ĥ�<���<��<<��<Ŗ�<H��<f��<�s�<�f�<VY�<�K�<>�<�/�<� �<��<���<��<fԉ<��<���<��<{^�<�v~</z<1�u<0�q<�^m<�!i<��d<�`<��\<}mX<PT<�6P<` L<7H<~�C<W�?<��;<̧7<�3<�e/<>A+<'<V�"<��<��<��<��<Wq<g
<*d<fh<X��;��;�=�;�{�;I��;U�;t�;���;�N�;Kз;�c�;G�;!ҡ;���;Q��;(��;
Y�;��;�hs;Z^g;j�[;�yP;��E;�;;��0;��&;�7;��;.�
;�;���:���:T}�:�y�:��:��:
S�:\9�:�!o:��T:{�::��!:Rz	:D�9n�9La�9�E.9��8y�"��"͸X6C��􏹌N���}칈(�V�#�j:�!�O�yce�aOz��`��-d���9�� ȑ��k0�� �����˺}|պ�ߺڮ����tp���|���	�<��d��������*$��[)��.��3���8�D�=��B��H��9M�fsR�ǿW�; ]�M�b��h�`�m��Vs�'�x�M�~�/������?����G���茻<}������������}���  �  >�=�S==^�=_[='=ï=}X= =-� =�O =-��<�?�<���<���<}9�<���<���<?�<a��<h��<�F�<��<���<�@�<���<���<�#�<
k�<��<Q��<�;�<^��<z��<��<a�<���<@ �<@R�<��<}��<�H�<N��<���<C-�<sq�<��<���<�!�<>S�<c��<���<���<��<p�<T*�<gA�<2T�<>b�<�j�<�l�<%g�<=Y�<�A�<��<n��<���<s�<c �<T��<,V�<���<�^�<��<�@�<���<?�<<\�<_��<���<�A�<���<���<��<� �<�G�<ag�<��<���<���<���<��<R��<F��<���<���<w�<Fj�<)]�<.P�<BC�<P6�<>)�<l�<��<���<L�<ԉ<���<��<8��<<c�<Ƃ~<X=z<��u<�q<�rm<6i<X�d<��`<��\<@�X<aT<�EP<-L<�H<N�C<��?<[�;<ۧ7<n�3<3`/<V9+<�'<n�"<!�<H�<�<dn<z]<�S
<�Q<�V<i��;���;(�;�j�;���;�;s�;���;X�;{޷;w�;%�;��;�ך;!�;>�;y��;��;-�s;ɨg;
�[; �P;I�E;?7;;�0;��&;(G;��;z�
;��;��:���:�!�:��:r�:-Z�:E��:���:��m:AyS:W�9:�� :��:ߠ�9�Ҳ9,��9�A-9�e�8����&˸ٙA��ڎ�*缹���A,���"��8���N��d�y�����u͐�/����s���)���ڷ�/���|m˺gaպr}ߺ-���$��e���(����	��P�Ħ�����<��w$��)�%�.���3�8�8�8	>��C��/H�mPM��R���W��]��b�� h�׍m��&s��x�o]~�����p����q���������U��:⑻�f���斻,e���  �  ��=�U=[=�=?[=>=�=V=\� =N� =NK =+��<�4�<G��<[��<U.�<��<,��<Y6�<���<z��<B�<��<��<�@�<S��<}��<5(�<�p�<E��<���<�E�<��<���<s �<�l�<H��<N�<i\�<��<e��<tO�<N��<B��<D/�<%r�<E��<v��<�<�M�<�y�<z��<���<���<��<�<6�<LI�<�W�<Va�<~d�<``�<	T�<>�<��<���<��<Ou�<Q$�<���<�\�<���<h�<���<uL�<5��<��<�h�<��<U�<GL�<7��<!ƻ<R��<�%�<:K�<di�<���<Ӑ�<���<���<���<P��<���<F��<y�<l�<�^�<�Q�<FE�<9�<3-�<9!�<��<i�<[��<$�<vӉ<̼�<G��<!��<|h�<v�~<�Mz<O
v<]�q<"�m<�Mi<me<��`<��\<��X<ltT<�VP<�;L<� H<D<9�?<��;<��7<��3<�Y/<�/+<�'<��"<�<ێ<�o<HW<�E<n<
<F;<�B<̣�;���;,�;�V�;���;��;#q�;,��;�a�;S�;X��;�@�;��;b��;�;,H�;#��;�B�;tt;�g;GM\;i�P;�F;�h;;�1;�';�T;
�;��
;��;g~�:\�:C��:��:Dܯ:v��:R�:u�:�|l:R:��8:��:��:t��9�t�9䏃9,9t�8̪�@Xɸ+�?�X���bR��@���@t!���7�SGM���b�f�w��	��� ��d��꣺����z��SO���;˺qIպ�yߺ��麩Q������2���2
�������J������$�~*�-#/��74�bB9�hH>�rMC��WH�lM���R���W��]�"ob���g�>cm�{�r��x�.~�E΁������B��ϐ���(��F���A���Ŗ��H���  �  ͩ=�W=�=i�=�Z==4�=HS=�� =� =nF =E��<#)�<z�<���<*"�<[y�<���<�,�<Ň�<���<�<�<���<��<S@�<���<W��<�,�<�v�<Ϳ�<��<�O�<S��<���<�,�<vy�<���<��<?g�<���<��<,V�<o��<���<D1�<�r�<���<���<��<�G�<3r�<���<���<���<���<��<�)�<`=�<�L�<>W�<�[�<�X�<	N�<�9�<��<���<���<�w�<.(�<��<d�<y��<&r�<��<�X�<��<��<�u�<@��<V�<jW�<��<tλ< �<+�<�N�<qk�<��<z��<���<�<g��<���<݆�<�z�<�m�<`�<�R�<�E�<Z9�<�-�<9#�<p�<��<��<&�<~�<e҉<u��<x��<���<�m�<s�~<�^z<0v<��q<Рm<�fi<�0e<��`<��\<T�X<�T<�hP<�JL<�,H<�D<��?<?�;<��7<�}3<3R/<�$+<��&<��"<5�<�x<�W<(><@,<>#
<#<1,<�{�;Ю�;%��;�?�;|��;���;�m�;7��;�j�;���;��;�\�;m0�;�#�;*9�;5v�;3ކ;?s�;Tot;NWh;��\;0FQ;�EF;��;;�?1;�/';�b;Q�;B�
;ss;H4�:���:V8�:E��:18�:���:�K�:� �:��j:��P:�7:�p:Xm:n��9,�9�e�9Q�*9Y��8W��^�Ǹ�(>�Bg������\�湒�	�/ �
6��K��a�?�u��H��Xk���j���W��,6��~�� ��?˺}1պ�{ߺL�����$?�����r
�����G�������6%��d*�M�/���4�d�9���>���C���H�c�M���R�(�W�\	]��\b��g��7m�%�r�->x���}�C����]��*��˼��_����������������",���  �  ��=�Y=�=��=[Z=�=�=nP=9� =�� =]A ='��<I�<�m�<_��<��<�m�<���< #�<]�<���<t7�<ő�<���<�?�<���<���<�0�<�|�<��<��<�Y�<g��<���<<9�<݅�<���<g"�<�q�<���<w�<�\�<]��<��<3�<�r�<l��<���<��<�A�<|j�<`��<:��<8��<���<\�<d�<N1�<eA�<�L�<eR�<EQ�<�G�< 5�<��<M��<���<�y�<�+�<V��<�j�<���<�{�<���<�d�<���<+�<��<���<2�<&b�<���<xֻ<��<�/�<R�<2m�<��<㍰<���<%��<���<���<p}�<Lp�<1b�<�S�<F�<(9�<a-�<�"�<��<j�<��<t��<��<��<�Љ<���<j��<i��<s�<߫~<�nz<d1v<�q<m�m<�i<Je<�a<��\<|�X<��T<�yP<�XL<.8H<�D<��?<��;<��7<�x3<�I/<'+<,�&<�"<��<�a<~?<�$<Y<�	
<�
<D<(R�;���;��;�'�;���;S��;eh�;���;�r�;I�;:��;jw�;OQ�;yI�;�c�;���;��;��;��t;�h;	�\;��Q;;�F;��;;�d1;�F';-n;_�;�x
;�X;~��:��:���:e_�:���:3E�:I��:�V�:�Zi:PO:��5:P:@:T��9�E�9C,�9w�(9�0�8\ ���Ÿ��<��8��������������,�4��=J�r�_��pt����e����ɘ��ɢ�;�������ؿ����ʺ:պ�ߺ�����l����;�δ
�j-�ߞ��XY �i�%�v�*���/���4���9���>��C���H�f�M���R�/�W�]��Kb���g�Fm��r�-�w�Fw}�dw���.��k������<.��tʎ��`��	�l���~���  �  �=5[=�=̰=�Y=z=��=�M=�� =�� =�< =���<��<�a�<|��<
�<b�<;��<��<Nw�<
��<62�<֍�<���<�>�<'��<���<Z4�<���<���<~�<�b�<���<���<�D�<O��<���<�,�<A{�<r��<��<Tb�<���<���<?4�<Tr�<ݫ�<g��<A�<�;�<�b�<���<j��<n��<��<���<��<�%�<�6�<�B�<�I�<�I�<�A�<�0�<��<���<���<�z�<�.�<���<�p�<X �<Մ�<���<�o�<u��<7�<��<z��<')�<�k�<H��<�ݻ<��<D4�<�T�<^n�<���<B��<'��<s��<���<
��<�t�<Hf�<AW�<@H�<1:�<R-�<�!�<��<%�<��<���<���<	�<�ދ<�ω<���<ݨ�<V��<�w�<ѷ~<~z<�Bv<�r<�m<"�i<Xae<�/a<�]<��X<�T<щP<�eL<0BH<�D<o�?<�;<��7<�s3<�A/<+<��&<�"<[w<wL<Y(<S<��<[�	<~�<��<P+�;�h�;���;��;�v�;��;�b�;���;�x�;m�;�ɰ;���;Io�;�k�;���;�͍;9�;(π;#"u;�i;j:];��Q;1�F;C�;;�1;<Z';�u;��;.j
;N=;���:8-�:{=�:�ҽ:��:���:`Ώ:ʗ�:��g:H�M:J4:��:%:a�9���9��9u''9�q�8���a�ĸ�_;��4��\���G*�Q��'���]3���H�0^�ws��ك�.���6���G���T���d��w����ʺ�պ/�ߺ�2�,��������p�t�
�(v�����\�� �|�%�>'+��<0��>5�j0:�2?���C�y�H���M�%�R�x�W�]�X?b���g�s�l��Pr��w��1}�3P���������>]��W��@����8���Γ��b�������  �  ް=�\=B=Ͱ=!Y=, =�=!K=�� =ߓ =o8 =a��<�<�W�<5��<���<�X�<-��<��<<p�<��<v-�<M��<B��<�=�<w��<���<B7�<��<���<�<�j�<6��<��< N�<��<$��<�5�<w��<���<��<
g�<��<��<#5�<�q�<��<f��<�<E6�<]\�<�<ƞ�<��<;��<`��<m�<��<,-�<M:�<B�<:C�<�<�<{,�<��<E��<i��<|�<1�<���<�u�<��<C��<��<y�<H��<5A�<��<8��<Z2�<at�<���<��<W�<�7�<&W�<Ao�<H��<n��<��<&��<*��<Yz�<�l�<~]�<�M�<N>�<�/�< #�<�<��<��<O��<��<E��<��<�ۋ<�͉<R��<海<œ�<K{�<��~<_�z<�Qv<�r<0�m<F�i<�te<�Ba<]<&�X<��T<ݖP<{pL<^JH<F#D<k�?<��;<C�7<~n3<:/<�+<[�&<C�"<Xf<�9<8<{�<��<��	<C�<��<��;�J�;!��;���;�f�;���;�\�;0��;�}�;J"�;|ذ;���;އ�;V��;^��;���;�]�;=�;:ju;�Ei;{y];�R;H�F;�<;ٝ1;j';�z;��;�Z
;�#;�Q�:%��:@��:hU�:Qa�:7��:.�:h�:�f:�UL:�3:�:�):�Z�9;P�9�}99�%9���8$m!��7ĸ�T:��_��ŗ��0�ṟ��ܡ��D2��G��\�M�q��F�����������ܡ���� ���S����ʺ�պ��ߺ3V��3��� �G���+����:8�/��_!��L&��x+��0�H�5�at:��S?�/D��I� �M��R�(�W�%]��5b�Zxg�f�l� )r���w���|��.��
���܍���6��Uۋ�{���������~I��+㘻�  �  J�=r]=�=��=�X='�=��=I=#� =�� =*5 =K��<x �<�O�<��<��<1Q�<5��<8�<�j�<h��<�)�<���<n��<�<�<���<���<O9�<���<��<$�<zp�<���<��<|U�<H��<w��<�<�<���<���<#!�<�j�<���<|��<�5�<q�<���<$��<��<�1�<JW�<y�<��<ô�<w��<i��<r��<-�<�%�<�3�<<�<*>�<38�<3)�<��<���<��<�|�<�2�<O��<�y�<X�<ܑ�<��<��<���<�H�<ʠ�<���<A9�<�z�<���<q�<��<W:�<�X�<�o�<��<���<ȋ�<���<ŀ�<u�<�f�<�V�<LF�<{6�<�'�<'�<U�<l�<���<_��<�<�<��<|ً<�̉< ��<���<j��<�}�<B�~<Ǔz<�\v<0%r<�m<*�i<ǃe<�Qa<:"]<�X<�T<ʠP<�xL<\PH<:'D<C�?<��;<9�7<�j3<=4/<��*<��&<��"<Y<7+<�<,�<�<0�	<��<:�<��;3�;���;��;�Z�;��;�W�; ��;N��;$)�;|�;���;���;H��;�Ô;%�;8z�;��;��u;/yi;=�];�-R;�G;5<;O�1;4t';"};	�;�M
;o;��:��:�:�:t��:]��: ��:Aq�:�e:CYK:�*2:��:�c:��92�9|9ba$9���8:�%���øȪ9��ň�,���0��*�R���p1���F���[���p��ӂ�� ���Z��񋡺Ӹ��~쵺�0���ʺ�	պ�ߺ�q�3]���4 �/��VW�)��{o�>���F!���&���+���0�w�5�=�:���?�~VD�-I�q
N��R���W��]��0b��jg���l��
r��hw�d�|�����ă�jp��W��꽋�__������<���I6���Ә��  �  (�=^=�=��=-X=p�=��=�G=�� =/� =3 =���<���<�J�<��<%��<mL�<���<9�<'g�<g��</'�<���<%��<(<�<���<O��<�:�<׊�<���</'�<t�<���<H�<�Y�<Ħ�<���<�@�<a��<B��<�#�<�l�<.��<r��<�5�<q�<���<y��<��<//�<�S�<Iu�<ѓ�<"��<���<��<���<U�<C!�<X/�<P8�<�:�<z5�<	'�</�<	��<ȹ�<#}�<�3�<���<�{�<I�<h��<��<u��<���<�M�<��<f��<�=�<�~�<p��<E�<�<�;�<�Y�<p�<o�<���<��<s��<�}�<�q�<�b�<`R�<�A�<�1�<�"�<7�<v�<��<���<���<��<S�<��<�׋<�ˉ<���<���<v��<��<��~<��z<�cv<-r<��m<�i<�e<�Za<�*]< �X<U�T<�P<w}L<TH<�)D<��?<��;<��7<�g3<"0/<��*<I�&<N�"<�P<�!<��<�<��<�	<��<��<A��;$�;{�;k��;�Q�;��;HT�;@��;C��;v-�;�;廩;\��;��;LӔ;��;M��;�!�;u�u;��i;��];ZGR;�G;hE<;��1;�z';;�;,E
;S;���:S_�:�H�:���:��:9<�:ga�:�!�:��d: �J:9�1:�Z:?�:3�9�|�9�z9p�#9��8P�)��øK99�Tg��l7����߹˿��h���0��=F��d[�cXp�����ߌ� ��dX������ε�[����ʺպ˳ߺ?��Q{���G ����Zs���ے�*��m!�]�&�I�+���0�1�5���:��?�2pD�BI�zN� S���W��
]��,b��ag�A�l���q�bQw���|��������^��e��+���ON���퐻���;*��=ʘ��  �  D�=mW=� =��=/Q=��=��=�B=�� =G� =/1 =j��<(��< I�<l��<���<E�<ĝ�<���<S�<g��<i	�<0c�<���<��<)f�<C��<_�<�V�<���<z��<�:�<*��<]��<��<�c�<��<~��<-?�<��<P��<��<�S�<��<���<j�<&:�<Yi�<���<y��<���<?��<��<�4�<�K�<�`�<�r�<��<?��<E��<̕�<֐�<c��<@o�<hP�<s'�<N��<��<�h�<��<!��<�D�<���<�L�<M��<�.�<Ò�<x��<IB�<ߎ�<%Ծ<h�<�I�<�z�<l��<yǵ<��<���<u	�<!�<��<��<�<��<v�<G��<�<�<K�<|ۙ<�՗<�Е<�˓<,Ǒ<���<��<���<_��<���<���<z{�<�h�<��~<�{z<�Nv<� r<�m<��i<-�e<oa<�F]<�Y<o�T<d�P<1�L<S�H<lD<H@<�!<<�7<+�3<"�/<�y+<�N'<�%#<Z <K�<��<n�<Ƭ<��
<�<��<���;`,�;��;���;�u�;J��;Ӓ�;"4�;���;y��;Tv�;�]�;h^�;�z�;���;1�;�;�5�;|;��o;x!d;�X;H�M;��B;�8;��-;��#;�;�};>2;`I�:J��:C~�:,��:P��:'�:��:K��:;{:�$`:'F:)�,:Qs:�*�9&h�9�W�9�|]99-�#8e2D���
��ud�C�ׅ˹x��������'�c�=��S�~lh�l�}�YT��O̓�h;�������������Ⱥ�Һ�wݺ{N��@�D��J��8
�����@�C��r ��d%�ћ*��/�l�4���9��>�ѾC�_�H�3�M�űR���W��\�b�iSg�M�l���q�qNw���|���������c��}�����5_��S��먓��M�����  �  ��=KW=� =��=BQ=��=�=(C= � =�� =�1 =���<I��<~J�<���<���<>F�<��<���<�S�<&��<�	�<�c�<Ի�<�<)f�<��<
�<;V�<���<���<�9�<��<B��<A�<*b�<��<b��<@>�<!��<���<0�<rS�<���<���<w�<K:�<�i�<���<��<j��<%��<��<�5�<)M�<b�<-t�<��<i��<^��<���<���< ��<�o�<�P�<�'�<T��<ӳ�<�h�<>�<w��<�C�<���<�K�<��<�-�<T��<��<A�<���<&Ӿ<��<&I�<�y�<���<Gǵ<��<���<�	�<��<>�<e�<��<��<��<f��<T��<��<��<�ܙ<�֗<�ѕ<�̓<ȑ<j<���<��<���<���<���<>{�<h�<_�~<�zz<Mv<�r<��m<x�i<c�e<ma<xD]<�Y<��T<��P<αL<$�H<�kD<�G@<�!<<J�7<��3<�/<�z+<CP'<�'#<�<��<#�<;�<�<S�
<]�<��<���;;0�;H��;��;x�;���;���;`4�;\��;a��;"t�;r[�;�[�;Ow�;|��;��;���;�0�;Y�{;H�o;hd;��X;�|M;�B;s8;x�-;��#;�;";�5;nQ�:v��:���:���:Hȸ:`/�:8"�:E��:�F{:�K`: @F:�-:�:nd�9@��9w�9��]9�!9��#8�?D�+�
�M�d�w����˹���{���'�W�=��=S��h���}�f��#ۓ�uG��򰨺���l����Ⱥ��Һ�uݺ�J�(9�0<������0
�����7�(��A �aX%���*��/�'�4�F�9���>��C�­H�+�M��R�q�W���\�b�`Ug���l��q�PTw�f�|��
��Z���\h���������c��^��Y����P��r����  �  I�=�V=� =��=�Q=|�=��=D=)� =� ==3 =���<���<N�<���<���<�I�<=��<���<�V�<]��<��<e�<���<v�<f�<���<�<�T�<��<R��<�6�<��<
��<��<�^�<���<7��<T;�<���<w��<��<3R�<��<9��<��<�:�<�j�<���<��<���<��<�<G9�<�P�<�e�<�w�<���<��<���<x��<&��<���<Eq�<�Q�<'(�<w��<h��<�g�<��<���<�A�<��<�H�<ǽ�<*�<ʍ�<���<�=�<a��< о<��<G�<;x�<���<qƵ<��<��<N
�<��<��<r�<c�<k�<�	�<� �<���<"�<=�<8��<Dڗ<�ԕ<�ϓ<qʑ<_ď</��<&��<!��<ћ�<-��<lz�<�f�<�~<vz<�Gv<�r<e�m<�i<��e<\fa<�=]<�Y<�T<"�P<�L<8�H< jD<�F@<�!<<2�7<��3<�/<�~+<�T'<	-#<�<��<{�<��<=�<��
<��<��<x��;N;�;Ϙ�;��;M~�;��;ו�;�4�;���;���;�n�;�T�;�R�;�l�;���;� �;J�;�#�;��{;��o; d;�X;�lM;ԖB;O8;��-;��#;�;��;�?;l�:���:ִ�:;�:v��:h�:�[�:jً:�{:��`:��F:�u-:��:��9J�9���9�S^9�z9�($8��D�S��De�񀟹�6̹y����r�ia(��>���S��i�k*~�����U��tn��Ш�6��¥��q'Ⱥ��ҺDpݺ�=躎#�5 ��E��T
����j��������;%�/t*�S�/���4���9��>�"�C�z�H�ٜM���R� �W��\��b�2\g�^�l��r�=fw���|����!ǃ�[u��[!��ʋ�mp�����9����Y�������  �  '�=V=M =��=�Q=9�=��=�E=�� =8� =�5 =#��<��<�S�<���<q��<wO�<J��<� �<�Z�<Դ�<��<g�<
��<�<�e�<���<^�<PR�<���<���<�2�<'|�<���<o�<OY�<<��<+��<�6�<}�<��<��<4P�<���<���<��<�;�<�l�<��<O��<���<t�<�#�<�>�<}V�<�k�<�}�<q��<@��<]��<���<���<'��<�s�<�S�<)�<���<ز�<�f�<��<ȫ�<>�<���<�C�<~��<T$�<���<���<�7�<,��<`˾<�
�<�C�<mu�<���<Bŵ<�<W��<\�<t�<q�<��<B�<��<��<h�<���<��<+�<�<�ߗ<�ٕ<ԓ<(Α<�Ǐ<���<ŵ�<��<���<���<y�<�d�<�~<�nz<]?v<hr<��m<��i<k�e<#[a<B3]<�Y<i�T<��P<ۧL<s�H<�fD<$E@<�!<<��7<��3<_�/<��+<+\'<�5#<c<�<6�<��<��<��
<��<y�<O�;�L�;���;]�;Q��;:
�;Q��;G5�;`��;f��;&f�;�H�;�D�;<\�;=��;(�;%j�;��;Z�{;(�o;}�c;JqX;�RM;	�B;��7;|�-;A�#;�	;�;�M;���:��:B��:=^�:�J�:���:���:�9�:Nz|:�za:`G:<.:O�:��9��9%��9�4_9-9f�$8��E����8f��+��4͹h���+�)��>��XT�}�i���~�)扺RO��뫞�e��&^�������5Ⱥ��ҺhݺN)�g����z�.�	�|�N��b�����%��D*�k/���4�"�9��>��C���H���M�A�R�g�W�(�\�(b�\gg���l�Kr���w��|��)���ۃ�a���n7��#���]����'��ȓ�+h���	���  �  ��=U=��=}�=SR=3�=$�=vG=A� =�� =�8 =���<��<n[�<-��<� �<�V�<���<��<�_�<@��<�<�i�<ſ�<��<�e�<Y��<�<O�<Ù�<���<�,�<�u�<ݾ�<U�<&R�<?��<���<�0�<z�<w��<	�<vM�<��< ��<�</=�<�n�< ��<T��<y��<.�<`*�<�E�<�]�<s�<(��<���</��<ǣ�<���<���<#��<�v�<�U�<B*�<���<��<�d�<��<٧�<19�<*��<R=�<���<��<j��<2��<�0�<F~�<ž<C�<�>�<�q�<靷<võ<H�<���<��<��<��<�!�<D �<��<9�<j�<��<���<���<?�<r�<��<�ٓ<�ґ<vˏ<�<뷋<&��<��<���<#w�<�a�<]�~<eez< 4v<�r<u�m<��i<�ve<�La<�%]<� Y<��T<��P<��L<�H<QbD<�B@<5!<<+�7<Z�3<�/<�+<me'<�@#<+<<��<�<f�<5�
<W�<z�<�;Cc�;Ϻ�;� �;*��;��;H��;?5�;i��;z��;|Z�;{9�;�1�;�E�;�z�;Ґ;�N�;'�;��{;ioo;�c;�GX;0M;fB;`�7;�-;��#;�;=�;�`;���:6I�:B�:���:o��:�/�:/�:���:in}:�eb:�AH:��.:[<:�<�9Y��92T�9�_`9��9�q%8��F�f����g�r��|+ι������)���?��=U�B�j�9���M���������H�����_轺MȺ�Һ�_ݺ��=��~���NW���	��K�0��6)������$��*�J1/��J4�EX9�j^>�nbC�gH��sM�։R�S�W���\�E%b�^wg� �l��<r�ݨw��}��B����������T��i���J����@���ޓ��{������  �  ѧ=�S= �=`�=�R=*�=��=�I=�� =� =J< =���<:�<*d�<��<�	�<�^�<���<��<�e�<Z��< �<�l�<g��<O�<e�<���<J �<'K�<���<x��<�%�<n�<���<���<�I�<���<���<Z)�<�s�<��<��<.J�<���<���<?�<O>�</q�<���<���<(��<��<�1�<�M�<6f�<�{�<ҍ�<,��<>��<��<��<^��<���<z�<�W�<@+�<���<���<+b�<L�<4��<`3�<j��<�5�<3��<G�<aw�</��<(�<v�<���<���<19�<2m�<���</��<7�<���<��</�<#�<�&�<&�<c"�<��<��<��<g�<c��<���<l�<E�<��<�ؑ<�Ϗ<�ō<��<0��<��<|��<�t�<9^�<,�~<�Yz<�&v<��q<>�m<��i<�ee<�;a<]<��X<�T<��P<��L<vyH<]D<d?@<� <<��7<�3<�/<`�+<9p'<MM#<z-<<*�<��<j�<6�
<��<�<�7�;�|�;���;2�;���;��;k��;�4�;��;	��;hL�;�&�;��;1,�;�]�;���;B.�;,҃;�@{;D2o;!zc;�X;�M;*EB;�7;V�-;��#;�;ȣ;[u;��:ӓ�:b��:$�:�*�:4��:��:�@�:�~:�zc:nHI:��/:x:���9��9\9�9��a9C]9K&8��H���Gi�
#��̅Ϲ������A�*��@��OV�F�k� \��8Ɋ����^`������Գ�����jȺ��Һ�Wݺ���>�������/��	�$������B?�Ɉ$���)���.�G4�(9�q,>��6C��DH�sYM�(yR��W�M�\��/b�Z�g�[�l��ar���w��L}�`�����Ɇ�bv��
�������^������
����,���  �  ��=ZR=$�=&�="S= �=S�=�K=�� =S� =@ =��<�<lm�<<��<��<�g�<׽�<��<Jl�<���<�<�o�<��<��<Qd�<���<!��<�F�<I��<���<[�<�e�<��<���<e@�<���<��<�!�<�l�<���<���<hF�<K��<���<?�<u?�<�s�<+��<~��<���<o�<9�<�U�<3o�<���<��<(��<���<��<���<"��<@��<�}�<;Z�<C,�<���< ��<�_�<N�<��< -�<��<�-�</��<�
�<�m�<���<��<1m�<���<p��<3�<%h�<Ж�<���<�߳<���<��<��<�&�<R+�<�+�<p)�<�$�<�<��<��<��<���<���<�<��<7ޑ<aԏ<aɍ<R��<;��<ۛ�<���<)r�<3Z�<��~<�Mz<zv<��q<��m<D�i<�Re<;)a<>]<�X<�T<~�P<ՊL<�pH<�VD<�;@<Q<<� 8<��3<v�/<�+<6{'<�Z#<�<<�"<@<��<��<C�
<�<�<�V�;��;l��;D�;��;'#�;k��;�3�;��;}�;J<�;��;9�;��;>�;��;F�;ٮ�;��z;%�n;>c;�W;��L;. B;�7;��-;��#;Z;��;��;"?�: ��:���:q��:ש�::�:
K�:�֍:��:՞d:XJ:��0:�:r/�9�U�9*�9@�b9l9Ug&8�K�����j��T����й�V��"���+�&�A�WtW���l�Zꀺ0O��Õ���˟��󩺕���K��|�Ⱥ�Һ�Pݺp��|��A����Sq	�!��|B�C�����7>$�ix)�7�.���3���8���=��	C��!H��>M��hR���W���\��<b�^�g��m���r�`x�*�}�����9��9톻:���SB���㎻�����`����A���  �  ��=�P=7�=ɨ=gS=�=Υ=�M=P� =�� =�C =@��<�%�<�v�<r��<��<Fp�<���<�<kr�<���<�<1r�<���<�<Tc�<���<���<:B�<���<#��<��<t]�<��<o��<7�<с�<y��<{�<pe�<۰�<���<B�<���<��<��<j@�<�u�<���<��<���<) �<A�<L^�<x�<��<��<��<��<y��<���<���<ƛ�<��<8\�<-�<��<t��<�\�< �<���<�&�<���<-%�<:��<2�<�c�<���<�<Jd�<@��<�<�,�<c�<ʒ�<���<^޳<a��<�<��<I*�< 0�<�1�<I0�<R,�<�&�<��<��<��<��<��<���<s�<��<�؏<�̍<U��<��<Z��<\��<9o�<$V�<�w~<�@z<�	v<n�q<�m<�mi<�?e<ra<S�\<>�X<��T<$�P<�L<�gH<5PD<�7@<�<<�8<'�3<M�/<~�+<߅'<�g#<�K<�3<? <�<�<�<�<^#<.u�;(��;l��;�U�;���;"+�;��;h1�;B��;q�;,�;���;��;��;�;�n�;��;�;$�z;i�n;? c;��W;��L;$�A;ږ7;�|-;��#;;�;؛;�w�:;-�:�Z�:z�:-%�:«:�ڜ:�i�:bm�:�e:iK:�1:��:�P :R��9��9id99��%8��M�g*�s�l������yҹ� ���.�,���B���X���m��z��bՋ����_9��P��Rg�������Ⱥ��Һ�Oݺ���%[���>��JA	������M]�Э���#��/)��_.���3�h�8���=���B�w�G��%M�zYR��W���\��Jb���g��2m���r�W;x�\�}�����[\��������Lg���������4��OƖ�W���  �  ��=<O=J�=e�=�S=��=�=�O=�� =y� =G =���<�-�<�~�<��<$�<Jx�<��<�"�<x�<0��<�!�<�t�<���<�<Yb�<^��<d��<�=�<��<���<r�<~U�<s��<���<R.�<'y�<6��<��<�^�<��<���<�>�<̈́�<���<c�<&A�<�w�<y��<&��<� �<P&�<�G�<f�<,��<{��<���<#��<���<[��<ͽ�<��<˟�<˃�<^�<�-�<]��<ի�<�Y�<&��<���<r �<���<9�<���<��<�Z�<��<�<�[�<x��<;�<�&�<$^�<�<;��<�ܳ<���<��<�!�<V-�<,4�<7�<�6�<a3�<e.�<�'�<X �<3�<��<��<V��<��<��<�܏<fύ<��<���<ɚ�<���<Rl�<>R�<;m~<�4z<��u<��q<;�m<\i<7.e<�a<2�\<?�X<\�T<}�P<�tL<U_H<�ID<�3@<�<<>8<�3<Y�/<�+<��'<ws#<bY<�B<�0<�#<U<I<|$<�2<ې�;w��;J�;ce�;���;�1�;ө�;/�;9��;ve�;>�;�;.Ѥ;Dם;���;N�;�ŉ;Ci�;`rz;�nn;��b;wW;�|L;�A;�z7;�h-;؛#;�;Q�;��;���:�p�:L��:3g�:j��:s?�:�^�:p�:%��:V�f:AeL:\�2:��:�� :���9�ӡ9�e9�9B%8igP��x���n������ӹY� �^��{�-�QD�ԶY��o�F��V��w���G�������Ǯ�����,�Ⱥ,Ӻ_QݺL�纞7����λ��	��o������hk��#���(��.�KJ3�Rp8�Ē=��B���G�^M�.LR���W���\�'Xb�P�g��Rm��r��kx�q�}�Ϳ���}���4��u㉻9���`(��[����P���ޖ�Ml���  �  ��=�M=W�=��=�S=`�=*�=6Q=�� =� =�I =��<�4�<��<.��<&+�<�~�<^��<(�<�|�<��<i$�<tv�<���<�<Ha�<F��<x��<:�<Z�<=��<	�<�N�<7��<)��<�&�<�q�<��<F�<�X�<ĥ�<���<e;�<U��<��<��<�A�<�x�<��<���<�<w+�<�M�<vl�<��<���<���<���<!��<T��<���<3��<0��<2��<h_�< .�<���<)��<�V�<���<��<�<E��<K�<"��<c��<�R�<���<i�<dT�<���< �<�!�<�Y�<���<���<]۳<w��<Y�<F#�<�/�<�7�<�;�<�;�<t9�<�4�<�.�<v'�<H�<q�<%�<<�<���<�<"��<�э<��<���<,��<��<�i�<�N�<\d~<*z<s�u<F�q<�m<Mi<�e<��`<��\<`�X<��T<P�P<JkL<�WH<�CD<�/@<�<<|8<V�3<��/<�+<��'<m}#<e<�O<�><�2<,<�+<d2<�?<\��;���;"�;Qr�;���;*7�;B��;F,�;=��;$[�;�;}׫;��;�;K�;_2�;降;�K�;�9z; 8n;��b;�HW;SUL;n�A;�a7;{V-;�#;�;��;��;)��:���:}��:���:���:���:Ν:Xf�:'j�:j�g:�7M:�p3:�>:u�:_x�9�y�9��e9�V9K�$8"4S�y���<p�pɦ��2չ2���b��.���D���Z�J�o�kw��`Ō����������y뾺,�Ⱥ,Ӻ5Sݺ���k����������JD�;����e3��v#��(�d�-��3��A8��j=�֕B�)�G�:�L��AR��W���\��fb���g�om��s���x��)~��ځ�d����R��������E���ڑ��i�������~���  �  :�=�L=��=��=�S=��=�=^R=C� =�� =L =���<�9�<���<���<�0�<��<��<=,�<Y��<���<�&�<�w�<Z��<��<d`�<���< ��<�6�<�{�<Ͽ�<7�<OI�<i��<7��<� �<�k�<���<G�<T�<̡�<-��<�8�<}��<���<t�<�A�<�y�<���<��<K�<S/�<[R�<Xq�<f��< ��<��<e��<��<���<���<f��<���<��<O`�<F.�<5��<Ȩ�<�T�<���<}��<��<Z��<�<`��<8��<TL�<?��<C��<�N�<l��<K޼<w�<DV�<ш�<ô�<ڳ<���<��<Q$�<�1�<[:�<�>�<�?�<>�<�9�<34�<�,�<�$�<��<�<��<c��<0�<��<vӍ<X<!��<���<���<�g�<�K�<j]~<�!z<��u<�q<mtm<Ai<�e<��`<��\<�X<ύT<�wP<�cL<|QH<w?D<~,@<V<<U8<��3<��/<��+<ݝ'<ӄ#<�m<�Y<jI<�=<�7<E7<=<�I<ֹ�;���;�.�;�{�;;��;d:�;ī�;�)�; ��;�R�;��;�ɫ;G��;���;і;�;��;�4�;cz;�n;�lb;%W;7L;ϚA;OM7;�H-;,�#;�;t�;�;:��:���:�,�:���:I?�:��:�%�:׾�:�:kVh:\�M:
4:�:��:!�94�9-cf9�9��#8�U�9��&�q����j*ֹ�0�N���/�(�E�j[�u�p��Ԃ�����<���B���3���!������ɺ(Ӻ�Vݺ{��`�~���:�����#��r���T��J#��(�ͽ-�4�2��8�M=��|B���G�J�L��;R���W���\��qb���g�K�m��s�Էx��O~����(j��-�������[���|����������  �  M�=L=$�=c�=�S=��=d�=S=*� =� =sM =���<$=�<͎�<
��<�3�<I��<��<�.�<���<���<�'�<�x�<���<��<�_�<���<���<�4�<Hy�<��<�<�E�<׋�<���< �<Yh�<��<�<7Q�<@��<��<�6�<(�<��<�<B�<�z�<Ϯ�<���<B
�<�1�<-U�<rt�<���<P��<n��<���<��<���<A��<_��<2��<��<�`�<m.�<���<��<�S�<���<A��<9�<S��<��<�}�<t��<�H�<���<���<K�<��<Tۼ<��<T�<��<u��<Yٳ<���<��<�$�<�2�<�;�<�@�<ZB�<�@�<=�<a7�<E0�<(�<��<�<g
�<���<�<�<}ԍ<�<@��<9��<ڀ�<]f�<J�<�X~<vz<��u<M�q<,mm<�9i<Me<X�`<��\<��X<��T< rP<1_L<�MH<i<D<z*@<J<<A8<��3<l�/<��+<�'<��#<Os<�_<�O<�D<g><�=<�C<�O<#��;]��;;6�;؁�;C��;�<�;���;:(�;d��;BM�;z��;���;���;Ƞ�;�Ö;]�;q��;'�;��y;�m;fSb;�W;�#L;��A;T@7;?-;��#;�;��;!�;�:��:�L�:�"�:Jm�:�*�:hY�:��:���:C�h:D<N:_4:�:]7:���9�=�9�f9�9I#8�V��,��br��"����ֹߋ�xh��/�`F���[��-q�z��}R���n��"o���Z���A��,���$ɺ�1Ӻ�Yݺ���~��6m���y������l[�w������/#��l(��-���2��8� :=�$nB�W�G�t�L�
7R���W��\��xb�h�Ĕm��/s���x�g~�w���g���rx��a(���͌�Dj������Έ��=����  �  �=�K=��=Q�=�S=�=��=]S=� =H� =�M =���<?>�<��<i��<5�<b��<��<�/�<L��<I��<`(�<�x�<���<��<�_�<A��<��<Y4�<ox�<(��< �<�D�<���<=��<��<g�<��<��<?P�<W��<X��<m6�<�~�<���<�<B�<�z�</��<<��<�
�<�2�<V�<�u�<���<���<ȹ�<���<:��<���<���<��<ɧ�<d��<
a�<g.�<���<���<S�<\��<���<D�<S��<w�<h|�<(��<�F�<���<B��<�I�<딾<[ڼ<��<lS�<���<��<$ٳ<���<��<$%�<N3�<<�<�A�<C�<�A�<$>�<�8�<�1�<X)�< �<*�<M�<���<��<��<�ԍ<$Ë<D��<��<���<�e�<�I�<oW~<�z<��u<�q<�jm<57i<4e<��`<]�\<��X<v�T<ApP<�]L<|LH<_;D<�)@<�<<78<��3<��/<��+<آ'<�#<u<�a<AR<(G<:A<u@<F<�Q<���;���;9�;3��;r��;q=�;��;�'�;"��;}K�;X��;���;���;���;r��;�	�;�~�;!�;"�y;/�m;�Jb;uW;�L;M�A;d<7;�;-;(�#;\;��;b�;�
�:Y��:+X�: /�:d|�:�<�:^k�:]
�:|�:f�h:�`N:}4:':UM:X��9�W�9/�f9��9+$#8�WW�	f�^�r�M��[׹���^���0��EF�d\�]q�q ��~e��l����}���h��_K���3���*ɺ
4Ӻ_Zݺp��U��e���t���e��S����a��%#�xb(�;�-�*�2��8�4=��hB���G���L��5R���W��\��zb�h��m��5s��x��o~� ���Ä��}���.��Lӌ��n��6�������� ����  �  M�=L=$�=c�=�S=��=d�=S=*� =� =sM =���<$=�<͎�<
��<�3�<I��<��<�.�<���<���<�'�<�x�<���<��<�_�<���<���<�4�<Hy�<��<�<�E�<׋�<���< �<Yh�<��<�<7Q�<@��<��<�6�<(�<��<�<B�<�z�<Ϯ�<���<B
�<�1�<-U�<rt�<���<P��<n��<���<��<���<A��<_��<2��<��<�`�<m.�<���<��<�S�<���<A��<9�<S��<��<�}�<u��<�H�<���<���<K�<��<Tۼ<��<T�<��<u��<Yٳ<���<��<�$�<�2�<�;�<�@�<ZB�<�@�<=�<a7�<E0�<(�<��<�<g
�<���<�<�<}ԍ<�<@��<9��<ڀ�<]f�<J�<�X~<uz<��u<M�q<,mm<�9i<Me<X�`<��\<��X<��T< rP<1_L<�MH<j<D<{*@<J<<B8<��3<m�/<��+<�'<��#<Os<�_<�O<�D<g><�=<�C<�O<#��;]��;;6�;؁�;B��;�<�;���;9(�;c��;AM�;z��;���;���;Ƞ�;�Ö;]�;p��;'�;��y;�m;fSb;�W;�#L;��A;T@7;?-;��#;�;��;!�;�:��:�L�:�"�:Jm�:�*�:hY�:��:���:C�h:D<N:_4:�:]7:���9�=�9�f9�9I#8�V��,��br��"����ֹߋ�xh��/�`F���[��-q�z��}R���n��"o���Z���A��,���$ɺ�1Ӻ�Yݺ���~��6m���y������l[�w������/#��l(��-���2��8� :=�$nB�W�G�t�L�
7R���W��\��xb�h�Ĕm��/s���x�g~�w���g���rx��a(���͌�Dj������Έ��=����  �  :�=�L=��=��=�S=��=�=^R=C� =�� =L =���<�9�<���<���<�0�<��<��<=,�<Y��<���<�&�<�w�<Z��<��<d`�<���< ��<�6�<�{�<Ͽ�<7�<OI�<i��<7��<� �<�k�<���<G�<T�<̡�<-��<�8�<}��<���<t�<�A�<�y�<���<��<K�<S/�<[R�<Xq�<f��< ��<��<e��<��<���<���<f��<���<��<O`�<F.�<5��<Ȩ�<�T�<���<}��<��<Z��<�<`��<8��<TL�<?��<C��<�N�<m��<K޼<w�<DV�<ш�<ô�<ڳ<���<��<Q$�<�1�<[:�<�>�<�?�<>�<�9�<34�<�,�<�$�<��<�<��<c��<0�<��<vӍ<X< ��<���<���<�g�<�K�<j]~<�!z<��u<�q<mtm<Ai<�e<��`<��\<�X<ύT<�wP<�cL<|QH<x?D<~,@<V<<U8<��3<��/<��+<ݝ'<ӄ#<�m<�Y<jI<�=<�7<E7<=<�I<ֹ�;���;�.�;�{�;:��;c:�;ë�;�)�;���;�R�;��;�ɫ;F��;���;і;�;��;�4�;az;�n;�lb;%W; 7L;ϚA;NM7;�H-;,�#;�;s�;�;:��:���:�,�:���:I?�:��:�%�:׾�:�:kVh:\�M:
4:�:��:!�94�9-cf9�9��#8�U�9��&�q����j*ֹ�0�N���/�(�E�j[�u�p��Ԃ�����<���B���3���!������ɺ(Ӻ�Vݺ{��`�~���:�����#��r���T��J#��(�ͽ-�4�2��8�M=��|B���G�J�L��;R���W���\��qb���g�K�m��s�Էx��O~����(j��-�������[���|����������  �  ��=�M=W�=��=�S=`�=*�=6Q=�� =� =�I =��<�4�<��<.��<&+�<�~�<^��<(�<�|�<��<i$�<tv�<���<�<Ha�<F��<x��<:�<Z�<=��<	�<�N�<7��<)��<�&�<�q�<��<F�<�X�<ĥ�<���<e;�<U��<��<��<�A�<�x�<��<���<�<w+�<�M�<vl�<��<���<���<���<!��<T��<���<3��<0��<2��<h_�< .�<���<)��<�V�<���<��<�<E��<K�<"��<d��<�R�<���<i�<dT�<���< �<�!�<�Y�<���<���<]۳<w��<Z�<G#�<�/�<�7�<�;�<�;�<t9�<�4�<�.�<v'�<H�<p�<%�<;�<���<�<"��<�э<~��<���<,��<��<�i�<�N�<[d~<*z<r�u<E�q<�m<Mi<�e<��`<��\<`�X<��T<Q�P<KkL<�WH<�CD<�/@<�<<}8<V�3<��/<�+<��'<m}#<e<�O<�><�2<,<�+<d2<�?<[��;���;"�;Pr�;���;)7�;A��;D,�;<��;#[�;�;|׫;��;�;J�;^2�;;�K�;�9z;8n;��b;�HW;SUL;m�A;�a7;zV-;�#;�;��;��;)��:���:}��:���:���:���:Ν:Xf�:'j�:j�g:�7M:�p3:�>:u�:_x�9�y�9��e9�V9K�$8"4S�y���<p�pɦ��2չ2���b��.���D���Z�J�o�kw��`Ō����������y뾺,�Ⱥ,Ӻ5Sݺ���k����������JD�;����e3��v#��(�d�-��3��A8��j=�֕B�)�G�:�L��AR��W���\��fb���g�om��s���x��)~��ځ�d����R��������E���ڑ��i�������~���  �  ��=<O=J�=e�=�S=��=�=�O=�� =y� =G =���<�-�<�~�<��<$�<Jx�<��<�"�<x�<0��<�!�<�t�<���<�<Yb�<^��<d��<�=�<��<���<r�<~U�<s��<���<R.�<'y�<6��<��<�^�<��<���<�>�<̈́�<���<c�<&A�<�w�<y��<&��<� �<P&�<�G�<f�<,��<{��<���<#��<���<[��<ͽ�<��<˟�<˃�<^�<�-�<]��<ի�<�Y�<&��<���<r �<���<9�<���<��<�Z�<��<�<�[�<x��<<�<�&�<$^�<�<;��<�ܳ<���<��<�!�<V-�<-4�<7�<�6�<a3�<e.�<�'�<X �<3�<��<��<U��<��<��<�܏<fύ<��<���<ɚ�<���<Ql�<>R�<;m~<�4z<��u<��q<;�m<\i<7.e<�a<2�\<?�X<\�T<~�P<�tL<U_H<�ID<�3@<�<<?8<�3<Z�/<�+<��'<ws#<cY<�B<�0<�#<U<I<{$<�2<ڐ�;u��;I�;ae�;���;�1�;ѩ�;/�;7��;te�;=�;�;-Ѥ;Bם;���;N�;�ŉ;Ai�;^rz;�nn;��b;wW;�|L;�A;�z7;�h-;כ#;�;Q�;��;���:�p�:L��:3g�:j��:s?�:�^�:p�:%��:V�f:AeL:\�2:��:�� :���9�ӡ9�e9�9B%8igP��x���n������ӹY� �^��{�-�QD�ԶY��o�F��V��w���G�������Ǯ�����,�Ⱥ,Ӻ_QݺL�纞7����λ��	��o������hk��#���(��.�KJ3�Rp8�Ē=��B���G�^M�.LR���W���\�'Xb�P�g��Rm��r��kx�q�}�Ϳ���}���4��u㉻9���`(��[����P���ޖ�Ml���  �  ��=�P=7�=ɨ=gS=�=Υ=�M=P� =�� =�C =@��<�%�<�v�<r��<��<Fp�<���<�<kr�<���<�<1r�<���<�<Tc�<���<���<:B�<���<#��<��<t]�<��<o��<7�<с�<y��<{�<pe�<۰�<���<B�<���<��<��<j@�<�u�<���<��<���<) �<A�<L^�<x�<��<��<��<��<y��<���<���<ƛ�<��<8\�<-�<��<t��<�\�< �<���<�&�<���<-%�<:��<2�<�c�<���<�<Jd�<@��<�<�,�<c�<ʒ�<���<^޳<a��<�<��<I*�<0�<�1�<I0�<S,�<�&�<��<��<��<��<��<���<r�<��<�؏<�̍<T��<��<Z��<[��<9o�<$V�<�w~<�@z<�	v<n�q<�m<�mi<�?e<ra<S�\<?�X<��T<%�P<�L<�gH<6PD<�7@<�<<�8<(�3<N�/<�+<��'<�g#<�K<�3<? <�<�<�<�<^#<-u�;&��;k��;�U�;���; +�;��;f1�;@��;q�;,�;���;��;��;�;�n�;��;�;"�z;g�n;= c;��W;��L;#�A;ٖ7;�|-;��#;;�;؛;�w�:;-�:�Z�:y�:-%�:«:�ڜ:�i�:bm�:�e:iK:�1:��:�P :R��9��9id99��%8��M�g*�s�l������yҹ� ���.�,���B���X���m��z��bՋ����_9��P��Rg�������Ⱥ��Һ�Oݺ���%[���>��JA	������M]�Э���#��/)��_.���3�h�8���=���B�w�G��%M�zYR��W���\��Jb���g��2m���r�W;x�\�}�����[\��������Lg���������4��OƖ�W���  �  ��=ZR=$�=&�="S= �=S�=�K=�� =S� =@ =��<�<lm�<<��<��<�g�<׽�<��<Jl�<���<�<�o�<��<��<Qd�<���<!��<�F�<I��<���<[�<�e�<��<���<e@�<���<��<�!�<�l�<���<���<hF�<K��<���<?�<u?�<�s�<+��<~��<���<o�<9�<�U�<3o�<���<��<)��<���<��<���<"��<@��<�}�<;Z�<C,�<���< ��<�_�<N�<��<!-�<��<�-�<0��<�
�<�m�<���<��<2m�<���<q��<3�<%h�<і�<���<�߳<���<��<��<�&�<R+�<�+�<p)�<�$�<�<��<��<��<���<���<�<��<6ޑ<aԏ<`ɍ<R��<:��<ۛ�<���<)r�<3Z�<��~<�Mz<yv<��q<��m<D�i<�Re<;)a<>]<�X<�T<�P<֊L<�pH<�VD<�;@<R<<� 8<��3<w�/<��+<7{'<�Z#<�<<�"<A<��<��<B�
<�<�<�V�;��;j��;D�;��;%#�;i��;�3�;��;}�;H<�;��;7�;��;>�;	��;E�;خ�;��z;#�n;>c;�W;��L;- B;�7;��-;��#;Y;��;��;"?�: ��:���:q��:֩�::�:
K�:�֍:��:՞d:XJ:��0:�:r/�9�U�9*�9@�b9l9Ug&8�K�����j��T����й�V��"���+�&�A�WtW���l�Zꀺ0O��Õ���˟��󩺕���K��|�Ⱥ�Һ�Pݺp��|��A����Sq	�!��|B�C�����7>$�ix)�7�.���3���8���=��	C��!H��>M��hR���W���\��<b�^�g��m���r�`x�*�}�����9��9톻:���SB���㎻�����`����A���  �  ѧ=�S= �=`�=�R=*�=��=�I=�� =� =J< =���<:�<*d�<��<�	�<�^�<���<��<�e�<Z��< �<�l�<g��<O�<e�<���<J �<'K�<���<x��<�%�<n�<���<���<�I�<���<���<Z)�<�s�<��<��<.J�<���<���<?�<O>�</q�<���<���<(��<��<�1�<�M�<6f�<�{�<ҍ�<,��<>��<��<��<^��<���<z�<�W�<@+�<���<���<+b�<L�<4��<`3�<j��<�5�<3��<H�<aw�</��<(�<v�<���<���<29�<2m�<���<0��<8�<���<��<0�<#�<�&�<&�<c"�<��<��<��<g�<c��<���<l�<E�<��<�ؑ<�Ϗ<�ō<��<0��<��<|��<�t�<8^�<,�~<�Yz<�&v<��q<>�m<��i<�ee<�;a<]<��X<�T<��P<��L<vyH<]D<e?@<� <<��7<�3<�/<a�+<9p'<NM#<{-<<*�<��<j�<6�
<��<�<�7�;�|�;���;2�;���;��;i��;�4�;��;��;fL�;�&�;��;/,�;�]�;���;A.�;+҃;�@{;B2o;zc;�X;�M;)EB;�7;U�-;��#;�;ǣ;[u;��:ғ�:a��:$�:�*�:3��:��:�@�:�~:�zc:nHI:��/:x:���9��9\9�9��a9C]9J&8��H���Gi�
#��̅Ϲ������A�*��@��OV�F�k� \��8Ɋ����^`������Գ�����jȺ��Һ�Wݺ���>�������/��	�$������B?�Ɉ$���)���.�G4�(9�q,>��6C��DH�sYM�(yR��W�M�\��/b�Z�g�[�l��ar���w��L}�`�����Ɇ�bv��
�������^������
����,���  �  ��=U=��=}�=SR=3�=$�=vG=A� =�� =�8 =���<��<n[�<-��<� �<�V�<���<��<�_�<@��<�<�i�<ſ�<��<�e�<Y��<�<O�<Ù�<���<�,�<�u�<ݾ�<U�<&R�<?��<���<�0�<z�<w��<	�<vM�<��< ��<�</=�<�n�< ��<T��<y��<.�<`*�<�E�<�]�<s�<(��<���</��<ǣ�<���<���<#��<�v�<�U�<B*�<���<��<�d�<��<٧�<19�<+��<R=�<���<��<j��<3��<�0�<G~�<ž<D�<�>�<�q�<靷<võ<I�<���<��<��<��<�!�<D �<��<9�<k�<��<���<���<?�<r�<��<�ٓ<�ґ<vˏ<�<뷋<&��<��<���<"w�<�a�<]�~<dez< 4v<�r<u�m<��i<�ve<�La<�%]<� Y<��T<��P<��L<�H<QbD<�B@<6!<<+�7<Z�3<�/<�+<me'<�@#<+<<��<�<f�<5�
<V�<z�<�;Bc�;κ�;� �;(��;��;F��;=5�;g��;x��;zZ�;y9�;�1�;�E�;�z�;Ґ;�N�;&�;��{;hoo;�c;�GX;0M;fB;_�7;�-;��#;�;=�;�`;���:5I�:B�:���:o��:�/�:/�:���:in}:�eb:�AH:��.:[<:�<�9Y��92T�9�_`9��9�q%8��F�f����g�r��|+ι������)���?��=U�B�j�9���M���������H�����_轺MȺ�Һ�_ݺ��=��~���NW���	��K�0��6)������$��*�J1/��J4�EX9�j^>�nbC�gH��sM�։R�S�W���\�E%b�^wg� �l��<r�ݨw��}��B����������T��i���J����@���ޓ��{������  �  '�=V=M =��=�Q=9�=��=�E=�� =8� =�5 =#��<��<�S�<���<q��<wO�<J��<� �<�Z�<Դ�<��<g�<
��<�<�e�<���<^�<PR�<���<���<�2�<'|�<���<o�<OY�<<��<+��<�6�<}�<��<��<4P�<���<���<��<�;�<�l�<��<O��<���<t�<�#�<�>�<}V�<�k�<�}�<q��<@��<]��<���<���<'��<�s�<�S�<)�<���<ز�<�f�<��<ȫ�<>�<���<�C�<~��<T$�<���<���<�7�<,��<`˾<�
�<�C�<mu�<���<Cŵ<�<X��<\�<u�<q�<��<B�<��<��<h�<���<��<+�<�<�ߗ<�ٕ<ԓ<(Α<�Ǐ<���<ĵ�<��<���<���<y�<�d�<�~<�nz<\?v<hr<��m<��i<k�e<#[a<B3]<�Y<i�T<��P<ۧL<s�H<�fD<$E@<�!<<��7<��3<_�/<��+<+\'<�5#<c<�<6�<��<��<��
<��<y�<N�;�L�;���;\�;O��;9
�;P��;F5�;^��;d��;$f�;�H�;�D�;;\�;<��;'�;$j�;��;X�{;'�o;|�c;IqX;�RM;�B;��7;|�-;A�#;�	;�;�M;���:��:B��:=^�:�J�:���:���:�9�:Nz|:�za:`G:<.:N�:��9��9%��9�4_9-9f�$8��E����8f��+��4͹h���+�)��>��XT�}�i���~�)扺RO��뫞�e��&^�������5Ⱥ��ҺhݺN)�g����z�.�	�|�N��b�����%��D*�k/���4�"�9��>��C���H���M�A�R�g�W�(�\�(b�\gg���l�Kr���w��|��)���ۃ�a���n7��#���]����'��ȓ�+h���	���  �  I�=�V=� =��=�Q=|�=��=D=)� =� ==3 =���<���<N�<���<���<�I�<=��<���<�V�<]��<��<e�<���<v�<f�<���<�<�T�<��<R��<�6�<��<
��<��<�^�<���<7��<T;�<���<w��<��<3R�<��<9��<��<�:�<�j�<���<��<���<��<�<G9�<�P�<�e�<�w�<���<��<���<x��<&��<���<Eq�<�Q�<'(�<w��<h��<�g�<��<���<�A�<��<�H�<Ƚ�<*�<ʍ�<���<�=�<a��<!о<��<G�<;x�<���<qƵ<��<��<N
�<��<��<r�<c�<k�<�	�<� �<���<"�<=�<8��<Dڗ<�ԕ<�ϓ<pʑ<_ď</��<&��<!��<Л�<-��<kz�<�f�<�~<vz<�Gv<�r<e�m<�i<��e<\fa<�=]<�Y<�T<"�P<�L<8�H<jD<�F@<�!<<3�7<��3<�/<�~+<�T'<	-#<�<��<{�<��<=�<��
<��<��<w��;N;�;Θ�;��;L~�;��;֕�;�4�;���;���;�n�;�T�;�R�;�l�;���;� �;I�;�#�;��{;��o; d;�X;�lM;ԖB;O8;��-;��#;�;��;�?;l�:���:մ�::�:v��:h�:�[�:jً:�{:��`:��F:�u-:��:��9J�9���9�S^9�z9�($8��D�S��De�񀟹�6̹y����r�ia(��>���S��i�k*~�����U��tn��Ш�6��¥��q'Ⱥ��ҺDpݺ�=躎#�5 ��E��T
����j��������;%�/t*�S�/���4���9��>�"�C�z�H�ٜM���R� �W��\��b�2\g�^�l��r�=fw���|����!ǃ�[u��[!��ʋ�mp�����9����Y�������  �  ��=KW=� =��=BQ=��=�=(C= � =�� =�1 =���<I��<~J�<���<���<>F�<��<���<�S�<&��<�	�<�c�<Ի�<�<)f�<��<
�<;V�<���<���<�9�<��<B��<A�<*b�<��<b��<@>�<!��<���<0�<rS�<���<���<w�<K:�<�i�<���<��<j��<%��<��<�5�<)M�<b�<-t�<��<i��<^��<���<���< ��<�o�<�P�<�'�<T��<ӳ�<�h�<>�<w��<�C�<���<�K�<��<�-�<T��<��<A�<���<&Ӿ<��<&I�<�y�<���<Gǵ<��<���<�	�<��<>�<e�<��<��<��<f��<T��<��<��<�ܙ<�֗<�ѕ<�̓<ȑ<j<���<��<���<���<���<>{�<h�<^�~<�zz<Mv<�r<��m<x�i<c�e<ma<xD]<�Y<��T<��P<αL<$�H<�kD<�G@<�!<<J�7<��3<�/<�z+<CP'<�'#<�<��<#�<;�<�<S�
<]�<��<���;:0�;G��;��;x�;���;���;_4�;\��;`��;!t�;r[�;�[�;Ow�;{��;��;���;�0�;Y�{;G�o;gd;��X;�|M;�B;s8;x�-;��#;�;";�5;nQ�:v��:���:���:Hȸ:`/�:8"�:E��:�F{:�K`: @F:�-:�:nd�9@��9w�9��]9�!9��#8�?D�+�
�M�d�w����˹���{���'�W�=��=S��h���}�f��#ۓ�uG��򰨺���l����Ⱥ��Һ�uݺ�J�(9�0<������0
�����7�(��A �aX%���*��/�'�4�F�9���>��C�­H�+�M��R�q�W���\�b�`Ug���l��q�PTw�f�|��
��Z���\h���������c��^��Y����P��r����  �  �=�Q=��=7�=�J=��=(�=�==h� =ڈ =]. =���<���<cD�<���<��<;�<���<���<>�<&��<���<�A�<u��<b��<�:�<��<���<6$�<o�<��<��<>J�<��<}��<� �</g�<A��<<��<B6�<�x�<F��<v��<�2�<�j�<^��<(��<���<�%�<�J�<�k�<n��<���<ú�<���<���<��<��<���<y��<���<O��<���<Ϳ�<��<�n�<+7�<b��<��<R�<���<��<��<Ɛ�<	�<ax�<���<�>�<���<.�<�0�<@s�</��<��<J�<�;�<�]�<�y�<��<Ǡ�<���<:��<^��<���<���<\��<B��<˯�<���<���<���<b��<̡�<���<���<���<��<���<�|�<up�<ob�<S�<*�~<|`z</;v<kr<��m<o�i<7�e<%�a<�a]<�AY<#U<�Q<3�L<!�H<��D<�@<�v<<=X8<?94<�0<��+<��'<��#<��<Ŗ<ĉ<��<x�<7�<��<��<���;P#�;���;��;���;�!�; ��;Vu�;$6�;m�;��;�;m��;)-�; z�;~�;ut�;U&�;���;'�u;5j;��^;)�S;��H;i2>;��3;��);	 ;|z;�';f;'m�:�2�:�t�:X2�:�o�:-�:�f�:x�:��t:*�Y:�?:�X&:�:�y�9R��9]�9�99��8C�ܴ<)��mE8��̉��:���f�V������4���J� �`�o5v��х�|����'���9N����i�ź�Wкm&ۺr��������
	�T��h�=r�o��S,$��p)���.���3���8�$�=��C�$#H�9M�0VR��}W�)�\��a�8g��l�S�q�$Ew�1�|����淃��h��o���ċ��o��I��ē��m������  �  ��=�Q=��=4�=�J=��=_�=9>=�� =+� =�. =q��<���<iE�<ԕ�<��<�;�<K��<���<�>�<̕�<~��<7B�<���<}��<�:�<��<���<�#�<�n�<N��<,�<qI�<=��<���<��<Rf�<`��<���<�5�<4x�<Ǹ�<��<�2�<�j�<f��<I��<7��<-&�<'K�<il�<��<p��<���<���<���<��<���<u��<@��<L��<���<+��<@��<Q��<�n�<17�<E��<���<�Q�<��<~��<�<��<�<ww�<���<�=�<���<H�<�/�<�r�<���<�<��<�;�<�]�<�y�<3��<��<$��<Ҵ�<���<.��<f��<��<1��<߰�<���<���<ħ�<)��<n��<F��<J��<��<`��<ᆉ<�|�<Yp�<Lb�<�R�<+�~<N_z<�9v<	r<�m<��i<p�e<t�a<`]<8@Y<�!U<�Q<"�L<7�H<H�D<Г@<v<<qX8<�94<�0<��+<<�'<��#<?�<_�<i�<ǅ<��<;�<6�<X�<���;�%�;l��;��;\��;�"�;���;ju�;�5�;��;��;.�;��;�*�;w�;:�;Pq�;�"�;_��;d�u;0j;��^;�S;+�H;�/>;��3;��);�	 ;�{;i*;;;w�:�=�:�~�:?�:�|�:F;�:�w�:�-�:��t:�Y:t�?:�m&:&�:u��9���9�r�9�+99�(�8��*E��p8�쉹	]�����m��*��K5��K�R�`�Qv�!߅������#������?V��������ź�Xк�$ۺ��2��U���{���ڀ� ��l�����#$��h)�!�.�Q�3�j�8�$�=�C��H�n5M�TR��|W�>�\���a�>9g�t�l�W�q��Iw��|�r	��Y���l�����ȋ�5s��,���Ɠ�#p������  �  .�=/Q=��=7�=(K=V�=�=�>=�� =+� =�/ =���<<��<H�<{��<���<�>�<ɓ�<���<�@�<v��<���<,C�<@��<���<�:�<���<���<�"�<m�<q��<��<"G�<ˎ�<(��<)�<�c�<��<h��<�3�<�v�<���<��<�1�<�j�<���<���<��<K'�<�L�<>n�<'��<Ѧ�<��<K��<:��<���<���< �<� �<e��<���<���<[��<��<:o�<U7�<���<��<�P�<���<���<��<ȍ�<��<�t�<���<J;�<$��<��<�-�<�p�<���<��<�<�:�<w]�<�y�<���<�<E��<^��<Ӻ�<W��<ӻ�<���<޶�<���<S��<0��<Q��<���<{��<��<���<1��<"��<Y��<�|�<�o�<�a�<�Q�<��~<�[z<�5v<�r<#�m<��i<<�e<f|a<[]<�;Y<�U<� Q<T�L<��H<ƮD<ޒ@<yv<<,Y8<;4<�0<u�+<��'<	�#<�<��<א<R�<2�<З<��<��<N��;<.�;���;o�;���;�%�;g��;�u�;|4�;(�;��;��;��;�"�;In�;�ٓ;�g�; �;��;��u;pj;��^;[�S;��H;o(>;��3;5�);� ;�;`1;�;O��:�[�:5��:�e�:%��:[f�:Ţ�:�X�:�u::.Z:@:ղ&:A�:��9"�9���9`l99�d�8�l�۹���8�j;���ķ�	�	���K��f5�ASK��a�
�v�Y�����:B���ԥ�i�����2�ź8[к� ۺ���������n����o�Y��W�C��\$��R)�Љ.���3���8���=��B��H�-M�CNR�&yW���\��a��>g���l���q��Ww�S�|�a��8Ń� v��4%���ы�}��5&���Γ�Ww��� ���  �  L�=�P=3�=0�=eK=��=��=�?=�� =ċ =�1 =ӯ�<s��<jL�<��<��<�B�<���<g��<�C�<��<���<�D�<?��<(��<^:�<���<���<� �<�j�<���<���<C�<܊�<	��<�<�_�</��<���<�0�<�s�<`��<���<�0�<j�<���<x��<I��<)�<�N�<q�<���<a��<��<���<���<��<���<�</�<���<���<���< ��<N��<�o�<X7�<h��<ݦ�<�N�<x��<��<�	�<��<��<�p�<���<�6�<��<�߿<�)�<\m�<0��<��<e�<�9�<
]�<z�<h��<9��<$��<���<���<���<s��<½�<��<㷝<���<m��<>��<��<ȧ�<ѣ�<���<���<X��<���<�|�<to�<x`�<�O�<|~<LVz<�/v<br<n�m<t�i<іe<ta<3S]<F4Y<�U<&�P<u�L<E�H<�D<t�@<=v<<Z8<-=4<�0<�,<�'<��#<�<e�<x�<-�<E�<��<V�<j�<��;Q;�;���;��;���;T*�;���;�u�;2�;l �;�;�ٮ;H�;e�;y`�;�ʓ;�W�;9	�;t��;�u;�j;3�^;'|S;��H;�>;��3;��);( ;u�;3<;�-;ӵ�:���:���:��:�:���::�:��:��u:��Z:��@:�':;:���9���9��9k�99W��8�=E��ߺ���9��hl��b�幡k	����G�5���K�K�a��w��>���ݐ�Gq��?���0������G�ź�^к�ۺ���'�𺁻��Z����\S����'6�$��4�#�X0)��g.���3�g�8���=�`�B��H�bM�ER��tW���\���a�NHg�l�l�+r��mw���|�� ��|ԃ�O����5��Y⋻v����4���ۓ�����Y*���  �  "�=�O=��=�=�K=��=��=eA=�� =ɍ =�3 =��<��<�Q�<���<���<H�<���<���<�G�<H��<x��<�F�<p��<���<:�<���<���<;�<ig�<���<^��<�>�<���<���<��<�Z�<0��<C��<�,�<fp�<���<t��</�<yi�<���<Q��<� �<c+�<�Q�<�t�<���< ��<H��<���<��<���<!�<2	�<��<��<��<���<^��<˟�<�p�<K7�<���<b��<�L�<w��<>|�<c�<7��<S��<k�<���<I1�<e��<�ڿ<3%�<0i�<���<�ݸ<<�<s8�<p\�<*z�<L��<ͤ�<���<ɻ�<`��<ĥ<Kģ<�¡<��<���<,��<Ͷ�<j��<Я�<�<X��<�<#��<ڒ�<���<�|�<�n�<�^�<�M�<v~<Oz<'v<��q<7�m<��i<
�e<>ia<�H]<}*Y<3U<��P<�L<g�H<��D<��@<�u<<[8<�?4<�#0<�,<��'<��#<��<̯<q�<��<�<�<j�<��<��;�K�;���;O"�;,��;00�;W��;�u�;6/�;I��;;ٵ;�ͮ;ܧ;��;N�;��;�C�;��;̀;��u;�i;&{^;�aS;^�H;}>;�3;	�);� ;E�;�I;�@;5��:���:K�:P��:�;�::�:�C�:��::=v:Z[:$-A:(�':2�:e�9��9i�9�L:9��8�c��� ����:��n��fF����湧�	��a �M�6���L�0=b���w�G����%������1��1����6��W�źYdк�ۺ��庍�𺍒��[@� ���/�#����wk���#�)��<.��j3��8��=���B���G�yM��9R�2oW�L�\���a��Tg�T�l�r���w�_�|��3���胻����K������ࠎ��G���쓻/����6���  �  ��=�N=5�=��=L=M�=�=�B=�� =� =�6 =���<	�<iX�<��<���<%N�<?��<��<$L�<��<o��<�H�<���<��<�9�<h��<���<7�<�c�<3��<;��<�8�<��<^��<W�<]T�<R��<���<�'�<Kl�<-��<���<�-�<�h�<П�<5��<��<�-�<aU�<�x�<���<���<.��<1��<���<�<q
�<�<f�<��<D��<J��<���<~��<uq�<F7�<���<���<�I�<���<�w�<M �<��<*��<�d�<5��<�*�<��<�Կ<��<2d�<l��<;ڸ<��<�6�<�[�<Ez�<5��<���<*��<J��<�ŧ<�ȥ<�ɣ<�ȡ<�Ɵ<ĝ<���<��<K��<:��<���<|��<B��<���<���<���<�|�<�m�<!]�<�J�<o~<�Fz< v<��q<.�m<�i<!e<|\a<�<]<Y<�U<��P<��L<l�H<_�D<�@<u<<>\8<�B4<�(0<�,<��'<�#<G�<��<:�<լ<r�<_�<4�<��<^ <_�;2��;n/�;)��;�6�;���;u�;)+�;��;dε;&��;˧;M�;a8�;ܟ�;-+�;e܆;i��;�hu;�i;OV^;�BS;zH;N�=;Կ3;L�);� ;��;�X;�V;� �:�	�:9l�:�F�:���:�h�:d��:�b�:�
w:o\:��A:�H(:M;:�F�9�ʼ9�9��:9��8�q��T���]�;��?��>F�����"�
��!�]T7��MM�	c���x��膺�x������n���ⰺ>[���ź�mк�ۺ���3��d���"����Q��t���
8���#��(��
.��;3��d8�-�=��B���G��L��,R�`iW�E�\�b��cg�u�l�%:r���w�!}��I��� �������d�����与��]��� �������D���  �  "�=�M=��=Ȣ=FL=	�=�=�D=�� =�� =j9 =���<��<N_�<��<��<�T�<K��<���<�P�<��<~��<�J�<���<^��<�8�<��<��<��<|_�<A��<���<�2�<y�<���<��<�M�<��<���<e"�<�g�<r��<��<�+�<�g�<���<��<j�<�0�<�X�<:}�<���<d��<e��<���<l��<��<!�<Q�<-�<��<���<���<���<8��<$r�<7�<x��<u��<�F�<���<*s�<���<Zy�<`��<�]�<��<`#�<�{�<�Ϳ<��<�^�<ȝ�<eָ<��<�4�<{Z�<5z�<	��<���<緫<�©<'ʧ<-Υ<�ϣ<Pϡ<�͟<�ʝ<�Ǜ<�Ù<~��<�<Ƶ�<ί�<���<G��<-��<8��<d|�<�l�<[�<�G�<Rg~<(=z<=v<��q<�m<��i<Cqe<�Na<M/]<�Y<��T<��P<c�L<ܴH<ǟD<>�@<t<<]8<zE4<c-0<J,<L�'<�#<��<&�<��<�<��<��<��<��<� <xs�;G��;=�;���;�<�;A��;�s�;{&�;~�;+µ;���;���;�ܠ;} �;ц�;L�;*;Ӛ�;7u;��i;�-^;A S;�]H;�=;Z�3;a�);L ;M�;�h;Zm;�Z�:JR�:���:��:� �:�զ:��:"҉:��w:��\:R�B:��(:K�:X0�9O�9�]�9�A;9��8L�𵳂���E=��'���a��OJ鹾c���!��(8��'N���c�Zy�N��Eԑ�pI�������������ź�yк�ۺ*���k��4���p�9���D����T�ER#�Θ(���-�m
3��78�Sa=�,�B���G���L�R R��dW���\��b�Ytg���l�gYr���w�pL}��a�����Eφ�����+���Ҏ�rv�����ҵ���T���  �  ��=rL=��=��=�L=��=:�=/F=�� =�� =/< =��<'�<f�<ٶ�<��<[�<T��<��<�U�<��<��<�L�<!��<���<S8�<C��<���<s�<3[�<=��<���<�,�<gr�<���<���<�F�<z��<���<�<c�<���<��<�)�<xf�<���<���<
�<73�<a\�<���<���<��<���<h��<$�<��<��<��<��<��<��<3��<��<¤�<�r�<�6�<D��<4��<�C�<���<?n�<#��<s�<���<WV�<���<�<�t�<=ǿ<W�<PY�<��<�Ҹ<��<�2�<cY�<z�<ה�<.��<���<wƩ<�Χ<Vӥ<�գ<�ա<9ԟ<�ѝ<DΛ<Iʙ<�ŗ<���<���<��<��<���<���<劉<|�<fk�<�X�<�D�<__~<�3z<5v<[�q<��m<��i<6ce<�@a<�!]<Y<2�T<��P<��L<0�H<��D<2�@<�r<<�]8<H4<�10<�,<l(<��#<��<��<�<��<��<t�<4�<+�<M <\��;��;dJ�;��;C�;���;�r�;D!�;t�;뵵;ڠ�;���;BǠ;��;Sm�;���;���;���;�u;�\i;^;��R;qAH;8�=;(�3;T�); ;�;�v;�;Ĕ�:֘�:�:��:�g�:�?�:2��:�?�:��x:n�]:�XC:��):�Z:	�9,�9�͍9�;9�ݸ8\v��z���>����7�����&!��"��9��O��d��0z������0��Қ��N����Q��D����ƺޅк�
ۺ���4M�������K����	��s����#��b(�U�-���2��
8�:=�-iB�b�G��L��R��_W�۶\�-b���g���l�byr���w�ox}�z���4���ꆻ����!G��*펻鎑�-��Sɖ�ae���  �  ��=KK="�=>�=�L=O�=@�=�G=�� =/� =�> =���<-�<Ql�<7��<��<a�<ʳ�<��<�Y�<\��<7��<�N�<&��<���<�7�<���<��<,�<W�<}��<u��<�&�<l�<5��<��<u@�<h��<X��<�<�^�<��<<��<�'�<Ve�<+��<l��<~�<�5�<~_�<\��<T��<M��<h��<t��<w�<�<��<R!�<�<�<��<G��<O��<#��<^s�<G6�<���<��<�@�<��<�i�<���<$m�<J��<�O�<յ�<2�<$n�<���<~�<"T�<x��<�θ<��<�0�<;X�<�y�<���<���<���<�ɩ<�ҧ<إ<�ڣ<wۡ<Wڟ<؝<�ԛ<ZЙ<q˗<�ŕ<O��<˷�<'��<<��<c��<�{�<#j�<�V�<�A�<�W~<{*z<��u<��q<��m<�{i<Ve<�3a<A]<K�X<t�T<6�P<��L<��H<ܕD<�@<�q<<]^8<[J4<�50<�!,<�(<��#<7�<,�<m�<��< �<W�<��<�	<�' <���;4��;�V�;���;`H�;/��;�p�;�;�ؼ;��;���;ٓ�;���;��;(U�;�݌;���;�g�;/�t;T1i;��];0�R;�%H;�=;K�3;��);x ;�;|�;��;���:K��:^�:6W�:�Ķ:R��:�:o��:�~y:�m^:^D:�.*:��:7��9=ɾ9(2�9+<9!��8q�7�6hø`@�����~���!�����?t#���9���O��e���z�c�������眺R<������׻�F.ƺ}�к2ۺ��41�i������Z*�Њ�����D������"�I0(��p-�I�2���7�=�wKB���G���L�p
R�}\W���\��#b���g��m�)�r�Ox���}� ���9M���������a��������B���ۖ�$u���  �  ��=NJ=z�=��=�L=��=�=�H=� =� =�@ =i��<L!�<�q�<���<�<f�<���<�<_]�<M��<h �<UP�<מ�<���<�6�<,��<���<9�<�S�<U��<���<u!�<�f�<���<f��<;�<��<l��<��<�Z�<Ѡ�<���<&�<@d�<��<���<��<p7�<b�<���<3��<���<J��<���<��<B�<�"�<1&�<�#�<Z�<
�<���<&��<1��<�s�<�5�<���<��<>�<���<�e�<:��<�g�<���<�I�<گ�<K�<nh�<j��<m�<�O�<���<�˸<K �<�.�<(W�<py�<㕯<ᬭ<澫<^̩<�է<ܥ<eߣ<f�<�ߟ<Gݝ<�ٛ<�ՙ<MЗ</ʕ< Ó<��<���<æ�<��<���<D{�<�h�<�T�<B?�<(Q~<�"z<��u<��q<Ùm<{pi<vJe<�(a<Y
]<��X<�T<��P<ɲL<��H<��D<P�@<Np<<�^8<L4<!90<9&,<�(<C$<�<��<��<��<��<d�<�<�<�0 <ب�;��;d`�;���;<L�;u��;�n�;>�;@Ѽ;F��;���;9��;堠;�ޙ;�@�;�Ȍ;�x�;�R�;v�t;�i;¼];z�R;�H;G�=;|�3;�);c ; �;A�;��;���:l�:���:[��:&�:���:�E�:���:I(z:�_:#�D:�*:8F:z��9�H�9B��9_R<9�q�8�QW�aŸ�EA�����h���[�칍o��$�q|:�$�P��Af�S�{��c���Ԓ�z+��hu���������Fƺ��к�ۺ�庼𺣺��ȳ�J��i������p�?�"��(��G-���2�Ծ7���<�2B�6pG�شL��R��ZW�}�\��-b���g�W*m���r��<x�"�}�����b�����p̉�	w��t��G����T���떻�����  �  ��=�I=��=��=�L=�=��=�I=D� =q� =}B =��<+%�<�u�<���<#�<�i�<��<#�<`�<���<�<�Q�<c��<���<:6�<�~�<*��<��<�P�<
��<6��<��<zb�<Q��<��<�6�<�<���<'�<�W�<V��<���<�$�<Wc�<���<��<�	�<�8�<d�<.��<#��<'��<���<���<��<]�<�&�<�)�<�&�<G�<��<���<���<��<�s�<�5�<���<���<�;�<��<�b�<���<d�<j��<ZE�<:��<�
�<�c�</��<��<L�<���<�ȸ<H��<\-�<IV�<.y�<1��<ح�<[��<jΩ<pا<ߥ<��<�<��<f�<�ݛ<oٙ<�ӗ<�͕<
Ɠ<���<���<-��<<勉<�z�<�g�<WS�<+=�<	L~<mz<��u<�q<V�m<�gi<�Ae<�a<�]<�X<��T<y�P<Z�L<m�H<T�D<	@<Ko<<�^8<NM4<�;0<�),<�(<�$<��<T�<��<-�<��<��<	<�<<7 <���;��;�g�;P��;FO�;C��;gm�;P�;˼;���;qz�;�w�;|��;�ϙ;T0�;׷�;�g�;�B�;�t;=�h;S�];ԧR;��G;f�=;�|3;��);  ;�;G�;�;p�:H8�:���:t��:�O�:S7�:f��:�>�:��z:�_:�E:f+:ϙ:��9M��9ӿ�9�}<9�C�8"�q�kpƸ�9B��Z���B�����!��G�$��;�}Q��f�R0|��������a��֡��!ݱ�����Zƺ@�к�ۺg�庺�����]�����CQ�w������O��"���'�R(-��g2�o�7���<�{B�?aG���L���Q�kYW���\��5b��g�E;m�(�r��Ux�#�}�7���Ds���+��މ�>���D,���ɑ��b��n�������  �  ܛ=�H=��=��=�L=N�=�=BJ=�� =[� =�C =G��<�'�<;x�<=��<��<Zl�<C��<)�<�a�<۲�<�<+R�<���<���<�5�<>~�<��<�
�<O�<���<���<��<�_�<���<W��<
4�<d|�<G��<��<V�<���<���<�#�<�b�<_��<:��<
�<�9�<;e�<���<��<?��<D��<�<U�<� �<J)�<.,�<)�<1�<�<���<]��<���<�s�<>5�<0��<���<�:�<k��<�`�<M��<�a�<���<�B�<i��<��<a�<w��<�<�I�<���<aǸ<
��<p,�<�U�<�x�<c��<[��<B��<�ϩ<ڧ<��<��<��<�<��<}��<�ۙ<@֗<�ϕ<�Ǔ<���<���<���<p��<���<�z�<dg�<dR�<�;�<�H~<�z<)�u<�q<�m<\bi<,<e<Ja<f�\<��X<�T<c�P<թL<H<6�D<�}@<vn<<�^8<)N4<=0< ,,<�(<�$<��<��<��<J�<��<��<.
<�<�; <���;��;�l�;k��;<Q�;Q��;!l�;��;_Ǽ;���;�s�; p�;���;	ƙ;&�;w��;�]�;!8�;�zt;U�h;h�];-�R;��G;U�=;\v3;�);� ;ߴ;�;��;A(�:�Q�:��:���:�u�:�^�:��:�g�:	�z:��_:_HE:}M+:1�:�e�9f�9$�9�<9�8����!OǸv�B�G���G���>S��1�B�$�Z;��kQ�&#g���|��̈��3��g���󾧺0���^)��zgƺ�к|ۺ�}�������.��a��0A�������<���"���'��-�EU2��7�'�<�=B�LXG��L���Q��XW�D�\��:b�ۻg�JEm���r�2ex�>�}�7����}��6���艻	����6���ӑ��k��a ��쓙��  �  ��=�H=�=��=�L=^�=0�={J=5� =�� =�C =��<{(�<y�<��<w�<8m�<��<��<ib�<Z��<��<NR�<۟�<���<�5�<�}�<���<�	�<fN�<`��<��<0�<�^�<���<D��<3�<�{�<~��<D�<jU�<��<
��<S#�<�b�<J��<G��< 
�<�9�<�e�<=��<���<���<��<��<'�<�!�<%*�<-�<�)�<��<��<n��<���<���<t�<%5�<��<9��<:�<���<�_�<���<�`�<���<�A�<K��<��<2`�<���<?�<I�<抺<�Ƹ<���<,�<�U�<�x�<s��<s��<���<Щ<�ڧ<��<��<a�<��<��<Q�<�ܙ<ח<=Е<�ȓ<}��<4��<.��<���<	��<�z�<1g�<�Q�<l;�<bG~<Iz<��u<��q<t�m<^`i<�9e<<a<��\<\�X<��T<�P<w�L<��H<U�D<}@<7n<<�^8<dN4<{=0<�,,<�(<�$< <z�<��<��<��<��<�<!<�< <u��;��;Xn�;&��;�Q�;���;�k�;��;�ż;ҏ�;Lq�;�m�;���;
Ù;�"�;r��;fY�;�4�;�tt;M�h;:�];d�R;��G;��=;�s3;ϟ); ;m�;ߚ;0�;~0�:KZ�:���:R�:p��:�l�:y��:u�:�{:��_:r]E:a+:��:���9d��9��9��<9/��8A4����ǸC��䐹9俹~�K��
%��w;�׍Q��Dg�T�|�Cو�5@��l����ɧ������0��dlƺ��к�ۺ�{����ފ��;�����R<�������(5�y�"�&�'��-�O2�؎7�%�<�B�~TG�L�L��Q��XW�%�\�o<b��g�fIm���r�'jx���}�\���ꀄ�r:��퉻���:���֑��n����������  �  ܛ=�H=��=��=�L=N�=�=BJ=�� =[� =�C =G��<�'�<;x�<=��<��<Zl�<C��<)�<�a�<۲�<�<+R�<���<���<�5�<>~�<��<�
�<O�<���<���<��<�_�<���<W��<
4�<d|�<G��<��<V�<���<���<�#�<�b�<_��<:��<
�<�9�<;e�<���<��<?��<D��<�<U�<� �<J)�<.,�<)�<1�<�<���<]��<���<�s�<>5�<1��<���<�:�<k��<�`�<M��<�a�<���<�B�<i��<��<a�<w��<�<�I�<���<aǸ<
��<p,�<�U�<�x�<c��<[��<B��<�ϩ<ڧ<��<��<��<�<��<}��<�ۙ<@֗<�ϕ<�Ǔ<���<���<���<p��<���<�z�<dg�<dR�<�;�<�H~<�z<)�u<�q<�m<\bi<,<e<Ja<g�\<��X<�T<c�P<թL<H<6�D<�}@<vn<<�^8<)N4<=0< ,,<�(<�$<��<��<��<J�<��<��<-
<�<�; <���;��;�l�;k��;<Q�;Q��;!l�;��;_Ǽ;���;�s�; p�;���;	ƙ;&�;w��;�]�; 8�;�zt;U�h;g�];-�R;��G;U�=;\v3;�);� ;ߴ;�;��;A(�:�Q�:��:���:�u�:�^�:��:�g�:	�z:��_:_HE:}M+:1�:�e�9f�9$�9�<9�8����!OǸv�B�G���G���>S��1�B�$�Z;��kQ�&#g���|��̈��3��g���󾧺0���^)��zgƺ�к|ۺ�}�������.��a��0A�������<���"���'��-�EU2��7�'�<�=B�LXG��L���Q��XW�D�\��:b�ۻg�JEm���r�2ex�>�}�7����}��6���艻	����6���ӑ��k��a ��쓙��  �  ��=�I=��=��=�L=�=��=�I=D� =q� =}B =��<+%�<�u�<���<#�<�i�<��<#�<`�<���<�<�Q�<c��<���<:6�<�~�<*��<��<�P�<
��<6��<��<zb�<Q��<��<�6�<�<���<'�<�W�<V��<���<�$�<Wc�<���<��<�	�<�8�<d�<.��<#��<'��<���<���<��<]�<�&�<�)�<�&�<G�<��<���<���<��<�s�<�5�<���<���<�;�<��<�b�<���<d�<j��<ZE�<:��<�
�<�c�</��<��<L�<���<�ȸ<H��<]-�<IV�</y�<1��<ح�<[��<jΩ<pا<ߥ<��<�<��<f�<�ݛ<oٙ<�ӗ<�͕<
Ɠ<���<���<-��<<勉<�z�<�g�<WS�<*=�<	L~<mz<��u<�q<V�m<�gi<�Ae<�a<�]<�X<��T<y�P<Z�L<m�H<T�D<	@<Ko<<�^8<NM4<�;0<�),<�(<�$<��<T�<��<-�<��<��<	<�<<7 <���;��;�g�;O��;FO�;C��;fm�;O�;˼;���;qz�;�w�;|��;�ϙ;S0�;׷�;�g�;�B�;�t;<�h;R�];ӧR;��G;e�=;�|3;��);  ;�;G�;�;p�:H8�:���:t��:�O�:S7�:f��:�>�:��z:�_:�E:f+:ϙ:��9M��9ӿ�9�}<9�C�8"�q�kpƸ�9B��Z���B�����!��G�$��;�}Q��f�R0|��������a��֡��!ݱ�����Zƺ@�к�ۺg�庺�����]�����CQ�w������O��"���'�R(-��g2�o�7���<�{B�?aG���L���Q�kYW���\��5b��g�E;m�(�r��Ux�#�}�7���Ds���+��މ�>���D,���ɑ��b��n�������  �  ��=NJ=z�=��=�L=��=�=�H=� =� =�@ =i��<L!�<�q�<���<�<f�<���<�<_]�<M��<h �<UP�<מ�<���<�6�<,��<���<9�<�S�<U��<���<u!�<�f�<���<f��<;�<��<l��<��<�Z�<Ѡ�<���<&�<@d�<��<���<��<p7�<b�<���<3��<���<J��<���<��<B�<�"�<1&�<�#�<Z�<
�<���<&��<2��<�s�<�5�<���<��<>�<���<�e�<;��<�g�<���<�I�<گ�<K�<nh�<k��<m�<�O�<���<�˸<K �<�.�<)W�<qy�<㕯<ᬭ<澫<^̩<�է<ܥ<eߣ<f�<�ߟ<Gݝ<�ٛ<�ՙ<MЗ<.ʕ< Ó<��<���<¦�<��<���<D{�<�h�<�T�<A?�<(Q~<�"z<��u<��q<Ùm<{pi<uJe<�(a<Y
]<��X<�T<��P<ʲL<��H<��D<Q�@<Op<<�^8<L4<!90<9&,< (<C$<�<��<��<��<��<c�<�<�<�0 <ب�;��;c`�;���;;L�;t��;�n�;=�;?Ѽ;E��;���;8��;䠠;�ޙ;�@�;�Ȍ;�x�;�R�;t�t;�i;��];y�R;�H;F�=;{�3;�);c ; �;@�;��;���:k�:���:[��:&�:���:�E�:���:I(z:�_:#�D:�*:8F:z��9�H�9B��9_R<9�q�8�QW�aŸ�EA�����h���[�칍o��$�q|:�$�P��Af�S�{��c���Ԓ�z+��hu���������Fƺ��к�ۺ�庼𺣺��ȳ�J��i������p�?�"��(��G-���2�Ծ7���<�2B�6pG�شL��R��ZW�}�\��-b���g�W*m���r��<x�"�}�����b�����p̉�	w��t��G����T���떻�����  �  ��=KK="�=>�=�L=O�=@�=�G=�� =/� =�> =���<-�<Ql�<7��<��<a�<ʳ�<��<�Y�<\��<7��<�N�<&��<���<�7�<���<��<,�<W�<}��<u��<�&�<l�<5��<��<u@�<h��<X��<�<�^�<��<<��<�'�<Ve�<+��<l��<~�<�5�<~_�<\��<T��<M��<h��<t��<w�<�<��<R!�<�<�<��<G��<O��<#��<^s�<G6�<���<��<�@�<��<�i�<���<%m�<K��<�O�<յ�<2�<$n�<���<~�<"T�<x��<�θ<��<�0�<;X�<�y�<���<���<���<�ɩ<�ҧ<إ<�ڣ<wۡ<Wڟ<؝<�ԛ<ZЙ<q˗<�ŕ<N��<ʷ�<'��<<��<c��<�{�<"j�<�V�<�A�<�W~<z*z<��u<��q<��m<�{i<Ve<�3a<A]<K�X<t�T<6�P<��L<��H<ݕD<�@<�q<<^^8<\J4<�50<�!,<�(<��#<7�<,�<m�<��< �<W�<��<�	<�' <���;3��;�V�;���;_H�;-��;�p�;�;�ؼ;��;���;ؓ�;���;��;'U�;�݌;���;�g�;.�t;S1i;��];/�R;�%H;�=;J�3;��);w ;�;|�;��;���:K��:^�:6W�:�Ķ:R��:�:o��:�~y:�m^:^D:�.*:��:7��9=ɾ9(2�9+<9!��8q�7�6hø`@�����~���!�����?t#���9���O��e���z�c�������眺R<������׻�F.ƺ}�к2ۺ��41�i������Z*�Њ�����D������"�I0(��p-�I�2���7�=�wKB���G���L�p
R�}\W���\��#b���g��m�)�r�Ox���}� ���9M���������a��������B���ۖ�$u���  �  ��=rL=��=��=�L=��=:�=/F=�� =�� =/< =��<'�<f�<ٶ�<��<[�<T��<��<�U�<��<��<�L�<!��<���<S8�<C��<���<s�<3[�<=��<���<�,�<gr�<���<���<�F�<z��<���<�<c�<���<��<�)�<xf�<���<���<
�<73�<a\�<���<���<��<���<h��<$�<��<��<��<��<��<��<3��<��<ä�<�r�<�6�<D��<4��<�C�<���<?n�<#��<s�<���<WV�<���<�<�t�<=ǿ<X�<PY�<��<�Ҹ<��<�2�<cY�<z�<ؔ�<.��<���<xƩ<�Χ<Vӥ<�գ<�ա<9ԟ<�ѝ<DΛ<Iʙ<�ŗ<���<���<��<��<���<���<劉<|�<fk�<�X�<�D�<__~<�3z<4v<Z�q<��m<��i<6ce<�@a<�!]<Y<2�T<��P<��L<1�H<��D<2�@<�r<<�]8<H4<�10<�,<l(<��#<��<��<�<��<��<t�<3�<*�<M <[��;��;cJ�;��; C�;���;�r�;B!�;s�;굵;٠�;���;AǠ;��;Rm�;���;���;���;�u;�\i;^;��R;pAH;7�=;'�3;S�); ;�;�v;�;Ĕ�:֘�:�:��:�g�:�?�:2��:�?�:��x:n�]:�XC:��):�Z:	�9,�9�͍9�;9�ݸ8]v��z���>����7�����&!��"��9��O��d��0z������0��Қ��N����Q��D����ƺޅк�
ۺ���4M�������K����	��s����#��b(�U�-���2��
8�:=�-iB�b�G��L��R��_W�۶\�-b���g���l�byr���w�ox}�z���4���ꆻ����!G��*펻鎑�-��Sɖ�ae���  �  "�=�M=��=Ȣ=FL=	�=�=�D=�� =�� =j9 =���<��<N_�<��<��<�T�<K��<���<�P�<��<~��<�J�<���<^��<�8�<��<��<��<|_�<A��<���<�2�<y�<���<��<�M�<��<���<e"�<�g�<r��<��<�+�<�g�<���<��<j�<�0�<�X�<:}�<���<d��<e��<���<l��<��<!�<Q�<-�<��<���<���<���<8��<$r�<7�<y��<u��<�F�<���<*s�<���<Zy�<`��<�]�<��<`#�<�{�<�Ϳ<��<�^�<ȝ�<fָ<��<�4�<{Z�<5z�<
��<���<緫<�©<'ʧ<-Υ<�ϣ<Pϡ<�͟<�ʝ<�Ǜ<�Ù<}��<�<Ƶ�<ͯ�<���<F��<-��<8��<d|�<�l�<[�<�G�<Rg~<(=z<<v<��q<�m<��i<Cqe<�Na<M/]<�Y<��T<��P<d�L<ݴH<ȟD<?�@<t<< ]8<{E4<c-0<K,<M�'<�#<��<'�<��<�<��<��<��<��<� <ws�;F��;=�;���;�<�;?��;�s�;y&�;|�;*µ;���;���;�ܠ;| �;І�;K�;);Қ�;�6u;��i;�-^;@ S;�]H;�=;Y�3;a�);L ;M�;�h;Zm;�Z�:IR�:���:��:� �:�զ:��:"҉:��w:��\:R�B:��(:K�:X0�9O�9�]�9�A;9��8N�𵳂���E=��'���a��OJ鹾c���!��(8��'N���c�Zy�N��Eԑ�pI�������������ź�yк�ۺ*���k��4���p�9���D����T�ER#�Θ(���-�m
3��78�Sa=�,�B���G���L�R R��dW���\��b�Ytg���l�gYr���w�pL}��a�����Eφ�����+���Ҏ�rv�����ҵ���T���  �  ��=�N=5�=��=L=M�=�=�B=�� =� =�6 =���<	�<iX�<��<���<%N�<?��<��<$L�<��<o��<�H�<���<��<�9�<h��<���<7�<�c�<3��<;��<�8�<��<^��<W�<]T�<R��<���<�'�<Kl�<-��<���<�-�<�h�<П�<5��<��<�-�<aU�<�x�<���<���<.��<1��<���<�<q
�<�<f�<��<D��<J��<���<~��<uq�<F7�<���<���<�I�<���<�w�<M �<��<*��<�d�<6��<�*�<���<�Կ<��<3d�<m��<<ڸ<��<�6�<�[�<Ez�<6��<���<*��<J��<�ŧ<�ȥ<�ɣ<�ȡ<�Ɵ<ĝ<���<��<K��<:��<���<|��<B��<���<���<���<�|�<�m�<!]�<�J�<o~<�Fz< v<��q<.�m<�i<!e<|\a<�<]<Y<�U<��P<��L<l�H<`�D<�@<u<<>\8<�B4<�(0<�,<��'<�#<G�<��<:�<լ<r�<_�<3�<��<^ <_�;1��;m/�;(��;�6�;���;u�;(+�;��;bε;%��;˧;L�;`8�;۟�;,+�;d܆;i��;hu;	�i;NV^;�BS;zH;M�=;Կ3;L�);� ;��;�X;�V;� �:�	�:9l�:�F�:���:�h�:d��:�b�:�
w:o\:��A:�H(:M;:�F�9�ʼ9�9��:9��8�q��U���]�;��?��>F�����"�
��!�]T7��MM�	c���x��膺�x������n���ⰺ>[���ź�mк�ۺ���3��d���"����Q��t���
8���#��(��
.��;3��d8�-�=��B���G��L��,R�`iW�E�\�b��cg�u�l�%:r���w�!}��I��� �������d�����与��]��� �������D���  �  "�=�O=��=�=�K=��=��=eA=�� =ɍ =�3 =��<��<�Q�<���<���<H�<���<���<�G�<H��<x��<�F�<p��<���<:�<���<���<;�<ig�<���<^��<�>�<���<���<��<�Z�<0��<C��<�,�<fp�<���<t��</�<yi�<���<Q��<� �<c+�<�Q�<�t�<���< ��<H��<���<��<���<!�<2	�<��<��<��<���<^��<˟�<�p�<L7�<���<b��<�L�<w��<>|�<c�<7��<S��<k�<���<I1�<e��<�ڿ<3%�<0i�<���<�ݸ<=�<s8�<p\�<*z�<M��<Τ�<���<ɻ�<`��<ĥ<Lģ<�¡<��<���<,��<Ͷ�<j��<Я�<�<X��<�<#��<ڒ�<���<�|�<�n�<�^�<�M�<v~<Oz<'v<��q<7�m<��i<
�e<>ia<�H]<}*Y<3U<��P<�L<h�H<��D<��@<�u<<[8<�?4<�#0<�,<��'<��#<��<̯<q�<��<�<�<j�<��<��;�K�;���;N"�;+��;/0�;U��;�u�;5/�;H��;:ٵ;�ͮ;ܧ;��; N�;��;�C�;��;̀;��u;�i;%{^;�aS;^�H;}>;
�3;	�);� ;D�;�I;�@;5��:���:K�:P��:�;�::�:�C�:��::=v:Z[:$-A:(�':2�:e�9��9i�9�L:9��8�c��� ����:��n��fF����湧�	��a �M�6���L�0=b���w�G����%������1��1����6��W�źYdк�ۺ��庍�𺍒��[@� ���/�#����wk���#�)��<.��j3��8��=���B���G�yM��9R�2oW�L�\���a��Tg�T�l�r���w�_�|��3���胻����K������ࠎ��G���쓻/����6���  �  L�=�P=3�=0�=eK=��=��=�?=�� =ċ =�1 =ӯ�<s��<jL�<��<��<�B�<���<g��<�C�<��<���<�D�<?��<(��<^:�<���<���<� �<�j�<���<���<C�<܊�<	��<�<�_�</��<���<�0�<�s�<`��<���<�0�<j�<���<x��<I��<)�<�N�<q�<���<a��<��<���<���<��<���<�</�<���<���<���< ��<N��<�o�<X7�<h��<ݦ�<�N�<x��<��<�	�<��<��<�p�<���<�6�<��<�߿<�)�<\m�<0��<��<f�<�9�<
]�<z�<h��<:��<%��<���<���<���<s��<½�<��<㷝<���<m��<>��<��<ȧ�<ѣ�<���<�<X��<���<�|�<to�<x`�<�O�<|~<LVz<�/v<br<n�m<t�i<іe<ta<3S]<G4Y<�U<&�P<u�L<E�H<�D<t�@<>v<<Z8<.=4<�0<�,<�'<��#<�<e�<x�<-�<E�<��<V�<j�<��;P;�;���;��;���;S*�;���;�u�;2�;k �;
�;�ٮ;G�;d�;x`�;�ʓ;�W�;8	�;s��;�u;�j;2�^;&|S;��H;�>;��3;��);( ;u�;3<;�-;ӵ�:���:���:��:�:���::�:��:��u:��Z:��@:�':;:���9���9��9k�99W��8�=E��ߺ���9��hl��b�幡k	����G�5���K�K�a��w��>���ݐ�Gq��?���0������G�ź�^к�ۺ���'�𺁻��Z����\S����'6�$��4�#�X0)��g.���3�g�8���=�`�B��H�bM�ER��tW���\���a�NHg�l�l�+r��mw���|�� ��|ԃ�O����5��Y⋻v����4���ۓ�����Y*���  �  .�=/Q=��=7�=(K=V�=�=�>=�� =+� =�/ =���<<��<H�<{��<���<�>�<ɓ�<���<�@�<v��<���<,C�<@��<���<�:�<���<���<�"�<m�<q��<��<"G�<ˎ�<(��<)�<�c�<��<h��<�3�<�v�<���<��<�1�<�j�<���<���<��<K'�<�L�<>n�<'��<Ѧ�<��<K��<:��<���<���< �<� �<e��<���<���<[��<��<:o�<U7�<���<��<�P�<���<���<��<ȍ�<��<�t�<���<J;�<$��<��<�-�<�p�<���<��<�<�:�<x]�<�y�<���<�<E��<^��<Ӻ�<W��<ӻ�<���<޶�<���<S��<0��<Q��<���<z��<��<���<1��<!��<Y��<�|�<�o�<�a�<�Q�<��~<�[z<�5v<�r<#�m<��i<<�e<f|a<[]<�;Y<�U<� Q<T�L<��H<ƮD<ޒ@<zv<<,Y8<;4<�0<u�+<��'<	�#<�<��<א<R�<2�<З<��<��<M��;;.�;���;n�;���;�%�;f��;�u�;{4�;'�;��;��;��;�"�;Hn�;�ٓ;�g�;�;��;��u;pj;��^;Z�S;��H;o(>;��3;5�);� ;�;`1;�;O��:�[�:5��:�e�:%��:[f�:Ţ�:�X�:�u::.Z:@:ղ&:A�:��9"�9���9`l99�d�8�l�۹���8�j;���ķ�	�	���K��f5�ASK��a�
�v�Y�����:B���ԥ�i�����2�ź8[к� ۺ���������n����o�Y��W�C��\$��R)�Љ.���3���8���=��B��H�-M�CNR�&yW���\��a��>g���l���q��Ww�S�|�a��8Ń� v��4%���ы�}��5&���Γ�Ww��� ���  �  ��=�Q=��=4�=�J=��=_�=9>=�� =+� =�. =q��<���<iE�<ԕ�<��<�;�<K��<���<�>�<̕�<~��<7B�<���<}��<�:�<��<���<�#�<�n�<N��<,�<qI�<=��<���<��<Rf�<`��<���<�5�<4x�<Ǹ�<��<�2�<�j�<f��<I��<7��<-&�<'K�<il�<��<p��<���<���<���<��<���<u��<@��<L��<���<+��<@��<Q��<�n�<17�<E��<���<�Q�<��<~��<�<��<�<ww�<���<�=�<���<H�<�/�<�r�<���<�<��<�;�<�]�<�y�<3��<��<$��<Ҵ�<���<.��<f��<��<1��<߰�<���<���<ħ�<)��<n��<F��<J��<��<`��<ᆉ<�|�<Yp�<Lb�<�R�<+�~<N_z<�9v<	r<�m<��i<p�e<t�a<`]<8@Y<�!U<�Q<"�L<7�H<I�D<Г@<v<<qX8<�94<�0<��+<<�'<��#<?�<_�<i�<ǅ<��<;�<6�<X�<���;�%�;l��;��;\��;�"�;���;ju�;�5�;��;��;-�;��;�*�;w�;9�;Pq�;�"�;_��;c�u;0j;��^;�S;+�H;�/>;��3;��);�	 ;�{;i*;;;w�:�=�:�~�:?�:�|�:F;�:�w�:�-�:��t:�Y:t�?:�m&:&�:u��9���9�r�9�+99�(�8��*E��p8�쉹	]�����m��*��K5��K�R�`�Qv�!߅������#������?V��������ź�Xк�$ۺ��2��U���{���ڀ� ��l�����#$��h)�!�.�Q�3�j�8�$�=�C��H�n5M�TR��|W�>�\���a�>9g�t�l�W�q��Iw��|�r	��Y���l�����ȋ�5s��,���Ɠ�#p������  �  P�=�L=P�=��=%E=8�=��=�8=�� =�� =Y* =���<��<<�<���< ��<�-�<x��<���<�'�<3{�<���<� �<Er�<0��<��<�]�<<��<d��<,<�<��<���<�<�V�<a��<���<;#�< f�<���<#��<�&�<�c�<��<���<}
�<�;�<yi�<{��<���<4��<��<+�<�-�<�A�<�R�<�_�<
i�<n�<�n�<.j�<`�<[O�<}7�<��<���<��<���<�@�<���<���<K:�<���<�[�<���<Y�<;��<d5�<��<F��<bG�<���<hۻ<j�<=U�<���<��<wݲ<���<9�<<2�<�D�<S�<�]�<�e�<Xk�<@o�<�q�<�s�<�t�<�u�<^v�<�v�<�v�<�u�<�s�<�p�<wl�<�f�<_�<�U�<,K�<:?�<�c~<�Gz<�*v<�r<��m<��i<F�e<��a<0~]<�dY<MU<[6Q<S M<"I<��D<��@<��<<��8<s�4<x�0<�x,<�f(<]W$<DK <D<2B<�F<�R<�e<�<�<d� <w�;�z�;���;��;w5�;L��;l��;�x�;�\�;�T�;!b�;���;�ȣ;�%�;���; =�;s��;�ڃ;��{;}p;��d;��Y;�N;�D;4�9;��/;!�%;�;;��;?�	;�� ;`�:��:�:�/�:��:���:�#�:���:%wl:ЦQ:��7:V�:k�:4-�9ce�9�Qn9#�9�B?8�(:�x=�*fi�\���!�й��������f,�-�B�j�X�#�n�)H���!���헺G����y���@��dú��ͺ��غ���c��ǯ���[�����^�����K�a��#�7c(���-�Y�2��8��B=�zmB�]�G���L���Q�f0W�kr\�h�a�[g��kl�(�q�Z2w�Z�|����嵃��i������̋�E|��|+��ړ�1����9���  �  #�=rL=B�=��=.E=L�=ߒ=9=�� =�� =�* =���<���<�<�<!��<���<o.�<��<j��<(�<�{�<���<&!�<lr�<D��<��<�]�< ��<��<�;�<���<h��<}�<�U�<Ӛ�<��<�"�<de�<"��<���<f&�<Dc�<Ý�<���<L
�<�;�<�i�<���<��<���<s��<��<N.�<�B�<6S�<J`�<�i�<�n�<]o�<�j�<�`�<�O�<�7�<=�<��<��<���<�@�<���<1��<�9�<��<[�<��<pX�<���<�4�<\��<���<�F�<#��<�ڻ<�<�T�<h��<յ�<Kݲ<��<[�<2�<E�<}S�<a^�<Uf�<�k�<�o�<jr�<2t�<ku�<]v�<�v�<'w�<�v�<v�<0t�<q�<�l�<�f�<_�<�U�<K�<�>�<@c~<�Fz<�)v<�r<j�m<��i<�e<X�a<�|]<�cY<LU<^5Q<�M<d
I<��D<��@<��<<��8<��4<�0<�y,<�g(<=X$<jL <@E<�C<H<�S<�f<1�<^�<�� <Q�;�|�;z�;F��;36�;���;+��;Vx�;�[�;;S�;�`�;���;ǣ;�#�;��;�:�;J��;H؃;�{;�p;d�d;m~Y;أN;�D;9�9;9�/;W�%;�<;��;�	;r� ;dg�:��:�%�:}8�:R��:`��:�,�:F�:ǈl:�Q:ɒ7:��:W�:�C�9�t�9edn9��9A�>8vw:��a���i�1��ѹ���h�D{,��B���X�x�n�=Q��&)�������������D���ú3�ͺ��غd��˪�����W����hZ����3G�ί��#�^(�Q�-���2�"8�/?=��iB��G���L��Q��/W��r\�z�a��g�]nl���q�6w�t�|����u����k����ϋ��~���-��ܓ����Z;���  �  ��=,L=�=��=OE=��=?�=�9=�� =z� =�+ =h��<���<�>�<*��<���<X0�<��<��<{)�<�|�<���<�!�<�r�<|��<��<=]�<b��<��<�:�<"��<���<��<T�<ܘ�<��<� �<�c�<���<��<4%�<Ib�< ��<)��<
�<�;�<�i�<C��<ܺ�<���<���</�< 0�<ZD�<DU�<\b�<�k�<�p�<.q�<�l�<b�<Q�<�8�<��<���<P��<���<I@�<P��<b��<�8�<���<sY�<Z��<�V�<���<�2�<C��<���<�D�<v��<@ٻ<��<�S�<���<_��<ݲ<%��<��<3�<�E�<�T�<�_�<�g�<�m�<�q�<�t�<8v�<�w�<[x�<�x�<�x�<ox�<Tw�</u�<�q�<.m�<�f�<_�<�U�<�J�<>�<Ca~<aDz<�&v<$r<��m<��i<�e<h�a<y]<T`Y<�HU<�2Q<yM<�I<b�D<�@<��<<%�8<��4<��0<|{,< j(<)[$<�O < I<�G<hL<�W<]k<+�<7�<� <G�;	��;W�;���;-8�;��;N��;^w�;�Y�;�O�;�\�;]��;5��;-�;ߗ�;`3�;}��; у;��{;_�o;�d;huY;��N;D;h�9;ĥ/;��%;k?;p�;��	;� ;�|�:���:1C�:-V�:��:�:N�:(�:�l: �Q:4�7:�#:��:�w�9��90�n9R�9
{>8�9;�w��Vj�!a���sѹ= ���=�o�,��C�RY�go�sm��B�����Y͢�r���`O���ú��ͺT�غ�����~����N�y��GM���8�����"�3M(�a�-��2��8�i3=�J_B�(�G��L��Q��-W�Ir\���a��g�ul���q�b@w���|��
���s��1&���֋�j���v4��6⓻w���l?���  �  	�=�K=��=x�=yE=��=�=^:=�� =�� =�, =L��<���<B�<k��<���<_3�<���<���<�+�<�~�<P��<#�<�s�<���<s�<�\�<V��<���<�8�<��<R��<��<.Q�<ԕ�<��<��<�`�<��<���<'#�<�`�<ɛ�<H��<�	�<�;�<[j�<B��<;��<n��<���<��<�2�<WG�<AX�<�e�<�n�<�s�<*t�<Eo�<td�<2S�<�:�<U�<���<���<���<�?�<Y��<��<7�<���<W�<���<�S�<x��<m/�<��<���<�A�<���<�ֻ<��<!R�<d��<{��<�ܲ<)��<)�<4�<JG�<dV�<�a�<[j�<xp�<�t�<�w�<ry�<�z�<^{�<�{�<�{�<�z�<ly�<�v�<;s�<n�<Yg�<_�<U�<�I�<�<�<�]~<1@z<�!v<�r<��m<��i<˨e<S�a<Gs]<�ZY<�CU<@.Q<�M<�I<O�D<��@<o�<<��8<P�4<�0<�~,<0n(<�_$<EU <�N<�M<�R<�^<�q<{�<�<w� <�;a��;6�;���;�;�;���;@��;Vu�;*V�;�J�;�U�;_y�;���;��;��;�'�;��;�Ń;��{;1�o;��d;�eY;��N;�C;�9;��/;W�%;�C;��;Q�	;�� ;)��:���:�n�:߆�:j�:��:ʁ�:�X�:�%m:�MR:|8:�j:�7:��9ߧ9�n98�9��=8�<��S�5�j�9⣹-ҹ�������-�eC��Y��lo����ak���/���좺A����`��D"ú	�ͺ��غ��㺃��1���v?�W��>9�����d����"��3(�J{-���2���7� =��NB��~G�^�L���Q��*W��r\���a�%g�Sl�+�q�$Qw�˽|�o��"˃�`��Q2���⋻����F?���듻ꘖ��F���  �  *�=K=��=e�=�E=o�=��=l;=�� =0� =~. =��<���<*F�<���<��<p7�<u��<���<�.�<E��<L��<`$�<ft�<���<.�<�[�<���<���<`6�<$}�<���<V�<AM�<ё�<��<��<�\�<^��<���<~ �<x^�<3��<-��<A	�<�;�< k�<]��<��<���<��<��<B6�<=K�<M\�<�i�<�r�<�w�<x�<�r�<�g�<�U�<�<�<�<���<Q��<���<P?�<#��<Z��<�4�<���<�S�<���<�O�<6��<6+�<ȍ�<L��<�=�<��<�ӻ<��<�O�<���<d��<7ܲ<-��<��<:5�<I�<�X�<�d�<�m�<t�<�x�<�{�<�}�<�~�<t�<��<�<�}�<|�< y�<�t�<,o�<�g�<_�<�T�<wH�< ;�<6Y~<�:z<Mv<��q<@�m<Ľi<Ġe<#�a<fk]<sSY<D=U<�(Q<�M<%I<��D<d�@<�<<��8<'�4<�0<��,<Ls(<%f$<"\ <�V<V<\[<gg<Lz<�<�<� <�#�;���;��;��;@�;���;��;�r�;�Q�;.D�;�L�;�n�;��;��;	~�;o�;�Չ;O��;�w{;T�o;�jd;�QY;�N;n�C;<�9;�/;t�%;�I;��;�	;u;<��:���:c��:kƿ:IU�:SW�:�Œ:r��:?�m:~�R:�|8:5�:s�:�E�9�*�9a.o9��9�=8��>�J���k����f�ҹ�R ���B�-�@�C�� Z�q�o��Ԃ�7���V^����Uŭ��w��U0úF�ͺ}�غ��Iy�}e��5,�n�����������e���"��(��Z-�ؙ2��7�u=�6:B�PmG��L���Q��&W��s\�*�a��'g�Ռl�Z�q��fw�V�|��#��wڃ�����$B����!����M������񣖻P���  �  �=DJ=�=K�=�E=��=|�=�<=Q� =�� =�0 =_��<R��<�J�<o��<���<�;�<���<���<2�<��<���<�%�<bu�<Y��<��<�Z�<9��<s��<�3�<�y�<��<%�<�H�<&��<W��<(�<�X�<W��<��<f�<�[�<.��<���<��<�;�<�k�<���<߿�<=��<��<w!�<\:�<�O�<�`�<nn�<�w�<�|�<`|�<�v�<Jk�<�X�<k?�<��<���<���<���<�>�<���<1��<2�<���<�O�<���<K�<U��<<&�<Ԉ�<x��<~9�<䇽<�ϻ<��<LM�<���<��<�۲<@��<��<�6�<K�<D[�<�g�<Sq�<)x�<}�<L��<f��<���<��<ꃗ<$��<���<�<�{�<�v�<fp�<�h�<�^�<�S�<�F�<�8�<�S~<@4z<�v<S�q<U�m<_�i<+�e<�{a<Qb]<KY<y5U<�!Q<2M<��H<P�D<y�@<z�<<c�8<H�4<w�0<��,</y(<@m$<Td <e_<�_<4e<Fq<-�<L�<��<�� <2�;'��;��;a��;�D�;���;���;�o�;yK�;�;�;_B�;�a�;n��;���;�l�;��;�É;���;pV{;��o;�Nd;H:Y;�lN;p�C;ԟ9;�/;��%;;P;�;��	;�;���:<�:e��:��:_��:���:��:��:�1n:ES:��8:U(:��:���9���9m�o9��9��;8i]A���%m�gK����ӹ�� ����(.��zD�N�Z��|p�d���ߍ�2���yC���뭺����HAú��ͺָغ^��Ca��B��5��������p�����?�m�"�^�'��5-�qw2���7���<�p"B��YG���L���Q�"W��t\���a��3g��l��r��w�o�|�4��$샻%���U��{������,^�� ��L����Z���  �  �=rI=��= �=F=��=h�=�==�� =�� =�2 =���<:�<P�<���<���<�@�<8��<���<�5�<��<���<�'�<Pv�<���<P�<�Y�<l��<���<]0�<�u�<��<x��<�C�<��<+��<3�<�S�<��<��<��<Y�<��<k��<��<�;�<Cl�<��<���<���<��<=%�<�>�<=T�<�e�<}s�<�|�<|��<��<${�<	o�<3\�<B�<��<-��<n��<P��<�=�<&��<��</�<���<�K�<���<�E�<��<� �<f��<>��<w4�<Z��<�˻<8�<qJ�<���<���<�ڲ<$��<!�<�7�<M�<�]�<+k�<-u�<�|�<Ɓ�<S��<|��<���<��<���<k��<Y��<T��<0~�<�x�<�q�<i�<�^�<�R�<vE�<�6�<N~<&-z<�v<@�q<��m<;�i<��e<nqa<hX]<�AY<$-U<EQ<�M<��H<��D<K�@<��<< �8<r�4<�0<��,<(<�t$<�l <�h<�i<�o<�{<��<j�<J�<X� <)A�;��;#)�;F��;�I�;���;���;[l�;NE�;�2�;�6�;�S�;���;"�;Z�;�;���;���;�1{;��o;�0d; Y;mWN;��C;��9;@�/;��%;�U;�;�
;�2;y5�:�y�:51�:2Y�:�:���:,e�:�7�:p�n:��S:6q9:˕:*.:�N�9��9{�o9t�9@}:8�D���"�n��#����Թu]��0�}�.��E�E:[�Sq��c���#��TӘ�Ow�����Ĳ���Tú� κҶغ�x�G�.�����o���M�P����tq"�u�'�-�AR2��7�X�<��B��EG�J�L���Q��W��v\�6�a�J@g�.�l�]%r�X�w��}�F������2����i�����eƎ�ip��_������g���  �  ��=�H=�=��=NF=�=?�=?=i� =�� =�4 =���<�<U�<���<���<�E�<���<���<'9�<���<��<2)�<4w�<���<��<\X�<��<j��<-�<<r�<���<���<�>�<���<��<"�<O�<v��<%��<y�<=V�<ݓ�<���<��<�;�<�l�<G��<���<x��<7�<�(�<�B�<�X�<�j�<�x�<��<Y��<�<^�<�r�<o_�<�D�<�!�<[��<���< ��<�<�<g��<���<,�<B��<�G�<J��<�@�<ı�<Y�<�}�<���<u/�<�~�<�ǻ<�
�<�G�<A~�<���<�ٲ<
��<��<>9�<O�<�`�<�n�<y�<倣<���<<��<���<Í�<퍙<@��<���<��<���<���<~z�<�r�<�i�<�^�<�Q�<�C�<q4�<H~<&z<zv<�q<��m<�i<H�e<ga<pN]<I8Y<�$U<�Q<�M<��H<�D<��@<��<<��8<t�4<q�0<`�,<��(<�{$<1u <3r<�s<z<��<�<��<��<�� <@P�;���;3�;q��;WN�;���;ʤ�;]h�;�>�;�)�;�*�;�E�;|�;jќ;/G�;vߏ;��;&~�;�{;�io;�d;�Y;�AN;x�C;׉9;�/;-�%;�[;�;
;%H;(k�:q��:Vv�:ѥ�:�A�:�I�:O��::�do:�]T:6�9:l :H�:���9�7�9fAp9��9�98�$G��#�"�o�����$�չ&������g/���E���[���q�%����h�����h����>���Ҹ�fjú9	κ��غ�k㺎/�����I��-T�s���)����H"�Ӛ'���,�-2��o7�ѯ<���A�%2G�6yL���Q��W��x\���a�:Ng���l�x=r�۹w�P6}�]X�����ʆ�F~��.���َ�҂��
)��%Ζ�us���  �  ��=�G=~�=��=nF=��=�=#@=�� =C� =�6 =���<�
�<�Y�<v��<��<J�<ƚ�<���<_<�<���<.��<�*�< x�<���<>�<(W�<���<���<*�<�n�<���<~��<;:�<'~�<E��<a�<�J�<E��<L��<2�<�S�<���<W��<�<q;�<Ym�<Z��<���<���<!�<�,�<�F�<&]�<Uo�<8}�<���<���<���<E��<Qv�<Sb�<�F�<�#�<_��<[��<ʃ�<�;�<���<J��<7)�<պ�<�C�<���<5<�<���<I�<�x�<���<�*�<Qz�<�û<I�<�D�<|�<z��<ٲ<���<@�<k:�<�P�<c�<�q�<�|�<؄�<ˊ�<Ύ�<P��<j��<n��<r��<��<���<`��<��<C|�<�s�<�i�<8^�<�P�<,B�<52�<eB~<6z<��u<��q<��m<J�i<�xe<U]a<$E]<�/Y<gU<�Q<��L<��H<p�D<��@<��<<
�8<5�4<��0<�,<;�(<Ԃ$<�| <�z<�|<��<S�<��<��<A�<�<^�;E��;�<�;H��;�R�;��;V��;�d�;!8�;� �;��;h8�;m�;��;b5�;!͏;É�;�k�;��z;lIo;p�c;��X;m-N;��C;=9;�/; �%;b`;($;�#
;1\;A��:���:B��:���:B��:h��:��:�Ѕ:g�o:��T:ua::�a :��:,K�9K��9��p9��9vy787�I�F,�g9q��ʧ���ֹip�dV�L�/��\F�w\��Or�u�˪��SJ��-ݣ�/g���񸺯~ú�κ��غ0`㺻��������!;�͢�8	��k�(��H""�u'���,��2��P7�@�<�>�A��G��kL�&�Q�KW��{\�'�a�=[g�	�l�Tr��w��U}�Ii��%���݆�b���.A��9쎻Փ��9��	ܖ��~���  �  z�=�F=�=��=�F=��=��=A=�� =�� =/8 =U��<r�<�]�<k��<���<�M�<T��<���<?�<؎�<���<�+�<�x�<���<��<"V�<��<���<�'�<�k�<)��<���<%6�<�y�<��<G�<�F�<���< ��<]�<Q�<Տ�<��<I�<B;�<�m�<E��<��<���<��<x/�<3J�<�`�<Fs�<*��<u��<Վ�<���<���<>y�<�d�<�H�<�$�<B��<���<���<�:�<t��<I��<�&�<ڷ�<@�<��<�7�<m��<��<zt�<���<�&�<�v�<v��<d�<EB�<0z�<.��<3ز<���<��<b;�<kR�<'e�<t�<��<J��<���<ђ�<A��<k��<W��<��<Ԓ�<n��<܊�<���<�}�<�t�<7j�<�]�<%P�<�@�<70�<y=~<Oz<��u<�q<f�m<��i< pe<�Ta<�<]<�'Y<�U<�Q<_�L<s�H<o�D<��@<��<<L�8<��4<.�0<r�,<�(<v�$<�� <�<��<��<��<"�<��<��<o<�i�;	��;D�;���;�U�;'��;��;>a�;�2�;��; �;�,�;`�;A��;�%�;%��;{y�;$\�;��z;�-o;?�c;9�X;aN;p�C;>v9;��/;��%;�c;?,;�/
;�l;*��:�!�:N��:D&�:w˱:�բ:D�:Q�:,fp:cLU:�::`� :S:��9`é9e�p9��9�68�HL��Zer�U|��g_׹�������0���F��\�X�r��2��3⎺}�����"������ú�κ��غyX㺫����;���%�ۉ� ���M�����"�ZU'���,���1��67��}<���A��G��`L��Q�lW�O~\�/�a�fg�*�l��gr���w��p}�?x��[5��W����Q����������{F��薻����  �  ��=YF=��=b�=�F='�=2�=�A=�� =�� =k9 =��<E�<�`�<t��<� �<�P�<��<4��<'A�<���<��<�,�<�x�<���<M�<6U�<���<��<p%�<i�<���<���<"3�<�v�<˺�<9��<�C�<އ�<���<�<@O�<V��<���<��< ;�<�m�<��<+��<Z��<��<�1�<�L�<�c�<v�<1��<y��<���<a��<3��<`{�<�f�<iJ�<�%�<���<���<W��<:�<;��<���<�$�<y��<|=�<(��<�4�<7��<k�<q�<u��<�#�<�s�<׽�<�<W@�<�x�<��<�ײ<���<��<'<�<�S�<�f�<v�<܁�<ኣ<E��<���<E��<o��<0��<ڗ�<]��<���<Ɍ�<e��<�~�<bu�<jj�<�]�<iO�<�?�<�.�<�9~<�z<��u<Q�q<K�m<��i<iie<�Na<�6]< "Y<3U<� Q<?�L<�H<��D<��@<7�<<�8<��4<&�0<#�,<��(<Ì$<�� <��<z�<-�<Ȟ<G�<��<X�<v<�r�;���;�I�;*��;�W�;���;��;2^�;�-�;u�;H�;�#�;V�;��;D�;���;m�;pP�;u�z;]o;3�c;�X;<N;C�C;�m9;%�/;�%;2f;�2;89
;'y;w��:E�:W�:rS�:���:��:4u�:�?�:�p:W�U:�;:�� :sI:h��9f��9V�p9�9��48LwN�3���Ns�L
����׹R:��6��0��JG��b]��2s��b����� ����)��0����!����ú�$κd�غuR�j��������G�Xw����C7�J��C�!�*='��,���1�d"7��l<���A��G��XL���Q�"W�?�\�N�a��og���l��wr�_�w�
�}�����uA�����Z���+^�����s����P��������  �  5�=�E=c�=B�=�F=O�=z�=$B=j� =c� =/: =���<)�<�b�<~��<g�<}R�<���<���<mB�<���<���<=-�<By�<���<�<�T�<��<��<#$�<�g�<���<���<1�<�t�<���<��<�A�<��<���<��<N�<���<N��<M�<�:�<n�<`��<���<H��<��<3�<TN�<Xe�< x�<*��<w��<���<(��<�<�|�<�g�<RK�<�&�<I��<���<��<�9�<���<͉�<}#�<��<�;�<6��<�2�<���<=�<�n�<I��<�!�<�q�<4��<� �<3?�<�w�<e��<5ײ<O��<��<�<�<?T�<�g�<2w�<Q��<x��<��<���<J��<a��<��<���<ꖕ<��<ۍ�<T��<W�<�u�<}j�<�]�<O�<�>�<�-�<*7~<�z<W�u<��q<n�m<h�i<Iee<LJa<�2]<@Y<�U<��P<��L<*�H<B�D<��@<��<<z�8<8�4<C�0<�,<ҕ(<��$<Ë < �<Z�<-�<��<9�<e�<��<�<x�;	��;fM�;���;tY�;"��;[��;�\�;=+�;��;y	�;�;7O�;��;��;䨏;1e�;KH�;��z;<
o;ļc;��X;|N;�C;i9;�/;��%;�g;6;�>
;�;���:]�:�0�:9p�:��:'�:���:c^�:4�p:��U:^8;:`!:=h:g#�9r�9��p9�9:48�O��5���s��`���bعu�hr�}&1���G�!�]�Xts�%���#*��V����>�������.��o�ú�)κ�غ�N㺊����������Kk����z(�����!��-'��},���1�7�ca<�2�A�v�F��SL�D�Q��W��\���a��ug���l�>�r��
x���}�늁�I�����~����f��e��˵���W��?�������  �   �=�E=Q�=9�=�F=]�=��=SB=�� =�� =m: =P��<��<Pc�<��<��<S�</��<>��<�B�<��<E��<c-�<hy�<���<��<T�<���<���<�#�<(g�<��<E��<r0�<t�<6��<h��<A�<h��<Z��<O�<�M�<%��<��<"�<�:�<-n�<���<��<���<�<�3�<�N�<�e�<�x�<���<��<1��<���<5��<^}�<;h�<�K�<�&�<m��<
��<��<�9�<B��<k��<#�<���<@;�<���<72�<>��<��<Bn�<���<� �<*q�<���<+ �<�>�<bw�<%��<ײ<I��< �<�<�<�T�<h�<�w�<ڃ�<���<���<)��<ܚ�<�<���<)��<b��<���<7��<���<��<�u�<�j�<v]�<�N�<�>�<g-�<06~<�z<8�u<`�q<+�m<�i<0de<�Ha<g1]<Y<�U<��P<��L<O�H<��D<��@<��<<��8<q�4<��0<��,<��(<��$<�� <@�<��<]�<4�<k�<��<��<�<�y�;���;�N�;7��;/Z�;^��;)��;�[�;*�;N�;��;i�; M�;㝜;��;���;*c�;�E�;��z;}o;��c;f�X;N;b�C;g9;�~/;}�%;�h;r7;A
;�;v��:�e�:*8�:}y�:9#�:�/�:���:�h�:�q:R�U:FJ;:w&!:zs:5�9��9�q9��9P�38n-P��b��t��{����ع��0��.=1�F�G��]�_�s�܈���3���Ù�
F��u����3��ݫúf+κ�غ�K�<��Ҝ������f�����#�t~�g�!�)'�xx,�@�1�a7�O]<�a�A�y�F�RL�-�Q�!W���\���a�xg���l�)�r�x��}�e����K���������\i�����7����Y�����������  �  5�=�E=c�=B�=�F=O�=z�=$B=j� =c� =/: =���<)�<�b�<~��<g�<}R�<���<���<mB�<���<���<=-�<By�<���<�<�T�<��<��<#$�<�g�<���<���<1�<�t�<���<��<�A�<��<���<��<N�<���<N��<M�<�:�<n�<`��<���<H��<��<3�<TN�<Xe�< x�<*��<w��<���<(��<�<�|�<�g�<RK�<�&�<I��<���<��<�9�<���<͉�<}#�<��<�;�<6��<�2�<���<=�<�n�<I��<�!�<�q�<4��<� �<4?�<�w�<e��<5ײ<O��<��<�<�<@T�<�g�<2w�<Q��<x��<��<���<J��<a��<��<���<ꖕ<��<ۍ�<T��<W�<�u�<}j�<�]�<O�<�>�<�-�<*7~<�z<W�u<��q<n�m<h�i<Iee<LJa<�2]<@Y<�U<��P<��L<+�H<C�D<��@<��<<z�8<8�4<C�0<�,<ҕ(<��$<Ë < �<Z�<-�<��<9�<e�<��<�<x�;	��;fM�;��;tY�;!��;[��;�\�;<+�;��;y	�;�;7O�;��;��;䨏;1e�;JH�;��z;<
o;ļc;��X;|N;�C;i9;�/;��%;�g;6;�>
;�;���:]�:�0�:9p�:��:'�:���:b^�:4�p:��U:^8;:`!:=h:g#�9r�9��p9�9:48�O��5���s��`���bعu�hr�}&1���G�!�]�Xts�%���#*��V����>�������.��o�ú�)κ�غ�N㺊����������Kk����z(�����!��-'��},���1�7�ca<�2�A�v�F��SL�D�Q��W��\���a��ug���l�>�r��
x���}�늁�I�����~����f��e��˵���W��?�������  �  ��=YF=��=b�=�F='�=2�=�A=�� =�� =k9 =��<E�<�`�<t��<� �<�P�<��<4��<'A�<���<��<�,�<�x�<���<M�<6U�<���<��<p%�<i�<���<���<"3�<�v�<˺�<9��<�C�<އ�<���<�<@O�<V��<���<��< ;�<�m�<��<+��<Z��<��<�1�<�L�<�c�<v�<1��<y��<���<a��<3��<`{�<�f�<iJ�<�%�<���<���<W��<:�<;��<���<�$�<y��<|=�<(��<�4�<7��<k�<q�<u��<�#�<�s�<ؽ�<�<W@�<�x�<��<�ײ<���<��<'<�<�S�<�f�<v�<܁�<ኣ<E��<���<E��<o��</��<ڗ�<]��<���<Ɍ�<e��<�~�<au�<jj�<�]�<hO�<�?�<�.�<�9~<�z<��u<Q�q<K�m<��i<iie<�Na<�6]< "Y<3U<� Q<?�L<�H<��D<��@<7�<<�8<��4<&�0<$�,<��(<Ì$<�� <��<z�<-�<Ȟ<G�<��<X�<v<�r�;���;�I�;)��;�W�;���;��;2^�;�-�;u�;H�;�#�;V�;��;D�;���;m�;pP�;t�z;\o;2�c;�X;<N;C�C;�m9;%�/;�%;1f;�2;89
;'y;w��:E�:W�:rS�:���:��:4u�:�?�:�p:W�U:�;:�� :sI:h��9f��9V�p9�9��48LwN�3���Ns�L
����׹R:��6��0��JG��b]��2s��b����� ����)��0����!����ú�$κd�غuR�j��������G�Xw����C7�J��C�!�*='��,���1�d"7��l<���A��G��XL���Q�"W�?�\�N�a��og���l��wr�_�w�
�}�����uA�����Z���+^�����s����P��������  �  z�=�F=�=��=�F=��=��=A=�� =�� =/8 =U��<r�<�]�<k��<���<�M�<T��<���<?�<؎�<���<�+�<�x�<���<��<"V�<��<���<�'�<�k�<)��<���<%6�<�y�<��<G�<�F�<���< ��<]�<Q�<Տ�<��<I�<B;�<�m�<E��<��<���<��<x/�<3J�<�`�<Fs�<*��<u��<Վ�<���<���<>y�<�d�<�H�<�$�<B��<���<���<�:�<t��<I��<�&�<ڷ�<@�<��<�7�<m��<��<zt�<���<�&�<�v�<v��<d�<EB�<0z�<.��<3ز<���<��<c;�<kR�<'e�<t�<��<J��<���<ђ�<A��<k��<W��<��<Ԓ�<n��<܊�<���<�}�<�t�<7j�<�]�<$P�<�@�<70�<y=~<Nz<��u<�q<f�m<��i< pe<�Ta<�<]<�'Y<�U<�Q<`�L<s�H<p�D<��@<��<<L�8<��4<.�0<r�,<�(<v�$<�� <�<��<��<��<"�<��<��<n<�i�;��;D�;���;�U�;'��;��;=a�;�2�;��;��;�,�;`�;@��;�%�;%��;zy�;#\�;��z;�-o;?�c;9�X;`N;p�C;=v9;��/;��%;�c;?,;�/
;�l;*��:�!�:N��:D&�:w˱:�բ:D�:Q�:,fp:cLU:�::`� :S:��9`é9e�p9��9�68�HL��Zer�U|��g_׹�������0���F��\�X�r��2��3⎺}�����"������ú�κ��غyX㺫����;���%�ۉ� ���M�����"�ZU'���,���1��67��}<���A��G��`L��Q�lW�O~\�/�a�fg�*�l��gr���w��p}�?x��[5��W����Q����������{F��薻����  �  ��=�G=~�=��=nF=��=�=#@=�� =C� =�6 =���<�
�<�Y�<v��<��<J�<ƚ�<���<_<�<���<.��<�*�< x�<���<>�<(W�<���<���<*�<�n�<���<~��<;:�<'~�<E��<a�<�J�<E��<L��<2�<�S�<���<W��<�<q;�<Ym�<Z��<���<���<!�<�,�<�F�<&]�<Uo�<8}�<���<���<���<E��<Qv�<Sb�<�F�<�#�<_��<[��<ʃ�<�;�<���<J��<7)�<պ�<�C�<���<5<�<���<I�<�x�<���<�*�<Qz�<�û<J�<�D�<|�<z��<ٲ<���<@�<k:�<�P�<c�<�q�<�|�<؄�<ˊ�<Ύ�<Q��<j��<n��<r��<��<���<`��<��<C|�<�s�<�i�<7^�<�P�<,B�<52�<eB~<6z<��u<��q<��m<J�i<�xe<U]a<$E]<�/Y<gU<�Q<��L<��H<q�D<��@<��<<�8<5�4<��0<�,<;�(<Ղ$<�| <�z<�|<��<S�<��<��<A�<�<^�;D��;�<�;G��;�R�;��;U��;�d�; 8�;� �;��;g8�;m�;��;b5�; ͏;É�;�k�;��z;kIo;o�c;��X;l-N;��C;<9;�/;�%;a`;'$;�#
;0\;A��:���:B��:���:B��:h��:��:�Ѕ:g�o:��T:ua::�a :��:,K�9K��9��p9��9vy787�I�F,�g9q��ʧ���ֹip�dV�L�/��\F�w\��Or�u�˪��SJ��-ݣ�/g���񸺯~ú�κ��غ0`㺻��������!;�͢�8	��k�(��H""�u'���,��2��P7�@�<�>�A��G��kL�&�Q�KW��{\�'�a�=[g�	�l�Tr��w��U}�Ii��%���݆�b���.A��9쎻Փ��9��	ܖ��~���  �  ��=�H=�=��=NF=�=?�=?=i� =�� =�4 =���<�<U�<���<���<�E�<���<���<'9�<���<��<2)�<4w�<���<��<\X�<��<j��<-�<<r�<���<���<�>�<���<��<"�<O�<v��<%��<y�<=V�<ݓ�<���<��<�;�<�l�<G��<���<x��<7�<�(�<�B�<�X�<�j�<�x�<��<Y��<�<^�<�r�<o_�<�D�<�!�<[��<���< ��<�<�<g��<���<,�<C��<�G�<J��<�@�<ı�<Y�<�}�<���<u/�<�~�<�ǻ<�
�<�G�<A~�<���<�ٲ<��<��<>9�<O�<�`�<�n�<y�<倣<���<<��<���<Í�<썙<@��<���<��<���<���<~z�<�r�<�i�<�^�<�Q�<�C�<q4�<H~<&z<yv<�q<��m<�i<H�e<ga<pN]<I8Y<�$U<�Q<�M<��H<�D<��@<��<<��8<u�4<q�0<`�,<��(<�{$<1u <3r<�s<z<��<�<��<��<�� <?P�;���;3�;p��;VN�;���;ɤ�;\h�;�>�;�)�;�*�;�E�;~|�;iќ;.G�;vߏ;��;%~�;�{;�io;�d;�Y;�AN;w�C;։9;�/;,�%;�[;�;
;%H;(k�:q��:Vv�:ѥ�:�A�:�I�:O��::�do:�]T:6�9:l :H�:���9�7�9eAp9��9�98�$G��#�"�o�����$�չ&������g/���E���[���q�%����h�����h����>���Ҹ�fjú9	κ��غ�k㺎/�����I��-T�s���)����H"�Ӛ'���,�-2��o7�ѯ<���A�%2G�6yL���Q��W��x\���a�:Ng���l�x=r�۹w�P6}�]X�����ʆ�F~��.���َ�҂��
)��%Ζ�us���  �  �=rI=��= �=F=��=h�=�==�� =�� =�2 =���<:�<P�<���<���<�@�<8��<���<�5�<��<���<�'�<Pv�<���<P�<�Y�<l��<���<]0�<�u�<��<x��<�C�<��<+��<3�<�S�<��<��<��<Y�<��<k��<��<�;�<Cl�<��<���<���<��<=%�<�>�<=T�<�e�<}s�<�|�<|��<��<${�<	o�<3\�<B�<��<-��<n��<P��<�=�<&��<��</�<���<�K�<���<�E�<��<� �<f��<>��<x4�<Z��<�˻<8�<qJ�<���<���<�ڲ<$��<!�<�7�<M�<�]�<+k�<-u�<�|�<Ɓ�<S��<|��<���<��<���<j��<Y��<S��<0~�<�x�<�q�<i�<�^�<�R�<vE�<�6�<N~<&-z<�v<@�q<��m<;�i<��e<nqa<hX]<�AY<$-U<FQ<�M<��H<��D<L�@<��<<�8<r�4<�0<��,<(<�t$<�l <�h<�i<�o<�{<��<i�<J�<W� <(A�;��;")�;E��;�I�;���;���;Yl�;ME�;�2�;�6�;�S�;���;!�;Z�;�;���;���;�1{;��o;�0d; Y;lWN;��C;��9;@�/;��%;�U;�;�
;�2;x5�:�y�:51�:2Y�:�:���:,e�:�7�:p�n:��S:6q9:˕:*.:�N�9��9{�o9t�9@}:8�D���"�n��#����Թu]��0�}�.��E�E:[�Sq��c���#��TӘ�Ow�����Ĳ���Tú� κҶغ�x�G�.�����o���M�P����tq"�u�'�-�AR2��7�X�<��B��EG�J�L���Q��W��v\�6�a�J@g�.�l�]%r�X�w��}�F������2����i�����eƎ�ip��_������g���  �  �=DJ=�=K�=�E=��=|�=�<=Q� =�� =�0 =_��<R��<�J�<o��<���<�;�<���<���<2�<��<���<�%�<bu�<Y��<��<�Z�<9��<s��<�3�<�y�<��<%�<�H�<&��<W��<(�<�X�<W��<��<f�<�[�<.��<���<��<�;�<�k�<���<߿�<=��<��<w!�<\:�<�O�<�`�<nn�<�w�<�|�<`|�<�v�<Jk�<�X�<k?�<��<���<���<���<�>�<���<2��<2�<���<�O�<���<K�<U��<<&�<Ԉ�<x��<~9�<䇽<�ϻ<��<LM�<���<��<�۲<@��<��<�6�<K�<D[�<�g�<Tq�<*x�<}�<L��<f��<���<��<ꃗ<$��<���<�<�{�<�v�<fp�<�h�<�^�<�S�<�F�<�8�<�S~<?4z<�v<S�q<U�m<_�i<+�e<�{a<Qb]<KY<z5U<�!Q<2M<��H<P�D<y�@<{�<<d�8<H�4<x�0<��,</y(<@m$<Td <e_<�_<4e<Fq<,�<L�<��<�� <2�;&��;��;`��;�D�;���;���;�o�;xK�;�;�;^B�;�a�;m��;���;�l�;��;�É;���;oV{;��o;�Nd;G:Y;�lN;o�C;ӟ9;�/;��%;;P;�;��	;�;���:<�:e��:��:_��:���:��:��:�1n:ES:��8:U(:��:���9���9m�o9��9��;8i]A���%m�gK����ӹ�� ����(.��zD�N�Z��|p�d���ߍ�2���yC���뭺����HAú��ͺָغ^��Ca��B��5��������p�����?�m�"�^�'��5-�qw2���7���<�p"B��YG���L���Q�"W��t\���a��3g��l��r��w�o�|�4��$샻%���U��{������,^�� ��L����Z���  �  *�=K=��=e�=�E=o�=��=l;=�� =0� =~. =��<���<*F�<���<��<p7�<u��<���<�.�<E��<L��<`$�<ft�<���<.�<�[�<���<���<`6�<$}�<���<V�<AM�<ё�<��<��<�\�<^��<���<~ �<x^�<3��<-��<A	�<�;�< k�<]��<��<���<��<��<B6�<=K�<M\�<�i�<�r�<�w�<x�<�r�<�g�<�U�<�<�<�<���<Q��<���<P?�<#��<Z��<�4�<���<�S�<���<�O�<6��<6+�<ȍ�<M��<�=�<��<�ӻ<��<�O�<���<e��<7ܲ<.��<��<:5�<I�<�X�<�d�<�m�<t�<�x�<�{�<�}�<�~�<t�<��<�<�}�<
|�< y�<�t�<,o�<�g�<_�<�T�<wH�<;�<5Y~<�:z<Mv<��q<@�m<Ľi<Ġe<#�a<fk]<sSY<D=U<�(Q<�M<%I<��D<e�@<�<<��8<'�4<�0<��,<Ms(<%f$<"\ <�V<V<\[<gg<Lz<�<�<~� <�#�;���;��;��;@�;���;��;�r�;�Q�;-D�;�L�;�n�;��;��;~�;n�;�Չ;N��;�w{;S�o;�jd;�QY;�N;m�C;<�9;�/;t�%;�I;��;�	;u;;��:���:c��:kƿ:IU�:SW�:�Œ:r��:?�m:~�R:�|8:5�:s�:�E�9�*�9a.o9��9�=8��>�J���k����f�ҹ�R ���B�-�@�C�� Z�q�o��Ԃ�7���V^����Uŭ��w��U0úF�ͺ}�غ��Iy�}e��5,�n�����������e���"��(��Z-�ؙ2��7�u=�6:B�PmG��L���Q��&W��s\�*�a��'g�Ռl�Z�q��fw�V�|��#��wڃ�����$B����!����M������񣖻P���  �  	�=�K=��=x�=yE=��=�=^:=�� =�� =�, =L��<���<B�<k��<���<_3�<���<���<�+�<�~�<P��<#�<�s�<���<s�<�\�<V��<���<�8�<��<R��<��<.Q�<ԕ�<��<��<�`�<��<���<'#�<�`�<ɛ�<H��<�	�<�;�<[j�<B��<;��<n��<���<��<�2�<WG�<AX�<�e�<�n�<�s�<*t�<Eo�<td�<2S�<�:�<U�<���<���<���<�?�<Y��<��<7�<���<W�<���<�S�<x��<n/�<��<���<�A�<���<�ֻ<��<!R�<e��<|��<�ܲ<)��<)�< 4�<JG�<dV�<�a�<[j�<xp�<�t�<�w�<ry�<�z�<^{�<�{�<�{�<�z�<ly�<�v�<;s�<n�<Xg�<_�<U�<�I�<�<�<�]~<1@z<�!v<�r<��m<��i<˨e<S�a<Gs]<�ZY<�CU<@.Q<�M<�I<O�D<��@<o�<<��8<P�4<�0<�~,<0n(< `$<EU <�N<�M<�R<�^<�q<{�<�<w� <�;`��;5�;��;�;�;���;?��;Vu�;*V�;�J�;�U�;_y�;���;��;��;�'�;��;�Ń;��{;1�o;��d;�eY;��N;�C;�9;��/;W�%;�C;��;Q�	;�� ;)��:���:�n�:߆�:j�:��:ʁ�:�X�:�%m:�MR:|8:�j:�7:��9ߧ9�n98�9��=8�<��S�5�j�9⣹-ҹ�������-�eC��Y��lo����ak���/���좺A����`��D"ú	�ͺ��غ��㺃��1���v?�W��>9�����d����"��3(�J{-���2���7� =��NB��~G�^�L���Q��*W��r\���a�%g�Sl�+�q�$Qw�˽|�o��"˃�`��Q2���⋻����F?���듻ꘖ��F���  �  ��=,L=�=��=OE=��=?�=�9=�� =z� =�+ =h��<���<�>�<*��<���<X0�<��<��<{)�<�|�<���<�!�<�r�<|��<��<=]�<b��<��<�:�<"��<���<��<T�<ܘ�<��<� �<�c�<���<��<4%�<Ib�< ��<)��<
�<�;�<�i�<C��<ܺ�<���<���</�< 0�<ZD�<DU�<\b�<�k�<�p�<.q�<�l�<b�<Q�<�8�<��<���<P��<���<I@�<P��<b��<�8�<���<sY�<Z��<�V�<���<�2�<C��<���<�D�<v��<@ٻ<��<�S�<���<_��<ݲ<%��<��<3�<�E�<�T�<�_�<�g�<�m�<�q�<�t�<8v�<�w�<[x�<�x�<�x�<ox�<Tw�<.u�<�q�<.m�<�f�<_�<�U�<�J�<>�<Ca~<aDz<�&v<$r<��m<��i<�e<h�a<y]<T`Y<�HU<�2Q<zM<�I<b�D<�@<��<<&�8<��4<��0<|{,< j(<)[$<�O < I<�G<hL<�W<]k<+�<7�<� <G�;��;W�;���;-8�;��;N��;]w�;�Y�;�O�;�\�;]��;5��;,�;ޗ�;`3�;|��; у;��{;_�o;�d;huY;��N;D;g�9;ĥ/;��%;k?;p�;��	;� ;�|�:���:1C�:-V�:��:�:N�:(�:�l: �Q:4�7:�#:��:�w�9��90�n9R�9
{>8�9;�w��Vj�!a���sѹ= ���=�o�,��C�RY�go�sm��B�����Y͢�r���`O���ú��ͺT�غ�����~����N�y��GM���8�����"�3M(�a�-��2��8�i3=�J_B�(�G��L��Q��-W�Ir\���a��g�ul���q�b@w���|��
���s��1&���֋�j���v4��6⓻w���l?���  �  #�=rL=B�=��=.E=L�=ߒ=9=�� =�� =�* =���<���<�<�<!��<���<o.�<��<j��<(�<�{�<���<&!�<lr�<D��<��<�]�< ��<��<�;�<���<h��<}�<�U�<Ӛ�<��<�"�<de�<"��<���<f&�<Dc�<Ý�<���<L
�<�;�<�i�<���<��<���<s��<��<N.�<�B�<6S�<J`�<�i�<�n�<]o�<�j�<�`�<�O�<�7�<=�<��<��<���<�@�<���<1��<�9�<��<[�<��<pX�<���<�4�<\��<���<�F�<#��<�ڻ<�<�T�<h��<յ�<Kݲ<	��<[�<2�<E�<}S�<a^�<Uf�<�k�<�o�<jr�<2t�<ku�<]v�<�v�<'w�<�v�<v�<0t�<q�<�l�<�f�<_�<�U�<K�<�>�<@c~<�Fz<�)v<�r<j�m<��i<�e<X�a<�|]<�cY<LU<^5Q<�M<d
I<��D<��@<��<<��8<��4<�0<�y,<�g(<=X$<jL <@E<�C<H<�S<�f<1�<^�<�� <Q�;�|�;z�;E��;36�;���;+��;Vx�;�[�;;S�;�`�;���;ǣ;�#�;��;�:�;J��;G؃;�{;�p;d�d;m~Y;ףN;�D;9�9;9�/;W�%;�<;��;�	;r� ;dg�:��:�%�:|8�:R��:`��:�,�:F�:ǈl:�Q:ɒ7:��:W�:�C�9�t�9edn9��9A�>8vw:��a���i�1��ѹ���h�D{,��B���X�x�n�=Q��&)�������������D���ú3�ͺ��غd��˪�����W����hZ����3G�ί��#�^(�Q�-���2�"8�/?=��iB��G���L��Q��/W��r\�z�a��g�]nl���q�6w�t�|����u����k����ϋ��~���-��ܓ����Z;���  �  A�=H=f�=V�=�?=��=V�=�3=�� =� =w% =��<���<>1�<��<^��<6�<}n�<;��<�<�`�<���<U �<�N�<��<1��<�2�<|�<!��<�
�<�P�<���<s��<��<�^�<v��<��<� �<)_�<>��<^��<��<�G�<�{�<!��<"��<��<-�<�P�<mp�<}��<��<���<���<-��<���<A��<���<H��<��<3��<��<ƚ�<w�<�K�<��<���<6��<SF�<j��<b��<S#�<���<g5�<��<�&�<y��<��<{W�<
��<���<hJ�<N��<C̷<�<6�<bb�<��<ƪ�<�Ǭ<�ߪ<J��<*�<�<j�<�'�<�/�<_6�<�;�<z@�<�D�<�G�<�J�<GL�<M�<{L�<�J�<yG�<�B�<�<�<h5�<�,�<wF~<�1z<"v<�r<=�m<��i<��e<��a<R�]<�Y<�wU<ygQ<!XM<�II<�;E<'.A<	!=<39<;5<
�0<��,<��(<B�$<
� <S�<��< <Y<�0<�S	<>~<p�<d��;�V�;���;��;L9�;���;!��;d��;���;g��;�ų;���;*M�;��;WB�;.�;]��;?��;5��;�u;�Dj;�%_;�JT;رI;�X?;f?5;�a+;��!;�[;<0;�>;��:�:���:i�:a��:Ԁ�:ì�:|8�:XR~:��b:  H:ʰ-:��:���9��9�G�9��@9�ܾ8��w�&(����?�{⎹ƚ��칅�G�#���:�;�P�Mg�y}���˻��������������u��.g˺�aֺ�`�xg캲p���>����F���-:�r��@"�]l'��,�T2�7R7���<���A�G�WPL���Q�_�V�.\���a���f�wDl�u�q��w�{�|���������^g������ы�����'9��i쓻�����U���  �  !�=�G=R�=O�=�?=��=r�=�3=�� =� =�% =���<]��<�1�<��<���<��<�n�<���<s�<a�<3��<� �<�N�<+��<��<�2�<�{�<���<�
�<UP�<#��<��<!�<y^�<��<���<[ �<�^�<Û�<��<f�<OG�<�{�<���<.��<��<2-�<�P�<�p�<׌�<q��<>��<l��<���<,��<���<���<���<���<���<<��<
��<Sw�<�K�<��<���<��<(F�<(��<��<#�<>��<�4�<���<&�<��<���<W�<���<���<�I�<	��<�˷<��<�5�<5b�< ��<ߪ�<�Ǭ<(�<���<��<�<��<_(�<0�<�6�<0<�<A�<E�<qH�<K�<�L�<MM�<�L�<�J�<�G�<�B�<�<�<@5�<�,�<�E~<1z<;v<�r<]�m< �i<��e<�a<p�]<�Y<�vU<�fQ<�WM<)II<S;E<�-A<� =<b9<�5<z�0<�,<��(<�$<�� <O�<��<� <�<�1<�T	<F<g�<���;RX�;���;��;�9�;��;���;ש�;��;���;ų;?��;�K�;~��;�@�;��;���;ř�;���;�u;Aj;*#_;!IT;�I;�W?;5>5;ib+;g�!;H];2;
A;��:��:҉�:=p�:�Ĺ:��:o��:�A�:�`~:(�b:�H:[�-:��:���9d��9�N�9��@9���8\���c���?�*������� ���H�#���:��
Q�L[g���}�ɉ�PÔ�곟�������x���i˺�`ֺ�^��c��l��<����{B���[6���*"�-i'���,��2�`N7�}�<���A�WG��NL�6�Q���V�9.\�օa��f��Fl�_�q��w��|�I���R����h�����wӋ�\����:��&/����V���  �  Ǟ=�G=6�=J�=�?=�=��=4=D� =F� =S& =��<���<N3�<x��<���< �<Np�<���<~�<�a�<��<�<=O�<J��<���<e2�<o{�<"��<�	�<BO�<���<���<��<]�<���<>��<��<�]�<���<%��<��<�F�<O{�<Ǭ�<>��<!�<�-�<cQ�<�q�<ލ�<���<���<���<O��<���<��<��<���<���<���<?��<ܛ�<�w�<L�<��<���<Δ�<�E�<���<=��<"�<��<�3�<��<�$�<j��< ��<~U�<(��<>��<�H�<��<˷<C�<�5�<b�<)��<��<+Ȭ<��<r��<��<��<4 �<�)�<�1�<48�<�=�<�B�<hF�<�I�<L�<�M�<N�<VM�<@K�<�G�<�B�<y<�<�4�<�+�<gD~</z<�v<Qr<��m<9�i<}�e<�a<��]<r�Y<�tU<�dQ<�UM<�GI<x:E<V-A<� =<�9<&	5<��0<��,<��(<4�$<�� <��<��<V<<�4<�W	<�<�<u��;`\�;���;���;3;�;���;���;G��;���;ӣ�;³;>��;NG�;y��;D;�;�;ު�;?��;I��;��u;�8j;a_;(CT;��I;�U?;=5;=c+;�!;�`;p7;�G;�"�:s'�:��:��:޹:��:I˛:i[�:}�~:�c:L1H:��-:F:j#�9���9�Z�9��@9���8Eϕ�O����@�y,��� ��m�i@�!$���:��9Q�ӈg�b�}��ۉ��Ԕ�8���$���.����{��Wk˺_ֺ.[Ẍ[�b���4����!9�^���+���u�!�1\'���,�9�1�-D7��<���A�:G��IL�K�Q�f�V�8.\�x�a��f��Kl���q�F"w��|�H ����n���$��*ً�򌎻�?����%���Z���  �  E�=[G=�=C�=@=P�=0�=�4=� =%� =O' =%��<��<�5�<؃�<���<T"�<yr�<���<5�<hc�<��<��<�O�<y��<���<�1�<�z�<��<f�<�M�<��<���<��<�Z�<J��<��<��<�[�<��<���<Y�<�E�<�z�<���<C��<��<W.�<dR�<�r�<x��<N��<���<���<y��<��<s��<B��<9��<���<y��<ֹ�<��<�x�<�L�<�<���<��<E�<���<��<j �<5��<�1�<ȭ�<?"�<��<���<8S�<骾<$��<�F�<��<�ɷ<K�<�4�<�a�<1��<i��<�Ȭ<��<���<%�<y�<M"�<�+�<�3�<�:�<@�<�D�<�H�<�K�<�M�<1O�<YO�<KN�<�K�<H�<�B�<%<�<-4�<�*�<�A~<�+z<Sv<(�q<0�m<��i<�e<{�a<1�]<4�Y<�pU<caQ<SM<�EI<�8E<|,A<� =<9<L
5<k 1<��,<��(<��$<�� <��<Y�<	<<�9<c\	<��<�<���;�b�;���;d��;�=�;��;���;ҧ�;���;�;���;V�;
@�;���; 3�;�ڒ;i��;Ջ�;��;�u;;+j;�_;�9T;ˤI;�P?;�;5;�c+;��!;.g;�?;�R;=�:�D�:x��:ة�:j�:�Ū:3�:�~�:e�~:�Tc:LlH:�.:�.:�f�9D'�9-v�9͝@9�R�8s����¸��@����bn�����Ą�Y]$��;�ĀQ���g���}�B�����؟�5������������m˺�\ֺOSẠN캝P���)����)�4����D����!��I'���,�5�1�347��x<���A�X�F�EBL�3�Q��V�o.\�B�a���f��Sl���q��.w���|���������w���-��#⋻����;H��!���f����_���  �  ��=�F=��=/�=*@=��=��=|5=�� =M� =�( =��<��<�8�<���<���<T%�<'u�<C��<l�<2e�<}��<��<pP�<���<���<<1�<�y�<���<{�<�K�<���<���<��<�W�<:��<��<�<�X�<���<���<��<�D�<�y�<��<8��<��<)/�<�S�<ft�<y��<���<��<���<���<1��<���<I��<��<_��<���<Ի�<���< z�<�M�<��<���<��<!D�<5��<.��<C�<˪�<�.�<��<�<ˋ�<Z��<P�<	��<q��<�D�<`��<6ȷ<�<�3�<Qa�<2��<竮<�ɬ<�<g��<:
�<��<�$�<�.�<�6�<�=�<3C�<�G�<K�<AN�<FP�<(Q�<�P�<|O�<�L�<|H�<�B�<�;�<;3�<�)�<3>~<�'z<�v<��q<{�m<��i<Ӵe<>�a<Z�]<�{Y<�kU<]Q<WOM<�BI<�6E<A+A<; =<�9<�5<�1<�,<[�(<p�$<�� <7�<� <m<y$<@<�b	<:�<3�<>��;Pj�;\��;$��;$A�;���;c��;ȥ�;��;Қ�;���;U�;�6�;f��;�'�;�Β;���;F��;���;^vu;�j;s_;X-T;�I;�J?;�85;<d+;�!;Vn;WJ;`; ^�:Cl�:���:���:�2�:]��:�#�:)��:�1:{�c:h�H:	U.:�c:,��9�^�9l��9ݡ@9���87o�ĸ�kA����G���ԑ������$�)j;���Q�,h��J~��#���������ժ�ᱵ�j���Kr˺XZֺ<I�1?��9�������a�%�����n���!��0'���,���1�8 7��e<�.�A���F�9L�	�Q���V�p/\�W�a���f�%^l���q�=?w���|����˃�̓���9��k
����R�����Ŵ���f���  �  Ĝ=HF=f�=�=S@=�=j�=_6=� =�� =* =��<p��<C<�<���<j��<�(�<Rx�<.��<��<Lg�<*��<(�<Q�<��<K��<z0�<Ex�<վ�<`�<�H�<���<���<?�<JT�<Õ�<���<��<�U�<֓�<B��<�
�<C�<�x�<���</��<y�<0�<U�<Uv�<���<k��<*��<��<���<���<��<���<O��<i��<���<��<���<�{�<tN�<��<���<]��<C�<���<��<��<ߧ�<�+�<b��<j�<#��<���<mL�<���<?��<�A�<��<-Ʒ<��<�2�<�`�<-��<a��<�ʬ<��<Y��<��<��<�'�<2�<r:�<3A�<�F�<3K�<�N�<KQ�<�R�<iS�<�R�<�P�<�M�<�H�<�B�<;�<12�<(�<9:~<�"z<�
v<��q<��m<��i<­e<T�a<��]<huY<�eU<�WQ<#KM<L?I<S4E<�)A<�=<=9<I5<E1<��,<��(<��$<�� <��<�<�<�+<sG<�i	<��<^�<���;ps�;���;���;�D�;$��;���;|��;���;r��;ﭳ;�߬;�+�;Q��; �;���;r��;.s�;��;	_u;�j;��^;�T;��I;�C?;V55;�d+;��!;�v;�V;p;σ�:���:��:F�:Zk�:�1�:]�:��:��:Qd:I:��.:[�:��9���9���9W�@9}w�8����{Ÿ�`B�Ꝑ�Ŭ��%S�6E�Q+%�7�;�
QR�A�h�ݱ~�S��`<��\��󪺊ǵ�7���Qx˺�Wֺ?�-캵��;���]���u�R��$R���!�G'�Mk,�(�1�7��P<�q�A�1�F��-L�1~Q���V��0\�S�a�.�f�kl���q��Rw�T�|�|��5ك�f����G�����o���P_��L��׾��o���  �  ޛ=�E=�=��=z@=}�=�=L7==� =�� =�+ =���<��<@�<X��<1��<I,�<�{�<6��<��<�i�<��<o�<�Q�<��<���<�/�<�v�<���<�<F�<���<P��<��<P�<��<���<+�<�R�<ސ�<���<��<lA�<�w�<���<+��<��<!1�<�V�<Xx�<D��<=��<m��<���<���<}��<���<q��<���<���<^��<���<���<}�<qO�<Y�<���<���<�A�<���<߄�<�<���</(�<���<��<��<���<�H�<⠾<��<�>�<a��<	ķ<���<�1�<.`�<"��<٬�<�ˬ<#�<p��<�<��<E+�<�5�<,>�<�D�<�J�<�N�<=R�<�T�<�U�<�U�<�T�<bR�<�N�<LI�<�B�<a:�<�0�<`&�<�5~<�z<�v<��q<i�m<�i<�e<��a<]<�nY<�_U<ARQ<vFM<�;I<�1E<(A<9=<�9<�5<�1<M-<��(<$�$<� <�<<�<�3<LO<*q	<�<��<6�;P}�;��;���;7H�;���;d��;���;��;���;I��;լ;��;H��;�;:��;�z�;e�;4r�;>Fu;�i;?�^;T;��I;�;?;�15;qe+;��!;�;�c;ـ;E��:��:&Q�:�F�:t��:[o�:���:%�:��:�vd:�pI:��.:��:U��9���9ݑ9��@9��8�8��
ǸNdC��?���h��t ﹘����%�qS<��R��i�� �'���&j���@������޵������~˺�Uֺ�4�i������ �=q�����Z�n�� 4���!���&��M,��1�~�6��:<�݅A���F��"L�	wQ�5�V��1\�2�a�g��xl�?�q�jhw���|��,���烻T���*W��������l��}���ɖ�x���  �  ��=�D=��=ؗ=�@=��=��=58=a� =R� =%- =���<���<�C�<5��<���<�/�<�<8��<6�<�k�<���<��<�R�<,��<���<�.�<mu�<��<���<PC�<J��<���<�
�<�L�<��<)��<��<?O�<��<��<x�<�?�<wv�<Y��<��<T�<2�<X�<Hz�<���<��<���<	��<J��<G��<���<��<L��<���<6��<���<���<x~�<^P�<��<R��<���<�@�<��<���<S�<���<�$�<ϟ�<��<��<���<�D�<��<c�<�;�<���<���<��<�0�<�_�<���<N��<�̬<��<m��<��<h!�<v.�<+9�<�A�<�H�<UN�<�R�<�U�<�W�<�X�<DX�<�V�<�S�<|O�<�I�<dB�<�9�<�/�<�$�<F1~<Iz<��u<��q<�m<s�i<?�e<��a<�w]<lgY<:YU<�LQ<�AM<�7I<�.E<e&A<�=<9<n5<�
1<�-<1)<�%<V!<�<�<^&<�;<W<�x	<�<,�<��;Ć�;3�;>��;�K�;� �;���;���;��;���;%��;�ʬ;��;�y�;���;���;l�;�V�;cd�;V,u;��i;��^;��S;qxI;3?;y-5;Pe+;�!;*�;4p; �;Z��:��:S��:v�:��:��:�؜:`�:�?�:L�d:��I::C/:�':E��9H*�9:��9t�@9fj�8D)]�C�ȸtsD�䑹�"����`)�X&���<�)ES�W�i����i���3���/i���1����������O�˺Uֺ�*��_����� �_\�����@����u��y!���&�s0,���1���6��$<�<sA��F��L�pQ���V�z3\��a�g��l��r��}w��|��:��F���w���Pf��6���ˎ��z���'��Ԗ�|����  �  �=PD=;�=��=�@=?�=X�=9=g� =�� =�. = ��< ��<;G�<���<Q��<=3�<%��<��<��<�m�<3��<��<S�<K��<2��<�-�<t�<(��<Q��<�@�<B��<���<s�<I�<���<���<E�<L�<��<���<k�<$>�<[u�<���<���<��<�2�<zY�<|�<ښ�<���<���<B��<���<���<��<p��<���<���<���< ��<Q��<��<#Q�<�<"��<H��<T?�<Q��<]��<��<���<M!�<V��<��<;|�<���<�@�<���<�<�8�<(�<���<r��<�/�<�^�<∰<���<�ͬ<�<D �<��<$�<t1�<o<�<2E�<@L�<�Q�<�U�<�X�<�Z�<*[�<dZ�<uX�<U�<FP�<�I�<4B�<9�<�.�<�"�<-~<=z<��u<��q<P�m<4�i<��e<��a<�p]<�`Y<"SU<zGQ<=M< 4I<,E<�$A<�=<�9<�5<�1<S	-<T)<�%<:!<8<s<a-<�B<^<�	<��<-�<�;m��;E�;&��;O�;,�;���;���;���;��;퓳;���;I�;�m�;��;���;i^�;I�;�W�;Pu;��i;M�^;/�S;[lI;+?;^)5;e+;��!;a�;�{;Z�;	��:�!�:Ҵ�:	��:�::�:��:R��:pt�:>e:�%J:�/:e:�C�98c�9��9��@9ڻ8�m~��5ʸ$vE�B{��r���S��ݑ�|�&�m?=��S�n�i����HꊺW�����kP��c������˺/Tֺ�!�I�������� �xI�X�� (� �� ���]!�F�&�l,�3k1�v�6��<��bA��F��L�jQ���V�J5\���a�Ug���l��r�w��}�9G�����̽���t���(��,َ�b����3���ޖ�(����  �  S�=�C=��=��=�@=��=ۑ=�9=R� =�� =�/ =ƭ�<��<NJ�<���<Z��<6�<Ä�<f��<�!�<wo�<}��<��<�S�<g��<���<�,�<�r�<���<[��<G>�<���<���<e�<�E�<f��<���<L	�<~I�<���<���<��<�<�<kt�<��<���<	�<�3�<�Z�<�}�<˜�<��<��<���<���<���< �<g �</��<;��<��<��<ʧ�<݀�<�Q�<H�<���<���<R>�<���<�~�<��<��<��<6��<��<�x�<���<�=�<���<d�<6�<�|�<뽷<��<�.�<N^�<͈�<��<bά<,�<��<��<W&�<�3�<'?�<.H�<IO�<�T�<�X�<�[�<]�<R]�<P\�<�Y�<.V�<�P�<;J�<B�<Z8�<{-�<z!�<o)~<�z<��u<+�q<>�m<��i<��e<r|a<�j]<M[Y<NU<�BQ<A9M<�0I<�)E<2#A<9=<�9<�5<�1<-<)<.%<1!<�<_#<�3<4I<fd<��	<�<'�<��;��;�;���;�Q�;D�;���;y��;�~�;Wz�;���;ݷ�;���;�b�;.�;��;oR�;8=�;eL�;[ u; �i;��^;$�S;bI;K$?;6%5;�d+;�!;�;�;��;!�:�E�:���:���:EJ�:H�:�A�:�ǎ:��:Ïe:�mJ:��/:�:_��9p��9�0�9�@9�M�82����˸�LF�� ��Tr¹'c�!����&���=�VT�TVj�+������蕺����j���!�������˺(Sֺ�������� �=9���^��|����sE!���&��+��U1���6���;�mSA���F�:L��dQ���V�&7\�2�a��"g���l�(!r���w�,%}�	R�����ʆ�/����4��K去h����=���疻�����  �  ��=TC=��=o�=�@=��=?�=@:=� =n� =�0 =گ�<+��<�L�<��<���<18�<ц�<3��<>#�<�p�<p��<X	�<�S�<k��<x��<P,�<�q�<R��<���<�<�<�~�<x��<1�<�C�<
��<Q��<�<\G�<���<���<S�<�;�<�s�<���<���<0	�<@4�<g[�<�~�<G��<���<���<��<���<���<C�<��<G��<4��<���<���<��<���<eR�<f�<���<��<o=�<���<}�<��<��<Q�<ϖ�<6
�<kv�<��<N;�<+��<4�<#4�<A{�<���<���<�-�<�]�<���<0��<�ά<�<�<;�<(�<�5�<AA�<]J�<zQ�<W�<[�<�]�<�^�<�^�<�]�<[�<W�<pQ�<ZJ�<�A�<�7�<�,�<V �<�&~<Sz<��u<��q<��m<i�i<ϋe<�wa<f]<�VY<JU<5?Q<<6M<�.I<�'E<�!A<�=<�9<�5<�1<$-<�)<a%<!<�<�'<U8<�M<
i<
�	<X�<��<~&�;Ȝ�;X �;��;^S�;��;��;P��;�{�;�u�;��;9��;7��;KZ�;�ݘ;6��;fI�;�4�;�C�;�t;Ġi;#�^;��S; ZI;s?;�!5;Kd+;��!;��;C�;I�;�1�:{`�:���:��:�l�::�:be�:Y�:b:��e:D�J:��/:>�:���97��9�=�9��@9ݺ8Ӱ���̸��F��j��}�¹���8�2'���=��eT�`�j�ZO���3������Ơ��~���1��������˺LSֺr����5���I� ��,�Ę���k�C���3!���&���+�#E1�S�6��;��GA�7�F���K�PaQ���V��8\���a�~)g�Ʃl��,r�i�w��4}��Z�����$ӆ�����>��3?����E���y����  �  ^�=
C=n�=]�=�@=��=t�=�:=n� =� =R1 =%��<���<�M�<y��<��<�9�<��<Q��<0$�<�q�<��<�	�< T�<e��<P��<�+�<Bq�<���<���<o;�<s}�<-��<� �<B�<q��<���<��<F�<���<���<n �<�:�<s�<p��<���<O	�<w4�<�[�<��<��<���<)��<b��<*��<b��<��<��<���<`��<���<R��<���<4��<�R�<��<���<ӏ�<�<�<���<&|�<��<՘�<��<n��<��<�t�<Y��<�9�<ʒ�<��<�2�<#z�<���<9��<7-�<�]�<���<Q��<>Ϭ<��<��<�< )�<,7�<�B�<�K�<�R�<vX�<h\�<�^�<'`�<�_�<�^�<�[�<~W�<�Q�<tJ�<�A�<�7�<,�<��<�$~<8	z<�u<�q<�m<�i<��e<zta<(c]<TY<�GU<=Q<<4M<�,I<�&E<T!A<\=<�9<!5<S1<�-<�)<l%<Y!<�<�*<F;<�P<l<��	<�<Y�<�*�;F��;P#�;���;�T�;�;���;��;gy�;�r�;D��;:��;]�;eU�;ؘ;�{�;BC�;�.�;�>�;��t;��i;E�^;'�S;�TI;�?;� 5;�c+;	�!;��;ǐ;ʼ;d?�:�r�:<�:'�:ԃ�:�Q�:}�:g�:�؀:�e:�J:�0:��:���9���9�G�9k�@9���8Y2��"@͸�eG�����A0ù�>��a�se'�@">���T���j��c��vH�����aנ������;��b�����˺/Tֺ[�������� ��%�ۏ�G���`�����'!�-�&���+��:1��6���;�bAA�E�F��K��_Q�O�V��9\���a��-g�c�l�>4r�Թw�]>}�`��6���ن������D���󎻄����J���Y����  �  B�=�B=\�=Q�=�@=��=��=�:=�� =$� =�1 =���<���<`N�<��<i��<:�<w��<���<�$�<�q�<Z��<�	�<IT�<e��<8��<�+�<q�<R��<t��<	;�<�|�<���< �<�A�<+��<"��<>�<�E�<!��<l��< �<�:�<�r�<Q��<~��<v	�<�4�<'\�<��<\��<'��<���<���<���<���<,�<W�<��<���<9��<���<��<k��<�R�<��<���<���<�<�<���<�{�<>�<`��<\�<��<��<jt�<���<9�<P��<H�<�2�<�y�<U��<���<-�<v]�<���<t��<^Ϭ<��<�<l�<�)�<�7�<C�<,L�<oS�<�X�<�\�<__�<�`�<l`�<�^�<\�<�W�<�Q�<�J�<�A�<x7�<�+�<n�<$~<vz<��u<�q<�m<�i<%�e<�sa<b]<SY<�FU<9<Q<�3M<�,I<<&E<!A<(=<9<r5<�1<-<�)<B%<8!<c<�+<<<�Q<�l<�	<Ѵ<O�<,�;U��;k$�;`��;?U�;*�;}��;���;�x�;/r�;�;���;��;�S�;�՘;�z�;@B�;a,�;�<�;��t;��i;w�^;��S;-SI;(?;�5;Nc+;`�!;_�;��;ݾ;�C�:Wz�:[�:��:؊�:�X�:���:�:�ހ:)f:��J:�0:�:i��9���9uR�9�z@9���8�l��7{͸ފG��ē��Kù�_�p��w'�E+>�t�T�z�j�k��mP��`��ݠ�����m?��.����˺�Tֺ��q��N����� ��"���	��M]���� $!��&� �+�F71�ӎ6�4�;��?A�T�F���K�E^Q�x�V��:\���a��/g��l��6r�ܼw�B}�b��@ ���ۆ�葉�SF�� ���z���cL�����������  �  ^�=
C=n�=]�=�@=��=t�=�:=n� =� =R1 =%��<���<�M�<y��<��<�9�<��<Q��<0$�<�q�<��<�	�< T�<e��<P��<�+�<Bq�<���<���<o;�<s}�<-��<� �<B�<q��<���<��<F�<���<���<n �<�:�<s�<p��<���<O	�<w4�<�[�<��<��<���<)��<b��<*��<b��<��<��<���<`��<���<R��<���<4��<�R�<��<���<ӏ�<�<�<���<&|�<��<՘�<��<n��<��<�t�<Y��<�9�<ʒ�<��<�2�<#z�<���<9��<7-�<�]�<���<Q��<>Ϭ<��<��<�< )�<,7�<�B�<�K�<�R�<vX�<h\�<�^�<'`�<�_�<�^�<�[�<~W�<�Q�<tJ�<�A�<�7�<,�<��<�$~<8	z<�u<�q<�m<�i<��e<zta<(c]<TY<�GU<=Q<<4M<�,I<�&E<T!A<\=<�9<!5<S1<�-<�)<l%<Y!<�<�*<F;<�P<l<��	<�<Y�<�*�;F��;P#�;���;�T�;�;���;��;gy�;�r�;C��;:��;]�;eU�;ؘ;�{�;BC�;�.�;�>�;��t;��i;E�^;&�S;�TI;�?;� 5;�c+;	�!;��;ǐ;ʼ;d?�:�r�:<�:'�:ԃ�:�Q�:}�:g�:�؀:�e:�J:�0:��:���9���9�G�9k�@9���8Y2��"@͸�eG�����A0ù�>��a�se'�@">���T���j��c��vH�����aנ������;��b�����˺/Tֺ[�������� ��%�ۏ�G���`�����'!�-�&���+��:1��6���;�bAA�E�F��K��_Q�O�V��9\���a��-g�c�l�>4r�Թw�]>}�`��6���ن������D���󎻄����J���Y����  �  ��=TC=��=o�=�@=��=?�=@:=� =n� =�0 =گ�<+��<�L�<��<���<18�<ц�<3��<>#�<�p�<p��<X	�<�S�<k��<x��<P,�<�q�<R��<���<�<�<�~�<x��<1�<�C�<
��<Q��<�<\G�<���<���<S�<�;�<�s�<���<���<0	�<@4�<g[�<�~�<G��<���<���<��<���<���<C�<��<G��<4��<���<���<��<���<eR�<f�<���<��<o=�<���<}�<��<	��<R�<ϖ�<6
�<kv�<��<N;�<+��<4�<#4�<A{�<���<���<�-�<�]�<���<0��<�ά<�<�<;�<(�<�5�<AA�<]J�<zQ�<W�<[�<�]�<�^�<�^�<�]�<[�<W�<pQ�<ZJ�<�A�<�7�<�,�<U �<�&~<Sz<��u<��q<��m<i�i<ϋe<�wa<f]<�VY<JU<5?Q<<6M<�.I<�'E<�!A<�=<�9<�5<�1<$-<�)<a%<!<�<�'<U8<�M<
i<
�	<X�<��<~&�;Ȝ�;X �;��;]S�;��;��;P��;�{�;�u�;��;8��;7��;KZ�;�ݘ;5��;eI�;�4�;�C�;�t;ài;#�^;��S;�YI;r?;�!5;Kd+;��!;��;B�;H�;�1�:{`�:���:��:�l�::�:be�:Y�:b:��e:D�J:��/:>�:���97��9�=�9��@9ݺ8Ӱ���̸��F��j��}�¹���8�2'���=��eT�`�j�ZO���3������Ơ��~���1��������˺LSֺr����5���I� ��,�Ę���k�C���3!���&���+�#E1�S�6��;��GA�7�F���K�PaQ���V��8\���a�~)g�Ʃl��,r�i�w��4}��Z�����$ӆ�����>��3?����E���y����  �  S�=�C=��=��=�@=��=ۑ=�9=R� =�� =�/ =ƭ�<��<NJ�<���<Z��<6�<Ä�<f��<�!�<wo�<}��<��<�S�<g��<���<�,�<�r�<���<[��<G>�<���<���<e�<�E�<f��<���<L	�<~I�<���<���<��<�<�<kt�<��<���<	�<�3�<�Z�<�}�<˜�<��<��<���<���<���< �<g �</��<;��<��<��<ʧ�<݀�<�Q�<H�<���<���<R>�<���<�~�<��<��<��<6��<��<�x�<���<�=�<���<e�<6�<�|�<콷<��<�.�<N^�<͈�<��<bά<,�<��<��<W&�<�3�<'?�<.H�<IO�<�T�<�X�<�[�<]�<R]�<O\�<�Y�<.V�<�P�<;J�<B�<Z8�<{-�<z!�<n)~<�z<��u<+�q<>�m<��i<��e<r|a<�j]<N[Y<NU<�BQ<A9M<�0I<�)E<2#A<9=<�9<�5<�1<-<)<.%<1!<�<_#<�3<4I<fd<��	<�<'�<��;��;�;���;�Q�;C�;���;y��;�~�;Vz�;���;ݷ�;���;�b�;.�;��;nR�;8=�;eL�;Z u;�i;��^;$�S;bI;K$?;6%5;�d+;�!;�;�;��;!�:�E�:���:���:EJ�:H�:�A�:�ǎ:��:Ïe:�mJ:��/:�:_��9p��9�0�9�@9�M�82����˸�LF�� ��Tr¹'c�!����&���=�VT�TVj�+������蕺����j���!�������˺(Sֺ�������� �=9���^��|����sE!���&��+��U1���6���;�mSA���F�:L��dQ���V�&7\�2�a��"g���l�(!r���w�,%}�	R�����ʆ�/����4��K去h����=���疻�����  �  �=PD=;�=��=�@=?�=X�=9=g� =�� =�. = ��< ��<;G�<���<Q��<=3�<%��<��<��<�m�<3��<��<S�<K��<2��<�-�<t�<(��<Q��<�@�<B��<���<s�<I�<���<���<E�<L�<��<���<k�<$>�<[u�<���<���<��<�2�<zY�<|�<ښ�<���<���<B��<���<���<��<p��<���<���<���< ��<Q��<��<#Q�<�<"��<H��<T?�<Q��<]��<��<���<M!�<V��<��<;|�<���<�@�<���<�<�8�<)�<���<s��<�/�<�^�<∰<���<�ͬ<�<D �<��<$�<t1�<o<�<2E�<@L�<�Q�<�U�<�X�<�Z�<)[�<cZ�<uX�<U�<EP�<�I�<4B�<9�<�.�<�"�<-~<<z<��u<��q<P�m<4�i<��e<��a<�p]<�`Y<"SU<zGQ<=M<!4I<,E<�$A<�=<�9<�5<�1<S	-<T)<�%<:!<9<s<a-<�B<^<�	<��<,�<�;l��;E�;%��;O�;+�;���;���;���;��;쓳;���;H�;�m�;��;���;i^�;I�;�W�;Pu;��i;M�^;/�S;[lI;+?;])5;e+;��!;a�;�{;Z�;	��:�!�:Ҵ�:	��:�::�:��:R��:pt�:>e:�%J:�/:e:�C�98c�9��9��@9ڻ8�m~��5ʸ$vE�B{��r���S��ݑ�|�&�m?=��S�n�i����HꊺW�����kP��c������˺/Tֺ�!�I�������� �xI�X�� (� �� ���]!�F�&�l,�3k1�v�6��<��bA��F��L�jQ���V�J5\���a�Ug���l��r�w��}�9G�����̽���t���(��,َ�b����3���ޖ�(����  �  ��=�D=��=ؗ=�@=��=��=58=a� =R� =%- =���<���<�C�<5��<���<�/�<�<8��<6�<�k�<���<��<�R�<,��<���<�.�<mu�<��<���<PC�<J��<���<�
�<�L�<��<)��<��<?O�<��<��<x�<�?�<wv�<Y��<��<T�<2�<X�<Hz�<���<��<���<	��<J��<G��<���<��<L��<���<6��<���<���<x~�<^P�<��<R��<���<�@�<��<���<T�<���<�$�<ϟ�<��<��<���<�D�<��<c�<�;�<���<���<��<�0�<�_�<���<N��<�̬<��<m��<��<h!�<v.�<+9�<�A�<�H�<UN�<�R�<�U�<�W�<�X�<DX�<�V�<�S�<|O�<�I�<dB�<�9�<�/�<�$�<F1~<Iz<��u<��q<�m<s�i<?�e<��a<�w]<lgY<:YU<�LQ<�AM<�7I<�.E<e&A<�=<9<o5<�
1<�-<2)<�%<V!<�<�<^&<�;<W<�x	<�<,�<��;Æ�;2�;=��;�K�;� �;���;���;��;���;$��;�ʬ;��;�y�;���;���;l�;�V�;bd�;U,u;��i;��^;��S;qxI;3?;y-5;Pe+;�!;)�;4p; �;Z��:��:S��:v�:��:��:�؜:`�:�?�:L�d:��I::C/:�':E��9H*�9:��9t�@9fj�8E)]�C�ȸtsD�䑹�"����`)�X&���<�)ES�W�i����i���3���/i���1����������O�˺Uֺ�*��_����� �_\�����@����u��y!���&�s0,���1���6��$<�<sA��F��L�pQ���V�z3\��a�g��l��r��}w��|��:��F���w���Pf��6���ˎ��z���'��Ԗ�|����  �  ޛ=�E=�=��=z@=}�=�=L7==� =�� =�+ =���<��<@�<X��<1��<I,�<�{�<6��<��<�i�<��<o�<�Q�<��<���<�/�<�v�<���<�<F�<���<P��<��<P�<��<���<+�<�R�<ސ�<���<��<lA�<�w�<���<+��<��<!1�<�V�<Xx�<D��<=��<m��<���<���<}��<���<q��<���<���<^��<���<���<}�<qO�<Y�<���<���<�A�<���<߄�<�<���</(�<���<��<��<���<�H�<⠾<��<�>�<a��<	ķ<���<�1�<.`�<"��<ڬ�<�ˬ<#�<p��<�<��<F+�<�5�<,>�<�D�<�J�<�N�<=R�<�T�<�U�<�U�<�T�<bR�<�N�<LI�<�B�<a:�<�0�<`&�<�5~<�z<�v<��q<i�m<�i<�e<��a<]<�nY<�_U<ARQ<vFM<�;I<�1E<(A<9=<�9<�5<�1<M-<��(<%�$<� <�<<�<�3<LO<*q	<�<��<6�;O}�;��;���;6H�;���;c��;���;��;���;H��;լ;��;G��;�;:��;�z�;e�;3r�;=Fu;�i;>�^;T;��I;�;?;�15;pe+;��!;�;�c;ـ;E��:��:&Q�:�F�:t��:[o�:���:%�:��:�vd:�pI:��.:��:U��9���9ݑ9��@9��8�8��
ǸNdC��?���h��t ﹘����%�qS<��R��i�� �'���&j���@������޵������~˺�Uֺ�4�i������ �=q�����Z�n�� 4���!���&��M,��1�~�6��:<�݅A���F��"L�	wQ�5�V��1\�2�a�g��xl�?�q�jhw���|��,���烻T���*W��������l��}���ɖ�x���  �  Ĝ=HF=f�=�=S@=�=j�=_6=� =�� =* =��<p��<C<�<���<j��<�(�<Rx�<.��<��<Lg�<*��<(�<Q�<��<K��<z0�<Ex�<վ�<`�<�H�<���<���<?�<JT�<Õ�<���<��<�U�<֓�<B��<�
�<C�<�x�<���</��<y�<0�<U�<Uv�<���<k��<*��<��<���<���<��<���<O��<i��<���<��<���<�{�<tN�<��<���<]��<C�<���<��<��<ߧ�<�+�<b��<k�<#��<���<mL�<���<@��<�A�<��<-Ʒ<��<�2�<�`�<-��<a��<�ʬ<��<Y��<��<��<�'�<2�<r:�<3A�<�F�<3K�<�N�<KQ�<�R�<iS�<�R�<�P�<�M�<�H�<�B�<;�<02�<(�<8:~<�"z<�
v<��q<��m<��i<­e<T�a<��]<huY<�eU<�WQ<#KM<L?I<S4E<�)A<�=<=9<I5<F1<��,<��(<��$<�� <��<�<�<�+<sG<�i	<��<^�<���;os�;���;���;�D�;#��;���;{��;���;r��;;�߬;�+�;P��;��;���;r��;-s�;��;_u;�j;��^;�T;��I;�C?;V55;�d+;��!;�v;�V;p;΃�:���:��:F�:Zk�:�1�:]�:��:��:Qd:I:��.:[�:��9���9���9W�@9}w�8����{Ÿ�`B�Ꝑ�Ŭ��%S�6E�Q+%�7�;�
QR�A�h�ݱ~�S��`<��\��󪺊ǵ�7���Qx˺�Wֺ?�-캵��;���]���u�R��$R���!�G'�Mk,�(�1�7��P<�q�A�1�F��-L�1~Q���V��0\�S�a�.�f�kl���q��Rw�T�|�|��5ك�f����G�����o���P_��L��׾��o���  �  ��=�F=��=/�=*@=��=��=|5=�� =M� =�( =��<��<�8�<���<���<T%�<'u�<C��<l�<2e�<}��<��<pP�<���<���<<1�<�y�<���<{�<�K�<���<���<��<�W�<:��<��<�<�X�<���<���<��<�D�<�y�<��<8��<��<)/�<�S�<ft�<y��<���<��<���<���<1��<���<I��<��<_��<���<Ի�<���< z�<�M�<��<���<��<!D�<5��<.��<C�<˪�<�.�<��<�<ˋ�<Z��<P�<	��<q��<�D�<`��<6ȷ<�<�3�<Qa�<3��<竮<�ɬ<�<g��<:
�<��<�$�<�.�<�6�<�=�<3C�<�G�<K�<AN�<FP�<(Q�<�P�<|O�<�L�<|H�<�B�<�;�<;3�<�)�<3>~<�'z<�v<��q<{�m<��i<Ӵe<>�a<Z�]<�{Y<�kU<]Q<WOM<�BI<�6E<A+A<; =<�9<�5<�1<�,<[�(<p�$<�� <8�<� <m<y$<@<�b	<:�<2�<>��;Pj�;[��;#��;#A�;���;c��;ǥ�;��;њ�;���;T�;�6�;f��;�'�;�Β;���;E��;���;]vu;�j;r_;X-T;�I;�J?;�85;<d+;�!;Vn;VJ;`; ^�:Cl�:���:���:�2�:]��:�#�:)��:�1:{�c:h�H:	U.:�c:,��9�^�9l��9ݡ@9���88o�ĸ�kA����G���ԑ������$�)j;���Q�,h��J~��#���������ժ�ᱵ�j���Kr˺XZֺ<I�1?��9�������a�%�����n���!��0'���,���1�8 7��e<�.�A���F�9L�	�Q���V�p/\�W�a���f�%^l���q�=?w���|����˃�̓���9��k
����R�����Ŵ���f���  �  E�=[G=�=C�=@=P�=0�=�4=� =%� =O' =%��<��<�5�<؃�<���<T"�<yr�<���<5�<hc�<��<��<�O�<y��<���<�1�<�z�<��<f�<�M�<��<���<��<�Z�<J��<��<��<�[�<��<���<Y�<�E�<�z�<���<C��<��<W.�<dR�<�r�<x��<N��<���<���<y��<��<s��<B��<9��<���<y��<ֹ�<��<�x�<�L�<�<���<��<E�<���<��<k �<5��<�1�<ȭ�<@"�<��<���<8S�<骾<%��<�F�<���<�ɷ<L�<�4�<�a�<1��<i��<�Ȭ<��<���<&�<y�<M"�<�+�<�3�<�:�<@�<�D�<�H�<�K�<�M�<1O�<YO�<KN�<�K�<H�<�B�<%<�<,4�<�*�<�A~<�+z<Sv<(�q<0�m<��i<�e<{�a<1�]<4�Y<�pU<caQ<SM<�EI<�8E<|,A<� =<9<M
5<k 1<��,<��(<��$<�� <��<Y�<	<<�9<c\	<��<�<���;�b�;���;c��;�=�;��;���;ҧ�;���;�;���;U�;	@�;���;3�;�ڒ;i��;ԋ�;��;�u;;+j;�_;�9T;ˤI;�P?;�;5;�c+;��!;.g;�?;�R;=�:�D�:x��:ة�:j�:�Ū:3�:�~�:e�~:�Tc:LlH:�.:�.:�f�9D'�9-v�9͝@9�R�8s����¸��@����bn�����Ą�Y]$��;�ĀQ���g���}�B�����؟�5������������m˺�\ֺOSẠN캝P���)����)�4����D����!��I'���,�5�1�347��x<���A�X�F�EBL�3�Q��V�o.\�B�a���f��Sl���q��.w���|���������w���-��#⋻����;H��!���f����_���  �  Ǟ=�G=6�=J�=�?=�=��=4=D� =F� =S& =��<���<N3�<x��<���< �<Np�<���<~�<�a�<��<�<=O�<J��<���<e2�<o{�<"��<�	�<BO�<���<���<��<]�<���<>��<��<�]�<���<%��<��<�F�<O{�<Ǭ�<>��<!�<�-�<cQ�<�q�<ލ�<���<���<���<O��<���<��<��<���<���<���<?��<ܛ�<�w�<L�<��<���<Δ�<�E�<���<=��<"�<��<�3�<��<�$�<j��<��<~U�<(��<?��<�H�<��<˷<C�<�5�<b�<)��<��<+Ȭ<��<s��<��<��<4 �<�)�<�1�<48�<�=�<�B�<hF�<�I�<L�<�M�<N�<UM�<@K�<�G�<�B�<y<�<�4�<�+�<fD~</z<�v<Pr<��m<9�i<}�e<�a<��]<r�Y<�tU<�dQ<�UM<�GI<x:E<V-A<� =<�9<&	5<��0<��,<��(<4�$<�� <��<��<V<<�4<�W	<�<�<u��;`\�;���;���;3;�;���;���;G��;���;ӣ�;³;>��;MG�;y��;C;�;�;ު�;?��;I��;��u;�8j;`_;(CT;��I;�U?;=5;<c+;�!;�`;p7;�G;�"�:s'�:��:��:޹:��:I˛:i[�:|�~:�c:L1H:��-:F:j#�9���9�Z�9��@9���8Eϕ�O����@�y,��� ��m�i@�!$���:��9Q�ӈg�b�}��ۉ��Ԕ�8���$���.����{��Wk˺_ֺ.[Ẍ[�b���4����!9�^���+���u�!�1\'���,�9�1�-D7��<���A�:G��IL�K�Q�f�V�8.\�x�a��f��Kl���q�F"w��|�H ����n���$��*ً�򌎻�?����%���Z���  �  !�=�G=R�=O�=�?=��=r�=�3=�� =� =�% =���<]��<�1�<��<���<��<�n�<���<s�<a�<3��<� �<�N�<+��<��<�2�<�{�<���<�
�<UP�<#��<��<!�<y^�<��<���<[ �<�^�<Û�<��<f�<OG�<�{�<���<.��<��<2-�<�P�<�p�<׌�<q��<>��<l��<���<,��<���<���<���<���<���<<��<
��<Sw�<�K�<��<���<��<(F�<(��<��<#�<>��<�4�<���<&�<��<���<W�<���<���<�I�<	��<�˷<��<�5�<5b�< ��<ߪ�<�Ǭ<(�<���<��<�<��<_(�<0�<�6�<0<�<A�<E�<qH�<K�<�L�<MM�<�L�<�J�<�G�<�B�<�<�<@5�<�,�<�E~<1z<;v<�r<]�m< �i<��e<�a<p�]<�Y<�vU<�fQ<�WM<)II<S;E<�-A<� =<b9<�5<z�0<�,<��(<�$<�� <O�<��<� <�<�1<�T	<F<g�<���;QX�;���;��;�9�;��;���;ש�;��;���;ų;?��;�K�;~��;�@�;��;���;ř�;���;�u;Aj;*#_;!IT;�I;�W?;5>5;ib+;g�!;H];2;
A;��:��:҉�:=p�:�Ĺ:��:o��:�A�:�`~:(�b:�H:[�-:��:���9d��9�N�9��@9���8\���c���?�*������� ���H�#���:��
Q�L[g���}�ɉ�PÔ�곟�������x���i˺�`ֺ�^��c��l��<����{B���[6���*"�-i'���,��2�`N7�}�<���A�WG��NL�6�Q���V�9.\�օa��f��Fl�_�q��w��|�I���R����h�����wӋ�\����:��&/����V���  �  ��=�C=��=x�=�:=��=�=G.=?� =z =� =Ƌ�<���<w$�<�q�<���<��<[�<���<���<�E�<���<I��<0,�<�v�<���<	�<AP�<3��<��<��<�a�<D��<��<�#�<�b�<���<f��<��<jR�<L��<��<���<�$�<�R�<�}�<C��<���<8��<e�<� �<m6�<;H�<_V�<{`�<�f�<Hh�<Re�<�]�<CP�<n=�<$�<[�<3��<���<x�<(9�<��<P��<�I�<��<��<F�<���<�<É�<I��<�a�<�¿<��<�q�<ƿ�<s�<0I�<��<l��<>�<��<>�<�`�<@~�<��<`��<���<]Ң<��<|�<���<U�<�
�<��<�<��<B#�<�&�<�(�<�)�<p)�<�'�<�$�<� �<��<
+~<�z<:v< r<�m<��i<��e<��a< �]<�Y<w�U<͘Q<�M<�I<-�E<�zA<gu=<�p9<_m5<@k1<)k-<"m)<$r%<�z!<��<��<�<��<��<y
<6O<��<��;"�;��;o�;�,�;c��;���;m��;1��;h�;��;�Z�;͹�;�3�;Qɛ;�|�;�N�;z?�;*Q�;{;��o;ڎd;�Y;�O;'�D;�:;S�0;';,�;�f;�h;��;�"�:an�:�(�:cK�:Iֳ:�ä:f�:Ƴ�:�Ts:��W:�<:7{":�n:��9@٪9hnq9�=9�/8V��"�/�u��~���ٹ�1�ae��c2��8I���_�hv�g��M���'�������ʲ�jؽ�i�Ⱥ��Ӻ+ߺa"�u9���' �����8�t���8�	���!�r�&���+��C1���6�|�;��;A�ƊF���K�O0Q�ʈV��[��Ea���f��l���q���v��i|�ɨ���b������ԋ�H���tD��:���Ǵ���n���  �  ��=�C=��=}�=�:=��=�=P.=Z� =Ez =&  =(��<Z��<�$�<�q�<a��<Y�<�[�<��<-��<(F�<���<l��<A,�<w�<���<��<)P�<��<���<��<.a�<��<���<�#�<b�<S��<��<B�<R�<��<���<���<~$�<�R�<�}�<U��<���<]��<��<� �<�6�<�H�<�V�<�`�<�f�<�h�<�e�<�]�<�P�<�=�<j$�<{�<R��<���<x�<B9�<���<2��<�I�<���<��<��<!��<��<q��<���<-a�<�¿<G�<yq�<l��<?�<I�<���<N��<6�<��<�>�<�`�<S~�<D��<���<¤<�Ң<O�<��<���<��<Y�<��<w�<	�<}#�<�&�<
)�<�)�<�)�<�'�<�$�<� �<p�<�*~<z<�v<X�q<D�m</�i<��e<��a<A�]<Y�Y<ġU<-�Q<��M<͇I<�E<�zA<xu=<�p9<�m5<�k1<Mk-<�m)<�r%<�{!<��<��<ױ<L�<Z�<E
<P<;�<?��;�"�;l��;�o�;2-�;��;���;��;���;��;B�;�Y�;���;2�;!ț;:{�;M�;L>�;�O�;M{;g�o;�d;)�Y;�O;p�D;��:;0�0;�';y�;.h;�i;ݢ;�'�:�t�:�.�:BR�:k۳:�Ȥ:3�:
��:�as:K�W:��<:�":+s:��9�ܪ90}q9K;9�/8�BV�83��v�����Ծٹ�>��n��o2�jDI��_��sv�yl������������I̲�ڽ���Ⱥ��ӺRߺF �8���& ���Y6�8���5�����!���&�o�+��@1���6���;��9A��F�y�K�c/Q�އV���[��Fa�[�f��l��q�	�v�wl|�����E���d�����Ջ������E������ ���Uo���  �  @�=�C=��=t�=�:=��=V�=�.=�� =�z =�  =��<[��<&�<s�<���<O�<u\�<���<���<�F�<.��<���<w,�<$w�<���<��<�O�<|��</��<��<a`�<��<���<~"�<ba�<G��<���<p�<NQ�<P��<Z��<��<:$�<fR�<�}�<s��<��<���<"�<�!�<�7�<�I�<�W�<�a�<
h�<�i�<�f�<�^�<�Q�<{>�<2%�<�<���<��<$x�<?9�<���<��<RI�<C��<�~�<�<D��<��<T��<���<`�<~��<8�<�p�<���<y�<_H�<���<��<�<��<�>�<�`�<�~�<혨<q��<�¤<�Ӣ<<�< �<��<��<`�<��<]�<��<H$�<{'�<�)�<F*�<�)�<�'�<�$�<e �<��<t)~<�z<�v<��q<-�m<
�i<}�e<��a<!�]<��Y<%�U<��Q<B�M<��I<H�E<KzA<Lu=<!q9<n5<|l1<�l-<o)<ht%<R}!<t�<��<?�<��<��<I 
<R<��<���;&�;���;�q�;H.�;���;t��;���;���;��;��;�V�;���;{.�;+ě;w�;�H�;K:�;�K�;�z;��o;k�d;M�Y;~O;��D;��:;k�0;�';I�;fl;	o;��;�4�:%��:">�:�c�:Y�:�ۤ:�&�:ɇ:8�s:yX:�=:�":�:���9��9F�q9�%9�!/8�$W�M��#pv��Ū�
�ٹ$_�P����2��gI�G`���v�y��꜑�T����Ƨ�ZҲ�lݽ���Ⱥ��Ӻ[ߺ��/��! �����/����C.����3!�Y{&�9�+�791�|�6���;��3A� �F���K�B-Q��V���[�fHa���f��l�\�q�%�v��r|���h���Xh���!��ڋ�둎�qI��� �����r���  �  �=cC=��=i�=�:=��=��=/=@� =O{ =V! =͎�<��<�'�<�t�<:��<�<#^�<7��<3��<�G�<��<c��<�,�<?w�<c��<b�<O�<���<"��<z�<�^�<`��<��<� �<�_�<���<c��<��<�O�<*��<x��<Z��<�#�<(R�<�}�<ť�<p��<���<	�<�"�<�8�<K�<gY�<�c�<�i�<sk�<h�<�`�<)S�<�?�<J&�<�<���<l��<ox�<49�<w��<K��<�H�<S��<�}�<��<���<��<{��<���<9^�<���<��<o�<,��<J�<{G�<Ã�<}��<��<��<�>�<ia�<��<ܙ�<���<FĤ<Nբ<��<��<���<��<�<��<��<)!�<Z%�<h(�<2*�<�*�<�)�<�'�<^$�<��<9�<�'~<1z<
v<r�q<��m<��i<2�e<R�a<Ĳ]<S�Y<$�U<�Q<4�M<0�I<�~E<�yA<u=<wq9<�n5<�m1<Qn-<0q)< w%<b�!<��<)�<ȷ<Q�<F�<�#
<�U<�<��;g*�;���;"t�;<0�;n��;?��;N��;V��;9�;��;R�;���;�(�;���;�p�;�B�;�3�;�E�;>�z;ږo;�~d;��Y;jO;��D;�:;ʸ0;�';�;fr;�v;��;�J�:���:<Z�:_�:+
�:g��:XB�:)�:׳s:�/X:v4=:�":��:z��9q��9��q9�9N.8�X����4 w����bSڹԑ����Z�2�-�I�GF`���v����������Ɯ�`ӧ�nݲ��佺��Ⱥy�Ӻߺ���!�� ���=$�]��2 ���G!��m&�d�+�n+1�`�6�!�;�+A��}F���K��)Q�/�V�b�[��Ja�g�f�z"l��q��w�`~|�A���ﴃ�4o��(�����������O�����񽖻v���  �  _�=�B=`�=]�=�:=2�=�=�/=�� =/| =E" =А�<I��<*�<w�<���<;�<`�<��<���<=I�<(��<0��<V-�<`w�<D��<��<DN�<���<���<��<
]�<m��<���<��<t]�<Z��<a��<��<1N�<���<0��<f��<#�<�Q�<�}�<��<��<���<O
�<Z$�<�:�<�L�<z[�<�e�<
l�<�m�<�j�<�b�<U�<�A�<�'�<:�<~��<��<�x�< 9�<,��<���<�G�<���<�{�<�	�<���<��<)��<���<�[�<]��<o�<�l�<_��<��<4F�<���<ֹ�<}�<��<Q?�<b�<���<��<(��<Ƥ<-ע<�<��<��<��<Q�<��<��<�"�<�&�<�)�<$+�<U+�<4*�<�'�<$�<�<:�<�$~<z<�v<��q<��m<�i<��e<��a<��]<^�Y<t�U<ϐQ<X�M<�I<F}E<�xA<�t=<�q9<�o5<eo1<�p-<t)<�z%<2�!<�<��<��<%�<�<w(
<�Y<�<��;J0�;���;�w�;�2�;s��;D��;���;m��;Nݼ;~�;L�;���;7!�;���;h�;�9�;J+�;>�;��z;�o;:sd;&�Y;fO;�D;��:;�0;�';��;�z;/�;�;ch�:P��:#|�:ţ�:�/�:��:�f�:U�:��s:8jX:�f=:O�":�:���9��9��q9��9z�,8[Z�l��q�w�����ڹg�����3���I�*�`�xw����H̑�ޜ��姺v벺���Ⱥ��Ӻ�޺��>��l � ��������σ��� �%[&���+�1�^t6���;�cA�!tF�(�K�+%Q�-�V���[��Ma���f��*l�Ǟq�;w�z�|����$���%x��M1���鋻Ӡ��nW�����OĖ��{���  �  ��=�B=�=G�=;=}�=��=L0=�� = } =a# =H��<���<�,�<�y�<'��<��<�b�<0��<���<�J�<^��<!��<�-�<�w�<��<P�<cM�<C��<��<��<�Z�<��<P��<��<�Z�<֘�<���<��<&L�<��<���<E��<M"�<xQ�<�}�<j��<���<���<��<&�<�<�<OO�<�]�<ph�<�n�<^p�<Im�<
e�<WW�<�C�<�)�<��<���<���< y�<
9�<���<ȟ�<SF�<[��<z�<��<'��< �<}��<���<Y�<���<��<�j�<J��<��<�D�<���<��<	�<��<�?�<�b�<���<���<賦<Ȥ<�٢<��<���<� �<�
�<��<�< �<�$�<�(�<+�<4,�< ,�<{*�<�'�<�#�<T�<�<�!~<rz<Lv<��q<��m<��i<(�e<��a<E�]<e�Y<�U<�Q<'�M<T�I<�{E<�wA<mt=<6r9<q5<dq1<Fs-<uw)<]~%<��!<�<�<�<��<�<�-
<�^<��<���;C7�;,��;.|�;25�;���;���;��;y��;^ؼ;��;E�;���;��;׫�;C^�;�/�;�!�;4�;��z;_zo;fd;��Y; O;�D;��:;��0;';�;��;�;��;���:D��:3��:R��:�Z�:�G�:���:,/�:Y=t:��X:��=:�#:��:�&�9�,�9S�q9ؼ9��+8X|\�K�ۚx��	��S`۹�#�^�e3�*8J���`�<Uw��҆��ꑺ���i���{���������Ⱥ��Ӻ��޺�麃���� �`����}�����n�a� ��E&�?�+�a1�?b6���;��A��iF���K� Q�.�V���[�PQa���f�j4l��q��#w�9�|����ǃ�;����;���(���,a��K���˖������  �  �=B=��=9�=8;=��=�=�0=�� =&~ =�$ =ԕ�<���<�/�<�|�<���<k�<e�<u��<���<�L�<���<��<[.�<�w�<Ŀ�<��<HL�<ɐ�<Z��<��<�X�<j��<���<(�<�W�<��<#��<G�<�I�<���<&��<���<k!�<�P�<�}�<Ȧ�<���<���<8�<�'�<�>�<�Q�<�`�<2k�<|q�<+s�<p�<�g�<�Y�<�E�<_+�<
�<���<m��<Ly�<9�< ��<ў�<�D�<���<x�<0�<���<4�<�~�<���<V�<���<�<h�<䶺<���<�B�<^��<(��<��<��<�?�<�c�<Ȃ�<)��<͵�<;ʤ<ܢ<"�<S��<��<U�<��<��<s"�<�&�<o*�<n,�<C-�<�,�<�*�<�'�<#�<c�<��<�~<ez<��u<��q<�m<M�i<C�e<�a<ģ]<b�Y<U�U<ǈQ<��M<j}I<�yE<@vA<"t=<�r9<@r5<\s1<�u-<{)<��%<{�!<R�<w�<��<v�<c	<N3
<d<X�<���;�>�;���;`��;�7�; �;y��;���;���;Ӽ;O��;�<�;���;=�;}��;|S�;�$�;�;�)�;�z;�ho;�Wd;e�Y;�N;��D;��:;��0;�';��;B�;z�;�;��:�	�:���:Z��:���:zu�:���:zY�:M�t:��X:��=:>#:^	:MX�9�F�9Ӗq9��9��)8��^���W�y�������۹�w�P��D�3�%�J�	4a���w�3���������L���������Ⱥ��Ӻ!�޺h��A�������t���
�em����8X��� �/&�g�+���0�<O6�*�;�A�`^F���K��Q��~V�C�[�Va�F�f�e?l��q��3w�ү|�;��=҃�b����G��<��������j������Ӗ�R����  �  _�=�A=��=�=J;= �=��=�1=�� =3 =�% =L��<@��<S2�<u�<���<�<xg�<ƴ�<��<+N�<���<���<�.�<�w�<p��<��<>K�<]��<���<��<V�<Ӗ�<���<S�<U�<?��<|��<��<�G�<��<}��<���<� �<�P�<r}�<��<O��<���<��<�)�<�@�<T�<c�<�m�<Nt�<v�<�r�</j�<\�<�G�<)-�<��<���<(��<�y�<�8�<���<��<�C�<���<�u�<��< ��<f�<�{�<���<S�<ȴ�<:�<we�<���<���<SA�<�<I��<�<��<_@�<ad�<���<���<���<w̤<Tޢ<��<��<j�<#�<P�<*�<�$�<%)�<.,�<�-�<a.�<l-�<+�<m'�<|"�<~�<f�<$~<a
z<�u<��q<��m<��i<��e<)�a<@�]<1�Y<��U<��Q<M<�zI<wwE<�tA<�s=<�r9<�s5<ku1<�x-<z~)<͆%<<�!<`�<�<��<v�<+<�8
<-i<B�<��;�E�;���;���;�:�;� �;���;���;��;�ͼ;��; 5�;���;l�;
��;�H�;��;N�;��;Ȫz;�Wo;�Hd;�zY;��N;��D;��:;��0;�';F�;��;�;��;���:0�:L��:�&�:���:ʣ�: �:���:#�t:T9Y:�>:�n#:#-	:4��9i_�9�q9�S9/I(8Ca�H��7�z��'����ܹ���8��4���J�Ҍa�.�w���E0���2���+��������^�Ⱥ��Ӻ�޺��,������e���
�fZ����	B��� ��&��}+���0��<6��;�N�@��RF��K�DQ��|V�/�[�|Za���f�~Il���q��Cw��|�Y���܃������R���
������$u���(��ܖ�u����  �  ��=A=9�=��=c;=d�=��=U2=Q� =� =�& =���<���<�4�<��<I��<��<�i�<ܶ�<�<�O�<,��<���<b/�<�w�<*��<B�<2J�<��<���<��<�S�<[��<J��<��<sR�<���< ��<Y
�<�E�<0�<���<���<��<P�<_}�<n��<���<���<"�<i+�<�B�<GV�<�e�<kp�<�v�<�x�<<u�<�l�<D^�<�I�<�.�<��<���<���<�y�<�8�<��<��<iB�<S��<	t�<� �<s��<��<�x�<���<1P�<��<��<�b�<~��<���<�?�<�}�<l��<��<��<�@�<�d�<��<��<V��<uΤ<��<L�<���<	�<��<��<�!�<�&�<+�<�-�<N/�<C/�<.�<V+�<J'�< "�<��<.�<�~<�z<��u<��q<��m<8�i<.�e<Ĥa<�]<'�Y<�U<��Q<�{M<xI<buE<�sA<s=<Hs9<�t5<�v1<o{-<��)<��%<��!<d�<T�<��<��<j<O>
<+n<��<���;YL�;-��;H��;A=�;��;E��;���;���;"ɼ;/�;.�;R��;��;U��;w>�;��;K�;V�;4�z;/Ho;�:d;ioY;2�N;1�D;��:;ù0;�"';��;*�;ɱ;��;\��:�T�:U!�:�O�:=�:�ͥ:��:���:Q!u:'yY:�O>:��#:}N	:Y��9%x�9[�q9%!9�&8c�����f{������-ݹ�Uc��p4�ICK���a�EIx�1D��jO���N��UB��/�����ɺ=�Ӻ��޺��麴���)����V��
��G�����-��� �,&��h+���0�++6��;���@��GF�8�K��Q�{V��[��^a�P�f�YSl���q��Rw�K�|�/)��烻K���b]��0���ʎ����1���㖻%����  �  '�=�@=��=�=p;=��=d�=�2=� =� =�' =���<���<7�<g��<���<��<�k�<���<�<Q�<)��<s��<�/�<�w�<��<��<@I�<Ȍ�<L��<��<�Q�<L��<��<V�< P�<Y��<���<p�<�C�<�}�<���<���<��<�O�<K}�<���<z��<���<K�<�,�<�D�<)X�<�g�<�r�<y�<�z�<`w�<�n�<"`�<pK�<80�<�<��<?��<�y�<�8�<���<$��<?A�<���<Ur�<���<k��< �<fv�<b��<�M�<���<\�<�`�<���<R��<`>�<�|�<���<6�<��<�@�<�e�<셪<?��<κ�<Ф<{�<F�<���<P�<��< �<�#�<�(�<�,�<>/�<i0�< 0�<�.�<{+�<+'�<�!�<��<�<,~<Iz<�u<��q<5�m<��i<r�e<�a<��]<�Y<C�U</}Q<�xM<�uI<�sE<�rA<�r=<ss9<au5<�x1<�}-<s�)<͍%<L�!<\�<��<�<��<<�B
<7r<b�<{��;#R�;���;Ƌ�;?�;��;���;ż�;3��;�ļ;��;I'�;F�;H�;ۄ�;�5�;��;���;"�;��z;L:o;�.d;�eY;�N;�D;ۈ:;��0;�$';��;��;}�;�;�
�:[s�:.A�:�r�:�:��:�5�:�̈:�^u:9�Y:�>:��#:�k	:���9у�9�q9/�9;9%8=�e��<�l1|������ݹ6_����4�z�K��&b��x�7b��Wl���f��\V���>���#��Oɺ��Ӻ��޺s��?���m����J�\�
�U8����>�0� ��%�!X+�[�0�o6��|;�5�@�6?F���K��Q�*zV���[��ba���f��\l���q�A`w��|�
1���q����f��^���ӎ�����9��yꖻ�����  �  ��=f@=��=В=|;=��=��=93=�� =�� =m( =?��<���<�8�<��<;��<Y �<Um�<��<<�<�Q�<ߜ�<	��<�/�<�w�<���<:�<�H�<ߋ�<<��<��<oP�<���<V��<��<bN�<���<��<��<HB�<a|�<���<���<y�<EO�<:}�<§�<���<j��<�<�-�<�E�<�Y�<i�<Et�<�z�<u|�<y�<1p�<�a�<�L�<K1�<��<"��<���< z�<m8�<(��<���<a@�<���<q�<8��<���<���<�t�<���<�K�<խ�<�	�<K_�<��<!��<Z=�<�{�<%��<��<w�<	A�<f�<���<��<黦<|Ѥ<�<��<n�<��<��<��<,%�<U*�<�-�<K0�<,1�<�0�<�.�<�+�<'�<$!�<:�<4�<(~<� z<�u<y�q<��m< �i<�e<��a<�]<��Y<0�U<�zQ<�vM<�sI<drE<�qA<;r=<�s9<v5<�y1<-<|�)<G�%<L�!<��<
�< �<�<�<�E
<�u<p�<���;CV�;���;���;�@�;�;
��;n��;��;m��;��;d"�;�y�;��;F~�;/�;B �;�;d�;}z;B/o;�%d;^Y;�N;y�D;$�:;��0;o&';��;�;8�;�; �:���:�Z�:���:��:7�:�Q�:�:��u:��Y:�>:��#:��	:���9I��9{q9*�9Q$8)g�#����|�;x��޹>�����s�4���K��]b�K�x�{��򁒺Ox��e���I���*��-ɺn�Ӻ��޺���������hA��
��+����s�*{ ���%��J+�ޮ0��6��r;���@�K9F�)�K��	Q�yV���[��ea��f�Scl���q�5jw��|��7������L����m��;%���ڎ�ȍ��?���ڟ���  �  h�=)@=��==�;=��=ߋ=3=�� =� =�( =(��<���<�9�<'��<I��<a!�<0n�<Ժ�<��<�R�<b��<Q��</0�<�w�<���<��<H�<>��<q��<��<�O�<���<L��<s�<3M�<���<)��<��<|A�<�{�<���<,��<�<O�<)}�<��<(��<���<��<�.�<�F�<lZ�<j�<Mu�<�{�<�}�<z�<1q�<bb�<�M�<�1�<z�<���<��<?z�<X8�<���<1��<�?�<'��<8p�<`��<���<���<is�<K��<�J�<���<��<K^�<9��<@��<�<�<m{�<ƴ�<��<m�<-A�<Jf�<���<���<���<=Ҥ<��<���<w�<�<��<��<&�<"+�<�.�<1�<�1�<.1�</�<�+�<�&�<� �<��<��<�~<5�y<Z�u<��q<��m<ζi<��e<?�a<�]<��Y<o~U<�xQ<uM<�rI<cqE<=qA<�q=<�s9<gv5<�z1<�-<߇)<ܑ%<�!<k�<0�<6�<c�<�< H
<Rw<�<���;&Y�;��;ڏ�;�A�;r�;���;���;B��;$��;��;k�;v�;6�;Tz�;�*�;���;��;��;�uz;:)o;�d;�XY;��N;��D;�:;C�0;�'';��;Я;D�;f;�,�:���:�j�:h��:�1�:3�:�b�:j��:�u:��Y:�>:��#:��	:.�9˜�9vq94�9�#8k8h���,}�J���'L޹����,5��K�nb��x�񉇺����G���o��R���/���ɺ5�Ӻ��޺D��]�������];�ư
�1%����
�Br ���%�DB+�S�0�;
6��l;�W�@��4F�_�K�iQ�3xV��[��ga���f�hl���q��pw���|��;������ⷆ�^r���)���ގ������B����ߢ���  �  `�=@=��=��=�;=��=�=�3=�� =� =�( =���<���<9:�<���<���<�!�<�n�<,��<E�<�R�<~��<i��<E0�<�w�<o��<��<�G�<'��<3��<��<!O�<@��<���<�<�L�<��<���<n�<*A�<D{�<ͳ�<��<��<O�<
}�<��<A��<���<��<�.�<�F�<�Z�<tj�<�u�<6|�<�}�<fz�<�q�<�b�<�M�<22�<��<���<���<@z�<78�<���<��<�?�<���<�o�<��<@��<;��<�r�<���<OJ�<@��<�<�]�<歺<���<�<�<B{�<���<��<Q�<7A�<_f�<��<ң�<޼�<�Ҥ<(�<<��<��<n�<�< �<|&�<z+�</�<(1�<�1�<H1�<;/�<�+�<�&�<� �<��<��<U~<��y<��u<��q<��m<�i<��e<z�a<?�]<�Y<�}U<HxQ<�tM<frI<qE<qA<�q=<�s9<�v5<�z1<[�-<)�)<}�%<��!<%�<��<��<8�<y<�H
<x<ح<���;�Y�;���;Q��;B�;;�;���;!��;ʱ�;ܾ�;��;7�;�t�;��;�x�;W)�;���;'�;R�;�rz;�&o;#d;�WY;G�N;��D;��:;^�0;(';z�;��;P�;�;-2�:��:q�:��:�7�:B%�:8g�:���:c�u:��Y:	�>:��#:W�	:w�99hgq9�9�H#89vh����S}�齮�f޹������!5�_�K�A�b���x�[���t��������p��XT��J2��5ɺ��Ӻ��޺���k�������d9��
�c"������o ��%��?+�g�0��6�-j;�%�@��3F���K��Q�9xV���[�#ha���f��hl�D�q�
sw�f�|�=��-���q����s��i+��4�������C����������  �  h�=)@=��==�;=��=ߋ=3=�� =� =�( =(��<���<�9�<'��<I��<a!�<0n�<Ժ�<��<�R�<b��<Q��</0�<�w�<���<��<H�<>��<q��<��<�O�<���<L��<s�<3M�<���<)��<��<|A�<�{�<���<,��<�<O�<)}�<��<(��<���<��<�.�<�F�<lZ�<j�<Mu�<�{�<�}�<z�<1q�<bb�<�M�<�1�<z�<���<��<?z�<X8�<���<1��<�?�<'��<8p�<`��<���<���<is�<K��<�J�<���<��<K^�<9��<@��<�<�<m{�<ƴ�<��<m�<-A�<Jf�<���<���<���<=Ҥ<��<���<w�<�<��<��<&�<"+�<�.�<1�<�1�<.1�</�<�+�<�&�<� �<��<��<�~<5�y<Z�u<��q<��m<ζi<��e<?�a<�]<��Y<o~U<�xQ<uM<�rI<cqE<=qA<�q=<�s9<gv5<�z1<�-<��)<ܑ%<�!<k�<0�<6�<c�<�< H
<Rw<�<���;%Y�;��;ڏ�;�A�;q�;���;���;B��;#��;��;j�;v�;6�;Tz�;�*�;���;��;��;�uz;:)o;�d;�XY;��N;��D;�:;C�0;�'';��;Я;D�;f;�,�:���:�j�:h��:�1�:3�:�b�:j��:�u:��Y:�>:��#:��	:.�9˜�9vq94�9�#8k8h���,}�J���'L޹����,5��K�nb��x�񉇺����G���o��R���/���ɺ5�Ӻ��޺D��]�������];�ư
�1%����
�Br ���%�DB+�S�0�;
6��l;�W�@��4F�_�K�iQ�3xV��[��ga���f�hl���q��pw���|��;������ⷆ�^r���)���ގ������B����ߢ���  �  ��=f@=��=В=|;=��=��=93=�� =�� =m( =?��<���<�8�<��<;��<Y �<Um�<��<<�<�Q�<ߜ�<	��<�/�<�w�<���<:�<�H�<ߋ�<<��<��<oP�<���<V��<��<bN�<���<��<��<HB�<a|�<���<���<y�<EO�<:}�<§�<���<j��<�<�-�<�E�<�Y�<i�<Et�<�z�<u|�<y�<1p�<�a�<�L�<K1�<��<"��<���< z�<m8�<(��<���<a@�<���<q�<8��<���<���<�t�<���<�K�<խ�<�	�<K_�<��<!��<Z=�<�{�<%��<��<x�<	A�<f�<���<��<黦<|Ѥ<�<��<n�<��<��<��<,%�<T*�<�-�<K0�<,1�<�0�<�.�<�+�<'�<$!�<:�<4�<(~<� z<�u<y�q<��m< �i<�e<��a<�]<��Y<0�U<�zQ<�vM<�sI<drE<�qA<;r=<�s9<v5<�y1<-<|�)<G�%<L�!<��<
�< �<�<�<�E
<�u<p�<���;CV�;���;��;�@�;�;
��;n��;��;l��;��;d"�;�y�;��;F~�;/�;A �;�;c�;}z;B/o;�%d;^Y;�N;y�D;$�:;��0;o&';��;�;8�;�; �:���:�Z�:���:��:7�:�Q�:�:��u:��Y:�>:��#:��	:���9I��9{q9*�9Q$8)g�#����|�;x��޹>�����s�4���K��]b�K�x�{��򁒺Ox��e���I���*��-ɺn�Ӻ��޺���������hA��
��+����s�*{ ���%��J+�ޮ0��6��r;���@�K9F�)�K��	Q�yV���[��ea��f�Scl���q�5jw��|��7������L����m��;%���ڎ�ȍ��?���ڟ���  �  '�=�@=��=�=p;=��=d�=�2=� =� =�' =���<���<7�<g��<���<��<�k�<���<�<Q�<)��<s��<�/�<�w�<��<��<@I�<Ȍ�<L��<��<�Q�<L��<��<V�< P�<Y��<���<p�<�C�<�}�<���<���<��<�O�<K}�<���<z��<���<K�<�,�<�D�<)X�<�g�<�r�<y�<�z�<`w�<�n�<"`�<pK�<80�<�<��<?��<�y�<�8�<���<$��<?A�<���<Ur�<���<k��< �<fv�<b��<�M�<���<\�<�`�<���<R��<`>�<�|�<���<6�<��<�@�<�e�<셪<@��<κ�<Ф<{�<F�<���<P�<��< �<�#�<�(�<�,�<>/�<i0�< 0�<�.�<{+�<+'�<�!�<��<�<,~<Iz<�u<��q<5�m<��i<r�e<�a<��]<�Y<C�U</}Q<�xM<�uI<�sE<�rA<�r=<ts9<bu5<�x1<�}-<t�)<͍%<L�!<\�<��<�<��<<�B
<6r<b�<z��;"R�;���;Ƌ�;?�;�;���;ļ�;3��;�ļ;��;I'�;F�;H�;ڄ�;�5�;��;���;"�;��z;L:o;�.d;�eY;�N;�D;ۈ:;��0;�$';��;��;}�;�;�
�:[s�:.A�:�r�:�:��:�5�:�̈:�^u:9�Y:�>:��#:�k	:���9у�9�q9/�9;9%8=�e��<�l1|������ݹ6_����4�z�K��&b��x�7b��Wl���f��\V���>���#��Oɺ��Ӻ��޺s��?���m����J�\�
�U8����>�0� ��%�!X+�[�0�o6��|;�5�@�6?F���K��Q�*zV���[��ba���f��\l���q�A`w��|�
1���q����f��^���ӎ�����9��yꖻ�����  �  ��=A=9�=��=c;=d�=��=U2=Q� =� =�& =���<���<�4�<��<I��<��<�i�<ܶ�<�<�O�<,��<���<b/�<�w�<*��<B�<2J�<��<���<��<�S�<[��<J��<��<sR�<���< ��<Y
�<�E�<0�<���<���<��<P�<_}�<n��<���<���<"�<i+�<�B�<GV�<�e�<kp�<�v�<�x�<<u�<�l�<D^�<�I�<�.�<��<���<���<�y�<�8�<��<��<iB�<S��<	t�<� �<s��<��<�x�<���<1P�<��<��<�b�<~��<���<�?�<�}�<l��<��<��<�@�<�d�<��<��<W��<uΤ<��<L�<���<	�<��<��<�!�<�&�<+�<�-�<N/�<C/�<.�<V+�<J'�< "�<��<.�<�~<�z<��u<��q<��m<8�i<.�e<Ĥa<�]<'�Y<�U<��Q<�{M<xI<buE<�sA<	s=<Is9<�t5< w1<o{-<��)<��%<��!<d�<T�<��<��<j<O>
<+n<��<���;YL�;,��;H��;@=�;��;D��;���;��;!ɼ;.�;.�;R��;��;U��;v>�;��;J�;V�;3�z;.Ho;�:d;hoY;2�N;0�D;��:;¹0;�"';��;*�;ɱ;��;\��:�T�:U!�:�O�:=�:�ͥ:��:���:Q!u:'yY:�O>:��#:}N	:Y��9%x�9[�q9%!9�&8c�����f{������-ݹ�Uc��p4�ICK���a�EIx�1D��jO���N��UB��/�����ɺ=�Ӻ��޺��麴���)����V��
��G�����-��� �,&��h+���0�++6��;���@��GF�8�K��Q�{V��[��^a�P�f�YSl���q��Rw�K�|�/)��烻K���b]��0���ʎ����1���㖻%����  �  _�=�A=��=�=J;= �=��=�1=�� =3 =�% =L��<@��<S2�<u�<���<�<xg�<ƴ�<��<+N�<���<���<�.�<�w�<p��<��<>K�<]��<���<��<V�<Ӗ�<���<S�<U�<?��<|��<��<�G�<��<}��<���<� �<�P�<r}�<��<O��<���<��<�)�<�@�<T�<c�<�m�<Nt�<v�<�r�</j�<\�<�G�<)-�<��<���<(��<�y�<�8�<���<��<�C�<���<�u�<��< ��<f�<�{�<���<S�<ȴ�<:�<we�<���<���<SA�<�<I��<�<��<_@�<ad�<���<���<���<w̤<Tޢ<��<��<j�<#�<P�<*�<�$�<%)�<.,�<�-�<a.�<k-�<+�<m'�<|"�<}�<f�<#~<a
z<�u<��q<��m<��i<��e<)�a<@�]<1�Y<��U<��Q<M<�zI<wwE<�tA<�s=<�r9<�s5<ku1<�x-<{~)<͆%<<�!<`�<�<��<v�<+<�8
<,i<A�<��;�E�;���;���;�:�;� �;���;���;��;�ͼ;��; 5�;;l�;	��;�H�;��;M�;��;Ȫz;�Wo;�Hd;�zY;��N;��D;��:;��0;�';F�;��;�;��;���:0�:L��:�&�:���:ʣ�: �:���:#�t:T9Y:�>:�n#:#-	:4��9i_�9�q9�S9/I(8Ca�H��7�z��'����ܹ���8��4���J�Ҍa�.�w���E0���2���+��������^�Ⱥ��Ӻ�޺��,������e���
�fZ����	B��� ��&��}+���0��<6��;�N�@��RF��K�DQ��|V�/�[�|Za���f�~Il���q��Cw��|�Y���܃������R���
������$u���(��ܖ�u����  �  �=B=��=9�=8;=��=�=�0=�� =&~ =�$ =ԕ�<���<�/�<�|�<���<k�<e�<u��<���<�L�<���<��<[.�<�w�<Ŀ�<��<HL�<ɐ�<Z��<��<�X�<j��<���<(�<�W�<��<#��<G�<�I�<���<&��<���<k!�<�P�<�}�<Ȧ�<���<���<8�<�'�<�>�<�Q�<�`�<2k�<|q�<+s�<p�<�g�<�Y�<�E�<_+�<
�<���<n��<Ly�<9�< ��<ў�<�D�<���<x�<0�<���<4�<�~�<���<V�<���<�<h�<䶺<���<�B�<^��<(��<��<��<�?�<�c�<Ȃ�<)��<͵�<;ʤ<ܢ<"�<S��<��<U�<��<��<s"�<�&�<o*�<n,�<C-�<�,�<�*�<�'�<#�<c�<��<�~<ez<��u<��q<�m<M�i<C�e<�a<ģ]<b�Y<U�U<ǈQ<��M<j}I<�yE<AvA<"t=<�r9<Ar5<\s1<�u-<{)<��%<{�!<R�<w�<��<v�<c	<N3
<d<X�<���;�>�;���;_��;�7�; �;x��;���;���;Ӽ;O��;�<�;���;=�;|��;|S�;�$�;�;�)�;߽z;�ho;�Wd;e�Y;~�N;��D;��:;��0;�';��;B�;z�;�;��:�	�:���:Z��:���:zu�:���:zY�:M�t:��X:��=:>#:^	:MX�9�F�9Ӗq9��9��)8��^���W�y�������۹�w�P��D�3�%�J�	4a���w�3���������L���������Ⱥ��Ӻ!�޺h��A�������t���
�em����8X��� �/&�g�+���0�<O6�*�;�A�`^F���K��Q��~V�C�[�Va�F�f�e?l��q��3w�ү|�;��=҃�b����G��<��������j������Ӗ�R����  �  ��=�B=�=G�=;=}�=��=L0=�� = } =a# =H��<���<�,�<�y�<'��<��<�b�<0��<���<�J�<^��<!��<�-�<�w�<��<P�<cM�<C��<��<��<�Z�<��<P��<��<�Z�<֘�<���<��<&L�<��<���<E��<M"�<xQ�<�}�<j��<���<���<��<&�<�<�<OO�<�]�<ph�<�n�<^p�<Im�<
e�<WW�<�C�<�)�<��<���<���< y�<
9�<���<ȟ�<SF�<[��<z�<��<'��< �<}��<���<Y�<���<��<�j�<J��<��<�D�<���<��<	�<��<�?�<�b�<���<���<賦<Ȥ<�٢<��<���<� �<�
�<��<�< �<�$�<�(�<+�<4,�<�+�<{*�<�'�<�#�<T�<�<�!~<rz<Lv<��q<��m<��i<(�e<��a<E�]<e�Y<�U<�Q<'�M<T�I<�{E<�wA<mt=<6r9<q5<dq1<Fs-<uw)<]~%<��!<�<�<�<��<�<�-
<�^<��<���;C7�;+��;-|�;15�;���;���;��;y��;]ؼ;��;E�;���;��;׫�;B^�;�/�;�!�;4�;��z;^zo;fd;��Y; O;�D;��:;��0;';�;��;�;��;���:D��:3��:Q��:�Z�:�G�:���:,/�:Y=t:��X:��=:�#:��:�&�9�,�9S�q9ؼ9��+8X|\�K�ۚx��	��S`۹�#�^�e3�*8J���`�<Uw��҆��ꑺ���i���{���������Ⱥ��Ӻ��޺�麃���� �`����}�����n�a� ��E&�?�+�a1�?b6���;��A��iF���K� Q�.�V���[�PQa���f�j4l��q��#w�9�|����ǃ�;����;���(���,a��K���˖������  �  _�=�B=`�=]�=�:=2�=�=�/=�� =/| =E" =А�<I��<*�<w�<���<;�<`�<��<���<=I�<(��<0��<V-�<`w�<D��<��<DN�<���<���<��<
]�<m��<���<��<t]�<Z��<a��<��<1N�<���<0��<f��<#�<�Q�<�}�<��<��<���<O
�<Z$�<�:�<�L�<z[�<�e�<
l�<�m�<�j�<�b�<U�<�A�<�'�<:�<~��<��<�x�< 9�<,��<���<�G�<���<�{�<�	�<���<��<)��<���<�[�<]��<o�<�l�<_��<��<4F�<���<ֹ�<}�<��<Q?�<b�<���<��<)��<Ƥ<-ע<�<��<��<��<Q�<��<��<�"�<�&�<�)�<$+�<U+�<3*�<�'�<$�<�<:�<�$~<z<�v<��q<��m<�i<��e<��a<��]<_�Y<t�U<АQ<Y�M<�I<G}E<�xA<�t=<�q9<�o5<eo1<�p-<t)<�z%<3�!<�<��<��<%�<�<w(
<�Y<�<��;J0�;���;�w�;�2�;s��;D��;���;m��;Mݼ;}�;L�;���;7!�;���;h�;�9�;J+�;>�;��z;�o;9sd;%�Y;fO;�D;��:;�0;�';��;�z;/�;�;ch�:P��:#|�:ţ�:�/�:��:�f�:U�:��s:8jX:�f=:O�":�:���9��9��q9��9z�,8[Z�l��q�w�����ڹg�����3���I�*�`�xw����H̑�ޜ��姺v벺���Ⱥ��Ӻ�޺��>��l � ��������σ��� �%[&���+�1�^t6���;�cA�!tF�(�K�+%Q�-�V���[��Ma���f��*l�Ǟq�;w�z�|����$���%x��M1���鋻Ӡ��nW�����OĖ��{���  �  �=cC=��=i�=�:=��=��=/=@� =O{ =V! =͎�<��<�'�<�t�<:��<�<#^�<7��<3��<�G�<��<c��<�,�<?w�<c��<b�<O�<���<"��<z�<�^�<`��<��<� �<�_�<���<c��<��<�O�<*��<x��<Z��<�#�<(R�<�}�<ť�<p��<���<	�<�"�<�8�<K�<gY�<�c�<�i�<sk�<h�<�`�<)S�<�?�<J&�<�<���<l��<ox�<49�<w��<K��<�H�<S��<�}�<��<���<��<|��<���<9^�<���<��<o�<,��<J�<{G�<Ã�<}��<��<��<�>�<ia�<��<ܙ�<���<FĤ<Nբ<��<��<���<��<�<��<��<)!�<Z%�<h(�<1*�<�*�<�)�<�'�<^$�<��<9�<�'~<0z<

v<r�q<��m<��i<2�e<R�a<Ĳ]<S�Y<$�U<�Q<5�M<0�I<�~E<�yA<u=<wq9<�n5<�m1<Qn-<0q)< w%<b�!<�<)�<ȷ<Q�<F�<�#
<�U<�<��;g*�;���;"t�;;0�;m��;?��;M��;U��;9�;��;R�;�;�(�;���;�p�;�B�;�3�;�E�;>�z;ږo;�~d;��Y;jO;��D;�:;ʸ0;�';�;fr;�v;��;�J�:���:<Z�:_�:+
�:g��:XB�:)�:׳s:�/X:v4=:�":��:z��9q��9��q9�9N.8�X����4 w����bSڹԑ����Z�2�-�I�GF`���v����������Ɯ�`ӧ�nݲ��佺��Ⱥy�Ӻߺ���!�� ���=$�]��2 ���G!��m&�d�+�n+1�`�6�!�;�+A��}F���K��)Q�/�V�b�[��Ja�g�f�z"l��q��w�`~|�A���ﴃ�4o��(�����������O�����񽖻v���  �  @�=�C=��=t�=�:=��=V�=�.=�� =�z =�  =��<[��<&�<s�<���<O�<u\�<���<���<�F�<.��<���<w,�<$w�<���<��<�O�<|��</��<��<a`�<��<���<~"�<ba�<G��<���<p�<NQ�<P��<Z��<��<:$�<fR�<�}�<s��<��<���<"�<�!�<�7�<�I�<�W�<�a�<
h�<�i�<�f�<�^�<�Q�<{>�<2%�<�<���<��<$x�<?9�<���<��<RI�<C��<�~�<�<D��<��<T��<���<`�<~��<8�<�p�<���<y�<_H�<���<��<�<��<�>�<�`�<�~�<혨<q��<�¤<�Ӣ<<�< �<��<��<_�<��<]�<��<H$�<{'�<�)�<F*�<�)�<�'�<�$�<e �<��<t)~<�z<�v<��q<-�m<
�i<}�e<��a<!�]<��Y<%�U<��Q<B�M<��I<H�E<KzA<Lu=<!q9<n5<}l1<�l-<o)<it%<R}!<t�<��<?�<��<��<I 
<R<��<���;&�;���;�q�;G.�;���;t��;���;���;��;��;�V�;���;{.�;+ě;w�;�H�;K:�;�K�;�z;��o;j�d;L�Y;~O;��D;��:;k�0;�';I�;fl;	o;��;�4�:%��:">�:�c�:Y�:�ۤ:�&�:ɇ:8�s:yX:�=:�":�:���9��9F�q9�%9�!/8�$W�M��#pv��Ū�
�ٹ$_�P����2��gI�G`���v�y��꜑�T����Ƨ�ZҲ�lݽ���Ⱥ��Ӻ[ߺ��/��! �����/����C.����3!�Y{&�9�+�791�|�6���;��3A� �F���K�B-Q��V���[�fHa���f��l�\�q�%�v��r|���h���Xh���!��ڋ�둎�qI��� �����r���  �  ��=�C=��=}�=�:=��=�=P.=Z� =Ez =&  =(��<Z��<�$�<�q�<a��<Y�<�[�<��<-��<(F�<���<l��<A,�<w�<���<��<)P�<��<���<��<.a�<��<���<�#�<b�<S��<��<B�<R�<��<���<���<~$�<�R�<�}�<U��<���<]��<��<� �<�6�<�H�<�V�<�`�<�f�<�h�<�e�<�]�<�P�<�=�<j$�<{�<R��<���<x�<B9�<���<2��<�I�<���<��<��<!��<��<q��<���<-a�<�¿<G�<yq�<l��<?�<I�<���<N��<6�<��<�>�<�`�<S~�<D��<���<¤<�Ң<O�<��<���<��<Y�<��<w�<�<}#�<�&�<
)�<�)�<�)�<�'�<�$�<� �<p�<�*~<z<�v<X�q<D�m</�i<��e<��a<A�]<Y�Y<ġU<-�Q<��M<͇I<�E<�zA<xu=<�p9<�m5<�k1<Mk-<�m)<�r%<�{!<��<��<ױ<L�<Z�<E
<P<;�<>��;�"�;l��;�o�;2-�;��;���;��;���;��;B�;�Y�;���;2�;!ț;:{�;M�;L>�;�O�;M{;f�o;�d;)�Y;�O;p�D;��:;0�0;�';y�;.h;�i;ݢ;�'�:�t�:�.�:BR�:k۳:�Ȥ:3�:
��:�as:K�W:��<:�":+s:��9�ܪ90}q9K;9�/8�BV�83��v�����Ծٹ�>��n��o2�jDI��_��sv�yl������������I̲�ڽ���Ⱥ��ӺRߺF �8���& ���Y6�8���5�����!���&�o�+��@1���6���;��9A��F�y�K�c/Q�އV���[��Fa�[�f��l��q�	�v�wl|�����E���d�����Ջ������E������ ���Uo���  �  Q�='@=��=�=�5=z�=��=�(=�� =at = =Q�<���<a�<4b�<I��<���<�F�<6��<?��<+�<;v�<���<C
�<�R�<-��<���<�%�<�i�<o��<*��<�.�<un�<��<Z��<�&�<�a�<ƛ�<��<�
�<a?�<r�<\��<$��<���<�"�<�G�<�h�<Ά�<.��<���<���<���<���<���<j��<���<_��<���<&��<���<��<�s�<�I�<��<���<U��<�V�<]�<���<�L�<D��<�s�<���<�{�<l��<@f�<��<(5�<撽<+�<H;�<q��<�˶<��<�E�<�z�<���<S֭<��<��<�>�<�Y�<+r�<���<К�<���<I��<ɚ<h՘<x��<b�<�<���<� �<�<�	�<{�<��<�<3�<]�<d~<�
z<�v<��q<��m<=�i<��e<��a<��]<^�Y<�U<��Q<s�M<W�I<+�E<��A<��=<�9<��5<��1<]�-<X�)<Y�%<
"<�<�:<�Z<Y�<I�<��
<�<,X<�>�;���;��;gD�;B�;���;���;���;��;��;�N�;���;K�;���;�6�;D��;iϑ;�ǋ;�߅;��;��t;��i;��^;[GT;��I;��?;U�5;#,;��";pe;�Y;��;���:���:�x�:�l�:+��:�t�:���:��:���:J'g:>�K:=�0::`��9��9寐9�1<9U:�8��1�v�ڸ��N�릗� �ǹ1����	��_*�d�A��X�eo����F^�����;ڤ�&���9���fƺ��Ѻk�ܺ��續
�>/�����5
����D�����< �5�%��+�}�0���5�{K;��@��	F�jK�G�P��/V��[�va�urf�,�k��Zq�g�v��J|�l※J����\������Ջ�L���rM���	��ǖ�����  �  H�=@=��=�=�5=x�=͂=�(=�� =xt =) =��<��<��<�b�<���<���<0G�<r��<v��<*+�<Ev�<���<5
�<�R�<9��<s��<�%�<�i�<Y��<���<�.�<n�<���<��<t&�<�a�<a��<���<k
�<;?�<�q�<E��<��<���<�"�<�G�<
i�<��<<��<޷�<���<���<���<���<���<��<���<C��<u��<��<5��<t�<�I�<��<���<_��<�V�<7�<���<�L�<��<~s�<#��<Q{�<)��<�e�<���<�4�<|��<��<;�<P��<�˶<~�<�E�<�z�<
��<B֭<#��<��<�>�<Z�<_r�<���<'��<K��<���<_ɚ<�՘<���<��<H�<���<�<�<�	�<��<��<��<�<J�<S~<�
z<v<��q<��m<��i<;�e<�a<�]<��Y<��U<R�Q<\�M<.�I<��E<��A<��=<�9<��5<�1<y�-<��)<��%<�
"<� <H;<P[<�<��<W�
<�<�X<�?�;��;&��;�D�;�;5��;6��;,��;���;��;YN�;ס�;#�;6��;�5�;2�;-Α;�Ƌ;;ޅ;c�;��t;޼i;��^;�FT;�I;��?;��5;�",;5�";Bf;uZ;e�;i��:���:�~�:�q�:�Ƽ:z�:���:�:���:�,g:٨K:1�0:�:�9D��9D��9�1<9P�8�=2���ڸ�N�1����ǹb��L��i*���A�E�X��qo�����a��Ѣ��Uۤ�����;��kfƺ��ѺA�ܺ����	�.��\��54
�R���A����W: ���%�F+���0�_�5�4J;�ҩ@�1	F�0iK�(�P��/V���[��a�Lsf���k�9[q���v�M|��〻�����]��2���֋������N���
���ǖ�G����  �  	�=�?=��=�=�5=��=��=)=� =�t =} =e��<���<|�<Zc�<_��<���<�G�<��<��<�+�<�v�<��<\
�<�R�<$��<H��<I%�<i�<ë�<c��<�-�<gm�<��<I��<�%�<�`�<���<��<�	�<�>�<rq�<��<���<���<�"�<�G�<Li�<J��<���<~��<`��<���<���<���<���<���<d��<���<%��<|��<ӗ�<�t�<TJ�<��<���<T��<�V�<��<.��<TL�<x��<�r�<|��<�z�<l��<e�<���<!4�<���</�<k:�<���<0˶<"�<�E�<�z�<	��<]֭<s��<& �<"?�<�Z�<�r�<���<ܛ�<��<j��<*ʚ<p֘<��<T�<��<d��<��<��<&
�<��<��<��<��<�
�<5~<e	z<�v<��q<m�m<D�i<��e<��a<��]<Q�Y<Z�U<!�Q</�M<-�I<m�E<}�A<��=<%�9<��5<��1<d�-<��)<��%<�"<"<�<<�\<��<��<��
<<�Y<oB�;f��;��;}F�;��;���;��;���;���;��;/L�;���;��;���;3�;5�;ˑ;.ċ;�ۅ;�;��t;R�i;��^;�CT;��I;ҿ?;��5;�#,;t�";�i;]^;��;���:���:/��:&}�:�Ӽ:@��:O��:���:��:�@g:a�K:v�0:�:ª�9���9���9�#<9K�8�5�|Q۸$O��ڗ���ǹ:<��='���*�j�A���X��o�!���j��C���[㤺����>���gƺ�Ѻ��ܺY���%��A��N/
����8<�����3 �1�%��+��}0� �5�1E;� �@�tF�fK�v�P�C/V��[�a�,uf�{�k��_q���v��Q|�`总�����`������ً�����wQ��-��ʖ������  �  Ɨ=�?=z�=܎=�5=��=1�=k)=h� =Fu = =���<'��<��<�d�<���<���<I�<+��< ��<s,�<Yw�<o��<�
�<�R�<��<��<�$�<�h�<��<u��<�,�<4l�<���<���<c$�<}_�<x��<���<��<�=�<�p�<^��<x��<���<�"�<H�<�i�<Ӈ�<l��<F��<q��<���<���<��<���<-��<���<;��<?��<���<���<3u�<�J�<;�<:��<?��<lV�<��<���<�K�<���<�q�<9��<Ly�<���<�c�<���<�2�<w��<��<^9�<Մ�<�ʶ<�
�<CE�<�z�<���<�֭<���<� �<�?�<t[�<t�<ʉ�<)��<\��<���<{˚<�ט<��<t�<���<)��<:�<��<�
�<��<��<��<y�<O
�<�~<�z<��u<J�q<��m<��i<�e<��a<��]<��Y<�U<]�Q<��M<�I<�E<�A<��=<r�9<��5<��1<��-<K�)<��%<1"<�$<�?<�_<r�<T�<��
<�<R\<VF�;���;��;6H�;��;"��;���;��;��;��;vI�;J��;��;��;.�;H�;OƑ;�;�օ;��;��t;U�i;��^;@T;=�I;ľ?;��5;�&,;1�";n;bd;�;��:'�:���:s��:�:���:p��:g
�:(��:�cg:N�K:�0:	#:ν�93��9㰐9u<9��8$9���۸�O�D���
ȹ5��� S���*�r�A���X��o�1��}z��]���r줺����B��	jƺ��Ѻ�ܺ5�������X���&
�n���1�1��=) ���%��
+�
t0��5�=;��@���E��bK���P��-V���[��a�jxf���k�Leq�$�v�sZ|�(뀻����f���"��
ߋ�����?V������͖�q����  �  d�=p?=U�=׎=
6=��=��=�)=�� =�u =� =��<���<��<jf�<f��<z��<�J�<���<A��<|-�<7x�<���<�<�R�<��<���<$�<�g�<��<9��<i+�<�j�<��<\��<�"�<�]�<��<o��<�<�<�<�o�<���<���<��<�"�<9H�<j�<���<f��<g��<���<	��<o��<���<���<���<]��<���<���<ڶ�<���<&v�<�K�<��<e��<,��<6V�< �<ǫ�<�J�<a��<fp�<���<�w�<=��<�a�<���< 1�<���<e�<8�<���<�ɶ<�	�<�D�<kz�<�<�֭<+��<!�<�@�<�\�<^u�</��<���<��<r��<+͚<g٘<@�<��<B��<B��<2�<��<�
�<��<��<o�<��<�	�<�~<Oz<�u<^�q<��m<8�i<��e<��a<��]<��Y<F�U<��Q<��M<x�I<)�E<b�A<`�=<��9<y�5<��1<��-<q�)<��%<"<�'<�B<'c<�<״<��
<�<C_<�K�;%��;�;�J�;e�;���;���;���;���;�
�;fE�;���;W�;���;(�;�;���;���;#х;�;νt;��i;��^;�:T;!�I;Ͻ?;��5;�(,;A�";ot;�l;a�;���:�#�:>��:��:��:4��:�Þ:�"�:�ρ:ǎg:�K:8�0:|<:	��9U��9���9�;9��8h�>���ܸ�P�n���gȹi�����R�*�mB��
Y��o��G��Z���Pʙ�����&���I��qkƺ,�ѺU�ܺ��纠��	�����n
����%�Ԣ�X ��%���*�Mh0���5��2;�P�@�d�E�.]K�P�P�a,V���[��a�Q}f���k��mq���v�1e|�����®���l��$)���勻Ϡ��\����jҖ������  �  �=$?=�=Î=!6=,�=�=U*=�� =�v =� =��<���<z�<ah�<X��<Z �<dL�< ��<���<�.�<y�<���<r�<S�<���<&��<~#�<�f�<���<���<�)�<�h�<&��<h��<� �<\�<��<���<��<O;�<�n�<؟�<Y��<��<�"�<tH�<�j�<O��<^��<»�<3��<���<M��<���<���<���<B��<���<m��<H��<��<w�<KL�<G�<���<��<�U�<]�<���<eI�<���<�n�<���<�u�<E��<�_�<���<�.�<܌�<��<n6�<3��<eȶ<��<D�<z�<�<"׭<���<:"�<�A�<�]�<�v�<��<���<�<g��<$Ϛ<Pۘ<&�<��<���<���<&�<t�<�<1�<��<�<M�<��<n
~<�z<��u<��q<��m<l�i<��e<��a<��]<9�Y<�U<��Q<�M<v�I<��E<`�A<�=<��9<`�5<\�1<k�-<��)<q&<m"<k+<�F<7g<#�<�<��
<�#<�b<�Q�;L��;���;<N�;]�;���;f��;F��;���;H�;�@�;[��;f��;���;� �;�ݗ;/��;���;�Ʌ;��;=�t;H�i;4�^;�4T;@�I;=�?;D�5;�*,;��";�z;�t;��;��:QA�:���:���:%�:�ح:��:*A�:��:M�g:�)L: 1:�T:t	�9"�9���9��;9!��8q�D���ݸh�P�,Θ���ȹ1d�����!+�LB�rFY��p�Ma�������ޙ�0��e0��5R��pƺ��Ѻߧܺ�级��q���S��<
����$�C��� �/%�|�*�)Y0�=�5�R';�׋@���E�WK�$�P��*V�ݙ[�7a���f���k��vq���v��q|����}���4t��K1��:틻����Bc��S��ؖ�v����  �  ^�=�>=��=��=76=a�=H�=�*=?� =aw =p =ֆ�<���<��<wj�<���<Z�<?N�<Ι�<"��<�/�<z�<r��<��<?S�<���<���<�"�<�e�<j��<!��<(�<�f�<��<R��<��<�Y�<��<���<4�<�9�<�m�<מ�<���<���<�"�<�H�<7k�<4��<���<&��<���<���<2��<���<���<���<\��<w��<2��<׹�<p��<Cx�<(M�<��<���<��<WU�<��<��<!H�<y��<�l�< ��<�s�<��<�]�<m��<�,�<ˊ�<��<�4�<ʀ�<!Ƕ<�<rC�<�y�<���<[׭<c��<#�<
C�<`_�<lx�<͎�<x��<��<uÜ<Bњ<dݘ<�<V�<@��<���<9�<N	�<��<j�<��<��<�
�<��<~<��y<f�u<&�q<��m<D�i<1�e<x�a<��]<w�Y<o�U<½Q<��M<;�I<^�E<a�A<��=<L�9</�5<��1<x�-<��)<�&<�"<H/<�J<�k<u�<^�<�
<g'<+f<X�;���;��;�Q�;<�;���;��;���;���;I�;Q<�;4��;���;cy�;�;�՗;��;ة�;(;��;ɤt;Ҕi;{�^;~-T;��I;��?;��5;C-,;V�";U�;J~;�;W*�:^�:���:/��:�F�:���:b�:c`�:�
�:��g:�WL:�.1:�r: .�9z �9+��9Z�;9�8�rL�;#߸^pQ��=��Bɹ������Qe+�
�B�E�Y�EWp��}������B�T��)>���Z���sƺ��Ѻ¢ܺj�纁��"����z�
�L��T������(n%���*�J0�7�5��;�Հ@���E�ePK�u�P�.)V�H�[��a�x�f�kl�b�q���v��|�L�������k|���9����������j��p$��Aޖ�B����  �  ݕ=c>=��=��=G6=��=��=c+=�� =*x =T =���<���<� �<�l�<���<]�<P�<���<���<$1�<{�<��<5�<GS�<I��<*��<�!�<qd�<��<���<I&�<e�<��<3��<|�<�W�<��<!��<��<v8�<Fl�<��<��<l��<�"�<�H�<�k�<��<���<o��<v��<\��<��<���<���<���<b��<e��<���<���<���<[y�<N�<E�<��<��<�T�<��<٨�<�F�<���<-k�<��<rq�<���<W[�<0��<�*�<���<��<�2�<D�<�Ŷ<��<�B�<Sy�<ת�<�׭<���<$�<"D�<�`�<#z�<���<o��<��<�Ŝ<VӚ<kߘ<��<!�<���<:�<Z�<
�<~�<��<��<?�<�	�<��<u~<��y<��u<f�q<��m<��i<��e<�a<��]<��Y<�U<��Q<ȺM< �I<��E<��A<c�=<�9<�5<m�1<��-<-�)<�&<�"<3<O<�o<�<��<@�
<;+<�i<_^�;��;���;�T�;a�;f��;���;L��;���;r��;?7�;m��;�;Dr�;*�;�͗;*��;���;���;��;s�t;͉i;�^;�&T;L�I;Ѷ?;��5;�/,;�";ȉ;ɇ;Ǻ;9F�:;{�:E�:��:�h�:��:�&�:��:'�:�)h:e�L:1T1:А:�R�9�5�9)��9#�;9�Y�8��S�I\��'R�ߤ����ɹ_��\H�|�+�A�B���Y��p�����َ��	��~/��bL���b���wƺˊѺ��ܺY��2��b���?o���	��v�T���q����v]%���*�;0���5��;�w@���E�JK���P��'V�q�[��a�R�f�Gl��q��w�T�|�����ƃ����,B���������!r��Y+��T䖻�����  �  k�=>=r�=��=]6=��=��=�+=u� =�x = =���<���<�"�<�n�<k��<L�<�Q�<��<���<M2�<�{�<���<��<^S�<��<���<!�<~c�<���<&��<�$�<4c�<��<4��<��<�U�<-��<B��<�<7�<)k�<��<\��<��<�"�<@I�<Il�<���<���<���<���<���<���<���<���<���<4��<E��<���<���<���<^z�<�N�<��<E��<͞�<�T�<5�<���<�E�<k��<�i�<��<so�<���<6Y�<��<�(�<���<�޻<T1�<�}�<�Ķ<"�<B�<�x�<Ǫ�<�׭<e �<�$�<0E�<b�<�{�<7��<S��<淞<�ǜ<B՚<S�<��<���<W��<{�<c�<�
�<�<��<a�<��<-	�<��<~<��y<��u<��q<��m<��i<��e<�a<��]<ºY<��U<ɷQ<9�M<E�I<(�E<��A<��=<��9<�5<��1<��-<��)<�
&<�"<�6<S<�s<�<��<J�
<�.<5m<Nd�;)��;���;nW�;��;3��;W��;���;U��;��;[2�;'��;��;k�;�	�;Ɨ;���;.��;���;]�;�t;.i;��^;� T;�I;��?;X�5;�2,;��";~�;t�;m�;O^�:���:3�:�.�:8��:�<�:gD�:۞�:{A�:�Yh:߬L:�v1:��:�u�9�J�98��9=`;9(��8�Y��h�D�R�����-ʹ
�������+�dC��Z�]�p���������?���>��KX��|l��E{ƺ'�Ѻ"�ܺq��=��l���\d���	�Fi�����b����N%�X�*�=,0�Q�5�t;�"m@���E�-EK�~�P�&V���[��a�\�f� l�z�q�w��|�N��΃�،��	J�����T����y���1���閻�����  �  ��=�==C�=}�=d6=�=H�=F,=�� =}y =� =���<5��<>$�<Mp�<��<��<@S�<t��</��<Q3�<�|�<J��<��<eS�<��<3��<a �<�b�<���<���<'#�<�a�<|��<���<��<1T�<���<���<���<�5�<%j�<D��<���<���<�"�<XI�<�l�<v��<���<���<)��<`��<y��<��<B��<���<���<���<���<3��<��<A{�<[O�<2�<U��<���<IT�<��<��<�D�<"��<!h�<���<�m�<���<aW�<=��<�&�< ��<jݻ<�/�<�|�<�ö<L�<�A�<�x�<���<ح<� �<o%�<F�<%c�<�|�<���<է�<���<>ɜ<�֚<��<=�<��<���<��<<�<u�<g�<��<O�<��<��<��<� ~<:�y<��u<��q<��m<��i<j�e<��a<y�]<зY<��U<$�Q<
�M<c�I<�E<��A<��=<��9<��5<��1<7�-<��)< &<�!"<�9<EV<>w<��<��<��
<�1<	p<xi�;� �;ܥ�;9Z�;��;���;��;D��;���;���;\.�;I|�;Y�;�e�;��;���;���;ד�;���;}�;��t;�ui; �^;�T;H�I;ز?;��5;�3,;��";��;�;��;�r�:¬�:<K�:�H�:���:XW�:l^�::��:�X�:��h:h�L:��1:K�:���9S�9��9�@;9l'�89m`�i�orS�0Z��3�ʹ�8��Ϻ��,��HC�=Z�y q�̓�%��"1��N��d���s��E~ƺ�Ѻ�ܺ��c�򺛮���Z�7�	��]�����U�?���@%�Ա*�� 0�>�5���:�\d@���E��?K���P��%V�G�[�wa��f�/l�ܜq�%!w�1�|���xԃ�����Q������Ǝ�y��z7��Ϧ���  �  ��=�==�=k�=t6=!�=��=�,=[� =�y =]  ='��<{��<�%�<�q�<i��<	�<sT�<���<��<4�<7}�<���<�<{S�<���<���<��<�a�<٢�<���<	"�<y`�<��</��<r�<�R�<O��<���<���<�4�<ji�<���<���<t��<�"�<}I�<�l�<��<)��<���<#��<���<���<w��<���<���<$��<���<��</��<Ѡ�<�{�<�O�<q�<p��<���<�S�<C�<q��<�C�<>��<�f�<[��<ql�<���<�U�<���<O%�<ǃ�<6ܻ<�.�<�{�<�¶<��<&A�<\x�<���<,ح<6�<�%�<�F�<�c�<�}�<ʔ�<��<ݺ�<{ʜ<.ؚ<1�<q�<G��<���<Y�<��<��<��<�<<�<+�<A�<I�<��}<`�y<��u<X�q<�m<��i<��e<��a<��]<\�Y<k�U<(�Q<~�M< �I<
�E<��A<f�=<�9<�5<��1<G�-<C�)<�&<�#"<9<<�X<�y<�<��<�
<{4<Xr<m�;��;=��;\�;��;W��;t��;%��;Z��;)��;�+�;hx�;'ߪ;�`�;���;���;�;���;���;��;,zt;�oi;��^;�T;+�I;S�?;��5;E5,;	�";��;͜;��;҂�:���:i^�:}^�:��:�k�:yt�:Dʐ:�k�:*�h:g�L:��1:�:z��93]�9�9;9�ܫ8f"e��#��S����F�ʹ��������H,�sC�iZ��(q��ރ�6���=���Y��gl���x��ÂƺވѺR�ܺS����֣��zT���	�(T�����J�B���6%�]�*��0���5�Y�:�h^@���E��;K�ȮP��$V���[��a��f�bl�ɢq��(w���|�����ك�����MV����̎�G����;����ͩ���  �  h�=S==��=e�={6=3�=��=�,=�� =7z =�  =э�<5��<P&�<`r�<"��<�	�<U�<��<���<�4�<�}�<���<2�<�S�<���<���<��<_a�<=��<.��<Z!�<�_�<g��<a��<��<R�<���<���<���<Z4�<�h�<;��<0��<O��<�"�<�I�</m�<C��<���<.��<���<"��<U��<'��<P��<���<���<���<���<���<e��<V|�<!P�<��<���<���<�S�<� �<���<7C�<���<Lf�<���<�k�<���<U�<���<�$�<��<wۻ<.�<{�<b¶<C�<�@�<7x�<���<Dح<a�<F&�<AG�<{d�<v~�<c��<���<���<J˜<�ؚ<��<�<���<��<��<I	�<:�<��<*�<3�<�<��<��<f�}<�y<��u<��q<��m<I�i<�e<f�a<B�]<ݳY<�U<߱Q<O�M<�I<J�E<��A<I�=<4�9<^�5<T�1<B�-<n�)<&<%"<�=<bZ<�{<ס<C�<��
<�5<�s<�o�;�;3��;$]�;��;���;Q��;m��;���;o��;Q)�;v�;�ܪ;^�;���;w��;ӑ�;Ջ�;ѥ�;b�;�ut;�ji;ҟ^;�T;��I;c�?;��5;!6,;��";h�;��;��;<��:���:�i�:�i�:%Ž:�x�:��:�Ր:�u�:��h:��L:Z�1:d�:S��9�c�9ð�9�;9a��8�^h����,T��ǚ���ʹ۹�����c,��C��Z��?q�
ꃺ$!���G���a���r���|��Z�ƺ9�Ѻ7�ܺ�纜��=����O�"�	�7O�@��%E����W0%���*��0�T5���:��Y@���E��9K���P��#V�Z�[��a�ǝf��!l�8�q��-w�	�|�����܃�����Y�����Ύ�6���z>��b�������  �  a�=E==��=b�=s6==�=��=�,=�� =Oz =�  =+��<���<�&�<�r�<`��<(
�<nU�<`��<���<�4�<�}�<��<@�<tS�<���<���<k�<Ra�<��<��<!�<i_�<��<��<N�<�Q�<=��<���<���<#4�<�h�<.��<��<\��<�"�<�I�<Qm�<]��<���<L��<���<w��<���<f��<���<���<��<��<��<���<���<_|�<6P�<��<}��<���<�S�<� �<��<"C�<T��<f�<D��<Mk�<m��<�T�<���<7$�<���<&ۻ<�-�<�z�<P¶<&�<�@�<7x�<���<Hح<~�<Z&�<FG�<�d�<�~�<���<��<ͻ�<�˜<8ٚ<3�<|�<)��<H��<�<]	�<Y�<��<�<)�<�<��<��<2�}<��y<�u<'�q<��m<��i<j�e<��a<��]<%�Y<��U<z�Q<�M<��I<�E<��A<=�=<�9<��5<��1<j�-<��)<v&<�%"<M><
[<|<{�<��<]�
<�6<t<Kp�;8�;���;�]�;��;z��;\��;W��;���;L��;�(�;�u�;�۪;�\�;���;5��;���;���;x��;ʽ;tt;ii;Q�^;�T;��I;ٯ?;\�5;�5,;��";F�;��;��;��:��:Jp�:�m�:�ɽ:�}�:o��:,ܐ:{�:�h:�M:ʺ1:O�:;��9c�9n��9�	;9ur�8J�h�r���GT��Қ��˹�����m,�ΗC�щZ��Jq���#��J��fb��9t���}���ƺF�Ѻܺ��+�򺳚��~N��	�^L�$��.C�)��%.%�R�*��0��|5�$�:�-Y@��E��8K���P�S$V���[�ja���f�<"l��q�H/w���|���	ރ�T����Z��r��CЎ�����}?��%��������  �  h�=S==��=e�={6=3�=��=�,=�� =7z =�  =э�<5��<P&�<`r�<"��<�	�<U�<��<���<�4�<�}�<���<2�<�S�<���<���<��<_a�<=��<.��<Z!�<�_�<g��<a��<��<R�<���<���<���<Z4�<�h�<;��<0��<O��<�"�<�I�</m�<C��<���<.��<���<"��<U��<'��<P��<���<���<���<���<���<e��<V|�<!P�<��<���<���<�S�<� �<���<7C�<���<Lf�<���<�k�<���<U�<���<�$�<��<wۻ<.�<{�<b¶<C�<�@�<7x�<���<Dح<a�<F&�<AG�<{d�<v~�<c��<���<���<J˜<�ؚ<��<�<���<��<��<I	�<:�<��<*�<2�<�<��<��<f�}<�y<��u<��q<��m<I�i<�e<f�a<B�]<ݳY<�U<߱Q<O�M<�I<J�E<��A<I�=<4�9<^�5<T�1<C�-<n�)<&<%"<�=<bZ<�{<ס<C�<��
<�5<�s<�o�;�;3��;$]�;��;���;P��;m��;���;o��;Q)�;v�;�ܪ;^�;���;w��;ӑ�;Ջ�;ѥ�;b�;�ut;�ji;ҟ^;�T;��I;c�?;��5;!6,;��";h�;��;��;<��:���:�i�:�i�:%Ž:�x�:��:�Ր:�u�:��h:��L:Z�1:d�:S��9�c�9ð�9�;9a��8�^h����,T��ǚ���ʹ۹�����c,��C��Z��?q�
ꃺ$!���G���a���r���|��Z�ƺ9�Ѻ7�ܺ�纜��=����O�"�	�7O�@��%E����W0%���*��0�T5���:��Y@���E��9K���P��#V�Z�[��a�ǝf��!l�8�q��-w�	�|�����܃�����Y�����Ύ�6���z>��b�������  �  ��=�==�=k�=t6=!�=��=�,=[� =�y =]  ='��<{��<�%�<�q�<i��<	�<sT�<���<��<4�<7}�<���<�<{S�<���<���<��<�a�<٢�<���<	"�<y`�<��</��<r�<�R�<O��<���<���<�4�<ji�<���<���<t��<�"�<}I�<�l�<��<)��<���<#��<���<���<w��<���<���<$��<���<��</��<Ѡ�<�{�<�O�<q�<p��<���<�S�<C�<q��<�C�<>��<�f�<[��<ql�<���<�U�<���<O%�<ǃ�<6ܻ<�.�<�{�<�¶<��<&A�<\x�<���<,ح<6�<�%�<�F�<�c�<�}�<ʔ�<��<ݺ�<{ʜ<.ؚ<1�<q�<G��<���<Y�<��<��<��<�<<�<+�<A�<I�<��}<`�y<��u<X�q<�m<��i<��e<��a<��]<\�Y<k�U<(�Q<~�M< �I<�E<��A<f�=<�9<�5<��1<G�-<C�)<�&<�#"<9<<�X<�y<�<��<�
<{4<Xr<m�;��;=��;\�;��;V��;t��;%��;Y��;)��;�+�;hx�;'ߪ;�`�;���;���;�;���;���;��;,zt;�oi;��^;�T;+�I;S�?;��5;E5,;	�";��;͜;��;҂�:���:i^�:}^�:��:�k�:yt�:Dʐ:�k�:*�h:g�L:��1:~�:z��93]�9�9;9�ܫ8f"e��#��S����F�ʹ��������H,�sC�iZ��(q��ރ�6���=���Y��gl���x��ÂƺވѺR�ܺS����֣��zT���	�(T�����J�B���6%�]�*��0���5�Y�:�h^@���E��;K�ȮP��$V���[��a��f�bl�ɢq��(w���|�����ك�����MV����̎�G����;����ͩ���  �  ��=�==C�=}�=d6=�=H�=F,=�� =}y =� =���<5��<>$�<Mp�<��<��<@S�<t��</��<Q3�<�|�<J��<��<eS�<��<3��<a �<�b�<���<���<'#�<�a�<|��<���<��<1T�<���<���<���<�5�<%j�<D��<���<���<�"�<XI�<�l�<v��<���<���<)��<`��<y��<��<B��<���<���<���<���<3��<��<A{�<[O�<2�<U��<���<IT�<��<��<�D�<"��<!h�<���<�m�<���<aW�<=��<�&�< ��<jݻ<�/�<�|�<�ö<L�<�A�<�x�<���<ح<� �<o%�<F�<%c�<�|�<���<է�<���<>ɜ<�֚<��<=�<��<���<��<<�<u�<g�<��<O�<��<��<��<� ~<:�y<��u<��q<��m<��i<j�e<��a<y�]<зY<��U<$�Q<
�M<c�I<�E<��A<��=<��9<��5<��1<7�-<��)< &<�!"<�9<EV<>w<��<��<��
<�1<	p<xi�;� �;ܥ�;9Z�;��;���;��;D��;���;���;\.�;H|�;Y�;�e�;��;���;���;ד�;���;|�;��t;�ui; �^;�T;H�I;ز?;��5;�3,;��";��;�;��;�r�:¬�:<K�:�H�:���:XW�:l^�::��:�X�:��h:h�L:��1:K�:���9S�9��9�@;9l'�89m`�i�orS�0Z��3�ʹ�8��Ϻ��,��HC�=Z�y q�̓�%��"1��N��d���s��E~ƺ�Ѻ�ܺ��c�򺛮���Z�7�	��]�����U�?���@%�Ա*�� 0�>�5���:�\d@���E��?K���P��%V�G�[�wa��f�/l�ܜq�%!w�1�|���xԃ�����Q������Ǝ�y��z7��Ϧ���  �  k�=>=r�=��=]6=��=��=�+=u� =�x = =���<���<�"�<�n�<k��<L�<�Q�<��<���<M2�<�{�<���<��<^S�<��<���<!�<~c�<���<&��<�$�<4c�<��<4��<��<�U�<-��<B��<�<7�<)k�<��<\��<��<�"�<@I�<Il�<���<���<���<���<���<���<���<���<���<4��<E��<���<���<���<^z�<�N�<��<E��<͞�<�T�<5�<���<�E�<k��<�i�<��<so�<���<6Y�<��<�(�<���<�޻<T1�<�}�<�Ķ<"�<B�<�x�<Ȫ�<�׭<e �<�$�<0E�<b�<�{�<7��<S��<淞<�ǜ<B՚<S�<��<���<W��<z�<c�<�
�<�<��<a�<��<-	�<��<~<��y<��u<��q<��m<��i<��e<�a<��]<ºY<��U<ɷQ<9�M<F�I<)�E<��A<��=<��9<�5<��1<��-<��)<�
&<�"<�6<S<�s<�<��<J�
<�.<5m<Md�;)��;���;nW�;��;2��;W��;���;U��;��;Z2�;'��;��;k�;�	�;Ɨ;���;.��;���;\�;�t;-i;��^;� T;�I;��?;X�5;�2,;��";~�;t�;m�;O^�:���:3�:�.�:8��:�<�:gD�:۞�:{A�:�Yh:߬L:�v1:��:�u�9�J�98��9=`;9(��8�Y��h�D�R�����-ʹ
�������+�dC��Z�]�p���������?���>��KX��|l��E{ƺ'�Ѻ"�ܺq��=��l���\d���	�Fi�����b����N%�X�*�=,0�Q�5�t;�"m@���E�-EK�~�P�&V���[��a�\�f� l�z�q�w��|�N��΃�،��	J�����T����y���1���閻�����  �  ݕ=c>=��=��=G6=��=��=c+=�� =*x =T =���<���<� �<�l�<���<]�<P�<���<���<$1�<{�<��<5�<GS�<I��<*��<�!�<qd�<��<���<I&�<e�<��<3��<|�<�W�<��<!��<��<v8�<Fl�<��<��<l��<�"�<�H�<�k�<��<���<o��<v��<\��<��<���<���<���<b��<e��<���<���<���<[y�<N�<E�<��<��<�T�<��<٨�<�F�<���<.k�<��<rq�<���<W[�<0��<�*�<���<��<�2�<D�<�Ŷ<��<�B�<Sy�<ת�<�׭<���<$�<"D�<�`�<#z�<���<o��<��<�Ŝ<VӚ<kߘ<��<!�<���<:�<Z�<
�<~�<��<��<>�<�	�<��<u~<��y<��u<f�q<��m<��i<��e<�a<��]<��Y<�U<��Q<ɺM< �I<��E<��A<c�=<�9<�5<m�1<��-<-�)<�&<�"<3<O<�o<�<��<@�
<;+<�i<^^�;��;���;�T�;`�;f��;���;K��;���;r��;?7�;m��;�;Cr�;)�;�͗;)��;���;���;��;s�t;̉i;�^;�&T;L�I;Ѷ?;��5;�/,;�";ȉ;ȇ;Ǻ;9F�:;{�:E�:��:�h�:��:�&�:��:'�:�)h:e�L:1T1:А:�R�9�5�9)��9#�;9�Y�8��S�I\��'R�ߤ����ɹ_��\H�|�+�A�B���Y��p�����َ��	��~/��bL���b���wƺˊѺ��ܺY��2��b���?o���	��v�T���q����v]%���*�;0���5��;�w@���E�JK���P��'V�q�[��a�R�f�Gl��q��w�T�|�����ƃ����,B���������!r��Y+��T䖻�����  �  ^�=�>=��=��=76=a�=H�=�*=?� =aw =p =ֆ�<���<��<wj�<���<Z�<?N�<Ι�<"��<�/�<z�<r��<��<?S�<���<���<�"�<�e�<j��<!��<(�<�f�<��<R��<��<�Y�<��<���<4�<�9�<�m�<מ�<���<���<�"�<�H�<7k�<4��<���<&��<���<���<2��<���<���<���<\��<w��<2��<׹�<p��<Cx�<(M�<��<���<��<WU�<��<��<!H�<z��<�l�< ��<�s�<��<�]�<m��<�,�<ˊ�<��<�4�<ʀ�<"Ƕ<�<rC�<�y�<���<[׭<c��<#�<
C�<`_�<lx�<͎�<x��<��<uÜ<Bњ<dݘ<�<V�<?��<���<9�<N	�<��<j�<��<��<�
�<��<~<��y<f�u<%�q<��m<D�i<1�e<x�a<��]<w�Y<o�U<½Q<��M<;�I<_�E<b�A<��=<L�9</�5<��1<x�-<��)<�&<�"<H/<�J<�k<u�<^�<�
<g'<+f<X�;���;��;�Q�;;�;���;��;���;���;H�;P<�;3��;���;by�;�;�՗;��;ة�;(;��;Ȥt;єi;{�^;}-T;��I;��?;��5;C-,;U�";U�;J~;�;V*�:^�:���:/��:�F�:���:b�:c`�:�
�:��g:�WL:�.1:�r: .�9z �9+��9Z�;9�8�rL�;#߸^pQ��=��Bɹ������Qe+�
�B�E�Y�EWp��}������B�T��)>���Z���sƺ��Ѻ¢ܺj�纁��"����z�
�L��T������(n%���*�J0�7�5��;�Հ@���E�ePK�u�P�.)V�H�[��a�x�f�kl�b�q���v��|�L�������k|���9����������j��p$��Aޖ�B����  �  �=$?=�=Î=!6=,�=�=U*=�� =�v =� =��<���<z�<ah�<X��<Z �<dL�< ��<���<�.�<y�<���<r�<S�<���<&��<~#�<�f�<���<���<�)�<�h�<&��<h��<� �<\�<��<���<��<O;�<�n�<؟�<Y��<��<�"�<tH�<�j�<O��<^��<»�<3��<���<M��<���<���<���<B��<���<m��<H��<��<w�<KL�<G�<���<��<�U�<]�<���<eI�<���<�n�<���<�u�<E��<�_�<���<�.�<܌�<��<n6�<3��<eȶ<��<D�<z�<�<"׭<���<;"�<�A�<�]�<�v�<��<���<�<g��<$Ϛ<Pۘ<&�<��<���<���<%�<t�<�<1�<��<�<M�<��<n
~<�z<��u<��q<��m<l�i<��e<��a<��]<:�Y<�U<��Q<	�M<v�I<��E<a�A<�=<��9<`�5<\�1<k�-<��)<q&<m"<k+<�F<7g<#�<�<��
<�#<�b<�Q�;L��;���;;N�;]�;���;f��;F��;���;H�;�@�;[��;e��;���;� �;�ݗ;/��;���;�Ʌ;��;<�t;G�i;3�^;�4T;?�I;=�?;D�5;�*,;��";�z;�t;��;��:QA�:���:���:%�:�ح:��:*A�:��:M�g:�)L: 1:�T:t	�9"�9���9��;9!��8q�D���ݸh�P�,Θ���ȹ1d�����!+�LB�rFY��p�Ma�������ޙ�0��e0��5R��pƺ��Ѻߧܺ�级��q���S��<
����$�C��� �/%�|�*�)Y0�=�5�R';�׋@���E�WK�$�P��*V�ݙ[�7a���f���k��vq���v��q|����}���4t��K1��:틻����Bc��S��ؖ�v����  �  d�=p?=U�=׎=
6=��=��=�)=�� =�u =� =��<���<��<jf�<f��<z��<�J�<���<A��<|-�<7x�<���<�<�R�<��<���<$�<�g�<��<9��<i+�<�j�<��<\��<�"�<�]�<��<o��<�<�<�<�o�<���<���<��<�"�<9H�<j�<���<f��<g��<���<	��<o��<���<���<���<]��<���<���<ڶ�<���<&v�<�K�<��<e��<,��<6V�< �<ǫ�<�J�<a��<fp�<���<�w�<=��<�a�<���< 1�<Ꮍ<e�<8�<���<�ɶ<�	�<�D�<kz�<�<�֭<+��<!�<�@�<�\�<^u�</��<���<��<r��<+͚<g٘<@�<��<A��<B��<2�<��<�
�<��<��<o�<��<�	�<�~<Oz<�u<^�q<��m<8�i<��e<��a<��]<��Y<F�U<��Q<��M<y�I<)�E<b�A<`�=<��9<z�5<��1<��-<q�)<��%<"<�'<�B<'c<�<״<��
<�<C_<�K�;$��;�;�J�;d�;���;���;���;���;�
�;eE�;���;W�;���;(�;�;���;���;#х;�;νt;��i;��^;�:T;!�I;Ͻ?;��5;�(,;A�";ot;�l;a�;���:�#�:>��:��:��:4��:�Þ:�"�:�ρ:ǎg:�K:8�0:|<:	��9U��9���9�;9��8h�>���ܸ�P�n���gȹi�����R�*�mB��
Y��o��G��Z���Pʙ�����&���I��qkƺ,�ѺU�ܺ��纠��	�����n
����%�Ԣ�X ��%���*�Mh0���5��2;�P�@�d�E�.]K�P�P�a,V���[��a�Q}f���k��mq���v�1e|�����®���l��$)���勻Ϡ��\����jҖ������  �  Ɨ=�?=z�=܎=�5=��=1�=k)=h� =Fu = =���<'��<��<�d�<���<���<I�<+��< ��<s,�<Yw�<o��<�
�<�R�<��<��<�$�<�h�<��<u��<�,�<4l�<���<���<c$�<}_�<x��<���<��<�=�<�p�<^��<x��<���<�"�<H�<�i�<Ӈ�<l��<F��<q��<���<���<��<���<-��<���<;��<?��<���<���<3u�<�J�<;�<:��<?��<lV�<��<���<�K�<���<�q�<9��<Ly�<���<�c�<���<�2�<w��<��<^9�<Մ�<�ʶ<�
�<CE�<�z�<���<�֭<���<� �<�?�<t[�<t�<ʉ�<)��<\��<���<{˚<�ט<��<t�<���<)��<:�<��<�
�<��<��<��<y�<O
�<�~<�z<��u<J�q<��m<��i<�e<��a<��]<��Y<�U<]�Q<��M<�I<�E<�A<��=<r�9<��5<��1<��-<K�)<��%<1"<�$<�?<�_<r�<T�<��
<�<R\<VF�;���;��;6H�;��;"��;���;��;��;��;vI�;I��;��;��; .�;H�;OƑ;�;�օ;��;��t;U�i;��^;@T;<�I;ľ?;��5;�&,;1�";n;bd;�;��:'�:���:s��:�:���:p��:g
�:(��:�cg:N�K:�0:	#:ν�93��9㰐9u<9��8$9���۸�O�D���
ȹ5��� S���*�r�A���X��o�1��}z��]���r줺����B��	jƺ��Ѻ�ܺ5�������X���&
�n���1�1��=) ���%��
+�
t0��5�=;��@���E��bK���P��-V���[��a�jxf���k�Leq�$�v�sZ|�(뀻����f���"��
ߋ�����?V������͖�q����  �  	�=�?=��=�=�5=��=��=)=� =�t =} =e��<���<|�<Zc�<_��<���<�G�<��<��<�+�<�v�<��<\
�<�R�<$��<H��<I%�<i�<ë�<c��<�-�<gm�<��<I��<�%�<�`�<���<��<�	�<�>�<rq�<��<���<���<�"�<�G�<Li�<J��<���<~��<`��<���<���<���<���<���<d��<���<%��<}��<ӗ�<�t�<TJ�<��<���<T��<�V�<��<.��<TL�<x��<�r�<|��<�z�<l��<e�<���<!4�<���</�<k:�<���<0˶<"�<�E�<�z�<	��<]֭<s��<& �<"?�<�Z�<�r�<���<ܛ�<��<j��<*ʚ<p֘<��<T�<��<d��<��<��<&
�<��<��<��<��<�
�<5~<e	z<�v<��q<m�m<D�i<��e<��a<��]<Q�Y<Z�U<!�Q</�M<.�I<m�E<}�A<��=<%�9<��5<��1<d�-<��)<��%<�"<"<�<<�\<��<��<��
<<�Y<oB�;f��;��;|F�;��;���;��;���;���;��;/L�;���;��;���;3�;5�;ˑ;.ċ;�ۅ;�;��t;R�i;��^;�CT;��I;ҿ?;��5;�#,;t�";�i;]^;��;���:���:/��:&}�:�Ӽ:@��:O��:���:��:�@g:a�K:v�0:�:ª�9���9���9�#<9K�8�5�|Q۸$O��ڗ���ǹ:<��='���*�j�A���X��o�!���j��C���[㤺����>���gƺ�Ѻ��ܺY���%��A��N/
����8<�����3 �1�%��+��}0� �5�1E;� �@�tF�fK�v�P�C/V��[�a�,uf�{�k��_q���v��Q|�`总�����`������ً�����wQ��-��ʖ������  �  H�=@=��=�=�5=x�=͂=�(=�� =xt =) =��<��<��<�b�<���<���<0G�<r��<v��<*+�<Ev�<���<5
�<�R�<9��<s��<�%�<�i�<Y��<���<�.�<n�<���<��<t&�<�a�<a��<���<k
�<;?�<�q�<E��<��<���<�"�<�G�<
i�<��<<��<޷�<���<���<���<���<���<��<���<C��<u��<��<5��<t�<�I�<��<���<_��<�V�<7�<���<�L�<��<~s�<#��<Q{�<)��<�e�<���<�4�<|��<��<;�<P��<�˶<~�<�E�<�z�<
��<B֭<#��<��<�>�<Z�<_r�<���<'��<K��<���<_ɚ<�՘<���<��<H�<���<�<�<�	�<��<��<��<�<J�<S~<�
z<v<��q<��m<��i<;�e<�a<�]<��Y<��U<R�Q<\�M<.�I<��E<��A<��=<�9<��5<�1<y�-<��)<��%<�
"<� <H;<P[<�<��<W�
<�<�X<�?�;��;&��;�D�;�;5��;6��;,��;���;��;YN�;ס�;#�;6��;�5�;1�;-Α;�Ƌ;;ޅ;c�;��t;޼i;��^;�FT;�I;��?;��5;�",;5�";Bf;uZ;e�;i��:���:�~�:�q�:�Ƽ:z�:���:�:���:�,g:٨K:1�0:�:�9D��9D��9�1<9P�8�=2���ڸ�N�1����ǹb��L��i*���A�E�X��qo�����a��Ѣ��Uۤ�����;��kfƺ��ѺA�ܺ����	�.��\��54
�R���A����W: ���%�F+���0�_�5�4J;�ҩ@�1	F�0iK�(�P��/V���[��a�Lsf���k�9[q���v�M|��〻�����]��2���֋������N���
���ǖ�G����  �  G�=�<=��=��=31=�=�}=X#=�� =qn =� =,r�<ļ�<a�<R�<���<e��<�1�<m|�<���<�<*Y�<_��<���<V/�<�t�<��<2��<->�<�<Ⱦ�<]��<�:�<w�<,��<��<�$�<�[�<'��<���<���<B&�<�S�<J~�< ��<��<���<T�<\&�<�=�<�Q�<�a�<�m�<v�<z�<�y�<�t�<`k�<�\�<�H�<)/�<y�<���<��<f��<�N�<��<��<�q�<��<n��<GP�<���<�i�<w��<%f�<��<%G�<ڭ�<4�<ah�<���<�<�S�<4��<Xղ<G�<uB�<r�<��<Nĩ<��<��<�$�<�>�<V�<gk�<�~�<c��<i��<�<)��<Ȓ<�Ґ<�ێ<��<��<`��<��<*��<���<���<;�}<��y<	�u<��q<��m<�i<=�e<��a<�]<�Y<9�U<K�Q<Y�M<�J<9
F<�B<�><e%:<�16<�?2<QP.<�c*<z&<,�"<g�<\�<m�<+<�^<T�<��<�<n <׆�;�@�;_	�;���;H��; ��;���;���;R)�;hs�;�Գ;YM�;1ߦ;?��;$R�;s5�;5�;HR�;���;��y;F�n;J�c;0>Y;��N;��D;�:;U1;�|';.;�;=/;~;���:�a�:9'�:�J�:2ȵ:���:���:V4�:_�u:�Y:�I>:%+#:~q:G)�9�9�-i9j\9���7ܴ��kE(�� ��2��� ��q�
�-{"�2�9�xOQ�1|h����Z8��&��������Q��b�����ú�+Ϻ�lں*��l�����3��j;	�3��Z�c���e���$��\*���/�'C5���:�T@�n�E���J�UfP�*�U��H[���`�;5f��k��,q�f�v��)|�Հ������U��U���Ջ�A����U�����ז�o����  �  ?�=�<=��=��=21=��=�}=e#=� =}n =� =gr�<���<��<AR�<���<���<42�<�|�<���<<�<CY�<���<���<W/�<�t�<���<��<#>�<�~�<���<,��<�:�<�v�<���<���<^$�<u[�<���<���<���<?&�<sS�<(~�<��<��<���<d�<u&�<�=�<�Q�<�a�<n�<Mv�<Vz�<z�<:u�<�k�<�\�<�H�<=/�<��<���<���<z��<�N�<��<��<�q�<��<f��<1P�<���<xi�</��<�e�<���<�F�<���<��</h�<r��<�
�<�S�<��<9ղ<>�<qB�<�q�<@��<cĩ<��<��<�$�<�>�<IV�<�k�<�<���<���</��<U��<'Ȓ<�Ґ<܎<�<��<[��<��<��<i��<���<;�}<T�y<��u<d�q<�m<��i<��e<?�a<��]<��Y<��U<��Q<V�M<�J<
F<�B<�><`%:<�16<�?2<�P.<�c*<Nz&<~�"<�<��<��<{+<_<˘<�<! <Qn <W��;A�; 
�;���;Z��;&��;3��;n��;6)�;Zs�;�ӳ;�L�;(ަ;>��;hQ�;�4�;?4�;?Q�;֋�;��y;��n;D�c;�=Y;��N;��D;d�:;)1;Q}';�.;c;g0;�~;- �:Se�:+�:�N�:7̵:ş�:aŗ:�7�:�u::�Y:�L>:�-#:Ct:D'�9��9,(i9iK9���7^���4O(�+��쿵�����
���"��:��WQ�>�h�X���:��¡��E���S�����G�ú�+Ϻ�lں��������K���:	�v��^X�q���c���$�[*��/��A5��:�2@���E���J��eP�U�U��H[�0�`�6f�|�k��,q�x�v��*|��Հ����PV��<��a֋�Q���rV������ז�p����  �  �=�<=��=��=<1=��=�}=�#=;� =�n =  =�r�<���<8�<�R�<���<)��<�2�<}�<��<��<�Y�<á�< ��<f/�<�t�<ٸ�<���<�=�<�~�<��<���<:�<Uv�<j��<;��<�#�<�Z�<|��<A��<��<�%�<+S�<~�<���<��<���<��<�&�<L>�<HR�<Zb�<�n�<�v�<�z�<�z�<�u�<)l�<~]�<yI�<�/�<�<���<A��<���<�N�<��<���<�q�<��<���<�O�<���<�h�<���<Te�<��<OF�<��<_�<�g�<껹<|
�<cS�<ݖ�<ղ<-�<sB�<
r�<p��<�ĩ<*�<<�<%�<A?�<�V�<9l�<��<:��</��<���<ڼ�<�Ȓ<)Ӑ<M܎<K�<��<p��<��<���<C��<���<q�}<W�y<��u<j�q<��m<��i<p�e<&�a<p�]<��Y<��U<��Q<��M<�J<�	F<�B<�><�%:<�16<n@2<Q.<�d*<E{&<��"<��<��<(�<�,<J`<�<H�<4!<[o <"��;9B�; �;c��;���;0��;���;���;�'�;�q�;ҳ;�J�;Uܦ;E��;EO�;,2�;42�;8O�;��;��y;��n;O�c;�;Y;z�N;)�D;ּ:;1;�~'; 1;E;K4;��;��:Dn�:'4�:X�:xյ:㨦:7Η:Q@�:��u:��Y:�X>:�6#:�z:U-�9��9:!i9�79��7����(��J�� ߵ�c���
� �"�,:�vhQ��h����B������5���V��p�����ú.+Ϻ�kں�庽����\���6	���T�����^���$��V*���/��=5��:��@�Z�E���J��dP���U��H[��`�F7f���k��/q�i�v��.|��׀�6���yX������؋�o���eX������ٖ�����  �  ݔ=]<=��=��=I1=��=�}=�#=�� =o =� =�s�<���<4	�<�S�<���<#��<�3�<�}�<���</�<Z�<	��<K��<q/�<�t�<���<���<N=�<�}�<|��<���</9�<cu�<k��<F��<�"�<Z�<���<���<}��<M%�<�R�<�}�<إ�<��< ��<��<'�<�>�<�R�<(c�<mo�<�w�<�{�<�{�<�v�<%m�<l^�<BJ�<�0�<��<t��<���<ۉ�<�N�<��<���<Qq�<+�<b��<O�<8��<�g�<���<Ed�<��<AE�<���<q�<�f�<2��<�	�<�R�<s��<�Բ< �<iB�<Gr�<���<ũ<��<��<�%�<@�<�W�<1m�<���<6��</��<���<���<fɒ<�Ӑ<�܎<��<A�<���<��<���<���<$��<H�}<%�y<&�u<��q<�m<��i<��e<�a<��]<��Y<5�U<��Q<F�M<�J<	F<B<�><�%:<z26<A2<R.<�e*<�|&<4�"<ε<��<0<�.<Rb<��<�<�"<�p <}��;jD�;q�;���;!��;���;+��;���;>&�;�o�;�ϳ;�G�;٦;���;|K�;�.�;a.�;�K�;���;F�y;��n;1�c;�8Y;��N;:�D;n�:;�1;�';f4;�;�8;M�;��:_}�:MD�:Th�:��: ��:�ݗ:JM�:�v:��Y:�i>:0D#:U�:=�9��9�i9�92 �7]���v�(�x��[���C湵��"��4:�G�Q���h�(��OM��L���&��2\�������ú�*Ϻ�fں��9����H���/	����AL�����V���$��N*�|�/�075���:�@�&�E���J��bP���U�rI[�{�`��9f�>�k�v4q�-�v�!5|�Zۀ�⛃�~\������܋�%����[�����ܖ�q����  �  ��=<={�=��=Q1=��=~=&$=�� =�o = =�t�<ƿ�<l
�<"U�<���<_��<�4�<�~�<���<��<�Z�<q��<���<w/�<t�<W��<��<�<�<!}�<���<���<8�<%t�<+��<��<�!�<�X�<���<���<���<�$�<?R�<F}�<���<���<F��<#�<�'�<�?�<�S�<!d�<�p�<�x�<}�<�|�<x�<Sn�<�_�<TK�<|1�<q�<(��<(��<(��<O�<��<���<�p�<��<���<N�<.��<�f�<w��<�b�<���<�C�<���<:�<�e�<1��<��<R�<ו�<XԲ<��<\B�<tr�<���<�ũ<^�<�	�<�&�<"A�<�X�<_n�<ځ�<p��<h��<α�<���<_ʒ<�Ԑ<�ݎ<!�<��<���<��<���<x��<���<��}<^�y<�u<i�q<��m<�i< �e<��a<�]<��Y<�U<��Q<��M<� J<�F<�B<{><�%:<�26<�A2<�S.<ag*<�~&<\�"<,�<��<�<s1<�d<��<l�<.%<�r <ӎ�;aG�;[�;	��;���;���;F��;���;
$�;�l�;a̳;�C�;�Ԧ;��;�F�;*�;�)�;vG�;���;��y;�n;��c;�4Y;A�N;i�D;��:;l1;�';�8;�";�?;V�;�'�:Ԑ�:�W�:P|�:���:`̦:�:�^�:�,v:�Z:��>:eV#:~�:I�9��9� i9��9��7�V��MD)�̵��l\��\��o-���"��\:�4�Q���h�k��\��ڿ������d������J�ú�*Ϻcں�������� ���'	����xB�H���L�
�$��D*�(�/��.5�G�:��@�U~E�$�J�V`P���U��I[���`��=f�κk��:q�K�v�E=|��߀������a��c!���ዻ�]`������ߖ������  �  :�=�;=N�=�=h1=	�=]~=y$=^� =p =� =Vv�<*��<��<�V�<:��<���<6�<��<���<��<K[�<���<���<�/�<[t�<���<���<�;�<6|�<o��<���<�6�<�r�<���<���<0 �<xW�<J��<d��<���<�#�<�Q�<�|�<q��<��<r��<��<2(�<I@�<�T�<2e�<�q�<Nz�<�~�<T~�<�y�<�o�<�`�<�L�<�2�<t�<���<���<���<=O�<��<G��<Up�<��<���<M�<���<�e�<���<va�<,��<YB�<*��<�	�<Ld�<�<��<AQ�<7��<�Ӳ<��<kB�<�r�<o��<2Ʃ<&�<�
�<�'�<uB�<OZ�<�o�<X��<ꔚ<Ф�<*��<��<s˒<�Ր<Cގ<��<��<���<��<U��<��<���<�}<?�y<��u<��q<��m<(�i<��e<��a<D�]<��Y<��U<��Q<��M<X�I<�F<�B<G><!&:<�36<C2<�T.<Ii*<ۀ&<�"<�<f�<�<�4<�g<o�<G�<�'<u <���;(J�;��;~��;u��;���;��;$��;l!�;=i�;(ȳ;M?�;�Ϧ;�z�;,A�;$�;V$�;B�;�}�;"�y;a�n;��c;I0Y;D�N;��D; �:;#1;�';�=;�(;UH;�;�<�:���:No�:���:/�:�:��:bt�:BOv:�:Z:��>:ji#:s�:�T�9��9��h9��9���7'��M�)���������a���Y��#���:���Q�� i�q��Xn���Ζ��"��Am��ӱ����ú�(Ϻk_ں���9���������	�����7�V���@�(�$��9*�M�/��$5���:��@��xE���J�$]P�^�U�	J[�{�`�ZAf�!�k��Aq���v��F|��䀻.���/g���'��W狻�����e���$���㖻����  �  ԓ=�;=$�=q�=u1=1�=�~=�$=�� =�p =S =�w�<���<��<2X�<٢�<6��<u7�<]��<���<��<\�<���<��<�/�<-t�<���<���<;�<G{�<>��<F��<95�<<q�<-��<���<��<�U�<��<��<���<�"�<�P�<n|�<"��<��<���<�<�(�<&A�<�U�<cf�<#s�<�{�<��<��<{�<Wq�<Pb�<�M�<�3�<��<���<[��<���<`O�<x�<���<�o�< �<���<�K�<���<d�<U��<�_�<���<�@�<���<%�<�b�<���<��<LP�<|��<mӲ<I�<bB�<�r�<鞫<�Ʃ<�<��<1)�<�C�<�[�<oq�<ᄜ<���<X��<���<S��<�̒<�֐<ߎ<e�<S�<
�<��<��<���<(��<9�}<
�y<&�u<��q<��m<�i<��e<��a<!�]<��Y< �U<R�Q<��M<��I<�F<1B<><P&:<M46<ZD2<uV.<fk*<.�&<��"<ʽ<��<
<�7<Lk<��<1�<`*<ow <��;�M�;��;���;��;a��;��;��;g�;�e�;�ó;K:�; ʦ;�t�;_;�;*�;��;5<�;�x�;A�y;��n;��c;�*Y;a�N;��D;y�:;�1;��';�C;,0;BQ;��;�R�:���:҈�:J��:�+�:���:|�:b��:�vv:^Z:5�>:A�#:6�:�a�9�9-�h9�{9��7$��6B*��P�����GH���6>#��:�R��0i�C��􁋺�ݖ�K0��mw��f���\�ú�'Ϻ�[ں���b���������	����,�p��24�M�$�E-*�+�/�	5���:�^�?�`rE�C�J�_ZP�a�U��J[��`�Ef�O�k��Hq���v�Q|��ꀻZ���8m���-��f틻����^k���)���薻�����  �  o�=O;=��=d�=�1=[�=�~=G%=Z� =>q =� =0y�<6��<�<�Y�<Z��<���<�8�<���<���<��<�\�<��<a��<�/�<
t�<@��<C��<D:�<6z�<��<���<�3�<�o�<���<k��<�<�T�<��<׾�<s��<�!�<+P�<�{�<��<���<���<\�<�)�<B�<�V�<�g�<{t�<.}�<���<i��<�|�<�r�<�c�<MO�<�4�<p�<���<���<P��<�O�<`�<���<Qo�<T�<ų�<�J�<?��<�b�<���<&^�<���<?�<ॾ<��<ga�<T��<��<VO�<���<�Ҳ<�<RB�< s�<E��<�ǩ<��<��<s*�<-E�<<]�<�r�<m��<��<ݧ�<��<�<�͒<�א<�ߎ<��<��<7�<��<���<���<b��<<�}<��y<��u<+�q<��m<��i<��e<D�a<�]<�Y<]�U<��Q<��M<�I<�F<�B<�><�&:<�46<`E2<X.<Em*<��&<;�"<��<��<><;<on<��<0�<%-<�y <��;�P�;��;���;���;6��;���;���;n�;�a�;n��;W5�;�Ħ;o�;E5�;@�;y�;�6�;Cs�;ěy;6�n;ۻc;�%Y;��N;P�D;��:;01;ʎ';I;W7;Y;�;�h�:��:L��:��:�D�:�:6�:���:��v:b}Z:��>:`�#:9�:�s�9��9>�h9�>9 �7@�����*�����sZ��'��"���p#���:�>R�b]i��*������N>�����������ú�'Ϻ�Vں�庇�����Y{�#
	�d����m���'��$�!*�Q�/�a5��:���?��kE���J��WP��U�]K[�-�`��If���k��Pq���v�@[|�"���A����s��4���󋻫����p���.��햻߫���  �  �=;=��=O�=�1=��=/=�%=�� =�q =� =z�<���<{�<O[�<å�<(��<%:�<҃�<��<��<x]�<v��<���<�/�<�s�<ն�<���<�9�<5y�<��<���<x2�<En�<��<���<��<$S�<%��<���<d��<!�<�O�<b{�<���<���<��<��<*�<�B�<�W�<�h�<�u�<�~�<��<��<~�<.t�</e�<zP�<6�<b�<S��<���<���<�O�<9�<b��<�n�<��<��<�I�<��<(a�<`��<�\�<=��<j=�<U��</�<�_�<(��<��<�N�<	��<eҲ<��<=B�<4s�<���<ȩ<��<��<�+�<aF�<�^�<Lt�<���<y��<B��<a��<�Ô<�Β<vؐ<���<~�<�<]�<f�<{��<p��<���<u�}<��y<0�u<s�q<�m<��i<��e<=�a<A�]<V�Y<��U<��Q<��M<��I<kF<�B<f><�&:<�56<WF2<�Y.<	o*<��&<��"<x�<��<6<@><`q<��<��<�/<| <���;�S�;��;��;.��;���;���;���;�;F^�;v��;�0�;ÿ�;�i�;�/�;��;��;�1�;n�;W�y;9�n;��c;!Y;��N;��D;޼:;�1;=�';�M;�=;�`;|�;R|�:���:ŷ�:3��:&]�:s,�:�L�:���:��v:+�Z:Y�>:�#:S�:ˀ�9��9��h9T�9ç�7����U+�冹���
��i���#��;�BlR�
�i��?����������I������Ÿ���ú�'Ϻ\Rں}庆�����Cs�	����j�2��E�x�$��*���/�5�{:���?��eE���J��TP��U��L[���`�NNf�s�k��Wq��v��d|�����ŷ���y��:������4���Qv���3��T񖻐����  �  =�:=��=H�=�1=��=q=�%=0� =?r = =�{�<���<��<~\�<��<T��<>;�<ք�<���<S�<^�<��<���<�/�<�s�<���<7��<�8�<jx�<��<���<L1�<m�<٧�<���<b�<�Q�<��<���<���<U �<�N�<{�<v��<���<��<�<�*�<kC�<�X�<�i�<�v�<��<)��<��<E�<gu�<Kf�<�Q�<�6�<;�<���<��<��<�O�<*�< ��<Sn�<�<��<�H�<���<�_�<��<J[�<���<<�<	��<��<�^�<��<��<�M�<s��<Ҳ<��<1B�<Js�<
��<�ȩ<]�<��<�,�<pG�<�_�<�u�<#��<���<}��<���<�Ĕ<�ϒ<Gِ<Q�<�<\�<p�<a�<@��<	��<��<��}<��y<�u<*�q<��m<_�i<�e<��a<��]<��Y<��U<��Q<P�M<@�I<~F<EB<E><�&:<66<^G2<�Z.<�p*<��&<��"<��<�<�<�@<�s<�<.�<�1<�} <���;sV�;�;��;���;���;���;4��;_�;a[�;ⷳ;�,�;U��;e�;�*�;��;9�;�,�;�i�;��y;�n;�c;wY;4�N;r�D;�:;�1;y�';BR;2C;
h;�;���:���:���: ��:�p�:�@�:�^�:ŉ:0�v:�Z:?:��#:��:���9��9|th9Q�9Q�7�x����+�6%�������F�����#�SG;��R��i��P��Ƶ�����{U��͓��ʸ���úQ'ϺPں�u�ٙ�ú��!l����σ�%�B����o�$�*���/���4��s:�C�?��`E���J�vRP���U��L[���`��Qf���k�	^q��v�$m|��������y~��)?������(����z��8����������  �  ��=�:=��==�=�1=��=�=%&=}� =�r =� =}|�<���<��<p]�<��<<��<<�<���<|��<��<p^�<B��<��<�/�<�s�<F��<���<Q8�<�w�<C��<���<d0�<l�<ۦ�<���<e�<�P�<9��<߻�<���<��<zN�<�z�<.��<���<?��<X�<�*�<�C�<Y�<Uj�<�w�<���< ��<��<;��<av�<&g�<bR�<�7�<��<t��<V��<>��<�O�<,�<���<n�<��<���<	H�<��<_�<��<;Z�<���<;�<���<��<�]�<:��<��<M�<��<�Ѳ<Q�<:B�<fs�<H��<�ȩ<��<"�<<-�<MH�<�`�<�v�<��<���<m��<_��<�Ŕ<|В<�ِ<��<b�<��<��<T�<���<���<���<��}<s�y<l�u<r�q<��m<e�i<��e<��a<��]<6�Y<�U<d�Q<1�M<4�I<�F<�B<><�&:<w66<H2<�[.<�q*<Պ&<l�"<��<��<�<�B<v<�<�<c3<8 <y��;KX�;��;���;/��;D��;���;��;x�;WY�;���;�)�;跦;Ka�;%'�;�	�;v
�;>)�;�f�;F�y;�zn;2�c;Y;~�N;p�D;d�:;.1;�';GU;bG;�l;��;��:��:���:�:��:�P�:m�:{Ӊ:��v:E�Z:�?:��#:��:��9��9�Sh9=�9@��7����,�XZ���)��-�蹼2���#�Tg;�вR���i��]��������]��ș��'θ�"�ú�%ϺzMں
q庐��ձ��tg����|���@��2
�s�$��*��~/���4��n:�`�?�A]E���J��PP���U�KM[���`��Sf���k�Obq���v��s|�{�������b���@C�����!���f~��V;������ִ���  �  _�=�:=}�=4�=�1=��=�=P&=�� =�r =� =�|�<F��<J�<^�<���<���<�<�<��<���<J�<�^�<h��< ��<�/�<�s�<��<���<8�<cw�<ʵ�<F��<�/�<k�<D��<��<��<hP�<���<\��<e��<g�<5N�<�z�<��<���<G��<~�</+�<KD�<�Y�<�j�<x�<��<���<���<Ҁ�<�v�<�g�<�R�<"8�<7�<���<���<`��<�O�<�<���<�m�<9�<��<�G�<���<�^�<y��<�Y�<5��<h:�<`��<S�<g]�<���<x�<�L�<���<|Ѳ<2�<)B�<ss�<h��<8ɩ<B�<��<�-�<�H�<&a�<
w�<���<E��<���<ܹ�<;Ɣ<�В<Sڐ<%�<��<��<��<E�<���<���<X��<�}<|�y<g�u<W�q<q�m<1�i<��e<��a<��]<�Y<��U<i�Q<J�M<��I<bF<dB<�><�&:<�66<ZH2<B\.<�r*<Ջ&<h�"<��<�<<D<3w<'�<�<m4<B� <,��;�Y�;G�;��;;��;��;t��;2��;g�;�W�;5��;�'�;ϵ�;4_�;�$�;��;>�;.'�;�d�;`�y;*wn;$�c;Y;��N;��D;<�:;�1;͘';8W;�J;�p;��;���:�:1��:k�:(��:Y�:Mu�:Kۉ:�	w:��Z:� ?:��#:��:��9�9aHh9D�9��7Xa���M,�Zz���L�����D�d�#��y;���R�]�i�f��/ʋ�]��>c��띭��и���ú|&Ϻ6Lں�n��𺎫���c� ���x���������$�S *��z/��4��j:��?�~ZE�^�J��OP�~�U��M[���`��Uf���k��eq���v��w|������������E�����MÎ�����h=�����������  �  R�=v:=y�=3�=�1=��=�=W&=�� =�r =� =7}�<���<w�<S^�<���<��<�<�<C��<��<K�<�^�<���<4��<�/�<�s�<��<~��<�7�<>w�<���<��<�/�<Ek�<��<���<��<1P�<u��<E��<G��<L�<N�<gz�<��<���<O��<��<A+�<SD�<�Y�<�j�<;x�<L��<��<܅�<��<#w�<�g�<S�<H8�<H�<���<���<��<�O�<�<���<�m�< �<���<aG�<y��<O^�<<��<_Y�<���<":�<!��<�<2]�<���<O�<�L�<���<kѲ<6�<B�<�s�<���<Jɩ<B�<��<�-�<�H�<la�<<w�<�<t��<7��<��<mƔ<'ђ<Xڐ<1�<��<��<��<D�<���<^��<?��<��}<F�y<*�u<��q<��m<��i<P�e<�a<#�]<��Y<��U<6�Q<�M<l�I<F<TB<�><�&:<�66<�H2<]\.<�r*<$�&<ƨ"<
�<��<a<D<�w<��<��<�4<�� <;��;�Y�;��;���;3��;@��;S��;���;�;W�;겳;�&�;촦;W^�;�#�;��;P�;Z&�;�c�;��y;Mvn;^�c;tY;ؾN;/�D;I�:;�1;ę';�W;�J;�p;��;���:��:W��:��:׍�:�\�:�y�:�݉:�w:��Z:k!?:5�#:��:���9#�9XLh9�9�)�7(z���],����Z��p�蹀L�b$�1�;�)�R���i� i���ˋ�����d�������Ѹ��ú'Ϻ*Kں�l庯��l����b����Fw����\��9�{�$�:�)��x/�u�4��i:���?�"ZE���J��NP�~�U��M[���`�Wf���k��fq���v��x|�� ���Ã�����F�����7Ď������=��=�������  �  _�=�:=}�=4�=�1=��=�=P&=�� =�r =� =�|�<F��<J�<^�<���<���<�<�<��<���<J�<�^�<h��< ��<�/�<�s�<��<���<8�<cw�<ʵ�<F��<�/�<k�<D��<��<��<hP�<���<\��<e��<g�<5N�<�z�<��<���<G��<~�</+�<LD�<�Y�<�j�<x�<��<���<���<Ҁ�<�v�<�g�<�R�<"8�<7�<���<���<`��<�O�<�<���<�m�<9�<��<�G�<���<�^�<y��<�Y�<5��<h:�<`��<S�<g]�<���<x�<�L�<���<|Ѳ<2�<)B�<ss�<h��<8ɩ<B�<��<�-�<�H�<&a�<
w�<���<E��<���<ܹ�<;Ɣ<�В<Sڐ<%�<��<��<��<E�<���<���<X��<�}<|�y<g�u<W�q<q�m<1�i<��e<��a<��]<�Y<��U<i�Q<J�M<��I<bF<dB<�><�&:<�66<ZH2<B\.<�r*<Ջ&<h�"<��<�<<D<3w<'�<�<m4<B� <,��;�Y�;F�;��;;��;��;t��;2��;g�;�W�;5��;�'�;ϵ�;4_�;�$�;��;>�;.'�;�d�;_�y;*wn;$�c;Y;��N;��D;<�:;�1;͘';8W;�J;�p;��;���:�:1��:k�:(��:Y�:Mu�:Kۉ:�	w:��Z:� ?:��#:��:��9�9aHh9D�9��7Xa���M,�Zz���L�����D�d�#��y;���R�]�i�f��/ʋ�]��>c��띭��и���ú|&Ϻ6Lں�n��𺎫���c� ���x���������$�S *��z/��4��j:��?�~ZE�^�J��OP�~�U��M[���`��Uf���k��eq���v��w|������������E�����MÎ�����h=�����������  �  ��=�:=��==�=�1=��=�=%&=}� =�r =� =}|�<���<��<p]�<��<<��<<�<���<|��<��<p^�<B��<��<�/�<�s�<F��<���<Q8�<�w�<C��<���<d0�<l�<ۦ�<���<e�<�P�<9��<߻�<���<��<zN�<�z�<.��<���<?��<X�<�*�<�C�<Y�<Uj�<�w�<���< ��<��<;��<av�<&g�<bR�<�7�<��<t��<V��<>��<�O�<,�<���<n�<��<���<	H�<��<_�<��<;Z�<���<;�<���<��<�]�<:��<��<M�<��<�Ѳ<Q�<:B�<fs�<H��<�ȩ<��<"�<<-�<MH�<�`�<�v�<��<���<m��<_��<�Ŕ<|В<�ِ<��<b�<��<��<T�<���<���<���<��}<s�y<l�u<r�q<��m<e�i<��e<��a<��]<6�Y<�U<d�Q<1�M<4�I<�F<�B<><�&:<w66<H2<�[.<�q*<Պ&<l�"<��<��<�<�B<v<�<�<c3<8 <x��;KX�;��;���;/��;D��;���;��;x�;WY�;���;�)�;跦;Ka�;$'�;�	�;v
�;>)�;�f�;F�y;�zn;1�c;Y;~�N;p�D;d�:;.1;�';GU;bG;�l;��;��:��:���:�:��:�P�:m�:{Ӊ:��v:E�Z:�?:��#:��:��9��9�Sh9=�9@��7����,�XZ���)��-�蹼2���#�Tg;�вR���i��]��������]��ș��'θ�"�ú�%ϺzMں
q庐��ձ��tg����|���@��2
�s�$��*��~/���4��n:�`�?�A]E���J��PP���U�KM[���`��Sf���k�Obq���v��s|�{�������b���@C�����!���f~��V;������ִ���  �  =�:=��=H�=�1=��=q=�%=0� =?r = =�{�<���<��<~\�<��<T��<>;�<ք�<���<S�<^�<��<���<�/�<�s�<���<7��<�8�<jx�<��<���<L1�<m�<٧�<���<b�<�Q�<��<���<���<U �<�N�<{�<v��<���<��<�<�*�<kC�<�X�<�i�<�v�<��<)��<��<E�<gu�<Kf�<�Q�<�6�<;�<���<��<��<�O�<*�< ��<Sn�<�<��<�H�<���<�_�<��<J[�<���<<�<	��<��<�^�<��<��<�M�<s��<Ҳ<��<1B�<Js�<
��<�ȩ<]�<��<�,�<pG�<�_�<�u�<#��<���<}��<���<�Ĕ<�ϒ<Gِ<Q�<�<\�<p�<a�<@��<	��<��<��}<��y<�u<*�q<��m<_�i<�e<��a<��]<��Y<��U<��Q<P�M<@�I<~F<EB<E><�&:<66<^G2<�Z.<�p*<��&<��"<��<�<�<�@<�s<�<.�<�1<�} <���;sV�;�;��;���;���;���;4��;^�;a[�;ⷳ;�,�;U��;e�;�*�;��;9�;�,�;�i�;��y;�n;�c;wY;4�N;r�D;�:;�1;y�';BR;2C;
h;�;���:���:���: ��:�p�:�@�:�^�:ŉ:0�v:�Z:?:��#:��:���9��9|th9Q�9Q�7�x����+�6%�������F�����#�SG;��R��i��P��Ƶ�����{U��͓��ʸ���úQ'ϺPں�u�ٙ�ú��!l����σ�%�B����o�$�*���/���4��s:�C�?��`E���J�vRP���U��L[���`��Qf���k�	^q��v�$m|��������y~��)?������(����z��8����������  �  �=;=��=O�=�1=��=/=�%=�� =�q =� =z�<���<{�<O[�<å�<(��<%:�<҃�<��<��<x]�<v��<���<�/�<�s�<ն�<���<�9�<5y�<��<���<x2�<En�<��<���<��<$S�<%��<���<d��<!�<�O�<b{�<���<���<��<��<*�<�B�<�W�<�h�<�u�<�~�<��<��<~�<.t�</e�<zP�<6�<b�<S��<���<���<�O�<9�<b��<�n�<��<��<�I�<��<(a�<`��<�\�<=��<j=�<U��</�<�_�<(��<��<�N�<	��<eҲ<��<=B�<4s�<���<ȩ<��<��<�+�<aF�<�^�<Lt�<���<y��<B��<a��<�Ô<�Β<vؐ<���<~�<�<]�<f�<{��<p��<���<u�}<��y<0�u<s�q<�m<��i<��e<=�a<A�]<V�Y<��U<��Q<��M<��I<kF<�B<g><�&:<�56<WF2<�Y.<	o*<��&<��"<x�<��<6<@><`q<��<��<�/<| <���;�S�;��;��;.��;���;���;���;�;F^�;v��;�0�;¿�;�i�;�/�;��;��;�1�;n�;V�y;9�n;��c;!Y;��N;��D;޼:;�1;=�';�M;�=;�`;|�;R|�:���:ŷ�:3��:&]�:s,�:�L�:���:��v:+�Z:Y�>:�#:S�:ˀ�9��9��h9T�9ç�7����U+�冹���
��i���#��;�BlR�
�i��?����������I������Ÿ���ú�'Ϻ\Rں}庆�����Cs�	����j�2��E�x�$��*���/�5�{:���?��eE���J��TP��U��L[���`�NNf�s�k��Wq��v��d|�����ŷ���y��:������4���Qv���3��T񖻐����  �  o�=O;=��=d�=�1=[�=�~=G%=Z� =>q =� =0y�<6��<�<�Y�<Z��<���<�8�<���<���<��<�\�<��<a��<�/�<
t�<@��<C��<D:�<6z�<��<���<�3�<�o�<���<k��<�<�T�<��<׾�<s��<�!�<+P�<�{�<��<���<���<\�<�)�<B�<�V�<�g�<{t�<.}�<���<i��<�|�<�r�<�c�<MO�<�4�<p�<���<���<P��<�O�<`�<���<Qo�<T�<ų�<�J�<?��<�b�<���<&^�<���<?�<ॾ<��<ga�<T��<��<VO�<���<�Ҳ<�<RB�< s�<E��<�ǩ<��<��<s*�<-E�<<]�<�r�<m��<��<ݧ�<��<�<�͒<�א<�ߎ<��<��<7�<��<���<���<b��<<�}<��y<��u<+�q<��m<��i<��e<D�a<�]<�Y<]�U<��Q<��M<�I<�F<�B<�><�&:<�46<aE2<X.<Em*<��&<;�"<��<��<><;<on<��<0�<%-<�y <��;�P�;��;���;���;5��;���;���;n�;�a�;m��;W5�;�Ħ;o�;D5�;@�;y�;�6�;Cs�;ěy;6�n;ۻc;�%Y;��N;O�D;��:;01;ʎ';I;W7;Y;�;�h�:��:L��:��:�D�:�:6�:���:��v:b}Z:��>:`�#:9�:�s�9��9>�h9�>9 �7@�����*�����sZ��'��"���p#���:�>R�b]i��*������N>�����������ú�'Ϻ�Vں�庇�����Y{�#
	�d����m���'��$�!*�Q�/�a5��:���?��kE���J��WP��U�]K[�-�`��If���k��Pq���v�@[|�"���A����s��4���󋻫����p���.��햻߫���  �  ԓ=�;=$�=q�=u1=1�=�~=�$=�� =�p =S =�w�<���<��<2X�<٢�<6��<u7�<]��<���<��<\�<���<��<�/�<-t�<���<���<;�<G{�<>��<F��<95�<<q�<-��<���<��<�U�<��<��<���<�"�<�P�<n|�<"��<��<���<�<�(�<&A�<�U�<cf�<#s�<�{�<��<��<{�<Wq�<Pb�<�M�<�3�<��<���<[��<���<`O�<x�<���<�o�< �<���<�K�<���<d�<U��<�_�<���<�@�<���<%�<�b�<���<��<LP�<|��<mӲ<I�<bB�<�r�<鞫<�Ʃ<�<��<1)�<�C�<�[�<oq�<ᄜ<���<X��<���<S��<�̒<�֐<ߎ<e�<R�<
�<��<��<���<'��<9�}<	�y<&�u<��q<��m<�i<��e<��a<!�]<��Y< �U<R�Q<��M<��I<�F<1B<><P&:<M46<ZD2<uV.<gk*<.�&<��"<ʽ<��<
<�7<Lk<��<1�<`*<ow <��;�M�;��;���;��;a��;��;��;g�;�e�;�ó;J:�; ʦ;�t�;_;�;*�;��;5<�;�x�;@�y;��n;��c;�*Y;a�N;��D;y�:;�1;��';�C;,0;BQ;��;�R�:���:҈�:J��:�+�:���:|�:b��:�vv:^Z:5�>:A�#:6�:�a�9�9-�h9�{9��7$��6B*��P�����GH���6>#��:�R��0i�C��􁋺�ݖ�K0��mw��f���\�ú�'Ϻ�[ں���b���������	����,�p��24�M�$�E-*�+�/�	5���:�^�?�`rE�C�J�_ZP�a�U��J[��`�Ef�O�k��Hq���v�Q|��ꀻZ���8m���-��f틻����^k���)���薻�����  �  :�=�;=N�=�=h1=	�=]~=y$=^� =p =� =Vv�<*��<��<�V�<:��<���<6�<��<���<��<K[�<���<���<�/�<[t�<���<���<�;�<6|�<o��<���<�6�<�r�<���<���<0 �<xW�<J��<d��<���<�#�<�Q�<�|�<q��<��<r��<��<2(�<I@�<�T�<2e�<�q�<Nz�<�~�<T~�<�y�<�o�<�`�<�L�<�2�<t�<���<���<���<=O�<��<G��<Up�<��<���<M�<���<�e�<���<va�<,��<YB�<*��<�	�<Ld�<�<��<AQ�<7��<�Ӳ<��<kB�<�r�<o��<2Ʃ<&�<�
�<�'�<uB�<OZ�<�o�<X��<ꔚ<Ф�<*��<��<s˒<�Ր<Cގ<��<��<���<��<U��<��<���<�}<?�y<��u<��q<��m<(�i<��e<��a<D�]<��Y<��U<��Q<��M<X�I<�F<�B<G><!&:<�36<C2<�T.<Ii*<܀&<�"<�<f�<�<�4<�g<o�<G�<�'<u <���;(J�;��;~��;u��;���;��;#��;l!�;=i�;(ȳ;M?�;�Ϧ;�z�;+A�;$�;V$�;B�;�}�;"�y;a�n;��c;I0Y;D�N;��D; �:;#1;�';�=;�(;UH;�;�<�:���:No�:���:/�:�:��:bt�:BOv:�:Z:��>:ji#:s�:�T�9��9��h9��9���7'��M�)���������a���Y��#���:���Q�� i�q��Xn���Ζ��"��Am��ӱ����ú�(Ϻk_ں���9���������	�����7�V���@�(�$��9*�M�/��$5���:��@��xE���J�$]P�^�U�	J[�{�`�ZAf�!�k��Aq���v��F|��䀻.���/g���'��W狻�����e���$���㖻����  �  ��=<={�=��=Q1=��=~=&$=�� =�o = =�t�<ƿ�<l
�<"U�<���<_��<�4�<�~�<���<��<�Z�<q��<���<w/�<t�<W��<��<�<�<!}�<���<���<8�<%t�<+��<��<�!�<�X�<���<���<���<�$�<?R�<F}�<���<���<F��<#�<�'�<�?�<�S�<!d�<�p�<�x�<}�<�|�<x�<Sn�<�_�<TK�<|1�<q�<(��<(��<(��<O�<��<���<�p�<��<���<N�<.��<�f�<w��<�b�<���<�C�<���<:�<�e�<1��<��<R�<ו�<XԲ<��<\B�<tr�<���<�ũ<^�<�	�<�&�<"A�<�X�<_n�<ځ�<p��<h��<α�<���<_ʒ<�Ԑ<�ݎ<!�<��<���<��<���<x��<���<��}<]�y<�u<i�q<��m<�i< �e<��a<�]<��Y<�U<��Q<��M<� J<�F<�B<{><�%:<�26<�A2<�S.<ag*<�~&<\�"<,�<��<�<s1<�d<��<l�<.%<�r <Ҏ�;aG�;Z�;	��;���;���;F��;���;
$�;�l�;a̳;�C�;�Ԧ;��;�F�;*�;�)�;vG�;���;��y;�n;��c;�4Y;A�N;i�D;��:;k1;�';�8;�";�?;V�;�'�:Ԑ�:�W�:P|�:���:`̦:�:�^�:�,v:�Z:��>:eV#:~�:I�9��9� i9��9��7�V��MD)�̵��l\��\��o-���"��\:�4�Q���h�k��\��ڿ������d������J�ú�*Ϻcں�������� ���'	����xB�H���L�
�$��D*�(�/��.5�G�:��@�U~E�$�J�V`P���U��I[���`��=f�κk��:q�K�v�E=|��߀������a��c!���ዻ�]`������ߖ������  �  ݔ=]<=��=��=I1=��=�}=�#=�� =o =� =�s�<���<4	�<�S�<���<#��<�3�<�}�<���</�<Z�<	��<K��<q/�<�t�<���<���<N=�<�}�<|��<���</9�<cu�<k��<F��<�"�<Z�<���<���<}��<M%�<�R�<�}�<إ�<��< ��<��<'�<�>�<�R�<(c�<mo�<�w�<�{�<�{�<�v�<%m�<l^�<BJ�<�0�<��<t��<���<ۉ�<�N�<��<���<Qq�<+�<b��<O�<8��<�g�<���<Ed�<��<AE�<���<q�<�f�<2��<�	�<�R�<s��<�Բ< �<iB�<Gr�<���<ũ<��<��<�%�<@�<�W�<1m�<���<6��</��<���<���<fɒ<�Ӑ<�܎<��<A�<���<��<���<���<$��<G�}<%�y<&�u<��q<�m<��i<��e<�a<��]<��Y<5�U<��Q<F�M<�J<	F<B<�><�%:<z26<A2<R.<�e*<�|&<4�"<ε<��<0<�.<Rb<��<�<�"<�p <}��;jD�;q�;���;!��;���;*��;���;>&�;�o�;�ϳ;�G�;٦;���;|K�;�.�;a.�;�K�;���;E�y;��n;1�c;�8Y;��N;:�D;n�:;�1;�';f4;�;�8;M�;��:_}�:MD�:Th�:��: ��:�ݗ:JM�:�v:��Y:�i>:0D#:U�:=�9��9�i9�92 �7]���v�(�x��[���C湵��"��4:�G�Q���h�(��OM��L���&��2\�������ú�*Ϻ�fں��9����H���/	����AL�����V���$��N*�|�/�075���:�@�&�E���J��bP���U�rI[�{�`��9f�>�k�v4q�-�v�!5|�Zۀ�⛃�~\������܋�%����[�����ܖ�q����  �  �=�<=��=��=<1=��=�}=�#=;� =�n =  =�r�<���<8�<�R�<���<)��<�2�<}�<��<��<�Y�<á�< ��<f/�<�t�<ٸ�<���<�=�<�~�<��<���<:�<Uv�<j��<;��<�#�<�Z�<|��<A��<��<�%�<+S�<~�<���<��<���<��<�&�<L>�<HR�<Zb�<�n�<�v�<�z�<�z�<�u�<)l�<~]�<yI�<�/�<�<���<A��<���<�N�<��<���<�q�<��<���<�O�<���<�h�<���<Te�<��<OF�<��<_�<�g�<껹<|
�<cS�<ݖ�<ղ<-�<sB�<
r�<p��<�ĩ<*�<<�<%�<A?�<�V�<9l�<��<:��</��<���<ڼ�<�Ȓ<)Ӑ<M܎<K�<��<p��<��<���<C��<���<q�}<W�y<��u<j�q<��m<��i<p�e<&�a<p�]<��Y<��U<��Q<��M<�J<�	F<�B<�><�%:<�16<o@2<Q.<�d*<E{&<��"<��<��<(�<�,<J`<�<H�<4!<Zo <"��;9B�;�;b��;���;0��;���;���;�'�;�q�;ҳ;�J�;Uܦ;E��;EO�;,2�;42�;8O�;��;��y;��n;O�c;�;Y;z�N;)�D;ּ:;1;�~'; 1;E;K4;��;��:Dn�:'4�:X�:xյ:㨦:7Η:Q@�:��u:��Y:�X>:�6#:�z:U-�9��9:!i9�79��7����(��J�� ߵ�c���
� �"�,:�vhQ��h����B������5���V��p�����ú.+Ϻ�kں�庽����\���6	���T�����^���$��V*���/��=5��:��@�Z�E���J��dP���U��H[��`�F7f���k��/q�i�v��.|��׀�6���yX������؋�o���eX������ٖ�����  �  ?�=�<=��=��=21=��=�}=e#=� =}n =� =gr�<���<��<AR�<���<���<42�<�|�<���<<�<CY�<���<���<W/�<�t�<���<��<#>�<�~�<���<,��<�:�<�v�<���<���<^$�<u[�<���<���<���<?&�<sS�<(~�<��<��<���<d�<u&�<�=�<�Q�<�a�<n�<Mv�<Vz�<z�<:u�<�k�<�\�<�H�<=/�<��<���<���<z��<�N�<��<��<�q�<��<f��<1P�<���<xi�</��<�e�<���<�F�<���<��</h�<r��<�
�<�S�<��<9ղ<>�<qB�<�q�<@��<cĩ<��<��<�$�<�>�<IV�<�k�<�<���<���</��<U��<'Ȓ<�Ґ<܎<�<��<[��<��<��<i��<���<;�}<T�y<��u<d�q<�m<��i<��e<?�a<��]<��Y<��U<��Q<V�M<�J<
F<�B<�><`%:<�16<�?2<�P.<�c*<Nz&<~�"<�<��<��<{+<_<˘<�<! <Pn <W��;A�; 
�;���;Z��;&��;3��;n��;6)�;Zs�;�ӳ;�L�;'ަ;=��;hQ�;�4�;?4�;?Q�;֋�;��y;��n;D�c;�=Y;��N;��D;d�:;)1;Q}';�.;c;g0;�~;- �:Se�:+�:�N�:7̵:ş�:aŗ:�7�:�u::�Y:�L>:�-#:Ct:D'�9��9,(i9iK9���7^���4O(�+��쿵�����
���"��:��WQ�>�h�X���:��¡��E���S�����G�ú�+Ϻ�lں��������K���:	�v��^X�q���c���$�[*��/��A5��:�2@���E���J��eP�U�U��H[�0�`�6f�|�k��,q�x�v��*|��Հ����PV��<��a֋�Q���rV������ז�p����  �  }�=[9=�=��=�,=��=Ux=�=&� =Yh =U =�d�<:��<���<OA�<���<���<��<oe�<���<R��<}<�<���<2��<��<7P�<���<���<��<�R�<���<��<j�<�B�<W{�<ز�<���<`�<P�<��<��<���<�<�.�<�S�<�u�<��<���<���<���<���<��<q�<�
�<�<��<�<���<	��<��<���<]��<�d�<6�<� �<;��<Ӏ�<[6�<~��<m��<+�<l��<�T�<���<b�<t��<4T�<�ÿ<�,�<r��<O�<�C�<���<�<�'�<Si�<��<�ݮ<�<�@�<l�<���<<�أ<-��<��<,�<gC�<�X�<@l�<=~�<���<���<B��<���<�<s̊<Ո<�܆<�<��<H�<h�}<E�y<(�u<��q<��m<��i<�f<_
b<^<JZ<� V<"*R<z4N<C@J<MF<~[B<Kk><�|:<,�6<��2<�.<��*<v�&<S#<�?<Bj<�<�<�	<�J<�<�<�4<�!�;���;k��;դ�;���;��;���;X��;-�;n��;��;^t�;�;!Ǣ;���;���;ه�;��;6�;^�~;Svs;��h;�];j�S;hI;An?;�5;,;S�";��;�;c�;ܩ�:���:��:�v�:X½:y`�:�O�:���: �:��g:f�K:��/:�:���9�۾9��9&�-9�[�8E������e�=B���չ��p��#�2�I0J��a��y����e����'��ܝ��.
���m���̺�&غ�{㺓��8����RH����"x�N
�Ζ��$��)��$/���4�N:�l�?��E�ЈJ��P�|U��Z��u`�b�e��wk���p�t�v��|��ƀ�׉���M�����ԋ�*����\��� ���喻����  �  i�=U9=�=z�=�,=��=hx=�=8� =dh =d =�d�<[��<���<cA�<�<���<��<�e�<̭�<s��<�<�<ڂ�<K��<��<#P�<���<���<��<�R�<p��<���<T�<iB�<:{�<���<���<?�<P�<��<��<���<�<�.�<�S�<�u�<��<���<���<���<���<-��<��<�
�<.�<��<<�<���<��<;��<ï�<s��<�d�<"6�<� �<F��<Ԁ�<F6�<|��<Z��<�*�<S��<�T�<���<�a�<F��<T�<cÿ<k,�<X��<K�<iC�<䔷<��<�'�<Oi�< ��<�ݮ<��<�@�<.l�<���<���<
٣<L��<��<J,�<C�<�X�<bl�<R~�<���<ʝ�<h��<���<�<�̊< Ո<�܆<�<��<"�<<�}<�y<�u<t�q<��m<��i<.f<
b<�^<*Z<� V<�)R<O4N<�?J<�LF<U[B<-k><�|:<b�6<�2<=�.<8�*<��&<�#<�?<�j<<�<H�<'
<K<V�<5�<#5<"�;��;(��;D��;���;���;��;-��;�,�;;��;"�;Vt�;��;aƢ;=��;��;H��;���;@�;��~;�us;��h;X�];b�S;\gI;*n?;2�5;�,;�";��;�;B�;]��:���:���:�x�:�Ľ:Kc�:�P�:4��:��:��g:��K:*�/:��:��9�ܾ9���9h�-9�K�8��)����e�A���չ]�������2�m6J�	�a��y���V����)������J
��,o����̺Z%غ7y�p�� ������G�����w������$��)��#/���4�~:�9�?��E���J�P��{U�|�Z��v`���e�yk�m�p�X�v�$|��ƀ�����#N�����KՋ������\�� !��<斻U����  �  M�=I9=��=~�=�,=��=zx==b� =�h =� =e�<Ѯ�<s��<�A�<I��<]��<[�<�e�<��<���<�<�<���<Q��<��< P�<g��<���<��<yR�<��<���<��<�A�<�z�<9��<M��<��<�O�<���<���<t��<��<�.�<�S�<�u�<���<���<��<���<'��<���<	�<b�<��<o	�<��<7��<���<���<��<���<:e�<F6�<� �<G��<���</6�<Z��<(��<�*�<��<T�<B��<^a�<���<�S�<�¿<�+�<؎�<��<�B�<���<��<}'�<-i�<�<ޮ<��<�@�<Kl�<��<J��<m٣<���<[�<�,�<�C�<NY�<�l�<�~�<0��<��<���<뷎<�<�̊<+Ո<�܆<��<m�<��<��}<U�y<:�u<��q<��m<��i<.f<?	b<�^<MZ<�V<)R<�3N<?J<�LF<"[B<;k><�|:<u�6<I�2<��.<��*<I�&<v#<�@<xk<J�<-�<?<�K<J�<�<�5<l#�;���;���;w��; ��;���;���;���;�+�;v��;��;�r�;�;Ģ;���;-�;���;���;��;f�~;Uss;�h; �];��S;�fI;�n?;t�5;�,;r�";��;��;��;���:���:Ό�:U��:�˽:�k�:JW�:���:5�:��g:�K:&�/:7�:`��9��9���9�-9 �8��򷗸��6f�^[��4չ��������2��EJ��a�:y�%������-��𠪺����o����̺%غ�w�W��G�����D����5t�������$�6�)�o /��4��:���?�pE���J�� P��{U��Z�Bw`�h�e��zk��p�2�v�p
|��Ȁ�|����O������֋�󚎻x^���"���疻)����  �  $�=#9=��=y�=�,=��=�x=8=�� =�h =� =�e�<y��<"��<�B�<��<��<��<�f�<���<0��<=�<<��<{��<��<P�<)��<J��<+�<�Q�<���< ��<;�<GA�<z�<���<���<�<O�<��<#��<��<��<v.�<�S�<�u�<��<���<r��<\��<���<��<��<�<P�<-
�<n�<���<0��<:��<���<4��<�e�<�6�<� �<Z��<р�<6�<��<Ҋ�<>*�<~��<�S�<���<�`�<��<�R�<$¿<5+�<$��<4�<nB�<��<7�<&'�<�h�<ץ�<ޮ<��<,A�<�l�<l��<���<�٣<T��<�<u-�<�D�<Z�<�m�<h�<Ï�<���<,��<[��<9Ì<�̊<=Ո<�܆<��<#�<��<��}<]�y<�u<X�q<J�m<t�i<�f<�b<h^<Z<�V<(R<�2N<�>J<'LF<�ZB<#k><�|:<Ԑ6<�2<m�.<��*<Z�&<�#<�A<�l<��<��<�<eM<��<T�<�6<F%�;���;���;J��;F��;���;Լ�;���;o*�;���;��;�p�;��;¢;ؑ�;}|�;��;T��;Y�;�~;�os;Șh;��];��S;2fI;�n?;Q�5;�,;E�";�;��;��;��:���:*��:���:ؽ:�u�:�b�:���:q�:��g:<�K:��/:4�:F��9A߾9}�9�]-9Iԍ8�O�����tf�����A]չ�����9�2��ZJ���a��&y�},��9����3������$���p��a�̺�"غIs����-���?�#���n�r��X��$� �)�./�z�4��:�2�?��	E��J���O�"{U�_�Z��x`���e�}k��q��v��|�ˀ�
����R��m���ً�y����`��%���閻����  �  �=�8=��=o�=�,=��=�x=y=�� =.i =I =�f�<o��<
��<�C�<Ռ�<��<��<Ig�<R��<���<�=�<���<���<��<�O�<���<���<��<XQ�<ގ�<,��<c�<Y@�<!y�<���<���<@�<,N�<O�<z��<{��<0�<2.�<�S�<�u�<8��<=��<���<���<;��<���<h�<��<6�<!�<d�<���< ��<��<m��<Ԏ�<#f�<�6�<)�<���<���<�5�<���<m��<�)�<���<�R�<���<�_�<��<�Q�<&��<3*�<<��<L�<�A�<`��<�ߵ<�&�<�h�<���<�ݮ<��<jA�<m�<�<k��<�ڣ<&��< �<S.�<�E�<�Z�<sn�<S��<���<k��<Ĭ�<㸎<�Ì<͊<XՈ<�܆<��<��<<�<��}<�y<��u<��q<��m<}�i< f<�b<�^<AZ<�V<�&R<�1N<�=J<{KF<nZB<�j><}:<P�6<��2<q�.<��*<��&<;#<�C<�n<��<��<{<nO<c�<��<k8<�'�;���;m��;k��;���;���;a��;���;�(�;V~�;U�;�m�;t	�;���;F��;!y�;]�;	��;�;�y~;�js;ߔh;J�];ĒS;�eI;�n?;ܭ5;!",;��";��;��;�;6��:�:��:%��:��:_��:�q�:��:-#�:�g:�K:�0:��:���9oݾ9)w�9�?-9�|�8P���L�n�f����!�չ��?���2��xJ���a��Ay��7��S���;��ݪ��,��r����̺Gغ�n�ܷ���������9�c���f�f��w���$�o�)��/�3�4��:�}�?��E�9�J���O�^zU���Z��y`�3�e�?�k�~q�H�v�C|��΀������V������݋����od��=(��Q얻~����  �  ��=�8=��=h�=�,=
�=�x=�==� =�i =� =�g�<}��<)��<�D�<���<��<��<*h�<��<o��<>�<��<���<��<�O�<���<��<!�<�P�<��<F��<h�<K?�<x�<���<���<7�<9M�<h~�<ĭ�<���<��<�-�<cS�<�u�<X��<���<Q��<���<���<���<U�<��<R�<0�<o�<���<��<���<8��<���<�f�<s7�<k�<���<���<�5�<c��<щ�<)�<��<�Q�<���<�^�<���<�P�< ��<)�<,��<P�<�@�<���<ߵ<1&�<Lh�<���<�ݮ<��<�A�<�m�<���<%��<�ۣ<��<��<p/�<�F�<\�<�o�<J��<{��<8��<|��<s��<Č<Z͊<yՈ<�܆<w�<t�<��<~�}<~�y<��u<��q<n�m<S�i<��e<�b<y
^<FZ<	V<%R<Z0N<�<J<�JF<�YB<�j><K}:<��6<_�2<��.<[�*<x�&<#<�E<�p<�<�<�<�Q<l�<��<:<�*�;���;"��;f��;0��;z��;���;��;�&�;�{�;#�;*j�;��;���;B��;�t�;C{�;��;~݄;�r~;ees;E�h;�];R�S;�dI;�n?;"�5;�$,;��";��;��;��;p��:��:��:|��:���:���:���:S��:[0�:��g:��K:0:g�:x��9�߾9wl�9�-9r�8������*Gg�]�����չ $�\&��2���J�Nb�_y��E���ʓ��D��粪�a���s��y�̺�غ<i㺢���������2�����^�X���{��$�؉)�/�ȋ4�;	:�Ѕ?�hE��}J���O�hyU�:�Z�5{`�S�e��k�qq���v�l|�dҀ������Z��{���ዻ1���Qh���+��������  �  X�=�8=��=Y�=�,=+�=:y= =�� = j =B =�h�<���<Z��<�E�<%��<��<� �<&i�<��<��<�>�<U��<��<��<�O�<p��<��<��<�O�<$��<T��<H�<+>�<�v�<K��<v��<�<:L�<�}�<��<+��<�<�-�<#S�<�u�<x��<ڱ�<���<��<���<���<e	�<�<q�<[�<��<���<��< ��<��<S��<Ig�<�7�<��<���<���<k5�<��<D��<C(�<!��<�P�<���<r]�<���<\O�<���<�'�<�<F�<�?�<đ�<J޵<�%�<�g�<=��<�ݮ<�<B�<�m�<.��<�<{ܣ<!��<�<�0�<�G�<8]�<�p�<[��<���<��<D��< ��<�Č<�͊<�Ո<p܆<4�<�<�<�}<��y<��u<��q<�m<�i<8�e<Rb<"^<Z<'V<J#R<�.N<�;J<�IF<[YB<�j><r}:<>�6<H�2<��.<��*<.�&<2!#<H<>s<\�<w�<L<�S<��<��<�;<�-�;>��; ��;���;���;��;���;���;�$�;'y�;��;�f�;��;[��;ą�;=p�;w�;Ù�;�ل;=l~;_s;�h;g�];�S;�bI;�n?;n�5;�',;��";`�;K�;;���:.,�:~��:���:��:Q��:咟:�ǐ:?�:F�g:I�K:�+0:��:���9߾9�]�9J�,9�r�8��3�H�g�4��uֹ�G�jM��3���J��3b��}y��S���ד�SO�����P��Vw����̺�غ�b㺪����ܐ�1+���FV�����r�#�#��)��/�g�4�c:��?��D�zJ���O��xU���Z�g}`�@f�k�k�Rq�r�v��#|��ր�P���b_��a#���拻˩���l��/��������  �  �=[8=r�=P�=�,=P�=my=M=�� =oj =� =�i�<���<���<	G�<I��<G��<�!�<j�<Ǳ�<���<&?�<���<]��<�<�O�<(��<���<��<!O�<F��<F��<7�<=�<�u�<#��<G��<�<'K�<�|�<��<���<��<-�<�R�<�u�<���<)��<8��<���<���<d �<Y
�<%�<��<��<��<��<=��<���<��<��<�g�<O8�<�<���<���<45�<���<���<�'�<;��<�O�<y��<L\�<v��<N�<q��<�&�<͉�<�<�>�<ᐷ<�ݵ<%%�<�g�<��<�ݮ<J�<XB�<qn�<֖�<���<Vݣ<��<%�<�1�<I�<b^�<�q�<x��<{��<���<��<���<�Č<�͊<�Ո<c܆<��<��<��<��}<�y<��u<c�q<��m<��i<��e<��a<�^<�Z<V<�!R<N-N<q:J<�HF<�XB<`j><�}:<Β6<�2<��.<b�*<��&<##<<J<�u<¥<��<�<<V<�<��<�=<�0�;���;���;��;G��;ܢ�;޹�; ��;�"�;Fv�;��;�b�;���; ��;1��;�k�;�r�;���;�Մ;e~;�Xs;[�h;��];�S;�aI;�n?;q�5;X*,;o�";�;��;
;���:�>�:���:G��:��:i��:K��:Zא:3M�:�	h:�K:x;0:��:}�9�޾9�S�9q�,9m��8�����w�v-h��x���bֹAm��r��C3���J��Ub�ݟy��a���䓺X��D���d!��Py����̺�غ@]�y��P�����$���M�����h���#��w)���.��{4�p�9�|y?�*�D��vJ�Y�O�5wU�d�Z�"`��f�{�k��q��v��+|��ڀ�����d���'��V닻*����p���3��[���幙��  �  Ӑ=(8=V�=A�=�,=m�=�y=�=M� =�j =+ =�j�<Ǵ�<���<.H�<\��<N��<�"�<�j�<���<w��<�?�<��<���<
�<zO�<��<*��<e�<kN�<z��<X��<@�<�;�<�t�<��<%��<�<0J�<�{�<W��<���<�<�,�<�R�<�u�<ϕ�<m��<���<U��<5��<C�<B�< �<��<��<��<��<;��<���<δ�<���<�h�<�8�<G�<���<���<5�<0��<*��<�&�<m��<�N�<s��<@[�<A��<�L�<I��<v%�<�<�<�=�<��< ݵ<�$�<0g�<ݤ�<�ݮ<j�<�B�<�n�<k��<n��<4ޣ<	��<(�<�2�<2J�<o_�<�r�<t��<`��<Т�<���<=��<dŌ<4Ί<�Ո<I܆<��<M�<�<<�}<��y<�u<r�q<��m<R�i<��e<��a<�^<�Z<7V<�R<�+N<[9J<HF<`XB<j><�}:<?�6<�2<��.<��*<�'<�$#<=L<�w<��<^�<�<eX<�<��<\?<�3�;I��;���;���;���;���;��;���;� �;�s�;�ݵ;5_�;���;��;}�;�g�;2n�;���;�ф;�^~;#Ss;j�h;�];ÈS;�`I;�n?;��5;�,,;��";	�;i�;K;�	�:�N�:���:���:=1�:�̮:���:k�:v[�:Dh:�K:�L0::�:��9�ܾ9gK�9��,9�x�8'< ���[�h�����:�ֹ{�����Bf3�+K��tb���y��n����a���Ȫ��%��E{���̺�غ�W�H��b���N����l���D�D���_�J�#�|o)���.��t4���9�Qt?�Y�D�'sJ�j�O��vU�E�Z���`��f���k��q�D�v��2|��ހ������h��A,���_����t��07�����������  �  ��=�7=7�=:�=-=�=�y=�=�� =.k =� =�k�<���<���<I�<T��</��<�#�<�k�<2��<��<@�<]��<���<�<]O�<���<���<��<�M�<���<���<S�<;�<�s�<��<C��<�<YI�<�z�<���<P��<��<�,�<�R�<�u�<��<���<��<���<���<��<�<��<��<��<��<��<��<���<���<c��<�h�<9�<x�<
��<���<�4�<���<���<I&�<���<N�<���<:Z�<M��<�K�<C��<y$�<�<@�<=�<j��<dܵ<($�<�f�<���<�ݮ<x�<�B�<Jo�<ꗧ<��<�ޣ<���<�<�3�<K�<a`�<�s�<L��<4��<���<R��<���<�Ō<_Ί<�Ո<G܆<��<��<��< �}<"�y<��u<��q<��m<��i<��e<��a<�^<
Z<�V<vR<�*N<U8J<]GF<�WB<�i><�}:<��6<��2<��.<��*<�'<�&#<�M<�y<�</�<�<=Z<��<q�<�@<6�;��;��;���;��;h��;L��;\��;��;�q�;�ڵ;A\�;f��;t��;~y�;d�;�j�;C��;�΄;�X~;�Ms;K}h;��];ՆS;`_I;o?;��5;�.,;��";�;��;1;c�:~\�:B��:���:�?�:ܮ:dß:
��:~g�:�4h:�L:�W0:�:�9r޾9�>�92u,9��8{U��*�Z�h��ꥹ��ֹ�����3��#K�Βb�O�y�{������fj��	Ϫ��)���}��S�̺	غS㺍�������������=�����X���#�h)��.�$n4�'�9�mo?���D��pJ�!�O��uU�h�Z���`�:f�k�k�� q��v��8|�7※����.l��20��l�9���Tx��B:��l��������  �  ^�=�7= �=5�=-=��=�y=�=�� =jk =� =7l�<P��<A �<�I�<��<���<W$�<Hl�<���<~��<i@�<���<���<#�<KO�<o��<|��<p�<aM�<)��<���<� �<`:�<�r�<M��<���<V�<�H�<_z�<)��<���<G�<<,�<sR�<�u�<���<��<Y��<-��<Y��<p�<��<��<.�<=�<w	�<���<���<K��<���<ޒ�<\i�<e9�<��<��<~��<�4�<���<J��<�%�<-��<{M�<���<zY�<���<K�<x��<�#�<��<��<w<�<鎷<�۵<�#�<�f�<���<�ݮ<��<#C�<�o�<W��<���<uߣ<y��<��<f4�<�K�<a�<[t�<<ϕ�<���<հ�<��<ƌ<�Ί<ֈ<A܆<l�<��<3�<G�}<�y<c�u<u�q<~�m<-�i<�e<i�a<q ^<�Z<rV<bR<�)N<u7J<�FF<zWB<�i><~:<�6<#�2<z�.<��*<�'<�'#<KO<�z<k�<��<g<�[<	�<��<�A<8�;h��;]��;h��;m��;L��;���;C��;3�;�o�;�ص;Z�;��;��;�v�;a�;[h�;���;�̄;hT~;EJs;.zh;��];�S;m^I;Co?;_�5;�0,;�";!�;��;;~!�: g�:��:O �:�K�:��:�͟:��:(o�:�Dh:)L:}a0:�:>"�9�߾97�9�T,9T��8)��h�}Ei�m���׹k�������3�8K���b���y�-���+��q��CԪ��-�� ����̺غ�N㺳����3{�x�����8�
��?S���#�c)���.�Pi4�i�9�]k?�"�D�4nJ�J�O��uU���Z��`�wf���k�_$q��v��=|��䀻`����n��`3��%���㸎��z���<�����������  �  J�=�7=�=/�=-=��=�y= =�� =�k = =�l�<϶�<� �<;J�<s��<P��<�$�<�l�<��<���<�@�<���<���<�<CO�<\��<U��<?�<M�<؉�<���<; �<�9�<sr�<ߩ�<��<��<LH�<�y�<۩�<���<%�<!,�<nR�<�u�< ��<���<��<i��<���<��<�<�<��<��<�	�<'��<,��<���<j��<��<�i�<�9�<��<!��<h��<�4�<t��<��<�%�<ؼ�<M�<s��<Y�<��<�J�<���<A#�<���<&�<<�<���<�۵<�#�<zf�<}��<�ݮ<��<5C�<�o�<���<ѽ�<�ߣ<���<�<�4�<>L�<�a�<�t�<b��<2��<a��<��<E��<&ƌ<�Ί<ֈ<3܆<g�<��<�<��}<w�y<��u<��q<��m<�i<;�e<[�a<��]<�Z<�V<�R<)N< 7J<vFF<dWB<�i><�}:<�6<V�2<��.<O�*<�'<�(#<,P<�{<L�<��<G<�\<�<~�<�B<9�;T��;���;׭�;S��;H��;u��;���;��;�n�;�׵;xX�;J�;1��;�t�;p_�;Yf�;���;�ʄ;vQ~;�Gs;�wh;��];1�S;h^I;�n?;̵5;�1,;c�";�;��;�;�'�:�n�:~�:o�:�R�:!�:�՟:z�:<v�:�Lh:�#L:�f0:0:&�9j۾9�5�9�F,9͊�8������ti��,��q&׹������3�HK�<�b���y�^���"��qt���֪�%/��O����̺�غM㺠��	����x��J���4����WO�z�#�_)�h�.�:f4�4�9��i?�D�D�CmJ���O�|uU�!�Z��`�df��k��&q���v��@|�~总$����p��5��9��������|��V>��������  �  @�=�7=�=,�=-=��=z=) =�� =�k = =�l�<��<� �<dJ�<���<y��<�$�<�l�< ��<���<�@�<ǅ�<���< �<?O�<@��<3��<'�<�L�<���<d��<& �<�9�<Mr�<ĩ�<���<��<*H�<�y�<ɩ�<z��<�<�+�<YR�<�u�<��<���<���<���<���<�<�<+�<��<��<
�<U��<G��<���<���<0��<�i�<�9�<��<2��<a��<�4�<T��<	��<j%�<���<�L�<K��<�X�<���<�J�<ҹ�<#�<~��<��<�;�<k��<�۵<{#�<]f�<u��<�ݮ<��<9C�<�o�<���<꽥<�ߣ<���<A�<�4�<bL�<�a�<u�<v��<9��<���<��<l��<3ƌ<�Ί<ֈ<0܆<M�<n�<��<`�}<V�y<Z�u<[�q<k�m<��i<�e<�a<F�]<�Z<UV<�R<�(N<�6J<(FF<1WB<�i><~:<<�6<o�2<<�.<v�*<'<�(#<QP<W|<��<��<�<�\<��<��<�B<t9�;���;���;7��;���;@��;��;F��;5�;0n�;\׵;�W�;��;���;`t�;_�;�e�;���;Nʄ;�P~;xGs;
wh;}�];�S;�]I;�n?;~�5;�1,;��";+�;j�;�;�'�:`p�:��:�	�:U�:�:]ן:E�:=x�:�Oh:b'L:�h0:,:�*�9)ھ9,2�9�7,9�x�8�����Ui�
6��p*׹�������3�	MK�R�b���y�-���[���u���ت��0�����C�̺Xغ�L������w�v�;���3�}��2N���#�}])���.�f4��9�*i?��D��lJ�5�O��tU�=�Z��`��f���k��'q��v��A|��总�����q��f5������/����|���>�� �����  �  J�=�7=�=/�=-=��=�y= =�� =�k = =�l�<϶�<� �<;J�<s��<P��<�$�<�l�<��<���<�@�<���<���<�<CO�<\��<U��<?�<M�<؉�<���<; �<�9�<sr�<ߩ�<��<��<LH�<�y�<۩�<���<%�<!,�<nR�<�u�< ��<���<��<i��<���<��<�<�<��<��<�	�<'��<,��<���<j��<��<�i�<�9�<��<!��<h��<�4�<t��<��<�%�<ؼ�<M�<s��<Y�<��<�J�<���<A#�<���<&�<<�<���<�۵<�#�<zf�<}��<�ݮ<��<5C�<�o�<���<ѽ�<�ߣ<���<�<�4�<>L�<�a�<�t�<b��<2��<a��<��<E��<&ƌ<�Ί<ֈ<3܆<g�<��<�<��}<w�y<��u<��q<��m<�i<;�e<[�a<��]<�Z<�V<�R<)N< 7J<wFF<dWB<�i><�}:<�6<V�2<��.<O�*<�'<�(#<,P<�{<L�<��<G<�\<�<~�<�B<9�;T��;���;׭�;S��;H��;u��;���;��;�n�;�׵;xX�;J�;1��;�t�;p_�;Yf�;���;�ʄ;vQ~;�Gs;�wh;��];1�S;h^I;�n?;̵5;�1,;c�";�;��;�;�'�:�n�:~�:o�:�R�:!�:�՟:z�:<v�:�Lh:�#L:�f0:0:&�9j۾9�5�9�F,9͊�8������ti��,��q&׹������3�HK�<�b���y�^���"��qt���֪�%/��O����̺�غM㺠��	����x��J���4����WO�z�#�_)�h�.�:f4�4�9��i?�D�D�CmJ���O�|uU�!�Z��`�df��k��&q���v��@|�~总$����p��5��9��������|��V>��������  �  ^�=�7= �=5�=-=��=�y=�=�� =jk =� =7l�<P��<A �<�I�<��<���<W$�<Hl�<���<~��<i@�<���<���<#�<KO�<o��<|��<p�<aM�<)��<���<� �<`:�<�r�<M��<���<V�<�H�<_z�<)��<���<G�<<,�<sR�<�u�<���<��<Y��<-��<Y��<p�<��<��<.�<=�<w	�<���<���<K��<���<ޒ�<\i�<e9�<��<��<~��<�4�<���<J��<�%�<-��<{M�<���<zY�<���<K�<x��<�#�<��<��<w<�<鎷<�۵<�#�<�f�<���<�ݮ<��<#C�<�o�<W��<���<uߣ<y��<��<f4�<�K�<a�<[t�<<ϕ�<���<հ�<��<ƌ<�Ί<ֈ<A܆<l�<��<3�<G�}<�y<c�u<u�q<~�m<-�i<�e<i�a<q ^<�Z<rV<bR<�)N<u7J<�FF<zWB<�i><~:<�6<#�2<z�.<��*<�'<�'#<KO<�z<k�<��<g<�[<	�<��<�A<8�;h��;]��;h��;m��;L��;���;B��;2�;�o�;�ص;Z�;��;��;�v�;a�;Zh�;���;�̄;hT~;DJs;.zh;��];�S;m^I;Co?;_�5;�0,;�";!�;��;;~!�: g�:��:O �:�K�:��:�͟:��:(o�:�Dh:)L:}a0:�:>"�9�߾97�9�T,9T��8)��h�}Ei�m���׹k�������3�8K���b���y�-���+��q��CԪ��-�� ����̺غ�N㺳����3{�x�����8�
��?S���#�c)���.�Pi4�i�9�]k?�"�D�4nJ�J�O��uU���Z��`�wf���k�_$q��v��=|��䀻`����n��`3��%���㸎��z���<�����������  �  ��=�7=7�=:�=-=�=�y=�=�� =.k =� =�k�<���<���<I�<T��</��<�#�<�k�<2��<��<@�<]��<���<�<]O�<���<���<��<�M�<���<���<S�<;�<�s�<��<C��<�<YI�<�z�<���<P��<��<�,�<�R�<�u�<��<���<��<���<���<��<�<��<��<��<��<��<��<���<���<c��<�h�<9�<x�<
��<���<�4�<���<���<I&�<���<N�<���<:Z�<M��<�K�<C��<y$�<�<@�<=�<k��<dܵ<($�<�f�<���<�ݮ<x�<�B�<Jo�<ꗧ<��<�ޣ<���<�<�3�<K�<a`�<�s�<L��<4��<���<R��<���<�Ō<_Ί<�Ո<G܆<��<��<��<�}<"�y<��u<��q<��m<��i<��e<��a<�^<
Z<�V<vR<�*N<U8J<]GF<�WB<�i><�}:<��6<��2<��.<��*<�'<�&#<�M<�y<�</�<�<=Z<��<q�<�@<6�;��;��;���;��;g��;L��;\��;��;�q�;�ڵ;A\�;f��;t��;}y�;d�;�j�;B��;�΄;�X~;�Ms;K}h;��];ՆS;`_I;o?;��5;�.,;��";�;��;1;c�:~\�:B��:���:�?�:ܮ:dß:
��:~g�:�4h:�L:�W0:�:�9r޾9�>�92u,9��8{U��*�Z�h��ꥹ��ֹ�����3��#K�Βb�O�y�{������fj��	Ϫ��)���}��S�̺	غS㺍�������������=�����X���#�h)��.�$n4�'�9�mo?���D��pJ�!�O��uU�h�Z���`�:f�k�k�� q��v��8|�7※����.l��20��l�9���Tx��B:��l��������  �  Ӑ=(8=V�=A�=�,=m�=�y=�=M� =�j =+ =�j�<Ǵ�<���<.H�<\��<N��<�"�<�j�<���<w��<�?�<��<���<
�<zO�<��<*��<e�<kN�<z��<X��<@�<�;�<�t�<��<%��<�<0J�<�{�<W��<���<�<�,�<�R�<�u�<ϕ�<m��<���<U��<5��<C�<B�< �<��<��<��<��<;��<���<δ�<���<�h�<�8�<G�<���<���<5�<0��<*��<�&�<m��<�N�<s��<@[�<A��<�L�<I��<v%�<�<�<�=�<��< ݵ<�$�<0g�<ݤ�<�ݮ<j�<�B�<�n�<k��<n��<4ޣ<	��<(�<�2�<2J�<o_�<�r�<t��<`��<Т�<���<=��<dŌ<4Ί<�Ո<I܆<��<M�<�<<�}<��y<�u<r�q<��m<R�i<��e<��a<�^<�Z<7V<�R<�+N<[9J<HF<`XB<j><�}:<?�6<�2<��.<��*<�'<�$#<=L<�w<��<^�<�<eX<�<��<\?<�3�;I��;���;���;���;���;��;���;� �;�s�;�ݵ;5_�;���;��;}�;�g�;2n�;���;�ф;�^~;#Ss;j�h;�];ÈS;�`I;�n?;��5;�,,;��";	�;i�;K;�	�:�N�:���:���:=1�:�̮:���:k�:v[�:Dh:�K:�L0::�:��9�ܾ9gK�9��,9�x�8'< ���[�h�����:�ֹ{�����Bf3�+K��tb���y��n����a���Ȫ��%��E{���̺�غ�W�H��b���N����l���D�D���_�J�#�|o)���.��t4���9�Qt?�Y�D�'sJ�j�O��vU�E�Z���`��f���k��q�D�v��2|��ހ������h��A,���_����t��07�����������  �  �=[8=r�=P�=�,=P�=my=M=�� =oj =� =�i�<���<���<	G�<I��<G��<�!�<j�<Ǳ�<���<&?�<���<]��<�<�O�<(��<���<��<!O�<F��<F��<7�<=�<�u�<#��<G��<�<'K�<�|�<��<���<��<-�<�R�<�u�<���<)��<8��<���<���<d �<Y
�<%�<��<��<��<��<=��<���<��<��<�g�<O8�<�<���<���<55�<���<���<�'�<;��<�O�<y��<L\�<v��<N�<q��<�&�<͉�<�<�>�<␷<�ݵ<%%�<�g�<��<�ݮ<J�<XB�<rn�<֖�<���<Vݣ<��<%�<�1�<I�<b^�<�q�<x��<{��<���<��<���<�Č<�͊<�Ո<c܆<��<��<��<��}<�y<��u<c�q<��m<��i<��e<��a<�^<�Z<V<�!R<N-N<q:J<�HF<�XB<`j><�}:<Β6<�2<��.<b�*<��&<##<<J<�u<å<��<�<<V<�<��<�=<�0�;���;���;��;G��;ܢ�;޹�; ��;�"�;Fv�;��;�b�;���; ��;1��;�k�;�r�;���;�Մ;e~;�Xs;[�h;��];�S;�aI;�n?;q�5;X*,;o�";�;��;
;���:�>�:���:G��:��:i��:K��:Zא:3M�:�	h:�K:x;0:��:}�9�޾9�S�9q�,9m��8�����w�v-h��x���bֹAm��r��C3���J��Ub�ݟy��a���䓺X��D���d!��Py����̺�غ@]�y��P�����$���M�����h���#��w)���.��{4�p�9�|y?�*�D��vJ�Y�O�5wU�d�Z�"`��f�{�k��q��v��+|��ڀ�����d���'��V닻*����p���3��[���幙��  �  X�=�8=��=Y�=�,=+�=:y= =�� = j =B =�h�<���<Z��<�E�<%��<��<� �<&i�<��<��<�>�<U��<��<��<�O�<p��<��<��<�O�<$��<T��<H�<+>�<�v�<K��<v��<�<:L�<�}�<��<+��<�<�-�<#S�<�u�<x��<ڱ�<���<��<���<���<e	�<�<q�<[�<��<���<��< ��<��<S��<Ig�<�7�<��<���<���<k5�<��<D��<C(�<!��<�P�<���<r]�<���<\O�<���<�'�<���<F�<�?�<đ�<K޵<�%�<�g�<=��<�ݮ<�<B�<�m�<.��<�<{ܣ<!��<�<�0�<�G�<8]�<�p�<[��<���<��<D��< ��<�Č<�͊<�Ո<p܆<3�<�<�<�}<��y<��u<��q<�m<�i<8�e<Rb<"^<Z<'V<J#R<�.N<�;J<�IF<[YB<�j><r}:<>�6<H�2<��.<��*<.�&<2!#<H<>s<\�<w�<L<�S<��<��<�;<�-�;>��; ��;���;���;��;���;���;�$�;&y�;��;�f�;��;[��;ą�;<p�;w�;Ù�;�ل;=l~;_s;�h;g�];�S;�bI;�n?;n�5;�',;��";`�;K�;;���:.,�:~��:���:��:Q��:咟:�ǐ:?�:F�g:I�K:�+0:��:���9߾9�]�9J�,9�r�8��3�H�g�4��uֹ�G�jM��3���J��3b��}y��S���ד�SO�����P��Vw����̺�غ�b㺪����ܐ�1+���FV�����r�#�#��)��/�g�4�c:��?��D�zJ���O��xU���Z�g}`�@f�k�k�Rq�r�v��#|��ր�P���b_��a#���拻˩���l��/��������  �  ��=�8=��=h�=�,=
�=�x=�==� =�i =� =�g�<}��<)��<�D�<���<��<��<*h�<��<o��<>�<��<���<��<�O�<���<��<!�<�P�<��<F��<h�<K?�<x�<���<���<7�<9M�<h~�<ĭ�<���<��<�-�<cS�<�u�<X��<���<Q��<���<���<���<U�<��<R�<0�<o�<���<��<���<8��<���<�f�<s7�<k�<���<���<�5�<c��<щ�<)�<��<�Q�<���<�^�<���<�P�< ��<)�<,��<P�<�@�<���<ߵ<1&�<Lh�<���<�ݮ<��<�A�<�m�<���<%��<�ۣ<��<��<p/�<�F�<\�<�o�<J��<{��<8��<|��<s��<Č<Z͊<yՈ<�܆<w�<t�<��<~�}<~�y<��u<��q<n�m<S�i<��e<�b<y
^<FZ<
V<%R<Z0N<�<J<�JF<�YB<�j><K}:<��6<_�2<��.<[�*<x�&<#<�E<�p<�<�<�<�Q<l�<��<:<�*�;���;"��;f��;0��;y��;���;��;�&�;�{�;"�;)j�;��;���;A��;�t�;C{�;��;~݄;�r~;ees;D�h;�];R�S;�dI;�n?;"�5;�$,;��";��;��;��;p��:��:��:{��:���:���:���:S��:[0�:��g:��K:0:g�:x��9�߾9wl�9�-9r�8������*Gg�]�����չ $�\&��2���J�Nb�_y��E���ʓ��D��粪�a���s��y�̺�غ<i㺢���������2�����^�X���{��$�؉)�/�ȋ4�;	:�Ѕ?�hE��}J���O�hyU�:�Z�5{`�S�e��k�qq���v�l|�dҀ������Z��{���ዻ1���Qh���+��������  �  �=�8=��=o�=�,=��=�x=y=�� =.i =I =�f�<o��<
��<�C�<Ռ�<��<��<Ig�<R��<���<�=�<���<���<��<�O�<���<���<��<XQ�<ގ�<,��<c�<Y@�<!y�<���<���<@�<,N�<O�<z��<{��<0�<2.�<�S�<�u�<8��<=��<���<���<;��<���<h�<��<6�<!�<d�<���< ��<��<m��<Ԏ�<#f�<�6�<)�<���<���<�5�<���<m��<�)�<���<�R�<���<�_�<��<�Q�<&��<3*�<<��<L�<�A�<`��<�ߵ<�&�<�h�<���<�ݮ<��<jA�<m�<�<k��<�ڣ<&��<�<S.�<�E�<�Z�<sn�<S��<���<k��<Ĭ�<㸎<�Ì<͊<XՈ<�܆<��<��<<�<��}<�y<��u<��q<��m<}�i< f<�b<�^<AZ<�V<�&R<�1N<�=J<{KF<nZB<�j><}:<P�6<��2<q�.<��*<��&<;#<�C<�n<��<��<{<nO<c�<��<k8<�'�;���;m��;k��;���;���;a��;���;�(�;V~�;U�;�m�;t	�;���;F��;!y�;]�;	��;�;�y~;�js;ߔh;I�];ĒS;�eI;�n?;ܭ5;!",;��";��;��;�;6��:�:��:%��:��:_��:�q�:��:-#�:�g:�K:�0:��:���9oݾ9)w�9�?-9�|�8P���L�n�f����!�չ��?���2��xJ���a��Ay��7��S���;��ݪ��,��r����̺Gغ�n�ܷ���������9�c���f�f��w���$�o�)��/�3�4��:�}�?��E�9�J���O�^zU���Z��y`�3�e�?�k�~q�H�v�C|��΀������V������݋����od��=(��Q얻~����  �  $�=#9=��=y�=�,=��=�x=8=�� =�h =� =�e�<y��<"��<�B�<��<��<��<�f�<���<0��<=�<<��<{��<��<P�<)��<J��<+�<�Q�<���< ��<;�<GA�<z�<���<���<�<O�<��<#��<��<��<v.�<�S�<�u�<��<���<r��<\��<���<��<��<�<P�<-
�<n�<���<0��<:��<���<4��<�e�<�6�<� �<Z��<р�<6�<��<ӊ�<>*�<~��<�S�<���<�`�<��<�R�<$¿<5+�<$��<4�<nB�<��<7�<''�<�h�<ץ�<ޮ<��<,A�<�l�<l��<���<�٣<T��<�<u-�<�D�<Z�<�m�<h�<Ï�<���<,��<[��<9Ì<�̊<=Ո<�܆<��<#�<��<��}<]�y<�u<X�q<J�m<t�i<�f<�b<h^<Z<�V<(R<�2N<�>J<'LF<�ZB<#k><�|:<Ր6<�2<m�.<��*<Z�&<�#<�A<�l<��<��<�<eM<��<T�<�6<F%�;���;���;J��;F��;���;Լ�;���;o*�;���;��;�p�;��;¢;ؑ�;}|�;��;T��;Y�;�~;�os;Șh;��];��S;2fI;�n?;Q�5;�,;E�";�;��;��;��:���:*��:���:ؽ:�u�:�b�:���:q�:��g:<�K:��/:4�:F��9A߾9}�9�]-9Iԍ8�O�����tf�����A]չ�����9�2��ZJ���a��&y�},��9����3������$���p��a�̺�"غIs����-���?�#���n�r��X��$� �)�./�z�4��:�2�?��	E��J���O�"{U�_�Z��x`���e�}k��q��v��|�ˀ�
����R��m���ً�y����`��%���閻����  �  M�=I9=��=~�=�,=��=zx==b� =�h =� =e�<Ѯ�<s��<�A�<I��<]��<[�<�e�<��<���<�<�<���<Q��<��< P�<g��<���<��<yR�<��<���<��<�A�<�z�<9��<M��<��<�O�<���<���<t��<��<�.�<�S�<�u�<���<���<��<���<'��<���<	�<b�<��<o	�<��<7��<���<���<��<���<:e�<F6�<� �<G��<���</6�<Z��<(��<�*�<��<T�<B��<^a�<���<�S�<�¿<�+�<؎�<��<�B�<���<��<}'�<-i�<�<ޮ<��<�@�<Kl�<��<J��<m٣<���<[�<�,�<�C�<NY�<�l�<�~�<0��<��<���<뷎<�<�̊<+Ո<�܆<��<m�<��<��}<U�y<:�u<��q<��m<��i<.f<?	b<�^<MZ<�V<)R<�3N<?J<�LF<"[B<;k><�|:<u�6<I�2<��.<��*<I�&<v#<�@<xk<J�<-�<?<�K<J�<�<�5<l#�;���;���;w��; ��;���;���;���;�+�;v��;��;�r�;�;Ģ;���;,�;���;���;��;f�~;Uss;�h; �];��S;�fI;�n?;t�5;�,;r�";��;��;��;���:���:Ό�:U��:�˽:�k�:JW�:���:5�:��g:�K:&�/:7�:`��9��9���9�-9 �8��򷗸��6f�^[��4չ��������2��EJ��a�:y�%������-��𠪺����o����̺%غ�w�W��G�����D����5t�������$�6�)�o /��4��:���?�pE���J�� P��{U��Z�Bw`�h�e��zk��p�2�v�p
|��Ȁ�|����O������֋�󚎻x^���"���疻)����  �  i�=U9=�=z�=�,=��=hx=�=8� =dh =d =�d�<[��<���<cA�<�<���<��<�e�<̭�<s��<�<�<ڂ�<K��<��<#P�<���<���<��<�R�<p��<���<T�<iB�<:{�<���<���<?�<P�<��<��<���<�<�.�<�S�<�u�<��<���<���<���<���<-��<��<�
�<.�<��<<�<���<��<;��<ï�<s��<�d�<"6�<� �<G��<Ԁ�<F6�<|��<Z��<�*�<S��<�T�<���<�a�<F��<T�<cÿ<k,�<X��<K�<iC�<䔷<��<�'�<Oi�< ��<�ݮ<��<�@�<.l�<���<���<
٣<L��<��<J,�<C�<�X�<bl�<R~�<���<ʝ�<h��<���<�<�̊< Ո<�܆<�<��<"�<<�}<�y<�u<t�q<��m<��i<.f<
b<�^<*Z<� V<�)R<O4N<�?J<�LF<U[B<.k><�|:<b�6<�2<=�.<8�*<��&<�#<�?<�j<<�<H�<'
<K<V�<5�<#5<"�;��;(��;D��;���;���;��;-��;�,�;;��;"�;Vt�;��;aƢ;=��;��;H��;���;@�;��~;�us;��h;X�];b�S;[gI;*n?;2�5;�,;�";��;�;B�;]��:���:���:�x�:�Ľ:Kc�:�P�:4��:��:��g:��K:*�/:��:��9�ܾ9���9h�-9�K�8��)����e�A���չ]�������2�m6J�	�a��y���V����)������J
��,o����̺Z%غ7y�p�� ������G�����w������$��)��#/���4�~:�9�?��E���J�P��{U�|�Z��v`���e�yk�m�p�X�v�$|��ƀ�����#N�����KՋ������\�� !��<斻U����  �  ߏ=76=z�=��=R(=��=Bs=t=Z� =.b =� =�V�<Q��<���</0�<%x�<��<j�<bN�<���<���<; �<�d�<?��<���<�,�<�l�<b��<���<�'�<�c�<���<L��<I�<�E�<"{�<���<���<��<B?�<zk�<���<&��<���<X�<�#�<�?�<�X�<kn�<~��<��<���<U��<.��<���<���<<��<��<�m�<1T�<@5�<��<���<#��<�}�<@�<���<E��<�]�<��<���<J=�<R��<kZ�<��<�\�<���<�E�<��<e�<�u�<�ϸ<$�<<s�<��<��< B�<�}�<δ�<��<�<wB�<�j�<���<ʱ�<Yџ<R�<L	�<"�<9�<tN�<�a�<6t�<ۄ�<J��<E��<��<���<Dņ<�΄<Eׂ<J߀<��}<��y<	�u<��q<o�m<�j<�f<� b<z-^<�:Z<UIV<�XR<iN<�{J<w�F<G�B<ٹ><��:<g�6<	3<�(/<�J+<�p'<љ#<��<��<s0<�l<t�<h�<aD	<ј<T�<@��;]��;�c�;�V�;�Y�;o�;%��;��;'�;�~�;.��;d��;�+�;��;�;���;���; �;)*�;(��;�x;>,m;�b;& X;��M;��C;<!:;)�0;�$';��;��;\;�{;��:B��:�J�:�g�:�ӵ:c��:.��:Cو:��t:-KX:F<:9� :`h:��9��9�V9���8�-7j[��oB�j)��^�Ĺ����#��D+��7C�\�Z�@�r��������^[����~��f���Xwʺ�պ+T��������r\����K��6:�R���c#���(��}.��4���9��?��D��J���O�"U��Z��-`���e�+>k���p�LUv�5�{�����C~��GE��	��uӋ������b���*��p�s����  �  ď=;6=y�=��=V(=��=Js=x=i� =8b =� =�V�<Z��<���<?0�<Jx�<��<�<�N�<��<���<A �<�d�<M��<���<r,�<�l�<Z��<���<�'�<bc�<���<N��<;�<�E�<{�<���<���<��<.?�<ak�<W��<��<��<B�<�#�<�?�<�X�<yn�<���<��<���<u��<"��<���<ƛ�<N��<��<�m�<NT�<[5�<��<��<0��<�}�<%@�<���<+��<�]�<��<L��<.=�<4��<mZ�<���<�\�<���<�E�<��<b�<�u�<�ϸ<�#�<�r�<���<��<B�<�}�<۴�<��<�<�B�<�j�<���<㱡<Xџ<w�<Z	�<3"�<%9�<rN�<b�<Kt�<���<T��<T��<'��<���<5ņ<�΄<Rׂ<߀<O�}<��y<��u<��q<B�m<�j<mf<� b<R-^<�:Z<KIV<�XR<7iN<4{J<��F<C�B<��><�:<��6<'	3<�(/<�J+<�p'<�#<��<��<�0<�l<®<p�<�D	<�<��<­�;x��;d�;W�;Z�;�n�;K��;��;4�;u~�;���;x��;�+�;t�;j;E��;w��;��;=*�;߇�;�x;�*m;�b;� X;8�M;a�C;�!:;�0;%';4�;l�; ;�|;��:΂�:>L�: i�:�յ:���:��:�ڈ:�t:�NX:�G<:s� :7j:�9{�9��V9���8�R 7Ru���|B�^(���Ĺd���&'��F+�&9C�|�Z�ɟr����?���b_����G}�����Ewʺ�պ�Rẅ�����)���[����I��9�����b#�U�(��}.��4��9�?���D��J��O��!U�h�Z�.`��e��?k���p�;Vv���{������~���E������Ӌ�
����b���*���� ����  �  ��=16=p�=��=X(=��=[s=�=�� =Ob =� = W�<���<V��<�0�<�x�<]��<��<�N�<C��<3��<] �<�d�<N��<���<f,�<�l�<@��<W��<t'�<c�<���<���<��<�E�<�z�<T��<@��<��<�>�<:k�<>��<ټ�<���<*�<�#�<�?�<�X�<�n�<���<=��<��<נ�<u��<��<��<���<x��<n�<�T�<�5�<��<0��<D��< ~�<!@�<���<��<�]�<q�<*��<
=�<���<Z�<���<�\�<��<vE�<���<��<yu�<Kϸ<�#�<�r�<Ѽ�<��<�A�<�}�<մ�<��<+�<�B�<�j�<��<A��<�џ<��<�	�<�"�<�9�<�N�<yb�<|t�<3��<z��<v��<2��<���<:ņ<�΄<Cׂ<�ހ<*�}<!�y<F�u<�q<u�m<!j<�f<�b<�,^<(:Z<�HV<3XR<iN<�zJ<]�F<�B<��><�:<��6<k	3<�(/<hK+<q'<Ě#<\�<m�<�1<�m<��<+�<SE	<��<��<���;���;�d�;-W�;KZ�;�n�;��;���;��;F~�;���;<��;d*�;�;,��;ܲ�;[��;@�;�(�;|��;� x;�)m;ǉb;� X;��M;��C;�!:;��0;�%';��;B�;� ;�;L�:��:�Q�:Hn�:ݵ:ٔ�:X��:�ވ:"�t:�TX:�J<:�� :$j:��9Fߟ9�V9���8���6����T�B�:>���Ĺ�����2�CR+�+DC��[�R�r����a����a������]~��C���qvʺ;�պ�P���n�����<Y��������5�����_#���(�{.��4�\�9�2?���D�zJ���O��!U�C�Z��.`���e�Ak�x�p��Wv�>�{�-���2����F�����ԋ�����d��;,������B����  �  ��=6=`�=��=](=	�={s=�=�� =�b =4 =yW�<;��<���<1�<+y�<���<K�<7O�<���<���<� �<e�<h��<���<m,�<�l�<��<��<'�<�b�<@��<o��<l�<�D�<z�<ԭ�<���< �<w>�<�j�<��<���<���<"�<�#�<�?�<Y�<�n�<��<���<V��<;��<���<��<���<(��<��<�n�<U�<�5�<F�<��<���<2~�<%@�<���<��<�]�<*�<̣�<�<�<q��<�Y�<��<\�<���<�D�<3��<o�<u�<�θ<^#�<}r�<���<��<�A�<�}�<ߴ�<+�<u�<C�<Yk�<j��<���<,ҟ<T�<6
�<#�<:�<HO�<�b�<�t�<���<Δ�<���<[��<ʺ�<@ņ<�΄<ׂ<�ހ<^�}<W�y<��u<1�q<��m<j<�f<�b<�+^<=9Z<�GV<gWR<9hN<KzJ<ӍF<٢B<��>< �:<��6<�	3<�)/< L+<�q'<��#<U�<o�<�2<�n<��<:�<<F	<��<��<8��;\��;�e�;�W�;�Z�;�n�;���;���;��;�|�;7��;ɂ�;�(�;k�;!��;ɰ�;{��;��;Q'�;+��;l�w;A'm;�b;�X;u�M;B�C;F":;M�0;C(';`�;��;E$;�;��:��:MZ�:w�:��:v��:П�:Z�:��t:#_X:�S<:�� :vk:�
�98ߟ9A�V9�U�8�y�6���,�B�	X����Ĺ����wD�tc+�YRC��[�Ͷr�����Ɛ�=f������H�������7vʺ"�պ M���'
��/���U�r�����2�����[#�K�(�$w.�p 4���9�9?� �D��J�c�O�A!U�#�Z�}/`���e�1Ck���p�[v�:�{�캀������H��?��׋�Z����e���-��t���꿙��  �  h�=�5=P�=w�=i(=%�=�s=�=� =�b =~ = X�<��<���<�1�<�y�<���<��<�O�<;��<���<� �<.e�<���<���<O,�<�l�<ë�<���<�&�<9b�<���<���<��<=D�<cy�<��<!��<x�<�=�<Sj�<x��<V��<���<�<�#�<@�<JY�<o�<b��<��<��<͡�<���<.��<]��<��<���<Mo�<�U�<�6�<��<���<���<V~�<M@�<t��<߯�<W]�<��<^��<<�<���<�X�<P��<A[�<���<D�<k��<��<Yt�<Zθ<�"�<r�<=��<]�<�A�<�}�<��<K�<��<lC�<�k�<���<A��<�ҟ<��<�
�<�#�<�:�<�O�<vc�<�u�<���<��<䢌<���<꺈<'ņ<p΄<�ւ<gހ<}�}<^�y<^�u<��q<1�m<j<)f<Pb<<*^<�7Z<�FV<iVR<IgN<�yJ<d�F<��B<y�><N�:<G�6<>
3<*/<�L+<'s'<˜#<��<��<�3<_p<�<��<�G	<��<�<ձ�;���;�f�;�X�;�Z�;�n�;/��;��;��;�z�;m�;r��;4&�;��;X��;��;���;�;�$�;2��;��w;/$m;�b;�X;��M;��C;�#:;ݍ0;*';�;'�;H);Շ;V*�:G��:Lf�:V��:�:��:*��:4�:�t:�iX:[<:� :zq:@�9�ן9�V9��8�E�6�}��cC������ŹE��C[��z+��iC�l/[�m�r��!��Hΐ��k����������� ��Fvʺ��պrJ�@�캃��
��%Q��������,����V#���(��q.���3�"�9�
?���D�J���O�K U���Z�l0`�+�e�OEk�/�p��^v���{����������K����ڋ����h��!0��`��������  �  -�=�5=:�=p�=s(=5�=�s==/� =c =� =�X�<���<V��<�2�<�z�<[��<�	�<}P�<Ŗ�<u��<d!�<|e�<���<���<5,�<bl�<f��<I��<&�<�a�<��<��<��<wC�<�x�<K��<g��<��<<=�<�i�<��<��<J��<��<�#�<.@�<sY�<qo�<��<���<���<~��<]��<��<%��<���<j��<�o�<RV�<47�<1�<M��<��<~~�<f@�<p��<���<]�<e�<��<�;�<"��<&X�<���<gZ�<���<FC�<���<��<�s�<�͸<W"�<�q�<ϻ�<�<�A�<�}�<&��<��<�<�C�<Vl�<���<ﳡ<�ӟ<��<��<�$�<�;�<�P�<%d�<v�<���<���<H��<���<��< ņ<E΄<�ւ<�݀<��}<3�y<��u<h�q<��m<�j<�f<�b<�(^<i6Z<1EV<)UR<ffN<�xJ<��F<3�B<Z�><r�:<��6<�
3<+/<N+<Mt'<.�#<�<��<�5<�q<ų<Y�<I	<K�<-�<A��;���;�g�;uY�;5[�;Nn�;���;���;��;Zy�;�;�}�;z#�;��;m��;#��;���;Cߌ;"�;���;��w;!m;΂b;�X;��M;��C;�$:;]�0;l-';b�;z�;~.;��;�5�:+��:'s�:��:��:9��:���:���:��t:�zX:Yh<:� :�u:��9I͟9�jV9���8}�6����rC�	���W0Ź�B��rt���+��C�]F[�6�r�:,��gՐ��r������������yuʺv�պ"F�������צ��K����ԋ��%�����O#��(�$l.�n�3�s~9��?���D�J���O��U�8�Z��1`���e��Hk���p��cv�V�{�s���ȇ���N����(݋�B���ek���2������qÙ��  �  ��=�5=!�=l�=|(=N�=�s=G=t� =fc =; =�Y�<���<<��<�3�<�{�<.��<y
�<=Q�<]��<���<�!�<�e�<��<��<$,�<,l�<��<���<z%�<�`�<?��<=��<�<�B�<�w�<u��<���<�<�<�<i�<���<���<��<��<�#�<A@�<�Y�<�o�<T��<.��<7��<R��<0��<ڤ�<��<���<?��<�p�<(W�<�7�<��<���<x��<�~�<s@�<o��<���<�\�<�<W��<�:�<n��<cW�<���<�Y�<���<SB�<���<�<�r�<�̸<�!�<q�<s��<� �<uA�<�}�<8��<��<j�<gD�<�l�<S��<Ĵ�<lԟ<��<��<{%�<`<�<|Q�<�d�<�v�<��<��<���<���<��<ņ<΄<Gւ<�݀<��}<��y<��u<��q<��m<=j<�f<b<�&^<�4Z<�CV<�SR<7eN<�wJ<)�F<ȡB<C�><��:<��6<�3<�+/<)O+<�u'<џ#<��<> <�7<�s<��<�<�J	<�<v�<{��;U��;�i�;BZ�;�[�;Cn�;��;���;_�;w�;��;S{�;h �;{ޤ;��;���;x��;�ی;_�;~�;��w;3m;+�b;X;��M;I�C;�%:;��0;�0';� ;l;�3;Z�;0C�:���:u��:���:�
�:���:K:m�:3u:��X:�t<:�� :�x:G
�9Rǟ9gKV9�P�8�q�6&����C��ܓ�YgŹ�x��V����+���C�3a[��r��6���ߐ�tz��|��v�������tʺ��պ�@���������#F���!�������cH#�k�(��e.���3�ry9�
?�_�D�J���O�U�c�Z�,3`���e�'Lk��p�iv���{�wÀ�;���aR�������������zn���5�������ř��  �  ǎ=|5=
�=d�=�(=g�=t=}=�� =�c =� =qZ�<l��<��<p4�<q|�<��<8�<�Q�<��<���<*"�<f�<��<��<,�<�k�<���<o��<�$�<H`�<l��<j��<:�<�A�<�v�<���<���<,�<�;�<�h�<	��<&��<���<��<�#�<U@�<�Y�<"p�<͂�<ב�<ۜ�<���<��<���<��<j��<��<�q�<�W�<v8�<p�<3��<¶�<�~�<�@�<Z��<c��<f\�<��<ҡ�<:�<���<xV�<���<�X�<
��<_A�<���<+�<�q�<7̸<� �<�p�< ��<~ �<TA�<{}�<M��<�<��<�D�<�m�<�<z��<F՟<��<�<[&�<9=�<IR�<�e�<iw�<���<y��<���<,��<(��<ņ<�̈́<�Ղ<.݀<��}<��y<!�u</�q<<�m<l j<�f<0b<6%^<3Z<9BV<�RR<dN<wJ<f�F<g�B<�><��:<L�6<@3<�,/<WP+<�v'<-�#<n�< <Q9<�u<j�<��<lL	<K�<��<߸�;��;�j�;[�;�[�;,n�;;��;���;��;�t�;E�;=x�;N�;Zۤ;���;k��;��;�،;�;q{�;@�w;�m;d}b;�X;<�M;)�C;�&:;��0;b3';�;�;9;�;�P�:;��:��:���:C�:�Ϧ:w͗:��:h#u:��X:T<:\� :�{:��95��9{!V9���8���6�E��D������Ź�������s�+�g�C��{[��s��@��P鐺+������������tʺ��պ�<���\�������@�3��,~���Y��UA#���(�_.���3�t9�0�>�݄D��J��O��U�ߨZ�j4`�}�e�)Ok�#�p��mv���{��ƀ������U��E��1䋻�����q���8�������Ǚ��  �  ��=P5=��=[�=�(=~�=;t=�=�� =d =� =+[�<8��<���<75�<2}�<���<��<�R�<���<���<�"�<`f�<7��<��<�+�<�k�<V��<���<[$�<�_�<���<���<d
�<�@�<v�<���<���<x�<9;�<�g�<��<���<s��<v�<t#�<x@�<-Z�<�p�<<��<H��<���<���<���<|��<���<0��<ۆ�<Ur�<�X�<!9�<��<���<%��<.�<�@�<I��<5��<&\�<�<=��<�9�<���<�U�<���<�W�<4��<�@�<׫�<k�<1q�<�˸<c �<p�<���<I �<,A�<q}�<m��<C�<)�<HE�<n�<���<-��<�՟<J�<D�<'�<>�<S�<Wf�<x�<+��<�<S��<_��<@��<ņ<�̈́<�Ղ<�܀<b�}<��y<��u<��q<��m<��i<q
f<~b<�#^<�1Z<�@V<_QR<�bN<vJ<��F<"�B<�><��:<��6<�3<�-/<7Q+</x'<��#<��<�<�:<Dw<��<~ <�M	<ġ<)�<���;��;2l�;�[�;:\�;n�;ڑ�;.��;�;�r�;�;�u�;��;2ؤ;���;���;Э�;֌;x�;�x�;X�w;�m;%zb;�X;L�M;�C;�':;ӕ0;�6';�;�;�>;��;�\�:���:���:7��:I%�:ۦ:�ؗ:��:a2u:[�X:��<:�� :؀:��9l��94V9U��8�x�6zɾ�:oD��@��n�ŹC�������+�n�C���[��(s��J�������'����������tʺ��պX8���캣���D��K;�t��Fx�����3;#�1�(�HY.���3�o9���>�+�D��	J���O��U�b�Z�l5`��e�Sk���p�=rv�|��ɀ�����[Y��E ���狻����t��e;��/��ʙ��  �  c�=;5=��=P�=�(=��=Vt=�=1� =Jd =5	 =�[�<��<���<�5�<�}�<z��<��<%S�<��<^��<�"�<�f�<V��</��<�+�<�k�<)��<���<�#�<_�<*��<��<�	�<+@�<Hu�<	��<<��<��<�:�<|g�<%��<z��<J��<A�<x#�<�@�<SZ�<�p�<���<���<��<Y��<^��<7��<`��<��<���<�r�<+Y�<�9�<T�<���<a��<N�<�@�<N��<���<�[�<��<ݠ�<	9�<U��<U�<1��<�V�<b��<�?�<��<��<�p�<�ʸ<��<�o�<O��< �<�@�<�}�<���<e�<b�<�E�<�n�<%��<Ѷ�<�֟<��<��<�'�<�>�<�S�<�f�<�x�<���<E��<���<���<`��<�Ć<�̈́<sՂ<r܀<��}<p�y<��u<}�q<8�m<V�i<�f<b<$"^<_0Z<�?V<5PR<+bN<zuJ<T�F<��B<Ÿ><��:<��6<S3<E./<'R+<,y'<ϣ#<F�<<v<<�x<��<�<VO	<��<6�<���;R��;m�;�\�;�\�;�m�;:��;���;�;�q�;��;�s�;�;�դ;�;���;F��;=ӌ;&�;�v�;��w;�m;�xb;�X;��M;U�C;�(:;3�0;�8';�;�;�B;�;g�:���:9��:���:l1�:��:��:B"�:�Au:��X:�<:z� :s�:V	�9F��9 �U9I�8��6]?��A�D��f����Ź���T��K�+���C���[�%;s��T��l���z���I��v���a	�� sʺ��պ�5�Ќ�����p��7�4���r���~��<5#���(�T.���3�'k9���>��~D�J�}�O��U���Z�7`�S�e�Uk���p��vv��|�3̀�{���\��}#��Eꋻ����9w���=��u���˙��  �  <�=5=��=L�=�(=��=wt=�=g� ={d =g	 =H\�<Z��<+��<s6�<}~�<���<	�<�S�<���<���<"#�<�f�<h��<)��<�+�<ik�<��<K��<�#�<�^�<���<���<=	�<�?�<�t�<���<���<r�<5:�<g�<ґ�<-��<��<2�<t#�<�@�<�Z�<q�<��<4��<^��<���<ը�<���<��<n��<��<ms�<�Y�<�9�<��<C��<���<��<�@�<B��<��<�[�<��<���<�8�<���<�T�<���<vV�<���<.?�<���<�< p�<kʸ<{�<Jo�<��<���<�@�<q}�<���<��<��<F�<�n�<|��<9��<ן<���<��<d(�<+?�<#T�<Zg�<�x�<��<���<Ѥ�<���<[��<�Ć<�̈́<4Ղ<"܀<��}<��y<��u<��q<3�m<j�i<�f<"b<#!^<l/Z<�>V<UOR<saN<�tJ<щF<h�B<��><��:<*�6<�3<�./< S+<�y'<��#<7�<�<�=<�y<��<�<AP	<��<�<Z��;}��;@n�;]�;�\�;�m�;���;���;��;!p�;>�;r�;<�;�Ӥ;	��;c��;���;Jь;��;u�;k�w;�m;Fvb;�X;��M;^�C;�(:;ޘ0;�:';;D;�E;@�;�n�:���:��:���:�8�:3�:�:�'�:6Pu:�X:�<:�� :D�:��9���9��U9P �8#��6���	�D�g���zƹ).������,���C��[��Gs�M[�������������z����	���sʺ*�պ�1ẵ��������%4����Ro���!���0#���(�PP.���3�3h9�r�>��|D�J�K�O�U��Z�8`�T�e��Wk�I�p�zv�|��̀�����]���%��+싻����y��a?��+��͙��  �  ,�=
5=��=I�=�(=��=�t==o� =�d =�	 =�\�<���<x��<�6�<�~�<T��<g�<�S�<���<���<N#�<�f�<���<"��<�+�<]k�<ɩ�<$��<X#�<v^�<d��<1��<��<F?�<jt�<(��<d��<�<�9�<�f�<���<��<���<4�<f#�<�@�<�Z�<#q�<��<H��<���<��<?��<���<C��<ʗ�<Y��<�s�<�Y�<M:�<��<_��<���<��<�@�<0��<��<�[�<j�<L��<X8�<���<;T�<H��<�U�<t��<�>�<'��<��<�o�<1ʸ<=�<o�<๳<���<�@�<`}�<���<��<��<F�<o�<Ք�<���<~ן<���<��<�(�<�?�<�T�<�g�<6y�<'��<���<뤌<���<e��<�Ć<�̈́<Ղ<܀<��}<4�y<&�u<��q<y�m<��i<f<Ob<[ ^<�.Z< >V<�NR<�`N<�tJ<��F<\�B<��><��:<L�6<3<%//<!S+<{z'<L�#<�<�<7><�z<Q�<�<Q	<{�<��<���;@��;�n�;�]�;�\�;�m�;���;]��;_�;To�;��;�p�;��;8Ҥ;���;A��;�;
Ќ;*�;t�;��w;m;�ub;X;��M;�C;�):;{�0;�;';>;�;gH;�;yu�:(��:ö�:���:�=�:��:{�:�-�:�Su:��X:C�<:�� :]�:��9��9��U9���8���6�⿸�E����2/ƹ�J����e,��D���[�Ts��^��t��h���C������
��Xtʺ��պ�0��캒������G1����l�D�!��c.#�
�(� M.�4�3��e9���>�9{D�RJ���O��U�7�Z�8`�T�e�~Xk�$�p��{v��|�gπ�𗃻�_���&���틻~����z���@������͙��  �  )�=5=��=F�=�(=��=t=2=� =�d =�	 =�\�<ͥ�<���<�6�<�~�<j��<d�<�S�<Й�<��<|#�<�f�<���<0��<�+�<Hk�<���<��<;#�<`^�<E��<6��<��<+?�<[t�<��<g��<�
�<�9�<�f�<{��<	��<���<%�<e#�<�@�<�Z�<7q�<C��<b��<՞�<��<C��<	��<X��<��<h��<�s�<�Y�<l:�<��<���<Է�<y�<�@�<2��<׮�<w[�<[�<,��<<8�<���<T�<P��<�U�<`��<�>�<��<��<�o�<ʸ< �<o�<ѹ�<���<�@�<h}�<���<��<��<JF�</o�<唣<���<�ן<���< �<�(�<�?�<�T�<�g�<Wy�<E��<�<奈<���<|��<�Ć<v̈́<Ղ< ܀<G�}<�y<��u<��q<q�m<F�i<�f<b<L ^<�.Z<�=V<�NR<�`N<�tJ<g�F<;�B<��><�:<K�6<�3<�//<eS+<�z'<R�#<�<�<X><�z<z�<�<Q	<��<��<s��;��;an�;�]�;]�;�m�;K��;+��;8�;�n�;<�;6p�;�;�Ѥ;(��;
��;f��;Ќ;��;�s�;�w;�m;Hub;qX;C�M;�C;�*:;�0;�<';?;�;zI;֪;�u�:��: ��:��:�>�:���:?�:~/�:�Vu:z�X:��<:E� :��:F�9t��9w�U9���8��6����E�d����,ƹ�R��F��M,��	D�F�[�Xs�`����������󙳺���sʺl�պ�1ẝ��~������0���ck������-#���(�3M.�?�3��d9��>�QyD�2J��O�U�U�Z��8`���e��Xk��p�4|v��|��π�����&`��&'��L�����z��9A��5��{Ι��  �  ,�=
5=��=I�=�(=��=�t==o� =�d =�	 =�\�<���<x��<�6�<�~�<T��<g�<�S�<���<���<N#�<�f�<���<"��<�+�<]k�<ɩ�<$��<X#�<v^�<d��<1��<��<F?�<jt�<(��<d��<�<�9�<�f�<���<��<���<4�<f#�<�@�<�Z�<#q�<��<H��<���<��<?��<���<C��<ʗ�<Y��<�s�<�Y�<M:�<��<_��<���<��<�@�<0��<��<�[�<j�<L��<X8�<���<;T�<H��<�U�<t��<�>�<'��<��<�o�<1ʸ<=�<o�<๳<���<�@�<`}�<���<��<��<F�<o�<Ք�<���<~ן<���<��<�(�<�?�<�T�<�g�<6y�<'��<���<뤌<���<e��<�Ć<�̈́<Ղ<܀<��}<4�y<&�u<��q<y�m<��i<f<Ob<[ ^<�.Z< >V<�NR<�`N<�tJ<��F<\�B<��><��:<L�6<3<&//<!S+<{z'<L�#<�<�<7><�z<Q�<�<Q	<{�<��<���;@��;�n�;�]�;�\�;�m�;���;]��;_�;So�;��;�p�;��;8Ҥ;���;A��;�;	Ќ;*�;t�;��w;m;�ub;X;��M;�C;�):;{�0;�;';>;�;gH;�;yu�:'��:ö�:���:�=�:��:{�:�-�:�Su:��X:C�<:�� :]�:��9��9��U9���8���6�⿸�E����2/ƹ�J����e,��D���[�Ts��^��t��h���C������
��Xtʺ��պ�0��캒������G1����l�D�!��c.#�
�(� M.�4�3��e9���>�9{D�RJ���O��U�7�Z�8`�T�e�~Xk�$�p��{v��|�gπ�𗃻�_���&���틻~����z���@������͙��  �  <�=5=��=L�=�(=��=wt=�=g� ={d =g	 =H\�<Z��<+��<s6�<}~�<���<	�<�S�<���<���<"#�<�f�<h��<)��<�+�<ik�<��<K��<�#�<�^�<���<���<=	�<�?�<�t�<���<���<r�<5:�<g�<ґ�<-��<��<2�<t#�<�@�<�Z�<q�<��<4��<^��<���<ը�<���<��<n��<��<ms�<�Y�<�9�<��<C��<���<��<�@�<B��<��<�[�<��<���<�8�<���<�T�<���<vV�<���<.?�<���<�< p�<kʸ<{�<Jo�<��<���<�@�<q}�<���<��<��<F�<�n�<|��<9��<ן<���<��<d(�<+?�<#T�<Zg�<�x�<��<���<Ѥ�<���<[��<�Ć<�̈́<4Ղ<"܀<��}<��y<��u<��q<3�m<j�i<�f<"b<#!^<l/Z<�>V<UOR<saN<�tJ<щF<h�B<��><��:<*�6<�3<�./< S+<�y'<��#<7�<�<�=<�y<��<�<AP	<��<�<Z��;}��;@n�;]�;�\�;�m�;���;���;��;!p�;>�;r�;<�;�Ӥ;	��;c��;���;Jь;��;u�;k�w;�m;Fvb;�X;��M;^�C;�(:;ޘ0;�:';;D;�E;@�;�n�:���:��:���:�8�:3�:�:�'�:6Pu:�X:�<:�� :D�:��9���9��U9P �8#��6���	�D�g���zƹ).������,���C��[��Gs�M[�������������z����	���sʺ*�պ�1ẵ��������%4����Ro���!���0#���(�PP.���3�3h9�r�>��|D�J�K�O�U��Z�8`�T�e��Wk�I�p�zv�|��̀�����]���%��+싻����y��a?��+��͙��  �  c�=;5=��=P�=�(=��=Vt=�=1� =Jd =5	 =�[�<��<���<�5�<�}�<z��<��<%S�<��<^��<�"�<�f�<V��</��<�+�<�k�<)��<���<�#�<_�<*��<��<�	�<+@�<Hu�<	��<<��<��<�:�<|g�<%��<z��<J��<A�<x#�<�@�<SZ�<�p�<���<���<��<Y��<^��<7��<`��<��<���<�r�<+Y�<�9�<T�<���<a��<N�<�@�<N��<���<�[�<��<ݠ�<	9�<U��<U�<1��<�V�<b��<�?�<��<��<�p�<�ʸ<��<�o�<O��< �<�@�<�}�<���<e�<b�<�E�<�n�<%��<Ѷ�<�֟<��<��<�'�<�>�<�S�<�f�<�x�<���<E��<���<���<`��<�Ć<�̈́<sՂ<r܀<��}<p�y<��u<}�q<8�m<V�i<�f<b<$"^<_0Z<�?V<5PR<+bN<zuJ<T�F<��B<Ÿ><��:<��6<S3<E./<'R+<,y'<ϣ#<F�<<w<<�x<��<�<UO	<��<6�<���;R��;m�;�\�;�\�;�m�;:��;���;�;�q�;��;�s�;�;�դ;�;���;F��;=ӌ;&�;�v�;��w;�m;�xb;�X;��M;U�C;�(:;3�0;�8';�;�;�B;�;g�:���:9��:���:l1�:��:��:B"�:�Au:��X:�<:z� :s�:V	�9F��9 �U9I�8��6]?��A�D��f����Ź���T��K�+���C���[�%;s��T��l���z���I��v���a	�� sʺ��պ�5�Ќ�����p��7�4���r���~��<5#���(�T.���3�'k9���>��~D�J�}�O��U���Z�7`�S�e�Uk���p��vv��|�3̀�{���\��}#��Eꋻ����9w���=��u���˙��  �  ��=P5=��=[�=�(=~�=;t=�=�� =d =� =+[�<8��<���<75�<2}�<���<��<�R�<���<���<�"�<`f�<7��<��<�+�<�k�<V��<���<[$�<�_�<���<���<d
�<�@�<v�<���<���<x�<9;�<�g�<��<���<s��<v�<t#�<x@�<-Z�<�p�<<��<H��<���<���<���<|��<���<0��<ۆ�<Ur�<�X�<!9�<��<���<%��<.�<�@�<I��<5��<&\�<�<=��<�9�<���<�U�<���<�W�<4��<�@�<׫�<k�<1q�<�˸<c �<p�<���<I �<,A�<q}�<m��<C�<)�<HE�<n�<���<-��<�՟<J�<D�<'�<>�<S�<Wf�<x�<+��<�<S��<_��<@��<ņ<�̈́<�Ղ<�܀<b�}<��y<��u<��q<��m<��i<p
f<~b<�#^<�1Z<�@V<_QR<�bN<vJ<��F<"�B<�><��:<��6<�3<�-/<7Q+</x'<��#<��<�<�:<Dw<��<~ <�M	<ġ<)�<���;��;2l�;�[�;:\�;n�;ڑ�;-��;�;�r�;�;�u�;��;2ؤ;���;���;Э�;֌;x�;�x�;X�w;�m;%zb;�X;K�M;�C;�':;ӕ0;�6';�;�;�>;��;�\�:���:���:7��:I%�:ۦ:�ؗ:��:a2u:[�X:��<:�� :؀:��9l��94V9U��8�x�6zɾ�:oD��@��n�ŹC�������+�n�C���[��(s��J�������'����������tʺ��պX8���캣���D��K;�t��Fx�����3;#�1�(�HY.���3�o9���>�+�D��	J���O��U�b�Z�l5`��e�Sk���p�=rv�|��ɀ�����[Y��E ���狻����t��e;��/��ʙ��  �  ǎ=|5=
�=d�=�(=g�=t=}=�� =�c =� =qZ�<l��<��<p4�<q|�<��<8�<�Q�<��<���<*"�<f�<��<��<,�<�k�<���<o��<�$�<H`�<l��<j��<:�<�A�<�v�<���<���<,�<�;�<�h�<	��<&��<���<��<�#�<U@�<�Y�<"p�<͂�<ב�<ۜ�<���<��<���<��<j��<��<�q�<�W�<v8�<p�<3��<¶�<�~�<�@�<Z��<c��<f\�<��<ҡ�<:�<���<yV�<���<�X�<
��<_A�<���<+�<�q�<7̸<� �<�p�< ��<~ �<TA�<{}�<M��<�<��<�D�<�m�<�<{��<F՟<��<�<[&�<9=�<IR�<�e�<iw�<���<y��<���<,��<(��<ņ<�̈́<�Ղ<.݀<��}<��y<!�u</�q<<�m<l j<�f<0b<6%^<3Z<9BV<�RR<dN<wJ<f�F<g�B<�><��:<L�6<@3<�,/<WP+<�v'<-�#<n�< <Q9<�u<j�<��<kL	<K�<��<߸�;��;�j�;[�;�[�;,n�;;��;���;��;�t�;E�;=x�;N�;Zۤ;���;k��;��;�،;�;q{�;@�w;�m;d}b;�X;;�M;)�C;�&:;��0;b3';�;�;9;�;�P�:;��:��:���:C�:�Ϧ:w͗:��:h#u:��X:T<:\� :�{:��95��9{!V9���8���6�E��D������Ź�������s�+�g�C��{[��s��@��P鐺+������������tʺ��պ�<���\�������@�3��,~���Y��UA#���(�_.���3�t9�0�>�݄D��J��O��U�ߨZ�j4`�}�e�)Ok�#�p��mv���{��ƀ������U��E��1䋻�����q���8�������Ǚ��  �  ��=�5=!�=l�=|(=N�=�s=G=t� =fc =; =�Y�<���<<��<�3�<�{�<.��<y
�<=Q�<]��<���<�!�<�e�<��<��<$,�<,l�<��<���<z%�<�`�<?��<=��<�<�B�<�w�<u��<���<�<�<�<i�<���<���<��<��<�#�<A@�<�Y�<�o�<T��<.��<7��<R��<0��<ڤ�<��<���<?��<�p�<(W�<�7�<��<���<x��<�~�<s@�<o��<���<�\�<�<W��<�:�<n��<cW�<���<�Y�<���<SB�<���<�<�r�<�̸<�!�<q�<s��<� �<uA�<�}�<8��<��<j�<gD�<�l�<S��<Ĵ�<lԟ<��<��<{%�<`<�<|Q�<�d�<�v�<��<��<���<���<��<ņ<΄<Gւ<�݀<��}<��y<��u<��q<��m<=j<�f<b<�&^<�4Z<�CV<�SR<7eN<�wJ<)�F<ȡB<C�><��:<��6<�3<�+/<)O+<�u'<џ#<��<> <�7<�s<��<�<�J	<�<v�<{��;T��;�i�;BZ�;�[�;Cn�;��;���;^�;w�;��;S{�;h �;zޤ;��;���;w��;�ی;_�;~�;��w;3m;+�b;X;��M;I�C;�%:;��0;�0';� ;l;�3;Z�;0C�:���:u��:���:�
�:���:K:m�:3u:��X:�t<:�� :�x:G
�9Rǟ9gKV9�P�8�q�6&����C��ܓ�YgŹ�x��V����+���C�3a[��r��6���ߐ�tz��|��v�������tʺ��պ�@���������#F���!�������cH#�k�(��e.���3�ry9�
?�_�D�J���O�U�c�Z�,3`���e�'Lk��p�iv���{�wÀ�;���aR�������������zn���5�������ř��  �  -�=�5=:�=p�=s(=5�=�s==/� =c =� =�X�<���<V��<�2�<�z�<[��<�	�<}P�<Ŗ�<u��<d!�<|e�<���<���<5,�<bl�<f��<I��<&�<�a�<��<��<��<wC�<�x�<K��<g��<��<<=�<�i�<��<��<J��<��<�#�<.@�<sY�<qo�<��<���<���<~��<]��<��<%��<���<j��<�o�<RV�<47�<1�<M��<��<~~�<f@�<p��<���<]�<e�<��<�;�<"��<&X�<���<gZ�<���<FC�<���<��<�s�<�͸<W"�<�q�<ϻ�<�<�A�<�}�<&��<��<�<�C�<Vl�<���<ﳡ<�ӟ<��<��<�$�<�;�<�P�<%d�<v�<���<���<H��<���<��< ņ<E΄<�ւ<�݀<��}<3�y<��u<h�q<��m<�j<�f<�b<�(^<i6Z<1EV<)UR<ffN<�xJ<��F<3�B<Z�><r�:<��6<�
3<+/<N+<Mt'<.�#<�<��<�5<�q<ų<Y�<I	<K�<-�<A��;���;�g�;uY�;5[�;Nn�;���;���;��;Zy�;�;�}�;y#�;��;m��;#��;���;Cߌ;"�;���;��w;!m;͂b;�X;��M;��C;�$:;]�0;l-';b�;z�;~.;��;�5�:+��:'s�:��:��:9��:���:���:��t:�zX:Yh<:� :�u:��9I͟9�jV9���8}�6����rC�	���W0Ź�B��rt���+��C�]F[�6�r�:,��gՐ��r������������yuʺv�պ"F�������צ��K����ԋ��%�����O#��(�$l.�n�3�s~9��?���D�J���O��U�8�Z��1`���e��Hk���p��cv�V�{�s���ȇ���N����(݋�B���ek���2������qÙ��  �  h�=�5=P�=w�=i(=%�=�s=�=� =�b =~ = X�<��<���<�1�<�y�<���<��<�O�<;��<���<� �<.e�<���<���<O,�<�l�<ë�<���<�&�<9b�<���<���<��<=D�<cy�<��<!��<x�<�=�<Sj�<x��<V��<���<�<�#�<@�<JY�<o�<b��<��<��<͡�<���<.��<]��<��<���<Mo�<�U�<�6�<��<���<���<V~�<M@�<t��<߯�<W]�<��<^��<<�<���<�X�<P��<A[�<���<D�<k��<��<Yt�<Zθ<�"�<r�<=��<]�<�A�<�}�<��<K�<��<lC�<�k�< ��<A��<�ҟ<��<�
�<�#�<�:�<�O�<vc�<�u�<���<��<䢌<���<꺈<'ņ<p΄<�ւ<gހ<}�}<^�y<^�u<��q<1�m<j<)f<Pb<<*^<�7Z<�FV<iVR<IgN<�yJ<d�F<��B<y�><O�:<G�6<>
3<*/<�L+<'s'<˜#<��<��<�3<_p<�<��<�G	<��<�<ձ�;���;�f�;�X�;�Z�;�n�;/��;��;��;�z�;l�;r��;3&�;��;X��;��;���;�;�$�;2��;��w;/$m;�b;�X;��M;��C;�#:;ݍ0;*';�;'�;H);Շ;V*�:G��:Lf�:V��:�:��:*��:4�:�t:�iX:[<:� :zq:@�9�ן9�V9��8�E�6�}��cC������ŹE��C[��z+��iC�l/[�m�r��!��Hΐ��k����������� ��Fvʺ��պrJ�@�캃��
��%Q��������,����V#���(��q.���3�"�9�
?���D�J���O�K U���Z�l0`�+�e�OEk�/�p��^v���{����������K����ڋ����h��!0��`��������  �  ��=6=`�=��=](=	�={s=�=�� =�b =4 =yW�<;��<���<1�<+y�<���<K�<7O�<���<���<� �<e�<h��<���<m,�<�l�<��<��<'�<�b�<@��<o��<l�<�D�<z�<ԭ�<���< �<w>�<�j�<��<���<���<"�<�#�<�?�<Y�<�n�<��<���<V��<;��<���<��<���<(��<��<�n�<U�<�5�<F�<��<���<2~�<%@�<���<��<�]�<*�<̣�<�<�<q��<�Y�<��<\�<���<�D�<3��<p�<u�<�θ<^#�<}r�<���<��<�A�<�}�<ߴ�<+�<u�<C�<Yk�<j��<���<,ҟ<T�<6
�<#�<:�<HO�<�b�<�t�<���<͔�<���<[��<ʺ�<@ņ<�΄<ׂ<�ހ<^�}<W�y<��u<1�q<��m<j<�f<�b<�+^<=9Z<�GV<gWR<9hN<KzJ<ӍF<٢B<��>< �:<��6<�	3<�)/< L+<�q'<��#<U�<o�<�2<�n<��<:�<<F	<��<��<8��;\��;�e�;�W�;�Z�;�n�;���;���;��;�|�;7��;ɂ�;�(�;k�;!��;ɰ�;{��;��;Q'�;+��;l�w;A'm;�b;�X;u�M;B�C;E":;M�0;C(';`�;��;E$;�;��:��:MZ�:w�:��:v��:П�:Z�:��t:#_X:�S<:�� :vk:�
�98ߟ9A�V9�U�8�y�6���,�B�	X����Ĺ����wD�tc+�YRC��[�Ͷr�����Ɛ�=f������H�������7vʺ"�պ M���'
��/���U�r�����2�����[#�K�(�$w.�p 4���9�9?� �D��J�c�O�A!U�#�Z�}/`���e�1Ck���p�[v�:�{�캀������H��?��׋�Z����e���-��t���꿙��  �  ��=16=p�=��=X(=��=[s=�=�� =Ob =� = W�<���<V��<�0�<�x�<]��<��<�N�<C��<3��<] �<�d�<N��<���<f,�<�l�<@��<W��<t'�<c�<���<���<��<�E�<�z�<T��<@��<��<�>�<:k�<>��<ټ�<���<*�<�#�<�?�<�X�<�n�<���<=��<��<נ�<u��<��<��<���<x��<n�<�T�<�5�<��<0��<D��< ~�<!@�<���<��<�]�<q�<*��<
=�<���<Z�<���<�\�<��<vE�<���<��<yu�<Kϸ<�#�<�r�<Ѽ�<��<�A�<�}�<մ�<��<,�<�B�<�j�<��<A��<�џ<��<�	�<�"�<�9�<�N�<yb�<|t�<3��<z��<v��<2��<���<:ņ<�΄<Cׂ<�ހ<*�}<!�y<F�u<�q<u�m<!j<�f<�b<�,^<(:Z<�HV<3XR<iN<�zJ<]�F<�B<��><�:<��6<k	3<�(/<hK+<q'<Ě#<\�<m�<�1<�m<��<+�<SE	<��<��<���;���;�d�;-W�;KZ�;�n�;��;���;��;F~�;���;<��;d*�;�;,��;ܲ�;[��;?�;�(�;|��;� x;�)m;ǉb;� X;��M;��C;�!:;��0;�%';��;B�;� ;�;L�:��:�Q�:Hn�:ݵ:ٔ�:X��:�ވ:"�t:�TX:�J<:�� :$j:��9Fߟ9�V9���8���6����T�B�:>���Ĺ�����2�CR+�+DC��[�R�r����a����a������]~��C���qvʺ;�պ�P���n�����<Y��������5�����_#���(�{.��4�\�9�2?���D�zJ���O��!U�C�Z��.`���e�Ak�x�p��Wv�>�{�-���2����F�����ԋ�����d��;,������B����  �  ď=;6=y�=��=V(=��=Js=x=i� =8b =� =�V�<Z��<���<?0�<Jx�<��<�<�N�<��<���<A �<�d�<M��<���<r,�<�l�<Z��<���<�'�<bc�<���<N��<;�<�E�<{�<���<���<��<.?�<ak�<W��<��<��<B�<�#�<�?�<�X�<yn�<���<��<���<u��<"��<���<ƛ�<N��<��<�m�<NT�<[5�<��<��<0��<�}�<%@�<���<+��<�]�<��<L��<.=�<4��<mZ�<���<�\�<���<�E�<��<b�<�u�<�ϸ<�#�<�r�<���<��<B�<�}�<۴�<��<�<�B�<�j�<���<㱡<Xџ<w�<Z	�<3"�<%9�<rN�<b�<Kt�<���<T��<T��<'��<���<5ņ<�΄<Rׂ<߀<O�}<��y<��u<��q<B�m<�j<mf<� b<R-^<�:Z<KIV<�XR<7iN<4{J<��F<C�B<��><�:<��6<'	3<�(/<�J+<�p'<�#<��<��<�0<�l<®<p�<�D	<�<��<���;x��;d�;W�;Z�;�n�;K��;��;4�;u~�;���;x��;�+�;t�;j;E��;w��;��;=*�;߇�;�x;�*m;�b;� X;8�M;a�C;�!:;�0;%';3�;l�; ;�|;��:΂�:>L�: i�:�յ:���:��:�ڈ:�t:�NX:�G<:s� :7j:�9{�9��V9���8�R 7Ru���|B�^(���Ĺd���&'��F+�&9C�|�Z�ɟr����?���b_����G}�����Ewʺ�պ�Rẅ�����)���[����I��9�����b#�U�(��}.��4��9�?���D��J��O��!U�h�Z�.`��e��?k���p�;Vv���{������~���E������Ӌ�
����b���*���� ����  �  K�=;3=�=�~=$=N�=@n=
=�� =�[ =)  =~H�<D��<���<��<�e�<��<��<�7�<�|�<���<[�<G�<���<���<�	�<XH�<��<q��<���<�7�<-p�<���<h��<��<�D�<&v�<Υ�<���<W��<)�<hP�<bu�<���<S��<���<���<��<��<o&�<U2�<�:�<�>�<�>�<�:�<Y2�<Z%�<��<��<��<��<��<gl�<�9�<�<��<o|�<t0�<���<U��<F$�<���<BP�<d��<:b�<���<�Z�<ξ<V;�<ࢻ<��<a�<��<
�<�V�<���<9�<!�<�[�<H��<Ũ<1��< �<�H�<�n�<���<;��<�Л<��<5�<��<r6�<�K�<h_�<�q�<͂�<���< ��<���<1��<�Ƃ<�р<��}<�y<��u<n�q<$n<�j<�$f<�6b<`I^<�\Z<:qV<ÆR<<�N<7�J<Z�F<��B<F?<�$;<
F7<[i3<��/<��+<��'<�$<�J <��<K�<@<�L<h�<��	<�J<��<*�;S
�;K��;���;_�;d(�;�Z�;���;���;�e�;q�;ǀ�;R0�;Q��;�֠;�Ϛ;�;�;�R�;��;�[|;�q;��f;�v\;5?R;�8H;hf>;z�4;V+;�";�;�';�t;���:�)�:���:��:%��:!��:V�:;l�:x��:C�d:�4H:@/,:+�:���9m��9��~9�9��58F�f�s��Ez��'���O7���#$��`<��nT��Wl�a��ݍ�����hR������땼��*Ⱥ��Ӻ�5ߺ��꺙!��4� �Cv�
#�Q���p�}�3�"�<G(�3�-�Zq3��9��>�}D�'�I�9:O�7�T�GVZ���_��ue�Nk�C�p�,)v�̼{�K���>r���<������ы�}����g���3��0 ��Ι��  �  <�=C3=�=�~=$=K�=Bn==�� =\ =7  =�H�<E��<���<��<�e�<��<!��<�7�<�|�<���<e�<G�<��<���<�	�<aH�<���<L��<���<z7�< p�<p��<[��<��<�D�<v�<���<{��<D��<�(�<?P�<Eu�<���<J��<���<���<��<��<�&�<o2�<�:�<�>�<�>�<�:�<r2�<q%�<��<���<#��<��<#��<�l�<�9�<�<
��<r|�<i0�<���<;��<$�<v��<,P�<[��< b�<���<�Z�<ξ<I;�<ɢ�<��<�`�<��<�	�<�V�<͞�<2�<
!�<�[�<J��< Ũ<M��<' �<�H�<�n�<���<Y��<�Л<��<;�<��<�6�<�K�<�_�<�q�<т�<���<(��<���<0��<�Ƃ<�р<p�}<��y<b�u<]�q< n<�j<V$f<�6b<CI^<�\Z<qV<��R<�N<��J<{�F<��B<B?<�$;<�E7<bi3<��/<��+<��'<$<�J <��<��<�<M<e�<��	<�J<��<�*�;
�;Z��;h��;��;V(�;�Z�;���;M��;�e�;�;���;0�; ��;�֠;�Κ;���;��;�R�;Ҳ�;[|;��q;�f;�w\;�>R;�8H;tf>;��4;gV+;�";�;?(;}u;{��:�*�:H��:`��:���:���:�W�: m�:
:��d:�6H:�/,:k�:���9���9�~99�9058g����(|�����c:���i&$��a<��qT�VYl����zލ�=����R�����H���2*Ⱥ��Ӻ�5ߺ�����z� ��u�n"�j���o���@�"�G(��-�|p3�K9��>�*D��I�`:O���T�2VZ���_��te�(k�3�p�*v�H�{�m����r���<��<���ы�����h���3��� ��nΙ��  �  /�=83=�=�~= $=T�=Tn==�� =\ =S  =�H�<���<��<�<f�<Y��<b��<�7�<�|�<���<y�<8G�<���<���<�	�<BH�<߅�<6��<w��<D7�<�o�<(��<��<��<|D�<�u�<o��<I��<
��<�(�<7P�<*u�<���<(��<���<���<�<�<�&�<�2�<�:�<?�<#?�<$;�<�2�<�%�<��<7��<g��<��<E��<�l�<�9�<3�<��<�|�<H0�<���<��<$�<]��<�O�<&��<�a�<Q��<�Z�<�;<;�<x��<g�<�`�<ﷶ<�	�<�V�<���<�<!�<�[�<l��<0Ũ<f��<G �<�H�<�n�<鑟<���<�Л<<�<��<��<�6�<�K�<�_�<�q�<�<���<4��<���<��<�Ƃ<xр<`�}<��y<��u<��q<r n<"j<�#f<6b<�H^<=\Z<�pV<)�R<�N<ĴJ<M�F<9�B<-?<%;< F7<�i3<��/<E�+<��'<�$<#K <�<�<�<�M<�<��	<QK<��<#+�;�
�;��;���;��;(�;UZ�;���;��;ge�;D�;��;�.�;+��;�ՠ;�͚;	��;��;�Q�;���;8Z|;{�q;W�f;	w\;�=R;Y9H;�f>;M�4;#W+;j";�	;o);�w;W��:�/�:6��:��:� �:���:�[�:Vo�:QĀ:ɧd:�8H:!3,:��:̍�9���9��~9�t9�58Eg����]���w����H�����.$��i<��zT��_l�I��]ߍ�T���T�����������(Ⱥ��Ӻ>3ߺ����k� �Lt�_ ����nm���0�"��D(��-��n3�@ 9���>�kD���I��9O���T�MVZ��_��ue��k�q�p�o+v��{�Z����s���=��^���ҋ�ʝ��
i���4��\���Ι��  �  �="3=�=�~=$=]�=gn=9=׷ =D\ =z  =I�<��<p��<��<bf�<¬�<���<"8�<}�<<��<��<XG�<��<���<�	�<5H�<���<��<��<�6�<�o�<Ԧ�<���<*�<D�<uu�<��<���<���<t(�<�O�< u�<o��<)��<���<���<!�<D�<�&�<�2�<;�<P?�<�?�<~;�<3�<&�<T�<���<���<j��<���<�l�<+:�<M�<��<x|�<B0�<j��<��<�#�<���<�O�<���<ta�<���<Z�<N;<�:�<��<�<j`�<���<�	�<uV�<���<�<!�<�[�<���<bŨ<���<� �<KI�<*o�<O��<���<Vћ<��<��<Y �<7�<NL�<�_�<4r�<��<���<3��<���<��<�Ƃ<Lр<Ŷ}<��y<P�u<1�q<��m<Kj<#f<35b<�G^<�[Z<	pV<��R<D�N<e�J<��F<3�B<*?<%;<EF7<�i3<_�/<չ+<��'<"$<�K <��<��<�<zN<Ŝ<8�	<L<��<M,�;��;���;��;��;7(�;;Z�;��;T��;d�; �;�~�;�-�;���;Ԡ;�̚;rޔ;M
�;�P�;Ű�;iW|;��q;*�f; v\;>R;f9H;�f>;Q�4;�X+;�";Y;L,;1z;k��:�5�:��:*��:=�::�`�: u�:wɀ:W�d:g?H:�6,:b�:��9n��9]�~99`9ן48%h�v! �����!���Pc����2;$�:v<���T��il�W��^卺�����V������ϗ��g)Ⱥ�Ӻe1ߺ�������� ��q���=���j�j��"��A(�B�-�/l3�s�8�_�>�oD���I�9O���T�WVZ���_��ve�dk�ޚp�.v���{������t��S?���	��iԋ�:���ij��6������ϙ��  �  ��=3=��=�~=%$=q�=|n=^=�� =u\ =�  =�I�<w��<���<  �<�f�<M��<6��<�8�<f}�<���<��<zG�<5��<���<�	�<H�<z��<���<���<�6�<o�<R��<4��<��<�C�<�t�<���<e��<\��<(�<�O�<�t�<C��<��<���<���<I�<|�<('�<)3�<v;�<�?�<@�< <�<�3�<�&�<��<'��<(��<���<ڙ�<m�<c:�<o�<,��<g|�<'0�<7��<���<v#�<���<6O�<8��<�`�<N��<�Y�<�̾<:�<���<��<`�<(��<8	�<4V�<h��<��<
!�<�[�<���<�Ũ<���<� �<�I�<�o�<ے�<w��<�ћ<�<i�<� �<�7�<�L�<@`�<�r�<L��<钊<J��<���<�<WƂ<р<�}<9�y<}�u<#�q<��m<6j<"f<4b<�F^<~ZZ<#oV<фR<��N<�J<��F<��B<?<,%;<�F7<Ij3<��/<b�+<u�'<$<�L <
�<��<<{O<�<E�	<M<l�<�-�;$�;J��;���;D�;(�;�Y�;:��;��;�b�;��;�|�;�+�;��;Ҡ;�ʚ;nܔ;w�;wN�;j��;�T|;I�q;��f;�t\;�=R;9H;
h>;��4;�Z+;�";�;�/;�};���:�=�:Y��:���:L�:'��:sh�:�{�:!΀:��d:GH:�;,:��:���9`��9ͤ~9�C9�48��h��L �����hڴ�7�湷���K$�C�<���T�,zl�x���ꍺ֨��oZ�����
���)Ⱥ��ӺE/ߺ ����9� ��m�������f����"��=(���-��h3�Q�8�8�>�D�F�I��7O���T��VZ���_��xe� 
k���p��0v���{�٬���v��yA������֋�)���wl���7�����?љ��  �  ό=�2=��=�~=,$=}�=�n=�=0� =�\ =�  =&J�<��<���<� �<g�<ۭ�<���<9�<�}�<���<D�<�G�<F��<���<p	�<�G�<@��<o��<i��<6�<�n�<Х�<���<�<�B�<Ut�<��<���<���<�'�<RO�<yt�<��<���<���<���<j�<��<�'�<�3�<�;�<H@�<�@�<�<�<14�<2'�<o�<���<���<O��<K��<~m�<�:�<��<9��<k|�<0�<��<[��<#�<��<�N�<���<W`�<���<�X�<̾<h9�<��<��<~_�<���<��<�U�<6��<��<!�<�[�<͒�<�Ũ<N��<O!�<6J�<p�<b��<��<wқ<��<	�<e!�<8�<(M�<�`�<�r�<���<��<[��<���<Ϻ�<'Ƃ<�Ѐ<v�}<I�y<r�u<�q<��m<�j<� f<�2b<�E^<sYZ<nV<ӃR<�N<8�J<�F<��B<�?<G%;<�F7<�j3<��/<>�+<[�'<'$<�M <>�<4�<;<�P<�<Z�	<N<[�<W/�;p�;Y��;/��;��;�'�;cY�;}��;L��;�a�;�;�z�;�)�;��;�Ϡ;EȚ;.ڔ;T�;�L�;t��;�Q|;�}q;S�f;�s\;�<R;�9H;�h>;��4;�\+; ";s;�3;2�;���:�G�:
��:A��:�:_��:�p�:���:�Հ:\�d:�OH:�@,:��:���9���9��~9�9T\38��i�"� ��߂�G���ª����k_$�љ<��T�g�l��#������\���@^�����Y���](Ⱥ��Ӻ�+ߺ��꺔���� ��i���u���a�B��"��8(���-�Ld3���8���>�sD�K�I� 7O��T��VZ��_�ze��k��p��4v���{�߮��Gy���C��W���؋�����n���9������ҙ��  �  ��=�2=��=�~=5$=��=�n=�=g� =�\ =A =�J�<���<<��<\!�<+h�<q��<R��<�9�<K~�<T��<��<�G�<c��<���<b	�<�G�<��<��<���<�5�<n�<-��<���<g�<PB�<�s�<\��<U��<T��<7'�<�N�<*t�<��<ζ�<���<���<��<�<�'�<4�<c<�<�@�<%A�<:=�<�4�<�'�<�<6��<=��<���<���<�m�<�:�<��<C��<f|�<�/�<���<
��<�"�<���<N�<��<�_�<���<2X�<i˾<�8�<O��<`�<�^�<B��<i�<�U�<��<��<	!�<�[�<��<ƨ<���<�!�<�J�<�p�<�<���< ӛ<g�<�	�<�!�<�8�<�M�<a�<s�<ԃ�<5��<m��<���<���<�ł<fЀ<��}<V�y<h�u<��q<;�m<�j<[f<�1b<qD^<6XZ<mV<ԂR<�N<z�J<��F<N�B<�?<e%;<G7<Sk3<�/<�+<I�'<M$<0O <|�<��<�	<5R<N�<��	<7O<[�<1�;��;���;���;��;�'�;�X�;���;���;�_�;.�; y�;�'�;(�;r͠;�Ś;�ה;��;wJ�;���;/N|;{q;�f;^r\;�;R;�9H;�i>;��4;_+;�"";�;j7;�;r�:R�:Z��:p��:�"�:���:jz�:{��:<܀:+�d:AXH:LH,:<�:h��9���9�y~9��9�28)sj�9� �|���(�����	��s$�]�<���T���l�(,������Z���Db��5��_����'Ⱥ�Ӻ�'ߺל꺋��&� ��e����h\������"��3(��-��_3��8�V�>�WD��I�{5O���T��VZ�B�_�{{e��k�K�p�L8v��{�:����{��RF����cۋ�.����p���;�����.ԙ��  �  ��=�2=��=�~=9$=��=�n=�=�� =&] =� =]K�<P��<���<
"�<�h�<��<���<&:�<�~�<���<��<(H�<���<���<R	�<�G�<���<���<���<(5�<m�<���<[��<��<�A�<s�<͢�<���<���<�&�<�N�<�s�<���<���<���<���<��<A�<3(�<v4�<�<�<gA�<�A�<�=�<�5�<�(�<��<���<���<C��<��<%n�<;�<��<X��<Z|�<�/�<���<���<H"�<,��<�M�<m��< _�<O��<wW�<�ʾ<	8�<���<��<k^�<˵�<�<OU�<���<��<!�<\�<0��<cƨ<��<,"�<4K�<Cq�<���<Y��<�ӛ<�<D
�<�"�<.9�<N�<�a�<}s�<��<`��<{��<���<���<�ł<)Ѐ<ٳ}<g�y<N�u<��q<
�m<cj<�f<E0b<9C^<�VZ<�kV<�R<-�N<��J<�F<��B<�?<u%;<fG7<�k3<ђ/<��+<J�'<[$<sP <ډ<��<<}S<��<��	<QP<`�<�2�;�;���;���;-	�;�'�;GX�;ɛ�;��;z^�;�߹;�v�;U%�;��;�ʠ;)Ú;`Ք;��;)H�;���;�J|;Kxq;V�f;�p\;O;R;�9H;Kj>;C�4;Ha+;�%";�;�;;s�;?�:�\�:���:���:-�:���:^��:瓏:Z�:��d:�`H:�M,:�:���9
��9(\~9��9��18QIk��!��)��M��1������$���<���T�_�l�f3��h�������f�����s����'Ⱥ��Ӻ�$ߺ���J��l� ��a�t���iW�x��Ĕ"��.(��-��[3�
�8��>�ID�S�I�/4O���T�YWZ�L�_��}e��k���p�<v�~�{�����Q~��I�����ދ�����Us��5>���	���ՙ��  �  [�=�2=��=�~==$=��=�n= =Ƹ =f] =� =�K�<��<s��<�"�<ai�<���<h��<�:�<9�<��<-�<VH�<���<���<A	�<wG�<���<p��<��<�4�<�l�<��<���<�<A�<kr�<D��<8��<O��<U&�<*N�<�s�<w��<���<���<��<��<��<�(�<�4�<n=�<�A�<QB�<o>�<6�< )�<B�<e �<C��<���<���<zn�<^;�<�<k��<H|�<�/�<W��<q��<�!�<���<M�<���<q^�<���<�V�<ʾ<b7�<��<*�<�]�<J��<��<U�<���<��<� �<4\�<Q��<�ƨ<Q��<�"�<�K�<�q�<(��<ﵝ<oԛ<��<�
�<!#�<�9�<�N�<�a�<�s�<H��<���<���<|��<x��<ył<�π<�}<��y<O�u<��q<��m<j<�f<�.b<B^<�UZ<�jV<��R<P�N<V�J<��F<��B<�?<�%;<�G7<&l3<��/<��+<M�'<m$<�Q <�<!�<c<�T<�<��	<kQ<\�<G4�;��;^��;O��;C	�;�'�;X�;���;���;�\�;�ݹ;�t�;m#�;��;�Ƞ;���;�Ҕ;���;@F�;���;�G|;Euq;R�f;8o\;�:R;�9H;!k>;��4;nc+;�(";�;@;��;��:�e�:��:��:�6�:>��:t��:��:3�:K�d:�iH:S,:#�:ي�9���9�F~9ɸ95#18�3l��O!�J���m���$��1��$��<�b�T�U�l�;����������j��	������O(Ⱥ��Ӻ5"ߺ������ܯ ��]������R�Q���"��)(���-�]W3���8�-~>��D���I��2O�,�T��WZ���_��e��k��p�x?v�w�{����������K���������㪎�au��C@��p���י��  �  6�=2=��=�~=F$=��=o==� =�] =� =bL�<d��<���<-#�<�i�<.��<���<;�<��<`��<e�<�H�<ɉ�<��<(	�<MG�<O��<%��<���<L4�<�l�<���<;��<��<�@�<�q�<���<���<���<&�<�M�<`s�<T��<���<���<��<�<��<�(�</5�<�=�<iB�<�B�<�>�<�6�<�)�<��<� �<���<��<՛�<�n�<�;�<1�<y��<H|�<|/�<)��<)��<�!�<Y��<�L�<`��<�]�<��<BV�<yɾ<�6�<���<� �<s]�<���<V�<�T�<f��<]�<� �<D\�<w��<�ƨ<���<�"�<L�<Fr�<���<w��<�ԛ<%�<Z�<�#�</:�<�N�<=b�<t�<~��<���<���<o��<Q��<Xł<�π<u�}<��y<^�u<��q<��m<!
j<�f<.b<�@^<�TZ<�iV<8�R<��N<��J<G�F<u�B<?<�%;<�G7<�l3<��/<N�+<��'<Y$<�R <�<<�<g<�U<��<	�	<GR<�<�5�;��;F �;���;�	�;s'�;�W�;X��;���;�[�;aܹ;)s�;`!�;��;�Ơ;ؾ�;є;v��;yD�;��;SE|;sq;Y�f;En\;:R;�9H;�k>;�4;Ie+;�*";�;�B;ȓ;��:�n�:��:6�:?�:+ƭ:�:ʡ�:��:_�d:�pH:~X,:��:���93�9�3~9)�9��08f�l��!�2h������vD��B�G�$���<�'�T���l��A��
���Ù��m�� ��v���Z'Ⱥ3�Ӻhߺ,�����0� ��Z�&���PN�p����"��%(��-��S3�_�8�v{>��D��I��1O���T�6XZ��_���e�%k�$�p�>Bv�3�{���������{M��C���⋻���nw��#B������ؙ��  �  �=m2=��=�~=F$=��=$o=5=� =�] =% =�L�<���<f��<�#�<Vj�<���<I��<_;�<��<���<��<�H�<ɉ�<��<*	�<2G�<#��<��<���<�3�<8l�<*��<���<5�<@�<�q�<L��<l��<���<�%�<�M�<+s�<6��<u��<���<��<0�<��<)�<�5�<>�<�B�<#C�<Y?�<�6�<�)�<-�<3�<��<e��<3��<�n�<�;�<L�<v��<F|�<o/�<��<��<<!�< ��<,L�<��<i]�<���<�U�<ɾ<o6�<��<Z �<]�<���<�<�T�<B��<V�<� �<>\�<���<Ǩ<���<B#�<[L�<�r�<���<ඝ<E՛<��<��<�#�<z:�<EO�<�b�<Dt�<���<���<���<y��<B��<7ł<]π<�}<%�y<��u<�q<��m<b	j<�f<>-b<!@^<5TZ<:iV<�R<0�N<?�J<��F<Q�B<�?<�%;<�G7<�l3<W�/<�+<��'<�$<=S <Ԍ<�<$<�V<��<��	<�R<ѳ<�6�;W�;�;���;�	�;�'�;7W�;ę�;���;�Z�;۹;r�;
 �;2�;(Š;#��;�ϔ;���;AC�;���;�B|;qq;��f;xm\;�9R;�9H;l>;��4;�f+;�,";�";LE;^�;B%�:u�:�:J�:�E�:�˭:8��:規:���:��d:WvH:[\,:�:���9>}�9�$~99708Iom��!��|�������Z��P���$�&�<���T�'�l�+G������Ǚ��p���������S'Ⱥ>�Ӻ�ߺ�������Q� �X�^�R���J����h�"��"(�I�-�,Q3���8��x>�+D�m�I��1O���T��WZ���_���e��k�E�p�Ev���{����_����N����䋻�����x��bC��U���ٙ��  �  �=Z2=��=�~=M$=��=/o=A="� =�] =A =�L�<��<���<�#�<�j�<˰�<���<�;�<��<���<��<�H�<��<��<	�< G�<��<̿�<c��<�3�<�k�<��<���<��<�?�<Eq�<��<)��<]��<�%�<~M�<s�<��<j��<���<1��<E�<��<)�<�5�<F>�<�B�<nC�<�?�<B7�<D*�<h�<}�<H��<���<C��<�n�<�;�<Z�<���<1|�<b/�<���<ف�<!�<ٹ�<L�<���<)]�<d��<�U�<�Ⱦ<6�<ܝ�< �<�\�<z��<��<tT�<+��<I�<� �<]\�<���<Ǩ<���<`#�<�L�<�r�<<��<��<�՛<��<��<>$�<�:�<zO�<�b�<\t�<Ǆ�<֓�<���<f��<4��<ł<Iπ<��}<��y<W�u<��q<z�m<�j<bf<�,b<�?^<�SZ<�hV<AR<�N<�J<��F<-�B<d?<�%;<7H7<m3<��/<�+<�'<i$<�S <`�<��<�<3W<@�<@�	<kS<,�<%7�;��;e�;���;�	�;z'�;�V�;X��;���;@Z�;�ڹ;q�;�;�;4Ġ;d��;�Δ;��;@B�;!��;�A|;Upq;N�f;ql\;o9R;[9H;�l>;��4;�g+;=-";)#;G;�;*�:y�:y�:��:zI�:ZЭ:X��:���:���:i�d:�yH:|^,:o�:��9�z�9n~9�u9��/8˴m���!�����ĺ���n�X�[�$���<��U��l�pI��y��,ə�}r��'������'Ⱥ�Ӻ�ߺي�[���N� �;V������CI�^��g�"�� (��-�mO3�8�8�>x>�sD���I��0O��T��XZ��_���e��k�[�p��Ev�N�{����_���P�����+勻�����y��3D�����Xڙ��  �  	�=X2=��=|~=N$=��='o=Q=.� =�] =H =	M�<��<���<�#�<�j�<��<���<�;�<+��<���<��<�H�<��< ��<	�<"G�<��<���<G��<�3�<�k�<��<���<��<�?�<)q�<��<��<K��<x%�<bM�<s�<��<x��<���<9��<6�<�<@)�<�5�<\>�<�B�<�C�<�?�<]7�<b*�<r�<��<O��<���<U��<*o�<�;�<H�<���<*|�<i/�<���<ˁ�<!�<���<�K�<���<+]�<J��<sU�<�Ⱦ<6�<ޝ�<���<�\�<^��<��<iT�<(��<D�<� �<b\�<���<8Ǩ<��<w#�<�L�<�r�<S��<$��<�՛<��<�<N$�<�:�<�O�<�b�<�t�<���<Г�<���<Y��<>��<ł<?π<e�}<��y<#�u<a�q<��m<�j<f<l,b<�?^<�SZ<�hV<R<��N<��J<��F<9�B<K?<�%;<2H7<�l3<Ȕ/<F�+<8�'<�$<�S <}�<��<<RW<l�<S�	<�S<g�<�7�;G�;�;���;�	�;d'�;W�;O��;]��;�Y�;nڹ;�p�;�;��;�à;���;+Δ;��;�A�;ݣ�;A|;{oq;�f;el\;�9R;9H;%m>;�4;�g+;�.";�#;�G;V�;w+�:�y�:/�:��:$J�:�ѭ:؜�:ګ�:	��:��d:|H:g\,:æ:���9}�9�~9�o9.�/8s�m���!����������t�[���$���<�-U�O�l�1J����gʙ�s��C��K����'Ⱥ��Ӻ%ߺ��������� ��U�~��^���H�.����"�{ (���-�O3�l�8��w>�R
D��I��0O���T��XZ���_��e��k�f�p��Fv��{�B���S����P��h���勻�����y���D�����ڙ��  �  �=Z2=��=�~=M$=��=/o=A="� =�] =A =�L�<��<���<�#�<�j�<˰�<���<�;�<��<���<��<�H�<��<��<	�< G�<��<̿�<c��<�3�<�k�<��<���<��<�?�<Eq�<��<)��<]��<�%�<~M�<s�<��<j��<���<1��<E�<��<)�<�5�<F>�<�B�<nC�<�?�<B7�<D*�<h�<}�<H��<���<C��<�n�<�;�<Z�<���<1|�<b/�<���<ف�<!�<ٹ�<L�<���<)]�<d��<�U�<�Ⱦ<6�<ܝ�< �<�\�<z��<��<tT�<+��<I�<� �<]\�<���<Ǩ<���<`#�<�L�<�r�<<��<��<�՛<��<��<>$�<�:�<zO�<�b�<\t�<Ǆ�<֓�<���<f��<4��<ł<Iπ<��}<��y<W�u<��q<z�m<�j<bf<�,b<�?^<�SZ<�hV<AR<�N<�J<��F<-�B<d?<�%;<7H7<m3<��/<�+<�'<i$<�S <`�<��<�<3W<@�<@�	<kS<+�<$7�;��;e�;���;�	�;z'�;�V�;X��;���;@Z�;�ڹ;q�;�;�;4Ġ;d��;�Δ;��;@B�;!��;�A|;Upq;N�f;ql\;n9R;[9H;�l>;��4;�g+;=-";)#;G;�;*�:y�:y�:��:zI�:ZЭ:X��:���:���:i�d:�yH:|^,:o�:��9�z�9n~9�u9��/8˴m���!�����ĺ���n�X�[�$���<��U��l�pI��y��,ə�}r��'������'Ⱥ�Ӻ�ߺي�[���N� �;V������CI�^��g�"�� (��-�mO3�8�8�>x>�sD���I��0O��T��XZ��_���e��k�[�p��Ev�N�{����_���P�����+勻�����y��3D�����Xڙ��  �  �=m2=��=�~=F$=��=$o=5=� =�] =% =�L�<���<f��<�#�<Vj�<���<I��<_;�<��<���<��<�H�<ɉ�<��<*	�<2G�<#��<��<���<�3�<8l�<*��<���<5�<@�<�q�<L��<l��<���<�%�<�M�<+s�<6��<u��<���<��<0�<��<)�<�5�<>�<�B�<#C�<Y?�<�6�<�)�<-�<3�<��<e��<3��<�n�<�;�<L�<v��<F|�<o/�<��<��<<!�< ��<,L�<��<i]�<���<�U�<ɾ<o6�<��<Z �<]�<���<�<�T�<B��<V�<� �<>\�<���<Ǩ<���<B#�<[L�<�r�<���<ඝ<E՛<��<��<�#�<z:�<EO�<�b�<Dt�<���<���<���<y��<B��<7ł<]π<�}<%�y<��u<�q<��m<b	j<�f<>-b<!@^<5TZ<:iV<�R<0�N<?�J<��F<Q�B<�?<�%;<�G7<�l3<W�/<�+<��'<�$<=S <Ԍ<�<$<�V<��<��	<�R<ѳ<�6�;W�;�;���;�	�;�'�;7W�;ę�;���;�Z�;۹;r�;
 �;2�;(Š;#��;�ϔ;���;AC�;���;�B|;qq;��f;xm\;�9R;�9H;l>;��4;�f+;�,";�";LE;^�;B%�:u�:�:J�:�E�:�˭:8��:規:���:��d:WvH:[\,:�:���9>}�9�$~99708Jom��!��|�������Z��P���$�&�<���T�'�l�+G������Ǚ��p���������S'Ⱥ>�Ӻ�ߺ�������Q� �X�^�R���J����h�"��"(�I�-�,Q3���8��x>�+D�m�I��1O���T��WZ���_���e��k�E�p�Ev���{����_����N����䋻�����x��bC��U���ٙ��  �  6�=2=��=�~=F$=��=o==� =�] =� =bL�<d��<���<-#�<�i�<.��<���<;�<��<`��<e�<�H�<ɉ�<��<(	�<MG�<O��<%��<���<L4�<�l�<���<;��<��<�@�<�q�<���<���<���<&�<�M�<`s�<T��<���<���<��<�<��<�(�</5�<�=�<iB�<�B�<�>�<�6�<�)�<��<� �<���<��<՛�<�n�<�;�<1�<y��<H|�<|/�<)��<)��<�!�<Y��<�L�<`��<�]�<��<BV�<yɾ<�6�<���<� �<s]�<���<V�<�T�<f��<]�<� �<D\�<w��<�ƨ<���<�"�<L�<Fr�<���<w��<�ԛ<%�<Z�<�#�</:�<�N�<=b�<t�<~��<���<���<o��<Q��<Xł<�π<u�}<��y<^�u<��q<��m<!
j<�f<.b<�@^<�TZ<�iV<8�R<��N<��J<G�F<u�B<?<�%;<�G7<�l3<��/<N�+<��'<Y$<�R <�<<�<g<�U<��<	�	<GR<�<�5�;��;F �;���;�	�;s'�;�W�;X��;���;�[�;aܹ;)s�;`!�;��;�Ơ;ؾ�;є;v��;yD�;��;SE|;sq;Y�f;En\;:R;�9H;�k>;�4;Ie+;�*";�;�B;ȓ;��:�n�:��:6�:?�:+ƭ:�:ʡ�:��:_�d:�pH:~X,:��:���93�9�3~9)�9��08f�l��!�2h������vD��B�G�$���<�'�T���l��A��
���Ù��m�� ��v���Z'Ⱥ3�Ӻhߺ,�����0� ��Z�&���PN�p����"��%(��-��S3�_�8�v{>��D��I��1O���T�6XZ��_���e�%k�$�p�>Bv�3�{���������{M��C���⋻���nw��#B������ؙ��  �  [�=�2=��=�~==$=��=�n= =Ƹ =f] =� =�K�<��<s��<�"�<ai�<���<h��<�:�<9�<��<-�<VH�<���<���<A	�<wG�<���<p��<��<�4�<�l�<��<���<�<A�<kr�<D��<8��<O��<U&�<*N�<�s�<w��<���<���<��<��<��<�(�<�4�<n=�<�A�<QB�<o>�<6�< )�<B�<e �<C��<���<���<zn�<^;�<�<k��<H|�<�/�<W��<q��<�!�<���<M�<���<q^�<���<�V�<ʾ<b7�<��<*�<�]�<J��<��<U�<���<��<� �<5\�<Q��<�ƨ<Q��<�"�<�K�<�q�<(��<ﵝ<oԛ<��<�
�<!#�<�9�<�N�<�a�<�s�<H��<���<���<|��<x��<ył<�π<�}<��y<O�u<��q<��m<j<�f<�.b<B^<�UZ<�jV<��R<Q�N<V�J<��F<��B<�?<�%;<�G7<&l3<��/<��+<M�'<m$<�Q <�<!�<c<�T<�<��	<kQ<\�<G4�;��;^��;O��;C	�;�'�;X�;���;���;�\�;�ݹ;�t�;m#�;��;�Ƞ;���;�Ҕ;���;@F�;���;�G|;Euq;R�f;8o\;�:R;�9H;!k>;��4;mc+;�(";�;@;��;��:�e�:��:��:�6�:>��:t��:��:3�:K�d:�iH:S,:#�:ي�9���9�F~9ɸ95#18�3l��O!�J���m���$��1��$��<�b�T�U�l�;����������j��	������O(Ⱥ��Ӻ5"ߺ������ܯ ��]������R�Q���"��)(���-�]W3���8�-~>��D���I��2O�,�T��WZ���_��e��k��p�x?v�w�{����������K���������㪎�au��C@��p���י��  �  ��=�2=��=�~=9$=��=�n=�=�� =&] =� =]K�<P��<���<
"�<�h�<��<���<&:�<�~�<���<��<(H�<���<���<R	�<�G�<���<���<���<(5�<m�<���<[��<��<�A�<s�<͢�<���<���<�&�<�N�<�s�<���<���<���<���<��<A�<3(�<v4�<�<�<gA�<�A�<�=�<�5�<�(�<��<���<���<C��<��<%n�<;�<��<X��<Z|�<�/�<���<���<H"�<,��<�M�<m��< _�<O��<wW�<�ʾ<
8�<���<��<k^�<˵�<�<PU�<���<��<!�<\�<0��<cƨ<��<,"�<4K�<Cq�<���<Y��<�ӛ<�<D
�<�"�<.9�<N�<�a�<}s�<��<`��<{��<���<���<�ł<)Ѐ<ٳ}<g�y<N�u<��q<
�m<cj<�f<E0b<9C^<�VZ<�kV<�R<-�N<��J< �F<��B<�?<u%;<fG7<�k3<Ғ/<��+<J�'<[$<sP <ډ<��<<}S<��<��	<QP<`�<�2�;�;���;���;-	�;�'�;GX�;ț�;��;z^�;�߹;�v�;U%�;��;�ʠ;)Ú;`Ք;��;)H�;���;�J|;Kxq;U�f;�p\;O;R;�9H;Kj>;C�4;Ha+;�%";�;�;;s�;?�:�\�:���:���:-�:���:^��:瓏:Z�:��d:�`H:�M,:�:���9
��9(\~9��9��18QIk��!��)��M��1������$���<���T�_�l�f3��h�������f�����s����'Ⱥ��Ӻ�$ߺ���J��l� ��a�t���iW�x��Ĕ"��.(��-��[3�
�8��>�ID�S�I�/4O���T�YWZ�L�_��}e��k���p�<v�~�{�����Q~��I�����ދ�����Us��5>���	���ՙ��  �  ��=�2=��=�~=5$=��=�n=�=g� =�\ =A =�J�<���<<��<\!�<+h�<q��<R��<�9�<K~�<T��<��<�G�<c��<���<b	�<�G�<��<��<���<�5�<n�<-��<���<g�<PB�<�s�<\��<U��<T��<7'�<�N�<*t�<��<ζ�<���<���<��<�<�'�<4�<c<�<�@�<%A�<:=�<�4�<�'�<�<6��<=��<���<���<�m�<�:�<��<C��<f|�<�/�<���<
��<�"�<���<N�<��<�_�<���<2X�<i˾<�8�<O��<`�<�^�<B��<i�<�U�<��<��<
!�<�[�<��<ƨ<���<�!�<�J�<�p�<�<���< ӛ<g�<�	�<�!�<�8�<�M�<a�<s�<ԃ�<5��<m��<���<���<�ł<fЀ<��}<U�y<h�u<��q<;�m<�j<[f<�1b<qD^<6XZ<mV<ԂR<�N<z�J<��F<N�B<�?<e%;<G7<Sk3<�/<�+<I�'<M$<0O <|�<��<�	<5R<N�<��	<7O<[�<1�;��;���;���;��;�'�;�X�;���;���;�_�;.�; y�;�'�;(�;r͠;�Ś;�ה;��;wJ�;���;.N|;{q;�f;]r\;�;R;�9H;�i>;��4;_+;�"";�;j7;�;r�:R�:Z��:p��:�"�:���:jz�:{��:<܀:+�d:AXH:LH,:<�:h��9���9�y~9��9�28)sj�9� �|���(�����	��s$�]�<���T���l�(,������Z���Db��5��_����'Ⱥ�Ӻ�'ߺל꺋��&� ��e����h\������"��3(��-��_3��8�V�>�WD��I�{5O���T��VZ�B�_�{{e��k�K�p�L8v��{�:����{��RF����cۋ�.����p���;�����.ԙ��  �  ό=�2=��=�~=,$=}�=�n=�=0� =�\ =�  =&J�<��<���<� �<g�<ۭ�<���<9�<�}�<���<D�<�G�<F��<���<p	�<�G�<@��<o��<i��<6�<�n�<Х�<���<�<�B�<Ut�<��<���<���<�'�<RO�<yt�<��<���<���<���<j�<��<�'�<�3�<�;�<H@�<�@�<�<�<14�<2'�<o�<���<���<O��<K��<~m�<�:�<��<9��<k|�<0�<��<[��<#�<��<�N�<���<W`�<���<�X�<̾<h9�<��<��<~_�<���<��<�U�<6��<��<!�<�[�<͒�<�Ũ<N��<O!�<6J�<p�<b��<��<wқ<��<	�<e!�<8�<(M�<�`�<�r�<���<��<[��<���<Ϻ�<'Ƃ<�Ѐ<v�}<I�y<r�u<�q<��m<�j<� f<�2b<�E^<sYZ<nV<ӃR<�N<8�J<�F<��B<�?<G%;<�F7<�j3<��/<>�+<[�'<'$<�M <>�<4�<;<�P<�<Z�	<N<[�<W/�;p�;Y��;.��;��;�'�;cY�;}��;L��;�a�;�;�z�;�)�;��;�Ϡ;EȚ;.ڔ;T�;�L�;t��;�Q|;�}q;S�f;�s\;�<R;�9H;�h>;��4;�\+; ";s;�3;2�;���:�G�:
��:A��:�:_��:�p�:���:�Հ:\�d:�OH:�@,:��:���9���9��~9�9T\38��i�"� ��߂�G���ª����k_$�љ<��T�g�l��#������\���@^�����Y���](Ⱥ��Ӻ�+ߺ��꺔���� ��i���u���a�B��"��8(���-�Ld3���8���>�sD�K�I� 7O��T��VZ��_�ze��k��p��4v���{�߮��Gy���C��W���؋�����n���9������ҙ��  �  ��=3=��=�~=%$=q�=|n=^=�� =u\ =�  =�I�<w��<���<  �<�f�<M��<6��<�8�<f}�<���<��<zG�<5��<���<�	�<H�<z��<���<���<�6�<o�<R��<4��<��<�C�<�t�<���<e��<\��<(�<�O�<�t�<C��<��<���<���<I�<|�<('�<)3�<v;�<�?�<@�< <�<�3�<�&�<��<'��<(��<���<ڙ�<m�<c:�<o�<,��<g|�<'0�<7��<���<v#�<���<6O�<8��<�`�<N��<�Y�<�̾<:�<���<��<`�<(��<8	�<4V�<h��<��<
!�<�[�<���<�Ũ<���<� �<�I�<�o�<ے�<w��<�ћ<�<i�<� �<�7�<�L�<@`�<�r�<L��<钊<J��<���<�<WƂ<р<�}<9�y<}�u<#�q<��m<6j<"f<4b<�F^<~ZZ<#oV<фR<��N<�J<��F<��B<?<,%;<�F7<Jj3<��/<b�+<u�'<$<�L <
�<��<<{O<�<E�	<M<l�<�-�;$�;J��;���;D�;(�;�Y�;:��;��;�b�;��;�|�;�+�;��;Ҡ;�ʚ;nܔ;w�;wN�;j��;�T|;I�q;��f;�t\;�=R;9H;
h>;��4;�Z+;�";�;�/;�};���:�=�:Y��:���:L�:'��:sh�:�{�:!΀:��d:GH:�;,:��:���9`��9ͤ~9�C9�48��h��L �����hڴ�7�湷���K$�C�<���T�,zl�x���ꍺ֨��oZ�����
���)Ⱥ��ӺE/ߺ ����9� ��m�������f����"��=(���-��h3�Q�8�8�>�D�F�I��7O���T��VZ���_��xe� 
k���p��0v���{�٬���v��yA������֋�)���wl���7�����?љ��  �  �="3=�=�~=$=]�=gn=9=׷ =D\ =z  =I�<��<p��<��<bf�<¬�<���<"8�<}�<<��<��<XG�<��<���<�	�<5H�<���<��<��<�6�<�o�<Ԧ�<���<*�<D�<uu�<��<���<���<t(�<�O�< u�<o��<)��<���<���<!�<D�<�&�<�2�<;�<P?�<�?�<~;�<3�<&�<T�<���<���<j��<���<�l�<+:�<M�<��<x|�<B0�<j��<��<�#�<���<�O�<���<ta�<���<Z�<N;<�:�<��<�<j`�<���<�	�<uV�<���<�<!�<�[�<���<bŨ<���<� �<KI�<*o�<O��<���<Vћ<��<��<Y �<7�<NL�<�_�<4r�<��<���<3��<���<��<�Ƃ<Lр<Ŷ}<��y<P�u<1�q<��m<Kj<#f<35b<�G^<�[Z<	pV<��R<D�N<e�J<��F<3�B<*?<%;<FF7<�i3<_�/<չ+<��'<"$<�K <��<��<�<zN<Ŝ<8�	<L<��<M,�;��;���;��;��;7(�;;Z�;��;T��;d�; �;�~�;�-�;���;Ԡ;�̚;rޔ;M
�;�P�;Ű�;iW|;��q;*�f; v\;>R;f9H;�f>;Q�4;�X+;�";Y;L,;1z;k��:�5�:��:*��:=�::�`�: u�:wɀ:W�d:g?H:�6,:b�:��9n��9]�~99`9ן48%h�v! �����!���Pc����2;$�:v<���T��il�W��^卺�����V������ϗ��g)Ⱥ�Ӻe1ߺ�������� ��q���=���j�j��"��A(�B�-�/l3�s�8�_�>�oD���I�9O���T�WVZ���_��ve�dk�ޚp�.v���{������t��S?���	��iԋ�:���ij��6������ϙ��  �  /�=83=�=�~= $=T�=Tn==�� =\ =S  =�H�<���<��<�<f�<Y��<b��<�7�<�|�<���<y�<8G�<���<���<�	�<BH�<߅�<6��<w��<D7�<�o�<(��<��<��<|D�<�u�<o��<I��<
��<�(�<7P�<*u�<���<(��<���<���<�<�<�&�<�2�<�:�<?�<#?�<$;�<�2�<�%�<��<7��<g��<��<E��<�l�<�9�<4�<��<�|�<H0�<���<��<$�<]��<�O�<&��<�a�<Q��<�Z�<�;<;�<y��<g�<�`�<ﷶ<�	�<�V�<���<�<!�<�[�<l��<0Ũ<f��<G �<�H�<�n�<鑟<���<�Л<<�<��<��<�6�<�K�<�_�<�q�<�<���<4��<���<��<�Ƃ<xр<`�}<��y<��u<��q<r n<"j<�#f<6b<�H^<=\Z<�pV<)�R<�N<ĴJ<M�F<9�B<-?<%;< F7<�i3<��/<E�+<��'<�$<#K <�<�<�<�M<�<��	<QK<��<#+�;�
�;��;���;��;(�;UZ�;���;��;ge�;D�;��;�.�;+��;�ՠ;�͚;	��;��;�Q�;���;8Z|;{�q;W�f;	w\;�=R;Y9H;�f>;M�4;#W+;j";�	;o);�w;W��:�/�:6��:��:� �:���:�[�:Vo�:QĀ:ɧd:�8H:!3,:��:̍�9���9��~9�t9�58Eg����]���w����H�����.$��i<��zT��_l�I��]ߍ�T���T�����������(Ⱥ��Ӻ>3ߺ����k� �Lt�_ ����nm���0�"��D(��-��n3�@ 9���>�kD���I��9O���T�MVZ��_��ue��k�q�p�o+v��{�Z����s���=��^���ҋ�ʝ��
i���4��\���Ι��  �  <�=C3=�=�~=$=K�=Bn==�� =\ =7  =�H�<E��<���<��<�e�<��<!��<�7�<�|�<���<e�<G�<��<���<�	�<aH�<���<L��<���<z7�< p�<p��<[��<��<�D�<v�<���<{��<D��<�(�<?P�<Eu�<���<J��<���<���<��<��<�&�<o2�<�:�<�>�<�>�<�:�<r2�<q%�<��<���<#��<��<#��<�l�<�9�<�<
��<r|�<i0�<���<;��<$�<v��<,P�<[��< b�<���<�Z�<ξ<I;�<ɢ�<��<�`�<��<�	�<�V�<͞�<2�<
!�<�[�<J��< Ũ<M��<' �<�H�<�n�<���<Y��<�Л<��<;�<��<�6�<�K�<�_�<�q�<т�<���<(��<���<0��<�Ƃ<�р<p�}<��y<b�u<]�q< n<�j<V$f<�6b<CI^<�\Z<qV<��R<�N<��J<{�F<��B<B?<�$;<�E7<bi3<��/<��+<��'<$<�J <��<��<�<M<e�<��	<�J<��<�*�;
�;Z��;h��;��;U(�;�Z�;���;M��;�e�;�;���;0�; ��;�֠;�Κ;���;��;�R�;Ҳ�;[|;��q;�f;�w\;�>R;�8H;tf>;��4;gV+;�";�;?(;}u;{��:�*�:H��:`��:���:���:�W�: m�:
:��d:�6H:�/,:k�:���9���9�~99�9058g����(|�����c:���i&$��a<��qT�VYl����zލ�=����R�����H���2*Ⱥ��Ӻ�5ߺ�����z� ��u�n"�j���o���@�"�G(��-�|p3�K9��>�*D��I�`:O���T�2VZ���_��te�(k�3�p�*v�H�{�m����r���<��<���ы�����h���3��� ��nΙ��  �  ݊=d0=��=�z=�=��=Qi=�=ұ =�U =$��<N:�<��<|��<z�<S�<8��<���<� �<Td�<��<
��<!*�<nj�<���<���<�$�<�`�<B��<���<��<�C�<�x�<��<G��<�<3?�<�l�<���<\��<���<v�<�/�<�O�<�l�<��<'��<���<���<���<���<���<t��<6��<���<���<���<���<���<�r�<cO�<�&�<I��<"��<��<�I�<M�<���<�c�<

�< ��<�C�<B��<\d�<I��<l�<��<�[�<�ʼ<�4�<���<Q��<�P�<c��<��<�?�<N��<Qȭ<Q�<@�<?v�<ɨ�<ؤ<6�<h-�<�S�<�w�<���<��<�֗<9�<�<b$�<;�<YP�<>d�<�v�<t��<Ę�<C��<Ͷ�<�Ā<��}<�y<Y�u<_�q<�n<cj<4f<Lb<�d^<�}Z< �V<8�R<��N<u�J<�G<�-C<wP?<�u;<�7<��3<a�/<#,<{V(<u�$<�� <E<�L<$�<.�<�9<��
<��<�]<A��;X��;'�;"��;���;S��;��;�]�;v��;�8�;�Ļ;yf�;��;O�;�Ӣ;BҜ;B�;�;�b�;BŅ;yA�;�u;^k;`;`V;�TL;�{B;�8;YX/;5&;��;$;�A;r�;y~�:]��:��:���:~3�:Pפ:l��:��:��p:�S:KW7:�X:�a�9T��9ܒ9j;9�+�8�/��;���qd�0褹�(׹\{�p/���5��N��3f�F9~����i햺G���6���X;��K�ź��Ѻ�"ݺf���9������Y��M�I��z��MX���!�֡'�B-���2�z8�
>�R�C��BI�Y�N��nT�/Z���_�=4e���j�vdp���u�v�{������e���3��B��oϋ������l��Q<������ݙ��  �  ؊=k0=��=�z=�=��=Si=�=� =�U =5��<e:�<#��<���<��<2S�<A��<���<� �<ed�< ��<��<!*�<Hj�<���<���<�$�<�`�<8��<���<��<�C�<�x�<Ѭ�<1��<��<,?�<vl�<��<G��<���<p�<�/�<�O�<�l�<���<��<��<���<���<��<���<���<I��<���<��<���<���<���<�r�<iO�<�&�<[��<+��<���<�I�<\�<���<�c�<
�<��<�C�<-��<Fd�<&��<�k�<��<�[�<�ʼ<e4�<���<B��<�P�<[��<
��<�?�<X��<Wȭ<*�<@�<Jv�<ߨ�<#ؤ<@�<�-�<�S�<
x�<���<8��<�֗<Q�<*�<i$�<!;�<hP�<Fd�<�v�<i��<֘�<J��<ٶ�<�Ā<��}<̼y<=�u<'�q<�n<Nj<�3f<�Kb<zd^<�}Z<�V<�R<��N<^�J<�G<�-C<�P?<�u;<��7<��3<|�/<K#,<�V(<��$<�� <\<�L<g�<`�<�9<ϔ
<��<�]<���;���;)�;���;���;���;�;7^�;R��;�8�;�Ļ;Cf�;�;�;ZӢ;�ќ;*�;�;Lb�;�ą;8A�;ǭu;Hk;�`;^`V;UL;�zB;��8;�X/;�&;��;S;}B;�;��:���:0��:��:�4�:�ؤ:ؾ�:��:�p:2�S:�U7:U:�e�9'��9�ݒ96;9�'�8ax���N���|d����*׹�~�l2�D�5��N��5f��:~�����햺����򂮺�:����ź݊Ѻ!#ݺ���q8��=�����QL����Ь�/W���!�p�'�IA-���2��y8�	>�ݪC�FBI�'�N�<oT��Z�i�_��3e���j��dp��u��{����Tf���3������ϋ����m���<������ݙ��  �  Ǌ=\0=��=�z=�=��=gi=�=� =�U =^��<�:�<R��<���<��<YS�<q��<��<!�<�d�<4��<%��<K*�<\j�<���<���<�$�<|`�<��<���<��<fC�<�x�<���<��<��<?�<El�<Ǘ�<)��<c��<W�<�/�<�O�<�l�< ��<��<��<���<���<1��<���<���<x��<���<*��<ѽ�<ϩ�<��<�r�<�O�<�&�<f��<D��<��<�I�<b�<���<jc�<�	�<���<�C�<	��<&d�<���<�k�<��<�[�<�ʼ<:4�<h��<��<�P�<;��<���<�?�<E��<dȭ<;�<>@�<[v�<�<Aؤ<^�<�-�<(T�<2x�<љ�<]��<�֗<��<U�<�$�<>;�<pP�<ld�<�v�<x��<Ԙ�<)��<���<�Ā<\�}<��y<�u<��q<cn<�j<�3f<�Kb<d^<o}Z<��V<ϲR<\�N<�J<�G<v-C<�P?<�u;<�7<��3<��/<}#,<�V(<�$<:� <�<:M<��<��<X:<;�
<*�<�]<��;ӄ�;��;��;��;c��;��;�]�;���;88�;Ļ;�e�;z�;o�;�Ң;Iќ;��;N�;�a�;�ą;�@�;�u;Rk;c�`;�_V;AUL;�{B;��8;�Y/;&;��;8;�C;��;E��:���:"��:���:�7�:�ۤ:���:��:��p:��S:�Z7:'W:�g�9���9�ג9~;9��8����o����d������4׹a���6�~�5��N�I9f�H?~���������܄���;����ź��Ѻ� ݺv��27��C���	���J�������NV���!��'��?-���2��x8�'>���C�AI�G�N��nT��Z�n�_��4e��j��ep�,�u�Ø{�����g��l4��S��MЋ�̞���m���<��c��Wޙ��  �  ��=P0=��=�z=�=��=hi=�=� =V =���<�:�<���<��<�<�S�<���<W��<_!�<�d�<e��<E��<G*�<mj�<���<���<�$�<]`�<���<M��<X�<C�<ux�<P��<���<��<�>�<
l�<x��<���<(��<$�<�/�<�O�<�l�<��<+��<��<���<���<d��<+��<���<���<M��<���</��<��<��<s�<�O�<'�<���<X��<��<�I�<N�<���<ac�<�	�<ɩ�<mC�<���<�c�<���<fk�<A�<*[�<Sʼ<�3�<��<���<uP�<��<���<�?�<9��<Pȭ<J�<3@�<tv�<"��<~ؤ<��<�-�<rT�<�x�<3��<���<'ח<��<��<�$�<l;�<�P�<rd�<w�<|��<˘�<7��<���<fĀ<�}<�y<z�u<P�q<�n</j< 3f<�Jb<�c^<�|Z<�V<X�R<��N<��J<TG<�-C<vP?<�u;<�7<��3<��/<�#,<hW(<p�$<�� <b	<�M<n�<_�<�:<��
<��<�^<��;h��;��;E��;���;Z��;��;f]�;s��;l7�;9û;�d�;��;)�;�Ѣ;(М;��;r�;�`�;�Å;�?�;��u;}
k;6�`;�_V;�TL;|B;��8;EZ/;�&;��;�;�E;��;j��:;�:��:���:�;�:Dߤ:�ŕ:��:�p:��S:�Z7:XY:�c�9[��9�֒9��:9�ݢ8E�W�����d��	��ZN׹��qA�7�5��N��Cf�G~������¢�~���<����źv�Ѻ� ݺ����3��H�������H�)����7S� �!�y�'��=-���2��v8��>�T�C��@I��N��nT�Z�	�_�J5e���j�>gp�v��{�����'h��6��q���ы������n��>��K��4ߙ��  �  ��=40=��=�z= =��=i=�= � =(V =���<1;�<��<j��<~�<�S�<��<���<�!�<�d�<���<���<p*�<�j�<���<���<|$�<*`�<͚�<��<"�<�B�<x�<���<U��<3�<?>�<�k�<��<���<���<��</�<gO�<�l�<���<<��<5��<���< ��<���<p��<D��<��<���<���<���<r��<���<js�<P�<3'�<���<���<9��<�I�<J�<s��<*c�<�	�<���<*C�<���<_c�<\��<k�<��<�Z�<�ɼ<�3�<���<���</P�<ޤ�<���<�?�<)��<Qȭ<a�<W@�<�v�<U��<�ؤ<��<;.�<�T�<�x�<���<��<�ח<�<��<%�<�;�<�P�<�d�<-w�<���<Ę�<��<u��<:Ā<z�}<��y<��u<|�q<.n<qj<O2f<Jb<�b^<|Z<i�V<�R<k�N<��J<�G<M-C<eP?<�u;<N�7<[�3<~�/<J$,<�W(<�$<u� <'
<�N<?�<�<�;<l�
<n�<�^<��;���;���;��;��;J��;j�;�\�;޿�;�6�;|»;Rc�;*�;��;Т;�Μ;��;G�;!_�;�;?�;$�u;.	k;��`;W_V;�TL;�|B;�8;\/;�&;�;
;�H;��;-��:c�:?��:2��:"B�:��:{ʕ:��: �p:��S:_7:
\:d�9���9*ʒ9�:9.��8:۸�����-�d���:e׹d��>M��5�w#N�6Pf��M~��������Ţ�܆���<��l�ź��ѺhݺH��v0��N���-��JF�'��n��(P�>�!���'��:-���2��t8�>��C�^?I���N�:nT�DZ���_�	7e�I�j�ip��v�Y�{�Y���si��y7�����DӋ�O���Lp��l?��!��,����  �  ��=*0=��=�z= =��=�i==K� =WV =W��<�;�<v��<���<��<T�<���<��<"�<ae�<��<���<�*�<�j�<���<���<_$�<`�<���<���<��<dB�<�w�<���<���<��<�=�<@k�<���<E��<���<��<O/�<QO�<�l�<���<7��<_��<��<N��<���<���<���<���<��<W��< ��<��<���<�s�<mP�<�'�<��<���<e��<�I�<O�<a��<
c�<^	�<I��<�B�<��<c�<���<�j�<R�<;Z�<}ɼ<!3�<L��<,��<�O�<���<`��<�?�<��<Vȭ<[�<�@�<�v�<���<٤<L�<�.�<GU�<Oy�<��<���<�ח<��<P�<o%�<�;�<Q�<�d�<Iw�<���<̘�<��<a��<Ā<�}<ͺy<�u<��q<@n<�j<51f<(Ib<�a^<W{Z<��V<�R<��N<�J<�G<-C<hP?<�u;<s�7<��3<��/<�$,<�X(<�$<L� <<�O<,�<�<�<<Q�
<<�<�_<)��;=��;���;��;J��;W��;�;X\�;���;U5�;���;)b�;��;<�;D΢;�̜;��;x�;�]�;+��;�=�;+�u;�k;�`;�^V;oUL;�|B;v�8;L]/;o&;Q�;�;�K;D�;Ɣ�:��:���:���:�I�:��:�ϕ:j�:��p:��S:7e7:�[:�f�9���9�Ò9z�:9�k�89^��+M���e�-=��ۀ׹��T]���5�&1N� Zf��Z~���������Ǣ�����'=����ź��Ѻ.ݺ��>,�����N���B�V��q���L�Q�!��'��7-���2��q8�;>�ʥC�>I��N�>nT�Z���_��7e��j�Kkp�
v�U�{�����Lk��M9����� Ջ�#����q���@�����Xᙻ�  �  [�=0=��=�z=	 =��=�i=$=y� =�V =���<<�<��<k��<l�<�T�<��<���<p"�<�e�<A��<���<�*�<�j�<���<r��<@$�<�_�<7��<��<Y�<�A�</w�<��<i��<5�<]=�<�j�<O��<տ�<H��<e�</�<7O�<ul�<��<C��<���<C��<���<Q��<!��<��<���<���<���<{��<e��<Z��<At�<�P�<�'�<H��<���<���<�I�<F�<1��<�b�<	�<���<B�<���<�b�<S��<j�<��<�Y�<�ȼ<�2�<ٖ�<���<�O�<6��<��<Y?�<�<Rȭ<j�<�@�<�v�<䩦<_٤<��</�<�U�<�y�<���<��<nؗ<��<��<�%�<Z<�<KQ�<e�<hw�<���<���<ৄ<B��<�À<m�}<8�y<B�u<��q<9n<�j<?0f<MHb<�`^<_zZ<ДV<h�R<T�N<]�J<bG<�,C<DP?<�u;<��7<%�3<.�/<�%,<QY(<��$<0� <<�P<1�<#�<�=<B�
<�<�`<���;#��;y��;���;z��;��;��;�[�;ɽ�;�4�;���;�`�;��;X�;�̢;˜;R�;��;X\�;���;�<�;�u;�k;f�`;�]V;eUL;*}B;��8;�^/;�&;;�;�;�O;��;���:��:���:���:+P�:��:֕:.��:�p:9�S:j7:y]:f�9���9���9#�:9��8�G��7���Ee��\����׹���k���5�"AN�&gf��g~� �����]ˢ�����:?����źN�Ѻ+ݺl���&��s���F��k?����~���H�K�!�6�'�&4-�d�2��n8�Z	>��C�f<I��N��mT�pZ�џ_��8e���j�Kmp�]v���{�����Tm���:������֋�+����s���B����G♻�  �  ?�=�/=��=�z= =�=�i=O=�� =�V =*��<�<�<k��<���<��<jU�<���< ��<�"�<�e�<���</��<�*�<�j�<���<g��< $�<�_�<���<#��<�
�<�A�<�v�<���<���<��<�<�<Tj�<ݕ�<t��<���<�<�.�<	O�<al�<��<g��<���<���<���<���<���<���<n��<��<C��<��<٫�<ג�<�t�<6Q�<#(�<���<��<���<J�<A�<��<�b�<��<���<B�<5��<b�<���<�i�<I�<8Y�<rȼ<#2�<a��<T��<)O�<룴<��</?�<݅�<Qȭ<��<�@�<@w�<%��<�٤<�<}/�<0V�<7z�<���<p��<�ؗ<s��<%�<(&�<�<�<�Q�<6e�<�w�<���<���<ʧ�<��<|À<��}<��y<{�u< �q<Y n<�j<?/f<IGb<�_^<{yZ< �V<��R<��N<��J<�
G<�,C<4P?<�u;<�7<u�3<��/<+&,< Z(<��$</� <<�Q<0�<�<�><8�
<��<$a<О�;���;��;O��;ť�;��;[�;[�;��;?3�;L��;_�;>�;��;�ʢ;2ɜ;p��;��;�Z�;��;L;�;��u;=k;�`;X]V;sUL;m~B;��8;�`/;V&;�;H;�R;��;a��:#�:��:P��:;X�:R��:�ܕ:���:�p:��S:�m7:�b:�f�9���9g��9��:94ҡ8^�������}e�bw��i�׹���={���5��NN��tf�Cs~��%��<��w΢������?���źɂѺ�ݺ��躊"��G���ц��;�������D���!�6�'�20-�
�2�l8��>�@�C��:I��N�*mT��Z���_�Y:e�B�j�pp�v�٦{�F���o���<���
���؋�즎�Vu�� D��v���㙻�  �  2�=�/=�=�z= =�=�i=m=�� =�V =���<�<�<ރ�<O��<q�<�U�<���<S��<?#�<if�<ɨ�<g��<	+�<�j�<���<h��< $�<}_�<ә�<���<�
�<&A�<Yv�<��<m��<C�<_<�<�i�<q��<��<���<��<�.�<�N�<cl�<��<o��<���<���<'��<���<���<���<���<{��<���<r��<D��<K��<�t�<�Q�<}(�<���<<��<���<J�<0�<��<b�<��<a��<�A�<���<�a�<_��<i�<��<�X�<�Ǽ<�1�<<���<�N�<���<��< ?�<څ�<@ȭ<��<�@�<nw�<d��< ڤ<r�<�/�<�V�<�z�<��<껙<`ٗ<���<y�<�&�<�<�<�Q�<Se�<�w�<���<���<ħ�<ܵ�<dÀ<!�}<��y<��u<%�q<i�m<�j<X.f<BFb<_^<�xZ<5�V<�R<��N<��J<�
G<x,C<+P?<�u;<�7<��3<T�/<�&,<�Z(<O�$<�� <�<�R<O�<��<�?<�
<��<b<��;���;���;ƌ�;ť�;'��;��;~Z�;w��;�1�;	��;�]�;��;��;�Ȣ;�ǜ;�ޖ;*�;Y�;ɼ�;�9�;ءu;tk;��`;�]V;4UL;�~B;��8;@b/;�&;�;{;SU;O�;U��:h&�:i��:>�:�_�:>��:�:��:��p:-�S:�p7:�c:�c�9���9���9�}:9�82P��Rt����e�q���[�׹��I���6�
\N�7�f��}~��+������Т�/����?����ź��Ѻ=ݺe��J��Ȗ�����^9���s���@��!���'�*--�o�2��h8�>�H�C�:I�:�N�mT��Z���_��;e��j�}rp�4v��{������p���>������ڋ����� w���E�����噻�  �  �=�/=l�=�z= =#�=�i=�=ܲ =�V =���<F=�<6��<���<��<;V�<N��<���<�#�<�f�< ��<���<@+�<�j�<���<Z��<�#�<I_�<���<���<d
�<�@�<�u�<���<��<��<<�<yi�<��<˾�<Z��<��<p.�<�N�<Hl�<���<x��<��<���<Q��<��<$��<6��<7��<���<!��<���<���<���<Yu�<�Q�<�(�<���<b��<ۊ�<J�<)�<���<Ub�<m�<��<xA�<���<Ia�<���<�h�<d�<OX�<�Ǽ<E1�<���<���<�N�<h��<x�<�>�<Å�<=ȭ<��<A�<�w�<���<5ڤ<��<30�<�V�<{�<Ԝ�<H��<�ٗ<7��<��<�&�<'=�<R�<�e�<�w�<���<���<���<���<À<��}<[�y<�u<s�q<��m<�j<�-f<�Eb<H^^<�wZ<��V<~�R<|�N<�J<2
G<,,C<P?<�u;<Z�7<�3<��/<G',<F[(<�$<�� <�<ES<�<��<^@<ƚ
<h�<b<���;O��;x��;?��;���;
��;��;�Y�;_��;11�;��;G\�;K�;��;�Ǣ;Ɯ;eݖ;��;�W�;���;9�;3�u;�k;��`;�\V;/UL;7B;�8;�c/;&;�;D;�X;:�;��:j,�:;��:��:Ae�:��:��:��:C�p:y�S:�v7:5e:pc�9��9���9=`:9�]�8b	������w�e�N���)�׹:��F��%6�2hN��f�{�~��.��q	��CԢ�]����@����źu�Ѻ�ݺ�����F������
6��������=��!��'�*-�x�2�g8�>��C�a8I�(�N��lT�3Z�ۡ_�7=e���j�Ctp��v�a�{�Z���fr��I@��2��&܋�A���qx���F������噻�  �  ��=�/=e�=�z= =�=�i=�=�� =W =&��<�=�<���<
��<�<�V�<���<	��<�#�<�f�<6��<���<O+�<�j�<���<T��<�#�<B_�<]��<d��<
�<�@�<�u�<j��<���<�<�;�</i�<��<}��<��<d�<U.�<�N�<4l�<���<~��<߲�<���<x��<U��<b��<���<l��<2��<r��<��< ��<Փ�<�u�<R�<�(�<'��<���<ۊ�<J�<6�<��<Tb�<P�<��<<A�<.��<a�<���<Ph�<��<�W�<7Ǽ<�0�<O��<R��<NN�<5��<f�<�>�<���<Eȭ<��<A�<�w�<Ū�<mڤ<��<0�<.W�<j{�<��<���<	ڗ<v��<&�<'�<`=�<,R�<�e�<�w�<ǈ�<���<���<���<�<N�}<ͷy<��u<�q<
�m<Vj<�,f<�Db<�]^<qwZ<�V<�R<�N<��J<-
G<,C<P?<v;<C�7<F�3<��/<�',<�[(<��$<H� <R<T<��<��<�@<h�
<��< c<��;΋�;Ȅ�;+��;9��;	��;��;�Y�;κ�;�0�;ﺻ;l[�;j�;F�;SƢ;�Ĝ;+ܖ;��;W�;v��;78�;��u;� k;Ε`;Q\V;�UL;xB;�8;�d/;O&;�;E;D[;��;��:�1�:+��:P�:�h�:
�:��:!
�:�p:��S:w7:�e:�g�9N��9k��9T:9�)�8y濷%��;�e�龥��عG��Z��d!6�.pN�u�f���~�2��I��բ�����uA����ź܀Ѻ�ݺØ躾���������3����J���;�7�!�M�'�(-��2�6e8�B>��C�u7I�{�N��lT��Z�R�_� =e���j��up�v���{�6����s���A�����f݋�����Ty��H������晻�  �  �=�/=[�=�z= =-�=j=�=� =-W =@��<�=�<���<2��<7�<�V�<�<'��<�#�<�f�<O��<���<k+�<k�<���<E��<�#�<_�<T��<F��<�	�<g@�<�u�<@��<���<b�<�;�< i�<���<^��<���<Q�<?.�<�N�<"l�<��<���<���<��<���<w��<���<���<���<[��<���<;��<'��<���<�u�<)R�<)�<?��<���<��<0J�<)�<ҵ�<*b�<3�<ӧ�<A�<��<�`�<y��<#h�<��<�W�<Ǽ<�0�<��<3��<-N�<(��<A�<�>�<���<@ȭ<��<$A�<�w�<۪�<�ڤ<�<�0�<^W�<�{�<C��<ȼ�<3ڗ<���<@�<&'�<|=�<MR�<�e�<�w�<҈�<���<~��<���<�<$�}<��y<=�u<��q<��m<j<�,f<�Db<E]^<wZ<��V<��R<��N<��J<�	G<�+C<�O?<v;<��7<��3<'�/<�',<\(<ԓ$<�� <�<XT<�<��<QA<��
<3�<Kc<V��;g��;D��;���;I��;���;�;:Y�;���;$0�;���;�Z�;��;�ߨ;�Ţ;9Ĝ;�ۖ;��;FV�;��;�7�; �u;% k;��`;�[V;[UL;�B;�8;�e/;5&;�;a;#\;>�;���:�3�:l��:��:fk�:��:��:b�:H�p:��S:Iz7:�h:�d�9/��9z��9@G:9R�8�c���-��f��ʥ��ع��P��&6�;vN���f�&�~��3�����*ע�����iB����źѺ]ݺ���:��U����~��2�6����]:�
�!���'��&-�8�2�d8�_ >��C��6I���N�1lT�YZ���_�r>e���j�qvp��v�Ư{����bt��-B��*��ދ�=���&z���H��l���晻�  �  �=�/=l�=�z= =*�=j=�=� =5W =P��<�=�<ń�<C��<T�<�V�<ݛ�<B��<�#�<g�<W��<���<_+�<k�<���<U��<�#�<_�<E��<'��<�	�<R@�<su�<1��<v��<>�<~;�<�h�<���<U��<���<=�<5.�<�N�<Fl�<؆�<���<���<
��<���<���<���<���<���<f��<���<W��<0��<!��<�u�<:R�< )�<D��<���<��<%J�<�<��<2b�<*�<���<�@�<��<�`�<g��<h�<��<�W�<�Ƽ<�0�<	��<,��<N�<��<6�<�>�<���<-ȭ<��<A�<�w�<⪦<�ڤ< �<�0�<|W�<�{�<`��<ܼ�<Fڗ<���<O�<2'�<�=�<YR�<�e�<�w�<ň�<���<���<���<�<�}<p�y<$�u<n�q<��m<�j<J,f<fDb</]^<�vZ<��V<��R<��N<��J<�	G<&,C<�O?<�u;<v�7<h�3<?�/<	(,<#\(<��$<�� <�<{T<)�<��<�A<�
<T�<gc<{��;���;��;���;��;��;v�;Y�;��;�/�;v��;yZ�;[�;sߨ;HŢ;�Ü;?ۖ;��;�U�;久;i7�;��u;��j;Ô`;�\V;UL;�B;��8;�e/;w&;p;�;�\;Y�;t��:o5�:0��:v�:�m�:�:�:}�:��p:s�S:uy7:Bg:{a�90��9疒9C:9��8E����5���f�ϥ�!عO��ǩ��(6��xN���f���~��5������ע�����A����ź�Ѻݺ=�����e���~��1�A��Ə�s9�l�!�e�'��%-���2��c8���=���C�7I���N��lT�aZ�ԡ_�p>e�[�j�^wp�rv�'�{�_����t���B�����}ދ�e����z���H�����t登�  �  �=�/=[�=�z= =-�=j=�=� =-W =@��<�=�<���<2��<7�<�V�<�<'��<�#�<�f�<O��<���<k+�<k�<���<E��<�#�<_�<T��<F��<�	�<g@�<�u�<@��<���<b�<�;�< i�<���<^��<���<Q�<?.�<�N�<"l�<��<���<���<��<���<w��<���<���<���<[��<���<;��<'��<���<�u�<)R�<)�<?��<���<��<0J�<)�<ҵ�<*b�<3�<ӧ�<A�<��<�`�<y��<#h�<��<�W�<Ǽ<�0�<��<3��<-N�<(��<A�<�>�<���<@ȭ<��<$A�<�w�<۪�<�ڤ<�<�0�<^W�<�{�<C��<ȼ�<3ڗ<���<@�<&'�<|=�<MR�<�e�<�w�<҈�<���<~��<���<�<$�}<��y<=�u<��q<��m<j<�,f<�Db<E]^<wZ<��V<��R<��N<��J<�	G<�+C<�O?<v;<��7<��3<'�/<�',<\(<ԓ$<�� <�<XT<�<��<QA<��
<3�<Kc<V��;g��;D��;���;I��;���;�;:Y�;���;$0�;���;�Z�;��;�ߨ;�Ţ;9Ĝ;�ۖ;��;FV�;��;�7�; �u;% k;��`;�[V;[UL;�B;�8;�e/;5&;�;a;#\;>�;���:�3�:l��:��:fk�:��:��:b�:H�p:��S:Iz7:�h:�d�9/��9z��9@G:9R�8�c���-��f��ʥ��ع��P��&6�;vN���f�&�~��3�����*ע�����iB����źѺ]ݺ���:��U����~��2�6����]:�
�!���'��&-�8�2�d8�_ >��C��6I���N�1lT�YZ���_�r>e���j�qvp��v�Ư{����bt��-B��*��ދ�=���&z���H��l���晻�  �  ��=�/=e�=�z= =�=�i=�=�� =W =&��<�=�<���<
��<�<�V�<���<	��<�#�<�f�<6��<���<O+�<�j�<���<T��<�#�<B_�<]��<d��<
�<�@�<�u�<j��<���<�<�;�</i�<��<}��<��<d�<U.�<�N�<4l�<���<~��<߲�<���<x��<U��<b��<���<l��<2��<r��<��< ��<Փ�<�u�<R�<�(�<'��<���<ۊ�<J�<6�<��<Tb�<P�<��<<A�<.��<a�<���<Ph�<��<�W�<7Ǽ<�0�<O��<R��<NN�<5��<f�<�>�<���<Eȭ<��<A�<�w�<Ū�<mڤ<��<0�<.W�<j{�<��<���<	ڗ<v��<&�<'�<`=�<,R�<�e�<�w�<ǈ�<���<���<���<�<N�}<ͷy<��u<�q<
�m<Vj<�,f<�Db<�]^<qwZ<�V<�R<�N<��J<-
G<,C<P?<v;<C�7<F�3<��/<�',<�[(<��$<H� <R<T<��<��<�@<h�
<��< c<��;΋�;Ǆ�;+��;9��;	��;��;�Y�;κ�;�0�;ﺻ;l[�;j�;F�;SƢ;�Ĝ;+ܖ;��;W�;v��;78�;��u;� k;Ε`;Q\V;�UL;xB;�8;�d/;O&;�;E;D[;��;��:�1�:+��:P�:�h�:
�:��:!
�:�p:��S:w7:�e:�g�9N��9k��9T:9�)�8y濷%��;�e�龥��عG��Z��d!6�.pN�u�f���~�2��I��բ�����uA����ź܀Ѻ�ݺØ躾���������3����J���;�7�!�M�'�(-��2�6e8�B>��C�u7I�{�N��lT��Z�R�_� =e���j��up�v���{�6����s���A�����f݋�����Ty��H������晻�  �  �=�/=l�=�z= =#�=�i=�=ܲ =�V =���<F=�<6��<���<��<;V�<N��<���<�#�<�f�< ��<���<@+�<�j�<���<Z��<�#�<I_�<���<���<d
�<�@�<�u�<���<��<��<<�<yi�<��<˾�<Z��<��<p.�<�N�<Hl�<���<x��<��<���<Q��<��<$��<6��<7��<���<!��<���<���<���<Yu�<�Q�<�(�<���<b��<ۊ�<J�<)�<���<Ub�<m�<��<xA�<���<Ia�<���<�h�<d�<OX�<�Ǽ<E1�<���<���<�N�<h��<x�<�>�<Å�<=ȭ<��<A�<�w�<���<5ڤ<��<30�<�V�<{�<Ԝ�<H��<�ٗ<7��<��<�&�<'=�<R�<�e�<�w�<���<���<���<���<À<��}<[�y<�u<s�q<��m<�j<�-f<�Eb<H^^<�wZ<��V<~�R<|�N<�J<2
G<,,C<P?<�u;<Z�7<�3<��/<G',<F[(<�$<�� <�<ES<�<��<^@<ƚ
<h�<b<���;O��;x��;?��;���;
��;��;�Y�;_��;01�;��;G\�;K�;��;�Ǣ;Ɯ;eݖ;��;�W�;���;9�;3�u;�k;��`;�\V;/UL;7B;�8;�c/;&;�;D;�X;:�;��:j,�:;��:��:Ae�:��:��:��:C�p:y�S:�v7:5e:pc�9��9���9=`:9�]�8b	������w�e�N���)�׹:��F��%6�2hN��f�{�~��.��q	��CԢ�]����@����źu�Ѻ�ݺ�����F������
6��������=��!��'�*-�x�2�g8�>��C�a8I�(�N��lT�3Z�ۡ_�7=e���j�Ctp��v�a�{�Z���fr��I@��2��&܋�A���qx���F������噻�  �  2�=�/=�=�z= =�=�i=m=�� =�V =���<�<�<ރ�<O��<q�<�U�<���<S��<?#�<if�<ɨ�<g��<	+�<�j�<���<h��< $�<}_�<ә�<���<�
�<&A�<Yv�<��<m��<C�<_<�<�i�<q��<��<���<��<�.�<�N�<cl�<��<o��<���<���<'��<���<���<���<���<{��<���<r��<D��<K��<�t�<�Q�<}(�<���<<��<���<J�<0�<��<b�<��<a��<�A�<���<�a�<_��<i�<��<�X�<�Ǽ<�1�<<���<�N�<���<��< ?�<څ�<@ȭ<��<�@�<nw�<d��< ڤ<r�<�/�<�V�<�z�<��<껙<`ٗ<���<y�<�&�<�<�<�Q�<Se�<�w�<���<���<ħ�<ܵ�<dÀ<!�}<��y<��u<%�q<i�m<�j<X.f<BFb<_^<�xZ<5�V<�R<��N<��J<�
G<x,C<+P?<�u;<�7<��3<T�/<�&,<�Z(<O�$<�� <�<�R<O�<��<�?<�
<��<b<��;���;���;Ō�;ť�;'��;��;~Z�;w��;�1�;	��;�]�;��;��;�Ȣ;�ǜ;�ޖ;*�;Y�;ɼ�;�9�;ءu;tk;��`;�]V;4UL;�~B;��8;@b/;�&;�;{;SU;O�;U��:h&�:i��:>�:�_�:>��:�:��:��p:-�S:�p7:�c:�c�9���9���9�}:9�82P��Rt����e�q���[�׹��I���6�
\N�7�f��}~��+������Т�/����?����ź��Ѻ=ݺe��J��Ȗ�����^9���s���@��!���'�*--�o�2��h8�>�H�C�:I�:�N�mT��Z���_��;e��j�}rp�4v��{������p���>������ڋ����� w���E�����噻�  �  ?�=�/=��=�z= =�=�i=O=�� =�V =*��<�<�<k��<���<��<jU�<���< ��<�"�<�e�<���</��<�*�<�j�<���<g��< $�<�_�<���<#��<�
�<�A�<�v�<���<���<��<�<�<Tj�<ݕ�<t��<���<�<�.�<	O�<al�<��<g��<���<���<���<���<���<���<n��<��<C��<��<٫�<ג�<�t�<6Q�<#(�<���<��<���<J�<A�<��<�b�<��<���<B�<5��<b�<���<�i�<I�<8Y�<rȼ<#2�<a��<T��<)O�<룴<��</?�<ޅ�<Qȭ<��<�@�<@w�<%��<�٤<�<}/�<0V�<7z�<���<p��<�ؗ<s��<%�<(&�<�<�<�Q�<6e�<�w�<���<���<ʧ�<��<|À<��}<��y<{�u< �q<Y n<�j<?/f<IGb<�_^<{yZ< �V<��R<��N<��J<�
G<�,C<4P?<�u;<�7<u�3<��/<+&,< Z(<��$</� <<�Q<0�<�<�><8�
<��<$a<О�;���;��;O��;ť�;��;[�;[�;��;?3�;L��;_�;>�;��;�ʢ;2ɜ;p��;��;�Z�;��;K;�;��u;=k;�`;X]V;sUL;m~B;��8;�`/;V&;�;H;�R;��;a��:"�:��:P��:;X�:R��:�ܕ:���:�p:��S:�m7:�b:�f�9���9g��9��:94ҡ8^�������}e�bw��i�׹���={���5��NN��tf�Cs~��%��<��w΢������?���źɂѺ�ݺ��躊"��G���ц��;�������D���!�6�'�20-�
�2�l8��>�@�C��:I��N�*mT��Z���_�Y:e�B�j�pp�v�٦{�F���o���<���
���؋�즎�Vu�� D��v���㙻�  �  [�=0=��=�z=	 =��=�i=$=y� =�V =���<<�<��<k��<l�<�T�<��<���<p"�<�e�<A��<���<�*�<�j�<���<r��<@$�<�_�<7��<��<Y�<�A�</w�<��<i��<5�<]=�<�j�<O��<տ�<H��<e�</�<7O�<ul�<��<C��<���<C��<���<Q��<!��<��<���<���<���<{��<e��<Z��<At�<�P�<�'�<H��<���<���<�I�<F�<1��<�b�<	�<���<B�<���<�b�<S��<j�<��<�Y�<�ȼ<�2�<ٖ�<���<�O�<6��<��<Y?�<�<Rȭ<j�<�@�<�v�<䩦<_٤<��</�<�U�<�y�<���<��<nؗ<��<��<�%�<Z<�<KQ�<e�<hw�<���<���<ৄ<B��<�À<m�}<8�y<B�u<��q<9n<�j<?0f<MHb<�`^<_zZ<ДV<h�R<T�N<]�J<cG<�,C<DP?<�u;<��7<%�3<.�/<�%,<QY(<��$<0� <<�P<1�<#�<�=<B�
<�<�`<���;#��;y��;���;z��;��;��;�[�;ɽ�;�4�;���;�`�;��;X�;�̢;˜;R�;��;X\�;���;�<�;�u;�k;f�`;�]V;eUL;*}B;��8;�^/;�&;;�;�;�O;��;���:��:���:���:+P�:��:֕:.��:�p:9�S:j7:y]:f�9���9���9#�:9��8�G��7���Ee��\����׹���k���5�"AN�&gf��g~� �����]ˢ�����:?����źN�Ѻ+ݺl���&��s���F��k?����~���H�K�!�6�'�&4-�d�2��n8�Z	>��C�f<I��N��mT�pZ�џ_��8e���j�Kmp�]v���{�����Tm���:������֋�+����s���B����G♻�  �  ��=*0=��=�z= =��=�i==K� =WV =W��<�;�<v��<���<��<T�<���<��<"�<ae�<��<���<�*�<�j�<���<���<_$�<`�<���<���<��<dB�<�w�<���<���<��<�=�<@k�<���<E��<���<��<O/�<QO�<�l�<���<7��<_��<��<N��<���<���<���<���<��<W��< ��<��<���<�s�<mP�<�'�<��<���<e��<�I�<O�<a��<
c�<^	�<I��<�B�<��<c�<���<�j�<R�<;Z�<}ɼ<!3�<L��<,��<�O�<���<`��<�?�<��<Vȭ<[�<�@�<�v�<���<٤<L�<�.�<GU�<Oy�<��<���<�ח<��<P�<o%�<�;�<Q�<�d�<Iw�<���<̘�<��<a��<Ā<�}<ͺy<�u<��q<@n<�j<51f<(Ib<�a^<W{Z<��V<�R<��N<�J<�G<-C<hP?<�u;<s�7<��3<��/<�$,<�X(<�$<L� <<�O<,�<�<�<<Q�
<<�<�_<(��;=��;���;��;I��;W��;�;X\�;���;T5�;���;)b�;��;<�;D΢;�̜;��;x�;�]�;+��;�=�;+�u;�k;�`;�^V;nUL;�|B;v�8;L]/;o&;Q�;�;�K;D�;Ɣ�:��:���:���:�I�:��:�ϕ:j�:��p:��S:7e7:�[:�f�9���9�Ò9z�:9�k�89^��+M���e�-=��ۀ׹��T]���5�&1N� Zf��Z~���������Ǣ�����'=����ź��Ѻ.ݺ��>,�����N���B�V��q���L�Q�!��'��7-���2��q8�;>�ʥC�>I��N�>nT�Z���_��7e��j�Kkp�
v�U�{�����Lk��M9����� Ջ�#����q���@�����Xᙻ�  �  ��=40=��=�z= =��=i=�= � =(V =���<1;�<��<j��<~�<�S�<��<���<�!�<�d�<���<���<p*�<�j�<���<���<|$�<*`�<͚�<��<"�<�B�<x�<���<U��<3�<?>�<�k�<��<���<���<��</�<gO�<�l�<���<<��<5��<���< ��<���<p��<D��<��<���<���<���<r��<���<js�<P�<3'�<���<���<9��<�I�<J�<s��<*c�<�	�<���<*C�<���<_c�<\��<k�<��<�Z�<�ɼ<�3�<���<���</P�<ޤ�<���<�?�<)��<Qȭ<a�<W@�<�v�<U��<�ؤ<��<;.�<�T�<�x�<���<��<�ח<�<��<%�<�;�<�P�<�d�<-w�<���<Ę�<��<u��<:Ā<z�}<��y<��u<|�q<.n<qj<O2f<Jb<�b^<|Z<i�V<�R<k�N<��J<�G<M-C<eP?<�u;<N�7<[�3<~�/<J$,<�W(<�$<u� <'
<�N<?�<�<�;<l�
<n�<�^<��;���;���;��;��;I��;j�;�\�;޿�;�6�;{»;Rc�;*�;��;Т;�Μ;��;G�;!_�;�;?�;$�u;-	k;��`;V_V;�TL;�|B;�8;\/;�&;�;
;�H;��;-��:c�:?��:2��:"B�:��:{ʕ:��: �p:��S:_7:
\:d�9���9*ʒ9�:9.��8:۸�����-�d���:e׹d��>M��5�w#N�6Pf��M~��������Ţ�܆���<��l�ź��ѺhݺH��v0��N���-��JF�'��n��(P�>�!���'��:-���2��t8�>��C�^?I���N�:nT�DZ���_�	7e�I�j�ip��v�Y�{�Y���si��y7�����DӋ�O���Lp��l?��!��,����  �  ��=P0=��=�z=�=��=hi=�=� =V =���<�:�<���<��<�<�S�<���<W��<_!�<�d�<e��<E��<G*�<mj�<���<���<�$�<]`�<���<M��<X�<C�<ux�<P��<���<��<�>�<
l�<x��<���<(��<$�<�/�<�O�<�l�<��<+��<��<���<���<d��<+��<���<���<M��<���</��<��<��<s�<�O�<'�<���<X��<��<�I�<N�<���<ac�<�	�<ɩ�<mC�<���<�c�<���<fk�<A�<*[�<Sʼ<�3�<��<���<uP�<��<���<�?�<9��<Pȭ<J�<3@�<tv�<"��<~ؤ<��<�-�<rT�<�x�<3��<���<'ח<��<��<�$�<l;�<�P�<qd�<w�<|��<˘�<7��<���<fĀ<�}<�y<z�u<P�q<�n</j< 3f<�Jb<�c^<�|Z<�V<X�R<��N<��J<TG<�-C<vP?<�u;<�7<��3<��/<�#,<hW(<p�$<�� <b	<�M<n�<_�<�:<��
<��<�^<��;h��;��;E��;���;Z��;��;f]�;s��;l7�;9û;�d�;��;)�;�Ѣ;(М;��;r�;�`�;�Å;�?�;��u;}
k;6�`;�_V;�TL;|B;��8;EZ/;�&;��;�;�E;��;j��:;�:��:���:�;�:Dߤ:�ŕ:��:�p:��S:�Z7:XY:�c�9[��9�֒9��:9�ݢ8E�W�����d��	��ZN׹��qA�7�5��N��Cf�G~������¢�~���<����źv�Ѻ� ݺ����3��H�������H�)����7S� �!�y�'��=-���2��v8��>�T�C��@I��N��nT�Z�	�_�J5e���j�>gp�v��{�����'h��6��q���ы������n��>��K��4ߙ��  �  Ǌ=\0=��=�z=�=��=gi=�=� =�U =^��<�:�<R��<���<��<YS�<q��<��<!�<�d�<4��<%��<K*�<\j�<���<���<�$�<|`�<��<���<��<fC�<�x�<���<��<��<?�<El�<Ǘ�<)��<c��<W�<�/�<�O�<�l�< ��<��<��<���<���<1��<���<���<x��<���<*��<ѽ�<ϩ�<��<�r�<�O�<�&�<f��<D��<��<�I�<b�<���<jc�<�	�<���<�C�<	��<&d�<���<�k�<��<�[�<�ʼ<:4�<h��<��<�P�<;��<���<�?�<E��<dȭ<;�<>@�<[v�<�<Aؤ<^�<�-�<(T�<2x�<љ�<]��<�֗<��<U�<�$�<>;�<pP�<ld�<�v�<x��<Ԙ�<)��<���<�Ā<\�}<��y<�u<��q<cn<�j<�3f<�Kb<d^<o}Z<��V<ϲR<\�N<�J<�G<v-C<�P?<�u;<�7<��3<��/<}#,<�V(<�$<:� <�<:M<��<��<X:<;�
<*�<�]<��;҄�;��;��;��;c��;��;�]�;���;88�;Ļ;�e�;z�;o�;�Ң;Iќ;��;N�;�a�;�ą;�@�;�u;Rk;c�`;�_V;AUL;�{B;��8;�Y/;&;��;8;�C;��;E��:���:"��:���:�7�:�ۤ:���:��:��p:��S:�Z7:'W:�g�9���9�ג9~;9��8����o����d������4׹a���6�~�5��N�I9f�H?~���������܄���;����ź��Ѻ� ݺv��27��C���	���J�������NV���!��'��?-���2��x8�'>���C�AI�G�N��nT��Z�n�_��4e��j��ep�,�u�Ø{�����g��l4��S��MЋ�̞���m���<��c��Wޙ��  �  ؊=k0=��=�z=�=��=Si=�=� =�U =5��<e:�<#��<���<��<2S�<A��<���<� �<ed�< ��<��<!*�<Hj�<���<���<�$�<�`�<8��<���<��<�C�<�x�<Ѭ�<1��<��<,?�<vl�<��<G��<���<p�<�/�<�O�<�l�<���<��<��<���<���<��<���<���<I��<���<��<���<���<���<�r�<iO�<�&�<[��<+��<���<�I�<\�<���<�c�<
�<��<�C�<-��<Fd�<&��<�k�<��<�[�<�ʼ<e4�<���<B��<�P�<[��<
��<�?�<X��<Wȭ<*�<@�<Jv�<ߨ�<#ؤ<@�<�-�<�S�<
x�<���<8��<�֗<Q�<*�<i$�<!;�<hP�<Fd�<�v�<i��<֘�<J��<ٶ�<�Ā<��}<̼y<=�u<'�q<�n<Nj<�3f<�Kb<zd^<�}Z<�V<�R<��N<^�J<�G<�-C<�P?<�u;<��7<��3<|�/<K#,<�V(<��$<�� <\<�L<g�<`�<�9<ϔ
<��<�]<���;���;)�;���;���;���;�;7^�;R��;�8�;�Ļ;Cf�;�;�;ZӢ;�ќ;*�;�;Lb�;�ą;8A�;ǭu;Hk;�`;^`V;UL;�zB;��8;�X/;�&;��;S;}B;�;��:���:0��:��:�4�:�ؤ:ؾ�:��:�p:2�S:�U7:U:�e�9'��9�ݒ96;9�'�8ax���N���|d����*׹�~�l2�D�5��N��5f��:~�����햺����򂮺�:����ź݊Ѻ!#ݺ���q8��=�����QL����Ь�/W���!�p�'�IA-���2��y8�	>�ݪC�FBI�'�N�<oT��Z�i�_��3e���j��dp��u��{����Tf���3������ϋ����m���<������ݙ��  �  ��=�-=��=[w=�=Y�=xd=r=(� =�O =��<D,�<r�<b��<H��<�@�<���<���<�
�<�L�<֍�<R��<��<�L�<��<���<��<(<�<!u�<׬�<3��<-�<�K�<�}�<��<���<�	�<5�<?^�<U��<:��<���<���<E
�<�$�<�<�<zQ�<�b�<q�<�{�<܂�<M��<ą�</��<�x�<mk�<�Y�<�C�<�(�<��<���<5��<V��<�S�<m�<;��<��<�B�<;��<���<�5�<��<d�< ��<�y�<���<Jx�<��<�_�<?˺<i1�<Z��<G�<=E�<��<.�<_.�<]s�<O��<6�<�*�<L`�<���<(¢<��<R�<�?�<Od�<톙<���<%ƕ<�<2��<��<�/�<�F�<=\�<�p�<���<	��<p��<��<P�}<g�y<��u<_�q<�n<�%j<WCf<�`b<^<��Z<½V<��R<� O<$K<IG<�oC<��?<��;<�7<� 4<�S0<��,<n�(<� %<.B!<�<��<b"<vw<G�<3<�<�<| <���;��;}�;
1�;rg�;���;�	�;�v�;���;��;07�;��;�̪;﹤;Y��;�٘;�;�Z�;g��;�<�;�y;�o;��d;�QZ;�AP;�aF;^�<;`-3;��);� ;��;f�;�=;F��:(��:z�:Yh�:ל�:��:4қ:wʌ: |:#�^:%B:��%:L�	:�M�9���9�z_9Dw�8Ð27Vź�O�D�����u�ȹ�����h��1/�N�G�l6`��{x�?M��5L��\:�����W췺ʱú0kϺ6ۺ
��;]�����W���|
��8��������T!�2'���,��Q2��7�2�=��9C���H�dxN�<T�Q�Y��T_���d���j� 2p���u��q{�.����Y���*��q���2͋�����:q��AD��.���왻�  �  ��=�-=��=bw=�=K�=xd=p=2� =�O =��<T,�<r�<|��<_��<�@�<���<���<�
�<�L�<��<K��<��<kL�<��<���<��<3<�<%u�<Ԭ�<'��<�<�K�<�}�<	��<���<�	�<�4�<-^�<E��<1��<���<���<I
�<�$�<�<�<`Q�<�b�<q�<�{�<���<O��<҅�<A��<�x�<�k�<	Z�<�C�<�(�<��<���<L��<U��<�S�<_�< ��<���<�B�<9��<���<�5�<��<�c�<���<�y�<���<#x�<��<�_�<$˺<Z1�<M��<A�<EE�<���<+�<g.�<`s�<3��<2�<�*�<S`�<В�<+¢<��<^�<�?�<ld�<��<���<5ƕ<�<2��<��<�/�<�F�<$\�<zp�<˃�<��<{��<"��<[�}<W�y<��u<(�q<�n<�%j<	Cf<�`b<�~^<ŝZ<��V<u�R<� O<$K< IG<�oC<��?<��;<��7<� 4<�S0<�,<o�(<� %<NB!<-�<��<�"<�w<b�<,3<!�<�<3| <y��;y��;�;�0�;�g�;���;�	�;
w�;���;׌�;�6�;���;�̪;���;���;�٘;��;NZ�;+��;�<�;]�y;o;��d;-RZ;BP;�`F;¯<;-3;w�);Ӱ ;�;��;u>;��:Z��:0|�:3i�:���:��:Nқ:�ˌ:��{:��^:�B:;�%:�	:�O�9&��9_9��8�527Ӻ��D�F����ȹ����-l��2/���G�18`�c}x��M���K���9������뷺��ú�lϺwۺ����\�����<��2|
�T8��������S!�� '�q�,�_Q2�
�7�s�=��9C���H�)yN��T�׵Y��T_�Y�d���j��1p���u�@r{�����Z���*�����b͋�4����q��yD��S���왻�  �  v�=�-=��=_w=�=X�=�d=w=?� =�O =1��<u,�<7r�<���<s��<�@�<���<��<�
�<�L�<���<]��<��<~L�<��<���<��<<�<u�<���<
��<�<yK�<�}�<��<���<�	�<�4�<^�<0��<��<���<���<2
�<�$�<�<�<iQ�<
c�<8q�<�{�<��<b��<��<b��<�x�<�k�< Z�<�C�<�(�<	�<���<g��<b��<�S�<��<&��<��<�B�<!��<���<�5�<���<�c�<���<�y�<���<x�<��<�_�<˺<=1�<2��<!�<&E�<q��<�<Y.�<^s�<?��<Y�<�*�<d`�<璤<@¢<��<|�<�?�<}d�<&��<���<Uƕ<(�<F��<��<�/�<�F�<A\�<�p�<Ń�<���<j��<��<,�}<�y<b�u<��q<Bn<�%j<�Bf<�`b<�~^<��Z<t�V<:�R<f O<�#K<�HG<�oC<��?<��;<	�7<2!4<�S0<�,<��(<%<�B!<e�<�<�"<�w<��<t3<X�<�<b| <���;.��;X�;1�;�g�;]��;�	�;�v�;t��;k��;�6�;*��;`̪;G��;X��;�٘;I�;�Y�;ᾇ;b<�;��y;o;�d;�QZ;�AP;QaF;�<;7.3;��);�� ;��;��;�?;���:���:�}�:�j�:͟�:��:�ӛ:�͌:�|:��^:vB:P�%:��	:VK�9߱�9�r_9�k�8617庸��D�iÕ���ȹg���o�6/�}�G��;`�u�x�aO��fM��;������췺��úlϺ�ۺF�溔[�s������"{
�_7���)���R!� '�p�,�~P2�k�7���=�_9C���H�IxN��T��Y�8U_���d�w�j��2p���u��r{�
����Z��7+��y����͋�����!r���D�����M홻�  �  m�=�-=��=Xw=�=\�=�d=�=N� =�O =e��<�,�<|r�<׷�<���<$A�< ��<C��<�
�<�L�<��<}��<��<�L�<��<���<��<<�<�t�<���<���<��<QK�<@}�<���<s��<k	�<�4�<�]�<��<��<���<���<5
�<�$�<�<�<Q�< c�<@q�<|�<-��<���<��<���<�x�<�k�<[Z�<8D�<7)�<+	�<��<���<���<�S�<v�<<��<��<�B�<&��<r��<�5�<���<�c�<���<�y�<~��<�w�<K�<>_�<�ʺ<�0�<	��<��<E�<Y��<�<V.�<Ts�<O��<K�<�*�<�`�<��<v¢<��<��<�?�<�d�<b��<�<�ƕ<Y�<���<
�<$0�<�F�<C\�<�p�<���<��<`��<���<�}<ͮy<��u<��q<�n<�$j<]Bf<�_b<E~^<)�Z<��V<��R< O<�#K<�HG<�oC<��?<��;<�7<%!4<1T0<\�,<	�(<n%<�B!<�<��<P#<kx<'�<�3<˚<Q<�| <Z��;��;��;&1�;�g�;���;w	�;av�;��;ዽ;�5�;���;[˪;/��;���;Pؘ;��;�X�;5��;�;�;��y;�o;9�d;�QZ;�AP;bF;��<;�.3;^�);�� ;��;3�;�A;g��:���:���:ko�:��:x�:Vכ:�ό:&|:��^:�B:M�%:I�	:M�9���9�h_9�L�8�J07���;E��˕�<�ȹ�����w��?/�1�G��C`��x�\Q���N��J<��M���췺�ú�jϺ�ۺ���;Y����ǹ��y
�^5������Q!���&�˧,��N2���7���=��7C���H�;xN�T�s�Y�U_�4�d��j��3p�$�u��t{�Ԋ��N[��z,��`����΋�}����r���E��d���홻�  �  \�=�-=��=Tw=�=h�=�d=�=b� =�O =���<�,�<�r�<��<��<aA�<H��<���<.�<M�<C��<���<�<�L�<��<��<��<�;�<�t�<Z��<���<��<K�<}�<d��<0��<"	�<r4�<�]�<΄�<���<]��<���<
�<�$�<�<�<�Q�<c�<aq�<?|�<Y��<܆�<W��<ށ�<-y�<&l�<�Z�<sD�<t)�<g	�<I��<���<���<T�<��<L��<ݏ�<�B�<���<I��<{5�<|��<{c�<;��<My�<3��<|w�<�<�^�<�ʺ<�0�<Ց�<��<�D�<(��<��<C.�<Ps�<a��<a�<�*�<�`�<:��<�¢</�<��<0@�<e�<���<3��<�ƕ<��<���<3�<U0�<�F�<\\�<�p�<���<땄<2��<з�<z�}<w�y<��u<��q<kn<a$j<�Af<`_b<�}^<��Z<|�V<��R<��N<]#K<HG<�oC<��?<��;<J�7<V!4<�T0<��,<v�(<�%<~C!<��< �<�#<�x<��<Z4<W�<�<
} <"��;���;�;91�;dg�;��;��;�u�;��;M��;�4�;���;�ʪ;0��;���;=ט;��;�W�;o��;;�;L�y;�o;�d;eQZ;�AP;�bF;u�<;�/3;��);� ;��;*�;�C;:��:��:/��:<s�:��:a �:�ۛ:�Ҍ:�|:Z�^:� B:��%:�	:�H�9Z��9�V_92!�8Tl.7�C���;E��ڕ���ȹ��,��-G/�Q�G�LL`�Ҋx�mU��IQ��?�����h��úoiϺ�ۺѻ溒V���������w
�63�	�����O!���&���,�M2���7�i�=�x6C���H�uwN��T���Y��U_���d�%�j�y5p�{�u��v{����D\���-��g���Ћ�u���t���F������  �  H�=w-=|�=Xw=�=p�=�d=�=�� =P =���<=-�<s�<u��<Z��<�A�<���<���<p�<]M�<z��<���<=�<�L�<��<���<��<�;�<�t�<��<j��<M�<�J�<�|�<
��<���<��<4�<I]�<���<p��<+��<c��<�	�<�$�<�<�<�Q�<Cc�<�q�<V|�<���<��<���<1��<�y�<�l�<�Z�<�D�<�)�<�	�<x��<��<׉�<"T�<��<<��<��<lB�<���<&��<F5�<1��<-c�<���<�x�<���<w�<��<�^�<!ʺ<m0�<��<r�<�D�<	��<��<8.�<Us�<W��<��<�*�<�`�<~��<�¢<��<N�<�@�<be�<���<���<!Ǖ<��<���<w�<h0�<G�<x\�<�p�<���<ו�<!��<���<�}<ԭy<�u<d�q<�n<�#j<Af<�^b<�|^<��Z<�V<��R<0�N<
#K<[HG<loC<��?<��;<k�7<�!4<�T0<6�,<��(<�%<.D!<1�<��<�$<�y<l�<5<�<W	<�} <���;c��;=�;o1�;g�;ݮ�;��;Gu�;:��;$��;�3�;-�;-ɪ;ߵ�;'��;֘;G
�;�V�;o��;:�;ءy;� o;f�d;�PZ;
BP;obF;��<;�03;��);_� ;D�;��;5F;���:��:��:�x�:H��:�%�:�ޛ:�֌:�|:V�^:�&B:q�%:v�	:�D�9���9�G_9���8(A,7����XE�����>�ȹb#������Q/�s�G�`S`���x�QY��
T���@��$����F�ú�iϺ�ۺ��溏S�q���ҵ�)u
��0�<���� L!���&��,��J2��7�I�=��5C���H��vN��T�U�Y�_V_�0�d�U�j�%7p��u�vx{�����]���.������Nы� ���.u���G��H����  �  +�=j-=n�=Tw==v�=�d=�=�� =5P =;��<�-�<ls�<ո�<���<$B�<��<-��<��<�M�<Î�<���<b�<�L�<.��<n��<��<�;�<mt�<��<��<��<\J�<U|�<���<n��<��<�3�<�\�<(��<B��< ��<,��<�	�<�$�<�<�<�Q�<Wc�<�q�<�|�<��<O��<���<}��<�y�<�l�<U[�<.E�<*�<
�<���<6��<��<HT�<��<D��<��<QB�<���<��<5�<��<�b�<���<zx�<���<�v�<;�<E^�<�ɺ<0�<��<P�<oD�<ݖ�<��<.�<`s�<\��<��<+�<a�<���<2â<��<��<�@�<�e�<\��<娗<oǕ<4�<1��<��<�0�<BG�<�\�<�p�<���<���<��<r��<Ɏ}<R�y<H�u<��q<�n<#j<D@f<
^b<B|^<W�Z<K�V<Y�R<��N<�"K<"HG<3oC<~�?<��;<��7<"4<-U0<Ƌ,<p�(<$%<�D!<�<��<V%<�z<�<�5<~�<�	< ~ <f��;��;�;�1�;Qg�;���;.�;�t�;���;;�2�;�;�Ǫ;���;���;�Ԙ;��;�U�;���;[9�;��y;"�n;�d;CPZ;�BP;�bF;��<;@23;��);и ;b�;��;�H;M��:���:���:F�:N��:+�:��:zی:�|:��^:*B:�%:��	:B?�9���9�._9��8��*7W컸~E������ȹ�;��A��K\/���G��\`�ßx��Z��cW���B��2��ﷺ0�úiϺ�ۺ���O��������r
�!.����!��2I!�&�&���,�H2��7���=��3C�0�H�/vN�T�T�Y�9W_���d��j�>8p��u�Z{{�U���Z_��*0������ҋ�p���iv��I��p��$��  �  �=V-=i�=Lw==��=�d=�=�� =\P =���<�-�<�s�<.��<��<yB�<G��<z��<�<�M�<��<'��<v�<�L�<*��<c��<��<};�<-t�<���<���<��<J�<�{�<T��<��<�<Z3�<�\�<��<��<���<���<�	�<�$�<�<�<�Q�<ec�<�q�<�|�<��<���<H��<Ђ�<;z�<8m�<�[�<~E�<e*�<S
�<��<X��<F��<sT�<��<V��<ُ�<?B�<���<���<�4�<���<}b�<O��<"x�<��<Ov�<��<�]�<rɺ<�/�<א�<��<&D�<���<��<.�<Qs�<n��<��<D+�<Ba�<瓤<�â<�<��<=A�<f�<���<;��<�Ǖ<��<���<��<�0�<bG�<�\�<�p�<���<���<概<?��<7�}<߬y<��u<�q<:n<I"j<�?f<E]b<�{^<��Z<��V<��R<_�N<)"K<�GG<oC<]�?<��;<��7<;"4<�U0<�,<�(<�%<{E!<��<c�<2&<6{<��<d6<E�<Y
<u~ <]��;w��;��;�1�;<g�;~��;��;�s�;���;��;�1�;��;�ƪ;3��;[��;bӘ;��;�T�;��;j8�;��y;��n;1�d;PZ;BP;�cF;D�<;�33;��);ʹ ;H�;��;ZK;���:���:З�:���:���:�/�:��:�݌:h |:��^:�+B:��%:w�	::<�9��9�_9�~�8��(7�.��էE������ȹ�Q��w��ih/�n�G�zg`��x��_���[��E��a ���ﷺʰú�gϺ�ۺ�溚L�u������,p
�E+�t����iF!�q�&��,�}E2���7� �=�N2C�6�H�yuN�T��Y��W_��d���j��:p���u��}{������`���1�����5ԋ�å���w��;J��W��=��  �  �=?-=c�=Kw==��=�d=�=Ӭ =�P =���</.�<'t�<��<y��<�B�<���<���<U�<#N�<��<M��<��<�L�<��<k��<s�<U;�<t�<r��<���<Z�<�I�<�{�<���<���<��<	3�<T\�<���<���<���<���<�	�<�$�<�<�<�Q�<zc�<�q�<�|�<E��<���<���<;��<�z�<�m�<\�<�E�<�*�<�
�<\��<���<p��<�T�<��<`��<ɏ�<EB�<o��<���<�4�<j��<Db�<���<�w�<���<�u�<t�<z]�<ɺ<c/�<���<��<
D�<���<s�<.�<@s�<��<��<b+�<ra�<1��<�â<X�<`�<�A�<{f�<��<���<ȕ<��<���<�<	1�<xG�<�\�<�p�<���<���<���<-��<ō}<T�y<,�u<t�q<�n<�!j<�>f<�\b<�z^<��Z<�V<[�R<��N<�!K<oGG<oC<V�?<��;<��7<^"4<�U0<z�,<��(<O%< F!<f�<�<�&<�{<��<�6<Ν<<�~ <
��;���;k�;�1�;tg�;��;�;ts�;���;B��;q0�;��;@Ū;˱�;��;Ҙ;��;\S�;4��;[7�;Y�y;H�n;ɍd;`PZ;�AP;�cF; �<;w43;-�);ڻ ;��;��;�N;��:���:���:���:���:r3�:��:�:&&|:�^:�.B:��%:�	:�>�9ٌ�9�_9�[�8E�&7a����E�4��2	ɹ�h��c���s/�	H��q`�v�x�6d���\���G���"��ﷺ��úCfϺ�ۺ��iI�������;n
��'������C!���&�?�,��C2�	�7�4�=��0C���H��tN�T��Y��W_���d�K�j�Q<p� �u��{������a��03��,���Ջ����y��bK��^��A��  �  �=3-=W�=Hw==��=�d=
	=� =�P =	��<x.�<et�<ǹ�<���<C�<��<
��<��<PN�<O��<q��<��<�L�<%��<]��<[�<:;�<�s�<I��<e��<�<vI�<_{�<���<o��<��<�2�<\�<g��<���<`��<���<y	�<�$�<�<�<�Q�<�c�<r�<!}�<���<'��<ć�<y��<�z�<�m�<O\�<F�<+�<�
�<���<Ժ�<���<�T�<�<m��<Ǐ�<+B�<T��<p��<f4�<4��<�a�<���<�w�<u��<�u�<+�<7]�<�Ⱥ< /�<X��<~�<�C�<\��<Y�<�-�<?s�<���<��<�+�<�a�<`��<Ģ<��<��<�A�<�f�<O��<ҩ�<`ȕ< �<���<Y�<-1�<�G�<�\�<�p�<���<���<���<���<w�}<�y<��u<��q<n<!j<N>f<\b<^z^<y�Z<��V<��R<��N<�!K<>GG<�nC<I�?<��;<�7<�"4<9V0<�,<�(<�%<�F!<�<��<}'<m|<5�<�7<D�<g<X <���;���;��;�1�;Qg�;ͭ�;��;�r�;J��;p��;�/�;��;VĪ;ڰ�;촞;-ј;��;hR�;.��;�6�;	�y;�n;�d;�OZ;�AP;�dF;i�<;�53;��);� ;a�;�;�P;է�:���:ˡ�:ʍ�:rº:�7�:��:��:�+|:��^:E4B:��%:>�	:�9�9��9��^9-)�8�%7������E�iD���ɹ�{�����v{/��H��y`�8�x��f���_���I��R$���U�ú�dϺ�ۺͯ�xF�x������k
�&�������A!���&��,��A2���7�I�=��/C�+�H��sN��T��Y�gX_�X�d���j��=p���u�ǁ{�����c��'4��`���֋�'���z��_L��/�����  �  ܇=7-=Q�=Ew==��=�d=	=� =�P =I��<�.�<�t�<��<���<]C�<��<@��<��<wN�<s��<���<��<�L�<3��<K��<[�<8;�<�s�<*��<*��<��<@I�<{�<x��<,��<@�<�2�<�[�<-��<e��<:��<���<�	�<z$�<�<�<�Q�<�c�<.r�<:}�<���<J��<��<���<{�<n�<�\�<^F�<++�<�<���<��<���<�T�<�<e��<Ώ�<B�<]��<Z��<:4�<��<�a�<���<<w�<(��<Xu�<��<�\�<�Ⱥ<�.�<��<\�<�C�<R��<Z�<�-�<Ks�<���<��<�+�<�a�<���</Ģ<��<��< B�<�f�<���<��<�ȕ<A�<# �<{�<?1�<�G�<�\�<�p�<���<���<���<ݶ�<1�}<��y<?�u<��q<~n<� j<�=f<�[b<�y^<�Z<1�V<��R<F�N<O!K<MGG<�nC<<�?< �;<�7<�"4<\V0<;�,<T�(<M%<G!<Y�<B�<�'<}<��<	8<��<�<� <��;���;��;:2�;g�;߭�;��;r�;���;���;�.�;��;@ê;���;�;&И;��;�Q�;S��;$6�;�y;_�n;��d;-OZ;=BP;�dF;1�<;�63;Y�);�� ;��;"�;�Q;٬�:	�:Х�:��:�ĺ:-<�:m�:��:F/|:��^:)3B:�%:��	:�3�9:��9��^9h �8�1$7�Ἰ�F�dU���*ɹI��� ����/��H�=`�|�x��h���b��4J���#��a�S�ú|eϺ�ۺ���DD�<���f���i
��$�?��-��-?!���&���,��?2���7�>�=�D/C���H�tN��T�/�Y��X_��d�˜j��>p��u�q�{�����d��5�����׋�9����z��-M�����^��  �  Շ=!-=E�=Bw==��= e="	=� =�P =`��<�.�<�t�<*��<��<tC�<7��<\��<��<�N�<���<���<��<M�<7��<B��<=�<;�<�s�<��<��<��<I�<�z�<]��<��<&�<c2�<�[�<��<K��<)��<���<\	�<p$�<�<�<�Q�<�c�<Er�<T}�<Ä�<a��<!��<���<0{�<-n�<�\�<tF�<M+�<-�<���<��<ˊ�<�T�<�<s��<Џ�<B�<2��<<��<(4�<���<�a�<_��<w�<��<@u�<��<�\�<lȺ<�.�<��<?�<�C�<+��<5�<�-�<Ls�<���<��<�+�<�a�<���<DĢ<��<��<5B�<g�<���</��<�ȕ<W�<A �<��<^1�<�G�<�\�<�p�<���<t��<|��<Ͷ�<�}<d�y<	�u<P�q<Cn<T j<�=f<K[b<�y^<ԘZ<��V<Y�R<�N<0!K<�FG<�nC</�?<�;</�7<�"4<�V0<i�,<��(<}%<OG!<��<n�<-(<D}<��<C8<�<�<� <|��; ��;+�;U2�;g�;p��;2�;�q�;��;O��;x.�;i�;�ª;���;���;�Ϙ;!�;UQ�;	��;�5�;q�y;��n;H�d;�NZ;QBP;�dF;ʶ<;T73;2�);�� ;H�;��;�R;y��:��:z��:o��:�ƺ:�=�:���:��:�2|:��^:�5B:�%:�	:�1�9��9��^9=��8/Z#7�����F��]���0ɹ����`����/��H���`�տx�lj���c��wL��&����'�ú/dϺuۺԬ溩B�S������i
��#����O��w>!���&�͖,�?2���7�v�=�P.C���H�jsN�LT�V�Y��Y_�h�d�Q�j�W?p���u�E�{�7���d���5�����؋�����V{���M��T �����  �  ׇ=!-=S�=Hw=
=��=�d=!	=� =�P =n��<�.�<�t�<8��<6��<{C�<I��<u��<��<�N�<���<���<��< M�<(��<X��<V�<;�<�s�<���<��<��<I�<�z�<>��<���<�<W2�<�[�<��<8��<#��<���<a	�<�$�<�<�<�Q�<�c�<9r�<I}�<Ʉ�<l��<0��<փ�<6{�<Nn�<�\�<xF�<f+�<<�<���<��<���<�T�<�<j��<���<!B�<;��<F��<&4�<���<�a�<N��<
w�<���<u�<��<�\�<YȺ<�.�<���<$�<�C�<1��<K�<�-�<:s�<���<��<�+�<�a�<���<TĢ<�<��<9B�<6g�<É�<8��<�ȕ<e�<M �<��<\1�<�G�<�\�<�p�<���<���<��<Ӷ�<�}<X�y<�u<0�q<,n<" j<e=f<[b<�y^<��Z<�V<U�R<��N<8!K<�FG<�nC<D�?<��;<'�7<�"4<�V0<e�,<��(<�%<�G!<��<��<|(<T}<��<x8<�<<� <l��;���;�;2�;^g�;֭�;C�;r�;��;N��;W.�;(�;�ª;��;3��;xϘ;��;Q�;���;{5�;I�y;��n;u�d;�OZ;BP;�dF;�<;�63;��);*� ;��;z�;�S;Ԯ�:��:ʩ�:���:bȺ:�>�:l��:��:�0|:t�^:76B:�%:P�	:�8�9���9F�^9>��8��"7*���{F��`���4ɹ5������c�/��H�S�`�I�x�l��ec��
L���$��X�;�ú�dϺ�ۺc��zC�����2��nh
�8#�l�����=!�|�&��,��>2�B�7�t�=�c.C�W�H�lsN��T� �Y��X_�W�d��j��?p���u�\�{�x����d���5��-���؋�ԩ���{���M��] ������  �  Շ=!-=E�=Bw==��= e="	=� =�P =`��<�.�<�t�<*��<��<tC�<7��<\��<��<�N�<���<���<��<M�<7��<B��<=�<;�<�s�<��<��<��<I�<�z�<]��<��<&�<c2�<�[�<��<K��<)��<���<\	�<p$�<�<�<�Q�<�c�<Er�<T}�<Ä�<a��<!��<���<0{�<-n�<�\�<tF�<M+�<-�<���<��<ˊ�<�T�<�<s��<Џ�<B�<2��<<��<(4�<���<�a�<_��<w�<��<@u�<��<�\�<lȺ<�.�<��<?�<�C�<+��<5�<�-�<Ls�<���<��<�+�<�a�<���<DĢ<��<��<5B�<g�<���</��<�ȕ<W�<A �<��<^1�<�G�<�\�<�p�<���<t��<|��<Ͷ�<�}<d�y<	�u<P�q<Cn<T j<�=f<K[b<�y^<ԘZ<��V<Y�R<�N<0!K<�FG<�nC</�?<�;</�7<�"4<�V0<i�,<��(<}%<OG!<��<n�<-(<D}<��<C8<�<�<� <|��; ��;+�;U2�;g�;p��;2�;�q�;��;O��;x.�;i�;�ª;���;���;�Ϙ;!�;UQ�;	��;�5�;q�y;��n;G�d;�NZ;QBP;�dF;ʶ<;T73;2�);�� ;H�;��;�R;y��:��:z��:o��:�ƺ:�=�:���:��:�2|:��^:�5B:�%:�	:�1�9��9��^9=��8/Z#7�����F��]���0ɹ����`����/��H���`�տx�lj���c��wL��&����'�ú/dϺuۺԬ溩B�S������i
��#����O��w>!���&�͖,�?2���7�v�=�P.C���H�jsN�LT�V�Y��Y_�h�d�Q�j�W?p���u�E�{�7���d���5�����؋�����V{���M��T �����  �  ܇=7-=Q�=Ew==��=�d=	=� =�P =I��<�.�<�t�<��<���<]C�<��<@��<��<wN�<s��<���<��<�L�<3��<K��<[�<8;�<�s�<*��<*��<��<@I�<{�<x��<,��<@�<�2�<�[�<-��<e��<:��<���<�	�<z$�<�<�<�Q�<�c�<.r�<:}�<���<J��<��<���<{�<n�<�\�<^F�<++�<�<���<��<���<�T�<�<e��<Ώ�<B�<]��<Z��<:4�<��<�a�<���<<w�<(��<Xu�<��<�\�<�Ⱥ<�.�<��<\�<�C�<R��<Z�<�-�<Ks�<���<��<�+�<�a�<���</Ģ<��<��< B�<�f�<���<��<�ȕ<A�<# �<{�<?1�<�G�<�\�<�p�<���<���<���<ݶ�<1�}<��y<?�u<��q<~n<� j<�=f<�[b<�y^<�Z<1�V<��R<F�N<O!K<MGG<�nC<<�?< �;<�7<�"4<\V0<;�,<T�(<N%<G!<Y�<B�<�'<}<��<	8<��<�<� <��;���;��;:2�;g�;߭�;��;r�;���;���;�.�;��;@ê;���;�;&И;��;�Q�;S��;$6�;�y;_�n;��d;-OZ;=BP;�dF;1�<;�63;Y�);�� ;��;"�;�Q;٬�:	�:Х�:��:�ĺ:-<�:m�:��:F/|:��^:)3B:�%:��	:�3�9:��9��^9h �8�1$7�Ἰ�F�dU���*ɹI��� ����/��H�=`�|�x��h���b��4J���#��a�S�ú|eϺ�ۺ���DD�<���f���i
��$�?��-��-?!���&���,��?2���7�>�=�D/C���H�tN��T�/�Y��X_��d�˜j��>p��u�q�{�����d��5�����׋�9����z��-M�����^��  �  �=3-=W�=Hw==��=�d=
	=� =�P =	��<x.�<et�<ǹ�<���<C�<��<
��<��<PN�<O��<q��<��<�L�<%��<]��<[�<:;�<�s�<I��<e��<�<vI�<_{�<���<o��<��<�2�<\�<g��<���<`��<���<y	�<�$�<�<�<�Q�<�c�<r�<!}�<���<'��<ć�<y��<�z�<�m�<O\�<F�<+�<�
�<���<Ժ�<���<�T�<�<m��<Ǐ�<+B�<T��<p��<f4�<4��<�a�<���<�w�<u��<�u�<+�<7]�<�Ⱥ< /�<X��<~�<�C�<\��<Y�<�-�<?s�<���<��<�+�<�a�<`��<Ģ<��<��<�A�<�f�<O��<ҩ�<`ȕ< �<���<Y�<-1�<�G�<�\�<�p�<���<���<���<���<w�}<�y<��u<��q<n<!j<N>f<\b<^z^<y�Z<��V<��R<��N<�!K<>GG<�nC<I�?<��;<�7<�"4<9V0<�,<�(<�%<�F!<�<��<}'<m|<5�<�7<D�<g<X <���;���;��;�1�;Qg�;ͭ�;��;�r�;I��;o��;�/�;��;VĪ;ڰ�;촞;-ј;��;hR�;.��;�6�;	�y;�n;�d;�OZ;�AP;�dF;i�<;�53;��);� ;a�;�;�P;է�:���:ˡ�:ʍ�:rº:�7�:��:��:�+|:��^:E4B:��%:>�	:�9�9��9��^9-)�8�%7������E�iD���ɹ�{�����v{/��H��y`�8�x��f���_���I��R$���U�ú�dϺ�ۺͯ�xF�x������k
�&�������A!���&��,��A2���7�I�=��/C�+�H��sN��T��Y�gX_�X�d���j��=p���u�ǁ{�����c��'4��`���֋�'���z��_L��/�����  �  �=?-=c�=Kw==��=�d=�=Ӭ =�P =���</.�<'t�<��<y��<�B�<���<���<U�<#N�<��<M��<��<�L�<��<k��<s�<U;�<t�<r��<���<Z�<�I�<�{�<���<���<��<	3�<T\�<���<���<���<���<�	�<�$�<�<�<�Q�<zc�<�q�<�|�<E��<���<���<;��<�z�<�m�<\�<�E�<�*�<�
�<\��<���<p��<�T�<��<`��<ɏ�<EB�<o��<���<�4�<j��<Db�<���<�w�<���<�u�<t�<z]�<ɺ<c/�<���<��<
D�<���<s�<.�<@s�<��<��<b+�<ra�<1��<�â<X�<`�<�A�<{f�<��<���<ȕ<��<���<�<1�<xG�<�\�<�p�<���<���<���<-��<ō}<T�y<,�u<t�q<�n<�!j<�>f<�\b<�z^<��Z<�V<[�R<��N<�!K<oGG<oC<V�?<��;<��7<^"4<�U0<z�,<��(<O%< F!<f�<�<�&<�{<��<�6<Ν<<�~ <
��;���;k�;�1�;tg�;��;�;ts�;���;B��;q0�;��;@Ū;˱�;��;Ҙ;��;[S�;4��;[7�;Y�y;H�n;ɍd;`PZ;�AP;�cF; �<;w43;-�);ڻ ;��;��;�N;��:���:���:���:���:r3�:��:�:&&|:�^:�.B:��%:�	:�>�9ٌ�9�_9�[�8E�&7a����E�4��2	ɹ�h��c���s/�	H��q`�v�x�6d���\���G���"��ﷺ��úCfϺ�ۺ��iI�������;n
��'������C!���&�?�,��C2�	�7�4�=��0C���H��tN�T��Y��W_���d�K�j�Q<p� �u��{������a��03��,���Ջ����y��bK��^��A��  �  �=V-=i�=Lw==��=�d=�=�� =\P =���<�-�<�s�<.��<��<yB�<G��<z��<�<�M�<��<'��<v�<�L�<*��<c��<��<};�<-t�<���<���<��<J�<�{�<T��<��<�<Z3�<�\�<��<��<���<���<�	�<�$�<�<�<�Q�<ec�<�q�<�|�<��<���<H��<Ђ�<;z�<8m�<�[�<~E�<e*�<S
�<��<X��<F��<sT�<��<V��<ُ�<?B�<���<���<�4�<���<}b�<O��<"x�<��<Ov�<��<�]�<rɺ<�/�<א�<��<&D�<���<��<.�<Qs�<n��<��<D+�<Ba�<瓤<�â<�<��<=A�<f�<���<;��<�Ǖ<��<���<��<�0�<bG�<�\�<�p�<���<���<概<?��<7�}<߬y<��u<�q<:n<I"j<�?f<E]b<�{^<��Z<��V<��R<_�N<)"K<�GG<oC<]�?<��;<��7<;"4<�U0<�,<�(<�%<{E!<��<c�<2&<6{<��<d6<E�<Y
<u~ <]��;w��;��;�1�;<g�;~��;��;�s�;���;��;�1�;��;�ƪ;3��;[��;bӘ;��;�T�;��;i8�;��y;��n;1�d;PZ;BP;�cF;D�<;�33;��);ʹ ;H�;��;ZK;���:���:З�:���:���:�/�:��:�݌:h |:��^:�+B:��%:w�	::<�9��9�_9�~�8��(7�.��էE������ȹ�Q��w��ih/�n�G�zg`��x��_���[��E��a ���ﷺʰú�gϺ�ۺ�溚L�u������,p
�E+�t����iF!�q�&��,�}E2���7� �=�N2C�6�H�yuN�T��Y��W_��d���j��:p���u��}{������`���1�����5ԋ�å���w��;J��W��=��  �  +�=j-=n�=Tw==v�=�d=�=�� =5P =;��<�-�<ls�<ո�<���<$B�<��<-��<��<�M�<Î�<���<b�<�L�<.��<n��<��<�;�<mt�<��<��<��<\J�<U|�<���<n��<��<�3�<�\�<(��<B��< ��<,��<�	�<�$�<�<�<�Q�<Wc�<�q�<�|�<��<O��<���<}��<�y�<�l�<U[�<.E�<*�<
�<���<6��<��<HT�<��<D��<��<QB�<���<��<5�<��<�b�<���<zx�<���<�v�<;�<E^�<�ɺ<0�<��<P�<oD�<ޖ�<��<.�<`s�<\��<��<+�<a�<���<2â<��<��<�@�<�e�<\��<娗<oǕ<4�<0��<��<�0�<BG�<�\�<�p�<���<���<��<r��<Ɏ}<R�y<H�u<��q<�n<#j<D@f<
^b<B|^<W�Z<K�V<Y�R<��N<�"K<"HG<3oC<~�?<��;<��7<"4<-U0<Ƌ,<p�(<$%<�D!<�<��<V%<�z<�<�5<~�<�	< ~ <f��;��;�;�1�;Qg�;���;-�;�t�;���;;�2�;�;�Ǫ;���;���;�Ԙ;��;�U�;���;Z9�;��y;"�n;�d;CPZ;�BP;�bF;��<;@23;��);и ;b�;��;�H;M��:���:���:F�:N��:+�:��:zی:�|:��^:*B:�%:��	:B?�9���9�._9��8��*7W컸~E������ȹ�;��A��K\/���G��\`�ßx��Z��cW���B��2��ﷺ0�úiϺ�ۺ���O��������r
�!.����!��2I!�&�&���,�H2��7���=��3C�0�H�/vN�T�T�Y�9W_���d��j�>8p��u�Z{{�U���Z_��*0������ҋ�p���iv��I��p��$��  �  H�=w-=|�=Xw=�=p�=�d=�=�� =P =���<=-�<s�<u��<Z��<�A�<���<���<p�<]M�<z��<���<=�<�L�<��<���<��<�;�<�t�<��<j��<M�<�J�<�|�<
��<���<��<4�<I]�<���<p��<+��<c��<�	�<�$�<�<�<�Q�<Cc�<�q�<V|�<���<��<���<1��<�y�<�l�<�Z�<�D�<�)�<�	�<x��<��<׉�<"T�<��<<��<��<lB�<���<&��<F5�<1��<-c�<���<�x�<���<w�<��<�^�<!ʺ<m0�<��<r�<�D�<	��<��<8.�<Us�<W��<��<�*�<�`�<~��<�¢<��<N�<�@�<be�<���<���<!Ǖ<��<���<w�<h0�<G�<x\�<�p�<���<ו�<!��<���<�}<ԭy<�u<d�q<�n<�#j<Af<�^b<�|^<��Z<�V<��R<0�N<
#K<[HG<loC<��?<��;<k�7<�!4<�T0<6�,<��(<�%<.D!<1�<��<�$<�y<l�<5<�<W	<�} <���;c��;=�;o1�;g�;ݮ�;��;Gu�;:��;$��;�3�;-�;-ɪ;ߵ�;'��;֘;G
�;�V�;o��;:�;ءy;� o;f�d;�PZ;
BP;obF;��<;�03;��);_� ;D�;��;5F;���:��:��:�x�:H��:�%�:�ޛ:�֌:�|:V�^:�&B:q�%:v�	:�D�9���9�G_9���8'A,7����XE�����>�ȹb#������Q/�s�G�`S`���x�QY��
T���@��$����F�ú�iϺ�ۺ��溏S�q���ҵ�)u
��0�<���� L!���&��,��J2��7�I�=��5C���H��vN��T�U�Y�_V_�0�d�U�j�%7p��u�vx{�����]���.������Nы� ���.u���G��H����  �  \�=�-=��=Tw=�=h�=�d=�=b� =�O =���<�,�<�r�<��<��<aA�<H��<���<.�<M�<C��<���<�<�L�<��<��<��<�;�<�t�<Z��<���<��<K�<}�<d��<0��<"	�<r4�<�]�<΄�<���<]��<���<
�<�$�<�<�<�Q�<c�<aq�<?|�<Y��<܆�<W��<ށ�<-y�<&l�<�Z�<sD�<t)�<g	�<I��<���<���<T�<��<L��<ݏ�<�B�<���<I��<{5�<|��<{c�<;��<My�<3��<|w�<�<�^�<�ʺ<�0�<Ց�<��<�D�<(��<��<C.�<Ps�<a��<a�<�*�<�`�<:��<�¢</�<��<0@�<e�<���<3��<�ƕ<��<���<3�<U0�<�F�<\\�<�p�<���<땄<2��<з�<z�}<w�y<�u<��q<kn<a$j<�Af<`_b<�}^<��Z<}�V<��R<��N<]#K<HG<�oC<��?<��;<J�7<V!4<�T0<��,<v�(<�%<~C!<��< �<�#<�x<��<Z4<W�<�<
} <"��;���;�;91�;dg�;��;��;�u�;��;M��;�4�;���;�ʪ;0��;���;=ט;��;�W�;o��;;�;L�y;�o;�d;eQZ;�AP;�bF;u�<;�/3;��);� ;��;*�;�C;:��:��:/��:<s�:��:a �:�ۛ:�Ҍ:�|:Z�^:� B:��%:�	:�H�9Z��9�V_92!�8Tl.7�C���;E��ڕ���ȹ��,��-G/�Q�G�LL`�Ҋx�mU��IQ��?�����h��úoiϺ�ۺѻ溒V���������w
�63�	�����O!���&���,�M2���7�i�=�x6C���H�uwN��T���Y��U_���d�%�j�y5p�{�u��v{����D\���-��g���Ћ�u���t���F������  �  m�=�-=��=Xw=�=\�=�d=�=N� =�O =e��<�,�<|r�<׷�<���<$A�< ��<C��<�
�<�L�<��<}��<��<�L�<��<���<��<<�<�t�<���<���<��<QK�<@}�<���<s��<k	�<�4�<�]�<��<��<���<���<5
�<�$�<�<�<Q�< c�<@q�<|�<-��<���<��<���<�x�<�k�<[Z�<8D�<7)�<+	�<��<���<���<�S�<v�<<��<��<�B�<&��<r��<�5�<���<�c�<���<�y�<~��<�w�<K�<>_�<�ʺ<�0�<	��<��<E�<Y��<�<V.�<Ts�<O��<K�<�*�<�`�<��<v¢<��<��<�?�<�d�<b��<�<�ƕ<Y�<���<
�<$0�<�F�<C\�<�p�<���<��<`��<���<�}<ͮy<��u<��q<�n<�$j<]Bf<�_b<E~^<)�Z<��V<��R< O<�#K<�HG<�oC<��?<��;<�7<%!4<1T0<\�,<	�(<n%<�B!<�<��<P#<kx<'�<�3<˚<Q<�| <Z��;��;��;&1�;�g�;���;w	�;av�;��;ዽ;�5�;���;[˪;/��;���;Pؘ;��;�X�;5��;�;�;��y;�o;9�d;�QZ;�AP;bF;��<;�.3;^�);�� ;��;3�;�A;g��:���:���:ko�:��:x�:Vכ:�ό:&|:��^:�B:M�%:I�	:M�9���9�h_9�L�8�J07���;E��˕�<�ȹ�����w��?/�1�G��C`��x�\Q���N��J<��M���췺�ú�jϺ�ۺ���;Y����ǹ��y
�^5������Q!���&�˧,��N2���7���=��7C���H�;xN�T�s�Y�U_�4�d��j��3p�$�u��t{�Ԋ��N[��z,��`����΋�}����r���E��d���홻�  �  v�=�-=��=_w=�=X�=�d=w=?� =�O =1��<u,�<7r�<���<s��<�@�<���<��<�
�<�L�<���<]��<��<~L�<��<���<��<<�<u�<���<
��<�<yK�<�}�<��<���<�	�<�4�<^�<0��<��<���<���<2
�<�$�<�<�<iQ�<
c�<8q�<�{�<��<b��<��<b��<�x�<�k�< Z�<�C�<�(�<	�<���<g��<b��<�S�<��<&��<��<�B�<!��<���<�5�<���<�c�<���<�y�<���<x�<��<�_�<˺<=1�<2��<"�<&E�<q��<�<Y.�<^s�<?��<Y�<�*�<d`�<璤<@¢<��<|�<�?�<}d�<&��<���<Uƕ<(�<F��<��<�/�<�F�<A\�<�p�<Ń�<���<j��<��<,�}<�y<b�u<��q<Bn<�%j<�Bf<�`b<�~^<��Z<t�V<:�R<f O<�#K<�HG<�oC<��?<��;<	�7<2!4<�S0<�,<��(<%<�B!<e�<�<�"<�w<��<t3<X�<�<b| <���;-��;X�;1�;�g�;]��;�	�;�v�;t��;k��;�6�;*��;`̪;G��;X��;�٘;I�;�Y�;ᾇ;b<�;��y;o;�d;�QZ;�AP;QaF;�<;7.3;��);�� ;��;��;�?;���:���:�}�:�j�:͟�:��:�ӛ:�͌:�|:��^:vB:P�%:��	:VK�9߱�9�r_9�k�8617庸��D�iÕ���ȹg���o�6/�}�G��;`�u�x�aO��fM��;������췺��úlϺ�ۺF�溔[�s������"{
�_7���)���R!� '�p�,�~P2�k�7���=�_9C���H�IxN��T��Y�8U_���d�w�j��2p���u��r{�
����Z��7+��y����͋�����!r���D�����M홻�  �  ��=�-=��=bw=�=K�=xd=p=2� =�O =��<T,�<r�<|��<_��<�@�<���<���<�
�<�L�<��<K��<��<kL�<��<���<��<3<�<%u�<Ԭ�<'��<�<�K�<�}�<	��<���<�	�<�4�<-^�<E��<1��<���<���<I
�<�$�<�<�<`Q�<�b�<q�<�{�<���<O��<҅�<A��<�x�<�k�<	Z�<�C�<�(�<��<���<L��<U��<�S�<_�< ��<���<�B�<9��<���<�5�<��<�c�<���<�y�<���<#x�<��<�_�<$˺<Z1�<M��<A�<EE�<���<+�<g.�<`s�<3��<2�<�*�<S`�<В�<+¢<��<^�<�?�<ld�<��<���<5ƕ<�<2��<��<�/�<�F�<$\�<zp�<˃�<��<{��<"��<[�}<W�y<��u<(�q<�n<�%j<	Cf<�`b<�~^<ŝZ<��V<u�R<� O<$K< IG<�oC<��?<��;<��7<� 4<�S0<�,<o�(<� %<NB!<-�<��<�"<�w<b�<,3<!�<�<3| <y��;y��;�;�0�;�g�;���;�	�;
w�;���;׌�;�6�;���;�̪;���;���;�٘;��;NZ�;+��;�<�;]�y;o;��d;-RZ;BP;�`F;¯<;-3;w�);Ӱ ;�;��;u>;��:Z��:0|�:3i�:���:��:Nқ:�ˌ:��{:��^:�B:;�%:�	:�O�9&��9_9��8�527Ӻ��D�F����ȹ����-l��2/���G�18`�c}x��M���K���9������뷺��ú�lϺwۺ����\�����<��2|
�T8��������S!�� '�q�,�_Q2�
�7�s�=��9C���H�)yN��T�׵Y��T_�Y�d���j��1p���u�@r{�����Z���*�����b͋�4����q��yD��S���왻�  �  K�=�*=��=�s= =��=�_=M=�� =�I =��<Y�<2c�<v��<T��<�.�<Dq�<C��<���<N5�<#u�<;��<B��<\/�<bk�<i��<=��<��<*P�<$��<ں�<���<��<�O�<c~�<B��<#��<D��<D&�<FK�<�m�<E��<��<@��<���<��<��<��<�"�<;+�<0�<E1�<�.�<�'�<�<��<_��<8��<c��<���<�|�<�P�<c�<���<��<�i�<�!�<=��<���<�&�<L��<�a�<d��<��<�<4��<��<ㆽ<z��<�f�<�θ<2�< ��<~�<2>�<j��<Kڮ<�!�<�e�<���<��<��<P�<���<��<�ޞ<	�<�0�<pV�<�y�<y��<-��<8ّ<���<��<*�<YB�<dY�<no�<���<���<!��<�}}<�y<=�u<]�q<Sn<�.j<Rf<�tb<��^<�Z<0�V<�S<0O<YK<��G<�C<p�?<<<8B8<x4<�0<��,<U,)<�o%<
�!<�<vS<3�<�<�d<�<�7<�<�$<$L�;�\�;�|�;ͬ�;���;�?�;���;�;���;cA�;�;e��;��;���;͓�;۳�;��;�:�;B��;$!�;�o};	�r;�Yh;^;� T;�J;Sa@;��6;w-;�C$;�;;U];ʨ	;�;�k�:���:���:l��:��:]��:�w�:���:��i:x|L:��/:2�:�)�9N�9�_�9[�9K$08އv�K&���O��;.�����(���A��cZ�1�r�����7���Lĝ���������g����[ͺ�!ٺ����4��{����	��w�i9���կ ��e&��,���1��u7��!=���B�XsH��N���S��gY�}_���d��Yj���o��u��L{�0z���M���!�������ʋ������u��#L��-#�������  �  H�=�*=��=�s==��=�_=C=�� =�I =��<d�<;c�<���<Q��<�.�<Iq�<M��<���<U5�<-u�<&��<D��<d/�<qk�<k��<6��<��<)P�<*��<ɺ�<���<��<�O�<U~�<��<"��<A��<K&�<<K�<�m�<C��<��<A��<���<'��<��<��<�"�<3+�<0�<A1�<�.�<�'�<�<��<c��<H��<h��<���<�|�<�P�<^�<���<��<�i�<	"�<5��<���<�&�<L��<�a�<Y��<��<�<5��<��<φ�<y��<�f�<�θ<�1�<#��<{�<->�<e��<Jڮ<�!�<�e�<���<��<��<$P�<���<��<�ޞ<	�<�0�<zV�< z�<���<8��<8ّ<���<��<*�<\B�<kY�<uo�<v��<���<��<�}}<d�y</�u<f�q<Wn<�.j<�Qf<�tb<��^<��Z<(�V<qS<
0O<YK<��G<��C<y�?<<<AB8<�w4<İ0<��,<Y,)<�o%<!�!<<�S<.�<"<�d< �<�7< �<�$<�K�;�\�;�|�;��;���;�?�;���;�;���;"A�;�;Q��;��;Ɖ�;A��;ٳ�;��;
;�;��;!�;�o};��r;�Yh;�^;T;J;na@;��6;�v-;�C$;�;;�];�	;7;$l�:���:���:���:m�:��:�x�:Y��:��i:}L:t�/:D�:�'�9V�9�^�9��9W 08ʜv��G&�􆹁N���5�U��'�(�R�A��cZ��r�]���R����ĝ������J���<[ͺ�!ٺQ��}���3��~��f�	�w��8����� �7e&�.,�6�1��u7�!=��B��sH��N�~�S��gY��_���d��Yj���o�|�u�-M{�z���M���!��^���ˋ�ퟎ��u��3L��l#��v����  �  =�=�*={�=�s== �=�_=F=�� =�I =?��<z�<Jc�<���<n��<�.�<Tq�<h��<���<i5�<Gu�<0��<V��<b/�<ok�<c��</��<��<P�<��<���<���<��<�O�<C~�<��<��<��<6&�<%K�<�m�<.��<���<>��<���<)��<��<��<�"�<B+�<90�<W1�<�.�<�'�<(�<�<���<`��<s��<���<�|�<�P�<q�<���<(��<�i�<	"�<)��<��<�&�<4��<�a�<>��<���<��<��<��<���<]��<�f�<�θ<�1�<��<`�< >�<]��<>ڮ<�!�<�e�<���<��<��<:P�<���<,��<�ޞ<7	�<1�<�V�<z�<���<Z��<Lّ<���<��<!*�<cB�<kY�<vo�<l��<���<��<�}}<6�y<
�u</�q<n<�.j<�Qf<�tb<[�^<��Z<�V<>S<�/O<�XK<��G<�C<r�?<<<GB8< x4<Ӱ0<�,<~,)<�o%<N�!<-<�S<i�<l<�d<Y�<8<*�<'%<L�;]�;�|�;��;���;�?�;|��;��;���;�@�;��;ƹ�;���;���;֒�;���;&�;�:�;ɡ�;� �;'o};r�r;�Yh;j^;"T;�J;�a@;0�6;Vw-;�D$;\<;�^;n�	;�;In�:���:���:���:��:���:nz�:���:�i:L:��/:z�:1%�9i�97Z�9^�9��/8��v�&R&������S��<�}��R�(��A��eZ�m�r�w���޻��Gŝ�L���O���c���{[ͺz ٺ�����2�����w�	� w��7�%��^� ��d&��,�!�1�u7�2 =���B� sH�eN���S��gY�6_���d�gZj�P p�6�u��M{��z��bN��G"������Lˋ�����=v��vL���#�������  �  6�=�*=x�=�s=	=�=�_=Z=�� =�I =[��<��<|c�<˧�<���<�.�<�q�<���<���<}5�<Xu�<U��<Z��<i/�<tk�<d��<��<��<�O�<���<���<���<t�<�O�<~�<��<���<���<&�<K�<�m�<!��<��<#��<���< ��<��<��<�"�<^+�<?0�<v1�<�.�<%(�<U�<:�<���<���<���<֣�<�|�<�P�<��<���<(��<�i�<"�<)��<e��<�&�<&��<�a�<��<τ�<��<��<��<���<)��<�f�<�θ<�1�<돵<P�<>�<G��<=ڮ<�!�<�e�<���<��<��<KP�<ǂ�<M��<ߞ<U	�<(1�<�V�<Bz�<ě�<w��<hّ<���<��<1*�<hB�<rY�<po�<j��<���<���<�}}<��y<��u<��q<�n<m.j<QQf<atb<�^<r�Z<��V<S<�/O<�XK<e�G<ٯC<m�?<%<<QB8<9x4<"�0<)�,<�,)<.p%<��!<�<&T<��<�<?e<��<Q8<Y�<N%<�L�;/]�;&}�;,��;���;i?�;<��;|�;
��;f@�;Q�;U��;畬;ڈ�;p��;ز�;��;$:�;M��;K �;�n};�r;Yh;�^;� T;NJ;b@;��6;Ex-;E$;b=;�_;�	;R;q�:���:���:���:c�:���:{�:��:ʐi:hL:��/:��:�%�9��9/W�9��9��/8?w��g&�o�� `��/D���c�(���A�]kZ���r���������0Ɲ�����@�������ZͺF ٺ���	��\1�����c�	�yu��6����:� �"c&�,,�9�1�>t7��=���B�{rH�AN�M�S��gY�C_���d��Zj�p��u��N{�{���N��#��8���̋�2����v��M��9$������  �  ,�=�*=w�=�s=
=�=�_=i=�� =�I =���<��<�c�<���<���</�<�q�<���<��<�5�<yu�<q��<g��<~/�<rk�<a��<��<��<�O�<΅�<m��<���<F�<]O�<�}�<���<���<���<�%�<�J�<�m�<���<ث�<��<���<��<��<��<�"�<�+�<i0�<�1�<�.�<](�<��<p�<���<���<���<���<2}�<Q�<��<���<4��<j�<�!�<#��<R��<�&�<���<Ya�<���<���<��<���<F�<M��<���<Sf�<oθ<�1�<���<2�<�=�<8��<4ڮ<�!�<�e�<���<�<��<{P�<���<x��<^ߞ<�	�<k1�<�V�<wz�<���<���<�ّ<���<��<D*�<zB�<|Y�<jo�<j��<���<嫀<8}}<��y<Z�u<}�q<Xn<�-j<�Pf<�sb<��^<�Z<N�V<�S<Y/O<�XK<:�G<ԯC<`�?<)<<uB8<Zx4<^�0<h�,<,-)<�p%<
�!<<�T<K�<<�e<�<�8<ͫ<�%<"M�;t]�;�}�;4��;���;Z?�;���;7�;c��;�?�;��;���;0��;�;���;ޱ�;
�;Z9�;���;��;�m};d�r;�Xh;�^;� T;�J;�b@;��6;ky-;rF$;H?;�`;Ϭ	;�;~t�:Z��:J��:r��:��:1��:�}�:[��:�i:C�L:��/:�:f%�9��9EQ�9_�9�V/8�aw�+�&�L���o��mR�4���(�p�A��qZ���r�u���X����ǝ�:�������^����Yͺ�ٺ��亶��9.������	�zs�5������ �va&��,���1�pr7��=���B��qH��N��S��gY�E_��d�r[j�fp�c�u�zP{��{���O��$��(���͋�㡎��w���M���$�������  �  �=�*=o�=�s=	=�=�_=v=Ӧ =�I =���<�<�c�<G��<��<S/�<�q�<���<L��<�5�<�u�<���<���<�/�<rk�<V��<��<��<�O�<���<:��<a��<��<O�<�}�<j��<k��<{��<�%�<�J�<km�<э�<���<	��<���<��<��<�<#�<�+�<�0�<�1�<:/�<�(�<��<��<(��<���<��<B��<[}�<:Q�<��<���<G��<�i�<�!�<��<H��<|&�<���<7a�<���<_��<4�<m��< �<��<���<�e�<=θ<\1�<���<�<�=�<-��<$ڮ<�!�<�e�<ѥ�<)�<�<�P�<#��<���<�ߞ<�	�<�1�<=W�<�z�<1��<໓<�ّ<��<��<j*�<�B�<wY�<io�<U��<m��<���<�|}<^�y<�u<��q<�
n<�-j<JPf<{sb<�^<z�Z<��V<`S</O<5XK<�G<��C<X�?<#<<�B8<�x4<��0<��,<x-)<q%<��!<x<(U<Ѫ<�<&f<��<"9<�<�%<�M�;^�;�}�;G��;���;D?�;���;��;���;?�;��;���;B��; ��;���;+��;��;�8�;���;'�;�l};`�r;jXh;^;� T;�J;5c@;��6;Qz-;�G$;�@;+c;y�	;�!;�x�:���:U��:���:b �:�:���:[��:�i:�L:��/:d�:� �9�9;I�9B�9?/8��w���&�9%���|���b����(�p�A�KwZ��r�H�������qɝ�����M���Z����Yͺvٺ �����+������	�$r��2����\� ��_&��,���1�4q7�E=���B��pH�<N�+�S��gY��_���d��\j�}p���u��Q{��|���P���$��>����͋�����x���N��%��O����  �  �=�*=a�=�s==�=�_=�=� =
J =���<W�<3d�<���<L��<�/�<9r�<C��<���<6�<�u�<���<���<�/�<�k�<I��<���<h�<�O�<���<��<,��<��<�N�<T}�<��<+��<:��<p%�<fJ�<2m�<���<���<���<i��<,��<��<�<##�<�+�<�0�<�1�<�/�<�(�<�<��<`��<G��<K��<���<�}�<lQ�<��<���<W��<�i�<	"�<���<%��<V&�<���< a�<m��<'��<��<)��<��<���<l��<�e�<θ<1�<e��<��<�=�<	��<ڮ<"�<�e�<ᥩ<<�<8�<�P�<W��<���<�ߞ<
�<�1�<�W�<�z�<s��<!��<�ّ<S��<�<~*�<�B�<�Y�<qo�<=��<S��<���<�|}<ؠy<��u<��q<A
n<-j<�Of<�rb<��^<�Z<x�V<�S<�.O<�WK<ւG<y�C<Y�?<L<<�B8<�x4<̱0<5�,<�-)<q%<�!<<�U<9�<W<�f<*�<�9<��<e&<N�;r^�;�}�;���;���;�>�;@��;	�;g��;>�;$�;���;[��;��;P��;<��;��;�7�;���;Q�;�k};d�r;�Wh;`^;�T;4J;�c@;c�6;�{-;�I$;�A;ee;��	;|$;�|�:?��:x��:���:�$�:|��:���:팃:��i:l�L:��/:�:v�9�޷9�@�9҅9,�.8�Lx���&�	5��C����w�x���(���A��}Z�; s������Ñ�[˝��é�F���ȇ��LYͺ0ٺ���6���(�������	�p�d0�4��=� �R]&��,���1�p7��=���B�&pH��N���S��gY��_�{�d��]j��p���u��S{��}���Q���%�������΋� ���oy��O���&�������  �  ��=�*=_�=�s=="�=�_=�=� =-J =8��<��<rd�<֨�<���<�/�<yr�<s��<���<G6�<�u�<ɴ�<���<�/�<�k�<;��<���<U�<sO�<Q��<ι�<���<~�<�N�<}�<ߩ�<���<���<(%�<2J�< m�<���<|��<���<c��<��<��<1�<C#�<�+�<�0�<E2�<�/�<	)�<O�<=�<���<���<���<���<�}�<�Q�< �<��<r��<j�<�!�<���<��<<&�<w��<�`�<=��<ۃ�<��<ҏ�<i�<r��<��<xe�<�͸<�0�<*��<��<�=�<���< ڮ<�!�<�e�<���<[�<W�<Q�<���<-��<��<[
�<32�<�W�<9{�<���<X��<6ڑ<|��<:�<�*�<�B�<�Y�<Yo�<;��<B��<~��<F|}<��y<�u<�q<�	n<c,j<8Of<Xrb<�^<��Z<��V<}S<X.O<�WK<��G<m�C<+�?<O<<�B8<�x4<�0<��,<Z.)<�q%<~�!<�<QV<�<�<>g<��<(:<�<�&<�N�;�^�;H~�;���;o��;�>�;��;��;���;�=�;)�;µ�;7��;��;���;��;��;�6�;>��;��;:j};��r;Wh;J^;� T;�J;�d@;q�6;�|-;)K$;D;g;i�	;h&;���:}�:`��:y��:$(�:��:��:k��:Ӟi:A�L:L�/:<�:��9�ٷ9S;�9�p9�M.8�x���&�4E������k��y��)���A���Z��s�H����ő��̝�qĩ����������Wͺvٺ�����%�����&�	�n�h.�u��� �Y[&��,�3�1��m7�Z=���B�RoH�N�Y�S�zhY��_��d��^j�2p��u��U{��~���R��'��Z���Ћ�#����z��mP��:'�������  �  �=�*=Y�=�s==+�=`=�=� =CJ =g��<��<�d�<��<���<0�<�r�<���<���<k6�<v�<��<���<�/�<�k�<@��<���<0�<ZO�<��<���<���<F�<WN�<�|�<���<���<���<�$�<J�<�l�<Z��<a��<���<d��<��<��<5�<a#�<,�<1�<w2�<�/�<Y)�<��<y�<���<���<���<��<�}�<�Q�<7 �<$��<u��<j�<�!�<���<��<&�<P��<�`�<��<���<v�<���< �<)��<���<>e�<o͸<�0�<���<��<o=�<���<ڮ<�!�<�e�<��<}�<{�<$Q�<���<e��<R��<�
�<u2�<�W�<{{�<���<���<fڑ<���<e�<�*�<�B�<�Y�<Yo�<3��<��<c��<�{}<8�y<��u<��q<V	n<�+j<�Nf<�qb<��^<	�Z<��V<2S<�-O<tWK<a�G<S�C<-�?<Y<<�B8<2y4<v�0<��,<�.)<Tr%<�!<$<�V<|�<E<�g<�<�:<^�<'<eO�;G_�;�~�;���;���;�>�;���;F�;��;=�;5�;���;]��;��;���;��;\�;�5�;���;�;i};�r;1Vh;k^;� T;LJ;e@;u�6;A~-;L$;�E;�h;��	;?(;���:��:���:���:E+�:��:爒:���:Ţi:�L:��/:$�:�9yӷ9)4�9&_9^�-8��x���&��P��ΰ��L��	��)�j�A��Z��	s�V���pǑ��Ν��ũ�����܈��RVͺ�ٺ;�亯~��"�����X�	��k��,�`��8� �JY&��,�ɽ1�Sl7�^=�7�B�ynH��N��S�zhY�_�8�d��_j��p�&�u�6W{�����S��,(��X���2ы�쥎�z{��MQ���'��w����  �  م=�*=O�=�s==,�=`=�=(� =WJ =���< �<�d�<H��<#��<W0�<�r�<��<$��<�6�<Hv�<��<���<�/�<�k�<4��<���<�<:O�<���<l��<��<�<#N�<�|�<Z��<`��<���<�$�<�I�<�l�<4��<D��<���<Q��<��<��<B�<w#�<.,�<C1�<�2�<0�<�)�<��<��<(��<���<���<��<~�<�Q�<V �<:��<���<j�<�!�<���<��<�%�<(��<f`�<���<b��<7�<R��<��<���<���<e�<C͸<w0�<Ȏ�<e�<S=�<̍�<�ٮ<�!�<�e�<��<��<��<PQ�<<���<}��<�
�<�2�<<X�<�{�<$��<���<�ڑ<���<z�<�*�<�B�<�Y�<[o�<��<��<G��<�{}<ȟy<J�u<,�q<�n<j+j</Nf<[qb<&�^<��Z<.�V<�S<�-O<7WK<@�G<*�C<*�?<b<<�B8<Zy4<��0<"�,</)<�r%<z�!<�<=W<��<�<;h<��<�:<��<a'<�O�;�_�;�~�;��;t��;i>�;H��;��;n��;*<�;��;/��;���;A��;���;;��;l�;5�;ќ�;T�;�g};?�r;�Uh;�^;&T;�J;�e@;;�6;2-;�M$;G;'j;Q�	;*;z��:0	�:���:9��:c.�:���:勒:%��:եi:��L:��/:�:(�9з9]-�9.M9K�-8>my��'�m_��I�������+)�V�A��Z�s�ײ���ɑ�!Н��Ʃ�����q���bVͺ�ٺ���|� �������	�Bj��*����J� ��W&�!,��1�k7��=���B��mH�}N���S�nhY��_���d�h`j��p��u��X{������T���(��e���ҋ�٦��;|��R���(�������  �  ƅ=�*=M�=�s==0�=`=�=7� =dJ =���<$ �<e�<x��<=��<�0�<s�<��<F��<�6�<\v�<��<���<�/�<�k�<-��<���<�<O�<��<O��<b��<��<�M�<p|�<4��<A��<Z��<�$�<�I�<�l�<"��<&��<���<F��<��<��<V�<�#�<:,�<c1�<�2�<>0�<�)�<��<��<J��<$��<��<D��<9~�< R�<` �<E��<���<j�<�!�<���<��<�%�<��<W`�<���<A��<��<+��<��<�<i��<�d�<"͸<T0�<���<B�<>=�<ō�<�ٮ<�!�<�e�<'��<��<��<jQ�<��<���<���<�
�<�2�<jX�<�{�<C��<㼓<�ڑ<���<��<�*�<�B�<�Y�<Vo�<��<	��<"��<�{}<��y<�u<��q<on<*+j<�Mf<qb<��^<Q�Z<��V<�S<�-O<�VK<*�G<�C<�?<d<<C8<�y4<��0<^�,<:/)<s%<��!<�<�W<0�<0<�h<��<;;<��<�'<
P�;`�;�~�;��;e��;e>�;��;K�;X��;�;�;:�;��;㏬;���;��;Ȭ�;��;�4�;V��;�;|g};]�r;�Uh;�^;T;�J;2f@;��6;�-;�N$;�G;�k;_�	;�+;��:g�:���:M��:?1�:���:֍�:ؔ�:a�i:ďL:��/:*�:s�9gϷ9l'�9�B9��-8��y�h'��l��Ǻ������)�c�A���Z��s�J����ˑ�>ѝ��Ʃ�*���Ї���Vͺٺ���2{�X�����t�	�:i�\)����ӟ �aV&�#
,�غ1�?j7��=��B�0mH�N���S��hY��_�ոd��aj�	p���u��Y{� ���tU��u)������ҋ������|��vR��)��* ���  �  =�*=L�=�s==6�=`=�=>� =qJ =���<F �<6e�<���<Y��<�0�<As�<%��<Y��<�6�<mv�<'��<���<�/�<�k�</��<���<��<O�<ׄ�<;��<?��<��<�M�<K|�<��< ��<N��<x$�<�I�<�l�<��<��<���<J��<��<��<[�<�#�<S,�<w1�<�2�<Q0�<�)�<�<��<a��<8��<F��<W��<Q~�<R�<w �<T��<���<$j�<�!�<���<��<�%�<���<:`�<���<��<��<��<��<���<S��<�d�<�̸<=0�<���<3�<*=�<���<�ٮ<�!�<�e�<)��<��<��<Q�<"��<Գ�<���<�<�2�<|X�<�{�<h��<�<�ڑ<���<��<�*�<�B�<�Y�<Yo�<��<���<��<U{}<t�y<��u<��q<Wn<�*j<�Mf<�pb<��^<#�Z<��V<`S<c-O<�VK<�G<�C<�?<l<<C8<�y4<�0<y�,<n/)<0s%<�!<'<�W<k�<X<�h<�<d;<'�<�'<dP�;+`�;�~�;��;u��;G>�;Ҡ�;3�;��;y;�;��;B��;���;$��;���;L��;x�;/4�;���;��;�f};�r;VUh;�^;&T;�J;`f@;!�6;l�-;PO$;�H;3l;��	;R,;$��:��:��:���:}2�:¡:G��:[��:��i:K�L: �/:�:��9#˷9�#�9�79�O-8K�y�6/'��o���ͺ����O��)��A��Z��s����`̑�[ҝ��ǩ����������Uͺ�ٺ����y����I����	��g��(����E� �\U&�	,�b�1�ki7��=�?�B�mH��N�ÿS��hY��_�c�d��aj��	p�3�u��Z{������U��*�����Ӌ�ڧ��<}���R��f)��� ���  �  ̅=�*=I�=�s==;�=`=�=<� =yJ =���<E �<5e�<���<���<�0�<As�<��<b��<�6�<mv�<,��<���<�/�<�k�<)��<���< �<O�<Ą�<<��<4��<��<�M�<D|�<��<��<J��<m$�<�I�<vl�<��<,��<���<C��<��<��<^�<�#�<T,�<s1�<�2�<M0�<�)�<�<�<{��<6��<K��<P��<\~�<R�<v �<X��<���<)j�<�!�<���<��<�%�<���<0`�<���<��<��<���<��<���<G��<�d�<�̸<?0�<���<<�<1=�<���<�ٮ<�!�<�e�<&��<��<��<�Q�<,��<γ�<���<�<
3�<�X�<�{�<l��<�<�ڑ<���<��<�*�<�B�<�Y�<Jo�<��<���<-��<>{}<h�y<��u<��q<Kn<�*j<�Mf<�pb<��^<�Z<��V<ZS<G-O<WK<�G<�C<�?<f<<3C8<�y4<��0<r�,<�/)<6s%<�!<%<�W<��<a<�h<�<v;<A�<�'<wP�;'`�;2�;��;^��;?>�;��;i�;���;~;�;��;��;{��;
��;���;��;j�;4�;���;��;�f};��r;KUh;�^;� T;�J;�f@;N�6;s�-;7O$;+I;l;ɸ	;S,;���:��:���:-��:2�:�¡:I��:Q��:�i:h�L:��/:̓:a�9Lʷ9�'�9�89t=-8A�y��4'��p��_Һ������)�?�A�W�Z�]s������ˑ��ѝ��ǩ�7���Ĉ��Uͺ�ٺ����y�j������	��g��(����� �dU&��,�[�1��h7��=�/�B�mH��N�ܿS��hY�_�d�d�8aj�P
p�c�u��Z{������U��Q*��s���VӋ�����h}��S��s)��� ���  �  =�*=L�=�s==6�=`=�=>� =qJ =���<F �<6e�<���<Y��<�0�<As�<%��<Y��<�6�<mv�<'��<���<�/�<�k�</��<���<��<O�<ׄ�<;��<?��<��<�M�<K|�<��< ��<N��<x$�<�I�<�l�<��<��<���<J��<��<��<[�<�#�<S,�<w1�<�2�<Q0�<�)�<�<��<a��<8��<F��<W��<Q~�<R�<w �<T��<���<$j�<�!�<���<��<�%�<���<:`�<���<��<��<��<��<���<S��<�d�<�̸<=0�<���<3�<*=�<���<�ٮ<�!�<�e�<)��<��<��<Q�<"��<Գ�<���<�<�2�<|X�<�{�<h��<�<�ڑ<���<��<�*�<�B�<�Y�<Yo�<��<���<��<U{}<t�y<��u<��q<Wn<�*j<�Mf<�pb<��^<#�Z<��V<`S<c-O<�VK<�G<�C<�?<l<<C8<�y4<�0<y�,<n/)<0s%<�!<'<�W<k�<X<�h<�<d;<'�<�'<dP�;+`�;�~�;��;u��;G>�;Ҡ�;3�;��;y;�;��;B��;���;$��;���;L��;x�;/4�;���;��;�f};�r;VUh;�^;&T;�J;`f@;!�6;l�-;PO$;�H;3l;��	;R,;$��:��:��:���:}2�:¡:G��:[��:��i:K�L: �/:�:��9#˷9�#�9�79�O-8K�y�6/'��o���ͺ����O��)��A��Z��s����`̑�[ҝ��ǩ����������Uͺ�ٺ����y����I����	��g��(����E� �\U&�	,�b�1�ki7��=�?�B�mH��N�ÿS��hY��_�c�d��aj��	p�3�u��Z{������U��*�����Ӌ�ڧ��<}���R��f)��� ���  �  ƅ=�*=M�=�s==0�=`=�=7� =dJ =���<$ �<e�<x��<=��<�0�<s�<��<F��<�6�<\v�<��<���<�/�<�k�<-��<���<�<O�<��<O��<b��<��<�M�<p|�<4��<A��<Z��<�$�<�I�<�l�<"��<&��<���<F��<��<��<V�<�#�<:,�<c1�<�2�<>0�<�)�<��<��<J��<$��<��<D��<9~�< R�<` �<E��<���<j�<�!�<���<��<�%�<��<W`�<���<A��<��<+��<��<�<i��<�d�<"͸<T0�<���<B�<>=�<ō�<�ٮ<�!�<�e�<'��<��<��<jQ�<��<���<���<�
�<�2�<jX�<�{�<C��<㼓<�ڑ<���<��<�*�<�B�<�Y�<Vo�<��<	��<"��<�{}<��y<�u<��q<on<*+j<�Mf<qb<��^<R�Z<��V<�S<�-O<�VK<*�G<�C<�?<d<<C8<�y4<��0<^�,<:/)<s%<��!<�<�W<0�<0<�h<��<;;<��<�'<
P�;`�;�~�;��;e��;e>�;��;K�;X��;�;�;:�;��;⏬;���;��;Ȭ�;��;�4�;V��;�;|g};]�r;�Uh;�^;T;�J;2f@;��6;�-;�N$;�G;�k;_�	;�+;��:g�:���:M��:?1�:���:֍�:ؔ�:a�i:ďL:��/:*�:s�9gϷ9l'�9�B9��-8��y�h'��l��Ǻ������)�c�A���Z��s�J����ˑ�>ѝ��Ʃ�*���Ї���Vͺٺ���2{�X�����t�	�:i�\)����ӟ �aV&�#
,�غ1�?j7��=��B�0mH�N���S��hY��_�ոd��aj�	p���u��Y{� ���tU��u)������ҋ������|��vR��)��* ���  �  م=�*=O�=�s==,�=`=�=(� =WJ =���< �<�d�<H��<#��<W0�<�r�<��<$��<�6�<Hv�<��<���<�/�<�k�<4��<���<�<:O�<���<l��<��<�<#N�<�|�<Z��<`��<���<�$�<�I�<�l�<4��<D��<���<Q��<��<��<B�<w#�<.,�<C1�<�2�<0�<�)�<��<��<(��<���<���<��<~�<�Q�<V �<:��<���<j�<�!�<���<��<�%�<(��<f`�<���<b��<7�<R��<��<���<���<e�<C͸<w0�<Ȏ�<e�<S=�<̍�<�ٮ<�!�<�e�<��<��<��<PQ�<<���<}��<�
�<�2�<<X�<�{�<$��<���<�ڑ<���<z�<�*�<�B�<�Y�<[o�<��<��<G��<�{}<ȟy<J�u<,�q<�n<j+j</Nf<[qb<&�^<��Z<.�V<�S<�-O<7WK<@�G<*�C<*�?<b<<�B8<Zy4<��0<"�,</)<�r%<z�!<�<=W<��<�<;h<��<�:<��<a'<�O�;�_�;�~�;��;t��;i>�;H��;��;m��;*<�;��;/��;���;A��;���;;��;l�;5�;ќ�;T�;�g};?�r;�Uh;�^;&T;�J;�e@;;�6;2-;�M$;G;'j;Q�	;*;z��:0	�:���:9��:c.�:���:勒:%��:եi:��L:��/:�:(�9з9]-�9.M9K�-8>my��'�m_��I�������+)�V�A��Z�s�ײ���ɑ�!Н��Ʃ�����q���bVͺ�ٺ���|� �������	�Bj��*����J� ��W&�!,��1�k7��=���B��mH�}N���S�nhY��_���d�h`j��p��u��X{������T���(��e���ҋ�٦��;|��R���(�������  �  �=�*=Y�=�s==+�=`=�=� =CJ =g��<��<�d�<��<���<0�<�r�<���<���<k6�<v�<��<���<�/�<�k�<@��<���<0�<ZO�<��<���<���<F�<WN�<�|�<���<���<���<�$�<J�<�l�<Z��<a��<���<d��<��<��<5�<a#�<,�<1�<w2�<�/�<Y)�<��<y�<���<���<���<��<�}�<�Q�<7 �<$��<u��<j�<�!�<���<��<&�<P��<�`�<��<���<v�<���< �<)��<���<>e�<o͸<�0�<���<��<o=�<���<ڮ<�!�<�e�<��<}�<{�<$Q�<���<e��<R��<�
�<u2�<�W�<{{�<���<���<fڑ<���<e�<�*�<�B�<�Y�<Yo�<3��<��<c��<�{}<8�y<��u<��q<V	n<�+j<�Nf<�qb<��^<	�Z<��V<2S<�-O<tWK<a�G<S�C<-�?<Y<<�B8<2y4<v�0<��,<�.)<Tr%<�!<$<�V<|�<E<�g<�<�:<^�<'<eO�;G_�;�~�;���;���;�>�;���;F�;��;=�;5�;���;]��;��;���;��;\�;�5�;���;�;i};�r;1Vh;k^;� T;LJ;e@;u�6;A~-;L$;�E;�h;��	;?(;���:��:���:���:E+�:��:爒:���:Ţi:�L:��/:$�:�9yӷ9)4�9&_9^�-8��x���&��P��ΰ��L��	��)�j�A��Z��	s�V���pǑ��Ν��ũ�����܈��RVͺ�ٺ;�亯~��"�����X�	��k��,�`��8� �JY&��,�ɽ1�Sl7�^=�7�B�ynH��N��S�zhY�_�8�d��_j��p�&�u�6W{�����S��,(��X���2ы�쥎�z{��MQ���'��w����  �  ��=�*=_�=�s=="�=�_=�=� =-J =8��<��<rd�<֨�<���<�/�<yr�<s��<���<G6�<�u�<ɴ�<���<�/�<�k�<;��<���<U�<sO�<Q��<ι�<���<~�<�N�<}�<ߩ�<���<���<(%�<2J�< m�<���<|��<���<c��<��<��<1�<C#�<�+�<�0�<E2�<�/�<	)�<O�<=�<���<���<���<���<�}�<�Q�< �<��<r��<j�<�!�<���<��<<&�<w��<�`�<=��<ۃ�<��<ҏ�<i�<r��<��<xe�<�͸<�0�<*��<��<�=�<���< ڮ<�!�<�e�<���<[�<W�<Q�<���<-��<��<[
�<32�<�W�<9{�<���<X��<6ڑ<|��<:�<�*�<�B�<�Y�<Yo�<:��<B��<~��<F|}<��y<�u<�q<�	n<c,j<8Of<Xrb<�^<��Z<��V<}S<X.O<�WK<��G<m�C<+�?<O<<�B8<�x4<�0<��,<Z.)<�q%<~�!<�<QV<�<�<>g<��<(:<�<�&<�N�;�^�;H~�;���;o��;�>�;��;��;���;�=�;)�;���;6��;��;���;��;��;�6�;>��;��;:j};��r;Wh;J^;� T;�J;�d@;q�6;�|-;)K$;D;g;i�	;h&;���:}�:`��:y��:$(�:��:��:k��:Ӟi:A�L:L�/:<�:��9�ٷ9S;�9�p9�M.8�x���&�4E������k��y��)���A���Z��s�H����ő��̝�qĩ����������Wͺvٺ�����%�����&�	�n�h.�u��� �Y[&��,�3�1��m7�Z=���B�RoH�N�Y�S�zhY��_��d��^j�2p��u��U{��~���R��'��Z���Ћ�#����z��mP��:'�������  �  �=�*=a�=�s==�=�_=�=� =
J =���<W�<3d�<���<L��<�/�<9r�<C��<���<6�<�u�<���<���<�/�<�k�<I��<���<h�<�O�<���<��<,��<��<�N�<T}�<��<+��<:��<p%�<fJ�<2m�<���<���<���<i��<,��<��<�<##�<�+�<�0�<�1�<�/�<�(�<�<��<`��<G��<K��<���<�}�<lQ�<��<���<W��<�i�<	"�<���<%��<V&�<���< a�<m��<'��<��<)��<��<���<l��<�e�<θ<1�<e��<��<�=�<	��<ڮ<"�<�e�<ᥩ<<�<8�<�P�<W��<���<�ߞ<
�<�1�<�W�<�z�<s��<!��<�ّ<S��<�<~*�<�B�<�Y�<qo�<=��<S��<���<�|}<ؠy<��u<��q<A
n<-j<�Of<�rb<��^<�Z<x�V<�S<�.O<�WK<ւG<y�C<Y�?<L<<�B8<�x4<̱0<5�,<�-)<q%<�!<<�U<9�<W<�f<*�<�9<��<e&<N�;r^�;�}�;���;���;�>�;@��;	�;g��;>�;$�;���;[��;��;P��;<��;��;�7�;���;Q�;�k};d�r;�Wh;`^;�T;4J;�c@;c�6;�{-;�I$;�A;ee;��	;|$;�|�:?��:x��:���:�$�:|��:���:팃:��i:l�L:��/:�:v�9�޷9�@�9҅9,�.8�Lx���&�	5��C����w�x���(���A��}Z�; s������Ñ�[˝��é�F���ȇ��LYͺ0ٺ���6���(�������	�p�d0�4��=� �R]&��,���1�p7��=���B�&pH��N���S��gY��_�{�d��]j��p���u��S{��}���Q���%�������΋� ���oy��O���&�������  �  �=�*=o�=�s=	=�=�_=v=Ӧ =�I =���<�<�c�<G��<��<S/�<�q�<���<L��<�5�<�u�<���<���<�/�<rk�<V��<��<��<�O�<���<:��<a��<��<O�<�}�<j��<k��<{��<�%�<�J�<km�<э�<���<	��<���<��<��<�<#�<�+�<�0�<�1�<:/�<�(�<��<��<(��<���<��<B��<[}�<:Q�<��<���<G��<�i�<�!�<��<H��<|&�<���<7a�<���<_��<4�<m��< �<��<���<�e�<=θ<\1�<���<�<�=�<-��<$ڮ<�!�<�e�<ѥ�<)�<�<�P�<#��<���<�ߞ<�	�<�1�<=W�<�z�<1��<໓<�ّ<��<��<j*�<�B�<wY�<io�<U��<m��<���<�|}<^�y<�u<��q<�
n<�-j<JPf<{sb<�^<z�Z<��V<`S</O<5XK<�G<��C<X�?<#<<�B8<�x4<��0<��,<x-)<q%<��!<x<(U<Ѫ<�<&f<��<"9<�<�%<�M�;^�;�}�;G��;���;D?�;���;��;���;?�;��;���;B��; ��;���;+��;��;�8�;���;'�;�l};`�r;jXh;^;� T;�J;5c@;��6;Qz-;�G$;�@;+c;y�	;�!;�x�:���:U��:���:b �:�:���:[��:�i:�L:��/:d�:� �9�9;I�9B�9?/8��w���&�9%���|���b����(�p�A�KwZ��r�H�������qɝ�����M���Z����Yͺvٺ �����+������	�$r��2����\� ��_&��,���1�4q7�E=���B��pH�<N�+�S��gY��_���d��\j�}p���u��Q{��|���P���$��>����͋�����x���N��%��O����  �  ,�=�*=w�=�s=
=�=�_=i=�� =�I =���<��<�c�<���<���</�<�q�<���<��<�5�<yu�<q��<g��<~/�<rk�<a��<��<��<�O�<΅�<m��<���<F�<]O�<�}�<���<���<���<�%�<�J�<�m�<���<ث�<��<���<��<��<��<�"�<�+�<i0�<�1�<�.�<](�<��<p�<���<���<���<���<2}�<Q�<��<���<4��<j�<�!�<#��<R��<�&�<���<Ya�<���<���<��<���<F�<M��<���<Sf�<oθ<�1�<���<2�<�=�<8��<4ڮ<�!�<�e�<���<�<��<{P�<���<x��<^ߞ<�	�<k1�<�V�<wz�<���<���<�ّ<���<��<D*�<zB�<|Y�<jo�<j��<���<嫀<8}}<��y<Z�u<}�q<Xn<�-j<�Pf<�sb<��^<�Z<N�V<�S<Y/O<�XK<:�G<ԯC<`�?<)<<uB8<Zx4<^�0<h�,<,-)<�p%<
�!<<�T<K�<<�e<�<�8<ͫ<�%<"M�;t]�;�}�;4��;���;Z?�;���;7�;c��;�?�;��;���;/��;�;���;ޱ�;
�;Z9�;���;��;�m};d�r;�Xh;�^;� T;�J;�b@;��6;ky-;rF$;H?;�`;Ϭ	;�;~t�:Z��:J��:r��:��:1��:�}�:[��:�i:C�L:��/:�:f%�9��9EQ�9_�9�V/8�aw�+�&�L���o��mR�4���(�p�A��qZ���r�u���X����ǝ�:�������^����Yͺ�ٺ��亶��9.������	�zs�5������ �va&��,���1�pr7��=���B��qH��N��S��gY�E_��d�r[j�fp�c�u�zP{��{���O��$��(���͋�㡎��w���M���$�������  �  6�=�*=x�=�s=	=�=�_=Z=�� =�I =[��<��<|c�<˧�<���<�.�<�q�<���<���<}5�<Xu�<U��<Z��<i/�<tk�<d��<��<��<�O�<���<���<���<t�<�O�<~�<��<���<���<&�<K�<�m�<!��<��<#��<���< ��<��<��<�"�<^+�<?0�<v1�<�.�<%(�<U�<:�<���<���<���<֣�<�|�<�P�<��<���<(��<�i�<"�<)��<e��<�&�<&��<�a�<��<τ�<��<��<��<���<)��<�f�<�θ<�1�<돵<P�<>�<G��<=ڮ<�!�<�e�<���<��<��<KP�<ǂ�<M��<ߞ<U	�<(1�<�V�<Bz�<ě�<w��<hّ<���<��<1*�<hB�<rY�<po�<j��<���<���<�}}<��y<��u<��q<�n<m.j<QQf<atb<�^<r�Z<��V<S<�/O<�XK<e�G<ٯC<m�?<%<<QB8<9x4<"�0<)�,<�,)<.p%<��!<�<&T<��<�<?e<��<Q8<Y�<N%<�L�;/]�;%}�;,��;���;i?�;;��;|�;
��;f@�;P�;U��;畬;ڈ�;p��;ز�;��;$:�;M��;K �;�n};�r;Yh;�^;� T;NJ;b@;��6;Ex-;E$;b=;�_;�	;R;q�:���:���:���:c�:���:{�:��:ʐi:hL:��/:��:�%�9��9/W�9��9��/8?w��g&�o�� `��/D���c�(���A�]kZ���r���������0Ɲ�����@�������ZͺF ٺ���	��\1�����c�	�yu��6����:� �"c&�,,�9�1�>t7��=���B�{rH�AN�M�S��gY�C_���d��Zj�p��u��N{�{���N��#��8���̋�2����v��M��9$������  �  =�=�*={�=�s== �=�_=F=�� =�I =?��<z�<Jc�<���<n��<�.�<Tq�<h��<���<i5�<Gu�<0��<V��<b/�<ok�<c��</��<��<P�<��<���<���<��<�O�<C~�<��<��<��<6&�<%K�<�m�<.��<���<>��<���<)��<��<��<�"�<B+�<90�<W1�<�.�<�'�<(�<�<���<`��<s��<���<�|�<�P�<q�<���<(��<�i�<	"�<)��<��<�&�<4��<�a�<>��<���<��<��<��<���<]��<�f�<�θ<�1�<��<`�< >�<]��<>ڮ<�!�<�e�<���<��<��<:P�<���<,��<�ޞ<7	�<1�<�V�<z�<���<Z��<Lّ<���<��<!*�<cB�<kY�<vo�<l��<���<��<�}}<6�y<
�u</�q<n<�.j<�Qf<�tb<[�^<��Z<�V<>S<�/O<�XK<��G<�C<r�?<<<HB8< x4<Ӱ0<�,<~,)<�o%<N�!<-<�S<i�<l<�d<Y�<8<*�<'%<L�;]�;�|�;��;���;�?�;{��;��;���;�@�;��;ƹ�;���;���;֒�;���;&�;�:�;ɡ�;� �;'o};r�r;�Yh;j^;"T;�J;�a@;0�6;Vw-;�D$;\<;�^;n�	;�;In�:���:���:���:��:���:nz�:���:�i:L:��/:z�:1%�9i�97Z�9^�9��/8��v�&R&������S��<�}��R�(��A��eZ�m�r�w���޻��Gŝ�L���O���c���{[ͺz ٺ�����2�����w�	� w��7�%��^� ��d&��,�!�1�u7�2 =���B� sH�eN���S��gY�6_���d�gZj�P p�6�u��M{��z��bN��G"������Lˋ�����=v��vL���#�������  �  H�=�*=��=�s==��=�_=C=�� =�I =��<d�<;c�<���<Q��<�.�<Iq�<M��<���<U5�<-u�<&��<D��<d/�<qk�<k��<6��<��<)P�<*��<ɺ�<���<��<�O�<U~�<��<"��<A��<K&�<<K�<�m�<C��<��<A��<���<'��<��<��<�"�<3+�<0�<A1�<�.�<�'�<�<��<c��<H��<h��<���<�|�<�P�<^�<���<��<�i�<	"�<5��<���<�&�<L��<�a�<Y��<��<�<5��<��<φ�<y��<�f�<�θ<�1�<#��<{�<->�<e��<Jڮ<�!�<�e�<���<��<��<$P�<���<��<�ޞ<	�<�0�<zV�< z�<���<8��<8ّ<���<��<*�<\B�<kY�<uo�<v��<���<��<�}}<d�y</�u<f�q<Wn<�.j<�Qf<�tb<��^<��Z<(�V<qS<
0O<YK<��G<��C<y�?<<<AB8<�w4<İ0<��,<Y,)<�o%<!�!<<�S<.�<"<�d< �<�7< �<�$<�K�;�\�;�|�;��;���;�?�;���;�;���;"A�;�;Q��;��;Ɖ�;A��;ٳ�;��;
;�;��;!�;�o};��r;�Yh;�^;T;J;na@;��6;�v-;�C$;�;;�];�	;7;$l�:���:���:���:m�:��:�x�:Y��:��i:}L:t�/:D�:�'�9V�9�^�9��9W 08ʜv��G&�􆹁N���5�U��'�(�R�A��cZ��r�]���R����ĝ������J���<[ͺ�!ٺQ��}���3��~��f�	�w��8����� �7e&�.,�6�1��u7�!=��B��sH��N�~�S��gY��_���d��Yj���o�|�u�-M{�z���M���!��^���ˋ�ퟎ��u��3L��l#��v����  �  %�=g(=��=vp=0=��=[=7� =� =�C =V��<��<�T�<͗�<���<��<?^�<��<:��<��<]�<���<R��<�<�M�<,��<u��<���<P,�<�`�<���<��<��<#�<$P�<{�<��<I��<:��<?�<�3�<R�<�m�<���<���<1��<t��<���<W��<���<z��<���<���<#��<<��<V��<��<Ȅ�<Ef�<�B�<��<���<O��<P��<�D�<��<Z��<8k�<+�<���<!^�<���<$��<r�<d��<�+�<|��<�#�<"��<'�<q�<7ֶ<H6�<�<��<�;�<�<(Ԭ<��<]�<0��<�ץ<)�<zE�<�w�<���<�Ԝ<d��<�'�<�M�<Nr�<���<���<�ԏ<D�<k�<^)�<"C�<�[�<�s�<p��<���<l}<�y<5�u<��q<�n<�7j<&`f<c�b<q�^<��Z<�W<*1S<�]O<R�K<+�G<�C<�!@<�W<<��8<��4<t
1<�K-<_�)<G�%<l'"<�x<&�<�*<Ҋ<�<�\<
�<�G<��<��;���;���;��;_c�;���;�+�;ժ�;J<�;4��;��;+i�;3L�;�D�;S�;�w�;N��;�;�n�;l�;��;;iv;��k;a�a; �W;��M;��C;S:;��0;�';��;W�;�;�O;;��:��:˹�:���:Ӷ:B�:3�:�ψ:��s:�xV:�9:^�:{� :��9Qi�9{�79o��8���r��EOq�����w�߹�s	��"�/�;��T�erm�?���9���^���s���w���o���X˺�5׺<������n�x��������fL�� ���%�F�+�C1���6�g�<��^B��H�&�M�imS��Y���^��td�O!j���o�X{u�F({�2k���A��L��g����ȋ�Ơ���y��S���-���	���  �  �=b(=�=tp=9=Ƿ=[=8� =� =�C =[��<��<�T�<Η�<���<��<F^�<��<6��<��<]�<���<g��<�<�M�<!��<g��<r��<?,�<�`�<���<#��<#��<|#�<*P�<{�< ��<D��<F��<.�<�3�<�Q�<�m�<���<֜�<3��<���<���<d��<���<x��<���<���<+��<V��<<��<͞�<���<Jf�<�B�<q�<���<V��<Y��<�D�<��<^��<k�<,�<}��<^�<���<��<|�<^��<�+�<���<�#�<��<'�<q�< ֶ<T6�<味<��<};�<���<6Ԭ<��</]�<3��<�ץ< �<qE�<�w�<���<�Ԝ<<��<�'�<N�<Vr�<Ɣ�<���<�ԏ<G�<~�<v)�<2C�<�[�<�s�<h��<���<l}<��y<'�u<��q<�n<�7j<!`f<t�b<q�^<�Z<�W<1S<�]O</�K<�G<��C<�!@<X<<��8<�4<v
1<L-<E�)<Q�%<{'"<y<)�<e*<�<�<�\<�<tG<��<��;��;7��;�;3c�;j��;D+�;���;n<�;���;4��;?i�;)L�;�D�;.S�;�w�;=��;5�;ln�;��;���;�hv;��k;\�a;.�W;)�M;_�C;yS:;
�0;�';]�;��;[�;�P;���:��:F��:��:�Ӷ:A�:��:Ј:��s:?{V:#�9:��:ު :r��9d�9��79ܪ�8n��X���Qq�}���,�߹s	�V�"��;���T�Cum�y���:��&`��Pt��y���n��yW˺r4׺�I��w�����#�����T���M� �]�%��+��B1�!�6��<��^B�[H�e�M��lS��Y�n�^�ud��!j�m�o��{u�~({��j���A��%��q����ȋ�Ǡ���y���S��.��{	���  �  �=l(=��=wp=3=��=[=9� =&� =�C =y��<��<�T�<���<���<��<O^�<.��<O��<��<.]�<���<h��<�<�M�< ��<w��<��<,,�<�`�<���<��<��<b#�<P�<�z�<��<��<8��<�<�3�<�Q�<�m�<���<ל�<?��<u��<���<a��<���<���<���<���<.��<w��<^��<��<��<Kf�<�B�<��<��<g��<V��<�D�<��<g��<k�<F�<x��<^�<���<��<r�<7��<�+�<\��<�#�<��<�<q�< ֶ<Q6�<ё�<��<�;�<܉�<2Ԭ<��<-]�<3��<�ץ<2�<�E�<�w�<���<�Ԝ<^��<�'�<N�<_r�<攓<���<�ԏ<M�<�<j)�<'C�<�[�<�s�<~��<y��<l}<ٕy<��u<��q<�n<�7j<�_f<T�b<,�^<��Z<\W<�0S<�]O<�K<?�G<��C<�!@<�W<<��8<�4<z
1<IL-<]�)<��%<�'"<,y<}�<�*<:�<'�<"]<6�<�G<��<��;��;���; �;6c�;���;+�;L��;o<�;t��;��;�h�;�K�;YD�;�R�;�w�;���;�;�m�;q�;���;ehv;��k;r�a;��W;��M;�C;hS:;y�0;ޭ';��;��;}�;�Q;Ϸ�:��:ӽ�:3��:�ն:rB�:j�:9ш:��s:�zV:�9:0�:�� :&��9c�9J�79Ѧ�83���u���dq�������߹\v	���"�1�;�t�T� ym�����;���_��&s��4y��o���X˺p4׺�����Q�����-��\�����L�� ���%���+��A1���6�3�<��^B�UH�˾M�HmS��Y�/�^�ntd�V"j���o�|u�,){�Sk��fB��c����ȋ�P���0z���S��h.���	���  �  �=[(=z�=vp=6=ȷ=%[=C� =)� =�C =���<��<�T�<��<���<��<p^�<H��<c��<��<0]�<Ϛ�<��<�<�M�<!��<W��<i��<,�<�`�<z��<���<���<O#�<�O�<�z�<���<��<��<�<�3�<�Q�<�m�<���<Ҝ�<=��<{��<���<t��<���<���<���<��<P��<��<x��<��<��<mf�<C�<��< ��<o��<j��<�D�<��<e��<k�<�<j��<�]�<���<ߍ�<T�<��<v+�<>��<�#�<<��<�p�<�ն<16�<���<��<f;�<ډ�<4Ԭ<��<C]�<G��<�ץ<I�<�E�<x�<���<�Ԝ<��<�'�<-N�<�r�<���<���<�ԏ<^�<��<~)�<,C�<�[�<~s�<W��<n��<�k}<��y<׾u<K�q<mn<�7j<�_f<�b<��^<��Z<2W<�0S<�]O<�K<��G<��C<�!@<�W<<��8<<�4<�
1<UL-<��)<��%<�'"<fy<��<�*<U�<m�<Z]<a�<�G<��<Q��;V��;5��;�;Ac�;8��;1+�;��;<�;O��;���;Yh�;�K�;�C�;AR�;/w�;C��;��;�m�;�;{��;"hv;�k;P�a;��W;�M;��C;
T:;��0;^�';Ś;Y�;��;R;���:��:7��:^��:L׶:D�:��:�ш:�s:�}V:��9:3�:�� :f��9&`�9��795��8A�����qq�������߹�y	���"���;��T�]zm�c���<���`���u��1y���n���W˺�2׺�㺞��Ă��L�t��F������K�4 ��%���+�hA1���6���<�^B��H�*�M�mS��Y���^��ud��"j�w�o��|u��){��k���B�����g�2ɋ������z��T���.���	���  �  
�=T(={�=sp=9=η=$[=M� =5� =�C =���<�<�T�<-��<���<�<�^�<e��<���<��<G]�<��<|��<(�<�M�<!��<U��<[��<,�<d`�<U��<���<���<#�<�O�<�z�<���<���<���<��<~3�<�Q�<m�<���<ڜ�</��<���<���<}��<���<���<���<��<���<���<���<:��<9��<�f�<C�<��<=��<���<s��<�D�<��<V��<k�<�<Y��<�]�<���<���<&�<���<:+�<��<�#�<���<��<�p�<�ն<6�<���<��<b;�<ۉ�<(Ԭ<��<=]�<T��<�ץ<p�<�E�<x�<觞<�Ԝ<���<
(�<bN�<�r�<��<ٵ�<�ԏ<r�<��<�)�<6C�<�[�<�s�<J��<g��<�k}<l�y<�u<�q<+n<7j<P_f<��b<��^<^�Z<�W<v0S<f]O<�K<ݻG<��C<�!@<X<<Ґ8<9�4<�
1<�L-<��)<��%<2("<�y<��<P+<��<��<�]<��<.H<*�<���;U��;���;�;Qc�;=��;+�;��;�;�;���;���;�g�;�J�;C�;�Q�;Mv�;б�;�;Bm�;��;��;�gv;��k;��a;/�W;c�M;�C;^T:;��0;Q�';�;��;��;�S;k��:��:��:Z��:�ض:IF�:��:$ӈ:��s: ~V:��9:��:W� :ԃ�9�\�9%�79�i�8��������q����2๢�	�l�"�?�;�G�T��~m�U���=���a���u���x��To���V˺/3׺��?��4���G����i��{��J�� �u�%��+��@1�a�6�$�<�{]B��H��M��lS��Y�x�^�vd��"j�w�o��}u�+{�5l��NC������ʋ�K���{���T��9/��}
���  �  ��=N(=u�=lp=;=ӷ=1[=\� =F� =�C =���<4�<U�<f��<-��<G�<�^�<���<���<��<j]�<���<���<5�<�M�<��<P��<D��<�+�<V`�<6��<���<���<�"�<�O�<�z�<���<���<���<��<n3�<�Q�<\m�<���<Ɯ�<,��<���<���<���<
��<���<��<O��<���<���<״�<i��<k��<�f�<IC�<��<W��<���<���<E�<
�<S��<k�<	�<6��<�]�<���<���<��<Ǧ�<+�<ݩ�<V#�<���<��<�p�<�ն<�5�<���<��<[;�<É�<&Ԭ<��<P]�<q��<إ<��<�E�<Mx�< ��<!՜<���<A(�<�N�<�r�<@��<���<�ԏ<��<��<�)�<?C�<�[�<ts�<D��<A��<gk}<D�y<%�u<��q<�n<�6j<�^f<\�b<H�^<��Z<�W<E0S<>]O<��K<ŻG<��C<�!@<X<<�8<m�4<1<�L-<)�)<K�%<~("<z<f�<�+<�<�<�]<�<`H<v�<+��;���;���;%�;c�;7��;�*�;e��;o;�;W��;r��;Cg�;J�;�B�;�P�;�u�;*��;X�;�l�;\�;���;�fv;��k;�a;-�W;�M;R�C;qU:;��0;O�';L�;��;X�;U;���:��:L��:��:�۶:�H�:m�:6Ո:p�s:cV:߅9:��:˨ :���9�T�9��79�Z�8 Z��8��{�q������p�	���"� �;���T�h�m�"	��,@��yc���u��:z��Ho���U˺�1׺� �3���~����*���������H�, �a�%�-�+�?1��6��<�y\B��H���M��lS�;Y���^�?vd�$j�2�o�d~u��,{�m��D��M���򈻰ʋ�����{��xU���/���
���  �  �=F(=n�=pp=>=׷=>[=d� =Z� =D =��<j�<HU�<���<N��<��<�^�<͟�<���<�<�]�<��<���<3�<�M�<��<?��<5��<�+�<)`�<��<���<g��<�"�<iO�<Bz�<g��<���<���<��<93�<�Q�<Gm�<n��<���<7��<���<���<���<��<��<&��<���<���<��<��<���<���<�f�<C�<�<��<���<���<E�< �<Z��<�j�<��< ��<�]�<X��<]��<��<���<�*�<���<#�<R��<X�<hp�<oն<�5�<c��<��<B;�<���<0Ԭ<��<c]�<|��<5إ<��<F�<�x�<4��<]՜<���<x(�<�N�<s�<t��<��<&Տ<��<��<�)�<BC�<�[�<is�<0��<(��<%k}<��y<�u<V�q<an<s6j<e^f<��b<�^<��Z<<W<�/S<�\O<a�K<��G<��C<�!@<X<<��8<��4<)1<M-<k�)<��%<�("<�z<��<�+<��<��<s^<\�<�H<��<m��;.��;���;f�;3c�;��;�*�;��;�:�;���;���;�f�;fI�;�A�; P�;u�;]��;��;	l�;��;D��;8fv;V�k;�a;��W;ۧM;��C;$V:;K�0;��';"�;l�;��;�V;���:;!�:��:��:F߶:�J�:��:�ֈ:��s:�V:�9:��:� :f~�9P�9i�79�&�8��������q������"�^�	���"���;�M�T�P�m�1���A��cd��w��,z��un��UV˺y0׺���?��m|����f����ƀ��G�p	 ���%���+��=1���6�ݨ<�\B��H�L�M�rlS��Y�J�^��vd��$j�7�o��u��-{��m���D�� ����lˋ�ѣ���|�� V��Y0��T���  �  �=8(=k�=lp=;=޷=G[=q� =l� = D ='��<��<yU�<ј�<���<��<._�<���<���<N�<�]�<%��<���<=�<�M�<��<1��<��<�+�<`�<��<P��<5��<�"�<3O�<z�<*��<M��<g��<m�<3�<eQ�<7m�<X��<Ɯ�<+��<���<���<���<7��<8��<R��<���<
��<D��<=��<̟�<Ӆ�<'g�<�C�<)�<���<Ϻ�<���<.E�<�<M��<�j�<��<
��<y]�<+��<=��<��<Z��<�*�<p��<�"�<��<$�<+p�<Sն<�5�<N��<r�<-;�<���<!Ԭ<��<v]�<���<Sإ<��<(F�<�x�<i��<�՜<< �<�(�<�N�<5s�<���<B��<QՏ<��<��<�)�<>C�<�[�<is�<��<��<�j}<��y<��u<��q<�n<�5j<!^f<��b<v�^<0�Z<�W<�/S<�\O<B�K<h�G<��C<�!@<X<<�8<��4<]1<gM-<͒)<��%<K)"<�z<D�<�,<��<��<�^<��<I<�<ߛ�;���;��;P�;9c�;ܽ�;A*�;��;;:�;H��;0��;�e�;�H�;
A�;�O�;.t�;���;��;�k�;�;؃�;�ev;��k;6�a;C�W;�M;��C;�V:;+�0;8�';��;��;��;iX;:��: %�:��:r��:��:BM�:=��:f؈:�s:�V:ǅ9:��:�� :Cy�9�K�9�t79���8�g���	�,�q��Ĭ�?,๊�	�?�"���;�c�T�^�m�����B���e��0x��$z��)o���U˺/׺d��<��y����-��@��^��E�� ��%��+�o<1��6���<�4[B�~H�ȼM��lS�TY�Q�^��wd�I%j�N�o��u��.{��n���E�����b�]̋�����i}���V���0������  �  ԃ=,(=g�=kp=B=�=N[=�� =u� =-D =P��<��<�U�<���<���<��<]_�<)��<&��<^�<�]�<K��<���<N�<�M�<��<)��<���<�+�<�_�<͒�<��<��<`"�<�N�<�y�<��<2��<4��<=�<�2�<EQ�<m�<D��<���<*��<���<���<���<[��<D��<x��<���<7��<o��<d��<���<���<Rg�<�C�<R�<���<��<̂�<+E�<�<J��<�j�<��<��<U]�<��<��<X�<:��<a*�<=��<�"�<喻<�<�o�<+ն<y5�<(��<M�<";�<���<"Ԭ<��<t]�<���<jإ<��<VF�<�x�<���<�՜<j �<�(�<O�<es�<���<`��<_Տ<��<��<�)�<OC�<�[�<]s�< ��<���<�j}<j�y</�u<��q<�n<�5j<�]f<�b<7�^<��Z<yW<l/S<c\O<�K<7�G<w�C<�!@<*X<<#�8<��4<�1<�M-<�)<I�%<�)"<Q{<��<�,<L�<`�<7_<�<EI<=�<���;���;S��;}�; c�;ƽ�;�)�;k��;�9�;���;q��;ge�;H�;:@�;�N�;Vs�;>��;4�;�j�;��;`��;�dv;0�k;��a;M�W;��M;��C;�W:;Z�0;��';Р;׶;�;�Y;���:�'�:���:H��:h�:�O�:(��:�ڈ:��s:��V:]�9:��:�� :�u�9�C�9ld79O�8v���,	���q�Ҭ�8��	���"��;���T�֐m����E���g���x���z���n���T˺/׺ �⺩��1x��8����ڳ�+~�	D�� ���%���+�7;1�.�6��<�ZB��H���M�lS�[Y���^�exd�5&j�d�o�ǁu�R0{�Ao��)F��������D͋�'���	~��}W��?1��s���  �  ʃ=-(=`�=ip=D=�=U[=�� =�� =AD =}��<��<�U�<0��<���<�<|_�<G��<Q��<��<�]�<R��<���<H�<�M�<���<#��<���<�+�<�_�<���<��<���<+"�<�N�<�y�<ʢ�<���<��<�<�2�</Q�<	m�<G��<���<3��<���<���<���<n��<d��<���<��<T��<���<���<$��<2��<pg�<�C�<t�<���<��<؂�<-E�<	�<T��<�j�<��<ټ�<>]�<���<��<B�<���<3*�<
��<|"�<���<��<�o�<�Զ<Z5�<��<B�<;�<���<,Ԭ<��<|]�<���<�إ<
�<{F�<�x�<���<�՜<� �<)�<LO�<�s�<앓<���<�Տ<��< �<�)�<QC�<�[�<Ns�<��<Ꟁ<lj}<�y<��u<I�q<Ln<55j<_]f<��b<ʮ^<��Z<DW<	/S<0\O<܊K<;�G<\�C<�!@<1X<< �8<��4<�1<�M-<R�)<��%<�)"<�{<�<=-<Ǎ<��<w_<a�<�I<��<���;��;K��;��;c�;���;�)�;(��;d9�;/��;%��;�d�;<G�;�?�;&N�;�r�;W��;� �;oj�;�;��;�dv;W�k;F�a;��W;��M;��C;X:;��0;��';��;e�;�;w[;��:�*�:.��:G��:B�:-R�::��:�ۈ:��s:��V:�9:�:ä :�u�9�@�9`Z79�Ö8����6	��q��ܬ��C๠�	���"�q�;�N�T�.�m�i��KF��=h���x���{��n��U˺g.׺z�����u��������R|��B�� ��%���+��91���6��<��YB�eH���M�	lS�FY�(�^�Jxd��&j��o�9�u�<1{��o��G��u�������͋������~���W��2������  �  ��="(=W�=fp=E=�=d[=�� =�� =GD =���<�<�U�<K��<��<-�<�_�<c��<b��<��<�]�<]��<���<R�<�M�<���<��<���<|+�<�_�<���<���<���<"�<�N�<�y�<â�<���<	��<�<�2�<+Q�<�l�</��<���</��<���<��<���<}��<���<���<��<o��<���<���<?��<D��<�g�<D�<~�<���<��<��<ZE�<�<Q��<�j�<��<ü�<4]�<���<͌�<*�<ӥ�<+*�<騾<`"�<���<��<�o�<�Զ<J5�<��<-�<;�<���<,Ԭ<��<�]�<�<�إ<!�<�F�<y�<ʨ�<֜<� �<")�<_O�<�s�<��<���<�Տ<��<�<�)�<PC�<�[�<=s�<쉂<ӟ�<fj}<ٓy<μu<�q<n<5j<]f<��b<��^<N�Z<W<�.S<&\O<��K<�G<6�C<�!@<5X<<Q�8<<�4<�1<N-<k�)<��%<)*"<�{<B�<s-<��<��<�_<��<�I<��<ߜ�;���;{��;��;�b�;p��;�)�;��;G9�;���;斺;d�;G�;L?�;�M�;�r�;ѭ�;� �;j�;��;
��;�cv;��k;��a;��W;��M;@�C;�X:;|�0;��';W�;Q�;��;\;���:t,�:j��:���:�:�R�:��:�܈:e�s:N�V:��9:��:� :Vo�9�;�9rV79��8���@	��r�%ެ��K�š	�#�"���;���T�q�m�:��G��ni��Tz��|���m���T˺z+׺���ͼ�qt����������{��A� �w�%��+��81���6�?�<�:YB��
H���M�lS�rY���^�yd��'j�1�o��u��1{�0p���G�����s���΋�u���$��,X��i2������  �  ��=!(=`�=kp=C=�=[[=�� =�� =RD =���<�<	V�<\��<)��<=�<�_�<y��<z��<��<^�<i��<���<L�<�M�<��<��<���<u+�<�_�<u��<���<���<"�<�N�<~y�<���<���<���<��<�2�<Q�<�l�</��<���</��<���<���<���<���<���<���<#��<���<���<ϵ�<`��<[��<�g�<D�<��<���<#��<��<?E�<�<H��<�j�<��<¼�<]�<���<���<�<ϥ�<�)�<Ũ�<:"�<���<��<�o�<�Զ<+5�<���<-�<;�<���<Ԭ<��<�]�<ʜ�<�إ<(�<�F�<&y�<�<֜<� �<5)�<zO�<�s�<��<���<�Տ<�<	�<�)�<PC�<�[�<Qs�<쉂<ԟ�<6j}<��y<��u<��q<�n<�4j<�\f<N�b<r�^<,�Z<�W<�.S<�[O<��K<�G<Z�C<�!@<*X<<9�8<�4<�1<N-<��)<��%<a*"<|<e�<�-<�<0�<�_<��<�I<��<��;D��;i��;��;/c�;���;�)�;ۧ�;�8�;���;h��;d�;�F�;�>�;#M�;r�;ƭ�; �;�i�;y�;���;�cv;��k;��a;��W;��M;��C;�X:;�0;��';T�;}�;��;�\;���:�.�:���:;��:m�:�T�:B��:ވ:��s:�V:�9:�:'� :Hp�9�;�9tL79x��8 Z��-R	��	r��謹�S�A�	���"�Q�;��T���m����G��Gi���y��{���n���T˺-׺\��ֻ��s����)��Ͱ�{��@�w ���%��~+��81���6�-�<��XB�H��M�lS�/Y��^�yd��'j���o�~�u��2{��p���G��R�������΋�����e���X���2��S���  �  ��=(=T�=cp=F=�=a[=�� =�� =[D =���<�<
V�<T��<*��<2�<�_�<h��<���<��<^�<}��<���<k�<�M�<��<��<���<q+�<�_�<���<���<���<�!�<�N�<�y�<���<���<���<��<�2�<Q�<�l�<��<���<$��<���<���<
��<���<t��<���<��<���<���<ȵ�<Z��<X��<�g�<D�<��<���<*��<���<=E�<(�<B��<�j�<��<���<]�<���<Ì�<��<̥�<�)�<稾<P"�<i��<��<�o�<�Զ<*5�<<�<�:�<���<Ԭ<��<�]�<ߜ�<�إ<&�<�F�<y�<���<֜<� �<.)�<|O�<�s�<��<���<�Տ<!�<�<�)�<YC�<�[�<8s�<։�<ҟ�<j}<Гy<��u<��q<�n<�4j<+]f<G�b<Z�^<�Z<�W<�.S<�[O<��K<ݺG<*�C<�!@<7X<<b�8<-�4<1<�M-<��)<��%<L*"<|<U�<�-<
�<0�<�_<��<�I<��<f��;`��;���;��;�b�;F��;C)�;̧�;�8�;���;T��;�c�;\F�;�>�;�M�;�q�;���;���;�i�;��;���;�cv;�k;�a;A�W;P�M;��C;#Y:;o�0;F�';�;1�;��;�\;K��:;.�:���:s��:��:SV�:V��:�ވ:M�s:��V:m�9:O�:�� :'k�9(:�9"H79���8�%���W	�5r�+bKไ�	���"�U�;���T��m���(H��Kj��C{��<|���n���R˺�,׺	��z��t��=�������[{��@�� ���%��~+��81�/�6�i�<�XB��
H���M��kS��Y���^��yd��'j�g�o�-�u��2{��p���G��q��F����΋�٦������X��e2������  �  ��=!(=`�=kp=C=�=[[=�� =�� =RD =���<�<	V�<\��<)��<=�<�_�<y��<z��<��<^�<i��<���<L�<�M�<��<��<���<u+�<�_�<u��<���<���<"�<�N�<~y�<���<���<���<��<�2�<Q�<�l�</��<���</��<���<���<���<���<���<���<#��<���<���<ϵ�<`��<[��<�g�<D�<��<���<#��<��<?E�<�<H��<�j�<��<¼�<]�<���<���<�<ϥ�<�)�<Ũ�<:"�<���<��<�o�<�Զ<+5�<���<.�<;�<���<Ԭ<��<�]�<ʜ�<�إ<(�<�F�<&y�<�<֜<� �<5)�<zO�<�s�<��<���<�Տ<�<	�<�)�<PC�<�[�<Qs�<쉂<ԟ�<6j}<��y<��u<��q<�n<�4j<�\f<N�b<r�^<,�Z<�W<�.S<�[O<��K<�G<Z�C<�!@<*X<<9�8<�4<�1<N-<��)<��%<a*"<|<e�<�-<�<0�<�_<��<�I<��<��;D��;i��;��;/c�;���;�)�;ۧ�;�8�;���;h��;d�;�F�;�>�;#M�;r�;ƭ�; �;�i�;y�;���;�cv;��k;��a;��W;��M;��C;�X:;�0;��';T�;}�;��;�\;���:�.�:���:;��:m�:�T�:B��:ވ:��s:�V:�9:�:'� :Hp�9�;�9tL79x��8 Z��-R	��	r��謹�S�A�	���"�Q�;��T���m����G��Gi���y��{���n���T˺-׺\��ֻ��s����)��Ͱ�{��@�w ���%��~+��81���6�-�<��XB�H��M�lS�/Y��^�yd��'j���o�~�u��2{��p���G��R�������΋�����e���X���2��S���  �  ��="(=W�=fp=E=�=d[=�� =�� =GD =���<�<�U�<K��<��<-�<�_�<c��<b��<��<�]�<]��<���<R�<�M�<���<��<���<|+�<�_�<���<���<���<"�<�N�<�y�<â�<���<	��<�<�2�<+Q�<�l�</��<���</��<���<��<���<}��<���<���<��<o��<���<���<?��<D��<�g�<D�<~�<���<��<��<ZE�<�<Q��<�j�<��<ü�<4]�<���<͌�<*�<ӥ�<+*�<騾<`"�<���<��<�o�<�Զ<J5�<��<-�<;�<���<,Ԭ<��<�]�<�<�إ<!�<�F�<y�<ʨ�<֜<� �<")�<_O�<�s�<��<���<�Տ<��<�<�)�<PC�<�[�<=s�<쉂<ӟ�<fj}<ٓy<μu<�q<n<5j<]f<��b<��^<N�Z<W<�.S<&\O<��K<�G<6�C<�!@<5X<<Q�8<<�4<�1<N-<k�)<��%<)*"<�{<B�<s-<��<��<�_<��<�I<��<ߜ�;���;{��;��;�b�;p��;�)�;��;G9�;���;斺;d�;G�;L?�;�M�;�r�;ѭ�;� �;j�;��;
��;�cv;��k;��a;��W;��M;@�C;�X:;|�0;��';W�;Q�;��;\;���:t,�:j��:���:�:�R�:��:�܈:e�s:N�V:��9:��:� :Vo�9�;�9rV79��8���@	��r�%ެ��K�š	�#�"���;���T�q�m�:��G��ni��Tz��|���m���T˺z+׺���ͼ�qt����������{��A� �w�%��+��81���6�?�<�:YB��
H���M�lS�rY���^�yd��'j�1�o��u��1{�0p���G�����s���΋�u���$��,X��i2������  �  ʃ=-(=`�=ip=D=�=U[=�� =�� =AD =}��<��<�U�<0��<���<�<|_�<G��<Q��<��<�]�<R��<���<H�<�M�<���<#��<���<�+�<�_�<���<��<���<+"�<�N�<�y�<ʢ�<���<��<�<�2�</Q�<	m�<G��<���<3��<���<���<���<n��<d��<���<��<T��<���<���<$��<2��<pg�<�C�<t�<���<��<؂�<-E�<	�<T��<�j�<��<ټ�<>]�<���<��<B�<���<3*�<
��<|"�<���<��<�o�<�Զ<Z5�<��<B�<;�<���<,Ԭ<��<|]�<���<�إ<
�<{F�<�x�<���<�՜<� �<)�<LO�<�s�<앓<���<�Տ<��<��<�)�<QC�<�[�<Ns�<��<Ꟁ<lj}<�y<��u<I�q<Ln<55j<_]f<��b<ʮ^<��Z<DW<	/S<0\O<܊K<;�G<\�C<�!@<1X<< �8<��4<�1<�M-<R�)<��%<�)"<�{<�<=-<Ǎ<��<w_<a�<�I<��<���;��;K��;��;c�;���;�)�;(��;d9�;/��;%��;�d�;<G�;�?�;&N�;�r�;W��;� �;oj�;�;��;�dv;W�k;F�a;��W;��M;��C;X:;��0;��';��;e�;�;w[;��:�*�:.��:G��:B�:-R�::��:�ۈ:��s:��V:�9:�:ä :�u�9�@�9`Z79�Ö8����6	��q��ܬ��C๠�	���"�q�;�N�T�.�m�i��KF��=h���x���{��n��U˺g.׺z�����u��������R|��B�� ��%���+��91���6��<��YB�eH���M�	lS�FY�(�^�Jxd��&j��o�9�u�<1{��o��G��u�������͋������~���W��2������  �  ԃ=,(=g�=kp=B=�=N[=�� =u� =-D =P��<��<�U�<���<���<��<]_�<)��<&��<^�<�]�<K��<���<N�<�M�<��<)��<���<�+�<�_�<͒�<��<��<`"�<�N�<�y�<��<2��<4��<=�<�2�<EQ�<m�<D��<���<*��<���<���<���<[��<D��<x��<���<7��<o��<d��<���<���<Rg�<�C�<R�<���<��<̂�<+E�<�<J��<�j�<��<��<U]�<��<��<X�<:��<a*�<=��<�"�<喻<�<�o�<+ն<y5�<(��<M�<";�<���<"Ԭ<��<t]�<���<jإ<��<VF�<�x�<���<�՜<j �<�(�<O�<es�<���<`��<_Տ<��<��<�)�<OC�<�[�<]s�< ��<���<�j}<j�y</�u<��q<�n<�5j<�]f<�b<7�^<��Z<yW<l/S<c\O<�K<7�G<w�C<�!@<*X<<#�8<��4<�1<�M-<�)<I�%<�)"<Q{<��<�,<L�<`�<7_<�<EI<=�<���;���;S��;}�; c�;ƽ�;�)�;k��;�9�;���;q��;ge�;H�;:@�;�N�;Vs�;>��;4�;�j�;��;`��;�dv;0�k;��a;M�W;��M;��C;�W:;Z�0;��';Р;׶;�;�Y;���:�'�:���:H��:h�:�O�:(��:�ڈ:��s:��V:]�9:��:�� :�u�9�C�9ld79O�8v���,	���q�Ҭ�8��	���"��;���T�֐m����E���g���x���z���n���T˺/׺ �⺩��1x��8����ڳ�+~�	D�� ���%���+�7;1�.�6��<�ZB��H���M�lS�[Y���^�exd�5&j�d�o�ǁu�R0{�Ao��)F��������D͋�'���	~��}W��?1��s���  �  �=8(=k�=lp=;=޷=G[=q� =l� = D ='��<��<yU�<ј�<���<��<._�<���<���<N�<�]�<%��<���<=�<�M�<��<1��<��<�+�<`�<��<P��<5��<�"�<3O�<z�<*��<M��<g��<m�<3�<eQ�<7m�<X��<Ɯ�<+��<���<���<���<7��<8��<R��<���<
��<D��<=��<̟�<Ӆ�<'g�<�C�<)�<���<Ϻ�<���<.E�<�<M��<�j�<��<
��<y]�<+��<=��<��<Z��<�*�<p��<�"�<��<$�<+p�<Sն<�5�<N��<r�<-;�<���<!Ԭ<��<v]�<���<Sإ<��<(F�<�x�<i��<�՜<< �<�(�<�N�<5s�<���<B��<QՏ<��<��<�)�<>C�<�[�<is�<��<��<�j}<��y<��u<��q<�n<�5j<!^f<��b<v�^<0�Z<�W<�/S<�\O<B�K<h�G<��C<�!@<X<<�8<��4<]1<gM-<͒)<��%<K)"<�z<D�<�,<��<��<�^<��<I<�<ߛ�;���;��;P�;9c�;ܽ�;A*�;��;;:�;H��;0��;�e�;�H�;	A�;�O�;.t�;���;��;�k�;�;؃�;�ev;��k;6�a;C�W;�M;��C;�V:;+�0;8�';��;��;��;iX;:��: %�:��:r��:��:BM�:=��:f؈:�s:�V:ǅ9:��:�� :Cy�9�K�9�t79���8�g���	�,�q��Ĭ�?,๊�	�?�"���;�c�T�^�m�����B���e��0x��$z��)o���U˺/׺d��<��y����-��@��^��E�� ��%��+�o<1��6���<�4[B�~H�ȼM��lS�TY�Q�^��wd�I%j�N�o��u��.{��n���E�����b�]̋�����i}���V���0������  �  �=F(=n�=pp=>=׷=>[=d� =Z� =D =��<j�<HU�<���<N��<��<�^�<͟�<���<�<�]�<��<���<3�<�M�<��<?��<5��<�+�<)`�<��<���<g��<�"�<iO�<Bz�<g��<���<���<��<93�<�Q�<Gm�<n��<���<7��<���<���<���<��<��<&��<���<���<��<��<���<���<�f�<C�<�<��<���<���<E�< �<Z��<�j�<��< ��<�]�<X��<]��<��<���<�*�<���<#�<R��<X�<hp�<oն<�5�<c��<��<B;�<���<0Ԭ<��<c]�<|��<5إ<��<F�<�x�<4��<]՜<���<x(�<�N�<s�<t��<��<&Տ<��<��<�)�<BC�<�[�<is�<0��<(��<%k}<��y<�u<V�q<an<s6j<e^f<��b<�^<��Z<<W<�/S<�\O<b�K<��G<��C<�!@<X<<��8<��4<)1<M-<k�)<��%<�("<�z<��<�+<��<��<s^<\�<�H<��<m��;.��;���;f�;3c�;��;�*�;��;�:�;���;���;�f�;fI�;�A�; P�;u�;]��;��;	l�;��;D��;8fv;V�k;�a;��W;ۧM;��C;#V:;K�0;��';"�;l�;��;�V;���:;!�:��:��:F߶:�J�:��:�ֈ:��s:�V:�9:��:� :f~�9P�9i�79�&�8��������q������"�^�	���"���;�M�T�P�m�1���A��cd��w��,z��un��UV˺y0׺���?��m|����f����ƀ��G�p	 ���%���+��=1���6�ݨ<�\B��H�L�M�rlS��Y�J�^��vd��$j�7�o��u��-{��m���D�� ����lˋ�ѣ���|�� V��Y0��T���  �  ��=N(=u�=lp=;=ӷ=1[=\� =F� =�C =���<4�<U�<f��<-��<G�<�^�<���<���<��<j]�<���<���<5�<�M�<��<P��<D��<�+�<V`�<6��<���<���<�"�<�O�<�z�<���<���<���<��<n3�<�Q�<\m�<���<Ɯ�<,��<���<���<���<
��<���<��<O��<���<���<״�<i��<k��<�f�<IC�<��<W��<���<���<E�<
�<S��<k�<	�<6��<�]�<���<���<��<Ǧ�<+�<ݩ�<V#�<���<��<�p�<�ն<�5�<���<��<[;�<É�<&Ԭ<��<P]�<q��<إ<��<�E�<Mx�< ��<!՜<���<A(�<�N�<�r�<@��<���<�ԏ<��<��<�)�<?C�<�[�<ts�<D��<A��<gk}<D�y<%�u<��q<�n<�6j<�^f<\�b<H�^<��Z<�W<E0S<>]O<��K<ŻG<��C<�!@<X<<�8<m�4<1<�L-<)�)<K�%<~("<z<f�<�+<�<�<�]<�<`H<v�<+��;���;���;%�;c�;7��;�*�;e��;n;�;W��;r��;Cg�;J�;�B�;�P�;�u�;)��;W�;�l�;\�;���;�fv;��k;�a;-�W;�M;R�C;qU:;��0;O�';L�;��;X�;U;���:��:L��:��:�۶:�H�:m�:6Ո:p�s:cV:߅9:��:˨ :���9�T�9��79�Z�8 Z��8��{�q������p�	���"� �;���T�h�m�"	��,@��yc���u��:z��Ho���U˺�1׺� �3���~����*���������H�, �a�%�-�+�?1��6��<�y\B��H���M��lS�;Y���^�?vd�$j�2�o�d~u��,{�m��D��M���򈻰ʋ�����{��xU���/���
���  �  
�=T(={�=sp=9=η=$[=M� =5� =�C =���<�<�T�<-��<���<�<�^�<e��<���<��<G]�<��<|��<(�<�M�<!��<U��<[��<,�<d`�<U��<���<���<#�<�O�<�z�<���<���<���<��<~3�<�Q�<m�<���<ڜ�</��<���<���<}��<���<���<���<��<���<���<���<:��<9��<�f�<C�<��<=��<���<s��<�D�<��<V��<k�<�<Y��<�]�<���<���<&�<���<:+�<��<�#�<���<��<�p�<�ն<6�<���<��<b;�<ۉ�<(Ԭ<��<=]�<T��<�ץ<p�<�E�<x�<觞<�Ԝ<���<
(�<bN�<�r�<��<ٵ�<�ԏ<r�<��<�)�<6C�<�[�<�s�<J��<g��<�k}<l�y<�u<�q<+n<7j<P_f<��b<��^<^�Z<�W<v0S<f]O<�K<ݻG<��C<�!@<X<<Ґ8<9�4<�
1<�L-<��)<��%<2("<�y<��<P+<��<��<�]<��<.H<*�<���;U��;���;�;Qc�;=��;+�;��;�;�;���;���;�g�;�J�;C�;�Q�;Mv�;б�;�;Bm�;��;��;�gv;��k;��a;.�W;c�M;�C;^T:;��0;Q�';�;��;��;�S;k��:��:��:Z��:�ض:IF�:��:$ӈ:��s: ~V:��9:��:W� :ԃ�9�\�9%�79�i�8��������q����2๢�	�l�"�?�;�G�T��~m�U���=���a���u���x��To���V˺/3׺��?��4���G����i��{��J�� �u�%��+��@1�a�6�$�<�{]B��H��M��lS��Y�x�^�vd��"j�w�o��}u�+{�5l��NC������ʋ�K���{���T��9/��}
���  �  �=[(=z�=vp=6=ȷ=%[=C� =)� =�C =���<��<�T�<��<���<��<p^�<H��<c��<��<0]�<Ϛ�<��<�<�M�<!��<W��<i��<,�<�`�<z��<���<���<O#�<�O�<�z�<���<��<��<�<�3�<�Q�<�m�<���<Ҝ�<=��<{��<���<t��<���<���<���<��<P��<��<x��<��<��<mf�<C�<��< ��<o��<j��<�D�<��<e��<k�<�<j��<�]�<���<ߍ�<T�<��<v+�<>��<�#�<<��<�p�<�ն<16�<���<��<f;�<ډ�<4Ԭ<��<C]�<G��<�ץ<I�<�E�<x�<���<�Ԝ<��<�'�<-N�<�r�<���<���<�ԏ<^�<��<~)�<,C�<�[�<~s�<W��<n��<�k}<��y<׾u<K�q<mn<�7j<�_f<�b<��^<��Z<2W<�0S<�]O<�K<��G<��C<�!@<�W<<��8<<�4<�
1<UL-<��)<��%<�'"<fy<��<�*<U�<m�<Z]<a�<�G<��<Q��;V��;5��;�;Ac�;8��;1+�;��;<�;O��;���;Yh�;�K�;�C�;@R�;/w�;C��;��;�m�;�;{��;"hv;�k;P�a;��W;�M;��C;
T:;��0;^�';Ś;Y�;��;R;���:��:7��:^��:L׶:D�:��:�ш:�s:�}V:��9:3�:�� :f��9&`�9��795��8A�����qq�������߹�y	���"���;��T�]zm�c���<���`���u��1y���n���W˺�2׺�㺞��Ă��L�t��F������K�4 ��%���+�hA1���6���<�^B��H�*�M�mS��Y���^��ud��"j�w�o��|u��){��k���B�����g�2ɋ������z��T���.���	���  �  �=l(=��=wp=3=��=[=9� =&� =�C =y��<��<�T�<���<���<��<O^�<.��<O��<��<.]�<���<h��<�<�M�< ��<w��<��<,,�<�`�<���<��<��<b#�<P�<�z�<��<��<8��<�<�3�<�Q�<�m�<���<ל�<?��<u��<���<a��<���<���<���<���<.��<w��<^��<��<��<Kf�<�B�<��<��<g��<V��<�D�<��<g��<k�<F�<x��<^�<���<��<r�<7��<�+�<\��<�#�<��<�<q�< ֶ<Q6�<ё�<��<�;�<܉�<2Ԭ<��<-]�<3��<�ץ<2�<�E�<�w�<���<�Ԝ<^��<�'�<N�<_r�<攓<���<�ԏ<M�<�<j)�<'C�<�[�<�s�<~��<y��<l}<ٕy<��u<��q<�n<�7j<�_f<T�b<,�^<��Z<\W<�0S<�]O<�K<?�G<��C<�!@<�W<<��8<�4<z
1<IL-<]�)<��%<�'"<,y<}�<�*<:�<'�<"]<6�<�G<��<��;��;���; �;6c�;���;+�;L��;o<�;t��;��;�h�;�K�;YD�;�R�;�w�;���;�;�m�;q�;���;ehv;��k;r�a;��W;��M;�C;hS:;y�0;ޭ';��;��;}�;�Q;Ϸ�:��:ӽ�:3��:�ն:rB�:j�:9ш:��s:�zV:�9:0�:�� :&��9c�9J�79Ѧ�83���u���dq�������߹\v	���"�1�;�t�T� ym�����;���_��&s��4y��o���X˺p4׺�����Q�����-��\�����L�� ���%���+��A1���6�3�<��^B�UH�˾M�HmS��Y�/�^�ntd�V"j���o�|u�,){�Sk��fB��c����ȋ�P���0z���S��h.���	���  �  �=b(=�=tp=9=Ƿ=[=8� =� =�C =[��<��<�T�<Η�<���<��<F^�<��<6��<��<]�<���<g��<�<�M�<!��<g��<r��<?,�<�`�<���<#��<#��<|#�<*P�<{�< ��<D��<F��<.�<�3�<�Q�<�m�<���<֜�<3��<���<���<d��<���<x��<���<���<+��<V��<<��<͞�<���<Jf�<�B�<q�<���<V��<Y��<�D�<��<^��<k�<,�<}��<^�<���<��<|�<^��<�+�<���<�#�<��<'�<q�< ֶ<T6�<味<��<};�<���<6Ԭ<��</]�<3��<�ץ< �<qE�<�w�<���<�Ԝ<<��<�'�<N�<Vr�<Ɣ�<���<�ԏ<G�<~�<v)�<2C�<�[�<�s�<h��<���<l}<��y<'�u<��q<�n<�7j<!`f<t�b<q�^<�Z<�W<1S<�]O</�K<�G<��C<�!@<X<<��8<�4<v
1<L-<E�)<Q�%<{'"<y<)�<e*<�<�<�\<�<tG<��<��;��;7��;�;3c�;j��;D+�;���;n<�;���;4��;?i�;)L�;�D�;.S�;�w�;=��;5�;ln�;��;���;�hv;��k;\�a;.�W;)�M;_�C;yS:;
�0;�';]�;��;[�;�P;���:��:F��:��:�Ӷ:A�:��:Ј:��s:?{V:#�9:��:ު :r��9d�9��79ܪ�8n��X���Qq�}���,�߹s	�V�"��;���T�Cum�y���:��&`��Pt��y���n��yW˺r4׺�I��w�����#�����T���M� �]�%��+��B1�!�6��<��^B�[H�e�M��lS��Y�n�^�ud��!j�m�o��{u�~({��j���A��%��q����ȋ�Ǡ���y���S��.��{	���  �  �=�%=��=(m=~=��=�V=A� =�� =�= =ӿ�<H�<$F�<p��<B��<0�<�K�<M��<D��<f�<�E�<��<7��<���<�0�<�h�<���<C��<�	�<B<�<�m�<���<���<���<w#�<�L�<�s�<��<��</��<���<��<�1�<�H�<�\�<�m�<4|�<4��<���<]��<'��<V��<���<��<Fq�<^�<WG�<�+�<u�<f��<���<��<Z�<� �<���<���<�U�<X�<��<lY�<��<1��< +�<���<�E�<˿<K�<�ż<y;�<��<��<�~�<��<p>�<���<{�<7=�<ۉ�<�Ҫ<��<�Y�<Ɨ�<�ң<�
�<�?�<Zr�<��<�Ϛ<���<�#�<�J�<�o�<,��<մ�<Ս<��<b�<�-�<I�<dc�<�|�<}��<�Z}<�y<��u<��q<�n<@j<�mf<B�b<y�^<��Z<�'W<FXS<�O<��K<��G<�)D<�b@<+�<<�8<�5<�`1<��-<c�)<�@&<G�"<,�<�E<��<<�w<��<�_	<p�<�a<O��;���;�1�;�t�;x��;�,�;��;@)�;��;�o�;�/�;�;��;h�;s��;&�;e�;\��;�$�;ʥ�;�=�;�y;bo;�e;Z�Z;�Q;�AG;k�=;�54;�*;��!;a�;�	;�_;���:M��:�}�:�I�:JS�:���:�$�:M�:0�}:�`:��B:��%:�q	:;��9/Ԣ9�W9=�8�1���ظϩU��5��gӹ3G�@��>6�><O��,h��}��͌�����8���U��vd���cɺ�Vպx;Ẳ�e����R�!0�V�d��E��!u��<%�} +���0��6�$<<��A�׮G�CeM��S���X��^�V7d�g�i�Z�o�iQu�,{�M\���5�����눻+Ƌ�D����}��wZ��C8��9���  �  �=�%=��=$m=�=��=�V=E� =�� =�= =ֿ�<I�<-F�<s��<$��<;�<�K�<V��<C��<Y�<�E�<��<P��<���<�0�<�h�<���</��<y	�<S<�<�m�<���<���<���<�#�<�L�<�s�<��<%��<��<���<��<1�<zH�<�\�<�m�<8|�<J��<��<b��<$��<N��<���<��<Uq�<q^�<?G�<�+�<n�<s��<���<ߍ�<Z�<	!�<���<��<�U�<6�<��<RY�<��<@��<�*�<��<�E�<˿<K�<�ż<p;�<��<��<�~�<��<f>�<���<i�<=�<މ�<�Ҫ<��<�Y�<ʗ�<�ң<�
�<�?�<[r�<��<�Ϛ<���<�#�<�J�<�o�<��<Դ�<Ս<��<q�<�-�<�H�<Fc�<�|�<j��<[}<�y<f�u<�q<Xn<�@j<�mf<N�b<E�^<��Z<�'W<@XS<<�O<��K<��G<�)D<�b@<3�<<.�8<�5<�`1<��-<C�)<�@&<H�"<?�<�E<N�<"<�w<��<�_	<V�<�a<~��;G��;�1�;�t�;,��;S,�;���;)�;���;o�;�/�;��;��;��;���;$&�;�d�;|��;�$�;���;>�;B�y;�ao;�e;C�Z;�Q;�BG;)�=;�54;��*;��!;��;v	;`;���:���:�~�:)I�:T�:���:�$�:��:�}:�`:*�B:��%:Bm	:<��9�͢9��W9��8�����ظ��U�V6��ӹ,E�N��t6��;O�~/h��|���͌�3���9��W��<d��KcɺUպ�:�t����S��/�N���8��$u�_<%�� +���0� �6�.<<���A���G��dM��S���X��^��7d���i�ϝo�\Qu��{�E\��>6��}���ꈻƋ������}���Z��P8������  �  ��=�%=��=)m=~=��=�V=B� =Û =�= =��<P�<9F�<���<7��<^�<�K�<d��<O��<d�<�E�<��<H��<���<�0�<�h�<���<=��<i	�<T<�<�m�<���<���<|��<e#�<L�<�s�<���<*��<���<���<��<w1�<�H�<�\�<n�<)|�<;��<��<d��<6��<R��<���< ��<rq�<�^�<YG�<�+�<h�<���<���<��<Z�<� �<���<��<�U�<4�<"��<PY�<��<@��<�*�<
��<�E�<�ʿ<�J�<�ż<a;�<���<��<~~�<��<U>�<���<{�<=�<艬<�Ҫ<��<�Y�<՗�<�ң<�
�< @�<Xr�<A��<�Ϛ<���<�#�<�J�<�o�<#��<鴏<Ս<��<^�<�-�<I�<Kc�<�|�<^��<�Z}<��y<:�u< �q<9n<i@j<�mf<)�b<(�^<��Z<y'W<XS<0�O<y�K<��G<�)D<�b@<*�<<	�8<�5<�`1<ϧ-<S�)<�@&<X�"<V�<F<v�<i<�w<��<�_	<n�<�a<e��;,��;�1�;u�;E��;�,�;ա�;�(�;���;o�;�/�;��;z�;$�;"��;�%�;�d�;���;0$�;���;�=�;�y;�bo;�e;��Z;lQ;#BG;̦=;�54;��*;��!;~�;]	;a;���:w��:���:�H�:LU�:؞�:�%�:�:F�}:`:.�B:��%:3m	:]��9q͢9zW9w�8!����׸m�U��9�� ӹCI����6�X<O�M3h��|���Ό�|���8���V���c��Vdɺ�Uպ_;Ặ�J����R�4/�`�������;t��;%�i +��0��6��;<���A�<�G�beM��S�`�X�ʃ^��6d�b�i��o��Qu�E{�I\��{6�����{눻[Ƌ�衎��}���Z���8������  �  ��=�%=��=$m=�=��=�V=K� =Ǜ => =���<l�<KF�<���<X��<c�<�K�<}��<_��<�<�E�<���<a��<���<�0�<�h�<���<-��<a	�<><�<�m�<|��<���<u��<X#�<hL�<�s�<��<��<���<���<��<y1�<rH�<�\�<�m�<8|�<\��<��<v��<G��<e��<Ê�<$��<xq�<�^�<nG�<�+�<��<���<���<���<Z�<!�<���<��<�U�</�< ��<MY�<���<*��<�*�<��<�E�<�ʿ<�J�<�ż<W;�<߫�<��<}~�<��<G>�<~��<\�<=�<ቬ<�Ҫ< �<�Y�<���<�ң<�
�<@�<vr�<G��<�Ϛ<���<�#�<�J�<�o�<<��<���<(Ս<��<�<�-�<�H�<=c�<�|�<^��<�Z}<�y<�u<��q<"n<O@j<Wmf<�b<�^<��Z<O'W<XS<��O<p�K<��G<�)D<�b@<3�<<G�8<
5<�`1<�-<��)<�@&<��"<}�<F<��<v<�w<��<`	<��<�a<���;���;2�;u�;B��;1,�;���;�(�;|��;o�;B/�;O�;c�;��;���;�%�;=d�;���;$�;���;�=�;!�y;�ao;�e;��Z;�Q;8CG;��=;�64;�*;^�!;�;�
;;a;���:���:��:K�:�V�:��:�&�:��:�}:,`:J�B:G�%:�l	:I~�9͢9�nW9���8E����$ظ��U�A;���$ӹ�J���e 6��?O�&3h�~��nό�D���:��W���c���bɺ�Sպ:�������7R�q.�l��������s�d;%�l�*���0�6�$;<�O�A���G�]dM��S���X�9�^��7d�c�i��o�Ru��{��\���6������눻�Ƌ�
���u~��%[���8��`���  �  ��=�%=��=&m=}=��=�V=X� =Λ => =��<��<tF�<���<~��<�<�K�<���<u��<��<�E�<��<S��<���<�0�<�h�<���<"��<X	�<<�<�m�<`��<���<F��<4#�<YL�<�s�<Ř�<��<���<���<��<x1�<gH�<�\�<�m�<5|�<N��<��<���<W��<���<ϊ�<O��<�q�<�^�<�G�<�+�<��<���<߼�<��<4Z�<!�<���<���<�U�<?�<���<GY�<���<��<�*�<º�<sE�<�ʿ<�J�<�ż<$;�<ɫ�<{�<e~�<��<:>�<s��<X�<)=�<ω�<�Ҫ<��<�Y�<<ӣ<�<)@�<�r�<a��<�Ϛ<���<�#�<�J�<�o�<[��<��<?Ս<��<x�<�-�<�H�<Lc�<�|�<Z��<�Z}<��y<�u<��q<�n<�?j<Cmf<��b<��^<{�Z<'W<�WS<ȉO<g�K<w�G<�)D<�b@<%�<<<�8<�5<�`1<��-<��)<A&<ӓ"<��<YF<�<�<)x<!�<?`	<��<�a<%��;e��;
2�;�t�;x��;B,�;v��;�(�;���;�n�;�.�;�;��;q�;���;#%�;�c�;���;�#�;Q��;:=�;&�y;Iao;be;G�Z;�Q;�BG;��=;074;��*;d�!;y�;�;=b;׼�:5��:Ԃ�:�M�:�W�:��:(�:X�:<�}:;`:��B:U�%:�n	::|�97̢9\gW9��8_ݯ��BظI�U��G��8*ӹ�N����"6�cCO��5h����Ќ�����:��V���d���bɺ�Tպ�8���m���gQ��-������v���r�):%�Q�*�$�0�~6��:<���A���G��dM��S���X�Ń^�o8d��i���o��Ru�z{�4]��C7�����숻Aǋ������~���[��
9������  �  �=�%=��=!m=�=��=�V=b� =ڛ => =5��<��<�F�<��<���<��<L�<���<���<��<�E�<+��<]��<���<�0�<�h�<���<��<;	�<<�<fm�<=��<���<#��<#�<3L�<`s�<���<λ�<���<m��<��<X1�<\H�<�\�<�m�<O|�<W��<2��<���<i��<���<���<d��<�q�<�^�<�G�<,�<��<���<���<!��<HZ�<-!�<���<��<�U�<"�<��<(Y�<���<���<*�<���<QE�<�ʿ<�J�<`ż<�:�<���<W�<=~�<z�<>�<\��<B�<=�<܉�<�Ҫ<��<�Y�<��<ӣ<-�<K@�<�r�<���<�Ϛ<��<$�<K�<p�<o��<��<SՍ<�<��<�-�<�H�<6c�<�|�<;��<sZ}<��y<��u<U�q<�n<�?j<�lf<r�b<y�^<G�Z<�&W<�WS<��O<&�K<c�G<|)D<�b@<N�<<Q�8<5<a1<,�-<��)<tA&<�"<�<�F<<�<<Yx<n�<�`	<�<!b<��;���;Y2�;9u�;@��;,�;F��;7(�;���;Ln�;Z.�;��;-�;��;	��;�$�;Zc�;:��;1#�;��;�<�;7�y; ao;�e;Y�Z;�	Q;&CG;g�=;�74;@�*;V�!;��;�;gc;��:��::��:0O�:�Y�:%��:2)�:��:�}:=`:A�B:(�%:�k	:�x�9�Ģ9�\W9���8`��^\ظw�U�
Q��,3ӹS�p��v&6�oGO�u:h�����ь�
���;��sW���c���aɺNTպy7ẙ�.���%P��,�Q��������q�;9%�^�*�ξ0�u}6�:<���A�%�G�]dM�S���X�x�^��8d�x�i�G�o��Su��{��]���7��#���숻�ǋ�>���)��\��9�����  �  �=�%=��="m=�=��=�V=g� =� =*> =T��<��<�F�<��<���<��<+L�<ڋ�<���<��<�E�<8��<|��<���<�0�<�h�<���<
��<,	�<�;�<Gm�<!��<_��<��<�"�<L�<Ds�<v��<���<���<O��<��<K1�<TH�<�\�<�m�<E|�<f��<L��<���<���<���<��<���<�q�<_�<�G�<3,�<��<���<��<B��<WZ�<A!�<���<
��<�U�<�<޲�<Y�<���<Ԕ�<e*�<���<E�<qʿ<iJ�<5ż<�:�<w��<8�<~�<]�<	>�<S��<;�<=�<؉�<�Ҫ<�<�Y�<��<8ӣ<@�<p@�<�r�<���<К<=��<0$�<&K�<<p�<���<;��<_Ս<%�<��<�-�<�H�<-c�<�|�<+��<NZ}<F�y<b�u<�q<5n<p?j<�lf<1�b<$�^<��Z<�&W<bWS<t�O<�K<U�G<h)D<�b@<D�<<Z�8<W5<3a1<j�-<(�)<�A&<V�"<R�<G<��<i<�x<��<�`	<L�<\b<���;��;V2�;<u�;N��;�+�;0��;(�;z��;�m�;�-�;��;��;h�;O��;($�;�b�;���;�"�;���;�<�;��y;�`o;qe;s�Z;{	Q;�CG;C�=;c84;f�*;�!;�;�;�d;���:��:��:Q�:�\�:���:b+�:��:��}:�`:��B:7�%:!k	:ww�9�¢9�SW9 ��8����}ظp�U��X���>ӹ�W�{��B,6��JO�>h������Ҍ�t��!<��jW��d��+bɺ�Rպ�6�����O��+�o�+��w��Sp�8%�e�*���0��|6��8<���A�0�G�dM�FS���X���^��8d���i�ڠo��Tu��{�<^��~8�����y툻Bȋ�棎�����\��:��n���  �  ܁=�%=��=$m=�=��=�V=p� =� =:> =p��<��<�F�<0��<���<��<WL�<��<���<��<F�<G��<���<���<�0�<�h�<w��<���<	�<�;�<,m�<���<A��<���<�"�<�K�<s�<Z��<���<���<-��<y�<;1�<;H�<�\�<�m�<E|�<i��<R��<���<���<ӑ�<:��<���<r�<4_�<H�<Q,�<�<��<+��<^��<fZ�<G!�<���<
��<�U�<$�<Ų�<Y�<���<���<K*�<T��<�D�<Bʿ<<J�<ż<�:�<V��<�<~�<6�<�=�<4��<*�<=�<Ӊ�<�Ҫ<�<�Y�<'��<Vӣ<Y�<�@�<�r�<Ң�<GК<`��<S$�<RK�<Xp�<���<Q��<pՍ<.�<��<�-�<�H�<0c�<r|�<��<Z}<�y<1�u<��q<�n<?j<Glf<ҙb<��^<��Z<\&W<#WS<9�O<�K<�G<b)D<�b@<B�<<o�8<e5<Ua1<��-<i�)<�A&<��"<��<QG<��<�<�x<	�<a	<��<�b<��;B��;�2�;>u�;m��;�+�;Ġ�;�'�;���;{m�;n-�;��;"�;��;���;�#�;Bb�;��;�"�;��;j<�;l�y;`o;�e;��Z;�	Q;�CG;�=;�84;H�*;��!;��;;�e;R��:��:���: T�:�^�:��:6-�:��:��}:+`:Q�B:H�%:}l	:r�9o��9FKW9P��8��ŵ�ظL
V��c���Hӹ�]�����/6��OO�Ah�񄀺�ӌ�7�� =���V��,d���aɺ$Rպ�5������N�n*��F����5o��6%��*�ռ0��{6�L8<��A��G��cM�KS���X���^��9d�W�i���o��Uu�b	{��^���8��[���ȋ�i���R��� ]��|:������  �  ҁ=�%=��=m=�=��=�V=� =�� =I> =���<�<�F�<Q��<��<�<zL�<��<���<	�<F�<f��<���<���<�0�<�h�<o��<���<	�<�;�<m�<М�<$��<���<�"�<�K�<�r�<F��<`��<a��<��<c�<%1�<4H�<�\�<�m�<]|�<|��<h��<֓�<���<���<X��<̀�<%r�<U_�<%H�<t,�<2�<,��<S��<o��<{Z�<a!�<���<"��<�U�<�<���<�X�<���<���<%*�<.��<�D�<ʿ<J�<�ļ<�:�<;��<��<�}�< �<�=�<��<�<�<�<Ӊ�<�Ҫ<�<�Y�<9��<iӣ<��<�@�<s�<���<lК<���<u$�<nK�<}p�<ʓ�<b��<�Ս<:�<��<�-�<�H�< c�<g|�<��<�Y}<߈y<޶u<z�q<�n<�>j<lf<�b<��^<i�Z<&W<�VS<	�O<üK<��G<I)D<�b@<V�<<��8<y5<�a1<��-<��)<<B&<�"<��<�G<A�<�<<y<A�<^a	<��<�b<���;i��;�2�;`u�;#��;�+�;���;�'�;���;2m�;�,�;'�;��;6�;]��;�"�;�a�;���;�!�;ͣ�;<�;��y;�_o;$e;/�Z;P
Q;pDG;<�=;�94;��*;-�!;��;�;�f;s��:��:K��:�U�:>`�:���:^.�:E�:X�}:5`:��B:4�%:9i	:;p�9��9m@W9`|�8�yε�ظ�V��m���Oӹ�a�����26��TO�ZDh�'����Ԍ�j���=��xX��d��`ɺ�Qպ�3�������JM��)�� ������*n��5%�!�*���0��z6��7<�%�A���G�;cM��S�O�X�)�^�(:d���i�l�o�.Vu��
{�L_��R9����c�ɋ�Ф��݀���]���:��=���  �  ā=�%=��=m=�=��=�V=�� =� =T> =���<%�<(G�<{��<��<G�<�L�<3��<��<	�<2F�<i��<���<���<�0�<�h�<y��<���<��<�;�<�l�<Ü�<���<���<z"�<�K�<�r�<��<N��<E��<��<Q�<1�<BH�<�\�<�m�<M|�<��<o��<��<֔�<��<u��<���<Vr�<q_�<=H�<�,�<G�<J��<g��<���<�Z�<d!�<���<��<�U�<�<ʲ�<�X�<u��<���<*�<��<�D�<�ɿ<�I�<�ļ<d:�<��<��<�}�<�<�=�<��<)�<�<�<؉�<�Ҫ<'�<�Y�<M��<�ӣ<��<�@�<>s�<&��<yК<���<�$�<�K�<�p�<ᓑ<���<�Ս<G�<��<�-�<�H�<#c�<s|�<�<�Y}<��y<��u<G�q<on<�>j<�kf<E�b<W�^<,�Z<�%W<�VS<�O<��K<�G<P)D<�b@<L�<<��8<�5<�a1<��-<��)<nB&<�"<F�<�G<X�<T<�y<s�<�a	<��<�b<���;���;�2�;uu�;<��;�+�;���;F'�;��;�l�;�,�;� �;�;��;���;�"�;Fa�;[��;�!�;{��;�;�;F�y;j`o;<e;��Z;�	Q;�DG;~�=;":4;��*;��!;��;�;jh;A��:Q�:u��:eW�:+b�:��:B0�:�:��}:!`:��B:<�%:�i	:Zt�9���9�5W9^g�8�ֵ�ظ�*V�t��_YӹSf�'�� 86��VO�UHh����7֌�����<��XX���c��1aɺ�Pպ�3��8����L��(�������H���l�o4%���*��0��y6��6<���A�"�G�YcM�S���X��^��9d���i�ܢo��Vu�M{��_��:��t���ʋ�w���T����]��1;��v���  �  ��=�%=x�=m=�=ų=�V=�� =� =V> =���<G�<0G�<���<9��<R�<�L�<X��<��<$	�<LF�<g��<���<���<�0�<�h�<X��<���<��<�;�<�l�<���<���<���<p"�<|K�<�r�<���<6��<5��<���<D�<�0�<%H�<u\�<�m�<N|�<���<x��<��<��<��<���<���<]r�<_�<OH�<�,�<^�<k��<f��<���<�Z�<g!�<��<��<�U�<��<���<�X�<f��<l��<�)�<��<�D�<�ɿ<�I�<�ļ<Z:�<骹<��<�}�<�ߴ<�=�<���<�<�<�<މ�<�Ҫ<E�<�Y�<g��<�ӣ<��<�@�<Os�</��<�К<���<�$�<�K�<�p�<ⓑ<���<�Ս<Z�<��<�-�<�H�<c�<]|�<ߔ�<�Y}<x�y<��u<�q<<n<w>j<�kf<1�b<,�^<��Z<�%W<�VS<܈O<i�K<��G<)D<�b@<\�<<��8<�5<�a1<)�-<��)<�B&<V�"<W�<
H<��<m<�y<��<�a	<�<c<���;: �;�2�;�u�;��;p+�;E��;�&�;P��;gl�;o,�; �;��;��;X��;k"�;�`�;��;Q!�;(��;�;�;��y;�_o;�e;��Z;�	Q;�EG;Ѫ=;�:4;��*;��!;��;y;�h;5��:r	�:��:�X�:Ld�:��:�1�:d�:��}:+!`:��B:��%:ag	:Fl�9_��9�.W9�S�8'�ڵ��ظn<V��u���_ӹ�g����<6�gXO��Jh����r׌�	���>��,Y��c���`ɺ�Nպ�3��	�5���vL��'�q��P������l�84%���*�%�0��y6�6<���A���G��bM��S���X���^�x:d�Y�i� �o��Wu��{�`��j:������:ʋ�̥������,^���;������  �  ��=�%=��=m=�=��=�V=�� =� =b> =���<O�<>G�<���<f��<_�<�L�<W��<6��</	�<VF�<r��<���<���<�0�<�h�<j��<���<��<�;�<�l�<���<���<u��<S"�<iK�<�r�<���<%��<.��<���<:�<
1�<.H�<�\�<�m�<L|�<���<o��<���<��<+��<���<��<kr�<�_�<uH�<�,�<r�<f��<���<���<�Z�<e!�<���<��<�U�<�<���<�X�<_��<_��<�)�<��<�D�<�ɿ<�I�<�ļ<>:�<骹<��<�}�<�ߴ<�=�<
��<�<�<�<Љ�<�Ҫ<*�<�Y�<q��<�ӣ<��<�@�<_s�<;��<�К<���<�$�<�K�<�p�<���<���<�Ս<I�<��<�-�<�H�<c�<e|�<攀<�Y}<b�y<y�u<��q<6n<3>j<bkf<�b<�^<��Z<�%W<|VS<��O<v�K<��G<9)D<�b@<K�<<��8<�5<�a1<2�-<�)<�B&<f�"<u�<3H<�<�<�y<��<�a	<)�<2c<���;���;�2�;vu�;>��;�+�;r��;'�;��;Tl�;,�; �;��;'�;��;�!�;�`�;µ�;:!�;���;�;�;�y;�_o;$e;��Z;�	Q;�DG;��=;;4;��*;��!;��;; i;c��:��:Ð�:-Z�:d�:��:�1�:E��:K�}:.`:��B:��%:ki	:-o�9²�9�+W9hG�8ӌ۵\ٸ�9V�i~��eeӹ�k�w��m<6�s[O�|Kh�N���r׌�O���=��NX���c���`ɺbPպ73�	������K��'�������)���k��3%�(�*�ι0� y6��5<�4�A��G��bM�-S���X�e�^�;:d��i���o�#Xu�?{�P`��w:������ʋ��け�y^���;������  �  ��=�%={�=m=�=γ=�V=�� =� =e> =���<S�<XG�<���<O��<\�<�L�<S��<F��<*	�<FF�<���<���<���<�0�<�h�<Z��<���<��<�;�<�l�<���<���<g��<V"�<�K�<�r�<���<��<.��<���<5�<�0�<H�<\�<�m�<h|�<���<���<��<ڔ�<C��<���<��<rr�<�_�<_H�<�,�<��<a��<���<���<�Z�<~!�<���<1��<�U�<��<���<�X�<X��<c��<�)�<��<�D�<�ɿ<�I�<�ļ</:�<�<��<�}�<�ߴ<�=�<�< �<�<�<҉�<�Ҫ<7�<Z�<e��<�ӣ<��<�@�<vs�<9��<�К<���<�$�<�K�<�p�<��<���<�Ս<\�<��<�-�<�H�<c�<I|�<۔�<�Y}<�y<y�u<��q<.n< >j<�kf<�b<�^<��Z<�%W<�VS<��O<e�K<��G< )D<�b@<c�<<��8<�5<�a1<�-<�)<�B&<n�"<��<%H<��<�<�y<��<�a	< �<c<#��;	 �;a3�;�u�;0��;+�;	��;�&�;
��;�l�;�+�;% �;r�;1�;���;�!�;�`�;���;:!�;��;s;�;��y;_o;�e;y�Z;�
Q;uEG;C�=;X;4;��*;��!;��;�;Vi;9��:~
�:��:Q[�:�c�:���:�0�:d��:p�}:�`:��B:��%:�h	:�h�9㭢9�(W9�K�8۵Uٸ07V�B����^ӹ�j�Q���;6��\O�GJh�0����׌����?���X���c���^ɺ�Oպ�1��	�����J��'�2�����֠�l�3%��*�޹0��x6��6<���A�}�G�DbM��S��X���^�;d�w�i�ңo��Wu�>{�i`���:��;��V�ʋ�
�����^���;������  �  ��=�%=��=m=�=��=�V=�� =� =b> =���<O�<>G�<���<f��<_�<�L�<W��<6��</	�<VF�<r��<���<���<�0�<�h�<j��<���<��<�;�<�l�<���<���<u��<S"�<iK�<�r�<���<%��<.��<���<:�<
1�<.H�<�\�<�m�<L|�<���<o��<���<��<+��<���<��<kr�<�_�<uH�<�,�<r�<f��<���<���<�Z�<e!�<���<��<�U�<�<���<�X�<_��<_��<�)�<��<�D�<�ɿ<�I�<�ļ<>:�<骹<��<�}�<�ߴ<�=�<
��<�<�<�<Љ�<�Ҫ<*�<�Y�<q��<�ӣ<��<�@�<_s�<;��<�К<���<�$�<�K�<�p�<���<���<�Ս<I�<��<�-�<�H�<c�<e|�<攀<�Y}<b�y<y�u<��q<6n<3>j<bkf<�b<�^<��Z<�%W<|VS<��O<v�K<��G<9)D<�b@<K�<<��8<�5<�a1<2�-<�)<�B&<f�"<u�<3H<�<�<�y<��<�a	<)�<2c<���;���;�2�;vu�;>��;�+�;r��;'�;��;Tl�;,�; �;��;'�;��;�!�;�`�;µ�;:!�;���;�;�;�y;�_o;$e;��Z;�	Q;�DG;��=;;4;��*;��!;��;; i;c��:��:Ð�:-Z�:d�:��:�1�:E��:K�}:.`:��B:��%:ki	:-o�9²�9�+W9hG�8ӌ۵\ٸ�9V�i~��eeӹ�k�w��m<6�s[O�|Kh�N���r׌�O���=��NX���c���`ɺbPպ73�	������K��'�������)���k��3%�(�*�ι0� y6��5<�4�A��G��bM�-S���X�e�^�;:d��i���o�#Xu�?{�P`��w:������ʋ��け�y^���;������  �  ��=�%=x�=m=�=ų=�V=�� =� =V> =���<G�<0G�<���<9��<R�<�L�<X��<��<$	�<LF�<g��<���<���<�0�<�h�<X��<���<��<�;�<�l�<���<���<���<p"�<|K�<�r�<���<6��<5��<���<D�<�0�<%H�<u\�<�m�<N|�<���<x��<��<��<��<���<���<]r�<_�<OH�<�,�<^�<k��<f��<���<�Z�<g!�<��<��<�U�<��<���<�X�<f��<l��<�)�<��<�D�<�ɿ<�I�<�ļ<Z:�<骹<��<�}�<�ߴ<�=�<���<�<�<�<މ�<�Ҫ<E�<�Y�<g��<�ӣ<��<�@�<Os�</��<�К<���<�$�<�K�<�p�<ⓑ<���<�Ս<Z�<��<�-�<�H�<c�<]|�<ߔ�<�Y}<x�y<��u<�q<<n<w>j<�kf<1�b<,�^<��Z<�%W<�VS<܈O<i�K<��G<)D<�b@<\�<<��8<�5<�a1<)�-<��)<�B&<V�"<W�<
H<��<m<�y<��<�a	<�<c<���;: �;�2�;�u�;��;p+�;E��;�&�;P��;gl�;o,�; �;��;��;X��;j"�;�`�;��;Q!�;(��;�;�;��y;�_o;�e;��Z;�	Q;�EG;Ѫ=;�:4;��*;��!;��;y;�h;5��:r	�:��:�X�:Ld�:��:�1�:d�:��}:+!`:��B:��%:ag	:Fl�9_��9�.W9�S�8'�ڵ��ظn<V��u���_ӹ�g����<6�gXO��Jh����r׌�	���>��,Y��c���`ɺ�Nպ�3��	�5���vL��'�q��P������l�84%���*�%�0��y6�6<���A���G��bM��S���X���^�x:d�Y�i� �o��Wu��{�`��j:������:ʋ�̥������,^���;������  �  ā=�%=��=m=�=��=�V=�� =� =T> =���<%�<(G�<{��<��<G�<�L�<3��<��<	�<2F�<i��<���<���<�0�<�h�<y��<���<��<�;�<�l�<Ü�<���<���<z"�<�K�<�r�<��<N��<E��<��<Q�<1�<BH�<�\�<�m�<M|�<��<o��<��<֔�<��<u��<���<Vr�<q_�<=H�<�,�<G�<J��<g��<���<�Z�<d!�<���<��<�U�<�<ʲ�<�X�<u��<���<*�<��<�D�<�ɿ<�I�<�ļ<d:�<��<��<�}�<�<�=�<��<)�<�<�<؉�<�Ҫ<'�<�Y�<M��<�ӣ<��<�@�<>s�<&��<yК<���<�$�<�K�<�p�<ᓑ<���<�Ս<G�<��<�-�<�H�<#c�<s|�<�<�Y}<��y<��u<G�q<on<�>j<�kf<E�b<W�^<,�Z<�%W<�VS<�O<��K<�G<P)D<�b@<L�<<��8<�5<�a1<��-<��)<nB&<�"<G�<�G<X�<T<�y<s�<�a	<��<�b<���;���;�2�;tu�;<��;�+�;���;F'�;��;�l�;�,�;� �;�;��;���;�"�;Fa�;[��;�!�;{��;�;�;F�y;j`o;<e;��Z;�	Q;�DG;~�=;":4;��*;��!;��;�;jh;A��:Q�:u��:eW�:+b�:��:B0�:�:��}:!`:��B:<�%:�i	:Zt�9���9�5W9^g�8�ֵ�ظ�*V�t��_YӹSf�'�� 86��VO�UHh����7֌�����<��XX���c��1aɺ�Pպ�3��8����L��(�������H���l�o4%���*��0��y6��6<���A�"�G�YcM�S���X��^��9d���i�ܢo��Vu�M{��_��:��t���ʋ�w���T����]��1;��v���  �  ҁ=�%=��=m=�=��=�V=� =�� =I> =���<�<�F�<Q��<��<�<zL�<��<���<	�<F�<f��<���<���<�0�<�h�<o��<���<	�<�;�<m�<М�<$��<���<�"�<�K�<�r�<F��<`��<a��<��<c�<%1�<4H�<�\�<�m�<]|�<|��<h��<֓�<���<���<X��<̀�<%r�<U_�<%H�<t,�<2�<,��<S��<o��<{Z�<a!�<���<"��<�U�<�<���<�X�<���<���<%*�<.��<�D�<ʿ<J�<�ļ<�:�<;��<��<�}�< �<�=�<��<�<�<�<Ӊ�<�Ҫ<�<�Y�<9��<iӣ<��<�@�<s�<���<lК<���<u$�<nK�<}p�<ʓ�<b��<�Ս<:�<��<�-�<�H�< c�<g|�<��<�Y}<߈y<޶u<z�q<�n<�>j<lf<�b<��^<i�Z<&W<�VS<	�O<üK<��G<I)D<�b@<V�<<��8<y5<�a1<��-<��)<<B&<�"<��<�G<A�<�<<y<A�<^a	<��<�b<���;i��;�2�;`u�;#��;�+�;���;�'�;���;2m�;�,�;'�;��;6�;]��;�"�;�a�;���;�!�;ͣ�;<�;��y;�_o;$e;/�Z;P
Q;pDG;<�=;�94;��*;-�!;��;�;�f;s��:��:K��:�U�:>`�:���:^.�:E�:X�}:5`:��B:4�%:9i	:;p�9��9m@W9`|�8�yε�ظ�V��m���Oӹ�a�����26��TO�ZDh�'����Ԍ�j���=��xX��d��`ɺ�Qպ�3�������JM��)�� ������*n��5%�!�*���0��z6��7<�%�A���G�;cM��S�O�X�)�^�(:d���i�l�o�.Vu��
{�L_��R9����c�ɋ�Ф��݀���]���:��=���  �  ܁=�%=��=$m=�=��=�V=p� =� =:> =p��<��<�F�<0��<���<��<WL�<��<���<��<F�<G��<���<���<�0�<�h�<w��<���<	�<�;�<,m�<���<A��<���<�"�<�K�<s�<Z��<���<���<-��<y�<;1�<;H�<�\�<�m�<E|�<i��<R��<���<���<ӑ�<:��<���<r�<4_�<H�<Q,�<�<��<+��<^��<fZ�<G!�<���<
��<�U�<$�<Ų�<Y�<���<���<K*�<T��<�D�<Bʿ<<J�<ż<�:�<V��<�<~�<6�<�=�<4��<*�<=�<Ӊ�<�Ҫ<�<�Y�<'��<Vӣ<Y�<�@�<�r�<Ң�<GК<`��<S$�<RK�<Xp�<���<Q��<pՍ<.�<��<�-�<�H�<0c�<r|�<��<Z}<�y<1�u<��q<�n<?j<Glf<ҙb<��^<��Z<\&W<#WS<9�O<�K<�G<b)D<�b@<B�<<o�8<e5<Ua1<��-<i�)<�A&<��"<��<QG<��<�<�x<	�<a	<��<�b<��;B��;�2�;>u�;m��;�+�;Ġ�;�'�;���;{m�;n-�;��;"�;��;���;�#�;Bb�;��;�"�;��;j<�;l�y;`o;�e;��Z;�	Q;�CG;�=;�84;H�*;��!;��;;�e;R��:��:���: T�:�^�:��:6-�:��:��}:+`:Q�B:H�%:}l	:r�9o��9FKW9P��8��ŵ�ظL
V��c���Hӹ�]�����/6��OO�Ah�񄀺�ӌ�7�� =���V��,d���aɺ$Rպ�5������N�n*��F����5o��6%��*�ռ0��{6�L8<��A��G��cM�KS���X���^��9d�W�i���o��Uu�b	{��^���8��[���ȋ�i���R��� ]��|:������  �  �=�%=��="m=�=��=�V=g� =� =*> =T��<��<�F�<��<���<��<+L�<ڋ�<���<��<�E�<8��<|��<���<�0�<�h�<���<
��<,	�<�;�<Gm�<!��<_��<��<�"�<L�<Ds�<v��<���<���<O��<��<K1�<TH�<�\�<�m�<E|�<f��<L��<���<���<���<��<���<�q�<_�<�G�<3,�<��<���<��<B��<WZ�<A!�<���<
��<�U�<�<޲�<Y�<���<Ԕ�<e*�<���<E�<qʿ<iJ�<5ż<�:�<w��<8�<~�<]�<	>�<S��<;�<=�<؉�<�Ҫ<�<�Y�<��<8ӣ<@�<p@�<�r�<���<К<=��<0$�<&K�<<p�<���<;��<_Ս<%�<��<�-�<�H�<-c�<�|�<+��<NZ}<F�y<b�u<�q<5n<p?j<�lf<1�b<$�^<��Z<�&W<bWS<t�O<�K<U�G<h)D<�b@<D�<<Z�8<W5<3a1<j�-<(�)<�A&<V�"<R�<G<��<i<�x<��<�`	<K�<\b<���;��;V2�;<u�;N��;�+�;0��;(�;y��;�m�;�-�;��;��;h�;O��;($�;�b�;���;�"�;���;�<�;��y;�`o;qe;s�Z;{	Q;�CG;C�=;c84;f�*;�!;�;�;�d;���:��:��:Q�:�\�:���:b+�:��:��}:�`:��B:7�%:!k	:ww�9�¢9�SW9 ��8����}ظp�U��X���>ӹ�W�{��B,6��JO�>h������Ҍ�t��!<��jW��d��+bɺ�Rպ�6�����O��+�o�+��w��Sp�8%�e�*���0��|6��8<���A�0�G�dM�FS���X���^��8d���i�ڠo��Tu��{�<^��~8�����y툻Bȋ�棎�����\��:��n���  �  �=�%=��=!m=�=��=�V=b� =ڛ => =5��<��<�F�<��<���<��<L�<���<���<��<�E�<+��<]��<���<�0�<�h�<���<��<;	�<<�<fm�<=��<���<#��<#�<3L�<`s�<���<λ�<���<m��<��<X1�<\H�<�\�<�m�<O|�<W��<2��<���<i��<���<���<d��<�q�<�^�<�G�<,�<��<���<���<!��<HZ�<-!�<���<��<�U�<"�<��<(Y�<���<���<*�<���<RE�<�ʿ<�J�<`ż<�:�<���<W�<=~�<z�<>�<\��<B�<=�<܉�<�Ҫ<��<�Y�<��<ӣ<-�<K@�<�r�<���<�Ϛ<��<$�<K�<p�<o��<��<SՍ<�<��<�-�<�H�<6c�<�|�<;��<sZ}<��y<��u<U�q<�n<�?j<�lf<r�b<y�^<G�Z<�&W<�WS<��O<&�K<c�G<|)D<�b@<N�<<Q�8<5<a1<,�-<��)<tA&<�"<�<�F<<�<<Yx<n�<�`	<�<!b<��;���;X2�;9u�;@��;,�;F��;7(�;���;Ln�;Z.�;��;-�;��;	��;�$�;Zc�;:��;1#�;��;�<�;7�y; ao;�e;Y�Z;�	Q;&CG;g�=;�74;@�*;V�!;��;�;gc;��:��::��:0O�:�Y�:%��:2)�:��:�}:=`:A�B:(�%:�k	:�x�9�Ģ9�\W9���8`��^\ظw�U�
Q��,3ӹS�p��v&6�oGO�u:h�����ь�
���;��sW���c���aɺNTպy7ẙ�.���%P��,�Q��������q�;9%�^�*�ξ0�u}6�:<���A�%�G�]dM�S���X�x�^��8d�x�i�G�o��Su��{��]���7��#���숻�ǋ�>���)��\��9�����  �  ��=�%=��=&m=}=��=�V=X� =Λ => =��<��<tF�<���<~��<�<�K�<���<u��<��<�E�<��<S��<���<�0�<�h�<���<"��<X	�<<�<�m�<`��<���<F��<4#�<YL�<�s�<Ř�<��<���<���<��<x1�<gH�<�\�<�m�<5|�<N��<��<���<W��<���<ϊ�<O��<�q�<�^�<�G�<�+�<��<���<߼�<��<4Z�<!�<���<���<�U�<?�<���<GY�<���<��<�*�<º�<sE�<�ʿ<�J�<�ż<$;�<ɫ�<{�<e~�<��<:>�<s��<X�<)=�<ω�<�Ҫ<��<�Y�<<ӣ<�<)@�<�r�<a��<�Ϛ<���<�#�<�J�<�o�<[��<��<?Ս<��<x�<�-�<�H�<Lc�<�|�<Z��<�Z}<��y<�u<��q<�n<�?j<Cmf<��b<��^<{�Z<'W<�WS<ȉO<g�K<w�G<�)D<�b@<%�<<<�8<�5<�`1<��-<��)<A&<ӓ"<��<YF<�<�<)x<!�<?`	<��<�a<%��;e��;
2�;�t�;x��;B,�;v��;�(�;���;�n�;�.�;�;��;q�;���;#%�;�c�;���;�#�;Q��;:=�;&�y;Iao;be;G�Z;�Q;�BG;��=;074;��*;d�!;y�;�;=b;׼�:5��:Ԃ�:�M�:�W�:��:(�:X�:<�}:;`:��B:U�%:�n	::|�97̢9\gW9��8`ݯ��BظI�U��G��8*ӹ�N����"6�cCO��5h����Ќ�����:��V���d���bɺ�Tպ�8���m���gQ��-������v���r�):%�Q�*�$�0�~6��:<���A���G��dM��S���X�Ń^�o8d��i���o��Ru�z{�4]��C7�����숻Aǋ������~���[��
9������  �  ��=�%=��=$m=�=��=�V=K� =Ǜ => =���<l�<KF�<���<X��<c�<�K�<}��<_��<�<�E�<���<a��<���<�0�<�h�<���<-��<a	�<><�<�m�<|��<���<u��<X#�<hL�<�s�<��<��<���<���<��<y1�<rH�<�\�<�m�<8|�<\��<��<v��<G��<e��<Ê�<$��<xq�<�^�<nG�<�+�<��<���<���<���<Z�<!�<���<��<�U�</�< ��<MY�<���<*��<�*�<��<�E�<�ʿ<�J�<�ż<W;�<߫�<��<}~�<��<G>�<~��<\�<=�<ቬ<�Ҫ< �<�Y�<���<�ң<�
�<@�<vr�<G��<�Ϛ<���<�#�<�J�<�o�<<��<���<(Ս<��<�<�-�<�H�<=c�<�|�<^��<�Z}<�y<�u<��q<"n<O@j<Wmf<�b<�^<��Z<O'W<XS<��O<p�K<��G<�)D<�b@<3�<<G�8<
5<�`1<�-<��)<�@&<��"<}�<F<��<v<�w<��<`	<��<�a<���;���;2�;u�;B��;1,�;���;�(�;{��;o�;B/�;O�;c�;��;���;�%�;=d�;���;$�;���;�=�;!�y;�ao;�e;��Z;�Q;8CG;��=;�64;�*;^�!;�;�
;;a;���:���:��:K�:�V�:��:�&�:��:�}:,`:J�B:G�%:�l	:I~�9͢9�nW9���8E����$ظ��U�A;���$ӹ�J���e 6��?O�&3h�~��nό�D���:��W���c���bɺ�Sպ:�������7R�q.�l��������s�d;%�l�*���0�6�$;<�O�A���G�]dM��S���X�9�^��7d�c�i��o�Ru��{��\���6������눻�Ƌ�
���u~��%[���8��`���  �  ��=�%=��=)m=~=��=�V=B� =Û =�= =��<P�<9F�<���<7��<^�<�K�<d��<O��<d�<�E�<��<H��<���<�0�<�h�<���<=��<i	�<T<�<�m�<���<���<|��<e#�<L�<�s�<���<*��<���<���<��<w1�<�H�<�\�<n�<)|�<;��<��<d��<6��<R��<���< ��<rq�<�^�<YG�<�+�<h�<���<���<��<Z�<� �<���<��<�U�<4�<"��<PY�<��<@��<�*�<
��<�E�<�ʿ<�J�<�ż<a;�<���<��<~~�<��<V>�<���<{�<=�<艬<�Ҫ<��<�Y�<՗�<�ң<�
�< @�<Xr�<A��<�Ϛ<���<�#�<�J�<�o�<#��<鴏<Ս<��<^�<�-�<I�<Kc�<�|�<^��<�Z}<��y<:�u< �q<9n<i@j<�mf<)�b<(�^<��Z<y'W<XS<0�O<y�K<��G<�)D<�b@<*�<<	�8<�5<�`1<ϧ-<S�)<�@&<X�"<V�<F<v�<i<�w<��<�_	<n�<�a<e��;,��;�1�;u�;E��;�,�;ԡ�;�(�;���;o�;�/�;��;z�;$�;"��;�%�;�d�;���;0$�;���;�=�;�y;�bo;�e;��Z;lQ;#BG;̦=;�54;��*;��!;~�;]	;a;���:w��:���:�H�:LU�:؞�:�%�:�:F�}:`:.�B:��%:3m	:]��9q͢9zW9w�8!����׸m�U��9�� ӹCI����6�X<O�M3h��|���Ό�|���8���V���c��Vdɺ�Uպ_;Ặ�J����R�4/�`�������;t��;%�i +��0��6��;<���A�<�G�beM��S�`�X�ʃ^��6d�b�i��o��Qu�E{�I\��{6�����{눻[Ƌ�衎��}���Z���8������  �  �=�%=��=$m=�=��=�V=E� =�� =�= =ֿ�<I�<-F�<s��<$��<;�<�K�<V��<C��<Y�<�E�<��<P��<���<�0�<�h�<���</��<y	�<S<�<�m�<���<���<���<�#�<�L�<�s�<��<%��<��<���<��<1�<zH�<�\�<�m�<8|�<J��<��<b��<$��<N��<���<��<Uq�<q^�<?G�<�+�<n�<s��<���<ߍ�<Z�<	!�<���<��<�U�<6�<��<RY�<��<@��<�*�<��<�E�<˿<K�<�ż<p;�<��<��<�~�<��<f>�<���<i�<=�<މ�<�Ҫ<��<�Y�<ʗ�<�ң<�
�<�?�<[r�<��<�Ϛ<���<�#�<�J�<�o�<��<Դ�<Ս<��<q�<�-�<�H�<Fc�<�|�<j��<[}<�y<f�u<�q<Xn<�@j<�mf<N�b<E�^<��Z<�'W<@XS<<�O<��K<��G<�)D<�b@<3�<<.�8<�5<�`1<��-<C�)<�@&<H�"<?�<�E<N�<"<�w<��<�_	<V�<�a<~��;G��;�1�;�t�;,��;S,�;���;)�;���;o�;�/�;��;��;��;���;$&�;�d�;|��;�$�;���;>�;B�y;�ao;�e;C�Z;�Q;�BG;)�=;�54;��*;��!;��;v	;`;���:���:�~�:)I�:T�:���:�$�:��:�}:�`:*�B:��%:Bm	:<��9�͢9��W9��8�����ظ��U�V6��ӹ,E�N��t6��;O�~/h��|���͌�3���9��W��<d��KcɺUպ�:�t����S��/�N���8��$u�_<%�� +���0� �6�.<<���A���G��dM��S���X��^��7d���i�ϝo�\Qu��{�E\��>6��}���ꈻƋ������}���Z��P8������  �  �={#=��=�i=�=��=!R=t� =|� =G8 =���<(��<8�<ky�<'��<(��<�9�<x�<ҵ�<���<�.�<�i�<��<���<��<|K�<��<��<���<(�<I�<dw�<'��<+��<[��<��<=E�<�h�<��<��<���<��<���<��<�<Z.�<�:�<�C�<�I�<&L�<K�<IF�<�=�<z1�<!�<t�<���<v��<���<Q��<=c�<H3�<k��<c��<<��<�@�<B��<U��<�S�<H��<��<�6�<���<y]�<��<Do�<X�<[l�<c�<�U�<�·<[+�<N��<��<J�<��<��<�B�<5��<�ը<��<�Z�<��<�ҡ<U
�<Z?�<�q�<���<\Ϙ<���<�$�<L�<r�<E��<��<Fڋ<T��<*�<�6�<�S�<�o�<Ί�<�J}<�~y<�u<��q<�n<�Hj<�zf<h�b<��^<�[<mHW<�}S<��O<:�K<0'H<<cD<4�@<��<<�$9<pj5<r�1<��-<LO*<Ϣ&<��"<�V<O�< <ć<0�<#n<5�	<�l<��<�
�;�8�;au�;J��;4�;���;��;ؕ�;�6�;X��;�;^��;�y�;�{�;D��;���;��;pX�;�Ŏ;H�;^��;�};��r;Yh;#7^;�@T;tJ;`�@;{X7;=.;E�$;5�;�;sK
;|�;ϖ�:���:,��:c��:}��:%�:�Ē:*��:JIi:E�K:�.:��:f��9I��9hv9�9k��7�Р�( ;��Y����ƹ����R
�C�0�	�I�c��|�t���˖����D��?i���}Ǻ�Ӻ'ߺ�k��M�����w�X�v4�������$� {*��D0��
6���;���A�PG��M�z�R���X��@^�o�c�ߴi�oo�.(u�x�z��M��D*�����刻�Ë�㡎�p���_a��=B��9$���  �  �=z#=��=�i=�=��=+R=o� =|� =K8 =���<,��<8�<{y�<-��<9��<�9�<x�<��<���<�.�<�i�<���<���<��<wK�<��<��<���<;�<I�<cw�<��<��<`��<��<5E�<�h�<��<��<���<��<���<��<�<d.�<�:�<�C�<�I�<L�<K�<YF�<�=�<s1�<
!�<��<���<y��<���<j��<Pc�<U3�<b��<p��<Q��<�@�<K��<N��<�S�<@��<&��<�6�<���<}]�<���<=o�<a�<_l�<W�<mU�<�·<V+�<[��<��<J�<��<��<�B�<-��<�ը<��<�Z�<(��<�ҡ<f
�<Y?�<�q�<���<oϘ<���<�$�<,L�<r�<H��< ��<[ڋ<Y��<%�<�6�<�S�<�o�<Ǌ�<�J}<�~y<ڱu<m�q<�n<�Hj<{f<j�b<D�^<�[<]HW<�}S<ݴO<-�K<-'H<'cD<7�@<��<<�$9<�j5<^�1<��-<ZO*<��&<��"<�V<p�<<�<,�<?n<`�	<�l<��<�
�;�8�;Fu�;M��;"�;���;��;ݕ�;�6�;Q��;鰽;��;Sy�;|�;t��;���;>�;rX�;eŎ;H�;���;�};{�r;�Xh;v7^;�@T;�tJ;��@;;X7;�.;��$;�;q;WK
;�;���:���:���:���:���:�%�:^Ē:���:�Ki:��K:>�.:��:F��9���9v9�9Y��7�̠�t;��[��Q�ƹ�������0���I��c�|� t���˖����E��i��T~ǺN�Ӻ�~ߺIl�8M��f��Bw�X��3������$�={*�5D0��
6�}�;��A�lOG��M���R�W�X�7A^�w�c��i�~no�5(u���z��M���*����|刻�Ë�f��������a��FB���#���  �  �=~#=��=�i=�=��=)R=o� =�� =L8 =���<5��<#8�<�y�<.��<I��<�9�<#x�<��<���<�.�<�i�<���<���<��<|K�<��<��<���<.�< I�<fw�<��<��<R��<��<3E�<�h�<���<���<���<��<���<��<
�<q.�<�:�<�C�<�I�<!L�<!K�<TF�<�=�<v1�<!�<��<���<���<´�<s��<Kc�<h3�<i��<m��<J��<�@�<X��<M��<�S�<9��<��<�6�<���<�]�<���<;o�<I�<Kl�<W�<lU�<�·<C+�<O��<��<J�<��<��<C�< ��<�ը<��<�Z�<7��<�ҡ<k
�<X?�<�q�<���<|Ϙ<���<�$�<6L�<r�<^��< ��<Zڋ<P��<*�<�6�<�S�<�o�<���<�J}<�~y<ӱu<��q<�n<�Hj<�zf<Y�b<>�^<�[<[HW<�}S<ŴO<
�K<:'H<cD<K�@<��<<�$9<�j5<^�1<��-<bO*<
�&<��"<�V<��<<	�<,�<On<d�	<�l<��<�
�;�8�;(u�;���;9�;���;��;���;�6�;��;���;%��;Vy�;�{�;��;���;*�;�X�;7Ŏ;�G�;k��;0};��r;�Xh;�7^;�@T;ZtJ;��@;UX7;(.;��$;d�;�;�K
;8�;��:� �:;��:���:`��:	'�:�Ē:ܚ�:/Ki::�K:�.:��:g��9��9�v9j9KC�7t���;��[���ƹ[������0���I��c�}|�#u���˖�����D���g��Ǻ��Ӻ�~ߺlk�@L��x��w� X�w3������ݮ$�{*��C0��
6���;��A�wOG��M�z�R���X�jA^�P�c���i��no��(u���z��M���*��'���刻�Ë�q���j����a���B��"$���  �  �=u#=��=�i=�=��=*R=w� =�� =S8 =���<N��<<8�<�y�<B��<Q��<�9�<<x�<���<���<�.�<�i�<���<���<��<qK�<ހ�< ��<���< �<�H�<Iw�<���<��<F��<��<E�<�h�<Ӊ�<��<���<���<���<��<�<_.�<�:�<�C�<�I�<-L�< K�<gF�<�=�<�1�<+!�<��<���<���<ߴ�<���<^c�<h3�<u��<u��<R��<�@�<D��<E��<�S�<4��<��<�6�<���<^]�<���<"o�<;�<?l�<=�<RU�<�·<;+�<A��<��<J�<��<��<�B�<8��<�ը<��<�Z�<=��<�ҡ<�
�<t?�<�q�<ϡ�<�Ϙ<��<�$�<AL�<r�<[��<��<\ڋ<`��<3�<�6�<�S�<�o�<���<uJ}<�~y<��u<@�q<�n<�Hj<�zf<:�b<�^<�[</HW<�}S<��O<�K<'H<cD<0�@<��<<�$9<�j5<�1<��-<~O*<"�&<��"<�V<��<:<�<g�<�n<��	<�l<��<�;�8�;�u�;f��;�;[��;��;���;x6�;���;���;���;�x�;�{�;蒥;J��;� �;X�;Ŏ;�G�;8��;7};%�r;�Xh;W7^;(AT;�tJ;�@;�X7;!.;B�$;��;�;mL
;��;ݘ�:��:��:���:���:'�:�Œ:k��:bLi:�K:��.:��:���9���9d	v9`9o#�7v頸&;��a��X�ƹ�����&�0��I��c�|�cu��|̖�����E���h��~}Ǻ��Ӻ5~ߺ�j��K����Wv�=W�!3��c���$�%z*��C0�
6���;���A�eOG�qM�6�R�~�X��A^���c���i�boo��(u�~�z�4N��3+��k��戻ċ����������a���B��g$���  �  �=l#=��=�i=�=��=.R=�� =�� =a8 =г�<T��<K8�<�y�<g��<e��<�9�<Bx�<��<���<�.�<j�<���<���<��<�K�<��<���<���<�<�H�<8w�<��<���<)��<��<�D�<}h�<�<��<���<���<���<��<�<[.�<�:�<�C�<�I�<AL�<)K�<�F�<�=�<�1�<8!�<��<���<���<��<���<|c�<p3�<���<���<N��<�@�<;��<Z��<�S�<.��<���<r6�<���<L]�<���<�n�<#�<"l�<�<HU�<�·<0+�<'��<��<�I�< ��<��<�B�<;��<�ը<��<�Z�<J��<�ҡ<�
�<�?�<�q�<���<�Ϙ<"��<�$�<PL�<=r�<b��<(��<fڋ<`��<$�<�6�<�S�<xo�<���<MJ}<`~y<��u<�q<Yn<bHj<�zf<��b<��^<�[<HW<�}S<x�O<�K<�&H<1cD<=�@<��<<�$9<�j5<��1<��-<�O*<E�&<��"<W<ط<�<E�<��<�n<��	<m<��<��;�8�;�u�;.��;[�;~��;��;���;!6�;���;L��;���;�x�;6{�;���;ʾ�;� �;�W�;�Ď;�G�;��;"};��r;bYh;>7^;AT;�tJ;��@;dY7;q.;X�$;%�;�;�L
;��;B��:��:���:���:�ñ:�'�:�ƒ:m��:Li:)�K:��.:��:Z��9���9�v9�
9 �7����;�;j����ƹ������%�0��I��c�|��u���̖����ED���i��:}Ǻ��Ӻ�|ߺIj��J��)��v��V��2��	�|����$�z*�C0�	6���;�ݎA�OG�pM���R�m�X��@^�b�c���i�po�P)u���z�{N���+�����Q戻�ċ����:���b���B���$���  �  �=k#=��=�i=�=��=4R=�� =�� =g8 =��<z��<i8�<�y�<s��<���<�9�<dx�< ��<��<�.�<j�<	��<��<��<xK�<р�<��<���<��<�H�<w�<գ�<���<
��<q�<�D�<\h�<���<Ũ�<���<���<���<��<
�<b.�<�:�<�C�<�I�<IL�<@K�<�F�<>�<�1�<Z!�<��<���<���<��<���<�c�<�3�<���<���<X��<�@�<E��<J��<�S�<��<��<a6�<t��<;]�<���<�n�<��<�k�<�<&U�<p·<+�<��<��<�I�<<��<�B�<A��<�ը<��<�Z�<\��<�ҡ<�
�<�?�<r�<���<�Ϙ<A��<�$�<oL�<Fr�<{��<+��<pڋ<o��<4�<�6�<�S�<to�<���<3J}<6~y<X�u<�q<*n<7Hj<Szf<Ǭb<��^<e[<�GW<�}S<b�O<��K<�&H<cD<5�@<��<<�$9<�j5<��1<��-<�O*<��&<A�"<KW<�<�<��<��<�n<��	</m<�<��;-9�;�u�;���;=�;4��;|�;=��;�5�;~��;;-��;Rx�;�z�;��;���;I �;�W�;yĎ;EG�;�߃;�};��r;�Xh;�7^;XAT; uJ;��@;�Y7;4	.;��$;<�;�;�M
;D�;;��:�:��:A��:&ı:)�:&ǒ:ݜ�:�Mi:��K:4�.:��:���9���9��u9�9��79��M1;��n���ƹ�����
�0���I�,c��|��v��g͖�����D���h���|Ǻ؃Ӻk|ߺVi��I�����u��U��1�z	������$��x*�B0��6���;���A��NG��M�*�R�j�X��A^���c�:�i�hpo��)u���z��N���+��D	���戻�ċ�n��������b��&C���$���  �  �=k#=��=�i=�=��==R=�� =�� =t8 = ��<���<�8�<�y�<���<���<�9�<�x�<4��< ��</�<j�<��<��<��<lK�<΀�<��<���<��<�H�<w�<���<���<���<V�<�D�<5h�<���<���<��<���<���<��<��<`.�<�:�<�C�<�I�<SL�<`K�<�F�<7>�<�1�<y!�<��<��<���<��<ǎ�<�c�<�3�<���<���<g��<�@�<B��<9��<�S�<
��<Ԛ�<S6�<X��<"]�<���<�n�<��<�k�<��<�T�<Z·<�*�<��<��<�I�<�<��<�B�<:��<�ը<�<�Z�<x��<ӡ<�
�<�?�<4r�<!��<�Ϙ<]��<�$�<�L�<]r�<���<4��<�ڋ<n��</�<�6�<�S�<wo�<���<J}<~y<&�u<��q<�n<Hj<zf<��b<p�^< [<�GW<Y}S<L�O<��K<�&H<�bD<)�@<��<<�$9<�j5<ȳ1<. .<P*<��&<g�"<}W<\�<�<ۈ<��<o<	�	<hm<:�<��;�9�;�u�;y��;�;4��;e�;ޔ�;�5�;&��;���;���;�w�;xz�;���;Q��;���;OW�;Ď;G�;�߃; };ۤr;�Xh;{7^;6AT;nuJ;;�@;Z7;>
.;E�$;
�;|;�N
;>�;H��:>�:��:��:�ű:+�:Ȓ:���:Oi:m�K:��.:�:	��9��9�u9��9!�7���D;��r����ƹ������0�r�I�r c�v|��x��HΖ�����E���h��
}Ǻ��Ӻ�{ߺh��G����t�@U�d0�g����ī$�Mx*�wA0�6���;�}�A�<NG�
M�Y�R���X��A^�g�c���i��po�*u���z�,O���,���	��t爻4ŋ����
����b��rC��%���  �  �=c#=��=�i=�=��==R=�� =�� =~8 =��<���<�8�<�y�<���<���<:�<�x�<M��</��<!/�<)j�<��<��<��<rK�<π�<ش�<���<��<�H�<�v�<���<���<���<3�<�D�<%h�<~��<���<_��<���<���<��<��<d.�<�:�<�C�<�I�<mL�<gK�<�F�<K>�<�1�<�!�<�<2��<���<>��<ێ�<�c�<�3�<���<���<a��<A�<B��<;��<�S�<���<Ú�<16�<@��<]�<u��<�n�<��<�k�<��<�T�<?·<�*�<쎴<��<�I�<堯<��<�B�<G��<�ը<�<�Z�<���<ӡ<�
�<�?�<Dr�<=��<�Ϙ<~��<%�<�L�<ur�<���<O��<�ڋ<q��<9�<�6�<�S�<fo�<���<�I}<�}y<��u<��q<�n<�Gj<�yf<b�b<A�^<�[<�GW<#}S<�O<��K<�&H<�bD<3�@<��<<�$9<�j5<��1<B .<-P*<У&<��"<�W<~�< <��<G�<Xo<>�	<�m<W�<$�;v9�;v�;���;9�;?��;,�;Ô�;w5�;���;a��;m��;rw�;�y�;4��;½�;}��;�V�;�Î;�F�;B߃;�};7�r;�Xh;�7^;�AT;puJ;��@;�Z7;{
.;'�$;��;�;�O
;�;���:Y�:V��:o��:.Ǳ:�+�:�ɒ:���:Oi:S�K:E�.:{�:P��9���9��u9��9���7�<��8K;�\{���ƹ׿������0�j�I�U#c��|�7y��1ϖ�����E���h��|Ǻ�Ӻ�zߺg�!G��?��?s��S��/�������$�8w*��@0�Y6���;���A�NG��M��R�a�X��A^���c�@�i��qo�O+u�5�z��O���,��
���爻�ŋ�b���]���-c���C��z%���  �  �=\#=��=�i=�=��=?R=�� =�� =�8 =/��<���<�8�<z�<ٺ�<���<&:�<�x�<i��<D��<./�<>j�<��<$��<��<cK�<���<д�<���<��<�H�<�v�<|��<x��<���<(�<�D�<h�<[��<���<L��<���<���<��<��<R.�<�:�<�C�<�I�<�L�<tK�<�F�<`>�<2�<�!�<"�<R��<��<`��<��<�c�<�3�<���<���<i��<A�<3��<4��<�S�<���<���<6�<4��<�\�<P��<�n�<��<�k�<��<�T�<·<�*�<Ҏ�<�<�I�<Ԡ�<��<�B�<W��<�ը<$�<�Z�<���<8ӡ<�
�<�?�<Tr�<`��<И<���<%�<�L�<�r�<���<e��<�ڋ<���<B�<�6�<�S�<Yo�<���<�I}<�}y<Ӱu<G�q<xn<�Gj<�yf<!�b<�^<�[<JGW<}S<�O<��K<�&H<�bD<�@<��<<%9<�j5<*�1<W .<[P*<	�&<��"<�W<��<s<&�<}�<oo<y�	<�m<u�<|�;�9�;^v�;���;�;	��;�;���;5�;���;뮽;㈷;�v�;�y�;��;=��;���;XV�;�Î;YF�;߃;�};��r;�Xh;&7^; BT;�uJ;�@;�[7;�
.;�$;e�;�;BP
;�;	��:�	�:���:���:ɱ:�,�:�ʒ:���:.Pi:�K:��.:��:���9P��9m�u9�9 ��7B`��];�����i�ƹI���% �B�0���I�$c�~"|��y���ϖ����5F��,i��{Ǻ��Ӻjyߺf��E��U���r� S�S/�j�+���$�dv*�@0��6�d�;���A��MG�AM���R��X�B^�^�c�U�i�&ro��+u���z�"P��H-���
�� 舻>Ƌ�Ԥ��񃑻�c��D���%���  �  �=Y#=��=�i=�=��=GR=�� =�� =�8 =A��<���<�8�<6z�<��<���<9:�<�x�<x��<V��<A/�<?j�<-��<��<��<pK�<���<Ĵ�<q��<��<�H�<�v�<x��<l��<���<�<�D�<�g�<T��<o��<@��<���<l��<��<��<_.�<�:�<�C�<�I�<�L�<�K�<�F�<o>�<2�<�!�<;�<i��<-��<f��<���<�c�<�3�<���<���<m��<�@�<;��<0��<�S�<���<���<6�<��<�\�<A��<zn�<��<�k�<��<�T�<·<�*�<ǎ�<g�<�I�<ՠ�<��<�B�<=��<�ը<%�<�Z�<���<Eӡ<�
�<@�<tr�<r��<(И<���<'%�<�L�<�r�<�<f��<�ڋ<}��<3�<�6�<�S�<Uo�<f��<�I}<�}y<��u<;�q<Un<_Gj<tyf<�b<��^<�[<&GW<�|S<ܳO<d�K<�&H<�bD<2�@<��<<�$9<k5<,�1<� .<sP*<.�&<��"<$X<��<�<j�<��<�o<��	<�m<��<��;�9�;v�;���;?�;��;��;d��;5�;;��;���;ڈ�;�v�;>y�;y��;��;���;?V�;<Î;1F�;�ރ;};�r;jXh;�7^;AT;�uJ;P�@;�[7;�.;V�$;��;�;KQ
;�;���:��:���:���:�ɱ:�-�:D˒:ݟ�:�Pi:=�K:Ġ.:��:Z��9∲9+�u9��9=,�7>g��:c;�,����ƹ�����!���0� J�k(c��#|�{��tЖ�����E��i���|Ǻ��ӺDyߺ'e뺿D����]r��R�P.���@��_�$�v*��?0�M6���;��A��MG��M�9�R��X�-B^���c�'�i�_ro��,u���z�:P���-���
���舻�Ƌ��������c��wD���%���  �  �=X#=��=�i=�=��=PR=�� =�� =�8 =Y��<���<�8�<Dz�<���<��<I:�<�x�<���<Y��<Q/�<<j�<>��<��<��<eK�<���<���<c��<��<pH�<�v�<Y��<Q��<���<��<wD�<�g�<>��<\��<;��<���<a��<��<��<p.�<�:�<D�<J�<�L�<�K�<�F�<�>�<22�<�!�<F�<t��<D��<y��<%��<�c�<�3�<���<���<��<�@�<M��<��<�S�<���<���<6�< ��<�\�<#��<in�<t�<}k�<{�<�T�< ·<�*�<Ȏ�<Y�<�I�<Ƞ�<��<�B�<B��< ֨<#�<[�<���<Pӡ<(�<@�<�r�<���<5И<���<D%�<�L�<�r�<і�<g��<�ڋ<���<?�<�6�<uS�<Vo�<X��<�I}<}}y<��u<	�q<n<NGj<Myf<ܫb<��^<j[<GW<�|S<ڳO<@�K<�&H<�bD<1�@<��<<%9<,k5<(�1<� .<{P*<^�&<>�"<NX<�<�<��<��<�o<��	<�m<��<��;&:�;v�;���;�;��;��;2��;5�;��;���;e��;fv�;y�;0��;߼�;^��;�U�;�; F�;�ރ;�};��r;�Wh;8^;�AT;�vJ;��@;�[7;.;��$;�;�;R
;I�;H��:"�:7��:?��: ʱ:�.�:�˒:E��:MSi:I�K:�.:��:e��9���9��u9��9O��7�x��yq;�#���2�ƹz����$��0��J��*c�X#|��{���Ж�]���F���g��%|Ǻv�ӺQyߺ=d뺌D������p�R��-�b������$�u*��>0�'6�9�;��A�MG�7M���R�>�X��B^�u�c���i�vro��,u���z��P���-�����舻�Ƌ�~���n���d���D���%���  �  �=Y#=��=�i=�=��=MR=�� =Ŗ =�8 =Y��<���<�8�<Nz�<��<��<M:�<�x�<���<h��<^/�<Oj�<9��<��<��<bK�<���<´�<b��<��<qH�<�v�<T��<H��<���<��<hD�<�g�<8��<_��<*��<���<d��<��<��<_.�<�:�<D�<J�<�L�<�K�<�F�<�>�<42�<�!�<Z�<���<C��<}��<��<�c�<�3�<���<���<{��<�@�<=��<"��<�S�<���<���<�5�<��<�\�<��<[n�<o�<qk�<q�<�T�<���<�*�<���<W�<�I�<Π�<��<�B�<E��<�ը<2�<[�<���<Yӡ<�<@�<�r�<���<@И<���<=%�<�L�<�r�<ݖ�<{��<�ڋ<���<9�<�6�<|S�<Xo�<X��<�I}<i}y<��u<��q<n<,Gj<Hyf<��b<��^<W[<GW<�|S<��O<A�K<�&H<�bD<�@<��<<%9< k5<M�1<� .<�P*<^�&<%�"<UX<'�<�<��<��<�o<��	<n<��<��;:�;7v�;���;�;��;��;3��;�4�;
��;m��;S��;Fv�;�x�;.��;���;a��;�U�;Î;�E�;�ރ;�};#�r;Xh;�7^;�AT;lvJ;��@;r\7;h.;!�$;��;�;R
;��;���:�:���:d��:˱:W/�:�̒:q��:�Ri:5�K:J�.:�:��9<��9��u9[�9���7t����r;�k���<�ƹ,���"&�k�0��J�5*c��%|��{���Ж�����F���h���{Ǻ݀Ӻ_xߺc뺚C��<���q��Q��-���y����$�Ou*��>0��6���;�H�A�.MG�.M��R���X��B^�f�c���i� so�'-u�	�z��P���-��S��鈻�Ƌ���������(d���D��<&���  �  �=P#=��=�i=�=��=MR=�� =�� =�8 =_��<���<9�<Kz�<��<��<u:�<�x�<���<i��<L/�<Vj�<;��<��<��<hK�<���<���<m��<��<fH�<�v�<Z��<L��<w��<��<YD�<�g�<%��<K��<��<���<[��<�<��<[.�<�:�<D�<	J�<�L�<�K�<G�<�>�<L2�<�!�<U�<���<J��<���<��<�c�<�3�<���<���<���<A�<4��<(��<�S�<���<���<�5�<���<�\�< ��<Sn�<c�<ak�<v�<�T�<���<�*�<���<_�<�I�<���<��<�B�<K��<�ը<7�<[�<���<gӡ<�<@@�<�r�<���<;И<���<O%�<�L�<�r�<ʖ�<{��<�ڋ<���<<�<�6�<�S�<Co�<\��<�I}<[}y<`�u<��q<n<Gj<>yf<��b<��^<H[<�FW<�|S<��O<T�K<|&H<�bD< �@<��<<%%9< k5<T�1<� .<�P*<k�&<C�"<�X<#�<�<��<#�<�o<��	<
n<��<��;:�;Vv�;���;)�;��;��;_��;�4�;���;	��;m��;Yv�;�x�;��;k��;a��;�U�;�;�E�;�ރ;�};Y�r;JXh;}7^;BT;�vJ;��@;r\7;.;T�$;��;};RR
;��;:��:��:b��:��:�˱:/�:s̒:ޠ�:�Si:'�K:7�.:��:@��9I��9��u9��9���7Ϙ��Ur;�J����ƹ*���v%�x�0�-J�,c��&|�V{���і����7F��Ji���{ǺӀӺ�wߺud�tC��ȋ��q��P�K-������$��t*��>0��6�q�;�G�A�6MG��M���R���X�tB^��c�v�i��ro�`-u���z��P���-�����鈻<ǋ���������zd���D��0&���  �  �=Y#=��=�i=�=��=MR=�� =Ŗ =�8 =Y��<���<�8�<Nz�<��<��<M:�<�x�<���<h��<^/�<Oj�<9��<��<��<bK�<���<´�<b��<��<qH�<�v�<T��<H��<���<��<hD�<�g�<8��<_��<*��<���<d��<��<��<_.�<�:�<D�<J�<�L�<�K�<�F�<�>�<42�<�!�<Z�<���<C��<}��<��<�c�<�3�<���<���<{��<�@�<=��<"��<�S�<���<���<�5�<��<�\�<��<[n�<o�<qk�<q�<�T�<���<�*�<���<W�<�I�<Π�<��<�B�<E��<�ը<2�<[�<���<Yӡ<�<@�<�r�<���<@И<���<=%�<�L�<�r�<ݖ�<{��<�ڋ<���<9�<�6�<|S�<Xo�<X��<�I}<i}y<��u<��q<n<,Gj<Hyf<��b<��^<W[<GW<�|S<��O<A�K<�&H<�bD<�@<��<<%9< k5<M�1<� .<�P*<^�&<%�"<UX<'�<�<��<��<�o<��	<n<��<��;:�;7v�;���;�;��;��;3��;�4�;
��;m��;S��;Fv�;�x�;.��;���;a��;�U�;Î;�E�;�ރ;�};#�r;Xh;�7^;�AT;lvJ;��@;r\7;h.;!�$;��;�;R
;��;���:�:���:d��:˱:W/�:�̒:q��:�Ri:5�K:J�.:�:��9<��9��u9[�9���7t����r;�k���<�ƹ,���"&�k�0��J�5*c��%|��{���Ж�����F���h���{Ǻ݀Ӻ_xߺc뺚C��<���q��Q��-���y����$�Ou*��>0��6���;�H�A�.MG�.M��R���X��B^�f�c���i� so�'-u�	�z��P���-��S��鈻�Ƌ���������(d���D��<&���  �  �=X#=��=�i=�=��=PR=�� =�� =�8 =Y��<���<�8�<Dz�<���<��<I:�<�x�<���<Y��<Q/�<<j�<>��<��<��<eK�<���<���<c��<��<pH�<�v�<Y��<Q��<���<��<wD�<�g�<>��<\��<;��<���<a��<��<��<p.�<�:�<D�<J�<�L�<�K�<�F�<�>�<22�<�!�<F�<t��<D��<y��<%��<�c�<�3�<���<���<��<�@�<M��<��<�S�<���<���<6�< ��<�\�<#��<in�<t�<}k�<{�<�T�< ·<�*�<Ȏ�<Y�<�I�<Ƞ�<��<�B�<B��< ֨<#�<[�<���<Pӡ<(�<@�<�r�<���<5И<���<D%�<�L�<�r�<і�<g��<�ڋ<���<?�<�6�<uS�<Vo�<X��<�I}<}}y<��u<	�q<n<NGj<Myf<ܫb<��^<j[<GW<�|S<ڳO<@�K<�&H<�bD<1�@<��<<%9<,k5<(�1<� .<{P*<^�&<>�"<NX<�<�<��<��<�o<��	<�m<��<��;&:�;v�;���;�;��;��;2��;5�;��;���;e��;fv�;y�;0��;߼�;^��;�U�;�; F�;�ރ;�};��r;�Wh;8^;�AT;�vJ;��@;�[7;.;��$;�;�;R
;I�;H��:"�:7��:?��: ʱ:�.�:�˒:E��:MSi:I�K:�.:��:e��9���9��u9��9O��7�x��yq;�#���2�ƹz����$��0��J��*c�X#|��{���Ж�]���F���g��%|Ǻv�ӺQyߺ=d뺌D������p�R��-�b������$�u*��>0�'6�9�;��A�MG�7M���R�>�X��B^�u�c���i�vro��,u���z��P���-�����舻�Ƌ�~���n���d���D���%���  �  �=Y#=��=�i=�=��=GR=�� =�� =�8 =A��<���<�8�<6z�<��<���<9:�<�x�<x��<V��<A/�<?j�<-��<��<��<pK�<���<Ĵ�<q��<��<�H�<�v�<x��<l��<���<�<�D�<�g�<T��<o��<@��<���<l��<��<��<_.�<�:�<�C�<�I�<�L�<�K�<�F�<o>�<2�<�!�<;�<i��<-��<f��<���<�c�<�3�<���<���<m��<�@�<;��<0��<�S�<���<���<6�<��<�\�<A��<zn�<��<�k�<��<�T�<·<�*�<ǎ�<g�<�I�<ՠ�<��<�B�<=��<�ը<%�<�Z�<���<Eӡ<�
�<@�<tr�<r��<(И<���<'%�<�L�<�r�<�<f��<�ڋ<}��<3�<�6�<�S�<Uo�<f��<�I}<�}y<��u<;�q<Un<_Gj<tyf<�b<��^<�[<&GW<�|S<ܳO<d�K<�&H<�bD<2�@<��<<�$9<k5<,�1<� .<sP*<.�&<��"<$X<��<�<j�<��<�o<��	<�m<��<��;�9�;v�;���;?�;��;��;d��;5�;;��;���;ڈ�;�v�;>y�;y��;��;���;?V�;<Î;1F�;�ރ;};�r;jXh;�7^;AT;�uJ;P�@;�[7;�.;V�$;��;�;KQ
;�;���:��:���:���:�ɱ:�-�:D˒:ݟ�:�Pi:=�K:Ġ.:��:Z��9∲9+�u9��9=,�7>g��:c;�,����ƹ�����!���0� J�k(c��#|�{��tЖ�����E��i���|Ǻ��ӺDyߺ'e뺿D����]r��R�P.���@��_�$�v*��?0�M6���;��A��MG��M�9�R��X�-B^���c�'�i�_ro��,u���z�:P���-���
���舻�Ƌ��������c��wD���%���  �  �=\#=��=�i=�=��=?R=�� =�� =�8 =/��<���<�8�<z�<ٺ�<���<&:�<�x�<i��<D��<./�<>j�<��<$��<��<cK�<���<д�<���<��<�H�<�v�<|��<x��<���<(�<�D�<h�<[��<���<L��<���<���<��<��<R.�<�:�<�C�<�I�<�L�<tK�<�F�<`>�<2�<�!�<"�<R��<��<`��<��<�c�<�3�<���<���<i��<A�<3��<4��<�S�<���<���<6�<4��<�\�<P��<�n�<��<�k�<��<�T�<·<�*�<Ҏ�<�<�I�<Ԡ�<��<�B�<W��<�ը<$�<�Z�<���<8ӡ<�
�<�?�<Tr�<`��<И<���<%�<�L�<�r�<���<e��<�ڋ<���<B�<�6�<�S�<Yo�<���<�I}<�}y<Ӱu<G�q<xn<�Gj<�yf<!�b<�^<�[<JGW<}S<�O<��K<�&H<�bD<�@<��<<%9<�j5<*�1<X .<[P*<	�&<��"<�W<��<s<&�<}�<oo<y�	<�m<u�<|�;�9�;^v�;���;�;	��;�;���;5�;���;뮽;㈷;�v�;�y�;��;=��;���;XV�;�Î;YF�;߃;�};��r;�Xh;&7^; BT;�uJ;�@;�[7;�
.;�$;e�;�;BP
;�;	��:�	�:���:���:ɱ:�,�:�ʒ:���:.Pi:�K:��.:��:���9P��9m�u9�9 ��7B`��];�����i�ƹI���% �B�0���I�$c�~"|��y���ϖ����5F��,i��{Ǻ��Ӻjyߺf��E��U���r� S�S/�j�+���$�dv*�@0��6�d�;���A��MG�AM���R��X�B^�^�c�U�i�&ro��+u���z�"P��H-���
�� 舻>Ƌ�Ԥ��񃑻�c��D���%���  �  �=c#=��=�i=�=��==R=�� =�� =~8 =��<���<�8�<�y�<���<���<:�<�x�<M��</��<!/�<)j�<��<��<��<rK�<π�<ش�<���<��<�H�<�v�<���<���<���<3�<�D�<%h�<~��<���<_��<���<���<��<��<d.�<�:�<�C�<�I�<mL�<gK�<�F�<K>�<�1�<�!�<�<2��<���<>��<ێ�<�c�<�3�<���<���<a��<A�<B��<;��<�S�<���<Ú�<16�<@��<]�<u��<�n�<��<�k�<��<�T�<?·<�*�<쎴<��<�I�<堯<��<�B�<G��<�ը<�<�Z�<���<ӡ<�
�<�?�<Dr�<=��<�Ϙ<~��<%�<�L�<ur�<���<O��<�ڋ<q��<9�<�6�<�S�<fo�<���<�I}<�}y<��u<��q<�n<�Gj<�yf<b�b<A�^<�[<�GW<#}S<�O<��K<�&H<�bD<3�@<��<<�$9<�j5<��1<B .<-P*<У&<��"<�W<~�< <��<G�<Xo<>�	<�m<W�<$�;v9�;v�;���;9�;?��;,�;Ô�;w5�;���;a��;l��;rw�;�y�;4��;½�;}��;�V�;�Î;�F�;B߃;�};7�r;�Xh;�7^;�AT;puJ;��@;�Z7;{
.;'�$;��;�;�O
;�;���:Y�:V��:o��:.Ǳ:�+�:�ɒ:���:Oi:S�K:E�.:{�:P��9���9��u9��9���7�<��8K;�\{���ƹ׿������0�j�I�U#c��|�7y��1ϖ�����E���h��|Ǻ�Ӻ�zߺg�!G��?��?s��S��/�������$�8w*��@0�Y6���;���A�NG��M��R�a�X��A^���c�@�i��qo�O+u�5�z��O���,��
���爻�ŋ�b���]���-c���C��z%���  �  �=k#=��=�i=�=��==R=�� =�� =t8 = ��<���<�8�<�y�<���<���<�9�<�x�<4��< ��</�<j�<��<��<��<lK�<΀�<��<���<��<�H�<w�<���<���<���<V�<�D�<5h�<���<���<��<���<���<��<��<`.�<�:�<�C�<�I�<SL�<`K�<�F�<7>�<�1�<y!�<��<��<���<��<ǎ�<�c�<�3�<���<���<g��<�@�<B��<9��<�S�<
��<Ԛ�<S6�<X��<"]�<���<�n�<��<�k�<��<�T�<Z·<�*�<��<��<�I�<�<��<�B�<:��<�ը<�<�Z�<x��<ӡ<�
�<�?�<4r�<!��<�Ϙ<]��<�$�<�L�<]r�<���<4��<�ڋ<n��</�<�6�<�S�<wo�<���<J}<~y<&�u<��q<�n<Hj<zf<��b<p�^< [<�GW<Y}S<L�O<��K<�&H<�bD<)�@<��<<�$9<�j5<ȳ1<. .<P*<��&<g�"<}W<\�<�<ۈ<��<o<	�	<hm<:�<��;�9�;�u�;x��;�;4��;e�;ޔ�;�5�;&��;���;���;�w�;xz�;���;Q��;���;OW�;Ď;G�;�߃; };ۤr;�Xh;{7^;6AT;nuJ;;�@;Z7;>
.;E�$;
�;|;�N
;>�;H��:>�:��:��:�ű:+�:Ȓ:���:Oi:m�K:��.:�:	��9��9�u9��9!�7���D;��r����ƹ������0�r�I�r c�v|��x��HΖ�����E���h��
}Ǻ��Ӻ�{ߺh��G����t�@U�d0�g����ī$�Mx*�wA0�6���;�}�A�<NG�
M�Y�R���X��A^�g�c���i��po�*u���z�,O���,���	��t爻4ŋ����
����b��rC��%���  �  �=k#=��=�i=�=��=4R=�� =�� =g8 =��<z��<i8�<�y�<s��<���<�9�<dx�< ��<��<�.�<j�<	��<��<��<xK�<р�<��<���<��<�H�<w�<գ�<���<
��<q�<�D�<\h�<���<Ũ�<���<���<���<��<
�<b.�<�:�<�C�<�I�<IL�<@K�<�F�<>�<�1�<Z!�<��<���<���<��<���<�c�<�3�<���<���<X��<�@�<E��<J��<�S�<��<��<a6�<t��<;]�<���<�n�<��<�k�<�<&U�<p·<+�<��<��<�I�<<��<�B�<A��<�ը<��<�Z�<\��<�ҡ<�
�<�?�<r�<���<�Ϙ<A��<�$�<oL�<Fr�<{��<+��<pڋ<o��<4�<�6�<�S�<to�<���<3J}<6~y<X�u<�q<*n<7Hj<Szf<Ǭb<��^<e[<�GW<�}S<b�O<��K<�&H<cD<5�@<��<<�$9<�j5<��1<��-<�O*<��&<A�"<KW<�<�<��<��<�n<��	</m<�<��;-9�;�u�;���;=�;4��;|�;=��;�5�;~��;;-��;Rx�;�z�;��;���;I �;�W�;yĎ;EG�;�߃;�};��r;�Xh;�7^;XAT; uJ;��@;�Y7;4	.;��$;<�;�;�M
;D�;;��:�:��:A��:&ı:)�:&ǒ:ݜ�:�Mi:��K:4�.:��:���9���9��u9�9��79��M1;��n���ƹ�����
�0���I�,c��|��v��g͖�����D���h���|Ǻ؃Ӻk|ߺVi��I�����u��U��1�z	������$��x*�B0��6���;���A��NG��M�*�R�j�X��A^���c�:�i�hpo��)u���z��N���+��D	���戻�ċ�n��������b��&C���$���  �  �=l#=��=�i=�=��=.R=�� =�� =a8 =г�<T��<K8�<�y�<g��<e��<�9�<Bx�<��<���<�.�<j�<���<���<��<�K�<��<���<���<�<�H�<8w�<��<���<)��<��<�D�<}h�<�<��<���<���<���<��<�<[.�<�:�<�C�<�I�<AL�<)K�<�F�<�=�<�1�<8!�<��<���<���<��<���<|c�<p3�<���<���<N��<�@�<;��<Z��<�S�<.��<���<r6�<���<L]�<���<�n�<#�<"l�<�<HU�<�·<0+�<'��<��<�I�< ��<��<�B�<;��<�ը<��<�Z�<J��<�ҡ<�
�<�?�<�q�<���<�Ϙ<"��<�$�<PL�<=r�<b��<(��<fڋ<`��<$�<�6�<�S�<xo�<���<MJ}<`~y<��u<�q<Yn<bHj<�zf<��b<��^<�[<HW<�}S<x�O<�K<�&H<1cD<=�@<��<<�$9<�j5<��1<��-<�O*<E�&<��"<W<ط<�<E�<��<�n<��	<m<��<��;�8�;�u�;.��;[�;}��;��;���;!6�;���;L��;���;�x�;6{�;���;ʾ�;� �;�W�;�Ď;�G�;��;"};��r;bYh;>7^;AT;�tJ;��@;dY7;q.;X�$;%�;�;�L
;��;B��:��:���:���:�ñ:�'�:�ƒ:m��:Li:)�K:��.:��:Z��9���9�v9�
9 �7����;�;j����ƹ������%�0��I��c�|��u���̖����ED���i��:}Ǻ��Ӻ�|ߺIj��J��)��v��V��2��	�|����$�z*�C0�	6���;�ݎA�OG�pM���R�m�X��@^�b�c���i�po�P)u���z�{N���+�����Q戻�ċ����:���b���B���$���  �  �=u#=��=�i=�=��=*R=w� =�� =S8 =���<N��<<8�<�y�<B��<Q��<�9�<<x�<���<���<�.�<�i�<���<���<��<qK�<ހ�< ��<���< �<�H�<Iw�<���<��<F��<��<E�<�h�<Ӊ�<��<���<���<���<��<�<_.�<�:�<�C�<�I�<-L�< K�<gF�<�=�<�1�<+!�<��<���<���<ߴ�<���<^c�<h3�<u��<u��<R��<�@�<D��<E��<�S�<4��<��<�6�<���<^]�<���<"o�<;�<?l�<=�<RU�<�·<;+�<A��<��<J�<��<��<�B�<8��<�ը<��<�Z�<=��<�ҡ<�
�<t?�<�q�<ϡ�<�Ϙ<��<�$�<AL�<r�<[��<��<\ڋ<`��<3�<�6�<�S�<�o�<���<uJ}<�~y<��u<@�q<�n<�Hj<�zf<:�b<�^<�[</HW<�}S<��O<�K<'H<cD<0�@<��<<�$9<�j5<�1<��-<~O*<"�&<��"<�V<��<:<�<g�<�n<��	<�l<��<�;�8�;�u�;f��;�;[��;��;���;x6�;���;���;���;�x�;�{�;璥;J��;� �;X�;Ŏ;�G�;8��;7};%�r;�Xh;W7^;(AT;�tJ;�@;�X7;!.;B�$;��;�;mL
;��;ݘ�:��:��:���:���:'�:�Œ:k��:bLi:�K:��.:��:���9���9d	v9`9o#�7v頸&;��a��X�ƹ�����&�0��I��c�|�cu��|̖�����E���h��~}Ǻ��Ӻ5~ߺ�j��K����Wv�=W�!3��c���$�%z*��C0�
6���;���A�eOG�qM�6�R�~�X��A^���c���i�boo��(u�~�z�4N��3+��k��戻ċ����������a���B��g$���  �  �=~#=��=�i=�=��=)R=o� =�� =L8 =���<5��<#8�<�y�<.��<I��<�9�<#x�<��<���<�.�<�i�<���<���<��<|K�<��<��<���<.�< I�<fw�<��<��<R��<��<3E�<�h�<���<���<���<��<���<��<
�<q.�<�:�<�C�<�I�<!L�<!K�<TF�<�=�<v1�<!�<��<���<���<´�<s��<Kc�<h3�<i��<m��<J��<�@�<X��<M��<�S�<9��<��<�6�<���<�]�<���<;o�<I�<Kl�<W�<lU�<�·<C+�<O��<��<J�<��<��<C�< ��<�ը<��<�Z�<7��<�ҡ<k
�<X?�<�q�<���<|Ϙ<���<�$�<6L�<r�<^��< ��<Zڋ<P��<*�<�6�<�S�<�o�<���<�J}<�~y<ӱu<��q<�n<�Hj<�zf<Y�b<>�^<�[<[HW<�}S<ŴO<
�K<:'H<cD<K�@<��<<�$9<�j5<^�1<��-<bO*<
�&<��"<�V<��<<	�<,�<On<d�	<�l<��<�
�;�8�;(u�;���;9�;���;��;���;�6�;��;���;%��;Vy�;�{�;��;���;*�;�X�;7Ŏ;�G�;k��;0};��r;�Xh;�7^;�@T;ZtJ;��@;UX7;(.;��$;d�;�;�K
;8�;��:� �:;��:���:`��:	'�:�Ē:ܚ�:/Ki::�K:�.:��:g��9��9�v9j9KC�7t���;��[���ƹ[������0���I��c�}|�#u���˖�����D���g��Ǻ��Ӻ�~ߺlk�@L��x��w� X�w3������ݮ$�{*��C0��
6���;��A�wOG��M�z�R���X�jA^�P�c���i��no��(u���z��M���*��'���刻�Ë�q���j����a���B��"$���  �  �=z#=��=�i=�=��=+R=o� =|� =K8 =���<,��<8�<{y�<-��<9��<�9�<x�<��<���<�.�<�i�<���<���<��<wK�<��<��<���<;�<I�<cw�<��<��<`��<��<5E�<�h�<��<��<���<��<���<��<�<d.�<�:�<�C�<�I�<L�<K�<YF�<�=�<s1�<
!�<��<���<y��<���<j��<Pc�<U3�<b��<p��<Q��<�@�<K��<N��<�S�<@��<&��<�6�<���<}]�<���<=o�<a�<_l�<W�<mU�<�·<V+�<[��<��<J�<��<��<�B�<-��<�ը<��<�Z�<(��<�ҡ<f
�<Y?�<�q�<���<oϘ<���<�$�<,L�<r�<H��< ��<[ڋ<Y��<%�<�6�<�S�<�o�<Ǌ�<�J}<�~y<ڱu<m�q<�n<�Hj<{f<j�b<D�^<�[<]HW<�}S<ݴO<-�K<-'H<'cD<7�@<��<<�$9<�j5<^�1<��-<ZO*<��&<��"<�V<p�<<�<,�<?n<`�	<�l<��<�
�;�8�;Fu�;M��;"�;���;��;ݕ�;�6�;Q��;鰽;��;Sy�;|�;t��;���;>�;rX�;eŎ;H�;���;�};{�r;�Xh;v7^;�@T;�tJ;��@;;X7;�.;��$;�;q;WK
;�;���:���:���:���:���:�%�:^Ē:���:�Ki:��K:>�.:��:F��9���9v9�9Y��7�̠�t;��[��Q�ƹ�������0���I��c�|� t���˖����E��i��T~ǺN�Ӻ�~ߺIl�8M��f��Bw�X��3������$�={*�5D0��
6�}�;��A�lOG��M���R�W�X�7A^�w�c��i�~no�5(u���z��M���*����|刻�Ë�f��������a��FB���#���  �  ~=!!=�=�f=i	=��=�M=�� =e� =�2 =���<a��<u*�<�j�<���<���<�'�<be�<��<���<��<�R�<a��<4��<���</�<;c�<���<c��<P��<�%�<�R�<�}�<6��<���<���<^�</:�<�Y�<�v�<���<h��<V��<���<���<{��<���<@�<S�<�<"�<���<y��<f��<i��<A��<��<M��<-b�<�:�<E�<0��<^��<ul�<�,�<���<���<>N�<���< ��<A�<���<bs�<��<��<$�<J��<q�<���<D�<r�<4ܵ<�A�<@��<V �<TY�<Q��<v��<�L�<���<ݦ<8 �<`�<��<$ן<��<cC�<�u�<�<�Ӗ<���<�)�<NR�<�x�<'��<���</�<p�<�%�<�D�<�b�<���<�:}<�sy<��u<!�q<n<�Pj<чf<ξb<|�^<�.[<�gW<?�S<��O<�L<�YH<W�D<7�@<�"=<Qj9<�5<�2<�S.<g�*<� '<u]#<z�<�#<g�<�<s<��<�n
<s�<
�<A <�d�;��;E��;b�;1��;�Z�;��;Ҙ�;�R�;��;���;��;���;*�;�D�;���;�;hQ�;PՊ;n�;L�;K�u;{pk;jKa;`PW;�}M;��C;3T:;%�0;	�';��;��;&;�t;N��:�?�:���:��:���:��:�n�:'$�:�r:�YT:��6:��:�|�9���9ɹ�9�$9<[8%9W��Y!�����Xú� ��� =+�+�D�2(^��Xw�Y/������m����D��?~��Чź��Ѻ��ݺ�麪����� �t�����7��As��N�@&$���)���/�0�5��d;��,A�X�F�+�L�_|R�?X�c ^�M�c��i��@o���t�w�z�k?��p������!���j���Ϣ��ᄑ��g���K���0���  �  ~=)!=�=�f=c	=��=�M=�� =b� =�2 =Χ�<i��<p*�<�j�<���<���<�'�<qe�< ��<���<��<�R�<q��<)��<���<"/�<>c�<��<g��<T��<�%�<�R�<�}�<.��<���<���<b�<:�<�Y�<�v�<���<n��<]��<���<���<���<���<F�<O�<��<$�<���<���<p��<k��<T��<���<Q��<3b�<�:�<H�<2��<=��<jl�<�,�<���<���<@N�<���<
��<	A�<���<cs�<��<���<$�<=��<g�<���<"�<�q�<1ܵ<�A�<E��<b �<YY�<T��<v��<�L�<���<ݦ<  �<`�<��<3ן<��<kC�<�u�<���<�Ӗ<���<*�<SR�<�x�<	��<���</�<c�<�%�<�D�<c�<���<�:}<�sy<��u<�q<�n<�Pj<��f<վb<h�^<�.[<�gW<4�S<��O<�L<�YH<b�D<B�@<r"=<Jj9<��5<�2<�S.<y�*<'<�]#<o�<	$<�<�<s<��<�n
<��<�< <�d�;��;6��;!b�;>��; [�;!��;��;�R�;v�;��;u�;���;��;�D�;<��;��;hQ�;<Պ;n�;l�;��u;�pk;�Ka;�OW;~M;��C;@S:;8�0;�';:�;#�;5;@u;���:@�:6��:��:槶:��:�l�:#�:�r:<XT:Y�6:V�:�~�9K��9޺�9��$9S>[8�KW��i!������ƺ�~���CA+�D�D�{(^��Xw��.����������D��@~����ź��Ѻ��ݺ���L���� �����������r�nN�l&$�s�)���/��5��d;��-A��F�)�L��|R��>X�= ^���c��i��@o� u���z��?���������Y���[�������0���h���K���0���  �  ~='!=�=�f=d	=��=�M=�� =n� =�2 =���<l��<q*�<�j�<���<���<�'�<re�<��<���<��<�R�<���<&��<���< /�<5c�<��<X��<J��<�%�<�R�<�}�<2��<���<���<n�<:�<�Y�<�v�<��<g��<Q��<���<���<���<���<L�<b�< �<<�<���<���<y��<m��<S��<���<S��<9b�<�:�<7�<D��<M��<|l�<�,�<���<���<8N�<���<���<A�<���<_s�<��<���<,�<2��<`�<���<#�<�q�<)ܵ<�A�<8��<\ �<RY�<P��<{��<�L�<���<ݦ<2 �<#`�<��<5ן<��<oC�<�u�<��<�Ӗ<���< *�<GR�<y�<��<���<2�<b�<�%�<�D�<�b�<��<�:}<�sy<��u<�q<�n<�Pj<��f<Ӿb<f�^<�.[<�gW< �S<��O<�L<�YH<O�D<>�@<t"=<Jj9<$�5<�2<�S.<l�*<� '<�]#<q�<$<u�<&�<!s<��<�n
<��<�<9 <&e�;ݩ�;K��;b�;��;[�;���;���;�R�;��;��;��;���;��;�D�;8��;��;dQ�;Պ;n�;;�;i�u;6pk;�Ka;�OW;8~M;2�C;�S:;��0;��';�;k�;P;:u;}��::@�:���:ٜ�:ᦶ:�:�m�:�$�:r:�WT:|�6:`�:}�9���9���9%�$9�6[8�FW��i!�g���ɺ�3�
��&A+���D�z)^��Yw��/�����|����D���}���ź��Ѻ��ݺ�������� �������֒��r�MN�g&$�G�)�S�/�e�5��c;�*-A�q�F��L��|R��>X�� ^���c�Z�i��@o�g u�¿z��?�������������_�������*���h���K���0���  �  ~=$!=�=�f=h	=��=�M=�� =j� =�2 =ԧ�<���<�*�<�j�<���<���<(�<�e�<%��<���<��<�R�<l��<3��<���</�<>c�<���<^��<G��<�%�<yR�<�}�<��<���<���<F�<:�<�Y�<�v�<��<f��<O��<���<���<u��<��<>�<Z�<�<5�<���<���<���<���<_��<��<j��<Pb�<�:�<T�<>��<S��<yl�<�,�<���<���<?N�<���<���< A�<���<Ss�<��<��<�<-��<R�<���<�<�q�<ܵ<�A�<:��<T �<YY�<N��<r��<�L�<���<ݦ<1 �<#`�<��<Dן<��<�C�<�u�<��<Ԗ< �<*�<]R�<y�<"��<���<.�<p�<�%�<�D�<�b�<���<�:}<�sy<��u<��q<�n<�Pj<��f<��b<1�^<�.[<�gW<�S<��O<�L<�YH<_�D<*�@<�"=<Oj9<��5<�2<�S.<��*<'<�]#<��<2$<��<L�<Zs<�<�n
<��<�<J <�d�;��;D��;b�;G��;�Z�;��;���;�R�;%�;���;��;W��;��;aD�;��;{�;7Q�;Պ;n�;7�;��u;�pk;DKa;�PW;�}M;��C;T:;��0;��';m�;�;;�u;m��:�A�:��:���:Ĩ�:��:5n�:�$�:�r:^ZT:��6:S�:�}�9���9��9�$9�![8B}W�m!�p��!ʺ�*!ﹺ��B+�,�D��*^�Zw��/��y��� ����D��e~���ź%�Ѻw�ݺ��麵���:� �i�����0��br��M��%$���)���/���5��c;��,A���F�0�L�a|R�>?X�M ^��c�;�i��@o�| u�=�z��?�� ��8 ����������e���p���ch��L���0���  �  ~=!=�=�f=g	=ī=�M=�� =m� =�2 =��<���<�*�< k�<���<���<
(�<�e�<;��<��<��<�R�<w��<A��<���</�<4c�<��<T��<1��<�%�<gR�<�}�<��<���<x��<6�<:�<�Y�<�v�<ӑ�<U��<F��<{��<���<o��<��<J�<j�<�<;�<���<���<���<���<r��<��<r��<Ub�<�:�<m�<I��<]��<�l�<�,�<���<x��<?N�<���<��<�@�<���<Is�<��<��<��<��<A�<���<�<�q�<ܵ<�A�<+��<? �<IY�<O��<i��<�L�<���<*ݦ<7 �<:`�<6��<Bן<��<�C�<�u�<��<Ԗ< �<*�<yR�<	y�<1��<���<;�<p�<z%�<�D�<�b�<{��<�:}<sy<i�u<��q<�n<|Pj<p�f<�b<4�^<�.[<�gW<��S<y�O<�L<gYH<X�D<'�@<�"=<kj9<�5<�2<�S.<ɨ*<1'<�]#<��<Q$<͎<d�<es<�<�n
<��<�<m <e�;V��;/��;b�;%��;�Z�;���;a��;�R�;��;���;��;��;��;&D�;!��;S�;
Q�;�Ԋ;�m�;�;۾u;�pk;Ka;�PW;3~M;y�C;pT:;��0;V�';��;-�;X;8v;���:CB�:l��: ��:`��:��:�n�:�%�:#r:�[T:
�6:}�:y�9���9���9�}$9k[8�W�;m!�c���ͺ�/%�p���B+�x�D��+^��\w�e0�����������D���~���ź}�Ѻo�ݺb��D���s� �t�����ۑ��q�qM�N%$���)�a�/�ԗ5��c;�e,A���F�ʸL�b|R�k?X�` ^���c�z�i��Ao�� u���z�@�����| �������\��������h��<L��91���  �  �}=!=�=�f=f	=ë=�M=�� =|� =�2 =��<���<�*�<k�<Ū�<���<%(�<�e�<;��<��<��<�R�<���<4��<���</�<*c�<��<I��<)��<�%�<]R�<�}�< ��<���<W��<4�<�9�<tY�<�v�<ɑ�<N��<E��<|��<���<|��<���<X�<m�<�<[�<���<���<���<���<���<+��<���<ub�<�:�<_�<g��<j��<�l�<�,�<���<���<1N�<���<��<�@�<���<-s�<��<���<��<���<'�<{��<��<�q�<�۵<�A�<��<D �<AY�<H��<o��<�L�<���<&ݦ<I �<K`�<0��<gן<��<�C�<v�<4��</Ԗ<- �<.*�<oR�<(y�<1��<���<A�<l�<�%�<�D�<�b�<u��<�:}<asy<?�u<��q<�n<jPj<(�f<d�b<��^<D.[<}gW<ءS<m�O<�L<wYH<>�D<2�@<~"=<gj9<$�5<�2<.T.<��*<D'<^#<�<�$<ڎ<��<�s<e�<�n
<��<N�<h <Ae�;(��;K��;b�;��;�Z�;���;H��;DR�;��;b��;��;���;�;"D�;u��;�;�P�;�Ԋ;�m�;�;�u;&pk;�Ka;TPW;�~M;��C;�T:;�0;��';��;;�;$;�v;���:�C�:x��:��:���:��:�o�:�%�:$ r:7YT:��6:��:�x�9���9/��9Ly$9c�Z8H�W���!�E��Vպ�+�]���G+���D�H.^��]w�1��H���E���E��k~���ź��Ѻ��ݺ4������� �H�������nq��L�|$$�v�)���/�&�5��b;�d,A�W�F���L��|R�?X�� ^���c���i��Ao�ou�H�z��@��� ��� ��oሻ:�ˣ�������h���L��Q1���  �  �}=!=�=�f=h	=ƫ=�M=�� =�� =�2 =
��<���<�*�<5k�<��<���<%(�<�e�<R��<��<��<�R�<���<5��<���</�<*c�<��<,��<*��<s%�<UR�<l}�<ަ�<���<C��<�<�9�<rY�<�v�<đ�<:��<,��<���<���<���<���<d�<u�<�<m�<���<���<���<���<���<E��<���<pb�<�:�<q�<w��<l��<�l�<�,�<���<���<#N�<���<֟�<�@�<���<s�<��<���<��<晽<�<Z��<��<�q�<�۵<�A�<��<7 �<AY�<>��<y��<�L�<ϖ�<)ݦ<Q �<Z`�<D��<zן<��<�C�<v�<P��<;Ԗ<2 �<L*�<�R�<7y�<4��<���<G�<l�<�%�<�D�<�b�<W��<�:}<?sy<�u<��q<En<IPj<��f<H�b<��^<..[<`gW<��S<e�O<gL<wYH</�D<1�@<�"=<qj9<K�5<�2<HT.<�*<�'<!^#<��<�$<�<��<�s<��<o
<�<i�<t <�e�;1��;v��;b�;	��;�Z�;N��;R��;�Q�;��;��;L�;���;��;�C�;���;�;RP�;�Ԋ;am�;��;%�u;�ok;�Ka;FPW;M;��C;�T:;��0;��';s�;7�;�;�w;B��:GE�:C��:���:���:��:�o�:�%�:"r:�XT:��6:f�:Az�9���9���9 y$9S�Z8޽W�N�!���uں�./�A���J+�[�D�-2^��]w��2�����*����E���}��"�źb�ѺU�ݺ���&����� �������;���p��K�$$�J�)���/���5�_b;�O,A���F�p�L�~|R��>X�^��c���i�Bo��u���z��@��!��� ���ሻr�W���*���i���L��`1���  �  �}=!=	�=�f=i	=ɫ=�M=�� =�� =�2 =��<���<�*�<Bk�<���<��<G(�<�e�<f��<,��<��<�R�<���<?��<���</�<#c�<ٕ�<)��<��<`%�<7R�<i}�<Ц�<r��<(��<�<�9�<]Y�<�v�<���<3��<(��<p��<���<x��< ��<`�<��<7�<h�<��<���<���<���<���<X��<���<�b�<�:�<��<t��<���<�l�<�,�<���<��<$N�<���<џ�<�@�<���<�r�<i�<���<��<ʙ�<��<E��<��<�q�<�۵<�A�< ��<, �<6Y�<>��<q��<�L�<ǖ�<Cݦ<b �<a`�<[��<|ן<��<�C�<1v�<\��<]Ԗ<F �<V*�<�R�<7y�<Q��<���<I�<q�<�%�<�D�<�b�<S��<t:}<sy<�u<d�q<@n<Pj<Ȇf<�b<��^<.[<$gW<��S<K�O<`L<OYH<&�D<&�@<�"=<|j9<N�5<32<MT.<�*<�'<>^#<C�<�$<=�<��<�s<��<Ao
<,�<��<� <�e�;`��;k��;b�;���;�Z�;K��;��;�Q�;6�;��;�;1��;U�;dC�;��;��;P�;LԊ;Jm�;��;��u;�ok;vKa;�PW;�~M;W�C;�U:;x�0;��';��;	�;�;7x;���:G�:��:���:���:q�:gq�:'�:T!r:�ZT:q�6:��:@v�92��9l��9q$9}Z8��W�J�!����ẹ�5﹕���J+���D��4^��_w��2����������|E��~��s�ź��Ѻ��ݺ��麦���9� �����������o�kK�#$���)���/���5�^b;�d+A���F�`�L�Y|R�@?X�)^��c���i��Bo�uu���z��@��!��U��-∻��r���c����i�� M���1���  �  �}=!=�=�f=g	=ϫ=�M=�� =�� =�2 =%��<���<�*�<Qk�<��<��<n(�<�e�<{��<:��< �<�R�<���<M��<���</�<c�<ҕ�<(��<���<l%�<$R�<G}�<���<Z��< ��<��<�9�<8Y�<�v�<���<!��<)��<a��<���<n��<��<e�<|�<A�<r�<��<���<���<���<Ǿ�<t��<���<�b�<�:�<��<}��<���<�l�<�,�<���<r��<6N�<���<ϟ�<�@�<r��<s�<E�<}��<��<���<��<*��<��<q�<�۵<�A�<���<% �<(Y�<H��<c��<�L�<Ŗ�<Dݦ<g �<j`�<p��<�ן<�<�C�<Sv�<p��<mԖ<g �<`*�<�R�<>y�<\��<���<U�<r�<}%�<�D�<�b�<W��<C:}<sy<�u<�q<n<�Oj<��f<۽b<x�^<�-[<gW<��S<�O<dL<7YH<0�D<%�@<�"=<�j9<>�5<E2<YT.<?�*<�'<{^#<u�<�$<��<	�<8t<��<no
<I�<��<� <ze�;���;C��;0b�;���;qZ�;K��;���;�Q�;��;���;��;���;9�;C�;���;#�;(P�;�ӊ;m�;��;)�u;�pk;2Ka;�PW;$M;*�C;�U:;��0;K�';�;b�;�; y;J��:NG�:���:���:L��:�:�q�:�&�:�!r:�[T:�6:(�:;r�9ӿ�9���9�b$9>�Z8*1X�=�!�)���㺹�:�ː��N+� �D�3^��cw�23��ꠔ������D���~����ź��Ѻ��ݺ������� ����c��x���n��J��"$���)�I�/���5�%b;�+A���F��L�U|R�Z?X�� ^���c���i�DCo��u���z�vA��z!�����A∻HË�Ϥ��􆑻�i��M��2���  �  �}=!=�=�f=h	=ѫ=�M=�� =�� =�2 =4��<���<�*�<ck�<*��<$��<i(�<�e�<���<J��<�<�R�<���<O��<���</�<c�<ƕ�<��<���<Q%�<R�<C}�<���<J��<	��<��<�9�<:Y�<�v�<���<��<��<U��<���<v��<��<u�<��<O�<��<��<���<���<���<׾�<���<ȅ�<�b�<�:�<��<���<���<�l�<�,�<���<x��<*N�<}��<���<�@�<b��<�r�<B�<v��<��<���<��< ��<��<sq�<�۵<~A�<碲< �<Y�<C��<i��<�L�<ۖ�<Kݦ<x �<}`�<|��<�ן<�<�C�<dv�<���<mԖ<m �<r*�<�R�<Vy�<f��<<\�<p�<�%�<�D�<�b�<H��<7:}<�ry<��u<�q<n<�Oj<��f<��b<i�^<�-[<�fW<P�S<�O<HL<&YH<�D<+�@<�"=<�j9<n�5<W2<�T.<Z�*<�'<�^#<t�<!%<��<,�</t<��<�o
<l�<��<� <�e�;���;d��;2b�;���;EZ�;��;���;SQ�;��;~��;��;���;��;�B�;���;/�;�O�;�ӊ;�l�;u�;ؽu;pk;xKa;�PW;�M;��C;lV:;��0;��';��;x�;1;�y;?��:�G�:���:���:Ǯ�:���:�r�:�'�:$r:�[T:��6:��:>o�9���9U��9[[$9�`Z8�4X�Ԣ!�o��?麹�?�ӑ�GO+�G�D�!6^�ndw�4��ܡ��[���E��x~����źs�Ѻ �ݺ���Ǿ��!� ���������]n�@J��"$�j�)���/���5�ga;��*A�3�F�ȷL�f|R�0?X�A^���c��i�vCo�{u�J�z�xA���!������∻�Ë�줎������i���M��2���  �  �}=!=�=�f=l	=ͫ=�M=�� =�� = 3 =H��<���<+�<xk�<&��<F��<{(�<�e�<���<M��<�<�R�<���<E��<���<
/�<c�<ӕ�<��<���<8%�<R�</}�<���<?��<���<��<�9�<+Y�<qv�<���<��<��<k��<���<���<��<n�<��<M�<��<)��<��<���<
��<��<���<��<�b�<;�<��<���<���<�l�<�,�<���<���<N�<���<���<�@�<d��<�r�<3�<]��<|�<���<��<��<��<eq�<�۵<�A�<ߢ�< �<%Y�<.��<t��<�L�<ؖ�<Jݦ<z �<`�<���<�ן<�<D�<cv�<���<�Ԗ<y �<�*�<�R�<Yy�<_��<<S�<v�<�%�<�D�<�b�<?��<A:}<�ry<��u<��q<�n<�Oj<g�f<��b<2�^<�-[<�fW<4�S<�O<4L<NYH<�D<�@<�"=<�j9<{�5<I2<�T.<b�*<'<�^#<��<M%<��<q�<Ut<�<�o
<t�<ȃ<� <�e�;���;���;�a�;���;�Z�;���;���;�P�;��;3��;6�;q��;��;�B�;'��;���;^O�;�ӊ;�l�;n�;��u;�ok;�Ka;�PW;|M;��C;cV:;��0;��';k�;��;g;�y;���:�J�:F��:Y��:k��:���:�r�:)(�:�#r:�ZT:��6:�:yt�9���9�9]$9&Z8QX��!�> ��*�rB�
���Q+���D��9^�zcw��4��0�������FF���}��/�ź��Ѻ �ݺ��麟����� ���������gn��I�o!$��)��/�w�5�Ma;��*A��F��L�5|R�,?X��^�*�c�U�i�KCo��u���z��A���!��+���∻�Ë�X���P���3j���M�� 2���  �  �}=!=�=�f=m	=ҫ=�M=�� =�� =3 =I��<���<+�<{k�<9��<?��<}(�<�e�<���<Y��<�<�R�<���<Q��<���</�<c�<���< ��<���<F%�<R�<)}�<���<<��<���<��<9�<)Y�<�v�<���<��<��<^��<���<{��<	��<s�<��<X�<��<0��<��<���<��<��<���<��<�b�<;�<��<���<���<�l�<�,�<���<���<N�<���<���<�@�<T��<�r�<3�<V��<y�<���<��<��<��<lq�<�۵<jA�<͢�<	 �<Y�</��<s��<�L�<ݖ�<Wݦ< �<�`�<���<�ן<�<D�<rv�<���<�Ԗ<u �<�*�<�R�<by�<n��<<]�<y�<~%�<�D�<�b�</��<:}<�ry<��u<��q<�n<�Oj<p�f<��b<1�^<�-[<�fW<;�S<��O<L<&YH<�D<�@<�"=<�j9<��5<h2<�T.<s�*<'<�^#<��<S%<ˏ<e�<Yt<�<�o
<��<҃<� <f�;���;���;�a�;���;0Z�;���;P��;/Q�;��;��;3�;g��;��;�B�;��;���;�O�;�ӊ;�l�;)�;&�u;�ok;�Ka;�PW;�M;0�C;�V:;��0;�';B�;��;0;z;2��:J�:W��: ��:¯�:K��:ks�:�(�:V$r:�[T:F�6:��:r�93��9���9bU$9BFZ8BNX���!�� ���캹�B�Z���R+���D��7^��fw��5��v�������.F���}��k�ź4�Ѻ1�ݺ���׽���� ���������m��I��!$�*�)��/�5�5�a;�}*A���F���L�|R�M?X��^���c�ڃi��Co��u�s�z��A��"��H���∻�Ë�[���X����i���M��]2���  �  �}=!=�=�f=j	=ϫ=�M=�� =�� =3 =S��<	��<+�<zk�<G��<9��<�(�<f�<���<a��<�<�R�<���<N��<���</�<c�<���<��<���<B%�<�Q�<}�<���<+��<���<��<�9�<Y�<zv�<{��< ��<��<O��<���<y��<��<m�<��<R�<��<2��<��<��<��<��<���<��<�b�<;�<��<���<���<�l�<�,�<���<}��<$N�<y��<���<�@�<R��<�r�<$�<S��<t�<���<��<��<{�<Wq�<�۵<gA�<좲<
 �<Y�<>��<m��<�L�<Җ�<Oݦ<x �<�`�<���<�ן<5�<�C�<�v�<���<�Ԗ<� �<�*�<�R�<_y�<l��<<Z�<u�<�%�<�D�<�b�<F��<2:}<�ry<��u<��q<�n<}Oj<[�f<t�b<7�^<-[<�fW<&�S<��O<GL<
YH<�D</�@<�"=<�j9<c�5<e2<�T.<}�*<'<�^#<��<Q%<�<X�<|t<,�<�o
<��<ƃ<� <�e�;���;���;8b�;���; Z�;4��;R��;"Q�;\�;���;F�;'��;u�;oB�;��;���;�O�;tӊ;m�;c�;��u;(pk;�Ka;�PW;uM;��C;�V:;��0;%�';��;��;T;lz;��:J�:a��:���:���:c��:&s�:(�:R#r:H[T:��6:E�:�n�9!��9���9cT$9�?Z8�lX���!�
"��z�*G�E��BT+���D�8^��fw��3��c���!���5E��~����ź��Ѻ��ݺ���g����� �m��M��E��rm�pI�O!$�B�)���/��5�a;��*A�N�F�ڷL�<|R�?X�4^�/�c�!�i��Co�u���z�B���!��r��㈻ċ�M�������Gj���M��92���  �  �}=!=�=�f=m	=ҫ=�M=�� =�� =3 =I��<���<+�<{k�<9��<?��<}(�<�e�<���<Y��<�<�R�<���<Q��<���</�<c�<���< ��<���<F%�<R�<)}�<���<<��<���<��<9�<)Y�<�v�<���<��<��<^��<���<{��<	��<s�<��<X�<��<0��<��<���<��<��<���<��<�b�<;�<��<���<���<�l�<�,�<���<���<N�<���<���<�@�<T��<�r�<3�<V��<y�<���<��<��<��<lq�<�۵<jA�<͢�<	 �<Y�</��<s��<�L�<ݖ�<Wݦ< �<�`�<���<�ן<�<D�<rv�<���<�Ԗ<u �<�*�<�R�<by�<n��<<]�<y�<~%�<�D�<�b�</��<:}<�ry<��u<��q<�n<�Oj<p�f<��b<1�^<�-[<�fW<;�S<��O<L<&YH<�D<�@<�"=<�j9<��5<h2<�T.<s�*<'<�^#<��<S%<ˏ<e�<Yt<�<�o
<��<҃<� <f�;���;���;�a�;���;0Z�;���;P��;/Q�;��;��;3�;g��;��;�B�;��;���;�O�;�ӊ;�l�;)�;&�u;�ok;�Ka;�PW;�M;0�C;�V:;��0;�';B�;��;0;z;2��:J�:W��: ��:¯�:K��:ks�:�(�:V$r:�[T:F�6:��:r�93��9���9bU$9BFZ8BNX���!�� ���캹�B�Z���R+���D��7^��fw��5��v�������.F���}��k�ź4�Ѻ1�ݺ���׽���� ���������m��I��!$�*�)��/�5�5�a;�}*A���F���L�|R�M?X��^���c�ڃi��Co��u�s�z��A��"��H���∻�Ë�[���X����i���M��]2���  �  �}=!=�=�f=l	=ͫ=�M=�� =�� = 3 =H��<���<+�<xk�<&��<F��<{(�<�e�<���<M��<�<�R�<���<E��<���<
/�<c�<ӕ�<��<���<8%�<R�</}�<���<?��<���<��<�9�<+Y�<qv�<���<��<��<k��<���<���<��<n�<��<M�<��<)��<��<���<
��<��<���<��<�b�<;�<��<���<���<�l�<�,�<���<���<N�<���<���<�@�<d��<�r�<3�<]��<|�<���<��<��<��<eq�<�۵<�A�<ߢ�< �<%Y�<.��<t��<�L�<ؖ�<Jݦ<z �<`�<���<�ן<�<D�<cv�<���<�Ԗ<y �<�*�<�R�<Yy�<_��<<S�<v�<�%�<�D�<�b�<?��<A:}<�ry<��u<��q<�n<�Oj<g�f<��b<2�^<�-[<�fW<4�S<�O<4L<NYH<�D<�@<�"=<�j9<{�5<I2<�T.<b�*<'<�^#<��<M%<��<q�<Ut<�<�o
<t�<ȃ<� <�e�;���;���;�a�;���;�Z�;���;���;�P�;��;3��;6�;q��;��;�B�;'��;���;^O�;�ӊ;�l�;n�;��u;�ok;�Ka;�PW;|M;��C;cV:;��0;��';k�;��;g;�y;���:�J�:F��:Y��:k��:���:�r�:)(�:�#r:�ZT:��6:�:yt�9���9�9]$9&Z8QX��!�> ��*�rB�
���Q+���D��9^�zcw��4��0�������FF���}��/�ź��Ѻ �ݺ��麟����� ���������gn��I�o!$��)��/�w�5�Ma;��*A��F��L�5|R�,?X��^�*�c�U�i�KCo��u���z��A���!��+���∻�Ë�X���P���3j���M�� 2���  �  �}=!=�=�f=h	=ѫ=�M=�� =�� =�2 =4��<���<�*�<ck�<*��<$��<i(�<�e�<���<J��<�<�R�<���<O��<���</�<c�<ƕ�<��<���<Q%�<R�<C}�<���<J��<	��<��<�9�<:Y�<�v�<���<��<��<U��<���<v��<��<u�<��<O�<��<��<���<���<���<׾�<���<ȅ�<�b�<�:�<��<���<���<�l�<�,�<���<x��<*N�<}��<���<�@�<b��<�r�<B�<v��<��<���<��< ��<��<sq�<�۵<~A�<碲< �<Y�<C��<i��<�L�<ۖ�<Kݦ<x �<}`�<|��<�ן<�<�C�<dv�<���<mԖ<m �<r*�<�R�<Vy�<f��<<\�<p�<�%�<�D�<�b�<H��<7:}<�ry<��u<�q<n<�Oj<��f<��b<i�^<�-[<�fW<P�S<�O<HL<&YH<�D<+�@<�"=<�j9<n�5<W2<�T.<Z�*<�'<�^#<t�<!%<��<,�</t<��<�o
<l�<��<� <�e�;���;d��;2b�;���;EZ�;��;���;SQ�;��;~��;��;���;��;�B�;���;/�;�O�;�ӊ;�l�;u�;ؽu;pk;xKa;�PW;�M;��C;lV:;��0;��';��;x�;1;�y;?��:�G�:���:���:Ǯ�:���:�r�:�'�:$r:�[T:��6:��:>o�9���9U��9[[$9�`Z8�4X�Ԣ!�o��?麹�?�ӑ�GO+�G�D�!6^�ndw�4��ܡ��[���E��x~����źs�Ѻ �ݺ���Ǿ��!� ���������]n�@J��"$�j�)���/���5�ga;��*A�3�F�ȷL�f|R�0?X�A^���c��i�vCo�{u�J�z�xA���!������∻�Ë�줎������i���M��2���  �  �}=!=�=�f=g	=ϫ=�M=�� =�� =�2 =%��<���<�*�<Qk�<��<��<n(�<�e�<{��<:��< �<�R�<���<M��<���</�<c�<ҕ�<(��<���<l%�<$R�<G}�<���<Z��< ��<��<�9�<8Y�<�v�<���<!��<)��<a��<���<n��<��<e�<|�<A�<r�<��<���<���<���<Ǿ�<t��<���<�b�<�:�<��<}��<���<�l�<�,�<���<r��<6N�<���<ϟ�<�@�<r��<s�<E�<}��<��<���<��<*��<��<q�<�۵<�A�<���<% �<(Y�<H��<c��<�L�<Ŗ�<Dݦ<g �<j`�<p��<�ן<�<�C�<Sv�<p��<mԖ<g �<`*�<�R�<>y�<\��<���<U�<r�<}%�<�D�<�b�<W��<C:}<sy<�u<�q<n<�Oj<��f<۽b<x�^<�-[<gW<��S<�O<dL<7YH<0�D<%�@<�"=<�j9<>�5<E2<YT.<?�*<�'<{^#<u�<�$<��<	�<8t<��<no
<I�<��<� <ze�;���;C��;0b�;���;qZ�;K��;���;�Q�;��;���;��;���;9�;C�;���;#�;(P�;�ӊ;m�;��;)�u;�pk;2Ka;�PW;$M;*�C;�U:;��0;K�';�;b�;�; y;J��:NG�:���:���:L��:�:�q�:�&�:�!r:�[T:�6:(�:;r�9ӿ�9���9�b$9>�Z8*1X�=�!�)���㺹�:�ː��N+� �D�3^��cw�23��ꠔ������D���~����ź��Ѻ��ݺ������� ����c��x���n��J��"$���)�I�/���5�%b;�+A���F��L�U|R�Z?X�� ^���c���i�DCo��u���z�vA��z!�����A∻HË�Ϥ��􆑻�i��M��2���  �  �}=!=	�=�f=i	=ɫ=�M=�� =�� =�2 =��<���<�*�<Bk�<���<��<G(�<�e�<f��<,��<��<�R�<���<?��<���</�<#c�<ٕ�<)��<��<`%�<7R�<i}�<Ц�<r��<(��<�<�9�<]Y�<�v�<���<3��<(��<p��<���<x��< ��<`�<��<7�<h�<��<���<���<���<���<X��<���<�b�<�:�<��<t��<���<�l�<�,�<���<��<$N�<���<џ�<�@�<���<�r�<i�<���<��<ʙ�<��<E��<��<�q�<�۵<�A�< ��<, �<6Y�<>��<q��<�L�<ǖ�<Cݦ<b �<a`�<[��<|ן<��<�C�<1v�<\��<]Ԗ<F �<V*�<�R�<7y�<Q��<���<I�<q�<�%�<�D�<�b�<S��<t:}<sy<�u<d�q<@n<Pj<Ȇf<�b<��^<.[<$gW<��S<K�O<`L<OYH<&�D<&�@<�"=<|j9<N�5<32<MT.<�*<�'<>^#<C�<�$<=�<��<�s<��<Ao
<,�<��<� <�e�;`��;k��;b�;���;�Z�;K��;��;�Q�;6�;��;�;1��;U�;dC�;��;��;P�;LԊ;Jm�;��;��u;�ok;vKa;�PW;�~M;W�C;�U:;x�0;��';��;	�;�;7x;���:G�:��:���:���:q�:gq�:'�:T!r:�ZT:q�6:��:@v�92��9l��9q$9}Z8��W�J�!����ẹ�5﹕���J+���D��4^��_w��2����������|E��~��s�ź��Ѻ��ݺ��麦���9� �����������o�kK�#$���)���/���5�^b;�d+A���F�`�L�Y|R�@?X�)^��c���i��Bo�uu���z��@��!��U��-∻��r���c����i�� M���1���  �  �}=!=�=�f=h	=ƫ=�M=�� =�� =�2 =
��<���<�*�<5k�<��<���<%(�<�e�<R��<��<��<�R�<���<5��<���</�<*c�<��<,��<*��<s%�<UR�<l}�<ަ�<���<C��<�<�9�<rY�<�v�<đ�<:��<,��<���<���<���<���<d�<u�<�<m�<���<���<���<���<���<E��<���<pb�<�:�<q�<w��<l��<�l�<�,�<���<���<#N�<���<֟�<�@�<���<s�<��<���<��<晽<�<Z��<��<�q�<�۵<�A�<��<7 �<AY�<>��<y��<�L�<ϖ�<)ݦ<Q �<Z`�<D��<zן<��<�C�<v�<P��<;Ԗ<2 �<L*�<�R�<7y�<4��<���<G�<l�<�%�<�D�<�b�<W��<�:}<?sy<�u<��q<En<IPj<��f<H�b<��^<..[<`gW<��S<e�O<gL<wYH</�D<1�@<�"=<qj9<K�5<�2<HT.<�*<�'<!^#<��<�$<�<��<�s<��<o
<�<i�<t <�e�;1��;v��;b�;	��;�Z�;N��;R��;�Q�;��;��;L�;���;��;�C�;���;�;RP�;�Ԋ;am�;��;%�u;�ok;�Ka;FPW;M;��C;�T:;��0;��';s�;7�;�;�w;B��:GE�:C��:���:���:��:�o�:�%�:"r:�XT:��6:f�:Az�9���9���9 y$9S�Z8޽W�N�!���uں�./�A���J+�[�D�-2^��]w��2�����*����E���}��"�źb�ѺU�ݺ���&����� �������;���p��K�$$�J�)���/���5�_b;�O,A���F�p�L�~|R��>X�^��c���i�Bo��u���z��@��!��� ���ሻr�W���*���i���L��`1���  �  �}=!=�=�f=f	=ë=�M=�� =|� =�2 =��<���<�*�<k�<Ū�<���<%(�<�e�<;��<��<��<�R�<���<4��<���</�<*c�<��<I��<)��<�%�<]R�<�}�< ��<���<W��<4�<�9�<tY�<�v�<ɑ�<N��<E��<|��<���<|��<���<X�<m�<�<[�<���<���<���<���<���<+��<���<ub�<�:�<_�<g��<j��<�l�<�,�<���<���<1N�<���<��<�@�<���<-s�<��<���<��<���<'�<{��<��<�q�<�۵<�A�<��<D �<AY�<H��<o��<�L�<���<&ݦ<I �<K`�<0��<gן<��<�C�<v�<4��</Ԗ<- �<.*�<oR�<(y�<1��<���<A�<l�<�%�<�D�<�b�<u��<�:}<asy<?�u<��q<�n<jPj<(�f<d�b<��^<D.[<}gW<ءS<m�O<�L<wYH<>�D<2�@<~"=<gj9<$�5<�2<.T.<��*<D'<^#<�<�$<ڎ<��<�s<e�<�n
<��<N�<h <Ae�;(��;J��;b�;��;�Z�;���;H��;DR�;��;b��;��;���;�;"D�;u��;�;�P�;�Ԋ;�m�;�;�u;&pk;�Ka;TPW;�~M;��C;�T:;�0;��';��;;�;$;�v;���:�C�:x��:��:���:��:�o�:�%�:$ r:7YT:��6:��:�x�9���9/��9Ly$9c�Z8H�W���!�E��Vպ�+�]���G+���D�H.^��]w�1��H���E���E��k~���ź��Ѻ��ݺ4������� �H�������nq��L�|$$�v�)���/�&�5��b;�d,A�W�F���L��|R�?X�� ^���c���i��Ao�ou�H�z��@��� ��� ��oሻ:�ˣ�������h���L��Q1���  �  ~=!=�=�f=g	=ī=�M=�� =m� =�2 =��<���<�*�< k�<���<���<
(�<�e�<;��<��<��<�R�<w��<A��<���</�<4c�<��<T��<1��<�%�<gR�<�}�<��<���<x��<6�<:�<�Y�<�v�<ӑ�<U��<F��<{��<���<o��<��<J�<j�<�<;�<���<���<���<���<r��<��<r��<Ub�<�:�<m�<I��<]��<�l�<�,�<���<x��<?N�<���<��<�@�<���<Is�<��<��<��<��<A�<���<�<�q�<ܵ<�A�<+��<? �<IY�<O��<i��<�L�<���<*ݦ<7 �<:`�<6��<Bן<��<�C�<�u�<��<Ԗ< �<*�<yR�<	y�<1��<���<;�<p�<z%�<�D�<�b�<{��<�:}<sy<i�u<��q<�n<|Pj<p�f<�b<4�^<�.[<�gW<��S<y�O<�L<gYH<X�D<'�@<�"=<kj9<�5<�2<�S.<ɨ*<1'<�]#<��<Q$<͎<d�<es<�<�n
<��<�<m <e�;V��;/��;b�;%��;�Z�;���;a��;�R�;��;���;��;��;��;&D�;!��;S�;
Q�;�Ԋ;�m�;�;۾u;�pk;Ka;�PW;3~M;y�C;pT:;��0;V�';��;-�;X;8v;���:CB�:l��: ��:`��:��:�n�:�%�:#r:�[T:
�6:}�:y�9���9���9�}$9k[8�W�;m!�c���ͺ�/%�p���B+�x�D��+^��\w�e0�����������D���~���ź}�Ѻo�ݺb��D���s� �t�����ۑ��q�qM�N%$���)�a�/�ԗ5��c;�e,A���F�ʸL�b|R�k?X�` ^���c�z�i��Ao�� u���z�@�����| �������\��������h��<L��91���  �  ~=$!=�=�f=h	=��=�M=�� =j� =�2 =ԧ�<���<�*�<�j�<���<���<(�<�e�<%��<���<��<�R�<l��<3��<���</�<>c�<���<^��<G��<�%�<yR�<�}�<��<���<���<F�<:�<�Y�<�v�<��<f��<O��<���<���<u��<��<>�<Z�<�<5�<���<���<���<���<_��<��<j��<Pb�<�:�<T�<>��<S��<yl�<�,�<���<���<?N�<���<���< A�<���<Ss�<��<��<�<-��<R�<���<�<�q�<ܵ<�A�<:��<T �<YY�<N��<r��<�L�<���<ݦ<1 �<#`�<��<Dן<��<�C�<�u�<��<Ԗ< �<*�<]R�<y�<"��<���<.�<p�<�%�<�D�<�b�<���<�:}<�sy<��u<��q<�n<�Pj<��f<��b<1�^<�.[<�gW<�S<��O<�L<�YH<_�D<*�@<�"=<Oj9<��5<�2<�S.<��*<'<�]#<��<2$<��<L�<Zs<�<�n
<��<�<J <�d�;��;D��;b�;G��;�Z�;��;���;�R�;%�;���;��;W��;��;aD�;��;{�;7Q�;Պ;n�;7�;��u;�pk;DKa;�PW;�}M;��C;T:;��0;��';m�;�;;�u;m��:�A�:��:���:Ĩ�:��:5n�:�$�:�r:^ZT:��6:S�:�}�9���9��9�$9�![8B}W�m!�p��!ʺ�*!ﹺ��B+�,�D��*^�Zw��/��y��� ����D��e~���ź%�Ѻw�ݺ��麵���:� �i�����0��br��M��%$���)���/���5��c;��,A���F�0�L�a|R�>?X�M ^��c�;�i��@o�| u�=�z��?�� ��8 ����������e���p���ch��L���0���  �  ~='!=�=�f=d	=��=�M=�� =n� =�2 =���<l��<q*�<�j�<���<���<�'�<re�<��<���<��<�R�<���<&��<���< /�<5c�<��<X��<J��<�%�<�R�<�}�<2��<���<���<n�<:�<�Y�<�v�<��<g��<Q��<���<���<���<���<L�<b�< �<<�<���<���<y��<m��<S��<���<S��<9b�<�:�<7�<D��<M��<|l�<�,�<���<���<8N�<���<���<A�<���<_s�<��<���<,�<2��<`�<���<#�<�q�<)ܵ<�A�<8��<\ �<RY�<P��<{��<�L�<���<ݦ<2 �<#`�<��<5ן<��<oC�<�u�<��<�Ӗ<���< *�<GR�<y�<��<���<2�<b�<�%�<�D�<�b�<��<�:}<�sy<��u<�q<�n<�Pj<��f<Ӿb<f�^<�.[<�gW< �S<��O<�L<�YH<O�D<>�@<t"=<Jj9<$�5<�2<�S.<l�*<� '<�]#<q�<$<u�<&�<!s<��<�n
<��<�<9 <&e�;ݩ�;K��;b�;��;[�;���;���;�R�;��;��;��;���;��;�D�;8��;��;dQ�;Պ;n�;;�;i�u;6pk;�Ka;�OW;8~M;2�C;�S:;��0;��';�;k�;P;:u;}��::@�:���:ٜ�:ᦶ:�:�m�:�$�:r:�WT:|�6:`�:}�9���9���9%�$9�6[8�FW��i!�g���ɺ�3�
��&A+���D�z)^��Yw��/�����|����D���}���ź��Ѻ��ݺ�������� �������֒��r�MN�g&$�G�)�S�/�e�5��c;�*-A�q�F��L��|R��>X�� ^���c�Z�i��@o�g u�¿z��?�������������_�������*���h���K���0���  �  ~=)!=�=�f=c	=��=�M=�� =b� =�2 =Χ�<i��<p*�<�j�<���<���<�'�<qe�< ��<���<��<�R�<q��<)��<���<"/�<>c�<��<g��<T��<�%�<�R�<�}�<.��<���<���<b�<:�<�Y�<�v�<���<n��<]��<���<���<���<���<F�<O�<��<$�<���<���<p��<k��<T��<���<Q��<3b�<�:�<H�<2��<=��<jl�<�,�<���<���<@N�<���<
��<	A�<���<cs�<��<���<$�<=��<g�<���<"�<�q�<1ܵ<�A�<E��<b �<YY�<T��<v��<�L�<���<ݦ<  �<`�<��<3ן<��<kC�<�u�<���<�Ӗ<���<*�<SR�<�x�<	��<���</�<c�<�%�<�D�<c�<���<�:}<�sy<��u<�q<�n<�Pj<��f<վb<h�^<�.[<�gW<4�S<��O<�L<�YH<b�D<B�@<r"=<Jj9<��5<�2<�S.<y�*<'<�]#<o�<	$<�<�<s<��<�n
<��<�< <�d�;��;6��;!b�;>��; [�;!��;��;�R�;v�;��;u�;���;��;�D�;<��;��;hQ�;<Պ;n�;l�;��u;�pk;�Ka;�OW;~M;��C;@S:;8�0;�';:�;#�;5;@u;���:@�:6��:��:槶:��:�l�:#�:�r:<XT:Y�6:W�:�~�9K��9޺�9��$9S>[8�KW��i!������ƺ�~���CA+�D�D�{(^��Xw��.����������D��@~����ź��Ѻ��ݺ���L���� �����������r�nN�l&$�s�)���/��5��d;��-A��F�)�L��|R��>X�= ^���c��i��@o� u���z��?���������Y���[�������0���h���K���0���  �  )|=�=t�=�c==��=�I=A� =r� =n- =4��<���<1�<�\�<���<���<��<DS�<���<���<d�<6<�<�s�<\��<���<��<�F�<x�<$��<���<��</�<�X�<Ȁ�<��<2��<P��<r�<h+�<�F�<L`�<w�<E��<���<{��<2��<��<���<���<��<k��<`��<���<��<h��<�s�<X�<8�<��<���<~��<e��<�T�<�<q��<���<eH�<���<6��<�J�<���<���<��<���<�=�<�ž<�H�<�ƻ<Q@�<0��<V%�<��<i��<s[�<S��<+�<l�<2��<��<�Z�<E��<�<�*�<�i�<<��<��<�<�K�<Q~�<���<�ܔ<I	�<�3�<�\�<g��<R��<ω<~�<��<Z6�<�V�<�v�<�+}<@iy<��u<��q<"n<sXj<�f<��b<�_<�H[<�W<��S<�P<�FL<�H<;�D<�A<~`=<�9<A�5<�N2<U�.<��*<�Z'<�#<�! <��<��<�n<n�<wg<��
<�w<�	<6� <���;���;�+�;F��;��;x��;N;�;y��;o��;�{�;�`�;zX�;�c�;K��;��;Z��;!Y�;ɑ;N�;��;���;��x;�_n; 7d;�7Z;y`P;)�F;`)=;0�3;I�*;v!;Q�;=�;9;��:�?�:���:Le�:*U�:=~�:��:z�:��z:d�\:/�>:D�!:��:pV�9�ӗ9��?9�a�8�Zⷲ���*t�YH��N
�.��&���?��iY�:�r�������������BV��z�����ú%к1ܺ�D�K��@" ����
����v��@��y�#��~)��V/�`+5�	�:���@�B�F��fL�11R�G�W�y�]���c�3Ni��o�,�t�ܞz��1����������ڈ� �������g����n��U���<���  �  *|=�=u�=�c==��=�I=1� =r� =n- =@��<��<1�<�\�<|��<���<��<SS�<��<���<\�<<�<�s�<S��<���<��<�F�<x�<$��<���<��</�<�X�<̀�<��<��<Z��<l�<e+�<G�<M`�<w�<J��<ɜ�<z��<;��<���<���<���<���<o��<Z��<���<���<o��<�s�<X�<8�<��<���<z��<j��<�T�<��<k��<��<kH�<���<B��<�J�<���<���<��<���<�=�<�ž<�H�<�ƻ<X@�<��<V%�<��<e��<s[�<]��<4�<!l�<7��<��<�Z�<&��<s�<�*�<�i�<H��<�ߝ<$�<�K�<S~�<���<�ܔ<U	�<�3�<�\�<F��<G��<�Ή<{�<��<Y6�<�V�<�v�<�+}<:iy<��u<��q<%n<�Xj<ϓf<��b<�_<qH[<�W<��S<�P<�FL<��H<=�D<�A<|`=<��9<8�5<�N2<S�.<��*<�Z'<��#<�! <��<��<�n<m�<�g<��
<�w<�	<�� <���;���;�+�;b��;��;���;K;�;e��;W��;�{�;�`�;�X�;�c�;;+��;C��;Y�;(ɑ;N�;n�;���;�x;�_n;G7d;�7Z;M`P;��F;(=;K�3;�*;lv!;��;u�;>;��:O@�:ٳ�:�e�:�T�:�~�:R��:�x�:ʌz:��\:��>:�!:G�:�X�9�җ9S�?9Dg�8�i�3��>&t�	M���-��&���?��jY���r�������������U��(���H�úbк3ܺ�E��J��C" �a��
�������.��_�#�~)�MV/��+5��:���@���F�gL�K1R���W���]�.�c�2Ni�o�C�t���z��1���������]ۈ����{�������gn��$U���<���  �  #|=�=k�=�c==��=�I=4� =|� =n- =?��<��<1�<�\�<~��<���<��<[S�<���<���<p�<<�<�s�<S��<���<��<�F�<x�<��<���<��</�<�X�<π�<��<��<^��<i�<Y+�<�F�<F`�<w�<<��<���<i��<@��<���<���<���<���<���<Y��<���<���<q��<�s�<X�<8�<��<���<y��<}��<�T�<��<|��<��<pH�<���<2��<xJ�<���<���<��<���<�=�<�ž<�H�<�ƻ<]@�<��<V%�<��<b��<i[�<I��< �<l�<;��<��<�Z�</��<��<�*�<�i�<S��<�ߝ<-�<�K�<_~�<���<�ܔ<W	�<�3�<�\�<L��<Z��<ω<|�<��<F6�<�V�<�v�<�+}<,iy<��u<��q<n<�Xj<��f<��b<�_<]H[<�W<��S<�P<�FL<߉H<�D<�A<�`=<��9<[�5<�N2<}�.<��*<�Z'<	�#<�! <Ƌ<��<�n<k�<�g<��
<x<�	<� <���;���;�+�;E��;��;a��;,;�;k��;A��;�{�;q`�;�X�;�c�;���;>��;7��;�X�;ɑ;�M�;e�;y��;��x;9_n;u7d;�7Z;�`P;=�F;�(=;��3;�*;�v!;k�;��;i;&�:t@�:���:�f�:�T�:��:@�:�y�:�z:h�\:��>:��!:M�:}T�9�З91�?9B^�8������#t�CO��r乂,��&���?��kY���r�o���.���V����V��ޤ���ú-кs2ܺzD�'J��T" ���g��t�����P�#��})�>V/��+5�Z�:���@��F��fL�@1R���W��]���c��Ni�o�y�t���z�2����������ۈ�������������nn��@U���<���  �  $|=�=w�=�c==��=�I=9� =v� =w- =N��<��<;�<�\�<���<���<��<aS�<��<���<h�<)<�<�s�<S��<���<��<�F�<x�<��<���<��</�<�X�<���<ަ�<��<;��<e�<Q+�<�F�<<`�<w�<<��<Ü�<|��<9��<��<���<���<���<x��<n��<���< ��<y��<�s�<.X�<&8�<��<���<���<s��<�T�< �<g��<���<hH�<���<=��<yJ�<���<���<��<���<�=�<vž<�H�<�ƻ<>@�<��<E%�<��<X��<l[�<O��<2�<l�<7��<��<�Z�<8��<��<�*�<�i�<W��<��<2�<�K�<i~�<���<�ܔ<e	�<4�<�\�<V��<R��<�Ή<��<��<]6�<�V�<�v�<�+}<iy<��u<��q<n<UXj<Ɠf<b�b<}_<\H[<��W<��S<�P<�FL<�H<F�D<�A<�`=<�9<A�5<�N2<e�.<��*<�Z'<�#<�! <Ӌ<��<�n<��<�g<��
<x<�	<� <���;���;�+�;T��;��;z��;>;�;I��;9��;\{�;�`�;;X�;�c�;ڂ�;���;,��;�X�;�ȑ;�M�;g�;z��;Ѱx;�_n;=7d;�7Z;B`P;,�F;)=;��3;Ì*;�v!;��;Ǹ;�;w�: A�:���:g�:$V�:,�:B�:z�:y�z:B�\:��>:>�!:׿:U�9�ї9��?9jX�8������6t��N��q�A0�}&���?��kY��r�6�������2���JV�������ú^к�1ܺ�D� J���! ����
�?�����|���#��})��U/��*5���:���@�D�F�5gL�1R��W�b�]�o�c��Ni�6o���t��z�2����"���mۈ�Z���ƣ�������n��WU��=���  �  !|=�=q�=�c=	=�=�I=B� =v� =}- =P��<��<L�<�\�<���<���<��<fS�<
��<���<k�<8<�<�s�<b��<���<��<�F�<x�<��<���<��<�.�<�X�<���<Φ�<��</��<_�<A+�<�F�<1`�<�v�<4��<���<u��<1��<��<���<��<��<|��<y��<���<��<���<�s�<2X�<08�<��<���<���<y��<�T�<�<o��<���<bH�<���<-��<oJ�<���<���<��<���<�=�<kž<�H�<�ƻ<4@�<��<3%�<��<D��<a[�<@��<!�<l�<6��<��<�Z�<G��<��<�*�<�i�<Y��<��<:�<L�<l~�<Į�<
ݔ<d	�<4�<�\�<e��<]��<	ω<��<��<S6�<�V�<�v�<�+}<iy<��u<n�q<�n<1Xj<��f<=�b<w_<@H[<�W<��S<�P<�FL<ʉH</�D<�A<�`=<�9<Y�5<�N2<e�.<��*<�Z'<2�#<�! <�<�<o<��<�g<��
<)x<�	<?� <ׂ�;��;�+�;>��;��;>��;;�;���;?��;){�;S`�;X�;�c�;���;���;��;�X�;�ȑ;�M�;#�;]��;i�x;�_n;7d;O8Z;�`P;��F;V)=;��3;�*; w!;q�;2�;;��:�A�:ϵ�:g�:�V�:��:��:�z�:��z:��\:�>:G�!:�:�R�90Η9,�?9�Y�8��ⷨ��N;t�DQ����F1�� &���?��kY�k�r���������&����V��	����ú�к�0ܺ�D躘I��i! ���
�������f����#�H})��U/��*5���:��@��F��fL��0R�S�W���]��c��Ni��o���t�E�z�V2����i����ۈ�����ң��舑��n��VU��K=���  �  |=�=n�=�c==��=�I=A� =�� =|- =Y��<3��<X�<�\�<���<���<�<�S�<	��<���<��<5<�<�s�<P��<���<��<�F�<x�<��<���<��<�.�<�X�<���<���<���<2��<D�<7+�<�F�<+`�<�v�<4��<���<k��<C��<���<���<��<��<���<v��<���<��<���<t�<GX�<@8�<��<��<���<���<�T�<�<v��<��<rH�<���</��<pJ�<���<���<��<���<i=�<lž<kH�<�ƻ<-@�<<2%�<ꐵ<@��<][�<C��<�<l�<;��<��<�Z�<B��<��<�*�<�i�<t��<'��<O�<L�<�~�<Ϯ�<ݔ<s	�<4�<
]�<d��<a��<�Ή<|�<��<K6�<�V�<�v�<�+}<�hy<w�u<A�q<�n<1Xj<}�f<6�b<G_<H[<ׅW<��S<�P<uFL<ӉH<"�D<�A<�`=<��9<g�5<�N2<��.<��*<['<]�#<�! <�<�<;o<��<�g<��
<8x<�	<;� <��;���;�+�;P��;��;[��;;�; ��;��;*{�;�_�;�W�;Oc�;F��;���;���;jX�;�ȑ;�M�;�;a��;��x;Y_n;�7d;�7Z;�`P;��F;l)=;��3;�*;�w!;Æ;��;�;�:�B�:N��:�h�:�V�:
��:8�:�z�:��z:=�\::�>:;�!:A�::S�9�͗9��?9rJ�8�����9t��X����	2��$&���?�`nY���r�����\���O����V������:�ú&к1ܺEC��H���! ����	�J�������0�#��|)�_U/��*5���:��@�ȚF�!gL�@1R���W���]���c��Ni��o�-�t���z��2��x��g����ۈ�����0���R����n���U��L=���  �  |=�=k�=�c==��=�I=?� =�� =- ={��<A��<]�<�\�<���<���<�<�S�<%��<���<��<1<�<�s�<V��<���<��<�F�<x�<���<���<~�< /�<�X�<���<���<���<��<*�<>+�<�F�<`�<�v�<��<���<`��<O��<���<���<��<��<���<��<ݮ�<"��<���<t�<RX�<S8�<��</��<���<���<�T�<�<���<��<H�<���</��<\J�<���<���<�<���<O=�<Už<_H�<�ƻ<@�<ܴ�<5%�<ϐ�<;��<B[�<:��<�<l�<J��<��<�Z�<?��<��<�*�<j�<���<'��<e�<L�<�~�<֮�<%ݔ<�	�<4�<]�<c��<m��<ω<��<��<C6�<�V�<�v�<�+}<�hy<a�u<P�q<�n<Xj<Y�f<�b<_<H[<˅W<|�S<�P<CFL<։H<�D<�A<�`=<	�9<��5<�N2<��.<��*<H['<z�#<�! <C�<,�<lo<��<*h<�
<Ix<�	<5� <R��;���;1,�;?��;��;T��;�:�;���;���;:{�;�_�;�W�;.c�;��;L��;L��;�X�;jȑ;XM�;��;��;��x;_n;8d;�7Z;$aP;бF;�)=;��3;W�*;�x!;ކ;�;V;��:�C�:���:�j�:�W�:r��:��:�z�:��z:`�\:�>:�!:n�:�N�9�ȗ9��?930�8�����dDt�p[����=5��&&�R�?��qY�9�r����҅��r���+W������(�ú5кH1ܺ�B�kH���  ���	������������#�u|)�AT/�u*5�h�:��@�h�F��fL�1R���W�4�]���c��Oi�o���t��z��2���������D܈�࿋�����H���o���U��_=���  �  |=�=f�=�c==�=�I=L� =�� =�- =}��<A��<u�<�\�<Û�<���<�<�S�<3��<���<��<G<�<�s�<_��<���<��<�F�<�w�<���<���<y�<�.�<�X�<���<���<���<	��<)�< +�<�F�<`�<�v�<!��<���<`��<?��<��<���<��<"��<���<���<خ�<4��<���<t�<[X�<i8�<��<'��<���<���<�T�<�<���<���<oH�<���<��<YJ�<x��<���<n�<g��<K=�<@ž<TH�<�ƻ<@�<״�<%�<Ɛ�<5��<<[�<.��<
�<l�<>��<��<�Z�<R��<��<�*�<%j�<���<?��<w�<'L�<�~�<ﮖ<-ݔ<�	�<(4�<]�<~��<o��<ω<��<��<;6�<�V�<�v�<�+}<�hy<%�u<$�q<�n<�Wj<E�f<��b<_<�G[<��W<o�S<�P<LFL<��H< �D<�A<�`=<�9<��5<�N2<��.<"�*<N['<{�#<!" <[�<P�<�o<��<h<=�
<rx<
<d� <J��; ��;,�;0��;T�;+��;�:�;���;���;�z�;�_�;wW�;�b�;���;���;M��;X�;ȑ;AM�;��;��;-�x;_n;�7d;8Z;)aP;&�F;l*=;��3;0�*;�x!;x�;�;�;x�:QE�:��:�j�:0Y�:Ł�:	�:�{�:7�z:��\:4�>:�!:��:7N�9
Ǘ9��?9��8�t�M���Nt��]����6�&'&���?�}rY���r����}���a���oW��[�����úMк�/ܺ5B�pG��,  �S�����Y�����'�#�5|)�MT/��)5�\�:�B�@�W�F��fL��0R��W�r�]� �c��Oi�9o��t�۠z��2���������k܈�?������������o��	V��~=���  �  |=�=n�=�c==�=�I=O� =�� =�- =���<^��<��<]�<ޛ�<���<9�<�S�<>��<���<��<K<�<�s�<h��<���<��<�F�<�w�<���<k��<{�<�.�<�X�<v��<���<���<���< �<+�<�F�<	`�<�v�<%��<���<r��<6��<
��<���<��<$��<���<���<֮�<R��<���<1t�<wX�<g8�<�<'��<˽�<���<�T�<�<��<���<_H�<���<��<\J�<l��<t��<q�<K��<B=�<-ž<>H�<uƻ<�?�<ʴ�<�$�<ǐ�<��<:[�<.��<�<l�<+��<��<�Z�<R��<��<�*�<2j�<���<Z��<s�<EL�<�~�<���<Iݔ<�	�<>4�<]�<���<i��<ω<��<��<N6�<�V�<�v�<Z+}<�hy<!�u<��q<zn<�Wj<1�f<��b<�
_<�G[<}�W<p�S<nP<NFL<��H<"�D<�A<�`=<!�9<u�5<	O2<��.<E�*<Y['<��#<L" <g�<��<�o<3�<Dh<U�
<�x<
<n� <8��;I��;�+�;z��;z�;&��;�:�;e��;���;qz�;j_�;OW�;�b�;���;���;,��;�W�;/ȑ;
M�;��;1��;ϯx;�_n;E7d;K8Z;>aP;�F;�*=;$�3;َ*;�x!;h�;�;R;H�:FE�:���:�j�:DZ�:��:4�:�{�:�z:|�\:P�>:M�!:M�:ZO�9Pė9ô?9�$�8����<Wt��b��9$�a8��(&�u�?�DrY���r����o���3���GV��w�����ú�к�/ܺ B��F��� ����%��b��L����#�N{)�?T/�)5�h�:�,�@���F�lfL�1R��W���]�w�c�vOi�o�,�t��z�Q3����[����܈�����Ԥ��㉑��o��V���=���  �  |=�=f�=�c==�=�I=R� =�� =�- =���<l��<��<]�<��<���<;�<�S�<C��<���<��<P<�<�s�<q��<���<��<}F�<�w�<��<i��<q�<�.�<tX�<g��<���<���<���<�<+�<�F�< `�<�v�<��<���<f��<7��<��<���< ��<.��<���<���<��<\��<ŋ�<=t�<�X�<p8�<�<;��<ɽ�<���<�T�< �<���< ��<cH�<���<��<NJ�<e��<k��<d�<I��<,=�<!ž<7H�<qƻ<�?�<���<�$�<���<��<.[�<"��<��<l�<3��<��<�Z�<Y��<��<�*�<3j�<���<_��<��<ML�<�~�<��<Wݔ<�	�<<4�<(]�<���<y��<#ω<��<��<>6�<�V�<�v�<T+}<�hy<�u<��q<Un<�Wj<�f<��b<�
_<�G[<v�W<U�S<lP<+FL<��H<�D<�A<�`=<;�9<��5<O2<�.<B�*<p['<Ҽ#<U" <��<��<�o<8�<ch<`�
<�x<:
<{� <w��;s��;,�;S��;N�;���;�:�;c��;i��;yz�;%_�;W�;zb�;���;���;���;�W�;ȑ;�L�;��;���;��x;H_n;W7d;r8Z;�aP;w�F;�*=;��3;Ў*;My!;��;I�;�;�:�E�:M��:�k�:0Z�:��:��:h|�:*�z:\�\:��>: �!:T�:L�9�9��?9��8���j��X\t��d���$�:�C+&�[�?��sY�N�r������������V����c�ú�кv/ܺ�@�iF��� �f������&��ʿ���#��z)��S/�)5���:���@��F� fL��0R�0�W�^�]���c��Oi�.o���t�
�z�h3��]��|����܈������������o��<V���=���  �  |=�=h�=�c== �=�I=Q� =�� =�- =���<i��<��<*]�<ڛ�<��<D�<�S�<O��<���<��<P<�<�s�<[��<���<��<�F�<�w�<��<v��<Z�<�.�<mX�<^��<{��<���<���<��<�*�<�F�<`�<�v�<��<���<c��<;��<��<���<��<*��<���<���<���<Y��<��<Gt�<�X�<�8�<�<F��<ͽ�<���<�T�<�<���<��<hH�<���<��<IJ�<f��<s��<P�<B��<=�<ž<"H�<`ƻ<�?�<���<�$�<���<��<&[�<$��<�<l�<8��<��<�Z�<X��<��<�*�<;j�<���<c��<��<AL�<�~�<��<Tݔ<�	�<@4�<1]�<���<t��<ω<��<��<?6�<�V�<�v�<f+}<�hy<�u<��q<?n<�Wj<�f<��b<�
_<�G[<U�W<7�S<�P<FL<��H<�D<�A<�`=<�9<��5<O2<��.<N�*<�['<μ#<v" <��<��<�o<K�<mh<y�
<�x<C
<|� <f��;��;,�;@��;}�;��;e:�;���;��;Gz�;_�;�V�;Lb�;R��;|��;���;�W�;�Ǒ;�L�;��;ڔ�;=�x;4_n;{7d;8Z;6aP;C�F;�*=;��3;�*;�y!;��;P�;;�:+H�:7��:�l�:rZ�:���:��:(|�:S�z:E�\:��>:F�!:�:K�92×9�?9��88�����"`t�|i���(�;�b,&���?�@vY���r���ꆒ�����VW��������ú)кt/ܺ�@��E��q �4���������A��Ӟ#��z)�HS/��(5�y�:���@�1�F��fL��0R�6�W�X�]�<�c�RPi��o���t���z��3���������݈�����A���*����o��wV���=���  �  |=�=g�=�c=	=	�=�I=W� =�� =�- =���<s��<��<(]�<��<
��<K�<�S�<R��<���<��<`<�<�s�<m��<���<��<�F�<�w�<ڧ�<`��<\�<�.�<lX�<\��<p��<���<���<�<�*�<�F�<�_�<�v�<��<���<^��<6��<��<���<.��<4��<���<���<���<`��<��<It�<�X�<�8�<!�<K��<ֽ�<���<�T�<.�<���< ��<bH�<���<��<8J�<V��<`��<P�<7��< =�<ž<H�<Xƻ<�?�<���<�$�<���<��<[�<��< �<�k�<3��<��<�Z�<g��<��<�*�<Aj�<���<h��<��<QL�<�~�<��<[ݔ<�	�<G4�<0]�<���<���< ω<��<��<?6�<�V�<{v�<?+}<�hy<��u<��q<Bn<�Wj<�f<��b<�
_<�G[<W�W<3�S<ZP<	FL<��H<�D<�A<�`=<0�9<��5<)O2<�.<\�*<�['<�#<~" <��<��<�o<Y�<�h<��
<�x<E
<�� <���;h��;,�;=��;_�;ϝ�;M:�;E��;��;=z�;_�;�V�;$b�;>��;_��;���;nW�;�Ǒ;�L�;K�;���;��x;_n;T7d;�8Z;�aP;�F;+=;�3;)�*;�y!;�;(�;;z�:�G�:���:�l�:[�:
��:L�:Q}�:}�z:t�\:��>:��!:��:�F�92��9��?9X�8�%����bt��j���*�\;�,&���?�vY�g�r����1�������yW��ͤ����ú\к�.ܺ�@�oE��A �����������A��֞#��z)�ES/��(5���:���@���F�fL��0R�Q�W�W�]�ˉc��Pi��o���t���z��3���������݈����>���C����o��~V��>���  �  |=�=i�=�c==�=�I=W� =�� =�- =���<��<��<$]�<��<���<K�<�S�<H��< ��<��<_<�<�s�<o��<���<��<�F�<�w�<���<_��<b�<�.�<]X�<W��<p��<���<���<�<�*�<�F�<�_�<�v�< ��<���<j��<0��<��<���<$��<3��<���<���<���<p��<׋�<St�<�X�<�8�<.�<O��<Խ�<���<�T�<$�<���< ��<]H�<���<��<PJ�<h��<Z��<T�<,��<=�<ž<H�<Wƻ<�?�<���<�$�<���<��<<[�< ��<�<l�<*��<��<�Z�<d��<��<�*�<7j�<���<l��<��<kL�<�~�<��<jݔ<�	�<J4�<4]�<���<y��<ω<��<��<E6�<�V�<�v�<I+}<�hy<�u<��q<An<yWj<��f<}�b<�
_<uG[<E�W<1�S<_P<IFL<��H<�D<�A<�`=<-�9<��5<*O2<��.<a�*<�['<��#<v" <��<��<�o<Z�<�h<n�
<�x<O
<�� <d��;o��;�+�;Q��;u�;��;�:�;B��;3��;z�;�^�;�V�;"b�;L��;J��;���;<W�;�Ǒ;�L�;��;$��;̯x;r_n;&7d;~8Z;|aP;��F;+=;,�3;L�*;�y!;c�;ܻ;k;y�:6G�:W��:m�:�Z�:���:e�:�|�:�z:h�\:G�>:L�!:`�:�L�9�×9��?9�	�8"O�t��Ret�;j���*�2<�L-&���?�ZuY���r�������v����V��c�����ú0к�.ܺr@�dE��� ���s���-��H����#�Ez)�lS/��(5�[�:���@��F�<fL��0R�d�W�!�]���c��Oi�Yo��t���z��3��������� ݈����?���x���p���V��>���  �  |=�=g�=�c=	=	�=�I=W� =�� =�- =���<s��<��<(]�<��<
��<K�<�S�<R��<���<��<`<�<�s�<m��<���<��<�F�<�w�<ڧ�<`��<\�<�.�<lX�<\��<p��<���<���<�<�*�<�F�<�_�<�v�<��<���<^��<6��<��<���<.��<4��<���<���<���<`��<��<It�<�X�<�8�<!�<K��<ֽ�<���<�T�<.�<���< ��<bH�<���<��<8J�<V��<`��<P�<7��< =�<ž<H�<Xƻ<�?�<���<�$�<���<��<[�<��< �<�k�<3��<��<�Z�<g��<��<�*�<Aj�<���<h��<��<QL�<�~�<��<[ݔ<�	�<G4�<0]�<���<���< ω<��<��<?6�<�V�<{v�<?+}<�hy<��u<��q<Bn<�Wj<�f<��b<�
_<�G[<W�W<3�S<ZP<	FL<��H<�D<�A<�`=<0�9<��5<)O2<�.<\�*<�['<�#<~" <��<��<�o<Y�<�h<��
<�x<E
<�� <���;h��;,�;=��;_�;ϝ�;M:�;E��;��;=z�;_�;�V�;$b�;>��;_��;���;nW�;�Ǒ;�L�;K�;���;��x;_n;S7d;�8Z;�aP;�F;+=;�3;)�*;�y!;�;(�;;z�:�G�:���:�l�:[�:
��:L�:Q}�:}�z:t�\:��>:��!:��:�F�92��9��?9X�8�%����bt��j���*�\;�,&���?�vY�g�r����1�������yW��ͤ����ú\к�.ܺ�@�oE��A �����������A��֞#��z)�ES/��(5���:���@���F�fL��0R�Q�W�W�]�ˉc��Pi��o���t���z��3���������݈����>���C����o��~V��>���  �  |=�=h�=�c== �=�I=Q� =�� =�- =���<i��<��<*]�<ڛ�<��<D�<�S�<O��<���<��<P<�<�s�<[��<���<��<�F�<�w�<��<v��<Z�<�.�<mX�<^��<{��<���<���<��<�*�<�F�<`�<�v�<��<���<c��<;��<��<���<��<*��<���<���<���<Y��<��<Gt�<�X�<�8�<�<F��<ͽ�<���<�T�<�<���<��<hH�<���<��<IJ�<f��<s��<P�<B��<=�<ž<"H�<`ƻ<�?�<���<�$�<���<��<&[�<$��<�<l�<8��<��<�Z�<X��<��<�*�<;j�<���<c��<��<AL�<�~�<��<Tݔ<�	�<@4�<1]�<���<t��<ω<��<��<?6�<�V�<�v�<f+}<�hy<�u<��q<?n<�Wj<�f<��b<�
_<�G[<U�W<7�S<�P<FL<��H<�D<�A<�`=<�9<��5<O2<��.<N�*<�['<μ#<v" <��<��<�o<K�<mh<y�
<�x<C
<|� <f��;��;,�;@��;}�;��;e:�;���;��;Gz�;_�;�V�;Lb�;R��;|��;���;�W�;�Ǒ;�L�;��;ڔ�;=�x;4_n;{7d;8Z;6aP;B�F;�*=;��3;�*;�y!;��;P�;;�:+H�:7��:�l�:rZ�:���:��:(|�:S�z:E�\:��>:F�!:�:K�92×9�?9��88�����"`t�|i���(�;�b,&���?�@vY���r���ꆒ�����VW��������ú)кt/ܺ�@��E��q �4���������A��Ӟ#��z)�HS/��(5�y�:���@�1�F��fL��0R�6�W�X�]�<�c�RPi��o���t���z��3���������݈�����A���*����o��wV���=���  �  |=�=f�=�c==�=�I=R� =�� =�- =���<l��<��<]�<��<���<;�<�S�<C��<���<��<P<�<�s�<q��<���<��<}F�<�w�<��<i��<q�<�.�<tX�<g��<���<���<���<�<+�<�F�< `�<�v�<��<���<f��<7��<��<���< ��<.��<���<���<��<\��<ŋ�<=t�<�X�<p8�<�<;��<ɽ�<���<�T�< �<���< ��<cH�<���<��<NJ�<e��<k��<d�<I��<,=�<!ž<7H�<qƻ<�?�<���<�$�<���<��<.[�<"��<��<l�<3��<��<�Z�<Y��<��<�*�<3j�<���<_��<��<ML�<�~�<��<Wݔ<�	�<<4�<(]�<���<y��<#ω<��<��<>6�<�V�<�v�<T+}<�hy<�u<��q<Un<�Wj<�f<��b<�
_<�G[<v�W<U�S<lP<+FL<��H<�D<�A<�`=<;�9<��5<O2<�.<B�*<p['<Ҽ#<U" <��<��<�o<8�<ch<`�
<�x<:
<{� <w��;s��;,�;S��;N�;���;�:�;c��;i��;yz�;%_�;W�;zb�;���;���;���;�W�;ȑ;�L�;��;���;��x;H_n;W7d;r8Z;�aP;w�F;�*=;��3;Ў*;My!;��;I�;�;�:�E�:M��:�k�:0Z�:��:��:h|�:*�z:\�\:��>: �!:T�:L�9�9��?9��8���j��X\t��d���$�:�C+&�[�?��sY�N�r������������V����c�ú�кv/ܺ�@�iF��� �f������&��ʿ���#��z)��S/�)5���:���@��F� fL��0R�0�W�^�]���c��Oi�.o���t�
�z�h3��]��|����܈������������o��<V���=���  �  |=�=n�=�c==�=�I=O� =�� =�- =���<^��<��<]�<ޛ�<���<9�<�S�<>��<���<��<K<�<�s�<h��<���<��<�F�<�w�<���<k��<{�<�.�<�X�<v��<���<���<���< �<+�<�F�<	`�<�v�<%��<���<r��<6��<
��<���<��<$��<���<���<֮�<R��<���<1t�<wX�<g8�<�<'��<˽�<���<�T�<�<��<���<_H�<���<��<\J�<l��<t��<q�<K��<B=�<-ž<>H�<uƻ<�?�<ʴ�<�$�<ǐ�<��<:[�<.��<�<l�<+��<��<�Z�<R��<��<�*�<2j�<���<Z��<s�<EL�<�~�<���<Iݔ<�	�<>4�<]�<���<i��<ω<��<��<N6�<�V�<�v�<Z+}<�hy<!�u<��q<zn<�Wj<1�f<��b<�
_<�G[<}�W<p�S<nP<NFL<��H<"�D<�A<�`=<!�9<u�5<	O2<��.<E�*<Y['<��#<L" <g�<��<�o<3�<Dh<U�
<�x<
<n� <8��;I��;�+�;z��;z�;&��;�:�;e��;���;qz�;j_�;OW�;�b�;���;���;,��;�W�;/ȑ;
M�;��;1��;ϯx;�_n;E7d;K8Z;>aP;�F;�*=;$�3;َ*;�x!;h�;�;R;H�:FE�:���:�j�:DZ�:��:4�:�{�:�z:|�\:P�>:M�!:M�:ZO�9Pė9ô?9�$�8����<Wt��b��9$�a8��(&�u�?�DrY���r����o���3���GV��w�����ú�к�/ܺ B��F��� ����%��b��L����#�N{)�?T/�)5�h�:�,�@���F�lfL�1R��W���]�w�c�vOi�o�,�t��z�Q3����[����܈�����Ԥ��㉑��o��V���=���  �  |=�=f�=�c==�=�I=L� =�� =�- =}��<A��<u�<�\�<Û�<���<�<�S�<3��<���<��<G<�<�s�<_��<���<��<�F�<�w�<���<���<y�<�.�<�X�<���<���<���<	��<)�< +�<�F�<`�<�v�<!��<���<`��<?��<��<���<��<"��<���<���<خ�<4��<���<t�<[X�<i8�<��<'��<���<���<�T�<�<���<���<oH�<���<��<YJ�<x��<���<n�<g��<K=�<@ž<TH�<�ƻ<@�<״�<%�<Ɛ�<5��<<[�<.��<
�<l�<>��<��<�Z�<R��<��<�*�<%j�<���<?��<w�<'L�<�~�<ﮖ<-ݔ<�	�<(4�<]�<~��<o��<ω<��<��<;6�<�V�<�v�<�+}<�hy<%�u<$�q<�n<�Wj<E�f<��b<_<�G[<��W<o�S<�P<LFL<��H< �D<�A<�`=<�9<��5<�N2<��.<"�*<N['<{�#<!" <[�<P�<�o<��<h<=�
<rx<
<d� <J��;��;,�;/��;T�;+��;�:�;���;���;�z�;�_�;wW�;�b�;���;���;M��;X�;ȑ;AM�;��;��;-�x;_n;�7d;8Z;)aP;&�F;l*=;��3;0�*;�x!;x�;�;�;x�:QE�:��:�j�:0Y�:Ł�:	�:�{�:7�z:��\:4�>:�!:��:7N�9
Ǘ9��?9��8�t�M���Nt��]����6�&'&���?�}rY���r����}���a���oW��[�����úMк�/ܺ5B�pG��,  �S�����Y�����'�#�5|)�MT/��)5�\�:�B�@�W�F��fL��0R��W�r�]� �c��Oi�9o��t�۠z��2���������k܈�?������������o��	V��~=���  �  |=�=k�=�c==��=�I=?� =�� =- ={��<A��<]�<�\�<���<���<�<�S�<%��<���<��<1<�<�s�<V��<���<��<�F�<x�<���<���<~�< /�<�X�<���<���<���<��<*�<>+�<�F�<`�<�v�<��<���<`��<O��<���<���<��<��<���<��<ݮ�<"��<���<t�<RX�<S8�<��</��<���<���<�T�<�<���<��<H�<���</��<\J�<���<���<�<���<O=�<Už<_H�<�ƻ<@�<ܴ�<5%�<ϐ�<;��<B[�<:��<�<l�<J��<��<�Z�<?��<��<�*�<j�<���<'��<e�<L�<�~�<֮�<%ݔ<�	�<4�<]�<c��<m��<ω<��<��<C6�<�V�<�v�<�+}<�hy<a�u<P�q<�n<Xj<Y�f<�b<_<H[<˅W<|�S<�P<CFL<։H<�D<�A<�`=<	�9<��5<�N2<��.<��*<H['<z�#<�! <C�<,�<lo<��<*h<�
<Ix<�	<5� <R��;���;1,�;?��;��;T��;�:�;���;���;:{�;�_�;�W�;.c�;��;L��;L��;�X�;jȑ;XM�;��;��;��x;_n;8d;�7Z;$aP;бF;�)=;��3;W�*;�x!;ކ;�;V;��:�C�:���:�j�:�W�:r��:��:�z�:��z:`�\:�>:�!:n�:�N�9�ȗ9��?930�8�����dDt�p[����=5��&&�R�?��qY�9�r����҅��r���+W������(�ú5кH1ܺ�B�kH���  ���	������������#�u|)�AT/�u*5�h�:��@�h�F��fL�1R���W�4�]���c��Oi�o���t��z��2���������D܈�࿋�����H���o���U��_=���  �  |=�=n�=�c==��=�I=A� =�� =|- =Y��<3��<X�<�\�<���<���<�<�S�<	��<���<��<5<�<�s�<P��<���<��<�F�<x�<��<���<��<�.�<�X�<���<���<���<2��<D�<7+�<�F�<+`�<�v�<4��<���<k��<C��<���<���<��<��<���<v��<���<��<���<t�<GX�<@8�<��<��<���<���<�T�<�<v��<��<rH�<���</��<pJ�<���<���<��<���<i=�<lž<kH�<�ƻ<-@�<<2%�<ꐵ<@��<][�<C��<�<l�<;��<��<�Z�<B��<��<�*�<�i�<t��<'��<O�<L�<�~�<Ϯ�<ݔ<s	�<4�<
]�<d��<a��<�Ή<|�<��<K6�<�V�<�v�<�+}<�hy<w�u<A�q<�n<1Xj<}�f<6�b<G_<H[<ׅW<��S<�P<uFL<ӉH<"�D<�A<�`=<��9<g�5<�N2<��.<��*<['<]�#<�! <�<�<;o<��<�g<��
<8x<�	<;� <��;���;�+�;P��;��;[��;;�; ��;��;*{�;�_�;�W�;Oc�;F��;���;���;jX�;�ȑ;�M�;�;a��;��x;Y_n;�7d;�7Z;�`P;��F;l)=;��3;�*;�w!;Æ;��;�;�:�B�:N��:�h�:�V�:
��:8�:�z�:��z:=�\::�>:;�!:A�::S�9�͗9��?9rJ�8�����9t��X����	2��$&���?�`nY���r�����\���O����V������:�ú&к1ܺEC��H���! ����	�J�������0�#��|)�_U/��*5���:��@�ȚF�!gL�@1R���W���]���c��Ni��o�-�t���z��2��x��g����ۈ�����0���R����n���U��L=���  �  !|=�=q�=�c=	=�=�I=B� =v� =}- =P��<��<L�<�\�<���<���<��<fS�<
��<���<k�<8<�<�s�<b��<���<��<�F�<x�<��<���<��<�.�<�X�<���<Φ�<��</��<_�<A+�<�F�<1`�<�v�<4��<���<u��<1��<��<���<��<��<|��<y��<���<��<���<�s�<2X�<08�<��<���<���<y��<�T�<�<o��<���<bH�<���<-��<oJ�<���<���<��<���<�=�<kž<�H�<�ƻ<4@�<��<3%�<��<D��<a[�<@��<!�<l�<6��<��<�Z�<G��<��<�*�<�i�<Y��<��<:�<L�<l~�<Į�<
ݔ<d	�<4�<�\�<e��<]��<	ω<��<��<S6�<�V�<�v�<�+}<iy<��u<n�q<�n<1Xj<��f<=�b<w_<@H[<�W<��S<�P<�FL<ʉH</�D<�A<�`=<�9<Y�5<�N2<e�.<��*<�Z'<2�#<�! <�<�<o<��<�g<��
<)x<�	<?� <ׂ�;��;�+�;>��;��;>��;;�;���;?��;){�;S`�;X�;�c�;���;���;��;�X�;�ȑ;�M�;#�;]��;i�x;�_n;7d;O8Z;�`P;��F;V)=;��3;�*; w!;q�;2�;;��:�A�:ϵ�:g�:�V�:��:��:�z�:��z:��\:�>:G�!:�:�R�90Η9,�?9�Y�8��ⷨ��N;t�DQ����F1�� &���?��kY�k�r���������&����V��	����ú�к�0ܺ�D躘I��i! ���
�������f����#�H})��U/��*5���:��@��F��fL��0R�S�W���]��c��Ni��o���t�E�z�V2����i����ۈ�����ң��舑��n��VU��K=���  �  $|=�=w�=�c==��=�I=9� =v� =w- =N��<��<;�<�\�<���<���<��<aS�<��<���<h�<)<�<�s�<S��<���<��<�F�<x�<��<���<��</�<�X�<���<ަ�<��<;��<e�<Q+�<�F�<<`�<w�<<��<Ü�<|��<9��<��<���<���<���<x��<n��<���< ��<y��<�s�<.X�<&8�<��<���<���<s��<�T�< �<g��<���<hH�<���<=��<yJ�<���<���<��<���<�=�<vž<�H�<�ƻ<>@�<��<E%�<��<X��<l[�<O��<2�<l�<7��<��<�Z�<8��<��<�*�<�i�<W��<��<2�<�K�<i~�<���<�ܔ<e	�<4�<�\�<V��<R��<�Ή<��<��<]6�<�V�<�v�<�+}<iy<��u<��q<n<UXj<Ɠf<b�b<}_<\H[<��W<��S<�P<�FL<�H<F�D<�A<�`=<�9<A�5<�N2<e�.<��*<�Z'<�#<�! <Ӌ<��<�n<��<�g<��
<x<�	<� <���;���;�+�;T��;��;z��;>;�;I��;9��;\{�;�`�;;X�;�c�;ڂ�;���;,��;�X�;�ȑ;�M�;g�;z��;Ѱx;�_n;=7d;�7Z;B`P;,�F;)=;��3;Ì*;�v!;��;Ǹ;�;w�: A�:���:g�:$V�:,�:B�:z�:y�z:B�\:��>:>�!:׿:U�9�ї9��?9jX�8������6t��N��q�A0�}&���?��kY��r�6�������2���JV�������ú^к�1ܺ�D� J���! ����
�?�����|���#��})��U/��*5���:���@�D�F�5gL�1R��W�b�]�o�c��Ni�6o���t��z�2����"���mۈ�Z���ƣ�������n��WU��=���  �  #|=�=k�=�c==��=�I=4� =|� =n- =?��<��<1�<�\�<~��<���<��<[S�<���<���<p�<<�<�s�<S��<���<��<�F�<x�<��<���<��</�<�X�<π�<��<��<^��<i�<Y+�<�F�<F`�<w�<<��<���<i��<@��<���<���<���<���<���<Y��<���<���<q��<�s�<X�<8�<��<���<y��<}��<�T�<��<|��<��<pH�<���<2��<xJ�<���<���<��<���<�=�<�ž<�H�<�ƻ<]@�<��<V%�<��<b��<i[�<I��< �<l�<;��<��<�Z�</��<��<�*�<�i�<S��<�ߝ<-�<�K�<_~�<���<�ܔ<W	�<�3�<�\�<L��<Z��<ω<|�<��<F6�<�V�<�v�<�+}<,iy<��u<��q<n<�Xj<��f<��b<�_<]H[<�W<��S<�P<�FL<߉H<�D<�A<�`=<��9<[�5<�N2<}�.<��*<�Z'<	�#<�! <Ƌ<��<�n<k�<�g<��
<x<�	<� <���;���;�+�;E��;��;a��;,;�;k��;A��;�{�;q`�;�X�;�c�;���;>��;7��;�X�;ɑ;�M�;e�;y��;��x;9_n;u7d;�7Z;�`P;=�F;�(=;��3;�*;�v!;k�;��;i;&�:t@�:���:�f�:�T�:��:@�:�y�:�z:h�\:��>:��!:M�:}T�9�З91�?9B^�8������#t�CO��r乂,��&���?��kY���r�o���.���V����V��ޤ���ú-кs2ܺzD�'J��T" ���g��t�����P�#��})�>V/��+5�Z�:���@��F��fL�@1R���W��]���c��Ni�o�y�t���z�2����������ۈ�������������nn��@U���<���  �  *|=�=u�=�c==��=�I=1� =r� =n- =@��<��<1�<�\�<|��<���<��<SS�<��<���<\�<<�<�s�<S��<���<��<�F�<x�<$��<���<��</�<�X�<̀�<��<��<Z��<l�<e+�<G�<M`�<w�<J��<ɜ�<z��<;��<���<���<���<���<o��<Z��<���<���<o��<�s�<X�<8�<��<���<z��<j��<�T�<��<k��<��<kH�<���<B��<�J�<���<���<��<���<�=�<�ž<�H�<�ƻ<X@�<��<V%�<��<e��<s[�<]��<4�<!l�<7��<��<�Z�<&��<s�<�*�<�i�<H��<�ߝ<$�<�K�<S~�<���<�ܔ<U	�<�3�<�\�<F��<G��<�Ή<{�<��<Y6�<�V�<�v�<�+}<:iy<��u<��q<%n<�Xj<ϓf<��b<�_<qH[<�W<��S<�P<�FL<��H<=�D<�A<|`=<��9<8�5<�N2<S�.<��*<�Z'<��#<�! <��<��<�n<m�<�g<��
<�w<�	<�� <���;���;�+�;b��;��;���;K;�;e��;W��;�{�;�`�;�X�;�c�;;+��;C��;Y�;(ɑ;N�;n�;���;�x;�_n;G7d;�7Z;M`P;��F;(=;K�3;�*;lv!;��;u�;>;��:O@�:ٳ�:�e�:�T�:�~�:R��:�x�:ʌz:��\:��>:�!:G�:�X�9�җ9S�?9Dg�8�i�3��>&t�	M���-��&���?��jY���r�������������U��(���H�úbк3ܺ�E��J��C" �a��
�������.��_�#�~)�MV/��+5��:���@���F�gL�K1R���W���]�.�c�2Ni�o�C�t���z��1���������]ۈ����{�������gn��$U���<���  �  Vz=�=�=�`=�=[�=�E=�� =�� =E( =��<	��<[�<�N�<��<���<f�<�A�<}|�<(��<���<{&�<�\�<n��<���<���<+�<M[�<��<_��<��<�<p5�<�[�<���<`��<��<���< ��<�<�0�<�E�<�X�<Zh�<�u�<��<ц�<Ȋ�<���<��<ۂ�<Wy�<�k�< [�<�E�<-�<�<���<E��<B��<�p�<�=�<4�<���<���<�B�<���<��<>S�<���<��<=7�<���<a�<��<iw�<d��<�z�<.��<7k�<�ܶ<�I�<���<\�<�w�<oԮ<@-�<7��<�ө<�!�<.l�<v��<���<79�<�w�<���<��<�#�<�X�<��<���<�<��<B�<�k�<ړ�<º�<k��<��<�(�<RK�<km�<�}<F_y<�u<H�q<* n<�_j<��f<t�b<�_<a[<�W<4�S<�*P<|pL<�H<�E<�MA<ƛ=<��9<J@6<�2<�.<�N+<y�'<$<� <t�<�a<)�<$X<j�<�d<�<��<&<n��;B��;_J�;��;?�;���;�t�;�(�;���;���;���;﫵;>��;�ݩ;��;�]�;G��;-�;ﲍ;�L�;��;	z{;�'q;��f;��\;lS;%gI;8�?;)o6;v,-;1$; ;�:;��	;f� ; �:�\�:���:�ɿ:ׯ:��:���:�L�:@bd:)�F:4):��:�@�9N�9��Y9���8�y�(B�%[]��I���nٹ���1!�(!;��T�Khn� 䃺�������z���ݵ�".º�pκۢں��溯�����$t�Em��b�NQ��<��##�H)���.���4���:��q@��EF��L�`�Q���W���]�Rc�>i���n�p�t��~z��$��?
��$���2ֈ�����㋑��t���]���H���  �  Uz=�=�=�`=�=U�=�E=�� =�� =?( =��<��<X�<�N�<݌�<���<^�<�A�<t|�<"��<���<z&�<�\�<e��<���<���<!+�<][�<��<[��<��<!�<w5�<�[�<���<\��<��<���<��<�<�0�<�E�<�X�<ph�<�u�<��<Ȇ�<���<���<���<��<My�<�k�<�Z�<�E�<
-�<�<���<:��<C��<�p�<�=�<D�<���<���<�B�<���<��<US�<���<ߚ�<>7�<���<a�<��<qw�<^��<�z�<4��<>k�<�ܶ<�I�<���<V�<�w�<�Ԯ<B-�<=��<�ө<�!�<-l�<���<���<,9�<�w�<���<��<�#�<�X�<	��<���<�<��<B�<�k�<ٓ�<���<k��<�<�(�<fK�<em�<w}<:_y<�u<X�q<! n<�_j<x�f<��b<�_<a[<�W<#�S<{*P<vpL<,�H<�E<�MA<ɛ=<��9<F@6<%�2<A�.<�N+<p�'<$<� <r�<�a<=�<X<l�<�d<�<ǉ<&<g��; ��;xJ�;��;Q?�;���;�t�;�(�;a��;���;���;���;b��;�ݩ;�;�]�;���;'-�;鲍;�L�;��;�z{;�'q;�f;��\;/S;gI;��?;�o6;-,-;4$;�;6;;C�	;
� ;� �:�[�:��:ɿ:�ׯ:��:���:IL�:�`d:b�F:>):w�:�A�9-L�9�Y9	��8��v�>�BW]��J��Mnٹ���0!�T;��T�zhn�䃺�~��M��xz��]ݵ��.ºqκ�ںf�����b���t��m�Fb��Q��<��##��)���.��4���:�zq@��EF�)L�]�Q�:�W���]�uQc�gi���n���t�i~z��$��R
�����^ֈ�Ѽ�����͋��st���]���H���  �  Sz=�=�=�`=�=X�=�E=�� =�� =>( =��<��<^�<O�<ߌ�<��<]�<�A�<|�< ��<���<p&�<	]�<g��<���<���<+�<T[�<��<h��<��<�<a5�<�[�<���<V��<��<���<��<�<�0�<�E�<�X�<ph�<vu�<��<ǆ�<Ί�<���<��<��<Ny�<l�<�Z�<F�<-�<�<���<7��<[��<�p�<�=�<>�<���<È�<�B�<���<��<RS�<���<��<A7�<���<a�<��<hw�<X��<�z�<(��<&k�<�ܶ<�I�<���<U�<�w�<}Ԯ<:-�<F��<�ө<�!�<$l�<���<���<39�<�w�<���<�<�#�<�X�<��<���<*�<��<B�<�k�<䓋<���<n��<
�<�(�<fK�<am�<�}<._y<
�u<E�q<�n<�_j<n�f<��b<�_<�`[<�W<�S<�*P<ppL<&�H<�E<�MA<ԛ=<��9<^@6<�2<O�.<�N+<��'<$<� <��<�a<j�<X<��<�d<�<щ<
&<���;+��;�J�;��;6?�;���;�t�;�(�;2��;���;d��;���;]��;�ݩ;��;t]�;j��;�,�;貍;�L�;���;�z{;$'q;j�f;��\;�S;,gI;`�?;�o6;1,-;�$;�;�;;{�	;)� ;%�:�[�:���:@ɿ:�ׯ:��:w��:7M�:�`d:ЉF:�):�:�?�9�L�9�Y9w��8��w��S�7[]�SL���oٹK��3!��;���T��fn��䃺�������z���ܵ��.ºpκy�ںW����������s��m��a��Q��<�H##��)�l�.��4�̚:��q@��EF��L�G�Q��W�/�]�vQc��i���n�ѳt��~z��$���
�����rֈ�˼��_��� ����t��&^���H���  �  Rz=�=�=�`=�=W�=�E=�� =�� =D( =��<��<a�<O�<��<��<f�<�A�<�|�<*��<���<|&�<]�<c��<���<���<+�<Q[�<��<S��<��<�<g5�<�[�<���<W��<	��<���<��<�<�0�<�E�<�X�<dh�<~u�<��<���<ʊ�<���<���<��<Ry�<l�<�Z�<F�<-�<�<���<@��<R��<�p�<�=�<C�<���<���<�B�<���<��<IS�<���<���<17�<���<a�<��<`w�<V��<�z�<)��<-k�<�ܶ<�I�<���<S�<�w�<{Ԯ<=-�<=��<�ө<�!�<-l�<���<���<69�<�w�<���<��<�#�<�X�<��<���<(�<��<B�<�k�<���<���<c��<�<�(�<[K�<`m�<v}<_y<��u<G�q< n<�_j<u�f<c�b<�_<�`[<�W<�S<q*P<lpL<�H<�E<�MA<��=<��9<Z@6</�2<O�.<�N+<��'<$<� <��<�a<Z�<&X<~�<�d<�<ω<"&<���;��;wJ�;��;C?�;���;�t�;�(�;3��;���;|��;֫�;��;�ݩ;��;�]�;c��;�,�;���;�L�;���;dz{;h'q;#�f;\�\;zS;(gI;��?;�o6;T,-;�$;�;�;;φ	;�� ;��:S\�:	��:wɿ:=د:��:���:M�:�_d:^�F:�):*�:�?�9�L�9Y�Y9��8�-x�pI��^]��L���rٹ��2!�� ;���T��in��䃺������z��Rݵ�+/º&pκڢںU��=������s�Ym��a�KQ�r<�G##�c)�u�.���4�ؚ:�Xq@��EF��L���Q�J�W���]��Qc��i���n��t��~z��$��q
��D���cֈ����<���󋑻�t��<^���H���  �  Tz=�=�=�`=�=[�=�E=�� =�� =I( =!��<"��<w�<O�<���<��<��<�A�<�|�<2��<���<�&�<]�<q��<���<~��<+�<N[�<��<H��<��<�<Z5�<�[�<���<Q��<���<���<���<�<�0�<�E�<�X�<]h�<}u�<��<φ�<Њ�<���<��<��<by�<l�<[�<F�<-�<�<���<^��<U��<�p�<�=�<N�<���<È�<�B�<���<��<AS�<���<ٚ�<)7�<���<�`�<��<Mw�<O��<�z�<��<!k�<�ܶ<�I�<���<Q�<�w�<tԮ<9-�<;��<�ө<�!�<7l�<���<���<C9�<�w�<ó�<��<�#�<�X�<&��<���<(�<��<B�<�k�<ᓋ<ƺ�<p��<��<�(�<VK�<em�<a}<_y<�u<�q<�n<�_j<o�f<8�b<�_<�`[<٢W<�S<Y*P<rpL<�H<�E<�MA<ϛ=<��9<U@6<G�2<D�.<O+<��'<C$<?� <��<b<`�<bX<��<�d<+�<щ<8&<���;V��;J�;���;6?�;���;�t�;p(�;Y��;{��;J��;���;⺯;�ݩ;��;x]�;뺘;�,�;���;�L�;���;/z{;g'q;��f;��\;�S;ngI;�?;�o6;�,-;�$;�;�;;��	;�� ;!�:?^�:A��:ʿ:�د:��:V��:FM�:�ad:��F:x):=�:�>�9K�9��Y9���8��{�mS�h]�N���tٹ�*4!��";���T�kn��䃺���)���z��gݵ�9.º[pκ?�ں���������\s�^l��a��P�K<��"#��)�{�.�[�4��:��p@��EF��L�:�Q���W��]��Qc�ni�S�n��t�z�'%���
������nֈ�e���g���J����t��+^���H���  �  Mz=�=�=�`=�=[�=�E=�� =�� =R( =3��<��<u�<O�<��<$��<u�<�A�<�|�<?��<���<�&�<]�<o��<���<���<+�<@[�<��<N��<���<��<Q5�<�[�<���<<��<���<���<���<��<�0�<�E�<vX�<bh�<yu�<��<Ɇ�<ӊ�<���<��<���<sy�<l�<[�<F�<.-�<&�<���<O��<^��<q�<�=�<N�<���<ǈ�<�B�<���<��<GS�<��<Ӛ�<"7�<���<�`�<��<Hw�<;��<zz�<��<k�<�ܶ<�I�<���<I�<�w�<wԮ<9-�<<��<�ө<�!�<2l�<���<���<P9�<�w�<���<�<$�<�X�<'��<���<7�<�<&B�<�k�<�<Ⱥ�<n��<�<�(�<SK�<Tm�<b}<�^y<؟u<�q<�n<�_j<?�f<6�b<�_<�`[<ȢW<��S<a*P<UpL<��H<�E<�MA<ϛ=<��9<q@6<7�2<`�.<4O+<��'<<$<;� <��<.b<��<GX<��<�d<F�<�<1&<Β�;S��;�J�;��;:?�;]��;�t�;�(�;���;`��;+��;���;ں�;\ݩ;{�;f]�;�;�,�;���;�L�;���;[z{;J'q;/�f;��\;�S;�gI;��?;Sp6;c--; $;�;X<;o�	;@� ;T�:_]�:���:o˿:$ٯ:��:i��:�M�:"ad:��F:):�:;�9�I�9��Y9���8� |�&\��i]�S���vٹ��>5!�K#;���T�ejn�,僺̀������z��Dݵ�V.º�oκz�ں_��@�����Ns��l�$a�nP��;��"#��)���.���4�|�:�2q@�GEF��L�J�Q�H�W��]�Rc��i�K�n���t�cz�'%���
�������ֈ�h���q���W����t���^���H���  �  Ez=�=�=�`=�=\�=�E=�� =�� =M( ==��<0��<��<'O�< ��<8��<��<B�<�|�<=��<���<�&�<]�<j��<���<z��<+�<G[�<���<F��<���<��<C5�<�[�<y��<*��<���<y��<���<��<�0�<�E�<oX�<fh�<mu�<��<ņ�<ڊ�<���<��<	��<fy�<,l�<[�<4F�<6-�<)�<���<]��<q��<�p�<�=�<Z�<���<Ј�<�B�<���<���<HS�<|��<Ϛ�<7�<t��<�`�<y�<Ew�<(��<iz�<
��<k�<�ܶ<�I�<���<;�<�w�<vԮ<.-�<<��<�ө<�!�<3l�<���<���<O9�<�w�<���<%�<$�<�X�<:��<���<F�<�<6B�<�k�<���<̺�<l��<��<�(�<YK�<Fm�<_}<�^y<Ɵu<��q<�n<_j<�f<%�b<�_<�`[<��W<��S<[*P<6pL<�H<�E<�MA<˛=<��9<~@6<9�2<��.<"O+<˰'<b$<^� <��< b<��<iX<��<e<C�<�<5&<��;A��;�J�;��;5?�;}��;Dt�;s(�;���;S��;���;o��;���;ݩ;t�;]�;޺�;�,�;^��;�L�;���;�z{;�&q;#�f;��\;S;�gI;9�?;�p6;--;�$;;=;��	;[� ;��:=^�:��:�ʿ:�ٯ:� �:���:/N�:D`d:d�F:a):Z�:V:�9I�94�Y9���8��|�Qr⸸j]�UW���zٹ��7!��#;���T��kn��僺r�������{��7ݵ��.ºoκ`�ںb��������r�dl�z`��P�H;�	"#�9)���.�&�4���:�#q@�(EF��L�\�Q�c�W�Z�]��Qc�di�Y�n���t��z�[%���
������3׈�������������u���^���H���  �  Dz=�=�=�`=�=_�=�E=�� =�� =T( =C��<?��<��<1O�<��<=��<��<B�<�|�<G��<���<�&�<]�<s��<���<}��<+�<D[�<���<8��<���<��<05�<�[�<i��<-��<���<i��<���<��<�0�<�E�<mX�<]h�<uu�<��<ц�<ڊ�<���<��<��<uy�<1l�<,[�<8F�<F-�<9�<���<q��<u��<q�<>�<_�<���<Έ�<�B�<���<��<>S�<x��<���<7�<x��<�`�<k�</w�<&��<]z�<���<�j�<ܶ<�I�<���<2�<�w�<nԮ<0-�<>��<�ө<�!�<<l�<���<���<X9�<�w�<׳�<(�<$�<�X�<F��<���<I�<�<=B�<�k�<쓋<Ϻ�<t��<��<�(�<RK�<Em�<=}<�^y<��u<��q<�n<Y_j<�f<�b<p_<�`[<��W<��S<5*P<3pL<��H<�E<�MA<؛=<��9<p@6<[�2<��.<<O+<ְ'<�$<� <��<Pb<��<�X<��<e<[�<�<R&<ߒ�;m��;�J�;��;(?�;w��;8t�;<(�;���;��;���;��;o��;)ݩ;�;�\�;���;�,�;M��;dL�;���;=z{;0'q; �f;��\;S;�gI;��?;�p6;--;�$;�;+=;:�	;�� ;��:�_�:[��:�˿:Mگ:� �:���:N�:bd:��F:V):1�:�9�9xE�9�Y9���8M�~�y�ku]��W���}ٹ3�]9!�P&;�+�T��ln�u惺����R��V{��
ݵ�.ºYoκ��ںK��o��~���br��k�[`��O��:��!#��)�l�.���4�Ǚ:��p@�cEF�wL��Q�c�W�A�]�Rc�hi���n�ִt��z��%��<���׈�ͽ������ތ��4u���^��8I���  �  Hz=�=�=�`=�=`�=�E=�� =�� =`( =K��<D��<��<2O�</��<>��<��<B�<�|�<X��<���<�&�<]�<z��<���<���<+�<6[�< ��<+��<���<��<85�<�[�<Z��< ��<���<z��<���<��<�0�<�E�<oX�<Rh�<wu�<��<І�<Ԋ�<���<��<��<�y�<4l�<3[�<=F�<Q-�<J�<���<z��<v��<q�<	>�<c�<���<ƈ�<�B�<���<��<6S�<w��<���<7�<i��<�`�<y�<w�<��<Mz�<���<�j�<rܶ<�I�<}��<6�<�w�<lԮ<5-�<5��<�ө<�!�<Ml�<���<��<f9�<�w�<۳�<)�<+$�<�X�<J��<û�<R�</�<7B�<�k�<���<к�<n��<��<�(�<DK�<Jm�<!}<�^y<��u<��q<�n<._j<�f<��b<x_<�`[<��W<��S<*P<BpL<�H<�E<�MA<̛=<��9<�@6<w�2<��.<oO+<�'<�$<�� <��<�b<��<�X<��<,e<~�<�<u&<��;���;�J�;��;#?�;A��;Yt�;(�;���;���;Ѯ�;��;8��;�ܩ;��;]�;}��;a,�;*��;?L�;���;�y{;H'q;�f;��\;�S;.hI;��?;�p6;?.-;$;�;X=;��	;n� ;�:(`�:���:$Ϳ:�گ:"!�:���:�M�:Rbd:ǇF:�):S�:�9�9�D�9�Y9F��8E��ep⸇]�:[���ٹZ�8!��';�a�T�\nn�惺P���n���z���ݵ��-º�oκ��ں*�溠�����kr��k�O`�NO��:��!#��)�$�.�տ4���:�2p@�EF�mL�I�Q�p�W�5�]��Rc�Ci�N�n�F�t�R�z��%����[�>׈����礎�Ќ��}u���^��oI���  �  Cz=�=�=�`=�=c�=�E=�� =Ň =]( =V��<W��<��<GO�<2��<U��<��<+B�<�|�<Y��<��<�&�<]�<y��<���<r��<+�<3[�<��<+��<���<��<5�<�[�<U��<��<���<Z��<���<��<�0�<�E�<fX�<Th�<hu�<��<ӆ�<ۊ�<���<��<��<�y�<Il�<?[�<NF�<W-�<O�<��<���<���<q�<>�<g�<��<͈�<�B�<���<���<4S�<l��<���<�6�<Y��<�`�<X�<w�<��<Gz�<���<�j�<uܶ<�I�<x��<)�<�w�<cԮ<$-�<;��<�ө<�!�<Ll�<���<��<j9�<x�<糝<?�<0$�<�X�<W��<ӻ�<^�<&�<BB�<�k�<���<պ�<u��<��<�(�<IK�<Am�<&}<�^y<��u<��q<�n<*_j<�f<��b<I_<e`[<y�W<��S<#*P<+pL<�H<�E<~MA<ڛ=<��9<�@6<p�2<��.<bO+<��'<�$<�� <&�<�b<��<�X<�<<e<��<,�<q&<��;���;�J�;ܼ�;?�;;��;,t�;(�;v��;���;n��;Ӫ�;%��;�ܩ;��;�\�;N��;*,�;��;.L�;���;�y{;�&q;#�f;�\;S;jhI;��?;7q6;.-;�$;2;�=;ˈ	;�� ;'�:�`�:.��:�̿:ۯ:w!�:��:!N�:ybd:Q�F:�
):�:$7�9>B�9g�Y9���8�Y�����3�]��]��U�ٹ
��;!�\';�T�T��nn��惺��������{��ݵ��-º!oκ��ں��溄��J���vq�)k��_�&O�N:� !#�)���.��4���:�Pp@��DF�IL��Q���W���]�_Rc��i�;�n���t���z��%����a񅻂׈�&���E�������u�� _��ZI���  �  <z=�=�=�`=�=^�=�E=�� =͇ =_( =c��<S��<��<YO�<0��<a��<��<+B�<�|�<b��<
��<�&�<$]�<p��<���<}��<+�<7[�<��<,��<���<��<5�<�[�<O��<��<���<Q��<���<��<�0�<�E�<]X�<Vh�<mu�<��<Ά�<݊�<���< ��<.��<�y�<Ul�<6[�<NF�<a-�<S�<��<y��<���<q�<">�<i�<��<ӈ�<�B�<���<���<5S�<f��<���<�6�<T��<�`�<P�<w�<���<=z�<���<�j�<wܶ<�I�<x��< �<�w�<gԮ<,-�<C��<�ө<�!�<Jl�<���<��<k9�<x�<ڳ�<I�<0$�<�X�<P��<ͻ�<m�<'�<VB�<�k�<��<Ϻ�<u��<�<�(�<JK�<3m�<'}<�^y<��u<��q<yn<8_j<ɞf<��b<?_<h`[<}�W<��S<#*P<pL<�H<�E<�MA<ߛ=<��9<�@6<u�2<��.<lO+<�'<�$<�� <J�<�b<�<�X<�<He<��<>�<q&</��;g��;�J�;��;?�;I��;t�;(�;Q��;���;V��;ڪ�;��;�ܩ;��;|\�;q��;,�;���;'L�;]��;z{;'q;j�f;��\;7S;\hI;��?;�q6;.-;$;�;�=;�	;�� ;u�:)`�:���:�̿:"ܯ:�!�:���:�N�:�ad:��F:�):\�:�5�91A�9(�Y9���8��4���}]��`����ٹ���<!��&;��T��nn�i烺�������k{���ܵ�N.ºinκĠںn�����.���kq��k�R_�'O��9�W!#�=)�P�.��4���:�>p@��DF�sL��Q�9�W�w�]�TRc��i�6�n��t���z��%�����F񅻷׈����X�������u��2_��[I���  �  @z=�=޾=�`=�=e�=�E=�� =Ǉ =e( =e��<b��<��<WO�<5��<b��<��<3B�<�|�<g��< ��<�&�<#]�<~��<���<|��<+�<.[�<��<(��<���<��<5�<�[�<D��<��<���<T��<���<��<�0�<�E�<eX�<Fh�<mu�<��<؆�<��<���< ��<#��<�y�<Yl�<M[�<XF�<g-�<Y�<��<���<���<#q�<>�<g�<
��<ֈ�<�B�<���<���<&S�<j��<���<�6�<Q��<�`�<Q�<w�<���<4z�<���<�j�<_ܶ<�I�<t��<&�<�w�<ZԮ<--�<:��<�ө<�!�<Pl�<���<��<w9�<x�<<N�<5$�<�X�<a��<໔<p�<3�<IB�<�k�<	��<ٺ�<y��<��<�(�<<K�<>m�<}<�^y<q�u<��q<wn<_j<ƞf<��b<6_<T`[<a�W<��S<*P<!pL<ѷH<�E<�MA<ݛ=<��9<�@6<z�2<��.<�O+<�'<�$<�� <G�<�b<�<�X<.�<Ze<��<+�<|&<.��;���;�J�;��;�>�;)��;#t�;(�;Z��;���;a��;���;幯;�ܩ;��;�\�;+��;,�;���;.L�;~��;�y{;'q;�f;@�\;eS;�hI;��?;�q6;w.-;5$;�;5>;N�	;�� ;��:�a�:���:�Ϳ:�ۯ:z!�:n��:�N�:3cd:K�F:�):t�:�6�9{B�9w�Y9���8�7�����0�]�la��͆ٹw�A<!��);���T�8on�烺灐�e��]{��"ݵ�i-ºonκi�ں��溡��i���7q��j�&_�O��9�� #��)�2�.���4�`�:�(p@��DF�(L���Q�r�W���]��Rc��i�]�n�εt���z�	&������񅻼׈�f���j���<����u��%_��vI���  �  ?z=�=�=�`=�=c�=�E=�� =ʇ =i( =T��<]��<��<NO�<>��<]��<��<*B�<�|�<k��<��<�&�<]�<���<���<{��<
+�</[�<��<��<���<��<#5�<�[�<J��<��<���<^��<���<��<�0�<�E�<fX�<Jh�<zu�<��<Ն�<͊�<���<'��<#��<�y�<Cl�<G[�<QF�<i-�<_�<��<���<���<&q�<>�<n�<��<���<�B�<���<
��<-S�<k��<���<�6�<]��<�`�<\�<�v�<��<>z�<���<�j�<_ܶ<�I�<a��<�<�w�<bԮ<1-�<0��<�ө<�!�<Sl�<���<��<s9�< x�<�<I�<:$�<�X�<`��<ڻ�<Z�<=�<NB�<�k�<���<κ�<w��<��<�(�<<K�<>m�<�}<�^y<��u<��q<�n<�^j<�f<��b<?_<V`[<m�W<��S<�)P<pL<ַH<�E<�MA<֛=<��9<|@6<��2<��.<�O+<��'<�$<�� <5�<�b<�<�X<�<Je<��<:�<�&<ܒ�;���;�J�;��;?�;-��;t�;�'�;~��;���;���;���; ��;�ܩ;_�;�\�;!��;4,�;���;�K�;���;�y{;k'q;��f;,�\;�S;ShI;�?;�q6;�.-;�$;{;�=;`�	;� ;��:La�:���:�Ϳ:�ۯ:�!�: ��:[M�:	cd:!�F:r):o�:D7�9�=�9"�Y9���8�S�����w�]�0^��y�ٹ���:!��);���T��qn��烺́�����{���ݵ�G-º�oκ4�ںL��w������q��j�M_��N�:�� #��)���.�`�4�9�:��o@�EF�|L� �Q���W�E�]��Rc��i��n���t���z�&�������}׈�n���W���7����u���^���I���  �  @z=�=޾=�`=�=e�=�E=�� =Ǉ =e( =e��<b��<��<WO�<5��<b��<��<3B�<�|�<g��< ��<�&�<#]�<~��<���<|��<+�<.[�<��<(��<���<��<5�<�[�<D��<��<���<T��<���<��<�0�<�E�<eX�<Fh�<mu�<��<؆�<��<���< ��<#��<�y�<Yl�<M[�<XF�<g-�<Y�<��<���<���<#q�<>�<g�<
��<ֈ�<�B�<���<���<&S�<j��<���<�6�<Q��<�`�<Q�<w�<���<4z�<���<�j�<_ܶ<�I�<t��<&�<�w�<ZԮ<--�<:��<�ө<�!�<Pl�<���<��<w9�<x�<<N�<5$�<�X�<a��<໔<p�<3�<IB�<�k�<	��<ٺ�<y��<��<�(�<<K�<>m�<}<�^y<q�u<��q<wn<_j<ƞf<��b<6_<T`[<a�W<��S<*P<!pL<ѷH<�E<�MA<ݛ=<��9<�@6<z�2<��.<�O+<�'<�$<�� <G�<�b<�<�X<.�<Ze<��<+�<|&<.��;���;�J�;��;�>�;)��;#t�;(�;Z��;���;a��;���;幯;�ܩ;��;�\�;+��;,�;���;.L�;~��;�y{;'q;�f;@�\;eS;�hI;��?;�q6;w.-;5$;�;5>;N�	;�� ;��:�a�:���:�Ϳ:�ۯ:z!�:n��:�N�:3cd:K�F:�):t�:�6�9{B�9w�Y9���8�7�����0�]�la��͆ٹw�A<!��);���T�8on�烺灐�e��]{��"ݵ�i-ºonκi�ں��溡��i���7q��j�&_�O��9�� #��)�2�.���4�`�:�(p@��DF�(L���Q�r�W���]��Rc��i�]�n�εt���z�	&������񅻼׈�f���j���<����u��%_��vI���  �  <z=�=�=�`=�=^�=�E=�� =͇ =_( =c��<S��<��<YO�<0��<a��<��<+B�<�|�<b��<
��<�&�<$]�<p��<���<}��<+�<7[�<��<,��<���<��<5�<�[�<O��<��<���<Q��<���<��<�0�<�E�<]X�<Vh�<mu�<��<Ά�<݊�<���< ��<.��<�y�<Ul�<6[�<NF�<a-�<S�<��<y��<���<q�<">�<i�<��<ӈ�<�B�<���<���<5S�<f��<���<�6�<T��<�`�<P�<w�<���<=z�<���<�j�<wܶ<�I�<x��< �<�w�<gԮ<,-�<C��<�ө<�!�<Jl�<���<��<k9�<x�<ڳ�<I�<0$�<�X�<P��<ͻ�<m�<'�<VB�<�k�<��<Ϻ�<u��<�<�(�<JK�<3m�<'}<�^y<��u<��q<yn<8_j<ɞf<��b<?_<h`[<}�W<��S<#*P<pL<�H<�E<�MA<ߛ=<��9<�@6<u�2<��.<lO+<�'<�$<�� <J�<�b<�<�X<�<He<��<>�<q&</��;g��;�J�;��;?�;I��;t�;(�;P��;���;V��;ڪ�;��;�ܩ;��;|\�;q��;,�;���;'L�;]��;z{;'q;j�f;��\;7S;\hI;��?;�q6;.-;$;�;�=;�	;�� ;u�:)`�:���:�̿:"ܯ:�!�:���:�N�:�ad:��F:�):\�:�5�91A�9(�Y9���8��4���}]��`����ٹ���<!��&;��T��nn�i烺�������k{���ܵ�N.ºinκĠںn�����.���kq��k�R_�'O��9�W!#�=)�P�.��4���:�>p@��DF�sL��Q�9�W�w�]�TRc��i�6�n��t���z��%�����F񅻷׈����X�������u��2_��[I���  �  Cz=�=�=�`=�=c�=�E=�� =Ň =]( =V��<W��<��<GO�<2��<U��<��<+B�<�|�<Y��<��<�&�<]�<y��<���<r��<+�<3[�<��<+��<���<��<5�<�[�<U��<��<���<Z��<���<��<�0�<�E�<fX�<Th�<hu�<��<ӆ�<ۊ�<���<��<��<�y�<Il�<?[�<NF�<W-�<O�<��<���<���<q�<>�<g�<��<͈�<�B�<���<���<4S�<l��<���<�6�<Y��<�`�<X�<w�<��<Gz�<���<�j�<uܶ<�I�<x��<)�<�w�<cԮ<$-�<;��<�ө<�!�<Ll�<���<��<j9�<x�<糝<?�<0$�<�X�<W��<ӻ�<^�<&�<BB�<�k�<���<պ�<u��<��<�(�<IK�<Am�<&}<�^y<��u<��q<�n<*_j<�f<��b<I_<e`[<y�W<��S<#*P<+pL<�H<�E<~MA<ڛ=<��9<�@6<p�2<��.<bO+<��'<�$<�� <&�<�b<��<�X<�<<e<��<,�<q&<��;���;�J�;ܼ�;?�;;��;,t�;(�;v��;���;n��;Ӫ�;%��;�ܩ;��;�\�;N��;*,�;��;.L�;���;�y{;�&q;#�f;�\;S;jhI;��?;7q6;.-;�$;2;�=;ˈ	;�� ;'�:�`�:.��:�̿:ۯ:w!�:��:!N�:ybd:Q�F:�
):�:$7�9>B�9g�Y9���8�Y�����3�]��]��U�ٹ
��;!�\';�T�T��nn��惺��������{��ݵ��-º!oκ��ں��溄��J���vq�)k��_�&O�N:� !#�)���.��4���:�Pp@��DF�IL��Q���W���]�_Rc��i�;�n���t���z��%����a񅻂׈�&���E�������u�� _��ZI���  �  Hz=�=�=�`=�=`�=�E=�� =�� =`( =K��<D��<��<2O�</��<>��<��<B�<�|�<X��<���<�&�<]�<z��<���<���<+�<6[�< ��<+��<���<��<85�<�[�<Z��< ��<���<z��<���<��<�0�<�E�<oX�<Rh�<wu�<��<І�<Ԋ�<���<��<��<�y�<4l�<3[�<=F�<Q-�<J�<���<z��<v��<q�<	>�<c�<���<ƈ�<�B�<���<��<6S�<w��<���<7�<i��<�`�<y�<w�<��<Mz�<���<�j�<rܶ<�I�<}��<6�<�w�<lԮ<5-�<5��<�ө<�!�<Ml�<���<��<f9�<�w�<۳�<)�<+$�<�X�<J��<û�<R�</�<7B�<�k�<���<к�<n��<��<�(�<DK�<Jm�<!}<�^y<��u<��q<�n<._j<�f<��b<x_<�`[<��W<��S<*P<BpL<�H<�E<�MA<̛=<��9<�@6<w�2<��.<oO+<�'<�$<�� <��<�b<��<�X<��<,e<~�<�<u&<��;���;�J�;��;#?�;A��;Yt�;(�;���;���;Ѯ�;��;8��;�ܩ;��;]�;}��;a,�;*��;?L�;���;�y{;H'q;�f;��\;�S;.hI;��?;�p6;?.-;$;�;X=;��	;n� ;�:(`�:���:$Ϳ:�گ:"!�:���:�M�:Rbd:ǇF:�):S�:�9�9�D�9�Y9F��8E��ep⸇]�:[���ٹZ�8!��';�a�T�\nn�惺P���n���z���ݵ��-º�oκ��ں*�溠�����kr��k�O`�NO��:��!#��)�$�.�տ4���:�2p@�EF�mL�I�Q�p�W�5�]��Rc�Ci�N�n�F�t�R�z��%����[�>׈����礎�Ќ��}u���^��oI���  �  Dz=�=�=�`=�=_�=�E=�� =�� =T( =C��<?��<��<1O�<��<=��<��<B�<�|�<G��<���<�&�<]�<s��<���<}��<+�<D[�<���<8��<���<��<05�<�[�<i��<-��<���<i��<���<��<�0�<�E�<mX�<]h�<uu�<��<ц�<ڊ�<���<��<��<uy�<1l�<,[�<8F�<F-�<9�<���<q��<u��<q�<>�<_�<���<Έ�<�B�<���<��<>S�<x��<���<7�<x��<�`�<k�</w�<&��<]z�<���<�j�<ܶ<�I�<���<2�<�w�<nԮ<0-�<>��<�ө<�!�<<l�<���<���<X9�<�w�<׳�<(�<$�<�X�<F��<���<I�<�<=B�<�k�<쓋<Ϻ�<t��<��<�(�<RK�<Em�<=}<�^y<��u<��q<�n<Y_j<�f<�b<p_<�`[<��W<��S<5*P<3pL<��H<�E<�MA<؛=<��9<p@6<[�2<��.<<O+<ְ'<�$<� <��<Pb<��<�X<��<e<[�<�<R&<ߒ�;m��;�J�;��;(?�;w��;8t�;<(�;���;��;���;��;o��;)ݩ;�;�\�;���;�,�;M��;dL�;���;=z{;0'q; �f;��\;S;�gI;��?;�p6;--;�$;�;+=;:�	;�� ;��:�_�:[��:�˿:Mگ:� �:���:N�:bd:��F:V):1�:�9�9xE�9�Y9���8M�~�y�ku]��W���}ٹ3�]9!�P&;�+�T��ln�u惺����R��V{��
ݵ�.ºYoκ��ںK��o��~���br��k�[`��O��:��!#��)�l�.���4�Ǚ:��p@�cEF�wL��Q�c�W�A�]�Rc�hi���n�ִt��z��%��<���׈�ͽ������ތ��4u���^��8I���  �  Ez=�=�=�`=�=\�=�E=�� =�� =M( ==��<0��<��<'O�< ��<8��<��<B�<�|�<=��<���<�&�<]�<j��<���<z��<+�<G[�<���<F��<���<��<C5�<�[�<y��<*��<���<y��<���<��<�0�<�E�<oX�<fh�<mu�<��<ņ�<ڊ�<���<��<	��<fy�<,l�<[�<4F�<6-�<)�<���<]��<q��<�p�<�=�<Z�<���<Ј�<�B�<���<���<HS�<|��<Ϛ�<7�<t��<�`�<y�<Ew�<(��<iz�<
��<k�<�ܶ<�I�<���<;�<�w�<vԮ<.-�<<��<�ө<�!�<3l�<���<���<O9�<�w�<���<%�<$�<�X�<:��<���<F�<�<6B�<�k�<���<̺�<l��<��<�(�<YK�<Fm�<_}<�^y<Ɵu<��q<�n<_j<�f<%�b<�_<�`[<��W<��S<[*P<6pL<�H<�E<�MA<˛=<��9<~@6<9�2<��.<"O+<˰'<b$<^� <��< b<��<iX<��<e<C�<�<5&<��;A��;�J�;��;5?�;}��;Dt�;s(�;���;S��;���;o��;���;ݩ;t�;]�;޺�;�,�;^��;�L�;���;�z{;�&q;#�f;��\;S;�gI;9�?;�p6;--;�$;;=;��	;[� ;��:=^�:��:�ʿ:�ٯ:� �:���:/N�:D`d:d�F:a):Z�:V:�9I�94�Y9���8��|�Qr⸸j]�UW���zٹ��7!��#;���T��kn��僺r�������{��7ݵ��.ºoκ`�ںb��������r�dl�z`��P�H;�	"#�9)���.�&�4���:�#q@�(EF��L�\�Q�c�W�Z�]��Qc�di�Y�n���t��z�[%���
������3׈�������������u���^���H���  �  Mz=�=�=�`=�=[�=�E=�� =�� =R( =3��<��<u�<O�<��<$��<u�<�A�<�|�<?��<���<�&�<]�<o��<���<���<+�<@[�<��<N��<���<��<Q5�<�[�<���<<��<���<���<���<��<�0�<�E�<vX�<bh�<yu�<��<Ɇ�<ӊ�<���<��<���<sy�<l�<[�<F�<.-�<&�<���<O��<^��<q�<�=�<N�<���<ǈ�<�B�<���<��<GS�<��<Ӛ�<"7�<���<�`�<��<Hw�<;��<zz�<��<k�<�ܶ<�I�<���<I�<�w�<wԮ<9-�<<��<�ө<�!�<2l�<���<���<P9�<�w�<���<�<$�<�X�<'��<���<7�<�<&B�<�k�<�<Ⱥ�<n��<�<�(�<SK�<Tm�<b}<�^y<؟u<�q<�n<�_j<?�f<6�b<�_<�`[<ȢW<��S<a*P<UpL<��H<�E<�MA<ϛ=<��9<q@6<7�2<`�.<4O+<��'<<$<;� <��<.b<��<GX<��<�d<F�<�<1&<Β�;S��;�J�;��;:?�;]��;�t�;�(�;���;`��;+��;���;ں�;\ݩ;{�;f]�;�;�,�;���;�L�;���;[z{;J'q;/�f;��\;�S;�gI;��?;Sp6;c--; $;�;X<;o�	;@� ;T�:_]�:���:o˿:$ٯ:��:i��:�M�:"ad:��F:):�:;�9�I�9��Y9���8� |�&\��i]�S���vٹ��>5!�K#;���T�ejn�,僺̀������z��Dݵ�V.º�oκz�ں_��@�����Ns��l�$a�nP��;��"#��)���.���4�|�:�2q@�GEF��L�J�Q�H�W��]�Rc��i�K�n���t�cz�'%���
�������ֈ�h���q���W����t���^���H���  �  Tz=�=�=�`=�=[�=�E=�� =�� =I( =!��<"��<w�<O�<���<��<��<�A�<�|�<2��<���<�&�<]�<q��<���<~��<+�<N[�<��<H��<��<�<Z5�<�[�<���<Q��<���<���<���<�<�0�<�E�<�X�<]h�<}u�<��<φ�<Њ�<���<��<��<by�<l�<[�<F�<-�<�<���<^��<U��<�p�<�=�<N�<���<È�<�B�<���<��<AS�<���<ٚ�<)7�<���<�`�<��<Mw�<O��<�z�<��<!k�<�ܶ<�I�<���<Q�<�w�<tԮ<9-�<;��<�ө<�!�<7l�<���<���<C9�<�w�<ó�<��<�#�<�X�<&��<���<(�<��<B�<�k�<ᓋ<ƺ�<p��<��<�(�<VK�<em�<a}<_y<�u<�q<�n<�_j<o�f<8�b<�_<�`[<٢W<�S<Y*P<rpL<�H<�E<�MA<ϛ=<��9<U@6<G�2<D�.<O+<��'<C$<?� <��<b<`�<bX<��<�d<+�<щ<8&<���;V��;J�;���;6?�;���;�t�;p(�;Y��;{��;J��;���;⺯;�ݩ;��;x]�;뺘;�,�;���;�L�;���;/z{;g'q;��f;��\;�S;ngI;�?;�o6;�,-;�$;�;�;;��	;�� ;!�:?^�:A��:ʿ:�د:��:V��:FM�:�ad:��F:x):=�:�>�9K�9��Y9���8��{�mS�h]�N���tٹ�*4!��";���T�kn��䃺���)���z��gݵ�9.º[pκ?�ں���������\s�^l��a��P�K<��"#��)�{�.�[�4��:��p@��EF��L�:�Q���W��]��Qc�ni�S�n��t�z�'%���
������nֈ�e���g���J����t��+^���H���  �  Rz=�=�=�`=�=W�=�E=�� =�� =D( =��<��<a�<O�<��<��<f�<�A�<�|�<*��<���<|&�<]�<c��<���<���<+�<Q[�<��<S��<��<�<g5�<�[�<���<W��<	��<���<��<�<�0�<�E�<�X�<dh�<~u�<��<���<ʊ�<���<���<��<Ry�<l�<�Z�<F�<-�<�<���<@��<R��<�p�<�=�<C�<���<���<�B�<���<��<IS�<���<���<17�<���<a�<��<`w�<V��<�z�<)��<-k�<�ܶ<�I�<���<S�<�w�<{Ԯ<=-�<=��<�ө<�!�<-l�<���<���<69�<�w�<���<��<�#�<�X�<��<���<(�<��<B�<�k�<���<���<c��<�<�(�<[K�<`m�<v}<_y<��u<G�q< n<�_j<u�f<c�b<�_<�`[<�W<�S<q*P<lpL<�H<�E<�MA<��=<��9<Z@6</�2<O�.<�N+<��'<$<� <��<�a<Z�<&X<~�<�d<�<ω<"&<���;��;wJ�;��;C?�;���;�t�;�(�;3��;���;|��;֫�;��;�ݩ;��;�]�;c��;�,�;���;�L�;���;dz{;h'q;#�f;\�\;zS;(gI;��?;�o6;T,-;�$;�;�;;φ	;�� ;��:S\�:	��:wɿ:=د:��:���:M�:�_d:^�F:�):*�:�?�9�L�9Y�Y9��8�-x�pI��^]��L���rٹ��2!�� ;���T��in��䃺������z��Rݵ�+/º&pκڢںU��=������s�Ym��a�KQ�r<�G##�c)�u�.���4�ؚ:�Xq@��EF��L���Q�J�W���]��Qc��i���n��t��~z��$��q
��D���cֈ����<���󋑻�t��<^���H���  �  Sz=�=�=�`=�=X�=�E=�� =�� =>( =��<��<^�<O�<ߌ�<��<]�<�A�<|�< ��<���<p&�<	]�<g��<���<���<+�<T[�<��<h��<��<�<a5�<�[�<���<V��<��<���<��<�<�0�<�E�<�X�<ph�<vu�<��<ǆ�<Ί�<���<��<��<Ny�<l�<�Z�<F�<-�<�<���<7��<[��<�p�<�=�<>�<���<È�<�B�<���<��<RS�<���<��<A7�<���<a�<��<hw�<X��<�z�<(��<&k�<�ܶ<�I�<���<U�<�w�<}Ԯ<:-�<F��<�ө<�!�<$l�<���<���<39�<�w�<���<�<�#�<�X�<��<���<*�<��<B�<�k�<䓋<���<n��<
�<�(�<fK�<am�<�}<._y<
�u<E�q<�n<�_j<n�f<��b<�_<�`[<�W<�S<�*P<ppL<&�H<�E<�MA<ԛ=<��9<^@6<�2<O�.<�N+<��'<$<� <��<�a<j�<X<��<�d<�<щ<
&<���;+��;�J�;��;6?�;���;�t�;�(�;2��;���;d��;���;]��;�ݩ;��;t]�;j��;�,�;貍;�L�;���;�z{;$'q;j�f;��\;�S;,gI;`�?;�o6;1,-;�$;�;�;;{�	;)� ;%�:�[�:���:@ɿ:�ׯ:��:w��:7M�:�`d:ЉF:�):�:�?�9�L�9�Y9w��8��w��S�7[]�SL���oٹK��3!��;���T��fn��䃺�������z���ܵ��.ºpκy�ںW����������s��m��a��Q��<�H##��)�l�.��4�̚:��q@��EF��L�G�Q��W�/�]�vQc��i���n�ѳt��~z��$���
�����rֈ�˼��_��� ����t��&^���H���  �  Uz=�=�=�`=�=U�=�E=�� =�� =?( =��<��<X�<�N�<݌�<���<^�<�A�<t|�<"��<���<z&�<�\�<e��<���<���<!+�<][�<��<[��<��<!�<w5�<�[�<���<\��<��<���<��<�<�0�<�E�<�X�<ph�<�u�<��<Ȇ�<���<���<���<��<My�<�k�<�Z�<�E�<
-�<�<���<:��<C��<�p�<�=�<D�<���<���<�B�<���<��<US�<���<ߚ�<>7�<���<a�<��<qw�<^��<�z�<4��<>k�<�ܶ<�I�<���<V�<�w�<�Ԯ<B-�<=��<�ө<�!�<-l�<���<���<,9�<�w�<���<��<�#�<�X�<	��<���<�<��<B�<�k�<ٓ�<���<k��<�<�(�<fK�<em�<w}<:_y<�u<X�q<! n<�_j<x�f<��b<�_<a[<�W<#�S<{*P<vpL<,�H<�E<�MA<ɛ=<��9<F@6<%�2<A�.<�N+<p�'<$<� <r�<�a<=�<X<l�<�d<�<ǉ<&<g��; ��;xJ�;��;Q?�;���;�t�;�(�;a��;���;���;���;b��;�ݩ;�;�]�;���;'-�;鲍;�L�;��;�z{;�'q;�f;��\;/S;gI;��?;�o6;-,-;4$;�;6;;C�	;
� ;� �:�[�:��:ɿ:�ׯ:��:���:IL�:�`d:b�F:>):w�:�A�9-L�9�Y9	��8��v�>�BW]��J��Mnٹ���0!�T;��T�zhn�䃺�~��M��xz��]ݵ��.ºqκ�ںf�����b���t��m�Fb��Q��<��##��)���.��4���:�zq@��EF�)L�]�Q�:�W���]�uQc�gi���n���t�i~z��$��R
�����^ֈ�Ѽ�����͋��st���]���H���  �  �x=�=|�=$^=��=۠=�A=�� =
� =J# =T��<���<��<�A�<�~�<��<���<1�<�j�<h��<���<��<G�<|{�<��<X��<��<�?�<em�<Q��<���<w��<��<�8�<\�<\}�<���<ȹ�<���<O��<t�< �<?(�<z6�<!B�<�J�<WP�<�R�<R�<�M�<zF�<�;�<�,�<w�<�<���<���<6��<���<�W�<c(�<z��<��<�<\=�<���<���<�[�<��<4��<�N�<1��<��<��<��<�-�<]��<�2�<'��<J%�<��<��<�p�<�ֱ<9�<=��<��<oH�<���<p�<�7�<1��<�Ǣ<�
�<{K�<y��<�ě<���<�4�<#i�<ě�<a̒<T��<x(�<(T�<z~�<v��<9χ<���<��<W@�<�d�<�}<�Uy<��u<��q<#n<�fj<��f<��b<A3_<ex[<��W<�T<FNP<��L<�H<2E<�A<T�=<^):<#�6<
�2<P:/<g�+<(<�k$<�� <jL<��<L@<F�<�I<��<�i</<Q�<X��;L��;=Z�;���; \�;���;ٝ�;W�;O"�;*��;��;�;0 �;&�;�^�;��;R
�;�}�;y�;잉;MM�;O~;�s;s�i;��_;��U;)�K;�bB;P�8;�/;p�&;|~;��;��;�?;S��:��:H�:9�:���:&�:��:!�:��k:��M:�0:��:#��9..�9��r9��9W��7����G����FϹ�*��z�Җ6�~zP��5j��ށ�"����*��o���/(��'����̺b$ٺ�Z庽��^�������
����(��޻���"��(��y.�\4��<:��@���E���K���Q�wW�(J]�3c���h�0�n�3�t��_z�%��- ���腻rш�Ѻ������<���yz��tf�� T���  �  �x=�=y�= ^=��=Ԡ=�A=�� =� =D# =K��<t��<��<�A�<�~�<��<v��<1�<�j�<`��<��<��< G�<n{�<���<G��<��<�?�<Nm�<P��<���<���<��<�8�<	\�<Y}�<���<Ϲ�<���<A��<q�<�<+(�<�6�<B�<�J�<QP�<�R�<R�<N�<�F�<z;�<�,�<]�<�<���<���<>��<���<�W�<R(�<���<*��<!�<\=�<���<���<�[�<��<$��<�N�<-��<��<��<(��<�-�<[��<�2�<,��<[%�<��<��<�p�<�ֱ<9�<?��<��<rH�<���<t�<8�<X��<�Ǣ<�
�<vK�<c��<�ě<���<�4�< i�<���<[̒<I��<�(�<CT�<�~�<i��<3χ<���<��<b@�<ud�<�}<�Uy<��u<�q<
#n<�fj<��f<��b<E3_<�x[<��W<�T<=NP<Y�L<-�H<�1E<߁A<P�=<A):<2�6<=�2<�:/<P�+<�(<�k$<�� <xL<��<a@<�<wI<��<�i<{<�<g��;��;FZ�;h��;!\�;���;}��;W�;�!�;f��;��;*�;3 �;�%�;�^�;/��;�
�;�}�;j�;ƞ�;M�;�~;��s;��i;{�_;��U;��K;�cB;��8;��/;D�&;�};��;��;�?;у�:P��:�G�:+�:H��::(�:��:"!�:��k:l�M:�0:��:!��9G*�9��r9�9��7P��)�G��Ù�oFϹJ*��x�U�6�/}P��5j����U����*�������'��������̺�"ٺ3X��� ���>����
����k�����ĩ"�˓(��y.�e\4��;:��@�K�E�	�K�-�Q�>wW��J]��c�c�h�T�n���t��_z����" ���腻�ш�������������wz���f��T���  �  �x=�=w�=!^=��=ՠ=�A=�� =� =A# =g��<���<��<�A�<�~�<��<x��<1�<�j�<V��<��<��<)G�<i{�<���<B��<��<�?�<Jm�<g��<���<���<|�<�8�<\�<V}�<���<���<���<5��<|�<!�<'(�<�6�<B�<�J�<LP�<�R�<R�<�M�<�F�<v;�<�,�<`�<1�<���<���<T��<���<�W�<T(�<y��<��<�<h=�<���<«�<�[�<��<"��<�N�<;��<��<��<��<�-�<Z��<�2�<��<?%�<��<w�<�p�<�ֱ<9�<E��<��<|H�<���<~�<�7�<D��<�Ǣ<�
�<�K�<c��<�ě<���<�4�<0i�<���<x̒<B��<�(�<)T�<�~�<n��<2χ<���<��<r@�<pd�<�}<�Uy<��u<�q<�"n<�fj<��f<��b<3_<rx[<{�W<�T<hNP<K�L<G�H<�1E<�A<R�=<E):<<�6<�2<n:/<D�+<*(<�k$<�� <�L<��<�@<$�<�I<��<�i<[<K�<���;��;jZ�;W��;0\�;���;n��;rW�;�!�;^��;u�;��;$ �;�%�;�^�;���;�
�;s}�;��;�;�L�;
~;8�s;Кi;T�_;�U;;�K;cB;��8;k�/;.�&;�};c�;��;�?;1��:D��:�I�:Q�:���:�&�:&��:�!�:��k:��M:�0:1�:���9,�9��r9p�9!�7�.����G��Ù��FϹ,�a|���6��~P�43j�/������<*�����W'��V���,�̺t$ٺkY庫����������
������r��B�"��(��x.��\4�%<:�y@�R�E���K�7�Q�wW��J]�_c���h�ɾn���t�(`z����~ ���腻�ш�����פ��!����z���f���S���  �  �x=�=v�=%^=��=۠=�A=�� =� =H# =\��<}��<�<�A�<�~�<��<���<1�<�j�<j��<��<��</G�<m{�<���<N��<��<�?�<Im�<Q��<���<���<��<�8�<�[�<I}�<���<���<���<>��<k�<�<&(�<�6�<B�<�J�<IP�<�R�<R�<N�<�F�<�;�<�,�<f�<&�<���<���<J��<���<�W�<Y(�<���<&��<�<p=�<���<«�<�[�<��<��<�N�<'��<��<��<��<�-�<K��<y2�</��<F%�<��<~�<�p�<�ֱ< 9�<9��<��<xH�<���<��<�7�<U��<�Ǣ<�
�<|K�<o��<�ě<���<�4�<+i�<���<j̒<L��<�(�<;T�<�~�<{��<.χ<���<��<]@�<pd�<�}<�Uy<��u<��q<�"n<�fj<o�f<��b<B3_<kx[<��W<�T<ANP<N�L< �H<�1E<�A<F�=<[):<?�6<&�2<�:/<a�+<(<�k$<�� <�L<��<t@<:�<�I<��<�i<~<e�<���;��;[Z�;���;\�;���;o��;W�;�!�;U��;��;?�;���;�%�;�^�;쪟;�
�;�}�;W�;���;�L�;�~;��s;�i;9�_;6�U;Y�K;�cB;A�8;��/;��&;�};�;��;�?;���:���:H�:��:��:(�:���:c"�:��k:��M:�0:{�:��9�(�9
�r9��9�͛7,#����G�Ǚ�[JϹ�)�T{��6��}P��5j�u���Ï���*��=����'��;�����̺�#ٺZX�J��c�����D�
�D��)�����g�"�h�(�my.�I\4��;:��@�I�E�w�K�[�Q��vW��J]�
c���h�i�n���t��_z���9 ���腻�ш�溋�����/����z���f��	T���  �  �x=�=y�="^=��=۠=�A=�� =� =J# =`��<���<�<�A�<�~�<��<���<1�<�j�<g��<��<��<G�<v{�<���<K��<��<�?�<Um�<E��<���<r��<s�<�8�<�[�<O}�<���<���<���<=��<i�<�<2(�<6�<B�<�J�<TP�<�R�<R�<N�<�F�<�;�<�,�<��<(�<���<���<H��<�<�W�<d(�<���<)��<�<c=�<���<���<�[�<��<(��<�N�<#��<��<��<��<{-�<K��<s2�<��<=%�<���<��<�p�<�ֱ<9�<9��<��<qH�<���<t�<�7�<V��<�Ǣ<�
�<�K�<���<�ě<���<�4�<6i�<Л�<o̒<U��<�(�<GT�<r~�<x��<3χ<���<��<Z@�<|d�<�}<�Uy<��u<��q<�"n<�fj<��f<��b<'3_<@x[<s�W<�T<-NP<e�L< �H<�1E<�A<L�=<^):<�6<?�2<�:/<h�+<(<�k$<� <�L< �<f@<n�<�I<��<�i<~<y�<`��;8��;LZ�;~��;\�;���;���;�V�;�!�;��;V�;��;���;�%�;�^�;窟;4
�;�}�;O�;���;M�;|~;��s;��i;��_;�U;�K;�cB;��8;�/;ځ&;�~;&�;g�;�@;���:���:�H�:X�:1��:=(�:8��:�!�:7�k:��M:(0:?�:���92*�9Y�r98�9�w�7$����G��ƙ��KϹ�,�j|�Q�6�Z}P�7j��߁�`����*��{����'�������̺m#ٺ;X庤��ך�����h�
�v�����j��
�"���(�Ey.�\4��;:��@���E���K�0�Q�wW�uJ]�c�/�h���n���t�`z�f��c ��酻�ш����ä�������z���f��1T���  �  �x=�=x�=#^=��=ܠ=�A=�� =� =O# =q��<���<�<�A�<�~�<$��<���<1�<�j�<m��<��<��<*G�<x{�<���<K��<��<�?�<@m�<I��<���<t��<w�<�8�<�[�<N}�<z��<���<���<3��<_�<�<(�<�6�<B�<�J�<WP�<�R�<R�<N�<�F�<�;�<�,�<w�<6�<��<���<W��<���<�W�<w(�<���<+��<�<g=�<���<���<�[�<��<��<�N�<��<���<��<
��<g-�<M��<t2�<��<=%�<���<q�<�p�<�ֱ<�8�<>��<��<sH�<���<}�<�7�<R��<�Ǣ<�<�K�<���<�ě<���<�4�<?i�<ś�<|̒<a��<�(�<GT�<�~�<w��<7χ<���<��<Z@�<gd�<�}<�Uy<��u<��q<�"n<�fj<��f<s�b<3_<Ux[<s�W<�T<2NP<<�L<�H<�1E<�A<T�=<_):<?�6<?�2<�:/<|�+<?(<�k$<� <�L<#�<�@<d�<�I<��<�i<t<|�<���;B��;[Z�;���;)\�;u��;N��;�V�;�!�;#��;i�;��;���;�%�;N^�;˪�;W
�;s}�;+�;���;�L�;�~;��s;��i;��_;��U;��K;�cB;��8;��/;5�&;�~;��;��;~@;s��:��:yI�:��:��:k(�::�!�:_�k:��M:�0:��:���9�'�97�r9��9I��7o)���G�fƙ�WKϹ]/�N|�+�6�:P��6j� ၺ�����*�������'��o����̺F#ٺrX�l��s��������
���������Ȩ"��(��x.��[4��;:��@�<�E���K��Q�wW��J]�c���h���n�"�t�<`z�<��� ��:酻�ш�A�������[����z���f��$T���  �  �x=�=s�="^=��=٠=�A=�� =#� =M# =p��<���< �<�A�<�~�<4��<���<$1�<�j�<s��<-��<��<2G�<p{�<���<G��<��<�?�<Fm�<J��<���<g��<h�<�8�<�[�<2}�<���<���<���<+��<X�<�<(�<�6�<B�<�J�<QP�<�R�< R�<N�<�F�<�;�<�,�<��<D�<��<���<f��<Ă�<�W�<n(�<���<6��< �<l=�<���<���<�[�<��<��<�N�<��<ׂ�<��<���<q-�<0��<_2�<	��<.%�<<g�<�p�<�ֱ<�8�<2��<��<vH�<���<��<�7�<d��<�Ǣ<�<�K�<���<�ě<���<�4�<Ii�<ԛ�<̒<\��<�(�<LT�<�~�<u��<3χ<���<��<^@�<gd�<�}<kUy<l�u<��q<�"n<�fj<N�f<o�b<3_<*x[<X�W<�T<?NP<;�L<#�H<�1E<�A<N�=<T):<P�6<E�2<�:/<w�+<>(<�k$<&� <�L<#�<�@<y�<�I<��<j<�<��<���;(��;fZ�;v��; \�;���;i��;W�;�!�;���;/�;��;���;g%�;|^�;���;
�;R}�;�;Ş�;�L�;�~;M�s;Ți;��_;�U;��K;8dB;��8;o�/;n�&;�~;�;��;�@;v��:���:J�:�:w��:)�:%��:K"�:��k:}�M:�0:a�:��9*�9��r9U�9�X�7:7����G�O͙�TPϹF.�~�̘6�b�P�17j�x���K���@+��Ͳ���'������̺�"ٺUW������G��_�
�I�����ĺ�s�"���(��x.��[4�&;:�b@���E���K�2�Q�wW��J]��c���h�R�n�t�t��`z����� ��,酻҈�H�����������z��'g��
T���  �  �x=�=v�=#^=��=ޠ=�A=�� = � =S# =~��<���<!�<�A�<�<.��<���<91�<�j�<}��<%��<��</G�<{{�<���<K��<��<�?�<@m�<0��<���<c��<Z�<�8�<�[�</}�<t��<���<~��<2��<J�<�<(�<x6�<B�<�J�<VP�<�R�<R�<N�<�F�<�;�<�,�<��<:�<��<���<\��<҂�<�W�<w(�<���<+��<�<q=�<���<���<�[�<��<��<~N�<��<ނ�<��<<`-�<+��<X2�<���<%�<闶<m�<�p�<�ֱ<�8�</��<��<sH�<���<��<�7�<[��<�Ǣ<�<�K�<���<�ě<��<�4�<Ei�<䛔<�̒<g��<�(�<GT�<�~�<���<6χ<���<��<V@�<dd�<�}<cUy<{�u<��q<�"n<lfj<Q�f<R�b<�2_<x[<^�W<�T<NP<5�L<�H<�1E<�A<S�=<j):<E�6<D�2<�:/<��+<Z(<&l$<)� <�L<[�<�@<��<�I<��<j<�<��<���;X��;cZ�;���;\�;v��;W��;�V�;�!�;���;��;��;{��;`%�;9^�;u��;�	�;s}�;��;���;�L�;R~;��s;��i;��_;l�U;��K;�cB;��8;��/;ׂ&;a;��;`�;wA;؅�:���:�J�:��:���:t(�:��:�"�:_�k:��M:�0:\�:��9'�9��r9C�9�-�70C���G�BΙ��QϹ�/���r�6��P��:j���������i+�������'��M�����̺#ٺ�W�=�J������
�
�������g����"�
�(�^x.�q[4�>;:��@�/�E�U�K��Q�wW��J]�@c���h��n���t�b`z����� ��l酻҈�����1���ޏ���z��g��iT���  �  �x=�=v�=!^=��=ޠ=�A=�� =� =\# =|��<���</�<�A�<	�<;��<���<.1�<�j�<���<$��<��<-G�<}{�<���<G��<��<�?�<@m�<7��<���<V��<d�<�8�<�[�<3}�<`��<���<{��<��<G�<�<(�<q6�<B�<�J�<XP�<�R�<1R�<$N�<�F�<�;�<�,�<��<N�<��<���<n��<Ղ�<�W�<�(�<���<7��<3�<l=�<���<���<�[�<��<��<|N�< ��<Ȃ�<��<���<O-�<-��<S2�<�<)%�<ݗ�<\�<�p�<�ֱ<�8�<.��<��<pH�<���<��<8�<^��<�Ǣ<�<�K�<���<�ě<	��<�4�<Wi�<ݛ�<�̒<w��<�(�<\T�<�~�<~��<6χ<���<��<G@�<cd�<�}<VUy<O�u<��q<�"n<Ffj<M�f<3�b<�2_<#x[<:�W<xT<NP<6�L<��H<�1E<�A<Q�=<i):<R�6<m�2<�:/<��+<X(<l$<G� <�L<c�<�@<��<�I<�<=j<�<��<���;_��;_Z�;}��;\�;1��;V��;�V�;!�;���;&�;m�;`��;o%�;�]�;���;�	�;}�;��;���;�L�;~;��s;��i;ē_;:�U;8�K;sdB;��8;&�/;Ȃ&;k;`�;M�;cA;���:��:�J�:f�:&��:@)�:o��:R"�:��k:��M:�0:��:�~�9�&�9��r9�9N�7/9��+�G��͙��RϹ�1�x~���6���P��9j�ၺ����k+�������'�������̺�!ٺ�W庄~����������
������F����"�A�(�kx.��Z4�d;:��@���E�_�K��Q�+wW��J]��c���h��n�ʐt�az����� ���酻҈�����7�������{��Bg��^T���  �  �x=�=t�= ^=��=ܠ=�A=�� =$� =[# =���<���<?�<�A�<�~�<N��<���<F1�<�j�<���<(��<��<0G�<x{�<���<A��<��<�?�<4m�<@��<���<Q��<L�<~8�<�[�< }�<f��<���<r��<��<O�<�<(�<�6�< B�<�J�<[P�<�R�<*R�<N�<�F�<�;�<-�<��<h�<��<���<���<ׂ�<�W�<�(�<���<0��<*�<l=�<���<���<�[�<��<��<xN�<��<���<��<ۣ�<Q-�<��<D2�<筹<%�<֗�<P�<�p�<�ֱ<�8�<6��<��<zH�<���<��<	8�<]��<�Ǣ<�<�K�<���<ś<���<�4�<ji�<훔<�̒<u��<�(�<PT�<�~�<{��<:χ<���<��<Z@�<Xd�<�}<YUy<@�u<��q<�"n<Vfj<&�f<>�b<�2_<�w[<-�W<uT<NP<�L<�H<�1E<߁A<Z�=<a):<O�6<U�2<�:/<��+<i(<:l$<f� <�L<G�<�@<��< J<�<<j<�<��<���;P��;�Z�;e��;'\�;u��;+��;�V�;Z!�;���;��;I�;A��;&%�;^�;3��;�	�;�|�;��;���;�L�;�~;2�s;Ӛi;ߓ_;8�U;�K;2dB;��8;	�/;\�&;�;2�;q�;pA;���:,��:�K�:C�:y��:�(�:狔:c"�:��k:��M:0:q�:z�9�%�9��r9΃9Z��7�U����G�ҙ�zVϹ"2����6���P�08j��ၺِ���*��T���6'��[�����̺G"ٺ�W�c~񺪘��E����
�g�������g�"�(�x.�[4� ;:�>@���E�w�K���Q�wW��J]�!c�L�h�ܿn���t�Oaz����$���酻n҈������������/{��Hg��TT���  �  |x=�=o�=#^=��=ޠ=�A=�� =.� =Z# =���<���<,�<B�<
�<S��<���<K1�<�j�<���<=��<��<EG�<t{�<���<D��<��<�?�<"m�<+��<���<`��<H�<�8�<�[�<}�<m��<~��<���<��<9�<��<(�<x6�< B�<�J�<NP�<�R�<2R�<"N�<�F�<�;�<
-�<��<W�<,��<���<}��<̂�<�W�<w(�<���<:��<.�<y=�<���<���<�[�<��<���<eN�<���<���<��<ϣ�<Y-�<��<B2�<�<%�<时<F�<�p�<�ֱ<�8�<*��<��<vH�<���<��<	8�<p��<�Ǣ<�<�K�<���<ś<��<�4�<Ui�<뛔<�̒<p��<�(�<PT�<�~�<���</χ<���<{�<U@�<Jd�<�}<4Uy<U�u<��q<u"n<bfj<��f<E�b<�2_<x[<C�W<UT<�MP<�L<�H<�1E<�A<K�=<i):<s�6<S�2<�:/<��+<f(<?l$<A� <M<g�<�@<��<J<�<Ij<�<��<��;A��;tZ�;s��;�[�;n��;��;�V�;4!�;���;��;h�;L��;�$�;&^�; ��;
�;}�;��;G��;tL�;]~;/�s;�i;��_;��U;L�K;edB;��8;ʩ/;~�&;R;��;��;�A;���:w��:8L�:��:���:t)�:,��:=#�:G�k:��M:60:��:�}�9K!�9��r9�9�7�7a��X�G��ԙ��VϹ�0�u����6�=�P�	;j��⁺����+�����k'�������̺A"ٺsV床}�=������
�m���������"�Б(��w.�+[4�M::�C@�o�E�F�K�Q�Q��vW�K]�Ic���h�a�n�P�t��`z����J��~酻�҈�������������{���g���T���  �  �x=�=o�="^=��=ߠ=�A=�� ="� =\# =���<���<>�<	B�<�<T��<���<P1�<�j�<���<-��<��<6G�<|{�<���<G��<��<�?�<<m�<9��<���<D��<@�<s8�<�[�<}�<Z��<��<j��<��<E�<�<(�<n6�<B�<�J�<UP�<�R�<0R�<!N�<�F�<�;�<-�<��<d�<+��<���<���<��<�W�<�(�<���<5��</�<p=�<���<���<�[�<��<��<{N�<���<���<��<У�<D-�<��<?2�<ܭ�<%�<ɗ�<K�<�p�<�ֱ<�8�<!��<��<mH�<���<��<8�<d��<�Ǣ<�<�K�<���<ś<��<�4�<hi�<���<�̒<x��<�(�<UT�<�~�<���<2χ<���<�<M@�<ed�<�}<EUy<&�u<|�q<o"n<Afj<�f<)�b<�2_<�w[<�W<aT<NP<7�L<�H<�1E<�A<H�=<m):<\�6<b�2<�:/<��+<s(<Yl$<f� <
M<t�<�@<��<J<�<Hj<�<��<Ք�;b��;WZ�;���;�[�;~��;L��;�V�;R!�;r��;��;!�;2��;%�;�]�;��;�	�;�|�;��;���;�L�;~;e�s;��i;��_;l�U;7�K;_dB;��8;<�/;��&;C�;�;��;�A;���:���:gL�:��:���:')�:5��:�"�:��k:t�M:0:�:��9�&�9��r9�9fǚ7=_����G��ә�xWϹr3���)�6���P��9j�2ၺ����/,��ٲ���'��<���i�̺�!ٺ4W�~�}������,�
�X��b�����}�"�;�(��w.��Z4�;:�@���E�N�K�9�Q�1wW��J]��c���h��n��t��az���V���酻�҈�ӻ������,���m{��pg��YT���  �  }x=�=w�="^=��=�=�A=�� =$� =e# =���<���<=�<B�<�<L��<���<<1�<�j�<���<2��<��<+G�<�{�<���<M��<��<�?�<m�< ��<���<G��<W�<t8�<�[�< }�<Q��<���<o��<��<E�<��<(�<j6�<B�<�J�<hP�<�R�<6R�<7N�<�F�<�;�<�,�<��<_�<+��<���<��<߂�<�W�<�(�<���<G��<<�<i=�<��<���<�[�<��<���<WN�<���<Ă�<��<룿<<-�<��<=2�<٭�<%�<͗�<Z�<�p�<�ֱ<�8�<)��<��<mH�<Û�<{�<"8�<k��<�Ǣ<%�<�K�<���<
ś<��<�4�<fi�<월<�̒<���<�(�<mT�<�~�<���<@χ<���<��<H@�<Nd�<V}<XUy<<�u<��q<�"n<0fj<)�f<�b<�2_<
x[< �W<wT<�MP<�L<��H<�1E<�A<[�=<t):<J�6<��2<�:/<՜+<l(<8l$<d� <M<|�<�@<��<�I<+�<Zj<�<أ<���;���;hZ�;���;\�;[��;؜�;mV�;�!�;���;��;"�;��;*%�;�]�;e��;�	�;}�;��;���;tL�;�~;��s;��i;K�_;N�U;k�K;eB;�8;�/;�&;�;�;��;�A;"��:���:�J�:��:���:T*�:��:A"�:��k:��M:.0:��:r}�9��9��r9��9ۚ7�C��ͱG��ҙ��WϹ�3�����6���P�
<j�;ぺ/����+��y����'��8����̺� ٺ�V庿}񺴗�����^�
����F�������"�ɑ(�4x.�FZ4��::�Y@���E�H�K�ɡQ�?wW��J]��c���h��n���t�\az�������酻f҈�򻋻����폑�I{��Cg���T���  �  �x=�=o�="^=��=ߠ=�A=�� ="� =\# =���<���<>�<	B�<�<T��<���<P1�<�j�<���<-��<��<6G�<|{�<���<G��<��<�?�<<m�<9��<���<D��<@�<s8�<�[�<}�<Z��<��<j��<��<E�<�<(�<n6�<B�<�J�<UP�<�R�<0R�<!N�<�F�<�;�<-�<��<d�<+��<���<���<��<�W�<�(�<���<5��</�<p=�<���<���<�[�<��<��<{N�<���<���<��<У�<D-�<��<?2�<ܭ�<%�<ɗ�<K�<�p�<�ֱ<�8�<!��<��<mH�<���<��<8�<d��<�Ǣ<�<�K�<���<ś<��<�4�<hi�<���<�̒<x��<�(�<UT�<�~�<���<2χ<���<�<M@�<ed�<�}<EUy<&�u<|�q<o"n<Afj<�f<)�b<�2_<�w[<�W<aT<NP<7�L<�H<�1E<�A<H�=<m):<\�6<b�2<�:/<��+<s(<Yl$<f� <
M<t�<�@<��<J<�<Hj<�<��<Ք�;b��;WZ�;���;�[�;~��;L��;�V�;R!�;r��;��;!�;2��;%�;�]�;��;�	�;�|�;��;���;�L�;~;e�s;��i;��_;l�U;7�K;_dB;��8;<�/;��&;C�;�;��;�A;���:���:gL�:��:���:')�:5��:�"�:��k:t�M:0:�:��9�&�9��r9�9fǚ7=_����G��ә�xWϹr3���)�6���P��9j�2ၺ����/,��ٲ���'��<���i�̺�!ٺ4W�~�}������,�
�X��b�����}�"�;�(��w.��Z4�;:�@���E�N�K�9�Q�1wW��J]��c���h��n��t��az���V���酻�҈�ӻ������,���m{��pg��YT���  �  |x=�=o�=#^=��=ޠ=�A=�� =.� =Z# =���<���<,�<B�<
�<S��<���<K1�<�j�<���<=��<��<EG�<t{�<���<D��<��<�?�<"m�<+��<���<`��<H�<�8�<�[�<}�<m��<~��<���<��<9�<��<(�<x6�< B�<�J�<NP�<�R�<2R�<"N�<�F�<�;�<
-�<��<W�<,��<���<}��<̂�<�W�<w(�<���<:��<.�<y=�<���<���<�[�<��<���<eN�<���<���<��<ϣ�<Y-�<��<B2�<�<%�<时<F�<�p�<�ֱ<�8�<*��<��<vH�<���<��<	8�<p��<�Ǣ<�<�K�<���<ś<��<�4�<Ui�<뛔<�̒<p��<�(�<PT�<�~�<���</χ<���<{�<U@�<Jd�<�}<4Uy<U�u<��q<u"n<bfj<��f<E�b<�2_<x[<C�W<UT<�MP<�L<�H<�1E<�A<K�=<i):<s�6<S�2<�:/<��+<f(<?l$<A� <M<g�<�@<��<J<�<Ij<�<��<��;A��;tZ�;s��;�[�;n��;��;�V�;4!�;���;��;h�;L��;�$�;&^�; ��;
�;}�;��;G��;tL�;]~;/�s;�i;��_;��U;L�K;edB;��8;ʩ/;~�&;R;��;��;�A;���:w��:8L�:��:���:t)�:,��:=#�:G�k:��M:60:��:�}�9K!�9��r9�9�7�7a��X�G��ԙ��VϹ�0�u����6�=�P�	;j��⁺����+�����k'�������̺A"ٺsV床}�=������
�m���������"�Б(��w.�+[4�M::�C@�o�E�F�K�Q�Q��vW�K]�Ic���h�a�n�P�t��`z����J��~酻�҈�������������{���g���T���  �  �x=�=t�= ^=��=ܠ=�A=�� =$� =[# =���<���<?�<�A�<�~�<N��<���<F1�<�j�<���<(��<��<0G�<x{�<���<A��<��<�?�<4m�<@��<���<Q��<L�<~8�<�[�< }�<f��<���<r��<��<O�<�<(�<�6�< B�<�J�<[P�<�R�<*R�<N�<�F�<�;�<-�<��<h�<��<���<���<ׂ�<�W�<�(�<���<0��<*�<l=�<���<���<�[�<��<��<xN�<��<���<��<ۣ�<Q-�<��<D2�<筹<%�<֗�<P�<�p�<�ֱ<�8�<6��<��<zH�<���<��<	8�<]��<�Ǣ<�<�K�<���<ś<���<�4�<ji�<훔<�̒<u��<�(�<PT�<�~�<{��<:χ<���<��<Z@�<Xd�<�}<YUy<@�u<��q<�"n<Vfj<&�f<>�b<�2_<�w[<-�W<uT<NP<�L<�H<�1E<߁A<Z�=<a):<O�6<U�2<�:/<��+<i(<:l$<f� <�L<G�<�@<��< J<�<<j<�<��<���;P��;�Z�;e��;'\�;u��;+��;�V�;Z!�;���;��;I�;A��;&%�;^�;3��;�	�;�|�;��;���;�L�;�~;2�s;Ӛi;ߓ_;8�U;�K;2dB;��8;	�/;\�&;�;2�;q�;pA;���:,��:�K�:C�:y��:�(�:狔:c"�:��k:��M:0:q�:z�9�%�9��r9΃9Z��7�U����G�ҙ�zVϹ"2����6���P�08j��ၺِ���*��T���6'��[�����̺G"ٺ�W�c~񺪘��E����
�g�������g�"�(�x.�[4� ;:�>@���E�w�K���Q�wW��J]�!c�L�h�ܿn���t�Oaz����$���酻n҈������������/{��Hg��TT���  �  �x=�=v�=!^=��=ޠ=�A=�� =� =\# =|��<���</�<�A�<	�<;��<���<.1�<�j�<���<$��<��<-G�<}{�<���<G��<��<�?�<@m�<7��<���<V��<d�<�8�<�[�<3}�<`��<���<{��<��<G�<�<(�<q6�<B�<�J�<XP�<�R�<1R�<$N�<�F�<�;�<�,�<��<N�<��<���<n��<Ղ�<�W�<�(�<���<7��<3�<l=�<���<���<�[�<��<��<|N�< ��<Ȃ�<��<���<O-�<-��<S2�<�<)%�<ݗ�<\�<�p�<�ֱ<�8�<.��<��<pH�<���<��<8�<^��<�Ǣ<�<�K�<���<�ě<	��<�4�<Wi�<ݛ�<�̒<w��<�(�<\T�<�~�<~��<6χ<���<��<G@�<cd�<�}<VUy<O�u<��q<�"n<Ffj<M�f<3�b<�2_<#x[<:�W<xT<NP<6�L<��H<�1E<�A<Q�=<i):<R�6<m�2<�:/<��+<X(<l$<G� <�L<c�<�@<��<�I<�<=j<�<��<���;_��;_Z�;}��;\�;1��;V��;�V�;!�;���;&�;m�;`��;o%�;�]�;���;�	�;}�;��;���;�L�;~;��s;��i;ē_;:�U;8�K;sdB;��8;&�/;Ȃ&;k;`�;M�;cA;���:��:�J�:f�:&��:@)�:o��:R"�:��k:��M:�0:��:�~�9�&�9��r9�9N�7/9��+�G��͙��RϹ�1�x~���6���P��9j�ၺ����k+�������'�������̺�!ٺ�W庄~����������
������F����"�A�(�kx.��Z4�d;:��@���E�_�K��Q�+wW��J]��c���h��n�ʐt�az����� ���酻҈�����7�������{��Bg��^T���  �  �x=�=v�=#^=��=ޠ=�A=�� = � =S# =~��<���<!�<�A�<�<.��<���<91�<�j�<}��<%��<��</G�<{{�<���<K��<��<�?�<@m�<0��<���<c��<Z�<�8�<�[�</}�<t��<���<~��<2��<J�<�<(�<x6�<B�<�J�<VP�<�R�<R�<N�<�F�<�;�<�,�<��<:�<��<���<\��<҂�<�W�<w(�<���<+��<�<q=�<���<���<�[�<��<��<~N�<��<ނ�<��<<`-�<+��<X2�<���<%�<闶<m�<�p�<�ֱ<�8�</��<��<sH�<���<��<�7�<[��<�Ǣ<�<�K�<���<�ě<��<�4�<Ei�<䛔<�̒<g��<�(�<GT�<�~�<���<6χ<���<��<V@�<dd�<�}<cUy<{�u<��q<�"n<lfj<Q�f<R�b<�2_<x[<^�W<�T<NP<5�L<�H<�1E<�A<S�=<j):<E�6<D�2<�:/<��+<Z(<&l$<)� <�L<[�<�@<��<�I<��<j<�<��<���;X��;cZ�;���;\�;v��;W��;�V�;�!�;���;��;��;{��;`%�;9^�;u��;�	�;s}�;��;���;�L�;R~;��s;��i;��_;l�U;��K;�cB;��8;��/;ׂ&;a;��;`�;wA;؅�:���:�J�:��:���:t(�:��:�"�:_�k:��M:�0:\�:��9'�9��r9C�9�-�70C���G�BΙ��QϹ�/���r�6��P��:j���������i+�������'��M�����̺#ٺ�W�=�J������
�
�������g����"�
�(�^x.�q[4�>;:��@�/�E�U�K��Q�wW��J]�@c���h��n���t�b`z����� ��l酻҈�����1���ޏ���z��g��iT���  �  �x=�=s�="^=��=٠=�A=�� =#� =M# =p��<���< �<�A�<�~�<4��<���<$1�<�j�<s��<-��<��<2G�<p{�<���<G��<��<�?�<Fm�<J��<���<g��<h�<�8�<�[�<2}�<���<���<���<+��<X�<�<(�<�6�<B�<�J�<QP�<�R�< R�<N�<�F�<�;�<�,�<��<D�<��<���<f��<Ă�<�W�<n(�<���<6��< �<l=�<���<���<�[�<��<��<�N�<��<ׂ�<��<���<q-�<0��<_2�<	��<.%�<<g�<�p�<�ֱ<�8�<2��<��<vH�<���<��<�7�<d��<�Ǣ<�<�K�<���<�ě<���<�4�<Ii�<ԛ�<̒<\��<�(�<LT�<�~�<u��<3χ<���<��<^@�<gd�<�}<kUy<l�u<��q<�"n<�fj<N�f<o�b<3_<*x[<X�W<�T<?NP<;�L<#�H<�1E<�A<N�=<T):<P�6<E�2<�:/<w�+<>(<�k$<&� <�L<#�<�@<y�<�I<��<j<�<��<���;(��;fZ�;v��; \�;���;i��;W�;�!�;���;/�;��;���;g%�;|^�;���;
�;R}�;�;Ş�;�L�;�~;M�s;Ți;��_;�U;��K;8dB;��8;o�/;n�&;�~;�;��;�@;v��:���:J�:�:w��:)�:%��:K"�:��k:}�M:�0:a�:��9*�9��r9U�9�X�7:7����G�O͙�TPϹF.�~�̘6�b�P�17j�x���K���@+��Ͳ���'������̺�"ٺUW������G��_�
�I�����ĺ�s�"���(��x.��[4�&;:�b@���E���K�2�Q�wW��J]��c���h�R�n�t�t��`z����� ��,酻҈�H�����������z��'g��
T���  �  �x=�=x�=#^=��=ܠ=�A=�� =� =O# =q��<���<�<�A�<�~�<$��<���<1�<�j�<m��<��<��<*G�<x{�<���<K��<��<�?�<@m�<I��<���<t��<w�<�8�<�[�<N}�<z��<���<���<3��<_�<�<(�<�6�<B�<�J�<WP�<�R�<R�<N�<�F�<�;�<�,�<w�<6�<��<���<W��<���<�W�<w(�<���<+��<�<g=�<���<���<�[�<��<��<�N�<��<���<��<
��<h-�<M��<t2�<��<=%�<���<q�<�p�<�ֱ<�8�<>��<��<sH�<���<}�<�7�<R��<�Ǣ<�<�K�<���<�ě<���<�4�<?i�<ś�<|̒<a��<�(�<GT�<�~�<w��<7χ<���<��<Z@�<gd�<�}<�Uy<��u<��q<�"n<�fj<��f<s�b<3_<Ux[<s�W<�T<2NP<<�L<�H<�1E<�A<T�=<_):<?�6<?�2<�:/<|�+<?(<�k$<� <�L<#�<�@<d�<�I<��<�i<t<|�<���;B��;[Z�;���;)\�;u��;N��;�V�;�!�;#��;i�;��;���;�%�;N^�;˪�;W
�;s}�;+�;���;�L�;�~;��s;��i;��_;��U;��K;�cB;��8;��/;5�&;�~;��;��;~@;s��:��:yI�:��:��:k(�::�!�:_�k:��M:�0:��:���9�'�97�r9��9I��7o)���G�fƙ�WKϹ]/�N|�+�6�:P��6j� ၺ�����*�������'��o����̺F#ٺrX�l��s��������
���������Ȩ"��(��x.��[4��;:��@�<�E���K��Q�wW��J]�c���h���n�"�t�<`z�<��� ��:酻�ш�A�������[����z���f��$T���  �  �x=�=y�="^=��=۠=�A=�� =� =J# =`��<���<�<�A�<�~�<��<���<1�<�j�<g��<��<��<G�<v{�<���<K��<��<�?�<Um�<E��<���<r��<s�<�8�<�[�<O}�<���<���<���<=��<i�<�<2(�<6�<B�<�J�<TP�<�R�<R�<N�<�F�<�;�<�,�<��<(�<���<���<H��<�<�W�<d(�<���<)��<�<c=�<���<���<�[�<��<(��<�N�<#��<��<��<��<{-�<K��<s2�<��<=%�<���<��<�p�<�ֱ<9�<9��<��<qH�<���<t�<�7�<V��<�Ǣ<�
�<�K�<���<�ě<���<�4�<6i�<Л�<o̒<U��<�(�<GT�<r~�<x��<3χ<���<��<Z@�<|d�<�}<�Uy<��u<��q<�"n<�fj<��f<��b<'3_<@x[<s�W<�T<-NP<e�L< �H<�1E<�A<L�=<^):<�6<?�2<�:/<h�+<(<�k$<� <�L< �<f@<n�<�I<��<�i<~<y�<`��;8��;LZ�;~��;\�;���;���;�V�;�!�;��;V�;��;���;�%�;�^�;窟;4
�;�}�;O�;���;M�;|~;��s;��i;��_;�U;�K;�cB;��8;�/;ځ&;�~;&�;g�;�@;���:���:�H�:X�:1��:=(�:8��:�!�:7�k:��M:(0:?�:���92*�9Y�r98�9�w�7$����G��ƙ��KϹ�,�j|�Q�6�Z}P�7j��߁�`����*��{����'�������̺m#ٺ;X庤��ך�����h�
�v�����j��
�"���(�Ey.�\4��;:��@���E���K�0�Q�wW�uJ]�c�/�h���n���t�`z�f��c ��酻�ш����ä�������z���f��1T���  �  �x=�=v�=%^=��=۠=�A=�� =� =H# =\��<}��<�<�A�<�~�<��<���<1�<�j�<j��<��<��</G�<m{�<���<N��<��<�?�<Im�<Q��<���<���<��<�8�<�[�<I}�<���<���<���<>��<k�<�<&(�<�6�<B�<�J�<IP�<�R�<R�<N�<�F�<�;�<�,�<f�<&�<���<���<J��<���<�W�<Y(�<���<&��<�<p=�<���<«�<�[�<��<��<�N�<'��<��<��<��<�-�<K��<y2�</��<F%�<��<~�<�p�<�ֱ< 9�<9��<��<xH�<���<��<�7�<U��<�Ǣ<�
�<|K�<o��<�ě<���<�4�<+i�<���<j̒<L��<�(�<;T�<�~�<{��<.χ<���<��<]@�<pd�<�}<�Uy<��u<��q<�"n<�fj<o�f<��b<B3_<kx[<��W<�T<ANP<N�L< �H<�1E<�A<F�=<[):<?�6<&�2<�:/<a�+<(<�k$<�� <�L<��<t@<:�<�I<��<�i<~<e�<���;��;[Z�;���;\�;���;o��;W�;�!�;U��;��;?�;���;�%�;�^�;쪟;�
�;�}�;W�;���;�L�;�~;��s;�i;9�_;6�U;Y�K;�cB;A�8;��/;��&;�};�;��;�?;���:���:H�:��:��:(�:���:c"�:��k:��M:�0:{�:��9�(�9
�r9��9�͛7,#����G�Ǚ�[JϹ�)�T{��6��}P��5j�u���Ï���*��=����'��;�����̺�#ٺZX�J��c�����D�
�D��)�����g�"�h�(�my.�I\4��;:��@�I�E�w�K�[�Q��vW��J]�
c���h�i�n���t��_z���9 ���腻�ш�溋�����/����z���f��	T���  �  �x=�=w�=!^=��=ՠ=�A=�� =� =A# =g��<���<��<�A�<�~�<��<x��<1�<�j�<V��<��<��<)G�<i{�<���<B��<��<�?�<Jm�<g��<���<���<|�<�8�<\�<V}�<���<���<���<5��<|�<!�<'(�<�6�<B�<�J�<LP�<�R�<R�<�M�<�F�<v;�<�,�<`�<1�<���<���<T��<���<�W�<T(�<y��<��<�<h=�<���<«�<�[�<��<"��<�N�<;��<��<��<��<�-�<Z��<�2�<��<?%�<��<w�<�p�<�ֱ<9�<E��<��<|H�<���<~�<�7�<D��<�Ǣ<�
�<�K�<c��<�ě<���<�4�<0i�<���<x̒<B��<�(�<)T�<�~�<n��<2χ<���<��<r@�<pd�<�}<�Uy<��u<�q<�"n<�fj<��f<��b<3_<rx[<{�W<�T<hNP<K�L<G�H<�1E<�A<R�=<E):<<�6<�2<n:/<D�+<*(<�k$<�� <�L<��<�@<$�<�I<��<�i<[<K�<���;��;jZ�;W��;0\�;���;n��;rW�;�!�;^��;u�;��;$ �;�%�;�^�;���;�
�;s}�;��;�;�L�;
~;8�s;Кi;T�_;�U;;�K;cB;��8;k�/;.�&;�};c�;��;�?;1��:D��:�I�:Q�:���:�&�:&��:�!�:��k:��M:�0:1�:���9,�9��r9p�9!�7�.����G��Ù��FϹ,�a|���6��~P�43j�/������<*�����W'��V���,�̺t$ٺkY庫����������
������r��B�"��(��x.��\4�%<:�y@�R�E���K�7�Q�wW��J]�_c���h�ɾn���t�(`z����~ ���腻�ш�����פ��!����z���f���S���  �  �x=�=y�= ^=��=Ԡ=�A=�� =� =D# =K��<t��<��<�A�<�~�<��<v��<1�<�j�<`��<��<��< G�<n{�<���<G��<��<�?�<Nm�<P��<���<���<��<�8�<	\�<Y}�<���<Ϲ�<���<A��<q�<�<+(�<�6�<B�<�J�<QP�<�R�<R�<N�<�F�<z;�<�,�<]�<�<���<���<>��<���<�W�<R(�<���<*��<!�<\=�<���<���<�[�<��<$��<�N�<-��<��<��<(��<�-�<[��<�2�<,��<[%�<��<��<�p�<�ֱ<9�<?��<��<rH�<���<t�<8�<X��<�Ǣ<�
�<vK�<c��<�ě<���<�4�< i�<���<[̒<I��<�(�<CT�<�~�<i��<3χ<���<��<b@�<ud�<�}<�Uy<��u<�q<
#n<�fj<��f<��b<E3_<�x[<��W<�T<=NP<Y�L<-�H<�1E<߁A<P�=<A):<2�6<=�2<�:/<P�+<�(<�k$<�� <xL<��<a@<�<wI<��<�i<{<�<g��;��;FZ�;h��;!\�;���;}��;W�;�!�;f��;��;*�;3 �;�%�;�^�;/��;�
�;�}�;j�;ƞ�;M�;�~;��s;��i;{�_;��U;��K;�cB;��8;��/;D�&;�};��;��;�?;у�:P��:�G�:+�:H��::(�:��:"!�:��k:l�M:�0:��:!��9G*�9��r9�9��7P��)�G��Ù�oFϹJ*��x�U�6�/}P��5j����U����*�������'��������̺�"ٺ3X��� ���>����
����k�����ĩ"�˓(��y.�e\4��;:��@�K�E�	�K�-�Q�>wW��J]��c�c�h�T�n���t��_z����" ���腻�ш�������������wz���f��T���  �  �v=�=(�=u[=��=z�=!>=�� =�~ ={ =�{�<j��<��<5�<Bq�<���<I��<� �<�Y�<f��<��<���<*2�<ye�<j��<4��<���<e%�<�Q�<�|�<��<f��<'��<�<9�<)Y�<�v�<˒�<H��<���<I��<���<;��<�<B�<Y�<��<��<��<�<8�<� �<���<G��<���<T��<���<�g�<�?�<��<���<(��<
v�<z8�<E��<q��<�c�<��<���<e�<��<t��<�;�<���<�]�<��<�m�<��<k�<U�<;W�<Ǵ<w2�<��<���<f]�<p��<��<�f�<A��<��<�Q�<͙�<ߠ<�!�<ma�<���<�ٙ<V�<�H�<�}�<!��<�<.�<�=�<&j�<��<ξ�<p�<2�<�5�<\�<�}<�Ly<��u<��q<�%n<_mj<N�f<'�b<�E_<��[<��W<�#T<FpP<��L<
I<�_E<��A<�	><�b:<;6<�3<�/<��+<mO(<0�$< /!<��<� <#�<�&<ݱ<�B<��<iv<<���;���;J[�;��;�i�;��;���;�t�; E�;�%�;�;K�;�2�;\�;!��;��;�F�;���;C�;�݊;W��;jM�;�Dv;Pl;J	b;_$X;�dN;��D;T;;E2;.�(;��;��;�;�l;���:���:�a�:��:"�:1��:F�:�Ĉ:��r:��T:k�6:�D:a+�9�n�9wO�9��9��&8����2�쳏�M�Ź�������(?2��ML�Z2f�(������b������/��������_˺ʹ׺���;2�\���<�lE
�!I�5G��@��4"��$(�.� �3�u�9�V�?���E�łK��^Q��9W��]�Z�b��h�]�n��lt��Az���������ᅻ�̈�ʸ��6���[�������n���^���  �  �v=�="�=t[=��=x�=#>=�� =�~ =y =�{�<_��<��<5�<Mq�<���<;��<� �<�Y�<f��<#��<���<-2�<re�<~��<+��<���<]%�<�Q�<�|�<��<d��<3��<�<9�<Y�<w�<Ԓ�<W��<���<D��<���<#��<�<5�<f�<��<��<��<$�<K�<� �<���<5��<���<_��< ��<�g�<�?�<�<���<8��<"v�<~8�<D��<r��<�c�<��<���<e�<��<s��<�;�<��<�]�<��<wm�<��<#k�<a�<?W�<�ƴ<~2�<��<���<Z]�<b��<��<�f�<C��<��<�Q�<ә�<	ߠ<�!�<^a�<���<�ٙ<g�<�H�<y}�<!��< �<E�<�=�<+j�<��<ھ�<s�<%�<�5�<�[�<�}<�Ly<}�u<��q<�%n<hmj<�f<$�b<�E_<Ԏ[<��W<�#T<XpP<X�L<I<�_E<��A<
><�b:<־6<�3<�/<��+<fO(<�$</!<��<� <?�<�&<ұ<�B<��<�v<<���;���;�[�;���;�i�;��;4��;u�;�D�;�%�;A�;y�;�2�;�[�;>��;��;G�;S��;�B�;�݊;���;mM�;MDv;�l;p	b;J$X;�dN;��D;�T;;�2;T�(;*�;s�;�;m;���:v��:b�:!�:*�:���:ZF�:�Ĉ:��r:q�T:��6:�D:&�9�k�9O�9 �9H�&8s����2������Ź�������>2�[PL�l1f���ŵ��nc������ꄲ������_˺W�׺����1�\��=��E
��H��F�@��4"�%(�.�>�3���9���?�g�E�݂K��^Q�p9W�;]�^�b��h�*�n��lt�.Bz����q����ᅻ͈�и������������n���^���  �  �v=�= �=u[=��=u�=%>=� =�~ =w =|�<j��<��<5�<:q�<���<?��<� �<�Y�<a��<��<���<82�<he�<���<&��<���<r%�<�Q�<�|�<ץ�<g��<#��<�<9�<Y�<w�<���<\��<z��<O��<���<&��<%�<*�<l�<��<��<��<�<B�<� �< ��<9��<���<[��<���<�g�<�?�<�<���<1��<v�<r8�<H��<h��<�c�<��<˾�<e�<��<���<�;�<��<�]�<��<{m�<��<k�<N�<DW�<�ƴ<�2�<��<���<e]�<Z��<��<�f�<K��<{�<�Q�<Ι�<ߠ<�!�<aa�<Ş�<�ٙ<h�<�H�<�}�<6��<���<?�<�=�<+j�<��<ؾ�<v�<�<�5�<�[�<�}<�Ly<v�u<��q<�%n<{mj<)�f<7�b<�E_<Ŏ[<��W<�#T<|pP<L�L<4I<�_E<��A<
><�b:<޾6<�3<�/<��+<�O(<0�$</!<��<� <G�<�&<��<�B<y�<�v<�<���;���;�[�;���;�i�;�;%��;Vu�;�D�;�%�;�;\�;�2�;�[�;\��;g�;G�;8��;C�;ފ;��;�M�;�Cv;�l;*	b;]$X;�dN;��D;^T;;2;�(;Q�;��;�;�l;g��:���:�c�:Q�:��:���:�E�:ň:��r:8�T:!�6:�F:>(�9�n�9.S�9��9�'8<���2�����ՔŹ���Y���=2��QL�/f���������b��8���h���v���6_˺��׺���*2��[��x<��E
��H�WG�@��4"�3%(�l.�J�3���9���?�g�E��K��^Q�U9W��]���b�?�h���n��lt�KBz��������xᅻ�̈�����V���0���%����n���^���  �  �v=�=�=z[=��=y�=(>=�� =�~ =} = |�<c��<��<5�<Sq�<���<H��<� �<�Y�<m��<#��<���<=2�<ne�<z��<0��<���<b%�<�Q�<�|�<٥�<m��<��<�<9�<
Y�<w�<���<Q��<���<@��<���<"��<�<0�<n�<��<��<��<�<N�<� �<���<>��<���<c��<��<�g�<�?�<�<���<<��<!v�<�8�<M��<g��<�c�<��<���<e�<��<o��<�;�<��<�]�<��<nm�<�<k�<L�<EW�<�ƴ<z2�<���<���<[]�<e��<��<�f�<N��<��<�Q�<ٙ�<ߠ<�!�<ja�<Ş�<�ٙ<j�<�H�<}�<%��<�<J�<�=�<4j�<��<ξ�<�<�<�5�<�[�<�}<�Ly<��u<��q<�%n<fmj<�f<$�b<�E_<��[<��W<�#T<KpP<V�L<I<�_E<ǳA<
><�b:<�6<�3<�/<��+<uO(<!�$<(/!<��<� <H�<�&<۱<�B<��<�v<<Ј�;���;�[�;��;�i�;��;)��;�t�;�D�;�%�;��;\�;�2�;�[�;9��;o�;�F�;R��;�B�;�݊;���;}M�;/Dv;�l;	b;�$X;EeN;��D;�T;;z2;c�(;x�;��;!;:m;|��:��:Mb�:�:n�:���:�F�:pň:��r:"�T:Y�6:�D:&�9�j�9UN�9��9�&8���ٽ2����s�Ź�������=2�/QL��1f��������Wc��}������A����^˺��׺���1�[���<�E
��H��F��?��4"�Q%(��.���3���9�	�?�!�E���K��^Q�9W�u]�'�b��h�_�n��lt�Bz���������ᅻ&͈�и��D���L������	o���^���  �  �v=�= �=u[=��=�= >=�� =�~ =} =|�<n��<"��<5�<dq�<���<P��<� �<�Y�<e��<��<���<,2�<|e�<w��<,��<~��<a%�<�Q�<�|�<٥�<S��<��<�<9�<Y�<�v�<ɒ�<>��<{��<B��<���<.��<�<2�<`�<��<��<��<$�<<�<� �<���<P��<���<i��<��<�g�<�?�<�<���<+��<!v�<y8�<G��<q��<�c�<��<���<e�<��<p��<�;�<���<�]�<��<nm�<y�<k�<I�<+W�<�ƴ<x2�<��<���<W]�<c��<��<�f�<@��<��<�Q�<͙�<ߠ<�!�<ta�<���<�ٙ<g�<�H�<�}�<.��<�<;�<�=�<'j�<��<о�<s�<!�<�5�<\�<�}<�Ly<g�u<��q<�%n<Qmj<�f<�b<�E_<��[<��W<�#T<NpP<m�L<
I<�_E<��A<
><c:<ʾ6<�3<�/<��+<�O(<9�$<2/!<��<!<.�<�&<�<�B<��<�v<<���;��;�[�;���;�i�;��;^��;�t�;�D�;Y%�;��;N�;�2�;�[�;��;��;�F�;?��;�B�;�݊;'��;\M�;BDv;�l;M	b;�$X;�dN;��D;1T;;�2;��(;�;��;S;�m;���:��:�b�:x�:k�:���:F�:ň:��r:��T:`�6:D:�(�9Qm�9�N�9�9.�&8m����2�ͺ��Ź��������@2�@QL�2f����S����c������M���j����_˺��׺��32�G[���<�4E
�I�:F�@��4"��$(��.���3��9���?���E�t�K��^Q�r9W�Z]�\�b���h�P�n��lt��Bz��������ᅻ͈�����*�������Q����n���^���  �  �v=�=�=s[=��=|�='>=�� =�~ = =|�<n��</��<!5�<]q�<���<Z��<� �<�Y�<k��<$��<���<82�<se�<z��<&��<���<g%�<�Q�<�|�<ӥ�<\��<��<��<�8�<Y�<�v�<���<G��<y��<;��<{��<��<�<.�<c�<��<��<��<0�<E�<� �<���<J��<���<q��<��<�g�<�?�<�<���<5��<+v�<�8�<O��<l��<�c�<��<���<e�<��<g��<�;�<���<�]�<��<om�<s�<k�<K�<4W�<�ƴ<o2�<���<���<\]�<Z��<��<�f�<K��<��<�Q�<ՙ�<%ߠ<�!�<{a�<ʞ�<�ٙ<v�<
I�<�}�<9��<�<C�<�=�</j�<��<Ӿ�<r�<�<�5�<�[�<�}<vLy<k�u<��q<�%n<1mj<�f<��b<pE_<��[<��W<�#T<HpP<7�L<I<�_E<��A<
><c:<�6<�3<�/<��+<�O(<9�$<M/!<��<!<Q�<�&<�<�B<��<�v<-<���;���;�[�;���;�i�;��;���;�t�;�D�;�%�;��;�;�2�;�[�;Ж�;U�;�F�;7��;�B�;�݊;鋅;M�;!Dv;�l;F	b;�$X;0eN;�D;{T;;�2;��(;��;	�;�;�m;���:���:�b�:��:�:S��:�F�:�ň:F�r:
�T:��6:E: &�9Ei�9�L�9��9��&8r����2�q����Ź�������?2�RL�*3f����7���*c��)�����������)_˺ܳ׺��㺳1��Z���<��D
�zH�aF��?�4"��$(�X.���3���9���?�G�E���K��^Q�y9W�k]��b��h���n�/mt�vBz��������ⅻ͈�0�������k���?���o���^���  �  �v=�=�=y[=��=w�=)>=�� =�~ =� =|�<v��<3��<-5�<aq�<ͬ�<[��< !�<�Y�<t��</��<���<=2�<le�<���<+��<u��<c%�<�Q�<�|�<ʥ�<S��<��<��<�8�<�X�<�v�<���<;��<m��<6��<}��<��<�<$�<w�<��<��<��<)�<U�<� �<���<O��<���<t��<��<�g�<�?�<�<���<A��<(v�<�8�<M��<i��<�c�<��<���<�d�<��<e��<~;�<���<�]�<��<_m�<k�<	k�<9�<)W�<�ƴ<t2�<���<���<Q]�<[��<��<�f�<O��<��<�Q�<ߙ�<ߠ<�!�<{a�<מ�<�ٙ<~�<I�<�}�<<��<�<V�<�=�<6j�<��<׾�<��<�<�5�<�[�<�}<jLy<[�u<��q<�%n<>mj<��f<��b<vE_<��[<��W<�#T<TpP<3�L<I<�_E<ƳA<
><�b:<�6<�3<1�/<��+<�O(<I�$<T/!<ե<!<n�<�&<�<�B<��<�v<<؈�;���;�[�;���;ji�;��;��;�t�;lD�;^%�;��;�;�2�;`[�;���;>�;�F�;��;�B�;�݊;ދ�;M�;�Cv;Ml;1	b;�$X;6eN;��D;�T;;�2;�(;�;e�;�;�m;���:9��:�c�:��:��:#��:�F�:�ň:��r:��T:��6:�D:�$�9�i�9`L�9r�9�&8-(����2�[���ޛŹ������A2��RL�j2f�A�������c��������_����^˺7�׺9��1�[��=<��D
�H�;F�Q?��3"��$(�=.���3�7�9���?��E�˂K��^Q� 9W��]�+�b���h�G�n�]mt��Bz�#�������ᅻY͈����w�������\���Bo���^���  �  �v=�=�=t[=��=�=*>=�� =�~ =� =|�<���</��<)5�<sq�<Ŭ�<\��<!�<�Y�<z��<)��<���<?2�<{e�<w��<*��<|��<]%�<�Q�<�|�<ɥ�<O��<��<��<�8�<�X�<�v�<���<2��<s��<,��<y��< ��<�<)�<h�<��<��<��<%�<Q�<� �<
��<^��<���<~��<"��<�g�<@�<"�<���<A��<%v�<�8�<Q��<k��<�c�<��<���<e�<��<Z��<�;�<���<�]�<��<Ym�<f�<�j�<3�<"W�<�ƴ<b2�<���<���<V]�<]��<��<�f�<O��<��<�Q�<㙢<*ߠ<�!�<a�<Ξ�<�ٙ<~�<
I�<�}�<D��<�<P�<�=�<9j�<#��<о�<u�<�<�5�<�[�<�}<XLy<Y�u<��q<�%n<#mj<�f<��b<qE_<|�[<��W<�#T<3pP<D�L<
I<�_E<��A<
><c:<�6<�3<'�/< �+<�O(<e�$<M/!<Υ<?!<`�< '< �<�B<��<�v<$<���;
��;�[�;���;�i�;��;#��;�t�;lD�;P%�;��;�;q2�;O[�;ɖ�;A�;uF�;$��;�B�;�݊;�;oM�;�Cv;�l;,	b;�$X;seN;��D;�T;;�2;o�(;��;8�;�;;n;>��:���:Od�:,	�:��:��:G�:�ň:C�r:9�T:N�6:�D:�%�9�i�9�I�9�9�&8�*���2�����ٜŹ���j���A2��RL��4f�s��˵��c������J��������^˺�׺w���0�rZ���;��D
�WH��E�N?�4"�5$(��.�O�3�f�9���?���E�N�K��^Q�b9W��]�Z�b�O�h���n��mt��Bz�K������(ⅻg͈�R�����������j���Yo��_���  �  �v=�= �=s[=��=�='>=�� =�~ =� =|�<��<E��<65�<sq�<լ�<p��<!�<�Y�<���<0��<���<62�<}e�<v��<'��<}��<U%�<�Q�<�|�<ǥ�<E��<	��<��<�8�<�X�<�v�<���<*��<l��<#��<r��<��<�<1�<b�<��<��<��<<�<Z�<�<��<_��<���<���<"��<�g�<
@�<�<���<H��<8v�<�8�<I��<r��<�c�<��<���<�d�<��<N��<|;�<���<�]�<��<Wm�<\�<�j�<8�<W�<�ƴ<X2�<�<���<Q]�<]��<��<�f�<F��<��<�Q�<Ꙣ<*ߠ<�!�<�a�<ݞ�<�ٙ<��<I�<�}�<=��<#�<U�<>�<1j�<��<վ�<s�< �<�5�<�[�<�}<QLy<G�u<��q<r%n<mj<��f<��b<XE_<{�[<��W<�#T<'pP<:�L<�I<�_E<��A<
><c:<�6<�3<,�/<�+<�O(<\�$<y/!<�<?!<��<*'<�<�B<��<�v<V<�;��;�[�;���;�i�;��;��;�t�;eD�;+%�;��;��;;2�;\[�;{��;-�;XF�;��;xB�;�݊;ʋ�;FM�;EDv;�l;y	b;�$X;�eN;}�D;*U;;(2;)�(;��;��;;:n;0��:C��:�c�:o	�:Q�::��:�G�:Xň:2�r:��T:&�6:_C:#�9gg�9�F�9;�9��&8J+��@�2�տ��W�Ź�������B2�?SL��5f����Z����c������t���U���R_˺�׺���R0�`Z�� <�DD
��G��E�?�}3"�Z$(�8.�(�3�@�9���?�9�E�r�K��^Q�u9W�`]���b���h�חn��mt�Cz�Y�����hⅻL͈���������������do��1_���  �  �v=�=�=t[=��=~�=)>=�� =�~ =� =-|�<���<A��<@5�<mq�<��<f��<!�<�Y�<���<-��<���<>2�<ze�<���<$��<w��<b%�<�Q�<�|�<¥�<;��<���<��<�8�<�X�<�v�<���<&��<e��<0��<v��<��<�<$�<f�<��<��<��<-�<[�<�<��<_��<���<���<"��<�g�<@�<1�<���<G��<+v�<�8�<O��<r��<�c�<��<���<�d�<��<]��<t;�<���<�]�<��<Lm�<W�<�j�<%�<W�<�ƴ<i2�<꙱<���<Q]�<V��<��<�f�<N��<��<�Q�<虢<2ߠ<�!�<�a�<螛<�ٙ<��<I�<�}�<U��<#�<U�<�=�<4j�<��<۾�<u�<�<�5�<�[�<�}<\Ly<:�u<t�q<b%n<mj<ٴf<��b<KE_<g�[<z�W<�#T<6pP<)�L<I<�_E<��A<
><c:<�6<�3<+�/<�+<�O(<u�$<r/!<��<4!<��<'<1�<C<��<�v<?<߈�;	��;�[�;���;xi�;��;��;�t�;TD�;%�;n�;��;=2�;0[�;���;�;IF�;�;�B�;�݊;ʋ�;{M�;�Cv;�l;�	b;�$X;SeN;�D;2U;;62;��(;��;��;6;;n;���:+��:=e�:�	�:F�:f��:�F�:�ň:Y�r:�T:��6:oD:L$�9�g�9�J�9e�9��&899����2���e�Źt�����D2��SL��3f���������c��H������������^˺��׺5��g0��Y���;��D
��G��E��>�p3"�!$(�v.�&�3�:�9�j�?��E�i�K��^Q�^9W��]�1�b���h���n��mt�7Cz�u��3���9ⅻ�͈�h���ʥ��꒑�����]o��_���  �  �v=�=�=y[=��=��=1>=�� =�~ =� =&|�<���<<��<I5�<yq�<��<a��<!�<�Y�<���<D��<���<M2�<we�<|��<-��<p��<X%�<�Q�<�|�<���<O��<���<��<�8�<�X�<�v�<���<5��<`��<%��<g��<��<�<"�<p�<��<��<��<5�<q�<� �<��<`��<���<���<-��<�g�<@�<5�<���<\��<:v�<�8�<]��<g��<�c�<��<���<�d�<y�<S��<k;�<���<�]�<��<=m�<P�<�j�<"�<%W�<�ƴ<]2�<ؙ�<���<I]�<[��<��<�f�<^��<��<�Q�<���<+ߠ<�!�<�a�<�<�ٙ<��<I�<�}�<N��<$�<m�<�=�<Ej�<&��<Ѿ�<��<�<�5�<�[�<�}<BLy<@�u<��q<Q%n<mj<��f<��b<=E_<x�[<��W<�#T<"pP<�L<I<�_E<ĳA<	
><c:<�6<�3<\�/<�+<�O(<��$<j/!<�<M!<��<'<E�<�B<��<�v<6<��;���;�[�;��;]i�;��;���;�t�;D�;V%�;u�;��;02�;�Z�;���;��;�F�;ܺ�;�B�;p݊;���;hM�;�Cv; l;%	b;&%X;�eN;J�D;�U;;2;��(;��;��;�;�n;��:��:�e�:Q	�:��:Z��:�G�:�ƈ:��r:_�T:��6:�C:f �9�c�9UH�9�9)�&8�A��R�2�Ə��Ź5��T��-A2��UL��4f����Y���4d������Ą�������]˺��׺��㺓/�TZ��?;��D
�3G�rE�w>�s3"��#(��.��3�z�9�z�?���E�6�K��^Q�9W�]�R�b�1�h��n��mt�"Cz�E��T���9ⅻ�͈�i���祎�Ȓ�������o��;_���  �  �v=�=�=x[=��=��=&>=�� =�~ =� ='|�<���<L��<?5�<uq�<��<y��<!!�<�Y�<���<4��<���<72�<e�<w��<0��<p��<Y%�<�Q�<�|�<���<9��<���<��<�8�<�X�<�v�<���<"��<W��<*��<t��<��<�<+�<h�<��<��<��<2�<]�<�<��<s��<���<���<)��<�g�<@�</�<���<J��<0v�<�8�<L��<q��<�c�<��<���<�d�<��<X��<f;�<���<�]�<��<Gm�<R�<�j�<�<W�<�ƴ<d2�<�<���<G]�<b��<��<�f�<I��<��<�Q�<왢<1ߠ<�!�<�a�<ꞛ<�ٙ<��<'I�<�}�<M��<+�<Z�<>�</j�<"��<վ�<{�<�<�5�<�[�<�}<LLy<�u<l�q<J%n<mj<дf<��b<5E_<_�[<g�W<�#T<6pP<6�L<�I<�_E<��A<
><c:<�6<�3<7�/<"�+<�O(<��$<�/!<��<C!<��<<'<J�<C<��<�v<A<Ɉ�;"��;�[�;��;_i�;��;��;�t�;D�;�$�;U�;��;02�;[�;���;��;<F�;���;�B�;�݊;ڋ�;NM�;Dv;�l;h	b;�$X;GeN;2�D;JU;;`2;��(;1�;�;Y;yn;���:_��:'e�:�	�:x�:���:�F�:�ň:J�r:��T:��6:-C:�#�9�g�9�I�9��9E�&8>D����2��Ï�y�Ź'	�� �D2��UL�4f�������Vd��v���.���?���_˺��׺���0��Y��R;��C
�wG��E��>�*3"��#(��.���3��9�L�?�F�E�T�K��^Q�49W��]���b�}�h���n��mt��Cz����d���Gⅻ�͈�r�����������ـ��|o��_���  �  �v=�=�=o[=��=��='>=�� =�~ =� =-|�<���<B��<C5�<�q�<۬�<o��<!�<�Y�<���<0��<���<72�<�e�<r��<'��<s��<S%�<�Q�<||�<���<7��<��<��<�8�<�X�<�v�<���<$��<`��<"��<Y��<��<�<.�<U�<��<��<��<F�<X�<�<��<g��<���<���<;��<�g�<@�<$�<��<I��<?v�<�8�<Q��<���<�c�<��<���<�d�<p�<I��<m;�<���<�]�<��<<m�<E�<�j�<.�<
W�<�ƴ<Q2�<ܙ�<���<J]�<\��<��<�f�<I��<��<�Q�<�<Cߠ<�!�<�a�<㞛<�ٙ<��<I�<�}�<Q��<9�<Q�<>�<5j�</��<۾�<g�<�<�5�<�[�<o}<NLy</�u<y�q<`%n<�lj<��f<��b<EE_<r�[<q�W<�#T<�oP<�L<�I<�_E<��A<
><1c:<�6<+3<#�/<4�+<�O(<q�$<u/!<�<s!<��<)'<&�<C<��<�v<|<ʈ�;Z��;[�;���;ki�;��;���;qt�;ED�;�$�;��;��;�1�;�Z�;{��;�;CF�;޺�;wB�;:݊;���;KM�;0Dv;Jl;�	b;%X;�eN;��D;"U;;2;��(;��;��;�;o;���:���:vd�:&�:l�:���:H�:�ň:Q�r:��T:��6:'C:�"�9da�9�E�9N�9[�&8�2����2�8Ə���Źl������D2��TL�l6f�b��X���$d������Ӆ��]���'_˺��׺����/��X���;�AD
��G��D��>��3"��#(��.�p�3�]�9�i�?��E��K��^Q��9W�~]���b���h���n��mt�dCz�j��8����ⅻ�͈�����֥��Ւ��Ā��no���_���  �  �v=�=�=x[=��=��=&>=�� =�~ =� ='|�<���<L��<?5�<uq�<��<y��<!!�<�Y�<���<4��<���<72�<e�<w��<0��<p��<Y%�<�Q�<�|�<���<9��<���<��<�8�<�X�<�v�<���<"��<W��<*��<t��<��<�<+�<h�<��<��<��<2�<]�<�<��<s��<���<���<)��<�g�<@�</�<���<J��<0v�<�8�<L��<q��<�c�<��<���<�d�<��<X��<f;�<���<�]�<��<Gm�<R�<�j�<�<W�<�ƴ<d2�<�<���<G]�<b��<��<�f�<I��<��<�Q�<왢<1ߠ<�!�<�a�<ꞛ<�ٙ<��<'I�<�}�<M��<+�<Z�<>�</j�<"��<վ�<{�<�<�5�<�[�<�}<LLy<�u<l�q<J%n<mj<дf<��b<5E_<_�[<g�W<�#T<6pP<6�L<�I<�_E<��A<
><c:<�6<�3<7�/<"�+<�O(<��$<�/!<��<C!<��<<'<J�<C<��<�v<A<Ɉ�;"��;�[�;��;_i�;��;��;�t�;D�;�$�;U�;��;02�;[�;���;��;<F�;���;�B�;�݊;ڋ�;NM�;Dv;�l;h	b;�$X;GeN;2�D;JU;;`2;��(;1�;�;Y;yn;���:_��:'e�:�	�:x�:���:�F�:�ň:J�r:��T:��6:-C:�#�9�g�9�I�9��9E�&8>D����2��Ï�y�Ź'	�� �D2��UL�4f�������Vd��v���.���?���_˺��׺���0��Y��R;��C
�wG��E��>�*3"��#(��.���3��9�L�?�F�E�T�K��^Q�49W��]���b�}�h���n��mt��Cz����d���Gⅻ�͈�r�����������ـ��|o��_���  �  �v=�=�=y[=��=��=1>=�� =�~ =� =&|�<���<<��<I5�<yq�<��<a��<!�<�Y�<���<D��<���<M2�<we�<|��<-��<p��<X%�<�Q�<�|�<���<O��<���<��<�8�<�X�<�v�<���<5��<`��<%��<g��<��<�<"�<p�<��<��<��<5�<q�<� �<��<`��<���<���<-��<�g�<@�<5�<���<\��<:v�<�8�<]��<g��<�c�<��<���<�d�<y�<S��<k;�<���<�]�<��<=m�<P�<�j�<"�<%W�<�ƴ<]2�<ؙ�<���<I]�<[��<��<�f�<^��<��<�Q�<���<+ߠ<�!�<�a�<�<�ٙ<��<I�<�}�<N��<$�<m�<�=�<Ej�<&��<Ѿ�<��<�<�5�<�[�<�}<BLy<@�u<��q<Q%n<mj<��f<��b<=E_<x�[<��W<�#T<"pP<�L<I<�_E<ĳA<	
><c:<�6<�3<\�/<�+<�O(<��$<j/!<�<M!<��<'<E�<�B<��<�v<6<��;���;�[�;��;]i�;��;���;�t�;D�;V%�;u�;��;02�;�Z�;���;��;�F�;ܺ�;�B�;p݊;���;hM�;�Cv; l;%	b;&%X;�eN;J�D;�U;;2;��(;��;��;�;�n;��:��:�e�:Q	�:��:Z��:�G�:�ƈ:��r:_�T:��6:�C:f �9�c�9UH�9�9)�&8�A��R�2�Ə��Ź5��T��-A2��UL��4f����Y���4d������Ą�������]˺��׺��㺓/�TZ��?;��D
�3G�rE�w>�s3"��#(��.��3�z�9�z�?���E�6�K��^Q�9W�]�R�b�1�h��n��mt�"Cz�E��T���9ⅻ�͈�i���祎�Ȓ�������o��;_���  �  �v=�=�=t[=��=~�=)>=�� =�~ =� =-|�<���<A��<@5�<mq�<��<f��<!�<�Y�<���<-��<���<>2�<ze�<���<$��<w��<b%�<�Q�<�|�<¥�<;��<���<��<�8�<�X�<�v�<���<&��<e��<0��<v��<��<�<$�<f�<��<��<��<-�<[�<�<��<_��<���<���<"��<�g�<@�<1�<���<G��<+v�<�8�<O��<r��<�c�<��<���<�d�<��<]��<t;�<���<�]�<��<Lm�<W�<�j�<%�<W�<�ƴ<i2�<꙱<���<Q]�<V��<��<�f�<N��<��<�Q�<虢<2ߠ<�!�<�a�<螛<�ٙ<��<I�<�}�<U��<#�<U�<�=�<4j�<��<۾�<u�<�<�5�<�[�<�}<\Ly<:�u<t�q<b%n<mj<ٴf<��b<KE_<g�[<z�W<�#T<6pP<)�L<I<�_E<��A<
><c:<�6<�3<+�/<�+<�O(<u�$<r/!<��<4!<��<'<1�<C<��<�v<?<߈�;	��;�[�;���;xi�;��;��;�t�;TD�;%�;n�;��;=2�;0[�;���;�;IF�;�;�B�;�݊;ʋ�;{M�;�Cv;�l;�	b;�$X;SeN;�D;2U;;62;��(;��;��;6;;n;���:+��:=e�:�	�:F�:f��:�F�:�ň:Y�r:�T:��6:oD:L$�9�g�9�J�9e�9��&899����2���e�Źt�����D2��SL��3f���������c��H������������^˺��׺5��g0��Y���;��D
��G��E��>�p3"�!$(�v.�&�3�:�9�j�?��E�i�K��^Q�^9W��]�1�b���h���n��mt�7Cz�u��3���9ⅻ�͈�h���ʥ��꒑�����]o��_���  �  �v=�= �=s[=��=�='>=�� =�~ =� =|�<��<E��<65�<sq�<լ�<p��<!�<�Y�<���<0��<���<62�<}e�<v��<'��<}��<U%�<�Q�<�|�<ǥ�<E��<	��<��<�8�<�X�<�v�<���<*��<l��<#��<r��<��<�<1�<b�<��<��<��<<�<Z�<�<��<_��<���<���<"��<�g�<
@�<�<���<H��<8v�<�8�<I��<r��<�c�<��<���<�d�<��<N��<|;�<���<�]�<��<Wm�<\�<�j�<8�<W�<�ƴ<X2�<�<���<Q]�<]��<��<�f�<F��<��<�Q�<Ꙣ<*ߠ<�!�<�a�<ݞ�<�ٙ<��<I�<�}�<=��<#�<U�<>�<1j�<��<վ�<s�< �<�5�<�[�<�}<QLy<G�u<��q<r%n<mj<��f<��b<XE_<{�[<��W<�#T<'pP<:�L<�I<�_E<��A<
><c:<�6<�3<,�/<�+<�O(<\�$<y/!<�<?!<��<*'<�<�B<��<�v<V<�;��;�[�;���;�i�;��;��;�t�;eD�;+%�;��;��;;2�;\[�;{��;-�;XF�;��;xB�;�݊;ʋ�;FM�;EDv;�l;y	b;�$X;�eN;}�D;*U;;(2;)�(;��;��;;:n;0��:C��:�c�:o	�:Q�::��:�G�:Xň:2�r:��T:&�6:_C:#�9gg�9�F�9;�9��&8J+��@�2�տ��W�Ź�������B2�?SL��5f����Z����c������t���U���R_˺�׺���R0�`Z�� <�DD
��G��E�?�}3"�Z$(�8.�(�3�@�9���?�9�E�r�K��^Q�u9W�`]���b���h�חn��mt�Cz�Y�����hⅻL͈���������������do��1_���  �  �v=�=�=t[=��=�=*>=�� =�~ =� =|�<���</��<)5�<sq�<Ŭ�<\��<!�<�Y�<z��<)��<���<?2�<{e�<w��<*��<|��<]%�<�Q�<�|�<ɥ�<O��<��<��<�8�<�X�<�v�<���<2��<s��<,��<y��< ��<�<)�<h�<��<��<��<%�<Q�<� �<
��<^��<���<~��<"��<�g�<@�<"�<���<A��<%v�<�8�<Q��<k��<�c�<��<���<e�<��<Z��<�;�<���<�]�<��<Ym�<f�<�j�<3�<"W�<�ƴ<b2�<���<���<V]�<]��<��<�f�<O��<��<�Q�<㙢<*ߠ<�!�<a�<Ξ�<�ٙ<~�<
I�<�}�<D��<�<P�<�=�<9j�<#��<о�<u�<�<�5�<�[�<�}<XLy<Y�u<��q<�%n<#mj<�f<��b<qE_<|�[<��W<�#T<3pP<D�L<
I<�_E<��A<
><c:<�6<�3<'�/< �+<�O(<e�$<M/!<Υ<?!<`�< '< �<�B<��<�v<$<���;
��;�[�;���;�i�;��;#��;�t�;lD�;P%�;��;�;q2�;O[�;ɖ�;A�;uF�;$��;�B�;�݊;�;oM�;�Cv;�l;,	b;�$X;seN;��D;�T;;�2;o�(;��;8�;�;;n;>��:���:Od�:,	�:��:��:G�:�ň:C�r:9�T:N�6:�D:�%�9�i�9�I�9�9�&8�*���2�����ٜŹ���j���A2��RL��4f�s��˵��c������J��������^˺�׺w���0�rZ���;��D
�WH��E�N?�4"�5$(��.�O�3�f�9���?���E�N�K��^Q�b9W��]�Z�b�O�h���n��mt��Bz�K������(ⅻg͈�R�����������j���Yo��_���  �  �v=�=�=y[=��=w�=)>=�� =�~ =� =|�<v��<3��<-5�<aq�<ͬ�<[��< !�<�Y�<t��</��<���<=2�<le�<���<+��<u��<c%�<�Q�<�|�<ʥ�<S��<��<��<�8�<�X�<�v�<���<;��<m��<6��<}��<��<�<$�<w�<��<��<��<)�<U�<� �<���<O��<���<t��<��<�g�<�?�<�<���<A��<(v�<�8�<M��<i��<�c�<��<���<�d�<��<e��<~;�<���<�]�<��<_m�<k�<	k�<9�<)W�<�ƴ<t2�<���<���<Q]�<[��<��<�f�<O��<��<�Q�<ߙ�<ߠ<�!�<{a�<מ�<�ٙ<~�<I�<�}�<<��<�<V�<�=�<6j�<��<׾�<��<�<�5�<�[�<�}<jLy<[�u<��q<�%n<>mj<��f<��b<vE_<��[<��W<�#T<TpP<3�L<I<�_E<ƳA<
><�b:<�6<�3<1�/<��+<�O(<I�$<T/!<ե<!<n�<�&<�<�B<��<�v<<؈�;���;�[�;���;ji�;��;��;�t�;lD�;^%�;��;�;�2�;`[�;���;>�;�F�;��;�B�;�݊;ދ�;M�;�Cv;Ml;1	b;�$X;6eN;��D;�T;;�2;�(;�;e�;�;�m;���:9��:�c�:��:��:#��:�F�:�ň:��r:��T:��6:�D:�$�9�i�9`L�9r�9�&8-(����2�[���ޛŹ������A2��RL�j2f�A�������c��������_����^˺7�׺9��1�[��=<��D
�H�;F�Q?��3"��$(�=.���3�7�9���?��E�˂K��^Q� 9W��]�+�b���h�G�n�]mt��Bz�#�������ᅻY͈����w�������\���Bo���^���  �  �v=�=�=s[=��=|�='>=�� =�~ = =|�<n��</��<!5�<]q�<���<Z��<� �<�Y�<k��<$��<���<82�<se�<z��<&��<���<g%�<�Q�<�|�<ӥ�<\��<��<��<�8�<Y�<�v�<���<G��<y��<;��<{��<��<�<.�<c�<��<��<��<0�<E�<� �<���<J��<���<q��<��<�g�<�?�<�<���<5��<+v�<�8�<O��<l��<�c�<��<���<e�<��<g��<�;�<���<�]�<��<om�<s�<k�<K�<4W�<�ƴ<o2�<���<���<\]�<Z��<��<�f�<K��<��<�Q�<ՙ�<%ߠ<�!�<{a�<ʞ�<�ٙ<v�<
I�<�}�<9��<�<C�<�=�</j�<��<Ӿ�<r�<�<�5�<�[�<�}<vLy<k�u<��q<�%n<1mj<�f<��b<pE_<��[<��W<�#T<HpP<7�L<I<�_E<��A<
><c:<�6<�3<�/<��+<�O(<9�$<M/!<��<!<Q�<�&<�<�B<��<�v<-<���;���;�[�;���;�i�;��;���;�t�;�D�;�%�;��;�;�2�;�[�;Ж�;U�;�F�;7��;�B�;�݊;鋅;M�;!Dv;�l;F	b;�$X;0eN;�D;{T;;�2;��(;��;	�;�;�m;���:���:�b�:��:�:S��:�F�:�ň:F�r:
�T:��6:E: &�9Ei�9�L�9��9��&8r����2�q����Ź�������?2�RL�*3f����7���*c��)�����������)_˺ܳ׺��㺳1��Z���<��D
�zH�aF��?�4"��$(�X.���3���9���?�G�E���K��^Q�y9W�k]��b��h���n�/mt�vBz��������ⅻ͈�0�������k���?���o���^���  �  �v=�= �=u[=��=�= >=�� =�~ =} =|�<n��<"��<5�<dq�<���<P��<� �<�Y�<e��<��<���<,2�<|e�<w��<,��<~��<a%�<�Q�<�|�<٥�<S��<��<�<9�<Y�<�v�<ɒ�<>��<{��<B��<���<.��<�<2�<`�<��<��<��<$�<<�<� �<���<P��<���<i��<��<�g�<�?�<�<���<+��<!v�<y8�<G��<q��<�c�<��<���<e�<��<p��<�;�<���<�]�<��<nm�<y�<k�<I�<+W�<�ƴ<x2�<��<���<W]�<c��<��<�f�<@��<��<�Q�<͙�<ߠ<�!�<ta�<���<�ٙ<g�<�H�<�}�<.��<�<;�<�=�<'j�<��<о�<s�<!�<�5�<\�<�}<�Ly<g�u<��q<�%n<Qmj<�f<�b<�E_<��[<��W<�#T<NpP<m�L<
I<�_E<��A<
><c:<ʾ6<�3<�/<��+<�O(<9�$<2/!<��<!<.�<�&<�<�B<��<�v<<���;��;�[�;���;�i�;��;^��;�t�;�D�;Y%�;��;N�;�2�;�[�;��;��;�F�;?��;�B�;�݊;'��;\M�;BDv;�l;M	b;�$X;�dN;��D;1T;;�2;��(;�;��;S;�m;���:��:�b�:x�:k�:���:F�:ň:��r:��T:`�6:D:�(�9Qm�9�N�9�9.�&8m����2�ͺ��Ź��������@2�@QL�2f����S����c������M���j����_˺��׺��32�G[���<�4E
�I�:F�@��4"��$(��.���3��9���?���E�t�K��^Q�r9W�Z]�\�b���h�P�n��lt��Bz��������ᅻ͈�����*�������Q����n���^���  �  �v=�=�=z[=��=y�=(>=�� =�~ =} = |�<c��<��<5�<Sq�<���<H��<� �<�Y�<m��<#��<���<=2�<ne�<z��<0��<���<b%�<�Q�<�|�<٥�<m��<��<�<9�<
Y�<w�<���<Q��<���<@��<���<"��<�<0�<n�<��<��<��<�<N�<� �<���<>��<���<c��<��<�g�<�?�<�<���<<��<!v�<�8�<M��<g��<�c�<��<���<e�<��<o��<�;�<��<�]�<��<nm�<�<k�<L�<EW�<�ƴ<z2�<���<���<[]�<e��<��<�f�<N��<��<�Q�<ٙ�<ߠ<�!�<ja�<Ş�<�ٙ<j�<�H�<}�<%��<�<J�<�=�<4j�<��<ξ�<�<�<�5�<�[�<�}<�Ly<��u<��q<�%n<fmj<�f<$�b<�E_<��[<��W<�#T<KpP<V�L<I<�_E<ǳA<
><�b:<�6<�3<�/<��+<uO(<!�$<(/!<��<� <H�<�&<۱<�B<��<�v<<Ј�;���;�[�;��;�i�;��;)��;�t�;�D�;�%�;��;\�;�2�;�[�;9��;o�;�F�;R��;�B�;�݊;���;}M�;/Dv;�l;	b;�$X;EeN;��D;�T;;z2;c�(;x�;��;!;:m;|��:��:Mb�:�:n�:���:�F�:pň:��r:"�T:Y�6:�D:&�9�j�9UN�9��9�&8���ٽ2����s�Ź�������=2�/QL��1f��������Wc��}������A����^˺��׺���1�[���<�E
��H��F��?��4"�Q%(��.���3���9�	�?�!�E���K��^Q�9W�u]�'�b��h�_�n��lt�Bz���������ᅻ&͈�и��D���L������	o���^���  �  �v=�= �=u[=��=u�=%>=� =�~ =w =|�<j��<��<5�<:q�<���<?��<� �<�Y�<a��<��<���<82�<he�<���<&��<���<r%�<�Q�<�|�<ץ�<g��<#��<�<9�<Y�<w�<���<\��<z��<O��<���<&��<%�<*�<l�<��<��<��<�<B�<� �< ��<9��<���<[��<���<�g�<�?�<�<���<1��<v�<r8�<H��<h��<�c�<��<˾�<e�<��<���<�;�<��<�]�<��<{m�<��<k�<N�<DW�<�ƴ<�2�<��<���<e]�<Z��<��<�f�<K��<{�<�Q�<Ι�<ߠ<�!�<aa�<Ş�<�ٙ<h�<�H�<�}�<6��<���<?�<�=�<+j�<��<ؾ�<v�<�<�5�<�[�<�}<�Ly<v�u<��q<�%n<{mj<)�f<7�b<�E_<Ŏ[<��W<�#T<|pP<L�L<4I<�_E<��A<
><�b:<޾6<�3<�/<��+<�O(<0�$</!<��<� <G�<�&<��<�B<y�<�v<�<���;���;�[�;���;�i�;�;%��;Vu�;�D�;�%�;�;\�;�2�;�[�;\��;g�;G�;8��;C�;ފ;��;�M�;�Cv;�l;*	b;]$X;�dN;��D;^T;;2;�(;Q�;��;�;�l;g��:���:�c�:Q�:��:���:�E�:ň:��r:8�T:!�6:�F:>(�9�n�9.S�9��9�'8<���2�����ՔŹ���Y���=2��QL�/f���������b��8���h���v���6_˺��׺���*2��[��x<��E
��H�WG�@��4"�3%(�l.�J�3���9���?�g�E��K��^Q�U9W��]���b�?�h���n��lt�KBz��������xᅻ�̈�����V���0���%����n���^���  �  �v=�="�=t[=��=x�=#>=�� =�~ =y =�{�<_��<��<5�<Mq�<���<;��<� �<�Y�<f��<#��<���<-2�<re�<~��<+��<���<]%�<�Q�<�|�<��<d��<3��<�<9�<Y�<w�<Ԓ�<W��<���<D��<���<#��<�<5�<f�<��<��<��<$�<K�<� �<���<5��<���<_��< ��<�g�<�?�<�<���<8��<"v�<~8�<D��<r��<�c�<��<���<e�<��<s��<�;�<��<�]�<��<wm�<��<#k�<a�<?W�<�ƴ<~2�<��<���<Z]�<b��<��<�f�<C��<��<�Q�<ә�<	ߠ<�!�<^a�<���<�ٙ<g�<�H�<y}�<!��< �<E�<�=�<+j�<��<ھ�<s�<%�<�5�<�[�<�}<�Ly<}�u<��q<�%n<hmj<�f<$�b<�E_<Ԏ[<��W<�#T<XpP<X�L<I<�_E<��A<
><�b:<־6<�3<�/<��+<fO(<�$</!<��<� <?�<�&<ұ<�B<��<�v<<���;���;�[�;���;�i�;��;4��;u�;�D�;�%�;A�;y�;�2�;�[�;>��;��;G�;S��;�B�;�݊;���;mM�;MDv;�l;p	b;J$X;�dN;��D;�T;;�2;T�(;*�;s�;�;m;���:v��:b�:!�:*�:���:ZF�:�Ĉ:��r:q�T:��6:�D:&�9�k�9O�9 �9H�&8s����2������Ź�������>2�[PL�l1f���ŵ��nc������ꄲ������_˺W�׺����1�\��=��E
��H��F�@��4"�%(�.�>�3���9���?�g�E�݂K��^Q�p9W�;]�^�b��h�*�n��lt�.Bz����q����ᅻ͈�и������������n���^���  �  Ou=�=�=�X=��=C�=�:=�� =ez =� =r�<���<���<�(�<Rd�<��<���<{�<`I�<2��<���<���<(�<�P�<r��<"��<z��<D�<�7�<Ba�<n��<ï�<[��<��<��<�6�<@S�<�m�<���<��<R��<:��<���<��<���<���<���<X��<���<3��<��<���<N��<n��<Ԋ�<Sn�<�M�<{)�<� �<3��<<��<�m�<'4�<��<K��<l�<@ �<���<�z�<>!�<���<�_�<y��<K��<��<W��<�,�<���< ,�<?��<5�<��<���<�`�<�ů<�&�<D��<5ު<�4�<懧<�ץ<�$�<�n�<���<���<�;�<�z�<z��<�<z*�<�`�<e��<*Ȑ<0��<�(�<�V�<���<F��<�م<`�<�+�<�S�<\�|<Dy<��u<��q<R(n<�sj<e�f<�
c<W_<�[<��W<�@T<��P<�L<�5I<`�E<��A<�<><��:<9�6<�[3<��/<y+,<Ϙ(<
%<�!<��<�x<��<�<v<Ҩ<�B	<U�<F�<o�;���;-N�;r��;�g�;g�;'��;T��;�V�;�;�;W2�;&:�;�S�;��;q��;�;�p�;��;o�;f
�;���;�y�;�x;�gn;�Zd;�qZ;�P;"G;ܑ=;�94;�+;��!;��;,;{;���:���:�B�:T��:���:���:�ϛ:�6�:��y:^4[:�&=:=q:�:��9{��9`y/9�{8O.B�����%���Y��q򹈮��.�UH��_b�;4|���������f]��O����{����ɺlUֺ��⺙���*�������	�������[��(�!�=�'�ٮ-�Н3�5�9��r?�YE��<K��Q���V�]�\��b�,�h�*qn�0Kt��%z� ��;킻�څ�+Ȉ�˶������'��������v��ai���  �  Hu=�=�=�X=��=B�=�:=�� =jz =� =r�<¯�<���<�(�<bd�<���<���<��<\I�<7��<���<���<*�<yP�<���<+��<v��<B�<�7�<Sa�<m��<���<W��<��<��<�6�<AS�<�m�<���<���<Q��<9��<���<��<���<���<���<[��<���<3��<��<y��<T��<q��<֊�<bn�<�M�<�)�<� �<;��<2��<�m�<(4�<���<L��<l�<R �<���<�z�<4!�<���<�_�<u��<H��<��<[��<�,�<|��<,�<9��<0�<��<���<�`�<�ů<�&�<M��<Iު<�4�<燧<�ץ<�$�<�n�<���<���<�;�<�z�<���<�<v*�<�`�<f��<Ȑ<<��<�(�<�V�<���<Q��<�م<b�< ,�<�S�<t�|<�Cy<��u<��q<N(n<�sj<�f<�
c<W_<�[<��W<�@T<��P<e�L<�5I<Y�E<��A<=><��:<5�6<�[3<��/<l+,<̘(<)
%<�!<�<�x<��<�<�<ɨ<C	<b�<%�<o�;���;|N�;���;�g�;a�;��;���;�V�;�;�;J2�;9:�;�S�;\�;v��;��;�p�;��;o�;a
�;���;�y�;,�x;Ahn;�Zd;�qZ;�P; G;X�=;b94;�+;��!;��;�,;|{;,��:���:AC�:���:���:���:ϛ:�6�:<�y:�6[:_'=:�q:F:!�9|��9w/9x�{8�?B�x��V,��^�� �9��4.�QUH��]b��5|�����Ű���\�����D|����ɺoVֺ�����K+����z�	�z�������D�!��'�̮-�*�3�։9��r?�YE��<K�<Q�B�V�Q�\�͹b���h��pn�NKt��%z� ��E킻�څ��Ȉ�䶋�����&��������v��&i���  �  Fu=�=�=�X=��=@�=�:=�� =oz =� =r�<ǯ�<���<�(�<Sd�<��<���<��<TI�<5��<��<���<<�<pP�<���<!��<r��<Q�<�7�<Wa�<b��<ǯ�<Q��<��<��<�6�<OS�<�m�<���<ޛ�<L��<=��<���<!��<���<���<���<`��<���<0��<!��<q��<W��<r��<Ҋ�<[n�<�M�<~)�<� �<;��<'��<�m�<$4�<���<U��<l�<S �<���<�z�<8!�<���<�_�<o��<N��<��<e��<�,�<���<,�<3��<7�<��<���<�`�<�ů<�&�<C��<Hު<�4�<���<�ץ<�$�<�n�<���<���<�;�<�z�<z��<�<p*�<�`�<h��<Ȑ<E��<�(�<�V�<���<M��<�م<T�<,�<�S�<��|<�Cy<��u<��q<5(n<�sj<$�f<c<W_<�[<��W<w@T<��P<]�L<�5I<C�E<��A<=><��:<S�6<�[3<��/<b+,<ɘ(<3
%<�!<��<�x<��<�<�<��<C	<s�<%�<ao�;���;xN�;p��;�g�;��;��;���;�V�;�;�;22�;*:�;�S�;~�;���;��;�p�;��;o�;r
�;���;�y�;Śx;1hn;sZd;rZ;�P;G;��=;"94;�+;��!;��;U,;"{;���:���:OC�:��:Û�:~��:Mϛ:�7�:X�y:�6[:�%=:�r:�:��90��9Rt/9��{8mSB�m��q*��[�������h.�VH�]b�.6|����ɰ��s]������|����ɺHVֺK�����+��y����	�������%��t�!���'���-�X�3���9��r?��XE��<K�\Q�r�V���\�_�b���h��pn��Kt��%z� ��v킻�څ��Ȉ�����¥��7��������v��i���  �  Hu=�=�=�X=��=>�=�:=�� =kz =� =r�<ǯ�<���<�(�<ad�<���<���<��<^I�<2��<��<���</�<tP�<z��<'��<v��<F�<�7�<Ga�<a��<ʯ�<T��<���<��<�6�<8S�<�m�<���<���<G��<8��<���<��<���<���<���<S��<���<7��<��<���<L��<y��<���<en�<�M�<�)�<� �<2��<8��<�m�<)4�<��<H��<l�<K �<���<�z�<4!�<���<�_�<p��<M��<��<O��<�,�<��<�+�<4��<8�<��<���<�`�<�ů<�&�<I��<<ު<�4�<뇧<�ץ<�$�<�n�<���<���<�;�<�z�<���<�<�*�<�`�<c��<'Ȑ<:��<�(�<�V�<���<J��<�م<X�<,�<�S�<i�|<�Cy<��u<��q<.(n<�sj<*�f<�
c<�V_<�[<��W<u@T<��P<b�L<�5I<L�E<��A<�<><��:<E�6<�[3<��/<t+,<ɘ(<3
%<�!<�<�x<��<�<�<Ϩ<�B	<o�<:�<-o�;���;PN�;���;�g�;s�;��;m��;�V�;
<�;>2�;�9�;�S�;{�;T��;��;�p�;��;�n�;_
�;���;�y�;�x;$hn;�Zd;�qZ;-�P;>G;&�=;�94;�+;	�!;�;�,;~{;���:~��:�B�:��:&��:˚�:�ϛ:�6�:(�y:�5[:�&=:�q:<:�99u/9��{8FOB�_��+��8]����̯�9.��VH�_b�'6|�����ʰ��]������H|��l�ɺ�Uֺ?�⺄���*������	�j��&�������!��'��-��3��9��r?��XE�=K�rQ�R�V���\���b���h��pn��Kt��%z� ���킻�څ��Ȉ�붋�륎�3���o����v��Gi���  �  Iu=�=�=�X=��=G�=�:=�� =gz =� =%r�<ʯ�<���<�(�<id�<��<���<��<mI�<9��<���<���<)�<�P�<{��<-��<u��<9�<�7�<Oa�<j��<���<U��<��<��<�6�<:S�<�m�<��<ڛ�<I��<9��<���<��<���<���<���<\��<���<;��<��<���<Q��<���<ڊ�<^n�<�M�<�)�<�<8��<F��<�m�<,4�<���<L��<$l�<H �<���<�z�<.!�<���<�_�<p��<;��<��<T��<�,�<|��<�+�<5��<"�<��<���<�`�<�ů<�&�<Q��<<ު<�4�<燧<�ץ<�$�<�n�<���<���<�;�<�z�<���<
�<�*�<�`�<k��<1Ȑ<3��<�(�<�V�<���<P��<�م<_�<�+�<�S�<s�|<�Cy<��u<��q<N(n<�sj<&�f<�
c<W_<�[<��W<�@T<��P<g�L<�5I<T�E<��A<=><��:<3�6<�[3<��/<�+,<ߘ(<:
%<�!<��<y<��<�<�<�<C	<d�<8�<o�;���;SN�;���;�g�;>�;��;���;�V�;�;�;C2�;$:�;�S�;{�;^��;��;�p�;��;�n�;b
�;���;zy�;K�x;hn;�Zd;�qZ;�P;cG;�=;
:4;�+;Z�!;��;r,;g{;M��:"��:C�:���:<��:��:Rϛ:7�:��y:�5[:+(=:�p:�:r�9�9!u/9�m{8�?B�}���*���]���򹢯��.��UH�I^b�|5|�������\������O{����ɺ�Uֺu��,��*��{���	�������.����!���'���-���3��9��r?�YE��<K�GQ�U�V�i�\��b���h��pn��Kt�&z�7 ��D킻�څ��Ȉ�	�������G��������v��2i���  �  Cu=�=�=�X=��=E�=�:=�� =qz =� =&r�<ʯ�<���<�(�<id�< ��<���<��<dI�<C��<��<���<:�<xP�<}��<$��<r��<J�<�7�<Ja�<^��<���<K��<��<��<�6�<=S�<�m�<��<՛�<C��<5��<���<��<���<���<���<k��<���<;��<*��<���<Y��<���<��<in�<�M�<�)�< �<?��<;��<�m�</4�<���<\��<l�<K �<���<�z�<3!�<���<�_�<g��<@��<��<S��<�,�<n��<�+�<)��<)�<��<���<�`�<�ů<�&�<E��<?ު<�4�<���<�ץ<�$�<�n�<���<���<�;�<�z�<���<�<�*�<�`�<p��<+Ȑ<K��<�(�<�V�<���<H��<�م<W�<,�<�S�<m�|<�Cy<��u<��q<-(n<�sj<�f<�
c<�V_<ԣ[<��W<j@T<��P<Q�L<�5I<J�E<��A<�<><��:<J�6<�[3<�/<�+,<��(<9
%<�!<�<y<��<�<�<ܨ<!C	<��<5�<\o�;���;\N�;~��;�g�;��;Ծ�;}��;�V�;�;�;2�;:�;�S�;D�;h��;��;�p�;r�;�n�;R
�;���;�y�;	�x;hn;jZd;erZ;�P;fG;ϒ=;�94;�+;K�!;-�;�,;�{;��:���:�C�:G��:z��:=��:>ϛ:8�:t�y:�5[:'=:�q:T:��9���9�p/99z{8z`B�����.��"a��I����.��VH��^b��6|���������F]������b|����ɺVֺȪ�8���*��P���	�#����������!���'��-�͝3�W�9��r?��XE�{<K��Q�u�V���\���b�Еh��pn��Kt�&z�C ���킻�څ��Ȉ����Х��^��������v��>i���  �  =u=�=ܷ=�X=��=A�=�:=�� =sz =� =.r�<ѯ�<���<)�<dd�<��<���<��<iI�<?��<��<���<>�<pP�<���<%��<n��<C�<�7�<Pa�<O��<���<A��< ��<��<~6�<9S�<�m�<���<ț�<G��<0��<r��<��<���<���<���<g��<���<4��<*��<���<e��<|��<��<ln�<�M�<�)�<� �<L��<9��<�m�<+4�<���<Y��<l�<Z �<���<�z�<'!�<���<�_�<Y��<C��<z�<O��<�,�<n��<�+�<��<*�<�<���<�`�<�ů<�&�<?��<Mު<�4�<���<�ץ<�$�<�n�<���<���<�;�<�z�<���<!�<�*�<�`�<x��<%Ȑ<M��<�(�<�V�<���<L��<�م<J�<
,�<�S�<m�|<�Cy<��u<��q<(n<�sj<��f<�
c<�V_<ɣ[<��W<[@T<��P<8�L<�5I<3�E<��A<=><��:<Z�6<�[3<�/<z+,<�(<H
%<�!<*�<�x<��<�<�<�<C	<��<'�<oo�;���;�N�;���;�g�;j�;���;���;vV�;�;�;�1�;�9�;�S�;&�;\��;��;�p�;A�;�n�;B
�;O��;�y�;~�x;�hn;\Zd;JrZ;�P;3G;Ւ=;�94;W+;&�!;{�;�,;�{;���:���:cD�:0��:���:���:Lϛ:�7�:נy:�7[:�$=:�q:�:�9���9j/9��{8�yB����0���`��u�q���.�YH�^b��8|�,������]�������|��w�ɺuVֺĪ�Y�*��ت�$�	������w����!���'�:�-���3�L�9��r?��XE��<K�aQ���V��\�{�b�@�h��pn��Kt�B&z�M ���킻�څ� Ɉ����󥎻t�������w��0i���  �  Bu=�=�=�X=��=F�=�:=�� =qz =� =-r�<د�<���<)�<od�<��<���<��<pI�<A��<��<���<;�<~P�<y��<$��<v��<=�<�7�<Oa�<T��<���<A��<���<��<�6�<.S�<�m�<��<Ǜ�<H��<0��<x��<��<���<���<���<e��<���<A��<$��<���<c��<���<��<ln�<N�<�)�<�<I��<G��<�m�<34�<��<X��<l�<J �<���<�z�<(!�<���<�_�<Y��<5��<��<E��<�,�<i��<�+�< ��<�<���<���<�`�<�ů<�&�<@��<;ު<�4�<���<�ץ<�$�<�n�<���<���<�;�<�z�<���< �<�*�<�`�<v��<3Ȑ<F��<�(�<�V�<���<G��<�م<R�<,�<�S�<f�|<�Cy<u�u<p�q<"(n<�sj<�f<�
c<�V_<��[<��W<f@T<��P<J�L<�5I<B�E<��A<�<><��:<]�6<�[3<�/<�+,<�(<V
%<	�!<*�<y<�<�<�<��<C	<��<E�<fo�;���;QN�;���;�g�;U�;ľ�;���;�V�;�;�;�1�;�9�;{S�;7�;3��;��;�p�;@�;�n�;E
�;h��;�y�;��x;-hn;�Zd;?rZ;\�P;�G;��=;-:4;I+;��!;��;�,;�{;���:e��::D�:��:0��:���:�ϛ:�7�:��y:�5[:�%=:r::��9ؕ�9jj/9hf{8�lB�o���/��)b������M.��XH�^b��7|�|񊺠����]�������{����ɺ�Uֺ���w���)����̺	����������Z�!�b�'�L�-���3���9��r?�|XE��<K��Q�b�V���\���b���h�qn��Kt�r&z�} ���킻*ۅ��Ȉ�9���񥎻����΅��w��Di���  �  Cu=�=�=�X=��=H�=�:=�� =sz =� =,r�<ޯ�<���<)�<yd�<��<���<��<qI�<K��<��<���<+�<�P�<|��<.��<m��<9�<�7�<7a�<[��<���<B��<���<��<~6�< S�<�m�<���<ӛ�<7��<'��<y��<
��<���<���<���<b��<���<J��<(��<���<\��<���<��<{n�<N�<�)�<�<B��<P��<�m�<;4�<���<Q��<$l�<G �<���<�z�<)!�<���<�_�<d��<.��<��<6��<�,�<\��<�+�<"��<�<���<���<�`�<�ů<�&�<O��<<ު<�4�<釧<�ץ<�$�<�n�<���<���<�;�<�z�<���<&�<�*�<�`�<s��<?Ȑ<K��<�(�<�V�<���<P��<�م<^�<�+�<�S�<G�|<�Cy<��u<l�q<"(n<lsj<�f<�
c<�V_<��[<��W<e@T<z�P<N�L<�5I<P�E<��A<=><Ù:<7�6<\3<	�/<�+,<�(<d
%<�!</�<'y<��<;�<�<��<2C	<��<R�<(o�;���;aN�;���;�g�;F�;о�;3��;�V�;�;�; 2�;�9�;GS�;+�;���;��;yp�;r�;�n�;!
�;m��;ky�;F�x;hn;�Zd;(rZ;��P;�G;ǒ=;z:4;+;��!;��;c-;L|;��:`��:�C�:���:x��:���:kϛ:y7�:أy:�5[:(=:�o:3:�
�92��98p/9�W{8IhB�b�c1��e��򹹱�8 .�yWH�ab�_7|��񊺉����\������={��h�ɺ_UֺI������)����@�	����Z��N��-�!��'�c�-�&�3�Y�9�r?�YE�n<K�HQ�_�V�n�\�)�b��h��qn�Lt�>&z�� ���킻`ۅ��Ȉ�n�����������ȅ��w���i���  �  Cu=�=۷=�X=��=G�=�:=�� =pz =� =>r�<��<���<)�<{d�<��<���<��<{I�<F��<��<���<9�<P�<|��<'��<`��<@�<�7�<<a�<Q��<���<;��<���<��<{6�<%S�<�m�<ۅ�<ě�<3��<)��<}��<��<���<���<���<h��<���<E��<"��<���<o��<���<��<|n�<N�<�)�<�<T��<N��<�m�<84�<��<Y��<l�<I �<���<�z�<.!�<���<�_�<U��<'��<y�<<��<�,�<e��<�+�<��<�<�<���<�`�<�ů<�&�<E��<=ު<�4�<���<�ץ<�$�<�n�<���<��<�;�<�z�<���<,�<�*�<�`�<���<6Ȑ<D��<�(�<�V�<���<K��<�م<L�<�+�<�S�<T�|<�Cy<f�u<f�q<(n<ysj<��f<�
c<�V_<��[<p�W<Q@T<��P<P�L<�5I</�E<��A<�<><��:<R�6<\3<��/<�+,<�(<j
%<�!<>�<,y<�<�<�<�<)C	<��<P�<_o�;���;cN�;���;�g�;c�;���;L��;�V�;z;�;�1�;�9�;pS�;�;��;��;hp�;6�;�n�;+
�;|��;wy�;՚x;hn;�Zd;ZrZ;\�P;�G;��=;L:4;�+;��!;[�;l-;F|;���:���:�D�:���:*��:֛�:�ϛ:�7�:^�y:�5[:g&=:�o:�:�	�9���9�h/95L{8MzB�v�=1���b������� .��XH��`b�8|��-��� ]�������{����ɺTUֺd��3��N)�������	����S������!��'���-�o�3���9�Kr?��XE�n<K�nQ�j�V���\��b��h�Kqn�LLt��&z�� ���킻Dۅ�Ɉ�O��������������0w��mi���  �  =u=�=۷=�X=��=D�=�:=�� =wz =� =8r�<��<���<)�<yd�<$��<���<��<xI�<I��<��<���<B�<{P�<{��<(��<j��<B�<�7�<Ia�<C��<���<7��<���<��<l6�<S�<�m�<���<���<:��<'��<u��<��<���<���<���<j��<��<F��<1��<���<n��<���<���<�n�<N�<�)�<�<T��<M��<�m�<:4�<
��<]��<l�<R �<���<�z�<&!�<���<�_�<E��</��<o�<3��<x,�<Z��<�+�<��<�<ኴ<���<�`�<�ů<�&�<B��<<ު<�4�<���<�ץ<�$�<�n�<���<��<�;�<�z�<���<;�<�*�<�`�<���<7Ȑ<S��<�(�<�V�<���<E��<�م<I�<,�<�S�<\�|<�Cy<V�u<k�q<�'n<nsj<׾f<�
c<�V_<��[<k�W<D@T<��P<5�L<�5I</�E<��A<�<><��:<i�6<\3<�/<�+,<�(<g
%<�!<b�<'y<1�<"�<�<�</C	<��<M�<�o�;���;]N�;���;�g�;m�;���;~��;LV�;�;�;�1�;�9�;MS�;�~�;���;]�;|p�;��;�n�;#
�;]��;�y�;��x;zhn;�Zd;irZ;��P;�G;�=;N:4;�+;��!;��;�-;c|;���:���:�D�:y��:朻:��:FЛ:>8�:��y:�6[:�%=:[q:�:	�9���9�`/9�[{8��B���v4���e��� 򹻳��.��ZH�_b��8|�-�g���R]������$|��&�ɺ\Uֺ������b)�������	���Q�����1�!�3�'�ۭ-�j�3��9�]r?�IXE��<K��Q�&�V��\���b�D�h�-qn�MLt��&z�� ���킻Zۅ�EɈ�h���O����������Kw��Ui���  �  =u=�=޷=�X=��=I�=�:=�� =uz =� =4r�<��<���<)�<pd�<��<���<��<xI�<R��<��<���<5�<�P�<���<-��<j��<8�<�7�<?a�<H��<���<3��<���<��<|6�<"S�<�m�<���<���<9��<$��<q��<
��<���<���<���<h��<���<H��<.��<���<i��<���<���<xn�<N�<�)�<�<N��<R��<�m�<94�<��<X��<l�<Q �<���<�z�<"!�<���<�_�<O��<.��<o�<6��<�,�<a��<�+�<��<�<芴<���<�`�<�ů<�&�<I��<@ު<�4�<�<�ץ<�$�<�n�<���<���<�;�<�z�<���<*�<�*�<a�<~��<CȐ<O��<�(�<�V�<���<M��<�م<Q�<�+�<�S�<H�|<�Cy<b�u<g�q< (n<wsj<��f<�
c<�V_<��[<q�W<M@T<��P<9�L<�5I<:�E<��A< =><ș:<J�6<
\3<�/<�+,<��(<r
%<&�!<@�<y<�<:�<�<�<AC	<��<U�<Ro�;���;rN�;���;�g�;D�;���;X��;bV�;�;�;�1�;�9�;nS�;$�;��;c�;zp�;&�;�n�;
�;O��;ly�;њx;|hn;�Zd;[rZ;C�P;�G;��=;�:4;|+;�!;��;Q-;&|;i��:y��:�D�:���:���:�:�ϛ:�7�:�y:�6[:j&=:�o:m:�	�9M��9,f/9y[{8��B�C� 1���c��c�����.�	ZH��_b�z8|��񊺖����\��x���K{����ɺGUֺF�⺋��Q)�����R�	�������*����!���'��-�	�3�9�9�6r?��XE�h<K�XQ��V���\�#�b�B�h�yqn�4Lt��&z�� ���킻Hۅ�Ɉ�P���7�����������8w��}i���  �  Eu=�=�=�X=��=K�=�:=�� =mz =� =6r�<��<���<)�<�d�<��<���<��<}I�<V��<
��<���</�<�P�<q��<$��<j��<;�<�7�<4a�<U��<���<0��<���<��<n6�<S�<�m�<م�<Ǜ�<0��<$��<���<	��<���<���<���<h��<���<S��<!��<���<m��<���<��<�n�<$N�<�)�<�<Q��<W��<�m�<A4�<��<U��<l�<= �<���<�z�<.!�<���<�_�<Y��<'��<k�<-��<x,�<R��<�+�<��<�<�<���<�`�<�ů<�&�<D��<0ު<�4�<퇧<�ץ<�$�<�n�<���<���<�;�<�z�<���<5�<�*�<a�<���<DȐ<>��<�(�<�V�<���<E��<�م<X�<�+�<�S�<9�|<�Cy<j�u<Z�q<(n<[sj<׾f<�
c<�V_<��[<v�W<S@T<n�P<V�L<�5I<B�E<��A<�<><Й:<C�6<$\3<��/<�+,<�(<r
%<�!<N�<ey<�<B�<�<�<JC	<��<n�<7o�;���;7N�;���;�g�;Q�;���;+��;�V�;�;�;�1�;�9�;7S�;�~�;ؼ�;Y�;`p�;C�;�n�;
�;���;jy�;�x;�gn;�Zd;\rZ;m�P;4G;��=;�:4;�+;5�!;��;�-;�|;��:���:�D�:%��:q��:j��:WЛ:�7�:o�y:n4[:�&=:�o:�:q	�9J��9k/9;M{8ܓB�c
�w4��ng��a�U��� .�sXH��ab�W8|�[񊺷���(]��u���d{��$�ɺTֺh��k��
)�����	�	�����������!��'���-��3���9��q?��XE�><K��Q���V���\�$�b���h��qn�HLt��&z�� ���킻�ۅ�FɈ�����)���˕��셔�+w���i���  �  =u=�=޷=�X=��=I�=�:=�� =uz =� =4r�<��<���<)�<pd�<��<���<��<xI�<R��<��<���<5�<�P�<���<-��<j��<8�<�7�<?a�<H��<���<3��<���<��<|6�<"S�<�m�<���<���<9��<$��<q��<
��<���<���<���<h��<���<H��<.��<���<i��<���<���<xn�<N�<�)�<�<N��<R��<�m�<94�<��<X��<l�<Q �<���<�z�<"!�<���<�_�<O��<.��<o�<6��<�,�<a��<�+�<��<�<芴<���<�`�<�ů<�&�<I��<@ު<�4�<�<�ץ<�$�<�n�<���<���<�;�<�z�<���<*�<�*�<a�<~��<CȐ<O��<�(�<�V�<���<M��<�م<Q�<�+�<�S�<H�|<�Cy<b�u<g�q< (n<wsj<��f<�
c<�V_<��[<q�W<M@T<��P<9�L<�5I<:�E<��A< =><ș:<J�6<
\3<�/<�+,<��(<r
%<&�!<@�<y<�<:�<�<�<AC	<��<U�<Ro�;���;rN�;���;�g�;D�;���;X��;bV�;�;�;�1�;�9�;nS�;$�;��;c�;zp�;&�;�n�;
�;O��;ly�;њx;|hn;�Zd;[rZ;C�P;�G;��=;�:4;|+;�!;��;Q-;&|;i��:y��:�D�:���:���:�:�ϛ:�7�:�y:�6[:j&=:�o:m:�	�9M��9,f/9y[{8��B�C� 1���c��c�����.�	ZH��_b�z8|��񊺖����\��x���K{����ɺGUֺF�⺋��Q)�����R�	�������*����!���'��-�	�3�9�9�6r?��XE�h<K�XQ��V���\�#�b�B�h�yqn�4Lt��&z�� ���킻Hۅ�Ɉ�P���7�����������8w��}i���  �  =u=�=۷=�X=��=D�=�:=�� =wz =� =8r�<��<���<)�<yd�<$��<���<��<xI�<I��<��<���<B�<{P�<{��<(��<j��<B�<�7�<Ia�<C��<���<7��<���<��<l6�<S�<�m�<���<���<:��<'��<u��<��<���<���<���<j��<��<F��<1��<���<n��<���<���<�n�<N�<�)�<�<T��<M��<�m�<:4�<
��<]��<l�<R �<���<�z�<&!�<���<�_�<E��</��<o�<3��<x,�<Z��<�+�<��<�<ኴ<���<�`�<�ů<�&�<B��<<ު<�4�<���<�ץ<�$�<�n�<���<��<�;�<�z�<���<;�<�*�<�`�<���<7Ȑ<S��<�(�<�V�<���<E��<�م<I�<,�<�S�<\�|<�Cy<V�u<k�q<�'n<nsj<׾f<�
c<�V_<��[<k�W<D@T<��P<5�L<�5I</�E<��A<�<><��:<i�6<\3<�/<�+,<�(<g
%<�!<b�<'y<1�<"�<�<�</C	<��<M�<�o�;���;]N�;���;�g�;m�;���;~��;LV�;�;�;�1�;�9�;MS�;�~�;���;]�;|p�;��;�n�;#
�;]��;�y�;��x;zhn;�Zd;irZ;��P;�G;�=;N:4;�+;��!;��;�-;c|;���:���:�D�:y��:朻:��:FЛ:>8�:��y:�6[:�%=:[q:�:	�9���9�`/9�[{8��B���v4���e��� 򹻳��.��ZH�_b��8|�-�g���R]������$|��&�ɺ\Uֺ������b)�������	���Q�����1�!�3�'�ۭ-�j�3��9�]r?�IXE��<K��Q�&�V��\���b�D�h�-qn�MLt��&z�� ���킻Zۅ�EɈ�h���O����������Kw��Ui���  �  Cu=�=۷=�X=��=G�=�:=�� =pz =� =>r�<��<���<)�<{d�<��<���<��<{I�<F��<��<���<9�<P�<|��<'��<`��<@�<�7�<<a�<Q��<���<;��<���<��<{6�<%S�<�m�<ۅ�<ě�<3��<)��<}��<��<���<���<���<h��<���<E��<"��<���<o��<���<��<|n�<N�<�)�<�<T��<N��<�m�<84�<��<Y��<l�<I �<���<�z�<.!�<���<�_�<U��<'��<y�<<��<�,�<e��<�+�<��<�<�<���<�`�<�ů<�&�<E��<=ު<�4�<���<�ץ<�$�<�n�<���<��<�;�<�z�<���<,�<�*�<�`�<���<6Ȑ<D��<�(�<�V�<���<K��<�م<L�<�+�<�S�<T�|<�Cy<f�u<f�q<(n<ysj<��f<�
c<�V_<��[<p�W<Q@T<��P<P�L<�5I</�E<��A<�<><��:<R�6<\3<��/<�+,<�(<j
%<�!<>�<,y<�<�<�<�<)C	<��<P�<_o�;���;cN�;���;�g�;c�;���;L��;�V�;z;�;�1�;�9�;pS�;�;��;��;hp�;6�;�n�;+
�;|��;wy�;՚x;hn;�Zd;ZrZ;\�P;�G;��=;L:4;�+;��!;[�;l-;F|;���:���:�D�:���:*��:֛�:�ϛ:�7�:^�y:�5[:g&=:�o:�:�	�9���9�h/95L{8MzB�v�=1���b������� .��XH��`b�8|��-��� ]�������{����ɺTUֺd��3��N)�������	����S������!��'���-�o�3���9�Kr?��XE�n<K�nQ�j�V���\��b��h�Kqn�LLt��&z�� ���킻Dۅ�Ɉ�O��������������0w��mi���  �  Cu=�=�=�X=��=H�=�:=�� =sz =� =,r�<ޯ�<���<)�<yd�<��<���<��<qI�<K��<��<���<+�<�P�<|��<.��<m��<9�<�7�<7a�<[��<���<B��<���<��<~6�< S�<�m�<���<ӛ�<7��<'��<y��<
��<���<���<���<b��<���<J��<(��<���<\��<���<��<{n�<N�<�)�<�<B��<P��<�m�<;4�<���<Q��<$l�<G �<���<�z�<)!�<���<�_�<d��<.��<��<6��<�,�<\��<�+�<"��<�<���<���<�`�<�ů<�&�<O��<<ު<�4�<釧<�ץ<�$�<�n�<���<���<�;�<�z�<���<&�<�*�<�`�<s��<?Ȑ<K��<�(�<�V�<���<P��<�م<^�<�+�<�S�<G�|<�Cy<��u<l�q<"(n<lsj<�f<�
c<�V_<��[<��W<e@T<z�P<N�L<�5I<P�E<��A<=><Ù:<7�6<\3<	�/<�+,<�(<d
%<�!</�<'y<��<;�<�<��<2C	<��<R�<(o�;���;aN�;���;�g�;F�;о�;3��;�V�;�;�; 2�;�9�;GS�;+�;���;��;yp�;r�;�n�;!
�;m��;ky�;F�x;hn;�Zd;(rZ;��P;�G;ǒ=;z:4;+;��!;��;c-;L|;��:`��:�C�:���:x��:���:kϛ:y7�:أy:�5[:(=:�o:3:�
�92��98p/9�W{8IhB�b�c1��e��򹹱�8 .�yWH�ab�_7|��񊺉����\������={��h�ɺ_UֺI������)����@�	����Z��N��-�!��'�c�-�&�3�Y�9�r?�YE�n<K�HQ�_�V�n�\�)�b��h��qn�Lt�>&z�� ���킻`ۅ��Ȉ�n�����������ȅ��w���i���  �  Bu=�=�=�X=��=F�=�:=�� =qz =� =-r�<د�<���<)�<od�<��<���<��<pI�<A��<��<���<;�<~P�<y��<$��<v��<=�<�7�<Oa�<T��<���<A��<���<��<�6�<.S�<�m�<��<Ǜ�<H��<0��<x��<��<���<���<���<e��<���<A��<$��<���<c��<���<��<ln�<N�<�)�<�<I��<G��<�m�<34�<��<X��<l�<J �<���<�z�<(!�<���<�_�<Y��<5��<��<E��<�,�<i��<�+�< ��<�<���<���<�`�<�ů<�&�<@��<;ު<�4�<���<�ץ<�$�<�n�<���<���<�;�<�z�<���< �<�*�<�`�<v��<3Ȑ<F��<�(�<�V�<���<G��<�م<R�<,�<�S�<f�|<�Cy<u�u<p�q<"(n<�sj<�f<�
c<�V_<��[<��W<f@T<��P<J�L<�5I<B�E<��A<�<><��:<]�6<�[3<�/<�+,<�(<V
%<	�!<*�<y<�<�<�<��<C	<��<E�<fo�;���;QN�;���;�g�;U�;ľ�;���;�V�;�;�;�1�;�9�;{S�;7�;3��;��;�p�;@�;�n�;E
�;h��;�y�;��x;-hn;�Zd;?rZ;\�P;�G;��=;-:4;I+;��!;��;�,;�{;���:e��::D�:��:0��:���:�ϛ:�7�:��y:�5[:�%=:r::��9ؕ�9jj/9hf{8�lB�o���/��)b������M.��XH�^b��7|�|񊺠����]�������{����ɺ�Uֺ���w���)����̺	����������Z�!�b�'�L�-���3���9��r?�|XE��<K��Q�b�V���\���b���h�qn��Kt�r&z�} ���킻*ۅ��Ȉ�9���񥎻����΅��w��Di���  �  =u=�=ܷ=�X=��=A�=�:=�� =sz =� =.r�<ѯ�<���<)�<dd�<��<���<��<iI�<?��<��<���<>�<pP�<���<%��<n��<C�<�7�<Pa�<O��<���<A��< ��<��<~6�<9S�<�m�<���<ț�<G��<0��<r��<��<���<���<���<g��<���<4��<*��<���<e��<|��<��<ln�<�M�<�)�<� �<L��<9��<�m�<+4�<���<Y��<l�<Z �<���<�z�<'!�<���<�_�<Y��<C��<z�<O��<�,�<n��<�+�<��<*�<�<���<�`�<�ů<�&�<?��<Mު<�4�<���<�ץ<�$�<�n�<���<���<�;�<�z�<���<!�<�*�<�`�<x��<%Ȑ<M��<�(�<�V�<���<L��<�م<J�<
,�<�S�<m�|<�Cy<��u<��q<(n<�sj<��f<�
c<�V_<ɣ[<��W<[@T<��P<8�L<�5I<3�E<��A<=><��:<Z�6<�[3<�/<z+,<�(<H
%<�!<*�<�x<��<�<�<�<C	<��<'�<oo�;���;�N�;���;�g�;j�;���;���;vV�;�;�;�1�;�9�;�S�;&�;\��;��;�p�;A�;�n�;B
�;O��;�y�;~�x;�hn;\Zd;JrZ;�P;3G;Ւ=;�94;W+;&�!;{�;�,;�{;���:���:cD�:0��:���:���:Lϛ:�7�:נy:�7[:�$=:�q:�:�9���9j/9��{8�yB����0���`��u�q���.�YH�^b��8|�,������]�������|��w�ɺuVֺĪ�Y�*��ت�$�	������w����!���'�:�-���3�L�9��r?��XE��<K�aQ���V��\�{�b�@�h��pn��Kt�B&z�M ���킻�څ� Ɉ����󥎻t�������w��0i���  �  Cu=�=�=�X=��=E�=�:=�� =qz =� =&r�<ʯ�<���<�(�<id�< ��<���<��<dI�<C��<��<���<:�<xP�<}��<$��<r��<J�<�7�<Ja�<^��<���<K��<��<��<�6�<=S�<�m�<��<՛�<C��<5��<���<��<���<���<���<k��<���<;��<*��<���<Y��<���<��<in�<�M�<�)�< �<?��<;��<�m�</4�<���<\��<l�<K �<���<�z�<3!�<���<�_�<g��<@��<��<S��<�,�<n��<�+�<)��<)�<��<���<�`�<�ů<�&�<E��<?ު<�4�<���<�ץ<�$�<�n�<���<���<�;�<�z�<���<�<�*�<�`�<p��<+Ȑ<K��<�(�<�V�<���<H��<�م<W�<,�<�S�<m�|<�Cy<��u<��q<-(n<�sj<�f<�
c<�V_<ԣ[<��W<j@T<��P<Q�L<�5I<J�E<��A<�<><��:<J�6<�[3<�/<�+,<��(<9
%<�!<�<y<��<�<�<ܨ<!C	<��<5�<\o�;���;\N�;~��;�g�;��;Ծ�;}��;�V�;�;�;2�;:�;�S�;D�;h��;��;�p�;r�;�n�;R
�;���;�y�;	�x;hn;jZd;erZ;�P;fG;ϒ=;�94;�+;K�!;-�;�,;�{;��:���:�C�:G��:z��:=��:>ϛ:8�:t�y:�5[:'=:�q:T:��9���9�p/99z{8z`B�����.��"a��I����.��VH��^b��6|���������F]������b|����ɺVֺȪ�8���*��P���	�#����������!���'��-�͝3�W�9��r?��XE�{<K��Q�u�V���\���b�Еh��pn��Kt�&z�C ���킻�څ��Ȉ����Х��^��������v��>i���  �  Iu=�=�=�X=��=G�=�:=�� =gz =� =%r�<ʯ�<���<�(�<id�<��<���<��<mI�<9��<���<���<)�<�P�<{��<-��<u��<9�<�7�<Oa�<j��<���<U��<��<��<�6�<:S�<�m�<��<ڛ�<I��<9��<���<��<���<���<���<\��<���<;��<��<���<Q��<���<ڊ�<^n�<�M�<�)�<�<8��<F��<�m�<,4�<���<L��<$l�<H �<���<�z�<.!�<���<�_�<p��<;��<��<T��<�,�<|��<�+�<5��<"�<��<���<�`�<�ů<�&�<Q��<<ު<�4�<燧<�ץ<�$�<�n�<���<���<�;�<�z�<���<
�<�*�<�`�<k��<1Ȑ<3��<�(�<�V�<���<P��<�م<_�<�+�<�S�<s�|<�Cy<��u<��q<N(n<�sj<&�f<�
c<W_<�[<��W<�@T<��P<g�L<�5I<T�E<��A<=><��:<3�6<�[3<��/<�+,<ߘ(<:
%<�!<��<y<��<�<�<�<C	<d�<8�<o�;���;SN�;���;�g�;>�;��;���;�V�;�;�;C2�;$:�;�S�;{�;^��;��;�p�;��;�n�;b
�;���;zy�;K�x;hn;�Zd;�qZ;�P;cG;�=;
:4;�+;Z�!;��;r,;g{;M��:"��:C�:���:<��:��:Rϛ:7�:��y:�5[:+(=:�p:�:r�9�9!u/9�m{8�?B�}���*���]���򹢯��.��UH�I^b�|5|�������\������O{����ɺ�Uֺu��,��*��{���	�������.����!���'���-���3��9��r?�YE��<K�GQ�U�V�i�\��b���h��pn��Kt�&z�7 ��D킻�څ��Ȉ�	�������G��������v��2i���  �  Hu=�=�=�X=��=>�=�:=�� =kz =� =r�<ǯ�<���<�(�<ad�<���<���<��<^I�<2��<��<���</�<tP�<z��<'��<v��<F�<�7�<Ga�<a��<ʯ�<T��<���<��<�6�<8S�<�m�<���<���<G��<8��<���<��<���<���<���<S��<���<7��<��<���<L��<y��<���<en�<�M�<�)�<� �<2��<8��<�m�<)4�<��<H��<l�<K �<���<�z�<4!�<���<�_�<p��<M��<��<O��<�,�<��<�+�<4��<8�<��<���<�`�<�ů<�&�<I��<<ު<�4�<뇧<�ץ<�$�<�n�<���<���<�;�<�z�<���<�<�*�<�`�<c��<'Ȑ<:��<�(�<�V�<���<J��<�م<X�<,�<�S�<i�|<�Cy<��u<��q<.(n<�sj<*�f<�
c<�V_<�[<��W<u@T<��P<b�L<�5I<L�E<��A<�<><��:<E�6<�[3<��/<t+,<ɘ(<3
%<�!<�<�x<��<�<�<Ϩ<�B	<o�<:�<-o�;���;PN�;���;�g�;s�;��;m��;�V�;
<�;>2�;�9�;�S�;{�;T��;��;�p�;��;�n�;_
�;���;�y�;�x;$hn;�Zd;�qZ;-�P;>G;&�=;�94;�+;	�!;�;�,;~{;���:~��:�B�:��:&��:˚�:�ϛ:�6�:(�y:�5[:�&=:�q:<:�99u/9��{8FOB�_��+��8]����̯�9.��VH�_b�'6|�����ʰ��]������H|��l�ɺ�Uֺ?�⺄���*������	�j��&�������!��'��-��3��9��r?��XE�=K�rQ�R�V���\���b���h��pn��Kt��%z� ���킻�څ��Ȉ�붋�륎�3���o����v��Gi���  �  Fu=�=�=�X=��=@�=�:=�� =oz =� =r�<ǯ�<���<�(�<Sd�<��<���<��<TI�<5��<��<���<<�<pP�<���<!��<r��<Q�<�7�<Wa�<b��<ǯ�<Q��<��<��<�6�<OS�<�m�<���<ޛ�<L��<=��<���<!��<���<���<���<`��<���<0��<!��<q��<W��<r��<Ҋ�<[n�<�M�<~)�<� �<;��<'��<�m�<$4�<���<U��<l�<S �<���<�z�<8!�<���<�_�<o��<N��<��<e��<�,�<���<,�<3��<7�<��<���<�`�<�ů<�&�<C��<Hު<�4�<���<�ץ<�$�<�n�<���<���<�;�<�z�<z��<�<p*�<�`�<h��<Ȑ<E��<�(�<�V�<���<M��<�م<T�<,�<�S�<��|<�Cy<��u<��q<5(n<�sj<$�f<c<W_<�[<��W<w@T<��P<]�L<�5I<C�E<��A<=><��:<S�6<�[3<��/<b+,<ɘ(<3
%<�!<��<�x<��<�<�<��<C	<s�<%�<ao�;���;xN�;p��;�g�;��;��;���;�V�;�;�;22�;*:�;�S�;~�;���;��;�p�;��;o�;r
�;���;�y�;Śx;1hn;sZd;rZ;�P;G;��=;"94;�+;��!;��;U,;"{;���:���:OC�:��:Û�:~��:Mϛ:�7�:X�y:�6[:�%=:�r:�:��90��9Rt/9��{8mSB�m��q*��[�������h.�VH�]b�.6|����ɰ��s]������|����ɺHVֺK�����+��y����	�������%��t�!���'���-�X�3���9��r?��XE��<K�\Q�r�V���\�_�b���h��pn��Kt��%z� ��v킻�څ��Ȉ�����¥��7��������v��i���  �  Hu=�=�=�X=��=B�=�:=�� =jz =� =r�<¯�<���<�(�<bd�<���<���<��<\I�<7��<���<���<*�<yP�<���<+��<v��<B�<�7�<Sa�<m��<���<W��<��<��<�6�<AS�<�m�<���<���<Q��<9��<���<��<���<���<���<[��<���<3��<��<y��<T��<q��<֊�<bn�<�M�<�)�<� �<;��<2��<�m�<(4�<���<L��<l�<R �<���<�z�<4!�<���<�_�<u��<H��<��<[��<�,�<|��<,�<9��<0�<��<���<�`�<�ů<�&�<M��<Iު<�4�<燧<�ץ<�$�<�n�<���<���<�;�<�z�<���<�<v*�<�`�<f��<Ȑ<<��<�(�<�V�<���<Q��<�م<b�< ,�<�S�<t�|<�Cy<��u<��q<N(n<�sj<�f<�
c<W_<�[<��W<�@T<��P<e�L<�5I<Y�E<��A<=><��:<5�6<�[3<��/<l+,<̘(<)
%<�!<�<�x<��<�<�<ɨ<C	<b�<%�<o�;���;|N�;���;�g�;a�;��;���;�V�;�;�;J2�;9:�;�S�;\�;v��;��;�p�;��;o�;a
�;���;�y�;,�x;Ahn;�Zd;�qZ;�P; G;X�=;b94;�+;��!;��;�,;|{;,��:���:AC�:���:���:���:ϛ:�6�:<�y:�6[:_'=:�q:F:!�9|��9w/9x�{8�?B�x��V,��^�� �9��4.�QUH��]b��5|�����Ű���\�����D|����ɺoVֺ�����K+����z�	�z�������D�!��'�̮-�*�3�։9��r?�YE��<K�<Q�B�V�Q�\�͹b���h��pn�NKt��%z� ��E킻�څ��Ȉ�䶋�����&��������v��&i���  �  �s=�=��=oV=��=4�=.7=�� =^v =� =�h�<���<���<M�<X�<ԑ�<���<��<�9�<�o�<Ǥ�<���<�<�<�<�l�<F��<���<c��<��<ZG�<bn�<���<&��<���<P��<��<Y1�<�J�<�a�<Hv�<���<.��<?��<���<��<���<`��<׻�<=��<W��<���<F��<��<�l�<SS�<�5�<w�<��<���<%��<|f�<t0�<8��<���<ct�<�,�<���<A��<+;�<���<\��<� �<a��<�M�<�ݾ<�h�<��<kr�<��<�j�<��<�R�<���<�*�<쐯<t�<TR�<���<��<bZ�<���<g��<�E�<���<mԞ<��<�X�<>��<|ӗ<��<�E�<|�<���<s�<��<�D�<Bs�<���<�̅<2��<�"�<]L�<��|<�;y<�u<��q<�*n<�yj<��f<�c<�g_<�[<%	X<�[T<7�P<�M<n[I<g�E<�B<9m><n�:<k07<Ė3< 0<2m,<��(<�R%<�!<�I<��<#S<��<bq<	<j�	<�I<��<8H�;ض�;�2�;���;	W�;���; ��;
��;�X�;}A�;�;�;�F�;hc�;ّ�;�Ѩ;{$�;܈�;y��;숒;�$�;�҇;���;��z;��p;��f;�\;�R;�/I;��?;]O6;Y-;��#;��;]$;�j	;+� ;��:���:/g�:��:��:�%�:"x�:��:ca:�(C:�H%:��:i�9sD�9�"D9�ܥ8�'鷘7��1z�-���W�鹚���0*��D�n�^���x�C����Ѣ��y��=��O�Ⱥ պil�O��		���!��7	��H��S�Z�[!�.X'��P-�[E3�'79��$?��E���J���P�+�V�h�\�p�b�lh�rLn�h+t�z�x��j䂻eԅ�?Ĉ�������җ��ъ��7~��s���  �  �s=�=��=tV=��=-�=.7=�� =\v =� =�h�<���<���<R�<X�<ב�<���<��<�9�<�o�<���<���<&�<~<�<�l�<P��<���<n��<��<`G�<en�<���<��<���<N��<��<a1�<�J�<�a�<Xv�<���<6��<F��<���<��<���<N��<ٻ�<2��<?��<���<<��<��<m�<]S�<�5�<}�<%��<���<1��<uf�<w0�<$��<y��<gt�<�,�<���<F��<3;�<���<a��<� �<p��<�M�<qݾ<�h�<��<gr�<��<�j�<��<�R�<���<�*�<���<}�<^R�<���<��<jZ�<䫥<W��<�E�<���<Ԟ<��<�X�<>��<�ӗ<��<�E�<|�<���<s�<��<�D�<7s�<���<�̅<:��<�"�<`L�<��|<�;y<��u<��q<�*n<�yj<��f<�c<�g_<�[<5	X<�[T<C�P<�M<�[I<w�E<�B< m><S�:<k07<��3< 0<*m,<�(<�R%<�!<�I<��<*S<��<�q<	<m�	<�I<��<QH�;���;�2�;���;/W�;���;���;$��;�X�;�A�;�;�;�F�;cc�;���;�Ѩ;/$�;ʈ�;���;��;�$�;Ӈ;���;��z;��p;�f;��\;��R;�.I;��?;O6;�-;��#;)�;�$;�j	;h� ;g��:���:�f�:��:c�:)%�:^x�:-�:Jca:s)C:xI%:��:��9�F�9*D9�ۥ8Jw鷜4�W6z�@�����ӝ��0*�2�D���^���x�kB�����nТ��y�����ٔȺa	պem�$�����9!��7	��H��S��Y��Z!��W'�xP-��E3�(79��%?�%E�I�J�+�P���V�-�\�/�b��kh�9Ln�+t��
z�����䂻Gԅ��Ĉ� ���F����������@~��s���  �  �s=�=��=sV=��=1�=77=�� =dv =� =�h�<���<���<X�<X�<ۑ�<���<��<�9�<�o�<ɤ�<���<6�<�<�<�l�<J��<���<e��<��<^G�<[n�<���<��<���<T��<��<n1�<�J�<�a�<Sv�<���</��<:��<���<��<���<N��<��<<��<F��<��<8��<��<�l�<US�<�5�<x�<!��<���<4��<rf�<�0�<-��<���<vt�<�,�<���<>��<&;�<���<W��<� �<i��<�M�<sݾ<�h�<��<kr�<��<�j�<��<�R�<���<�*�<퐯<k�<WR�<���<��<zZ�<ꫥ<d��<�E�<���<�Ԟ<��<�X�<=��<�ӗ<��<�E�<|�<���<��<��<�D�<As�<���<�̅<0��<�"�<RL�<��|<�;y<�u<��q<�*n<�yj<��f<�c<�g_<��[<8	X<�[T<@�P<lM<q[I<b�E<�B<$m><a�:<�07<��3<8 0<,m,<
�(<�R%<��!<�I<��<2S<��<�q<	<x�	< J<��<�H�;���;�2�;���;�V�;���;׷�;��;wX�;�A�;�;�;�F�;zc�;���;,Ҩ;:$�;ƈ�;���;݈�;�$�;�҇;���;v�z;Șp;�f;j�\;�R;./I;Q�?;�N6;�-;��#;��;o$;�j	;L� ;ۧ�:���:�f�:�:��:�%�:Ry�:�:�ca:q(C:�G%:�:R�9�C�9�&D9sܥ8�m�.��6z�1���S��]���0*�X�D�I�^��x�C������Т��y�����ϓȺ�պ�lẉ��	��+!�8	��H��S��Y�[!��W'�yP-��E3��69��%?��E���J�%�P���V�|�\�q�b�Ylh�@Ln��+t��
z�����䂻ԅ��Ĉ�ϴ��#�����������g~��s���  �  �s=�=��=pV=��=2�=-7=�� =\v =� =�h�<���<���<[�<
X�<ۑ�<���<��<�9�<�o�<���<���<�<�<�<�l�<J��<���<i��<��<_G�<bn�<���<!��<���<H��<��<S1�<�J�<�a�<Mv�<���<6��<B��<���<��<���<_��<ֻ�<5��<J��<���<G��<���<m�<YS�<�5�<��<$��<���<6��<�f�<z0�<,��<��<_t�<�,�<���<C��<0;�<���<d��<� �<f��<�M�<zݾ<�h�<��<br�<��<�j�<��<�R�<���<�*�<���<v�<YR�<���<��<]Z�<<^��<�E�<���<|Ԟ<��<�X�<D��<�ӗ<��<�E�<%|�<���<s�<��<�D�<?s�<���<�̅<:��<�"�<[L�<��|<�;y<�u<��q<�*n<�yj<��f<�c<�g_<��[<	X<�[T<D�P<�M<y[I<w�E<�B<4m><f�:<e07<��3< 0<7m,<�(<�R%<�!<�I<��<2S<��<�q<	<o�	<�I<��<%H�;ɶ�;3�;���;!W�;���;��;��;�X�;^A�;�;�;�F�;Lc�;���;�Ѩ;T$�;���;���;���;�$�;�҇;���;��z;r�p;��f;ޛ\;��R;N/I;ĭ?;gO6;�-;��#;�;�$;k	;g� ;]��:���:�g�:%�:��:�%�:�w�:E�:�ba:!)C:0I%:n�:|�99E�9n%D9Sԥ8R�x;�H6z�S�����h��2*���D���^��x�}B������Т��y�������Ⱥ�պ�l���Z��N!��7	��H�S��Y��Z!��W'�HP-�TE3�+79�b%?�)E��J���P�5�V�)�\�<�b�lh�0Ln��+t�z����}䂻tԅ�}Ĉ�!���,�������䊔�C~��s���  �  �s=�=µ=qV=��=3�=.7=�� =\v =� =�h�<���<���<T�<X�<֑�<���<��<�9�<�o�<¤�<���<�<�<�<�l�<M��<���<]��<��<JG�<hn�<���<��<���<G��<��<N1�<�J�<�a�<Wv�<���<'��<;��<���<��<���<`��<׻�<>��<U��<���<L��<���<m�<YS�<�5�<��<"��<���<-��<�f�<z0�<6��<���<`t�<�,�<���<H��<&;�<���<T��<� �<n��<�M�<yݾ<�h�<��<ar�<��<�j�<��<�R�<���<�*�<鐯<u�<]R�<���<��<`Z�<���<c��<�E�<���<xԞ<��<�X�<F��<�ӗ<��<�E�<|�<���<t�<��<�D�<>s�<���<�̅<>��<�"�<VL�<��|<�;y<�u<�q<�*n<�yj<��f<�c<�g_<�[<	X<�[T< �P<{M<_[I<{�E<�B<+m><i�:<i07<Ė3< 0<Dm,<�(<�R%<�!<�I<��<)S<��<~q<	<|�	<�I<��<;H�;׶�;�2�;���;$W�;���;��;��;�X�;ZA�;�;�;�F�;Ic�;ʑ�;�Ѩ;I$�;���;���;ڈ�;$�;�҇;���;��z;N�p;��f;�\;(�R;�/I;ʭ?;�O6;�-;��#;�;�$;/k	;X� ;���:o��:�g�:0�:��:C&�:�w�:��:�aa:�)C:�G%:g�:��9�B�9�)D9IΥ8GS�d=��4z����� �鹃��}2*�܍D�2�^��x�/C�����{Т�oz��X��h�Ⱥ�պ�lằ��c��t!��7	��H�sS��Y��Z!��W'��P-�E3�!79��$?�E��J���P�4�V��\���b�?lh��Ln��+t��
z����䂻�ԅ�TĈ�:���7������ߊ��?~��Ns���  �  �s=�=��=sV=��=2�=37=�� =dv =� =�h�<���<���<a�<X�<��<���<��<�9�<�o�<Ȥ�<���<.�<�<�<�l�<N��<���<e��<��<SG�<Yn�<���<��<���<G��<��<^1�<�J�<�a�<Pv�<}��<1��<B��<���<��<���<N��<��<9��<H��<	��<<��<���<m�<_S�<�5�<��<*��<���<?��<rf�<�0�<+��<���<mt�<�,�<���<B��<#;�<���<[��<� �<c��<�M�<gݾ<�h�<��<\r�<��<�j�<��<�R�<���<�*�<�<l�<[R�<���<��<rZ�<뫥<b��<�E�<���<�Ԟ<��<�X�<L��<�ӗ<��<�E�<#|�<���<��<��<�D�<@s�<���<�̅<2��<�"�<[L�<��|<�;y<��u<s�q<�*n<�yj<��f<�c<}g_<շ[</	X<�[T<2�P<�M<m[I<c�E<�B<"m><d�:<|07<��3<7 0<4m,<�(<�R%<�!<�I<�<CS<��<�q<
	<��	<�I<��<yH�;���;�2�;���;�V�;���;��;��;rX�;�A�;F;�;�F�;Ic�;}��;�Ѩ;
$�;���;���;ǈ�;�$�;�҇;���;��z;��p;�f;4�\;��R;=/I;.�?;O6;
-;�#;:�;�$;Qk	;�� ;���:���:�f�:��:��:�%�:�x�:��:Xca:)C:�G%:'�:|�9vB�9$D9�ҥ8���6��;z����������y1*�͏D�F�^���x��B������Т��y��K��O�Ⱥ�պ�l�w��>	��� ��7	�EH�BS�iY��Z!�sW'�XP-��E3��69�j%?��E��J�,�P���V�g�\�w�b�lh�_Ln��+t��
z�@���䂻Wԅ��Ĉ����Y���?�������v~��*s���  �  �s=�=��=sV=��=0�=67=�� =hv =� =�h�<���<���<l�<X�<��<���<��<�9�<�o�<Ф�<���<5�<<�<�l�<G��<���<j��<��<^G�<Jn�<���<��<���<G��<��<Z1�<�J�<�a�<Dv�<���<-��<2��<���<��<»�<P��<��<?��<N��<��<=��<��<m�<cS�<�5�<��<1��<���<Q��<wf�<�0�<2��<���<qt�<�,�<���<8��<.;�<���<T��<� �<U��<�M�<[ݾ<�h�<��<]r�<��<�j�<��<�R�<���<�*�<�<r�<SR�<ɭ�<��<wZ�<쫥<j��<�E�<���<�Ԟ<��<�X�<B��<�ӗ<��<�E�<8|�<���<��<��<�D�<?s�<���<�̅<+��<�"�<HL�<��|<�;y<�u<��q<�*n<�yj<w�f<�c<gg_<�[<-	X<j[T<A�P<[M<{[I<[�E<�B<)m><]�:<�07<��3<G 0<0m,<3�(<S%<	�!<�I<��<[S<��<�q<$	<z�	<J<��<�H�;���;#3�;���;W�;���;ŷ�; ��;8X�;�A�;X;�;}F�;Lc�;k��;�Ѩ;�#�;舝;l��;Ո�;�$�;�҇;���;C�z;�p; �f;K�\;/�R;p/I;i�?;O6;�-;��#;_�;%;Tk	;�� ; ��:���:�f�:7�:^�:
&�:y�:Y�:�da:�'C:I%:�:��9D�9�D9o�81�鷫8��<z�e��� �鹹��v/*�ؑD��^�f�x��B����Ѣ��x�������Ⱥ�պ-l�p��}��k ��7	��G��S�Y��Z!�pW'��O-�E3�k69�c%?��E��J��P���V���\�/�b��lh�HLn�5,t�z�����䂻bԅ��Ĉ��������"��������~��s���  �  �s=�=��=qV=��=0�=37=�� =cv =� =�h�<���<���<m�<X�<��<���<��<�9�<�o�<Ϥ�<���<+�<�<�<�l�<B��<���<b��<��<XG�<Jn�<���<��<���<>��<��<O1�<�J�<�a�<9v�<}��<%��<1��<���<��<���<Y��<ܻ�<A��<Z��<��<L��<��<	m�<gS�<�5�<��<5��<���<?��<�f�<�0�<;��<���<gt�<�,�<���<<��<);�<~��<L��<� �<M��<�M�<aݾ<�h�<��<Ur�<��<�j�<��<�R�<���<�*�<鐯<o�<OR�<���<��<kZ�<���<k��<�E�<���<�Ԟ<��<�X�<H��<�ӗ<��<�E�</|�<���<�<��<�D�<<s�<���<�̅<.��<�"�<JL�<��|<�;y<׋u<y�q<�*n<�yj<��f<�c<qg_<ڷ[<	X<p[T<2�P<aM<l[I<c�E<�B<+m><`�:<�07<Ŗ3<3 0<Im,</�(<�R%<�!<�I<�<bS<��<�q<3	<��	<J<��<nH�;���;�2�;~��;
W�;���;���;��;9X�;_A�;b;�;xF�;'c�;���;�Ѩ;�#�;���;A��;Ɉ�;z$�;�҇;���;j�z;��p;k�f;�\;@�R;�/I;#�?;�O6;%-;�#;��; %;ck	;�� ;Ũ�:���:�g�:��:��:o&�:sx�:��:Lca:O(C:zH%:h�:��9VB�9�D92ӥ8?���<��;z��������2*�ۑD��^��x�"C��H��NѢ��y�������Ⱥ�պl������� ��7	��G�^S�Y��Z!��W'��O-�E3��69��$?��E�"�J���P��V���\�d�b��lh��Ln�,t�oz�+���䂻�ԅ��Ĉ�C���p���3�������~��*s���  �  �s=�=��=rV=��=7�=07=�� =^v =� =�h�<���<���<e�<%X�<��<���<��<�9�<�o�<ä�<���<%�<�<�<�l�<Q��<���<^��<��<HG�<Xn�<���<��<���<5��<��<E1�<�J�<�a�<Gv�<y��<(��<A��<���<��<���<[��<��<:��<S��<��<\��<���< m�<cS�<�5�<��<*��<���<9��<�f�<�0�<3��<���<kt�<�,�<���<K��<;�<���<U��<� �<\��<�M�<cݾ<�h�<��<Nr�<��<�j�<��<�R�<���<�*�<됯<g�<`R�<���<��<gZ�<���<`��<�E�<���<�Ԟ<��<�X�<]��<�ӗ<��<�E�<%|�<���<v�<��<�D�<Hs�<���<�̅<9��<�"�<\L�<��|<�;y<�u<Z�q<�*n<oyj<��f<�c<ug_<��[<	X<{[T<�P<�M<W[I<p�E<�B<%m><y�:<q07<��3<! 0<gm,<�(<S%<,�!<�I<.�<DS<��<�q<3	<��	<�I<��<UH�;��;�2�;���;�V�;���;���;��;rX�;?A�;>;�;rF�;c�;y��;�Ѩ;$�;]��;|��;���;�$�;�҇;a��;��z;M�p;�f;T�\;�R;�/I;��?;P6;�-;��#;b�;N%;�k	;�� ;���:8��:�h�:��:t�:&�:�x�:(�:�aa:?*C:�F%:پ:+�9�@�9o!D9���8Ĥ�(A��=z�������ş��3*�͏D���^�5�x��B�����6Т�Tz��_���Ⱥ0պ�l������ �7	�LH��R�*Y�eZ!�W'�IP-��D3�79��$?�E���J���P�/�V�0�\�ԋb�lh��Ln�,t�Az�����䂻�ԅ��Ĉ�x���g���j�������~��bs���  �  �s=�=��=uV=��=6�=67=�� =hv =� =�h�<���<���<j�<X�<��<���<��<�9�<�o�<Ԥ�<���<3�<�<�<�l�<T��<���<[��<��<FG�<Pn�<���<��<���<8��<��<G1�<�J�<�a�<Hv�<t��<"��<2��<|��<��<���<U��<��<E��<`��<��<U��<���< m�<eS�<�5�<��<-��<���<>��<�f�<�0�<B��<���<rt�<�,�<���<F��<;�<}��<K��<� �<]��<�M�<_ݾ<�h�<��<Nr�<��<�j�<��<�R�<���<�*�<㐯<g�<`R�<���<��<tZ�<���<p��<�E�<���<�Ԟ<��<�X�<T��<�ӗ<��<�E�<&|�<���<��<��<�D�<Hs�<���<�̅<6��<�"�<LL�<��|<�;y<�u<_�q<�*n<{yj<��f<�c<ig_<��[<	X<l[T<�P<^M<P[I<j�E<�B<"m><v�:<�07<Ŗ3<I 0<am,<�(<S%<1�!<�I<�<RS<��<�q<'	<��	<J<��<�H�;۶�;�2�;Ƚ�;W�;���;ŷ�;��;VX�;bA�;=;�;fF�;c�;q��;�Ѩ;�#�;x��;��;���;q$�;�҇;T��;��z;��p;T�f;e�\;a�R;	0I;w�?;�O6;-;��#;p�;L%;�k	;�� ;��:���:%h�:m�:i�:�&�:4y�:{�:�ba:�)C:hF%:a�:��9@�9�!D9�ȥ8U��M@��>z�����i�����2*���D�ֽ^�¸x�oC�����,Т�z������Ⱥ�պ�kẨ����� ��6	�H��R�Y�RZ!��V'�BP-��D3�g69��$?��E���J��P���V�I�\���b��lh��Ln�O,t�+z�����䂻�ԅ��Ĉ�_�������i���는��~��as���  �  �s=�=��=qV=��=1�=47=�� =gv =� =�h�<���<���<|�<X�<��<���<��<�9�<�o�<Ҥ�<���<+�<�<�<�l�<C��<���<g��<��<YG�<Fn�<���< ��<���<2��<��<E1�<�J�<�a�<<v�<~��<'��<1��<���<
��<���<S��<ۻ�<:��<P��<��<R��<	��<m�<yS�<�5�<��<F��<���<H��<�f�<�0�<3��<���<gt�<�,�<���<5��<1;�<��<M��<� �<N��<�M�<Vݾ<�h�<��<Er�<��<�j�<��<�R�<���<�*�<됯<t�<OR�<���<��<kZ�<�<k��<�E�<���<�Ԟ<��<�X�<L��<�ӗ<��<�E�<6|�<���<��<��<�D�<=s�<���<�̅<-��<�"�<DL�<��|<�;y<Ջu<d�q<w*n<yyj<u�f<�c<Vg_<·[<		X<h[T<3�P<OM<|[I<_�E<�B<.m><a�:<�07<��3<E 0<Om,<:�(<S%<:�!<�I<�<�S<��<�q<:	<��	<J<��<rH�;���;3�;���;W�;���;���;��;+X�;KA�;3;�;QF�;�b�;Q��;�Ѩ;�#�;���;N��;Ј�;�$�;�҇;ȓ�;@�z;p;>�f;�\;�R;�/I;^�?;�O6;e-;��#;�;�%;�k	;�� ;���:.��:2h�:!�:x�:�%�:�x�:��:�ca:�'C:�I%:��:n�9SC�9�D9�ȥ8��鷱A��Cz�㣳�Q�鹠��A3*�~�D�~�^�n�x��B�����=Ѣ�xy������ȺGպl������ �(7	�HG�?S��X�Z!��V'��O-�E3�o69�(%?��E��J���P��V���\�%�b��lh�xLn�5,t�tz�|���䂻�ԅ��Ĉ�g�������d�������~��&s���  �  �s=�=��=pV=��=6�=87=�� =gv =� =�h�<���<���<q�<X�<���<���<��<�9�<�o�<Ӥ�<���<4�<�<�<�l�<B��<���<Y��<��<GG�<Hn�<���<��<���<2��<��<E1�<�J�<�a�<>v�<r��<��<)��<���<��<���<[��<��<E��<[��<��<Z��<��<m�<nS�<�5�<��<9��<���<F��<�f�<�0�<=��<���<vt�<�,�<���<6��<!;�<u��<C��<� �<P��<�M�<_ݾ<�h�<��<Ir�<��<�j�<��<�R�<���<�*�<ᐯ<g�<NR�<���<��<sZ�< ��<p��<�E�<���<�Ԟ<��<�X�<S��<�ӗ<��<�E�<5|�<���<��<��<�D�<Js�<���<�̅<*��<�"�<AL�<��|<�;y<ڋu<c�q<�*n<pyj<s�f<�c<kg_<÷[<	X<c[T<�P<MM<\[I<U�E<�B<2m><w�:<�07<ɖ3<H 0<cm,<8�(<S%<)�!<�I<�<jS<��<�q<8	<��	<J<��<�H�;ٶ�;
3�;���;�V�;���;���;��;8X�;JA�;J;�;zF�;�b�;Z��;�Ѩ;�#�;{��;[��;���;W$�;�҇;���;M�z;��p;~�f;��\;g�R;�/I;��?;P6;X-;n�#;��;i%;�k	;� ;Z��:��:�h�:��:�:�&�:yy�:��:Gca:�'C:�G%:e�:�
�9N?�9�D9�ĥ8P�鷾@��Az�����
�鹹��c3*��D�½^�.�x��C�����JѢ��y�����#�Ⱥ{պ�k�y��t��� �?7	��G�S��X�VZ!�W'��O-��D3�_69��$?��E���J���P�#�V���\���b��lh��Ln�V,t�bz����䂻�ԅ��Ĉ�~���z���a�������~��cs���  �  �s=�=��=uV=��=2�=37=�� =ev =� =�h�<ĥ�<���<n�<,X�<��<���<��<�9�<�o�<̤�<���<+�<�<�<�l�<S��<���<`��<��<GG�<Pn�<���<���<���<(��<��<@1�<�J�<�a�<>v�<o��<,��<<��<���< ��<���<Q��<��<<��<\��<��<S��<��<(m�<oS�<�5�<��<6��<���<F��<�f�<�0�<;��<���<nt�<�,�<���<J��<;�<���<U��<� �<U��<�M�<\ݾ<�h�<��<@r�<��<�j�<��<�R�<���<�*�<됯<h�<`R�<���<��<lZ�<���<h��<�E�<���<�Ԟ<��<�X�<b��<�ӗ<��<�E�<,|�<���<��<��<�D�<Bs�<���<�̅<:��<�"�<]L�<��|<�;y<͋u<?�q<�*n<jyj<{�f<�c<ig_<��[<�X<h[T<!�P<�M<V[I<r�E<�B<m><e�:<07<ʖ3<= 0<fm,<(�(<0S%<:�!<�I<<�<[S<��<�q<$	<��	<J<��<rH�;���;�2�;Ƚ�;W�;���; ��;��;WX�;&A�;;�;PF�;�b�;T��;{Ѩ;�#�;7��;X��;���;�$�;�҇;l��;��z;��p;.�f;R�\;"�R;�/I;Y�?;�O6;K-;�#;��;�%;�k	; � ;���:��:�g�::�:��:6&�:�x�:
�:*ca:I*C:�F%:*�:o�9�>�9'D9�8���zD��Cz�,���	��B���4*���D���^��x��B�����*Т��y�������Ⱥ�պAlẾ��R��_ ��6	��G��R��X�Z!��V'�P-��D3��69��$?��E���J��P���V�)�\�ҋb�lh��Ln�X,t��z����䂻�ԅ��Ĉ�����������������~��Ks���  �  �s=�=��=pV=��=6�=87=�� =gv =� =�h�<���<���<q�<X�<���<���<��<�9�<�o�<Ӥ�<���<4�<�<�<�l�<B��<���<Y��<��<GG�<Hn�<���<��<���<2��<��<E1�<�J�<�a�<>v�<r��<��<)��<���<��<���<[��<��<E��<[��<��<Z��<��<m�<nS�<�5�<��<9��<���<F��<�f�<�0�<=��<���<vt�<�,�<���<6��<!;�<u��<C��<� �<P��<�M�<_ݾ<�h�<��<Ir�<��<�j�<��<�R�<���<�*�<ᐯ<g�<NR�<���<��<sZ�< ��<p��<�E�<���<�Ԟ<��<�X�<S��<�ӗ<��<�E�<5|�<���<��<��<�D�<Js�<���<�̅<*��<�"�<AL�<��|<�;y<ڋu<c�q<�*n<pyj<s�f<�c<kg_<÷[<	X<c[T<�P<MM<\[I<U�E<�B<2m><w�:<�07<ɖ3<H 0<cm,<8�(<S%<)�!<�I<�<jS<��<�q<8	<��	<J<��<�H�;ٶ�;
3�;���;�V�;���;���;��;8X�;JA�;J;�;zF�;�b�;Z��;�Ѩ;�#�;{��;[��;���;W$�;�҇;���;M�z;��p;~�f;��\;g�R;�/I;��?;P6;X-;n�#;��;i%;�k	;� ;Z��:��:�h�:��:�:�&�:yy�:��:Gca:�'C:�G%:e�:�
�9N?�9�D9�ĥ8P�鷾@��Az�����
�鹹��c3*��D�½^�.�x��C�����JѢ��y�����#�Ⱥ{պ�k�y��t��� �?7	��G�S��X�VZ!�W'��O-��D3�_69��$?��E���J���P�#�V���\���b��lh��Ln�V,t�bz����䂻�ԅ��Ĉ�~���z���a�������~��cs���  �  �s=�=��=qV=��=1�=47=�� =gv =� =�h�<���<���<|�<X�<��<���<��<�9�<�o�<Ҥ�<���<+�<�<�<�l�<C��<���<g��<��<YG�<Fn�<���< ��<���<2��<��<E1�<�J�<�a�<<v�<~��<'��<1��<���<
��<���<S��<ۻ�<:��<P��<��<R��<	��<m�<yS�<�5�<��<F��<���<H��<�f�<�0�<3��<���<gt�<�,�<���<5��<1;�<��<M��<� �<N��<�M�<Vݾ<�h�<��<Er�<��<�j�<��<�R�<���<�*�<됯<t�<OR�<���<��<kZ�<�<k��<�E�<���<�Ԟ<��<�X�<L��<�ӗ<��<�E�<6|�<���<��<��<�D�<=s�<���<�̅<-��<�"�<DL�<��|<�;y<Ջu<d�q<w*n<yyj<u�f<�c<Vg_<·[<		X<h[T<3�P<OM<|[I<_�E<�B<.m><a�:<�07<��3<E 0<Om,<:�(<S%<:�!<�I<�<�S<��<�q<:	<��	<J<��<rH�;���;3�;���;W�;���;���;��;+X�;KA�;3;�;QF�;�b�;Q��;�Ѩ;�#�;���;N��;Ј�;�$�;�҇;ȓ�;@�z;p;>�f;�\;�R;�/I;^�?;�O6;e-;��#;�;�%;�k	;�� ;���:.��:2h�:!�:x�:�%�:�x�:��:�ca:�'C:�I%:��:n�9SC�9�D9�ȥ8��鷱A��Cz�㣳�Q�鹠��A3*�~�D�~�^�n�x��B�����=Ѣ�xy������ȺGպl������ �(7	�HG�?S��X�Z!��V'��O-�E3�o69�(%?��E��J���P��V���\�%�b��lh�xLn�5,t�tz�|���䂻�ԅ��Ĉ�g�������d�������~��&s���  �  �s=�=��=uV=��=6�=67=�� =hv =� =�h�<���<���<j�<X�<��<���<��<�9�<�o�<Ԥ�<���<3�<�<�<�l�<T��<���<[��<��<FG�<Pn�<���<��<���<8��<��<G1�<�J�<�a�<Hv�<t��<"��<2��<|��<��<���<U��<��<E��<`��<��<U��<���< m�<eS�<�5�<��<-��<���<>��<�f�<�0�<B��<���<rt�<�,�<���<F��<;�<}��<K��<� �<]��<�M�<_ݾ<�h�<��<Nr�<��<�j�<��<�R�<���<�*�<㐯<g�<`R�<���<��<tZ�<���<p��<�E�<���<�Ԟ<��<�X�<T��<�ӗ<��<�E�<&|�<���<��<��<�D�<Hs�<���<�̅<6��<�"�<LL�<��|<�;y<�u<_�q<�*n<{yj<��f<�c<ig_<��[<	X<l[T<�P<^M<P[I<j�E<�B<"m><v�:<�07<Ŗ3<I 0<am,<�(<S%<1�!<�I<�<RS<��<�q<'	<��	<J<��<�H�;۶�;�2�;Ƚ�;W�;���;ŷ�;��;VX�;bA�;=;�;fF�;c�;q��;�Ѩ;�#�;x��;��;���;q$�;�҇;T��;��z;��p;T�f;e�\;a�R;	0I;w�?;�O6;-;��#;p�;L%;�k	;�� ;��:���:%h�:m�:i�:�&�:4y�:{�:�ba:�)C:hF%:a�:��9@�9�!D9�ȥ8U��M@��>z�����i�����2*���D�ֽ^�¸x�oC�����,Т�z������Ⱥ�պ�kẨ����� ��6	�H��R�Y�RZ!��V'�BP-��D3�g69��$?��E���J��P���V�I�\���b��lh��Ln�O,t�+z�����䂻�ԅ��Ĉ�_�������i���는��~��as���  �  �s=�=��=rV=��=7�=07=�� =^v =� =�h�<���<���<e�<%X�<��<���<��<�9�<�o�<ä�<���<%�<�<�<�l�<Q��<���<^��<��<HG�<Xn�<���<��<���<5��<��<E1�<�J�<�a�<Gv�<y��<(��<A��<���<��<���<[��<��<:��<S��<��<\��<���< m�<cS�<�5�<��<*��<���<9��<�f�<�0�<3��<���<kt�<�,�<���<K��<;�<���<U��<� �<\��<�M�<cݾ<�h�<��<Nr�<��<�j�<��<�R�<���<�*�<됯<g�<`R�<���<��<gZ�<���<`��<�E�<���<�Ԟ<��<�X�<]��<�ӗ<��<�E�<%|�<���<v�<��<�D�<Hs�<���<�̅<9��<�"�<\L�<��|<�;y<�u<Z�q<�*n<oyj<��f<�c<ug_<��[<	X<{[T<�P<�M<W[I<p�E<�B<%m><y�:<q07<��3<! 0<gm,<�(<S%<,�!<�I<.�<DS<��<�q<3	<��	<�I<��<UH�;��;�2�;���;�V�;���;���;��;rX�;?A�;>;�;rF�;c�;y��;�Ѩ;$�;]��;|��;���;�$�;�҇;a��;��z;M�p;�f;T�\;�R;�/I;��?;P6;�-;��#;b�;N%;�k	;�� ;���:8��:�h�:��:t�:&�:�x�:(�:�aa:?*C:�F%:پ:+�9�@�9o!D9���8Ĥ�(A��=z�������ş��3*�͏D���^�5�x��B�����6Т�Tz��_���Ⱥ0պ�l������ �7	�LH��R�*Y�eZ!�W'�IP-��D3�79��$?�E���J���P�/�V�0�\�ԋb�lh��Ln�,t�Az�����䂻�ԅ��Ĉ�x���g���j�������~��bs���  �  �s=�=��=qV=��=0�=37=�� =cv =� =�h�<���<���<m�<X�<��<���<��<�9�<�o�<Ϥ�<���<+�<�<�<�l�<B��<���<b��<��<XG�<Jn�<���<��<���<>��<��<O1�<�J�<�a�<9v�<}��<%��<1��<���<��<���<Y��<ܻ�<A��<Z��<��<L��<��<	m�<gS�<�5�<��<5��<���<?��<�f�<�0�<;��<���<gt�<�,�<���<<��<);�<~��<L��<� �<M��<�M�<aݾ<�h�<��<Ur�<��<�j�<��<�R�<���<�*�<鐯<o�<OR�<���<��<kZ�<���<k��<�E�<���<�Ԟ<��<�X�<H��<�ӗ<��<�E�</|�<���<�<��<�D�<<s�<���<�̅<.��<�"�<JL�<��|<�;y<׋u<y�q<�*n<�yj<��f<�c<qg_<ڷ[<	X<p[T<2�P<aM<l[I<c�E<�B<+m><`�:<�07<Ŗ3<3 0<Im,</�(<�R%<�!<�I<�<bS<��<�q<3	<��	<J<��<nH�;���;�2�;~��;
W�;���;���;��;9X�;_A�;b;�;xF�;'c�;���;�Ѩ;�#�;���;A��;Ɉ�;z$�;�҇;���;j�z;��p;k�f;�\;@�R;�/I;#�?;�O6;%-;�#;��; %;ck	;�� ;Ũ�:���:�g�:��:��:o&�:sx�:��:Lca:O(C:zH%:h�:��9VB�9�D92ӥ8?���<��;z��������2*�ۑD��^��x�"C��H��NѢ��y�������Ⱥ�պl������� ��7	��G�^S�Y��Z!��W'��O-�E3��69��$?��E�"�J���P��V���\�d�b��lh��Ln�,t�oz�+���䂻�ԅ��Ĉ�C���p���3�������~��*s���  �  �s=�=��=sV=��=0�=67=�� =hv =� =�h�<���<���<l�<X�<��<���<��<�9�<�o�<Ф�<���<5�<<�<�l�<G��<���<j��<��<^G�<Jn�<���<��<���<G��<��<Z1�<�J�<�a�<Dv�<���<-��<2��<���<��<»�<P��<��<?��<N��<��<=��<��<m�<cS�<�5�<��<1��<���<Q��<wf�<�0�<2��<���<qt�<�,�<���<8��<.;�<���<T��<� �<U��<�M�<[ݾ<�h�<��<]r�<��<�j�<��<�R�<���<�*�<�<r�<SR�<ɭ�<��<wZ�<쫥<j��<�E�<���<�Ԟ<��<�X�<B��<�ӗ<��<�E�<8|�<���<��<��<�D�<?s�<���<�̅<+��<�"�<HL�<��|<�;y<�u<��q<�*n<�yj<w�f<�c<gg_<�[<-	X<j[T<A�P<[M<{[I<[�E<�B<)m><]�:<�07<��3<G 0<0m,<3�(<S%<	�!<�I<��<[S<��<�q<$	<z�	<J<��<�H�;���;#3�;���;W�;���;ŷ�; ��;8X�;�A�;X;�;}F�;Lc�;k��;�Ѩ;�#�;舝;l��;Ո�;�$�;�҇;���;C�z;�p; �f;K�\;/�R;p/I;i�?;O6;�-;��#;_�;%;Tk	;�� ; ��:���:�f�:7�:^�:
&�:y�:Y�:�da:�'C:I%:�:��9D�9�D9o�81�鷫8��<z�e��� �鹹��v/*�ؑD��^�f�x��B����Ѣ��x�������Ⱥ�պ-l�p��}��k ��7	��G��S�Y��Z!�pW'��O-�E3�k69�c%?��E��J��P���V���\�/�b��lh�HLn�5,t�z�����䂻bԅ��Ĉ��������"��������~��s���  �  �s=�=��=sV=��=2�=37=�� =dv =� =�h�<���<���<a�<X�<��<���<��<�9�<�o�<Ȥ�<���<.�<�<�<�l�<N��<���<e��<��<SG�<Yn�<���<��<���<G��<��<^1�<�J�<�a�<Pv�<}��<1��<B��<���<��<���<N��<��<9��<H��<	��<<��<���<m�<_S�<�5�<��<*��<���<?��<rf�<�0�<+��<���<mt�<�,�<���<B��<#;�<���<[��<� �<c��<�M�<gݾ<�h�<��<\r�<��<�j�<��<�R�<���<�*�<�<l�<[R�<���<��<rZ�<뫥<b��<�E�<���<�Ԟ<��<�X�<L��<�ӗ<��<�E�<#|�<���<��<��<�D�<@s�<���<�̅<2��<�"�<[L�<��|<�;y<��u<s�q<�*n<�yj<��f<�c<}g_<շ[</	X<�[T<2�P<�M<m[I<c�E<�B<"m><d�:<|07<��3<7 0<4m,<�(<�R%<�!<�I<�<CS<��<�q<
	<��	<�I<��<yH�;���;�2�;���;�V�;���;��;��;rX�;�A�;F;�;�F�;Ic�;}��;�Ѩ;
$�;���;���;ǈ�;�$�;�҇;���;��z;��p;�f;4�\;��R;=/I;.�?;O6;
-;�#;:�;�$;Qk	;�� ;���:���:�f�:��:��:�%�:�x�:��:Xca:)C:�G%:'�:|�9vB�9$D9�ҥ8���6��;z����������y1*�͏D�F�^���x��B������Т��y��K��O�Ⱥ�պ�l�w��>	��� ��7	�EH�BS�iY��Z!�sW'�XP-��E3��69�j%?��E��J�,�P���V�g�\�w�b�lh�_Ln��+t��
z�@���䂻Wԅ��Ĉ����Y���?�������v~��*s���  �  �s=�=µ=qV=��=3�=.7=�� =\v =� =�h�<���<���<T�<X�<֑�<���<��<�9�<�o�<¤�<���<�<�<�<�l�<M��<���<]��<��<JG�<hn�<���<��<���<G��<��<N1�<�J�<�a�<Wv�<���<'��<;��<���<��<���<`��<׻�<>��<U��<���<L��<���<m�<YS�<�5�<��<"��<���<-��<�f�<z0�<6��<���<`t�<�,�<���<H��<&;�<���<T��<� �<n��<�M�<yݾ<�h�<��<ar�<��<�j�<��<�R�<���<�*�<鐯<u�<]R�<���<��<`Z�<���<c��<�E�<���<xԞ<��<�X�<F��<�ӗ<��<�E�<|�<���<t�<��<�D�<>s�<���<�̅<>��<�"�<VL�<��|<�;y<�u<�q<�*n<�yj<��f<�c<�g_<�[<	X<�[T< �P<{M<_[I<{�E<�B<+m><i�:<i07<Ė3< 0<Dm,<�(<�R%<�!<�I<��<)S<��<~q<	<|�	<�I<��<;H�;׶�;�2�;���;$W�;���;��;��;�X�;ZA�;�;�;�F�;Ic�;ʑ�;�Ѩ;I$�;���;���;ڈ�;$�;�҇;���;��z;N�p;��f;�\;(�R;�/I;ʭ?;�O6;�-;��#;�;�$;/k	;X� ;���:o��:�g�:0�:��:C&�:�w�:��:�aa:�)C:�G%:g�:��9�B�9�)D9IΥ8GS�d=��4z����� �鹃��}2*�܍D�2�^��x�/C�����{Т�oz��X��h�Ⱥ�պ�lằ��c��t!��7	��H�sS��Y��Z!��W'��P-�E3�!79��$?�E��J���P�4�V��\���b�?lh��Ln��+t��
z����䂻�ԅ�TĈ�:���7������ߊ��?~��Ns���  �  �s=�=��=pV=��=2�=-7=�� =\v =� =�h�<���<���<[�<
X�<ۑ�<���<��<�9�<�o�<���<���<�<�<�<�l�<J��<���<i��<��<_G�<bn�<���<!��<���<H��<��<S1�<�J�<�a�<Mv�<���<6��<B��<���<��<���<_��<ֻ�<5��<J��<���<G��<���<m�<YS�<�5�<��<$��<���<6��<�f�<z0�<,��<��<_t�<�,�<���<C��<0;�<���<d��<� �<f��<�M�<zݾ<�h�<��<br�<��<�j�<��<�R�<���<�*�<���<v�<YR�<���<��<]Z�<<^��<�E�<���<|Ԟ<��<�X�<D��<�ӗ<��<�E�<%|�<���<s�<��<�D�<?s�<���<�̅<:��<�"�<[L�<��|<�;y<�u<��q<�*n<�yj<��f<�c<�g_<��[<	X<�[T<D�P<�M<y[I<w�E<�B<4m><f�:<e07<��3< 0<7m,<�(<�R%<�!<�I<��<2S<��<�q<	<o�	<�I<��<%H�;ɶ�;3�;���;!W�;���;��;��;�X�;^A�;�;�;�F�;Lc�;���;�Ѩ;T$�;���;���;���;�$�;�҇;���;��z;r�p;��f;ޛ\;��R;N/I;ĭ?;gO6;�-;��#;�;�$;k	;g� ;]��:���:�g�:%�:��:�%�:�w�:E�:�ba:!)C:0I%:n�:|�99E�9n%D9Sԥ8R�x;�H6z�S�����h��2*���D���^��x�}B������Т��y�������Ⱥ�պ�l���Z��N!��7	��H�S��Y��Z!��W'�HP-�TE3�+79�b%?�)E��J���P�5�V�)�\�<�b�lh�0Ln��+t�z����}䂻tԅ�}Ĉ�!���,�������䊔�C~��s���  �  �s=�=��=sV=��=1�=77=�� =dv =� =�h�<���<���<X�<X�<ۑ�<���<��<�9�<�o�<ɤ�<���<6�<�<�<�l�<J��<���<e��<��<^G�<[n�<���<��<���<T��<��<n1�<�J�<�a�<Sv�<���</��<:��<���<��<���<N��<��<<��<F��<��<8��<��<�l�<US�<�5�<x�<!��<���<4��<rf�<�0�<-��<���<vt�<�,�<���<>��<&;�<���<W��<� �<i��<�M�<sݾ<�h�<��<kr�<��<�j�<��<�R�<���<�*�<퐯<k�<WR�<���<��<zZ�<ꫥ<d��<�E�<���<�Ԟ<��<�X�<=��<�ӗ<��<�E�<|�<���<��<��<�D�<As�<���<�̅<0��<�"�<RL�<��|<�;y<�u<��q<�*n<�yj<��f<�c<�g_<��[<8	X<�[T<@�P<lM<q[I<b�E<�B<$m><a�:<�07<��3<8 0<,m,<
�(<�R%<��!<�I<��<2S<��<�q<	<x�	< J<��<�H�;���;�2�;���;�V�;���;׷�;��;wX�;�A�;�;�;�F�;zc�;���;,Ҩ;:$�;ƈ�;���;݈�;�$�;�҇;���;v�z;Șp;�f;j�\;�R;./I;Q�?;�N6;�-;��#;��;o$;�j	;L� ;ۧ�:���:�f�:�:��:�%�:Ry�:�:�ca:q(C:�G%:�:R�9�C�9�&D9sܥ8�m�.��6z�1���S��]���0*�X�D�I�^��x�C������Т��y�����ϓȺ�պ�lẉ��	��+!�8	��H��S��Y�[!��W'�yP-��E3��69��%?��E���J�%�P���V�|�\�q�b�Ylh�@Ln��+t��
z�����䂻ԅ��Ĉ�ϴ��#�����������g~��s���  �  �s=�=��=tV=��=-�=.7=�� =\v =� =�h�<���<���<R�<X�<ב�<���<��<�9�<�o�<���<���<&�<~<�<�l�<P��<���<n��<��<`G�<en�<���<��<���<N��<��<a1�<�J�<�a�<Xv�<���<6��<F��<���<��<���<N��<ٻ�<2��<?��<���<<��<��<m�<]S�<�5�<}�<%��<���<1��<uf�<w0�<$��<y��<gt�<�,�<���<F��<3;�<���<a��<� �<p��<�M�<qݾ<�h�<��<gr�<��<�j�<��<�R�<���<�*�<���<}�<^R�<���<��<jZ�<䫥<W��<�E�<���<Ԟ<��<�X�<>��<�ӗ<��<�E�<|�<���<s�<��<�D�<7s�<���<�̅<:��<�"�<`L�<��|<�;y<��u<��q<�*n<�yj<��f<�c<�g_<�[<5	X<�[T<C�P<�M<�[I<w�E<�B< m><S�:<k07<��3< 0<*m,<�(<�R%<�!<�I<��<*S<��<�q<	<m�	<�I<��<QH�;���;�2�;���;/W�;���;���;$��;�X�;�A�;�;�;�F�;cc�;���;�Ѩ;/$�;ʈ�;���;��;�$�;Ӈ;���;��z;��p;�f;��\;��R;�.I;��?;O6;�-;��#;)�;�$;�j	;h� ;g��:���:�f�:��:c�:)%�:^x�:-�:Jca:s)C:xI%:��:��9�F�9*D9�ۥ8Jw鷜4�W6z�@�����ӝ��0*�2�D���^���x�kB�����nТ��y�����ٔȺa	պem�$�����9!��7	��H��S��Y��Z!��W'�xP-��E3�(79��%?�%E�I�J�+�P���V�-�\�/�b��kh�9Ln�+t��
z�����䂻Gԅ��Ĉ� ���F����������@~��s���  �  Dr==��= T=T�=G�=�3=i� =�r =Z =�_�<���<���<O�<aL�<_��<���<���<!+�<P`�<n��<d��<��<�)�<�X�<���<��<���<�<�.�<�T�< y�<���<���<y��<���<Y�<�)�<i?�<�R�<�c�<lr�<H~�<x��<܍�<H��<ґ�<&��<^��<h��<�s�<+d�<�P�<�9�</�<� �<���<S��<7��<�_�<�-�<���<)��<�|�<{9�<���<^��<�T�<���<��<�G�<^��<f~�<�<U��<1/�<ƶ�<:�<@��<G4�<��<�<	��<&��<�_�<Kí<�#�<=��<�٨<�/�<���<�ң<��<�i�<J��<R��<�8�<�x�<˶�<��<g,�<Nd�<}��<�Ύ<�<y3�<�c�<Ғ�<���<��<��<"E�<��|<24y<��u<��q<-n<<j<��f<$c<9w_<��[<LX<uT<�P<�$M<�~I<,�E<�9B<��><�:<cd7<�3<�:0<�,<2)<L�%<�"<q�<'<W�<4<��<�c<�
<P�<W<
 <��;�	�;D��;k7�;���;X��;�m�;5J�;�6�;h4�;�B�;�a�;���;�ԩ;)�;��;��;��;�,�;5ۈ;���;��|;��r;E�h;b�^;T�T;�.K;�A;�C8;� /;��%;n�;�;�<;'�;�)�:GY�:���:�e�:k>�:�I�:ǈ�:d��:a4g:�H:��*:?:[q�9]X�9z�W9���8ht-�����i��X���������{&���@�+J[��hu�[���{���%Y���������KǺd�Ӻ]>�|��-������ĺ�;�����:��M� ���&�%�,�[�2�M�8���>���D�ɺJ�Y�P���V��x\��_b�2Eh��)n�Ct���y�R��܂�@΅�����\���}�������Џ��d����|���  �  Lr==��= T=L�=C�=�3=b� =�r =Y =�_�<���<���<L�<GL�<^��<���<���<+�<J`�<g��<X��<#��<�)�<�X�<���<��<���<"�<�.�<�T�<y�<p��<��<���<
��<d�<|)�<l?�<�R�<�c�<xr�<_~�<���<֍�<H��<���<(��<]��<Q��<�s�<)d�<�P�<�9�<8�<� �<���<Y��</��<�_�<�-�<���<��<�|�<�9�<���<[��<�T�<���<���<�G�<`��<k~�<�<B��<5/�<Ѷ�<#:�<7��<44�<'��<
�<��<5��<�_�<Wí<�#�<5��<�٨<�/�<���<�ң<��<�i�<T��<H��<�8�<�x�<Ŷ�<��<g,�<Ud�<{��<�Ύ<��<�3�<�c�<���<���<��<��<3E�<��|<%4y<��u<��q<�,n<_j<��f<<$c<w_<��[<jX<uT<�P<�$M<�~I<+�E<�9B<y�><�:<�d7<��3<�:0<�,<<)<S�%<�"<k�<�<V�<4<��<�c<�
<B�<�V<.
 <��;d	�;>��;�7�;���;���;�m�;J�;�6�; 4�;KB�;�a�;���;	թ;�(�;��;��;��;.-�;�ۈ;;��|;��r;��h;w�^;M�T;(.K;��A;�C8;/;��%;��;��;:<;Z�;o)�:/Z�:���:Ge�:=�:uI�:B��:P��:4g:F�H:��*:�:u�9�X�9�W9˺�8.�u����i��U��0��9���y&��@��I[�gu�Ъ��Ì��eY��&��h���JǺ�Ӻ�>��캊���H����9��g��j��� ���&���,�c�2�b�8��>���D��J�ܦP���V��x\�&_b��Dh�~)n�wt��y����T܂��ͅ�X������Ҧ�������������w|���  �  Er==��=%T=Q�=B�=�3=c� =�r =W =�_�<���<���<[�<JL�<r��<���<���<+�<L`�<w��<Z��<*��<�)�<�X�<���<��<���<�<�.�<�T�<y�<r��<���<���<���<c�<)�<r?�<�R�<�c�<nr�<O~�<y��<֍�<Y��<���<,��<b��<[��<t�<!d�<�P�<�9�<@�<� �<���<f��<#��<�_�<�-�<���<!��<�|�<�9�<���<j��<�T�<���<��<�G�<Y��<d~�<�<E��<6/�<���<:�<=��<64�<.��<�<��<(��<�_�<Pí<�#�<@��<�٨<�/�<���<�ң<��<�i�<Y��<?��<�8�<�x�<ж�<��<^,�<Sd�<v��<ώ<��<�3�<�c�<ƒ�<���<��<��<%E�<��|<4y<��u<��q<�,n<Wj<v�f<.$c<w_<��[<tX<uT<�P<�$M<�~I< �E<�9B<��><�:<�d7<��3<�:0<�,<3)<H�%<�"<��<�<~�<�3<��<qc<�
<c�<�V<<
 <��;�	�;V��;x7�;���;V��;�m�;J�;7�;,4�;eB�;�a�;b��;թ;�(�;+��;��;쐓;-�;Sۈ;ě�;��|;@�r;��h;��^;z�T;{.K;H�A;�C8;+/;H�%;��;��;n<;��;�(�:zZ�:���:8f�:�=�:�I�:v��:��:�5g:��H:��*:|:r�9)W�9��W9��8W�-�����#i�X���������x&���@��J[��hu�ͫ��,���'Y��n�������IǺ��Ӻ >�x��3���!��U�����8����� ���&���,���2���8���>�\�D��J���P��V��x\��_b�Eh��)n��t���y�q��N܂�΅�����2���˦��������������~|���  �  Lr==��=T=Q�=F�=�3=d� =�r =X =�_�<��<���<U�<LL�<i��<���<���<!+�<N`�<e��<]��<��<�)�<�X�<���<��<���<"�<�.�<�T�<�x�<r��<���<��<��<\�<�)�<a?�<�R�<�c�<wr�<W~�<~��<ݍ�<E��<Ǒ�<&��<Z��<T��<�s�<#d�<�P�<�9�<;�<� �<���<^��<2��<�_�<�-�<���<��<�|�<{9�<���<\��<�T�<���<��<�G�<d��<e~�<�<N��<1/�<˶�<:�<:��<74�<��<�<��<3��<�_�<Ví<�#�<9��<�٨<�/�<���<�ң<��<�i�<[��<J��<�8�<�x�<̶�<��<k,�<Zd�<x��<�Ύ<��<{3�<�c�<ɒ�<���<��<��<3E�<��|<24y<��u<��q< -n<Bj<��f<$c<$w_<��[<FX< uT<�P<�$M<�~I<3�E<�9B<��><�:<hd7<��3<�:0<�,<B)<[�%<�"<|�<�<m�<4<��<�c<�
<?�<�V<
 <��;�	�;2��;�7�;���;���;�m�;GJ�;�6�;,4�;gB�;�a�;���;�ԩ;)�;뎞;��;��;)-�;tۈ;ڛ�;��|;��r;�h;d�^;3�T;E.K;ЧA;�C8;G/;��%;��;��;O<;��;�)�:�Z�:��:|e�:+=�:fI�:ӈ�:���:$4g:2�H:�*:4:dt�9Z�9�W9��8��-�����i�gW��f�����Y|&�z�@��I[�Egu�����ь��OY�����ն���JǺ��Ӻ#?຦�캒�����������7��3��4� ���&���,���2�R�8���>���D�κJ���P���V��x\�Q_b��Dh�y)n�Ct���y����%܂�5΅�i���Y�����������ݏ��b���r|���  �  Mr==��=T=O�=E�=�3=n� =�r =` =�_�<���<���<W�<WL�<g��<���<���<+�<Y`�<f��<r��<��<�)�<�X�<���<��<���< �<�.�<�T�<y�<{��<��<w��<��<M�<�)�<c?�<�R�<�c�<hr�<Y~�<t��<ߍ�<?��<ʑ�<$��<l��<_��<�s�<1d�<�P�<�9�<=�<� �<���<_��<6��<�_�<�-�<���<��<}�<z9�<���<R��<�T�<���<��<�G�<S��<n~�<�<R��<#/�<̶�<:�</��<A4�<��<�<�<,��<�_�<Qí<�#�<.��<�٨<�/�<���<�ң<��<�i�<Q��<S��<�8�<�x�<Ѷ�<��<j,�<Od�<���<�Ύ<�<�3�<�c�<Ȓ�<���<��<��<6E�<��|<%4y<��u<��q<�,n<)j<��f<$c<w_<��[<\X<uT<��P<�$M<�~I<5�E<�9B<��><�:<{d7<�3<�:0</�,<0)<X�%<�"<��<<i�<4<��<}c<�
<A�<!W<
 <��;Z	�;,��;�7�;���;���;qm�;PJ�;�6�;P4�;>B�;�a�;���;�ԩ;)�;�;��;萓;�,�;}ۈ;���;��|;m�r;
�h;Z�^;��T;�.K;��A;	D8;� /;��%;��;�;�<;��;�)�:�Y�:���:f�:�=�:�J�:���:C��:�2g:I�H:�*:�:�p�9�U�9�W9��8]�-�3	��Li��X���ṑ���{&���@��L[�(hu��������qY����������JǺe�Ӻ�>���v���_�������������� ���&��,���2�[�8�j�>���D�ѺJ���P�אV��x\��_b��Dh�,*n�wt�6�y����'܂�g΅�K�������������������n����|���  �  Lr==��=#T=S�=D�=�3=c� =�r =^ =�_�<��<���<Z�<TL�<n��<���<���<+�<X`�<k��<]��<��<�)�<�X�<���<��<���< �<�.�<�T�<y�<o��<��<���<���<\�<�)�<Z?�<�R�<�c�<qr�<V~�<s��<؍�<P��<ɑ�<$��<g��<U��<�s�<*d�<�P�<�9�<B�<� �<���<g��<3��<�_�<�-�<���<��<�|�<z9�<���<a��<�T�<}��<��<�G�<Z��<a~�< �<G��<//�<���<:�<8��<44�<��<�<��<.��<�_�<Jí<�#�<<��<�٨<�/�<���<�ң<��<�i�<f��<L��<�8�<�x�<Ҷ�<��<r,�<Vd�<���<�Ύ<��<�3�<�c�<̒�<���<��<��<0E�<��|<4y<��u<r�q<�,n<Ej<q�f<!$c<w_<��[<VX<
uT<�P<�$M<�~I<(�E<�9B<��><�:<}d7<��3<�:0<)�,<;)<r�%<�"<��<<x�<4<�<�c<�
<K�<�V<%
 <��;�	�;V��;x7�;���;���;�m�;J�;�6�;!4�;^B�;�a�;`��;�ԩ;�(�;ώ�;��;;-�;pۈ;���;��|;��r; �h;X�^;��T;L.K;2�A;�C8;F/;��%;�;��;k<;Ι;�)�:�Z�:���:nf�:S=�:J�:ƈ�:���:�4g:��H:��*::�r�9�W�9��W9���8�-�h���xi�
X�����$���{&���@��J[��gu�꫇�����Y�����󶺺�JǺ��Ӻ�>���캉�����������	�����	� �W�&���,�!�2�<�8��>�~�D�غJ���P�H�V��x\��_b��Dh��)n��t�b�y����1܂�.΅�����K�������ښ�����������|���  �  Br==��=T=P�=G�=�3=b� =�r =[ =�_�<��<���<i�<JL�<}��<���<���<+�<W`�<w��<\��<)��<�)�<�X�<���<��<���<�<�.�<�T�<y�<i��<��<~��<���<`�<r)�<d?�<�R�<�c�<pr�<O~�<���<э�<H��<�<-��<g��<V��<t�<$d�<�P�<�9�<G�<� �<���<o��<,��<�_�<�-�< ��<��<�|�<�9�<���<[��<�T�<���<��<�G�<\��<Y~�<�<7��<1/�<���<:�<3��<*4�<��<��<��<!��<�_�<Rí<}#�<7��<�٨<�/�<���<�ң<��<�i�<e��<D��<�8�<�x�<޶�<��<n,�<]d�<}��<ώ<��<�3�<�c�<Œ�<���<��<��< E�<��|<4y<��u<�q<�,n<Lj<k�f<&$c<w_<��[<RX<�tT<�P<$M<�~I<*�E<�9B<��><�:<�d7<��3<�:0<�,<F)<j�%<�"<��<�<��<�3<�<�c<�
<c�<�V<=
 <���;~	�;'��;�7�;���;D��;�m�;�I�;�6�;4�;BB�;�a�;S��;�ԩ;�(�;���;��;�;-�;Tۈ;;��|;��r;ɒh;��^;��T;[.K;~�A;�C8;�/;��%;/�;)�;�<;�;B)�:>[�:&��:�f�:�=�:J�:���:���:$4g:��H:y�*:�:~q�9EX�9c�W9R��8 a.�����i�!Y��ū�g���z&���@��I[�uiu���������Y�����R����IǺ��Ӻ3>�ڠ캛������0��H��9�����
� �x�&���,�Z�2���8��>�^�D���J���P���V��x\�-_b�BEh�u)n��t�z�y����t܂�!΅�����B���즎�Ϛ��ŏ������o|���  �  Cr==��=!T=V�=E�=�3=l� =�r =_ =�_�<��<���<h�<NL�<z��<���<���<"+�<Z`�<q��<j��<��<�)�<�X�<���<��<���<�<�.�<�T�<�x�<l��<��<s��<���<R�<z)�<d?�<�R�<�c�<hr�<O~�<s��<׍�<M��<ˑ�<#��<d��<a��< t�<-d�<�P�<�9�<I�<� �<���<n��<:��<�_�<�-�<���<"��<�|�<x9�<���<`��<�T�<}��<��<�G�<X��<_~�<�<>��<&/�<���<:�<0��<.4�<��< �<���<��<�_�<Ií<�#�<@��<�٨<�/�<���<�ң<��<�i�<[��<V��<�8�<�x�<߶�<��<s,�<Zd�<���<ώ<�<3�<�c�<ђ�<���<��<��<"E�<��|<4y<��u<��q<�,n</j<��f<$c<w_<��[<HX<uT<��P<�$M<�~I<#�E<�9B<��><�:<nd7<�3<�:0<,�,<G)<i�%<�"<��<<��<4<��<�c<�
<Y�<W<
 <��;�	�;H��;u7�;���;A��;�m�;J�;�6�;4�;>B�;�a�;a��;�ԩ;�(�;���;��;琓;�,�;Tۈ;���;��|;�r;�h;W�^;��T;�.K;J�A;�C8;A/;�%;D�;T�;�<;�;,*�:�Z�:���:f�:	>�:7J�:���:)��:�4g:��H:��*:�:6p�9W�9��W9��8�&.�A���i�K[���������{&�!�@�;K[��iu���������/Y��c��߶���JǺ�ӺG>�۠�]��������l��������� �N�&���,��2� �8�s�>���D�ɺJ�b�P�k�V��x\��_b�6Eh��)n��t���y����a܂�[΅���������㦎�����ُ�������|���  �  Nr==��=T=N�=I�=�3=m� =�r =d =�_�<��<���<[�<kL�<k��<���<���<)+�<]`�<b��<p��<��<�)�<�X�<���<��<���< �<�.�<�T�<�x�<f��<��<t��<���<I�<�)�<O?�<�R�<�c�<gr�<`~�<r��<ݍ�<>��<Ǒ�<)��<h��<^��<�s�<;d�<�P�<�9�<>�<� �<���<b��<F��<�_�<�-�<���<��<}�<}9�<���<P��<�T�<}��<���<�G�<R��<b~�<��<C��</�<���<:�<-��<+4�<��<�<���<+��<�_�<Jí<�#�<-��<�٨<�/�<���<�ң<��<�i�<e��<]��<�8�< y�<ն�<��<,�<[d�<���<�Ύ<�<�3�<�c�<Œ�<���<��<��<7E�<��|<4y<��u<]�q<�,n<!j<��f<�#c<w_<��[<?X<uT<��P<�$M<�~I<'�E<�9B<��>< �:<vd7<�3<�:0<B�,<J)<��%<�"<��<=<q�<&4<�<�c<�
<<�<W<#
 <'��;[	�;A��;z7�;���;���;�m�;*J�;�6�;�3�;BB�;�a�;j��;�ԩ;�(�;���;��;ᐓ;�,�;�ۈ;���;��|;j�r;��h;��^;��T;�.K;֧A;bD8;C/;z�%;��;b�;=;��;�*�:�Z�:���:�e�:�=�:fJ�:���:0��:�2g:L�H:��*:X:Eq�9�U�9��W9���8%�-�"��i��Z����$���}&�:�@��K[�(hu�z���q���0Y�����q����JǺ��Ӻ�>�Ԡ��������e�����V������� ���&���,���2���8�q�>���D���J���P�אV��x\��_b��Dh� *n��t���y�K��B܂�u΅���������̦������ꏔ������|���  �  Dr==��=T=O�=H�=�3=l� =�r =e =�_�<��<���<d�<fL�<x��<���<���<+�<e`�<w��<m��<%��<�)�<�X�<���<��<���<�<�.�<�T�<y�<g��<��<m��<���<K�<w)�<Z?�<�R�<�c�<cr�<J~�<r��<ٍ�<J��<ɑ�</��<h��<g��<	t�<6d�<�P�<�9�<J�<� �<���<o��<@��<�_�<�-�<��<(��<�|�<�9�<���<\��<�T�<~��<��<�G�<H��<W~�<��<<��</�<���<:�<)��<*4�<��<��<���<��<�_�<Kí<�#�<2��<�٨<�/�<���<�ң<��<�i�<c��<Z��<�8�<�x�<ܶ�<��<w,�<Rd�<���<ώ<�<�3�<�c�<ƒ�<���<��<��<"E�<��|<4y<��u<j�q<�,n<$j<n�f<�#c<w_<��[<QX<�tT<��P<�$M<�~I<)�E<�9B<��><�:<�d7<�3<�:0<D�,<7)<u�%<�"<��<1<��<$4<�<�c<	
<f�<W<6
 <%��;q	�;:��;z7�;���;P��;�m�;�I�;�6�;4�;*B�;�a�;M��;�ԩ;�(�;Ў�;��;���;�,�;Aۈ;���;��|;ѥr;�h;��^;��T;�.K;��A;7D8;3/;/�%;J�;�;
=;�;�*�:�Z�:���:g�:l>�:GJ�:g��:2��:[4g:��H:��*:�:To�9jS�9R�W9���8E,.�A��ki�Z\����8���{&��@�ML[��iu�|���f���mY��4������
JǺ��Ӻ�=���u���ɝ���n��q������� �2�&��,���2���8�q�>�i�D���J���P���V��x\��_b�4Eh� *n��t�m�y���c܂�q΅���������覎��Ə��Å���|���  �  Cr==��=T=V�=D�=�3=f� =�r =^ =�_�<��<���<m�<QL�<���<���<���</+�<Z`�<q��<_��<��<�)�<�X�<���<��<���<�<�.�<�T�<�x�<X��<��<q��<���<V�<l)�<X?�<�R�<�c�<tr�<G~�<���<̍�<S��<ȑ�<*��<d��<]��< t�<,d�<�P�<�9�<M�<� �<���<s��<9��<	`�<�-�<���<��<�|�<9�<���<h��<�T�<���<��<�G�<R��<S~�<��<.��<&/�<���<	:�<-��<4�<��<��<��<$��<�_�<Oí<w#�<H��<�٨<�/�<���<�ң<��<�i�<q��<P��<�8�<�x�<㶗<��<x,�<ld�<���<	ώ<��<�3�<�c�<ђ�<���<��<��<E�<��|<�3y<|�u<a�q<�,n<4j<l�f<
$c<w_<��[<@X<�tT<�P<�$M<�~I<�E<�9B<��><�:<{d7<��3<�:0<)�,<i)<z�%<�"<��<<��<4<$�<�c<�
<Y�<�V<*
 <��;�	�;*��;|7�;���;S��;�m�;�I�;�6�;�3�;:B�;�a�;V��;�ԩ;�(�;ˎ�;��;ϐ�;"-�;:ۈ;ꛃ;h�|;�r;�h;��^;��T;�.K;K�A;�C8;/;�%;h�;Q�;�<;7�;"*�:#\�:���:{f�:�=�:�I�:$��:���:�5g:��H:]�*:�:�r�9�U�9�W9O��8�.�[��|i�{[����L��L|&�[�@�_J[� iu�˫��"����Y��������dJǺ��Ӻq>�Ӡ�����W��ͺ�*��	��w���� �*�&�.�,�0�2���8���>���D�ԺJ�\�P�{�V��x\�*_b�HEh�s)n�t���y�;��x܂�Q΅�����y���즎����揔�΅��m|���  �  Ar==��=T=R�=G�=�3=l� =�r =a =�_�<��<���<t�<jL�<���<���<���<-+�<_`�<v��<n��<+��<�)�<�X�<���<��<���<�<�.�<�T�<�x�<b��<��<g��<���<C�<v)�<S?�<�R�<�c�<er�<F~�<}��<ύ�<F��<ő�<1��<t��<i��<t�<3d�<�P�<�9�<H�<� �<���<q��<5��<`�<�-�< ��<+��<}�<�9�<���<Y��<�T�<���<ߥ�<�G�<D��<]~�<��<:��</�<���<:�<'��<&4�<��<��<�<��<�_�<Lí<w#�<6��<�٨<�/�<���<�ң<��<�i�<m��<N��<�8�<y�<궗<��<u,�<hd�<���<ώ<�<�3�<�c�<˒�<���<��<��<E�<��|<�3y<��u<b�q<�,n<j<d�f<�#c<w_<��[<KX<�tT<��P<{$M<�~I<�E<�9B<��><�:<�d7<�3<�:0<3�,<^)<r�%<�"<��<;<��<4<�<�c< 
<e�<W<C
 <��;�	�;$��;w7�;���;C��;�m�;�I�;�6�;�3�;6B�;pa�;<��;�ԩ;�(�;���;��;���;�,�;4ۈ;ܛ�;��|;��r;�h;ƣ^;�T;�.K;x�A;&D8;�/;�%;=�;��;7=;!�;�)�:�[�:0��:�f�:�>�:K�:���:���:4g:d�H:��*:p:�o�9�R�9��W9ˡ�8�=.����� i�a]����ṷ��c|&�q�@��L[�ju�*���Q����Y���������IǺ��Ӻ�=�c�캰���{��޺�#��D��A���� �?�&�U�,��2���8�u�>�!�D���J���P�ɐV��x\�`_b�VEh��)n�t���y�5��`܂��΅���������ߦ�� ���ҏ��ǅ���|���  �  Hr==��="T=R�=F�=�3=e� =�r =d =�_�<��<���<c�<XL�<t��<���<���< +�<d`�<p��<\��<��<�)�<�X�<���<��<���<!�<�.�<�T�<�x�<d��<��<n��<���<A�<)�<H?�<�R�<�c�<qr�<P~�<n��<ڍ�<M��<ʑ�<$��<Z��<Y��<t�<4d�<�P�<�9�<N�<� �<���<r��<I��<�_�<�-�<���<��<�|�<y9�<���<^��<�T�<|��<��<�G�<M��<d~�<��<C��</�<���<
:�<��<*4�<��<��<���<1��<�_�<Jí<�#�<6��<�٨<�/�<���<�ң<��<�i�<k��<^��<�8�<�x�<׶�<��<�,�<Yd�<���<
ώ<��<3�<�c�<˒�<���<��<��<)E�<��|<4y<��u<T�q<�,n<j<��f<�#c<w_<��[<EX<�tT<��P<�$M<�~I<1�E<�9B<��><�:<sd7<��3<�:0<B�,<@)<��%<�"<��<<��<34<&�<�c<
<W�<�V<*
 <!��;�	�;i��;z7�;���;���;�m�;�I�;�6�;�3�;B�;�a�;���;�ԩ;�(�;���;��;ǐ�;-�;^ۈ;���;��|;�r;�h;_�^;B�T;w.K;`�A;*D8;c/;��%;o�;X�;�<;*�;,+�:5[�:���:�f�:�=�:WI�:�:+��:�4g:E�H:��*::t�9�T�9��W9��8U�-����Ji�Q[�����?��~&�R�@��K[�Qgu�U���r����X���������[JǺ��Ӻ�>�6��E������]�����������p� ���&���,���2���8���>���D�ߺJ���P�]�V��x\��_b��Dh��)n��t���y�p��U܂��΅�w�������禎����ݏ�������|���  �  Ar==��=T=R�=G�=�3=l� =�r =a =�_�<��<���<t�<jL�<���<���<���<-+�<_`�<v��<n��<+��<�)�<�X�<���<��<���<�<�.�<�T�<�x�<b��<��<g��<���<C�<v)�<S?�<�R�<�c�<er�<F~�<}��<ύ�<F��<ő�<1��<t��<i��<t�<3d�<�P�<�9�<H�<� �<���<q��<5��<`�<�-�< ��<+��<}�<�9�<���<Y��<�T�<���<ߥ�<�G�<D��<]~�<��<:��</�<���<:�<'��<&4�<��<��<�<��<�_�<Lí<w#�<6��<�٨<�/�<���<�ң<��<�i�<m��<N��<�8�<y�<궗<��<u,�<hd�<���<ώ<�<�3�<�c�<˒�<���<��<��<E�<��|<�3y<��u<b�q<�,n<j<d�f<�#c<w_<��[<KX<�tT<��P<{$M<�~I<�E<�9B<��><�:<�d7<�3<�:0<3�,<^)<r�%<�"<��<;<��<4<�<�c< 
<e�<W<C
 <��;�	�;$��;w7�;���;C��;�m�;�I�;�6�;�3�;6B�;pa�;<��;�ԩ;�(�;���;��;���;�,�;4ۈ;ܛ�;��|;��r;�h;ƣ^;�T;�.K;x�A;&D8;�/;�%;=�;��;7=;!�;�)�:�[�:0��:�f�:�>�:K�:���:���:4g:d�H:��*:p:�o�9�R�9��W9ˡ�8�=.����� i�a]����ṷ��c|&�q�@��L[�ju�*���Q����Y���������IǺ��Ӻ�=�c�캰���{��޺�#��D��A���� �?�&�U�,��2���8�u�>�!�D���J���P�ɐV��x\�`_b�VEh��)n�t���y�5��`܂��΅���������ߦ�� ���ҏ��ǅ���|���  �  Cr==��=T=V�=D�=�3=f� =�r =^ =�_�<��<���<m�<QL�<���<���<���</+�<Z`�<q��<_��<��<�)�<�X�<���<��<���<�<�.�<�T�<�x�<X��<��<q��<���<V�<l)�<X?�<�R�<�c�<tr�<G~�<���<̍�<S��<ȑ�<*��<d��<]��< t�<,d�<�P�<�9�<M�<� �<���<s��<9��<	`�<�-�<���<��<�|�<9�<���<h��<�T�<���<��<�G�<R��<S~�<��<.��<&/�<���<	:�<-��<4�<��<��<��<$��<�_�<Oí<w#�<H��<�٨<�/�<���<�ң<��<�i�<q��<P��<�8�<�x�<㶗<��<x,�<ld�<���<	ώ<��<�3�<�c�<ђ�<���<��<��<E�<��|<�3y<|�u<a�q<�,n<4j<l�f<
$c<w_<��[<@X<�tT<�P<�$M<�~I<�E<�9B<��><�:<{d7<��3<�:0<)�,<i)<z�%<�"<��<<��<4<$�<�c<�
<Y�<�V<*
 <��;�	�;*��;|7�;���;S��;�m�;�I�;�6�;�3�;:B�;�a�;V��;�ԩ;�(�;ˎ�;��;ϐ�;"-�;:ۈ;ꛃ;h�|;�r;�h;��^;��T;�.K;K�A;�C8;/;�%;h�;Q�;�<;7�;"*�:#\�:���:{f�:�=�:�I�:$��:���:�5g:��H:]�*:�:�r�9�U�9�W9O��8�.�[��|i�{[����L��L|&�[�@�_J[� iu�˫��"����Y��������dJǺ��Ӻq>�Ӡ�����W��ͺ�*��	��w���� �*�&�.�,�0�2���8���>���D�ԺJ�\�P�{�V��x\�*_b�HEh�s)n�t���y�;��x܂�Q΅�����y���즎����揔�΅��m|���  �  Dr==��=T=O�=H�=�3=l� =�r =e =�_�<��<���<d�<fL�<x��<���<���<+�<e`�<w��<m��<%��<�)�<�X�<���<��<���<�<�.�<�T�<y�<g��<��<m��<���<K�<w)�<Z?�<�R�<�c�<cr�<J~�<r��<ٍ�<J��<ɑ�</��<h��<g��<	t�<6d�<�P�<�9�<J�<� �<���<o��<@��<�_�<�-�<��<(��<�|�<�9�<���<\��<�T�<~��<��<�G�<H��<W~�<��<<��</�<���<:�<)��<*4�<��<��<���<��<�_�<Kí<�#�<2��<�٨<�/�<���<�ң<��<�i�<c��<Z��<�8�<�x�<ܶ�<��<w,�<Rd�<���<ώ<�<�3�<�c�<ƒ�<���<��<��<"E�<��|<4y<��u<j�q<�,n<$j<n�f<�#c<w_<��[<QX<�tT<��P<�$M<�~I<)�E<�9B<��><�:<�d7<�3<�:0<D�,<7)<u�%<�"<��<1<��<$4<�<�c<	
<f�<W<6
 <%��;q	�;:��;z7�;���;P��;�m�;�I�;�6�;4�;*B�;�a�;M��;�ԩ;�(�;Ў�;��;���;�,�;Aۈ;���;��|;ѥr;�h;��^;��T;�.K;��A;7D8;3/;/�%;J�;�;
=;�;�*�:�Z�:���:g�:l>�:GJ�:g��:2��:[4g:��H:��*:�:To�9jS�9R�W9���8E,.�A��ki�Z\����8���{&��@�ML[��iu�|���f���mY��4������
JǺ��Ӻ�=���u���ɝ���n��q������� �2�&��,���2���8�q�>�i�D���J���P���V��x\��_b�4Eh� *n��t�m�y���c܂�q΅���������覎��Ə��Å���|���  �  Nr==��=T=N�=I�=�3=m� =�r =d =�_�<��<���<[�<kL�<k��<���<���<)+�<]`�<b��<p��<��<�)�<�X�<���<��<���< �<�.�<�T�<�x�<f��<��<t��<���<I�<�)�<O?�<�R�<�c�<gr�<`~�<r��<ݍ�<>��<Ǒ�<)��<h��<^��<�s�<;d�<�P�<�9�<>�<� �<���<b��<F��<�_�<�-�<���<��<}�<}9�<���<P��<�T�<}��<���<�G�<R��<b~�<��<C��</�<���<:�<-��<+4�<��<�<���<+��<�_�<Jí<�#�<-��<�٨<�/�<���<�ң<��<�i�<e��<]��<�8�< y�<ն�<��<,�<[d�<���<�Ύ<�<�3�<�c�<Œ�<���<��<��<7E�<��|<4y<��u<]�q<�,n<!j<��f<�#c<w_<��[<?X<uT<��P<�$M<�~I<'�E<�9B<��>< �:<vd7<�3<�:0<B�,<J)<��%<�"<��<=<q�<&4<�<�c<�
<<�<W<#
 <'��;[	�;A��;z7�;���;���;�m�;*J�;�6�;�3�;BB�;�a�;j��;�ԩ;�(�;���;��;ᐓ;�,�;�ۈ;���;��|;j�r;��h;��^;��T;�.K;֧A;bD8;C/;z�%;��;b�;=;��;�*�:�Z�:���:�e�:�=�:fJ�:���:0��:�2g:L�H:��*:X:Eq�9�U�9��W9���8%�-�"��i��Z����$���}&�:�@��K[�(hu�z���q���0Y�����q����JǺ��Ӻ�>�Ԡ��������e�����V������� ���&���,���2���8�q�>���D���J���P�אV��x\��_b��Dh� *n��t���y�K��B܂�u΅���������̦������ꏔ������|���  �  Cr==��=!T=V�=E�=�3=l� =�r =_ =�_�<��<���<h�<NL�<z��<���<���<"+�<Z`�<q��<j��<��<�)�<�X�<���<��<���<�<�.�<�T�<�x�<l��<��<s��<���<R�<z)�<d?�<�R�<�c�<hr�<O~�<s��<׍�<M��<ˑ�<#��<d��<a��< t�<-d�<�P�<�9�<I�<� �<���<n��<:��<�_�<�-�<���<"��<�|�<x9�<���<`��<�T�<}��<��<�G�<X��<_~�<�<>��<&/�<���<:�<0��<.4�<��< �<���<��<�_�<Ií<�#�<@��<�٨<�/�<���<�ң<��<�i�<[��<V��<�8�<�x�<߶�<��<s,�<Zd�<���<ώ<�<3�<�c�<ђ�<���<��<��<"E�<��|<4y<��u<��q<�,n</j<��f<$c<w_<��[<HX<uT<��P<�$M<�~I<#�E<�9B<��><�:<nd7<�3<�:0<,�,<G)<i�%<�"<��<<��<4<��<�c<�
<Y�<W<
 <��;�	�;H��;u7�;���;A��;�m�;J�;�6�;4�;>B�;�a�;a��;�ԩ;�(�;���;��;琓;�,�;Tۈ;���;��|;�r;�h;W�^;��T;�.K;J�A;�C8;A/;�%;D�;T�;�<;�;,*�:�Z�:���:f�:	>�:7J�:���:)��:�4g:��H:��*:�:6p�9W�9��W9��8�&.�A���i�K[���������{&�!�@�;K[��iu���������/Y��c��߶���JǺ�ӺG>�۠�]��������l��������� �N�&���,��2� �8�s�>���D�ɺJ�b�P�k�V��x\��_b�6Eh��)n��t���y����a܂�[΅���������㦎�����ُ�������|���  �  Br==��=T=P�=G�=�3=b� =�r =[ =�_�<��<���<i�<JL�<}��<���<���<+�<W`�<w��<\��<)��<�)�<�X�<���<��<���<�<�.�<�T�<y�<i��<��<~��<���<`�<r)�<d?�<�R�<�c�<pr�<O~�<���<э�<H��<�<-��<g��<V��<t�<$d�<�P�<�9�<G�<� �<���<o��<,��<�_�<�-�< ��<��<�|�<�9�<���<[��<�T�<���<��<�G�<\��<Y~�<�<7��<1/�<���<:�<3��<*4�<��<��<��<!��<�_�<Rí<}#�<7��<�٨<�/�<���<�ң<��<�i�<e��<D��<�8�<�x�<޶�<��<n,�<]d�<}��<ώ<��<�3�<�c�<Œ�<���<��<��< E�<��|<4y<��u<�q<�,n<Lj<k�f<&$c<w_<��[<RX<�tT<�P<$M<�~I<*�E<�9B<��><�:<�d7<��3<�:0<�,<F)<j�%<�"<��<�<��<�3<�<�c<�
<c�<�V<=
 <���;~	�;'��;�7�;���;D��;�m�;�I�;�6�;4�;BB�;�a�;S��;�ԩ;�(�;���;��;�;-�;Tۈ;;��|;��r;ɒh;��^;��T;[.K;~�A;�C8;�/;��%;/�;)�;�<;�;B)�:>[�:&��:�f�:�=�:J�:���:���:$4g:��H:y�*:�:~q�9EX�9c�W9R��8 a.�����i�!Y��ū�g���z&���@��I[�uiu���������Y�����R����IǺ��Ӻ3>�ڠ캛������0��H��9�����
� �x�&���,�Z�2���8��>�^�D���J���P���V��x\�-_b�BEh�u)n��t�z�y����t܂�!΅�����B���즎�Ϛ��ŏ������o|���  �  Lr==��=#T=S�=D�=�3=c� =�r =^ =�_�<��<���<Z�<TL�<n��<���<���<+�<X`�<k��<]��<��<�)�<�X�<���<��<���< �<�.�<�T�<y�<o��<��<���<���<\�<�)�<Z?�<�R�<�c�<qr�<V~�<s��<؍�<P��<ɑ�<$��<g��<U��<�s�<*d�<�P�<�9�<B�<� �<���<g��<3��<�_�<�-�<���<��<�|�<z9�<���<a��<�T�<}��<��<�G�<Z��<a~�< �<G��<//�<���<:�<8��<44�<��<�<��<.��<�_�<Jí<�#�<<��<�٨<�/�<���<�ң<��<�i�<f��<L��<�8�<�x�<Ҷ�<��<r,�<Vd�<���<�Ύ<��<�3�<�c�<̒�<���<��<��<0E�<��|<4y<��u<r�q<�,n<Ej<q�f<!$c<w_<��[<VX<
uT<�P<�$M<�~I<(�E<�9B<��><�:<}d7<��3<�:0<)�,<;)<r�%<�"<��<<x�<4<�<�c<�
<K�<�V<%
 <��;�	�;V��;x7�;���;���;�m�;J�;�6�;!4�;^B�;�a�;`��;�ԩ;�(�;ώ�;��;;-�;pۈ;���;��|;��r; �h;X�^;��T;L.K;2�A;�C8;F/;��%;�;��;k<;Ι;�)�:�Z�:���:nf�:S=�:J�:ƈ�:���:�4g:��H:��*::�r�9�W�9��W9���8�-�h���xi�
X�����$���{&���@��J[��gu�꫇�����Y�����󶺺�JǺ��Ӻ�>���캉�����������	�����	� �W�&���,�!�2�<�8��>�~�D�غJ���P�H�V��x\��_b��Dh��)n��t�b�y����1܂�.΅�����K�������ښ�����������|���  �  Mr==��=T=O�=E�=�3=n� =�r =` =�_�<���<���<W�<WL�<g��<���<���<+�<Y`�<f��<r��<��<�)�<�X�<���<��<���< �<�.�<�T�<y�<{��<��<w��<��<M�<�)�<c?�<�R�<�c�<hr�<Y~�<t��<ߍ�<?��<ʑ�<$��<l��<_��<�s�<1d�<�P�<�9�<=�<� �<���<_��<6��<�_�<�-�<���<��<}�<z9�<���<R��<�T�<���<��<�G�<S��<n~�<�<R��<#/�<̶�<:�</��<A4�<��<�<�<,��<�_�<Qí<�#�<.��<�٨<�/�<���<�ң<��<�i�<Q��<S��<�8�<�x�<Ѷ�<��<j,�<Od�<���<�Ύ<�<�3�<�c�<Ȓ�<���<��<��<6E�<��|<%4y<��u<��q<�,n<)j<��f<$c<w_<��[<\X<uT<��P<�$M<�~I<5�E<�9B<��><�:<{d7<�3<�:0</�,<0)<X�%<�"<��<<i�<4<��<}c<�
<A�<!W<
 <��;Z	�;,��;�7�;���;���;qm�;PJ�;�6�;P4�;>B�;�a�;���;�ԩ;)�;�;��;萓;�,�;}ۈ;���;��|;m�r;
�h;Z�^;��T;�.K;��A;	D8;� /;��%;��;�;�<;��;�)�:�Y�:���:f�:�=�:�J�:���:C��:�2g:I�H:�*:�:�p�9�U�9�W9��8]�-�3	��Li��X���ṑ���{&���@��L[�(hu��������qY����������JǺe�Ӻ�>���v���_�������������� ���&��,���2�[�8�j�>���D�ѺJ���P�אV��x\��_b��Dh�,*n�wt�6�y����'܂�g΅�K�������������������n����|���  �  Lr==��=T=Q�=F�=�3=d� =�r =X =�_�<��<���<U�<LL�<i��<���<���<!+�<N`�<e��<]��<��<�)�<�X�<���<��<���<"�<�.�<�T�<�x�<r��<���<��<��<\�<�)�<a?�<�R�<�c�<wr�<W~�<~��<ݍ�<E��<Ǒ�<&��<Z��<T��<�s�<#d�<�P�<�9�<;�<� �<���<^��<2��<�_�<�-�<���<��<�|�<{9�<���<\��<�T�<���<��<�G�<d��<e~�<�<N��<1/�<˶�<:�<:��<74�<��<�<��<3��<�_�<Ví<�#�<9��<�٨<�/�<���<�ң<��<�i�<[��<J��<�8�<�x�<̶�<��<k,�<Zd�<x��<�Ύ<��<{3�<�c�<ɒ�<���<��<��<3E�<��|<24y<��u<��q< -n<Bj<��f<$c<$w_<��[<FX< uT<�P<�$M<�~I<3�E<�9B<��><�:<hd7<��3<�:0<�,<B)<[�%<�"<|�<�<m�<4<��<�c<�
<?�<�V<
 <��;�	�;2��;�7�;���;���;�m�;GJ�;�6�;,4�;gB�;�a�;���;�ԩ;)�;뎞;��;��;)-�;tۈ;ڛ�;��|;��r;�h;d�^;3�T;E.K;ЧA;�C8;G/;��%;��;��;O<;��;�)�:�Z�:��:|e�:+=�:fI�:ӈ�:���:$4g:2�H:�*:4:dt�9Z�9�W9��8��-�����i�gW��f�����Y|&�z�@��I[�Egu�����ь��OY�����ն���JǺ��Ӻ#?຦�캒�����������7��3��4� ���&���,���2�R�8���>���D�κJ���P���V��x\�Q_b��Dh�y)n�Ct���y����%܂�5΅�i���Y�����������ݏ��b���r|���  �  Er==��=%T=Q�=B�=�3=c� =�r =W =�_�<���<���<[�<JL�<r��<���<���<+�<L`�<w��<Z��<*��<�)�<�X�<���<��<���<�<�.�<�T�<y�<r��<���<���<���<c�<)�<r?�<�R�<�c�<nr�<O~�<y��<֍�<Y��<���<,��<b��<[��<t�<!d�<�P�<�9�<@�<� �<���<f��<#��<�_�<�-�<���<!��<�|�<�9�<���<j��<�T�<���<��<�G�<Y��<d~�<�<E��<6/�<���<:�<=��<64�<.��<�<��<(��<�_�<Pí<�#�<@��<�٨<�/�<���<�ң<��<�i�<Y��<?��<�8�<�x�<ж�<��<^,�<Sd�<v��<ώ<��<�3�<�c�<ƒ�<���<��<��<%E�<��|<4y<��u<��q<�,n<Wj<v�f<.$c<w_<��[<tX<uT<�P<�$M<�~I< �E<�9B<��><�:<�d7<��3<�:0<�,<3)<H�%<�"<��<�<~�<�3<��<qc<�
<c�<�V<<
 <��;�	�;V��;x7�;���;V��;�m�;J�;7�;,4�;eB�;�a�;b��;թ;�(�;+��;��;쐓;-�;Sۈ;ě�;��|;@�r;��h;��^;z�T;{.K;H�A;�C8;+/;H�%;��;��;n<;��;�(�:zZ�:���:8f�:�=�:�I�:v��:��:�5g:��H:��*:|:r�9)W�9��W9��8W�-�����#i�X���������x&���@��J[��hu�ͫ��,���'Y��n�������IǺ��Ӻ >�x��3���!��U�����8����� ���&���,���2���8���>�\�D��J���P��V��x\��_b�Eh��)n��t���y�q��N܂�΅�����2���˦��������������~|���  �  Lr==��= T=L�=C�=�3=b� =�r =Y =�_�<���<���<L�<GL�<^��<���<���<+�<J`�<g��<X��<#��<�)�<�X�<���<��<���<"�<�.�<�T�<y�<p��<��<���<
��<d�<|)�<l?�<�R�<�c�<xr�<_~�<���<֍�<H��<���<(��<]��<Q��<�s�<)d�<�P�<�9�<8�<� �<���<Y��</��<�_�<�-�<���<��<�|�<�9�<���<[��<�T�<���<���<�G�<`��<k~�<�<B��<5/�<Ѷ�<#:�<7��<44�<'��<
�<��<5��<�_�<Wí<�#�<5��<�٨<�/�<���<�ң<��<�i�<T��<H��<�8�<�x�<Ŷ�<��<g,�<Ud�<{��<�Ύ<��<�3�<�c�<���<���<��<��<3E�<��|<%4y<��u<��q<�,n<_j<��f<<$c<w_<��[<jX<uT<�P<�$M<�~I<+�E<�9B<y�><�:<�d7<��3<�:0<�,<<)<S�%<�"<k�<�<V�<4<��<�c<�
<B�<�V<.
 <��;d	�;>��;�7�;���;���;�m�;J�;�6�; 4�;KB�;�a�;���;	թ;�(�;��;��;��;.-�;�ۈ;;��|;��r;��h;w�^;M�T;(.K;��A;�C8;/;��%;��;��;:<;Z�;o)�:/Z�:���:Ge�:=�:uI�:B��:P��:4g:F�H:��*:�:u�9�X�9�W9˺�8.�u����i��U��0��9���y&��@��I[�gu�Ъ��Ì��eY��&��h���JǺ�Ӻ�>��캊���H����9��g��j��� ���&���,�c�2�b�8��>���D��J�ܦP���V��x\�&_b��Dh�~)n�wt��y����T܂��ͅ�X������Ҧ�������������w|���  �  �p=l=б=�Q=��=��=�0=� =�n =j =,W�<ߒ�<���<��<MA�<�y�<0��<���<2�<�Q�<���<(��<��<��<F�<s�<���<|��<���<��<�<�<�_�<m��<���<j��<���<>��<h
�<(�<�1�<�A�<�N�<�Y�<�a�<3g�<}i�<�h�<4e�<`^�<_T�<�F�<)6�<�!�<	
�<n��<<��<-��<��<OZ�<B+�<V��<+��<��<KF�<r�<Z��<�m�<$�<���<Pn�<[�<��<kG�<Tܿ<m�<l��<���<��<r��<<�<�x�<��<�\�<�Ȱ<w1�<\��<���<�U�<Q��<��<\�<e��<���<wG�<_��<�֜<��<�\�<⛗<2ٕ<��<�M�<���<Ȼ�<R��<Z#�<1U�<ʅ�<P��<��<|�<p>�<j�|<�,y<��u<��q<=/n<��j<��f<�/c<Ӆ_<��[<64X<�T<�P<�BM<!�I<��E<+aB<�><�+;<+�7<�4<�q0<&�,<E\)<�%<�V"<��<Rc<i�<�<�<3�<M[
<t<Գ<wi <�K�;��;�f�;�	�;��;�{�;�K�;%,�;��;��;�-�;IO�;E��;�ƪ;��;���;���;���;$�;]҉;m��;��~;3�t;�zj;g�`;ȸV;$M;ԀC;�:;��0;8�';A�;�;e�;!E;^r�:ؐ�:J��:${�:�A�:};�:2h�:ǅ:��l:�%N:d�/:�:�5�9Ѯ9
j9�E�8r��6.�Ӹ��X������#ڹB"�j�"���=��X��Ir��+�����d���c����q��^ƺ3�Һi!ߺZ�뺧����"��D�xb�Fx�p��� ���&���,��2�ȝ8�C�>�r�D�J��oP��]V�J\�6b��h��n���s���y����Ԃ�pȅ����ֱ������C���V������v����  �  �p=r=Ǳ=�Q=��=��=�0=� =�n =i =9W�<ْ�<���<��<4A�<�y�<%��<���<8�<�Q�<���< ��<��<��<F�<�r�<~��<���<���<��<�<�<�_�<c��<��<���<���<I��<Z
�<*�<�1�<�A�<O�<�Y�<�a�<g�<}i�<�h�<De�<k^�<UT�<�F�<,6�<�!�<�	�<p��<&��<��<#��<AZ�<U+�<Y��<%��<ۅ�<OF�<��<`��<�m�<�<���<Un�<_�<��<XG�<Xܿ<m�<t��<���<��<n��</�<�x�<��<�\�<�Ȱ<|1�<T��<���<�U�<X��<��<\�<a��<���<{G�<i��<�֜<��<n\�<ٛ�<1ٕ<��<N�<���<���<F��<n#�<<U�<΅�<G��<��<��<x>�<{�|<�,y<��u<��q<"/n<��j<
�f<�/c<��_<��[<64X< �T<,�P<�BM<8�I<��E<aB<)�><�+;<R�7<�4<�q0<&�,<_\)<s�%<�V"<��< c<w�<�<�<>�<K[
<r<ĳ<�i <�K�;<��;zf�;Z	�;��;�{�;�K�;�+�;��;\�;�-�;�O�;���;�ƪ;|�;˃�;���;|��;$�;x҉;���;��~;5�t;{j;�`;&�V;�M;��C;�:;k�0;Ƨ';N�;^�;��;HE;~q�:��:u��:�z�:TA�:�;�:Yi�:�ǅ:��l:�"N:~�/:I:�6�9�Ю9�
j9QJ�8��6��Ӹ�X�[����$ڹ�#���"��=��X��Hr�*+��t������뽬�;q��Gƺ��Һ�!ߺ���o���w"�3E�;b�y����� ��&�6�,��2��8���>�ԋD��~J�ioP�6^V��J\��5b�uh�{n�
�s���y����EԂ�+ȅ�����}���&���K���U���Q���M����  �  �p=u=Ǳ=�Q=��=|�=�0=
� =�n =e =8W�<֒�<���<��<5A�<�y�<��<���</�<�Q�<��<��<��<��<!F�<s�<���<���<���<��<�<�<`�<g��<��<t��<���<C��<S
�<;�<�1�<�A�<�N�<�Y�<�a�<g�<�i�<�h�<8e�<i^�<_T�<�F�<6�<�!�<�	�<���<6��<!��<7��<2Z�<Z+�<K��<4��<��<LF�<{�<T��<�m�<	�<���<Mn�<X�<��<SG�<iܿ<�l�<q��<���<��<o��</�<y�<��<�\�<�Ȱ<x1�<^��<���<�U�<G��<��<
\�<q��<���<oG�<r��<�֜<��<r\�<뛗<:ٕ<��<	N�<���<ϻ�<H��<j#�<+U�<υ�<V��<��<��<k>�<x�|<�,y<��u<��q</n<��j<��f<�/c<��_<��[<B4X<�T<,�P<�BM<A�I<��E<*aB<1�><�+;<J�7<�4<�q0<�,<]\)<m�%<�V"<��<#c<��<�<�<,�<K[
<�<��<�i <�K�;c��;�f�;u	�;��;�{�;L�;�+�;7�;m�;�-�;rO�;,��;�ƪ;`�;��;���;���;�#�;S҉;���;��~;��t;�zj;��`;�V;,M;�C;=:;��0;Z�';٠;۸;�;�E;�p�:g��:���:�{�:GB�:�;�:�h�:�ƅ:'�l:W"N:��/:R:�4�9
Ү9Yj9H[�8
`�6��Ӹ`�X�َ���$ڹ�#���"�,�=�!X��Ir�l+���������F���Er���ƺڢҺ� ߺ1��#���3"��E�za��x�*��ϖ �.�&�%�,�:�2���8���>��D�6J�coP��]V��J\�h5b��h��n��s���y�H��QԂ�Mȅ�$�������,���,���=���m���J����  �  �p=n=ɱ=�Q=��=��=�0=� =�n =g =8W�<��<���<��<1A�<�y�<!��<���<1�<�Q�<���<"��<��<��<F�<s�<���<y��<���<��<�<�<�_�<_��<��<z��<���<K��<Q
�<+�<�1�<�A�<�N�<�Y�<�a�<g�<i�<�h�<Ce�<i^�<WT�<�F�< 6�<�!�< 
�<r��<-��<��<%��<BZ�<Z+�<N��<4��<ޅ�<PF�<��<Z��<�m�<�<���<Mn�<Y�<��<YG�<Xܿ<�l�<v��<���<��<t��<)�<�x�<��<�\�<�Ȱ<q1�<Z��<���<�U�<P��<��<\�<a��<���<rG�<v��<�֜<��<l\�<ݛ�<2ٕ<��<N�<���<˻�<G��<i#�<7U�<˅�<N��<��<�<n>�<l�|<�,y<��u<��q<"/n<��j<��f<�/c<��_<��[<24X<�T<�P<�BM<&�I<��E< aB<&�><�+;<L�7<�4<�q0<�,<^\)<��%<�V"<��<c<|�<��<�<0�<U[
<u<ɳ<�i <�K�;3��;�f�;r	�;���;�{�;�K�;�+�;��;L�;�-�;�O�;���;�ƪ;[�;΃�;���;���;�#�;]҉;x��;��~;G�t;�zj;ۈ`;�V;�M;�C;K:;~�0;�';]�;��;��;ZE;�q�:`��:���:�{�:�A�:�;�:Xi�:%ǅ:(�l:�"N:B�/:Q:=5�9�Ѯ9nj91J�8�-�6L�Ӹ��X�����7#ڹ}$���"�؝=�X��Ir��+�������=����q��$ƺV�Һ�!ߺ������"�KE�#b�#y����� ���&�8�,�(�2���8���>���D��~J��oP��]V��J\��5b��h��n���s��y����DԂ�;ȅ������������`���]���B���j����  �  �p=k=̱=�Q=��=��=�0=� =�n =p =-W�<ߒ�<���<��<EA�<�y�<,��<���<.�<�Q�<��<*��<��<��<F�<s�<���<y��<���<��<�<�<�_�<k��<��<l��<���<4��<Z
�<+�<�1�<�A�<�N�<�Y�<�a�<-g�<|i�<�h�<9e�<k^�<VT�<�F�<26�<�!�<
�<s��<9��<)��<(��<JZ�<L+�<[��<4��<؅�<UF�<x�<a��<�m�<�<���<Wn�<Z�<��<^G�<Xܿ<m�<b��<���<��<b��<4�<�x�<��<�\�<�Ȱ<v1�<U��<���<�U�<Y��<��<\�<Z��<���<tG�<e��<�֜<��<�\�<盗<6ٕ<��<�M�<�<���<M��<h#�<6U�<υ�<M��<��<z�<}>�<]�|<�,y<��u<��q</n<q�j<��f<�/c<��_<��[<74X<�T<�P<�BM<�I<��E<!aB<(�><�+;<C�7<�4<�q0<A�,<H\)<�%<�V"<��<Dc<��<�<�<,�<n[
<g<ٳ<�i <�K�;4��;�f�;s	�;���;�{�;�K�;�+�;��;|�;d-�;UO�;u��;�ƪ;}�;у�;���;k��;�#�;�҉;c��;_�~;,�t;{j;��`;'�V;�M;��C;�:;�0;�';j�;��;B�;qE;r�:���:���:�{�:$A�:<�:�h�:�ǅ:�l:�$N:��/:�:�5�9Qή9�j9yJ�8]��6��Ӹ��X������'ڹ#���"��=�rX�CHr��+��O������B���0q��ƺ�Һ"ߺf�������"��D��a�~x�E��� ���&���,���2���8�f�>��D��~J�coP�^V�HJ\�"6b�Ph��n���s���y����JԂ��ȅ�ļ��ޱ��/���?���U���;��������  �  �p=m=ɱ=�Q=��=�=�0=� =�n =o =6W�<��<���<��<4A�<�y�<$��<���<3�<�Q�<���<+��<��<��<F�<s�<���<x��<���<��<�<�<�_�<i��<��<t��<���<=��<\
�<(�<�1�<�A�<�N�<�Y�<�a�<%g�<�i�<�h�<2e�<l^�<\T�<�F�<-6�<�!�<
�<z��<5��<!��<.��<DZ�<Z+�<V��<2��<���<VF�<q�<f��<�m�<�<���<Ln�<W�<��<XG�<Uܿ<m�<i��<���<��<g��<3�<�x�<��<�\�<�Ȱ<s1�<X��<���<�U�<Z��<��<\�<f��<���<vG�<t��<�֜<��<r\�<⛗<7ٕ<��<N�<���<ƻ�<U��<g#�<+U�<ׅ�<P��<��<��<m>�<j�|<�,y<w�u<��q<$/n<��j<��f<�/c<��_<��[<4X<�T<�P<�BM<"�I<��E<#aB<7�><�+;<@�7<�4<�q0<;�,<Y\)<��%<�V"<��<!c<��<�<�<5�<^[
<z<ڳ<~i <�K�;Z��;�f�;w	�;���;�{�;�K�;�+�;��;v�;t-�;wO�;X��;�ƪ;��;ƃ�;���;���;�#�;R҉;v��;"�~;V�t;S{j;V�`;.�V;M;�C;�:;~�0;��';��;Ҹ;�;�E;�q�:c��:O��:�{�:�A�:,<�:'h�:�ǅ:ƪl:$N:�/:D:�4�9�Ѯ9j9gH�8���6d�Ӹ&�X�����c&ڹG#���"�ם=�|X��Ir��+�� ���������q��aƺ�ҺO!ߺ̐뺯���#"�9E��a��x�q��� ���&�D�,���2�՝8�,�>��D�/J�#oP��]V��J\��5b��h��n���s�8�y����AԂ�]ȅ���������(���R�������H���g����  �  �p=u=Ǳ=�Q=��=��=�0=� =�n =k =6W�<��<���<��<9A�<�y�<��<���<2�<�Q�<���<#��<$��<��<F�<�r�<���<���<���<��<�<�<�_�<_��<��<r��<���<C��<J
�<*�<�1�<�A�<�N�<�Y�<�a�< g�<ti�<�h�<Ce�<q^�<RT�<�F�<'6�<�!�<�	�<}��<9��<#��<5��<=Z�<_+�<P��<7��<څ�<UF�<��<[��<�m�<�<���<Kn�<Q�<��<OG�<Xܿ<�l�<m��<���<��<e��<&�<�x�<��<�\�<�Ȱ<x1�<\��<���<�U�<T��<��<\�<c��<���<tG�<w��<�֜<��<u\�<<4ٕ<��<N�<���<λ�<I��<r#�<7U�<Ņ�<F��<��<��<i>�<h�|<�,y<{�u<��q</n<��j<��f<�/c<��_<��[<(4X<��T<�P<�BM<A�I<��E<aB<�><�+;<a�7<�4<�q0<.�,<Z\)<��%<�V"<��<-c<��<��<�<4�<_[
<~<̳<�i <�K�;��;~f�;w	�;��;�{�;�K�;�+�;��;N�;W-�;oO�;P��;�ƪ;@�;̓�;���;x��;�#�;N҉;���;��~;�t;�zj;�`;U�V;�M;(�C;~:;��0;Ƨ';��;��;�;�E;Dq�:���:���:�{�:FA�:%<�:_i�:>ǅ:�l:9#N:1�/:1:e3�9�Ϯ9�j9�K�8p��6�Ӹ�X� ����&ڹ�$��"��=�#X��Jr�\+���������ᾬ�wq���ƺL�Һt!ߺ�������	"�iE�ha��x����� ���&�?�,�ޡ2���8���>���D��~J��oP�<^V��J\�o5b��h��n�$�s�)�y�����Ԃ�=ȅ���������`���Z���q���d���l����  �  �p=l=Ʊ=�Q=��=��=�0=� =�n =o =2W�<��<���<��<;A�<�y�<0��<���<2�<�Q�<���<&��<��<��<F�<s�<w��<w��<���<��<�<�<�_�<d��<��<h��<���<8��<P
�<&�<�1�<�A�<�N�<�Y�<�a�<(g�<�i�<�h�<=e�<m^�<[T�<G�<06�<�!�<
�<}��<:��<#��<2��<LZ�<[+�<Z��<>��<��<TF�<|�<b��<�m�<�<���<Nn�<V�<��<TG�<Sܿ<�l�<e��<���<��<c��<,�<�x�<��<�\�<�Ȱ<q1�<K��<���<�U�<Y��<��<\�<e��<���<xG�<u��<�֜<��<x\�<<=ٕ<��<N�<���<ѻ�<N��<g#�<8U�<̅�<X��<��<z�<p>�<_�|<�,y<|�u<��q</n<z�j<��f<�/c<��_<��[<'4X< �T<�P<�BM<�I<��E<5aB<#�><�+;<D�7<�4<�q0<<�,<Q\)<��%<�V"<��<0c<��<�<�<5�<q[
<�<ҳ<�i <�K�;@��;�f�;B	�;��;�{�;�K�;�+�;��;b�;^-�;HO�;I��;�ƪ;X�;���;���;m��;�#�;c҉;J��;9�~;|�t;%{j;��`;:�V;M;\�C;�:;s�0;2�';��;��;�;�E;8r�:u��:���:`|�:�A�:<�:�h�:�ǅ:�l:r$N:��/::�4�9�ή9^	j9�E�8�G�6��Ӹ��X�o���B'ڹ$�W�"��=�X�dIr��+������������*q���ƺ8�ҺZ!ߺ�뺓���"��D��a��x����� �h�&�f�,���2��8�^�>�
�D��~J��oP��]V��J\�6b��h��n��s�$�y����pԂ�~ȅ����ձ��R���]���r���Q��������  �  �p=m=ɱ=�Q=��=��=�0=� =�n =q ==W�<��<���<��<FA�<�y�<-��<���<;�<�Q�<���<7��<��<��<F�<s�<���<x��<���<��<�<�<�_�<`��<��<n��<���<3��<Y
�<�<�1�<�A�<�N�<�Y�<�a�<%g�<|i�<�h�<:e�<r^�<eT�<�F�<66�<�!�<

�<w��<9��<&��<+��<MZ�<]+�<`��<0��<��<]F�<y�<g��<�m�<�<���<Mn�<L�<��<WG�<Dܿ<m�<^��<���<��<\��<,�<�x�<��<�\�<�Ȱ<p1�<T��<���<�U�<`��<��<"\�<d��<���<~G�<x��<�֜<��<�\�<囗<:ٕ<��<
N�<Ņ�<»�<^��<g#�<9U�<υ�<O��<��<|�<o>�<O�|<�,y<q�u<q�q</n<w�j<��f<�/c<��_<o�[<4X<	�T< �P<�BM< �I<��E<&aB<$�><�+;<>�7<�4<�q0<E�,<h\)<��%<�V"<��<Fc<��<�<�<G�<i[
<x<��<�i <L�;.��;�f�;m	�;���;�{�;�K�;�+�;��;R�;S-�;^O�;}��;�ƪ;|�;���;���;���;�#�;d҉;d��;$�~;8�t;D{j;��`;^�V;]M;��C; :;��0;C�';��;��;4�;�E;Fr�:���:���:}{�:B�:�<�:�h�:�ǅ:�l:�#N:r�/:n:I2�9�Ϯ9)j9�7�8��6ҰӸ��X�;����(ڹ�#���"���=�,X�Jr��+��`�� ���i����p��ƺB�Һe!ߺ���6����!��D��a��x�U��ɖ �U�&��,�x�2��8�ߕ>�	�D��~J�goP��]V��J\�6b��h�-	n���s�Q�y���PԂ��ȅ�ʼ��ɱ��<�����������?��������  �  �p=p=ȱ=�Q=��=��=�0=� =�n =p =<W�<��<���<��<HA�<�y�<-��<���<7�<�Q�< ��<(��<��<��<F�<s�<���<x��<���<��<�<�<�_�<b��<ݠ�<c��<���<.��<N
�<)�<�1�<�A�<�N�<�Y�<�a�<g�<~i�<�h�<?e�<j^�<\T�<�F�<06�<�!�<�	�<���<C��<.��<?��<AZ�<^+�<Z��<=��<��<SF�<~�<Y��<�m�<�<���<Hn�<S�<��<LG�<Sܿ<�l�<Z��<���<�<Z��<*�<�x�<��<�\�<�Ȱ<o1�<Z��<���<�U�<R��<��<\�<g��<���<zG�<w��<�֜<��<�\�<���<Eٕ<��<N�<���<˻�<Q��<j#�<8U�<˅�<P��<��<��<h>�<_�|<�,y<{�u<��q</n<g�j<��f<}/c<��_<��[<+4X<�T<�P<�BM<-�I<��E<%aB<!�><�+;<H�7<�4<�q0<?�,<f\)<��%<�V"<��<Kc<��<�<�<?�<r[
<�<׳<�i <�K�;8��;�f�;w	�;���;�{�;�K�;�+�;��;^�;I-�;5O�;0��;�ƪ;R�;˃�;���;l��;�#�;L҉;���;��~;C�t;�zj;Ĉ`;&�V;M;>�C;�:;��0;�';)�;H�;p�;/F;�q�:���:���:N|�:�A�:<�: i�: ǅ:0�l:�"N:�/:�:#4�9Ϯ9�j9�F�84/�6q�ӸW Y�[���S)ڹA$�E�"��=��X�EJr��+�����q���!����q���ƺ�Һ7!ߺ*��m���"� E�9a�gx�݉�v� ���&��,���2���8�J�>��D��~J��oP��]V��J\��5b��h��n�Q�s�*�y����~Ԃ��ȅ����󱋻b���X���k�������{����  �  �p=o=��=�Q=��=��=�0=� =�n =j =FW�<��<���<��</A�<�y�<+��<���<9�<�Q�<��<%��<&��<��<F�<s�<y��<y��<���<��<�<�<�_�<O��<��<o��<���<B��<D
�<&�<�1�<�A�<O�<�Y�<�a�<g�<�i�<�h�<Ee�<o^�<ZT�<G�<%6�<�!�<
�<���<7��<��<:��<EZ�<o+�<Q��<@��<߅�<UF�<��<T��<�m�<�<���<An�<a�<��<IG�<Rܿ<�l�<m��<���<��<i��<�<�x�<��<�\�<�Ȱ<o1�<O��<���<�U�<L��<��<\�<j��<���<yG�<���<�֜<��<k\�<<@ٕ<��<N�<���<ֻ�<M��<t#�<7U�<˅�<Y��<��<��<a>�<y�|<�,y<v�u<r�q</n<��j<��f<�/c<��_<e�[<'4X<ߌT<'�P<�BM<*�I<u�E<3aB<(�><�+;<a�7<�4<�q0<)�,<{\)<��%<�V"<��<c<��<�<<D�<f[
<�<ѳ<�i <�K�;\��;�f�;J	�;���;�{�;�K�;�+�;��;�;r-�;fO�;E��;�ƪ;)�;���;���;]��;%$�;.҉;z��;��~;��t;�zj;��`;L�V;M;q�C;w:;1�0;�';�;�;��;F;�q�:���:��:x|�:�A�:)<�:�i�:�ƅ:-�l:"N:�/::|7�9�ή9)j95F�8H�6[�Ӹ��X�ʏ���%ڹ�&���"�!�=��X��Ir��+���������V����q���ƺ1�Һ!ߺM�뺀����!�E�ta�*y����� �d�&���,��2�O�8�j�>���D��~J��oP��]V�K\��5b�0 h��n�t�s�<�y����Ԃ�Yȅ�
�������]�������r�������U����  �  �p=q=ʱ=�Q=��=��=�0=� =�n =n =>W�<��<���<�<NA�<�y�</��<���<9�<�Q�<��<2��<��<��<F�<s�<���<}��<���<��<�<�<�_�<U��<۠�<^��<���<*��<Q
�<�<�1�<�A�<�N�<�Y�<�a�<#g�<�i�<�h�<;e�<u^�<dT�<G�</6�<�!�<
�<���<L��<7��<<��<IZ�<^+�<Y��<;��<��<[F�<~�<U��<�m�<�<���<En�<P�<���<VG�<Kܿ<�l�<W��<��<y�<Y��<"�<�x�<��<�\�<�Ȱ<r1�<\��<���<�U�<O��<��<\�<o��<���<xG�<v��<�֜<��<�\�<���<Bٕ<��<N�<���<Ի�<Y��<r#�<3U�<Ņ�<Q��<��<��<f>�<Y�|<�,y<��u<k�q</n<c�j<��f<z/c<��_<g�[</4X<�T<�P<�BM<2�I<��E<'aB<�><�+;<Y�7<�4<�q0<8�,<i\)<��%<�V"<��<Wc<��<�<�<C�<g[
<�<�<�i <�K�;��;�f�;�	�;��;�{�;�K�;�+�;��;*�;C-�; O�;+��;vƪ;^�;���;���;>��;�#�;?҉;���;�~;h�t;�zj;��`;x�V;VM;P�C;�:;��0;�';��;��;��;F;r�:���:���:-|�:7B�:�<�:	i�:�ƅ:��l:�#N:�/:k:s3�9rˮ9�
j9K?�8�)�69�Ӹ)Y���)ڹH%�r�"���=�cX��Jr��+�����H���m����q��Pƺ��Һ� ߺ��뺇���"��D�=a�:x������ ���&��,���2�i�8��>���D��~J��oP��]V�|J\��5b� h�	n�`�s���y�*��iԂ��ȅ��������T�������c���x��������  �  �p=g=Ʊ=�Q=��=��=�0=� =�n =u =;W�<��<���<��<6A�<�y�<=��<���<A�<�Q�<��<)��<��<��<F�<s�<|��<j��<���<��<�<�<�_�<b��<۠�<k��<���<#��<_
�<�<�1�<�A�<�N�<�Y�<�a�<g�<{i�<�h�<Ae�<p^�<]T�<�F�<A6�<�!�<
�<���<2��<��<5��<VZ�<Y+�<k��<9��<��<VF�<�<n��<�m�<�<���<Dn�<X�<���<TG�<9ܿ<m�<Q��<���<��<X��<0�<�x�<��<�\�<�Ȱ<c1�<N��<���<�U�<g��<��<\�<j��<���<�G�<t��<�֜<��<r\�<㛗<Kٕ<��<N�<υ�<ǻ�<R��<j#�<@U�<օ�<J��<��<v�<n>�<\�|<�,y<x�u<f�q</n<X�j<�f<w/c<��_<l�[<4X<�T<�P<�BM<�I<��E<aB<0�><�+;<D�7<�4<�q0<V�,<e\)<��%<W"<��<'c<��<4�<�<S�<y[
<�<ٳ<�i <0L�;8��;�f�;W	�;º�;�{�;�K�;�+�;��;[�;D-�;TO�;���;\ƪ;��;d��;���;L��;�#�;P҉;Q��;��~;0�t;�{j;׈`;O�V;M;�C;V:;z�0;��';��;Ÿ;��;�E;�r�:`��:���:|�:�A�:B<�: i�:vȅ:��l:�"N:��/:O:�5�9�̮9�	j9*-�8�6b�Ӹ��X�����)ڹ�#���"�Ӟ=�YX�FIr��,�����h���G���>p���ƺ�Һ!ߺ!�뺣���"�yD��a��x�d��A� �N�&�.�,�*�2�̝8�C�>��D��~J�+oP�^V��J\�=6b��h��n�`�s�5�y�@��JԂ��ȅ���������D�����������x��������  �  �p=q=ʱ=�Q=��=��=�0=� =�n =n =>W�<��<���<�<NA�<�y�</��<���<9�<�Q�<��<2��<��<��<F�<s�<���<}��<���<��<�<�<�_�<U��<۠�<^��<���<*��<Q
�<�<�1�<�A�<�N�<�Y�<�a�<#g�<�i�<�h�<;e�<u^�<dT�<G�</6�<�!�<
�<���<L��<7��<<��<IZ�<^+�<Y��<;��<��<[F�<~�<U��<�m�<�<���<En�<P�<���<VG�<Kܿ<�l�<W��<��<y�<Y��<"�<�x�<��<�\�<�Ȱ<r1�<\��<���<�U�<O��<��<\�<o��<���<xG�<v��<�֜<��<�\�<���<Bٕ<��<N�<���<Ի�<Y��<r#�<3U�<Ņ�<Q��<��<��<f>�<Y�|<�,y<��u<k�q</n<c�j<��f<z/c<��_<g�[</4X<�T<�P<�BM<2�I<��E<'aB<�><�+;<Y�7<�4<�q0<8�,<i\)<��%<�V"<��<Wc<��<�<�<C�<g[
<�<�<�i <�K�;��;�f�;�	�;��;�{�;�K�;�+�;��;*�;C-�; O�;+��;vƪ;^�;���;���;>��;�#�;?҉;���;�~;h�t;�zj;��`;x�V;VM;P�C;�:;��0;�';��;��;��;F;r�:���:���:-|�:7B�:�<�:	i�:�ƅ:��l:�#N:�/:k:s3�9rˮ9�
j9K?�8�)�69�Ӹ)Y���)ڹH%�r�"���=�cX��Jr��+�����H���m����q��Pƺ��Һ� ߺ��뺇���"��D�=a�:x������ ���&��,���2�i�8��>���D��~J��oP��]V�|J\��5b� h�	n�`�s���y�*��iԂ��ȅ��������T�������c���x��������  �  �p=o=��=�Q=��=��=�0=� =�n =j =FW�<��<���<��</A�<�y�<+��<���<9�<�Q�<��<%��<&��<��<F�<s�<y��<y��<���<��<�<�<�_�<O��<��<o��<���<B��<D
�<&�<�1�<�A�<O�<�Y�<�a�<g�<�i�<�h�<Ee�<o^�<ZT�<G�<%6�<�!�<
�<���<7��<��<:��<EZ�<o+�<Q��<@��<߅�<UF�<��<T��<�m�<�<���<An�<a�<��<IG�<Rܿ<�l�<m��<���<��<i��<�<�x�<��<�\�<�Ȱ<o1�<O��<���<�U�<L��<��<\�<j��<���<yG�<���<�֜<��<k\�<<@ٕ<��<N�<���<ֻ�<M��<t#�<7U�<˅�<Y��<��<��<a>�<y�|<�,y<v�u<r�q</n<��j<��f<�/c<��_<e�[<'4X<ߌT<'�P<�BM<*�I<u�E<3aB<(�><�+;<a�7<�4<�q0<)�,<{\)<��%<�V"<��<c<��<�<<D�<f[
<�<ѳ<�i <�K�;\��;�f�;J	�;���;�{�;�K�;�+�;��;�;r-�;fO�;E��;�ƪ;)�;���;���;]��;%$�;.҉;z��;��~;��t;�zj;��`;L�V;M;q�C;w:;1�0;�';�;�;��;F;�q�:���:��:x|�:�A�:)<�:�i�:�ƅ:-�l:"N:�/::|7�9�ή9)j95F�8H�6[�Ӹ��X�ʏ���%ڹ�&���"�!�=��X��Ir��+���������V����q���ƺ1�Һ!ߺM�뺀����!�E�ta�*y����� �d�&���,��2�O�8�j�>���D��~J��oP��]V�K\��5b�0 h��n�t�s�<�y����Ԃ�Yȅ�
�������]�������r�������U����  �  �p=p=ȱ=�Q=��=��=�0=� =�n =p =<W�<��<���<��<HA�<�y�<-��<���<7�<�Q�< ��<(��<��<��<F�<s�<���<x��<���<��<�<�<�_�<b��<ݠ�<c��<���<.��<N
�<)�<�1�<�A�<�N�<�Y�<�a�<g�<~i�<�h�<?e�<j^�<\T�<�F�<06�<�!�<�	�<���<C��<.��<?��<AZ�<^+�<Z��<=��<��<SF�<~�<Y��<�m�<�<���<Hn�<S�<��<LG�<Sܿ<�l�<Z��<���<�<Z��<*�<�x�<��<�\�<�Ȱ<o1�<Z��<���<�U�<R��<��<\�<g��<���<zG�<w��<�֜<��<�\�<���<Eٕ<��<N�<���<˻�<Q��<j#�<8U�<˅�<P��<��<��<h>�<_�|<�,y<{�u<��q</n<g�j<��f<}/c<��_<��[<+4X<�T<�P<�BM<-�I<��E<%aB<!�><�+;<H�7<�4<�q0<?�,<f\)<��%<�V"<��<Kc<��<�<�<?�<r[
<�<׳<�i <�K�;8��;�f�;w	�;���;�{�;�K�;�+�;��;^�;I-�;5O�;0��;�ƪ;R�;˃�;���;l��;�#�;L҉;���;��~;C�t;�zj;Ĉ`;&�V;M;>�C;�:;��0;�';)�;H�;p�;/F;�q�:���:���:N|�:�A�:<�: i�: ǅ:0�l:�"N:�/:�:#4�9Ϯ9�j9�F�84/�6q�ӸW Y�[���S)ڹA$�E�"��=��X�EJr��+�����q���!����q���ƺ�Һ7!ߺ*��m���"� E�9a�gx�݉�v� ���&��,���2���8�J�>��D��~J��oP��]V��J\��5b��h��n�Q�s�*�y����~Ԃ��ȅ����󱋻b���X���k�������{����  �  �p=m=ɱ=�Q=��=��=�0=� =�n =q ==W�<��<���<��<FA�<�y�<-��<���<;�<�Q�<���<7��<��<��<F�<s�<���<x��<���<��<�<�<�_�<`��<��<n��<���<3��<Y
�<�<�1�<�A�<�N�<�Y�<�a�<%g�<|i�<�h�<:e�<r^�<eT�<�F�<66�<�!�<

�<w��<9��<&��<+��<MZ�<]+�<`��<0��<��<]F�<y�<g��<�m�<�<���<Mn�<L�<��<WG�<Dܿ<m�<^��<���<��<\��<,�<�x�<��<�\�<�Ȱ<p1�<T��<���<�U�<`��<��<"\�<d��<���<~G�<x��<�֜<��<�\�<囗<:ٕ<��<
N�<Ņ�<»�<^��<g#�<9U�<υ�<O��<��<|�<o>�<O�|<�,y<q�u<q�q</n<w�j<��f<�/c<��_<o�[<4X<	�T< �P<�BM< �I<��E<&aB<$�><�+;<>�7<�4<�q0<E�,<h\)<��%<�V"<��<Fc<��<�<�<G�<i[
<x<��<�i <L�;.��;�f�;m	�;���;�{�;�K�;�+�;��;R�;S-�;^O�;}��;�ƪ;|�;���;���;���;�#�;d҉;d��;$�~;8�t;D{j;��`;^�V;]M;��C; :;��0;C�';��;��;4�;�E;Fr�:���:���:}{�:B�:�<�:�h�:�ǅ:�l:�#N:r�/:n:I2�9�Ϯ9)j9�7�8��6ҰӸ��X�;����(ڹ�#���"���=�,X�Jr��+��`�� ���i����p��ƺB�Һe!ߺ���6����!��D��a��x�U��ɖ �U�&��,�x�2��8�ߕ>�	�D��~J�goP��]V��J\�6b��h�-	n���s�Q�y���PԂ��ȅ�ʼ��ɱ��<�����������?��������  �  �p=l=Ʊ=�Q=��=��=�0=� =�n =o =2W�<��<���<��<;A�<�y�<0��<���<2�<�Q�<���<&��<��<��<F�<s�<w��<w��<���<��<�<�<�_�<d��<��<h��<���<8��<P
�<&�<�1�<�A�<�N�<�Y�<�a�<(g�<�i�<�h�<=e�<m^�<[T�<G�<06�<�!�<
�<}��<:��<#��<2��<LZ�<[+�<Z��<>��<��<TF�<|�<b��<�m�<�<���<Nn�<V�<��<TG�<Sܿ<�l�<e��<���<��<c��<,�<�x�<��<�\�<�Ȱ<q1�<K��<���<�U�<Y��<��<\�<e��<���<xG�<u��<�֜<��<x\�<<=ٕ<��<N�<���<ѻ�<N��<g#�<8U�<̅�<X��<��<z�<p>�<_�|<�,y<|�u<��q</n<z�j<��f<�/c<��_<��[<'4X< �T<�P<�BM<�I<��E<5aB<#�><�+;<D�7<�4<�q0<<�,<Q\)<��%<�V"<��<0c<��<�<�<5�<q[
<�<ҳ<�i <�K�;@��;�f�;B	�;��;�{�;�K�;�+�;��;b�;^-�;HO�;I��;�ƪ;X�;���;���;m��;�#�;c҉;J��;9�~;|�t;%{j;��`;:�V;M;\�C;�:;s�0;2�';��;��;�;�E;8r�:u��:���:`|�:�A�:<�:�h�:�ǅ:�l:r$N:��/::�4�9�ή9^	j9�E�8�G�6��Ӹ��X�o���B'ڹ$�W�"��=�X�dIr��+������������*q���ƺ8�ҺZ!ߺ�뺓���"��D��a��x����� �h�&�f�,���2��8�^�>�
�D��~J��oP��]V��J\�6b��h��n��s�$�y����pԂ�~ȅ����ձ��R���]���r���Q��������  �  �p=u=Ǳ=�Q=��=��=�0=� =�n =k =6W�<��<���<��<9A�<�y�<��<���<2�<�Q�<���<#��<$��<��<F�<�r�<���<���<���<��<�<�<�_�<_��<��<r��<���<C��<J
�<*�<�1�<�A�<�N�<�Y�<�a�< g�<ti�<�h�<Ce�<q^�<RT�<�F�<'6�<�!�<�	�<}��<9��<#��<5��<=Z�<_+�<P��<7��<څ�<UF�<��<[��<�m�<�<���<Kn�<Q�<��<OG�<Xܿ<�l�<m��<���<��<e��<&�<�x�<��<�\�<�Ȱ<x1�<\��<���<�U�<T��<��<\�<c��<���<tG�<w��<�֜<��<u\�<<4ٕ<��<N�<���<λ�<I��<r#�<7U�<Ņ�<F��<��<��<i>�<h�|<�,y<{�u<��q</n<��j<��f<�/c<��_<��[<(4X<��T<�P<�BM<A�I<��E<aB<�><�+;<a�7<�4<�q0<.�,<Z\)<��%<�V"<��<-c<��<��<�<4�<_[
<~<̳<�i <�K�;��;~f�;w	�;��;�{�;�K�;�+�;��;N�;W-�;oO�;P��;�ƪ;@�;̓�;���;x��;�#�;N҉;���;��~;�t;�zj;�`;U�V;�M;(�C;~:;��0;Ƨ';��;��;�;�E;Dq�:���:���:�{�:FA�:%<�:_i�:>ǅ:�l:9#N:1�/:1:e3�9�Ϯ9�j9�K�8p��6�Ӹ�X� ����&ڹ�$��"��=�#X��Jr�\+���������ᾬ�wq���ƺL�Һt!ߺ�������	"�iE�ha��x����� ���&�?�,�ޡ2���8���>���D��~J��oP�<^V��J\�o5b��h��n�$�s�)�y�����Ԃ�=ȅ���������`���Z���q���d���l����  �  �p=m=ɱ=�Q=��=�=�0=� =�n =o =6W�<��<���<��<4A�<�y�<$��<���<3�<�Q�<���<+��<��<��<F�<s�<���<x��<���<��<�<�<�_�<i��<��<t��<���<=��<\
�<(�<�1�<�A�<�N�<�Y�<�a�<%g�<�i�<�h�<2e�<l^�<\T�<�F�<-6�<�!�<
�<z��<5��<!��<.��<DZ�<Z+�<V��<2��<���<VF�<q�<f��<�m�<�<���<Ln�<W�<��<XG�<Uܿ<m�<i��<���<��<g��<3�<�x�<��<�\�<�Ȱ<s1�<X��<���<�U�<Z��<��<\�<f��<���<vG�<t��<�֜<��<r\�<⛗<7ٕ<��<N�<���<ƻ�<U��<g#�<+U�<ׅ�<P��<��<��<m>�<j�|<�,y<w�u<��q<$/n<��j<��f<�/c<��_<��[<4X<�T<�P<�BM<"�I<��E<#aB<7�><�+;<@�7<�4<�q0<;�,<Y\)<��%<�V"<��<!c<��<�<�<5�<^[
<z<ڳ<~i <�K�;Z��;�f�;w	�;���;�{�;�K�;�+�;��;v�;t-�;wO�;X��;�ƪ;��;ƃ�;���;���;�#�;R҉;v��;"�~;V�t;S{j;V�`;.�V;M;�C;�:;~�0;��';��;Ҹ;�;�E;�q�:c��:O��:�{�:�A�:,<�:'h�:�ǅ:ƪl:$N:�/:D:�4�9�Ѯ9j9gH�8���6d�Ӹ&�X�����c&ڹG#���"�ם=�|X��Ir��+�� ���������q��aƺ�ҺO!ߺ̐뺯���#"�9E��a��x�q��� ���&�D�,���2�՝8�,�>��D�/J�#oP��]V��J\��5b��h��n���s�8�y����AԂ�]ȅ���������(���R�������H���g����  �  �p=k=̱=�Q=��=��=�0=� =�n =p =-W�<ߒ�<���<��<EA�<�y�<,��<���<.�<�Q�<��<*��<��<��<F�<s�<���<y��<���<��<�<�<�_�<k��<��<l��<���<4��<Z
�<+�<�1�<�A�<�N�<�Y�<�a�<-g�<|i�<�h�<9e�<k^�<VT�<�F�<26�<�!�<
�<s��<9��<)��<(��<JZ�<L+�<[��<4��<؅�<UF�<x�<a��<�m�<�<���<Wn�<Z�<��<^G�<Xܿ<m�<b��<���<��<b��<4�<�x�<��<�\�<�Ȱ<v1�<U��<���<�U�<Y��<��<\�<Z��<���<tG�<e��<�֜<��<�\�<盗<6ٕ<��<�M�<�<���<M��<h#�<6U�<υ�<M��<��<z�<}>�<]�|<�,y<��u<��q</n<q�j<��f<�/c<��_<��[<74X<�T<�P<�BM<�I<��E<!aB<(�><�+;<C�7<�4<�q0<A�,<H\)<�%<�V"<��<Dc<��<�<�<,�<n[
<g<ٳ<�i <�K�;4��;�f�;s	�;���;�{�;�K�;�+�;��;|�;d-�;UO�;u��;�ƪ;}�;у�;���;k��;�#�;�҉;c��;_�~;,�t;{j;��`;'�V;�M;��C;�:;�0;�';j�;��;B�;qE;r�:���:���:�{�:$A�:<�:�h�:�ǅ:�l:�$N:��/:�:�5�9Qή9�j9yJ�8]��6��Ӹ��X������'ڹ#���"��=�rX�CHr��+��O������B���0q��ƺ�Һ"ߺf�������"��D��a�~x�E��� ���&���,���2���8�f�>��D��~J�coP�^V�HJ\�"6b�Ph��n���s���y����JԂ��ȅ�ļ��ޱ��/���?���U���;��������  �  �p=n=ɱ=�Q=��=��=�0=� =�n =g =8W�<��<���<��<1A�<�y�<!��<���<1�<�Q�<���<"��<��<��<F�<s�<���<y��<���<��<�<�<�_�<_��<��<z��<���<K��<Q
�<+�<�1�<�A�<�N�<�Y�<�a�<g�<i�<�h�<Ce�<i^�<WT�<�F�< 6�<�!�< 
�<r��<-��<��<%��<BZ�<Z+�<N��<4��<ޅ�<PF�<��<Z��<�m�<�<���<Mn�<Y�<��<YG�<Xܿ<�l�<v��<���<��<t��<)�<�x�<��<�\�<�Ȱ<q1�<Z��<���<�U�<P��<��<\�<a��<���<rG�<v��<�֜<��<l\�<ݛ�<2ٕ<��<N�<���<˻�<G��<i#�<7U�<˅�<N��<��<�<n>�<l�|<�,y<��u<��q<"/n<��j<��f<�/c<��_<��[<24X<�T<�P<�BM<&�I<��E< aB<&�><�+;<L�7<�4<�q0<�,<^\)<��%<�V"<��<c<|�<��<�<0�<U[
<u<ɳ<�i <�K�;3��;�f�;r	�;���;�{�;�K�;�+�;��;L�;�-�;�O�;���;�ƪ;[�;΃�;���;���;�#�;]҉;x��;��~;G�t;�zj;ۈ`;�V;�M;�C;K:;~�0;�';]�;��;��;ZE;�q�:`��:���:�{�:�A�:�;�:Xi�:%ǅ:(�l:�"N:B�/:Q:=5�9�Ѯ9nj91J�8�-�6L�Ӹ��X�����7#ڹ}$���"�؝=�X��Ir��+�������=����q��$ƺV�Һ�!ߺ������"�KE�#b�#y����� ���&�8�,�(�2���8���>���D��~J��oP��]V��J\��5b��h��n���s��y����DԂ�;ȅ������������`���]���B���j����  �  �p=u=Ǳ=�Q=��=|�=�0=
� =�n =e =8W�<֒�<���<��<5A�<�y�<��<���</�<�Q�<��<��<��<��<!F�<s�<���<���<���<��<�<�<`�<g��<��<t��<���<C��<S
�<;�<�1�<�A�<�N�<�Y�<�a�<g�<�i�<�h�<8e�<i^�<_T�<�F�<6�<�!�<�	�<���<6��<!��<7��<2Z�<Z+�<K��<4��<��<LF�<{�<T��<�m�<	�<���<Mn�<X�<��<SG�<iܿ<�l�<q��<���<��<o��</�<y�<��<�\�<�Ȱ<x1�<^��<���<�U�<G��<��<
\�<q��<���<oG�<r��<�֜<��<r\�<뛗<:ٕ<��<	N�<���<ϻ�<H��<j#�<+U�<υ�<V��<��<��<k>�<x�|<�,y<��u<��q</n<��j<��f<�/c<��_<��[<B4X<�T<,�P<�BM<A�I<��E<*aB<1�><�+;<J�7<�4<�q0<�,<]\)<m�%<�V"<��<#c<��<�<�<,�<K[
<�<��<�i <�K�;c��;�f�;u	�;��;�{�;L�;�+�;7�;m�;�-�;rO�;,��;�ƪ;`�;��;���;���;�#�;S҉;���;��~;��t;�zj;��`;�V;,M;�C;=:;��0;Z�';٠;۸;�;�E;�p�:g��:���:�{�:GB�:�;�:�h�:�ƅ:'�l:W"N:��/:R:�4�9
Ү9Yj9H[�8
`�6��Ӹ`�X�َ���$ڹ�#���"�,�=�!X��Ir�l+���������F���Er���ƺڢҺ� ߺ1��#���3"��E�za��x�*��ϖ �.�&�%�,�:�2���8���>��D�6J�coP��]V��J\�h5b��h��n��s���y�H��QԂ�Mȅ�$�������,���,���=���m���J����  �  �p=r=Ǳ=�Q=��=��=�0=� =�n =i =9W�<ْ�<���<��<4A�<�y�<%��<���<8�<�Q�<���< ��<��<��<F�<�r�<~��<���<���<��<�<�<�_�<c��<��<���<���<I��<Z
�<*�<�1�<�A�<O�<�Y�<�a�<g�<}i�<�h�<De�<k^�<UT�<�F�<,6�<�!�<�	�<p��<&��<��<#��<AZ�<U+�<Y��<%��<ۅ�<OF�<��<`��<�m�<�<���<Un�<_�<��<XG�<Xܿ<m�<t��<���<��<n��</�<�x�<��<�\�<�Ȱ<|1�<T��<���<�U�<X��<��<\�<a��<���<{G�<i��<�֜<��<n\�<ٛ�<1ٕ<��<N�<���<���<F��<n#�<<U�<΅�<G��<��<��<x>�<{�|<�,y<��u<��q<"/n<��j<
�f<�/c<��_<��[<64X< �T<,�P<�BM<8�I<��E<aB<)�><�+;<R�7<�4<�q0<&�,<_\)<s�%<�V"<��< c<w�<�<�<>�<K[
<r<ĳ<�i <�K�;<��;zf�;Z	�;��;�{�;�K�;�+�;��;\�;�-�;�O�;���;�ƪ;|�;˃�;���;|��;$�;x҉;���;��~;5�t;{j;�`;&�V;�M;��C;�:;k�0;Ƨ';N�;^�;��;HE;~q�:��:u��:�z�:TA�:�;�:Yi�:�ǅ:��l:�"N:~�/:I:�6�9�Ю9�
j9QJ�8��6��Ӹ�X�[����$ڹ�#���"��=��X��Hr�*+��t������뽬�;q��Gƺ��Һ�!ߺ���o���w"�3E�;b�y����� ��&�6�,��2��8���>�ԋD��~J�ioP�6^V��J\��5b�uh�{n�
�s���y����EԂ�+ȅ�����}���&���K���U���Q���M����  �  �o=�=��=�O={�=�=.=�� =wk =�	 ='O�<I��<���<��<�6�<�n�<u��<7��<�<�C�<yv�<��<
��<��<z4�<�`�<`��<y��<��<��<%&�<wH�< i�<���<!��<���<���<7��<� �<��<]!�<�-�<�7�<�>�<C�<MD�<�B�<	>�<G6�<L+�<��<E�<��<`��<���<���<)}�<nU�<�)�<L��<���<+��<kS�<w�<I��<���<C:�<o��<"��<�:�<���<�z�<E�<w��<�:�<eǼ<!P�<�Թ<9U�<�Ѷ<NJ�<��<�/�<��<��<�l�<ϫ< .�<≨<~�<8�<���<kڡ<a'�<�q�<���<���<�A�<���<���<G��<9�<Rr�<ҩ�<�ߌ<S�<�G�<�y�<���<�ڃ<�	�<=8�<��|<,&y<�u<��q<:1n<`�j<��f<R:c<u�_<�[<�GX<w�T<J Q<+_M<<�I<�!F<�B<��><nV;<��7<m24<�0<c-<O�)<k&<��"<<��<p7<��<g<<�
<�X<b
<e� <E�;���;&�;��;y��;JG�;o�;Q��;D��;���;;�;m,�;�a�;���;5��;kg�;��;�l�;�	�;n��;�w�;�I�;�Xv;Al;�Kb;<yX;��N;I9E;M�;;H}2;�P);VC ;�U;4�;9�;���:U��:&��:�\�:��:���:��:�e�::�q:�S:t�4:��:(Y�9���9�I{9�K9�M�7�o��?�I�
C���ӹt��
��&r:��U�ZYo���6���ɩ������?��P�ĺщѺ,޺"������x����#����,�H= �1J&�FS,�W2��W8��T>�qOD��FJ��;P�:.V��\��b���g�,�m� �s���y����̂�Å�#���G�����������������������  �  �o=�=��=�O=��=�=.=�� =uk =�	 =;O�<H��<���<��<�6�<�n�<l��<A��<!�<�C�<rv�<��<��< �<�4�<�`�<Q��<k��<��<��<&�<qH�<�h�<���<.��<���<��<.��<� �<n�<e!�<�-�<�7�<�>�<�B�<RD�<�B�<>�<Q6�<F+�<��<D�<��<X��<���<��<}�<vU�<�)�<]��<���<*��<eS�<}�<^��<���<M:�<Y��<��<�:�<���<�z�</�<y��<�:�<nǼ</P�<�Թ<<U�<�Ѷ<JJ�<���<�/�<��<z�<tl�<�Ϋ<.�<艨<��<8�<���<mڡ<o'�<�q�<���<���<�A�<���<���<B��<.9�<Qr�<Ω�<�ߌ<a�<�G�<�y�<���<�ڃ<�	�<!8�<��|<,&y<�u<��q<,1n<w�j<��f<f:c<j�_<�[<�GX<l�T<j Q<�^M<5�I<�!F<�B<	�><�V;<��7<V24<�0<e-<w�)<g&<��"<&<h�<�7<��<,g<?<�
<�X<U
<�� <l�;I��;�%�;���;@��;�F�;��;��;*��;���;;�;�,�;�a�;���;��;vg�;u�;�l�;�	�;���;�w�;mI�;�Xv;kAl;lLb;�yX;v�N;89E;H�;;�}2;�P);uC ;U;��;v�;��:o��:k��:r\�:"�:\��:��:(f�:��q: S:S�4:��:FW�9v��9�>{99M9�)�7�f���I�.?���ӹ?��q��bt:�� U��[o��Ä� ������~��J?���ĺ�Ѻ�޺������	��R������,�[= �YJ&��R,�$W2��W8�U>�OD�oFJ�J;P�j.V�P\��b���g���m� �s�	�y�׭��̂�����������������Ø������Ӎ���  �  �o=�=��=�O=��=ߎ=.=�� ={k =�	 =;O�<C��<���<(��<�6�<�n�<`��<E��<�<�C�<yv�<٧�<��<��<�4�<�`�<a��<���<���<��<&�<zH�<�h�<���<&��<���<��<'��<
�<g�<r!�<�-�<�7�<�>�<�B�<YD�<�B�<
>�<B6�<A+�<��<8�<��<N��<	��<���<}�<�U�<�)�<b��<���<,��<bS�<o�<N��<��<W:�<W��<7��<�:�<���<�z�<(�<���<�:�<tǼ<P�<�Թ<=U�<�Ѷ<WJ�<���<�/�<���<��<�l�<�Ϋ<.�<҉�<��<8�<���<jڡ<d'�<�q�<w��<���<�A�<Ƃ�<���<:��<29�<Er�<ک�<�ߌ<Z�<�G�<�y�<���<�ڃ<�	�<8�<��|<1&y<�u<��q<$1n<��j<��f<h:c<f�_<-�[<�GX<f�T<� Q<�^M<l�I<�!F<�B<�><]V;<��7<I24<+�0<R-<w�)<^&<��"<I<i�<�7<��<4g<1<ڬ
<�X<A
<}� <�;_��;�%�;��;���;�F�;�;���;P��;���;9�;�,�;�a�;ߧ�;���;�g�;Y�;m�;�	�;��;gx�;gI�;�Xv;�@l;�Kb;yX;P�N;f9E;��;;~2;oP);�C ;rU;�;��;<��:Ē�:���:�\�:��:|��:��:�d�:��q:�S:�4:��:�W�9\��96;{9�V9-�7�`����I��B���ӹ������u:���T�.\o����������;~���@����ĺ��Ѻ`޺<�꺨��������9����+�W= ��J&��R,�W2��W8�AU>�;OD�GJ�y;P�T.V�?\��b��g�o�m��s�"�y�~���̂���w���������������������������  �  �o=�=��=�O=��=�=.=�� ={k =�	 =6O�<N��<���<��<�6�<�n�<f��<L��<�<�C�<zv�<��<$��<��<�4�<�`�<R��<v��<��<��<&�<{H�<�h�<���</��<���<��<#��<� �<m�<e!�<�-�<�7�<�>�<�B�<VD�<�B�<>�<Q6�<F+�<��<A�<��<\��<���<��<}�<sU�<�)�<c��<���<0��<fS�<|�<^��<��<R:�<Y��<��<�:�<���<�z�<.�<���<�:�<zǼ<"P�<�Թ<CU�<�Ѷ<TJ�<���<�/�<��<��<wl�<�Ϋ<.�<䉨<��<8�<���<pڡ<c'�<�q�<���<���<�A�<���<y��<F��<-9�<Or�<ܩ�<�ߌ<g�<�G�<�y�<���<�ڃ<�	�<%8�<��|<+&y<�u<��q<!1n<��j<��f<v:c<g�_<�[<�GX<e�T<k Q<�^M<D�I<�!F<�B<��><�V;<��7<V24<,�0<_-<m�)<t&<��"<0<q�<�7<��<Bg<(<�
<�X<U
<�� <[�;A��;�%�;���;n��;�F�;��;��;T��;q��;O�;�,�;�a�;���;���;�g�;q�;�l�;�	�;��;x�;iI�;�Xv;7Al;mLb;�yX;t�N;{9E;2�;;~2;�P);RC ;JU;Ӆ;d�;��:Ӓ�:��:�\�:5�:N��: �:�e�:�q:)S:2�4:��:W�9̭�9;>{9�Q9���7(Z��t�I��@��;ӹ���4���t:�� U�v[o�$Ä����������~���?����ĺ�Ѻ<޺ݐ��������������	��+��= �4J&��R,�2W2�~W8�U>��ND�pFJ�p;P�I.V�^\��b���g���m� �s���y����̂���\�����������՟����������э���  �  �o=�=��=�O=}�=�=	.=�� =uk =�	 =1O�<I��<���<��<�6�<�n�<n��<A��<�<�C�<qv�<��<��<��<4�<�`�<W��<s��<��<��<&�<sH�<�h�<���<&��<���<��<*��<� �<n�<b!�<�-�<�7�<�>�<�B�<JD�<�B�<>�<J6�<F+�<��<H�<
��<_��<���<���<)}�<tU�<�)�<T��<���<*��<dS�<x�<O��<��<C:�<j��<��<�:�<���<�z�</�<}��<�:�<kǼ<P�<�Թ<:U�<�Ѷ<LJ�<���<�/�<��<��<xl�<�Ϋ<.�<䉨<��<8�<���<rڡ<h'�<�q�<���<���<�A�<�<}��<D��<$9�<Yr�<ͩ�<�ߌ<W�<�G�<�y�<���<�ڃ<�	�<28�<��|<%&y<�u<��q<(1n<r�j<��f<[:c<k�_<�[<�GX<e�T<c Q<_M<>�I<�!F<�B<��><�V;<��7<W24<�0<t-<c�)<i&<��"<8<��<�7<��<+g</<�
<�X<X
<p� <\�;��;&�;���;a��;%G�;��;��;2��;���;7�;�,�;�a�;���;��;�g�;t�;�l�;�	�;B��;�w�;�I�;vXv;"Al;Lb;[yX;v�N;'9E;g�;;�}2;�P);\C ;�U;6�;h�;]��:���:k��:p\�:�:
��:	�:�e�:M�q:JS:��4:��:>X�9]��9�>{9O9��7'i���I��A��sӹ���8���t:��U�]Zo�:Ä������������?����ĺ��Ѻ�޺���p�����=��������+�u= �CJ&��R,��V2��W8�U>�SOD��FJ��;P�.V��\��b�J�g���m�9�s��y����̂���Y���6���������Ę������ፚ��  �  �o=�=��=�O=��=�=	.=�� =xk =�	 =8O�<O��<���<$��<�6�<�n�<l��<I��<�<�C�<zv�<��<��<��<�4�<�`�<T��<z��<���<��<&�<qH�<�h�<���<*��<���<��<$��<� �<f�<l!�<�-�<�7�<�>�<�B�<KD�<�B�<>�<O6�<W+�<��<?�<��<\��<��<��<}�<xU�<�)�<d��<���<*��<sS�<��<O��<���<F:�<V��<��<�:�<���<�z�<'�<z��<�:�<mǼ<%P�<�Թ<6U�<�Ѷ<JJ�<���<�/�<���<��<vl�<�Ϋ<.�<牨<��<&8�<���<kڡ<h'�<�q�<���<���<�A�<Ă�<���<G��<-9�<Lr�<Щ�<�ߌ<W�<�G�<�y�<���<�ڃ<�	�< 8�<��|<2&y<�u<��q<1n<v�j<��f<a:c<[�_<"�[<�GX<o�T<i Q<�^M<N�I<�!F<��B<
�><|V;<��7<~24<�0<[-<q�)<u&<��"<B<g�<�7<��<;g<4<�
<�X<t
<p� <]�;?��;�%�;���;���;�F�;��;��;.��;���;�;�,�;�a�;���;���;�g�;V�;�l�;�	�;��;x�;gI�;�Xv;�Al;�Kb;~yX;��N;39E;!�;;~2;�P);�C ;dU;��;��;'��:ڒ�:���:n\�:�:���:
�:Yf�:��q:�S:�4:��:$V�9Ϯ�9R;{9�M9��7�g����I��@��Iӹ���j���t:�� U�]\o�Ä�����6�����a?����ĺ%�Ѻ޺+��u������W�������+�== �-J&��R,�CW2��W8�{T>�VOD��FJ�:;P��.V�L\��b���g���m��s�G�y�����̂���H���*�����������Ԙ������Ս���  �  �o=�=��=�O=��=�=.=�� =xk =�	 =BO�<S��<���<*��<�6�<�n�<b��<S��<�<�C�<wv�<��<��<��<�4�<�`�<T��<|��< ��<��<&�<}H�<�h�<���<*��<���<	��<��<�<g�<c!�<�-�<�7�<�>�<�B�<ZD�<�B�<>�<Q6�<H+�<��<?�<#��<X��<��<���<&}�<~U�<�)�<n��<���<2��<fS�<}�<V��<��<T:�<[��<"��<�:�<���<�z�<(�<���<�:�<nǼ<P�<�Թ<6U�<�Ѷ<VJ�<���<�/�< ��<��<wl�<�Ϋ<.�<ቨ<��<8�<���<pڡ<h'�<�q�<}��<���<�A�<ʂ�<}��<I��<89�<Pr�<ԩ�<�ߌ<a�<�G�<�y�<���<�ڃ<�	�< 8�<��|<!&y<�u<��q<
1n<~�j<��f<h:c<M�_<%�[<�GX<\�T<e Q<�^M<Q�I<�!F<!�B<�><{V;<��7<U24<�0<e-<��)<&<��"<N<t�<�7<��<Og<:<�
<�X<V
<�� <L�;Y��;&�;���;���;�F�;��;���;^��;}��;�;�,�;�a�;ȧ�;���;�g�;[�;�l�;�	�;��;x�;tI�;�Xv;<Al;*Lb;�yX;��N;w9E;#�;;\~2;�P);�C ;�U;�;��;�:���:
��:�\�:>�:f��:|�:�e�:[�q:�S:��4:��:?V�9���9|;{9�T9�7/f����I��A��Eӹ���ڲ�}u:�� U�\o�����������i~���?��[�ĺ׉Ѻg޺А�s���q�����U����h+�v= � J&�TR,�&W2��W8�U>��ND��FJ�V;P�.V�g\�{b���g���m�H�s�
�y����	͂���r������ϧ����������˒��ݍ���  �  �o=�=��=�O=z�=�=.=�� =yk =�	 =6O�<R��<���<&��<�6�<�n�<l��<N��<�<�C�<yv�<��<��<��<|4�<�`�<O��<s��<��<��<&�<rH�<�h�<���<$��<���<��<$��<� �<h�<]!�<�-�<�7�<�>�<�B�<ND�<�B�<>�<N6�<D+�<��<B�<��<`��<��<���<,}�<}U�<�)�<`��<���<4��<dS�<{�<R��<��<F:�<e��<��<�:�<���<�z�<&�<}��<�:�<gǼ<P�<�Թ<7U�<�Ѷ<LJ�<���<�/�<��<��<rl�<�Ϋ<.�<މ�<��<8�<���<xڡ<e'�<�q�<���<���<�A�<Ȃ�<~��<K��<,9�<Yr�<֩�<�ߌ<`�<�G�<�y�<���<�ڃ<�	�<28�<��|<&y<�u<��q<1n<s�j<��f<]:c<e�_<�[<�GX<R�T<f Q<_M<;�I<�!F< �B<��><�V;<��7<P24<#�0<w-<m�)<~&<��"<F<��<�7<��<Gg</<��
<�X<Y
<�� <S�;��;&�;���;c��;.G�;��;���;2��;��;5�;z,�;ya�;���;���;�g�;^�;�l�;�	�;A��;�w�;�I�;�Xv;�@l;"Lb;wyX;n�N;�9E;>�;;�}2;Q);�C ;�U;K�;��;H��:���:��:]�:�:;��:G�:Xe�:��q:�S:��4:��:&Y�9���9�:{9VO9a �7m����I�.C��ӹC��,���u:��U�Zo�<Ä�6�!���t���?����ĺ��ѺV޺L�꺒������Z��l����}+�r= �J&��R,��V2��W8�*U>�OD��FJ��;P�+.V�E\��b�O�g���m�n�s�2�y����̂�������1�������ȟ��͘��ߒ��ۍ���  �  �o=�=��=�O=��=�=
.=�� =xk =�	 =9O�<P��<���<#��<�6�<�n�<q��<I��<�<�C�<wv�<���<��<
�<�4�<�`�<S��<r��<���<��<&�<gH�<�h�<���<#��<���<���<(��<� �<i�<d!�<�-�<�7�<�>�<�B�<ID�<�B�<>�<O6�<S+�<��<F�<��<c��<��<���<%}�<{U�<�)�<c��<���<+��<oS�<�<P��<���<C:�<]��<��<�:�<���<�z�<+�<n��<�:�<bǼ<#P�<�Թ<0U�<�Ѷ<?J�<���<�/�<���<��<vl�<�Ϋ<.�<���<��<(8�<���<pڡ<m'�<�q�<���<���<�A�<ł�<���<J��<.9�<Wr�<ө�<�ߌ<W�<�G�<�y�<���<�ڃ<�	�<"8�<��|<,&y<�u<��q< 1n<g�j<��f<R:c<_�_<
�[<�GX<j�T<X Q<�^M<:�I<�!F<�B<��><�V;<��7<|24<�0<o-<t�)<x&<��"<A<��<�7<��<=g<<<�
<�X<x
<r� <��;��;�%�;���;a��;�F�;��;��;��;|��;�;w,�;�a�;���;���;Yg�;d�;�l�;�	�;��;�w�;|I�;sXv;�Al;%Lb;�yX;��N;:9E;_�;;~2;Q);�C ;�U;�;��;���:Ӓ�:t��:�\�:��:~��:'�:�f�:L�q:�S:}�4:Z�:�U�9M��9�={9�G9E�7�q��7�I�'B���ӹ��ɵ�it:�1U�<\o�lÄ�����爵�q���>����ĺ �Ѻ@޺א����ȭ�/��t�����+�2= �J&��R,��V2��W8��T>�ROD�gFJ�Z;P��.V�?\��b���g��m��s�J�y�!���̂�Å�D���G�������⟑��������������  �  �o=�=��=�O=��=�=.=�� =zk =�	 =BO�<J��<���<1��<�6�<�n�<l��<I��<#�<�C�<yv�<��<��<��<�4�<�`�<Y��<���<���<��<&�<qH�<�h�<���<��<���<���< ��<� �<d�<c!�<�-�<�7�<�>�<�B�<WD�<�B�<>�<N6�<K+�<��<E�< ��<Z��<��<���<)}�<�U�<�)�<i��<���<1��<iS�<|�<S��<��<Q:�<\��<*��<�:�<���<�z�<'�<}��<�:�<aǼ<P�<�Թ<.U�<�Ѷ<KJ�<���<�/�<���<��<l�<�Ϋ<.�<߉�<��<8�<���<rڡ<m'�<�q�<���<���<�A�<ς�<���<D��<79�<Tr�<ة�<�ߌ<Z�<�G�<�y�<���<�ڃ<�	�<!8�<��|<&y<�u<��q<1n<a�j<��f<J:c<S�_<�[<�GX<U�T<p Q<�^M<a�I<�!F<�B<��><|V;<��7<a24<'�0<n-<��)<n&<��"<\<�<�7<��<>g<E<��
<�X<^
<~� <R�;A��;�%�;���;���;�F�;��;���;1��;|��;�;`,�;|a�;���;���;�g�;P�;�l�;�	�;��;5x�;{I�;�Xv;Al;'Lb;yX;��N;�9E;Q�;;?~2;�P);�C ;�U;4�;�;��:>��:k��:�\�:u�:U��:S�:|e�:�q:�S:��4:��:OV�9#��9�;{9�O9���7;r����I�FD��Eӹa��D��Nu:�� U�[\o���^��������~���?����ĺ��ѺE޺���������a�������@+�= �GJ&�_R,�W2��W8��T>�;OD��FJ��;P�G.V�B\�>b���g���m�f�s�Z�y�ʭ��̂�Å�t���V���ħ����֘��ْ��ō���  �  �o=�=�=�O=~�=�=.=�� =�k =�	 =>O�<X��<���<)��<�6�<�n�<o��<W��<�<�C�<�v�<ݧ�<-��<��<�4�<�`�<C��<s��<���<��<&�<wH�<�h�<���<&��<���<��<��<� �<c�<]!�<�-�<�7�<�>�<�B�<^D�<�B�<(>�<S6�<G+�<�<?�<$��<`��<	��<���<!}�<�U�<�)�<q��<���<@��<iS�<}�<i��<��<W:�<M��<��<�:�<���<�z�<!�<z��<{:�<qǼ<P�<�Թ<<U�<�Ѷ<NJ�<쾳<�/�<���<{�<jl�<�Ϋ<.�<މ�<��<8�<���<|ڡ<g'�<�q�<���<���<�A�<ǂ�<���<P��<59�<Or�<驎<�ߌ<i�<�G�<�y�<���<�ڃ<�	�<8�<��|<&y<�u<��q<1n<~�j<��f<e:c<V�_<�[<�GX<K�T<p Q<�^M<I�I<o!F<�B<��><�V;<�7<I24<E�0<k-<}�)<�&<��"<L<r�<�7<��<Yg<7<��
<�X<L
<�� <Y�;?��;�%�;���;f��;�F�;��;���;F��;J��;3�;�,�;|a�;ا�;���;xg�;M�;�l�;�	�;귊;x�;7I�;Yv;Al;�Lb;�yX;��N;:E;"�;;f~2;Q);�C ;oU;��;��;\��:���:��:�]�:x�:c��:��:ne�:��q:�S:��4:Y�:{U�9
��9�8{9N9ĳ7b��W�I��B���ӹ���ٳ��v:�� U��\o��Ä�������~���?���ĺ�Ѻ�޺��y���P��?��&�����+�:= ��I&�mR,�+W2�W8�8U>��ND�5FJ��;P�.V��\��b�!�g���m���s�1�y���͂������� �������쟑�Ę���ƍ���  �  �o=�=��=�O=}�=�=.=�� =zk =�	 =9O�<R��<���<*��<�6�<�n�<s��<J��< �<�C�<yv�<��<��<��<�4�<�`�<X��<|��<���<��<&�<rH�<�h�<���<��<���<���<%��<� �<o�<_!�<�-�<�7�<�>�<�B�<SD�<�B�<>�<B6�<J+�<��<H�<��<d��<��<��<4}�<~U�<�)�<_��<���<0��<iS�<p�<L��<��<M:�<b��<(��<�:�<���<�z�<.�<u��<�:�<cǼ<P�<�Թ<4U�<�Ѷ<HJ�<���<�/�<���<��<~l�<�Ϋ<.�<���<��<8�<���<rڡ<n'�<�q�<���<���<�A�<̂�<���<M��<-9�<Xr�<ة�<�ߌ<P�<�G�<�y�<���<�ڃ<�	�<!8�<��|<&y<�u<��q<1n<\�j<��f<B:c<_�_<
�[<�GX<\�T<Y Q<�^M<R�I<�!F<"�B<��><~V;<��7<^24<&�0<u-<u�)<~&<��"<O<��<�7<��<?g<@<�
<�X<V
<n� <W�;3��;&�;���;���;�F�;��;���;1��;o��;(�;C,�;ta�;���;���;gg�;|�;�l�;�	�;��;)x�;�I�;�Xv;Al;Lb;yX;��N;w9E;n�;;�}2;$Q);�C ;�U;��;��;Ɂ�:���:���:�\�:o�:���:��:{e�:��q:kS:f�4:��:�U�9 ��9�>{9�K9���7qp���I�F���ӹӽ����u:��U�3\o���i���H������?���ĺ�Ѻ1޺������֭���i��>�U+�3= ��I&��R,��V2��W8��T>��OD��FJ��;P�.V�#\�{b���g��m�_�s��y� ���̂�Å�����f�������⟑�����˒��􍚻�  �  �o=�=�=�O=��=�=
.=�� =qk =�	 =EO�<Q��<���< ��<�6�<�n�<{��<G��<2�<�C�<pv�<���<��<�<�4�<�`�<K��<o��<��<��<&�<]H�<�h�<���<��<���<���</��<� �<b�<]!�<�-�<�7�<�>�<�B�<CD�<�B�<>�<X6�<Z+�<��<[�<��<l��<��<���<%}�<vU�<�)�<]��<���<#��<tS�<��<X��<��<@:�<Z��<��<�:�<���<�z�<&�<d��<�:�<ZǼ<$P�<�Թ<1U�<�Ѷ<5J�<���<�/�<��<}�<ll�<�Ϋ<.�<���<��<48�<���<kڡ<�'�<�q�<���<���<�A�<���<���<N��<69�<fr�<ĩ�<�ߌ<\�<�G�<�y�<���<�ڃ<�	�<)8�<��|<&y<�u<��q<-1n<M�j<��f<8:c<k�_<�[<�GX<W�T<b Q<_M<.�I<�!F<��B<�><�V;<��7<�24<�0<�-<��)<{&<��"<:<��<�7<��<9g<d<�
<�X<�
<p� <��;C��;�%�;���;U��;G�;��;��;���;���;*�;R,�;�a�;i��;��;)g�;K�;�l�;�	�;��;�w�;yI�;FXv;�Al;oLb;�yX;�N;�8E;�;;�}2;cQ);�C ;�U;�;��;L��:u��:���:	\�:�::��:��:�f�:�q:mS:��4:T�:�W�9ݫ�9;{9:C9�!�7�y����I�uC��aӹ�����t:��U�k[o��Ä��������d>����ĺ=�ѺP޺�꺪��������������+�$= ��I&�gR,�vV2�:X8�;T>�.OD�&FJ�9;P��.V�{\�b���g���m�k�s���y�W���̂�=Å�A���{�������柑����Ԓ��⍚��  �  �o=�=��=�O=}�=�=.=�� =zk =�	 =9O�<R��<���<*��<�6�<�n�<s��<J��< �<�C�<yv�<��<��<��<�4�<�`�<X��<|��<���<��<&�<rH�<�h�<���<��<���<���<%��<� �<o�<_!�<�-�<�7�<�>�<�B�<SD�<�B�<>�<B6�<J+�<��<H�<��<d��<��<��<4}�<~U�<�)�<_��<���<0��<iS�<p�<L��<��<M:�<b��<(��<�:�<���<�z�<.�<u��<�:�<cǼ<P�<�Թ<4U�<�Ѷ<HJ�<���<�/�<���<��<~l�<�Ϋ<.�<���<��<8�<���<rڡ<n'�<�q�<���<���<�A�<̂�<���<M��<-9�<Xr�<ة�<�ߌ<P�<�G�<�y�<���<�ڃ<�	�<!8�<��|<&y<�u<��q<1n<\�j<��f<B:c<_�_<
�[<�GX<\�T<Y Q<�^M<R�I<�!F<"�B<��><~V;<��7<^24<&�0<u-<u�)<~&<��"<O<��<�7<��<?g<@<�
<�X<V
<n� <W�;3��;&�;���;���;�F�;��;���;1��;o��;(�;C,�;ta�;���;���;gg�;|�;�l�;�	�;��;)x�;�I�;�Xv;Al;Lb;yX;��N;w9E;n�;;�}2;$Q);�C ;�U;��;��;Ɂ�:���:���:�\�:o�:���:��:{e�:��q:kS:f�4:��:�U�9 ��9�>{9�K9���7qp���I�F���ӹӽ����u:��U�3\o���i���H������?���ĺ�Ѻ1޺������֭���i��>�U+�3= ��I&��R,��V2��W8��T>��OD��FJ��;P�.V�#\�{b���g��m�_�s��y� ���̂�Å�����f�������⟑�����˒��􍚻�  �  �o=�=�=�O=~�=�=.=�� =�k =�	 =>O�<X��<���<)��<�6�<�n�<o��<W��<�<�C�<�v�<ݧ�<-��<��<�4�<�`�<C��<s��<���<��<&�<wH�<�h�<���<&��<���<��<��<� �<c�<]!�<�-�<�7�<�>�<�B�<^D�<�B�<(>�<S6�<G+�<�<?�<$��<`��<	��<���<!}�<�U�<�)�<q��<���<@��<iS�<}�<i��<��<W:�<M��<��<�:�<���<�z�<!�<z��<{:�<qǼ<P�<�Թ<<U�<�Ѷ<NJ�<쾳<�/�<���<{�<jl�<�Ϋ<.�<މ�<��<8�<���<|ڡ<g'�<�q�<���<���<�A�<ǂ�<���<P��<59�<Or�<驎<�ߌ<i�<�G�<�y�<���<�ڃ<�	�<8�<��|<&y<�u<��q<1n<~�j<��f<e:c<V�_<�[<�GX<K�T<p Q<�^M<I�I<o!F<�B<��><�V;<�7<I24<E�0<k-<}�)<�&<��"<L<r�<�7<��<Yg<7<��
<�X<L
<�� <Y�;?��;�%�;���;f��;�F�;��;���;F��;J��;3�;�,�;|a�;ا�;���;xg�;M�;�l�;�	�;귊;x�;7I�;Yv;Al;�Lb;�yX;��N;:E;"�;;f~2;Q);�C ;oU;��;��;\��:���:��:�]�:x�:c��:��:ne�:��q:�S:��4:Y�:{U�9
��9�8{9N9ĳ7b��W�I��B���ӹ���ٳ��v:�� U��\o��Ä�������~���?���ĺ�Ѻ�޺��y���P��?��&�����+�:= ��I&�mR,�+W2�W8�8U>��ND�5FJ��;P�.V��\��b�!�g���m���s�1�y���͂������� �������쟑�Ę���ƍ���  �  �o=�=��=�O=��=�=.=�� =zk =�	 =BO�<J��<���<1��<�6�<�n�<l��<I��<#�<�C�<yv�<��<��<��<�4�<�`�<Y��<���<���<��<&�<qH�<�h�<���<��<���<���< ��<� �<d�<c!�<�-�<�7�<�>�<�B�<WD�<�B�<>�<N6�<K+�<��<E�< ��<Z��<��<���<)}�<�U�<�)�<i��<���<1��<iS�<|�<S��<��<Q:�<\��<*��<�:�<���<�z�<'�<}��<�:�<aǼ<P�<�Թ<.U�<�Ѷ<KJ�<���<�/�<���<��<l�<�Ϋ<.�<߉�<��<8�<���<rڡ<m'�<�q�<���<���<�A�<ς�<���<D��<79�<Tr�<ة�<�ߌ<Z�<�G�<�y�<���<�ڃ<�	�<!8�<��|<&y<�u<��q<1n<a�j<��f<J:c<S�_<�[<�GX<U�T<p Q<�^M<a�I<�!F<�B<��><|V;<��7<a24<'�0<n-<��)<n&<��"<\<�<�7<��<>g<E<��
<�X<^
<~� <R�;A��;�%�;���;���;�F�;��;���;1��;|��;�;`,�;|a�;���;���;�g�;P�;�l�;�	�;��;5x�;{I�;�Xv;Al;'Lb;yX;��N;�9E;Q�;;?~2;�P);�C ;�U;4�;�;��:>��:k��:�\�:u�:U��:S�:|e�:�q:�S:��4:��:OV�9#��9�;{9�O9���7;r����I�FD��Eӹa��D��Nu:�� U�[\o���^��������~���?����ĺ��ѺE޺���������a�������@+�= �GJ&�_R,�W2��W8��T>�;OD��FJ��;P�G.V�B\�>b���g���m�f�s�Z�y�ʭ��̂�Å�t���V���ħ����֘��ْ��ō���  �  �o=�=��=�O=��=�=
.=�� =xk =�	 =9O�<P��<���<#��<�6�<�n�<q��<I��<�<�C�<wv�<���<��<
�<�4�<�`�<S��<r��<���<��<&�<gH�<�h�<���<#��<���<���<(��<� �<i�<d!�<�-�<�7�<�>�<�B�<ID�<�B�<>�<O6�<S+�<��<F�<��<c��<��<���<%}�<{U�<�)�<c��<���<+��<oS�<�<P��<���<C:�<]��<��<�:�<���<�z�<+�<n��<�:�<bǼ<#P�<�Թ<0U�<�Ѷ<?J�<���<�/�<���<��<vl�<�Ϋ<.�<���<��<(8�<���<pڡ<m'�<�q�<���<���<�A�<ł�<���<J��<.9�<Wr�<ө�<�ߌ<W�<�G�<�y�<���<�ڃ<�	�<"8�<��|<,&y<�u<��q< 1n<g�j<��f<R:c<_�_<
�[<�GX<j�T<X Q<�^M<:�I<�!F<�B<��><�V;<��7<|24<�0<o-<t�)<x&<��"<A<��<�7<��<=g<<<�
<�X<x
<r� <��;��;�%�;���;a��;�F�;��;��;��;|��;�;w,�;�a�;���;���;Yg�;d�;�l�;�	�;��;�w�;|I�;sXv;�Al;%Lb;�yX;��N;:9E;_�;;~2;Q);�C ;�U;�;��;���:Ӓ�:t��:�\�:��:~��:'�:�f�:L�q:�S:}�4:Z�:�U�9M��9�={9�G9E�7�q��7�I�'B���ӹ��ɵ�it:�1U�<\o�lÄ�����爵�q���>����ĺ �Ѻ@޺א����ȭ�/��t�����+�2= �J&��R,��V2��W8��T>�ROD�gFJ�Z;P��.V�?\��b���g��m��s�J�y�!���̂�Å�D���G�������⟑��������������  �  �o=�=��=�O=z�=�=.=�� =yk =�	 =6O�<R��<���<&��<�6�<�n�<l��<N��<�<�C�<yv�<��<��<��<|4�<�`�<O��<s��<��<��<&�<rH�<�h�<���<$��<���<��<$��<� �<h�<]!�<�-�<�7�<�>�<�B�<ND�<�B�<>�<N6�<D+�<��<B�<��<`��<��<���<,}�<}U�<�)�<`��<���<4��<dS�<{�<R��<��<F:�<e��<��<�:�<���<�z�<&�<}��<�:�<gǼ<P�<�Թ<7U�<�Ѷ<LJ�<���<�/�<��<��<rl�<�Ϋ<.�<މ�<��<8�<���<xڡ<e'�<�q�<���<���<�A�<Ȃ�<~��<K��<,9�<Yr�<֩�<�ߌ<`�<�G�<�y�<���<�ڃ<�	�<28�<��|<&y<�u<��q<1n<s�j<��f<]:c<e�_<�[<�GX<R�T<f Q<_M<;�I<�!F< �B<��><�V;<��7<P24<#�0<w-<m�)<~&<��"<F<��<�7<��<Gg</<��
<�X<Y
<�� <S�;��;&�;���;c��;.G�;��;���;2��;��;5�;z,�;ya�;���;���;�g�;^�;�l�;�	�;A��;�w�;�I�;�Xv;�@l;"Lb;wyX;n�N;�9E;>�;;�}2;Q);�C ;�U;K�;��;H��:���:��:]�:�:;��:G�:Xe�:��q:�S:��4:��:&Y�9���9�:{9VO9a �7m����I�.C��ӹC��,���u:��U�Zo�<Ä�6�!���t���?����ĺ��ѺV޺L�꺒������Z��l����}+�r= �J&��R,��V2��W8�*U>�OD��FJ��;P�+.V�E\��b�O�g���m�n�s�2�y����̂�������1�������ȟ��͘��ߒ��ۍ���  �  �o=�=��=�O=��=�=.=�� =xk =�	 =BO�<S��<���<*��<�6�<�n�<b��<S��<�<�C�<wv�<��<��<��<�4�<�`�<T��<|��< ��<��<&�<}H�<�h�<���<*��<���<	��<��<�<g�<c!�<�-�<�7�<�>�<�B�<ZD�<�B�<>�<Q6�<H+�<��<?�<#��<X��<��<���<&}�<~U�<�)�<n��<���<2��<fS�<}�<V��<��<T:�<[��<"��<�:�<���<�z�<(�<���<�:�<nǼ<P�<�Թ<6U�<�Ѷ<VJ�<���<�/�< ��<��<wl�<�Ϋ<.�<ቨ<��<8�<���<pڡ<h'�<�q�<}��<���<�A�<ʂ�<}��<I��<89�<Pr�<ԩ�<�ߌ<a�<�G�<�y�<���<�ڃ<�	�< 8�<��|<!&y<�u<��q<
1n<~�j<��f<h:c<M�_<%�[<�GX<\�T<e Q<�^M<Q�I<�!F<!�B<�><{V;<��7<U24<�0<e-<��)<&<��"<N<t�<�7<��<Og<:<�
<�X<V
<�� <L�;Y��;&�;���;���;�F�;��;���;^��;}��;�;�,�;�a�;ȧ�;���;�g�;[�;�l�;�	�;��;x�;tI�;�Xv;<Al;*Lb;�yX;��N;w9E;#�;;\~2;�P);�C ;�U;�;��;�:���:
��:�\�:>�:f��:|�:�e�:[�q:�S:��4:��:?V�9���9|;{9�T9�7/f����I��A��Eӹ���ڲ�}u:�� U�\o�����������i~���?��[�ĺ׉Ѻg޺А�s���q�����U����h+�v= � J&�TR,�&W2��W8�U>��ND��FJ�V;P�.V�g\�{b���g���m�H�s�
�y����	͂���r������ϧ����������˒��ݍ���  �  �o=�=��=�O=��=�=	.=�� =xk =�	 =8O�<O��<���<$��<�6�<�n�<l��<I��<�<�C�<zv�<��<��<��<�4�<�`�<T��<z��<���<��<&�<qH�<�h�<���<*��<���<��<$��<� �<f�<l!�<�-�<�7�<�>�<�B�<KD�<�B�<>�<O6�<W+�<��<?�<��<\��<��<��<}�<xU�<�)�<d��<���<*��<sS�<��<O��<���<F:�<V��<��<�:�<���<�z�<'�<z��<�:�<mǼ<%P�<�Թ<6U�<�Ѷ<JJ�<���<�/�<���<��<vl�<�Ϋ<.�<牨<��<&8�<���<kڡ<h'�<�q�<���<���<�A�<Ă�<���<G��<-9�<Lr�<Щ�<�ߌ<W�<�G�<�y�<���<�ڃ<�	�< 8�<��|<2&y<�u<��q<1n<v�j<��f<a:c<[�_<"�[<�GX<o�T<i Q<�^M<N�I<�!F<��B<
�><|V;<��7<~24<�0<[-<q�)<u&<��"<B<g�<�7<��<;g<4<�
<�X<t
<p� <]�;?��;�%�;���;���;�F�;��;��;.��;���;�;�,�;�a�;���;���;�g�;V�;�l�;�	�;��;x�;gI�;�Xv;�Al;�Kb;~yX;��N;39E;!�;;~2;�P);�C ;dU;��;��;'��:ڒ�:���:n\�:�:���:
�:Yf�:��q:�S:�4:��:$V�9Ϯ�9R;{9�M9��7�g����I��@��Iӹ���j���t:�� U�]\o�Ä�����6�����a?����ĺ%�Ѻ޺+��u������W�������+�== �-J&��R,�CW2��W8�{T>�VOD��FJ�:;P��.V�L\��b���g���m��s�G�y�����̂���H���*�����������Ԙ������Ս���  �  �o=�=��=�O=}�=�=	.=�� =uk =�	 =1O�<I��<���<��<�6�<�n�<n��<A��<�<�C�<qv�<��<��<��<4�<�`�<W��<s��<��<��<&�<sH�<�h�<���<&��<���<��<*��<� �<n�<b!�<�-�<�7�<�>�<�B�<JD�<�B�<>�<J6�<F+�<��<H�<
��<_��<���<���<)}�<tU�<�)�<T��<���<*��<dS�<x�<O��<��<C:�<j��<��<�:�<���<�z�</�<}��<�:�<kǼ<P�<�Թ<:U�<�Ѷ<LJ�<���<�/�<��<��<xl�<�Ϋ<.�<䉨<��<8�<���<rڡ<h'�<�q�<���<���<�A�<�<}��<D��<$9�<Yr�<ͩ�<�ߌ<W�<�G�<�y�<���<�ڃ<�	�<28�<��|<%&y<�u<��q<(1n<r�j<��f<[:c<k�_<�[<�GX<e�T<c Q<_M<>�I<�!F<�B<��><�V;<��7<W24<�0<t-<c�)<i&<��"<8<��<�7<��<+g</<�
<�X<X
<p� <\�;��;&�;���;a��;%G�;��;��;2��;���;7�;�,�;�a�;���;��;�g�;t�;�l�;�	�;B��;�w�;�I�;vXv;"Al;Lb;[yX;v�N;'9E;g�;;�}2;�P);\C ;�U;6�;h�;]��:���:k��:p\�:�:
��:	�:�e�:M�q:JS:��4:��:>X�9]��9�>{9O9��7'i���I��A��sӹ���8���t:��U�]Zo�:Ä������������?����ĺ��Ѻ�޺���p�����=��������+�u= �CJ&��R,��V2��W8�U>�SOD��FJ��;P�.V��\��b�J�g���m�9�s��y����̂���Y���6���������Ę������ፚ��  �  �o=�=��=�O=��=�=.=�� ={k =�	 =6O�<N��<���<��<�6�<�n�<f��<L��<�<�C�<zv�<��<$��<��<�4�<�`�<R��<v��<��<��<&�<{H�<�h�<���</��<���<��<#��<� �<m�<e!�<�-�<�7�<�>�<�B�<VD�<�B�<>�<Q6�<F+�<��<A�<��<\��<���<��<}�<sU�<�)�<c��<���<0��<fS�<|�<^��<��<R:�<Y��<��<�:�<���<�z�<.�<���<�:�<zǼ<"P�<�Թ<CU�<�Ѷ<TJ�<���<�/�<��<��<wl�<�Ϋ<.�<䉨<��<8�<���<pڡ<c'�<�q�<���<���<�A�<���<y��<F��<-9�<Or�<ܩ�<�ߌ<g�<�G�<�y�<���<�ڃ<�	�<%8�<��|<+&y<�u<��q<!1n<��j<��f<v:c<g�_<�[<�GX<e�T<k Q<�^M<D�I<�!F<�B<��><�V;<��7<V24<,�0<_-<m�)<t&<��"<0<q�<�7<��<Bg<(<�
<�X<U
<�� <[�;A��;�%�;���;n��;�F�;��;��;T��;q��;O�;�,�;�a�;���;���;�g�;q�;�l�;�	�;��;x�;iI�;�Xv;7Al;mLb;�yX;t�N;{9E;2�;;~2;�P);RC ;JU;Ӆ;d�;��:Ӓ�:��:�\�:5�:N��: �:�e�:�q:)S:2�4:��:W�9̭�9;>{9�Q9���7(Z��t�I��@��;ӹ���4���t:�� U�v[o�$Ä����������~���?����ĺ�Ѻ<޺ݐ��������������	��+��= �4J&��R,�2W2�~W8�U>��ND�pFJ�p;P�I.V�^\��b���g���m� �s���y����̂���\�����������՟����������э���  �  �o=�=��=�O=��=ߎ=.=�� ={k =�	 =;O�<C��<���<(��<�6�<�n�<`��<E��<�<�C�<yv�<٧�<��<��<�4�<�`�<a��<���<���<��<&�<zH�<�h�<���<&��<���<��<'��<
�<g�<r!�<�-�<�7�<�>�<�B�<YD�<�B�<
>�<B6�<A+�<��<8�<��<N��<	��<���<}�<�U�<�)�<b��<���<,��<bS�<o�<N��<��<W:�<W��<7��<�:�<���<�z�<(�<���<�:�<tǼ<P�<�Թ<=U�<�Ѷ<WJ�<���<�/�<���<��<�l�<�Ϋ<.�<҉�<��<8�<���<jڡ<d'�<�q�<w��<���<�A�<Ƃ�<���<:��<29�<Er�<ک�<�ߌ<Z�<�G�<�y�<���<�ڃ<�	�<8�<��|<1&y<�u<��q<$1n<��j<��f<h:c<f�_<-�[<�GX<f�T<� Q<�^M<l�I<�!F<�B<�><]V;<��7<I24<+�0<R-<w�)<^&<��"<I<i�<�7<��<4g<1<ڬ
<�X<A
<}� <�;_��;�%�;��;���;�F�;�;���;P��;���;9�;�,�;�a�;ߧ�;���;�g�;Y�;m�;�	�;��;gx�;gI�;�Xv;�@l;�Kb;yX;P�N;f9E;��;;~2;oP);�C ;rU;�;��;<��:Ē�:���:�\�:��:|��:��:�d�:��q:�S:�4:��:�W�9\��96;{9�V9-�7�`����I��B���ӹ������u:���T�.\o����������;~���@����ĺ��Ѻ`޺<�꺨��������9����+�W= ��J&��R,�W2��W8�AU>�;OD�GJ�y;P�T.V�?\��b��g�o�m��s�"�y�~���̂���w���������������������������  �  �o=�=��=�O=��=�=.=�� =uk =�	 =;O�<H��<���<��<�6�<�n�<l��<A��<!�<�C�<rv�<��<��< �<�4�<�`�<Q��<k��<��<��<&�<qH�<�h�<���<.��<���<��<.��<� �<n�<e!�<�-�<�7�<�>�<�B�<RD�<�B�<>�<Q6�<F+�<��<D�<��<X��<���<��<}�<vU�<�)�<]��<���<*��<eS�<}�<^��<���<M:�<Y��<��<�:�<���<�z�</�<y��<�:�<nǼ</P�<�Թ<<U�<�Ѷ<JJ�<���<�/�<��<z�<tl�<�Ϋ<.�<艨<��<8�<���<mڡ<o'�<�q�<���<���<�A�<���<���<B��<.9�<Qr�<Ω�<�ߌ<a�<�G�<�y�<���<�ڃ<�	�<!8�<��|<,&y<�u<��q<,1n<w�j<��f<f:c<j�_<�[<�GX<l�T<j Q<�^M<5�I<�!F<�B<	�><�V;<��7<V24<�0<e-<w�)<g&<��"<&<h�<�7<��<,g<?<�
<�X<U
<�� <l�;I��;�%�;���;@��;�F�;��;��;*��;���;;�;�,�;�a�;���;��;vg�;u�;�l�;�	�;���;�w�;mI�;�Xv;kAl;lLb;�yX;v�N;89E;H�;;�}2;�P);uC ;U;��;v�;��:o��:k��:r\�:"�:\��:��:(f�:��q: S:S�4:��:FW�9v��9�>{99M9�)�7�f���I�.?���ӹ?��q��bt:�� U��[o��Ä� ������~��J?���ĺ�Ѻ�޺������	��R������,�[= �YJ&��R,�$W2��W8�U>�OD�oFJ�J;P�j.V�P\��b���g���m� �s�	�y�׭��̂�����������������Ø������Ӎ���  �  qn=j=I�=�M=M�=w�=W+=�� ==h =? =�G�<8��< ��<���<-�<'d�<p��<���<��<�6�<�h�<���<��<T��<$�<�O�<oy�<ȡ�<���<���<�<~2�<5R�<�o�<���<S��<���<	��<���<q��<g�<��<��<��<L!�<�!�<A�<��<��<�<���<m��<j��<��<ɖ�<
v�<�Q�<2)�<��<���<��<�`�<�$�<\��<��<`W�<~
�<���<>d�<�
�<��<�J�<���<bz�<��<%��<i"�<���<�(�<֥�<�<���<5�<ht�<�ޮ<�E�<,��<L	�<Hf�<�<��<�j�<n��<�	�<4U�<I��<��<N)�<^k�<u��<��<�%�<M`�<��<rЌ<T�<�:�<^n�<���<҃<��<i2�<��|<�y<1|u<��q</3n<��j<8�f<ZDc<C�_<��[<�YX<K�T<�Q<yM<=�I<PAF<c�B<�?<=~;<>�7<r_4<��0<�M-<v�)<K&<��"<	Y<�<ny<7<�<�P<��
<��<�Z<�<���;�:�;V��;?��;h;�;��;��;���;���;ݼ�;�ҽ;Y��;�0�;	x�;Ѧ;>:�;p��;A�;uސ;;��;�L�;��;!�w;#�m;$�c;�Z;odP;	�F;(_=;�4;��*;��!;/�;��;�F;dX�:�[�:���:��:ݯ�:`��:���:�Պ:ȃv:��W:�K9:#4:���9��9$��9�9,Y8�H��W�;��q��4�̹ ��@���7��+R��l�r���}���s��3U��!����ú��к�ݺʡ����4A��n�������b�����i�%�i,��2��8��>�zD��J��
P�V�y�[���a���g�"�m��s���y�_���ł�轅�ϵ��Ю��ç�����؜������핚��  �  `n=e=F�=�M=R�=y�=^+=�� =Bh =; =�G�<=��< ��<���<-�</d�<n��<���<��<�6�<�h�<���<%��<O��<"$�<�O�<my�<���<���<���< �<�2�<8R�<�o�<���<I��<���<���<���<j��<t�<��<��<��<H!�<�!�<C�<��<
�<!�<���<g��<p��<��<і�<v�<�Q�<<)�<��<���<��<�`�<�$�<g��<���<[W�<�
�<���<8d�<�
�<��<K�<���<jz�<��<"��<_"�<~��<�(�<ե�<�<���<E�<Tt�<�ޮ<�E�<+��<W	�<@f�<��<��<�j�<r��<�	�<9U�<G��<��<C)�<bk�<x��<��<�%�<F`�<"��<sЌ<a�<�:�<fn�<���<҃<��<E2�<��|<�y<*|u<��q<3n<��j<$�f<VDc<-�_<��[<�YX<N�T<�Q<;yM<(�I<CAF<k�B<?<C~;<Z�7<q_4<��0<�M-<��)<K&<��"<Y<��<~y<2<!�<�P<��
<��<�Z<
<���;�:�;Z��;4��;6;�;h�;^��;���;ʶ�;��;�ҽ;M��;x0�;x�;�Ц;j:�;T��;EA�;�ސ;���;�L�;��;~�w;/�m;��c;�Z;�dP;|�F;�^=;4;��*;!�!;B�;��;�F;PX�:(\�:T��:n	�:%��:��:Ǘ�:�Պ:&�v:�W:*K9:1:���9��9֣�91�9dD8�K��a�;�xr���̹B�����S�7��)R���l�
s��~���s���T���!��n�ú��к�ݺ������
A��n�8��Z��@�����D�%�2,�-2�38��>�D��J��
P��V���[�A�a�
�g���m�¼s���y�"���ł�轅�����ڮ��������圔����������  �  ^n=t=F�=�M=P�=r�=^+=�� =Fh =7 =�G�<9��<���<���<�,�<5d�<g��<���<��<�6�<�h�<���<&��<<��<"$�<|O�<uy�<ա�<���<���<��<�2�<4R�<�o�<���<H��<���<���<���<^��<p�<��<��<��<C!�<�!�<3�<��<�<�<���<^��<q��<��<ϖ�<v�<�Q�<>)�<	��<���<���<�`�<�$�<`��<���<JW�<�
�<{��<Ld�<�
�< ��<K�<���<uz�<��<+��<^"�<���<�(�<Х�<�<���<L�<Lt�<�ޮ<�E�<%��<Y	�<,f�<
��<��<�j�<s��<�	�<7U�<?��<��<7)�<fk�<s��<��<�%�<<`�<)��<iЌ<a�<�:�<^n�<���<҃<��<C2�<��|<�y<#|u<��q<�2n<�j<$�f<pDc<�_<��[<�YX<8�T<Q<1yM<b�I<EAF<j�B<?<'~;<[�7<`_4<��0<�M-<�)<K&<��"<Y<��<�y<%<�<�P<��
<��<�Z<<_��;�:�;H��;U��;�;�;A�;���;���;߶�;ۼ�;�ҽ;l��;s0�;3x�;�Ц;�:�;$��;3A�;�ސ;֌�;�L�;��;��w;��m;y�c;�Z;WdP;��F;�^=; 4;��*;�!;;�;��;�F;�W�:1\�:���:�	�:ϯ�:���:���:jԊ:��v:�W:�M9:v2:���9��9V��9��9N28�B����;��q����̹Տ����܁7��(R���l��q��M}��?t��cT���"��M�ú�к�ݺ���]��A�o�����������l�%�3,��2��8�!>�D�J��
P��V���[�l�a��g���m��s�ìy����ł����������������ꡑ�㜔�Ę�������  �  cn=j=>�=�M=S�=x�=^+=�� =Bh =9 =�G�<?��<��<���<-�<4d�<t��<���<��<�6�<�h�<���<��<P��<"$�<~O�<^y�<ǡ�<���<���<��<�2�</R�<�o�<���<A��<���<���<���<f��<n�<��<��<��<?!�<�!�<B�<��<
�<#�<���<i��<l��<��<і�<v�<�Q�<=)�<��<���<��<�`�<�$�<e��<���<]W�<�
�<x��<3d�<�
�<���<�J�<���<lz�<��<'��<\"�<���<�(�<ͥ�<�<���<C�<Ot�<�ޮ<�E�<$��<Y	�<Af�<��<��<�j�<p��<�	�<:U�<L��<��<A)�<fk�<z��<��<�%�<D`�<��<pЌ<b�<�:�<gn�<���<҃<��<O2�<��|<�y<5|u<��q<�2n<�j<�f<hDc<�_<��[<�YX<=�T<�Q<EyM<;�I<#AF<r�B<?<=~;<Y�7<j_4<��0<�M-<z�)<K&<��"<Y<��<�y<><!�<�P<��
<��<�Z<�<���;�:�;O��;���;d;�;b�;[��;���;��;ļ�;�ҽ;i��;U0�;x�;�Ц;t:�;E��;,A�;mސ;茋;�L�;w�;��w;*�m;��c;�Z;�dP;X�F;_=;�4;��*;"�!;B�;��;�F;�X�:\�:_��:	�:b��:ꊪ:���:�Պ:օv:��W:�J9:12:���9q�9_��9C�9�18%F����;��q����̹M����ހ7��)R�1�l�er���~��Jt��`T��~!����ú׃кDݺ�����A��n���i����}��%�%�S,�C2�K8��>�D��J��
P��V��[��a���g���m��s�{�y�#���ł�Ƚ���������������Ĝ�����������  �  dn=g=I�=�M=L�=x�=X+=�� =@h =? =�G�<A��<��<���<-�<)d�<r��<���<��<�6�<�h�<���<��<S��<$�<�O�<ry�<ġ�<���<���<��<2�<7R�<�o�<���<E��<���<��<���<k��<u�<��<��<��<Y!�<�!�<=�<��<��<$�<���<u��<e��<��<Ӗ�<v�<�Q�<<)�<��<���<���<�`�<�$�<^��<��<ZW�<�
�<���<:d�<�
�<���<K�<���<iz�<��<$��<Z"�<~��<�(�<֥�<�<���<C�<Tt�<�ޮ<�E�<<��<H	�<Cf�<���<��<�j�<p��<�	�<3U�<J��<��<C)�<^k�<y��<��<�%�<Q`�<��<wЌ<V�<�:�<\n�<���<҃<��<P2�<��|<�y<,|u<��q<3n<
�j<�f<aDc<0�_<��[<�YX<G�T<�Q<JyM<.�I<RAF<{�B<�?<@~;<A�7<x_4<��0<�M-<��)<!K&<��"<Y<��<ry<:<�<�P<��
<��<�Z<�<���;x:�;���;I��;V;�;q�;J��;���;Ķ�;��;�ҽ;Y��;f0�;x�;�Ц;o:�;Y��;FA�;fސ;茋;�L�;��;T�w;�m;a�c;�Z;�dP;4�F;e_=;�4;�*;-�!;9�;��;�F;�X�:�[�:��:��:Y��:���:3��:fՊ:�v:$�W:wK9:;2:m��9��9Z��9��9 O8kI����;�nr����̹�����7��)R���l�~r���}���r��nU��`!���ú��к�ݺ���o��9A��n�^��[��^������%�F,��2�m8��>�mD��J�P��V�=�[�@�a���g��m�߼s���y�!���ł�ѽ�����î��駎�������������ϕ���  �  an=n=D�=�M=N�=|�=\+=�� =Bh =; =�G�<;��<��<���<-�<9d�<s��<���<��<�6�<�h�<���<#��<S��<$�<|O�<jy�<͡�<���<���<��<~2�<2R�<�o�<���<B��<���<���<���<]��<q�<��<��<��<E!�<�!�<?�<��<�<!�<���<m��<o��<��<ז�<v�<�Q�<D)�<��<���<��<�`�<�$�<^��<���<ZW�<�
�<~��<@d�<�
�<���<K�<���<jz�<��<'��<W"�<y��<�(�<ϥ�<�<���<H�<Lt�<�ޮ<�E�<%��<N	�<Bf�<
��<��<�j�<u��<�	�<6U�<I��<��<@)�<hk�<y��<��<�%�<H`�<!��<uЌ<\�<;�<`n�<���<҃<��<K2�<��|<�y<|u<��q<3n<	�j<�f<`Dc<�_<��[<�YX<C�T<�Q<>yM<I�I<>AF<]�B< ?<P~;<Q�7<w_4<��0<�M-<��)<K&<��"<"Y<��<�y<=<�<�P<��
<��<�Z<<���;�:�;H��;+��;|;�;W�;j��;���;���;Ӽ�;�ҽ;H��;]0�; x�;�Ц;s:�;��;8A�;Zސ;�;�L�;��;J�w;�m;��c;�Z;�dP;w�F;$_=;4;��*;R�!;A�;��;G;}X�:\�:���:a	�:��:���:��:qՊ:b�v:w�W:JL9:�2:���9��9⠅9V�9�58�F����;��s����̹���ʤ�N�7�&)R���l�
r���}��5t��U��o!��I�ú��к�ݺb����� A��n���m�������W�%�3,�#2�78��>�@D�xJ��
P��V���[���a���g���m��s�ݬy����ł�ӽ�����Ů����������������������  �  \n=l=A�=�M=R�=u�=\+=�� =Gh =; =�G�<>��<��<���<�,�<;d�<l��<���<��<�6�<�h�<���< ��<D��<,$�<�O�<dy�<š�<���<���<��<�2�<(R�<�o�<���<8��<���<���<���<]��<x�<��<��<��<=!�<�!�<8�<��<�<�< ��<f��<u��<��<ۖ�<v�<�Q�<H)�<��<��<��<�`�<�$�<_��<��<PW�<�
�<w��<:d�<�
�<���<	K�<���<pz�<��<-��<Q"�<y��<�(�<ť�<�<���<N�<Ht�<�ޮ<�E�<&��<e	�<4f�<��<��<�j�<}��<�	�<?U�<C��<��<9)�<jk�<{��<��<�%�<E`�<+��<mЌ<\�<�:�<bn�<���<҃<��<@2�<��|<�y<|u<��q<�2n<�j<�f<hDc<�_<��[<�YX<;�T<Q<*yM<A�I</AF<}�B<?<2~;<S�7<f_4<��0<�M-<��)<K&<��"<&Y<��<�y<0<,�<�P<��
<��<�Z<<���;�:�;`��;��;\;�;>�;���;���;ݶ�;���;�ҽ;S��;40�;<x�;�Ц;�:�;��;SA�;fސ;Ɍ�;�L�;r�; x;��m;�c;�Z;gdP;��F;�^=;C4;��*;m�!;:�;��;3G;X�:�\�:.��:�	�:寺:���:���:�Ԋ:��v:��W:|K9:�1:���9-�92��9��9g&8�?���;��s��V�̹5��ģ�
�7�R(R��l�zr��N~��!t���S��B"����ú$�к�ݺ��.���@��n�ȕ������r��F�%�!,�62��8�>�AD�J��
P�QV���[���a�4�g���m���s�Ԭy�.���ł�����=�������������휔����������  �  `n=k=H�=�M=L�=x�=_+=�� =Dh => =�G�<E��<��<���<-�<6d�<p��<���<��<�6�<�h�<���<#��<M��<$�<�O�<uy�<š�<���<���<��<�2�<'R�<�o�<���<>��<���<���<���<c��<o�<��<��<��<J!�<�!�<9�<��<
�<�<���<l��<m��<��<Ԗ�<v�<�Q�<A)�<��<���<��<�`�<�$�<h��<���<VW�<�
�<���<Ad�<�
�<���<K�<���<hz�<��<)��<T"�<x��<�(�<ƥ�<�<���<D�<Mt�<�ޮ<�E�<+��<L	�<=f�<��<��<�j�<w��<�	�<=U�<G��<��<E)�<fk�<{��<��<�%�<J`�<$��<uЌ<c�<�:�<Zn�<���<҃<��<I2�<��|<�y<%|u<��q<3n<�j<�f<cDc< �_<{�[<�YX<9�T<�Q<:yM<A�I<MAF<h�B<�?<?~;<]�7<y_4<��0<�M-<z�)<)K&<��"<Y<��<�y<7<,�<�P<��
<��<�Z<<���;�:�;b��;Y��;[;�;Z�;a��;���;Ͷ�;���;�ҽ;M��;M0�;)x�;�Ц;]:�;;��;3A�;Xސ;ڌ�;�L�;��;W�w;��m;��c;Z;�dP;��F;#_=;4;�*;=�!;H�;��;�F;�X�:!\�:}��:�	�:��: ��:嗚:,Պ:r�v:�W:fL9:�1:���9�9�9��948�C��t�;��s��?�̹�����[�7��)R�f�l��r���}���s��*U���!��\�úq�к�ݺ<��<���@��n����G����u����%�T,�2�"8��>�D��J�P��V�v�[���a���g���m��s���y�b���ł�ǽ������������$���朔�Ø�������  �  `n=g=E�=�M=T�=|�=X+=�� =?h =? =�G�<G��<��<���<-�<6d�<}��<���<��<�6�<�h�<���<��<\��<$�<O�<hy�<���<���<���<��<}2�<2R�<�o�<���<@��<���<���<���<i��<i�<��<��<��<K!�<�!�<O�<��<�<(�<���<x��<l��<���<Ӗ�<v�<�Q�<>)�<!��<���<���<�`�<�$�<b��<���<kW�<~
�<���<4d�<�
�<���<�J�<���<`z�<��<��<V"�<v��<�(�<ϥ�<�<���<<�<Pt�<�ޮ<�E�<)��<P	�<Of�<���<��<�j�<{��<�	�<<U�<V��<��<G)�<jk�<~��<��<�%�<P`�<��<|Ќ<X�< ;�<nn�<���<҃<��<H2�<��|<�y</|u<��q<3n<�j<�f<BDc<�_<��[<�YX<C�T<�Q<;yM<.�I<AAF<\�B<?<Q~;<C�7<�_4<��0<�M-<��)<-K&<��"<!Y<��<�y<R<+�<�P<��
<��<�Z<�<��;�:�;W��;#��;K;�;f�;E��;���;���;Լ�;�ҽ;5��;W0�;�w�;�Ц;J:�;R��;A�;fސ;݌�;�L�;��;,�w;��m;��c;�Z;�dP;{�F;}_=;�4;N�*;6�!;k�;��;�F;VY�:
\�:G��:�	�:���:ʊ�:���:�֊:�v:��W:�J9:�1:��9E�9���9��9�;8�M��o�;�It����̹ۏ����C�7��*R��l��r��a~���s���T��� ���ú~�к�ݺ���m���@�Cn���9�����\����%�:,��2�c8��>�[D��J�s
P�V�{�[�7�a���g�	�m��s���y�`���ł�	������ ���������ܜ������ϕ���  �  ]n=m=E�=�M=P�=r�=[+=�� =Bh == =�G�<C��<��<���<-�<8d�<n��<���<��<�6�<�h�<���<��<B��< $�<�O�<gy�<̡�<���<���<��<}2�<.R�<�o�<���<>��<���<���<���<_��<j�<��<��<��<J!�<�!�<6�<��<�<#�<���<o��<q��<��<Ֆ�<v�<�Q�<B)�<��<���<��<�`�<�$�<b��<��<PW�<�
�<���<;d�<�
�<���<�J�<���<hz�<��<#��<T"�<x��<�(�<˥�<�<���<@�<Mt�<�ޮ<�E�<.��<W	�<5f�<���<��<�j�<t��<�	�<=U�<F��<��<A)�<nk�<v��<��<�%�<L`�<!��<xЌ<^�<�:�<^n�<���<҃<��<C2�<��|<�y<|u<��q<3n<�j<�f<YDc<"�_<��[<�YX<2�T<�Q</yM<G�I<?AF<y�B<?<&~;<P�7<�_4<��0<�M-<��)<%K&<��"<(Y<��<�y<4<+�<�P<��
<��<�Z<�<{��;�:�;z��;#��;x;�;M�;U��;���;���;ļ�;�ҽ;M��;O0�;x�;�Ц;j:�;+��;A�;|ސ;݌�;�L�;��;��w;��m;=�c;�Z;�dP;r�F;;_=;*4;��*;B�!;��;��;G;�X�:H\�:ė�:>	�:8��:���:��:�Ԋ:хv:N�W:�K9:O2:u��9��9䠅9��978,I��k�;��s���̹k�� ����7�*R�n�l�r��.~���s���T��;"��	�ú��кݺj�麔���@��n����h���������%��,��2�88��>�0D�'J��
P��V���[���a��g���m�*�s�׬y�P���ł�ܽ�����Ү������������И�������  �  [n=n=>�=�M=N�=z�=d+=�� =Hh =; =�G�<I��<��<���<-�<?d�<n��<���<��<�6�<�h�<���<0��<M��<$�<~O�<by�<ʡ�<~��<���<��<�2�<#R�<�o�<���<6��<���<���<���<Y��<n�<��<��<��<5!�<�!�<8�<��<�<"�<���<h��<x��<��<ٖ�<v�<�Q�<D)�<��<��<��<�`�<�$�<g��<��<SW�<�
�<o��<<d�<�
�<���<K�<���<hz�<��<$��<O"�<w��<�(�<���<�<��<K�<Et�<�ޮ<�E�<"��<T	�<;f�<��<��<�j�<u��<�	�<FU�<F��<��<J)�<pk�<y��<��<�%�<F`�<+��<nЌ<m�<;�<\n�<���<�у<��<A2�<��|<�y<|u<��q<�2n<	�j<��f<_Dc<�_<w�[<�YX<(�T<Q<%yM<K�I<"AF<q�B< ?<I~;<t�7<k_4<��0<�M-<��)<2K&<��"</Y<��<�y<3<=�<�P<��
<��<�Z<"<���;�:�;T��;��;q;�;2�;���;���;Ӷ�;���;�ҽ;H��;.0�;x�;�Ц;b:�;��;.A�;^ސ;Ќ�;�L�;R�;��w;��m; �c;#Z;�dP;��F;�^=;a4;�*;b�!;��;��;G;�X�:�\�:=��:�	�:{��:��:���:Պ:Åv:��W:�K9:�1:A��9}�9���9��9�8�H����;��s��G�̹ő�H��+�7��(R�c�l�Or��_~��^t���T���!����ú�к
ݺY�����@��n�ɕ������}����%�,�,2��8��>��D��J�P��V�*�[���a�/�g���m�8�s�ݬy�l��Ƃ�ӽ��H���Ǯ��*���-����䘗������  �  _n=m=E�=�M=O�=y�=V+=�� =Ch =A =�G�<G��<
��<���<-�<1d�<z��<���<��<�6�<�h�<���<��<O��<$�<�O�<my�<ˡ�<���<���<��<�2�<)R�<�o�<���<A��<���<���<���<a��<n�<��<��<��<H!�<�!�<?�<��<��<)�<���<t��<o��<���<Ֆ�<v�<�Q�<=)�<��<���<���<�`�<�$�<Y��<��<YW�<�
�<���<=d�<�
�<���<K�<���<iz�<��< ��<V"�<w��<�(�<ǥ�<�<���<D�<Lt�<�ޮ<�E�<0��<S	�<@f�<���<��<�j�<|��<�	�<;U�<R��<��<K)�<fk�<~��<��<�%�<R`�<!��<xЌ<R�<�:�<_n�<���<҃<��<G2�<��|<�y<#|u<��q<�2n<��j<�f<RDc<�_<~�[<�YX<5�T<�Q<7yM<I�I<AAF<u�B<?<D~;<;�7<z_4<��0<�M-<��)<.K&<��"<Y<��<�y<K<*�<�P<��
<��<�Z<�<���;�:�;z��;:��;u;�;S�;`��;���;Ѷ�;���;�ҽ;>��;Y0�;x�;�Ц;h:�;4��;-A�;cސ;쌋;�L�;��;��w;�m;~�c;�Z;�dP;�F;c_=;4;=�*;B�!;q�;��;�F;Y�:&\�:��:�	�:���:/��:_��:nՊ:<�v:��W:�K9:�2:G��9S�9項9S�9�.8sL���;��s��l�̹Ԑ�t��
�7��)R�x�l�r���}��|s���T���!���ú0�кEݺ��w���@�gn�4������U����%�<,��2�58��>��D��J��
P��V���[���a���g���m�*�s���y�M���ł�����ᮋ�������蜔�˘�������  �  ^n=e=E�=�M=N�=}�=[+=� =;h =A =�G�<C��<��<���<-�<0d�<���<���<��<�6�<�h�<���<"��<R��<$�<�O�<cy�<���<���<���<��<{2�<%R�<�o�<���<I��<���<���<���<b��<f�<��<��<��<P!�<�!�<A�<��<�<8�<���<|��<h��<���<Ֆ�<v�<�Q�<@)�<&��<���<���<�`�<�$�<o��<���<^W�<~
�<���<+d�<�
�<���<�J�<���<cz�<��<��<Z"�<s��<�(�<ƥ�<�<���<5�<It�<�ޮ<�E�<,��<F	�<Cf�<��<��<�j�<p��<�	�<0U�<_��<��<U)�<hk�<���<��<�%�<U`�<��<�Ќ<^�<�:�<^n�<���<҃<~�<C2�<��|<�y<|u<��q<3n<�j<1�f<IDc<�_<x�[<�YX<C�T<�Q<4yM<)�I<AAF<b�B<�?<R~;<O�7<�_4<��0<�M-<��)<%K&<�"<Y<�<�y<g<�<�P<��
<��<�Z<<���;x:�;^��;��;G;�;N�;)��;���;���;���;�ҽ;,��;{0�;�w�;�Ц;R:�;7��;A�;]ސ;ό�;YL�;��;;�w;*�m;��c;Z;IeP;�F;�_=;�4;b�*;E�!;��;;�;�F;�Y�:�[�:���:~�:!��:���:Ɨ�:�Պ:ۃv:üW:�I9:1:2��9t�9u��9F�9?18�V��b�;��t����̹���:���7�f+R�ןl��r���~���s���U��U!����ú
�к�ݺ�����NA��m�3��ʶ���8����%�A,��2��8��>�,D��J��
P��V�x�[�h�a��g���m��s�Ьy�b���ł�	���ݵ��󮋻���*�����������ܕ���  �  _n=m=E�=�M=O�=y�=V+=�� =Ch =A =�G�<G��<
��<���<-�<1d�<z��<���<��<�6�<�h�<���<��<O��<$�<�O�<my�<ˡ�<���<���<��<�2�<)R�<�o�<���<A��<���<���<���<a��<n�<��<��<��<H!�<�!�<?�<��<��<)�<���<t��<o��<���<Ֆ�<v�<�Q�<=)�<��<���<���<�`�<�$�<Y��<��<YW�<�
�<���<=d�<�
�<���<K�<���<iz�<��< ��<V"�<w��<�(�<ǥ�<�<���<D�<Lt�<�ޮ<�E�<0��<S	�<@f�<���<��<�j�<|��<�	�<;U�<R��<��<K)�<fk�<~��<��<�%�<R`�<!��<xЌ<R�<�:�<_n�<���<҃<��<G2�<��|<�y<#|u<��q<�2n<��j<�f<RDc<�_<~�[<�YX<5�T<�Q<7yM<I�I<AAF<u�B<?<D~;<;�7<z_4<��0<�M-<��)<.K&<��"<Y<��<�y<K<*�<�P<��
<��<�Z<�<���;�:�;z��;:��;u;�;S�;`��;���;Ѷ�;���;�ҽ;>��;Y0�;x�;�Ц;h:�;4��;-A�;cސ;쌋;�L�;��;��w;�m;~�c;�Z;�dP;�F;c_=;4;=�*;B�!;q�;��;�F;Y�:&\�:��:�	�:���:/��:_��:nՊ:<�v:��W:�K9:�2:G��9S�9項9S�9�.8sL���;��s��l�̹Ԑ�t��
�7��)R�x�l�r���}��|s���T���!���ú0�кEݺ��w���@�gn�4������U����%�<,��2�58��>��D��J��
P��V���[���a���g���m�*�s���y�M���ł�����ᮋ�������蜔�˘�������  �  [n=n=>�=�M=N�=z�=d+=�� =Hh =; =�G�<I��<��<���<-�<?d�<n��<���<��<�6�<�h�<���<0��<M��<$�<~O�<by�<ʡ�<~��<���<��<�2�<#R�<�o�<���<6��<���<���<���<Y��<n�<��<��<��<5!�<�!�<8�<��<�<"�<���<h��<x��<��<ٖ�<v�<�Q�<D)�<��<��<��<�`�<�$�<g��<��<SW�<�
�<o��<<d�<�
�<���<K�<���<hz�<��<$��<O"�<w��<�(�<���<�<��<K�<Et�<�ޮ<�E�<"��<T	�<;f�<��<��<�j�<u��<�	�<FU�<F��<��<J)�<pk�<y��<��<�%�<F`�<+��<nЌ<m�<;�<\n�<���<�у<��<A2�<��|<�y<|u<��q<�2n<	�j<��f<_Dc<�_<w�[<�YX<(�T<Q<%yM<K�I<"AF<q�B< ?<I~;<t�7<k_4<��0<�M-<��)<2K&<��"</Y<��<�y<3<=�<�P<��
<��<�Z<"<���;�:�;T��;��;q;�;2�;���;���;Ӷ�;���;�ҽ;H��;.0�;x�;�Ц;b:�;��;.A�;^ސ;Ќ�;�L�;R�;��w;��m; �c;#Z;�dP;��F;�^=;a4;�*;b�!;��;��;G;�X�:�\�:=��:�	�:{��:��:���:Պ:Åv:��W:�K9:�1:A��9}�9���9��9�8�H����;��s��G�̹ő�H��+�7��(R�c�l�Or��_~��^t���T���!����ú�к
ݺY�����@��n�ɕ������}����%�,�,2��8��>��D��J�P��V�*�[���a�/�g���m�8�s�ݬy�l��Ƃ�ӽ��H���Ǯ��*���-����䘗������  �  ]n=m=E�=�M=P�=r�=[+=�� =Bh == =�G�<C��<��<���<-�<8d�<n��<���<��<�6�<�h�<���<��<B��< $�<�O�<gy�<̡�<���<���<��<}2�<.R�<�o�<���<>��<���<���<���<_��<j�<��<��<��<J!�<�!�<6�<��<�<#�<���<o��<q��<��<Ֆ�<v�<�Q�<B)�<��<���<��<�`�<�$�<b��<��<PW�<�
�<���<;d�<�
�<���<�J�<���<hz�<��<#��<T"�<x��<�(�<˥�<�<���<@�<Mt�<�ޮ<�E�<.��<W	�<5f�<���<��<�j�<t��<�	�<=U�<F��<��<A)�<nk�<v��<��<�%�<L`�<!��<xЌ<^�<�:�<^n�<���<҃<��<C2�<��|<�y<|u<��q<3n<�j<�f<YDc<"�_<��[<�YX<2�T<�Q</yM<G�I<?AF<y�B<?<&~;<P�7<�_4<��0<�M-<��)<%K&<��"<(Y<��<�y<4<+�<�P<��
<��<�Z<�<{��;�:�;z��;#��;x;�;M�;U��;���;���;ļ�;�ҽ;M��;O0�;x�;�Ц;j:�;+��;A�;|ސ;݌�;�L�;��;��w;��m;=�c;�Z;�dP;r�F;;_=;*4;��*;B�!;��;��;G;�X�:H\�:ė�:>	�:8��:���:��:�Ԋ:хv:N�W:�K9:O2:u��9��9䠅9��978,I��k�;��s���̹k�� ����7�*R�n�l�r��.~���s���T��;"��	�ú��кݺj�麔���@��n����h���������%��,��2�88��>�0D�'J��
P��V���[���a��g���m�*�s�׬y�P���ł�ܽ�����Ү������������И�������  �  `n=g=E�=�M=T�=|�=X+=�� =?h =? =�G�<G��<��<���<-�<6d�<}��<���<��<�6�<�h�<���<��<\��<$�<O�<hy�<���<���<���<��<}2�<2R�<�o�<���<@��<���<���<���<i��<i�<��<��<��<K!�<�!�<O�<��<�<(�<���<x��<l��<���<Ӗ�<v�<�Q�<>)�<!��<���<���<�`�<�$�<b��<���<kW�<~
�<���<4d�<�
�<���<�J�<���<`z�<��<��<V"�<v��<�(�<ϥ�<�<���<<�<Pt�<�ޮ<�E�<)��<P	�<Of�<���<��<�j�<{��<�	�<<U�<V��<��<G)�<jk�<~��<��<�%�<P`�<��<|Ќ<X�< ;�<nn�<���<҃<��<H2�<��|<�y</|u<��q<3n<�j<�f<BDc<�_<��[<�YX<C�T<�Q<;yM<.�I<AAF<\�B<?<Q~;<C�7<�_4<��0<�M-<��)<-K&<��"<!Y<��<�y<R<+�<�P<��
<��<�Z<�<��;�:�;W��;#��;K;�;f�;E��;���;���;Լ�;�ҽ;5��;W0�;�w�;�Ц;J:�;R��;A�;fސ;݌�;�L�;��;,�w;��m;��c;�Z;�dP;{�F;}_=;�4;N�*;6�!;k�;��;�F;VY�:
\�:G��:�	�:���:ʊ�:���:�֊:�v:��W:�J9:�1:��9E�9���9��9�;8�M��o�;�It����̹ۏ����C�7��*R��l��r��a~���s���T��� ���ú~�к�ݺ���m���@�Cn���9�����\����%�:,��2�c8��>�[D��J�s
P�V�{�[�7�a���g�	�m��s���y�`���ł�	������ ���������ܜ������ϕ���  �  `n=k=H�=�M=L�=x�=_+=�� =Dh => =�G�<E��<��<���<-�<6d�<p��<���<��<�6�<�h�<���<#��<M��<$�<�O�<uy�<š�<���<���<��<�2�<'R�<�o�<���<>��<���<���<���<c��<o�<��<��<��<J!�<�!�<9�<��<
�<�<���<l��<m��<��<Ԗ�<v�<�Q�<A)�<��<���<��<�`�<�$�<h��<���<VW�<�
�<���<Ad�<�
�<���<K�<���<hz�<��<)��<T"�<x��<�(�<ƥ�<�<���<D�<Mt�<�ޮ<�E�<+��<L	�<=f�<��<��<�j�<w��<�	�<=U�<G��<��<E)�<fk�<{��<��<�%�<J`�<$��<uЌ<c�<�:�<Zn�<���<҃<��<I2�<��|<�y<%|u<��q<3n<�j<�f<cDc< �_<{�[<�YX<9�T<�Q<:yM<A�I<MAF<h�B<�?<?~;<]�7<y_4<��0<�M-<z�)<)K&<��"<Y<��<�y<7<,�<�P<��
<��<�Z<<���;�:�;b��;Y��;[;�;Z�;a��;���;Ͷ�;���;�ҽ;M��;M0�;)x�;�Ц;]:�;;��;3A�;Xސ;ڌ�;�L�;��;W�w;��m;��c;Z;�dP;��F;#_=;4;�*;=�!;H�;��;�F;�X�:!\�:}��:�	�:��: ��:嗚:,Պ:r�v:�W:fL9:�1:���9�9�9��948�C��t�;��s��?�̹�����[�7��)R�f�l��r���}���s��*U���!��\�úq�к�ݺ<��<���@��n����G����u����%�T,�2�"8��>�D��J�P��V�v�[���a���g���m��s���y�b���ł�ǽ������������$���朔�Ø�������  �  \n=l=A�=�M=R�=u�=\+=�� =Gh =; =�G�<>��<��<���<�,�<;d�<l��<���<��<�6�<�h�<���< ��<D��<,$�<�O�<dy�<š�<���<���<��<�2�<(R�<�o�<���<8��<���<���<���<]��<x�<��<��<��<=!�<�!�<8�<��<�<�< ��<f��<u��<��<ۖ�<v�<�Q�<H)�<��<��<��<�`�<�$�<_��<��<PW�<�
�<w��<:d�<�
�<���<	K�<���<pz�<��<-��<Q"�<y��<�(�<ť�<�<���<N�<Ht�<�ޮ<�E�<&��<e	�<4f�<��<��<�j�<}��<�	�<?U�<C��<��<9)�<jk�<{��<��<�%�<E`�<+��<mЌ<\�<�:�<bn�<���<҃<��<@2�<��|<�y<|u<��q<�2n<�j<�f<hDc<�_<��[<�YX<;�T<Q<*yM<A�I</AF<}�B<?<2~;<S�7<f_4<��0<�M-<��)<K&<��"<&Y<��<�y<0<,�<�P<��
<��<�Z<<���;�:�;`��;��;\;�;>�;���;���;ݶ�;���;�ҽ;S��;40�;<x�;�Ц;�:�;��;SA�;fސ;Ɍ�;�L�;r�; x;��m;�c;�Z;gdP;��F;�^=;C4;��*;m�!;:�;��;3G;X�:�\�:.��:�	�:寺:���:���:�Ԋ:��v:��W:|K9:�1:���9-�92��9��9g&8�?���;��s��V�̹5��ģ�
�7�R(R��l�zr��N~��!t���S��B"����ú$�к�ݺ��.���@��n�ȕ������r��F�%�!,�62��8�>�AD�J��
P�QV���[���a�4�g���m���s�Ԭy�.���ł�����=�������������휔����������  �  an=n=D�=�M=N�=|�=\+=�� =Bh =; =�G�<;��<��<���<-�<9d�<s��<���<��<�6�<�h�<���<#��<S��<$�<|O�<jy�<͡�<���<���<��<~2�<2R�<�o�<���<B��<���<���<���<]��<q�<��<��<��<E!�<�!�<?�<��<�<!�<���<m��<o��<��<ז�<v�<�Q�<D)�<��<���<��<�`�<�$�<^��<���<ZW�<�
�<~��<@d�<�
�<���<K�<���<jz�<��<'��<W"�<y��<�(�<ϥ�<�<���<H�<Lt�<�ޮ<�E�<%��<N	�<Bf�<
��<��<�j�<u��<�	�<6U�<I��<��<@)�<hk�<y��<��<�%�<H`�<!��<uЌ<\�<;�<`n�<���<҃<��<K2�<��|<�y<|u<��q<3n<	�j<�f<`Dc<�_<��[<�YX<C�T<�Q<>yM<I�I<>AF<]�B< ?<P~;<Q�7<w_4<��0<�M-<��)<K&<��"<"Y<��<�y<=<�<�P<��
<��<�Z<<���;�:�;H��;+��;|;�;W�;j��;���;���;Ӽ�;�ҽ;H��;]0�; x�;�Ц;s:�;��;8A�;Zސ;�;�L�;��;J�w;�m;��c;�Z;�dP;w�F;$_=;4;��*;R�!;A�;��;G;}X�:\�:���:a	�:��:���:��:qՊ:b�v:w�W:JL9:�2:���9��9⠅9V�9�58�F����;��s����̹���ʤ�N�7�&)R���l�
r���}��5t��U��o!��I�ú��к�ݺb����� A��n���m�������W�%�3,�#2�78��>�@D�xJ��
P��V���[���a���g���m��s�ݬy����ł�ӽ�����Ů����������������������  �  dn=g=I�=�M=L�=x�=X+=�� =@h =? =�G�<A��<��<���<-�<)d�<r��<���<��<�6�<�h�<���<��<S��<$�<�O�<ry�<ġ�<���<���<��<2�<7R�<�o�<���<E��<���<��<���<k��<u�<��<��<��<Y!�<�!�<=�<��<��<$�<���<u��<e��<��<Ӗ�<v�<�Q�<<)�<��<���<���<�`�<�$�<^��<��<ZW�<�
�<���<:d�<�
�<���<K�<���<iz�<��<$��<Z"�<~��<�(�<֥�<�<���<C�<Tt�<�ޮ<�E�<<��<H	�<Cf�<���<��<�j�<p��<�	�<3U�<J��<��<C)�<^k�<y��<��<�%�<Q`�<��<wЌ<V�<�:�<\n�<���<҃<��<P2�<��|<�y<,|u<��q<3n<
�j<�f<aDc<0�_<��[<�YX<G�T<�Q<JyM<.�I<RAF<{�B<�?<@~;<A�7<x_4<��0<�M-<��)<!K&<��"<Y<��<ry<:<�<�P<��
<��<�Z<�<���;x:�;���;I��;V;�;q�;J��;���;Ķ�;��;�ҽ;Y��;f0�;x�;�Ц;o:�;Y��;FA�;fސ;茋;�L�;��;T�w;�m;a�c;�Z;�dP;4�F;e_=;�4;�*;-�!;9�;��;�F;�X�:�[�:��:��:Y��:���:3��:fՊ:�v:$�W:wK9:;2:m��9��9Z��9��9 O8kI����;�nr����̹�����7��)R���l�~r���}���r��nU��`!���ú��к�ݺ���o��9A��n�^��[��^������%�F,��2�m8��>�mD��J�P��V�=�[�@�a���g��m�߼s���y�!���ł�ѽ�����î��駎�������������ϕ���  �  cn=j=>�=�M=S�=x�=^+=�� =Bh =9 =�G�<?��<��<���<-�<4d�<t��<���<��<�6�<�h�<���<��<P��<"$�<~O�<^y�<ǡ�<���<���<��<�2�</R�<�o�<���<A��<���<���<���<f��<n�<��<��<��<?!�<�!�<B�<��<
�<#�<���<i��<l��<��<і�<v�<�Q�<=)�<��<���<��<�`�<�$�<e��<���<]W�<�
�<x��<3d�<�
�<���<�J�<���<lz�<��<'��<\"�<���<�(�<ͥ�<�<���<C�<Ot�<�ޮ<�E�<$��<Y	�<Af�<��<��<�j�<p��<�	�<:U�<L��<��<A)�<fk�<z��<��<�%�<D`�<��<pЌ<b�<�:�<gn�<���<҃<��<O2�<��|<�y<5|u<��q<�2n<�j<�f<hDc<�_<��[<�YX<=�T<�Q<EyM<;�I<#AF<r�B<?<=~;<Y�7<j_4<��0<�M-<z�)<K&<��"<Y<��<�y<><!�<�P<��
<��<�Z<�<���;�:�;O��;���;d;�;b�;[��;���;��;ļ�;�ҽ;i��;U0�;x�;�Ц;t:�;E��;,A�;mސ;茋;�L�;w�;��w;*�m;��c;�Z;�dP;X�F;_=;�4;��*;"�!;B�;��;�F;�X�:\�:_��:	�:b��:ꊪ:���:�Պ:օv:��W:�J9:12:���9q�9_��9C�9�18%F����;��q����̹M����ހ7��)R�1�l�er���~��Jt��`T��~!����ú׃кDݺ�����A��n���i����}��%�%�S,�C2�K8��>�D��J��
P��V��[��a���g���m��s�{�y�#���ł�Ƚ���������������Ĝ�����������  �  ^n=t=F�=�M=P�=r�=^+=�� =Fh =7 =�G�<9��<���<���<�,�<5d�<g��<���<��<�6�<�h�<���<&��<<��<"$�<|O�<uy�<ա�<���<���<��<�2�<4R�<�o�<���<H��<���<���<���<^��<p�<��<��<��<C!�<�!�<3�<��<�<�<���<^��<q��<��<ϖ�<v�<�Q�<>)�<	��<���<���<�`�<�$�<`��<���<JW�<�
�<{��<Ld�<�
�< ��<K�<���<uz�<��<+��<^"�<���<�(�<Х�<�<���<L�<Lt�<�ޮ<�E�<%��<Y	�<,f�<
��<��<�j�<s��<�	�<7U�<?��<��<7)�<fk�<s��<��<�%�<<`�<)��<iЌ<a�<�:�<^n�<���<҃<��<C2�<��|<�y<#|u<��q<�2n<�j<$�f<pDc<�_<��[<�YX<8�T<Q<1yM<b�I<EAF<j�B<?<'~;<[�7<`_4<��0<�M-<�)<K&<��"<Y<��<�y<%<�<�P<��
<��<�Z<<_��;�:�;H��;U��;�;�;A�;���;���;߶�;ۼ�;�ҽ;l��;s0�;3x�;�Ц;�:�;$��;3A�;�ސ;֌�;�L�;��;��w;��m;y�c;�Z;WdP;��F;�^=; 4;��*;�!;;�;��;�F;�W�:1\�:���:�	�:ϯ�:���:���:jԊ:��v:�W:�M9:v2:���9��9V��9��9N28�B����;��q����̹Տ����܁7��(R���l��q��M}��?t��cT���"��M�ú�к�ݺ���]��A�o�����������l�%�3,��2��8�!>�D�J��
P��V���[�l�a��g���m��s�ìy����ł����������������ꡑ�㜔�Ę�������  �  `n=e=F�=�M=R�=y�=^+=�� =Bh =; =�G�<=��< ��<���<-�</d�<n��<���<��<�6�<�h�<���<%��<O��<"$�<�O�<my�<���<���<���< �<�2�<8R�<�o�<���<I��<���<���<���<j��<t�<��<��<��<H!�<�!�<C�<��<
�<!�<���<g��<p��<��<і�<v�<�Q�<<)�<��<���<��<�`�<�$�<g��<���<[W�<�
�<���<8d�<�
�<��<K�<���<jz�<��<"��<_"�<~��<�(�<ե�<�<���<E�<Tt�<�ޮ<�E�<+��<W	�<@f�<��<��<�j�<r��<�	�<9U�<G��<��<C)�<bk�<x��<��<�%�<F`�<"��<sЌ<a�<�:�<fn�<���<҃<��<E2�<��|<�y<*|u<��q<3n<��j<$�f<VDc<-�_<��[<�YX<N�T<�Q<;yM<(�I<CAF<k�B<?<C~;<Z�7<q_4<��0<�M-<��)<K&<��"<Y<��<~y<2<!�<�P<��
<��<�Z<
<���;�:�;Z��;4��;6;�;h�;^��;���;ʶ�;��;�ҽ;M��;x0�;x�;�Ц;j:�;T��;EA�;�ސ;���;�L�;��;~�w;/�m;��c;�Z;�dP;|�F;�^=;4;��*;!�!;B�;��;�F;PX�:(\�:T��:n	�:%��:��:Ǘ�:�Պ:&�v:�W:*K9:1:���9��9֣�91�9dD8�K��a�;�xr���̹B�����S�7��)R���l�
s��~���s���T���!��n�ú��к�ݺ������
A��n�8��Z��@�����D�%�2,�-2�38��>�D��J��
P��V���[�A�a�
�g���m�¼s���y�"���ł�轅�����ڮ��������圔����������  �  >m==��=L=H�=5�=�(=9� =Ae = =�@�<�z�<���<Z��<�#�<�Z�<5��<���<z��<�*�<=\�<c��<0��<���<��<�?�<�h�<e��<r��<���<j��<�<=�< Z�<�t�<�<Z��<˸�<���<���<���<P��<U��<���<$�<��<w��<��<���<���<���<���<��<���<�o�<lN�<M)�<n �<���< ��<�n�<6�<���<��<Gt�<�+�<���<j��<!8�<���<���<&�<8��<	O�<��<�n�<:��<�}�<���<X}�<@��<�m�<�߱<�N�<��<�!�<M��<o�<eE�<$��<���<�L�<՞�<8�<�:�<��<�̚<q�<�U�<��<c֓<��<�O�<���<H<h��<G/�<�c�<{��<'ʃ<���<�,�<[�|<y<�xu<��q<�4n<P�j<��f<�Mc<��_<�
\<�jX<��T<�-Q<��M<�I<�^F<$�B<W4?<�;<�8<2�4<� 1<}|-<��)<�~&<�#<F�<v!<c�<oP<��<O�<�><��<Ϥ<a<�G�;���;�z�;�)�;���;��;���;~t�;�l�;cu�;���;0��;�;+8�;I��;���;lx�;��;T��;�P�;��;�;؄y;>jo;pe;ܗ[;��Q;�IH;��>;*}5;UF,;�.#;F5;1Z;��;���:���:�:���:>�:7�:I�:��:��z:n\:�v=:?:\:ѓ�9��9	7&9�N8��x�ͯ.�N ��Bjƹ(;�������4��O�j��9���P��zS���?��t��{�º��Ϻ�1ܺ'���C���� �k��:��`������̱%���+���1���7���=�P�C���I�\�O�~�U���[���a�i�g�7�m�p�s�֘y�݋�@��� �������l���T���4���ɠ��5���2����  �  >m==��=L=E�=/�=�(=7� =He =� =�@�<�z�< ��<g��<�#�<�Z�<9��<���<l��<�*�<D\�<\��<5��<���<��<�?�<�h�<h��<w��<���<j��<*�<=�<�Y�<�t�<���<X��<¸�<���<���<���<_��<V��<���<%�<��<h��<��<���<���<���<���<��<���<�o�<wN�<W)�<v �<���<"��<�n�<6�<���<���<Ht�<|+�<���<l��<!8�<���<��<0�<7��<O�<��<�n�<&��<�}�<���<R}�<J��<�m�<�߱<�N�<��<�!�<Q��<v�<WE�<(��<���<�L�<֞�<&�<�:�<!��<�̚<{�<�U�<��<i֓<��<�O�<���<A<g��<A/�<�c�<���<$ʃ<���<�,�<~�|< y<�xu<	�q<�4n<J�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<��M<�I<�^F<9�B<L4?<��;<�8<)�4<1<]|-<��)<�~&<�#<`�<�!<�<xP<��<4�<z><��<��<#a<�G�;���;{�;o)�;���;-��;1��;|t�;m�;]u�;���; ��;��;%8�;%��;���;wx�;��;���;�P�;��;!�;@�y;�io;�oe;��[;d�Q;�IH;H�>;"}5;qF,;�.#;�5;�Z;�;��:��:�:��:6�:��:T�:�:D�z:�\:�v=:$?:�]:.��9~�9�<&95N8��x�	�.��#���jƹ�<�������4�`�O�j��9��DQ��6S��l?��M��=�º*�Ϻ�1ܺ��E���� �M�k:�]`���������%��+�a�1��7���=�V�C���I���O��U���[���a�a�g���m�b�s���y����\������$���z���d����������5���󜚻�  �  ;m==��=L=D�=2�=�(=0� =Je =� =�@�<�z�<���<c��<�#�<�Z�<1��<���<w��<�*�<D\�<R��<A��<���<��<�?�<�h�<n��<r��<���<]��<-�<=�< Z�<�t�<���<h��<���<���<���<���<W��<W��<���<�<��<d��<��<���<���<���<���<��<���<�o�<pN�<N)�<n �<���<-��<�n�<%6�<���<���<Xt�<x+�<���<d��<#8�<���<���<(�<2��<O�<��<�n�<3��<�}�<���<M}�<O��<tm�<�߱<�N�<��<�!�<O��<y�<WE�<6��<���<�L�<ߞ�</�<�:�<��<�̚<q�<�U�<��<i֓<��<�O�<���<5<q��<I/�<�c�<���<ʃ<���<�,�<x�|<y<�xu<�q<�4n<k�j<��f<�Mc<�_<�
\<�jX<y�T<�-Q<��M<�I<�^F<<�B<G4?<�;<�8<�4<"1<k|-<��)<�~&<�#<Y�<x!<t�<hP<��<I�<�><��<��<;a<�G�;���;{�;V)�;���;��;&��;Ht�;m�;Ru�;���;A��;��;g8�;��;���;hx�;��;r��;�P�;��; �;Z�y;�io;ipe;ɗ[;"�Q;JH;d�>;�}5;XF,;�.#;g5;;Z;��;���:���:O�:���:��:��:M�:��:��z:�\:�v=:;?:�\:R��9*�91@&9�M8�lx�O�.�����iƹ�=�����O�4�؅O��j��9��wQ��SS��??��V��W�º��Ϻ�1ܺ��躍D���� ����:��`�΀�����%���+�/�1���7�B�=��C���I���O�"�U���[���a�o�g�±m�٥s���y����g���˸������5���m����������q��������  �  >m==��=L=F�=3�=�(=7� =Ce =� =�@�<�z�<��<e��<�#�<�Z�<;��<���<y��<�*�<@\�<_��</��<���<��<�?�<�h�<n��<v��<���<f��<$�<=�<�Y�<�t�<���<T��<ĸ�<���<���<���<X��<^��<���<�<��<o��<��<���<���<���<���<��<���<�o�<yN�<Z)�<t �<���<��<�n�<6�<���<���<Gt�<�+�<���<g��<!8�<���<��<-�<9��<O�<��<�n�<,��<�}�<���<X}�<D��<}m�<�߱<�N�<��<�!�<Q��<q�<`E�<$��<���<�L�<Ӟ�<4�<�:�<"��<�̚<~�<�U�<��<c֓<��<�O�<���<D<g��<D/�<�c�<���< ʃ<���<�,�<s�|<y<�xu<�q<�4n<D�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<��M<�I<�^F<1�B<P4?<�;<�8<,�4<1<q|-<��)<�~&<�#<^�<�!<y�<}P<��<M�<|><��<Ǥ<a<�G�;���;{�;V)�;���;(��;"��;mt�;�l�;tu�;���;��;��;8�;.��;���;yx�;��;t��;Q�;��;�;�y; jo;�oe;��[;~�Q;�IH;��>;"}5;oF,;�.#;�5;�Z;ޜ;��:���:��:���:c�:��:H�:Q�:��z:\:�v=:"@:]:���9��9_:&9�N8F�x��.�R"��Elƹ�:��K��;�4�؅O�Sj�u9��tQ��.S���?�����}�º�Ϻ�1ܺG��1D��� �G�u:�C`�������ʱ%���+���1�h�7���=�U�C���I��O�J�U���[���a�L�g�ױm�i�s�Řy����P���������x���h������Ġ��:�������  �  >m==��=L=D�=3�=�(=?� =Ce =� =�@�<�z�<��<Y��<�#�<}Z�<>��<���<y��<�*�<C\�<k��<*��<���<��<�?�<�h�<f��<v��<���<m��<�<=�<�Y�<�t�<���<Q��<ɸ�<���<���<���<V��<Y��<���<+�<��<s��<��<���<���<���<���<ݧ�<���<�o�<qN�<U)�<h �<���<��<�n�<6�<���<���<Ft�<�+�<���<r��<8�<���<��<(�<7��<O�<��<�n�<9��<�}�<���<[}�<;��<�m�<�߱<�N�<��<�!�<X��<j�<fE�<��<���<�L�<Ҟ�<7�<�:�<&��<�̚<�<�U�<��<j֓<��<�O�<���<R<c��<D/�<�c�<���<'ʃ<���<�,�<i�|<'y<�xu<��q<�4n<<�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<��M<��I<�^F<<�B<H4?<�;<}8<K�4<1<r|-<��)<�~&<�#<E�<�!<Y�<�P<��<O�<y><��<ޤ<a< H�;���;({�;^)�;���;'��;	��;�t�;�l�;vu�;���;��;�;8�;D��;���;ix�;��;o��;�P�;f�;5�;�y;jo;�oe;��[;��Q;�IH;��>; }5;�F,;�.#;r5;qZ;��;v��:���:?�:l��:��:��:9�:��:��z:v\:iu=:�?:�\:>��9y�95&9�N8�x�_�.�� ��olƹ:��a����4���O�>j��9���Q���R��+@��j����º}�Ϻ`1ܺ]���C��� �!��:�?`�
�������%�0�+���1�f�7�V�=�w�C���I���O�5�U���[��a�K�g���m�C�s��y���B���)���ʲ������a���0���Ӡ��!�������  �  ?m==��=L=B�=5�=�(=2� =Ee =  =�@�<�z�<���<e��<�#�<�Z�<9��<���<u��<�*�<B\�<W��<<��<���<��<�?�<�h�<n��<u��<���<a��<*�<	=�<�Y�<�t�<���<V��<���<���<���<���<U��<Z��<���<"�<��<d��<��<���<���<���<���<��<���<�o�<|N�<^)�<o �<���<$��<�n�<6�<���<���<Xt�<y+�<���<j��<8�<���<���<$�<5��<O�<��<�n�<0��<�}�<���<P}�<K��<xm�<�߱<�N�<��<�!�<T��<r�<[E�<1��<���<�L�<ڞ�</�<�:�<!��<�̚<��<�U�<��<j֓<��<�O�<���<9<n��<N/�<�c�<���<ʃ<���<�,�<i�|<
y<�xu<�q<�4n<H�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<��M<�I<�^F<A�B<>4?<�;<�8<�4<1<v|-<��)<�~&<�#<]�<�!<s�<wP<��<F�<�><��<��<1a<�G�;���;${�;X)�;���;#��;��;Zt�;m�;Vu�;���;��;��;8�;��;���;vx�;��;i��;Q�;��;�; �y;�io;�pe;ɗ[;J�Q;�IH;��>;V}5;sF,;�.#;�5;�Z;��;��:3��:��:��:�:��:_�:��:��z:r\:6v=:�?:�\:T��9�9)?&9��M8n�x���.��!���kƹ=��l����4���O��j�s9���Q���R���?������ºm�Ϻ�1ܺ��躋D���� �J��:�`���������%���+��1�8�7�$�=��C�m�I���O��U���[���a�9�g���m���s���y����o����������y���v���#�������`�������  �  :m==��=L=E�=.�=�(=4� =Ke =� =�@�<�z�<��<j��<�#�<�Z�<6��<���<s��<�*�<J\�<Y��<?��<���<��<�?�<�h�<p��<l��<���<U��<-�<=�<�Y�<�t�<���<_��<���<���<x��<���<\��<T��<���<�<��<^��<��<���<���<���<���<��<���<�o�<xN�<T)�<y �<���<,��<�n�<#6�<���<���<Qt�<o+�<���<Z��<#8�<���<��<1�<&��<O�<��<�n�<)��<�}�<���<K}�<N��<jm�<�߱<�N�<��<�!�<F��<}�<NE�<2��<���<�L�<ܞ�<+�<�:�<��<�̚<q�<�U�<��<i֓<��<�O�<���<<<q��<A/�<�c�<���<ʃ<���<�,�<��|<y<�xu<�q<�4n<X�j<��f<�Mc<�_<�
\<�jX<}�T<�-Q<z�M<�I<u^F<;�B<L4?<�;<�8<�4<&1<g|-<��)<�~&<�#<f�<v!<��<rP<��<C�<�><��<��<7a<�G�;���;�z�;S)�;��; ��;O��;*t�;m�;Mu�;���;��;��;B8�;���;���;Hx�;��;���;�P�;��;���;��y;xio;;pe;ؗ[;g�Q;JH;7�>;�}5;KF,;/#;�5;lZ;�;���:���:��:���:��:��:��:5�:��z:�\:�v=:S?:6]:���9j�9)?&9��M8�~x�i�.��!���iƹ'>������4�ʄO�[j�u9��uQ���S���>�������ºA�Ϻ-1ܺ��躾D���� �}�1:��`����q����%���+�Q�1���7��=��C���I���O� �U�:�[���a���g���m���s�˘y����c���񸅻-���a���e���%�������i���䜚��  �  8m==��=L=H�=1�=�(=9� =De =� =�@�<�z�<���<e��<�#�<�Z�<3��<���<{��<�*�<@\�<c��<9��<���<��<�?�<�h�<m��<h��<���<^��<*�<
=�<�Y�<�t�<���<U��<���<���<|��<���<R��<Q��<���< �<��<l��<
��<���<���<���<���<��<���<�o�<xN�<Y)�<s �<���<+��<�n�<6�<���<���<Lt�<~+�<���<f��<)8�<���<���<*�<.��<O�<��<�n�<6��<�}�<���<P}�<I��<tm�<�߱<�N�<��<�!�<I��<r�<]E�<,��<���<�L�<՞�<5�<�:�<��<�̚<}�<�U�<��<j֓<��<�O�<���<F<m��<D/�<�c�<���<"ʃ<���<�,�<n�|<y<�xu<��q<�4n<>�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<r�M<�I<�^F<*�B<W4?<��;<�8<4�4<
1<p|-<��)<�~&<�#<]�<�!<}�<mP<��<R�<�><��<Ф<,a<�G�;���;�z�;�)�;���;��;��;Nt�;m�;Yu�;���;��;�;8�;��;���;Zx�;��;`��;�P�;��;�;'�y;�io;"pe;�[;��Q;�IH;��>;p}5;tF,;�.#;�5;�Z;؜;%��:���:��:���:i�:�:��:%�:��z:�\:�w=:?:	\:Ӕ�9^�9�:&9��M8U�x�ֱ.�/!���lƹ=�����@�4��O��j��9���P���S���?�������ºǏϺ�1ܺ/��D���� �t�{:�K`���������%���+��1�C�7���=�#�C���I�j�O�W�U���[���a���g��m���s�Řy�ҋ�`���%���ᲈ�����w���2�������N�������  �  Dm=
=��=L=G�=4�=�(=9� =Ce = =�@�<�z�<��<d��< $�<�Z�<A��<���<s��<�*�<@\�<b��<-��<���<��<�?�<�h�<d��<���<���<d��<�<
=�<�Y�<�t�<���<I��<ĸ�<���<���<���<[��<^��<���<+�<��<r��<��<���<���<���<���<ڧ�<���<�o�<~N�<a)�<n �<���<��<�n�<6�<���<���<Gt�<�+�<��<r��<8�<���<��< �<9��<O�<��<{n�<-��<�}�<}��<T}�<>��<}m�<�߱<�N�<��<�!�<Y��<l�<eE�<"��<���<�L�<ߞ�<1�<�:�<+��<�̚<��<�U�<��<o֓<��<�O�<���<G<e��<G/�<�c�<}��<'ʃ<���<�,�<n�|<y<�xu<��q<�4n<%�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<��M<��I<�^F<.�B<S4?<�;<�8<2�4<1<�|-<��)<�~&<�#<[�<�!<p�<�P<��<C�<�><��<ͤ<a< H�;���;!{�;R)�;���;U��;��;ft�;�l�;\u�;���;�;��;�7�;/��;���;�x�;��;���;Q�;[�;7�;߄y;jo;pe;��[;��Q;�IH;��>;�|5;�F,;�.#;�5;�Z;��;���:r��:'�:ʁ�:��:��:K�:��:��z:�\:=u=:�?:�]:i��9"�9�6&9N80�x��.�$���mƹ<�����4��O�!j��9���Q���R��@��t����º܏Ϻ�1ܺ���eD��� ����:��_�������k�%�.�+���1�\�7���=�d�C���I�k�O�n�U���[�"�a��g��m�˥s���y����G���V���㲈�����[���<���ʠ��`�������  �  =m==��=L=D�=2�=�(=8� =Ge = =�@�<�z�<��<f��<�#�<�Z�<=��<���<w��<�*�<D\�<b��<9��<���<��<�?�<�h�<g��<s��<���<`��<#�<=�<�Y�<�t�<���<W��<���<���<���<���<U��<U��<���<%�<��<j��<��<���<���<���<���<��<���<�o�<uN�<U)�<p �<���<!��<�n�<6�<���<��<Pt�<{+�<���<l��<8�<���<���<#�<3��<O�<��<�n�<0��<�}�<���<M}�<B��<wm�<�߱<�N�<��<�!�<V��<p�<ZE�<,��<���<�L�<ޞ�<5�<�:�<&��<�̚<y�<�U�<��<q֓<��<�O�<���<F<n��<C/�<�c�<���<#ʃ<���<�,�<j�|<y<�xu<��q<�4n<E�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<��M<�I<�^F<;�B<H4?<��;<�8</�4<1<�|-<��)<�~&<�#<`�<�!<y�<�P<��<J�<�><��<Τ<,a<�G�;���;!{�;R)�;���;��;��;Yt�;�l�;Bu�;���;��;��;%8�;��;���;sx�;��;j��;�P�;k�;!�;�y;�io;=pe;�[;��Q;�IH;��>;3}5;�F,;�.#;�5;rZ;��;���:��:.�::��:��:6�:��: �:��z:�\:Yu=:�>:�\:+��9��98&9�M8��x���.��!���kƹ�=��u����4��O��j��9���Q���R���?������º��Ϻ�1ܺ���"D���� �'��:�l`�������]�%���+���1�'�7���=��C���I���O�&�U���[��a�^�g���m�ås���y���P����������w���a���S�������]�������  �  6m==��=L=F�=1�=�(=6� =Ge =� =�@�<�z�<��<u��<�#�<�Z�<5��<���<x��<�*�<F\�<^��<<��<���<��<�?�<�h�<p��<d��<���<Z��<.�<	=�<�Y�<�t�<���<R��<���<���<{��<���<S��<N��<���<�<��<g��<��<���<���<���<���<��<���<�o�<�N�<^)�<� �<���<-��<�n�<6�<���<���<Qt�<x+�<���<d��<(8�<���<���<2�<+��<O�<��<�n�<#��<�}�<}��<M}�<O��<om�<�߱<�N�<��<�!�<J��<x�<YE�</��<���<�L�<Ӟ�<2�<�:�<��<͚<|�<�U�<��<j֓<��<�O�<���<B<n��<B/�<�c�<���<ʃ<���<�,�<w�|<y<�xu<�q<�4n<A�j<��f<�Mc<ԫ_<�
\<�jX<��T<�-Q<l�M<�I<�^F<6�B<P4?<��;<�8<%�4<1<h|-<��)<�~&<�#<~�<�!<��<qP<��<M�<z><��<Ƥ<1a<�G�;���;�z�;x)�;��;��;I��;?t�; m�;Vu�;���;��;��;8�;���;���;Vx�;��;e��;�P�;��;���;X�y;�io;;pe;͗[;z�Q;�IH;��>;�}5;aF,;/#;�5;�Z;K�;��:���:��:���:S�:��:��:��:��z:�\:�w=:�>:�[:��9��9�?&9��M8��x�Ժ.��#���mƹ�=�������4�ׄO�\j�}9��Q���S��F?��3����º��Ϻp1ܺK��LD��|� �i��9�P`�J��n����%���+��1��7���=��C���I���O��U� �[�x�a�ƽg�űm���s���y����������,�����������(�������c�����  �  =m==��=L=F�=4�=�(=9� =Ie = =�@�<�z�<��<d��<�#�<�Z�<:��<���<{��<�*�<J\�<^��<4��<���<��<�?�<�h�<g��<p��<���<U��<!�<=�<�Y�<�t�<���<X��<���<���<s��<���<U��<U��<���<�<��<k��<��<���<���<���<���<��<���<�o�<qN�<P)�<u �<���<&��<�n�< 6�<���<���<Pt�<+�<���<g��<8�<���<���<)�<%��<O�<��<�n�<-��<�}�<���<O}�<B��<lm�<�߱<�N�<��<�!�<O��<u�<`E�<)��<���<�L�<���<5�<�:�<#��<�̚<p�<�U�<��<l֓<��<�O�<���<H<g��<J/�<�c�<���<ʃ<���<�,�<s�|<y<�xu<��q<�4n<K�j<��f<�Mc<�_<�
\<�jX<s�T<�-Q<��M<�I<}^F<8�B<N4?<�;<�8<2�4<1<�|-<��)<�~&<�#<[�<y!<�<zP<��<R�<�><��<Ƥ<"a<�G�;���;{�;N)�;���;��;1��;+t�;�l�;Tu�;���;��;��;)8�;��;���;6x�;��;j��;�P�;{�;�;B�y;�io;Ipe;��[;��Q;�IH;��>;`}5;�F,;�.#;v5;NZ;�;i��:b��:�:X��:��:��:��:6�::�z:9\:�u=:)?:]\:���9#�9�9&9��M8.�x�.�.��!��kƹ+=�����?�4�~�O�2j��9���Q��ES��p?������º�Ϻ1ܺs��D���� �7�l:��`�΀�x����%���+���1��7���=�W�C���I���O�'�U��[���a�p�g�Աm�ڥs��y�ԋ�^���
������q���n���/���ޠ��~��������  �  >m==��=L=A�=7�=�(=8� =Ae = =�@�<�z�<��<i��<$�<�Z�<B��<���<t��<�*�<9\�<]��<6��<���<��<�?�<�h�<j��<w��<���<e��<(�<=�<�Y�<�t�<���<P��<���<���<���<���<P��<^��<���<,�<��<g��<��<���<���<���<���<ާ�<���<�o�<N�<b)�<u �<���<��<�n�<6�<���<���<Qt�<|+�<���<u��<8�<���<���<"�<7��<O�<��<�n�<#��<�}�<���<J}�<D��<}m�<�߱<�N�<��<�!�<]��<h�<`E�<+��<���<�L�<ڞ�<1�<�:�<-��<�̚<��<�U�<!��<k֓<��<�O�<���<D<d��<P/�<�c�<���<'ʃ<���<�,�<b�|<y<�xu<��q<�4n</�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<��M< �I<�^F<@�B<:4?<�;<�8<0�4<� 1<�|-<��)<�~&<�#<e�<�!<��<�P<��<D�<�><��<ä<&a<�G�;���;7{�;^)�;���;/��;���;kt�;m�;=u�;���;ᵸ;��;8�;��;���;�x�;��;W��;Q�;m�;=�;��y;�io;npe;��[;_�Q;�IH;��>;	}5;�F,;�.#;�5;�Z;�;���:���:=�:���:�:��:��:�:��z:�\:Wu=:.@:.\:��9��9�8&97�M8$�x��.�7%���lƹD>��5��(�4�;�O��j��9���Q��pR��8@����� �º"�Ϻ2ܺ���dD���� ���X:��_����c����%��+���1���7���=�l�C�_�I���O�$�U���[���a�C�g��m���s���y���l���B���-�������v���I�������@���/����  �  =m==��=L=F�=4�=�(=9� =Ie = =�@�<�z�<��<d��<�#�<�Z�<:��<���<{��<�*�<J\�<^��<4��<���<��<�?�<�h�<g��<p��<���<U��<!�<=�<�Y�<�t�<���<X��<���<���<s��<���<U��<U��<���<�<��<k��<��<���<���<���<���<��<���<�o�<qN�<P)�<u �<���<&��<�n�< 6�<���<���<Pt�<+�<���<g��<8�<���<���<)�<%��<O�<��<�n�<-��<�}�<���<O}�<B��<lm�<�߱<�N�<��<�!�<O��<u�<`E�<)��<���<�L�<���<5�<�:�<#��<�̚<p�<�U�<��<l֓<��<�O�<���<H<g��<J/�<�c�<���<ʃ<���<�,�<s�|<y<�xu<��q<�4n<K�j<��f<�Mc<�_<�
\<�jX<s�T<�-Q<��M<�I<}^F<8�B<N4?<�;<�8<2�4<1<�|-<��)<�~&<�#<[�<y!<�<zP<��<R�<�><��<Ƥ<"a<�G�;���;{�;N)�;���;��;1��;+t�;�l�;Tu�;���;��;��;)8�;��;���;6x�;��;j��;�P�;{�;�;B�y;�io;Ipe;��[;��Q;�IH;��>;`}5;�F,;�.#;v5;NZ;�;i��:b��:�:X��:��:��:��:6�::�z:9\:�u=:)?:]\:���9#�9�9&9��M8.�x�.�.��!��kƹ+=�����?�4�~�O�2j��9���Q��ES��p?������º�Ϻ1ܺs��D���� �7�l:��`�΀�x����%���+���1��7���=�W�C���I���O�'�U��[���a�p�g�Աm�ڥs��y�ԋ�^���
������q���n���/���ޠ��~��������  �  6m==��=L=F�=1�=�(=6� =Ge =� =�@�<�z�<��<u��<�#�<�Z�<5��<���<x��<�*�<F\�<^��<<��<���<��<�?�<�h�<p��<d��<���<Z��<.�<	=�<�Y�<�t�<���<R��<���<���<{��<���<S��<N��<���<�<��<g��<��<���<���<���<���<��<���<�o�<�N�<^)�<� �<���<-��<�n�<6�<���<���<Qt�<x+�<���<d��<(8�<���<���<2�<+��<O�<��<�n�<#��<�}�<}��<M}�<O��<om�<�߱<�N�<��<�!�<J��<x�<YE�</��<���<�L�<Ӟ�<2�<�:�<��<͚<|�<�U�<��<j֓<��<�O�<���<B<n��<B/�<�c�<���<ʃ<���<�,�<w�|<y<�xu<�q<�4n<A�j<��f<�Mc<ԫ_<�
\<�jX<��T<�-Q<l�M<�I<�^F<6�B<P4?<��;<�8<%�4<1<h|-<��)<�~&<�#<~�<�!<��<qP<��<M�<z><��<Ƥ<1a<�G�;���;�z�;x)�;��;��;I��;?t�; m�;Vu�;���;��;��;8�;���;���;Vx�;��;e��;�P�;��;���;X�y;�io;;pe;͗[;z�Q;�IH;��>;�}5;aF,;/#;�5;�Z;K�;��:���:��:���:S�:��:��:��:��z:�\:�w=:�>:�[:��9��9�?&9��M8��x�Ժ.��#���mƹ�=�������4�ׄO�\j�}9��Q���S��F?��3����º��Ϻp1ܺK��LD��|� �i��9�P`�J��n����%���+��1��7���=��C���I���O��U� �[�x�a�ƽg�űm���s���y����������,�����������(�������c�����  �  =m==��=L=D�=2�=�(=8� =Ge = =�@�<�z�<��<f��<�#�<�Z�<=��<���<w��<�*�<D\�<b��<9��<���<��<�?�<�h�<g��<s��<���<`��<#�<=�<�Y�<�t�<���<W��<���<���<���<���<U��<U��<���<%�<��<j��<��<���<���<���<���<��<���<�o�<uN�<U)�<p �<���<!��<�n�<6�<���<��<Pt�<{+�<���<l��<8�<���<���<#�<3��<O�<��<�n�<0��<�}�<���<M}�<B��<wm�<�߱<�N�<��<�!�<V��<p�<ZE�<,��<���<�L�<ޞ�<5�<�:�<&��<�̚<y�<�U�<��<q֓<��<�O�<���<F<n��<C/�<�c�<���<#ʃ<���<�,�<j�|<y<�xu<��q<�4n<E�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<��M<�I<�^F<;�B<H4?<��;<�8</�4<1<�|-<��)<�~&<�#<`�<�!<y�<�P<��<J�<�><��<Τ<,a<�G�;���;!{�;R)�;���;��;��;Yt�;�l�;Bu�;���;��;��;%8�;��;���;sx�;��;j��;�P�;k�;!�;�y;�io;=pe;�[;��Q;�IH;��>;3}5;�F,;�.#;�5;rZ;��;���:��:.�::��:��:6�:��: �:��z:�\:Yu=:�>:�\:+��9��98&9�M8��x���.��!���kƹ�=��u����4��O��j��9���Q���R���?������º��Ϻ�1ܺ���"D���� �'��:�l`�������]�%���+���1�'�7���=��C���I���O�&�U���[��a�^�g���m�ås���y���P����������w���a���S�������]�������  �  Dm=
=��=L=G�=4�=�(=9� =Ce = =�@�<�z�<��<d��< $�<�Z�<A��<���<s��<�*�<@\�<b��<-��<���<��<�?�<�h�<d��<���<���<d��<�<
=�<�Y�<�t�<���<I��<ĸ�<���<���<���<[��<^��<���<+�<��<r��<��<���<���<���<���<ڧ�<���<�o�<~N�<a)�<n �<���<��<�n�<6�<���<���<Gt�<�+�<��<r��<8�<���<��< �<9��<O�<��<{n�<-��<�}�<}��<T}�<>��<}m�<�߱<�N�<��<�!�<Y��<l�<eE�<"��<���<�L�<ߞ�<1�<�:�<+��<�̚<��<�U�<��<o֓<��<�O�<���<G<e��<G/�<�c�<}��<'ʃ<���<�,�<n�|<y<�xu<��q<�4n<%�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<��M<��I<�^F<.�B<S4?<�;<�8<2�4<1<�|-<��)<�~&<�#<[�<�!<p�<�P<��<C�<�><��<ͤ<a< H�;���;!{�;R)�;���;U��;��;ft�;�l�;\u�;���;�;��;�7�;/��;���;�x�;��;���;Q�;[�;7�;߄y;jo;pe;��[;��Q;�IH;��>;�|5;�F,;�.#;�5;�Z;��;���:r��:'�:ʁ�:��:��:K�:��:��z:�\:=u=:�?:�]:i��9"�9�6&9N80�x��.�$���mƹ<�����4��O�!j��9���Q���R��@��t����º܏Ϻ�1ܺ���eD��� ����:��_�������k�%�.�+���1�\�7���=�d�C���I�k�O�n�U���[�"�a��g��m�˥s���y����G���V���㲈�����[���<���ʠ��`�������  �  8m==��=L=H�=1�=�(=9� =De =� =�@�<�z�<���<e��<�#�<�Z�<3��<���<{��<�*�<@\�<c��<9��<���<��<�?�<�h�<m��<h��<���<^��<*�<
=�<�Y�<�t�<���<U��<���<���<|��<���<R��<Q��<���< �<��<l��<
��<���<���<���<���<��<���<�o�<xN�<Y)�<s �<���<+��<�n�<6�<���<���<Lt�<~+�<���<f��<)8�<���<���<*�<.��<O�<��<�n�<6��<�}�<���<P}�<I��<tm�<�߱<�N�<��<�!�<I��<r�<]E�<,��<���<�L�<՞�<5�<�:�<��<�̚<}�<�U�<��<j֓<��<�O�<���<F<m��<D/�<�c�<���<"ʃ<���<�,�<n�|<y<�xu<��q<�4n<>�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<r�M<�I<�^F<*�B<W4?<��;<�8<4�4<
1<p|-<��)<�~&<�#<]�<�!<}�<mP<��<R�<�><��<Ф<,a<�G�;���;�z�;�)�;���;��;��;Nt�;m�;Yu�;���;��;�;8�;��;���;Zx�;��;`��;�P�;��;�;'�y;�io;"pe;�[;��Q;�IH;��>;p}5;tF,;�.#;�5;�Z;؜;%��:���:��:���:i�:�:��:%�:��z:�\:�w=:?:	\:Ӕ�9^�9�:&9��M8U�x�ֱ.�/!���lƹ=�����@�4��O��j��9���P���S���?�������ºǏϺ�1ܺ/��D���� �t�{:�K`���������%���+��1�C�7���=�#�C���I�j�O�W�U���[���a���g��m���s�Řy�ҋ�`���%���ᲈ�����w���2�������N�������  �  :m==��=L=E�=.�=�(=4� =Ke =� =�@�<�z�<��<j��<�#�<�Z�<6��<���<s��<�*�<J\�<Y��<?��<���<��<�?�<�h�<p��<l��<���<U��<-�<=�<�Y�<�t�<���<_��<���<���<x��<���<\��<T��<���<�<��<^��<��<���<���<���<���<��<���<�o�<xN�<T)�<y �<���<,��<�n�<#6�<���<���<Qt�<o+�<���<Z��<#8�<���<��<1�<&��<O�<��<�n�<)��<�}�<���<K}�<N��<jm�<�߱<�N�<��<�!�<F��<}�<NE�<2��<���<�L�<ܞ�<+�<�:�<��<�̚<q�<�U�<��<i֓<��<�O�<���<<<q��<A/�<�c�<���<ʃ<���<�,�<��|<y<�xu<�q<�4n<X�j<��f<�Mc<�_<�
\<�jX<}�T<�-Q<z�M<�I<u^F<;�B<L4?<�;<�8<�4<&1<g|-<��)<�~&<�#<f�<v!<��<rP<��<C�<�><��<��<7a<�G�;���;�z�;S)�;��; ��;O��;*t�;m�;Mu�;���;��;��;B8�;���;���;Hx�;��;���;�P�;��;���;��y;xio;;pe;ؗ[;g�Q;JH;7�>;�}5;KF,;/#;�5;lZ;�;���:���:��:���:��:��:��:5�:��z:�\:�v=:S?:6]:���9j�9)?&9��M8�~x�i�.��!���iƹ'>������4�ʄO�[j�u9��uQ���S���>�������ºA�Ϻ-1ܺ��躾D���� �}�1:��`����q����%���+�Q�1���7��=��C���I���O� �U�:�[���a���g���m���s�˘y����c���񸅻-���a���e���%�������i���䜚��  �  ?m==��=L=B�=5�=�(=2� =Ee =  =�@�<�z�<���<e��<�#�<�Z�<9��<���<u��<�*�<B\�<W��<<��<���<��<�?�<�h�<n��<u��<���<a��<*�<	=�<�Y�<�t�<���<V��<���<���<���<���<U��<Z��<���<"�<��<d��<��<���<���<���<���<��<���<�o�<|N�<^)�<o �<���<$��<�n�<6�<���<���<Xt�<y+�<���<j��<8�<���<���<$�<5��<O�<��<�n�<0��<�}�<���<P}�<K��<xm�<�߱<�N�<��<�!�<T��<r�<[E�<1��<���<�L�<ڞ�</�<�:�<!��<�̚<��<�U�<��<j֓<��<�O�<���<9<n��<N/�<�c�<���<ʃ<���<�,�<i�|<
y<�xu<�q<�4n<H�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<��M<�I<�^F<A�B<>4?<�;<�8<�4<1<v|-<��)<�~&<�#<]�<�!<s�<wP<��<F�<�><��<��<1a<�G�;���;${�;X)�;���;#��;��;Zt�;m�;Vu�;���;��;��;8�;��;���;vx�;��;i��;Q�;��;�; �y;�io;�pe;ɗ[;J�Q;�IH;��>;V}5;sF,;�.#;�5;�Z;��;��:3��:��:��:�:��:_�:��:��z:r\:6v=:�?:�\:T��9�9)?&9��M8n�x���.��!���kƹ=��l����4���O��j�s9���Q���R���?������ºm�Ϻ�1ܺ��躋D���� �J��:�`���������%���+��1�8�7�$�=��C�m�I���O��U���[���a�9�g���m���s���y����o����������y���v���#�������`�������  �  >m==��=L=D�=3�=�(=?� =Ce =� =�@�<�z�<��<Y��<�#�<}Z�<>��<���<y��<�*�<C\�<k��<*��<���<��<�?�<�h�<f��<v��<���<m��<�<=�<�Y�<�t�<���<Q��<ɸ�<���<���<���<V��<Y��<���<+�<��<s��<��<���<���<���<���<ݧ�<���<�o�<qN�<U)�<h �<���<��<�n�<6�<���<���<Ft�<�+�<���<r��<8�<���<��<(�<7��<O�<��<�n�<9��<�}�<���<[}�<;��<�m�<�߱<�N�<��<�!�<X��<j�<fE�<��<���<�L�<Ҟ�<7�<�:�<&��<�̚<�<�U�<��<j֓<��<�O�<���<R<c��<D/�<�c�<���<'ʃ<���<�,�<i�|<'y<�xu<��q<�4n<<�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<��M<��I<�^F<<�B<H4?<�;<}8<K�4<1<r|-<��)<�~&<�#<E�<�!<Y�<�P<��<O�<y><��<ޤ<a< H�;���;({�;^)�;���;'��;	��;�t�;�l�;vu�;���;��;�;8�;D��;���;ix�;��;o��;�P�;f�;5�;�y;jo;�oe;��[;��Q;�IH;��>; }5;�F,;�.#;r5;qZ;��;v��:���:?�:l��:��:��:9�:��:��z:v\:iu=:�?:�\:>��9y�95&9�N8�x�_�.�� ��olƹ:��a����4���O�>j��9���Q���R��+@��j����º}�Ϻ`1ܺ]���C��� �!��:�?`�
�������%�0�+���1�f�7�V�=�w�C���I���O�5�U���[��a�K�g���m�C�s��y���B���)���ʲ������a���0���Ӡ��!�������  �  >m==��=L=F�=3�=�(=7� =Ce =� =�@�<�z�<��<e��<�#�<�Z�<;��<���<y��<�*�<@\�<_��</��<���<��<�?�<�h�<n��<v��<���<f��<$�<=�<�Y�<�t�<���<T��<ĸ�<���<���<���<X��<^��<���<�<��<o��<��<���<���<���<���<��<���<�o�<yN�<Z)�<t �<���<��<�n�<6�<���<���<Gt�<�+�<���<g��<!8�<���<��<-�<9��<O�<��<�n�<,��<�}�<���<X}�<D��<}m�<�߱<�N�<��<�!�<Q��<q�<`E�<$��<���<�L�<Ӟ�<4�<�:�<"��<�̚<~�<�U�<��<c֓<��<�O�<���<D<g��<D/�<�c�<���< ʃ<���<�,�<s�|<y<�xu<�q<�4n<D�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<��M<�I<�^F<1�B<P4?<�;<�8<,�4<1<q|-<��)<�~&<�#<^�<�!<y�<}P<��<M�<|><��<Ǥ<a<�G�;���;{�;V)�;���;(��;"��;mt�;�l�;tu�;���;��;��;8�;.��;���;yx�;��;t��;Q�;��;�;�y; jo;�oe;��[;~�Q;�IH;��>;"}5;oF,;�.#;�5;�Z;ޜ;��:���:��:���:c�:��:H�:Q�:��z:\:�v=:"@:]:���9��9_:&9�N8F�x��.�R"��Elƹ�:��K��;�4�؅O�Sj�u9��tQ��.S���?�����}�º�Ϻ�1ܺG��1D��� �G�u:�C`�������ʱ%���+���1�h�7���=�U�C���I��O�J�U���[���a�L�g�ױm�i�s�Řy����P���������x���h������Ġ��:�������  �  ;m==��=L=D�=2�=�(=0� =Je =� =�@�<�z�<���<c��<�#�<�Z�<1��<���<w��<�*�<D\�<R��<A��<���<��<�?�<�h�<n��<r��<���<]��<-�<=�< Z�<�t�<���<h��<���<���<���<���<W��<W��<���<�<��<d��<��<���<���<���<���<��<���<�o�<pN�<N)�<n �<���<-��<�n�<%6�<���<���<Xt�<x+�<���<d��<#8�<���<���<(�<2��<O�<��<�n�<3��<�}�<���<M}�<O��<tm�<�߱<�N�<��<�!�<O��<y�<WE�<6��<���<�L�<ߞ�</�<�:�<��<�̚<q�<�U�<��<i֓<��<�O�<���<5<q��<I/�<�c�<���<ʃ<���<�,�<x�|<y<�xu<�q<�4n<k�j<��f<�Mc<�_<�
\<�jX<y�T<�-Q<��M<�I<�^F<<�B<G4?<�;<�8<�4<"1<k|-<��)<�~&<�#<Y�<x!<t�<hP<��<I�<�><��<��<;a<�G�;���;{�;V)�;���;��;&��;Ht�;m�;Ru�;���;A��;��;g8�;��;���;hx�;��;r��;�P�;��; �;Z�y;�io;ipe;ɗ[;"�Q;JH;d�>;�}5;XF,;�.#;g5;;Z;��;���:���:O�:���:��:��:M�:��:��z:�\:�v=:;?:�\:R��9*�91@&9�M8�lx�O�.�����iƹ�=�����O�4�؅O��j��9��wQ��SS��??��V��W�º��Ϻ�1ܺ��躍D���� ����:��`�΀�����%���+�/�1���7�B�=��C���I���O�"�U���[���a�o�g�±m�٥s���y����g���˸������5���m����������q��������  �  >m==��=L=E�=/�=�(=7� =He =� =�@�<�z�< ��<g��<�#�<�Z�<9��<���<l��<�*�<D\�<\��<5��<���<��<�?�<�h�<h��<w��<���<j��<*�<=�<�Y�<�t�<���<X��<¸�<���<���<���<_��<V��<���<%�<��<h��<��<���<���<���<���<��<���<�o�<wN�<W)�<v �<���<"��<�n�<6�<���<���<Ht�<|+�<���<l��<!8�<���<��<0�<7��<O�<��<�n�<&��<�}�<���<R}�<J��<�m�<�߱<�N�<��<�!�<Q��<v�<WE�<(��<���<�L�<֞�<&�<�:�<!��<�̚<{�<�U�<��<i֓<��<�O�<���<A<g��<A/�<�c�<���<$ʃ<���<�,�<~�|< y<�xu<	�q<�4n<J�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<��M<�I<�^F<9�B<L4?<��;<�8<)�4<1<]|-<��)<�~&<�#<`�<�!<�<xP<��<4�<z><��<��<#a<�G�;���;{�;o)�;���;-��;1��;|t�;m�;]u�;���; ��;��;%8�;%��;���;wx�;��;���;�P�;��;!�;@�y;�io;�oe;��[;d�Q;�IH;H�>;"}5;qF,;�.#;�5;�Z;�;��:��:�:��:6�:��:T�:�:D�z:�\:�v=:$?:�]:.��9~�9�<&95N8��x�	�.��#���jƹ�<�������4�`�O�j��9��DQ��6S��l?��M��=�º*�Ϻ�1ܺ��E���� �M�k:�]`���������%��+�a�1��7���=�V�C���I���O��U���[���a�a�g���m�b�s���y����\������$���z���d����������5���󜚻�  �  *l=�=:�=hJ=e�=�=�&=�� =|b =  =U:�<�s�<���<y��<�<�Q�<ǆ�<ں�<���<��<�P�<)��<d��<L��<��<�0�<oY�<c��<���<o��<R��<`�<�)�<�E�<�_�<x�<��<���<ݲ�<���</��<��<=��<���<���<T��<K��<,��<���<���<а�<��<p��<�j�<'L�<"*�<q�<��<׭�<�|�<�G�<��<��<I��<[L�<]�<8��<e�<��<F��<�X�<��<D��<g'�<|��<�G�<�Ѻ<�W�<�ٷ<KX�<�Ҵ<�I�<ټ�<a,�<u��<�<bf�<bȩ<='�<���<�ۤ<�1�<���<՟<�"�<
n�<鶚<���<�A�<e��<�ē<q�<T@�<w{�<>��<��<�$�<^Z�<��<�<���<�'�<ʲ|<�y<�uu<b�q<O6n<5�j<5�f<5Vc<��_<
\<	zX<M�T<�AQ<ɧM<�J<�yF<c�B<�S?<��;<�88<��4<�)1<`�-<�(*<ڭ&<K7#<��<HW<e�<��<�+<��<�~<�0<��<�<=��;vm�;�;���;2��;0P�;(-�;��;��;��;�8�;$c�;���;�;C�;箢;)+�;<��;�U�;w�;�Ç;,��;��z;��p;��f;��\;�<S;��I;z)@;��6;ٓ-;{w$;�y;S�;g�	;P0;�K�:�o�:��:�S�:��:U�:�(�:��~:8�_:�JA:O�":b�:Ӡ�9g�9�}39��8��F�6�"�LM��8�������f.�^=2�YM��g�c���;���H��@��["������v�κ[ۺ���9���~ �I�����a��4��S��m%���+�r�1�&�7���=��C� �I�|�O��U���[�`�a�j�g��m�ˏs�l�y�0|�v��������'���娎�����^���s���ѣ���  �  5l=�=7�=mJ=b�=�=�&=�� =�b =���<C:�<�s�<���<���<��<�Q�<ņ�<ݺ�<���<��<�P�<��<W��<<��<��<�0�<mY�<r��<˥�<p��<J��<h�<�)�<�E�<�_�<�w�<��<���<޲�<���<,��<��<O��<���<~��<]��<:��<��<���<~��<԰�<Ϝ�<j��<�j�<,L�<**�<z�<��<ӭ�<�|�<�G�<��<��<7��<JL�<K�<A��<e�<��<V��<�X�<��<?��<m'�<x��<�G�<�Ѻ<�W�<�ٷ<CX�<�Ҵ<�I�<ټ�<q,�<���< �<bf�<gȩ<.'�<<�ۤ<�1�<���<�ԟ<�"�<n�<�<���<B�<d��<�ē<b�<<@�<�{�<3��<~�<{$�<SZ�<��<�<���<�'�<ֲ|<�y<�uu<Z�q<U6n<A�j<��f<>Vc<��_<\<zX<@�T<�AQ<��M<�J<wyF<w�B<�S?<��;<�88<{�4<�)1<8�-<�(*<ޭ&<K7#<�<_W<x�<��<�+<[�<�~<�0<��<�<���;sm�;"�;���;n��;uP�;--�;��;�;��;�8�;c�;E��;%�;C�;ﮢ;+�;.��;V�;��;ć;��;(�z;��p;<�f;z�\;}<S;��I;�(@;��6;��-;�w$;�y;��;��	;)0;�K�:1n�:���:�S�:x�::�:�'�:+�~:��_:�KA:e�":��:���9�9}�39��8�F�	�"��P��w�������`-�6>2�LM�(�g�b���;���H���?��P#�������κ;Zۺ~������p~ �f������v4��S��m%�2�+�,�1� 7�N�=�r�C���I�гO���U���[���a�Šg���m���s�M�y�O|�h�������]������Ҩ��	���>������������  �  -l=�=3�=oJ=b�=�=�&=�� =�b =���<Q:�<�s�<���<}��<��<�Q�<���<��<���<��<�P�<��<l��<G��<��<�0�<dY�<`��<���<n��<H��<m�<�)�<�E�<�_�<�w�<���<z��<ز�<���<,��<��<<��<���<v��<e��<=��<0��<���<|��<ܰ�<ќ�<{��<�j�<*L�< *�<p�<
��<ϭ�<�|�<�G�<��<��<>��<aL�<P�<G��<e�<��<B��<�X�<��<>��<i'�<i��<�G�<�Ѻ<�W�<�ٷ<6X�<�Ҵ<�I�<ؼ�<f,�<s��<�<_f�<iȩ<5'�<��<�ۤ<�1�<���<�ԟ<�"�<�m�<춚<���<�A�<`��<�ē<r�<>@�<�{�<.��<��<�$�<TZ�<��<�<���<�'�<ʲ|<�y<�uu<E�q<I6n<R�j<��f<JVc<��_<�\<%zX<@�T<�AQ<קM<�J<eyF<��B<�S?<��;<�88<k�4<�)1<=�-<�(*<�&<>7#<�<MW<i�<p�<�+<n�<�~<�0<��<�<&��;vm�;%�;���;(��;CP�;#-�;��;�;P�;�8�;-c�;V��;K�;�B�;ծ�;+�;0��;�U�;s�;�Ç;���;f�z;�p;��f;��\;o<S;�I;�(@;�6;��-;�w$;|y;I�;��	;0;�L�:zn�:S��:�S�:��:��:�'�:��~:��_:�JA:��":��:���9��9f~39x��8��F���"�+N��K��� ����,�J>2�{M��g����p<���H���?���"��7�����κ&Zۺ<��m����} �������K��4��S��m%���+��1���7�y�=���C� �I�ʳO��U�7�[�b�a�L�g��m���s�)�y��|����g���_�������먎�8���)�������ʣ���  �  .l=�=?�=jJ=a�=�=�&=�� =~b =  =N:�<�s�<���<|��<��<�Q�<ǆ�<պ�<���<��<�P�<#��<[��<C��<��<�0�<|Y�<k��<¥�<o��<T��<a�<�)�<�E�<�_�< x�<��<���<ڲ�<���<1��<��<B��<���<���<V��<>��< ��<���<���<Ѱ�<ڜ�<k��<�j�<0L�<)*�<y�<��<ԭ�<�|�<�G�<��<��<<��<PL�<O�<;��<e�<��<I��<�X�<��<G��<h'�<���<�G�<�Ѻ<�W�<�ٷ<KX�<�Ҵ<�I�<ټ�<k,�<}��<-�<if�<^ȩ<4'�<�<�ۤ<�1�<���<�ԟ<�"�<	n�<<���<�A�<i��<�ē<k�<J@�<z{�<;��<~�<�$�<SZ�<��<�<���<�'�<̲|<�y<�uu<X�q<d6n<+�j<�f<#Vc<Ŷ_<\<zX<R�T<�AQ<ܧM<�J<�yF<l�B<�S?<��;<�88<��4<�)1<M�-<�(*<Э&<S7#<�<_W<m�<��<�+<p�<�~<�0<��<��<��;Qm�;5�;���;Q��;SP�;*-�;��;��;��;�8�;�b�;\��;��;MC�;߮�;4+�;A��;�U�;��;ć;Q��;��z;�p;k�f;��\;�<S;��I;)@;��6;��-;�w$;�y;��;��	;40;�K�:�n�:���:�S�:��:��:�'�:`�~:?�_:�LA:��":]�:n��97�9�}39���8��F�i�"�fQ��[�������:.��<2�OM�ռg����;��?H��?@���"��;����κ�Zۺ���:����~ �S�����	��4�wS��m%��+���1��7��=�o�C�]�I�γO��U�s�[��a�:�g��m���s�\�y�[|�I�������.���L�����������U���j���ƣ���  �  4l=�=7�=eJ=f�=�=�&=�� =~b =  =I:�<�s�<���<s��<��<�Q�<ֆ�<ۺ�<���<��<�P�<*��<R��<Q��<��<�0�<eY�<e��<ʥ�<d��<W��<V�<�)�<�E�<�_�<x�<ۍ�<���<ʲ�<���<%��<
��<H��<���<��<R��<O��<"��<���<���<Ͱ�<ޜ�<i��<�j�<'L�<#*�<v�<��<��<�|�<�G�<��<$��<B��<NL�<b�<9��<e�<��<K��<�X�<��<E��<V'�<���<~G�<�Ѻ<�W�<�ٷ<IX�<�Ҵ<�I�<˼�<p,�<x��<�<Zf�<bȩ<D'�<낦<�ۤ<�1�<���< ՟<�"�<n�<ᶚ<���<�A�<k��<�ē<f�<L@�<x{�<D��<|�<�$�<_Z�<��<�<���<�'�<Ų|<�y<�uu<F�q<m6n<"�j<1�f< Vc<̶_<�\<zX<O�T<�AQ<�M<�J<uyF<V�B<�S?<��;<�88<��4<�)1<N�-<�(*<�&<`7#<��<kW<Z�<��<�+<s�<�~<�0<��<�<R��;om�;��;���;<��;qP�;�,�;��;��;��;�8�;�b�;���;��;]C�;���;!+�;��;�U�;��;�Ç;��;��z;��p;y�f;��\;�<S;w�I;.)@;~�6;)�-;~w$;�y;}�;N�	;�0;�K�:Mo�:���:XT�:(�:��:)�:%�~:y�_:7JA:�":��:[��9��9Qu39K��8��F�ק"��O��E���]����/�<2�M�?�g�3���<��2I��@���!������z�κfZۺP������~ �Ĵ�8�����4�kS�{m%��+���1�#�7�̩=���C�)�I�r�O�C�U��[�Y�a��g��m��s���y��|�8���Ǵ������R����������m���o���棚��  �  /l=�=8�=pJ=a�=�=�&=�� =�b =  =N:�<�s�<���<{��<��<�Q�<ņ�<��<���<��<�P�<��<a��<B��<��<�0�<lY�<d��<å�<e��<Q��<n�<�)�<�E�<�_�<x�<��<���<ײ�<���<&��<��<>��<���<���<d��<<��<!��<���<|��<װ�<֜�<s��<�j�<'L�<)*�<z�<��<ڭ�<�|�<�G�<��<��<9��<RL�<M�<E��<e�<��<D��<�X�<��<M��<g'�<t��<�G�<�Ѻ<�W�<�ٷ<;X�<�Ҵ<�I�<ϼ�<l,�<v��<�<if�<eȩ<1'�<���<�ۤ<�1�<���<�ԟ<�"�<
n�<㶚<���<�A�<b��<�ē<m�<F@�<�{�</��<��<�$�<QZ�<��<�<���<�'�<Ȳ|<�y<�uu<J�q<V6n<7�j<�f</Vc<��_<�\<-zX<C�T<�AQ<ߧM<�J<{yF<��B<�S?<��;<�88<p�4<�)1<I�-<�(*<�&<F7#<�<iW<^�<��<�+<o�<�~<�0<��<�<��;nm�;E�;���;9��;VP�;-�;��;�;`�;�8�;c�;_��;�; C�;Ѯ�;S+�;��;V�;~�;�Ç;-��;e�z;�p;q�f;��\;l<S;̢I;�(@;��6;��-;{w$;�y;��;]�	;i0;<L�:�n�:'��:�S�:��:��:�'�:��~:n�_:{KA:%�":��:m��9��9�}39��8��F���"�{P���������� -��<2��M���g�R���;��BH���?��"#��������κbZۺD��B���.~ �F��-�����4��S��m%�Ղ+��1���7�p�=�8�C�o�I��O�w�U��[�P�a�7�g���m��s��y��|�f�������?���3���ը��1����������ᣚ��  �  ,l=�=5�=nJ=d�=�=�&=�� =�b =���<Q:�<�s�<���<���<~�<�Q�<���<��<���<��<�P�<��<k��<<��<��<�0�<lY�<m��<���<w��<A��<i�<�)�<�E�<�_�<�w�<��<���<ٲ�<���<%��<��<:��<���<u��<e��<=��<)��<���<���<��<͜�<{��<�j�<2L�<"*�<p�<��<ҭ�<�|�<�G�<��<!��<8��<]L�<L�<H��<e�<��<B��<�X�<��<9��<j'�<r��<�G�<�Ѻ<�W�<�ٷ<9X�<�Ҵ<�I�<߼�<i,�<z��< �<^f�<mȩ<,'�<��<�ۤ<�1�<���<�ԟ<�"�<n�<���<���<B�<h��<�ē<s�<8@�<�{�<2��<��<�$�<WZ�<��<�<���<�'�<�|<�y<�uu<K�q<Q6n<F�j<��f<:Vc<��_<�\<zX<0�T<�AQ<ҧM<�J<kyF<z�B<�S?<��;<�88<u�4<�)1<1�-<�(*<߭&<M7#<�<HW<��<z�<�+<l�<�~<�0<��<�<���;�m�;$�;���;\��;EP�;H-�;��;�;Z�;�8�;c�;;��;/�;C�;ۮ�;+�;��;V�;o�;-ć;���;h�z;�p;��f;��\;�<S;�I;�(@;�6;��-;�w$;�y;K�;��	;#0;�L�:>n�:o��:(T�:��:z�:�'�:�~:��_:�LA:��":��:|��9���9!39̩�8 �F��"�dQ������H���K-��>2�~M��g����;���H��H?��o#��8�����κ�Yۺ��纕���-~ �~�����b�|4��S��m%���+�O�1�q�7�U�=��C�W�I���O���U�0�[�ӧa�d�g���m�7�s�V�y��|�p������^������ը��+���@������������  �  +l=�=6�=jJ=g�=�=�&=�� =�b =   =Z:�<�s�<���<���<��<�Q�<ņ�<��<���<��<�P�<��<Z��<G��<��<�0�<hY�<h��<���<m��<O��<b�<�)�<�E�<�_�<x�<ٍ�<���<ز�<���<)��<	��<;��<���<x��<]��<I��<&��<���<���<Ұ�<ޜ�<z��<�j�<-L�<&*�<w�<��<ҭ�<�|�<�G�<��<!��<8��<VL�<Y�<C��<e�<��<C��<�X�<
��<C��<e'�<{��<{G�<�Ѻ<�W�<�ٷ<CX�<�Ҵ<�I�<ռ�<c,�<y��<�<\f�<oȩ<9'�<�<�ۤ<�1�<���<	՟<�"�<n�<�<���<B�<f��<�ē<z�<G@�<|{�<7��<��<�$�<^Z�<��<�<���<�'�<Ͳ|<�y<�uu<K�q<V6n<"�j<�f< Vc<��_<�\<zX<E�T<�AQ<ͧM<�J<ryF<k�B<�S?<��;<�88<��4<�)1<G�-<�(*<ܭ&<K7#<�<XW<v�<��<�+<��<�~<�0<��<��<+��;�m�;�;���;G��;6P�;%-�;��;��;��;�8�;�b�;v��;��;0C�;خ�;"+�;#��;�U�;s�;ć;��;+�z;r�p;��f;��\;�<S;��I;/)@;
�6;��-;�w$;�y;��;��	;*0;oL�:io�:���:0T�:��:�:�(�:t�~:��_:?KA:�":�:3��9.�9�|39���8��F���"�P��"�������G.��=2��M�νg�$��D<��I��1?���"��D���O�κ5Zۺv��q��=~ �]�������4��S��m%�t�+�ד1���7�/�=�U�C�J�I�w�O�رU��[�"�a�t�g��m��s�U�y��|�f���Ǵ�����R���ۨ��!���J�������ˣ���  �  7l=�=<�=nJ=\�=�=�&=�� =�b =  =D:�<�s�<���<{��<��<�Q�<ц�<ݺ�<���<��<�P�<'��<Y��<E��<��<�0�<oY�<a��<Υ�<`��<V��<Z�<�)�<�E�<�_�<x�<؍�<���<β�<���<'��<
��<J��<���<���<W��<<��<��<���<���<Ͱ�<ߜ�<e��<�j�<*L�<,*�<��<��<��<�|�<�G�<��<!��<>��<KL�<P�<:��<e�<��<N��<�X�<��<J��<['�<���<yG�<�Ѻ<�W�<�ٷ<HX�<�Ҵ<�I�<ɼ�<r,�<x��<�<nf�<Yȩ<7'�<<�ۤ<�1�<���<�ԟ<�"�<n�<嶚<���<�A�<j��<�ē<b�<N@�<|{�<>��<��<�$�<KZ�<��<�<���<�'�<��|<�y<�uu<>�q<w6n<�j<!�f<Vc<Ӷ_<�\<zX<J�T<�AQ<��M<�J<�yF<}�B<�S?<��;<�88<��4<�)1<V�-<�(*<�&<[7#<�<yW<_�<��<�+<e�<�~<�0<��<�<"��;4m�;O�;���;-��;�P�;�,�;��;��;��;�8�;�b�;n��;��;mC�;���;;+�;��; V�;��;�Ç;T��;��z;�p;G�f;��\;�<S;~�I;1)@;`�6;,�-;�w$;�y;Ι;r�	;�0;\K�:o�:���:6T�:��:[�:�'�:H�~:��_:cJA:e�":��:���9��9�w390��8��F���"��Q������w���/��<2�2M��g�,��<���G���@���"��������κ`Zۺx��]����~ ��������4�sS�nm%�3�+���1��7���=�N�C�s�I��O���U���[���a� g��m��s�R�y��|�#���մ�����l�������+���T���z�����  �  1l=�=6�=iJ=b�=�=�&=�� =�b =  =K:�<�s�<���<{��<��<�Q�<̆�<��<���<��<�P�<��<e��<T��<��<�0�<iY�<b��<ť�<d��<T��<`�<�)�<�E�<�_�<x�<��<���<Ȳ�<���<$��<��<D��<���<|��<V��<J��<2��<���<���<۰�<ݜ�<s��<�j�<*L�<$*�<t�<	��<��<�|�<�G�<��< ��<>��<`L�<^�<;��<e�<��<H��<�X�<��<C��<X'�<t��<�G�<�Ѻ<�W�<�ٷ<9X�<�Ҵ<�I�<μ�<j,�<t��<�<^f�<_ȩ<D'�<���<�ۤ<�1�<���<�ԟ<�"�<n�<붚<���<�A�<h��<�ē<j�<J@�<�{�<6��<��<�$�<XZ�<��<�<���<�'�<��|<�y<�uu<2�q<[6n<-�j<�f<#Vc<��_<�\<zX<G�T<�AQ<�M<�J<syF<g�B<�S?<��;<�88<~�4<�)1<S�-<�(*<��&<T7#<�<`W<j�<��<�+<p�<�~<�0<��<�<_��;`m�;�;���;1��;aP�;�,�;��;��;Y�;�8�;�b�;h��;�;"C�;���;$+�;��;�U�;��;�Ç;��;��z;z�p;�f;��\;�<S;�I;%)@;��6;1�-;�w$;�y;n�;{�	;�0;dL�:&o�:s��:T�:��:��:�(�:y�~:D�_:�JA:��":��:���9E�9,v39e��81�F���"�#P�����)���/�=2��M���g�g��><���H��+@���!�������κyZۺ������~ �
�������4�}S�Am%��+���1���7�7�=�!�C�˲I���O��U���[�W�a��g�*�m��s�N�y��|�[�������1���K���Ũ��Q���I������񣚻�  �  *l=�=:�=kJ=f�=�=�&=�� =�b =���<W:�<�s�<���<���<�<�Q�<���<��<���<��<�P�<��<Y��<;��<��<�0�<sY�<o��<���<r��<G��<h�<�)�<�E�<�_�<�w�<��<~��<��<���<+��<��<<��<���<|��<a��<=��<��<���<}��<ڰ�<ќ�<|��<�j�<5L�<.*�<{�<��<ɭ�<�|�<�G�<��<��<6��<ML�<M�<F��<e�<��<G��<�X�<��<=��<n'�<n��<�G�<�Ѻ<�W�<�ٷ<;X�<�Ҵ<�I�<ڼ�<c,�<��<'�<]f�<nȩ<-'�<���<�ۤ<�1�<���<�ԟ<�"�<�m�<���<���<B�<e��<�ē<w�<?@�<�{�<3��<}�<~$�<XZ�<��<�<���<�'�<ֲ|<�y<�uu<X�q<D6n<*�j<�f<&Vc<��_<�\<zX<;�T<�AQ<ɧM<�J<�yF<p�B<�S?<��;<�88<y�4<�)1<A�-<�(*<ح&<C7#<)�<JW<��<s�<�+<w�<�~<�0<��<�<���;�m�;�;���;e��;3P�;5-�;��;�;t�;�8�;�b�;G��;�;C�;���;+�;+��;V�;x�;2ć;��;J�z;�p;V�f;w�\;z<S;�I;�(@;�6;��-;�w$;�y;��;��	;�/;�L�:�n�:L��:�S�:u�:z�:�'�:��~:?�_:	MA:��":�:ğ�9��9��39H��8��F���"��Q����������`-�N>2�M�νg����T;���H��C?��W#��m���q�κ�Zۺ ��;���8~ ����F��;�-4��S��m%���+��1���7�Q�=�s�C���I���O�ǱU�֭[�ʧa���g���m��s�W�y�W|���������S���E���𨎻���B������������  �  .l=�=3�=lJ=c�=�=�&=�� =�b =���<R:�<�s�<���<���<�<�Q�<Æ�<��<���<��<�P�<,��<e��<D��<��<�0�<aY�<a��<���<m��<E��<W�<�)�<�E�<�_�<x�<��<���<в�<���<&��<
��<;��<���<v��<^��<B��<'��<���<���<۰�<Ҝ�<{��<�j�</L�<%*�<s�<��<׭�<�|�<�G�<��<$��<J��<WL�<T�<A��<e�<��<B��<�X�<��<7��<\'�<s��<�G�<�Ѻ<�W�<�ٷ<;X�<�Ҵ<�I�<Ӽ�<f,�<s��<�<Zf�<fȩ<5'�<���<�ۤ<�1�<���<�ԟ<�"�<n�<���<���<B�<e��<�ē<s�<@@�<�{�<A��<��<�$�<VZ�<��<�<���<�'�<Ӳ|<�y<�uu<C�q<W6n<:�j<�f<3Vc<��_<�\<�yX<7�T<�AQ<اM<�J<eyF<r�B<�S?<��;<�88<��4<�)1<B�-<�(*<�&<L7#<�<JW<��<�<�+<p�<�~<�0<��<�<��;ym�;�;���;,��;FP�;#-�;��;��;g�;�8�;c�;j��;�;C�;���;�*�;��;�U�;s�;�Ç;���;2�z;;�p;��f;�\;�<S;�I;�(@;�6;�-;�w$;�y;i�;��	;T0;�L�:�n�:_��:aT�:��:�:?(�:>�~:��_:JA:��":�:=��9:��9�x39���8��F�ƫ"��O��?�������p/��>2�M�q�g�����<��-I���?���"������@�κZۺ*��R����} �r�����T�h4��S�xm%���+��1���7��=��C�>�I���O�űU�1�[�n�a�O�g�˘m��s���y��|�d�������-���*���Ө��1���u�������ȣ���  �  4l=�=:�=nJ=_�=�=�&=�� =�b =  =J:�<�s�<���<���<��<�Q�<���<��<���<��<�P�<��<X��<L��<��<�0�<qY�<n��<ȥ�<a��<]��<d�<�)�<�E�<�_�<�w�<���<���<ϲ�<���<-��<��<M��<���<���<W��<A��<#��<���<y��<ܰ�<؜�<s��<�j�<'L�<4*�<��<��<ݭ�<�|�<�G�<��<��<:��<OL�<V�<8��<e�<��<T��<�X�<��<U��<]'�<x��<G�<�Ѻ<�W�<�ٷ<?X�<�Ҵ<�I�<˼�<m,�<���<$�<kf�<]ȩ<<'�<���<�ۤ<�1�<���<�ԟ<�"�<n�<�<���<	B�<_��<�ē<k�<I@�<�{�<-��<�<�$�<QZ�<��<�<���<�'�<��|<�y<�uu<;�q<[6n<&�j<��f<Vc<��_<�\<$zX<Y�T<�AQ<�M<�J<�yF<|�B<�S?<��;<�88<k�4<�)1<P�-<�(*<��&<A7#<�<�W<r�<x�<�+<n�<�~<�0<��<�<=��;Um�;K�;���;b��;lP�;�,�;�;��;u�;�8�;�b�;=��;��;+C�;���;h+�;5��;�U�;��;ć;;��;��z;6�p;��f;��\;V<S;�I; )@;��6;�-;�w$;z;�;q�	;0;RL�:�n�:���:�S�:��:��:T(�:�~:��_:LA:-�":��:`��9��9y39���8��F�j�"��Q���������p.��;2�M���g�����;��H��F@��q"��c���n�κ�Zۺ���$��� ~ �z�������L4��S�.m%��+�Ǔ1���7�|�=�g�C�0�I��O���U���[��a�ؠg�]�m�Əs���y��|�\�������^���W���Ш��>���*���[�������  �  .l=�=3�=lJ=c�=�=�&=�� =�b =���<R:�<�s�<���<���<�<�Q�<Æ�<��<���<��<�P�<,��<e��<D��<��<�0�<aY�<a��<���<m��<E��<W�<�)�<�E�<�_�<x�<��<���<в�<���<&��<
��<;��<���<v��<^��<B��<'��<���<���<۰�<Ҝ�<{��<�j�</L�<%*�<s�<��<׭�<�|�<�G�<��<$��<J��<WL�<T�<A��<e�<��<B��<�X�<��<7��<\'�<s��<�G�<�Ѻ<�W�<�ٷ<;X�<�Ҵ<�I�<Ӽ�<f,�<s��<�<Zf�<fȩ<5'�<���<�ۤ<�1�<���<�ԟ<�"�<n�<���<���<B�<e��<�ē<s�<@@�<�{�<A��<��<�$�<VZ�<��<�<���<�'�<Ӳ|<�y<�uu<C�q<W6n<:�j<�f<3Vc<��_<�\<�yX<7�T<�AQ<اM<�J<eyF<r�B<�S?<��;<�88<��4<�)1<B�-<�(*<�&<L7#<�<JW<��<�<�+<p�<�~<�0<��<�<��;ym�;�;���;,��;FP�;#-�;��;��;g�;�8�;c�;j��;�;C�;���;�*�;��;�U�;s�;�Ç;���;2�z;;�p;��f;�\;�<S;�I;�(@;�6;�-;�w$;�y;i�;��	;T0;�L�:�n�:_��:aT�:��:�:?(�:>�~:��_:JA:��":�:=��9:��9�x39���8��F�ƫ"��O��?�������p/��>2�M�q�g�����<��-I���?���"������@�κZۺ*��R����} �r�����T�h4��S�xm%���+��1���7��=��C�>�I���O�űU�1�[�n�a�O�g�˘m��s���y��|�d�������-���*���Ө��1���u�������ȣ���  �  *l=�=:�=kJ=f�=�=�&=�� =�b =���<W:�<�s�<���<���<�<�Q�<���<��<���<��<�P�<��<Y��<;��<��<�0�<sY�<o��<���<r��<G��<h�<�)�<�E�<�_�<�w�<��<~��<��<���<+��<��<<��<���<|��<a��<=��<��<���<}��<ڰ�<ќ�<|��<�j�<5L�<.*�<{�<��<ɭ�<�|�<�G�<��<��<6��<ML�<M�<F��<e�<��<G��<�X�<��<=��<n'�<n��<�G�<�Ѻ<�W�<�ٷ<;X�<�Ҵ<�I�<ڼ�<c,�<��<'�<]f�<nȩ<-'�<���<�ۤ<�1�<���<�ԟ<�"�<�m�<���<���<B�<e��<�ē<w�<?@�<�{�<3��<}�<~$�<XZ�<��<�<���<�'�<ֲ|<�y<�uu<X�q<D6n<*�j<�f<&Vc<��_<�\<zX<;�T<�AQ<ɧM<�J<�yF<p�B<�S?<��;<�88<y�4<�)1<A�-<�(*<ح&<C7#<)�<JW<��<s�<�+<w�<�~<�0<��<�<���;�m�;�;���;e��;3P�;5-�;��;�;t�;�8�;�b�;G��;�;C�;���;+�;+��;V�;x�;2ć;��;J�z;�p;V�f;w�\;z<S;�I;�(@;�6;��-;�w$;�y;��;��	;�/;�L�:�n�:L��:�S�:u�:z�:�'�:��~:?�_:	MA:��":�:ß�9��9��39H��8��F���"��Q����������`-�N>2�M�νg����T;���H��C?��W#��m���q�κ�Zۺ ��;���8~ ����F��;�-4��S��m%���+��1���7�Q�=�s�C���I���O�ǱU�֭[�ʧa���g���m��s�W�y�W|���������S���E���𨎻���B������������  �  1l=�=6�=iJ=b�=�=�&=�� =�b =  =K:�<�s�<���<{��<��<�Q�<̆�<��<���<��<�P�<��<e��<T��<��<�0�<iY�<b��<ť�<d��<T��<`�<�)�<�E�<�_�<x�<��<���<Ȳ�<���<$��<��<D��<���<|��<V��<J��<2��<���<���<۰�<ݜ�<s��<�j�<*L�<$*�<t�<	��<��<�|�<�G�<��< ��<>��<`L�<^�<;��<e�<��<H��<�X�<��<C��<X'�<t��<�G�<�Ѻ<�W�<�ٷ<9X�<�Ҵ<�I�<μ�<j,�<t��<�<^f�<_ȩ<D'�<���<�ۤ<�1�<���<�ԟ<�"�<n�<붚<���<�A�<h��<�ē<j�<J@�<�{�<6��<��<�$�<XZ�<��<�<���<�'�<��|<�y<�uu<2�q<[6n<-�j<�f<#Vc<��_<�\<zX<G�T<�AQ<�M<�J<syF<g�B<�S?<��;<�88<~�4<�)1<S�-<�(*<��&<T7#<�<`W<j�<��<�+<p�<�~<�0<��<�<_��;`m�;�;���;1��;aP�;�,�;��;��;Y�;�8�;�b�;h��;�;"C�;���;$+�;��;�U�;��;�Ç;��;��z;z�p;�f;��\;�<S;�I;%)@;��6;1�-;�w$;�y;n�;{�	;�0;dL�:&o�:s��:T�:��:��:�(�:y�~:D�_:�JA:��":��:���9E�9,v39e��81�F���"�#P�����)���/�=2��M���g�g��><���H��+@���!�������κyZۺ������~ �
�������4�}S�Am%��+���1���7�7�=�!�C�˲I���O��U���[�W�a��g�*�m��s�N�y��|�[�������1���K���Ũ��Q���I������񣚻�  �  7l=�=<�=nJ=\�=�=�&=�� =�b =  =D:�<�s�<���<{��<��<�Q�<ц�<ݺ�<���<��<�P�<'��<Y��<E��<��<�0�<oY�<a��<Υ�<`��<V��<Z�<�)�<�E�<�_�<x�<؍�<���<β�<���<'��<
��<J��<���<���<W��<<��<��<���<���<Ͱ�<ߜ�<e��<�j�<*L�<,*�<��<��<��<�|�<�G�<��<!��<>��<KL�<P�<:��<e�<��<N��<�X�<��<J��<['�<���<yG�<�Ѻ<�W�<�ٷ<HX�<�Ҵ<�I�<ɼ�<r,�<x��<�<nf�<Yȩ<7'�<<�ۤ<�1�<���<�ԟ<�"�<n�<嶚<���<�A�<j��<�ē<b�<N@�<|{�<>��<��<�$�<KZ�<��<�<���<�'�<��|<�y<�uu<>�q<w6n<�j<!�f<Vc<Ӷ_<�\<zX<J�T<�AQ<��M<�J<�yF<}�B<�S?<��;<�88<��4<�)1<V�-<�(*<�&<[7#<�<yW<_�<��<�+<e�<�~<�0<��<�<"��;4m�;O�;���;-��;�P�;�,�;��;��;��;�8�;�b�;n��;��;mC�;���;;+�;��; V�;��;�Ç;T��;��z;�p;G�f;��\;�<S;~�I;1)@;`�6;,�-;�w$;�y;Ι;r�	;�0;\K�:o�:���:6T�:��:[�:�'�:H�~:��_:cJA:e�":��:���9��9�w390��8��F���"��Q������w���/��<2�2M��g�,��<���G���@���"��������κ`Zۺx��]����~ ��������4�sS�nm%�3�+���1��7���=�N�C�s�I��O���U���[���a� g��m��s�R�y��|�#���մ�����l�������+���T���z�����  �  +l=�=6�=jJ=g�=�=�&=�� =�b =   =Z:�<�s�<���<���<��<�Q�<ņ�<��<���<��<�P�<��<Z��<G��<��<�0�<hY�<h��<���<m��<O��<b�<�)�<�E�<�_�<x�<ٍ�<���<ز�<���<)��<	��<;��<���<x��<]��<I��<&��<���<���<Ұ�<ޜ�<z��<�j�<-L�<&*�<w�<��<ҭ�<�|�<�G�<��<!��<8��<VL�<Y�<C��<e�<��<C��<�X�<
��<C��<e'�<{��<{G�<�Ѻ<�W�<�ٷ<CX�<�Ҵ<�I�<ռ�<c,�<y��<�<\f�<oȩ<9'�<�<�ۤ<�1�<���<	՟<�"�<n�<�<���<B�<f��<�ē<z�<G@�<|{�<7��<��<�$�<^Z�<��<�<���<�'�<Ͳ|<�y<�uu<K�q<V6n<"�j<�f< Vc<��_<�\<zX<E�T<�AQ<ͧM<�J<ryF<k�B<�S?<��;<�88<��4<�)1<G�-<�(*<ܭ&<K7#<�<XW<v�<��<�+<��<�~<�0<��<��<+��;�m�;�;���;G��;6P�;%-�;��;��;��;�8�;�b�;v��;��;0C�;خ�;"+�;#��;�U�;s�;ć;��;+�z;r�p;��f;��\;�<S;��I;/)@;
�6;��-;�w$;�y;��;��	;*0;oL�:io�:���:0T�:��:�:�(�:t�~:��_:?KA:�":�:3��9.�9�|39���8��F���"�P��"�������G.��=2��M�νg�$��D<��I��1?���"��D���O�κ5Zۺv��q��=~ �]�������4��S��m%�t�+�ד1���7�/�=�U�C�J�I�w�O�رU��[�"�a�t�g��m��s�U�y��|�f���Ǵ�����R���ۨ��!���J�������ˣ���  �  ,l=�=5�=nJ=d�=�=�&=�� =�b =���<Q:�<�s�<���<���<~�<�Q�<���<��<���<��<�P�<��<k��<<��<��<�0�<lY�<m��<���<w��<A��<i�<�)�<�E�<�_�<�w�<��<���<ٲ�<���<%��<��<:��<���<u��<e��<=��<)��<���<���<��<͜�<{��<�j�<2L�<"*�<p�<��<ҭ�<�|�<�G�<��<!��<8��<]L�<L�<H��<e�<��<B��<�X�<��<9��<j'�<r��<�G�<�Ѻ<�W�<�ٷ<9X�<�Ҵ<�I�<߼�<i,�<z��< �<^f�<mȩ<,'�<��<�ۤ<�1�<���<�ԟ<�"�<n�<���<���<B�<h��<�ē<s�<8@�<�{�<2��<��<�$�<WZ�<��<�<���<�'�<�|<�y<�uu<K�q<Q6n<F�j<��f<:Vc<��_<�\<zX<0�T<�AQ<ҧM<�J<kyF<z�B<�S?<��;<�88<u�4<�)1<1�-<�(*<߭&<M7#<�<HW<��<z�<�+<l�<�~<�0<��<�<���;�m�;$�;���;\��;EP�;H-�;��;�;Z�;�8�;c�;;��;/�;C�;ۮ�;+�;��;V�;o�;-ć;���;h�z;�p;��f;��\;�<S;�I;�(@;�6;��-;�w$;�y;K�;��	;#0;�L�:>n�:o��:(T�:��:z�:�'�:�~:��_:�LA:��":��:|��9���9!39̩�8 �F��"�dQ������H���K-��>2�~M��g����;���H��H?��o#��8�����κ�Yۺ��纕���-~ �~�����b�|4��S��m%���+�O�1�q�7�U�=��C�W�I���O���U�0�[�ӧa�d�g���m�7�s�V�y��|�p������^������ը��+���@������������  �  /l=�=8�=pJ=a�=�=�&=�� =�b =  =N:�<�s�<���<{��<��<�Q�<ņ�<��<���<��<�P�<��<a��<B��<��<�0�<lY�<d��<å�<e��<Q��<n�<�)�<�E�<�_�<x�<��<���<ײ�<���<&��<��<>��<���<���<d��<<��<!��<���<|��<װ�<֜�<s��<�j�<'L�<)*�<z�<��<ڭ�<�|�<�G�<��<��<9��<RL�<M�<E��<e�<��<D��<�X�<��<M��<g'�<t��<�G�<�Ѻ<�W�<�ٷ<;X�<�Ҵ<�I�<ϼ�<l,�<v��<�<if�<eȩ<1'�<���<�ۤ<�1�<���<�ԟ<�"�<
n�<㶚<���<�A�<b��<�ē<m�<F@�<�{�</��<��<�$�<QZ�<��<�<���<�'�<Ȳ|<�y<�uu<J�q<V6n<7�j<�f</Vc<��_<�\<-zX<C�T<�AQ<ߧM<�J<{yF<��B<�S?<��;<�88<p�4<�)1<I�-<�(*<�&<F7#<�<iW<^�<��<�+<o�<�~<�0<��<�<��;nm�;E�;���;9��;VP�;-�;��;�;`�;�8�;c�;_��;�; C�;Ѯ�;S+�;��;V�;~�;�Ç;-��;e�z;�p;q�f;��\;l<S;̢I;�(@;��6;��-;{w$;�y;��;]�	;i0;<L�:�n�:'��:�S�:��:��:�'�:��~:n�_:{KA:%�":��:m��9��9�}39��8��F���"�{P���������� -��<2��M���g�R���;��BH���?��"#��������κbZۺD��B���.~ �F��-�����4��S��m%�Ղ+��1���7�p�=�8�C�o�I��O�w�U��[�P�a�7�g���m��s��y��|�f�������?���3���ը��1����������ᣚ��  �  4l=�=7�=eJ=f�=�=�&=�� =~b =  =I:�<�s�<���<s��<��<�Q�<ֆ�<ۺ�<���<��<�P�<*��<R��<Q��<��<�0�<eY�<e��<ʥ�<d��<W��<V�<�)�<�E�<�_�<x�<ۍ�<���<ʲ�<���<%��<
��<H��<���<��<R��<O��<"��<���<���<Ͱ�<ޜ�<i��<�j�<'L�<#*�<v�<��<��<�|�<�G�<��<$��<B��<NL�<b�<9��<e�<��<K��<�X�<��<E��<V'�<���<~G�<�Ѻ<�W�<�ٷ<IX�<�Ҵ<�I�<˼�<p,�<x��<�<Zf�<bȩ<D'�<낦<�ۤ<�1�<���< ՟<�"�<n�<ᶚ<���<�A�<k��<�ē<f�<L@�<x{�<D��<|�<�$�<_Z�<��<�<���<�'�<Ų|<�y<�uu<F�q<m6n<"�j<1�f< Vc<̶_<�\<zX<O�T<�AQ<�M<�J<uyF<V�B<�S?<��;<�88<��4<�)1<N�-<�(*<�&<`7#<��<kW<Z�<��<�+<s�<�~<�0<��<�<R��;om�;��;���;<��;qP�;�,�;��;��;��;�8�;�b�;���;��;]C�;���;!+�;��;�U�;��;�Ç;��;��z;��p;y�f;��\;�<S;w�I;.)@;~�6;)�-;~w$;�y;}�;N�	;�0;�K�:Mo�:���:XT�:(�:��:)�:%�~:y�_:7JA:�":��:[��9��9Qu39K��8��F�ק"��O��E���]����/�<2�M�?�g�3���<��2I��@���!������z�κfZۺP������~ �Ĵ�8�����4�kS�{m%��+���1�#�7�̩=���C�)�I�r�O�C�U��[�Y�a��g��m��s���y��|�8���Ǵ������R����������m���o���棚��  �  .l=�=?�=jJ=a�=�=�&=�� =~b =  =N:�<�s�<���<|��<��<�Q�<ǆ�<պ�<���<��<�P�<#��<[��<C��<��<�0�<|Y�<k��<¥�<o��<T��<a�<�)�<�E�<�_�< x�<��<���<ڲ�<���<1��<��<B��<���<���<V��<>��< ��<���<���<Ѱ�<ڜ�<k��<�j�<0L�<)*�<y�<��<ԭ�<�|�<�G�<��<��<<��<PL�<O�<;��<e�<��<I��<�X�<��<G��<h'�<���<�G�<�Ѻ<�W�<�ٷ<KX�<�Ҵ<�I�<ټ�<k,�<}��<-�<if�<^ȩ<4'�<�<�ۤ<�1�<���<�ԟ<�"�<	n�<<���<�A�<i��<�ē<k�<J@�<z{�<;��<~�<�$�<SZ�<��<�<���<�'�<̲|<�y<�uu<X�q<d6n<+�j<�f<#Vc<Ŷ_<\<zX<R�T<�AQ<ܧM<�J<�yF<l�B<�S?<��;<�88<��4<�)1<M�-<�(*<Э&<S7#<�<_W<m�<��<�+<p�<�~<�0<��<��<��;Qm�;5�;���;Q��;SP�;*-�;��;��;��;�8�;�b�;\��;��;MC�;߮�;4+�;A��;�U�;��;ć;Q��;��z;�p;k�f;��\;�<S;��I;)@;��6;��-;�w$;�y;��;��	;40;�K�:�n�:���:�S�:��:��:�'�:`�~:?�_:�LA:��":]�:n��97�9�}39���8��F�i�"�fQ��[�������:.��<2�OM�ռg����;��?H��?@���"��;����κ�Zۺ���:����~ �S�����	��4�wS��m%��+���1��7��=�o�C�]�I�γO��U�s�[��a�:�g��m���s�\�y�[|�I�������.���L�����������U���j���ƣ���  �  -l=�=3�=oJ=b�=�=�&=�� =�b =���<Q:�<�s�<���<}��<��<�Q�<���<��<���<��<�P�<��<l��<G��<��<�0�<dY�<`��<���<n��<H��<m�<�)�<�E�<�_�<�w�<���<z��<ز�<���<,��<��<<��<���<v��<e��<=��<0��<���<|��<ܰ�<ќ�<{��<�j�<*L�< *�<p�<
��<ϭ�<�|�<�G�<��<��<>��<aL�<P�<G��<e�<��<B��<�X�<��<>��<i'�<i��<�G�<�Ѻ<�W�<�ٷ<6X�<�Ҵ<�I�<ؼ�<f,�<s��<�<_f�<iȩ<5'�<��<�ۤ<�1�<���<�ԟ<�"�<�m�<춚<���<�A�<`��<�ē<r�<>@�<�{�<.��<��<�$�<TZ�<��<�<���<�'�<ʲ|<�y<�uu<E�q<I6n<R�j<��f<JVc<��_<�\<%zX<@�T<�AQ<קM<�J<eyF<��B<�S?<��;<�88<k�4<�)1<=�-<�(*<�&<>7#<�<MW<i�<p�<�+<n�<�~<�0<��<�<&��;vm�;%�;���;(��;CP�;#-�;��;�;P�;�8�;-c�;V��;K�;�B�;ծ�;+�;0��;�U�;s�;�Ç;���;f�z;�p;��f;��\;o<S;�I;�(@;�6;��-;�w$;|y;I�;��	;0;�L�:zn�:S��:�S�:��:��:�'�:��~:��_:�JA:��":��:���9��9f~39x��8��F���"�+N��K��� ����,�J>2�{M��g����p<���H���?���"��7�����κ&Zۺ<��m����} �������K��4��S��m%���+��1���7�y�=���C� �I�ʳO��U�7�[�b�a�L�g��m���s�)�y��|����g���_�������먎�8���)�������ʣ���  �  5l=�=7�=mJ=b�=�=�&=�� =�b =���<C:�<�s�<���<���<��<�Q�<ņ�<ݺ�<���<��<�P�<��<W��<<��<��<�0�<mY�<r��<˥�<p��<J��<h�<�)�<�E�<�_�<�w�<��<���<޲�<���<,��<��<O��<���<~��<]��<:��<��<���<~��<԰�<Ϝ�<j��<�j�<,L�<**�<z�<��<ӭ�<�|�<�G�<��<��<7��<JL�<K�<A��<e�<��<V��<�X�<��<?��<m'�<x��<�G�<�Ѻ<�W�<�ٷ<CX�<�Ҵ<�I�<ټ�<q,�<���< �<bf�<gȩ<.'�<<�ۤ<�1�<���<�ԟ<�"�<n�<�<���<B�<d��<�ē<b�<<@�<�{�<3��<~�<{$�<SZ�<��<�<���<�'�<ֲ|<�y<�uu<Z�q<U6n<A�j<��f<>Vc<��_<\<zX<@�T<�AQ<��M<�J<wyF<w�B<�S?<��;<�88<{�4<�)1<8�-<�(*<ޭ&<K7#<�<_W<x�<��<�+<[�<�~<�0<��<�<���;sm�;"�;���;n��;uP�;--�;��;�;��;�8�;c�;E��;%�;C�;ﮢ;+�;.��;V�;��;ć;��;(�z;��p;<�f;z�\;}<S;��I;�(@;��6;��-;�w$;�y;��;��	;)0;�K�:1n�:���:�S�:x�::�:�'�:+�~:��_:�KA:e�":��:���9�9}�39��8�F�	�"��P��w�������`-�6>2�LM�(�g�b���;���H���?��P#�������κ;Zۺ~������p~ �f������v4��S��m%�2�+�,�1� 7�N�=�r�C���I�гO���U���[���a�Šg���m���s�M�y�O|�h�������]������Ҩ��	���>������������  �  7k=�
=�=�H=��=/�=i$=[� =�_ =���<^4�<~m�<̥�<=��<��<lI�<$~�<���<K��<��<�E�<�t�<���<���<���<h#�<PK�<�q�<|��<���<���<.��<��<<3�<�L�<2d�<Zy�<Q��<��<��<��<��<���<G��<k��<���<���<���<��<���<���<~�<
f�<�J�<�+�<	�<���<���<i��<�Y�<�$�<T��<1��<m�< (�<���<���<e@�<���<���<4�<���<�l�<M�<���<$�<���<5�<���<�6�<���< )�<<&�<�y�<6�<YI�<��<��<bh�<¤<��<�l�<��<��<	Y�<բ�<��<�/�<Us�<Ѵ�<c��<U2�<n�<R��<��<��<�Q�<W��<4��<��<V#�<٫|<�y<su<��q<�7n<��j<��f<�]c<��_<�#\<�X<��T<)TQ<A�M<&J<�F< C<�p?<��;<�Y8<��4<�N1<f�-<�Q*<�&<kd#<�<{�<\!<x�<�b<<�<�l<�&<��<�Y�;���;˙�;�M�;f�;2��;���;���;���;a��;5Կ;A �;(<�;凮;"�;�P�;�͝;V[�;:��;᧍;�f�;$7�;�.|;�r;h;�5^;6yT;;�J;�_A;�8;��.;��%;��;
�;��
;�I;s�:܋�:��:�Y�:��:���:]�:+Q�:��c:��D:�`&:�J:��9a �9��?9/'�84e����O���������������/���J��e�r��I?��dT��"V��uA�������ͺ�ں#9�;��( �sc����V�������!/%�fH+�w\1��m7��y=�C�C�p�I�T�O�ЎU���[�ԋa�G�g��m��{s��uy��n�������������6���F���ا��������������  �  :k=�
=�=�H=��=)�=d$=W� =�_ =���<^4�<zm�<ĥ�<=��<��<qI�<~�<���<B��<��<�E�<�t�<���<���<���<j#�<aK�<�q�<{��<���<���<8��<��<N3�<�L�<%d�<ky�<Z��<���<��<۶�<���<���<d��<e��<���<���<��<��<��<���<~�<f�<�J�<�+�<	�<���<���<Y��<�Y�<�$�<]��<>��<m�<�'�<���<���<`@�<��<���<4�<���<�l�<_�<���<$�<v��<5�<���<�6�<���<)�<圱<"�<�y�<M�<XI�<"��<��<Yh�<���<��<�l�<��<��<�X�<ܢ�<{�<�/�<Ps�<ʴ�<g��<Q2�<�n�<O��<��<��<�Q�<]��<1��</��<\#�<��|<�y<su<��q<�7n<יj<��f<^c<��_<$\<#�X<w�T<TQ<K�M<G&J<�F<  C<�p?<��;<zY8<s�4<�N1<b�-<�Q*<��&<[d#<�<e�<f!<]�<�b<<�<�l<�&<��<�Y�;��;ә�;8N�;��;-��;i��;���;ī�;g��;}Կ;S �;�;�;)��;I�;�P�;�͝;&[�;��;��;Gg�;7�;�.|;Wr;�h;�5^;cyT;��J;�_A;�8;;�.;̢%;Ƞ;�;+�
;I;>s�:%��:���:�Z�:��:���:��:�Q�:�c:\�D:�b&:"J:�9��9ڝ?9�.�8�@����_���������2��
�/���J���e�
���=��iT���U��<B��Z��6�ͺ�ں9����( ��c�c����������V/%�HH+��\1�m7��y=�v�C�׉I�b�O���U���[���a��g�Z�m�|s��uy�_n�ó��v���ĭ���������ϧ������F���*����  �  6k=�
=ک=�H=��=,�=m$=U� =�_ =|��<c4�<m�<ʥ�<D��<��<~I�<~�<Ʊ�<D��<��<�E�<�t�<���<���<���<_#�<UK�<�q�<y��<���<���<@��<��<I3�<�L�<'d�<iy�<D��<���<��<��<��<���<[��<R��<���<���<���<��<���<���<~�<f�<�J�<�+�<	�<���<��<S��<�Y�<�$�<`��<<��<m�<(�<���<���<L@�<��<���< 4�<���<�l�<]�<���<$�<y��<5�<���<�6�<���<)�<�<!�<�y�<B�<II�<(��<��<jh�<���<��<�l�<��<��<�X�<袚<t�<�/�<Ys�<̴�<p��<D2�<�n�<L��<��<��<�Q�<b��< ��<&��<T#�<׫|<�y<su<��q<�7n<ڙj<��f<^c<��_<�#\<1�X<��T<'TQ<=�M<2&J<��F< C<�p?<��;<�Y8<h�4<�N1<J�-<�Q*<	�&<gd#<,�<X�<�!<\�<�b<<�<�l<�&<��<�Y�;��;���;	N�;��;$��;���;���;��;#��;gԿ;] �;�;�; ��;��;�P�;�͝;N[�;B��;ӧ�;&g�;�6�;�.|;kr;&h;
6^;LyT;��J;a_A;^8;�.;%�%;��;�;��
;�H;At�:��:���:�Z�:��:���:��:#R�:��c:F�D:�`&:UK:��9��9��?9Y�8�A����Z�������1�����O�/�q�J���e�����>��aU��GU��&B��7��A�ͺ�ںH9����,( �
d� ����������I/%�H+��\1� m7�z=��C���I�L�O�w�U�@�[�*�a�Y�g��m��{s�vuy��n����p��������?�����������2��������  �  9k=�
=�=�H=��='�=f$=X� =�_ =���<_4�<wm�<˥�<?��<��<uI�<~�<���<E��<��<�E�<�t�<���<���<���<h#�<dK�<�q�<|��<���<���<:��<��<H3�<�L�<5d�<^y�<S��<���<��<ڶ�<��<���<\��<i��<���<���<��<	��<���<���<~�<f�<�J�<�+�<	�<���<���<V��<�Y�<�$�<b��<7��<m�<�'�<���<���<a@�<��<���< 4�<���<�l�<[�<���<$�<���<5�<���<�6�<���<)�<朱<%�<�y�<M�<VI�<"��<��<\h�<���<��<�l�<��<��<�X�<ߢ�<{�<�/�<Ys�<Ŵ�<g��<L2�<�n�<R��<��<��<�Q�<`��<7��<��<X#�<ҫ|<�y<su<��q<�7n<��j<��f<�]c<��_<$\<,�X<v�T<TQ<G�M<'&J<"�F<% C<�p?<��;<�Y8<x�4<�N1<]�-<�Q*<��&<jd#<!�<i�<m!<e�<�b<
<$�<�l<�&<��<pY�;��;ʙ�;DN�;��;0��;y��;���;ͫ�;X��;cԿ;D �;7<�;�;-�;�P�;�͝;![�;D��;٧�;)g�;7�;�.|;&r;�h;�5^;CyT;��J;�_A;�8;�.;��%;��;��;B�
;�H;@s�:T��:���:@Z�:��:���:>�:�Q�:.�c:��D:�`&:bK:��9��9r�?9�*�8`U����s������V��m���/���J�=�e����=���T���U���B���� �ͺt�ں�8纨��( ��c�I����������}/%�GH+��\1�/m7��y=�|�C��I���O���U���[�\�a�6�g��m�(|s�tuy�Vn�泂���������%���)���ԧ������H�������  �  >k=�
=�=�H=��=/�=f$=Z� =�_ =���<a4�<|m�<Υ�<9��<��<kI�<%~�<���<G��<��<�E�<�t�<���< ��<���<^#�<[K�<�q�<���<���<���</��<��<K3�<�L�<5d�<Wy�<\��<��<*��<ֶ�<��<���<V��<_��<���<���<���<��<���<���<~�<f�<�J�<�+�<	�<���<���<f��<�Y�<�$�<Z��<7��<m�<�'�<���<���<V@�<���<���< 4�<���< m�<K�<���<$�<���<5�<���<�6�<���<")�<���<,�<�y�<F�<MI�<&��<��<\h�<¤<��<�l�<��<��<Y�<֢�<��<�/�<Ys�<ϴ�<g��<U2�<�n�<U��<��<��<�Q�<T��</��<��<b#�<ī|<�y<su<��q<�7n<��j<��f<�]c<��_<�#\<'�X<~�T<TQ<[�M<!&J<�F<
 C<�p?<��;<Y8<��4<�N1<k�-<�Q*<�&<qd#<�<w�<Z!<y�<�b<<$�<�l<�&<��<�Y�;'��;���;"N�;��;W��;Z��;���;���;O��;pԿ;1 �;5<�;ه�;P�;�P�;�͝;[�;4��;���;g�;�6�;~.|;�r;�h;6^;FyT;l�J;�_A;�8;��.;�%;��;�;�
;kI;�r�:���:t��:IZ�:�:0��:��:gQ�:щc:��D:�a&:mK:��9�"�9��?9Q1�8�b�������槻�?������/���J�U�e����N>��U��mU��_A������ͺʕں�8����( �uc����>������2/%�FH+�r\1��m7��y=�Z�C�p�I��O��U�ʍ[�y�a��g�=�m�|s�cuy��n�������������>��������������7���.����  �  7k=�
=�=�H=��=(�=k$=W� =�_ =���<b4�<ym�<ɥ�<@��<��<tI�<~�<���<J��<��<�E�<�t�<���<���<���<e#�<eK�<�q�<��<���<���<;��<��<M3�<�L�<)d�<`y�<T��<��<)��<۶�<��<���<a��<b��<���<���<��<��<���<���<~�<f�<�J�<�+�<	�<���< ��<V��<�Y�<�$�<_��<8��<m�<�'�<���<���<Z@�<��<���<#4�<���<�l�<P�<���<$�<z��<5�<���<�6�<���<)�<朱<'�<�y�<Q�<SI�<��<��<ch�<���<��<�l�<��<��<�X�<ޢ�<��<�/�<Ws�<Ǵ�<h��<P2�<�n�<N��<��<��<�Q�<b��<3��<$��<R#�<׫|<�y<su<��q<�7n<ęj<��f<�]c<��_<�#\<5�X<�T<$TQ<>�M<-&J<�F< C<�p?<��;<�Y8<q�4<�N1<]�-<�Q*<��&<gd#<#�<p�<m!<d�<�b<<�<�l<�&<��<�Y�;���;�;JN�;��;<��;��;���;ҫ�;>��;|Կ;A �;<�;���;2�;�P�;�͝;%[�;G��;̧�;=g�;�6�;�.|;>r;�h;
6^;0yT;��J;�_A;�8;$�.;�%;ʠ;"�;I�
;�H;s�:���:���:LZ�: �:��:m�:�Q�:a�c:��D:�`&:�K:��9�!�9'�?9�(�8�Q������������������/���J�ۗe�#���=���T���U��{B������ͺH�ں�8�C��( ��c�M��U�������k/%�BH+��\1�m7�z=��C��I�y�O�w�U���[�;�a�j�g��m��{s�Muy��n�ҳ����������������
���~���6��������  �  2k=�
=ީ=�H=��=)�=k$=S� =�_ =y��<c4�<zm�<˥�<H��<��<�I�<~�<���<D��<��<�E�<�t�<���<���<���<_#�<]K�<�q�<v��<���<���<;��<��<M3�<�L�<'d�<ly�<N��<��<��<׶�<��<��<g��<X��<���<���<���<��<���<���<~�<f�<�J�<�+�<	�<���<��<V��<�Y�<�$�<^��<9��<m�<(�<���<���<Q@�<��<���<!4�<���<�l�<V�<���<$�<y��<5�<���<�6�<���<)�<뜱< �<�y�<M�<KI�<"��<��<mh�<���<��<�l�<��<��<�X�<뢚<w�<�/�<\s�<Ǵ�<n��<B2�<�n�<I��<��<��<�Q�<[��<'��<.��<K#�<�|<�y<su<��q<�7n<ՙj<��f<^c<��_<�#\<*�X<c�T<6TQ<-�M<?&J<�F< C<�p?<��;<�Y8<b�4<�N1<D�-<�Q*<��&<jd#<2�<[�<�!<c�<�b<	<�<m<�&<��<}Y�;���;���;+N�;��;��;���;c��;Ы�;2��;{Կ;K �;�;�;-��;�;�P�;�͝;[�;T��;���;Vg�;�6�;�.|;*r;h;�5^;.yT;��J;Y_A;(8;�.;E�%; ;�;��
;�H;�s�:��:���:aZ�:��:���:E�:�Q�:=�c:��D:`&:|K:b�9��9t�?9V#�8�=�y��5���������@��-�/��J�ǘe�����=��5U���U���B������ͺ˔ںB9线��( ��c���������v�m/%�H+�
]1��l7�0z=�4�C���I�z�O���U��[��a���g���m�\|s��uy��n��z���ǭ������-�����������n���۩���  �  6k=�
=ݩ=�H=��=.�=g$=W� =�_ =���<h4�<wm�<ϥ�<C��<��<vI�<!~�<���<M��<��<�E�<�t�<���<���<���<a#�<UK�<�q�<{��<���<���<3��<��<G3�<�L�<0d�<^y�<M��<��<'��<ڶ�<��<���<]��<Z��<���<���<���<��< ��<���<~�<f�<�J�<�+�<	�<���<��<[��<�Y�<�$�<_��<=��<m�<(�<���<���<S@�<��<���<4�<���<�l�<L�<���<$�<~��<5�<���<�6�<���<)�<眱<!�<�y�<B�<NI�<%��<��<eh�<���<��<�l�<��<��<Y�<࢚<z�<�/�<]s�<ȴ�<p��<N2�<�n�<R��<��<��<�Q�<X��<(��<(��<T#�<ϫ|<�y<su<��q<�7n<��j<��f<�]c<��_<�#\<+�X<y�T<TQ<=�M<:&J<�F< C<�p?<��;<�Y8<u�4<�N1<`�-<�Q*<��&<qd#<)�<b�<q!<r�<b<< �<�l<�&<��<�Y�;��;���;N�;��;+��;~��;���;���;6��;`Կ;9 �;%<�;���;�;�P�;�͝;#[�;<��;ק�;,g�;�6�;�.|;jr;4h;�5^;^yT;��J;�_A;8;>�.;%�%;��;�;b�
;I;Ss�:���:���:�Z�:��:���:��:�Q�:��c:[�D:a&:(K:��9�!�9?�?9�"�8W����n���٧��v��n��#�/���J���e�����>��U��{U���A�����L�ͺ�ں�8� ���( ��c�A��������n�c/%��G+��\1�m7��y=�`�C�t�I�S�O�ÎU���[��a�V�g��m�|s�auy��n�쳂������������0�����������A�������  �  :k=�
=�=�H=��=+�=e$=^� =�_ =���<_4�<{m�<ҥ�<9��<��<mI�<&~�<���<L��<��<�E�<�t�<���<���<���<p#�<dK�<�q�<���<|��<���<2��<��<H3�<�L�<3d�<Wy�<\��<��<$��<ٶ�<���<���<X��<m��<���<���<��<��<��<���<~�<f�<�J�<�+�<	�<���<���<c��<�Y�<�$�<[��<<��<m�<�'�<���<���<f@�<��<���<4�<���<�l�<I�<���<$�<��<�4�<���<�6�<���<)�<ݜ�<&�<�y�<L�<]I�<��<��<[h�<¤<��<�l�<��<��<	Y�<֢�<��<�/�<]s�<̴�<e��<S2�<�n�<[��<��<��<�Q�<g��<9��<��<[#�<��|<�y<su<��q<�7n<��j<��f<�]c<��_<�#\<(�X<��T<TQ<L�M<$&J<!�F<2 C<p?<��;<}Y8<��4<�N1<d�-<�Q*< �&<xd#<�<{�<_!<|�<�b<<�<�l<�&<��<�Y�;���;��;EN�;��;C��;L��;���;���;Y��;eԿ;* �;0<�;ۇ�;S�;�P�;�͝; [�;��;맍;g�;,7�;�.|;<r;�h;�5^;oyT;��J;`A;�8;x�.;�%;Š;"�;"�
;YI;�r�:��:���:�Z�:�:���:�:�Q�:�c:^�D:Ga&:�J:��9x!�9В?9r3�8�b�{�����`����������/���J�
�e�����=��T��:V��B��1��w�ͺs�ں,9����( �rc����,�����p�C/%�[H+��\1�am7��y=�e�C���I���O�L�U�{�[�m�a��g�e�m��{s�zuy��n�ų��Ȱ������A��������������#���>����  �  8k=�
=۩=�H=��=0�=f$=Y� =�_ =���<d4�<�m�<˥�<>��<��<tI�<~�<Ʊ�<F��<��<�E�<�t�<���<���<���<^#�<VK�<�q�<~��<���<���<4��<��<H3�<�L�<*d�<_y�<O��<��<!��<߶�<��<���<W��<V��<���<���<���<��<���<���<~�<f�<�J�<�+�<	�<���< ��<^��<�Y�<�$�<^��<:��<m�<�'�<���<���<P@�<��<���<4�<���<�l�<O�<���<$�<y��<�4�<���<�6�<���<)�<眱<%�<�y�<B�<JI�<"��<��<`h�<���<��<�l�<��<��<�X�<ܢ�<��<�/�<Xs�<д�<n��<M2�<�n�<Q��<��<��<�Q�<\��<$��< ��<U#�<˫|<�y<su<��q<�7n<��j<��f<�]c<��_<�#\<#�X<|�T<TQ<C�M<(&J<��F< C<�p?<��;<�Y8<z�4<�N1<Y�-<�Q*<�&<jd#< �<~�<l!<i�<�b<<�<�l<�&<��<�Y�;��;���;N�;s�;8��;u��;���;���;.��;gԿ;9 �;<�;���;�;�P�;�͝;6[�;0��;֧�;g�;�6�;�.|;�r;h;�5^;FyT;��J;�_A;*8;k�.;��%;�;>�;M�
;4I;�s�:)��:���:pZ�:��:l��:'�:�Q�:�c:%�D:}`&:�J:��9@ �9�?9�#�8>W�~��0���������*����/���J�+�e�T���>��FU���U���A������ͺ�ں�8线��J( ��c�[��*�������#/%�H+��\1�m7��y=�_�C�l�I�<�O���U� �[�U�a�L�g�"�m��{s��uy��n�곂���������"���+����������;�������  �  4k=�
=�=�H=��=%�=i$=W� =�_ =���<h4�<xm�<ǥ�<K��<��<�I�<~�<���<D��<��<�E�<�t�<���<���<���<f#�<aK�<�q�<y��<���<���<>��<��<J3�<�L�<#d�<hy�<I��<���<��<׶�<��<���<e��<_��<���<���<��<��<���<���<~�<f�<�J�<�+�<	�<���<	��<L��<�Y�<�$�<j��<8��<m�<�'�<���<���<X@�<��<���<!4�<���<�l�<`�<���<$�<u��<�4�<���<�6�<���<)�<眱<$�<�y�<N�<SI�<)��<��<bh�<���<��<�l�<���<��<�X�<颚<v�<�/�<Ws�<Ĵ�<s��<N2�<�n�<M��<��<��<�Q�<`��</��<.��<N#�<ݫ|<�y<su<��q<�7n<ҙj<��f<�]c<��_<�#\<(�X<h�T<)TQ<3�M<C&J<�F<  C<�p?<��;<�Y8<s�4<�N1<b�-<�Q*<��&<cd#<:�<\�<�!<W�<�b<	<.�<�l<�&<��<^Y�; ��;Ǚ�;9N�;��;&��;���;f��;ܫ�;A��;nԿ;B �;�;�;��;�;�P�;�͝;[�;H��;ӧ�;Ng�;�6�;�.|;r;�h;�5^;.yT;��J;�_A;N8;��.;3�%;ڠ;�;��
;�H;t�:���:s��:[Z�:��: ��:�
�:$R�:%�c:��D:�`&:�K:��9��9^�?9	 �8�E�K���������_�����/���J�B�e�����=���T��/U��
C�����/�ͺ'�ںE8����_( �&d�������������/%��G+��\1��l7�z=�F�C���I�{�O���U�ʍ[��a���g�فm�R|s��uy�Xn���������ɭ�����4���ߧ������b��������  �  6k=�
=ީ=�H=��=,�=n$=Y� =�_ =���<_4�<�m�<ѥ�<H��<��<�I�<%~�<ı�<A��<��<�E�<�t�<���<���<���<d#�<WK�<�q�<|��<���<���<4��<��<@3�<�L�<+d�<\y�<L��<��<��<ض�<	��<���<S��<^��<���<���<���<��<���<���<~�<f�<�J�<�+�<	�<���<	��<a��<�Y�<�$�<_��<1��<&m�< (�<���<���<W@�<���<���<#4�<���<�l�<O�<���<$�<{��<5�<���<�6�<���<)�<䜱<'�<�y�<A�<QI�<"��<��<jh�<¤<��<�l�< ��<��<Y�<뢚<u�<�/�<_s�<մ�<j��<L2�<�n�<Q��<��<��<�Q�<]��<+��<��<T#�<٫|<�y<su<��q<�7n<��j<��f<�]c<��_<�#\<!�X<~�T<#TQ<=�M<&J<�F< C<�p?<��;<�Y8<|�4<�N1<Y�-<�Q*<�&<wd#<3�<Z�<�!<{�<�b<<�<�l<�&<��<�Y�;��;���;N�;z�;3��;{��;���;���;A��;FԿ;> �;<�;���;�;�P�;�͝;[�;K��;̧�;g�;�6�;�.|;�r;h;d6^;$yT;��J;�_A;@8;w�.;?�%;��;�;��
;GI;#t�:8��:���:�Y�:��:���::�:�Q�:
�c:|�D:`&:�K:v�95�9�?9*%�8]�4��c����������V����/���J�ϗe�a���>���T���U���A��1��s�ͺ�ں�8����7( �|c���������`�/%�1H+��\1�@m7��y=�܂C���I�5�O���U��[���a�\�g��m�|s��uy��n�������������.���F�����������7��� ����  �  ;k=�
=�=�H=��=)�=a$=X� =�_ =���<Z4�<�m�<¥�<;��<��<qI�<~�<���<A��<��<�E�<�t�<���<���<���<g#�<dK�<�q�<}��<u��<���</��<��<C3�<�L�</d�<Uy�<]��<��<(��<ն�<���<���<^��<k��<���<���<��<��<���<���<~�<f�<�J�<�+�<	�<���<���<[��<�Y�<�$�<i��<6��<m�<�'�<���<���<c@�<
��<���<4�<���<�l�<L�<���<$�<|��<5�<���<�6�<���< )�<ל�<$�<�y�<N�<WI�<��<��<Lh�< ¤<��<�l�<��<��<�X�<ڢ�<��<�/�<Ls�<Ӵ�<a��<[2�<�n�<P��<��<��<�Q�<X��<7��<%��<\#�<��|<�y<su<��q<�7n<��j<��f<�]c<��_<�#\<'�X<��T<�SQ<Q�M<3&J<�F< C<�p?<��;<nY8<v�4<�N1<z�-<�Q*<�&<Xd#<�<s�<e!<e�<�b<<7�<�l<�&<q�<�Y�;���;ș�;FN�;��;3��;2��;���;���;f��;TԿ;C �;<�;Ӈ�;T�;�P�;�͝;[�;
��;觍;2g�;%7�;�.|;�r;Kh;�5^;HyT;��J;�_A;�8;Z�.;��%;�;H�;�
;I;s�:s��:m��:;Z�:��:��:v�:#Q�:��c:D�D:�`&:�I:�
�9*"�9��?95�8�j����{�������e�������/���J�5�e����=���T��0V���A������ͺ3�ں#8����( ��c�m��U�������/%�zH+�D\1��l7��y=���C���I�J�O�ƎU���[�2�a��g���m�|s�`uy��n�̳����������/������六�����0���Y����  �  6k=�
=ީ=�H=��=,�=n$=Y� =�_ =���<_4�<�m�<ѥ�<H��<��<�I�<%~�<ı�<A��<��<�E�<�t�<���<���<���<d#�<WK�<�q�<|��<���<���<4��<��<@3�<�L�<+d�<\y�<L��<��<��<ض�<	��<���<S��<^��<���<���<���<��<���<���<~�<f�<�J�<�+�<	�<���<	��<a��<�Y�<�$�<_��<1��<&m�< (�<���<���<W@�<���<���<#4�<���<�l�<O�<���<$�<{��<5�<���<�6�<���<)�<䜱<'�<�y�<A�<QI�<"��<��<jh�<¤<��<�l�< ��<��<Y�<뢚<u�<�/�<_s�<մ�<j��<L2�<�n�<Q��<��<��<�Q�<]��<+��<��<T#�<٫|<�y<su<��q<�7n<��j<��f<�]c<��_<�#\<!�X<~�T<#TQ<=�M<&J<�F< C<�p?<��;<�Y8<|�4<�N1<Y�-<�Q*<�&<wd#<3�<Z�<�!<{�<�b<<�<�l<�&<��<�Y�;��;���;N�;z�;3��;{��;���;���;A��;FԿ;> �;<�;���;�;�P�;�͝;[�;K��;̧�;g�;�6�;�.|;�r;h;d6^;$yT;��J;�_A;@8;w�.;?�%;��;�;��
;GI;#t�:8��:���:�Y�:��:���::�:�Q�:
�c:|�D:`&:�K:v�95�9�?9*%�8]�4��c����������V����/���J�ϗe�a���>���T���U���A��1��s�ͺ�ں�8����7( �|c���������`�/%�1H+��\1�@m7��y=�܂C���I�5�O���U��[���a�\�g��m�|s��uy��n�������������.���F�����������7��� ����  �  4k=�
=�=�H=��=%�=i$=W� =�_ =���<h4�<xm�<ǥ�<K��<��<�I�<~�<���<D��<��<�E�<�t�<���<���<���<f#�<aK�<�q�<y��<���<���<>��<��<J3�<�L�<#d�<hy�<I��<���<��<׶�<��<���<e��<_��<���<���<��<��<���<���<~�<f�<�J�<�+�<	�<���<	��<L��<�Y�<�$�<j��<8��<m�<�'�<���<���<X@�<��<���<!4�<���<�l�<`�<���<$�<u��<�4�<���<�6�<���<)�<眱<$�<�y�<N�<SI�<)��<��<bh�<���<��<�l�<���<��<�X�<颚<v�<�/�<Ws�<Ĵ�<s��<N2�<�n�<M��<��<��<�Q�<`��</��<.��<N#�<ݫ|<�y<su<��q<�7n<ҙj<��f<�]c<��_<�#\<(�X<h�T<)TQ<3�M<C&J<�F<  C<�p?<��;<�Y8<s�4<�N1<b�-<�Q*<��&<cd#<:�<\�<�!<W�<�b<	<.�<�l<�&<��<^Y�; ��;Ǚ�;9N�;��;&��;���;f��;ܫ�;A��;nԿ;B �;�;�;��;�;�P�;�͝;[�;H��;ӧ�;Ng�;�6�;�.|;r;�h;�5^;.yT;��J;�_A;N8;��.;3�%;ڠ;�;��
;�H;t�:���:s��:[Z�:��: ��:�
�:$R�:%�c:��D:�`&:�K:��9��9^�?9	 �8�E�K���������_�����/���J�B�e�����=���T��/U��
C�����/�ͺ'�ںE8����_( �&d�������������/%��G+��\1��l7�z=�F�C���I�{�O���U�ʍ[��a���g�فm�R|s��uy�Xn���������ɭ�����4���ߧ������b��������  �  8k=�
=۩=�H=��=0�=f$=Y� =�_ =���<d4�<�m�<˥�<>��<��<tI�<~�<Ʊ�<F��<��<�E�<�t�<���<���<���<^#�<VK�<�q�<~��<���<���<4��<��<H3�<�L�<*d�<_y�<O��<��<!��<߶�<��<���<W��<V��<���<���<���<��<���<���<~�<f�<�J�<�+�<	�<���< ��<^��<�Y�<�$�<^��<:��<m�<�'�<���<���<P@�<��<���<4�<���<�l�<O�<���<$�<y��<�4�<���<�6�<���<)�<眱<%�<�y�<B�<JI�<"��<��<`h�<���<��<�l�<��<��<�X�<ܢ�<��<�/�<Xs�<д�<n��<M2�<�n�<Q��<��<��<�Q�<\��<$��< ��<U#�<˫|<�y<su<��q<�7n<��j<��f<�]c<��_<�#\<#�X<|�T<TQ<C�M<(&J<��F< C<�p?<��;<�Y8<z�4<�N1<Y�-<�Q*<�&<jd#< �<~�<l!<i�<�b<<�<�l<�&<��<�Y�;��;���;N�;s�;8��;u��;���;���;.��;gԿ;9 �;<�;���;�;�P�;�͝;6[�;0��;֧�;g�;�6�;�.|;�r;h;�5^;FyT;��J;�_A;*8;k�.;��%;�;>�;M�
;4I;�s�:)��:���:pZ�:��:l��:'�:�Q�:�c:%�D:}`&:�J:��9@ �9�?9�#�8>W�~��0���������*����/���J�+�e�T���>��FU���U���A������ͺ�ں�8线��J( ��c�[��*�������#/%�H+��\1�m7��y=�_�C�l�I�<�O���U� �[�U�a�L�g�"�m��{s��uy��n�곂���������"���+����������;�������  �  :k=�
=�=�H=��=+�=e$=^� =�_ =���<_4�<{m�<ҥ�<9��<��<mI�<&~�<���<L��<��<�E�<�t�<���<���<���<p#�<dK�<�q�<���<|��<���<2��<��<H3�<�L�<3d�<Wy�<\��<��<$��<ٶ�<���<���<X��<m��<���<���<��<��<��<���<~�<f�<�J�<�+�<	�<���<���<c��<�Y�<�$�<[��<<��<m�<�'�<���<���<f@�<��<���<4�<���<�l�<I�<���<$�<��<�4�<���<�6�<���<)�<ݜ�<&�<�y�<L�<]I�<��<��<[h�<¤<��<�l�<��<��<	Y�<֢�<��<�/�<]s�<̴�<e��<S2�<�n�<[��<��<��<�Q�<g��<9��<��<[#�<��|<�y<su<��q<�7n<��j<��f<�]c<��_<�#\<(�X<��T<TQ<L�M<$&J<!�F<2 C<p?<��;<}Y8<��4<�N1<d�-<�Q*< �&<xd#<�<{�<_!<|�<�b<<�<�l<�&<��<�Y�;���;��;EN�;��;C��;L��;���;���;Y��;eԿ;* �;0<�;ۇ�;S�;�P�;�͝; [�;��;맍;g�;,7�;�.|;<r;�h;�5^;oyT;��J;`A;�8;x�.;�%;Š;"�;"�
;YI;�r�:��:���:�Z�:�:���:�:�Q�:�c:^�D:Ga&:�J:��9x!�9В?9r3�8�b�{�����`����������/���J�
�e�����=��T��:V��B��1��w�ͺs�ں,9����( �rc����,�����p�C/%�[H+��\1�am7��y=�e�C���I���O�L�U�{�[�m�a��g�e�m��{s�zuy��n�ų��Ȱ������A��������������#���>����  �  6k=�
=ݩ=�H=��=.�=g$=W� =�_ =���<h4�<wm�<ϥ�<C��<��<vI�<!~�<���<M��<��<�E�<�t�<���<���<���<a#�<UK�<�q�<{��<���<���<3��<��<G3�<�L�<0d�<^y�<M��<��<'��<ڶ�<��<���<]��<Z��<���<���<���<��< ��<���<~�<f�<�J�<�+�<	�<���<��<[��<�Y�<�$�<_��<=��<m�<(�<���<���<S@�<��<���<4�<���<�l�<L�<���<$�<~��<5�<���<�6�<���<)�<眱<!�<�y�<B�<NI�<%��<��<eh�<���<��<�l�<��<��<Y�<࢚<z�<�/�<]s�<ȴ�<p��<N2�<�n�<R��<��<��<�Q�<X��<(��<(��<T#�<ϫ|<�y<su<��q<�7n<��j<��f<�]c<��_<�#\<+�X<y�T<TQ<=�M<:&J<�F< C<�p?<��;<�Y8<u�4<�N1<`�-<�Q*<��&<qd#<)�<b�<q!<r�<b<< �<�l<�&<��<�Y�;��;���;N�;��;+��;~��;���;���;6��;`Կ;9 �;%<�;���;�;�P�;�͝;#[�;<��;ק�;+g�;�6�;�.|;jr;4h;�5^;^yT;��J;�_A;8;>�.;%�%;��;�;b�
;I;Ss�:���:���:�Z�:��:���:��:�Q�:��c:[�D:a&:(K:��9�!�9?�?9�"�8W����n���٧��v��n��#�/���J���e�����>��U��{U���A�����L�ͺ�ں�8� ���( ��c�A��������n�c/%��G+��\1�m7��y=�`�C�t�I�S�O�ÎU���[��a�V�g��m�|s�auy��n�쳂������������0�����������A�������  �  2k=�
=ީ=�H=��=)�=k$=S� =�_ =y��<c4�<zm�<˥�<H��<��<�I�<~�<���<D��<��<�E�<�t�<���<���<���<_#�<]K�<�q�<v��<���<���<;��<��<M3�<�L�<'d�<ly�<N��<��<��<׶�<��<��<g��<X��<���<���<���<��<���<���<~�<f�<�J�<�+�<	�<���<��<V��<�Y�<�$�<^��<9��<m�<(�<���<���<Q@�<��<���<!4�<���<�l�<V�<���<$�<y��<5�<���<�6�<���<)�<뜱< �<�y�<M�<KI�<"��<��<mh�<���<��<�l�<��<��<�X�<뢚<w�<�/�<\s�<Ǵ�<n��<B2�<�n�<I��<��<��<�Q�<[��<'��<.��<K#�<�|<�y<su<��q<�7n<ՙj<��f<^c<��_<�#\<*�X<c�T<6TQ<-�M<?&J<�F< C<�p?<��;<�Y8<b�4<�N1<D�-<�Q*<��&<jd#<2�<[�<�!<c�<�b<	<�<m<�&<��<}Y�;���;���;+N�;��;��;���;c��;Ы�;2��;{Կ;K �;�;�;-��;�;�P�;�͝;[�;T��;���;Vg�;�6�;�.|;*r;h;�5^;.yT;��J;Y_A;(8;�.;E�%; ;�;��
;�H;�s�:��:���:aZ�:��:���:E�:�Q�:=�c:��D:`&:|K:b�9��9t�?9V#�8�=�y��5���������@��-�/��J�ǘe�����=��5U���U���B������ͺ˔ںB9线��( ��c���������v�m/%�H+�
]1��l7�0z=�4�C���I�z�O���U��[��a���g���m�\|s��uy��n��z���ǭ������-�����������n���۩���  �  7k=�
=�=�H=��=(�=k$=W� =�_ =���<b4�<ym�<ɥ�<@��<��<tI�<~�<���<J��<��<�E�<�t�<���<���<���<e#�<eK�<�q�<��<���<���<;��<��<M3�<�L�<)d�<`y�<T��<��<)��<۶�<��<���<a��<b��<���<���<��<��<���<���<~�<f�<�J�<�+�<	�<���< ��<V��<�Y�<�$�<_��<8��<m�<�'�<���<���<Z@�<��<���<#4�<���<�l�<P�<���<$�<z��<5�<���<�6�<���<)�<朱<'�<�y�<Q�<SI�<��<��<ch�<���<��<�l�<��<��<�X�<ޢ�<��<�/�<Ws�<Ǵ�<h��<P2�<�n�<N��<��<��<�Q�<b��<3��<$��<R#�<׫|<�y<su<��q<�7n<ęj<��f<�]c<��_<�#\<5�X<�T<$TQ<>�M<-&J<�F< C<�p?<��;<�Y8<q�4<�N1<]�-<�Q*<��&<gd#<#�<p�<m!<d�<�b<<�<�l<�&<��<�Y�;���;�;JN�;��;<��;��;���;ҫ�;>��;|Կ;A �;<�;���;2�;�P�;�͝;%[�;G��;̧�;=g�;�6�;�.|;>r;�h;
6^;0yT;��J;�_A;�8;$�.;�%;ʠ;"�;I�
;�H;s�:���:���:LZ�: �:��:m�:�Q�:a�c:��D:�`&:�K:��9�!�9'�?9�(�8�Q������������������/���J�ۗe�#���=���T���U��{B������ͺH�ں�8�C��( ��c�M��U�������k/%�BH+��\1�m7�z=��C��I�y�O�w�U���[�;�a�j�g��m��{s�Muy��n�ҳ����������������
���~���6��������  �  >k=�
=�=�H=��=/�=f$=Z� =�_ =���<a4�<|m�<Υ�<9��<��<kI�<%~�<���<G��<��<�E�<�t�<���< ��<���<^#�<[K�<�q�<���<���<���</��<��<K3�<�L�<5d�<Wy�<\��<��<*��<ֶ�<��<���<V��<_��<���<���<���<��<���<���<~�<f�<�J�<�+�<	�<���<���<f��<�Y�<�$�<Z��<7��<m�<�'�<���<���<V@�<���<���< 4�<���< m�<K�<���<$�<���<5�<���<�6�<���<")�<���<,�<�y�<F�<MI�<&��<��<\h�<¤<��<�l�<��<��<Y�<֢�<��<�/�<Ys�<ϴ�<g��<U2�<�n�<U��<��<��<�Q�<T��</��<��<b#�<ī|<�y<su<��q<�7n<��j<��f<�]c<��_<�#\<'�X<~�T<TQ<[�M<!&J<�F<
 C<�p?<��;<Y8<��4<�N1<k�-<�Q*<�&<qd#<�<w�<Z!<y�<�b<<$�<�l<�&<��<�Y�;'��;���;"N�;��;W��;Z��;���;���;O��;pԿ;1 �;5<�;ه�;P�;�P�;�͝;[�;4��;���;g�;�6�;~.|;�r;�h;6^;FyT;l�J;�_A;�8;��.;�%;��;�;�
;kI;�r�:���:t��:IZ�:�:0��:��:gQ�:щc:��D:�a&:mK:��9�"�9��?9Q1�8�b�������槻�?������/���J�U�e����N>��U��mU��_A������ͺʕں�8����( �uc����>������2/%�FH+�r\1��m7��y=�Z�C�p�I��O��U�ʍ[�y�a��g�=�m�|s�cuy��n�������������>��������������7���.����  �  9k=�
=�=�H=��='�=f$=X� =�_ =���<_4�<wm�<˥�<?��<��<uI�<~�<���<E��<��<�E�<�t�<���<���<���<h#�<dK�<�q�<|��<���<���<:��<��<H3�<�L�<5d�<^y�<S��<���<��<ڶ�<��<���<\��<i��<���<���<��<	��<���<���<~�<f�<�J�<�+�<	�<���<���<V��<�Y�<�$�<b��<7��<m�<�'�<���<���<a@�<��<���< 4�<���<�l�<[�<���<$�<���<5�<���<�6�<���<)�<朱<%�<�y�<M�<VI�<"��<��<\h�<���<��<�l�<��<��<�X�<ߢ�<{�<�/�<Ys�<Ŵ�<g��<L2�<�n�<R��<��<��<�Q�<`��<7��<��<X#�<ҫ|<�y<su<��q<�7n<��j<��f<�]c<��_<$\<,�X<v�T<TQ<G�M<'&J<"�F<% C<�p?<��;<�Y8<x�4<�N1<]�-<�Q*<��&<jd#<!�<i�<m!<e�<�b<
<$�<�l<�&<��<pY�;��;ʙ�;DN�;��;0��;y��;���;ͫ�;X��;cԿ;D �;7<�;�;-�;�P�;�͝;![�;D��;٧�;)g�;7�;�.|;&r;�h;�5^;CyT;��J;�_A;�8;�.;��%;��;��;B�
;�H;@s�:T��:���:@Z�:��:���:>�:�Q�:.�c:��D:�`&:bK:��9��9r�?9�*�8`U����s������V��m���/���J�=�e����=���T���U���B���� �ͺt�ں�8纨��( ��c�I����������}/%�GH+��\1�/m7��y=�|�C��I���O���U���[�\�a�6�g��m�(|s�tuy�Vn�泂���������%���)���ԧ������H�������  �  6k=�
=ک=�H=��=,�=m$=U� =�_ =|��<c4�<m�<ʥ�<D��<��<~I�<~�<Ʊ�<D��<��<�E�<�t�<���<���<���<_#�<UK�<�q�<y��<���<���<@��<��<I3�<�L�<'d�<iy�<D��<���<��<��<��<���<[��<R��<���<���<���<��<���<���<~�<f�<�J�<�+�<	�<���<��<S��<�Y�<�$�<`��<<��<m�<(�<���<���<L@�<��<���< 4�<���<�l�<]�<���<$�<y��<5�<���<�6�<���<)�<�<!�<�y�<B�<II�<(��<��<jh�<���<��<�l�<��<��<�X�<袚<t�<�/�<Ys�<̴�<p��<D2�<�n�<L��<��<��<�Q�<b��< ��<&��<T#�<׫|<�y<su<��q<�7n<ڙj<��f<^c<��_<�#\<1�X<��T<'TQ<=�M<2&J<��F< C<�p?<��;<�Y8<h�4<�N1<J�-<�Q*<	�&<gd#<,�<X�<�!<\�<�b<<�<�l<�&<��<�Y�;��;���;	N�;��;$��;���;���;��;#��;gԿ;] �;�;�; ��;��;�P�;�͝;N[�;B��;ӧ�;&g�;�6�;�.|;kr;&h;
6^;LyT;��J;a_A;^8;�.;%�%;��;�;��
;�H;At�:��:���:�Z�:��:���:��:#R�:��c:F�D:�`&:UK:��9��9��?9Y�8�A����Z�������1�����O�/�q�J���e�����>��aU��GU��&B��7��A�ͺ�ںH9����,( �
d� ����������I/%�H+��\1� m7�z=��C���I�L�O�w�U�@�[�*�a�Y�g��m��{s�vuy��n����p��������?�����������2��������  �  :k=�
=�=�H=��=)�=d$=W� =�_ =���<^4�<zm�<ĥ�<=��<��<qI�<~�<���<B��<��<�E�<�t�<���<���<���<j#�<aK�<�q�<{��<���<���<8��<��<N3�<�L�<%d�<ky�<Z��<���<��<۶�<���<���<d��<e��<���<���<��<��<��<���<~�<f�<�J�<�+�<	�<���<���<Y��<�Y�<�$�<]��<>��<m�<�'�<���<���<`@�<��<���<4�<���<�l�<_�<���<$�<v��<5�<���<�6�<���<)�<圱<"�<�y�<M�<XI�<"��<��<Yh�<���<��<�l�<��<��<�X�<ܢ�<{�<�/�<Ps�<ʴ�<g��<Q2�<�n�<O��<��<��<�Q�<]��<1��</��<\#�<��|<�y<su<��q<�7n<יj<��f<^c<��_<$\<#�X<w�T<TQ<K�M<G&J<�F<  C<�p?<��;<zY8<s�4<�N1<b�-<�Q*<��&<[d#<�<e�<f!<]�<�b<<�<�l<�&<��<�Y�;��;ә�;8N�;��;-��;i��;���;ī�;g��;}Կ;S �;�;�;)��;H�;�P�;�͝;&[�;��;��;Gg�;7�;�.|;Wr;�h;�5^;cyT;��J;�_A;�8;;�.;̢%;Ƞ;�;+�
;I;>s�:%��:���:�Z�:��:���:��:�Q�:�c:\�D:�b&:"J:�9��9ڝ?9�.�8�@����_���������2��
�/���J���e�
���=��iT���U��<B��Z��6�ͺ�ں9����( ��c�c����������V/%�HH+��\1�m7��y=�v�C�׉I�b�O���U���[���a��g�Z�m�|s��uy�_n�ó��v���ĭ���������ϧ������F���*����  �  ej=�	=��=}G=�=p�=t"=@� =�] =���<�.�<�g�<���<���<��<�A�<Pv�<l��<w��<u�<.<�<�j�<��<���<(��<8�<�>�<pd�<���<��<���<���<��<�"�<s;�<<R�<�f�< y�<��<���<ˡ�<U��<C��<C��<γ�<=��<��<}��<���<Y��<iw�<Hb�<�I�<�-�<H�<E��<���<F��<Nl�<^:�<��<<��<܍�<�L�<3�<��<�p�<U�<���<�p�<2�<���<IL�<��<pu�<�<ߎ�<��<՘�<.�<���<��<��<	�<^^�<TȬ<)/�<���<�<[P�<ժ�<U�<&W�<D��<���<F�<���<Q٘<��<�c�<]��<��<�%�<�b�<���<�؊<��<�I�<b��<2��<��<V�<��|<�y<�pu<��q<9n<�j<� g<�dc<��_<�.\<�X<9�T<�dQ<��M<_:J<L�F<;C<��?<��;<3w8<)�4<p1<��-<�v*<
 '<?�#<� <״<hO<N�< �<><��<2�<�^<�<���;Ok�;%�;���;ɐ�;Ad�;GE�;�5�;~4�;�B�;�`�;��;9˴;�;Pu�;_�;:`�;1�;���;h;�;���;�Ƀ;�R};4s;�4i;�U_;�U;Z�K;�wB;�9;��/;�&;"�;l�;"�;
G;Hd�:�s�:���:�.�:*ٲ:´�:���:��:]�f:t�G:w):`K:���9%ȟ9ĆJ90j�8d෎���W~�L ���V�Y���-�|�H��c��B~��X���v��J���ou��*X���%ͺ��ٺ9���)����8�)R�?��������H�$�}+��*1��>7��M=��ZC��cI�xjO��nU�qp[��qa��ng�Amm��is�fy�6b�殂���� ������}�����������_���ȯ���  �  Tj=�	=��=}G=�=j�=u"=>� =�] =���</�<�g�<���<���<��<B�<<v�<j��<���<}�<8<�<�j�<��<���<0��<6�<�>�<vd�<���<��<���<���<��<�"�<t;�<7R�<�f�<!y�<��<���<ġ�<8��<-��<_��<̳�<F��<��<w��<���<\��<yw�<Pb�<�I�<�-�<E�<@��<���<G��<:l�<i:�<��<L��<��<�L�<0�<��<�p�<R�<���<�p�<�<���<DL�<��<ru�< �<܎�<��<ᘷ<2�<ȓ�<��<��<��<]^�<hȬ<&/�<���<
�<^P�<ժ�<_�<2W�<T��<���<�E�<���<A٘<��<�c�<O��<��<�%�<�b�<���<�؊<��<�I�<e��<3��<�<6�<[�|<|y<�pu<�q<#9n<�j<� g<ec<��_<�.\<�X<(�T<�dQ<��M<�:J<X�F<=C<��?<��;<7w8<!�4<(p1<��-<�v*<��&<"�#<� <��<uO<&�<��<5><��<F�<�^<�<Q��;ok�;�;��;��;�c�;)E�;�5�;�4�;C�;�`�;��;(˴;F�;Vu�;��;3`�;�;��;;�;F��;�Ƀ;@S};�3s;�4i;�U_;�U;��K;4xB;9;��/; �&;��;(�;#�;hF;�d�:$t�:���:0/�:Kٲ:���:/��:���:��f:��G:u):rG:���9�Ɵ9�J9Bl�8R.���W~�/����U�����-�>�H��c��B~�~W���v��ց��>v���W���%ͺS�ٺy��)�ܵ�����Q�ă���������$��+�b*1�!>7��M=��ZC��cI�ojO��nU�ip[��pa��og��mm��is�fy��a�ۮ��鬅�B������n��������������������  �  Uj=�	=��=zG=�=j�=|"=6� =�] =|��</�<�g�<���<���<��<B�<:v�<o��<���<m�<1<�<�j�<���<���<?��<(�<�>�<}d�<���<1��<���<���<��<�"�<o;�<0R�<�f�<y�<$��<���<ѡ�<P��<.��<h��<���<N��<��<|��<���<H��<qw�<=b�<�I�<�-�<V�<C��<���<Y��<7l�<s:�<��<A��<Ѝ�<�L�<8�<��<�p�<>�<���<�p�<&�<ı�<<L�<��<du�<�<Վ�<��<ژ�<%�<̓�<��<.��<��<a^�<cȬ</�<���<�<kP�<Ǫ�<S�<"W�<H��<���<�E�<Ր�<:٘<��<�c�<M��<��<�%�<�b�<���<�؊<��<�I�<b��< ��<�<5�<��|<�y<�pu<�q<9n<�j<� g<ec<��_<�.\<��X<*�T<�dQ<��M<�:J<:�F<.C<��?<�;<Rw8<�4<!p1<��-<�v*<��&<(�#<� <��<�O<"�<�<,><��<7�<�^<	 <@��;�k�;��;���;���;�c�;�E�;x5�;�4�;�B�;�`�;��;˴;M�;!u�;��;`�;H�;x��;;�;i��;�Ƀ;S};�3s;�4i;�U_;�U;��K;�wB;`9;��/;��&;�; �;��;UF;�e�:�r�:��:�-�:�ز:��:��:j��:p�f:X�G:4u):�I:f��9�ğ98�J9�^�8{1෍���Y~������X�o��!�-���H�j�c�;B~��W���w��Ӏ��mv��(W��b&ͺ�ٺn�溺)�~�����JQ����'�������$��+��*1�A>7�uN=�YZC��cI�]jO��nU�q[��pa��og��lm��is�Pfy��a����嬅�f������������������|��������  �  Yj=�	=��=}G=�=g�={"=:� =�] =���<�.�<�g�<���<���<��<B�<8v�<s��<��<{�<><�<�j�<��<���<9��<1�<�>�<ud�<���<��<���<���<��<�"�<r;�<9R�<�f�<y�<��<���<���<K��<0��<Y��<ų�<P��<��<{��<���<V��<~w�<Bb�<�I�<�-�<F�<C��<���<G��<:l�<q:�<��<N��<ߍ�<�L�<6�<��<�p�<M�<���<�p�<#�<���<=L�<��<ou�<�<ݎ�<��<ݘ�</�<͓�<��<��<��<\^�<aȬ<"/�<���<�<hP�<˪�<c�<1W�<H��<���<�E�<���<C٘<��<�c�<Q��<��<�%�<�b�<���<�؊<��<�I�<i��<-��<�<=�<}�|<dy<�pu<�q<!9n<�j<� g<ec<��_<�.\<�X<�T<�dQ<��M<~:J<M�F<<C<��?<u�;<Mw8<�4<8p1<��-<�v*<  '<�#<� <��<zO<�<�<#><��<Q�<�^< <2��;�k�;�;���;ސ�;�c�;EE�;f5�;�4�;C�;�`�;��;-˴;G�;Pu�;��;`�;��;b��;;�;/��;�Ƀ;�S};�3s;�4i;�U_;�U;�K;�wB;A9;��/;�&;�;H�;)�;mF;ue�:Ws�:���:�.�:ٲ:���:���:O��:[�f:�G:Ku):�I:���9Kş9~�J9Ji�8�:෕���W~�U����V�E����-���H�$�c��B~��W��<w��,����v��_W�� &ͺ�ٺ��溺)�G������Q����n�������$��+��*1��=7� N=�rZC��cI��jO��nU��p[�qa��og�Smm�Fjs�-fy��a�߮��⬅�H���
���s���������������ȯ���  �  \j=�	=��={G=�=k�=x"=<� =�] =���<�.�<�g�<���<���<��<B�<Cv�<p��<��<s�<1<�<�j�<��<���<2��</�<�>�<pd�<���<��<���<���<��<�"�<i;�<;R�<�f�<%y�<��<���<ǡ�<G��<3��<W��<ȳ�<F��<��<y��<���<V��<lw�<Fb�<�I�<�-�<E�<E��<���<E��<Gl�<l:�<��<>��<܍�<�L�<3�<��<�p�<P�<���<�p�<!�<���<RL�<��<ru�<�<ߎ�<��<٘�<.�<Ó�<��<��<��<Y^�<dȬ<!/�<���<�<bP�<Ѫ�<X�<$W�<K��<���<F�<���<L٘<��<�c�<V��<��<�%�<�b�<���<�؊<��<�I�<b��<0��<
�<B�<m�|<�y<�pu<��q<*9n<�j<� g<�dc<��_<�.\<�X<9�T<�dQ<��M<q:J<S�F<2C<��?<��;<Aw8<�4<p1<��-<�v*<  '<+�#<� <ȴ<pO<6�<�<"><��<8�<�^<�<W��;vk�;�;
��;Ȑ�;�c�;?E�;�5�;�4�;�B�;�`�;���;7˴;�;fu�;h�;e`�;!�;S��;,;�;'��;�Ƀ;>S};4s;�4i;�U_;�U;w�K;�wB;9;E�/;�&;#�;v�;�;�F;(e�:�s�:���:�.�:�ز:ʹ�:Y��:���:��f:��G:�u):WI:=��9Wʟ96�J9�l�8\����Z~�J����V����-���H��c�2C~��W��Bw������%v���W���%ͺ��ٺZ�溉)󺅵����R�l��{�������$��+��*1�i>7� N=��ZC��cI�gjO��nU��p[�:qa�|og��mm��is��ey�Pb�ͮ�����;���3���j�������|���`���௚��  �  Xj=�	=��={G=�=h�=z"=<� =�] =���</�<�g�<���<���<��<B�<@v�<i��<���<v�<:<�<�j�<��<���<:��<+�<�>�<sd�<���< ��<���<���<��<�"�<n;�<?R�<�f�<%y�<��<���<���<K��<-��<a��<���<J��<��<y��< ��<Y��<sw�<Jb�<�I�<�-�<M�<>��<���<N��<=l�<j:�<��<D��<��<�L�<5�<��<�p�<E�<���<�p�<$�<���<<L�<��<tu�<�<⎺<��<ט�</�<Ɠ�<��<��<��<W^�<bȬ</�<���<�<aP�<Ӫ�<`�<'W�<S��<���<�E�<Ȑ�<?٘<��<�c�<M��<��<�%�<�b�<���<�؊<��<�I�<a��<(��<�<<�<|�|<qy<�pu<�q<(9n<��j<� g<�dc<��_<�.\<۔X<�T<�dQ<��M<�:J<I�F<2C<��?<x�;<Iw8<�4<%p1<��-<�v*<��&<4�#<� <��<�O</�<��<6><��<J�<�^<�<E��;�k�;��;��;Ԑ�;�c�;bE�;v5�;�4�;C�;�`�;��;I˴;�;fu�;��;`�;�;e��;;�;M��;�Ƀ;aS};�3s;�4i;�U_;�U;��K;xB;9;��/;A�&;�;%�;^�;�F;e�:�s�:��: /�:Nٲ:ᴢ:��:,��:h�f:g�G:�t):�I:���9�ğ9Z�J9�n�8k`�����X~�����vV�,��;�-���H� �c�vC~��W���w��
���hv���W���%ͺF�ٺ(��)�������Q�̃�s�������$��+��*1�G>7�N=�iZC� dI�fjO��nU��p[��pa��og�Tmm�js�Pfy��a�Ю�����#���%���q��������������������  �  Rj=�	=��=�G=�=h�={"=6� =�] =���<	/�<�g�<���<���<��<	B�<:v�<y��<���<r�<<<�<�j�<��<���<A��<1�<�>�<xd�<���<!��<���<���<��<�"�<p;�<5R�<�f�<y�<'��<���<���<P��<(��<a��<���<X��<��<}��<���<T��<vw�<Cb�<�I�<�-�<H�<C��<���<H��<<l�<z:�<��<G��<ߍ�<�L�<8�<��<�p�<B�<���<�p�<'�<���<AL�<��<iu�<�<ڎ�<��<ؘ�<*�<Փ�<��<��<��<]^�<dȬ</�<���<�<hP�<ƪ�<b�<&W�<N��<���<�E�<���<C٘<��<�c�<U��<��<�%�<�b�<���<�؊<��<�I�<n��<&��<�<1�<��|<jy<�pu<!�q<9n<��j<� g<�dc<��_<�.\<��X<�T<�dQ<��M<�:J<>�F<HC<��?<y�;<Mw8< �4<,p1<��-<�v*< '<"�#<� <��<~O<$�<�<4><��<M�<�^< <>��;�k�;	�;��;��;�c�;eE�;k5�;�4�;C�;�`�;��; ˴;&�;:u�;��;+`�;�;v��;�:�;N��;�Ƀ;�S};�3s;�4i;�U_;ݖU;��K;�wB;�9;��/;�&;�;E�;3�;yF;f�:~s�:I��:�.�:�ز:��:���:���:�f:��G:�t):J:h��99Ɵ9�J9Bd�8NY����X~������W�:��e�-���H��c��B~��W���w�������v��UW��z&ͺ$�ٺ:��U)�ִ�����Q����i�������$��+��*1�>7�]N=�iZC��cI�[jO�_nU��p[��pa�pg�2mm�.js��ey��a�����󬅻\��� �������u���y������������  �  Zj=�	=��=~G=�=k�=y"=;� =�] =���<�.�<�g�<���<���<��<B�<Fv�<n��<~��<t�<7<�<�j�<��<���<3��<1�<�>�<yd�<���<��<���<���<��<�"�<m;�<1R�<�f�<y�<��<���<���<N��<3��<[��<���<O��<߫�<z��<���<X��<tw�<Bb�<�I�<�-�<H�<F��<���<H��<Fl�<m:�<��<C��<ލ�<�L�<5�<��<�p�<I�<���<�p�<&�<���<HL�<��<lu�<�<׎�<��<ܘ�<(�<Ǔ�<��<��<��<_^�<_Ȭ<!/�<���<�<iP�<ͪ�<]�<&W�<G��<���<F�<���<O٘<��<�c�<S��<��<�%�<�b�<���<�؊<��<�I�<h��<'��<�<@�<��|<ty<�pu<�q<9n<�j<� g<ec<��_<�.\<�X< �T<�dQ<��M<�:J<?�F<@C<��?<��;<Hw8<�4<%p1<��-<�v*<  '</�#<� <д<rO<;�<�<!><��<D�<�^< <D��;{k�;	�;���;��;�c�;OE�;�5�;�4�;�B�;�`�;��;˴;@�;Iu�;��;@`�;�;m��;-;�;6��;�Ƀ;�S};�3s;�4i;�U_;�U;��K;�wB;#9;5�/;�&;)�;u�;.�;�F;9e�:Gs�:��:�.�:�ز:㴢:���:?��:��f:I�G:�u):�I:���9ȟ9��J9f�8�Aෙ��D[~�|���?X���_�-�?�H��c�xB~�X��Hw��n����v��GW��&ͺm�ٺ4���)󺤵����R�Q��z�������$�+��*1�)>7�N=��ZC��cI��jO��nU��p[�
qa��og�<mm�js�fy�b�宂�ଅ�g������s��������������������  �  Yj=�	=��={G=�=m�=t"=?� =�] =���</�<�g�<���<���<��<B�<Gv�<a��<���<�<0<�<�j�<��<���<4��<1�<�>�<rd�<���<��<���<���<��<�"�<n;�<=R�<�f�<%y�<��<���<���<F��<1��<[��<Ƴ�<E��<��<|��<���<Y��<pw�<Vb�<�I�<�-�<I�<B��<���<I��<Cl�<c:�<��<D��<ݍ�<�L�<3�<��<�p�<N�<���<�p�<!�<���<BL�<��<uu�<�<⎺<��<՘�<2�<œ�<��<��<��<X^�<`Ȭ<#/�<���<�<]P�<Ӫ�<X�</W�<\��<���<F�<���<J٘<��<�c�<M��<��<�%�<�b�<���<�؊<��<�I�<a��<+��<�<@�<q�|<oy<�pu<�q<#9n<�j<� g<�dc<��_<�.\<۔X<�T<�dQ<��M<:J<I�F<5C<��?<��;<3w8<&�4<p1<��-<�v*<��&<5�#<� <Ŵ<uO<>�<�<E><��<6�<�^<�<g��;}k�;�; ��;Ґ�;�c�;@E�;�5�;�4�;C�;�`�;��;A˴;�;fu�;��;&`�;��;Q��;%;�;8��;�Ƀ;:S};�3s;�4i;�U_;�U;��K;`xB;�9;$�/;#�&;�;S�;6�;�F;�d�:�t�:��:�.�:4ٲ:ʹ�:l��:���:z�f:!�G:u):[I:F��9�Ɵ9&�J9�o�8mj����X~�- ���U�D����-�
�H�>�c�IC~��W��"w�������u��X���%ͺ��ٺ���~(�e���}� R�u����������$��+�$*1�p>7��M=��ZC��cI�|jO��nU��p[�qa��og��mm�js�Wfy��a�ۮ�����2���+���z���������������د���  �  Vj=�	=��=|G=�=k�=x"=<� =�] =���</�<�g�<���<���<��<B�<Bv�<r��<���<m�<8<�<�j�<��<���<;��<*�<�>�<wd�<���<+��<���<���<��<�"�<o;�<5R�<�f�<y�<��<���<ˡ�<P��<-��<_��<���<N��<��<z��<���<W��<nw�<@b�<�I�<�-�<N�<F��<���<P��<Al�<r:�<��<@��<ݍ�<�L�<4�<��<�p�<C�<���<�p�<'�<���<>L�<��<gu�<�<ێ�<��<Ԙ�<'�<ʓ�<��<%��<��<\^�<bȬ</�<���<�<`P�<Ϫ�<]�< W�<J��<���<F�<ɐ�<H٘<��<�c�<R��<��<�%�<�b�<���<�؊<��<�I�<f��<"��<�<8�<��|<|y<�pu<�q<9n<��j<� g<�dc<|�_<�.\<�X<$�T<�dQ<��M<�:J<9�F<6C<��?<��;<Aw8<�4<p1<��-<�v*<��&<3�#<� <��<�O<2�<�<)><��<E�<�^<�<[��;�k�;��;���;��;�c�;�E�;}5�;�4�;�B�;�`�;
��;!˴;�;0u�;��;`�;2�;v��;;�;G��;�Ƀ;~S};�3s;�4i;�U_;��U;��K;�wB;U9;%�/;H�&;(�;U�;o�;�F;�e�:Vs�:ض�:�.�:&ٲ:ٴ�:I��:L��:�f:n�G:�t):J:;��9iş9ΏJ9b�8\a෉��Y~�� ��VX��,�-���H�[�c��B~��W���w�� ���)v���W���%ͺp�ٺ��溛)�[������Q����Z�������$��+��*1�`>7��M=��ZC��cI�fjO��nU��p[��pa��og�mm��is�Hfy��a��������X���������������������������  �  Sj=�	=��=�G=�=g�=~"=8� =�] =���<�.�<�g�<���<���<��<B�<7v�<w��<~��<�<C<�<�j�<���<���<5��<0�<�>�<yd�<���<��<���<���<��<�"�<v;�<-R�<�f�<y�<��<���<���<@��<)��<c��<³�<S��<ܫ�<}��<��<W��<�w�<Cb�<�I�<�-�<M�<@��<���<Q��<7l�<v:�<��<W��<ߍ�<�L�<<�<޽�<�p�<J�<���<�p�<�<���<8L�<��<eu�<&�<Վ�<��<☷<$�<ϓ�<��<��<��<\^�<bȬ</�<���<��<pP�<̪�<d�<5W�<H��<���<�E�<ʐ�<?٘<��<�c�<P��<��<�%�<�b�<���<�؊<��<�I�<m��<&��<�<3�<t�|<`y<�pu<�q<9n<�j<� g<ec<��_<�.\<�X<�T<�dQ<��M<�:J<C�F<GC<��?<u�;<Zw8<�4<Ap1<��-<�v*< '<&�#<� <��<�O<�<�<"><��<\�<�^< <"��;�k�;�;��;��;�c�;VE�;W5�;�4�;�B�;�`�;$��;�ʴ;s�;(u�;��;`�;��;8��;;�;V��;�Ƀ;�S};�3s;�4i;�U_;��U;N�K;�wB;Y9;��/;A�&;��;�;|�;TF;�e�:Es�:O��:�.�:2ٲ:T��:Y��:���:��f:��G:�t):H:���9ğ98�J9�_�8U෫���W~�����Y����-�b�H���c��B~��W��pw��4���0w���V��&ͺ�ٺ?�溿)�������Q�у�l�������$��+��*1��=7�'N=�<ZC�dI��jO�dnU��p[��pa��og�wmm�Sjs�fy��a�������������㩋�����������������ů���  �  Zj=�	=��={G=�=n�=y"=7� =�] =���< /�<�g�<���<���<��<B�<Bv�<s��<���<z�<&<�<�j�<��<���<6��<0�<�>�<qd�<���<"��<���<���<��<�"�<l;�<2R�<�f�<y�<��<���<̡�<N��<5��<W��<ų�<B��<��<���<���<G��<mw�<Kb�<�I�<�-�<R�<F��<���<S��<Dl�<o:�<��<B��<͍�<�L�<9�<��<�p�<L�<���<�p�<*�<���<JL�<��<hu�<�<׎�<��<Ԙ�<'�<Ó�<��<��<��<[^�<^Ȭ< /�<���<�<fP�<˪�<J�<+W�<P��<���<F�<Ȑ�<G٘<��<�c�<X��<��<�%�<�b�<���<�؊<��<�I�<_��<*��<�<A�<��|<�y<�pu<�q<9n<�j<� g<�dc<��_<�.\<�X<,�T<�dQ<��M<t:J<H�F<4C<��?<��;<Fw8<�4<p1<��-<�v*< '<4�#<� <��<�O<4�<�<3><��<#�<�^<�<v��;�k�;�;���;А�;d�;hE�;�5�;�4�;�B�;�`�;���;˴;!�;8u�;��;G`�;5�;q��;2;�;$��;�Ƀ; S};4s;�4i;�U_;x�U;|�K;xB;-9;>�/;l�&;.�;W�;��;�F;`e�:�s�:���:�-�:ٲ:$��:��:���:7�f:��G:�u):cJ:��9�ȟ9b�J9�b�8�_�`��vZ~�� ��_X�m��}�-���H���c�C~�X��Tw��}����u��xW��%&ͺ��ٺލ�8)�[������Q����N�����p�$��+�n*1��>7�cN=��ZC��cI�AjO��nU��p[�/qa��og�Gmm��is�fy�b��������e���.���������������z��������  �  \j=�	=��=xG=�=j�=q"=H� =�] =���<�.�<�g�<���<���<��<B�<@v�<e��<���<~�<;<�<�j�<ԗ�<���<1��<0�<�>�<nd�<���<��<���<���<��<�"�<m;�<@R�<�f�<.y�<��<���<���<E��<4��<U��<г�<:��<��<j��<��<h��<tw�<Sb�<�I�<�-�<E�<F��<���<E��<Bl�<_:�<��<I��<��<�L�< �<���<�p�<S�<���<�p�< �<���<AL�<��<|u�<�<⎺<��<ט�<:�<���<��<��<��<W^�<eȬ<"/�<���<�<JP�<䪤<e�<1W�<Q��<���< F�<���<L٘<��<�c�<O��<��<�%�<�b�<���<�؊<��<�I�<W��<7��<�<C�<j�|<ry<tpu<�q<;9n<�j<� g<�dc<��_<�.\<ŔX<�T<�dQ<��M<q:J<`�F<&C<��?<�;<(w8<K�4<p1<��-<�v*<��&<*�#<� <Ѵ<qO<1�<�<3><��<M�<�^<�<w��;rk�;�;��;Ð�;d�;(E�;|5�;S4�;/C�;�`�;���;M˴;�;�u�;v�;`�;��;J��;1;�;��; ʃ;�R};84s;14i; V_;~�U;��K;LxB;�9;(�/;�&;+�;j�;�;�F;jd�:+t�:p��:�/�:�ٲ:���:���:��:)�f:��G:�u):4I:��9"Ɵ9��J9Hw�82g�L��Y~������S����-���H�ӥc�iC~��W��.w������u��:Y���$ͺ��ٺ���-)�a�����R�f��U�������$�#+�*1�c>7�RM=��ZC�dI�6jO�oU�Hp[�Bqa�tog��mm�js��fy��a�����������?���P�������ت������쯚��  �  Zj=�	=��={G=�=n�=y"=7� =�] =���< /�<�g�<���<���<��<B�<Bv�<s��<���<z�<&<�<�j�<��<���<6��<0�<�>�<qd�<���<"��<���<���<��<�"�<l;�<2R�<�f�<y�<��<���<̡�<N��<5��<W��<ų�<B��<��<���<���<G��<mw�<Kb�<�I�<�-�<R�<F��<���<S��<Dl�<o:�<��<B��<͍�<�L�<9�<��<�p�<L�<���<�p�<*�<���<JL�<��<hu�<�<׎�<��<Ԙ�<'�<Ó�<��<��<��<[^�<^Ȭ< /�<���<�<fP�<˪�<J�<+W�<P��<���<F�<Ȑ�<G٘<��<�c�<X��<��<�%�<�b�<���<�؊<��<�I�<_��<*��<�<A�<��|<�y<�pu<�q<9n<�j<� g<�dc<��_<�.\<�X<,�T<�dQ<��M<t:J<H�F<4C<��?<��;<Fw8<�4<p1<��-<�v*< '<4�#<� <��<�O<4�<�<3><��<#�<�^<�<v��;�k�;�;���;А�;d�;hE�;�5�;�4�;�B�;�`�;���;˴;!�;8u�;��;G`�;5�;q��;2;�;$��;�Ƀ; S};4s;�4i;�U_;x�U;|�K;xB;-9;>�/;l�&;.�;W�;��;�F;`e�:�s�:���:�-�:ٲ:$��:��:���:7�f:��G:�u):cJ:��9�ȟ9b�J9�b�8�_�`��vZ~�� ��_X�m��}�-���H���c�C~�X��Tw��}����u��xW��%&ͺ��ٺލ�8)�[������Q����N�����p�$��+�n*1��>7�cN=��ZC��cI�AjO��nU��p[�/qa��og�Gmm��is�fy�b��������e���.���������������z��������  �  Sj=�	=��=�G=�=g�=~"=8� =�] =���<�.�<�g�<���<���<��<B�<7v�<w��<~��<�<C<�<�j�<���<���<5��<0�<�>�<yd�<���<��<���<���<��<�"�<v;�<-R�<�f�<y�<��<���<���<@��<)��<c��<³�<S��<ܫ�<}��<��<W��<�w�<Cb�<�I�<�-�<M�<@��<���<Q��<7l�<v:�<��<W��<ߍ�<�L�<<�<޽�<�p�<J�<���<�p�<�<���<8L�<��<eu�<&�<Վ�<��<☷<$�<ϓ�<��<��<��<\^�<bȬ</�<���<��<pP�<̪�<d�<5W�<H��<���<�E�<ʐ�<?٘<��<�c�<P��<��<�%�<�b�<���<�؊<��<�I�<m��<&��<�<3�<t�|<`y<�pu<�q<9n<�j<� g<ec<��_<�.\<�X<�T<�dQ<��M<�:J<C�F<GC<��?<u�;<Zw8<�4<Ap1<��-<�v*< '<&�#<� <��<�O<�<�<"><��<\�<�^< <"��;�k�;�;��;��;�c�;VE�;W5�;�4�;�B�;�`�;$��;�ʴ;s�;(u�;��;`�;��;8��;;�;V��;�Ƀ;�S};�3s;�4i;�U_;��U;N�K;�wB;Y9;��/;A�&;��;�;|�;TF;�e�:Es�:O��:�.�:2ٲ:T��:Y��:���:��f:��G:�t):H:���9ğ98�J9�_�8U෫���W~�����Y����-�b�H���c��B~��W��pw��4���0w���V��&ͺ�ٺ?�溿)�������Q�у�l�������$��+��*1��=7�'N=�<ZC�dI��jO�dnU��p[��pa��og�wmm�Sjs�fy��a�������������㩋�����������������ů���  �  Vj=�	=��=|G=�=k�=x"=<� =�] =���</�<�g�<���<���<��<B�<Bv�<r��<���<m�<8<�<�j�<��<���<;��<*�<�>�<wd�<���<+��<���<���<��<�"�<o;�<5R�<�f�<y�<��<���<ˡ�<P��<-��<_��<���<N��<��<z��<���<W��<nw�<@b�<�I�<�-�<N�<F��<���<P��<Al�<r:�<��<@��<ݍ�<�L�<4�<��<�p�<C�<���<�p�<'�<���<>L�<��<gu�<�<ێ�<��<Ԙ�<'�<ʓ�<��<%��<��<\^�<bȬ</�<���<�<`P�<Ϫ�<]�< W�<J��<���<F�<ɐ�<H٘<��<�c�<R��<��<�%�<�b�<���<�؊<��<�I�<f��<"��<�<8�<��|<|y<�pu<�q<9n<��j<� g<�dc<|�_<�.\<�X<$�T<�dQ<��M<�:J<9�F<6C<��?<��;<Aw8<�4<p1<��-<�v*<��&<3�#<� <��<�O<2�<�<)><��<E�<�^<�<[��;�k�;��;���;��;�c�;�E�;}5�;�4�;�B�;�`�;
��;!˴;�;0u�;��;`�;2�;v��;;�;G��;�Ƀ;~S};�3s;�4i;�U_;��U;��K;�wB;U9;%�/;H�&;(�;U�;o�;�F;�e�:Vs�:ض�:�.�:&ٲ:ٴ�:I��:L��:�f:n�G:�t):J:;��9iş9ΏJ9b�8\a෉��Y~�� ��VX��,�-���H�[�c��B~��W���w�� ���)v���W���%ͺp�ٺ��溛)�[������Q����Z�������$��+��*1�`>7��M=��ZC��cI�fjO��nU��p[��pa��og�mm��is�Hfy��a��������X���������������������������  �  Yj=�	=��={G=�=m�=t"=?� =�] =���</�<�g�<���<���<��<B�<Gv�<a��<���<�<0<�<�j�<��<���<4��<1�<�>�<rd�<���<��<���<���<��<�"�<n;�<=R�<�f�<%y�<��<���<���<F��<1��<[��<Ƴ�<E��<��<|��<���<Y��<pw�<Vb�<�I�<�-�<I�<B��<���<I��<Cl�<c:�<��<D��<ݍ�<�L�<3�<��<�p�<N�<���<�p�<!�<���<BL�<��<uu�<�<⎺<��<՘�<2�<œ�<��<��<��<X^�<`Ȭ<#/�<���<�<]P�<Ӫ�<X�</W�<\��<���<F�<���<J٘<��<�c�<M��<��<�%�<�b�<���<�؊<��<�I�<a��<+��<�<@�<q�|<oy<�pu<�q<#9n<�j<� g<�dc<��_<�.\<۔X<�T<�dQ<��M<:J<I�F<5C<��?<��;<3w8<&�4<p1<��-<�v*<��&<5�#<� <Ŵ<uO<>�<�<E><��<6�<�^<�<g��;}k�;�; ��;Ґ�;�c�;@E�;�5�;�4�;C�;�`�;��;A˴;�;fu�;��;&`�;��;Q��;%;�;8��;�Ƀ;:S};�3s;�4i;�U_;�U;��K;`xB;�9;$�/;#�&;�;S�;6�;�F;�d�:�t�:��:�.�:4ٲ:ʹ�:l��:���:z�f:!�G:u):[I:F��9�Ɵ9&�J9�o�8mj����X~�- ���U�D����-�
�H�>�c�IC~��W��"w�������u��X���%ͺ��ٺ���~(�e���}� R�u����������$��+�$*1�p>7��M=��ZC��cI�|jO��nU��p[�qa��og��mm�js�Wfy��a�ۮ�����2���+���z���������������د���  �  Zj=�	=��=~G=�=k�=y"=;� =�] =���<�.�<�g�<���<���<��<B�<Fv�<n��<~��<t�<7<�<�j�<��<���<3��<1�<�>�<yd�<���<��<���<���<��<�"�<m;�<1R�<�f�<y�<��<���<���<N��<3��<[��<���<O��<߫�<z��<���<X��<tw�<Bb�<�I�<�-�<H�<F��<���<H��<Fl�<m:�<��<C��<ލ�<�L�<5�<��<�p�<I�<���<�p�<&�<���<HL�<��<lu�<�<׎�<��<ܘ�<(�<Ǔ�<��<��<��<_^�<_Ȭ<!/�<���<�<iP�<ͪ�<]�<&W�<G��<���<F�<���<O٘<��<�c�<S��<��<�%�<�b�<���<�؊<��<�I�<h��<'��<�<@�<��|<ty<�pu<�q<9n<�j<� g<ec<��_<�.\<�X< �T<�dQ<��M<�:J<?�F<@C<��?<��;<Hw8<�4<%p1<��-<�v*<  '</�#<� <д<rO<;�<�<!><��<D�<�^< <D��;{k�;	�;���;��;�c�;OE�;�5�;�4�;�B�;�`�;��;˴;@�;Iu�;��;@`�;�;m��;-;�;6��;�Ƀ;�S};�3s;�4i;�U_;�U;��K;�wB;#9;5�/;�&;)�;u�;.�;�F;9e�:Gs�:��:�.�:�ز:㴢:���:?��:��f:I�G:�u):�I:���9ȟ9��J9f�8�Aෙ��D[~�|���?X���_�-�?�H��c�xB~�X��Hw��n����v��GW��&ͺm�ٺ4���)󺤵����R�Q��z�������$�+��*1�)>7�N=��ZC��cI��jO��nU��p[�
qa��og�<mm�js�fy�b�宂�ଅ�g������s��������������������  �  Rj=�	=��=�G=�=h�={"=6� =�] =���<	/�<�g�<���<���<��<	B�<:v�<y��<���<r�<<<�<�j�<��<���<A��<1�<�>�<xd�<���<!��<���<���<��<�"�<p;�<5R�<�f�<y�<'��<���<���<P��<(��<a��<���<X��<��<}��<���<T��<vw�<Cb�<�I�<�-�<H�<C��<���<H��<<l�<z:�<��<G��<ߍ�<�L�<8�<��<�p�<B�<���<�p�<'�<���<AL�<��<iu�<�<ڎ�<��<ؘ�<*�<Փ�<��<��<��<]^�<dȬ</�<���<�<hP�<ƪ�<b�<&W�<N��<���<�E�<���<C٘<��<�c�<U��<��<�%�<�b�<���<�؊<��<�I�<n��<&��<�<1�<��|<jy<�pu<!�q<9n<��j<� g<�dc<��_<�.\<��X<�T<�dQ<��M<�:J<>�F<HC<��?<y�;<Mw8< �4<,p1<��-<�v*< '<"�#<� <��<~O<$�<�<4><��<M�<�^< <>��;�k�;	�;��;��;�c�;eE�;k5�;�4�;C�;�`�;��; ˴;&�;:u�;��;+`�;�;v��;�:�;N��;�Ƀ;�S};�3s;�4i;�U_;ݖU;��K;�wB;�9;��/;�&;�;E�;3�;yF;f�:~s�:I��:�.�:�ز:��:���:���:�f:��G:�t):J:h��99Ɵ9�J9Bd�8NY����X~������W�:��e�-���H��c��B~��W���w�������v��UW��z&ͺ$�ٺ:��U)�ִ�����Q����i�������$��+��*1�>7�]N=�iZC��cI�[jO�_nU��p[��pa�pg�2mm�.js��ey��a�����󬅻\��� �������u���y������������  �  Xj=�	=��={G=�=h�=z"=<� =�] =���</�<�g�<���<���<��<B�<@v�<i��<���<v�<:<�<�j�<��<���<:��<+�<�>�<sd�<���< ��<���<���<��<�"�<n;�<?R�<�f�<%y�<��<���<���<K��<-��<a��<���<J��<��<y��< ��<Y��<sw�<Jb�<�I�<�-�<M�<>��<���<N��<=l�<j:�<��<D��<��<�L�<5�<��<�p�<E�<���<�p�<$�<���<<L�<��<tu�<�<⎺<��<ט�</�<Ɠ�<��<��<��<W^�<bȬ</�<���<�<aP�<Ӫ�<`�<'W�<S��<���<�E�<Ȑ�<?٘<��<�c�<M��<��<�%�<�b�<���<�؊<��<�I�<a��<(��<�<<�<|�|<qy<�pu<�q<(9n<��j<� g<�dc<��_<�.\<۔X<�T<�dQ<��M<�:J<I�F<2C<��?<x�;<Iw8<�4<%p1<��-<�v*<��&<4�#<� <��<�O</�<��<6><��<J�<�^<�<E��;�k�;��;��;Ԑ�;�c�;bE�;v5�;�4�;C�;�`�;��;I˴;�;fu�;��;`�;�;e��;;�;M��;�Ƀ;aS};�3s;�4i;�U_;�U;��K;xB;9;��/;A�&;�;%�;^�;�F;e�:�s�:��: /�:Nٲ:ᴢ:��:,��:h�f:g�G:�t):�I:���9�ğ9Z�J9�n�8k`�����X~�����vV�,��;�-���H� �c�vC~��W���w��
���hv���W���%ͺF�ٺ(��)�������Q�̃�s�������$��+��*1�G>7�N=�iZC� dI�fjO��nU��p[��pa��og�Tmm�js�Pfy��a�Ю�����#���%���q��������������������  �  \j=�	=��={G=�=k�=x"=<� =�] =���<�.�<�g�<���<���<��<B�<Cv�<p��<��<s�<1<�<�j�<��<���<2��</�<�>�<pd�<���<��<���<���<��<�"�<i;�<;R�<�f�<%y�<��<���<ǡ�<G��<3��<W��<ȳ�<F��<��<y��<���<V��<lw�<Fb�<�I�<�-�<E�<E��<���<E��<Gl�<l:�<��<>��<܍�<�L�<3�<��<�p�<P�<���<�p�<!�<���<RL�<��<ru�<�<ߎ�<��<٘�<.�<Ó�<��<��<��<Y^�<dȬ<!/�<���<�<bP�<Ѫ�<X�<$W�<K��<���<F�<���<L٘<��<�c�<V��<��<�%�<�b�<���<�؊<��<�I�<b��<0��<
�<B�<m�|<�y<�pu<��q<*9n<�j<� g<�dc<��_<�.\<�X<9�T<�dQ<��M<q:J<S�F<2C<��?<��;<Aw8<�4<p1<��-<�v*<  '<+�#<� <ȴ<pO<6�<�<"><��<8�<�^<�<W��;vk�;�;
��;Ȑ�;�c�;?E�;�5�;�4�;�B�;�`�;���;7˴;�;fu�;h�;e`�;!�;S��;,;�;'��;�Ƀ;>S};4s;�4i;�U_;�U;w�K;�wB;9;E�/;�&;#�;v�;�;�F;(e�:�s�:���:�.�:�ز:ʹ�:Y��:���:��f:��G:�u):WI:=��9Wʟ96�J9�l�8\����Z~�J����V����-���H��c�2C~��W��Bw������%v���W���%ͺ��ٺZ�溉)󺅵����R�l��{�������$��+��*1�i>7� N=��ZC��cI�gjO��nU��p[�:qa�|og��mm��is��ey�Pb�ͮ�����;���3���j�������|���`���௚��  �  Yj=�	=��=}G=�=g�={"=:� =�] =���<�.�<�g�<���<���<��<B�<8v�<s��<��<{�<><�<�j�<��<���<9��<1�<�>�<ud�<���<��<���<���<��<�"�<r;�<9R�<�f�<y�<��<���<���<K��<0��<Y��<ų�<P��<��<{��<���<V��<~w�<Bb�<�I�<�-�<F�<C��<���<G��<:l�<q:�<��<N��<ߍ�<�L�<6�<��<�p�<M�<���<�p�<#�<���<=L�<��<ou�<�<ݎ�<��<ݘ�</�<͓�<��<��<��<\^�<aȬ<"/�<���<�<hP�<˪�<c�<1W�<H��<���<�E�<���<C٘<��<�c�<Q��<��<�%�<�b�<���<�؊<��<�I�<i��<-��<�<=�<}�|<dy<�pu<�q<!9n<�j<� g<ec<��_<�.\<�X<�T<�dQ<��M<~:J<M�F<<C<��?<u�;<Mw8<�4<8p1<��-<�v*<  '<�#<� <��<zO<�<�<#><��<Q�<�^< <2��;�k�;�;���;ސ�;�c�;EE�;f5�;�4�;C�;�`�;��;-˴;G�;Pu�;��;`�;��;b��;;�;/��;�Ƀ;�S};�3s;�4i;�U_;�U;�K;�wB;A9;��/;�&;�;H�;)�;mF;ue�:Ws�:���:�.�:ٲ:���:���:O��:[�f:�G:Ku):�I:���9Kş9~�J9Ji�8�:෕���W~�U����V�E����-���H�$�c��B~��W��<w��,����v��_W�� &ͺ�ٺ��溺)�G������Q����n�������$��+��*1��=7� N=�rZC��cI��jO��nU��p[�qa��og�Smm�Fjs�-fy��a�߮��⬅�H���
���s���������������ȯ���  �  Uj=�	=��=zG=�=j�=|"=6� =�] =|��</�<�g�<���<���<��<B�<:v�<o��<���<m�<1<�<�j�<���<���<?��<(�<�>�<}d�<���<1��<���<���<��<�"�<o;�<0R�<�f�<y�<$��<���<ѡ�<P��<.��<h��<���<N��<��<|��<���<H��<qw�<=b�<�I�<�-�<V�<C��<���<Y��<7l�<s:�<��<A��<Ѝ�<�L�<8�<��<�p�<>�<���<�p�<&�<ı�<<L�<��<du�<�<Վ�<��<ژ�<%�<̓�<��<.��<��<a^�<cȬ</�<���<�<kP�<Ǫ�<S�<"W�<H��<���<�E�<Ր�<:٘<��<�c�<M��<��<�%�<�b�<���<�؊<��<�I�<b��< ��<�<5�<��|<�y<�pu<�q<9n<�j<� g<ec<��_<�.\<��X<*�T<�dQ<��M<�:J<:�F<.C<��?<�;<Rw8<�4<!p1<��-<�v*<��&<(�#<� <��<�O<"�<�<,><��<7�<�^<	 <@��;�k�;��;���;���;�c�;�E�;x5�;�4�;�B�;�`�;��;˴;M�;!u�;��;`�;H�;x��;;�;i��;�Ƀ;S};�3s;�4i;�U_;�U;��K;�wB;`9;��/;��&;�; �;��;UF;�e�:�r�:��:�-�:�ز:��:��:j��:p�f:X�G:4u):�I:f��9�ğ98�J9�^�8{1෍���Y~������X�o��!�-���H�j�c�;B~��W���w��Ӏ��mv��(W��b&ͺ�ٺn�溺)�~�����JQ����'�������$��+��*1�A>7�uN=�YZC��cI�]jO��nU�q[��pa��og��lm��is�Pfy��a����嬅�f������������������|��������  �  Tj=�	=��=}G=�=j�=u"=>� =�] =���</�<�g�<���<���<��<B�<<v�<j��<���<}�<8<�<�j�<��<���<0��<6�<�>�<vd�<���<��<���<���<��<�"�<t;�<7R�<�f�<!y�<��<���<ġ�<8��<-��<_��<̳�<F��<��<w��<���<\��<yw�<Pb�<�I�<�-�<E�<@��<���<G��<:l�<i:�<��<L��<��<�L�<0�<��<�p�<R�<���<�p�<�<���<DL�<��<ru�< �<܎�<��<ᘷ<2�<ȓ�<��<��<��<]^�<hȬ<&/�<���<
�<^P�<ժ�<_�<2W�<T��<���<�E�<���<A٘<��<�c�<O��<��<�%�<�b�<���<�؊<��<�I�<e��<3��<�<6�<[�|<|y<�pu<�q<#9n<�j<� g<ec<��_<�.\<�X<(�T<�dQ<��M<�:J<X�F<=C<��?<��;<7w8<!�4<(p1<��-<�v*<��&<"�#<� <��<uO<&�<��<5><��<F�<�^<�<Q��;ok�;�;��;��;�c�;)E�;�5�;�4�;C�;�`�;��;(˴;F�;Vu�;��;3`�;�;��;;�;F��;�Ƀ;@S};�3s;�4i;�U_;�U;��K;4xB;9;��/; �&;��;(�;#�;hF;�d�:$t�:���:0/�:Kٲ:���:/��:���:��f:��G:u):rG:���9�Ɵ9�J9Bl�8R.���W~�/����U�����-�>�H��c��B~�~W���v��ց��>v���W���%ͺS�ٺy��)�ܵ�����Q�ă���������$��+�b*1�!>7��M=��ZC��cI�ojO��nU�ip[��pa��og��mm��is�fy��a�ۮ��鬅�B������n��������������������  �  �i=�=��=9F=��=݂=� =T� =�[ =��<#*�<�b�<��<���<��<R;�<:o�<���<���<0�<x3�<�a�<H��<ӹ�<���<A�<03�<�X�<`|�<)��<j��<���<%��<��<�+�<#B�<%V�<h�<\w�<i��<ێ�<��<I��<���<���<���<���<���<���<q�<_�<vI�<i0�<�<��<���<���<�~�<�P�<S�<f��<���<�p�<s/�<���<���<%S�<��<f��<)S�<���<^��<(/�<�ž<�X�<��<�r�<���<W}�< ��<y�<��<ff�<�ׯ<�E�<`��<��<�{�<ݧ<�:�<��<S�<�C�<���< �<5�<���<�ɘ<�<0V�<e��<�ڑ<l�<^X�<���<
Њ<�	�<�B�<"z�<Ѱ�<�<��<̟|<}y<\nu<��q<m:n<ԟj<vg<Akc<��_<y8\<T�X<8	U<^sQ<{�M<�LJ<2�F<�-C<ɡ?<�<<��8<Y5<�1<J.<��*<�"'<��#<�D <g�<�x<�</�<�k<�<��<��<S<�8�;��;��;M<�;\�;��;���;��;���;Ǿ�;���;r�;�J�;���;��;�d�;��;�p�;��;;�;=}�;�L�;X~;8t;7j;fV`;��V;��L;rC;H:;��0;D�';͘;��;��;V);{!�:�'�:�a�:���:^r�:^D�:�H�:�x�:G�i:o�J:�8,:�:��9�פ9�]T9�8r������%�u�Բ��L�_����+��	G���a�Ĕ|�����q���4å�e���w���~̺�Bٺ���ȗ�P*������[G��v�ǟ���$�M�*�Z�0��7��&=�>6C��AI�#KO�5RU�LV[��Ya�Yg��Zm��Ys�AXy��V�&���©��8���B����������8���v�������  �  �i=�=��=:F=��=ׂ=� =X� =�[ =��<2*�<�b�<��<���<��<];�<-o�<���<���<8�<3�<�a�<W��<Ź�<���<9�<23�<�X�<9|�<0��<h��<���<#��<��<�+�<&B�<(V�<�g�<Yw�<^��<��<Ԗ�<)��<Ȟ�<���<���<���<���<���<�q�<$_�<{I�<t0�<��<��<���<���<�~�<yP�<]�<p��<���< q�<�/�<���<���<*S�<��<l��<S�<���<c��</�<�ž<�X�<��<�r�<���<W}�<��<!y�<��<jf�<�ׯ<�E�<b��<��<�{�<�ܧ<�:�<#��<[�<�C�<Ӗ�<&�<5�<���<�ɘ<�<(V�<Y��<�ڑ<j�<kX�<���<Њ<�	�<�B�<)z�<ΰ�<��<��<̟|<�y<Wnu<��q<J:n<ܟj<~g<Ekc<��_<�8\<Q�X<=	U<isQ<-�M<�LJ<1�F<�-C<ʡ?<k<<ߑ8<e5<�1<F.<�*<�"'<��#<�D <T�<�x<�<2�<�k<<��<��<1S<s8�;��;���;U<�;:�;i��;Ի�;���;ɮ�;���;���;}�;�J�;���;���;�d�;��;q�;��;N��;Y}�;�L�;YX~;�7t;7j;�V`;̕V;c�L;/rC;�:;=�0;"�';И;g�;��;�(;"�:4(�:c�:H��:*s�:�D�:+H�:=y�:��i:)�J:85,:S�:��9�Ԥ9�\T9l�8P������u��Ӳ��N�ݪ���+��	G��a�ǖ|��������å�M��������}̺MBٺ�废���)��o�����G��v����$���*�k�0�!7��&=��5C��AI�%KO��QU�eV[��Ya��Zg��Zm��Ys�WXy��V�n�������'���<���ϩ�����<���l���괚��  �  �i=�=��=;F=��=҂=� =O� =�[ =��<.*�<�b�<��<���<w�<k;�<,o�<���<���<*�<3�<�a�<]��<���<���<6�<13�<�X�<8|�<H��<]��<���<!��<��<�+�<B�<1V�<�g�<cw�<V��<��<��<*��<מ�<���<���<���<���<���<xq�<$_�<gI�<t0�<��<��<���<���<�~�<yP�<^�<]��<���<�p�<x/�<���<���<4S�<��<x��<S�<���<t��</�<�ž<�X�<��<�r�<���<Y}�<��<(y�<��<�f�<�ׯ<�E�<g��<��<�{�<�ܧ<�:�<��<Y�<�C�<Ė�<&�<5�<���<�ɘ<�<.V�<Z��<�ڑ<V�<mX�<锌<Њ<�	�<�B�<.z�<°�<��<��<��|<�y<Inu<��q<;:n<�j<og<Skc<~�_<�8\<G�X<4	U<�sQ<%�M<�LJ< �F<�-C<ݡ?<X<<�8<D5<
�1<".<�*<�"'<��#<�D <*�<�x<�<0�<�k<�<��<r�<<S<;8�;>��;��;T<�;u�;h��;4��;խ�;Ԯ�;���;���;��;�J�;ᘯ;���;�d�;��;:q�;��;S��;�}�;�L�;�X~;�7t;7j;�V`;W�V;d�L;�qC;�:;9�0;��';��;0�;��;�(;."�:'�:�b�:���:�r�:�D�:~G�:�y�:��i:��J:�5,:)�:�9~Ҥ9GaT9�g�8���c��X�u�tӲ��O���)�+��G�M�a�4�|�8���d���N¥�!���n���b~̺{Bٺ��应���)��o��G�%H�Sv�؟�	�$���*��0�7�'=��5C�4BI�
KO��QU��V[��Xa��Zg�%Zm��Ys��Xy�TV���������G������橎�󪑻P���~��������  �  �i=�=��=;F=��=ق=� =Q� =�[ =��<+*�<�b�<��<���<��<_;�<,o�<���<���<6�<�3�<�a�<_��<Ĺ�<���<=�</3�<�X�<;|�<0��<_��<���<��<��<�+�<B�<.V�<�g�<\w�<`��<ێ�<Ֆ�<.��<˞�<���<���<���<���<���<�q�<-_�<uI�<q0�<��<��<���<���<�~�<{P�<[�<i��<���<q�<}/�<��<���<-S�<��<k��<S�<���<_��</�<�ž<�X�<��<�r�<���<_}�<��<'y�<��<if�<�ׯ<�E�<a��<��<�{�<�ܧ<;�<��<g�<�C�<ǖ�<)�<5�<���<�ɘ<�<(V�<c��<�ڑ<e�<uX�<<Њ<�	�<�B�<*z�<ǰ�<��<��<Ο|<vy<]nu<��q<Q:n<�j<bg<Zkc<��_<8\<U�X<*	U<esQ<2�M<�LJ<$�F<�-C<ӡ?<r<<�8<I5<�1<B.<�*<�"'<��#<�D <K�<�x<�<;�<�k<<��<r�<AS<l8�;��;��;I<�;_�;t��;Ի�;ۭ�;ܮ�;���;���;��;�J�;Ԙ�;���;�d�;��;�p�;��;b��;g}�;�L�;pX~;�7t;a7j;�V`;V;��L;rC;�:;O�0;>�';��;]�;��;�(;�!�:�'�:_c�:���:s�:oE�:�G�:yy�:|�i:
�J:*6,:��:��9�Ԥ9_T9�p�8����J���u�Ҳ�MO�8����+��	G���a���|����������¥�s���&���P~̺�Aٺ8��Y���)��s�����G��v�����$��*���0��7��&=��5C��AI�!KO��QU��V[�JYa��Zg��Zm�Zs�?Xy��V�`�������`�������������4�������𴚻�  �  �i=�=��=;F=��=ق=� =T� =�[ =��<**�<�b�<��<���<��<Z;�<5o�<���<���<.�<|3�<�a�<U��<ɹ�<���<A�<53�<�X�<D|�<1��<s��<���<��<��<�+�< B�<&V�<�g�<Nw�<i��<��<ۖ�<5��<ƞ�<���<���<���<���<���<�q�<_�<xI�<m0�<�<��<���<���<�~�<�P�<V�<m��<���< q�<q/�<���<���<"S�<��<k��<S�<���<k��<)/�<�ž<�X�<��<�r�<���<]}�<��<y�<��<lf�<�ׯ<�E�<f��<��<�{�<�ܧ<�:�<��<Z�<�C�<Ζ�<$�<5�<���<�ɘ<�<,V�<c��<�ڑ<d�<cX�<���<Њ<�	�<�B�<(z�<԰�<��<��<П|<�y<anu<v�q<X:n<ԟj<ug<Akc<��_<u8\<R�X<S	U<hsQ<E�M<�LJ<<�F<�-C<š?<s<<ϑ8<W5<��1<9.<
�*<�"'<��#<�D <_�<�x<�<:�<�k<�<��<v�<,S<�8�;���;��;c<�;P�;���;ػ�;-��;���;���;���;q�;�J�;���;���;�d�;��;1q�;��;}��;R}�;�L�;)X~;�7t;7j;nV`;��V;	�L;rC;j:;��0;5�';ݘ;��;v�;);�!�:(�:.b�:N��:Br�:�D�:&H�:�x�:��i:��J:�6,:��:��97ؤ9�WT9�r�8
������o�u�}Ҳ�bO�ʫ�2�+�D	G���a���|�I��������å����Ĩ��o~̺fBٺ�����*��&����vG��v�����$�(�*���0�]7��&=�6C��AI�5KO�RU�5V[��Ya�\Zg��Zm�wYs�.Xy��V�R�������9���C�������$���:���A���봚��  �  �i=�=��=8F=��=ق=� =W� =�[ =��<-*�<�b�<��<���<~�<e;�<5o�<��<���<2�<�3�<�a�<U��<ƹ�<���<6�<+3�<�X�<@|�<4��<_��<���<'��<��<�+�<*B�<&V�<�g�<^w�<T��<��<ܖ�<0��<͞�<���<���<���<���<���<�q�<"_�<uI�<i0�<��<��<���<���<�~�<�P�<Q�<i��<���<q�<s/�<���<���<+S�<��<q��<S�<���<g��</�<�ž<�X�<��<�r�<���<[}�<��<y�<��<nf�<�ׯ<�E�<b��<��<�{�<�ܧ<�:�<��<`�<�C�<̖�<�<5�<���<�ɘ<�<2V�<X��<�ڑ<e�<oX�<���<Њ<�	�<�B�<%z�<ư�<��<��<ן|<~y<=nu<��q<T:n<ϟj<�g<<kc<��_<�8\<6�X<4	U<psQ<;�M<�LJ<!�F<�-C<ڡ?<q<<Б8<b5<�1<;.<�*<�"'<��#<�D <8�<�x<�<�<�k<�<��<��<,S<u8�;-��;��;<<�;e�;���;��;ݭ�;���;Ͼ�;���;o�;�J�;���;���;�d�;��;q�;��;h��;n}�;�L�;YX~;�7t;07j;�V`;ՕV;W�L;�qC;N:;d�0;��';��;E�;��;);b!�:�'�:�b�:p��:`r�:E�:H�:Yy�:x�i:��J:E6,:i�:��9�Ҥ9y]T9u�8���������u��Ҳ��M�m����+��G� �a�i�|�~���;����¥�e�������~̺Bٺ������*��&��m��G�v�����$��*���0��7��&=�6C��AI��JO�RU��V[�ZYa�|Zg��Zm��Ys��Xy�PV�Z���˩�����N�������񪑻s���~���ܴ���  �  �i=�=��=;F=��=ւ=� =Q� =�[ =��<2*�<�b�<��<���<��<`;�<(o�<���<���<4�<�3�<�a�<`��<���<���<7�</3�<�X�<8|�<<��<c��<���<��<��<�+�<!B�<*V�<�g�<^w�<\��<��<ז�<+��<Ԟ�<���<���<���<���<���<~q�<(_�<sI�<u0�<��<��<���<���<�~�<vP�<]�<g��<���<�p�<t/�<��<���<3S�<��<x��<S�<���<m��</�<�ž<�X�<��<�r�<���<Y}�<��<(y�<��<vf�<�ׯ<�E�<g��<��<�{�<�ܧ<;�<��<^�<�C�<̖�<'�<�4�<���<�ɘ<�<'V�<Z��<�ڑ<c�<rX�<<Њ<�	�<�B�<.z�<Ű�<��<��<ן|<�y<Xnu<��q<8:n<�j<wg<Qkc<~�_<x8\<U�X<?	U<vsQ<*�M<�LJ< �F<�-C<ˡ?<e<<�8<L5<�1<>.<�*<�"'<��#<�D <T�<�x<�<7�<�k<<��<r�<CS<S8�;0��;��;I<�;r�;f��;��;��;߮�;���;���;��;�J�;Ƙ�;���;�d�;��;,q�;��;T��;�}�;�L�;�X~;�7t;b7j;�V`;��V;��L;�qC;�:;-�0;E�';�;x�;��;�(;!"�:�'�:c�:��:xr�:�E�:yG�:�y�:��i:��J:�5,:��:a�9Ԥ9�^T9Ue�8������͵u��Ӳ�Q���P�+��G��a�R�|�4���b���{¥�쿲�
����~̺&BٺY�����)��������G�vv����$���*���0��7��&=��5C�BI�<KO��QU��V[�,Ya��Zg��Zm��Ys�SXy��V���������5���$���穎����4���i���Ѵ���  �  �i=�=��=>F=��=ւ=� =U� =�[ =
��<"*�<�b�<��<���<��<W;�<8o�<��<���<-�<�3�<�a�<Z��<���<���<@�<03�<�X�<B|�<9��<e��<���<��<��<�+�<B�<2V�<�g�<Pw�<^��<��<ۖ�<0��<ɞ�<���<���<���<���<���<�q�<!_�<pI�<k0�<�<��<���<���<�~�<�P�<Y�<c��<���<q�<v/�<���<���<,S�<��<n��<S�<���<h��</�<�ž<�X�<��<�r�<���<c}�<��<y�<��<qf�<�ׯ<�E�<c��<��<�{�<�ܧ<�:�<��<a�<�C�<�<)�<5�<���<�ɘ<
�<0V�<g��<�ڑ<_�<jX�<���<Њ<�	�<�B�</z�<Ͱ�<��<��<՟|<�y<Tnu<o�q<S:n<�j<[g<Rkc<��_<i8\<N�X<;	U<rsQ<?�M<�LJ<.�F<�-C<��?<e<<ߑ8<]5<	�1<4.<��*<�"'<��#<�D <h�<�x<�<C�<�k<�<��<��<8S<W8�;
��;��;N<�;M�;���;���;���;���;���;���;�;�J�;蘯;���;�d�;��;q�;��;j��;_}�;�L�;}X~;�7t;77j;�V`;ЕV;M�L;�qC;^:;��0;E�';ʘ;��;��;6);�!�:o'�:�b�:n��:�r�:9E�:�G�:fy�:��i:`�J:�5,:k�:�9�Ԥ9�XT9�r�8n�����u��в��O�p���+��G���a��|�u���Ͱ��å�����q���*~̺�Aٺ��庳��)��
����PG��v�ɟ���$�Q�*���0�#7��&=��5C�BI�SKO��QU�iV[��Ya�qZg��Zm��Ys�cXy��V�\�������m���"�������<���C���p���״���  �  �i=�=��=8F=��=܂=� =X� =�[ =��<.*�<�b�<��<���<��<Y;�<9o�<��<���<:�<�3�<�a�<S��<̹�<���<:�</3�<�X�<=|�<,��<e��<���<"��<��<�+�<%B�<#V�<�g�<Yw�<`��<ߎ�<֖�<+��<Ȟ�<���<���<���<���<���<�q�<_�<�I�<f0�<�<��<���<���<�~�<�P�<O�<x��<���<q�<z/�<���<���<!S�<��<k��<S�<���<`��</�<�ž<�X�<��<�r�<���<Z}�<��<y�<��<ff�<�ׯ<�E�<`��<��<�{�<�ܧ<�:�< ��<_�<�C�<ז�<�<5�<���<�ɘ<
�<2V�<]��<�ڑ<s�<hX�<���<Њ<�	�<�B�< z�<Ѱ�<��<��<Ɵ|<�y<Unu<��q<P:n<ןj<�g<Akc<��_<�8\<J�X<7	U<`sQ<4�M<�LJ<1�F<�-C<С?<�<<͑8<h5<�1<V.<�*<�"'<��#<�D <R�<�x<�<�<�k<<��<��<(S<�8�;��;���;J<�;B�;}��;ǻ�;���;���;���;���;x�;�J�;���;���;�d�;��;q�;��;U��;Y}�;�L�;X~;8t;97j;�V`;�V;?�L;~rC;5:;o�0;W�';͘;q�;��;);<!�:�(�:�b�:���:�r�:�D�:�H�:�x�:�i:�J:�5,:�::�9xդ9�[T9gr�8����?����u�dӲ�jN�5����+��	G�H�a�[�|��������Jå�ʾ��⨿��}̺Bٺ,��\���*�������G��v������$��*�#�0�77�w&=�
6C��AI�KO�CRU�NV[��Ya��Zg��Zm��Ys�^Xy�rV�a����������D���ũ������K���y��������  �  �i=�=��==F=��=ׂ=� =S� =�[ =��<2*�<�b�<��<���<��<e;�<5o�<���<���<)�<�3�<�a�<\��<���<���<;�<43�<�X�<9|�<?��<e��<���<!��<��<�+�<B�<)V�<�g�<^w�<Y��<��<��</��<Ҟ�<���<���<���<���<���<�q�<_�<sI�<t0�< �<��<���<���<�~�<�P�<^�<i��<���<�p�<v/�<���<���<-S�<��<u��<S�<���<q��</�<�ž<�X�<��<�r�<���<X}�<��<#y�<��<zf�<�ׯ<�E�<i��<��<�{�<�ܧ<�:�<��<[�<�C�<Ж�<%�<5�<���<�ɘ<�<0V�<_��<�ڑ<^�<gX�<�<Њ<�	�<�B�<,z�<̰�<��<��<�|<�y<Mnu<��q<>:n<ߟj<ng<Hkc<~�_<�8\<H�X<C	U<�sQ<&�M<�LJ<-�F<�-C<͡?<j<<ܑ8<T5<�1<+.<�*<�"'<��#<�D <>�<�x<�<2�<�k<�<��<x�<;S<_8�;"��; ��;_<�;|�;m��;��;��;ɮ�;���;���;r�;�J�;Ř�;���;�d�;��;6q�;��;f��;�}�;�L�;dX~;�7t;7j;�V`;��V;�L;�qC;�:;l�0;n�';��;]�;��;);("�:�'�:2b�:��:�r�:�D�:�G�:xy�:��i:A�J:�6,:��:t�9CԤ9�]T9�j�8ܒ�����?�u��Ӳ��O깭���+�dG�z�a���|��������¥�����s���M~̺XBٺ1��Җ��)��2�����G�Uv�ǟ���$���*���0�=7��&=��5C��AI�KO��QU�rV[�0Ya��Zg�bZm��Ys�Xy�sV���������H���6���婎�����N���a��������  �  �i=�=��=@F=��=ׂ=� =P� =�[ =	��<,*�<�b�<��<���<��<f;�<*o�<��<���<2�<�3�<�a�<f��<���<���<<�<(3�<�X�<1|�<7��<V��<���<��<��<�+�<B�<6V�<�g�<^w�<T��<��<Җ�<.��<̞�<���<���<���<���<���<�q�<1_�<lI�<v0�<��<��<���<���<�~�<xP�<a�<`��<���<q�<v/�<��<���<4S�<��<n��<S�<���<g��</�<�ž<�X�<��<�r�<���<a}�<��<%y�<��<rf�<�ׯ<�E�<]��<��<�{�<�ܧ<;�<��<m�<�C�<Ŗ�<,�<5�<���<�ɘ<�<(V�<c��<�ڑ<^�<�X�<<Њ<�	�<�B�<3z�<���<��<��<П|<ty<Qnu<��q<A:n<��j<Mg<ckc<��_<t8\<N�X<#	U<msQ<$�M<�LJ<�F<�-C<ɡ?<i<<�8<G5<4�1<2.<�*<�"'<��#<�D <K�<�x<�<D�<�k<�<��<j�<OS<E8�;0��;��;0<�;o�;M��;��;���;Ѯ�;���;���;��;�J�;���;���;�d�;��;q�;z�;a��;j}�;�L�;�X~;�7t;\7j;�V`;ЕV;��L;�qC;�:;T�0;N�';��;k�;��;�(;\"�:<'�:�c�:���:�r�:�E�:wG�:�y�:��i:Y�J:I6,:��:��9�Ѥ9_T9@i�8�b�����A�u��Ѳ��P�Z����+�|G���a��|�ȉ��/���v¥����ɧ���~̺7Aٺ?�庁��)�����m��G�iv�����$���*���0�z7��&=��5C��AI�LKO��QU��V[�>Ya��Zg��Zm�Zs�mXy��V�����w�����������ש��%���C�������ᴚ��  �  �i=�=��=:F=��=ڂ=� =R� =�[ =��<0*�<�b�<��<���<��<];�<2o�<���<���<0�<~3�<�a�<S��<ƹ�<���<<�</3�<�X�<A|�<5��<j��<���<��<��<�+�< B�<%V�<�g�<]w�<d��<��<ז�<9��<Ȟ�<���<���<���<���<���<~q�<_�<vI�<o0�<�<��<���<���<�~�<~P�<X�<j��<���<�p�<n/�<���<���<)S�<��<k��<S�<���<n��<!/�<�ž<�X�<��<�r�<���<U}�<��<%y�<��<pf�<�ׯ<�E�<a��<��<�{�<�ܧ<�:�<��<Y�<�C�<͖�<#�<5�<���<�ɘ<�<)V�<c��<�ڑ<g�<gX�<�<Њ<�	�<�B�<'z�<̰�<��<��<͟|<�y<bnu<��q<@:n<ޟj<yg<Kkc<��_<u8\<Z�X<F	U<jsQ<E�M<�LJ<)�F<�-C<ʡ?<w<<͑8<O5<�1<@.<�*<�"'<��#<�D <[�<�x<�<2�<�k<�<��<s�<*S<u8�;��;��;I<�;l�;���;��;	��;Ү�;���;���;}�;�J�;���;���;�d�;��;8q�;��;���;Z}�;�L�;KX~;�7t;#7j;VV`;��V;"�L;
rC;y:;y�0;5�';��;��;��;�(;�!�:�'�:gb�:���:r�:�D�:H�:3y�:�i:�J:a7,:�:��9b֤9�^T9>h�8�������u�lԲ��P�]��b�+��G���a�Ô|�����ఘ� å�:���ͨ���~̺pBٺ�����$*��R����{G��v������$���*���0�=7��&=�)6C��AI�9KO�	RU�nV[�iYa�TZg��Zm��Ys�*Xy��V���������1���/���ک��%���+���Z���級��  �  �i=�=��=9F=��=ق=� =f� =�[ =��</*�<�b�<��<���<��<X;�<Do�<���<���<+�<�3�<�a�<N��<˹�<���<>�<53�<�X�<<|�<'��<l��<���<'��<��<�+�<)B�<"V�<�g�<Uw�<S��<ݎ�<͖�<0��<���<���<���<���<���<���<�q�<_�<�I�<k0�<�<��<���<���<�~�<�P�<Y�<w��<���<q�<�/�<���<���<&S�<��<b��<S�<���<\��</�<�ž<�X�<��<�r�<���<Z}�< ��<y�<��<`f�<�ׯ<�E�<`��<��<�{�< ݧ<�:�<7��<c�<�C�<֖�<$�<5�<���<�ɘ<�<2V�<d��<�ڑ<h�<`X�<��<Њ<�	�<�B�<&z�<۰�<y�<��<��|<�y<;nu<��q<Z:n<ğj<�g<*kc<��_<�8\<7�X<G	U<YsQ<6�M<�LJ<B�F<�-C<ɡ?<s<<͑8<�5<��1<<.<�*<�"'<��#<�D <T�<�x<<-�<�k<�<��<��<S<�8�;���;��;d<�;6�;x��;���;��;���;о�;���;[�;�J�;���;���;�d�;��;�p�;h�;k��;.}�;M�;AX~;$8t;
7j;�V`;��V;�L;YrC;^:;��0;&�';��;e�;��;});�!�:�(�:b�:t��:�s�:�D�:�H�:	y�:g�i:��J:�5,:��:@�9PӤ9�YT9lx�8P������i�u�Ӳ��L깬����+��
G���a���|����������å�����4���c|̺�Aٺ*��s��*��������G��v������$��*�|�0�y7��%=��5C��AI�KO�RU��U[��Ya��Zg�[m��Ys��Xy��V�N���ᩅ����q����������o���Y���	����  �  �i=�=��=:F=��=ڂ=� =R� =�[ =��<0*�<�b�<��<���<��<];�<2o�<���<���<0�<~3�<�a�<S��<ƹ�<���<<�</3�<�X�<A|�<5��<j��<���<��<��<�+�< B�<%V�<�g�<]w�<d��<��<ז�<9��<Ȟ�<���<���<���<���<���<~q�<_�<vI�<o0�<�<��<���<���<�~�<~P�<X�<j��<���<�p�<n/�<���<���<)S�<��<k��<S�<���<n��<!/�<�ž<�X�<��<�r�<���<U}�<��<%y�<��<pf�<�ׯ<�E�<a��<��<�{�<�ܧ<�:�<��<Y�<�C�<͖�<#�<5�<���<�ɘ<�<)V�<c��<�ڑ<g�<gX�<�<Њ<�	�<�B�<'z�<̰�<��<��<͟|<�y<bnu<��q<@:n<ޟj<yg<Kkc<��_<u8\<Z�X<F	U<jsQ<E�M<�LJ<)�F<�-C<ʡ?<w<<͑8<O5<�1<@.<�*<�"'<��#<�D <[�<�x<�<2�<�k<�<��<s�<*S<u8�;��;��;I<�;l�;���;��;	��;Ү�;���;���;}�;�J�;���;���;�d�;��;8q�;��;���;Z}�;�L�;KX~;�7t;#7j;VV`;��V;"�L;
rC;y:;y�0;5�';��;��;��;�(;�!�:�'�:gb�:���:r�:�D�:H�:3y�:�i:�J:a7,:�:��9b֤9�^T9>h�8�������u�lԲ��P�]��b�+��G���a�Ô|�����ఘ� å�:���ͨ���~̺pBٺ�����$*��R����{G��v������$���*���0�=7��&=�)6C��AI�9KO�	RU�nV[�iYa�TZg��Zm��Ys�*Xy��V���������1���/���ک��%���+���Z���級��  �  �i=�=��=@F=��=ׂ=� =P� =�[ =	��<,*�<�b�<��<���<��<f;�<*o�<��<���<2�<�3�<�a�<f��<���<���<<�<(3�<�X�<1|�<7��<V��<���<��<��<�+�<B�<6V�<�g�<^w�<T��<��<Җ�<.��<̞�<���<���<���<���<���<�q�<1_�<lI�<v0�<��<��<���<���<�~�<xP�<a�<`��<���<q�<v/�<��<���<4S�<��<n��<S�<���<g��</�<�ž<�X�<��<�r�<���<a}�<��<%y�<��<rf�<�ׯ<�E�<]��<��<�{�<�ܧ<;�<��<m�<�C�<Ŗ�<,�<5�<���<�ɘ<�<(V�<c��<�ڑ<^�<�X�<<Њ<�	�<�B�<3z�<���<��<��<П|<ty<Qnu<��q<A:n<��j<Mg<ckc<��_<t8\<N�X<#	U<msQ<$�M<�LJ<�F<�-C<ɡ?<i<<�8<G5<4�1<2.<�*<�"'<��#<�D <K�<�x<�<D�<�k<�<��<j�<OS<E8�;0��;��;0<�;o�;M��;��;���;Ѯ�;���;���;��;�J�;���;���;�d�;��;q�;z�;a��;j}�;�L�;�X~;�7t;\7j;�V`;ЕV;��L;�qC;�:;T�0;N�';��;k�;��;�(;\"�:<'�:�c�:���:�r�:�E�:wG�:�y�:��i:Y�J:I6,:��:��9�Ѥ9_T9@i�8�b�����A�u��Ѳ��P�Z����+�|G���a��|�ȉ��/���v¥����ɧ���~̺7Aٺ?�庁��)�����m��G�iv�����$���*���0�z7��&=��5C��AI�LKO��QU��V[�>Ya��Zg��Zm�Zs�mXy��V�����w�����������ש��%���C�������ᴚ��  �  �i=�=��==F=��=ׂ=� =S� =�[ =��<2*�<�b�<��<���<��<e;�<5o�<���<���<)�<�3�<�a�<\��<���<���<;�<43�<�X�<9|�<?��<e��<���<!��<��<�+�<B�<)V�<�g�<^w�<Y��<��<��</��<Ҟ�<���<���<���<���<���<�q�<_�<sI�<t0�< �<��<���<���<�~�<�P�<^�<i��<���<�p�<v/�<���<���<-S�<��<u��<S�<���<q��</�<�ž<�X�<��<�r�<���<X}�<��<#y�<��<zf�<�ׯ<�E�<i��<��<�{�<�ܧ<�:�<��<[�<�C�<Ж�<%�<5�<���<�ɘ<�<0V�<_��<�ڑ<^�<gX�<�<Њ<�	�<�B�<,z�<̰�<��<��<�|<�y<Mnu<��q<>:n<ߟj<ng<Hkc<~�_<�8\<H�X<C	U<�sQ<&�M<�LJ<-�F<�-C<͡?<j<<ܑ8<T5<�1<+.<�*<�"'<��#<�D <>�<�x<�<2�<�k<�<��<x�<;S<_8�;"��; ��;_<�;|�;m��;��;��;ɮ�;���;���;r�;�J�;Ř�;���;�d�;��;6q�;��;f��;�}�;�L�;dX~;�7t;7j;�V`;��V;�L;�qC;�:;l�0;n�';��;]�;��;);("�:�'�:2b�:��:�r�:�D�:�G�:xy�:��i:A�J:�6,:��:t�9CԤ9�]T9�j�8ܒ�����?�u��Ӳ��O깭���+�dG�z�a���|��������¥�����s���M~̺XBٺ1��Җ��)��2�����G�Uv�ǟ���$���*���0�=7��&=��5C��AI�KO��QU�rV[�0Ya��Zg�bZm��Ys�Xy�sV���������H���6���婎�����N���a��������  �  �i=�=��=8F=��=܂=� =X� =�[ =��<.*�<�b�<��<���<��<Y;�<9o�<��<���<:�<�3�<�a�<S��<̹�<���<:�</3�<�X�<=|�<,��<e��<���<"��<��<�+�<%B�<#V�<�g�<Yw�<`��<ߎ�<֖�<+��<Ȟ�<���<���<���<���<���<�q�<_�<�I�<f0�<�<��<���<���<�~�<�P�<O�<x��<���<q�<z/�<���<���<!S�<��<k��<S�<���<`��</�<�ž<�X�<��<�r�<���<Z}�<��<y�<��<ff�<�ׯ<�E�<`��<��<�{�<�ܧ<�:�< ��<_�<�C�<ז�<�<5�<���<�ɘ<
�<2V�<]��<�ڑ<s�<hX�<���<Њ<�	�<�B�< z�<Ѱ�<��<��<Ɵ|<�y<Unu<��q<P:n<ןj<�g<Akc<��_<�8\<J�X<7	U<`sQ<4�M<�LJ<1�F<�-C<С?<�<<͑8<h5<�1<V.<�*<�"'<��#<�D <R�<�x<�<�<�k<<��<��<(S<�8�;��;���;J<�;B�;}��;ǻ�;���;���;���;���;x�;�J�;���;���;�d�;��;q�;��;U��;Y}�;�L�;X~;8t;97j;�V`;�V;?�L;~rC;5:;o�0;W�';͘;q�;��;);<!�:�(�:�b�:���:�r�:�D�:�H�:�x�:�i:�J:�5,:�::�9xդ9�[T9gr�8����?����u�dӲ�jN�5����+��	G�H�a�[�|��������Jå�ʾ��⨿��}̺Bٺ,��\���*�������G��v������$��*�#�0�77�w&=�
6C��AI�KO�CRU�NV[��Ya��Zg��Zm��Ys�^Xy�rV�a����������D���ũ������K���y��������  �  �i=�=��=>F=��=ւ=� =U� =�[ =
��<"*�<�b�<��<���<��<W;�<8o�<��<���<-�<�3�<�a�<Z��<���<���<@�<03�<�X�<B|�<9��<e��<���<��<��<�+�<B�<2V�<�g�<Pw�<^��<��<ۖ�<0��<ɞ�<���<���<���<���<���<�q�<!_�<pI�<k0�<�<��<���<���<�~�<�P�<Y�<c��<���<q�<v/�<���<���<,S�<��<n��<S�<���<h��</�<�ž<�X�<��<�r�<���<c}�<��<y�<��<qf�<�ׯ<�E�<c��<��<�{�<�ܧ<�:�<��<a�<�C�<�<)�<5�<���<�ɘ<
�<0V�<g��<�ڑ<_�<jX�<���<Њ<�	�<�B�</z�<Ͱ�<��<��<՟|<�y<Tnu<o�q<S:n<�j<[g<Rkc<��_<i8\<N�X<;	U<rsQ<?�M<�LJ<.�F<�-C<��?<e<<ߑ8<]5<	�1<4.<��*<�"'<��#<�D <h�<�x<�<C�<�k<�<��<��<8S<W8�;
��;��;N<�;M�;���;���;���;���;���;���;�;�J�;蘯;���;�d�;��;q�;��;j��;_}�;�L�;}X~;�7t;77j;�V`;ЕV;M�L;�qC;^:;��0;E�';ʘ;��;��;6);�!�:o'�:�b�:n��:�r�:9E�:�G�:fy�:��i:`�J:�5,:k�:�9�Ԥ9�XT9�r�8	n�����u��в��O�p���+��G���a��|�u���Ͱ��å�����q���*~̺�Aٺ��庳��)��
����PG��v�ɟ���$�Q�*���0�#7��&=��5C�BI�SKO��QU�iV[��Ya�qZg��Zm��Ys�cXy��V�\�������m���"�������<���C���p���״���  �  �i=�=��=;F=��=ւ=� =Q� =�[ =��<2*�<�b�<��<���<��<`;�<(o�<���<���<4�<�3�<�a�<`��<���<���<7�</3�<�X�<8|�<<��<c��<���<��<��<�+�<!B�<*V�<�g�<^w�<\��<��<ז�<+��<Ԟ�<���<���<���<���<���<~q�<(_�<sI�<u0�<��<��<���<���<�~�<vP�<]�<g��<���<�p�<t/�<��<���<3S�<��<x��<S�<���<m��</�<�ž<�X�<��<�r�<���<Y}�<��<(y�<��<vf�<�ׯ<�E�<g��<��<�{�<�ܧ<;�<��<^�<�C�<̖�<'�<�4�<���<�ɘ<�<'V�<Z��<�ڑ<c�<rX�<<Њ<�	�<�B�<.z�<Ű�<��<��<ן|<�y<Xnu<��q<8:n<�j<wg<Qkc<~�_<x8\<U�X<?	U<vsQ<*�M<�LJ< �F<�-C<ˡ?<e<<�8<L5<�1<>.<�*<�"'<��#<�D <T�<�x<�<7�<�k<<��<r�<CS<S8�;0��;��;I<�;r�;f��;��;��;߮�;���;���;��;�J�;Ƙ�;���;�d�;��;,q�;��;T��;�}�;�L�;�X~;�7t;b7j;�V`;��V;��L;�qC;�:;-�0;E�';�;x�;��;�(;!"�:�'�:c�:��:xr�:�E�:yG�:�y�:��i:��J:�5,:��:a�9Ԥ9�^T9Ue�8������͵u��Ӳ�Q���P�+��G��a�R�|�4���b���{¥�쿲�
����~̺&BٺY�����)��������G�vv����$���*���0��7��&=��5C�BI�<KO��QU��V[�,Ya��Zg��Zm��Ys�SXy��V���������5���$���穎����4���i���Ѵ���  �  �i=�=��=8F=��=ق=� =W� =�[ =��<-*�<�b�<��<���<~�<e;�<5o�<��<���<2�<�3�<�a�<U��<ƹ�<���<6�<+3�<�X�<@|�<4��<_��<���<'��<��<�+�<*B�<&V�<�g�<^w�<T��<��<ܖ�<0��<͞�<���<���<���<���<���<�q�<"_�<uI�<i0�<��<��<���<���<�~�<�P�<Q�<i��<���<q�<s/�<���<���<+S�<��<q��<S�<���<g��</�<�ž<�X�<��<�r�<���<[}�<��<y�<��<nf�<�ׯ<�E�<b��<��<�{�<�ܧ<�:�<��<`�<�C�<̖�<�<5�<���<�ɘ<�<2V�<X��<�ڑ<e�<oX�<���<Њ<�	�<�B�<%z�<ư�<��<��<ן|<~y<=nu<��q<T:n<ϟj<�g<<kc<��_<�8\<6�X<4	U<psQ<;�M<�LJ<!�F<�-C<ڡ?<q<<Б8<b5<�1<;.<�*<�"'<��#<�D <8�<�x<�<�<�k<�<��<��<,S<u8�;-��;��;<<�;e�;���;��;ݭ�;���;Ͼ�;���;o�;�J�;���;���;�d�;��;q�;��;h��;n}�;�L�;YX~;�7t;07j;�V`;ՕV;W�L;�qC;N:;d�0;��';��;E�;��;);b!�:�'�:�b�:p��:`r�:E�:H�:Yy�:x�i:��J:E6,:i�:��9�Ҥ9y]T9u�8���������u��Ҳ��M�m����+��G� �a�i�|�~���;����¥�e�������~̺Bٺ������*��&��m��G�v�����$��*���0��7��&=�6C��AI��JO�RU��V[�ZYa�|Zg��Zm��Ys��Xy�PV�Z���˩�����N�������񪑻s���~���ܴ���  �  �i=�=��=;F=��=ق=� =T� =�[ =��<**�<�b�<��<���<��<Z;�<5o�<���<���<.�<|3�<�a�<U��<ɹ�<���<A�<53�<�X�<D|�<1��<s��<���<��<��<�+�< B�<&V�<�g�<Nw�<i��<��<ۖ�<5��<ƞ�<���<���<���<���<���<�q�<_�<xI�<m0�<�<��<���<���<�~�<�P�<V�<m��<���< q�<q/�<���<���<"S�<��<k��<S�<���<k��<)/�<�ž<�X�<��<�r�<���<]}�<��<y�<��<lf�<�ׯ<�E�<f��<��<�{�<�ܧ<�:�<��<Z�<�C�<Ζ�<$�<5�<���<�ɘ<�<,V�<c��<�ڑ<d�<cX�<���<Њ<�	�<�B�<(z�<԰�<��<��<П|<�y<anu<v�q<X:n<ԟj<ug<Akc<��_<u8\<R�X<S	U<hsQ<E�M<�LJ<<�F<�-C<š?<s<<ϑ8<W5<��1<9.<
�*<�"'<��#<�D <_�<�x<�<:�<�k<�<��<v�<,S<�8�;���;��;c<�;P�;���;ػ�;-��;���;���;���;q�;�J�;���;���;�d�;��;1q�;��;}��;R}�;�L�;)X~;�7t;7j;nV`;��V;	�L;rC;j:;��0;5�';ݘ;��;v�;);�!�:(�:.b�:N��:Br�:�D�:&H�:�x�:��i:��J:�6,:��:��97ؤ9�WT9�r�8
������o�u�}Ҳ�bO�ʫ�2�+�D	G���a���|�I��������å����Ĩ��o~̺fBٺ�����*��&����vG��v�����$�(�*���0�]7��&=�6C��AI�5KO�RU�5V[��Ya�\Zg��Zm�wYs�.Xy��V�R�������9���C�������$���:���A���봚��  �  �i=�=��=;F=��=ق=� =Q� =�[ =��<+*�<�b�<��<���<��<_;�<,o�<���<���<6�<�3�<�a�<_��<Ĺ�<���<=�</3�<�X�<;|�<0��<_��<���<��<��<�+�<B�<.V�<�g�<\w�<`��<ێ�<Ֆ�<.��<˞�<���<���<���<���<���<�q�<-_�<uI�<q0�<��<��<���<���<�~�<{P�<[�<i��<���<q�<}/�<��<���<-S�<��<k��<S�<���<_��</�<�ž<�X�<��<�r�<���<_}�<��<'y�<��<if�<�ׯ<�E�<a��<��<�{�<�ܧ<;�<��<g�<�C�<ǖ�<)�<5�<���<�ɘ<�<(V�<c��<�ڑ<e�<uX�<<Њ<�	�<�B�<*z�<ǰ�<��<��<Ο|<vy<]nu<��q<Q:n<�j<bg<Zkc<��_<8\<U�X<*	U<esQ<2�M<�LJ<$�F<�-C<ӡ?<r<<�8<I5<�1<B.<�*<�"'<��#<�D <K�<�x<�<;�<�k<<��<r�<AS<l8�;��;��;I<�;_�;t��;Ի�;ۭ�;ܮ�;���;���;��;�J�;Ԙ�;���;�d�;��;�p�;��;b��;g}�;�L�;pX~;�7t;a7j;�V`;V;��L;rC;�:;O�0;>�';��;]�;��;�(;�!�:�'�:_c�:���:s�:oE�:�G�:yy�:|�i:
�J:*6,:��:��9�Ԥ9_T9�p�8����J���u�Ҳ�MO�8����+��	G���a���|����������¥�s���&���P~̺�Aٺ8��Y���)��s�����G��v�����$��*���0��7��&=��5C��AI�!KO��QU��V[�JYa��Zg��Zm�Zs�?Xy��V�`�������`�������������4�������𴚻�  �  �i=�=��=;F=��=҂=� =O� =�[ =��<.*�<�b�<��<���<w�<k;�<,o�<���<���<*�<3�<�a�<]��<���<���<6�<13�<�X�<8|�<H��<]��<���<!��<��<�+�<B�<1V�<�g�<cw�<V��<��<��<*��<מ�<���<���<���<���<���<xq�<$_�<gI�<t0�<��<��<���<���<�~�<yP�<^�<]��<���<�p�<x/�<���<���<4S�<��<x��<S�<���<t��</�<�ž<�X�<��<�r�<���<Y}�<��<(y�<��<�f�<�ׯ<�E�<g��<��<�{�<�ܧ<�:�<��<Y�<�C�<Ė�<&�<5�<���<�ɘ<�<.V�<Z��<�ڑ<V�<mX�<锌<Њ<�	�<�B�<.z�<°�<��<��<��|<�y<Inu<��q<;:n<�j<og<Skc<~�_<�8\<G�X<4	U<�sQ<%�M<�LJ< �F<�-C<ݡ?<X<<�8<D5<
�1<".<�*<�"'<��#<�D <*�<�x<�<0�<�k<�<��<r�<<S<;8�;>��;��;T<�;u�;h��;4��;խ�;Ԯ�;���;���;��;�J�;ᘯ;���;�d�;��;:q�;��;S��;�}�;�L�;�X~;�7t;7j;�V`;W�V;d�L;�qC;�:;9�0;��';��;0�;��;�(;."�:'�:�b�:���:�r�:�D�:~G�:�y�:��i:��J:�5,:)�:�9~Ҥ9GaT9�g�8���c��X�u�tӲ��O���)�+��G�M�a�4�|�8���d���N¥�!���n���b~̺{Bٺ��应���)��o��G�%H�Sv�؟�	�$���*��0�7�'=��5C�4BI�
KO��QU��V[��Xa��Zg�%Zm��Ys��Xy�TV���������G������橎�󪑻P���~��������  �  �i=�=��=:F=��=ׂ=� =X� =�[ =��<2*�<�b�<��<���<��<];�<-o�<���<���<8�<3�<�a�<W��<Ź�<���<9�<23�<�X�<9|�<0��<h��<���<#��<��<�+�<&B�<(V�<�g�<Yw�<^��<��<Ԗ�<)��<Ȟ�<���<���<���<���<���<�q�<$_�<{I�<t0�<��<��<���<���<�~�<yP�<]�<p��<���< q�<�/�<���<���<*S�<��<l��<S�<���<c��</�<�ž<�X�<��<�r�<���<W}�<��<!y�<��<jf�<�ׯ<�E�<b��<��<�{�<�ܧ<�:�<#��<[�<�C�<Ӗ�<&�<5�<���<�ɘ<�<(V�<Y��<�ڑ<j�<kX�<���<Њ<�	�<�B�<)z�<ΰ�<��<��<̟|<�y<Wnu<��q<J:n<ܟj<~g<Ekc<��_<�8\<Q�X<=	U<isQ<-�M<�LJ<1�F<�-C<ʡ?<k<<ߑ8<e5<�1<F.<�*<�"'<��#<�D <T�<�x<�<2�<�k<<��<��<1S<s8�;��;���;U<�;:�;i��;Ի�;���;ɮ�;���;���;}�;�J�;���;���;�d�;��;q�;��;N��;Y}�;�L�;YX~;�7t;7j;�V`;̕V;c�L;/rC;�:;=�0;"�';И;g�;��;�(;"�:4(�:c�:H��:*s�:�D�:+H�:=y�:��i:)�J:85,:S�:��9�Ԥ9�\T9l�8P������u��Ӳ��N�ݪ���+��	G��a�ǖ|��������å�M��������}̺MBٺ�废���)��o�����G��v����$���*�k�0�!7��&=��5C��AI�%KO��QU�eV[��Ya��Zg��Zm��Ys�WXy��V�n�������'���<���ϩ�����<���l���괚��  �  �h=�=��=E=l�=r�=-=�� =�Y =��<�%�<�]�<3��<|��<� �<p5�<�h�<a��<���<���<�+�<�Y�<օ�<��<s��<��<)�<�M�<Fq�<���<���<`��<\��<S�<)�<�3�<vG�<�X�<�g�<<t�<=~�<���<���<���<��<{��<��<�x�<%l�<�\�<�I�<�3�<�<O��<��<'��<���<�f�<8�<��<q��<v��<�W�<��<?��<ǆ�<B9�<���<���<)9�<���<�z�<~�<U��<q?�<�λ<�Y�<f�<3e�<K�<�a�<�ڲ<�O�<���< 0�<L��<-�<�g�<�ɧ<(�<䃤<�ܢ<�2�<~��<�ם<&�<Qr�<S��<)�<J�<���<Б<w�<0O�<|��<PȊ<��<Z<�<�t�<��<��<M�<Ś|<y<blu<�q<o;n<\�j<�	g<�pc<��_<A\<]�X<�U<l�Q<��M<�\J<��F<�@C<T�?<d.<<7�8<C'5<`�1<-.<E�*<zA'<��#<f </�<Ӝ<{?<�<�<�F<|�<w�<;�<���;�5�;���;H��;h�;?�;$�;�;&�;�+�;L�;�{�;��;�	�;�h�;	פ;�U�;^�;�;�1�;���;��;�=;�u;kk;}8a;vW;��M;5ND;��:;��1;�v(;�i;Wz;�;��;\��:��:���:KB�:z۵:T��:͠�:BɅ:9Bl:�GM:�.:�S:��9�L�9� ]9%G�8��*�#����n��!���湸��OK*��pE�2^`��{��Ҋ�[��������Q����˺5�غ�l庾򺘮��e��������D�p��$��*���0���6��=��C��#I�[/O��8U�?[��Da��Gg��Jm�?Ks�Ly��L�A���অ�T�������ܩ��p�������˳�������  �  �h=�=��=E=j�=t�=7=�� =�Y =��<�%�<�]�<*��<���< �<{5�<�h�<d��<���<���<�+�<�Y�<��<��<w��<��<)�<N�<Eq�<В�<���<d��<S��<I�<,�<�3�<xG�<�X�<�g�<5t�<A~�<���<���<���< ��<���<��<�x�<0l�<�\�<�I�<�3�<)�<K��< ��<5��<ϑ�<�f�<8�<��<k��<w��<�W�<��<N��<ņ�<H9�<���<��<'9�<���<�z�<x�<^��<b?�<�λ<�Y�<f�<,e�<?�<�a�<�ڲ<�O�<���<#0�<F��<#�<�g�<�ɧ<*(�<⃤<�ܢ<�2�<{��<�ם<&�<Wr�<\��<:�<J�<���<Б<l�<6O�<{��<cȊ<��<W<�<�t�<	��<��<K�<�|<y<_lu<	�q<P;n<j�j<�	g<�pc<��_<A\<]�X<�U<��Q<��M<�\J<��F<�@C<K�?<j.<<a�8<A'5<j�1<-.<R�*<}A'<��#<<f <?�<�<j?<#�<�<vF<�<p�<c�<��;�5�;���;-��;h�;?�;Q$�;��;4�;u+�;�K�;�{�;��;�	�;�h�;%פ;�U�;m�;!��;�1�;���;޿�;>;�u;�k;�8a;�uW;��M;�MD;N�:;f�1;�v(;Vj;�z;��;K�;��:���:���:B�:�۵:A��:���:�Ʌ:�@l:�GM:��.:�T:��9FK�9+]9e8�8��*������n��#��k�����L*�6oE��]`�>{��Ҋ� ��W�����.����˺H�غ�l���X���������c�D�Np���$���*���0���6��=�2C��#I�z/O��8U�q?[�mDa�Hg�Jm�YKs�%Ly��L����Ŧ��M���e������s�������ݳ��G����  �  �h=�=��="E=k�=m�=4=�� =�Y =��<�%�<�]�<(��<���<� �<}5�<�h�<j��<���<���<�+�<}Y�<��<ذ�<��<��<)�<N�<@q�<Ԓ�<~��<l��<Y��<M�<3�<�3�<�G�<�X�<�g�</t�<=~�<���<���<���<���<���<��<�x�<(l�<�\�<�I�<�3�</�<M��<��<.��<Ƒ�<�f�<8�<��<f��<~��<�W�<��<F��<���<U9�<���<���<,9�<���<�z�<p�<m��<c?�<�λ<�Y�<g�<3e�<C�<�a�<ڲ<�O�<���<.0�<L��<&�<�g�<xɧ<&(�<ۃ�<�ܢ<�2�<z��<�ם<&�<Yr�<L��<7�<	J�<���<Б<i�<DO�<t��<\Ȋ<��<W<�<�t�<��<��<H�<�|<�y<^lu<�q<N;n<��j<s	g<�pc<��_<A\<a�X<�U<��Q<��M<�\J<��F<�@C<N�?<O.<<V�8<0'5<��1<-.<W�*<�A'<��#<:f <�<�<k?</�<�<qF<��<_�<[�<���;�5�;���;2��;Ph�;?�;`$�;��;V�;�+�;L�;�{�;躵;
�;�h�;aפ;�U�;]�;+��;�1�;�;ֿ�;x>;Uu;|k;�8a;�uW;��M;�MD;~�:;v�1;�v(;j;z;��;K�;5��:f��:��:B�:l۵:���:��:oʅ:�@l:�HM:S�.:�T:��97I�9�]9L9�8U�*�]���=n��!����湢���M*��nE�l^`��{�~Ҋ����������r���˺޳غ�l��� �����������4D�^p�ؖ$�|�*��0�[�6�=�fC�-$I�x/O�<8U��?[�Da�%Hg��Im��Ks�)Ly�QL���������}���9������Q����������:����  �  �h=�=��=E=k�=s�=3=�� =�Y =��<�%�<�]�<0��<���<� �<|5�<�h�<`��<���<���<�+�<�Y�<��<��<u��<��<)�<N�<Bq�<Β�<���<i��<V��<C�<0�<�3�<{G�<�X�<�g�<9t�<>~�<���<���<���<��<��<��<�x�<(l�<�\�<�I�<�3�<#�<N��<��</��<ˑ�<�f�<8�<��<r��<p��<�W�<��<G��<ǆ�<H9�<���<��<+9�<���<�z�<z�<`��<a?�<�λ<�Y�<g�<*e�<@�<�a�<�ڲ<�O�<���<%0�<B��<%�<�g�<�ɧ<#(�<���<�ܢ<�2�<���<�ם<&�<Zr�<Y��<5�<J�<���<	Б<t�<2O�<z��<\Ȋ<��<Y<�<�t�<��<��<O�<ښ|<y<jlu<�q<K;n<q�j<u	g<�pc<��_<
A\<h�X<�U<~�Q<��M<�\J<��F<�@C<L�?<g.<<S�8<?'5<g�1<-.<D�*<vA'<��#<9f <;�<�<u?<�<�<sF<��<m�<T�<��;�5�;���;��;%h�;?�;H$�;��;I�;�+�;�K�;�{�;���;�	�;�h�;-פ;�U�;`�;	��;�1�;���;ῄ;>;�u;�k;�8a;�uW;��M;!ND;�:;��1;�v(;%j;�z;��;y�;y��:&��:A��:�A�:s۵:֥�:ʠ�:�Ʌ:Al:�GM:L�.:�S:R��9�K�9]9i7�8��*�q���Vn�$��N�湢��,L*�YoE��^`��{�*ӊ����o����������˺S�غm庇򺦮��������|�ED�!p���$��*���0���6��=�hC��#I�i/O��8U��?[�^Da��Gg�6Jm�rKs��Ky��L���������y���X���&���i�������޳��^����  �  �h=�=��=E=g�=u�=0=�� =�Y =��<�%�<�]�<*��<���<�<m5�<�h�<\��<���<���<�+�<�Y�<م�<��<n��<��<)�< N�<Nq�<ǒ�<���<^��<Z��<G�<-�<�3�<vG�<�X�<�g�<6t�<9~�<���<���<���<��<y��<��<�x�<*l�<�\�<�I�<�3�<!�<O��<���<0��<͑�<�f�<8�<��<~��<k��<�W�<��<E��<̆�<@9�<���<x��</9�<���<�z�<x�<Z��<j?�<�λ<�Y�<h�<*e�<F�<�a�<�ڲ<�O�<���<%0�<A��<0�<�g�<�ɧ<(�<僤<�ܢ<�2�<���<~ם<&�<Kr�<_��</�<	J�<���<Б<}�<(O�<���<WȊ<��<U<�<�t�<��<��<Y�<ך|<	y<Ulu<�q<Y;n<g�j<�	g<�pc<��_<A\<P�X<�U<x�Q<��M<�\J<��F<�@C<?�?<o.<<D�8<U'5<U�1<-.<S�*<wA'<��#<&f <I�<͜<q?<�<�<{F<w�<~�<B�<��;�5�;���;&��;h�;;?�;-$�;��;�;�+�;�K�;�{�;#��;�	�;�h�;פ;�U�;N�;��;2�;���;��;�=;�u;�k;�8a;%vW;F�M;�ND;�:;��1;jv(;+j;�z;C�;��;.��:ب�:���:OB�:�۵:���:��:,Ʌ:�Bl:�FM:��.:�T:4��9\K�9a]9�?�8d+������n�6$����湕���K*�(pE�]`�{�*ӊ�(�����G������˺[�غ	m�1�����|����J�uD�ap��$���*�u�0�3�6��=��C��#I��/O��8U�?[��Da��Gg�?Jm�}Ks�NLy��L�n���ʦ��2���k������f�������۳��j����  �  �h=�=��=!E=k�=t�=0=�� =�Y =��<�%�<�]�</��<���<� �<w5�<�h�<e��<���<���<�+�<�Y�<߅�<��<v��<��<)�<N�<Dq�<ʒ�<���<h��<]��<N�<'�<�3�<{G�<�X�<�g�<3t�<>~�<���<���<���<��<���<��<�x�<+l�<�\�<�I�<�3�<'�<S��< ��<.��<Ǒ�<�f�<8�<��<r��<t��<�W�<��<I��<Ć�<M9�<���<{��<+9�<���<�z�<u�<f��<e?�<�λ<�Y�<a�<1e�<G�<�a�<�ڲ<�O�<���<&0�<C��<-�<�g�<�ɧ<"(�<䃤<�ܢ<�2�<~��<�ם<&�<Ur�<R��<7�<J�<���<Б<m�<6O�<}��<WȊ<��<Y<�<�t�<��<��<M�<ۚ|<y<Wlu<�q<T;n<h�j<u	g<�pc<��_<A\<[�X<�U<|�Q<��M<�\J<��F<�@C<N�?<l.<<E�8<G'5<l�1<-.<T�*<�A'<��#<8f <)�<�<�?<'�<�<pF<��<{�<N�<��;�5�;���;"��;*h�;?�;:$�;��;F�;�+�;L�;�{�;ẵ;�	�;�h�;Mפ;�U�;b�;��;�1�;���;���;A>;�u;�k;�8a;'vW;��M;ND;>�:;��1;�v(;j;�z;��;��;���:��:���:�B�:�۵:���:���:�Ʌ:nAl:GM:2�.:&T:��9�J�9�	]9�;�8a�*�#���%n�_"��V��J��|L*��oE�-^`��{�ӊ�\��]����������˺�غm庸�V���N�������8D�3p�Ö$���*���0���6��=��C��#I�b/O�i8U�D?[��Da��Gg�/Jm�bKs�CLy�VL�x���Ȧ��x���{������J�������ڳ��a����  �  �h=�=��=E=i�=s�=7=�� =�Y =��<�%�<�]�<+��<���<� �<�5�<�h�<c��<���<���<�+�<Y�<��<ݰ�<r��<��<)�<	N�<:q�<Ғ�<���<k��<Q��<J�<2�<�3�<�G�<�X�<�g�<3t�<C~�<���<���<���<���<���<��<�x�<,l�<~\�<�I�<�3�<+�<E��<��<2��<ʑ�<�f�<8�<��<p��<x��<�W�<��<P��<���<N9�<���<���<*9�<���<�z�<u�<f��<Y?�<�λ<�Y�<i�</e�<9�<�a�<�ڲ<�O�<���<(0�<I��< �<�g�<{ɧ</(�<܃�<�ܢ<�2�<���<�ם<&�<br�<Q��<<�<J�<�<Б<m�<;O�<p��<aȊ<��<S<�<�t�<��<��<J�<ښ|<y<^lu<�q<H;n<��j<u	g<�pc<��_<A\<c�X<�U<��Q<��M<�\J<��F<�@C<E�?<f.<<a�8<-'5<q�1<-.<[�*<tA'<��#<If <(�<��<e?<!�<�<~F<�<b�<k�<̔�;�5�;���;,��;?h�;�>�;X$�;��;P�;n+�;�K�;�{�;뺵;
�;jh�;Cפ;�U�;v�;���;�1�;�;ο�;.>;/u;�k;�8a;�uW;��M;ND;^�:;9�1;�v(;>j;�z;ǧ;�; ��:���:���:�A�:�۵:b��:ݟ�:ʅ:@l:�HM:+�.:WS:���9oJ�9,	]9u/�8L�*�����:n��"�����)��M*��nE�W_`��{��Ҋ�-��k��r������˺r�غ�l府�S���ל�^����	D�@p��$���*���0���6�8=�>C��#I��/O��8U��?[�Da�Hg�4Jm�\Ks�'Ly��L���������y���<������l�������賗�T����  �  �h=�=��=E=m�=s�=1=�� =�Y =��<�%�<�]�<.��<���<� �<x5�<�h�<h��<���<���<�+�<�Y�<݅�<��<z��<��<)�<N�<Hq�<̒�<���<g��<]��<K�<-�<�3�<{G�<�X�<�g�<3t�<=~�<���<���<���<��<���<��<�x�<*l�<�\�<�I�<�3�<*�<S��<��<,��<Ƒ�<�f�<8�<��<q��<r��<�W�<��<F��<Æ�<L9�<���<~��</9�<���<�z�<v�<a��<i?�<�λ<�Y�<e�<-e�<G�<�a�<�ڲ<�O�<���<%0�<G��<*�<�g�<�ɧ<(�<ރ�<�ܢ<�2�<~��<�ם<&�<Vr�<O��</�<J�<���<Б<t�<4O�<y��<ZȊ<��<^<�<�t�<��<��<W�<ښ|<y<Wlu<�q<`;n<i�j<t	g<�pc<��_<A\<\�X<�U<�Q<��M<�\J<��F<�@C<V�?<g.<<H�8<;'5<i�1<-.<S�*<�A'<��#<+f <(�<�<s?<+�<�<{F<��<g�<J�<���;�5�;���;3��;h�;#?�;B$�;��;C�;�+�;�K�;�{�;�;�	�;�h�;<פ;�U�;^�;��;�1�;���;�;&>;�u;�k;�8a;�uW;��M;ND;W�:;��1;�v(;j;|z;��;��;���:��:c��:,B�:�۵:ƥ�:���:�Ʌ:�Al:}GM:��.:�T:��9�J�9�]93?�8#�*������n�]#��|�湟���L*��oE��]`��{��Ҋ����"����������˺,�غ�l庵������������rD�&p���$���*���0���6��=�vC��#I�B/O��8U�a?[��Da��Gg�4Jm��Ks�DLy�lL�_���Ǧ��z���g�������Y�����������[����  �  �h=�=��=E=k�=v�=/=�� =�Y =��<�%�<�]�<+��<���<�<v5�<�h�<_��<���<���<�+�<�Y�<څ�<��<q��<��<)�<N�<Nq�<���<���<c��<W��<E�<'�<�3�<pG�<�X�<�g�<<t�<9~�<���<���<���<��<z��<��<�x�<+l�<�\�<�I�<�3�< �<T��<���<3��<Б�<�f�<8�<��<v��<o��<�W�<��<B��<̆�<A9�<���<y��<.9�<���<�z�<��<Y��<f?�<�λ<�Y�<d�<'e�<B�<�a�<�ڲ<�O�<���<%0�<E��<,�<�g�<�ɧ<(�<胤<�ܢ<�2�<���<�ם<&�<Qr�<a��<6�<
J�<���<Б<t�<0O�<���<VȊ<��<^<�<�t�<��<��<Z�<̚|<y<clu<�q<P;n<U�j<�	g<�pc<��_<A\<`�X<�U<k�Q<��M<�\J<��F<�@C<P�?<r.<<B�8<S'5<b�1<-.<E�*<{A'<��#<6f <L�<ߜ<{?<�<�<qF<��<~�<D�<��;�5�;���;-��;#h�;=?�;$�;�;1�;�+�;�K�;�{�;��;�	�;�h�;פ;�U�;P�;��;�1�;���;��;�=;�u;�k;�8a;3vW;u�M;OND;�:;��1;�v(;Ij;�z;d�;��;?��:X��:-��:uB�:�۵:���:��:2Ʌ:�Bl:�FM:��.:9T:b��9jM�9�]9,<�8�>+�v����n��$�����M��K*�qE�M]`��{��Ҋ�n�����Z����U�˺*�غ;m庚�̮��[�����7�9D�Yp���$��*���0���6��=��C��#I�B/O��8U�#?[��Da��Gg�jJm�XKs�Ly��L����礪�6����������p�������ɳ�������  �  �h=�=��=E=i�=p�=3=�� =�Y =��<�%�<�]�<%��<���<� �<{5�<�h�<_��<���<���<�+�<�Y�<��<ݰ�<s��<��<)�<N�<Dq�<ɒ�<���<a��<V��<N�<,�<�3�<~G�<�X�<�g�<6t�<<~�<���<���<���<��<���<��<�x�<*l�<�\�<�I�<�3�<&�<L��<���<0��<ʑ�<�f�<8�<��<u��<t��<�W�<��<H��<���<H9�<���<~��<)9�<���<�z�<w�<^��<e?�<�λ<�Y�<e�<1e�<B�<�a�<�ڲ<�O�<���<$0�<D��<+�<�g�<}ɧ<%(�<ރ�<�ܢ<�2�<���<�ם<&�<Wr�<T��<9�<J�<���<Б<r�<7O�<x��<ZȊ<��<U<�<�t�<��<��<P�<ٚ|<y<Tlu<�q<W;n<q�j<�	g<�pc<��_<A\<P�X<�U<|�Q<��M<�\J<��F<�@C<H�?<Z.<<R�8<<'5<k�1<-.<]�*<xA'<��#<?f <*�<�<l?<�<�<vF<��<i�<Z�<˔�;�5�;���;!��;,h�;?�;3$�;��;(�;�+�;L�;�{�;��;�	�;�h�;*פ;�U�;X�;��;�1�;���;���;>;ju;�k;�8a;�uW;��M;8ND;6�:;r�1;�v(;0j;�z;��;b�;���:T��:{��:�A�:�۵:⥥:h��:�Ʌ:�Al:nGM:�.:�S:���9K�97]9D;�8i�*�:���`n�V"��ÿ�&��{L*��oE��^`�{�ӊ�x�����G��}����˺:�غ�l�<򺥮����������"D�|p���$���*���0���6��=�zC�$I��/O��8U�Z?[�qDa��Gg�7Jm�Ks�QLy��L�q�������U���_�������l�������೗�a����  �  �h=�=��= E=l�=q�=8=�� =�Y =��<�%�<�]�<,��<���<� �<�5�<�h�<i��<���<���<�+�<|Y�<��<ݰ�<���<��<)�<N�<@q�<ڒ�<��<m��<Y��<G�<.�<�3�<}G�<�X�<�g�<-t�<B~�<���<���<���<���<���<��<�x�<0l�<�\�<�I�<�3�<0�<N��<��<0��<ɑ�<�f�<8�<��<k��<x��<�W�<��<S��<���<T9�<���<}��<(9�<���<�z�<l�<i��<^?�<�λ<�Y�<e�<,e�<B�<�a�<|ڲ<�O�<���<%0�<>��<%�<�g�<|ɧ<0(�<ك�<�ܢ<�2�<|��<�ם<&�<_r�<P��<>�<J�<���<Б<g�<>O�<t��<eȊ<��<Y<�<�t�<���<��<I�<�|<y<Tlu<�q<M;n<r�j<d	g<�pc<��_<A\<\�X<�U<��Q<��M<�\J<��F<�@C<T�?<_.<<f�8</'5<}�1<�,.<Z�*<�A'<��#<Mf <&�<��<m?</�<�<iF<��<^�<n�<˔�; 6�;���;��;.h�;?�;y$�;��;Z�;�+�;�K�;�{�;׺�;�	�;h�;Tפ;�U�;q�;��;�1�;���;Ŀ�;v>;iu;�k;�8a;�uW;��M;�MD;��:;��1;�v(;-j;�z;ѧ;m�;_��:���:���:\B�:�۵:���:M��:lʅ:K@l:^GM:�.:T:���98H�9]9�4�8 �*�T���2n��#����湨��
N*��mE��^`��{�aӊ�������\�����;�˺��غ$m���ۭ�����w�����C�0p�ؖ$�}�*�"�0���6�=�!C��#I�h/O�Q8U��?[�UDa�"Hg��Im��Ks�QLy�KL�������������^������K�����������,����  �  �h=�=��=E=h�=s�=2=�� =�Y =��<�%�<�]�<,��<���<� �<w5�<�h�<^��<���<���<�+�<Y�<��<��<t��<��<)�<N�<Fq�<͒�<���<g��<U��<H�<1�<�3�<|G�<�X�<�g�<.t�<?~�<���<���<���<��<���<��<�x�<'l�<�\�<�I�<�3�<%�<L��< ��<1��<ˑ�<�f�<8�<��<u��<w��<�W�<��<I��<���<H9�<���<���<09�<���<�z�<n�<e��<_?�<�λ<�Y�<k�<+e�<>�<�a�<�ڲ<�O�<���<+0�<H��<*�<�g�<ɧ<%(�<ۃ�<�ܢ<�2�<���<�ם<&�<Sr�<Y��<6�<J�<�<Б<t�<:O�<x��<XȊ<��<R<�<�t�<��<��<R�<ך|<	y<Wlu<�q<M;n<o�j<�	g<�pc<��_<A\<[�X<�U<}�Q<��M<�\J<��F<�@C<D�?<e.<<M�8<8'5<u�1<-.<S�*<rA'<��#<7f <=�<�<p?<�<�<~F<��<c�<W�<ߔ�;�5�;���;5��;Ih�;?�;C$�;��;B�;�+�;�K�;�{�;��;�	�;�h�;@פ;�U�;f�;��;�1�;���;���;#>;Ou;�k;�8a;vW;��M;=ND;0�:;o�1;�v(;3j;�z;�;b�;���:M��:���:hB�:R۵:���:6��:�Ʌ:�Al:CHM:ڤ.:�S:��9�H�9�]9a5�8��*�����/n��#�����h��EM*�=oE�'^`�.{��Ҋ�������,������˺سغ�l应򺿮��������|�@D�Bp��$���*���0���6��=��C��#I��/O�|8U�b?[�:Da��Gg�>Jm�~Ks�FLy�yL���������J���^������^�������򳗻_����  �  �h=�=��= E=j�=w�=0=�� =�Y =��<�%�<�]�<8��<���<� �<r5�<i�<Y��<���<���<�+�<�Y�<���<��<r��<��<)�<�M�<Hq�<Ȓ�<���<^��<W��<O�<"�<�3�<xG�<�X�<�g�<3t�<C~�<���<���<���<��<|��<��<�x�<&l�<�\�<�I�<�3�<�<X��<��<1��<ˑ�<�f�<8�<��<{��<m��<�W�<��<K��<Ȇ�<A9�<���<u��<+9�<���<�z�<t�<]��<g?�<�λ<�Y�<]�</e�<B�<�a�<�ڲ<�O�<���<0�<>��<.�<�g�<�ɧ<"(�<ރ�<�ܢ<�2�<���<{ם<%&�<Pr�<Y��<0�<J�<���<
Б<y�<+O�<{��<RȊ<��<X<�<�t�<	��<��<V�<Қ|<y<Qlu<�q<^;n<W�j<|	g<�pc<��_<A\<N�X<�U<t�Q<��M<�\J<��F<�@C<K�?<x.<<C�8<?'5<W�1<-.<O�*<vA'<��#<&f <:�<ל<�?<�<�<�F<l�<g�<Q�<��;�5�;���;��;h�;"?�;/$�;��;�;�+�;L�;�{�;캵;�	�;�h�;,פ;�U�;u�;��;�1�;���;���;�=;�u;�k;�8a;�uW;W�M;kND;��:;Ѡ1;�v(;6j;�z;��;��;��:���:��:�A�:n۵:��:⠕:;Ʌ:�Al:UFM:N�.:WT:n��9aJ�9]9=�8)�*�����an��"����湡��L*��oE��]`��{�_ӊ�O�����a�������˺��غ�l�.�$��������|�mD��o��$�Ѹ*���0��6��=��C��#I�k/O��8U�s?[��Da��Gg�SJm�MKs�\Ly��L�c���ꦅ�j�������祈�f�������ҳ��q����  �  �h=�=��=E=h�=s�=2=�� =�Y =��<�%�<�]�<,��<���<� �<w5�<�h�<^��<���<���<�+�<Y�<��<��<t��<��<)�<N�<Fq�<͒�<���<g��<U��<H�<1�<�3�<|G�<�X�<�g�<.t�<?~�<���<���<���<��<���<��<�x�<'l�<�\�<�I�<�3�<%�<L��< ��<1��<ˑ�<�f�<8�<��<u��<w��<�W�<��<I��<���<H9�<���<���<09�<���<�z�<n�<e��<_?�<�λ<�Y�<k�<+e�<>�<�a�<�ڲ<�O�<���<+0�<H��<*�<�g�<ɧ<%(�<ۃ�<�ܢ<�2�<���<�ם<&�<Sr�<Y��<6�<J�<�<Б<t�<:O�<x��<XȊ<��<R<�<�t�<��<��<R�<ך|<	y<Wlu<�q<M;n<o�j<�	g<�pc<��_<A\<[�X<�U<}�Q<��M<�\J<��F<�@C<D�?<e.<<M�8<8'5<u�1<-.<S�*<rA'<��#<7f <=�<�<p?<�<�<~F<��<c�<W�<ߔ�;�5�;���;5��;Ih�;?�;C$�;��;B�;�+�;�K�;�{�;��;�	�;�h�;@פ;�U�;f�;��;�1�;���;���;#>;Ou;�k;�8a;vW;��M;=ND;0�:;o�1;�v(;3j;�z;�;b�;���:M��:���:hB�:R۵:���:6��:�Ʌ:�Al:CHM:ڤ.:�S:��9�H�9�]9a5�8��*�����/n��#�����h��EM*�=oE�'^`�.{��Ҋ�������,������˺سغ�l应򺿮��������|�@D�Bp��$���*���0���6��=��C��#I��/O�|8U�b?[�:Da��Gg�>Jm�~Ks�FLy�yL���������J���^������^�������򳗻_����  �  �h=�=��= E=l�=q�=8=�� =�Y =��<�%�<�]�<,��<���<� �<�5�<�h�<i��<���<���<�+�<|Y�<��<ݰ�<���<��<)�<N�<@q�<ڒ�<��<m��<Y��<G�<.�<�3�<}G�<�X�<�g�<-t�<B~�<���<���<���<���<���<��<�x�<0l�<�\�<�I�<�3�<0�<N��<��<0��<ɑ�<�f�<8�<��<k��<x��<�W�<��<S��<���<T9�<���<}��<(9�<���<�z�<l�<i��<^?�<�λ<�Y�<e�<,e�<B�<�a�<|ڲ<�O�<���<%0�<>��<%�<�g�<|ɧ<0(�<ك�<�ܢ<�2�<|��<�ם<&�<_r�<P��<>�<J�<���<Б<g�<>O�<t��<eȊ<��<Y<�<�t�<���<��<I�<�|<y<Tlu<�q<M;n<r�j<d	g<�pc<��_<A\<\�X<�U<��Q<��M<�\J<��F<�@C<T�?<_.<<f�8</'5<}�1<�,.<Z�*<�A'<��#<Mf <&�<��<m?</�<�<iF<��<^�<n�<˔�; 6�;���;��;.h�;?�;y$�;��;Z�;�+�;�K�;�{�;׺�;�	�;h�;Tפ;�U�;q�;��;�1�;���;Ŀ�;v>;iu;�k;�8a;�uW;��M;�MD;��:;��1;�v(;-j;�z;ѧ;m�;_��:���:���:\B�:�۵:���:M��:lʅ:K@l:^GM:�.:T:���98H�9]9�4�8 �*�T���2n��#����湨��
N*��mE��^`��{�aӊ�������\�����;�˺��غ$m���ۭ�����w�����C�0p�ؖ$�}�*�"�0���6�=�!C��#I�h/O�Q8U��?[�UDa�"Hg��Im��Ks�QLy�KL�������������^������K�����������,����  �  �h=�=��=E=i�=p�=3=�� =�Y =��<�%�<�]�<%��<���<� �<{5�<�h�<_��<���<���<�+�<�Y�<��<ݰ�<s��<��<)�<N�<Dq�<ɒ�<���<a��<V��<N�<,�<�3�<~G�<�X�<�g�<6t�<<~�<���<���<���<��<���<��<�x�<*l�<�\�<�I�<�3�<&�<L��<���<0��<ʑ�<�f�<8�<��<u��<t��<�W�<��<H��<���<H9�<���<~��<)9�<���<�z�<w�<^��<e?�<�λ<�Y�<e�<1e�<B�<�a�<�ڲ<�O�<���<$0�<D��<+�<�g�<}ɧ<%(�<ރ�<�ܢ<�2�<���<�ם<&�<Wr�<T��<9�<J�<���<Б<r�<7O�<x��<ZȊ<��<U<�<�t�<��<��<P�<ٚ|<y<Tlu<�q<W;n<q�j<�	g<�pc<��_<A\<P�X<�U<|�Q<��M<�\J<��F<�@C<H�?<Z.<<R�8<<'5<k�1<-.<]�*<xA'<��#<?f <*�<�<l?<�<�<vF<��<i�<Z�<˔�;�5�;���;!��;,h�;?�;3$�;��;(�;�+�;L�;�{�;��;�	�;�h�;*פ;�U�;X�;��;�1�;���;���;>;ju;�k;�8a;�uW;��M;8ND;6�:;r�1;�v(;0j;�z;��;b�;���:T��:{��:�A�:�۵:⥥:h��:�Ʌ:�Al:nGM:�.:�S:���9K�97]9D;�8i�*�:���`n�V"��ÿ�&��{L*��oE��^`�{�ӊ�x�����G��}����˺:�غ�l�<򺥮����������"D�|p���$���*���0���6��=�zC�$I��/O��8U�Z?[�qDa��Gg�7Jm�Ks�QLy��L�q�������U���_�������l�������೗�a����  �  �h=�=��=E=k�=v�=/=�� =�Y =��<�%�<�]�<+��<���<�<v5�<�h�<_��<���<���<�+�<�Y�<څ�<��<q��<��<)�<N�<Nq�<���<���<c��<W��<E�<'�<�3�<pG�<�X�<�g�<<t�<9~�<���<���<���<��<z��<��<�x�<+l�<�\�<�I�<�3�< �<T��<���<3��<Б�<�f�<8�<��<v��<o��<�W�<��<B��<̆�<A9�<���<y��<.9�<���<�z�<��<Y��<f?�<�λ<�Y�<d�<'e�<B�<�a�<�ڲ<�O�<���<%0�<E��<,�<�g�<�ɧ<(�<胤<�ܢ<�2�<���<�ם<&�<Qr�<a��<6�<
J�<���<Б<t�<0O�<���<VȊ<��<^<�<�t�<��<��<Z�<̚|<y<clu<�q<P;n<U�j<�	g<�pc<��_<A\<`�X<�U<k�Q<��M<�\J<��F<�@C<P�?<r.<<B�8<S'5<b�1<-.<E�*<{A'<��#<6f <L�<ߜ<{?<�<�<qF<��<~�<D�<��;�5�;���;-��;#h�;=?�;$�;�;1�;�+�;�K�;�{�;��;�	�;�h�;פ;�U�;P�;��;�1�;���;��;�=;�u;�k;�8a;3vW;u�M;OND;�:;��1;�v(;Ij;�z;d�;��;?��:X��:-��:uB�:�۵:���:��:2Ʌ:�Bl:�FM:��.:9T:b��9jM�9�]9,<�8�>+�v����n��$�����M��K*�qE�M]`��{��Ҋ�n�����Z����U�˺*�غ;m庚�̮��[�����7�9D�Yp���$��*���0���6��=��C��#I�B/O��8U�#?[��Da��Gg�jJm�XKs�Ly��L����礪�6����������p�������ɳ�������  �  �h=�=��=E=m�=s�=1=�� =�Y =��<�%�<�]�<.��<���<� �<x5�<�h�<h��<���<���<�+�<�Y�<݅�<��<z��<��<)�<N�<Hq�<̒�<���<g��<]��<K�<-�<�3�<{G�<�X�<�g�<3t�<=~�<���<���<���<��<���<��<�x�<*l�<�\�<�I�<�3�<*�<S��<��<,��<Ƒ�<�f�<8�<��<q��<r��<�W�<��<F��<Æ�<L9�<���<~��</9�<���<�z�<v�<a��<i?�<�λ<�Y�<e�<-e�<G�<�a�<�ڲ<�O�<���<%0�<G��<*�<�g�<�ɧ<(�<ރ�<�ܢ<�2�<~��<�ם<&�<Vr�<O��</�<J�<���<Б<t�<4O�<y��<ZȊ<��<^<�<�t�<��<��<W�<ښ|<y<Wlu<�q<`;n<i�j<t	g<�pc<��_<A\<\�X<�U<�Q<��M<�\J<��F<�@C<V�?<g.<<H�8<;'5<i�1<-.<S�*<�A'<��#<+f <(�<�<s?<+�<�<{F<��<g�<J�<���;�5�;���;3��;h�;#?�;B$�;��;C�;�+�;�K�;�{�;�;�	�;�h�;<פ;�U�;^�;��;�1�;���;�;&>;�u;�k;�8a;�uW;��M;ND;W�:;��1;�v(;j;|z;��;��;���:��:c��:,B�:�۵:ƥ�:���:�Ʌ:�Al:}GM:��.:�T:��9�J�9�]93?�8#�*������n�]#��|�湟���L*��oE��]`��{��Ҋ����"����������˺,�غ�l庵������������rD�&p���$���*���0���6��=�vC��#I�B/O��8U�a?[��Da��Gg�4Jm��Ks�DLy�lL�_���Ǧ��z���g�������Y�����������[����  �  �h=�=��=E=i�=s�=7=�� =�Y =��<�%�<�]�<+��<���<� �<�5�<�h�<c��<���<���<�+�<Y�<��<ݰ�<r��<��<)�<	N�<:q�<Ғ�<���<k��<Q��<J�<2�<�3�<�G�<�X�<�g�<3t�<C~�<���<���<���<���<���<��<�x�<,l�<~\�<�I�<�3�<+�<E��<��<2��<ʑ�<�f�<8�<��<p��<x��<�W�<��<P��<���<N9�<���<���<*9�<���<�z�<u�<f��<Y?�<�λ<�Y�<i�</e�<9�<�a�<�ڲ<�O�<���<(0�<I��< �<�g�<{ɧ</(�<܃�<�ܢ<�2�<���<�ם<&�<br�<Q��<<�<J�<�<Б<m�<;O�<p��<aȊ<��<S<�<�t�<��<��<J�<ښ|<y<^lu<�q<H;n<��j<u	g<�pc<��_<A\<c�X<�U<��Q<��M<�\J<��F<�@C<E�?<f.<<a�8<-'5<q�1<-.<[�*<tA'<��#<If <(�<��<e?<!�<�<~F<�<b�<k�<̔�;�5�;���;,��;?h�;�>�;X$�;��;P�;n+�;�K�;�{�;뺵;
�;jh�;Cפ;�U�;v�;���;�1�;�;ο�;.>;/u;�k;�8a;�uW;��M;ND;^�:;9�1;�v(;>j;�z;ǧ;�; ��:���:���:�A�:�۵:b��:ݟ�:ʅ:@l:�HM:+�.:WS:���9oJ�9,	]9u/�8L�*�����:n��"�����)��M*��nE�W_`��{��Ҋ�-��k��r������˺r�غ�l府�S���ל�^����	D�@p��$���*���0���6�8=�>C��#I��/O��8U��?[�Da�Hg�4Jm�\Ks�'Ly��L���������y���<������l�������賗�T����  �  �h=�=��=!E=k�=t�=0=�� =�Y =��<�%�<�]�</��<���<� �<w5�<�h�<e��<���<���<�+�<�Y�<߅�<��<v��<��<)�<N�<Dq�<ʒ�<���<h��<]��<N�<'�<�3�<{G�<�X�<�g�<3t�<>~�<���<���<���<��<���<��<�x�<+l�<�\�<�I�<�3�<'�<S��< ��<.��<Ǒ�<�f�<8�<��<r��<t��<�W�<��<I��<Ć�<M9�<���<{��<+9�<���<�z�<u�<f��<e?�<�λ<�Y�<a�<1e�<G�<�a�<�ڲ<�O�<���<&0�<C��<-�<�g�<�ɧ<"(�<䃤<�ܢ<�2�<~��<�ם<&�<Ur�<R��<7�<J�<���<Б<m�<6O�<}��<WȊ<��<Y<�<�t�<��<��<M�<ۚ|<y<Wlu<�q<T;n<h�j<u	g<�pc<��_<A\<[�X<�U<|�Q<��M<�\J<��F<�@C<N�?<l.<<E�8<G'5<l�1<-.<T�*<�A'<��#<8f <)�<�<�?<'�<�<pF<��<{�<N�<��;�5�;���;"��;*h�;?�;:$�;��;F�;�+�;L�;�{�;ẵ;�	�;�h�;Mפ;�U�;b�;��;�1�;���;���;A>;�u;�k;�8a;'vW;��M;ND;>�:;��1;�v(;j;�z;��;��;���:��:���:�B�:�۵:���:���:�Ʌ:nAl:GM:2�.:&T:��9�J�9�	]9�;�8a�*�#���%n�_"��V��J��|L*��oE�-^`��{�ӊ�\��]����������˺�غm庸�V���N�������8D�3p�Ö$���*���0���6��=��C��#I�b/O�i8U�D?[��Da��Gg�/Jm�bKs�CLy�VL�x���Ȧ��x���{������J�������ڳ��a����  �  �h=�=��=E=g�=u�=0=�� =�Y =��<�%�<�]�<*��<���<�<m5�<�h�<\��<���<���<�+�<�Y�<م�<��<n��<��<)�< N�<Nq�<ǒ�<���<^��<Z��<G�<-�<�3�<vG�<�X�<�g�<6t�<9~�<���<���<���<��<y��<��<�x�<*l�<�\�<�I�<�3�<!�<O��<���<0��<͑�<�f�<8�<��<~��<k��<�W�<��<E��<̆�<@9�<���<x��</9�<���<�z�<x�<Z��<j?�<�λ<�Y�<h�<*e�<F�<�a�<�ڲ<�O�<���<%0�<A��<0�<�g�<�ɧ<(�<僤<�ܢ<�2�<���<~ם<&�<Kr�<_��</�<	J�<���<Б<}�<(O�<���<WȊ<��<U<�<�t�<��<��<Y�<ך|<	y<Ulu<�q<Y;n<g�j<�	g<�pc<��_<A\<P�X<�U<x�Q<��M<�\J<��F<�@C<?�?<o.<<D�8<U'5<U�1<-.<S�*<wA'<��#<&f <I�<͜<q?<�<�<{F<w�<~�<B�<��;�5�;���;&��;h�;;?�;-$�;��;�;�+�;�K�;�{�;#��;�	�;�h�;פ;�U�;N�;��;2�;���;��;�=;�u;�k;�8a;%vW;F�M;�ND;�:;��1;jv(;+j;�z;C�;��;.��:ب�:���:OB�:�۵:���:��:,Ʌ:�Bl:�FM:��.:�T:4��9\K�9a]9�?�8d+������n�6$����湕���K*�(pE�]`�{�*ӊ�(�����G������˺[�غ	m�1�����|����J�uD�ap��$���*�u�0�3�6��=��C��#I��/O��8U�?[��Da��Gg�?Jm�}Ks�NLy��L�n���ʦ��2���k������f�������۳��j����  �  �h=�=��=E=k�=s�=3=�� =�Y =��<�%�<�]�<0��<���<� �<|5�<�h�<`��<���<���<�+�<�Y�<��<��<u��<��<)�<N�<Bq�<Β�<���<i��<V��<C�<0�<�3�<{G�<�X�<�g�<9t�<>~�<���<���<���<��<��<��<�x�<(l�<�\�<�I�<�3�<#�<N��<��</��<ˑ�<�f�<8�<��<r��<p��<�W�<��<G��<ǆ�<H9�<���<��<+9�<���<�z�<z�<`��<a?�<�λ<�Y�<g�<*e�<@�<�a�<�ڲ<�O�<���<%0�<B��<%�<�g�<�ɧ<#(�<���<�ܢ<�2�<���<�ם<&�<Zr�<Y��<5�<J�<���<	Б<t�<2O�<z��<\Ȋ<��<Y<�<�t�<��<��<O�<ښ|<y<jlu<�q<K;n<q�j<u	g<�pc<��_<
A\<h�X<�U<~�Q<��M<�\J<��F<�@C<L�?<g.<<S�8<?'5<g�1<-.<D�*<vA'<��#<9f <;�<�<u?<�<�<sF<��<m�<T�<��;�5�;���;��;%h�;?�;H$�;��;I�;�+�;�K�;�{�;���;�	�;�h�;-פ;�U�;`�;	��;�1�;���;ῄ;>;�u;�k;�8a;�uW;��M;!ND;�:;��1;�v(;%j;�z;��;y�;y��:&��:A��:�A�:s۵:֥�:ʠ�:�Ʌ:Al:�GM:L�.:�S:R��9�K�9]9i7�8��*�q���Vn�$��N�湢��,L*�YoE��^`��{�*ӊ����o����������˺S�غm庇򺦮��������|�ED�!p���$��*���0���6��=�hC��#I�i/O��8U��?[�^Da��Gg�6Jm�rKs��Ky��L���������y���X���&���i�������޳��^����  �  �h=�=��="E=k�=m�=4=�� =�Y =��<�%�<�]�<(��<���<� �<}5�<�h�<j��<���<���<�+�<}Y�<��<ذ�<��<��<)�<N�<@q�<Ԓ�<~��<l��<Y��<M�<3�<�3�<�G�<�X�<�g�</t�<=~�<���<���<���<���<���<��<�x�<(l�<�\�<�I�<�3�</�<M��<��<.��<Ƒ�<�f�<8�<��<f��<~��<�W�<��<F��<���<U9�<���<���<,9�<���<�z�<p�<m��<c?�<�λ<�Y�<g�<3e�<C�<�a�<ڲ<�O�<���<.0�<L��<&�<�g�<xɧ<&(�<ۃ�<�ܢ<�2�<z��<�ם<&�<Yr�<L��<7�<	J�<���<Б<i�<DO�<t��<\Ȋ<��<W<�<�t�<��<��<H�<�|<�y<^lu<�q<N;n<��j<s	g<�pc<��_<A\<a�X<�U<��Q<��M<�\J<��F<�@C<N�?<O.<<V�8<0'5<��1<-.<W�*<�A'<��#<:f <�<�<k?</�<�<qF<��<_�<[�<���;�5�;���;2��;Ph�;?�;`$�;��;V�;�+�;L�;�{�;躵;
�;�h�;aפ;�U�;]�;+��;�1�;�;ֿ�;x>;Uu;|k;�8a;�uW;��M;�MD;~�:;v�1;�v(;j;z;��;K�;5��:f��:��:B�:l۵:���:��:oʅ:�@l:�HM:S�.:�T:��97I�9�]9L9�8U�*�]���=n��!����湢���M*��nE�l^`��{�~Ҋ����������r���˺޳غ�l��� �����������4D�^p�ؖ$�|�*��0�[�6�=�fC�-$I�x/O�<8U��?[�Da�%Hg��Im��Ks�)Ly�QL���������}���9������Q����������:����  �  �h=�=��=E=j�=t�=7=�� =�Y =��<�%�<�]�<*��<���< �<{5�<�h�<d��<���<���<�+�<�Y�<��<��<w��<��<)�<N�<Eq�<В�<���<d��<S��<I�<,�<�3�<xG�<�X�<�g�<5t�<A~�<���<���<���< ��<���<��<�x�<0l�<�\�<�I�<�3�<)�<K��< ��<5��<ϑ�<�f�<8�<��<k��<w��<�W�<��<N��<ņ�<H9�<���<��<'9�<���<�z�<x�<^��<b?�<�λ<�Y�<f�<,e�<?�<�a�<�ڲ<�O�<���<#0�<F��<#�<�g�<�ɧ<*(�<⃤<�ܢ<�2�<{��<�ם<&�<Wr�<\��<:�<J�<���<Б<l�<6O�<{��<cȊ<��<W<�<�t�<	��<��<K�<�|<y<_lu<	�q<P;n<j�j<�	g<�pc<��_<A\<]�X<�U<��Q<��M<�\J<��F<�@C<K�?<j.<<a�8<A'5<j�1<-.<R�*<}A'<��#<<f <?�<�<j?<#�<�<vF<�<p�<c�<��;�5�;���;-��;h�;?�;Q$�;��;4�;u+�;�K�;�{�;��;�	�;�h�;%פ;�U�;m�;!��;�1�;���;޿�;>;�u;�k;�8a;�uW;��M;�MD;N�:;f�1;�v(;Vj;�z;��;K�;��:���:���:B�:�۵:A��:���:�Ʌ:�@l:�GM:��.:�T:��9FK�9+]9e8�8��*������n��#��k�����L*�6oE��]`�>{��Ҋ� ��W�����.����˺H�غ�l���X���������c�D�Np���$���*���0���6��=�2C��#I�z/O��8U�q?[�mDa�Hg�Jm�YKs�%Ly��L����Ŧ��M���e������s�������ݳ��G����  �  ;h==��=(D=V�=6�=�=6� =.X =���<4"�<�Y�<��<���<��<U0�<�c�<���<���<���<&%�<�R�<�~�<)��<m��<%��<W �<�D�<�g�<��<A��<���<H��<���<C�<�'�<�:�<�K�<Z�<4f�<�o�<�v�<<{�<�|�<�{�<�w�<q�<@g�<dZ�<hJ�<(7�<� �<��<���<��<��</}�<�Q�<�"�<@��<��<��<�A�<���<��<rp�<�"�<|��<|�<�"�<���<]d�<Q��<P��<�)�<ḻ<wD�<8̸<IP�<�е<fM�<�Ʋ<J<�<���<m�<��<_�<�V�<���<��<!t�<�͢<P$�<tx�<�ɝ<+�<�e�<���<��<�?�<��<�Ƒ<��<@G�<5��<���<���<�6�<�o�<�<߁<{�<��|<y<�ju<��q<L<n<��j<)g<�uc<��_<xH\<�X<�U<ɋQ<L�M<�jJ<��F<FQC<�?<UA<<��8<�<5<H�1<3E.<��*< \'<��#<1� <W<?�<
`<�<�<hj<�#	<��<V�<���;͇�;�7�;���;M��;���;h~�;�s�;w�;���;5��;�ۻ;8�;�k�;(˪;�9�;��;H�;��;���;�T�;�#�;c�;C�u;%�k;�a;I8X;�N;�E;e�;;�Z2;`.); ;�,;"W;��;X��:���:�!�:F��:U�: צ:�ʖ:&�:-zn:�qO:��0:�_:��9�)�9��d9|��8�]h�q��yg�A�æ��u���(�0D��_��y�/4��=i��������\����h˺�8غ���L��C��ai�Q��������F��o$��*��0�;�6��<�}�B�&
I�,O�R"U�.+[�:2a��7g��;m� ?s��Ay��C�䢂�]���z���ܧ��(�������ű��ᶗ�Q����  �  Bh==��='D=T�=?�=�=(� =+X =���<-"�<�Y�<��<��<)��<]0�<�c�<���<���<z��<%�<rR�<�~�<2��<m��<!��<K �<�D�<�g�<��<>��<���<=��<���<D�<�'�<�:�<�K�< Z�<8f�<�o�<�v�<H{�<�|�<�{�<�w�<q�<Og�<`Z�<PJ�<7�<� �<��<���<��<��<7}�<�Q�<�"�<G��<չ�<��<�A�<���<��<qp�<�"�<q��<|�<�"�<���<cd�<R��<_��<�)�<⸻<pD�<6̸<FP�<�е<rM�<�Ʋ<X<�<���<u�< ��<Y�<�V�<���<��<t�<�͢<A$�<`x�<�ɝ<(�<f�<���<��<�?�<��<�Ƒ<��<7G�<��<���<���<�6�<�o�<姃<߁<��<��|< y<�ju<��q<8<n<��j<g<�uc<��_<sH\<�X<�U<��Q<h�M<�jJ<��F<AQC<�?<zA<<��8<�<5<<�1<E.<��*<
\'<z�#<@� <m<O�<�_<�<ζ<Lj<u#	<U�<q�<���;̇�;�7�;���;c��;���;�~�;�s�;>w�;���;!��;�ۻ;�;�k�;˪;5:�;-��;
H�;�;ە�;�T�;g#�;\�;�u;��k;��a;�7X;��N;HE;��;;�Z2;t.);] ;-;YW;�;���:`��:!�:��:��:
ئ:�ʖ:>�:�xn:wqO:�0:�a:���9*�9��d9���8:h��#�{g����[t���(�D�|_��y��4���i��򇤺����p����i˺L9غ��亗��nC��si���a��l��F��o$��*���0���6���<�5�B��	I�kO�~"U��+[�2a�o7g�{;m�?s�wAy��C�
���N�������ǧ��I�����������𶗻#����  �  :h==��=-D=R�==�=�=(� =4X =���<6"�<�Y�<ݐ�<���<#��<W0�<zc�<���<���<���<0%�<sR�<�~�<)��<k��<)��<M �<�D�<�g�<��<2��<���<=��<���<G�<�'�<�:�<�K�<"Z�</f�<�o�<�v�<:{�<�|�<�{�<�w�<q�<Ng�<cZ�<^J�<37�<� �<��<���<��<��<1}�<�Q�<�"�<O��<ٹ�<��<�A�<���<��<jp�<�"�<r��<|�<�"�<}��<Wd�<G��<b��<�)�<<jD�<7̸<RP�<�е<vM�<�Ʋ<L<�<���<n�<��<]�<�V�<���<��<t�<�͢<Q$�<gx�<ʝ<�<�e�<���<��<�?�<��<�Ƒ<��<KG�<��<���<���<�6�<�o�<꧃<߁<x�<��|<� y<�ju<��q<=<n<��j<�g<�uc<��_<sH\<�X<�U<ɋQ<I�M<�jJ<��F<YQC<�?<qA<<��8<�<5<b�1<E.<��*<\'<g�#<6� <a<B�<�_<�<޶<fj<�#	<W�<p�<���;Ƈ�;�7�;���;X��;���;k~�;Vs�;Ew�;���;J��;�ۻ;��;�k�;�ʪ;;:�;��;�G�;��;���;�T�;s#�;~�;��u;��k;�a;�7X;P�N;lE;Ԥ;;TZ2;$.);. ;�,;W;��;A��:���:R"�:
��:��:�צ:rʖ:��:
yn:�qO:T�0:x_:���9;'�9̋d9���87�f�*츠zg���B���s�`�(��D�	_���y��4��bi��􇤺U���|����i˺"8غ���$���B���i�@�������?G��o$���*�_�0���6���<�?�B��	I��O�""U�m+[�2a��7g��;m�a?s��Ay��C� ��������������9��������������R����  �  >h==��=(D=U�=>�=�=2� =%X =���<0"�<�Y�<��<���<$��<X0�<�c�<���<���<{��<%�<�R�<�~�<4��<j��<%��<Q �<�D�<�g�<��<F��<���<E��<���<@�<�'�<�:�<�K�<Z�<5f�<�o�<�v�<A{�<�|�<�{�<�w�<!q�<Gg�<bZ�<`J�<7�<� �<��<���<��<��<4}�<�Q�<�"�<B��<ݹ�<��<�A�<���<��<vp�<�"�<v��<|�<�"�<���<nd�<R��<U��<�)�<⸻<oD�<4̸<FP�<�е<jM�<�Ʋ<[<�<���<s�<��<]�<�V�<���<��<t�<�͢<B$�<jx�<�ɝ<0�<f�<���<��<�?�<��<�Ƒ<��<.G�<*��<���<���<�6�<�o�<<߁<�<��|< y<�ju<��q<;<n<��j<g<�uc<��_<xH\<�X<�U<܋Q<V�M<�jJ<��F<FQC<�?<uA<<��8<�<5<#�1<E.<��*<\'<��#<6� <d<E�<`<�<�<Oj<d#	<}�<\�<���;�;�7�;���;`��;՗�;�~�;�s�;w�;���;'��;�ۻ;�;�k�; ˪;:�;!��;;H�;��;���;�T�;�#�;T�;V�u;]�k;�a;	8X;��N;~E;o�;;�Z2;�.);@ ; -;?W;+�;t��:���:� �:���:7�:�צ:5˖:��:myn:EqO:e�0:�`:Y��9%*�9��d9	��8�Fh��$�!|g���E��Hu�s�(�D��_�Q�y�q4��Xi��4�����������h˺y9غ������C��5i�,��������F��o$���*�M�0���6�i�<�x�B��	I�;O�g"U�L+[�B2a��7g��;m��>s��Ay��C����L���ǥ��ͧ��F�������ñ������-����  �  Ch==��=&D=S�=@�=�=5� ='X =���<,"�<�Y�<��<���</��<N0�<�c�<���<���<���<%�<�R�<|~�<:��<b��<&��<Q �<�D�<�g�<܈�<;��<���<N��<���<G�<�'�<�:�<�K�<Z�<0f�<�o�<�v�<G{�<�|�<�{�<�w�<!q�<Cg�<bZ�<eJ�<!7�<� �<��<���<��<��<9}�<�Q�<�"�<9��<��<��<�A�<���<��<wp�<�"�<���<|�<�"�<���<Xd�<L��<[��<�)�<ܸ�<yD�<;̸<AP�<�е<iM�<�Ʋ<G<�<���<r�<��<b�<�V�<���<��<&t�<�͢<O$�<kx�<�ɝ<3�<�e�<���<��<�?�<��<�Ƒ<��<4G�<2��<���<���<�6�<�o�<���<߁<��<y�|<y<�ju<��q<F<n<��j< g<�uc<��_<�H\<�X<�U<��Q<j�M<�jJ<��F<=QC<	�?<zA<<��8<�<5<.�1<BE.<��*<\'<��#<#� <y<1�<`<�<ݶ<pj<t#	<��<E�<��;���;�7�;���;R��;��;U~�;ys�;w�;ԉ�;��;�ۻ;6�;�k�;0˪;1:�;��;�G�;��;ו�;�T�;�#�;3�;Z�u;:�k;�a;88X;��N;�E;�;;�Z2;9.);J ;/-;�V;S�;���:���:�!�:���:^�:"צ:K˖:r�:�zn:�pO:��0:-`:��9}(�9��d9x��8 i�\�wxg�8򫹢��ru�{�(��D��_�{�y��4��i��Ɉ��6�������Wh˺�8غ���ڤ�D��"i����3�����F��o$��*���0���6�(�<���B��	I�\O��"U�+[�i2a�c7g�<m�?s��Ay��C��X�������ǧ��8���k���ձ��򶗻t����  �  @h==��=+D=R�=<�=�=,� =.X =���<,"�<Z�<��<���<.��<R0�<�c�<���<���<��<$%�<zR�<�~�<4��<i��<*��<J �<�D�<�g�<��<A��<���<8��<���<I�<�'�<�:�<�K�<Z�<5f�<�o�<�v�<D{�<�|�<�{�<�w�<q�<Dg�<^Z�<YJ�<$7�<� �<��<���<��<��<8}�<�Q�<�"�<K��<չ�<��<�A�<���<��<rp�<�"�<w��<|�<�"�<���<dd�<P��<\��<�)�<鸻<iD�<8̸<GP�<�е<pM�<�Ʋ<U<�<���<p�<���<a�<�V�<���<��<t�<�͢<G$�<`x�<ʝ<(�<�e�<���<��<�?�<"��<�Ƒ<��<?G�< ��<���<���<�6�<�o�<맃<߁<��<��|<y<�ju<��q<0<n<��j<�g<�uc<��_<jH\< �X<�U<ϋQ<_�M<�jJ<��F<RQC<�?<nA<<��8<�<5<J�1<E.<��*<#\'<s�#<2� <w<9�<�_<�<ζ<Xj<�#	<e�<V�<���;���;�7�;���;N��;ؗ�;�~�;�s�;?w�;}��;#��;�ۻ;��;�k�;�ʪ;':�; ��;H�;��;̕�;�T�;#�;e�;2�u;I�k;��a;�7X;גN;IE;��;;�Z2;.);X ;"-;�V;2�;��:]��:s!�:{��:��:`צ:�ʖ:A�:�yn:�pO:Q�0:�`:��9~)�9�d9O��8�`g��*��yg�����xt���(��D��_���y��4��i��/�������M���`i˺�8غa�云��B��ui�{��F���� G��o$���*�w�0�H�6���<�[�B��	I�uO�H"U�d+[�X2a��7g��;m��>s�nAy��C���������������S�����������׶��F����  �  :h==��=)D=U�=9�=�=*� =1X =���<2"�<�Y�<��<��<��<g0�<yc�<���<���<~��<'%�<yR�<�~�<+��<q��<%��<M �<�D�<�g�<��<2��<���<:��<���<M�<�'�<�:�<�K�<#Z�<)f�<�o�<�v�<>{�<�|�<�{�<�w�<q�<Ig�<fZ�<ZJ�<-7�<� �<��<���<��<��</}�<�Q�<�"�<O��<ҹ�<��<�A�<���<��<mp�<�"�<o��<|�<�"�<���<cd�<D��<c��<~)�<�<hD�<:̸<JP�<�е<uM�<�Ʋ<Z<�<���<v�<��<[�<�V�<���<��<t�<�͢<J$�<^x�<ʝ<�<f�<���< ��<�?�<��<�Ƒ<��<GG�<��<���<���<�6�<�o�<秃<"߁<y�<��|<� y<�ju<��q<"<n<��j<�g<�uc<��_<tH\<�X<�U<�Q<I�M<�jJ<��F<KQC<�?<`A<<��8<�<5<W�1<E.<��*<\'<p�#<L� <M<c�<�_<�<Ѷ<Vj<�#	<d�<s�<���;އ�;�7�;���;t��;���;�~�;Us�;;w�;���;'��;ܻ;��;�k�;�ʪ;B:�;�;H�;��;���;�T�;e#�;��;#�u;l�k;%�a;�7X;�N;/E;ͤ;;UZ2;�.);H ;�,;vW;��;B��:6��:�!�:���:�:�צ:�ʖ:��:�xn:rO:��0:�`:���9�&�9��d9���8/�f��+��xg��﫹ª��s�t�(�3D�=_���y�y4���i������$�������\i˺�8غ:�享���B���i�������D��F�p$���*���0��6���<���B��	I�QO�A"U��+[��1a��7g��;m�,?s��Ay��C�8��������������m��������������"����  �  <h==��=&D=W�=:�=�=/� =-X =���<7"�<�Y�<��<��<��<`0�<�c�<���<���<���<"%�<�R�<�~�</��<n��<!��<N �<�D�<�g�<��<6��<���<L��<���<E�<�'�<�:�<�K�<'Z�<,f�<�o�<�v�<={�<�|�<�{�<�w�<!q�<Cg�<bZ�<^J�<*7�<� �<��<���<��<��<0}�<�Q�<�"�<H��<޹�<��<�A�<���<��<tp�<�"�<v��<|�<�"�<���<\d�<F��<b��<�)�<۸�<rD�<9̸<@P�<�е<oM�<�Ʋ<P<�<���<m�<��<[�<�V�<���<��<t�<�͢<P$�<ix�<�ɝ<!�<f�<���<��<�?�<��<�Ƒ<��<?G�<%��<���<���<�6�<�o�<�<߁<{�<��|<y<�ju<��q<6<n<��j<g<�uc<��_<�H\<�X<�U<ՋQ<N�M<�jJ<��F<?QC<�?<dA<<��8<�<5<E�1<*E.<��*<�['<z�#<C� <N<U�<�_<�<�<hj<~#	<w�<X�<���;҇�;�7�;���;G��;ʗ�;�~�;fs�;#w�;Ή�;
��;�ۻ;�;�k�;˪;N:�;���;�G�;��;���;�T�;�#�;[�;V�u;<�k;�a;�7X;�N;�E;��;;TZ2;b.);A ;�,;KW;ǜ;���:���:�!�:ց�:!�:Yצ:˖:5�:�yn:�pO:��0:N`:��96'�9��d9x��8�%i��!츻yg���]�㹶t��(�jD�7_��y��4���i������͑��I����h˺�8غ������TC���i�������g��F�$p$���*� �0�E�6���<�N�B��	I�*O�z"U�5+[�b2a��7g��;m�?s��Ay�jC����T�������ɧ��Y���Y���ͱ������8����  �  Eh==��=&D=S�=>�=�=2� ='X =���<("�< Z�<��<���<4��<Q0�<�c�<���<���<~��<%�<�R�<�~�<8��<b��<%��<Q �<�D�<�g�<ވ�<N��<���<B��<���<@�<�'�<�:�<�K�<Z�<9f�<�o�<�v�<L{�<�|�<�{�<�w�<$q�<Eg�<dZ�<]J�<7�<� �<��<���<��<��<=}�<�Q�<�"�<E��<ڹ�<��<�A�<���<��<|p�<�"�<|��<|�<�"�<���<_d�<X��<N��<�)�<ݸ�<uD�<6̸<DP�<�е<aM�<�Ʋ<K<�<���<n�<��<`�<�V�<���<��<!t�<�͢<F$�<cx�<ʝ<2�<�e�<���<��<�?�<#��<�Ƒ<��<2G�<)��<���<���<�6�<�o�<���<
߁<��<�|<y<�ju<��q<L<n<��j<g<�uc<��_<fH\<�X<�U<��Q<u�M<�jJ<��F<=QC<�?<sA<<��8<�<5<-�1<E.<��*<\'<��#<4� <�<6�<`<�<Ѷ<Vj<m#	<��<T�<	��;���;�7�;���;5��;��;^~�;�s�;w�;���;&��;�ۻ;&�;�k�;-˪;�9�;3��;H�;��;앏;vT�;�#�;1�;p�u;Q�k;�a;�7X;��N;kE;j�;;�Z2;.);r ;H-;�V;o�;���:���:"!�:���:B�:cצ:�˖:l�:0zn:0pO:�0:a:���9�+�9�d9���8��h���!{g�g�ڧ�^v�W�(�D��_��y��4��-i���������V����h˺X9غv��\��C��&i�r�������F��o$��*�R�0���6�q�<�L�B��	I�]O��"U�+[��2a�;7g�<m��>s��Ay�'D�䢂�g�������⧋�.���������������p����  �  Bh==��=(D=U�=<�=�=-� =0X =���<."�<�Y�<��<���<%��<V0�<�c�<���<���<���<(%�<~R�<�~�<1��<j��<)��<S �<�D�<�g�<و�<<��<���<?��<���<E�<�'�<�:�<�K�<Z�<5f�<�o�<�v�<E{�<�|�<�{�<�w�<q�<Gg�<eZ�<]J�<17�<� �<��<���<	��<��<4}�<�Q�<�"�<@��<��<��<�A�<���<��<sp�<�"�<y��<|�<�"�<���<Vd�<O��<W��<�)�<渻<nD�<7̸<NP�<�е<jM�<�Ʋ<E<�<���<o�<��<a�<�V�<���<��<t�<�͢<X$�<hx�<�ɝ<(�<�e�<���<��<�?�<��<�Ƒ<��<EG�<$��<���<���<�6�<�o�<�<߁<��<p�|<� y<�ju<��q<L<n<��j< g<�uc<��_<kH\<�X<�U<��Q<g�M<�jJ<��F<HQC<�?<mA<<��8<�<5<Q�1<;E.<��*<\'<�#<,� <g<A�<�_<�<ٶ<vj<�#	<m�<_�<���;Ň�;�7�;���;>��;��;I~�;s�;w�;���;J��;�ۻ; �;�k�;!˪;:�;!��;�G�;��;Е�;�T�;�#�;V�;<�u;a�k;�a;�7X;?�N;�E;m�;;�Z2;N.);5 ;-;W;
�;V��: ��:z"�:́�:8�:�צ: ˖:��:�yn:%qO:}�0:M`:Y��9>)�9D�d9���80�g�&츁zg�﫹���Su�9�(��D�W_���y�s4��i��/���������� i˺�8غU����C��wi�=��z�����F��o$���*��0��6���<�(�B��	I�QO�j"U�5+[�V2a�w7g�@<m�5?s��Ay��C�䢂�?���˥������$��������������������  �  8h==��=&D=Y�=:�=�=*� =+X =���<6"�<�Y�<��<��<��<b0�<�c�<���<���<v��< %�<vR�<�~�<,��<s��<��<U �<�D�<�g�<���<9��<���<>��<���<D�<�'�<�:�<�K�<#Z�<1f�<�o�<�v�<8{�<�|�<�{�<�w�<q�<Fg�<^Z�<SJ�< 7�<� �<��<���<��<��<1}�<�Q�<�"�<N��<Թ�<��<�A�<���<��<op�<�"�<m��<|�<�"�<���<id�<J��<d��<~)�<฻<kD�<5̸<@P�<�е<vM�<�Ʋ<_<�<���<r�<	��<T�<�V�<���<��<t�<�͢<?$�<ex�<ʝ<$�<
f�<���<��<�?�<��<�Ƒ<��<8G�<��<���<���<�6�<�o�<駃< ߁<t�<��|<y<�ju<��q<"<n<��j<�g<�uc<��_<~H\<�X<�U<�Q<A�M<�jJ<��F<>QC< �?<eA<<��8<�<5<<�1<E.<��*<\'<��#<A� <N<Y�<�_<�<ݶ<Ej<x#	<^�<l�<���;��;n7�;���;S��;���;�~�;ss�;Ew�;���;���;�ۻ;��;�k�;�ʪ;@:�;��;#H�;	�;���;�T�;\#�;n�;(�u;T�k;��a;�7X;��N;6E;Ϥ;;kZ2;�.);; ;�,;xW;ٜ;+��:M��:!�:��:��:�צ:�ʖ:��:`xn:"rO:��0:�a:I��90(�9͌d9$��8sh�)츋{g��򫹕���s���(��
D�_���y�%4���i���������������i˺G9غ���8��C���i������z��F��o$���*���0�{�6���<�$�B��	I�&O�k"U�x+[�2a�8g�Z;m��>s��Ay��C�7���G���ѥ������x���z�������궗�����  �  8h==��=(D=S�=9�=�=2� =0X =���<7"�<�Y�<��<���<)��<U0�<�c�<���<���<��<.%�<�R�<�~�<'��<h��<"��<W �<�D�<�g�<���<4��<���<C��<���<I�<�'�<�:�<�K�<Z�<+f�<�o�<�v�<6{�<�|�<�{�<�w�<q�<Eg�<gZ�<gJ�<+7�<� �<��<���<	��<��<5}�<�Q�<�"�<K��<߹�<��<�A�<���<��<np�<�"�<u��<|�<�"�<{��<Ud�<F��<\��<�)�<븻<rD�<:̸<IP�<�е<mM�<�Ʋ<I<�<���<p�<��<Y�<�V�<���<��<!t�<�͢<J$�<lx�<ʝ<'�<�e�<���<��<�?�<��<�Ƒ<��<DG�<.��<���<���<�6�<�o�<�< ߁<s�<��|<� y<�ju<��q<7<n<��j<	g<�uc<��_<rH\<�X<�U<ǋQ<?�M<�jJ<��F<EQC<	�?<^A<<��8<�<5<S�1<E.<��*<\'<}�#<2� <n<>�<�_<�<�<Xj<�#	<��<i�<���;���;�7�;���;U��;���;g~�;]s�;&w�;���;&��;�ۻ;�;�k�;˪;#:�;���;�G�;��;���;�T�;�#�;j�;�u;Q�k;-�a;I8X;�N;�E;��;;uZ2;H.);: ;	-;W;��;���:	��:�!�:U��:h�:�צ:�ʖ:T�:cyn:/rO::�0:0_:A��9'�9݈d9���8\g�"�yg�𫹐���t��(�JD�l	_���y��3���i��1���-���ʆ���h˺F8غ,��Ԥ�C��~i�A��S�����F��o$���*�E�0��6�N�<��B��	I�vO�X"U�9+[� 2a�8g��;m�D?s��Ay��C����.�����������R�������ű�����T����  �  Fh==��=)D=T�=@�=�=+� =+X =���<."�<�Y�<��<���<8��<Q0�<�c�<���<���<���<%�<zR�<�~�<5��<m��<*��<E �<�D�<�g�<��<H��<���<>��<���<@�<�'�<�:�<�K�<Z�<@f�<�o�<�v�<H{�<�|�<�{�<�w�< q�<Lg�<_Z�<UJ�<7�<� �<��<���<��<��<;}�<�Q�<�"�<;��<߹�<��<�A�<���<��<wp�<�"�<s��<|�<�"�<���<ed�<[��<U��<�)�<⸻<hD�<1̸<IP�<�е<iM�<�Ʋ<S<�<���<p�<���<_�<�V�<���<��<t�<�͢<J$�<fx�<�ɝ<1�<�e�<���<��<�?�<��<�Ƒ<��<8G�<��<���<���<�6�<�o�<姃<߁<��<��|<y<�ju<��q<G<n<��j<�g<�uc<��_<hH\<�X<�U<ӋQ<v�M<�jJ<��F<KQC<�?<{A<<��8<�<5<>�1<(E.<��*<\'<��#<(� <�<7�<`<�<ֶ<]j<v#	<e�<`�<���;χ�;�7�;x��;:��;��;�~�;�s�;w�;���;1��;�ۻ;��;�k�;˪;:�;O��;H�;��;ܕ�;�T�;l#�;X�;S�u;��k;��a;�7X;��N;�E;G�;;�Z2;_.);V ;;-;W;[�;
��:��:g!�:F��:��:�צ:M˖: �: yn:NpO:ο0:�a:N��9�,�9��d9!��8�0h�Q,�J}g�J�&��tu���(�D�R_���y��4��Ai������T������ki˺Q9غ*��,���C��-i�c�� �����F��o$���*��0���6���<�I�B��	I�YO�V"U��+[�h2a�O7g��;m��>s�LAy��C�좂�I���䥈�ç��2�����������ɶ��?����  �  8h==��=(D=S�=9�=�=2� =0X =���<7"�<�Y�<��<���<)��<U0�<�c�<���<���<��<.%�<�R�<�~�<'��<h��<"��<W �<�D�<�g�<���<4��<���<C��<���<I�<�'�<�:�<�K�<Z�<+f�<�o�<�v�<6{�<�|�<�{�<�w�<q�<Eg�<gZ�<gJ�<+7�<� �<��<���<	��<��<5}�<�Q�<�"�<K��<߹�<��<�A�<���<��<np�<�"�<u��<|�<�"�<{��<Ud�<F��<\��<�)�<븻<rD�<:̸<IP�<�е<mM�<�Ʋ<I<�<���<p�<��<Y�<�V�<���<��<!t�<�͢<J$�<lx�<ʝ<'�<�e�<���<��<�?�<��<�Ƒ<��<DG�<.��<���<���<�6�<�o�<�< ߁<s�<��|<� y<�ju<��q<7<n<��j<	g<�uc<��_<rH\<�X<�U<ǋQ<?�M<�jJ<��F<EQC<	�?<^A<<��8<�<5<S�1<E.<��*<\'<}�#<2� <n<>�<�_<�<�<Xj<�#	<��<i�<���;���;�7�;���;U��;���;g~�;]s�;&w�;���;&��;�ۻ;�;�k�;˪;#:�;���;�G�;��;���;�T�;�#�;j�;�u;Q�k;-�a;I8X;�N;�E;��;;uZ2;H.);: ;	-;W;��;���:	��:�!�:U��:h�:�צ:�ʖ:T�:cyn:/rO::�0:0_:A��9'�9݈d9���8\g�"�yg�𫹐���t��(�JD�l	_���y��3���i��1���-���ʆ���h˺F8غ,��Ԥ�C��~i�A��S�����F��o$���*�E�0��6�N�<��B��	I�vO�X"U�9+[� 2a�8g��;m�D?s��Ay��C����.�����������R�������ű�����T����  �  8h==��=&D=Y�=:�=�=*� =+X =���<6"�<�Y�<��<��<��<b0�<�c�<���<���<v��< %�<vR�<�~�<,��<s��<��<U �<�D�<�g�<���<9��<���<>��<���<D�<�'�<�:�<�K�<#Z�<1f�<�o�<�v�<8{�<�|�<�{�<�w�<q�<Fg�<^Z�<SJ�< 7�<� �<��<���<��<��<1}�<�Q�<�"�<N��<Թ�<��<�A�<���<��<op�<�"�<m��<|�<�"�<���<id�<J��<d��<~)�<฻<kD�<5̸<@P�<�е<vM�<�Ʋ<_<�<���<r�<	��<T�<�V�<���<��<t�<�͢<?$�<ex�<ʝ<$�<
f�<���<��<�?�<��<�Ƒ<��<8G�<��<���<���<�6�<�o�<駃< ߁<t�<��|<y<�ju<��q<"<n<��j<�g<�uc<��_<~H\<�X<�U<�Q<A�M<�jJ<��F<>QC< �?<eA<<��8<�<5<<�1<E.<��*<\'<��#<A� <N<Y�<�_<�<ݶ<Ej<x#	<^�<l�<���;��;n7�;���;S��;���;�~�;ss�;Ew�;���;���;�ۻ;��;�k�;�ʪ;@:�;��;#H�;	�;���;�T�;\#�;n�;(�u;T�k;��a;�7X;��N;6E;Ϥ;;kZ2;�.);; ;�,;xW;ٜ;+��:M��:!�:��:��:�צ:�ʖ:��:`xn:"rO:��0:�a:I��90(�9͌d9$��8sh�)츋{g��򫹕���s���(��
D�_���y�%4���i���������������i˺G9غ���8��C���i������z��F��o$���*���0�{�6���<�$�B��	I�&O�k"U�x+[�2a�8g�Z;m��>s��Ay��C�7���G���ѥ������x���z�������궗�����  �  Bh==��=(D=U�=<�=�=-� =0X =���<."�<�Y�<��<���<%��<V0�<�c�<���<���<���<(%�<~R�<�~�<1��<j��<)��<S �<�D�<�g�<و�<<��<���<?��<���<E�<�'�<�:�<�K�<Z�<5f�<�o�<�v�<E{�<�|�<�{�<�w�<q�<Gg�<eZ�<]J�<17�<� �<��<���<	��<��<4}�<�Q�<�"�<@��<��<��<�A�<���<��<sp�<�"�<y��<|�<�"�<���<Vd�<O��<W��<�)�<渻<nD�<7̸<NP�<�е<jM�<�Ʋ<E<�<���<o�<��<a�<�V�<���<��<t�<�͢<X$�<hx�<�ɝ<(�<�e�<���<��<�?�<��<�Ƒ<��<EG�<$��<���<���<�6�<�o�<�<߁<��<p�|<� y<�ju<��q<L<n<��j< g<�uc<��_<kH\<�X<�U<��Q<g�M<�jJ<��F<HQC<�?<mA<<��8<�<5<Q�1<;E.<��*<\'<�#<,� <g<A�<�_<�<ٶ<vj<�#	<m�<_�<���;Ň�;�7�;���;>��;��;I~�;s�;w�;���;J��;�ۻ; �;�k�;!˪;:�;!��;�G�;��;Е�;�T�;�#�;V�;<�u;a�k;�a;�7X;?�N;�E;m�;;�Z2;N.);5 ;-;W;
�;V��: ��:z"�:́�:8�:�צ: ˖:��:�yn:%qO:}�0:M`:Y��9>)�9D�d9���80�g�&츁zg�﫹���Su�9�(��D�W_���y�s4��i��/���������� i˺�8غU����C��wi�=��z�����F��o$���*��0��6���<�(�B��	I�QO�j"U�5+[�V2a�w7g�@<m�5?s��Ay��C�䢂�?���˥������$��������������������  �  Eh==��=&D=S�=>�=�=2� ='X =���<("�< Z�<��<���<4��<Q0�<�c�<���<���<~��<%�<�R�<�~�<8��<b��<%��<Q �<�D�<�g�<ވ�<N��<���<B��<���<@�<�'�<�:�<�K�<Z�<9f�<�o�<�v�<L{�<�|�<�{�<�w�<$q�<Eg�<dZ�<]J�<7�<� �<��<���<��<��<=}�<�Q�<�"�<E��<ڹ�<��<�A�<���<��<|p�<�"�<|��<|�<�"�<���<_d�<X��<N��<�)�<ݸ�<uD�<6̸<DP�<�е<aM�<�Ʋ<K<�<���<n�<��<`�<�V�<���<��<!t�<�͢<F$�<cx�<ʝ<2�<�e�<���<��<�?�<#��<�Ƒ<��<2G�<)��<���<���<�6�<�o�<���<
߁<��<�|<y<�ju<��q<L<n<��j<g<�uc<��_<fH\<�X<�U<��Q<u�M<�jJ<��F<=QC<�?<sA<<��8<�<5<-�1<E.<��*<\'<��#<4� <�<6�<`<�<Ѷ<Vj<m#	<��<T�<	��;���;�7�;���;5��;��;^~�;�s�;w�;���;&��;�ۻ;&�;�k�;-˪;�9�;3��;H�;��;앏;vT�;�#�;1�;p�u;Q�k;�a;�7X;��N;kE;j�;;�Z2;.);r ;H-;�V;o�;���:���:"!�:���:B�:cצ:�˖:l�:0zn:0pO:�0:a:���9�+�9�d9���8��h���!{g�g�ڧ�^v�W�(�D��_��y��4��-i���������V����h˺X9غv��\��C��&i�r�������F��o$��*�R�0���6�q�<�L�B��	I�]O��"U�+[��2a�;7g�<m��>s��Ay�'D�䢂�g�������⧋�.���������������p����  �  <h==��=&D=W�=:�=�=/� =-X =���<7"�<�Y�<��<��<��<`0�<�c�<���<���<���<"%�<�R�<�~�</��<n��<!��<N �<�D�<�g�<��<6��<���<L��<���<E�<�'�<�:�<�K�<'Z�<,f�<�o�<�v�<={�<�|�<�{�<�w�<!q�<Cg�<bZ�<^J�<*7�<� �<��<���<��<��<0}�<�Q�<�"�<H��<޹�<��<�A�<���<��<tp�<�"�<v��<|�<�"�<���<\d�<F��<b��<�)�<۸�<rD�<9̸<@P�<�е<oM�<�Ʋ<P<�<���<m�<��<[�<�V�<���<��<t�<�͢<P$�<ix�<�ɝ<!�<f�<���<��<�?�<��<�Ƒ<��<?G�<%��<���<���<�6�<�o�<�<߁<{�<��|<y<�ju<��q<6<n<��j<g<�uc<��_<�H\<�X<�U<ՋQ<N�M<�jJ<��F<?QC<�?<dA<<��8<�<5<E�1<*E.<��*<�['<z�#<C� <N<U�<�_<�<�<hj<~#	<w�<X�<���;҇�;�7�;���;G��;ʗ�;�~�;fs�;#w�;Ή�;
��;�ۻ;�;�k�;˪;N:�;���;�G�;��;���;�T�;�#�;[�;V�u;<�k;�a;�7X;�N;�E;��;;TZ2;b.);A ;�,;KW;ǜ;���:���:�!�:ց�:!�:Yצ:˖:5�:�yn:�pO:��0:N`:��96'�9��d9x��8�%i��!츻yg���]�㹶t��(�jD�7_��y��4���i������͑��I����h˺�8غ������TC���i�������g��F�$p$���*� �0�E�6���<�N�B��	I�*O�z"U�5+[�b2a��7g��;m�?s��Ay�jC����T�������ɧ��Y���Y���ͱ������8����  �  :h==��=)D=U�=9�=�=*� =1X =���<2"�<�Y�<��<��<��<g0�<yc�<���<���<~��<'%�<yR�<�~�<+��<q��<%��<M �<�D�<�g�<��<2��<���<:��<���<M�<�'�<�:�<�K�<#Z�<)f�<�o�<�v�<>{�<�|�<�{�<�w�<q�<Ig�<fZ�<ZJ�<-7�<� �<��<���<��<��</}�<�Q�<�"�<O��<ҹ�<��<�A�<���<��<mp�<�"�<o��<|�<�"�<���<cd�<D��<c��<~)�<�<hD�<:̸<JP�<�е<uM�<�Ʋ<Z<�<���<v�<��<[�<�V�<���<��<t�<�͢<J$�<^x�<ʝ<�<f�<���< ��<�?�<��<�Ƒ<��<GG�<��<���<���<�6�<�o�<秃<"߁<y�<��|<� y<�ju<��q<"<n<��j<�g<�uc<��_<tH\<�X<�U<�Q<I�M<�jJ<��F<KQC<�?<`A<<��8<�<5<W�1<E.<��*<\'<p�#<L� <M<c�<�_<�<Ѷ<Vj<�#	<d�<s�<���;އ�;�7�;���;t��;���;�~�;Us�;;w�;���;'��;ܻ;��;�k�;�ʪ;B:�;�;H�;��;���;�T�;e#�;��;#�u;l�k;%�a;�7X;�N;/E;ͤ;;UZ2;�.);H ;�,;vW;��;B��:6��:�!�:���:�:�צ:�ʖ:��:�xn:rO:��0:�`:���9�&�9��d9���8/�f��+��xg��﫹ª��s�t�(�3D�=_���y�y4���i������$�������\i˺�8غ:�享���B���i�������D��F�p$���*���0��6���<���B��	I�QO�A"U��+[��1a��7g��;m�,?s��Ay��C�8��������������m��������������"����  �  @h==��=+D=R�=<�=�=,� =.X =���<,"�<Z�<��<���<.��<R0�<�c�<���<���<��<$%�<zR�<�~�<4��<i��<*��<J �<�D�<�g�<��<A��<���<8��<���<I�<�'�<�:�<�K�<Z�<5f�<�o�<�v�<D{�<�|�<�{�<�w�<q�<Dg�<^Z�<YJ�<$7�<� �<��<���<��<��<8}�<�Q�<�"�<K��<չ�<��<�A�<���<��<rp�<�"�<w��<|�<�"�<���<dd�<P��<\��<�)�<鸻<iD�<8̸<GP�<�е<pM�<�Ʋ<U<�<���<p�<���<a�<�V�<���<��<t�<�͢<G$�<`x�<ʝ<(�<�e�<���<��<�?�<"��<�Ƒ<��<?G�< ��<���<���<�6�<�o�<맃<߁<��<��|<y<�ju<��q<0<n<��j<�g<�uc<��_<jH\< �X<�U<ϋQ<_�M<�jJ<��F<RQC<�?<nA<<��8<�<5<J�1<E.<��*<#\'<s�#<2� <w<9�<�_<�<ζ<Xj<�#	<e�<V�<���;���;�7�;���;N��;ؗ�;�~�;�s�;?w�;}��;#��;�ۻ;��;�k�;�ʪ;':�; ��;H�;��;̕�;�T�;#�;e�;2�u;I�k;��a;�7X;גN;IE;��;;�Z2;.);X ;"-;�V;2�;��:]��:s!�:{��:��:`צ:�ʖ:A�:�yn:�pO:Q�0:�`:��9~)�9�d9O��8�`g��*��yg�����xt���(��D��_���y��4��i��/�������M���`i˺�8غa�云��B��ui�{��F���� G��o$���*�w�0�H�6���<�[�B��	I�uO�H"U�d+[�X2a��7g��;m��>s�nAy��C���������������S�����������׶��F����  �  Ch==��=&D=S�=@�=�=5� ='X =���<,"�<�Y�<��<���</��<N0�<�c�<���<���<���<%�<�R�<|~�<:��<b��<&��<Q �<�D�<�g�<܈�<;��<���<N��<���<G�<�'�<�:�<�K�<Z�<0f�<�o�<�v�<G{�<�|�<�{�<�w�<!q�<Cg�<bZ�<eJ�<!7�<� �<��<���<��<��<9}�<�Q�<�"�<9��<��<��<�A�<���<��<wp�<�"�<���<|�<�"�<���<Xd�<L��<[��<�)�<ܸ�<yD�<;̸<AP�<�е<iM�<�Ʋ<G<�<���<r�<��<b�<�V�<���<��<&t�<�͢<O$�<kx�<�ɝ<3�<�e�<���<��<�?�<��<�Ƒ<��<4G�<2��<���<���<�6�<�o�<���<߁<��<y�|<y<�ju<��q<F<n<��j< g<�uc<��_<�H\<�X<�U<��Q<j�M<�jJ<��F<=QC<	�?<zA<<��8<�<5<.�1<BE.<��*<\'<��#<#� <y<1�<`<�<ݶ<pj<t#	<��<E�<��;���;�7�;���;R��;��;U~�;ys�;w�;ԉ�;��;�ۻ;6�;�k�;0˪;1:�;��;�G�;��;ו�;�T�;�#�;3�;Z�u;:�k;�a;88X;��N;�E;�;;�Z2;9.);J ;/-;�V;S�;���:���:�!�:���:^�:"צ:K˖:r�:�zn:�pO:��0:-`:��9}(�9��d9x��8 i�\�wxg�8򫹢��ru�{�(��D��_�{�y��4��i��Ɉ��6�������Wh˺�8غ���ڤ�D��"i����3�����F��o$��*���0���6�(�<���B��	I�\O��"U�+[�i2a�c7g�<m�?s��Ay��C��X�������ǧ��8���k���ձ��򶗻t����  �  >h==��=(D=U�=>�=�=2� =%X =���<0"�<�Y�<��<���<$��<X0�<�c�<���<���<{��<%�<�R�<�~�<4��<j��<%��<Q �<�D�<�g�<��<F��<���<E��<���<@�<�'�<�:�<�K�<Z�<5f�<�o�<�v�<A{�<�|�<�{�<�w�<!q�<Gg�<bZ�<`J�<7�<� �<��<���<��<��<4}�<�Q�<�"�<B��<ݹ�<��<�A�<���<��<vp�<�"�<v��<|�<�"�<���<nd�<R��<U��<�)�<⸻<oD�<4̸<FP�<�е<jM�<�Ʋ<[<�<���<s�<��<]�<�V�<���<��<t�<�͢<B$�<jx�<�ɝ<0�<f�<���<��<�?�<��<�Ƒ<��<.G�<*��<���<���<�6�<�o�<<߁<�<��|< y<�ju<��q<;<n<��j<g<�uc<��_<xH\<�X<�U<܋Q<V�M<�jJ<��F<FQC<�?<uA<<��8<�<5<#�1<E.<��*<\'<��#<6� <d<E�<`<�<�<Oj<d#	<}�<\�<���;�;�7�;���;`��;՗�;�~�;�s�;w�;���;'��;�ۻ;�;�k�; ˪;:�;!��;;H�;��;���;�T�;�#�;T�;V�u;]�k;�a;	8X;��N;~E;o�;;�Z2;�.);@ ; -;?W;+�;t��:���:� �:���:7�:�צ:5˖:��:myn:EqO:e�0:�`:Y��9%*�9��d9	��8�Fh��$�!|g���E��Hu�s�(�D��_�Q�y�q4��Xi��4�����������h˺y9غ������C��5i�,��������F��o$���*�M�0���6�i�<�x�B��	I�;O�g"U�L+[�B2a��7g��;m��>s��Ay��C����L���ǥ��ͧ��F�������ñ������-����  �  :h==��=-D=R�==�=�=(� =4X =���<6"�<�Y�<ݐ�<���<#��<W0�<zc�<���<���<���<0%�<sR�<�~�<)��<k��<)��<M �<�D�<�g�<��<2��<���<=��<���<G�<�'�<�:�<�K�<"Z�</f�<�o�<�v�<:{�<�|�<�{�<�w�<q�<Ng�<cZ�<^J�<37�<� �<��<���<��<��<1}�<�Q�<�"�<O��<ٹ�<��<�A�<���<��<jp�<�"�<r��<|�<�"�<}��<Wd�<G��<b��<�)�<<jD�<7̸<RP�<�е<vM�<�Ʋ<L<�<���<n�<��<]�<�V�<���<��<t�<�͢<Q$�<gx�<ʝ<�<�e�<���<��<�?�<��<�Ƒ<��<KG�<��<���<���<�6�<�o�<꧃<߁<x�<��|<� y<�ju<��q<=<n<��j<�g<�uc<��_<sH\<�X<�U<ɋQ<I�M<�jJ<��F<YQC<�?<qA<<��8<�<5<b�1<E.<��*<\'<g�#<6� <a<B�<�_<�<޶<fj<�#	<W�<p�<���;Ƈ�;�7�;���;X��;���;k~�;Vs�;Ew�;���;J��;�ۻ;��;�k�;�ʪ;;:�;��;�G�;��;���;�T�;s#�;~�;��u;��k;�a;�7X;P�N;lE;Ԥ;;TZ2;$.);. ;�,;W;��;A��:���:R"�:
��:��:�צ:rʖ:��:
yn:�qO:T�0:x_:���9;'�9̋d9���87�f�*츠zg���B���s�`�(��D�	_���y��4��bi��􇤺U���|����i˺"8غ���$���B���i�@�������?G��o$���*�_�0���6���<�?�B��	I��O�""U�m+[�2a��7g��;m�a?s��Ay��C� ��������������9��������������R����  �  Bh==��='D=T�=?�=�=(� =+X =���<-"�<�Y�<��<��<)��<]0�<�c�<���<���<z��<%�<rR�<�~�<2��<m��<!��<K �<�D�<�g�<��<>��<���<=��<���<D�<�'�<�:�<�K�< Z�<8f�<�o�<�v�<H{�<�|�<�{�<�w�<q�<Og�<`Z�<PJ�<7�<� �<��<���<��<��<7}�<�Q�<�"�<G��<չ�<��<�A�<���<��<qp�<�"�<q��<|�<�"�<���<cd�<R��<_��<�)�<⸻<pD�<6̸<FP�<�е<rM�<�Ʋ<X<�<���<u�< ��<Y�<�V�<���<��<t�<�͢<A$�<`x�<�ɝ<(�<f�<���<��<�?�<��<�Ƒ<��<7G�<��<���<���<�6�<�o�<姃<߁<��<��|< y<�ju<��q<8<n<��j<g<�uc<��_<sH\<�X<�U<��Q<h�M<�jJ<��F<AQC<�?<zA<<��8<�<5<<�1<E.<��*<
\'<z�#<@� <m<O�<�_<�<ζ<Lj<u#	<U�<q�<���;̇�;�7�;���;c��;���;�~�;�s�;>w�;���;!��;�ۻ;�;�k�;˪;5:�;-��;
H�;�;ە�;�T�;g#�;\�;�u;��k;��a;�7X;��N;HE;��;;�Z2;t.);] ;-;YW;�;���:`��:!�:��:��:
ئ:�ʖ:>�:�xn:wqO:�0:�a:���9*�9��d9���8:h��#�{g����[t���(�D�|_��y��4���i��򇤺����p����i˺L9غ��亗��nC��si���a��l��F��o$��*���0���6���<�5�B��	I�kO�~"U��+[�2a�o7g�{;m�?s�wAy��C�
���N�������ǧ��I�����������𶗻#����  �  �g=y=�=TC=i�=5=�=�� =�V =���<�<�V�<F��< ��<��<�+�<�^�<���<���<��<}�<�L�<Fx�<���<���<��<��< =�<�_�<{��<���<���<���<��<-�<3�<�/�<�@�<�N�<XZ�<�c�<>j�<Nn�<�o�<An�<�i�<�b�<�X�<^K�<;�<p'�<��<���<��<��<̓�<�k�<8@�<�<0��<���<Am�<1/�<+��<K��<�]�<�<���<%i�<��<���<�Q�<��<���<&�<���<\2�<T��<�>�<R��<K<�<ѵ�<�+�<c��<��<�y�<R�<�G�<���<
�<�f�<���<��<�l�<���<=�<�[�<���<��<�6�<�{�<��<� �<u@�<�<���<���<`2�<�k�<{��<)܁<�<ؒ|<m�x<2iu<I�q<=n<e�j<g<�yc<��_<�N\<g�X<5'U<P�Q<�N<^vJ<��F<-_C<�?<�Q<<��8<7O5<��1<�Y.<(�*<tr'<�$<�� <7<��<�{<(%<a�<��<�B	<�<I�<�(�;���;B~�;�<�;��;���;���;���;x��;3��;���;-�;n�;��;a�;���;��;���;;�;��;ڨ�;�w�;0V�;F�v;N�l; �b;c�X;5O;ɭE;lC<;��2;�);�� ;�;�;�.;��:�:�4�:א�:��:�٧:�Ǘ:��:=Zp:PEQ:��2:+:.�9Ao�9��j9$,�86 6p��9�a�\<��\�O2��'���B���]��x�!����薺�����}��)�ʺ��׺����D�U���>�c����d��$��N$��t*���0�&�6�Z�<�b�B���H��O��U�[��"a�*g��/m��4s��8y��<�����H���=���K���J��������������������  �  �g=y=�=WC=g�=8=�=� =�V =���<�<�V�<S��< ��<��<�+�<�^�<ʐ�<���<��<w�<�L�<Ox�<���<���<��<��< =�<�_�<���<���<���<���<��<1�<1�<�/�<w@�<�N�<^Z�<�c�<Sj�<Vn�<�o�<9n�<�i�<�b�<�X�<SK�<�:�<l'�<��<���<��</��<���<�k�<I@�<"�<7��<���<:m�</�<��<T��<�]�<
�<���<&i�<��<���<�Q�<��<ȃ�<�<���<[2�<W��<�>�<F��<X<�<ѵ�<�+�<t��<��<�y�<U�<�G�<}��<
�<�f�<���<��<~l�<���<F�<�[�<���<��<�6�<�{�<���<� �<u@�<�~�<���<���<\2�<�k�<q��<)܁<"�<��|<z�x<Giu<G�q<=n<s�j<�g<�yc<��_<�N\<��X<?'U<o�Q<	N<_vJ<��F<:_C<�?<�Q<<��8<�N5<��1<vY.<�*<�r'<$<�� <�6<��<�{<D%<E�<��<�B	<|<]�<�(�;���;S~�;�<�;��;���;���;���;���;��;���;-�;�m�;5��;$�;���;�;+��;X;�;�;٨�;�w�;CV�;�v;��l;Πb;��X;�4O;=�E;C<;�2;��);#� ;��;��;;/;�:�:~4�:|��:��:8ڧ:AǗ:��:�Yp:qEQ:��2:�:$�9�o�9��j9s�8a�6 ���a�G<��LṸ0� �'���B���]�j�x�F���_薺��������s�ʺ��׺,�人E�w����=����������#��N$��t*��0�!�6�7�<�s�B�u�H��O��U�Z[��"a��)g�`/m�x4s�X8y��<����,���c���5���u�������P���u���}����  �  �g={=�=ZC=b�=5=�=� =�V =���<�<�V�<H��<)��<��<,�<�^�<ʐ�<���<��<��<�L�<Wx�<���<���<��<��<=�<�_�<���<~��<���<���<��<6�<-�<�/�<o@�<�N�<YZ�<�c�<Bj�<Kn�<�o�<:n�<�i�<�b�<�X�<YK�<;�<�'�<��<���<��<-��<Ǔ�<�k�<K@�<�<<��<���<Pm�<)/�<!��<W��<�]�<�<���<,i�<��<���<�Q�<��<˃�<�<���<X2�<Y��<�>�<=��<]<�<ɵ�<�+�<c��<��<�y�<W�<�G�<s��<
�<�f�<���<��<~l�<���<2�<�[�<���<��<�6�<�{�< ��<� �<�@�<�~�<��<���<P2�<�k�<r��<.܁<�<�|<n�x<Ciu<G�q<�<n<��j<�g<�yc<��_<�N\<��X<0'U<[�Q<�N<fvJ<��F<C_C<��?<�Q<<��8<O5<��1<Y.<�*<zr'<�$<ț <�6<��<r{<D%<D�<��<�B	<�<k�<l(�;���;[~�;�<�;��;���;���;���;���;���;���;,-�;�m�;i��;�;���;��;	��;;�;��;�;�w�;SV�;ƈv;��l;��b;��X;�5O;C�E;�C<;|�2;��);i� ;��;��;�.;b�:�:�5�:_��:#�:mڧ:�Ɨ:��:�Yp:0FQ:}�2:�:��9n�9@�j9��8�K6��ฌ�a�:��m�"0��'���B���]��x����K薺D��p��g��K�ʺ@�׺$�亹E�L���k>���Q��P���#��N$��t*��0�S�6���<�>�B���H�[O�jU�N[��"a�,*g��/m��4s�i8y��<� �������m������v�������Z������������  �  �g=z=�=UC=h�=7=�=�� =�V =���<�<�V�<N��< ��<��<�+�<�^�<Ȑ�<���<��<p�<�L�<Gx�<���<���<��<��<"=�<�_�<���<���<���<���<��<1�<3�<�/�<}@�<�N�<YZ�<�c�<Mj�<Xn�<�o�<:n�<�i�<�b�<�X�<VK�< ;�<h'�<��<���<��<*��<Ó�<�k�<E@�<�<<��<���<9m�</�< ��<O��<�]�<	�<���<$i�<��<���<�Q�<��<�<�<���<Z2�<V��<�>�<E��<M<�<ֵ�<�+�<p��<��<�y�<S�<�G�<���<
�<�f�<���<��<�l�<���<@�<�[�<���<��<�6�<�{�<��<� �<p@�<�~�<���<���<\2�<�k�<t��<*܁<#�<�|<��x<(iu<M�q<=n<q�j<g<�yc<��_<�N\<b�X<O'U<k�Q<N<cvJ<��F<0_C<�?<�Q<<��8<%O5<{�1<wY.<$�*<�r'<$<�� <�6<��<�{<?%<L�<��<�B	<�<L�<�(�;��;F~�;�<�;��;���;���;��;���;��;���;-�;n�;<��;<�;���;��;D��;A;�;'�;ڨ�;�w�;1V�;;�v;|�l;�b;��X;�4O;D�E;�C<;��2;w�);H� ;��;l�;/;^�:�:h4�:���:�:�٧:�Ǘ:��:�Yp:EEQ:��2:+:f�9�o�9��j9�#�876+����a�o;����2�k�'�]�B�B�]�
�x�N����薺���n��?����ʺ��׺�亣E�����=�,��j������#��N$�qt*�	�0�O�6���<���B���H��O��U�D[��"a��)g�v/m�24s��8y�v<����/���=���7���h�����������T��������  �  �g=x=�=TC=h�=9=�=�� =�V =���<�<�V�<V��<��<��<�+�<�^�<���<���<'��<r�<�L�<Cx�<���<���<��<��<=�<�_�<x��<���<���<���<��<,�<3�<�/�<�@�<�N�<XZ�<�c�<;j�<Un�<�o�<Hn�<�i�<�b�<�X�<ZK�<;�<w'�<��<���<��<)��<���<�k�<C@�< �<,��<���<Km�<"/�<(��<M��<�]�< �<���<!i�<��<���<�Q�<��<Ã�<$�<���<[2�<U��<�>�<S��<N<�<Ե�<�+�<g��<��<�y�<Z�<�G�<���<
�<�f�<���<��<�l�<���<J�<�[�<���<��<�6�<�{�<���<� �<v@�<�~�<���<���<_2�<�k�<~��<%܁<$�<˒|<�x<0iu<X�q<=n<Z�j<	g<�yc<��_<�N\<m�X<G'U<E�Q<N<XvJ<��F<-_C<�?<�Q<<��8<'O5<��1<�Y.<�*<zr'<$<�� <�6<��<�{<.%<E�<ƈ<�B	<�<D�<�(�;���;W~�;�<�;��;���;���;���;���;B��;��;-�;n�;
��;P�;���;��;��;�:�;�;˨�;�w�;V�;T�v;x�l;�b;��X;E5O;��E;/C<;��2;p�);/� ;��;\�;2/;W�:��:�5�:��:��:�٧:�Ǘ:�:>[p:�DQ:l�2:I:��9io�9I�j9�*�8 �6:��f�a��<�����1���'���B�]�]�Ϲx�4���薺���M�����h�ʺ��׺Ғ�tE�F����=�/��;������#��N$�u*���0��6���<���B�o�H��O��U��[�#a��)g�0m�c4s��8y�I<� ���^���L���_���n���k�������e��������  �  �g={=�=WC=e�=7=�=� =�V =���<�<�V�<E��<"��<��<�+�<�^�<ΐ�<���< ��<x�<�L�<Tx�<���<���<��<��<"=�<�_�<���<���<���<���<��<8�<+�< 0�<q@�<�N�<\Z�<�c�<Ej�<Tn�<�o�<:n�<�i�<�b�<�X�<\K�<�:�<y'�<��<���<��<&��<ȓ�<�k�<C@�<�<;��<���<Im�</�<#��<U��<�]�<�<���<(i�<��<���<�Q�<��<���<�<���<V2�<Z��<�>�<?��<Q<�<Ե�<�+�<i��<��<�y�<T�<�G�<���<
�<�f�<���<��<{l�<���<5�<�[�<���<��<�6�<�{�<���<� �<�@�<�~�<��<���<Z2�<�k�<q��<+܁<$�<�|<��x<;iu<B�q<�<n<��j<�g<�yc<��_<�N\<y�X<F'U<a�Q<N<dvJ<��F<7_C<�?<�Q<<��8<�N5<��1<�Y.<�*<�r'<�$<�� <�6<��<o{<L%<>�<��<�B	<<f�<�(�;���;L~�;�<�;��;���;���;���;���;���;���;4-�;�m�;j��;�;���;	�;:��;;�;�;娊;�w�;"V�;&�v;��l;�b;}�X;Q5O;G�E;�C<;��2;V�);s� ;��;b�;�.;S�:��:k5�:V��:<�:Iڧ:�Ǘ:D�:�Yp:�EQ:i�2:;:��9�o�9��j9��8�>6E����a��:���ṏ1���'���B��]�n�x�L���p薺���q�����F�ʺ��׺*���E�M���Z>���'��p��$��N$��t*�ٕ0�в6�5�<�4�B���H�O��U�\[��"a��)g��/m�Y4s��8y��<����񡅻��������x�������h���h��������  �  �g== �=XC=i�=1=�=� =�V =���<�<�V�<I��<-��<���<,�<�^�<֐�<���<��<��<�L�<Vx�<���<���<��<��<)=�<�_�<���<{��<���<���<��<5�< �<0�<o@�<�N�<SZ�<�c�<Kj�<On�<�o�<5n�<�i�<�b�<�X�<_K�<�:�<}'�<��<���<��<4��<�<�k�<S@�<�<F��<���<Lm�< /�<%��<V��<�]�<�<���<.i�<��<���<�Q�<��<у�<�<���<M2�<V��<�>�<D��<]<�<ŵ�<�+�<e��<��<�y�<S�<�G�<v��<
�<�f�<���<��<xl�<���<4�<�[�<���<��<�6�<�{�<	��<� �<�@�<�~�<	��<���<^2�<�k�<k��<3܁<�<��|<k�x<3iu<c�q<�<n<��j<�g<�yc<��_<�N\<w�X</'U<s�Q<�N<vvJ<��F<<_C<�?<vQ<<��8<�N5<��1<oY.< �*<�r'<�$<ћ <�6<��<s{<[%<>�<��<�B	<�<i�<a(�;��;N~�;�<�;	�;���;���;���;���;��;���;'-�;�m�;���;�;㍥;��;(��;8;�;�;���;w�;HV�;�v;��l;-�b;��X;o5O;�E;�C<;��2;��);;� ;��;��;�.;�:l�:�5�:Ï�:a�:Sڧ:Ǘ:��:PYp:wFQ:
�2:�:Q�9�l�9��j9��8�6����a��9����0���'���B���]��x�?����薺���G�����.�ʺ�׺k��!F����Z>����߽�M���#��N$�^t*�B�0���6�6�<��B���H��O��U��[��"a�#*g�V/m��4s��8y�<�2���ꡅ�������������l���j�������t����  �  �g=~=�=SC=h�=4=�=� =�V =���<�<�V�<K��<.��<��<
,�<�^�<Ő�<���<!��<w�<�L�<Nx�<���<���<��<��<$=�<�_�<���<���<���<���<��<4�<5�<�/�<q@�<�N�<WZ�<�c�<Aj�<Nn�<�o�<Bn�<�i�<�b�<�X�<]K�< ;�<{'�<��<���<��<0��<Ɠ�<�k�<N@�<�<7��<���<Lm�</�<&��<P��<�]�<�<���<,i�<��<���<�Q�<��<ƃ�<�<���<]2�<[��<�>�<F��<P<�<ѵ�<�+�<b��<��<�y�<S�<�G�<{��<
�<�f�<���<��<�l�<���<7�<�[�<���<��<�6�<�{�<��<� �<�@�<�~�< ��<���<^2�<�k�<y��<1܁<�<�|<��x</iu<Y�q<�<n<v�j<
g<�yc<��_<�N\<h�X<F'U<`�Q<�N<qvJ<��F<'_C<�?<�Q<<��8<O5<��1<�Y.<�*<qr'<�$<қ <�6<��<{<9%<I�<��<�B	<�<Z�<w(�;���;B~�;�<�;��;���;���;���;���;��;p��;#-�;n�;<��;�;���;��;1��;;�;��;���;�w�;V�;&�v;v�l;�b;��X;d5O;g�E;�C<;��2;��);`� ;��;��;�.;�:H�:�5�:���:v�:�٧:VǗ:<�:uZp:DFQ:ˆ2:�:��9|n�9��j9��8��6��ม�a�=��.Ṻ1��'�7�B���]�p�x�����{薺e����������ʺ��׺�亠E����D>����y��8���#�O$��t*��0�̲6���<�Y�B���H��O��U�[��"a�(*g��/m�_4s��8y�E<�9���&���J���'�������o�������g��������  �  �g=t=	�=UC=g�=9=�=� =�V =���<�<�V�<L��<��<��<�+�<�^�<͐�<���<��<k�<�L�<Gx�<���<���<��<��<=�<�_�<}��<���<���<���<��<-�<2�<�/�<�@�<�N�<`Z�<�c�<Dj�<Yn�<�o�<Dn�<�i�<�b�<�X�<ZK�<�:�<l'�<��<���<"��<%��<ē�<�k�<=@�<$�<8��<���<<m�</�<%��<K��<�]�< �<���<"i�<��<���<�Q�<��<���<"�<���<X2�<R��<�>�<L��<D<�<ߵ�<�+�<p��<��<�y�<X�<�G�<���<
�<�f�<���<��<|l�<���<E�<�[�<���<��<�6�<�{�<���<� �<r@�<�~�<���<���<^2�<�k�<}��<܁<+�<ג|<��x<1iu<<�q<=n<m�j< g<�yc<��_<�N\<e�X<['U<O�Q<N<KvJ<��F<1_C<�?<�Q<<��8<O5<z�1<�Y.<�*<�r'<�$<�� <�6<��<�{<J%<?�<��<�B	<�<L�<�(�;���;W~�;�<�;��;���;���;��;l��; ��;���;-�;n�;5��;Z�;t��;�;E��;;�;+�;Ĩ�;�w�;V�;]�v;o�l;�b;��X;�4O;c�E;�C<;1�2;N�);P� ;��;/�;Q/;�:.�:�4�:L��:l�:�٧:�Ǘ:�:�Zp:�DQ:̇2:x:��9�q�9��j9+(�8��6J����a��;���	�)3�T�'���B�.�]���x�#���/薺�����h����ʺ�׺����E�b����=����2������#�xN$��t*�Е0�<�6���<���B�s�H��O��U��[�2#a��)g��/m�4s��8y��<�����9���_���A���H�����������=��������  �  �g=v=�=VC=f�=6=�=� =�V =���<�<�V�<P��<��<��<�+�<�^�<Ȑ�<���<&��<~�<�L�<Mx�<���<���<��<��<=�<�_�<u��<���<���<���<��<0�<-�<�/�<z@�<�N�<[Z�<�c�<@j�<Pn�<�o�<Bn�<�i�<�b�<�X�<`K�<;�<�'�<��<���<��<+��<ē�<�k�<G@�<�<7��<���<Om�<%/�<*��<N��<�]�<	�<���<&i�<��<���<�Q�<��<Ń�<�<���<V2�<U��<�>�<J��<W<�<ϵ�<�+�<k��<��<�y�<U�<�G�<|��<
�<�f�<���<��<{l�<���<A�<�[�<���<��<�6�<�{�<���<� �<�@�<�~�< ��<���<[2�<�k�<y��<#܁<&�<Ԓ|<m�x<@iu<K�q<=n<r�j<�g<�yc<��_<�N\<�X<6'U<H�Q<N<PvJ<��F<4_C<�?<�Q<<��8<O5<��1<�Y.<�*<r'<$<�� <7<��<�{<A%<:�<ň<�B	<�<X�<�(�;���;L~�;�<�;��;���;w��;���;���;&��;���;-�;�m�;6��;3�;���;�;���;;�;�;٨�;�w�;?V�;!�v;q�l;5�b;��X;�5O;r�E;�C<;��2;��);M� ;��;{�;	/;�::�:�5�:"��:��:�٧:WǗ:��:�Zp:sEQ:��2:�:��9o�9��j9�!�8�6���\�a��;��6
��0�F�'�P�B���]�O�x�#���\薺N����� ����ʺ��׺֒��E�����=���.������#��N$��t*���0���6���<�V�B���H� O��U�[�#a��)g��/m��4s�v8y�~<����.���q���3���m�������[������������  �  �g=}=�=PC=k�=5=�=� =�V =���<�<�V�<N��<*��<��<	,�<�^�<ǐ�<���<��<u�<�L�<Rx�<���<���<���<��<#=�<�_�<���<���<���<���<��<7�</�<�/�<m@�<�N�<[Z�<�c�<Wj�<Mn�<�o�<1n�<�i�<�b�<�X�<WK�<�:�<s'�<��<���<��<3��<œ�<�k�<O@�<�<B��<���<Bm�</�< ��<T��<�]�<�<~��</i�<��<���<�Q�<��<ǃ�<�<���<Y2�<[��<�>�<>��<S<�<е�<�+�<o��<��<�y�<H�<�G�<|��<
�<�f�<���<��<l�<���<6�<�[�<���<��<�6�<�{�<	��<� �<{@�<�~�<���<���<a2�<�k�<n��<2܁<�<�|<y�x<6iu<M�q<�<n<��j< g<�yc<��_<�N\<s�X<?'U<��Q<�N<nvJ<��F<_C< �?<�Q<<��8<O5<��1<qY.<%�*<tr'<$<ʛ <�6<��<z{<>%<N�<��<�B	<|<a�<�(�;��;~�;�<�;��;���;���;���;���;���;���;.-�;�m�;X��;��;���;�;7��;h;�;��;��;nw�;5V�;5�v;��l;�b;��X;5O;�E;�C<;}�2;��);Y� ;��;��;�.;��:��:�4�:_��:�:>ڧ:jǗ:��:�Xp:�FQ:��2:�:P�9zo�9��j9��8�65����a�w;��F�Y1�:�'���B�V�]���x��/閺���������h�ʺ��׺œ亮E�f���Q>����j��J���#�O$�^t*�+�0��6�5�<�t�B���H��O��U�n[��"a�*g�/m�z4s��8y�t<�3������_��������������t���v���U����  �  �g=z=�=UC=i�=3=�=� =�V =���<�<�V�<L��<��<��<�+�<�^�<ǐ�<���<��<��<�L�<Lx�<���<���<��<��<=�<�_�<z��<���<���<���<��<0�<'�<�/�<�@�<�N�<ZZ�<�c�<Dj�<Jn�<�o�<;n�<�i�<�b�<�X�<]K�<;�<|'�<��<���<��<)��<œ�<�k�<C@�<�<>��<���<Km�<+/�<(��<O��<�]�<
�<���<+i�<��<���<�Q�<��<�<!�<���<P2�<S��<�>�<P��<N<�<ϵ�<�+�<e��<��<�y�<S�<�G�<z��<
�<�f�<���<��<�l�<���<<�<�[�<���<��<�6�<�{�<��<� �<�@�<�~�<���<���<_2�<�k�<v��<+܁<�<�|<d�x<5iu<Q�q<=n<w�j<�g<�yc<��_<�N\<m�X<2'U<T�Q<�N<avJ<��F<1_C<�?<~Q<<��8<O5<��1<Y.<'�*<}r'<�$<�� <�6<��<�{<=%<T�<��<�B	<�<V�<|(�;��;G~�;�<�;��;���;���;���;���;4��;���;-�;�m�;G��;L�;���;�;�;;�;��;�;�w�;?V�;/�v;v�l;�b;�X;m5O;S�E;�C<;��2;k�);[� ;��;c�;�.;x�:7�:�5�:}��:��:�٧:RǗ:��:�Yp:FQ:L�2:�:(�9;o�9��j9�'�8�6�����a��:�����1�Z�'���B���]�n�x������薺�����-����ʺ��׺B��kE�v���>�%��Q������#��N$�kt*���0���6���<�k�B���H��O��U�/[��"a�3*g��/m��4s��8y�f<�򟂻#�������-���U�������������������  �  �g=x=�=WC=f�=8=�=� =�V =���<�<�V�<U��<��<��<�+�<�^�<Ɛ�<���<��<q�<�L�<Lx�<���<���<��<��<!=�<�_�<{��<���<���<���<��<7�<:�<�/�<w@�<�N�<hZ�<�c�<Oj�<^n�<�o�<@n�<�i�<�b�<�X�<WK�<�:�<m'�<��<���<!��<'��<Ó�<�k�<?@�<&�<5��<���<;m�</�<��<N��<�]�<�<���<"i�<��<���<�Q�<��<���<�<���<b2�<^��<�>�<E��<N<�<൲<�+�<��<��<�y�<W�<�G�<���<
�<�f�<���<��<|l�<���<K�<�[�<���<��<�6�<�{�<���<� �<u@�<�~�<���<���<[2�<�k�<v��<#܁</�<�|<}�x<Qiu<6�q<�<n<j�j<g<�yc<��_<�N\<��X<O'U<V�Q<&N<YvJ<��F<7_C<�?<�Q<<��8<O5<��1<vY.<�*<�r'<$<�� < 7<��<�{<<%<B�<��<�B	<�<V�<�(�;���;V~�;�<�;��;��;���;��;���;��;]��;.-�;"n�;��;'�;y��;9�;��;K;�;<�;ʨ�;�w�;6V�;#�v;w�l;�b;~�X;�4O;]�E;lC<;*�2;Z�);I� ;��;@�;Z/;��: �:�4�:&��:��:�٧:qǗ:��:�Zp:�DQ:A�2:,:��9�r�9��j9u�8{6b���a�F?��s��1�,�'�Q�B�X�]�q�x�����C薺R��u��&��/�ʺ��׺����E�����=�e��/������#��N$��t*��0�&�6�*�<�j�B�z�H�O��U�2[�#a�q)g��/m�k4s�28y��<����>���F���8�����������J���T��������  �  �g=z=�=UC=i�=3=�=� =�V =���<�<�V�<L��<��<��<�+�<�^�<ǐ�<���<��<��<�L�<Lx�<���<���<��<��<=�<�_�<z��<���<���<���<��<0�<'�<�/�<�@�<�N�<ZZ�<�c�<Dj�<Jn�<�o�<;n�<�i�<�b�<�X�<]K�<;�<|'�<��<���<��<)��<œ�<�k�<C@�<�<>��<���<Km�<+/�<(��<O��<�]�<
�<���<+i�<��<���<�Q�<��<�<!�<���<P2�<S��<�>�<P��<N<�<ϵ�<�+�<e��<��<�y�<S�<�G�<z��<
�<�f�<���<��<�l�<���<<�<�[�<���<��<�6�<�{�<��<� �<�@�<�~�<���<���<_2�<�k�<v��<+܁<�<�|<d�x<5iu<Q�q<=n<w�j<�g<�yc<��_<�N\<m�X<2'U<T�Q<�N<avJ<��F<1_C<�?<~Q<<��8<O5<��1<Y.<'�*<}r'<�$<�� <�6<��<�{<=%<T�<��<�B	<�<V�<|(�;��;G~�;�<�;��;���;���;���;���;4��;���;-�;�m�;G��;L�;���;�;�;;�;��;�;�w�;?V�;/�v;v�l;�b;�X;m5O;S�E;�C<;��2;k�);[� ;��;c�;�.;x�:7�:�5�:}��:��:�٧:RǗ:��:�Yp:FQ:L�2:�:(�9;o�9��j9�'�8�6�����a��:�����1�Z�'���B���]�n�x������薺�����-����ʺ��׺B��kE�v���>�%��Q������#��N$�kt*���0���6���<�k�B���H��O��U�/[��"a�3*g��/m��4s��8y�f<�򟂻#�������-���U�������������������  �  �g=}=�=PC=k�=5=�=� =�V =���<�<�V�<N��<*��<��<	,�<�^�<ǐ�<���<��<u�<�L�<Rx�<���<���<���<��<#=�<�_�<���<���<���<���<��<7�</�<�/�<m@�<�N�<[Z�<�c�<Wj�<Mn�<�o�<1n�<�i�<�b�<�X�<WK�<�:�<s'�<��<���<��<3��<œ�<�k�<O@�<�<B��<���<Bm�</�< ��<T��<�]�<�<~��</i�<��<���<�Q�<��<ǃ�<�<���<Y2�<[��<�>�<>��<S<�<е�<�+�<o��<��<�y�<H�<�G�<|��<
�<�f�<���<��<l�<���<6�<�[�<���<��<�6�<�{�<	��<� �<{@�<�~�<���<���<a2�<�k�<n��<2܁<�<�|<y�x<6iu<M�q<�<n<��j< g<�yc<��_<�N\<s�X<?'U<��Q<�N<nvJ<��F<_C< �?<�Q<<��8<O5<��1<qY.<%�*<tr'<$<ʛ <�6<��<z{<>%<N�<��<�B	<|<a�<�(�;��;~�;�<�;��;���;���;���;���;���;���;.-�;�m�;X��;��;���;�;7��;h;�;��;��;nw�;5V�;5�v;��l;�b;��X;5O;�E;�C<;}�2;��);Y� ;��;��;�.;��:��:�4�:_��:�:>ڧ:jǗ:��:�Xp:�FQ:��2:�:P�9zo�9��j9��8�65����a�w;��F�Y1�:�'���B�V�]���x��/閺���������h�ʺ��׺œ亮E�f���Q>����j��J���#�O$�^t*�+�0��6�5�<�t�B���H��O��U�n[��"a�*g�/m�z4s��8y�t<�3������_��������������t���v���U����  �  �g=v=�=VC=f�=6=�=� =�V =���<�<�V�<P��<��<��<�+�<�^�<Ȑ�<���<&��<~�<�L�<Mx�<���<���<��<��<=�<�_�<u��<���<���<���<��<0�<-�<�/�<z@�<�N�<[Z�<�c�<@j�<Pn�<�o�<Bn�<�i�<�b�<�X�<`K�<;�<�'�<��<���<��<+��<ē�<�k�<G@�<�<7��<���<Om�<%/�<*��<N��<�]�<	�<���<&i�<��<���<�Q�<��<Ń�<�<���<V2�<U��<�>�<J��<W<�<ϵ�<�+�<k��<��<�y�<U�<�G�<|��<
�<�f�<���<��<{l�<���<A�<�[�<���<��<�6�<�{�<���<� �<�@�<�~�< ��<���<[2�<�k�<y��<#܁<&�<Ԓ|<m�x<@iu<K�q<=n<r�j<�g<�yc<��_<�N\<�X<6'U<H�Q<N<PvJ<��F<4_C<�?<�Q<<��8<O5<��1<�Y.<�*<r'<$<�� <7<��<�{<A%<:�<ň<�B	<�<X�<�(�;���;L~�;�<�;��;���;w��;���;���;&��;���;-�;�m�;6��;3�;���;�;���;;�;�;٨�;�w�;?V�;!�v;q�l;5�b;��X;�5O;r�E;�C<;��2;��);M� ;��;{�;	/;�::�:�5�:"��:��:�٧:WǗ:��:�Zp:sEQ:��2:�:��9o�9��j9�!�8�6���\�a��;��6
��0�F�'�P�B���]�O�x�#���\薺N����� ����ʺ��׺֒��E�����=���.������#��N$��t*���0���6���<�V�B���H� O��U�[�#a��)g��/m��4s�v8y�~<����.���q���3���m�������[������������  �  �g=t=	�=UC=g�=9=�=� =�V =���<�<�V�<L��<��<��<�+�<�^�<͐�<���<��<k�<�L�<Gx�<���<���<��<��<=�<�_�<}��<���<���<���<��<-�<2�<�/�<�@�<�N�<`Z�<�c�<Dj�<Yn�<�o�<Dn�<�i�<�b�<�X�<ZK�<�:�<l'�<��<���<"��<%��<ē�<�k�<=@�<$�<8��<���<<m�</�<%��<K��<�]�< �<���<"i�<��<���<�Q�<��<���<"�<���<X2�<R��<�>�<L��<D<�<ߵ�<�+�<p��<��<�y�<X�<�G�<���<
�<�f�<���<��<|l�<���<E�<�[�<���<��<�6�<�{�<���<� �<r@�<�~�<���<���<^2�<�k�<}��<܁<+�<ג|<��x<1iu<<�q<=n<m�j< g<�yc<��_<�N\<e�X<['U<O�Q<N<KvJ<��F<1_C<�?<�Q<<��8<O5<z�1<�Y.<�*<�r'<�$<�� <�6<��<�{<J%<?�<��<�B	<�<L�<�(�;���;W~�;�<�;��;���;���;��;l��; ��;���;-�;n�;5��;Z�;t��;�;E��;;�;+�;Ĩ�;�w�;V�;]�v;o�l;�b;��X;�4O;c�E;�C<;1�2;N�);P� ;��;/�;Q/;�:.�:�4�:L��:l�:�٧:�Ǘ:�:�Zp:�DQ:̇2:x:��9�q�9��j9+(�8��6J����a��;���	�)3�T�'���B�.�]���x�#���/薺�����h����ʺ�׺����E�b����=����2������#�xN$��t*�Е0�<�6���<���B�s�H��O��U��[�2#a��)g��/m�4s��8y��<�����9���_���A���H�����������=��������  �  �g=~=�=SC=h�=4=�=� =�V =���<�<�V�<K��<.��<��<
,�<�^�<Ő�<���<!��<w�<�L�<Nx�<���<���<��<��<$=�<�_�<���<���<���<���<��<4�<5�<�/�<q@�<�N�<WZ�<�c�<Aj�<Nn�<�o�<Bn�<�i�<�b�<�X�<]K�< ;�<{'�<��<���<��<0��<Ɠ�<�k�<N@�<�<7��<���<Lm�</�<&��<P��<�]�<�<���<,i�<��<���<�Q�<��<ƃ�<�<���<]2�<[��<�>�<F��<P<�<ѵ�<�+�<b��<��<�y�<S�<�G�<{��<
�<�f�<���<��<�l�<���<7�<�[�<���<��<�6�<�{�<��<� �<�@�<�~�< ��<���<^2�<�k�<y��<1܁<�<�|<��x</iu<Y�q<�<n<v�j<
g<�yc<��_<�N\<h�X<F'U<`�Q<�N<qvJ<��F<'_C<�?<�Q<<��8<O5<��1<�Y.<�*<qr'<�$<қ <�6<��<{<9%<I�<��<�B	<�<Z�<w(�;���;B~�;�<�;��;���;���;���;���;��;p��;#-�;n�;<��;�;���;��;1��;;�;��;���;�w�;V�;&�v;v�l;�b;��X;d5O;g�E;�C<;��2;��);`� ;��;��;�.;�:H�:�5�:���:v�:�٧:VǗ:<�:uZp:DFQ:ˆ2:�:��9|n�9��j9��8��6��ม�a�=��.Ṻ1��'�7�B���]�p�x�����{薺e����������ʺ��׺�亠E����D>����y��8���#�O$��t*��0�̲6���<�Y�B���H��O��U�[��"a�(*g��/m�_4s��8y�E<�9���&���J���'�������o�������g��������  �  �g== �=XC=i�=1=�=� =�V =���<�<�V�<I��<-��<���<,�<�^�<֐�<���<��<��<�L�<Vx�<���<���<��<��<)=�<�_�<���<{��<���<���<��<5�< �<0�<o@�<�N�<SZ�<�c�<Kj�<On�<�o�<5n�<�i�<�b�<�X�<_K�<�:�<}'�<��<���<��<4��<�<�k�<S@�<�<F��<���<Lm�< /�<%��<V��<�]�<�<���<.i�<��<���<�Q�<��<у�<�<���<M2�<V��<�>�<D��<]<�<ŵ�<�+�<e��<��<�y�<S�<�G�<v��<
�<�f�<���<��<xl�<���<4�<�[�<���<��<�6�<�{�<	��<� �<�@�<�~�<	��<���<^2�<�k�<k��<3܁<�<��|<k�x<3iu<c�q<�<n<��j<�g<�yc<��_<�N\<w�X</'U<s�Q<�N<vvJ<��F<<_C<�?<vQ<<��8<�N5<��1<oY.< �*<�r'<�$<ћ <�6<��<s{<[%<>�<��<�B	<�<i�<a(�;��;N~�;�<�;	�;���;���;���;���;��;���;'-�;�m�;���;�;㍥;��;(��;8;�;�;���;w�;HV�;�v;��l;-�b;��X;o5O;�E;�C<;��2;��);;� ;��;��;�.;�:l�:�5�:Ï�:a�:Sڧ:Ǘ:��:PYp:wFQ:
�2:�:Q�9�l�9��j9��8�6����a��9����0���'���B���]��x�?����薺���G�����.�ʺ�׺k��!F����Z>����߽�M���#��N$�^t*�B�0���6�6�<��B���H��O��U��[��"a�#*g�V/m��4s��8y�<�2���ꡅ�������������l���j�������t����  �  �g={=�=WC=e�=7=�=� =�V =���<�<�V�<E��<"��<��<�+�<�^�<ΐ�<���< ��<x�<�L�<Tx�<���<���<��<��<"=�<�_�<���<���<���<���<��<8�<+�< 0�<q@�<�N�<\Z�<�c�<Ej�<Tn�<�o�<:n�<�i�<�b�<�X�<\K�<�:�<y'�<��<���<��<&��<ȓ�<�k�<C@�<�<;��<���<Im�</�<#��<U��<�]�<�<���<(i�<��<���<�Q�<��<���<�<���<V2�<Z��<�>�<?��<Q<�<Ե�<�+�<i��<��<�y�<T�<�G�<���<
�<�f�<���<��<{l�<���<5�<�[�<���<��<�6�<�{�<���<� �<�@�<�~�<��<���<Z2�<�k�<q��<+܁<$�<�|<��x<;iu<B�q<�<n<��j<�g<�yc<��_<�N\<y�X<F'U<a�Q<N<dvJ<��F<7_C<�?<�Q<<��8<�N5<��1<�Y.<�*<�r'<�$<�� <�6<��<o{<L%<>�<��<�B	<<f�<�(�;���;L~�;�<�;��;���;���;���;���;���;���;4-�;�m�;j��;�;���;	�;:��;;�;�;娊;�w�;"V�;&�v;��l;�b;}�X;Q5O;G�E;�C<;��2;V�);s� ;��;b�;�.;S�:��:k5�:V��:<�:Iڧ:�Ǘ:D�:�Yp:�EQ:i�2:;:��9�o�9��j9��8�>6E����a��:���ṏ1���'���B��]�n�x�L���p薺���q�����F�ʺ��׺*���E�M���Z>���'��p��$��N$��t*�ٕ0�в6�5�<�4�B���H�O��U�\[��"a��)g��/m�Y4s��8y��<����񡅻��������x�������h���h��������  �  �g=x=�=TC=h�=9=�=�� =�V =���<�<�V�<V��<��<��<�+�<�^�<���<���<'��<r�<�L�<Cx�<���<���<��<��<=�<�_�<x��<���<���<���<��<,�<3�<�/�<�@�<�N�<XZ�<�c�<;j�<Un�<�o�<Hn�<�i�<�b�<�X�<ZK�<;�<w'�<��<���<��<)��<���<�k�<C@�< �<,��<���<Km�<"/�<(��<M��<�]�< �<���<!i�<��<���<�Q�<��<Ã�<$�<���<[2�<U��<�>�<S��<N<�<Ե�<�+�<g��<��<�y�<Z�<�G�<���<
�<�f�<���<��<�l�<���<J�<�[�<���<��<�6�<�{�<���<� �<v@�<�~�<���<���<_2�<�k�<~��<%܁<$�<˒|<�x<0iu<X�q<=n<Z�j<	g<�yc<��_<�N\<m�X<G'U<E�Q<N<XvJ<��F<-_C<�?<�Q<<��8<'O5<��1<�Y.<�*<zr'<$<�� <�6<��<�{<.%<E�<ƈ<�B	<�<D�<�(�;���;W~�;�<�;��;���;���;���;���;B��;��;-�;n�;
��;P�;���;��;��;�:�;�;˨�;�w�;V�;T�v;x�l;�b;��X;E5O;��E;/C<;��2;p�);/� ;��;\�;2/;W�:��:�5�:��:��:�٧:�Ǘ:�:>[p:�DQ:l�2:I:��9io�9I�j9�*�8 �6:��f�a��<�����1���'���B�]�]�Ϲx�4���薺���M�����h�ʺ��׺Ғ�tE�F����=�/��;������#��N$�u*���0��6���<���B�o�H��O��U��[�#a��)g�0m�c4s��8y�I<� ���^���L���_���n���k�������e��������  �  �g=z=�=UC=h�=7=�=�� =�V =���<�<�V�<N��< ��<��<�+�<�^�<Ȑ�<���<��<p�<�L�<Gx�<���<���<��<��<"=�<�_�<���<���<���<���<��<1�<3�<�/�<}@�<�N�<YZ�<�c�<Mj�<Xn�<�o�<:n�<�i�<�b�<�X�<VK�< ;�<h'�<��<���<��<*��<Ó�<�k�<E@�<�<<��<���<9m�</�< ��<O��<�]�<	�<���<$i�<��<���<�Q�<��<�<�<���<Z2�<V��<�>�<E��<M<�<ֵ�<�+�<p��<��<�y�<S�<�G�<���<
�<�f�<���<��<�l�<���<@�<�[�<���<��<�6�<�{�<��<� �<p@�<�~�<���<���<\2�<�k�<t��<*܁<#�<�|<��x<(iu<M�q<=n<q�j<g<�yc<��_<�N\<b�X<O'U<k�Q<N<cvJ<��F<0_C<�?<�Q<<��8<%O5<{�1<wY.<$�*<�r'<$<�� <�6<��<�{<?%<L�<��<�B	<�<L�<�(�;��;F~�;�<�;��;���;���;��;���;��;���;-�;n�;<��;<�;���;��;D��;A;�;'�;ڨ�;�w�;1V�;;�v;|�l;�b;��X;�4O;D�E;�C<;��2;w�);H� ;��;l�;/;^�:�:h4�:���:�:�٧:�Ǘ:��:�Yp:EEQ:��2:+:f�9�o�9��j9�#�876+����a�o;����2�k�'�]�B�B�]�
�x�N����薺���n��?����ʺ��׺�亣E�����=�,��j������#��N$�qt*�	�0�O�6���<���B���H��O��U�D[��"a��)g�v/m�24s��8y�v<����/���=���7���h�����������T��������  �  �g={=�=ZC=b�=5=�=� =�V =���<�<�V�<H��<)��<��<,�<�^�<ʐ�<���<��<��<�L�<Wx�<���<���<��<��<=�<�_�<���<~��<���<���<��<6�<-�<�/�<o@�<�N�<YZ�<�c�<Bj�<Kn�<�o�<:n�<�i�<�b�<�X�<YK�<;�<�'�<��<���<��<-��<Ǔ�<�k�<K@�<�<<��<���<Pm�<)/�<!��<W��<�]�<�<���<,i�<��<���<�Q�<��<˃�<�<���<X2�<Y��<�>�<=��<]<�<ɵ�<�+�<c��<��<�y�<W�<�G�<s��<
�<�f�<���<��<~l�<���<2�<�[�<���<��<�6�<�{�< ��<� �<�@�<�~�<��<���<P2�<�k�<r��<.܁<�<�|<n�x<Ciu<G�q<�<n<��j<�g<�yc<��_<�N\<��X<0'U<[�Q<�N<fvJ<��F<C_C<��?<�Q<<��8<O5<��1<Y.<�*<zr'<�$<ț <�6<��<r{<D%<D�<��<�B	<�<k�<l(�;���;[~�;�<�;��;���;���;���;���;���;���;,-�;�m�;i��;�;���;��;	��;;�;��;�;�w�;SV�;ƈv;��l;��b;��X;�5O;C�E;�C<;|�2;��);i� ;��;��;�.;b�:�:�5�:_��:#�:mڧ:�Ɨ:��:�Yp:0FQ:}�2:�:��9n�9@�j9��8�K6��ฌ�a�:��m�"0��'���B���]��x����K薺D��p��g��K�ʺ@�׺$�亹E�L���k>���Q��P���#��N$��t*��0�S�6���<�>�B���H�[O�jU�N[��"a�,*g��/m��4s�i8y��<� �������m������v�������Z������������  �  �g=y=�=WC=g�=8=�=� =�V =���<�<�V�<S��< ��<��<�+�<�^�<ʐ�<���<��<w�<�L�<Ox�<���<���<��<��< =�<�_�<���<���<���<���<��<1�<1�<�/�<w@�<�N�<^Z�<�c�<Sj�<Vn�<�o�<9n�<�i�<�b�<�X�<SK�<�:�<l'�<��<���<��</��<���<�k�<I@�<"�<7��<���<:m�</�<��<T��<�]�<
�<���<&i�<��<���<�Q�<��<ȃ�<�<���<[2�<W��<�>�<F��<X<�<ѵ�<�+�<t��<��<�y�<U�<�G�<}��<
�<�f�<���<��<~l�<���<F�<�[�<���<��<�6�<�{�<���<� �<u@�<�~�<���<���<\2�<�k�<q��<)܁<"�<��|<z�x<Giu<G�q<=n<s�j<�g<�yc<��_<�N\<��X<?'U<o�Q<	N<_vJ<��F<:_C<�?<�Q<<��8<�N5<��1<vY.<�*<�r'<$<�� <�6<��<�{<D%<E�<��<�B	<|<]�<�(�;���;S~�;�<�;��;���;���;���;���;��;���;-�;�m�;5��;$�;���;�;+��;X;�;�;٨�;�w�;CV�;�v;��l;Πb;��X;�4O;=�E;C<;�2;��);#� ;��;��;;/;�:�:~4�:|��:��:8ڧ:AǗ:��:�Yp:qEQ:��2:�:$�9�o�9��j9s�8a�6 ���a�G<��LṸ0� �'���B���]�j�x�F���_薺��������s�ʺ��׺,�人E�w����=����������#��N$��t*��0�!�6�7�<�s�B�u�H��O��U�Z[��"a��)g�`/m�x4s�X8y��<����,���c���5���u�������P���u���}����  �  Pg=�=s�=�B=��=c~=�=� =�U =U��<k�<�S�<N��<���<���<d(�<+[�<���<W��<���<��<�G�<(s�<\��<���<+��<��<�6�<Y�<�y�<r��<=��<0��<��<���<��<'�<d7�<,E�<�P�<�Y�<�_�<�c�<�d�<c�<t^�<W�<�L�<?�<}.�<��<��<.��<���<S��<Յ�<�]�<�1�<��<m��<ǘ�<7^�< �<���<���<@N�<� �<��<�Y�<o �<?��<3B�<cݿ<�t�<�<���<�#�<���<;0�<��<P.�<&��<R�<7��<� �<m�<֪<�;�<잧<���<�[�</��<��<�b�<+��<S�< S�<���<�<a/�<�t�<���<���<�:�<�y�<U��<��<�.�<�h�<���<�ف<3�<܏|<i�x<hu<��q<�=n<�j<vg<�|c<1�_<�S\<��X<8.U<!�Q<�N< �J<H�F<�jC<O�?<�^<<��8<^5<I�1<1j.<��*<Մ'<&$<�� <L<b�<�<i<<O�<��<A\	<�<6�<�_�;Z�;��;�w�;E�; �;��;P �;��;	�;A=�;\o�;���;��;.b�;�ѥ;�Q�;���;��;�.�;��;c��;q��;�w;1m;�'c;�aY;��O;1F;�<;^x3;�G*;�5!;�?;Cd;q�;��:|��:�:m�:��:��:"��:E��:��q:��R:��3:Ԇ:Q��9m �9~p9�@�8�?�6q׸L]����s�޹�)���&�d�A���\���w��?���~��n���ڸ��F���<�ʺ�z׺�A�r�����y��_�7����i��3$�r[*��}0���6�z�<��B�7�H�Q�N�� U��[�0a�yg��%m��+s��0y��6���������0���٦��z���l���ٴ��q���yÚ��  �  Mg=�=n�=�B=��=^~=�=� =�U =T��<s�<�S�<_��<��<���<f(�<4[�<ь�<]��<���<��<�G�<1s�<S��<��<2��<��<�6�<Y�<�y�<c��<=��<,��<��<���<��<$'�<\7�<+E�<�P�<�Y�<`�<�c�<�d�<c�<�^�<W�<�L�<?�<u.�<��<��<:��<���<d��<���<�]�<�1�<��<x��<Ř�<>^�<��<���<��<<N�<� �<��<�Y�<g �<J��<>B�<Tݿ<�t�<	�<���<�#�<���<=0�<��<S.�<��<a�<<��<� �<�l�<֪< <�<䞧<���<�[�<,��<��<�b�<;��<X�<S�<���<��<t/�<�t�<���<���<�:�<�y�<W��<��<�.�<�h�<���<�ف<-�<��|<e�x<	hu<��q<�=n<�j<wg<	}c<(�_<�S\<x�X<,.U<A�Q<�N<�J<4�F<�jC<_�?<�^<<��8< ^5<W�1<0j.<��*<�'<H$<�� <�K<f�<�<�<<\�<{�<?\	<�<H�<�_�;��;'��;�w�;E�; �;	�; �;��;��;==�;so�;���;��;b�;�ѥ;�Q�;���;��;�.�;��;:��;���;�w;Im;�'c;�aY;��O;�0F;m�<;�x3;UH*; 5!;�>;�d;��;/�:X��:u�:�l�:+��:���:하:,��:��q:��R:��3:G�:��9��9Kp9�6�8���6�׸�I]�a����޹�)���&���A�7�\�}�w�[@���~������`���������ʺ�z׺�A�=�����Q��_���������W3$�3[*��}0�u�6�ж<���B�n�H��N�9 U�P[�Ea��g�k%m��+s�81y��6�����]���/�����������n���鴔�����:Ú��  �  Ig=�=l�=�B=��=[~=�=� =�U =L��<s�<�S�<U��< ��<���<{(�<![�<ˌ�<U��<���<��<�G�<;s�<L��<��<,��<��<�6�<Y�<�y�<Y��<L��<0��<��<���<��<%'�<W7�<?E�<�P�<�Y�<�_�<�c�<�d�<c�<�^�<W�<�L�<?�<t.�<��<��<>��<~��<h��<ȅ�<�]�<�1�<z�<z��<���<D^�<��<���<��<2N�<� �<��<�Y�<f �<@��<;B�<Sݿ<�t�<�<���<�#�<���<<0�<��<e.�<��<`�<3��<� �<	m�<
֪<<�<ڞ�<���<�[�<2��<��<�b�<9��<B�<S�<���<
�<n/�<�t�<���<���<�:�<�y�<b��<��<�.�<�h�<���<�ف<'�<�|<U�x<hu<�q<�=n<��j<Tg<}c<�_<�S\<��X<.U<<�Q<�N<�J<.�F<�jC<[�?<�^<<��8<�]5<f�1< j.<��*<ӄ'<2$<ӯ <�K<��<�<�<<K�<u�<M\	<�<]�<�_�;��;��;�w�;1E�;��;	�;���;��;�;0=�;^o�;���;��;�a�;ҥ;�Q�;���;��;�.�;��;.��;̚�;Ww;Bm;�'c;�aY;�O;�0F;��<;�w3;vH*;�5!;?; e;إ;\�:���:��:�l�:H��:���:L��:���:r�q:u�R:��3:��:H��9��9�p9�2�8���6�!׸9N]������޹8'�~�&���A�P�\���w��?���~��Z����������ޢʺ�z׺�A����!������^�G�������3$�)[*�~0�/�6��<���B���H�2�N�" U��[��a��g��%m�,s�1y�86�����b���t�����������I���Ĵ������BÚ��  �  Pg=�=k�=�B=��=`~=�=� =�U =N��<y�<�S�<L��<���<���<j(�<"[�<֌�<Y��<���<��<�G�</s�<V��<��<'��<��<�6�<Y�<�y�<`��<A��<,��<��<���<��<"'�<Z7�<3E�<�P�<�Y�<�_�<�c�<�d�<c�<�^�<W�<�L�<?�<q.�<��<��<F��<���<Z��<ą�<�]�<�1�<��<���<���<<^�<��<���<���<=N�<� �<��<�Y�<m �<D��<5B�<Tݿ<�t�<�<���<�#�<���<=0�<��<W.�<��<Y�<;��<� �<�l�<֪<<�<垧<���<�[�<0��<��<�b�<D��<H�<S�<���<�<b/�<�t�<���<���<�:�<�y�<[��<��<�.�<�h�<���<�ف<4�<�|<X�x<
hu<�q<�=n<��j<sg<}c<$�_<�S\<{�X<$.U<3�Q<�N<�J<+�F<�jC<^�?<�^<<��8<�]5<X�1<$j.<��*<�'<"$<�� <�K<n�<�<�<<S�<z�<H\	<�<E�<�_�;��;���;�w�;E�; �;��;	 �;��;��;:=�;uo�;���;��;b�;�ѥ;�Q�;���;��;�.�;��;-��;���;�w;2m;�'c;{aY;ǹO;�0F;��<;Ix3;H*;\5!;?;�d;0�;�:���:d�:|l�:*��:R��:���:��:��q:��R:j�3:x�:���9��9lp9S4�8V��6�׸�I]����Q�޹�(���&�y�A�H�\���w��@��4������E���������ʺ�z׺�A云��r�����|_�<��3��d��3$��Z*��}0�w�6���<���B�Y�H��N�f U�z[�2a�ug��%m� ,s�61y�h6�����e���6�����������c���ⴔ�����VÚ��  �  Rg=�=r�=�B=��=]~=�=� =�U =T��<m�<�S�<Z��<���<���<j(�</[�<̌�<V��<���<��<�G�<+s�<R��<���<7��<��<�6�<Y�<�y�<m��<?��<3��<��<���<��<'�<a7�<-E�<�P�<�Y�<�_�<�c�<�d�<c�<�^�<
W�<�L�<?�<x.�<��<��<5��<���<e��<ą�<�]�<�1�<��<s��<�<>^�<��<���<���<=N�<� �<"��<�Y�<n �<F��<7B�<]ݿ<�t�<�<���<�#�<���<60�<��<U.�<!��<U�<@��<� �<�l�<֪<�;�<㞧<���<�[�<,��<��<�b�<6��<U�<S�<���<�<q/�<�t�<���<���<�:�<�y�<Y��<��<�.�<�h�<���<�ف<5�<�|<p�x<hu<��q<�=n<�j<}g<�|c<(�_<�S\<}�X<:.U<'�Q<�N<�J<E�F<�jC<T�?<�^<<��8<^5<S�1<1j.<��*<�'<>$<�� <�K<n�<
�<�<<N�<~�<<\	<�<<�<�_�;z�;<��;�w�;�D�;" �;��;> �;��;�;*=�;Ko�;���;��;"b�;�ѥ;�Q�;���;��;�.�;��;o��;���;�w;�m;�'c;�aY;��O;�0F;A�<;rx3;]H*;`5!;?;�d;i�;��:,��:{�:�l�:���:ެ�:��:���:��q:��R:��3:͇:w��9(�9p9�<�83
�6�׸�M]�2����޹;)�S�&��A���\���w�x@��~��񦣺d���,���١ʺ�z׺�A云��P���j�y_�L��2�����3$�`[*��}0�|�6���<���B�}�H�;�N�W U��[��a�jg��%m��+s�1y��6���������"���ڦ������[���ߴ��n���nÚ��  �  Ng=�=p�=�B=��=^~=�=� =�U =R��<w�<�S�<Q��<���<���<u(�<$[�<̌�<Y��<���<��<�G�<6s�<S��< ��<0��<��<�6�<Y�<�y�<c��<<��<-��<��<���<��<%'�<Y7�<3E�<�P�<�Y�<�_�<�c�<�d�<c�<�^�<
W�<�L�<?�<r.�<��<��<B��<���<b��<Ņ�<�]�<�1�<�<��<���<@^�<��<���<���<=N�<� �<��<�Y�<n �<@��<:B�<Vݿ<�t�<	�<���<�#�<���<:0�<��<V.�<��<]�<:��<� �<m�<֪<�;�<䞧<���<�[�<*��<��<�b�<:��<I�<S�<���<�<j/�<�t�<���<���<�:�<�y�<a��<��<�.�<�h�<���<�ف</�<�|<e�x<hu< �q<�=n<�j<tg<	}c<�_<�S\<p�X<).U<3�Q<�N<�J<>�F<�jC<W�?<�^<<��8<^5<R�1<,j.<��*<ڄ'<+$<ͯ <�K<��<��<�<<T�<|�<<\	<�<R�<�_�;~�;��;�w�;E�; �;��; �;��;��;0=�;po�;���;��;b�;�ѥ;�Q�;���;��;�.�;��;O��;���;�w;m;�'c;�aY;׹O;�0F;��<;x3;JH*;k5!;?;�d; �;��:��:��:ul�:���:6��:���:��:Z�q:�R:�3:
�:��9/�9�p96�8���6�׸�J]�C����޹%)���&���A�k�\���w�@���~��Ȧ��^�������<�ʺ{׺�A争�������*_�P����!��3$�[*��}0�}�6�ܶ<���B�u�H�7�N�o U� [�'a��g��%m��+s�K1y�{6�����[���4�����������^�����������VÚ��  �  Jg=�=k�=�B=��=[~=�=� =�U =I��<x�<�S�<S��<���<���<u(�<%[�<ٌ�<V��<���<��<�G�<4s�<K��<	��<0��<��<�6�<Y�<�y�<Y��<H��<.��<��<���<��<&'�<R7�<BE�<�P�<�Y�< `�<�c�<�d�<c�<�^�<W�<�L�<?�<o.�<��<��<I��<���<d��<���<�]�<�1�<�<���<���<C^�<��<���<���<6N�<� �<��<�Y�<h �<C��<:B�<Kݿ<�t�<�<���<�#�<���<:0�<��<b.�<��<a�<4��<� �<�l�<֪<<�<ܞ�<���<�[�<2��<��<�b�<G��<G�<S�<���<�<k/�<�t�<���<���< ;�<�y�<^��<��<�.�<�h�<���<�ف<&�<��|<Z�x<hu<�q<�=n<�j<Jg<}c<�_<�S\<}�X<.U<A�Q<�N<�J<*�F<�jC<c�?<�^<<��8<�]5<l�1<j.<��*<�'</$<̯ <�K<��<��<�<<M�<v�<R\	<�<N�<�_�;��;��;�w�;E�;��;	�;���;��;�;-=�;io�;���;��;�a�;ҥ;gQ�;���;��;�.�;��;+��;Ӛ�;{w;�m;�'c;gaY;�O;[0F;��<;$x3;UH*;:5!;�>;�d; �;0�:U��:��:sl�:>��:��:���:���:|�q:f�R:��3:Z�:7��9��9Rp9�.�86��6"׸�L]����޹�'�ڥ&�u�A�&�\�-�w��@���~��+���⹰�����ޢʺ�z׺�A����6�����1_������ ��3$��Z*�&~0�'�6�$�<���B���H��N�" U�y[�'a��g�s%m��+s�>1y�6�����G���������������:���ߴ������:Ú��  �  Og=�=n�=�B=��=`~=�=� =�U =O��<p�<�S�<V��<���<���<p(�<&[�<ˌ�<V��<���<��<�G�<5s�<W��< ��</��<��<�6�<Y�<�y�<e��<D��<*��<��<���<��<''�<U7�<5E�<�P�<�Y�<�_�<�c�<�d�<c�<�^�<
W�<�L�<?�<s.�<��<��<<��<���<b��<ƅ�<�]�<�1�<��<z��<���<A^�<��<���<��<<N�<� �<��<�Y�<q �<A��<8B�<Vݿ<�t�<�<���<�#�<���<90�<��<\.�<��<Z�<9��<� �<�l�<֪<�;�<枧<���<�[�<,��<��<�b�<9��<L�<S�<���<�<l/�<�t�<���<���<�:�<�y�<`��<��<�.�<�h�<���<�ف<1�<�|<e�x<hu< �q<�=n<
�j<eg<}c<�_<�S\<}�X</.U<&�Q<�N<�J<4�F<�jC<V�?<�^<<��8<�]5<_�1<&j.<��*<݄'<5$<ǯ <�K<z�<��<�<<N�<��<C\	<�<Q�<�_�;}�;��;�w�;$E�; �;��; �;��;��;)=�;zo�;尶;��;�a�;�ѥ;�Q�;���;��;�.�;��;I��;���;�w;2m;�'c;�aY;�O;�0F;y�<;=x3;JH*;o5!;"?;�d;4�;Y�:��:��:el�:���:k��::��:d�q:��R:��3:�:���9f�9`p90�8]��6*׸J]�w����޹K(�:�&�Y�A���\�n�w�X@���~��Ŧ��>�������g�ʺ�z׺�A亢��$�����F_�������3$�=[*��}0�G�6�ٶ<���B�O�H�,�N�d U�H[�a��g��%m��+s�(1y�z6�ȝ��J���S�����������d���޴������oÚ��  �  Tg=�=n�=�B=��=a~=�=� =�U =X��<w�<�S�<Y��<��<���<f(�<0[�<ʌ�<\��<���<��<�G�<&s�<^��<��</��<��<�6�<Y�<�y�<g��<7��<3��<��<���<��<'�<a7�</E�<�P�<�Y�<�_�<�c�<�d�<c�<^�<W�<�L�<?�<y.�<��<��<9��<���<^��<���<�]�<�1�<��<t��<Ș�<=^�<  �<���<���<FN�<� �<��<�Y�<s �<C��<7B�<Wݿ<�t�<�<���<�#�<���<<0�<��<O.�<��<W�<@��<� �<�l�<֪<�;�<<���<�[�<.��<��<�b�<4��<U�<S�<���<��<m/�<�t�<���<���<�:�<�y�<T��<��<�.�<�h�<���<�ف<;�<�|<g�x<hu<�q<�=n<��j<pg<}c<(�_<�S\<j�X<3.U<'�Q<�N<�J<4�F<�jC<`�?<�^<<��8<^5<Q�1<9j.<��*<�'<<$<�� <�K<g�<�<~<<Y�<��<?\	<�<3�<�_�;��;��;�w�;E�;% �;��;' �;��;�;>=�;do�;ⰶ;��;"b�;�ѥ;�Q�;���;��;/�;��;J��;���;�w;�m;�'c;�aY;��O;�0F;a�<;{x3;%H*;A5!;?;�d;j�;��:���:r�:�l�:���:㬨:���:���:g�q:��R:�3:d�:p��9��9sp9.=�8�u�6׸�K]�����޹�)��&���A���\���w��@���~��Ѧ������g���.�ʺ�z׺�A�6��k���j��_���i���{3$�[*��}0���6���<��B�_�H���N�i U�I[�va�<g��%m��+s�X1y�g6�����p���<�����������S������}���mÚ��  �  Lg=�=p�=�B=��=[~=�=� =�U =L��<w�<�S�<Y��<���<���<m(�<+[�<Ό�<X��<���<��<�G�<3s�<K��< ��<1��<��<�6�<Y�<�y�<a��<H��<1��<��<���<��<'�<U7�<?E�<�P�<�Y�<�_�<�c�<�d�<c�<�^�<W�<�L�<?�<u.�<��<��<<��<���<e��<ǅ�<�]�<�1�<��<y��<���<=^�<��<���<���<5N�<� �<��<�Y�<h �<B��<5B�<Sݿ<�t�<�<���<�#�<���<00�<��<`.�<��<X�<8��<� �<m�<֪<�;�<ܞ�<���<�[�</��<��<�b�<:��<N�<S�<���<�<n/�<�t�<���<���<�:�<�y�<^��<��<�.�<�h�<���<�ف<+�<�|<a�x<hu<�q<�=n<��j<qg<}c<�_<�S\<�X<(.U<.�Q<�N<�J<>�F<�jC<Q�?<�^<<��8<^5<\�1<!j.<��*<؄'<;$<ɯ <�K<u�<�<�<<R�<p�<F\	<�<L�<�_�;}�;$��;�w�;E�;��;��; �;��;�;=�;eo�;찶;��;�a�;ҥ;�Q�;���;��;�.�;��;Q��;���;Yw;m;�'c;�aY;˹O;�0F;y�<;$x3;^H*;y5!;%?;�d;�;B�:���:m�:�l�:���:2��:|��:��:v�q:��R:��3:P�:��9��9�p9�4�8�)�6�׸�K]�����޹�'��&���A���\�j�w�&@���~��¦��۹������H�ʺ�z׺�A二�������\_���
����3$�[*�~0�n�6���<���B���H�e�N�7 U�'[�Sa��g��%m��+s�01y�(6�ѝ��q���;�������Ī��=���ܴ������^Ú��  �  Kg=�=k�=�B=��=]~=�=� =�U =G��<�<�S�<T��<���<���<n(�<%[�<Ռ�<]��<���<��<�G�<As�<K��<
��<.��<��<�6�<Y�<�y�<^��<?��<%��<��<���<��</'�<N7�<3E�<�P�<�Y�< `�<�c�<�d�<	c�<�^�<W�<�L�<?�<m.�<��<��<K��<���<e��<���<�]�<�1�<��<���<���<C^�<��<���<��<6N�<� �<��<�Y�<h �<E��<;B�<Pݿ<�t�<��<���<�#�<ë�<>0�<��<X.�<��<b�<9��<� �<m�<֪<<�<ܞ�<���<�[�</��<��<�b�<C��<J�<S�<���<�<k/�<�t�<���<���< ;�<�y�<g��<��<�.�<�h�<���<�ف<)�<�|<]�x<hu<��q<�=n<�j<bg<}c<�_<�S\<t�X<%.U<:�Q<�N<�J<+�F<�jC<]�?<�^<<��8<�]5<h�1<j.<��*<�'<1$<į <�K<w�<��<�<<[�<r�<L\	<�<i�<�_�;��;��;�w�;E�;��;	�; �;��;��;<=�;�o�;鰶;��;�a�;�ѥ;oQ�;���;��;�.�;��;!��;Ś�;jw;nm;�'c;YaY;�O;~0F;��<;3x3;^H*;)5!;�>;�d;�;.�:���:��:El�:5��:��:���:���:
�q:��R:��3:��:���9��97p9�*�8�.�6�׸yH]�.����޹�(�,�&�Z�A���\���w�+@����6���׹�������ʺ�z׺�A���x�����G_����1����3$��Z*�2~0�*�6��<���B�N�H�7�N�: U�r[��a��g��%m��+s�N1y��6�˝��3���Y�����������o���񴔻����GÚ��  �  Og=�=n�=�B=��=]~=�=� =�U =Q��<t�<�S�<Z��<���<���<p(�<.[�<ƌ�<X��<���<��<�G�<1s�<P��<��<2��<��<�6�<Y�<�y�<g��<<��<8��< ��<���<��<'�<d7�<3E�<�P�<�Y�<�_�<�c�<�d�<c�<�^�<W�<�L�<?�<v.�<��<��<7��<���<e��<ǅ�<�]�<�1�<��<s��<���<E^�< �<���<���<9N�<� �<��<�Y�<g �<D��<6B�<Zݿ<�t�<�<���<�#�<���<<0�<��<T.�<��<V�<<��<� �<m�<֪<<�<���<���<�[�<6��<��<�b�<1��<P�<S�<���<�<p/�<�t�<���<���< ;�<�y�<\��<��<�.�<�h�<���<�ف<0�<�|<e�x<hu<�q<�=n<�j<Qg<�|c<2�_<�S\<x�X<2.U<+�Q<�N<�J<7�F<�jC<`�?<�^<<��8<�]5<k�1<*j.<��*<ք'<=$<ǯ <�K<z�<�<v<<R�<�<V\	<�<I�<�_�;��;(��;�w�;�D�;
 �;��;% �;��;(�;J=�;4o�;���;��;/b�;�ѥ;�Q�;���;��;�.�;��;I��;���;�w;m;�'c;�aY;�O;�0F;W�<;Bx3;cH*;u5!;?;�d;4�;��:���:��:�l�:2��:<��:���:!��:O�q:4�R:��3:��:K��9\�9,p9�@�8�@�6k&׸RQ]������޹C)��&���A�4�\���w�	@���~��������������ʢʺEz׺iA亠�𺜞����C_�)�������3$�-[*��}0�'�6�۶<���B�s�H��N�C U�9[�Ga��g��%m��+s�1y�C6���������y���ަ��w���?���鴔����dÚ��  �  Sg=�=s�=�B=��=b~=�=� =�U =Y��<w�<�S�<^��<��<���<c(�<4[�<ƌ�<c��<���<��<�G�<5s�<\��<���<,��<��<�6�<#Y�<�y�<k��<4��<.��<��<���<��<'�<a7�<%E�<�P�<�Y�< `�<�c�<�d�<c�<w^�<	W�<�L�<?�<p.�<��<��<5��<���<a��<Å�<�]�<�1�<��<r��<͘�<8^�<��<���<��<?N�<� �<��<�Y�<h �<J��<2B�<[ݿ<�t�<�<���<�#�<˫�<*0�<��<J.�<!��<O�<D��<� �<m�<֪<�;�<랧<���<�[�<'��<��<�b�<2��<W�<S�<���<��<r/�<�t�<���<���<�:�<�y�<_��<��<�.�<�h�<���<�ف<8�<�|<i�x<hu<��q<�=n<�j<�g<�|c<�_<�S\<g�X<3.U<!�Q<�N<�J<K�F<�jC<I�?<�^<<��8<^5<J�1<9j.<��*<؄'<F$<�� <�K<a�<�<w<<g�<}�<6\	<�<P�<�_�;L�;��;�w�;�D�;2 �;��;4 �;��;�;�<�;o�;d��;{�;#b�;�ѥ;�Q�;���;��;�.�;��;i��;{��;�w;Qm;�'c;oaY;��O;%1F;A�<;ox3;?H*;V5!;�>;�d;~�;��:���:�:Ol�:���:���:��:A��:�q:�R:��3:?�:/��9��9�p9?�8���6K�ָmD]�.����޹�*�G�&���A�'�\���w�@���~������񸰺M���J�ʺ>{׺�A���𺇞��W��_���B�����3$�*[*�x}0���6�Զ<���B�K�H�T�N�� U��[��a�Ug��%m��+s�Q1y��6�������������Ʀ������s���
���~���yÚ��  �  Og=�=n�=�B=��=]~=�=� =�U =Q��<t�<�S�<Z��<���<���<p(�<.[�<ƌ�<X��<���<��<�G�<1s�<P��<��<2��<��<�6�<Y�<�y�<g��<<��<8��< ��<���<��<'�<d7�<3E�<�P�<�Y�<�_�<�c�<�d�<c�<�^�<W�<�L�<?�<v.�<��<��<7��<���<e��<ǅ�<�]�<�1�<��<s��<���<E^�< �<���<���<9N�<� �<��<�Y�<g �<D��<6B�<Zݿ<�t�<�<���<�#�<���<<0�<��<T.�<��<V�<<��<� �<m�<֪<<�<���<���<�[�<6��<��<�b�<1��<P�<S�<���<�<p/�<�t�<���<���< ;�<�y�<\��<��<�.�<�h�<���<�ف<0�<�|<e�x<hu<�q<�=n<�j<Qg<�|c<2�_<�S\<x�X<2.U<+�Q<�N<�J<7�F<�jC<`�?<�^<<��8<�]5<k�1<*j.<��*<ք'<=$<ǯ <�K<z�<�<v<<R�<�<V\	<�<I�<�_�;��;(��;�w�;�D�;
 �;��;% �;��;(�;J=�;4o�;���;��;/b�;�ѥ;�Q�;���;��;�.�;��;I��;���;�w;m;�'c;�aY;�O;�0F;W�<;Bx3;cH*;u5!;?;�d;4�;��:���:��:�l�:2��:<��:���:!��:O�q:4�R:��3:��:K��9\�9,p9�@�8�@�6k&׸RQ]������޹C)��&���A�4�\���w�	@���~��������������ʢʺEz׺iA亠�𺜞����C_�)�������3$�-[*��}0�'�6�۶<���B�s�H��N�C U�9[�Ga��g��%m��+s�1y�C6���������y���ަ��w���?���鴔����dÚ��  �  Kg=�=k�=�B=��=]~=�=� =�U =G��<�<�S�<T��<���<���<n(�<%[�<Ռ�<]��<���<��<�G�<As�<K��<
��<.��<��<�6�<Y�<�y�<^��<?��<%��<��<���<��</'�<N7�<3E�<�P�<�Y�< `�<�c�<�d�<	c�<�^�<W�<�L�<?�<m.�<��<��<K��<���<e��<���<�]�<�1�<��<���<���<C^�<��<���<��<6N�<� �<��<�Y�<h �<E��<;B�<Pݿ<�t�<��<���<�#�<ë�<>0�<��<X.�<��<b�<9��<� �<m�<֪<<�<ܞ�<���<�[�</��<��<�b�<C��<J�<S�<���<�<k/�<�t�<���<���< ;�<�y�<g��<��<�.�<�h�<���<�ف<)�<�|<]�x<hu<��q<�=n<�j<bg<}c<�_<�S\<t�X<%.U<:�Q<�N<�J<+�F<�jC<]�?<�^<<��8<�]5<h�1<j.<��*<�'<1$<į <�K<w�<��<�<<[�<r�<L\	<�<i�<�_�;��;��;�w�;E�;��;	�; �;��;��;<=�;�o�;鰶;��;�a�;�ѥ;oQ�;���;��;�.�;��;!��;Ś�;jw;nm;�'c;YaY;�O;~0F;��<;3x3;^H*;)5!;�>;�d;�;.�:���:��:El�:5��:��:���:���:
�q:��R:��3:��:���9��97p9�*�8�.�6�׸yH]�.����޹�(�,�&�Z�A���\���w�+@����6���׹�������ʺ�z׺�A���x�����G_����1����3$��Z*�2~0�*�6��<���B�N�H�7�N�: U�r[��a��g��%m��+s�N1y��6�˝��3���Y�����������o���񴔻����GÚ��  �  Lg=�=p�=�B=��=[~=�=� =�U =L��<w�<�S�<Y��<���<���<m(�<+[�<Ό�<X��<���<��<�G�<3s�<K��< ��<1��<��<�6�<Y�<�y�<a��<H��<1��<��<���<��<'�<U7�<?E�<�P�<�Y�<�_�<�c�<�d�<c�<�^�<W�<�L�<?�<u.�<��<��<<��<���<e��<ǅ�<�]�<�1�<��<y��<���<=^�<��<���<���<5N�<� �<��<�Y�<h �<B��<5B�<Sݿ<�t�<�<���<�#�<���<00�<��<`.�<��<X�<8��<� �<m�<֪<�;�<ܞ�<���<�[�</��<��<�b�<:��<N�<S�<���<�<n/�<�t�<���<���<�:�<�y�<^��<��<�.�<�h�<���<�ف<+�<�|<a�x<hu<�q<�=n<��j<qg<}c<�_<�S\<�X<(.U<.�Q<�N<�J<>�F<�jC<Q�?<�^<<��8<^5<\�1<!j.<��*<؄'<;$<ɯ <�K<u�<�<�<<R�<p�<F\	<�<L�<�_�;}�;$��;�w�;E�;��;��; �;��;�;=�;eo�;찶;��;�a�;ҥ;�Q�;���;��;�.�;��;Q��;���;Yw;m;�'c;�aY;˹O;�0F;y�<;$x3;^H*;y5!;%?;�d;�;B�:���:m�:�l�:���:2��:|��:��:v�q:��R:��3:P�:��9��9�p9�4�8�)�6�׸�K]�����޹�'��&���A���\�j�w�&@���~��¦��۹������H�ʺ�z׺�A二�������\_���
����3$�[*�~0�n�6���<���B���H�e�N�7 U�'[�Sa��g��%m��+s�01y�(6�ѝ��q���;�������Ī��=���ܴ������^Ú��  �  Tg=�=n�=�B=��=a~=�=� =�U =X��<w�<�S�<Y��<��<���<f(�<0[�<ʌ�<\��<���<��<�G�<&s�<^��<��</��<��<�6�<Y�<�y�<g��<7��<3��<��<���<��<'�<a7�</E�<�P�<�Y�<�_�<�c�<�d�<c�<^�<W�<�L�<?�<y.�<��<��<9��<���<^��<���<�]�<�1�<��<t��<Ș�<=^�<  �<���<���<FN�<� �<��<�Y�<s �<C��<7B�<Wݿ<�t�<�<���<�#�<���<<0�<��<O.�<��<W�<@��<� �<�l�<֪<�;�<<���<�[�<.��<��<�b�<4��<U�<S�<���<��<m/�<�t�<���<���<�:�<�y�<T��<��<�.�<�h�<���<�ف<;�<�|<g�x<hu<�q<�=n<��j<pg<}c<(�_<�S\<j�X<3.U<'�Q<�N<�J<4�F<�jC<`�?<�^<<��8<^5<Q�1<9j.<��*<�'<<$<�� <�K<g�<�<~<<Y�<��<?\	<�<3�<�_�;��;��;�w�;E�;% �;��;' �;��;�;>=�;do�;ⰶ;��;"b�;�ѥ;�Q�;���;��;/�;��;J��;���;�w;�m;�'c;�aY;��O;�0F;a�<;{x3;%H*;A5!;?;�d;j�;��:���:r�:�l�:���:㬨:���:���:g�q:��R:�3:d�:p��9��9sp9.=�8�u�6׸�K]�����޹�)��&���A���\���w��@���~��Ѧ������g���.�ʺ�z׺�A�6��k���j��_���i���{3$�[*��}0���6���<��B�_�H���N�i U�I[�va�<g��%m��+s�X1y�g6�����p���<�����������S������}���mÚ��  �  Og=�=n�=�B=��=`~=�=� =�U =O��<p�<�S�<V��<���<���<p(�<&[�<ˌ�<V��<���<��<�G�<5s�<W��< ��</��<��<�6�<Y�<�y�<e��<D��<*��<��<���<��<''�<U7�<5E�<�P�<�Y�<�_�<�c�<�d�<c�<�^�<
W�<�L�<?�<s.�<��<��<<��<���<b��<ƅ�<�]�<�1�<��<z��<���<A^�<��<���<��<<N�<� �<��<�Y�<q �<A��<8B�<Vݿ<�t�<�<���<�#�<���<90�<��<\.�<��<Z�<9��<� �<�l�<֪<�;�<枧<���<�[�<,��<��<�b�<9��<L�<S�<���<�<l/�<�t�<���<���<�:�<�y�<`��<��<�.�<�h�<���<�ف<1�<�|<e�x<hu< �q<�=n<
�j<eg<}c<�_<�S\<}�X</.U<&�Q<�N<�J<4�F<�jC<V�?<�^<<��8<�]5<_�1<&j.<��*<݄'<5$<ǯ <�K<z�<��<�<<N�<��<C\	<�<Q�<�_�;}�;��;�w�;$E�; �;��; �;��;��;)=�;zo�;尶;��;�a�;�ѥ;�Q�;���;��;�.�;��;I��;���;�w;2m;�'c;�aY;�O;�0F;y�<;=x3;JH*;o5!;"?;�d;4�;Y�:��:��:el�:���:k��::��:d�q:��R:��3:�:���9f�9`p90�8]��6*׸J]�w����޹K(�:�&�Y�A���\�n�w�X@���~��Ŧ��>�������g�ʺ�z׺�A亢��$�����F_�������3$�=[*��}0�G�6�ٶ<���B�O�H�,�N�d U�H[�a��g��%m��+s�(1y�z6�ȝ��J���S�����������d���޴������oÚ��  �  Jg=�=k�=�B=��=[~=�=� =�U =I��<x�<�S�<S��<���<���<u(�<%[�<ٌ�<V��<���<��<�G�<4s�<K��<	��<0��<��<�6�<Y�<�y�<Y��<H��<.��<��<���<��<&'�<R7�<BE�<�P�<�Y�< `�<�c�<�d�<c�<�^�<W�<�L�<?�<o.�<��<��<I��<���<d��<���<�]�<�1�<�<���<���<C^�<��<���<���<6N�<� �<��<�Y�<h �<C��<:B�<Kݿ<�t�<�<���<�#�<���<:0�<��<b.�<��<a�<4��<� �<�l�<֪<<�<ܞ�<���<�[�<2��<��<�b�<G��<G�<S�<���<�<k/�<�t�<���<���< ;�<�y�<^��<��<�.�<�h�<���<�ف<&�<��|<Z�x<hu<�q<�=n<�j<Jg<}c<�_<�S\<}�X<.U<A�Q<�N<�J<*�F<�jC<c�?<�^<<��8<�]5<l�1<j.<��*<�'</$<̯ <�K<��<��<�<<M�<v�<R\	<�<N�<�_�;��;��;�w�;E�;��;	�;���;��;�;-=�;io�;���;��;�a�;ҥ;gQ�;���;��;�.�;��;+��;Ӛ�;{w;�m;�'c;gaY;�O;[0F;��<;$x3;UH*;:5!;�>;�d; �;0�:U��:��:sl�:>��:��:���:���:|�q:f�R:��3:Z�:7��9��9Rp9�.�86��6"׸�L]����޹�'�ڥ&�u�A�&�\�-�w��@���~��+���⹰�����ޢʺ�z׺�A����6�����1_������ ��3$��Z*�&~0�'�6�$�<���B���H��N�" U�y[�'a��g�s%m��+s�>1y�6�����G���������������:���ߴ������:Ú��  �  Ng=�=p�=�B=��=^~=�=� =�U =R��<w�<�S�<Q��<���<���<u(�<$[�<̌�<Y��<���<��<�G�<6s�<S��< ��<0��<��<�6�<Y�<�y�<c��<<��<-��<��<���<��<%'�<Y7�<3E�<�P�<�Y�<�_�<�c�<�d�<c�<�^�<
W�<�L�<?�<r.�<��<��<B��<���<b��<Ņ�<�]�<�1�<�<��<���<@^�<��<���<���<=N�<� �<��<�Y�<n �<@��<:B�<Vݿ<�t�<	�<���<�#�<���<:0�<��<V.�<��<]�<:��<� �<m�<֪<�;�<䞧<���<�[�<*��<��<�b�<:��<I�<S�<���<�<j/�<�t�<���<���<�:�<�y�<a��<��<�.�<�h�<���<�ف</�<�|<e�x<hu< �q<�=n<�j<tg<	}c<�_<�S\<p�X<).U<3�Q<�N<�J<>�F<�jC<W�?<�^<<��8<^5<R�1<,j.<��*<ڄ'<+$<ͯ <�K<��<��<�<<T�<|�<<\	<�<R�<�_�;~�;��;�w�;E�; �;��; �;��;��;0=�;po�;���;��;b�;�ѥ;�Q�;���;��;�.�;��;O��;���;�w;m;�'c;�aY;׹O;�0F;��<;x3;JH*;k5!;?;�d; �;��:��:��:ul�:���:6��:���:��:Z�q:�R:�3:
�:��9/�9�p96�8���6�׸�J]�C����޹%)���&���A�k�\���w�@���~��Ȧ��^�������<�ʺ{׺�A争�������*_�P����!��3$�[*��}0�}�6�ܶ<���B�u�H�7�N�o U� [�'a��g��%m��+s�K1y�{6�����[���4�����������^�����������VÚ��  �  Rg=�=r�=�B=��=]~=�=� =�U =T��<m�<�S�<Z��<���<���<j(�</[�<̌�<V��<���<��<�G�<+s�<R��<���<7��<��<�6�<Y�<�y�<m��<?��<3��<��<���<��<'�<a7�<-E�<�P�<�Y�<�_�<�c�<�d�<c�<�^�<
W�<�L�<?�<x.�<��<��<5��<���<e��<ą�<�]�<�1�<��<s��<�<>^�<��<���<���<=N�<� �<"��<�Y�<n �<F��<7B�<]ݿ<�t�<�<���<�#�<���<60�<��<U.�<!��<U�<@��<� �<�l�<֪<�;�<㞧<���<�[�<,��<��<�b�<6��<U�<S�<���<�<q/�<�t�<���<���<�:�<�y�<Y��<��<�.�<�h�<���<�ف<5�<�|<p�x<hu<��q<�=n<�j<}g<�|c<(�_<�S\<}�X<:.U<'�Q<�N<�J<E�F<�jC<T�?<�^<<��8<^5<S�1<1j.<��*<�'<>$<�� <�K<n�<
�<�<<N�<~�<<\	<�<<�<�_�;z�;<��;�w�;�D�;" �;��;> �;��;�;*=�;Ko�;���;��;"b�;�ѥ;�Q�;���;��;�.�;��;o��;���;�w;�m;�'c;�aY;��O;�0F;A�<;rx3;]H*;`5!;?;�d;i�;��:,��:{�:�l�:���:ެ�:��:���:��q:��R:��3:͇:w��9(�9p9�<�83
�6�׸�M]�2����޹;)�S�&��A���\���w�x@��~��񦣺d���,���١ʺ�z׺�A云��P���j�y_�L��2�����3$�`[*��}0�|�6���<���B�}�H�;�N�W U��[��a�jg��%m��+s�1y��6���������"���ڦ������[���ߴ��n���nÚ��  �  Pg=�=k�=�B=��=`~=�=� =�U =N��<y�<�S�<L��<���<���<j(�<"[�<֌�<Y��<���<��<�G�</s�<V��<��<'��<��<�6�<Y�<�y�<`��<A��<,��<��<���<��<"'�<Z7�<3E�<�P�<�Y�<�_�<�c�<�d�<c�<�^�<W�<�L�<?�<q.�<��<��<F��<���<Z��<ą�<�]�<�1�<��<���<���<<^�<��<���<���<=N�<� �<��<�Y�<m �<D��<5B�<Tݿ<�t�<�<���<�#�<���<=0�<��<W.�<��<Y�<;��<� �<�l�<֪<<�<垧<���<�[�<0��<��<�b�<D��<H�<S�<���<�<b/�<�t�<���<���<�:�<�y�<[��<��<�.�<�h�<���<�ف<4�<�|<X�x<
hu<�q<�=n<��j<sg<}c<$�_<�S\<{�X<$.U<3�Q<�N<�J<+�F<�jC<^�?<�^<<��8<�]5<X�1<$j.<��*<�'<"$<�� <�K<n�<�<�<<S�<z�<H\	<�<E�<�_�;��;���;�w�;E�; �;��;	 �;��;��;:=�;uo�;���;��;b�;�ѥ;�Q�;���;��;�.�;��;-��;���;�w;2m;�'c;{aY;ǹO;�0F;��<;Ix3;H*;\5!;?;�d;0�;�:���:d�:|l�:*��:R��:���:��:��q:��R:j�3:x�:���9��9lp9S4�8V��6�׸�I]����Q�޹�(���&�y�A�H�\���w��@��4������E���������ʺ�z׺�A云��r�����|_�<��3��d��3$��Z*��}0�w�6���<���B�Y�H��N�f U�z[�2a�ug��%m� ,s�61y�h6�����e���6�����������c���ⴔ�����VÚ��  �  Ig=�=l�=�B=��=[~=�=� =�U =L��<s�<�S�<U��< ��<���<{(�<![�<ˌ�<U��<���<��<�G�<;s�<L��<��<,��<��<�6�<Y�<�y�<Y��<L��<0��<��<���<��<%'�<W7�<?E�<�P�<�Y�<�_�<�c�<�d�<c�<�^�<W�<�L�<?�<t.�<��<��<>��<~��<h��<ȅ�<�]�<�1�<z�<z��<���<D^�<��<���<��<2N�<� �<��<�Y�<f �<@��<;B�<Sݿ<�t�<�<���<�#�<���<<0�<��<e.�<��<`�<3��<� �<	m�<
֪<<�<ڞ�<���<�[�<2��<��<�b�<9��<B�<S�<���<
�<n/�<�t�<���<���<�:�<�y�<b��<��<�.�<�h�<���<�ف<'�<�|<U�x<hu<�q<�=n<��j<Tg<}c<�_<�S\<��X<.U<<�Q<�N<�J<.�F<�jC<[�?<�^<<��8<�]5<f�1< j.<��*<ӄ'<2$<ӯ <�K<��<�<�<<K�<u�<M\	<�<]�<�_�;��;��;�w�;1E�;��;	�;���;��;�;0=�;^o�;���;��;�a�;ҥ;�Q�;���;��;�.�;��;.��;̚�;Ww;Bm;�'c;�aY;�O;�0F;��<;�w3;vH*;�5!;?; e;إ;\�:���:��:�l�:H��:���:L��:���:r�q:u�R:��3:��:H��9��9�p9�2�8���6�!׸9N]������޹8'�~�&���A�P�\���w��?���~��Z����������ޢʺ�z׺�A����!������^�G�������3$�)[*�~0�/�6��<���B���H�2�N�" U��[��a��g��%m�,s�1y�86�����b���t�����������I���Ĵ������BÚ��  �  Mg=�=n�=�B=��=^~=�=� =�U =T��<s�<�S�<_��<��<���<f(�<4[�<ь�<]��<���<��<�G�<1s�<S��<��<2��<��<�6�<Y�<�y�<c��<=��<,��<��<���<��<$'�<\7�<+E�<�P�<�Y�<`�<�c�<�d�<c�<�^�<W�<�L�<?�<u.�<��<��<:��<���<d��<���<�]�<�1�<��<x��<Ř�<>^�<��<���<��<<N�<� �<��<�Y�<g �<J��<>B�<Tݿ<�t�<	�<���<�#�<���<=0�<��<S.�<��<a�<<��<� �<�l�<֪< <�<䞧<���<�[�<,��<��<�b�<;��<X�<S�<���<��<t/�<�t�<���<���<�:�<�y�<W��<��<�.�<�h�<���<�ف<-�<��|<e�x<	hu<��q<�=n<�j<wg<	}c<(�_<�S\<x�X<,.U<A�Q<�N<�J<4�F<�jC<_�?<�^<<��8< ^5<W�1<0j.<��*<�'<H$<�� <�K<f�<�<�<<\�<{�<?\	<�<H�<�_�;��;'��;�w�;E�; �;	�; �;��;��;==�;so�;���;��;b�;�ѥ;�Q�;���;��;�.�;��;:��;���;�w;Im;�'c;�aY;��O;�0F;m�<;�x3;UH*; 5!;�>;�d;��;/�:X��:u�:�l�:+��:���:하:,��:��q:��R:��3:G�:��9��9Kp9�6�8���6�׸�I]�a����޹�)���&���A�7�\�}�w�[@���~������`���������ʺ�z׺�A�=�����Q��_���������W3$�3[*��}0�u�6�ж<���B�n�H��N�9 U�P[�Ea��g�k%m��+s�81y��6�����]���/�����������n���鴔�����:Ú��  �  g=�=��=%B=	�=�}==!� =�T =v��<e�<�Q�<��<|��<+��<�%�<FX�<���<��<A��<-�<�C�<2o�<8��<���<���<�<�1�<T�<;t�<��<���<8��<���<y��<�<9 �<I0�<�=�<2I�<�Q�<�W�<�[�<V\�<qZ�<�U�<�M�<?C�<|5�<�$�<��<t��<���<��<���<�z�<�R�<�&�<;��<���<0��<�R�<8�<��<��<KB�<���<%��<�M�<x��<R��<F6�<�ѿ<�h�<]��<��<�<^��<%�<��<�#�<���<��<	��<���<;c�<�̪<�2�<앧<��<oS�<���<��<)[�<���<i��<aL�<b��<�<�)�<�o�<���<���<�6�<�u�<���<`��<�+�<f�<o��<�ׁ<��<��|<��x<?gu<��q<">n<�j<Vg<|c<k�_<�W\<H�X<�3U<*�Q<�N<l�J<l�F<xsC<��?<
i<<��8<�i5<��1<"w.<+<-�'<,'$<L� <5\<7�<��<�N<��<´<	p	<21<.�<��;51�;*��;���;�s�;�O�;9�;n1�;�7�;~L�;p�;���;��;�5�;Ԗ�;��;��;�;m��;�d�;#�;��;�π;u{w;�vm;D�c;s�Y;� P;ݖF;*=;S�3;��*;��!;�;��;;���:æ�:?��:�:��:�Q�:�6�:4I�:ss:��S:z5:\�:���9A8�9�"t9��8eR07��ϸ��Y�fL��3:ݹ�Y
�$�%�>+A��=\�^"w�xꈺ�+���X���l��?o���\ʺ�8׺�N��Ed�����tE����������T$��G*�k0��6�i�<��B���H�Z�N�_�T�[��a�Ng�9m� %s��*y��1�ț��F���W�����������﯑�ʵ��
����Ś��  �  �f=�=��=%B=�=�}==%� =�T =z��<z�<�Q�<��<~��<��<�%�<:X�<���<��<I��<6�<�C�<8o�<(��<���<���<�<�1�<�S�<It�<Β�<r��<0��<���<���<�<H �<G0�<�=�<I�<�Q�< X�<[�<S\�<`Z�<�U�<�M�<>C�<�5�<�$�<��<x��<���<���<���<�z�<�R�<�&�<3��<��<6��<�R�<=�<��<��<HB�<���<��<�M�<h��<N��<F6�<rѿ<�h�<X��<��<"�<m��<%�<��<w#�<h��<��<���<���<-c�<�̪<�2�<ߕ�<��<wS�<��<��<7[�<���<^��<hL�<F��<�<�)�<�o�<���<���<�6�<�u�<ĳ�<U��<�+�<f�<a��<�ׁ<��<��|<��x<gu<��q<'>n<4�j<dg<�c<r�_<�W\<�X<3U<J�Q<zN<p�J<S�F<zsC<��?<�h<<��8<�i5<��1<,w.<F+<&�'<$'$<Q� <�[<D�<x�<�N<�<Ѵ<p	<C1<9�<���;1�;��;���;�s�;�O�;99�;1�;R7�;^L�;9p�; ��; �;6�;˖�;��;���;�;t��;Nd�;#�;��;�π;o{w;�vm;��c;��Y;� P;��F;�*=;�3;Ī*;C�!;��;��;�;���:$��:���:g�:���:�Q�:H6�:DJ�:gs:��S:�5:ء:��9�0�9�t9#�8��07��ϸ^�Y�]J���;ݹ�[
�[�%��)A�u?\��#w�b눺n,��mW���m���n��k\ʺ8׺n�n���c�����9E�����������$��F*��j0�Ɋ6�5�<���B�O�H�*�N�D�T��[��a��g��m�T%s��+y��1���������<���F����������5���J���sŚ��  �  �f=�=��=#B=�=�}==� =�T =i��<v�<�Q�<��<���<��<�%�</X�<���<��<=��<1�<�C�<Ao�<��<���<���<�<�1�<�S�<\t�<Ғ�<���<5��<���<���<��<G �<?0�<�=�<I�<�Q�<X�<|[�<i\�<XZ�<�U�<�M�<;C�<�5�<�$�<��<f��<���<���<���<�z�<�R�<�&�<'��<��<#��<�R�<1�<��<��<>B�<���<��<�M�<l��<Q��<V6�<wѿ<�h�<S��<��<�<c��<%�<��<�#�<j��<��<�<���<>c�<|̪<�2�<ӕ�<��<kS�<���<��<+[�<���<S��<~L�<E��<�<�)�<�o�<���<���<�6�<�u�<ͳ�<N��<�+�<f�<_��<�ׁ<��<��|<��x<#gu<��q<>n<4�j<8g<�c<_�_<�W\<4�X<�3U<h�Q<\N<��J<S�F<psC<��?<�h<<��8<�i5<��1<	w.<@+<�'<'$<w� <�[<q�<c�<�N<��<��<p	<(1<K�<{��;�1�;���;���;�s�;[O�;�9�;1�;�7�;rL�; p�;㢼;��;6�;���;�;���;F�;���;Bd�;h#�;i�;�π;5{w;rvm;��c;"�Y;� P;h�F;�*=;��3;��*;��!;��;D�;;��:���:���:��:Z��:�Q�:�5�:�J�:/s:q�S:5:*�:���9�1�9�(t9��8۪07o�ϸ�Y�;K���;ݹOY
�"�%�{'A��@\�z"w�Tꈺ�,���V��Zn��~n��$]ʺ�8׺��1���c��O���D���� ������$��F*�}k0��6�Ȧ<�B�B���H�'�N�^�T��[��a�]g�sm�%s�k+y�Z1�雂���������P���Ҫ��ׯ��񵔻6���7Ś��  �  �f=�=��=%B=�=�}==� =�T =v��<o�<�Q�<��<���<��<�%�<7X�<���<��<I��<?�<�C�<Co�<*��<���<���<�<�1�<�S�<Kt�<ђ�<}��<-��<���<���<�<K �<>0�<�=�<I�<�Q�<�W�<|[�<\\�<dZ�<�U�<�M�<CC�<�5�<�$�<��<p��<���<��<���<�z�<�R�<�&�<2��<��<,��<�R�<>�<��< ��<JB�<���<��<�M�<g��<M��<I6�<yѿ<�h�<R��<��<�<k��<%�<	��<#�<k��<��<���<���<<c�<�̪<�2�<���< ��<lS�<��<��<-[�<��<\��<nL�<G��<�<�)�<�o�<���<���<�6�<�u�<ʳ�<W��<�+�<f�<h��<�ׁ<��<��|<��x<'gu<��q<>n<>�j<Ig<�c<j�_<�W\<2�X<�3U<F�Q<vN<z�J<`�F<xsC<��?<�h<<��8<�i5<��1<#w.<1+<;�'<'$<[� <�[<R�<r�<�N<��<Ѵ<,p	<&1<P�<���;l1�;��;ĥ�;�s�;�O�;A9�;1�;~7�;TL�;8p�;���;��;&6�;���;��;���;�;m��;Bd�;3#�;��;�π;�{w;�vm;��c;v�Y;b!P;��F;�*=;�3;��*;_�!;��;��;�;��:���:���:u�:���:�Q�:g6�:�I�:�s:#�S:v5:��:���9a2�93 t9�
�8��07��ϸ��Y��I���<ݹ�Z
��%��)A��?\��#w�iꈺv,���W���m��]n��]ʺ�7׺:�	��Tc����
E����u�����B$�8G*�k0�V�6���<�V�B�:�H�'�N�J�T�U[�Oa�	g��m�E%s�\+y��1�ڛ��䞅�s���5��������������H���zŚ��  �  �f=�=��=%B=�=�}=="� =�T =u��<k�<�Q�<��<���<��<�%�<;X�<���<��<@��<2�<�C�<4o�<-��<���<���<�<�1�<�S�<Ct�<ޒ�<x��<3��<���<���<�<A �<Q0�<�=�<&I�<�Q�<X�<�[�<P\�<oZ�<�U�<�M�<6C�<�5�<�$�<��<r��<���< ��<���<�z�<�R�<�&�<5��<���<-��<�R�<7�<��<��<NB�<���<#��<�M�<o��<V��<L6�<�ѿ<�h�<b��<��<�<a��<%�<��<z#�<x��<��<��<���<6c�<�̪<�2�<啧<��<rS�<���<��<-[�<���<_��<lL�<Q��<�<�)�<�o�<���<���<�6�<�u�<���<R��<�+�<	f�<m��<�ׁ<��<��|<��x<(gu<��q<5>n<#�j<Mg<�c<��_<�W\<.�X<�3U<>�Q<�N<c�J<j�F<xsC<��?<�h<<��8<�i5<��1<!w.<)+<-�'<$'$<Y� <\<L�<y�<�N<��<��<p	<71<2�<���;^1�;��;���;�s�;�O�;"9�;Q1�;i7�;kL�;Cp�;֢�;��;�5�;�;��;↠;)�;���;rd�;#�;��;�π;�{w;Jvm;~�c;l�Y;� P;ǖF;>*=;�3;̪*;��!;؞;��;�;��:���:���:��:h��:'Q�:�6�:AI�:4s:��S:`5:Ѣ:[��95�9�t9��8F�07��ϸ'�Y�WJ���:ݹH[
�k�%�9*A�>\��#w��ꈺ�+��X��<m��8o���\ʺl8׺���;d�����E�.��s�����c$�nG*�k0��6�e�<���B�c�H�)�N�q�T�+[��a�yg��m�
%s�T+y��1��������j���g������������������Ś��  �  �f=�=��=B=�=�}==$� =�T =t��<z�<�Q�<��<���<��<�%�<:X�<���<��<C��<3�<�C�<4o�<.��<���<���<�<�1�<�S�<Gt�<ؒ�<z��<7��<���<���<
�<> �<H0�<�=�<I�<�Q�<�W�<�[�<^\�<cZ�<�U�<�M�<<C�<�5�<�$�<��<r��<���<���<���<�z�<�R�<�&�<1��<��<1��<�R�<8�<��<��<PB�<���<��<�M�<p��<H��<L6�<wѿ<�h�<\��<��< �<i��<%�<��<}#�<o��<��<���<���<:c�<|̪<�2�<啧<��<sS�<��<��<6[�<���<]��<sL�<G��<�<�)�<�o�<���<���<�6�<�u�<���<V��<�+�< f�<g��<�ׁ<��<��|<��x<gu<��q<>n<�j<cg<�c<g�_<�W\<%�X<�3U<<�Q<}N<��J<c�F<[sC<��?<�h<<��8<�i5<��1<w.<F+<�'<%'$<b� <�[<[�<y�<�N<�<Ŵ<p	<;1<1�<���;�1�;���;���;�s�;O�;29�;:1�;p7�;|L�;,p�;颼;��;�5�;Ζ�;��;���;&�;[��;dd�;;#�;��;�π;�{w;{vm;��c;{�Y;� P;͖F;�*=;��3;�*;f�!;��;�;�;���:ڦ�:���:�:���:pQ�:�6�:nI�:ys:Q�S:�5:�:M��92�9$!t9i�8ju07�ϸ:�Y�K���:ݹ�Z
�v�%��)A�M@\��"w��ꈺ�,���W��Am��!o���\ʺ>8׺��v���c������D����s������$��F*�#k0��6�G�<���B�D�H���N���T�^[�6a��g�m�!%s��+y��1�ӛ��*���>���t���ê��ᯑ����$����Ś��  �  �f=�=��=$B=�=�}== � =�T =q��<p�<�Q�<��<���<��<�%�<5X�<���<��<C��<=�<�C�<<o�<&��<���<���<�<�1�<�S�<Xt�<В�<}��</��<���<���<�<H �<=0�<�=�<I�<�Q�<X�<�[�<\\�<aZ�<�U�<�M�<@C�<�5�<�$�<��<i��<���<���<���<�z�<�R�<�&�<-��<��<&��<�R�<;�<��<��<FB�<���<��<�M�<m��<O��<X6�<qѿ<�h�<Q��<��<�<j��<%�<	��<�#�<g��<��<���<���<:c�<�̪<�2�<ܕ�<��<lS�<	��<��<*[�<���<W��<qL�<N��<�<�)�<�o�<���<���<�6�<�u�<ó�<T��<�+�<f�<e��<�ׁ<��<��|<��x<gu<��q<>n<6�j<Ng<�c<c�_<�W\<"�X<�3U<Y�Q<}N<z�J<^�F<vsC<��?<�h<<��8<�i5<��1<w.<3+<$�'<'$<e� <	\<X�<n�<�N<��<ƴ<)p	<,1<C�<���;�1�;���;���;�s�;�O�;v9�;1�;{7�;]L�;*p�;���;��;6�;���;��;���;O�;}��;Qd�;3#�;��;�π;h{w;�vm;��c;m�Y;L!P;�F;�*=;��3;�*;��!;̞;	�;�;���:$��:���:B�:Z��:�Q�:-6�:#J�:ms:�S:%5:�:x��9e0�9�"t9/	�8@�07v�ϸ̸Y�HJ���<ݹ�Z
���%��'A��?\�5#w��ꈺ�,��OW���m���n��]ʺ�7׺��<���c��.���D�F��R������$�1G*�Jk0�t�6��<���B�P�H�+�N�A�T�q[�Ka��g��m�%s��+y��1�䛂�����i���<���ʪ���������+���UŚ��  �  �f=�=��='B=	�=�}== � =�T =t��<p�<�Q�<��<|��<��<�%�<;X�<���<��<>��<2�<�C�<>o�<(��<���<���<�<�1�<�S�<Et�<֒�<���<0��<���<���<��<J �<C0�<�=�<!I�<�Q�<�W�<�[�<U\�<kZ�<�U�<�M�<@C�<�5�<�$�<��<q��<���<��<���<�z�<�R�<�&�<7��<��<-��<�R�<5�<��<��<EB�<���<��<�M�<q��<K��<N6�<|ѿ<�h�<V��<��<�<d��<%�<��<�#�<o��<��<���<���<7c�<�̪<�2�<ޕ�<��<pS�< ��<��<0[�<���<a��<fL�<T��<�<�)�<�o�<���<���<�6�<�u�<ȳ�<V��<�+�<f�<k��<�ׁ<��<��|<��x<*gu<��q<>n<:�j<<g<�c<k�_<�W\<7�X<�3U<9�Q<�N<l�J<h�F<�sC<��?<�h<<��8<�i5<��1< w.<3+<1�'<"'$<L� <\<?�<z�<�N<��<��<p	<31<F�<���;G1�;��;���;�s�;�O�;+9�;/1�;�7�;`L�;.p�;뢼;��;%6�;���;��;ˆ�;7�;f��;ld�;#�;��;�π;F{w;�vm;��c;P�Y;� P;��F;p*=;$�3;��*;��!;�;��;�;c��:���:���:��:���:�Q�:6�:|I�:�s:l�S:�5:z�:���9E3�9d#t9x�8�07R�ϸ��Y�5J��K<ݹ�Y
�x�%��)A�t?\�##w��ꈺ�+��>X���m���n���\ʺa8׺�ں��c�����HE���������V$�CG*�k0���6���<�j�B�D�H���N�3�T�@[��a��g�m�%s�O+y��1�қ��힅�����=����������뵔�#����Ś��  �  �f=�=��="B=�=�}==&� =�T =x��<s�<�Q�<��<~��<��<�%�<FX�<���<��<A��<9�<�C�<.o�<1��<���<���<�<�1�<�S�<Ht�<ؒ�<s��<6��<���<���<�<D �<E0�<�=�<I�<�Q�<�W�<�[�<S\�<kZ�<�U�<�M�<;C�<�5�<�$�<��<{��<���<��<���<�z�<�R�<�&�<<��<��<9��<�R�<C�<��<��<TB�<���<��<�M�<o��<I��<J6�<wѿ<�h�<Y��<��<�<i��<
%�<��<v#�<p��<��<���<���<1c�<�̪<�2�<镧<��<vS�<	��<��<;[�<�<k��<iL�<K��<�<�)�<�o�<���<���<�6�<�u�<���<V��<�+�<f�<j��<�ׁ<��<��|<��x<gu<��q<>n<+�j<Ug<�c<i�_<�W\<�X<�3U<=�Q<�N<r�J<c�F<msC<��?<�h<<��8<�i5<��1<'w.<8+<�'<:'$<O� <\<G�<��<�N<�<��<!p	<F1<%�<ϊ�;b1�;��;���;�s�;�O�;59�;71�;V7�;xL�;0p�;�;��;6�;Ė�;��;���;$�;Y��;id�;#�;��;�π;�{w;lvm;p�c;��Y;� P;�F;W*=;5�3;ɪ*;Y�!;��;��;%;��:X��:���:��:U��:BQ�:7�:HI�:�s:��S:r5:3�:���9�1�9�t9��8�07Y�ϸ��Y��J��;ݹ�[
�^�%�*A��?\�g#w�눺W,��X���l��so��|\ʺ�7׺��-��hd�����2E�^�����r���$�HG*��j0��6��<�ʾB�@�H�	�N���T�G[��a��g�m�%s��+y��1�ӛ��
���Z���V�������ꯑ�"���!����Ś��  �  �f=�=��=#B=�=�}==� =�T =l��<w�<�Q�<��<���<��<�%�<7X�<���<��<:��<7�<�C�<<o�<+��<���<���<�<�1�<�S�<[t�<֒�<|��<8��<���<���<��<E �<B0�<�=�<I�<�Q�<X�<�[�<`\�<eZ�<�U�<�M�<AC�<�5�<�$�<��<n��<���<���<���<�z�<�R�<�&�<.��<��<-��<�R�<9�<��<��<FB�<���<��<�M�<p��<S��<\6�<wѿ<�h�<V��<��<�<d��<%�<��<�#�<n��<��<���<���<<c�<�̪<�2�<ߕ�<��<hS�<��<��<3[�<�<Y��<tL�<M��<�<�)�<�o�<���<���<�6�<�u�<³�<X��<�+�<	f�<g��<�ׁ<��<��|<��x<gu<��q<>n<0�j<@g<�c<a�_<�W\< �X<�3U<`�Q<mN<��J<a�F<qsC<��?<�h<<��8<�i5<��1<w.<@+<�'<''$<f� <\<`�<q�<�N<�<��<p	<$1<B�<���;~1�;��;���;�s�;xO�;�9�;11�;x7�;�L�;!p�;뢼;��;6�;���;�;���;`�;���;Yd�;A#�;��;�π;q{w;�vm;k�c;e�Y;� P;��F;�*=;��3;��*;��!;�;�;�;^��:���:���:&�:��:�Q�:36�:�I�:�s:��S:�5:o�:|��9�1�9�%t9_�8��07�ϸһY�K���:ݹgZ
���%��'A��?\��"w�jꈺT,���W���m���n��R]ʺ8׺:亦��{d��$���D�K��U������$�G*�Jk0�׊6���<���B�5�H��N�q�T�_[�a�g��m��$s��+y�G1�⛂� �������N���Ϫ��ȯ��������GŚ��  �  �f=�=�='B=�=�}==� =�T =o��<x�<�Q�<��<���<��<�%�<5X�<���<��<B��<C�<�C�<Ko�< ��<���<���<
�<�1�<�S�<Jt�<ʒ�<���<*��<���<���<��<T �<90�<�=�<I�<�Q�<�W�<�[�<^\�<YZ�<�U�<�M�<FC�<�5�<�$�<��<l��<���<���<���<�z�<�R�<�&�</��<��<*��<�R�<;�<��<%��<<B�<���<��<�M�<l��<E��<K6�<oѿ<�h�<L��<"��<�<l��<%�<��<�#�<c��<��<���<���<4c�<}̪<�2�<ӕ�<)��<fS�<��<��<1[�<��<Y��<pL�<C��<	�<�)�<�o�<���<���<�6�<�u�<γ�<S��<�+�<f�<Z��<�ׁ<��<��|<��x<gu<��q<	>n<P�j<<g<�c<\�_<�W\<-�X<�3U<@�Q<qN<��J<J�F<�sC<��?<�h<<��8<ri5<��1<w.<C+<4�'<'$<Y� <�[<W�<n�<�N<�<ô<5p	<1<a�<���;{1�;���;���;�s�;gO�;=9�;1�;�7�;FL�;6p�;��;��;M6�;���;��;���;*�;O��;Rd�;:#�;o�;Ѐ;.{w;�vm;��c;P�Y;W!P;��F;�*=;��3;��*;a�!;��;��;�;Z��:p��:n��:<�:f��:WR�:�5�:�J�:rs:�S:5:��:G��9�/�9�$t9��8�17��ϸ��Y�hI��Y>ݹ�Y
���%��)A�A\��"w��ꈺ�,��AW��Zn���m��]ʺ�7׺��ú�/c��!���D����������_$��F*�Ck0�K�6��<�<�B�X�H�^�N��T��[�a�g�m�6%s��+y��1����������������ת���������I����Ś��  �  �f=�=��=$B=�=�}==� =�T =k��<g�<�Q�<��<���< ��<�%�<?X�<���<��<8��<:�<�C�<5o�<$��<���<���<�<�1�<�S�<Mt�<ݒ�<���<3��<���<��<��<A �<D0�<�=�<"I�<�Q�<�W�<�[�<Y\�<eZ�<�U�<�M�<3C�<~5�<�$�<��<j��<���<���<���<�z�<�R�<�&�<3��<��<'��<�R�<;�<��<��<FB�<���<��<�M�<s��<P��<Q6�<�ѿ<�h�<W��<��<�<^��<
%�<��<�#�<w��<��< ��<���<8c�<�̪<�2�<ڕ�<��<kS�<��<��<([�<���<a��<qL�<V��<�<�)�<�o�<���<���<�6�<�u�<���<K��<�+�<f�<e��<�ׁ<��<��|<��x<&gu<��q<>n<"�j<@g<�c<i�_<�W\<6�X<�3U<F�Q<�N<v�J<^�F<vsC<��?<�h<<��8<�i5<��1<w.< +< �'<-'$<`� <\<V�<��<�N<��<��<"p	<+1<3�<���;�1�;���;���;�s�;�O�;I9�;M1�;�7�;iL�;/p�;Ѣ�;��;�5�;�;��;ц�;F�;q��;|d�;&#�;��;�π;w{w;2vm;Z�c;��Y;� P;��F;C*=;	�3;٪*;��!;��;�;�;��:8��:i��:A�:���:	Q�:/6�:8J�:�s:��S:�5:�:���9k4�9M#t9)�8�07��ϸw�Y��J���;ݹ0Z
���%�S)A�?\��"w��ꈺ�,��AW���m��3o��#]ʺ�7׺p�W��8d������D���V������$��G*�ak0��6���<���B���H�"�N�L�T�k[�pa��g��m��$s�]+y��1�ԛ���������d�������󯑻�����{Ś��  �  �f=�= �=B=�=�}==)� =�T =}��<��<�Q�<��<r��<��<�%�<=X�<���<$��<A��</�<�C�<3o�<3��<���<���<�<�1�<�S�<Bt�<ْ�<p��<9��<���<���<�<9 �<N0�<�=�<I�<�Q�<�W�<�[�<S\�<pZ�<�U�<�M�<@C�<�5�<�$�<��<���<���<��<���<�z�<�R�<�&�<9��<��<E��<�R�<B�<��<��<WB�<���<��<�M�<j��<J��<F6�<yѿ<�h�<_��<��<(�<h��<	%�<��<q#�<s��<��<���<���<<c�<�̪<�2�<땧<��<}S�<��<��<F[�<���<b��<aL�<N��<��<�)�<�o�<���<��<�6�<�u�<ó�<X��<�+�<�e�<v��<�ׁ<��<��|<��x<gu<��q<1>n<�j<zg<�c<s�_<�W\<�X<�3U<4�Q<�N<c�J<~�F<YsC<��?<�h<<��8<�i5<��1<1w.<T+<,�'<$'$<8� <\<1�<~�<�N<"�<��<p	<R1<0�<֊�;s1�;���;ڥ�;�s�;�O�;!9�;>1�;I7�;�L�;3p�;�;.�;�5�;薫;��;���;�;W��;[d�;#�;��;�π;�{w;�vm;Ðc;��Y; P;e�F;�*=;?�3;��*;R�!;��;��;;���:��:6��:��::�Q�:@7�:"I�:|s:z�S:�5:b�:���9v2�9+t9��8�h07ǫϸp�Y��J��{9ݹg\
���%��*A��?\�X$w�kꈺ�,���W���l�� o��\ʺ68׺�{���c�����xE�G�������T$��F*��j0�R�6��<���B�3�H���N���T�� [��a��g�;m�%s��+y��1�����5������u���������=�������Ś��  �  �f=�=��=$B=�=�}==� =�T =k��<g�<�Q�<��<���< ��<�%�<?X�<���<��<8��<:�<�C�<5o�<$��<���<���<�<�1�<�S�<Mt�<ݒ�<���<3��<���<��<��<A �<D0�<�=�<"I�<�Q�<�W�<�[�<Y\�<eZ�<�U�<�M�<3C�<~5�<�$�<��<j��<���<���<���<�z�<�R�<�&�<3��<��<'��<�R�<;�<��<��<FB�<���<��<�M�<s��<P��<Q6�<�ѿ<�h�<W��<��<�<^��<
%�<��<�#�<w��<��< ��<���<8c�<�̪<�2�<ڕ�<��<kS�<��<��<([�<���<a��<qL�<V��<�<�)�<�o�<���<���<�6�<�u�<���<K��<�+�<f�<e��<�ׁ<��<��|<��x<&gu<��q<>n<"�j<@g<�c<i�_<�W\<6�X<�3U<F�Q<�N<v�J<^�F<vsC<��?<�h<<��8<�i5<��1<w.< +< �'<-'$<`� <\<V�<��<�N<��<��<"p	<+1<3�<���;�1�;���;���;�s�;�O�;I9�;M1�;�7�;iL�;/p�;Ѣ�;��;�5�;�;��;ц�;F�;q��;|d�;&#�;��;�π;w{w;2vm;Z�c;��Y;� P;��F;C*=;	�3;٪*;��!;��;�;�;��:8��:i��:A�:���:	Q�:/6�:8J�:�s:��S:�5:�:���9k4�9M#t9)�8�07��ϸw�Y��J���;ݹ0Z
���%�S)A�?\��"w��ꈺ�,��AW���m��3o��#]ʺ�7׺p�W��8d������D���V������$��G*�ak0��6���<���B���H�"�N�L�T�k[�pa��g��m��$s�]+y��1�ԛ���������d�������󯑻�����{Ś��  �  �f=�=�='B=�=�}==� =�T =o��<x�<�Q�<��<���<��<�%�<5X�<���<��<B��<C�<�C�<Ko�< ��<���<���<
�<�1�<�S�<Jt�<ʒ�<���<*��<���<���<��<T �<90�<�=�<I�<�Q�<�W�<�[�<^\�<YZ�<�U�<�M�<FC�<�5�<�$�<��<l��<���<���<���<�z�<�R�<�&�</��<��<*��<�R�<;�<��<%��<<B�<���<��<�M�<l��<E��<K6�<oѿ<�h�<L��<"��<�<l��<%�<��<�#�<c��<��<���<���<4c�<}̪<�2�<ӕ�<)��<fS�<��<��<1[�<��<Y��<pL�<C��<	�<�)�<�o�<���<���<�6�<�u�<γ�<S��<�+�<f�<Z��<�ׁ<��<��|<��x<gu<��q<	>n<P�j<<g<�c<\�_<�W\<-�X<�3U<@�Q<qN<��J<J�F<�sC<��?<�h<<��8<ri5<��1<w.<C+<4�'<'$<Y� <�[<W�<n�<�N<�<ô<5p	<1<a�<���;{1�;���;���;�s�;gO�;=9�;1�;�7�;FL�;6p�;��;��;M6�;���;��;���;*�;O��;Rd�;:#�;o�;Ѐ;.{w;�vm;��c;P�Y;W!P;��F;�*=;��3;��*;a�!;��;��;�;Z��:p��:n��:<�:f��:WR�:�5�:�J�:rs:�S:5:��:G��9�/�9�$t9��8�17��ϸ��Y�hI��Y>ݹ�Y
���%��)A�A\��"w��ꈺ�,��AW��Zn���m��]ʺ�7׺��ú�/c��!���D����������_$��F*�Ck0�K�6��<�<�B�X�H�^�N��T��[�a�g�m�6%s��+y��1����������������ת���������I����Ś��  �  �f=�=��=#B=�=�}==� =�T =l��<w�<�Q�<��<���<��<�%�<7X�<���<��<:��<7�<�C�<<o�<+��<���<���<�<�1�<�S�<[t�<֒�<|��<8��<���<���<��<E �<B0�<�=�<I�<�Q�<X�<�[�<`\�<eZ�<�U�<�M�<AC�<�5�<�$�<��<n��<���<���<���<�z�<�R�<�&�<.��<��<-��<�R�<9�<��<��<FB�<���<��<�M�<p��<S��<\6�<wѿ<�h�<V��<��<�<d��<%�<��<�#�<n��<��<���<���<<c�<�̪<�2�<ߕ�<��<hS�<��<��<3[�<�<Y��<tL�<M��<�<�)�<�o�<���<���<�6�<�u�<³�<X��<�+�<	f�<g��<�ׁ<��<��|<��x<gu<��q<>n<0�j<@g<�c<a�_<�W\< �X<�3U<`�Q<mN<��J<a�F<qsC<��?<�h<<��8<�i5<��1<w.<@+<�'<''$<f� <\<`�<q�<�N<�<��<p	<$1<B�<���;~1�;��;���;�s�;xO�;�9�;11�;x7�;�L�;!p�;뢼;��;6�;���;�;���;`�;���;Yd�;A#�;��;�π;q{w;�vm;k�c;e�Y;� P;��F;�*=;��3;��*;��!;�;�;�;^��:���:���:&�:��:�Q�:36�:�I�:�s:��S:�5:o�:|��9�1�9�%t9_�8��07�ϸһY�K���:ݹgZ
���%��'A��?\��"w�jꈺT,���W���m���n��R]ʺ8׺:亦��{d��$���D�K��U������$�G*�Jk0�׊6���<���B�5�H��N�q�T�_[�a�g��m��$s��+y�G1�⛂� �������N���Ϫ��ȯ��������GŚ��  �  �f=�=��="B=�=�}==&� =�T =x��<s�<�Q�<��<~��<��<�%�<FX�<���<��<A��<9�<�C�<.o�<1��<���<���<�<�1�<�S�<Ht�<ؒ�<s��<6��<���<���<�<D �<E0�<�=�<I�<�Q�<�W�<�[�<S\�<kZ�<�U�<�M�<;C�<�5�<�$�<��<{��<���<��<���<�z�<�R�<�&�<<��<��<9��<�R�<C�<��<��<TB�<���<��<�M�<o��<I��<J6�<wѿ<�h�<Y��<��<�<i��<
%�<��<v#�<p��<��<���<���<1c�<�̪<�2�<镧<��<vS�<	��<��<;[�<�<k��<iL�<K��<�<�)�<�o�<���<���<�6�<�u�<���<V��<�+�<f�<j��<�ׁ<��<��|<��x<gu<��q<>n<+�j<Ug<�c<i�_<�W\<�X<�3U<=�Q<�N<r�J<c�F<msC<��?<�h<<��8<�i5<��1<'w.<8+<�'<:'$<O� <\<G�<��<�N<�<��<!p	<F1<%�<ϊ�;b1�;��;���;�s�;�O�;59�;71�;V7�;xL�;0p�;�;��;6�;Ė�;��;���;$�;Y��;id�;#�;��;�π;�{w;lvm;p�c;��Y;� P;�F;W*=;5�3;ɪ*;Y�!;��;��;%;��:X��:���:��:U��:BQ�:7�:HI�:�s:��S:r5:3�:���9�1�9�t9��8�07Y�ϸ��Y��J��;ݹ�[
�^�%�*A��?\�g#w�눺W,��X���l��so��|\ʺ�7׺��-��hd�����2E�^�����r���$�HG*��j0��6��<�ʾB�@�H�	�N���T�G[��a��g�m�%s��+y��1�ӛ��
���Z���V�������ꯑ�"���!����Ś��  �  �f=�=��='B=	�=�}== � =�T =t��<p�<�Q�<��<|��<��<�%�<;X�<���<��<>��<2�<�C�<>o�<(��<���<���<�<�1�<�S�<Et�<֒�<���<0��<���<���<��<J �<C0�<�=�<!I�<�Q�<�W�<�[�<U\�<kZ�<�U�<�M�<@C�<�5�<�$�<��<q��<���<��<���<�z�<�R�<�&�<7��<��<-��<�R�<5�<��<��<EB�<���<��<�M�<q��<K��<N6�<|ѿ<�h�<V��<��<�<d��<%�<��<�#�<o��<��<���<���<7c�<�̪<�2�<ޕ�<��<pS�< ��<��<0[�<���<a��<fL�<T��<�<�)�<�o�<���<���<�6�<�u�<ȳ�<V��<�+�<f�<k��<�ׁ<��<��|<��x<*gu<��q<>n<:�j<<g<�c<k�_<�W\<7�X<�3U<9�Q<�N<l�J<h�F<�sC<��?<�h<<��8<�i5<��1< w.<3+<1�'<"'$<L� <\<?�<z�<�N<��<��<p	<31<F�<���;G1�;��;���;�s�;�O�;+9�;/1�;�7�;`L�;.p�;뢼;��;%6�;���;��;ˆ�;7�;e��;ld�;#�;��;�π;F{w;�vm;��c;P�Y;� P;��F;p*=;$�3;��*;��!;�;��;�;c��:���:���:��:���:�Q�:6�:|I�:�s:l�S:�5:z�:���9E3�9d#t9x�8�07R�ϸ��Y�5J��K<ݹ�Y
�x�%��)A�t?\�##w��ꈺ�+��>X���m���n���\ʺa8׺�ں��c�����HE���������V$�CG*�k0���6���<�j�B�D�H���N�3�T�@[��a��g�m�%s�O+y��1�қ��힅�����=����������뵔�#����Ś��  �  �f=�=��=$B=�=�}== � =�T =q��<p�<�Q�<��<���<��<�%�<5X�<���<��<C��<=�<�C�<<o�<&��<���<���<�<�1�<�S�<Xt�<В�<}��</��<���<���<�<H �<=0�<�=�<I�<�Q�<X�<�[�<\\�<aZ�<�U�<�M�<@C�<�5�<�$�<��<i��<���<���<���<�z�<�R�<�&�<-��<��<&��<�R�<;�<��<��<FB�<���<��<�M�<m��<O��<X6�<qѿ<�h�<Q��<��<�<j��<%�<	��<�#�<g��<��<���<���<:c�<�̪<�2�<ܕ�<��<lS�<	��<��<*[�<���<W��<qL�<N��<�<�)�<�o�<���<���<�6�<�u�<ó�<T��<�+�<f�<e��<�ׁ<��<��|<��x<gu<��q<>n<6�j<Ng<�c<c�_<�W\<"�X<�3U<Y�Q<}N<z�J<^�F<vsC<��?<�h<<��8<�i5<��1<w.<3+<$�'<'$<e� <	\<X�<n�<�N<��<ƴ<)p	<,1<C�<���;�1�;���;���;�s�;�O�;v9�;1�;{7�;]L�;*p�;���;��;6�;���;��;���;O�;}��;Qd�;3#�;��;�π;h{w;�vm;��c;m�Y;L!P;�F;�*=;��3;�*;��!;̞;	�;�;���:$��:���:B�:Z��:�Q�:-6�:#J�:ms:�S:%5:�:x��9e0�9�"t9/	�8@�07v�ϸ̸Y�HJ���<ݹ�Z
���%��'A��?\�5#w��ꈺ�,��OW���m���n��]ʺ�7׺��<���c��.���D�F��R������$�1G*�Jk0�t�6��<���B�P�H�+�N�A�T�q[�Ka��g��m�%s��+y��1�䛂�����i���<���ʪ���������+���UŚ��  �  �f=�=��=B=�=�}==$� =�T =t��<z�<�Q�<��<���<��<�%�<:X�<���<��<C��<3�<�C�<4o�<.��<���<���<�<�1�<�S�<Gt�<ؒ�<z��<7��<���<���<
�<> �<H0�<�=�<I�<�Q�<�W�<�[�<^\�<cZ�<�U�<�M�<<C�<�5�<�$�<��<r��<���<���<���<�z�<�R�<�&�<1��<��<1��<�R�<8�<��<��<PB�<���<��<�M�<p��<H��<L6�<wѿ<�h�<\��<��< �<i��<%�<��<}#�<o��<��<���<���<:c�<|̪<�2�<啧<��<sS�<��<��<6[�<���<]��<sL�<G��<�<�)�<�o�<���<���<�6�<�u�<���<V��<�+�< f�<g��<�ׁ<��<��|<��x<gu<��q<>n<�j<cg<�c<g�_<�W\<%�X<�3U<<�Q<}N<��J<c�F<[sC<��?<�h<<��8<�i5<��1<w.<F+<�'<%'$<b� <�[<[�<y�<�N<�<Ŵ<p	<;1<1�<���;�1�;���;���;�s�;O�;29�;:1�;p7�;|L�;,p�;颼;��;�5�;Ζ�;��;���;&�;[��;dd�;;#�;��;�π;�{w;{vm;��c;{�Y;� P;͖F;�*=;��3;�*;f�!;��;�;�;���:ڦ�:���:�:���:pQ�:�6�:nI�:ys:Q�S:�5:�:M��92�9$!t9i�8ju07�ϸ:�Y�K���:ݹ�Z
�v�%��)A�M@\��"w��ꈺ�,���W��Am��!o���\ʺ>8׺��v���c������D����s������$��F*�#k0��6�G�<���B�D�H���N���T�^[�6a��g�m�!%s��+y��1�ӛ��*���>���t���ê��ᯑ����$����Ś��  �  �f=�=��=%B=�=�}=="� =�T =u��<k�<�Q�<��<���<��<�%�<;X�<���<��<@��<2�<�C�<4o�<-��<���<���<�<�1�<�S�<Ct�<ޒ�<x��<3��<���<���<�<A �<Q0�<�=�<&I�<�Q�<X�<�[�<P\�<oZ�<�U�<�M�<6C�<�5�<�$�<��<r��<���< ��<���<�z�<�R�<�&�<5��<���<-��<�R�<7�<��<��<NB�<���<#��<�M�<o��<V��<L6�<�ѿ<�h�<b��<��<�<a��<%�<��<z#�<x��<��<��<���<6c�<�̪<�2�<啧<��<rS�<���<��<-[�<���<_��<lL�<Q��<�<�)�<�o�<���<���<�6�<�u�<���<R��<�+�<	f�<m��<�ׁ<��<��|<��x<(gu<��q<5>n<#�j<Mg<�c<��_<�W\<.�X<�3U<>�Q<�N<c�J<j�F<xsC<��?<�h<<��8<�i5<��1<!w.<)+<-�'<$'$<Y� <\<L�<y�<�N<��<��<p	<71<2�<���;^1�;��;���;�s�;�O�;"9�;Q1�;i7�;kL�;Cp�;֢�;��;�5�;�;��;↠;)�;���;rd�;#�;��;�π;�{w;Jvm;~�c;l�Y;� P;ǖF;>*=;�3;̪*;��!;؞;��;�;��:���:���:��:h��:'Q�:�6�:AI�:4s:��S:`5:Ѣ:[��95�9�t9��8F�07��ϸ'�Y�WJ���:ݹH[
�k�%�9*A�>\��#w��ꈺ�+��X��<m��8o���\ʺl8׺���;d�����E�.��s�����c$�nG*�k0��6�e�<���B�c�H�)�N�q�T�+[��a�yg��m�
%s�T+y��1��������j���g������������������Ś��  �  �f=�=��=%B=�=�}==� =�T =v��<o�<�Q�<��<���<��<�%�<7X�<���<��<I��<?�<�C�<Co�<*��<���<���<�<�1�<�S�<Kt�<ђ�<}��<-��<���<���<�<K �<>0�<�=�<I�<�Q�<�W�<|[�<\\�<dZ�<�U�<�M�<CC�<�5�<�$�<��<p��<���<��<���<�z�<�R�<�&�<2��<��<,��<�R�<>�<��< ��<JB�<���<��<�M�<g��<M��<I6�<yѿ<�h�<R��<��<�<k��<%�<	��<#�<k��<��<���<���<<c�<�̪<�2�<���< ��<lS�<��<��<-[�<��<\��<nL�<G��<�<�)�<�o�<���<���<�6�<�u�<ʳ�<W��<�+�<f�<h��<�ׁ<��<��|<��x<'gu<��q<>n<>�j<Ig<�c<j�_<�W\<2�X<�3U<F�Q<vN<z�J<`�F<xsC<��?<�h<<��8<�i5<��1<#w.<1+<;�'<'$<[� <�[<R�<r�<�N<��<Ѵ<,p	<&1<P�<���;l1�;��;ĥ�;�s�;�O�;A9�;1�;~7�;TL�;8p�;���;��;&6�;���;��;���;�;m��;Bd�;3#�;��;�π;�{w;�vm;��c;v�Y;b!P;��F;�*=;�3;��*;_�!;��;��;�;��:���:���:u�:���:�Q�:g6�:�I�:�s:#�S:v5:��:���9a2�93 t9�
�8��07��ϸ��Y��I���<ݹ�Z
��%��)A��?\��#w�iꈺv,���W���m��]n��]ʺ�7׺:�	��Tc����
E����u�����B$�8G*�k0�V�6���<�V�B�:�H�'�N�J�T�U[�Oa�	g��m�E%s�\+y��1�ڛ��䞅�s���5��������������H���zŚ��  �  �f=�=��=#B=�=�}==� =�T =i��<v�<�Q�<��<���<��<�%�</X�<���<��<=��<1�<�C�<Ao�<��<���<���<�<�1�<�S�<\t�<Ғ�<���<5��<���<���<��<G �<?0�<�=�<I�<�Q�<X�<|[�<i\�<XZ�<�U�<�M�<;C�<�5�<�$�<��<f��<���<���<���<�z�<�R�<�&�<'��<��<#��<�R�<1�<��<��<>B�<���<��<�M�<l��<Q��<V6�<wѿ<�h�<S��<��<�<c��<%�<��<�#�<j��<��<�<���<>c�<|̪<�2�<ӕ�<��<kS�<���<��<+[�<���<S��<~L�<E��<�<�)�<�o�<���<���<�6�<�u�<ͳ�<N��<�+�<f�<_��<�ׁ<��<��|<��x<#gu<��q<>n<4�j<8g<�c<_�_<�W\<4�X<�3U<h�Q<\N<��J<S�F<psC<��?<�h<<��8<�i5<��1<	w.<@+<�'<'$<w� <�[<q�<c�<�N<��<��<p	<(1<K�<{��;�1�;���;���;�s�;[O�;�9�;1�;�7�;rL�; p�;㢼;��;6�;���;�;���;F�;���;Bd�;h#�;i�;�π;5{w;rvm;��c;"�Y;� P;h�F;�*=;��3;��*;��!;��;D�;;��:���:���:��:Z��:�Q�:�5�:�J�:/s:q�S:5:*�:���9�1�9�(t9��8۪07o�ϸ�Y�;K���;ݹOY
�"�%�{'A��@\�z"w�Tꈺ�,���V��Zn��~n��$]ʺ�8׺��1���c��O���D���� ������$��F*�}k0��6�Ȧ<�B�B���H�'�N�^�T��[��a�]g�sm�%s�k+y�Z1�雂���������P���Ҫ��ׯ��񵔻6���7Ś��  �  �f=�=��=%B=�=�}==%� =�T =z��<z�<�Q�<��<~��<��<�%�<:X�<���<��<I��<6�<�C�<8o�<(��<���<���<�<�1�<�S�<It�<Β�<r��<0��<���<���<�<H �<G0�<�=�<I�<�Q�< X�<[�<S\�<`Z�<�U�<�M�<>C�<�5�<�$�<��<x��<���<���<���<�z�<�R�<�&�<3��<��<6��<�R�<=�<��<��<HB�<���<��<�M�<h��<N��<F6�<rѿ<�h�<X��<��<"�<m��<%�<��<w#�<h��<��<���<���<-c�<�̪<�2�<ߕ�<��<wS�<��<��<7[�<���<^��<hL�<F��<�<�)�<�o�<���<���<�6�<�u�<ĳ�<U��<�+�<f�<a��<�ׁ<��<��|<��x<gu<��q<'>n<4�j<dg<�c<r�_<�W\<�X<3U<J�Q<zN<p�J<S�F<zsC<��?<�h<<��8<�i5<��1<,w.<F+<&�'<$'$<Q� <�[<D�<x�<�N<�<Ѵ<p	<C1<9�<���;1�;��;���;�s�;�O�;99�;1�;R7�;^L�;9p�; ��; �;6�;˖�;��;���;�;t��;Nd�;#�;��;�π;o{w;�vm;��c;��Y;� P;��F;�*=;�3;Ī*;C�!;��;��;�;���:$��:���:g�:���:�Q�:H6�:DJ�:gs:��S:�5:ء:��9�0�9�t9#�8��07��ϸ^�Y�]J���;ݹ�[
�[�%��)A�u?\��#w�b눺n,��mW���m���n��k\ʺ8׺n�n���c�����9E�����������$��F*��j0�Ɋ6�5�<���B�O�H�*�N�D�T��[��a��g��m�T%s��+y��1���������<���F����������5���J���sŚ��  �  �f=F=��=�A=��=D}=�=�� =7T =��<��<"P�<k��<���<-��<�#�<(V�<���<���<���<��<-A�<Xl�<?��<{��<q��<�
�<G.�<RP�<sp�<��<^��<���<y��<���<F	�<T�<:+�<�8�<�C�<KL�<KR�<�U�<CV�<;T�<9O�<gG�<�<�<�.�<��<�	�<,��<z��<���<
��<s�<�J�<��<%��<ֻ�<��<:J�<��<���<���<�9�<��<���<E�<���<͎�<�-�<ɿ<``�<��<ʃ�<��<K��<�<5��<��<ޕ�<i�<��<��<;\�<�Ū<,�<~��<��<gM�<'��<D �<�U�<˨�<p��<�G�<œ�<�ݖ<�%�<�k�<��<��<�3�<s�<*��<�<�)�<;d�<ٝ�<�ց<��<��|<��x<�fu<��q<>n<��j<�g<h�c<��_<�Z\<��X<�7U<��Q<wN<��J<AG<�yC<��?<Vp<<}�8<�q5<U�1<^�.<�+<f�'<�1$<g� <�g<M	< �<�[<I<��<1~	<�?<<���;�P�;@�;u��;���;�q�;�[�;^T�;[�;rp�;���;�Ǽ;�	�;H[�;w��;�,�;֬�;T<�;�ە;���;I�;��;���;�w;��m;�c;�Z;7jP;w�F;\r=;�#4;7�*;��!;��;3;;E;=�:&�:pB�:���:0�:�Ʃ:^��:۸�:L�s:|�T:"�5:bl:t�9.��9�w9�9��[7�uʸv0W����d	ܹ��	�!N%�!�@�h�[���v�������K ���6��w;��+ʺ	׺��㺏��:����k2��r���d��$�>9*��]0��~6�ښ<�޳B���H��N���T�b�Z��a�g��m��s�'y�l.�i���"�������,���Ȫ��q�������%���*ǚ��  �  �f=M=��=�A=��=?}=�=�� ==T =��<�<P�<Y��<ǻ�<7��<�#�<V�<~��<���<���<��<4A�<]l�<2��<���<e��<�
�<T.�<EP�<xp�<َ�<Z��<���<~��<���<G	�<^�<3+�<�8�<�C�<BL�<CR�<�U�<OV�<3T�<EO�<fG�<�<�<�.�<��<�	�</��<���<o��<��<#s�<�J�<��<��<��<��<IJ�<��<���<���<�9�<��<���<%E�<���<���<�-�<�ȿ<c`�< ��<Ӄ�<��<U��<�<0��<��<Ε�<m�<��<��<<\�<�Ū<,�<r��<��<oM�<5��<M �<�U�<Ψ�<_��<�G�<ѓ�<�ݖ<�%�<�k�<��<��<�3�< s�<2��<�<�)�<<d�<ӝ�<�ց<��<�|<��x<jfu<��q<u>n<�j<�g<|�c<��_<�Z\<u�X<c7U<��Q<UN<ӌJ<5G<�yC<��?<@p<<��8<�q5<j�1<[�.<�+<M�'<�1$<�� <�g<i	<ܯ<�[<U<��<M~	<�?<$<[��;�P�;�;f��;*��;{q�;�[�;#T�;�Z�;ap�;���;�Ǽ;�	�;o[�;\��;�,�;���;2<�;}ە;���;GI�;��;���;�w;��m;^�c;�Z;�jP;��F;�r=;�"4;�*;�!;,�;A;�D;�=�:C&�:aC�:<��:��:�Ʃ:�:ù�:5�s:��T:h�5:�j:s�9(��9gw9��9�1\7�rʸ�+W�2���
ܹ��	�)P%���@��[�ޣv�������P��O7��;;���*ʺ'׺���B��c:�����2�ar�Y������$��8*��]0�-~6���<���B�#�H���N���T���Z�Fa��g�om�I s��'y�V.�~���	���ϡ�����Ϫ��t����]���ǚ��  �  �f=T=��=�A=��=:}=�=�� =>T =��<�<P�<Z��<ͻ�<&��<�#�<V�<���<���<���<��<(A�<dl�<'��<���<^��<�
�<^.�<<P�<�p�<َ�<h��<���<v��<���<>	�<c�<)+�<�8�<�C�<OL�<NR�<�U�<ZV�<&T�<JO�<aG�<�<�<�.�<��<�	�< ��<���<q��<��<!s�<�J�<��<��<��<���<BJ�<��<���<���<�9�<��<}��</E�<���<Ȏ�<�-�< ɿ<o`�<��<Ճ�<��<Q��<�<+��<��<͕�<}�<��<��<A\�<�Ū<#,�<h��<��<dM�<+��<D �<�U�<֨�<]��<�G�<���<�ݖ<�%�<�k�<!��<��<�3�<s�<4��<��<�)�<:d�<˝�<�ց<��<�|<��x<zfu<��q<a>n<�j<�g<��c<��_<�Z\<��X<f7U<��Q<=N<�J<+G<�yC<��?<.p<<��8<�q5<m�1<?�.<�+<Y�'<�1$<�� <|g<u	<ܯ<�[<M<u�<A~	<�?<2<.��;�P�;��;g��;S��;Xq�;\�;$T�;)[�;\p�;���;�Ǽ;�	�;�[�;3��;�,�;���;c<�;�ە;z��;rI�;z�;���;��w;��m;:�c;XZ;~jP;�F;�r=;�"4;W�*;��!;��;�;�D;3>�:]%�:�B�::��:4�:�Ʃ:x��:W��:��s:��T:��5:�k:�v�9���9�
w9N�9�;\7d{ʸZ-W�Y��ܹ�	�6P%���@�}�[���v�=���.�y���7���:��C+ʺ�׺���ŏ��9������1��r�E�����t$��8*�<^0�%~6��<���B�[�H���N���T���Z��a��g��m�2 s�T'y�.�����񝅻案���������S�������Y����ƚ��  �  �f=L=��=�A=��=<}=�=�� =AT =��<��< P�<_��<»�<)��<�#�<V�<���<���<���<��<)A�<fl�<.��<���<h��<�
�<N.�<CP�<zp�<׎�<`��<���<z��<���<C	�<d�<1+�<�8�<�C�<AL�<HR�<�U�<OV�<3T�<CO�<eG�<�<�<�.�<��<�	�<-��<��<|��<
��<s�<�J�<��<��<ݻ�<��<JJ�<��<���<���<�9�<��<���<%E�<���<Ď�<�-�< ɿ<e`�<��<փ�<��<Q��<�<-��<��<Ε�<n�<��<��<=\�<�Ū<,�<p��<��<fM�<1��<O �<�U�<Ϩ�<h��<�G�<Ó�<�ݖ<�%�<�k�<��<��<�3�<s�<6��< �<�)�<:d�<ӝ�<�ց<��<�|<��x<{fu<��q<n>n<�j<�g<��c<��_<�Z\<��X<X7U<��Q<PN<όJ<7G<�yC<��?<8p<<��8<�q5<|�1<[�.<�+<a�'<�1$<}� <�g<_	<�<�[<H<��<M~	<�?<6<J��;�P�;�;l��;��;uq�;�[�;T�;[�;Xp�;���;�Ǽ;�	�;�[�;T��;�,�;���;,<�;�ە;t��;EI�;��;���;�w;��m;U�c;�Z;�jP;{�F;�r=;Z#4;7�*;��!;��;[;E;x=�:&�:gC�:���:b�:ǩ:騙:ǹ�:0�s:��T:��5:]k:�r�9���9�w97�9�G\7�vʸ�-W�����ܹ%�	�P%���@�ڻ[�|�v�|�����V��q7���:��!+ʺh׺��㺝��L:��G��/2��r�������1$�9*��]0��}6��<���B�>�H���N���T���Z�Pa��g�Qm�q s�R'y�^.�����񝅻ʡ������䪎�t���ɶ��s����ƚ��  �  �f=H=��=�A=��=?}=�=�� =6T =!��<��<P�<[��<���<C��<�#�<V�<x��<���<���<��<.A�<[l�<8��<���<i��<�
�<L.�<TP�<up�<��<Y��<���<|��<���<D	�<V�<:+�<�8�<�C�<@L�<JR�<�U�<HV�<;T�<<O�<lG�<�<�<�.�<��<�	�<7��<|��<z��<���<$s�<�J�<��<��<ػ�<��<<J�<��<���<���<�9�<��<���<E�<���<ʎ�<�-�<ɿ<^`�<��<̃�<��<N��<�<2��<��<ە�<j�<��<��<:\�<�Ū<,�<z��<��<iM�<*��<G �<�U�<ƨ�<h��<�G�<ړ�<�ݖ<�%�<�k�<��<��<�3�<s�<2��<�<�)�<6d�<؝�<�ց<��<�|<��x<yfu<��q<�>n<��j<�g<i�c<��_<�Z\<��X<o7U<��Q<pN<��J<;G<�yC<��?<Cp<<��8<�q5<Q�1<c�.<�+<R�'<�1$<x� <�g<V	<�<{[<R<��<8~	<�?<!<s��;�P�;�;g��;��;�q�;�[�;RT�;�Z�;bp�;���;�Ǽ;�	�;Q[�;y��;�,�;Ȭ�;+<�;�ە;���;)I�;��;���;C�w;��m;H�c;�Z;0jP;��F;jr=;H#4;��*;�!;Q�;;
E;"=�:�&�:�B�:���:n�:�Ʃ:s��:K��:B�s:��T:�5:l:Lr�9\��9�w9��9��[7�vʸ�.W����D
ܹ*�	��N%���@�"�[�I�v�����B񕺡���6��d;���*ʺ�׺d��8���:��H��X2�r�������e$�9*��]0��~6�Ú<���B�%�H���N���T�k�Z��a�.g�jm�< s�X'y�z.�^���/���ϡ��)�������}���ض��F���ǚ��  �  �f=M=��=�A=��==}=�=�� =:T =��<�<P�<d��<���<+��<�#�<"V�<���<���<���<��<2A�<^l�<0��<���<a��<�
�<R.�<@P�<tp�<ߎ�<a��<���<t��<���<F	�<X�<3+�<�8�<�C�<FL�<BR�<�U�<NV�<2T�<@O�<jG�<�<�<�.�<��<�	�<1��<���<y��<��<s�<�J�<��<��<��<��<AJ�<��<���<���<�9�<��<���<#E�<���<���<�-�<ɿ<e`�<��<̃�<��<N��<
�<2��<��<֕�<k�<��<��<?\�<�Ū<,�<q��<��<lM�<.��<G �<�U�<Ϩ�<i��<�G�<Ó�<�ݖ<�%�<�k�<��<��<�3�<s�</��<�<�)�<6d�<՝�<�ց<��<�|<��x<xfu<��q<y>n<��j<�g<m�c<��_<�Z\<��X<p7U<��Q<JN<ӌJ<:G<�yC<��?<;p<<��8<�q5<_�1<^�.<�+<\�'<�1$<s� <�g<S	<��<�[<^<��<@~	<�?<&<S��;�P�;��;{��;#��;fq�;�[�;=T�;[�;sp�;}��;�Ǽ;�	�;X[�;\��;�,�;���;?<�;|ە;{��;CI�;��;���;.�w;��m;N�c;�Z;ajP;��F;�r=;@#4;*�*;��!;��;2;�D;�=�:K&�:�B�:ޒ�:��:�Ʃ:'��:���:��s:p�T:q�5:�j:�s�9$��9�w9��9��[7�uʸ�.W�	��>
ܹ	�	�%O%��@���[��v�V�������U7��;���*ʺ�׺d����D:��:��[2��r�������X$��8*��]0�f~6���<���B�5�H���N���T���Z�Ka��g�~m�' s�['y�3.�v����������"���ݪ��\���϶��E���ǚ��  �  �f=N=��=�A=��==}=�=�� =?T =��<��<P�<`��<Ļ�<3��<�#�<V�<}��<���<���<��<(A�<il�<*��<���<a��<�
�<S.�<BP�<�p�<֎�<]��<���<|��<���<B	�<f�</+�<�8�<�C�<KL�<FR�<�U�<VV�<,T�<HO�<`G�<�<�<�.�<��<�	�<(��<���<t��<��<s�<�J�<��<��<��<��<JJ�<��<���<���<�9�<��<���<*E�<���<�<�-�<�ȿ<h`�<��<ڃ�<��<P��<�<,��<��<˕�<z�<��<��<@\�<�Ū<,�<j��<��<cM�<1��<K �<�U�<ͨ�<f��<�G�<˓�<�ݖ<�%�<�k�<��<��<�3�<s�<4��<�<�)�<;d�<͝�<�ց<��<��|<��x<jfu<��q<q>n<�j<�g<�c<��_<�Z\<w�X<a7U<��Q<LN<،J<0G<�yC<��?<;p<<��8<�q5<t�1<R�.<�+<V�'<�1$<�� <�g<e	<�<�[<J<��<L~	<�?<<<:��;�P�; �;u��;(��;nq�;�[�;T�;�Z�;\p�;���;�Ǽ;�	�;�[�;L��;�,�;���;S<�;�ە;y��;bI�;��;���;��w;��m;E�c;�Z;�jP;T�F;�r=;#4;K�*;��!;
�;z;�D;�=�:�%�:rC�:���:6�:=ǩ:���:	��:�s:M�T:>�5:k:�u�9ޭ�9_w9��9�g\7Fwʸ.W����ܹ1�	�}P%��@� �[�ѣv�I���������7��n:��Q+ʺi׺#�㺤��k:��Y��2��r�v�����d$��8*��]0��}6��<���B��H���N���T���Z�$a��g�7m�@ s��'y�H.���������ա������۪��m���궔�a����ƚ��  �  �f=I=��=�A=��=?}=�=�� =9T = ��<�<P�<]��<���<=��<�#�<#V�<��<���<���<��<&A�<bl�<1��<���<j��<�
�<P.�<JP�<vp�<ߎ�<a��<���<|��<���<:	�<[�<3+�<�8�<�C�<EL�<FR�<�U�<LV�<4T�<BO�<bG�<�<�<�.�<��<�	�<2��<���<{��<��<s�<�J�<��<��<ݻ�<���<>J�<��<���<���<�9�<��<���<"E�<���<Ǝ�<�-�<ɿ<i`�<��<Ѓ�<��<L��<�<0��<��<ԕ�<m�<��<��<=\�<�Ū<,�<p��<��<cM�<,��<H �<�U�<̨�<j��<�G�<ѓ�<�ݖ<�%�<�k�<��<��<�3�<s�<3��<�<�)�<<d�<ӝ�<�ց<��<�|<��x<~fu<��q<y>n<�j<�g<q�c<��_<�Z\<��X<i7U<��Q<dN<ŌJ<4G<�yC<��?<Bp<<��8<�q5<\�1<b�.<�+<`�'<�1$<p� <�g<O	<��<�[<Y<��<=~	<�?</<W��;�P�;"�;h��;��;�q�;�[�;=T�;[�;dp�;���;�Ǽ;�	�;d[�;Z��;�,�;���;=<�;�ە;���;:I�;��;���;��w;��m;D�c;mZ;PjP;��F;�r=;O#4;�*;��!;�;;E;�=�:e&�:�B�:l��:R�:�Ʃ:Ҩ�:���:��s:M�T:��5:�k:�s�9ϯ�9�w9��9�\7�}ʸ�/W�����
ܹ��	�gO%���@�>�[��v�����]�G��d7���:��K+ʺ�׺W����:��3��m2�`r�������8$��8*��]0�t~6���<���B��H���N���T���Z�ta�Og�sm�G s�C'y�'.�u�������������̪��a���Ŷ��R���ǚ��  �  �f=J=��=�A=��=?}=�=�� =;T =!��< �<P�<f��<���<5��<�#�<)V�<v��<���<���<��<6A�<Zl�<6��<���<g��<�
�<R.�<FP�<np�<��<X��<���<r��<���<P	�<[�<2+�<�8�<�C�<DL�<AR�<�U�<GV�<<T�<:O�<mG�<�<�<�.�<��<�	�<7��<z��<|��<��<s�<�J�<��<#��<ջ�<���<:J�<��<���<���<�9�<��<���<E�<���<���<�-�<ɿ<_`�<��<̃�<��<U��<�<0��<��<ە�<g�<��<��<<\�<�Ū<,�<y��<��<nM�<1��<C �<�U�<Ũ�<q��<�G�<͓�<�ݖ<�%�<�k�<��<��<�3�<)s�<,��<�<�)�<2d�<ڝ�<�ց<��<�|<��x<pfu<��q<m>n<�j<�g<u�c<��_<�Z\<y�X<n7U<��Q<[N<ɌJ<@G<�yC<��?<Ap<<�8<�q5<b�1<d�.<�+<Q�'<�1$<p� <�g<E	<�<x[<\<��<C~	<�?<<m��;�P�;�;k��;$��;�q�;�[�;OT�;�Z�;ap�;v��;�Ǽ;"
�;c[�;X��;�,�;���;9<�;yە;���;&I�;��;���;H�w;��m;8�c;�Z;BjP;��F;ar=;Y#4;�*;��!;
�; ;'E;=�:�&�:lB�:5��:{�:�Ʃ:���:B��:9�s:��T:��5:�j:�r�9���9�w9��9�[7?mʸ�+W�����
ܹ�	��N%�s�@���[�أv�����R񕺆���6��`;���*ʺ_׺������:������2�}r�������h$�
9*��]0�`~6�R�<�ͳB�(�H���N���T�[�Z��a�ug��m�- s�{'y�k.�����������������y���趔�G���(ǚ��  �  �f=N=��=�A=��=>}=�=�� ==T =��<�<P�<^��<Ż�<6��<�#�<V�<z��<���<���<��<(A�<bl�</��<���<a��<�
�<U.�<CP�<�p�<ێ�<Z��<���<y��<���<:	�<a�<2+�<�8�<�C�<ML�<FR�<�U�<RV�<2T�<@O�<gG�<�<�<�.�<��<�	�<+��<���<v��<	��<s�<�J�<��<��<ݻ�<��<=J�<��<���<���<�9�<��<���<'E�<���<�<�-�<�ȿ<f`�<��<փ�<��<M��<�<4��<��<Е�<y�<��<��<>\�<�Ū<,�<q��<��<bM�<1��<B �<�U�<ʨ�<g��<�G�<͓�<�ݖ<�%�<�k�<��<��<�3�<s�<0��<�<�)�<3d�<ѝ�<�ց<��<��|<��x<hfu<��q<r>n<�j<�g<|�c<��_<�Z\<v�X<k7U<��Q<PN<،J<1G<�yC<��?<=p<<��8<�q5<j�1<K�.<�+<S�'<�1$<�� <�g<f	<�<�[<Y<w�<G~	<�?</<P��;�P�; �;c��;0��;rq�;�[�;,T�;�Z�;zp�;���;�Ǽ;�	�;y[�;X��;�,�;���;_<�;�ە;���;OI�;��;���;�w;��m;�c;�Z;_jP;l�F;�r=;(#4;,�*;��!;�;[;�D;}=�:&�:�B�:���:�:�Ʃ:��:���:�s:��T:��5:k:�u�9���9)w9��9]D\7�|ʸ�/W�����	ܹ��	��O%�,�@��[���v�r�������_7���:��b+ʺj׺���S��:��L��2�~r�v�����n$��8*��]0�?~6�ۚ<���B�'�H���N���T���Z�.a��g�*m� s��'y� .���������������ݪ��W�����M����ƚ��  �  �f=M=��=�A=��=;}=�=�� =ET =��<	�<P�<Z��<ƻ�</��<�#�<V�<���<���<���<��<"A�<ol�<&��<���<d��<�
�<R.�<>P�<~p�<͎�<h��<���<x��<���<8	�<g�<&+�<�8�<�C�<DL�<AR�<�U�<PV�<)T�<MO�<\G�<�<�<�.�<��<�	�<*��<���<s��<��<s�<�J�<��<��<��<��<NJ�<��<���<���<�9�< ��<���<%E�<���<���<�-�<�ȿ<p`�<��<ڃ�<��<T��<�<)��<��<Õ�<r�<��<��<;\�<�Ū<,�<e��<��<aM�<9��<N �<�U�<ը�<_��<�G�<Ǔ�<�ݖ<�%�<�k�<!��<��<�3�<s�<@��< �<�)�<Bd�<ʝ�<�ց<��<��|<��x<sfu<��q<a>n<%�j<�g<��c<��_<�Z\<��X<O7U<��Q<LN<ӌJ<&G<�yC<��?<3p<<��8<�q5<��1<W�.<�+<`�'<�1$<�� <�g<e	<ܯ<�[<Y<��<_~	<�?<I<-��;�P�;�;Y��;%��;_q�;�[�;�S�;)[�;Rp�;���;�Ǽ;�	�;�[�;)��;�,�;���;8<�;wە;|��;JI�;��;���;��w;��m;��c;{Z;�jP;f�F;�r=;#4; �*;��!;��;K;�D;!>�:�%�:�C�:В�:��:�ǩ:D��:b��:�s:��T:,�5:oj:�s�9C��9Jw9��9j\7�|ʸ,W����ܹ��	�~Q%���@�ż[��v������񕺵��!8��-:��k+ʺ�׺���H���9�����2��r�m�����\$��8*��]0��}6��<�/�B�=�H���N�~�T���Z�?a��g�[m�� s�p'y�.�����ϝ�����٥������_���Ƕ�������ƚ��  �  �f=K=��=�A=��=>}=�=�� =;T =��<��<P�<d��<Ļ�<6��<�#�< V�<{��<���<���<��<*A�<cl�<0��<���<a��<�
�<R.�<LP�<~p�<܎�<a��<���<t��<���<H	�<c�<)+�<�8�<�C�<LL�<LR�<�U�<KV�<3T�<@O�<fG�<�<�<�.�<��<�	�<+��<}��<y��<
��<#s�<�J�<��<��<ڻ�<��<>J�<��<���<���<�9�<��<���<"E�<���<̎�<�-�<ɿ<i`�<��<Ӄ�<��<U��<�<%��<��<ҕ�<w�<��<��<>\�<�Ū<,�<q��<��<fM�<,��<D �<�U�<ɨ�<i��<�G�<ϓ�<�ݖ<�%�<�k�<��<��<�3�<s�<4��<�<�)�<5d�<՝�<�ց<��<��|<��x<vfu<��q<`>n<�j<�g<��c<��_<�Z\<��X<i7U<��Q<eN<ʌJ<;G<�yC<��?<=p<<��8<�q5<e�1<U�.<�+<S�'<�1$<�� <�g<X	<�<�[<J<�<?~	<�?<1<S��;�P�; �;n��;$��;�q�;�[�;3T�;[�;<p�;~��;�Ǽ;
�;�[�;4��;�,�;���;Z<�;�ە;���;4I�;��;���;�w;��m;@�c;Z;VjP;i�F;yr=;A#4;:�*;�!;0�;N; E;P=�:�%�:�B�:~��:G�:�Ʃ:�:���:�s:P�T:B�5:Gl:�u�9���9�w9�92\7�rʸ]+W�����ܹ��	��O%�o�@���[���v�i��������\7���:��'+ʺ�׺��㺗��:��>��H2�pr�d�����g$�
9*��]0�K~6�˚<���B�/�H���N���T���Z�{a�Fg�?m�& s�e'y�J.�����ꝅ�ʡ��󥋻����z���ж��R����ƚ��  �  �f=G=��=�A=��=@}=�=�� =7T =(��<�<P�<d��<���<9��<�#�<'V�<x��<Ƿ�<���<��<8A�<Vl�<6��<���<^��<�
�<J.�<DP�<op�<܎�<T��<���<���<���<;	�<Y�<:+�<�8�<�C�<AL�<?R�<�U�<HV�<?T�<0O�<rG�<�<�<�.�<��<�	�<;��<��<~��<��<s�<�J�<��<"��<ػ�<���<@J�<��<���<���<�9�<��<���<!E�<���<���<�-�<�ȿ<_`�<��<σ�<��<H��<�<8��<��<ϕ�<g�<��<��<A\�<�Ū<,�<y��<��<oM�<1��<O �<�U�<Ũ�<p��<�G�<ϓ�<�ݖ<�%�<�k�<��<��<�3�<(s�<'��<�<�)�<'d�<㝃<�ց<��<݋|<��x<gfu<��q<�>n<��j<�g<f�c<��_<�Z\<p�X<k7U<��Q<WN<��J<RG<�yC<��?<Fp<<u�8<�q5<S�1<q�.<�+<W�'<�1$<j� <�g<M	<��<{[<j<��<;~	<�?<<m��;�P�;��;���;��;vq�;�[�;2T�;�Z�;�p�;���;�Ǽ;�	�;][�;x��;�,�;���;-<�;pە;���;*I�;��;���;m�w;��m;+�c;�Z;JjP;��F;�r=;i#4;��*;��!;�;;!E;.=�:�&�:�B�:I��:w�:~Ʃ:���:ø�:2�s:/�T:Z�5:�j:Mr�9���9�w9��9f\7�|ʸ�1W�����ܹb�	��O%�q�@��[���v�:����񕺓���6���;���*ʺf׺��㺦���:�� ���2�or�ͬ����F$��8*�t]0��~6�U�<���B��H�g�N�T�T��Z��a�yg��m�4 s��'y�.�[���"����0�������S�������M���)ǚ��  �  �f=K=��=�A=��=>}=�=�� =;T =��<��<P�<d��<Ļ�<6��<�#�< V�<{��<���<���<��<*A�<cl�<0��<���<a��<�
�<R.�<LP�<~p�<܎�<a��<���<t��<���<H	�<c�<)+�<�8�<�C�<LL�<LR�<�U�<KV�<3T�<@O�<fG�<�<�<�.�<��<�	�<+��<}��<y��<
��<#s�<�J�<��<��<ڻ�<��<>J�<��<���<���<�9�<��<���<"E�<���<̎�<�-�<ɿ<i`�<��<Ӄ�<��<U��<�<%��<��<ҕ�<w�<��<��<>\�<�Ū<,�<q��<��<fM�<,��<D �<�U�<ɨ�<i��<�G�<ϓ�<�ݖ<�%�<�k�<��<��<�3�<s�<4��<�<�)�<5d�<՝�<�ց<��<��|<��x<vfu<��q<`>n<�j<�g<��c<��_<�Z\<��X<i7U<��Q<eN<ʌJ<;G<�yC<��?<=p<<��8<�q5<e�1<U�.<�+<S�'<�1$<�� <�g<X	<�<�[<J<�<?~	<�?<1<S��;�P�; �;n��;$��;�q�;�[�;3T�;[�;<p�;~��;�Ǽ;
�;�[�;4��;�,�;���;Z<�;�ە;���;4I�;��;���;�w;��m;@�c;Z;VjP;i�F;yr=;A#4;:�*;�!;0�;N; E;P=�:�%�:�B�:~��:G�:�Ʃ:�:���:�s:P�T:B�5:Gl:�u�9���9�w9�92\7�rʸ]+W�����ܹ��	��O%�o�@���[���v�i��������\7���:��'+ʺ�׺��㺗��:��>��H2�pr�d�����g$�
9*��]0�K~6�˚<���B�/�H���N���T���Z�{a�Fg�?m�& s�e'y�J.�����ꝅ�ʡ��󥋻����z���ж��R����ƚ��  �  �f=M=��=�A=��=;}=�=�� =ET =��<	�<P�<Z��<ƻ�</��<�#�<V�<���<���<���<��<"A�<ol�<&��<���<d��<�
�<R.�<>P�<~p�<͎�<h��<���<x��<���<8	�<g�<&+�<�8�<�C�<DL�<AR�<�U�<PV�<)T�<MO�<\G�<�<�<�.�<��<�	�<*��<���<s��<��<s�<�J�<��<��<��<��<NJ�<��<���<���<�9�< ��<���<%E�<���<���<�-�<�ȿ<p`�<��<ڃ�<��<T��<�<)��<��<Õ�<r�<��<��<;\�<�Ū<,�<e��<��<aM�<9��<N �<�U�<ը�<_��<�G�<Ǔ�<�ݖ<�%�<�k�<!��<��<�3�<s�<@��< �<�)�<Bd�<ʝ�<�ց<��<��|<��x<sfu<��q<a>n<%�j<�g<��c<��_<�Z\<��X<O7U<��Q<LN<ӌJ<&G<�yC<��?<3p<<��8<�q5<��1<W�.<�+<`�'<�1$<�� <�g<e	<ܯ<�[<Y<��<_~	<�?<I<-��;�P�;�;Y��;%��;_q�;�[�;�S�;)[�;Rp�;���;�Ǽ;�	�;�[�;)��;�,�;���;8<�;wە;|��;JI�;��;���;��w;��m;��c;{Z;�jP;f�F;�r=;#4; �*;��!;��;K;�D;!>�:�%�:�C�:В�:��:�ǩ:D��:b��:�s:��T:,�5:oj:�s�9C��9Jw9��9j\7�|ʸ,W����ܹ��	�~Q%���@�ż[��v������񕺵��!8��-:��k+ʺ�׺���H���9�����2��r�m�����\$��8*��]0��}6��<�/�B�=�H���N�~�T���Z�?a��g�[m�� s�p'y�.�����ϝ�����٥������_���Ƕ�������ƚ��  �  �f=N=��=�A=��=>}=�=�� ==T =��<�<P�<^��<Ż�<6��<�#�<V�<z��<���<���<��<(A�<bl�</��<���<a��<�
�<U.�<CP�<�p�<ێ�<Z��<���<y��<���<:	�<a�<2+�<�8�<�C�<ML�<FR�<�U�<RV�<2T�<@O�<gG�<�<�<�.�<��<�	�<+��<���<v��<	��<s�<�J�<��<��<ݻ�<��<=J�<��<���<���<�9�<��<���<'E�<���<�<�-�<�ȿ<f`�<��<փ�<��<M��<�<4��<��<Е�<y�<��<��<>\�<�Ū<,�<q��<��<bM�<1��<B �<�U�<ʨ�<g��<�G�<͓�<�ݖ<�%�<�k�<��<��<�3�<s�<0��<�<�)�<3d�<ѝ�<�ց<��<��|<��x<hfu<��q<r>n<�j<�g<|�c<��_<�Z\<v�X<k7U<��Q<PN<،J<1G<�yC<��?<=p<<��8<�q5<j�1<K�.<�+<S�'<�1$<�� <�g<f	<�<�[<Y<w�<G~	<�?</<P��;�P�; �;c��;0��;rq�;�[�;,T�;�Z�;zp�;���;�Ǽ;�	�;y[�;X��;�,�;���;_<�;�ە;���;OI�;��;���;�w;��m;�c;�Z;_jP;l�F;�r=;(#4;,�*;��!;�;[;�D;}=�:&�:�B�:���:�:�Ʃ:��:���:�s:��T:��5:k:�u�9���9)w9��9]D\7�|ʸ�/W�����	ܹ��	��O%�,�@��[���v�r�������_7���:��b+ʺj׺���S��:��L��2�~r�v�����n$��8*��]0�?~6�ۚ<���B�'�H���N���T���Z�.a��g�*m� s��'y� .���������������ݪ��W�����M����ƚ��  �  �f=J=��=�A=��=?}=�=�� =;T =!��< �<P�<f��<���<5��<�#�<)V�<v��<���<���<��<6A�<Zl�<6��<���<g��<�
�<R.�<FP�<np�<��<X��<���<r��<���<P	�<[�<2+�<�8�<�C�<DL�<AR�<�U�<GV�<<T�<:O�<mG�<�<�<�.�<��<�	�<7��<z��<|��<��<s�<�J�<��<#��<ջ�<���<:J�<��<���<���<�9�<��<���<E�<���<���<�-�<ɿ<_`�<��<̃�<��<U��<�<0��<��<ە�<g�<��<��<<\�<�Ū<,�<y��<��<nM�<1��<C �<�U�<Ũ�<q��<�G�<͓�<�ݖ<�%�<�k�<��<��<�3�<)s�<,��<�<�)�<2d�<ڝ�<�ց<��<�|<��x<pfu<��q<m>n<�j<�g<u�c<��_<�Z\<y�X<n7U<��Q<[N<ɌJ<@G<�yC<��?<Ap<<�8<�q5<b�1<d�.<�+<Q�'<�1$<p� <�g<E	<�<x[<\<��<C~	<�?<<m��;�P�;�;k��;$��;�q�;�[�;OT�;�Z�;ap�;v��;�Ǽ;"
�;c[�;X��;�,�;���;9<�;yە;���;&I�;��;���;H�w;��m;8�c;�Z;BjP;��F;ar=;Y#4;�*;��!;
�; ;'E;=�:�&�:lB�:5��:{�:�Ʃ:���:B��:9�s:��T:��5:�j:�r�9���9�w9��9�[7?mʸ�+W�����
ܹ�	��N%�s�@���[�أv�����R񕺆���6��`;���*ʺ_׺������:������2�}r�������h$�
9*��]0�`~6�R�<�ͳB�(�H���N���T�[�Z��a�ug��m�- s�{'y�k.�����������������y���趔�G���(ǚ��  �  �f=I=��=�A=��=?}=�=�� =9T = ��<�<P�<]��<���<=��<�#�<#V�<��<���<���<��<&A�<bl�<1��<���<j��<�
�<P.�<JP�<vp�<ߎ�<a��<���<|��<���<:	�<[�<3+�<�8�<�C�<EL�<FR�<�U�<LV�<4T�<BO�<bG�<�<�<�.�<��<�	�<2��<���<{��<��<s�<�J�<��<��<ݻ�<���<>J�<��<���<���<�9�<��<���<"E�<���<Ǝ�<�-�<ɿ<i`�<��<Ѓ�<��<L��<�<0��<��<ԕ�<m�<��<��<=\�<�Ū<,�<p��<��<cM�<,��<H �<�U�<̨�<j��<�G�<ѓ�<�ݖ<�%�<�k�<��<��<�3�<s�<3��<�<�)�<<d�<ӝ�<�ց<��<�|<��x<~fu<��q<y>n<�j<�g<q�c<��_<�Z\<��X<i7U<��Q<dN<ŌJ<4G<�yC<��?<Bp<<��8<�q5<\�1<b�.<�+<`�'<�1$<p� <�g<O	<��<�[<Y<��<=~	<�?</<W��;�P�;"�;h��;��;�q�;�[�;=T�;[�;dp�;���;�Ǽ;�	�;d[�;Z��;�,�;���;=<�;�ە;���;:I�;��;���;��w;��m;D�c;mZ;PjP;��F;�r=;O#4;�*;��!;�;;E;�=�:e&�:�B�:l��:R�:�Ʃ:Ҩ�:���:��s:M�T:��5:�k:�s�9ϯ�9�w9��9�\7�}ʸ�/W�����
ܹ��	�gO%���@�>�[��v�����]�G��d7���:��K+ʺ�׺W����:��3��m2�`r�������8$��8*��]0�t~6���<���B��H���N���T���Z�ta�Og�sm�G s�C'y�'.�u�������������̪��a���Ŷ��R���ǚ��  �  �f=N=��=�A=��==}=�=�� =?T =��<��<P�<`��<Ļ�<3��<�#�<V�<}��<���<���<��<(A�<il�<*��<���<a��<�
�<S.�<BP�<�p�<֎�<]��<���<|��<���<B	�<f�</+�<�8�<�C�<KL�<FR�<�U�<VV�<,T�<HO�<`G�<�<�<�.�<��<�	�<(��<���<t��<��<s�<�J�<��<��<��<��<JJ�<��<���<���<�9�<��<���<*E�<���<�<�-�<�ȿ<h`�<��<ڃ�<��<P��<�<,��<��<˕�<z�<��<��<@\�<�Ū<,�<j��<��<cM�<1��<K �<�U�<ͨ�<f��<�G�<˓�<�ݖ<�%�<�k�<��<��<�3�<s�<4��<�<�)�<;d�<͝�<�ց<��<��|<��x<jfu<��q<q>n<�j<�g<�c<��_<�Z\<w�X<a7U<��Q<LN<،J<0G<�yC<��?<;p<<��8<�q5<t�1<R�.<�+<V�'<�1$<�� <�g<e	<�<�[<J<��<L~	<�?<<<:��;�P�; �;u��;(��;nq�;�[�;T�;�Z�;\p�;���;�Ǽ;�	�;�[�;L��;�,�;���;S<�;�ە;y��;bI�;��;���;��w;��m;E�c;�Z;�jP;T�F;�r=;#4;K�*;��!;
�;z;�D;�=�:�%�:rC�:���:6�:=ǩ:���:	��:�s:M�T:>�5:k:�u�9ޭ�9_w9��9�g\7Fwʸ.W����ܹ1�	�}P%��@� �[�ѣv�I���������7��n:��Q+ʺi׺#�㺤��k:��Y��2��r�v�����d$��8*��]0��}6��<���B��H���N���T���Z�$a��g�7m�@ s��'y�H.���������ա������۪��m���궔�a����ƚ��  �  �f=M=��=�A=��==}=�=�� =:T =��<�<P�<d��<���<+��<�#�<"V�<���<���<���<��<2A�<^l�<0��<���<a��<�
�<R.�<@P�<tp�<ߎ�<a��<���<t��<���<F	�<X�<3+�<�8�<�C�<FL�<BR�<�U�<NV�<2T�<@O�<jG�<�<�<�.�<��<�	�<1��<���<y��<��<s�<�J�<��<��<��<��<AJ�<��<���<���<�9�<��<���<#E�<���<���<�-�<ɿ<e`�<��<̃�<��<N��<
�<2��<��<֕�<k�<��<��<?\�<�Ū<,�<q��<��<lM�<.��<G �<�U�<Ϩ�<i��<�G�<Ó�<�ݖ<�%�<�k�<��<��<�3�<s�</��<�<�)�<6d�<՝�<�ց<��<�|<��x<xfu<��q<y>n<��j<�g<m�c<��_<�Z\<��X<p7U<��Q<JN<ӌJ<:G<�yC<��?<;p<<��8<�q5<_�1<^�.<�+<\�'<�1$<s� <�g<S	<��<�[<^<��<@~	<�?<&<S��;�P�;��;{��;#��;fq�;�[�;=T�;[�;sp�;}��;�Ǽ;�	�;X[�;\��;�,�;���;?<�;|ە;{��;CI�;��;���;.�w;��m;N�c;�Z;ajP;��F;�r=;@#4;*�*;��!;��;2;�D;�=�:K&�:�B�:ޒ�:��:�Ʃ:'��:���:��s:p�T:q�5:�j:�s�9$��9�w9��9��[7�uʸ�.W�	��>
ܹ	�	�%O%��@���[��v�V�������U7��;���*ʺ�׺d����D:��:��[2��r�������X$��8*��]0�f~6���<���B�5�H���N���T���Z�Ka��g�~m�' s�['y�3.�v����������"���ݪ��\���϶��E���ǚ��  �  �f=H=��=�A=��=?}=�=�� =6T =!��<��<P�<[��<���<C��<�#�<V�<x��<���<���<��<.A�<[l�<8��<���<i��<�
�<L.�<TP�<up�<��<Y��<���<|��<���<D	�<V�<:+�<�8�<�C�<@L�<JR�<�U�<HV�<;T�<<O�<lG�<�<�<�.�<��<�	�<7��<|��<z��<���<$s�<�J�<��<��<ػ�<��<<J�<��<���<���<�9�<��<���<E�<���<ʎ�<�-�<ɿ<^`�<��<̃�<��<N��<�<2��<��<ە�<j�<��<��<:\�<�Ū<,�<z��<��<iM�<*��<G �<�U�<ƨ�<h��<�G�<ړ�<�ݖ<�%�<�k�<��<��<�3�<s�<2��<�<�)�<6d�<؝�<�ց<��<�|<��x<yfu<��q<�>n<��j<�g<i�c<��_<�Z\<��X<o7U<��Q<pN<��J<;G<�yC<��?<Cp<<��8<�q5<Q�1<c�.<�+<R�'<�1$<x� <�g<V	<�<{[<R<��<8~	<�?<!<s��;�P�;�;g��;��;�q�;�[�;RT�;�Z�;bp�;���;�Ǽ;�	�;Q[�;y��;�,�;Ȭ�;+<�;�ە;���;)I�;��;���;C�w;��m;H�c;�Z;0jP;��F;jr=;H#4;��*;�!;Q�;;
E;"=�:�&�:�B�:���:n�:�Ʃ:s��:K��:B�s:��T:�5:l:Lr�9\��9�w9��9��[7�vʸ�.W����D
ܹ*�	��N%���@�"�[�I�v�����B񕺡���6��d;���*ʺ�׺d��8���:��H��X2�r�������e$�9*��]0��~6�Ú<���B�%�H���N���T�k�Z��a�.g�jm�< s�X'y�z.�^���/���ϡ��)�������}���ض��F���ǚ��  �  �f=L=��=�A=��=<}=�=�� =AT =��<��< P�<_��<»�<)��<�#�<V�<���<���<���<��<)A�<fl�<.��<���<h��<�
�<N.�<CP�<zp�<׎�<`��<���<z��<���<C	�<d�<1+�<�8�<�C�<AL�<HR�<�U�<OV�<3T�<CO�<eG�<�<�<�.�<��<�	�<-��<��<|��<
��<s�<�J�<��<��<ݻ�<��<JJ�<��<���<���<�9�<��<���<%E�<���<Ď�<�-�< ɿ<e`�<��<փ�<��<Q��<�<-��<��<Ε�<n�<��<��<=\�<�Ū<,�<p��<��<fM�<1��<O �<�U�<Ϩ�<h��<�G�<Ó�<�ݖ<�%�<�k�<��<��<�3�<s�<6��< �<�)�<:d�<ӝ�<�ց<��<�|<��x<{fu<��q<n>n<�j<�g<��c<��_<�Z\<��X<X7U<��Q<PN<όJ<7G<�yC<��?<8p<<��8<�q5<|�1<[�.<�+<a�'<�1$<}� <�g<_	<�<�[<H<��<M~	<�?<6<J��;�P�;�;l��;��;uq�;�[�;T�;[�;Xp�;���;�Ǽ;�	�;�[�;T��;�,�;���;,<�;�ە;t��;EI�;��;���;�w;��m;U�c;�Z;�jP;{�F;�r=;Z#4;7�*;��!;��;[;E;x=�:&�:gC�:���:b�:ǩ:騙:ǹ�:0�s:��T:��5:]k:�r�9���9�w97�9�G\7�vʸ�-W�����ܹ%�	�P%���@�ڻ[�|�v�|�����V��q7���:��!+ʺh׺��㺝��L:��G��/2��r�������1$�9*��]0��}6��<���B�>�H���N���T���Z�Pa��g�Qm�q s�R'y�^.�����񝅻ʡ������䪎�t���ɶ��s����ƚ��  �  �f=T=��=�A=��=:}=�=�� =>T =��<�<P�<Z��<ͻ�<&��<�#�<V�<���<���<���<��<(A�<dl�<'��<���<^��<�
�<^.�<<P�<�p�<َ�<h��<���<v��<���<>	�<c�<)+�<�8�<�C�<OL�<NR�<�U�<ZV�<&T�<JO�<aG�<�<�<�.�<��<�	�< ��<���<q��<��<!s�<�J�<��<��<��<���<BJ�<��<���<���<�9�<��<}��</E�<���<Ȏ�<�-�< ɿ<o`�<��<Ճ�<��<Q��<�<+��<��<͕�<}�<��<��<A\�<�Ū<#,�<h��<��<dM�<+��<D �<�U�<֨�<]��<�G�<���<�ݖ<�%�<�k�<!��<��<�3�<s�<4��<��<�)�<:d�<˝�<�ց<��<�|<��x<zfu<��q<a>n<�j<�g<��c<��_<�Z\<��X<f7U<��Q<=N<�J<+G<�yC<��?<.p<<��8<�q5<m�1<?�.<�+<Y�'<�1$<�� <|g<u	<ܯ<�[<M<u�<A~	<�?<2<.��;�P�;��;g��;S��;Xq�;\�;$T�;)[�;\p�;���;�Ǽ;�	�;�[�;3��;�,�;���;c<�;�ە;z��;rI�;z�;���;��w;��m;:�c;XZ;~jP;�F;�r=;�"4;W�*;��!;��;�;�D;3>�:]%�:�B�::��:4�:�Ʃ:x��:W��:��s:��T:��5:�k:�v�9���9�
w9N�9�;\7d{ʸZ-W�Y��ܹ�	�6P%���@�}�[���v�=���.�y���7���:��C+ʺ�׺���ŏ��9������1��r�E�����t$��8*�<^0�%~6��<���B�[�H���N���T���Z��a��g��m�2 s�T'y�.�����񝅻案���������S�������Y����ƚ��  �  �f=M=��=�A=��=?}=�=�� ==T =��<�<P�<Y��<ǻ�<7��<�#�<V�<~��<���<���<��<4A�<]l�<2��<���<e��<�
�<T.�<EP�<xp�<َ�<Z��<���<~��<���<G	�<^�<3+�<�8�<�C�<BL�<CR�<�U�<OV�<3T�<EO�<fG�<�<�<�.�<��<�	�</��<���<o��<��<#s�<�J�<��<��<��<��<IJ�<��<���<���<�9�<��<���<%E�<���<���<�-�<�ȿ<c`�< ��<Ӄ�<��<U��<�<0��<��<Ε�<m�<��<��<<\�<�Ū<,�<r��<��<oM�<5��<M �<�U�<Ψ�<_��<�G�<ѓ�<�ݖ<�%�<�k�<��<��<�3�< s�<2��<�<�)�<<d�<ӝ�<�ց<��<�|<��x<jfu<��q<u>n<�j<�g<|�c<��_<�Z\<u�X<c7U<��Q<UN<ӌJ<5G<�yC<��?<@p<<��8<�q5<j�1<[�.<�+<M�'<�1$<�� <�g<i	<ܯ<�[<U<��<M~	<�?<$<[��;�P�;�;f��;*��;{q�;�[�;#T�;�Z�;ap�;���;�Ǽ;�	�;o[�;\��;�,�;���;2<�;}ە;���;GI�;��;���;�w;��m;^�c;�Z;�jP;��F;�r=;�"4;�*;�!;,�;A;�D;�=�:C&�:aC�:<��:��:�Ʃ:�:ù�:5�s:��T:h�5:�j:s�9(��9gw9��9�1\7�rʸ�+W�2���
ܹ��	�)P%���@��[�ޣv�������P��O7��;;���*ʺ'׺���B��c:�����2�ar�Y������$��8*��]0�-~6���<���B�#�H���N���T���Z�Fa��g�om�I s��'y�V.�~���	���ϡ�����Ϫ��t����]���ǚ��  �  �f==q�=�A=b�=�|=;=>� =�S =[��<#�<3O�<c��<���<��<}"�<�T�<(��<Y��<X��<�<�?�<�j�<r��<���<s��<��<*,�<N�<2n�<~��<֨�<Z��<���<2��<x�<k�<1(�<}5�<v@�<�H�<�N�<!R�<�R�<�P�<gK�<�C�<�8�<�*�<��<G�<���<��<���<p��<qn�<�E�<��<P��<���<��<@E�<��<���<}~�<�4�<���<o��<�?�<���<���<�(�<�ÿ<N[�<�<�~�<�<z��<E�<w��<�<E��<��<M{�<E�<X�<���<(�<���<�<�I�<���<���<�R�<���<u��<�D�<��<5ۖ<X#�<�i�<���<���<�1�<sq�<���<��<j(�<c�<ᜃ<�Ձ<��<��|<��x<�eu<��q<�>n<��j<�g<��c<2�_<_\\<g�X<�9U<8�Q<LN<�J<�G<�}C<��?<�t<<-�8<�v5<��1<��.<�+<��'<28$<#� <{n<�<l�<Cc<]<��<��	<�H<<߻�;�c�;H�;���;���;��;�p�;Bi�;p�;��;d��;�ݼ;d �;�q�;
ӫ;6C�;Yà;%S�;p�;x��;�_�;�.�;c�;��w;��m;,d;�?Z;S�P;�G;��=;:N4;<+;J";�;�.;�l;H��:=s�:���:���:�\�:��:��:>��:st:�AU:j6:��:?`�9��9c�x9��9*0v7�BǸv�U��Q��T۹�p	���$�tM@��k[�8Xv�u���#Ε��������O��ʺx�ֺ��㺵t�!��<���&�h������$�x0*�WU0��v6�u�<��B��H��N���T���Z�qa��g�
m�8s�W%y�e,�����j���>���ܥ��ժ���������������ǚ��  �  �f=#=t�=�A=a�=�|===8� =�S =R��<�<0O�<[��<���<��<�"�<�T�<*��<M��<T��<�<�?�<�j�<l��<���<s��<��<9,�<N�</n�<}��<��<]��<���<)��<c�<m�<)(�<�5�<�@�<�H�<�N�< R�<�R�<�P�<kK�<�C�<�8�<�*�<��<Q�<���<��<��<o��<}n�<�E�<��<@��<���<��<GE�<��<���<�~�<�4�<���<m��<@�<���<���<�(�<�ÿ<a[�< �<�~�<�
�<p��<F�<y��<%�<F��<��<B{�<Q�<X�<���<(�<���<�<�I�<���<���<�R�<���<g��<�D�<��<Aۖ<R#�<�i�<�<���<�1�<jq�<���<��<f(�<c�<䜃<�Ձ<��<�|<��x<fu<��q<�>n<��j<`g<��c<'�_<m\\<��X<�9U<0�Q<<N<�J<�G<�}C<��?<�t<<4�8<�v5<��1<�.<�+<y�'<#8$<6� <�n<�<W�<Gc<D<��<��	<H<<Ļ�;�c�;J�;��;6��;���;xp�;<i�;lp�;���;\��;�ݼ; �;�q�;�ҫ;uC�;�à;"S�;J�;t��;<`�;�.�;t�;s�w;��m;�d;�?Z;��P;G;ɝ=;�M4;;+;�";6;�.;�l;f��:Zr�:#��:	��:3\�:	�:��:i��:�rt:�CU:Yj6:M�:N`�9W��9��x9��9�Av7�TǸ��U��Q���S۹n	���$��M@�9m[��Vv�l���Ε�����������$ʺ�ֺҸ㺘u�~!������&��g�(��@��?$��0*��U0��v6���<�*�B� �H�>�N���T���Z�� a��g�6m�Gs��$y�,�����q�������祋�쪎�����:��������ǚ��  �  �f=!=n�=�A=c�=�|=@=4� =�S =N��<'�<9O�<]��<���<��<�"�<�T�<7��<R��<S��<�<�?�<�j�<i��<���<r��<��<7,�<N�<6n�<m��<��<T��<���<4��<e�<x�<(�<�5�<t@�<�H�<�N�<R�<�R�<uP�<wK�<~C�<�8�<�*�<��<W�<���<��<��<r��<nn�<�E�<��<?��<��<��<ME�<��<���<�~�<�4�<���<a��<�?�<���<���<�(�<�ÿ<_[�<��<�~�< �<z��<J�<o��<#�<8��<��<D{�<L�<X�<���<$(�<���<%�<�I�<���<���<�R�<���<g��<�D�<��<9ۖ<V#�<�i�<���<���<�1�<dq�<���<��<i(�<$c�<ל�<�Ձ<��<��|<��x<	fu<��q<�>n<��j<dg<��c<"�_<`\\<��X<�9U<B�Q<9N<�J<�G<�}C<��?<�t<<A�8<�v5<��1<�.<�+<��'<(8$<)� <pn<�<Y�<`c<M<��<Ȇ	<qH<1<���;�c�;E�;���;/��;Ņ�;�p�;�h�;^p�;Յ�;f��;�ݼ; �;r�;�ҫ;lC�;Pà;S�;e�;`��;`�;h.�;��;b�w;�m;d;@Z;ٖP;G;,�=;�M4;O+;/";�;�.;ul;>��:Er�:|��:2��:F\�:��:��:#��:Zqt:�BU:zi6:��:�`�9���9��x9�~9��v7�OǸ̤U�nP��V۹On	���$��L@��l[�RWv�/����Ε��������7��mʺ��ֺ���{u� ������&�0h�g��"��$�70*��U0�zv6��<�
�B���H�"�N���T�1�Z�a��g��m��s�%y�7,�̙��F�������������������T���,����ǚ��  �  �f= =r�=�A=b�=�|=<=;� =�S =Q��<%�<+O�<a��<���<��<�"�<�T�<#��<V��<R��<�<�?�<�j�<h��<���<u��<��<5,�<N�<-n�<x��<��<b��<���<+��<h�<j�<+(�<�5�<{@�<�H�<�N�< R�<�R�<}P�<qK�<{C�<�8�<�*�<��<J�<���<��<��<q��<yn�<�E�<��<B��<��<��<AE�<��<���<�~�<�4�<���<j��<@�<���<���<�(�<�ÿ<a[�<�<�~�< �<s��<D�<}��<"�<B��<��<H{�<L�<	X�<���<(�<���<�<�I�<���<���<�R�<���<m��<�D�<��<=ۖ<W#�<�i�<���<���<�1�<nq�<���<��<e(�< c�<���<�Ձ<��<�|<��x<fu<��q<�>n<��j<sg<��c<.�_<u\\<��X<�9U<5�Q<AN<�J<�G<�}C<��?<�t<<1�8<�v5<��1<�.<�+<n�'</8$</� <�n<�<d�<8c<V<��<��	<�H<<���;�c�;P�;���;$��;ԅ�;mp�;*i�;\p�;��;`��;�ݼ;! �;�q�;�ҫ;�C�;mà;S�;a�;v��;`�;�.�;��;G�w;��m;d;)@Z;o�P;MG;��=;�M4;I+;�";;�.;�l;��:�r�:Ǎ�:@��:y\�:�:��:���:vrt:CU:j6:�:�_�9��9��x9}�9�0v7�PǸB�U��Q���R۹cn	�]�$�5N@��l[�ZWv����Ε�g���������ʺ�ֺ���u��!��z���&��g�E����d$�p0*��U0��v6���<�*�B�$�H�?�N���T���Z�'a��g�m�Zs��$y��+���������q�������ު������P���	����ǚ��  �  �f==s�=�A=b�=�|=:=>� =�S =W��<%�<1O�<e��<���<��<s"�<�T�<'��<Z��<S��<�<�?�<�j�<s��<���<s��<��<2,�<N�<*n�<���<ݨ�<_��<���<1��<w�<h�<,(�<5�<�@�<�H�<�N�<%R�<�R�<P�<iK�<�C�<�8�<�*�<��<D�<���<��<��<i��<xn�<�E�<��<P��<��<��<=E�<��<���<�~�<�4�<���<k��<�?�<���<���<�(�<�ÿ<Q[�<�<�~�<�<{��<B�<|��<�<K��<��<L{�<L�<X�<���<(�<���<�<�I�<���<���<�R�<���<y��<�D�<"��<6ۖ<W#�<�i�<���<���<�1�<uq�<���<��<h(�<c�<圃<�Ձ<��<�|<��x<fu<��q<�>n<~�j<�g<��c<.�_<b\\<{�X<�9U<.�Q<KN<��J<�G<�}C<��?<�t<<)�8<�v5<��1<��.<�+<|�'<78$<� <�n<~<z�<@c<_<��<��	<�H<<��;�c�;I�;���;��;��;ap�;Vi�;.p�;��;[��;�ݼ;_ �;�q�;�ҫ;=C�;�à; S�;`�;���;`�;�.�;l�;��w;��m;d;X@Z;B�P;�G;��=;JN4;	+;|";;E.;�l;#��:Ns�:���:���:�\�:��:N�:9��:�rt:�BU:�j6:S�:�_�9Ε�9��x9%�9}v7�BǸ$�U�cR���R۹<p	�@�$��N@�l[�hWv�툈�!Ε�����	��[���ʺ��ֺ
�㺻t�!����I'��g������$�k0*�rU0�	w6�^�<�>�B���H�*�N���T���Z�;a��g�3m�(s��$y�`,���������3�������ݪ������c����Ț��  �  �f==r�=�A=`�=�|=?=9� =�S =P��< �<0O�<d��<���<��<{"�<�T�<)��<O��<Q��<�<�?�<�j�<b��<���<y��<��<0,�<N�<4n�<w��<��<[��<���<2��<i�<p�<((�<�5�<~@�<�H�<�N�<R�<�R�<P�<xK�<wC�<�8�<�*�<��<O�<���<��<���<s��<yn�<�E�<��<D��<��<��<DE�<��<���<�~�<�4�<���<m��<�?�<���<���<�(�<�ÿ<\[�<��<�~�<�<w��<E�<x��<�<@��<��<N{�<J�<X�<���<!(�<���<�<�I�<���<���<�R�<���<p��<�D�<��<:ۖ<[#�<�i�<�<���<�1�<kq�<���<��<_(�<&c�<✃<�Ձ<��<��|<��x<fu<��q<�>n<��j<jg<��c<+�_<b\\<��X<�9U<G�Q<BN<��J<�G<�}C<��?<�t<<=�8<�v5<��1<�.<�+<x�'<58$<#� <�n<�<l�<Dc<I<��<Ɔ	<}H<'<���;�c�;b�;���;��;��;�p�;'i�;Np�;��;^��;�ݼ;% �;�q�;�ҫ;eC�;wà;S�;��;n��;`�;�.�;��;+�w;��m; d;(@Z;��P;,G;��=;�M4;W+;�";;�.;�l;6��:tr�:���:d��:@\�:,�:O�:��:�rt:�BU:j6:	�:�_�9(��9l�x9�9�Sv7�NǸl�U��Q���S۹�n	���$��M@��k[��Wv�∈��͕�$���/�����$ʺ��ֺ��}u�!��d���&��g�`�����I$��0*��U0��v6���<��B�8�H�q�N�w�T���Z�1a��g��m�cs��$y�P,�����c�������ե��㪎�����N�������ǚ��  �  �f=&=o�=�A=b�=�|=C=3� =�S =G��<+�<-O�<^��<���<��<�"�<�T�<,��<V��<L��<�<�?�<�j�<]��<���<k��<��<8,�<
N�<4n�<r��<��<V��<���<3��<d�<v�<(�<�5�<z@�<�H�<�N�<R�<�R�<pP�<{K�<wC�<�8�<�*�<��<Q�<���<��<��<u��<un�<�E�<��<:��<��<��<EE�<��<���<�~�<�4�<���<^��<	@�<���<���<�(�<�ÿ<d[�<��<�~�<�
�<w��<H�<p��<(�<:��<��<C{�<L�<X�<���<((�<���<(�<�I�<���<���<�R�<���<f��<�D�<��<>ۖ<V#�<�i�<���<���<�1�<aq�<���<��<b(�<$c�<؜�<�Ձ<��<��|<��x<fu<��q<�>n<��j<_g<��c<�_<f\\<��X<�9U<G�Q<-N<�J<�G<�}C<��?<�t<<N�8<�v5<��1<օ.<�+<s�'<)8$<2� <zn<�<X�<Kc<U<��<ʆ	<kH<9<���;�c�;+�;���;0��;���;�p�;i�;lp�;݅�;`��;�ݼ; �;�q�;�ҫ;�C�;eà;S�;m�;X��;F`�;U.�;��;*�w;��m;d;�?Z;��P;�
G;�=;�M4;j+;k";�;�.;Ql;��:?r�:���:���:-\�:��:2�:t��:�pt:DU:�i6:
�:D_�9i��9��x9�~9�~v7�QǸ.�U�Q���U۹�m	�P�$��M@�m[�OWv�ǈ���Ε�����������ʺ��ֺ0��Gu� !������&�	h�@�� ��s$�*0*��U0��v6���<�ݬB�6�H�]�N���T�.�Z�� a�	g��m��s��$y�*,�֙��P�������ɥ����������;���$����ǚ��  �  �f=!=p�=�A=f�=�|===9� =�S =K��<&�<-O�<c��<���<��<�"�<�T�<&��<V��<Q��<�<�?�<�j�<i��<���<j��<��<2,�<N�<3n�<|��<ߨ�<\��<���<1��<m�<l�<((�<�5�<w@�<�H�<�N�<R�<�R�<tP�<tK�<�C�<�8�<�*�<��<Q�<���<��<���<q��<vn�<�E�<��<E��<���<��<FE�<��<���<�~�<�4�<���<a��<@�<���<���<�(�<�ÿ<X[�<��<�~�<�<y��<G�<y��<�<B��<��<K{�<H�<
X�<���<&(�<���<�<�I�<���<���<�R�<���<o��<�D�<��<<ۖ<W#�<�i�<���<���<�1�<mq�<���<��<o(�<c�<ܜ�<�Ձ<��<��|<��x<fu<��q<�>n<��j<}g<��c<,�_<h\\<{�X<�9U<B�Q<@N<�J<�G<�}C<��?<�t<<4�8<�v5<��1<ޅ.<�+<s�'<48$<.� <�n<�<i�<?c<W<��<φ	<}H<<���;�c�;'�;���;��;߅�;�p�;8i�;6p�;���;l��;�ݼ;7 �;�q�;�ҫ;\C�;]à;S�;v�;l��;!`�;f.�;��;��w;��m;d;:@Z;��P;*G;ٝ=;�M4;H+;o";�;�.;�l;���:�r�:��:���:b\�:�:�:��:Rqt:CU:�i6:��:q_�9Ғ�9`�x9��9M=v7$KǸ'�U�4Q���S۹�o	�\�$��M@� l[��Wv������Ε�����������!ʺy�ֺ��u�!��j���&��g�Q����P$�Z0*��U0��v6���<�-�B�(�H���N���T��Z�a��g��m�Vs�%y�5,�����x���\���륋�⪎�����c�������ǚ��  �  �f==w�=�A=a�=�|===;� =�S =V��< �</O�<d��<���<%��<v"�<�T�<"��<T��<V��<�<�?�<�j�<k��<���<u��<��</,�<N�<$n�<���<��<c��<���<-��<q�<b�<2(�<�5�<�@�<�H�<�N�<'R�<�R�<�P�<iK�<�C�<�8�<�*�<��<J�<���<��<���<n��<}n�<F�<��<I��<��<��<CE�<��<���<�~�<�4�<���<q��<�?�<���<���<�(�<�ÿ<W[�<�<�~�<�<v��<>�<���<�<M��<��<R{�<H�<X�<���<(�<���<�<�I�<���<���<�R�<���<s��<�D�<(��<9ۖ<W#�<�i�<�<���<�1�<oq�<���<��<f(�<c�<휃<�Ձ<��<�|<��x<fu<��q<�>n<y�j<�g<��c<2�_<i\\<��X<�9U<'�Q<VN<�J<�G<�}C<��?<�t<<4�8<�v5<��1<�.<�+<w�'<58$< � <�n<�<r�<8c<S<��<��	<�H<<Ļ�;�c�;P�;��;��;��;Mp�;Zi�;Bp�;��;R��;�ݼ;G �;�q�;ӫ;ZC�;�à;S�;n�;���;�_�;�.�;m�;��w;��m;*d;&@Z;q�P;yG;u�=;N4;1+;�";Q;v.;�l;Ɗ�:/s�:��:M��:�\�:�:��:9��:^st:dBU:�j6:��:#^�9k��9ݿx9n�9a�u7�IǸy�U�qS��MQ۹�o	��$�KO@�Bk[��Wv�ʈ���͕�����������ʺ�ֺǸ�u�"��L��$'�^g�k����3$��0*�|U0��v6���<�'�B�+�H�:�N���T���Z�xa�dg�>m�<s��$y�B,���������D�������ժ������J���ﾗ�Ț��  �  �f==s�=�A=c�=�|=?=8� =�S =N��<&�<6O�<d��<���<��<w"�<�T�<2��<T��<Q��<�<�?�<�j�<f��<���<p��<��<0,�<N�<)n�<|��<��<X��<���<4��<m�<q�<&(�<�5�<~@�<�H�<�N�<$R�<�R�<{P�<pK�<�C�<�8�<�*�<��<M�<���<��<���<p��<sn�<�E�<��<H��<���<��<DE�<��<���<�~�<�4�<���<f��<�?�<���<���<�(�<�ÿ<V[�<��<�~�<�<z��<D�<u��<�<E��<��<L{�<I�<	X�<���<(�<���<�<�I�<���<���<�R�<���<r��<�D�<��<4ۖ<X#�<�i�<���<���<�1�<iq�<���<��<i(�<c�<㜃<�Ձ<��<�|<��x<fu<��q<�>n<��j<wg<��c<'�_<\\\<��X<�9U<+�Q<KN<��J<�G<�}C<��?<�t<<;�8<�v5<��1<�.<�+<��'<58$<� <�n<�<r�<Vc<R<��<��	<�H<!<���;�c�;@�;���;��;��;ap�;<i�;Ap�;��;]��;�ݼ;7 �;�q�;�ҫ;OC�;wà;S�;b�;���;`�;�.�;��;��w;��m;d;@Z;��P;6G;�=;N4;B+;W";�;�.;�l;ċ�:�r�:���:#��:`\�:$�:��:���:�qt:�BU:lj6:Q�:�^�9p��94�x9�9FYv70KǸϤU��Q���T۹�o	���$��N@�l[��Wv�����Ε�K����������ʺ
�ֺ��@u�!��O��'��g������$�G0*��U0��v6���<��B�C�H�%�N���T���Z�Ua��g�/m�Qs��$y�h,�����a���i���ѥ��몎�����O������Ț��  �  �f=#=t�=�A=d�=�|=@=6� =�S =E��<'�<*O�<_��<���<��<�"�<�T�<*��<O��<K��<�<�?�<�j�<^��<���<u��<��<4,�<N�<7n�<u��<��<_��<���<.��<_�<s�< (�<�5�<v@�<�H�<�N�<R�<�R�<|P�<wK�<zC�<�8�<�*�<��<U�<���<��<��<x��<yn�<�E�<��<;��<���<��<IE�<��<���<�~�<�4�<���<g��<@�<���<���<�(�<�ÿ<i[�<��<�~�<�
�<q��<E�<w��<(�<=��< �<F{�<K�<X�<���<%(�<���<�<�I�<���<���<�R�<���<f��<�D�<��<?ۖ<X#�<�i�<���<���<�1�<eq�<���<��<h(�<"c�<㜃<�Ձ<��<��|<��x<fu<��q<�>n<��j<Vg<��c<�_<|\\<��X<�9U<E�Q<1N<�J<�G<�}C<��?<�t<<?�8<�v5<��1<҅.<�+<m�'<,8$<8� <~n<�<\�<Fc<I<��<ǆ	<|H<%<���;�c�;P�;��; ��;�;�p�; i�;hp�;��;\��;�ݼ;��;�q�;�ҫ;�C�;Yà;)S�;n�;]��;D`�;�.�;��;D�w;��m;d;�?Z;ʖP;�
G;��=;�M4;�+;�";;�.;Wl;���:r�:H��:���:#\�:��:_�:%��:rt:nDU:�i6:i�:la�9Z��9��x9��9u^v7�XǸa�U��Q��T۹�m	��$��L@��l[��Wv�X���MΕ�����>�����Hʺ��ֺ�㺠u�n!������&��g�7�����$�?0*�(V0��v6�ߓ<��B�d�H�.�N���T���Z�� a��g��m�Os�%y��+�֙��c�������ۥ�� ������M�������ǚ��  �  �f==t�=�A=a�=�|=A=7� =�S =Q��<,�<2O�<a��<���<��<|"�<�T�<-��<Y��<S��<�<�?�<�j�<k��<���<r��<��<0,�<N�<1n�<z��<��<]��<���<7��<o�<r�<!(�<�5�<v@�<�H�<�N�<R�<�R�<P�<mK�<�C�<�8�<�*�<��<P�<���<��<���<r��<on�<�E�<��<G��<���<��<GE�<��<���<�~�<�4�<���<k��<�?�<���<���<�(�<�ÿ<[[�<��<�~�<�<}��<B�<v��<�<@��<��<G{�<H�<
X�<���<(�<���<$�<�I�<���<���<�R�<���<q��<�D�<��<4ۖ<W#�<�i�<���<���<�1�<eq�<���<��<f(�<c�<圃<�Ձ<��<�|<��x<fu<��q<�>n<��j<zg<��c<�_<i\\<v�X<�9U<9�Q<@N<��J<�G<�}C<��?<�t<<D�8<�v5<��1<�.<�+<|�'<.8$<"� <{n<�<j�<Lc<]<��<��	<�H<-<»�;�c�;G�;��;��;؅�;p�;2i�;Ap�;���;O��;�ݼ;A �;�q�;�ҫ;cC�;Wà; S�;c�;h��;`�;�.�;}�;��w; �m;Bd;�?Z;��P;YG;�=;�M4;Q+;:";�;�.;�l;Ћ�: s�:!��:���:�\�:��:�:z��:�rt:�BU:�i6:�:A`�9���9��x9��9kMv7�GǸ	�U�iR��YT۹�n	���$��M@��l[��Wv�����@Ε�����s��O��ʺ`�ֺԸ��t�F!��_���&�h������<$�0*��U0��v6��<��B��H�9�N���T���Z�=a��g�m�Fs�.%y�+,�ڙ��P���c���ť���������m��������ǚ��  �  �f==u�=�A=`�=�|=:=;� =�S =T��<�<+O�<e��<���<#��<}"�<�T�<!��<I��<U��<�<�?�<�j�<h��<���<w��<��<3,�<N�<(n�<���<��<f��<���<+��<`�<l�<0(�<�5�<�@�<�H�<�N�<&R�<�R�<�P�<lK�<�C�<�8�<�*�<��<Q�<���<��<���<p��<|n�<F�<��<J��<��<��<GE�<��<���<{~�<�4�<���<w��<�?�<���<���<�(�<�ÿ<Y[�<	�<�~�<�
�<r��<D�<���<�<M��<��<G{�<L�<	X�<���<(�<���<�<�I�<���<���<�R�<���<y��<�D�<)��<;ۖ<Z#�<�i�<譑<���<�1�<mq�<���<��<e(�<c�<꜃<�Ձ<��<ڊ|<��x<fu<��q<�>n<��j<bg<��c<+�_<l\\<��X<�9U<'�Q<XN<�J<�G<�}C<��?<�t<<(�8<�v5<��1<��.<�+<p�'<88$<+� <�n<�<{�<5c<=<��<��	<�H<<���;vc�;Z�;��;��;��;Zp�;fi�;Cp�;��;a��;�ݼ; �;�q�;ӫ;WC�;�à;!S�;H�;���;�_�;�.�;w�;��w;x�m;�d;7@Z;��P;=G;Y�=;�M4;D+;�";N;�.;�l;���:�r�:!��:k��:H\�:��:#�:P��:tt:BU:�j6:m�:_�9��9��x9ԉ9�0v7�TǸ�U�R��}Q۹ o	��$��N@��l[�OWv�����͕��������_���ʺ��ֺ��㺡u�9"�����&�Sg�U����`$��0*��U0��v6���<�a�B�]�H�C�N���T���Z�ta�Yg�`m�s��$y�<,�����n�������䥋�㪎�����P���ܾ��Ț��  �  �f==t�=�A=a�=�|=A=7� =�S =Q��<,�<2O�<a��<���<��<|"�<�T�<-��<Y��<S��<�<�?�<�j�<k��<���<r��<��<0,�<N�<1n�<z��<��<]��<���<7��<o�<r�<!(�<�5�<v@�<�H�<�N�<R�<�R�<P�<mK�<�C�<�8�<�*�<��<P�<���<��<���<r��<on�<�E�<��<G��<���<��<GE�<��<���<�~�<�4�<���<k��<�?�<���<���<�(�<�ÿ<[[�<��<�~�<�<}��<B�<v��<�<@��<��<G{�<H�<
X�<���<(�<���<$�<�I�<���<���<�R�<���<q��<�D�<��<4ۖ<W#�<�i�<���<���<�1�<eq�<���<��<f(�<c�<圃<�Ձ<��<�|<��x<fu<��q<�>n<��j<zg<��c<�_<i\\<v�X<�9U<9�Q<@N<��J<�G<�}C<��?<�t<<D�8<�v5<��1<�.<�+<|�'<.8$<"� <{n<�<j�<Lc<]<��<��	<�H<-<»�;�c�;G�;��;��;؅�;p�;2i�;Ap�;���;O��;�ݼ;A �;�q�;�ҫ;cC�;Wà; S�;c�;h��;`�;�.�;}�;��w; �m;Bd;�?Z;��P;YG;�=;�M4;Q+;:";�;�.;�l;Ћ�: s�:!��:���:�\�:��:�:z��:�rt:�BU:�i6:�:A`�9���9��x9��9kMv7�GǸ	�U�iR��YT۹�n	���$��M@��l[��Wv�����@Ε�����s��O��ʺ`�ֺԸ��t�F!��_���&�h������<$�0*��U0��v6��<��B��H�9�N���T���Z�=a��g�m�Fs�.%y�+,�ڙ��P���c���ť���������m��������ǚ��  �  �f=#=t�=�A=d�=�|=@=6� =�S =E��<'�<*O�<_��<���<��<�"�<�T�<*��<O��<K��<�<�?�<�j�<^��<���<u��<��<4,�<N�<7n�<u��<��<_��<���<.��<_�<s�< (�<�5�<v@�<�H�<�N�<R�<�R�<|P�<wK�<zC�<�8�<�*�<��<U�<���<��<��<x��<yn�<�E�<��<;��<���<��<IE�<��<���<�~�<�4�<���<g��<@�<���<���<�(�<�ÿ<i[�<��<�~�<�
�<q��<E�<w��<(�<=��< �<F{�<K�<X�<���<%(�<���<�<�I�<���<���<�R�<���<f��<�D�<��<?ۖ<X#�<�i�<���<���<�1�<eq�<���<��<h(�<"c�<㜃<�Ձ<��<��|<��x<fu<��q<�>n<��j<Vg<��c<�_<|\\<��X<�9U<E�Q<1N<�J<�G<�}C<��?<�t<<?�8<�v5<��1<҅.<�+<m�'<,8$<8� <~n<�<\�<Fc<I<��<ǆ	<|H<%<���;�c�;P�;��; ��;�;�p�; i�;hp�;��;\��;�ݼ;��;�q�;�ҫ;�C�;Yà;)S�;n�;]��;D`�;�.�;��;D�w;��m;d;�?Z;ʖP;�
G;��=;�M4;�+;�";;�.;Wl;���:r�:H��:���:#\�:��:_�:%��:rt:nDU:�i6:i�:la�9Z��9��x9��9u^v7�XǸa�U��Q��T۹�m	��$��L@��l[��Wv�X���MΕ�����>�����Hʺ��ֺ�㺠u�n!������&��g�7�����$�?0*�(V0��v6�ߓ<��B�d�H�.�N���T���Z�� a��g��m�Os�%y��+�֙��c�������ۥ�� ������M�������ǚ��  �  �f==s�=�A=c�=�|=?=8� =�S =N��<&�<6O�<d��<���<��<w"�<�T�<2��<T��<Q��<�<�?�<�j�<f��<���<p��<��<0,�<N�<)n�<|��<��<X��<���<4��<m�<q�<&(�<�5�<~@�<�H�<�N�<$R�<�R�<{P�<pK�<�C�<�8�<�*�<��<M�<���<��<���<p��<sn�<�E�<��<H��<���<��<DE�<��<���<�~�<�4�<���<f��<�?�<���<���<�(�<�ÿ<V[�<��<�~�<�<z��<D�<u��<�<E��<��<L{�<I�<	X�<���<(�<���<�<�I�<���<���<�R�<���<r��<�D�<��<4ۖ<X#�<�i�<���<���<�1�<iq�<���<��<i(�<c�<㜃<�Ձ<��<�|<��x<fu<��q<�>n<��j<wg<��c<'�_<\\\<��X<�9U<+�Q<KN<��J<�G<�}C<��?<�t<<;�8<�v5<��1<�.<�+<��'<58$<� <�n<�<r�<Vc<R<��<��	<�H<!<���;�c�;@�;���;��;��;ap�;<i�;Ap�;��;]��;�ݼ;7 �;�q�;�ҫ;OC�;wà;S�;b�;���;`�;�.�;��;��w;��m;d;@Z;��P;6G;�=;N4;B+;W";�;�.;�l;ċ�:�r�:���:#��:`\�:$�:��:���:�qt:�BU:lj6:Q�:�^�9p��94�x9�9FYv70KǸϤU��Q���T۹�o	���$��N@�l[��Wv�����Ε�K����������ʺ
�ֺ��@u�!��O��'��g������$�G0*��U0��v6���<��B�C�H�%�N���T���Z�Ua��g�/m�Qs��$y�h,�����a���i���ѥ��몎�����O������Ț��  �  �f==w�=�A=a�=�|===;� =�S =V��< �</O�<d��<���<%��<v"�<�T�<"��<T��<V��<�<�?�<�j�<k��<���<u��<��</,�<N�<$n�<���<��<c��<���<-��<q�<b�<2(�<�5�<�@�<�H�<�N�<'R�<�R�<�P�<iK�<�C�<�8�<�*�<��<J�<���<��<���<n��<}n�<F�<��<I��<��<��<CE�<��<���<�~�<�4�<���<q��<�?�<���<���<�(�<�ÿ<W[�<�<�~�<�<v��<>�<���<�<M��<��<R{�<H�<X�<���<(�<���<�<�I�<���<���<�R�<���<s��<�D�<(��<9ۖ<W#�<�i�<�<���<�1�<oq�<���<��<f(�<c�<휃<�Ձ<��<�|<��x<fu<��q<�>n<y�j<�g<��c<2�_<i\\<��X<�9U<'�Q<VN<�J<�G<�}C<��?<�t<<4�8<�v5<��1<�.<�+<w�'<58$< � <�n<�<r�<8c<S<��<��	<�H<<Ļ�;�c�;P�;��;��;��;Mp�;Zi�;Bp�;��;R��;�ݼ;G �;�q�;ӫ;ZC�;�à;S�;n�;���;�_�;�.�;m�;��w;��m;*d;&@Z;q�P;yG;u�=;N4;1+;�";Q;v.;�l;Ɗ�:/s�:��:M��:�\�:�:��:9��:^st:dBU:�j6:��:#^�9k��9ݿx9n�9a�u7�IǸy�U�qS��MQ۹�o	��$�KO@�Bk[��Wv�ʈ���͕�����������ʺ�ֺǸ�u�"��L��$'�^g�k����3$��0*�|U0��v6���<�'�B�+�H�:�N���T���Z�xa�dg�>m�<s��$y�B,���������D�������ժ������J���ﾗ�Ț��  �  �f=!=p�=�A=f�=�|===9� =�S =K��<&�<-O�<c��<���<��<�"�<�T�<&��<V��<Q��<�<�?�<�j�<i��<���<j��<��<2,�<N�<3n�<|��<ߨ�<\��<���<1��<m�<l�<((�<�5�<w@�<�H�<�N�<R�<�R�<tP�<tK�<�C�<�8�<�*�<��<Q�<���<��<���<q��<vn�<�E�<��<E��<���<��<FE�<��<���<�~�<�4�<���<a��<@�<���<���<�(�<�ÿ<X[�<��<�~�<�<y��<G�<y��<�<B��<��<K{�<H�<
X�<���<&(�<���<�<�I�<���<���<�R�<���<o��<�D�<��<<ۖ<W#�<�i�<���<���<�1�<mq�<���<��<o(�<c�<ܜ�<�Ձ<��<��|<��x<fu<��q<�>n<��j<}g<��c<,�_<h\\<{�X<�9U<B�Q<@N<�J<�G<�}C<��?<�t<<4�8<�v5<��1<ޅ.<�+<s�'<48$<.� <�n<�<i�<?c<W<��<φ	<}H<<���;�c�;'�;���;��;߅�;�p�;8i�;6p�;���;l��;�ݼ;7 �;�q�;�ҫ;\C�;]à;S�;v�;l��;!`�;f.�;��;��w;��m;d;:@Z;��P;*G;ٝ=;�M4;H+;o";�;�.;�l;���:�r�:��:���:b\�:�:�:��:Rqt:CU:�i6:��:q_�9Ғ�9`�x9��9M=v7$KǸ'�U�4Q���S۹�o	�\�$��M@� l[��Wv������Ε�����������!ʺy�ֺ��u�!��j���&��g�Q����P$�Z0*��U0��v6���<�-�B�(�H���N���T��Z�a��g��m�Vs�%y�5,�����x���\���륋�⪎�����c�������ǚ��  �  �f=&=o�=�A=b�=�|=C=3� =�S =G��<+�<-O�<^��<���<��<�"�<�T�<,��<V��<L��<�<�?�<�j�<]��<���<k��<��<8,�<
N�<4n�<r��<��<V��<���<3��<d�<v�<(�<�5�<z@�<�H�<�N�<R�<�R�<pP�<{K�<wC�<�8�<�*�<��<Q�<���<��<��<u��<un�<�E�<��<:��<��<��<EE�<��<���<�~�<�4�<���<^��<	@�<���<���<�(�<�ÿ<d[�<��<�~�<�
�<w��<H�<p��<(�<:��<��<C{�<L�<X�<���<((�<���<(�<�I�<���<���<�R�<���<f��<�D�<��<>ۖ<V#�<�i�<���<���<�1�<aq�<���<��<b(�<$c�<؜�<�Ձ<��<��|<��x<fu<��q<�>n<��j<_g<��c<�_<f\\<��X<�9U<G�Q<-N<�J<�G<�}C<��?<�t<<N�8<�v5<��1<օ.<�+<s�'<)8$<2� <zn<�<X�<Kc<U<��<ʆ	<kH<9<���;�c�;+�;���;0��;���;�p�;i�;lp�;݅�;`��;�ݼ; �;�q�;�ҫ;�C�;eà;S�;m�;X��;F`�;U.�;��;*�w;��m;d;�?Z;��P;�
G;�=;�M4;j+;k";�;�.;Ql;��:?r�:���:���:-\�:��:2�:t��:�pt:DU:�i6:
�:D_�9i��9��x9�~9�~v7�QǸ.�U�Q���U۹�m	�P�$��M@�m[�OWv�ǈ���Ε�����������ʺ��ֺ0��Gu� !������&�	h�@�� ��s$�*0*��U0��v6���<�ݬB�6�H�]�N���T�.�Z�� a�	g��m��s��$y�*,�֙��P�������ɥ����������;���$����ǚ��  �  �f==r�=�A=`�=�|=?=9� =�S =P��< �<0O�<d��<���<��<{"�<�T�<)��<O��<Q��<�<�?�<�j�<b��<���<y��<��<0,�<N�<4n�<w��<��<[��<���<2��<i�<p�<((�<�5�<~@�<�H�<�N�<R�<�R�<P�<xK�<wC�<�8�<�*�<��<O�<���<��<���<s��<yn�<�E�<��<D��<��<��<DE�<��<���<�~�<�4�<���<m��<�?�<���<���<�(�<�ÿ<\[�<��<�~�<�<w��<E�<x��<�<@��<��<N{�<J�<X�<���<!(�<���<�<�I�<���<���<�R�<���<p��<�D�<��<:ۖ<[#�<�i�<�<���<�1�<kq�<���<��<_(�<&c�<✃<�Ձ<��<��|<��x<fu<��q<�>n<��j<jg<��c<+�_<b\\<��X<�9U<G�Q<BN<��J<�G<�}C<��?<�t<<=�8<�v5<��1<�.<�+<x�'<58$<#� <�n<�<l�<Dc<I<��<Ɔ	<}H<'<���;�c�;b�;���;��;��;�p�;'i�;Np�;��;^��;�ݼ;% �;�q�;�ҫ;eC�;wà;S�;��;n��;`�;�.�;��;+�w;��m; d;(@Z;��P;,G;��=;�M4;W+;�";;�.;�l;6��:tr�:���:d��:@\�:,�:O�:��:�rt:�BU:j6:	�:�_�9(��9l�x9�9�Sv7�NǸl�U��Q���S۹�n	���$��M@��k[��Wv�∈��͕�$���/�����$ʺ��ֺ��}u�!��d���&��g�`�����I$��0*��U0��v6���<��B�8�H�q�N�w�T���Z�1a��g��m�cs��$y�P,�����c�������ե��㪎�����N�������ǚ��  �  �f==s�=�A=b�=�|=:=>� =�S =W��<%�<1O�<e��<���<��<s"�<�T�<'��<Z��<S��<�<�?�<�j�<s��<���<s��<��<2,�<N�<*n�<���<ݨ�<_��<���<1��<w�<h�<,(�<5�<�@�<�H�<�N�<%R�<�R�<P�<iK�<�C�<�8�<�*�<��<D�<���<��<��<i��<xn�<�E�<��<P��<��<��<=E�<��<���<�~�<�4�<���<k��<�?�<���<���<�(�<�ÿ<Q[�<�<�~�<�<{��<B�<|��<�<K��<��<L{�<L�<X�<���<(�<���<�<�I�<���<���<�R�<���<y��<�D�<"��<6ۖ<W#�<�i�<���<���<�1�<uq�<���<��<h(�<c�<圃<�Ձ<��<�|<��x<fu<��q<�>n<~�j<�g<��c<.�_<b\\<{�X<�9U<.�Q<KN<��J<�G<�}C<��?<�t<<)�8<�v5<��1<��.<�+<|�'<78$<� <�n<~<z�<@c<_<��<��	<�H<<��;�c�;I�;���;��;��;ap�;Vi�;.p�;��;[��;�ݼ;_ �;�q�;�ҫ;=C�;�à; S�;`�;���;`�;�.�;l�;��w;��m;d;X@Z;B�P;�G;��=;JN4;	+;|";;E.;�l;#��:Ns�:���:���:�\�:��:N�:9��:�rt:�BU:�j6:S�:�_�9Ε�9��x9%�9}v7�BǸ$�U�cR���R۹<p	�@�$��N@�l[�hWv�툈�!Ε�����	��[���ʺ��ֺ
�㺻t�!����I'��g������$�k0*�rU0�	w6�^�<�>�B���H�*�N���T���Z�;a��g�3m�(s��$y�`,���������3�������ݪ������c����Ț��  �  �f= =r�=�A=b�=�|=<=;� =�S =Q��<%�<+O�<a��<���<��<�"�<�T�<#��<V��<R��<�<�?�<�j�<h��<���<u��<��<5,�<N�<-n�<x��<��<b��<���<+��<h�<j�<+(�<�5�<{@�<�H�<�N�< R�<�R�<}P�<qK�<{C�<�8�<�*�<��<J�<���<��<��<q��<yn�<�E�<��<B��<��<��<AE�<��<���<�~�<�4�<���<j��<@�<���<���<�(�<�ÿ<a[�<�<�~�< �<s��<D�<}��<"�<B��<��<H{�<L�<	X�<���<(�<���<�<�I�<���<���<�R�<���<m��<�D�<��<=ۖ<W#�<�i�<���<���<�1�<nq�<���<��<e(�< c�<���<�Ձ<��<�|<��x<fu<��q<�>n<��j<sg<��c<.�_<u\\<��X<�9U<5�Q<AN<�J<�G<�}C<��?<�t<<1�8<�v5<��1<�.<�+<n�'</8$</� <�n<�<d�<8c<V<��<��	<�H<<���;�c�;P�;���;$��;ԅ�;mp�;*i�;\p�;��;`��;�ݼ;! �;�q�;�ҫ;�C�;mà;S�;a�;v��;`�;�.�;��;G�w;��m;d;)@Z;o�P;MG;��=;�M4;I+;�";;�.;�l;��:�r�:Ǎ�:@��:y\�:�:��:���:vrt:CU:j6:�:�_�9��9��x9}�9�0v7�PǸB�U��Q���R۹cn	�]�$�5N@��l[�ZWv����Ε�g���������ʺ�ֺ���u��!��z���&��g�E����d$�p0*��U0��v6���<�*�B�$�H�?�N���T���Z�'a��g�m�Zs��$y��+���������q�������ު������P���	����ǚ��  �  �f=!=n�=�A=c�=�|=@=4� =�S =N��<'�<9O�<]��<���<��<�"�<�T�<7��<R��<S��<�<�?�<�j�<i��<���<r��<��<7,�<N�<6n�<m��<��<T��<���<4��<e�<x�<(�<�5�<t@�<�H�<�N�<R�<�R�<uP�<wK�<~C�<�8�<�*�<��<W�<���<��<��<r��<nn�<�E�<��<?��<��<��<ME�<��<���<�~�<�4�<���<a��<�?�<���<���<�(�<�ÿ<_[�<��<�~�< �<z��<J�<o��<#�<8��<��<D{�<L�<X�<���<$(�<���<%�<�I�<���<���<�R�<���<g��<�D�<��<9ۖ<V#�<�i�<���<���<�1�<dq�<���<��<i(�<$c�<ל�<�Ձ<��<��|<��x<	fu<��q<�>n<��j<dg<��c<"�_<`\\<��X<�9U<B�Q<9N<�J<�G<�}C<��?<�t<<A�8<�v5<��1<�.<�+<��'<(8$<)� <pn<�<Y�<`c<M<��<Ȇ	<qH<1<���;�c�;E�;���;/��;Ņ�;�p�;�h�;^p�;Յ�;f��;�ݼ; �;r�;�ҫ;lC�;Pà;S�;e�;`��;`�;h.�;��;b�w;�m;d;@Z;ٖP;G;,�=;�M4;O+;/";�;�.;ul;>��:Er�:|��:2��:F\�:��:��:#��:Zqt:�BU:zi6:��:�`�9���9��x9�~9��v7�OǸ̤U�nP��V۹On	���$��L@��l[�RWv�/����Ε��������7��mʺ��ֺ���{u� ������&�0h�g��"��$�70*��U0�zv6��<�
�B���H�"�N���T�1�Z�a��g��m��s�%y�7,�̙��F�������������������T���,����ǚ��  �  �f=#=t�=�A=a�=�|===8� =�S =R��<�<0O�<[��<���<��<�"�<�T�<*��<M��<T��<�<�?�<�j�<l��<���<s��<��<9,�<N�</n�<}��<��<]��<���<)��<c�<m�<)(�<�5�<�@�<�H�<�N�< R�<�R�<�P�<kK�<�C�<�8�<�*�<��<Q�<���<��<��<o��<}n�<�E�<��<@��<���<��<GE�<��<���<�~�<�4�<���<m��<@�<���<���<�(�<�ÿ<a[�< �<�~�<�
�<p��<F�<y��<%�<F��<��<B{�<Q�<X�<���<(�<���<�<�I�<���<���<�R�<���<g��<�D�<��<Aۖ<R#�<�i�<�<���<�1�<jq�<���<��<f(�<c�<䜃<�Ձ<��<�|<��x<fu<��q<�>n<��j<`g<��c<'�_<m\\<��X<�9U<0�Q<<N<�J<�G<�}C<��?<�t<<4�8<�v5<��1<�.<�+<y�'<#8$<6� <�n<�<W�<Gc<D<��<��	<H<<Ļ�;�c�;J�;��;6��;���;xp�;<i�;lp�;���;\��;�ݼ; �;�q�;�ҫ;uC�;�à;"S�;J�;t��;<`�;�.�;t�;s�w;��m;�d;�?Z;��P;G;ɝ=;�M4;;+;�";6;�.;�l;f��:Zr�:#��:	��:3\�:	�:��:i��:�rt:�CU:Yj6:M�:N`�9W��9��x9��9�Av7�TǸ��U��Q���S۹n	���$��M@�9m[��Vv�l���Ε�����������$ʺ�ֺҸ㺘u�~!������&��g�(��@��?$��0*��U0��v6���<�*�B� �H�>�N���T���Z�� a��g�6m�Gs��$y�,�����q�������祋�쪎�����:��������ǚ��  �  �f==b�=uA=U�=�|="=%� =�S =��<��<�N�<��<]��<���<"�<vT�<���<��<���<��<?�<j�<ӓ�<��<���<��<�+�<\M�<jm�<���<��<���<���<K��<��<h�<''�<t4�<[?�<�G�<�M�<�P�<hQ�<CO�<,J�<DB�<17�<T)�<.�<��<v��<���<{��<��<�l�<bD�<K�<���<O��<f~�<�C�<&�<���<�|�<3�<>��<���<9>�<��<��<�&�<5¿<�Y�<W�</}�<q	�<㑸<��<藵<��<���<u�<�y�<��<�V�<H��<�&�<R��<��<�H�<��<���<�Q�<���<x��<�C�<1��<fږ<�"�<�h�<>��<��<1�<�p�<%��<!�<(�<�b�<���<{Ձ<��<��|<��x<�eu<��q<�>n<��j<�g<�c<��_<�\\<�X<v:U<�Q<<N<	�J<�G<�~C<L�?<v<<��8<�x5<F�1<ׇ.<�+<��'<E:$<i� <�p<�<�<�e<<��<��	<�K<
<���;j�;��;b��;��;���;Uw�;p�;(w�;.��;���;+�;�'�;(y�;oګ;�J�;�ʠ;�Z�;��;��;vg�;16�;$�;x;n�m;�d;'OZ;8�P;dG; �=;X\4;)+;/";�;�;;z;��:L��:'��:���:�u�:�#�:��:�:}�t:UkU:6:�:Ϭ�9uݷ9�Py9e9�~7/Ƹ�U����5۹�R	���$�)3@�wQ[��=v��}��g��񢺛������ʺ��ֺj���k�b��@��V#�Xd�˞�$��$��-*��R0��t6���<�֪B�?�H���N��T�6�Z� a�c
g��m��s��$y��+�}���_������ޥ����������ӷ��N���+Ț��  �  �f==f�=wA=K�=�|=#=� =�S =��<��<�N�<��<_��<���<"�<oT�<���<ε�<���<��<�>�<j�<̓�<��<���<��<�+�<OM�<jm�<���<"��<���<���<=��<n�<n�<#'�<�4�<t?�<�G�<�M�<�P�<{Q�<DO�<%J�<0B�<37�<@)�<!�<��<[��<���<w��<��<�l�<mD�<S�<���<O��<K~�<�C�<�<���<�|�<�2�<7��<���<N>�<��<��<'�<H¿<�Y�<R�<1}�<W	�<Б�<��<闵<��<���<x�<�y�<��<�V�<M��<�&�<I��<��<�H�<���<���<kQ�<���<n��<�C�<5��<gږ<�"�<�h�<6��<��<&1�<�p�<"��<!�<�'�<�b�<���<�Ձ<��<��|<��x<
fu<��q<�>n<��j<�g<�c<��_<]\<L�X<�:U<�Q<4N<�J<�G<�~C<'�?<v<<��8<zx5<[�1<.<�+<��'<G:$<n� <�p<�<�<�e<�<��<��	<dK<<���;�i�;��;���;��;���;Uw�;Ap�;�w�;9��;���;��;p'�;@y�;aګ;!K�;3ˠ;�Z�;���;$��;�g�;56�;�;vx;{�m;d;�NZ;%�P;�G;�=;6\4;X)+;�";�;<;�y;��:���:ͦ�:I��:`t�:$$�:��:��:��t:�mU:��6:C:���9`�90\y9�9�~7|HƸ�(U�<��۹xO	�w�$��2@��R[�=v�M|�� �p�0�����Dʺ��ֺկ�dm�-�����9#�4d�Ğ���$��-*�S0�qt6�|�<���B�B�H�h�N��T��Z���`�
g�m�.s��#y�8+�����E���p���᥋��������B���+���EȚ��  �  �f==_�={A=H�=�|=(=� =�S =��<��<�N�<��<X��<���<"�<mT�<ą�<յ�<���<��<�>�<%j�<Γ�<��<���<��<x+�<TM�<wm�<���<��<r��<���<T��<{�<��<'�<y4�<[?�<�G�<�M�<�P�<qQ�<<O�<0J�<-B�<F7�<A)�<$�<��<_��<���<v��<��<�l�<`D�<Y�<���<b��<P~�<�C�<!�<���<�|�<�2�<D��<���<B>�<��<���<'�<1¿<�Y�<F�<D}�<g	�<䑸<��<ח�<��<���<��<�y�<��<�V�<J��<�&�<K��<��<�H�<���<���<rQ�<���<n��<�C�<)��<\ږ<�"�<�h�<A��<��<41�<�p�<,��<+�<�'�<�b�<���<Ձ<��<��|<��x<�eu<s�q<�>n<ڪj<�g<�c<��_<�\\<%�X<p:U<"�Q<>N<�J<�G<�~C<�?<v<<��8<tx5<v�1<ʇ.<�+<��'<M:$<_� <�p<�<�<�e<�<��<��	<ZK<4<���;�i�;��;a��;���;���;�w�;p�;`w�;��;ñ�;L�;�'�;�y�;=ګ;�J�;�ʠ;�Z�;��;��;�g�;6�;3�;ax;�m;d;�NZ;v�P;�G;u�=;4\4;t)+;&";};-<;�y;?��:��:o��:���:.t�:8%�:|�:p�:t:wlU:��6::d��9mܷ9=Uy9�9wc7A9Ƹ�U�_���۹�Q	���$�v1@�
R[��>v�J}��L�/�������ʺ�ֺ0���l�`�����#��d������$��-*��R0�t6�z�<���B���H���N���T�l�Z���`�m
g��m�ls�U$y��+���������W�������򪎻��������Y���$Ț��  �  �f==d�=xA=J�=�|= =!� =�S =��<��<�N�<��<^��<���<"�<rT�<���<ݵ�<���<��<?�<j�<Г�<��<���<��<�+�<VM�<om�<���<��<���<���<?��<t�<i�<''�<�4�<g?�<�G�<�M�<�P�<|Q�<FO�<-J�</B�<77�<=)�<)�<��<i��<���<n��<��<�l�<oD�<U�<���<K��<X~�<�C�<"�<���<�|�<�2�<?��<���<O>�<��<��<	'�<@¿<�Y�<W�<.}�<[	�<ӑ�<��<뗵<��<ď�<|�<�y�<��<�V�<Q��<�&�<M��<��<�H�<���<���<zQ�<���<o��<�C�<=��<gږ<�"�<�h�<=��<	��< 1�<�p�<��<#�<�'�<�b�<���<�Ձ<��<��|<��x<�eu<��q<�>n<��j<�g<ނc<��_< ]\<+�X<�:U<�Q<<N<�J<�G<�~C<!�?<v<<��8<�x5<O�1<Ƈ.<�+<g�'<Q:$<l� <�p<<�<�e<�<|�<��	<|K<	<���;�i�;��;���;��;���;iw�;Wp�;nw�;5��;���;��;�'�;,y�;sګ;K�;ˠ;�Z�;���;��;�g�;<6�;'�;rx;��m;�d;�NZ;�P;�G;�=;�[4;d)+;�";�;<;�y;Ӥ�:v��:o��:���:Jt�:*$�:��:+�:�t:nU:L�6:�:���9q�9Zy9�9�~7�DƸ�&U�X���۹Q	��$�62@��Q[��<v�T|������2��������ʺ��ֺ��sl������#��c��������$��-*��R0��t6��<��B�.�H�~�N���T��Z���`�h
g��m��s�4$y�a+�f���l���[�������ߪ�������������>Ț��  �  �f==d�=sA=M�=�|=="� =�S =��<��<�N�<��<H��<���<"�<�T�<���<��<���<��<
?�<j�<���<��<���<��<�+�<MM�<`m�<���<��<���<���<A��<��<l�<*'�<r4�<h?�<�G�<�M�<�P�<wQ�<?O�<!J�<?B�<A7�<9)�<-�<��<m��<���<���<��<�l�<_D�<I�<���<M��<^~�<�C�<$�<���<�|�<3�<4��<���<H>�<
��<��<'�<A¿<�Y�<Y�<.}�<g	�<ّ�<��<뗵<��<Ǐ�<r�<�y�<��<�V�<C��<�&�<`��<��<�H�<���<���<�Q�<���<���<�C�<-��<Rږ<�"�<�h�<>��<��<$1�<�p�<��<0�<(�<�b�<���<�Ձ<��<��|<��x<�eu<��q<�>n<��j<�g<�c<��_<�\\<$�X<�:U<��Q<1N<�J<�G<�~C<.�?<.v<<��8<�x5<X�1<͇.<�+<��'<d:$<?� <�p<�<
�<�e<<��<��	<{K<<��;�i�;��;���;ү�;���;-w�;[p�;6w�;/��;���;�;�'�;:y�;~ګ;�J�;ˠ;�Z�;���;��;�g�;!6�;��;�x;��m;�d;!OZ;�P;G;��=;�\4;)+;";u;�;;dz;��:،�:���:���:)t�:�$�:��:q�:ҝt:DmU:K�6::���9��9�Oy9�9ȵ~79Ƹ�#U���x۹�R	���$�3@�0S[��=v��|�������
������ʺ��ֺ���l�m������#�rd�k������$��-*��R0��t6���<�]�B���H�&�N�M�T�9�Z���`��
g�Mm�,s�F$y��+�e���V������񥋻�̰������!���qȚ��  �  �f==_�={A=J�=�|=%=� =�S =	��<��<�N�<��<Y��<���<"�<qT�<���<ӵ�<���<��<�>�< j�<͓�<��<���<��<{+�<[M�<qm�<���<��<���<���<G��<j�<v�<('�<4�<c?�<�G�<�M�<�P�<wQ�<AO�</J�<*B�<E7�<;)�<#�<��<c��<���<t��<��<�l�<kD�<X�<���<N��<S~�<�C�<�<���<�|�<�2�<B��<���<H>�<	��<���<'�<9¿<�Y�<V�<9}�<W	�<ّ�<��<藵<��<���<~�<�y�<��<�V�<K��<�&�<J��<��<�H�<���<���<sQ�<���<q��<�C�<?��<`ږ<�"�<�h�<8��<��<11�<�p�<#��<,�<�'�<�b�<���<�Ձ<��<��|<��x<�eu<��q<�>n<��j<�g<��c<��_<�\\<5�X<g:U<)�Q<@N<�J<�G<�~C<�?<v<<��8<jx5<q�1<��.<�+<z�'<P:$<b� <�p<�<�<�e<�<��<��	<QK<+<���;�i�;��;s��;���;���;sw�;p�;hw�;'��;���;�;`'�;^y�;uګ;�J�;�ʠ;�Z�; ��;��;�g�;(6�;/�;Jx;�m;�d;�NZ;g�P;�G;�=;$\4;U)+;a";�;%<;�y;��:&��:X��:���:�s�:%�:X�:R�:J�t:=mU:)�6:N:���9�޷9Wy99J7�HƸ$U�v��f۹YQ	���$��1@�IQ[��>v��|��4��������ʺ)�ֺg���l���w��#��c�������A$��-*�#S0�t6���<��B���H���N���T�y�Z���`�U
g��m��s�$y�~+�k���+�������å��᪎�Ȱ��o���l���Ț��  �  �f==_�=xA=M�=�|=+=� =�S =��<��<�N�<��<b��<���<""�<eT�<���<��<���<��<�>�<*j�<Ɠ�<��<���<��<�+�<KM�<mm�<���<&��<{��<���<I��<n�<y�<'�<�4�<k?�<�G�<�M�<�P�<�Q�<3O�<1J�<)B�<G7�<C)�< �<��<^��<���<j��<��<�l�<bD�<X�<���<f��<R~�<�C�<�<���<�|�<�2�<D��<���<Y>�<��<��<'�<?¿<�Y�<D�<;}�<Y	�<ۑ�<��<ܗ�<��<���<{�<�y�<��<�V�<A��<�&�<B��<��<�H�<���<���<}Q�<���<c��<�C�<*��<fږ<�"�<�h�<V��<��<01�<�p�<0��<&�<�'�<�b�<���<�Ձ<��<��|<��x<fu<��q<�>n<Ϫj<�g<
�c<��_<�\\<N�X<m:U<"�Q<N<0�J<�G<�~C<,�?<v<<��8<bx5<s�1<��.<�+<}�'<C:$<t� <�p<<Ϲ<�e<<x�<��	<NK<><���;�i�;��;���;���;v��;bw�;p�;�w�;��;���;!�;n'�;ly�;(ګ; K�;ˠ;�Z�;��;稐;�g�;�5�;6�;Cx;�m;#d;�NZ;P�P;�G;��=;�[4;r)+;U";�;'<;ky;w��:��:!��:���:\t�:q%�:�:��:^�t:YoU:�6:�:���9�9�]y9�9�7�FƸ #U�M��d۹<O	�d�$�\2@�S[�Z=v�|�����񢺟��_���ʺ�ֺ���<l�������"��d�Ϟ�
��[$��,*�:S0�$t6���<���B��H�k�N���T���Z�>�`��
g��m��s��#y�T+�������������������°��=���`���$Ț��  �  �f==c�=tA=Q�=�|="=� =�S =��<��<�N�<��<]��<���<"�<sT�<���<ݵ�<���<��<?�<j�<̓�<��<���<��<}+�<PM�<om�<���<��<���<���<E��<��<w�<%'�<v4�<c?�<�G�<�M�<�P�<�Q�<;O�<+J�<6B�<77�<<)�<+�<��<[��<���<x��<��<�l�<`D�<W�<���<W��<M~�<�C�<&�<���<�|�<�2�<A��<���<S>�<��<��<	'�<=¿<�Y�<T�<;}�<f	�<ڑ�<��<嗵<��<���<~�<�y�<��<�V�<@��<�&�<N��<��<�H�<���<���<uQ�<���<u��<�C�<%��<bږ<�"�<�h�<B��<��<41�<�p�<!��< �<(�<�b�<���<�Ձ<��<��|<��x<�eu<~�q<�>n<��j<�g<�c<��_<�\\<�X<|:U< �Q<"N<�J<�G<�~C<=�?<
v<<��8<�x5<y�1<��.<�+<|�'<\:$<i� <�p<<�<�e<�<l�<��	<oK<<���;�i�;��;���;¯�;���;mw�;,p�;@w�;"��;���;�;�'�;dy�;kګ;�J�;�ʠ;�Z�;��;ި�;�g�;6�;�;�x;��m;�d;OZ;[�P;�G;:�=;?\4;{)+;?";;!<;�y;���:���:��:���:+t�:i$�:��:E�:>�t:�nU:Q�6:�:���9�߷9�Ry9�9�7�9ƸO#U����,۹�R	���$��1@�iR[��>v�|���������{��#ʺ��ֺF�㺻l���]��#��d������A$�}-*�CS0�t6�+�<���B�M�H��N�&�T�W�Z���`��
g��m�6s�|$y��+�s���>���!���ӥ��񪎻԰������A���)Ț��  �  �f=
=i�=vA=I�=�|=%=� =�S =��<��<�N�<��<Q��<���<"�<uT�<���<ٵ�<���<��<?�<j�<ғ�<��<���<��<q+�<aM�<bm�<���<��<���<���<9��<q�<a�<5'�<w4�<o?�<�G�<�M�<�P�<tQ�<RO�<!J�<.B�<:7�<@)�<�<��<k��<���<|��<��<�l�<lD�<M�<���<I��<X~�<�C�<�<���<�|�<�2�<4��<ē�<I>�<��<��<�&�<I¿<�Y�<d�<)}�<Y	�<ϑ�<��<���<��<Ǐ�<o�<�y�<��<�V�<R��<�&�<N��<��<�H�<x��<���<xQ�<���<w��<�C�<A��<Zږ<�"�<�h�<7��<��<!1�<�p�<'��<)�<�'�<�b�<���<wՁ<��<��|<��x<�eu<��q<�>n<��j<�g<̂c<��_<]\<.�X<�:U<�Q<SN<�J<�G<�~C<�?<v<<��8<vx5<N�1<҇.<�+<~�'<P:$<Q� <�p<�<�<�e<�<��<�	<gK<<���;�i�;��;���;���;ь�;6w�;Rp�;Sw�;Z��;���;��;{'�;y�;�ګ;�J�;!ˠ;�Z�;���;��;�g�;k6�;��;ix;��m;
d;�NZ;�P;G;ҫ=;a\4;%)+;_";�;�;;z;���:p��:̦�:���:@t�:|$�:��:v�:�t:jmU:]�6:�:c��9��9BRy99��~7GƸ�(U�����۹dR	���$��3@��P[�'?v�;|��������������ʺ=�ֺ��㺓l����I��[#��c�*�����6$��-*��R0��t6���<�ʪB��H�|�N�,�T���Z�) a�
g�(m�Ls�$y��+�5�������k���"�����������|���*���ZȚ��  �  �f==a�=tA=N�=�|='=� =�S =��<��<�N�<��<O��<���<"�<sT�<���<ڵ�<���<��<?�<j�<ٓ�<��<���<��<z+�<]M�<_m�<���<��<w��<���<M��<��<u�< '�<o4�<j?�<�G�<�M�<�P�<pQ�<>O�<(J�<<B�<A7�<H)�<&�<��<g��<���<{��<��<�l�<aD�<M�<���<]��<V~�<�C�<!�<���<�|�<�2�<?��<���<B>�<��<��<�&�<B¿<�Y�<M�<7}�<h	�<䑸<��<ޗ�<��<ŏ�<n�<�y�<��<�V�<D��<�&�<U��<��<�H�<���<���<xQ�<���<t��<�C�<1��<Yږ<�"�<�h�<C��<��<11�<�p�<-��<+�<(�<�b�<���<{Ձ<��<��|<��x<�eu<o�q<�>n<��j<�g<��c<��_<�\\<*�X<:U<��Q<RN<��J<�G<�~C<3�?<v<<��8<�x5<k�1<ه.<�+<��'<Z:$<N� <�p<�<�<�e<�<��<��	<kK<#<���;�i�;��;���;���;���;+w�;Np�;Pw�;���;���;3�;�'�;_y�;Vګ;�J�;ˠ;�Z�;���;��;�g�;6�;�;�x;��m;Md;�NZ;U�P;�G;Y�=;Y\4;7)+;$";�;�;;z;��:X��:J��:���:�t�:�$�:G�:!�:��t:{lU:q�6:�:3��9��9?Py9�9��~7R7Ƹ�U�H���۹mR	���$��3@�oQ[��>v��|������r��3���ʺ��ֺ'�㺒l���`���#�Ud�2����� $�s-*��R0�t6�e�<���B���H�"�N��T�J�Z� a�
g�Bm�ms�$y��+�p���+���*���å��𪎻��������;���mȚ��  �  �f==b�=rA=Q�=�|=!=� =�S =��<��<�N�<��<h��<���<)"�<jT�<���<յ�<���<��< ?�<j�<̓�<��<���<��<�+�<SM�<rm�<���<��<���<���<@��<m�<v�<!'�<�4�<c?�<�G�<�M�<�P�<�Q�<<O�<*J�<3B�<27�<<)�<'�<��<S��<���<f��<���<�l�<nD�<`�<���<T��<E~�<�C�<$�<���<�|�<�2�<A��<���<U>�<��<��<
'�<;¿<�Y�<Q�<;}�<X	�<ӑ�<��<藵<��<���<��<�y�<��<�V�<B��<�&�<J��<��<�H�<���<���<mQ�<���<h��<�C�<7��<oږ<�"�<�h�<?��<��<91�<�p�<��<�<(�<�b�<���<�Ձ<��<��|<��x<�eu<��q<�>n<��j<�g<�c<��_<]\<�X<�:U<$�Q<,N<&�J<�G<�~C<=�?<v<<��8<�x5<y�1<��.<�+<e�'<V:$<�� <�p<<ڹ<�e<�<��<��	<gK<<���;�i�;��;���;��;���;vw�;:p�;lw�;8��;���;��;j'�;by�;Zګ;+K�;�ʠ;�Z�;��;�;�g�;6�;�;�x;v�m;�d;�NZ;q�P;NG;&�=;�[4;�)+;�";�;h<;py;V��:I��:+��:���:\t�:$�:��:R�:u�t:�nU:��6:�:���9߷9�\y9�9�7RHƸ�&U����^۹�P	��$��1@�YR[��=v�|������!�����-ʺ�ֺϯ�Am�������"�'d��������$��-*�cS0��s6�l�<��B�f�H��N�<�T�[�Z�i�`��
g��m�s�d$y�3+�����:���q���ӥ��������������'���"Ț��  �  �f==`�=uA=N�=�|='=� =�S =��<��<�N�<	��<T��<���<"�<nT�<Å�<��<���<��<?�<j�<ؓ�<
��<���<��<}+�<RM�<dm�<���<��<���<���<K��<z�<p�<!'�<{4�<[?�<�G�<�M�<�P�<uQ�<;O�<%J�<7B�<A7�<H)�< �<��<g��<���<w��<��<�l�<^D�<O�<���<b��<\~�<�C�<�<���<�|�<�2�<7��<���<D>�<��<��<�&�<5¿<�Y�<O�<5}�<e	�<ޑ�<��<藵<��<���<u�<�y�<��<�V�<E��<�&�<T��<��<�H�<���<���<�Q�<���<p��<�C�<+��<Xږ<�"�<�h�<Q��<��<,1�<�p�<-��<+�<(�<�b�<���<�Ձ<��<��|<��x<�eu<��q<�>n<��j<�g<��c<��_<]\<�X<:U<	�Q<2N<�J<�G<�~C</�?<"v<<��8<yx5<f�1<ɇ.<�+<��'<J:$<W� <�p<�<�<�e<<��<��	<hK<#<���;�i�;��;q��;ï�;���;Aw�;'p�;8w�;5��;���;+�;�'�;Iy�;Xګ;�J�;�ʠ;�Z�;���;��;�g�;6�;�;�x;��m;Kd;�NZ;B�P;�G;��=;<\4;>)+;";m;�;;�y;9��:���:��:w��:�t�:�$�:�:��:{�t:�lU:{�6:�:��9�ݷ9mSy9�9�~7�:Ƹ(!U����N۹�R	���$�3@��R[�>v�.}����^򢺅��N���ʺz�ֺ��㺽k�{�����Q#��d�>�����
$�-*��R0�Ct6���<���B���H�,�N�$�T�f�Z���`��
g�m�Is��$y�]+�y���5���R������������������<���WȚ��  �  �f==a�=~A=L�=�|=#=� =�S =	��<��<�N�<��<Y��<���<"�<pT�<���<̵�<���<��<?�<j�<ԓ�<��<���<��<�+�<aM�<am�<���<��<���<���<J��<u�<l�<+'�<y4�<t?�<�G�<�M�<Q�<oQ�<DO�<.J�<3B�<,7�<A)�<(�<��<Z��<���<y��<��<�l�<wD�<N�<���<J��<K~�<�C�<#�<���<�|�<�2�<>��<���<@>�<$��<��<'�<P¿<�Y�<X�<.}�<]	�<ב�<��<ꗵ<��<я�<v�<�y�<��<�V�<Z��<�&�<R��<��<�H�<���<���<jQ�<���<s��<�C�<E��<cږ<�"�<�h�<0��< ��<.1�<�p�<(��<�<�'�<�b�<���<{Ձ<��<��|<��x<�eu<��q<�>n<��j<�g<��c<��_<�\\<2�X<�:U<��Q<`N<�J<�G<�~C<(�?<v<<��8<�x5<r�1<��.<�+<��'<Q:$<a� <�p<�<�<�e<�<z�<��	<nK<<���;�i�;��;s��;߯�;Ќ�;1w�;tp�;Mw�;1��;���;$�;�'�;8y�;�ګ;�J�;4ˠ;�Z�;���;f��;�g�;56�;*�;�x;F�m;d;�NZ;#�P;�G;۫=;G\4;K)+;�";6;�;;�y;���:���:���:���:qt�:�#�:��:�:Q�t:MlU:y�6:�:��9a�9Sy909{�~7RCƸ�$U�r���۹lR	�v�$��2@��P[�<v�0}��R���򢺚��Z���ʺ)�ֺ5��{m���o���#��c�������-$�.*�'S0�1t6�9�<���B�Z�H�P�N���T�A�Z� a��	g�Tm�s�$y��+�m���G���s���ͥ���������t������|Ț��  �  �f==`�=uA=N�=�|='=� =�S =��<��<�N�<	��<T��<���<"�<nT�<Å�<��<���<��<?�<j�<ؓ�<
��<���<��<}+�<RM�<dm�<���<��<���<���<K��<z�<p�<!'�<{4�<[?�<�G�<�M�<�P�<uQ�<;O�<%J�<7B�<A7�<H)�< �<��<g��<���<w��<��<�l�<^D�<O�<���<b��<\~�<�C�<�<���<�|�<�2�<7��<���<D>�<��<��<�&�<5¿<�Y�<O�<5}�<e	�<ޑ�<��<藵<��<���<u�<�y�<��<�V�<E��<�&�<T��<��<�H�<���<���<�Q�<���<p��<�C�<+��<Xږ<�"�<�h�<Q��<��<,1�<�p�<-��<+�<(�<�b�<���<�Ձ<��<��|<��x<�eu<��q<�>n<��j<�g<��c<��_<]\<�X<:U<	�Q<2N<�J<�G<�~C</�?<"v<<��8<yx5<f�1<ɇ.<�+<��'<J:$<W� <�p<�<�<�e<<��<��	<hK<#<���;�i�;��;q��;ï�;���;Aw�;'p�;8w�;5��;���;+�;�'�;Iy�;Xګ;�J�;�ʠ;�Z�;���;��;�g�;6�;�;�x;��m;Kd;�NZ;B�P;�G;��=;<\4;>)+;";m;�;;�y;9��:���:��:w��:�t�:�$�:�:��:{�t:�lU:{�6:�:��9�ݷ9mSy9�9�~7�:Ƹ(!U����N۹�R	���$�3@��R[�>v�.}����^򢺅��N���ʺz�ֺ��㺽k�{�����Q#��d�>�����
$�-*��R0�Ct6���<���B���H�,�N�$�T�f�Z���`��
g�m�Is��$y�]+�y���5���R������������������<���WȚ��  �  �f==b�=rA=Q�=�|=!=� =�S =��<��<�N�<��<h��<���<)"�<jT�<���<յ�<���<��< ?�<j�<̓�<��<���<��<�+�<SM�<rm�<���<��<���<���<@��<m�<v�<!'�<�4�<c?�<�G�<�M�<�P�<�Q�<<O�<*J�<3B�<27�<<)�<'�<��<S��<���<f��<���<�l�<nD�<`�<���<T��<E~�<�C�<$�<���<�|�<�2�<A��<���<U>�<��<��<
'�<;¿<�Y�<Q�<;}�<X	�<ӑ�<��<藵<��<���<��<�y�<��<�V�<B��<�&�<J��<��<�H�<���<���<mQ�<���<h��<�C�<7��<oږ<�"�<�h�<?��<��<91�<�p�<��<�<(�<�b�<���<�Ձ<��<��|<��x<�eu<��q<�>n<��j<�g<�c<��_<]\<�X<�:U<$�Q<,N<&�J<�G<�~C<=�?<v<<��8<�x5<y�1<��.<�+<e�'<V:$<�� <�p<<ڹ<�e<�<��<��	<gK<<���;�i�;��;���;��;���;vw�;:p�;lw�;8��;���;��;j'�;by�;Zګ;+K�;�ʠ;�Z�;��;�;�g�;6�;�;�x;v�m;�d;�NZ;q�P;NG;&�=;�[4;�)+;�";�;h<;py;V��:I��:+��:���:\t�:$�:��:R�:u�t:�nU:��6:�:���9߷9�\y9�9�7RHƸ�&U����^۹�P	��$��1@�YR[��=v�|������!�����-ʺ�ֺϯ�Am�������"�'d��������$��-*�cS0��s6�l�<��B�f�H��N�<�T�[�Z�i�`��
g��m�s�d$y�3+�����:���q���ӥ��������������'���"Ț��  �  �f==a�=tA=N�=�|='=� =�S =��<��<�N�<��<O��<���<"�<sT�<���<ڵ�<���<��<?�<j�<ٓ�<��<���<��<z+�<]M�<_m�<���<��<w��<���<M��<��<u�< '�<o4�<j?�<�G�<�M�<�P�<pQ�<>O�<(J�<<B�<A7�<H)�<&�<��<g��<���<{��<��<�l�<aD�<M�<���<]��<V~�<�C�<!�<���<�|�<�2�<?��<���<B>�<��<��<�&�<B¿<�Y�<M�<7}�<h	�<䑸<��<ޗ�<��<ŏ�<n�<�y�<��<�V�<D��<�&�<U��<��<�H�<���<���<xQ�<���<t��<�C�<1��<Yږ<�"�<�h�<C��<��<11�<�p�<-��<+�<(�<�b�<���<{Ձ<��<��|<��x<�eu<o�q<�>n<��j<�g<��c<��_<�\\<*�X<:U<��Q<RN<��J<�G<�~C<3�?<v<<��8<�x5<k�1<ه.<�+<��'<Z:$<N� <�p<�<�<�e<�<��<��	<kK<#<���;�i�;��;���;���;���;+w�;Np�;Pw�;���;���;3�;�'�;_y�;Vګ;�J�;ˠ;�Z�;���;��;�g�;6�;�;�x;��m;Md;�NZ;U�P;�G;Y�=;Y\4;7)+;$";�;�;;z;��:X��:J��:���:�t�:�$�:G�:!�:��t:{lU:q�6:�:3��9��9?Py9�9��~7R7Ƹ�U�H���۹mR	���$��3@�oQ[��>v��|������r��3���ʺ��ֺ'�㺒l���`���#�Ud�2����� $�s-*��R0�t6�e�<���B���H�"�N��T�J�Z� a�
g�Bm�ms�$y��+�p���+���*���å��𪎻��������;���mȚ��  �  �f=
=i�=vA=I�=�|=%=� =�S =��<��<�N�<��<Q��<���<"�<uT�<���<ٵ�<���<��<?�<j�<ғ�<��<���<��<q+�<aM�<bm�<���<��<���<���<9��<q�<a�<5'�<w4�<o?�<�G�<�M�<�P�<tQ�<RO�<!J�<.B�<:7�<@)�<�<��<k��<���<|��<��<�l�<lD�<M�<���<I��<X~�<�C�<�<���<�|�<�2�<4��<ē�<I>�<��<��<�&�<I¿<�Y�<d�<)}�<Y	�<ϑ�<��<���<��<Ǐ�<o�<�y�<��<�V�<R��<�&�<N��<��<�H�<x��<���<xQ�<���<w��<�C�<A��<Zږ<�"�<�h�<7��<��<!1�<�p�<'��<)�<�'�<�b�<���<wՁ<��<��|<��x<�eu<��q<�>n<��j<�g<̂c<��_<]\<.�X<�:U<�Q<SN<�J<�G<�~C<�?<v<<��8<vx5<N�1<҇.<�+<~�'<P:$<Q� <�p<�<�<�e<�<��<�	<gK<<���;�i�;��;���;���;ь�;6w�;Rp�;Sw�;Z��;���;��;{'�;y�;�ګ;�J�;!ˠ;�Z�;���;��;�g�;k6�;��;ix;��m;
d;�NZ;�P;G;ҫ=;a\4;%)+;_";�;�;;z;���:p��:̦�:���:@t�:|$�:��:v�:�t:jmU:]�6:�:c��9��9BRy99��~7GƸ�(U�����۹dR	���$��3@��P[�'?v�;|��������������ʺ=�ֺ��㺓l����I��[#��c�*�����6$��-*��R0��t6���<�ʪB��H�|�N�,�T���Z�) a�
g�(m�Ls�$y��+�5�������k���"�����������|���*���ZȚ��  �  �f==c�=tA=Q�=�|="=� =�S =��<��<�N�<��<]��<���<"�<sT�<���<ݵ�<���<��<?�<j�<̓�<��<���<��<}+�<PM�<om�<���<��<���<���<E��<��<w�<%'�<v4�<c?�<�G�<�M�<�P�<�Q�<;O�<+J�<6B�<77�<<)�<+�<��<[��<���<x��<��<�l�<`D�<W�<���<W��<M~�<�C�<&�<���<�|�<�2�<A��<���<S>�<��<��<	'�<=¿<�Y�<T�<;}�<f	�<ڑ�<��<嗵<��<���<~�<�y�<��<�V�<@��<�&�<N��<��<�H�<���<���<uQ�<���<u��<�C�<%��<bږ<�"�<�h�<B��<��<41�<�p�<!��< �<(�<�b�<���<�Ձ<��<��|<��x<�eu<~�q<�>n<��j<�g<�c<��_<�\\<�X<|:U< �Q<"N<�J<�G<�~C<=�?<
v<<��8<�x5<y�1<��.<�+<|�'<\:$<i� <�p<<�<�e<�<l�<��	<oK<<���;�i�;��;���;¯�;���;mw�;,p�;@w�;"��;���;�;�'�;dy�;kګ;�J�;�ʠ;�Z�;��;ި�;�g�;6�;�;�x;��m;�d;OZ;[�P;�G;:�=;?\4;{)+;?";;!<;�y;���:���:��:���:+t�:i$�:��:E�:>�t:�nU:Q�6:�:���9�߷9�Ry9�9�7�9ƸO#U����,۹�R	���$��1@�iR[��>v�|���������{��#ʺ��ֺF�㺻l���]��#��d������A$�}-*�CS0�t6�+�<���B�M�H��N�&�T�W�Z���`��
g��m�6s�|$y��+�s���>���!���ӥ��񪎻԰������A���)Ț��  �  �f==_�=xA=M�=�|=+=� =�S =��<��<�N�<��<b��<���<""�<eT�<���<��<���<��<�>�<*j�<Ɠ�<��<���<��<�+�<KM�<mm�<���<&��<{��<���<I��<n�<y�<'�<�4�<k?�<�G�<�M�<�P�<�Q�<3O�<1J�<)B�<G7�<C)�< �<��<^��<���<j��<��<�l�<bD�<X�<���<f��<R~�<�C�<�<���<�|�<�2�<D��<���<Y>�<��<��<'�<?¿<�Y�<D�<;}�<Y	�<ۑ�<��<ܗ�<��<���<{�<�y�<��<�V�<A��<�&�<B��<��<�H�<���<���<}Q�<���<c��<�C�<*��<fږ<�"�<�h�<V��<��<01�<�p�<0��<&�<�'�<�b�<���<�Ձ<��<��|<��x<fu<��q<�>n<Ϫj<�g<
�c<��_<�\\<N�X<m:U<"�Q<N<0�J<�G<�~C<,�?<v<<��8<bx5<s�1<��.<�+<}�'<C:$<t� <�p<<Ϲ<�e<<x�<��	<NK<><���;�i�;��;���;���;v��;bw�;p�;�w�;��;���;!�;n'�;ly�;(ګ; K�;ˠ;�Z�;��;稐;�g�;�5�;6�;Cx;�m;#d;�NZ;P�P;�G;��=;�[4;r)+;U";�;'<;ky;w��:��:!��:���:\t�:q%�:�:��:^�t:YoU:�6:�:���9�9�]y9�9�7�FƸ #U�M��d۹<O	�d�$�\2@�S[�Z=v�|�����񢺟��_���ʺ�ֺ���<l�������"��d�Ϟ�
��[$��,*�:S0�$t6���<���B��H�k�N���T���Z�>�`��
g��m��s��#y�T+�������������������°��=���`���$Ț��  �  �f==_�={A=J�=�|=%=� =�S =	��<��<�N�<��<Y��<���<"�<qT�<���<ӵ�<���<��<�>�< j�<͓�<��<���<��<{+�<[M�<qm�<���<��<���<���<G��<j�<v�<('�<4�<c?�<�G�<�M�<�P�<wQ�<AO�</J�<*B�<E7�<;)�<#�<��<c��<���<t��<��<�l�<kD�<X�<���<N��<S~�<�C�<�<���<�|�<�2�<B��<���<H>�<	��<���<'�<9¿<�Y�<V�<9}�<W	�<ّ�<��<藵<��<���<~�<�y�<��<�V�<K��<�&�<J��<��<�H�<���<���<sQ�<���<q��<�C�<?��<`ږ<�"�<�h�<8��<��<11�<�p�<#��<,�<�'�<�b�<���<�Ձ<��<��|<��x<�eu<��q<�>n<��j<�g<��c<��_<�\\<5�X<g:U<)�Q<@N<�J<�G<�~C<�?<v<<��8<jx5<q�1<��.<�+<z�'<P:$<b� <�p<�<�<�e<�<��<��	<QK<+<���;�i�;��;s��;���;���;sw�;p�;hw�;'��;���;�;`'�;^y�;uګ;�J�;�ʠ;�Z�; ��;��;�g�;(6�;/�;Jx;�m;�d;�NZ;g�P;�G;�=;$\4;U)+;a";�;%<;�y;��:&��:X��:���:�s�:%�:X�:R�:J�t:=mU:)�6:N:���9�޷9Wy99J7�HƸ$U�v��f۹YQ	���$��1@�IQ[��>v��|��4��������ʺ)�ֺg���l���w��#��c�������A$��-*�#S0�t6���<��B���H���N���T�y�Z���`�U
g��m��s�$y�~+�k���+�������å��᪎�Ȱ��o���l���Ț��  �  �f==d�=sA=M�=�|=="� =�S =��<��<�N�<��<H��<���<"�<�T�<���<��<���<��<
?�<j�<���<��<���<��<�+�<MM�<`m�<���<��<���<���<A��<��<l�<*'�<r4�<h?�<�G�<�M�<�P�<wQ�<?O�<!J�<?B�<A7�<9)�<-�<��<m��<���<���<��<�l�<_D�<I�<���<M��<^~�<�C�<$�<���<�|�<3�<4��<���<H>�<
��<��<'�<A¿<�Y�<Y�<.}�<g	�<ّ�<��<뗵<��<Ǐ�<r�<�y�<��<�V�<C��<�&�<`��<��<�H�<���<���<�Q�<���<���<�C�<-��<Rږ<�"�<�h�<>��<��<$1�<�p�<��<0�<(�<�b�<���<�Ձ<��<��|<��x<�eu<��q<�>n<��j<�g<�c<��_<�\\<$�X<�:U<��Q<1N<�J<�G<�~C<.�?<.v<<��8<�x5<X�1<͇.<�+<��'<d:$<?� <�p<�<
�<�e<<��<��	<{K<<��;�i�;��;���;ү�;���;-w�;[p�;6w�;/��;���;�;�'�;:y�;~ګ;�J�;ˠ;�Z�;���;��;�g�;!6�;��;�x;��m;�d;!OZ;�P;G;��=;�\4;)+;";u;�;;dz;��:،�:���:���:)t�:�$�:��:q�:ҝt:DmU:K�6::���9��9�Oy9�9ȵ~79Ƹ�#U���x۹�R	���$�3@�0S[��=v��|�������
������ʺ��ֺ���l�m������#�rd�k������$��-*��R0��t6���<�]�B���H�&�N�M�T�9�Z���`��
g�Mm�,s�F$y��+�e���V������񥋻�̰������!���qȚ��  �  �f==d�=xA=J�=�|= =!� =�S =��<��<�N�<��<^��<���<"�<rT�<���<ݵ�<���<��<?�<j�<Г�<��<���<��<�+�<VM�<om�<���<��<���<���<?��<t�<i�<''�<�4�<g?�<�G�<�M�<�P�<|Q�<FO�<-J�</B�<77�<=)�<)�<��<i��<���<n��<��<�l�<oD�<U�<���<K��<X~�<�C�<"�<���<�|�<�2�<?��<���<O>�<��<��<	'�<@¿<�Y�<W�<.}�<[	�<ӑ�<��<뗵<��<ď�<|�<�y�<��<�V�<Q��<�&�<M��<��<�H�<���<���<zQ�<���<o��<�C�<=��<gږ<�"�<�h�<=��<	��< 1�<�p�<��<#�<�'�<�b�<���<�Ձ<��<��|<��x<�eu<��q<�>n<��j<�g<ނc<��_< ]\<+�X<�:U<�Q<<N<�J<�G<�~C<!�?<v<<��8<�x5<O�1<Ƈ.<�+<g�'<Q:$<l� <�p<<�<�e<�<|�<��	<|K<	<���;�i�;��;���;��;���;iw�;Wp�;nw�;5��;���;��;�'�;,y�;sګ;K�;ˠ;�Z�;���;��;�g�;<6�;'�;rx;��m;�d;�NZ;�P;�G;�=;�[4;d)+;�";�;<;�y;Ӥ�:v��:o��:���:Jt�:*$�:��:+�:�t:nU:L�6:�:���9q�9Zy9�9�~7�DƸ�&U�X���۹Q	��$�62@��Q[��<v�T|������2��������ʺ��ֺ��sl������#��c��������$��-*��R0��t6��<��B�.�H�~�N���T��Z���`�h
g��m��s�4$y�a+�f���l���[�������ߪ�������������>Ț��  �  �f==_�={A=H�=�|=(=� =�S =��<��<�N�<��<X��<���<"�<mT�<ą�<յ�<���<��<�>�<%j�<Γ�<��<���<��<x+�<TM�<wm�<���<��<r��<���<T��<{�<��<'�<y4�<[?�<�G�<�M�<�P�<qQ�<<O�<0J�<-B�<F7�<A)�<$�<��<_��<���<v��<��<�l�<`D�<Y�<���<b��<P~�<�C�<!�<���<�|�<�2�<D��<���<B>�<��<���<'�<1¿<�Y�<F�<D}�<g	�<䑸<��<ח�<��<���<��<�y�<��<�V�<J��<�&�<K��<��<�H�<���<���<rQ�<���<n��<�C�<)��<\ږ<�"�<�h�<A��<��<41�<�p�<,��<+�<�'�<�b�<���<Ձ<��<��|<��x<�eu<s�q<�>n<ڪj<�g<�c<��_<�\\<%�X<p:U<"�Q<>N<�J<�G<�~C<�?<v<<��8<tx5<v�1<ʇ.<�+<��'<M:$<_� <�p<�<�<�e<�<��<��	<ZK<4<���;�i�;��;a��;���;���;�w�;p�;`w�;��;ñ�;L�;�'�;�y�;=ګ;�J�;�ʠ;�Z�;��;��;�g�;6�;3�;ax;�m;d;�NZ;v�P;�G;u�=;4\4;t)+;&";};-<;�y;?��:��:o��:���:.t�:8%�:|�:p�:t:wlU:��6::d��9mܷ9=Uy9�9wc7A9Ƹ�U�_���۹�Q	���$�v1@�
R[��>v�J}��L�/�������ʺ�ֺ0���l�`�����#��d������$��-*��R0�t6�z�<���B���H���N���T�l�Z���`�m
g��m�ls�U$y��+���������W�������򪎻��������Y���$Ț��  �  �f==f�=wA=K�=�|=#=� =�S =��<��<�N�<��<_��<���<"�<oT�<���<ε�<���<��<�>�<j�<̓�<��<���<��<�+�<OM�<jm�<���<"��<���<���<=��<n�<n�<#'�<�4�<t?�<�G�<�M�<�P�<{Q�<DO�<%J�<0B�<37�<@)�<!�<��<[��<���<w��<��<�l�<mD�<S�<���<O��<K~�<�C�<�<���<�|�<�2�<7��<���<N>�<��<��<'�<H¿<�Y�<R�<1}�<W	�<Б�<��<闵<��<���<x�<�y�<��<�V�<M��<�&�<I��<��<�H�<���<���<kQ�<���<n��<�C�<5��<gږ<�"�<�h�<6��<��<&1�<�p�<"��<!�<�'�<�b�<���<�Ձ<��<��|<��x<
fu<��q<�>n<��j<�g<�c<��_<]\<L�X<�:U<�Q<4N<�J<�G<�~C<'�?<v<<��8<zx5<[�1<.<�+<��'<G:$<n� <�p<�<�<�e<�<��<��	<dK<<���;�i�;��;���;��;���;Uw�;Ap�;�w�;9��;���;��;p'�;@y�;aګ;!K�;3ˠ;�Z�;���;$��;�g�;56�;�;vx;{�m;d;�NZ;%�P;�G;�=;6\4;X)+;�";�;<;�y;��:���:ͦ�:I��:`t�:$$�:��:��:��t:�mU:��6:C:���9`�90\y9�9�~7|HƸ�(U�<��۹xO	�w�$��2@��R[�=v�M|�� �p�0�����Dʺ��ֺկ�dm�-�����9#�4d�Ğ���$��-*�S0�qt6�|�<���B�B�H�h�N��T��Z���`�
g�m�.s��#y�8+�����E���p���᥋��������B���+���EȚ��  �  �f==q�=�A=b�=�|=;=>� =�S =[��<#�<3O�<c��<���<��<}"�<�T�<(��<Y��<X��<�<�?�<�j�<r��<���<s��<��<*,�<N�<2n�<~��<֨�<Z��<���<2��<x�<k�<1(�<}5�<v@�<�H�<�N�<!R�<�R�<�P�<gK�<�C�<�8�<�*�<��<G�<���<��<���<p��<qn�<�E�<��<P��<���<��<@E�<��<���<}~�<�4�<���<o��<�?�<���<���<�(�<�ÿ<N[�<�<�~�<�<z��<E�<w��<�<E��<��<M{�<E�<X�<���<(�<���<�<�I�<���<���<�R�<���<u��<�D�<��<5ۖ<X#�<�i�<���<���<�1�<sq�<���<��<j(�<c�<ᜃ<�Ձ<��<��|<��x<�eu<��q<�>n<��j<�g<��c<2�_<_\\<g�X<�9U<8�Q<LN<�J<�G<�}C<��?<�t<<-�8<�v5<��1<��.<�+<��'<28$<#� <{n<�<l�<Cc<]<��<��	<�H<<߻�;�c�;H�;���;���;��;�p�;Bi�;p�;��;d��;�ݼ;d �;�q�;
ӫ;6C�;Yà;%S�;p�;x��;�_�;�.�;c�;��w;��m;,d;�?Z;S�P;�G;��=;:N4;<+;J";�;�.;�l;H��:=s�:���:���:�\�:��:��:>��:st:�AU:j6:��:?`�9��9c�x9��9*0v7�BǸv�U��Q��T۹�p	���$�tM@��k[�8Xv�u���#Ε��������O��ʺx�ֺ��㺵t�!��<���&�h������$�x0*�WU0��v6�u�<��B��H��N���T���Z�qa��g�
m�8s�W%y�e,�����j���>���ܥ��ժ���������������ǚ��  �  �f=#=t�=�A=a�=�|===8� =�S =R��<�<0O�<[��<���<��<�"�<�T�<*��<M��<T��<�<�?�<�j�<l��<���<s��<��<9,�<N�</n�<}��<��<]��<���<)��<c�<m�<)(�<�5�<�@�<�H�<�N�< R�<�R�<�P�<kK�<�C�<�8�<�*�<��<Q�<���<��<��<o��<}n�<�E�<��<@��<���<��<GE�<��<���<�~�<�4�<���<m��<@�<���<���<�(�<�ÿ<a[�< �<�~�<�
�<p��<F�<y��<%�<F��<��<B{�<Q�<X�<���<(�<���<�<�I�<���<���<�R�<���<g��<�D�<��<Aۖ<R#�<�i�<�<���<�1�<jq�<���<��<f(�<c�<䜃<�Ձ<��<�|<��x<fu<��q<�>n<��j<`g<��c<'�_<m\\<��X<�9U<0�Q<<N<�J<�G<�}C<��?<�t<<4�8<�v5<��1<�.<�+<y�'<#8$<6� <�n<�<W�<Gc<D<��<��	<H<<Ļ�;�c�;J�;��;6��;���;xp�;<i�;lp�;���;\��;�ݼ; �;�q�;�ҫ;uC�;�à;"S�;J�;t��;<`�;�.�;t�;s�w;��m;�d;�?Z;��P;G;ɝ=;�M4;;+;�";6;�.;�l;f��:Zr�:#��:	��:3\�:	�:��:i��:�rt:�CU:Yj6:M�:N`�9W��9��x9��9�Av7�TǸ��U��Q���S۹n	���$��M@�9m[��Vv�l���Ε�����������$ʺ�ֺҸ㺘u�~!������&��g�(��@��?$��0*��U0��v6���<�*�B� �H�>�N���T���Z�� a��g�6m�Gs��$y�,�����q�������祋�쪎�����:��������ǚ��  �  �f=!=n�=�A=c�=�|=@=4� =�S =N��<'�<9O�<]��<���<��<�"�<�T�<7��<R��<S��<�<�?�<�j�<i��<���<r��<��<7,�<N�<6n�<m��<��<T��<���<4��<e�<x�<(�<�5�<t@�<�H�<�N�<R�<�R�<uP�<wK�<~C�<�8�<�*�<��<W�<���<��<��<r��<nn�<�E�<��<?��<��<��<ME�<��<���<�~�<�4�<���<a��<�?�<���<���<�(�<�ÿ<_[�<��<�~�< �<z��<J�<o��<#�<8��<��<D{�<L�<X�<���<$(�<���<%�<�I�<���<���<�R�<���<g��<�D�<��<9ۖ<V#�<�i�<���<���<�1�<dq�<���<��<i(�<$c�<ל�<�Ձ<��<��|<��x<	fu<��q<�>n<��j<dg<��c<"�_<`\\<��X<�9U<B�Q<9N<�J<�G<�}C<��?<�t<<A�8<�v5<��1<�.<�+<��'<(8$<)� <pn<�<Y�<`c<M<��<Ȇ	<qH<1<���;�c�;E�;���;/��;Ņ�;�p�;�h�;^p�;Յ�;f��;�ݼ; �;r�;�ҫ;lC�;Pà;S�;e�;`��;`�;h.�;��;b�w;�m;d;@Z;ٖP;G;,�=;�M4;O+;/";�;�.;ul;>��:Er�:|��:2��:F\�:��:��:#��:Zqt:�BU:zi6:��:�`�9���9��x9�~9��v7�OǸ̤U�nP��V۹On	���$��L@��l[�RWv�/����Ε��������7��mʺ��ֺ���{u� ������&�0h�g��"��$�70*��U0�zv6��<�
�B���H�"�N���T�1�Z�a��g��m��s�%y�7,�̙��F�������������������T���,����ǚ��  �  �f= =r�=�A=b�=�|=<=;� =�S =Q��<%�<+O�<a��<���<��<�"�<�T�<#��<V��<R��<�<�?�<�j�<h��<���<u��<��<5,�<N�<-n�<x��<��<b��<���<+��<h�<j�<+(�<�5�<{@�<�H�<�N�< R�<�R�<}P�<qK�<{C�<�8�<�*�<��<J�<���<��<��<q��<yn�<�E�<��<B��<��<��<AE�<��<���<�~�<�4�<���<j��<@�<���<���<�(�<�ÿ<a[�<�<�~�< �<s��<D�<}��<"�<B��<��<H{�<L�<	X�<���<(�<���<�<�I�<���<���<�R�<���<m��<�D�<��<=ۖ<W#�<�i�<���<���<�1�<nq�<���<��<e(�< c�<���<�Ձ<��<�|<��x<fu<��q<�>n<��j<sg<��c<.�_<u\\<��X<�9U<5�Q<AN<�J<�G<�}C<��?<�t<<1�8<�v5<��1<�.<�+<n�'</8$</� <�n<�<d�<8c<V<��<��	<�H<<���;�c�;P�;���;$��;ԅ�;mp�;*i�;\p�;��;`��;�ݼ;! �;�q�;�ҫ;�C�;mà;S�;a�;v��;`�;�.�;��;G�w;��m;d;)@Z;o�P;MG;��=;�M4;I+;�";;�.;�l;��:�r�:Ǎ�:@��:y\�:�:��:���:vrt:CU:j6:�:�_�9��9��x9}�9�0v7�PǸB�U��Q���R۹cn	�]�$�5N@��l[�ZWv����Ε�g���������ʺ�ֺ���u��!��z���&��g�E����d$�p0*��U0��v6���<�*�B�$�H�?�N���T���Z�'a��g�m�Zs��$y��+���������q�������ު������P���	����ǚ��  �  �f==s�=�A=b�=�|=:=>� =�S =W��<%�<1O�<e��<���<��<s"�<�T�<'��<Z��<S��<�<�?�<�j�<s��<���<s��<��<2,�<N�<*n�<���<ݨ�<_��<���<1��<w�<h�<,(�<5�<�@�<�H�<�N�<%R�<�R�<P�<iK�<�C�<�8�<�*�<��<D�<���<��<��<i��<xn�<�E�<��<P��<��<��<=E�<��<���<�~�<�4�<���<k��<�?�<���<���<�(�<�ÿ<Q[�<�<�~�<�<{��<B�<|��<�<K��<��<L{�<L�<X�<���<(�<���<�<�I�<���<���<�R�<���<y��<�D�<"��<6ۖ<W#�<�i�<���<���<�1�<uq�<���<��<h(�<c�<圃<�Ձ<��<�|<��x<fu<��q<�>n<~�j<�g<��c<.�_<b\\<{�X<�9U<.�Q<KN<��J<�G<�}C<��?<�t<<)�8<�v5<��1<��.<�+<|�'<78$<� <�n<~<z�<@c<_<��<��	<�H<<��;�c�;I�;���;��;��;ap�;Vi�;.p�;��;[��;�ݼ;_ �;�q�;�ҫ;=C�;�à; S�;`�;���;`�;�.�;l�;��w;��m;d;X@Z;B�P;�G;��=;JN4;	+;|";;E.;�l;#��:Ns�:���:���:�\�:��:N�:9��:�rt:�BU:�j6:S�:�_�9Ε�9��x9%�9}v7�BǸ$�U�cR���R۹<p	�@�$��N@�l[�hWv�툈�!Ε�����	��[���ʺ��ֺ
�㺻t�!����I'��g������$�k0*�rU0�	w6�^�<�>�B���H�*�N���T���Z�;a��g�3m�(s��$y�`,���������3�������ݪ������c����Ț��  �  �f==r�=�A=`�=�|=?=9� =�S =P��< �<0O�<d��<���<��<{"�<�T�<)��<O��<Q��<�<�?�<�j�<b��<���<y��<��<0,�<N�<4n�<w��<��<[��<���<2��<i�<p�<((�<�5�<~@�<�H�<�N�<R�<�R�<P�<xK�<wC�<�8�<�*�<��<O�<���<��<���<s��<yn�<�E�<��<D��<��<��<DE�<��<���<�~�<�4�<���<m��<�?�<���<���<�(�<�ÿ<\[�<��<�~�<�<w��<E�<x��<�<@��<��<N{�<J�<X�<���<!(�<���<�<�I�<���<���<�R�<���<p��<�D�<��<:ۖ<[#�<�i�<�<���<�1�<kq�<���<��<_(�<&c�<✃<�Ձ<��<��|<��x<fu<��q<�>n<��j<jg<��c<+�_<b\\<��X<�9U<G�Q<BN<��J<�G<�}C<��?<�t<<=�8<�v5<��1<�.<�+<x�'<58$<#� <�n<�<l�<Dc<I<��<Ɔ	<}H<'<���;�c�;b�;���;��;��;�p�;'i�;Np�;��;^��;�ݼ;% �;�q�;�ҫ;eC�;wà;S�;��;n��;`�;�.�;��;+�w;��m; d;(@Z;��P;,G;��=;�M4;W+;�";;�.;�l;6��:tr�:���:d��:@\�:,�:O�:��:�rt:�BU:j6:	�:�_�9(��9l�x9�9�Sv7�NǸl�U��Q���S۹�n	���$��M@��k[��Wv�∈��͕�$���/�����$ʺ��ֺ��}u�!��d���&��g�`�����I$��0*��U0��v6���<��B�8�H�q�N�w�T���Z�1a��g��m�cs��$y�P,�����c�������ե��㪎�����N�������ǚ��  �  �f=&=o�=�A=b�=�|=C=3� =�S =G��<+�<-O�<^��<���<��<�"�<�T�<,��<V��<L��<�<�?�<�j�<]��<���<k��<��<8,�<
N�<4n�<r��<��<V��<���<3��<d�<v�<(�<�5�<z@�<�H�<�N�<R�<�R�<pP�<{K�<wC�<�8�<�*�<��<Q�<���<��<��<u��<un�<�E�<��<:��<��<��<EE�<��<���<�~�<�4�<���<^��<	@�<���<���<�(�<�ÿ<d[�<��<�~�<�
�<w��<H�<p��<(�<:��<��<C{�<L�<X�<���<((�<���<(�<�I�<���<���<�R�<���<f��<�D�<��<>ۖ<V#�<�i�<���<���<�1�<aq�<���<��<b(�<$c�<؜�<�Ձ<��<��|<��x<fu<��q<�>n<��j<_g<��c<�_<f\\<��X<�9U<G�Q<-N<�J<�G<�}C<��?<�t<<N�8<�v5<��1<օ.<�+<s�'<)8$<2� <zn<�<X�<Kc<U<��<ʆ	<kH<9<���;�c�;+�;���;0��;���;�p�;i�;lp�;݅�;`��;�ݼ; �;�q�;�ҫ;�C�;eà;S�;m�;X��;F`�;U.�;��;*�w;��m;d;�?Z;��P;�
G;�=;�M4;j+;k";�;�.;Ql;��:?r�:���:���:-\�:��:2�:t��:�pt:DU:�i6:
�:D_�9i��9��x9�~9�~v7�QǸ.�U�Q���U۹�m	�P�$��M@�m[�OWv�ǈ���Ε�����������ʺ��ֺ0��Gu� !������&�	h�@�� ��s$�*0*��U0��v6���<�ݬB�6�H�]�N���T�.�Z�� a�	g��m��s��$y�*,�֙��P�������ɥ����������;���$����ǚ��  �  �f=!=p�=�A=f�=�|===9� =�S =K��<&�<-O�<c��<���<��<�"�<�T�<&��<V��<Q��<�<�?�<�j�<i��<���<j��<��<2,�<N�<3n�<|��<ߨ�<\��<���<1��<m�<l�<((�<�5�<w@�<�H�<�N�<R�<�R�<tP�<tK�<�C�<�8�<�*�<��<Q�<���<��<���<q��<vn�<�E�<��<E��<���<��<FE�<��<���<�~�<�4�<���<a��<@�<���<���<�(�<�ÿ<X[�<��<�~�<�<y��<G�<y��<�<B��<��<K{�<H�<
X�<���<&(�<���<�<�I�<���<���<�R�<���<o��<�D�<��<<ۖ<W#�<�i�<���<���<�1�<mq�<���<��<o(�<c�<ܜ�<�Ձ<��<��|<��x<fu<��q<�>n<��j<}g<��c<,�_<h\\<{�X<�9U<B�Q<@N<�J<�G<�}C<��?<�t<<4�8<�v5<��1<ޅ.<�+<s�'<48$<.� <�n<�<i�<?c<W<��<φ	<}H<<���;�c�;'�;���;��;߅�;�p�;8i�;6p�;���;l��;�ݼ;7 �;�q�;�ҫ;\C�;]à;S�;v�;l��;!`�;f.�;��;��w;��m;d;:@Z;��P;*G;ٝ=;�M4;H+;o";�;�.;�l;���:�r�:��:���:b\�:�:�:��:Rqt:CU:�i6:��:q_�9Ғ�9`�x9��9M=v7$KǸ'�U�4Q���S۹�o	�\�$��M@� l[��Wv������Ε�����������!ʺy�ֺ��u�!��j���&��g�Q����P$�Z0*��U0��v6���<�-�B�(�H���N���T��Z�a��g��m�Vs�%y�5,�����x���\���륋�⪎�����c�������ǚ��  �  �f==w�=�A=a�=�|===;� =�S =V��< �</O�<d��<���<%��<v"�<�T�<"��<T��<V��<�<�?�<�j�<k��<���<u��<��</,�<N�<$n�<���<��<c��<���<-��<q�<b�<2(�<�5�<�@�<�H�<�N�<'R�<�R�<�P�<iK�<�C�<�8�<�*�<��<J�<���<��<���<n��<}n�<F�<��<I��<��<��<CE�<��<���<�~�<�4�<���<q��<�?�<���<���<�(�<�ÿ<W[�<�<�~�<�<v��<>�<���<�<M��<��<R{�<H�<X�<���<(�<���<�<�I�<���<���<�R�<���<s��<�D�<(��<9ۖ<W#�<�i�<�<���<�1�<oq�<���<��<f(�<c�<휃<�Ձ<��<�|<��x<fu<��q<�>n<y�j<�g<��c<2�_<i\\<��X<�9U<'�Q<VN<�J<�G<�}C<��?<�t<<4�8<�v5<��1<�.<�+<w�'<58$< � <�n<�<r�<8c<S<��<��	<�H<<Ļ�;�c�;P�;��;��;��;Mp�;Zi�;Bp�;��;R��;�ݼ;G �;�q�;ӫ;ZC�;�à;S�;n�;���;�_�;�.�;m�;��w;��m;*d;&@Z;q�P;yG;u�=;N4;1+;�";Q;v.;�l;Ɗ�:/s�:��:M��:�\�:�:��:9��:^st:dBU:�j6:��:#^�9k��9ݿx9n�9a�u7�IǸy�U�qS��MQ۹�o	��$�KO@�Bk[��Wv�ʈ���͕�����������ʺ�ֺǸ�u�"��L��$'�^g�k����3$��0*�|U0��v6���<�'�B�+�H�:�N���T���Z�xa�dg�>m�<s��$y�B,���������D�������ժ������J���ﾗ�Ț��  �  �f==s�=�A=c�=�|=?=8� =�S =N��<&�<6O�<d��<���<��<w"�<�T�<2��<T��<Q��<�<�?�<�j�<f��<���<p��<��<0,�<N�<)n�<|��<��<X��<���<4��<m�<q�<&(�<�5�<~@�<�H�<�N�<$R�<�R�<{P�<pK�<�C�<�8�<�*�<��<M�<���<��<���<p��<sn�<�E�<��<H��<���<��<DE�<��<���<�~�<�4�<���<f��<�?�<���<���<�(�<�ÿ<V[�<��<�~�<�<z��<D�<u��<�<E��<��<L{�<I�<	X�<���<(�<���<�<�I�<���<���<�R�<���<r��<�D�<��<4ۖ<X#�<�i�<���<���<�1�<iq�<���<��<i(�<c�<㜃<�Ձ<��<�|<��x<fu<��q<�>n<��j<wg<��c<'�_<\\\<��X<�9U<+�Q<KN<��J<�G<�}C<��?<�t<<;�8<�v5<��1<�.<�+<��'<58$<� <�n<�<r�<Vc<R<��<��	<�H<!<���;�c�;@�;���;��;��;ap�;<i�;Ap�;��;]��;�ݼ;7 �;�q�;�ҫ;OC�;wà;S�;b�;���;`�;�.�;��;��w;��m;d;@Z;��P;6G;�=;N4;B+;W";�;�.;�l;ċ�:�r�:���:#��:`\�:$�:��:���:�qt:�BU:lj6:Q�:�^�9p��94�x9�9FYv70KǸϤU��Q���T۹�o	���$��N@�l[��Wv�����Ε�K����������ʺ
�ֺ��@u�!��O��'��g������$�G0*��U0��v6���<��B�C�H�%�N���T���Z�Ua��g�/m�Qs��$y�h,�����a���i���ѥ��몎�����O������Ț��  �  �f=#=t�=�A=d�=�|=@=6� =�S =E��<'�<*O�<_��<���<��<�"�<�T�<*��<O��<K��<�<�?�<�j�<^��<���<u��<��<4,�<N�<7n�<u��<��<_��<���<.��<_�<s�< (�<�5�<v@�<�H�<�N�<R�<�R�<|P�<wK�<zC�<�8�<�*�<��<U�<���<��<��<x��<yn�<�E�<��<;��<���<��<IE�<��<���<�~�<�4�<���<g��<@�<���<���<�(�<�ÿ<i[�<��<�~�<�
�<q��<E�<w��<(�<=��< �<F{�<K�<X�<���<%(�<���<�<�I�<���<���<�R�<���<f��<�D�<��<?ۖ<X#�<�i�<���<���<�1�<eq�<���<��<h(�<"c�<㜃<�Ձ<��<��|<��x<fu<��q<�>n<��j<Vg<��c<�_<|\\<��X<�9U<E�Q<1N<�J<�G<�}C<��?<�t<<?�8<�v5<��1<҅.<�+<m�'<,8$<8� <~n<�<\�<Fc<I<��<ǆ	<|H<%<���;�c�;P�;��; ��;�;�p�; i�;hp�;��;\��;�ݼ;��;�q�;�ҫ;�C�;Yà;)S�;n�;]��;D`�;�.�;��;D�w;��m;d;�?Z;ʖP;�
G;��=;�M4;�+;�";;�.;Wl;���:r�:H��:���:#\�:��:_�:%��:rt:nDU:�i6:i�:la�9Z��9��x9��9u^v7�XǸa�U��Q��T۹�m	��$��L@��l[��Wv�X���MΕ�����>�����Hʺ��ֺ�㺠u�n!������&��g�7�����$�?0*�(V0��v6�ߓ<��B�d�H�.�N���T���Z�� a��g��m�Os�%y��+�֙��c�������ۥ�� ������M�������ǚ��  �  �f==t�=�A=a�=�|=A=7� =�S =Q��<,�<2O�<a��<���<��<|"�<�T�<-��<Y��<S��<�<�?�<�j�<k��<���<r��<��<0,�<N�<1n�<z��<��<]��<���<7��<o�<r�<!(�<�5�<v@�<�H�<�N�<R�<�R�<P�<mK�<�C�<�8�<�*�<��<P�<���<��<���<r��<on�<�E�<��<G��<���<��<GE�<��<���<�~�<�4�<���<k��<�?�<���<���<�(�<�ÿ<[[�<��<�~�<�<}��<B�<v��<�<@��<��<G{�<H�<
X�<���<(�<���<$�<�I�<���<���<�R�<���<q��<�D�<��<4ۖ<W#�<�i�<���<���<�1�<eq�<���<��<f(�<c�<圃<�Ձ<��<�|<��x<fu<��q<�>n<��j<zg<��c<�_<i\\<v�X<�9U<9�Q<@N<��J<�G<�}C<��?<�t<<D�8<�v5<��1<�.<�+<|�'<.8$<"� <{n<�<j�<Lc<]<��<��	<�H<-<»�;�c�;G�;��;��;؅�;p�;2i�;Ap�;���;O��;�ݼ;A �;�q�;�ҫ;cC�;Wà; S�;c�;h��;`�;�.�;}�;��w; �m;Bd;�?Z;��P;YG;�=;�M4;Q+;:";�;�.;�l;Ћ�: s�:!��:���:�\�:��:�:z��:�rt:�BU:�i6:�:A`�9���9��x9��9jMv7�GǸ	�U�iR��YT۹�n	���$��M@��l[��Wv�����@Ε�����s��O��ʺ`�ֺԸ��t�F!��_���&�h������<$�0*��U0��v6��<��B��H�9�N���T���Z�=a��g�m�Fs�.%y�+,�ڙ��P���c���ť���������m��������ǚ��  �  �f==u�=�A=`�=�|=:=;� =�S =T��<�<+O�<e��<���<#��<}"�<�T�<!��<I��<U��<�<�?�<�j�<h��<���<w��<��<3,�<N�<(n�<���<��<f��<���<+��<`�<l�<0(�<�5�<�@�<�H�<�N�<&R�<�R�<�P�<lK�<�C�<�8�<�*�<��<Q�<���<��<���<p��<|n�<F�<��<J��<��<��<GE�<��<���<{~�<�4�<���<w��<�?�<���<���<�(�<�ÿ<Y[�<	�<�~�<�
�<r��<D�<���<�<M��<��<G{�<L�<	X�<���<(�<���<�<�I�<���<���<�R�<���<y��<�D�<)��<;ۖ<Z#�<�i�<譑<���<�1�<mq�<���<��<e(�<c�<꜃<�Ձ<��<ڊ|<��x<fu<��q<�>n<��j<bg<��c<+�_<l\\<��X<�9U<'�Q<XN<�J<�G<�}C<��?<�t<<(�8<�v5<��1<��.<�+<p�'<88$<+� <�n<�<{�<5c<=<��<��	<�H<<���;vc�;Z�;��;��;��;Zp�;fi�;Cp�;��;a��;�ݼ; �;�q�;ӫ;WC�;�à;!S�;H�;���;�_�;�.�;w�;��w;x�m;�d;7@Z;��P;=G;Y�=;�M4;D+;�";N;�.;�l;���:�r�:!��:k��:H\�:��:#�:P��:tt:BU:�j6:m�:_�9��9��x9ԉ9�0v7�TǸ�U�R��}Q۹ o	��$��N@��l[�OWv�����͕��������_���ʺ��ֺ��㺡u�9"�����&�Sg�U����`$��0*��U0��v6���<�a�B�]�H�C�N���T���Z�ta�Yg�`m�s��$y�<,�����n�������䥋�㪎�����P���ܾ��Ț��  �  �f==t�=�A=a�=�|=A=7� =�S =Q��<,�<2O�<a��<���<��<|"�<�T�<-��<Y��<S��<�<�?�<�j�<k��<���<r��<��<0,�<N�<1n�<z��<��<]��<���<7��<o�<r�<!(�<�5�<v@�<�H�<�N�<R�<�R�<P�<mK�<�C�<�8�<�*�<��<P�<���<��<���<r��<on�<�E�<��<G��<���<��<GE�<��<���<�~�<�4�<���<k��<�?�<���<���<�(�<�ÿ<[[�<��<�~�<�<}��<B�<v��<�<@��<��<G{�<H�<
X�<���<(�<���<$�<�I�<���<���<�R�<���<q��<�D�<��<4ۖ<W#�<�i�<���<���<�1�<eq�<���<��<f(�<c�<圃<�Ձ<��<�|<��x<fu<��q<�>n<��j<zg<��c<�_<i\\<v�X<�9U<9�Q<@N<��J<�G<�}C<��?<�t<<D�8<�v5<��1<�.<�+<|�'<.8$<"� <{n<�<j�<Lc<]<��<��	<�H<-<»�;�c�;G�;��;��;؅�;p�;2i�;Ap�;���;O��;�ݼ;A �;�q�;�ҫ;cC�;Wà; S�;c�;h��;`�;�.�;}�;��w; �m;Bd;�?Z;��P;YG;�=;�M4;Q+;:";�;�.;�l;Ћ�: s�:!��:���:�\�:��:�:z��:�rt:�BU:�i6:�:A`�9���9��x9��9jMv7�GǸ	�U�iR��YT۹�n	���$��M@��l[��Wv�����@Ε�����s��O��ʺ`�ֺԸ��t�F!��_���&�h������<$�0*��U0��v6��<��B��H�9�N���T���Z�=a��g�m�Fs�.%y�+,�ڙ��P���c���ť���������m��������ǚ��  �  �f=#=t�=�A=d�=�|=@=6� =�S =E��<'�<*O�<_��<���<��<�"�<�T�<*��<O��<K��<�<�?�<�j�<^��<���<u��<��<4,�<N�<7n�<u��<��<_��<���<.��<_�<s�< (�<�5�<v@�<�H�<�N�<R�<�R�<|P�<wK�<zC�<�8�<�*�<��<U�<���<��<��<x��<yn�<�E�<��<;��<���<��<IE�<��<���<�~�<�4�<���<g��<@�<���<���<�(�<�ÿ<i[�<��<�~�<�
�<q��<E�<w��<(�<=��< �<F{�<K�<X�<���<%(�<���<�<�I�<���<���<�R�<���<f��<�D�<��<?ۖ<X#�<�i�<���<���<�1�<eq�<���<��<h(�<"c�<㜃<�Ձ<��<��|<��x<fu<��q<�>n<��j<Vg<��c<�_<|\\<��X<�9U<E�Q<1N<�J<�G<�}C<��?<�t<<?�8<�v5<��1<҅.<�+<m�'<,8$<8� <~n<�<\�<Fc<I<��<ǆ	<|H<%<���;�c�;P�;��; ��;�;�p�; i�;hp�;��;\��;�ݼ;��;�q�;�ҫ;�C�;Yà;)S�;n�;]��;D`�;�.�;��;D�w;��m;d;�?Z;ʖP;�
G;��=;�M4;�+;�";;�.;Wl;���:r�:H��:���:#\�:��:_�:%��:rt:nDU:�i6:i�:la�9Z��9��x9��9u^v7�XǸa�U��Q��T۹�m	��$��L@��l[��Wv�X���MΕ�����>�����Hʺ��ֺ�㺠u�n!������&��g�7�����$�?0*�(V0��v6�ߓ<��B�d�H�.�N���T���Z�� a��g��m�Os�%y��+�֙��c�������ۥ�� ������M�������ǚ��  �  �f==s�=�A=c�=�|=?=8� =�S =N��<&�<6O�<d��<���<��<w"�<�T�<2��<T��<Q��<�<�?�<�j�<f��<���<p��<��<0,�<N�<)n�<|��<��<X��<���<4��<m�<q�<&(�<�5�<~@�<�H�<�N�<$R�<�R�<{P�<pK�<�C�<�8�<�*�<��<M�<���<��<���<p��<sn�<�E�<��<H��<���<��<DE�<��<���<�~�<�4�<���<f��<�?�<���<���<�(�<�ÿ<V[�<��<�~�<�<z��<D�<u��<�<E��<��<L{�<I�<	X�<���<(�<���<�<�I�<���<���<�R�<���<r��<�D�<��<4ۖ<X#�<�i�<���<���<�1�<iq�<���<��<i(�<c�<㜃<�Ձ<��<�|<��x<fu<��q<�>n<��j<wg<��c<'�_<\\\<��X<�9U<+�Q<KN<��J<�G<�}C<��?<�t<<;�8<�v5<��1<�.<�+<��'<58$<� <�n<�<r�<Vc<R<��<��	<�H<!<���;�c�;@�;���;��;��;ap�;<i�;Ap�;��;]��;�ݼ;7 �;�q�;�ҫ;OC�;wà;S�;b�;���;`�;�.�;��;��w;��m;d;@Z;��P;6G;�=;N4;B+;W";�;�.;�l;ċ�:�r�:���:#��:`\�:$�:��:���:�qt:�BU:lj6:Q�:�^�9p��94�x9�9FYv70KǸϤU��Q���T۹�o	���$��N@�l[��Wv�����Ε�K����������ʺ
�ֺ��@u�!��O��'��g������$�G0*��U0��v6���<��B�C�H�%�N���T���Z�Ua��g�/m�Qs��$y�h,�����a���i���ѥ��몎�����O������Ț��  �  �f==w�=�A=a�=�|===;� =�S =V��< �</O�<d��<���<%��<v"�<�T�<"��<T��<V��<�<�?�<�j�<k��<���<u��<��</,�<N�<$n�<���<��<c��<���<-��<q�<b�<2(�<�5�<�@�<�H�<�N�<'R�<�R�<�P�<iK�<�C�<�8�<�*�<��<J�<���<��<���<n��<}n�<F�<��<I��<��<��<CE�<��<���<�~�<�4�<���<q��<�?�<���<���<�(�<�ÿ<W[�<�<�~�<�<v��<>�<���<�<M��<��<R{�<H�<X�<���<(�<���<�<�I�<���<���<�R�<���<s��<�D�<(��<9ۖ<W#�<�i�<�<���<�1�<oq�<���<��<f(�<c�<휃<�Ձ<��<�|<��x<fu<��q<�>n<y�j<�g<��c<2�_<i\\<��X<�9U<'�Q<VN<�J<�G<�}C<��?<�t<<4�8<�v5<��1<�.<�+<w�'<58$< � <�n<�<r�<8c<S<��<��	<�H<<Ļ�;�c�;P�;��;��;��;Mp�;Zi�;Bp�;��;R��;�ݼ;G �;�q�;ӫ;ZC�;�à;S�;n�;���;�_�;�.�;m�;��w;��m;*d;&@Z;q�P;yG;u�=;N4;1+;�";Q;v.;�l;Ɗ�:/s�:��:M��:�\�:�:��:9��:^st:dBU:�j6:��:#^�9k��9ݿx9n�9a�u7�IǸy�U�qS��MQ۹�o	��$�KO@�Bk[��Wv�ʈ���͕�����������ʺ�ֺǸ�u�"��L��$'�^g�k����3$��0*�|U0��v6���<�'�B�+�H�:�N���T���Z�xa�dg�>m�<s��$y�B,���������D�������ժ������J���ﾗ�Ț��  �  �f=!=p�=�A=f�=�|===9� =�S =K��<&�<-O�<c��<���<��<�"�<�T�<&��<V��<Q��<�<�?�<�j�<i��<���<j��<��<2,�<N�<3n�<|��<ߨ�<\��<���<1��<m�<l�<((�<�5�<w@�<�H�<�N�<R�<�R�<tP�<tK�<�C�<�8�<�*�<��<Q�<���<��<���<q��<vn�<�E�<��<E��<���<��<FE�<��<���<�~�<�4�<���<a��<@�<���<���<�(�<�ÿ<X[�<��<�~�<�<y��<G�<y��<�<B��<��<K{�<H�<
X�<���<&(�<���<�<�I�<���<���<�R�<���<o��<�D�<��<<ۖ<W#�<�i�<���<���<�1�<mq�<���<��<o(�<c�<ܜ�<�Ձ<��<��|<��x<fu<��q<�>n<��j<}g<��c<,�_<h\\<{�X<�9U<B�Q<@N<�J<�G<�}C<��?<�t<<4�8<�v5<��1<ޅ.<�+<s�'<48$<.� <�n<�<i�<?c<W<��<φ	<}H<<���;�c�;'�;���;��;߅�;�p�;8i�;6p�;���;l��;�ݼ;7 �;�q�;�ҫ;\C�;]à;S�;v�;l��;!`�;f.�;��;��w;��m;d;:@Z;��P;*G;ٝ=;�M4;H+;o";�;�.;�l;���:�r�:��:���:b\�:�:�:��:Rqt:CU:�i6:��:q_�9Ғ�9`�x9��9M=v7$KǸ'�U�4Q���S۹�o	�\�$��M@� l[��Wv������Ε�����������!ʺy�ֺ��u�!��j���&��g�Q����P$�Z0*��U0��v6���<�-�B�(�H���N���T��Z�a��g��m�Vs�%y�5,�����x���\���륋�⪎�����c�������ǚ��  �  �f=&=o�=�A=b�=�|=C=3� =�S =G��<+�<-O�<^��<���<��<�"�<�T�<,��<V��<L��<�<�?�<�j�<]��<���<k��<��<8,�<
N�<4n�<r��<��<V��<���<3��<d�<v�<(�<�5�<z@�<�H�<�N�<R�<�R�<pP�<{K�<wC�<�8�<�*�<��<Q�<���<��<��<u��<un�<�E�<��<:��<��<��<EE�<��<���<�~�<�4�<���<^��<	@�<���<���<�(�<�ÿ<d[�<��<�~�<�
�<w��<H�<p��<(�<:��<��<C{�<L�<X�<���<((�<���<(�<�I�<���<���<�R�<���<f��<�D�<��<>ۖ<V#�<�i�<���<���<�1�<aq�<���<��<b(�<$c�<؜�<�Ձ<��<��|<��x<fu<��q<�>n<��j<_g<��c<�_<f\\<��X<�9U<G�Q<-N<�J<�G<�}C<��?<�t<<N�8<�v5<��1<օ.<�+<s�'<)8$<2� <zn<�<X�<Kc<U<��<ʆ	<kH<9<���;�c�;+�;���;0��;���;�p�;i�;lp�;݅�;`��;�ݼ; �;�q�;�ҫ;�C�;eà;S�;m�;X��;F`�;U.�;��;*�w;��m;d;�?Z;��P;�
G;�=;�M4;j+;k";�;�.;Ql;��:?r�:���:���:-\�:��:2�:t��:�pt:DU:�i6:
�:D_�9i��9��x9�~9�~v7�QǸ.�U�Q���U۹�m	�P�$��M@�m[�OWv�ǈ���Ε�����������ʺ��ֺ0��Gu� !������&�	h�@�� ��s$�*0*��U0��v6���<�ݬB�6�H�]�N���T�.�Z�� a�	g��m��s��$y�*,�֙��P�������ɥ����������;���$����ǚ��  �  �f==r�=�A=`�=�|=?=9� =�S =P��< �<0O�<d��<���<��<{"�<�T�<)��<O��<Q��<�<�?�<�j�<b��<���<y��<��<0,�<N�<4n�<w��<��<[��<���<2��<i�<p�<((�<�5�<~@�<�H�<�N�<R�<�R�<P�<xK�<wC�<�8�<�*�<��<O�<���<��<���<s��<yn�<�E�<��<D��<��<��<DE�<��<���<�~�<�4�<���<m��<�?�<���<���<�(�<�ÿ<\[�<��<�~�<�<w��<E�<x��<�<@��<��<N{�<J�<X�<���<!(�<���<�<�I�<���<���<�R�<���<p��<�D�<��<:ۖ<[#�<�i�<�<���<�1�<kq�<���<��<_(�<&c�<✃<�Ձ<��<��|<��x<fu<��q<�>n<��j<jg<��c<+�_<b\\<��X<�9U<G�Q<BN<��J<�G<�}C<��?<�t<<=�8<�v5<��1<�.<�+<x�'<58$<#� <�n<�<l�<Dc<I<��<Ɔ	<}H<'<���;�c�;b�;���;��;��;�p�;'i�;Np�;��;^��;�ݼ;% �;�q�;�ҫ;eC�;wà;S�;��;n��;`�;�.�;��;+�w;��m; d;(@Z;��P;,G;��=;�M4;W+;�";;�.;�l;6��:tr�:���:d��:@\�:,�:O�:��:�rt:�BU:j6:	�:�_�9(��9l�x9�9�Sv7�NǸl�U��Q���S۹�n	���$��M@��k[��Wv�∈��͕�$���/�����$ʺ��ֺ��}u�!��d���&��g�`�����I$��0*��U0��v6���<��B�8�H�q�N�w�T���Z�1a��g��m�cs��$y�P,�����c�������ե��㪎�����N�������ǚ��  �  �f==s�=�A=b�=�|=:=>� =�S =W��<%�<1O�<e��<���<��<s"�<�T�<'��<Z��<S��<�<�?�<�j�<s��<���<s��<��<2,�<N�<*n�<���<ݨ�<_��<���<1��<w�<h�<,(�<5�<�@�<�H�<�N�<%R�<�R�<P�<iK�<�C�<�8�<�*�<��<D�<���<��<��<i��<xn�<�E�<��<P��<��<��<=E�<��<���<�~�<�4�<���<k��<�?�<���<���<�(�<�ÿ<Q[�<�<�~�<�<{��<B�<|��<�<K��<��<L{�<L�<X�<���<(�<���<�<�I�<���<���<�R�<���<y��<�D�<"��<6ۖ<W#�<�i�<���<���<�1�<uq�<���<��<h(�<c�<圃<�Ձ<��<�|<��x<fu<��q<�>n<~�j<�g<��c<.�_<b\\<{�X<�9U<.�Q<KN<��J<�G<�}C<��?<�t<<)�8<�v5<��1<��.<�+<|�'<78$<� <�n<~<z�<@c<_<��<��	<�H<<��;�c�;I�;���;��;��;ap�;Vi�;.p�;��;[��;�ݼ;_ �;�q�;�ҫ;=C�;�à; S�;`�;���;`�;�.�;l�;��w;��m;d;X@Z;B�P;�G;��=;JN4;	+;|";;E.;�l;#��:Ns�:���:���:�\�:��:N�:9��:�rt:�BU:�j6:S�:�_�9Ε�9��x9%�9}v7�BǸ$�U�cR���R۹<p	�@�$��N@�l[�hWv�툈�!Ε�����	��[���ʺ��ֺ
�㺻t�!����I'��g������$�k0*�rU0�	w6�^�<�>�B���H�*�N���T���Z�;a��g�3m�(s��$y�`,���������3�������ݪ������c����Ț��  �  �f= =r�=�A=b�=�|=<=;� =�S =Q��<%�<+O�<a��<���<��<�"�<�T�<#��<V��<R��<�<�?�<�j�<h��<���<u��<��<5,�<N�<-n�<x��<��<b��<���<+��<h�<j�<+(�<�5�<{@�<�H�<�N�< R�<�R�<}P�<qK�<{C�<�8�<�*�<��<J�<���<��<��<q��<yn�<�E�<��<B��<��<��<AE�<��<���<�~�<�4�<���<j��<@�<���<���<�(�<�ÿ<a[�<�<�~�< �<s��<D�<}��<"�<B��<��<H{�<L�<	X�<���<(�<���<�<�I�<���<���<�R�<���<m��<�D�<��<=ۖ<W#�<�i�<���<���<�1�<nq�<���<��<e(�< c�<���<�Ձ<��<�|<��x<fu<��q<�>n<��j<sg<��c<.�_<u\\<��X<�9U<5�Q<AN<�J<�G<�}C<��?<�t<<1�8<�v5<��1<�.<�+<n�'</8$</� <�n<�<d�<8c<V<��<��	<�H<<���;�c�;P�;���;$��;ԅ�;mp�;*i�;\p�;��;`��;�ݼ;! �;�q�;�ҫ;�C�;mà;S�;a�;v��;`�;�.�;��;G�w;��m;d;)@Z;o�P;MG;��=;�M4;I+;�";;�.;�l;��:�r�:Ǎ�:@��:y\�:�:��:���:vrt:CU:j6:�:�_�9��9��x9}�9�0v7�PǸB�U��Q���R۹cn	�]�$�5N@��l[�ZWv����Ε�g���������ʺ�ֺ���u��!��z���&��g�E����d$�p0*��U0��v6���<�*�B�$�H�?�N���T���Z�'a��g�m�Zs��$y��+���������q�������ު������P���	����ǚ��  �  �f=!=n�=�A=c�=�|=@=4� =�S =N��<'�<9O�<]��<���<��<�"�<�T�<7��<R��<S��<�<�?�<�j�<i��<���<r��<��<7,�<N�<6n�<m��<��<T��<���<4��<e�<x�<(�<�5�<t@�<�H�<�N�<R�<�R�<uP�<wK�<~C�<�8�<�*�<��<W�<���<��<��<r��<nn�<�E�<��<?��<��<��<ME�<��<���<�~�<�4�<���<a��<�?�<���<���<�(�<�ÿ<_[�<��<�~�< �<z��<J�<o��<#�<8��<��<D{�<L�<X�<���<$(�<���<%�<�I�<���<���<�R�<���<g��<�D�<��<9ۖ<V#�<�i�<���<���<�1�<dq�<���<��<i(�<$c�<ל�<�Ձ<��<��|<��x<	fu<��q<�>n<��j<dg<��c<"�_<`\\<��X<�9U<B�Q<9N<�J<�G<�}C<��?<�t<<A�8<�v5<��1<�.<�+<��'<(8$<)� <pn<�<Y�<`c<M<��<Ȇ	<qH<1<���;�c�;E�;���;/��;Ņ�;�p�;�h�;^p�;Յ�;f��;�ݼ; �;r�;�ҫ;lC�;Pà;S�;e�;`��;`�;h.�;��;b�w;�m;d;@Z;ٖP;G;,�=;�M4;O+;/";�;�.;ul;>��:Er�:|��:2��:F\�:��:��:#��:Zqt:�BU:zi6:��:�`�9���9��x9�~9��v7�OǸ̤U�nP��V۹On	���$��L@��l[�RWv�/����Ε��������7��mʺ��ֺ���{u� ������&�0h�g��"��$�70*��U0�zv6��<�
�B���H�"�N���T�1�Z�a��g��m��s�%y�7,�̙��F�������������������T���,����ǚ��  �  �f=#=t�=�A=a�=�|===8� =�S =R��<�<0O�<[��<���<��<�"�<�T�<*��<M��<T��<�<�?�<�j�<l��<���<s��<��<9,�<N�</n�<}��<��<]��<���<)��<c�<m�<)(�<�5�<�@�<�H�<�N�< R�<�R�<�P�<kK�<�C�<�8�<�*�<��<Q�<���<��<��<o��<}n�<�E�<��<@��<���<��<GE�<��<���<�~�<�4�<���<m��<@�<���<���<�(�<�ÿ<a[�< �<�~�<�
�<p��<F�<y��<%�<F��<��<B{�<Q�<X�<���<(�<���<�<�I�<���<���<�R�<���<g��<�D�<��<Aۖ<R#�<�i�<�<���<�1�<jq�<���<��<f(�<c�<䜃<�Ձ<��<�|<��x<fu<��q<�>n<��j<`g<��c<'�_<m\\<��X<�9U<0�Q<<N<�J<�G<�}C<��?<�t<<4�8<�v5<��1<�.<�+<y�'<#8$<6� <�n<�<W�<Gc<D<��<��	<H<<Ļ�;�c�;J�;��;6��;���;xp�;<i�;lp�;���;\��;�ݼ; �;�q�;�ҫ;uC�;�à;"S�;J�;t��;<`�;�.�;t�;s�w;��m;�d;�?Z;��P;G;ɝ=;�M4;;+;�";6;�.;�l;f��:Zr�:#��:	��:3\�:	�:��:i��:�rt:�CU:Yj6:M�:N`�9W��9��x9��9�Av7�TǸ��U��Q���S۹n	���$��M@�9m[��Vv�l���Ε�����������$ʺ�ֺҸ㺘u�~!������&��g�(��@��?$��0*��U0��v6���<�*�B� �H�>�N���T���Z�� a��g�6m�Gs��$y�,�����q�������祋�쪎�����:��������ǚ��  �  �f=F=��=�A=��=D}=�=�� =7T =��<��<"P�<k��<���<-��<�#�<(V�<���<���<���<��<-A�<Xl�<?��<{��<q��<�
�<G.�<RP�<sp�<��<^��<���<y��<���<F	�<T�<:+�<�8�<�C�<KL�<KR�<�U�<CV�<;T�<9O�<gG�<�<�<�.�<��<�	�<,��<z��<���<
��<s�<�J�<��<%��<ֻ�<��<:J�<��<���<���<�9�<��<���<E�<���<͎�<�-�<ɿ<``�<��<ʃ�<��<K��<�<5��<��<ޕ�<i�<��<��<;\�<�Ū<,�<~��<��<gM�<'��<D �<�U�<˨�<p��<�G�<œ�<�ݖ<�%�<�k�<��<��<�3�<s�<*��<�<�)�<;d�<ٝ�<�ց<��<��|<��x<�fu<��q<>n<��j<�g<h�c<��_<�Z\<��X<�7U<��Q<wN<��J<AG<�yC<��?<Vp<<}�8<�q5<U�1<^�.<�+<f�'<�1$<g� <�g<M	< �<�[<I<��<1~	<�?<<���;�P�;@�;u��;���;�q�;�[�;^T�;[�;rp�;���;�Ǽ;�	�;H[�;w��;�,�;֬�;T<�;�ە;���;I�;��;���;�w;��m;�c;�Z;7jP;w�F;\r=;�#4;7�*;��!;��;3;;E;=�:&�:pB�:���:0�:�Ʃ:^��:۸�:L�s:|�T:"�5:bl:t�9.��9�w9�9��[7�uʸv0W����d	ܹ��	�!N%�!�@�h�[���v�������K ���6��w;��+ʺ	׺��㺏��:����k2��r���d��$�>9*��]0��~6�ښ<�޳B���H��N���T�b�Z��a�g��m��s�'y�l.�i���"�������,���Ȫ��q�������%���*ǚ��  �  �f=M=��=�A=��=?}=�=�� ==T =��<�<P�<Y��<ǻ�<7��<�#�<V�<~��<���<���<��<4A�<]l�<2��<���<e��<�
�<T.�<EP�<xp�<َ�<Z��<���<~��<���<G	�<^�<3+�<�8�<�C�<BL�<CR�<�U�<OV�<3T�<EO�<fG�<�<�<�.�<��<�	�</��<���<o��<��<#s�<�J�<��<��<��<��<IJ�<��<���<���<�9�<��<���<%E�<���<���<�-�<�ȿ<c`�< ��<Ӄ�<��<U��<�<0��<��<Ε�<m�<��<��<<\�<�Ū<,�<r��<��<oM�<5��<M �<�U�<Ψ�<_��<�G�<ѓ�<�ݖ<�%�<�k�<��<��<�3�< s�<2��<�<�)�<<d�<ӝ�<�ց<��<�|<��x<jfu<��q<u>n<�j<�g<|�c<��_<�Z\<u�X<c7U<��Q<UN<ӌJ<5G<�yC<��?<@p<<��8<�q5<j�1<[�.<�+<M�'<�1$<�� <�g<i	<ܯ<�[<U<��<M~	<�?<$<[��;�P�;�;f��;*��;{q�;�[�;#T�;�Z�;ap�;���;�Ǽ;�	�;o[�;\��;�,�;���;2<�;}ە;���;GI�;��;���;�w;��m;^�c;�Z;�jP;��F;�r=;�"4;�*;�!;,�;A;�D;�=�:C&�:aC�:<��:��:�Ʃ:�:ù�:5�s:��T:h�5:�j:s�9(��9gw9��9�1\7�rʸ�+W�2���
ܹ��	�)P%���@��[�ޣv�������P��O7��;;���*ʺ'׺���B��c:�����2�ar�Y������$��8*��]0�-~6���<���B�#�H���N���T���Z�Fa��g�om�I s��'y�V.�~���	���ϡ�����Ϫ��t����]���ǚ��  �  �f=T=��=�A=��=:}=�=�� =>T =��<�<P�<Z��<ͻ�<&��<�#�<V�<���<���<���<��<(A�<dl�<'��<���<^��<�
�<^.�<<P�<�p�<َ�<h��<���<v��<���<>	�<c�<)+�<�8�<�C�<OL�<NR�<�U�<ZV�<&T�<JO�<aG�<�<�<�.�<��<�	�< ��<���<q��<��<!s�<�J�<��<��<��<���<BJ�<��<���<���<�9�<��<}��</E�<���<Ȏ�<�-�< ɿ<o`�<��<Ճ�<��<Q��<�<+��<��<͕�<}�<��<��<A\�<�Ū<#,�<h��<��<dM�<+��<D �<�U�<֨�<]��<�G�<���<�ݖ<�%�<�k�<!��<��<�3�<s�<4��<��<�)�<:d�<˝�<�ց<��<�|<��x<zfu<��q<a>n<�j<�g<��c<��_<�Z\<��X<f7U<��Q<=N<�J<+G<�yC<��?<.p<<��8<�q5<m�1<?�.<�+<Y�'<�1$<�� <|g<u	<ܯ<�[<M<u�<A~	<�?<2<.��;�P�;��;g��;S��;Xq�;\�;$T�;)[�;\p�;���;�Ǽ;�	�;�[�;3��;�,�;���;c<�;�ە;z��;rI�;z�;���;��w;��m;:�c;XZ;~jP;�F;�r=;�"4;W�*;��!;��;�;�D;3>�:]%�:�B�::��:4�:�Ʃ:x��:W��:��s:��T:��5:�k:�v�9���9�
w9N�9�;\7d{ʸZ-W�Y��ܹ�	�6P%���@�}�[���v�=���.�y���7���:��C+ʺ�׺���ŏ��9������1��r�E�����t$��8*�<^0�%~6��<���B�[�H���N���T���Z��a��g��m�2 s�T'y�.�����񝅻案���������S�������Y����ƚ��  �  �f=L=��=�A=��=<}=�=�� =AT =��<��< P�<_��<»�<)��<�#�<V�<���<���<���<��<)A�<fl�<.��<���<h��<�
�<N.�<CP�<zp�<׎�<`��<���<z��<���<C	�<d�<1+�<�8�<�C�<AL�<HR�<�U�<OV�<3T�<CO�<eG�<�<�<�.�<��<�	�<-��<��<|��<
��<s�<�J�<��<��<ݻ�<��<JJ�<��<���<���<�9�<��<���<%E�<���<Ď�<�-�< ɿ<e`�<��<փ�<��<Q��<�<-��<��<Ε�<n�<��<��<=\�<�Ū<,�<p��<��<fM�<1��<O �<�U�<Ϩ�<h��<�G�<Ó�<�ݖ<�%�<�k�<��<��<�3�<s�<6��< �<�)�<:d�<ӝ�<�ց<��<�|<��x<{fu<��q<n>n<�j<�g<��c<��_<�Z\<��X<X7U<��Q<PN<όJ<7G<�yC<��?<8p<<��8<�q5<|�1<[�.<�+<a�'<�1$<}� <�g<_	<�<�[<H<��<M~	<�?<6<J��;�P�;�;l��;��;uq�;�[�;T�;[�;Xp�;���;�Ǽ;�	�;�[�;T��;�,�;���;,<�;�ە;t��;EI�;��;���;�w;��m;U�c;�Z;�jP;{�F;�r=;Z#4;7�*;��!;��;[;E;x=�:&�:gC�:���:b�:ǩ:騙:ǹ�:0�s:��T:��5:]k:�r�9���9�w97�9�G\7�vʸ�-W�����ܹ%�	�P%���@�ڻ[�|�v�|�����V��q7���:��!+ʺh׺��㺝��L:��G��/2��r�������1$�9*��]0��}6��<���B�>�H���N���T���Z�Pa��g�Qm�q s�R'y�^.�����񝅻ʡ������䪎�t���ɶ��s����ƚ��  �  �f=H=��=�A=��=?}=�=�� =6T =!��<��<P�<[��<���<C��<�#�<V�<x��<���<���<��<.A�<[l�<8��<���<i��<�
�<L.�<TP�<up�<��<Y��<���<|��<���<D	�<V�<:+�<�8�<�C�<@L�<JR�<�U�<HV�<;T�<<O�<lG�<�<�<�.�<��<�	�<7��<|��<z��<���<$s�<�J�<��<��<ػ�<��<<J�<��<���<���<�9�<��<���<E�<���<ʎ�<�-�<ɿ<^`�<��<̃�<��<N��<�<2��<��<ە�<j�<��<��<:\�<�Ū<,�<z��<��<iM�<*��<G �<�U�<ƨ�<h��<�G�<ړ�<�ݖ<�%�<�k�<��<��<�3�<s�<2��<�<�)�<6d�<؝�<�ց<��<�|<��x<yfu<��q<�>n<��j<�g<i�c<��_<�Z\<��X<o7U<��Q<pN<��J<;G<�yC<��?<Cp<<��8<�q5<Q�1<c�.<�+<R�'<�1$<x� <�g<V	<�<{[<R<��<8~	<�?<!<s��;�P�;�;g��;��;�q�;�[�;RT�;�Z�;bp�;���;�Ǽ;�	�;Q[�;y��;�,�;Ȭ�;+<�;�ە;���;)I�;��;���;C�w;��m;H�c;�Z;0jP;��F;jr=;H#4;��*;�!;Q�;;
E;"=�:�&�:�B�:���:n�:�Ʃ:r��:K��:B�s:��T:�5:l:Lr�9\��9�w9��9��[7�vʸ�.W����D
ܹ*�	��N%���@�"�[�I�v�����B񕺡���6��d;���*ʺ�׺d��8���:��H��X2�r�������e$�9*��]0��~6�Ú<���B�%�H���N���T�k�Z��a�.g�jm�< s�X'y�z.�^���/���ϡ��)�������}���ض��F���ǚ��  �  �f=M=��=�A=��==}=�=�� =:T =��<�<P�<d��<���<+��<�#�<"V�<���<���<���<��<2A�<^l�<0��<���<a��<�
�<R.�<@P�<tp�<ߎ�<a��<���<t��<���<F	�<X�<3+�<�8�<�C�<FL�<BR�<�U�<NV�<2T�<@O�<jG�<�<�<�.�<��<�	�<1��<���<y��<��<s�<�J�<��<��<��<��<AJ�<��<���<���<�9�<��<���<#E�<���<���<�-�<ɿ<e`�<��<̃�<��<N��<
�<2��<��<֕�<k�<��<��<?\�<�Ū<,�<q��<��<lM�<.��<G �<�U�<Ϩ�<i��<�G�<Ó�<�ݖ<�%�<�k�<��<��<�3�<s�</��<�<�)�<6d�<՝�<�ց<��<�|<��x<xfu<��q<y>n<��j<�g<m�c<��_<�Z\<��X<p7U<��Q<JN<ӌJ<:G<�yC<��?<;p<<��8<�q5<_�1<^�.<�+<\�'<�1$<s� <�g<S	<��<�[<^<��<@~	<�?<&<S��;�P�;��;{��;#��;fq�;�[�;=T�;[�;sp�;}��;�Ǽ;�	�;X[�;\��;�,�;���;?<�;|ە;{��;CI�;��;���;.�w;��m;N�c;�Z;ajP;��F;�r=;@#4;*�*;��!;��;2;�D;�=�:K&�:�B�:ޒ�:��:�Ʃ:'��:���:��s:p�T:q�5:�j:�s�9$��9�w9��9��[7�uʸ�.W�	��>
ܹ	�	�%O%��@���[��v�V�������U7��;���*ʺ�׺d����D:��:��[2��r�������X$��8*��]0�f~6���<���B�5�H���N���T���Z�Ka��g�~m�' s�['y�3.�v����������"���ݪ��\���϶��E���ǚ��  �  �f=N=��=�A=��==}=�=�� =?T =��<��<P�<`��<Ļ�<3��<�#�<V�<}��<���<���<��<(A�<il�<*��<���<a��<�
�<S.�<BP�<�p�<֎�<]��<���<|��<���<B	�<f�</+�<�8�<�C�<KL�<FR�<�U�<VV�<,T�<HO�<`G�<�<�<�.�<��<�	�<(��<���<t��<��<s�<�J�<��<��<��<��<JJ�<��<���<���<�9�<��<���<*E�<���<�<�-�<�ȿ<h`�<��<ڃ�<��<P��<�<,��<��<˕�<z�<��<��<@\�<�Ū<,�<j��<��<cM�<1��<K �<�U�<ͨ�<f��<�G�<˓�<�ݖ<�%�<�k�<��<��<�3�<s�<4��<�<�)�<;d�<͝�<�ց<��<��|<��x<jfu<��q<q>n<�j<�g<�c<��_<�Z\<w�X<a7U<��Q<LN<،J<0G<�yC<��?<;p<<��8<�q5<t�1<R�.<�+<V�'<�1$<�� <�g<e	<�<�[<J<��<L~	<�?<<<:��;�P�; �;u��;(��;nq�;�[�;T�;�Z�;\p�;���;�Ǽ;�	�;�[�;L��;�,�;���;S<�;�ە;y��;bI�;��;���;��w;��m;E�c;�Z;�jP;T�F;�r=;#4;K�*;��!;
�;z;�D;�=�:�%�:rC�:���:6�:=ǩ:���:	��:�s:M�T:>�5:k:�u�9ޭ�9_w9��9�g\7Fwʸ.W����ܹ1�	�}P%��@� �[�ѣv�I���������7��n:��Q+ʺi׺#�㺤��k:��Y��2��r�v�����d$��8*��]0��}6��<���B��H���N���T���Z�$a��g�7m�@ s��'y�H.���������ա������۪��m���궔�a����ƚ��  �  �f=I=��=�A=��=?}=�=�� =9T = ��<�<P�<]��<���<=��<�#�<#V�<��<���<���<��<&A�<bl�<1��<���<j��<�
�<P.�<JP�<vp�<ߎ�<a��<���<|��<���<:	�<[�<3+�<�8�<�C�<EL�<FR�<�U�<LV�<4T�<BO�<bG�<�<�<�.�<��<�	�<2��<���<{��<��<s�<�J�<��<��<ݻ�<���<>J�<��<���<���<�9�<��<���<"E�<���<Ǝ�<�-�<ɿ<i`�<��<Ѓ�<��<L��<�<0��<��<ԕ�<m�<��<��<=\�<�Ū<,�<p��<��<cM�<,��<H �<�U�<̨�<j��<�G�<ѓ�<�ݖ<�%�<�k�<��<��<�3�<s�<3��<�<�)�<<d�<ӝ�<�ց<��<�|<��x<~fu<��q<y>n<�j<�g<q�c<��_<�Z\<��X<i7U<��Q<dN<ŌJ<4G<�yC<��?<Bp<<��8<�q5<\�1<b�.<�+<`�'<�1$<p� <�g<O	<��<�[<Y<��<=~	<�?</<W��;�P�;"�;h��;��;�q�;�[�;=T�;[�;dp�;���;�Ǽ;�	�;d[�;Z��;�,�;���;=<�;�ە;���;:I�;��;���;��w;��m;D�c;mZ;PjP;��F;�r=;O#4;�*;��!;�;;E;�=�:e&�:�B�:l��:R�:�Ʃ:Ҩ�:���:��s:M�T:��5:�k:�s�9ϯ�9�w9��9�\7�}ʸ�/W�����
ܹ��	�gO%���@�>�[��v�����]�G��d7���:��K+ʺ�׺W����:��3��m2�`r�������8$��8*��]0�t~6���<���B��H���N���T���Z�ta�Og�sm�G s�C'y�'.�u�������������̪��a���Ŷ��R���ǚ��  �  �f=J=��=�A=��=?}=�=�� =;T =!��< �<P�<f��<���<5��<�#�<)V�<v��<���<���<��<6A�<Zl�<6��<���<g��<�
�<R.�<FP�<np�<��<X��<���<r��<���<P	�<[�<2+�<�8�<�C�<DL�<AR�<�U�<GV�<<T�<:O�<mG�<�<�<�.�<��<�	�<7��<z��<|��<��<s�<�J�<��<#��<ջ�<���<:J�<��<���<���<�9�<��<���<E�<���<���<�-�<ɿ<_`�<��<̃�<��<U��<�<0��<��<ە�<g�<��<��<<\�<�Ū<,�<y��<��<nM�<1��<C �<�U�<Ũ�<q��<�G�<͓�<�ݖ<�%�<�k�<��<��<�3�<)s�<,��<�<�)�<2d�<ڝ�<�ց<��<�|<��x<pfu<��q<m>n<�j<�g<u�c<��_<�Z\<y�X<n7U<��Q<[N<ɌJ<@G<�yC<��?<Ap<<�8<�q5<b�1<d�.<�+<Q�'<�1$<p� <�g<E	<�<x[<\<��<C~	<�?<<m��;�P�;�;k��;$��;�q�;�[�;OT�;�Z�;ap�;v��;�Ǽ;"
�;c[�;X��;�,�;���;9<�;yە;���;&I�;��;���;H�w;��m;8�c;�Z;BjP;��F;ar=;Y#4;�*;��!;
�; ;'E;=�:�&�:lB�:5��:{�:�Ʃ:���:B��:9�s:��T:��5:�j:�r�9���9�w9��9~�[7?mʸ�+W�����
ܹ�	��N%�s�@���[�أv�����R񕺆���6��`;���*ʺ_׺������:������2�}r�������h$�
9*��]0�`~6�R�<�ͳB�(�H���N���T�[�Z��a�ug��m�- s�{'y�k.�����������������y���趔�G���(ǚ��  �  �f=N=��=�A=��=>}=�=�� ==T =��<�<P�<^��<Ż�<6��<�#�<V�<z��<���<���<��<(A�<bl�</��<���<a��<�
�<U.�<CP�<�p�<ێ�<Z��<���<y��<���<:	�<a�<2+�<�8�<�C�<ML�<FR�<�U�<RV�<2T�<@O�<gG�<�<�<�.�<��<�	�<+��<���<v��<	��<s�<�J�<��<��<ݻ�<��<=J�<��<���<���<�9�<��<���<'E�<���<�<�-�<�ȿ<f`�<��<փ�<��<M��<�<4��<��<Е�<y�<��<��<>\�<�Ū<,�<q��<��<bM�<1��<B �<�U�<ʨ�<g��<�G�<͓�<�ݖ<�%�<�k�<��<��<�3�<s�<0��<�<�)�<3d�<ѝ�<�ց<��<��|<��x<hfu<��q<r>n<�j<�g<|�c<��_<�Z\<v�X<k7U<��Q<PN<،J<1G<�yC<��?<=p<<��8<�q5<j�1<K�.<�+<S�'<�1$<�� <�g<f	<�<�[<Y<w�<G~	<�?</<P��;�P�; �;c��;0��;rq�;�[�;,T�;�Z�;zp�;���;�Ǽ;�	�;y[�;X��;�,�;���;_<�;�ە;���;OI�;��;���;�w;��m;�c;�Z;_jP;l�F;�r=;(#4;,�*;��!;�;[;�D;}=�:&�:�B�:���:�:�Ʃ:��:���:�s:��T:��5:k:�u�9���9)w9��9]D\7�|ʸ�/W�����	ܹ��	��O%�,�@��[���v�r�������_7���:��b+ʺj׺���S��:��L��2�~r�v�����n$��8*��]0�?~6�ۚ<���B�'�H���N���T���Z�.a��g�*m� s��'y� .���������������ݪ��W�����M����ƚ��  �  �f=M=��=�A=��=;}=�=�� =ET =��<	�<P�<Z��<ƻ�</��<�#�<V�<���<���<���<��<"A�<ol�<&��<���<d��<�
�<R.�<>P�<~p�<͎�<h��<���<x��<���<8	�<g�<&+�<�8�<�C�<DL�<AR�<�U�<PV�<)T�<MO�<\G�<�<�<�.�<��<�	�<*��<���<s��<��<s�<�J�<��<��<��<��<NJ�<��<���<���<�9�< ��<���<%E�<���<���<�-�<�ȿ<p`�<��<ڃ�<��<T��<�<)��<��<Õ�<r�<��<��<;\�<�Ū<,�<e��<��<aM�<9��<N �<�U�<ը�<_��<�G�<Ǔ�<�ݖ<�%�<�k�<!��<��<�3�<s�<@��< �<�)�<Bd�<ʝ�<�ց<��<��|<��x<sfu<��q<a>n<%�j<�g<��c<��_<�Z\<��X<O7U<��Q<LN<ӌJ<&G<�yC<��?<3p<<��8<�q5<��1<W�.<�+<`�'<�1$<�� <�g<e	<ܯ<�[<Y<��<_~	<�?<I<-��;�P�;�;Y��;%��;_q�;�[�;�S�;)[�;Rp�;���;�Ǽ;�	�;�[�;)��;�,�;���;8<�;wە;|��;JI�;��;���;��w;��m;��c;{Z;�jP;f�F;�r=;#4; �*;��!;��;K;�D;!>�:�%�:�C�:В�:��:�ǩ:D��:b��:�s:��T:,�5:oj:�s�9C��9Jw9��9j\7�|ʸ,W����ܹ��	�~Q%���@�ż[��v������񕺵��!8��-:��k+ʺ�׺���H���9�����2��r�m�����\$��8*��]0��}6��<�/�B�=�H���N�~�T���Z�?a��g�[m�� s�p'y�.�����ϝ�����٥������_���Ƕ�������ƚ��  �  �f=K=��=�A=��=>}=�=�� =;T =��<��<P�<d��<Ļ�<6��<�#�< V�<{��<���<���<��<*A�<cl�<0��<���<a��<�
�<R.�<LP�<~p�<܎�<a��<���<t��<���<H	�<c�<)+�<�8�<�C�<LL�<LR�<�U�<KV�<3T�<@O�<fG�<�<�<�.�<��<�	�<+��<}��<y��<
��<#s�<�J�<��<��<ڻ�<��<>J�<��<���<���<�9�<��<���<"E�<���<̎�<�-�<ɿ<i`�<��<Ӄ�<��<U��<�<%��<��<ҕ�<w�<��<��<>\�<�Ū<,�<q��<��<fM�<,��<D �<�U�<ɨ�<i��<�G�<ϓ�<�ݖ<�%�<�k�<��<��<�3�<s�<4��<�<�)�<5d�<՝�<�ց<��<��|<��x<vfu<��q<`>n<�j<�g<��c<��_<�Z\<��X<i7U<��Q<eN<ʌJ<;G<�yC<��?<=p<<��8<�q5<e�1<U�.<�+<S�'<�1$<�� <�g<X	<�<�[<J<�<?~	<�?<1<S��;�P�; �;n��;$��;�q�;�[�;3T�;[�;<p�;~��;�Ǽ;
�;�[�;4��;�,�;���;Z<�;�ە;���;4I�;��;���;�w;��m;@�c;Z;VjP;i�F;yr=;A#4;:�*;�!;0�;N; E;P=�:�%�:�B�:~��:G�:�Ʃ:�:���:�s:P�T:B�5:Gl:�u�9���9�w9�92\7�rʸ]+W�����ܹ��	��O%�o�@���[���v�i��������\7���:��'+ʺ�׺��㺗��:��>��H2�pr�d�����g$�
9*��]0�K~6�˚<���B�/�H���N���T���Z�{a�Fg�?m�& s�e'y�J.�����ꝅ�ʡ��󥋻����z���ж��R����ƚ��  �  �f=G=��=�A=��=@}=�=�� =7T =(��<�<P�<d��<���<9��<�#�<'V�<x��<Ƿ�<���<��<8A�<Vl�<6��<���<^��<�
�<J.�<DP�<op�<܎�<T��<���<���<���<;	�<Y�<:+�<�8�<�C�<AL�<?R�<�U�<HV�<?T�<0O�<rG�<�<�<�.�<��<�	�<;��<��<~��<��<s�<�J�<��<"��<ػ�<���<@J�<��<���<���<�9�<��<���<!E�<���<���<�-�<�ȿ<_`�<��<σ�<��<H��<�<8��<��<ϕ�<g�<��<��<A\�<�Ū<,�<y��<��<oM�<1��<O �<�U�<Ũ�<p��<�G�<ϓ�<�ݖ<�%�<�k�<��<��<�3�<(s�<'��<�<�)�<'d�<㝃<�ց<��<݋|<��x<gfu<��q<�>n<��j<�g<f�c<��_<�Z\<p�X<k7U<��Q<WN<��J<RG<�yC<��?<Fp<<u�8<�q5<S�1<q�.<�+<W�'<�1$<j� <�g<M	<��<{[<j<��<;~	<�?<<m��;�P�;��;���;��;vq�;�[�;2T�;�Z�;�p�;���;�Ǽ;�	�;][�;x��;�,�;���;-<�;pە;���;*I�;��;���;m�w;��m;+�c;�Z;JjP;��F;�r=;i#4;��*;��!;�;;!E;.=�:�&�:�B�:I��:w�:~Ʃ:���:ø�:2�s:/�T:Z�5:�j:Mr�9���9�w9��9f\7�|ʸ�1W�����ܹb�	��O%�q�@��[���v�:����񕺓���6���;���*ʺf׺��㺦���:�� ���2�or�ͬ����F$��8*�t]0��~6�U�<���B��H�g�N�T�T��Z��a�yg��m�4 s��'y�.�[���"����0�������S�������M���)ǚ��  �  �f=K=��=�A=��=>}=�=�� =;T =��<��<P�<d��<Ļ�<6��<�#�< V�<{��<���<���<��<*A�<cl�<0��<���<a��<�
�<R.�<LP�<~p�<܎�<a��<���<t��<���<H	�<c�<)+�<�8�<�C�<LL�<LR�<�U�<KV�<3T�<@O�<fG�<�<�<�.�<��<�	�<+��<}��<y��<
��<#s�<�J�<��<��<ڻ�<��<>J�<��<���<���<�9�<��<���<"E�<���<̎�<�-�<ɿ<i`�<��<Ӄ�<��<U��<�<%��<��<ҕ�<w�<��<��<>\�<�Ū<,�<q��<��<fM�<,��<D �<�U�<ɨ�<i��<�G�<ϓ�<�ݖ<�%�<�k�<��<��<�3�<s�<4��<�<�)�<5d�<՝�<�ց<��<��|<��x<vfu<��q<`>n<�j<�g<��c<��_<�Z\<��X<i7U<��Q<eN<ʌJ<;G<�yC<��?<=p<<��8<�q5<e�1<U�.<�+<S�'<�1$<�� <�g<X	<�<�[<J<�<?~	<�?<1<S��;�P�; �;n��;$��;�q�;�[�;3T�;[�;<p�;~��;�Ǽ;
�;�[�;4��;�,�;���;Z<�;�ە;���;4I�;��;���;�w;��m;@�c;Z;VjP;i�F;yr=;A#4;:�*;�!;0�;N; E;P=�:�%�:�B�:~��:G�:�Ʃ:�:���:�s:P�T:B�5:Gl:�u�9���9�w9�92\7�rʸ]+W�����ܹ��	��O%�o�@���[���v�i��������\7���:��'+ʺ�׺��㺗��:��>��H2�pr�d�����g$�
9*��]0�K~6�˚<���B�/�H���N���T���Z�{a�Fg�?m�& s�e'y�J.�����ꝅ�ʡ��󥋻����z���ж��R����ƚ��  �  �f=M=��=�A=��=;}=�=�� =ET =��<	�<P�<Z��<ƻ�</��<�#�<V�<���<���<���<��<"A�<ol�<&��<���<d��<�
�<R.�<>P�<~p�<͎�<h��<���<x��<���<8	�<g�<&+�<�8�<�C�<DL�<AR�<�U�<PV�<)T�<MO�<\G�<�<�<�.�<��<�	�<*��<���<s��<��<s�<�J�<��<��<��<��<NJ�<��<���<���<�9�< ��<���<%E�<���<���<�-�<�ȿ<p`�<��<ڃ�<��<T��<�<)��<��<Õ�<r�<��<��<;\�<�Ū<,�<e��<��<aM�<9��<N �<�U�<ը�<_��<�G�<Ǔ�<�ݖ<�%�<�k�<!��<��<�3�<s�<@��< �<�)�<Bd�<ʝ�<�ց<��<��|<��x<sfu<��q<a>n<%�j<�g<��c<��_<�Z\<��X<O7U<��Q<LN<ӌJ<&G<�yC<��?<3p<<��8<�q5<��1<W�.<�+<`�'<�1$<�� <�g<e	<ܯ<�[<Y<��<_~	<�?<I<-��;�P�;�;Y��;%��;_q�;�[�;�S�;)[�;Rp�;���;�Ǽ;�	�;�[�;)��;�,�;���;8<�;wە;|��;JI�;��;���;��w;��m;��c;{Z;�jP;f�F;�r=;#4; �*;��!;��;K;�D;!>�:�%�:�C�:В�:��:�ǩ:D��:b��:�s:��T:,�5:oj:�s�9C��9Jw9��9j\7�|ʸ,W����ܹ��	�~Q%���@�ż[��v������񕺵��!8��-:��k+ʺ�׺���H���9�����2��r�m�����\$��8*��]0��}6��<�/�B�=�H���N�~�T���Z�?a��g�[m�� s�p'y�.�����ϝ�����٥������_���Ƕ�������ƚ��  �  �f=N=��=�A=��=>}=�=�� ==T =��<�<P�<^��<Ż�<6��<�#�<V�<z��<���<���<��<(A�<bl�</��<���<a��<�
�<U.�<CP�<�p�<ێ�<Z��<���<y��<���<:	�<a�<2+�<�8�<�C�<ML�<FR�<�U�<RV�<2T�<@O�<gG�<�<�<�.�<��<�	�<+��<���<v��<	��<s�<�J�<��<��<ݻ�<��<=J�<��<���<���<�9�<��<���<'E�<���<�<�-�<�ȿ<f`�<��<փ�<��<M��<�<4��<��<Е�<y�<��<��<>\�<�Ū<,�<q��<��<bM�<1��<B �<�U�<ʨ�<g��<�G�<͓�<�ݖ<�%�<�k�<��<��<�3�<s�<0��<�<�)�<3d�<ѝ�<�ց<��<��|<��x<hfu<��q<r>n<�j<�g<|�c<��_<�Z\<v�X<k7U<��Q<PN<،J<1G<�yC<��?<=p<<��8<�q5<j�1<K�.<�+<S�'<�1$<�� <�g<f	<�<�[<Y<w�<G~	<�?</<P��;�P�; �;c��;0��;rq�;�[�;,T�;�Z�;zp�;���;�Ǽ;�	�;y[�;X��;�,�;���;_<�;�ە;���;OI�;��;���;�w;��m;�c;�Z;_jP;l�F;�r=;(#4;,�*;��!;�;[;�D;}=�:&�:�B�:���:�:�Ʃ:��:���:�s:��T:��5:k:�u�9���9)w9��9]D\7�|ʸ�/W�����	ܹ��	��O%�,�@��[���v�r�������_7���:��b+ʺj׺���S��:��L��2�~r�v�����n$��8*��]0�?~6�ۚ<���B�'�H���N���T���Z�.a��g�*m� s��'y� .���������������ݪ��W�����M����ƚ��  �  �f=J=��=�A=��=?}=�=�� =;T =!��< �<P�<f��<���<5��<�#�<)V�<v��<���<���<��<6A�<Zl�<6��<���<g��<�
�<R.�<FP�<np�<��<X��<���<r��<���<P	�<[�<2+�<�8�<�C�<DL�<AR�<�U�<GV�<<T�<:O�<mG�<�<�<�.�<��<�	�<7��<z��<|��<��<s�<�J�<��<#��<ջ�<���<:J�<��<���<���<�9�<��<���<E�<���<���<�-�<ɿ<_`�<��<̃�<��<U��<�<0��<��<ە�<g�<��<��<<\�<�Ū<,�<y��<��<nM�<1��<C �<�U�<Ũ�<q��<�G�<͓�<�ݖ<�%�<�k�<��<��<�3�<)s�<,��<�<�)�<2d�<ڝ�<�ց<��<�|<��x<pfu<��q<m>n<�j<�g<u�c<��_<�Z\<y�X<n7U<��Q<[N<ɌJ<@G<�yC<��?<Ap<<�8<�q5<b�1<d�.<�+<Q�'<�1$<p� <�g<E	<�<x[<\<��<C~	<�?<<m��;�P�;�;k��;$��;�q�;�[�;OT�;�Z�;ap�;v��;�Ǽ;"
�;c[�;X��;�,�;���;9<�;yە;���;&I�;��;���;H�w;��m;8�c;�Z;BjP;��F;ar=;Y#4;�*;��!;
�; ;'E;=�:�&�:lB�:5��:{�:�Ʃ:���:B��:9�s:��T:��5:�j:�r�9���9�w9��9~�[7?mʸ�+W�����
ܹ�	��N%�s�@���[�أv�����R񕺆���6��`;���*ʺ_׺������:������2�}r�������h$�
9*��]0�`~6�R�<�ͳB�(�H���N���T�[�Z��a�ug��m�- s�{'y�k.�����������������y���趔�G���(ǚ��  �  �f=I=��=�A=��=?}=�=�� =9T = ��<�<P�<]��<���<=��<�#�<#V�<��<���<���<��<&A�<bl�<1��<���<j��<�
�<P.�<JP�<vp�<ߎ�<a��<���<|��<���<:	�<[�<3+�<�8�<�C�<EL�<FR�<�U�<LV�<4T�<BO�<bG�<�<�<�.�<��<�	�<2��<���<{��<��<s�<�J�<��<��<ݻ�<���<>J�<��<���<���<�9�<��<���<"E�<���<Ǝ�<�-�<ɿ<i`�<��<Ѓ�<��<L��<�<0��<��<ԕ�<m�<��<��<=\�<�Ū<,�<p��<��<cM�<,��<H �<�U�<̨�<j��<�G�<ѓ�<�ݖ<�%�<�k�<��<��<�3�<s�<3��<�<�)�<<d�<ӝ�<�ց<��<�|<��x<~fu<��q<y>n<�j<�g<q�c<��_<�Z\<��X<i7U<��Q<dN<ŌJ<4G<�yC<��?<Bp<<��8<�q5<\�1<b�.<�+<`�'<�1$<p� <�g<O	<��<�[<Y<��<=~	<�?</<W��;�P�;"�;h��;��;�q�;�[�;=T�;[�;dp�;���;�Ǽ;�	�;d[�;Z��;�,�;���;=<�;�ە;���;:I�;��;���;��w;��m;D�c;mZ;PjP;��F;�r=;O#4;�*;��!;�;;E;�=�:e&�:�B�:l��:R�:�Ʃ:Ҩ�:���:��s:M�T:��5:�k:�s�9ϯ�9�w9��9�\7�}ʸ�/W�����
ܹ��	�gO%���@�>�[��v�����]�G��d7���:��K+ʺ�׺W����:��3��m2�`r�������8$��8*��]0�t~6���<���B��H���N���T���Z�ta�Og�sm�G s�C'y�'.�u�������������̪��a���Ŷ��R���ǚ��  �  �f=N=��=�A=��==}=�=�� =?T =��<��<P�<`��<Ļ�<3��<�#�<V�<}��<���<���<��<(A�<il�<*��<���<a��<�
�<S.�<BP�<�p�<֎�<]��<���<|��<���<B	�<f�</+�<�8�<�C�<KL�<FR�<�U�<VV�<,T�<HO�<`G�<�<�<�.�<��<�	�<(��<���<t��<��<s�<�J�<��<��<��<��<JJ�<��<���<���<�9�<��<���<*E�<���<�<�-�<�ȿ<h`�<��<ڃ�<��<P��<�<,��<��<˕�<z�<��<��<@\�<�Ū<,�<j��<��<cM�<1��<K �<�U�<ͨ�<f��<�G�<˓�<�ݖ<�%�<�k�<��<��<�3�<s�<4��<�<�)�<;d�<͝�<�ց<��<��|<��x<jfu<��q<q>n<�j<�g<�c<��_<�Z\<w�X<a7U<��Q<LN<،J<0G<�yC<��?<;p<<��8<�q5<t�1<R�.<�+<V�'<�1$<�� <�g<e	<�<�[<J<��<L~	<�?<<<:��;�P�; �;u��;(��;nq�;�[�;T�;�Z�;\p�;���;�Ǽ;�	�;�[�;L��;�,�;���;S<�;�ە;y��;bI�;��;���;��w;��m;E�c;�Z;�jP;T�F;�r=;#4;K�*;��!;
�;z;�D;�=�:�%�:rC�:���:6�:=ǩ:���:	��:�s:M�T:>�5:k:�u�9ޭ�9_w9��9�g\7Fwʸ.W����ܹ1�	�}P%��@� �[�ѣv�I���������7��n:��Q+ʺi׺#�㺤��k:��Y��2��r�v�����d$��8*��]0��}6��<���B��H���N���T���Z�$a��g�7m�@ s��'y�H.���������ա������۪��m���궔�a����ƚ��  �  �f=M=��=�A=��==}=�=�� =:T =��<�<P�<d��<���<+��<�#�<"V�<���<���<���<��<2A�<^l�<0��<���<a��<�
�<R.�<@P�<tp�<ߎ�<a��<���<t��<���<F	�<X�<3+�<�8�<�C�<FL�<BR�<�U�<NV�<2T�<@O�<jG�<�<�<�.�<��<�	�<1��<���<y��<��<s�<�J�<��<��<��<��<AJ�<��<���<���<�9�<��<���<#E�<���<���<�-�<ɿ<e`�<��<̃�<��<N��<
�<2��<��<֕�<k�<��<��<?\�<�Ū<,�<q��<��<lM�<.��<G �<�U�<Ϩ�<i��<�G�<Ó�<�ݖ<�%�<�k�<��<��<�3�<s�</��<�<�)�<6d�<՝�<�ց<��<�|<��x<xfu<��q<y>n<��j<�g<m�c<��_<�Z\<��X<p7U<��Q<JN<ӌJ<:G<�yC<��?<;p<<��8<�q5<_�1<^�.<�+<\�'<�1$<s� <�g<S	<��<�[<^<��<@~	<�?<&<S��;�P�;��;{��;#��;fq�;�[�;=T�;[�;sp�;}��;�Ǽ;�	�;X[�;\��;�,�;���;?<�;|ە;{��;CI�;��;���;.�w;��m;N�c;�Z;ajP;��F;�r=;@#4;*�*;��!;��;2;�D;�=�:K&�:�B�:ޒ�:��:�Ʃ:'��:���:��s:p�T:q�5:�j:�s�9$��9�w9��9��[7�uʸ�.W�	��>
ܹ	�	�%O%��@���[��v�V�������U7��;���*ʺ�׺d����D:��:��[2��r�������X$��8*��]0�f~6���<���B�5�H���N���T���Z�Ka��g�~m�' s�['y�3.�v����������"���ݪ��\���϶��E���ǚ��  �  �f=H=��=�A=��=?}=�=�� =6T =!��<��<P�<[��<���<C��<�#�<V�<x��<���<���<��<.A�<[l�<8��<���<i��<�
�<L.�<TP�<up�<��<Y��<���<|��<���<D	�<V�<:+�<�8�<�C�<@L�<JR�<�U�<HV�<;T�<<O�<lG�<�<�<�.�<��<�	�<7��<|��<z��<���<$s�<�J�<��<��<ػ�<��<<J�<��<���<���<�9�<��<���<E�<���<ʎ�<�-�<ɿ<^`�<��<̃�<��<N��<�<2��<��<ە�<j�<��<��<:\�<�Ū<,�<z��<��<iM�<*��<G �<�U�<ƨ�<h��<�G�<ړ�<�ݖ<�%�<�k�<��<��<�3�<s�<2��<�<�)�<6d�<؝�<�ց<��<�|<��x<yfu<��q<�>n<��j<�g<i�c<��_<�Z\<��X<o7U<��Q<pN<��J<;G<�yC<��?<Cp<<��8<�q5<Q�1<c�.<�+<R�'<�1$<x� <�g<V	<�<{[<R<��<8~	<�?<!<s��;�P�;�;g��;��;�q�;�[�;RT�;�Z�;bp�;���;�Ǽ;�	�;Q[�;y��;�,�;Ȭ�;+<�;�ە;���;)I�;��;���;C�w;��m;H�c;�Z;0jP;��F;jr=;H#4;��*;�!;Q�;;
E;"=�:�&�:�B�:���:n�:�Ʃ:s��:K��:B�s:��T:�5:l:Lr�9\��9�w9��9��[7�vʸ�.W����D
ܹ*�	��N%���@�"�[�I�v�����B񕺡���6��d;���*ʺ�׺d��8���:��H��X2�r�������e$�9*��]0��~6�Ú<���B�%�H���N���T�k�Z��a�.g�jm�< s�X'y�z.�^���/���ϡ��)�������}���ض��F���ǚ��  �  �f=L=��=�A=��=<}=�=�� =AT =��<��< P�<_��<»�<)��<�#�<V�<���<���<���<��<)A�<fl�<.��<���<h��<�
�<N.�<CP�<zp�<׎�<`��<���<z��<���<C	�<d�<1+�<�8�<�C�<AL�<HR�<�U�<OV�<3T�<CO�<eG�<�<�<�.�<��<�	�<-��<��<|��<
��<s�<�J�<��<��<ݻ�<��<JJ�<��<���<���<�9�<��<���<%E�<���<Ď�<�-�< ɿ<e`�<��<փ�<��<Q��<�<-��<��<Ε�<n�<��<��<=\�<�Ū<,�<p��<��<fM�<1��<O �<�U�<Ϩ�<h��<�G�<Ó�<�ݖ<�%�<�k�<��<��<�3�<s�<6��< �<�)�<:d�<ӝ�<�ց<��<�|<��x<{fu<��q<n>n<�j<�g<��c<��_<�Z\<��X<X7U<��Q<PN<όJ<7G<�yC<��?<8p<<��8<�q5<|�1<[�.<�+<a�'<�1$<}� <�g<_	<�<�[<H<��<M~	<�?<6<J��;�P�;�;l��;��;uq�;�[�;T�;[�;Xp�;���;�Ǽ;�	�;�[�;T��;�,�;���;,<�;�ە;t��;EI�;��;���;�w;��m;U�c;�Z;�jP;{�F;�r=;Z#4;7�*;��!;��;[;E;x=�:&�:gC�:���:b�:ǩ:騙:ǹ�:0�s:��T:��5:]k:�r�9���9�w97�9�G\7�vʸ�-W�����ܹ%�	�P%���@�ڻ[�|�v�|�����V��q7���:��!+ʺh׺��㺝��L:��G��/2��r�������1$�9*��]0��}6��<���B�>�H���N���T���Z�Pa��g�Qm�q s�R'y�^.�����񝅻ʡ������䪎�t���ɶ��s����ƚ��  �  �f=T=��=�A=��=:}=�=�� =>T =��<�<P�<Z��<ͻ�<&��<�#�<V�<���<���<���<��<(A�<dl�<'��<���<^��<�
�<^.�<<P�<�p�<َ�<h��<���<v��<���<>	�<c�<)+�<�8�<�C�<OL�<NR�<�U�<ZV�<&T�<JO�<aG�<�<�<�.�<��<�	�< ��<���<q��<��<!s�<�J�<��<��<��<���<BJ�<��<���<���<�9�<��<}��</E�<���<Ȏ�<�-�< ɿ<o`�<��<Ճ�<��<Q��<�<+��<��<͕�<}�<��<��<A\�<�Ū<#,�<h��<��<dM�<+��<D �<�U�<֨�<]��<�G�<���<�ݖ<�%�<�k�<!��<��<�3�<s�<4��<��<�)�<:d�<˝�<�ց<��<�|<��x<zfu<��q<a>n<�j<�g<��c<��_<�Z\<��X<f7U<��Q<=N<�J<+G<�yC<��?<.p<<��8<�q5<m�1<?�.<�+<Y�'<�1$<�� <|g<u	<ܯ<�[<M<u�<A~	<�?<2<.��;�P�;��;g��;S��;Xq�;\�;$T�;)[�;\p�;���;�Ǽ;�	�;�[�;3��;�,�;���;c<�;�ە;z��;rI�;z�;���;��w;��m;:�c;XZ;~jP;�F;�r=;�"4;W�*;��!;��;�;�D;3>�:]%�:�B�::��:4�:�Ʃ:x��:W��:��s:��T:��5:�k:�v�9���9�
w9N�9�;\7d{ʸZ-W�Y��ܹ�	�6P%���@�}�[���v�=���.�y���7���:��C+ʺ�׺���ŏ��9������1��r�E�����t$��8*�<^0�%~6��<���B�[�H���N���T���Z��a��g��m�2 s�T'y�.�����񝅻案���������S�������Y����ƚ��  �  �f=M=��=�A=��=?}=�=�� ==T =��<�<P�<Y��<ǻ�<7��<�#�<V�<~��<���<���<��<4A�<]l�<2��<���<e��<�
�<T.�<EP�<xp�<َ�<Z��<���<~��<���<G	�<^�<3+�<�8�<�C�<BL�<CR�<�U�<OV�<3T�<EO�<fG�<�<�<�.�<��<�	�</��<���<o��<��<#s�<�J�<��<��<��<��<IJ�<��<���<���<�9�<��<���<%E�<���<���<�-�<�ȿ<c`�< ��<Ӄ�<��<U��<�<0��<��<Ε�<m�<��<��<<\�<�Ū<,�<r��<��<oM�<5��<M �<�U�<Ψ�<_��<�G�<ѓ�<�ݖ<�%�<�k�<��<��<�3�< s�<2��<�<�)�<<d�<ӝ�<�ց<��<�|<��x<jfu<��q<u>n<�j<�g<|�c<��_<�Z\<u�X<c7U<��Q<UN<ӌJ<5G<�yC<��?<@p<<��8<�q5<j�1<[�.<�+<M�'<�1$<�� <�g<i	<ܯ<�[<U<��<M~	<�?<$<[��;�P�;�;f��;*��;{q�;�[�;#T�;�Z�;ap�;���;�Ǽ;�	�;o[�;\��;�,�;���;2<�;}ە;���;GI�;��;���;�w;��m;^�c;�Z;�jP;��F;�r=;�"4;�*;�!;,�;A;�D;�=�:C&�:aC�:<��:��:�Ʃ:�:ù�:5�s:��T:h�5:�j:s�9(��9gw9��9�1\7�rʸ�+W�2���
ܹ��	�)P%���@��[�ޣv�������P��O7��;;���*ʺ'׺���B��c:�����2�ar�Y������$��8*��]0�-~6���<���B�#�H���N���T���Z�Fa��g�om�I s��'y�V.�~���	���ϡ�����Ϫ��t����]���ǚ��  �  g=�=��=%B=	�=�}==!� =�T =v��<e�<�Q�<��<|��<+��<�%�<FX�<���<��<A��<-�<�C�<2o�<8��<���<���<�<�1�<T�<;t�<��<���<8��<���<y��<�<9 �<I0�<�=�<2I�<�Q�<�W�<�[�<V\�<qZ�<�U�<�M�<?C�<|5�<�$�<��<t��<���<��<���<�z�<�R�<�&�<;��<���<0��<�R�<8�<��<��<KB�<���<%��<�M�<x��<R��<F6�<�ѿ<�h�<]��<��<�<^��<%�<��<�#�<���<��<	��<���<;c�<�̪<�2�<앧<��<oS�<���<��<)[�<���<i��<aL�<b��<�<�)�<�o�<���<���<�6�<�u�<���<`��<�+�<f�<o��<�ׁ<��<��|<��x<?gu<��q<">n<�j<Vg<|c<k�_<�W\<H�X<�3U<*�Q<�N<l�J<l�F<xsC<��?<
i<<��8<�i5<��1<"w.<+<-�'<,'$<L� <5\<7�<��<�N<��<´<	p	<21<.�<��;51�;*��;���;�s�;�O�;9�;n1�;�7�;~L�;p�;���;��;�5�;Ԗ�;��;��;�;m��;�d�;#�;��;�π;u{w;�vm;D�c;s�Y;� P;ݖF;*=;S�3;��*;��!;�;��;;���:æ�:?��:�:��:�Q�:�6�:4I�:ss:��S:z5:\�:���9A8�9�"t9��8dR07��ϸ��Y�fL��3:ݹ�Y
�$�%�>+A��=\�^"w�xꈺ�+���X���l��?o���\ʺ�8׺�N��Ed�����tE����������T$��G*�k0��6�i�<��B���H�Z�N�_�T�[��a�Ng�9m� %s��*y��1�ț��F���W�����������﯑�ʵ��
����Ś��  �  �f=�=��=%B=�=�}==%� =�T =z��<z�<�Q�<��<~��<��<�%�<:X�<���<��<I��<6�<�C�<8o�<(��<���<���<�<�1�<�S�<It�<Β�<r��<0��<���<���<�<H �<G0�<�=�<I�<�Q�< X�<[�<S\�<`Z�<�U�<�M�<>C�<�5�<�$�<��<x��<���<���<���<�z�<�R�<�&�<3��<��<6��<�R�<=�<��<��<HB�<���<��<�M�<h��<N��<F6�<rѿ<�h�<X��<��<"�<m��<%�<��<w#�<h��<��<���<���<-c�<�̪<�2�<ߕ�<��<wS�<��<��<7[�<���<^��<hL�<F��<�<�)�<�o�<���<���<�6�<�u�<ĳ�<U��<�+�<f�<a��<�ׁ<��<��|<��x<gu<��q<'>n<4�j<dg<�c<r�_<�W\<�X<3U<J�Q<zN<p�J<S�F<zsC<��?<�h<<��8<�i5<��1<,w.<F+<&�'<$'$<Q� <�[<D�<x�<�N<�<Ѵ<p	<C1<9�<���;1�;��;���;�s�;�O�;99�;1�;R7�;^L�;9p�; ��; �;6�;˖�;��;���;�;t��;Nd�;#�;��;�π;o{w;�vm;��c;��Y;� P;��F;�*=;�3;Ī*;C�!;��;��;�;���:$��:���:g�:���:�Q�:H6�:DJ�:gs:��S:�5:ء:��9�0�9�t9#�8��07��ϸ^�Y�^J���;ݹ�[
�[�%��)A�u?\��#w�b눺n,��mW���m���n��k\ʺ8׺n�n���c�����9E�����������$��F*��j0�Ɋ6�5�<���B�O�H�*�N�D�T��[��a��g��m�T%s��+y��1���������<���F����������5���J���sŚ��  �  �f=�=��=#B=�=�}==� =�T =i��<v�<�Q�<��<���<��<�%�</X�<���<��<=��<1�<�C�<Ao�<��<���<���<�<�1�<�S�<\t�<Ғ�<���<5��<���<���<��<G �<?0�<�=�<I�<�Q�<X�<|[�<i\�<XZ�<�U�<�M�<;C�<�5�<�$�<��<f��<���<���<���<�z�<�R�<�&�<'��<��<#��<�R�<1�<��<��<>B�<���<��<�M�<l��<Q��<V6�<wѿ<�h�<S��<��<�<c��<%�<��<�#�<j��<��<�<���<>c�<|̪<�2�<ӕ�<��<kS�<���<��<+[�<���<S��<~L�<E��<�<�)�<�o�<���<���<�6�<�u�<ͳ�<N��<�+�<f�<_��<�ׁ<��<��|<��x<#gu<��q<>n<4�j<8g<�c<_�_<�W\<4�X<�3U<h�Q<\N<��J<S�F<psC<��?<�h<<��8<�i5<��1<	w.<@+<�'<'$<w� <�[<q�<c�<�N<��<��<p	<(1<K�<{��;�1�;���;���;�s�;[O�;�9�;1�;�7�;rL�; p�;㢼;��;6�;���;�;���;F�;���;Bd�;h#�;i�;�π;5{w;rvm;��c;"�Y;� P;h�F;�*=;��3;��*;��!;��;D�;;��:���:���:��:Z��:�Q�:�5�:�J�:/s:q�S:5:*�:���9�1�9�(t9��8ڪ07o�ϸ�Y�;K���;ݹOY
�"�%�{'A��@\�z"w�Tꈺ�,���V��Zn��~n��$]ʺ�8׺��1���c��O���D���� ������$��F*�}k0��6�Ȧ<�B�B���H�'�N�^�T��[��a�]g�sm�%s�k+y�Z1�雂���������P���Ҫ��ׯ��񵔻6���7Ś��  �  �f=�=��=%B=�=�}==� =�T =v��<o�<�Q�<��<���<��<�%�<7X�<���<��<I��<?�<�C�<Co�<*��<���<���<�<�1�<�S�<Kt�<ђ�<}��<-��<���<���<�<K �<>0�<�=�<I�<�Q�<�W�<|[�<\\�<dZ�<�U�<�M�<CC�<�5�<�$�<��<p��<���<��<���<�z�<�R�<�&�<2��<��<,��<�R�<>�<��< ��<JB�<���<��<�M�<g��<M��<I6�<yѿ<�h�<R��<��<�<k��<%�<	��<#�<k��<��<���<���<<c�<�̪<�2�<���< ��<lS�<��<��<-[�<��<\��<nL�<G��<�<�)�<�o�<���<���<�6�<�u�<ʳ�<W��<�+�<f�<h��<�ׁ<��<��|<��x<'gu<��q<>n<>�j<Ig<�c<j�_<�W\<2�X<�3U<F�Q<vN<z�J<`�F<xsC<��?<�h<<��8<�i5<��1<#w.<1+<;�'<'$<[� <�[<R�<r�<�N<��<Ѵ<,p	<&1<P�<���;l1�;��;ĥ�;�s�;�O�;A9�;1�;~7�;TL�;8p�;���;��;&6�;���;��;���;�;m��;Bd�;3#�;��;�π;�{w;�vm;��c;v�Y;b!P;��F;�*=;�3;��*;_�!;��;��;�;��:���:���:u�:���:�Q�:g6�:�I�:�s:#�S:v5:��:���9a2�93 t9�
�8��07��ϸ��Y��I���<ݹ�Z
��%��)A��?\��#w�iꈺv,���W���m��]n��]ʺ�7׺:�	��Tc����
E����u�����B$�8G*�k0�V�6���<�V�B�:�H�'�N�J�T�U[�Oa�	g��m�E%s�\+y��1�ڛ��䞅�s���5��������������H���zŚ��  �  �f=�=��=%B=�=�}=="� =�T =u��<k�<�Q�<��<���<��<�%�<;X�<���<��<@��<2�<�C�<4o�<-��<���<���<�<�1�<�S�<Ct�<ޒ�<x��<3��<���<���<�<A �<Q0�<�=�<&I�<�Q�<X�<�[�<P\�<oZ�<�U�<�M�<6C�<�5�<�$�<��<r��<���< ��<���<�z�<�R�<�&�<5��<���<-��<�R�<7�<��<��<NB�<���<#��<�M�<o��<V��<L6�<�ѿ<�h�<b��<��<�<a��<%�<��<z#�<x��<��<��<���<6c�<�̪<�2�<啧<��<rS�<���<��<-[�<���<_��<lL�<Q��<�<�)�<�o�<���<���<�6�<�u�<���<R��<�+�<	f�<m��<�ׁ<��<��|<��x<(gu<��q<5>n<#�j<Mg<�c<��_<�W\<.�X<�3U<>�Q<�N<c�J<j�F<xsC<��?<�h<<��8<�i5<��1<!w.<)+<-�'<$'$<Y� <\<L�<y�<�N<��<��<p	<71<2�<���;^1�;��;���;�s�;�O�;"9�;Q1�;i7�;kL�;Cp�;֢�;��;�5�;�;��;↠;)�;���;rd�;#�;��;�π;�{w;Jvm;~�c;l�Y;� P;ǖF;>*=;�3;̪*;��!;؞;��;�;��:���:���:��:h��:'Q�:�6�:AI�:3s:��S:_5:Ѣ:[��95�9�t9��8F�07��ϸ'�Y�WJ���:ݹH[
�k�%�9*A�>\��#w��ꈺ�+��X��<m��8o���\ʺl8׺���;d�����E�.��s�����c$�nG*�k0��6�e�<���B�c�H�)�N�q�T�+[��a�yg��m�
%s�T+y��1��������j���g������������������Ś��  �  �f=�=��=B=�=�}==$� =�T =t��<z�<�Q�<��<���<��<�%�<:X�<���<��<C��<3�<�C�<4o�<.��<���<���<�<�1�<�S�<Gt�<ؒ�<z��<7��<���<���<
�<> �<H0�<�=�<I�<�Q�<�W�<�[�<^\�<cZ�<�U�<�M�<<C�<�5�<�$�<��<r��<���<���<���<�z�<�R�<�&�<1��<��<1��<�R�<8�<��<��<PB�<���<��<�M�<p��<H��<L6�<wѿ<�h�<\��<��< �<i��<%�<��<}#�<o��<��<���<���<:c�<|̪<�2�<啧<��<sS�<��<��<6[�<���<]��<sL�<G��<�<�)�<�o�<���<���<�6�<�u�<���<V��<�+�< f�<g��<�ׁ<��<��|<��x<gu<��q<>n<�j<cg<�c<g�_<�W\<%�X<�3U<<�Q<}N<��J<c�F<[sC<��?<�h<<��8<�i5<��1<w.<F+<�'<%'$<b� <�[<[�<y�<�N<�<Ŵ<p	<;1<1�<���;�1�;���;���;�s�;O�;29�;:1�;p7�;|L�;,p�;颼;��;�5�;Ζ�;��;���;&�;[��;dd�;;#�;��;�π;�{w;{vm;��c;{�Y;� P;͖F;�*=;��3;�*;f�!;��;�;�;���:ڦ�:���:�:���:pQ�:�6�:nI�:ys:Q�S:�5:�:M��92�9$!t9i�8iu07�ϸ:�Y�K���:ݹ�Z
�v�%��)A�M@\��"w��ꈺ�,���W��Am��!o���\ʺ>8׺��v���c������D����s������$��F*�#k0��6�G�<���B�D�H���N���T�^[�6a��g�m�!%s��+y��1�ӛ��*���>���t���ê��ᯑ����$����Ś��  �  �f=�=��=$B=�=�}== � =�T =q��<p�<�Q�<��<���<��<�%�<5X�<���<��<C��<=�<�C�<<o�<&��<���<���<�<�1�<�S�<Xt�<В�<}��</��<���<���<�<H �<=0�<�=�<I�<�Q�<X�<�[�<\\�<aZ�<�U�<�M�<@C�<�5�<�$�<��<i��<���<���<���<�z�<�R�<�&�<-��<��<&��<�R�<;�<��<��<FB�<���<��<�M�<m��<O��<X6�<qѿ<�h�<Q��<��<�<j��<%�<	��<�#�<g��<��<���<���<:c�<�̪<�2�<ܕ�<��<lS�<	��<��<*[�<���<W��<qL�<N��<�<�)�<�o�<���<���<�6�<�u�<ó�<T��<�+�<f�<e��<�ׁ<��<��|<��x<gu<��q<>n<6�j<Ng<�c<c�_<�W\<"�X<�3U<Y�Q<}N<z�J<^�F<vsC<��?<�h<<��8<�i5<��1<w.<3+<$�'<'$<e� <	\<X�<n�<�N<��<ƴ<)p	<,1<C�<���;�1�;���;���;�s�;�O�;v9�;1�;{7�;]L�;*p�;���;��;6�;���;��;���;O�;}��;Qd�;3#�;��;�π;h{w;�vm;��c;m�Y;L!P;�F;�*=;��3;�*;��!;̞;	�;�;���:$��:���:B�:Z��:�Q�:-6�:#J�:ms:�S:%5:�:x��9e0�9�"t9/	�8@�07v�ϸ̸Y�HJ���<ݹ�Z
���%��'A��?\�5#w��ꈺ�,��OW���m���n��]ʺ�7׺��<���c��.���D�F��R������$�1G*�Jk0�t�6��<���B�P�H�+�N�A�T�q[�Ka��g��m�%s��+y��1�䛂�����i���<���ʪ���������+���UŚ��  �  �f=�=��='B=	�=�}== � =�T =t��<p�<�Q�<��<|��<��<�%�<;X�<���<��<>��<2�<�C�<>o�<(��<���<���<�<�1�<�S�<Et�<֒�<���<0��<���<���<��<J �<C0�<�=�<!I�<�Q�<�W�<�[�<U\�<kZ�<�U�<�M�<@C�<�5�<�$�<��<q��<���<��<���<�z�<�R�<�&�<7��<��<-��<�R�<5�<��<��<EB�<���<��<�M�<q��<K��<N6�<|ѿ<�h�<V��<��<�<d��<%�<��<�#�<o��<��<���<���<7c�<�̪<�2�<ޕ�<��<pS�< ��<��<0[�<���<a��<fL�<T��<�<�)�<�o�<���<���<�6�<�u�<ȳ�<V��<�+�<f�<k��<�ׁ<��<��|<��x<*gu<��q<>n<:�j<<g<�c<k�_<�W\<7�X<�3U<9�Q<�N<l�J<h�F<�sC<��?<�h<<��8<�i5<��1< w.<3+<1�'<"'$<L� <\<?�<z�<�N<��<��<p	<31<F�<���;G1�;��;���;�s�;�O�;+9�;/1�;�7�;`L�;.p�;뢼;��;%6�;���;��;ˆ�;7�;e��;ld�;#�;��;�π;F{w;�vm;��c;P�Y;� P;��F;p*=;$�3;��*;��!;�;��;�;c��:���:���:��:���:�Q�:6�:|I�:�s:l�S:�5:z�:���9E3�9d#t9x�8�07R�ϸ��Y�5J��K<ݹ�Y
�x�%��)A�t?\�##w��ꈺ�+��>X���m���n���\ʺa8׺�ں��c�����HE���������V$�CG*�k0���6���<�j�B�D�H���N�3�T�@[��a��g�m�%s�O+y��1�қ��힅�����=����������뵔�#����Ś��  �  �f=�=��="B=�=�}==&� =�T =x��<s�<�Q�<��<~��<��<�%�<FX�<���<��<A��<9�<�C�<.o�<1��<���<���<�<�1�<�S�<Ht�<ؒ�<s��<6��<���<���<�<D �<E0�<�=�<I�<�Q�<�W�<�[�<S\�<kZ�<�U�<�M�<;C�<�5�<�$�<��<{��<���<��<���<�z�<�R�<�&�<<��<��<9��<�R�<C�<��<��<TB�<���<��<�M�<o��<I��<J6�<wѿ<�h�<Y��<��<�<i��<
%�<��<v#�<p��<��<���<���<1c�<�̪<�2�<镧<��<vS�<	��<��<;[�<�<k��<iL�<K��<�<�)�<�o�<���<���<�6�<�u�<���<V��<�+�<f�<j��<�ׁ<��<��|<��x<gu<��q<>n<+�j<Ug<�c<i�_<�W\<�X<�3U<=�Q<�N<r�J<c�F<msC<��?<�h<<��8<�i5<��1<'w.<8+<�'<:'$<O� <\<G�<��<�N<�<��<!p	<F1<%�<ϊ�;b1�;��;���;�s�;�O�;59�;71�;V7�;xL�;0p�;�;��;6�;Ė�;��;���;$�;Y��;id�;#�;��;�π;�{w;lvm;p�c;��Y;� P;�F;W*=;5�3;ɪ*;Y�!;��;��;%;��:X��:���:��:U��:BQ�:7�:HI�:�s:��S:r5:3�:���9�1�9�t9��8�07Y�ϸ��Y��J��;ݹ�[
�^�%�*A��?\�g#w�눺W,��X���l��so��|\ʺ�7׺��-��hd�����2E�^�����r���$�HG*��j0��6��<�ʾB�@�H�	�N���T�G[��a��g�m�%s��+y��1�ӛ��
���Z���V�������ꯑ�"���!����Ś��  �  �f=�=��=#B=�=�}==� =�T =l��<w�<�Q�<��<���<��<�%�<7X�<���<��<:��<7�<�C�<<o�<+��<���<���<�<�1�<�S�<[t�<֒�<|��<8��<���<���<��<E �<B0�<�=�<I�<�Q�<X�<�[�<`\�<eZ�<�U�<�M�<AC�<�5�<�$�<��<n��<���<���<���<�z�<�R�<�&�<.��<��<-��<�R�<9�<��<��<FB�<���<��<�M�<p��<S��<\6�<wѿ<�h�<V��<��<�<d��<%�<��<�#�<n��<��<���<���<<c�<�̪<�2�<ߕ�<��<hS�<��<��<3[�<�<Y��<tL�<M��<�<�)�<�o�<���<���<�6�<�u�<³�<X��<�+�<	f�<g��<�ׁ<��<��|<��x<gu<��q<>n<0�j<@g<�c<a�_<�W\< �X<�3U<`�Q<mN<��J<a�F<qsC<��?<�h<<��8<�i5<��1<w.<@+<�'<''$<f� <\<`�<q�<�N<�<��<p	<$1<B�<���;~1�;��;���;�s�;xO�;�9�;11�;x7�;�L�;!p�;뢼;��;6�;���;�;���;`�;���;Yd�;A#�;��;�π;q{w;�vm;k�c;e�Y;� P;��F;�*=;��3;��*;��!;�;�;�;^��:���:���:&�:��:�Q�:36�:�I�:�s:��S:�5:o�:|��9�1�9�%t9_�8��07�ϸһY�K���:ݹgZ
���%��'A��?\��"w�jꈺT,���W���m���n��R]ʺ8׺:亦��{d��$���D�K��U������$�G*�Jk0�׊6���<���B�5�H��N�q�T�_[�a�g��m��$s��+y�G1�⛂� �������N���Ϫ��ȯ��������GŚ��  �  �f=�=�='B=�=�}==� =�T =o��<x�<�Q�<��<���<��<�%�<5X�<���<��<B��<C�<�C�<Ko�< ��<���<���<
�<�1�<�S�<Jt�<ʒ�<���<*��<���<���<��<T �<90�<�=�<I�<�Q�<�W�<�[�<^\�<YZ�<�U�<�M�<FC�<�5�<�$�<��<l��<���<���<���<�z�<�R�<�&�</��<��<*��<�R�<;�<��<%��<<B�<���<��<�M�<l��<E��<K6�<oѿ<�h�<L��<"��<�<l��<%�<��<�#�<c��<��<���<���<4c�<}̪<�2�<ӕ�<)��<fS�<��<��<1[�<��<Y��<pL�<C��<	�<�)�<�o�<���<���<�6�<�u�<γ�<S��<�+�<f�<Z��<�ׁ<��<��|<��x<gu<��q<	>n<P�j<<g<�c<\�_<�W\<-�X<�3U<@�Q<qN<��J<J�F<�sC<��?<�h<<��8<ri5<��1<w.<C+<4�'<'$<Y� <�[<W�<n�<�N<�<ô<5p	<1<a�<���;{1�;���;���;�s�;gO�;=9�;1�;�7�;FL�;6p�;��;��;M6�;���;��;���;*�;O��;Rd�;:#�;o�;Ѐ;.{w;�vm;��c;P�Y;W!P;��F;�*=;��3;��*;a�!;��;��;�;Z��:p��:n��:<�:f��:WR�:�5�:�J�:rs:�S:5:��:G��9�/�9�$t9��8�17��ϸ��Y�hI��Y>ݹ�Y
���%��)A�A\��"w��ꈺ�,��AW��Zn���m��]ʺ�7׺��ú�/c��!���D����������_$��F*�Ck0�K�6��<�<�B�X�H�^�N��T��[�a�g�m�6%s��+y��1����������������ת���������I����Ś��  �  �f=�=��=$B=�=�}==� =�T =k��<g�<�Q�<��<���< ��<�%�<?X�<���<��<8��<:�<�C�<5o�<$��<���<���<�<�1�<�S�<Mt�<ݒ�<���<3��<���<��<��<A �<D0�<�=�<"I�<�Q�<�W�<�[�<Y\�<eZ�<�U�<�M�<3C�<~5�<�$�<��<j��<���<���<���<�z�<�R�<�&�<3��<��<'��<�R�<;�<��<��<FB�<���<��<�M�<s��<P��<Q6�<�ѿ<�h�<W��<��<�<^��<
%�<��<�#�<w��<��< ��<���<8c�<�̪<�2�<ڕ�<��<kS�<��<��<([�<���<a��<qL�<V��<�<�)�<�o�<���<���<�6�<�u�<���<K��<�+�<f�<e��<�ׁ<��<��|<��x<&gu<��q<>n<"�j<@g<�c<i�_<�W\<6�X<�3U<F�Q<�N<v�J<^�F<vsC<��?<�h<<��8<�i5<��1<w.< +< �'<-'$<`� <\<V�<��<�N<��<��<"p	<+1<3�<���;�1�;���;���;�s�;�O�;I9�;M1�;�7�;iL�;/p�;Ѣ�;��;�5�;�;��;ц�;F�;q��;|d�;&#�;��;�π;w{w;2vm;Z�c;��Y;� P;��F;C*=;	�3;٪*;��!;��;�;�;��:8��:i��:A�:���:	Q�:/6�:8J�:�s:��S:�5:�:���9k4�9M#t9)�8�07��ϸw�Y��J���;ݹ0Z
���%�S)A�?\��"w��ꈺ�,��AW���m��3o��#]ʺ�7׺p�W��8d������D���V������$��G*�ak0��6���<���B���H�"�N�L�T�k[�pa��g��m��$s�]+y��1�ԛ���������d�������󯑻�����{Ś��  �  �f=�= �=B=�=�}==)� =�T =}��<��<�Q�<��<r��<��<�%�<=X�<���<$��<A��</�<�C�<3o�<3��<���<���<�<�1�<�S�<Bt�<ْ�<p��<9��<���<���<�<9 �<N0�<�=�<I�<�Q�<�W�<�[�<S\�<pZ�<�U�<�M�<@C�<�5�<�$�<��<���<���<��<���<�z�<�R�<�&�<9��<��<E��<�R�<B�<��<��<WB�<���<��<�M�<j��<J��<F6�<yѿ<�h�<_��<��<(�<h��<	%�<��<q#�<s��<��<���<���<<c�<�̪<�2�<땧<��<}S�<��<��<F[�<���<b��<aL�<N��<��<�)�<�o�<���<��<�6�<�u�<ó�<X��<�+�<�e�<v��<�ׁ<��<��|<��x<gu<��q<1>n<�j<zg<�c<s�_<�W\<�X<�3U<4�Q<�N<c�J<~�F<YsC<��?<�h<<��8<�i5<��1<1w.<T+<,�'<$'$<8� <\<1�<~�<�N<"�<��<p	<R1<0�<֊�;s1�;���;ڥ�;�s�;�O�;!9�;>1�;I7�;�L�;3p�;�;.�;�5�;薫;��;���;�;W��;[d�;#�;��;�π;�{w;�vm;Ðc;��Y; P;e�F;�*=;?�3;��*;R�!;��;��;;���:��:6��:��::�Q�:@7�:"I�:|s:z�S:�5:b�:���9v2�9+t9��8�h07ǫϸp�Y��J��{9ݹg\
���%��*A��?\�X$w�kꈺ�,���W���l�� o��\ʺ68׺�{���c�����xE�G�������T$��F*��j0�R�6��<���B�3�H���N���T�� [��a��g�;m�%s��+y��1�����5������u���������=�������Ś��  �  �f=�=��=$B=�=�}==� =�T =k��<g�<�Q�<��<���< ��<�%�<?X�<���<��<8��<:�<�C�<5o�<$��<���<���<�<�1�<�S�<Mt�<ݒ�<���<3��<���<��<��<A �<D0�<�=�<"I�<�Q�<�W�<�[�<Y\�<eZ�<�U�<�M�<3C�<~5�<�$�<��<j��<���<���<���<�z�<�R�<�&�<3��<��<'��<�R�<;�<��<��<FB�<���<��<�M�<s��<P��<Q6�<�ѿ<�h�<W��<��<�<^��<
%�<��<�#�<w��<��< ��<���<8c�<�̪<�2�<ڕ�<��<kS�<��<��<([�<���<a��<qL�<V��<�<�)�<�o�<���<���<�6�<�u�<���<K��<�+�<f�<e��<�ׁ<��<��|<��x<&gu<��q<>n<"�j<@g<�c<i�_<�W\<6�X<�3U<F�Q<�N<v�J<^�F<vsC<��?<�h<<��8<�i5<��1<w.< +< �'<-'$<`� <\<V�<��<�N<��<��<"p	<+1<3�<���;�1�;���;���;�s�;�O�;I9�;M1�;�7�;iL�;/p�;Ѣ�;��;�5�;�;��;ц�;F�;q��;|d�;&#�;��;�π;w{w;2vm;Z�c;��Y;� P;��F;C*=;	�3;٪*;��!;��;�;�;��:8��:i��:A�:���:	Q�:/6�:8J�:�s:��S:�5:�:���9k4�9M#t9)�8�07��ϸw�Y��J���;ݹ0Z
���%�S)A�?\��"w��ꈺ�,��AW���m��3o��#]ʺ�7׺p�W��8d������D���V������$��G*�ak0��6���<���B���H�"�N�L�T�k[�pa��g��m��$s�]+y��1�ԛ���������d�������󯑻�����{Ś��  �  �f=�=�='B=�=�}==� =�T =o��<x�<�Q�<��<���<��<�%�<5X�<���<��<B��<C�<�C�<Ko�< ��<���<���<
�<�1�<�S�<Jt�<ʒ�<���<*��<���<���<��<T �<90�<�=�<I�<�Q�<�W�<�[�<^\�<YZ�<�U�<�M�<FC�<�5�<�$�<��<l��<���<���<���<�z�<�R�<�&�</��<��<*��<�R�<;�<��<%��<<B�<���<��<�M�<l��<E��<K6�<oѿ<�h�<L��<"��<�<l��<%�<��<�#�<c��<��<���<���<4c�<}̪<�2�<ӕ�<)��<fS�<��<��<1[�<��<Y��<pL�<C��<	�<�)�<�o�<���<���<�6�<�u�<γ�<S��<�+�<f�<Z��<�ׁ<��<��|<��x<gu<��q<	>n<P�j<<g<�c<\�_<�W\<-�X<�3U<@�Q<qN<��J<J�F<�sC<��?<�h<<��8<ri5<��1<w.<C+<4�'<'$<Y� <�[<W�<n�<�N<�<ô<5p	<1<a�<���;{1�;���;���;�s�;gO�;=9�;1�;�7�;FL�;6p�;��;��;M6�;���;��;���;*�;O��;Rd�;:#�;o�;Ѐ;.{w;�vm;��c;P�Y;W!P;��F;�*=;��3;��*;a�!;��;��;�;Z��:p��:n��:<�:f��:WR�:�5�:�J�:rs:�S:5:��:G��9�/�9�$t9��8�17��ϸ��Y�hI��Y>ݹ�Y
���%��)A�A\��"w��ꈺ�,��AW��Zn���m��]ʺ�7׺��ú�/c��!���D����������_$��F*�Ck0�K�6��<�<�B�X�H�^�N��T��[�a�g�m�6%s��+y��1����������������ת���������I����Ś��  �  �f=�=��=#B=�=�}==� =�T =l��<w�<�Q�<��<���<��<�%�<7X�<���<��<:��<7�<�C�<<o�<+��<���<���<�<�1�<�S�<[t�<֒�<|��<8��<���<���<��<E �<B0�<�=�<I�<�Q�<X�<�[�<`\�<eZ�<�U�<�M�<AC�<�5�<�$�<��<n��<���<���<���<�z�<�R�<�&�<.��<��<-��<�R�<9�<��<��<FB�<���<��<�M�<p��<S��<\6�<wѿ<�h�<V��<��<�<d��<%�<��<�#�<n��<��<���<���<<c�<�̪<�2�<ߕ�<��<hS�<��<��<3[�<�<Y��<tL�<M��<�<�)�<�o�<���<���<�6�<�u�<³�<X��<�+�<	f�<g��<�ׁ<��<��|<��x<gu<��q<>n<0�j<@g<�c<a�_<�W\< �X<�3U<`�Q<mN<��J<a�F<qsC<��?<�h<<��8<�i5<��1<w.<@+<�'<''$<f� <\<`�<q�<�N<�<��<p	<$1<B�<���;~1�;��;���;�s�;xO�;�9�;11�;x7�;�L�;!p�;뢼;��;6�;���;�;���;`�;���;Yd�;A#�;��;�π;q{w;�vm;k�c;e�Y;� P;��F;�*=;��3;��*;��!;�;�;�;^��:���:���:&�:��:�Q�:36�:�I�:�s:��S:�5:o�:|��9�1�9�%t9_�8��07�ϸһY�K���:ݹgZ
���%��'A��?\��"w�jꈺT,���W���m���n��R]ʺ8׺:亦��{d��$���D�K��U������$�G*�Jk0�׊6���<���B�5�H��N�q�T�_[�a�g��m��$s��+y�G1�⛂� �������N���Ϫ��ȯ��������GŚ��  �  �f=�=��="B=�=�}==&� =�T =x��<s�<�Q�<��<~��<��<�%�<FX�<���<��<A��<9�<�C�<.o�<1��<���<���<�<�1�<�S�<Ht�<ؒ�<s��<6��<���<���<�<D �<E0�<�=�<I�<�Q�<�W�<�[�<S\�<kZ�<�U�<�M�<;C�<�5�<�$�<��<{��<���<��<���<�z�<�R�<�&�<<��<��<9��<�R�<C�<��<��<TB�<���<��<�M�<o��<I��<J6�<wѿ<�h�<Y��<��<�<i��<
%�<��<v#�<p��<��<���<���<1c�<�̪<�2�<镧<��<vS�<	��<��<;[�<�<k��<iL�<K��<�<�)�<�o�<���<���<�6�<�u�<���<V��<�+�<f�<j��<�ׁ<��<��|<��x<gu<��q<>n<+�j<Ug<�c<i�_<�W\<�X<�3U<=�Q<�N<r�J<c�F<msC<��?<�h<<��8<�i5<��1<'w.<8+<�'<:'$<O� <\<G�<��<�N<�<��<!p	<F1<%�<ϊ�;b1�;��;���;�s�;�O�;59�;71�;V7�;xL�;0p�;�;��;6�;Ė�;��;���;$�;Y��;id�;#�;��;�π;�{w;lvm;p�c;��Y;� P;�F;W*=;5�3;ɪ*;Y�!;��;��;%;��:X��:���:��:U��:BQ�:7�:HI�:�s:��S:r5:3�:���9�1�9�t9��8�07Y�ϸ��Y��J��;ݹ�[
�^�%�*A��?\�g#w�눺W,��X���l��so��|\ʺ�7׺��-��hd�����2E�^�����r���$�HG*��j0��6��<�ʾB�@�H�	�N���T�G[��a��g�m�%s��+y��1�ӛ��
���Z���V�������ꯑ�"���!����Ś��  �  �f=�=��='B=	�=�}== � =�T =t��<p�<�Q�<��<|��<��<�%�<;X�<���<��<>��<2�<�C�<>o�<(��<���<���<�<�1�<�S�<Et�<֒�<���<0��<���<���<��<J �<C0�<�=�<!I�<�Q�<�W�<�[�<U\�<kZ�<�U�<�M�<@C�<�5�<�$�<��<q��<���<��<���<�z�<�R�<�&�<7��<��<-��<�R�<5�<��<��<EB�<���<��<�M�<q��<K��<N6�<|ѿ<�h�<V��<��<�<d��<%�<��<�#�<o��<��<���<���<7c�<�̪<�2�<ޕ�<��<pS�< ��<��<0[�<���<a��<fL�<T��<�<�)�<�o�<���<���<�6�<�u�<ȳ�<V��<�+�<f�<k��<�ׁ<��<��|<��x<*gu<��q<>n<:�j<<g<�c<k�_<�W\<7�X<�3U<9�Q<�N<l�J<h�F<�sC<��?<�h<<��8<�i5<��1< w.<3+<1�'<"'$<L� <\<?�<z�<�N<��<��<p	<31<F�<���;G1�;��;���;�s�;�O�;+9�;/1�;�7�;`L�;.p�;뢼;��;%6�;���;��;ˆ�;7�;e��;ld�;#�;��;�π;F{w;�vm;��c;P�Y;� P;��F;p*=;$�3;��*;��!;�;��;�;c��:���:���:��:���:�Q�:6�:|I�:�s:l�S:�5:z�:���9E3�9d#t9x�8�07R�ϸ��Y�5J��K<ݹ�Y
�x�%��)A�t?\�##w��ꈺ�+��>X���m���n���\ʺa8׺�ں��c�����HE���������V$�CG*�k0���6���<�j�B�D�H���N�3�T�@[��a��g�m�%s�O+y��1�қ��힅�����=����������뵔�#����Ś��  �  �f=�=��=$B=�=�}== � =�T =q��<p�<�Q�<��<���<��<�%�<5X�<���<��<C��<=�<�C�<<o�<&��<���<���<�<�1�<�S�<Xt�<В�<}��</��<���<���<�<H �<=0�<�=�<I�<�Q�<X�<�[�<\\�<aZ�<�U�<�M�<@C�<�5�<�$�<��<i��<���<���<���<�z�<�R�<�&�<-��<��<&��<�R�<;�<��<��<FB�<���<��<�M�<m��<O��<X6�<qѿ<�h�<Q��<��<�<j��<%�<	��<�#�<g��<��<���<���<:c�<�̪<�2�<ܕ�<��<lS�<	��<��<*[�<���<W��<qL�<N��<�<�)�<�o�<���<���<�6�<�u�<ó�<T��<�+�<f�<e��<�ׁ<��<��|<��x<gu<��q<>n<6�j<Ng<�c<c�_<�W\<"�X<�3U<Y�Q<}N<z�J<^�F<vsC<��?<�h<<��8<�i5<��1<w.<3+<$�'<'$<e� <	\<X�<n�<�N<��<ƴ<)p	<,1<C�<���;�1�;���;���;�s�;�O�;v9�;1�;{7�;]L�;*p�;���;��;6�;���;��;���;O�;}��;Qd�;3#�;��;�π;h{w;�vm;��c;m�Y;L!P;�F;�*=;��3;�*;��!;̞;	�;�;���:$��:���:B�:Z��:�Q�:-6�:#J�:ms:�S:%5:�:x��9e0�9�"t9/	�8@�07v�ϸ̸Y�HJ���<ݹ�Z
���%��'A��?\�5#w��ꈺ�,��OW���m���n��]ʺ�7׺��<���c��.���D�F��R������$�1G*�Jk0�t�6��<���B�P�H�+�N�A�T�q[�Ka��g��m�%s��+y��1�䛂�����i���<���ʪ���������+���UŚ��  �  �f=�=��=B=�=�}==$� =�T =t��<z�<�Q�<��<���<��<�%�<:X�<���<��<C��<3�<�C�<4o�<.��<���<���<�<�1�<�S�<Gt�<ؒ�<z��<7��<���<���<
�<> �<H0�<�=�<I�<�Q�<�W�<�[�<^\�<cZ�<�U�<�M�<<C�<�5�<�$�<��<r��<���<���<���<�z�<�R�<�&�<1��<��<1��<�R�<8�<��<��<PB�<���<��<�M�<p��<H��<L6�<wѿ<�h�<\��<��< �<i��<%�<��<}#�<o��<��<���<���<:c�<|̪<�2�<啧<��<sS�<��<��<6[�<���<]��<sL�<G��<�<�)�<�o�<���<���<�6�<�u�<���<V��<�+�< f�<g��<�ׁ<��<��|<��x<gu<��q<>n<�j<cg<�c<g�_<�W\<%�X<�3U<<�Q<}N<��J<c�F<[sC<��?<�h<<��8<�i5<��1<w.<F+<�'<%'$<b� <�[<[�<y�<�N<�<Ŵ<p	<;1<1�<���;�1�;���;���;�s�;O�;29�;:1�;p7�;|L�;,p�;颼;��;�5�;Ζ�;��;���;&�;[��;dd�;;#�;��;�π;�{w;{vm;��c;{�Y;� P;͖F;�*=;��3;�*;f�!;��;�;�;���:ڦ�:���:�:���:pQ�:�6�:nI�:ys:Q�S:�5:�:M��92�9$!t9i�8iu07�ϸ:�Y�K���:ݹ�Z
�v�%��)A�M@\��"w��ꈺ�,���W��Am��!o���\ʺ>8׺��v���c������D����s������$��F*�#k0��6�G�<���B�D�H���N���T�^[�6a��g�m�!%s��+y��1�ӛ��*���>���t���ê��ᯑ����$����Ś��  �  �f=�=��=%B=�=�}=="� =�T =u��<k�<�Q�<��<���<��<�%�<;X�<���<��<@��<2�<�C�<4o�<-��<���<���<�<�1�<�S�<Ct�<ޒ�<x��<3��<���<���<�<A �<Q0�<�=�<&I�<�Q�<X�<�[�<P\�<oZ�<�U�<�M�<6C�<�5�<�$�<��<r��<���< ��<���<�z�<�R�<�&�<5��<���<-��<�R�<7�<��<��<NB�<���<#��<�M�<o��<V��<L6�<�ѿ<�h�<b��<��<�<a��<%�<��<z#�<x��<��<��<���<6c�<�̪<�2�<啧<��<rS�<���<��<-[�<���<_��<lL�<Q��<�<�)�<�o�<���<���<�6�<�u�<���<R��<�+�<	f�<m��<�ׁ<��<��|<��x<(gu<��q<5>n<#�j<Mg<�c<��_<�W\<.�X<�3U<>�Q<�N<c�J<j�F<xsC<��?<�h<<��8<�i5<��1<!w.<)+<-�'<$'$<Y� <\<L�<y�<�N<��<��<p	<71<2�<���;^1�;��;���;�s�;�O�;"9�;Q1�;i7�;kL�;Cp�;֢�;��;�5�;�;��;↠;)�;���;rd�;#�;��;�π;�{w;Jvm;~�c;l�Y;� P;ǖF;>*=;�3;̪*;��!;؞;��;�;��:���:���:��:h��:'Q�:�6�:AI�:3s:��S:_5:Ѣ:[��95�9�t9��8F�07��ϸ'�Y�WJ���:ݹH[
�k�%�9*A�>\��#w��ꈺ�+��X��<m��8o���\ʺl8׺���;d�����E�.��s�����c$�nG*�k0��6�e�<���B�c�H�)�N�q�T�+[��a�yg��m�
%s�T+y��1��������j���g������������������Ś��  �  �f=�=��=%B=�=�}==� =�T =v��<o�<�Q�<��<���<��<�%�<7X�<���<��<I��<?�<�C�<Co�<*��<���<���<�<�1�<�S�<Kt�<ђ�<}��<-��<���<���<�<K �<>0�<�=�<I�<�Q�<�W�<|[�<\\�<dZ�<�U�<�M�<CC�<�5�<�$�<��<p��<���<��<���<�z�<�R�<�&�<2��<��<,��<�R�<>�<��< ��<JB�<���<��<�M�<g��<M��<I6�<yѿ<�h�<R��<��<�<k��<%�<	��<#�<k��<��<���<���<<c�<�̪<�2�<���< ��<lS�<��<��<-[�<��<\��<nL�<G��<�<�)�<�o�<���<���<�6�<�u�<ʳ�<W��<�+�<f�<h��<�ׁ<��<��|<��x<'gu<��q<>n<>�j<Ig<�c<j�_<�W\<2�X<�3U<F�Q<vN<z�J<`�F<xsC<��?<�h<<��8<�i5<��1<#w.<1+<;�'<'$<[� <�[<R�<r�<�N<��<Ѵ<,p	<&1<P�<���;l1�;��;ĥ�;�s�;�O�;A9�;1�;~7�;TL�;8p�;���;��;&6�;���;��;���;�;m��;Bd�;3#�;��;�π;�{w;�vm;��c;v�Y;b!P;��F;�*=;�3;��*;_�!;��;��;�;��:���:���:u�:���:�Q�:g6�:�I�:�s:#�S:v5:��:���9a2�93 t9�
�8��07��ϸ��Y��I���<ݹ�Z
��%��)A��?\��#w�iꈺv,���W���m��]n��]ʺ�7׺:�	��Tc����
E����u�����B$�8G*�k0�V�6���<�V�B�:�H�'�N�J�T�U[�Oa�	g��m�E%s�\+y��1�ڛ��䞅�s���5��������������H���zŚ��  �  �f=�=��=#B=�=�}==� =�T =i��<v�<�Q�<��<���<��<�%�</X�<���<��<=��<1�<�C�<Ao�<��<���<���<�<�1�<�S�<\t�<Ғ�<���<5��<���<���<��<G �<?0�<�=�<I�<�Q�<X�<|[�<i\�<XZ�<�U�<�M�<;C�<�5�<�$�<��<f��<���<���<���<�z�<�R�<�&�<'��<��<#��<�R�<1�<��<��<>B�<���<��<�M�<l��<Q��<V6�<wѿ<�h�<S��<��<�<c��<%�<��<�#�<j��<��<�<���<>c�<|̪<�2�<ӕ�<��<kS�<���<��<+[�<���<S��<~L�<E��<�<�)�<�o�<���<���<�6�<�u�<ͳ�<N��<�+�<f�<_��<�ׁ<��<��|<��x<#gu<��q<>n<4�j<8g<�c<_�_<�W\<4�X<�3U<h�Q<\N<��J<S�F<psC<��?<�h<<��8<�i5<��1<	w.<@+<�'<'$<w� <�[<q�<c�<�N<��<��<p	<(1<K�<{��;�1�;���;���;�s�;[O�;�9�;1�;�7�;rL�; p�;㢼;��;6�;���;�;���;F�;���;Bd�;h#�;i�;�π;5{w;rvm;��c;"�Y;� P;h�F;�*=;��3;��*;��!;��;D�;;��:���:���:��:Z��:�Q�:�5�:�J�:/s:q�S:5:*�:���9�1�9�(t9��8ڪ07o�ϸ�Y�;K���;ݹOY
�"�%�{'A��@\�z"w�Tꈺ�,���V��Zn��~n��$]ʺ�8׺��1���c��O���D���� ������$��F*�}k0��6�Ȧ<�B�B���H�'�N�^�T��[��a�]g�sm�%s�k+y�Z1�雂���������P���Ҫ��ׯ��񵔻6���7Ś��  �  �f=�=��=%B=�=�}==%� =�T =z��<z�<�Q�<��<~��<��<�%�<:X�<���<��<I��<6�<�C�<8o�<(��<���<���<�<�1�<�S�<It�<Β�<r��<0��<���<���<�<H �<G0�<�=�<I�<�Q�< X�<[�<S\�<`Z�<�U�<�M�<>C�<�5�<�$�<��<x��<���<���<���<�z�<�R�<�&�<3��<��<6��<�R�<=�<��<��<HB�<���<��<�M�<h��<N��<F6�<rѿ<�h�<X��<��<"�<m��<%�<��<w#�<h��<��<���<���<-c�<�̪<�2�<ߕ�<��<wS�<��<��<7[�<���<^��<hL�<F��<�<�)�<�o�<���<���<�6�<�u�<ĳ�<U��<�+�<f�<a��<�ׁ<��<��|<��x<gu<��q<'>n<4�j<dg<�c<r�_<�W\<�X<3U<J�Q<zN<p�J<S�F<zsC<��?<�h<<��8<�i5<��1<,w.<F+<&�'<$'$<Q� <�[<D�<x�<�N<�<Ѵ<p	<C1<9�<���;1�;��;���;�s�;�O�;99�;1�;R7�;^L�;9p�; ��; �;6�;˖�;��;���;�;t��;Nd�;#�;��;�π;o{w;�vm;��c;��Y;� P;��F;�*=;�3;Ī*;C�!;��;��;�;���:$��:���:g�:���:�Q�:H6�:DJ�:gs:��S:�5:ء:��9�0�9�t9#�8��07��ϸ^�Y�^J���;ݹ�[
�[�%��)A�u?\��#w�b눺n,��mW���m���n��k\ʺ8׺n�n���c�����9E�����������$��F*��j0�Ɋ6�5�<���B�O�H�*�N�D�T��[��a��g��m�T%s��+y��1���������<���F����������5���J���sŚ��  �  Pg=�=s�=�B=��=c~=�=� =�U =U��<k�<�S�<N��<���<���<d(�<+[�<���<W��<���<��<�G�<(s�<\��<���<+��<��<�6�<Y�<�y�<r��<=��<0��<��<���<��<'�<d7�<,E�<�P�<�Y�<�_�<�c�<�d�<c�<t^�<W�<�L�<?�<}.�<��<��<.��<���<S��<Յ�<�]�<�1�<��<m��<ǘ�<7^�< �<���<���<@N�<� �<��<�Y�<o �<?��<3B�<cݿ<�t�<�<���<�#�<���<;0�<��<P.�<&��<R�<7��<� �<m�<֪<�;�<잧<���<�[�</��<��<�b�<+��<S�< S�<���<�<a/�<�t�<���<���<�:�<�y�<U��<��<�.�<�h�<���<�ف<3�<܏|<i�x<hu<��q<�=n<�j<vg<�|c<1�_<�S\<��X<8.U<!�Q<�N< �J<H�F<�jC<O�?<�^<<��8<^5<I�1<1j.<��*<Մ'<&$<�� <L<b�<�<i<<O�<��<A\	<�<6�<�_�;Z�;��;�w�;E�; �;��;P �;��;	�;A=�;\o�;���;��;.b�;�ѥ;�Q�;���;��;�.�;��;c��;q��;�w;1m;�'c;�aY;��O;1F;�<;^x3;�G*;�5!;�?;Cd;q�;��:|��:�:m�:��:��:"��:E��:��q:��R:��3:Ԇ:Q��9m �9~p9�@�8�?�6q׸L]����s�޹�)���&�d�A���\���w��?���~��n���ڸ��F���<�ʺ�z׺�A�r�����y��_�7����i��3$�r[*��}0���6�z�<��B�7�H�R�N�� U��[�0a�yg��%m��+s��0y��6���������0���٦��z���l���ٴ��q���yÚ��  �  Mg=�=n�=�B=��=^~=�=� =�U =T��<s�<�S�<_��<��<���<f(�<4[�<ь�<]��<���<��<�G�<1s�<S��<��<2��<��<�6�<Y�<�y�<c��<=��<,��<��<���<��<$'�<\7�<+E�<�P�<�Y�<`�<�c�<�d�<c�<�^�<W�<�L�<?�<u.�<��<��<:��<���<d��<���<�]�<�1�<��<x��<Ř�<>^�<��<���<��<<N�<� �<��<�Y�<g �<J��<>B�<Tݿ<�t�<	�<���<�#�<���<=0�<��<S.�<��<a�<<��<� �<�l�<֪< <�<䞧<���<�[�<,��<��<�b�<;��<X�<S�<���<��<t/�<�t�<���<���<�:�<�y�<W��<��<�.�<�h�<���<�ف<-�<��|<e�x<	hu<��q<�=n<�j<wg<	}c<(�_<�S\<x�X<,.U<A�Q<�N<�J<4�F<�jC<_�?<�^<<��8< ^5<W�1<0j.<��*<�'<H$<�� <�K<f�<�<�<<\�<{�<?\	<�<H�<�_�;��;'��;�w�;E�; �;	�; �;��;��;==�;so�;���;��;b�;�ѥ;�Q�;���;��;�.�;��;:��;���;�w;Im;�'c;�aY;��O;�0F;m�<;�x3;UH*; 5!;�>;�d;��;/�:X��:u�:�l�:+��:���:하:,��:��q:��R:��3:G�:��9��9Kp9�6�8���6�׸�I]�a����޹�)���&���A�7�\�}�w�[@���~������`���������ʺ�z׺�A�=�����Q��_���������W3$�3[*��}0�u�6�ж<���B�n�H��N�9 U�P[�Ea��g�k%m��+s�81y��6�����]���/�����������n���鴔�����:Ú��  �  Ig=�=l�=�B=��=[~=�=� =�U =L��<s�<�S�<U��< ��<���<{(�<![�<ˌ�<U��<���<��<�G�<;s�<L��<��<,��<��<�6�<Y�<�y�<Y��<L��<0��<��<���<��<%'�<W7�<?E�<�P�<�Y�<�_�<�c�<�d�<c�<�^�<W�<�L�<?�<t.�<��<��<>��<~��<h��<ȅ�<�]�<�1�<z�<z��<���<D^�<��<���<��<2N�<� �<��<�Y�<f �<@��<;B�<Sݿ<�t�<�<���<�#�<���<<0�<��<e.�<��<`�<3��<� �<	m�<
֪<<�<ڞ�<���<�[�<2��<��<�b�<9��<B�<S�<���<
�<n/�<�t�<���<���<�:�<�y�<b��<��<�.�<�h�<���<�ف<'�<�|<U�x<hu<�q<�=n<��j<Tg<}c<�_<�S\<��X<.U<<�Q<�N<�J<.�F<�jC<[�?<�^<<��8<�]5<f�1< j.<��*<ӄ'<2$<ӯ <�K<��<�<�<<K�<u�<M\	<�<]�<�_�;��;��;�w�;1E�;��;	�;���;��;�;0=�;^o�;���;��;�a�;ҥ;�Q�;���;��;�.�;��;.��;̚�;Ww;Bm;�'c;�aY;�O;�0F;��<;�w3;vH*;�5!;?; e;إ;\�:���:��:�l�:H��:���:L��:���:r�q:u�R:��3:��:H��9��9�p9�2�8���6�!׸9N]������޹8'�~�&���A�P�\���w��?���~��Z����������ޢʺ�z׺�A����!������^�G�������3$�)[*�~0�/�6��<���B���H�2�N�" U��[��a��g��%m�,s�1y�86�����b���t�����������I���Ĵ������BÚ��  �  Pg=�=k�=�B=��=`~=�=� =�U =N��<y�<�S�<L��<���<���<j(�<"[�<֌�<Y��<���<��<�G�</s�<V��<��<'��<��<�6�<Y�<�y�<`��<A��<,��<��<���<��<"'�<Z7�<3E�<�P�<�Y�<�_�<�c�<�d�<c�<�^�<W�<�L�<?�<q.�<��<��<F��<���<Z��<ą�<�]�<�1�<��<���<���<<^�<��<���<���<=N�<� �<��<�Y�<m �<D��<5B�<Tݿ<�t�<�<���<�#�<���<=0�<��<W.�<��<Y�<;��<� �<�l�<֪<<�<垧<���<�[�<0��<��<�b�<D��<H�<S�<���<�<b/�<�t�<���<���<�:�<�y�<[��<��<�.�<�h�<���<�ف<4�<�|<X�x<
hu<�q<�=n<��j<sg<}c<$�_<�S\<{�X<$.U<3�Q<�N<�J<+�F<�jC<^�?<�^<<��8<�]5<X�1<$j.<��*<�'<"$<�� <�K<n�<�<�<<S�<z�<H\	<�<E�<�_�;��;���;�w�;E�; �;��;	 �;��;��;:=�;uo�;���;��;b�;�ѥ;�Q�;���;��;�.�;��;-��;���;�w;2m;�'c;{aY;ǹO;�0F;��<;Ix3;H*;\5!;?;�d;0�;�:���:d�:|l�:*��:R��:���:��:��q:��R:j�3:x�:���9��9lp9S4�8T��6�׸�I]����Q�޹�(���&�y�A�H�\���w��@��4������E���������ʺ�z׺�A云��r�����|_�<��3��d��3$��Z*��}0�w�6���<���B�Y�H��N�f U�z[�2a�ug��%m� ,s�61y�h6�����e���6�����������c���ⴔ�����VÚ��  �  Rg=�=r�=�B=��=]~=�=� =�U =T��<m�<�S�<Z��<���<���<j(�</[�<̌�<V��<���<��<�G�<+s�<R��<���<7��<��<�6�<Y�<�y�<m��<?��<3��<��<���<��<'�<a7�<-E�<�P�<�Y�<�_�<�c�<�d�<c�<�^�<
W�<�L�<?�<x.�<��<��<5��<���<e��<ą�<�]�<�1�<��<s��<�<>^�<��<���<���<=N�<� �<"��<�Y�<n �<F��<7B�<]ݿ<�t�<�<���<�#�<���<60�<��<U.�<!��<U�<@��<� �<�l�<֪<�;�<㞧<���<�[�<,��<��<�b�<6��<U�<S�<���<�<q/�<�t�<���<���<�:�<�y�<Y��<��<�.�<�h�<���<�ف<5�<�|<p�x<hu<��q<�=n<�j<}g<�|c<(�_<�S\<}�X<:.U<'�Q<�N<�J<E�F<�jC<T�?<�^<<��8<^5<S�1<1j.<��*<�'<>$<�� <�K<n�<
�<�<<N�<~�<<\	<�<<�<�_�;z�;<��;�w�;�D�;" �;��;> �;��;�;*=�;Ko�;���;��;"b�;�ѥ;�Q�;���;��;�.�;��;o��;���;�w;�m;�'c;�aY;��O;�0F;A�<;rx3;]H*;`5!;?;�d;i�;��:,��:{�:�l�:���:ެ�:��:���:��q:��R:��3:͇:w��9(�9p9�<�82
�6�׸�M]�2����޹;)�S�&��A���\���w�x@��~��񦣺d���,���١ʺ�z׺�A云��P���j�y_�L��2�����3$�`[*��}0�|�6���<���B�}�H�;�N�W U��[��a�jg��%m��+s�1y��6���������"���ڦ������[���ߴ��n���nÚ��  �  Ng=�=p�=�B=��=^~=�=� =�U =R��<w�<�S�<Q��<���<���<u(�<$[�<̌�<Y��<���<��<�G�<6s�<S��< ��<0��<��<�6�<Y�<�y�<c��<<��<-��<��<���<��<%'�<Y7�<3E�<�P�<�Y�<�_�<�c�<�d�<c�<�^�<
W�<�L�<?�<r.�<��<��<B��<���<b��<Ņ�<�]�<�1�<�<��<���<@^�<��<���<���<=N�<� �<��<�Y�<n �<@��<:B�<Vݿ<�t�<	�<���<�#�<���<:0�<��<V.�<��<]�<:��<� �<m�<֪<�;�<䞧<���<�[�<*��<��<�b�<:��<I�<S�<���<�<j/�<�t�<���<���<�:�<�y�<a��<��<�.�<�h�<���<�ف</�<�|<e�x<hu< �q<�=n<�j<tg<	}c<�_<�S\<p�X<).U<3�Q<�N<�J<>�F<�jC<W�?<�^<<��8<^5<R�1<,j.<��*<ڄ'<+$<ͯ <�K<��<��<�<<T�<|�<<\	<�<R�<�_�;~�;��;�w�;E�; �;��; �;��;��;0=�;po�;���;��;b�;�ѥ;�Q�;���;��;�.�;��;O��;���;�w;m;�'c;�aY;׹O;�0F;��<;x3;JH*;k5!;?;�d; �;��:��:��:ul�:���:6��:���:��:Z�q:�R:�3:
�:��9/�9�p96�8���6�׸�J]�C����޹%)���&���A�k�\���w�@���~��Ȧ��^�������<�ʺ{׺�A争�������*_�P����!��3$�[*��}0�}�6�ܶ<���B�u�H�7�N�o U� [�'a��g��%m��+s�K1y�{6�����[���4�����������^�����������VÚ��  �  Jg=�=k�=�B=��=[~=�=� =�U =I��<x�<�S�<S��<���<���<u(�<%[�<ٌ�<V��<���<��<�G�<4s�<K��<	��<0��<��<�6�<Y�<�y�<Y��<H��<.��<��<���<��<&'�<R7�<BE�<�P�<�Y�< `�<�c�<�d�<c�<�^�<W�<�L�<?�<o.�<��<��<I��<���<d��<���<�]�<�1�<�<���<���<C^�<��<���<���<6N�<� �<��<�Y�<h �<C��<:B�<Kݿ<�t�<�<���<�#�<���<:0�<��<b.�<��<a�<4��<� �<�l�<֪<<�<ܞ�<���<�[�<2��<��<�b�<G��<G�<S�<���<�<k/�<�t�<���<���< ;�<�y�<^��<��<�.�<�h�<���<�ف<&�<��|<Z�x<hu<�q<�=n<�j<Jg<}c<�_<�S\<}�X<.U<A�Q<�N<�J<*�F<�jC<c�?<�^<<��8<�]5<l�1<j.<��*<�'</$<̯ <�K<��<��<�<<M�<v�<R\	<�<N�<�_�;��;��;�w�;E�;��;	�;���;��;�;-=�;io�;���;��;�a�;ҥ;gQ�;���;��;�.�;��;+��;Ӛ�;{w;�m;�'c;gaY;�O;[0F;��<;$x3;UH*;:5!;�>;�d; �;0�:U��:��:sl�:>��:��:���:���:|�q:f�R:��3:Z�:7��9��9Rp9�.�84��6"׸�L]����޹�'�ڥ&�u�A�&�\�-�w��@���~��+���⹰�����ޢʺ�z׺�A����6�����1_������ ��3$��Z*�&~0�'�6�$�<���B���H��N�" U�y[�'a��g�s%m��+s�>1y�6�����G���������������:���ߴ������:Ú��  �  Og=�=n�=�B=��=`~=�=� =�U =O��<p�<�S�<V��<���<���<p(�<&[�<ˌ�<V��<���<��<�G�<5s�<W��< ��</��<��<�6�<Y�<�y�<e��<D��<*��<��<���<��<''�<U7�<5E�<�P�<�Y�<�_�<�c�<�d�<c�<�^�<
W�<�L�<?�<s.�<��<��<<��<���<b��<ƅ�<�]�<�1�<��<z��<���<A^�<��<���<��<<N�<� �<��<�Y�<q �<A��<8B�<Vݿ<�t�<�<���<�#�<���<90�<��<\.�<��<Z�<9��<� �<�l�<֪<�;�<枧<���<�[�<,��<��<�b�<9��<L�<S�<���<�<l/�<�t�<���<���<�:�<�y�<`��<��<�.�<�h�<���<�ف<1�<�|<e�x<hu< �q<�=n<
�j<eg<}c<�_<�S\<}�X</.U<&�Q<�N<�J<4�F<�jC<V�?<�^<<��8<�]5<_�1<&j.<��*<݄'<5$<ǯ <�K<z�<��<�<<N�<��<C\	<�<Q�<�_�;}�;��;�w�;$E�; �;��; �;��;��;)=�;zo�;尶;��;�a�;�ѥ;�Q�;���;��;�.�;��;I��;���;�w;2m;�'c;�aY;�O;�0F;y�<;=x3;JH*;o5!;"?;�d;4�;Y�:��:��:el�:���:k��::��:d�q:��R:��3:�:���9f�9`p90�8\��6*׸J]�w����޹K(�:�&�Y�A���\�o�w�X@���~��Ŧ��>�������g�ʺ�z׺�A亢��$�����F_�������3$�=[*��}0�G�6�ٶ<���B�O�H�,�N�d U�H[�a��g��%m��+s�(1y�z6�ȝ��J���S�����������d���޴������oÚ��  �  Tg=�=n�=�B=��=a~=�=� =�U =X��<w�<�S�<Y��<��<���<f(�<0[�<ʌ�<\��<���<��<�G�<&s�<^��<��</��<��<�6�<Y�<�y�<g��<7��<3��<��<���<��<'�<a7�</E�<�P�<�Y�<�_�<�c�<�d�<c�<^�<W�<�L�<?�<y.�<��<��<9��<���<^��<���<�]�<�1�<��<t��<Ș�<=^�<  �<���<���<FN�<� �<��<�Y�<s �<C��<7B�<Wݿ<�t�<�<���<�#�<���<<0�<��<O.�<��<W�<@��<� �<�l�<֪<�;�<<���<�[�<.��<��<�b�<4��<U�<S�<���<��<m/�<�t�<���<���<�:�<�y�<T��<��<�.�<�h�<���<�ف<;�<�|<g�x<hu<�q<�=n<��j<pg<}c<(�_<�S\<j�X<3.U<'�Q<�N<�J<4�F<�jC<`�?<�^<<��8<^5<Q�1<9j.<��*<�'<<$<�� <�K<g�<�<~<<Y�<��<?\	<�<3�<�_�;��;��;�w�;E�;% �;��;' �;��;�;>=�;do�;ⰶ;��;"b�;�ѥ;�Q�;���;��;/�;��;J��;���;�w;�m;�'c;�aY;��O;�0F;a�<;{x3;%H*;A5!;?;�d;j�;��:���:r�:�l�:���:㬨:���:���:g�q:��R:�3:d�:p��9��9sp9.=�8�u�6׸�K]�����޹�)��&���A���\���w��@���~��Ѧ������g���.�ʺ�z׺�A�6��k���j��_���i���{3$�[*��}0���6���<��B�_�H���N�i U�I[�va�<g��%m��+s�X1y�g6�����p���<�����������S������}���mÚ��  �  Lg=�=p�=�B=��=[~=�=� =�U =L��<w�<�S�<Y��<���<���<m(�<+[�<Ό�<X��<���<��<�G�<3s�<K��< ��<1��<��<�6�<Y�<�y�<a��<H��<1��<��<���<��<'�<U7�<?E�<�P�<�Y�<�_�<�c�<�d�<c�<�^�<W�<�L�<?�<u.�<��<��<<��<���<e��<ǅ�<�]�<�1�<��<y��<���<=^�<��<���<���<5N�<� �<��<�Y�<h �<B��<5B�<Sݿ<�t�<�<���<�#�<���<00�<��<`.�<��<X�<8��<� �<m�<֪<�;�<ܞ�<���<�[�</��<��<�b�<:��<N�<S�<���<�<n/�<�t�<���<���<�:�<�y�<^��<��<�.�<�h�<���<�ف<+�<�|<a�x<hu<�q<�=n<��j<qg<}c<�_<�S\<�X<(.U<.�Q<�N<�J<>�F<�jC<Q�?<�^<<��8<^5<\�1<!j.<��*<؄'<;$<ɯ <�K<u�<�<�<<R�<p�<F\	<�<L�<�_�;}�;$��;�w�;E�;��;��; �;��;�;=�;eo�;찶;��;�a�;ҥ;�Q�;���;��;�.�;��;Q��;���;Yw;m;�'c;�aY;˹O;�0F;y�<;$x3;^H*;y5!;%?;�d;�;B�:���:m�:�l�:���:2��:|��:��:v�q:��R:��3:P�:��9��9�p9�4�8�)�6�׸�K]�����޹�'��&���A���\�j�w�&@���~��¦��۹������H�ʺ�z׺�A二�������\_���
����3$�[*�~0�n�6���<���B���H�e�N�7 U�'[�Sa��g��%m��+s�01y�(6�ѝ��q���;�������Ī��=���ܴ������^Ú��  �  Kg=�=k�=�B=��=]~=�=� =�U =G��<�<�S�<T��<���<���<n(�<%[�<Ռ�<]��<���<��<�G�<As�<K��<
��<.��<��<�6�<Y�<�y�<^��<?��<%��<��<���<��</'�<N7�<3E�<�P�<�Y�< `�<�c�<�d�<	c�<�^�<W�<�L�<?�<m.�<��<��<K��<���<e��<���<�]�<�1�<��<���<���<C^�<��<���<��<6N�<� �<��<�Y�<h �<E��<;B�<Pݿ<�t�<��<���<�#�<ë�<>0�<��<X.�<��<b�<9��<� �<m�<֪<<�<ܞ�<���<�[�</��<��<�b�<C��<J�<S�<���<�<k/�<�t�<���<���< ;�<�y�<g��<��<�.�<�h�<���<�ف<)�<�|<]�x<hu<��q<�=n<�j<bg<}c<�_<�S\<t�X<%.U<:�Q<�N<�J<+�F<�jC<]�?<�^<<��8<�]5<h�1<j.<��*<�'<1$<į <�K<w�<��<�<<[�<r�<L\	<�<i�<�_�;��;��;�w�;E�;��;	�; �;��;��;<=�;�o�;鰶;��;�a�;�ѥ;oQ�;���;��;�.�;��;!��;Ś�;jw;nm;�'c;YaY;�O;~0F;��<;3x3;^H*;)5!;�>;�d;�;.�:���:��:El�:5��:��:���:���:
�q:��R:��3:��:���9��97p9�*�8�.�6�׸yH]�.����޹�(�,�&�Z�A���\���w�+@����6���׹�������ʺ�z׺�A���x�����G_����1����3$��Z*�2~0�*�6��<���B�N�H�7�N�: U�r[��a��g��%m��+s�N1y��6�˝��3���Y�����������o���񴔻����GÚ��  �  Og=�=n�=�B=��=]~=�=� =�U =Q��<t�<�S�<Z��<���<���<p(�<.[�<ƌ�<X��<���<��<�G�<1s�<P��<��<2��<��<�6�<Y�<�y�<g��<<��<8��< ��<���<��<'�<d7�<3E�<�P�<�Y�<�_�<�c�<�d�<c�<�^�<W�<�L�<?�<v.�<��<��<7��<���<e��<ǅ�<�]�<�1�<��<s��<���<E^�< �<���<���<9N�<� �<��<�Y�<g �<D��<6B�<Zݿ<�t�<�<���<�#�<���<<0�<��<T.�<��<V�<<��<� �<m�<֪<<�<���<���<�[�<6��<��<�b�<1��<P�<S�<���<�<p/�<�t�<���<���< ;�<�y�<\��<��<�.�<�h�<���<�ف<0�<�|<e�x<hu<�q<�=n<�j<Qg<�|c<2�_<�S\<x�X<2.U<+�Q<�N<�J<7�F<�jC<`�?<�^<<��8<�]5<k�1<*j.<��*<ք'<=$<ǯ <�K<z�<�<v<<R�<�<V\	<�<I�<�_�;��;(��;�w�;�D�;
 �;��;% �;��;(�;J=�;4o�;���;��;/b�;�ѥ;�Q�;���;��;�.�;��;I��;���;�w;m;�'c;�aY;�O;�0F;W�<;Bx3;cH*;u5!;?;�d;4�;��:���:��:�l�:2��:<��:���:!��:O�q:4�R:��3:��:K��9\�9,p9�@�8�@�6k&׸RQ]������޹C)��&���A�4�\���w�	@���~��������������ʢʺEz׺iA亠�𺜞����C_�)�������3$�-[*��}0�'�6�۶<���B�s�H��N�C U�9[�Ga��g��%m��+s�1y�C6���������y���ަ��w���?���鴔����dÚ��  �  Sg=�=s�=�B=��=b~=�=� =�U =Y��<w�<�S�<^��<��<���<c(�<4[�<ƌ�<c��<���<��<�G�<5s�<\��<���<,��<��<�6�<#Y�<�y�<k��<4��<.��<��<���<��<'�<a7�<%E�<�P�<�Y�< `�<�c�<�d�<c�<w^�<	W�<�L�<?�<p.�<��<��<5��<���<a��<Å�<�]�<�1�<��<r��<͘�<8^�<��<���<��<?N�<� �<��<�Y�<h �<J��<2B�<[ݿ<�t�<�<���<�#�<˫�<*0�<��<J.�<!��<O�<D��<� �<m�<֪<�;�<랧<���<�[�<'��<��<�b�<2��<W�<S�<���<��<r/�<�t�<���<���<�:�<�y�<_��<��<�.�<�h�<���<�ف<8�<�|<i�x<hu<��q<�=n<�j<�g<�|c<�_<�S\<g�X<3.U<!�Q<�N<�J<K�F<�jC<I�?<�^<<��8<^5<J�1<9j.<��*<؄'<F$<�� <�K<a�<�<w<<g�<}�<6\	<�<P�<�_�;L�;��;�w�;�D�;2 �;��;4 �;��;�;�<�;o�;d��;{�;#b�;�ѥ;�Q�;���;��;�.�;��;i��;{��;�w;Qm;�'c;oaY;��O;%1F;A�<;ox3;?H*;V5!;�>;�d;~�;��:���:�:Ol�:���:���:��:A��:�q:�R:��3:?�:/��9��9�p9?�8���6K�ָmD]�.����޹�*�G�&���A�'�\���w�@���~������񸰺M���J�ʺ>{׺�A���𺇞��W��_���B�����3$�*[*�x}0���6�Զ<���B�K�H�T�N�� U��[��a�Ug��%m��+s�Q1y��6�������������Ʀ������s���
���~���yÚ��  �  Og=�=n�=�B=��=]~=�=� =�U =Q��<t�<�S�<Z��<���<���<p(�<.[�<ƌ�<X��<���<��<�G�<1s�<P��<��<2��<��<�6�<Y�<�y�<g��<<��<8��< ��<���<��<'�<d7�<3E�<�P�<�Y�<�_�<�c�<�d�<c�<�^�<W�<�L�<?�<v.�<��<��<7��<���<e��<ǅ�<�]�<�1�<��<s��<���<E^�< �<���<���<9N�<� �<��<�Y�<g �<D��<6B�<Zݿ<�t�<�<���<�#�<���<<0�<��<T.�<��<V�<<��<� �<m�<֪<<�<���<���<�[�<6��<��<�b�<1��<P�<S�<���<�<p/�<�t�<���<���< ;�<�y�<\��<��<�.�<�h�<���<�ف<0�<�|<e�x<hu<�q<�=n<�j<Qg<�|c<2�_<�S\<x�X<2.U<+�Q<�N<�J<7�F<�jC<`�?<�^<<��8<�]5<k�1<*j.<��*<ք'<=$<ǯ <�K<z�<�<v<<R�<�<V\	<�<I�<�_�;��;(��;�w�;�D�;
 �;��;% �;��;(�;J=�;4o�;���;��;/b�;�ѥ;�Q�;���;��;�.�;��;I��;���;�w;m;�'c;�aY;�O;�0F;W�<;Bx3;cH*;u5!;?;�d;4�;��:���:��:�l�:2��:<��:���:!��:O�q:4�R:��3:��:K��9\�9,p9�@�8�@�6k&׸RQ]������޹C)��&���A�4�\���w�	@���~��������������ʢʺEz׺iA亠�𺜞����C_�)�������3$�-[*��}0�'�6�۶<���B�s�H��N�C U�9[�Ga��g��%m��+s�1y�C6���������y���ަ��w���?���鴔����dÚ��  �  Kg=�=k�=�B=��=]~=�=� =�U =G��<�<�S�<T��<���<���<n(�<%[�<Ռ�<]��<���<��<�G�<As�<K��<
��<.��<��<�6�<Y�<�y�<^��<?��<%��<��<���<��</'�<N7�<3E�<�P�<�Y�< `�<�c�<�d�<	c�<�^�<W�<�L�<?�<m.�<��<��<K��<���<e��<���<�]�<�1�<��<���<���<C^�<��<���<��<6N�<� �<��<�Y�<h �<E��<;B�<Pݿ<�t�<��<���<�#�<ë�<>0�<��<X.�<��<b�<9��<� �<m�<֪<<�<ܞ�<���<�[�</��<��<�b�<C��<J�<S�<���<�<k/�<�t�<���<���< ;�<�y�<g��<��<�.�<�h�<���<�ف<)�<�|<]�x<hu<��q<�=n<�j<bg<}c<�_<�S\<t�X<%.U<:�Q<�N<�J<+�F<�jC<]�?<�^<<��8<�]5<h�1<j.<��*<�'<1$<į <�K<w�<��<�<<[�<r�<L\	<�<i�<�_�;��;��;�w�;E�;��;	�; �;��;��;<=�;�o�;鰶;��;�a�;�ѥ;oQ�;���;��;�.�;��;!��;Ś�;jw;nm;�'c;YaY;�O;~0F;��<;3x3;^H*;)5!;�>;�d;�;.�:���:��:El�:5��:��:���:���:
�q:��R:��3:��:���9��97p9�*�8�.�6�׸yH]�.����޹�(�,�&�Z�A���\���w�+@����6���׹�������ʺ�z׺�A���x�����G_����1����3$��Z*�2~0�*�6��<���B�N�H�7�N�: U�r[��a��g��%m��+s�N1y��6�˝��3���Y�����������o���񴔻����GÚ��  �  Lg=�=p�=�B=��=[~=�=� =�U =L��<w�<�S�<Y��<���<���<m(�<+[�<Ό�<X��<���<��<�G�<3s�<K��< ��<1��<��<�6�<Y�<�y�<a��<H��<1��<��<���<��<'�<U7�<?E�<�P�<�Y�<�_�<�c�<�d�<c�<�^�<W�<�L�<?�<u.�<��<��<<��<���<e��<ǅ�<�]�<�1�<��<y��<���<=^�<��<���<���<5N�<� �<��<�Y�<h �<B��<5B�<Sݿ<�t�<�<���<�#�<���<00�<��<`.�<��<X�<8��<� �<m�<֪<�;�<ܞ�<���<�[�</��<��<�b�<:��<N�<S�<���<�<n/�<�t�<���<���<�:�<�y�<^��<��<�.�<�h�<���<�ف<+�<�|<a�x<hu<�q<�=n<��j<qg<}c<�_<�S\<�X<(.U<.�Q<�N<�J<>�F<�jC<Q�?<�^<<��8<^5<\�1<!j.<��*<؄'<;$<ɯ <�K<u�<�<�<<R�<p�<F\	<�<L�<�_�;}�;$��;�w�;E�;��;��; �;��;�;=�;eo�;찶;��;�a�;ҥ;�Q�;���;��;�.�;��;Q��;���;Yw;m;�'c;�aY;˹O;�0F;y�<;$x3;^H*;y5!;%?;�d;�;B�:���:m�:�l�:���:2��:|��:��:v�q:��R:��3:P�:��9��9�p9�4�8�)�6�׸�K]�����޹�'��&���A���\�j�w�&@���~��¦��۹������H�ʺ�z׺�A二�������\_���
����3$�[*�~0�n�6���<���B���H�e�N�7 U�'[�Sa��g��%m��+s�01y�(6�ѝ��q���;�������Ī��=���ܴ������^Ú��  �  Tg=�=n�=�B=��=a~=�=� =�U =X��<w�<�S�<Y��<��<���<f(�<0[�<ʌ�<\��<���<��<�G�<&s�<^��<��</��<��<�6�<Y�<�y�<g��<7��<3��<��<���<��<'�<a7�</E�<�P�<�Y�<�_�<�c�<�d�<c�<^�<W�<�L�<?�<y.�<��<��<9��<���<^��<���<�]�<�1�<��<t��<Ș�<=^�<  �<���<���<FN�<� �<��<�Y�<s �<C��<7B�<Wݿ<�t�<�<���<�#�<���<<0�<��<O.�<��<W�<@��<� �<�l�<֪<�;�<<���<�[�<.��<��<�b�<4��<U�<S�<���<��<m/�<�t�<���<���<�:�<�y�<T��<��<�.�<�h�<���<�ف<;�<�|<g�x<hu<�q<�=n<��j<pg<}c<(�_<�S\<j�X<3.U<'�Q<�N<�J<4�F<�jC<`�?<�^<<��8<^5<Q�1<9j.<��*<�'<<$<�� <�K<g�<�<~<<Y�<��<?\	<�<3�<�_�;��;��;�w�;E�;% �;��;' �;��;�;>=�;do�;ⰶ;��;"b�;�ѥ;�Q�;���;��;/�;��;J��;���;�w;�m;�'c;�aY;��O;�0F;a�<;{x3;%H*;A5!;?;�d;j�;��:���:r�:�l�:���:㬨:���:���:g�q:��R:�3:d�:p��9��9sp9.=�8�u�6׸�K]�����޹�)��&���A���\���w��@���~��Ѧ������g���.�ʺ�z׺�A�6��k���j��_���i���{3$�[*��}0���6���<��B�_�H���N�i U�I[�va�<g��%m��+s�X1y�g6�����p���<�����������S������}���mÚ��  �  Og=�=n�=�B=��=`~=�=� =�U =O��<p�<�S�<V��<���<���<p(�<&[�<ˌ�<V��<���<��<�G�<5s�<W��< ��</��<��<�6�<Y�<�y�<e��<D��<*��<��<���<��<''�<U7�<5E�<�P�<�Y�<�_�<�c�<�d�<c�<�^�<
W�<�L�<?�<s.�<��<��<<��<���<b��<ƅ�<�]�<�1�<��<z��<���<A^�<��<���<��<<N�<� �<��<�Y�<q �<A��<8B�<Vݿ<�t�<�<���<�#�<���<90�<��<\.�<��<Z�<9��<� �<�l�<֪<�;�<枧<���<�[�<,��<��<�b�<9��<L�<S�<���<�<l/�<�t�<���<���<�:�<�y�<`��<��<�.�<�h�<���<�ف<1�<�|<e�x<hu< �q<�=n<
�j<eg<}c<�_<�S\<}�X</.U<&�Q<�N<�J<4�F<�jC<V�?<�^<<��8<�]5<_�1<&j.<��*<݄'<5$<ǯ <�K<z�<��<�<<N�<��<C\	<�<Q�<�_�;}�;��;�w�;$E�; �;��; �;��;��;)=�;zo�;尶;��;�a�;�ѥ;�Q�;���;��;�.�;��;I��;���;�w;2m;�'c;�aY;�O;�0F;y�<;=x3;JH*;o5!;"?;�d;4�;Y�:��:��:el�:���:k��::��:d�q:��R:��3:�:���9f�9`p90�8\��6*׸J]�w����޹K(�:�&�Y�A���\�o�w�X@���~��Ŧ��>�������g�ʺ�z׺�A亢��$�����F_�������3$�=[*��}0�G�6�ٶ<���B�O�H�,�N�d U�H[�a��g��%m��+s�(1y�z6�ȝ��J���S�����������d���޴������oÚ��  �  Jg=�=k�=�B=��=[~=�=� =�U =I��<x�<�S�<S��<���<���<u(�<%[�<ٌ�<V��<���<��<�G�<4s�<K��<	��<0��<��<�6�<Y�<�y�<Y��<H��<.��<��<���<��<&'�<R7�<BE�<�P�<�Y�< `�<�c�<�d�<c�<�^�<W�<�L�<?�<o.�<��<��<I��<���<d��<���<�]�<�1�<�<���<���<C^�<��<���<���<6N�<� �<��<�Y�<h �<C��<:B�<Kݿ<�t�<�<���<�#�<���<:0�<��<b.�<��<a�<4��<� �<�l�<֪<<�<ܞ�<���<�[�<2��<��<�b�<G��<G�<S�<���<�<k/�<�t�<���<���< ;�<�y�<^��<��<�.�<�h�<���<�ف<&�<��|<Z�x<hu<�q<�=n<�j<Jg<}c<�_<�S\<}�X<.U<A�Q<�N<�J<*�F<�jC<c�?<�^<<��8<�]5<l�1<j.<��*<�'</$<̯ <�K<��<��<�<<M�<v�<R\	<�<N�<�_�;��;��;�w�;E�;��;	�;���;��;�;-=�;io�;���;��;�a�;ҥ;gQ�;���;��;�.�;��;+��;Ӛ�;{w;�m;�'c;gaY;�O;[0F;��<;$x3;UH*;:5!;�>;�d; �;0�:U��:��:sl�:>��:��:���:���:|�q:f�R:��3:Z�:7��9��9Rp9�.�84��6"׸�L]����޹�'�ڥ&�u�A�&�\�-�w��@���~��+���⹰�����ޢʺ�z׺�A����6�����1_������ ��3$��Z*�&~0�'�6�$�<���B���H��N�" U�y[�'a��g�s%m��+s�>1y�6�����G���������������:���ߴ������:Ú��  �  Ng=�=p�=�B=��=^~=�=� =�U =R��<w�<�S�<Q��<���<���<u(�<$[�<̌�<Y��<���<��<�G�<6s�<S��< ��<0��<��<�6�<Y�<�y�<c��<<��<-��<��<���<��<%'�<Y7�<3E�<�P�<�Y�<�_�<�c�<�d�<c�<�^�<
W�<�L�<?�<r.�<��<��<B��<���<b��<Ņ�<�]�<�1�<�<��<���<@^�<��<���<���<=N�<� �<��<�Y�<n �<@��<:B�<Vݿ<�t�<	�<���<�#�<���<:0�<��<V.�<��<]�<:��<� �<m�<֪<�;�<䞧<���<�[�<*��<��<�b�<:��<I�<S�<���<�<j/�<�t�<���<���<�:�<�y�<a��<��<�.�<�h�<���<�ف</�<�|<e�x<hu< �q<�=n<�j<tg<	}c<�_<�S\<p�X<).U<3�Q<�N<�J<>�F<�jC<W�?<�^<<��8<^5<R�1<,j.<��*<ڄ'<+$<ͯ <�K<��<��<�<<T�<|�<<\	<�<R�<�_�;~�;��;�w�;E�; �;��; �;��;��;0=�;po�;���;��;b�;�ѥ;�Q�;���;��;�.�;��;O��;���;�w;m;�'c;�aY;׹O;�0F;��<;x3;JH*;k5!;?;�d; �;��:��:��:ul�:���:6��:���:��:Z�q:�R:�3:
�:��9/�9�p96�8���6�׸�J]�C����޹%)���&���A�k�\���w�@���~��Ȧ��^�������<�ʺ{׺�A争�������*_�P����!��3$�[*��}0�}�6�ܶ<���B�u�H�7�N�o U� [�'a��g��%m��+s�K1y�{6�����[���4�����������^�����������VÚ��  �  Rg=�=r�=�B=��=]~=�=� =�U =T��<m�<�S�<Z��<���<���<j(�</[�<̌�<V��<���<��<�G�<+s�<R��<���<7��<��<�6�<Y�<�y�<m��<?��<3��<��<���<��<'�<a7�<-E�<�P�<�Y�<�_�<�c�<�d�<c�<�^�<
W�<�L�<?�<x.�<��<��<5��<���<e��<ą�<�]�<�1�<��<s��<�<>^�<��<���<���<=N�<� �<"��<�Y�<n �<F��<7B�<]ݿ<�t�<�<���<�#�<���<60�<��<U.�<!��<U�<@��<� �<�l�<֪<�;�<㞧<���<�[�<,��<��<�b�<6��<U�<S�<���<�<q/�<�t�<���<���<�:�<�y�<Y��<��<�.�<�h�<���<�ف<5�<�|<p�x<hu<��q<�=n<�j<}g<�|c<(�_<�S\<}�X<:.U<'�Q<�N<�J<E�F<�jC<T�?<�^<<��8<^5<S�1<1j.<��*<�'<>$<�� <�K<n�<
�<�<<N�<~�<<\	<�<<�<�_�;z�;<��;�w�;�D�;" �;��;> �;��;�;*=�;Ko�;���;��;"b�;�ѥ;�Q�;���;��;�.�;��;o��;���;�w;�m;�'c;�aY;��O;�0F;A�<;rx3;]H*;`5!;?;�d;i�;��:,��:{�:�l�:���:ެ�:��:���:��q:��R:��3:͇:w��9(�9p9�<�82
�6�׸�M]�2����޹;)�S�&��A���\���w�x@��~��񦣺d���,���١ʺ�z׺�A云��P���j�y_�L��2�����3$�`[*��}0�|�6���<���B�}�H�;�N�W U��[��a�jg��%m��+s�1y��6���������"���ڦ������[���ߴ��n���nÚ��  �  Pg=�=k�=�B=��=`~=�=� =�U =N��<y�<�S�<L��<���<���<j(�<"[�<֌�<Y��<���<��<�G�</s�<V��<��<'��<��<�6�<Y�<�y�<`��<A��<,��<��<���<��<"'�<Z7�<3E�<�P�<�Y�<�_�<�c�<�d�<c�<�^�<W�<�L�<?�<q.�<��<��<F��<���<Z��<ą�<�]�<�1�<��<���<���<<^�<��<���<���<=N�<� �<��<�Y�<m �<D��<5B�<Tݿ<�t�<�<���<�#�<���<=0�<��<W.�<��<Y�<;��<� �<�l�<֪<<�<垧<���<�[�<0��<��<�b�<D��<H�<S�<���<�<b/�<�t�<���<���<�:�<�y�<[��<��<�.�<�h�<���<�ف<4�<�|<X�x<
hu<�q<�=n<��j<sg<}c<$�_<�S\<{�X<$.U<3�Q<�N<�J<+�F<�jC<^�?<�^<<��8<�]5<X�1<$j.<��*<�'<"$<�� <�K<n�<�<�<<S�<z�<H\	<�<E�<�_�;��;���;�w�;E�; �;��;	 �;��;��;:=�;uo�;���;��;b�;�ѥ;�Q�;���;��;�.�;��;-��;���;�w;2m;�'c;{aY;ǹO;�0F;��<;Ix3;H*;\5!;?;�d;0�;�:���:d�:|l�:*��:R��:���:��:��q:��R:j�3:x�:���9��9lp9S4�8T��6�׸�I]����Q�޹�(���&�y�A�H�\���w��@��4������E���������ʺ�z׺�A云��r�����|_�<��3��d��3$��Z*��}0�w�6���<���B�Y�H��N�f U�z[�2a�ug��%m� ,s�61y�h6�����e���6�����������c���ⴔ�����VÚ��  �  Ig=�=l�=�B=��=[~=�=� =�U =L��<s�<�S�<U��< ��<���<{(�<![�<ˌ�<U��<���<��<�G�<;s�<L��<��<,��<��<�6�<Y�<�y�<Y��<L��<0��<��<���<��<%'�<W7�<?E�<�P�<�Y�<�_�<�c�<�d�<c�<�^�<W�<�L�<?�<t.�<��<��<>��<~��<h��<ȅ�<�]�<�1�<z�<z��<���<D^�<��<���<��<2N�<� �<��<�Y�<f �<@��<;B�<Sݿ<�t�<�<���<�#�<���<<0�<��<e.�<��<`�<3��<� �<	m�<
֪<<�<ڞ�<���<�[�<2��<��<�b�<9��<B�<S�<���<
�<n/�<�t�<���<���<�:�<�y�<b��<��<�.�<�h�<���<�ف<'�<�|<U�x<hu<�q<�=n<��j<Tg<}c<�_<�S\<��X<.U<<�Q<�N<�J<.�F<�jC<[�?<�^<<��8<�]5<f�1< j.<��*<ӄ'<2$<ӯ <�K<��<�<�<<K�<u�<M\	<�<]�<�_�;��;��;�w�;1E�;��;	�;���;��;�;0=�;^o�;���;��;�a�;ҥ;�Q�;���;��;�.�;��;.��;̚�;Ww;Bm;�'c;�aY;�O;�0F;��<;�w3;vH*;�5!;?; e;إ;\�:���:��:�l�:H��:���:L��:���:r�q:u�R:��3:��:H��9��9�p9�2�8���6�!׸9N]������޹8'�~�&���A�P�\���w��?���~��Z����������ޢʺ�z׺�A����!������^�G�������3$�)[*�~0�/�6��<���B���H�2�N�" U��[��a��g��%m�,s�1y�86�����b���t�����������I���Ĵ������BÚ��  �  Mg=�=n�=�B=��=^~=�=� =�U =T��<s�<�S�<_��<��<���<f(�<4[�<ь�<]��<���<��<�G�<1s�<S��<��<2��<��<�6�<Y�<�y�<c��<=��<,��<��<���<��<$'�<\7�<+E�<�P�<�Y�<`�<�c�<�d�<c�<�^�<W�<�L�<?�<u.�<��<��<:��<���<d��<���<�]�<�1�<��<x��<Ř�<>^�<��<���<��<<N�<� �<��<�Y�<g �<J��<>B�<Tݿ<�t�<	�<���<�#�<���<=0�<��<S.�<��<a�<<��<� �<�l�<֪< <�<䞧<���<�[�<,��<��<�b�<;��<X�<S�<���<��<t/�<�t�<���<���<�:�<�y�<W��<��<�.�<�h�<���<�ف<-�<��|<e�x<	hu<��q<�=n<�j<wg<	}c<(�_<�S\<x�X<,.U<A�Q<�N<�J<4�F<�jC<_�?<�^<<��8< ^5<W�1<0j.<��*<�'<H$<�� <�K<f�<�<�<<\�<{�<?\	<�<H�<�_�;��;'��;�w�;E�; �;	�; �;��;��;==�;so�;���;��;b�;�ѥ;�Q�;���;��;�.�;��;:��;���;�w;Im;�'c;�aY;��O;�0F;m�<;�x3;UH*; 5!;�>;�d;��;/�:X��:u�:�l�:+��:���:하:,��:��q:��R:��3:G�:��9��9Kp9�6�8���6�׸�I]�a����޹�)���&���A�7�\�}�w�[@���~������`���������ʺ�z׺�A�=�����Q��_���������W3$�3[*��}0�u�6�ж<���B�n�H��N�9 U�P[�Ea��g�k%m��+s�81y��6�����]���/�����������n���鴔�����:Ú��  �  �g=y=�=TC=i�=5=�=�� =�V =���<�<�V�<F��< ��<��<�+�<�^�<���<���<��<}�<�L�<Fx�<���<���<��<��< =�<�_�<{��<���<���<���<��<-�<3�<�/�<�@�<�N�<XZ�<�c�<>j�<Nn�<�o�<An�<�i�<�b�<�X�<^K�<;�<p'�<��<���<��<��<̓�<�k�<8@�<�<0��<���<Am�<1/�<+��<K��<�]�<�<���<%i�<��<���<�Q�<��<���<&�<���<\2�<T��<�>�<R��<K<�<ѵ�<�+�<c��<��<�y�<R�<�G�<���<
�<�f�<���<��<�l�<���<=�<�[�<���<��<�6�<�{�<��<� �<u@�<�<���<���<`2�<�k�<{��<)܁<�<ؒ|<m�x<2iu<I�q<=n<e�j<g<�yc<��_<�N\<g�X<5'U<P�Q<�N<^vJ<��F<-_C<�?<�Q<<��8<7O5<��1<�Y.<(�*<tr'<�$<�� <7<��<�{<(%<a�<��<�B	<�<I�<�(�;���;B~�;�<�;��;���;���;���;x��;3��;���;-�;n�;��;a�;���;��;���;;�;��;ڨ�;�w�;0V�;F�v;N�l; �b;c�X;5O;ɭE;lC<;��2;�);�� ;�;�;�.;��:�:�4�:א�:��:�٧:�Ǘ:��:=Zp:PEQ:��2:+:.�9Ao�9��j9$,�83 6p��9�a�\<��\�O2��'���B���]��x�!����薺�����}��)�ʺ��׺����D�U���>�c����d��$��N$��t*���0�&�6�Z�<�b�B���H��O��U�[��"a�*g��/m��4s��8y��<�����H���=���K���J��������������������  �  �g=y=�=WC=g�=8=�=� =�V =���<�<�V�<S��< ��<��<�+�<�^�<ʐ�<���<��<w�<�L�<Ox�<���<���<��<��< =�<�_�<���<���<���<���<��<1�<1�<�/�<w@�<�N�<^Z�<�c�<Sj�<Vn�<�o�<9n�<�i�<�b�<�X�<SK�<�:�<l'�<��<���<��</��<���<�k�<I@�<"�<7��<���<:m�</�<��<T��<�]�<
�<���<&i�<��<���<�Q�<��<ȃ�<�<���<[2�<W��<�>�<F��<X<�<ѵ�<�+�<t��<��<�y�<U�<�G�<}��<
�<�f�<���<��<~l�<���<F�<�[�<���<��<�6�<�{�<���<� �<u@�<�~�<���<���<\2�<�k�<q��<)܁<"�<��|<z�x<Giu<G�q<=n<s�j<�g<�yc<��_<�N\<��X<?'U<o�Q<	N<_vJ<��F<:_C<�?<�Q<<��8<�N5<��1<vY.<�*<�r'<$<�� <�6<��<�{<D%<E�<��<�B	<|<]�<�(�;���;S~�;�<�;��;���;���;���;���;��;���;-�;�m�;5��;$�;���;�;+��;X;�;�;٨�;�w�;CV�;�v;��l;Πb;��X;�4O;=�E;C<;�2;��);#� ;��;��;;/;�:�:~4�:|��:��:8ڧ:AǗ:��:�Yp:qEQ:��2:�:$�9�o�9��j9s�8]�6 ���a�G<��LṸ0� �'���B���]�j�x�F���_薺��������s�ʺ��׺,�人E�w����=����������#��N$��t*��0�!�6�7�<�s�B�u�H��O��U�Z[��"a��)g�`/m�x4s�X8y��<����,���c���5���u�������P���u���}����  �  �g={=�=ZC=b�=5=�=� =�V =���<�<�V�<H��<)��<��<,�<�^�<ʐ�<���<��<��<�L�<Wx�<���<���<��<��<=�<�_�<���<~��<���<���<��<6�<-�<�/�<o@�<�N�<YZ�<�c�<Bj�<Kn�<�o�<:n�<�i�<�b�<�X�<YK�<;�<�'�<��<���<��<-��<Ǔ�<�k�<K@�<�<<��<���<Pm�<)/�<!��<W��<�]�<�<���<,i�<��<���<�Q�<��<˃�<�<���<X2�<Y��<�>�<=��<]<�<ɵ�<�+�<c��<��<�y�<W�<�G�<s��<
�<�f�<���<��<~l�<���<2�<�[�<���<��<�6�<�{�< ��<� �<�@�<�~�<��<���<P2�<�k�<r��<.܁<�<�|<n�x<Ciu<G�q<�<n<��j<�g<�yc<��_<�N\<��X<0'U<[�Q<�N<fvJ<��F<C_C<��?<�Q<<��8<O5<��1<Y.<�*<zr'<�$<ț <�6<��<r{<D%<D�<��<�B	<�<k�<l(�;���;[~�;�<�;��;���;���;���;���;���;���;,-�;�m�;i��;�;���;��;	��;;�;��;�;�w�;SV�;ƈv;��l;��b;��X;�5O;C�E;�C<;|�2;��);i� ;��;��;�.;b�:�:�5�:_��:#�:mڧ:�Ɨ:��:�Yp:0FQ:}�2:�:��9n�9@�j9��8�K6��ฌ�a�:��m�"0��'���B���]��x����K薺D��p��g��K�ʺ@�׺$�亹E�L���k>���Q��P���#��N$��t*��0�S�6���<�>�B���H�[O�jU�N[��"a�,*g��/m��4s�i8y��<� �������m������v�������Z������������  �  �g=z=�=UC=h�=7=�=�� =�V =���<�<�V�<N��< ��<��<�+�<�^�<Ȑ�<���<��<p�<�L�<Gx�<���<���<��<��<"=�<�_�<���<���<���<���<��<1�<3�<�/�<}@�<�N�<YZ�<�c�<Mj�<Xn�<�o�<:n�<�i�<�b�<�X�<VK�< ;�<h'�<��<���<��<*��<Ó�<�k�<E@�<�<<��<���<9m�</�< ��<O��<�]�<	�<���<$i�<��<���<�Q�<��<�<�<���<Z2�<V��<�>�<E��<M<�<ֵ�<�+�<p��<��<�y�<S�<�G�<���<
�<�f�<���<��<�l�<���<@�<�[�<���<��<�6�<�{�<��<� �<p@�<�~�<���<���<\2�<�k�<t��<*܁<#�<�|<��x<(iu<M�q<=n<q�j<g<�yc<��_<�N\<b�X<O'U<k�Q<N<cvJ<��F<0_C<�?<�Q<<��8<%O5<{�1<wY.<$�*<�r'<$<�� <�6<��<�{<?%<L�<��<�B	<�<L�<�(�;��;F~�;�<�;��;���;���;��;���;��;���;-�;n�;<��;<�;���;��;D��;A;�;'�;ڨ�;�w�;1V�;;�v;|�l;�b;��X;�4O;D�E;�C<;��2;w�);H� ;��;l�;/;^�:�:h4�:���:�:�٧:�Ǘ:��:�Yp:EEQ:��2:+:f�9�o�9��j9�#�846,����a�o;����2�k�'�]�B�B�]��x�N����薺���n��?����ʺ��׺�亣E�����=�,��j������#��N$�qt*�	�0�O�6���<���B���H��O��U�D[��"a��)g�v/m�24s��8y�v<����/���=���7���h�����������T��������  �  �g=x=�=TC=h�=9=�=�� =�V =���<�<�V�<V��<��<��<�+�<�^�<���<���<'��<r�<�L�<Cx�<���<���<��<��<=�<�_�<x��<���<���<���<��<,�<3�<�/�<�@�<�N�<XZ�<�c�<;j�<Un�<�o�<Hn�<�i�<�b�<�X�<ZK�<;�<w'�<��<���<��<)��<���<�k�<C@�< �<,��<���<Km�<"/�<(��<M��<�]�< �<���<!i�<��<���<�Q�<��<Ã�<$�<���<[2�<U��<�>�<S��<N<�<Ե�<�+�<g��<��<�y�<Z�<�G�<���<
�<�f�<���<��<�l�<���<J�<�[�<���<��<�6�<�{�<���<� �<v@�<�~�<���<���<_2�<�k�<~��<%܁<$�<˒|<�x<0iu<X�q<=n<Z�j<	g<�yc<��_<�N\<m�X<G'U<E�Q<N<XvJ<��F<-_C<�?<�Q<<��8<'O5<��1<�Y.<�*<zr'<$<�� <�6<��<�{<.%<E�<ƈ<�B	<�<D�<�(�;���;W~�;�<�;��;���;���;���;���;B��;��;-�;n�;
��;P�;���;��;��;�:�;�;˨�;�w�;V�;T�v;x�l;�b;��X;E5O;��E;/C<;��2;p�);/� ;��;\�;2/;W�:��:�5�:��:��:�٧:�Ǘ:�:>[p:�DQ:l�2:I:��9io�9I�j9�*�8��6:��f�a��<�����1���'���B�]�]�Ϲx�4���薺���M�����h�ʺ��׺Ғ�tE�F����=�/��;������#��N$�u*���0��6���<���B�o�H��O��U��[�#a��)g�0m�c4s��8y�I<� ���^���L���_���n���k�������e��������  �  �g={=�=WC=e�=7=�=� =�V =���<�<�V�<E��<"��<��<�+�<�^�<ΐ�<���< ��<x�<�L�<Tx�<���<���<��<��<"=�<�_�<���<���<���<���<��<8�<+�< 0�<q@�<�N�<\Z�<�c�<Ej�<Tn�<�o�<:n�<�i�<�b�<�X�<\K�<�:�<y'�<��<���<��<&��<ȓ�<�k�<C@�<�<;��<���<Im�</�<#��<U��<�]�<�<���<(i�<��<���<�Q�<��<���<�<���<V2�<Z��<�>�<?��<Q<�<Ե�<�+�<i��<��<�y�<T�<�G�<���<
�<�f�<���<��<{l�<���<5�<�[�<���<��<�6�<�{�<���<� �<�@�<�~�<��<���<Z2�<�k�<q��<+܁<$�<�|<��x<;iu<B�q<�<n<��j<�g<�yc<��_<�N\<y�X<F'U<a�Q<N<dvJ<��F<7_C<�?<�Q<<��8<�N5<��1<�Y.<�*<�r'<�$<�� <�6<��<o{<L%<>�<��<�B	<<f�<�(�;���;L~�;�<�;��;���;���;���;���;���;���;4-�;�m�;j��;�;���;	�;:��;;�;�;娊;�w�;"V�;&�v;��l;�b;}�X;Q5O;G�E;�C<;��2;V�);s� ;��;b�;�.;S�:��:k5�:V��:<�:Iڧ:�Ǘ:D�:�Yp:�EQ:i�2:;:��9�o�9��j9��8�>6E����a��:���ṏ1���'���B��]�n�x�L���p薺���q�����F�ʺ��׺*���E�M���Z>���'��p��$��N$��t*�ٕ0�в6�5�<�4�B���H�O��U�\[��"a��)g��/m�Y4s��8y��<����񡅻��������x�������h���h��������  �  �g== �=XC=i�=1=�=� =�V =���<�<�V�<I��<-��<���<,�<�^�<֐�<���<��<��<�L�<Vx�<���<���<��<��<)=�<�_�<���<{��<���<���<��<5�< �<0�<o@�<�N�<SZ�<�c�<Kj�<On�<�o�<5n�<�i�<�b�<�X�<_K�<�:�<}'�<��<���<��<4��<�<�k�<S@�<�<F��<���<Lm�< /�<%��<V��<�]�<�<���<.i�<��<���<�Q�<��<у�<�<���<M2�<V��<�>�<D��<]<�<ŵ�<�+�<e��<��<�y�<S�<�G�<v��<
�<�f�<���<��<xl�<���<4�<�[�<���<��<�6�<�{�<	��<� �<�@�<�~�<	��<���<^2�<�k�<k��<3܁<�<��|<k�x<3iu<c�q<�<n<��j<�g<�yc<��_<�N\<w�X</'U<s�Q<�N<vvJ<��F<<_C<�?<vQ<<��8<�N5<��1<oY.< �*<�r'<�$<ћ <�6<��<s{<[%<>�<��<�B	<�<i�<a(�;��;N~�;�<�;	�;���;���;���;���;��;���;'-�;�m�;���;�;㍥;��;(��;8;�;�;���;w�;HV�;�v;��l;-�b;��X;o5O;�E;�C<;��2;��);;� ;��;��;�.;�:k�:�5�:Ï�:a�:Sڧ:Ǘ:��:PYp:wFQ:
�2:�:Q�9�l�9��j9��8�6����a��9����0���'���B���]��x�?����薺���G�����.�ʺ�׺k��!F����Z>����߽�M���#��N$�^t*�B�0���6�6�<��B���H��O��U��[��"a�#*g�V/m��4s��8y�<�2���ꡅ�������������l���j�������t����  �  �g=~=�=SC=h�=4=�=� =�V =���<�<�V�<K��<.��<��<
,�<�^�<Ő�<���<!��<w�<�L�<Nx�<���<���<��<��<$=�<�_�<���<���<���<���<��<4�<5�<�/�<q@�<�N�<WZ�<�c�<Aj�<Nn�<�o�<Bn�<�i�<�b�<�X�<]K�< ;�<{'�<��<���<��<0��<Ɠ�<�k�<N@�<�<7��<���<Lm�</�<&��<P��<�]�<�<���<,i�<��<���<�Q�<��<ƃ�<�<���<]2�<[��<�>�<F��<P<�<ѵ�<�+�<b��<��<�y�<S�<�G�<{��<
�<�f�<���<��<�l�<���<7�<�[�<���<��<�6�<�{�<��<� �<�@�<�~�< ��<���<^2�<�k�<y��<1܁<�<�|<��x</iu<Y�q<�<n<v�j<
g<�yc<��_<�N\<h�X<F'U<`�Q<�N<qvJ<��F<'_C<�?<�Q<<��8<O5<��1<�Y.<�*<qr'<�$<қ <�6<��<{<9%<I�<��<�B	<�<Z�<w(�;���;B~�;�<�;��;���;���;���;���;��;p��;#-�;n�;<��;�;���;��;1��;;�;��;���;�w�;V�;&�v;v�l;�b;��X;d5O;g�E;�C<;��2;��);`� ;��;��;�.;�:H�:�5�:���:v�:�٧:VǗ:<�:uZp:DFQ:ˆ2:�:��9|n�9��j9��8��6��ม�a�=��.Ṻ1��'�7�B���]�p�x�����{薺e����������ʺ��׺�亠E����D>����y��8���#�O$��t*��0�̲6���<�Y�B���H��O��U�[��"a�(*g��/m�_4s��8y�E<�9���&���J���'�������o�������g��������  �  �g=t=	�=UC=g�=9=�=� =�V =���<�<�V�<L��<��<��<�+�<�^�<͐�<���<��<k�<�L�<Gx�<���<���<��<��<=�<�_�<}��<���<���<���<��<-�<2�<�/�<�@�<�N�<`Z�<�c�<Dj�<Yn�<�o�<Dn�<�i�<�b�<�X�<ZK�<�:�<l'�<��<���<"��<%��<ē�<�k�<=@�<$�<8��<���<<m�</�<%��<K��<�]�< �<���<"i�<��<���<�Q�<��<���<"�<���<X2�<R��<�>�<L��<D<�<ߵ�<�+�<p��<��<�y�<X�<�G�<���<
�<�f�<���<��<|l�<���<E�<�[�<���<��<�6�<�{�<���<� �<r@�<�~�<���<���<^2�<�k�<}��<܁<+�<ג|<��x<1iu<<�q<=n<m�j< g<�yc<��_<�N\<e�X<['U<O�Q<N<KvJ<��F<1_C<�?<�Q<<��8<O5<z�1<�Y.<�*<�r'<�$<�� <�6<��<�{<J%<?�<��<�B	<�<L�<�(�;���;W~�;�<�;��;���;���;��;l��; ��;���;-�;n�;5��;Z�;t��;�;E��;;�;+�;Ĩ�;�w�;V�;]�v;o�l;�b;��X;�4O;c�E;�C<;1�2;N�);P� ;��;/�;Q/;�:.�:�4�:L��:l�:�٧:�Ǘ:�:�Zp:�DQ:̇2:x:��9�q�9��j9+(�8��6J����a��;���	�)3�T�'���B�.�]���x�#���/薺�����h����ʺ�׺����E�b����=����2������#�xN$��t*�Е0�<�6���<���B�s�H��O��U��[�2#a��)g��/m�4s��8y��<�����9���_���A���H�����������=��������  �  �g=v=�=VC=f�=6=�=� =�V =���<�<�V�<P��<��<��<�+�<�^�<Ȑ�<���<&��<~�<�L�<Mx�<���<���<��<��<=�<�_�<u��<���<���<���<��<0�<-�<�/�<z@�<�N�<[Z�<�c�<@j�<Pn�<�o�<Bn�<�i�<�b�<�X�<`K�<;�<�'�<��<���<��<+��<ē�<�k�<G@�<�<7��<���<Om�<%/�<*��<N��<�]�<	�<���<&i�<��<���<�Q�<��<Ń�<�<���<V2�<U��<�>�<J��<W<�<ϵ�<�+�<k��<��<�y�<U�<�G�<|��<
�<�f�<���<��<{l�<���<A�<�[�<���<��<�6�<�{�<���<� �<�@�<�~�< ��<���<[2�<�k�<y��<#܁<&�<Ԓ|<m�x<@iu<K�q<=n<r�j<�g<�yc<��_<�N\<�X<6'U<H�Q<N<PvJ<��F<4_C<�?<�Q<<��8<O5<��1<�Y.<�*<r'<$<�� <7<��<�{<A%<:�<ň<�B	<�<X�<�(�;���;L~�;�<�;��;���;w��;���;���;&��;���;-�;�m�;6��;3�;���;�;���;;�;�;٨�;�w�;?V�;!�v;q�l;5�b;��X;�5O;r�E;�C<;��2;��);M� ;��;{�;	/;�::�:�5�:"��:��:�٧:WǗ:��:�Zp:sEQ:��2:�:��9o�9��j9�!�8�6���\�a��;��6
��0�F�'�P�B���]�O�x�#���\薺N����� ����ʺ��׺֒��E�����=���.������#��N$��t*���0���6���<�V�B���H� O��U�[�#a��)g��/m��4s�v8y�~<����.���q���3���m�������[������������  �  �g=}=�=PC=k�=5=�=� =�V =���<�<�V�<N��<*��<��<	,�<�^�<ǐ�<���<��<u�<�L�<Rx�<���<���<���<��<#=�<�_�<���<���<���<���<��<7�</�<�/�<m@�<�N�<[Z�<�c�<Wj�<Mn�<�o�<1n�<�i�<�b�<�X�<WK�<�:�<s'�<��<���<��<3��<œ�<�k�<O@�<�<B��<���<Bm�</�< ��<T��<�]�<�<~��</i�<��<���<�Q�<��<ǃ�<�<���<Y2�<[��<�>�<>��<S<�<е�<�+�<o��<��<�y�<H�<�G�<|��<
�<�f�<���<��<l�<���<6�<�[�<���<��<�6�<�{�<	��<� �<{@�<�~�<���<���<a2�<�k�<n��<2܁<�<�|<y�x<6iu<M�q<�<n<��j< g<�yc<��_<�N\<s�X<?'U<��Q<�N<nvJ<��F<_C< �?<�Q<<��8<O5<��1<qY.<%�*<tr'<$<ʛ <�6<��<z{<>%<N�<��<�B	<|<a�<�(�;��;~�;�<�;��;���;���;���;���;���;���;.-�;�m�;X��;��;���;�;7��;h;�;��;��;nw�;5V�;5�v;��l;�b;��X;5O;�E;�C<;}�2;��);Y� ;��;��;�.;��:��:�4�:_��:�:>ڧ:jǗ:��:�Xp:�FQ:��2:�:P�9zo�9��j9��8�65����a�w;��F�Y1�:�'���B�V�]���x��/閺���������h�ʺ��׺œ亮E�f���Q>����j��J���#�O$�^t*�+�0��6�5�<�t�B���H��O��U�n[��"a�*g�/m�z4s��8y�t<�3������_��������������t���v���U����  �  �g=z=�=UC=i�=3=�=� =�V =���<�<�V�<L��<��<��<�+�<�^�<ǐ�<���<��<��<�L�<Lx�<���<���<��<��<=�<�_�<z��<���<���<���<��<0�<'�<�/�<�@�<�N�<ZZ�<�c�<Dj�<Jn�<�o�<;n�<�i�<�b�<�X�<]K�<;�<|'�<��<���<��<)��<œ�<�k�<C@�<�<>��<���<Km�<+/�<(��<O��<�]�<
�<���<+i�<��<���<�Q�<��<�<!�<���<P2�<S��<�>�<P��<N<�<ϵ�<�+�<e��<��<�y�<S�<�G�<z��<
�<�f�<���<��<�l�<���<<�<�[�<���<��<�6�<�{�<��<� �<�@�<�~�<���<���<_2�<�k�<v��<+܁<�<�|<d�x<5iu<Q�q<=n<w�j<�g<�yc<��_<�N\<m�X<2'U<T�Q<�N<avJ<��F<1_C<�?<~Q<<��8<O5<��1<Y.<'�*<}r'<�$<�� <�6<��<�{<=%<T�<��<�B	<�<V�<|(�;��;G~�;�<�;��;���;���;���;���;4��;���;-�;�m�;G��;L�;���;�;�;;�;��;�;�w�;?V�;/�v;v�l;�b;�X;m5O;S�E;�C<;��2;k�);[� ;��;c�;�.;x�:7�:�5�:}��:��:�٧:RǗ:��:�Yp:FQ:L�2:�:(�9;o�9��j9�'�8�6�����a��:�����1�Z�'���B���]�n�x������薺�����-����ʺ��׺C��kE�v���>�%��Q������#��N$�kt*���0���6���<�k�B���H��O��U�/[��"a�3*g��/m��4s��8y�f<�򟂻#�������-���U�������������������  �  �g=x=�=WC=f�=8=�=� =�V =���<�<�V�<U��<��<��<�+�<�^�<Ɛ�<���<��<q�<�L�<Lx�<���<���<��<��<!=�<�_�<{��<���<���<���<��<7�<:�<�/�<w@�<�N�<hZ�<�c�<Oj�<^n�<�o�<@n�<�i�<�b�<�X�<WK�<�:�<m'�<��<���<!��<'��<Ó�<�k�<?@�<&�<5��<���<;m�</�<��<N��<�]�<�<���<"i�<��<���<�Q�<��<���<�<���<b2�<^��<�>�<E��<N<�<൲<�+�<��<��<�y�<W�<�G�<���<
�<�f�<���<��<|l�<���<K�<�[�<���<��<�6�<�{�<���<� �<u@�<�~�<���<���<[2�<�k�<v��<#܁</�<�|<}�x<Qiu<6�q<�<n<j�j<g<�yc<��_<�N\<��X<O'U<V�Q<&N<YvJ<��F<7_C<�?<�Q<<��8<O5<��1<vY.<�*<�r'<$<�� < 7<��<�{<<%<B�<��<�B	<�<V�<�(�;���;V~�;�<�;��;��;���;��;���;��;]��;.-�;"n�;��;'�;y��;9�;��;K;�;<�;ʨ�;�w�;6V�;#�v;w�l;�b;~�X;�4O;]�E;lC<;*�2;Z�);I� ;��;@�;Z/;��: �:�4�:&��:��:�٧:qǗ:��:�Zp:�DQ:A�2:,:��9�r�9��j9u�8{6b���a�F?��s��1�,�'�Q�B�X�]�q�x�����C薺R��u��&��/�ʺ��׺����E�����=�e��/������#��N$��t*��0�&�6�*�<�j�B�z�H�O��U�2[�#a�q)g��/m�k4s�28y��<����>���F���8�����������J���T��������  �  �g=z=�=UC=i�=3=�=� =�V =���<�<�V�<L��<��<��<�+�<�^�<ǐ�<���<��<��<�L�<Lx�<���<���<��<��<=�<�_�<z��<���<���<���<��<0�<'�<�/�<�@�<�N�<ZZ�<�c�<Dj�<Jn�<�o�<;n�<�i�<�b�<�X�<]K�<;�<|'�<��<���<��<)��<œ�<�k�<C@�<�<>��<���<Km�<+/�<(��<O��<�]�<
�<���<+i�<��<���<�Q�<��<�<!�<���<P2�<S��<�>�<P��<N<�<ϵ�<�+�<e��<��<�y�<S�<�G�<z��<
�<�f�<���<��<�l�<���<<�<�[�<���<��<�6�<�{�<��<� �<�@�<�~�<���<���<_2�<�k�<v��<+܁<�<�|<d�x<5iu<Q�q<=n<w�j<�g<�yc<��_<�N\<m�X<2'U<T�Q<�N<avJ<��F<1_C<�?<~Q<<��8<O5<��1<Y.<'�*<}r'<�$<�� <�6<��<�{<=%<T�<��<�B	<�<V�<|(�;��;G~�;�<�;��;���;���;���;���;4��;���;-�;�m�;G��;L�;���;�;�;;�;��;�;�w�;?V�;/�v;v�l;�b;�X;m5O;S�E;�C<;��2;k�);[� ;��;c�;�.;x�:7�:�5�:}��:��:�٧:RǗ:��:�Yp:FQ:L�2:�:(�9;o�9��j9�'�8�6�����a��:�����1�Z�'���B���]�n�x������薺�����-����ʺ��׺C��kE�v���>�%��Q������#��N$�kt*���0���6���<�k�B���H��O��U�/[��"a�3*g��/m��4s��8y�f<�򟂻#�������-���U�������������������  �  �g=}=�=PC=k�=5=�=� =�V =���<�<�V�<N��<*��<��<	,�<�^�<ǐ�<���<��<u�<�L�<Rx�<���<���<���<��<#=�<�_�<���<���<���<���<��<7�</�<�/�<m@�<�N�<[Z�<�c�<Wj�<Mn�<�o�<1n�<�i�<�b�<�X�<WK�<�:�<s'�<��<���<��<3��<œ�<�k�<O@�<�<B��<���<Bm�</�< ��<T��<�]�<�<~��</i�<��<���<�Q�<��<ǃ�<�<���<Y2�<[��<�>�<>��<S<�<е�<�+�<o��<��<�y�<H�<�G�<|��<
�<�f�<���<��<l�<���<6�<�[�<���<��<�6�<�{�<	��<� �<{@�<�~�<���<���<a2�<�k�<n��<2܁<�<�|<y�x<6iu<M�q<�<n<��j< g<�yc<��_<�N\<s�X<?'U<��Q<�N<nvJ<��F<_C< �?<�Q<<��8<O5<��1<qY.<%�*<tr'<$<ʛ <�6<��<z{<>%<N�<��<�B	<|<a�<�(�;��;~�;�<�;��;���;���;���;���;���;���;.-�;�m�;X��;��;���;�;7��;h;�;��;��;nw�;5V�;5�v;��l;�b;��X;5O;�E;�C<;}�2;��);Y� ;��;��;�.;��:��:�4�:_��:�:>ڧ:jǗ:��:�Xp:�FQ:��2:�:P�9zo�9��j9��8�65����a�w;��F�Y1�:�'���B�V�]���x��/閺���������h�ʺ��׺œ亮E�f���Q>����j��J���#�O$�^t*�+�0��6�5�<�t�B���H��O��U�n[��"a�*g�/m�z4s��8y�t<�3������_��������������t���v���U����  �  �g=v=�=VC=f�=6=�=� =�V =���<�<�V�<P��<��<��<�+�<�^�<Ȑ�<���<&��<~�<�L�<Mx�<���<���<��<��<=�<�_�<u��<���<���<���<��<0�<-�<�/�<z@�<�N�<[Z�<�c�<@j�<Pn�<�o�<Bn�<�i�<�b�<�X�<`K�<;�<�'�<��<���<��<+��<ē�<�k�<G@�<�<7��<���<Om�<%/�<*��<N��<�]�<	�<���<&i�<��<���<�Q�<��<Ń�<�<���<V2�<U��<�>�<J��<W<�<ϵ�<�+�<k��<��<�y�<U�<�G�<|��<
�<�f�<���<��<{l�<���<A�<�[�<���<��<�6�<�{�<���<� �<�@�<�~�< ��<���<[2�<�k�<y��<#܁<&�<Ԓ|<m�x<@iu<K�q<=n<r�j<�g<�yc<��_<�N\<�X<6'U<H�Q<N<PvJ<��F<4_C<�?<�Q<<��8<O5<��1<�Y.<�*<r'<$<�� <7<��<�{<A%<:�<ň<�B	<�<X�<�(�;���;L~�;�<�;��;���;w��;���;���;&��;���;-�;�m�;6��;3�;���;�;���;;�;�;٨�;�w�;?V�;!�v;q�l;5�b;��X;�5O;r�E;�C<;��2;��);M� ;��;{�;	/;�::�:�5�:"��:��:�٧:WǗ:��:�Zp:sEQ:��2:�:��9o�9��j9�!�8�6���\�a��;��6
��0�F�'�P�B���]�O�x�#���\薺N����� ����ʺ��׺֒��E�����=���.������#��N$��t*���0���6���<�V�B���H� O��U�[�#a��)g��/m��4s�v8y�~<����.���q���3���m�������[������������  �  �g=t=	�=UC=g�=9=�=� =�V =���<�<�V�<L��<��<��<�+�<�^�<͐�<���<��<k�<�L�<Gx�<���<���<��<��<=�<�_�<}��<���<���<���<��<-�<2�<�/�<�@�<�N�<`Z�<�c�<Dj�<Yn�<�o�<Dn�<�i�<�b�<�X�<ZK�<�:�<l'�<��<���<"��<%��<ē�<�k�<=@�<$�<8��<���<<m�</�<%��<K��<�]�< �<���<"i�<��<���<�Q�<��<���<"�<���<X2�<R��<�>�<L��<D<�<ߵ�<�+�<p��<��<�y�<X�<�G�<���<
�<�f�<���<��<|l�<���<E�<�[�<���<��<�6�<�{�<���<� �<r@�<�~�<���<���<^2�<�k�<}��<܁<+�<ג|<��x<1iu<<�q<=n<m�j< g<�yc<��_<�N\<e�X<['U<O�Q<N<KvJ<��F<1_C<�?<�Q<<��8<O5<z�1<�Y.<�*<�r'<�$<�� <�6<��<�{<J%<?�<��<�B	<�<L�<�(�;���;W~�;�<�;��;���;���;��;l��; ��;���;-�;n�;5��;Z�;t��;�;E��;;�;+�;Ĩ�;�w�;V�;]�v;o�l;�b;��X;�4O;c�E;�C<;1�2;N�);P� ;��;/�;Q/;�:.�:�4�:L��:l�:�٧:�Ǘ:�:�Zp:�DQ:̇2:x:��9�q�9��j9+(�8��6J����a��;���	�)3�T�'���B�.�]���x�#���/薺�����h����ʺ�׺����E�b����=����2������#�xN$��t*�Е0�<�6���<���B�s�H��O��U��[�2#a��)g��/m�4s��8y��<�����9���_���A���H�����������=��������  �  �g=~=�=SC=h�=4=�=� =�V =���<�<�V�<K��<.��<��<
,�<�^�<Ő�<���<!��<w�<�L�<Nx�<���<���<��<��<$=�<�_�<���<���<���<���<��<4�<5�<�/�<q@�<�N�<WZ�<�c�<Aj�<Nn�<�o�<Bn�<�i�<�b�<�X�<]K�< ;�<{'�<��<���<��<0��<Ɠ�<�k�<N@�<�<7��<���<Lm�</�<&��<P��<�]�<�<���<,i�<��<���<�Q�<��<ƃ�<�<���<]2�<[��<�>�<F��<P<�<ѵ�<�+�<b��<��<�y�<S�<�G�<{��<
�<�f�<���<��<�l�<���<7�<�[�<���<��<�6�<�{�<��<� �<�@�<�~�< ��<���<^2�<�k�<y��<1܁<�<�|<��x</iu<Y�q<�<n<v�j<
g<�yc<��_<�N\<h�X<F'U<`�Q<�N<qvJ<��F<'_C<�?<�Q<<��8<O5<��1<�Y.<�*<qr'<�$<қ <�6<��<{<9%<I�<��<�B	<�<Z�<w(�;���;B~�;�<�;��;���;���;���;���;��;p��;#-�;n�;<��;�;���;��;1��;;�;��;���;�w�;V�;&�v;v�l;�b;��X;d5O;g�E;�C<;��2;��);`� ;��;��;�.;�:H�:�5�:���:v�:�٧:VǗ:<�:uZp:DFQ:ˆ2:�:��9|n�9��j9��8��6��ม�a�=��.Ṻ1��'�7�B���]�p�x�����{薺e����������ʺ��׺�亠E����D>����y��8���#�O$��t*��0�̲6���<�Y�B���H��O��U�[��"a�(*g��/m�_4s��8y�E<�9���&���J���'�������o�������g��������  �  �g== �=XC=i�=1=�=� =�V =���<�<�V�<I��<-��<���<,�<�^�<֐�<���<��<��<�L�<Vx�<���<���<��<��<)=�<�_�<���<{��<���<���<��<5�< �<0�<o@�<�N�<SZ�<�c�<Kj�<On�<�o�<5n�<�i�<�b�<�X�<_K�<�:�<}'�<��<���<��<4��<�<�k�<S@�<�<F��<���<Lm�< /�<%��<V��<�]�<�<���<.i�<��<���<�Q�<��<у�<�<���<M2�<V��<�>�<D��<]<�<ŵ�<�+�<e��<��<�y�<S�<�G�<v��<
�<�f�<���<��<xl�<���<4�<�[�<���<��<�6�<�{�<	��<� �<�@�<�~�<	��<���<^2�<�k�<k��<3܁<�<��|<k�x<3iu<c�q<�<n<��j<�g<�yc<��_<�N\<w�X</'U<s�Q<�N<vvJ<��F<<_C<�?<vQ<<��8<�N5<��1<oY.< �*<�r'<�$<ћ <�6<��<s{<[%<>�<��<�B	<�<i�<a(�;��;N~�;�<�;	�;���;���;���;���;��;���;'-�;�m�;���;�;㍥;��;(��;8;�;�;���;w�;HV�;�v;��l;-�b;��X;o5O;�E;�C<;��2;��);;� ;��;��;�.;�:k�:�5�:Ï�:a�:Sڧ:Ǘ:��:PYp:wFQ:
�2:�:Q�9�l�9��j9��8�6����a��9����0���'���B���]��x�?����薺���G�����.�ʺ�׺k��!F����Z>����߽�M���#��N$�^t*�B�0���6�6�<��B���H��O��U��[��"a�#*g�V/m��4s��8y�<�2���ꡅ�������������l���j�������t����  �  �g={=�=WC=e�=7=�=� =�V =���<�<�V�<E��<"��<��<�+�<�^�<ΐ�<���< ��<x�<�L�<Tx�<���<���<��<��<"=�<�_�<���<���<���<���<��<8�<+�< 0�<q@�<�N�<\Z�<�c�<Ej�<Tn�<�o�<:n�<�i�<�b�<�X�<\K�<�:�<y'�<��<���<��<&��<ȓ�<�k�<C@�<�<;��<���<Im�</�<#��<U��<�]�<�<���<(i�<��<���<�Q�<��<���<�<���<V2�<Z��<�>�<?��<Q<�<Ե�<�+�<i��<��<�y�<T�<�G�<���<
�<�f�<���<��<{l�<���<5�<�[�<���<��<�6�<�{�<���<� �<�@�<�~�<��<���<Z2�<�k�<q��<+܁<$�<�|<��x<;iu<B�q<�<n<��j<�g<�yc<��_<�N\<y�X<F'U<a�Q<N<dvJ<��F<7_C<�?<�Q<<��8<�N5<��1<�Y.<�*<�r'<�$<�� <�6<��<o{<L%<>�<��<�B	<<f�<�(�;���;L~�;�<�;��;���;���;���;���;���;���;4-�;�m�;j��;�;���;	�;:��;;�;�;娊;�w�;"V�;&�v;��l;�b;}�X;Q5O;G�E;�C<;��2;V�);s� ;��;b�;�.;S�:��:k5�:V��:<�:Iڧ:�Ǘ:D�:�Yp:�EQ:i�2:;:��9�o�9��j9��8�>6E����a��:���ṏ1���'���B��]�n�x�L���p薺���q�����F�ʺ��׺*���E�M���Z>���'��p��$��N$��t*�ٕ0�в6�5�<�4�B���H�O��U�\[��"a��)g��/m�Y4s��8y��<����񡅻��������x�������h���h��������  �  �g=x=�=TC=h�=9=�=�� =�V =���<�<�V�<V��<��<��<�+�<�^�<���<���<'��<r�<�L�<Cx�<���<���<��<��<=�<�_�<x��<���<���<���<��<,�<3�<�/�<�@�<�N�<XZ�<�c�<;j�<Un�<�o�<Hn�<�i�<�b�<�X�<ZK�<;�<w'�<��<���<��<)��<���<�k�<C@�< �<,��<���<Km�<"/�<(��<M��<�]�< �<���<!i�<��<���<�Q�<��<Ã�<$�<���<[2�<U��<�>�<S��<N<�<Ե�<�+�<g��<��<�y�<Z�<�G�<���<
�<�f�<���<��<�l�<���<J�<�[�<���<��<�6�<�{�<���<� �<v@�<�~�<���<���<_2�<�k�<~��<%܁<$�<˒|<�x<0iu<X�q<=n<Z�j<	g<�yc<��_<�N\<m�X<G'U<E�Q<N<XvJ<��F<-_C<�?<�Q<<��8<'O5<��1<�Y.<�*<zr'<$<�� <�6<��<�{<.%<E�<ƈ<�B	<�<D�<�(�;���;W~�;�<�;��;���;���;���;���;B��;��;-�;n�;
��;P�;���;��;��;�:�;�;˨�;�w�;V�;T�v;x�l;�b;��X;E5O;��E;/C<;��2;p�);/� ;��;\�;2/;W�:��:�5�:��:��:�٧:�Ǘ:�:>[p:�DQ:l�2:I:��9io�9I�j9�*�8��6:��f�a��<�����1���'���B�]�]�Ϲx�4���薺���M�����h�ʺ��׺Ғ�tE�F����=�/��;������#��N$�u*���0��6���<���B�o�H��O��U��[�#a��)g�0m�c4s��8y�I<� ���^���L���_���n���k�������e��������  �  �g=z=�=UC=h�=7=�=�� =�V =���<�<�V�<N��< ��<��<�+�<�^�<Ȑ�<���<��<p�<�L�<Gx�<���<���<��<��<"=�<�_�<���<���<���<���<��<1�<3�<�/�<}@�<�N�<YZ�<�c�<Mj�<Xn�<�o�<:n�<�i�<�b�<�X�<VK�< ;�<h'�<��<���<��<*��<Ó�<�k�<E@�<�<<��<���<9m�</�< ��<O��<�]�<	�<���<$i�<��<���<�Q�<��<�<�<���<Z2�<V��<�>�<E��<M<�<ֵ�<�+�<p��<��<�y�<S�<�G�<���<
�<�f�<���<��<�l�<���<@�<�[�<���<��<�6�<�{�<��<� �<p@�<�~�<���<���<\2�<�k�<t��<*܁<#�<�|<��x<(iu<M�q<=n<q�j<g<�yc<��_<�N\<b�X<O'U<k�Q<N<cvJ<��F<0_C<�?<�Q<<��8<%O5<{�1<wY.<$�*<�r'<$<�� <�6<��<�{<?%<L�<��<�B	<�<L�<�(�;��;F~�;�<�;��;���;���;��;���;��;���;-�;n�;<��;<�;���;��;D��;A;�;'�;ڨ�;�w�;1V�;;�v;|�l;�b;��X;�4O;D�E;�C<;��2;w�);H� ;��;l�;/;^�:�:h4�:���:�:�٧:�Ǘ:��:�Yp:EEQ:��2:+:f�9�o�9��j9�#�846,����a�o;����2�k�'�]�B�B�]��x�N����薺���n��?����ʺ��׺�亣E�����=�,��j������#��N$�qt*�	�0�O�6���<���B���H��O��U�D[��"a��)g�v/m�24s��8y�v<����/���=���7���h�����������T��������  �  �g={=�=ZC=b�=5=�=� =�V =���<�<�V�<H��<)��<��<,�<�^�<ʐ�<���<��<��<�L�<Wx�<���<���<��<��<=�<�_�<���<~��<���<���<��<6�<-�<�/�<o@�<�N�<YZ�<�c�<Bj�<Kn�<�o�<:n�<�i�<�b�<�X�<YK�<;�<�'�<��<���<��<-��<Ǔ�<�k�<K@�<�<<��<���<Pm�<)/�<!��<W��<�]�<�<���<,i�<��<���<�Q�<��<˃�<�<���<X2�<Y��<�>�<=��<]<�<ɵ�<�+�<c��<��<�y�<W�<�G�<s��<
�<�f�<���<��<~l�<���<2�<�[�<���<��<�6�<�{�< ��<� �<�@�<�~�<��<���<P2�<�k�<r��<.܁<�<�|<n�x<Ciu<G�q<�<n<��j<�g<�yc<��_<�N\<��X<0'U<[�Q<�N<fvJ<��F<C_C<��?<�Q<<��8<O5<��1<Y.<�*<zr'<�$<ț <�6<��<r{<D%<D�<��<�B	<�<k�<l(�;���;[~�;�<�;��;���;���;���;���;���;���;,-�;�m�;i��;�;���;��;	��;;�;��;�;�w�;SV�;ƈv;��l;��b;��X;�5O;C�E;�C<;|�2;��);i� ;��;��;�.;b�:�:�5�:_��:#�:mڧ:�Ɨ:��:�Yp:0FQ:}�2:�:��9n�9@�j9��8�K6��ฌ�a�:��m�"0��'���B���]��x����K薺D��p��g��K�ʺ@�׺$�亹E�L���k>���Q��P���#��N$��t*��0�S�6���<�>�B���H�[O�jU�N[��"a�,*g��/m��4s�i8y��<� �������m������v�������Z������������  �  �g=y=�=WC=g�=8=�=� =�V =���<�<�V�<S��< ��<��<�+�<�^�<ʐ�<���<��<w�<�L�<Ox�<���<���<��<��< =�<�_�<���<���<���<���<��<1�<1�<�/�<w@�<�N�<^Z�<�c�<Sj�<Vn�<�o�<9n�<�i�<�b�<�X�<SK�<�:�<l'�<��<���<��</��<���<�k�<I@�<"�<7��<���<:m�</�<��<T��<�]�<
�<���<&i�<��<���<�Q�<��<ȃ�<�<���<[2�<W��<�>�<F��<X<�<ѵ�<�+�<t��<��<�y�<U�<�G�<}��<
�<�f�<���<��<~l�<���<F�<�[�<���<��<�6�<�{�<���<� �<u@�<�~�<���<���<\2�<�k�<q��<)܁<"�<��|<z�x<Giu<G�q<=n<s�j<�g<�yc<��_<�N\<��X<?'U<o�Q<	N<_vJ<��F<:_C<�?<�Q<<��8<�N5<��1<vY.<�*<�r'<$<�� <�6<��<�{<D%<E�<��<�B	<|<]�<�(�;���;S~�;�<�;��;���;���;���;���;��;���;-�;�m�;5��;$�;���;�;+��;X;�;�;٨�;�w�;CV�;�v;��l;Πb;��X;�4O;=�E;C<;�2;��);#� ;��;��;;/;�:�:~4�:|��:��:8ڧ:AǗ:��:�Yp:qEQ:��2:�:$�9�o�9��j9s�8]�6 ���a�G<��LṸ0� �'���B���]�j�x�F���_薺��������s�ʺ��׺,�人E�w����=����������#��N$��t*��0�!�6�7�<�s�B�u�H��O��U�Z[��"a��)g�`/m�x4s�X8y��<����,���c���5���u�������P���u���}����  �  ;h==��=(D=V�=6�=�=6� =.X =���<4"�<�Y�<��<���<��<U0�<�c�<���<���<���<&%�<�R�<�~�<)��<m��<%��<W �<�D�<�g�<��<A��<���<H��<���<C�<�'�<�:�<�K�<Z�<4f�<�o�<�v�<<{�<�|�<�{�<�w�<q�<@g�<dZ�<hJ�<(7�<� �<��<���<��<��</}�<�Q�<�"�<@��<��<��<�A�<���<��<rp�<�"�<|��<|�<�"�<���<]d�<Q��<P��<�)�<ḻ<wD�<8̸<IP�<�е<fM�<�Ʋ<J<�<���<m�<��<_�<�V�<���<��<!t�<�͢<P$�<tx�<�ɝ<+�<�e�<���<��<�?�<��<�Ƒ<��<@G�<5��<���<���<�6�<�o�<�<߁<{�<��|<y<�ju<��q<L<n<��j<)g<�uc<��_<xH\<�X<�U<ɋQ<L�M<�jJ<��F<FQC<�?<UA<<��8<�<5<H�1<3E.<��*< \'<��#<1� <W<?�<
`<�<�<hj<�#	<��<V�<���;͇�;�7�;���;M��;���;h~�;�s�;w�;���;5��;�ۻ;8�;�k�;(˪;�9�;��;H�;��;���;�T�;�#�;c�;C�u;%�k;�a;I8X;�N;�E;e�;;�Z2;`.); ;�,;"W;��;X��:���:�!�:F��:U�: צ:�ʖ:&�:-zn:�qO:��0:�_:��9�)�9��d9|��8�]h�q��yg�A�æ��u���(�0D��_��y�/4��=i��������\����h˺�8غ���L��C��ai�Q��������F��o$��*��0�;�6��<�}�B�&
I�,O�R"U�.+[�:2a��7g��;m� ?s��Ay��C�䢂�]���z���ܧ��(�������ű��ᶗ�Q����  �  Bh==��='D=T�=?�=�=(� =+X =���<-"�<�Y�<��<��<)��<]0�<�c�<���<���<z��<%�<rR�<�~�<2��<m��<!��<K �<�D�<�g�<��<>��<���<=��<���<D�<�'�<�:�<�K�< Z�<8f�<�o�<�v�<H{�<�|�<�{�<�w�<q�<Og�<`Z�<PJ�<7�<� �<��<���<��<��<7}�<�Q�<�"�<G��<չ�<��<�A�<���<��<qp�<�"�<q��<|�<�"�<���<cd�<R��<_��<�)�<⸻<pD�<6̸<FP�<�е<rM�<�Ʋ<X<�<���<u�< ��<Y�<�V�<���<��<t�<�͢<A$�<`x�<�ɝ<(�<f�<���<��<�?�<��<�Ƒ<��<7G�<��<���<���<�6�<�o�<姃<߁<��<��|< y<�ju<��q<8<n<��j<g<�uc<��_<sH\<�X<�U<��Q<h�M<�jJ<��F<AQC<�?<zA<<��8<�<5<<�1<E.<��*<
\'<z�#<@� <m<O�<�_<�<ζ<Lj<u#	<U�<q�<���;̇�;�7�;���;c��;���;�~�;�s�;>w�;���;!��;�ۻ;�;�k�;˪;5:�;-��;
H�;�;ە�;�T�;g#�;\�;�u;��k;��a;�7X;��N;HE;��;;�Z2;t.);] ;-;YW;�;���:`��:!�:��:��:
ئ:�ʖ:>�:�xn:wqO:�0:�a:���9*�9��d9���8:h��#�{g����[t���(�D�|_��y��4���i��򇤺����p����i˺L9غ��亗��nC��si���a��l��F��o$��*���0���6���<�5�B��	I�kO�~"U��+[�2a�o7g�{;m�?s�wAy��C�
���N�������ǧ��I�����������𶗻#����  �  :h==��=-D=R�==�=�=(� =4X =���<6"�<�Y�<ݐ�<���<#��<W0�<zc�<���<���<���<0%�<sR�<�~�<)��<k��<)��<M �<�D�<�g�<��<2��<���<=��<���<G�<�'�<�:�<�K�<"Z�</f�<�o�<�v�<:{�<�|�<�{�<�w�<q�<Ng�<cZ�<^J�<37�<� �<��<���<��<��<1}�<�Q�<�"�<O��<ٹ�<��<�A�<���<��<jp�<�"�<r��<|�<�"�<}��<Wd�<G��<b��<�)�<<jD�<7̸<RP�<�е<vM�<�Ʋ<L<�<���<n�<��<]�<�V�<���<��<t�<�͢<Q$�<gx�<ʝ<�<�e�<���<��<�?�<��<�Ƒ<��<KG�<��<���<���<�6�<�o�<꧃<߁<x�<��|<� y<�ju<��q<=<n<��j<�g<�uc<��_<sH\<�X<�U<ɋQ<I�M<�jJ<��F<YQC<�?<qA<<��8<�<5<b�1<E.<��*<\'<g�#<6� <a<B�<�_<�<޶<fj<�#	<W�<p�<���;Ƈ�;�7�;���;X��;���;k~�;Vs�;Ew�;���;J��;�ۻ;��;�k�;�ʪ;;:�;��;�G�;��;���;�T�;s#�;~�;��u;��k;�a;�7X;P�N;lE;Ԥ;;TZ2;$.);. ;�,;W;��;A��:���:R"�:
��:��:�צ:rʖ:��:
yn:�qO:T�0:x_:���9;'�9̋d9���8:�f�*츠zg���B���s�`�(��D�	_���y��4��bi��􇤺U���|����i˺"8غ���$���B���i�@�������?G��o$���*�_�0���6���<�?�B��	I��O�""U�m+[�2a��7g��;m�a?s��Ay��C� ��������������9��������������R����  �  >h==��=(D=U�=>�=�=2� =%X =���<0"�<�Y�<��<���<$��<X0�<�c�<���<���<{��<%�<�R�<�~�<4��<j��<%��<Q �<�D�<�g�<��<F��<���<E��<���<@�<�'�<�:�<�K�<Z�<5f�<�o�<�v�<A{�<�|�<�{�<�w�<!q�<Gg�<bZ�<`J�<7�<� �<��<���<��<��<4}�<�Q�<�"�<B��<ݹ�<��<�A�<���<��<vp�<�"�<v��<|�<�"�<���<nd�<R��<U��<�)�<⸻<oD�<4̸<FP�<�е<jM�<�Ʋ<[<�<���<s�<��<]�<�V�<���<��<t�<�͢<B$�<jx�<�ɝ<0�<f�<���<��<�?�<��<�Ƒ<��<.G�<*��<���<���<�6�<�o�<<߁<�<��|< y<�ju<��q<;<n<��j<g<�uc<��_<xH\<�X<�U<܋Q<V�M<�jJ<��F<FQC<�?<uA<<��8<�<5<#�1<E.<��*<\'<��#<6� <d<E�<`<�<�<Oj<d#	<}�<\�<���;�;�7�;���;`��;՗�;�~�;�s�;w�;���;'��;�ۻ;�;�k�; ˪;:�;!��;;H�;��;���;�T�;�#�;T�;V�u;]�k;�a;	8X;��N;~E;o�;;�Z2;�.);@ ; -;?W;+�;t��:���:� �:���:7�:�צ:5˖:��:myn:EqO:d�0:�`:Y��9%*�9��d9	��8�Fh��$�!|g���E��Hu�s�(�D��_�Q�y�q4��Xi��4�����������h˺y9غ������C��5i�,��������F��o$���*�M�0���6�i�<�x�B��	I�;O�g"U�L+[�B2a��7g��;m��>s��Ay��C����L���ǥ��Χ��F�������ñ������-����  �  Ch==��=&D=S�=@�=�=5� ='X =���<,"�<�Y�<��<���</��<N0�<�c�<���<���<���<%�<�R�<|~�<:��<b��<&��<Q �<�D�<�g�<܈�<;��<���<N��<���<G�<�'�<�:�<�K�<Z�<0f�<�o�<�v�<G{�<�|�<�{�<�w�<!q�<Cg�<bZ�<eJ�<!7�<� �<��<���<��<��<9}�<�Q�<�"�<9��<��<��<�A�<���<��<wp�<�"�<���<|�<�"�<���<Xd�<L��<[��<�)�<ܸ�<yD�<;̸<AP�<�е<iM�<�Ʋ<G<�<���<r�<��<b�<�V�<���<��<&t�<�͢<O$�<kx�<�ɝ<3�<�e�<���<��<�?�<��<�Ƒ<��<4G�<2��<���<���<�6�<�o�<���<߁<��<y�|<y<�ju<��q<F<n<��j< g<�uc<��_<�H\<�X<�U<��Q<j�M<�jJ<��F<=QC<	�?<zA<<��8<�<5<.�1<BE.<��*<\'<��#<#� <y<1�<`<�<ݶ<pj<t#	<��<E�<��;���;�7�;���;R��;��;U~�;ys�;w�;ԉ�;��;�ۻ;6�;�k�;0˪;1:�;��;�G�;��;ו�;�T�;�#�;3�;Z�u;:�k;�a;88X;��N;�E;�;;�Z2;9.);J ;/-;�V;S�;���:���:�!�:���:^�:"צ:K˖:r�:�zn:�pO:��0:-`:��9}(�9��d9x��8 i�\�wxg�8򫹢��ru�{�(��D��_�{�y��4��i��Ɉ��6�������Wh˺�8غ���ڤ�D��"i����3�����F��o$��*���0���6�(�<���B��	I�\O��"U�+[�i2a�c7g�<m�?s��Ay��C��X�������ǧ��8���k���ձ��򶗻t����  �  @h==��=+D=R�=<�=�=,� =.X =���<,"�<Z�<��<���<.��<R0�<�c�<���<���<��<$%�<zR�<�~�<4��<i��<*��<J �<�D�<�g�<��<A��<���<8��<���<I�<�'�<�:�<�K�<Z�<5f�<�o�<�v�<D{�<�|�<�{�<�w�<q�<Dg�<^Z�<YJ�<$7�<� �<��<���<��<��<8}�<�Q�<�"�<K��<չ�<��<�A�<���<��<rp�<�"�<w��<|�<�"�<���<dd�<P��<\��<�)�<鸻<iD�<8̸<GP�<�е<pM�<�Ʋ<U<�<���<p�<���<a�<�V�<���<��<t�<�͢<G$�<`x�<ʝ<(�<�e�<���<��<�?�<"��<�Ƒ<��<?G�< ��<���<���<�6�<�o�<맃<߁<��<��|<y<�ju<��q<0<n<��j<�g<�uc<��_<jH\< �X<�U<ϋQ<_�M<�jJ<��F<RQC<�?<nA<<��8<�<5<J�1<E.<��*<#\'<s�#<2� <w<9�<�_<�<ζ<Xj<�#	<e�<V�<���;���;�7�;���;N��;ؗ�;�~�;�s�;?w�;}��;#��;�ۻ;��;�k�;�ʪ;':�; ��;H�;��;̕�;�T�;#�;e�;2�u;I�k;��a;�7X;גN;IE;��;;�Z2;.);X ;"-;�V;2�;��:]��:s!�:{��:��:`צ:�ʖ:A�:�yn:�pO:Q�0:�`:��9~)�9�d9O��8�`g��*��yg�����xt���(��D��_���y��4��i��/�������M���`i˺�8غa�云��B��ui�{��F���� G��o$���*�w�0�H�6���<�[�B��	I�uO�H"U�d+[�X2a��7g��;m��>s�nAy��C���������������S�����������׶��F����  �  :h==��=)D=U�=9�=�=*� =1X =���<2"�<�Y�<��<��<��<g0�<yc�<���<���<~��<'%�<yR�<�~�<+��<q��<%��<M �<�D�<�g�<��<2��<���<:��<���<M�<�'�<�:�<�K�<#Z�<)f�<�o�<�v�<>{�<�|�<�{�<�w�<q�<Ig�<fZ�<ZJ�<-7�<� �<��<���<��<��</}�<�Q�<�"�<O��<ҹ�<��<�A�<���<��<mp�<�"�<o��<|�<�"�<���<cd�<D��<c��<~)�<�<hD�<:̸<JP�<�е<uM�<�Ʋ<Z<�<���<v�<��<[�<�V�<���<��<t�<�͢<J$�<^x�<ʝ<�<f�<���< ��<�?�<��<�Ƒ<��<GG�<��<���<���<�6�<�o�<秃<"߁<y�<��|<� y<�ju<��q<"<n<��j<�g<�uc<��_<tH\<�X<�U<�Q<I�M<�jJ<��F<KQC<�?<`A<<��8<�<5<W�1<E.<��*<\'<p�#<L� <M<c�<�_<�<Ѷ<Vj<�#	<d�<s�<���;އ�;�7�;���;t��;���;�~�;Us�;;w�;���;'��;ܻ;��;�k�;�ʪ;B:�;�;H�;��;���;�T�;e#�;��;#�u;l�k;%�a;�7X;�N;/E;ͤ;;UZ2;�.);H ;�,;vW;��;B��:6��:�!�:���:�:�צ:�ʖ:��:�xn:rO:��0:�`:���9�&�9��d9���82�f��+��xg��﫹ª��s�u�(�3D�=_���y�y4���i������$�������\i˺�8غ:�享���B���i�������D��F�p$���*���0��6���<���B��	I�QO�A"U��+[��1a��7g��;m�,?s��Ay��C�8��������������m��������������"����  �  <h==��=&D=W�=:�=�=/� =-X =���<7"�<�Y�<��<��<��<`0�<�c�<���<���<���<"%�<�R�<�~�</��<n��<!��<N �<�D�<�g�<��<6��<���<L��<���<E�<�'�<�:�<�K�<'Z�<,f�<�o�<�v�<={�<�|�<�{�<�w�<!q�<Cg�<bZ�<^J�<*7�<� �<��<���<��<��<0}�<�Q�<�"�<H��<޹�<��<�A�<���<��<tp�<�"�<v��<|�<�"�<���<\d�<F��<b��<�)�<۸�<rD�<9̸<@P�<�е<oM�<�Ʋ<P<�<���<m�<��<[�<�V�<���<��<t�<�͢<P$�<ix�<�ɝ<!�<f�<���<��<�?�<��<�Ƒ<��<?G�<%��<���<���<�6�<�o�<�<߁<{�<��|<y<�ju<��q<6<n<��j<g<�uc<��_<�H\<�X<�U<ՋQ<N�M<�jJ<��F<?QC<�?<dA<<��8<�<5<E�1<*E.<��*<�['<z�#<C� <N<U�<�_<�<�<hj<~#	<w�<X�<���;҇�;�7�;���;G��;ʗ�;�~�;fs�;#w�;Ή�;
��;�ۻ;�;�k�;˪;N:�;���;�G�;��;���;�T�;�#�;[�;V�u;<�k;�a;�7X;�N;�E;��;;TZ2;b.);A ;�,;KW;ǜ;���:���:�!�:ց�:!�:Yצ:˖:5�:�yn:�pO:��0:N`:��96'�9��d9x��8�%i��!츻yg���]�㹶t��(�jD�7_��y��4���i������͑��I����h˺�8غ������TC���i�������g��F�$p$���*� �0�E�6���<�N�B��	I�*O�z"U�5+[�b2a��7g��;m�?s��Ay�jC����T�������ɧ��Y���Y���ͱ������8����  �  Eh==��=&D=S�=>�=�=2� ='X =���<("�< Z�<��<���<4��<Q0�<�c�<���<���<~��<%�<�R�<�~�<8��<b��<%��<Q �<�D�<�g�<ވ�<N��<���<B��<���<@�<�'�<�:�<�K�<Z�<9f�<�o�<�v�<L{�<�|�<�{�<�w�<$q�<Eg�<dZ�<]J�<7�<� �<��<���<��<��<=}�<�Q�<�"�<E��<ڹ�<��<�A�<���<��<|p�<�"�<|��<|�<�"�<���<_d�<X��<N��<�)�<ݸ�<uD�<6̸<DP�<�е<aM�<�Ʋ<K<�<���<n�<��<`�<�V�<���<��<!t�<�͢<F$�<cx�<ʝ<2�<�e�<���<��<�?�<#��<�Ƒ<��<2G�<)��<���<���<�6�<�o�<���<
߁<��<�|<y<�ju<��q<L<n<��j<g<�uc<��_<fH\<�X<�U<��Q<u�M<�jJ<��F<=QC<�?<sA<<��8<�<5<-�1<E.<��*<\'<��#<4� <�<6�<`<�<Ѷ<Vj<m#	<��<T�<	��;���;�7�;���;5��;��;^~�;�s�;w�;���;&��;�ۻ;&�;�k�;-˪;�9�;3��;H�;��;앏;vT�;�#�;1�;p�u;Q�k;�a;�7X;��N;kE;j�;;�Z2;.);r ;H-;�V;o�;���:���:"!�:���:B�:cצ:�˖:l�:0zn:0pO:�0:a:���9�+�9�d9���8��h���!{g�g�ڧ�^v�W�(�D��_��y��4��-i���������V����h˺X9غv��\��C��&i�r�������F��o$��*�R�0���6�q�<�L�B��	I�]O��"U�+[��2a�;7g�<m��>s��Ay�'D�䢂�g�������⧋�.���������������p����  �  Bh==��=(D=U�=<�=�=-� =0X =���<."�<�Y�<��<���<%��<V0�<�c�<���<���<���<(%�<~R�<�~�<1��<j��<)��<S �<�D�<�g�<و�<<��<���<?��<���<E�<�'�<�:�<�K�<Z�<5f�<�o�<�v�<E{�<�|�<�{�<�w�<q�<Gg�<eZ�<]J�<17�<� �<��<���<	��<��<4}�<�Q�<�"�<@��<��<��<�A�<���<��<sp�<�"�<y��<|�<�"�<���<Vd�<O��<W��<�)�<渻<nD�<7̸<NP�<�е<jM�<�Ʋ<E<�<���<o�<��<a�<�V�<���<��<t�<�͢<X$�<hx�<�ɝ<(�<�e�<���<��<�?�<��<�Ƒ<��<EG�<$��<���<���<�6�<�o�<�<߁<��<p�|<� y<�ju<��q<L<n<��j< g<�uc<��_<kH\<�X<�U<��Q<g�M<�jJ<��F<HQC<�?<mA<<��8<�<5<Q�1<;E.<��*<\'<�#<,� <g<A�<�_<�<ٶ<vj<�#	<m�<_�<���;Ň�;�7�;���;>��;��;I~�;s�;w�;���;J��;�ۻ; �;�k�;!˪;:�;!��;�G�;��;Е�;�T�;�#�;V�;<�u;a�k;�a;�7X;?�N;�E;m�;;�Z2;N.);5 ;-;W;
�;V��: ��:z"�:́�:8�:�צ: ˖:��:�yn:%qO:}�0:M`:Y��9>)�9D�d9���83�g�&츁zg�﫹���Su�9�(��D�W_���y�s4��i��/���������� i˺�8غU����C��wi�=��z�����F��o$���*��0��6���<�(�B��	I�QO�j"U�5+[�V2a�w7g�@<m�5?s��Ay��C�䢂�?���˥������$��������������������  �  8h==��=&D=Y�=:�=�=*� =+X =���<6"�<�Y�<��<��<��<b0�<�c�<���<���<v��< %�<vR�<�~�<,��<s��<��<U �<�D�<�g�<���<9��<���<>��<���<D�<�'�<�:�<�K�<#Z�<1f�<�o�<�v�<8{�<�|�<�{�<�w�<q�<Fg�<^Z�<SJ�< 7�<� �<��<���<��<��<1}�<�Q�<�"�<N��<Թ�<��<�A�<���<��<op�<�"�<m��<|�<�"�<���<id�<J��<d��<~)�<฻<kD�<5̸<@P�<�е<vM�<�Ʋ<_<�<���<r�<	��<T�<�V�<���<��<t�<�͢<?$�<ex�<ʝ<$�<
f�<���<��<�?�<��<�Ƒ<��<8G�<��<���<���<�6�<�o�<駃< ߁<t�<��|<y<�ju<��q<"<n<��j<�g<�uc<��_<~H\<�X<�U<�Q<A�M<�jJ<��F<>QC< �?<eA<<��8<�<5<<�1<E.<��*<\'<��#<A� <N<Y�<�_<�<ݶ<Ej<x#	<^�<l�<���;��;n7�;���;S��;���;�~�;ss�;Ew�;���;���;�ۻ;��;�k�;�ʪ;@:�;��;#H�;	�;���;�T�;\#�;n�;(�u;T�k;��a;�7X;��N;6E;Ϥ;;kZ2;�.);; ;�,;xW;ٜ;+��:M��:!�:��:��:�צ:�ʖ:��:`xn:"rO:��0:�a:I��90(�9͌d9$��8sh�)츋{g��򫹕���s���(��
D�_���y�%4���i���������������i˺G9غ���8��C���i������z��F��o$���*���0�{�6���<�$�B��	I�&O�k"U�x+[�2a�8g�Z;m��>s��Ay��C�7���G���ѥ������x���z�������궗�����  �  8h==��=(D=S�=9�=�=2� =0X =���<7"�<�Y�<��<���<)��<U0�<�c�<���<���<��<.%�<�R�<�~�<'��<h��<"��<W �<�D�<�g�<���<4��<���<C��<���<I�<�'�<�:�<�K�<Z�<+f�<�o�<�v�<6{�<�|�<�{�<�w�<q�<Eg�<gZ�<gJ�<+7�<� �<��<���<	��<��<5}�<�Q�<�"�<K��<߹�<��<�A�<���<��<np�<�"�<u��<|�<�"�<{��<Ud�<F��<\��<�)�<븻<rD�<:̸<IP�<�е<mM�<�Ʋ<I<�<���<p�<��<Y�<�V�<���<��<!t�<�͢<J$�<lx�<ʝ<'�<�e�<���<��<�?�<��<�Ƒ<��<DG�<.��<���<���<�6�<�o�<�< ߁<s�<��|<� y<�ju<��q<7<n<��j<	g<�uc<��_<rH\<�X<�U<ǋQ<?�M<�jJ<��F<EQC<	�?<^A<<��8<�<5<S�1<E.<��*<\'<}�#<2� <n<>�<�_<�<�<Xj<�#	<��<i�<���;���;�7�;���;U��;���;g~�;]s�;&w�;���;&��;�ۻ;�;�k�;˪;#:�;���;�G�;��;���;�T�;�#�;j�;�u;Q�k;-�a;I8X;�N;�E;��;;uZ2;H.);: ;	-;W;��;���:	��:�!�:U��:h�:�צ:�ʖ:T�:cyn:/rO::�0:0_:A��9'�9݈d9���8`g�"�yg�𫹐���t��(�JD�l	_���y��3���i��1���-���ʆ���h˺F8غ,��Ԥ�C��~i�A��S�����F��o$���*�E�0��6�N�<��B��	I�vO�Y"U�9+[�2a�8g��;m�D?s��Ay��C����.�����������R�������ű�����T����  �  Fh==��=)D=T�=@�=�=+� =+X =���<."�<�Y�<��<���<8��<Q0�<�c�<���<���<���<%�<zR�<�~�<5��<m��<*��<E �<�D�<�g�<��<H��<���<>��<���<@�<�'�<�:�<�K�<Z�<@f�<�o�<�v�<H{�<�|�<�{�<�w�< q�<Lg�<_Z�<UJ�<7�<� �<��<���<��<��<;}�<�Q�<�"�<;��<߹�<��<�A�<���<��<wp�<�"�<s��<|�<�"�<���<ed�<[��<U��<�)�<⸻<hD�<1̸<IP�<�е<iM�<�Ʋ<S<�<���<p�<���<_�<�V�<���<��<t�<�͢<J$�<fx�<�ɝ<1�<�e�<���<��<�?�<��<�Ƒ<��<8G�<��<���<���<�6�<�o�<姃<߁<��<��|<y<�ju<��q<G<n<��j<�g<�uc<��_<hH\<�X<�U<ӋQ<v�M<�jJ<��F<KQC<�?<{A<<��8<�<5<>�1<(E.<��*<\'<��#<(� <�<7�<`<�<ֶ<]j<v#	<e�<`�<���;χ�;�7�;x��;:��;��;�~�;�s�;w�;���;1��;�ۻ;��;�k�;˪;:�;O��;H�;��;ܕ�;�T�;l#�;X�;S�u;��k;��a;�7X;��N;�E;G�;;�Z2;_.);V ;;-;W;[�;
��:��:g!�:F��:��:�צ:M˖: �: yn:NpO:ο0:�a:N��9�,�9��d9!��8�0h�Q,�J}g�J�&��tu���(�D�R_���y��4��Ai������T������ki˺Q9غ*��,���C��-i�c�� �����F��o$���*��0���6���<�I�B��	I�YO�V"U��+[�h2a�O7g��;m��>s�LAy��C�좂�I���䥈�ç��2�����������ɶ��?����  �  8h==��=(D=S�=9�=�=2� =0X =���<7"�<�Y�<��<���<)��<U0�<�c�<���<���<��<.%�<�R�<�~�<'��<h��<"��<W �<�D�<�g�<���<4��<���<C��<���<I�<�'�<�:�<�K�<Z�<+f�<�o�<�v�<6{�<�|�<�{�<�w�<q�<Eg�<gZ�<gJ�<+7�<� �<��<���<	��<��<5}�<�Q�<�"�<K��<߹�<��<�A�<���<��<np�<�"�<u��<|�<�"�<{��<Ud�<F��<\��<�)�<븻<rD�<:̸<IP�<�е<mM�<�Ʋ<I<�<���<p�<��<Y�<�V�<���<��<!t�<�͢<J$�<lx�<ʝ<'�<�e�<���<��<�?�<��<�Ƒ<��<DG�<.��<���<���<�6�<�o�<�< ߁<s�<��|<� y<�ju<��q<7<n<��j<	g<�uc<��_<rH\<�X<�U<ǋQ<?�M<�jJ<��F<EQC<	�?<^A<<��8<�<5<S�1<E.<��*<\'<}�#<2� <n<>�<�_<�<�<Xj<�#	<��<i�<���;���;�7�;���;U��;���;g~�;]s�;&w�;���;&��;�ۻ;�;�k�;˪;#:�;���;�G�;��;���;�T�;�#�;j�;�u;Q�k;-�a;I8X;�N;�E;��;;uZ2;H.);: ;	-;W;��;���:	��:�!�:U��:h�:�צ:�ʖ:T�:cyn:/rO::�0:0_:A��9'�9݈d9���8`g�"�yg�𫹐���t��(�JD�l	_���y��3���i��1���-���ʆ���h˺F8غ,��Ԥ�C��~i�A��S�����F��o$���*�E�0��6�N�<��B��	I�vO�Y"U�9+[�2a�8g��;m�D?s��Ay��C����.�����������R�������ű�����T����  �  8h==��=&D=Y�=:�=�=*� =+X =���<6"�<�Y�<��<��<��<b0�<�c�<���<���<v��< %�<vR�<�~�<,��<s��<��<U �<�D�<�g�<���<9��<���<>��<���<D�<�'�<�:�<�K�<#Z�<1f�<�o�<�v�<8{�<�|�<�{�<�w�<q�<Fg�<^Z�<SJ�< 7�<� �<��<���<��<��<1}�<�Q�<�"�<N��<Թ�<��<�A�<���<��<op�<�"�<m��<|�<�"�<���<id�<J��<d��<~)�<฻<kD�<5̸<@P�<�е<vM�<�Ʋ<_<�<���<r�<	��<T�<�V�<���<��<t�<�͢<?$�<ex�<ʝ<$�<
f�<���<��<�?�<��<�Ƒ<��<8G�<��<���<���<�6�<�o�<駃< ߁<t�<��|<y<�ju<��q<"<n<��j<�g<�uc<��_<~H\<�X<�U<�Q<A�M<�jJ<��F<>QC< �?<eA<<��8<�<5<<�1<E.<��*<\'<��#<A� <N<Y�<�_<�<ݶ<Ej<x#	<^�<l�<���;��;n7�;���;S��;���;�~�;ss�;Ew�;���;���;�ۻ;��;�k�;�ʪ;@:�;��;#H�;	�;���;�T�;\#�;n�;(�u;T�k;��a;�7X;��N;6E;Ϥ;;kZ2;�.);; ;�,;xW;ٜ;+��:M��:!�:��:��:�צ:�ʖ:��:`xn:"rO:��0:�a:I��90(�9͌d9$��8sh�)츋{g��򫹕���s���(��
D�_���y�%4���i���������������i˺G9غ���8��C���i������z��F��o$���*���0�{�6���<�$�B��	I�&O�k"U�x+[�2a�8g�Z;m��>s��Ay��C�7���G���ѥ������x���z�������궗�����  �  Bh==��=(D=U�=<�=�=-� =0X =���<."�<�Y�<��<���<%��<V0�<�c�<���<���<���<(%�<~R�<�~�<1��<j��<)��<S �<�D�<�g�<و�<<��<���<?��<���<E�<�'�<�:�<�K�<Z�<5f�<�o�<�v�<E{�<�|�<�{�<�w�<q�<Gg�<eZ�<]J�<17�<� �<��<���<	��<��<4}�<�Q�<�"�<@��<��<��<�A�<���<��<sp�<�"�<y��<|�<�"�<���<Vd�<O��<W��<�)�<渻<nD�<7̸<NP�<�е<jM�<�Ʋ<E<�<���<o�<��<a�<�V�<���<��<t�<�͢<X$�<hx�<�ɝ<(�<�e�<���<��<�?�<��<�Ƒ<��<EG�<$��<���<���<�6�<�o�<�<߁<��<p�|<� y<�ju<��q<L<n<��j< g<�uc<��_<kH\<�X<�U<��Q<g�M<�jJ<��F<HQC<�?<mA<<��8<�<5<Q�1<;E.<��*<\'<�#<,� <g<A�<�_<�<ٶ<vj<�#	<m�<_�<���;Ň�;�7�;���;>��;��;I~�;s�;w�;���;J��;�ۻ; �;�k�;!˪;:�;!��;�G�;��;Е�;�T�;�#�;V�;<�u;a�k;�a;�7X;?�N;�E;m�;;�Z2;N.);5 ;-;W;
�;V��: ��:z"�:́�:8�:�צ: ˖:��:�yn:%qO:}�0:M`:Y��9>)�9D�d9���84�g�&츁zg�﫹���Su�9�(��D�W_���y�s4��i��/���������� i˺�8غU����C��wi�=��z�����F��o$���*��0��6���<�(�B��	I�QO�j"U�5+[�V2a�w7g�@<m�5?s��Ay��C�䢂�?���˥������$��������������������  �  Eh==��=&D=S�=>�=�=2� ='X =���<("�< Z�<��<���<4��<Q0�<�c�<���<���<~��<%�<�R�<�~�<8��<b��<%��<Q �<�D�<�g�<ވ�<N��<���<B��<���<@�<�'�<�:�<�K�<Z�<9f�<�o�<�v�<L{�<�|�<�{�<�w�<$q�<Eg�<dZ�<]J�<7�<� �<��<���<��<��<=}�<�Q�<�"�<E��<ڹ�<��<�A�<���<��<|p�<�"�<|��<|�<�"�<���<_d�<X��<N��<�)�<ݸ�<uD�<6̸<DP�<�е<aM�<�Ʋ<K<�<���<n�<��<`�<�V�<���<��<!t�<�͢<F$�<cx�<ʝ<2�<�e�<���<��<�?�<#��<�Ƒ<��<2G�<)��<���<���<�6�<�o�<���<
߁<��<�|<y<�ju<��q<L<n<��j<g<�uc<��_<fH\<�X<�U<��Q<u�M<�jJ<��F<=QC<�?<sA<<��8<�<5<-�1<E.<��*<\'<��#<4� <�<6�<`<�<Ѷ<Vj<m#	<��<T�<	��;���;�7�;���;5��;��;^~�;�s�;w�;���;&��;�ۻ;&�;�k�;-˪;�9�;3��;H�;��;앏;vT�;�#�;1�;p�u;Q�k;�a;�7X;��N;kE;j�;;�Z2;.);r ;H-;�V;o�;���:���:"!�:���:B�:cצ:�˖:l�:0zn:0pO:�0:a:���9�+�9�d9���8��h���!{g�g�ڧ�^v�W�(�D��_��y��4��-i���������V����h˺X9غv��\��C��&i�r�������F��o$��*�R�0���6�q�<�L�B��	I�]O��"U�+[��2a�;7g�<m��>s��Ay�'D�䢂�g�������⧋�.���������������p����  �  <h==��=&D=W�=:�=�=/� =-X =���<7"�<�Y�<��<��<��<`0�<�c�<���<���<���<"%�<�R�<�~�</��<n��<!��<N �<�D�<�g�<��<6��<���<L��<���<E�<�'�<�:�<�K�<'Z�<,f�<�o�<�v�<={�<�|�<�{�<�w�<!q�<Cg�<bZ�<^J�<*7�<� �<��<���<��<��<0}�<�Q�<�"�<H��<޹�<��<�A�<���<��<tp�<�"�<v��<|�<�"�<���<\d�<F��<b��<�)�<۸�<rD�<9̸<@P�<�е<oM�<�Ʋ<P<�<���<m�<��<[�<�V�<���<��<t�<�͢<P$�<ix�<�ɝ<!�<f�<���<��<�?�<��<�Ƒ<��<?G�<%��<���<���<�6�<�o�<�<߁<{�<��|<y<�ju<��q<6<n<��j<g<�uc<��_<�H\<�X<�U<ՋQ<N�M<�jJ<��F<?QC<�?<dA<<��8<�<5<E�1<*E.<��*<�['<z�#<C� <N<U�<�_<�<�<hj<~#	<w�<X�<���;҇�;�7�;���;G��;ʗ�;�~�;fs�;#w�;Ή�;
��;�ۻ;�;�k�;˪;N:�;���;�G�;��;���;�T�;�#�;[�;V�u;<�k;�a;�7X;�N;�E;��;;TZ2;b.);A ;�,;KW;ǜ;���:���:�!�:ց�:!�:Yצ:˖:5�:�yn:�pO:��0:N`:��96'�9��d9x��8�%i��!츻yg���]�㹶t��(�jD�7_��y��4���i������͑��I����h˺�8غ������TC���i�������g��F�$p$���*� �0�E�6���<�N�B��	I�*O�z"U�5+[�b2a��7g��;m�?s��Ay�jC����T�������ɧ��Y���Y���ͱ������8����  �  :h==��=)D=U�=9�=�=*� =1X =���<2"�<�Y�<��<��<��<g0�<yc�<���<���<~��<'%�<yR�<�~�<+��<q��<%��<M �<�D�<�g�<��<2��<���<:��<���<M�<�'�<�:�<�K�<#Z�<)f�<�o�<�v�<>{�<�|�<�{�<�w�<q�<Ig�<fZ�<ZJ�<-7�<� �<��<���<��<��</}�<�Q�<�"�<O��<ҹ�<��<�A�<���<��<mp�<�"�<o��<|�<�"�<���<cd�<D��<c��<~)�<�<hD�<:̸<JP�<�е<uM�<�Ʋ<Z<�<���<v�<��<[�<�V�<���<��<t�<�͢<J$�<^x�<ʝ<�<f�<���< ��<�?�<��<�Ƒ<��<GG�<��<���<���<�6�<�o�<秃<"߁<y�<��|<� y<�ju<��q<"<n<��j<�g<�uc<��_<tH\<�X<�U<�Q<I�M<�jJ<��F<KQC<�?<`A<<��8<�<5<W�1<E.<��*<\'<p�#<L� <M<c�<�_<�<Ѷ<Vj<�#	<d�<s�<���;އ�;�7�;���;t��;���;�~�;Us�;;w�;���;'��;ܻ;��;�k�;�ʪ;B:�;�;H�;��;���;�T�;e#�;��;#�u;l�k;%�a;�7X;�N;/E;ͤ;;UZ2;�.);H ;�,;vW;��;B��:6��:�!�:���:�:�צ:�ʖ:��:�xn:rO:��0:�`:���9�&�9��d9���82�f��+��xg��﫹ª��s�u�(�3D�=_���y�y4���i������$�������\i˺�8غ:�享���B���i�������D��F�p$���*���0��6���<���B��	I�QO�A"U��+[��1a��7g��;m�,?s��Ay��C�8��������������m��������������"����  �  @h==��=+D=R�=<�=�=,� =.X =���<,"�<Z�<��<���<.��<R0�<�c�<���<���<��<$%�<zR�<�~�<4��<i��<*��<J �<�D�<�g�<��<A��<���<8��<���<I�<�'�<�:�<�K�<Z�<5f�<�o�<�v�<D{�<�|�<�{�<�w�<q�<Dg�<^Z�<YJ�<$7�<� �<��<���<��<��<8}�<�Q�<�"�<K��<չ�<��<�A�<���<��<rp�<�"�<w��<|�<�"�<���<dd�<P��<\��<�)�<鸻<iD�<8̸<GP�<�е<pM�<�Ʋ<U<�<���<p�<���<a�<�V�<���<��<t�<�͢<G$�<`x�<ʝ<(�<�e�<���<��<�?�<"��<�Ƒ<��<?G�< ��<���<���<�6�<�o�<맃<߁<��<��|<y<�ju<��q<0<n<��j<�g<�uc<��_<jH\< �X<�U<ϋQ<_�M<�jJ<��F<RQC<�?<nA<<��8<�<5<J�1<E.<��*<#\'<s�#<2� <w<9�<�_<�<ζ<Xj<�#	<e�<V�<���;���;�7�;���;N��;ؗ�;�~�;�s�;?w�;}��;#��;�ۻ;��;�k�;�ʪ;':�; ��;H�;��;̕�;�T�;#�;e�;2�u;I�k;��a;�7X;גN;IE;��;;�Z2;.);X ;"-;�V;2�;��:]��:s!�:{��:��:`צ:�ʖ:A�:�yn:�pO:Q�0:�`:��9~)�9�d9O��8�`g��*��yg�����xt���(��D��_���y��4��i��/�������M���`i˺�8غa�云��B��ui�{��F���� G��o$���*�w�0�H�6���<�[�B��	I�uO�H"U�d+[�X2a��7g��;m��>s�nAy��C���������������S�����������׶��F����  �  Ch==��=&D=S�=@�=�=5� ='X =���<,"�<�Y�<��<���</��<N0�<�c�<���<���<���<%�<�R�<|~�<:��<b��<&��<Q �<�D�<�g�<܈�<;��<���<N��<���<G�<�'�<�:�<�K�<Z�<0f�<�o�<�v�<G{�<�|�<�{�<�w�<!q�<Cg�<bZ�<eJ�<!7�<� �<��<���<��<��<9}�<�Q�<�"�<9��<��<��<�A�<���<��<wp�<�"�<���<|�<�"�<���<Xd�<L��<[��<�)�<ܸ�<yD�<;̸<AP�<�е<iM�<�Ʋ<G<�<���<r�<��<b�<�V�<���<��<&t�<�͢<O$�<kx�<�ɝ<3�<�e�<���<��<�?�<��<�Ƒ<��<4G�<2��<���<���<�6�<�o�<���<߁<��<y�|<y<�ju<��q<F<n<��j< g<�uc<��_<�H\<�X<�U<��Q<j�M<�jJ<��F<=QC<	�?<zA<<��8<�<5<.�1<BE.<��*<\'<��#<#� <y<1�<`<�<ݶ<pj<t#	<��<E�<��;���;�7�;���;R��;��;U~�;ys�;w�;ԉ�;��;�ۻ;6�;�k�;0˪;1:�;��;�G�;��;ו�;�T�;�#�;3�;Z�u;:�k;�a;88X;��N;�E;�;;�Z2;9.);J ;/-;�V;S�;���:���:�!�:���:^�:"צ:K˖:r�:�zn:�pO:��0:-`:��9}(�9��d9x��8 i�\�wxg�8򫹢��ru�{�(��D��_�{�y��4��i��Ɉ��6�������Wh˺�8غ���ڤ�D��"i����3�����F��o$��*���0���6�(�<���B��	I�\O��"U�+[�i2a�c7g�<m�?s��Ay��C��X�������ǧ��8���k���ձ��򶗻t����  �  >h==��=(D=U�=>�=�=2� =%X =���<0"�<�Y�<��<���<$��<X0�<�c�<���<���<{��<%�<�R�<�~�<4��<j��<%��<Q �<�D�<�g�<��<F��<���<E��<���<@�<�'�<�:�<�K�<Z�<5f�<�o�<�v�<A{�<�|�<�{�<�w�<!q�<Gg�<bZ�<`J�<7�<� �<��<���<��<��<4}�<�Q�<�"�<B��<ݹ�<��<�A�<���<��<vp�<�"�<v��<|�<�"�<���<nd�<R��<U��<�)�<⸻<oD�<4̸<FP�<�е<jM�<�Ʋ<[<�<���<s�<��<]�<�V�<���<��<t�<�͢<B$�<jx�<�ɝ<0�<f�<���<��<�?�<��<�Ƒ<��<.G�<*��<���<���<�6�<�o�<<߁<�<��|< y<�ju<��q<;<n<��j<g<�uc<��_<xH\<�X<�U<܋Q<V�M<�jJ<��F<FQC<�?<uA<<��8<�<5<#�1<E.<��*<\'<��#<6� <d<E�<`<�<�<Oj<d#	<}�<\�<���;�;�7�;���;`��;՗�;�~�;�s�;w�;���;'��;�ۻ;�;�k�; ˪;:�;!��;;H�;��;���;�T�;�#�;T�;V�u;]�k;�a;	8X;��N;~E;o�;;�Z2;�.);@ ; -;?W;+�;t��:���:� �:���:7�:�צ:5˖:��:myn:EqO:d�0:�`:Y��9%*�9��d9	��8�Fh��$�!|g���E��Hu�s�(�D��_�Q�y�q4��Xi��4�����������h˺y9غ������C��5i�,��������F��o$���*�M�0���6�i�<�x�B��	I�;O�g"U�L+[�B2a��7g��;m��>s��Ay��C����L���ǥ��Χ��F�������ñ������-����  �  :h==��=-D=R�==�=�=(� =4X =���<6"�<�Y�<ݐ�<���<#��<W0�<zc�<���<���<���<0%�<sR�<�~�<)��<k��<)��<M �<�D�<�g�<��<2��<���<=��<���<G�<�'�<�:�<�K�<"Z�</f�<�o�<�v�<:{�<�|�<�{�<�w�<q�<Ng�<cZ�<^J�<37�<� �<��<���<��<��<1}�<�Q�<�"�<O��<ٹ�<��<�A�<���<��<jp�<�"�<r��<|�<�"�<}��<Wd�<G��<b��<�)�<<jD�<7̸<RP�<�е<vM�<�Ʋ<L<�<���<n�<��<]�<�V�<���<��<t�<�͢<Q$�<gx�<ʝ<�<�e�<���<��<�?�<��<�Ƒ<��<KG�<��<���<���<�6�<�o�<꧃<߁<x�<��|<� y<�ju<��q<=<n<��j<�g<�uc<��_<sH\<�X<�U<ɋQ<I�M<�jJ<��F<YQC<�?<qA<<��8<�<5<b�1<E.<��*<\'<g�#<6� <a<B�<�_<�<޶<fj<�#	<W�<p�<���;Ƈ�;�7�;���;X��;���;k~�;Vs�;Ew�;���;J��;�ۻ;��;�k�;�ʪ;;:�;��;�G�;��;���;�T�;s#�;~�;��u;��k;�a;�7X;P�N;lE;Ԥ;;TZ2;$.);. ;�,;W;��;A��:���:R"�:
��:��:�צ:rʖ:��:
yn:�qO:T�0:x_:���9;'�9̋d9���8:�f�*츠zg���B���s�`�(��D�	_���y��4��bi��􇤺U���|����i˺"8غ���$���B���i�@�������?G��o$���*�_�0���6���<�?�B��	I��O�""U�m+[�2a��7g��;m�a?s��Ay��C� ��������������9��������������R����  �  Bh==��='D=T�=?�=�=(� =+X =���<-"�<�Y�<��<��<)��<]0�<�c�<���<���<z��<%�<rR�<�~�<2��<m��<!��<K �<�D�<�g�<��<>��<���<=��<���<D�<�'�<�:�<�K�< Z�<8f�<�o�<�v�<H{�<�|�<�{�<�w�<q�<Og�<`Z�<PJ�<7�<� �<��<���<��<��<7}�<�Q�<�"�<G��<չ�<��<�A�<���<��<qp�<�"�<q��<|�<�"�<���<cd�<R��<_��<�)�<⸻<pD�<6̸<FP�<�е<rM�<�Ʋ<X<�<���<u�< ��<Y�<�V�<���<��<t�<�͢<A$�<`x�<�ɝ<(�<f�<���<��<�?�<��<�Ƒ<��<7G�<��<���<���<�6�<�o�<姃<߁<��<��|< y<�ju<��q<8<n<��j<g<�uc<��_<sH\<�X<�U<��Q<h�M<�jJ<��F<AQC<�?<zA<<��8<�<5<<�1<E.<��*<
\'<z�#<@� <m<O�<�_<�<ζ<Lj<u#	<U�<q�<���;̇�;�7�;���;c��;���;�~�;�s�;>w�;���;!��;�ۻ;�;�k�;˪;5:�;-��;
H�;�;ە�;�T�;g#�;\�;�u;��k;��a;�7X;��N;HE;��;;�Z2;t.);] ;-;YW;�;���:`��:!�:��:��:
ئ:�ʖ:>�:�xn:wqO:�0:�a:���9*�9��d9���8:h��#�{g����[t���(�D�|_��y��4���i��򇤺����p����i˺L9غ��亗��nC��si���a��l��F��o$��*���0���6���<�5�B��	I�kO�~"U��+[�2a�o7g�{;m�?s�wAy��C�
���N�������ǧ��I�����������𶗻#����  �  �h=�=��=E=l�=r�=-=�� =�Y =��<�%�<�]�<3��<|��<� �<p5�<�h�<a��<���<���<�+�<�Y�<օ�<��<s��<��<)�<�M�<Fq�<���<���<`��<\��<S�<)�<�3�<vG�<�X�<�g�<<t�<=~�<���<���<���<��<{��<��<�x�<%l�<�\�<�I�<�3�<�<O��<��<'��<���<�f�<8�<��<q��<v��<�W�<��<?��<ǆ�<B9�<���<���<)9�<���<�z�<~�<U��<q?�<�λ<�Y�<f�<3e�<K�<�a�<�ڲ<�O�<���< 0�<L��<-�<�g�<�ɧ<(�<䃤<�ܢ<�2�<~��<�ם<&�<Qr�<S��<)�<J�<���<Б<w�<0O�<|��<PȊ<��<Z<�<�t�<��<��<M�<Ś|<y<blu<�q<o;n<\�j<�	g<�pc<��_<A\<]�X<�U<l�Q<��M<�\J<��F<�@C<T�?<d.<<7�8<C'5<`�1<-.<E�*<zA'<��#<f </�<Ӝ<{?<�<�<�F<|�<w�<;�<���;�5�;���;H��;h�;?�;$�;�;&�;�+�;L�;�{�;��;�	�;�h�;	פ;�U�;^�;�;�1�;���;��;�=;�u;kk;}8a;vW;��M;5ND;��:;��1;�v(;�i;Wz;�;��;\��:��:���:KB�:z۵:T��:͠�:BɅ:9Bl:�GM:�.:�S:��9�L�9� ]9%G�8��*�#����n��!���湸��OK*��pE�2^`��{��Ҋ�[��������Q����˺5�غ�l庾򺘮��e��������D�p��$��*���0���6��=��C��#I�[/O��8U�?[��Da��Gg��Jm�?Ks�Ly��L�A���অ�T�������ܩ��p�������˳�������  �  �h=�=��=E=j�=t�=7=�� =�Y =��<�%�<�]�<*��<���< �<{5�<�h�<d��<���<���<�+�<�Y�<��<��<w��<��<)�<N�<Eq�<В�<���<d��<S��<I�<,�<�3�<xG�<�X�<�g�<5t�<A~�<���<���<���< ��<���<��<�x�<0l�<�\�<�I�<�3�<)�<K��< ��<5��<ϑ�<�f�<8�<��<k��<w��<�W�<��<N��<ņ�<H9�<���<��<'9�<���<�z�<x�<^��<b?�<�λ<�Y�<f�<,e�<?�<�a�<�ڲ<�O�<���<#0�<F��<#�<�g�<�ɧ<*(�<⃤<�ܢ<�2�<{��<�ם<&�<Wr�<\��<:�<J�<���<Б<l�<6O�<{��<cȊ<��<W<�<�t�<	��<��<K�<�|<y<_lu<	�q<P;n<j�j<�	g<�pc<��_<A\<]�X<�U<��Q<��M<�\J<��F<�@C<K�?<j.<<a�8<A'5<j�1<-.<R�*<}A'<��#<<f <?�<�<j?<#�<�<vF<�<p�<c�<��;�5�;���;-��;h�;?�;Q$�;��;4�;u+�;�K�;�{�;��;�	�;�h�;%פ;�U�;m�;!��;�1�;���;޿�;>;�u;�k;�8a;�uW;��M;�MD;N�:;f�1;�v(;Vj;�z;��;K�;��:���:���:B�:�۵:A��:���:�Ʌ:�@l:�GM:��.:�T:��9FK�9+]9e8�8��*������n��#��k�����L*�6oE��]`�>{��Ҋ� ��W�����.����˺H�غ�l���X���������c�D�Np���$���*���0���6��=�2C��#I�z/O��8U�q?[�mDa�Hg�Jm�YKs�%Ly��L����Ŧ��M���e������s�������ݳ��G����  �  �h=�=��="E=k�=m�=4=�� =�Y =��<�%�<�]�<(��<���<� �<}5�<�h�<j��<���<���<�+�<}Y�<��<ذ�<��<��<)�<N�<@q�<Ԓ�<~��<l��<Y��<M�<3�<�3�<�G�<�X�<�g�</t�<=~�<���<���<���<���<���<��<�x�<(l�<�\�<�I�<�3�</�<M��<��<.��<Ƒ�<�f�<8�<��<f��<~��<�W�<��<F��<���<U9�<���<���<,9�<���<�z�<p�<m��<c?�<�λ<�Y�<g�<3e�<C�<�a�<ڲ<�O�<���<.0�<L��<&�<�g�<xɧ<&(�<ۃ�<�ܢ<�2�<z��<�ם<&�<Yr�<L��<7�<	J�<���<Б<i�<DO�<t��<\Ȋ<��<W<�<�t�<��<��<H�<�|<�y<^lu<�q<N;n<��j<s	g<�pc<��_<A\<a�X<�U<��Q<��M<�\J<��F<�@C<N�?<O.<<V�8<0'5<��1<-.<W�*<�A'<��#<:f <�<�<k?</�<�<qF<��<_�<[�<���;�5�;���;2��;Ph�;?�;`$�;��;V�;�+�;L�;�{�;躵;
�;�h�;aפ;�U�;]�;+��;�1�;�;ֿ�;x>;Uu;|k;�8a;�uW;��M;�MD;~�:;v�1;�v(;j;z;��;K�;5��:f��:��:B�:l۵:���:��:oʅ:�@l:�HM:S�.:�T:��97I�9�]9L9�8V�*�]���=n��!����湢���M*��nE�l^`��{�~Ҋ����������r���˺߳غ�l��� �����������4D�^p�ؖ$�|�*��0�[�6�=�fC�-$I�x/O�<8U��?[�Da�%Hg��Im��Ks�)Ly�QL���������}���9������Q����������:����  �  �h=�=��=E=k�=s�=3=�� =�Y =��<�%�<�]�<0��<���<� �<|5�<�h�<`��<���<���<�+�<�Y�<��<��<u��<��<)�<N�<Bq�<Β�<���<i��<V��<C�<0�<�3�<{G�<�X�<�g�<9t�<>~�<���<���<���<��<��<��<�x�<(l�<�\�<�I�<�3�<#�<N��<��</��<ˑ�<�f�<8�<��<r��<p��<�W�<��<G��<ǆ�<H9�<���<��<+9�<���<�z�<z�<`��<a?�<�λ<�Y�<g�<*e�<@�<�a�<�ڲ<�O�<���<%0�<B��<%�<�g�<�ɧ<#(�<���<�ܢ<�2�<���<�ם<&�<Zr�<Y��<5�<J�<���<	Б<t�<2O�<z��<\Ȋ<��<Y<�<�t�<��<��<O�<ښ|<y<jlu<�q<K;n<q�j<u	g<�pc<��_<
A\<h�X<�U<~�Q<��M<�\J<��F<�@C<L�?<g.<<S�8<?'5<g�1<-.<D�*<vA'<��#<9f <;�<�<u?<�<�<sF<��<m�<T�<��;�5�;���;��;%h�;?�;H$�;��;I�;�+�;�K�;�{�;���;�	�;�h�;-פ;�U�;`�;	��;�1�;���;ῄ;>;�u;�k;�8a;�uW;��M;!ND;�:;��1;�v(;%j;�z;��;y�;y��:&��:A��:�A�:s۵:֥�:ʠ�:�Ʌ:Al:�GM:L�.:�S:R��9�K�9]9i7�8��*�q���Vn�$��N�湢��,L*�YoE��^`��{�*ӊ����o����������˺S�غm庇򺦮��������|�ED�!p���$��*���0���6��=�hC��#I�i/O��8U��?[�^Da��Gg�6Jm�rKs��Ky��L���������y���X���&���i�������޳��^����  �  �h=�=��=E=g�=u�=0=�� =�Y =��<�%�<�]�<*��<���<�<m5�<�h�<\��<���<���<�+�<�Y�<م�<��<n��<��<)�< N�<Nq�<ǒ�<���<^��<Z��<G�<-�<�3�<vG�<�X�<�g�<6t�<9~�<���<���<���<��<y��<��<�x�<*l�<�\�<�I�<�3�<!�<O��<���<0��<͑�<�f�<8�<��<~��<k��<�W�<��<E��<̆�<@9�<���<x��</9�<���<�z�<x�<Z��<j?�<�λ<�Y�<h�<*e�<F�<�a�<�ڲ<�O�<���<%0�<A��<0�<�g�<�ɧ<(�<僤<�ܢ<�2�<���<~ם<&�<Kr�<_��</�<	J�<���<Б<}�<(O�<���<WȊ<��<U<�<�t�<��<��<Y�<ך|<	y<Ulu<�q<Y;n<g�j<�	g<�pc<��_<A\<P�X<�U<x�Q<��M<�\J<��F<�@C<?�?<o.<<D�8<U'5<U�1<-.<S�*<wA'<��#<&f <I�<͜<q?<�<�<{F<w�<~�<B�<��;�5�;���;&��;h�;;?�;-$�;��;�;�+�;�K�;�{�;#��;�	�;�h�;פ;�U�;N�;��;2�;���;��;�=;�u;�k;�8a;%vW;F�M;�ND;�:;��1;jv(;+j;�z;C�;��;.��:ب�:���:OB�:�۵:���:��:,Ʌ:�Bl:�FM:��.:�T:4��9\K�9a]9�?�8e+������n�6$����湕���K*�(pE�]`�{�*ӊ�(�����G������˺[�غ	m�1�����|����J�uD�ap��$���*�u�0�3�6��=��C��#I��/O��8U�?[��Da��Gg�?Jm�}Ks�NLy��L�n���ʦ��2���k������f�������۳��j����  �  �h=�=��=!E=k�=t�=0=�� =�Y =��<�%�<�]�</��<���<� �<w5�<�h�<e��<���<���<�+�<�Y�<߅�<��<v��<��<)�<N�<Dq�<ʒ�<���<h��<]��<N�<'�<�3�<{G�<�X�<�g�<3t�<>~�<���<���<���<��<���<��<�x�<+l�<�\�<�I�<�3�<'�<S��< ��<.��<Ǒ�<�f�<8�<��<r��<t��<�W�<��<I��<Ć�<M9�<���<{��<+9�<���<�z�<u�<f��<e?�<�λ<�Y�<a�<1e�<G�<�a�<�ڲ<�O�<���<&0�<C��<-�<�g�<�ɧ<"(�<䃤<�ܢ<�2�<~��<�ם<&�<Ur�<R��<7�<J�<���<Б<m�<6O�<}��<WȊ<��<Y<�<�t�<��<��<M�<ۚ|<y<Wlu<�q<T;n<h�j<u	g<�pc<��_<A\<[�X<�U<|�Q<��M<�\J<��F<�@C<N�?<l.<<E�8<G'5<l�1<-.<T�*<�A'<��#<8f <)�<�<�?<'�<�<pF<��<{�<N�<��;�5�;���;"��;*h�;?�;:$�;��;F�;�+�;L�;�{�;ẵ;�	�;�h�;Mפ;�U�;b�;��;�1�;���;���;A>;�u;�k;�8a;'vW;��M;ND;>�:;��1;�v(;j;�z;��;��;���:��:���:�B�:�۵:���:���:�Ʌ:nAl:GM:2�.:&T:��9�J�9�	]9�;�8b�*�#���%n�_"��V��J��|L*��oE�-^`��{�ӊ�\��]����������˺�غm庸�V���N�������8D�3p�Ö$���*���0���6��=��C��#I�b/O�i8U�D?[��Da��Gg�/Jm�bKs�CLy�VL�x���Ȧ��x���{������J�������ڳ��a����  �  �h=�=��=E=i�=s�=7=�� =�Y =��<�%�<�]�<+��<���<� �<�5�<�h�<c��<���<���<�+�<Y�<��<ݰ�<r��<��<)�<	N�<:q�<Ғ�<���<k��<Q��<J�<2�<�3�<�G�<�X�<�g�<3t�<C~�<���<���<���<���<���<��<�x�<,l�<~\�<�I�<�3�<+�<E��<��<2��<ʑ�<�f�<8�<��<p��<x��<�W�<��<P��<���<N9�<���<���<*9�<���<�z�<u�<f��<Y?�<�λ<�Y�<i�</e�<9�<�a�<�ڲ<�O�<���<(0�<I��< �<�g�<{ɧ</(�<܃�<�ܢ<�2�<���<�ם<&�<br�<Q��<<�<J�<�<Б<m�<;O�<p��<aȊ<��<S<�<�t�<��<��<J�<ښ|<y<^lu<�q<H;n<��j<u	g<�pc<��_<A\<c�X<�U<��Q<��M<�\J<��F<�@C<E�?<f.<<a�8<-'5<q�1<-.<[�*<tA'<��#<If <(�<��<e?<!�<�<~F<�<b�<k�<̔�;�5�;���;,��;?h�;�>�;X$�;��;P�;n+�;�K�;�{�;뺵;
�;jh�;Cפ;�U�;v�;���;�1�;�;ο�;.>;/u;�k;�8a;�uW;��M;ND;^�:;9�1;�v(;>j;�z;ǧ;�; ��:���:���:�A�:�۵:b��:ݟ�:ʅ:@l:�HM:+�.:WS:���9oJ�9,	]9u/�8M�*�����:n��"�����)��M*��nE�W_`��{��Ҋ�-��k��r������˺r�غ�l府�S���ל�^����	D�@p��$���*���0���6�8=�>C��#I��/O��8U��?[�Da�Hg�4Jm�\Ks�'Ly��L���������y���<������l�������賗�T����  �  �h=�=��=E=m�=s�=1=�� =�Y =��<�%�<�]�<.��<���<� �<x5�<�h�<h��<���<���<�+�<�Y�<݅�<��<z��<��<)�<N�<Hq�<̒�<���<g��<]��<K�<-�<�3�<{G�<�X�<�g�<3t�<=~�<���<���<���<��<���<��<�x�<*l�<�\�<�I�<�3�<*�<S��<��<,��<Ƒ�<�f�<8�<��<q��<r��<�W�<��<F��<Æ�<L9�<���<~��</9�<���<�z�<v�<a��<i?�<�λ<�Y�<e�<-e�<G�<�a�<�ڲ<�O�<���<%0�<G��<*�<�g�<�ɧ<(�<ރ�<�ܢ<�2�<~��<�ם<&�<Vr�<O��</�<J�<���<Б<t�<4O�<y��<ZȊ<��<^<�<�t�<��<��<W�<ښ|<y<Wlu<�q<`;n<i�j<t	g<�pc<��_<A\<\�X<�U<�Q<��M<�\J<��F<�@C<V�?<g.<<H�8<;'5<i�1<-.<S�*<�A'<��#<+f <(�<�<s?<+�<�<{F<��<g�<J�<���;�5�;���;3��;h�;#?�;B$�;��;C�;�+�;�K�;�{�;�;�	�;�h�;<פ;�U�;^�;��;�1�;���;�;&>;�u;�k;�8a;�uW;��M;ND;W�:;��1;�v(;j;|z;��;��;���:��:c��:,B�:�۵:ƥ�:���:�Ʌ:�Al:}GM:��.:�T:��9�J�9�]93?�8%�*������n�]#��}�湟���L*��oE��]`��{��Ҋ����"����������˺,�غ�l庵������������rD�&p���$���*���0���6��=�vC��#I�B/O��8U�a?[��Da��Gg�4Jm��Ks�DLy�lL�_���Ǧ��z���g�������Y�����������[����  �  �h=�=��=E=k�=v�=/=�� =�Y =��<�%�<�]�<+��<���<�<v5�<�h�<_��<���<���<�+�<�Y�<څ�<��<q��<��<)�<N�<Nq�<���<���<c��<W��<E�<'�<�3�<pG�<�X�<�g�<<t�<9~�<���<���<���<��<z��<��<�x�<+l�<�\�<�I�<�3�< �<T��<���<3��<Б�<�f�<8�<��<v��<o��<�W�<��<B��<̆�<A9�<���<y��<.9�<���<�z�<��<Y��<f?�<�λ<�Y�<d�<'e�<B�<�a�<�ڲ<�O�<���<%0�<E��<,�<�g�<�ɧ<(�<胤<�ܢ<�2�<���<�ם<&�<Qr�<a��<6�<
J�<���<Б<t�<0O�<���<VȊ<��<^<�<�t�<��<��<Z�<̚|<y<clu<�q<P;n<U�j<�	g<�pc<��_<A\<`�X<�U<k�Q<��M<�\J<��F<�@C<P�?<r.<<B�8<S'5<b�1<-.<E�*<{A'<��#<6f <L�<ߜ<{?<�<�<qF<��<~�<D�<��;�5�;���;-��;#h�;=?�;$�;�;1�;�+�;�K�;�{�;��;�	�;�h�;פ;�U�;P�;��;�1�;���;��;�=;�u;�k;�8a;3vW;u�M;OND;�:;��1;�v(;Ij;�z;d�;��;?��:X��:-��:uB�:�۵:���:��:2Ʌ:�Bl:�FM:��.:9T:b��9jM�9�]9,<�8�>+�v����n��$�����M��K*�qE�M]`��{��Ҋ�n�����Z����U�˺*�غ;m庚�̮��[�����7�9D�Yp���$��*���0���6��=��C��#I�B/O��8U�#?[��Da��Gg�jJm�XKs�Ly��L����礪�6����������p�������ɳ�������  �  �h=�=��=E=i�=p�=3=�� =�Y =��<�%�<�]�<%��<���<� �<{5�<�h�<_��<���<���<�+�<�Y�<��<ݰ�<s��<��<)�<N�<Dq�<ɒ�<���<a��<V��<N�<,�<�3�<~G�<�X�<�g�<6t�<<~�<���<���<���<��<���<��<�x�<*l�<�\�<�I�<�3�<&�<L��<���<0��<ʑ�<�f�<8�<��<u��<t��<�W�<��<H��<���<H9�<���<~��<)9�<���<�z�<w�<^��<e?�<�λ<�Y�<e�<1e�<B�<�a�<�ڲ<�O�<���<$0�<D��<+�<�g�<}ɧ<%(�<ރ�<�ܢ<�2�<���<�ם<&�<Wr�<T��<9�<J�<���<Б<r�<7O�<x��<ZȊ<��<U<�<�t�<��<��<P�<ٚ|<y<Tlu<�q<W;n<q�j<�	g<�pc<��_<A\<P�X<�U<|�Q<��M<�\J<��F<�@C<H�?<Z.<<R�8<<'5<k�1<-.<]�*<xA'<��#<?f <*�<�<l?<�<�<vF<��<i�<Z�<˔�;�5�;���;!��;,h�;?�;3$�;��;(�;�+�;L�;�{�;��;�	�;�h�;*פ;�U�;X�;��;�1�;���;���;>;ju;�k;�8a;�uW;��M;8ND;6�:;r�1;�v(;0j;�z;��;b�;���:T��:{��:�A�:�۵:⥥:h��:�Ʌ:�Al:nGM:�.:�S:���9K�97]9D;�8j�*�:���`n�V"��ÿ�&��{L*��oE��^`�{�ӊ�x�����G��}����˺:�غ�l�<򺥮����������"D�|p���$���*���0���6��=�zC�$I��/O��8U�Z?[�qDa��Gg�7Jm�Ks�QLy��L�q�������U���_�������l�������೗�a����  �  �h=�=��= E=l�=q�=8=�� =�Y =��<�%�<�]�<,��<���<� �<�5�<�h�<i��<���<���<�+�<|Y�<��<ݰ�<���<��<)�<N�<@q�<ڒ�<��<m��<Y��<G�<.�<�3�<}G�<�X�<�g�<-t�<B~�<���<���<���<���<���<��<�x�<0l�<�\�<�I�<�3�<0�<N��<��<0��<ɑ�<�f�<8�<��<k��<x��<�W�<��<S��<���<T9�<���<}��<(9�<���<�z�<l�<i��<^?�<�λ<�Y�<e�<,e�<B�<�a�<|ڲ<�O�<���<%0�<>��<%�<�g�<|ɧ<0(�<ك�<�ܢ<�2�<|��<�ם<&�<_r�<P��<>�<J�<���<Б<g�<>O�<t��<eȊ<��<Y<�<�t�<���<��<I�<�|<y<Tlu<�q<M;n<r�j<d	g<�pc<��_<A\<\�X<�U<��Q<��M<�\J<��F<�@C<T�?<_.<<f�8</'5<}�1<�,.<Z�*<�A'<��#<Mf <&�<��<m?</�<�<iF<��<^�<n�<˔�; 6�;���;��;.h�;?�;y$�;��;Z�;�+�;�K�;�{�;׺�;�	�;h�;Tפ;�U�;q�;��;�1�;���;Ŀ�;v>;iu;�k;�8a;�uW;��M;�MD;��:;��1;�v(;-j;�z;ѧ;m�;_��:���:���:\B�:�۵:���:M��:lʅ:K@l:^GM:�.:T:���98H�9]9�4�8�*�T���2n��#����湨��
N*��mE��^`��{�aӊ�������\�����;�˺��غ$m���ۭ�����w�����C�0p�ؖ$�}�*�"�0���6�=�!C��#I�h/O�Q8U��?[�UDa�"Hg��Im��Ks�QLy�KL�������������^������K�����������,����  �  �h=�=��=E=h�=s�=2=�� =�Y =��<�%�<�]�<,��<���<� �<w5�<�h�<^��<���<���<�+�<Y�<��<��<t��<��<)�<N�<Fq�<͒�<���<g��<U��<H�<1�<�3�<|G�<�X�<�g�<.t�<?~�<���<���<���<��<���<��<�x�<'l�<�\�<�I�<�3�<%�<L��< ��<1��<ˑ�<�f�<8�<��<u��<w��<�W�<��<I��<���<H9�<���<���<09�<���<�z�<n�<e��<_?�<�λ<�Y�<k�<+e�<>�<�a�<�ڲ<�O�<���<+0�<H��<*�<�g�<ɧ<%(�<ۃ�<�ܢ<�2�<���<�ם<&�<Sr�<Y��<6�<J�<�<Б<t�<:O�<x��<XȊ<��<R<�<�t�<��<��<R�<ך|<	y<Wlu<�q<M;n<o�j<�	g<�pc<��_<A\<[�X<�U<}�Q<��M<�\J<��F<�@C<D�?<e.<<M�8<8'5<u�1<-.<S�*<rA'<��#<7f <=�<�<p?<�<�<~F<��<c�<W�<ߔ�;�5�;���;5��;Ih�;?�;C$�;��;B�;�+�;�K�;�{�;��;�	�;�h�;@פ;�U�;f�;��;�1�;���;���;#>;Ou;�k;�8a;vW;��M;=ND;0�:;o�1;�v(;3j;�z;�;b�;���:M��:���:hB�:R۵:���:6��:�Ʌ:�Al:CHM:ڤ.:�S:��9�H�9�]9`5�8��*�����/n��#�����h��EM*�=oE�'^`�.{��Ҋ�������,������˺سغ�l应򺿮��������|�@D�Bp��$���*���0���6��=��C��#I��/O�|8U�b?[�:Da��Gg�>Jm�~Ks�FLy�yL���������J���^������^�������򳗻_����  �  �h=�=��= E=j�=w�=0=�� =�Y =��<�%�<�]�<8��<���<� �<r5�<i�<Y��<���<���<�+�<�Y�<���<��<r��<��<)�<�M�<Hq�<Ȓ�<���<^��<W��<O�<"�<�3�<xG�<�X�<�g�<3t�<C~�<���<���<���<��<|��<��<�x�<&l�<�\�<�I�<�3�<�<X��<��<1��<ˑ�<�f�<8�<��<{��<m��<�W�<��<K��<Ȇ�<A9�<���<u��<+9�<���<�z�<t�<]��<g?�<�λ<�Y�<]�</e�<B�<�a�<�ڲ<�O�<���<0�<>��<.�<�g�<�ɧ<"(�<ރ�<�ܢ<�2�<���<{ם<%&�<Pr�<Y��<0�<J�<���<
Б<y�<+O�<{��<RȊ<��<X<�<�t�<	��<��<V�<Қ|<y<Qlu<�q<^;n<W�j<|	g<�pc<��_<A\<N�X<�U<t�Q<��M<�\J<��F<�@C<K�?<x.<<C�8<?'5<W�1<-.<O�*<vA'<��#<&f <:�<ל<�?<�<�<�F<l�<g�<Q�<��;�5�;���;��;h�;"?�;/$�;��;�;�+�;L�;�{�;캵;�	�;�h�;,פ;�U�;u�;��;�1�;���;���;�=;�u;�k;�8a;�uW;W�M;kND;��:;Ѡ1;�v(;6j;�z;��;��;��:���:��:�A�:n۵:��:⠕:;Ʌ:�Al:UFM:N�.:WT:n��9aJ�9]9=�8*�*�����an��"����湡��L*��oE��]`��{�_ӊ�O�����a�������˺��غ�l�.�$��������|�mD��o��$�Ѹ*���0��6��=��C��#I�k/O��8U�s?[��Da��Gg�SJm�MKs�\Ly��L�c���ꦅ�j�������祈�f�������ҳ��q����  �  �h=�=��=E=h�=s�=2=�� =�Y =��<�%�<�]�<,��<���<� �<w5�<�h�<^��<���<���<�+�<Y�<��<��<t��<��<)�<N�<Fq�<͒�<���<g��<U��<H�<1�<�3�<|G�<�X�<�g�<.t�<?~�<���<���<���<��<���<��<�x�<'l�<�\�<�I�<�3�<%�<L��< ��<1��<ˑ�<�f�<8�<��<u��<w��<�W�<��<I��<���<H9�<���<���<09�<���<�z�<n�<e��<_?�<�λ<�Y�<k�<+e�<>�<�a�<�ڲ<�O�<���<+0�<H��<*�<�g�<ɧ<%(�<ۃ�<�ܢ<�2�<���<�ם<&�<Sr�<Y��<6�<J�<�<Б<t�<:O�<x��<XȊ<��<R<�<�t�<��<��<R�<ך|<	y<Wlu<�q<M;n<o�j<�	g<�pc<��_<A\<[�X<�U<}�Q<��M<�\J<��F<�@C<D�?<e.<<M�8<8'5<u�1<-.<S�*<rA'<��#<7f <=�<�<p?<�<�<~F<��<c�<W�<ߔ�;�5�;���;5��;Ih�;?�;C$�;��;B�;�+�;�K�;�{�;��;�	�;�h�;@פ;�U�;f�;��;�1�;���;���;#>;Ou;�k;�8a;vW;��M;=ND;0�:;o�1;�v(;3j;�z;�;b�;���:M��:���:hB�:R۵:���:6��:�Ʌ:�Al:CHM:ڤ.:�S:��9�H�9�]9`5�8��*�����/n��#�����h��EM*�=oE�'^`�.{��Ҋ�������,������˺سغ�l应򺿮��������|�@D�Bp��$���*���0���6��=��C��#I��/O�|8U�b?[�:Da��Gg�>Jm�~Ks�FLy�yL���������J���^������^�������򳗻_����  �  �h=�=��= E=l�=q�=8=�� =�Y =��<�%�<�]�<,��<���<� �<�5�<�h�<i��<���<���<�+�<|Y�<��<ݰ�<���<��<)�<N�<@q�<ڒ�<��<m��<Y��<G�<.�<�3�<}G�<�X�<�g�<-t�<B~�<���<���<���<���<���<��<�x�<0l�<�\�<�I�<�3�<0�<N��<��<0��<ɑ�<�f�<8�<��<k��<x��<�W�<��<S��<���<T9�<���<}��<(9�<���<�z�<l�<i��<^?�<�λ<�Y�<e�<,e�<B�<�a�<|ڲ<�O�<���<%0�<>��<%�<�g�<|ɧ<0(�<ك�<�ܢ<�2�<|��<�ם<&�<_r�<P��<>�<J�<���<Б<g�<>O�<t��<eȊ<��<Y<�<�t�<���<��<I�<�|<y<Tlu<�q<M;n<r�j<d	g<�pc<��_<A\<\�X<�U<��Q<��M<�\J<��F<�@C<T�?<_.<<f�8</'5<}�1<�,.<Z�*<�A'<��#<Mf <&�<��<m?</�<�<iF<��<^�<n�<˔�; 6�;���;��;.h�;?�;y$�;��;Z�;�+�;�K�;�{�;׺�;�	�;h�;Tפ;�U�;q�;��;�1�;���;Ŀ�;v>;iu;�k;�8a;�uW;��M;�MD;��:;��1;�v(;-j;�z;ѧ;m�;_��:���:���:\B�:�۵:���:M��:lʅ:K@l:^GM:�.:T:���98H�9]9�4�8�*�T���2n��#����湨��
N*��mE��^`��{�aӊ�������\�����;�˺��غ$m���ۭ�����w�����C�0p�ؖ$�}�*�"�0���6�=�!C��#I�h/O�Q8U��?[�UDa�"Hg��Im��Ks�QLy�KL�������������^������K�����������,����  �  �h=�=��=E=i�=p�=3=�� =�Y =��<�%�<�]�<%��<���<� �<{5�<�h�<_��<���<���<�+�<�Y�<��<ݰ�<s��<��<)�<N�<Dq�<ɒ�<���<a��<V��<N�<,�<�3�<~G�<�X�<�g�<6t�<<~�<���<���<���<��<���<��<�x�<*l�<�\�<�I�<�3�<&�<L��<���<0��<ʑ�<�f�<8�<��<u��<t��<�W�<��<H��<���<H9�<���<~��<)9�<���<�z�<w�<^��<e?�<�λ<�Y�<e�<1e�<B�<�a�<�ڲ<�O�<���<$0�<D��<+�<�g�<}ɧ<%(�<ރ�<�ܢ<�2�<���<�ם<&�<Wr�<T��<9�<J�<���<Б<r�<7O�<x��<ZȊ<��<U<�<�t�<��<��<P�<ٚ|<y<Tlu<�q<W;n<q�j<�	g<�pc<��_<A\<P�X<�U<|�Q<��M<�\J<��F<�@C<H�?<Z.<<R�8<<'5<k�1<-.<]�*<xA'<��#<?f <*�<�<l?<�<�<vF<��<i�<Z�<˔�;�5�;���;!��;,h�;?�;3$�;��;(�;�+�;L�;�{�;��;�	�;�h�;*פ;�U�;X�;��;�1�;���;���;>;ju;�k;�8a;�uW;��M;8ND;6�:;r�1;�v(;0j;�z;��;b�;���:T��:{��:�A�:�۵:⥥:h��:�Ʌ:�Al:nGM:�.:�S:���9K�97]9D;�8j�*�:���`n�V"��ÿ�&��{L*��oE��^`�{�ӊ�x�����G��}����˺:�غ�l�<򺥮����������"D�|p���$���*���0���6��=�zC�$I��/O��8U�Z?[�qDa��Gg�7Jm�Ks�QLy��L�q�������U���_�������l�������೗�a����  �  �h=�=��=E=k�=v�=/=�� =�Y =��<�%�<�]�<+��<���<�<v5�<�h�<_��<���<���<�+�<�Y�<څ�<��<q��<��<)�<N�<Nq�<���<���<c��<W��<E�<'�<�3�<pG�<�X�<�g�<<t�<9~�<���<���<���<��<z��<��<�x�<+l�<�\�<�I�<�3�< �<T��<���<3��<Б�<�f�<8�<��<v��<o��<�W�<��<B��<̆�<A9�<���<y��<.9�<���<�z�<��<Y��<f?�<�λ<�Y�<d�<'e�<B�<�a�<�ڲ<�O�<���<%0�<E��<,�<�g�<�ɧ<(�<胤<�ܢ<�2�<���<�ם<&�<Qr�<a��<6�<
J�<���<Б<t�<0O�<���<VȊ<��<^<�<�t�<��<��<Z�<̚|<y<clu<�q<P;n<U�j<�	g<�pc<��_<A\<`�X<�U<k�Q<��M<�\J<��F<�@C<P�?<r.<<B�8<S'5<b�1<-.<E�*<{A'<��#<6f <L�<ߜ<{?<�<�<qF<��<~�<D�<��;�5�;���;-��;#h�;=?�;$�;�;1�;�+�;�K�;�{�;��;�	�;�h�;פ;�U�;P�;��;�1�;���;��;�=;�u;�k;�8a;3vW;u�M;OND;�:;��1;�v(;Ij;�z;d�;��;?��:X��:-��:uB�:�۵:���:��:2Ʌ:�Bl:�FM:��.:9T:b��9jM�9�]9,<�8�>+�v����n��$�����M��K*�qE�M]`��{��Ҋ�n�����Z����U�˺*�غ;m庚�̮��[�����7�9D�Yp���$��*���0���6��=��C��#I�B/O��8U�#?[��Da��Gg�jJm�XKs�Ly��L����礪�6����������p�������ɳ�������  �  �h=�=��=E=m�=s�=1=�� =�Y =��<�%�<�]�<.��<���<� �<x5�<�h�<h��<���<���<�+�<�Y�<݅�<��<z��<��<)�<N�<Hq�<̒�<���<g��<]��<K�<-�<�3�<{G�<�X�<�g�<3t�<=~�<���<���<���<��<���<��<�x�<*l�<�\�<�I�<�3�<*�<S��<��<,��<Ƒ�<�f�<8�<��<q��<r��<�W�<��<F��<Æ�<L9�<���<~��</9�<���<�z�<v�<a��<i?�<�λ<�Y�<e�<-e�<G�<�a�<�ڲ<�O�<���<%0�<G��<*�<�g�<�ɧ<(�<ރ�<�ܢ<�2�<~��<�ם<&�<Vr�<O��</�<J�<���<Б<t�<4O�<y��<ZȊ<��<^<�<�t�<��<��<W�<ښ|<y<Wlu<�q<`;n<i�j<t	g<�pc<��_<A\<\�X<�U<�Q<��M<�\J<��F<�@C<V�?<g.<<H�8<;'5<i�1<-.<S�*<�A'<��#<+f <(�<�<s?<+�<�<{F<��<g�<J�<���;�5�;���;3��;h�;#?�;B$�;��;C�;�+�;�K�;�{�;�;�	�;�h�;<פ;�U�;^�;��;�1�;���;�;&>;�u;�k;�8a;�uW;��M;ND;W�:;��1;�v(;j;|z;��;��;���:��:c��:,B�:�۵:ƥ�:���:�Ʌ:�Al:}GM:��.:�T:��9�J�9�]93?�8%�*������n�]#��}�湟���L*��oE��]`��{��Ҋ����"����������˺,�غ�l庵������������rD�&p���$���*���0���6��=�vC��#I�B/O��8U�a?[��Da��Gg�4Jm��Ks�DLy�lL�_���Ǧ��z���g�������Y�����������[����  �  �h=�=��=E=i�=s�=7=�� =�Y =��<�%�<�]�<+��<���<� �<�5�<�h�<c��<���<���<�+�<Y�<��<ݰ�<r��<��<)�<	N�<:q�<Ғ�<���<k��<Q��<J�<2�<�3�<�G�<�X�<�g�<3t�<C~�<���<���<���<���<���<��<�x�<,l�<~\�<�I�<�3�<+�<E��<��<2��<ʑ�<�f�<8�<��<p��<x��<�W�<��<P��<���<N9�<���<���<*9�<���<�z�<u�<f��<Y?�<�λ<�Y�<i�</e�<9�<�a�<�ڲ<�O�<���<(0�<I��< �<�g�<{ɧ</(�<܃�<�ܢ<�2�<���<�ם<&�<br�<Q��<<�<J�<�<Б<m�<;O�<p��<aȊ<��<S<�<�t�<��<��<J�<ښ|<y<^lu<�q<H;n<��j<u	g<�pc<��_<A\<c�X<�U<��Q<��M<�\J<��F<�@C<E�?<f.<<a�8<-'5<q�1<-.<[�*<tA'<��#<If <(�<��<e?<!�<�<~F<�<b�<k�<̔�;�5�;���;,��;?h�;�>�;X$�;��;P�;n+�;�K�;�{�;뺵;
�;jh�;Cפ;�U�;v�;���;�1�;�;ο�;.>;/u;�k;�8a;�uW;��M;ND;^�:;9�1;�v(;>j;�z;ǧ;�; ��:���:���:�A�:�۵:b��:ݟ�:ʅ:@l:�HM:+�.:WS:���9oJ�9,	]9u/�8M�*�����:n��"�����)��M*��nE�W_`��{��Ҋ�-��k��r������˺r�غ�l府�S���ל�^����	D�@p��$���*���0���6�8=�>C��#I��/O��8U��?[�Da�Hg�4Jm�\Ks�'Ly��L���������y���<������l�������賗�T����  �  �h=�=��=!E=k�=t�=0=�� =�Y =��<�%�<�]�</��<���<� �<w5�<�h�<e��<���<���<�+�<�Y�<߅�<��<v��<��<)�<N�<Dq�<ʒ�<���<h��<]��<N�<'�<�3�<{G�<�X�<�g�<3t�<>~�<���<���<���<��<���<��<�x�<+l�<�\�<�I�<�3�<'�<S��< ��<.��<Ǒ�<�f�<8�<��<r��<t��<�W�<��<I��<Ć�<M9�<���<{��<+9�<���<�z�<u�<f��<e?�<�λ<�Y�<a�<1e�<G�<�a�<�ڲ<�O�<���<&0�<C��<-�<�g�<�ɧ<"(�<䃤<�ܢ<�2�<~��<�ם<&�<Ur�<R��<7�<J�<���<Б<m�<6O�<}��<WȊ<��<Y<�<�t�<��<��<M�<ۚ|<y<Wlu<�q<T;n<h�j<u	g<�pc<��_<A\<[�X<�U<|�Q<��M<�\J<��F<�@C<N�?<l.<<E�8<G'5<l�1<-.<T�*<�A'<��#<8f <)�<�<�?<'�<�<pF<��<{�<N�<��;�5�;���;"��;*h�;?�;:$�;��;F�;�+�;L�;�{�;ẵ;�	�;�h�;Mפ;�U�;b�;��;�1�;���;���;A>;�u;�k;�8a;'vW;��M;ND;>�:;��1;�v(;j;�z;��;��;���:��:���:�B�:�۵:���:���:�Ʌ:nAl:GM:2�.:&T:��9�J�9�	]9�;�8b�*�#���%n�_"��V��J��|L*��oE�-^`��{�ӊ�\��]����������˺�غm庸�V���N�������8D�3p�Ö$���*���0���6��=��C��#I�b/O�i8U�D?[��Da��Gg�/Jm�bKs�CLy�VL�x���Ȧ��x���{������J�������ڳ��a����  �  �h=�=��=E=g�=u�=0=�� =�Y =��<�%�<�]�<*��<���<�<m5�<�h�<\��<���<���<�+�<�Y�<م�<��<n��<��<)�< N�<Nq�<ǒ�<���<^��<Z��<G�<-�<�3�<vG�<�X�<�g�<6t�<9~�<���<���<���<��<y��<��<�x�<*l�<�\�<�I�<�3�<!�<O��<���<0��<͑�<�f�<8�<��<~��<k��<�W�<��<E��<̆�<@9�<���<x��</9�<���<�z�<x�<Z��<j?�<�λ<�Y�<h�<*e�<F�<�a�<�ڲ<�O�<���<%0�<A��<0�<�g�<�ɧ<(�<僤<�ܢ<�2�<���<~ם<&�<Kr�<_��</�<	J�<���<Б<}�<(O�<���<WȊ<��<U<�<�t�<��<��<Y�<ך|<	y<Ulu<�q<Y;n<g�j<�	g<�pc<��_<A\<P�X<�U<x�Q<��M<�\J<��F<�@C<?�?<o.<<D�8<U'5<U�1<-.<S�*<wA'<��#<&f <I�<͜<q?<�<�<{F<w�<~�<B�<��;�5�;���;&��;h�;;?�;-$�;��;�;�+�;�K�;�{�;#��;�	�;�h�;פ;�U�;N�;��;2�;���;��;�=;�u;�k;�8a;%vW;F�M;�ND;�:;��1;jv(;+j;�z;C�;��;.��:ب�:���:OB�:�۵:���:��:,Ʌ:�Bl:�FM:��.:�T:4��9\K�9a]9�?�8e+������n�6$����湕���K*�(pE�]`�{�*ӊ�(�����G������˺[�غ	m�1�����|����J�uD�ap��$���*�u�0�3�6��=��C��#I��/O��8U�?[��Da��Gg�?Jm�}Ks�NLy��L�n���ʦ��2���k������f�������۳��j����  �  �h=�=��=E=k�=s�=3=�� =�Y =��<�%�<�]�<0��<���<� �<|5�<�h�<`��<���<���<�+�<�Y�<��<��<u��<��<)�<N�<Bq�<Β�<���<i��<V��<C�<0�<�3�<{G�<�X�<�g�<9t�<>~�<���<���<���<��<��<��<�x�<(l�<�\�<�I�<�3�<#�<N��<��</��<ˑ�<�f�<8�<��<r��<p��<�W�<��<G��<ǆ�<H9�<���<��<+9�<���<�z�<z�<`��<a?�<�λ<�Y�<g�<*e�<@�<�a�<�ڲ<�O�<���<%0�<B��<%�<�g�<�ɧ<#(�<���<�ܢ<�2�<���<�ם<&�<Zr�<Y��<5�<J�<���<	Б<t�<2O�<z��<\Ȋ<��<Y<�<�t�<��<��<O�<ښ|<y<jlu<�q<K;n<q�j<u	g<�pc<��_<
A\<h�X<�U<~�Q<��M<�\J<��F<�@C<L�?<g.<<S�8<?'5<g�1<-.<D�*<vA'<��#<9f <;�<�<u?<�<�<sF<��<m�<T�<��;�5�;���;��;%h�;?�;H$�;��;I�;�+�;�K�;�{�;���;�	�;�h�;-פ;�U�;`�;	��;�1�;���;ῄ;>;�u;�k;�8a;�uW;��M;!ND;�:;��1;�v(;%j;�z;��;y�;y��:&��:A��:�A�:s۵:֥�:ʠ�:�Ʌ:Al:�GM:L�.:�S:R��9�K�9]9i7�8��*�q���Vn�$��N�湢��,L*�YoE��^`��{�*ӊ����o����������˺S�غm庇򺦮��������|�ED�!p���$��*���0���6��=�hC��#I�i/O��8U��?[�^Da��Gg�6Jm�rKs��Ky��L���������y���X���&���i�������޳��^����  �  �h=�=��="E=k�=m�=4=�� =�Y =��<�%�<�]�<(��<���<� �<}5�<�h�<j��<���<���<�+�<}Y�<��<ذ�<��<��<)�<N�<@q�<Ԓ�<~��<l��<Y��<M�<3�<�3�<�G�<�X�<�g�</t�<=~�<���<���<���<���<���<��<�x�<(l�<�\�<�I�<�3�</�<M��<��<.��<Ƒ�<�f�<8�<��<f��<~��<�W�<��<F��<���<U9�<���<���<,9�<���<�z�<p�<m��<c?�<�λ<�Y�<g�<3e�<C�<�a�<ڲ<�O�<���<.0�<L��<&�<�g�<xɧ<&(�<ۃ�<�ܢ<�2�<z��<�ם<&�<Yr�<L��<7�<	J�<���<Б<i�<DO�<t��<\Ȋ<��<W<�<�t�<��<��<H�<�|<�y<^lu<�q<N;n<��j<s	g<�pc<��_<A\<a�X<�U<��Q<��M<�\J<��F<�@C<N�?<O.<<V�8<0'5<��1<-.<W�*<�A'<��#<:f <�<�<k?</�<�<qF<��<_�<[�<���;�5�;���;2��;Ph�;?�;`$�;��;V�;�+�;L�;�{�;躵;
�;�h�;aפ;�U�;]�;+��;�1�;�;ֿ�;x>;Uu;|k;�8a;�uW;��M;�MD;~�:;v�1;�v(;j;z;��;K�;5��:f��:��:B�:l۵:���:��:oʅ:�@l:�HM:S�.:�T:��97I�9�]9L9�8V�*�]���=n��!����湢���M*��nE�l^`��{�~Ҋ����������r���˺߳غ�l��� �����������4D�^p�ؖ$�|�*��0�[�6�=�fC�-$I�x/O�<8U��?[�Da�%Hg��Im��Ks�)Ly�QL���������}���9������Q����������:����  �  �h=�=��=E=j�=t�=7=�� =�Y =��<�%�<�]�<*��<���< �<{5�<�h�<d��<���<���<�+�<�Y�<��<��<w��<��<)�<N�<Eq�<В�<���<d��<S��<I�<,�<�3�<xG�<�X�<�g�<5t�<A~�<���<���<���< ��<���<��<�x�<0l�<�\�<�I�<�3�<)�<K��< ��<5��<ϑ�<�f�<8�<��<k��<w��<�W�<��<N��<ņ�<H9�<���<��<'9�<���<�z�<x�<^��<b?�<�λ<�Y�<f�<,e�<?�<�a�<�ڲ<�O�<���<#0�<F��<#�<�g�<�ɧ<*(�<⃤<�ܢ<�2�<{��<�ם<&�<Wr�<\��<:�<J�<���<Б<l�<6O�<{��<cȊ<��<W<�<�t�<	��<��<K�<�|<y<_lu<	�q<P;n<j�j<�	g<�pc<��_<A\<]�X<�U<��Q<��M<�\J<��F<�@C<K�?<j.<<a�8<A'5<j�1<-.<R�*<}A'<��#<<f <?�<�<j?<#�<�<vF<�<p�<c�<��;�5�;���;-��;h�;?�;Q$�;��;4�;u+�;�K�;�{�;��;�	�;�h�;%פ;�U�;m�;!��;�1�;���;޿�;>;�u;�k;�8a;�uW;��M;�MD;N�:;f�1;�v(;Vj;�z;��;K�;��:���:���:B�:�۵:A��:���:�Ʌ:�@l:�GM:��.:�T:��9FK�9+]9e8�8��*������n��#��k�����L*�6oE��]`�>{��Ҋ� ��W�����.����˺H�غ�l���X���������c�D�Np���$���*���0���6��=�2C��#I�z/O��8U�q?[�mDa�Hg�Jm�YKs�%Ly��L����Ŧ��M���e������s�������ݳ��G����  �  �i=�=��=9F=��=݂=� =T� =�[ =��<#*�<�b�<��<���<��<R;�<:o�<���<���<0�<x3�<�a�<H��<ӹ�<���<A�<03�<�X�<`|�<)��<j��<���<%��<��<�+�<#B�<%V�<h�<\w�<i��<ێ�<��<I��<���<���<���<���<���<���<q�<_�<vI�<i0�<�<��<���<���<�~�<�P�<S�<f��<���<�p�<s/�<���<���<%S�<��<f��<)S�<���<^��<(/�<�ž<�X�<��<�r�<���<W}�< ��<y�<��<ff�<�ׯ<�E�<`��<��<�{�<ݧ<�:�<��<S�<�C�<���< �<5�<���<�ɘ<�<0V�<e��<�ڑ<l�<^X�<���<
Њ<�	�<�B�<"z�<Ѱ�<�<��<̟|<}y<\nu<��q<m:n<ԟj<vg<Akc<��_<y8\<T�X<8	U<^sQ<{�M<�LJ<2�F<�-C<ɡ?<�<<��8<Y5<�1<J.<��*<�"'<��#<�D <g�<�x<�</�<�k<�<��<��<S<�8�;��;��;M<�;\�;��;���;��;���;Ǿ�;���;r�;�J�;���;��;�d�;��;�p�;��;;�;=}�;�L�;X~;8t;7j;fV`;��V;��L;rC;H:;��0;D�';͘;��;��;V);{!�:�'�:�a�:���:^r�:^D�:�H�:�x�:G�i:o�J:�8,:�:��9�פ9�]T9�8r������%�u�Բ��L�_����+��	G���a�Ĕ|�����q���4å�e���w���~̺�Bٺ���ȗ�P*������[G��v�ǟ���$�M�*�Z�0��7��&=�>6C��AI�#KO�5RU�LV[��Ya�Yg��Zm��Ys�AXy��V�&���©��8���B����������8���v�������  �  �i=�=��=:F=��=ׂ=� =X� =�[ =��<2*�<�b�<��<���<��<];�<-o�<���<���<8�<3�<�a�<W��<Ź�<���<9�<23�<�X�<9|�<0��<h��<���<#��<��<�+�<&B�<(V�<�g�<Yw�<^��<��<Ԗ�<)��<Ȟ�<���<���<���<���<���<�q�<$_�<{I�<t0�<��<��<���<���<�~�<yP�<]�<p��<���< q�<�/�<���<���<*S�<��<l��<S�<���<c��</�<�ž<�X�<��<�r�<���<W}�<��<!y�<��<jf�<�ׯ<�E�<b��<��<�{�<�ܧ<�:�<#��<[�<�C�<Ӗ�<&�<5�<���<�ɘ<�<(V�<Y��<�ڑ<j�<kX�<���<Њ<�	�<�B�<)z�<ΰ�<��<��<̟|<�y<Wnu<��q<J:n<ܟj<~g<Ekc<��_<�8\<Q�X<=	U<isQ<-�M<�LJ<1�F<�-C<ʡ?<k<<ߑ8<e5<�1<F.<�*<�"'<��#<�D <T�<�x<�<2�<�k<<��<��<1S<s8�;��;���;U<�;:�;i��;Ի�;���;ɮ�;���;���;}�;�J�;���;���;�d�;��;q�;��;N��;Y}�;�L�;YX~;�7t;7j;�V`;̕V;c�L;/rC;�:;=�0;"�';И;f�;��;�(;"�:4(�:c�:H��:*s�:�D�:+H�:=y�:��i:)�J:85,:S�:��9�Ԥ9�\T9l�8Q������u��Ӳ��N�ݪ���+��	G��a�ǖ|��������å�M��������}̺MBٺ�废���)��o�����G��v����$���*�k�0�!7��&=��5C��AI�%KO��QU�eV[��Ya��Zg��Zm��Ys�WXy��V�n�������'���<���ϩ�����<���l���괚��  �  �i=�=��=;F=��=҂=� =O� =�[ =��<.*�<�b�<��<���<w�<k;�<,o�<���<���<*�<3�<�a�<]��<���<���<6�<13�<�X�<8|�<H��<]��<���<!��<��<�+�<B�<1V�<�g�<cw�<V��<��<��<*��<מ�<���<���<���<���<���<xq�<$_�<gI�<t0�<��<��<���<���<�~�<yP�<^�<]��<���<�p�<x/�<���<���<4S�<��<x��<S�<���<t��</�<�ž<�X�<��<�r�<���<Y}�<��<(y�<��<�f�<�ׯ<�E�<g��<��<�{�<�ܧ<�:�<��<Y�<�C�<Ė�<&�<5�<���<�ɘ<�<.V�<Z��<�ڑ<V�<mX�<锌<Њ<�	�<�B�<.z�<°�<��<��<��|<�y<Inu<��q<;:n<�j<og<Skc<~�_<�8\<G�X<4	U<�sQ<%�M<�LJ< �F<�-C<ݡ?<X<<�8<D5<
�1<".<�*<�"'<��#<�D <*�<�x<�<0�<�k<�<��<r�<<S<;8�;>��;��;T<�;u�;h��;4��;խ�;Ԯ�;���;���;��;�J�;ᘯ;���;�d�;��;:q�;��;S��;�}�;�L�;�X~;�7t;7j;�V`;W�V;d�L;�qC;�:;9�0;��';��;0�;��;�(;."�:'�:�b�:���:�r�:�D�:~G�:�y�:��i:��J:�5,:)�:�9~Ҥ9GaT9�g�8���c��X�u�tӲ��O���*�+��G�M�a�4�|�8���d���N¥�!���n���b~̺{Bٺ��应���)��o��G�%H�Sv�؟�	�$���*��0�7�'=��5C�4BI�
KO��QU��V[��Xa��Zg�%Zm��Ys��Xy�TV���������G������橎�󪑻P���~��������  �  �i=�=��=;F=��=ق=� =Q� =�[ =��<+*�<�b�<��<���<��<_;�<,o�<���<���<6�<�3�<�a�<_��<Ĺ�<���<=�</3�<�X�<;|�<0��<_��<���<��<��<�+�<B�<.V�<�g�<\w�<`��<ێ�<Ֆ�<.��<˞�<���<���<���<���<���<�q�<-_�<uI�<q0�<��<��<���<���<�~�<{P�<[�<i��<���<q�<}/�<��<���<-S�<��<k��<S�<���<_��</�<�ž<�X�<��<�r�<���<_}�<��<'y�<��<if�<�ׯ<�E�<a��<��<�{�<�ܧ<;�<��<g�<�C�<ǖ�<)�<5�<���<�ɘ<�<(V�<c��<�ڑ<e�<uX�<<Њ<�	�<�B�<*z�<ǰ�<��<��<Ο|<vy<]nu<��q<Q:n<�j<bg<Zkc<��_<8\<U�X<*	U<esQ<2�M<�LJ<$�F<�-C<ӡ?<r<<�8<I5<�1<B.<�*<�"'<��#<�D <K�<�x<�<;�<�k<<��<r�<AS<l8�;��;��;I<�;_�;t��;Ի�;ۭ�;ܮ�;���;���;��;�J�;Ԙ�;���;�d�;��;�p�;��;b��;g}�;�L�;pX~;�7t;a7j;�V`;V;��L;rC;�:;O�0;>�';��;]�;��;�(;�!�:�'�:_c�:���:s�:oE�:�G�:yy�:|�i:
�J:*6,:��:��9�Ԥ9_T9�p�8����J���u�Ҳ�MO�8����+��	G���a���|����������¥�s���&���P~̺�Aٺ8��Y���)��s�����G��v�����$��*���0��7��&=��5C��AI�!KO��QU��V[�JYa��Zg��Zm�Zs�?Xy��V�`�������`�������������4�������𴚻�  �  �i=�=��=;F=��=ق=� =T� =�[ =��<**�<�b�<��<���<��<Z;�<5o�<���<���<.�<|3�<�a�<U��<ɹ�<���<A�<53�<�X�<D|�<1��<s��<���<��<��<�+�< B�<&V�<�g�<Nw�<i��<��<ۖ�<5��<ƞ�<���<���<���<���<���<�q�<_�<xI�<m0�<�<��<���<���<�~�<�P�<V�<m��<���< q�<q/�<���<���<"S�<��<k��<S�<���<k��<)/�<�ž<�X�<��<�r�<���<]}�<��<y�<��<lf�<�ׯ<�E�<f��<��<�{�<�ܧ<�:�<��<Z�<�C�<Ζ�<$�<5�<���<�ɘ<�<,V�<c��<�ڑ<d�<cX�<���<Њ<�	�<�B�<(z�<԰�<��<��<П|<�y<anu<v�q<X:n<ԟj<ug<Akc<��_<u8\<R�X<S	U<hsQ<E�M<�LJ<<�F<�-C<š?<s<<ϑ8<W5<��1<9.<
�*<�"'<��#<�D <_�<�x<�<:�<�k<�<��<v�<,S<�8�;���;��;c<�;P�;���;ػ�;-��;���;���;���;q�;�J�;���;���;�d�;��;1q�;��;}��;R}�;�L�;)X~;�7t;7j;nV`;��V;	�L;rC;j:;��0;5�';ݘ;��;v�;);�!�:(�:.b�:N��:Br�:�D�:&H�:�x�:��i:��J:�6,:��:��97ؤ9�WT9�r�8
������o�u�}Ҳ�bO�ʫ�2�+�D	G���a���|�I��������å����Ĩ��p~̺fBٺ�����*��&����vG��v�����$�(�*���0�]7��&=�6C��AI�5KO�RU�5V[��Ya�\Zg��Zm�wYs�.Xy��V�R�������9���C�������$���:���A���봚��  �  �i=�=��=8F=��=ق=� =W� =�[ =��<-*�<�b�<��<���<~�<e;�<5o�<��<���<2�<�3�<�a�<U��<ƹ�<���<6�<+3�<�X�<@|�<4��<_��<���<'��<��<�+�<*B�<&V�<�g�<^w�<T��<��<ܖ�<0��<͞�<���<���<���<���<���<�q�<"_�<uI�<i0�<��<��<���<���<�~�<�P�<Q�<i��<���<q�<s/�<���<���<+S�<��<q��<S�<���<g��</�<�ž<�X�<��<�r�<���<[}�<��<y�<��<nf�<�ׯ<�E�<b��<��<�{�<�ܧ<�:�<��<`�<�C�<̖�<�<5�<���<�ɘ<�<2V�<X��<�ڑ<e�<oX�<���<Њ<�	�<�B�<%z�<ư�<��<��<ן|<~y<=nu<��q<T:n<ϟj<�g<<kc<��_<�8\<6�X<4	U<psQ<;�M<�LJ<!�F<�-C<ڡ?<q<<Б8<b5<�1<;.<�*<�"'<��#<�D <8�<�x<�<�<�k<�<��<��<,S<u8�;-��;��;<<�;e�;���;��;ݭ�;���;Ͼ�;���;o�;�J�;���;���;�d�;��;q�;��;h��;n}�;�L�;YX~;�7t;07j;�V`;ՕV;W�L;�qC;N:;d�0;��';��;E�;��;);b!�:�'�:�b�:p��:`r�:E�:H�:Yy�:x�i:��J:E6,:i�:��9�Ҥ9y]T9u�8���������u��Ҳ��M�m����+��G� �a�i�|�~���;����¥�f�������~̺Bٺ������*��&��m��G�v�����$��*���0��7��&=�6C��AI��JO�RU��V[�ZYa�|Zg��Zm��Ys��Xy�PV�Z���˩�����N�������񪑻s���~���ܴ���  �  �i=�=��=;F=��=ւ=� =Q� =�[ =��<2*�<�b�<��<���<��<`;�<(o�<���<���<4�<�3�<�a�<`��<���<���<7�</3�<�X�<8|�<<��<c��<���<��<��<�+�<!B�<*V�<�g�<^w�<\��<��<ז�<+��<Ԟ�<���<���<���<���<���<~q�<(_�<sI�<u0�<��<��<���<���<�~�<vP�<]�<g��<���<�p�<t/�<��<���<3S�<��<x��<S�<���<m��</�<�ž<�X�<��<�r�<���<Y}�<��<(y�<��<vf�<�ׯ<�E�<g��<��<�{�<�ܧ<;�<��<^�<�C�<̖�<'�<�4�<���<�ɘ<�<'V�<Z��<�ڑ<c�<rX�<<Њ<�	�<�B�<.z�<Ű�<��<��<ן|<�y<Xnu<��q<8:n<�j<wg<Qkc<~�_<x8\<U�X<?	U<vsQ<*�M<�LJ< �F<�-C<ˡ?<e<<�8<L5<�1<>.<�*<�"'<��#<�D <T�<�x<�<7�<�k<<��<r�<CS<S8�;0��;��;I<�;r�;f��;��;��;߮�;���;���;��;�J�;Ƙ�;���;�d�;��;,q�;��;T��;�}�;�L�;�X~;�7t;b7j;�V`;��V;��L;�qC;�:;-�0;E�';�;x�;��;�(;!"�:�'�:c�:��:xr�:�E�:yG�:�y�:��i:��J:�5,:��:a�9Ԥ9�^T9Ue�8������͵u��Ӳ�Q���P�+��G��a�R�|�4���b���{¥�쿲�
����~̺'BٺY�����)��������G�vv����$���*���0��7��&=��5C�BI�<KO��QU��V[�,Ya��Zg��Zm��Ys�SXy��V���������5���$���穎����4���i���Ѵ���  �  �i=�=��=>F=��=ւ=� =U� =�[ =
��<"*�<�b�<��<���<��<W;�<8o�<��<���<-�<�3�<�a�<Z��<���<���<@�<03�<�X�<B|�<9��<e��<���<��<��<�+�<B�<2V�<�g�<Pw�<^��<��<ۖ�<0��<ɞ�<���<���<���<���<���<�q�<!_�<pI�<k0�<�<��<���<���<�~�<�P�<Y�<c��<���<q�<v/�<���<���<,S�<��<n��<S�<���<h��</�<�ž<�X�<��<�r�<���<c}�<��<y�<��<qf�<�ׯ<�E�<c��<��<�{�<�ܧ<�:�<��<a�<�C�<�<)�<5�<���<�ɘ<
�<0V�<g��<�ڑ<_�<jX�<���<Њ<�	�<�B�</z�<Ͱ�<��<��<՟|<�y<Tnu<o�q<S:n<�j<[g<Rkc<��_<i8\<N�X<;	U<rsQ<?�M<�LJ<.�F<�-C<��?<e<<ߑ8<]5<	�1<4.<��*<�"'<��#<�D <h�<�x<�<C�<�k<�<��<��<8S<W8�;
��;��;N<�;M�;���;���;���;���;���;���;�;�J�;蘯;���;�d�;��;q�;��;j��;_}�;�L�;}X~;�7t;77j;�V`;ЕV;M�L;�qC;^:;��0;E�';ʘ;��;��;6);�!�:o'�:�b�:n��:�r�:9E�:�G�:fy�:��i:`�J:�5,:k�:�9�Ԥ9�XT9�r�8	n�����u��в��O�p���+��G���a��|�u���Ͱ��å�����q���*~̺�Aٺ��庳��)��
����PG��v�ɟ���$�Q�*���0�#7��&=��5C�BI�SKO��QU�iV[��Ya�qZg��Zm��Ys�cXy��V�\�������m���"�������<���C���p���״���  �  �i=�=��=8F=��=܂=� =X� =�[ =��<.*�<�b�<��<���<��<Y;�<9o�<��<���<:�<�3�<�a�<S��<̹�<���<:�</3�<�X�<=|�<,��<e��<���<"��<��<�+�<%B�<#V�<�g�<Yw�<`��<ߎ�<֖�<+��<Ȟ�<���<���<���<���<���<�q�<_�<�I�<f0�<�<��<���<���<�~�<�P�<O�<x��<���<q�<z/�<���<���<!S�<��<k��<S�<���<`��</�<�ž<�X�<��<�r�<���<Z}�<��<y�<��<ff�<�ׯ<�E�<`��<��<�{�<�ܧ<�:�< ��<_�<�C�<ז�<�<5�<���<�ɘ<
�<2V�<]��<�ڑ<s�<hX�<���<Њ<�	�<�B�< z�<Ѱ�<��<��<Ɵ|<�y<Unu<��q<P:n<ןj<�g<Akc<��_<�8\<J�X<7	U<`sQ<4�M<�LJ<1�F<�-C<С?<�<<͑8<h5<�1<V.<�*<�"'<��#<�D <R�<�x<�<�<�k<<��<��<(S<�8�;��;���;J<�;B�;}��;ǻ�;���;���;���;���;x�;�J�;���;���;�d�;��;q�;��;U��;Y}�;�L�;X~;8t;97j;�V`;�V;?�L;~rC;5:;o�0;W�';͘;q�;��;);<!�:�(�:�b�:���:�r�:�D�:�H�:�x�:�i:�J:�5,:�::�9xդ9�[T9fr�8����?����u�dӲ�jN�5����+��	G�H�a�[�|��������Jå�ʾ��⨿��}̺Bٺ,��\���*�������G��v������$��*�#�0�77�w&=�
6C��AI�KO�CRU�NV[��Ya��Zg��Zm��Ys�^Xy�rV�a����������D���ũ������L���y��������  �  �i=�=��==F=��=ׂ=� =S� =�[ =��<2*�<�b�<��<���<��<e;�<5o�<���<���<)�<�3�<�a�<\��<���<���<;�<43�<�X�<9|�<?��<e��<���<!��<��<�+�<B�<)V�<�g�<^w�<Y��<��<��</��<Ҟ�<���<���<���<���<���<�q�<_�<sI�<t0�< �<��<���<���<�~�<�P�<^�<i��<���<�p�<v/�<���<���<-S�<��<u��<S�<���<q��</�<�ž<�X�<��<�r�<���<X}�<��<#y�<��<zf�<�ׯ<�E�<i��<��<�{�<�ܧ<�:�<��<[�<�C�<Ж�<%�<5�<���<�ɘ<�<0V�<_��<�ڑ<^�<gX�<�<Њ<�	�<�B�<,z�<̰�<��<��<�|<�y<Mnu<��q<>:n<ߟj<ng<Hkc<~�_<�8\<H�X<C	U<�sQ<&�M<�LJ<-�F<�-C<͡?<j<<ܑ8<T5<�1<+.<�*<�"'<��#<�D <>�<�x<�<2�<�k<�<��<x�<;S<_8�;"��; ��;_<�;|�;m��;��;��;ɮ�;���;���;r�;�J�;Ř�;���;�d�;��;6q�;��;f��;�}�;�L�;dX~;�7t;7j;�V`;��V;�L;�qC;�:;l�0;n�';��;]�;��;);("�:�'�:2b�:��:�r�:�D�:�G�:wy�:��i:A�J:�6,:��:t�9CԤ9�]T9�j�8ݒ�����?�u��Ӳ��O깭���+�dG�z�a���|��������¥�����s���M~̺XBٺ1��Җ��)��2�����G�Uv�ǟ���$���*���0�=7��&=��5C��AI�KO��QU�rV[�0Ya��Zg�bZm��Ys�Xy�sV���������H���6���婎�����N���a��������  �  �i=�=��=@F=��=ׂ=� =P� =�[ =	��<,*�<�b�<��<���<��<f;�<*o�<��<���<2�<�3�<�a�<f��<���<���<<�<(3�<�X�<1|�<7��<V��<���<��<��<�+�<B�<6V�<�g�<^w�<T��<��<Җ�<.��<̞�<���<���<���<���<���<�q�<1_�<lI�<v0�<��<��<���<���<�~�<xP�<a�<`��<���<q�<v/�<��<���<4S�<��<n��<S�<���<g��</�<�ž<�X�<��<�r�<���<a}�<��<%y�<��<rf�<�ׯ<�E�<]��<��<�{�<�ܧ<;�<��<m�<�C�<Ŗ�<,�<5�<���<�ɘ<�<(V�<c��<�ڑ<^�<�X�<<Њ<�	�<�B�<3z�<���<��<��<П|<ty<Qnu<��q<A:n<��j<Mg<ckc<��_<t8\<N�X<#	U<msQ<$�M<�LJ<�F<�-C<ɡ?<i<<�8<G5<4�1<2.<�*<�"'<��#<�D <K�<�x<�<D�<�k<�<��<j�<OS<E8�;0��;��;0<�;o�;M��;��;���;Ѯ�;���;���;��;�J�;���;���;�d�;��;q�;z�;a��;j}�;�L�;�X~;�7t;\7j;�V`;ЕV;��L;�qC;�:;T�0;N�';��;k�;��;�(;\"�:<'�:�c�:���:�r�:�E�:wG�:�y�:��i:Y�J:I6,:��:��9�Ѥ9_T9?i�8�b�����A�u��Ѳ��P�Z����+�|G���a��|�ȉ��/���v¥����ɧ���~̺7Aٺ?�庁��)�����m��G�iv�����$���*���0�z7��&=��5C��AI�LKO��QU��V[�>Ya��Zg��Zm�Zs�mXy��V�����w�����������ש��%���C�������ᴚ��  �  �i=�=��=:F=��=ڂ=� =R� =�[ =��<0*�<�b�<��<���<��<];�<2o�<���<���<0�<~3�<�a�<S��<ƹ�<���<<�</3�<�X�<A|�<5��<j��<���<��<��<�+�< B�<%V�<�g�<]w�<d��<��<ז�<9��<Ȟ�<���<���<���<���<���<~q�<_�<vI�<o0�<�<��<���<���<�~�<~P�<X�<j��<���<�p�<n/�<���<���<)S�<��<k��<S�<���<n��<!/�<�ž<�X�<��<�r�<���<U}�<��<%y�<��<pf�<�ׯ<�E�<a��<��<�{�<�ܧ<�:�<��<Y�<�C�<͖�<#�<5�<���<�ɘ<�<)V�<c��<�ڑ<g�<gX�<�<Њ<�	�<�B�<'z�<̰�<��<��<͟|<�y<bnu<��q<@:n<ޟj<yg<Kkc<��_<u8\<Z�X<F	U<jsQ<E�M<�LJ<)�F<�-C<ʡ?<w<<͑8<O5<�1<@.<�*<�"'<��#<�D <[�<�x<�<2�<�k<�<��<s�<*S<u8�;��;��;I<�;l�;���;��;	��;Ү�;���;���;}�;�J�;���;���;�d�;��;8q�;��;���;Z}�;�L�;KX~;�7t;#7j;VV`;��V;"�L;
rC;y:;y�0;5�';��;��;��;�(;�!�:�'�:gb�:���:r�:�D�:H�:3y�:�i:�J:a7,:�:��9b֤9�^T9=h�8�������u�lԲ��P�]��b�+��G���a�Ô|�����ఘ� å�:���ͨ���~̺pBٺ�����$*��R����{G��v������$���*���0�=7��&=�)6C��AI�9KO�	RU�nV[�iYa�TZg��Zm��Ys�*Xy��V���������1���/���ک��%���+���Z���級��  �  �i=�=��=9F=��=ق=� =f� =�[ =��</*�<�b�<��<���<��<X;�<Do�<���<���<+�<�3�<�a�<N��<˹�<���<>�<53�<�X�<<|�<'��<l��<���<'��<��<�+�<)B�<"V�<�g�<Uw�<S��<ݎ�<͖�<0��<���<���<���<���<���<���<�q�<_�<�I�<k0�<�<��<���<���<�~�<�P�<Y�<w��<���<q�<�/�<���<���<&S�<��<b��<S�<���<\��</�<�ž<�X�<��<�r�<���<Z}�< ��<y�<��<`f�<�ׯ<�E�<`��<��<�{�< ݧ<�:�<7��<c�<�C�<֖�<$�<5�<���<�ɘ<�<2V�<d��<�ڑ<h�<`X�<��<Њ<�	�<�B�<&z�<۰�<y�<��<��|<�y<;nu<��q<Z:n<ğj<�g<*kc<��_<�8\<7�X<G	U<YsQ<6�M<�LJ<B�F<�-C<ɡ?<s<<͑8<�5<��1<<.<�*<�"'<��#<�D <T�<�x<<-�<�k<�<��<��<S<�8�;���;��;d<�;6�;x��;���;��;���;о�;���;[�;�J�;���;���;�d�;��;�p�;h�;k��;.}�;M�;AX~;$8t;
7j;�V`;��V;�L;YrC;^:;��0;&�';��;e�;��;});�!�:�(�:b�:t��:�s�:�D�:�H�:	y�:g�i:��J:�5,:��:@�9PӤ9�YT9lx�8Q������i�u�Ӳ��L깬����+��
G���a���|����������å�����4���c|̺�Aٺ*��s��*��������G��v������$��*�|�0�y7��%=��5C��AI�KO�RU��U[��Ya��Zg�[m��Ys��Xy��V�N���ᩅ����q����������o���Y���	����  �  �i=�=��=:F=��=ڂ=� =R� =�[ =��<0*�<�b�<��<���<��<];�<2o�<���<���<0�<~3�<�a�<S��<ƹ�<���<<�</3�<�X�<A|�<5��<j��<���<��<��<�+�< B�<%V�<�g�<]w�<d��<��<ז�<9��<Ȟ�<���<���<���<���<���<~q�<_�<vI�<o0�<�<��<���<���<�~�<~P�<X�<j��<���<�p�<n/�<���<���<)S�<��<k��<S�<���<n��<!/�<�ž<�X�<��<�r�<���<U}�<��<%y�<��<pf�<�ׯ<�E�<a��<��<�{�<�ܧ<�:�<��<Y�<�C�<͖�<#�<5�<���<�ɘ<�<)V�<c��<�ڑ<g�<gX�<�<Њ<�	�<�B�<'z�<̰�<��<��<͟|<�y<bnu<��q<@:n<ޟj<yg<Kkc<��_<u8\<Z�X<F	U<jsQ<E�M<�LJ<)�F<�-C<ʡ?<w<<͑8<O5<�1<@.<�*<�"'<��#<�D <[�<�x<�<2�<�k<�<��<s�<*S<u8�;��;��;I<�;l�;���;��;	��;Ү�;���;���;}�;�J�;���;���;�d�;��;8q�;��;���;Z}�;�L�;KX~;�7t;#7j;VV`;��V;"�L;
rC;y:;y�0;5�';��;��;��;�(;�!�:�'�:gb�:���:r�:�D�:H�:3y�:�i:�J:a7,:�:��9b֤9�^T9=h�8�������u�lԲ��P�]��b�+��G���a�Ô|�����ఘ� å�:���ͨ���~̺pBٺ�����$*��R����{G��v������$���*���0�=7��&=�)6C��AI�9KO�	RU�nV[�iYa�TZg��Zm��Ys�*Xy��V���������1���/���ک��%���+���Z���級��  �  �i=�=��=@F=��=ׂ=� =P� =�[ =	��<,*�<�b�<��<���<��<f;�<*o�<��<���<2�<�3�<�a�<f��<���<���<<�<(3�<�X�<1|�<7��<V��<���<��<��<�+�<B�<6V�<�g�<^w�<T��<��<Җ�<.��<̞�<���<���<���<���<���<�q�<1_�<lI�<v0�<��<��<���<���<�~�<xP�<a�<`��<���<q�<v/�<��<���<4S�<��<n��<S�<���<g��</�<�ž<�X�<��<�r�<���<a}�<��<%y�<��<rf�<�ׯ<�E�<]��<��<�{�<�ܧ<;�<��<m�<�C�<Ŗ�<,�<5�<���<�ɘ<�<(V�<c��<�ڑ<^�<�X�<<Њ<�	�<�B�<3z�<���<��<��<П|<ty<Qnu<��q<A:n<��j<Mg<ckc<��_<t8\<N�X<#	U<msQ<$�M<�LJ<�F<�-C<ɡ?<i<<�8<G5<4�1<2.<�*<�"'<��#<�D <K�<�x<�<D�<�k<�<��<j�<OS<E8�;0��;��;0<�;o�;M��;��;���;Ѯ�;���;���;��;�J�;���;���;�d�;��;q�;z�;a��;j}�;�L�;�X~;�7t;\7j;�V`;ЕV;��L;�qC;�:;T�0;N�';��;k�;��;�(;\"�:<'�:�c�:���:�r�:�E�:wG�:�y�:��i:Y�J:I6,:��:��9�Ѥ9_T9?i�8�b�����A�u��Ѳ��P�Z����+�|G���a��|�ȉ��/���v¥����ɧ���~̺7Aٺ?�庁��)�����m��G�iv�����$���*���0�z7��&=��5C��AI�LKO��QU��V[�>Ya��Zg��Zm�Zs�mXy��V�����w�����������ש��%���C�������ᴚ��  �  �i=�=��==F=��=ׂ=� =S� =�[ =��<2*�<�b�<��<���<��<e;�<5o�<���<���<)�<�3�<�a�<\��<���<���<;�<43�<�X�<9|�<?��<e��<���<!��<��<�+�<B�<)V�<�g�<^w�<Y��<��<��</��<Ҟ�<���<���<���<���<���<�q�<_�<sI�<t0�< �<��<���<���<�~�<�P�<^�<i��<���<�p�<v/�<���<���<-S�<��<u��<S�<���<q��</�<�ž<�X�<��<�r�<���<X}�<��<#y�<��<zf�<�ׯ<�E�<i��<��<�{�<�ܧ<�:�<��<[�<�C�<Ж�<%�<5�<���<�ɘ<�<0V�<_��<�ڑ<^�<gX�<�<Њ<�	�<�B�<,z�<̰�<��<��<�|<�y<Mnu<��q<>:n<ߟj<ng<Hkc<~�_<�8\<H�X<C	U<�sQ<&�M<�LJ<-�F<�-C<͡?<j<<ܑ8<T5<�1<+.<�*<�"'<��#<�D <>�<�x<�<2�<�k<�<��<x�<;S<_8�;"��; ��;_<�;|�;m��;��;��;ɮ�;���;���;r�;�J�;Ř�;���;�d�;��;6q�;��;f��;�}�;�L�;dX~;�7t;7j;�V`;��V;�L;�qC;�:;l�0;n�';��;]�;��;);("�:�'�:2b�:��:�r�:�D�:�G�:wy�:��i:A�J:�6,:��:t�9CԤ9�]T9�j�8ݒ�����?�u��Ӳ��O깭���+�dG�z�a���|��������¥�����s���M~̺XBٺ1��Җ��)��2�����G�Uv�ǟ���$���*���0�=7��&=��5C��AI�KO��QU�rV[�0Ya��Zg�bZm��Ys�Xy�sV���������H���6���婎�����N���a��������  �  �i=�=��=8F=��=܂=� =X� =�[ =��<.*�<�b�<��<���<��<Y;�<9o�<��<���<:�<�3�<�a�<S��<̹�<���<:�</3�<�X�<=|�<,��<e��<���<"��<��<�+�<%B�<#V�<�g�<Yw�<`��<ߎ�<֖�<+��<Ȟ�<���<���<���<���<���<�q�<_�<�I�<f0�<�<��<���<���<�~�<�P�<O�<x��<���<q�<z/�<���<���<!S�<��<k��<S�<���<`��</�<�ž<�X�<��<�r�<���<Z}�<��<y�<��<ff�<�ׯ<�E�<`��<��<�{�<�ܧ<�:�< ��<_�<�C�<ז�<�<5�<���<�ɘ<
�<2V�<]��<�ڑ<s�<hX�<���<Њ<�	�<�B�< z�<Ѱ�<��<��<Ɵ|<�y<Unu<��q<P:n<ןj<�g<Akc<��_<�8\<J�X<7	U<`sQ<4�M<�LJ<1�F<�-C<С?<�<<͑8<h5<�1<V.<�*<�"'<��#<�D <R�<�x<�<�<�k<<��<��<(S<�8�;��;���;J<�;B�;}��;ǻ�;���;���;���;���;x�;�J�;���;���;�d�;��;q�;��;U��;Y}�;�L�;X~;8t;97j;�V`;�V;?�L;~rC;5:;o�0;W�';͘;q�;��;);<!�:�(�:�b�:���:�r�:�D�:�H�:�x�:�i:�J:�5,:�::�9xդ9�[T9fr�8����?����u�dӲ�jN�5����+��	G�H�a�[�|��������Jå�ʾ��⨿��}̺Bٺ,��\���*�������G��v������$��*�#�0�77�w&=�
6C��AI�KO�CRU�NV[��Ya��Zg��Zm��Ys�^Xy�rV�a����������D���ũ������L���y��������  �  �i=�=��=>F=��=ւ=� =U� =�[ =
��<"*�<�b�<��<���<��<W;�<8o�<��<���<-�<�3�<�a�<Z��<���<���<@�<03�<�X�<B|�<9��<e��<���<��<��<�+�<B�<2V�<�g�<Pw�<^��<��<ۖ�<0��<ɞ�<���<���<���<���<���<�q�<!_�<pI�<k0�<�<��<���<���<�~�<�P�<Y�<c��<���<q�<v/�<���<���<,S�<��<n��<S�<���<h��</�<�ž<�X�<��<�r�<���<c}�<��<y�<��<qf�<�ׯ<�E�<c��<��<�{�<�ܧ<�:�<��<a�<�C�<�<)�<5�<���<�ɘ<
�<0V�<g��<�ڑ<_�<jX�<���<Њ<�	�<�B�</z�<Ͱ�<��<��<՟|<�y<Tnu<o�q<S:n<�j<[g<Rkc<��_<i8\<N�X<;	U<rsQ<?�M<�LJ<.�F<�-C<��?<e<<ߑ8<]5<	�1<4.<��*<�"'<��#<�D <h�<�x<�<C�<�k<�<��<��<8S<W8�;
��;��;N<�;M�;���;���;���;���;���;���;�;�J�;蘯;���;�d�;��;q�;��;j��;_}�;�L�;}X~;�7t;77j;�V`;ЕV;M�L;�qC;^:;��0;E�';ʘ;��;��;6);�!�:o'�:�b�:n��:�r�:9E�:�G�:fy�:��i:`�J:�5,:k�:�9�Ԥ9�XT9�r�8	n�����u��в��O�p���+��G���a��|�u���Ͱ��å�����q���*~̺�Aٺ��庳��)��
����PG��v�ɟ���$�Q�*���0�#7��&=��5C�BI�SKO��QU�iV[��Ya�qZg��Zm��Ys�cXy��V�\�������m���"�������<���C���p���״���  �  �i=�=��=;F=��=ւ=� =Q� =�[ =��<2*�<�b�<��<���<��<`;�<(o�<���<���<4�<�3�<�a�<`��<���<���<7�</3�<�X�<8|�<<��<c��<���<��<��<�+�<!B�<*V�<�g�<^w�<\��<��<ז�<+��<Ԟ�<���<���<���<���<���<~q�<(_�<sI�<u0�<��<��<���<���<�~�<vP�<]�<g��<���<�p�<t/�<��<���<3S�<��<x��<S�<���<m��</�<�ž<�X�<��<�r�<���<Y}�<��<(y�<��<vf�<�ׯ<�E�<g��<��<�{�<�ܧ<;�<��<^�<�C�<̖�<'�<�4�<���<�ɘ<�<'V�<Z��<�ڑ<c�<rX�<<Њ<�	�<�B�<.z�<Ű�<��<��<ן|<�y<Xnu<��q<8:n<�j<wg<Qkc<~�_<x8\<U�X<?	U<vsQ<*�M<�LJ< �F<�-C<ˡ?<e<<�8<L5<�1<>.<�*<�"'<��#<�D <T�<�x<�<7�<�k<<��<r�<CS<S8�;0��;��;I<�;r�;f��;��;��;߮�;���;���;��;�J�;Ƙ�;���;�d�;��;,q�;��;T��;�}�;�L�;�X~;�7t;b7j;�V`;��V;��L;�qC;�:;-�0;E�';�;x�;��;�(;!"�:�'�:c�:��:xr�:�E�:yG�:�y�:��i:��J:�5,:��:a�9Ԥ9�^T9Ue�8������͵u��Ӳ�Q���P�+��G��a�R�|�4���b���{¥�쿲�
����~̺'BٺY�����)��������G�vv����$���*���0��7��&=��5C�BI�<KO��QU��V[�,Ya��Zg��Zm��Ys�SXy��V���������5���$���穎����4���i���Ѵ���  �  �i=�=��=8F=��=ق=� =W� =�[ =��<-*�<�b�<��<���<~�<e;�<5o�<��<���<2�<�3�<�a�<U��<ƹ�<���<6�<+3�<�X�<@|�<4��<_��<���<'��<��<�+�<*B�<&V�<�g�<^w�<T��<��<ܖ�<0��<͞�<���<���<���<���<���<�q�<"_�<uI�<i0�<��<��<���<���<�~�<�P�<Q�<i��<���<q�<s/�<���<���<+S�<��<q��<S�<���<g��</�<�ž<�X�<��<�r�<���<[}�<��<y�<��<nf�<�ׯ<�E�<b��<��<�{�<�ܧ<�:�<��<`�<�C�<̖�<�<5�<���<�ɘ<�<2V�<X��<�ڑ<e�<oX�<���<Њ<�	�<�B�<%z�<ư�<��<��<ן|<~y<=nu<��q<T:n<ϟj<�g<<kc<��_<�8\<6�X<4	U<psQ<;�M<�LJ<!�F<�-C<ڡ?<q<<Б8<b5<�1<;.<�*<�"'<��#<�D <8�<�x<�<�<�k<�<��<��<,S<u8�;-��;��;<<�;e�;���;��;ݭ�;���;Ͼ�;���;o�;�J�;���;���;�d�;��;q�;��;h��;n}�;�L�;YX~;�7t;07j;�V`;ՕV;W�L;�qC;N:;d�0;��';��;E�;��;);b!�:�'�:�b�:p��:`r�:E�:H�:Yy�:x�i:��J:E6,:i�:��9�Ҥ9y]T9u�8���������u��Ҳ��M�m����+��G� �a�i�|�~���;����¥�f�������~̺Bٺ������*��&��m��G�v�����$��*���0��7��&=�6C��AI��JO�RU��V[�ZYa�|Zg��Zm��Ys��Xy�PV�Z���˩�����N�������񪑻s���~���ܴ���  �  �i=�=��=;F=��=ق=� =T� =�[ =��<**�<�b�<��<���<��<Z;�<5o�<���<���<.�<|3�<�a�<U��<ɹ�<���<A�<53�<�X�<D|�<1��<s��<���<��<��<�+�< B�<&V�<�g�<Nw�<i��<��<ۖ�<5��<ƞ�<���<���<���<���<���<�q�<_�<xI�<m0�<�<��<���<���<�~�<�P�<V�<m��<���< q�<q/�<���<���<"S�<��<k��<S�<���<k��<)/�<�ž<�X�<��<�r�<���<]}�<��<y�<��<lf�<�ׯ<�E�<f��<��<�{�<�ܧ<�:�<��<Z�<�C�<Ζ�<$�<5�<���<�ɘ<�<,V�<c��<�ڑ<d�<cX�<���<Њ<�	�<�B�<(z�<԰�<��<��<П|<�y<anu<v�q<X:n<ԟj<ug<Akc<��_<u8\<R�X<S	U<hsQ<E�M<�LJ<<�F<�-C<š?<s<<ϑ8<W5<��1<9.<
�*<�"'<��#<�D <_�<�x<�<:�<�k<�<��<v�<,S<�8�;���;��;c<�;P�;���;ػ�;-��;���;���;���;q�;�J�;���;���;�d�;��;1q�;��;}��;R}�;�L�;)X~;�7t;7j;nV`;��V;	�L;rC;j:;��0;5�';ݘ;��;v�;);�!�:(�:.b�:N��:Br�:�D�:&H�:�x�:��i:��J:�6,:��:��97ؤ9�WT9�r�8
������o�u�}Ҳ�bO�ʫ�2�+�D	G���a���|�I��������å����Ĩ��p~̺fBٺ�����*��&����vG��v�����$�(�*���0�]7��&=�6C��AI�5KO�RU�5V[��Ya�\Zg��Zm�wYs�.Xy��V�R�������9���C�������$���:���A���봚��  �  �i=�=��=;F=��=ق=� =Q� =�[ =��<+*�<�b�<��<���<��<_;�<,o�<���<���<6�<�3�<�a�<_��<Ĺ�<���<=�</3�<�X�<;|�<0��<_��<���<��<��<�+�<B�<.V�<�g�<\w�<`��<ێ�<Ֆ�<.��<˞�<���<���<���<���<���<�q�<-_�<uI�<q0�<��<��<���<���<�~�<{P�<[�<i��<���<q�<}/�<��<���<-S�<��<k��<S�<���<_��</�<�ž<�X�<��<�r�<���<_}�<��<'y�<��<if�<�ׯ<�E�<a��<��<�{�<�ܧ<;�<��<g�<�C�<ǖ�<)�<5�<���<�ɘ<�<(V�<c��<�ڑ<e�<uX�<<Њ<�	�<�B�<*z�<ǰ�<��<��<Ο|<vy<]nu<��q<Q:n<�j<bg<Zkc<��_<8\<U�X<*	U<esQ<2�M<�LJ<$�F<�-C<ӡ?<r<<�8<I5<�1<B.<�*<�"'<��#<�D <K�<�x<�<;�<�k<<��<r�<AS<l8�;��;��;I<�;_�;t��;Ի�;ۭ�;ܮ�;���;���;��;�J�;Ԙ�;���;�d�;��;�p�;��;b��;g}�;�L�;pX~;�7t;a7j;�V`;V;��L;rC;�:;O�0;>�';��;]�;��;�(;�!�:�'�:_c�:���:s�:oE�:�G�:yy�:|�i:
�J:*6,:��:��9�Ԥ9_T9�p�8����J���u�Ҳ�MO�8����+��	G���a���|����������¥�s���&���P~̺�Aٺ8��Y���)��s�����G��v�����$��*���0��7��&=��5C��AI�!KO��QU��V[�JYa��Zg��Zm�Zs�?Xy��V�`�������`�������������4�������𴚻�  �  �i=�=��=;F=��=҂=� =O� =�[ =��<.*�<�b�<��<���<w�<k;�<,o�<���<���<*�<3�<�a�<]��<���<���<6�<13�<�X�<8|�<H��<]��<���<!��<��<�+�<B�<1V�<�g�<cw�<V��<��<��<*��<מ�<���<���<���<���<���<xq�<$_�<gI�<t0�<��<��<���<���<�~�<yP�<^�<]��<���<�p�<x/�<���<���<4S�<��<x��<S�<���<t��</�<�ž<�X�<��<�r�<���<Y}�<��<(y�<��<�f�<�ׯ<�E�<g��<��<�{�<�ܧ<�:�<��<Y�<�C�<Ė�<&�<5�<���<�ɘ<�<.V�<Z��<�ڑ<V�<mX�<锌<Њ<�	�<�B�<.z�<°�<��<��<��|<�y<Inu<��q<;:n<�j<og<Skc<~�_<�8\<G�X<4	U<�sQ<%�M<�LJ< �F<�-C<ݡ?<X<<�8<D5<
�1<".<�*<�"'<��#<�D <*�<�x<�<0�<�k<�<��<r�<<S<;8�;>��;��;T<�;u�;h��;4��;խ�;Ԯ�;���;���;��;�J�;ᘯ;���;�d�;��;:q�;��;S��;�}�;�L�;�X~;�7t;7j;�V`;W�V;d�L;�qC;�:;9�0;��';��;0�;��;�(;."�:'�:�b�:���:�r�:�D�:~G�:�y�:��i:��J:�5,:)�:�9~Ҥ9GaT9�g�8���c��X�u�tӲ��O���*�+��G�M�a�4�|�8���d���N¥�!���n���b~̺{Bٺ��应���)��o��G�%H�Sv�؟�	�$���*��0�7�'=��5C�4BI�
KO��QU��V[��Xa��Zg�%Zm��Ys��Xy�TV���������G������橎�󪑻P���~��������  �  �i=�=��=:F=��=ׂ=� =X� =�[ =��<2*�<�b�<��<���<��<];�<-o�<���<���<8�<3�<�a�<W��<Ź�<���<9�<23�<�X�<9|�<0��<h��<���<#��<��<�+�<&B�<(V�<�g�<Yw�<^��<��<Ԗ�<)��<Ȟ�<���<���<���<���<���<�q�<$_�<{I�<t0�<��<��<���<���<�~�<yP�<]�<p��<���< q�<�/�<���<���<*S�<��<l��<S�<���<c��</�<�ž<�X�<��<�r�<���<W}�<��<!y�<��<jf�<�ׯ<�E�<b��<��<�{�<�ܧ<�:�<#��<[�<�C�<Ӗ�<&�<5�<���<�ɘ<�<(V�<Y��<�ڑ<j�<kX�<���<Њ<�	�<�B�<)z�<ΰ�<��<��<̟|<�y<Wnu<��q<J:n<ܟj<~g<Ekc<��_<�8\<Q�X<=	U<isQ<-�M<�LJ<1�F<�-C<ʡ?<k<<ߑ8<e5<�1<F.<�*<�"'<��#<�D <T�<�x<�<2�<�k<<��<��<1S<s8�;��;���;U<�;:�;i��;Ի�;���;ɮ�;���;���;}�;�J�;���;���;�d�;��;q�;��;N��;Y}�;�L�;YX~;�7t;7j;�V`;̕V;c�L;/rC;�:;=�0;"�';И;f�;��;�(;"�:4(�:c�:H��:*s�:�D�:+H�:=y�:��i:)�J:85,:S�:��9�Ԥ9�\T9l�8Q������u��Ӳ��N�ݪ���+��	G��a�ǖ|��������å�M��������}̺MBٺ�废���)��o�����G��v����$���*�k�0�!7��&=��5C��AI�%KO��QU�eV[��Ya��Zg��Zm��Ys�WXy��V�n�������'���<���ϩ�����<���l���괚��  �  ej=�	=��=}G=�=p�=t"=@� =�] =���<�.�<�g�<���<���<��<�A�<Pv�<l��<w��<u�<.<�<�j�<��<���<(��<8�<�>�<pd�<���<��<���<���<��<�"�<s;�<<R�<�f�< y�<��<���<ˡ�<U��<C��<C��<γ�<=��<��<}��<���<Y��<iw�<Hb�<�I�<�-�<H�<E��<���<F��<Nl�<^:�<��<<��<܍�<�L�<3�<��<�p�<U�<���<�p�<2�<���<IL�<��<pu�<�<ߎ�<��<՘�<.�<���<��<��<	�<^^�<TȬ<)/�<���<�<[P�<ժ�<U�<&W�<D��<���<F�<���<Q٘<��<�c�<]��<��<�%�<�b�<���<�؊<��<�I�<b��<2��<��<V�<��|<�y<�pu<��q<9n<�j<� g<�dc<��_<�.\<�X<9�T<�dQ<��M<_:J<L�F<;C<��?<��;<3w8<)�4<p1<��-<�v*<
 '<?�#<� <״<hO<N�< �<><��<2�<�^<�<���;Ok�;%�;���;ɐ�;Ad�;GE�;�5�;~4�;�B�;�`�;��;9˴;�;Pu�;_�;:`�;1�;���;h;�;���;�Ƀ;�R};4s;�4i;�U_;�U;Z�K;�wB;�9;��/;�&;"�;l�;"�;
G;Hd�:�s�:���:�.�:*ٲ:´�:���:��:]�f:t�G:w):`K:���9%ȟ9ĆJ90j�8�d෎���W~�L ���V�Y���-�|�H��c��B~��X���v��J���ou��*X���%ͺ��ٺ9���)����8�)R�?��������H�$�}+��*1��>7��M=��ZC��cI�xjO��nU�qp[��qa��ng�Amm��is�fy�6b�殂���� ������}�����������_���ȯ���  �  Tj=�	=��=}G=�=j�=u"=>� =�] =���</�<�g�<���<���<��<B�<<v�<j��<���<}�<8<�<�j�<��<���<0��<6�<�>�<vd�<���<��<���<���<��<�"�<t;�<7R�<�f�<!y�<��<���<ġ�<8��<-��<_��<̳�<F��<��<w��<���<\��<yw�<Pb�<�I�<�-�<E�<@��<���<G��<:l�<i:�<��<L��<��<�L�<0�<��<�p�<R�<���<�p�<�<���<DL�<��<ru�< �<܎�<��<ᘷ<2�<ȓ�<��<��<��<]^�<hȬ<&/�<���<
�<^P�<ժ�<_�<2W�<T��<���<�E�<���<A٘<��<�c�<O��<��<�%�<�b�<���<�؊<��<�I�<e��<3��<�<6�<[�|<|y<�pu<�q<#9n<�j<� g<ec<��_<�.\<�X<(�T<�dQ<��M<�:J<X�F<=C<��?<��;<7w8<!�4<(p1<��-<�v*<��&<"�#<� <��<uO<&�<��<5><��<F�<�^<�<Q��;ok�;�;��;��;�c�;)E�;�5�;�4�;C�;�`�;��;(˴;F�;Vu�;��;3`�;�;��;;�;F��;�Ƀ;@S};�3s;�4i;�U_;�U;��K;4xB;9;��/; �&;��;(�;#�;hF;�d�:$t�:���:0/�:Kٲ:���:/��:���:��f:��G:u):rG:���9�Ɵ9�J9Bl�8S.���W~�/����U�����-�>�H��c��B~�~W���v��ց��>v���W���%ͺS�ٺy��)�ܵ�����Q�ă���������$��+�b*1�!>7��M=��ZC��cI�ojO��nU�ip[��pa��og��mm��is�fy��a�ۮ��鬅�B������n��������������������  �  Uj=�	=��=zG=�=j�=|"=6� =�] =|��</�<�g�<���<���<��<B�<:v�<o��<���<m�<1<�<�j�<���<���<?��<(�<�>�<}d�<���<1��<���<���<��<�"�<o;�<0R�<�f�<y�<$��<���<ѡ�<P��<.��<h��<���<N��<��<|��<���<H��<qw�<=b�<�I�<�-�<V�<C��<���<Y��<7l�<s:�<��<A��<Ѝ�<�L�<8�<��<�p�<>�<���<�p�<&�<ı�<<L�<��<du�<�<Վ�<��<ژ�<%�<̓�<��<.��<��<a^�<cȬ</�<���<�<kP�<Ǫ�<S�<"W�<H��<���<�E�<Ր�<:٘<��<�c�<M��<��<�%�<�b�<���<�؊<��<�I�<b��< ��<�<5�<��|<�y<�pu<�q<9n<�j<� g<ec<��_<�.\<��X<*�T<�dQ<��M<�:J<:�F<.C<��?<�;<Rw8<�4<!p1<��-<�v*<��&<(�#<� <��<�O<"�<�<,><��<7�<�^<	 <@��;�k�;��;���;���;�c�;�E�;x5�;�4�;�B�;�`�;��;˴;M�;!u�;��;`�;H�;x��;;�;i��;�Ƀ;S};�3s;�4i;�U_;�U;��K;�wB;`9;��/;��&;�; �;��;UF;�e�:�r�:��:�-�:�ز:��:��:j��:p�f:X�G:4u):�I:f��9�ğ98�J9�^�8{1෍���Y~������X�o��!�-���H�j�c�;B~��W���w��Ӏ��mv��(W��b&ͺ�ٺn�溺)�~�����JQ����'�������$��+��*1�A>7�uN=�YZC��cI�]jO��nU�q[��pa��og��lm��is�Pfy��a����嬅�f������������������|��������  �  Yj=�	=��=}G=�=g�={"=:� =�] =���<�.�<�g�<���<���<��<B�<8v�<s��<��<{�<><�<�j�<��<���<9��<1�<�>�<ud�<���<��<���<���<��<�"�<r;�<9R�<�f�<y�<��<���<���<K��<0��<Y��<ų�<P��<��<{��<���<V��<~w�<Bb�<�I�<�-�<F�<C��<���<G��<:l�<q:�<��<N��<ߍ�<�L�<6�<��<�p�<M�<���<�p�<#�<���<=L�<��<ou�<�<ݎ�<��<ݘ�</�<͓�<��<��<��<\^�<aȬ<"/�<���<�<hP�<˪�<c�<1W�<H��<���<�E�<���<C٘<��<�c�<Q��<��<�%�<�b�<���<�؊<��<�I�<i��<-��<�<=�<}�|<dy<�pu<�q<!9n<�j<� g<ec<��_<�.\<�X<�T<�dQ<��M<~:J<M�F<<C<��?<u�;<Mw8<�4<8p1<��-<�v*<  '<�#<� <��<zO<�<�<#><��<Q�<�^< <2��;�k�;�;���;ސ�;�c�;EE�;f5�;�4�;C�;�`�;��;-˴;G�;Pu�;��;`�;��;b��;;�;/��;�Ƀ;�S};�3s;�4i;�U_;�U;�K;�wB;A9;��/;�&;�;H�;)�;mF;ue�:Ws�:���:�.�:ٲ:���:���:O��:[�f:�G:Ku):�I:���9Kş9~�J9Ji�8�:෕���W~�U����V�E����-���H�$�c��B~��W��<w��,����v��_W�� &ͺ�ٺ��溺)�G������Q����n�������$��+��*1��=7� N=�rZC��cI��jO��nU��p[�qa��og�Smm�Fjs�-fy��a�߮��⬅�H���
���s���������������ȯ���  �  \j=�	=��={G=�=k�=x"=<� =�] =���<�.�<�g�<���<���<��<B�<Cv�<p��<��<s�<1<�<�j�<��<���<2��</�<�>�<pd�<���<��<���<���<��<�"�<i;�<;R�<�f�<%y�<��<���<ǡ�<G��<3��<W��<ȳ�<F��<��<y��<���<V��<lw�<Fb�<�I�<�-�<E�<E��<���<E��<Gl�<l:�<��<>��<܍�<�L�<3�<��<�p�<P�<���<�p�<!�<���<RL�<��<ru�<�<ߎ�<��<٘�<.�<Ó�<��<��<��<Y^�<dȬ<!/�<���<�<bP�<Ѫ�<X�<$W�<K��<���<F�<���<L٘<��<�c�<V��<��<�%�<�b�<���<�؊<��<�I�<b��<0��<
�<B�<m�|<�y<�pu<��q<*9n<�j<� g<�dc<��_<�.\<�X<9�T<�dQ<��M<q:J<S�F<2C<��?<��;<Aw8<�4<p1<��-<�v*<  '<+�#<� <ȴ<pO<6�<�<"><��<8�<�^<�<W��;vk�;�;
��;Ȑ�;�c�;?E�;�5�;�4�;�B�;�`�;���;7˴;�;fu�;h�;e`�;!�;S��;,;�;'��;�Ƀ;>S};4s;�4i;�U_;�U;w�K;�wB;9;E�/;�&;#�;v�;�;�F;(e�:�s�:���:�.�:�ز:ʹ�:Y��:���:��f:��G:�u):WI:=��9Wʟ96�J9�l�8\����Z~�J����V����-���H��c�2C~��W��Bw������%v���W���%ͺ��ٺZ�溉)󺅵����R�l��{�������$��+��*1�i>7� N=��ZC��cI�gjO��nU��p[�:qa�|og��mm��is��ey�Pb�ͮ�����;���3���j�������|���`���௚��  �  Xj=�	=��={G=�=h�=z"=<� =�] =���</�<�g�<���<���<��<B�<@v�<i��<���<v�<:<�<�j�<��<���<:��<+�<�>�<sd�<���< ��<���<���<��<�"�<n;�<?R�<�f�<%y�<��<���<���<K��<-��<a��<���<J��<��<y��< ��<Y��<sw�<Jb�<�I�<�-�<M�<>��<���<N��<=l�<j:�<��<D��<��<�L�<5�<��<�p�<E�<���<�p�<$�<���<<L�<��<tu�<�<⎺<��<ט�</�<Ɠ�<��<��<��<W^�<bȬ</�<���<�<aP�<Ӫ�<`�<'W�<S��<���<�E�<Ȑ�<?٘<��<�c�<M��<��<�%�<�b�<���<�؊<��<�I�<a��<(��<�<<�<|�|<qy<�pu<�q<(9n<��j<� g<�dc<��_<�.\<۔X<�T<�dQ<��M<�:J<I�F<2C<��?<x�;<Iw8<�4<%p1<��-<�v*<��&<4�#<� <��<�O</�<��<6><��<J�<�^<�<E��;�k�;��;��;Ԑ�;�c�;bE�;v5�;�4�;C�;�`�;��;I˴;�;fu�;��;`�;�;e��;;�;M��;�Ƀ;aS};�3s;�4i;�U_;�U;��K;xB;9;��/;A�&;�;%�;^�;�F;e�:�s�:��: /�:Nٲ:ᴢ:��:,��:h�f:g�G:�t):�I:���9�ğ9Z�J9�n�8l`�����X~�����vV�,��;�-���H� �c�vC~��W���w��
���hv���W���%ͺF�ٺ(��)�������Q�̃�s�������$��+��*1�G>7�N=�iZC� dI�fjO��nU��p[��pa��og�Tmm�js�Pfy��a�Ю�����#���%���q��������������������  �  Rj=�	=��=�G=�=h�={"=6� =�] =���<	/�<�g�<���<���<��<	B�<:v�<y��<���<r�<<<�<�j�<��<���<A��<1�<�>�<xd�<���<!��<���<���<��<�"�<p;�<5R�<�f�<y�<'��<���<���<P��<(��<a��<���<X��<��<}��<���<T��<vw�<Bb�<�I�<�-�<H�<C��<���<H��<<l�<z:�<��<G��<ߍ�<�L�<8�<��<�p�<B�<���<�p�<'�<���<AL�<��<iu�<�<ڎ�<��<ؘ�<*�<Փ�<��<��<��<]^�<dȬ</�<���<�<hP�<ƪ�<b�<&W�<N��<���<�E�<���<C٘<��<�c�<U��<��<�%�<�b�<���<�؊<��<�I�<n��<&��<�<1�<��|<jy<�pu<!�q<9n<��j<� g<�dc<��_<�.\<��X<�T<�dQ<��M<�:J<>�F<HC<��?<y�;<Mw8< �4<,p1<��-<�v*< '<"�#<� <��<~O<$�<�<4><��<M�<�^< <>��;�k�;	�;��;��;�c�;eE�;k5�;�4�;C�;�`�;��; ˴;&�;:u�;��;+`�;�;v��;�:�;N��;�Ƀ;�S};�3s;�4i;�U_;ݖU;��K;�wB;�9;��/;�&;�;E�;3�;yF;f�:~s�:H��:�.�:�ز:��:���:���:�f:��G:�t):J:h��99Ɵ9�J9Bd�8OY����X~������W�:��e�-���H��c��B~��W���w�������v��UW��z&ͺ$�ٺ:��U)�ִ�����Q����i�������$��+��*1�>7�]N=�iZC��cI�[jO�_nU��p[��pa�pg�2mm�.js��ey��a�����󬅻\��� �������u���y������������  �  Zj=�	=��=~G=�=k�=y"=;� =�] =���<�.�<�g�<���<���<��<B�<Fv�<n��<~��<t�<7<�<�j�<��<���<3��<1�<�>�<yd�<���<��<���<���<��<�"�<m;�<1R�<�f�<y�<��<���<���<N��<3��<[��<���<O��<߫�<z��<���<X��<tw�<Bb�<�I�<�-�<H�<F��<���<H��<Fl�<m:�<��<C��<ލ�<�L�<5�<��<�p�<I�<���<�p�<&�<���<HL�<��<lu�<�<׎�<��<ܘ�<(�<Ǔ�<��<��<��<_^�<_Ȭ<!/�<���<�<iP�<ͪ�<]�<&W�<G��<���<F�<���<O٘<��<�c�<S��<��<�%�<�b�<���<�؊<��<�I�<h��<'��<�<@�<��|<ty<�pu<�q<9n<�j<� g<ec<��_<�.\<�X< �T<�dQ<��M<�:J<?�F<@C<��?<��;<Hw8<�4<%p1<��-<�v*<  '</�#<� <д<rO<;�<�<!><��<D�<�^< <D��;{k�;	�;���;��;�c�;OE�;�5�;�4�;�B�;�`�;��;˴;@�;Iu�;��;@`�;�;m��;-;�;6��;�Ƀ;�S};�3s;�4i;�U_;�U;��K;�wB;#9;5�/;�&;)�;u�;.�;�F;9e�:Gs�:��:�.�:�ز:㴢:���:?��:��f:I�G:�u):�I:���9ȟ9��J9f�8�Aෙ��D[~�|���?X���_�-�?�H��c�xB~�X��Hw��n����v��GW��&ͺm�ٺ4���)󺤵����R�Q��z�������$�+��*1�)>7�N=��ZC��cI��jO��nU��p[�
qa��og�<mm�js�fy�b�宂�ଅ�g������s��������������������  �  Yj=�	=��={G=�=m�=t"=?� =�] =���</�<�g�<���<���<��<B�<Gv�<a��<���<�<0<�<�j�<��<���<4��<1�<�>�<rd�<���<��<���<���<��<�"�<n;�<=R�<�f�<%y�<��<���<���<F��<1��<[��<Ƴ�<E��<��<|��<���<Y��<pw�<Vb�<�I�<�-�<I�<B��<���<I��<Cl�<c:�<��<D��<ݍ�<�L�<3�<��<�p�<N�<���<�p�<!�<���<BL�<��<uu�<�<⎺<��<՘�<2�<œ�<��<��<��<X^�<`Ȭ<#/�<���<�<]P�<Ӫ�<X�</W�<\��<���<F�<���<J٘<��<�c�<M��<��<�%�<�b�<���<�؊<��<�I�<a��<+��<�<@�<q�|<oy<�pu<�q<#9n<�j<� g<�dc<��_<�.\<۔X<�T<�dQ<��M<:J<I�F<5C<��?<��;<3w8<&�4<p1<��-<�v*<��&<5�#<� <Ŵ<uO<>�<�<E><��<6�<�^<�<g��;}k�;�; ��;Ґ�;�c�;@E�;�5�;�4�;C�;�`�;��;A˴;�;fu�;��;&`�;��;Q��;%;�;8��;�Ƀ;:S};�3s;�4i;�U_;�U;��K;`xB;�9;$�/;#�&;�;S�;6�;�F;�d�:�t�:��:�.�:4ٲ:ʹ�:l��:���:z�f:!�G:u):[I:F��9�Ɵ9&�J9�o�8nj����X~�- ���U�D����-�
�H�>�c�IC~��W��"w�������u��X���%ͺ��ٺ���~(�e���}� R�u����������$��+�%*1�p>7��M=��ZC��cI�|jO��nU��p[�qa��og��mm�js�Wfy��a�ۮ�����2���+���z���������������د���  �  Vj=�	=��=|G=�=k�=x"=<� =�] =���</�<�g�<���<���<��<B�<Bv�<r��<���<m�<8<�<�j�<��<���<;��<*�<�>�<wd�<���<+��<���<���<��<�"�<o;�<5R�<�f�<y�<��<���<ˡ�<P��<-��<_��<���<N��<��<z��<���<W��<nw�<@b�<�I�<�-�<N�<F��<���<P��<Al�<r:�<��<@��<ݍ�<�L�<4�<��<�p�<C�<���<�p�<'�<���<>L�<��<gu�<�<ێ�<��<Ԙ�<'�<ʓ�<��<%��<��<\^�<bȬ</�<���<�<`P�<Ϫ�<]�< W�<J��<���<F�<ɐ�<H٘<��<�c�<R��<��<�%�<�b�<���<�؊<��<�I�<f��<"��<�<8�<��|<|y<�pu<�q<9n<��j<� g<�dc<|�_<�.\<�X<$�T<�dQ<��M<�:J<9�F<6C<��?<��;<Aw8<�4<p1<��-<�v*<��&<3�#<� <��<�O<2�<�<)><��<E�<�^<�<[��;�k�;��;���;��;�c�;�E�;}5�;�4�;�B�;�`�;
��;!˴;�;0u�;��;`�;2�;v��;;�;G��;�Ƀ;~S};�3s;�4i;�U_;��U;��K;�wB;U9;%�/;H�&;(�;U�;o�;�F;�e�:Vs�:ض�:�.�:&ٲ:ٴ�:I��:L��:�f:n�G:�t):J:;��9iş9ΏJ9b�8\a෉��Y~�� ��VX��,�-���H�[�c��B~��W���w�� ���)v���W���%ͺp�ٺ��溛)�[������Q����Z�������$��+��*1�`>7��M=��ZC��cI�fjO��nU��p[��pa��og�mm��is�Hfy��a��������X���������������������������  �  Sj=�	=��=�G=�=g�=~"=8� =�] =���<�.�<�g�<���<���<��<B�<7v�<w��<~��<�<C<�<�j�<���<���<5��<0�<�>�<yd�<���<��<���<���<��<�"�<v;�<-R�<�f�<y�<��<���<���<@��<)��<c��<³�<S��<ܫ�<}��<��<W��<�w�<Cb�<�I�<�-�<M�<@��<���<Q��<7l�<v:�<��<W��<ߍ�<�L�<<�<޽�<�p�<J�<���<�p�<�<���<8L�<��<eu�<&�<Վ�<��<☷<$�<ϓ�<��<��<��<\^�<bȬ</�<���<��<pP�<̪�<d�<5W�<H��<���<�E�<ʐ�<?٘<��<�c�<P��<��<�%�<�b�<���<�؊<��<�I�<m��<&��<�<3�<t�|<`y<�pu<�q<9n<�j<� g<ec<��_<�.\<�X<�T<�dQ<��M<�:J<C�F<GC<��?<u�;<Zw8<�4<Ap1<��-<�v*< '<&�#<� <��<�O<�<�<"><��<\�<�^< <"��;�k�;�;��;��;�c�;VE�;W5�;�4�;�B�;�`�;$��;�ʴ;s�;(u�;��;`�;��;8��;;�;V��;�Ƀ;�S};�3s;�4i;�U_;��U;N�K;�wB;Y9;��/;A�&;��;�;|�;TF;�e�:Es�:O��:�.�:2ٲ:T��:Y��:���:��f:��G:�t):H:���9ğ98�J9�_�8U෫���W~�����Y����-�b�H���c��B~��W��pw��5���0w���V��&ͺ�ٺ?�溿)�������Q�у�l�������$��+��*1��=7�'N=�<ZC�dI��jO�dnU��p[��pa��og�wmm�Sjs�fy��a�������������㩋�����������������ů���  �  Zj=�	=��={G=�=n�=y"=7� =�] =���< /�<�g�<���<���<��<B�<Bv�<s��<���<z�<&<�<�j�<��<���<6��<0�<�>�<qd�<���<"��<���<���<��<�"�<l;�<2R�<�f�<y�<��<���<̡�<N��<5��<W��<ų�<B��<��<���<���<G��<mw�<Kb�<�I�<�-�<R�<F��<���<S��<Dl�<o:�<��<B��<͍�<�L�<9�<��<�p�<L�<���<�p�<*�<���<JL�<��<hu�<�<׎�<��<Ԙ�<'�<Ó�<��<��<��<[^�<^Ȭ< /�<���<�<fP�<˪�<J�<+W�<P��<���<F�<Ȑ�<G٘<��<�c�<X��<��<�%�<�b�<���<�؊<��<�I�<_��<*��<�<A�<��|<�y<�pu<�q<9n<�j<� g<�dc<��_<�.\<�X<,�T<�dQ<��M<t:J<H�F<4C<��?<��;<Fw8<�4<p1<��-<�v*< '<4�#<� <��<�O<4�<�<3><��<#�<�^<�<v��;�k�;�;���;А�;d�;hE�;�5�;�4�;�B�;�`�;���;˴;!�;8u�;��;G`�;5�;q��;2;�;$��;�Ƀ; S};4s;�4i;�U_;x�U;|�K;xB;-9;>�/;l�&;.�;W�;��;�F;`e�:�s�:���:�-�:ٲ:$��:��:���:7�f:��G:�u):cJ:��9�ȟ9a�J9�b�8�_�`��vZ~�� ��_X�m��}�-���H���c�C~�X��Tw��}����u��xW��%&ͺ��ٺލ�8)�[������Q����N�����p�$��+�n*1��>7�cN=��ZC��cI�AjO��nU��p[�/qa��og�Gmm��is�fy�b��������e���.���������������z��������  �  \j=�	=��=xG=�=j�=q"=H� =�] =���<�.�<�g�<���<���<��<B�<@v�<e��<���<~�<;<�<�j�<ԗ�<���<1��<0�<�>�<nd�<���<��<���<���<��<�"�<m;�<@R�<�f�<.y�<��<���<���<E��<4��<U��<г�<:��<��<j��<��<h��<tw�<Sb�<�I�<�-�<E�<F��<���<E��<Bl�<_:�<��<I��<��<�L�< �<���<�p�<S�<���<�p�< �<���<AL�<��<|u�<�<⎺<��<ט�<:�<���<��<��<��<W^�<eȬ<"/�<���<�<JP�<䪤<e�<1W�<Q��<���< F�<���<L٘<��<�c�<O��<��<�%�<�b�<���<�؊<��<�I�<W��<7��<�<C�<j�|<ry<tpu<�q<;9n<�j<� g<�dc<��_<�.\<ŔX<�T<�dQ<��M<q:J<`�F<&C<��?<�;<(w8<K�4<p1<��-<�v*<��&<*�#<� <Ѵ<qO<1�<�<3><��<M�<�^<�<w��;rk�;�;��;Ð�;d�;(E�;|5�;S4�;/C�;�`�;���;M˴;�;�u�;v�;`�;��;J��;1;�;��; ʃ;�R};84s;14i; V_;~�U;��K;LxB;�9;(�/;�&;+�;j�;�;�F;jd�:+t�:p��:�/�:�ٲ:���:���:��:)�f:��G:�u):4I:��9"Ɵ9��J9Hw�83g�L��Y~������S����-���H�ӥc�iC~��W��.w������u��:Y���$ͺ��ٺ���-)�a�����R�f��U�������$�#+�*1�c>7�RM=��ZC�dI�6jO�oU�Hp[�Bqa�tog��mm�js��fy��a�����������?���P�������ت������쯚��  �  Zj=�	=��={G=�=n�=y"=7� =�] =���< /�<�g�<���<���<��<B�<Bv�<s��<���<z�<&<�<�j�<��<���<6��<0�<�>�<qd�<���<"��<���<���<��<�"�<l;�<2R�<�f�<y�<��<���<̡�<N��<5��<W��<ų�<B��<��<���<���<G��<mw�<Kb�<�I�<�-�<R�<F��<���<S��<Dl�<o:�<��<B��<͍�<�L�<9�<��<�p�<L�<���<�p�<*�<���<JL�<��<hu�<�<׎�<��<Ԙ�<'�<Ó�<��<��<��<[^�<^Ȭ< /�<���<�<fP�<˪�<J�<+W�<P��<���<F�<Ȑ�<G٘<��<�c�<X��<��<�%�<�b�<���<�؊<��<�I�<_��<*��<�<A�<��|<�y<�pu<�q<9n<�j<� g<�dc<��_<�.\<�X<,�T<�dQ<��M<t:J<H�F<4C<��?<��;<Fw8<�4<p1<��-<�v*< '<4�#<� <��<�O<4�<�<3><��<#�<�^<�<v��;�k�;�;���;А�;d�;hE�;�5�;�4�;�B�;�`�;���;˴;!�;8u�;��;G`�;5�;q��;2;�;$��;�Ƀ; S};4s;�4i;�U_;x�U;|�K;xB;-9;>�/;l�&;.�;W�;��;�F;`e�:�s�:���:�-�:ٲ:$��:��:���:7�f:��G:�u):cJ:��9�ȟ9a�J9�b�8�_�`��vZ~�� ��_X�m��}�-���H���c�C~�X��Tw��}����u��xW��%&ͺ��ٺލ�8)�[������Q����N�����p�$��+�n*1��>7�cN=��ZC��cI�AjO��nU��p[�/qa��og�Gmm��is�fy�b��������e���.���������������z��������  �  Sj=�	=��=�G=�=g�=~"=8� =�] =���<�.�<�g�<���<���<��<B�<7v�<w��<~��<�<C<�<�j�<���<���<5��<0�<�>�<yd�<���<��<���<���<��<�"�<v;�<-R�<�f�<y�<��<���<���<@��<)��<c��<³�<S��<ܫ�<}��<��<W��<�w�<Cb�<�I�<�-�<M�<@��<���<Q��<7l�<v:�<��<W��<ߍ�<�L�<<�<޽�<�p�<J�<���<�p�<�<���<8L�<��<eu�<&�<Վ�<��<☷<$�<ϓ�<��<��<��<\^�<bȬ</�<���<��<pP�<̪�<d�<5W�<H��<���<�E�<ʐ�<?٘<��<�c�<P��<��<�%�<�b�<���<�؊<��<�I�<m��<&��<�<3�<t�|<`y<�pu<�q<9n<�j<� g<ec<��_<�.\<�X<�T<�dQ<��M<�:J<C�F<GC<��?<u�;<Zw8<�4<Ap1<��-<�v*< '<&�#<� <��<�O<�<�<"><��<\�<�^< <"��;�k�;�;��;��;�c�;VE�;W5�;�4�;�B�;�`�;$��;�ʴ;s�;(u�;��;`�;��;8��;;�;V��;�Ƀ;�S};�3s;�4i;�U_;��U;N�K;�wB;Y9;��/;A�&;��;�;|�;TF;�e�:Es�:O��:�.�:2ٲ:T��:Y��:���:��f:��G:�t):H:���9ğ98�J9�_�8U෫���W~�����Y����-�b�H���c��B~��W��pw��5���0w���V��&ͺ�ٺ?�溿)�������Q�у�l�������$��+��*1��=7�'N=�<ZC�dI��jO�dnU��p[��pa��og�wmm�Sjs�fy��a�������������㩋�����������������ů���  �  Vj=�	=��=|G=�=k�=x"=<� =�] =���</�<�g�<���<���<��<B�<Bv�<r��<���<m�<8<�<�j�<��<���<;��<*�<�>�<wd�<���<+��<���<���<��<�"�<o;�<5R�<�f�<y�<��<���<ˡ�<P��<-��<_��<���<N��<��<z��<���<W��<nw�<@b�<�I�<�-�<N�<F��<���<P��<Al�<r:�<��<@��<ݍ�<�L�<4�<��<�p�<C�<���<�p�<'�<���<>L�<��<gu�<�<ێ�<��<Ԙ�<'�<ʓ�<��<%��<��<\^�<bȬ</�<���<�<`P�<Ϫ�<]�< W�<J��<���<F�<ɐ�<H٘<��<�c�<R��<��<�%�<�b�<���<�؊<��<�I�<f��<"��<�<8�<��|<|y<�pu<�q<9n<��j<� g<�dc<|�_<�.\<�X<$�T<�dQ<��M<�:J<9�F<6C<��?<��;<Aw8<�4<p1<��-<�v*<��&<3�#<� <��<�O<2�<�<)><��<E�<�^<�<[��;�k�;��;���;��;�c�;�E�;}5�;�4�;�B�;�`�;
��;!˴;�;0u�;��;`�;2�;v��;;�;G��;�Ƀ;~S};�3s;�4i;�U_;��U;��K;�wB;U9;%�/;H�&;(�;U�;o�;�F;�e�:Vs�:ض�:�.�:&ٲ:ٴ�:I��:L��:�f:n�G:�t):J:;��9iş9ΏJ9b�8\a෉��Y~�� ��VX��,�-���H�[�c��B~��W���w�� ���)v���W���%ͺp�ٺ��溛)�[������Q����Z�������$��+��*1�`>7��M=��ZC��cI�fjO��nU��p[��pa��og�mm��is�Hfy��a��������X���������������������������  �  Yj=�	=��={G=�=m�=t"=?� =�] =���</�<�g�<���<���<��<B�<Gv�<a��<���<�<0<�<�j�<��<���<4��<1�<�>�<rd�<���<��<���<���<��<�"�<n;�<=R�<�f�<%y�<��<���<���<F��<1��<[��<Ƴ�<E��<��<|��<���<Y��<pw�<Vb�<�I�<�-�<I�<B��<���<I��<Cl�<c:�<��<D��<ݍ�<�L�<3�<��<�p�<N�<���<�p�<!�<���<BL�<��<uu�<�<⎺<��<՘�<2�<œ�<��<��<��<X^�<`Ȭ<#/�<���<�<]P�<Ӫ�<X�</W�<\��<���<F�<���<J٘<��<�c�<M��<��<�%�<�b�<���<�؊<��<�I�<a��<+��<�<@�<q�|<oy<�pu<�q<#9n<�j<� g<�dc<��_<�.\<۔X<�T<�dQ<��M<:J<I�F<5C<��?<��;<3w8<&�4<p1<��-<�v*<��&<5�#<� <Ŵ<uO<>�<�<E><��<6�<�^<�<g��;}k�;�; ��;Ґ�;�c�;@E�;�5�;�4�;C�;�`�;��;A˴;�;fu�;��;&`�;��;Q��;%;�;8��;�Ƀ;:S};�3s;�4i;�U_;�U;��K;`xB;�9;$�/;#�&;�;S�;6�;�F;�d�:�t�:��:�.�:4ٲ:ʹ�:l��:���:z�f:!�G:u):[I:F��9�Ɵ9&�J9�o�8nj����X~�- ���U�D����-�
�H�>�c�IC~��W��"w�������u��X���%ͺ��ٺ���~(�e���}� R�u����������$��+�%*1�p>7��M=��ZC��cI�|jO��nU��p[�qa��og��mm�js�Wfy��a�ۮ�����2���+���z���������������د���  �  Zj=�	=��=~G=�=k�=y"=;� =�] =���<�.�<�g�<���<���<��<B�<Fv�<n��<~��<t�<7<�<�j�<��<���<3��<1�<�>�<yd�<���<��<���<���<��<�"�<m;�<1R�<�f�<y�<��<���<���<N��<3��<[��<���<O��<߫�<z��<���<X��<tw�<Bb�<�I�<�-�<H�<F��<���<H��<Fl�<m:�<��<C��<ލ�<�L�<5�<��<�p�<I�<���<�p�<&�<���<HL�<��<lu�<�<׎�<��<ܘ�<(�<Ǔ�<��<��<��<_^�<_Ȭ<!/�<���<�<iP�<ͪ�<]�<&W�<G��<���<F�<���<O٘<��<�c�<S��<��<�%�<�b�<���<�؊<��<�I�<h��<'��<�<@�<��|<ty<�pu<�q<9n<�j<� g<ec<��_<�.\<�X< �T<�dQ<��M<�:J<?�F<@C<��?<��;<Hw8<�4<%p1<��-<�v*<  '</�#<� <д<rO<;�<�<!><��<D�<�^< <D��;{k�;	�;���;��;�c�;OE�;�5�;�4�;�B�;�`�;��;˴;@�;Iu�;��;@`�;�;m��;-;�;6��;�Ƀ;�S};�3s;�4i;�U_;�U;��K;�wB;#9;5�/;�&;)�;u�;.�;�F;9e�:Gs�:��:�.�:�ز:㴢:���:?��:��f:I�G:�u):�I:���9ȟ9��J9f�8�Aෙ��D[~�|���?X���_�-�?�H��c�xB~�X��Hw��n����v��GW��&ͺm�ٺ4���)󺤵����R�Q��z�������$�+��*1�)>7�N=��ZC��cI��jO��nU��p[�
qa��og�<mm�js�fy�b�宂�ଅ�g������s��������������������  �  Rj=�	=��=�G=�=h�={"=6� =�] =���<	/�<�g�<���<���<��<	B�<:v�<y��<���<r�<<<�<�j�<��<���<A��<1�<�>�<xd�<���<!��<���<���<��<�"�<p;�<5R�<�f�<y�<'��<���<���<P��<(��<a��<���<X��<��<}��<���<T��<vw�<Bb�<�I�<�-�<H�<C��<���<H��<<l�<z:�<��<G��<ߍ�<�L�<8�<��<�p�<B�<���<�p�<'�<���<AL�<��<iu�<�<ڎ�<��<ؘ�<*�<Փ�<��<��<��<]^�<dȬ</�<���<�<hP�<ƪ�<b�<&W�<N��<���<�E�<���<C٘<��<�c�<U��<��<�%�<�b�<���<�؊<��<�I�<n��<&��<�<1�<��|<jy<�pu<!�q<9n<��j<� g<�dc<��_<�.\<��X<�T<�dQ<��M<�:J<>�F<HC<��?<y�;<Mw8< �4<,p1<��-<�v*< '<"�#<� <��<~O<$�<�<4><��<M�<�^< <>��;�k�;	�;��;��;�c�;eE�;k5�;�4�;C�;�`�;��; ˴;&�;:u�;��;+`�;�;v��;�:�;N��;�Ƀ;�S};�3s;�4i;�U_;ݖU;��K;�wB;�9;��/;�&;�;E�;3�;yF;f�:~s�:H��:�.�:�ز:��:���:���:�f:��G:�t):J:h��99Ɵ9�J9Bd�8OY����X~������W�:��e�-���H��c��B~��W���w�������v��UW��z&ͺ$�ٺ:��U)�ִ�����Q����i�������$��+��*1�>7�]N=�iZC��cI�[jO�_nU��p[��pa�pg�2mm�.js��ey��a�����󬅻\��� �������u���y������������  �  Xj=�	=��={G=�=h�=z"=<� =�] =���</�<�g�<���<���<��<B�<@v�<i��<���<v�<:<�<�j�<��<���<:��<+�<�>�<sd�<���< ��<���<���<��<�"�<n;�<?R�<�f�<%y�<��<���<���<K��<-��<a��<���<J��<��<y��< ��<Y��<sw�<Jb�<�I�<�-�<M�<>��<���<N��<=l�<j:�<��<D��<��<�L�<5�<��<�p�<E�<���<�p�<$�<���<<L�<��<tu�<�<⎺<��<ט�</�<Ɠ�<��<��<��<W^�<bȬ</�<���<�<aP�<Ӫ�<`�<'W�<S��<���<�E�<Ȑ�<?٘<��<�c�<M��<��<�%�<�b�<���<�؊<��<�I�<a��<(��<�<<�<|�|<qy<�pu<�q<(9n<��j<� g<�dc<��_<�.\<۔X<�T<�dQ<��M<�:J<I�F<2C<��?<x�;<Iw8<�4<%p1<��-<�v*<��&<4�#<� <��<�O</�<��<6><��<J�<�^<�<E��;�k�;��;��;Ԑ�;�c�;bE�;v5�;�4�;C�;�`�;��;I˴;�;fu�;��;`�;�;e��;;�;M��;�Ƀ;aS};�3s;�4i;�U_;�U;��K;xB;9;��/;A�&;�;%�;^�;�F;e�:�s�:��: /�:Nٲ:ᴢ:��:,��:h�f:g�G:�t):�I:���9�ğ9Z�J9�n�8l`�����X~�����vV�,��;�-���H� �c�vC~��W���w��
���hv���W���%ͺF�ٺ(��)�������Q�̃�s�������$��+��*1�G>7�N=�iZC� dI�fjO��nU��p[��pa��og�Tmm�js�Pfy��a�Ю�����#���%���q��������������������  �  \j=�	=��={G=�=k�=x"=<� =�] =���<�.�<�g�<���<���<��<B�<Cv�<p��<��<s�<1<�<�j�<��<���<2��</�<�>�<pd�<���<��<���<���<��<�"�<i;�<;R�<�f�<%y�<��<���<ǡ�<G��<3��<W��<ȳ�<F��<��<y��<���<V��<lw�<Fb�<�I�<�-�<E�<E��<���<E��<Gl�<l:�<��<>��<܍�<�L�<3�<��<�p�<P�<���<�p�<!�<���<RL�<��<ru�<�<ߎ�<��<٘�<.�<Ó�<��<��<��<Y^�<dȬ<!/�<���<�<bP�<Ѫ�<X�<$W�<K��<���<F�<���<L٘<��<�c�<V��<��<�%�<�b�<���<�؊<��<�I�<b��<0��<
�<B�<m�|<�y<�pu<��q<*9n<�j<� g<�dc<��_<�.\<�X<9�T<�dQ<��M<q:J<S�F<2C<��?<��;<Aw8<�4<p1<��-<�v*<  '<+�#<� <ȴ<pO<6�<�<"><��<8�<�^<�<W��;vk�;�;
��;Ȑ�;�c�;?E�;�5�;�4�;�B�;�`�;���;7˴;�;fu�;h�;e`�;!�;S��;,;�;'��;�Ƀ;>S};4s;�4i;�U_;�U;w�K;�wB;9;E�/;�&;#�;v�;�;�F;(e�:�s�:���:�.�:�ز:ʹ�:Y��:���:��f:��G:�u):WI:=��9Wʟ96�J9�l�8\����Z~�J����V����-���H��c�2C~��W��Bw������%v���W���%ͺ��ٺZ�溉)󺅵����R�l��{�������$��+��*1�i>7� N=��ZC��cI�gjO��nU��p[�:qa�|og��mm��is��ey�Pb�ͮ�����;���3���j�������|���`���௚��  �  Yj=�	=��=}G=�=g�={"=:� =�] =���<�.�<�g�<���<���<��<B�<8v�<s��<��<{�<><�<�j�<��<���<9��<1�<�>�<ud�<���<��<���<���<��<�"�<r;�<9R�<�f�<y�<��<���<���<K��<0��<Y��<ų�<P��<��<{��<���<V��<~w�<Bb�<�I�<�-�<F�<C��<���<G��<:l�<q:�<��<N��<ߍ�<�L�<6�<��<�p�<M�<���<�p�<#�<���<=L�<��<ou�<�<ݎ�<��<ݘ�</�<͓�<��<��<��<\^�<aȬ<"/�<���<�<hP�<˪�<c�<1W�<H��<���<�E�<���<C٘<��<�c�<Q��<��<�%�<�b�<���<�؊<��<�I�<i��<-��<�<=�<}�|<dy<�pu<�q<!9n<�j<� g<ec<��_<�.\<�X<�T<�dQ<��M<~:J<M�F<<C<��?<u�;<Mw8<�4<8p1<��-<�v*<  '<�#<� <��<zO<�<�<#><��<Q�<�^< <2��;�k�;�;���;ސ�;�c�;EE�;f5�;�4�;C�;�`�;��;-˴;G�;Pu�;��;`�;��;b��;;�;/��;�Ƀ;�S};�3s;�4i;�U_;�U;�K;�wB;A9;��/;�&;�;H�;)�;mF;ue�:Ws�:���:�.�:ٲ:���:���:O��:[�f:�G:Ku):�I:���9Kş9~�J9Ji�8�:෕���W~�U����V�E����-���H�$�c��B~��W��<w��,����v��_W�� &ͺ�ٺ��溺)�G������Q����n�������$��+��*1��=7� N=�rZC��cI��jO��nU��p[�qa��og�Smm�Fjs�-fy��a�߮��⬅�H���
���s���������������ȯ���  �  Uj=�	=��=zG=�=j�=|"=6� =�] =|��</�<�g�<���<���<��<B�<:v�<o��<���<m�<1<�<�j�<���<���<?��<(�<�>�<}d�<���<1��<���<���<��<�"�<o;�<0R�<�f�<y�<$��<���<ѡ�<P��<.��<h��<���<N��<��<|��<���<H��<qw�<=b�<�I�<�-�<V�<C��<���<Y��<7l�<s:�<��<A��<Ѝ�<�L�<8�<��<�p�<>�<���<�p�<&�<ı�<<L�<��<du�<�<Վ�<��<ژ�<%�<̓�<��<.��<��<a^�<cȬ</�<���<�<kP�<Ǫ�<S�<"W�<H��<���<�E�<Ր�<:٘<��<�c�<M��<��<�%�<�b�<���<�؊<��<�I�<b��< ��<�<5�<��|<�y<�pu<�q<9n<�j<� g<ec<��_<�.\<��X<*�T<�dQ<��M<�:J<:�F<.C<��?<�;<Rw8<�4<!p1<��-<�v*<��&<(�#<� <��<�O<"�<�<,><��<7�<�^<	 <@��;�k�;��;���;���;�c�;�E�;x5�;�4�;�B�;�`�;��;˴;M�;!u�;��;`�;H�;x��;;�;i��;�Ƀ;S};�3s;�4i;�U_;�U;��K;�wB;`9;��/;��&;�; �;��;UF;�e�:�r�:��:�-�:�ز:��:��:j��:p�f:X�G:4u):�I:f��9�ğ98�J9�^�8{1෍���Y~������X�o��!�-���H�j�c�;B~��W���w��Ӏ��mv��(W��b&ͺ�ٺn�溺)�~�����JQ����'�������$��+��*1�A>7�uN=�YZC��cI�]jO��nU�q[��pa��og��lm��is�Pfy��a����嬅�f������������������|��������  �  Tj=�	=��=}G=�=j�=u"=>� =�] =���</�<�g�<���<���<��<B�<<v�<j��<���<}�<8<�<�j�<��<���<0��<6�<�>�<vd�<���<��<���<���<��<�"�<t;�<7R�<�f�<!y�<��<���<ġ�<8��<-��<_��<̳�<F��<��<w��<���<\��<yw�<Pb�<�I�<�-�<E�<@��<���<G��<:l�<i:�<��<L��<��<�L�<0�<��<�p�<R�<���<�p�<�<���<DL�<��<ru�< �<܎�<��<ᘷ<2�<ȓ�<��<��<��<]^�<hȬ<&/�<���<
�<^P�<ժ�<_�<2W�<T��<���<�E�<���<A٘<��<�c�<O��<��<�%�<�b�<���<�؊<��<�I�<e��<3��<�<6�<[�|<|y<�pu<�q<#9n<�j<� g<ec<��_<�.\<�X<(�T<�dQ<��M<�:J<X�F<=C<��?<��;<7w8<!�4<(p1<��-<�v*<��&<"�#<� <��<uO<&�<��<5><��<F�<�^<�<Q��;ok�;�;��;��;�c�;)E�;�5�;�4�;C�;�`�;��;(˴;F�;Vu�;��;3`�;�;��;;�;F��;�Ƀ;@S};�3s;�4i;�U_;�U;��K;4xB;9;��/; �&;��;(�;#�;hF;�d�:$t�:���:0/�:Kٲ:���:/��:���:��f:��G:u):rG:���9�Ɵ9�J9Bl�8S.���W~�/����U�����-�>�H��c��B~�~W���v��ց��>v���W���%ͺS�ٺy��)�ܵ�����Q�ă���������$��+�b*1�!>7��M=��ZC��cI�ojO��nU�ip[��pa��og��mm��is�fy��a�ۮ��鬅�B������n��������������������  �  7k=�
=�=�H=��=/�=i$=[� =�_ =���<^4�<~m�<̥�<=��<��<lI�<$~�<���<K��<��<�E�<�t�<���<���<���<h#�<PK�<�q�<|��<���<���<.��<��<<3�<�L�<2d�<Zy�<Q��<��<��<��<��<���<G��<k��<���<���<���<��<���<���<~�<
f�<�J�<�+�<	�<���<���<i��<�Y�<�$�<T��<1��<m�< (�<���<���<e@�<���<���<4�<���<�l�<M�<���<$�<���<5�<���<�6�<���< )�<<&�<�y�<6�<YI�<��<��<bh�<¤<��<�l�<��<��<	Y�<բ�<��<�/�<Us�<Ѵ�<c��<U2�<n�<R��<��<��<�Q�<W��<4��<��<V#�<٫|<�y<su<��q<�7n<��j<��f<�]c<��_<�#\<�X<��T<)TQ<A�M<&J<�F< C<�p?<��;<�Y8<��4<�N1<f�-<�Q*<�&<kd#<�<{�<\!<x�<�b<<�<�l<�&<��<�Y�;���;˙�;�M�;f�;2��;���;���;���;a��;5Կ;A �;(<�;凮;"�;�P�;�͝;V[�;:��;᧍;�f�;$7�;�.|;�r;h;�5^;6yT;;�J;�_A;�8;��.;��%;��;
�;��
;�I;s�:܋�:��:�Y�:��:���:]�:+Q�:��c:��D:�`&:�J:��9a �9��?9/'�84e����O���������������/���J��e�r��I?��dT��"V��uA�������ͺ�ں#9�;��( �sc����V�������!/%�fH+�w\1��m7��y=�C�C�p�I�T�O�ЎU���[�ԋa�G�g��m��{s��uy��n�������������6���F���ا��������������  �  :k=�
=�=�H=��=)�=d$=W� =�_ =���<^4�<zm�<ĥ�<=��<��<qI�<~�<���<B��<��<�E�<�t�<���<���<���<j#�<aK�<�q�<{��<���<���<8��<��<N3�<�L�<%d�<ky�<Z��<���<��<۶�<���<���<d��<e��<���<���<��<��<��<���<~�<f�<�J�<�+�<	�<���<���<Y��<�Y�<�$�<]��<>��<m�<�'�<���<���<`@�<��<���<4�<���<�l�<_�<���<$�<v��<5�<���<�6�<���<)�<圱<"�<�y�<M�<XI�<"��<��<Yh�<���<��<�l�<��<��<�X�<ܢ�<{�<�/�<Ps�<ʴ�<g��<Q2�<�n�<O��<��<��<�Q�<]��<1��</��<\#�<��|<�y<su<��q<�7n<יj<��f<^c<��_<$\<#�X<w�T<TQ<K�M<G&J<�F<  C<�p?<��;<zY8<s�4<�N1<b�-<�Q*<��&<[d#<�<e�<f!<]�<�b<<�<�l<�&<��<�Y�;��;ә�;8N�;��;-��;i��;���;ī�;g��;}Կ;S �;�;�;)��;H�;�P�;�͝;&[�;��;��;Gg�;7�;�.|;Wr;�h;�5^;cyT;��J;�_A;�8;;�.;̢%;Ƞ;�;+�
;I;>s�:%��:���:�Z�:��:���:��:�Q�:�c:\�D:�b&:"J:�9��9ڝ?9�.�8�@����_���������2��
�/���J���e�
���=��iT���U��=B��Z��6�ͺ�ں9����( ��c�c����������V/%�HH+��\1�m7��y=�v�C�׉I�b�O���U���[���a��g�Z�m�|s��uy�_n�ó��v���ĭ���������ϧ������F���*����  �  6k=�
=ک=�H=��=,�=m$=U� =�_ =|��<c4�<m�<ʥ�<D��<��<~I�<~�<Ʊ�<D��<��<�E�<�t�<���<���<���<_#�<UK�<�q�<y��<���<���<@��<��<I3�<�L�<'d�<iy�<D��<���<��<��<��<���<[��<R��<���<���<���<��<���<���<~�<f�<�J�<�+�<	�<���<��<S��<�Y�<�$�<`��<<��<m�<(�<���<���<L@�<��<���< 4�<���<�l�<]�<���<$�<y��<5�<���<�6�<���<)�<�<!�<�y�<B�<II�<(��<��<jh�<���<��<�l�<��<��<�X�<袚<t�<�/�<Ys�<̴�<p��<D2�<�n�<L��<��<��<�Q�<b��< ��<&��<T#�<׫|<�y<su<��q<�7n<ڙj<��f<^c<��_<�#\<1�X<��T<'TQ<=�M<2&J<��F< C<�p?<��;<�Y8<h�4<�N1<J�-<�Q*<	�&<gd#<,�<X�<�!<\�<�b<<�<�l<�&<��<�Y�;��;���;	N�;��;$��;���;���;��;#��;gԿ;] �;�;�; ��;��;�P�;�͝;N[�;B��;ӧ�;&g�;�6�;�.|;kr;&h;
6^;LyT;��J;a_A;^8;�.;%�%;��;�;��
;�H;At�:��:���:�Z�:��:���:��:#R�:��c:F�D:�`&:TK:��9��9��?9Y�8�A����Z�������1�����O�/�q�J���e�����>��aU��GU��&B��7��A�ͺ�ںH9����,( �
d� ����������I/%�H+��\1� m7�z=��C���I�L�O�w�U�@�[�*�a�Y�g��m��{s�vuy��n����p��������?�����������2��������  �  9k=�
=�=�H=��='�=f$=X� =�_ =���<_4�<wm�<˥�<?��<��<uI�<~�<���<E��<��<�E�<�t�<���<���<���<h#�<dK�<�q�<|��<���<���<:��<��<H3�<�L�<5d�<^y�<S��<���<��<ڶ�<��<���<\��<i��<���<���<��<	��<���<���<~�<f�<�J�<�+�<	�<���<���<V��<�Y�<�$�<b��<7��<m�<�'�<���<���<a@�<��<���< 4�<���<�l�<[�<���<$�<���<5�<���<�6�<���<)�<朱<%�<�y�<M�<VI�<"��<��<\h�<���<��<�l�<��<��<�X�<ߢ�<{�<�/�<Ys�<Ŵ�<g��<L2�<�n�<R��<��<��<�Q�<`��<7��<��<X#�<ҫ|<�y<su<��q<�7n<��j<��f<�]c<��_<$\<,�X<v�T<TQ<G�M<'&J<"�F<% C<�p?<��;<�Y8<x�4<�N1<]�-<�Q*<��&<jd#<!�<i�<m!<e�<�b<
<$�<�l<�&<��<pY�;��;ʙ�;DN�;��;0��;y��;���;ͫ�;X��;cԿ;D �;7<�;�;-�;�P�;�͝;![�;D��;٧�;)g�;7�;�.|;&r;�h;�5^;CyT;��J;�_A;�8;�.;��%;��;��;B�
;�H;@s�:T��:���:@Z�:��:���:>�:�Q�:.�c:��D:�`&:bK:��9��9r�?9�*�8aU����s������V��m���/���J�=�e����=���T���U���B���� �ͺt�ں�8纨��( ��c�I����������}/%�GH+��\1�/m7��y=�|�C��I���O���U���[�\�a�6�g��m�(|s�tuy�Vn�泂���������%���)���ԧ������H�������  �  >k=�
=�=�H=��=/�=f$=Z� =�_ =���<a4�<|m�<Υ�<9��<��<kI�<%~�<���<G��<��<�E�<�t�<���< ��<���<^#�<[K�<�q�<���<���<���</��<��<K3�<�L�<5d�<Wy�<\��<��<*��<ֶ�<��<���<V��<_��<���<���<���<��<���<���<~�<f�<�J�<�+�<	�<���<���<f��<�Y�<�$�<Z��<7��<m�<�'�<���<���<V@�<���<���< 4�<���< m�<K�<���<$�<���<5�<���<�6�<���<")�<���<,�<�y�<F�<MI�<&��<��<\h�<¤<��<�l�<��<��<Y�<֢�<��<�/�<Ys�<ϴ�<g��<U2�<�n�<U��<��<��<�Q�<T��</��<��<b#�<ī|<�y<su<��q<�7n<��j<��f<�]c<��_<�#\<'�X<~�T<TQ<[�M<!&J<�F<
 C<�p?<��;<Y8<��4<�N1<k�-<�Q*<�&<qd#<�<w�<Z!<y�<�b<<$�<�l<�&<��<�Y�;'��;���;"N�;��;W��;Z��;���;���;O��;pԿ;1 �;5<�;ه�;P�;�P�;�͝;[�;4��;���;g�;�6�;~.|;�r;�h;6^;FyT;l�J;�_A;�8;��.;�%;��;�;�
;kI;�r�:���:t��:IZ�:�:0��:��:gQ�:щc:��D:�a&:mK:��9�"�9��?9Q1�8�b�������槻�?������/���J�U�e����N>��U��mU��_A������ͺʕں�8����( �uc����>������2/%�FH+�r\1��m7��y=�Z�C�p�I��O��U�ʍ[�y�a��g�=�m�|s�cuy��n�������������>��������������7���.����  �  7k=�
=�=�H=��=(�=k$=W� =�_ =���<b4�<ym�<ɥ�<@��<��<tI�<~�<���<J��<��<�E�<�t�<���<���<���<e#�<eK�<�q�<��<���<���<;��<��<M3�<�L�<)d�<`y�<T��<��<)��<۶�<��<���<a��<b��<���<���<��<��<���<���<~�<f�<�J�<�+�<	�<���< ��<V��<�Y�<�$�<_��<8��<m�<�'�<���<���<Z@�<��<���<#4�<���<�l�<P�<���<$�<z��<5�<���<�6�<���<)�<朱<'�<�y�<Q�<SI�<��<��<ch�<���<��<�l�<��<��<�X�<ޢ�<��<�/�<Ws�<Ǵ�<h��<P2�<�n�<N��<��<��<�Q�<b��<3��<$��<R#�<׫|<�y<su<��q<�7n<ęj<��f<�]c<��_<�#\<5�X<�T<$TQ<>�M<-&J<�F< C<�p?<��;<�Y8<q�4<�N1<]�-<�Q*<��&<gd#<#�<p�<m!<d�<�b<<�<�l<�&<��<�Y�;���;�;JN�;��;<��;��;���;ҫ�;>��;|Կ;A �;<�;���;2�;�P�;�͝;%[�;G��;̧�;=g�;�6�;�.|;>r;�h;
6^;0yT;��J;�_A;�8;$�.;�%;ʠ;"�;I�
;�H;s�:���:���:LZ�: �:��:m�:�Q�:a�c:��D:�`&:�K:��9�!�9'�?9�(�8�Q� �����������������/���J�ۗe�#���=���T���U��{B������ͺH�ں�8�C��( ��c�M��U�������k/%�BH+��\1�m7�z=��C��I�y�O�w�U���[�;�a�j�g��m��{s�Muy��n�ҳ����������������
���~���6��������  �  2k=�
=ީ=�H=��=)�=k$=S� =�_ =y��<c4�<zm�<˥�<H��<��<�I�<~�<���<D��<��<�E�<�t�<���<���<���<_#�<]K�<�q�<v��<���<���<;��<��<M3�<�L�<'d�<ly�<N��<��<��<׶�<��<��<g��<X��<���<���<���<��<���<���<~�<f�<�J�<�+�<	�<���<��<V��<�Y�<�$�<^��<9��<m�<(�<���<���<Q@�<��<���<!4�<���<�l�<V�<���<$�<y��<5�<���<�6�<���<)�<뜱< �<�y�<M�<KI�<"��<��<mh�<���<��<�l�<��<��<�X�<뢚<w�<�/�<\s�<Ǵ�<n��<B2�<�n�<I��<��<��<�Q�<[��<'��<.��<K#�<�|<�y<su<��q<�7n<ՙj<��f<^c<��_<�#\<*�X<c�T<6TQ<-�M<?&J<�F< C<�p?<��;<�Y8<b�4<�N1<D�-<�Q*<��&<jd#<2�<[�<�!<c�<�b<	<�<m<�&<��<}Y�;���;���;+N�;��;��;���;c��;Ы�;2��;{Կ;K �;�;�;-��;�;�P�;�͝;[�;T��;���;Vg�;�6�;�.|;*r;h;�5^;.yT;��J;Y_A;(8;�.;E�%; ;�;��
;�H;�s�:��:���:aZ�:��:���:E�:�Q�:=�c:��D:`&:|K:b�9��9t�?9V#�8�=�y��5���������@��-�/��J�ǘe�����=��5U���U���B������ͺ˔ںB9线��( ��c���������v�m/%�H+�
]1��l7�0z=�4�C���I�z�O���U��[��a���g���m�\|s��uy��n��z���ǭ������-�����������n���۩���  �  6k=�
=ݩ=�H=��=.�=g$=W� =�_ =���<h4�<wm�<ϥ�<C��<��<vI�<!~�<���<M��<��<�E�<�t�<���<���<���<a#�<UK�<�q�<{��<���<���<3��<��<G3�<�L�<0d�<^y�<M��<��<'��<ڶ�<��<���<]��<Z��<���<���<���<��< ��<���<~�<f�<�J�<�+�<	�<���<��<[��<�Y�<�$�<_��<=��<m�<(�<���<���<S@�<��<���<4�<���<�l�<L�<���<$�<~��<5�<���<�6�<���<)�<眱<!�<�y�<B�<NI�<%��<��<eh�<���<��<�l�<��<��<Y�<࢚<z�<�/�<]s�<ȴ�<p��<N2�<�n�<R��<��<��<�Q�<X��<(��<(��<T#�<ϫ|<�y<su<��q<�7n<��j<��f<�]c<��_<�#\<+�X<y�T<TQ<=�M<:&J<�F< C<�p?<��;<�Y8<u�4<�N1<`�-<�Q*<��&<qd#<)�<b�<q!<r�<b<< �<�l<�&<��<�Y�;��;���;N�;��;+��;~��;���;���;6��;`Կ;9 �;%<�;���;�;�P�;�͝;#[�;<��;ק�;+g�;�6�;�.|;jr;4h;�5^;^yT;��J;�_A;8;>�.;%�%;��;�;b�
;I;Ss�:���:���:�Z�:��:���:��:�Q�:��c:[�D:a&:(K:��9�!�9?�?9�"�8W����n���٧��v��n��#�/���J���e�����>��U��{U���A�����L�ͺ�ں�8� ���( ��c�A��������n�c/%��G+��\1�m7��y=�`�C�t�I�S�O�ÎU���[��a�V�g��m�|s�auy��n�쳂������������0�����������A�������  �  :k=�
=�=�H=��=+�=e$=^� =�_ =���<_4�<{m�<ҥ�<9��<��<mI�<&~�<���<L��<��<�E�<�t�<���<���<���<p#�<dK�<�q�<���<|��<���<2��<��<H3�<�L�<3d�<Wy�<\��<��<$��<ٶ�<���<���<X��<m��<���<���<��<��<��<���<~�<f�<�J�<�+�<	�<���<���<c��<�Y�<�$�<[��<<��<m�<�'�<���<���<f@�<��<���<4�<���<�l�<I�<���<$�<��<�4�<���<�6�<���<)�<ݜ�<&�<�y�<L�<]I�<��<��<[h�<¤<��<�l�<��<��<	Y�<֢�<��<�/�<]s�<̴�<e��<S2�<�n�<[��<��<��<�Q�<g��<9��<��<[#�<��|<�y<su<��q<�7n<��j<��f<�]c<��_<�#\<(�X<��T<TQ<L�M<$&J<!�F<2 C<p?<��;<}Y8<��4<�N1<d�-<�Q*< �&<xd#<�<{�<_!<|�<�b<<�<�l<�&<��<�Y�;���;��;EN�;��;C��;L��;���;���;Y��;eԿ;* �;0<�;ۇ�;S�;�P�;�͝; [�;��;맍;g�;,7�;�.|;<r;�h;�5^;oyT;��J;`A;�8;x�.;�%;Š;"�;"�
;YI;�r�:��:���:�Z�:�:���:�:�Q�:�c:^�D:Ga&:�J:��9x!�9В?9r3�8�b�{�����`����������/���J�
�e�����=��T��:V��B��1��w�ͺs�ں,9����( �rc����,�����p�C/%�[H+��\1�am7��y=�e�C���I���O�L�U�{�[�m�a��g�e�m��{s�zuy��n�ų��Ȱ������A��������������#���>����  �  8k=�
=۩=�H=��=0�=f$=Y� =�_ =���<d4�<�m�<˥�<>��<��<tI�<~�<Ʊ�<F��<��<�E�<�t�<���<���<���<^#�<VK�<�q�<~��<���<���<4��<��<H3�<�L�<*d�<_y�<O��<��<!��<߶�<��<���<W��<V��<���<���<���<��<���<���<~�<f�<�J�<�+�<	�<���< ��<^��<�Y�<�$�<^��<:��<m�<�'�<���<���<P@�<��<���<4�<���<�l�<O�<���<$�<y��<�4�<���<�6�<���<)�<眱<%�<�y�<B�<JI�<"��<��<`h�<���<��<�l�<��<��<�X�<ܢ�<��<�/�<Xs�<д�<n��<M2�<�n�<Q��<��<��<�Q�<\��<$��< ��<U#�<˫|<�y<su<��q<�7n<��j<��f<�]c<��_<�#\<#�X<|�T<TQ<C�M<(&J<��F< C<�p?<��;<�Y8<z�4<�N1<Y�-<�Q*<�&<jd#< �<~�<l!<i�<�b<<�<�l<�&<��<�Y�;��;���;N�;s�;8��;u��;���;���;.��;gԿ;9 �;<�;���;�;�P�;�͝;6[�;0��;֧�;g�;�6�;�.|;�r;h;�5^;FyT;��J;�_A;*8;k�.;��%;�;>�;M�
;4I;�s�:)��:���:pZ�:��:l��:'�:�Q�:�c:%�D:}`&:�J:��9@ �9�?9�#�8>W�~��0���������*����/���J�+�e�T���>��FU���U���A������ͺ�ں�8线��J( ��c�[��*�������#/%�H+��\1�m7��y=�_�C�l�I�<�O���U� �[�U�a�L�g�"�m��{s��uy��n�곂���������"���+����������;�������  �  4k=�
=�=�H=��=%�=i$=W� =�_ =���<h4�<xm�<ǥ�<K��<��<�I�<~�<���<D��<��<�E�<�t�<���<���<���<f#�<aK�<�q�<y��<���<���<>��<��<J3�<�L�<#d�<hy�<I��<���<��<׶�<��<���<e��<_��<���<���<��<��<���<���<~�<f�<�J�<�+�<	�<���<	��<L��<�Y�<�$�<j��<8��<m�<�'�<���<���<X@�<��<���<!4�<���<�l�<`�<���<$�<u��<�4�<���<�6�<���<)�<眱<$�<�y�<N�<SI�<)��<��<bh�<���<��<�l�<���<��<�X�<颚<v�<�/�<Ws�<Ĵ�<s��<N2�<�n�<M��<��<��<�Q�<`��</��<.��<N#�<ݫ|<�y<su<��q<�7n<ҙj<��f<�]c<��_<�#\<(�X<h�T<)TQ<3�M<C&J<�F<  C<�p?<��;<�Y8<s�4<�N1<b�-<�Q*<��&<cd#<:�<\�<�!<W�<�b<	<.�<�l<�&<��<^Y�; ��;Ǚ�;9N�;��;&��;���;f��;ܫ�;A��;nԿ;B �;�;�;��;�;�P�;�͝;[�;H��;ӧ�;Ng�;�6�;�.|;r;�h;�5^;.yT;��J;�_A;N8;��.;3�%;ڠ;�;��
;�H;t�:���:s��:[Z�:��: ��:�
�:$R�:%�c:��D:�`&:�K:��9��9^�?9	 �8�E�K���������_�����/���J�B�e�����=���T��/U��
C�����/�ͺ'�ںE8����_( �&d�������������/%��G+��\1��l7�z=�F�C���I�{�O���U�ʍ[��a���g�فm�R|s��uy�Xn���������ɭ�����4���ߧ������b��������  �  6k=�
=ީ=�H=��=,�=n$=Y� =�_ =���<_4�<�m�<ѥ�<H��<��<�I�<%~�<ı�<A��<��<�E�<�t�<���<���<���<d#�<WK�<�q�<|��<���<���<4��<��<@3�<�L�<+d�<\y�<L��<��<��<ض�<	��<���<S��<^��<���<���<���<��<���<���<~�<f�<�J�<�+�<	�<���<	��<a��<�Y�<�$�<_��<1��<&m�< (�<���<���<W@�<���<���<#4�<���<�l�<O�<���<$�<{��<5�<���<�6�<���<)�<䜱<'�<�y�<A�<QI�<"��<��<jh�<¤<��<�l�< ��<��<Y�<뢚<u�<�/�<_s�<մ�<j��<L2�<�n�<Q��<��<��<�Q�<]��<+��<��<T#�<٫|<�y<su<��q<�7n<��j<��f<�]c<��_<�#\<!�X<~�T<#TQ<=�M<&J<�F< C<�p?<��;<�Y8<|�4<�N1<Y�-<�Q*<�&<wd#<3�<Z�<�!<{�<�b<<�<�l<�&<��<�Y�;��;���;N�;z�;3��;{��;���;���;A��;FԿ;> �;<�;���;�;�P�;�͝;[�;K��;̧�;g�;�6�;�.|;�r;h;d6^;$yT;��J;�_A;@8;w�.;?�%;��;�;��
;GI;#t�:8��:���:�Y�:��:���::�:�Q�:
�c:|�D:`&:�K:v�95�9�?9*%�8]�5��c����������V����/���J�ϗe�a���>���T���U���A��1��s�ͺ�ں�8����7( �|c���������`�/%�1H+��\1�@m7��y=�܂C���I�5�O���U��[���a�\�g��m�|s��uy��n�������������.���F�����������7��� ����  �  ;k=�
=�=�H=��=)�=a$=X� =�_ =���<Z4�<�m�<¥�<;��<��<qI�<~�<���<A��<��<�E�<�t�<���<���<���<g#�<dK�<�q�<}��<u��<���</��<��<C3�<�L�</d�<Uy�<]��<��<(��<ն�<���<���<^��<k��<���<���<��<��<���<���<~�<f�<�J�<�+�<	�<���<���<[��<�Y�<�$�<i��<6��<m�<�'�<���<���<c@�<
��<���<4�<���<�l�<L�<���<$�<|��<5�<���<�6�<���< )�<ל�<$�<�y�<N�<WI�<��<��<Lh�< ¤<��<�l�<��<��<�X�<ڢ�<��<�/�<Ls�<Ӵ�<a��<[2�<�n�<P��<��<��<�Q�<X��<7��<%��<\#�<��|<�y<su<��q<�7n<��j<��f<�]c<��_<�#\<'�X<��T<�SQ<Q�M<3&J<�F< C<�p?<��;<nY8<v�4<�N1<z�-<�Q*<�&<Xd#<�<s�<e!<e�<�b<<7�<�l<�&<q�<�Y�;���;ș�;FN�;��;3��;2��;���;���;f��;TԿ;C �;<�;Ӈ�;T�;�P�;�͝;[�;
��;觍;2g�;%7�;�.|;�r;Kh;�5^;HyT;��J;�_A;�8;Z�.;��%;�;H�;�
;I;s�:s��:m��:;Z�:��:��:v�:#Q�:��c:D�D:�`&:�I:�
�9)"�9��?95�8�j����{�������e�������/���J�5�e����=���T��0V���A������ͺ3�ں#8����( ��c�m��U�������/%�zH+�D\1��l7��y=���C���I�J�O�ƎU���[�2�a��g���m�|s�`uy��n�̳����������/������六�����0���Y����  �  6k=�
=ީ=�H=��=,�=n$=Y� =�_ =���<_4�<�m�<ѥ�<H��<��<�I�<%~�<ı�<A��<��<�E�<�t�<���<���<���<d#�<WK�<�q�<|��<���<���<4��<��<@3�<�L�<+d�<\y�<L��<��<��<ض�<	��<���<S��<^��<���<���<���<��<���<���<~�<f�<�J�<�+�<	�<���<	��<a��<�Y�<�$�<_��<1��<&m�< (�<���<���<W@�<���<���<#4�<���<�l�<O�<���<$�<{��<5�<���<�6�<���<)�<䜱<'�<�y�<A�<QI�<"��<��<jh�<¤<��<�l�< ��<��<Y�<뢚<u�<�/�<_s�<մ�<j��<L2�<�n�<Q��<��<��<�Q�<]��<+��<��<T#�<٫|<�y<su<��q<�7n<��j<��f<�]c<��_<�#\<!�X<~�T<#TQ<=�M<&J<�F< C<�p?<��;<�Y8<|�4<�N1<Y�-<�Q*<�&<wd#<3�<Z�<�!<{�<�b<<�<�l<�&<��<�Y�;��;���;N�;z�;3��;{��;���;���;A��;FԿ;> �;<�;���;�;�P�;�͝;[�;K��;̧�;g�;�6�;�.|;�r;h;d6^;$yT;��J;�_A;@8;w�.;?�%;��;�;��
;GI;#t�:8��:���:�Y�:��:���::�:�Q�:
�c:|�D:`&:�K:v�95�9�?9*%�8]�5��c����������V����/���J�ϗe�a���>���T���U���A��1��s�ͺ�ں�8����7( �|c���������`�/%�1H+��\1�@m7��y=�܂C���I�5�O���U��[���a�\�g��m�|s��uy��n�������������.���F�����������7��� ����  �  4k=�
=�=�H=��=%�=i$=W� =�_ =���<h4�<xm�<ǥ�<K��<��<�I�<~�<���<D��<��<�E�<�t�<���<���<���<f#�<aK�<�q�<y��<���<���<>��<��<J3�<�L�<#d�<hy�<I��<���<��<׶�<��<���<e��<_��<���<���<��<��<���<���<~�<f�<�J�<�+�<	�<���<	��<L��<�Y�<�$�<j��<8��<m�<�'�<���<���<X@�<��<���<!4�<���<�l�<`�<���<$�<u��<�4�<���<�6�<���<)�<眱<$�<�y�<N�<SI�<)��<��<bh�<���<��<�l�<���<��<�X�<颚<v�<�/�<Ws�<Ĵ�<s��<N2�<�n�<M��<��<��<�Q�<`��</��<.��<N#�<ݫ|<�y<su<��q<�7n<ҙj<��f<�]c<��_<�#\<(�X<h�T<)TQ<3�M<C&J<�F<  C<�p?<��;<�Y8<s�4<�N1<b�-<�Q*<��&<cd#<:�<\�<�!<W�<�b<	<.�<�l<�&<��<^Y�; ��;Ǚ�;9N�;��;&��;���;f��;ܫ�;A��;nԿ;B �;�;�;��;�;�P�;�͝;[�;H��;ӧ�;Ng�;�6�;�.|;r;�h;�5^;.yT;��J;�_A;N8;��.;3�%;ڠ;�;��
;�H;t�:���:s��:[Z�:��: ��:�
�:$R�:%�c:��D:�`&:�K:��9��9^�?9	 �8�E�K���������_�����/���J�B�e�����=���T��/U��
C�����/�ͺ'�ںE8����_( �&d�������������/%��G+��\1��l7�z=�F�C���I�{�O���U�ʍ[��a���g�فm�R|s��uy�Xn���������ɭ�����4���ߧ������b��������  �  8k=�
=۩=�H=��=0�=f$=Y� =�_ =���<d4�<�m�<˥�<>��<��<tI�<~�<Ʊ�<F��<��<�E�<�t�<���<���<���<^#�<VK�<�q�<~��<���<���<4��<��<H3�<�L�<*d�<_y�<O��<��<!��<߶�<��<���<W��<V��<���<���<���<��<���<���<~�<f�<�J�<�+�<	�<���< ��<^��<�Y�<�$�<^��<:��<m�<�'�<���<���<P@�<��<���<4�<���<�l�<O�<���<$�<y��<�4�<���<�6�<���<)�<眱<%�<�y�<B�<JI�<"��<��<`h�<���<��<�l�<��<��<�X�<ܢ�<��<�/�<Xs�<д�<n��<M2�<�n�<Q��<��<��<�Q�<\��<$��< ��<U#�<˫|<�y<su<��q<�7n<��j<��f<�]c<��_<�#\<#�X<|�T<TQ<C�M<(&J<��F< C<�p?<��;<�Y8<z�4<�N1<Y�-<�Q*<�&<jd#< �<~�<l!<i�<�b<<�<�l<�&<��<�Y�;��;���;N�;s�;8��;u��;���;���;.��;gԿ;9 �;<�;���;�;�P�;�͝;6[�;0��;֧�;g�;�6�;�.|;�r;h;�5^;FyT;��J;�_A;*8;k�.;��%;�;>�;M�
;4I;�s�:)��:���:pZ�:��:l��:'�:�Q�:�c:%�D:}`&:�J:��9@ �9�?9�#�8>W�~��0���������*����/���J�+�e�T���>��FU���U���A������ͺ�ں�8线��J( ��c�[��*�������#/%�H+��\1�m7��y=�_�C�l�I�<�O���U� �[�U�a�L�g�"�m��{s��uy��n�곂���������"���+����������;�������  �  :k=�
=�=�H=��=+�=e$=^� =�_ =���<_4�<{m�<ҥ�<9��<��<mI�<&~�<���<L��<��<�E�<�t�<���<���<���<p#�<dK�<�q�<���<|��<���<2��<��<H3�<�L�<3d�<Wy�<\��<��<$��<ٶ�<���<���<X��<m��<���<���<��<��<��<���<~�<f�<�J�<�+�<	�<���<���<c��<�Y�<�$�<[��<<��<m�<�'�<���<���<f@�<��<���<4�<���<�l�<I�<���<$�<��<�4�<���<�6�<���<)�<ݜ�<&�<�y�<L�<]I�<��<��<[h�<¤<��<�l�<��<��<	Y�<֢�<��<�/�<]s�<̴�<e��<S2�<�n�<[��<��<��<�Q�<g��<9��<��<[#�<��|<�y<su<��q<�7n<��j<��f<�]c<��_<�#\<(�X<��T<TQ<L�M<$&J<!�F<2 C<p?<��;<}Y8<��4<�N1<d�-<�Q*< �&<xd#<�<{�<_!<|�<�b<<�<�l<�&<��<�Y�;���;��;EN�;��;C��;L��;���;���;Y��;eԿ;* �;0<�;ۇ�;S�;�P�;�͝; [�;��;맍;g�;,7�;�.|;<r;�h;�5^;oyT;��J;`A;�8;x�.;�%;Š;"�;"�
;YI;�r�:��:���:�Z�:�:���:�:�Q�:�c:^�D:Ga&:�J:��9x!�9В?9r3�8�b�{�����`����������/���J�
�e�����=��T��:V��B��1��w�ͺs�ں,9����( �rc����,�����p�C/%�[H+��\1�am7��y=�e�C���I���O�L�U�{�[�m�a��g�e�m��{s�zuy��n�ų��Ȱ������A��������������#���>����  �  6k=�
=ݩ=�H=��=.�=g$=W� =�_ =���<h4�<wm�<ϥ�<C��<��<vI�<!~�<���<M��<��<�E�<�t�<���<���<���<a#�<UK�<�q�<{��<���<���<3��<��<G3�<�L�<0d�<^y�<M��<��<'��<ڶ�<��<���<]��<Z��<���<���<���<��< ��<���<~�<f�<�J�<�+�<	�<���<��<[��<�Y�<�$�<_��<=��<m�<(�<���<���<S@�<��<���<4�<���<�l�<L�<���<$�<~��<5�<���<�6�<���<)�<眱<!�<�y�<B�<NI�<%��<��<eh�<���<��<�l�<��<��<Y�<࢚<z�<�/�<]s�<ȴ�<p��<N2�<�n�<R��<��<��<�Q�<X��<(��<(��<T#�<ϫ|<�y<su<��q<�7n<��j<��f<�]c<��_<�#\<+�X<y�T<TQ<=�M<:&J<�F< C<�p?<��;<�Y8<u�4<�N1<`�-<�Q*<��&<qd#<)�<b�<q!<r�<b<< �<�l<�&<��<�Y�;��;���;N�;��;+��;~��;���;���;6��;`Կ;9 �;%<�;���;�;�P�;�͝;#[�;<��;ק�;+g�;�6�;�.|;jr;4h;�5^;^yT;��J;�_A;8;>�.;%�%;��;�;b�
;I;Ss�:���:���:�Z�:��:���:��:�Q�:��c:[�D:a&:(K:��9�!�9?�?9�"�8W����n���٧��v��n��#�/���J���e�����>��U��{U���A�����L�ͺ�ں�8� ���( ��c�A��������n�c/%��G+��\1�m7��y=�`�C�t�I�S�O�ÎU���[��a�V�g��m�|s�auy��n�쳂������������0�����������A�������  �  2k=�
=ީ=�H=��=)�=k$=S� =�_ =y��<c4�<zm�<˥�<H��<��<�I�<~�<���<D��<��<�E�<�t�<���<���<���<_#�<]K�<�q�<v��<���<���<;��<��<M3�<�L�<'d�<ly�<N��<��<��<׶�<��<��<g��<X��<���<���<���<��<���<���<~�<f�<�J�<�+�<	�<���<��<V��<�Y�<�$�<^��<9��<m�<(�<���<���<Q@�<��<���<!4�<���<�l�<V�<���<$�<y��<5�<���<�6�<���<)�<뜱< �<�y�<M�<KI�<"��<��<mh�<���<��<�l�<��<��<�X�<뢚<w�<�/�<\s�<Ǵ�<n��<B2�<�n�<I��<��<��<�Q�<[��<'��<.��<K#�<�|<�y<su<��q<�7n<ՙj<��f<^c<��_<�#\<*�X<c�T<6TQ<-�M<?&J<�F< C<�p?<��;<�Y8<b�4<�N1<D�-<�Q*<��&<jd#<2�<[�<�!<c�<�b<	<�<m<�&<��<}Y�;���;���;+N�;��;��;���;c��;Ы�;2��;{Կ;K �;�;�;-��;�;�P�;�͝;[�;T��;���;Vg�;�6�;�.|;*r;h;�5^;.yT;��J;Y_A;(8;�.;E�%; ;�;��
;�H;�s�:��:���:aZ�:��:���:E�:�Q�:=�c:��D:`&:|K:b�9��9t�?9V#�8�=�y��5���������@��-�/��J�ǘe�����=��5U���U���B������ͺ˔ںB9线��( ��c���������v�m/%�H+�
]1��l7�0z=�4�C���I�z�O���U��[��a���g���m�\|s��uy��n��z���ǭ������-�����������n���۩���  �  7k=�
=�=�H=��=(�=k$=W� =�_ =���<b4�<ym�<ɥ�<@��<��<tI�<~�<���<J��<��<�E�<�t�<���<���<���<e#�<eK�<�q�<��<���<���<;��<��<M3�<�L�<)d�<`y�<T��<��<)��<۶�<��<���<a��<b��<���<���<��<��<���<���<~�<f�<�J�<�+�<	�<���< ��<V��<�Y�<�$�<_��<8��<m�<�'�<���<���<Z@�<��<���<#4�<���<�l�<P�<���<$�<z��<5�<���<�6�<���<)�<朱<'�<�y�<Q�<SI�<��<��<ch�<���<��<�l�<��<��<�X�<ޢ�<��<�/�<Ws�<Ǵ�<h��<P2�<�n�<N��<��<��<�Q�<b��<3��<$��<R#�<׫|<�y<su<��q<�7n<ęj<��f<�]c<��_<�#\<5�X<�T<$TQ<>�M<-&J<�F< C<�p?<��;<�Y8<q�4<�N1<]�-<�Q*<��&<gd#<#�<p�<m!<d�<�b<<�<�l<�&<��<�Y�;���;�;JN�;��;<��;��;���;ҫ�;>��;|Կ;A �;<�;���;2�;�P�;�͝;%[�;G��;̧�;=g�;�6�;�.|;>r;�h;
6^;0yT;��J;�_A;�8;$�.;�%;ʠ;"�;I�
;�H;s�:���:���:LZ�: �:��:m�:�Q�:a�c:��D:�`&:�K:��9�!�9'�?9�(�8�Q� �����������������/���J�ۗe�#���=���T���U��{B������ͺH�ں�8�C��( ��c�M��U�������k/%�BH+��\1�m7�z=��C��I�y�O�w�U���[�;�a�j�g��m��{s�Muy��n�ҳ����������������
���~���6��������  �  >k=�
=�=�H=��=/�=f$=Z� =�_ =���<a4�<|m�<Υ�<9��<��<kI�<%~�<���<G��<��<�E�<�t�<���< ��<���<^#�<[K�<�q�<���<���<���</��<��<K3�<�L�<5d�<Wy�<\��<��<*��<ֶ�<��<���<V��<_��<���<���<���<��<���<���<~�<f�<�J�<�+�<	�<���<���<f��<�Y�<�$�<Z��<7��<m�<�'�<���<���<V@�<���<���< 4�<���< m�<K�<���<$�<���<5�<���<�6�<���<")�<���<,�<�y�<F�<MI�<&��<��<\h�<¤<��<�l�<��<��<Y�<֢�<��<�/�<Ys�<ϴ�<g��<U2�<�n�<U��<��<��<�Q�<T��</��<��<b#�<ī|<�y<su<��q<�7n<��j<��f<�]c<��_<�#\<'�X<~�T<TQ<[�M<!&J<�F<
 C<�p?<��;<Y8<��4<�N1<k�-<�Q*<�&<qd#<�<w�<Z!<y�<�b<<$�<�l<�&<��<�Y�;'��;���;"N�;��;W��;Z��;���;���;O��;pԿ;1 �;5<�;ه�;P�;�P�;�͝;[�;4��;���;g�;�6�;~.|;�r;�h;6^;FyT;l�J;�_A;�8;��.;�%;��;�;�
;kI;�r�:���:t��:IZ�:�:0��:��:gQ�:щc:��D:�a&:mK:��9�"�9��?9Q1�8�b�������槻�?������/���J�U�e����N>��U��mU��_A������ͺʕں�8����( �uc����>������2/%�FH+�r\1��m7��y=�Z�C�p�I��O��U�ʍ[�y�a��g�=�m�|s�cuy��n�������������>��������������7���.����  �  9k=�
=�=�H=��='�=f$=X� =�_ =���<_4�<wm�<˥�<?��<��<uI�<~�<���<E��<��<�E�<�t�<���<���<���<h#�<dK�<�q�<|��<���<���<:��<��<H3�<�L�<5d�<^y�<S��<���<��<ڶ�<��<���<\��<i��<���<���<��<	��<���<���<~�<f�<�J�<�+�<	�<���<���<V��<�Y�<�$�<b��<7��<m�<�'�<���<���<a@�<��<���< 4�<���<�l�<[�<���<$�<���<5�<���<�6�<���<)�<朱<%�<�y�<M�<VI�<"��<��<\h�<���<��<�l�<��<��<�X�<ߢ�<{�<�/�<Ys�<Ŵ�<g��<L2�<�n�<R��<��<��<�Q�<`��<7��<��<X#�<ҫ|<�y<su<��q<�7n<��j<��f<�]c<��_<$\<,�X<v�T<TQ<G�M<'&J<"�F<% C<�p?<��;<�Y8<x�4<�N1<]�-<�Q*<��&<jd#<!�<i�<m!<e�<�b<
<$�<�l<�&<��<pY�;��;ʙ�;DN�;��;0��;y��;���;ͫ�;X��;cԿ;D �;7<�;�;-�;�P�;�͝;![�;D��;٧�;)g�;7�;�.|;&r;�h;�5^;CyT;��J;�_A;�8;�.;��%;��;��;B�
;�H;@s�:T��:���:@Z�:��:���:>�:�Q�:.�c:��D:�`&:bK:��9��9r�?9�*�8aU����s������V��m���/���J�=�e����=���T���U���B���� �ͺt�ں�8纨��( ��c�I����������}/%�GH+��\1�/m7��y=�|�C��I���O���U���[�\�a�6�g��m�(|s�tuy�Vn�泂���������%���)���ԧ������H�������  �  6k=�
=ک=�H=��=,�=m$=U� =�_ =|��<c4�<m�<ʥ�<D��<��<~I�<~�<Ʊ�<D��<��<�E�<�t�<���<���<���<_#�<UK�<�q�<y��<���<���<@��<��<I3�<�L�<'d�<iy�<D��<���<��<��<��<���<[��<R��<���<���<���<��<���<���<~�<f�<�J�<�+�<	�<���<��<S��<�Y�<�$�<`��<<��<m�<(�<���<���<L@�<��<���< 4�<���<�l�<]�<���<$�<y��<5�<���<�6�<���<)�<�<!�<�y�<B�<II�<(��<��<jh�<���<��<�l�<��<��<�X�<袚<t�<�/�<Ys�<̴�<p��<D2�<�n�<L��<��<��<�Q�<b��< ��<&��<T#�<׫|<�y<su<��q<�7n<ڙj<��f<^c<��_<�#\<1�X<��T<'TQ<=�M<2&J<��F< C<�p?<��;<�Y8<h�4<�N1<J�-<�Q*<	�&<gd#<,�<X�<�!<\�<�b<<�<�l<�&<��<�Y�;��;���;	N�;��;$��;���;���;��;#��;gԿ;] �;�;�; ��;��;�P�;�͝;N[�;B��;ӧ�;&g�;�6�;�.|;kr;&h;
6^;LyT;��J;a_A;^8;�.;%�%;��;�;��
;�H;At�:��:���:�Z�:��:���:��:#R�:��c:F�D:�`&:TK:��9��9��?9Y�8�A����Z�������1�����O�/�q�J���e�����>��aU��GU��&B��7��A�ͺ�ںH9����,( �
d� ����������I/%�H+��\1� m7�z=��C���I�L�O�w�U�@�[�*�a�Y�g��m��{s�vuy��n����p��������?�����������2��������  �  :k=�
=�=�H=��=)�=d$=W� =�_ =���<^4�<zm�<ĥ�<=��<��<qI�<~�<���<B��<��<�E�<�t�<���<���<���<j#�<aK�<�q�<{��<���<���<8��<��<N3�<�L�<%d�<ky�<Z��<���<��<۶�<���<���<d��<e��<���<���<��<��<��<���<~�<f�<�J�<�+�<	�<���<���<Y��<�Y�<�$�<]��<>��<m�<�'�<���<���<`@�<��<���<4�<���<�l�<_�<���<$�<v��<5�<���<�6�<���<)�<圱<"�<�y�<M�<XI�<"��<��<Yh�<���<��<�l�<��<��<�X�<ܢ�<{�<�/�<Ps�<ʴ�<g��<Q2�<�n�<O��<��<��<�Q�<]��<1��</��<\#�<��|<�y<su<��q<�7n<יj<��f<^c<��_<$\<#�X<w�T<TQ<K�M<G&J<�F<  C<�p?<��;<zY8<s�4<�N1<b�-<�Q*<��&<[d#<�<e�<f!<]�<�b<<�<�l<�&<��<�Y�;��;ә�;8N�;��;-��;i��;���;ī�;g��;}Կ;S �;�;�;)��;H�;�P�;�͝;&[�;��;��;Gg�;7�;�.|;Wr;�h;�5^;cyT;��J;�_A;�8;;�.;̢%;Ƞ;�;+�
;I;>s�:%��:���:�Z�:��:���:��:�Q�:�c:\�D:�b&:"J:�9��9ڝ?9�.�8�@����_���������2��
�/���J���e�
���=��iT���U��=B��Z��6�ͺ�ں9����( ��c�c����������V/%�HH+��\1�m7��y=�v�C�׉I�b�O���U���[���a��g�Z�m�|s��uy�_n�ó��v���ĭ���������ϧ������F���*����  �  *l=�=:�=hJ=e�=�=�&=�� =|b =  =U:�<�s�<���<y��<�<�Q�<ǆ�<ں�<���<��<�P�<)��<d��<L��<��<�0�<oY�<c��<���<o��<R��<`�<�)�<�E�<�_�<x�<��<���<ݲ�<���</��<��<=��<���<���<T��<K��<,��<���<���<а�<��<p��<�j�<'L�<"*�<q�<��<׭�<�|�<�G�<��<��<I��<[L�<]�<8��<e�<��<F��<�X�<��<D��<g'�<|��<G�<�Ѻ<�W�<�ٷ<KX�<�Ҵ<�I�<ټ�<a,�<u��<�<bf�<bȩ<='�<���<�ۤ<�1�<���<՟<�"�<
n�<鶚<���<�A�<e��<�ē<q�<T@�<w{�<>��<��<�$�<^Z�<��<�<���<�'�<ʲ|<�y<�uu<b�q<O6n<5�j<5�f<5Vc<��_<
\<	zX<M�T<�AQ<ɧM<�J<�yF<c�B<�S?<��;<�88<��4<�)1<`�-<�(*<ڭ&<K7#<��<HW<e�<��<�+<��<�~<�0<��<�<=��;vm�;�;���;2��;0P�;(-�;��;��;��;�8�;$c�;���;�;C�;箢;)+�;<��;�U�;w�;�Ç;,��;��z;��p;��f;��\;�<S;��I;z)@;��6;ٓ-;{w$;�y;S�;g�	;P0;�K�:�o�:��:�S�:��:U�:�(�:��~:8�_:�JA:O�":b�:Ӡ�9g�9�}39��8��F�6�"�LM��8�������f.�^=2�YM��g�c���;���H��@��["������v�κ[ۺ���9���~ �I�����a��4��S��m%���+�r�1�&�7���=��C� �I�|�O��U���[�`�a�j�g��m�ˏs�l�y�0|�v��������'���娎�����^���s���ѣ���  �  5l=�=7�=mJ=b�=�=�&=�� =�b =���<C:�<�s�<���<���<��<�Q�<ņ�<ݺ�<���<��<�P�<��<W��<<��<��<�0�<mY�<r��<˥�<p��<J��<h�<�)�<�E�<�_�<�w�<��<���<޲�<���<,��<��<O��<���<~��<]��<:��<��<���<~��<԰�<Ϝ�<j��<�j�<,L�<**�<z�<��<ӭ�<�|�<�G�<��<��<7��<JL�<K�<A��<e�<��<V��<�X�<��<?��<m'�<x��<�G�<�Ѻ<�W�<�ٷ<CX�<�Ҵ<�I�<ټ�<q,�<���< �<bf�<gȩ<.'�<<�ۤ<�1�<���<�ԟ<�"�<n�<�<���<B�<d��<�ē<b�<<@�<�{�<3��<~�<{$�<SZ�<��<�<���<�'�<ֲ|<�y<�uu<Z�q<U6n<A�j<��f<>Vc<��_<\<zX<@�T<�AQ<��M<�J<wyF<w�B<�S?<��;<�88<{�4<�)1<8�-<�(*<ޭ&<K7#<�<_W<x�<��<�+<[�<�~<�0<��<�<���;sm�;"�;���;n��;uP�;--�;��;�;��;�8�;c�;E��;%�;C�;ﮢ;+�;.��;V�;��;ć;��;(�z;��p;<�f;z�\;}<S;��I;�(@;��6;��-;�w$;�y;��;��	;)0;�K�:1n�:���:�S�:x�:9�:�'�:+�~:��_:�KA:e�":��:���9�9}�39��8�F�	�"��P��w�������`-�6>2�LM�(�g�b���;���H���?��P#�������κ;Zۺ~������p~ �f������v4��S��m%�2�+�,�1� 7�N�=�r�C���I�гO���U���[���a�Šg���m���s�M�y�O|�h�������]������Ҩ��	���>������������  �  -l=�=3�=oJ=b�=�=�&=�� =�b =���<Q:�<�s�<���<}��<��<�Q�<���<��<���<��<�P�<��<l��<G��<��<�0�<dY�<`��<���<n��<H��<m�<�)�<�E�<�_�<�w�<���<z��<ز�<���<,��<��<<��<���<v��<e��<=��<0��<���<|��<ܰ�<ќ�<{��<�j�<*L�< *�<p�<
��<ϭ�<�|�<�G�<��<��<>��<aL�<P�<G��<e�<��<B��<�X�<��<>��<i'�<i��<�G�<�Ѻ<�W�<�ٷ<6X�<�Ҵ<�I�<ؼ�<f,�<s��<�<_f�<iȩ<5'�<��<�ۤ<�1�<���<�ԟ<�"�<�m�<춚<���<�A�<`��<�ē<r�<>@�<�{�<.��<��<�$�<TZ�<��<�<���<�'�<ʲ|<�y<�uu<E�q<I6n<R�j<��f<JVc<��_<�\<%zX<@�T<�AQ<קM<�J<eyF<��B<�S?<��;<�88<k�4<�)1<=�-<�(*<�&<>7#<�<MW<i�<p�<�+<n�<�~<�0<��<�<&��;vm�;%�;���;(��;CP�;#-�;��;�;P�;�8�;-c�;V��;K�;�B�;ծ�;+�;0��;�U�;s�;�Ç;���;f�z;�p;��f;��\;o<S;�I;�(@;�6;��-;�w$;|y;I�;��	;0;�L�:zn�:S��:�S�:��:��:�'�:��~:��_:�JA:��":��:���9��9f~39w��8��F���"�+N��K��� ����,�J>2�{M��g����p<���H���?���"��7�����κ&Zۺ<��m����} �������K��4��S��m%���+��1���7�y�=���C� �I�ʳO��U�7�[�b�a�L�g��m���s�)�y��|����g���_�������먎�8���)�������ʣ���  �  .l=�=?�=jJ=a�=�=�&=�� =~b =  =N:�<�s�<���<|��<��<�Q�<ǆ�<պ�<���<��<�P�<#��<[��<C��<��<�0�<|Y�<k��<¥�<o��<T��<a�<�)�<�E�<�_�< x�<��<���<ڲ�<���<1��<��<B��<���<���<V��<>��< ��<���<���<Ѱ�<ڜ�<k��<�j�<0L�<)*�<y�<��<ԭ�<�|�<�G�<��<��<<��<PL�<O�<;��<e�<��<I��<�X�<��<G��<h'�<���<�G�<�Ѻ<�W�<�ٷ<KX�<�Ҵ<�I�<ټ�<k,�<}��<-�<if�<^ȩ<4'�<�<�ۤ<�1�<���<�ԟ<�"�<	n�<<���<�A�<i��<�ē<k�<J@�<z{�<;��<~�<�$�<SZ�<��<�<���<�'�<̲|<�y<�uu<X�q<d6n<+�j<�f<#Vc<Ŷ_<\<zX<R�T<�AQ<ܧM<�J<�yF<l�B<�S?<��;<�88<��4<�)1<M�-<�(*<Э&<S7#<�<_W<m�<��<�+<p�<�~<�0<��<��<��;Qm�;5�;���;Q��;SP�;*-�;��;��;��;�8�;�b�;\��;��;MC�;߮�;4+�;A��;�U�;��;ć;Q��;��z;�p;k�f;��\;�<S;��I;)@;��6;��-;�w$;�y;��;��	;40;�K�:�n�:���:�S�:��:��:�'�:`�~:?�_:�LA:��":]�:n��97�9�}39���8��F�i�"�fQ��[�������:.��<2�OM�ռg����;��?H��?@���"��;����κ�Zۺ���:����~ �S�����	��4�wS��m%��+���1��7��=�o�C�]�I�γO��U�s�[��a�:�g��m���s�\�y�[|�I�������.���L�����������U���j���ƣ���  �  4l=�=7�=eJ=f�=�=�&=�� =~b =  =I:�<�s�<���<s��<��<�Q�<ֆ�<ۺ�<���<��<�P�<*��<R��<Q��<��<�0�<eY�<e��<ʥ�<d��<W��<V�<�)�<�E�<�_�<x�<ۍ�<���<ʲ�<���<%��<
��<H��<���<��<R��<O��<"��<���<���<Ͱ�<ޜ�<i��<�j�<'L�<#*�<v�<��<��<�|�<�G�<��<$��<B��<NL�<b�<9��<e�<��<K��<�X�<��<E��<V'�<���<~G�<�Ѻ<�W�<�ٷ<IX�<�Ҵ<�I�<˼�<p,�<x��<�<Zf�<bȩ<D'�<낦<�ۤ<�1�<���< ՟<�"�<n�<ᶚ<���<�A�<k��<�ē<f�<L@�<x{�<D��<|�<�$�<_Z�<��<�<���<�'�<Ų|<�y<�uu<F�q<m6n<"�j<1�f< Vc<̶_<�\<zX<O�T<�AQ<�M<�J<uyF<V�B<�S?<��;<�88<��4<�)1<N�-<�(*<�&<`7#<��<kW<Z�<��<�+<s�<�~<�0<��<�<R��;om�;��;���;<��;qP�;�,�;��;��;��;�8�;�b�;���;��;]C�;���;!+�;��;�U�;��;�Ç;��;��z;��p;y�f;��\;�<S;w�I;.)@;~�6;)�-;~w$;�y;}�;N�	;�0;�K�:Mo�:���:XT�:(�:��:)�:%�~:y�_:7JA:�":��:[��9��9Qu39K��8��F�ק"��O��E���]����/�<2�M�?�g�3���<��2I��@���!������z�κfZۺP������~ �Ĵ�8�����4�kS�{m%��+���1�#�7�̩=���C�)�I�r�O�C�U��[�Y�a��g��m��s���y��|�8���Ǵ������R����������m���o���棚��  �  /l=�=8�=pJ=a�=�=�&=�� =�b =  =N:�<�s�<���<{��<��<�Q�<ņ�<��<���<��<�P�<��<a��<B��<��<�0�<lY�<d��<å�<e��<Q��<n�<�)�<�E�<�_�<x�<��<���<ײ�<���<&��<��<>��<���<���<d��<<��<!��<���<|��<װ�<֜�<s��<�j�<'L�<)*�<z�<��<ڭ�<�|�<�G�<��<��<9��<RL�<M�<E��<e�<��<D��<�X�<��<M��<g'�<t��<�G�<�Ѻ<�W�<�ٷ<;X�<�Ҵ<�I�<ϼ�<l,�<v��<�<if�<eȩ<1'�<���<�ۤ<�1�<���<�ԟ<�"�<
n�<㶚<���<�A�<b��<�ē<m�<F@�<�{�</��<��<�$�<QZ�<��<�<���<�'�<Ȳ|<�y<�uu<J�q<V6n<7�j<�f</Vc<��_<�\<-zX<C�T<�AQ<ߧM<�J<{yF<��B<�S?<��;<�88<p�4<�)1<I�-<�(*<�&<F7#<�<iW<^�<��<�+<o�<�~<�0<��<�<��;nm�;E�;���;9��;VP�;-�;��;�;`�;�8�;c�;_��;�; C�;Ѯ�;S+�;��;V�;~�;�Ç;-��;e�z;�p;q�f;��\;l<S;̢I;�(@;��6;��-;{w$;�y;��;]�	;i0;<L�:�n�:'��:�S�:��:��:�'�:��~:n�_:{KA:%�":��:m��9��9�}39��8��F���"�{P���������� -��<2��M���g�R���;��BH���?��"#��������κbZۺD��B���.~ �F��-�����4��S��m%�Ղ+��1���7�p�=�8�C�o�I��O�w�U��[�P�a�7�g���m��s��y��|�f�������?���3���ը��1����������ᣚ��  �  ,l=�=5�=nJ=d�=�=�&=�� =�b =���<Q:�<�s�<���<���<~�<�Q�<���<��<���<��<�P�<��<k��<<��<��<�0�<lY�<m��<���<w��<A��<i�<�)�<�E�<�_�<�w�<��<���<ٲ�<���<%��<��<:��<���<u��<e��<=��<)��<���<���<��<͜�<{��<�j�<2L�<"*�<p�<��<ҭ�<�|�<�G�<��<!��<8��<]L�<L�<H��<e�<��<B��<�X�<��<9��<j'�<r��<�G�<�Ѻ<�W�<�ٷ<9X�<�Ҵ<�I�<߼�<i,�<z��< �<^f�<mȩ<,'�<��<�ۤ<�1�<���<�ԟ<�"�<n�<���<���<B�<h��<�ē<s�<8@�<�{�<2��<��<�$�<WZ�<��<�<���<�'�<�|<�y<�uu<K�q<Q6n<F�j<��f<:Vc<��_<�\<zX<0�T<�AQ<ҧM<�J<kyF<z�B<�S?<��;<�88<u�4<�)1<1�-<�(*<߭&<M7#<�<HW<��<z�<�+<l�<�~<�0<��<�<���;�m�;$�;���;\��;EP�;H-�;��;�;Z�;�8�;c�;;��;/�;C�;ۮ�;+�;��;V�;o�;-ć;���;h�z;�p;��f;��\;�<S;�I;�(@;�6;��-;�w$;�y;K�;��	;#0;�L�:>n�:o��:(T�:��:z�:�'�:�~:��_:�LA:��":��:|��9���9!39˩�8!�F��"�dQ������H���K-��>2�~M��g����;���H��H?��o#��8�����κ�Yۺ��纕���-~ �~�����b�|4��S��m%���+�O�1�q�7�U�=��C�W�I���O���U�0�[�ӧa�d�g���m�7�s�V�y��|�p������^������ը��+���@������������  �  +l=�=6�=jJ=g�=�=�&=�� =�b =   =Z:�<�s�<���<���<��<�Q�<ņ�<��<���<��<�P�<��<Z��<G��<��<�0�<hY�<h��<���<m��<O��<b�<�)�<�E�<�_�<x�<ٍ�<���<ز�<���<)��<	��<;��<���<x��<]��<I��<&��<���<���<Ұ�<ޜ�<z��<�j�<-L�<&*�<w�<��<ҭ�<�|�<�G�<��<!��<8��<VL�<Y�<C��<e�<��<C��<�X�<
��<C��<e'�<{��<{G�<�Ѻ<�W�<�ٷ<CX�<�Ҵ<�I�<ռ�<c,�<y��<�<\f�<oȩ<9'�<�<�ۤ<�1�<���<	՟<�"�<n�<�<���<B�<f��<�ē<z�<G@�<|{�<7��<��<�$�<^Z�<��<�<���<�'�<Ͳ|<�y<�uu<K�q<V6n<"�j<�f< Vc<��_<�\<zX<E�T<�AQ<ͧM<�J<ryF<k�B<�S?<��;<�88<��4<�)1<G�-<�(*<ܭ&<K7#<�<XW<v�<��<�+<��<�~<�0<��<��<+��;�m�;�;���;G��;6P�;%-�;��;��;��;�8�;�b�;v��;��;0C�;خ�;"+�;#��;�U�;s�;ć;��;+�z;r�p;��f;��\;�<S;��I;/)@;
�6;��-;�w$;�y;��;��	;*0;oL�:io�:���:0T�:��:�:�(�:t�~:��_:?KA:�":�:3��9.�9�|39���8��F���"�P��"�������G.��=2��M�νg�$��E<��I��1?���"��D���O�κ5Zۺv��q��=~ �]�������4��S��m%�t�+�ד1���7�/�=�U�C�J�I�w�O�رU��[�"�a�t�g��m��s�U�y��|�f���Ǵ�����R���ۨ��!���J�������ˣ���  �  7l=�=<�=nJ=\�=�=�&=�� =�b =  =D:�<�s�<���<{��<��<�Q�<ц�<ݺ�<���<��<�P�<'��<Y��<E��<��<�0�<oY�<a��<Υ�<`��<V��<Z�<�)�<�E�<�_�<x�<؍�<���<β�<���<'��<
��<J��<���<���<W��<<��<��<���<���<Ͱ�<ߜ�<e��<�j�<*L�<,*�<��<��<��<�|�<�G�<��<!��<>��<KL�<P�<:��<e�<��<N��<�X�<��<J��<['�<���<yG�<�Ѻ<�W�<�ٷ<HX�<�Ҵ<�I�<ɼ�<r,�<x��<�<nf�<Yȩ<7'�<<�ۤ<�1�<���<�ԟ<�"�<n�<嶚<���<�A�<j��<�ē<b�<N@�<|{�<>��<��<�$�<KZ�<��<�<���<�'�<��|<�y<�uu<>�q<w6n<�j<!�f<Vc<Ӷ_<�\<zX<J�T<�AQ<��M<�J<�yF<}�B<�S?<��;<�88<��4<�)1<V�-<�(*<�&<[7#<�<yW<_�<��<�+<e�<�~<�0<��<�<"��;4m�;O�;���;-��;�P�;�,�;��;��;��;�8�;�b�;n��;��;mC�;���;;+�;��; V�;��;�Ç;T��;��z;�p;G�f;��\;�<S;~�I;1)@;`�6;,�-;�w$;�y;Ι;r�	;�0;\K�:o�:���:6T�:��:[�:�'�:H�~:��_:cJA:e�":��:���9��9�w390��8��F���"��Q������w���/��<2�2M��g�,��<���G���@���"��������κ`Zۺx��]����~ ��������4�sS�nm%�3�+���1��7���=�N�C�s�I��O���U���[���a� g��m��s�R�y��|�#���մ�����l�������+���T���z�����  �  1l=�=6�=iJ=b�=�=�&=�� =�b =  =K:�<�s�<���<{��<��<�Q�<̆�<��<���<��<�P�<��<e��<T��<��<�0�<iY�<b��<ť�<d��<T��<`�<�)�<�E�<�_�<x�<��<���<Ȳ�<���<$��<��<D��<���<|��<V��<J��<2��<���<���<۰�<ݜ�<s��<�j�<*L�<$*�<t�<	��<��<�|�<�G�<��< ��<>��<`L�<^�<;��<e�<��<H��<�X�<��<C��<X'�<t��<�G�<�Ѻ<�W�<�ٷ<9X�<�Ҵ<�I�<μ�<j,�<t��<�<^f�<_ȩ<D'�<���<�ۤ<�1�<���<�ԟ<�"�<n�<붚<���<�A�<h��<�ē<j�<J@�<�{�<6��<��<�$�<XZ�<��<�<���<�'�<��|<�y<�uu<2�q<[6n<-�j<�f<#Vc<��_<�\<zX<G�T<�AQ<�M<�J<syF<g�B<�S?<��;<�88<~�4<�)1<S�-<�(*<��&<T7#<�<`W<j�<��<�+<p�<�~<�0<��<�<_��;`m�;�;���;1��;aP�;�,�;��;��;Y�;�8�;�b�;h��;�;"C�;���;$+�;��;�U�;��;�Ç;��;��z;z�p;�f;��\;�<S;�I;%)@;��6;1�-;�w$;�y;n�;{�	;�0;dL�:&o�:s��:T�:��:��:�(�:y�~:D�_:�JA:��":��:���9E�9+v39d��82�F���"�#P�����)���/�=2��M���g�g��><���H��+@���!�������κyZۺ������~ �
�������4�}S�Am%��+���1���7�7�=�!�C�˲I���O��U���[�W�a��g�*�m��s�N�y��|�[�������1���K���Ũ��Q���I������񣚻�  �  *l=�=:�=kJ=f�=�=�&=�� =�b =���<W:�<�s�<���<���<�<�Q�<���<��<���<��<�P�<��<Y��<;��<��<�0�<sY�<o��<���<r��<G��<h�<�)�<�E�<�_�<�w�<��<~��<��<���<+��<��<<��<���<|��<a��<=��<��<���<}��<ڰ�<ќ�<|��<�j�<5L�<.*�<{�<��<ɭ�<�|�<�G�<��<��<6��<ML�<M�<F��<e�<��<G��<�X�<��<=��<n'�<n��<�G�<�Ѻ<�W�<�ٷ<;X�<�Ҵ<�I�<ڼ�<c,�<��<'�<]f�<nȩ<-'�<���<�ۤ<�1�<���<�ԟ<�"�<�m�<���<���<B�<e��<�ē<w�<?@�<�{�<3��<}�<~$�<XZ�<��<�<���<�'�<ֲ|<�y<�uu<X�q<D6n<*�j<�f<&Vc<��_<�\<zX<;�T<�AQ<ɧM<�J<�yF<p�B<�S?<��;<�88<y�4<�)1<A�-<�(*<ح&<C7#<)�<JW<��<s�<�+<w�<�~<�0<��<�<���;�m�;�;���;e��;3P�;5-�;��;�;t�;�8�;�b�;G��;�;C�;���;+�;+��;V�;x�;2ć;��;J�z;�p;V�f;w�\;z<S;�I;�(@;�6;��-;�w$;�y;��;��	;�/;�L�:�n�:L��:�S�:u�:z�:�'�:��~:?�_:	MA:��":�:ß�9��9��39G��8��F���"��Q����������`-�N>2�M�νg����T;���H��C?��W#��m���q�κ�Zۺ ��;���8~ ����F��;�-4��S��m%���+��1���7�Q�=�s�C���I���O�ǱU�֭[�ʧa���g���m��s�W�y�W|���������T���E���𨎻���B������������  �  .l=�=3�=lJ=c�=�=�&=�� =�b =���<R:�<�s�<���<���<�<�Q�<Æ�<��<���<��<�P�<,��<e��<D��<��<�0�<aY�<a��<���<m��<E��<W�<�)�<�E�<�_�<x�<��<���<в�<���<&��<
��<;��<���<v��<^��<B��<'��<���<���<۰�<Ҝ�<{��<�j�</L�<%*�<s�<��<׭�<�|�<�G�<��<$��<J��<WL�<T�<A��<e�<��<B��<�X�<��<7��<\'�<s��<�G�<�Ѻ<�W�<�ٷ<;X�<�Ҵ<�I�<Ӽ�<f,�<s��<�<Zf�<fȩ<5'�<���<�ۤ<�1�<���<�ԟ<�"�<n�<���<���<B�<e��<�ē<s�<@@�<�{�<A��<��<�$�<VZ�<��<�<���<�'�<Ӳ|<�y<�uu<C�q<W6n<:�j<�f<3Vc<��_<�\<�yX<7�T<�AQ<اM<�J<eyF<r�B<�S?<��;<�88<��4<�)1<B�-<�(*<�&<L7#<�<JW<��<�<�+<p�<�~<�0<��<�<��;ym�;�;���;,��;FP�;#-�;��;��;g�;�8�;c�;j��;�;C�;���;�*�;��;�U�;s�;�Ç;���;2�z;;�p;��f;�\;�<S;�I;�(@;�6;�-;�w$;�y;i�;��	;T0;�L�:�n�:_��:aT�:��:�:?(�:>�~:��_:JA:��":�:=��9:��9�x39���8��F�ǫ"��O��?�������p/��>2�M�q�g�����<��-I���?���"������@�κZۺ*��R����} �r�����T�h4��S�xm%���+��1���7��=��C�>�I���O�űU�1�[�n�a�O�g�˘m��s���y��|�d�������-���*���Ө��1���u�������ȣ���  �  4l=�=:�=nJ=_�=�=�&=�� =�b =  =J:�<�s�<���<���<��<�Q�<���<��<���<��<�P�<��<X��<L��<��<�0�<qY�<n��<ȥ�<a��<]��<d�<�)�<�E�<�_�<�w�<���<���<ϲ�<���<-��<��<M��<���<���<W��<A��<#��<���<y��<ܰ�<؜�<s��<�j�<'L�<4*�<��<��<ݭ�<�|�<�G�<��<��<:��<OL�<V�<8��<e�<��<T��<�X�<��<U��<]'�<x��<G�<�Ѻ<�W�<�ٷ<?X�<�Ҵ<�I�<˼�<m,�<���<$�<kf�<]ȩ<<'�<���<�ۤ<�1�<���<�ԟ<�"�<n�<�<���<	B�<_��<�ē<k�<I@�<�{�<-��<�<�$�<QZ�<��<�<���<�'�<��|<�y<�uu<;�q<[6n<&�j<��f<Vc<��_<�\<$zX<Y�T<�AQ<�M<�J<�yF<|�B<�S?<��;<�88<k�4<�)1<P�-<�(*<��&<A7#<�<�W<r�<x�<�+<n�<�~<�0<��<�<=��;Um�;K�;���;b��;lP�;�,�;�;��;u�;�8�;�b�;=��;��;+C�;���;h+�;5��;�U�;��;ć;;��;��z;6�p;��f;��\;V<S;�I; )@;��6;�-;�w$;z;�;q�	;0;RL�:�n�:���:�S�:��:��:T(�:�~:��_:LA:-�":��:`��9��9y39���8 �F�j�"��Q���������p.��;2�M���g�����;��H��F@��q"��c���n�κ�Zۺ���$��� ~ �z�������L4��S�.m%��+�Ǔ1���7�|�=�g�C�0�I��O���U���[��a�ؠg�]�m�Əs���y��|�\�������^���W���Ш��>���*���[�������  �  .l=�=3�=lJ=c�=�=�&=�� =�b =���<R:�<�s�<���<���<�<�Q�<Æ�<��<���<��<�P�<,��<e��<D��<��<�0�<aY�<a��<���<m��<E��<W�<�)�<�E�<�_�<x�<��<���<в�<���<&��<
��<;��<���<v��<^��<B��<'��<���<���<۰�<Ҝ�<{��<�j�</L�<%*�<s�<��<׭�<�|�<�G�<��<$��<J��<WL�<T�<A��<e�<��<B��<�X�<��<7��<\'�<s��<�G�<�Ѻ<�W�<�ٷ<;X�<�Ҵ<�I�<Ӽ�<f,�<s��<�<Zf�<fȩ<5'�<���<�ۤ<�1�<���<�ԟ<�"�<n�<���<���<B�<e��<�ē<s�<@@�<�{�<A��<��<�$�<VZ�<��<�<���<�'�<Ӳ|<�y<�uu<C�q<W6n<:�j<�f<3Vc<��_<�\<�yX<7�T<�AQ<اM<�J<eyF<r�B<�S?<��;<�88<��4<�)1<B�-<�(*<�&<L7#<�<JW<��<�<�+<p�<�~<�0<��<�<��;ym�;�;���;,��;FP�;#-�;��;��;g�;�8�;c�;j��;�;C�;���;�*�;��;�U�;s�;�Ç;���;2�z;;�p;��f;�\;�<S;�I;�(@;�6;�-;�w$;�y;i�;��	;T0;�L�:�n�:_��:aT�:��:�:?(�:>�~:��_:JA:��":�:=��9:��9�x39���8��F�ǫ"��O��?�������p/��>2�M�q�g�����<��-I���?���"������@�κZۺ*��R����} �r�����T�h4��S�xm%���+��1���7��=��C�>�I���O�űU�1�[�n�a�O�g�˘m��s���y��|�d�������-���*���Ө��1���u�������ȣ���  �  *l=�=:�=kJ=f�=�=�&=�� =�b =���<W:�<�s�<���<���<�<�Q�<���<��<���<��<�P�<��<Y��<;��<��<�0�<sY�<o��<���<r��<G��<h�<�)�<�E�<�_�<�w�<��<~��<��<���<+��<��<<��<���<|��<a��<=��<��<���<}��<ڰ�<ќ�<|��<�j�<5L�<.*�<{�<��<ɭ�<�|�<�G�<��<��<6��<ML�<M�<F��<e�<��<G��<�X�<��<=��<n'�<n��<�G�<�Ѻ<�W�<�ٷ<;X�<�Ҵ<�I�<ڼ�<c,�<��<'�<]f�<nȩ<-'�<���<�ۤ<�1�<���<�ԟ<�"�<�m�<���<���<B�<e��<�ē<w�<?@�<�{�<3��<}�<~$�<XZ�<��<�<���<�'�<ֲ|<�y<�uu<X�q<D6n<*�j<�f<&Vc<��_<�\<zX<;�T<�AQ<ɧM<�J<�yF<p�B<�S?<��;<�88<y�4<�)1<A�-<�(*<ح&<C7#<)�<JW<��<s�<�+<w�<�~<�0<��<�<���;�m�;�;���;e��;3P�;5-�;��;�;t�;�8�;�b�;G��;�;C�;���;+�;+��;V�;x�;2ć;��;J�z;�p;V�f;w�\;z<S;�I;�(@;�6;��-;�w$;�y;��;��	;�/;�L�:�n�:L��:�S�:u�:z�:�'�:��~:?�_:	MA:��":�:ß�9��9��39G��8��F���"��Q����������`-�N>2�M�νg����T;���H��C?��W#��m���q�κ�Zۺ ��;���8~ ����F��;�-4��S��m%���+��1���7�Q�=�s�C���I���O�ǱU�֭[�ʧa���g���m��s�W�y�W|���������T���E���𨎻���B������������  �  1l=�=6�=iJ=b�=�=�&=�� =�b =  =K:�<�s�<���<{��<��<�Q�<̆�<��<���<��<�P�<��<e��<T��<��<�0�<iY�<b��<ť�<d��<T��<`�<�)�<�E�<�_�<x�<��<���<Ȳ�<���<$��<��<D��<���<|��<V��<J��<2��<���<���<۰�<ݜ�<s��<�j�<*L�<$*�<t�<	��<��<�|�<�G�<��< ��<>��<`L�<^�<;��<e�<��<H��<�X�<��<C��<X'�<t��<�G�<�Ѻ<�W�<�ٷ<9X�<�Ҵ<�I�<μ�<j,�<t��<�<^f�<_ȩ<D'�<���<�ۤ<�1�<���<�ԟ<�"�<n�<붚<���<�A�<h��<�ē<j�<J@�<�{�<6��<��<�$�<XZ�<��<�<���<�'�<��|<�y<�uu<2�q<[6n<-�j<�f<#Vc<��_<�\<zX<G�T<�AQ<�M<�J<syF<g�B<�S?<��;<�88<~�4<�)1<S�-<�(*<��&<T7#<�<`W<j�<��<�+<p�<�~<�0<��<�<_��;`m�;�;���;1��;aP�;�,�;��;��;Y�;�8�;�b�;h��;�;"C�;���;$+�;��;�U�;��;�Ç;��;��z;z�p;�f;��\;�<S;�I;%)@;��6;1�-;�w$;�y;n�;{�	;�0;dL�:&o�:s��:T�:��:��:�(�:y�~:D�_:�JA:��":��:���9E�9+v39d��82�F���"�#P�����)���/�=2��M���g�g��><���H��+@���!�������κyZۺ������~ �
�������4�}S�Am%��+���1���7�7�=�!�C�˲I���O��U���[�W�a��g�*�m��s�N�y��|�[�������1���K���Ũ��Q���I������񣚻�  �  7l=�=<�=nJ=\�=�=�&=�� =�b =  =D:�<�s�<���<{��<��<�Q�<ц�<ݺ�<���<��<�P�<'��<Y��<E��<��<�0�<oY�<a��<Υ�<`��<V��<Z�<�)�<�E�<�_�<x�<؍�<���<β�<���<'��<
��<J��<���<���<W��<<��<��<���<���<Ͱ�<ߜ�<e��<�j�<*L�<,*�<��<��<��<�|�<�G�<��<!��<>��<KL�<P�<:��<e�<��<N��<�X�<��<J��<['�<���<yG�<�Ѻ<�W�<�ٷ<HX�<�Ҵ<�I�<ɼ�<r,�<x��<�<nf�<Yȩ<7'�<<�ۤ<�1�<���<�ԟ<�"�<n�<嶚<���<�A�<j��<�ē<b�<N@�<|{�<>��<��<�$�<KZ�<��<�<���<�'�<��|<�y<�uu<>�q<w6n<�j<!�f<Vc<Ӷ_<�\<zX<J�T<�AQ<��M<�J<�yF<}�B<�S?<��;<�88<��4<�)1<V�-<�(*<�&<[7#<�<yW<_�<��<�+<e�<�~<�0<��<�<"��;4m�;O�;���;-��;�P�;�,�;��;��;��;�8�;�b�;n��;��;mC�;���;;+�;��; V�;��;�Ç;T��;��z;�p;G�f;��\;�<S;~�I;1)@;`�6;,�-;�w$;�y;Ι;r�	;�0;\K�:o�:���:6T�:��:[�:�'�:H�~:��_:cJA:e�":��:���9��9�w390��8��F���"��Q������w���/��<2�2M��g�,��<���G���@���"��������κ`Zۺx��]����~ ��������4�sS�nm%�3�+���1��7���=�N�C�s�I��O���U���[���a� g��m��s�R�y��|�#���մ�����l�������+���T���z�����  �  +l=�=6�=jJ=g�=�=�&=�� =�b =   =Z:�<�s�<���<���<��<�Q�<ņ�<��<���<��<�P�<��<Z��<G��<��<�0�<hY�<h��<���<m��<O��<b�<�)�<�E�<�_�<x�<ٍ�<���<ز�<���<)��<	��<;��<���<x��<]��<I��<&��<���<���<Ұ�<ޜ�<z��<�j�<-L�<&*�<w�<��<ҭ�<�|�<�G�<��<!��<8��<VL�<Y�<C��<e�<��<C��<�X�<
��<C��<e'�<{��<{G�<�Ѻ<�W�<�ٷ<CX�<�Ҵ<�I�<ռ�<c,�<y��<�<\f�<oȩ<9'�<�<�ۤ<�1�<���<	՟<�"�<n�<�<���<B�<f��<�ē<z�<G@�<|{�<7��<��<�$�<^Z�<��<�<���<�'�<Ͳ|<�y<�uu<K�q<V6n<"�j<�f< Vc<��_<�\<zX<E�T<�AQ<ͧM<�J<ryF<k�B<�S?<��;<�88<��4<�)1<G�-<�(*<ܭ&<K7#<�<XW<v�<��<�+<��<�~<�0<��<��<+��;�m�;�;���;G��;6P�;%-�;��;��;��;�8�;�b�;v��;��;0C�;خ�;"+�;#��;�U�;s�;ć;��;+�z;r�p;��f;��\;�<S;��I;/)@;
�6;��-;�w$;�y;��;��	;*0;oL�:io�:���:0T�:��:�:�(�:t�~:��_:?KA:�":�:3��9.�9�|39���8��F���"�P��"�������G.��=2��M�νg�$��E<��I��1?���"��D���O�κ5Zۺv��q��=~ �]�������4��S��m%�t�+�ד1���7�/�=�U�C�J�I�w�O�رU��[�"�a�t�g��m��s�U�y��|�f���Ǵ�����R���ۨ��!���J�������ˣ���  �  ,l=�=5�=nJ=d�=�=�&=�� =�b =���<Q:�<�s�<���<���<~�<�Q�<���<��<���<��<�P�<��<k��<<��<��<�0�<lY�<m��<���<w��<A��<i�<�)�<�E�<�_�<�w�<��<���<ٲ�<���<%��<��<:��<���<u��<e��<=��<)��<���<���<��<͜�<{��<�j�<2L�<"*�<p�<��<ҭ�<�|�<�G�<��<!��<8��<]L�<L�<H��<e�<��<B��<�X�<��<9��<j'�<r��<�G�<�Ѻ<�W�<�ٷ<9X�<�Ҵ<�I�<߼�<i,�<z��< �<^f�<mȩ<,'�<��<�ۤ<�1�<���<�ԟ<�"�<n�<���<���<B�<h��<�ē<s�<8@�<�{�<2��<��<�$�<WZ�<��<�<���<�'�<�|<�y<�uu<K�q<Q6n<F�j<��f<:Vc<��_<�\<zX<0�T<�AQ<ҧM<�J<kyF<z�B<�S?<��;<�88<u�4<�)1<1�-<�(*<߭&<M7#<�<HW<��<z�<�+<l�<�~<�0<��<�<���;�m�;$�;���;\��;EP�;H-�;��;�;Z�;�8�;c�;;��;/�;C�;ۮ�;+�;��;V�;o�;-ć;���;h�z;�p;��f;��\;�<S;�I;�(@;�6;��-;�w$;�y;K�;��	;#0;�L�:>n�:o��:(T�:��:z�:�'�:�~:��_:�LA:��":��:|��9���9!39˩�8!�F��"�dQ������H���K-��>2�~M��g����;���H��H?��o#��8�����κ�Yۺ��纕���-~ �~�����b�|4��S��m%���+�O�1�q�7�U�=��C�W�I���O���U�0�[�ӧa�d�g���m�7�s�V�y��|�p������^������ը��+���@������������  �  /l=�=8�=pJ=a�=�=�&=�� =�b =  =N:�<�s�<���<{��<��<�Q�<ņ�<��<���<��<�P�<��<a��<B��<��<�0�<lY�<d��<å�<e��<Q��<n�<�)�<�E�<�_�<x�<��<���<ײ�<���<&��<��<>��<���<���<d��<<��<!��<���<|��<װ�<֜�<s��<�j�<'L�<)*�<z�<��<ڭ�<�|�<�G�<��<��<9��<RL�<M�<E��<e�<��<D��<�X�<��<M��<g'�<t��<�G�<�Ѻ<�W�<�ٷ<;X�<�Ҵ<�I�<ϼ�<l,�<v��<�<if�<eȩ<1'�<���<�ۤ<�1�<���<�ԟ<�"�<
n�<㶚<���<�A�<b��<�ē<m�<F@�<�{�</��<��<�$�<QZ�<��<�<���<�'�<Ȳ|<�y<�uu<J�q<V6n<7�j<�f</Vc<��_<�\<-zX<C�T<�AQ<ߧM<�J<{yF<��B<�S?<��;<�88<p�4<�)1<I�-<�(*<�&<F7#<�<iW<^�<��<�+<o�<�~<�0<��<�<��;nm�;E�;���;9��;VP�;-�;��;�;`�;�8�;c�;_��;�; C�;Ѯ�;S+�;��;V�;~�;�Ç;-��;e�z;�p;q�f;��\;l<S;̢I;�(@;��6;��-;{w$;�y;��;]�	;i0;<L�:�n�:'��:�S�:��:��:�'�:��~:n�_:{KA:%�":��:m��9��9�}39��8��F���"�{P���������� -��<2��M���g�R���;��BH���?��"#��������κbZۺD��B���.~ �F��-�����4��S��m%�Ղ+��1���7�p�=�8�C�o�I��O�w�U��[�P�a�7�g���m��s��y��|�f�������?���3���ը��1����������ᣚ��  �  4l=�=7�=eJ=f�=�=�&=�� =~b =  =I:�<�s�<���<s��<��<�Q�<ֆ�<ۺ�<���<��<�P�<*��<R��<Q��<��<�0�<eY�<e��<ʥ�<d��<W��<V�<�)�<�E�<�_�<x�<ۍ�<���<ʲ�<���<%��<
��<H��<���<��<R��<O��<"��<���<���<Ͱ�<ޜ�<i��<�j�<'L�<#*�<v�<��<��<�|�<�G�<��<$��<B��<NL�<b�<9��<e�<��<K��<�X�<��<E��<V'�<���<~G�<�Ѻ<�W�<�ٷ<IX�<�Ҵ<�I�<˼�<p,�<x��<�<Zf�<bȩ<D'�<낦<�ۤ<�1�<���< ՟<�"�<n�<ᶚ<���<�A�<k��<�ē<f�<L@�<x{�<D��<|�<�$�<_Z�<��<�<���<�'�<Ų|<�y<�uu<F�q<m6n<"�j<1�f< Vc<̶_<�\<zX<O�T<�AQ<�M<�J<uyF<V�B<�S?<��;<�88<��4<�)1<N�-<�(*<�&<`7#<��<kW<Z�<��<�+<s�<�~<�0<��<�<R��;om�;��;���;<��;qP�;�,�;��;��;��;�8�;�b�;���;��;]C�;���;!+�;��;�U�;��;�Ç;��;��z;��p;y�f;��\;�<S;w�I;.)@;~�6;)�-;~w$;�y;}�;N�	;�0;�K�:Mo�:���:XT�:(�:��:)�:%�~:y�_:7JA:�":��:[��9��9Qu39K��8��F�ק"��O��E���]����/�<2�M�?�g�3���<��2I��@���!������z�κfZۺP������~ �Ĵ�8�����4�kS�{m%��+���1�#�7�̩=���C�)�I�r�O�C�U��[�Y�a��g��m��s���y��|�8���Ǵ������R����������m���o���棚��  �  .l=�=?�=jJ=a�=�=�&=�� =~b =  =N:�<�s�<���<|��<��<�Q�<ǆ�<պ�<���<��<�P�<#��<[��<C��<��<�0�<|Y�<k��<¥�<o��<T��<a�<�)�<�E�<�_�< x�<��<���<ڲ�<���<1��<��<B��<���<���<V��<>��< ��<���<���<Ѱ�<ڜ�<k��<�j�<0L�<)*�<y�<��<ԭ�<�|�<�G�<��<��<<��<PL�<O�<;��<e�<��<I��<�X�<��<G��<h'�<���<�G�<�Ѻ<�W�<�ٷ<KX�<�Ҵ<�I�<ټ�<k,�<}��<-�<if�<^ȩ<4'�<�<�ۤ<�1�<���<�ԟ<�"�<	n�<<���<�A�<i��<�ē<k�<J@�<z{�<;��<~�<�$�<SZ�<��<�<���<�'�<̲|<�y<�uu<X�q<d6n<+�j<�f<#Vc<Ŷ_<\<zX<R�T<�AQ<ܧM<�J<�yF<l�B<�S?<��;<�88<��4<�)1<M�-<�(*<Э&<S7#<�<_W<m�<��<�+<p�<�~<�0<��<��<��;Qm�;5�;���;Q��;SP�;*-�;��;��;��;�8�;�b�;\��;��;MC�;߮�;4+�;A��;�U�;��;ć;Q��;��z;�p;k�f;��\;�<S;��I;)@;��6;��-;�w$;�y;��;��	;40;�K�:�n�:���:�S�:��:��:�'�:`�~:?�_:�LA:��":]�:n��97�9�}39���8��F�i�"�fQ��[�������:.��<2�OM�ռg����;��?H��?@���"��;����κ�Zۺ���:����~ �S�����	��4�wS��m%��+���1��7��=�o�C�]�I�γO��U�s�[��a�:�g��m���s�\�y�[|�I�������.���L�����������U���j���ƣ���  �  -l=�=3�=oJ=b�=�=�&=�� =�b =���<Q:�<�s�<���<}��<��<�Q�<���<��<���<��<�P�<��<l��<G��<��<�0�<dY�<`��<���<n��<H��<m�<�)�<�E�<�_�<�w�<���<z��<ز�<���<,��<��<<��<���<v��<e��<=��<0��<���<|��<ܰ�<ќ�<{��<�j�<*L�< *�<p�<
��<ϭ�<�|�<�G�<��<��<>��<aL�<P�<G��<e�<��<B��<�X�<��<>��<i'�<i��<�G�<�Ѻ<�W�<�ٷ<6X�<�Ҵ<�I�<ؼ�<f,�<s��<�<_f�<iȩ<5'�<��<�ۤ<�1�<���<�ԟ<�"�<�m�<춚<���<�A�<`��<�ē<r�<>@�<�{�<.��<��<�$�<TZ�<��<�<���<�'�<ʲ|<�y<�uu<E�q<I6n<R�j<��f<JVc<��_<�\<%zX<@�T<�AQ<קM<�J<eyF<��B<�S?<��;<�88<k�4<�)1<=�-<�(*<�&<>7#<�<MW<i�<p�<�+<n�<�~<�0<��<�<&��;vm�;%�;���;(��;CP�;#-�;��;�;P�;�8�;-c�;V��;K�;�B�;ծ�;+�;0��;�U�;s�;�Ç;���;f�z;�p;��f;��\;o<S;�I;�(@;�6;��-;�w$;|y;I�;��	;0;�L�:zn�:S��:�S�:��:��:�'�:��~:��_:�JA:��":��:���9��9f~39w��8��F���"�+N��K��� ����,�J>2�{M��g����p<���H���?���"��7�����κ&Zۺ<��m����} �������K��4��S��m%���+��1���7�y�=���C� �I�ʳO��U�7�[�b�a�L�g��m���s�)�y��|����g���_�������먎�8���)�������ʣ���  �  5l=�=7�=mJ=b�=�=�&=�� =�b =���<C:�<�s�<���<���<��<�Q�<ņ�<ݺ�<���<��<�P�<��<W��<<��<��<�0�<mY�<r��<˥�<p��<J��<h�<�)�<�E�<�_�<�w�<��<���<޲�<���<,��<��<O��<���<~��<]��<:��<��<���<~��<԰�<Ϝ�<j��<�j�<,L�<**�<z�<��<ӭ�<�|�<�G�<��<��<7��<JL�<K�<A��<e�<��<V��<�X�<��<?��<m'�<x��<�G�<�Ѻ<�W�<�ٷ<CX�<�Ҵ<�I�<ټ�<q,�<���< �<bf�<gȩ<.'�<<�ۤ<�1�<���<�ԟ<�"�<n�<�<���<B�<d��<�ē<b�<<@�<�{�<3��<~�<{$�<SZ�<��<�<���<�'�<ֲ|<�y<�uu<Z�q<U6n<A�j<��f<>Vc<��_<\<zX<@�T<�AQ<��M<�J<wyF<w�B<�S?<��;<�88<{�4<�)1<8�-<�(*<ޭ&<K7#<�<_W<x�<��<�+<[�<�~<�0<��<�<���;sm�;"�;���;n��;uP�;--�;��;�;��;�8�;c�;E��;%�;C�;ﮢ;+�;.��;V�;��;ć;��;(�z;��p;<�f;z�\;}<S;��I;�(@;��6;��-;�w$;�y;��;��	;)0;�K�:1n�:���:�S�:x�:9�:�'�:+�~:��_:�KA:e�":��:���9�9}�39��8�F�	�"��P��w�������`-�6>2�LM�(�g�b���;���H���?��P#�������κ;Zۺ~������p~ �f������v4��S��m%�2�+�,�1� 7�N�=�r�C���I�гO���U���[���a�Šg���m���s�M�y�O|�h�������]������Ҩ��	���>������������  �  >m==��=L=H�=5�=�(=9� =Ae = =�@�<�z�<���<Z��<�#�<�Z�<5��<���<z��<�*�<=\�<c��<0��<���<��<�?�<�h�<e��<r��<���<j��<�<=�< Z�<�t�<�<Z��<˸�<���<���<���<P��<U��<���<$�<��<w��<��<���<���<���<���<��<���<�o�<lN�<M)�<n �<���< ��<�n�<6�<���<��<Gt�<�+�<���<j��<!8�<���<���<&�<8��<	O�<��<�n�<:��<�}�<���<X}�<@��<�m�<�߱<�N�<��<�!�<M��<o�<eE�<$��<���<�L�<՞�<8�<�:�<��<�̚<q�<�U�<��<c֓<��<�O�<���<H<h��<G/�<�c�<{��<'ʃ<���<�,�<[�|<y<�xu<��q<�4n<P�j<��f<�Mc<��_<�
\<�jX<��T<�-Q<��M<�I<�^F<$�B<W4?<�;<�8<2�4<� 1<}|-<��)<�~&<�#<F�<v!<c�<oP<��<O�<�><��<Ϥ<a<�G�;���;�z�;�)�;���;��;���;~t�;�l�;cu�;���;0��;�;+8�;I��;���;lx�;��;T��;�P�;��;�;؄y;>jo;pe;ܗ[;��Q;�IH;��>;*}5;UF,;�.#;F5;1Z;��;���:���:�:���:=�:7�:I�:��:��z:n\:�v=:?:\:ѓ�9��9	7&9�N8��x�ί.�N ��Bjƹ(;�������4��O�j��9���P��zS���?��t��{�º��Ϻ�1ܺ'���C���� �k��:��`������̱%���+���1���7���=�P�C���I�\�O�~�U���[���a�i�g�7�m�p�s�֘y�݋�@��� �������l���T���4���ɠ��5���2����  �  >m==��=L=E�=/�=�(=7� =He =� =�@�<�z�< ��<g��<�#�<�Z�<9��<���<l��<�*�<D\�<\��<5��<���<��<�?�<�h�<h��<w��<���<j��<*�<=�<�Y�<�t�<���<X��<¸�<���<���<���<_��<V��<���<%�<��<h��<��<���<���<���<���<��<���<�o�<wN�<W)�<v �<���<"��<�n�<6�<���<���<Ht�<|+�<���<l��<!8�<���<��<0�<7��<O�<��<�n�<&��<�}�<���<R}�<J��<�m�<�߱<�N�<��<�!�<Q��<v�<WE�<(��<���<�L�<֞�<&�<�:�<!��<�̚<{�<�U�<��<i֓<��<�O�<���<A<g��<A/�<�c�<���<$ʃ<���<�,�<~�|< y<�xu<	�q<�4n<J�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<��M<�I<�^F<9�B<L4?<��;<�8<)�4<1<]|-<��)<�~&<�#<`�<�!<�<xP<��<4�<z><��<��<#a<�G�;���;{�;o)�;���;-��;1��;|t�;m�;]u�;���; ��;��;%8�;%��;���;wx�;��;���;�P�;��;!�;@�y;�io;�oe;��[;d�Q;�IH;H�>;"}5;qF,;�.#;�5;�Z;�;��:��:�:��:6�:��:T�:�:D�z:�\:�v=:$?:�]:.��9~�9�<&95N8��x�	�.��#���jƹ�<�������4�`�O�j��9��DQ��6S��l?��M��=�º*�Ϻ�1ܺ��E���� �M�k:�]`���������%��+�a�1��7���=�V�C���I���O��U���[���a�a�g���m�b�s���y����\������$���z���d����������5���󜚻�  �  ;m==��=L=D�=2�=�(=0� =Je =� =�@�<�z�<���<c��<�#�<�Z�<1��<���<w��<�*�<D\�<R��<A��<���<��<�?�<�h�<n��<r��<���<]��<-�<=�< Z�<�t�<���<h��<���<���<���<���<W��<W��<���<�<��<d��<��<���<���<���<���<��<���<�o�<pN�<N)�<n �<���<-��<�n�<%6�<���<���<Xt�<x+�<���<d��<#8�<���<���<(�<2��<O�<��<�n�<3��<�}�<���<M}�<O��<tm�<�߱<�N�<��<�!�<O��<y�<WE�<6��<���<�L�<ߞ�</�<�:�<��<�̚<q�<�U�<��<i֓<��<�O�<���<5<q��<I/�<�c�<���<ʃ<���<�,�<x�|<y<�xu<�q<�4n<k�j<��f<�Mc<�_<�
\<�jX<y�T<�-Q<��M<�I<�^F<<�B<G4?<�;<�8<�4<"1<k|-<��)<�~&<�#<Y�<x!<t�<hP<��<I�<�><��<��<;a<�G�;���;{�;V)�;���;��;&��;Ht�;m�;Ru�;���;A��;��;g8�;��;���;hx�;��;r��;�P�;��; �;Z�y;�io;ipe;ɗ[;"�Q;JH;d�>;�}5;XF,;�.#;g5;;Z;��;���:���:O�:���:��:��:M�:��:��z:�\:�v=:;?:�\:R��9*�91@&9�M8�lx�O�.�����iƹ�=�����O�4�؅O��j��9��wQ��SS��??��V��W�º��Ϻ�1ܺ��躍D���� ����:��`�΀�����%���+�/�1���7�B�=��C���I���O�"�U���[���a�o�g�±m�٥s���y����g���˸������5���m����������q��������  �  >m==��=L=F�=3�=�(=7� =Ce =� =�@�<�z�<��<e��<�#�<�Z�<;��<���<y��<�*�<@\�<_��</��<���<��<�?�<�h�<n��<v��<���<f��<$�<=�<�Y�<�t�<���<T��<ĸ�<���<���<���<X��<^��<���<�<��<o��<��<���<���<���<���<��<���<�o�<yN�<Z)�<t �<���<��<�n�<6�<���<���<Gt�<�+�<���<g��<!8�<���<��<-�<9��<O�<��<�n�<,��<�}�<���<X}�<D��<}m�<�߱<�N�<��<�!�<Q��<q�<`E�<$��<���<�L�<Ӟ�<4�<�:�<"��<�̚<~�<�U�<��<c֓<��<�O�<���<D<g��<D/�<�c�<���< ʃ<���<�,�<s�|<y<�xu<�q<�4n<D�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<��M<�I<�^F<1�B<P4?<�;<�8<,�4<1<q|-<��)<�~&<�#<^�<�!<y�<}P<��<M�<|><��<Ǥ<a<�G�;���;{�;V)�;���;(��;"��;mt�;�l�;tu�;���;��;��;8�;.��;���;yx�;��;t��;Q�;��;�;�y; jo;�oe;��[;~�Q;�IH;��>;"}5;oF,;�.#;�5;�Z;ޜ;��:���:��:���:c�:��:H�:Q�:��z:\:�v=:"@:]:���9��9_:&9�N8G�x��.�S"��Elƹ�:��K��;�4�؅O�Sj�u9��tQ��.S���?�����}�º�Ϻ�1ܺG��1D��� �G�u:�C`�������ʱ%���+���1�h�7���=�U�C���I��O�J�U���[���a�M�g�ױm�i�s�Řy����P���������x���h������Ġ��:�������  �  >m==��=L=D�=3�=�(=?� =Ce =� =�@�<�z�<��<Y��<�#�<}Z�<>��<���<y��<�*�<C\�<k��<*��<���<��<�?�<�h�<f��<v��<���<m��<�<=�<�Y�<�t�<���<Q��<ɸ�<���<���<���<V��<Y��<���<+�<��<s��<��<���<���<���<���<ݧ�<���<�o�<qN�<U)�<h �<���<��<�n�<6�<���<���<Ft�<�+�<���<r��<8�<���<��<(�<7��<O�<��<�n�<9��<�}�<���<[}�<;��<�m�<�߱<�N�<��<�!�<X��<j�<fE�<��<���<�L�<Ҟ�<7�<�:�<&��<�̚<�<�U�<��<j֓<��<�O�<���<R<c��<D/�<�c�<���<'ʃ<���<�,�<i�|<'y<�xu<��q<�4n<<�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<��M<��I<�^F<<�B<H4?<�;<}8<K�4<1<r|-<��)<�~&<�#<E�<�!<Y�<�P<��<O�<y><��<ޤ<a< H�;���;({�;^)�;���;'��;	��;�t�;�l�;vu�;���;��;�;8�;D��;���;ix�;��;o��;�P�;f�;5�;�y;jo;�oe;��[;��Q;�IH;��>; }5;�F,;�.#;r5;qZ;��;v��:���:?�:k��:��:��:9�:��:��z:v\:iu=:�?:�\:>��9y�95&9�N8�x�_�.�� ��olƹ:��a����4���O�>j��9���Q���R��+@��j����º}�Ϻ`1ܺ]���C��� �!��:�?`�
�������%�0�+���1�f�7�V�=�w�C���I���O�5�U���[��a�K�g���m�C�s��y���B���)���ʲ������a���0���Ӡ��!�������  �  ?m==��=L=B�=5�=�(=2� =Ee =  =�@�<�z�<���<e��<�#�<�Z�<9��<���<u��<�*�<B\�<W��<<��<���<��<�?�<�h�<n��<u��<���<a��<*�<	=�<�Y�<�t�<���<V��<���<���<���<���<U��<Z��<���<"�<��<d��<��<���<���<���<���<��<���<�o�<|N�<^)�<o �<���<$��<�n�<6�<���<���<Xt�<y+�<���<j��<8�<���<���<$�<5��<O�<��<�n�<0��<�}�<���<P}�<K��<xm�<�߱<�N�<��<�!�<T��<r�<[E�<1��<���<�L�<ڞ�</�<�:�<!��<�̚<��<�U�<��<j֓<��<�O�<���<9<n��<N/�<�c�<���<ʃ<���<�,�<i�|<
y<�xu<�q<�4n<H�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<��M<�I<�^F<A�B<>4?<�;<�8<�4<1<v|-<��)<�~&<�#<]�<�!<s�<wP<��<F�<�><��<��<1a<�G�;���;${�;X)�;���;#��;��;Zt�;m�;Vu�;���;��;��;8�;��;���;vx�;��;i��;Q�;��;�; �y;�io;�pe;ɗ[;J�Q;�IH;��>;V}5;sF,;�.#;�5;�Z;��;��:3��:��:��:�:��:_�:��:��z:r\:6v=:�?:�\:T��9�9)?&9��M8o�x���.��!���kƹ=��l����4���O��j�s9���Q���R���?������ºm�Ϻ�1ܺ��躋D���� �J��:�`���������%���+��1�8�7�$�=��C�m�I���O��U���[���a�9�g���m���s���y����o����������y���v���#�������`�������  �  :m==��=L=E�=.�=�(=4� =Ke =� =�@�<�z�<��<j��<�#�<�Z�<6��<���<s��<�*�<J\�<Y��<?��<���<��<�?�<�h�<p��<l��<���<U��<-�<=�<�Y�<�t�<���<_��<���<���<x��<���<\��<T��<���<�<��<^��<��<���<���<���<���<��<���<�o�<xN�<T)�<y �<���<,��<�n�<#6�<���<���<Qt�<o+�<���<Z��<#8�<���<��<1�<&��<O�<��<�n�<)��<�}�<���<K}�<N��<jm�<�߱<�N�<��<�!�<F��<}�<NE�<2��<���<�L�<ܞ�<+�<�:�<��<�̚<q�<�U�<��<i֓<��<�O�<���<<<q��<A/�<�c�<���<ʃ<���<�,�<��|<y<�xu<�q<�4n<X�j<��f<�Mc<�_<�
\<�jX<}�T<�-Q<z�M<�I<u^F<;�B<L4?<�;<�8<�4<&1<g|-<��)<�~&<�#<f�<v!<��<rP<��<C�<�><��<��<7a<�G�;���;�z�;S)�;��; ��;O��;*t�;m�;Mu�;���;��;��;B8�;���;���;Hx�;��;���;�P�;��;���;��y;xio;;pe;ؗ[;g�Q;JH;7�>;�}5;KF,;/#;�5;lZ;�;���:���:��:���:��:��:��:5�:��z:�\:�v=:S?:6]:���9j�9)?&9��M8�~x�i�.��!���iƹ'>������4�ʄO�[j�u9��uQ���S���>�������ºA�Ϻ-1ܺ��躾D���� �}�1:��`����q����%���+�Q�1���7��=��C���I���O� �U�:�[���a���g���m���s�˘y����c���񸅻-���a���e���%�������i���䜚��  �  8m==��=L=H�=1�=�(=9� =De =� =�@�<�z�<���<e��<�#�<�Z�<3��<���<{��<�*�<@\�<c��<9��<���<��<�?�<�h�<m��<h��<���<^��<*�<
=�<�Y�<�t�<���<U��<���<���<|��<���<R��<Q��<���< �<��<l��<
��<���<���<���<���<��<���<�o�<xN�<Y)�<s �<���<+��<�n�<6�<���<���<Lt�<~+�<���<f��<)8�<���<���<*�<.��<O�<��<�n�<6��<�}�<���<P}�<I��<tm�<�߱<�N�<��<�!�<I��<r�<]E�<,��<���<�L�<՞�<5�<�:�<��<�̚<}�<�U�<��<j֓<��<�O�<���<F<m��<D/�<�c�<���<"ʃ<���<�,�<n�|<y<�xu<��q<�4n<>�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<r�M<�I<�^F<*�B<W4?<��;<�8<4�4<
1<p|-<��)<�~&<�#<]�<�!<}�<mP<��<R�<�><��<Ф<,a<�G�;���;�z�;�)�;���;��;��;Nt�;m�;Yu�;���;��;�;8�;��;���;Zx�;��;`��;�P�;��;�;'�y;�io;"pe;�[;��Q;�IH;��>;p}5;tF,;�.#;�5;�Z;؜;%��:���:��:���:i�:�:��:%�:��z:�\:�w=:?:	\:Ӕ�9^�9�:&9��M8U�x�ֱ.�/!���lƹ=�����@�4��O��j��9���P���S���?�������ºǏϺ�1ܺ0��D���� �t�{:�K`���������%���+��1�C�7���=�#�C���I�j�O�W�U���[���a���g��m���s�Řy�ҋ�`���%���ᲈ�����w���2�������N�������  �  Dm=
=��=L=G�=4�=�(=9� =Ce = =�@�<�z�<��<d��< $�<�Z�<A��<���<s��<�*�<@\�<b��<-��<���<��<�?�<�h�<d��<���<���<d��<�<
=�<�Y�<�t�<���<I��<ĸ�<���<���<���<[��<^��<���<+�<��<r��<��<���<���<���<���<ڧ�<���<�o�<~N�<a)�<n �<���<��<�n�<6�<���<���<Gt�<�+�<��<r��<8�<���<��< �<9��<O�<��<{n�<-��<�}�<}��<T}�<>��<}m�<�߱<�N�<��<�!�<Y��<l�<eE�<"��<���<�L�<ߞ�<1�<�:�<+��<�̚<��<�U�<��<o֓<��<�O�<���<G<e��<G/�<�c�<}��<'ʃ<���<�,�<n�|<y<�xu<��q<�4n<%�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<��M<��I<�^F<.�B<S4?<�;<�8<2�4<1<�|-<��)<�~&<�#<[�<�!<p�<�P<��<C�<�><��<ͤ<a< H�;���;!{�;R)�;���;U��;��;ft�;�l�;\u�;���;�;��;�7�;/��;���;�x�;��;���;Q�;[�;7�;߄y;jo;pe;��[;��Q;�IH;��>;�|5;�F,;�.#;�5;�Z;��;���:r��:'�:ʁ�:��:��:K�:��:��z:�\:=u=:�?:�]:i��9"�9�6&9N80�x��.�$���mƹ<�����4��O�!j��9���Q���R��@��t����º܏Ϻ�1ܺ���eD��� ����:��_�������k�%�.�+���1�\�7���=�d�C���I�k�O�n�U���[�"�a��g��m�̥s���y����G���V���㲈�����[���<���ʠ��`�������  �  =m==��=L=D�=2�=�(=8� =Ge = =�@�<�z�<��<f��<�#�<�Z�<=��<���<w��<�*�<D\�<b��<9��<���<��<�?�<�h�<g��<s��<���<`��<#�<=�<�Y�<�t�<���<W��<���<���<���<���<U��<U��<���<%�<��<j��<��<���<���<���<���<��<���<�o�<uN�<U)�<p �<���<!��<�n�<6�<���<��<Pt�<{+�<���<l��<8�<���<���<#�<3��<O�<��<�n�<0��<�}�<���<M}�<B��<wm�<�߱<�N�<��<�!�<V��<p�<ZE�<,��<���<�L�<ޞ�<5�<�:�<&��<�̚<y�<�U�<��<q֓<��<�O�<���<F<n��<C/�<�c�<���<#ʃ<���<�,�<j�|<y<�xu<��q<�4n<E�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<��M<�I<�^F<;�B<H4?<��;<�8</�4<1<�|-<��)<�~&<�#<`�<�!<y�<�P<��<J�<�><��<Τ<,a<�G�;���;!{�;R)�;���;��;��;Yt�;�l�;Bu�;���;��;��;%8�;��;���;sx�;��;j��;�P�;k�;!�;�y;�io;=pe;�[;��Q;�IH;��>;3}5;�F,;�.#;�5;rZ;��;���:��:.�::��:��:6�:��: �:��z:�\:Yu=:�>:�\:+��9��98&9�M8��x���.��!���kƹ�=��u����4��O��j��9���Q���R���?������º��Ϻ�1ܺ���"D���� �'��:�l`�������]�%���+���1�'�7���=��C���I���O�&�U���[��a�^�g���m�ås���y���P����������w���a���S�������]�������  �  6m==��=L=F�=1�=�(=6� =Ge =� =�@�<�z�<��<u��<�#�<�Z�<5��<���<x��<�*�<F\�<^��<<��<���<��<�?�<�h�<p��<d��<���<Z��<.�<	=�<�Y�<�t�<���<R��<���<���<{��<���<S��<N��<���<�<��<g��<��<���<���<���<���<��<���<�o�<�N�<^)�<� �<���<-��<�n�<6�<���<���<Qt�<x+�<���<d��<(8�<���<���<2�<+��<O�<��<�n�<#��<�}�<}��<M}�<O��<om�<�߱<�N�<��<�!�<J��<x�<YE�</��<���<�L�<Ӟ�<2�<�:�<��<͚<|�<�U�<��<j֓<��<�O�<���<B<n��<B/�<�c�<���<ʃ<���<�,�<w�|<y<�xu<�q<�4n<A�j<��f<�Mc<ԫ_<�
\<�jX<��T<�-Q<l�M<�I<�^F<6�B<P4?<��;<�8<%�4<1<h|-<��)<�~&<�#<~�<�!<��<qP<��<M�<z><��<Ƥ<1a<�G�;���;�z�;x)�;��;��;I��;?t�; m�;Vu�;���;��;��;8�;���;���;Vx�;��;e��;�P�;��;���;X�y;�io;;pe;͗[;z�Q;�IH;��>;�}5;aF,;/#;�5;�Z;K�;��:���:��:���:S�:��:��:��:��z:�\:�w=:�>:�[:��9��9�?&9��M8��x�Ժ.��#���mƹ�=�������4�ׄO�\j�}9��Q���S��F?��3����º��Ϻp1ܺK��LD��|� �i��9�P`�J��n����%���+��1��7���=��C���I���O��U� �[�x�a�ƽg�űm���s���y����������,�����������(�������c�����  �  =m==��=L=F�=4�=�(=9� =Ie = =�@�<�z�<��<d��<�#�<�Z�<:��<���<{��<�*�<J\�<^��<4��<���<��<�?�<�h�<g��<p��<���<U��<!�<=�<�Y�<�t�<���<X��<���<���<s��<���<U��<U��<���<�<��<k��<��<���<���<���<���<��<���<�o�<qN�<P)�<u �<���<&��<�n�< 6�<���<���<Pt�<+�<���<g��<8�<���<���<)�<%��<O�<��<�n�<-��<�}�<���<O}�<B��<lm�<�߱<�N�<��<�!�<O��<u�<`E�<)��<���<�L�<���<5�<�:�<#��<�̚<p�<�U�<��<l֓<��<�O�<���<H<g��<J/�<�c�<���<ʃ<���<�,�<s�|<y<�xu<��q<�4n<K�j<��f<�Mc<�_<�
\<�jX<s�T<�-Q<��M<�I<}^F<8�B<N4?<�;<�8<2�4<1<�|-<��)<�~&<�#<[�<y!<�<zP<��<R�<�><��<Ƥ<"a<�G�;���;{�;N)�;���;��;1��;+t�;�l�;Tu�;���;��;��;)8�;��;���;6x�;��;j��;�P�;z�;�;B�y;�io;Ipe;��[;��Q;�IH;��>;`}5;�F,;�.#;v5;NZ;�;i��:b��:�:X��:��:��:��:6�:9�z:9\:�u=:)?:]\:���9#�9�9&9��M8.�x�.�.��!��kƹ+=�����?�4�~�O�2j��9���Q��ES��p?������º�Ϻ1ܺs��D���� �7�l:��`�΀�x����%���+���1��7���=�W�C���I���O�'�U��[���a�p�g�Աm�ڥs��y�ԋ�^���
������q���n���/���ޠ��~��������  �  >m==��=L=A�=7�=�(=8� =Ae = =�@�<�z�<��<i��<$�<�Z�<B��<���<t��<�*�<9\�<]��<6��<���<��<�?�<�h�<j��<w��<���<e��<(�<=�<�Y�<�t�<���<P��<���<���<���<���<P��<^��<���<,�<��<g��<��<���<���<���<���<ާ�<���<�o�<N�<b)�<u �<���<��<�n�<6�<���<���<Qt�<|+�<���<u��<8�<���<���<"�<7��<O�<��<�n�<#��<�}�<���<J}�<D��<}m�<�߱<�N�<��<�!�<]��<h�<`E�<+��<���<�L�<ڞ�<1�<�:�<-��<�̚<��<�U�<!��<k֓<��<�O�<���<D<d��<P/�<�c�<���<'ʃ<���<�,�<b�|<y<�xu<��q<�4n</�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<��M< �I<�^F<@�B<:4?<�;<�8<0�4<� 1<�|-<��)<�~&<�#<e�<�!<��<�P<��<D�<�><��<ä<&a<�G�;���;7{�;^)�;���;/��;���;kt�;m�;=u�;���;ᵸ;��;8�;��;���;�x�;��;W��;Q�;m�;=�;��y;�io;npe;��[;_�Q;�IH;��>;	}5;�F,;�.#;�5;�Z;�;���:���:=�:���:�:��:��:�:��z:�\:Wu=:.@:.\:��9��9�8&96�M8%�x��.�7%���lƹD>��5��(�4�;�O��j��9���Q��pR��8@����� �º"�Ϻ2ܺ���dD���� ���X:��_����c����%��+���1���7���=�l�C�_�I���O�$�U���[���a�C�g��m���s���y���l���B���-�������v���I�������@���/����  �  =m==��=L=F�=4�=�(=9� =Ie = =�@�<�z�<��<d��<�#�<�Z�<:��<���<{��<�*�<J\�<^��<4��<���<��<�?�<�h�<g��<p��<���<U��<!�<=�<�Y�<�t�<���<X��<���<���<s��<���<U��<U��<���<�<��<k��<��<���<���<���<���<��<���<�o�<qN�<P)�<u �<���<&��<�n�< 6�<���<���<Pt�<+�<���<g��<8�<���<���<)�<%��<O�<��<�n�<-��<�}�<���<O}�<B��<lm�<�߱<�N�<��<�!�<O��<u�<`E�<)��<���<�L�<���<5�<�:�<#��<�̚<p�<�U�<��<l֓<��<�O�<���<H<g��<J/�<�c�<���<ʃ<���<�,�<s�|<y<�xu<��q<�4n<K�j<��f<�Mc<�_<�
\<�jX<s�T<�-Q<��M<�I<}^F<8�B<N4?<�;<�8<2�4<1<�|-<��)<�~&<�#<[�<y!<�<zP<��<R�<�><��<Ƥ<"a<�G�;���;{�;N)�;���;��;1��;+t�;�l�;Tu�;���;��;��;)8�;��;���;6x�;��;j��;�P�;z�;�;B�y;�io;Ipe;��[;��Q;�IH;��>;`}5;�F,;�.#;v5;NZ;�;i��:b��:�:X��:��:��:��:6�:9�z:9\:�u=:)?:]\:���9#�9�9&9��M8.�x�.�.��!��kƹ+=�����?�4�~�O�2j��9���Q��ES��p?������º�Ϻ1ܺs��D���� �7�l:��`�΀�x����%���+���1��7���=�W�C���I���O�'�U��[���a�p�g�Աm�ڥs��y�ԋ�^���
������q���n���/���ޠ��~��������  �  6m==��=L=F�=1�=�(=6� =Ge =� =�@�<�z�<��<u��<�#�<�Z�<5��<���<x��<�*�<F\�<^��<<��<���<��<�?�<�h�<p��<d��<���<Z��<.�<	=�<�Y�<�t�<���<R��<���<���<{��<���<S��<N��<���<�<��<g��<��<���<���<���<���<��<���<�o�<�N�<^)�<� �<���<-��<�n�<6�<���<���<Qt�<x+�<���<d��<(8�<���<���<2�<+��<O�<��<�n�<#��<�}�<}��<M}�<O��<om�<�߱<�N�<��<�!�<J��<x�<YE�</��<���<�L�<Ӟ�<2�<�:�<��<͚<|�<�U�<��<j֓<��<�O�<���<B<n��<B/�<�c�<���<ʃ<���<�,�<w�|<y<�xu<�q<�4n<A�j<��f<�Mc<ԫ_<�
\<�jX<��T<�-Q<l�M<�I<�^F<6�B<P4?<��;<�8<%�4<1<h|-<��)<�~&<�#<~�<�!<��<qP<��<M�<z><��<Ƥ<1a<�G�;���;�z�;x)�;��;��;I��;?t�; m�;Vu�;���;��;��;8�;���;���;Vx�;��;e��;�P�;��;���;X�y;�io;;pe;͗[;z�Q;�IH;��>;�}5;aF,;/#;�5;�Z;K�;��:���:��:���:S�:��:��:��:��z:�\:�w=:�>:�[:��9��9�?&9��M8��x�Ժ.��#���mƹ�=�������4�ׄO�\j�}9��Q���S��F?��3����º��Ϻp1ܺK��LD��|� �i��9�P`�J��n����%���+��1��7���=��C���I���O��U� �[�x�a�ƽg�űm���s���y����������,�����������(�������c�����  �  =m==��=L=D�=2�=�(=8� =Ge = =�@�<�z�<��<f��<�#�<�Z�<=��<���<w��<�*�<D\�<b��<9��<���<��<�?�<�h�<g��<s��<���<`��<#�<=�<�Y�<�t�<���<W��<���<���<���<���<U��<U��<���<%�<��<j��<��<���<���<���<���<��<���<�o�<uN�<U)�<p �<���<!��<�n�<6�<���<��<Pt�<{+�<���<l��<8�<���<���<#�<3��<O�<��<�n�<0��<�}�<���<M}�<B��<wm�<�߱<�N�<��<�!�<V��<p�<ZE�<,��<���<�L�<ޞ�<5�<�:�<&��<�̚<y�<�U�<��<q֓<��<�O�<���<F<n��<C/�<�c�<���<#ʃ<���<�,�<j�|<y<�xu<��q<�4n<E�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<��M<�I<�^F<;�B<H4?<��;<�8</�4<1<�|-<��)<�~&<�#<`�<�!<y�<�P<��<J�<�><��<Τ<,a<�G�;���;!{�;R)�;���;��;��;Yt�;�l�;Bu�;���;��;��;%8�;��;���;sx�;��;j��;�P�;k�;!�;�y;�io;=pe;�[;��Q;�IH;��>;3}5;�F,;�.#;�5;rZ;��;���:��:.�::��:��:6�:��: �:��z:�\:Yu=:�>:�\:+��9��98&9�M8��x���.��!���kƹ�=��u����4��O��j��9���Q���R���?������º��Ϻ�1ܺ���"D���� �'��:�l`�������]�%���+���1�'�7���=��C���I���O�&�U���[��a�^�g���m�ås���y���P����������w���a���S�������]�������  �  Dm=
=��=L=G�=4�=�(=9� =Ce = =�@�<�z�<��<d��< $�<�Z�<A��<���<s��<�*�<@\�<b��<-��<���<��<�?�<�h�<d��<���<���<d��<�<
=�<�Y�<�t�<���<I��<ĸ�<���<���<���<[��<^��<���<+�<��<r��<��<���<���<���<���<ڧ�<���<�o�<~N�<a)�<n �<���<��<�n�<6�<���<���<Gt�<�+�<��<r��<8�<���<��< �<9��<O�<��<{n�<-��<�}�<}��<T}�<>��<}m�<�߱<�N�<��<�!�<Y��<l�<eE�<"��<���<�L�<ߞ�<1�<�:�<+��<�̚<��<�U�<��<o֓<��<�O�<���<G<e��<G/�<�c�<}��<'ʃ<���<�,�<n�|<y<�xu<��q<�4n<%�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<��M<��I<�^F<.�B<S4?<�;<�8<2�4<1<�|-<��)<�~&<�#<[�<�!<p�<�P<��<C�<�><��<ͤ<a< H�;���;!{�;R)�;���;U��;��;ft�;�l�;\u�;���;�;��;�7�;/��;���;�x�;��;���;Q�;[�;7�;߄y;jo;pe;��[;��Q;�IH;��>;�|5;�F,;�.#;�5;�Z;��;���:r��:'�:ʁ�:��:��:K�:��:��z:�\:=u=:�?:�]:i��9"�9�6&9N80�x��.�$���mƹ<�����4��O�!j��9���Q���R��@��t����º܏Ϻ�1ܺ���eD��� ����:��_�������k�%�.�+���1�\�7���=�d�C���I�k�O�n�U���[�"�a��g��m�̥s���y����G���V���㲈�����[���<���ʠ��`�������  �  8m==��=L=H�=1�=�(=9� =De =� =�@�<�z�<���<e��<�#�<�Z�<3��<���<{��<�*�<@\�<c��<9��<���<��<�?�<�h�<m��<h��<���<^��<*�<
=�<�Y�<�t�<���<U��<���<���<|��<���<R��<Q��<���< �<��<l��<
��<���<���<���<���<��<���<�o�<xN�<Y)�<s �<���<+��<�n�<6�<���<���<Lt�<~+�<���<f��<)8�<���<���<*�<.��<O�<��<�n�<6��<�}�<���<P}�<I��<tm�<�߱<�N�<��<�!�<I��<r�<]E�<,��<���<�L�<՞�<5�<�:�<��<�̚<}�<�U�<��<j֓<��<�O�<���<F<m��<D/�<�c�<���<"ʃ<���<�,�<n�|<y<�xu<��q<�4n<>�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<r�M<�I<�^F<*�B<W4?<��;<�8<4�4<
1<p|-<��)<�~&<�#<]�<�!<}�<mP<��<R�<�><��<Ф<,a<�G�;���;�z�;�)�;���;��;��;Nt�;m�;Yu�;���;��;�;8�;��;���;Zx�;��;`��;�P�;��;�;'�y;�io;"pe;�[;��Q;�IH;��>;p}5;tF,;�.#;�5;�Z;؜;%��:���:��:���:i�:�:��:%�:��z:�\:�w=:?:	\:Ӕ�9^�9�:&9��M8U�x�ֱ.�/!���lƹ=�����@�4��O��j��9���P���S���?�������ºǏϺ�1ܺ0��D���� �t�{:�K`���������%���+��1�C�7���=�#�C���I�j�O�W�U���[���a���g��m���s�Řy�ҋ�`���%���ᲈ�����w���2�������N�������  �  :m==��=L=E�=.�=�(=4� =Ke =� =�@�<�z�<��<j��<�#�<�Z�<6��<���<s��<�*�<J\�<Y��<?��<���<��<�?�<�h�<p��<l��<���<U��<-�<=�<�Y�<�t�<���<_��<���<���<x��<���<\��<T��<���<�<��<^��<��<���<���<���<���<��<���<�o�<xN�<T)�<y �<���<,��<�n�<#6�<���<���<Qt�<o+�<���<Z��<#8�<���<��<1�<&��<O�<��<�n�<)��<�}�<���<K}�<N��<jm�<�߱<�N�<��<�!�<F��<}�<NE�<2��<���<�L�<ܞ�<+�<�:�<��<�̚<q�<�U�<��<i֓<��<�O�<���<<<q��<A/�<�c�<���<ʃ<���<�,�<��|<y<�xu<�q<�4n<X�j<��f<�Mc<�_<�
\<�jX<}�T<�-Q<z�M<�I<u^F<;�B<L4?<�;<�8<�4<&1<g|-<��)<�~&<�#<f�<v!<��<rP<��<C�<�><��<��<7a<�G�;���;�z�;S)�;��; ��;O��;*t�;m�;Mu�;���;��;��;B8�;���;���;Hx�;��;���;�P�;��;���;��y;xio;;pe;ؗ[;g�Q;JH;7�>;�}5;KF,;/#;�5;lZ;�;���:���:��:���:��:��:��:5�:��z:�\:�v=:S?:6]:���9j�9)?&9��M8�~x�i�.��!���iƹ'>������4�ʄO�[j�u9��uQ���S���>�������ºA�Ϻ-1ܺ��躾D���� �}�1:��`����q����%���+�Q�1���7��=��C���I���O� �U�:�[���a���g���m���s�˘y����c���񸅻-���a���e���%�������i���䜚��  �  ?m==��=L=B�=5�=�(=2� =Ee =  =�@�<�z�<���<e��<�#�<�Z�<9��<���<u��<�*�<B\�<W��<<��<���<��<�?�<�h�<n��<u��<���<a��<*�<	=�<�Y�<�t�<���<V��<���<���<���<���<U��<Z��<���<"�<��<d��<��<���<���<���<���<��<���<�o�<|N�<^)�<o �<���<$��<�n�<6�<���<���<Xt�<y+�<���<j��<8�<���<���<$�<5��<O�<��<�n�<0��<�}�<���<P}�<K��<xm�<�߱<�N�<��<�!�<T��<r�<[E�<1��<���<�L�<ڞ�</�<�:�<!��<�̚<��<�U�<��<j֓<��<�O�<���<9<n��<N/�<�c�<���<ʃ<���<�,�<i�|<
y<�xu<�q<�4n<H�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<��M<�I<�^F<A�B<>4?<�;<�8<�4<1<v|-<��)<�~&<�#<]�<�!<s�<wP<��<F�<�><��<��<1a<�G�;���;${�;X)�;���;#��;��;Zt�;m�;Vu�;���;��;��;8�;��;���;vx�;��;i��;Q�;��;�; �y;�io;�pe;ɗ[;J�Q;�IH;��>;V}5;sF,;�.#;�5;�Z;��;��:3��:��:��:�:��:_�:��:��z:r\:6v=:�?:�\:T��9�9)?&9��M8o�x���.��!���kƹ=��l����4���O��j�s9���Q���R���?������ºm�Ϻ�1ܺ��躋D���� �J��:�`���������%���+��1�8�7�$�=��C�m�I���O��U���[���a�9�g���m���s���y����o����������y���v���#�������`�������  �  >m==��=L=D�=3�=�(=?� =Ce =� =�@�<�z�<��<Y��<�#�<}Z�<>��<���<y��<�*�<C\�<k��<*��<���<��<�?�<�h�<f��<v��<���<m��<�<=�<�Y�<�t�<���<Q��<ɸ�<���<���<���<V��<Y��<���<+�<��<s��<��<���<���<���<���<ݧ�<���<�o�<qN�<U)�<h �<���<��<�n�<6�<���<���<Ft�<�+�<���<r��<8�<���<��<(�<7��<O�<��<�n�<9��<�}�<���<[}�<;��<�m�<�߱<�N�<��<�!�<X��<j�<fE�<��<���<�L�<Ҟ�<7�<�:�<&��<�̚<�<�U�<��<j֓<��<�O�<���<R<c��<D/�<�c�<���<'ʃ<���<�,�<i�|<'y<�xu<��q<�4n<<�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<��M<��I<�^F<<�B<H4?<�;<}8<K�4<1<r|-<��)<�~&<�#<E�<�!<Y�<�P<��<O�<y><��<ޤ<a< H�;���;({�;^)�;���;'��;	��;�t�;�l�;vu�;���;��;�;8�;D��;���;ix�;��;o��;�P�;f�;5�;�y;jo;�oe;��[;��Q;�IH;��>; }5;�F,;�.#;r5;qZ;��;v��:���:?�:k��:��:��:9�:��:��z:v\:iu=:�?:�\:>��9y�95&9�N8�x�_�.�� ��olƹ:��a����4���O�>j��9���Q���R��+@��j����º}�Ϻ`1ܺ]���C��� �!��:�?`�
�������%�0�+���1�f�7�V�=�w�C���I���O�5�U���[��a�K�g���m�C�s��y���B���)���ʲ������a���0���Ӡ��!�������  �  >m==��=L=F�=3�=�(=7� =Ce =� =�@�<�z�<��<e��<�#�<�Z�<;��<���<y��<�*�<@\�<_��</��<���<��<�?�<�h�<n��<v��<���<f��<$�<=�<�Y�<�t�<���<T��<ĸ�<���<���<���<X��<^��<���<�<��<o��<��<���<���<���<���<��<���<�o�<yN�<Z)�<t �<���<��<�n�<6�<���<���<Gt�<�+�<���<g��<!8�<���<��<-�<9��<O�<��<�n�<,��<�}�<���<X}�<D��<}m�<�߱<�N�<��<�!�<Q��<q�<`E�<$��<���<�L�<Ӟ�<4�<�:�<"��<�̚<~�<�U�<��<c֓<��<�O�<���<D<g��<D/�<�c�<���< ʃ<���<�,�<s�|<y<�xu<�q<�4n<D�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<��M<�I<�^F<1�B<P4?<�;<�8<,�4<1<q|-<��)<�~&<�#<^�<�!<y�<}P<��<M�<|><��<Ǥ<a<�G�;���;{�;V)�;���;(��;"��;mt�;�l�;tu�;���;��;��;8�;.��;���;yx�;��;t��;Q�;��;�;�y; jo;�oe;��[;~�Q;�IH;��>;"}5;oF,;�.#;�5;�Z;ޜ;��:���:��:���:c�:��:H�:Q�:��z:\:�v=:"@:]:���9��9_:&9�N8G�x��.�S"��Elƹ�:��K��;�4�؅O�Sj�u9��tQ��.S���?�����}�º�Ϻ�1ܺG��1D��� �G�u:�C`�������ʱ%���+���1�h�7���=�U�C���I��O�J�U���[���a�M�g�ױm�i�s�Řy����P���������x���h������Ġ��:�������  �  ;m==��=L=D�=2�=�(=0� =Je =� =�@�<�z�<���<c��<�#�<�Z�<1��<���<w��<�*�<D\�<R��<A��<���<��<�?�<�h�<n��<r��<���<]��<-�<=�< Z�<�t�<���<h��<���<���<���<���<W��<W��<���<�<��<d��<��<���<���<���<���<��<���<�o�<pN�<N)�<n �<���<-��<�n�<%6�<���<���<Xt�<x+�<���<d��<#8�<���<���<(�<2��<O�<��<�n�<3��<�}�<���<M}�<O��<tm�<�߱<�N�<��<�!�<O��<y�<WE�<6��<���<�L�<ߞ�</�<�:�<��<�̚<q�<�U�<��<i֓<��<�O�<���<5<q��<I/�<�c�<���<ʃ<���<�,�<x�|<y<�xu<�q<�4n<k�j<��f<�Mc<�_<�
\<�jX<y�T<�-Q<��M<�I<�^F<<�B<G4?<�;<�8<�4<"1<k|-<��)<�~&<�#<Y�<x!<t�<hP<��<I�<�><��<��<;a<�G�;���;{�;V)�;���;��;&��;Ht�;m�;Ru�;���;A��;��;g8�;��;���;hx�;��;r��;�P�;��; �;Z�y;�io;ipe;ɗ[;"�Q;JH;d�>;�}5;XF,;�.#;g5;;Z;��;���:���:O�:���:��:��:M�:��:��z:�\:�v=:;?:�\:R��9*�91@&9�M8�lx�O�.�����iƹ�=�����O�4�؅O��j��9��wQ��SS��??��V��W�º��Ϻ�1ܺ��躍D���� ����:��`�΀�����%���+�/�1���7�B�=��C���I���O�"�U���[���a�o�g�±m�٥s���y����g���˸������5���m����������q��������  �  >m==��=L=E�=/�=�(=7� =He =� =�@�<�z�< ��<g��<�#�<�Z�<9��<���<l��<�*�<D\�<\��<5��<���<��<�?�<�h�<h��<w��<���<j��<*�<=�<�Y�<�t�<���<X��<¸�<���<���<���<_��<V��<���<%�<��<h��<��<���<���<���<���<��<���<�o�<wN�<W)�<v �<���<"��<�n�<6�<���<���<Ht�<|+�<���<l��<!8�<���<��<0�<7��<O�<��<�n�<&��<�}�<���<R}�<J��<�m�<�߱<�N�<��<�!�<Q��<v�<WE�<(��<���<�L�<֞�<&�<�:�<!��<�̚<{�<�U�<��<i֓<��<�O�<���<A<g��<A/�<�c�<���<$ʃ<���<�,�<~�|< y<�xu<	�q<�4n<J�j<��f<�Mc<�_<�
\<�jX<��T<�-Q<��M<�I<�^F<9�B<L4?<��;<�8<)�4<1<]|-<��)<�~&<�#<`�<�!<�<xP<��<4�<z><��<��<#a<�G�;���;{�;o)�;���;-��;1��;|t�;m�;]u�;���; ��;��;%8�;%��;���;wx�;��;���;�P�;��;!�;@�y;�io;�oe;��[;d�Q;�IH;H�>;"}5;qF,;�.#;�5;�Z;�;��:��:�:��:6�:��:T�:�:D�z:�\:�v=:$?:�]:.��9~�9�<&95N8��x�	�.��#���jƹ�<�������4�`�O�j��9��DQ��6S��l?��M��=�º*�Ϻ�1ܺ��E���� �M�k:�]`���������%��+�a�1��7���=�V�C���I���O��U���[���a�a�g���m�b�s���y����\������$���z���d����������5���󜚻�  �  qn=j=I�=�M=M�=w�=W+=�� ==h =? =�G�<8��< ��<���<-�<'d�<p��<���<��<�6�<�h�<���<��<T��<$�<�O�<oy�<ȡ�<���<���<�<~2�<5R�<�o�<���<S��<���<	��<���<q��<g�<��<��<��<L!�<�!�<A�<��<��<�<���<m��<j��<��<ɖ�<
v�<�Q�<2)�<��<���<��<�`�<�$�<\��<��<`W�<~
�<���<>d�<�
�<��<�J�<���<bz�<��<%��<i"�<���<�(�<֥�<�<���<5�<ht�<�ޮ<�E�<,��<L	�<Hf�<�<��<�j�<n��<�	�<4U�<I��<��<N)�<^k�<u��<��<�%�<M`�<��<rЌ<T�<�:�<^n�<���<҃<��<i2�<��|<�y<1|u<��q</3n<��j<8�f<ZDc<C�_<��[<�YX<K�T<�Q<yM<=�I<PAF<c�B<�?<=~;<>�7<r_4<��0<�M-<v�)<K&<��"<	Y<�<ny<7<�<�P<��
<��<�Z<�<���;�:�;V��;?��;h;�;��;��;���;���;ݼ�;�ҽ;Y��;�0�;	x�;Ѧ;>:�;p��;A�;uސ;;��;�L�;��;!�w;#�m;$�c;�Z;ndP;	�F;(_=;�4;��*;��!;/�;��;�F;dX�:�[�:���:��:ݯ�:`��:���:�Պ:ȃv:��W:�K9:#4:���9��9$��9�9+Y8�H��W�;��q��4�̹ ��@���7��+R��l�r���}���s��3U��!����ú��к�ݺʡ����4A��n�������b�����i�%�i,��2��8��>�zD��J��
P�V�y�[���a���g�"�m��s���y�_���ł�轅�ϵ��Ю��ç�����؜������핚��  �  `n=e=F�=�M=R�=y�=^+=�� =Bh =; =�G�<=��< ��<���<-�</d�<n��<���<��<�6�<�h�<���<%��<O��<"$�<�O�<my�<���<���<���< �<�2�<8R�<�o�<���<I��<���<���<���<j��<t�<��<��<��<H!�<�!�<C�<��<
�<!�<���<g��<p��<��<і�<v�<�Q�<<)�<��<���<��<�`�<�$�<g��<���<[W�<�
�<���<8d�<�
�<��<K�<���<jz�<��<"��<_"�<~��<�(�<ե�<�<���<E�<Tt�<�ޮ<�E�<+��<W	�<@f�<��<��<�j�<r��<�	�<9U�<G��<��<C)�<bk�<x��<��<�%�<F`�<"��<sЌ<a�<�:�<fn�<���<҃<��<E2�<��|<�y<*|u<��q<3n<��j<$�f<VDc<-�_<��[<�YX<N�T<�Q<;yM<(�I<CAF<k�B<?<C~;<Z�7<q_4<��0<�M-<��)<K&<��"<Y<��<~y<2<!�<�P<��
<��<�Z<
<���;�:�;Z��;4��;6;�;h�;^��;���;ʶ�;��;�ҽ;M��;x0�;x�;�Ц;j:�;T��;EA�;�ސ;���;�L�;��;~�w;/�m;��c;�Z;�dP;|�F;�^=;4;��*;!�!;B�;��;�F;PX�:(\�:T��:n	�:%��:��:Ǘ�:�Պ:&�v:�W:*K9:1:���9��9֣�91�9dD8�K��a�;�xr���̹B�����S�7��)R���l�
s��~���s���T���!��n�ú��к�ݺ������
A��n�8��Z��@�����D�%�2,�-2�38��>�D��J��
P��V���[�A�a�
�g���m�¼s���y�"���ł�轅�����ڮ��������圔����������  �  ^n=t=F�=�M=P�=r�=^+=�� =Fh =7 =�G�<9��<���<���<�,�<5d�<g��<���<��<�6�<�h�<���<&��<<��<"$�<|O�<uy�<ա�<���<���<��<�2�<4R�<�o�<���<H��<���<���<���<^��<p�<��<��<��<C!�<�!�<3�<��<�<�<���<^��<q��<��<ϖ�<v�<�Q�<>)�<	��<���<���<�`�<�$�<`��<���<JW�<�
�<{��<Ld�<�
�< ��<K�<���<uz�<��<+��<^"�<���<�(�<Х�<�<���<L�<Lt�<�ޮ<�E�<%��<Y	�<,f�<
��<��<�j�<s��<�	�<7U�<?��<��<7)�<fk�<s��<��<�%�<<`�<)��<iЌ<a�<�:�<^n�<���<҃<��<C2�<��|<�y<#|u<��q<�2n<�j<$�f<pDc<�_<��[<�YX<8�T<Q<1yM<b�I<EAF<j�B<?<'~;<[�7<`_4<��0<�M-<�)<K&<��"<Y<��<�y<%<�<�P<��
<��<�Z<<_��;�:�;H��;U��;�;�;A�;���;���;߶�;ۼ�;�ҽ;l��;s0�;3x�;�Ц;�:�;$��;3A�;�ސ;֌�;�L�;��;��w;��m;y�c;�Z;WdP;��F;�^=; 4;��*;�!;;�;��;�F;�W�:1\�:���:�	�:ϯ�:���:���:jԊ:��v:�W:�M9:v2:���9��9V��9��9N28�B����;��q����̹Տ����܁7��(R���l��q��M}��?t��cT���"��M�ú�к�ݺ���]��A�o�����������l�%�3,��2��8�!>�D�J��
P��V���[�l�a��g���m��s�ìy����ł����������������ꡑ�㜔�Ę�������  �  cn=j=>�=�M=S�=x�=^+=�� =Bh =9 =�G�<?��<��<���<-�<4d�<t��<���<��<�6�<�h�<���<��<P��<"$�<~O�<^y�<ǡ�<���<���<��<�2�</R�<�o�<���<A��<���<���<���<f��<n�<��<��<��<?!�<�!�<B�<��<
�<#�<���<i��<l��<��<і�<v�<�Q�<=)�<��<���<��<�`�<�$�<e��<���<]W�<�
�<x��<3d�<�
�<���<�J�<���<lz�<��<'��<\"�<���<�(�<ͥ�<�<���<C�<Ot�<�ޮ<�E�<$��<Y	�<Af�<��<��<�j�<p��<�	�<:U�<L��<��<A)�<fk�<z��<��<�%�<D`�<��<pЌ<b�<�:�<gn�<���<҃<��<O2�<��|<�y<5|u<��q<�2n<�j<�f<hDc<�_<��[<�YX<=�T<�Q<EyM<;�I<#AF<r�B<?<=~;<Y�7<j_4<��0<�M-<z�)<K&<��"<Y<��<�y<><!�<�P<��
<��<�Z<�<���;�:�;O��;���;d;�;b�;[��;���;��;ļ�;�ҽ;i��;U0�;x�;�Ц;t:�;E��;,A�;mސ;茋;�L�;w�;��w;*�m;��c;�Z;�dP;X�F;_=;�4;��*;"�!;B�;��;�F;�X�:\�:_��:	�:b��:ꊪ:���:�Պ:օv:��W:�J9:12:���9q�9_��9C�9�18&F����;��q����̹M����ހ7��)R�1�l�er���~��Jt��`T��~!����ú׃кDݺ�����A��n���i����}��%�%�S,�C2�K8��>�D��J��
P��V��[��a���g���m��s�{�y�#���ł�Ƚ���������������Ĝ�����������  �  dn=g=I�=�M=L�=x�=X+=�� =@h =? =�G�<A��<��<���<-�<)d�<r��<���<��<�6�<�h�<���<��<S��<$�<�O�<ry�<ġ�<���<���<��<2�<7R�<�o�<���<E��<���<��<���<k��<u�<��<��<��<Y!�<�!�<=�<��<��<$�<���<u��<e��<��<Ӗ�<v�<�Q�<<)�<��<���<���<�`�<�$�<^��<��<ZW�<�
�<���<:d�<�
�<���<K�<���<iz�<��<$��<Z"�<~��<�(�<֥�<�<���<C�<Tt�<�ޮ<�E�<<��<H	�<Cf�<���<��<�j�<p��<�	�<3U�<J��<��<C)�<^k�<y��<��<�%�<Q`�<��<wЌ<V�<�:�<\n�<���<҃<��<P2�<��|<�y<,|u<��q<3n<
�j<�f<aDc<0�_<��[<�YX<G�T<�Q<JyM<.�I<RAF<{�B<�?<@~;<A�7<x_4<��0<�M-<��)<!K&<��"<Y<��<ry<:<�<�P<��
<��<�Z<�<���;x:�;���;I��;V;�;q�;J��;���;Ķ�;��;�ҽ;Y��;f0�;x�;�Ц;o:�;Y��;FA�;fސ;茋;�L�;��;T�w;�m;a�c;�Z;�dP;4�F;e_=;�4;�*;-�!;9�;��;�F;�X�:�[�:��:��:Y��:���:3��:fՊ:�v:$�W:wK9:;2:m��9��9Z��9��9 O8kI����;�nr����̹�����7��)R���l�~r���}���r��nU��`!���ú��к�ݺ���o��9A��n�^��[��^������%�F,��2�m8��>�mD��J�P��V�=�[�@�a���g��m�߼s���y�!���ł�ѽ�����î��駎�������������ϕ���  �  an=n=D�=�M=N�=|�=\+=�� =Bh =; =�G�<;��<��<���<-�<9d�<s��<���<��<�6�<�h�<���<#��<S��<$�<|O�<jy�<͡�<���<���<��<~2�<2R�<�o�<���<B��<���<���<���<]��<q�<��<��<��<E!�<�!�<?�<��<�<!�<���<m��<o��<��<ז�<v�<�Q�<D)�<��<���<��<�`�<�$�<^��<���<ZW�<�
�<~��<@d�<�
�<���<K�<���<jz�<��<'��<W"�<y��<�(�<ϥ�<�<���<H�<Lt�<�ޮ<�E�<%��<N	�<Bf�<
��<��<�j�<u��<�	�<6U�<I��<��<@)�<hk�<y��<��<�%�<H`�<!��<uЌ<\�<;�<`n�<���<҃<��<K2�<��|<�y<|u<��q<3n<	�j<�f<`Dc<�_<��[<�YX<C�T<�Q<>yM<I�I<>AF<]�B< ?<P~;<Q�7<w_4<��0<�M-<��)<K&<��"<"Y<��<�y<=<�<�P<��
<��<�Z<<���;�:�;H��;+��;|;�;W�;j��;���;���;Ӽ�;�ҽ;H��;]0�; x�;�Ц;s:�;��;8A�;Zސ;�;�L�;��;J�w;�m;��c;�Z;�dP;w�F;$_=;4;��*;R�!;A�;��;G;}X�:\�:���:a	�:��:���:��:qՊ:b�v:w�W:JL9:�2:���9��9⠅9U�9�58�F����;��s����̹���ʤ�N�7�&)R���l�
r���}��5t��U��o!��I�ú��к�ݺb����� A��n���m�������W�%�3,�#2�78��>�@D�xJ��
P��V���[���a���g���m��s�ݬy����ł�ӽ�����Ů����������������������  �  \n=l=A�=�M=R�=u�=\+=�� =Gh =; =�G�<>��<��<���<�,�<;d�<l��<���<��<�6�<�h�<���< ��<D��<,$�<�O�<dy�<š�<���<���<��<�2�<(R�<�o�<���<8��<���<���<���<]��<x�<��<��<��<=!�<�!�<8�<��<�<�< ��<f��<u��<��<ۖ�<v�<�Q�<H)�<��<��<��<�`�<�$�<_��<��<PW�<�
�<w��<:d�<�
�<���<	K�<���<pz�<��<-��<Q"�<y��<�(�<ť�<�<���<N�<Ht�<�ޮ<�E�<&��<e	�<4f�<��<��<�j�<}��<�	�<?U�<C��<��<9)�<jk�<{��<��<�%�<E`�<+��<mЌ<\�<�:�<bn�<���<҃<��<@2�<��|<�y<|u<��q<�2n<�j<�f<hDc<�_<��[<�YX<;�T<Q<*yM<A�I</AF<}�B<?<2~;<S�7<f_4<��0<�M-<��)<K&<��"<&Y<��<�y<0<,�<�P<��
<��<�Z<<���;�:�;`��;��;\;�;>�;���;���;ݶ�;���;�ҽ;S��;40�;<x�;�Ц;�:�;��;SA�;fސ;Ɍ�;�L�;r�; x;��m;�c;�Z;gdP;��F;�^=;C4;��*;m�!;:�;��;3G;X�:�\�:.��:�	�:寺:���:���:�Ԋ:��v:��W:|K9:�1:���9-�92��9��9g&8�?���;��s��V�̹5��ģ�
�7�R(R��l�zr��N~��!t���S��B"����ú$�к�ݺ��.���@��n�ȕ������r��F�%�!,�62��8�>�AD�J��
P�QV���[���a�4�g���m���s�Ԭy�.���ł�����=�������������휔����������  �  `n=k=H�=�M=L�=x�=_+=�� =Dh => =�G�<E��<��<���<-�<6d�<p��<���<��<�6�<�h�<���<#��<M��<$�<�O�<uy�<š�<���<���<��<�2�<'R�<�o�<���<>��<���<���<���<c��<o�<��<��<��<J!�<�!�<9�<��<
�<�<���<l��<m��<��<Ԗ�<v�<�Q�<A)�<��<���<��<�`�<�$�<h��<���<VW�<�
�<���<Ad�<�
�<���<K�<���<hz�<��<)��<T"�<x��<�(�<ƥ�<�<���<D�<Mt�<�ޮ<�E�<+��<L	�<=f�<��<��<�j�<w��<�	�<=U�<G��<��<E)�<fk�<{��<��<�%�<J`�<$��<uЌ<c�<�:�<Zn�<���<҃<��<I2�<��|<�y<%|u<��q<3n<�j<�f<cDc< �_<{�[<�YX<9�T<�Q<:yM<A�I<MAF<h�B<�?<?~;<]�7<y_4<��0<�M-<z�)<)K&<��"<Y<��<�y<7<,�<�P<��
<��<�Z<<���;�:�;b��;Y��;[;�;Z�;a��;���;Ͷ�;���;�ҽ;M��;M0�;)x�;�Ц;]:�;;��;3A�;Xސ;ڌ�;�L�;��;W�w;��m;��c;Z;�dP;��F;#_=;4;�*;=�!;H�;��;�F;�X�:!\�:}��:�	�:��: ��:嗚:,Պ:r�v:�W:fL9:�1:���9�9�9��948�C��t�;��s��?�̹�����[�7��)R�f�l��r���}���s��*U���!��\�úq�к�ݺ<��<���@��n����G����u����%�T,�2�"8��>�D��J�P��V�v�[���a���g���m��s���y�b���ł�ǽ������������$���朔�Ø�������  �  `n=g=E�=�M=T�=|�=X+=�� =?h =? =�G�<G��<��<���<-�<6d�<}��<���<��<�6�<�h�<���<��<\��<$�<O�<hy�<���<���<���<��<}2�<2R�<�o�<���<@��<���<���<���<i��<i�<��<��<��<K!�<�!�<O�<��<�<(�<���<x��<l��<���<Ӗ�<v�<�Q�<>)�<!��<���<���<�`�<�$�<b��<���<kW�<~
�<���<4d�<�
�<���<�J�<���<`z�<��<��<V"�<v��<�(�<ϥ�<�<���<<�<Pt�<�ޮ<�E�<)��<P	�<Of�<���<��<�j�<{��<�	�<<U�<V��<��<G)�<jk�<~��<��<�%�<P`�<��<|Ќ<X�< ;�<nn�<���<҃<��<H2�<��|<�y</|u<��q<3n<�j<�f<BDc<�_<��[<�YX<C�T<�Q<;yM<.�I<AAF<\�B<?<Q~;<C�7<�_4<��0<�M-<��)<-K&<��"<!Y<��<�y<R<+�<�P<��
<��<�Z<�<��;�:�;W��;#��;K;�;f�;E��;���;���;Լ�;�ҽ;5��;W0�;�w�;�Ц;J:�;R��;A�;fސ;݌�;�L�;��;,�w;��m;��c;�Z;�dP;{�F;}_=;�4;N�*;6�!;k�;��;�F;VY�:
\�:G��:�	�:���:ʊ�:���:�֊:�v:��W:�J9:�1:��9E�9���9��9�;8�M��o�;�It����̹ۏ����C�7��*R��l��r��a~���s���T��� ���ú~�к�ݺ���m���@�Cn���9�����\����%�:,��2�c8��>�[D��J�s
P�V�{�[�7�a���g�	�m��s���y�`���ł�	������ ���������ܜ������ϕ���  �  ]n=m=E�=�M=P�=r�=[+=�� =Bh == =�G�<C��<��<���<-�<8d�<n��<���<��<�6�<�h�<���<��<B��< $�<�O�<gy�<̡�<���<���<��<}2�<.R�<�o�<���<>��<���<���<���<_��<j�<��<��<��<J!�<�!�<6�<��<�<#�<���<o��<q��<��<Ֆ�<v�<�Q�<B)�<��<���<��<�`�<�$�<b��<��<PW�<�
�<���<;d�<�
�<���<�J�<���<hz�<��<#��<T"�<x��<�(�<˥�<�<���<@�<Mt�<�ޮ<�E�<.��<W	�<5f�<���<��<�j�<t��<�	�<=U�<F��<��<A)�<nk�<v��<��<�%�<L`�<!��<xЌ<^�<�:�<^n�<���<҃<��<C2�<��|<�y<|u<��q<3n<�j<�f<YDc<"�_<��[<�YX<2�T<�Q</yM<G�I<?AF<y�B<?<&~;<P�7<�_4<��0<�M-<��)<%K&<��"<(Y<��<�y<4<+�<�P<��
<��<�Z<�<{��;�:�;z��;#��;x;�;M�;U��;���;���;ļ�;�ҽ;M��;O0�;x�;�Ц;j:�;+��;A�;|ސ;݌�;�L�;��;��w;��m;=�c;�Z;�dP;r�F;;_=;*4;��*;B�!;��;��;G;�X�:H\�:ė�:>	�:8��:���:��:�Ԋ:хv:N�W:�K9:O2:u��9��9䠅9��978-I��k�;��s���̹k�� ����7�*R�n�l�r��.~���s���T��;"��	�ú��кݺj�麔���@��n����h���������%��,��2�88��>�0D�'J��
P��V���[���a��g���m�*�s�׬y�P���ł�ܽ�����Ү������������И�������  �  [n=n=>�=�M=N�=z�=d+=�� =Hh =; =�G�<I��<��<���<-�<?d�<n��<���<��<�6�<�h�<���<0��<M��<$�<~O�<by�<ʡ�<~��<���<��<�2�<#R�<�o�<���<6��<���<���<���<Y��<n�<��<��<��<5!�<�!�<8�<��<�<"�<���<h��<x��<��<ٖ�<v�<�Q�<D)�<��<��<��<�`�<�$�<g��<��<SW�<�
�<o��<<d�<�
�<���<K�<���<hz�<��<$��<O"�<w��<�(�<���<�<��<K�<Et�<�ޮ<�E�<"��<T	�<;f�<��<��<�j�<u��<�	�<FU�<F��<��<J)�<pk�<y��<��<�%�<F`�<+��<nЌ<m�<;�<\n�<���<�у<��<A2�<��|<�y<|u<��q<�2n<	�j<��f<_Dc<�_<w�[<�YX<(�T<Q<%yM<K�I<"AF<q�B< ?<I~;<t�7<k_4<��0<�M-<��)<2K&<��"</Y<��<�y<3<=�<�P<��
<��<�Z<"<���;�:�;T��;��;q;�;2�;���;���;Ӷ�;���;�ҽ;H��;.0�;x�;�Ц;b:�;��;.A�;^ސ;Ќ�;�L�;R�;��w;��m; �c;#Z;�dP;��F;�^=;a4;�*;b�!;��;��;G;�X�:�\�:=��:�	�:{��:��:���:Պ:Åv:��W:�K9:�1:A��9}�9���9��9�8�H����;��s��G�̹ő�H��+�7��(R�c�l�Or��_~��^t���T���!����ú�к
ݺY�����@��n�ɕ������}����%�,�,2��8��>��D��J�P��V�*�[���a�/�g���m�8�s�ݬy�l��Ƃ�ӽ��H���Ǯ��*���-����䘗������  �  _n=m=E�=�M=O�=y�=V+=�� =Ch =A =�G�<G��<
��<���<-�<1d�<z��<���<��<�6�<�h�<���<��<O��<$�<�O�<my�<ˡ�<���<���<��<�2�<)R�<�o�<���<A��<���<���<���<a��<n�<��<��<��<H!�<�!�<?�<��<��<)�<���<t��<o��<���<Ֆ�<v�<�Q�<=)�<��<���<���<�`�<�$�<Y��<��<YW�<�
�<���<=d�<�
�<���<K�<���<iz�<��< ��<V"�<w��<�(�<ǥ�<�<���<D�<Lt�<�ޮ<�E�<0��<S	�<@f�<���<��<�j�<|��<�	�<;U�<R��<��<K)�<fk�<~��<��<�%�<R`�<!��<xЌ<R�<�:�<_n�<���<҃<��<G2�<��|<�y<#|u<��q<�2n<��j<�f<RDc<�_<~�[<�YX<5�T<�Q<7yM<I�I<AAF<u�B<?<D~;<;�7<z_4<��0<�M-<��)<.K&<��"<Y<��<�y<K<*�<�P<��
<��<�Z<�<���;�:�;z��;:��;u;�;S�;`��;���;Ѷ�;���;�ҽ;>��;Y0�;x�;�Ц;h:�;4��;-A�;cސ;쌋;�L�;��;��w;�m;~�c;�Z;�dP;�F;c_=;4;=�*;B�!;q�;��;�F;Y�:&\�:��:�	�:���:/��:_��:nՊ:<�v:��W:�K9:�2:G��9S�9蠅9S�9�.8sL���;��s��l�̹Ԑ�t��
�7��)R�x�l�r���}��|s���T���!���ú0�кEݺ��w���@�gn�4������U����%�<,��2�58��>��D��J��
P��V���[���a���g���m�*�s���y�M���ł�����ᮋ�������蜔�˘�������  �  ^n=e=E�=�M=N�=}�=[+=� =;h =A =�G�<C��<��<���<-�<0d�<���<���<��<�6�<�h�<���<"��<R��<$�<�O�<cy�<���<���<���<��<{2�<%R�<�o�<���<I��<���<���<���<b��<f�<��<��<��<P!�<�!�<A�<��<�<8�<���<|��<h��<���<Ֆ�<v�<�Q�<@)�<&��<���<���<�`�<�$�<o��<���<^W�<~
�<���<+d�<�
�<���<�J�<���<cz�<��<��<Z"�<s��<�(�<ƥ�<�<���<5�<It�<�ޮ<�E�<,��<F	�<Cf�<��<��<�j�<p��<�	�<0U�<_��<��<U)�<hk�<���<��<�%�<U`�<��<�Ќ<^�<�:�<^n�<���<҃<~�<C2�<��|<�y<|u<��q<3n<�j<1�f<IDc<�_<x�[<�YX<C�T<�Q<4yM<)�I<AAF<b�B<�?<R~;<O�7<�_4<��0<�M-<��)<%K&<�"<Y<�<�y<g<�<�P<��
<��<�Z<<���;x:�;^��;��;G;�;N�;)��;���;���;���;�ҽ;,��;{0�;�w�;�Ц;R:�;7��;A�;]ސ;ό�;YL�;��;;�w;*�m;��c;Z;IeP;�F;�_=;�4;b�*;E�!;��;;�;�F;�Y�:�[�:���:~�:!��:���:Ɨ�:�Պ:ۃv:üW:�I9:1:2��9t�9u��9F�9?18�V��b�;��t����̹���:���7�f+R�ןl��r���~���s���U��U!����ú
�к�ݺ�����NA��m�3��ʶ���8����%�A,��2��8��>�,D��J��
P��V�x�[�h�a��g���m��s�Ьy�b���ł�	���ݵ��󮋻���*�����������ܕ���  �  _n=m=E�=�M=O�=y�=V+=�� =Ch =A =�G�<G��<
��<���<-�<1d�<z��<���<��<�6�<�h�<���<��<O��<$�<�O�<my�<ˡ�<���<���<��<�2�<)R�<�o�<���<A��<���<���<���<a��<n�<��<��<��<H!�<�!�<?�<��<��<)�<���<t��<o��<���<Ֆ�<v�<�Q�<=)�<��<���<���<�`�<�$�<Y��<��<YW�<�
�<���<=d�<�
�<���<K�<���<iz�<��< ��<V"�<w��<�(�<ǥ�<�<���<D�<Lt�<�ޮ<�E�<0��<S	�<@f�<���<��<�j�<|��<�	�<;U�<R��<��<K)�<fk�<~��<��<�%�<R`�<!��<xЌ<R�<�:�<_n�<���<҃<��<G2�<��|<�y<#|u<��q<�2n<��j<�f<RDc<�_<~�[<�YX<5�T<�Q<7yM<I�I<AAF<u�B<?<D~;<;�7<z_4<��0<�M-<��)<.K&<��"<Y<��<�y<K<*�<�P<��
<��<�Z<�<���;�:�;z��;:��;u;�;S�;`��;���;Ѷ�;���;�ҽ;>��;Y0�;x�;�Ц;h:�;4��;-A�;cސ;쌋;�L�;��;��w;�m;~�c;�Z;�dP;�F;c_=;4;=�*;B�!;q�;��;�F;Y�:&\�:��:�	�:���:/��:_��:nՊ:<�v:��W:�K9:�2:G��9S�9蠅9S�9�.8sL���;��s��l�̹Ԑ�t��
�7��)R�x�l�r���}��|s���T���!���ú0�кEݺ��w���@�gn�4������U����%�<,��2�58��>��D��J��
P��V���[���a���g���m�*�s���y�M���ł�����ᮋ�������蜔�˘�������  �  [n=n=>�=�M=N�=z�=d+=�� =Hh =; =�G�<I��<��<���<-�<?d�<n��<���<��<�6�<�h�<���<0��<M��<$�<~O�<by�<ʡ�<~��<���<��<�2�<#R�<�o�<���<6��<���<���<���<Y��<n�<��<��<��<5!�<�!�<8�<��<�<"�<���<h��<x��<��<ٖ�<v�<�Q�<D)�<��<��<��<�`�<�$�<g��<��<SW�<�
�<o��<<d�<�
�<���<K�<���<hz�<��<$��<O"�<w��<�(�<���<�<��<K�<Et�<�ޮ<�E�<"��<T	�<;f�<��<��<�j�<u��<�	�<FU�<F��<��<J)�<pk�<y��<��<�%�<F`�<+��<nЌ<m�<;�<\n�<���<�у<��<A2�<��|<�y<|u<��q<�2n<	�j<��f<_Dc<�_<w�[<�YX<(�T<Q<%yM<K�I<"AF<q�B< ?<I~;<t�7<k_4<��0<�M-<��)<2K&<��"</Y<��<�y<3<=�<�P<��
<��<�Z<"<���;�:�;T��;��;q;�;2�;���;���;Ӷ�;���;�ҽ;H��;.0�;x�;�Ц;b:�;��;.A�;^ސ;Ќ�;�L�;R�;��w;��m; �c;#Z;�dP;��F;�^=;a4;�*;b�!;��;��;G;�X�:�\�:=��:�	�:{��:��:���:Պ:Åv:��W:�K9:�1:A��9}�9���9��9�8�H����;��s��G�̹ő�H��+�7��(R�c�l�Or��_~��^t���T���!����ú�к
ݺY�����@��n�ɕ������}����%�,�,2��8��>��D��J�P��V�*�[���a�/�g���m�8�s�ݬy�l��Ƃ�ӽ��H���Ǯ��*���-����䘗������  �  ]n=m=E�=�M=P�=r�=[+=�� =Bh == =�G�<C��<��<���<-�<8d�<n��<���<��<�6�<�h�<���<��<B��< $�<�O�<gy�<̡�<���<���<��<}2�<.R�<�o�<���<>��<���<���<���<_��<j�<��<��<��<J!�<�!�<6�<��<�<#�<���<o��<q��<��<Ֆ�<v�<�Q�<B)�<��<���<��<�`�<�$�<b��<��<PW�<�
�<���<;d�<�
�<���<�J�<���<hz�<��<#��<T"�<x��<�(�<˥�<�<���<@�<Mt�<�ޮ<�E�<.��<W	�<5f�<���<��<�j�<t��<�	�<=U�<F��<��<A)�<nk�<v��<��<�%�<L`�<!��<xЌ<^�<�:�<^n�<���<҃<��<C2�<��|<�y<|u<��q<3n<�j<�f<YDc<"�_<��[<�YX<2�T<�Q</yM<G�I<?AF<y�B<?<&~;<P�7<�_4<��0<�M-<��)<%K&<��"<(Y<��<�y<4<+�<�P<��
<��<�Z<�<{��;�:�;z��;#��;x;�;M�;U��;���;���;ļ�;�ҽ;M��;O0�;x�;�Ц;j:�;+��;A�;|ސ;݌�;�L�;��;��w;��m;=�c;�Z;�dP;r�F;;_=;*4;��*;B�!;��;��;G;�X�:H\�:ė�:>	�:8��:���:��:�Ԋ:хv:N�W:�K9:O2:u��9��9䠅9��978-I��k�;��s���̹k�� ����7�*R�n�l�r��.~���s���T��;"��	�ú��кݺj�麔���@��n����h���������%��,��2�88��>�0D�'J��
P��V���[���a��g���m�*�s�׬y�P���ł�ܽ�����Ү������������И�������  �  `n=g=E�=�M=T�=|�=X+=�� =?h =? =�G�<G��<��<���<-�<6d�<}��<���<��<�6�<�h�<���<��<\��<$�<O�<hy�<���<���<���<��<}2�<2R�<�o�<���<@��<���<���<���<i��<i�<��<��<��<K!�<�!�<O�<��<�<(�<���<x��<l��<���<Ӗ�<v�<�Q�<>)�<!��<���<���<�`�<�$�<b��<���<kW�<~
�<���<4d�<�
�<���<�J�<���<`z�<��<��<V"�<v��<�(�<ϥ�<�<���<<�<Pt�<�ޮ<�E�<)��<P	�<Of�<���<��<�j�<{��<�	�<<U�<V��<��<G)�<jk�<~��<��<�%�<P`�<��<|Ќ<X�< ;�<nn�<���<҃<��<H2�<��|<�y</|u<��q<3n<�j<�f<BDc<�_<��[<�YX<C�T<�Q<;yM<.�I<AAF<\�B<?<Q~;<C�7<�_4<��0<�M-<��)<-K&<��"<!Y<��<�y<R<+�<�P<��
<��<�Z<�<��;�:�;W��;#��;K;�;f�;E��;���;���;Լ�;�ҽ;5��;W0�;�w�;�Ц;J:�;R��;A�;fސ;݌�;�L�;��;,�w;��m;��c;�Z;�dP;{�F;}_=;�4;N�*;6�!;k�;��;�F;VY�:
\�:G��:�	�:���:ʊ�:���:�֊:�v:��W:�J9:�1:��9E�9���9��9�;8�M��o�;�It����̹ۏ����C�7��*R��l��r��a~���s���T��� ���ú~�к�ݺ���m���@�Cn���9�����\����%�:,��2�c8��>�[D��J�s
P�V�{�[�7�a���g�	�m��s���y�`���ł�	������ ���������ܜ������ϕ���  �  `n=k=H�=�M=L�=x�=_+=�� =Dh => =�G�<E��<��<���<-�<6d�<p��<���<��<�6�<�h�<���<#��<M��<$�<�O�<uy�<š�<���<���<��<�2�<'R�<�o�<���<>��<���<���<���<c��<o�<��<��<��<J!�<�!�<9�<��<
�<�<���<l��<m��<��<Ԗ�<v�<�Q�<A)�<��<���<��<�`�<�$�<h��<���<VW�<�
�<���<Ad�<�
�<���<K�<���<hz�<��<)��<T"�<x��<�(�<ƥ�<�<���<D�<Mt�<�ޮ<�E�<+��<L	�<=f�<��<��<�j�<w��<�	�<=U�<G��<��<E)�<fk�<{��<��<�%�<J`�<$��<uЌ<c�<�:�<Zn�<���<҃<��<I2�<��|<�y<%|u<��q<3n<�j<�f<cDc< �_<{�[<�YX<9�T<�Q<:yM<A�I<MAF<h�B<�?<?~;<]�7<y_4<��0<�M-<z�)<)K&<��"<Y<��<�y<7<,�<�P<��
<��<�Z<<���;�:�;b��;Y��;[;�;Z�;a��;���;Ͷ�;���;�ҽ;M��;M0�;)x�;�Ц;]:�;;��;3A�;Xސ;ڌ�;�L�;��;W�w;��m;��c;Z;�dP;��F;#_=;4;�*;=�!;H�;��;�F;�X�:!\�:}��:�	�:��: ��:嗚:,Պ:r�v:�W:fL9:�1:���9�9�9��948�C��t�;��s��?�̹�����[�7��)R�f�l��r���}���s��*U���!��\�úq�к�ݺ<��<���@��n����G����u����%�T,�2�"8��>�D��J�P��V�v�[���a���g���m��s���y�b���ł�ǽ������������$���朔�Ø�������  �  \n=l=A�=�M=R�=u�=\+=�� =Gh =; =�G�<>��<��<���<�,�<;d�<l��<���<��<�6�<�h�<���< ��<D��<,$�<�O�<dy�<š�<���<���<��<�2�<(R�<�o�<���<8��<���<���<���<]��<x�<��<��<��<=!�<�!�<8�<��<�<�< ��<f��<u��<��<ۖ�<v�<�Q�<H)�<��<��<��<�`�<�$�<_��<��<PW�<�
�<w��<:d�<�
�<���<	K�<���<pz�<��<-��<Q"�<y��<�(�<ť�<�<���<N�<Ht�<�ޮ<�E�<&��<e	�<4f�<��<��<�j�<}��<�	�<?U�<C��<��<9)�<jk�<{��<��<�%�<E`�<+��<mЌ<\�<�:�<bn�<���<҃<��<@2�<��|<�y<|u<��q<�2n<�j<�f<hDc<�_<��[<�YX<;�T<Q<*yM<A�I</AF<}�B<?<2~;<S�7<f_4<��0<�M-<��)<K&<��"<&Y<��<�y<0<,�<�P<��
<��<�Z<<���;�:�;`��;��;\;�;>�;���;���;ݶ�;���;�ҽ;S��;40�;<x�;�Ц;�:�;��;SA�;fސ;Ɍ�;�L�;r�; x;��m;�c;�Z;gdP;��F;�^=;C4;��*;m�!;:�;��;3G;X�:�\�:.��:�	�:寺:���:���:�Ԋ:��v:��W:|K9:�1:���9-�92��9��9g&8�?���;��s��V�̹5��ģ�
�7�R(R��l�zr��N~��!t���S��B"����ú$�к�ݺ��.���@��n�ȕ������r��F�%�!,�62��8�>�AD�J��
P�QV���[���a�4�g���m���s�Ԭy�.���ł�����=�������������휔����������  �  an=n=D�=�M=N�=|�=\+=�� =Bh =; =�G�<;��<��<���<-�<9d�<s��<���<��<�6�<�h�<���<#��<S��<$�<|O�<jy�<͡�<���<���<��<~2�<2R�<�o�<���<B��<���<���<���<]��<q�<��<��<��<E!�<�!�<?�<��<�<!�<���<m��<o��<��<ז�<v�<�Q�<D)�<��<���<��<�`�<�$�<^��<���<ZW�<�
�<~��<@d�<�
�<���<K�<���<jz�<��<'��<W"�<y��<�(�<ϥ�<�<���<H�<Lt�<�ޮ<�E�<%��<N	�<Bf�<
��<��<�j�<u��<�	�<6U�<I��<��<@)�<hk�<y��<��<�%�<H`�<!��<uЌ<\�<;�<`n�<���<҃<��<K2�<��|<�y<|u<��q<3n<	�j<�f<`Dc<�_<��[<�YX<C�T<�Q<>yM<I�I<>AF<]�B< ?<P~;<Q�7<w_4<��0<�M-<��)<K&<��"<"Y<��<�y<=<�<�P<��
<��<�Z<<���;�:�;H��;+��;|;�;W�;j��;���;���;Ӽ�;�ҽ;H��;]0�; x�;�Ц;s:�;��;8A�;Zސ;�;�L�;��;J�w;�m;��c;�Z;�dP;w�F;$_=;4;��*;R�!;A�;��;G;}X�:\�:���:a	�:��:���:��:qՊ:b�v:w�W:JL9:�2:���9��9⠅9U�9�58�F����;��s����̹���ʤ�N�7�&)R���l�
r���}��5t��U��o!��I�ú��к�ݺb����� A��n���m�������W�%�3,�#2�78��>�@D�xJ��
P��V���[���a���g���m��s�ݬy����ł�ӽ�����Ů����������������������  �  dn=g=I�=�M=L�=x�=X+=�� =@h =? =�G�<A��<��<���<-�<)d�<r��<���<��<�6�<�h�<���<��<S��<$�<�O�<ry�<ġ�<���<���<��<2�<7R�<�o�<���<E��<���<��<���<k��<u�<��<��<��<Y!�<�!�<=�<��<��<$�<���<u��<e��<��<Ӗ�<v�<�Q�<<)�<��<���<���<�`�<�$�<^��<��<ZW�<�
�<���<:d�<�
�<���<K�<���<iz�<��<$��<Z"�<~��<�(�<֥�<�<���<C�<Tt�<�ޮ<�E�<<��<H	�<Cf�<���<��<�j�<p��<�	�<3U�<J��<��<C)�<^k�<y��<��<�%�<Q`�<��<wЌ<V�<�:�<\n�<���<҃<��<P2�<��|<�y<,|u<��q<3n<
�j<�f<aDc<0�_<��[<�YX<G�T<�Q<JyM<.�I<RAF<{�B<�?<@~;<A�7<x_4<��0<�M-<��)<!K&<��"<Y<��<ry<:<�<�P<��
<��<�Z<�<���;x:�;���;I��;V;�;q�;J��;���;Ķ�;��;�ҽ;Y��;f0�;x�;�Ц;o:�;Y��;FA�;fސ;茋;�L�;��;T�w;�m;a�c;�Z;�dP;4�F;e_=;�4;�*;-�!;9�;��;�F;�X�:�[�:��:��:Y��:���:3��:fՊ:�v:$�W:wK9:;2:m��9��9Z��9��9 O8kI����;�nr����̹�����7��)R���l�~r���}���r��nU��`!���ú��к�ݺ���o��9A��n�^��[��^������%�F,��2�m8��>�mD��J�P��V�=�[�@�a���g��m�߼s���y�!���ł�ѽ�����î��駎�������������ϕ���  �  cn=j=>�=�M=S�=x�=^+=�� =Bh =9 =�G�<?��<��<���<-�<4d�<t��<���<��<�6�<�h�<���<��<P��<"$�<~O�<^y�<ǡ�<���<���<��<�2�</R�<�o�<���<A��<���<���<���<f��<n�<��<��<��<?!�<�!�<B�<��<
�<#�<���<i��<l��<��<і�<v�<�Q�<=)�<��<���<��<�`�<�$�<e��<���<]W�<�
�<x��<3d�<�
�<���<�J�<���<lz�<��<'��<\"�<���<�(�<ͥ�<�<���<C�<Ot�<�ޮ<�E�<$��<Y	�<Af�<��<��<�j�<p��<�	�<:U�<L��<��<A)�<fk�<z��<��<�%�<D`�<��<pЌ<b�<�:�<gn�<���<҃<��<O2�<��|<�y<5|u<��q<�2n<�j<�f<hDc<�_<��[<�YX<=�T<�Q<EyM<;�I<#AF<r�B<?<=~;<Y�7<j_4<��0<�M-<z�)<K&<��"<Y<��<�y<><!�<�P<��
<��<�Z<�<���;�:�;O��;���;d;�;b�;[��;���;��;ļ�;�ҽ;i��;U0�;x�;�Ц;t:�;E��;,A�;mސ;茋;�L�;w�;��w;*�m;��c;�Z;�dP;X�F;_=;�4;��*;"�!;B�;��;�F;�X�:\�:_��:	�:b��:ꊪ:���:�Պ:օv:��W:�J9:12:���9q�9_��9C�9�18&F����;��q����̹M����ހ7��)R�1�l�er���~��Jt��`T��~!����ú׃кDݺ�����A��n���i����}��%�%�S,�C2�K8��>�D��J��
P��V��[��a���g���m��s�{�y�#���ł�Ƚ���������������Ĝ�����������  �  ^n=t=F�=�M=P�=r�=^+=�� =Fh =7 =�G�<9��<���<���<�,�<5d�<g��<���<��<�6�<�h�<���<&��<<��<"$�<|O�<uy�<ա�<���<���<��<�2�<4R�<�o�<���<H��<���<���<���<^��<p�<��<��<��<C!�<�!�<3�<��<�<�<���<^��<q��<��<ϖ�<v�<�Q�<>)�<	��<���<���<�`�<�$�<`��<���<JW�<�
�<{��<Ld�<�
�< ��<K�<���<uz�<��<+��<^"�<���<�(�<Х�<�<���<L�<Lt�<�ޮ<�E�<%��<Y	�<,f�<
��<��<�j�<s��<�	�<7U�<?��<��<7)�<fk�<s��<��<�%�<<`�<)��<iЌ<a�<�:�<^n�<���<҃<��<C2�<��|<�y<#|u<��q<�2n<�j<$�f<pDc<�_<��[<�YX<8�T<Q<1yM<b�I<EAF<j�B<?<'~;<[�7<`_4<��0<�M-<�)<K&<��"<Y<��<�y<%<�<�P<��
<��<�Z<<_��;�:�;H��;U��;�;�;A�;���;���;߶�;ۼ�;�ҽ;l��;s0�;3x�;�Ц;�:�;$��;3A�;�ސ;֌�;�L�;��;��w;��m;y�c;�Z;WdP;��F;�^=; 4;��*;�!;;�;��;�F;�W�:1\�:���:�	�:ϯ�:���:���:jԊ:��v:�W:�M9:v2:���9��9V��9��9N28�B����;��q����̹Տ����܁7��(R���l��q��M}��?t��cT���"��M�ú�к�ݺ���]��A�o�����������l�%�3,��2��8�!>�D�J��
P��V���[�l�a��g���m��s�ìy����ł����������������ꡑ�㜔�Ę�������  �  `n=e=F�=�M=R�=y�=^+=�� =Bh =; =�G�<=��< ��<���<-�</d�<n��<���<��<�6�<�h�<���<%��<O��<"$�<�O�<my�<���<���<���< �<�2�<8R�<�o�<���<I��<���<���<���<j��<t�<��<��<��<H!�<�!�<C�<��<
�<!�<���<g��<p��<��<і�<v�<�Q�<<)�<��<���<��<�`�<�$�<g��<���<[W�<�
�<���<8d�<�
�<��<K�<���<jz�<��<"��<_"�<~��<�(�<ե�<�<���<E�<Tt�<�ޮ<�E�<+��<W	�<@f�<��<��<�j�<r��<�	�<9U�<G��<��<C)�<bk�<x��<��<�%�<F`�<"��<sЌ<a�<�:�<fn�<���<҃<��<E2�<��|<�y<*|u<��q<3n<��j<$�f<VDc<-�_<��[<�YX<N�T<�Q<;yM<(�I<CAF<k�B<?<C~;<Z�7<q_4<��0<�M-<��)<K&<��"<Y<��<~y<2<!�<�P<��
<��<�Z<
<���;�:�;Z��;4��;6;�;h�;^��;���;ʶ�;��;�ҽ;M��;x0�;x�;�Ц;j:�;T��;EA�;�ސ;���;�L�;��;~�w;/�m;��c;�Z;�dP;|�F;�^=;4;��*;!�!;B�;��;�F;PX�:(\�:T��:n	�:%��:��:Ǘ�:�Պ:&�v:�W:*K9:1:���9��9֣�91�9dD8�K��a�;�xr���̹B�����S�7��)R���l�
s��~���s���T���!��n�ú��к�ݺ������
A��n�8��Z��@�����D�%�2,�-2�38��>�D��J��
P��V���[�A�a�
�g���m�¼s���y�"���ł�轅�����ڮ��������圔����������  �  �o=�=��=�O={�=�=.=�� =wk =�	 ='O�<I��<���<��<�6�<�n�<u��<7��<�<�C�<yv�<��<
��<��<z4�<�`�<`��<y��<��<��<%&�<wH�< i�<���<!��<���<���<7��<� �<��<]!�<�-�<�7�<�>�<C�<MD�<�B�<	>�<G6�<L+�<��<E�<��<`��<���<���<)}�<nU�<�)�<L��<���<+��<kS�<w�<I��<���<C:�<o��<"��<�:�<���<�z�<E�<w��<�:�<eǼ<!P�<�Թ<9U�<�Ѷ<NJ�<��<�/�<��<��<�l�<ϫ< .�<≨<~�<8�<���<kڡ<a'�<�q�<���<���<�A�<���<���<G��<9�<Rr�<ҩ�<�ߌ<S�<�G�<�y�<���<�ڃ<�	�<=8�<��|<,&y<�u<��q<:1n<`�j<��f<R:c<u�_<�[<�GX<w�T<J Q<+_M<<�I<�!F<�B<��><nV;<��7<m24<�0<c-<O�)<k&<��"<<��<p7<��<g<<�
<�X<b
<e� <E�;���;&�;��;y��;JG�;o�;Q��;D��;���;;�;m,�;�a�;���;5��;kg�;��;�l�;�	�;n��;�w�;�I�;�Xv;Al;�Kb;<yX;��N;I9E;M�;;H}2;�P);VC ;�U;4�;9�;���:U��:&��:�\�:��:���:��:�e�::�q:�S:t�4:��:'Y�9���9�I{9�K9�M�7�o��?�I�
C���ӹt��
��&r:��U�[Yo���6���ɩ������?��P�ĺщѺ,޺"������x����#����,�H= �1J&�FS,�W2��W8��T>�qOD��FJ��;P�:.V��\��b���g�,�m� �s���y����̂�Å�#���G�����������������������  �  �o=�=��=�O=��=�=.=�� =uk =�	 =;O�<H��<���<��<�6�<�n�<l��<A��<!�<�C�<rv�<��<��< �<�4�<�`�<Q��<k��<��<��<&�<qH�<�h�<���<.��<���<��<.��<� �<n�<e!�<�-�<�7�<�>�<�B�<RD�<�B�<>�<Q6�<F+�<��<D�<��<X��<���<��<}�<vU�<�)�<]��<���<*��<eS�<}�<^��<���<M:�<Y��<��<�:�<���<�z�</�<y��<�:�<nǼ</P�<�Թ<<U�<�Ѷ<JJ�<���<�/�<��<z�<tl�<�Ϋ<.�<艨<��<8�<���<mڡ<o'�<�q�<���<���<�A�<���<���<B��<.9�<Qr�<Ω�<�ߌ<a�<�G�<�y�<���<�ڃ<�	�<!8�<��|<,&y<�u<��q<,1n<w�j<��f<f:c<j�_<�[<�GX<l�T<j Q<�^M<5�I<�!F<�B<	�><�V;<��7<V24<�0<e-<w�)<g&<��"<&<h�<�7<��<,g<?<�
<�X<U
<�� <l�;I��;�%�;���;@��;�F�;��;��;*��;���;;�;�,�;�a�;���;��;vg�;u�;�l�;�	�;���;�w�;mI�;�Xv;kAl;lLb;�yX;v�N;89E;H�;;�}2;�P);uC ;U;��;v�;��:o��:k��:r\�:"�:\��:��:(f�:��q: S:S�4:��:FW�9v��9�>{99M9�)�7�f���I�.?���ӹ?��q��bt:�� U��[o��Ä� ������~��J?���ĺ�Ѻ�޺������	��R������,�[= �YJ&��R,�$W2��W8�U>�OD�oFJ�J;P�j.V�P\��b���g���m� �s�	�y�׭��̂�����������������Ø������Ӎ���  �  �o=�=��=�O=��=ߎ=.=�� ={k =�	 =;O�<C��<���<(��<�6�<�n�<`��<E��<�<�C�<yv�<٧�<��<��<�4�<�`�<a��<���<���<��<&�<zH�<�h�<���<&��<���<��<'��<
�<g�<r!�<�-�<�7�<�>�<�B�<YD�<�B�<
>�<B6�<A+�<��<8�<��<N��<	��<���<}�<�U�<�)�<b��<���<,��<bS�<o�<N��<��<W:�<W��<7��<�:�<���<�z�<(�<���<�:�<tǼ<P�<�Թ<=U�<�Ѷ<WJ�<���<�/�<���<��<�l�<�Ϋ<.�<҉�<��<8�<���<jڡ<d'�<�q�<w��<���<�A�<Ƃ�<���<:��<29�<Er�<ک�<�ߌ<Z�<�G�<�y�<���<�ڃ<�	�<8�<��|<1&y<�u<��q<$1n<��j<��f<h:c<f�_<-�[<�GX<f�T<� Q<�^M<l�I<�!F<�B<�><]V;<��7<I24<+�0<R-<w�)<^&<��"<I<i�<�7<��<4g<1<ڬ
<�X<A
<}� <�;_��;�%�;��;���;�F�;�;���;P��;���;9�;�,�;�a�;ߧ�;���;�g�;Y�;m�;�	�;��;gx�;gI�;�Xv;�@l;�Kb;yX;P�N;f9E;��;;~2;oP);�C ;rU;�;��;<��:Ē�:���:�\�:��:|��:��:�d�:��q:�S:�4:��:�W�9\��95;{9�V9,�7�`����I��B���ӹ������u:���T�.\o����������;~���@����ĺ��Ѻ`޺<�꺨��������9����+�W= ��J&��R,�W2��W8�AU>�;OD�GJ�y;P�T.V�?\��b��g�o�m��s�"�y�~���̂���w���������������������������  �  �o=�=��=�O=��=�=.=�� ={k =�	 =6O�<N��<���<��<�6�<�n�<f��<L��<�<�C�<zv�<��<$��<��<�4�<�`�<R��<v��<��<��<&�<{H�<�h�<���</��<���<��<#��<� �<m�<e!�<�-�<�7�<�>�<�B�<VD�<�B�<>�<Q6�<F+�<��<A�<��<\��<���<��<}�<sU�<�)�<c��<���<0��<fS�<|�<^��<��<R:�<Y��<��<�:�<���<�z�<.�<���<�:�<zǼ<"P�<�Թ<CU�<�Ѷ<TJ�<���<�/�<��<��<wl�<�Ϋ<.�<䉨<��<8�<���<pڡ<c'�<�q�<���<���<�A�<���<y��<F��<-9�<Or�<ܩ�<�ߌ<g�<�G�<�y�<���<�ڃ<�	�<%8�<��|<+&y<�u<��q<!1n<��j<��f<v:c<g�_<�[<�GX<e�T<k Q<�^M<D�I<�!F<�B<��><�V;<��7<V24<,�0<_-<m�)<t&<��"<0<q�<�7<��<Bg<(<�
<�X<U
<�� <[�;A��;�%�;���;n��;�F�;��;��;T��;q��;O�;�,�;�a�;���;���;�g�;q�;�l�;�	�;��;x�;iI�;�Xv;7Al;mLb;�yX;t�N;{9E;2�;;~2;�P);RC ;JU;Ӆ;d�;��:Ӓ�:��:�\�:5�:N��:��:�e�:�q:)S:2�4:��:W�9̭�9;>{9�Q9���7)Z��t�I��@��;ӹ���4���t:�� U�v[o�$Ä����������~���?����ĺ�Ѻ<޺ݐ��������������	��+��= �4J&��R,�2W2�~W8�U>��ND�pFJ�p;P�I.V�^\��b���g���m� �s���y����̂���\�����������՟����������э���  �  �o=�=��=�O=}�=�=	.=�� =uk =�	 =1O�<I��<���<��<�6�<�n�<n��<A��<�<�C�<qv�<��<��<��<4�<�`�<W��<s��<��<��<&�<sH�<�h�<���<&��<���<��<*��<� �<n�<b!�<�-�<�7�<�>�<�B�<JD�<�B�<>�<J6�<F+�<��<H�<
��<_��<���<���<)}�<tU�<�)�<T��<���<*��<dS�<x�<O��<��<C:�<j��<��<�:�<���<�z�</�<}��<�:�<kǼ<P�<�Թ<:U�<�Ѷ<LJ�<���<�/�<��<��<xl�<�Ϋ<.�<䉨<��<8�<���<rڡ<h'�<�q�<���<���<�A�<�<}��<D��<$9�<Yr�<ͩ�<�ߌ<W�<�G�<�y�<���<�ڃ<�	�<28�<��|<%&y<�u<��q<(1n<r�j<��f<[:c<k�_<�[<�GX<e�T<c Q<_M<>�I<�!F<�B<��><�V;<��7<W24<�0<t-<c�)<i&<��"<8<��<�7<��<+g</<�
<�X<X
<p� <\�;��;&�;���;a��;%G�;��;��;2��;���;7�;�,�;�a�;���;��;�g�;t�;�l�;�	�;B��;�w�;�I�;vXv;"Al;Lb;[yX;v�N;'9E;g�;;�}2;�P);\C ;�U;6�;h�;]��:���:k��:p\�:�:
��:	�:�e�:M�q:JS:��4:��:>X�9]��9�>{9O9��7'i���I��A��sӹ���8���t:��U�]Zo�:Ä������������?����ĺ��Ѻ�޺���p�����=��������+�u= �CJ&��R,��V2��W8�U>�SOD��FJ��;P�.V��\��b�J�g���m�9�s��y����̂���Y���6���������Ę������ፚ��  �  �o=�=��=�O=��=�=	.=�� =xk =�	 =8O�<O��<���<$��<�6�<�n�<l��<I��<�<�C�<zv�<��<��<��<�4�<�`�<T��<z��<���<��<&�<qH�<�h�<���<*��<���<��<$��<� �<f�<l!�<�-�<�7�<�>�<�B�<KD�<�B�<>�<O6�<W+�<��<?�<��<\��<��<��<}�<xU�<�)�<d��<���<*��<sS�<��<O��<���<F:�<V��<��<�:�<���<�z�<'�<z��<�:�<mǼ<%P�<�Թ<6U�<�Ѷ<JJ�<���<�/�<���<��<vl�<�Ϋ<.�<牨<��<&8�<���<kڡ<h'�<�q�<���<���<�A�<Ă�<���<G��<-9�<Lr�<Щ�<�ߌ<W�<�G�<�y�<���<�ڃ<�	�< 8�<��|<2&y<�u<��q<1n<v�j<��f<a:c<[�_<"�[<�GX<o�T<i Q<�^M<N�I<�!F<��B<
�><|V;<��7<~24<�0<[-<q�)<u&<��"<B<g�<�7<��<;g<4<�
<�X<t
<p� <]�;?��;�%�;���;���;�F�;��;��;.��;���;�;�,�;�a�;���;���;�g�;V�;�l�;�	�;��;x�;gI�;�Xv;�Al;�Kb;~yX;��N;39E;!�;;~2;�P);�C ;dU;��;��;'��:ڒ�:���:n\�:�:���:
�:Yf�:��q:�S:�4:��:$V�9Ϯ�9R;{9�M9��7�g����I��@��Iӹ���j���t:�� U�]\o�Ä�����6�����a?����ĺ%�Ѻ޺+��u������W�������+�== �-J&��R,�CW2��W8�{T>�VOD��FJ�:;P��.V�L\��b���g���m��s�G�y�����̂���H���*�����������Ԙ������Ս���  �  �o=�=��=�O=��=�=.=�� =xk =�	 =AO�<S��<���<*��<�6�<�n�<b��<S��<�<�C�<wv�<��<��<��<�4�<�`�<T��<|��< ��<��<&�<}H�<�h�<���<*��<���<	��<��<�<g�<c!�<�-�<�7�<�>�<�B�<ZD�<�B�<>�<Q6�<H+�<��<?�<#��<X��<��<���<&}�<~U�<�)�<n��<���<2��<fS�<}�<V��<��<T:�<[��<"��<�:�<���<�z�<(�<���<�:�<nǼ<P�<�Թ<6U�<�Ѷ<VJ�<���<�/�< ��<��<wl�<�Ϋ<.�<ቨ<��<8�<���<pڡ<h'�<�q�<}��<���<�A�<ʂ�<}��<I��<89�<Pr�<ԩ�<�ߌ<a�<�G�<�y�<���<�ڃ<�	�< 8�<��|<!&y<�u<��q<
1n<~�j<��f<h:c<M�_<%�[<�GX<\�T<e Q<�^M<Q�I<�!F<!�B<�><{V;<��7<U24<�0<e-<��)<&<��"<N<t�<�7<��<Og<:<�
<�X<V
<�� <L�;Y��;&�;���;���;�F�;��;���;^��;}��;�;�,�;�a�;ȧ�;���;�g�;[�;�l�;�	�;��;x�;tI�;�Xv;<Al;*Lb;�yX;��N;w9E;#�;;\~2;�P);�C ;�U;�;��;�:���:
��:�\�:>�:f��:|�:�e�:[�q:�S:��4:��:?V�9���9|;{9�T9�7/f����I��A��Eӹ���ڲ�}u:�� U�\o�����������i~���?��[�ĺ׉Ѻg޺А�s���q�����U����h+�v= � J&�TR,�&W2��W8�U>��ND��FJ�V;P�.V�h\�{b���g���m�H�s�
�y����	͂���r������ϧ����������˒��ݍ���  �  �o=�=��=�O=z�=�=.=�� =yk =�	 =6O�<R��<���<&��<�6�<�n�<l��<N��<�<�C�<yv�<��<��<��<|4�<�`�<O��<s��<��<��<&�<rH�<�h�<���<$��<���<��<$��<� �<h�<]!�<�-�<�7�<�>�<�B�<ND�<�B�<>�<N6�<D+�<��<B�<��<`��<��<���<,}�<}U�<�)�<`��<���<4��<dS�<{�<R��<��<F:�<e��<��<�:�<���<�z�<&�<}��<�:�<gǼ<P�<�Թ<7U�<�Ѷ<LJ�<���<�/�<��<��<rl�<�Ϋ<.�<މ�<��<8�<���<xڡ<e'�<�q�<���<���<�A�<Ȃ�<~��<K��<,9�<Yr�<֩�<�ߌ<`�<�G�<�y�<���<�ڃ<�	�<28�<��|<&y<�u<��q<1n<s�j<��f<]:c<e�_<�[<�GX<R�T<f Q<_M<;�I<�!F< �B<��><�V;<��7<P24<#�0<w-<m�)<~&<��"<F<��<�7<��<Gg</<��
<�X<Y
<�� <S�;��;&�;���;c��;.G�;��;���;2��;��;5�;z,�;ya�;���;���;�g�;^�;�l�;�	�;A��;�w�;�I�;�Xv;�@l;"Lb;wyX;n�N;�9E;>�;;�}2;Q);�C ;�U;K�;��;H��:���:��:]�:�:;��:G�:Xe�:��q:�S:��4:��:&Y�9���9�:{9VO9` �7m����I�.C��ӹC��,���u:��U�Zo�<Ä�6�!���t���?����ĺ��ѺV޺L�꺒������Z��l����}+�r= �J&��R,��V2��W8�*U>�OD��FJ��;P�+.V�E\��b�O�g���m�n�s�2�y����̂�������1�������ȟ��͘��ߒ��ۍ���  �  �o=�=��=�O=��=�=
.=�� =xk =�	 =9O�<P��<���<#��<�6�<�n�<q��<I��<�<�C�<wv�<���<��<
�<�4�<�`�<S��<r��<���<��<&�<gH�<�h�<���<#��<���<���<(��<� �<i�<d!�<�-�<�7�<�>�<�B�<ID�<�B�<>�<O6�<S+�<��<F�<��<c��<��<���<%}�<{U�<�)�<c��<���<+��<oS�<�<P��<���<C:�<]��<��<�:�<���<�z�<+�<n��<�:�<bǼ<#P�<�Թ<0U�<�Ѷ<?J�<���<�/�<���<��<vl�<�Ϋ<.�<���<��<(8�<���<pڡ<m'�<�q�<���<���<�A�<ł�<���<J��<.9�<Wr�<ө�<�ߌ<W�<�G�<�y�<���<�ڃ<�	�<"8�<��|<,&y<�u<��q< 1n<g�j<��f<R:c<_�_<
�[<�GX<j�T<X Q<�^M<:�I<�!F<�B<��><�V;<��7<|24<�0<o-<t�)<x&<��"<A<��<�7<��<=g<<<�
<�X<x
<r� <��;��;�%�;���;a��;�F�;��;��;��;|��;�;w,�;�a�;���;���;Yg�;d�;�l�;�	�;��;�w�;|I�;sXv;�Al;%Lb;�yX;��N;:9E;_�;;~2;Q);�C ;�U;�;��;���:Ӓ�:t��:�\�:��:~��:'�:�f�:L�q:�S:}�4:Z�:�U�9M��9�={9�G9D�7�q��7�I�'B���ӹ��ɵ�it:�1U�<\o�lÄ�����爵�q���>����ĺ �Ѻ@޺א����ȭ�/��t�����+�2= �J&��R,��V2��W8��T>�ROD�gFJ�Z;P��.V�?\��b���g��m��s�J�y�!���̂�Å�D���G�������⟑��������������  �  �o=�=��=�O=��=�=.=�� =zk =�	 =BO�<J��<���<1��<�6�<�n�<l��<I��<#�<�C�<yv�<��<��<��<�4�<�`�<Y��<���<���<��<&�<qH�<�h�<���<��<���<���< ��<� �<d�<c!�<�-�<�7�<�>�<�B�<WD�<�B�<>�<N6�<K+�<��<E�< ��<Z��<��<���<)}�<�U�<�)�<i��<���<1��<iS�<|�<S��<��<Q:�<\��<*��<�:�<���<�z�<'�<}��<�:�<aǼ<P�<�Թ<.U�<�Ѷ<KJ�<���<�/�<���<��<l�<�Ϋ<.�<߉�<��<8�<���<rڡ<m'�<�q�<���<���<�A�<ς�<���<D��<79�<Tr�<ة�<�ߌ<Z�<�G�<�y�<���<�ڃ<�	�<!8�<��|<&y<�u<��q<1n<a�j<��f<J:c<S�_<�[<�GX<U�T<p Q<�^M<a�I<�!F<�B<��><|V;<��7<a24<'�0<n-<��)<n&<��"<\<�<�7<��<>g<E<��
<�X<^
<~� <R�;A��;�%�;���;���;�F�;��;���;1��;|��;�;`,�;|a�;���;���;�g�;P�;�l�;�	�;��;5x�;{I�;�Xv;Al;'Lb;yX;��N;�9E;Q�;;?~2;�P);�C ;�U;4�;�;��:>��:k��:�\�:u�:U��:S�:|e�:�q:�S:��4:��:OV�9#��9�;{9O9���7<r����I�FD��Eӹa��D��Nu:�� U�[\o���^��������~���?����ĺ��ѺE޺���������a�������@+�= �GJ&�_R,�W2��W8��T>�;OD��FJ��;P�G.V�B\�>b���g���m�f�s�Z�y�ʭ��̂�Å�t���V���ħ����֘��ْ��ō���  �  �o=�=�=�O=~�=�=.=�� =�k =�	 =>O�<X��<���<)��<�6�<�n�<o��<W��<�<�C�<�v�<ݧ�<-��<��<�4�<�`�<C��<s��<���<��<&�<wH�<�h�<���<&��<���<��<��<� �<c�<]!�<�-�<�7�<�>�<�B�<^D�<�B�<(>�<S6�<G+�<�<?�<$��<`��<	��<���<!}�<�U�<�)�<q��<���<@��<iS�<}�<i��<��<W:�<M��<��<�:�<���<�z�<!�<z��<{:�<qǼ<P�<�Թ<<U�<�Ѷ<NJ�<쾳<�/�<���<{�<jl�<�Ϋ<.�<މ�<��<8�<���<|ڡ<g'�<�q�<���<���<�A�<ǂ�<���<P��<59�<Or�<驎<�ߌ<i�<�G�<�y�<���<�ڃ<�	�<8�<��|<&y<�u<��q<1n<~�j<��f<e:c<V�_<�[<�GX<K�T<p Q<�^M<I�I<o!F<�B<��><�V;<�7<I24<E�0<k-<}�)<�&<��"<L<r�<�7<��<Yg<7<��
<�X<L
<�� <Y�;?��;�%�;���;f��;�F�;��;���;F��;J��;3�;�,�;|a�;ا�;���;xg�;M�;�l�;�	�;귊;x�;7I�;Yv;Al;�Lb;�yX;��N;:E;"�;;f~2;Q);�C ;oU;��;��;\��:���:��:�]�:x�:c��:��:ne�:��q:�S:��4:Y�:zU�9
��9�8{9N9ĳ7b��W�I��B���ӹ���ٳ��v:�� U��\o��Ä�������~���?���ĺ�Ѻ�޺��y���P��?��&�����+�:= ��I&�mR,�+W2�W8�8U>��ND�5FJ��;P�.V��\��b�!�g���m���s�1�y���͂������� �������쟑�Ę���ƍ���  �  �o=�=��=�O=}�=�=.=�� =zk =�	 =9O�<R��<���<*��<�6�<�n�<s��<J��< �<�C�<yv�<��<��<��<�4�<�`�<X��<|��<���<��<&�<rH�<�h�<���<��<���<���<%��<� �<o�<_!�<�-�<�7�<�>�<�B�<SD�<�B�<>�<B6�<J+�<��<H�<��<d��<��<��<4}�<~U�<�)�<_��<���<0��<iS�<p�<L��<��<M:�<b��<(��<�:�<���<�z�<.�<u��<�:�<cǼ<P�<�Թ<4U�<�Ѷ<HJ�<���<�/�<���<��<~l�<�Ϋ<.�<���<��<8�<���<rڡ<n'�<�q�<���<���<�A�<̂�<���<M��<-9�<Xr�<ة�<�ߌ<P�<�G�<�y�<���<�ڃ<�	�<!8�<��|<&y<�u<��q<1n<\�j<��f<B:c<_�_<
�[<�GX<\�T<Y Q<�^M<R�I<�!F<"�B<��><~V;<��7<^24<&�0<u-<u�)<~&<��"<O<��<�7<��<?g<@<�
<�X<V
<n� <W�;3��;&�;���;���;�F�;��;���;1��;o��;(�;C,�;ta�;���;���;gg�;|�;�l�;�	�;��;)x�;�I�;�Xv;Al;Lb;yX;��N;w9E;n�;;�}2;$Q);�C ;�U;��;��;Ɂ�:���:���:�\�:o�:���:��:{e�:��q:kS:f�4:��:�U�9 ��9�>{9�K9���7rp���I�F���ӹӽ����u:��U�3\o���i���H������?���ĺ�Ѻ1޺������֭���i��>�U+�3= ��I&��R,��V2��W8��T>��OD��FJ��;P�.V�#\�{b���g��m�_�s��y� ���̂�Å�����f�������⟑�����˒��􍚻�  �  �o=�=�=�O=��=�=
.=�� =qk =�	 =EO�<Q��<���< ��<�6�<�n�<{��<G��<2�<�C�<pv�<���<��<�<�4�<�`�<K��<o��<��<��<&�<]H�<�h�<���<��<���<���</��<� �<b�<]!�<�-�<�7�<�>�<�B�<CD�<�B�<>�<X6�<Z+�<��<[�<��<l��<��<���<%}�<vU�<�)�<]��<���<#��<tS�<��<X��<��<@:�<Z��<��<�:�<���<�z�<&�<d��<�:�<ZǼ<$P�<�Թ<1U�<�Ѷ<5J�<���<�/�<��<}�<ll�<�Ϋ<.�<���<��<48�<���<kڡ<�'�<�q�<���<���<�A�<���<���<N��<69�<fr�<ĩ�<�ߌ<\�<�G�<�y�<���<�ڃ<�	�<)8�<��|<&y<�u<��q<-1n<M�j<��f<8:c<k�_<�[<�GX<W�T<b Q<_M<.�I<�!F<��B<�><�V;<��7<�24<�0<�-<��)<{&<��"<:<��<�7<��<9g<d<�
<�X<�
<p� <��;C��;�%�;���;U��;G�;��;��;���;���;*�;R,�;�a�;i��;��;)g�;K�;�l�;�	�;��;�w�;yI�;FXv;�Al;oLb;�yX;�N;�8E;�;;�}2;cQ);�C ;�U;�;��;L��:u��:���:	\�:�::��:��:�f�:�q:mS:��4:T�:�W�9ݫ�9;{9:C9�!�7�y����I�uC��aӹ�����t:��U�k[o��Ä��������d>����ĺ=�ѺP޺�꺪��������������+�$= ��I&�gR,�vV2�:X8�;T>�.OD�&FJ�9;P��.V�{\�b���g���m�k�s���y�W���̂�=Å�A���{�������柑����Ԓ��⍚��  �  �o=�=��=�O=}�=�=.=�� =zk =�	 =9O�<R��<���<*��<�6�<�n�<s��<J��< �<�C�<yv�<��<��<��<�4�<�`�<X��<|��<���<��<&�<rH�<�h�<���<��<���<���<%��<� �<o�<_!�<�-�<�7�<�>�<�B�<SD�<�B�<>�<B6�<J+�<��<H�<��<d��<��<��<4}�<~U�<�)�<_��<���<0��<iS�<p�<L��<��<M:�<b��<(��<�:�<���<�z�<.�<u��<�:�<cǼ<P�<�Թ<4U�<�Ѷ<HJ�<���<�/�<���<��<~l�<�Ϋ<.�<���<��<8�<���<rڡ<n'�<�q�<���<���<�A�<̂�<���<M��<-9�<Xr�<ة�<�ߌ<P�<�G�<�y�<���<�ڃ<�	�<!8�<��|<&y<�u<��q<1n<\�j<��f<B:c<_�_<
�[<�GX<\�T<Y Q<�^M<R�I<�!F<"�B<��><~V;<��7<^24<&�0<u-<u�)<~&<��"<O<��<�7<��<?g<@<�
<�X<V
<n� <W�;3��;&�;���;���;�F�;��;���;1��;o��;(�;C,�;ta�;���;���;gg�;|�;�l�;�	�;��;)x�;�I�;�Xv;Al;Lb;yX;��N;w9E;n�;;�}2;$Q);�C ;�U;��;��;Ɂ�:���:���:�\�:o�:���:��:{e�:��q:kS:f�4:��:�U�9 ��9�>{9�K9���7rp���I�F���ӹӽ����u:��U�3\o���i���H������?���ĺ�Ѻ1޺������֭���i��>�U+�3= ��I&��R,��V2��W8��T>��OD��FJ��;P�.V�#\�{b���g��m�_�s��y� ���̂�Å�����f�������⟑�����˒��􍚻�  �  �o=�=�=�O=~�=�=.=�� =�k =�	 =>O�<X��<���<)��<�6�<�n�<o��<W��<�<�C�<�v�<ݧ�<-��<��<�4�<�`�<C��<s��<���<��<&�<wH�<�h�<���<&��<���<��<��<� �<c�<]!�<�-�<�7�<�>�<�B�<^D�<�B�<(>�<S6�<G+�<�<?�<$��<`��<	��<���<!}�<�U�<�)�<q��<���<@��<iS�<}�<i��<��<W:�<M��<��<�:�<���<�z�<!�<z��<{:�<qǼ<P�<�Թ<<U�<�Ѷ<NJ�<쾳<�/�<���<{�<jl�<�Ϋ<.�<މ�<��<8�<���<|ڡ<g'�<�q�<���<���<�A�<ǂ�<���<P��<59�<Or�<驎<�ߌ<i�<�G�<�y�<���<�ڃ<�	�<8�<��|<&y<�u<��q<1n<~�j<��f<e:c<V�_<�[<�GX<K�T<p Q<�^M<I�I<o!F<�B<��><�V;<�7<I24<E�0<k-<}�)<�&<��"<L<r�<�7<��<Yg<7<��
<�X<L
<�� <Y�;?��;�%�;���;f��;�F�;��;���;F��;J��;3�;�,�;|a�;ا�;���;xg�;M�;�l�;�	�;귊;x�;7I�;Yv;Al;�Lb;�yX;��N;:E;"�;;f~2;Q);�C ;oU;��;��;\��:���:��:�]�:x�:c��:��:ne�:��q:�S:��4:Y�:zU�9
��9�8{9N9ĳ7b��W�I��B���ӹ���ٳ��v:�� U��\o��Ä�������~���?���ĺ�Ѻ�޺��y���P��?��&�����+�:= ��I&�mR,�+W2�W8�8U>��ND�5FJ��;P�.V��\��b�!�g���m���s�1�y���͂������� �������쟑�Ę���ƍ���  �  �o=�=��=�O=��=�=.=�� =zk =�	 =BO�<J��<���<1��<�6�<�n�<l��<I��<#�<�C�<yv�<��<��<��<�4�<�`�<Y��<���<���<��<&�<qH�<�h�<���<��<���<���< ��<� �<d�<c!�<�-�<�7�<�>�<�B�<WD�<�B�<>�<N6�<K+�<��<E�< ��<Z��<��<���<)}�<�U�<�)�<i��<���<1��<iS�<|�<S��<��<Q:�<\��<*��<�:�<���<�z�<'�<}��<�:�<aǼ<P�<�Թ<.U�<�Ѷ<KJ�<���<�/�<���<��<l�<�Ϋ<.�<߉�<��<8�<���<rڡ<m'�<�q�<���<���<�A�<ς�<���<D��<79�<Tr�<ة�<�ߌ<Z�<�G�<�y�<���<�ڃ<�	�<!8�<��|<&y<�u<��q<1n<a�j<��f<J:c<S�_<�[<�GX<U�T<p Q<�^M<a�I<�!F<�B<��><|V;<��7<a24<'�0<n-<��)<n&<��"<\<�<�7<��<>g<E<��
<�X<^
<~� <R�;A��;�%�;���;���;�F�;��;���;1��;|��;�;`,�;|a�;���;���;�g�;P�;�l�;�	�;��;5x�;{I�;�Xv;Al;'Lb;yX;��N;�9E;Q�;;?~2;�P);�C ;�U;4�;�;��:>��:k��:�\�:u�:U��:S�:|e�:�q:�S:��4:��:OV�9#��9�;{9O9���7<r����I�FD��Eӹa��D��Nu:�� U�[\o���^��������~���?����ĺ��ѺE޺���������a�������@+�= �GJ&�_R,�W2��W8��T>�;OD��FJ��;P�G.V�B\�>b���g���m�f�s�Z�y�ʭ��̂�Å�t���V���ħ����֘��ْ��ō���  �  �o=�=��=�O=��=�=
.=�� =xk =�	 =9O�<P��<���<#��<�6�<�n�<q��<I��<�<�C�<wv�<���<��<
�<�4�<�`�<S��<r��<���<��<&�<gH�<�h�<���<#��<���<���<(��<� �<i�<d!�<�-�<�7�<�>�<�B�<ID�<�B�<>�<O6�<S+�<��<F�<��<c��<��<���<%}�<{U�<�)�<c��<���<+��<oS�<�<P��<���<C:�<]��<��<�:�<���<�z�<+�<n��<�:�<bǼ<#P�<�Թ<0U�<�Ѷ<?J�<���<�/�<���<��<vl�<�Ϋ<.�<���<��<(8�<���<pڡ<m'�<�q�<���<���<�A�<ł�<���<J��<.9�<Wr�<ө�<�ߌ<W�<�G�<�y�<���<�ڃ<�	�<"8�<��|<,&y<�u<��q< 1n<g�j<��f<R:c<_�_<
�[<�GX<j�T<X Q<�^M<:�I<�!F<�B<��><�V;<��7<|24<�0<o-<t�)<x&<��"<A<��<�7<��<=g<<<�
<�X<x
<r� <��;��;�%�;���;a��;�F�;��;��;��;|��;�;w,�;�a�;���;���;Yg�;d�;�l�;�	�;��;�w�;|I�;sXv;�Al;%Lb;�yX;��N;:9E;_�;;~2;Q);�C ;�U;�;��;���:Ӓ�:t��:�\�:��:~��:'�:�f�:L�q:�S:}�4:Z�:�U�9M��9�={9�G9C�7�q��7�I�'B���ӹ��ɵ�it:�1U�<\o�lÄ�����爵�q���>����ĺ �Ѻ@޺א����ȭ�/��t�����+�2= �J&��R,��V2��W8��T>�ROD�gFJ�Z;P��.V�?\��b���g��m��s�J�y�!���̂�Å�D���G�������⟑��������������  �  �o=�=��=�O=z�=�=.=�� =yk =�	 =6O�<R��<���<&��<�6�<�n�<l��<N��<�<�C�<yv�<��<��<��<|4�<�`�<O��<s��<��<��<&�<rH�<�h�<���<$��<���<��<$��<� �<h�<]!�<�-�<�7�<�>�<�B�<ND�<�B�<>�<N6�<D+�<��<B�<��<`��<��<���<,}�<}U�<�)�<`��<���<4��<dS�<{�<R��<��<F:�<e��<��<�:�<���<�z�<&�<}��<�:�<gǼ<P�<�Թ<7U�<�Ѷ<LJ�<���<�/�<��<��<rl�<�Ϋ<.�<މ�<��<8�<���<xڡ<e'�<�q�<���<���<�A�<Ȃ�<~��<K��<,9�<Yr�<֩�<�ߌ<`�<�G�<�y�<���<�ڃ<�	�<28�<��|<&y<�u<��q<1n<s�j<��f<]:c<e�_<�[<�GX<R�T<f Q<_M<;�I<�!F< �B<��><�V;<��7<P24<#�0<w-<m�)<~&<��"<F<��<�7<��<Gg</<��
<�X<Y
<�� <S�;��;&�;���;c��;.G�;��;���;2��;��;5�;z,�;ya�;���;���;�g�;^�;�l�;�	�;A��;�w�;�I�;�Xv;�@l;"Lb;wyX;n�N;�9E;>�;;�}2;Q);�C ;�U;K�;��;H��:���:��:]�:�:;��:G�:Xe�:��q:�S:��4:��:&Y�9���9�:{9VO9` �7m����I�.C��ӹC��,���u:��U�Zo�<Ä�6�!���t���?����ĺ��ѺV޺L�꺒������Z��l����}+�r= �J&��R,��V2��W8�*U>�OD��FJ��;P�+.V�E\��b�O�g���m�n�s�2�y����̂�������1�������ȟ��͘��ߒ��ۍ���  �  �o=�=��=�O=��=�=.=�� =xk =�	 =AO�<S��<���<*��<�6�<�n�<b��<S��<�<�C�<wv�<��<��<��<�4�<�`�<T��<|��< ��<��<&�<}H�<�h�<���<*��<���<	��<��<�<g�<c!�<�-�<�7�<�>�<�B�<ZD�<�B�<>�<Q6�<H+�<��<?�<#��<X��<��<���<&}�<~U�<�)�<n��<���<2��<fS�<}�<V��<��<T:�<[��<"��<�:�<���<�z�<(�<���<�:�<nǼ<P�<�Թ<6U�<�Ѷ<VJ�<���<�/�< ��<��<wl�<�Ϋ<.�<ቨ<��<8�<���<pڡ<h'�<�q�<}��<���<�A�<ʂ�<}��<I��<89�<Pr�<ԩ�<�ߌ<a�<�G�<�y�<���<�ڃ<�	�< 8�<��|<!&y<�u<��q<
1n<~�j<��f<h:c<M�_<%�[<�GX<\�T<e Q<�^M<Q�I<�!F<!�B<�><{V;<��7<U24<�0<e-<��)<&<��"<N<t�<�7<��<Og<:<�
<�X<V
<�� <L�;Y��;&�;���;���;�F�;��;���;^��;}��;�;�,�;�a�;ȧ�;���;�g�;[�;�l�;�	�;��;x�;tI�;�Xv;<Al;*Lb;�yX;��N;w9E;#�;;\~2;�P);�C ;�U;�;��;�:���:
��:�\�:>�:f��:|�:�e�:[�q:�S:��4:��:?V�9���9|;{9�T9�7/f����I��A��Eӹ���ڲ�}u:�� U�\o�����������i~���?��[�ĺ׉Ѻg޺А�s���q�����U����h+�v= � J&�TR,�&W2��W8�U>��ND��FJ�V;P�.V�h\�{b���g���m�H�s�
�y����	͂���r������ϧ����������˒��ݍ���  �  �o=�=��=�O=��=�=	.=�� =xk =�	 =8O�<O��<���<$��<�6�<�n�<l��<I��<�<�C�<zv�<��<��<��<�4�<�`�<T��<z��<���<��<&�<qH�<�h�<���<*��<���<��<$��<� �<f�<l!�<�-�<�7�<�>�<�B�<KD�<�B�<>�<O6�<W+�<��<?�<��<\��<��<��<}�<xU�<�)�<d��<���<*��<sS�<��<O��<���<F:�<V��<��<�:�<���<�z�<'�<z��<�:�<mǼ<%P�<�Թ<6U�<�Ѷ<JJ�<���<�/�<���<��<vl�<�Ϋ<.�<牨<��<&8�<���<kڡ<h'�<�q�<���<���<�A�<Ă�<���<G��<-9�<Lr�<Щ�<�ߌ<W�<�G�<�y�<���<�ڃ<�	�< 8�<��|<2&y<�u<��q<1n<v�j<��f<a:c<[�_<"�[<�GX<o�T<i Q<�^M<N�I<�!F<��B<
�><|V;<��7<~24<�0<[-<q�)<u&<��"<B<g�<�7<��<;g<4<�
<�X<t
<p� <]�;?��;�%�;���;���;�F�;��;��;.��;���;�;�,�;�a�;���;���;�g�;V�;�l�;�	�;��;x�;gI�;�Xv;�Al;�Kb;~yX;��N;39E;!�;;~2;�P);�C ;dU;��;��;'��:ڒ�:���:n\�:�:���:
�:Yf�:��q:�S:�4:��:$V�9Ϯ�9R;{9�M9��7�g����I��@��Iӹ���j���t:�� U�]\o�Ä�����6�����a?����ĺ%�Ѻ޺+��u������W�������+�== �-J&��R,�CW2��W8�{T>�VOD��FJ�:;P��.V�L\��b���g���m��s�G�y�����̂���H���*�����������Ԙ������Ս���  �  �o=�=��=�O=}�=�=	.=�� =uk =�	 =1O�<I��<���<��<�6�<�n�<n��<A��<�<�C�<qv�<��<��<��<4�<�`�<W��<s��<��<��<&�<sH�<�h�<���<&��<���<��<*��<� �<n�<b!�<�-�<�7�<�>�<�B�<JD�<�B�<>�<J6�<F+�<��<H�<
��<_��<���<���<)}�<tU�<�)�<T��<���<*��<dS�<x�<O��<��<C:�<j��<��<�:�<���<�z�</�<}��<�:�<kǼ<P�<�Թ<:U�<�Ѷ<LJ�<���<�/�<��<��<xl�<�Ϋ<.�<䉨<��<8�<���<rڡ<h'�<�q�<���<���<�A�<�<}��<D��<$9�<Yr�<ͩ�<�ߌ<W�<�G�<�y�<���<�ڃ<�	�<28�<��|<%&y<�u<��q<(1n<r�j<��f<[:c<k�_<�[<�GX<e�T<c Q<_M<>�I<�!F<�B<��><�V;<��7<W24<�0<t-<c�)<i&<��"<8<��<�7<��<+g</<�
<�X<X
<p� <\�;��;&�;���;a��;%G�;��;��;2��;���;7�;�,�;�a�;���;��;�g�;t�;�l�;�	�;B��;�w�;�I�;vXv;"Al;Lb;[yX;v�N;'9E;g�;;�}2;�P);\C ;�U;6�;h�;]��:���:k��:p\�:�:
��:	�:�e�:M�q:JS:��4:��:>X�9]��9�>{9O9��7'i���I��A��sӹ���8���t:��U�]Zo�:Ä������������?����ĺ��Ѻ�޺���p�����=��������+�u= �CJ&��R,��V2��W8�U>�SOD��FJ��;P�.V��\��b�J�g���m�9�s��y����̂���Y���6���������Ę������ፚ��  �  �o=�=��=�O=��=�=.=�� ={k =�	 =6O�<N��<���<��<�6�<�n�<f��<L��<�<�C�<zv�<��<$��<��<�4�<�`�<R��<v��<��<��<&�<{H�<�h�<���</��<���<��<#��<� �<m�<e!�<�-�<�7�<�>�<�B�<VD�<�B�<>�<Q6�<F+�<��<A�<��<\��<���<��<}�<sU�<�)�<c��<���<0��<fS�<|�<^��<��<R:�<Y��<��<�:�<���<�z�<.�<���<�:�<zǼ<"P�<�Թ<CU�<�Ѷ<TJ�<���<�/�<��<��<wl�<�Ϋ<.�<䉨<��<8�<���<pڡ<c'�<�q�<���<���<�A�<���<y��<F��<-9�<Or�<ܩ�<�ߌ<g�<�G�<�y�<���<�ڃ<�	�<%8�<��|<+&y<�u<��q<!1n<��j<��f<v:c<g�_<�[<�GX<e�T<k Q<�^M<D�I<�!F<�B<��><�V;<��7<V24<,�0<_-<m�)<t&<��"<0<q�<�7<��<Bg<(<�
<�X<U
<�� <[�;A��;�%�;���;n��;�F�;��;��;T��;p��;O�;�,�;�a�;���;���;�g�;q�;�l�;�	�;��;x�;iI�;�Xv;7Al;mLb;�yX;t�N;{9E;2�;;~2;�P);RC ;JU;Ӆ;d�;��:Ӓ�:��:�\�:5�:N��:��:�e�:�q:)S:2�4:��:W�9̭�9;>{9�Q9���7)Z��t�I��@��;ӹ���4���t:�� U�v[o�$Ä����������~���?����ĺ�Ѻ<޺ݐ��������������	��+��= �4J&��R,�2W2�~W8�U>��ND�pFJ�p;P�I.V�^\��b���g���m� �s���y����̂���\�����������՟����������э���  �  �o=�=��=�O=��=ߎ=.=�� ={k =�	 =;O�<C��<���<(��<�6�<�n�<`��<E��<�<�C�<yv�<٧�<��<��<�4�<�`�<a��<���<���<��<&�<zH�<�h�<���<&��<���<��<'��<
�<g�<r!�<�-�<�7�<�>�<�B�<YD�<�B�<
>�<B6�<A+�<��<8�<��<N��<	��<���<}�<�U�<�)�<b��<���<,��<bS�<o�<N��<��<W:�<W��<7��<�:�<���<�z�<(�<���<�:�<tǼ<P�<�Թ<=U�<�Ѷ<WJ�<���<�/�<���<��<�l�<�Ϋ<.�<҉�<��<8�<���<jڡ<d'�<�q�<w��<���<�A�<Ƃ�<���<:��<29�<Er�<ک�<�ߌ<Z�<�G�<�y�<���<�ڃ<�	�<8�<��|<1&y<�u<��q<$1n<��j<��f<h:c<f�_<-�[<�GX<f�T<� Q<�^M<l�I<�!F<�B<�><]V;<��7<I24<+�0<R-<w�)<^&<��"<I<i�<�7<��<4g<1<ڬ
<�X<A
<}� <�;_��;�%�;��;���;�F�;�;���;P��;���;9�;�,�;�a�;ߧ�;���;�g�;Y�;m�;�	�;��;gx�;gI�;�Xv;�@l;�Kb;yX;P�N;f9E;��;;~2;oP);�C ;rU;�;��;<��:Ē�:���:�\�:��:|��:��:�d�:��q:�S:�4:��:�W�9\��95;{9�V9,�7�`����I��B���ӹ������u:���T�.\o����������;~���@����ĺ��Ѻ`޺<�꺨��������9����+�W= ��J&��R,�W2��W8�AU>�;OD�GJ�y;P�T.V�?\��b��g�o�m��s�"�y�~���̂���w���������������������������  �  �o=�=��=�O=��=�=.=�� =uk =�	 =;O�<H��<���<��<�6�<�n�<l��<A��<!�<�C�<rv�<��<��< �<�4�<�`�<Q��<k��<��<��<&�<qH�<�h�<���<.��<���<��<.��<� �<n�<e!�<�-�<�7�<�>�<�B�<RD�<�B�<>�<Q6�<F+�<��<D�<��<X��<���<��<}�<vU�<�)�<]��<���<*��<eS�<}�<^��<���<M:�<Y��<��<�:�<���<�z�</�<y��<�:�<nǼ</P�<�Թ<<U�<�Ѷ<JJ�<���<�/�<��<z�<tl�<�Ϋ<.�<艨<��<8�<���<mڡ<o'�<�q�<���<���<�A�<���<���<B��<.9�<Qr�<Ω�<�ߌ<a�<�G�<�y�<���<�ڃ<�	�<!8�<��|<,&y<�u<��q<,1n<w�j<��f<f:c<j�_<�[<�GX<l�T<j Q<�^M<5�I<�!F<�B<	�><�V;<��7<V24<�0<e-<w�)<g&<��"<&<h�<�7<��<,g<?<�
<�X<U
<�� <l�;I��;�%�;���;@��;�F�;��;��;*��;���;;�;�,�;�a�;���;��;vg�;u�;�l�;�	�;���;�w�;mI�;�Xv;kAl;lLb;�yX;v�N;89E;H�;;�}2;�P);uC ;U;��;v�;��:o��:k��:r\�:"�:\��:��:(f�:��q: S:S�4:��:FW�9v��9�>{99M9�)�7�f���I�.?���ӹ?��q��bt:�� U��[o��Ä� ������~��J?���ĺ�Ѻ�޺������	��R������,�[= �YJ&��R,�$W2��W8�U>�OD�oFJ�J;P�j.V�P\��b���g���m� �s�	�y�׭��̂�����������������Ø������Ӎ���  �  �p=l=б=�Q=��=��=�0=� =�n =j =,W�<ߒ�<���<��<MA�<�y�<0��<���<2�<�Q�<���<(��<��<��<F�<s�<���<|��<���<��<�<�<�_�<m��<���<j��<���<>��<h
�<(�<�1�<�A�<�N�<�Y�<�a�<3g�<}i�<�h�<4e�<`^�<_T�<�F�<)6�<�!�<	
�<n��<<��<-��<��<OZ�<B+�<V��<+��<��<KF�<r�<Z��<�m�<$�<���<Pn�<[�<��<kG�<Tܿ<m�<l��<���<��<r��<<�<�x�<��<�\�<�Ȱ<w1�<\��<���<�U�<Q��<��<\�<e��<���<wG�<_��<�֜<��<�\�<⛗<2ٕ<��<�M�<���<Ȼ�<R��<Z#�<1U�<ʅ�<P��<��<|�<p>�<j�|<�,y<��u<��q<=/n<��j<��f<�/c<Ӆ_<��[<64X<�T<�P<�BM<!�I<��E<+aB<�><�+;<+�7<�4<�q0<&�,<E\)<�%<�V"<��<Rc<i�<�<�<3�<M[
<t<Գ<wi <�K�;��;�f�;�	�;��;�{�;�K�;%,�;��;��;�-�;IO�;E��;�ƪ;��;���;���;���;$�;]҉;m��;��~;3�t;�zj;g�`;ȸV;$M;ԀC;�:;��0;8�';A�;�;e�;!E;^r�:ؐ�:J��:${�:�A�:};�:2h�:ǅ:��l:�%N:d�/:�:�5�9Ѯ9
j9�E�8m��6.�Ӹ��X������#ڹB"�j�"���=��X��Ir��+�����d���c����q��^ƺ3�Һi!ߺZ�뺧����"��D�xb�Fx�p��� ���&���,��2�ȝ8�D�>�r�D�J��oP��]V�J\�6b��h��n���s���y����Ԃ�pȅ����ֱ������C���V������v����  �  �p=r=Ǳ=�Q=��=��=�0=� =�n =i =9W�<ْ�<���<��<4A�<�y�<%��<���<8�<�Q�<���< ��<��<��<F�<�r�<~��<���<���<��<�<�<�_�<c��<��<���<���<I��<Z
�<*�<�1�<�A�<O�<�Y�<�a�<g�<}i�<�h�<De�<k^�<UT�<�F�<,6�<�!�<�	�<p��<&��<��<#��<AZ�<U+�<Y��<%��<ۅ�<OF�<��<`��<�m�<�<���<Un�<_�<��<XG�<Xܿ<m�<t��<���<��<n��</�<�x�<��<�\�<�Ȱ<|1�<T��<���<�U�<X��<��<\�<a��<���<{G�<i��<�֜<��<n\�<ٛ�<1ٕ<��<N�<���<���<F��<n#�<<U�<΅�<G��<��<��<x>�<{�|<�,y<��u<��q<"/n<��j<
�f<�/c<��_<��[<64X< �T<,�P<�BM<8�I<��E<aB<)�><�+;<R�7<�4<�q0<&�,<_\)<s�%<�V"<��< c<w�<�<�<>�<K[
<r<ĳ<�i <�K�;<��;zf�;Z	�;��;�{�;�K�;�+�;��;\�;�-�;�O�;���;�ƪ;|�;˃�;���;|��;$�;x҉;���;��~;5�t;{j;�`;&�V;�M;��C;�:;k�0;Ƨ';N�;^�;��;HE;~q�:��:u��:�z�:TA�:�;�:Yi�:�ǅ:��l:�"N:~�/:I:�6�9�Ю9�
j9PJ�8��6��Ӹ�X�[����$ڹ�#���"��=��X��Hr�*+��t������뽬�;q��Gƺ��Һ�!ߺ���o���w"�3E�;b�y����� ��&�6�,��2��8���>�ԋD��~J�ioP�6^V��J\��5b�uh�{n�
�s���y����EԂ�+ȅ�����}���&���K���U���Q���M����  �  �p=u=Ǳ=�Q=��=|�=�0=
� =�n =e =8W�<֒�<���<��<5A�<�y�<��<���</�<�Q�<��<��<��<��<!F�<s�<���<���<���<��<�<�<`�<g��<��<t��<���<C��<S
�<;�<�1�<�A�<�N�<�Y�<�a�<g�<�i�<�h�<8e�<i^�<_T�<�F�<6�<�!�<�	�<���<6��<!��<7��<2Z�<Z+�<K��<4��<��<LF�<{�<T��<�m�<	�<���<Mn�<X�<��<SG�<iܿ<�l�<q��<���<��<o��</�<y�<��<�\�<�Ȱ<x1�<^��<���<�U�<G��<��<
\�<q��<���<oG�<r��<�֜<��<r\�<뛗<:ٕ<��<	N�<���<ϻ�<H��<j#�<+U�<υ�<V��<��<��<k>�<x�|<�,y<��u<��q</n<��j<��f<�/c<��_<��[<B4X<�T<,�P<�BM<A�I<��E<*aB<1�><�+;<J�7<�4<�q0<�,<]\)<m�%<�V"<��<#c<��<�<�<,�<K[
<�<��<�i <�K�;c��;�f�;u	�;��;�{�;L�;�+�;7�;m�;�-�;rO�;,��;�ƪ;`�;��;���;���;�#�;S҉;���;��~;��t;�zj;��`;�V;,M;�C;=:;��0;Z�';٠;۸;�;�E;�p�:g��:���:�{�:GB�:�;�:�h�:�ƅ:'�l:W"N:��/:R:�4�9	Ү9Yj9G[�8`�6��Ӹ`�X�َ���$ڹ�#���"�,�=�!X��Ir�l+���������F���Er���ƺڢҺ� ߺ1��#���3"��E�za��x�*��ϖ �.�&�%�,�:�2���8���>��D�6J�coP��]V��J\�h5b��h��n��s���y�H��QԂ�Mȅ�$�������,���,���=���m���J����  �  �p=n=ɱ=�Q=��=��=�0=� =�n =g =8W�<��<���<��<1A�<�y�<!��<���<1�<�Q�<���<"��<��<��<F�<s�<���<y��<���<��<�<�<�_�<_��<��<z��<���<K��<Q
�<+�<�1�<�A�<�N�<�Y�<�a�<g�<i�<�h�<Ce�<i^�<WT�<�F�< 6�<�!�< 
�<r��<-��<��<%��<BZ�<Z+�<N��<4��<ޅ�<PF�<��<Z��<�m�<�<���<Mn�<Y�<��<YG�<Xܿ<�l�<v��<���<��<t��<)�<�x�<��<�\�<�Ȱ<q1�<Z��<���<�U�<P��<��<\�<a��<���<rG�<v��<�֜<��<l\�<ݛ�<2ٕ<��<N�<���<˻�<G��<i#�<7U�<˅�<N��<��<�<n>�<l�|<�,y<��u<��q<"/n<��j<��f<�/c<��_<��[<24X<�T<�P<�BM<&�I<��E< aB<&�><�+;<L�7<�4<�q0<�,<^\)<��%<�V"<��<c<|�<��<�<0�<U[
<u<ɳ<�i <�K�;3��;�f�;r	�;���;�{�;�K�;�+�;��;L�;�-�;�O�;���;�ƪ;[�;΃�;���;���;�#�;]҉;x��;��~;G�t;�zj;ۈ`;�V;�M;�C;K:;~�0;�';]�;��;��;ZE;�q�:`��:���:�{�:�A�:�;�:Xi�:%ǅ:(�l:�"N:B�/:Q:<5�9�Ѯ9nj91J�8�-�6L�Ӹ��X�����7#ڹ}$���"�؝=�X��Ir��+�������=����q��$ƺV�Һ�!ߺ������"�KE�#b�#y����� ���&�8�,�(�2���8���>���D��~J��oP��]V��J\��5b��h��n���s��y����DԂ�;ȅ������������`���]���B���j����  �  �p=k=̱=�Q=��=��=�0=� =�n =p =-W�<ߒ�<���<��<EA�<�y�<,��<���<.�<�Q�<��<*��<��<��<F�<s�<���<y��<���<��<�<�<�_�<k��<��<l��<���<4��<Z
�<+�<�1�<�A�<�N�<�Y�<�a�<-g�<|i�<�h�<9e�<k^�<VT�<�F�<26�<�!�<
�<s��<9��<)��<(��<JZ�<L+�<[��<4��<؅�<UF�<x�<a��<�m�<�<���<Wn�<Z�<��<^G�<Xܿ<m�<b��<���<��<b��<4�<�x�<��<�\�<�Ȱ<v1�<U��<���<�U�<Y��<��<\�<Z��<���<tG�<e��<�֜<��<�\�<盗<6ٕ<��<�M�<�<���<M��<h#�<6U�<υ�<M��<��<z�<}>�<]�|<�,y<��u<��q</n<q�j<��f<�/c<��_<��[<74X<�T<�P<�BM<�I<��E<!aB<(�><�+;<C�7<�4<�q0<A�,<H\)<�%<�V"<��<Dc<��<�<�<,�<n[
<g<ٳ<�i <�K�;4��;�f�;s	�;���;�{�;�K�;�+�;��;|�;d-�;UO�;u��;�ƪ;}�;у�;���;k��;�#�;�҉;c��;_�~;,�t;{j;��`;'�V;�M;��C;�:;�0;�';j�;��;B�;qE;r�:���:���:�{�:$A�:<�:�h�:�ǅ:�l:�$N:��/:�:�5�9Qή9�j9yJ�8X��6��Ӹ��X������'ڹ#���"��=�rX�DHr��+��O������B���0q��ƺ�Һ"ߺf�������"��D��a�~x�E��� ���&���,���2���8�f�>��D��~J�coP�^V�HJ\�"6b�Ph��n���s���y����JԂ��ȅ�ļ��ޱ��/���?���U���;��������  �  �p=m=ɱ=�Q=��=�=�0=� =�n =o =6W�<��<���<��<4A�<�y�<$��<���<3�<�Q�<���<+��<��<��<F�<s�<���<x��<���<��<�<�<�_�<i��<��<t��<���<=��<\
�<(�<�1�<�A�<�N�<�Y�<�a�<%g�<�i�<�h�<2e�<l^�<\T�<�F�<-6�<�!�<
�<z��<5��<!��<.��<DZ�<Z+�<V��<2��<���<VF�<q�<f��<�m�<�<���<Ln�<W�<��<XG�<Uܿ<m�<i��<���<��<g��<3�<�x�<��<�\�<�Ȱ<s1�<X��<���<�U�<Z��<��<\�<f��<���<vG�<t��<�֜<��<r\�<⛗<7ٕ<��<N�<���<ƻ�<U��<g#�<+U�<ׅ�<P��<��<��<m>�<j�|<�,y<w�u<��q<$/n<��j<��f<�/c<��_<��[<4X<�T<�P<�BM<"�I<��E<#aB<7�><�+;<@�7<�4<�q0<;�,<Y\)<��%<�V"<��<!c<��<�<�<5�<^[
<z<ڳ<~i <�K�;Z��;�f�;w	�;���;�{�;�K�;�+�;��;v�;t-�;wO�;X��;�ƪ;��;ƃ�;���;���;�#�;R҉;v��;"�~;V�t;S{j;V�`;.�V;M;�C;�:;~�0;��';��;Ҹ;�;�E;�q�:c��:O��:�{�:�A�:,<�:'h�:�ǅ:ƪl:$N:�/:D:�4�9�Ѯ9j9fH�8���6d�Ӹ&�X�����c&ڹG#���"�ם=�|X��Ir��+�� ���������q��aƺ�ҺO!ߺ͐뺯���#"�9E��a��x�q��� ���&�D�,���2�՝8�,�>��D�/J�#oP��]V��J\��5b��h��n���s�8�y����AԂ�]ȅ���������(���R�������H���g����  �  �p=u=Ǳ=�Q=��=��=�0=� =�n =k =6W�<��<���<��<9A�<�y�<��<���<2�<�Q�<���<#��<$��<��<F�<�r�<���<���<���<��<�<�<�_�<_��<��<r��<���<C��<J
�<*�<�1�<�A�<�N�<�Y�<�a�< g�<ti�<�h�<Ce�<q^�<RT�<�F�<'6�<�!�<�	�<}��<9��<#��<5��<=Z�<_+�<P��<7��<څ�<UF�<��<[��<�m�<�<���<Kn�<Q�<��<OG�<Xܿ<�l�<m��<���<��<e��<&�<�x�<��<�\�<�Ȱ<x1�<\��<���<�U�<T��<��<\�<c��<���<tG�<w��<�֜<��<u\�<<4ٕ<��<N�<���<λ�<I��<r#�<7U�<Ņ�<F��<��<��<i>�<h�|<�,y<{�u<��q</n<��j<��f<�/c<��_<��[<(4X<��T<�P<�BM<A�I<��E<aB<�><�+;<a�7<�4<�q0<.�,<Z\)<��%<�V"<��<-c<��<��<�<4�<_[
<~<̳<�i <�K�;��;~f�;w	�;��;�{�;�K�;�+�;��;N�;W-�;oO�;P��;�ƪ;@�;̓�;���;x��;�#�;N҉;���;��~;�t;�zj;�`;U�V;�M;(�C;~:;��0;Ƨ';��;��;�;�E;Dq�:���:���:�{�:FA�:$<�:_i�:>ǅ:�l:9#N:1�/:1:e3�9�Ϯ9�j9�K�8l��6�Ӹ�X� ����&ڹ�$��"��=�#X��Jr�\+���������ᾬ�wq���ƺL�Һt!ߺ�������	"�iE�ha��x����� ���&�?�,�ޡ2���8���>���D��~J��oP�<^V��J\�o5b��h��n�$�s�)�y�����Ԃ�=ȅ���������`���Z���q���d���l����  �  �p=l=Ʊ=�Q=��=��=�0=� =�n =o =2W�<��<���<��<;A�<�y�<0��<���<2�<�Q�<���<&��<��<��<F�<s�<w��<w��<���<��<�<�<�_�<d��<��<h��<���<8��<P
�<&�<�1�<�A�<�N�<�Y�<�a�<(g�<�i�<�h�<=e�<m^�<[T�<G�<06�<�!�<
�<}��<:��<#��<2��<LZ�<[+�<Z��<>��<��<TF�<|�<b��<�m�<�<���<Nn�<V�<��<TG�<Sܿ<�l�<e��<���<��<c��<,�<�x�<��<�\�<�Ȱ<q1�<K��<���<�U�<Y��<��<\�<e��<���<xG�<u��<�֜<��<x\�<<=ٕ<��<N�<���<ѻ�<N��<g#�<8U�<̅�<X��<��<z�<p>�<_�|<�,y<|�u<��q</n<z�j<��f<�/c<��_<��[<'4X< �T<�P<�BM<�I<��E<5aB<#�><�+;<D�7<�4<�q0<<�,<Q\)<��%<�V"<��<0c<��<�<�<5�<q[
<�<ҳ<�i <�K�;@��;�f�;B	�;��;�{�;�K�;�+�;��;b�;^-�;HO�;I��;�ƪ;X�;���;���;m��;�#�;c҉;J��;9�~;|�t;%{j;��`;:�V;M;\�C;�:;s�0;2�';��;��;�;�E;8r�:u��:���:`|�:�A�:<�:�h�:�ǅ:�l:r$N:��/::�4�9�ή9^	j9�E�8�G�6��Ӹ��X�o���B'ڹ$�W�"��=�X�dIr��+������������*q���ƺ8�ҺZ!ߺ�뺓���"��D��a��x����� �h�&�g�,���2��8�^�>�
�D��~J��oP��]V��J\�6b��h��n��s�$�y����pԂ�~ȅ����ձ��R���]���r���Q��������  �  �p=m=ɱ=�Q=��=��=�0=� =�n =q ==W�<��<���<��<FA�<�y�<-��<���<;�<�Q�<���<7��<��<��<F�<s�<���<x��<���<��<�<�<�_�<`��<��<n��<���<3��<Y
�<�<�1�<�A�<�N�<�Y�<�a�<%g�<|i�<�h�<:e�<r^�<eT�<�F�<66�<�!�<

�<w��<9��<&��<+��<MZ�<]+�<`��<0��<��<]F�<y�<g��<�m�<�<���<Mn�<L�<��<WG�<Dܿ<m�<^��<���<��<\��<,�<�x�<��<�\�<�Ȱ<p1�<T��<���<�U�<`��<��<"\�<d��<���<~G�<x��<�֜<��<�\�<囗<:ٕ<��<
N�<Ņ�<»�<^��<g#�<9U�<υ�<O��<��<|�<o>�<O�|<�,y<q�u<q�q</n<w�j<��f<�/c<��_<o�[<4X<	�T< �P<�BM< �I<��E<&aB<$�><�+;<>�7<�4<�q0<E�,<h\)<��%<�V"<��<Fc<��<�<�<G�<i[
<x<��<�i <L�;.��;�f�;m	�;���;�{�;�K�;�+�;��;R�;S-�;^O�;}��;�ƪ;|�;���;���;���;�#�;d҉;d��;$�~;8�t;D{j;��`;^�V;]M;��C; :;��0;C�';��;��;4�;�E;Fr�:���:���:}{�:B�:�<�:�h�:�ǅ:�l:�#N:r�/:n:I2�9�Ϯ9)j9�7�8��6ҰӸ��X�;����(ڹ�#���"���=�-X�Jr��+��`�� ���i����p��ƺB�Һe!ߺ���6����!��D��a��x�U��ɖ �U�&��,�x�2��8�ߕ>�	�D��~J�goP��]V��J\�6b��h�-	n���s�Q�y���PԂ��ȅ�ʼ��ɱ��<�����������?��������  �  �p=p=ȱ=�Q=��=��=�0=� =�n =p =<W�<��<���<��<HA�<�y�<-��<���<7�<�Q�< ��<(��<��<��<F�<s�<���<x��<���<��<�<�<�_�<b��<ݠ�<c��<���<.��<N
�<)�<�1�<�A�<�N�<�Y�<�a�<g�<~i�<�h�<?e�<j^�<\T�<�F�<06�<�!�<�	�<���<C��<.��<?��<AZ�<^+�<Z��<=��<��<SF�<~�<Y��<�m�<�<���<Hn�<S�<��<LG�<Sܿ<�l�<Z��<���<�<Z��<*�<�x�<��<�\�<�Ȱ<o1�<Z��<���<�U�<R��<��<\�<g��<���<zG�<w��<�֜<��<�\�<���<Eٕ<��<N�<���<˻�<Q��<j#�<8U�<˅�<P��<��<��<h>�<_�|<�,y<{�u<��q</n<g�j<��f<}/c<��_<��[<+4X<�T<�P<�BM<-�I<��E<%aB<!�><�+;<H�7<�4<�q0<?�,<f\)<��%<�V"<��<Kc<��<�<�<?�<r[
<�<׳<�i <�K�;8��;�f�;w	�;���;�{�;�K�;�+�;��;^�;I-�;5O�;0��;�ƪ;R�;˃�;���;l��;�#�;L҉;���;��~;C�t;�zj;Ĉ`;&�V;M;>�C;�:;��0;�';)�;H�;p�;/F;�q�:���:���:N|�:�A�:<�: i�: ǅ:0�l:�"N:�/:�:#4�9Ϯ9�j9�F�8//�6q�ӸW Y�[���S)ڹA$�E�"��=��X�EJr��+�����q���!����q���ƺ�Һ7!ߺ*��m���"� E�9a�gx�݉�v� ���&��,���2���8�J�>��D��~J��oP��]V��J\��5b��h��n�Q�s�*�y����~Ԃ��ȅ����󱋻b���X���k�������{����  �  �p=o=��=�Q=��=��=�0=� =�n =j =FW�<��<���<��</A�<�y�<+��<���<9�<�Q�<��<%��<&��<��<F�<s�<y��<y��<���<��<�<�<�_�<O��<��<o��<���<B��<D
�<&�<�1�<�A�<O�<�Y�<�a�<g�<�i�<�h�<Ee�<o^�<ZT�<G�<%6�<�!�<
�<���<7��<��<:��<EZ�<o+�<Q��<@��<߅�<UF�<��<T��<�m�<�<���<An�<a�<��<IG�<Rܿ<�l�<m��<���<��<i��<�<�x�<��<�\�<�Ȱ<o1�<O��<���<�U�<L��<��<\�<j��<���<yG�<���<�֜<��<k\�<<@ٕ<��<N�<���<ֻ�<M��<t#�<7U�<˅�<Y��<��<��<a>�<y�|<�,y<v�u<r�q</n<��j<��f<�/c<��_<e�[<'4X<ߌT<'�P<�BM<*�I<u�E<3aB<(�><�+;<a�7<�4<�q0<)�,<{\)<��%<�V"<��<c<��<�<<D�<f[
<�<ѳ<�i <�K�;\��;�f�;J	�;���;�{�;�K�;�+�;��;�;r-�;fO�;E��;�ƪ;)�;���;���;]��;%$�;.҉;z��;��~;��t;�zj;��`;L�V;M;q�C;w:;1�0;�';�;�;��;F;�q�:���:��:x|�:�A�:)<�:�i�:�ƅ:-�l:"N:�/::|7�9�ή9)j95F�8H�6[�Ӹ��X�ʏ���%ڹ�&���"�!�=��X��Ir��+���������V����q���ƺ1�Һ!ߺM�뺀����!�E�ta�*y����� �d�&���,��2�O�8�j�>���D��~J��oP��]V�K\��5b�0 h��n�t�s�<�y����Ԃ�Yȅ�
�������]�������r�������U����  �  �p=q=ʱ=�Q=��=��=�0=� =�n =n =>W�<��<���<�<NA�<�y�</��<���<9�<�Q�<��<2��<��<��<F�<s�<���<}��<���<��<�<�<�_�<U��<۠�<^��<���<*��<Q
�<�<�1�<�A�<�N�<�Y�<�a�<#g�<�i�<�h�<;e�<u^�<dT�<G�</6�<�!�<
�<���<L��<7��<<��<IZ�<^+�<Y��<;��<��<[F�<~�<U��<�m�<�<���<En�<P�<���<VG�<Kܿ<�l�<W��<��<y�<Y��<"�<�x�<��<�\�<�Ȱ<r1�<\��<���<�U�<O��<��<\�<o��<���<xG�<v��<�֜<��<�\�<���<Bٕ<��<N�<���<Ի�<Y��<r#�<3U�<Ņ�<Q��<��<��<f>�<Y�|<�,y<��u<k�q</n<c�j<��f<z/c<��_<g�[</4X<�T<�P<�BM<2�I<��E<'aB<�><�+;<Y�7<�4<�q0<8�,<i\)<��%<�V"<��<Wc<��<�<�<C�<g[
<�<�<�i <�K�;��;�f�;�	�;��;�{�;�K�;�+�;��;*�;C-�; O�;+��;vƪ;^�;���;���;>��;�#�;?҉;���;�~;h�t;�zj;��`;x�V;VM;P�C;�:;��0;�';��;��;��;F;r�:���:���:-|�:7B�:�<�:	i�:�ƅ:��l:�#N:�/:k:s3�9rˮ9�
j9K?�8�)�69�Ӹ*Y���)ڹH%�r�"���=�cX��Jr��+�����H���m����q��Pƺ��Һ� ߺ��뺇���"��D�=a�:x������ ���&��,���2�i�8��>���D��~J��oP��]V�|J\��5b� h�	n�`�s���y�*��iԂ��ȅ��������T�������c���x��������  �  �p=g=Ʊ=�Q=��=��=�0=� =�n =u =;W�<��<���<��<6A�<�y�<=��<���<A�<�Q�<��<)��<��<��<F�<s�<|��<j��<���<��<�<�<�_�<b��<۠�<k��<���<#��<_
�<�<�1�<�A�<�N�<�Y�<�a�<g�<{i�<�h�<Ae�<p^�<]T�<�F�<A6�<�!�<
�<���<2��<��<5��<VZ�<Y+�<k��<9��<��<VF�<�<n��<�m�<�<���<Dn�<X�<���<TG�<9ܿ<m�<Q��<���<��<X��<0�<�x�<��<�\�<�Ȱ<c1�<N��<���<�U�<g��<��<\�<j��<���<�G�<t��<�֜<��<r\�<㛗<Kٕ<��<N�<υ�<ǻ�<R��<j#�<@U�<օ�<J��<��<v�<n>�<\�|<�,y<x�u<f�q</n<X�j<�f<w/c<��_<l�[<4X<�T<�P<�BM<�I<��E<aB<0�><�+;<D�7<�4<�q0<V�,<e\)<��%<W"<��<'c<��<4�<�<S�<y[
<�<ٳ<�i <0L�;8��;�f�;W	�;º�;�{�;�K�;�+�;��;[�;D-�;TO�;���;\ƪ;��;d��;���;L��;�#�;P҉;Q��;��~;0�t;�{j;׈`;O�V;M;�C;V:;z�0;��';��;Ÿ;��;�E;�r�:`��:���:|�:�A�:B<�: i�:vȅ:��l:�"N:��/:O:�5�9�̮9�	j9)-�8�6b�Ӹ��X�����)ڹ�#���"�Ӟ=�ZX�FIr��,�����h���G���>p���ƺ�Һ!ߺ!�뺣���"�yD��a��x�d��A� �N�&�.�,�*�2�̝8�C�>��D��~J�+oP�^V��J\�>6b��h��n�`�s�5�y�@��JԂ��ȅ���������D�����������x��������  �  �p=q=ʱ=�Q=��=��=�0=� =�n =n =>W�<��<���<�<NA�<�y�</��<���<9�<�Q�<��<2��<��<��<F�<s�<���<}��<���<��<�<�<�_�<U��<۠�<^��<���<*��<Q
�<�<�1�<�A�<�N�<�Y�<�a�<#g�<�i�<�h�<;e�<u^�<dT�<G�</6�<�!�<
�<���<L��<7��<<��<IZ�<^+�<Y��<;��<��<[F�<~�<U��<�m�<�<���<En�<P�<���<VG�<Kܿ<�l�<W��<��<y�<Y��<"�<�x�<��<�\�<�Ȱ<r1�<\��<���<�U�<O��<��<\�<o��<���<xG�<v��<�֜<��<�\�<���<Bٕ<��<N�<���<Ի�<Y��<r#�<3U�<Ņ�<Q��<��<��<f>�<Y�|<�,y<��u<k�q</n<c�j<��f<z/c<��_<g�[</4X<�T<�P<�BM<2�I<��E<'aB<�><�+;<Y�7<�4<�q0<8�,<i\)<��%<�V"<��<Wc<��<�<�<C�<g[
<�<�<�i <�K�;��;�f�;�	�;��;�{�;�K�;�+�;��;*�;C-�; O�;+��;vƪ;^�;���;���;>��;�#�;?҉;���;�~;h�t;�zj;��`;x�V;VM;P�C;�:;��0;�';��;��;��;F;r�:���:���:-|�:7B�:�<�:	i�:�ƅ:��l:�#N:�/:k:s3�9rˮ9�
j9K?�8�)�69�Ӹ*Y���)ڹH%�r�"���=�cX��Jr��+�����H���m����q��Pƺ��Һ� ߺ��뺇���"��D�=a�:x������ ���&��,���2�i�8��>���D��~J��oP��]V�|J\��5b� h�	n�`�s���y�*��iԂ��ȅ��������T�������c���x��������  �  �p=o=��=�Q=��=��=�0=� =�n =j =FW�<��<���<��</A�<�y�<+��<���<9�<�Q�<��<%��<&��<��<F�<s�<y��<y��<���<��<�<�<�_�<O��<��<o��<���<B��<D
�<&�<�1�<�A�<O�<�Y�<�a�<g�<�i�<�h�<Ee�<o^�<ZT�<G�<%6�<�!�<
�<���<7��<��<:��<EZ�<o+�<Q��<@��<߅�<UF�<��<T��<�m�<�<���<An�<a�<��<IG�<Rܿ<�l�<m��<���<��<i��<�<�x�<��<�\�<�Ȱ<o1�<O��<���<�U�<L��<��<\�<j��<���<yG�<���<�֜<��<k\�<<@ٕ<��<N�<���<ֻ�<M��<t#�<7U�<˅�<Y��<��<��<a>�<y�|<�,y<v�u<r�q</n<��j<��f<�/c<��_<e�[<'4X<ߌT<'�P<�BM<*�I<u�E<3aB<(�><�+;<a�7<�4<�q0<)�,<{\)<��%<�V"<��<c<��<�<<D�<f[
<�<ѳ<�i <�K�;\��;�f�;J	�;���;�{�;�K�;�+�;��;�;r-�;fO�;E��;�ƪ;)�;���;���;]��;%$�;.҉;z��;��~;��t;�zj;��`;L�V;M;q�C;w:;1�0;�';�;�;��;F;�q�:���:��:x|�:�A�:)<�:�i�:�ƅ:-�l:"N:�/::|7�9�ή9)j95F�8H�6[�Ӹ��X�ʏ���%ڹ�&���"�!�=��X��Ir��+���������V����q���ƺ1�Һ!ߺM�뺀����!�E�ta�*y����� �d�&���,��2�O�8�j�>���D��~J��oP��]V�K\��5b�0 h��n�t�s�<�y����Ԃ�Yȅ�
�������]�������r�������U����  �  �p=p=ȱ=�Q=��=��=�0=� =�n =p =<W�<��<���<��<HA�<�y�<-��<���<7�<�Q�< ��<(��<��<��<F�<s�<���<x��<���<��<�<�<�_�<b��<ݠ�<c��<���<.��<N
�<)�<�1�<�A�<�N�<�Y�<�a�<g�<~i�<�h�<?e�<j^�<\T�<�F�<06�<�!�<�	�<���<C��<.��<?��<AZ�<^+�<Z��<=��<��<SF�<~�<Y��<�m�<�<���<Hn�<S�<��<LG�<Sܿ<�l�<Z��<���<�<Z��<*�<�x�<��<�\�<�Ȱ<o1�<Z��<���<�U�<R��<��<\�<g��<���<zG�<w��<�֜<��<�\�<���<Eٕ<��<N�<���<˻�<Q��<j#�<8U�<˅�<P��<��<��<h>�<_�|<�,y<{�u<��q</n<g�j<��f<}/c<��_<��[<+4X<�T<�P<�BM<-�I<��E<%aB<!�><�+;<H�7<�4<�q0<?�,<f\)<��%<�V"<��<Kc<��<�<�<?�<r[
<�<׳<�i <�K�;8��;�f�;w	�;���;�{�;�K�;�+�;��;^�;I-�;5O�;0��;�ƪ;R�;˃�;���;l��;�#�;L҉;���;��~;C�t;�zj;Ĉ`;&�V;M;>�C;�:;��0;�';)�;H�;p�;/F;�q�:���:���:N|�:�A�:<�: i�: ǅ:0�l:�"N:�/:�:#4�9Ϯ9�j9�F�8//�6q�ӸW Y�[���S)ڹA$�E�"��=��X�EJr��+�����q���!����q���ƺ�Һ7!ߺ*��m���"� E�9a�gx�݉�v� ���&��,���2���8�J�>��D��~J��oP��]V��J\��5b��h��n�Q�s�*�y����~Ԃ��ȅ����󱋻b���X���k�������{����  �  �p=m=ɱ=�Q=��=��=�0=� =�n =q ==W�<��<���<��<FA�<�y�<-��<���<;�<�Q�<���<7��<��<��<F�<s�<���<x��<���<��<�<�<�_�<`��<��<n��<���<3��<Y
�<�<�1�<�A�<�N�<�Y�<�a�<%g�<|i�<�h�<:e�<r^�<eT�<�F�<66�<�!�<

�<w��<9��<&��<+��<MZ�<]+�<`��<0��<��<]F�<y�<g��<�m�<�<���<Mn�<L�<��<WG�<Dܿ<m�<^��<���<��<\��<,�<�x�<��<�\�<�Ȱ<p1�<T��<���<�U�<`��<��<"\�<d��<���<~G�<x��<�֜<��<�\�<囗<:ٕ<��<
N�<Ņ�<»�<^��<g#�<9U�<υ�<O��<��<|�<o>�<O�|<�,y<q�u<q�q</n<w�j<��f<�/c<��_<o�[<4X<	�T< �P<�BM< �I<��E<&aB<$�><�+;<>�7<�4<�q0<E�,<h\)<��%<�V"<��<Fc<��<�<�<G�<i[
<x<��<�i <L�;.��;�f�;m	�;���;�{�;�K�;�+�;��;R�;S-�;^O�;}��;�ƪ;|�;���;���;���;�#�;d҉;d��;$�~;8�t;D{j;��`;^�V;]M;��C; :;��0;C�';��;��;4�;�E;Fr�:���:���:}{�:B�:�<�:�h�:�ǅ:�l:�#N:r�/:n:I2�9�Ϯ9)j9�7�8��6ҰӸ��X�;����(ڹ�#���"���=�-X�Jr��+��`�� ���i����p��ƺB�Һe!ߺ���6����!��D��a��x�U��ɖ �U�&��,�x�2��8�ߕ>�	�D��~J�goP��]V��J\�6b��h�-	n���s�Q�y���PԂ��ȅ�ʼ��ɱ��<�����������?��������  �  �p=l=Ʊ=�Q=��=��=�0=� =�n =o =2W�<��<���<��<;A�<�y�<0��<���<2�<�Q�<���<&��<��<��<F�<s�<w��<w��<���<��<�<�<�_�<d��<��<h��<���<8��<P
�<&�<�1�<�A�<�N�<�Y�<�a�<(g�<�i�<�h�<=e�<m^�<[T�<G�<06�<�!�<
�<}��<:��<#��<2��<LZ�<[+�<Z��<>��<��<TF�<|�<b��<�m�<�<���<Nn�<V�<��<TG�<Sܿ<�l�<e��<���<��<c��<,�<�x�<��<�\�<�Ȱ<q1�<K��<���<�U�<Y��<��<\�<e��<���<xG�<u��<�֜<��<x\�<<=ٕ<��<N�<���<ѻ�<N��<g#�<8U�<̅�<X��<��<z�<p>�<_�|<�,y<|�u<��q</n<z�j<��f<�/c<��_<��[<'4X< �T<�P<�BM<�I<��E<5aB<#�><�+;<D�7<�4<�q0<<�,<Q\)<��%<�V"<��<0c<��<�<�<5�<q[
<�<ҳ<�i <�K�;@��;�f�;B	�;��;�{�;�K�;�+�;��;b�;^-�;HO�;I��;�ƪ;X�;���;���;m��;�#�;c҉;J��;9�~;|�t;%{j;��`;:�V;M;\�C;�:;s�0;2�';��;��;�;�E;8r�:u��:���:`|�:�A�:<�:�h�:�ǅ:�l:r$N:��/::�4�9�ή9^	j9�E�8�G�6��Ӹ��X�o���B'ڹ$�W�"��=�X�dIr��+������������*q���ƺ8�ҺZ!ߺ�뺓���"��D��a��x����� �h�&�g�,���2��8�^�>�
�D��~J��oP��]V��J\�6b��h��n��s�$�y����pԂ�~ȅ����ձ��R���]���r���Q��������  �  �p=u=Ǳ=�Q=��=��=�0=� =�n =k =6W�<��<���<��<9A�<�y�<��<���<2�<�Q�<���<#��<$��<��<F�<�r�<���<���<���<��<�<�<�_�<_��<��<r��<���<C��<J
�<*�<�1�<�A�<�N�<�Y�<�a�< g�<ti�<�h�<Ce�<q^�<RT�<�F�<'6�<�!�<�	�<}��<9��<#��<5��<=Z�<_+�<P��<7��<څ�<UF�<��<[��<�m�<�<���<Kn�<Q�<��<OG�<Xܿ<�l�<m��<���<��<e��<&�<�x�<��<�\�<�Ȱ<x1�<\��<���<�U�<T��<��<\�<c��<���<tG�<w��<�֜<��<u\�<<4ٕ<��<N�<���<λ�<I��<r#�<7U�<Ņ�<F��<��<��<i>�<h�|<�,y<{�u<��q</n<��j<��f<�/c<��_<��[<(4X<��T<�P<�BM<A�I<��E<aB<�><�+;<a�7<�4<�q0<.�,<Z\)<��%<�V"<��<-c<��<��<�<4�<_[
<~<̳<�i <�K�;��;~f�;w	�;��;�{�;�K�;�+�;��;N�;W-�;oO�;P��;�ƪ;@�;̓�;���;x��;�#�;N҉;���;��~;�t;�zj;�`;U�V;�M;(�C;~:;��0;Ƨ';��;��;�;�E;Dq�:���:���:�{�:FA�:$<�:_i�:>ǅ:�l:9#N:1�/:1:e3�9�Ϯ9�j9�K�8l��6�Ӹ�X� ����&ڹ�$��"��=�#X��Jr�\+���������ᾬ�wq���ƺL�Һt!ߺ�������	"�iE�ha��x����� ���&�?�,�ޡ2���8���>���D��~J��oP�<^V��J\�o5b��h��n�$�s�)�y�����Ԃ�=ȅ���������`���Z���q���d���l����  �  �p=m=ɱ=�Q=��=�=�0=� =�n =o =6W�<��<���<��<4A�<�y�<$��<���<3�<�Q�<���<+��<��<��<F�<s�<���<x��<���<��<�<�<�_�<i��<��<t��<���<=��<\
�<(�<�1�<�A�<�N�<�Y�<�a�<%g�<�i�<�h�<2e�<l^�<\T�<�F�<-6�<�!�<
�<z��<5��<!��<.��<DZ�<Z+�<V��<2��<���<VF�<q�<f��<�m�<�<���<Ln�<W�<��<XG�<Uܿ<m�<i��<���<��<g��<3�<�x�<��<�\�<�Ȱ<s1�<X��<���<�U�<Z��<��<\�<f��<���<vG�<t��<�֜<��<r\�<⛗<7ٕ<��<N�<���<ƻ�<U��<g#�<+U�<ׅ�<P��<��<��<m>�<j�|<�,y<w�u<��q<$/n<��j<��f<�/c<��_<��[<4X<�T<�P<�BM<"�I<��E<#aB<7�><�+;<@�7<�4<�q0<;�,<Y\)<��%<�V"<��<!c<��<�<�<5�<^[
<z<ڳ<~i <�K�;Z��;�f�;w	�;���;�{�;�K�;�+�;��;v�;t-�;wO�;X��;�ƪ;��;ƃ�;���;���;�#�;R҉;v��;"�~;V�t;S{j;V�`;.�V;M;�C;�:;~�0;��';��;Ҹ;�;�E;�q�:c��:O��:�{�:�A�:,<�:'h�:�ǅ:ƪl:$N:�/:D:�4�9�Ѯ9j9fH�8���6d�Ӹ&�X�����c&ڹG#���"�ם=�|X��Ir��+�� ���������q��aƺ�ҺO!ߺ͐뺯���#"�9E��a��x�q��� ���&�D�,���2�՝8�,�>��D�/J�#oP��]V��J\��5b��h��n���s�8�y����AԂ�]ȅ���������(���R�������H���g����  �  �p=k=̱=�Q=��=��=�0=� =�n =p =-W�<ߒ�<���<��<EA�<�y�<,��<���<.�<�Q�<��<*��<��<��<F�<s�<���<y��<���<��<�<�<�_�<k��<��<l��<���<4��<Z
�<+�<�1�<�A�<�N�<�Y�<�a�<-g�<|i�<�h�<9e�<k^�<VT�<�F�<26�<�!�<
�<s��<9��<)��<(��<JZ�<L+�<[��<4��<؅�<UF�<x�<a��<�m�<�<���<Wn�<Z�<��<^G�<Xܿ<m�<b��<���<��<b��<4�<�x�<��<�\�<�Ȱ<v1�<U��<���<�U�<Y��<��<\�<Z��<���<tG�<e��<�֜<��<�\�<盗<6ٕ<��<�M�<�<���<M��<h#�<6U�<υ�<M��<��<z�<}>�<]�|<�,y<��u<��q</n<q�j<��f<�/c<��_<��[<74X<�T<�P<�BM<�I<��E<!aB<(�><�+;<C�7<�4<�q0<A�,<H\)<�%<�V"<��<Dc<��<�<�<,�<n[
<g<ٳ<�i <�K�;4��;�f�;r	�;���;�{�;�K�;�+�;��;|�;d-�;UO�;u��;�ƪ;}�;у�;���;k��;�#�;�҉;c��;_�~;,�t;{j;��`;'�V;�M;��C;�:;�0;�';j�;��;B�;qE;r�:���:���:�{�:$A�:<�:�h�:�ǅ:�l:�$N:��/:�:�5�9Qή9�j9yJ�8X��6��Ӹ��X������'ڹ#���"��=�rX�DHr��+��O������B���0q��ƺ�Һ"ߺf�������"��D��a�~x�E��� ���&���,���2���8�f�>��D��~J�coP�^V�HJ\�"6b�Ph��n���s���y����JԂ��ȅ�ļ��ޱ��/���?���U���;��������  �  �p=n=ɱ=�Q=��=��=�0=� =�n =g =8W�<��<���<��<1A�<�y�<!��<���<1�<�Q�<���<"��<��<��<F�<s�<���<y��<���<��<�<�<�_�<_��<��<z��<���<K��<Q
�<+�<�1�<�A�<�N�<�Y�<�a�<g�<i�<�h�<Ce�<i^�<WT�<�F�< 6�<�!�< 
�<r��<-��<��<%��<BZ�<Z+�<N��<4��<ޅ�<PF�<��<Z��<�m�<�<���<Mn�<Y�<��<YG�<Xܿ<�l�<v��<���<��<t��<)�<�x�<��<�\�<�Ȱ<q1�<Z��<���<�U�<P��<��<\�<a��<���<rG�<v��<�֜<��<l\�<ݛ�<2ٕ<��<N�<���<˻�<G��<i#�<7U�<˅�<N��<��<�<n>�<l�|<�,y<��u<��q<"/n<��j<��f<�/c<��_<��[<24X<�T<�P<�BM<&�I<��E< aB<&�><�+;<L�7<�4<�q0<�,<^\)<��%<�V"<��<c<|�<��<�<0�<U[
<u<ɳ<�i <�K�;3��;�f�;r	�;���;�{�;�K�;�+�;��;L�;�-�;�O�;���;�ƪ;[�;΃�;���;���;�#�;]҉;x��;��~;G�t;�zj;ۈ`;�V;�M;�C;K:;~�0;�';]�;��;��;ZE;�q�:`��:���:�{�:�A�:�;�:Xi�:%ǅ:(�l:�"N:B�/:Q:<5�9�Ѯ9nj91J�8�-�6L�Ӹ��X�����7#ڹ}$���"�؝=�X��Ir��+�������=����q��$ƺV�Һ�!ߺ������"�KE�#b�#y����� ���&�8�,�(�2���8���>���D��~J��oP��]V��J\��5b��h��n���s��y����DԂ�;ȅ������������`���]���B���j����  �  �p=u=Ǳ=�Q=��=|�=�0=
� =�n =e =8W�<֒�<���<��<5A�<�y�<��<���</�<�Q�<��<��<��<��<!F�<s�<���<���<���<��<�<�<`�<g��<��<t��<���<C��<S
�<;�<�1�<�A�<�N�<�Y�<�a�<g�<�i�<�h�<8e�<i^�<_T�<�F�<6�<�!�<�	�<���<6��<!��<7��<2Z�<Z+�<K��<4��<��<LF�<{�<T��<�m�<	�<���<Mn�<X�<��<SG�<iܿ<�l�<q��<���<��<o��</�<y�<��<�\�<�Ȱ<x1�<^��<���<�U�<G��<��<
\�<q��<���<oG�<r��<�֜<��<r\�<뛗<:ٕ<��<	N�<���<ϻ�<H��<j#�<+U�<υ�<V��<��<��<k>�<x�|<�,y<��u<��q</n<��j<��f<�/c<��_<��[<B4X<�T<,�P<�BM<A�I<��E<*aB<1�><�+;<J�7<�4<�q0<�,<]\)<m�%<�V"<��<#c<��<�<�<,�<K[
<�<��<�i <�K�;c��;�f�;u	�;��;�{�;L�;�+�;7�;m�;�-�;rO�;,��;�ƪ;`�;��;���;���;�#�;S҉;���;��~;��t;�zj;��`;�V;,M;�C;=:;��0;Z�';٠;۸;�;�E;�p�:g��:���:�{�:GB�:�;�:�h�:�ƅ:'�l:W"N:��/:R:�4�9	Ү9Yj9G[�8`�6��Ӹ`�X�َ���$ڹ�#���"�,�=�!X��Ir�l+���������F���Er���ƺڢҺ� ߺ1��#���3"��E�za��x�*��ϖ �.�&�%�,�:�2���8���>��D�6J�coP��]V��J\�h5b��h��n��s���y�H��QԂ�Mȅ�$�������,���,���=���m���J����  �  �p=r=Ǳ=�Q=��=��=�0=� =�n =i =9W�<ْ�<���<��<4A�<�y�<%��<���<8�<�Q�<���< ��<��<��<F�<�r�<~��<���<���<��<�<�<�_�<c��<��<���<���<I��<Z
�<*�<�1�<�A�<O�<�Y�<�a�<g�<}i�<�h�<De�<k^�<UT�<�F�<,6�<�!�<�	�<p��<&��<��<#��<AZ�<U+�<Y��<%��<ۅ�<OF�<��<`��<�m�<�<���<Un�<_�<��<XG�<Xܿ<m�<t��<���<��<n��</�<�x�<��<�\�<�Ȱ<|1�<T��<���<�U�<X��<��<\�<a��<���<{G�<i��<�֜<��<n\�<ٛ�<1ٕ<��<N�<���<���<F��<n#�<<U�<΅�<G��<��<��<x>�<{�|<�,y<��u<��q<"/n<��j<
�f<�/c<��_<��[<64X< �T<,�P<�BM<8�I<��E<aB<)�><�+;<R�7<�4<�q0<&�,<_\)<s�%<�V"<��< c<w�<�<�<>�<K[
<r<ĳ<�i <�K�;<��;zf�;Z	�;��;�{�;�K�;�+�;��;\�;�-�;�O�;���;�ƪ;|�;˃�;���;|��;$�;x҉;���;��~;5�t;{j;�`;&�V;�M;��C;�:;k�0;Ƨ';N�;^�;��;HE;~q�:��:u��:�z�:TA�:�;�:Yi�:�ǅ:��l:�"N:~�/:I:�6�9�Ю9�
j9PJ�8��6��Ӹ�X�[����$ڹ�#���"��=��X��Hr�*+��t������뽬�;q��Gƺ��Һ�!ߺ���o���w"�3E�;b�y����� ��&�6�,��2��8���>�ԋD��~J�ioP�6^V��J\��5b�uh�{n�
�s���y����EԂ�+ȅ�����}���&���K���U���Q���M����  �  Dr==��= T=T�=G�=�3=i� =�r =Z =�_�<���<���<O�<aL�<_��<���<���<!+�<P`�<n��<d��<��<�)�<�X�<���<��<���<�<�.�<�T�< y�<���<���<y��<���<Y�<�)�<i?�<�R�<�c�<lr�<H~�<x��<܍�<H��<ґ�<&��<^��<h��<�s�<+d�<�P�<�9�</�<� �<���<S��<7��<�_�<�-�<���<)��<�|�<{9�<���<^��<�T�<���<��<�G�<^��<f~�<�<U��<1/�<ƶ�<:�<@��<G4�<��<�<	��<&��<�_�<Kí<�#�<=��<�٨<�/�<���<�ң<��<�i�<J��<R��<�8�<�x�<˶�<��<g,�<Nd�<}��<�Ύ<�<y3�<�c�<Ғ�<���<��<��<"E�<��|<24y<��u<��q<-n<<j<��f<$c<9w_<��[<LX<uT<�P<�$M<�~I<,�E<�9B<��><�:<cd7<�3<�:0<�,<2)<L�%<�"<q�<'<W�<4<��<�c<�
<P�<W<
 <��;�	�;D��;k7�;���;X��;�m�;5J�;�6�;h4�;�B�;�a�;���;�ԩ;)�;��;��;��;�,�;5ۈ;���;��|;��r;E�h;b�^;T�T;�.K;�A;�C8;� /;��%;n�;�;�<;'�;�)�:GY�:���:�e�:k>�:�I�:ǈ�:d��:a4g:�H:��*:?:[q�9]X�9z�W9���8jt-�����i��X���������{&���@�+J[��hu�[���{���%Y���������KǺd�Ӻ]>�|��-������ĺ�;�����:��M� ���&�%�,�[�2�M�8���>���D�ɺJ�Y�P���V��x\��_b�2Eh��)n�Ct���y�R��܂�@΅�����\���}�������Џ��d����|���  �  Lr==��= T=L�=C�=�3=b� =�r =Y =�_�<���<���<L�<GL�<^��<���<���<+�<J`�<g��<X��<#��<�)�<�X�<���<��<���<"�<�.�<�T�<y�<p��<��<���<
��<d�<|)�<l?�<�R�<�c�<xr�<_~�<���<֍�<H��<���<(��<]��<Q��<�s�<)d�<�P�<�9�<8�<� �<���<Y��</��<�_�<�-�<���<��<�|�<�9�<���<[��<�T�<���<���<�G�<`��<k~�<�<B��<5/�<Ѷ�<#:�<7��<44�<'��<
�<��<5��<�_�<Wí<�#�<5��<�٨<�/�<���<�ң<��<�i�<T��<H��<�8�<�x�<Ŷ�<��<g,�<Ud�<{��<�Ύ<��<�3�<�c�<���<���<��<��<3E�<��|<%4y<��u<��q<�,n<_j<��f<<$c<w_<��[<jX<uT<�P<�$M<�~I<+�E<�9B<y�><�:<�d7<��3<�:0<�,<<)<S�%<�"<k�<�<V�<4<��<�c<�
<B�<�V<.
 <��;d	�;>��;�7�;���;���;�m�;J�;�6�; 4�;KB�;�a�;���;	թ;�(�;��;��;��;.-�;�ۈ;;��|;��r;��h;w�^;M�T;(.K;��A;�C8;/;��%;��;��;:<;Z�;o)�:/Z�:���:Ge�:=�:uI�:B��:P��:4g:F�H:��*:�:u�9�X�9�W9ʺ�8.�v����i��U��0��9���y&��@��I[�gu�Ъ��Ì��eY��&��h���JǺ�Ӻ�>��캊���H����9��g��j��� ���&���,�c�2�b�8��>���D��J�ܦP���V��x\�&_b��Dh�~)n�wt��y����T܂��ͅ�X������Ҧ�������������w|���  �  Er==��=%T=Q�=B�=�3=c� =�r =W =�_�<���<���<[�<JL�<r��<���<���<+�<L`�<w��<Z��<*��<�)�<�X�<���<��<���<�<�.�<�T�<y�<r��<���<���<���<c�<)�<r?�<�R�<�c�<nr�<O~�<y��<֍�<Y��<���<,��<b��<[��<t�<!d�<�P�<�9�<@�<� �<���<f��<#��<�_�<�-�<���<!��<�|�<�9�<���<j��<�T�<���<��<�G�<Y��<d~�<�<E��<6/�<���<:�<=��<64�<.��<�<��<(��<�_�<Pí<�#�<@��<�٨<�/�<���<�ң<��<�i�<Y��<?��<�8�<�x�<ж�<��<^,�<Sd�<v��<ώ<��<�3�<�c�<ƒ�<���<��<��<%E�<��|<4y<��u<��q<�,n<Wj<v�f<.$c<w_<��[<tX<uT<�P<�$M<�~I< �E<�9B<��><�:<�d7<��3<�:0<�,<3)<H�%<�"<��<�<~�<�3<��<qc<�
<c�<�V<<
 <��;�	�;V��;x7�;���;V��;�m�;J�;7�;,4�;eB�;�a�;b��;թ;�(�;+��;��;쐓;-�;Sۈ;ě�;��|;@�r;��h;��^;z�T;{.K;H�A;�C8;+/;H�%;��;��;n<;��;�(�:zZ�:���:7f�:�=�:�I�:v��:��:�5g:��H:��*:|:r�9)W�9��W9��8Y�-�����$i�X���������x&���@��J[��hu�ͫ��,���'Y��n�������IǺ��Ӻ >�x��3���!��U�����8����� ���&���,���2���8���>�\�D��J���P��V��x\��_b�Eh��)n��t���y�q��N܂�΅�����2���˦��������������~|���  �  Lr==��=T=Q�=F�=�3=d� =�r =X =�_�<��<���<U�<LL�<i��<���<���<!+�<N`�<e��<]��<��<�)�<�X�<���<��<���<"�<�.�<�T�<�x�<r��<���<��<��<\�<�)�<a?�<�R�<�c�<wr�<W~�<~��<ݍ�<E��<Ǒ�<&��<Z��<T��<�s�<#d�<�P�<�9�<;�<� �<���<^��<2��<�_�<�-�<���<��<�|�<{9�<���<\��<�T�<���<��<�G�<d��<e~�<�<N��<1/�<˶�<:�<:��<74�<��<�<��<3��<�_�<Ví<�#�<9��<�٨<�/�<���<�ң<��<�i�<[��<J��<�8�<�x�<̶�<��<k,�<Zd�<x��<�Ύ<��<{3�<�c�<ɒ�<���<��<��<3E�<��|<24y<��u<��q< -n<Bj<��f<$c<$w_<��[<FX< uT<�P<�$M<�~I<3�E<�9B<��><�:<hd7<��3<�:0<�,<B)<[�%<�"<|�<�<m�<4<��<�c<�
<?�<�V<
 <��;�	�;2��;�7�;���;���;�m�;GJ�;�6�;,4�;gB�;�a�;���;�ԩ;)�;뎞;��;��;)-�;tۈ;ڛ�;��|;��r;�h;d�^;3�T;E.K;ЧA;�C8;G/;��%;��;��;O<;��;�)�:�Z�:��:|e�:+=�:fI�:ӈ�:���:$4g:2�H:�*:4:dt�9Z�9�W9��8��-�����i�gW��f�����Y|&�z�@��I[�Egu�����ь��OY�����ն���JǺ��Ӻ$?຦�캒�����������7��3��4� ���&���,���2�R�8���>���D�κJ���P���V��x\�Q_b��Dh�y)n�Ct���y����%܂�5΅�i���Y�����������ݏ��b���r|���  �  Mr==��=T=O�=E�=�3=n� =�r =` =�_�<���<���<W�<WL�<g��<���<���<+�<Y`�<f��<r��<��<�)�<�X�<���<��<���< �<�.�<�T�<y�<{��<��<w��<��<M�<�)�<c?�<�R�<�c�<hr�<Y~�<t��<ߍ�<?��<ʑ�<$��<l��<_��<�s�<1d�<�P�<�9�<=�<� �<���<_��<6��<�_�<�-�<���<��<}�<z9�<���<R��<�T�<���<��<�G�<S��<n~�<�<R��<#/�<̶�<:�</��<A4�<��<�<�<,��<�_�<Qí<�#�<.��<�٨<�/�<���<�ң<��<�i�<Q��<S��<�8�<�x�<Ѷ�<��<j,�<Od�<���<�Ύ<�<�3�<�c�<Ȓ�<���<��<��<6E�<��|<%4y<��u<��q<�,n<)j<��f<$c<w_<��[<\X<uT<��P<�$M<�~I<5�E<�9B<��><�:<{d7<�3<�:0</�,<0)<X�%<�"<��<<i�<4<��<}c<�
<A�<!W<
 <��;Z	�;,��;�7�;���;���;qm�;PJ�;�6�;P4�;>B�;�a�;���;�ԩ;)�;�;��;萓;�,�;}ۈ;���;��|;m�r;
�h;Z�^;��T;�.K;��A;	D8;� /;��%;��;�;�<;��;�)�:�Y�:���:f�:�=�:�J�:���:C��:�2g:I�H:�*:�:�p�9�U�9�W9��8_�-�4	��Mi��X���ṑ���{&���@��L[�(hu��������qY����������JǺe�Ӻ�>���v���_�������������� ���&��,���2�[�8�j�>���D�ѺJ���P�אV��x\��_b��Dh�,*n�wt�6�y����'܂�g΅�K�������������������n����|���  �  Lr==��=#T=S�=D�=�3=c� =�r =^ =�_�<��<���<Z�<TL�<n��<���<���<+�<X`�<k��<]��<��<�)�<�X�<���<��<���< �<�.�<�T�<y�<o��<��<���<���<\�<�)�<Z?�<�R�<�c�<qr�<V~�<s��<؍�<P��<ɑ�<$��<g��<U��<�s�<*d�<�P�<�9�<B�<� �<���<g��<3��<�_�<�-�<���<��<�|�<z9�<���<a��<�T�<}��<��<�G�<Z��<a~�< �<G��<//�<���<:�<8��<44�<��<�<��<.��<�_�<Jí<�#�<<��<�٨<�/�<���<�ң<��<�i�<f��<L��<�8�<�x�<Ҷ�<��<r,�<Vd�<���<�Ύ<��<�3�<�c�<̒�<���<��<��<0E�<��|<4y<��u<r�q<�,n<Ej<q�f<!$c<w_<��[<VX<
uT<�P<�$M<�~I<(�E<�9B<��><�:<}d7<��3<�:0<)�,<;)<r�%<�"<��<<x�<4<�<�c<�
<K�<�V<%
 <��;�	�;V��;x7�;���;���;�m�;J�;�6�;!4�;^B�;�a�;`��;�ԩ;�(�;ώ�;��;;-�;pۈ;���;��|;��r; �h;X�^;��T;L.K;2�A;�C8;F/;��%;�;��;k<;Ι;�)�:�Z�:���:nf�:S=�:J�:ƈ�:���:�4g:��H:��*::�r�9�W�9��W9���8�-�h���xi�
X�����$���{&���@��J[��gu�꫇�����Y�����󶺺�JǺ��Ӻ�>���캉�����������	�����	� �W�&���,�!�2�=�8��>�~�D�غJ���P�H�V��x\��_b��Dh��)n��t�b�y����1܂�.΅�����K�������ښ�����������|���  �  Br==��=T=P�=G�=�3=b� =�r =[ =�_�<��<���<i�<JL�<}��<���<���<+�<W`�<w��<\��<)��<�)�<�X�<���<��<���<�<�.�<�T�<y�<i��<��<~��<���<`�<r)�<d?�<�R�<�c�<pr�<O~�<���<э�<H��<�<-��<g��<V��<t�<$d�<�P�<�9�<G�<� �<���<o��<,��<�_�<�-�< ��<��<�|�<�9�<���<[��<�T�<���<��<�G�<\��<Y~�<�<7��<1/�<���<:�<3��<*4�<��<��<��<!��<�_�<Rí<}#�<7��<�٨<�/�<���<�ң<��<�i�<e��<D��<�8�<�x�<޶�<��<n,�<]d�<}��<ώ<��<�3�<�c�<Œ�<���<��<��< E�<��|<4y<��u<�q<�,n<Lj<k�f<&$c<w_<��[<RX<�tT<�P<$M<�~I<*�E<�9B<��><�:<�d7<��3<�:0<�,<F)<j�%<�"<��<�<��<�3<�<�c<�
<c�<�V<=
 <���;~	�;'��;�7�;���;D��;�m�;�I�;�6�;4�;BB�;�a�;S��;�ԩ;�(�;���;��;�;-�;Tۈ;;��|;��r;Ȓh;��^;��T;[.K;~�A;�C8;�/;��%;/�;)�;�<;�;B)�:>[�:&��:�f�:�=�:J�:���:���:$4g:��H:y�*:�:~q�9EX�9c�W9R��8a.�����i�!Y��ū�g���z&���@��I[�uiu���������Y�����R����IǺ��Ӻ3>�ڠ캛������0��H��9�����
� �x�&���,�Z�2���8��>�^�D���J���P���V��x\�-_b�BEh�u)n��t�z�y����t܂�!΅�����B���즎�Ϛ��ŏ������o|���  �  Cr==��=!T=V�=E�=�3=l� =�r =_ =�_�<��<���<h�<NL�<z��<���<���<"+�<Z`�<q��<j��<��<�)�<�X�<���<��<���<�<�.�<�T�<�x�<l��<��<s��<���<R�<z)�<d?�<�R�<�c�<hr�<O~�<s��<׍�<M��<ˑ�<#��<d��<a��< t�<-d�<�P�<�9�<I�<� �<���<n��<:��<�_�<�-�<���<"��<�|�<x9�<���<`��<�T�<}��<��<�G�<X��<_~�<�<>��<&/�<���<:�<0��<.4�<��< �<���<��<�_�<Ií<�#�<@��<�٨<�/�<���<�ң<��<�i�<[��<V��<�8�<�x�<߶�<��<s,�<Zd�<���<ώ<�<3�<�c�<ђ�<���<��<��<"E�<��|<4y<��u<��q<�,n</j<��f<$c<w_<��[<HX<uT<��P<�$M<�~I<#�E<�9B<��><�:<nd7<�3<�:0<,�,<G)<i�%<�"<��<<��<4<��<�c<�
<Y�<W<
 <��;�	�;H��;u7�;���;A��;�m�;J�;�6�;4�;>B�;�a�;a��;�ԩ;�(�;���;��;琓;�,�;Tۈ;���;��|;�r;�h;W�^;��T;�.K;J�A;�C8;A/;�%;D�;T�;�<;�;,*�:�Z�:���:f�:	>�:7J�:���:)��:�4g:��H:��*:�:6p�9W�9��W9��8�&.�B���i�K[���������{&�"�@�;K[��iu���������/Y��c��߶���JǺ�ӺG>�۠�^��������l��������� �N�&���,��2� �8�s�>���D�ɺJ�b�P�k�V��x\��_b�6Eh��)n��t���y����a܂�[΅���������㦎�����ُ�������|���  �  Nr==��=T=N�=I�=�3=m� =�r =d =�_�<��<���<[�<kL�<k��<���<���<)+�<]`�<b��<p��<��<�)�<�X�<���<��<���< �<�.�<�T�<�x�<f��<��<t��<���<I�<�)�<O?�<�R�<�c�<gr�<`~�<r��<ݍ�<>��<Ǒ�<)��<h��<^��<�s�<;d�<�P�<�9�<>�<� �<���<b��<F��<�_�<�-�<���<��<}�<}9�<���<P��<�T�<}��<���<�G�<R��<b~�<��<C��</�<���<:�<-��<+4�<��<�<���<+��<�_�<Jí<�#�<-��<�٨<�/�<���<�ң<��<�i�<e��<]��<�8�< y�<ն�<��<,�<[d�<���<�Ύ<�<�3�<�c�<Œ�<���<��<��<7E�<��|<4y<��u<]�q<�,n<!j<��f<�#c<w_<��[<?X<uT<��P<�$M<�~I<'�E<�9B<��>< �:<vd7<�3<�:0<B�,<J)<��%<�"<��<=<q�<&4<�<�c<�
<<�<W<#
 <'��;[	�;A��;z7�;���;���;�m�;*J�;�6�;�3�;BB�;�a�;j��;�ԩ;�(�;���;��;ᐓ;�,�;�ۈ;���;��|;j�r;��h;��^;��T;�.K;֧A;bD8;C/;z�%;��;b�;=;��;�*�:�Z�:���:�e�:�=�:fJ�:���:0��:�2g:L�H:��*:X:Eq�9�U�9��W9���8'�-�"��i��Z����$���}&�:�@��K[�(hu�z���q���0Y�����q����JǺ��Ӻ�>�Ԡ��������e�����V������� ���&���,���2���8�q�>���D���J���P�אV��x\��_b��Dh� *n��t���y�K��B܂�u΅���������̦������ꏔ������|���  �  Dr==��=T=O�=H�=�3=l� =�r =e =�_�<��<���<d�<fL�<x��<���<���<+�<e`�<w��<m��<%��<�)�<�X�<���<��<���<�<�.�<�T�<y�<g��<��<m��<���<K�<w)�<Z?�<�R�<�c�<cr�<J~�<r��<ٍ�<J��<ɑ�</��<h��<g��<	t�<6d�<�P�<�9�<J�<� �<���<o��<@��<�_�<�-�<��<(��<�|�<�9�<���<\��<�T�<~��<��<�G�<H��<W~�<��<<��</�<���<:�<)��<*4�<��<��<���<��<�_�<Kí<�#�<2��<�٨<�/�<���<�ң<��<�i�<c��<Z��<�8�<�x�<ܶ�<��<w,�<Rd�<���<ώ<�<�3�<�c�<ƒ�<���<��<��<"E�<��|<4y<��u<j�q<�,n<$j<n�f<�#c<w_<��[<QX<�tT<��P<�$M<�~I<)�E<�9B<��><�:<�d7<�3<�:0<D�,<7)<u�%<�"<��<1<��<$4<�<�c<	
<f�<W<6
 <%��;q	�;:��;z7�;���;P��;�m�;�I�;�6�;4�;*B�;�a�;M��;�ԩ;�(�;Ў�;��;���;�,�;Aۈ;���;��|;ѥr;�h;��^;��T;�.K;��A;7D8;3/;/�%;J�;�;
=;�;�*�:�Z�:���:g�:l>�:GJ�:g��:2��:[4g:��H:��*:�:To�9jS�9R�W9���8G,.�A��ki�Z\����8���{&��@�ML[��iu�|���f���mY��4������
JǺ��Ӻ�=���u���ɝ���n��q������� �2�&��,���2���8�q�>�i�D���J���P���V��x\��_b�4Eh� *n��t�m�y���c܂�q΅���������覎��Ə��Å���|���  �  Cr==��=T=V�=D�=�3=f� =�r =^ =�_�<��<���<m�<QL�<���<���<���</+�<Z`�<q��<_��<��<�)�<�X�<���<��<���<�<�.�<�T�<�x�<X��<��<q��<���<V�<l)�<X?�<�R�<�c�<tr�<G~�<���<̍�<S��<ȑ�<*��<d��<]��< t�<,d�<�P�<�9�<M�<� �<���<s��<9��<	`�<�-�<���<��<�|�<9�<���<h��<�T�<���<��<�G�<R��<S~�<��<.��<&/�<���<	:�<-��<4�<��<��<��<$��<�_�<Oí<w#�<H��<�٨<�/�<���<�ң<��<�i�<q��<P��<�8�<�x�<㶗<��<x,�<ld�<���<	ώ<��<�3�<�c�<ђ�<���<��<��<E�<��|<�3y<|�u<a�q<�,n<4j<l�f<
$c<w_<��[<@X<�tT<�P<�$M<�~I<�E<�9B<��><�:<{d7<��3<�:0<)�,<i)<z�%<�"<��<<��<4<$�<�c<�
<Y�<�V<*
 <��;�	�;*��;|7�;���;S��;�m�;�I�;�6�;�3�;:B�;�a�;V��;�ԩ;�(�;ˎ�;��;ϐ�;"-�;:ۈ;ꛃ;h�|;�r;�h;��^;��T;�.K;K�A;�C8;/;�%;h�;Q�;�<;7�;"*�:#\�:���:{f�:�=�:�I�:$��:���:�5g:��H:]�*:�:�r�9�U�9�W9N��8�.�[��}i�{[����L��L|&�[�@�_J[� iu�˫��"����Y��������dJǺ��Ӻq>�Ӡ�����W��ͺ�+��	��w���� �*�&�.�,�0�2���8���>���D�ԺJ�\�P�{�V��x\�+_b�HEh�s)n�t���y�;��x܂�Q΅�����y���즎����揔�΅��m|���  �  Ar==��=T=R�=G�=�3=l� =�r =a =�_�<��<���<t�<jL�<���<���<���<-+�<_`�<v��<n��<+��<�)�<�X�<���<��<���<�<�.�<�T�<�x�<b��<��<g��<���<C�<v)�<S?�<�R�<�c�<er�<F~�<}��<ύ�<F��<ő�<1��<t��<i��<t�<3d�<�P�<�9�<H�<� �<���<q��<5��<`�<�-�< ��<+��<}�<�9�<���<Y��<�T�<���<ߥ�<�G�<D��<]~�<��<:��</�<���<:�<'��<&4�<��<��<�<��<�_�<Lí<w#�<6��<�٨<�/�<���<�ң<��<�i�<m��<N��<�8�<y�<궗<��<u,�<hd�<���<ώ<�<�3�<�c�<˒�<���<��<��<E�<��|<�3y<��u<b�q<�,n<j<d�f<�#c<w_<��[<KX<�tT<��P<{$M<�~I<�E<�9B<��><�:<�d7<�3<�:0<3�,<^)<r�%<�"<��<;<��<4<�<�c< 
<e�<W<C
 <��;�	�;$��;w7�;���;C��;�m�;�I�;�6�;�3�;6B�;pa�;<��;�ԩ;�(�;���;��;���;�,�;4ۈ;ܛ�;��|;��r;�h;ƣ^;�T;�.K;x�A;&D8;�/;�%;=�;��;7=;!�;�)�:�[�:0��:�f�:�>�:K�:���:���:4g:d�H:��*:p:�o�9�R�9��W9ˡ�8�=.����� i�a]����ṷ��c|&�q�@��L[�ju�*���Q����Y���������IǺ��Ӻ�=�c�캰���{��޺�#��D��A���� �?�&�U�,��2���8�u�>�!�D���J���P�ɐV��x\�`_b�VEh��)n�t���y�5��`܂��΅���������ߦ�� ���ҏ��ǅ���|���  �  Hr==��="T=R�=F�=�3=e� =�r =d =�_�<��<���<c�<XL�<t��<���<���< +�<d`�<p��<\��<��<�)�<�X�<���<��<���<!�<�.�<�T�<�x�<d��<��<n��<���<A�<)�<H?�<�R�<�c�<qr�<P~�<n��<ڍ�<M��<ʑ�<$��<Z��<Y��<t�<4d�<�P�<�9�<N�<� �<���<r��<I��<�_�<�-�<���<��<�|�<y9�<���<^��<�T�<|��<��<�G�<M��<d~�<��<C��</�<���<
:�<��<*4�<��<��<���<1��<�_�<Jí<�#�<6��<�٨<�/�<���<�ң<��<�i�<k��<^��<�8�<�x�<׶�<��<�,�<Yd�<���<
ώ<��<3�<�c�<˒�<���<��<��<)E�<��|<4y<��u<T�q<�,n<j<��f<�#c<w_<��[<EX<�tT<��P<�$M<�~I<1�E<�9B<��><�:<sd7<��3<�:0<B�,<@)<��%<�"<��<<��<34<&�<�c<
<W�<�V<*
 <!��;�	�;i��;z7�;���;���;�m�;�I�;�6�;�3�;B�;�a�;���;�ԩ;�(�;���;��;ǐ�;-�;^ۈ;���;��|;�r;�h;_�^;B�T;w.K;`�A;*D8;c/;��%;o�;X�;�<;*�;,+�:5[�:���:�f�:�=�:WI�:�:+��:�4g:E�H:��*::t�9�T�9��W9��8X�-����Ji�Q[�����?��~&�R�@��K[�Qgu�U���r����X���������[JǺ��Ӻ�>�6��E������]�����������p� ���&���,���2���8���>���D�ߺJ���P�]�V��x\��_b��Dh��)n��t���y�p��U܂��΅�w�������禎����ݏ�������|���  �  Ar==��=T=R�=G�=�3=l� =�r =a =�_�<��<���<t�<jL�<���<���<���<-+�<_`�<v��<n��<+��<�)�<�X�<���<��<���<�<�.�<�T�<�x�<b��<��<g��<���<C�<v)�<S?�<�R�<�c�<er�<F~�<}��<ύ�<F��<ő�<1��<t��<i��<t�<3d�<�P�<�9�<H�<� �<���<q��<5��<`�<�-�< ��<+��<}�<�9�<���<Y��<�T�<���<ߥ�<�G�<D��<]~�<��<:��</�<���<:�<'��<&4�<��<��<�<��<�_�<Lí<w#�<6��<�٨<�/�<���<�ң<��<�i�<m��<N��<�8�<y�<궗<��<u,�<hd�<���<ώ<�<�3�<�c�<˒�<���<��<��<E�<��|<�3y<��u<b�q<�,n<j<d�f<�#c<w_<��[<KX<�tT<��P<{$M<�~I<�E<�9B<��><�:<�d7<�3<�:0<3�,<^)<r�%<�"<��<;<��<4<�<�c< 
<e�<W<C
 <��;�	�;$��;w7�;���;C��;�m�;�I�;�6�;�3�;6B�;pa�;<��;�ԩ;�(�;���;��;���;�,�;4ۈ;ܛ�;��|;��r;�h;ƣ^;�T;�.K;x�A;&D8;�/;�%;=�;��;7=;!�;�)�:�[�:0��:�f�:�>�:K�:���:���:4g:d�H:��*:p:�o�9�R�9��W9ˡ�8�=.����� i�a]����ṷ��c|&�q�@��L[�ju�*���Q����Y���������IǺ��Ӻ�=�c�캰���{��޺�#��D��A���� �?�&�U�,��2���8�u�>�!�D���J���P�ɐV��x\�`_b�VEh��)n�t���y�5��`܂��΅���������ߦ�� ���ҏ��ǅ���|���  �  Cr==��=T=V�=D�=�3=f� =�r =^ =�_�<��<���<m�<QL�<���<���<���</+�<Z`�<q��<_��<��<�)�<�X�<���<��<���<�<�.�<�T�<�x�<X��<��<q��<���<V�<l)�<X?�<�R�<�c�<tr�<G~�<���<̍�<S��<ȑ�<*��<d��<]��< t�<,d�<�P�<�9�<M�<� �<���<s��<9��<	`�<�-�<���<��<�|�<9�<���<h��<�T�<���<��<�G�<R��<S~�<��<.��<&/�<���<	:�<-��<4�<��<��<��<$��<�_�<Oí<w#�<H��<�٨<�/�<���<�ң<��<�i�<q��<P��<�8�<�x�<㶗<��<x,�<ld�<���<	ώ<��<�3�<�c�<ђ�<���<��<��<E�<��|<�3y<|�u<a�q<�,n<4j<l�f<
$c<w_<��[<@X<�tT<�P<�$M<�~I<�E<�9B<��><�:<{d7<��3<�:0<)�,<i)<z�%<�"<��<<��<4<$�<�c<�
<Y�<�V<*
 <��;�	�;*��;|7�;���;S��;�m�;�I�;�6�;�3�;:B�;�a�;V��;�ԩ;�(�;ˎ�;��;ϐ�;"-�;:ۈ;ꛃ;h�|;�r;�h;��^;��T;�.K;K�A;�C8;/;�%;h�;Q�;�<;7�;"*�:#\�:���:{f�:�=�:�I�:$��:���:�5g:��H:]�*:�:�r�9�U�9�W9N��8�.�[��}i�{[����L��L|&�[�@�_J[� iu�˫��"����Y��������dJǺ��Ӻq>�Ӡ�����W��ͺ�+��	��w���� �*�&�.�,�0�2���8���>���D�ԺJ�\�P�{�V��x\�+_b�HEh�s)n�t���y�;��x܂�Q΅�����y���즎����揔�΅��m|���  �  Dr==��=T=O�=H�=�3=l� =�r =e =�_�<��<���<d�<fL�<x��<���<���<+�<e`�<w��<m��<%��<�)�<�X�<���<��<���<�<�.�<�T�<y�<g��<��<m��<���<K�<w)�<Z?�<�R�<�c�<cr�<J~�<r��<ٍ�<J��<ɑ�</��<h��<g��<	t�<6d�<�P�<�9�<J�<� �<���<o��<@��<�_�<�-�<��<(��<�|�<�9�<���<\��<�T�<~��<��<�G�<H��<W~�<��<<��</�<���<:�<)��<*4�<��<��<���<��<�_�<Kí<�#�<2��<�٨<�/�<���<�ң<��<�i�<c��<Z��<�8�<�x�<ܶ�<��<w,�<Rd�<���<ώ<�<�3�<�c�<ƒ�<���<��<��<"E�<��|<4y<��u<j�q<�,n<$j<n�f<�#c<w_<��[<QX<�tT<��P<�$M<�~I<)�E<�9B<��><�:<�d7<�3<�:0<D�,<7)<u�%<�"<��<1<��<$4<�<�c<	
<f�<W<6
 <%��;q	�;:��;z7�;���;P��;�m�;�I�;�6�;4�;*B�;�a�;M��;�ԩ;�(�;Ў�;��;���;�,�;Aۈ;���;��|;ѥr;�h;��^;��T;�.K;��A;7D8;3/;/�%;J�;�;
=;�;�*�:�Z�:���:g�:l>�:GJ�:g��:2��:[4g:��H:��*:�:To�9jS�9R�W9���8G,.�A��ki�Z\����8���{&��@�ML[��iu�|���f���mY��4������
JǺ��Ӻ�=���u���ɝ���n��q������� �2�&��,���2���8�q�>�i�D���J���P���V��x\��_b�4Eh� *n��t�m�y���c܂�q΅���������覎��Ə��Å���|���  �  Nr==��=T=N�=I�=�3=m� =�r =d =�_�<��<���<[�<kL�<k��<���<���<)+�<]`�<b��<p��<��<�)�<�X�<���<��<���< �<�.�<�T�<�x�<f��<��<t��<���<I�<�)�<O?�<�R�<�c�<gr�<`~�<r��<ݍ�<>��<Ǒ�<)��<h��<^��<�s�<;d�<�P�<�9�<>�<� �<���<b��<F��<�_�<�-�<���<��<}�<}9�<���<P��<�T�<}��<���<�G�<R��<b~�<��<C��</�<���<:�<-��<+4�<��<�<���<+��<�_�<Jí<�#�<-��<�٨<�/�<���<�ң<��<�i�<e��<]��<�8�< y�<ն�<��<,�<[d�<���<�Ύ<�<�3�<�c�<Œ�<���<��<��<7E�<��|<4y<��u<]�q<�,n<!j<��f<�#c<w_<��[<?X<uT<��P<�$M<�~I<'�E<�9B<��>< �:<vd7<�3<�:0<B�,<J)<��%<�"<��<=<q�<&4<�<�c<�
<<�<W<#
 <'��;[	�;A��;z7�;���;���;�m�;*J�;�6�;�3�;BB�;�a�;j��;�ԩ;�(�;���;��;ᐓ;�,�;�ۈ;���;��|;j�r;��h;��^;��T;�.K;֧A;bD8;C/;z�%;��;b�;=;��;�*�:�Z�:���:�e�:�=�:fJ�:���:0��:�2g:L�H:��*:X:Eq�9�U�9��W9���8'�-�"��i��Z����$���}&�:�@��K[�(hu�z���q���0Y�����q����JǺ��Ӻ�>�Ԡ��������e�����V������� ���&���,���2���8�q�>���D���J���P�אV��x\��_b��Dh� *n��t���y�K��B܂�u΅���������̦������ꏔ������|���  �  Cr==��=!T=V�=E�=�3=l� =�r =_ =�_�<��<���<h�<NL�<z��<���<���<"+�<Z`�<q��<j��<��<�)�<�X�<���<��<���<�<�.�<�T�<�x�<l��<��<s��<���<R�<z)�<d?�<�R�<�c�<hr�<O~�<s��<׍�<M��<ˑ�<#��<d��<a��< t�<-d�<�P�<�9�<I�<� �<���<n��<:��<�_�<�-�<���<"��<�|�<x9�<���<`��<�T�<}��<��<�G�<X��<_~�<�<>��<&/�<���<:�<0��<.4�<��< �<���<��<�_�<Ií<�#�<@��<�٨<�/�<���<�ң<��<�i�<[��<V��<�8�<�x�<߶�<��<s,�<Zd�<���<ώ<�<3�<�c�<ђ�<���<��<��<"E�<��|<4y<��u<��q<�,n</j<��f<$c<w_<��[<HX<uT<��P<�$M<�~I<#�E<�9B<��><�:<nd7<�3<�:0<,�,<G)<i�%<�"<��<<��<4<��<�c<�
<Y�<W<
 <��;�	�;H��;u7�;���;A��;�m�;J�;�6�;4�;>B�;�a�;a��;�ԩ;�(�;���;��;琓;�,�;Tۈ;���;��|;�r;�h;W�^;��T;�.K;J�A;�C8;A/;�%;D�;T�;�<;�;,*�:�Z�:���:f�:	>�:7J�:���:)��:�4g:��H:��*:�:6p�9W�9��W9��8�&.�B���i�K[���������{&�"�@�;K[��iu���������/Y��c��߶���JǺ�ӺG>�۠�^��������l��������� �N�&���,��2� �8�s�>���D�ɺJ�b�P�k�V��x\��_b�6Eh��)n��t���y����a܂�[΅���������㦎�����ُ�������|���  �  Br==��=T=P�=G�=�3=b� =�r =[ =�_�<��<���<i�<JL�<}��<���<���<+�<W`�<w��<\��<)��<�)�<�X�<���<��<���<�<�.�<�T�<y�<i��<��<~��<���<`�<r)�<d?�<�R�<�c�<pr�<O~�<���<э�<H��<�<-��<g��<V��<t�<$d�<�P�<�9�<G�<� �<���<o��<,��<�_�<�-�< ��<��<�|�<�9�<���<[��<�T�<���<��<�G�<\��<Y~�<�<7��<1/�<���<:�<3��<*4�<��<��<��<!��<�_�<Rí<}#�<7��<�٨<�/�<���<�ң<��<�i�<e��<D��<�8�<�x�<޶�<��<n,�<]d�<}��<ώ<��<�3�<�c�<Œ�<���<��<��< E�<��|<4y<��u<�q<�,n<Lj<k�f<&$c<w_<��[<RX<�tT<�P<$M<�~I<*�E<�9B<��><�:<�d7<��3<�:0<�,<F)<j�%<�"<��<�<��<�3<�<�c<�
<c�<�V<=
 <���;~	�;'��;�7�;���;D��;�m�;�I�;�6�;4�;BB�;�a�;S��;�ԩ;�(�;���;��;�;-�;Tۈ;;��|;��r;Ȓh;��^;��T;[.K;~�A;�C8;�/;��%;/�;)�;�<;�;B)�:>[�:&��:�f�:�=�:J�:���:���:$4g:��H:y�*:�:~q�9EX�9c�W9R��8a.�����i�!Y��ū�g���z&���@��I[�uiu���������Y�����R����IǺ��Ӻ3>�ڠ캛������0��H��9�����
� �x�&���,�Z�2���8��>�^�D���J���P���V��x\�-_b�BEh�u)n��t�z�y����t܂�!΅�����B���즎�Ϛ��ŏ������o|���  �  Lr==��=#T=S�=D�=�3=c� =�r =^ =�_�<��<���<Z�<TL�<n��<���<���<+�<X`�<k��<]��<��<�)�<�X�<���<��<���< �<�.�<�T�<y�<o��<��<���<���<\�<�)�<Z?�<�R�<�c�<qr�<V~�<s��<؍�<P��<ɑ�<$��<g��<U��<�s�<*d�<�P�<�9�<B�<� �<���<g��<3��<�_�<�-�<���<��<�|�<z9�<���<a��<�T�<}��<��<�G�<Z��<a~�< �<G��<//�<���<:�<8��<44�<��<�<��<.��<�_�<Jí<�#�<<��<�٨<�/�<���<�ң<��<�i�<f��<L��<�8�<�x�<Ҷ�<��<r,�<Vd�<���<�Ύ<��<�3�<�c�<̒�<���<��<��<0E�<��|<4y<��u<r�q<�,n<Ej<q�f<!$c<w_<��[<VX<
uT<�P<�$M<�~I<(�E<�9B<��><�:<}d7<��3<�:0<)�,<;)<r�%<�"<��<<x�<4<�<�c<�
<K�<�V<%
 <��;�	�;V��;x7�;���;���;�m�;J�;�6�;!4�;^B�;�a�;`��;�ԩ;�(�;ώ�;��;;-�;pۈ;���;��|;��r; �h;X�^;��T;L.K;2�A;�C8;F/;��%;�;��;k<;Ι;�)�:�Z�:���:nf�:S=�:J�:ƈ�:���:�4g:��H:��*::�r�9�W�9��W9���8�-�h���xi�
X�����$���{&���@��J[��gu�꫇�����Y�����󶺺�JǺ��Ӻ�>���캉�����������	�����	� �W�&���,�!�2�=�8��>�~�D�غJ���P�H�V��x\��_b��Dh��)n��t�b�y����1܂�.΅�����K�������ښ�����������|���  �  Mr==��=T=O�=E�=�3=n� =�r =` =�_�<���<���<W�<WL�<g��<���<���<+�<Y`�<f��<r��<��<�)�<�X�<���<��<���< �<�.�<�T�<y�<{��<��<w��<��<M�<�)�<c?�<�R�<�c�<hr�<Y~�<t��<ߍ�<?��<ʑ�<$��<l��<_��<�s�<1d�<�P�<�9�<=�<� �<���<_��<6��<�_�<�-�<���<��<}�<z9�<���<R��<�T�<���<��<�G�<S��<n~�<�<R��<#/�<̶�<:�</��<A4�<��<�<�<,��<�_�<Qí<�#�<.��<�٨<�/�<���<�ң<��<�i�<Q��<S��<�8�<�x�<Ѷ�<��<j,�<Od�<���<�Ύ<�<�3�<�c�<Ȓ�<���<��<��<6E�<��|<%4y<��u<��q<�,n<)j<��f<$c<w_<��[<\X<uT<��P<�$M<�~I<5�E<�9B<��><�:<{d7<�3<�:0</�,<0)<X�%<�"<��<<i�<4<��<}c<�
<A�<!W<
 <��;Z	�;,��;�7�;���;���;qm�;PJ�;�6�;P4�;>B�;�a�;���;�ԩ;)�;�;��;萓;�,�;}ۈ;���;��|;m�r;
�h;Z�^;��T;�.K;��A;	D8;� /;��%;��;�;�<;��;�)�:�Y�:���:f�:�=�:�J�:���:C��:�2g:I�H:�*:�:�p�9�U�9�W9��8_�-�4	��Mi��X���ṑ���{&���@��L[�(hu��������qY����������JǺe�Ӻ�>���v���_�������������� ���&��,���2�[�8�j�>���D�ѺJ���P�אV��x\��_b��Dh�,*n�wt�6�y����'܂�g΅�K�������������������n����|���  �  Lr==��=T=Q�=F�=�3=d� =�r =X =�_�<��<���<U�<LL�<i��<���<���<!+�<N`�<e��<]��<��<�)�<�X�<���<��<���<"�<�.�<�T�<�x�<r��<���<��<��<\�<�)�<a?�<�R�<�c�<wr�<W~�<~��<ݍ�<E��<Ǒ�<&��<Z��<T��<�s�<#d�<�P�<�9�<;�<� �<���<^��<2��<�_�<�-�<���<��<�|�<{9�<���<\��<�T�<���<��<�G�<d��<e~�<�<N��<1/�<˶�<:�<:��<74�<��<�<��<3��<�_�<Ví<�#�<9��<�٨<�/�<���<�ң<��<�i�<[��<J��<�8�<�x�<̶�<��<k,�<Zd�<x��<�Ύ<��<{3�<�c�<ɒ�<���<��<��<3E�<��|<24y<��u<��q< -n<Bj<��f<$c<$w_<��[<FX< uT<�P<�$M<�~I<3�E<�9B<��><�:<hd7<��3<�:0<�,<B)<[�%<�"<|�<�<m�<4<��<�c<�
<?�<�V<
 <��;�	�;2��;�7�;���;���;�m�;GJ�;�6�;,4�;gB�;�a�;���;�ԩ;)�;뎞;��;��;)-�;tۈ;ڛ�;��|;��r;�h;d�^;3�T;E.K;ЧA;�C8;G/;��%;��;��;O<;��;�)�:�Z�:��:|e�:+=�:fI�:ӈ�:���:$4g:2�H:�*:4:dt�9Z�9�W9��8��-�����i�gW��f�����Y|&�z�@��I[�Egu�����ь��OY�����ն���JǺ��Ӻ$?຦�캒�����������7��3��4� ���&���,���2�R�8���>���D�κJ���P���V��x\�Q_b��Dh�y)n�Ct���y����%܂�5΅�i���Y�����������ݏ��b���r|���  �  Er==��=%T=Q�=B�=�3=c� =�r =W =�_�<���<���<[�<JL�<r��<���<���<+�<L`�<w��<Z��<*��<�)�<�X�<���<��<���<�<�.�<�T�<y�<r��<���<���<���<c�<)�<r?�<�R�<�c�<nr�<O~�<y��<֍�<Y��<���<,��<b��<[��<t�<!d�<�P�<�9�<@�<� �<���<f��<#��<�_�<�-�<���<!��<�|�<�9�<���<j��<�T�<���<��<�G�<Y��<d~�<�<E��<6/�<���<:�<=��<64�<.��<�<��<(��<�_�<Pí<�#�<@��<�٨<�/�<���<�ң<��<�i�<Y��<?��<�8�<�x�<ж�<��<^,�<Sd�<v��<ώ<��<�3�<�c�<ƒ�<���<��<��<%E�<��|<4y<��u<��q<�,n<Wj<v�f<.$c<w_<��[<tX<uT<�P<�$M<�~I< �E<�9B<��><�:<�d7<��3<�:0<�,<3)<H�%<�"<��<�<~�<�3<��<qc<�
<c�<�V<<
 <��;�	�;V��;x7�;���;V��;�m�;J�;7�;,4�;eB�;�a�;b��;թ;�(�;+��;��;쐓;-�;Sۈ;ě�;��|;@�r;��h;��^;z�T;{.K;H�A;�C8;+/;H�%;��;��;n<;��;�(�:zZ�:���:7f�:�=�:�I�:v��:��:�5g:��H:��*:|:r�9)W�9��W9��8Y�-�����$i�X���������x&���@��J[��hu�ͫ��,���'Y��n�������IǺ��Ӻ >�x��3���!��U�����8����� ���&���,���2���8���>�\�D��J���P��V��x\��_b�Eh��)n��t���y�q��N܂�΅�����2���˦��������������~|���  �  Lr==��= T=L�=C�=�3=b� =�r =Y =�_�<���<���<L�<GL�<^��<���<���<+�<J`�<g��<X��<#��<�)�<�X�<���<��<���<"�<�.�<�T�<y�<p��<��<���<
��<d�<|)�<l?�<�R�<�c�<xr�<_~�<���<֍�<H��<���<(��<]��<Q��<�s�<)d�<�P�<�9�<8�<� �<���<Y��</��<�_�<�-�<���<��<�|�<�9�<���<[��<�T�<���<���<�G�<`��<k~�<�<B��<5/�<Ѷ�<#:�<7��<44�<'��<
�<��<5��<�_�<Wí<�#�<5��<�٨<�/�<���<�ң<��<�i�<T��<H��<�8�<�x�<Ŷ�<��<g,�<Ud�<{��<�Ύ<��<�3�<�c�<���<���<��<��<3E�<��|<%4y<��u<��q<�,n<_j<��f<<$c<w_<��[<jX<uT<�P<�$M<�~I<+�E<�9B<y�><�:<�d7<��3<�:0<�,<<)<S�%<�"<k�<�<V�<4<��<�c<�
<B�<�V<.
 <��;d	�;>��;�7�;���;���;�m�;J�;�6�; 4�;KB�;�a�;���;	թ;�(�;��;��;��;.-�;�ۈ;;��|;��r;��h;w�^;M�T;(.K;��A;�C8;/;��%;��;��;:<;Z�;o)�:/Z�:���:Ge�:=�:uI�:B��:P��:4g:F�H:��*:�:u�9�X�9�W9ʺ�8.�v����i��U��0��9���y&��@��I[�gu�Ъ��Ì��eY��&��h���JǺ�Ӻ�>��캊���H����9��g��j��� ���&���,�c�2�b�8��>���D��J�ܦP���V��x\�&_b��Dh�~)n�wt��y����T܂��ͅ�X������Ҧ�������������w|���  �  �s=�=��=oV=��=4�=.7=�� =^v =� =�h�<���<���<M�<X�<ԑ�<���<��<�9�<�o�<Ǥ�<���<�<�<�<�l�<F��<���<c��<��<ZG�<bn�<���<&��<���<P��<��<Y1�<�J�<�a�<Hv�<���<.��<?��<���<��<���<`��<׻�<=��<W��<���<F��<��<�l�<SS�<�5�<w�<��<���<%��<|f�<t0�<8��<���<ct�<�,�<���<A��<+;�<���<\��<� �<a��<�M�<�ݾ<�h�<��<kr�<��<�j�<��<�R�<���<�*�<쐯<t�<TR�<���<��<bZ�<���<g��<�E�<���<mԞ<��<�X�<>��<|ӗ<��<�E�<|�<���<s�<��<�D�<Bs�<���<�̅<2��<�"�<]L�<��|<�;y<�u<��q<�*n<�yj<��f<�c<�g_<�[<%	X<�[T<7�P<�M<n[I<g�E<�B<9m><n�:<k07<Ė3< 0<2m,<��(<�R%<�!<�I<��<#S<��<bq<	<j�	<�I<��<8H�;ض�;�2�;���;	W�;���; ��;
��;�X�;}A�;�;�;�F�;hc�;ّ�;�Ѩ;{$�;܈�;y��;숒;�$�;�҇;���;��z;��p;��f;�\;�R;�/I;��?;]O6;Y-;��#;��;]$;�j	;+� ;��:���:/g�:��:��:�%�:"x�:��:ca:�(C:�H%:��:i�9sD�9�"D9�ܥ8�'鷙7��1z�-���W�鹚���0*��D�n�^���x�C����Ѣ��y��=��O�Ⱥ պil�O��
	���!��7	��H��S�Z�[!�.X'��P-�[E3�'79��$?��E���J���P�+�V�h�\�p�b�lh�rLn�h+t�z�x��j䂻eԅ�?Ĉ�������җ��ъ��7~��s���  �  �s=�=��=tV=��=-�=.7=�� =\v =� =�h�<���<���<R�<X�<ב�<���<��<�9�<�o�<���<���<&�<~<�<�l�<P��<���<n��<��<`G�<en�<���<��<���<N��<��<a1�<�J�<�a�<Xv�<���<6��<F��<���<��<���<N��<ٻ�<2��<?��<���<<��<��<m�<]S�<�5�<}�<%��<���<1��<uf�<w0�<$��<y��<gt�<�,�<���<F��<3;�<���<a��<� �<p��<�M�<qݾ<�h�<��<gr�<��<�j�<��<�R�<���<�*�<���<}�<^R�<���<��<jZ�<䫥<W��<�E�<���<Ԟ<��<�X�<>��<�ӗ<��<�E�<|�<���<s�<��<�D�<7s�<���<�̅<:��<�"�<`L�<��|<�;y<��u<��q<�*n<�yj<��f<�c<�g_<�[<5	X<�[T<C�P<�M<�[I<w�E<�B< m><S�:<k07<��3< 0<*m,<�(<�R%<�!<�I<��<*S<��<�q<	<m�	<�I<��<QH�;���;�2�;���;/W�;���;���;$��;�X�;�A�;�;�;�F�;cc�;���;�Ѩ;/$�;ʈ�;���;��;�$�;Ӈ;���;��z;��p;�f;��\;��R;�.I;��?;O6;�-;��#;)�;�$;�j	;h� ;g��:���:�f�:��:c�:)%�:^x�:-�:Jca:s)C:xI%:��:��9�F�9*D9�ۥ8Kw鷜4�W6z�@�����ӝ��0*�2�D���^���x�kB�����nТ��y�����ٔȺa	պem�$�����9!��7	��H��S��Y��Z!��W'�xP-��E3�(79��%?�%E�I�J�+�P���V�-�\�/�b��kh�9Ln�+t��
z�����䂻Gԅ��Ĉ� ���F����������@~��s���  �  �s=�=��=sV=��=1�=77=�� =dv =� =�h�<���<���<X�<X�<ۑ�<���<��<�9�<�o�<ɤ�<���<6�<�<�<�l�<J��<���<e��<��<^G�<[n�<���<��<���<T��<��<n1�<�J�<�a�<Sv�<���</��<:��<���<��<���<N��<��<<��<F��<��<8��<��<�l�<US�<�5�<x�<!��<���<4��<rf�<�0�<-��<���<vt�<�,�<���<>��<&;�<���<W��<� �<i��<�M�<sݾ<�h�<��<kr�<��<�j�<��<�R�<���<�*�<퐯<k�<WR�<���<��<zZ�<ꫥ<d��<�E�<���<�Ԟ<��<�X�<=��<�ӗ<��<�E�<|�<���<��<��<�D�<As�<���<�̅<0��<�"�<RL�<��|<�;y<�u<��q<�*n<�yj<��f<�c<�g_<��[<8	X<�[T<@�P<lM<q[I<b�E<�B<$m><a�:<�07<��3<8 0<,m,<
�(<�R%<��!<�I<��<2S<��<�q<	<x�	< J<��<�H�;���;�2�;���;�V�;���;׷�;��;wX�;�A�;�;�;�F�;zc�;���;,Ҩ;:$�;ƈ�;���;݈�;�$�;�҇;���;v�z;Șp;�f;j�\;�R;./I;Q�?;�N6;�-;��#;��;o$;�j	;L� ;ۧ�:���:�f�:�:��:�%�:Ry�:�:�ca:q(C:�G%:�:R�9�C�9�&D9sܥ8�m�.��6z�1���S��]���0*�X�D�J�^��x�C������Т��y�����ϓȺ�պ�lẉ��	��+!�8	��H��S��Y�[!��W'�yP-��E3��69��%?��E���J�%�P���V�|�\�q�b�Ylh�@Ln��+t��
z�����䂻ԅ��Ĉ�ϴ��#�����������g~��s���  �  �s=�=��=pV=��=2�=-7=�� =\v =� =�h�<���<���<[�<
X�<ۑ�<���<��<�9�<�o�<���<���<�<�<�<�l�<J��<���<i��<��<_G�<bn�<���<!��<���<H��<��<S1�<�J�<�a�<Mv�<���<6��<B��<���<��<���<_��<ջ�<5��<J��<���<G��<���<m�<YS�<�5�<��<$��<���<6��<�f�<z0�<,��<��<_t�<�,�<���<C��<0;�<���<d��<� �<f��<�M�<zݾ<�h�<��<br�<��<�j�<��<�R�<���<�*�<���<v�<YR�<���<��<]Z�<<^��<�E�<���<|Ԟ<��<�X�<D��<�ӗ<��<�E�<%|�<���<s�<��<�D�<?s�<���<�̅<:��<�"�<[L�<��|<�;y<�u<��q<�*n<�yj<��f<�c<�g_<��[<	X<�[T<D�P<�M<y[I<w�E<�B<4m><f�:<e07<��3< 0<7m,<�(<�R%<�!<�I<��<2S<��<�q<	<o�	<�I<��<%H�;ɶ�;3�;���;!W�;���;��;��;�X�;^A�;�;�;�F�;Lc�;���;�Ѩ;T$�;���;���;���;�$�;�҇;���;��z;r�p;��f;ޛ\;��R;N/I;ĭ?;gO6;�-;��#;�;�$;k	;g� ;]��:���:�g�:%�:��:�%�:�w�:E�:�ba: )C:0I%:n�:{�99E�9n%D9Sԥ8R�x;�H6z�S�����h��2*���D���^��x�}B������Т��y�������Ⱥ�պ�l���Z��N!��7	��H�S��Y��Z!��W'�HP-�TE3�+79�b%?�)E��J���P�5�V�)�\�<�b�lh�0Ln��+t�z����}䂻tԅ�}Ĉ�!���,�������䊔�C~��s���  �  �s=�=µ=qV=��=3�=.7=�� =\v =� =�h�<���<���<T�<X�<֑�<���<��<�9�<�o�<¤�<���<�<�<�<�l�<M��<���<]��<��<JG�<hn�<���<��<���<G��<��<N1�<�J�<�a�<Wv�<���<'��<;��<���<��<���<`��<׻�<>��<U��<���<L��<���<m�<YS�<�5�<��<"��<���<-��<�f�<z0�<6��<���<`t�<�,�<���<H��<&;�<���<T��<� �<n��<�M�<yݾ<�h�<��<ar�<��<�j�<��<�R�<���<�*�<鐯<u�<]R�<���<��<`Z�<���<c��<�E�<���<xԞ<��<�X�<F��<�ӗ<��<�E�<|�<���<t�<��<�D�<>s�<���<�̅<>��<�"�<VL�<��|<�;y<�u<�q<�*n<�yj<��f<�c<�g_<�[<	X<�[T< �P<{M<_[I<{�E<�B<+m><i�:<i07<Ė3< 0<Dm,<�(<�R%<�!<�I<��<)S<��<~q<	<|�	<�I<��<;H�;׶�;�2�;���;$W�;���;��;��;�X�;ZA�;�;�;�F�;Ic�;ʑ�;�Ѩ;I$�;���;���;ڈ�;$�;�҇;���;��z;N�p;��f;�\;(�R;�/I;ʭ?;�O6;�-;��#;�;�$;/k	;X� ;���:o��:�g�:0�:��:C&�:�w�:��:�aa:�)C:�G%:g�:��9�B�9�)D9IΥ8HS�d=��4z����� �鹃��}2*�܍D�2�^��x�/C�����{Т�pz��X��h�Ⱥ�պ�lằ��c��t!��7	��H�sS��Y��Z!��W'��P-�E3�!79��$?�E��J���P�4�V��\���b�?lh��Ln��+t��
z����䂻�ԅ�TĈ�:���7������ߊ��?~��Ns���  �  �s=�=��=sV=��=2�=37=�� =dv =� =�h�<���<���<a�<X�<��<���<��<�9�<�o�<Ȥ�<���<.�<�<�<�l�<N��<���<e��<��<SG�<Yn�<���<��<���<G��<��<^1�<�J�<�a�<Pv�<}��<1��<B��<���<��<���<N��<��<9��<H��<	��<<��<���<m�<_S�<�5�<��<*��<���<?��<rf�<�0�<+��<���<mt�<�,�<���<B��<#;�<���<[��<� �<c��<�M�<gݾ<�h�<��<\r�<��<�j�<��<�R�<���<�*�<�<l�<[R�<���<��<rZ�<뫥<b��<�E�<���<�Ԟ<��<�X�<L��<�ӗ<��<�E�<#|�<���<��<��<�D�<@s�<���<�̅<2��<�"�<[L�<��|<�;y<��u<s�q<�*n<�yj<��f<�c<}g_<շ[</	X<�[T<2�P<�M<m[I<c�E<�B<"m><d�:<|07<��3<7 0<4m,<�(<�R%<�!<�I<�<CS<��<�q<
	<��	<�I<��<yH�;���;�2�;���;�V�;���;��;��;rX�;�A�;F;�;�F�;Ic�;}��;�Ѩ;
$�;���;���;ǈ�;�$�;�҇;���;��z;��p;�f;4�\;��R;=/I;.�?;O6;
-;�#;:�;�$;Qk	;�� ;���:���:�f�:��:��:�%�:�x�:��:Xca:)C:�G%:'�:|�9vB�9$D9�ҥ8���6��;z����������y1*�͏D�F�^���x��B������Т��y��K��O�Ⱥ�պ�l�w��>	��� ��7	�FH�BS�iY��Z!�sW'�XP-��E3��69�j%?��E��J�,�P���V�g�\�w�b�lh�_Ln��+t��
z�@���䂻Wԅ��Ĉ����Y���?�������v~��*s���  �  �s=�=��=sV=��=0�=67=�� =hv =� =�h�<���<���<l�<X�<��<���<��<�9�<�o�<Ф�<���<5�<<�<�l�<G��<���<j��<��<^G�<Jn�<���<��<���<G��<��<Z1�<�J�<�a�<Dv�<���<-��<2��<���<��<»�<P��<��<?��<N��<��<=��<��<m�<cS�<�5�<��<1��<���<Q��<wf�<�0�<2��<���<qt�<�,�<���<8��<.;�<���<T��<� �<U��<�M�<[ݾ<�h�<��<]r�<��<�j�<��<�R�<���<�*�<�<r�<SR�<ɭ�<��<wZ�<쫥<j��<�E�<���<�Ԟ<��<�X�<B��<�ӗ<��<�E�<8|�<���<��<��<�D�<?s�<���<�̅<+��<�"�<HL�<��|<�;y<�u<��q<�*n<�yj<w�f<�c<gg_<�[<-	X<j[T<A�P<[M<{[I<[�E<�B<)m><]�:<�07<��3<G 0<0m,<3�(<S%<	�!<�I<��<[S<��<�q<$	<z�	<J<��<�H�;���;#3�;���;W�;���;ŷ�; ��;8X�;�A�;X;�;}F�;Lc�;k��;�Ѩ;�#�;舝;l��;Ո�;�$�;�҇;���;C�z;�p; �f;K�\;/�R;p/I;i�?;O6;�-;��#;_�;%;Tk	;�� ; ��:���:�f�:7�:^�:
&�:y�:Y�:�da:�'C:I%:�:��9D�9�D9n�82�鷫8��<z�e��� �鹹��v/*�ؑD��^�f�x��B����Ѣ��x�������Ⱥ�պ-l�p��}��l ��7	��G��S�Y��Z!�pW'��O-�E3�k69�c%?��E��J��P���V���\�/�b��lh�HLn�5,t�z�����䂻bԅ��Ĉ��������"��������~��s���  �  �s=�=��=qV=��=0�=37=�� =cv =� =�h�<���<���<m�<X�<��<���<��<�9�<�o�<Ϥ�<���<+�<�<�<�l�<B��<���<b��<��<XG�<Jn�<���<��<���<>��<��<O1�<�J�<�a�<9v�<}��<%��<1��<���<��<���<Y��<ܻ�<A��<Z��<��<L��<��<	m�<gS�<�5�<��<5��<���<?��<�f�<�0�<;��<���<gt�<�,�<���<<��<);�<~��<L��<� �<M��<�M�<aݾ<�h�<��<Ur�<��<�j�<��<�R�<���<�*�<鐯<o�<OR�<���<��<kZ�<���<k��<�E�<���<�Ԟ<��<�X�<H��<�ӗ<��<�E�</|�<���<�<��<�D�<<s�<���<�̅<.��<�"�<JL�<��|<�;y<׋u<y�q<�*n<�yj<��f<�c<qg_<ڷ[<	X<p[T<2�P<aM<l[I<c�E<�B<+m><`�:<�07<Ŗ3<3 0<Im,</�(<�R%<�!<�I<�<bS<��<�q<3	<��	<J<��<nH�;���;�2�;~��;
W�;���;���;��;9X�;_A�;b;�;xF�;'c�;���;�Ѩ;�#�;���;A��;Ɉ�;z$�;�҇;���;j�z;��p;k�f;�\;@�R;�/I;#�?;�O6;%-;�#;��; %;ck	;�� ;Ũ�:���:�g�:��:��:o&�:sx�:��:Lca:O(C:zH%:h�:��9VB�9�D92ӥ8@���<��;z��������2*�ۑD��^��x�"C��H��NѢ��y�������Ⱥ�պl������� ��7	��G�^S�Y��Z!��W'��O-�E3��69��$?��E�"�J���P��V���\�d�b��lh��Ln�,t�oz�+���䂻�ԅ��Ĉ�C���q���3�������~��*s���  �  �s=�=��=rV=��=7�=07=�� =^v =� =�h�<���<���<e�<%X�<��<���<��<�9�<�o�<ä�<���<%�<�<�<�l�<Q��<���<^��<��<HG�<Xn�<���<��<���<5��<��<E1�<�J�<�a�<Gv�<y��<(��<A��<���<��<���<[��<��<:��<S��<��<\��<���< m�<cS�<�5�<��<*��<���<9��<�f�<�0�<3��<���<kt�<�,�<���<K��<;�<���<U��<� �<\��<�M�<cݾ<�h�<��<Nr�<��<�j�<��<�R�<���<�*�<됯<g�<`R�<���<��<gZ�<���<`��<�E�<���<�Ԟ<��<�X�<]��<�ӗ<��<�E�<%|�<���<v�<��<�D�<Hs�<���<�̅<9��<�"�<\L�<��|<�;y<�u<Z�q<�*n<oyj<��f<�c<ug_<��[<	X<{[T<�P<�M<W[I<p�E<�B<%m><y�:<q07<��3<! 0<gm,<�(<S%<,�!<�I<.�<DS<��<�q<3	<��	<�I<��<UH�;��;�2�;���;�V�;���;���;��;rX�;?A�;>;�;rF�;c�;y��;�Ѩ;$�;]��;|��;���;�$�;�҇;a��;��z;M�p;�f;T�\;�R;�/I;��?;P6;�-;��#;b�;N%;�k	;�� ;���:8��:�h�:��:t�:&�:�x�:(�:�aa:?*C:�F%:پ:+�9�@�9o!D9���8Ƥ�(A��=z�������ş��3*�͏D���^�5�x��B�����6Т�Tz��_���Ⱥ0պ�l������ �7	�LH��R�*Y�eZ!�W'�IP-��D3�79��$?�E���J���P�/�V�0�\�ԋb�lh��Ln�,t�Az�����䂻�ԅ��Ĉ�x���g���j�������~��bs���  �  �s=�=��=uV=��=6�=67=�� =hv =� =�h�<���<���<j�<X�<��<���<��<�9�<�o�<Ԥ�<���<3�<�<�<�l�<T��<���<[��<��<FG�<Pn�<���<��<���<8��<��<G1�<�J�<�a�<Hv�<t��<"��<2��<|��<��<���<U��<��<E��<`��<��<U��<���< m�<eS�<�5�<��<-��<���<>��<�f�<�0�<B��<���<rt�<�,�<���<F��<;�<}��<K��<� �<]��<�M�<_ݾ<�h�<��<Nr�<��<�j�<��<�R�<���<�*�<㐯<g�<`R�<���<��<tZ�<���<p��<�E�<���<�Ԟ<��<�X�<T��<�ӗ<��<�E�<&|�<���<��<��<�D�<Hs�<���<�̅<6��<�"�<LL�<��|<�;y<�u<_�q<�*n<{yj<��f<�c<ig_<��[<	X<l[T<�P<^M<P[I<j�E<�B<"m><v�:<�07<Ŗ3<I 0<am,<�(<S%<1�!<�I<�<RS<��<�q<'	<��	<J<��<�H�;۶�;�2�;Ƚ�;W�;���;ŷ�;��;VX�;bA�;=;�;fF�;c�;q��;�Ѩ;�#�;x��;��;���;q$�;�҇;T��;��z;��p;T�f;e�\;a�R;	0I;w�?;�O6;-;��#;p�;L%;�k	;�� ;��:���:%h�:m�:i�:�&�:4y�:{�:�ba:�)C:hF%:a�:��9@�9�!D9�ȥ8V��M@��>z�����i�����2*���D�׽^�¸x�oC�����,Т�z������Ⱥ�պ�kẨ����� ��6	�H��R�Y�RZ!��V'�BP-��D3�g69��$?��E���J��P���V�I�\���b��lh��Ln�O,t�+z�����䂻�ԅ��Ĉ�_�������i���는��~��as���  �  �s=�=��=qV=��=1�=47=�� =gv =� =�h�<���<���<|�<X�<��<���<��<�9�<�o�<Ҥ�<���<+�<�<�<�l�<C��<���<g��<��<YG�<Fn�<���< ��<���<2��<��<E1�<�J�<�a�<<v�<~��<'��<1��<���<
��<���<S��<ۻ�<:��<P��<��<R��<	��<m�<yS�<�5�<��<F��<���<H��<�f�<�0�<3��<���<gt�<�,�<���<5��<1;�<��<M��<� �<N��<�M�<Vݾ<�h�<��<Er�<��<�j�<��<�R�<���<�*�<됯<t�<OR�<���<��<kZ�<�<k��<�E�<���<�Ԟ<��<�X�<L��<�ӗ<��<�E�<6|�<���<��<��<�D�<=s�<���<�̅<-��<�"�<DL�<��|<�;y<Ջu<d�q<w*n<yyj<u�f<�c<Vg_<·[<		X<h[T<3�P<OM<|[I<_�E<�B<.m><a�:<�07<��3<E 0<Om,<:�(<S%<:�!<�I<�<�S<��<�q<:	<��	<J<��<rH�;���;3�;���;W�;���;���;��;+X�;KA�;3;�;QF�;�b�;Q��;�Ѩ;�#�;���;N��;Ј�;�$�;�҇;ȓ�;@�z;p;>�f;�\;�R;�/I;^�?;�O6;e-;��#;�;�%;�k	;�� ;���:.��:2h�:!�:x�:�%�:�x�:��:�ca:�'C:�I%:��:n�9SC�9�D9�ȥ8��鷱A��Cz�㣳�Q�鹠��A3*�~�D�~�^�n�x��B�����=Ѣ�xy������ȺGպl������ �(7	�HG�?S��X�Z!��V'��O-�E3�o69�(%?��E��J���P��V���\�%�b��lh�xLn�5,t�tz�|���䂻�ԅ��Ĉ�g�������d�������~��'s���  �  �s=�=��=pV=��=6�=87=�� =gv =� =�h�<���<���<q�<X�<���<���<��<�9�<�o�<Ӥ�<���<4�<�<�<�l�<B��<���<Y��<��<GG�<Hn�<���<��<���<2��<��<E1�<�J�<�a�<>v�<r��<��<)��<���<��<���<[��<��<E��<[��<��<Z��<��<m�<nS�<�5�<��<9��<���<F��<�f�<�0�<=��<���<vt�<�,�<���<6��<!;�<u��<C��<� �<P��<�M�<_ݾ<�h�<��<Ir�<��<�j�<��<�R�<���<�*�<ᐯ<g�<NR�<���<��<sZ�< ��<p��<�E�<���<�Ԟ<��<�X�<S��<�ӗ<��<�E�<5|�<���<��<��<�D�<Js�<���<�̅<*��<�"�<AL�<��|<�;y<ڋu<c�q<�*n<pyj<s�f<�c<kg_<÷[<	X<c[T<�P<MM<\[I<U�E<�B<2m><w�:<�07<ɖ3<H 0<cm,<8�(<S%<)�!<�I<�<jS<��<�q<8	<��	<J<��<�H�;ٶ�;
3�;���;�V�;���;���;��;8X�;JA�;J;�;zF�;�b�;Z��;�Ѩ;�#�;{��;[��;���;W$�;�҇;���;M�z;��p;~�f;��\;g�R;�/I;��?;P6;X-;n�#;��;i%;�k	;� ;Z��:��:�h�:��:�:�&�:yy�:��:Gca:�'C:�G%:e�:�
�9N?�9�D9�ĥ8Q�鷾@��Az�����
�鹹��c3*��D�½^�.�x��C�����JѢ��y�����#�Ⱥ{պ�k�y��t��� �?7	��G�S��X�WZ!�W'��O-��D3�_69��$?��E���J���P�#�V���\���b��lh��Ln�V,t�bz����䂻�ԅ��Ĉ�~���z���a�������~��cs���  �  �s=�=��=uV=��=2�=37=�� =ev =� =�h�<ĥ�<���<n�<,X�<��<���<��<�9�<�o�<̤�<���<+�<�<�<�l�<S��<���<`��<��<GG�<Pn�<���<���<���<(��<��<@1�<�J�<�a�<>v�<o��<,��<<��<���< ��<���<Q��<��<<��<\��<��<S��<��<(m�<oS�<�5�<��<6��<���<F��<�f�<�0�<;��<���<nt�<�,�<���<J��<;�<���<U��<� �<U��<�M�<\ݾ<�h�<��<@r�<��<�j�<��<�R�<���<�*�<됯<h�<`R�<���<��<lZ�<���<h��<�E�<���<�Ԟ<��<�X�<b��<�ӗ<��<�E�<,|�<���<��<��<�D�<Bs�<���<�̅<:��<�"�<]L�<��|<�;y<͋u<?�q<�*n<jyj<{�f<�c<ig_<��[<�X<h[T<!�P<�M<V[I<r�E<�B<m><e�:<07<ʖ3<= 0<fm,<(�(<0S%<:�!<�I<<�<[S<��<�q<$	<��	<J<��<rH�;���;�2�;Ƚ�;W�;���; ��;��;WX�;&A�;;�;PF�;�b�;T��;{Ѩ;�#�;7��;X��;���;�$�;�҇;l��;��z;��p;.�f;R�\;"�R;�/I;Y�?;�O6;K-;�#;��;�%;�k	; � ;���:��:�g�::�:��:6&�:�x�:
�:*ca:I*C:�F%:*�:n�9�>�9'D9�8���zD��Cz�,���	��B���4*���D���^��x��B�����*Т��y�������Ⱥ�պAlẾ��R��_ ��6	��G��R��X�Z!��V'�P-��D3��69��$?��E���J��P���V�)�\�ҋb�lh��Ln�X,t��z����䂻�ԅ��Ĉ�����������������~��Ks���  �  �s=�=��=pV=��=6�=87=�� =gv =� =�h�<���<���<q�<X�<���<���<��<�9�<�o�<Ӥ�<���<4�<�<�<�l�<B��<���<Y��<��<GG�<Hn�<���<��<���<2��<��<E1�<�J�<�a�<>v�<r��<��<)��<���<��<���<[��<��<E��<[��<��<Z��<��<m�<nS�<�5�<��<9��<���<F��<�f�<�0�<=��<���<vt�<�,�<���<6��<!;�<u��<C��<� �<P��<�M�<_ݾ<�h�<��<Ir�<��<�j�<��<�R�<���<�*�<ᐯ<g�<NR�<���<��<sZ�< ��<p��<�E�<���<�Ԟ<��<�X�<S��<�ӗ<��<�E�<5|�<���<��<��<�D�<Js�<���<�̅<*��<�"�<AL�<��|<�;y<ڋu<c�q<�*n<pyj<s�f<�c<kg_<÷[<	X<c[T<�P<MM<\[I<U�E<�B<2m><w�:<�07<ɖ3<H 0<cm,<8�(<S%<)�!<�I<�<jS<��<�q<8	<��	<J<��<�H�;ٶ�;
3�;���;�V�;���;���;��;8X�;JA�;J;�;zF�;�b�;Z��;�Ѩ;�#�;{��;[��;���;W$�;�҇;���;M�z;��p;~�f;��\;g�R;�/I;��?;P6;X-;n�#;��;i%;�k	;� ;Z��:��:�h�:��:�:�&�:yy�:��:Gca:�'C:�G%:e�:�
�9N?�9�D9�ĥ8Q�鷾@��Az�����
�鹹��c3*��D�½^�.�x��C�����JѢ��y�����#�Ⱥ{պ�k�y��t��� �?7	��G�S��X�WZ!�W'��O-��D3�_69��$?��E���J���P�#�V���\���b��lh��Ln�V,t�bz����䂻�ԅ��Ĉ�~���z���a�������~��cs���  �  �s=�=��=qV=��=1�=47=�� =gv =� =�h�<���<���<|�<X�<��<���<��<�9�<�o�<Ҥ�<���<+�<�<�<�l�<C��<���<g��<��<YG�<Fn�<���< ��<���<2��<��<E1�<�J�<�a�<<v�<~��<'��<1��<���<
��<���<S��<ۻ�<:��<P��<��<R��<	��<m�<yS�<�5�<��<F��<���<H��<�f�<�0�<3��<���<gt�<�,�<���<5��<1;�<��<M��<� �<N��<�M�<Vݾ<�h�<��<Er�<��<�j�<��<�R�<���<�*�<됯<t�<OR�<���<��<kZ�<�<k��<�E�<���<�Ԟ<��<�X�<L��<�ӗ<��<�E�<6|�<���<��<��<�D�<=s�<���<�̅<-��<�"�<DL�<��|<�;y<Ջu<d�q<w*n<yyj<u�f<�c<Vg_<·[<		X<h[T<3�P<OM<|[I<_�E<�B<.m><a�:<�07<��3<E 0<Om,<:�(<S%<:�!<�I<�<�S<��<�q<:	<��	<J<��<rH�;���;3�;���;W�;���;���;��;+X�;KA�;3;�;QF�;�b�;Q��;�Ѩ;�#�;���;N��;Ј�;�$�;�҇;ȓ�;@�z;p;>�f;�\;�R;�/I;^�?;�O6;e-;��#;�;�%;�k	;�� ;���:.��:2h�:!�:x�:�%�:�x�:��:�ca:�'C:�I%:��:n�9SC�9�D9�ȥ8��鷱A��Cz�㣳�Q�鹠��A3*�~�D�~�^�n�x��B�����=Ѣ�xy������ȺGպl������ �(7	�HG�?S��X�Z!��V'��O-�E3�o69�(%?��E��J���P��V���\�%�b��lh�xLn�5,t�tz�|���䂻�ԅ��Ĉ�g�������d�������~��'s���  �  �s=�=��=uV=��=6�=67=�� =hv =� =�h�<���<���<j�<X�<��<���<��<�9�<�o�<Ԥ�<���<3�<�<�<�l�<T��<���<[��<��<FG�<Pn�<���<��<���<8��<��<G1�<�J�<�a�<Hv�<t��<"��<2��<|��<��<���<U��<��<E��<`��<��<U��<���< m�<eS�<�5�<��<-��<���<>��<�f�<�0�<B��<���<rt�<�,�<���<F��<;�<}��<K��<� �<]��<�M�<_ݾ<�h�<��<Nr�<��<�j�<��<�R�<���<�*�<㐯<g�<`R�<���<��<tZ�<���<p��<�E�<���<�Ԟ<��<�X�<T��<�ӗ<��<�E�<&|�<���<��<��<�D�<Hs�<���<�̅<6��<�"�<LL�<��|<�;y<�u<_�q<�*n<{yj<��f<�c<ig_<��[<	X<l[T<�P<^M<P[I<j�E<�B<"m><v�:<�07<Ŗ3<I 0<am,<�(<S%<1�!<�I<�<RS<��<�q<'	<��	<J<��<�H�;۶�;�2�;Ƚ�;W�;���;ŷ�;��;VX�;bA�;=;�;fF�;c�;q��;�Ѩ;�#�;x��;��;���;q$�;�҇;T��;��z;��p;T�f;e�\;a�R;	0I;w�?;�O6;-;��#;p�;L%;�k	;�� ;��:���:%h�:m�:i�:�&�:4y�:{�:�ba:�)C:hF%:a�:��9@�9�!D9�ȥ8V��M@��>z�����i�����2*���D�׽^�¸x�oC�����,Т�z������Ⱥ�պ�kẨ����� ��6	�H��R�Y�RZ!��V'�BP-��D3�g69��$?��E���J��P���V�I�\���b��lh��Ln�O,t�+z�����䂻�ԅ��Ĉ�_�������i���는��~��as���  �  �s=�=��=rV=��=7�=07=�� =^v =� =�h�<���<���<e�<%X�<��<���<��<�9�<�o�<ä�<���<%�<�<�<�l�<Q��<���<^��<��<HG�<Xn�<���<��<���<5��<��<E1�<�J�<�a�<Gv�<y��<(��<A��<���<��<���<[��<��<:��<S��<��<\��<���< m�<cS�<�5�<��<*��<���<9��<�f�<�0�<3��<���<kt�<�,�<���<K��<;�<���<U��<� �<\��<�M�<cݾ<�h�<��<Nr�<��<�j�<��<�R�<���<�*�<됯<g�<`R�<���<��<gZ�<���<`��<�E�<���<�Ԟ<��<�X�<]��<�ӗ<��<�E�<%|�<���<v�<��<�D�<Hs�<���<�̅<9��<�"�<\L�<��|<�;y<�u<Z�q<�*n<oyj<��f<�c<ug_<��[<	X<{[T<�P<�M<W[I<p�E<�B<%m><y�:<q07<��3<! 0<gm,<�(<S%<,�!<�I<.�<DS<��<�q<3	<��	<�I<��<UH�;��;�2�;���;�V�;���;���;��;rX�;?A�;>;�;rF�;c�;y��;�Ѩ;$�;]��;|��;���;�$�;�҇;a��;��z;M�p;�f;T�\;�R;�/I;��?;P6;�-;��#;b�;N%;�k	;�� ;���:8��:�h�:��:t�:&�:�x�:(�:�aa:?*C:�F%:پ:+�9�@�9o!D9���8Ƥ�(A��=z�������ş��3*�͏D���^�5�x��B�����6Т�Tz��_���Ⱥ0պ�l������ �7	�LH��R�*Y�eZ!�W'�IP-��D3�79��$?�E���J���P�/�V�0�\�ԋb�lh��Ln�,t�Az�����䂻�ԅ��Ĉ�x���g���j�������~��bs���  �  �s=�=��=qV=��=0�=37=�� =cv =� =�h�<���<���<m�<X�<��<���<��<�9�<�o�<Ϥ�<���<+�<�<�<�l�<B��<���<b��<��<XG�<Jn�<���<��<���<>��<��<O1�<�J�<�a�<9v�<}��<%��<1��<���<��<���<Y��<ܻ�<A��<Z��<��<L��<��<	m�<gS�<�5�<��<5��<���<?��<�f�<�0�<;��<���<gt�<�,�<���<<��<);�<~��<L��<� �<M��<�M�<aݾ<�h�<��<Ur�<��<�j�<��<�R�<���<�*�<鐯<o�<OR�<���<��<kZ�<���<k��<�E�<���<�Ԟ<��<�X�<H��<�ӗ<��<�E�</|�<���<�<��<�D�<<s�<���<�̅<.��<�"�<JL�<��|<�;y<׋u<y�q<�*n<�yj<��f<�c<qg_<ڷ[<	X<p[T<2�P<aM<l[I<c�E<�B<+m><`�:<�07<Ŗ3<3 0<Im,</�(<�R%<�!<�I<�<bS<��<�q<3	<��	<J<��<nH�;���;�2�;~��;
W�;���;���;��;9X�;_A�;b;�;xF�;'c�;���;�Ѩ;�#�;���;A��;Ɉ�;z$�;�҇;���;j�z;��p;k�f;�\;@�R;�/I;#�?;�O6;%-;�#;��; %;ck	;�� ;Ũ�:���:�g�:��:��:o&�:sx�:��:Lca:O(C:zH%:h�:��9VB�9�D92ӥ8@���<��;z��������2*�ۑD��^��x�"C��H��NѢ��y�������Ⱥ�պl������� ��7	��G�^S�Y��Z!��W'��O-�E3��69��$?��E�"�J���P��V���\�d�b��lh��Ln�,t�oz�+���䂻�ԅ��Ĉ�C���q���3�������~��*s���  �  �s=�=��=sV=��=0�=67=�� =hv =� =�h�<���<���<l�<X�<��<���<��<�9�<�o�<Ф�<���<5�<<�<�l�<G��<���<j��<��<^G�<Jn�<���<��<���<G��<��<Z1�<�J�<�a�<Dv�<���<-��<2��<���<��<»�<P��<��<?��<N��<��<=��<��<m�<cS�<�5�<��<1��<���<Q��<wf�<�0�<2��<���<qt�<�,�<���<8��<.;�<���<T��<� �<U��<�M�<[ݾ<�h�<��<]r�<��<�j�<��<�R�<���<�*�<�<r�<SR�<ɭ�<��<wZ�<쫥<j��<�E�<���<�Ԟ<��<�X�<B��<�ӗ<��<�E�<8|�<���<��<��<�D�<?s�<���<�̅<+��<�"�<HL�<��|<�;y<�u<��q<�*n<�yj<w�f<�c<gg_<�[<-	X<j[T<A�P<[M<{[I<[�E<�B<)m><]�:<�07<��3<G 0<0m,<3�(<S%<	�!<�I<��<[S<��<�q<$	<z�	<J<��<�H�;���;#3�;���;W�;���;ŷ�; ��;8X�;�A�;X;�;}F�;Lc�;k��;�Ѩ;�#�;舝;l��;Ո�;�$�;�҇;���;C�z;�p; �f;K�\;/�R;p/I;i�?;O6;�-;��#;_�;%;Tk	;�� ; ��:���:�f�:7�:^�:
&�:y�:Y�:�da:�'C:I%:�:��9D�9�D9n�82�鷫8��<z�e��� �鹹��v/*�ؑD��^�f�x��B����Ѣ��x�������Ⱥ�պ-l�p��}��l ��7	��G��S�Y��Z!�pW'��O-�E3�k69�c%?��E��J��P���V���\�/�b��lh�HLn�5,t�z�����䂻bԅ��Ĉ��������"��������~��s���  �  �s=�=��=sV=��=2�=37=�� =dv =� =�h�<���<���<a�<X�<��<���<��<�9�<�o�<Ȥ�<���<.�<�<�<�l�<N��<���<e��<��<SG�<Yn�<���<��<���<G��<��<^1�<�J�<�a�<Pv�<}��<1��<B��<���<��<���<N��<��<9��<H��<	��<<��<���<m�<_S�<�5�<��<*��<���<?��<rf�<�0�<+��<���<mt�<�,�<���<B��<#;�<���<[��<� �<c��<�M�<gݾ<�h�<��<\r�<��<�j�<��<�R�<���<�*�<�<l�<[R�<���<��<rZ�<뫥<b��<�E�<���<�Ԟ<��<�X�<L��<�ӗ<��<�E�<#|�<���<��<��<�D�<@s�<���<�̅<2��<�"�<[L�<��|<�;y<��u<s�q<�*n<�yj<��f<�c<}g_<շ[</	X<�[T<2�P<�M<m[I<c�E<�B<"m><d�:<|07<��3<7 0<4m,<�(<�R%<�!<�I<�<CS<��<�q<
	<��	<�I<��<yH�;���;�2�;���;�V�;���;��;��;rX�;�A�;F;�;�F�;Ic�;}��;�Ѩ;
$�;���;���;ǈ�;�$�;�҇;���;��z;��p;�f;4�\;��R;=/I;.�?;O6;
-;�#;:�;�$;Qk	;�� ;���:���:�f�:��:��:�%�:�x�:��:Xca:)C:�G%:'�:|�9vB�9$D9�ҥ8���6��;z����������y1*�͏D�F�^���x��B������Т��y��K��O�Ⱥ�պ�l�w��>	��� ��7	�FH�BS�iY��Z!�sW'�XP-��E3��69�j%?��E��J�,�P���V�g�\�w�b�lh�_Ln��+t��
z�@���䂻Wԅ��Ĉ����Y���?�������v~��*s���  �  �s=�=µ=qV=��=3�=.7=�� =\v =� =�h�<���<���<T�<X�<֑�<���<��<�9�<�o�<¤�<���<�<�<�<�l�<M��<���<]��<��<JG�<hn�<���<��<���<G��<��<N1�<�J�<�a�<Wv�<���<'��<;��<���<��<���<`��<׻�<>��<U��<���<L��<���<m�<YS�<�5�<��<"��<���<-��<�f�<z0�<6��<���<`t�<�,�<���<H��<&;�<���<T��<� �<n��<�M�<yݾ<�h�<��<ar�<��<�j�<��<�R�<���<�*�<鐯<u�<]R�<���<��<`Z�<���<c��<�E�<���<xԞ<��<�X�<F��<�ӗ<��<�E�<|�<���<t�<��<�D�<>s�<���<�̅<>��<�"�<VL�<��|<�;y<�u<�q<�*n<�yj<��f<�c<�g_<�[<	X<�[T< �P<{M<_[I<{�E<�B<+m><i�:<i07<Ė3< 0<Dm,<�(<�R%<�!<�I<��<)S<��<~q<	<|�	<�I<��<;H�;׶�;�2�;���;$W�;���;��;��;�X�;ZA�;�;�;�F�;Ic�;ʑ�;�Ѩ;I$�;���;���;ڈ�;$�;�҇;���;��z;N�p;��f;�\;(�R;�/I;ʭ?;�O6;�-;��#;�;�$;/k	;X� ;���:o��:�g�:0�:��:C&�:�w�:��:�aa:�)C:�G%:g�:��9�B�9�)D9IΥ8HS�d=��4z����� �鹃��}2*�܍D�2�^��x�/C�����{Т�pz��X��h�Ⱥ�պ�lằ��c��t!��7	��H�sS��Y��Z!��W'��P-�E3�!79��$?�E��J���P�4�V��\���b�?lh��Ln��+t��
z����䂻�ԅ�TĈ�:���7������ߊ��?~��Ns���  �  �s=�=��=pV=��=2�=-7=�� =\v =� =�h�<���<���<[�<
X�<ۑ�<���<��<�9�<�o�<���<���<�<�<�<�l�<J��<���<i��<��<_G�<bn�<���<!��<���<H��<��<S1�<�J�<�a�<Mv�<���<6��<B��<���<��<���<_��<ջ�<5��<J��<���<G��<���<m�<YS�<�5�<��<$��<���<6��<�f�<z0�<,��<��<_t�<�,�<���<C��<0;�<���<d��<� �<f��<�M�<zݾ<�h�<��<br�<��<�j�<��<�R�<���<�*�<���<v�<YR�<���<��<]Z�<<^��<�E�<���<|Ԟ<��<�X�<D��<�ӗ<��<�E�<%|�<���<s�<��<�D�<?s�<���<�̅<:��<�"�<[L�<��|<�;y<�u<��q<�*n<�yj<��f<�c<�g_<��[<	X<�[T<D�P<�M<y[I<w�E<�B<4m><f�:<e07<��3< 0<7m,<�(<�R%<�!<�I<��<2S<��<�q<	<o�	<�I<��<%H�;ɶ�;3�;���;!W�;���;��;��;�X�;^A�;�;�;�F�;Lc�;���;�Ѩ;T$�;���;���;���;�$�;�҇;���;��z;r�p;��f;ޛ\;��R;N/I;ĭ?;gO6;�-;��#;�;�$;k	;g� ;]��:���:�g�:%�:��:�%�:�w�:E�:�ba: )C:0I%:n�:{�99E�9n%D9Sԥ8R�x;�H6z�S�����h��2*���D���^��x�}B������Т��y�������Ⱥ�պ�l���Z��N!��7	��H�S��Y��Z!��W'�HP-�TE3�+79�b%?�)E��J���P�5�V�)�\�<�b�lh�0Ln��+t�z����}䂻tԅ�}Ĉ�!���,�������䊔�C~��s���  �  �s=�=��=sV=��=1�=77=�� =dv =� =�h�<���<���<X�<X�<ۑ�<���<��<�9�<�o�<ɤ�<���<6�<�<�<�l�<J��<���<e��<��<^G�<[n�<���<��<���<T��<��<n1�<�J�<�a�<Sv�<���</��<:��<���<��<���<N��<��<<��<F��<��<8��<��<�l�<US�<�5�<x�<!��<���<4��<rf�<�0�<-��<���<vt�<�,�<���<>��<&;�<���<W��<� �<i��<�M�<sݾ<�h�<��<kr�<��<�j�<��<�R�<���<�*�<퐯<k�<WR�<���<��<zZ�<ꫥ<d��<�E�<���<�Ԟ<��<�X�<=��<�ӗ<��<�E�<|�<���<��<��<�D�<As�<���<�̅<0��<�"�<RL�<��|<�;y<�u<��q<�*n<�yj<��f<�c<�g_<��[<8	X<�[T<@�P<lM<q[I<b�E<�B<$m><a�:<�07<��3<8 0<,m,<
�(<�R%<��!<�I<��<2S<��<�q<	<x�	< J<��<�H�;���;�2�;���;�V�;���;׷�;��;wX�;�A�;�;�;�F�;zc�;���;,Ҩ;:$�;ƈ�;���;݈�;�$�;�҇;���;v�z;Șp;�f;j�\;�R;./I;Q�?;�N6;�-;��#;��;o$;�j	;L� ;ۧ�:���:�f�:�:��:�%�:Ry�:�:�ca:q(C:�G%:�:R�9�C�9�&D9sܥ8�m�.��6z�1���S��]���0*�X�D�J�^��x�C������Т��y�����ϓȺ�պ�lẉ��	��+!�8	��H��S��Y�[!��W'�yP-��E3��69��%?��E���J�%�P���V�|�\�q�b�Ylh�@Ln��+t��
z�����䂻ԅ��Ĉ�ϴ��#�����������g~��s���  �  �s=�=��=tV=��=-�=.7=�� =\v =� =�h�<���<���<R�<X�<ב�<���<��<�9�<�o�<���<���<&�<~<�<�l�<P��<���<n��<��<`G�<en�<���<��<���<N��<��<a1�<�J�<�a�<Xv�<���<6��<F��<���<��<���<N��<ٻ�<2��<?��<���<<��<��<m�<]S�<�5�<}�<%��<���<1��<uf�<w0�<$��<y��<gt�<�,�<���<F��<3;�<���<a��<� �<p��<�M�<qݾ<�h�<��<gr�<��<�j�<��<�R�<���<�*�<���<}�<^R�<���<��<jZ�<䫥<W��<�E�<���<Ԟ<��<�X�<>��<�ӗ<��<�E�<|�<���<s�<��<�D�<7s�<���<�̅<:��<�"�<`L�<��|<�;y<��u<��q<�*n<�yj<��f<�c<�g_<�[<5	X<�[T<C�P<�M<�[I<w�E<�B< m><S�:<k07<��3< 0<*m,<�(<�R%<�!<�I<��<*S<��<�q<	<m�	<�I<��<QH�;���;�2�;���;/W�;���;���;$��;�X�;�A�;�;�;�F�;cc�;���;�Ѩ;/$�;ʈ�;���;��;�$�;Ӈ;���;��z;��p;�f;��\;��R;�.I;��?;O6;�-;��#;)�;�$;�j	;h� ;g��:���:�f�:��:c�:)%�:^x�:-�:Jca:s)C:xI%:��:��9�F�9*D9�ۥ8Kw鷜4�W6z�@�����ӝ��0*�2�D���^���x�kB�����nТ��y�����ٔȺa	պem�$�����9!��7	��H��S��Y��Z!��W'�xP-��E3�(79��%?�%E�I�J�+�P���V�-�\�/�b��kh�9Ln�+t��
z�����䂻Gԅ��Ĉ� ���F����������@~��s���  �  Ou=�=�=�X=��=C�=�:=�� =ez =� =r�<���<���<�(�<Rd�<��<���<{�<`I�<2��<���<���<(�<�P�<r��<"��<z��<D�<�7�<Ba�<n��<ï�<[��<��<��<�6�<@S�<�m�<���<��<R��<:��<���<��<���<���<���<X��<���<3��<��<���<N��<n��<Ԋ�<Sn�<�M�<{)�<� �<3��<<��<�m�<'4�<��<K��<l�<@ �<���<�z�<>!�<���<�_�<y��<K��<��<W��<�,�<���< ,�<?��<5�<��<���<�`�<�ů<�&�<D��<5ު<�4�<懧<�ץ<�$�<�n�<���<���<�;�<�z�<z��<�<z*�<�`�<e��<*Ȑ<0��<�(�<�V�<���<F��<�م<`�<�+�<�S�<\�|<Dy<��u<��q<R(n<�sj<e�f<�
c<W_<�[<��W<�@T<��P<�L<�5I<`�E<��A<�<><��:<9�6<�[3<��/<y+,<Ϙ(<
%<�!<��<�x<��<�<v<Ҩ<�B	<U�<F�<o�;���;-N�;r��;�g�;g�;'��;T��;�V�;�;�;W2�;&:�;�S�;��;q��;�;�p�;��;o�;f
�;���;�y�;�x;�gn;�Zd;�qZ;�P;"G;ܑ=;�94;�+;��!;��;,;{;���:���:�B�:T��:���:���:�ϛ:�6�:��y:^4[:�&=:=q:�:��9{��9_y/9�{8P.B�����%���Y��q򹈮��.�UH��_b�;4|���������f]��O����{����ɺlUֺ��⺙���*�������	�������[��(�!�=�'�ٮ-�Н3�5�9��r?�YE��<K��Q���V�]�\��b�,�h�*qn�0Kt��%z� ��;킻�څ�+Ȉ�˶������'��������v��ai���  �  Hu=�=�=�X=��=B�=�:=�� =jz =� =r�<¯�<���<�(�<bd�<���<���<��<[I�<7��<���<���<*�<yP�<���<+��<v��<B�<�7�<Sa�<m��<���<W��<��<��<�6�<AS�<�m�<���<���<Q��<9��<���<��<���<���<���<[��<���<3��<��<y��<T��<q��<֊�<bn�<�M�<�)�<� �<;��<2��<�m�<(4�<���<L��<l�<R �<���<�z�<4!�<���<�_�<u��<H��<��<[��<�,�<|��<,�<9��<0�<��<���<�`�<�ů<�&�<M��<Iު<�4�<燧<�ץ<�$�<�n�<���<���<�;�<�z�<���<�<v*�<�`�<f��<Ȑ<<��<�(�<�V�<���<Q��<�م<b�< ,�<�S�<t�|<�Cy<��u<��q<N(n<�sj<�f<�
c<W_<�[<��W<�@T<��P<e�L<�5I<Y�E<��A<=><��:<5�6<�[3<��/<l+,<̘(<)
%<�!<�<�x<��<�<�<ɨ<C	<b�<%�<o�;���;|N�;���;�g�;a�;��;���;�V�;�;�;J2�;9:�;�S�;\�;v��;��;�p�;��;o�;a
�;���;�y�;,�x;Ahn;�Zd;�qZ;�P; G;X�=;b94;�+;��!;��;�,;|{;,��:���:AC�:���:���:���:ϛ:�6�:<�y:�6[:_'=:�q:F: �9|��9w/9x�{8�?B�x��W,��^�� �9��4.�QUH��]b��5|�����Ű���\�����D|����ɺoVֺ�����K+����z�	�z�������D�!��'�̮-�*�3�։9��r?�YE��<K�<Q�B�V�Q�\�͹b���h��pn�NKt��%z� ��E킻�څ��Ȉ�䶋�����&��������v��&i���  �  Fu=�=�=�X=��=@�=�:=�� =oz =� =r�<ǯ�<���<�(�<Sd�<��<���<��<TI�<5��<��<���<<�<pP�<���<!��<r��<Q�<�7�<Wa�<b��<ǯ�<Q��<��<��<�6�<OS�<�m�<���<ޛ�<L��<=��<���<!��<���<���<���<`��<���<0��<!��<q��<W��<r��<Ҋ�<[n�<�M�<~)�<� �<;��<'��<�m�<$4�<���<U��<l�<S �<���<�z�<8!�<���<�_�<o��<N��<��<e��<�,�<���<,�<3��<7�<��<���<�`�<�ů<�&�<C��<Hު<�4�<���<�ץ<�$�<�n�<���<���<�;�<�z�<z��<�<p*�<�`�<h��<Ȑ<E��<�(�<�V�<���<M��<�م<T�<,�<�S�<��|<�Cy<��u<��q<5(n<�sj<$�f<c<W_<�[<��W<w@T<��P<]�L<�5I<C�E<��A<=><��:<S�6<�[3<��/<b+,<ɘ(<3
%<�!<��<�x<��<�<�<��<C	<s�<%�<ao�;���;xN�;p��;�g�;��;��;���;�V�;�;�;22�;*:�;�S�;~�;���;��;�p�;��;o�;r
�;���;�y�;Śx;1hn;sZd;rZ;�P;G;��=;"94;�+;��!;��;U,;"{;���:���:OC�:��:Û�:~��:Mϛ:�7�:X�y:�6[:�%=:�r:�:��90��9Rt/9��{8nSB�n��q*��[�������h.�VH�]b�.6|����ɰ��s]������|����ɺHVֺK�����+��y����	�������%��t�!���'���-�X�3���9��r?��XE��<K�\Q�r�V���\�_�b���h��pn��Kt��%z� ��v킻�څ��Ȉ�����¥��7��������v��i���  �  Hu=�=�=�X=��=>�=�:=�� =kz =� =r�<ǯ�<���<�(�<ad�<���<���<��<^I�<2��<��<���</�<tP�<z��<'��<v��<F�<�7�<Ga�<a��<ʯ�<T��<���<��<�6�<8S�<�m�<���<���<G��<8��<���<��<���<���<���<S��<���<7��<��<���<L��<y��<���<en�<�M�<�)�<� �<2��<8��<�m�<)4�<��<H��<l�<K �<���<�z�<4!�<���<�_�<p��<M��<��<O��<�,�<��<�+�<4��<8�<��<���<�`�<�ů<�&�<I��<<ު<�4�<뇧<�ץ<�$�<�n�<���<���<�;�<�z�<���<�<�*�<�`�<c��<'Ȑ<:��<�(�<�V�<���<J��<�م<X�<,�<�S�<i�|<�Cy<��u<��q<.(n<�sj<*�f<�
c<�V_<�[<��W<u@T<��P<b�L<�5I<L�E<��A<�<><��:<E�6<�[3<��/<t+,<ɘ(<3
%<�!<�<�x<��<�<�<Ϩ<�B	<o�<:�<-o�;���;PN�;���;�g�;s�;��;m��;�V�;
<�;>2�;�9�;�S�;{�;T��;��;�p�;��;�n�;_
�;���;�y�;�x;$hn;�Zd;�qZ;-�P;>G;&�=;�94;�+;	�!;�;�,;~{;���:~��:�B�:��:&��:˚�:�ϛ:�6�:(�y:�5[:�&=:�q:<:�99u/9��{8GOB�`��+��8]����̯�9.��VH�_b�'6|�����ʰ��]������H|��m�ɺ�Uֺ?�⺄���*������	�j��'�������!��'��-��3��9��r?��XE�=K�rQ�R�V���\���b���h��pn��Kt��%z� ���킻�څ��Ȉ�붋�륎�3���o����v��Gi���  �  Iu=�=�=�X=��=G�=�:=�� =gz =� =%r�<ʯ�<���<�(�<id�<��<���<��<mI�<9��<���<���<)�<�P�<{��<-��<u��<9�<�7�<Oa�<j��<���<U��<��<��<�6�<:S�<�m�<��<ڛ�<I��<9��<���<��<���<���<���<\��<���<;��<��<���<Q��<���<ڊ�<^n�<�M�<�)�<�<8��<F��<�m�<,4�<���<L��<$l�<H �<���<�z�<.!�<���<�_�<p��<;��<��<T��<�,�<|��<�+�<5��<"�<��<���<�`�<�ů<�&�<Q��<<ު<�4�<燧<�ץ<�$�<�n�<���<���<�;�<�z�<���<
�<�*�<�`�<k��<1Ȑ<3��<�(�<�V�<���<P��<�م<_�<�+�<�S�<s�|<�Cy<��u<��q<N(n<�sj<&�f<�
c<W_<�[<��W<�@T<��P<g�L<�5I<T�E<��A<=><��:<3�6<�[3<��/<�+,<ߘ(<:
%<�!<��<y<��<�<�<�<C	<d�<8�<o�;���;SN�;���;�g�;>�;��;���;�V�;�;�;C2�;$:�;�S�;{�;^��;��;�p�;��;�n�;b
�;���;zy�;K�x;hn;�Zd;�qZ;�P;cG;�=;
:4;�+;Z�!;��;r,;g{;M��:"��:C�:���:<��:��:Rϛ:7�:��y:�5[:+(=:�p:�:q�9�9 u/9�m{8�?B�}���*���]���򹢯��.��UH�I^b�|5|�������\������O{����ɺ�Uֺu��,��*��{���	�������.����!���'���-���3��9��r?�YE��<K�GQ�U�V�i�\��b���h��pn��Kt�&z�7 ��D킻�څ��Ȉ�	�������G��������v��2i���  �  Cu=�=�=�X=��=E�=�:=�� =qz =� =&r�<ʯ�<���<�(�<id�< ��<���<��<dI�<C��<��<���<:�<xP�<}��<$��<r��<J�<�7�<Ja�<^��<���<K��<��<��<�6�<=S�<�m�<��<՛�<C��<5��<���<��<���<���<���<k��<���<;��<*��<���<Y��<���<��<in�<�M�<�)�< �<?��<;��<�m�</4�<���<\��<l�<K �<���<�z�<3!�<���<�_�<g��<@��<��<S��<�,�<n��<�+�<)��<)�<��<���<�`�<�ů<�&�<E��<?ު<�4�<���<�ץ<�$�<�n�<���<���<�;�<�z�<���<�<�*�<�`�<p��<+Ȑ<K��<�(�<�V�<���<H��<�م<W�<,�<�S�<m�|<�Cy<��u<��q<-(n<�sj<�f<�
c<�V_<ԣ[<��W<j@T<��P<Q�L<�5I<J�E<��A<�<><��:<J�6<�[3<�/<�+,<��(<9
%<�!<�<y<��<�<�<ܨ<!C	<��<5�<\o�;���;\N�;~��;�g�;��;Ծ�;}��;�V�;�;�;2�;:�;�S�;D�;h��;��;�p�;r�;�n�;R
�;���;�y�;	�x;hn;jZd;erZ;�P;fG;ϒ=;�94;�+;K�!;-�;�,;�{;��:���:�C�:G��:z��:=��:>ϛ:8�:t�y:�5[:'=:�q:T:��9���9�p/98z{8{`B�����.��"a��I����.��VH��^b��6|���������F]������b|����ɺVֺȪ�8���*��P���	�#����������!���'��-�͝3�W�9��r?��XE�{<K��Q�u�V���\���b�Еh��pn��Kt�&z�C ���킻�څ��Ȉ����Х��^��������v��>i���  �  =u=�=ܷ=�X=��=A�=�:=�� =sz =� =.r�<ѯ�<���<)�<dd�<��<���<��<iI�<?��<��<���<>�<pP�<���<%��<n��<C�<�7�<Pa�<O��<���<A��< ��<��<~6�<9S�<�m�<���<ț�<G��<0��<r��<��<���<���<���<g��<���<4��<*��<���<e��<|��<��<ln�<�M�<�)�<� �<L��<9��<�m�<+4�<���<Y��<l�<Z �<���<�z�<'!�<���<�_�<Y��<C��<z�<O��<�,�<n��<�+�<��<*�<�<���<�`�<�ů<�&�<?��<Mު<�4�<���<�ץ<�$�<�n�<���<���<�;�<�z�<���<!�<�*�<�`�<x��<%Ȑ<M��<�(�<�V�<���<L��<�م<J�<
,�<�S�<m�|<�Cy<��u<��q<(n<�sj<��f<�
c<�V_<ɣ[<��W<[@T<��P<8�L<�5I<3�E<��A<=><��:<Z�6<�[3<�/<z+,<�(<H
%<�!<*�<�x<��<�<�<�<C	<��<'�<oo�;���;�N�;���;�g�;j�;���;���;vV�;�;�;�1�;�9�;�S�;&�;\��;��;�p�;A�;�n�;B
�;O��;�y�;~�x;�hn;\Zd;JrZ;�P;3G;Ւ=;�94;W+;&�!;{�;�,;�{;���:���:cD�:0��:���:���:Lϛ:�7�:נy:�7[:�$=:�q:�:�9���9j/9��{8�yB����0���`��u�q���.�YH�^b��8|�,������]�������|��w�ɺuVֺĪ�Y�*��ت�$�	������w����!���'�:�-���3�L�9��r?��XE��<K�aQ���V��\�{�b�@�h��pn��Kt�B&z�M ���킻�څ� Ɉ����󥎻t�������w��0i���  �  Bu=�=�=�X=��=F�=�:=�� =qz =� =-r�<د�<���<)�<od�<��<���<��<pI�<A��<��<���<;�<~P�<y��<$��<v��<=�<�7�<Oa�<T��<���<A��<���<��<�6�<.S�<�m�<��<Ǜ�<H��<0��<x��<��<���<���<���<e��<���<A��<$��<���<c��<���<��<ln�<N�<�)�<�<I��<G��<�m�<34�<��<X��<l�<J �<���<�z�<(!�<���<�_�<Y��<5��<��<E��<�,�<i��<�+�< ��<�<���<���<�`�<�ů<�&�<@��<;ު<�4�<���<�ץ<�$�<�n�<���<���<�;�<�z�<���< �<�*�<�`�<v��<3Ȑ<F��<�(�<�V�<���<G��<�م<R�<,�<�S�<f�|<�Cy<u�u<p�q<"(n<�sj<�f<�
c<�V_<��[<��W<f@T<��P<J�L<�5I<B�E<��A<�<><��:<]�6<�[3<�/<�+,<�(<V
%<	�!<*�<y<�<�<�<��<C	<��<E�<fo�;���;QN�;���;�g�;U�;ľ�;���;�V�;�;�;�1�;�9�;{S�;7�;3��;��;�p�;@�;�n�;E
�;h��;�y�;��x;-hn;�Zd;?rZ;\�P;�G;��=;-:4;I+;��!;��;�,;�{;���:e��::D�:��:0��:���:�ϛ:�7�:��y:�5[:�%=:r::��9ؕ�9ij/9gf{8�lB�o���/��)b������M.��XH�^b��7|�|񊺠����]�������{����ɺ�Uֺ���w���)����̺	����������Z�!�b�'�L�-���3���9��r?�|XE��<K��Q�b�V���\���b���h�qn��Kt�r&z�} ���킻*ۅ��Ȉ�9���񥎻����΅��w��Di���  �  Cu=�=�=�X=��=H�=�:=�� =sz =� =,r�<ޯ�<���<)�<yd�<��<���<��<qI�<K��<��<���<+�<�P�<|��<.��<m��<9�<�7�<7a�<[��<���<B��<���<��<~6�< S�<�m�<���<ӛ�<7��<'��<y��<
��<���<���<���<b��<���<J��<(��<���<\��<���<��<{n�<N�<�)�<�<B��<P��<�m�<;4�<���<Q��<$l�<G �<���<�z�<)!�<���<�_�<d��<.��<��<6��<�,�<\��<�+�<"��<�<���<���<�`�<�ů<�&�<O��<<ު<�4�<釧<�ץ<�$�<�n�<���<���<�;�<�z�<���<&�<�*�<�`�<s��<?Ȑ<K��<�(�<�V�<���<P��<�م<^�<�+�<�S�<G�|<�Cy<��u<l�q<"(n<lsj<�f<�
c<�V_<��[<��W<e@T<z�P<N�L<�5I<P�E<��A<=><Ù:<7�6<\3<	�/<�+,<�(<d
%<�!</�<'y<��<;�<�<��<2C	<��<R�<(o�;���;aN�;���;�g�;F�;о�;3��;�V�;�;�; 2�;�9�;GS�;+�;���;��;yp�;r�;�n�;!
�;m��;ky�;F�x;hn;�Zd;(rZ;��P;�G;ǒ=;z:4;+;��!;��;c-;L|;��:`��:�C�:���:x��:���:kϛ:y7�:أy:�5[:(=:�o:3:�
�92��97p/9�W{8JhB�b�c1��e��򹹱�8 .�yWH�ab�_7|��񊺉����\������={��h�ɺ_UֺI������)����@�	����Z��N��-�!��'�c�-�&�3�Y�9�r?�YE�n<K�HQ�_�V�n�\�)�b��h��qn�Lt�>&z�� ���킻`ۅ��Ȉ�n�����������ȅ��w���i���  �  Cu=�=۷=�X=��=G�=�:=�� =pz =� =>r�<��<���<)�<{d�<��<���<��<{I�<F��<��<���<9�<P�<|��<'��<`��<@�<�7�<<a�<Q��<���<;��<���<��<{6�<%S�<�m�<ۅ�<ě�<3��<)��<}��<��<���<���<���<h��<���<E��<"��<���<o��<���<��<|n�<N�<�)�<�<T��<N��<�m�<84�<��<Y��<l�<I �<���<�z�<.!�<���<�_�<U��<'��<y�<<��<�,�<e��<�+�<��<�<�<���<�`�<�ů<�&�<E��<=ު<�4�<���<�ץ<�$�<�n�<���<��<�;�<�z�<���<,�<�*�<�`�<���<6Ȑ<D��<�(�<�V�<���<K��<�م<L�<�+�<�S�<T�|<�Cy<f�u<f�q<(n<ysj<��f<�
c<�V_<��[<p�W<Q@T<��P<P�L<�5I</�E<��A<�<><��:<R�6<\3<��/<�+,<�(<j
%<�!<>�<,y<�<�<�<�<)C	<��<P�<_o�;���;cN�;���;�g�;c�;���;L��;�V�;z;�;�1�;�9�;pS�;�;��;��;hp�;6�;�n�;+
�;|��;wy�;՚x;hn;�Zd;ZrZ;\�P;�G;��=;L:4;�+;��!;[�;l-;F|;���:���:�D�:���:*��:֛�:�ϛ:�7�:^�y:�5[:g&=:�o:�:�	�9���9�h/95L{8NzB�v�=1���b������� .��XH��`b�8|��-��� ]�������{����ɺTUֺd��3��N)�������	����S������!��'���-�o�3���9�Kr?��XE�n<K�nQ�j�V���\��b��h�Kqn�LLt��&z�� ���킻Dۅ�Ɉ�O��������������0w��mi���  �  =u=�=۷=�X=��=D�=�:=�� =wz =� =8r�<��<���<)�<yd�<$��<���<��<xI�<I��<��<���<B�<{P�<{��<(��<j��<B�<�7�<Ia�<C��<���<7��<���<��<l6�<S�<�m�<���<���<:��<'��<u��<��<���<���<���<j��<��<F��<1��<���<n��<���<���<�n�<N�<�)�<�<T��<M��<�m�<:4�<
��<]��<l�<R �<���<�z�<&!�<���<�_�<E��</��<o�<3��<x,�<Z��<�+�<��<�<ኴ<���<�`�<�ů<�&�<B��<<ު<�4�<���<�ץ<�$�<�n�<���<��<�;�<�z�<���<;�<�*�<�`�<���<7Ȑ<S��<�(�<�V�<���<E��<�م<I�<,�<�S�<\�|<�Cy<V�u<k�q<�'n<nsj<׾f<�
c<�V_<��[<k�W<D@T<��P<5�L<�5I</�E<��A<�<><��:<i�6<\3<�/<�+,<�(<g
%<�!<b�<'y<1�<"�<�<�</C	<��<M�<�o�;���;]N�;���;�g�;m�;���;~��;LV�;�;�;�1�;�9�;MS�;�~�;���;]�;|p�;��;�n�;#
�;]��;�y�;��x;zhn;�Zd;irZ;��P;�G;�=;N:4;�+;��!;��;�-;c|;���:���:�D�:y��:朻:��:FЛ:>8�:��y:�6[:�%=:[q:�:	�9���9�`/9�[{8��B���v4���e��� 򹻳��.��ZH�_b��8|�-�g���R]������$|��&�ɺ\Uֺ������b)�������	���Q�����1�!�3�'�ۭ-�j�3��9�]r?�IXE��<K��Q�&�V��\���b�D�h�-qn�MLt��&z�� ���킻Zۅ�EɈ�h���O����������Kw��Ui���  �  =u=�=޷=�X=��=I�=�:=�� =uz =� =4r�<��<���<)�<pd�<��<���<��<xI�<R��<��<���<5�<�P�<���<-��<j��<8�<�7�<?a�<H��<���<3��<���<��<|6�<"S�<�m�<���<���<9��<$��<q��<
��<���<���<���<h��<���<H��<.��<���<i��<���<���<xn�<N�<�)�<�<N��<R��<�m�<94�<��<X��<l�<Q �<���<�z�<"!�<���<�_�<O��<.��<o�<6��<�,�<a��<�+�<��<�<芴<���<�`�<�ů<�&�<I��<@ު<�4�<�<�ץ<�$�<�n�<���<���<�;�<�z�<���<*�<�*�<a�<~��<CȐ<O��<�(�<�V�<���<M��<�م<Q�<�+�<�S�<H�|<�Cy<b�u<g�q< (n<wsj<��f<�
c<�V_<��[<q�W<M@T<��P<9�L<�5I<:�E<��A< =><ș:<J�6<
\3<�/<�+,<��(<r
%<&�!<@�<y<�<:�<�<�<AC	<��<U�<Ro�;���;rN�;���;�g�;D�;���;X��;bV�;�;�;�1�;�9�;nS�;$�;��;c�;zp�;&�;�n�;
�;O��;ly�;њx;|hn;�Zd;[rZ;C�P;�G;��=;�:4;|+;�!;��;Q-;&|;i��:y��:�D�:���:���:�:�ϛ:�7�:�y:�6[:j&=:�o:m:�	�9M��9,f/9x[{8��B�D� 1���c��c�����.�	ZH��_b�z8|��񊺗����\��x���K{����ɺGUֺF�⺋��Q)�����R�	�������*����!���'��-�	�3�9�9�6r?��XE�h<K�XQ��V���\�#�b�B�h�yqn�4Lt��&z�� ���킻Hۅ�Ɉ�P���7�����������8w��}i���  �  Eu=�=�=�X=��=K�=�:=�� =mz =� =6r�<��<���<)�<�d�<��<���<��<}I�<V��<
��<���</�<�P�<q��<$��<j��<;�<�7�<4a�<U��<���<0��<���<��<n6�<S�<�m�<م�<Ǜ�<0��<$��<���<	��<���<���<���<h��<���<S��<!��<���<m��<���<��<�n�<$N�<�)�<�<Q��<W��<�m�<A4�<��<U��<l�<= �<���<�z�<.!�<���<�_�<Y��<'��<k�<-��<x,�<R��<�+�<��<�<�<���<�`�<�ů<�&�<D��<0ު<�4�<퇧<�ץ<�$�<�n�<���<���<�;�<�z�<���<5�<�*�<a�<���<DȐ<>��<�(�<�V�<���<E��<�م<X�<�+�<�S�<9�|<�Cy<j�u<Z�q<(n<[sj<׾f<�
c<�V_<��[<v�W<S@T<n�P<V�L<�5I<B�E<��A<�<><Й:<C�6<$\3<��/<�+,<�(<r
%<�!<N�<ey<�<B�<�<�<JC	<��<n�<7o�;���;7N�;���;�g�;Q�;���;+��;�V�;�;�;�1�;�9�;7S�;�~�;ؼ�;Y�;`p�;C�;�n�;
�;���;jy�;�x;�gn;�Zd;\rZ;m�P;4G;��=;�:4;�+;5�!;��;�-;�|;��:���:�D�:%��:q��:j��:WЛ:�7�:o�y:n4[:�&=:�o:�:q	�9J��9k/9;M{8ݓB�d
�w4��ng��a�U��� .�sXH��ab�W8|�[񊺷���(]��u���d{��$�ɺTֺh��k��
)�����	�	�����������!��'���-��3���9��q?��XE�><K��Q���V���\�$�b���h��qn�HLt��&z�� ���킻�ۅ�FɈ�����)���˕��셔�+w���i���  �  =u=�=޷=�X=��=I�=�:=�� =uz =� =4r�<��<���<)�<pd�<��<���<��<xI�<R��<��<���<5�<�P�<���<-��<j��<8�<�7�<?a�<H��<���<3��<���<��<|6�<"S�<�m�<���<���<9��<$��<q��<
��<���<���<���<h��<���<H��<.��<���<i��<���<���<xn�<N�<�)�<�<N��<R��<�m�<94�<��<X��<l�<Q �<���<�z�<"!�<���<�_�<O��<.��<o�<6��<�,�<a��<�+�<��<�<芴<���<�`�<�ů<�&�<I��<@ު<�4�<�<�ץ<�$�<�n�<���<���<�;�<�z�<���<*�<�*�<a�<~��<CȐ<O��<�(�<�V�<���<M��<�م<Q�<�+�<�S�<H�|<�Cy<b�u<g�q< (n<wsj<��f<�
c<�V_<��[<q�W<M@T<��P<9�L<�5I<:�E<��A< =><ș:<J�6<
\3<�/<�+,<��(<r
%<&�!<@�<y<�<:�<�<�<AC	<��<U�<Ro�;���;rN�;���;�g�;D�;���;X��;bV�;�;�;�1�;�9�;nS�;$�;��;c�;zp�;&�;�n�;
�;O��;ly�;њx;|hn;�Zd;[rZ;C�P;�G;��=;�:4;|+;�!;��;Q-;&|;i��:y��:�D�:���:���:�:�ϛ:�7�:�y:�6[:j&=:�o:m:�	�9M��9,f/9x[{8��B�D� 1���c��c�����.�	ZH��_b�z8|��񊺗����\��x���K{����ɺGUֺF�⺋��Q)�����R�	�������*����!���'��-�	�3�9�9�6r?��XE�h<K�XQ��V���\�#�b�B�h�yqn�4Lt��&z�� ���킻Hۅ�Ɉ�P���7�����������8w��}i���  �  =u=�=۷=�X=��=D�=�:=�� =wz =� =8r�<��<���<)�<yd�<$��<���<��<xI�<I��<��<���<B�<{P�<{��<(��<j��<B�<�7�<Ia�<C��<���<7��<���<��<l6�<S�<�m�<���<���<:��<'��<u��<��<���<���<���<j��<��<F��<1��<���<n��<���<���<�n�<N�<�)�<�<T��<M��<�m�<:4�<
��<]��<l�<R �<���<�z�<&!�<���<�_�<E��</��<o�<3��<x,�<Z��<�+�<��<�<ኴ<���<�`�<�ů<�&�<B��<<ު<�4�<���<�ץ<�$�<�n�<���<��<�;�<�z�<���<;�<�*�<�`�<���<7Ȑ<S��<�(�<�V�<���<E��<�م<I�<,�<�S�<\�|<�Cy<V�u<k�q<�'n<nsj<׾f<�
c<�V_<��[<k�W<D@T<��P<5�L<�5I</�E<��A<�<><��:<i�6<\3<�/<�+,<�(<g
%<�!<b�<'y<1�<"�<�<�</C	<��<M�<�o�;���;]N�;���;�g�;m�;���;~��;LV�;�;�;�1�;�9�;MS�;�~�;���;]�;|p�;��;�n�;#
�;]��;�y�;��x;zhn;�Zd;irZ;��P;�G;�=;N:4;�+;��!;��;�-;c|;���:���:�D�:y��:朻:��:FЛ:>8�:��y:�6[:�%=:[q:�:	�9���9�`/9�[{8��B���v4���e��� 򹻳��.��ZH�_b��8|�-�g���R]������$|��&�ɺ\Uֺ������b)�������	���Q�����1�!�3�'�ۭ-�j�3��9�]r?�IXE��<K��Q�&�V��\���b�D�h�-qn�MLt��&z�� ���킻Zۅ�EɈ�h���O����������Kw��Ui���  �  Cu=�=۷=�X=��=G�=�:=�� =pz =� =>r�<��<���<)�<{d�<��<���<��<{I�<F��<��<���<9�<P�<|��<'��<`��<@�<�7�<<a�<Q��<���<;��<���<��<{6�<%S�<�m�<ۅ�<ě�<3��<)��<}��<��<���<���<���<h��<���<E��<"��<���<o��<���<��<|n�<N�<�)�<�<T��<N��<�m�<84�<��<Y��<l�<I �<���<�z�<.!�<���<�_�<U��<'��<y�<<��<�,�<e��<�+�<��<�<�<���<�`�<�ů<�&�<E��<=ު<�4�<���<�ץ<�$�<�n�<���<��<�;�<�z�<���<,�<�*�<�`�<���<6Ȑ<D��<�(�<�V�<���<K��<�م<L�<�+�<�S�<T�|<�Cy<f�u<f�q<(n<ysj<��f<�
c<�V_<��[<p�W<Q@T<��P<P�L<�5I</�E<��A<�<><��:<R�6<\3<��/<�+,<�(<j
%<�!<>�<,y<�<�<�<�<)C	<��<P�<_o�;���;cN�;���;�g�;c�;���;L��;�V�;z;�;�1�;�9�;pS�;�;��;��;hp�;6�;�n�;+
�;|��;wy�;Ԛx;hn;�Zd;ZrZ;\�P;�G;��=;L:4;�+;��!;[�;l-;F|;���:���:�D�:���:*��:֛�:�ϛ:�7�:^�y:�5[:g&=:�o:�:�	�9���9�h/95L{8NzB�v�=1���b������� .��XH��`b�8|��-��� ]�������{����ɺTUֺd��3��N)�������	����S������!��'���-�o�3���9�Kr?��XE�n<K�nQ�j�V���\��b��h�Kqn�LLt��&z�� ���킻Dۅ�Ɉ�O��������������0w��mi���  �  Cu=�=�=�X=��=H�=�:=�� =sz =� =,r�<ޯ�<���<)�<yd�<��<���<��<qI�<K��<��<���<+�<�P�<|��<.��<m��<9�<�7�<7a�<[��<���<B��<���<��<~6�< S�<�m�<���<ӛ�<7��<'��<y��<
��<���<���<���<b��<���<J��<(��<���<\��<���<��<{n�<N�<�)�<�<B��<P��<�m�<;4�<���<Q��<$l�<G �<���<�z�<)!�<���<�_�<d��<.��<��<6��<�,�<\��<�+�<"��<�<���<���<�`�<�ů<�&�<O��<<ު<�4�<釧<�ץ<�$�<�n�<���<���<�;�<�z�<���<&�<�*�<�`�<s��<?Ȑ<K��<�(�<�V�<���<P��<�م<^�<�+�<�S�<G�|<�Cy<��u<l�q<"(n<lsj<�f<�
c<�V_<��[<��W<e@T<z�P<N�L<�5I<P�E<��A<=><Ù:<7�6<\3<	�/<�+,<�(<d
%<�!</�<'y<��<;�<�<��<2C	<��<R�<(o�;���;aN�;���;�g�;F�;о�;3��;�V�;�;�; 2�;�9�;GS�;+�;���;��;yp�;r�;�n�;!
�;m��;ky�;F�x;hn;�Zd;(rZ;��P;�G;ǒ=;z:4;+;��!;��;c-;L|;��:`��:�C�:���:x��:���:kϛ:y7�:أy:�5[:(=:�o:3:�
�92��97p/9�W{8JhB�b�c1��e��򹹱�8 .�yWH�ab�_7|��񊺉����\������={��h�ɺ_UֺI������)����@�	����Z��N��-�!��'�c�-�&�3�Y�9�r?�YE�n<K�HQ�_�V�n�\�)�b��h��qn�Lt�>&z�� ���킻`ۅ��Ȉ�n�����������ȅ��w���i���  �  Bu=�=�=�X=��=F�=�:=�� =qz =� =-r�<د�<���<)�<od�<��<���<��<pI�<A��<��<���<;�<~P�<y��<$��<v��<=�<�7�<Oa�<T��<���<A��<���<��<�6�<.S�<�m�<��<Ǜ�<H��<0��<x��<��<���<���<���<e��<���<A��<$��<���<c��<���<��<ln�<N�<�)�<�<I��<G��<�m�<34�<��<X��<l�<J �<���<�z�<(!�<���<�_�<Y��<5��<��<E��<�,�<i��<�+�< ��<�<���<���<�`�<�ů<�&�<@��<;ު<�4�<���<�ץ<�$�<�n�<���<���<�;�<�z�<���< �<�*�<�`�<v��<3Ȑ<F��<�(�<�V�<���<G��<�م<R�<,�<�S�<f�|<�Cy<u�u<p�q<"(n<�sj<�f<�
c<�V_<��[<��W<f@T<��P<J�L<�5I<B�E<��A<�<><��:<]�6<�[3<�/<�+,<�(<V
%<	�!<*�<y<�<�<�<��<C	<��<E�<fo�;���;QN�;���;�g�;U�;ľ�;���;�V�;�;�;�1�;�9�;{S�;7�;3��;��;�p�;@�;�n�;E
�;h��;�y�;��x;-hn;�Zd;?rZ;\�P;�G;��=;-:4;I+;��!;��;�,;�{;���:e��::D�:��:0��:���:�ϛ:�7�:��y:�5[:�%=:r::��9ؕ�9ij/9gf{8�lB�o���/��)b������M.��XH�^b��7|�|񊺠����]�������{����ɺ�Uֺ���w���)����̺	����������Z�!�b�'�L�-���3���9��r?�|XE��<K��Q�b�V���\���b���h�qn��Kt�r&z�} ���킻*ۅ��Ȉ�9���񥎻����΅��w��Di���  �  =u=�=ܷ=�X=��=A�=�:=�� =sz =� =.r�<ѯ�<���<)�<dd�<��<���<��<iI�<?��<��<���<>�<pP�<���<%��<n��<C�<�7�<Pa�<O��<���<A��< ��<��<~6�<9S�<�m�<���<ț�<G��<0��<r��<��<���<���<���<g��<���<4��<*��<���<e��<|��<��<ln�<�M�<�)�<� �<L��<9��<�m�<+4�<���<Y��<l�<Z �<���<�z�<'!�<���<�_�<Y��<C��<z�<O��<�,�<n��<�+�<��<*�<�<���<�`�<�ů<�&�<?��<Mު<�4�<���<�ץ<�$�<�n�<���<���<�;�<�z�<���<!�<�*�<�`�<x��<%Ȑ<M��<�(�<�V�<���<L��<�م<J�<
,�<�S�<m�|<�Cy<��u<��q<(n<�sj<��f<�
c<�V_<ɣ[<��W<[@T<��P<8�L<�5I<3�E<��A<=><��:<Z�6<�[3<�/<z+,<�(<H
%<�!<*�<�x<��<�<�<�<C	<��<'�<oo�;���;�N�;���;�g�;j�;���;���;vV�;�;�;�1�;�9�;�S�;&�;\��;��;�p�;A�;�n�;B
�;O��;�y�;~�x;�hn;\Zd;JrZ;�P;3G;Ւ=;�94;W+;&�!;{�;�,;�{;���:���:cD�:0��:���:���:Lϛ:�7�:נy:�7[:�$=:�q:�:�9���9j/9��{8�yB����0���`��u�q���.�YH�^b��8|�,������]�������|��w�ɺuVֺĪ�Y�*��ت�$�	������w����!���'�:�-���3�L�9��r?��XE��<K�aQ���V��\�{�b�@�h��pn��Kt�B&z�M ���킻�څ� Ɉ����󥎻t�������w��0i���  �  Cu=�=�=�X=��=E�=�:=�� =qz =� =&r�<ʯ�<���<�(�<id�< ��<���<��<dI�<C��<��<���<:�<xP�<}��<$��<r��<J�<�7�<Ja�<^��<���<K��<��<��<�6�<=S�<�m�<��<՛�<C��<5��<���<��<���<���<���<k��<���<;��<*��<���<Y��<���<��<in�<�M�<�)�< �<?��<;��<�m�</4�<���<\��<l�<K �<���<�z�<3!�<���<�_�<g��<@��<��<S��<�,�<n��<�+�<)��<)�<��<���<�`�<�ů<�&�<E��<?ު<�4�<���<�ץ<�$�<�n�<���<���<�;�<�z�<���<�<�*�<�`�<p��<+Ȑ<K��<�(�<�V�<���<H��<�م<W�<,�<�S�<m�|<�Cy<��u<��q<-(n<�sj<�f<�
c<�V_<ԣ[<��W<j@T<��P<Q�L<�5I<J�E<��A<�<><��:<J�6<�[3<�/<�+,<��(<9
%<�!<�<y<��<�<�<ܨ<!C	<��<5�<\o�;���;\N�;~��;�g�;��;Ծ�;}��;�V�;�;�;2�;:�;�S�;D�;h��;��;�p�;r�;�n�;R
�;���;�y�;	�x;hn;jZd;erZ;�P;fG;ϒ=;�94;�+;K�!;-�;�,;�{;��:���:�C�:G��:z��:=��:>ϛ:8�:t�y:�5[:'=:�q:T:��9���9�p/98z{8{`B�����.��"a��I����.��VH��^b��6|���������F]������b|����ɺVֺȪ�8���*��P���	�#����������!���'��-�͝3�W�9��r?��XE�{<K��Q�u�V���\���b�Еh��pn��Kt�&z�C ���킻�څ��Ȉ����Х��^��������v��>i���  �  Iu=�=�=�X=��=G�=�:=�� =gz =� =%r�<ʯ�<���<�(�<id�<��<���<��<mI�<9��<���<���<)�<�P�<{��<-��<u��<9�<�7�<Oa�<j��<���<U��<��<��<�6�<:S�<�m�<��<ڛ�<I��<9��<���<��<���<���<���<\��<���<;��<��<���<Q��<���<ڊ�<^n�<�M�<�)�<�<8��<F��<�m�<,4�<���<L��<$l�<H �<���<�z�<.!�<���<�_�<p��<;��<��<T��<�,�<|��<�+�<5��<"�<��<���<�`�<�ů<�&�<Q��<<ު<�4�<燧<�ץ<�$�<�n�<���<���<�;�<�z�<���<
�<�*�<�`�<k��<1Ȑ<3��<�(�<�V�<���<P��<�م<_�<�+�<�S�<s�|<�Cy<��u<��q<N(n<�sj<&�f<�
c<W_<�[<��W<�@T<��P<g�L<�5I<T�E<��A<=><��:<3�6<�[3<��/<�+,<ߘ(<:
%<�!<��<y<��<�<�<�<C	<d�<8�<o�;���;SN�;���;�g�;>�;��;���;�V�;�;�;C2�;$:�;�S�;{�;^��;��;�p�;��;�n�;b
�;���;zy�;K�x;hn;�Zd;�qZ;�P;cG;�=;
:4;�+;Z�!;��;r,;g{;M��:"��:C�:���:<��:��:Rϛ:7�:��y:�5[:+(=:�p:�:q�9�9 u/9�m{8�?B�}���*���]���򹢯��.��UH�I^b�|5|�������\������O{����ɺ�Uֺu��,��*��{���	�������.����!���'���-���3��9��r?�YE��<K�GQ�U�V�i�\��b���h��pn��Kt�&z�7 ��D킻�څ��Ȉ�	�������G��������v��2i���  �  Hu=�=�=�X=��=>�=�:=�� =kz =� =r�<ǯ�<���<�(�<ad�<���<���<��<^I�<2��<��<���</�<tP�<z��<'��<v��<F�<�7�<Ga�<a��<ʯ�<T��<���<��<�6�<8S�<�m�<���<���<G��<8��<���<��<���<���<���<S��<���<7��<��<���<L��<y��<���<en�<�M�<�)�<� �<2��<8��<�m�<)4�<��<H��<l�<K �<���<�z�<4!�<���<�_�<p��<M��<��<O��<�,�<��<�+�<4��<8�<��<���<�`�<�ů<�&�<I��<<ު<�4�<뇧<�ץ<�$�<�n�<���<���<�;�<�z�<���<�<�*�<�`�<c��<'Ȑ<:��<�(�<�V�<���<J��<�م<X�<,�<�S�<i�|<�Cy<��u<��q<.(n<�sj<*�f<�
c<�V_<�[<��W<u@T<��P<b�L<�5I<L�E<��A<�<><��:<E�6<�[3<��/<t+,<ɘ(<3
%<�!<�<�x<��<�<�<Ϩ<�B	<o�<:�<-o�;���;PN�;���;�g�;s�;��;m��;�V�;
<�;>2�;�9�;�S�;{�;T��;��;�p�;��;�n�;_
�;���;�y�;�x;$hn;�Zd;�qZ;-�P;>G;&�=;�94;�+;	�!;�;�,;~{;���:~��:�B�:��:&��:˚�:�ϛ:�6�:(�y:�5[:�&=:�q:<:�99u/9��{8GOB�`��+��8]����̯�9.��VH�_b�'6|�����ʰ��]������H|��m�ɺ�Uֺ?�⺄���*������	�j��'�������!��'��-��3��9��r?��XE�=K�rQ�R�V���\���b���h��pn��Kt��%z� ���킻�څ��Ȉ�붋�륎�3���o����v��Gi���  �  Fu=�=�=�X=��=@�=�:=�� =oz =� =r�<ǯ�<���<�(�<Sd�<��<���<��<TI�<5��<��<���<<�<pP�<���<!��<r��<Q�<�7�<Wa�<b��<ǯ�<Q��<��<��<�6�<OS�<�m�<���<ޛ�<L��<=��<���<!��<���<���<���<`��<���<0��<!��<q��<W��<r��<Ҋ�<[n�<�M�<~)�<� �<;��<'��<�m�<$4�<���<U��<l�<S �<���<�z�<8!�<���<�_�<o��<N��<��<e��<�,�<���<,�<3��<7�<��<���<�`�<�ů<�&�<C��<Hު<�4�<���<�ץ<�$�<�n�<���<���<�;�<�z�<z��<�<p*�<�`�<h��<Ȑ<E��<�(�<�V�<���<M��<�م<T�<,�<�S�<��|<�Cy<��u<��q<5(n<�sj<$�f<c<W_<�[<��W<w@T<��P<]�L<�5I<C�E<��A<=><��:<S�6<�[3<��/<b+,<ɘ(<3
%<�!<��<�x<��<�<�<��<C	<s�<%�<ao�;���;xN�;p��;�g�;��;��;���;�V�;�;�;22�;*:�;�S�;~�;���;��;�p�;��;o�;r
�;���;�y�;Śx;1hn;sZd;rZ;�P;G;��=;"94;�+;��!;��;U,;"{;���:���:OC�:��:Û�:~��:Mϛ:�7�:X�y:�6[:�%=:�r:�:��90��9Rt/9��{8nSB�n��q*��[�������h.�VH�]b�.6|����ɰ��s]������|����ɺHVֺK�����+��y����	�������%��t�!���'���-�X�3���9��r?��XE��<K�\Q�r�V���\�_�b���h��pn��Kt��%z� ��v킻�څ��Ȉ�����¥��7��������v��i���  �  Hu=�=�=�X=��=B�=�:=�� =jz =� =r�<¯�<���<�(�<bd�<���<���<��<[I�<7��<���<���<*�<yP�<���<+��<v��<B�<�7�<Sa�<m��<���<W��<��<��<�6�<AS�<�m�<���<���<Q��<9��<���<��<���<���<���<[��<���<3��<��<y��<T��<q��<֊�<bn�<�M�<�)�<� �<;��<2��<�m�<(4�<���<L��<l�<R �<���<�z�<4!�<���<�_�<u��<H��<��<[��<�,�<|��<,�<9��<0�<��<���<�`�<�ů<�&�<M��<Iު<�4�<燧<�ץ<�$�<�n�<���<���<�;�<�z�<���<�<v*�<�`�<f��<Ȑ<<��<�(�<�V�<���<Q��<�م<b�< ,�<�S�<t�|<�Cy<��u<��q<N(n<�sj<�f<�
c<W_<�[<��W<�@T<��P<e�L<�5I<Y�E<��A<=><��:<5�6<�[3<��/<l+,<̘(<)
%<�!<�<�x<��<�<�<ɨ<C	<b�<%�<o�;���;|N�;���;�g�;a�;��;���;�V�;�;�;J2�;9:�;�S�;\�;v��;��;�p�;��;o�;a
�;���;�y�;,�x;Ahn;�Zd;�qZ;�P; G;X�=;b94;�+;��!;��;�,;|{;,��:���:AC�:���:���:���:ϛ:�6�:<�y:�6[:_'=:�q:F: �9|��9w/9x�{8�?B�x��W,��^�� �9��4.�QUH��]b��5|�����Ű���\�����D|����ɺoVֺ�����K+����z�	�z�������D�!��'�̮-�*�3�։9��r?�YE��<K�<Q�B�V�Q�\�͹b���h��pn�NKt��%z� ��E킻�څ��Ȉ�䶋�����&��������v��&i���  �  �v=�=(�=u[=��=z�=!>=�� =�~ ={ =�{�<j��<��<5�<Bq�<���<I��<� �<�Y�<f��<��<���<*2�<ye�<j��<4��<���<e%�<�Q�<�|�<��<f��<'��<�<9�<)Y�<�v�<˒�<H��<���<I��<���<;��<�<B�<Y�<��<��<��<�<8�<� �<���<G��<���<T��<���<�g�<�?�<��<���<(��<
v�<z8�<E��<q��<�c�<��<���<e�<��<t��<�;�<���<�]�<��<�m�<��<k�<U�<;W�<Ǵ<w2�<��<���<f]�<p��<��<�f�<A��<��<�Q�<͙�<ߠ<�!�<ma�<���<�ٙ<V�<�H�<�}�<!��<�<.�<�=�<&j�<��<ξ�<p�<2�<�5�<\�<�}<�Ly<��u<��q<�%n<_mj<N�f<'�b<�E_<��[<��W<�#T<FpP<��L<
I<�_E<��A<�	><�b:<;6<�3<�/<��+<mO(<0�$< /!<��<� <#�<�&<ݱ<�B<��<iv<<���;���;J[�;��;�i�;��;���;�t�; E�;�%�;�;K�;�2�;\�;!��;��;�F�;���;C�;�݊;W��;jM�;�Dv;Pl;J	b;_$X;�dN;��D;T;;E2;.�(;��;��;�;�l;���:���:�a�:��:"�:1��:F�:�Ĉ:��r:��T:k�6:�D:a+�9�n�9wO�9��9��&8����2�쳏�M�Ź�������)?2��ML�[2f�(������b������/��������_˺δ׺���;2�\���<�lE
�!I�5G��@��4"��$(�.��3�u�9�V�?���E�łK��^Q��9W��]�Z�b��h�]�n��lt��Az���������ᅻ�̈�ʸ��6���[�������n���^���  �  �v=�="�=t[=��=x�=#>=�� =�~ =y =�{�<_��<��<5�<Mq�<���<;��<� �<�Y�<f��<#��<���<-2�<re�<~��<+��<���<]%�<�Q�<�|�<��<d��<3��<�<9�<Y�<w�<Ԓ�<W��<���<D��<���<#��<�<5�<f�<��<��<��<$�<K�<� �<���<5��<���<_��< ��<�g�<�?�<�<���<8��<"v�<~8�<D��<r��<�c�<��<���<e�<��<s��<�;�<��<�]�<��<wm�<��<#k�<a�<?W�<�ƴ<~2�<��<���<Z]�<b��<��<�f�<C��<��<�Q�<ә�<	ߠ<�!�<^a�<���<�ٙ<g�<�H�<y}�<!��< �<E�<�=�<+j�<��<ھ�<s�<%�<�5�<�[�<�}<�Ly<}�u<��q<�%n<hmj<�f<$�b<�E_<Ԏ[<��W<�#T<XpP<X�L<I<�_E<��A<
><�b:<־6<�3<�/<��+<fO(<�$</!<��<� <?�<�&<ұ<�B<��<�v<<���;���;�[�;���;�i�;��;4��;u�;�D�;�%�;A�;y�;�2�;�[�;>��;��;G�;S��;�B�;�݊;���;mM�;MDv;�l;p	b;J$X;�dN;��D;�T;;�2;T�(;*�;s�;�;m;���:v��:b�:!�:*�:���:ZF�:�Ĉ:��r:q�T:��6:�D:&�9�k�9O�9 �9G�&8s����2������Ź�������>2�[PL�l1f���ŵ��nc������ꄲ������_˺W�׺����1�\��=��E
��H��F�@��4"�%(�.�>�3���9���?�g�E�݂K��^Q�p9W�;]�^�b��h�*�n��lt�.Bz����q����ᅻ͈�и������������n���^���  �  �v=�= �=u[=��=u�=%>=� =�~ =w =|�<j��<��<5�<:q�<���<?��<� �<�Y�<a��<��<���<82�<he�<���<&��<���<r%�<�Q�<�|�<ץ�<g��<#��<�<9�<Y�<w�<���<\��<z��<O��<���<&��<%�<*�<l�<��<��<��<�<B�<� �< ��<9��<���<[��<���<�g�<�?�<�<���<1��<v�<r8�<H��<h��<�c�<��<˾�<e�<��<���<�;�<��<�]�<��<{m�<��<k�<N�<DW�<�ƴ<�2�<��<���<e]�<Z��<��<�f�<K��<{�<�Q�<Ι�<ߠ<�!�<aa�<Ş�<�ٙ<h�<�H�<�}�<6��<���<?�<�=�<+j�<��<ؾ�<v�<�<�5�<�[�<�}<�Ly<v�u<��q<�%n<{mj<)�f<7�b<�E_<Ŏ[<��W<�#T<|pP<L�L<4I<�_E<��A<
><�b:<޾6<�3<�/<��+<�O(<0�$</!<��<� <G�<�&<��<�B<y�<�v<�<���;���;�[�;���;�i�;�;%��;Vu�;�D�;�%�;�;\�;�2�;�[�;\��;g�;G�;8��;C�;ފ;��;�M�;�Cv;�l;*	b;]$X;�dN;��D;^T;;2;�(;Q�;��;�;�l;g��:���:�c�:Q�:��:���:�E�:ň:��r:8�T:!�6:�F:>(�9�n�9.S�9��9�'8<���2�����ՔŹ���Y���=2��QL�/f���������b��8���h���v���6_˺��׺���*2��[��x<��E
��H�WG�@��4"�3%(�l.�J�3���9���?�g�E��K��^Q�U9W��]���b�?�h���n��lt�KBz��������xᅻ�̈�����V���0���%����n���^���  �  �v=�=�=z[=��=y�=(>=�� =�~ =} = |�<c��<��<5�<Sq�<���<H��<� �<�Y�<m��<#��<���<=2�<ne�<z��<0��<���<b%�<�Q�<�|�<٥�<m��<��<�<9�<
Y�<w�<���<Q��<���<@��<���<"��<�<0�<n�<��<��<��<�<N�<� �<���<>��<���<c��<��<�g�<�?�<�<���<<��<!v�<�8�<M��<g��<�c�<��<���<e�<��<o��<�;�<��<�]�<��<nm�<�<k�<L�<EW�<�ƴ<z2�<���<���<[]�<e��<��<�f�<N��<��<�Q�<ٙ�<ߠ<�!�<ja�<Ş�<�ٙ<j�<�H�<}�<%��<�<J�<�=�<4j�<��<ξ�<�<�<�5�<�[�<�}<�Ly<��u<��q<�%n<fmj<�f<$�b<�E_<��[<��W<�#T<KpP<V�L<I<�_E<ǳA<
><�b:<�6<�3<�/<��+<uO(<!�$<(/!<��<� <H�<�&<۱<�B<��<�v<<Ј�;���;�[�;��;�i�;��;)��;�t�;�D�;�%�;��;\�;�2�;�[�;9��;o�;�F�;R��;�B�;�݊;���;}M�;/Dv;�l;	b;�$X;DeN;��D;�T;;z2;c�(;x�;��; ;:m;|��:��:Mb�:�:n�:���:�F�:pň:��r:"�T:Y�6:�D:&�9�j�9UN�9��9�&8���ٽ2����s�Ź�������=2�/QL��1f��������Wc��}������A����^˺��׺���1�[���<�E
��H��F��?��4"�Q%(��.���3���9�	�?�!�E���K��^Q�9W�u]�'�b��h�_�n��lt�Bz���������ᅻ&͈�и��D���L������	o���^���  �  �v=�= �=u[=��=�= >=�� =�~ =} =|�<n��<"��<5�<dq�<���<P��<� �<�Y�<e��<��<���<,2�<|e�<w��<,��<~��<a%�<�Q�<�|�<٥�<S��<��<�<9�<Y�<�v�<ɒ�<>��<{��<B��<���<.��<�<2�<`�<��<��<��<$�<<�<� �<���<P��<���<i��<��<�g�<�?�<�<���<+��<!v�<y8�<G��<q��<�c�<��<���<e�<��<p��<�;�<���<�]�<��<nm�<y�<k�<I�<+W�<�ƴ<x2�<��<���<W]�<c��<��<�f�<@��<��<�Q�<͙�<ߠ<�!�<ta�<���<�ٙ<g�<�H�<�}�<.��<�<;�<�=�<'j�<��<о�<s�<!�<�5�<\�<�}<�Ly<g�u<��q<�%n<Qmj<�f<�b<�E_<��[<��W<�#T<NpP<m�L<
I<�_E<��A<
><c:<ʾ6<�3<�/<��+<�O(<9�$<2/!<��<!<.�<�&<�<�B<��<�v<<���;��;�[�;���;�i�;��;^��;�t�;�D�;Y%�;��;N�;�2�;�[�;��;��;�F�;?��;�B�;�݊;'��;\M�;BDv;�l;M	b;�$X;�dN;��D;1T;;�2;��(;�;��;S;�m;���:��:�b�:x�:k�:���:F�:ň:��r:��T:`�6:D:�(�9Qm�9�N�9�9.�&8m����2�ͺ��Ź��������@2�@QL�2f����S����c������M���j����_˺��׺��32�G[���<�4E
�I�:F�@��4"��$(��.���3��9���?���E�t�K��^Q�r9W�Z]�\�b���h�P�n��lt��Bz��������ᅻ͈�����*�������Q����n���^���  �  �v=�=�=s[=��=|�='>=�� =�~ = =|�<n��</��<!5�<]q�<���<Z��<� �<�Y�<k��<$��<���<82�<se�<z��<&��<���<g%�<�Q�<�|�<ӥ�<\��<��<��<�8�<Y�<�v�<���<G��<y��<;��<{��<��<�<.�<c�<��<��<��<0�<E�<� �<���<J��<���<q��<��<�g�<�?�<�<���<5��<+v�<�8�<O��<l��<�c�<��<���<e�<��<g��<�;�<���<�]�<��<om�<s�<k�<K�<4W�<�ƴ<o2�<���<���<\]�<Z��<��<�f�<K��<��<�Q�<ՙ�<%ߠ<�!�<{a�<ʞ�<�ٙ<v�<
I�<�}�<9��<�<C�<�=�</j�<��<Ӿ�<r�<�<�5�<�[�<�}<vLy<k�u<��q<�%n<1mj<�f<��b<pE_<��[<��W<�#T<HpP<7�L<I<�_E<��A<
><c:<�6<�3<�/<��+<�O(<9�$<M/!<��<!<Q�<�&<�<�B<��<�v<-<���;���;�[�;���;�i�;��;���;�t�;�D�;�%�;��;�;�2�;�[�;Ж�;U�;�F�;7��;�B�;�݊;鋅;M�;!Dv;�l;F	b;�$X;0eN;�D;{T;;�2;��(;��;	�;�;�m;���:���:�b�:��:�:S��:�F�:�ň:F�r:
�T:��6:E: &�9Ei�9�L�9��9��&8r����2�q����Ź�������?2�RL�*3f����7���*c��)�����������)_˺ܳ׺��㺳1��Z���<��D
�zH�aF��?�4"��$(�X.���3���9���?�H�E���K��^Q�y9W�k]��b��h���n�/mt�vBz��������ⅻ͈�0�������k���?���o���^���  �  �v=�=�=y[=��=w�=)>=�� =�~ =� =|�<v��<3��<-5�<aq�<ͬ�<[��< !�<�Y�<t��</��<���<=2�<le�<���<+��<u��<c%�<�Q�<�|�<ʥ�<S��<��<��<�8�<�X�<�v�<���<;��<m��<6��<}��<��<�<$�<w�<��<��<��<)�<U�<� �<���<O��<���<t��<��<�g�<�?�<�<���<A��<(v�<�8�<M��<i��<�c�<��<���<�d�<��<e��<~;�<���<�]�<��<_m�<k�<	k�<9�<)W�<�ƴ<t2�<���<���<Q]�<[��<��<�f�<O��<��<�Q�<ߙ�<ߠ<�!�<{a�<מ�<�ٙ<~�<I�<�}�<<��<�<V�<�=�<6j�<��<׾�<��<�<�5�<�[�<�}<jLy<[�u<��q<�%n<>mj<��f<��b<vE_<��[<��W<�#T<TpP<3�L<I<�_E<ƳA<
><�b:<�6<�3<1�/<��+<�O(<I�$<T/!<ե<!<n�<�&<�<�B<��<�v<<؈�;���;�[�;���;ji�;��;��;�t�;lD�;^%�;��;�;�2�;`[�;���;>�;�F�;��;�B�;�݊;ދ�;M�;�Cv;Ml;1	b;�$X;6eN;��D;�T;;�2;�(;�;e�;�;�m;���:9��:�c�:��:��:#��:�F�:�ň:��r:��T:��6:�D:�$�9�i�9`L�9r�9�&8.(����2�[���ޛŹ������A2��RL�j2f�A�������c��������_����^˺7�׺9��1�[��=<��D
�H�;F�Q?��3"��$(�=.���3�7�9���?��E�˂K��^Q� 9W��]�+�b���h�G�n�]mt��Bz�#�������ᅻY͈����w�������\���Bo���^���  �  �v=�=�=t[=��=�=*>=�� =�~ =� =|�<���</��<)5�<sq�<Ŭ�<\��<!�<�Y�<z��<)��<���<?2�<{e�<w��<*��<|��<]%�<�Q�<�|�<ɥ�<O��<��<��<�8�<�X�<�v�<���<2��<s��<,��<y��< ��<�<)�<h�<��<��<��<%�<Q�<� �<
��<^��<���<~��<"��<�g�<@�<"�<���<A��<%v�<�8�<Q��<k��<�c�<��<���<e�<��<Z��<�;�<���<�]�<��<Ym�<f�<�j�<3�<"W�<�ƴ<b2�<���<���<V]�<]��<��<�f�<O��<��<�Q�<㙢<*ߠ<�!�<a�<Ξ�<�ٙ<~�<
I�<�}�<D��<�<P�<�=�<9j�<#��<о�<u�<�<�5�<�[�<�}<XLy<Y�u<��q<�%n<#mj<�f<��b<qE_<|�[<��W<�#T<3pP<D�L<
I<�_E<��A<
><c:<�6<�3<'�/< �+<�O(<e�$<M/!<Υ<?!<`�< '< �<�B<��<�v<$<���;
��;�[�;���;�i�;��;#��;�t�;lD�;P%�;��;�;q2�;O[�;ɖ�;A�;uF�;$��;�B�;�݊;�;oM�;�Cv;�l;,	b;�$X;seN;��D;�T;;�2;o�(;��;8�;�;;n;>��:���:Od�:,	�:��:��:G�:�ň:C�r:9�T:N�6:�D:�%�9�i�9�I�9�9�&8�*���2�����ٜŹ���j���A2��RL��4f�s��˵��c������J��������^˺�׺w���0�rZ���;��D
�WH��E�N?�4"�5$(��.�O�3�f�9���?���E�N�K��^Q�b9W��]�Z�b�O�h���n��mt��Bz�K������(ⅻg͈�R�����������j���Yo��_���  �  �v=�= �=s[=��=�='>=�� =�~ =� =|�<��<E��<65�<sq�<լ�<p��<!�<�Y�<���<0��<���<62�<}e�<v��<'��<}��<U%�<�Q�<�|�<ǥ�<E��<	��<��<�8�<�X�<�v�<���<*��<l��<#��<r��<��<�<1�<b�<��<��<��<<�<Z�<�<��<_��<���<���<"��<�g�<
@�<�<���<H��<8v�<�8�<I��<r��<�c�<��<���<�d�<��<N��<|;�<���<�]�<��<Wm�<\�<�j�<8�<W�<�ƴ<X2�<�<���<Q]�<]��<��<�f�<F��<��<�Q�<Ꙣ<*ߠ<�!�<�a�<ݞ�<�ٙ<��<I�<�}�<=��<#�<U�<>�<1j�<��<վ�<s�< �<�5�<�[�<�}<QLy<G�u<��q<r%n<mj<��f<��b<XE_<{�[<��W<�#T<'pP<:�L<�I<�_E<��A<
><c:<�6<�3<,�/<�+<�O(<\�$<y/!<�<?!<��<*'<�<�B<��<�v<V<�;��;�[�;���;�i�;��;��;�t�;eD�;+%�;��;��;;2�;\[�;{��;-�;XF�;��;xB�;�݊;ʋ�;FM�;EDv;�l;y	b;�$X;�eN;}�D;*U;;(2;)�(;��;��;;:n;0��:C��:�c�:o	�:Q�::��:�G�:Xň:2�r:��T:&�6:_C:#�9gg�9�F�9;�9��&8J+��@�2�տ��W�Ź�������B2�?SL��5f����Z����c������t���U���R_˺�׺���R0�`Z�� <�DD
��G��E�?�}3"�Z$(�8.�(�3�@�9���?�9�E�r�K��^Q�u9W�`]���b���h�ؗn��mt�Cz�Y�����hⅻL͈���������������do��1_���  �  �v=�=�=t[=��=~�=)>=�� =�~ =� =-|�<���<A��<@5�<mq�<��<f��<!�<�Y�<���<-��<���<>2�<ze�<���<$��<w��<b%�<�Q�<�|�<¥�<;��<���<��<�8�<�X�<�v�<���<&��<e��<0��<v��<��<�<$�<f�<��<��<��<-�<[�<�<��<_��<���<���<"��<�g�<@�<1�<���<G��<+v�<�8�<O��<r��<�c�<��<���<�d�<��<]��<t;�<���<�]�<��<Lm�<W�<�j�<%�<W�<�ƴ<i2�<꙱<���<Q]�<V��<��<�f�<N��<��<�Q�<虢<2ߠ<�!�<�a�<螛<�ٙ<��<I�<�}�<U��<#�<U�<�=�<4j�<��<۾�<u�<�<�5�<�[�<�}<\Ly<:�u<t�q<b%n<mj<ٴf<��b<KE_<g�[<z�W<�#T<6pP<)�L<I<�_E<��A<
><c:<�6<�3<+�/<�+<�O(<u�$<r/!<��<4!<��<'<1�<C<��<�v<?<߈�;	��;�[�;���;xi�;��;��;�t�;TD�;%�;n�;��;=2�;0[�;���;�;IF�;�;�B�;�݊;ʋ�;{M�;�Cv;�l;�	b;�$X;SeN;�D;2U;;62;��(;��;��;6;;n;���:+��:=e�:�	�:F�:f��:�F�:�ň:Y�r:�T:��6:oD:L$�9�g�9�J�9e�9��&899����2���e�Źt�����D2��SL��3f���������c��H������������^˺��׺5��g0��Y���;��D
��G��E��>�p3"�!$(�v.�&�3�:�9�j�?��E�i�K��^Q�^9W��]�1�b���h���n��mt�7Cz�u��3���9ⅻ�͈�h���ʥ��꒑�����]o��_���  �  �v=�=�=y[=��=��=1>=�� =�~ =� =&|�<���<<��<I5�<yq�<��<a��<!�<�Y�<���<D��<���<M2�<we�<|��<-��<p��<X%�<�Q�<�|�<���<O��<���<��<�8�<�X�<�v�<���<5��<`��<%��<g��<��<�<"�<p�<��<��<��<5�<q�<� �<��<`��<���<���<-��<�g�<@�<5�<���<\��<:v�<�8�<]��<g��<�c�<��<���<�d�<y�<S��<k;�<���<�]�<��<=m�<P�<�j�<"�<%W�<�ƴ<]2�<ؙ�<���<I]�<[��<��<�f�<^��<��<�Q�<���<+ߠ<�!�<�a�<�<�ٙ<��<I�<�}�<N��<$�<m�<�=�<Ej�<&��<Ѿ�<��<�<�5�<�[�<�}<BLy<@�u<��q<Q%n<mj<��f<��b<=E_<x�[<��W<�#T<"pP<�L<I<�_E<ĳA<	
><c:<�6<�3<\�/<�+<�O(<��$<j/!<�<M!<��<'<E�<�B<��<�v<6<��;���;�[�;��;]i�;��;���;�t�;D�;V%�;u�;��;02�;�Z�;���;��;�F�;ܺ�;�B�;p݊;���;hM�;�Cv; l;%	b;&%X;�eN;J�D;�U;;2;��(;��;��;�;�n;��:��:�e�:Q	�:��:Z��:�G�:�ƈ:��r:_�T:��6:�C:f �9�c�9UH�9�9(�&8�A��R�2�Ə��Ź5��T��.A2��UL��4f����Y���4d������Ą�������]˺��׺��㺓/�TZ��?;��D
�3G�rE�w>�s3"��#(��.��3�z�9�z�?���E�6�K��^Q�9W�]�R�b�1�h��n��mt�"Cz�E��T���9ⅻ�͈�i���祎�Ȓ�������o��;_���  �  �v=�=�=x[=��=��=&>=�� =�~ =� ='|�<���<L��<?5�<uq�<��<y��<!!�<�Y�<���<4��<���<72�<e�<w��<0��<p��<Y%�<�Q�<�|�<���<9��<���<��<�8�<�X�<�v�<���<"��<W��<*��<t��<��<�<+�<h�<��<��<��<2�<]�<�<��<s��<���<���<)��<�g�<@�</�<���<J��<0v�<�8�<L��<q��<�c�<��<���<�d�<��<X��<f;�<���<�]�<��<Gm�<R�<�j�<�<W�<�ƴ<d2�<�<���<G]�<b��<��<�f�<I��<��<�Q�<왢<1ߠ<�!�<�a�<ꞛ<�ٙ<��<'I�<�}�<M��<+�<Z�<>�</j�<"��<վ�<{�<�<�5�<�[�<�}<LLy<�u<l�q<J%n<mj<дf<��b<5E_<_�[<g�W<�#T<6pP<6�L<�I<�_E<��A<
><c:<�6<�3<7�/<"�+<�O(<��$<�/!<��<C!<��<<'<J�<C<��<�v<A<Ɉ�;"��;�[�;��;_i�;��;��;�t�;D�;�$�;U�;��;02�;[�;���;��;<F�;���;�B�;�݊;ڋ�;NM�;Dv;�l;h	b;�$X;GeN;2�D;JU;;`2;��(;1�;�;Y;yn;���:_��:'e�:�	�:x�:���:�F�:�ň:J�r:��T:��6:-C:�#�9�g�9�I�9��9D�&8>D����2��Ï�y�Ź'	�� �D2��UL�4f�������Vd��v���.���?���_˺��׺���0��Y��R;��C
�wG��E��>�*3"��#(��.���3��9�L�?�F�E�T�K��^Q�49W��]���b�}�h���n��mt��Cz����d���Hⅻ�͈�r�����������ـ��|o��_���  �  �v=�=�=o[=��=��='>=�� =�~ =� =-|�<���<B��<C5�<�q�<۬�<o��<!�<�Y�<���<0��<���<72�<�e�<r��<'��<s��<S%�<�Q�<||�<���<7��<��<��<�8�<�X�<�v�<���<$��<`��<"��<Y��<��<�<.�<U�<��<��<��<F�<X�<�<��<g��<���<���<;��<�g�<@�<$�<��<I��<?v�<�8�<Q��<���<�c�<��<���<�d�<p�<I��<m;�<���<�]�<��<<m�<E�<�j�<.�<
W�<�ƴ<Q2�<ܙ�<���<J]�<\��<��<�f�<I��<��<�Q�<�<Cߠ<�!�<�a�<㞛<�ٙ<��<I�<�}�<Q��<9�<Q�<>�<5j�</��<۾�<g�<�<�5�<�[�<o}<NLy</�u<y�q<`%n<�lj<��f<��b<EE_<r�[<q�W<�#T<�oP<�L<�I<�_E<��A<
><1c:<�6<+3<#�/<4�+<�O(<q�$<u/!<�<s!<��<)'<&�<C<��<�v<|<ʈ�;Z��;[�;���;ki�;��;���;qt�;ED�;�$�;��;��;�1�;�Z�;{��;�;CF�;޺�;wB�;:݊;���;KM�;0Dv;Jl;�	b;%X;�eN;��D;"U;;2;��(;��;��;�;o;���:���:vd�:&�:l�:���:H�:�ň:Q�r:��T:��6:'C:�"�9da�9�E�9N�9Z�&8�2����2�8Ə���Źl������D2��TL�l6f�b��X���$d������Ӆ��]���'_˺��׺����/��X���;�AD
��G��D��>��3"��#(��.�p�3�]�9�i�?��E��K��^Q��9W�~]���b���h���n��mt�dCz�j��8����ⅻ�͈�����֥��Ւ��Ā��no���_���  �  �v=�=�=x[=��=��=&>=�� =�~ =� ='|�<���<L��<?5�<uq�<��<y��<!!�<�Y�<���<4��<���<72�<e�<w��<0��<p��<Y%�<�Q�<�|�<���<9��<���<��<�8�<�X�<�v�<���<"��<W��<*��<t��<��<�<+�<h�<��<��<��<2�<]�<�<��<s��<���<���<)��<�g�<@�</�<���<J��<0v�<�8�<L��<q��<�c�<��<���<�d�<��<X��<f;�<���<�]�<��<Gm�<R�<�j�<�<W�<�ƴ<d2�<�<���<G]�<b��<��<�f�<I��<��<�Q�<왢<1ߠ<�!�<�a�<ꞛ<�ٙ<��<'I�<�}�<M��<+�<Z�<>�</j�<"��<վ�<{�<�<�5�<�[�<�}<LLy<�u<l�q<J%n<mj<дf<��b<5E_<_�[<g�W<�#T<6pP<6�L<�I<�_E<��A<
><c:<�6<�3<7�/<"�+<�O(<��$<�/!<��<C!<��<<'<J�<C<��<�v<A<Ɉ�;"��;�[�;��;_i�;��;��;�t�;D�;�$�;U�;��;02�;[�;���;��;<F�;���;�B�;�݊;ڋ�;NM�;Dv;�l;h	b;�$X;GeN;2�D;JU;;`2;��(;1�;�;Y;yn;���:_��:'e�:�	�:x�:���:�F�:�ň:J�r:��T:��6:-C:�#�9�g�9�I�9��9D�&8>D����2��Ï�y�Ź'	�� �D2��UL�4f�������Vd��v���.���?���_˺��׺���0��Y��R;��C
�wG��E��>�*3"��#(��.���3��9�L�?�F�E�T�K��^Q�49W��]���b�}�h���n��mt��Cz����d���Hⅻ�͈�r�����������ـ��|o��_���  �  �v=�=�=y[=��=��=1>=�� =�~ =� =&|�<���<<��<I5�<yq�<��<a��<!�<�Y�<���<D��<���<M2�<we�<|��<-��<p��<X%�<�Q�<�|�<���<O��<���<��<�8�<�X�<�v�<���<5��<`��<%��<g��<��<�<"�<p�<��<��<��<5�<q�<� �<��<`��<���<���<-��<�g�<@�<5�<���<\��<:v�<�8�<]��<g��<�c�<��<���<�d�<y�<S��<k;�<���<�]�<��<=m�<P�<�j�<"�<%W�<�ƴ<]2�<ؙ�<���<I]�<[��<��<�f�<^��<��<�Q�<���<+ߠ<�!�<�a�<�<�ٙ<��<I�<�}�<N��<$�<m�<�=�<Ej�<&��<Ѿ�<��<�<�5�<�[�<�}<BLy<@�u<��q<Q%n<mj<��f<��b<=E_<x�[<��W<�#T<"pP<�L<I<�_E<ĳA<	
><c:<�6<�3<\�/<�+<�O(<��$<j/!<�<M!<��<'<E�<�B<��<�v<6<��;���;�[�;��;]i�;��;���;�t�;D�;V%�;u�;��;02�;�Z�;���;��;�F�;ܺ�;�B�;p݊;���;hM�;�Cv; l;%	b;&%X;�eN;J�D;�U;;2;��(;��;��;�;�n;��:��:�e�:Q	�:��:Z��:�G�:�ƈ:��r:_�T:��6:�C:f �9�c�9UH�9�9(�&8�A��R�2�Ə��Ź5��T��.A2��UL��4f����Y���4d������Ą�������]˺��׺��㺓/�TZ��?;��D
�3G�rE�w>�s3"��#(��.��3�z�9�z�?���E�6�K��^Q�9W�]�R�b�1�h��n��mt�"Cz�E��T���9ⅻ�͈�i���祎�Ȓ�������o��;_���  �  �v=�=�=t[=��=~�=)>=�� =�~ =� =-|�<���<A��<@5�<mq�<��<f��<!�<�Y�<���<-��<���<>2�<ze�<���<$��<w��<b%�<�Q�<�|�<¥�<;��<���<��<�8�<�X�<�v�<���<&��<e��<0��<v��<��<�<$�<f�<��<��<��<-�<[�<�<��<_��<���<���<"��<�g�<@�<1�<���<G��<+v�<�8�<O��<r��<�c�<��<���<�d�<��<]��<t;�<���<�]�<��<Lm�<W�<�j�<%�<W�<�ƴ<i2�<꙱<���<Q]�<V��<��<�f�<N��<��<�Q�<虢<2ߠ<�!�<�a�<螛<�ٙ<��<I�<�}�<U��<#�<U�<�=�<4j�<��<۾�<u�<�<�5�<�[�<�}<\Ly<:�u<t�q<b%n<mj<ٴf<��b<KE_<g�[<z�W<�#T<6pP<)�L<I<�_E<��A<
><c:<�6<�3<+�/<�+<�O(<u�$<r/!<��<4!<��<'<1�<C<��<�v<?<߈�;	��;�[�;���;xi�;��;��;�t�;TD�;%�;n�;��;=2�;0[�;���;�;IF�;�;�B�;�݊;ʋ�;{M�;�Cv;�l;�	b;�$X;SeN;�D;2U;;62;��(;��;��;6;;n;���:+��:=e�:�	�:F�:f��:�F�:�ň:Y�r:�T:��6:oD:L$�9�g�9�J�9e�9��&899����2���e�Źt�����D2��SL��3f���������c��H������������^˺��׺5��g0��Y���;��D
��G��E��>�p3"�!$(�v.�&�3�:�9�j�?��E�i�K��^Q�^9W��]�1�b���h���n��mt�7Cz�u��3���9ⅻ�͈�h���ʥ��꒑�����]o��_���  �  �v=�= �=s[=��=�='>=�� =�~ =� =|�<��<E��<65�<sq�<լ�<p��<!�<�Y�<���<0��<���<62�<}e�<v��<'��<}��<U%�<�Q�<�|�<ǥ�<E��<	��<��<�8�<�X�<�v�<���<*��<l��<#��<r��<��<�<1�<b�<��<��<��<<�<Z�<�<��<_��<���<���<"��<�g�<
@�<�<���<H��<8v�<�8�<I��<r��<�c�<��<���<�d�<��<N��<|;�<���<�]�<��<Wm�<\�<�j�<8�<W�<�ƴ<X2�<�<���<Q]�<]��<��<�f�<F��<��<�Q�<Ꙣ<*ߠ<�!�<�a�<ݞ�<�ٙ<��<I�<�}�<=��<#�<U�<>�<1j�<��<վ�<s�< �<�5�<�[�<�}<QLy<G�u<��q<r%n<mj<��f<��b<XE_<{�[<��W<�#T<'pP<:�L<�I<�_E<��A<
><c:<�6<�3<,�/<�+<�O(<\�$<y/!<�<?!<��<*'<�<�B<��<�v<V<�;��;�[�;���;�i�;��;��;�t�;eD�;+%�;��;��;;2�;\[�;{��;-�;XF�;��;xB�;�݊;ʋ�;FM�;EDv;�l;y	b;�$X;�eN;}�D;*U;;(2;)�(;��;��;;:n;0��:C��:�c�:o	�:Q�::��:�G�:Xň:2�r:��T:&�6:_C:#�9gg�9�F�9;�9��&8J+��@�2�տ��W�Ź�������B2�?SL��5f����Z����c������t���U���R_˺�׺���R0�`Z�� <�DD
��G��E�?�}3"�Z$(�8.�(�3�@�9���?�9�E�r�K��^Q�u9W�`]���b���h�ؗn��mt�Cz�Y�����hⅻL͈���������������do��1_���  �  �v=�=�=t[=��=�=*>=�� =�~ =� =|�<���</��<)5�<sq�<Ŭ�<\��<!�<�Y�<z��<)��<���<?2�<{e�<w��<*��<|��<]%�<�Q�<�|�<ɥ�<O��<��<��<�8�<�X�<�v�<���<2��<s��<,��<y��< ��<�<)�<h�<��<��<��<%�<Q�<� �<
��<^��<���<~��<"��<�g�<@�<"�<���<A��<%v�<�8�<Q��<k��<�c�<��<���<e�<��<Z��<�;�<���<�]�<��<Ym�<f�<�j�<3�<"W�<�ƴ<b2�<���<���<V]�<]��<��<�f�<O��<��<�Q�<㙢<*ߠ<�!�<a�<Ξ�<�ٙ<~�<
I�<�}�<D��<�<P�<�=�<9j�<#��<о�<u�<�<�5�<�[�<�}<XLy<Y�u<��q<�%n<#mj<�f<��b<qE_<|�[<��W<�#T<3pP<D�L<
I<�_E<��A<
><c:<�6<�3<'�/< �+<�O(<e�$<M/!<Υ<?!<`�< '< �<�B<��<�v<$<���;
��;�[�;���;�i�;��;#��;�t�;lD�;P%�;��;�;q2�;O[�;ɖ�;A�;uF�;$��;�B�;�݊;�;oM�;�Cv;�l;,	b;�$X;seN;��D;�T;;�2;o�(;��;8�;�;;n;>��:���:Od�:,	�:��:��:G�:�ň:C�r:9�T:N�6:�D:�%�9�i�9�I�9�9�&8�*���2�����ٜŹ���j���A2��RL��4f�s��˵��c������J��������^˺�׺w���0�rZ���;��D
�WH��E�N?�4"�5$(��.�O�3�f�9���?���E�N�K��^Q�b9W��]�Z�b�O�h���n��mt��Bz�K������(ⅻg͈�R�����������j���Yo��_���  �  �v=�=�=y[=��=w�=)>=�� =�~ =� =|�<v��<3��<-5�<aq�<ͬ�<[��< !�<�Y�<t��</��<���<=2�<le�<���<+��<u��<c%�<�Q�<�|�<ʥ�<S��<��<��<�8�<�X�<�v�<���<;��<m��<6��<}��<��<�<$�<w�<��<��<��<)�<U�<� �<���<O��<���<t��<��<�g�<�?�<�<���<A��<(v�<�8�<M��<i��<�c�<��<���<�d�<��<e��<~;�<���<�]�<��<_m�<k�<	k�<9�<)W�<�ƴ<t2�<���<���<Q]�<[��<��<�f�<O��<��<�Q�<ߙ�<ߠ<�!�<{a�<מ�<�ٙ<~�<I�<�}�<<��<�<V�<�=�<6j�<��<׾�<��<�<�5�<�[�<�}<jLy<[�u<��q<�%n<>mj<��f<��b<vE_<��[<��W<�#T<TpP<3�L<I<�_E<ƳA<
><�b:<�6<�3<1�/<��+<�O(<I�$<T/!<ե<!<n�<�&<�<�B<��<�v<<؈�;���;�[�;���;ji�;��;��;�t�;lD�;^%�;��;�;�2�;`[�;���;>�;�F�;��;�B�;�݊;ދ�;M�;�Cv;Ml;1	b;�$X;6eN;��D;�T;;�2;�(;�;e�;�;�m;���:9��:�c�:��:��:#��:�F�:�ň:��r:��T:��6:�D:�$�9�i�9`L�9r�9�&8.(����2�[���ޛŹ������A2��RL�j2f�A�������c��������_����^˺7�׺9��1�[��=<��D
�H�;F�Q?��3"��$(�=.���3�7�9���?��E�˂K��^Q� 9W��]�+�b���h�G�n�]mt��Bz�#�������ᅻY͈����w�������\���Bo���^���  �  �v=�=�=s[=��=|�='>=�� =�~ = =|�<n��</��<!5�<]q�<���<Z��<� �<�Y�<k��<$��<���<82�<se�<z��<&��<���<g%�<�Q�<�|�<ӥ�<\��<��<��<�8�<Y�<�v�<���<G��<y��<;��<{��<��<�<.�<c�<��<��<��<0�<E�<� �<���<J��<���<q��<��<�g�<�?�<�<���<5��<+v�<�8�<O��<l��<�c�<��<���<e�<��<g��<�;�<���<�]�<��<om�<s�<k�<K�<4W�<�ƴ<o2�<���<���<\]�<Z��<��<�f�<K��<��<�Q�<ՙ�<%ߠ<�!�<{a�<ʞ�<�ٙ<v�<
I�<�}�<9��<�<C�<�=�</j�<��<Ӿ�<r�<�<�5�<�[�<�}<vLy<k�u<��q<�%n<1mj<�f<��b<pE_<��[<��W<�#T<HpP<7�L<I<�_E<��A<
><c:<�6<�3<�/<��+<�O(<9�$<M/!<��<!<Q�<�&<�<�B<��<�v<-<���;���;�[�;���;�i�;��;���;�t�;�D�;�%�;��;�;�2�;�[�;Ж�;U�;�F�;7��;�B�;�݊;鋅;M�;!Dv;�l;F	b;�$X;0eN;�D;{T;;�2;��(;��;	�;�;�m;���:���:�b�:��:�:S��:�F�:�ň:F�r:
�T:��6:E: &�9Ei�9�L�9��9��&8r����2�q����Ź�������?2�RL�*3f����7���*c��)�����������)_˺ܳ׺��㺳1��Z���<��D
�zH�aF��?�4"��$(�X.���3���9���?�H�E���K��^Q�y9W�k]��b��h���n�/mt�vBz��������ⅻ͈�0�������k���?���o���^���  �  �v=�= �=u[=��=�= >=�� =�~ =} =|�<n��<"��<5�<dq�<���<P��<� �<�Y�<e��<��<���<,2�<|e�<w��<,��<~��<a%�<�Q�<�|�<٥�<S��<��<�<9�<Y�<�v�<ɒ�<>��<{��<B��<���<.��<�<2�<`�<��<��<��<$�<<�<� �<���<P��<���<i��<��<�g�<�?�<�<���<+��<!v�<y8�<G��<q��<�c�<��<���<e�<��<p��<�;�<���<�]�<��<nm�<y�<k�<I�<+W�<�ƴ<x2�<��<���<W]�<c��<��<�f�<@��<��<�Q�<͙�<ߠ<�!�<ta�<���<�ٙ<g�<�H�<�}�<.��<�<;�<�=�<'j�<��<о�<s�<!�<�5�<\�<�}<�Ly<g�u<��q<�%n<Qmj<�f<�b<�E_<��[<��W<�#T<NpP<m�L<
I<�_E<��A<
><c:<ʾ6<�3<�/<��+<�O(<9�$<2/!<��<!<.�<�&<�<�B<��<�v<<���;��;�[�;���;�i�;��;^��;�t�;�D�;Y%�;��;N�;�2�;�[�;��;��;�F�;?��;�B�;�݊;'��;\M�;BDv;�l;M	b;�$X;�dN;��D;1T;;�2;��(;�;��;S;�m;���:��:�b�:x�:k�:���:F�:ň:��r:��T:`�6:D:�(�9Qm�9�N�9�9.�&8m����2�ͺ��Ź��������@2�@QL�2f����S����c������M���j����_˺��׺��32�G[���<�4E
�I�:F�@��4"��$(��.���3��9���?���E�t�K��^Q�r9W�Z]�\�b���h�P�n��lt��Bz��������ᅻ͈�����*�������Q����n���^���  �  �v=�=�=z[=��=y�=(>=�� =�~ =} = |�<c��<��<5�<Sq�<���<H��<� �<�Y�<m��<#��<���<=2�<ne�<z��<0��<���<b%�<�Q�<�|�<٥�<m��<��<�<9�<
Y�<w�<���<Q��<���<@��<���<"��<�<0�<n�<��<��<��<�<N�<� �<���<>��<���<c��<��<�g�<�?�<�<���<<��<!v�<�8�<M��<g��<�c�<��<���<e�<��<o��<�;�<��<�]�<��<nm�<�<k�<L�<EW�<�ƴ<z2�<���<���<[]�<e��<��<�f�<N��<��<�Q�<ٙ�<ߠ<�!�<ja�<Ş�<�ٙ<j�<�H�<}�<%��<�<J�<�=�<4j�<��<ξ�<�<�<�5�<�[�<�}<�Ly<��u<��q<�%n<fmj<�f<$�b<�E_<��[<��W<�#T<KpP<V�L<I<�_E<ǳA<
><�b:<�6<�3<�/<��+<uO(<!�$<(/!<��<� <H�<�&<۱<�B<��<�v<<Ј�;���;�[�;��;�i�;��;)��;�t�;�D�;�%�;��;\�;�2�;�[�;9��;o�;�F�;R��;�B�;�݊;���;}M�;/Dv;�l;	b;�$X;DeN;��D;�T;;z2;c�(;x�;��; ;:m;|��:��:Mb�:�:n�:���:�F�:pň:��r:"�T:Y�6:�D:&�9�j�9UN�9��9�&8���ٽ2����s�Ź�������=2�/QL��1f��������Wc��}������A����^˺��׺���1�[���<�E
��H��F��?��4"�Q%(��.���3���9�	�?�!�E���K��^Q�9W�u]�'�b��h�_�n��lt�Bz���������ᅻ&͈�и��D���L������	o���^���  �  �v=�= �=u[=��=u�=%>=� =�~ =w =|�<j��<��<5�<:q�<���<?��<� �<�Y�<a��<��<���<82�<he�<���<&��<���<r%�<�Q�<�|�<ץ�<g��<#��<�<9�<Y�<w�<���<\��<z��<O��<���<&��<%�<*�<l�<��<��<��<�<B�<� �< ��<9��<���<[��<���<�g�<�?�<�<���<1��<v�<r8�<H��<h��<�c�<��<˾�<e�<��<���<�;�<��<�]�<��<{m�<��<k�<N�<DW�<�ƴ<�2�<��<���<e]�<Z��<��<�f�<K��<{�<�Q�<Ι�<ߠ<�!�<aa�<Ş�<�ٙ<h�<�H�<�}�<6��<���<?�<�=�<+j�<��<ؾ�<v�<�<�5�<�[�<�}<�Ly<v�u<��q<�%n<{mj<)�f<7�b<�E_<Ŏ[<��W<�#T<|pP<L�L<4I<�_E<��A<
><�b:<޾6<�3<�/<��+<�O(<0�$</!<��<� <G�<�&<��<�B<y�<�v<�<���;���;�[�;���;�i�;�;%��;Vu�;�D�;�%�;�;\�;�2�;�[�;\��;g�;G�;8��;C�;ފ;��;�M�;�Cv;�l;*	b;]$X;�dN;��D;^T;;2;�(;Q�;��;�;�l;g��:���:�c�:Q�:��:���:�E�:ň:��r:8�T:!�6:�F:>(�9�n�9.S�9��9�'8<���2�����ՔŹ���Y���=2��QL�/f���������b��8���h���v���6_˺��׺���*2��[��x<��E
��H�WG�@��4"�3%(�l.�J�3���9���?�g�E��K��^Q�U9W��]���b�?�h���n��lt�KBz��������xᅻ�̈�����V���0���%����n���^���  �  �v=�="�=t[=��=x�=#>=�� =�~ =y =�{�<_��<��<5�<Mq�<���<;��<� �<�Y�<f��<#��<���<-2�<re�<~��<+��<���<]%�<�Q�<�|�<��<d��<3��<�<9�<Y�<w�<Ԓ�<W��<���<D��<���<#��<�<5�<f�<��<��<��<$�<K�<� �<���<5��<���<_��< ��<�g�<�?�<�<���<8��<"v�<~8�<D��<r��<�c�<��<���<e�<��<s��<�;�<��<�]�<��<wm�<��<#k�<a�<?W�<�ƴ<~2�<��<���<Z]�<b��<��<�f�<C��<��<�Q�<ә�<	ߠ<�!�<^a�<���<�ٙ<g�<�H�<y}�<!��< �<E�<�=�<+j�<��<ھ�<s�<%�<�5�<�[�<�}<�Ly<}�u<��q<�%n<hmj<�f<$�b<�E_<Ԏ[<��W<�#T<XpP<X�L<I<�_E<��A<
><�b:<־6<�3<�/<��+<fO(<�$</!<��<� <?�<�&<ұ<�B<��<�v<<���;���;�[�;���;�i�;��;4��;u�;�D�;�%�;A�;y�;�2�;�[�;>��;��;G�;S��;�B�;�݊;���;mM�;MDv;�l;p	b;J$X;�dN;��D;�T;;�2;T�(;*�;s�;�;m;���:v��:b�:!�:*�:���:ZF�:�Ĉ:��r:q�T:��6:�D:&�9�k�9O�9 �9G�&8s����2������Ź�������>2�[PL�l1f���ŵ��nc������ꄲ������_˺W�׺����1�\��=��E
��H��F�@��4"�%(�.�>�3���9���?�g�E�݂K��^Q�p9W�;]�^�b��h�*�n��lt�.Bz����q����ᅻ͈�и������������n���^���  �  �x=�=|�=$^=��=۠=�A=�� =
� =J# =T��<���<��<�A�<�~�<��<���<1�<�j�<h��<���<��<G�<|{�<��<X��<��<�?�<em�<Q��<���<w��<��<�8�<\�<\}�<���<ȹ�<���<O��<t�< �<?(�<z6�<!B�<�J�<WP�<�R�<R�<�M�<zF�<�;�<�,�<w�<�<���<���<6��<���<�W�<c(�<z��<��<�<\=�<���<���<�[�<��<4��<�N�<1��<��<��<��<�-�<]��<�2�<'��<J%�<��<��<�p�<�ֱ<9�<=��<��<oH�<���<p�<�7�<1��<�Ǣ<�
�<{K�<y��<�ě<���<�4�<#i�<ě�<a̒<T��<x(�<(T�<z~�<v��<9χ<���<��<W@�<�d�<�}<�Uy<��u<��q<#n<�fj<��f<��b<A3_<ex[<��W<�T<FNP<��L<�H<2E<�A<T�=<^):<#�6<
�2<P:/<g�+<(<�k$<�� <jL<��<L@<F�<�I<��<�i</<Q�<X��;L��;=Z�;���; \�;���;ٝ�;W�;O"�;*��;��;�;0 �;&�;�^�;��;R
�;�}�;y�;잉;MM�;O~;�s;s�i;��_;��U;)�K;�bB;P�8;�/;p�&;|~;��;��;�?;S��:��:H�:9�:���:&�:��:!�:��k:��M:�0:��:#��9..�9��r9��9U��7����G����FϹ�*��z�Җ6�~zP��5j��ށ�#����*��o���/(��'����̺b$ٺ�Z庽��^�������
����(��޻���"��(��y.�\4��<:��@���E���K���Q�wW�(J]�3c���h�0�n�3�t��_z�%��- ���腻rш�Ѻ������<���yz��tf�� T���  �  �x=�=y�= ^=��=Ԡ=�A=�� =� =D# =K��<t��<��<�A�<�~�<��<v��<1�<�j�<`��<��<��< G�<n{�<���<G��<��<�?�<Nm�<P��<���<���<��<�8�<	\�<Y}�<���<Ϲ�<���<A��<q�<�<+(�<�6�<B�<�J�<QP�<�R�<R�<N�<�F�<z;�<�,�<]�<�<���<���<>��<���<�W�<R(�<���<*��<!�<\=�<���<���<�[�<��<$��<�N�<-��<��<��<(��<�-�<[��<�2�<,��<[%�<��<��<�p�<�ֱ<9�<?��<��<rH�<���<t�<8�<X��<�Ǣ<�
�<vK�<c��<�ě<���<�4�< i�<���<[̒<I��<�(�<CT�<�~�<i��<3χ<���<��<b@�<ud�<�}<�Uy<��u<�q<
#n<�fj<��f<��b<E3_<�x[<��W<�T<=NP<Y�L<-�H<�1E<߁A<P�=<A):<2�6<=�2<�:/<P�+<�(<�k$<�� <xL<��<a@<�<wI<��<�i<{<�<g��;��;FZ�;h��;!\�;���;}��;W�;�!�;f��;��;*�;3 �;�%�;�^�;/��;�
�;�}�;j�;ƞ�;M�;�~;��s;��i;{�_;��U;��K;�cB;��8;��/;D�&;�};��;��;�?;у�:P��:�G�:+�:H��::(�:��:"!�:��k:l�M:�0:��: ��9G*�9��r9�9��7Q��)�G��Ù�oFϹJ*��x�U�6�/}P��5j����U����*�������'��������̺�"ٺ3X��� ���>����
����k�����ĩ"�˓(��y.�e\4��;:��@�K�E�	�K�-�Q�>wW��J]��c�c�h�T�n���t��_z����" ���腻�ш�������������wz���f��T���  �  �x=�=w�=!^=��=ՠ=�A=�� =� =A# =g��<���<��<�A�<�~�<��<x��<1�<�j�<V��<��<��<)G�<i{�<���<B��<��<�?�<Jm�<g��<���<���<|�<�8�<\�<V}�<���<���<���<5��<|�<!�<'(�<�6�<B�<�J�<LP�<�R�<R�<�M�<�F�<v;�<�,�<`�<1�<���<���<T��<���<�W�<T(�<y��<��<�<h=�<���<«�<�[�<��<"��<�N�<;��<��<��<��<�-�<Z��<�2�<��<?%�<��<w�<�p�<�ֱ<9�<E��<��<|H�<���<~�<�7�<D��<�Ǣ<�
�<�K�<c��<�ě<���<�4�<0i�<���<x̒<B��<�(�<)T�<�~�<n��<2χ<���<��<r@�<pd�<�}<�Uy<��u<�q<�"n<�fj<��f<��b<3_<rx[<{�W<�T<hNP<K�L<G�H<�1E<�A<R�=<E):<<�6<�2<n:/<D�+<*(<�k$<�� <�L<��<�@<$�<�I<��<�i<[<K�<���;��;jZ�;W��;0\�;���;n��;rW�;�!�;^��;u�;��;$ �;�%�;�^�;���;�
�;s}�;��;�;�L�;
~;8�s;Кi;T�_;�U;;�K;cB;��8;k�/;.�&;�};c�;��;�?;1��:D��:�I�:Q�:���:�&�:&��:�!�:��k:��M:�0:1�:���9,�9��r9p�9�7�.����G��Ù��FϹ,�a|���6��~P�43j�/������<*�����W'��V���,�̺t$ٺkY庫����������
������r��B�"��(��x.��\4�%<:�y@�R�E���K�7�Q�wW��J]�_c���h�ɾn���t�(`z����~ ���腻�ш�����פ��!����z���f���S���  �  �x=�=v�=%^=��=۠=�A=�� =� =H# =\��<}��<�<�A�<�~�<��<���<1�<�j�<j��<��<��</G�<m{�<���<N��<��<�?�<Im�<Q��<���<���<��<�8�<�[�<I}�<���<���<���<>��<k�<�<&(�<�6�<B�<�J�<IP�<�R�<R�<N�<�F�<�;�<�,�<f�<&�<���<���<J��<���<�W�<Y(�<���<&��<�<p=�<���<«�<�[�<��<��<�N�<'��<��<��<��<�-�<K��<y2�</��<F%�<��<~�<�p�<�ֱ< 9�<9��<��<xH�<���<��<�7�<U��<�Ǣ<�
�<|K�<o��<�ě<���<�4�<+i�<���<j̒<L��<�(�<;T�<�~�<{��<.χ<���<��<]@�<pd�<�}<�Uy<��u<��q<�"n<�fj<o�f<��b<B3_<kx[<��W<�T<ANP<N�L< �H<�1E<�A<F�=<[):<?�6<&�2<�:/<a�+<(<�k$<�� <�L<��<t@<:�<�I<��<�i<~<e�<���;��;[Z�;���;\�;���;o��;W�;�!�;U��;��;?�;���;�%�;�^�;쪟;�
�;�}�;W�;���;�L�;�~;��s;�i;9�_;6�U;Y�K;�cB;A�8;��/;��&;�};�;��;�?;���:���:H�:��:��:(�:���:c"�:��k:��M:�0:{�:��9�(�9
�r9��9�͛7-#����G�Ǚ�[JϹ�)�T{��6��}P��5j�u���Ï���*��=����'��;�����̺�#ٺZX�J��c�����D�
�D��)�����g�"�h�(�my.�I\4��;:��@�I�E�w�K�[�Q��vW��J]�
c���h�i�n���t��_z���9 ���腻�ш�溋�����/����z���f��	T���  �  �x=�=y�="^=��=۠=�A=�� =� =J# =`��<���<�<�A�<�~�<��<���<1�<�j�<g��<��<��<G�<v{�<���<K��<��<�?�<Um�<E��<���<r��<s�<�8�<�[�<O}�<���<���<���<=��<i�<�<2(�<6�<B�<�J�<TP�<�R�<R�<N�<�F�<�;�<�,�<��<(�<���<���<H��<�<�W�<d(�<���<)��<�<c=�<���<���<�[�<��<(��<�N�<#��<��<��<��<{-�<K��<s2�<��<=%�<���<��<�p�<�ֱ<9�<9��<��<qH�<���<t�<�7�<V��<�Ǣ<�
�<�K�<���<�ě<���<�4�<6i�<Л�<o̒<U��<�(�<GT�<r~�<x��<3χ<���<��<Z@�<|d�<�}<�Uy<��u<��q<�"n<�fj<��f<��b<'3_<@x[<s�W<�T<-NP<e�L< �H<�1E<�A<L�=<^):<�6<?�2<�:/<h�+<(<�k$<� <�L< �<f@<n�<�I<��<�i<~<y�<`��;8��;LZ�;~��;\�;���;���;�V�;�!�;��;V�;��;���;�%�;�^�;窟;4
�;�}�;O�;���;M�;|~;��s;��i;��_;�U;�K;�cB;��8;�/;ځ&;�~;&�;g�;�@;���:���:�H�:W�:1��:=(�:8��:�!�:7�k:��M:(0:?�:���92*�9Y�r98�9�w�7$����G��ƙ��KϹ�,�j|�Q�6�Z}P�7j��߁�`����*��{����'�������̺m#ٺ;X庤��ך�����h�
�v�����j��
�"���(�Ey.�\4��;:��@���E���K�0�Q�wW�uJ]� c�/�h���n���t�`z�f��c ��酻�ш����ä�������z���f��1T���  �  �x=�=x�=#^=��=ܠ=�A=�� =� =O# =q��<���<�<�A�<�~�<$��<���<1�<�j�<m��<��<��<*G�<x{�<���<K��<��<�?�<@m�<I��<���<t��<w�<�8�<�[�<N}�<z��<���<���<3��<_�<�<(�<�6�<B�<�J�<WP�<�R�<R�<N�<�F�<�;�<�,�<w�<6�<��<���<W��<���<�W�<w(�<���<+��<�<g=�<���<���<�[�<��<��<�N�<��<���<��<
��<g-�<M��<t2�<��<=%�<���<q�<�p�<�ֱ<�8�<>��<��<sH�<���<}�<�7�<R��<�Ǣ<�<�K�<���<�ě<���<�4�<?i�<ś�<|̒<a��<�(�<GT�<�~�<w��<7χ<���<��<Z@�<gd�<�}<�Uy<��u<��q<�"n<�fj<��f<s�b<3_<Ux[<s�W<�T<2NP<<�L<�H<�1E<�A<T�=<_):<?�6<?�2<�:/<|�+<?(<�k$<� <�L<#�<�@<d�<�I<��<�i<t<|�<���;B��;[Z�;���;)\�;u��;N��;�V�;�!�;#��;i�;��;���;�%�;N^�;˪�;W
�;s}�;+�;���;�L�;�~;��s;��i;��_;��U;��K;�cB;��8;��/;5�&;�~;��;��;~@;s��:��:yI�:��:��:k(�::�!�:_�k:��M:�0:��:���9�'�96�r9��9H��7p)���G�gƙ�WKϹ]/�N|�+�6�:P��6j� ၺ�����*�������'��o����̺F#ٺrX�l��s��������
���������Ȩ"��(��x.��[4��;:��@�<�E���K��Q�wW��J]�c���h���n�"�t�<`z�<��� ��:酻�ш�A�������[����z���f��$T���  �  �x=�=s�="^=��=٠=�A=�� =#� =M# =p��<���< �<�A�<�~�<4��<���<$1�<�j�<s��<-��<��<2G�<p{�<���<G��<��<�?�<Fm�<J��<���<g��<h�<�8�<�[�<2}�<���<���<���<+��<X�<�<(�<�6�<B�<�J�<QP�<�R�< R�<N�<�F�<�;�<�,�<��<D�<��<���<f��<Ă�<�W�<n(�<���<6��< �<l=�<���<���<�[�<��<��<�N�<��<ׂ�<��<���<q-�<0��<_2�<	��<.%�<<g�<�p�<�ֱ<�8�<2��<��<vH�<���<��<�7�<d��<�Ǣ<�<�K�<���<�ě<���<�4�<Ii�<ԛ�<̒<\��<�(�<LT�<�~�<u��<3χ<���<��<^@�<gd�<�}<kUy<l�u<��q<�"n<�fj<N�f<o�b<3_<*x[<X�W<�T<?NP<;�L<#�H<�1E<�A<N�=<T):<P�6<E�2<�:/<w�+<>(<�k$<&� <�L<#�<�@<y�<�I<��<j<�<��<���;(��;fZ�;v��; \�;���;i��;W�;�!�;���;/�;��;���;g%�;|^�;���;
�;R}�;�;Ş�;�L�;�~;M�s;Ți;��_;�U;��K;8dB;��8;o�/;n�&;�~;�;��;�@;v��:���:J�:�:w��:)�:%��:K"�:��k:}�M:�0:a�:��9*�9��r9U�9�X�7:7����G�O͙�TPϹF.�~�̘6�b�P�17j�x���K���@+��Ͳ���'������̺�"ٺUW������G��_�
�I�����ĺ�s�"���(��x.��[4�&;:�b@���E���K�2�Q�wW��J]��c���h�S�n�t�t��`z����� ��,酻҈�H�����������z��'g��
T���  �  �x=�=v�=#^=��=ޠ=�A=�� = � =S# =~��<���<!�<�A�<�<.��<���<91�<�j�<}��<%��<��</G�<{{�<���<K��<��<�?�<@m�<0��<���<c��<Z�<�8�<�[�</}�<t��<���<~��<2��<J�<�<(�<x6�<B�<�J�<VP�<�R�<R�<N�<�F�<�;�<�,�<��<:�<��<���<\��<҂�<�W�<w(�<���<+��<�<q=�<���<���<�[�<��<��<~N�<��<ނ�<��<<`-�<+��<X2�<���<%�<闶<m�<�p�<�ֱ<�8�</��<��<sH�<���<��<�7�<[��<�Ǣ<�<�K�<���<�ě<��<�4�<Ei�<䛔<�̒<g��<�(�<GT�<�~�<���<6χ<���<��<V@�<dd�<�}<cUy<{�u<��q<�"n<lfj<Q�f<R�b<�2_<x[<^�W<�T<NP<5�L<�H<�1E<�A<S�=<j):<E�6<D�2<�:/<��+<Z(<&l$<)� <�L<[�<�@<��<�I<��<j<�<��<���;X��;cZ�;���;\�;v��;W��;�V�;�!�;���;��;��;{��;`%�;9^�;u��;�	�;s}�;��;���;�L�;R~;��s;��i;��_;l�U;��K;�cB;��8;��/;ׂ&;a;��;`�;wA;؅�:���:�J�:��:���:t(�:��:�"�:_�k:��M:�0:\�:��9'�9��r9C�9�-�70C���G�BΙ��QϹ�/���r�6��P��:j���������i+�������'��M�����̺#ٺ�W�=�J������
�
�������g����"�
�(�^x.�q[4�>;:��@�/�E�U�K��Q�wW��J]�@c���h��n���t�b`z����� ��l酻҈�����1���ޏ���z��g��iT���  �  �x=�=v�=!^=��=ޠ=�A=�� =� =\# =|��<���</�<�A�<	�<;��<���<.1�<�j�<���<$��<��<-G�<}{�<���<G��<��<�?�<@m�<7��<���<V��<d�<�8�<�[�<3}�<`��<���<{��<��<G�<�<(�<q6�<B�<�J�<XP�<�R�<1R�<$N�<�F�<�;�<�,�<��<N�<��<���<n��<Ղ�<�W�<�(�<���<7��<3�<l=�<���<���<�[�<��<��<|N�< ��<Ȃ�<��<���<O-�<-��<S2�<�<)%�<ݗ�<\�<�p�<�ֱ<�8�<.��<��<pH�<���<��<8�<^��<�Ǣ<�<�K�<���<�ě<	��<�4�<Wi�<ݛ�<�̒<w��<�(�<\T�<�~�<~��<6χ<���<��<G@�<cd�<�}<VUy<O�u<��q<�"n<Ffj<M�f<3�b<�2_<#x[<:�W<xT<NP<6�L<��H<�1E<�A<Q�=<i):<R�6<m�2<�:/<��+<X(<l$<G� <�L<c�<�@<��<�I<�<=j<�<��<���;_��;_Z�;}��;\�;1��;V��;�V�;!�;���;&�;m�;`��;o%�;�]�;���;�	�;}�;��;���;�L�;~;��s;��i;ē_;:�U;8�K;sdB;��8;&�/;Ȃ&;k;`�;M�;cA;���:��:�J�:f�:&��:@)�:o��:R"�:��k:��M:�0:��:�~�9�&�9��r9�9L�709��+�G��͙��RϹ�1�x~���6���P��9j�ၺ����k+�������'�������̺�!ٺ�W庄~����������
������F����"�A�(�kx.��Z4�d;:��@���E�_�K��Q�+wW��J]��c���h��n�ʐt�az����� ���酻҈�����7�������{��Bg��^T���  �  �x=�=t�= ^=��=ܠ=�A=�� =$� =[# =���<���<?�<�A�<�~�<N��<���<F1�<�j�<���<(��<��<0G�<x{�<���<A��<��<�?�<4m�<@��<���<Q��<L�<~8�<�[�< }�<f��<���<r��<��<O�<�<(�<�6�< B�<�J�<[P�<�R�<*R�<N�<�F�<�;�<-�<��<h�<��<���<���<ׂ�<�W�<�(�<���<0��<*�<l=�<���<���<�[�<��<��<xN�<��<���<��<ۣ�<Q-�<��<D2�<筹<%�<֗�<P�<�p�<�ֱ<�8�<6��<��<zH�<���<��<	8�<]��<�Ǣ<�<�K�<���<ś<���<�4�<ji�<훔<�̒<u��<�(�<PT�<�~�<{��<:χ<���<��<Z@�<Xd�<�}<YUy<@�u<��q<�"n<Vfj<&�f<>�b<�2_<�w[<-�W<uT<NP<�L<�H<�1E<߁A<Z�=<a):<O�6<U�2<�:/<��+<i(<:l$<f� <�L<G�<�@<��< J<�<<j<�<��<���;P��;�Z�;e��;'\�;u��;+��;�V�;Z!�;���;��;I�;A��;&%�;^�;3��;�	�;�|�;��;���;�L�;�~;2�s;Ӛi;ߓ_;8�U;�K;2dB;��8;	�/;\�&;�;2�;q�;pA;���:,��:�K�:C�:y��:�(�:狔:c"�:��k:��M:0:p�:z�9�%�9��r9΃9X��7�U����G�ҙ�zVϹ"2����6���P�08j��ၺِ���*��T���6'��[�����̺G"ٺ�W�c~񺪘��E����
�g�������g�"�(�x.�[4� ;:�>@���E�w�K���Q�wW��J]�!c�L�h�ܿn���t�Oaz����$���酻n҈������������/{��Hg��TT���  �  |x=�=o�=#^=��=ޠ=�A=�� =.� =Z# =���<���<,�<B�<
�<S��<���<K1�<�j�<���<=��<��<EG�<t{�<���<D��<��<�?�<"m�<+��<���<`��<H�<�8�<�[�<}�<m��<~��<���<��<9�<��<(�<x6�< B�<�J�<NP�<�R�<2R�<"N�<�F�<�;�<
-�<��<W�<,��<���<}��<̂�<�W�<w(�<���<:��<.�<y=�<���<���<�[�<��<���<eN�<���<���<��<ϣ�<Y-�<��<B2�<�<%�<时<F�<�p�<�ֱ<�8�<*��<��<vH�<���<��<	8�<p��<�Ǣ<�<�K�<���<ś<��<�4�<Ui�<뛔<�̒<p��<�(�<PT�<�~�<���</χ<���<{�<U@�<Jd�<�}<4Uy<U�u<��q<u"n<bfj<��f<E�b<�2_<x[<C�W<UT<�MP<�L<�H<�1E<�A<K�=<i):<s�6<S�2<�:/<��+<f(<?l$<A� <M<g�<�@<��<J<�<Ij<�<��<��;A��;tZ�;s��;�[�;n��;��;�V�;4!�;���;��;h�;L��;�$�;&^�; ��;
�;}�;��;G��;tL�;]~;/�s;�i;��_;��U;L�K;edB;��8;ʩ/;~�&;R;��;��;�A;���:w��:8L�:��:���:t)�:,��:<#�:G�k:��M:60:��:�}�9K!�9��r9�9�7�7a��X�G��ԙ��VϹ�0�u����6�=�P�	;j��⁺����+�����k'�������̺A"ٺsV床}�=������
�m���������"�Б(��w.�+[4�M::�C@�o�E�F�K�Q�Q��vW�K]�Ic���h�a�n�P�t��`z����J��~酻�҈�������������{���g���T���  �  �x=�=o�="^=��=ߠ=�A=�� ="� =\# =���<���<>�<B�<�<T��<���<P1�<�j�<���<-��<��<6G�<|{�<���<G��<��<�?�<<m�<9��<���<D��<@�<s8�<�[�<}�<Z��<��<j��<��<E�<�<(�<n6�<B�<�J�<UP�<�R�<0R�<!N�<�F�<�;�<-�<��<d�<+��<���<���<��<�W�<�(�<���<5��</�<p=�<���<���<�[�<��<��<{N�<���<���<��<У�<D-�<��<?2�<ܭ�<%�<ɗ�<K�<�p�<�ֱ<�8�<!��<��<mH�<���<��<8�<d��<�Ǣ<�<�K�<���<ś<��<�4�<hi�<���<�̒<x��<�(�<UT�<�~�<���<2χ<���<�<M@�<ed�<�}<EUy<&�u<|�q<o"n<Afj<�f<)�b<�2_<�w[<�W<aT<NP<7�L<�H<�1E<�A<H�=<m):<\�6<b�2<�:/<��+<s(<Yl$<f� <
M<t�<�@<��<J<�<Hj<�<��<Ք�;b��;WZ�;���;�[�;~��;L��;�V�;R!�;r��;��;!�;2��;%�;�]�;��;�	�;�|�;��;���;�L�;~;e�s;��i;��_;l�U;7�K;_dB;��8;<�/;��&;C�;�;��;�A;���:���:gL�:��:���:')�:5��:�"�:��k:t�M:0:�:��9�&�9��r9�9dǚ7=_����G��ә�xWϹr3���)�6���P��9j�2ၺ����/,��ٲ���'��<���i�̺�!ٺ4W�~�}������,�
�X��b�����}�"�;�(��w.��Z4�;:�@���E�N�K�9�Q�1wW��J]��c���h��n��t��az���V���酻�҈�ӻ������,���m{��pg��YT���  �  }x=�=w�="^=��=�=�A=�� =$� =e# =���<���<=�<B�<�<L��<���<<1�<�j�<���<2��<��<+G�<�{�<���<M��<��<�?�<m�< ��<���<G��<W�<t8�<�[�< }�<Q��<���<o��<��<E�<��<(�<j6�<B�<�J�<hP�<�R�<6R�<7N�<�F�<�;�<�,�<��<_�<+��<���<��<߂�<�W�<�(�<���<G��<<�<i=�<��<���<�[�<��<���<WN�<���<Ă�<��<룿<<-�<��<=2�<٭�<%�<͗�<Z�<�p�<�ֱ<�8�<)��<��<mH�<Û�<{�<"8�<k��<�Ǣ<%�<�K�<���<
ś<��<�4�<fi�<월<�̒<���<�(�<mT�<�~�<���<@χ<���<��<H@�<Nd�<V}<XUy<<�u<��q<�"n<0fj<)�f<�b<�2_<
x[< �W<wT<�MP<�L<��H<�1E<�A<[�=<t):<J�6<��2<�:/<՜+<l(<8l$<d� <M<|�<�@<��<�I<+�<Zj<�<أ<���;���;hZ�;���;\�;[��;؜�;mV�;�!�;���;��;"�;��;*%�;�]�;e��;�	�;}�;��;���;tL�;�~;��s;��i;K�_;N�U;k�K;eB;�8;�/;�&;�;�;��;�A;"��:���:�J�:��:���:T*�:��:A"�:��k:��M:.0:��:r}�9��9��r9��9 ۚ7�C��ͱG��ҙ��WϹ�3�����6���P�
<j�;ぺ/����+��y����'��8����̺� ٺ�V庿}񺴗�����^�
����F�������"�ɑ(�4x.�FZ4��::�Y@���E�H�K�ɡQ�?wW��J]��c���h��n���t�\az�������酻f҈�򻋻����폑�I{��Cg���T���  �  �x=�=o�="^=��=ߠ=�A=�� ="� =\# =���<���<>�<B�<�<T��<���<P1�<�j�<���<-��<��<6G�<|{�<���<G��<��<�?�<<m�<9��<���<D��<@�<s8�<�[�<}�<Z��<��<j��<��<E�<�<(�<n6�<B�<�J�<UP�<�R�<0R�<!N�<�F�<�;�<-�<��<d�<+��<���<���<��<�W�<�(�<���<5��</�<p=�<���<���<�[�<��<��<{N�<���<���<��<У�<D-�<��<?2�<ܭ�<%�<ɗ�<K�<�p�<�ֱ<�8�<!��<��<mH�<���<��<8�<d��<�Ǣ<�<�K�<���<ś<��<�4�<hi�<���<�̒<x��<�(�<UT�<�~�<���<2χ<���<�<M@�<ed�<�}<EUy<&�u<|�q<o"n<Afj<�f<)�b<�2_<�w[<�W<aT<NP<7�L<�H<�1E<�A<H�=<m):<\�6<b�2<�:/<��+<s(<Yl$<f� <
M<t�<�@<��<J<�<Hj<�<��<Ք�;b��;WZ�;���;�[�;~��;L��;�V�;R!�;r��;��;!�;2��;%�;�]�;��;�	�;�|�;��;���;�L�;~;e�s;��i;��_;l�U;7�K;_dB;��8;<�/;��&;C�;�;��;�A;���:���:gL�:��:���:')�:5��:�"�:��k:t�M:0:�:��9�&�9��r9�9dǚ7=_����G��ә�xWϹr3���)�6���P��9j�2ၺ����/,��ٲ���'��<���i�̺�!ٺ4W�~�}������,�
�X��b�����}�"�;�(��w.��Z4�;:�@���E�N�K�9�Q�1wW��J]��c���h��n��t��az���V���酻�҈�ӻ������,���m{��pg��YT���  �  |x=�=o�=#^=��=ޠ=�A=�� =.� =Z# =���<���<,�<B�<
�<S��<���<K1�<�j�<���<=��<��<EG�<t{�<���<D��<��<�?�<"m�<+��<���<`��<H�<�8�<�[�<}�<m��<~��<���<��<9�<��<(�<x6�< B�<�J�<NP�<�R�<2R�<"N�<�F�<�;�<
-�<��<W�<,��<���<}��<̂�<�W�<w(�<���<:��<.�<y=�<���<���<�[�<��<���<eN�<���<���<��<ϣ�<Y-�<��<B2�<�<%�<时<F�<�p�<�ֱ<�8�<*��<��<vH�<���<��<	8�<p��<�Ǣ<�<�K�<���<ś<��<�4�<Ui�<뛔<�̒<p��<�(�<PT�<�~�<���</χ<���<{�<U@�<Jd�<�}<4Uy<U�u<��q<u"n<bfj<��f<E�b<�2_<x[<C�W<UT<�MP<�L<�H<�1E<�A<K�=<i):<s�6<S�2<�:/<��+<f(<?l$<A� <M<g�<�@<��<J<�<Ij<�<��<��;A��;tZ�;s��;�[�;n��;��;�V�;4!�;���;��;h�;L��;�$�;&^�; ��;
�;}�;��;G��;tL�;]~;/�s;�i;��_;��U;L�K;edB;��8;ʩ/;~�&;R;��;��;�A;���:w��:8L�:��:���:t)�:,��:<#�:G�k:��M:60:��:�}�9K!�9��r9�9�7�7a��X�G��ԙ��VϹ�0�u����6�=�P�	;j��⁺����+�����k'�������̺A"ٺsV床}�=������
�m���������"�Б(��w.�+[4�M::�C@�o�E�F�K�Q�Q��vW�K]�Ic���h�a�n�P�t��`z����J��~酻�҈�������������{���g���T���  �  �x=�=t�= ^=��=ܠ=�A=�� =$� =[# =���<���<?�<�A�<�~�<N��<���<F1�<�j�<���<(��<��<0G�<x{�<���<A��<��<�?�<4m�<@��<���<Q��<L�<~8�<�[�< }�<f��<���<r��<��<O�<�<(�<�6�< B�<�J�<[P�<�R�<*R�<N�<�F�<�;�<-�<��<h�<��<���<���<ׂ�<�W�<�(�<���<0��<*�<l=�<���<���<�[�<��<��<xN�<��<���<��<ۣ�<Q-�<��<D2�<筹<%�<֗�<P�<�p�<�ֱ<�8�<6��<��<zH�<���<��<	8�<]��<�Ǣ<�<�K�<���<ś<���<�4�<ji�<훔<�̒<u��<�(�<PT�<�~�<{��<:χ<���<��<Z@�<Xd�<�}<YUy<@�u<��q<�"n<Vfj<&�f<>�b<�2_<�w[<-�W<uT<NP<�L<�H<�1E<߁A<Z�=<a):<O�6<U�2<�:/<��+<i(<:l$<f� <�L<G�<�@<��< J<�<<j<�<��<���;P��;�Z�;e��;'\�;u��;+��;�V�;Z!�;���;��;I�;A��;&%�;^�;3��;�	�;�|�;��;���;�L�;�~;2�s;Ӛi;ߓ_;8�U;�K;2dB;��8;	�/;\�&;�;2�;q�;pA;���:,��:�K�:C�:y��:�(�:狔:c"�:��k:��M:0:p�:z�9�%�9��r9΃9X��7�U����G�ҙ�zVϹ"2����6���P�08j��ၺِ���*��T���6'��[�����̺G"ٺ�W�c~񺪘��E����
�g�������g�"�(�x.�[4� ;:�>@���E�w�K���Q�wW��J]�!c�L�h�ܿn���t�Oaz����$���酻n҈������������/{��Hg��TT���  �  �x=�=v�=!^=��=ޠ=�A=�� =� =\# =|��<���</�<�A�<	�<;��<���<.1�<�j�<���<$��<��<-G�<}{�<���<G��<��<�?�<@m�<7��<���<V��<d�<�8�<�[�<3}�<`��<���<{��<��<G�<�<(�<q6�<B�<�J�<XP�<�R�<1R�<$N�<�F�<�;�<�,�<��<N�<��<���<n��<Ղ�<�W�<�(�<���<7��<3�<l=�<���<���<�[�<��<��<|N�< ��<Ȃ�<��<���<O-�<-��<S2�<�<)%�<ݗ�<\�<�p�<�ֱ<�8�<.��<��<pH�<���<��<8�<^��<�Ǣ<�<�K�<���<�ě<	��<�4�<Wi�<ݛ�<�̒<w��<�(�<\T�<�~�<~��<6χ<���<��<G@�<cd�<�}<VUy<O�u<��q<�"n<Ffj<M�f<3�b<�2_<#x[<:�W<xT<NP<6�L<��H<�1E<�A<Q�=<i):<R�6<m�2<�:/<��+<X(<l$<G� <�L<c�<�@<��<�I<�<=j<�<��<���;_��;_Z�;}��;\�;1��;V��;�V�;!�;���;&�;m�;`��;o%�;�]�;���;�	�;}�;��;���;�L�;~;��s;��i;ē_;:�U;8�K;sdB;��8;&�/;Ȃ&;k;`�;M�;cA;���:��:�J�:f�:&��:@)�:o��:R"�:��k:��M:�0:��:�~�9�&�9��r9�9L�709��+�G��͙��RϹ�1�x~���6���P��9j�ၺ����k+�������'�������̺�!ٺ�W庄~����������
������F����"�A�(�kx.��Z4�d;:��@���E�_�K��Q�+wW��J]��c���h��n�ʐt�az����� ���酻҈�����7�������{��Bg��^T���  �  �x=�=v�=#^=��=ޠ=�A=�� = � =S# =~��<���<!�<�A�<�<.��<���<91�<�j�<}��<%��<��</G�<{{�<���<K��<��<�?�<@m�<0��<���<c��<Z�<�8�<�[�</}�<t��<���<~��<2��<J�<�<(�<x6�<B�<�J�<VP�<�R�<R�<N�<�F�<�;�<�,�<��<:�<��<���<\��<҂�<�W�<w(�<���<+��<�<q=�<���<���<�[�<��<��<~N�<��<ނ�<��<<`-�<+��<X2�<���<%�<闶<m�<�p�<�ֱ<�8�</��<��<sH�<���<��<�7�<[��<�Ǣ<�<�K�<���<�ě<��<�4�<Ei�<䛔<�̒<g��<�(�<GT�<�~�<���<6χ<���<��<V@�<dd�<�}<cUy<{�u<��q<�"n<lfj<Q�f<R�b<�2_<x[<^�W<�T<NP<5�L<�H<�1E<�A<S�=<j):<E�6<D�2<�:/<��+<Z(<&l$<)� <�L<[�<�@<��<�I<��<j<�<��<���;X��;cZ�;���;\�;v��;W��;�V�;�!�;���;��;��;{��;`%�;9^�;u��;�	�;s}�;��;���;�L�;R~;��s;��i;��_;l�U;��K;�cB;��8;��/;ׂ&;a;��;`�;wA;؅�:���:�J�:��:���:t(�:��:�"�:_�k:��M:�0:\�:��9'�9��r9C�9�-�70C���G�BΙ��QϹ�/���r�6��P��:j���������i+�������'��M�����̺#ٺ�W�=�J������
�
�������g����"�
�(�^x.�q[4�>;:��@�/�E�U�K��Q�wW��J]�@c���h��n���t�b`z����� ��l酻҈�����1���ޏ���z��g��iT���  �  �x=�=s�="^=��=٠=�A=�� =#� =M# =p��<���< �<�A�<�~�<4��<���<$1�<�j�<s��<-��<��<2G�<p{�<���<G��<��<�?�<Fm�<J��<���<g��<h�<�8�<�[�<2}�<���<���<���<+��<X�<�<(�<�6�<B�<�J�<QP�<�R�< R�<N�<�F�<�;�<�,�<��<D�<��<���<f��<Ă�<�W�<n(�<���<6��< �<l=�<���<���<�[�<��<��<�N�<��<ׂ�<��<���<q-�<0��<_2�<	��<.%�<<g�<�p�<�ֱ<�8�<2��<��<vH�<���<��<�7�<d��<�Ǣ<�<�K�<���<�ě<���<�4�<Ii�<ԛ�<̒<\��<�(�<LT�<�~�<u��<3χ<���<��<^@�<gd�<�}<kUy<l�u<��q<�"n<�fj<N�f<o�b<3_<*x[<X�W<�T<?NP<;�L<#�H<�1E<�A<N�=<T):<P�6<E�2<�:/<w�+<>(<�k$<&� <�L<#�<�@<y�<�I<��<j<�<��<���;(��;fZ�;v��; \�;���;i��;W�;�!�;���;/�;��;���;g%�;|^�;���;
�;R}�;�;Ş�;�L�;�~;M�s;Ți;��_;�U;��K;8dB;��8;o�/;n�&;�~;�;��;�@;v��:���:J�:�:w��:)�:%��:K"�:��k:}�M:�0:a�:��9*�9��r9U�9�X�7:7����G�O͙�TPϹF.�~�̘6�b�P�17j�x���K���@+��Ͳ���'������̺�"ٺUW������G��_�
�I�����ĺ�s�"���(��x.��[4�&;:�b@���E���K�2�Q�wW��J]��c���h�S�n�t�t��`z����� ��,酻҈�H�����������z��'g��
T���  �  �x=�=x�=#^=��=ܠ=�A=�� =� =O# =q��<���<�<�A�<�~�<$��<���<1�<�j�<m��<��<��<*G�<x{�<���<K��<��<�?�<@m�<I��<���<t��<w�<�8�<�[�<N}�<z��<���<���<3��<_�<�<(�<�6�<B�<�J�<WP�<�R�<R�<N�<�F�<�;�<�,�<w�<6�<��<���<W��<���<�W�<w(�<���<+��<�<g=�<���<���<�[�<��<��<�N�<��<���<��<
��<h-�<M��<t2�<��<=%�<���<q�<�p�<�ֱ<�8�<>��<��<sH�<���<}�<�7�<R��<�Ǣ<�<�K�<���<�ě<���<�4�<?i�<ś�<|̒<a��<�(�<GT�<�~�<w��<7χ<���<��<Z@�<gd�<�}<�Uy<��u<��q<�"n<�fj<��f<s�b<3_<Ux[<s�W<�T<2NP<<�L<�H<�1E<�A<T�=<_):<?�6<?�2<�:/<|�+<?(<�k$<� <�L<#�<�@<d�<�I<��<�i<t<|�<���;B��;[Z�;���;)\�;u��;N��;�V�;�!�;#��;i�;��;���;�%�;N^�;˪�;W
�;s}�;+�;���;�L�;�~;��s;��i;��_;��U;��K;�cB;��8;��/;5�&;�~;��;��;~@;s��:��:yI�:��:��:k(�::�!�:_�k:��M:�0:��:���9�'�96�r9��9H��7p)���G�gƙ�WKϹ]/�N|�+�6�:P��6j� ၺ�����*�������'��o����̺F#ٺrX�l��s��������
���������Ȩ"��(��x.��[4��;:��@�<�E���K��Q�wW��J]�c���h���n�"�t�<`z�<��� ��:酻�ш�A�������[����z���f��$T���  �  �x=�=y�="^=��=۠=�A=�� =� =J# =`��<���<�<�A�<�~�<��<���<1�<�j�<g��<��<��<G�<v{�<���<K��<��<�?�<Um�<E��<���<r��<s�<�8�<�[�<O}�<���<���<���<=��<i�<�<2(�<6�<B�<�J�<TP�<�R�<R�<N�<�F�<�;�<�,�<��<(�<���<���<H��<�<�W�<d(�<���<)��<�<c=�<���<���<�[�<��<(��<�N�<#��<��<��<��<{-�<K��<s2�<��<=%�<���<��<�p�<�ֱ<9�<9��<��<qH�<���<t�<�7�<V��<�Ǣ<�
�<�K�<���<�ě<���<�4�<6i�<Л�<o̒<U��<�(�<GT�<r~�<x��<3χ<���<��<Z@�<|d�<�}<�Uy<��u<��q<�"n<�fj<��f<��b<'3_<@x[<s�W<�T<-NP<e�L< �H<�1E<�A<L�=<^):<�6<?�2<�:/<h�+<(<�k$<� <�L< �<f@<n�<�I<��<�i<~<y�<`��;8��;LZ�;~��;\�;���;���;�V�;�!�;��;V�;��;���;�%�;�^�;窟;4
�;�}�;O�;���;M�;|~;��s;��i;��_;�U;�K;�cB;��8;�/;ځ&;�~;&�;g�;�@;���:���:�H�:W�:1��:=(�:8��:�!�:7�k:��M:(0:?�:���92*�9Y�r98�9�w�7$����G��ƙ��KϹ�,�j|�Q�6�Z}P�7j��߁�`����*��{����'�������̺m#ٺ;X庤��ך�����h�
�v�����j��
�"���(�Ey.�\4��;:��@���E���K�0�Q�wW�uJ]� c�/�h���n���t�`z�f��c ��酻�ш����ä�������z���f��1T���  �  �x=�=v�=%^=��=۠=�A=�� =� =H# =\��<}��<�<�A�<�~�<��<���<1�<�j�<j��<��<��</G�<m{�<���<N��<��<�?�<Im�<Q��<���<���<��<�8�<�[�<I}�<���<���<���<>��<k�<�<&(�<�6�<B�<�J�<IP�<�R�<R�<N�<�F�<�;�<�,�<f�<&�<���<���<J��<���<�W�<Y(�<���<&��<�<p=�<���<«�<�[�<��<��<�N�<'��<��<��<��<�-�<K��<y2�</��<F%�<��<~�<�p�<�ֱ< 9�<9��<��<xH�<���<��<�7�<U��<�Ǣ<�
�<|K�<o��<�ě<���<�4�<+i�<���<j̒<L��<�(�<;T�<�~�<{��<.χ<���<��<]@�<pd�<�}<�Uy<��u<��q<�"n<�fj<o�f<��b<B3_<kx[<��W<�T<ANP<N�L< �H<�1E<�A<F�=<[):<?�6<&�2<�:/<a�+<(<�k$<�� <�L<��<t@<:�<�I<��<�i<~<e�<���;��;[Z�;���;\�;���;o��;W�;�!�;U��;��;?�;���;�%�;�^�;쪟;�
�;�}�;W�;���;�L�;�~;��s;�i;9�_;6�U;Y�K;�cB;A�8;��/;��&;�};�;��;�?;���:���:H�:��:��:(�:���:c"�:��k:��M:�0:{�:��9�(�9
�r9��9�͛7-#����G�Ǚ�[JϹ�)�T{��6��}P��5j�u���Ï���*��=����'��;�����̺�#ٺZX�J��c�����D�
�D��)�����g�"�h�(�my.�I\4��;:��@�I�E�w�K�[�Q��vW��J]�
c���h�i�n���t��_z���9 ���腻�ш�溋�����/����z���f��	T���  �  �x=�=w�=!^=��=ՠ=�A=�� =� =A# =g��<���<��<�A�<�~�<��<x��<1�<�j�<V��<��<��<)G�<i{�<���<B��<��<�?�<Jm�<g��<���<���<|�<�8�<\�<V}�<���<���<���<5��<|�<!�<'(�<�6�<B�<�J�<LP�<�R�<R�<�M�<�F�<v;�<�,�<`�<1�<���<���<T��<���<�W�<T(�<y��<��<�<h=�<���<«�<�[�<��<"��<�N�<;��<��<��<��<�-�<Z��<�2�<��<?%�<��<w�<�p�<�ֱ<9�<E��<��<|H�<���<~�<�7�<D��<�Ǣ<�
�<�K�<c��<�ě<���<�4�<0i�<���<x̒<B��<�(�<)T�<�~�<n��<2χ<���<��<r@�<pd�<�}<�Uy<��u<�q<�"n<�fj<��f<��b<3_<rx[<{�W<�T<hNP<K�L<G�H<�1E<�A<R�=<E):<<�6<�2<n:/<D�+<*(<�k$<�� <�L<��<�@<$�<�I<��<�i<[<K�<���;��;jZ�;W��;0\�;���;n��;rW�;�!�;^��;u�;��;$ �;�%�;�^�;���;�
�;s}�;��;�;�L�;
~;8�s;Кi;T�_;�U;;�K;cB;��8;k�/;.�&;�};c�;��;�?;1��:D��:�I�:Q�:���:�&�:&��:�!�:��k:��M:�0:1�:���9,�9��r9p�9�7�.����G��Ù��FϹ,�a|���6��~P�43j�/������<*�����W'��V���,�̺t$ٺkY庫����������
������r��B�"��(��x.��\4�%<:�y@�R�E���K�7�Q�wW��J]�_c���h�ɾn���t�(`z����~ ���腻�ш�����פ��!����z���f���S���  �  �x=�=y�= ^=��=Ԡ=�A=�� =� =D# =K��<t��<��<�A�<�~�<��<v��<1�<�j�<`��<��<��< G�<n{�<���<G��<��<�?�<Nm�<P��<���<���<��<�8�<	\�<Y}�<���<Ϲ�<���<A��<q�<�<+(�<�6�<B�<�J�<QP�<�R�<R�<N�<�F�<z;�<�,�<]�<�<���<���<>��<���<�W�<R(�<���<*��<!�<\=�<���<���<�[�<��<$��<�N�<-��<��<��<(��<�-�<[��<�2�<,��<[%�<��<��<�p�<�ֱ<9�<?��<��<rH�<���<t�<8�<X��<�Ǣ<�
�<vK�<c��<�ě<���<�4�< i�<���<[̒<I��<�(�<CT�<�~�<i��<3χ<���<��<b@�<ud�<�}<�Uy<��u<�q<
#n<�fj<��f<��b<E3_<�x[<��W<�T<=NP<Y�L<-�H<�1E<߁A<P�=<A):<2�6<=�2<�:/<P�+<�(<�k$<�� <xL<��<a@<�<wI<��<�i<{<�<g��;��;FZ�;h��;!\�;���;}��;W�;�!�;f��;��;*�;3 �;�%�;�^�;/��;�
�;�}�;j�;ƞ�;M�;�~;��s;��i;{�_;��U;��K;�cB;��8;��/;D�&;�};��;��;�?;у�:P��:�G�:+�:H��::(�:��:"!�:��k:l�M:�0:��: ��9G*�9��r9�9��7Q��)�G��Ù�oFϹJ*��x�U�6�/}P��5j����U����*�������'��������̺�"ٺ3X��� ���>����
����k�����ĩ"�˓(��y.�e\4��;:��@�K�E�	�K�-�Q�>wW��J]��c�c�h�T�n���t��_z����" ���腻�ш�������������wz���f��T���  �  Vz=�=�=�`=�=[�=�E=�� =�� =E( =��<	��<[�<�N�<��<���<f�<�A�<}|�<(��<���<{&�<�\�<n��<���<���<+�<M[�<��<_��<��<�<p5�<�[�<���<`��<��<���< ��<�<�0�<�E�<�X�<Zh�<�u�<��<ц�<Ȋ�<���<��<ۂ�<Wy�<�k�< [�<�E�<-�<�<���<E��<B��<�p�<�=�<4�<���<���<�B�<���<��<>S�<���<��<=7�<���<a�<��<iw�<d��<�z�<.��<7k�<�ܶ<�I�<���<\�<�w�<oԮ<@-�<7��<�ө<�!�<.l�<v��<���<79�<�w�<���<��<�#�<�X�<��<���<�<��<B�<�k�<ړ�<º�<k��<��<�(�<RK�<km�<�}<F_y<�u<H�q<* n<�_j<��f<t�b<�_<a[<�W<4�S<�*P<|pL<�H<�E<�MA<ƛ=<��9<J@6<�2<�.<�N+<y�'<$<� <t�<�a<)�<$X<j�<�d<�<��<&<n��;B��;_J�;��;?�;���;�t�;�(�;���;���;���;﫵;>��;�ݩ;��;�]�;G��;-�;ﲍ;�L�;��;	z{;�'q;��f;��\;lS;%gI;8�?;)o6;v,-;1$; ;�:;��	;f� ; �:�\�:���:�ɿ:ׯ:��:���:�L�:@bd:)�F:4):��:�@�9N�9��Y9���8�y�)B�%[]��I���nٹ���1!�(!;��T�Khn� 䃺�������z���ݵ�".º�pκۢں��溯�����$t�Em��b�NQ��<��##�H)���.���4���:��q@��EF��L�`�Q���W���]�Rc�>i���n�p�t��~z��$��?
��$���2ֈ�����㋑��t���]���H���  �  Uz=�=�=�`=�=U�=�E=�� =�� =?( =��<��<X�<�N�<݌�<���<^�<�A�<t|�<"��<���<z&�<�\�<e��<���<���<!+�<][�<��<[��<��<!�<w5�<�[�<���<\��<��<���<��<�<�0�<�E�<�X�<ph�<�u�<��<Ȇ�<���<���<���<��<My�<�k�<�Z�<�E�<
-�<�<���<:��<C��<�p�<�=�<D�<���<���<�B�<���<��<US�<���<ߚ�<>7�<���<a�<��<qw�<^��<�z�<4��<>k�<�ܶ<�I�<���<V�<�w�<�Ԯ<B-�<=��<�ө<�!�<-l�<���<���<,9�<�w�<���<��<�#�<�X�<	��<���<�<��<B�<�k�<ٓ�<���<k��<�<�(�<fK�<em�<w}<:_y<�u<X�q<! n<�_j<x�f<��b<�_<a[<�W<#�S<{*P<vpL<,�H<�E<�MA<ɛ=<��9<F@6<%�2<A�.<�N+<p�'<$<� <r�<�a<=�<X<l�<�d<�<ǉ<&<g��; ��;xJ�;��;Q?�;���;�t�;�(�;a��;���;���;���;b��;�ݩ;�;�]�;���;'-�;鲍;�L�;��;�z{;�'q;�f;��\;/S;gI;��?;�o6;-,-;4$;�;6;;C�	;
� ;� �:�[�:��:ɿ:�ׯ:��:���:IL�:�`d:b�F:>):w�:�A�9-L�9�Y9	��8��v�>�BW]��J��Mnٹ���0!�T;��T�zhn�䃺�~��M��xz��]ݵ��.ºqκ�ںf�����b���t��m�Fb��Q��<��##��)���.��4���:�zq@��EF�)L�]�Q�:�W���]�uQc�gi���n���t�i~z��$��R
�����^ֈ�Ѽ�����͋��st���]���H���  �  Sz=�=�=�`=�=X�=�E=�� =�� =>( =��<��<^�<O�<ߌ�<��<]�<�A�<|�< ��<���<p&�<	]�<g��<���<���<+�<T[�<��<h��<��<�<a5�<�[�<���<V��<��<���<��<�<�0�<�E�<�X�<ph�<vu�<��<ǆ�<Ί�<���<��<��<Ny�<l�<�Z�<F�<-�<�<���<7��<[��<�p�<�=�<>�<���<È�<�B�<���<��<RS�<���<��<A7�<���<a�<��<hw�<X��<�z�<(��<&k�<�ܶ<�I�<���<U�<�w�<}Ԯ<:-�<F��<�ө<�!�<$l�<���<���<39�<�w�<���<�<�#�<�X�<��<���<*�<��<B�<�k�<䓋<���<n��<
�<�(�<fK�<am�<�}<._y<
�u<E�q<�n<�_j<n�f<��b<�_<�`[<�W<�S<�*P<ppL<&�H<�E<�MA<ԛ=<��9<^@6<�2<O�.<�N+<��'<$<� <��<�a<j�<X<��<�d<�<щ<
&<���;+��;�J�;��;6?�;���;�t�;�(�;2��;���;d��;���;]��;�ݩ;��;t]�;j��;�,�;貍;�L�;���;�z{;$'q;j�f;��\;�S;,gI;`�?;�o6;1,-;�$;�;�;;{�	;)� ;%�:�[�:���:@ɿ:�ׯ:��:w��:7M�:�`d:ЉF:�):�:�?�9�L�9�Y9w��8�w��S�7[]�TL���oٹK��3!��;���T��fn��䃺�������z���ܵ��.ºpκy�ںW����������s��m��a��Q��<�H##��)�l�.��4�̚:��q@��EF��L�G�Q��W�/�]�vQc��i���n�ҳt��~z��$���
�����rֈ�˼��_��� ����t��&^���H���  �  Rz=�=�=�`=�=W�=�E=�� =�� =D( =��<��<a�<O�<��<��<f�<�A�<�|�<*��<���<|&�<]�<c��<���<���<+�<Q[�<��<S��<��<�<g5�<�[�<���<W��<	��<���<��<�<�0�<�E�<�X�<dh�<~u�<��<���<ʊ�<���<���<��<Ry�<l�<�Z�<F�<-�<�<���<@��<R��<�p�<�=�<C�<���<���<�B�<���<��<IS�<���<���<17�<���<a�<��<`w�<V��<�z�<)��<-k�<�ܶ<�I�<���<S�<�w�<{Ԯ<=-�<=��<�ө<�!�<-l�<���<���<69�<�w�<���<��<�#�<�X�<��<���<(�<��<B�<�k�<���<���<c��<�<�(�<[K�<`m�<v}<_y<��u<G�q< n<�_j<u�f<c�b<�_<�`[<�W<�S<q*P<lpL<�H<�E<�MA<��=<��9<Z@6</�2<O�.<�N+<��'<$<� <��<�a<Z�<&X<~�<�d<�<ω<"&<���;��;wJ�;��;C?�;���;�t�;�(�;3��;���;|��;֫�;��;�ݩ;��;�]�;c��;�,�;���;�L�;���;dz{;h'q;#�f;\�\;zS;(gI;��?;�o6;T,-;�$;�;�;;φ	;�� ;��:S\�:	��:wɿ:=د:��:���:M�:�_d:^�F:�):*�:�?�9�L�9Y�Y9��8�-x�qI��^]��L���rٹ��2!�� ;���T��in��䃺�������z��Rݵ�+/º&pκڢںU��=������s�Ym��a�KQ�r<�G##�c)�u�.���4�ؚ:�Xq@��EF��L���Q�J�W���]��Qc��i���n��t��~z��$��q
��D���cֈ����<���󋑻�t��<^���H���  �  Tz=�=�=�`=�=[�=�E=�� =�� =I( =!��<"��<w�<O�<���<��<��<�A�<�|�<2��<���<�&�<]�<q��<���<~��<+�<N[�<��<H��<��<�<Z5�<�[�<���<Q��<���<���<���<�<�0�<�E�<�X�<]h�<}u�<��<φ�<Њ�<���<��<��<by�<l�<[�<F�<-�<�<���<^��<U��<�p�<�=�<N�<���<È�<�B�<���<��<AS�<���<ٚ�<)7�<���<�`�<��<Mw�<O��<�z�<��<!k�<�ܶ<�I�<���<Q�<�w�<tԮ<9-�<;��<�ө<�!�<7l�<���<���<C9�<�w�<ó�<��<�#�<�X�<&��<���<(�<��<B�<�k�<ᓋ<ƺ�<p��<��<�(�<VK�<em�<a}<_y<�u<�q<�n<�_j<o�f<8�b<�_<�`[<٢W<�S<Y*P<rpL<�H<�E<�MA<ϛ=<��9<U@6<G�2<D�.<O+<��'<C$<?� <��<b<`�<bX<��<�d<+�<щ<8&<���;V��;J�;���;6?�;���;�t�;p(�;Y��;{��;J��;���;⺯;�ݩ;��;x]�;뺘;�,�;���;�L�;���;/z{;g'q;��f;��\;�S;ngI;�?;�o6;�,-;�$;�;�;;��	;�� ;!�:?^�:A��:ʿ:�د:��:V��:FM�:�ad:��F:x):=�:�>�9K�9��Y9���8�{�mS�h]�N���tٹ�*4!��";���T�kn��䃺���)���z��gݵ�9.º[pκ?�ں���������\s�^l��a��P�K<��"#��)�{�.�[�4��:��p@��EF��L�:�Q���W��]��Qc�ni�S�n��t�z�'%���
������nֈ�e���g���J����t��+^���H���  �  Mz=�=�=�`=�=[�=�E=�� =�� =R( =3��<��<u�<O�<��<$��<u�<�A�<�|�<?��<���<�&�<]�<o��<���<���<+�<@[�<��<N��<���<��<Q5�<�[�<���<<��<���<���<���<��<�0�<�E�<vX�<bh�<yu�<��<Ɇ�<ӊ�<���<��<���<sy�<l�<[�<F�<.-�<&�<���<O��<^��<q�<�=�<N�<���<ǈ�<�B�<���<��<GS�<��<Ӛ�<"7�<���<�`�<��<Hw�<;��<zz�<��<k�<�ܶ<�I�<���<I�<�w�<wԮ<9-�<<��<�ө<�!�<2l�<���<���<P9�<�w�<���<�<$�<�X�<'��<���<7�<�<&B�<�k�<�<Ⱥ�<n��<�<�(�<SK�<Tm�<b}<�^y<؟u<�q<�n<�_j<?�f<6�b<�_<�`[<ȢW<��S<a*P<UpL<��H<�E<�MA<ϛ=<��9<q@6<7�2<`�.<4O+<��'<<$<;� <��<.b<��<GX<��<�d<F�<�<1&<Β�;S��;�J�;��;:?�;]��;�t�;�(�;���;`��;+��;���;ں�;\ݩ;{�;f]�;�;�,�;���;�L�;���;[z{;J'q;/�f;��\;�S;�gI;��?;Sp6;c--; $;�;X<;o�	;@� ;T�:_]�:���:o˿:$ٯ:��:i��:�M�:"ad:��F:):�:
;�9�I�9��Y9���8� |�&\��i]�S���vٹ��>5!�K#;���T�ejn�,僺̀������z��Dݵ�V.º�oκz�ں_��@�����Ns��l�$a�nP��;��"#��)���.���4�|�:�2q@�GEF��L�J�Q�H�W��]�Rc��i�K�n���t�cz�'%���
�������ֈ�h���q���W����t���^���H���  �  Ez=�=�=�`=�=\�=�E=�� =�� =M( ==��<0��<��<'O�< ��<8��<��<B�<�|�<=��<���<�&�<]�<j��<���<z��<+�<G[�<���<F��<���<��<C5�<�[�<y��<*��<���<y��<���<��<�0�<�E�<oX�<fh�<mu�<��<ņ�<ڊ�<���<��<	��<fy�<,l�<[�<4F�<6-�<)�<���<]��<q��<�p�<�=�<Z�<���<Ј�<�B�<���<���<HS�<|��<Ϛ�<7�<t��<�`�<y�<Ew�<(��<iz�<
��<k�<�ܶ<�I�<���<;�<�w�<vԮ<.-�<<��<�ө<�!�<3l�<���<���<O9�<�w�<���<%�<$�<�X�<:��<���<F�<�<6B�<�k�<���<̺�<l��<��<�(�<YK�<Fm�<_}<�^y<Ɵu<��q<�n<_j<�f<%�b<�_<�`[<��W<��S<[*P<6pL<�H<�E<�MA<˛=<��9<~@6<9�2<��.<"O+<˰'<b$<^� <��< b<��<iX<��<e<C�<�<5&<��;A��;�J�;��;5?�;}��;Dt�;s(�;���;S��;���;o��;���;ݩ;t�;]�;޺�;�,�;^��;�L�;���;�z{;�&q;#�f;��\;S;�gI;9�?;�p6;--;�$;;=;��	;[� ;��:=^�:��:�ʿ:�ٯ:� �:���:/N�:D`d:d�F:a):Z�:V:�9I�94�Y9���8��|�Rr⸸j]�UW���zٹ��7!��#;���T��kn��僺r�������{��8ݵ��.ºoκ`�ںb��������r�dl�z`��P�H;�	"#�9)���.�&�4���:�#q@�)EF��L�\�Q�c�W�Z�]��Qc�di�Y�n���t��z�[%���
������3׈�������������u���^���H���  �  Dz=�=�=�`=�=_�=�E=�� =�� =T( =C��<?��<��<1O�<��<=��<��<B�<�|�<G��<���<�&�<]�<s��<���<}��<+�<D[�<���<8��<���<��<05�<�[�<i��<-��<���<i��<���<��<�0�<�E�<mX�<]h�<uu�<��<ц�<ڊ�<���<��<��<uy�<1l�<,[�<8F�<F-�<9�<���<q��<u��<q�<>�<_�<���<Έ�<�B�<���<��<>S�<x��<���<7�<x��<�`�<k�</w�<&��<]z�<���<�j�<ܶ<�I�<���<2�<�w�<nԮ<0-�<>��<�ө<�!�<<l�<���<���<X9�<�w�<׳�<(�<$�<�X�<F��<���<I�<�<=B�<�k�<쓋<Ϻ�<t��<��<�(�<RK�<Em�<=}<�^y<��u<��q<�n<Y_j<�f<�b<p_<�`[<��W<��S<5*P<3pL<��H<�E<�MA<؛=<��9<p@6<[�2<��.<<O+<ְ'<�$<� <��<Pb<��<�X<��<e<[�<�<R&<ߒ�;m��;�J�;��;(?�;w��;8t�;<(�;���;��;���;��;o��;)ݩ;�;�\�;���;�,�;M��;dL�;���;=z{;0'q; �f;��\;S;�gI;��?;�p6;--;�$;�;+=;:�	;�� ;��:�_�:[��:�˿:Mگ:� �:���:N�:bd:��F:U):1�:�9�9xE�9�Y9���8Z�~�y�ku]��W���}ٹ3�]9!�P&;�+�T��ln�u惺����R��V{��
ݵ�.ºYoκ��ںK��o��~���br��k�[`��O��:��!#��)�l�.���4�Ǚ:��p@�cEF�wL��Q�c�W�A�]�Rc�hi���n�ִt��z��%��<���׈�ͽ������ތ��4u���^��8I���  �  Hz=�=�=�`=�=`�=�E=�� =�� =`( =K��<D��<��<2O�</��<>��<��<B�<�|�<X��<���<�&�<]�<z��<���<���<+�<6[�< ��<+��<���<��<85�<�[�<Z��< ��<���<z��<���<��<�0�<�E�<oX�<Rh�<wu�<��<І�<Ԋ�<���<��<��<�y�<4l�<3[�<=F�<Q-�<J�<���<z��<v��<q�<	>�<c�<���<ƈ�<�B�<���<��<6S�<w��<���<7�<i��<�`�<y�<w�<��<Mz�<���<�j�<rܶ<�I�<}��<6�<�w�<lԮ<5-�<5��<�ө<�!�<Ml�<���<��<f9�<�w�<۳�<)�<+$�<�X�<J��<û�<R�</�<7B�<�k�<���<к�<n��<��<�(�<DK�<Jm�<!}<�^y<��u<��q<�n<._j<�f<��b<x_<�`[<��W<��S<*P<BpL<�H<�E<�MA<̛=<��9<�@6<w�2<��.<oO+<�'<�$<�� <��<�b<��<�X<��<,e<~�<�<u&<��;���;�J�;��;#?�;A��;Yt�;(�;���;���;Ѯ�;��;8��;�ܩ;��;]�;}��;a,�;*��;?L�;���;�y{;H'q;�f;��\;�S;.hI;��?;�p6;?.-;$;�;X=;��	;n� ;�:(`�:���:$Ϳ:�گ:"!�:���:�M�:Rbd:ǇF:�):S�:�9�9�D�9�Y9F��8S��ep⸇]�:[���ٹZ�8!��';�a�T�\nn�惺Q���n���z���ݵ��-º�oκ��ں*�溠�����kr��k�O`�NO��:��!#��)�$�.�տ4���:�2p@�EF�nL�I�Q�p�W�5�]��Rc�Ci�N�n�F�t�S�z��%����[�>׈����礎�Ќ��}u���^��oI���  �  Cz=�=�=�`=�=c�=�E=�� =Ň =]( =V��<W��<��<GO�<2��<U��<��<+B�<�|�<Y��<��<�&�<]�<y��<���<r��<+�<3[�<��<+��<���<��<5�<�[�<U��<��<���<Z��<���<��<�0�<�E�<fX�<Th�<hu�<��<ӆ�<ۊ�<���<��<��<�y�<Il�<?[�<NF�<W-�<O�<��<���<���<q�<>�<g�<��<͈�<�B�<���<���<4S�<l��<���<�6�<Y��<�`�<X�<w�<��<Gz�<���<�j�<uܶ<�I�<x��<)�<�w�<cԮ<$-�<;��<�ө<�!�<Ll�<���<��<j9�<x�<糝<?�<0$�<�X�<W��<ӻ�<^�<&�<BB�<�k�<���<պ�<u��<��<�(�<IK�<Am�<&}<�^y<��u<��q<�n<*_j<�f<��b<I_<e`[<y�W<��S<#*P<+pL<�H<�E<~MA<ڛ=<��9<�@6<p�2<��.<bO+<��'<�$<�� <&�<�b<��<�X<�<<e<��<,�<q&<��;���;�J�;ܼ�;?�;;��;,t�;(�;v��;���;n��;Ӫ�;%��;�ܩ;��;�\�;N��;*,�;��;.L�;���;�y{;�&q;#�f;�\;S;jhI;��?;7q6;.-;�$;2;�=;ˈ	;�� ;'�:�`�:.��:�̿:ۯ:w!�:��:!N�:ybd:Q�F:�
):�:$7�9=B�9g�Y9���8�Y�����4�]��]��U�ٹ
��;!�\';�T�T��nn��惺��������{��ݵ��-º!oκ��ں��溄��J���vq�)k��_�&O�N:� !#�)���.��4���:�Pp@��DF�IL��Q���W���]�_Rc��i�;�n���t���z��%����a񅻂׈�&���E�������u�� _��[I���  �  <z=�=�=�`=�=^�=�E=�� =͇ =_( =c��<S��<��<YO�<0��<a��<��<+B�<�|�<b��<
��<�&�<$]�<p��<���<}��<+�<7[�<��<,��<���<��<5�<�[�<O��<��<���<Q��<���<��<�0�<�E�<]X�<Vh�<mu�<��<Ά�<݊�<���< ��<.��<�y�<Ul�<6[�<NF�<a-�<S�<��<y��<���<q�<">�<i�<��<ӈ�<�B�<���<���<5S�<f��<���<�6�<T��<�`�<P�<w�<���<=z�<���<�j�<wܶ<�I�<x��< �<�w�<gԮ<,-�<C��<�ө<�!�<Jl�<���<��<k9�<x�<ڳ�<I�<0$�<�X�<P��<ͻ�<m�<'�<VB�<�k�<��<Ϻ�<u��<�<�(�<JK�<3m�<'}<�^y<��u<��q<yn<8_j<ɞf<��b<?_<h`[<}�W<��S<#*P<pL<�H<�E<�MA<ߛ=<��9<�@6<u�2<��.<lO+<�'<�$<�� <J�<�b<�<�X<�<He<��<>�<q&</��;g��;�J�;��;?�;I��;t�;(�;Q��;���;V��;ڪ�;��;�ܩ;��;|\�;q��;,�;���;'L�;]��;z{;'q;j�f;��\;7S;\hI;��?;�q6;.-;$;�;�=;�	;�� ;u�:)`�:���:�̿:"ܯ:�!�:���:�N�:�ad:��F:�):\�:�5�91A�9'�Y9���8��4���}]��`����ٹ���<!��&;��T��nn�i烺�������k{���ܵ�N.ºinκĠںn�����.���kq��k�R_�'O��9�W!#�=)�P�.��4���:�>p@��DF�sL��Q�:�W�w�]�TRc��i�6�n��t���z��%�����F񅻷׈����X�������u��2_��[I���  �  @z=�=޾=�`=�=e�=�E=�� =Ǉ =e( =e��<b��<��<WO�<5��<b��<��<3B�<�|�<g��< ��<�&�<#]�<~��<���<|��<+�<.[�<��<(��<���<��<5�<�[�<D��<��<���<T��<���<��<�0�<�E�<eX�<Fh�<mu�<��<؆�<��<���< ��<#��<�y�<Yl�<M[�<XF�<g-�<Y�<��<���<���<#q�<>�<g�<
��<ֈ�<�B�<���<���<&S�<j��<���<�6�<Q��<�`�<Q�<w�<���<4z�<���<�j�<_ܶ<�I�<t��<&�<�w�<ZԮ<--�<:��<�ө<�!�<Pl�<���<��<w9�<x�<<N�<5$�<�X�<a��<໔<p�<3�<IB�<�k�<	��<ٺ�<y��<��<�(�<<K�<>m�<}<�^y<q�u<��q<wn<_j<ƞf<��b<6_<T`[<a�W<��S<*P<!pL<ѷH<�E<�MA<ݛ=<��9<�@6<z�2<��.<�O+<�'<�$<�� <G�<�b<�<�X<.�<Ze<��<+�<|&<.��;���;�J�;��;�>�;)��;#t�;(�;Z��;���;a��;���;幯;�ܩ;��;�\�;+��;,�;���;.L�;~��;�y{;'q;�f;@�\;eS;�hI;��?;�q6;w.-;5$;�;5>;N�	;�� ;��:�a�:���:�Ϳ:�ۯ:z!�:n��:�N�:3cd:K�F:�):t�:�6�9{B�9w�Y9���8�7�����1�]�la��͆ٹw�A<!��);���T�8on�烺灐�e��]{��"ݵ�i-ºonκi�ں��溡��i���7q��j�&_�O��9�� #��)�2�.���4�`�:�(p@��DF�(L���Q�r�W���]��Rc��i�]�n�εt���z�	&������񅻼׈�f���j���<����u��%_��vI���  �  ?z=�=�=�`=�=c�=�E=�� =ʇ =i( =T��<]��<��<NO�<>��<]��<��<*B�<�|�<k��<��<�&�<]�<���<���<{��<
+�</[�<��<��<���<��<#5�<�[�<J��<��<���<^��<���<��<�0�<�E�<fX�<Jh�<zu�<��<Ն�<͊�<���<'��<#��<�y�<Cl�<G[�<QF�<i-�<_�<��<���<���<&q�<>�<n�<��<���<�B�<���<
��<-S�<k��<���<�6�<]��<�`�<\�<�v�<��<>z�<���<�j�<_ܶ<�I�<a��<�<�w�<bԮ<1-�<0��<�ө<�!�<Sl�<���<��<s9�< x�<�<I�<:$�<�X�<`��<ڻ�<Z�<=�<NB�<�k�<���<κ�<w��<��<�(�<<K�<>m�<�}<�^y<��u<��q<�n<�^j<�f<��b<?_<V`[<m�W<��S<�)P<pL<ַH<�E<�MA<֛=<��9<|@6<��2<��.<�O+<��'<�$<�� <5�<�b<�<�X<�<Je<��<:�<�&<ܒ�;���;�J�;��;?�;-��;t�;�'�;~��;���;���;���; ��;�ܩ;_�;�\�;!��;4,�;���;�K�;���;�y{;k'q;��f;,�\;�S;ShI;�?;�q6;�.-;�$;{;�=;`�	;� ;��:La�:���:�Ϳ:�ۯ:�!�: ��:[M�:	cd:!�F:r):o�:C7�9�=�9!�Y9���8�S�����w�]�0^��y�ٹ���:!��);���T��qn��烺́�����{���ݵ�G-º�oκ4�ںL��w������q��j�M_��N�:�� #��)���.�`�4�9�:��o@�EF�|L� �Q���W�E�]��Rc��i��n���t���z�&�������}׈�n���W���7����u���^���I���  �  @z=�=޾=�`=�=e�=�E=�� =Ǉ =e( =e��<b��<��<WO�<5��<b��<��<3B�<�|�<g��< ��<�&�<#]�<~��<���<|��<+�<.[�<��<(��<���<��<5�<�[�<D��<��<���<T��<���<��<�0�<�E�<eX�<Fh�<mu�<��<؆�<��<���< ��<#��<�y�<Yl�<M[�<XF�<g-�<Y�<��<���<���<#q�<>�<g�<
��<ֈ�<�B�<���<���<&S�<j��<���<�6�<Q��<�`�<Q�<w�<���<4z�<���<�j�<_ܶ<�I�<t��<&�<�w�<ZԮ<--�<:��<�ө<�!�<Pl�<���<��<w9�<x�<<N�<5$�<�X�<a��<໔<p�<3�<IB�<�k�<	��<ٺ�<y��<��<�(�<<K�<>m�<}<�^y<q�u<��q<wn<_j<ƞf<��b<6_<T`[<a�W<��S<*P<!pL<ѷH<�E<�MA<ݛ=<��9<�@6<z�2<��.<�O+<�'<�$<�� <G�<�b<�<�X<.�<Ze<��<+�<|&<.��;���;�J�;��;�>�;)��;#t�;(�;Z��;���;a��;���;幯;�ܩ;��;�\�;+��;,�;���;.L�;~��;�y{;'q;�f;@�\;eS;�hI;��?;�q6;w.-;5$;�;5>;N�	;�� ;��:�a�:���:�Ϳ:�ۯ:z!�:n��:�N�:3cd:K�F:�):t�:�6�9{B�9w�Y9���8�7�����1�]�la��͆ٹw�A<!��);���T�8on�烺灐�e��]{��"ݵ�i-ºonκi�ں��溡��i���7q��j�&_�O��9�� #��)�2�.���4�`�:�(p@��DF�(L���Q�r�W���]��Rc��i�]�n�εt���z�	&������񅻼׈�f���j���<����u��%_��vI���  �  <z=�=�=�`=�=^�=�E=�� =͇ =_( =c��<S��<��<YO�<0��<a��<��<+B�<�|�<b��<
��<�&�<$]�<p��<���<}��<+�<7[�<��<,��<���<��<5�<�[�<O��<��<���<Q��<���<��<�0�<�E�<]X�<Vh�<mu�<��<Ά�<݊�<���< ��<.��<�y�<Ul�<6[�<NF�<a-�<S�<��<y��<���<q�<">�<i�<��<ӈ�<�B�<���<���<5S�<f��<���<�6�<T��<�`�<P�<w�<���<=z�<���<�j�<wܶ<�I�<x��< �<�w�<gԮ<,-�<C��<�ө<�!�<Jl�<���<��<k9�<x�<ڳ�<I�<0$�<�X�<P��<ͻ�<m�<'�<VB�<�k�<��<Ϻ�<u��<�<�(�<JK�<3m�<'}<�^y<��u<��q<yn<8_j<ɞf<��b<?_<h`[<}�W<��S<#*P<pL<�H<�E<�MA<ߛ=<��9<�@6<u�2<��.<lO+<�'<�$<�� <J�<�b<�<�X<�<He<��<>�<q&</��;g��;�J�;��;?�;I��;t�;(�;P��;���;V��;ڪ�;��;�ܩ;��;|\�;q��;,�;���;'L�;]��;z{;'q;j�f;��\;7S;\hI;��?;�q6;.-;$;�;�=;�	;�� ;u�:)`�:���:�̿:"ܯ:�!�:���:�N�:�ad:��F:�):\�:�5�91A�9'�Y9���8��4���}]��`����ٹ���<!��&;��T��nn�i烺�������k{���ܵ�N.ºinκĠںn�����.���kq��k�R_�'O��9�W!#�=)�P�.��4���:�>p@��DF�sL��Q�:�W�w�]�TRc��i�6�n��t���z��%�����F񅻷׈����X�������u��2_��[I���  �  Cz=�=�=�`=�=c�=�E=�� =Ň =]( =V��<W��<��<GO�<2��<U��<��<+B�<�|�<Y��<��<�&�<]�<y��<���<r��<+�<3[�<��<+��<���<��<5�<�[�<U��<��<���<Z��<���<��<�0�<�E�<fX�<Th�<hu�<��<ӆ�<ۊ�<���<��<��<�y�<Il�<?[�<NF�<W-�<O�<��<���<���<q�<>�<g�<��<͈�<�B�<���<���<4S�<l��<���<�6�<Y��<�`�<X�<w�<��<Gz�<���<�j�<uܶ<�I�<x��<)�<�w�<cԮ<$-�<;��<�ө<�!�<Ll�<���<��<j9�<x�<糝<?�<0$�<�X�<W��<ӻ�<^�<&�<BB�<�k�<���<պ�<u��<��<�(�<IK�<Am�<&}<�^y<��u<��q<�n<*_j<�f<��b<I_<e`[<y�W<��S<#*P<+pL<�H<�E<~MA<ڛ=<��9<�@6<p�2<��.<bO+<��'<�$<�� <&�<�b<��<�X<�<<e<��<,�<q&<��;���;�J�;ܼ�;?�;;��;,t�;(�;v��;���;n��;Ӫ�;%��;�ܩ;��;�\�;N��;*,�;��;.L�;���;�y{;�&q;#�f;�\;S;jhI;��?;7q6;.-;�$;2;�=;ˈ	;�� ;'�:�`�:.��:�̿:ۯ:w!�:��:!N�:ybd:Q�F:�
):�:$7�9=B�9g�Y9���8�Y�����4�]��]��U�ٹ
��;!�\';�T�T��nn��惺��������{��ݵ��-º!oκ��ں��溄��J���vq�)k��_�&O�N:� !#�)���.��4���:�Pp@��DF�IL��Q���W���]�_Rc��i�;�n���t���z��%����a񅻂׈�&���E�������u�� _��[I���  �  Hz=�=�=�`=�=`�=�E=�� =�� =`( =K��<D��<��<2O�</��<>��<��<B�<�|�<X��<���<�&�<]�<z��<���<���<+�<6[�< ��<+��<���<��<85�<�[�<Z��< ��<���<z��<���<��<�0�<�E�<oX�<Rh�<wu�<��<І�<Ԋ�<���<��<��<�y�<4l�<3[�<=F�<Q-�<J�<���<z��<v��<q�<	>�<c�<���<ƈ�<�B�<���<��<6S�<w��<���<7�<i��<�`�<y�<w�<��<Mz�<���<�j�<rܶ<�I�<}��<6�<�w�<lԮ<5-�<5��<�ө<�!�<Ml�<���<��<f9�<�w�<۳�<)�<+$�<�X�<J��<û�<R�</�<7B�<�k�<���<к�<n��<��<�(�<DK�<Jm�<!}<�^y<��u<��q<�n<._j<�f<��b<x_<�`[<��W<��S<*P<BpL<�H<�E<�MA<̛=<��9<�@6<w�2<��.<oO+<�'<�$<�� <��<�b<��<�X<��<,e<~�<�<u&<��;���;�J�;��;#?�;A��;Yt�;(�;���;���;Ѯ�;��;8��;�ܩ;��;]�;}��;a,�;*��;?L�;���;�y{;H'q;�f;��\;�S;.hI;��?;�p6;?.-;$;�;X=;��	;n� ;�:(`�:���:$Ϳ:�گ:"!�:���:�M�:Rbd:ǇF:�):S�:�9�9�D�9�Y9F��8S��ep⸇]�:[���ٹZ�8!��';�a�T�\nn�惺Q���n���z���ݵ��-º�oκ��ں*�溠�����kr��k�O`�NO��:��!#��)�$�.�տ4���:�2p@�EF�nL�I�Q�p�W�5�]��Rc�Ci�N�n�F�t�S�z��%����[�>׈����礎�Ќ��}u���^��oI���  �  Dz=�=�=�`=�=_�=�E=�� =�� =T( =C��<?��<��<1O�<��<=��<��<B�<�|�<G��<���<�&�<]�<s��<���<}��<+�<D[�<���<8��<���<��<05�<�[�<i��<-��<���<i��<���<��<�0�<�E�<mX�<]h�<uu�<��<ц�<ڊ�<���<��<��<uy�<1l�<,[�<8F�<F-�<9�<���<q��<u��<q�<>�<_�<���<Έ�<�B�<���<��<>S�<x��<���<7�<x��<�`�<k�</w�<&��<]z�<���<�j�<ܶ<�I�<���<2�<�w�<nԮ<0-�<>��<�ө<�!�<<l�<���<���<X9�<�w�<׳�<(�<$�<�X�<F��<���<I�<�<=B�<�k�<쓋<Ϻ�<t��<��<�(�<RK�<Em�<=}<�^y<��u<��q<�n<Y_j<�f<�b<p_<�`[<��W<��S<5*P<3pL<��H<�E<�MA<؛=<��9<p@6<[�2<��.<<O+<ְ'<�$<� <��<Pb<��<�X<��<e<[�<�<R&<ߒ�;m��;�J�;��;(?�;w��;8t�;<(�;���;��;���;��;o��;)ݩ;�;�\�;���;�,�;M��;dL�;���;=z{;0'q; �f;��\;S;�gI;��?;�p6;--;�$;�;+=;:�	;�� ;��:�_�:[��:�˿:Mگ:� �:���:N�:bd:��F:U):1�:�9�9xE�9�Y9���8Z�~�y�ku]��W���}ٹ3�]9!�P&;�+�T��ln�u惺����R��V{��
ݵ�.ºYoκ��ںK��o��~���br��k�[`��O��:��!#��)�l�.���4�Ǚ:��p@�cEF�wL��Q�c�W�A�]�Rc�hi���n�ִt��z��%��<���׈�ͽ������ތ��4u���^��8I���  �  Ez=�=�=�`=�=\�=�E=�� =�� =M( ==��<0��<��<'O�< ��<8��<��<B�<�|�<=��<���<�&�<]�<j��<���<z��<+�<G[�<���<F��<���<��<C5�<�[�<y��<*��<���<y��<���<��<�0�<�E�<oX�<fh�<mu�<��<ņ�<ڊ�<���<��<	��<fy�<,l�<[�<4F�<6-�<)�<���<]��<q��<�p�<�=�<Z�<���<Ј�<�B�<���<���<HS�<|��<Ϛ�<7�<t��<�`�<y�<Ew�<(��<iz�<
��<k�<�ܶ<�I�<���<;�<�w�<vԮ<.-�<<��<�ө<�!�<3l�<���<���<O9�<�w�<���<%�<$�<�X�<:��<���<F�<�<6B�<�k�<���<̺�<l��<��<�(�<YK�<Fm�<_}<�^y<Ɵu<��q<�n<_j<�f<%�b<�_<�`[<��W<��S<[*P<6pL<�H<�E<�MA<˛=<��9<~@6<9�2<��.<"O+<˰'<b$<^� <��< b<��<iX<��<e<C�<�<5&<��;A��;�J�;��;5?�;}��;Dt�;s(�;���;S��;���;o��;���;ݩ;t�;]�;޺�;�,�;^��;�L�;���;�z{;�&q;#�f;��\;S;�gI;9�?;�p6;--;�$;;=;��	;[� ;��:=^�:��:�ʿ:�ٯ:� �:���:/N�:D`d:d�F:a):Z�:V:�9I�94�Y9���8��|�Rr⸸j]�UW���zٹ��7!��#;���T��kn��僺r�������{��8ݵ��.ºoκ`�ںb��������r�dl�z`��P�H;�	"#�9)���.�&�4���:�#q@�)EF��L�\�Q�c�W�Z�]��Qc�di�Y�n���t��z�[%���
������3׈�������������u���^���H���  �  Mz=�=�=�`=�=[�=�E=�� =�� =R( =3��<��<u�<O�<��<$��<u�<�A�<�|�<?��<���<�&�<]�<o��<���<���<+�<@[�<��<N��<���<��<Q5�<�[�<���<<��<���<���<���<��<�0�<�E�<vX�<bh�<yu�<��<Ɇ�<ӊ�<���<��<���<sy�<l�<[�<F�<.-�<&�<���<O��<^��<q�<�=�<N�<���<ǈ�<�B�<���<��<GS�<��<Ӛ�<"7�<���<�`�<��<Hw�<;��<zz�<��<k�<�ܶ<�I�<���<I�<�w�<wԮ<9-�<<��<�ө<�!�<2l�<���<���<P9�<�w�<���<�<$�<�X�<'��<���<7�<�<&B�<�k�<�<Ⱥ�<n��<�<�(�<SK�<Tm�<b}<�^y<؟u<�q<�n<�_j<?�f<6�b<�_<�`[<ȢW<��S<a*P<UpL<��H<�E<�MA<ϛ=<��9<q@6<7�2<`�.<4O+<��'<<$<;� <��<.b<��<GX<��<�d<F�<�<1&<Β�;S��;�J�;��;:?�;]��;�t�;�(�;���;`��;+��;���;ں�;\ݩ;{�;f]�;�;�,�;���;�L�;���;[z{;J'q;/�f;��\;�S;�gI;��?;Sp6;c--; $;�;X<;o�	;@� ;T�:_]�:���:o˿:$ٯ:��:i��:�M�:"ad:��F:):�:
;�9�I�9��Y9���8� |�&\��i]�S���vٹ��>5!�K#;���T�ejn�,僺̀������z��Dݵ�V.º�oκz�ں_��@�����Ns��l�$a�nP��;��"#��)���.���4�|�:�2q@�GEF��L�J�Q�H�W��]�Rc��i�K�n���t�cz�'%���
�������ֈ�h���q���W����t���^���H���  �  Tz=�=�=�`=�=[�=�E=�� =�� =I( =!��<"��<w�<O�<���<��<��<�A�<�|�<2��<���<�&�<]�<q��<���<~��<+�<N[�<��<H��<��<�<Z5�<�[�<���<Q��<���<���<���<�<�0�<�E�<�X�<]h�<}u�<��<φ�<Њ�<���<��<��<by�<l�<[�<F�<-�<�<���<^��<U��<�p�<�=�<N�<���<È�<�B�<���<��<AS�<���<ٚ�<)7�<���<�`�<��<Mw�<O��<�z�<��<!k�<�ܶ<�I�<���<Q�<�w�<tԮ<9-�<;��<�ө<�!�<7l�<���<���<C9�<�w�<ó�<��<�#�<�X�<&��<���<(�<��<B�<�k�<ᓋ<ƺ�<p��<��<�(�<VK�<em�<a}<_y<�u<�q<�n<�_j<o�f<8�b<�_<�`[<٢W<�S<Y*P<rpL<�H<�E<�MA<ϛ=<��9<U@6<G�2<D�.<O+<��'<C$<?� <��<b<`�<bX<��<�d<+�<щ<8&<���;V��;J�;���;6?�;���;�t�;p(�;Y��;{��;J��;���;⺯;�ݩ;��;x]�;뺘;�,�;���;�L�;���;/z{;g'q;��f;��\;�S;ngI;�?;�o6;�,-;�$;�;�;;��	;�� ;!�:?^�:A��:ʿ:�د:��:V��:FM�:�ad:��F:x):=�:�>�9K�9��Y9���8�{�mS�h]�N���tٹ�*4!��";���T�kn��䃺���)���z��gݵ�9.º[pκ?�ں���������\s�^l��a��P�K<��"#��)�{�.�[�4��:��p@��EF��L�:�Q���W��]��Qc�ni�S�n��t�z�'%���
������nֈ�e���g���J����t��+^���H���  �  Rz=�=�=�`=�=W�=�E=�� =�� =D( =��<��<a�<O�<��<��<f�<�A�<�|�<*��<���<|&�<]�<c��<���<���<+�<Q[�<��<S��<��<�<g5�<�[�<���<W��<	��<���<��<�<�0�<�E�<�X�<dh�<~u�<��<���<ʊ�<���<���<��<Ry�<l�<�Z�<F�<-�<�<���<@��<R��<�p�<�=�<C�<���<���<�B�<���<��<IS�<���<���<17�<���<a�<��<`w�<V��<�z�<)��<-k�<�ܶ<�I�<���<S�<�w�<{Ԯ<=-�<=��<�ө<�!�<-l�<���<���<69�<�w�<���<��<�#�<�X�<��<���<(�<��<B�<�k�<���<���<c��<�<�(�<[K�<`m�<v}<_y<��u<G�q< n<�_j<u�f<c�b<�_<�`[<�W<�S<q*P<lpL<�H<�E<�MA<��=<��9<Z@6</�2<O�.<�N+<��'<$<� <��<�a<Z�<&X<~�<�d<�<ω<"&<���;��;wJ�;��;C?�;���;�t�;�(�;3��;���;|��;֫�;��;�ݩ;��;�]�;c��;�,�;���;�L�;���;dz{;h'q;#�f;\�\;zS;(gI;��?;�o6;T,-;�$;�;�;;φ	;�� ;��:S\�:	��:wɿ:=د:��:���:M�:�_d:^�F:�):*�:�?�9�L�9Y�Y9��8�-x�qI��^]��L���rٹ��2!�� ;���T��in��䃺�������z��Rݵ�+/º&pκڢںU��=������s�Ym��a�KQ�r<�G##�c)�u�.���4�ؚ:�Xq@��EF��L���Q�J�W���]��Qc��i���n��t��~z��$��q
��D���cֈ����<���󋑻�t��<^���H���  �  Sz=�=�=�`=�=X�=�E=�� =�� =>( =��<��<^�<O�<ߌ�<��<]�<�A�<|�< ��<���<p&�<	]�<g��<���<���<+�<T[�<��<h��<��<�<a5�<�[�<���<V��<��<���<��<�<�0�<�E�<�X�<ph�<vu�<��<ǆ�<Ί�<���<��<��<Ny�<l�<�Z�<F�<-�<�<���<7��<[��<�p�<�=�<>�<���<È�<�B�<���<��<RS�<���<��<A7�<���<a�<��<hw�<X��<�z�<(��<&k�<�ܶ<�I�<���<U�<�w�<}Ԯ<:-�<F��<�ө<�!�<$l�<���<���<39�<�w�<���<�<�#�<�X�<��<���<*�<��<B�<�k�<䓋<���<n��<
�<�(�<fK�<am�<�}<._y<
�u<E�q<�n<�_j<n�f<��b<�_<�`[<�W<�S<�*P<ppL<&�H<�E<�MA<ԛ=<��9<^@6<�2<O�.<�N+<��'<$<� <��<�a<j�<X<��<�d<�<щ<
&<���;+��;�J�;��;6?�;���;�t�;�(�;2��;���;d��;���;]��;�ݩ;��;t]�;j��;�,�;貍;�L�;���;�z{;$'q;j�f;��\;�S;,gI;`�?;�o6;1,-;�$;�;�;;{�	;)� ;%�:�[�:���:@ɿ:�ׯ:��:w��:7M�:�`d:ЉF:�):�:�?�9�L�9�Y9w��8�w��S�7[]�TL���oٹK��3!��;���T��fn��䃺�������z���ܵ��.ºpκy�ںW����������s��m��a��Q��<�H##��)�l�.��4�̚:��q@��EF��L�G�Q��W�/�]�vQc��i���n�ҳt��~z��$���
�����rֈ�˼��_��� ����t��&^���H���  �  Uz=�=�=�`=�=U�=�E=�� =�� =?( =��<��<X�<�N�<݌�<���<^�<�A�<t|�<"��<���<z&�<�\�<e��<���<���<!+�<][�<��<[��<��<!�<w5�<�[�<���<\��<��<���<��<�<�0�<�E�<�X�<ph�<�u�<��<Ȇ�<���<���<���<��<My�<�k�<�Z�<�E�<
-�<�<���<:��<C��<�p�<�=�<D�<���<���<�B�<���<��<US�<���<ߚ�<>7�<���<a�<��<qw�<^��<�z�<4��<>k�<�ܶ<�I�<���<V�<�w�<�Ԯ<B-�<=��<�ө<�!�<-l�<���<���<,9�<�w�<���<��<�#�<�X�<	��<���<�<��<B�<�k�<ٓ�<���<k��<�<�(�<fK�<em�<w}<:_y<�u<X�q<! n<�_j<x�f<��b<�_<a[<�W<#�S<{*P<vpL<,�H<�E<�MA<ɛ=<��9<F@6<%�2<A�.<�N+<p�'<$<� <r�<�a<=�<X<l�<�d<�<ǉ<&<g��; ��;xJ�;��;Q?�;���;�t�;�(�;a��;���;���;���;b��;�ݩ;�;�]�;���;'-�;鲍;�L�;��;�z{;�'q;�f;��\;/S;gI;��?;�o6;-,-;4$;�;6;;C�	;
� ;� �:�[�:��:ɿ:�ׯ:��:���:IL�:�`d:b�F:>):w�:�A�9-L�9�Y9	��8��v�>�BW]��J��Mnٹ���0!�T;��T�zhn�䃺�~��M��xz��]ݵ��.ºqκ�ںf�����b���t��m�Fb��Q��<��##��)���.��4���:�zq@��EF�)L�]�Q�:�W���]�uQc�gi���n���t�i~z��$��R
�����^ֈ�Ѽ�����͋��st���]���H���  �  )|=�=t�=�c==��=�I=A� =r� =n- =4��<���<1�<�\�<���<���<��<DS�<���<���<d�<6<�<�s�<\��<���<��<�F�<x�<$��<���<��</�<�X�<Ȁ�<��<2��<P��<r�<h+�<�F�<L`�<w�<E��<���<{��<2��<��<���<���<��<k��<`��<���<��<h��<�s�<X�<8�<��<���<~��<e��<�T�<�<q��<���<eH�<���<6��<�J�<���<���<��<���<�=�<�ž<�H�<�ƻ<Q@�<0��<V%�<��<i��<s[�<S��<+�<l�<2��<��<�Z�<E��<�<�*�<�i�<<��<��<�<�K�<Q~�<���<�ܔ<I	�<�3�<�\�<g��<R��<ω<~�<��<Z6�<�V�<�v�<�+}<@iy<��u<��q<"n<sXj<�f<��b<�_<�H[<�W<��S<�P<�FL<�H<;�D<�A<~`=<�9<A�5<�N2<U�.<��*<�Z'<�#<�! <��<��<�n<n�<wg<��
<�w<�	<6� <���;���;�+�;F��;��;x��;N;�;y��;o��;�{�;�`�;zX�;�c�;K��;��;Z��;!Y�;ɑ;N�;��;���;��x;�_n; 7d;�7Z;y`P;)�F;`)=;0�3;I�*;v!;Q�;=�;9;��:�?�:���:Le�:*U�:=~�:��:z�:��z:d�\:/�>:D�!:��:pV�9�ӗ9��?9�a�8�Zⷲ���*t�ZH��N
�.��&���?��iY�:�r�������������BV��z�����ú%к1ܺ�D�K��@" ����
����v��@��y�#��~)��V/�`+5�	�:���@�B�F��fL�11R�G�W�z�]���c�3Ni��o�,�t�ܞz��1����������ڈ� �������g����n��U���<���  �  *|=�=u�=�c==��=�I=1� =r� =n- =@��<��<1�<�\�<|��<���<��<SS�<��<���<\�<<�<�s�<S��<���<��<�F�<x�<$��<���<��</�<�X�<̀�<��<��<Z��<l�<e+�<G�<M`�<w�<J��<ɜ�<z��<;��<���<���<���<���<o��<Z��<���<���<o��<�s�<X�<8�<��<���<z��<j��<�T�<��<k��<��<kH�<���<B��<�J�<���<���<��<���<�=�<�ž<�H�<�ƻ<X@�<��<V%�<��<e��<s[�<]��<4�<!l�<7��<��<�Z�<&��<s�<�*�<�i�<H��<�ߝ<$�<�K�<S~�<���<�ܔ<U	�<�3�<�\�<F��<G��<�Ή<{�<��<Y6�<�V�<�v�<�+}<:iy<��u<��q<%n<�Xj<ϓf<��b<�_<qH[<�W<��S<�P<�FL<��H<=�D<�A<|`=<��9<8�5<�N2<S�.<��*<�Z'<��#<�! <��<��<�n<m�<�g<��
<�w<�	<�� <���;���;�+�;b��;��;���;K;�;e��;W��;�{�;�`�;�X�;�c�;;+��;C��;Y�;(ɑ;N�;n�;���;�x;�_n;G7d;�7Z;M`P;��F;(=;K�3;�*;lv!;��;u�;>;��:O@�:ٳ�:�e�:�T�:�~�:R��:�x�:ʌz:��\:��>:�!:G�:�X�9�җ9S�?9Dg�8�i�4��>&t�	M���-��&���?��jY���r�������������U��(���H�úbк3ܺ�E��J��C" �a��
�������.��_�#�~)�MV/��+5��:���@���F�gL�K1R���W���]�.�c�2Ni�o�C�t���z��1���������]ۈ����{�������gn��$U���<���  �  #|=�=k�=�c==��=�I=4� =|� =n- =?��<��<1�<�\�<~��<���<��<[S�<���<���<p�<<�<�s�<S��<���<��<�F�<x�<��<���<��</�<�X�<π�<��<��<^��<i�<Y+�<�F�<F`�<w�<<��<���<i��<@��<���<���<���<���<���<Y��<���<���<q��<�s�<X�<8�<��<���<y��<}��<�T�<��<|��<��<pH�<���<2��<xJ�<���<���<��<���<�=�<�ž<�H�<�ƻ<]@�<��<V%�<��<b��<i[�<I��< �<l�<;��<��<�Z�</��<��<�*�<�i�<S��<�ߝ<-�<�K�<_~�<���<�ܔ<W	�<�3�<�\�<L��<Z��<ω<|�<��<F6�<�V�<�v�<�+}<,iy<��u<��q<n<�Xj<��f<��b<�_<]H[<�W<��S<�P<�FL<߉H<�D<�A<�`=<��9<[�5<�N2<}�.<��*<�Z'<	�#<�! <Ƌ<��<�n<k�<�g<��
<x<�	<� <���;���;�+�;E��;��;a��;,;�;k��;A��;�{�;q`�;�X�;�c�;���;>��;7��;�X�;ɑ;�M�;e�;y��;��x;9_n;u7d;�7Z;�`P;=�F;�(=;��3;�*;�v!;k�;��;i;&�:t@�:���:�f�:�T�:��:@�:�y�:�z:h�\:��>:��!:M�:}T�9�З90�?9B^�8������#t�CO��r乂,��&���?��kY���r�o���.���V����V��ޤ���ú-кs2ܺzD�'J��T" ���g��t�����P�#��})�>V/��+5�Z�:���@��F��fL�@1R���W��]���c��Ni�o�y�t���z�2����������ۈ�������������nn��@U���<���  �  $|=�=w�=�c==��=�I=9� =v� =w- =N��<��<;�<�\�<���<���<��<aS�<��<���<h�<)<�<�s�<S��<���<��<�F�<x�<��<���<��</�<�X�<���<ަ�<��<;��<e�<Q+�<�F�<<`�<w�<<��<Ü�<|��<9��<��<���<���<���<x��<n��<���< ��<y��<�s�<.X�<&8�<��<���<���<s��<�T�< �<g��<���<hH�<���<=��<yJ�<���<���<��<���<�=�<vž<�H�<�ƻ<>@�<��<E%�<��<X��<l[�<O��<2�<l�<7��<��<�Z�<8��<��<�*�<�i�<W��<��<2�<�K�<i~�<���<�ܔ<e	�<4�<�\�<V��<R��<�Ή<��<��<]6�<�V�<�v�<�+}<iy<��u<��q<n<UXj<Ɠf<b�b<}_<\H[<��W<��S<�P<�FL<�H<F�D<�A<�`=<�9<A�5<�N2<e�.<��*<�Z'<�#<�! <Ӌ<��<�n<��<�g<��
<x<�	<� <���;���;�+�;T��;��;z��;>;�;I��;9��;\{�;�`�;;X�;�c�;ڂ�;���;,��;�X�;�ȑ;�M�;g�;z��;Ѱx;�_n;=7d;�7Z;B`P;,�F;)=;��3;Ì*;�v!;��;Ǹ;�;w�: A�:���:g�:$V�:,�:B�:z�:y�z:B�\:��>:>�!:׿:U�9�ї9��?9iX�8������6t��N��q�A0�}&���?��kY��r�6�������2���JV�������ú^к�1ܺ�D� J���! ����
�?�����|���#��})��U/��*5���:���@�D�F�5gL�1R��W�b�]�o�c��Ni�6o���t��z�2����"���mۈ�Z���ƣ�������n��WU��=���  �  !|=�=q�=�c=	=�=�I=B� =v� =}- =P��<��<L�<�\�<���<���<��<fS�<
��<���<k�<8<�<�s�<b��<���<��<�F�<x�<��<���<��<�.�<�X�<���<Φ�<��</��<_�<A+�<�F�<1`�<�v�<4��<���<u��<1��<��<���<��<��<|��<y��<���<��<���<�s�<2X�<08�<��<���<���<y��<�T�<�<o��<���<bH�<���<-��<oJ�<���<���<��<���<�=�<kž<�H�<�ƻ<4@�<��<3%�<��<D��<a[�<@��<!�<l�<6��<��<�Z�<G��<��<�*�<�i�<Y��<��<:�<L�<l~�<Į�<
ݔ<d	�<4�<�\�<e��<]��<	ω<��<��<S6�<�V�<�v�<�+}<iy<��u<n�q<�n<1Xj<��f<=�b<w_<@H[<�W<��S<�P<�FL<ʉH</�D<�A<�`=<�9<Y�5<�N2<e�.<��*<�Z'<2�#<�! <�<�<o<��<�g<��
<)x<�	<?� <ׂ�;��;�+�;>��;��;>��;;�;���;?��;){�;S`�;X�;�c�;���;���;��;�X�;�ȑ;�M�;#�;]��;i�x;�_n;7d;O8Z;�`P;��F;V)=;��3;�*; w!;q�;2�;;��:�A�:ϵ�:g�:�V�:��:��:�z�:��z:��\:�>:G�!:�:�R�90Η9+�?9�Y�8��ⷩ��O;t�DQ����F1�� &���?��kY�k�r���������&����V��	����ú�к�0ܺ�D躘I��i! ���
�������f����#�H})��U/��*5���:��@��F��fL��0R�S�W���]��c��Ni��o���t�E�z�V2����i����ۈ�����ң��舑��n��VU��K=���  �  |=�=n�=�c==��=�I=A� =�� =|- =Y��<3��<X�<�\�<���<���<�<�S�<	��<���<��<5<�<�s�<P��<���<��<�F�<x�<��<���<��<�.�<�X�<���<���<���<2��<D�<7+�<�F�<+`�<�v�<4��<���<k��<C��<���<���<��<��<���<v��<���<��<���<t�<GX�<@8�<��<��<���<���<�T�<�<v��<��<rH�<���</��<pJ�<���<���<��<���<i=�<lž<kH�<�ƻ<-@�<<2%�<ꐵ<@��<][�<C��<�<l�<;��<��<�Z�<B��<��<�*�<�i�<t��<'��<O�<L�<�~�<Ϯ�<ݔ<s	�<4�<
]�<d��<a��<�Ή<|�<��<K6�<�V�<�v�<�+}<�hy<w�u<A�q<�n<1Xj<}�f<6�b<G_<H[<ׅW<��S<�P<uFL<ӉH<"�D<�A<�`=<��9<g�5<�N2<��.<��*<['<]�#<�! <�<�<;o<��<�g<��
<8x<�	<;� <��;���;�+�;P��;��;[��;;�; ��;��;*{�;�_�;�W�;Oc�;F��;���;���;jX�;�ȑ;�M�;�;a��;��x;Y_n;�7d;�7Z;�`P;��F;l)=;��3;�*;�w!;Æ;��;�;�:�B�:N��:�h�:�V�:
��:8�:�z�:��z:=�\::�>:;�!:A�::S�9�͗9��?9rJ�8�����9t��X����	2��$&���?�`nY���r�����\���O����V������:�ú&к1ܺEC��H���! ����	�J�������0�#��|)�_U/��*5���:��@�ȚF�!gL�@1R���W���]���c��Ni��o�-�t���z��2��x��g����ۈ�����0���R����n���U��L=���  �  |=�=k�=�c==��=�I=?� =�� =- ={��<A��<]�<�\�<���<���<�<�S�<%��<���<��<1<�<�s�<V��<���<��<�F�<x�<���<���<~�< /�<�X�<���<���<���<��<*�<>+�<�F�<`�<�v�<��<���<`��<O��<���<���<��<��<���<��<ݮ�<"��<���<t�<RX�<S8�<��</��<���<���<�T�<�<���<��<H�<���</��<\J�<���<���<�<���<O=�<Už<_H�<�ƻ<@�<ܴ�<5%�<ϐ�<;��<B[�<:��<�<l�<J��<��<�Z�<?��<��<�*�<j�<���<'��<e�<L�<�~�<֮�<%ݔ<�	�<4�<]�<c��<m��<ω<��<��<C6�<�V�<�v�<�+}<�hy<a�u<P�q<�n<Xj<Y�f<�b<_<H[<˅W<|�S<�P<CFL<։H<�D<�A<�`=<	�9<��5<�N2<��.<��*<H['<z�#<�! <C�<,�<lo<��<*h<�
<Ix<�	<5� <R��;���;1,�;?��;��;T��;�:�;���;���;:{�;�_�;�W�;.c�;��;L��;L��;�X�;jȑ;XM�;��;��;��x;_n;8d;�7Z;$aP;бF;�)=;��3;W�*;�x!;ކ;�;V;��:�C�:���:�j�:�W�:r��:��:�z�:��z:`�\:�>:�!:n�:�N�9�ȗ9��?930�8�����dDt�p[����=5��&&�R�?��qY�9�r����҅��r���+W������(�ú5кH1ܺ�B�kH���  ���	������������#�u|)�AT/�u*5�h�:��@�h�F��fL�1R���W�4�]���c��Oi�o���t��z��2���������D܈�࿋�����H���o���U��_=���  �  |=�=f�=�c==�=�I=L� =�� =�- =}��<A��<u�<�\�<Û�<���<�<�S�<3��<���<��<G<�<�s�<_��<���<��<�F�<�w�<���<���<y�<�.�<�X�<���<���<���<	��<)�< +�<�F�<`�<�v�<!��<���<`��<?��<��<���<��<"��<���<���<خ�<4��<���<t�<[X�<i8�<��<'��<���<���<�T�<�<���<���<oH�<���<��<YJ�<x��<���<n�<g��<K=�<@ž<TH�<�ƻ<@�<״�<%�<Ɛ�<5��<<[�<.��<
�<l�<>��<��<�Z�<R��<��<�*�<%j�<���<?��<w�<'L�<�~�<ﮖ<-ݔ<�	�<(4�<]�<~��<o��<ω<��<��<;6�<�V�<�v�<�+}<�hy<%�u<$�q<�n<�Wj<E�f<��b<_<�G[<��W<o�S<�P<LFL<��H< �D<�A<�`=<�9<��5<�N2<��.<"�*<N['<{�#<!" <[�<P�<�o<��<h<=�
<rx<
<d� <J��; ��;,�;0��;T�;+��;�:�;���;���;�z�;�_�;wW�;�b�;���;���;M��;X�;ȑ;AM�;��;��;-�x;_n;�7d;8Z;)aP;&�F;l*=;��3;0�*;�x!;x�;�;�;x�:QE�:��:�j�:0Y�:Ł�:	�:�{�:7�z:��\:4�>:�!:��:6N�9
Ǘ9��?9��8�t�M���Nt��]����6�&'&���?�}rY���r����}���a���oW��[�����úMк�/ܺ5B�pG��,  �S�����Y�����'�#�5|)�MT/��)5�\�:�B�@�W�F��fL��0R��W�r�]� �c��Oi�9o��t�۠z��2���������k܈�?������������o��	V��~=���  �  |=�=n�=�c==�=�I=O� =�� =�- =���<^��<��<]�<ޛ�<���<9�<�S�<>��<���<��<K<�<�s�<h��<���<��<�F�<�w�<���<k��<{�<�.�<�X�<v��<���<���<���< �<+�<�F�<	`�<�v�<%��<���<r��<6��<
��<���<��<$��<���<���<֮�<R��<���<1t�<wX�<g8�<�<'��<˽�<���<�T�<�<��<���<_H�<���<��<\J�<l��<t��<q�<K��<B=�<-ž<>H�<uƻ<�?�<ʴ�<�$�<ǐ�<��<:[�<.��<�<l�<+��<��<�Z�<R��<��<�*�<2j�<���<Z��<s�<EL�<�~�<���<Iݔ<�	�<>4�<]�<���<i��<ω<��<��<N6�<�V�<�v�<Z+}<�hy<!�u<��q<zn<�Wj<1�f<��b<�
_<�G[<}�W<p�S<nP<NFL<��H<"�D<�A<�`=<!�9<u�5<	O2<��.<E�*<Y['<��#<L" <g�<��<�o<3�<Dh<U�
<�x<
<n� <8��;I��;�+�;z��;z�;&��;�:�;e��;���;qz�;j_�;OW�;�b�;���;���;,��;�W�;/ȑ;
M�;��;1��;ϯx;�_n;E7d;K8Z;>aP;�F;�*=;$�3;َ*;�x!;h�;�;R;H�:FE�:���:�j�:DZ�:��:4�:�{�:�z:|�\:P�>:M�!:M�:ZO�9Pė9´?9�$�8 ����=Wt��b��9$�a8��(&�u�?�DrY���r����o���3���GV��w�����ú�к�/ܺ B��F��� ����%��b��L����#�N{)�?T/�)5�h�:�,�@���F�lfL�1R��W���]�w�c�vOi�o�,�t��z�Q3����[����܈�����Ԥ��㉑��o��V���=���  �  |=�=f�=�c==�=�I=R� =�� =�- =���<l��<��<]�<��<���<;�<�S�<C��<���<��<P<�<�s�<q��<���<��<}F�<�w�<��<i��<q�<�.�<tX�<g��<���<���<���<�<+�<�F�< `�<�v�<��<���<f��<7��<��<���< ��<.��<���<���<��<\��<ŋ�<=t�<�X�<p8�<�<;��<ɽ�<���<�T�< �<���< ��<cH�<���<��<NJ�<e��<k��<d�<I��<,=�<!ž<7H�<qƻ<�?�<���<�$�<���<��<.[�<"��<��<l�<3��<��<�Z�<Y��<��<�*�<3j�<���<_��<��<ML�<�~�<��<Wݔ<�	�<<4�<(]�<���<y��<#ω<��<��<>6�<�V�<�v�<T+}<�hy<�u<��q<Un<�Wj<�f<��b<�
_<�G[<v�W<U�S<lP<+FL<��H<�D<�A<�`=<;�9<��5<O2<�.<B�*<p['<Ҽ#<U" <��<��<�o<8�<ch<`�
<�x<:
<{� <w��;s��;,�;S��;N�;���;�:�;c��;i��;yz�;%_�;W�;zb�;���;���;���;�W�;ȑ;�L�;��;���;��x;H_n;W7d;r8Z;�aP;w�F;�*=;��3;Ў*;My!;��;I�;�;�:�E�:M��:�k�:0Z�:��:��:h|�:*�z:\�\:��>: �!:T�:L�9�9��?9��8���j��X\t��d���$�:�C+&�[�?��sY�N�r������������V����c�ú�кv/ܺ�@�iF��� �f������&��ʿ���#��z)��S/�)5���:���@��F� fL��0R�0�W�^�]���c��Oi�.o���t�
�z�h3��]��|����܈������������o��<V���=���  �  |=�=h�=�c== �=�I=Q� =�� =�- =���<i��<��<*]�<ڛ�<��<D�<�S�<O��<���<��<P<�<�s�<[��<���<��<�F�<�w�<��<v��<Z�<�.�<mX�<^��<{��<���<���<��<�*�<�F�<`�<�v�<��<���<c��<;��<��<���<��<*��<���<���<���<Y��<��<Gt�<�X�<�8�<�<F��<ͽ�<���<�T�<�<���<��<hH�<���<��<IJ�<f��<s��<P�<B��<=�<ž<"H�<`ƻ<�?�<���<�$�<���<��<&[�<$��<�<l�<8��<��<�Z�<X��<��<�*�<;j�<���<c��<��<AL�<�~�<��<Tݔ<�	�<@4�<1]�<���<t��<ω<��<��<?6�<�V�<�v�<f+}<�hy<�u<��q<?n<�Wj<�f<��b<�
_<�G[<U�W<7�S<�P<FL<��H<�D<�A<�`=<�9<��5<O2<��.<N�*<�['<μ#<v" <��<��<�o<K�<mh<y�
<�x<C
<|� <f��;��;,�;@��;}�;��;e:�;���;��;Gz�;_�;�V�;Lb�;R��;|��;���;�W�;�Ǒ;�L�;��;ڔ�;=�x;4_n;{7d;8Z;6aP;B�F;�*=;��3;�*;�y!;��;P�;;�:+H�:7��:�l�:rZ�:���:��:(|�:S�z:E�\:��>:F�!:�:K�92×9�?9��8:�����"`t�|i���(�;�b,&���?�@vY���r���ꆒ�����VW��������ú)кt/ܺ�@��E��q �4���������A��Ӟ#��z)�HS/��(5�y�:���@�1�F��fL��0R�6�W�X�]�<�c�RPi��o���t���z��3���������݈�����A���*����o��wV���=���  �  |=�=g�=�c=	=	�=�I=W� =�� =�- =���<s��<��<(]�<��<
��<K�<�S�<R��<���<��<`<�<�s�<m��<���<��<�F�<�w�<ڧ�<`��<\�<�.�<lX�<\��<p��<���<���<�<�*�<�F�<�_�<�v�<��<���<^��<6��<��<���<.��<4��<���<���<���<`��<��<It�<�X�<�8�<!�<K��<ֽ�<���<�T�<-�<���< ��<bH�<���<��<8J�<V��<`��<P�<7��< =�<ž<H�<Xƻ<�?�<���<�$�<���<��<[�<��< �<�k�<3��<��<�Z�<g��<��<�*�<Aj�<���<h��<��<QL�<�~�<��<[ݔ<�	�<G4�<0]�<���<���< ω<��<��<?6�<�V�<{v�<?+}<�hy<��u<��q<Bn<�Wj<�f<��b<�
_<�G[<W�W<3�S<ZP<	FL<��H<�D<�A<�`=<0�9<��5<)O2<�.<\�*<�['<�#<~" <��<��<�o<Y�<�h<��
<�x<E
<�� <���;h��;,�;=��;_�;ϝ�;M:�;E��;��;=z�;_�;�V�;$b�;>��;_��;���;nW�;�Ǒ;�L�;K�;���;��x;_n;S7d;�8Z;�aP;�F;+=;�3;)�*;�y!;�;(�;;z�:�G�:���:�l�:[�:	��:L�:Q}�:}�z:t�\:��>:��!:��:�F�92��9��?9W�8�%����bt��j���*�\;�,&���?�vY�g�r����1�������yW��ͤ����ú\к�.ܺ�@�oE��A �����������A��֞#��z)�ES/��(5���:���@���F�fL��0R�Q�W�W�]�ˉc��Pi��o���t���z��3���������݈����>���C����o��~V��>���  �  |=�=i�=�c==�=�I=W� =�� =�- =���<��<��<$]�<��<���<K�<�S�<H��< ��<��<_<�<�s�<o��<���<��<�F�<�w�<���<_��<b�<�.�<]X�<W��<p��<���<���<�<�*�<�F�<�_�<�v�< ��<���<j��<0��<��<���<$��<3��<���<���<���<p��<׋�<St�<�X�<�8�<.�<O��<Խ�<���<�T�<$�<���< ��<]H�<���<��<PJ�<h��<Z��<T�<,��<=�<ž<H�<Wƻ<�?�<���<�$�<���<��<<[�< ��<�<l�<*��<��<�Z�<d��<��<�*�<7j�<���<l��<��<kL�<�~�<��<jݔ<�	�<J4�<4]�<���<y��<ω<��<��<E6�<�V�<�v�<I+}<�hy<�u<��q<An<yWj<��f<}�b<�
_<uG[<E�W<1�S<_P<IFL<��H<�D<�A<�`=<-�9<��5<*O2<��.<a�*<�['<��#<v" <��<��<�o<Z�<�h<n�
<�x<O
<�� <d��;o��;�+�;Q��;u�;��;�:�;B��;3��;z�;�^�;�V�;"b�;L��;J��;���;<W�;�Ǒ;�L�;��;$��;̯x;r_n;&7d;~8Z;|aP;��F;+=;,�3;L�*;�y!;c�;ܻ;k;y�:6G�:W��:m�:�Z�:���:e�:�|�:�z:h�\:G�>:L�!:`�:�L�9�×9��?9�	�8#O�t��Set�;j���*�2<�L-&���?�ZuY���r�������v����V��c�����ú0к�.ܺr@�eE��� ���s���-��H����#�Ez)�lS/��(5�[�:���@��F�<fL��0R�d�W�!�]���c��Oi�Yo��t���z��3��������� ݈����?���x���p���V��>���  �  |=�=g�=�c=	=	�=�I=W� =�� =�- =���<s��<��<(]�<��<
��<K�<�S�<R��<���<��<`<�<�s�<m��<���<��<�F�<�w�<ڧ�<`��<\�<�.�<lX�<\��<p��<���<���<�<�*�<�F�<�_�<�v�<��<���<^��<6��<��<���<.��<4��<���<���<���<`��<��<It�<�X�<�8�<!�<K��<ֽ�<���<�T�<-�<���< ��<bH�<���<��<8J�<V��<`��<P�<7��< =�<ž<H�<Xƻ<�?�<���<�$�<���<��<[�<��< �<�k�<3��<��<�Z�<g��<��<�*�<Aj�<���<h��<��<QL�<�~�<��<[ݔ<�	�<G4�<0]�<���<���< ω<��<��<?6�<�V�<{v�<?+}<�hy<��u<��q<Bn<�Wj<�f<��b<�
_<�G[<W�W<3�S<ZP<	FL<��H<�D<�A<�`=<0�9<��5<)O2<�.<\�*<�['<�#<~" <��<��<�o<Y�<�h<��
<�x<E
<�� <���;h��;,�;=��;_�;ϝ�;M:�;E��;��;=z�;_�;�V�;$b�;>��;_��;���;nW�;�Ǒ;�L�;K�;���;��x;_n;S7d;�8Z;�aP;�F;+=;�3;)�*;�y!;�;(�;;z�:�G�:���:�l�:[�:	��:L�:Q}�:}�z:t�\:��>:��!:��:�F�92��9��?9W�8�%����bt��j���*�\;�,&���?�vY�g�r����1�������yW��ͤ����ú\к�.ܺ�@�oE��A �����������A��֞#��z)�ES/��(5���:���@���F�fL��0R�Q�W�W�]�ˉc��Pi��o���t���z��3���������݈����>���C����o��~V��>���  �  |=�=h�=�c== �=�I=Q� =�� =�- =���<i��<��<*]�<ڛ�<��<D�<�S�<O��<���<��<P<�<�s�<[��<���<��<�F�<�w�<��<v��<Z�<�.�<mX�<^��<{��<���<���<��<�*�<�F�<`�<�v�<��<���<c��<;��<��<���<��<*��<���<���<���<Y��<��<Gt�<�X�<�8�<�<F��<ͽ�<���<�T�<�<���<��<hH�<���<��<IJ�<f��<s��<P�<B��<=�<ž<"H�<`ƻ<�?�<���<�$�<���<��<&[�<$��<�<l�<8��<��<�Z�<X��<��<�*�<;j�<���<c��<��<AL�<�~�<��<Tݔ<�	�<@4�<1]�<���<t��<ω<��<��<?6�<�V�<�v�<f+}<�hy<�u<��q<?n<�Wj<�f<��b<�
_<�G[<U�W<7�S<�P<FL<��H<�D<�A<�`=<�9<��5<O2<��.<N�*<�['<μ#<v" <��<��<�o<K�<mh<y�
<�x<C
<|� <f��;��;,�;@��;}�;��;e:�;���;��;Gz�;_�;�V�;Lb�;R��;|��;���;�W�;�Ǒ;�L�;��;ڔ�;=�x;4_n;{7d;8Z;6aP;B�F;�*=;��3;�*;�y!;��;P�;;�:+H�:7��:�l�:rZ�:���:��:(|�:S�z:E�\:��>:F�!:�:K�92×9�?9��8:�����"`t�|i���(�;�b,&���?�@vY���r���ꆒ�����VW��������ú)кt/ܺ�@��E��q �4���������A��Ӟ#��z)�HS/��(5�y�:���@�1�F��fL��0R�6�W�X�]�<�c�RPi��o���t���z��3���������݈�����A���*����o��wV���=���  �  |=�=f�=�c==�=�I=R� =�� =�- =���<l��<��<]�<��<���<;�<�S�<C��<���<��<P<�<�s�<q��<���<��<}F�<�w�<��<i��<q�<�.�<tX�<g��<���<���<���<�<+�<�F�< `�<�v�<��<���<f��<7��<��<���< ��<.��<���<���<��<\��<ŋ�<=t�<�X�<p8�<�<;��<ɽ�<���<�T�< �<���< ��<cH�<���<��<NJ�<e��<k��<d�<I��<,=�<!ž<7H�<qƻ<�?�<���<�$�<���<��<.[�<"��<��<l�<3��<��<�Z�<Y��<��<�*�<3j�<���<_��<��<ML�<�~�<��<Wݔ<�	�<<4�<(]�<���<y��<#ω<��<��<>6�<�V�<�v�<T+}<�hy<�u<��q<Un<�Wj<�f<��b<�
_<�G[<v�W<U�S<lP<+FL<��H<�D<�A<�`=<;�9<��5<O2<�.<B�*<p['<Ҽ#<U" <��<��<�o<8�<ch<`�
<�x<:
<{� <w��;s��;,�;S��;N�;���;�:�;c��;i��;yz�;%_�;W�;zb�;���;���;���;�W�;ȑ;�L�;��;���;��x;H_n;W7d;r8Z;�aP;w�F;�*=;��3;Ў*;My!;��;I�;�;�:�E�:M��:�k�:0Z�:��:��:h|�:*�z:\�\:��>: �!:T�:L�9�9��?9��8���j��X\t��d���$�:�C+&�[�?��sY�N�r������������V����c�ú�кv/ܺ�@�iF��� �f������&��ʿ���#��z)��S/�)5���:���@��F� fL��0R�0�W�^�]���c��Oi�.o���t�
�z�h3��]��|����܈������������o��<V���=���  �  |=�=n�=�c==�=�I=O� =�� =�- =���<^��<��<]�<ޛ�<���<9�<�S�<>��<���<��<K<�<�s�<h��<���<��<�F�<�w�<���<k��<{�<�.�<�X�<v��<���<���<���< �<+�<�F�<	`�<�v�<%��<���<r��<6��<
��<���<��<$��<���<���<֮�<R��<���<1t�<wX�<g8�<�<'��<˽�<���<�T�<�<��<���<_H�<���<��<\J�<l��<t��<q�<K��<B=�<-ž<>H�<uƻ<�?�<ʴ�<�$�<ǐ�<��<:[�<.��<�<l�<+��<��<�Z�<R��<��<�*�<2j�<���<Z��<s�<EL�<�~�<���<Iݔ<�	�<>4�<]�<���<i��<ω<��<��<N6�<�V�<�v�<Z+}<�hy<!�u<��q<zn<�Wj<1�f<��b<�
_<�G[<}�W<p�S<nP<NFL<��H<"�D<�A<�`=<!�9<u�5<	O2<��.<E�*<Y['<��#<L" <g�<��<�o<3�<Dh<U�
<�x<
<n� <8��;I��;�+�;z��;z�;&��;�:�;e��;���;qz�;j_�;OW�;�b�;���;���;,��;�W�;/ȑ;
M�;��;1��;ϯx;�_n;E7d;K8Z;>aP;�F;�*=;$�3;َ*;�x!;h�;�;R;H�:FE�:���:�j�:DZ�:��:4�:�{�:�z:|�\:P�>:M�!:M�:ZO�9Pė9´?9�$�8 ����=Wt��b��9$�a8��(&�u�?�DrY���r����o���3���GV��w�����ú�к�/ܺ B��F��� ����%��b��L����#�N{)�?T/�)5�h�:�,�@���F�lfL�1R��W���]�w�c�vOi�o�,�t��z�Q3����[����܈�����Ԥ��㉑��o��V���=���  �  |=�=f�=�c==�=�I=L� =�� =�- =}��<A��<u�<�\�<Û�<���<�<�S�<3��<���<��<G<�<�s�<_��<���<��<�F�<�w�<���<���<y�<�.�<�X�<���<���<���<	��<)�< +�<�F�<`�<�v�<!��<���<`��<?��<��<���<��<"��<���<���<خ�<4��<���<t�<[X�<i8�<��<'��<���<���<�T�<�<���<���<oH�<���<��<YJ�<x��<���<n�<g��<K=�<@ž<TH�<�ƻ<@�<״�<%�<Ɛ�<5��<<[�<.��<
�<l�<>��<��<�Z�<R��<��<�*�<%j�<���<?��<w�<'L�<�~�<ﮖ<-ݔ<�	�<(4�<]�<~��<o��<ω<��<��<;6�<�V�<�v�<�+}<�hy<%�u<$�q<�n<�Wj<E�f<��b<_<�G[<��W<o�S<�P<LFL<��H< �D<�A<�`=<�9<��5<�N2<��.<"�*<N['<{�#<!" <[�<P�<�o<��<h<=�
<rx<
<d� <J��;��;,�;/��;T�;+��;�:�;���;���;�z�;�_�;wW�;�b�;���;���;M��;X�;ȑ;AM�;��;��;-�x;_n;�7d;8Z;)aP;&�F;l*=;��3;0�*;�x!;x�;�;�;x�:QE�:��:�j�:0Y�:Ł�:	�:�{�:7�z:��\:4�>:�!:��:6N�9
Ǘ9��?9��8�t�M���Nt��]����6�&'&���?�}rY���r����}���a���oW��[�����úMк�/ܺ5B�pG��,  �S�����Y�����'�#�5|)�MT/��)5�\�:�B�@�W�F��fL��0R��W�r�]� �c��Oi�9o��t�۠z��2���������k܈�?������������o��	V��~=���  �  |=�=k�=�c==��=�I=?� =�� =- ={��<A��<]�<�\�<���<���<�<�S�<%��<���<��<1<�<�s�<V��<���<��<�F�<x�<���<���<~�< /�<�X�<���<���<���<��<*�<>+�<�F�<`�<�v�<��<���<`��<O��<���<���<��<��<���<��<ݮ�<"��<���<t�<RX�<S8�<��</��<���<���<�T�<�<���<��<H�<���</��<\J�<���<���<�<���<O=�<Už<_H�<�ƻ<@�<ܴ�<5%�<ϐ�<;��<B[�<:��<�<l�<J��<��<�Z�<?��<��<�*�<j�<���<'��<e�<L�<�~�<֮�<%ݔ<�	�<4�<]�<c��<m��<ω<��<��<C6�<�V�<�v�<�+}<�hy<a�u<P�q<�n<Xj<Y�f<�b<_<H[<˅W<|�S<�P<CFL<։H<�D<�A<�`=<	�9<��5<�N2<��.<��*<H['<z�#<�! <C�<,�<lo<��<*h<�
<Ix<�	<5� <R��;���;1,�;?��;��;S��;�:�;���;���;:{�;�_�;�W�;.c�;��;L��;L��;�X�;jȑ;XM�;��;��;��x;_n;8d;�7Z;$aP;бF;�)=;��3;W�*;�x!;ކ;�;V;��:�C�:���:�j�:�W�:r��:��:�z�:��z:`�\:�>:�!:n�:�N�9�ȗ9��?930�8�����dDt�p[����=5��&&�R�?��qY�9�r����҅��r���+W������(�ú5кH1ܺ�B�kH���  ���	������������#�u|)�AT/�u*5�h�:��@�h�F��fL�1R���W�4�]���c��Oi�o���t��z��2���������D܈�࿋�����H���o���U��_=���  �  |=�=n�=�c==��=�I=A� =�� =|- =Y��<3��<X�<�\�<���<���<�<�S�<	��<���<��<5<�<�s�<P��<���<��<�F�<x�<��<���<��<�.�<�X�<���<���<���<2��<D�<7+�<�F�<+`�<�v�<4��<���<k��<C��<���<���<��<��<���<v��<���<��<���<t�<GX�<@8�<��<��<���<���<�T�<�<v��<��<rH�<���</��<pJ�<���<���<��<���<i=�<lž<kH�<�ƻ<-@�<<2%�<ꐵ<@��<][�<C��<�<l�<;��<��<�Z�<B��<��<�*�<�i�<t��<'��<O�<L�<�~�<Ϯ�<ݔ<s	�<4�<
]�<d��<a��<�Ή<|�<��<K6�<�V�<�v�<�+}<�hy<w�u<A�q<�n<1Xj<}�f<6�b<G_<H[<ׅW<��S<�P<uFL<ӉH<"�D<�A<�`=<��9<g�5<�N2<��.<��*<['<]�#<�! <�<�<;o<��<�g<��
<8x<�	<;� <��;���;�+�;P��;��;[��;;�; ��;��;*{�;�_�;�W�;Oc�;F��;���;���;jX�;�ȑ;�M�;�;a��;��x;Y_n;�7d;�7Z;�`P;��F;l)=;��3;�*;�w!;Æ;��;�;�:�B�:N��:�h�:�V�:
��:8�:�z�:��z:=�\::�>:;�!:A�::S�9�͗9��?9rJ�8�����9t��X����	2��$&���?�`nY���r�����\���O����V������:�ú&к1ܺEC��H���! ����	�J�������0�#��|)�_U/��*5���:��@�ȚF�!gL�@1R���W���]���c��Ni��o�-�t���z��2��x��g����ۈ�����0���R����n���U��L=���  �  !|=�=q�=�c=	=�=�I=B� =v� =}- =P��<��<L�<�\�<���<���<��<fS�<
��<���<k�<8<�<�s�<b��<���<��<�F�<x�<��<���<��<�.�<�X�<���<Φ�<��</��<_�<A+�<�F�<1`�<�v�<4��<���<u��<1��<��<���<��<��<|��<y��<���<��<���<�s�<2X�<08�<��<���<���<y��<�T�<�<o��<���<bH�<���<-��<oJ�<���<���<��<���<�=�<kž<�H�<�ƻ<4@�<��<3%�<��<D��<a[�<@��<!�<l�<6��<��<�Z�<G��<��<�*�<�i�<Y��<��<:�<L�<l~�<Į�<
ݔ<d	�<4�<�\�<e��<]��<	ω<��<��<S6�<�V�<�v�<�+}<iy<��u<n�q<�n<1Xj<��f<=�b<w_<@H[<�W<��S<�P<�FL<ʉH</�D<�A<�`=<�9<Y�5<�N2<e�.<��*<�Z'<2�#<�! <�<�<o<��<�g<��
<)x<�	<?� <ׂ�;��;�+�;>��;��;>��;;�;���;?��;){�;S`�;X�;�c�;���;���;��;�X�;�ȑ;�M�;#�;]��;i�x;�_n;7d;O8Z;�`P;��F;V)=;��3;�*; w!;q�;2�;;��:�A�:ϵ�:g�:�V�:��:��:�z�:��z:��\:�>:G�!:�:�R�90Η9+�?9�Y�8��ⷩ��O;t�DQ����F1�� &���?��kY�k�r���������&����V��	����ú�к�0ܺ�D躘I��i! ���
�������f����#�H})��U/��*5���:��@��F��fL��0R�S�W���]��c��Ni��o���t�E�z�V2����i����ۈ�����ң��舑��n��VU��K=���  �  $|=�=w�=�c==��=�I=9� =v� =w- =N��<��<;�<�\�<���<���<��<aS�<��<���<h�<)<�<�s�<S��<���<��<�F�<x�<��<���<��</�<�X�<���<ަ�<��<;��<e�<Q+�<�F�<<`�<w�<<��<Ü�<|��<9��<��<���<���<���<x��<n��<���< ��<y��<�s�<.X�<&8�<��<���<���<s��<�T�< �<g��<���<hH�<���<=��<yJ�<���<���<��<���<�=�<vž<�H�<�ƻ<>@�<��<E%�<��<X��<l[�<O��<2�<l�<7��<��<�Z�<8��<��<�*�<�i�<W��<��<2�<�K�<i~�<���<�ܔ<e	�<4�<�\�<V��<R��<�Ή<��<��<]6�<�V�<�v�<�+}<iy<��u<��q<n<UXj<Ɠf<b�b<}_<\H[<��W<��S<�P<�FL<�H<F�D<�A<�`=<�9<A�5<�N2<e�.<��*<�Z'<�#<�! <Ӌ<��<�n<��<�g<��
<x<�	<� <���;���;�+�;T��;��;z��;>;�;I��;9��;\{�;�`�;;X�;�c�;ڂ�;���;,��;�X�;�ȑ;�M�;g�;z��;Ѱx;�_n;=7d;�7Z;B`P;,�F;)=;��3;Ì*;�v!;��;Ǹ;�;w�: A�:���:g�:$V�:,�:B�:z�:y�z:B�\:��>:>�!:׿:U�9�ї9��?9iX�8������6t��N��q�A0�}&���?��kY��r�6�������2���JV�������ú^к�1ܺ�D� J���! ����
�?�����|���#��})��U/��*5���:���@�D�F�5gL�1R��W�b�]�o�c��Ni�6o���t��z�2����"���mۈ�Z���ƣ�������n��WU��=���  �  #|=�=k�=�c==��=�I=4� =|� =n- =?��<��<1�<�\�<~��<���<��<[S�<���<���<p�<<�<�s�<S��<���<��<�F�<x�<��<���<��</�<�X�<π�<��<��<^��<i�<Y+�<�F�<F`�<w�<<��<���<i��<@��<���<���<���<���<���<Y��<���<���<q��<�s�<X�<8�<��<���<y��<}��<�T�<��<|��<��<pH�<���<2��<xJ�<���<���<��<���<�=�<�ž<�H�<�ƻ<]@�<��<V%�<��<b��<i[�<I��< �<l�<;��<��<�Z�</��<��<�*�<�i�<S��<�ߝ<-�<�K�<_~�<���<�ܔ<W	�<�3�<�\�<L��<Z��<ω<|�<��<F6�<�V�<�v�<�+}<,iy<��u<��q<n<�Xj<��f<��b<�_<]H[<�W<��S<�P<�FL<߉H<�D<�A<�`=<��9<[�5<�N2<}�.<��*<�Z'<	�#<�! <Ƌ<��<�n<k�<�g<��
<x<�	<� <���;���;�+�;E��;��;a��;,;�;k��;A��;�{�;q`�;�X�;�c�;���;>��;7��;�X�;ɑ;�M�;e�;y��;��x;9_n;u7d;�7Z;�`P;=�F;�(=;��3;�*;�v!;k�;��;i;&�:t@�:���:�f�:�T�:��:@�:�y�:�z:h�\:��>:��!:M�:}T�9�З90�?9B^�8������#t�CO��r乂,��&���?��kY���r�o���.���V����V��ޤ���ú-кs2ܺzD�'J��T" ���g��t�����P�#��})�>V/��+5�Z�:���@��F��fL�@1R���W��]���c��Ni�o�y�t���z�2����������ۈ�������������nn��@U���<���  �  *|=�=u�=�c==��=�I=1� =r� =n- =@��<��<1�<�\�<|��<���<��<SS�<��<���<\�<<�<�s�<S��<���<��<�F�<x�<$��<���<��</�<�X�<̀�<��<��<Z��<l�<e+�<G�<M`�<w�<J��<ɜ�<z��<;��<���<���<���<���<o��<Z��<���<���<o��<�s�<X�<8�<��<���<z��<j��<�T�<��<k��<��<kH�<���<B��<�J�<���<���<��<���<�=�<�ž<�H�<�ƻ<X@�<��<V%�<��<e��<s[�<]��<4�<!l�<7��<��<�Z�<&��<s�<�*�<�i�<H��<�ߝ<$�<�K�<S~�<���<�ܔ<U	�<�3�<�\�<F��<G��<�Ή<{�<��<Y6�<�V�<�v�<�+}<:iy<��u<��q<%n<�Xj<ϓf<��b<�_<qH[<�W<��S<�P<�FL<��H<=�D<�A<|`=<��9<8�5<�N2<S�.<��*<�Z'<��#<�! <��<��<�n<m�<�g<��
<�w<�	<�� <���;���;�+�;b��;��;���;K;�;e��;W��;�{�;�`�;�X�;�c�;;+��;C��;Y�;(ɑ;N�;n�;���;�x;�_n;G7d;�7Z;M`P;��F;(=;K�3;�*;lv!;��;u�;>;��:O@�:ٳ�:�e�:�T�:�~�:R��:�x�:ʌz:��\:��>:�!:G�:�X�9�җ9S�?9Dg�8�i�4��>&t�	M���-��&���?��jY���r�������������U��(���H�úbк3ܺ�E��J��C" �a��
�������.��_�#�~)�MV/��+5��:���@���F�gL�K1R���W���]�.�c�2Ni�o�C�t���z��1���������]ۈ����{�������gn��$U���<���  �  ~=!!=�=�f=i	=��=�M=�� =e� =�2 =���<a��<u*�<�j�<���<���<�'�<be�<��<���<��<�R�<a��<4��<���</�<;c�<���<c��<P��<�%�<�R�<�}�<6��<���<���<^�</:�<�Y�<�v�<���<h��<V��<���<���<{��<���<@�<S�<�<"�<���<y��<f��<i��<A��<��<M��<-b�<�:�<E�<0��<^��<ul�<�,�<���<���<>N�<���< ��<A�<���<bs�<��<��<$�<J��<q�<���<D�<r�<4ܵ<�A�<@��<V �<TY�<Q��<v��<�L�<���<ݦ<8 �<`�<��<$ן<��<cC�<�u�<�<�Ӗ<���<�)�<NR�<�x�<'��<���</�<p�<�%�<�D�<�b�<���<�:}<�sy<��u<!�q<n<�Pj<чf<ξb<|�^<�.[<�gW<?�S<��O<�L<�YH<W�D<7�@<�"=<Qj9<�5<�2<�S.<g�*<� '<u]#<z�<�#<g�<�<s<��<�n
<s�<
�<A <�d�;��;E��;b�;1��;�Z�;��;Ҙ�;�R�;��;���;��;���;*�;�D�;���;�;hQ�;PՊ;n�;L�;K�u;{pk;jKa;`PW;�}M;��C;3T:;%�0;	�';��;��;&;�t;M��:�?�:���:��:���:��:�n�:'$�:�r:�YT:��6:��:�|�9���9ɹ�9�$9<[8&9W��Y!�����Xú� ��� =+�+�D�2(^��Xw�Z/������m����D��?~��Чź��Ѻ��ݺ�麫����� �t�����7��As��N�@&$���)���/�0�5��d;��,A�X�F�+�L�_|R�?X�c ^�M�c��i��@o���t�w�z�k?��p������!���j���Ϣ��ᄑ��g���K���0���  �  ~=)!=�=�f=c	=��=�M=�� =b� =�2 =Χ�<i��<p*�<�j�<���<���<�'�<qe�< ��<���<��<�R�<q��<)��<���<"/�<>c�<��<g��<T��<�%�<�R�<�}�<.��<���<���<b�<:�<�Y�<�v�<���<n��<]��<���<���<���<���<F�<O�<��<$�<���<���<p��<k��<T��<���<Q��<3b�<�:�<H�<2��<=��<jl�<�,�<���<���<@N�<���<
��<	A�<���<cs�<��<���<$�<=��<g�<���<"�<�q�<1ܵ<�A�<E��<b �<YY�<T��<v��<�L�<���<ݦ<  �<`�<��<3ן<��<kC�<�u�<���<�Ӗ<���<*�<SR�<�x�<	��<���</�<c�<�%�<�D�<c�<���<�:}<�sy<��u<�q<�n<�Pj<��f<վb<h�^<�.[<�gW<4�S<��O<�L<�YH<b�D<B�@<r"=<Jj9<��5<�2<�S.<y�*<'<�]#<o�<	$<�<�<s<��<�n
<��<�< <�d�;��;6��;!b�;>��; [�;!��;��;�R�;v�;��;u�;���;��;�D�;<��;��;hQ�;<Պ;n�;l�;��u;�pk;�Ka;�OW;~M;��C;@S:;8�0;�';:�;#�;5;@u;���:@�:6��:��:槶:��:�l�:#�:�r:<XT:Y�6:V�:�~�9K��9޺�9��$9R>[8�KW��i!������ƺ�~���CA+�D�D�{(^��Xw��.����������D��@~����ź��Ѻ��ݺ���L���� �����������r�oN�l&$�s�)���/��5��d;��-A��F�)�L��|R��>X�= ^���c��i��@o� u���z��?���������Y���[�������0���h���K���0���  �  ~='!=�=�f=d	=��=�M=�� =n� =�2 =���<l��<q*�<�j�<���<���<�'�<re�<��<���<��<�R�<���<&��<���< /�<5c�<��<X��<J��<�%�<�R�<�}�<2��<���<���<n�<:�<�Y�<�v�<��<g��<Q��<���<���<���<���<L�<b�< �<<�<���<���<y��<m��<S��<���<S��<9b�<�:�<7�<D��<M��<|l�<�,�<���<���<8N�<���<���<A�<���<_s�<��<���<,�<2��<`�<���<#�<�q�<)ܵ<�A�<8��<\ �<RY�<P��<{��<�L�<���<ݦ<2 �<#`�<��<5ן<��<oC�<�u�<��<�Ӗ<���< *�<GR�<y�<��<���<2�<b�<�%�<�D�<�b�<��<�:}<�sy<��u<�q<�n<�Pj<��f<Ӿb<f�^<�.[<�gW< �S<��O<�L<�YH<O�D<>�@<t"=<Jj9<$�5<�2<�S.<l�*<� '<�]#<q�<$<u�<&�<!s<��<�n
<��<�<9 <&e�;ݩ�;K��;b�;��;[�;���;���;�R�;��;��;��;���;��;�D�;8��;��;dQ�;Պ;n�;;�;i�u;6pk;�Ka;�OW;8~M;2�C;�S:;��0;��';�;k�;P;:u;}��::@�:���:ٜ�:ᦶ:�:�m�:�$�:r:�WT:|�6:`�:}�9���9���9%�$9�6[8�FW��i!�g���ɺ�3�
��&A+���D�z)^��Yw��/�����|����D���}���ź��Ѻ��ݺ�������� �������֒��r�MN�g&$�G�)�S�/�e�5��c;�*-A�q�F��L��|R��>X�� ^���c�Z�i��@o�g u�¿z��?�������������_�������*���h���K���0���  �  ~=$!=�=�f=h	=��=�M=�� =j� =�2 =ԧ�<���<�*�<�j�<���<���<(�<�e�<%��<���<��<�R�<l��<3��<���</�<>c�<���<^��<G��<�%�<yR�<�}�<��<���<���<F�<:�<�Y�<�v�<��<f��<O��<���<���<u��<��<>�<Z�<�<5�<���<���<���<���<_��<��<j��<Pb�<�:�<T�<>��<S��<yl�<�,�<���<���<?N�<���<���< A�<���<Ss�<��<��<�<-��<R�<���<�<�q�<ܵ<�A�<:��<T �<YY�<N��<r��<�L�<���<ݦ<1 �<#`�<��<Dן<��<�C�<�u�<��<Ԗ< �<*�<]R�<y�<"��<���<.�<p�<�%�<�D�<�b�<���<�:}<�sy<��u<��q<�n<�Pj<��f<��b<1�^<�.[<�gW<�S<��O<�L<�YH<_�D<*�@<�"=<Oj9<��5<�2<�S.<��*<'<�]#<��<2$<��<L�<Zs<�<�n
<��<�<J <�d�;��;D��;b�;G��;�Z�;��;���;�R�;%�;���;��;W��;��;aD�;��;{�;7Q�;Պ;n�;7�;��u;�pk;DKa;�PW;�}M;��C;T:;��0;��';m�;�;;�u;m��:�A�:��:���:Ĩ�:��:5n�:�$�:�r:^ZT:��6:S�:�}�9���9��9�$9�![8C}W�m!�p��!ʺ�*!ﹺ��B+�,�D��*^�Zw��/��y��� ����D��e~���ź%�Ѻw�ݺ��麵���:� �i�����0��br��M��%$���)���/���5��c;��,A���F�0�L�a|R�>?X�M ^��c�;�i��@o�| u�=�z��?�� ��8 ����������e���p���ch��L���0���  �  ~=!=�=�f=g	=ī=�M=�� =m� =�2 =��<���<�*�< k�<���<���<
(�<�e�<;��<��<��<�R�<w��<A��<���</�<4c�<��<T��<1��<�%�<gR�<�}�<��<���<x��<6�<:�<�Y�<�v�<ӑ�<U��<F��<{��<���<o��<��<J�<j�<�<;�<���<���<���<���<r��<��<r��<Ub�<�:�<m�<I��<]��<�l�<�,�<���<x��<?N�<���<��<�@�<���<Is�<��<��<��<��<A�<���<�<�q�<ܵ<�A�<+��<? �<IY�<O��<i��<�L�<���<*ݦ<7 �<:`�<6��<Bן<��<�C�<�u�<��<Ԗ< �<*�<yR�<	y�<1��<���<;�<p�<z%�<�D�<�b�<{��<�:}<sy<i�u<��q<�n<|Pj<p�f<�b<4�^<�.[<�gW<��S<y�O<�L<gYH<X�D<'�@<�"=<kj9<�5<�2<�S.<ɨ*<1'<�]#<��<Q$<͎<d�<es<�<�n
<��<�<m <e�;V��;/��;b�;%��;�Z�;���;a��;�R�;��;���;��;��;��;&D�;!��;S�;
Q�;�Ԋ;�m�;�;۾u;�pk;Ka;�PW;3~M;y�C;pT:;��0;V�';��;-�;X;8v;���:CB�:l��: ��:`��:��:�n�:�%�:#r:�[T:
�6:}�:y�9���9���9�}$9j[8�W�;m!�c���ͺ�/%�p���B+�x�D��+^��\w�e0�����������D���~���ź}�Ѻo�ݺb��D���s� �t�����ۑ��q�qM�N%$���)�a�/�ԗ5��c;�e,A���F�ʸL�b|R�k?X�` ^���c�z�i��Ao�� u���z�@�����| �������\��������h��<L��91���  �  �}=!=�=�f=f	=ë=�M=�� =|� =�2 =��<���<�*�<k�<Ū�<���<%(�<�e�<;��<��<��<�R�<���<4��<���</�<*c�<��<I��<)��<�%�<]R�<�}�< ��<���<W��<4�<�9�<tY�<�v�<ɑ�<N��<E��<|��<���<|��<���<X�<m�<�<[�<���<���<���<���<���<+��<���<ub�<�:�<_�<g��<j��<�l�<�,�<���<���<1N�<���<��<�@�<���<-s�<��<���<��<���<'�<{��<��<�q�<�۵<�A�<��<D �<AY�<H��<o��<�L�<���<&ݦ<I �<K`�<0��<gן<��<�C�<v�<4��</Ԗ<- �<.*�<oR�<(y�<1��<���<A�<l�<�%�<�D�<�b�<u��<�:}<asy<?�u<��q<�n<jPj<(�f<d�b<��^<D.[<}gW<ءS<m�O<�L<wYH<>�D<2�@<~"=<gj9<$�5<�2<.T.<��*<D'<^#<�<�$<ڎ<��<�s<e�<�n
<��<N�<h <Ae�;(��;K��;b�;��;�Z�;���;H��;DR�;��;b��;��;���;�;"D�;u��;�;�P�;�Ԋ;�m�;�;�u;&pk;�Ka;TPW;�~M;��C;�T:;�0;��';��;;�;$;�v;���:�C�:x��:��:���:��:�o�:�%�:$ r:7YT:��6:��:�x�9���9.��9Ly$9b�Z8I�W���!�E��Vպ�+�]���G+���D�H.^��]w�1��H���E���E��k~���ź��Ѻ��ݺ4������� �H�������nq��L�|$$�v�)���/�&�5��b;�d,A�W�F���L��|R�?X�� ^���c���i��Ao�ou�H�z��@��� ��� ��oሻ:�ˣ�������h���L��Q1���  �  �}=!=�=�f=h	=ƫ=�M=�� =�� =�2 =
��<���<�*�<5k�<��<���<%(�<�e�<R��<��<��<�R�<���<5��<���</�<*c�<��<,��<*��<s%�<UR�<l}�<ަ�<���<C��<�<�9�<rY�<�v�<đ�<:��<,��<���<���<���<���<d�<u�<�<m�<���<���<���<���<���<E��<���<pb�<�:�<q�<w��<l��<�l�<�,�<���<���<#N�<���<֟�<�@�<���<s�<��<���<��<晽<�<Z��<��<�q�<�۵<�A�<��<7 �<AY�<>��<y��<�L�<ϖ�<)ݦ<Q �<Z`�<D��<zן<��<�C�<v�<P��<;Ԗ<2 �<L*�<�R�<7y�<4��<���<G�<l�<�%�<�D�<�b�<W��<�:}<?sy<�u<��q<En<IPj<��f<H�b<��^<..[<`gW<��S<e�O<gL<wYH</�D<1�@<�"=<qj9<K�5<�2<HT.<�*<�'<!^#<��<�$<�<��<�s<��<o
<�<i�<t <�e�;1��;v��;b�;	��;�Z�;N��;R��;�Q�;��;��;L�;���;��;�C�;���;�;RP�;�Ԋ;am�;��;%�u;�ok;�Ka;FPW;M;��C;�T:;��0;��';s�;7�;�;�w;B��:GE�:B��:���:���:��:�o�:�%�:"r:�XT:��6:f�:Az�9���9���9 y$9R�Z8߽W�N�!���vں�./�B���J+�[�D�-2^��]w��2�����*����E���}��"�źb�ѺU�ݺ���&����� �������;���p��K�$$�J�)���/���5�_b;�O,A���F�p�L�~|R��>X�^��c���i�Bo��u���z��@��!��� ���ሻr�W���*���i���L��`1���  �  �}=!=	�=�f=i	=ɫ=�M=�� =�� =�2 =��<���<�*�<Bk�<���<��<G(�<�e�<f��<,��<��<�R�<���<?��<���</�<#c�<ٕ�<)��<��<`%�<7R�<i}�<Ц�<r��<(��<�<�9�<]Y�<�v�<���<3��<(��<p��<���<x��< ��<`�<��<7�<h�<��<���<���<���<���<X��<���<�b�<�:�<��<t��<���<�l�<�,�<���<��<$N�<���<џ�<�@�<���<�r�<i�<���<��<ʙ�<��<E��<��<�q�<�۵<�A�< ��<, �<6Y�<>��<q��<�L�<ǖ�<Cݦ<b �<a`�<[��<|ן<��<�C�<1v�<\��<]Ԗ<F �<V*�<�R�<7y�<Q��<���<I�<q�<�%�<�D�<�b�<S��<t:}<sy<�u<d�q<@n<Pj<Ȇf<�b<��^<.[<$gW<��S<K�O<`L<OYH<&�D<&�@<�"=<|j9<N�5<32<MT.<�*<�'<>^#<C�<�$<=�<��<�s<��<Ao
<,�<��<� <�e�;`��;k��;b�;���;�Z�;K��;��;�Q�;6�;��;�;1��;U�;dC�;��;��;P�;LԊ;Jm�;��;��u;�ok;vKa;�PW;�~M;W�C;�U:;x�0;��';��;	�;�;7x;���:G�:��:���:���:q�:gq�:'�:T!r:�ZT:q�6:��:@v�92��9l��9q$9}Z8��W�J�!����ẹ�5﹕���J+���D��4^��_w��2����������|E��~��s�ź��Ѻ��ݺ��麦���9� �����������o�kK�#$���)���/���5�^b;�d+A���F�`�L�Y|R�@?X�)^��c���i��Bo�uu���z��@��!��U��-∻��r���c����i�� M���1���  �  �}=!=�=�f=g	=ϫ=�M=�� =�� =�2 =%��<���<�*�<Qk�<��<��<n(�<�e�<{��<:��< �<�R�<���<M��<���</�<c�<ҕ�<(��<���<l%�<$R�<G}�<���<Z��< ��<��<�9�<8Y�<�v�<���<!��<)��<a��<���<n��<��<e�<|�<A�<r�<��<���<���<���<Ǿ�<t��<���<�b�<�:�<��<}��<���<�l�<�,�<���<r��<6N�<���<ϟ�<�@�<r��<s�<E�<}��<��<���<��<*��<��<q�<�۵<�A�<���<% �<(Y�<H��<c��<�L�<Ŗ�<Dݦ<g �<j`�<p��<�ן<�<�C�<Sv�<p��<mԖ<g �<`*�<�R�<>y�<\��<���<U�<r�<}%�<�D�<�b�<W��<C:}<sy<�u<�q<n<�Oj<��f<۽b<x�^<�-[<gW<��S<�O<dL<7YH<0�D<%�@<�"=<�j9<>�5<E2<YT.<?�*<�'<{^#<u�<�$<��<	�<8t<��<no
<I�<��<� <ze�;���;C��;0b�;���;qZ�;K��;���;�Q�;��;���;��;���;9�;C�;���;#�;(P�;�ӊ;m�;��;)�u;�pk;2Ka;�PW;$M;*�C;�U:;��0;K�';�;b�;�; y;J��:NG�:���:���:L��:�:�q�:�&�:�!r:�[T:�6:(�:;r�9ӿ�9���9�b$9=�Z8+1X�=�!�)���㺹�:�ː��N+� �D�3^��cw�23��ꠔ������D���~����ź��Ѻ��ݺ ������� ����c��x���n��J��"$���)�I�/���5�%b;�+A���F��L�U|R�Z?X�� ^���c���i�DCo��u���z�vA��z!�����A∻HË�Ϥ��􆑻�i��M��2���  �  �}=!=�=�f=h	=ѫ=�M=�� =�� =�2 =4��<���<�*�<ck�<*��<$��<i(�<�e�<���<J��<�<�R�<���<O��<���</�<c�<ƕ�<��<���<Q%�<R�<C}�<���<J��<	��<��<�9�<:Y�<�v�<���<��<��<U��<���<v��<��<u�<��<O�<��<��<���<���<���<׾�<���<ȅ�<�b�<�:�<��<���<���<�l�<�,�<���<x��<*N�<}��<���<�@�<b��<�r�<B�<v��<��<���<��< ��<��<sq�<�۵<~A�<碲< �<Y�<C��<i��<�L�<ۖ�<Kݦ<x �<}`�<|��<�ן<�<�C�<dv�<���<mԖ<m �<r*�<�R�<Vy�<f��<<\�<p�<�%�<�D�<�b�<H��<7:}<�ry<��u<�q<n<�Oj<��f<��b<i�^<�-[<�fW<P�S<�O<HL<&YH<�D<+�@<�"=<�j9<n�5<W2<�T.<Z�*<�'<�^#<t�<!%<��<,�</t<��<�o
<l�<��<� <�e�;���;d��;2b�;���;EZ�;��;���;SQ�;��;~��;��;���;��;�B�;���;/�;�O�;�ӊ;�l�;u�;ؽu;pk;xKa;�PW;�M;��C;lV:;��0;��';��;x�;1;�y;?��:�G�:���:���:Ǯ�:���:�r�:�'�:$r:�[T:��6:��:>o�9���9U��9[[$9�`Z8�4X�Ԣ!�o��?麹�?�ԑ�GO+�H�D�!6^�ndw�4��ܡ��[���E��x~����źs�Ѻ �ݺ���Ǿ��!� ���������^n�@J��"$�j�)���/���5�ga;��*A�3�F�ȷL�f|R�0?X�A^���c��i�vCo�{u�J�z�xA���!������∻�Ë�줎������i���M��2���  �  �}=!=�=�f=l	=ͫ=�M=�� =�� = 3 =H��<���<+�<xk�<&��<F��<{(�<�e�<���<M��<�<�R�<���<E��<���<
/�<c�<ӕ�<��<���<8%�<R�</}�<���<?��<���<��<�9�<+Y�<qv�<���<��<��<k��<���<���<��<n�<��<M�<��<)��<��<���<
��<��<���<��<�b�<;�<��<���<���<�l�<�,�<���<���<N�<���<���<�@�<d��<�r�<3�<]��<|�<���<��<��<��<eq�<�۵<�A�<ߢ�< �<%Y�<.��<t��<�L�<ؖ�<Jݦ<z �<`�<���<�ן<�<D�<cv�<���<�Ԗ<y �<�*�<�R�<Yy�<_��<<S�<v�<�%�<�D�<�b�<?��<A:}<�ry<��u<��q<�n<�Oj<g�f<��b<2�^<�-[<�fW<4�S<�O<4L<NYH<�D<�@<�"=<�j9<{�5<I2<�T.<b�*<'<�^#<��<M%<��<q�<Ut<�<�o
<t�<ȃ<� <�e�;���;���;�a�;���;�Z�;���;���;�P�;��;3��;6�;q��;��;�B�;'��;���;^O�;�ӊ;�l�;n�;��u;�ok;�Ka;�PW;|M;��C;cV:;��0;��';k�;��;g;�y;���:�J�:F��:Y��:k��:���:�r�:)(�:�#r:�ZT:��6:�:yt�9���9�9]$9&Z8	QX��!�> ��*�rB�
���Q+���D��9^�{cw��4��0�������FF���}��/�ź��Ѻ �ݺ��麟����� ���������gn��I�o!$��)��/�w�5�Ma;��*A��F��L�5|R�,?X��^�*�c�U�i�KCo��u���z��A���!��+���∻�Ë�X���P���3j���M�� 2���  �  �}=!=�=�f=m	=ҫ=�M=�� =�� =3 =I��<���<+�<{k�<9��<?��<}(�<�e�<���<Y��<�<�R�<���<Q��<���</�<c�<���< ��<���<F%�<R�<)}�<���<<��<���<��<9�<)Y�<�v�<���<��<��<^��<���<{��<	��<s�<��<X�<��<0��<��<���<��<��<���<��<�b�<;�<��<���<���<�l�<�,�<���<���<N�<���<���<�@�<T��<�r�<3�<V��<y�<���<��<��<��<lq�<�۵<jA�<͢�<	 �<Y�</��<s��<�L�<ݖ�<Wݦ< �<�`�<���<�ן<�<D�<rv�<���<�Ԗ<u �<�*�<�R�<by�<n��<<]�<y�<~%�<�D�<�b�</��<:}<�ry<��u<��q<�n<�Oj<p�f<��b<1�^<�-[<�fW<;�S<��O<L<&YH<�D<�@<�"=<�j9<��5<h2<�T.<s�*<'<�^#<��<S%<ˏ<e�<Yt<�<�o
<��<҃<� <f�;���;���;�a�;���;0Z�;���;P��;/Q�;��;��;3�;g��;��;�B�;��;���;�O�;�ӊ;�l�;)�;&�u;�ok;�Ka;�PW;�M;0�C;�V:;��0;�';B�;��;0;z;2��:J�:W��: ��:���:J��:ks�:�(�:V$r:�[T:F�6:��:r�93��9���9bU$9BFZ8CNX���!�� ���캹�B�Z���R+���D��7^��fw��5��v�������.F���}��k�ź4�Ѻ1�ݺ���׽���� ���������m��I��!$�*�)��/�5�5�a;�}*A���F���L�|R�M?X��^���c�ڃi��Co��u�s�z��A��"��H���∻�Ë�[���X����i���M��]2���  �  �}=!=�=�f=j	=ϫ=�M=�� =�� =3 =S��<	��<+�<zk�<G��<9��<�(�<f�<���<a��<�<�R�<���<N��<���</�<c�<���<��<���<B%�<�Q�<}�<���<+��<���<��<�9�<Y�<zv�<{��< ��<��<O��<���<y��<��<m�<��<R�<��<2��<��<��<��<��<���<��<�b�<;�<��<���<���<�l�<�,�<���<}��<$N�<y��<���<�@�<R��<�r�<$�<S��<t�<���<��<��<{�<Wq�<�۵<gA�<좲<
 �<Y�<>��<m��<�L�<Җ�<Oݦ<x �<�`�<���<�ן<5�<�C�<�v�<���<�Ԗ<� �<�*�<�R�<_y�<l��<<Z�<u�<�%�<�D�<�b�<F��<2:}<�ry<��u<��q<�n<}Oj<[�f<t�b<7�^<-[<�fW<&�S<��O<GL<
YH<�D</�@<�"=<�j9<c�5<e2<�T.<}�*<'<�^#<��<Q%<�<X�<|t<,�<�o
<��<ƃ<� <�e�;���;���;8b�;���; Z�;4��;R��;"Q�;\�;���;F�;'��;u�;oB�;��;���;�O�;tӊ;m�;c�;��u;(pk;�Ka;�PW;uM;��C;�V:;��0;%�';��;��;T;lz;��:J�:a��:���:���:c��:&s�:(�:R#r:H[T:��6:E�:�n�9!��9���9cT$9�?Z8�lX���!�
"��z�*G�E��BT+���D�8^��fw��3��c���!���5E��~����ź��Ѻ��ݺ���g����� �m��M��E��rm�pI�O!$�B�)���/��5�a;��*A�N�F�ڷL�<|R�?X�4^�/�c�!�i��Co�u���z�B���!��r��㈻ċ�M�������Gj���M��92���  �  �}=!=�=�f=m	=ҫ=�M=�� =�� =3 =I��<���<+�<{k�<9��<?��<}(�<�e�<���<Y��<�<�R�<���<Q��<���</�<c�<���< ��<���<F%�<R�<)}�<���<<��<���<��<9�<)Y�<�v�<���<��<��<^��<���<{��<	��<s�<��<X�<��<0��<��<���<��<��<���<��<�b�<;�<��<���<���<�l�<�,�<���<���<N�<���<���<�@�<T��<�r�<3�<V��<y�<���<��<��<��<lq�<�۵<jA�<͢�<	 �<Y�</��<s��<�L�<ݖ�<Wݦ< �<�`�<���<�ן<�<D�<rv�<���<�Ԗ<u �<�*�<�R�<by�<n��<<]�<y�<~%�<�D�<�b�</��<:}<�ry<��u<��q<�n<�Oj<p�f<��b<1�^<�-[<�fW<;�S<��O<L<&YH<�D<�@<�"=<�j9<��5<h2<�T.<s�*<'<�^#<��<S%<ˏ<e�<Yt<�<�o
<��<҃<� <f�;���;���;�a�;���;0Z�;���;P��;/Q�;��;��;3�;g��;��;�B�;��;���;�O�;�ӊ;�l�;)�;&�u;�ok;�Ka;�PW;�M;0�C;�V:;��0;�';B�;��;0;z;2��:J�:W��: ��:���:J��:ks�:�(�:V$r:�[T:F�6:��:r�93��9���9bU$9BFZ8CNX���!�� ���캹�B�Z���R+���D��7^��fw��5��v�������.F���}��k�ź4�Ѻ1�ݺ���׽���� ���������m��I��!$�*�)��/�5�5�a;�}*A���F���L�|R�M?X��^���c�ڃi��Co��u�s�z��A��"��H���∻�Ë�[���X����i���M��]2���  �  �}=!=�=�f=l	=ͫ=�M=�� =�� = 3 =H��<���<+�<xk�<&��<F��<{(�<�e�<���<M��<�<�R�<���<E��<���<
/�<c�<ӕ�<��<���<8%�<R�</}�<���<?��<���<��<�9�<+Y�<qv�<���<��<��<k��<���<���<��<n�<��<M�<��<)��<��<���<
��<��<���<��<�b�<;�<��<���<���<�l�<�,�<���<���<N�<���<���<�@�<d��<�r�<3�<]��<|�<���<��<��<��<eq�<�۵<�A�<ߢ�< �<%Y�<.��<t��<�L�<ؖ�<Jݦ<z �<`�<���<�ן<�<D�<cv�<���<�Ԗ<y �<�*�<�R�<Yy�<_��<<S�<v�<�%�<�D�<�b�<?��<A:}<�ry<��u<��q<�n<�Oj<g�f<��b<2�^<�-[<�fW<4�S<�O<4L<NYH<�D<�@<�"=<�j9<{�5<I2<�T.<b�*<'<�^#<��<M%<��<q�<Ut<�<�o
<t�<ȃ<� <�e�;���;���;�a�;���;�Z�;���;���;�P�;��;3��;6�;q��;��;�B�;'��;���;^O�;�ӊ;�l�;n�;��u;�ok;�Ka;�PW;|M;��C;cV:;��0;��';k�;��;g;�y;���:�J�:F��:Y��:k��:���:�r�:)(�:�#r:�ZT:��6:�:yt�9���9�9]$9&Z8	QX��!�> ��*�rB�
���Q+���D��9^�{cw��4��0�������FF���}��/�ź��Ѻ �ݺ��麟����� ���������gn��I�o!$��)��/�w�5�Ma;��*A��F��L�5|R�,?X��^�*�c�U�i�KCo��u���z��A���!��+���∻�Ë�X���P���3j���M�� 2���  �  �}=!=�=�f=h	=ѫ=�M=�� =�� =�2 =4��<���<�*�<ck�<*��<$��<i(�<�e�<���<J��<�<�R�<���<O��<���</�<c�<ƕ�<��<���<Q%�<R�<C}�<���<J��<	��<��<�9�<:Y�<�v�<���<��<��<U��<���<v��<��<u�<��<O�<��<��<���<���<���<׾�<���<ȅ�<�b�<�:�<��<���<���<�l�<�,�<���<x��<*N�<}��<���<�@�<b��<�r�<B�<v��<��<���<��< ��<��<sq�<�۵<~A�<碲< �<Y�<C��<i��<�L�<ۖ�<Kݦ<x �<}`�<|��<�ן<�<�C�<dv�<���<mԖ<m �<r*�<�R�<Vy�<f��<<\�<p�<�%�<�D�<�b�<H��<7:}<�ry<��u<�q<n<�Oj<��f<��b<i�^<�-[<�fW<P�S<�O<HL<&YH<�D<+�@<�"=<�j9<n�5<W2<�T.<Z�*<�'<�^#<t�<!%<��<,�</t<��<�o
<l�<��<� <�e�;���;d��;2b�;���;EZ�;��;���;SQ�;��;~��;��;���;��;�B�;���;/�;�O�;�ӊ;�l�;u�;ؽu;pk;xKa;�PW;�M;��C;lV:;��0;��';��;x�;1;�y;?��:�G�:���:���:Ǯ�:���:�r�:�'�:$r:�[T:��6:��:>o�9���9U��9[[$9�`Z8�4X�Ԣ!�o��?麹�?�ԑ�GO+�H�D�!6^�ndw�4��ܡ��[���E��x~����źs�Ѻ �ݺ���Ǿ��!� ���������^n�@J��"$�j�)���/���5�ga;��*A�3�F�ȷL�f|R�0?X�A^���c��i�vCo�{u�J�z�xA���!������∻�Ë�줎������i���M��2���  �  �}=!=�=�f=g	=ϫ=�M=�� =�� =�2 =%��<���<�*�<Qk�<��<��<n(�<�e�<{��<:��< �<�R�<���<M��<���</�<c�<ҕ�<(��<���<l%�<$R�<G}�<���<Z��< ��<��<�9�<8Y�<�v�<���<!��<)��<a��<���<n��<��<e�<|�<A�<r�<��<���<���<���<Ǿ�<t��<���<�b�<�:�<��<}��<���<�l�<�,�<���<r��<6N�<���<ϟ�<�@�<r��<s�<E�<}��<��<���<��<*��<��<q�<�۵<�A�<���<% �<(Y�<H��<c��<�L�<Ŗ�<Dݦ<g �<j`�<p��<�ן<�<�C�<Sv�<p��<mԖ<g �<`*�<�R�<>y�<\��<���<U�<r�<}%�<�D�<�b�<W��<C:}<sy<�u<�q<n<�Oj<��f<۽b<x�^<�-[<gW<��S<�O<dL<7YH<0�D<%�@<�"=<�j9<>�5<E2<YT.<?�*<�'<{^#<u�<�$<��<	�<8t<��<no
<I�<��<� <ze�;���;C��;0b�;���;qZ�;K��;���;�Q�;��;���;��;���;9�;C�;���;#�;(P�;�ӊ;m�;��;)�u;�pk;2Ka;�PW;$M;*�C;�U:;��0;K�';�;b�;�; y;J��:NG�:���:���:L��:�:�q�:�&�:�!r:�[T:�6:(�:;r�9ӿ�9���9�b$9=�Z8+1X�=�!�)���㺹�:�ː��N+� �D�3^��cw�23��ꠔ������D���~����ź��Ѻ��ݺ ������� ����c��x���n��J��"$���)�I�/���5�%b;�+A���F��L�U|R�Z?X�� ^���c���i�DCo��u���z�vA��z!�����A∻HË�Ϥ��􆑻�i��M��2���  �  �}=!=	�=�f=i	=ɫ=�M=�� =�� =�2 =��<���<�*�<Bk�<���<��<G(�<�e�<f��<,��<��<�R�<���<?��<���</�<#c�<ٕ�<)��<��<`%�<7R�<i}�<Ц�<r��<(��<�<�9�<]Y�<�v�<���<3��<(��<p��<���<x��< ��<`�<��<7�<h�<��<���<���<���<���<X��<���<�b�<�:�<��<t��<���<�l�<�,�<���<��<$N�<���<џ�<�@�<���<�r�<i�<���<��<ʙ�<��<E��<��<�q�<�۵<�A�< ��<, �<6Y�<>��<q��<�L�<ǖ�<Cݦ<b �<a`�<[��<|ן<��<�C�<1v�<\��<]Ԗ<F �<V*�<�R�<7y�<Q��<���<I�<q�<�%�<�D�<�b�<S��<t:}<sy<�u<d�q<@n<Pj<Ȇf<�b<��^<.[<$gW<��S<K�O<`L<OYH<&�D<&�@<�"=<|j9<N�5<32<MT.<�*<�'<>^#<C�<�$<=�<��<�s<��<Ao
<,�<��<� <�e�;`��;k��;b�;���;�Z�;K��;��;�Q�;6�;��;�;1��;U�;dC�;��;��;P�;LԊ;Jm�;��;��u;�ok;vKa;�PW;�~M;W�C;�U:;x�0;��';��;	�;�;7x;���:G�:��:���:���:q�:gq�:'�:T!r:�ZT:q�6:��:@v�92��9l��9q$9}Z8��W�J�!����ẹ�5﹕���J+���D��4^��_w��2����������|E��~��s�ź��Ѻ��ݺ��麦���9� �����������o�kK�#$���)���/���5�^b;�d+A���F�`�L�Y|R�@?X�)^��c���i��Bo�uu���z��@��!��U��-∻��r���c����i�� M���1���  �  �}=!=�=�f=h	=ƫ=�M=�� =�� =�2 =
��<���<�*�<5k�<��<���<%(�<�e�<R��<��<��<�R�<���<5��<���</�<*c�<��<,��<*��<s%�<UR�<l}�<ަ�<���<C��<�<�9�<rY�<�v�<đ�<:��<,��<���<���<���<���<d�<u�<�<m�<���<���<���<���<���<E��<���<pb�<�:�<q�<w��<l��<�l�<�,�<���<���<#N�<���<֟�<�@�<���<s�<��<���<��<晽<�<Z��<��<�q�<�۵<�A�<��<7 �<AY�<>��<y��<�L�<ϖ�<)ݦ<Q �<Z`�<D��<zן<��<�C�<v�<P��<;Ԗ<2 �<L*�<�R�<7y�<4��<���<G�<l�<�%�<�D�<�b�<W��<�:}<?sy<�u<��q<En<IPj<��f<H�b<��^<..[<`gW<��S<e�O<gL<wYH</�D<1�@<�"=<qj9<K�5<�2<HT.<�*<�'<!^#<��<�$<�<��<�s<��<o
<�<i�<t <�e�;1��;v��;b�;	��;�Z�;N��;R��;�Q�;��;��;L�;���;��;�C�;���;�;RP�;�Ԋ;am�;��;%�u;�ok;�Ka;FPW;M;��C;�T:;��0;��';s�;7�;�;�w;B��:GE�:B��:���:���:��:�o�:�%�:"r:�XT:��6:f�:Az�9���9���9 y$9R�Z8߽W�N�!���vں�./�B���J+�[�D�-2^��]w��2�����*����E���}��"�źb�ѺU�ݺ���&����� �������;���p��K�$$�J�)���/���5�_b;�O,A���F�p�L�~|R��>X�^��c���i�Bo��u���z��@��!��� ���ሻr�W���*���i���L��`1���  �  �}=!=�=�f=f	=ë=�M=�� =|� =�2 =��<���<�*�<k�<Ū�<���<%(�<�e�<;��<��<��<�R�<���<4��<���</�<*c�<��<I��<)��<�%�<]R�<�}�< ��<���<W��<4�<�9�<tY�<�v�<ɑ�<N��<E��<|��<���<|��<���<X�<m�<�<[�<���<���<���<���<���<+��<���<ub�<�:�<_�<g��<j��<�l�<�,�<���<���<1N�<���<��<�@�<���<-s�<��<���<��<���<'�<{��<��<�q�<�۵<�A�<��<D �<AY�<H��<o��<�L�<���<&ݦ<I �<K`�<0��<gן<��<�C�<v�<4��</Ԗ<- �<.*�<oR�<(y�<1��<���<A�<l�<�%�<�D�<�b�<u��<�:}<asy<?�u<��q<�n<jPj<(�f<d�b<��^<D.[<}gW<ءS<m�O<�L<wYH<>�D<2�@<~"=<gj9<$�5<�2<.T.<��*<D'<^#<�<�$<ڎ<��<�s<e�<�n
<��<N�<h <Ae�;(��;J��;b�;��;�Z�;���;H��;DR�;��;b��;��;���;�;"D�;u��;�;�P�;�Ԋ;�m�;�;�u;&pk;�Ka;TPW;�~M;��C;�T:;�0;��';��;;�;$;�v;���:�C�:x��:��:���:��:�o�:�%�:$ r:7YT:��6:��:�x�9���9.��9Ly$9b�Z8I�W���!�E��Vպ�+�]���G+���D�H.^��]w�1��H���E���E��k~���ź��Ѻ��ݺ4������� �H�������nq��L�|$$�v�)���/�&�5��b;�d,A�W�F���L��|R�?X�� ^���c���i��Ao�ou�H�z��@��� ��� ��oሻ:�ˣ�������h���L��Q1���  �  ~=!=�=�f=g	=ī=�M=�� =m� =�2 =��<���<�*�< k�<���<���<
(�<�e�<;��<��<��<�R�<w��<A��<���</�<4c�<��<T��<1��<�%�<gR�<�}�<��<���<x��<6�<:�<�Y�<�v�<ӑ�<U��<F��<{��<���<o��<��<J�<j�<�<;�<���<���<���<���<r��<��<r��<Ub�<�:�<m�<I��<]��<�l�<�,�<���<x��<?N�<���<��<�@�<���<Is�<��<��<��<��<A�<���<�<�q�<ܵ<�A�<+��<? �<IY�<O��<i��<�L�<���<*ݦ<7 �<:`�<6��<Bן<��<�C�<�u�<��<Ԗ< �<*�<yR�<	y�<1��<���<;�<p�<z%�<�D�<�b�<{��<�:}<sy<i�u<��q<�n<|Pj<p�f<�b<4�^<�.[<�gW<��S<y�O<�L<gYH<X�D<'�@<�"=<kj9<�5<�2<�S.<ɨ*<1'<�]#<��<Q$<͎<d�<es<�<�n
<��<�<m <e�;V��;/��;b�;%��;�Z�;���;a��;�R�;��;���;��;��;��;&D�;!��;S�;
Q�;�Ԋ;�m�;�;۾u;�pk;Ka;�PW;3~M;y�C;pT:;��0;V�';��;-�;X;8v;���:CB�:l��: ��:`��:��:�n�:�%�:#r:�[T:
�6:}�:y�9���9���9�}$9j[8�W�;m!�c���ͺ�/%�p���B+�x�D��+^��\w�e0�����������D���~���ź}�Ѻo�ݺb��D���s� �t�����ۑ��q�qM�N%$���)�a�/�ԗ5��c;�e,A���F�ʸL�b|R�k?X�` ^���c�z�i��Ao�� u���z�@�����| �������\��������h��<L��91���  �  ~=$!=�=�f=h	=��=�M=�� =j� =�2 =ԧ�<���<�*�<�j�<���<���<(�<�e�<%��<���<��<�R�<l��<3��<���</�<>c�<���<^��<G��<�%�<yR�<�}�<��<���<���<F�<:�<�Y�<�v�<��<f��<O��<���<���<u��<��<>�<Z�<�<5�<���<���<���<���<_��<��<j��<Pb�<�:�<T�<>��<S��<yl�<�,�<���<���<?N�<���<���< A�<���<Ss�<��<��<�<-��<R�<���<�<�q�<ܵ<�A�<:��<T �<YY�<N��<r��<�L�<���<ݦ<1 �<#`�<��<Dן<��<�C�<�u�<��<Ԗ< �<*�<]R�<y�<"��<���<.�<p�<�%�<�D�<�b�<���<�:}<�sy<��u<��q<�n<�Pj<��f<��b<1�^<�.[<�gW<�S<��O<�L<�YH<_�D<*�@<�"=<Oj9<��5<�2<�S.<��*<'<�]#<��<2$<��<L�<Zs<�<�n
<��<�<J <�d�;��;D��;b�;G��;�Z�;��;���;�R�;%�;���;��;W��;��;aD�;��;{�;7Q�;Պ;n�;7�;��u;�pk;DKa;�PW;�}M;��C;T:;��0;��';m�;�;;�u;m��:�A�:��:���:Ĩ�:��:5n�:�$�:�r:^ZT:��6:S�:�}�9���9��9�$9�![8C}W�m!�p��!ʺ�*!ﹺ��B+�,�D��*^�Zw��/��y��� ����D��e~���ź%�Ѻw�ݺ��麵���:� �i�����0��br��M��%$���)���/���5��c;��,A���F�0�L�a|R�>?X�M ^��c�;�i��@o�| u�=�z��?�� ��8 ����������e���p���ch��L���0���  �  ~='!=�=�f=d	=��=�M=�� =n� =�2 =���<l��<q*�<�j�<���<���<�'�<re�<��<���<��<�R�<���<&��<���< /�<5c�<��<X��<J��<�%�<�R�<�}�<2��<���<���<n�<:�<�Y�<�v�<��<g��<Q��<���<���<���<���<L�<b�< �<<�<���<���<y��<m��<S��<���<S��<9b�<�:�<7�<D��<M��<|l�<�,�<���<���<8N�<���<���<A�<���<_s�<��<���<,�<2��<`�<���<#�<�q�<)ܵ<�A�<8��<\ �<RY�<P��<{��<�L�<���<ݦ<2 �<#`�<��<5ן<��<oC�<�u�<��<�Ӗ<���< *�<GR�<y�<��<���<2�<b�<�%�<�D�<�b�<��<�:}<�sy<��u<�q<�n<�Pj<��f<Ӿb<f�^<�.[<�gW< �S<��O<�L<�YH<O�D<>�@<t"=<Jj9<$�5<�2<�S.<l�*<� '<�]#<q�<$<u�<&�<!s<��<�n
<��<�<9 <&e�;ݩ�;K��;b�;��;[�;���;���;�R�;��;��;��;���;��;�D�;8��;��;dQ�;Պ;n�;;�;i�u;6pk;�Ka;�OW;8~M;2�C;�S:;��0;��';�;k�;P;:u;}��::@�:���:ٜ�:ᦶ:�:�m�:�$�:r:�WT:|�6:`�:}�9���9���9$�$9�6[8�FW��i!�g���ɺ�3�
��&A+���D�z)^��Yw��/�����|����D���}���ź��Ѻ��ݺ�������� �������֒��r�MN�g&$�G�)�S�/�e�5��c;�*-A�q�F��L��|R��>X�� ^���c�Z�i��@o�g u�¿z��?�������������_�������*���h���K���0���  �  ~=)!=�=�f=c	=��=�M=�� =b� =�2 =Χ�<i��<p*�<�j�<���<���<�'�<qe�< ��<���<��<�R�<q��<)��<���<"/�<>c�<��<g��<T��<�%�<�R�<�}�<.��<���<���<b�<:�<�Y�<�v�<���<n��<]��<���<���<���<���<F�<O�<��<$�<���<���<p��<k��<T��<���<Q��<3b�<�:�<H�<2��<=��<jl�<�,�<���<���<@N�<���<
��<	A�<���<cs�<��<���<$�<=��<g�<���<"�<�q�<1ܵ<�A�<E��<b �<YY�<T��<v��<�L�<���<ݦ<  �<`�<��<3ן<��<kC�<�u�<���<�Ӗ<���<*�<SR�<�x�<	��<���</�<c�<�%�<�D�<c�<���<�:}<�sy<��u<�q<�n<�Pj<��f<վb<h�^<�.[<�gW<4�S<��O<�L<�YH<b�D<B�@<r"=<Jj9<��5<�2<�S.<y�*<'<�]#<o�<	$<�<�<s<��<�n
<��<�< <�d�;��;6��;!b�;>��; [�;!��;��;�R�;v�;��;u�;���;��;�D�;<��;��;hQ�;<Պ;n�;l�;��u;�pk;�Ka;�OW;~M;��C;@S:;8�0;�';:�;#�;5;@u;���:@�:6��:��:槶:��:�l�:#�:�r:<XT:Y�6:V�:�~�9K��9޺�9��$9R>[8�KW��i!������ƺ�~���CA+�D�D�{(^��Xw��.����������D��@~����ź��Ѻ��ݺ���L���� �����������r�oN�l&$�s�)���/��5��d;��-A��F�)�L��|R��>X�= ^���c��i��@o� u���z��?���������Y���[�������0���h���K���0���  �  �={#=��=�i=�=��=!R=t� =|� =G8 =���<(��<8�<ky�<'��<(��<�9�<x�<ҵ�<���<�.�<�i�<��<���<��<|K�<��<��<���<(�<I�<dw�<'��<+��<[��<��<=E�<�h�<��<��<���<��<���<��<�<Z.�<�:�<�C�<�I�<&L�<K�<IF�<�=�<z1�<!�<t�<���<v��<���<Q��<=c�<H3�<k��<c��<<��<�@�<B��<U��<�S�<H��<��<�6�<���<y]�<��<Do�<X�<[l�<c�<�U�<�·<[+�<N��<��<J�<��<��<�B�<5��<�ը<��<�Z�<��<�ҡ<U
�<Z?�<�q�<���<\Ϙ<���<�$�<L�<r�<E��<��<Fڋ<T��<*�<�6�<�S�<�o�<Ί�<�J}<�~y<�u<��q<�n<�Hj<�zf<h�b<��^<�[<mHW<�}S<��O<:�K<0'H<<cD<4�@<��<<�$9<pj5<r�1<��-<LO*<Ϣ&<��"<�V<O�< <ć<0�<#n<5�	<�l<��<�
�;�8�;au�;J��;4�;���;��;ؕ�;�6�;X��;�;^��;�y�;�{�;D��;���;��;pX�;�Ŏ;H�;^��;�};��r;Yh;#7^;�@T;tJ;`�@;{X7;=.;E�$;5�;�;sK
;|�;ϖ�:���:,��:c��:}��:%�:�Ē:*��:JIi:E�K:�.:��:f��9I��9gv9�9i��7�Р�( ;��Y����ƹ����R
�C�0�	�I�c��|�t���˖����D��?i���}Ǻ�Ӻ'ߺ�k��M�����w�X�v4�������$� {*��D0��
6���;���A�PG��M�z�R���X��@^�o�c�ߴi�oo�.(u�x�z��M��D*�����刻�Ë�㡎�p���_a��=B��9$���  �  �=z#=��=�i=�=��=+R=o� =|� =K8 =���<,��<8�<{y�<-��<8��<�9�<x�<��<���<�.�<�i�<���<���<��<wK�<��<��<���<;�<I�<cw�<��<��<`��<��<5E�<�h�<��<��<���<��<���<��<�<d.�<�:�<�C�<�I�<L�<K�<YF�<�=�<s1�<
!�<��<���<y��<���<j��<Pc�<U3�<b��<p��<Q��<�@�<K��<N��<�S�<@��<&��<�6�<���<}]�<���<=o�<a�<_l�<W�<mU�<�·<V+�<[��<��<J�<��<��<�B�<-��<�ը<��<�Z�<(��<�ҡ<f
�<Y?�<�q�<���<oϘ<���<�$�<,L�<r�<H��< ��<[ڋ<Y��<%�<�6�<�S�<�o�<Ǌ�<�J}<�~y<ڱu<m�q<�n<�Hj<{f<j�b<D�^<�[<]HW<�}S<ݴO<-�K<-'H<'cD<7�@<��<<�$9<�j5<^�1<��-<ZO*<��&<��"<�V<p�<<�<,�<?n<`�	<�l<��<�
�;�8�;Fu�;M��;"�;���;��;ݕ�;�6�;Q��;鰽;��;Sy�;|�;t��;���;>�;rX�;eŎ;H�;���;�};{�r;�Xh;v7^;�@T;�tJ;��@;;X7;�.;��$;�;q;WK
;�;���:���:���:���:���:�%�:^Ē:���:�Ki:��K:>�.:��:E��9���9v9�9W��7�̠�t;��[��Q�ƹ�������0���I��c�|� t���˖����E��i��T~ǺN�Ӻ�~ߺIl�8M��f��Bw�X��3������$�={*�5D0��
6�}�;��A�lOG��M���R�W�X�7A^�w�c��i�~no�5(u���z��M���*����|刻�Ë�f��������a��FB���#���  �  �=~#=��=�i=�=��=)R=o� =�� =L8 =���<5��<#8�<�y�<.��<I��<�9�<#x�<��<���<�.�<�i�<���<���<��<|K�<��<��<���<.�< I�<fw�<��<��<R��<��<3E�<�h�<���<���<���<��<���<��<
�<q.�<�:�<�C�<�I�<!L�<!K�<TF�<�=�<v1�<!�<��<���<���<´�<s��<Kc�<h3�<i��<m��<J��<�@�<X��<M��<�S�<9��<��<�6�<���<�]�<���<;o�<I�<Kl�<W�<lU�<�·<C+�<O��<��<J�<��<��<C�< ��<�ը<��<�Z�<7��<�ҡ<k
�<X?�<�q�<���<|Ϙ<���<�$�<6L�<r�<^��< ��<Zڋ<P��<*�<�6�<�S�<�o�<���<�J}<�~y<ӱu<��q<�n<�Hj<�zf<Y�b<>�^<�[<[HW<�}S<ŴO<
�K<:'H<cD<K�@<��<<�$9<�j5<^�1<��-<bO*<
�&<��"<�V<��<<	�<,�<On<d�	<�l<��<�
�;�8�;(u�;���;9�;���;��;���;�6�;��;���;%��;Vy�;�{�;��;���;*�;�X�;7Ŏ;�G�;k��;0};��r;�Xh;�7^;�@T;ZtJ;��@;UX7;(.;��$;d�;�;�K
;8�;��:� �:;��:���:`��:	'�:�Ē:ܚ�:/Ki:9�K:�.:��:g��9��9�v9i9IC�7u���;��[���ƹ[������0���I��c�}|�#u���˖�����D���g��Ǻ��Ӻ�~ߺlk�@L��x��w� X�w3������ݮ$�{*��C0��
6���;��A�wOG��M�z�R���X�jA^�P�c���i��no��(u���z��M���*��'���刻�Ë�q���j����a���B��#$���  �  �=u#=��=�i=�=��=*R=w� =�� =S8 =���<N��<<8�<�y�<B��<Q��<�9�<<x�<���<���<�.�<�i�<���<���<��<qK�<ހ�< ��<���< �<�H�<Iw�<���<��<F��<��<E�<�h�<Ӊ�<��<���<���<���<��<�<_.�<�:�<�C�<�I�<-L�< K�<gF�<�=�<�1�<+!�<��<���<���<ߴ�<���<^c�<h3�<u��<u��<R��<�@�<D��<E��<�S�<4��<��<�6�<���<^]�<���<"o�<;�<?l�<=�<RU�<�·<;+�<A��<��<J�<��<��<�B�<8��<�ը<��<�Z�<=��<�ҡ<�
�<t?�<�q�<ϡ�<�Ϙ<��<�$�<AL�<r�<[��<��<\ڋ<`��<3�<�6�<�S�<�o�<���<uJ}<�~y<��u<@�q<�n<�Hj<�zf<:�b<�^<�[</HW<�}S<��O<�K<'H<cD<0�@<��<<�$9<�j5<�1<��-<~O*<"�&<��"<�V<��<:<�<g�<�n<��	<�l<��<�;�8�;�u�;f��;�;[��;��;���;x6�;���;���;���;�x�;�{�;蒥;J��;� �;X�;Ŏ;�G�;8��;7};%�r;�Xh;W7^;(AT;�tJ;�@;�X7;!.;B�$;��;�;mL
;��;ݘ�:��:��:���:���:'�:�Œ:k��:bLi:�K:��.:��:���9���9d	v9`9m#�7w頸&;��a��X�ƹ�����&�0��I��c�|�cu��|̖�����E���h��~}Ǻ��Ӻ5~ߺ�j��K����Wv�=W�!3��c���$�%z*��C0�
6���;���A�eOG�qM�6�R�~�X��A^���c���i�boo��(u�~�z�4N��3+��k��戻ċ����������a���B��g$���  �  �=l#=��=�i=�=��=.R=�� =�� =a8 =г�<T��<K8�<�y�<g��<e��<�9�<Bx�<��<���<�.�<j�<���<���<��<�K�<��<���<���<�<�H�<8w�<��<���<)��<��<�D�<}h�<�<��<���<���<���<��<�<[.�<�:�<�C�<�I�<AL�<)K�<�F�<�=�<�1�<8!�<��<���<���<��<���<|c�<p3�<���<���<N��<�@�<;��<Z��<�S�<.��<���<r6�<���<L]�<���<�n�<#�<"l�<�<HU�<�·<0+�<'��<��<�I�< ��<��<�B�<;��<�ը<��<�Z�<J��<�ҡ<�
�<�?�<�q�<���<�Ϙ<"��<�$�<PL�<=r�<b��<(��<fڋ<`��<$�<�6�<�S�<xo�<���<MJ}<`~y<��u<�q<Yn<bHj<�zf<��b<��^<�[<HW<�}S<x�O<�K<�&H<1cD<=�@<��<<�$9<�j5<��1<��-<�O*<E�&<��"<W<ط<�<E�<��<�n<��	<m<��<��;�8�;�u�;.��;[�;~��;��;���;!6�;���;L��;���;�x�;6{�;���;ʾ�;� �;�W�;�Ď;�G�;��;"};��r;bYh;>7^;AT;�tJ;��@;dY7;q.;X�$;%�;�;�L
;��;B��:��:���:���:�ñ:�'�:�ƒ:m��:Li:)�K:��.:��:Z��9���9�v9�
9���7 ����;�;j����ƹ������%�0��I��c�|��u���̖����ED���i��:}Ǻ��Ӻ�|ߺIj��J��)��v��V��2��	�|����$�z*�C0�	6���;�ݎA�OG�pM���R�m�X��@^�b�c���i�po�P)u���z�{N���+�����Q戻�ċ����:���b���B���$���  �  �=k#=��=�i=�=��=4R=�� =�� =g8 =��<z��<i8�<�y�<s��<���<�9�<dx�< ��<��<�.�<j�<	��<��<��<xK�<р�<��<���<��<�H�<w�<գ�<���<
��<q�<�D�<\h�<���<Ũ�<���<���<���<��<
�<b.�<�:�<�C�<�I�<IL�<@K�<�F�<>�<�1�<Z!�<��<���<���<��<���<�c�<�3�<���<���<X��<�@�<E��<J��<�S�<��<��<a6�<t��<;]�<���<�n�<��<�k�<�<&U�<p·<+�<��<��<�I�<<��<�B�<A��<�ը<��<�Z�<\��<�ҡ<�
�<�?�<r�<���<�Ϙ<A��<�$�<oL�<Fr�<{��<+��<pڋ<o��<4�<�6�<�S�<to�<���<3J}<6~y<X�u<�q<*n<7Hj<Szf<Ǭb<��^<e[<�GW<�}S<b�O<��K<�&H<cD<5�@<��<<�$9<�j5<��1<��-<�O*<��&<A�"<KW<�<�<��<��<�n<��	</m<�<��;-9�;�u�;���;=�;4��;|�;=��;�5�;~��;;-��;Rx�;�z�;��;���;I �;�W�;yĎ;EG�;�߃;�};��r;�Xh;�7^;XAT; uJ;��@;�Y7;4	.;��$;<�;�;�M
;D�;:��:�:��:A��:&ı:)�:&ǒ:ݜ�:�Mi:��K:4�.:��:���9���9��u9�9��79��M1;��n���ƹ�����
�0���I�,c��|��v��g͖�����D���h���|Ǻ؃Ӻk|ߺVi��I�����u��U��1�z	������$��x*�B0��6���;���A��NG��M�*�R�j�X��A^���c�:�i�hpo��)u���z��N���+��D	���戻�ċ�n��������b��&C���$���  �  �=k#=��=�i=�=��==R=�� =�� =t8 = ��<���<�8�<�y�<���<���<�9�<�x�<4��< ��</�<j�<��<��<��<lK�<΀�<��<���<��<�H�<w�<���<���<���<V�<�D�<5h�<���<���<��<���<���<��<��<`.�<�:�<�C�<�I�<SL�<`K�<�F�<7>�<�1�<y!�<��<��<���<��<ǎ�<�c�<�3�<���<���<g��<�@�<B��<9��<�S�<
��<Ԛ�<S6�<X��<"]�<���<�n�<��<�k�<��<�T�<Z·<�*�<��<��<�I�<�<��<�B�<:��<�ը<�<�Z�<x��<ӡ<�
�<�?�<4r�<!��<�Ϙ<]��<�$�<�L�<]r�<���<4��<�ڋ<n��</�<�6�<�S�<wo�<���<J}<~y<&�u<��q<�n<Hj<zf<��b<p�^< [<�GW<Y}S<L�O<��K<�&H<�bD<)�@<��<<�$9<�j5<ȳ1<. .<P*<��&<g�"<}W<\�<�<ۈ<��<o<	�	<hm<:�<��;�9�;�u�;y��;�;4��;e�;ޔ�;�5�;&��;���;���;�w�;xz�;���;Q��;���;OW�;Ď;G�;�߃; };ۤr;�Xh;{7^;6AT;nuJ;;�@;Z7;>
.;E�$;
�;|;�N
;>�;H��:>�:��:��:�ű:+�:Ȓ:���:Oi:m�K:��.:�:	��9��9�u9��9!�7���D;��r����ƹ������0�r�I�r c�v|��x��HΖ�����E���h��
}Ǻ��Ӻ�{ߺh��G����t�@U�d0�g����ī$�Mx*�wA0�6���;�}�A�<NG�
M�Y�R���X��A^�g�c���i��po�*u���z�,O���,���	��t爻4ŋ����
����b��rC��%���  �  �=c#=��=�i=�=��==R=�� =�� =~8 =��<���<�8�<�y�<���<���<:�<�x�<M��</��<!/�<)j�<��<��<��<rK�<π�<ش�<���<��<�H�<�v�<���<���<���<3�<�D�<%h�<~��<���<_��<���<���<��<��<d.�<�:�<�C�<�I�<mL�<gK�<�F�<K>�<�1�<�!�<�<2��<���<>��<ێ�<�c�<�3�<���<���<a��<A�<B��<;��<�S�<���<Ú�<16�<@��<]�<u��<�n�<��<�k�<��<�T�<?·<�*�<쎴<��<�I�<堯<��<�B�<G��<�ը<�<�Z�<���<ӡ<�
�<�?�<Dr�<=��<�Ϙ<~��<%�<�L�<ur�<���<O��<�ڋ<q��<9�<�6�<�S�<fo�<���<�I}<�}y<��u<��q<�n<�Gj<�yf<b�b<A�^<�[<�GW<#}S<�O<��K<�&H<�bD<3�@<��<<�$9<�j5<��1<B .<-P*<У&<��"<�W<~�< <��<G�<Xo<>�	<�m<W�<$�;v9�;v�;���;9�;?��;,�;Ô�;w5�;���;a��;m��;rw�;�y�;4��;½�;}��;�V�;�Î;�F�;B߃;�};7�r;�Xh;�7^;�AT;puJ;��@;�Z7;{
.;'�$;��;�;�O
;�;���:Y�:V��:o��:.Ǳ:�+�:�ɒ:���:Oi:R�K:E�.:{�:P��9���9��u9��9���7�<��8K;�\{���ƹ׿������0�j�I�U#c��|�7y��1ϖ�����E���h��|Ǻ�Ӻ�zߺg�!G��?��?s��S��/�������$�8w*��@0�Y6���;���A�NG��M��R�a�X��A^���c�@�i��qo�O+u�5�z��O���,��
���爻�ŋ�b���]���-c���C��z%���  �  �=\#=��=�i=�=��=?R=�� =�� =�8 =/��<���<�8�<z�<ٺ�<���<&:�<�x�<i��<D��<./�<>j�<��<$��<��<cK�<���<д�<���<��<�H�<�v�<|��<x��<���<(�<�D�<h�<[��<���<L��<���<���<��<��<R.�<�:�<�C�<�I�<�L�<tK�<�F�<`>�<2�<�!�<"�<R��<��<`��<��<�c�<�3�<���<���<i��<A�<3��<4��<�S�<���<���<6�<4��<�\�<P��<�n�<��<�k�<��<�T�<·<�*�<Ҏ�<�<�I�<Ԡ�<��<�B�<W��<�ը<$�<�Z�<���<8ӡ<�
�<�?�<Tr�<`��<И<���<%�<�L�<�r�<���<e��<�ڋ<���<B�<�6�<�S�<Yo�<���<�I}<�}y<Ӱu<G�q<xn<�Gj<�yf<!�b<�^<�[<JGW<}S<�O<��K<�&H<�bD<�@<��<<%9<�j5<*�1<W .<[P*<	�&<��"<�W<��<s<&�<}�<oo<y�	<�m<u�<|�;�9�;^v�;���;�;	��;�;���;5�;���;뮽;㈷;�v�;�y�;��;=��;���;XV�;�Î;YF�;߃;�};��r;�Xh;&7^; BT;�uJ;�@;�[7;�
.;�$;e�;�;BP
;�;	��:�	�:���:���:ɱ:�,�:�ʒ:���:.Pi:�K:��.:��:���9P��9m�u9�9���7B`��];�����i�ƹJ���% �C�0���I�$c�~"|��y���ϖ����5F��,i��{Ǻ��Ӻjyߺf��E��U���r� S�S/�j�+���$�dv*�@0��6�d�;���A��MG�AM���R��X�B^�^�c�U�i�&ro��+u���z�"P��H-���
�� 舻>Ƌ�Ԥ��񃑻�c��D���%���  �  �=Y#=��=�i=�=��=GR=�� =�� =�8 =A��<���<�8�<6z�<��<���<9:�<�x�<x��<V��<A/�<?j�<-��<��<��<pK�<���<Ĵ�<q��<��<�H�<�v�<x��<l��<���<�<�D�<�g�<T��<o��<@��<���<l��<��<��<_.�<�:�<�C�<�I�<�L�<�K�<�F�<o>�<2�<�!�<;�<i��<-��<f��<���<�c�<�3�<���<���<m��<�@�<;��<0��<�S�<���<���<6�<��<�\�<A��<zn�<��<�k�<��<�T�<·<�*�<ǎ�<g�<�I�<ՠ�<��<�B�<=��<�ը<%�<�Z�<���<Eӡ<�
�<@�<tr�<r��<(И<���<'%�<�L�<�r�<�<f��<�ڋ<}��<3�<�6�<�S�<Uo�<f��<�I}<�}y<��u<;�q<Un<_Gj<tyf<�b<��^<�[<&GW<�|S<ܳO<d�K<�&H<�bD<2�@<��<<�$9<k5<,�1<� .<sP*<.�&<��"<$X<��<�<j�<��<�o<��	<�m<��<��;�9�;v�;���;?�;��;��;d��;5�;;��;���;ڈ�;�v�;>y�;y��;��;���;?V�;<Î;1F�;�ރ;};�r;jXh;�7^;AT;�uJ;P�@;�[7;�.;V�$;��;�;KQ
;�;���:��:���:���:�ɱ:�-�:D˒:ݟ�:�Pi:=�K:Ġ.:��:Z��9∲9+�u9��9;,�7>g��:c;�,����ƹ�����!���0� J�k(c��#|�{��tЖ�����E��i���|Ǻ��ӺDyߺ'e뺿D����]r��R�P.���@��_�$�v*��?0�M6���;��A��MG��M�9�R��X�-B^���c�'�i�_ro��,u���z�:P���-���
���舻�Ƌ��������c��wD���%���  �  �=X#=��=�i=�=��=PR=�� =�� =�8 =Y��<���<�8�<Dz�<���<��<I:�<�x�<���<Y��<Q/�<<j�<>��<��<��<eK�<���<���<c��<��<pH�<�v�<Y��<Q��<���<��<wD�<�g�<>��<\��<;��<���<a��<��<��<p.�<�:�<D�<J�<�L�<�K�<�F�<�>�<22�<�!�<F�<t��<D��<y��<%��<�c�<�3�<���<���<��<�@�<M��<��<�S�<���<���<6�< ��<�\�<#��<in�<t�<}k�<{�<�T�< ·<�*�<Ȏ�<Y�<�I�<Ƞ�<��<�B�<B��< ֨<#�<[�<���<Pӡ<(�<@�<�r�<���<5И<���<D%�<�L�<�r�<і�<g��<�ڋ<���<?�<�6�<uS�<Vo�<X��<�I}<}}y<��u<	�q<n<NGj<Myf<ܫb<��^<j[<GW<�|S<ڳO<@�K<�&H<�bD<1�@<��<<%9<,k5<(�1<� .<{P*<^�&<>�"<NX<�<�<��<��<�o<��	<�m<��<��;&:�;v�;���;�;��;��;2��;5�;��;���;e��;fv�;y�;0��;߼�;^��;�U�;�; F�;�ރ;�};��r;�Wh;8^;�AT;�vJ;��@;�[7;.;��$;�;�;R
;I�;H��:"�:7��:?��: ʱ:�.�:�˒:E��:MSi:I�K:�.:��:e��9���9��u9��9M��7�x��yq;�#���2�ƹz����$��0��J��*c�X#|��{���Ж�]���F���g��%|Ǻv�ӺQyߺ=d뺌D������p�R��-�b������$�u*��>0�'6�9�;��A�MG�7M���R�>�X��B^�u�c���i�vro��,u���z��P���-�����舻�Ƌ�~���n���d���D���%���  �  �=Y#=��=�i=�=��=MR=�� =Ŗ =�8 =Y��<���<�8�<Nz�<��<��<M:�<�x�<���<h��<^/�<Oj�<9��<��<��<bK�<���<´�<b��<��<qH�<�v�<T��<H��<���<��<hD�<�g�<8��<_��<*��<���<d��<��<��<_.�<�:�<D�<J�<�L�<�K�<�F�<�>�<42�<�!�<Z�<���<C��<}��<��<�c�<�3�<���<���<{��<�@�<=��<"��<�S�<���<���<�5�<��<�\�<��<[n�<o�<qk�<q�<�T�<���<�*�<���<W�<�I�<Π�<��<�B�<E��<�ը<2�<[�<���<Yӡ<�<@�<�r�<���<@И<���<=%�<�L�<�r�<ݖ�<{��<�ڋ<���<9�<�6�<|S�<Xo�<X��<�I}<i}y<��u<��q<n<,Gj<Hyf<��b<��^<W[<GW<�|S<��O<A�K<�&H<�bD<�@<��<<%9< k5<M�1<� .<�P*<^�&<%�"<UX<'�<�<��<��<�o<��	<n<��<��;:�;7v�;���;�;��;��;3��;�4�;
��;m��;S��;Fv�;�x�;.��;���;a��;�U�;Î;�E�;�ރ;�};#�r;Xh;�7^;�AT;lvJ;��@;r\7;h.;!�$;��;�;R
;��;���:�:���:d��:˱:W/�:�̒:q��:�Ri:4�K:I�.:�:��9<��9��u9[�9���7t����r;�k���<�ƹ,���"&�k�0��J�5*c��%|��{���Ж�����F���h���{Ǻ݀Ӻ_xߺc뺚C��<���q��Q��-���y����$�Ou*��>0��6���;�H�A�.MG�.M��R���X��B^�f�c���i� so�'-u�	�z��P���-��S��鈻�Ƌ���������(d���D��<&���  �  �=P#=��=�i=�=��=MR=�� =�� =�8 =_��<���<9�<Kz�<��<��<u:�<�x�<���<i��<L/�<Vj�<;��<��<��<hK�<���<���<m��<��<fH�<�v�<Z��<L��<w��<��<YD�<�g�<%��<K��<��<���<[��<�<��<[.�<�:�<D�<	J�<�L�<�K�<G�<�>�<L2�<�!�<U�<���<J��<���<��<�c�<�3�<���<���<���<A�<4��<(��<�S�<���<���<�5�<���<�\�< ��<Sn�<c�<ak�<v�<�T�<���<�*�<���<_�<�I�<���<��<�B�<K��<�ը<7�<[�<���<gӡ<�<@@�<�r�<���<;И<���<O%�<�L�<�r�<ʖ�<{��<�ڋ<���<<�<�6�<�S�<Co�<\��<�I}<[}y<`�u<��q<n<Gj<>yf<��b<��^<H[<�FW<�|S<��O<T�K<|&H<�bD< �@<��<<%%9< k5<T�1<� .<�P*<k�&<C�"<�X<#�<�<��<#�<�o<��	<
n<��<��;:�;Vv�;���;)�;��;��;_��;�4�;���;	��;m��;Yv�;�x�;��;k��;a��;�U�;�;�E�;�ރ;�};Y�r;JXh;}7^;BT;�vJ;��@;r\7;.;T�$;��;};RR
;��;:��:��:b��:��:�˱:/�:s̒:ޠ�:�Si:'�K:7�.:��:@��9I��9��u9��9���7Ϙ��Ur;�J����ƹ*���w%�x�0�-J�,c��&|�V{���і����7F��Ji���{ǺӀӺ�wߺud�tC��ȋ��q��P�K-������$��t*��>0��6�q�;�G�A�6MG��M���R���X�tB^��c�v�i��ro�`-u���z��P���-�����鈻<ǋ���������zd���D��0&���  �  �=Y#=��=�i=�=��=MR=�� =Ŗ =�8 =Y��<���<�8�<Nz�<��<��<M:�<�x�<���<h��<^/�<Oj�<9��<��<��<bK�<���<´�<b��<��<qH�<�v�<T��<H��<���<��<hD�<�g�<8��<_��<*��<���<d��<��<��<_.�<�:�<D�<J�<�L�<�K�<�F�<�>�<42�<�!�<Z�<���<C��<}��<��<�c�<�3�<���<���<{��<�@�<=��<"��<�S�<���<���<�5�<��<�\�<��<[n�<o�<qk�<q�<�T�<���<�*�<���<W�<�I�<Π�<��<�B�<E��<�ը<2�<[�<���<Yӡ<�<@�<�r�<���<@И<���<=%�<�L�<�r�<ݖ�<{��<�ڋ<���<9�<�6�<|S�<Xo�<X��<�I}<i}y<��u<��q<n<,Gj<Hyf<��b<��^<W[<GW<�|S<��O<A�K<�&H<�bD<�@<��<<%9< k5<M�1<� .<�P*<^�&<%�"<UX<'�<�<��<��<�o<��	<n<��<��;:�;7v�;���;�;��;��;3��;�4�;
��;m��;S��;Fv�;�x�;.��;���;a��;�U�;Î;�E�;�ރ;�};#�r;Xh;�7^;�AT;lvJ;��@;r\7;h.;!�$;��;�;R
;��;���:�:���:d��:˱:W/�:�̒:q��:�Ri:4�K:I�.:�:��9<��9��u9[�9���7t����r;�k���<�ƹ,���"&�k�0��J�5*c��%|��{���Ж�����F���h���{Ǻ݀Ӻ_xߺc뺚C��<���q��Q��-���y����$�Ou*��>0��6���;�H�A�.MG�.M��R���X��B^�f�c���i� so�'-u�	�z��P���-��S��鈻�Ƌ���������(d���D��<&���  �  �=X#=��=�i=�=��=PR=�� =�� =�8 =Y��<���<�8�<Dz�<���<��<I:�<�x�<���<Y��<Q/�<<j�<>��<��<��<eK�<���<���<c��<��<pH�<�v�<Y��<Q��<���<��<wD�<�g�<>��<\��<;��<���<a��<��<��<p.�<�:�<D�<J�<�L�<�K�<�F�<�>�<22�<�!�<F�<t��<D��<y��<%��<�c�<�3�<���<���<��<�@�<M��<��<�S�<���<���<6�< ��<�\�<#��<in�<t�<}k�<{�<�T�< ·<�*�<Ȏ�<Y�<�I�<Ƞ�<��<�B�<B��< ֨<#�<[�<���<Pӡ<(�<@�<�r�<���<5И<���<D%�<�L�<�r�<і�<g��<�ڋ<���<?�<�6�<uS�<Vo�<X��<�I}<}}y<��u<	�q<n<NGj<Myf<ܫb<��^<j[<GW<�|S<ڳO<@�K<�&H<�bD<1�@<��<<%9<,k5<(�1<� .<{P*<^�&<>�"<NX<�<�<��<��<�o<��	<�m<��<��;&:�;v�;���;�;��;��;2��;5�;��;���;e��;fv�;y�;0��;߼�;^��;�U�;�; F�;�ރ;�};��r;�Wh;8^;�AT;�vJ;��@;�[7;.;��$;�;�;R
;I�;H��:"�:7��:?��: ʱ:�.�:�˒:E��:MSi:I�K:�.:��:e��9���9��u9��9M��7�x��yq;�#���2�ƹz����$��0��J��*c�X#|��{���Ж�]���F���g��%|Ǻv�ӺQyߺ=d뺌D������p�R��-�b������$�u*��>0�'6�9�;��A�MG�7M���R�>�X��B^�u�c���i�vro��,u���z��P���-�����舻�Ƌ�~���n���d���D���%���  �  �=Y#=��=�i=�=��=GR=�� =�� =�8 =A��<���<�8�<6z�<��<���<9:�<�x�<x��<V��<A/�<?j�<-��<��<��<pK�<���<Ĵ�<q��<��<�H�<�v�<x��<l��<���<�<�D�<�g�<T��<o��<@��<���<l��<��<��<_.�<�:�<�C�<�I�<�L�<�K�<�F�<o>�<2�<�!�<;�<i��<-��<f��<���<�c�<�3�<���<���<m��<�@�<;��<0��<�S�<���<���<6�<��<�\�<A��<zn�<��<�k�<��<�T�<·<�*�<ǎ�<g�<�I�<ՠ�<��<�B�<=��<�ը<%�<�Z�<���<Eӡ<�
�<@�<tr�<r��<(И<���<'%�<�L�<�r�<�<f��<�ڋ<}��<3�<�6�<�S�<Uo�<f��<�I}<�}y<��u<;�q<Un<_Gj<tyf<�b<��^<�[<&GW<�|S<ܳO<d�K<�&H<�bD<2�@<��<<�$9<k5<,�1<� .<sP*<.�&<��"<$X<��<�<j�<��<�o<��	<�m<��<��;�9�;v�;���;?�;��;��;d��;5�;;��;���;ڈ�;�v�;>y�;y��;��;���;?V�;<Î;1F�;�ރ;};�r;jXh;�7^;AT;�uJ;P�@;�[7;�.;V�$;��;�;KQ
;�;���:��:���:���:�ɱ:�-�:D˒:ݟ�:�Pi:=�K:Ġ.:��:Z��9∲9+�u9��9;,�7>g��:c;�,����ƹ�����!���0� J�k(c��#|�{��tЖ�����E��i���|Ǻ��ӺDyߺ'e뺿D����]r��R�P.���@��_�$�v*��?0�M6���;��A��MG��M�9�R��X�-B^���c�'�i�_ro��,u���z�:P���-���
���舻�Ƌ��������c��wD���%���  �  �=\#=��=�i=�=��=?R=�� =�� =�8 =/��<���<�8�<z�<ٺ�<���<&:�<�x�<i��<D��<./�<>j�<��<$��<��<cK�<���<д�<���<��<�H�<�v�<|��<x��<���<(�<�D�<h�<[��<���<L��<���<���<��<��<R.�<�:�<�C�<�I�<�L�<tK�<�F�<`>�<2�<�!�<"�<R��<��<`��<��<�c�<�3�<���<���<i��<A�<3��<4��<�S�<���<���<6�<4��<�\�<P��<�n�<��<�k�<��<�T�<·<�*�<Ҏ�<�<�I�<Ԡ�<��<�B�<W��<�ը<$�<�Z�<���<8ӡ<�
�<�?�<Tr�<`��<И<���<%�<�L�<�r�<���<e��<�ڋ<���<B�<�6�<�S�<Yo�<���<�I}<�}y<Ӱu<G�q<xn<�Gj<�yf<!�b<�^<�[<JGW<}S<�O<��K<�&H<�bD<�@<��<<%9<�j5<*�1<X .<[P*<	�&<��"<�W<��<s<&�<}�<oo<y�	<�m<u�<|�;�9�;^v�;���;�;	��;�;���;5�;���;뮽;㈷;�v�;�y�;��;=��;���;XV�;�Î;YF�;߃;�};��r;�Xh;&7^; BT;�uJ;�@;�[7;�
.;�$;e�;�;BP
;�;	��:�	�:���:���:ɱ:�,�:�ʒ:���:.Pi:�K:��.:��:���9P��9m�u9�9���7B`��];�����i�ƹJ���% �C�0���I�$c�~"|��y���ϖ����5F��,i��{Ǻ��Ӻjyߺf��E��U���r� S�S/�j�+���$�dv*�@0��6�d�;���A��MG�AM���R��X�B^�^�c�U�i�&ro��+u���z�"P��H-���
�� 舻>Ƌ�Ԥ��񃑻�c��D���%���  �  �=c#=��=�i=�=��==R=�� =�� =~8 =��<���<�8�<�y�<���<���<:�<�x�<M��</��<!/�<)j�<��<��<��<rK�<π�<ش�<���<��<�H�<�v�<���<���<���<3�<�D�<%h�<~��<���<_��<���<���<��<��<d.�<�:�<�C�<�I�<mL�<gK�<�F�<K>�<�1�<�!�<�<2��<���<>��<ێ�<�c�<�3�<���<���<a��<A�<B��<;��<�S�<���<Ú�<16�<@��<]�<u��<�n�<��<�k�<��<�T�<?·<�*�<쎴<��<�I�<堯<��<�B�<G��<�ը<�<�Z�<���<ӡ<�
�<�?�<Dr�<=��<�Ϙ<~��<%�<�L�<ur�<���<O��<�ڋ<q��<9�<�6�<�S�<fo�<���<�I}<�}y<��u<��q<�n<�Gj<�yf<b�b<A�^<�[<�GW<#}S<�O<��K<�&H<�bD<3�@<��<<�$9<�j5<��1<B .<-P*<У&<��"<�W<~�< <��<G�<Xo<>�	<�m<W�<$�;v9�;v�;���;9�;?��;,�;Ô�;w5�;���;a��;l��;rw�;�y�;4��;½�;}��;�V�;�Î;�F�;B߃;�};7�r;�Xh;�7^;�AT;puJ;��@;�Z7;{
.;'�$;��;�;�O
;�;���:Y�:V��:o��:.Ǳ:�+�:�ɒ:���:Oi:R�K:E�.:{�:P��9���9��u9��9���7�<��8K;�\{���ƹ׿������0�j�I�U#c��|�7y��1ϖ�����E���h��|Ǻ�Ӻ�zߺg�!G��?��?s��S��/�������$�8w*��@0�Y6���;���A�NG��M��R�a�X��A^���c�@�i��qo�O+u�5�z��O���,��
���爻�ŋ�b���]���-c���C��z%���  �  �=k#=��=�i=�=��==R=�� =�� =t8 = ��<���<�8�<�y�<���<���<�9�<�x�<4��< ��</�<j�<��<��<��<lK�<΀�<��<���<��<�H�<w�<���<���<���<V�<�D�<5h�<���<���<��<���<���<��<��<`.�<�:�<�C�<�I�<SL�<`K�<�F�<7>�<�1�<y!�<��<��<���<��<ǎ�<�c�<�3�<���<���<g��<�@�<B��<9��<�S�<
��<Ԛ�<S6�<X��<"]�<���<�n�<��<�k�<��<�T�<Z·<�*�<��<��<�I�<�<��<�B�<:��<�ը<�<�Z�<x��<ӡ<�
�<�?�<4r�<!��<�Ϙ<]��<�$�<�L�<]r�<���<4��<�ڋ<n��</�<�6�<�S�<wo�<���<J}<~y<&�u<��q<�n<Hj<zf<��b<p�^< [<�GW<Y}S<L�O<��K<�&H<�bD<)�@<��<<�$9<�j5<ȳ1<. .<P*<��&<g�"<}W<\�<�<ۈ<��<o<	�	<hm<:�<��;�9�;�u�;x��;�;4��;e�;ޔ�;�5�;%��;���;���;�w�;xz�;���;Q��;���;OW�;Ď;G�;�߃; };ۤr;�Xh;{7^;6AT;nuJ;;�@;Z7;>
.;E�$;
�;|;�N
;>�;H��:>�:��:��:�ű:+�:Ȓ:���:Oi:m�K:��.:�:	��9��9�u9��9!�7���D;��r����ƹ������0�r�I�r c�v|��x��HΖ�����E���h��
}Ǻ��Ӻ�{ߺh��G����t�@U�d0�g����ī$�Mx*�wA0�6���;�}�A�<NG�
M�Y�R���X��A^�g�c���i��po�*u���z�,O���,���	��t爻4ŋ����
����b��rC��%���  �  �=k#=��=�i=�=��=4R=�� =�� =g8 =��<z��<i8�<�y�<s��<���<�9�<dx�< ��<��<�.�<j�<	��<��<��<xK�<р�<��<���<��<�H�<w�<գ�<���<
��<q�<�D�<\h�<���<Ũ�<���<���<���<��<
�<b.�<�:�<�C�<�I�<IL�<@K�<�F�<>�<�1�<Z!�<��<���<���<��<���<�c�<�3�<���<���<X��<�@�<E��<J��<�S�<��<��<a6�<t��<;]�<���<�n�<��<�k�<�<&U�<p·<+�<��<��<�I�<<��<�B�<A��<�ը<��<�Z�<\��<�ҡ<�
�<�?�<r�<���<�Ϙ<A��<�$�<oL�<Fr�<{��<+��<pڋ<o��<4�<�6�<�S�<to�<���<3J}<6~y<X�u<�q<*n<7Hj<Szf<Ǭb<��^<e[<�GW<�}S<b�O<��K<�&H<cD<5�@<��<<�$9<�j5<��1<��-<�O*<��&<A�"<KW<�<�<��<��<�n<��	</m<�<��;-9�;�u�;���;=�;4��;|�;=��;�5�;}��;;-��;Rx�;�z�;��;���;I �;�W�;yĎ;EG�;�߃;�};��r;�Xh;�7^;XAT; uJ;��@;�Y7;4	.;��$;<�;�;�M
;D�;:��:�:��:A��:&ı:)�:&ǒ:ݜ�:�Mi:��K:4�.:��:���9���9��u9�9��79��M1;��n���ƹ�����
�0���I�,c��|��v��g͖�����D���h���|Ǻ؃Ӻk|ߺVi��I�����u��U��1�z	������$��x*�B0��6���;���A��NG��M�*�R�j�X��A^���c�:�i�hpo��)u���z��N���+��D	���戻�ċ�n��������b��&C���$���  �  �=l#=��=�i=�=��=.R=�� =�� =a8 =г�<T��<K8�<�y�<g��<e��<�9�<Bx�<��<���<�.�<j�<���<���<��<�K�<��<���<���<�<�H�<8w�<��<���<)��<��<�D�<}h�<�<��<���<���<���<��<�<[.�<�:�<�C�<�I�<AL�<)K�<�F�<�=�<�1�<8!�<��<���<���<��<���<|c�<p3�<���<���<N��<�@�<;��<Z��<�S�<.��<���<r6�<���<L]�<���<�n�<#�<"l�<�<HU�<�·<0+�<'��<��<�I�< ��<��<�B�<;��<�ը<��<�Z�<J��<�ҡ<�
�<�?�<�q�<���<�Ϙ<"��<�$�<PL�<=r�<b��<(��<fڋ<`��<$�<�6�<�S�<xo�<���<MJ}<`~y<��u<�q<Yn<bHj<�zf<��b<��^<�[<HW<�}S<x�O<�K<�&H<1cD<=�@<��<<�$9<�j5<��1<��-<�O*<E�&<��"<W<ط<�<E�<��<�n<��	<m<��<��;�8�;�u�;.��;[�;}��;��;���;!6�;���;L��;���;�x�;6{�;���;ʾ�;� �;�W�;�Ď;�G�;��;"};��r;bYh;>7^;AT;�tJ;��@;dY7;q.;X�$;%�;�;�L
;��;B��:��:���:���:�ñ:�'�:�ƒ:m��:Li:)�K:��.:��:Z��9���9�v9�
9���7 ����;�;j����ƹ������%�0��I��c�|��u���̖����ED���i��:}Ǻ��Ӻ�|ߺIj��J��)��v��V��2��	�|����$�z*�C0�	6���;�ݎA�OG�pM���R�m�X��@^�b�c���i�po�P)u���z�{N���+�����Q戻�ċ����:���b���B���$���  �  �=u#=��=�i=�=��=*R=w� =�� =S8 =���<N��<<8�<�y�<B��<Q��<�9�<<x�<���<���<�.�<�i�<���<���<��<qK�<ހ�< ��<���< �<�H�<Iw�<���<��<F��<��<E�<�h�<Ӊ�<��<���<���<���<��<�<_.�<�:�<�C�<�I�<-L�< K�<gF�<�=�<�1�<+!�<��<���<���<ߴ�<���<^c�<h3�<u��<u��<R��<�@�<D��<E��<�S�<4��<��<�6�<���<^]�<���<"o�<;�<?l�<=�<RU�<�·<;+�<A��<��<J�<��<��<�B�<8��<�ը<��<�Z�<=��<�ҡ<�
�<t?�<�q�<ϡ�<�Ϙ<��<�$�<AL�<r�<[��<��<\ڋ<`��<3�<�6�<�S�<�o�<���<uJ}<�~y<��u<@�q<�n<�Hj<�zf<:�b<�^<�[</HW<�}S<��O<�K<'H<cD<0�@<��<<�$9<�j5<�1<��-<~O*<"�&<��"<�V<��<:<�<g�<�n<��	<�l<��<�;�8�;�u�;f��;�;[��;��;���;x6�;���;���;���;�x�;�{�;璥;J��;� �;X�;Ŏ;�G�;8��;7};%�r;�Xh;W7^;(AT;�tJ;�@;�X7;!.;B�$;��;�;mL
;��;ݘ�:��:��:���:���:'�:�Œ:k��:bLi:�K:��.:��:���9���9d	v9`9m#�7w頸&;��a��X�ƹ�����&�0��I��c�|�cu��|̖�����E���h��~}Ǻ��Ӻ5~ߺ�j��K����Wv�=W�!3��c���$�%z*��C0�
6���;���A�eOG�qM�6�R�~�X��A^���c���i�boo��(u�~�z�4N��3+��k��戻ċ����������a���B��g$���  �  �=~#=��=�i=�=��=)R=o� =�� =L8 =���<5��<#8�<�y�<.��<I��<�9�<#x�<��<���<�.�<�i�<���<���<��<|K�<��<��<���<.�< I�<fw�<��<��<R��<��<3E�<�h�<���<���<���<��<���<��<
�<q.�<�:�<�C�<�I�<!L�<!K�<TF�<�=�<v1�<!�<��<���<���<´�<s��<Kc�<h3�<i��<m��<J��<�@�<X��<M��<�S�<9��<��<�6�<���<�]�<���<;o�<I�<Kl�<W�<lU�<�·<C+�<O��<��<J�<��<��<C�< ��<�ը<��<�Z�<7��<�ҡ<k
�<X?�<�q�<���<|Ϙ<���<�$�<6L�<r�<^��< ��<Zڋ<P��<*�<�6�<�S�<�o�<���<�J}<�~y<ӱu<��q<�n<�Hj<�zf<Y�b<>�^<�[<[HW<�}S<ŴO<
�K<:'H<cD<K�@<��<<�$9<�j5<^�1<��-<bO*<
�&<��"<�V<��<<	�<,�<On<d�	<�l<��<�
�;�8�;(u�;���;9�;���;��;���;�6�;��;���;%��;Vy�;�{�;��;���;*�;�X�;7Ŏ;�G�;k��;0};��r;�Xh;�7^;�@T;ZtJ;��@;UX7;(.;��$;d�;�;�K
;8�;��:� �:;��:���:`��:	'�:�Ē:ܚ�:/Ki:9�K:�.:��:g��9��9�v9i9IC�7u���;��[���ƹ[������0���I��c�}|�#u���˖�����D���g��Ǻ��Ӻ�~ߺlk�@L��x��w� X�w3������ݮ$�{*��C0��
6���;��A�wOG��M�z�R���X�jA^�P�c���i��no��(u���z��M���*��'���刻�Ë�q���j����a���B��#$���  �  �=z#=��=�i=�=��=+R=o� =|� =K8 =���<,��<8�<{y�<-��<8��<�9�<x�<��<���<�.�<�i�<���<���<��<wK�<��<��<���<;�<I�<cw�<��<��<`��<��<5E�<�h�<��<��<���<��<���<��<�<d.�<�:�<�C�<�I�<L�<K�<YF�<�=�<s1�<
!�<��<���<y��<���<j��<Pc�<U3�<b��<p��<Q��<�@�<K��<N��<�S�<@��<&��<�6�<���<}]�<���<=o�<a�<_l�<W�<mU�<�·<V+�<[��<��<J�<��<��<�B�<-��<�ը<��<�Z�<(��<�ҡ<f
�<Y?�<�q�<���<oϘ<���<�$�<,L�<r�<H��< ��<[ڋ<Y��<%�<�6�<�S�<�o�<Ǌ�<�J}<�~y<ڱu<m�q<�n<�Hj<{f<j�b<D�^<�[<]HW<�}S<ݴO<-�K<-'H<'cD<7�@<��<<�$9<�j5<^�1<��-<ZO*<��&<��"<�V<p�<<�<,�<?n<`�	<�l<��<�
�;�8�;Fu�;M��;"�;���;��;ݕ�;�6�;Q��;鰽;��;Sy�;|�;t��;���;>�;rX�;eŎ;H�;���;�};{�r;�Xh;v7^;�@T;�tJ;��@;;X7;�.;��$;�;q;WK
;�;���:���:���:���:���:�%�:^Ē:���:�Ki:��K:>�.:��:E��9���9v9�9W��7�̠�t;��[��Q�ƹ�������0���I��c�|� t���˖����E��i��T~ǺN�Ӻ�~ߺIl�8M��f��Bw�X��3������$�={*�5D0��
6�}�;��A�lOG��M���R�W�X�7A^�w�c��i�~no�5(u���z��M���*����|刻�Ë�f��������a��FB���#���  �  �=�%=��=(m=~=��=�V=A� =�� =�= =ӿ�<H�<$F�<p��<B��<0�<�K�<M��<D��<f�<�E�<��<7��<���<�0�<�h�<���<C��<�	�<B<�<�m�<���<���<���<w#�<�L�<�s�<��<��</��<���<��<�1�<�H�<�\�<�m�<4|�<4��<���<]��<'��<V��<���<��<Fq�<^�<WG�<�+�<u�<f��<���<��<Z�<� �<���<���<�U�<X�<��<lY�<��<1��< +�<���<�E�<˿<K�<�ż<y;�<��<��<�~�<��<p>�<���<{�<7=�<ۉ�<�Ҫ<��<�Y�<Ɨ�<�ң<�
�<�?�<Zr�<��<�Ϛ<���<�#�<�J�<�o�<,��<մ�<Ս<��<b�<�-�<I�<dc�<�|�<}��<�Z}<�y<��u<��q<�n<@j<�mf<B�b<y�^<��Z<�'W<FXS<�O<��K<��G<�)D<�b@<+�<<�8<�5<�`1<��-<c�)<�@&<G�"<,�<�E<��<<�w<��<�_	<p�<�a<O��;���;�1�;�t�;x��;�,�;��;@)�;��;�o�;�/�;�;��;h�;s��;&�;e�;\��;�$�;ʥ�;�=�;�y;bo;�e;Z�Z;�Q;�AG;k�=;�54;�*;��!;a�;�	;�_;���:M��:�}�:�I�:JS�:���:�$�:M�:0�}:�`:��B:��%:�q	::��9/Ԣ9�W9=�8�1���ظЩU��5��gӹ3G�@��>6�><O��,h��}��͌�����8���U��vd���cɺ�Vպx;Ẳ�e����R�!0�V�d��E��!u��<%�} +���0��6�$<<��A�׮G�CeM��S���X��^�V7d�g�i�Z�o�iQu�,{�M\���5�����눻+Ƌ�D����}��wZ��D8��9���  �  �=�%=��=$m=�=��=�V=E� =�� =�= =ֿ�<I�<-F�<s��<$��<;�<�K�<V��<C��<Y�<�E�<��<P��<���<�0�<�h�<���</��<y	�<S<�<�m�<���<���<���<�#�<�L�<�s�<��<%��<��<���<��<1�<zH�<�\�<�m�<8|�<J��<��<b��<$��<N��<���<��<Uq�<q^�<?G�<�+�<n�<s��<���<ߍ�<Z�<	!�<���<��<�U�<6�<��<RY�<��<@��<�*�<��<�E�<˿<K�<�ż<p;�<��<��<�~�<��<f>�<���<i�<=�<މ�<�Ҫ<��<�Y�<ʗ�<�ң<�
�<�?�<[r�<��<�Ϛ<���<�#�<�J�<�o�<��<Դ�<Ս<��<q�<�-�<�H�<Fc�<�|�<j��<[}<�y<f�u<�q<Xn<�@j<�mf<N�b<E�^<��Z<�'W<@XS<<�O<��K<��G<�)D<�b@<3�<<.�8<�5<�`1<��-<C�)<�@&<H�"<?�<�E<N�<"<�w<��<�_	<V�<�a<~��;G��;�1�;�t�;,��;S,�;���;)�;���;o�;�/�;��;��;��;���;$&�;�d�;|��;�$�;���;>�;B�y;�ao;�e;C�Z;�Q;�BG;)�=;�54;��*;��!;��;v	;`;���:���:�~�:)I�:T�:���:�$�:��:�}:�`:*�B:��%:Bm	:<��9�͢9��W9��8����ظ��U�W6��ӹ,E�N��t6��;O�~/h��|���͌�3���9��W��<d��KcɺUպ�:�t����S��/�N���8��$u�_<%�� +���0� �6�.<<���A���G��dM��S���X��^��7d���i�ϝo�\Qu��{�E\��>6��}���ꈻƋ������}���Z��P8������  �  ��=�%=��=)m=~=��=�V=B� =Û =�= =��<P�<9F�<���<7��<^�<�K�<d��<O��<d�<�E�<��<H��<���<�0�<�h�<���<=��<i	�<T<�<�m�<���<���<|��<e#�<L�<�s�<���<*��<���<���<��<w1�<�H�<�\�<n�<)|�<;��<��<d��<6��<R��<���< ��<rq�<�^�<YG�<�+�<h�<���<���<��<Z�<� �<���<��<�U�<4�<"��<PY�<��<@��<�*�<
��<�E�<�ʿ<�J�<�ż<a;�<���<��<~~�<��<U>�<���<{�<=�<艬<�Ҫ<��<�Y�<՗�<�ң<�
�< @�<Xr�<A��<�Ϛ<���<�#�<�J�<�o�<#��<鴏<Ս<��<^�<�-�<I�<Kc�<�|�<^��<�Z}<��y<:�u< �q<9n<i@j<�mf<)�b<(�^<��Z<y'W<XS<0�O<y�K<��G<�)D<�b@<*�<<	�8<�5<�`1<ϧ-<S�)<�@&<X�"<V�<F<v�<i<�w<��<�_	<n�<�a<e��;,��;�1�;u�;E��;�,�;ա�;�(�;���;o�;�/�;��;z�;$�;"��;�%�;�d�;���;0$�;���;�=�;�y;�bo;�e;��Z;lQ;#BG;̦=;�54;��*;��!;~�;]	;a;���:w��:���:�H�:LU�:؞�:�%�:�:F�}:`:.�B:��%:3m	:]��9q͢9zW9v�8-!����׸m�U��9�� ӹCI����6�X<O�M3h��|���Ό�|���8���V���c��Vdɺ�Uպ_;Ặ�J����R�4/�`�������;t��;%�i +��0��6��;<���A�<�G�beM��S�`�X�ʃ^��6d�b�i��o��Qu�E{�I\��{6�����{눻[Ƌ�衎��}���Z���8������  �  ��=�%=��=$m=�=��=�V=K� =Ǜ => =���<l�<KF�<���<X��<c�<�K�<}��<_��<�<�E�<���<a��<���<�0�<�h�<���<-��<a	�<><�<�m�<|��<���<u��<X#�<hL�<�s�<��<��<���<���<��<y1�<rH�<�\�<�m�<8|�<\��<��<v��<G��<e��<Ê�<$��<xq�<�^�<nG�<�+�<��<���<���<���<Z�<!�<���<��<�U�</�< ��<MY�<���<*��<�*�<��<�E�<�ʿ<�J�<�ż<W;�<߫�<��<}~�<��<G>�<~��<\�<=�<ቬ<�Ҫ< �<�Y�<���<�ң<�
�<@�<vr�<G��<�Ϛ<���<�#�<�J�<�o�<<��<���<(Ս<��<�<�-�<�H�<=c�<�|�<^��<�Z}<�y<�u<��q<"n<O@j<Wmf<�b<�^<��Z<O'W<XS<��O<p�K<��G<�)D<�b@<3�<<G�8<
5<�`1<�-<��)<�@&<��"<}�<F<��<v<�w<��<`	<��<�a<���;���;2�;u�;B��;1,�;���;�(�;|��;o�;B/�;O�;c�;��;���;�%�;=d�;���;$�;���;�=�;!�y;�ao;�e;��Z;�Q;8CG;��=;�64;�*;^�!;�;�
;;a;���:���:��:K�:�V�:��:�&�:��:�}:+`:J�B:G�%:�l	:I~�9͢9�nW9���8e����$ظ��U�A;���$ӹ�J���e 6��?O�&3h�~��nό�D���:��W���c���bɺ�Sպ:�������7R�q.�l��������s�d;%�l�*���0�6�$;<�O�A���G�]dM��S���X�9�^��7d�c�i��o�Ru��{��\���6������눻�Ƌ�
���v~��&[���8��`���  �  ��=�%=��=&m=}=��=�V=X� =Λ => =��<��<tF�<���<~��<�<�K�<���<u��<��<�E�<��<S��<���<�0�<�h�<���<"��<X	�<<�<�m�<`��<���<F��<4#�<YL�<�s�<Ř�<��<���<���<��<x1�<gH�<�\�<�m�<5|�<N��<��<���<W��<���<ϊ�<O��<�q�<�^�<�G�<�+�<��<���<߼�<��<4Z�<!�<���<���<�U�<?�<���<GY�<���<��<�*�<º�<sE�<�ʿ<�J�<�ż<$;�<ɫ�<{�<e~�<��<:>�<s��<X�<)=�<ω�<�Ҫ<��<�Y�<<ӣ<�<)@�<�r�<a��<�Ϛ<���<�#�<�J�<�o�<[��<��<?Ս<��<x�<�-�<�H�<Lc�<�|�<Z��<�Z}<��y<�u<��q<�n<�?j<Cmf<��b<��^<{�Z<'W<�WS<ȉO<g�K<w�G<�)D<�b@<%�<<<�8<�5<�`1<��-<��)<A&<ӓ"<��<YF<�<�<)x<!�<?`	<��<�a<%��;e��;
2�;�t�;x��;B,�;v��;�(�;���;�n�;�.�;�;��;q�;���;#%�;�c�;���;�#�;Q��;:=�;&�y;Iao;be;G�Z;�Q;�BG;��=;074;��*;d�!;y�;�;=b;׼�:5��:Ԃ�:�M�:�W�:��:(�:X�:<�}:;`:��B:U�%:�n	::|�96̢9\gW9��8ݯ��BظI�U��G��8*ӹ�N����"6�cCO��5h����Ќ�����:��V���d���bɺ�Tպ�8���m���gQ��-������v���r�):%�Q�*�$�0�~6��:<���A���G��dM��S���X�Ń^�o8d��i���o��Ru�z{�4]��C7�����숻Aǋ������~���[��
9������  �  �=�%=��=!m=�=��=�V=b� =ڛ => =5��<��<�F�<��<���<��<L�<���<���<��<�E�<+��<]��<���<�0�<�h�<���<��<;	�<<�<fm�<=��<���<#��<#�<3L�<`s�<���<λ�<���<m��<��<X1�<\H�<�\�<�m�<O|�<W��<2��<���<i��<���<���<d��<�q�<�^�<�G�<,�<��<���<���<!��<HZ�<-!�<���<��<�U�<"�<��<(Y�<���<���<*�<���<QE�<�ʿ<�J�<`ż<�:�<���<W�<=~�<z�<>�<\��<B�<=�<܉�<�Ҫ<��<�Y�<��<ӣ<-�<K@�<�r�<���<�Ϛ<��<$�<K�<p�<o��<��<SՍ<�<��<�-�<�H�<6c�<�|�<;��<sZ}<��y<��u<U�q<�n<�?j<�lf<r�b<y�^<G�Z<�&W<�WS<��O<&�K<c�G<|)D<�b@<N�<<Q�8<5<a1<,�-<��)<tA&<�"<�<�F<<�<<Yx<n�<�`	<�<!b<��;���;Y2�;9u�;@��;,�;F��;7(�;���;Ln�;Z.�;��;-�;��;	��;�$�;Zc�;:��;1#�;��;�<�;7�y; ao;�e;Y�Z;�	Q;&CG;g�=;�74;@�*;V�!;��;�;gc;��:��::��:0O�:�Y�:%��:2)�:��:�}:=`:A�B:(�%:�k	:�x�9�Ģ9�\W9���84`��_\ظw�U�
Q��,3ӹS�p��v&6�oGO�u:h�����ь�
���;��sW���c���aɺNTպy7ẙ�.���%P��,�Q��������q�;9%�^�*�ξ0�u}6�:<���A�%�G�]dM�S���X�x�^��8d�x�i�G�o��Su��{��]���7��#���숻�ǋ�>���)��\��9�����  �  �=�%=��="m=�=��=�V=g� =� =*> =T��<��<�F�<��<���<��<+L�<ڋ�<���<��<�E�<8��<|��<���<�0�<�h�<���<
��<,	�<�;�<Gm�<!��<_��<��<�"�<L�<Ds�<v��<���<���<O��<��<K1�<TH�<�\�<�m�<E|�<f��<L��<���<���<���<��<���<�q�<_�<�G�<3,�<��<���<��<B��<WZ�<A!�<���<
��<�U�<�<޲�<Y�<���<Ԕ�<e*�<���<E�<qʿ<iJ�<5ż<�:�<w��<8�<~�<]�<	>�<S��<;�<=�<؉�<�Ҫ<�<�Y�<��<8ӣ<@�<p@�<�r�<���<К<=��<0$�<&K�<<p�<���<;��<_Ս<%�<��<�-�<�H�<-c�<�|�<+��<NZ}<F�y<b�u<�q<5n<p?j<�lf<1�b<$�^<��Z<�&W<bWS<t�O<�K<U�G<h)D<�b@<D�<<Z�8<W5<3a1<j�-<(�)<�A&<V�"<R�<G<��<i<�x<��<�`	<L�<\b<���;��;V2�;<u�;N��;�+�;0��;(�;z��;�m�;�-�;��;��;h�;O��;($�;�b�;���;�"�;���;�<�;��y;�`o;qe;s�Z;{	Q;�CG;C�=;c84;f�*;�!;�;�;�d;���:��:��:Q�:�\�:���:b+�:��:��}:�`:��B:7�%:!k	:ww�9�¢9�SW9 ��8���}ظp�U��X���>ӹ�W�{��B,6��JO�>h������Ҍ�t��"<��jW��d��+bɺ�Rպ�6�����O��+�o�+��w��Sp�8%�e�*���0��|6��8<���A�0�G�dM�FS���X���^��8d���i�ڠo��Tu��{�<^��~8�����z툻Bȋ�棎�����\��:��n���  �  ܁=�%=��=$m=�=��=�V=p� =� =:> =p��<��<�F�<0��<���<��<WL�<��<���<��<F�<G��<���<���<�0�<�h�<w��<���<	�<�;�<,m�<���<A��<���<�"�<�K�<s�<Z��<���<���<-��<y�<;1�<;H�<�\�<�m�<E|�<i��<R��<���<���<ӑ�<:��<���<r�<4_�<H�<Q,�<�<��<+��<^��<fZ�<G!�<���<
��<�U�<$�<Ų�<Y�<���<���<K*�<T��<�D�<Bʿ<<J�<ż<�:�<V��<�<~�<6�<�=�<4��<*�<=�<Ӊ�<�Ҫ<�<�Y�<'��<Vӣ<Y�<�@�<�r�<Ң�<GК<`��<S$�<RK�<Xp�<���<Q��<pՍ<.�<��<�-�<�H�<0c�<r|�<��<Z}<�y<1�u<��q<�n<?j<Glf<ҙb<��^<��Z<\&W<#WS<9�O<�K<�G<b)D<�b@<B�<<o�8<e5<Ua1<��-<i�)<�A&<��"<��<QG<��<�<�x<	�<a	<��<�b<��;B��;�2�;>u�;m��;�+�;Ġ�;�'�;���;{m�;n-�;��;"�;��;���;�#�;Bb�;��;�"�;��;j<�;l�y;`o;�e;��Z;�	Q;�CG;�=;�84;H�*;��!;��;;�e;R��:��:���: T�:�^�:��:6-�:��:��}:+`:Q�B:H�%:}l	:r�9o��9FKW9O��8��ŵ�ظL
V��c���Hӹ�]�����/6��OO�Ah�񄀺�ӌ�7�� =���V��,d���aɺ$Rպ�5������N�n*��F����5o��6%�	�*�ּ0��{6�L8<��A��G��cM�KS���X���^��9d�W�i���o��Uu�b	{��^���8��[���ȋ�i���R��� ]��|:������  �  ҁ=�%=��=m=�=��=�V=� =�� =I> =���<�<�F�<Q��<��<�<zL�<��<���<	�<F�<f��<���<���<�0�<�h�<o��<���<	�<�;�<m�<М�<$��<���<�"�<�K�<�r�<F��<`��<a��<��<c�<%1�<4H�<�\�<�m�<]|�<|��<h��<֓�<���<���<X��<̀�<%r�<U_�<%H�<t,�<2�<,��<S��<o��<{Z�<a!�<���<"��<�U�<�<���<�X�<���<���<%*�<.��<�D�<ʿ<J�<�ļ<�:�<;��<��<�}�< �<�=�<��<�<�<�<Ӊ�<�Ҫ<�<�Y�<9��<iӣ<��<�@�<s�<���<lК<���<u$�<nK�<}p�<ʓ�<b��<�Ս<:�<��<�-�<�H�< c�<g|�<��<�Y}<߈y<޶u<z�q<�n<�>j<lf<�b<��^<i�Z<&W<�VS<	�O<üK<��G<I)D<�b@<V�<<��8<y5<�a1<��-<��)<<B&<�"<��<�G<A�<�<<y<A�<^a	<��<�b<���;i��;�2�;`u�;#��;�+�;���;�'�;���;2m�;�,�;'�;��;6�;]��;�"�;�a�;���;�!�;ͣ�;<�;��y;�_o;$e;/�Z;P
Q;pDG;<�=;�94;��*;-�!;��;�;�f;s��:��:K��:�U�:>`�:���:^.�:E�:X�}:5`:��B:4�%:9i	:;p�9��9m@W9`|�8�yε�ظ�V��m���Oӹ�a�����26��TO�ZDh�'����Ԍ�j���=��xX��d��`ɺ�Qպ�3�������JM��)�� ������*n��5%�!�*���0��z6��7<�%�A���G�;cM��S�O�X�)�^�(:d���i�l�o�.Vu��
{�L_��R9����c�ɋ�Ф��݀���]���:��=���  �  ā=�%=��=m=�=��=�V=�� =� =T> =���<%�<(G�<{��<��<G�<�L�<3��<��<	�<2F�<i��<���<���<�0�<�h�<y��<���<��<�;�<�l�<Ü�<���<���<z"�<�K�<�r�<��<N��<E��<��<Q�<1�<BH�<�\�<�m�<M|�<��<o��<��<֔�<��<u��<���<Vr�<q_�<=H�<�,�<G�<J��<g��<���<�Z�<d!�<���<��<�U�<�<ʲ�<�X�<u��<���<*�<��<�D�<�ɿ<�I�<�ļ<d:�<��<��<�}�<�<�=�<��<)�<�<�<؉�<�Ҫ<'�<�Y�<M��<�ӣ<��<�@�<>s�<&��<yК<���<�$�<�K�<�p�<ᓑ<���<�Ս<G�<��<�-�<�H�<#c�<s|�<�<�Y}<��y<��u<G�q<on<�>j<�kf<E�b<W�^<,�Z<�%W<�VS<�O<��K<�G<P)D<�b@<L�<<��8<�5<�a1<��-<��)<nB&<�"<F�<�G<X�<T<�y<s�<�a	<��<�b<���;���;�2�;uu�;<��;�+�;���;F'�;��;�l�;�,�;� �;�;��;���;�"�;Fa�;[��;�!�;{��;�;�;F�y;j`o;<e;��Z;�	Q;�DG;~�=;":4;��*;��!;��;�;jh;A��:Q�:u��:eW�:+b�:��:B0�:�:��}:!`:��B:<�%:�i	:Zt�9���9�5W9^g�8�ֵ�ظ�*V�t��_YӹSf�'�� 86��VO�UHh����7֌�����<��XX���c��1aɺ�Pպ�3��8����L��(�������H���l�o4%���*��0��y6��6<���A�"�G�YcM�S���X��^��9d���i�ܢo��Vu�M{��_��:��t���ʋ�w���T����]��1;��v���  �  ��=�%=x�=m=�=ų=�V=�� =� =V> =���<G�<0G�<���<9��<R�<�L�<X��<��<$	�<LF�<g��<���<���<�0�<�h�<X��<���<��<�;�<�l�<���<���<���<p"�<|K�<�r�<���<6��<5��<���<D�<�0�<%H�<u\�<�m�<N|�<���<x��<��<��<��<���<���<]r�<_�<OH�<�,�<^�<k��<f��<���<�Z�<g!�<��<��<�U�<��<���<�X�<f��<l��<�)�<��<�D�<�ɿ<�I�<�ļ<Z:�<骹<��<�}�<�ߴ<�=�<���<�<�<�<މ�<�Ҫ<E�<�Y�<g��<�ӣ<��<�@�<Os�</��<�К<���<�$�<�K�<�p�<ⓑ<���<�Ս<Z�<��<�-�<�H�<c�<]|�<ߔ�<�Y}<x�y<��u<�q<<n<w>j<�kf<1�b<,�^<��Z<�%W<�VS<܈O<i�K<��G<)D<�b@<\�<<��8<�5<�a1<)�-<��)<�B&<V�"<W�<
H<��<m<�y<��<�a	<�<c<���;: �;�2�;�u�;��;p+�;E��;�&�;P��;gl�;o,�; �;��;��;X��;k"�;�`�;��;Q!�;(��;�;�;��y;�_o;�e;��Z;�	Q;�EG;Ѫ=;�:4;��*;��!;��;y;�h;5��:r	�:��:�X�:Ld�:��:�1�:d�:��}:*!`:��B:��%:ag	:Fl�9_��9�.W9�S�8G�ڵ��ظn<V��u���_ӹ�g����<6�gXO��Jh����r׌�	���>��,Y��c���`ɺ�Nպ�3��	�5���vL��'�q��P������l�84%���*�%�0��y6�6<���A���G��bM��S���X���^�x:d�Y�i� �o��Wu��{�`��j:������:ʋ�̥������,^���;������  �  ��=�%=��=m=�=��=�V=�� =� =b> =���<O�<>G�<���<f��<_�<�L�<W��<6��</	�<VF�<r��<���<���<�0�<�h�<j��<���<��<�;�<�l�<���<���<u��<S"�<iK�<�r�<���<%��<.��<���<:�<
1�<.H�<�\�<�m�<L|�<���<o��<���<��<+��<���<��<kr�<�_�<uH�<�,�<r�<f��<���<���<�Z�<e!�<���<��<�U�<�<���<�X�<_��<_��<�)�<��<�D�<�ɿ<�I�<�ļ<>:�<骹<��<�}�<�ߴ<�=�<
��<�<�<�<Љ�<�Ҫ<*�<�Y�<q��<�ӣ<��<�@�<_s�<;��<�К<���<�$�<�K�<�p�<���<���<�Ս<I�<��<�-�<�H�<c�<e|�<攀<�Y}<b�y<y�u<��q<6n<3>j<bkf<�b<�^<��Z<�%W<|VS<��O<v�K<��G<9)D<�b@<K�<<��8<�5<�a1<2�-<�)<�B&<f�"<u�<3H<�<�<�y<��<�a	<)�<2c<���;���;�2�;vu�;>��;�+�;r��;'�;��;Tl�;,�; �;��;'�;��;�!�;�`�;µ�;:!�;���;�;�;�y;�_o;$e;��Z;�	Q;�DG;��=;;4;��*;��!;��;; i;c��:��:Ð�:-Z�:d�:��:�1�:E��:K�}:-`:��B:��%:ki	:-o�9²�9�+W9hG�8�۵\ٸ�9V�i~��eeӹ�k�w��m<6�s[O�|Kh�N���r׌�O���=��NX���c���`ɺbPպ73�	������K��'�������)���k��3%�(�*�Ϲ0� y6��5<�4�A��G��bM�-S���X�e�^�;:d��i���o�#Xu�?{�P`��w:������ʋ��け�y^���;������  �  ��=�%={�=m=�=γ=�V=�� =� =e> =���<S�<XG�<���<O��<\�<�L�<S��<F��<*	�<FF�<���<���<���<�0�<�h�<Z��<���<��<�;�<�l�<���<���<g��<V"�<�K�<�r�<���<��<.��<���<5�<�0�<H�<\�<�m�<h|�<���<���<��<ڔ�<C��<���<��<rr�<�_�<_H�<�,�<��<a��<���<���<�Z�<~!�<���<1��<�U�<��<���<�X�<X��<c��<�)�<��<�D�<�ɿ<�I�<�ļ</:�<�<��<�}�<�ߴ<�=�<�< �<�<�<҉�<�Ҫ<7�<Z�<e��<�ӣ<��<�@�<vs�<9��<�К<���<�$�<�K�<�p�<��<���<�Ս<\�<��<�-�<�H�<c�<I|�<۔�<�Y}<�y<y�u<��q<.n< >j<�kf<�b<�^<��Z<�%W<�VS<��O<e�K<��G< )D<�b@<c�<<��8<�5<�a1<�-<�)<�B&<n�"<��<%H<��<�<�y<��<�a	< �<c<#��;	 �;a3�;�u�;0��;+�;	��;�&�;
��;�l�;�+�;% �;r�;1�;���;�!�;�`�;���;:!�;��;s;�;��y;_o;�e;y�Z;�
Q;uEG;C�=;X;4;��*;��!;��;�;Vi;9��:~
�:��:Q[�:�c�:���:�0�:d��:p�}:�`:��B:��%:�h	:�h�9㭢9�(W9�K�8/۵Uٸ17V�B����^ӹ�j�Q���;6��\O�GJh�0����׌����?���X���c���^ɺ�Oպ�1��	�����J��'�2�����֠�l�3%��*�޹0��x6��6<���A�}�G�DbM��S��X���^�;d�w�i�ңo��Wu�>{�i`���:��;��V�ʋ�
�����^���;������  �  ��=�%=��=m=�=��=�V=�� =� =b> =���<O�<>G�<���<f��<_�<�L�<W��<6��</	�<VF�<r��<���<���<�0�<�h�<j��<���<��<�;�<�l�<���<���<u��<S"�<iK�<�r�<���<%��<.��<���<:�<
1�<.H�<�\�<�m�<L|�<���<o��<���<��<+��<���<��<kr�<�_�<uH�<�,�<r�<f��<���<���<�Z�<e!�<���<��<�U�<�<���<�X�<_��<_��<�)�<��<�D�<�ɿ<�I�<�ļ<>:�<骹<��<�}�<�ߴ<�=�<
��<�<�<�<Љ�<�Ҫ<*�<�Y�<q��<�ӣ<��<�@�<_s�<;��<�К<���<�$�<�K�<�p�<���<���<�Ս<I�<��<�-�<�H�<c�<e|�<攀<�Y}<b�y<y�u<��q<6n<3>j<bkf<�b<�^<��Z<�%W<|VS<��O<v�K<��G<9)D<�b@<K�<<��8<�5<�a1<2�-<�)<�B&<f�"<u�<3H<�<�<�y<��<�a	<)�<2c<���;���;�2�;vu�;>��;�+�;r��;'�;��;Tl�;,�; �;��;'�;��;�!�;�`�;µ�;9!�;���;�;�;�y;�_o;$e;��Z;�	Q;�DG;��=;;4;��*;��!;��;; i;c��:��:Ð�:-Z�:d�:��:�1�:E��:K�}:-`:��B:��%:ki	:-o�9²�9�+W9hG�8�۵\ٸ�9V�i~��eeӹ�k�w��m<6�s[O�|Kh�N���r׌�O���=��NX���c���`ɺbPպ73�	������K��'�������)���k��3%�(�*�Ϲ0� y6��5<�4�A��G��bM�-S���X�e�^�;:d��i���o�#Xu�?{�P`��w:������ʋ��け�y^���;������  �  ��=�%=x�=m=�=ų=�V=�� =� =V> =���<G�<0G�<���<9��<R�<�L�<X��<��<$	�<LF�<g��<���<���<�0�<�h�<X��<���<��<�;�<�l�<���<���<���<p"�<|K�<�r�<���<6��<5��<���<D�<�0�<%H�<u\�<�m�<N|�<���<x��<��<��<��<���<���<]r�<_�<OH�<�,�<^�<k��<f��<���<�Z�<g!�<��<��<�U�<��<���<�X�<f��<l��<�)�<��<�D�<�ɿ<�I�<�ļ<Z:�<骹<��<�}�<�ߴ<�=�<���<�<�<�<މ�<�Ҫ<E�<�Y�<g��<�ӣ<��<�@�<Os�</��<�К<���<�$�<�K�<�p�<ⓑ<���<�Ս<Z�<��<�-�<�H�<c�<]|�<ߔ�<�Y}<x�y<��u<�q<<n<w>j<�kf<1�b<,�^<��Z<�%W<�VS<܈O<i�K<��G<)D<�b@<\�<<��8<�5<�a1<)�-<��)<�B&<V�"<W�<
H<��<m<�y<��<�a	<�<c<���;: �;�2�;�u�;��;p+�;E��;�&�;P��;gl�;o,�; �;��;��;X��;j"�;�`�;��;Q!�;(��;�;�;��y;�_o;�e;��Z;�	Q;�EG;Ѫ=;�:4;��*;��!;��;y;�h;5��:r	�:��:�X�:Ld�:��:�1�:d�:��}:*!`:��B:��%:ag	:Fl�9_��9�.W9�S�8G�ڵ��ظn<V��u���_ӹ�g����<6�gXO��Jh����r׌�	���>��,Y��c���`ɺ�Nպ�3��	�5���vL��'�q��P������l�84%���*�%�0��y6�6<���A���G��bM��S���X���^�x:d�Y�i� �o��Wu��{�`��j:������:ʋ�̥������,^���;������  �  ā=�%=��=m=�=��=�V=�� =� =T> =���<%�<(G�<{��<��<G�<�L�<3��<��<	�<2F�<i��<���<���<�0�<�h�<y��<���<��<�;�<�l�<Ü�<���<���<z"�<�K�<�r�<��<N��<E��<��<Q�<1�<BH�<�\�<�m�<M|�<��<o��<��<֔�<��<u��<���<Vr�<q_�<=H�<�,�<G�<J��<g��<���<�Z�<d!�<���<��<�U�<�<ʲ�<�X�<u��<���<*�<��<�D�<�ɿ<�I�<�ļ<d:�<��<��<�}�<�<�=�<��<)�<�<�<؉�<�Ҫ<'�<�Y�<M��<�ӣ<��<�@�<>s�<&��<yК<���<�$�<�K�<�p�<ᓑ<���<�Ս<G�<��<�-�<�H�<#c�<s|�<�<�Y}<��y<��u<G�q<on<�>j<�kf<E�b<W�^<,�Z<�%W<�VS<�O<��K<�G<P)D<�b@<L�<<��8<�5<�a1<��-<��)<nB&<�"<G�<�G<X�<T<�y<s�<�a	<��<�b<���;���;�2�;tu�;<��;�+�;���;F'�;��;�l�;�,�;� �;�;��;���;�"�;Fa�;[��;�!�;{��;�;�;F�y;j`o;<e;��Z;�	Q;�DG;~�=;":4;��*;��!;��;�;jh;A��:Q�:u��:eW�:+b�:��:B0�:�:��}:!`:��B:<�%:�i	:Zt�9���9�5W9^g�8�ֵ�ظ�*V�t��_YӹSf�'�� 86��VO�UHh����7֌�����<��XX���c��1aɺ�Pպ�3��8����L��(�������H���l�o4%���*��0��y6��6<���A�"�G�YcM�S���X��^��9d���i�ܢo��Vu�M{��_��:��t���ʋ�w���T����]��1;��v���  �  ҁ=�%=��=m=�=��=�V=� =�� =I> =���<�<�F�<Q��<��<�<zL�<��<���<	�<F�<f��<���<���<�0�<�h�<o��<���<	�<�;�<m�<М�<$��<���<�"�<�K�<�r�<F��<`��<a��<��<c�<%1�<4H�<�\�<�m�<]|�<|��<h��<֓�<���<���<X��<̀�<%r�<U_�<%H�<t,�<2�<,��<S��<o��<{Z�<a!�<���<"��<�U�<�<���<�X�<���<���<%*�<.��<�D�<ʿ<J�<�ļ<�:�<;��<��<�}�< �<�=�<��<�<�<�<Ӊ�<�Ҫ<�<�Y�<9��<iӣ<��<�@�<s�<���<lК<���<u$�<nK�<}p�<ʓ�<b��<�Ս<:�<��<�-�<�H�< c�<g|�<��<�Y}<߈y<޶u<z�q<�n<�>j<lf<�b<��^<i�Z<&W<�VS<	�O<üK<��G<I)D<�b@<V�<<��8<y5<�a1<��-<��)<<B&<�"<��<�G<A�<�<<y<A�<^a	<��<�b<���;i��;�2�;`u�;#��;�+�;���;�'�;���;2m�;�,�;'�;��;6�;]��;�"�;�a�;���;�!�;ͣ�;<�;��y;�_o;$e;/�Z;P
Q;pDG;<�=;�94;��*;-�!;��;�;�f;s��:��:K��:�U�:>`�:���:^.�:E�:X�}:5`:��B:4�%:9i	:;p�9��9m@W9`|�8�yε�ظ�V��m���Oӹ�a�����26��TO�ZDh�'����Ԍ�j���=��xX��d��`ɺ�Qպ�3�������JM��)�� ������*n��5%�!�*���0��z6��7<�%�A���G�;cM��S�O�X�)�^�(:d���i�l�o�.Vu��
{�L_��R9����c�ɋ�Ф��݀���]���:��=���  �  ܁=�%=��=$m=�=��=�V=p� =� =:> =p��<��<�F�<0��<���<��<WL�<��<���<��<F�<G��<���<���<�0�<�h�<w��<���<	�<�;�<,m�<���<A��<���<�"�<�K�<s�<Z��<���<���<-��<y�<;1�<;H�<�\�<�m�<E|�<i��<R��<���<���<ӑ�<:��<���<r�<4_�<H�<Q,�<�<��<+��<^��<fZ�<G!�<���<
��<�U�<$�<Ų�<Y�<���<���<K*�<T��<�D�<Bʿ<<J�<ż<�:�<V��<�<~�<6�<�=�<4��<*�<=�<Ӊ�<�Ҫ<�<�Y�<'��<Vӣ<Y�<�@�<�r�<Ң�<GК<`��<S$�<RK�<Xp�<���<Q��<pՍ<.�<��<�-�<�H�<0c�<r|�<��<Z}<�y<1�u<��q<�n<?j<Glf<ҙb<��^<��Z<\&W<#WS<9�O<�K<�G<b)D<�b@<B�<<o�8<e5<Ua1<��-<i�)<�A&<��"<��<QG<��<�<�x<	�<a	<��<�b<��;B��;�2�;>u�;m��;�+�;Ġ�;�'�;���;{m�;n-�;��;"�;��;���;�#�;Bb�;��;�"�;��;j<�;l�y;`o;�e;��Z;�	Q;�CG;�=;�84;H�*;��!;��;;�e;R��:��:���: T�:�^�:��:6-�:��:��}:+`:Q�B:H�%:}l	:r�9o��9FKW9O��8��ŵ�ظL
V��c���Hӹ�]�����/6��OO�Ah�񄀺�ӌ�7�� =���V��,d���aɺ$Rպ�5������N�n*��F����5o��6%�	�*�ּ0��{6�L8<��A��G��cM�KS���X���^��9d�W�i���o��Uu�b	{��^���8��[���ȋ�i���R��� ]��|:������  �  �=�%=��="m=�=��=�V=g� =� =*> =T��<��<�F�<��<���<��<+L�<ڋ�<���<��<�E�<8��<|��<���<�0�<�h�<���<
��<,	�<�;�<Gm�<!��<_��<��<�"�<L�<Ds�<v��<���<���<O��<��<K1�<TH�<�\�<�m�<E|�<f��<L��<���<���<���<��<���<�q�<_�<�G�<3,�<��<���<��<B��<WZ�<A!�<���<
��<�U�<�<޲�<Y�<���<Ԕ�<e*�<���<E�<qʿ<iJ�<5ż<�:�<w��<8�<~�<]�<	>�<S��<;�<=�<؉�<�Ҫ<�<�Y�<��<8ӣ<@�<p@�<�r�<���<К<=��<0$�<&K�<<p�<���<;��<_Ս<%�<��<�-�<�H�<-c�<�|�<+��<NZ}<F�y<b�u<�q<5n<p?j<�lf<1�b<$�^<��Z<�&W<bWS<t�O<�K<U�G<h)D<�b@<D�<<Z�8<W5<3a1<j�-<(�)<�A&<V�"<R�<G<��<i<�x<��<�`	<K�<\b<���;��;V2�;<u�;N��;�+�;0��;(�;y��;�m�;�-�;��;��;h�;O��;($�;�b�;���;�"�;���;�<�;��y;�`o;qe;s�Z;{	Q;�CG;C�=;c84;f�*;�!;�;�;�d;���:��:��:Q�:�\�:���:b+�:��:��}:�`:��B:7�%:!k	:ww�9�¢9�SW9 ��8���}ظp�U��X���>ӹ�W�{��B,6��JO�>h������Ҍ�t��"<��jW��d��+bɺ�Rպ�6�����O��+�o�+��w��Sp�8%�e�*���0��|6��8<���A�0�G�dM�FS���X���^��8d���i�ڠo��Tu��{�<^��~8�����z툻Bȋ�棎�����\��:��n���  �  �=�%=��=!m=�=��=�V=b� =ڛ => =5��<��<�F�<��<���<��<L�<���<���<��<�E�<+��<]��<���<�0�<�h�<���<��<;	�<<�<fm�<=��<���<#��<#�<3L�<`s�<���<λ�<���<m��<��<X1�<\H�<�\�<�m�<O|�<W��<2��<���<i��<���<���<d��<�q�<�^�<�G�<,�<��<���<���<!��<HZ�<-!�<���<��<�U�<"�<��<(Y�<���<���<*�<���<RE�<�ʿ<�J�<`ż<�:�<���<W�<=~�<z�<>�<\��<B�<=�<܉�<�Ҫ<��<�Y�<��<ӣ<-�<K@�<�r�<���<�Ϛ<��<$�<K�<p�<o��<��<SՍ<�<��<�-�<�H�<6c�<�|�<;��<sZ}<��y<��u<U�q<�n<�?j<�lf<r�b<y�^<G�Z<�&W<�WS<��O<&�K<c�G<|)D<�b@<N�<<Q�8<5<a1<,�-<��)<tA&<�"<�<�F<<�<<Yx<n�<�`	<�<!b<��;���;X2�;9u�;@��;,�;F��;7(�;���;Ln�;Z.�;��;-�;��;	��;�$�;Zc�;:��;1#�;��;�<�;7�y; ao;�e;Y�Z;�	Q;&CG;g�=;�74;@�*;V�!;��;�;gc;��:��::��:0O�:�Y�:%��:2)�:��:�}:=`:A�B:(�%:�k	:�x�9�Ģ9�\W9���84`��_\ظw�U�
Q��,3ӹS�p��v&6�oGO�u:h�����ь�
���;��sW���c���aɺNTպy7ẙ�.���%P��,�Q��������q�;9%�^�*�ξ0�u}6�:<���A�%�G�]dM�S���X�x�^��8d�x�i�G�o��Su��{��]���7��#���숻�ǋ�>���)��\��9�����  �  ��=�%=��=&m=}=��=�V=X� =Λ => =��<��<tF�<���<~��<�<�K�<���<u��<��<�E�<��<S��<���<�0�<�h�<���<"��<X	�<<�<�m�<`��<���<F��<4#�<YL�<�s�<Ř�<��<���<���<��<x1�<gH�<�\�<�m�<5|�<N��<��<���<W��<���<ϊ�<O��<�q�<�^�<�G�<�+�<��<���<߼�<��<4Z�<!�<���<���<�U�<?�<���<GY�<���<��<�*�<º�<sE�<�ʿ<�J�<�ż<$;�<ɫ�<{�<e~�<��<:>�<s��<X�<)=�<ω�<�Ҫ<��<�Y�<<ӣ<�<)@�<�r�<a��<�Ϛ<���<�#�<�J�<�o�<[��<��<?Ս<��<x�<�-�<�H�<Lc�<�|�<Z��<�Z}<��y<�u<��q<�n<�?j<Cmf<��b<��^<{�Z<'W<�WS<ȉO<g�K<w�G<�)D<�b@<%�<<<�8<�5<�`1<��-<��)<A&<ӓ"<��<YF<�<�<)x<!�<?`	<��<�a<%��;e��;
2�;�t�;x��;B,�;v��;�(�;���;�n�;�.�;�;��;q�;���;#%�;�c�;���;�#�;Q��;:=�;&�y;Iao;be;G�Z;�Q;�BG;��=;074;��*;d�!;y�;�;=b;׼�:5��:Ԃ�:�M�:�W�:��:(�:X�:<�}:;`:��B:U�%:�n	::|�96̢9\gW9��8ݯ��BظI�U��G��8*ӹ�N����"6�cCO��5h����Ќ�����:��V���d���bɺ�Tպ�8���m���gQ��-������v���r�):%�Q�*�$�0�~6��:<���A���G��dM��S���X�Ń^�o8d��i���o��Ru�z{�4]��C7�����숻Aǋ������~���[��
9������  �  ��=�%=��=$m=�=��=�V=K� =Ǜ => =���<l�<KF�<���<X��<c�<�K�<}��<_��<�<�E�<���<a��<���<�0�<�h�<���<-��<a	�<><�<�m�<|��<���<u��<X#�<hL�<�s�<��<��<���<���<��<y1�<rH�<�\�<�m�<8|�<\��<��<v��<G��<e��<Ê�<$��<xq�<�^�<nG�<�+�<��<���<���<���<Z�<!�<���<��<�U�</�< ��<MY�<���<*��<�*�<��<�E�<�ʿ<�J�<�ż<W;�<߫�<��<}~�<��<G>�<~��<\�<=�<ቬ<�Ҫ< �<�Y�<���<�ң<�
�<@�<vr�<G��<�Ϛ<���<�#�<�J�<�o�<<��<���<(Ս<��<�<�-�<�H�<=c�<�|�<^��<�Z}<�y<�u<��q<"n<O@j<Wmf<�b<�^<��Z<O'W<XS<��O<p�K<��G<�)D<�b@<3�<<G�8<
5<�`1<�-<��)<�@&<��"<}�<F<��<v<�w<��<`	<��<�a<���;���;2�;u�;B��;1,�;���;�(�;{��;o�;B/�;O�;c�;��;���;�%�;=d�;���;$�;���;�=�;!�y;�ao;�e;��Z;�Q;8CG;��=;�64;�*;^�!;�;�
;;a;���:���:��:K�:�V�:��:�&�:��:�}:+`:J�B:G�%:�l	:I~�9͢9�nW9���8e����$ظ��U�A;���$ӹ�J���e 6��?O�&3h�~��nό�D���:��W���c���bɺ�Sպ:�������7R�q.�l��������s�d;%�l�*���0�6�$;<�O�A���G�]dM��S���X�9�^��7d�c�i��o�Ru��{��\���6������눻�Ƌ�
���v~��&[���8��`���  �  ��=�%=��=)m=~=��=�V=B� =Û =�= =��<P�<9F�<���<7��<^�<�K�<d��<O��<d�<�E�<��<H��<���<�0�<�h�<���<=��<i	�<T<�<�m�<���<���<|��<e#�<L�<�s�<���<*��<���<���<��<w1�<�H�<�\�<n�<)|�<;��<��<d��<6��<R��<���< ��<rq�<�^�<YG�<�+�<h�<���<���<��<Z�<� �<���<��<�U�<4�<"��<PY�<��<@��<�*�<
��<�E�<�ʿ<�J�<�ż<a;�<���<��<~~�<��<V>�<���<{�<=�<艬<�Ҫ<��<�Y�<՗�<�ң<�
�< @�<Xr�<A��<�Ϛ<���<�#�<�J�<�o�<#��<鴏<Ս<��<^�<�-�<I�<Kc�<�|�<^��<�Z}<��y<:�u< �q<9n<i@j<�mf<)�b<(�^<��Z<y'W<XS<0�O<y�K<��G<�)D<�b@<*�<<	�8<�5<�`1<ϧ-<S�)<�@&<X�"<V�<F<v�<i<�w<��<�_	<n�<�a<e��;,��;�1�;u�;E��;�,�;ԡ�;�(�;���;o�;�/�;��;z�;$�;"��;�%�;�d�;���;0$�;���;�=�;�y;�bo;�e;��Z;lQ;#BG;̦=;�54;��*;��!;~�;]	;a;���:w��:���:�H�:LU�:؞�:�%�:�:F�}:`:.�B:��%:3m	:]��9q͢9zW9v�8-!����׸m�U��9�� ӹCI����6�X<O�M3h��|���Ό�|���8���V���c��Vdɺ�Uպ_;Ặ�J����R�4/�`�������;t��;%�i +��0��6��;<���A�<�G�beM��S�`�X�ʃ^��6d�b�i��o��Qu�E{�I\��{6�����{눻[Ƌ�衎��}���Z���8������  �  �=�%=��=$m=�=��=�V=E� =�� =�= =ֿ�<I�<-F�<s��<$��<;�<�K�<V��<C��<Y�<�E�<��<P��<���<�0�<�h�<���</��<y	�<S<�<�m�<���<���<���<�#�<�L�<�s�<��<%��<��<���<��<1�<zH�<�\�<�m�<8|�<J��<��<b��<$��<N��<���<��<Uq�<q^�<?G�<�+�<n�<s��<���<ߍ�<Z�<	!�<���<��<�U�<6�<��<RY�<��<@��<�*�<��<�E�<˿<K�<�ż<p;�<��<��<�~�<��<f>�<���<i�<=�<މ�<�Ҫ<��<�Y�<ʗ�<�ң<�
�<�?�<[r�<��<�Ϛ<���<�#�<�J�<�o�<��<Դ�<Ս<��<q�<�-�<�H�<Fc�<�|�<j��<[}<�y<f�u<�q<Xn<�@j<�mf<N�b<E�^<��Z<�'W<@XS<<�O<��K<��G<�)D<�b@<3�<<.�8<�5<�`1<��-<C�)<�@&<H�"<?�<�E<N�<"<�w<��<�_	<V�<�a<~��;G��;�1�;�t�;,��;S,�;���;)�;���;o�;�/�;��;��;��;���;$&�;�d�;|��;�$�;���;>�;B�y;�ao;�e;C�Z;�Q;�BG;)�=;�54;��*;��!;��;v	;`;���:���:�~�:)I�:T�:���:�$�:��:�}:�`:*�B:��%:Bm	:<��9�͢9��W9��8����ظ��U�W6��ӹ,E�N��t6��;O�~/h��|���͌�3���9��W��<d��KcɺUպ�:�t����S��/�N���8��$u�_<%�� +���0� �6�.<<���A���G��dM��S���X��^��7d���i�ϝo�\Qu��{�E\��>6��}���ꈻƋ������}���Z��P8������  �  %�=g(=��=vp=0=��=[=7� =� =�C =V��<��<�T�<͗�<���<��<?^�<��<:��<��<]�<���<R��<�<�M�<,��<u��<���<P,�<�`�<���<��<��<#�<$P�<{�<��<I��<:��<?�<�3�<R�<�m�<���<���<1��<t��<���<W��<���<z��<���<���<#��<<��<V��<��<Ȅ�<Ef�<�B�<��<���<O��<P��<�D�<��<Z��<8k�<+�<���<!^�<���<$��<r�<d��<�+�<|��<�#�<"��<'�<q�<7ֶ<H6�<�<��<�;�<�<(Ԭ<��<]�<0��<�ץ<)�<zE�<�w�<���<�Ԝ<d��<�'�<�M�<Nr�<���<���<�ԏ<D�<k�<^)�<"C�<�[�<�s�<p��<���<l}<�y<5�u<��q<�n<�7j<&`f<c�b<q�^<��Z<�W<*1S<�]O<R�K<+�G<�C<�!@<�W<<��8<��4<t
1<�K-<_�)<G�%<l'"<�x<&�<�*<Ҋ<�<�\<
�<�G<��<��;���;���;��;_c�;���;�+�;ժ�;J<�;4��;��;+i�;3L�;�D�;S�;�w�;N��;�;�n�;l�;��;;iv;��k;a�a; �W;��M;��C;S:;��0;�';��;W�;�;�O;;��:��:˹�:���:Ӷ:B�:3�:�ψ:��s:�xV:�9:^�:{� :��9Qi�9z�79o��8���r��EOq�����w�߹�s	��"�/�;��T�erm�?���9���^���s���w���o���X˺�5׺<������n�x��������fL�� ���%�F�+�C1���6�g�<��^B��H�&�M�imS��Y���^��td�O!j���o�X{u�F({�2k���A��L��g����ȋ�Ơ���y��S���-���	���  �  �=b(=�=tp=9=Ƿ=[=8� =� =�C =[��<��<�T�<Η�<���<��<F^�<��<6��<��<]�<���<g��<�<�M�<!��<g��<r��<?,�<�`�<���<#��<#��<|#�<*P�<{�< ��<D��<F��<.�<�3�<�Q�<�m�<���<֜�<3��<���<���<d��<���<x��<���<���<+��<V��<<��<͞�<���<Jf�<�B�<q�<���<V��<Y��<�D�<��<^��<k�<,�<}��<^�<���<��<|�<^��<�+�<���<�#�<��<'�<q�< ֶ<T6�<味<��<};�<���<6Ԭ<��</]�<3��<�ץ< �<qE�<�w�<���<�Ԝ<<��<�'�<N�<Vr�<Ɣ�<���<�ԏ<G�<~�<v)�<2C�<�[�<�s�<h��<���<l}<��y<'�u<��q<�n<�7j<!`f<t�b<q�^<�Z<�W<1S<�]O</�K<�G<��C<�!@<X<<��8<�4<v
1<L-<E�)<Q�%<{'"<y<)�<e*<�<�<�\<�<tG<��<��;��;7��;�;3c�;j��;D+�;���;n<�;���;4��;?i�;)L�;�D�;.S�;�w�;=��;5�;ln�;��;���;�hv;��k;\�a;.�W;)�M;_�C;yS:;
�0;�';]�;��;[�;�P;���:��:F��:��:�Ӷ:A�:��:Ј:��s:?{V:#�9:��:ު :r��9d�9��79۪�8n��Y���Qq�}���,�߹s	�V�"��;���T�Cum�y���:��&`��Pt��y���n��yW˺r4׺�I��w�����#�����T���M� �]�%��+��B1�!�6��<��^B�[H�e�M��lS��Y�n�^�ud��!j�m�o��{u�~({��j���A��%��q����ȋ�Ǡ���y���S��.��{	���  �  �=l(=��=wp=3=��=[=9� =&� =�C =y��<��<�T�<���<���<��<O^�<.��<O��<��<.]�<���<h��<�<�M�< ��<w��<��<,,�<�`�<���<��<��<b#�<P�<�z�<��<��<8��<�<�3�<�Q�<�m�<���<ל�<?��<u��<���<a��<���<���<���<���<.��<w��<^��<��<��<Kf�<�B�<��<��<g��<V��<�D�<��<g��<k�<F�<x��<^�<���<��<r�<7��<�+�<\��<�#�<��<�<q�< ֶ<Q6�<ё�<��<�;�<܉�<2Ԭ<��<-]�<3��<�ץ<2�<�E�<�w�<���<�Ԝ<^��<�'�<N�<_r�<攓<���<�ԏ<M�<�<j)�<'C�<�[�<�s�<~��<y��<l}<ٕy<��u<��q<�n<�7j<�_f<T�b<,�^<��Z<\W<�0S<�]O<�K<?�G<��C<�!@<�W<<��8<�4<z
1<IL-<]�)<��%<�'"<,y<}�<�*<:�<'�<"]<6�<�G<��<��;��;���; �;6c�;���;+�;L��;o<�;t��;��;�h�;�K�;YD�;�R�;�w�;���;�;�m�;q�;���;ehv;��k;r�a;��W;��M;�C;hS:;y�0;ޭ';��;��;}�;�Q;Ϸ�:��:ӽ�:3��:�ն:rB�:j�:9ш:��s:�zV:�9:0�:�� :&��9c�9I�79Ѧ�85���u���dq�������߹]v	���"�1�;�t�T� ym�����;���_��&s��4y��o���X˺q4׺�����Q�����-��\�����L�� ���%���+��A1���6�3�<��^B�UH�˾M�HmS��Y�/�^�ntd�V"j���o�|u�,){�Sk��fB��c����ȋ�P���0z���S��h.���	���  �  �=[(=z�=vp=6=ȷ=%[=C� =)� =�C =���<��<�T�<��<���<��<p^�<H��<c��<��<0]�<Ϛ�<��<�<�M�<!��<W��<i��<,�<�`�<z��<���<���<O#�<�O�<�z�<���<��<��<�<�3�<�Q�<�m�<���<Ҝ�<=��<{��<���<t��<���<���<���<��<P��<��<x��<��<��<mf�<C�<��< ��<o��<j��<�D�<��<e��<k�<�<j��<�]�<���<ߍ�<T�<��<v+�<>��<�#�<<��<�p�<�ն<16�<���<��<f;�<ډ�<4Ԭ<��<C]�<G��<�ץ<I�<�E�<x�<���<�Ԝ<��<�'�<-N�<�r�<���<���<�ԏ<^�<��<~)�<,C�<�[�<~s�<W��<n��<�k}<��y<׾u<K�q<mn<�7j<�_f<�b<��^<��Z<2W<�0S<�]O<�K<��G<��C<�!@<�W<<��8<<�4<�
1<UL-<��)<��%<�'"<fy<��<�*<U�<m�<Z]<a�<�G<��<Q��;V��;5��;�;Ac�;8��;1+�;��;<�;O��;���;Yh�;�K�;�C�;AR�;/w�;C��;��;�m�;�;{��;"hv;�k;P�a;��W;�M;��C;
T:;��0;^�';Ś;Y�;��;R;���:��:7��:^��:L׶:D�:��:�ш:�s:�}V:��9:3�:�� :f��9&`�9��795��8C�����qq�������߹�y	���"���;��T�]zm�c���<���`���u��1y���n���W˺�2׺�㺞��Ă��L�t��F������K�4 ��%���+�hA1���6���<�^B��H�*�M�mS��Y���^��ud��"j�w�o��|u��){��k���B�����g�2ɋ������z��T���.���	���  �  
�=T(={�=sp=9=η=$[=M� =5� =�C =���<�<�T�<-��<���<�<�^�<e��<���<��<G]�<��<|��<(�<�M�<!��<U��<[��<,�<d`�<U��<���<���<#�<�O�<�z�<���<���<���<��<~3�<�Q�<m�<���<ڜ�</��<���<���<}��<���<���<���<��<���<���<���<:��<9��<�f�<C�<��<=��<���<s��<�D�<��<V��<k�<�<Y��<�]�<���<���<&�<���<:+�<��<�#�<���<��<�p�<�ն<6�<���<��<b;�<ۉ�<(Ԭ<��<=]�<T��<�ץ<p�<�E�<x�<觞<�Ԝ<���<
(�<bN�<�r�<��<ٵ�<�ԏ<r�<��<�)�<6C�<�[�<�s�<J��<g��<�k}<l�y<�u<�q<+n<7j<P_f<��b<��^<^�Z<�W<v0S<f]O<�K<ݻG<��C<�!@<X<<Ґ8<9�4<�
1<�L-<��)<��%<2("<�y<��<P+<��<��<�]<��<.H<*�<���;U��;���;�;Qc�;=��;+�;��;�;�;���;���;�g�;�J�;C�;�Q�;Mv�;б�;�;Bm�;��;��;�gv;��k;��a;/�W;c�M;�C;^T:;��0;Q�';�;��;��;�S;k��:��:��:Z��:�ض:IF�:��:$ӈ:��s: ~V:��9:��:W� :ԃ�9�\�9%�79�i�8��������q����2๣�	�l�"�?�;�G�T��~m�U���=���a���u���x��To���V˺/3׺��?��4���G����i��{��J�� �v�%��+��@1�a�6�$�<�{]B��H��M��lS��Y�x�^�vd��"j�w�o��}u�+{�6l��NC������ʋ�K���{���T��9/��}
���  �  ��=N(=u�=lp=;=ӷ=1[=\� =F� =�C =���<4�<U�<f��<-��<G�<�^�<���<���<��<j]�<���<���<5�<�M�<��<P��<D��<�+�<V`�<6��<���<���<�"�<�O�<�z�<���<���<���<��<n3�<�Q�<\m�<���<Ɯ�<,��<���<���<���<
��<���<��<O��<���<���<״�<i��<k��<�f�<IC�<��<W��<���<���<E�<
�<S��<k�<	�<6��<�]�<���<���<��<Ǧ�<+�<ݩ�<V#�<���<��<�p�<�ն<�5�<���<��<[;�<É�<&Ԭ<��<P]�<q��<إ<��<�E�<Mx�< ��<!՜<���<A(�<�N�<�r�<@��<���<�ԏ<��<��<�)�<?C�<�[�<ts�<D��<A��<gk}<D�y<%�u<��q<�n<�6j<�^f<\�b<H�^<��Z<�W<E0S<>]O<��K<ŻG<��C<�!@<X<<�8<m�4<1<�L-<)�)<K�%<~("<z<f�<�+<�<�<�]<�<`H<v�<+��;���;���;%�;c�;7��;�*�;e��;o;�;W��;r��;Cg�;J�;�B�;�P�;�u�;*��;X�;�l�;\�;���;�fv;��k;�a;-�W;�M;R�C;qU:;��0;O�';L�;��;X�;U;���:��:L��:��:�۶:�H�:m�:6Ո:p�s:cV:߅9:��:˨ :���9�T�9��79�Z�8Z��9��{�q������p�	���"� �;���T�h�m�"	��,@��yc���u��;z��Io���U˺�1׺� �3���~����*���������H�, �a�%�-�+�?1���6��<�y\B��H���M��lS�;Y���^�?vd�$j�2�o�d~u��,{�m��D��M���򈻰ʋ�����{��xU���/���
���  �  �=F(=n�=pp=>=׷=>[=d� =Z� =D =��<j�<HU�<���<N��<��<�^�<͟�<���<�<�]�<��<���<3�<�M�<��<?��<5��<�+�<)`�<��<���<g��<�"�<iO�<Bz�<g��<���<���<��<93�<�Q�<Gm�<n��<���<7��<���<���<���<��<��<&��<���<���<��<��<���<���<�f�<C�<�<��<���<���<E�< �<Z��<�j�<��< ��<�]�<X��<]��<��<���<�*�<���<#�<R��<X�<hp�<oն<�5�<c��<��<B;�<���<0Ԭ<��<c]�<|��<5إ<��<F�<�x�<4��<]՜<���<x(�<�N�<s�<t��<��<&Տ<��<��<�)�<BC�<�[�<is�<0��<(��<%k}<��y<�u<V�q<an<s6j<e^f<��b<�^<��Z<<W<�/S<�\O<a�K<��G<��C<�!@<X<<��8<��4<)1<M-<k�)<��%<�("<�z<��<�+<��<��<s^<\�<�H<��<m��;.��;���;f�;3c�;��;�*�;��;�:�;���;���;�f�;fI�;�A�; P�;u�;]��;��;	l�;��;D��;8fv;V�k;�a;��W;ۧM;��C;#V:;K�0;��';"�;l�;��;�V;���:;!�:��:��:F߶:�J�:��:�ֈ:��s:�V:�9:��:� :f~�9P�9h�79�&�8��������q������"�^�	���"���;�M�T�P�m�1���A��cd��w��,z��un��UV˺y0׺���?��m|����f����ƀ��G�p	 ���%���+��=1���6�ݨ<�\B��H�L�M�rlS��Y�J�^��vd��$j�7�o��u��-{��m���D�� ����lˋ�ѣ���|�� V��Y0��T���  �  �=8(=k�=lp=;=޷=G[=q� =l� = D ='��<��<yU�<ј�<���<��<._�<���<���<N�<�]�<%��<���<=�<�M�<��<1��<��<�+�<`�<��<P��<5��<�"�<3O�<z�<*��<M��<g��<m�<3�<eQ�<7m�<X��<Ɯ�<+��<���<���<���<7��<8��<R��<���<
��<D��<=��<̟�<Ӆ�<'g�<�C�<)�<���<Ϻ�<���<.E�<�<M��<�j�<��<
��<y]�<+��<=��<��<Z��<�*�<p��<�"�<��<$�<+p�<Sն<�5�<N��<r�<-;�<���<!Ԭ<��<v]�<���<Sإ<��<(F�<�x�<i��<�՜<< �<�(�<�N�<5s�<���<B��<QՏ<��<��<�)�<>C�<�[�<is�<��<��<�j}<��y<��u<��q<�n<�5j<!^f<��b<v�^<0�Z<�W<�/S<�\O<B�K<h�G<��C<�!@<X<<�8<��4<]1<gM-<͒)<��%<K)"<�z<D�<�,<��<��<�^<��<I<�<ߛ�;���;��;P�;9c�;ܽ�;A*�;��;;:�;H��;0��;�e�;�H�;
A�;�O�;.t�;���;��;�k�;�;؃�;�ev;��k;6�a;C�W;�M;��C;�V:;+�0;8�';��;��;��;iX;:��: %�:��:r��:��:BM�:=��:f؈:�s:�V:ǅ9:��:�� :Cy�9�K�9�t79���8�g���	�,�q��Ĭ�?,๊�	�?�"���;�c�T�^�m�����B���e��0x��$z��)o���U˺/׺d��<��y����-��@��^��E�� ��%��+�o<1��6���<�4[B�~H�ȼM��lS�TY�Q�^��wd�I%j�N�o��u��.{��n���E�����b�]̋�����i}���V���0������  �  ԃ=,(=g�=kp=B=�=N[=�� =u� =-D =P��<��<�U�<���<���<��<]_�<)��<&��<^�<�]�<K��<���<N�<�M�<��<)��<���<�+�<�_�<͒�<��<��<`"�<�N�<�y�<��<2��<4��<=�<�2�<EQ�<m�<D��<���<*��<���<���<���<[��<D��<x��<���<7��<o��<d��<���<���<Rg�<�C�<R�<���<��<̂�<+E�<�<J��<�j�<��<��<U]�<��<��<X�<:��<a*�<=��<�"�<喻<�<�o�<+ն<y5�<(��<M�<";�<���<"Ԭ<��<t]�<���<jإ<��<VF�<�x�<���<�՜<j �<�(�<O�<es�<���<`��<_Տ<��<��<�)�<OC�<�[�<]s�< ��<���<�j}<j�y</�u<��q<�n<�5j<�]f<�b<7�^<��Z<yW<l/S<c\O<�K<7�G<w�C<�!@<*X<<#�8<��4<�1<�M-<�)<I�%<�)"<Q{<��<�,<L�<`�<7_<�<EI<=�<���;���;S��;}�; c�;ƽ�;�)�;k��;�9�;���;q��;ge�;H�;:@�;�N�;Vs�;>��;4�;�j�;��;`��;�dv;0�k;��a;M�W;��M;��C;�W:;Z�0;��';Р;׶;�;�Y;���:�'�:���:H��:h�:�O�:(��:�ڈ:��s:��V:]�9:��:�� :�u�9�C�9ld79N�8x���,	���q�Ҭ�8��	���"��;���T�֐m����E���g���x���z���n���T˺/׺ �⺩��1x��8����ڳ�+~�	D�� ���%���+�7;1�.�6��<�ZB��H���M�lS�[Y���^�exd�5&j�d�o�ǁu�R0{�Ao��)F��������D͋�'���	~��}W��?1��s���  �  ʃ=-(=`�=ip=D=�=U[=�� =�� =AD =}��<��<�U�<0��<���<�<|_�<G��<Q��<��<�]�<R��<���<H�<�M�<���<#��<���<�+�<�_�<���<��<���<+"�<�N�<�y�<ʢ�<���<��<�<�2�</Q�<	m�<G��<���<3��<���<���<���<n��<d��<���<��<T��<���<���<$��<2��<pg�<�C�<t�<���<��<؂�<-E�<	�<T��<�j�<��<ټ�<>]�<���<��<B�<���<3*�<
��<|"�<���<��<�o�<�Զ<Z5�<��<B�<;�<���<,Ԭ<��<|]�<���<�إ<
�<{F�<�x�<���<�՜<� �<)�<LO�<�s�<앓<���<�Տ<��< �<�)�<QC�<�[�<Ns�<��<Ꟁ<lj}<�y<��u<I�q<Ln<55j<_]f<��b<ʮ^<��Z<DW<	/S<0\O<܊K<;�G<\�C<�!@<1X<< �8<��4<�1<�M-<R�)<��%<�)"<�{<�<=-<Ǎ<��<w_<a�<�I<��<���;��;K��;��;c�;���;�)�;(��;d9�;/��;%��;�d�;<G�;�?�;&N�;�r�;W��;� �;oj�;�;��;�dv;W�k;F�a;��W;��M;��C;X:;��0;��';��;e�;�;w[;��:�*�:.��:G��:B�:-R�::��:�ۈ:��s:��V:�9:�:ä :�u�9�@�9`Z79�Ö8����6	��q��ܬ��C๠�	���"�q�;�N�T�.�m�i��KF��=h���x���{��n��U˺g.׺z�����u��������R|��B�� ��%���+��91���6��<��YB�eH���M�	lS�FY�(�^�Jxd��&j��o�9�u�<1{��o��G��u�������͋������~���W��2������  �  ��="(=W�=fp=E=�=d[=�� =�� =GD =���<�<�U�<K��<��<-�<�_�<c��<b��<��<�]�<]��<���<R�<�M�<���<��<���<|+�<�_�<���<���<���<"�<�N�<�y�<â�<���<	��<�<�2�<+Q�<�l�</��<���</��<���<��<���<}��<���<���<��<o��<���<���<?��<D��<�g�<D�<~�<���<��<��<ZE�<�<Q��<�j�<��<ü�<4]�<���<͌�<*�<ӥ�<+*�<騾<`"�<���<��<�o�<�Զ<J5�<��<-�<;�<���<,Ԭ<��<�]�<�<�إ<!�<�F�<y�<ʨ�<֜<� �<")�<_O�<�s�<��<���<�Տ<��<�<�)�<PC�<�[�<=s�<쉂<ӟ�<fj}<ٓy<μu<�q<n<5j<]f<��b<��^<N�Z<W<�.S<&\O<��K<�G<6�C<�!@<5X<<Q�8<<�4<�1<N-<k�)<��%<)*"<�{<B�<s-<��<��<�_<��<�I<��<ߜ�;���;{��;��;�b�;p��;�)�;��;G9�;���;斺;d�;G�;L?�;�M�;�r�;ѭ�;� �;j�;��;
��;�cv;��k;��a;��W;��M;@�C;�X:;|�0;��';W�;Q�;��;\;���:t,�:j��:���:�:�R�:��:�܈:e�s:N�V:��9:��:� :Vo�9�;�9rV79��8���@	��r�%ެ��K�š	�#�"���;���T�q�m�:��G��ni��Tz��|���m���T˺z+׺���ͼ�qt����������{��A� �w�%��+��81���6�?�<�:YB��
H���M�lS�rY���^�yd��'j�1�o��u��1{�0p���G�����s���΋�u���$��,X��i2������  �  ��=!(=`�=kp=C=�=[[=�� =�� =RD =���<�<	V�<\��<)��<=�<�_�<y��<z��<��<^�<i��<���<L�<�M�<��<��<���<u+�<�_�<u��<���<���<"�<�N�<~y�<���<���<���<��<�2�<Q�<�l�</��<���</��<���<���<���<���<���<���<#��<���<���<ϵ�<`��<[��<�g�<D�<��<���<#��<��<?E�<�<H��<�j�<��<¼�<]�<���<���<�<ϥ�<�)�<Ũ�<:"�<���<��<�o�<�Զ<+5�<���<-�<;�<���<Ԭ<��<�]�<ʜ�<�إ<(�<�F�<&y�<�<֜<� �<5)�<zO�<�s�<��<���<�Տ<�<	�<�)�<PC�<�[�<Qs�<쉂<ԟ�<6j}<��y<��u<��q<�n<�4j<�\f<N�b<r�^<,�Z<�W<�.S<�[O<��K<�G<Z�C<�!@<*X<<9�8<�4<�1<N-<��)<��%<a*"<|<e�<�-<�<0�<�_<��<�I<��<��;D��;i��;��;/c�;���;�)�;ۧ�;�8�;���;h��;d�;�F�;�>�;#M�;r�;ƭ�; �;�i�;y�;���;�cv;��k;��a;��W;��M;��C;�X:;�0;��';T�;}�;��;�\;���:�.�:���:;��:m�:�T�:B��:ވ:��s:�V:�9:�:'� :Hp�9�;�9tL79x��8"Z��-R	��	r��謹�S�A�	���"�Q�;��T���m����G��Gi���y��{���n���T˺-׺\��ֻ��s����)��Ͱ�{��@�w ���%��~+��81���6�-�<��XB�H��M�lS�/Y��^�yd��'j���o�~�u��2{��p���G��R�������΋�����e���X���2��S���  �  ��=(=T�=cp=F=�=a[=�� =�� =[D =���<�<
V�<T��<*��<2�<�_�<h��<���<��<^�<}��<���<k�<�M�<��<��<���<q+�<�_�<���<���<���<�!�<�N�<�y�<���<���<���<��<�2�<Q�<�l�<��<���<$��<���<���<
��<���<t��<���<��<���<���<ȵ�<Z��<X��<�g�<D�<��<���<*��<���<=E�<(�<B��<�j�<��<���<]�<���<Ì�<��<̥�<�)�<稾<P"�<i��<��<�o�<�Զ<*5�<<�<�:�<���<Ԭ<��<�]�<ߜ�<�إ<&�<�F�<y�<���<֜<� �<.)�<|O�<�s�<��<���<�Տ<!�<�<�)�<YC�<�[�<8s�<։�<ҟ�<j}<Гy<��u<��q<�n<�4j<+]f<G�b<Z�^<�Z<�W<�.S<�[O<��K<ݺG<*�C<�!@<7X<<b�8<-�4<1<�M-<��)<��%<L*"<|<U�<�-<
�<0�<�_<��<�I<��<f��;`��;���;��;�b�;F��;C)�;̧�;�8�;���;T��;�c�;\F�;�>�;�M�;�q�;���;���;�i�;��;���;�cv;�k;�a;A�W;P�M;��C;#Y:;o�0;F�';�;1�;��;�\;K��:;.�:���:s��:��:SV�:V��:�ވ:M�s:��V:m�9:O�:�� :'k�9':�9!H79���8�%���W	�5r�+bKไ�	���"�U�;���T��m���(H��Lj��C{��<|���n���R˺�,׺	��{��t��=�������[{��@�� ���%��~+��81�/�6�i�<�XB��
H���M��kS��Y���^��yd��'j�g�o�-�u��2{��p���G��q��F����΋�٦������X��e2������  �  ��=!(=`�=kp=C=�=[[=�� =�� =RD =���<�<	V�<\��<)��<=�<�_�<y��<z��<��<^�<i��<���<L�<�M�<��<��<���<u+�<�_�<u��<���<���<"�<�N�<~y�<���<���<���<��<�2�<Q�<�l�</��<���</��<���<���<���<���<���<���<#��<���<���<ϵ�<`��<[��<�g�<D�<��<���<#��<��<?E�<�<H��<�j�<��<¼�<]�<���<���<�<ϥ�<�)�<Ũ�<:"�<���<��<�o�<�Զ<+5�<���<.�<;�<���<Ԭ<��<�]�<ʜ�<�إ<(�<�F�<&y�<�<֜<� �<5)�<zO�<�s�<��<���<�Տ<�<	�<�)�<PC�<�[�<Qs�<쉂<ԟ�<6j}<��y<��u<��q<�n<�4j<�\f<N�b<r�^<,�Z<�W<�.S<�[O<��K<�G<Z�C<�!@<*X<<9�8<�4<�1<N-<��)<��%<a*"<|<e�<�-<�<0�<�_<��<�I<��<��;D��;i��;��;/c�;���;�)�;ۧ�;�8�;���;h��;d�;�F�;�>�;#M�;r�;ƭ�; �;�i�;y�;���;�cv;��k;��a;��W;��M;��C;�X:;�0;��';T�;}�;��;�\;���:�.�:���:;��:m�:�T�:B��:ވ:��s:�V:�9:�:'� :Hp�9�;�9tL79x��8"Z��-R	��	r��謹�S�A�	���"�Q�;��T���m����G��Gi���y��{���n���T˺-׺\��ֻ��s����)��Ͱ�{��@�w ���%��~+��81���6�-�<��XB�H��M�lS�/Y��^�yd��'j���o�~�u��2{��p���G��R�������΋�����e���X���2��S���  �  ��="(=W�=fp=E=�=d[=�� =�� =GD =���<�<�U�<K��<��<-�<�_�<c��<b��<��<�]�<]��<���<R�<�M�<���<��<���<|+�<�_�<���<���<���<"�<�N�<�y�<â�<���<	��<�<�2�<+Q�<�l�</��<���</��<���<��<���<}��<���<���<��<o��<���<���<?��<D��<�g�<D�<~�<���<��<��<ZE�<�<Q��<�j�<��<ü�<4]�<���<͌�<*�<ӥ�<+*�<騾<`"�<���<��<�o�<�Զ<J5�<��<-�<;�<���<,Ԭ<��<�]�<�<�إ<!�<�F�<y�<ʨ�<֜<� �<")�<_O�<�s�<��<���<�Տ<��<�<�)�<PC�<�[�<=s�<쉂<ӟ�<fj}<ٓy<μu<�q<n<5j<]f<��b<��^<N�Z<W<�.S<&\O<��K<�G<6�C<�!@<5X<<Q�8<<�4<�1<N-<k�)<��%<)*"<�{<B�<s-<��<��<�_<��<�I<��<ߜ�;���;{��;��;�b�;p��;�)�;��;G9�;���;斺;d�;G�;L?�;�M�;�r�;ѭ�;� �;j�;��;
��;�cv;��k;��a;��W;��M;@�C;�X:;|�0;��';W�;Q�;��;\;���:t,�:j��:���:�:�R�:��:�܈:e�s:N�V:��9:��:� :Vo�9�;�9rV79��8���@	��r�%ެ��K�š	�#�"���;���T�q�m�:��G��ni��Tz��|���m���T˺z+׺���ͼ�qt����������{��A� �w�%��+��81���6�?�<�:YB��
H���M�lS�rY���^�yd��'j�1�o��u��1{�0p���G�����s���΋�u���$��,X��i2������  �  ʃ=-(=`�=ip=D=�=U[=�� =�� =AD =}��<��<�U�<0��<���<�<|_�<G��<Q��<��<�]�<R��<���<H�<�M�<���<#��<���<�+�<�_�<���<��<���<+"�<�N�<�y�<ʢ�<���<��<�<�2�</Q�<	m�<G��<���<3��<���<���<���<n��<d��<���<��<T��<���<���<$��<2��<pg�<�C�<t�<���<��<؂�<-E�<	�<T��<�j�<��<ټ�<>]�<���<��<B�<���<3*�<
��<|"�<���<��<�o�<�Զ<Z5�<��<B�<;�<���<,Ԭ<��<|]�<���<�إ<
�<{F�<�x�<���<�՜<� �<)�<LO�<�s�<앓<���<�Տ<��<��<�)�<QC�<�[�<Ns�<��<Ꟁ<lj}<�y<��u<I�q<Ln<55j<_]f<��b<ʮ^<��Z<DW<	/S<0\O<܊K<;�G<\�C<�!@<1X<< �8<��4<�1<�M-<R�)<��%<�)"<�{<�<=-<Ǎ<��<w_<a�<�I<��<���;��;K��;��;c�;���;�)�;(��;d9�;/��;%��;�d�;<G�;�?�;&N�;�r�;W��;� �;oj�;�;��;�dv;W�k;F�a;��W;��M;��C;
X:;��0;��';��;e�;�;w[;��:�*�:.��:G��:B�:-R�::��:�ۈ:��s:��V:�9:�:ä :�u�9�@�9`Z79�Ö8����6	��q��ܬ��C๠�	���"�q�;�N�T�.�m�i��KF��=h���x���{��n��U˺g.׺z�����u��������R|��B�� ��%���+��91���6��<��YB�eH���M�	lS�FY�(�^�Jxd��&j��o�9�u�<1{��o��G��u�������͋������~���W��2������  �  ԃ=,(=g�=kp=B=�=N[=�� =u� =-D =P��<��<�U�<���<���<��<]_�<)��<&��<^�<�]�<K��<���<N�<�M�<��<)��<���<�+�<�_�<͒�<��<��<`"�<�N�<�y�<��<2��<4��<=�<�2�<EQ�<m�<D��<���<*��<���<���<���<[��<D��<x��<���<7��<o��<d��<���<���<Rg�<�C�<R�<���<��<̂�<+E�<�<J��<�j�<��<��<U]�<��<��<X�<:��<a*�<=��<�"�<喻<�<�o�<+ն<y5�<(��<M�<";�<���<"Ԭ<��<t]�<���<jإ<��<VF�<�x�<���<�՜<j �<�(�<O�<es�<���<`��<_Տ<��<��<�)�<OC�<�[�<]s�< ��<���<�j}<j�y</�u<��q<�n<�5j<�]f<�b<7�^<��Z<yW<l/S<c\O<�K<7�G<w�C<�!@<*X<<#�8<��4<�1<�M-<�)<I�%<�)"<Q{<��<�,<L�<`�<7_<�<EI<=�<���;���;S��;}�; c�;ƽ�;�)�;k��;�9�;���;q��;ge�;H�;:@�;�N�;Vs�;>��;4�;�j�;��;`��;�dv;0�k;��a;M�W;��M;��C;�W:;Z�0;��';Р;׶;�;�Y;���:�'�:���:H��:h�:�O�:(��:�ڈ:��s:��V:]�9:��:�� :�u�9�C�9ld79N�8x���,	���q�Ҭ�8��	���"��;���T�֐m����E���g���x���z���n���T˺/׺ �⺩��1x��8����ڳ�+~�	D�� ���%���+�7;1�.�6��<�ZB��H���M�lS�[Y���^�exd�5&j�d�o�ǁu�R0{�Ao��)F��������D͋�'���	~��}W��?1��s���  �  �=8(=k�=lp=;=޷=G[=q� =l� = D ='��<��<yU�<ј�<���<��<._�<���<���<N�<�]�<%��<���<=�<�M�<��<1��<��<�+�<`�<��<P��<5��<�"�<3O�<z�<*��<M��<g��<m�<3�<eQ�<7m�<X��<Ɯ�<+��<���<���<���<7��<8��<R��<���<
��<D��<=��<̟�<Ӆ�<'g�<�C�<)�<���<Ϻ�<���<.E�<�<M��<�j�<��<
��<y]�<+��<=��<��<Z��<�*�<p��<�"�<��<$�<+p�<Sն<�5�<N��<r�<-;�<���<!Ԭ<��<v]�<���<Sإ<��<(F�<�x�<i��<�՜<< �<�(�<�N�<5s�<���<B��<QՏ<��<��<�)�<>C�<�[�<is�<��<��<�j}<��y<��u<��q<�n<�5j<!^f<��b<v�^<0�Z<�W<�/S<�\O<B�K<h�G<��C<�!@<X<<�8<��4<]1<gM-<͒)<��%<K)"<�z<D�<�,<��<��<�^<��<I<�<ߛ�;���;��;P�;9c�;ܽ�;A*�;��;;:�;H��;0��;�e�;�H�;	A�;�O�;.t�;���;��;�k�;�;؃�;�ev;��k;6�a;C�W;�M;��C;�V:;+�0;8�';��;��;��;iX;:��: %�:��:r��:��:BM�:=��:f؈:�s:�V:ǅ9:��:�� :Cy�9�K�9�t79���8�g���	�,�q��Ĭ�?,๊�	�?�"���;�c�T�^�m�����B���e��0x��$z��)o���U˺/׺d��<��y����-��@��^��E�� ��%��+�o<1��6���<�4[B�~H�ȼM��lS�TY�Q�^��wd�I%j�N�o��u��.{��n���E�����b�]̋�����i}���V���0������  �  �=F(=n�=pp=>=׷=>[=d� =Z� =D =��<j�<HU�<���<N��<��<�^�<͟�<���<�<�]�<��<���<3�<�M�<��<?��<5��<�+�<)`�<��<���<g��<�"�<iO�<Bz�<g��<���<���<��<93�<�Q�<Gm�<n��<���<7��<���<���<���<��<��<&��<���<���<��<��<���<���<�f�<C�<�<��<���<���<E�< �<Z��<�j�<��< ��<�]�<X��<]��<��<���<�*�<���<#�<R��<X�<hp�<oն<�5�<c��<��<B;�<���<0Ԭ<��<c]�<|��<5إ<��<F�<�x�<4��<]՜<���<x(�<�N�<s�<t��<��<&Տ<��<��<�)�<BC�<�[�<is�<0��<(��<%k}<��y<�u<V�q<an<s6j<e^f<��b<�^<��Z<<W<�/S<�\O<b�K<��G<��C<�!@<X<<��8<��4<)1<M-<k�)<��%<�("<�z<��<�+<��<��<s^<\�<�H<��<m��;.��;���;f�;3c�;��;�*�;��;�:�;���;���;�f�;fI�;�A�; P�;u�;]��;��;	l�;��;D��;8fv;V�k;�a;��W;ۧM;��C;#V:;K�0;��';"�;l�;��;�V;���:;!�:��:��:F߶:�J�:��:�ֈ:��s:�V:�9:��:� :f~�9P�9h�79�&�8��������q������"�^�	���"���;�M�T�P�m�1���A��cd��w��,z��un��UV˺y0׺���?��m|����f����ƀ��G�p	 ���%���+��=1���6�ݨ<�\B��H�L�M�rlS��Y�J�^��vd��$j�7�o��u��-{��m���D�� ����lˋ�ѣ���|�� V��Y0��T���  �  ��=N(=u�=lp=;=ӷ=1[=\� =F� =�C =���<4�<U�<f��<-��<G�<�^�<���<���<��<j]�<���<���<5�<�M�<��<P��<D��<�+�<V`�<6��<���<���<�"�<�O�<�z�<���<���<���<��<n3�<�Q�<\m�<���<Ɯ�<,��<���<���<���<
��<���<��<O��<���<���<״�<i��<k��<�f�<IC�<��<W��<���<���<E�<
�<S��<k�<	�<6��<�]�<���<���<��<Ǧ�<+�<ݩ�<V#�<���<��<�p�<�ն<�5�<���<��<[;�<É�<&Ԭ<��<P]�<q��<إ<��<�E�<Mx�< ��<!՜<���<A(�<�N�<�r�<@��<���<�ԏ<��<��<�)�<?C�<�[�<ts�<D��<A��<gk}<D�y<%�u<��q<�n<�6j<�^f<\�b<H�^<��Z<�W<E0S<>]O<��K<ŻG<��C<�!@<X<<�8<m�4<1<�L-<)�)<K�%<~("<z<f�<�+<�<�<�]<�<`H<v�<+��;���;���;%�;c�;7��;�*�;e��;n;�;W��;r��;Cg�;J�;�B�;�P�;�u�;)��;W�;�l�;\�;���;�fv;��k;�a;-�W;�M;R�C;qU:;��0;O�';L�;��;X�;U;���:��:L��:��:�۶:�H�:m�:5Ո:p�s:cV:߅9:��:˨ :���9�T�9��79�Z�8Z��9��{�q������p�	���"� �;���T�h�m�"	��,@��yc���u��;z��Io���U˺�1׺� �3���~����*���������H�, �a�%�-�+�?1���6��<�y\B��H���M��lS�;Y���^�?vd�$j�2�o�d~u��,{�m��D��M���򈻰ʋ�����{��xU���/���
���  �  
�=T(={�=sp=9=η=$[=M� =5� =�C =���<�<�T�<-��<���<�<�^�<e��<���<��<G]�<��<|��<(�<�M�<!��<U��<[��<,�<d`�<U��<���<���<#�<�O�<�z�<���<���<���<��<~3�<�Q�<m�<���<ڜ�</��<���<���<}��<���<���<���<��<���<���<���<:��<9��<�f�<C�<��<=��<���<s��<�D�<��<V��<k�<�<Y��<�]�<���<���<&�<���<:+�<��<�#�<���<��<�p�<�ն<6�<���<��<b;�<ۉ�<(Ԭ<��<=]�<T��<�ץ<p�<�E�<x�<觞<�Ԝ<���<
(�<bN�<�r�<��<ٵ�<�ԏ<r�<��<�)�<6C�<�[�<�s�<J��<g��<�k}<l�y<�u<�q<+n<7j<P_f<��b<��^<^�Z<�W<v0S<f]O<�K<ݻG<��C<�!@<X<<Ґ8<9�4<�
1<�L-<��)<��%<2("<�y<��<P+<��<��<�]<��<.H<*�<���;U��;���;�;Qc�;=��;+�;��;�;�;���;���;�g�;�J�;C�;�Q�;Mv�;б�;�;Bm�;��;��;�gv;��k;��a;.�W;c�M;�C;^T:;��0;Q�';�;��;��;�S;k��:��:��:Z��:�ض:IF�:��:$ӈ:��s: ~V:��9:��:W� :ԃ�9�\�9%�79�i�8��������q����2๣�	�l�"�?�;�G�T��~m�U���=���a���u���x��To���V˺/3׺��?��4���G����i��{��J�� �v�%��+��@1�a�6�$�<�{]B��H��M��lS��Y�x�^�vd��"j�w�o��}u�+{�6l��NC������ʋ�K���{���T��9/��}
���  �  �=[(=z�=vp=6=ȷ=%[=C� =)� =�C =���<��<�T�<��<���<��<p^�<H��<c��<��<0]�<Ϛ�<��<�<�M�<!��<W��<i��<,�<�`�<z��<���<���<O#�<�O�<�z�<���<��<��<�<�3�<�Q�<�m�<���<Ҝ�<=��<{��<���<t��<���<���<���<��<P��<��<x��<��<��<mf�<C�<��< ��<o��<j��<�D�<��<e��<k�<�<j��<�]�<���<ߍ�<T�<��<v+�<>��<�#�<<��<�p�<�ն<16�<���<��<f;�<ډ�<4Ԭ<��<C]�<G��<�ץ<I�<�E�<x�<���<�Ԝ<��<�'�<-N�<�r�<���<���<�ԏ<^�<��<~)�<,C�<�[�<~s�<W��<n��<�k}<��y<׾u<K�q<mn<�7j<�_f<�b<��^<��Z<2W<�0S<�]O<�K<��G<��C<�!@<�W<<��8<<�4<�
1<UL-<��)<��%<�'"<fy<��<�*<U�<m�<Z]<a�<�G<��<Q��;V��;5��;�;Ac�;8��;1+�;��;<�;O��;���;Yh�;�K�;�C�;@R�;/w�;C��;��;�m�;�;{��;"hv;�k;P�a;��W;�M;��C;
T:;��0;^�';Ś;Y�;��;R;���:��:7��:^��:L׶:D�:��:�ш:�s:�}V:��9:3�:�� :f��9&`�9��795��8C�����qq�������߹�y	���"���;��T�]zm�c���<���`���u��1y���n���W˺�2׺�㺞��Ă��L�t��F������K�4 ��%���+�hA1���6���<�^B��H�*�M�mS��Y���^��ud��"j�w�o��|u��){��k���B�����g�2ɋ������z��T���.���	���  �  �=l(=��=wp=3=��=[=9� =&� =�C =y��<��<�T�<���<���<��<O^�<.��<O��<��<.]�<���<h��<�<�M�< ��<w��<��<,,�<�`�<���<��<��<b#�<P�<�z�<��<��<8��<�<�3�<�Q�<�m�<���<ל�<?��<u��<���<a��<���<���<���<���<.��<w��<^��<��<��<Kf�<�B�<��<��<g��<V��<�D�<��<g��<k�<F�<x��<^�<���<��<r�<7��<�+�<\��<�#�<��<�<q�< ֶ<Q6�<ё�<��<�;�<܉�<2Ԭ<��<-]�<3��<�ץ<2�<�E�<�w�<���<�Ԝ<^��<�'�<N�<_r�<攓<���<�ԏ<M�<�<j)�<'C�<�[�<�s�<~��<y��<l}<ٕy<��u<��q<�n<�7j<�_f<T�b<,�^<��Z<\W<�0S<�]O<�K<?�G<��C<�!@<�W<<��8<�4<z
1<IL-<]�)<��%<�'"<,y<}�<�*<:�<'�<"]<6�<�G<��<��;��;���; �;6c�;���;+�;L��;o<�;t��;��;�h�;�K�;YD�;�R�;�w�;���;�;�m�;q�;���;ehv;��k;r�a;��W;��M;�C;hS:;y�0;ޭ';��;��;}�;�Q;Ϸ�:��:ӽ�:3��:�ն:rB�:j�:9ш:��s:�zV:�9:0�:�� :&��9c�9I�79Ѧ�85���u���dq�������߹]v	���"�1�;�t�T� ym�����;���_��&s��4y��o���X˺q4׺�����Q�����-��\�����L�� ���%���+��A1���6�3�<��^B�UH�˾M�HmS��Y�/�^�ntd�V"j���o�|u�,){�Sk��fB��c����ȋ�P���0z���S��h.���	���  �  �=b(=�=tp=9=Ƿ=[=8� =� =�C =[��<��<�T�<Η�<���<��<F^�<��<6��<��<]�<���<g��<�<�M�<!��<g��<r��<?,�<�`�<���<#��<#��<|#�<*P�<{�< ��<D��<F��<.�<�3�<�Q�<�m�<���<֜�<3��<���<���<d��<���<x��<���<���<+��<V��<<��<͞�<���<Jf�<�B�<q�<���<V��<Y��<�D�<��<^��<k�<,�<}��<^�<���<��<|�<^��<�+�<���<�#�<��<'�<q�< ֶ<T6�<味<��<};�<���<6Ԭ<��</]�<3��<�ץ< �<qE�<�w�<���<�Ԝ<<��<�'�<N�<Vr�<Ɣ�<���<�ԏ<G�<~�<v)�<2C�<�[�<�s�<h��<���<l}<��y<'�u<��q<�n<�7j<!`f<t�b<q�^<�Z<�W<1S<�]O</�K<�G<��C<�!@<X<<��8<�4<v
1<L-<E�)<Q�%<{'"<y<)�<e*<�<�<�\<�<tG<��<��;��;7��;�;3c�;j��;D+�;���;n<�;���;4��;?i�;)L�;�D�;.S�;�w�;=��;5�;ln�;��;���;�hv;��k;\�a;.�W;)�M;_�C;yS:;
�0;�';]�;��;[�;�P;���:��:F��:��:�Ӷ:A�:��:Ј:��s:?{V:#�9:��:ު :r��9d�9��79۪�8n��Y���Qq�}���,�߹s	�V�"��;���T�Cum�y���:��&`��Pt��y���n��yW˺r4׺�I��w�����#�����T���M� �]�%��+��B1�!�6��<��^B�[H�e�M��lS��Y�n�^�ud��!j�m�o��{u�~({��j���A��%��q����ȋ�Ǡ���y���S��.��{	���  �  K�=�*=��=�s= =��=�_=M=�� =�I =��<Y�<2c�<v��<T��<�.�<Dq�<C��<���<N5�<#u�<;��<B��<\/�<bk�<i��<=��<��<*P�<$��<ں�<���<��<�O�<c~�<B��<#��<D��<D&�<FK�<�m�<E��<��<@��<���<��<��<��<�"�<;+�<0�<E1�<�.�<�'�<�<��<_��<8��<c��<���<�|�<�P�<c�<���<��<�i�<�!�<=��<���<�&�<L��<�a�<d��<��<�<4��<��<ㆽ<z��<�f�<�θ<2�< ��<~�<2>�<j��<Kڮ<�!�<�e�<���<��<��<P�<���<��<�ޞ<	�<�0�<pV�<�y�<y��<-��<8ّ<���<��<*�<YB�<dY�<no�<���<���<!��<�}}<�y<=�u<]�q<Sn<�.j<Rf<�tb<��^<�Z<0�V<�S<0O<YK<��G<�C<p�?<<<8B8<x4<�0<��,<U,)<�o%<
�!<�<vS<3�<�<�d<�<�7<�<�$<$L�;�\�;�|�;ͬ�;���;�?�;���;�;���;cA�;�;e��;��;���;͓�;۳�;��;�:�;B��;$!�;�o};	�r;�Yh;^;� T;�J;Sa@;��6;w-;�C$;�;;U];ʨ	;�;�k�:���:���:l��:��:]��:�w�:���:��i:x|L:��/:2�:�)�9M�9�_�9[�9J$08߇v�K&���O��;.�����(���A��cZ�1�r�����7���Lĝ���������g����[ͺ�!ٺ����4��{����	��w�i9���կ ��e&��,���1��u7��!=���B�XsH��N���S��gY�}_���d��Yj���o��u��L{�0z���M���!�������ʋ������u��#L��-#�������  �  H�=�*=��=�s==��=�_=C=�� =�I =��<d�<;c�<���<Q��<�.�<Iq�<M��<���<U5�<-u�<&��<D��<d/�<qk�<k��<6��<��<)P�<*��<ɺ�<���<��<�O�<U~�<��<"��<A��<K&�<<K�<�m�<C��<��<A��<���<'��<��<��<�"�<3+�<0�<A1�<�.�<�'�<�<��<c��<H��<h��<���<�|�<�P�<^�<���<��<�i�<	"�<5��<���<�&�<L��<�a�<Y��<��<�<5��<��<φ�<y��<�f�<�θ<�1�<#��<{�<->�<e��<Jڮ<�!�<�e�<���<��<��<$P�<���<��<�ޞ<	�<�0�<zV�< z�<���<8��<8ّ<���<��<*�<\B�<kY�<uo�<v��<���<��<�}}<d�y</�u<f�q<Wn<�.j<�Qf<�tb<��^<��Z<(�V<qS<
0O<YK<��G<��C<y�?<<<AB8<�w4<İ0<��,<Y,)<�o%<!�!<<�S<.�<"<�d< �<�7< �<�$<�K�;�\�;�|�;��;���;�?�;���;�;���;"A�;�;Q��;��;Ɖ�;A��;ٳ�;��;
;�;��;!�;�o};��r;�Yh;�^;T;J;na@;��6;�v-;�C$;�;;�];�	;7;$l�:���:���:���:m�:��:�x�:Y��:��i:}L:t�/:D�:�'�9V�9�^�9��9V 08˜v��G&�􆹁N���5�U��(�(�R�A��cZ��r�]���R����ĝ������J���<[ͺ�!ٺQ��}���3��~��f�	�w��8����� �7e&�.,�6�1��u7�!=��B��sH��N�~�S��gY��_���d��Yj���o�|�u�-M{�z���M���!��^���ˋ�ퟎ��u��3L��l#��v����  �  =�=�*={�=�s== �=�_=F=�� =�I =?��<z�<Jc�<���<n��<�.�<Tq�<h��<���<i5�<Gu�<0��<V��<b/�<ok�<c��</��<��<P�<��<���<���<��<�O�<C~�<��<��<��<6&�<%K�<�m�<.��<���<>��<���<)��<��<��<�"�<B+�<90�<W1�<�.�<�'�<(�<�<���<`��<s��<���<�|�<�P�<q�<���<(��<�i�<	"�<)��<��<�&�<4��<�a�<>��<���<��<��<��<���<]��<�f�<�θ<�1�<��<`�< >�<]��<>ڮ<�!�<�e�<���<��<��<:P�<���<,��<�ޞ<7	�<1�<�V�<z�<���<Z��<Lّ<���<��<!*�<cB�<kY�<vo�<l��<���<��<�}}<6�y<
�u</�q<n<�.j<�Qf<�tb<[�^<��Z<�V<>S<�/O<�XK<��G<�C<r�?<<<GB8< x4<Ӱ0<�,<~,)<�o%<N�!<-<�S<i�<l<�d<Y�<8<*�<'%<L�;]�;�|�;��;���;�?�;{��;��;���;�@�;��;ƹ�;���;���;֒�;���;&�;�:�;ɡ�;� �;'o};r�r;�Yh;j^;"T;�J;�a@;0�6;Vw-;�D$;\<;�^;n�	;�;In�:���:���:���:��:���:nz�:���:�i:L:��/:z�:0%�9i�97Z�9^�9��/8��v�'R&������S��<�}��R�(��A��eZ�m�r�w���޻��Gŝ�L���O���c���{[ͺz ٺ�����2�����w�	� w��7�%��^� ��d&��,�!�1�u7�2 =���B� sH�eN���S��gY�6_���d�gZj�P p�6�u��M{��z��bN��G"������Lˋ�����=v��vL���#�������  �  6�=�*=x�=�s=	=�=�_=Z=�� =�I =[��<��<|c�<˧�<���<�.�<�q�<���<���<}5�<Xu�<U��<Z��<i/�<tk�<d��<��<��<�O�<���<���<���<t�<�O�<~�<��<���<���<&�<K�<�m�<!��<��<#��<���< ��<��<��<�"�<^+�<?0�<v1�<�.�<%(�<U�<:�<���<���<���<֣�<�|�<�P�<��<���<(��<�i�<"�<)��<e��<�&�<&��<�a�<��<τ�<��<��<��<���<)��<�f�<�θ<�1�<돵<P�<>�<G��<=ڮ<�!�<�e�<���<��<��<KP�<ǂ�<M��<ߞ<U	�<(1�<�V�<Bz�<ě�<w��<hّ<���<��<1*�<hB�<rY�<po�<j��<���<���<�}}<��y<��u<��q<�n<m.j<QQf<atb<�^<r�Z<��V<S<�/O<�XK<e�G<ٯC<m�?<%<<QB8<9x4<"�0<)�,<�,)<.p%<��!<�<&T<��<�<?e<��<Q8<Y�<N%<�L�;/]�;&}�;,��;���;i?�;<��;|�;
��;f@�;Q�;U��;畬;ڈ�;p��;ز�;��;$:�;M��;K �;�n};�r;Yh;�^;� T;NJ;b@;��6;Ex-;E$;b=;�_;�	;R;q�:���:���:���:c�:���:{�:��:ʐi:gL:��/:��:�%�9��9/W�9��9��/8@w��g&�o�� `��/D���c�(���A�]kZ���r���������0Ɲ�����@�������ZͺF ٺ���	��\1�����c�	�yu��6����:� �"c&�,,�9�1�?t7��=���B�{rH�AN�M�S��gY�C_���d��Zj�p��u��N{�{���N��#��8���̋�2����v��M��9$������  �  ,�=�*=w�=�s=
=�=�_=i=�� =�I =���<��<�c�<���<���</�<�q�<���<��<�5�<yu�<q��<g��<~/�<rk�<a��<��<��<�O�<΅�<m��<���<F�<]O�<�}�<���<���<���<�%�<�J�<�m�<���<ث�<��<���<��<��<��<�"�<�+�<i0�<�1�<�.�<](�<��<p�<���<���<���<���<2}�<Q�<��<���<4��<j�<�!�<#��<R��<�&�<���<Ya�<���<���<��<���<F�<M��<���<Sf�<oθ<�1�<���<2�<�=�<8��<4ڮ<�!�<�e�<���<�<��<{P�<���<x��<^ߞ<�	�<k1�<�V�<wz�<���<���<�ّ<���<��<D*�<zB�<|Y�<jo�<j��<���<嫀<8}}<��y<Z�u<}�q<Xn<�-j<�Pf<�sb<��^<�Z<N�V<�S<Y/O<�XK<:�G<ԯC<`�?<)<<uB8<Zx4<^�0<h�,<,-)<�p%<
�!<<�T<K�<<�e<�<�8<ͫ<�%<"M�;t]�;�}�;4��;���;Z?�;���;7�;c��;�?�;��;���;0��;�;���;ޱ�;
�;Z9�;���;��;�m};d�r;�Xh;�^;� T;�J;�b@;��6;ky-;rF$;H?;�`;Ϭ	;�;~t�:Z��:J��:r��:��:1��:�}�:[��:�i:C�L:��/:�:e%�9��9EQ�9_�9�V/8�aw�+�&�L���o��mR�4���(�p�A��qZ���r�u���X����ǝ�:�������^����Yͺ�ٺ��亶��:.������	�zs�5������ �va&��,���1�pr7��=���B��qH��N��S��gY�E_��d�r[j�fp�c�u�zP{��{���O��$��(���͋�㡎��w���M���$�������  �  �=�*=o�=�s=	=�=�_=v=Ӧ =�I =���<�<�c�<G��<��<S/�<�q�<���<L��<�5�<�u�<���<���<�/�<rk�<V��<��<��<�O�<���<:��<a��<��<O�<�}�<j��<k��<{��<�%�<�J�<km�<э�<���<	��<���<��<��<�<#�<�+�<�0�<�1�<:/�<�(�<��<��<(��<���<��<B��<[}�<:Q�<��<���<G��<�i�<�!�<��<H��<|&�<���<7a�<���<_��<4�<m��< �<��<���<�e�<=θ<\1�<���<�<�=�<-��<$ڮ<�!�<�e�<ѥ�<)�<�<�P�<#��<���<�ߞ<�	�<�1�<=W�<�z�<1��<໓<�ّ<��<��<j*�<�B�<wY�<io�<U��<m��<���<�|}<^�y<�u<��q<�
n<�-j<JPf<{sb<�^<z�Z<��V<`S</O<5XK<�G<��C<X�?<#<<�B8<�x4<��0<��,<x-)<q%<��!<x<(U<Ѫ<�<&f<��<"9<�<�%<�M�;^�;�}�;G��;���;D?�;���;��;���;?�;��;���;B��; ��;���;+��;��;�8�;���;'�;�l};`�r;jXh;^;� T;�J;5c@;��6;Qz-;�G$;�@;+c;y�	;�!;�x�:���:U��:���:b �:�:���:[��:�i:�L:��/:d�:� �9�9;I�9B�9>/8��w���&�9%���|���b����(�p�A�KwZ��r�H�������qɝ�����M���Z����Yͺvٺ �����+������	�$r��2����\� ��_&��,���1�4q7�E=���B��pH�<N�+�S��gY��_���d��\j�}p���u��Q{��|���P���$��>����͋�����x���N��%��O����  �  �=�*=a�=�s==�=�_=�=� =
J =���<W�<3d�<���<L��<�/�<9r�<C��<���<6�<�u�<���<���<�/�<�k�<I��<���<h�<�O�<���<��<,��<��<�N�<T}�<��<+��<:��<p%�<fJ�<2m�<���<���<���<i��<,��<��<�<##�<�+�<�0�<�1�<�/�<�(�<�<��<`��<G��<K��<���<�}�<lQ�<��<���<W��<�i�<	"�<���<%��<V&�<���< a�<m��<'��<��<)��<��<���<l��<�e�<θ<1�<e��<��<�=�<	��<ڮ<"�<�e�<ᥩ<<�<8�<�P�<W��<���<�ߞ<
�<�1�<�W�<�z�<s��<!��<�ّ<S��<�<~*�<�B�<�Y�<qo�<=��<S��<���<�|}<ؠy<��u<��q<A
n<-j<�Of<�rb<��^<�Z<x�V<�S<�.O<�WK<ւG<y�C<Y�?<L<<�B8<�x4<̱0<5�,<�-)<q%<�!<<�U<9�<W<�f<*�<�9<��<e&<N�;r^�;�}�;���;���;�>�;@��;	�;g��;>�;$�;���;[��;��;P��;<��;��;�7�;���;Q�;�k};d�r;�Wh;`^;�T;4J;�c@;c�6;�{-;�I$;�A;ee;��	;|$;�|�:?��:x��:���:�$�:|��:���:팃:��i:l�L:��/:�:v�9�޷9�@�9҅9+�.8�Lx���&�
5��D����w�x���(���A��}Z�< s������Ñ�[˝��é�F���ȇ��LYͺ0ٺ���6���(�������	�p�d0�4��=� �R]&��,���1�p7��=���B�&pH��N���S��gY��_�{�d��]j��p���u��S{��}���Q���%�������΋� ���oy��O���&�������  �  ��=�*=_�=�s=="�=�_=�=� =-J =8��<��<rd�<֨�<���<�/�<yr�<s��<���<G6�<�u�<ɴ�<���<�/�<�k�<;��<���<U�<sO�<Q��<ι�<���<~�<�N�<}�<ߩ�<���<���<(%�<2J�< m�<���<|��<���<c��<��<��<1�<C#�<�+�<�0�<E2�<�/�<	)�<O�<=�<���<���<���<���<�}�<�Q�< �<��<r��<j�<�!�<���<��<<&�<w��<�`�<=��<ۃ�<��<ҏ�<i�<r��<��<xe�<�͸<�0�<*��<��<�=�<���< ڮ<�!�<�e�<���<[�<W�<Q�<���<-��<��<[
�<32�<�W�<9{�<���<X��<6ڑ<|��<:�<�*�<�B�<�Y�<Yo�<;��<B��<~��<F|}<��y<�u<�q<�	n<c,j<8Of<Xrb<�^<��Z<��V<}S<X.O<�WK<��G<m�C<+�?<O<<�B8<�x4<�0<��,<Z.)<�q%<~�!<�<QV<�<�<>g<��<(:<�<�&<�N�;�^�;H~�;���;o��;�>�;��;��;���;�=�;)�;µ�;7��;��;���;��;��;�6�;>��;��;:j};��r;Wh;J^;� T;�J;�d@;q�6;�|-;)K$;D;g;i�	;h&;���:}�:`��:y��:$(�:��:��:k��:Ӟi:A�L:L�/:<�:��9�ٷ9S;�9�p9�M.8��x���&�5E������k��y��)���A���Z��s�H����ő��̝�qĩ����������Wͺvٺ�����%�����&�	�n�h.�u��� �Y[&��,�3�1��m7�Z=���B�RoH�N�Y�S�zhY��_��d��^j�2p��u��U{��~���R��'��Z���Ћ�#����z��mP��:'�������  �  �=�*=Y�=�s==+�=`=�=� =CJ =g��<��<�d�<��<���<0�<�r�<���<���<k6�<v�<��<���<�/�<�k�<@��<���<0�<ZO�<��<���<���<F�<WN�<�|�<���<���<���<�$�<J�<�l�<Z��<a��<���<d��<��<��<5�<a#�<,�<1�<w2�<�/�<Y)�<��<y�<���<���<���<��<�}�<�Q�<7 �<$��<u��<j�<�!�<���<��<&�<P��<�`�<��<���<v�<���< �<)��<���<>e�<o͸<�0�<���<��<o=�<���<ڮ<�!�<�e�<��<}�<{�<$Q�<���<e��<R��<�
�<u2�<�W�<{{�<���<���<fڑ<���<e�<�*�<�B�<�Y�<Yo�<3��<��<c��<�{}<8�y<��u<��q<V	n<�+j<�Nf<�qb<��^<	�Z<��V<2S<�-O<tWK<a�G<S�C<-�?<Y<<�B8<2y4<v�0<��,<�.)<Tr%<�!<$<�V<|�<E<�g<�<�:<^�<'<eO�;G_�;�~�;���;���;�>�;���;F�;��;=�;5�;���;]��;��;���;��;\�;�5�;���;�;i};�r;1Vh;k^;� T;LJ;e@;u�6;A~-;L$;�E;�h;��	;?(;���:��:���:���:E+�:��:爒:���:Ţi:�L:��/:$�:�9yӷ9)4�9&_9]�-8��x���&��P��ΰ��L��	��)�j�A��Z��	s�V���pǑ��Ν��ũ�����܈��RVͺ�ٺ;�亯~��"�����X�	��k��,�`��8� �JY&��,�ɽ1�Sl7�^=�7�B�ynH��N��S�zhY�_�8�d��_j��p�&�u�6W{�����S��,(��X���2ы�쥎�z{��MQ���'��w����  �  م=�*=O�=�s==,�=`=�=(� =WJ =���< �<�d�<H��<#��<W0�<�r�<��<$��<�6�<Hv�<��<���<�/�<�k�<4��<���<�<:O�<���<l��<��<�<#N�<�|�<Z��<`��<���<�$�<�I�<�l�<4��<D��<���<Q��<��<��<B�<w#�<.,�<C1�<�2�<0�<�)�<��<��<(��<���<���<��<~�<�Q�<V �<:��<���<j�<�!�<���<��<�%�<(��<f`�<���<b��<7�<R��<��<���<���<e�<C͸<w0�<Ȏ�<e�<S=�<̍�<�ٮ<�!�<�e�<��<��<��<PQ�<<���<}��<�
�<�2�<<X�<�{�<$��<���<�ڑ<���<z�<�*�<�B�<�Y�<[o�<��<��<G��<�{}<ȟy<J�u<,�q<�n<j+j</Nf<[qb<&�^<��Z<.�V<�S<�-O<7WK<@�G<*�C<*�?<b<<�B8<Zy4<��0<"�,</)<�r%<z�!<�<=W<��<�<;h<��<�:<��<a'<�O�;�_�;�~�;��;t��;i>�;H��;��;n��;*<�;��;/��;���;A��;���;;��;l�;5�;ќ�;T�;�g};?�r;�Uh;�^;&T;�J;�e@;;�6;2-;�M$;G;'j;Q�	;*;z��:0	�:���:9��:c.�:���:勒:%��:եi:��L:��/:�:'�9з9]-�9.M9J�-8?my� '�m_��I�������+)�V�A��Z�s�ز���ɑ�!Н��Ʃ�����q���bVͺ�ٺ���|� �������	�Bj��*����J� ��W&�",��1�k7��=���B��mH�}N���S�nhY��_���d�h`j��p��u��X{������T���(��e���ҋ�٦��;|��R���(�������  �  ƅ=�*=M�=�s==0�=`=�=7� =dJ =���<$ �<e�<x��<=��<�0�<s�<��<F��<�6�<\v�<��<���<�/�<�k�<-��<���<�<O�<��<O��<b��<��<�M�<p|�<4��<A��<Z��<�$�<�I�<�l�<"��<&��<���<F��<��<��<V�<�#�<:,�<c1�<�2�<>0�<�)�<��<��<J��<$��<��<D��<9~�< R�<` �<E��<���<j�<�!�<���<��<�%�<��<W`�<���<A��<��<+��<��<�<i��<�d�<"͸<T0�<���<B�<>=�<ō�<�ٮ<�!�<�e�<'��<��<��<jQ�<��<���<���<�
�<�2�<jX�<�{�<C��<㼓<�ڑ<���<��<�*�<�B�<�Y�<Vo�<��<	��<"��<�{}<��y<�u<��q<on<*+j<�Mf<qb<��^<Q�Z<��V<�S<�-O<�VK<*�G<�C<�?<d<<C8<�y4<��0<^�,<:/)<s%<��!<�<�W<0�<0<�h<��<;;<��<�'<
P�;`�;�~�;��;e��;e>�;��;K�;X��;�;�;:�;��;㏬;���;��;Ȭ�;��;�4�;V��;�;|g};]�r;�Uh;�^;T;�J;2f@;��6;�-;�N$;�G;�k;_�	;�+;��:g�:���:M��:?1�:���:֍�:ؔ�:a�i:ďL:��/:)�:s�9gϷ9l'�9�B9��-8��y�i'��l��Ǻ������)�c�A���Z��s�J����ˑ�>ѝ��Ʃ�+���Ї���Vͺٺ���2{�X�����t�	�:i�\)����ӟ �aV&�#
,�غ1�?j7��=��B�0mH�N���S��hY��_�ոd��aj�	p���u��Y{� ���tU��u)������ҋ������|��vR��)��* ���  �  =�*=L�=�s==6�=`=�=>� =qJ =���<F �<6e�<���<Y��<�0�<As�<%��<Y��<�6�<mv�<'��<���<�/�<�k�</��<���<��<O�<ׄ�<;��<?��<��<�M�<K|�<��< ��<N��<x$�<�I�<�l�<��<��<���<J��<��<��<[�<�#�<S,�<w1�<�2�<Q0�<�)�<�<��<a��<8��<F��<W��<Q~�<R�<w �<T��<���<$j�<�!�<���<��<�%�<���<:`�<���<��<��<��<��<���<S��<�d�<�̸<=0�<���<3�<*=�<���<�ٮ<�!�<�e�<)��<��<��<Q�<"��<Գ�<���<�<�2�<|X�<�{�<h��<�<�ڑ<���<��<�*�<�B�<�Y�<Yo�<��<���<��<U{}<t�y<��u<��q<Wn<�*j<�Mf<�pb<��^<#�Z<��V<`S<c-O<�VK<�G<�C<�?<l<<C8<�y4<�0<y�,<n/)<0s%<�!<'<�W<k�<X<�h<�<d;<'�<�'<dP�;+`�;�~�;��;u��;G>�;Ҡ�;3�;��;y;�;��;B��;���;$��;���;L��;x�;/4�;���;��;�f};�r;VUh;�^;&T;�J;`f@;!�6;l�-;PO$;�H;3l;��	;R,;$��:��:��:���:}2�:¡:G��:[��:��i:K�L: �/:�:��9#˷9�#�9�79�O-8M�y�7/'��o���ͺ����O��)��A��Z��s����`̑�[ҝ��ǩ����������Uͺ�ٺ����y����I����	��g��(����E� �\U&�	,�b�1�ki7��=�?�B�mH��N�ÿS��hY��_�c�d��aj��	p�4�u��Z{������U��*�����Ӌ�ڧ��<}���R��f)��� ���  �  ̅=�*=I�=�s==;�=`=�=<� =yJ =���<E �<5e�<���<���<�0�<As�<��<b��<�6�<mv�<,��<���<�/�<�k�<)��<���< �<O�<Ą�<<��<4��<��<�M�<D|�<��<��<J��<m$�<�I�<vl�<��<,��<���<C��<��<��<^�<�#�<T,�<s1�<�2�<M0�<�)�<�<�<{��<6��<K��<P��<\~�<R�<v �<X��<���<)j�<�!�<���<��<�%�<���<0`�<���<��<��<���<��<���<G��<�d�<�̸<?0�<���<<�<1=�<���<�ٮ<�!�<�e�<&��<��<��<�Q�<,��<γ�<���<�<
3�<�X�<�{�<l��<�<�ڑ<���<��<�*�<�B�<�Y�<Jo�<��<���<-��<>{}<h�y<��u<��q<Kn<�*j<�Mf<�pb<��^<�Z<��V<ZS<G-O<WK<�G<�C<�?<f<<3C8<�y4<��0<r�,<�/)<6s%<�!<%<�W<��<a<�h<�<v;<A�<�'<wP�;'`�;2�;��;^��;?>�;��;i�;���;~;�;��;��;{��;
��;���;��;j�;4�;���;��;�f};��r;KUh;�^;� T;�J;�f@;N�6;s�-;7O$;+I;l;ɸ	;S,;���:��:���:-��:2�:�¡:I��:Q��:�i:h�L:��/:̓:a�9Lʷ9�'�9�89s=-8B�y��4'��p��`Һ������)�?�A�X�Z�]s������ˑ��ѝ��ǩ�7���Ĉ��Uͺ�ٺ����y�j������	��g��(����� �dU&��,�[�1��h7��=�/�B�mH��N�ܿS��hY�_�d�d�8aj�P
p�c�u��Z{������U��Q*��s���VӋ�����h}��S��s)��� ���  �  =�*=L�=�s==6�=`=�=>� =qJ =���<F �<6e�<���<Y��<�0�<As�<%��<Y��<�6�<mv�<'��<���<�/�<�k�</��<���<��<O�<ׄ�<;��<?��<��<�M�<K|�<��< ��<N��<x$�<�I�<�l�<��<��<���<J��<��<��<[�<�#�<S,�<w1�<�2�<Q0�<�)�<�<��<a��<8��<F��<W��<Q~�<R�<w �<T��<���<$j�<�!�<���<��<�%�<���<:`�<���<��<��<��<��<���<S��<�d�<�̸<=0�<���<3�<*=�<���<�ٮ<�!�<�e�<)��<��<��<Q�<"��<Գ�<���<�<�2�<|X�<�{�<h��<�<�ڑ<���<��<�*�<�B�<�Y�<Yo�<��<���<��<U{}<t�y<��u<��q<Wn<�*j<�Mf<�pb<��^<#�Z<��V<`S<c-O<�VK<�G<�C<�?<l<<C8<�y4<�0<y�,<n/)<0s%<�!<'<�W<k�<X<�h<�<d;<'�<�'<dP�;+`�;�~�;��;t��;G>�;Ҡ�;3�;��;y;�;��;B��;���;$��;���;L��;x�;/4�;���;��;�f};�r;VUh;�^;&T;�J;`f@;!�6;l�-;PO$;�H;3l;��	;R,;$��:��:��:���:}2�:¡:G��:[��:��i:K�L: �/:�:��9#˷9�#�9�79�O-8M�y�7/'��o���ͺ����O��)��A��Z��s����`̑�[ҝ��ǩ����������Uͺ�ٺ����y����I����	��g��(����E� �\U&�	,�b�1�ki7��=�?�B�mH��N�ÿS��hY��_�c�d��aj��	p�4�u��Z{������U��*�����Ӌ�ڧ��<}���R��f)��� ���  �  ƅ=�*=M�=�s==0�=`=�=7� =dJ =���<$ �<e�<x��<=��<�0�<s�<��<F��<�6�<\v�<��<���<�/�<�k�<-��<���<�<O�<��<O��<b��<��<�M�<p|�<4��<A��<Z��<�$�<�I�<�l�<"��<&��<���<F��<��<��<V�<�#�<:,�<c1�<�2�<>0�<�)�<��<��<J��<$��<��<D��<9~�< R�<` �<E��<���<j�<�!�<���<��<�%�<��<W`�<���<A��<��<+��<��<�<i��<�d�<"͸<T0�<���<B�<>=�<ō�<�ٮ<�!�<�e�<'��<��<��<jQ�<��<���<���<�
�<�2�<jX�<�{�<C��<㼓<�ڑ<���<��<�*�<�B�<�Y�<Vo�<��<	��<"��<�{}<��y<�u<��q<on<*+j<�Mf<qb<��^<R�Z<��V<�S<�-O<�VK<*�G<�C<�?<d<<C8<�y4<��0<^�,<:/)<s%<��!<�<�W</�<0<�h<��<;;<��<�'<
P�;`�;�~�;��;e��;e>�;��;K�;X��;�;�;:�;��;⏬;���;��;Ȭ�;��;�4�;V��;�;|g};]�r;�Uh;�^;T;�J;2f@;��6;�-;�N$;�G;�k;_�	;�+;��:g�:���:M��:?1�:���:֍�:ؔ�:a�i:ďL:��/:)�:s�9gϷ9l'�9�B9��-8��y�i'��l��Ǻ������)�c�A���Z��s�J����ˑ�>ѝ��Ʃ�+���Ї���Vͺٺ���2{�X�����t�	�:i�\)����ӟ �aV&�#
,�غ1�?j7��=��B�0mH�N���S��hY��_�ոd��aj�	p���u��Y{� ���tU��u)������ҋ������|��vR��)��* ���  �  م=�*=O�=�s==,�=`=�=(� =WJ =���< �<�d�<H��<#��<W0�<�r�<��<$��<�6�<Hv�<��<���<�/�<�k�<4��<���<�<:O�<���<l��<��<�<#N�<�|�<Z��<`��<���<�$�<�I�<�l�<4��<D��<���<Q��<��<��<B�<w#�<.,�<C1�<�2�<0�<�)�<��<��<(��<���<���<��<~�<�Q�<V �<:��<���<j�<�!�<���<��<�%�<(��<f`�<���<b��<7�<R��<��<���<���<e�<C͸<w0�<Ȏ�<e�<S=�<̍�<�ٮ<�!�<�e�<��<��<��<PQ�<<���<}��<�
�<�2�<<X�<�{�<$��<���<�ڑ<���<z�<�*�<�B�<�Y�<[o�<��<��<G��<�{}<ȟy<J�u<,�q<�n<j+j</Nf<[qb<&�^<��Z<.�V<�S<�-O<7WK<@�G<*�C<*�?<b<<�B8<Zy4<��0<"�,</)<�r%<z�!<�<=W<��<�<;h<��<�:<��<a'<�O�;�_�;�~�;��;t��;i>�;H��;��;m��;*<�;��;/��;���;A��;���;;��;l�;5�;ќ�;T�;�g};?�r;�Uh;�^;&T;�J;�e@;;�6;2-;�M$;G;'j;Q�	;*;z��:0	�:���:9��:c.�:���:勒:%��:եi:��L:��/:�:'�9з9]-�9.M9J�-8?my� '�m_��I�������+)�V�A��Z�s�ز���ɑ�!Н��Ʃ�����q���bVͺ�ٺ���|� �������	�Bj��*����J� ��W&�",��1�k7��=���B��mH�}N���S�nhY��_���d�h`j��p��u��X{������T���(��e���ҋ�٦��;|��R���(�������  �  �=�*=Y�=�s==+�=`=�=� =CJ =g��<��<�d�<��<���<0�<�r�<���<���<k6�<v�<��<���<�/�<�k�<@��<���<0�<ZO�<��<���<���<F�<WN�<�|�<���<���<���<�$�<J�<�l�<Z��<a��<���<d��<��<��<5�<a#�<,�<1�<w2�<�/�<Y)�<��<y�<���<���<���<��<�}�<�Q�<7 �<$��<u��<j�<�!�<���<��<&�<P��<�`�<��<���<v�<���< �<)��<���<>e�<o͸<�0�<���<��<o=�<���<ڮ<�!�<�e�<��<}�<{�<$Q�<���<e��<R��<�
�<u2�<�W�<{{�<���<���<fڑ<���<e�<�*�<�B�<�Y�<Yo�<3��<��<c��<�{}<8�y<��u<��q<V	n<�+j<�Nf<�qb<��^<	�Z<��V<2S<�-O<tWK<a�G<S�C<-�?<Y<<�B8<2y4<v�0<��,<�.)<Tr%<�!<$<�V<|�<E<�g<�<�:<^�<'<eO�;G_�;�~�;���;���;�>�;���;F�;��;=�;5�;���;]��;��;���;��;\�;�5�;���;�;i};�r;1Vh;k^;� T;LJ;e@;u�6;A~-;L$;�E;�h;��	;?(;���:��:���:���:E+�:��:爒:���:Ţi:�L:��/:$�:�9yӷ9)4�9&_9]�-8��x���&��P��ΰ��L��	��)�j�A��Z��	s�V���pǑ��Ν��ũ�����܈��RVͺ�ٺ;�亯~��"�����X�	��k��,�`��8� �JY&��,�ɽ1�Sl7�^=�7�B�ynH��N��S�zhY�_�8�d��_j��p�&�u�6W{�����S��,(��X���2ы�쥎�z{��MQ���'��w����  �  ��=�*=_�=�s=="�=�_=�=� =-J =8��<��<rd�<֨�<���<�/�<yr�<s��<���<G6�<�u�<ɴ�<���<�/�<�k�<;��<���<U�<sO�<Q��<ι�<���<~�<�N�<}�<ߩ�<���<���<(%�<2J�< m�<���<|��<���<c��<��<��<1�<C#�<�+�<�0�<E2�<�/�<	)�<O�<=�<���<���<���<���<�}�<�Q�< �<��<r��<j�<�!�<���<��<<&�<w��<�`�<=��<ۃ�<��<ҏ�<i�<r��<��<xe�<�͸<�0�<*��<��<�=�<���< ڮ<�!�<�e�<���<[�<W�<Q�<���<-��<��<[
�<32�<�W�<9{�<���<X��<6ڑ<|��<:�<�*�<�B�<�Y�<Yo�<:��<B��<~��<F|}<��y<�u<�q<�	n<c,j<8Of<Xrb<�^<��Z<��V<}S<X.O<�WK<��G<m�C<+�?<O<<�B8<�x4<�0<��,<Z.)<�q%<~�!<�<QV<�<�<>g<��<(:<�<�&<�N�;�^�;H~�;���;o��;�>�;��;��;���;�=�;)�;���;6��;��;���;��;��;�6�;>��;��;:j};��r;Wh;J^;� T;�J;�d@;q�6;�|-;)K$;D;g;i�	;h&;���:}�:`��:y��:$(�:��:��:k��:Ӟi:A�L:L�/:<�:��9�ٷ9S;�9�p9�M.8��x���&�5E������k��y��)���A���Z��s�H����ő��̝�qĩ����������Wͺvٺ�����%�����&�	�n�h.�u��� �Y[&��,�3�1��m7�Z=���B�RoH�N�Y�S�zhY��_��d��^j�2p��u��U{��~���R��'��Z���Ћ�#����z��mP��:'�������  �  �=�*=a�=�s==�=�_=�=� =
J =���<W�<3d�<���<L��<�/�<9r�<C��<���<6�<�u�<���<���<�/�<�k�<I��<���<h�<�O�<���<��<,��<��<�N�<T}�<��<+��<:��<p%�<fJ�<2m�<���<���<���<i��<,��<��<�<##�<�+�<�0�<�1�<�/�<�(�<�<��<`��<G��<K��<���<�}�<lQ�<��<���<W��<�i�<	"�<���<%��<V&�<���< a�<m��<'��<��<)��<��<���<l��<�e�<θ<1�<e��<��<�=�<	��<ڮ<"�<�e�<ᥩ<<�<8�<�P�<W��<���<�ߞ<
�<�1�<�W�<�z�<s��<!��<�ّ<S��<�<~*�<�B�<�Y�<qo�<=��<S��<���<�|}<ؠy<��u<��q<A
n<-j<�Of<�rb<��^<�Z<x�V<�S<�.O<�WK<ւG<y�C<Y�?<L<<�B8<�x4<̱0<5�,<�-)<q%<�!<<�U<9�<W<�f<*�<�9<��<e&<N�;r^�;�}�;���;���;�>�;@��;	�;g��;>�;$�;���;[��;��;P��;<��;��;�7�;���;Q�;�k};d�r;�Wh;`^;�T;4J;�c@;c�6;�{-;�I$;�A;ee;��	;|$;�|�:?��:x��:���:�$�:|��:���:팃:��i:l�L:��/:�:v�9�޷9�@�9҅9+�.8�Lx���&�
5��D����w�x���(���A��}Z�< s������Ñ�[˝��é�F���ȇ��LYͺ0ٺ���6���(�������	�p�d0�4��=� �R]&��,���1�p7��=���B�&pH��N���S��gY��_�{�d��]j��p���u��S{��}���Q���%�������΋� ���oy��O���&�������  �  �=�*=o�=�s=	=�=�_=v=Ӧ =�I =���<�<�c�<G��<��<S/�<�q�<���<L��<�5�<�u�<���<���<�/�<rk�<V��<��<��<�O�<���<:��<a��<��<O�<�}�<j��<k��<{��<�%�<�J�<km�<э�<���<	��<���<��<��<�<#�<�+�<�0�<�1�<:/�<�(�<��<��<(��<���<��<B��<[}�<:Q�<��<���<G��<�i�<�!�<��<H��<|&�<���<7a�<���<_��<4�<m��< �<��<���<�e�<=θ<\1�<���<�<�=�<-��<$ڮ<�!�<�e�<ѥ�<)�<�<�P�<#��<���<�ߞ<�	�<�1�<=W�<�z�<1��<໓<�ّ<��<��<j*�<�B�<wY�<io�<U��<m��<���<�|}<^�y<�u<��q<�
n<�-j<JPf<{sb<�^<z�Z<��V<`S</O<5XK<�G<��C<X�?<#<<�B8<�x4<��0<��,<x-)<q%<��!<x<(U<Ѫ<�<&f<��<"9<�<�%<�M�;^�;�}�;G��;���;D?�;���;��;���;?�;��;���;B��; ��;���;+��;��;�8�;���;'�;�l};`�r;jXh;^;� T;�J;5c@;��6;Qz-;�G$;�@;+c;y�	;�!;�x�:���:U��:���:b �:�:���:[��:�i:�L:��/:d�:� �9�9;I�9B�9>/8��w���&�9%���|���b����(�p�A�KwZ��r�H�������qɝ�����M���Z����Yͺvٺ �����+������	�$r��2����\� ��_&��,���1�4q7�E=���B��pH�<N�+�S��gY��_���d��\j�}p���u��Q{��|���P���$��>����͋�����x���N��%��O����  �  ,�=�*=w�=�s=
=�=�_=i=�� =�I =���<��<�c�<���<���</�<�q�<���<��<�5�<yu�<q��<g��<~/�<rk�<a��<��<��<�O�<΅�<m��<���<F�<]O�<�}�<���<���<���<�%�<�J�<�m�<���<ث�<��<���<��<��<��<�"�<�+�<i0�<�1�<�.�<](�<��<p�<���<���<���<���<2}�<Q�<��<���<4��<j�<�!�<#��<R��<�&�<���<Ya�<���<���<��<���<F�<M��<���<Sf�<oθ<�1�<���<2�<�=�<8��<4ڮ<�!�<�e�<���<�<��<{P�<���<x��<^ߞ<�	�<k1�<�V�<wz�<���<���<�ّ<���<��<D*�<zB�<|Y�<jo�<j��<���<嫀<8}}<��y<Z�u<}�q<Xn<�-j<�Pf<�sb<��^<�Z<N�V<�S<Y/O<�XK<:�G<ԯC<`�?<)<<uB8<Zx4<^�0<h�,<,-)<�p%<
�!<<�T<K�<<�e<�<�8<ͫ<�%<"M�;t]�;�}�;4��;���;Z?�;���;7�;b��;�?�;��;���;/��;�;���;ޱ�;
�;Y9�;���;��;�m};d�r;�Xh;�^;� T;�J;�b@;��6;ky-;rF$;H?;�`;Ϭ	;�;~t�:Z��:J��:r��:��:1��:�}�:[��:�i:C�L:��/:�:e%�9��9EQ�9_�9�V/8�aw�+�&�L���o��mR�4���(�p�A��qZ���r�u���X����ǝ�:�������^����Yͺ�ٺ��亶��:.������	�zs�5������ �va&��,���1�pr7��=���B��qH��N��S��gY�E_��d�r[j�fp�c�u�zP{��{���O��$��(���͋�㡎��w���M���$�������  �  6�=�*=x�=�s=	=�=�_=Z=�� =�I =[��<��<|c�<˧�<���<�.�<�q�<���<���<}5�<Xu�<U��<Z��<i/�<tk�<d��<��<��<�O�<���<���<���<t�<�O�<~�<��<���<���<&�<K�<�m�<!��<��<#��<���< ��<��<��<�"�<^+�<?0�<v1�<�.�<%(�<U�<:�<���<���<���<֣�<�|�<�P�<��<���<(��<�i�<"�<)��<e��<�&�<&��<�a�<��<τ�<��<��<��<���<)��<�f�<�θ<�1�<돵<P�<>�<G��<=ڮ<�!�<�e�<���<��<��<KP�<ǂ�<M��<ߞ<U	�<(1�<�V�<Bz�<ě�<w��<hّ<���<��<1*�<hB�<rY�<po�<j��<���<���<�}}<��y<��u<��q<�n<m.j<QQf<atb<�^<r�Z<��V<S<�/O<�XK<e�G<ٯC<m�?<%<<QB8<9x4<"�0<)�,<�,)<.p%<��!<�<&T<��<�<?e<��<Q8<Y�<N%<�L�;/]�;%}�;,��;���;i?�;;��;|�;
��;f@�;P�;U��;畬;ڈ�;p��;ز�;��;$:�;M��;K �;�n};�r;Yh;�^;� T;NJ;b@;��6;Ex-;E$;b=;�_;�	;R;q�:���:���:���:c�:���:{�:��:ʐi:gL:��/:��:�%�9��9/W�9��9��/8@w��g&�o�� `��/D���c�(���A�]kZ���r���������0Ɲ�����@�������ZͺF ٺ���	��\1�����c�	�yu��6����:� �"c&�,,�9�1�?t7��=���B�{rH�AN�M�S��gY�C_���d��Zj�p��u��N{�{���N��#��8���̋�2����v��M��9$������  �  =�=�*={�=�s== �=�_=F=�� =�I =?��<z�<Jc�<���<n��<�.�<Tq�<h��<���<i5�<Gu�<0��<V��<b/�<ok�<c��</��<��<P�<��<���<���<��<�O�<C~�<��<��<��<6&�<%K�<�m�<.��<���<>��<���<)��<��<��<�"�<B+�<90�<W1�<�.�<�'�<(�<�<���<`��<s��<���<�|�<�P�<q�<���<(��<�i�<	"�<)��<��<�&�<4��<�a�<>��<���<��<��<��<���<]��<�f�<�θ<�1�<��<`�< >�<]��<>ڮ<�!�<�e�<���<��<��<:P�<���<,��<�ޞ<7	�<1�<�V�<z�<���<Z��<Lّ<���<��<!*�<cB�<kY�<vo�<l��<���<��<�}}<6�y<
�u</�q<n<�.j<�Qf<�tb<[�^<��Z<�V<>S<�/O<�XK<��G<�C<r�?<<<HB8< x4<Ӱ0<�,<~,)<�o%<N�!<-<�S<i�<l<�d<Y�<8<*�<'%<L�;]�;�|�;��;���;�?�;{��;��;���;�@�;��;ƹ�;���;���;֒�;���;&�;�:�;ɡ�;� �;'o};r�r;�Yh;j^;"T;�J;�a@;0�6;Vw-;�D$;\<;�^;n�	;�;In�:���:���:���:��:���:nz�:���:�i:L:��/:z�:0%�9i�97Z�9^�9��/8��v�'R&������S��<�}��R�(��A��eZ�m�r�w���޻��Gŝ�L���O���c���{[ͺz ٺ�����2�����w�	� w��7�%��^� ��d&��,�!�1�u7�2 =���B� sH�eN���S��gY�6_���d�gZj�P p�6�u��M{��z��bN��G"������Lˋ�����=v��vL���#�������  �  H�=�*=��=�s==��=�_=C=�� =�I =��<d�<;c�<���<Q��<�.�<Iq�<M��<���<U5�<-u�<&��<D��<d/�<qk�<k��<6��<��<)P�<*��<ɺ�<���<��<�O�<U~�<��<"��<A��<K&�<<K�<�m�<C��<��<A��<���<'��<��<��<�"�<3+�<0�<A1�<�.�<�'�<�<��<c��<H��<h��<���<�|�<�P�<^�<���<��<�i�<	"�<5��<���<�&�<L��<�a�<Y��<��<�<5��<��<φ�<y��<�f�<�θ<�1�<#��<{�<->�<e��<Jڮ<�!�<�e�<���<��<��<$P�<���<��<�ޞ<	�<�0�<zV�< z�<���<8��<8ّ<���<��<*�<\B�<kY�<uo�<v��<���<��<�}}<d�y</�u<f�q<Wn<�.j<�Qf<�tb<��^<��Z<(�V<qS<
0O<YK<��G<��C<y�?<<<AB8<�w4<İ0<��,<Y,)<�o%<!�!<<�S<.�<"<�d< �<�7< �<�$<�K�;�\�;�|�;��;���;�?�;���;�;���;"A�;�;Q��;��;Ɖ�;A��;ٳ�;��;
;�;��;!�;�o};��r;�Yh;�^;T;J;na@;��6;�v-;�C$;�;;�];�	;7;$l�:���:���:���:m�:��:�x�:Y��:��i:}L:t�/:D�:�'�9V�9�^�9��9V 08˜v��G&�􆹁N���5�U��(�(�R�A��cZ��r�]���R����ĝ������J���<[ͺ�!ٺQ��}���3��~��f�	�w��8����� �7e&�.,�6�1��u7�!=��B��sH��N�~�S��gY��_���d��Yj���o�|�u�-M{�z���M���!��^���ˋ�ퟎ��u��3L��l#��v����  �  ��=�-=��=[w=�=Y�=xd=r=(� =�O =��<D,�<r�<b��<H��<�@�<���<���<�
�<�L�<֍�<R��<��<�L�<��<���<��<(<�<!u�<׬�<3��<-�<�K�<�}�<��<���<�	�<5�<?^�<U��<:��<���<���<E
�<�$�<�<�<zQ�<�b�<q�<�{�<܂�<M��<ą�</��<�x�<mk�<�Y�<�C�<�(�<��<���<5��<V��<�S�<m�<;��<��<�B�<;��<���<�5�<��<d�< ��<�y�<���<Jx�<��<�_�<?˺<i1�<Z��<G�<=E�<��<.�<_.�<]s�<O��<6�<�*�<L`�<���<(¢<��<R�<�?�<Od�<톙<���<%ƕ<�<2��<��<�/�<�F�<=\�<�p�<���<	��<p��<��<P�}<g�y<��u<_�q<�n<�%j<WCf<�`b<^<��Z<½V<��R<� O<$K<IG<�oC<��?<��;<�7<� 4<�S0<��,<n�(<� %<.B!<�<��<b"<vw<G�<3<�<�<| <���;��;}�;
1�;rg�;���;�	�;�v�;���;��;07�;��;�̪;﹤;Y��;�٘;�;�Z�;g��;�<�;�y;�o;��d;�QZ;�AP;�aF;^�<;`-3;��);� ;��;f�;�=;F��:(��:z�:Yh�:ל�:��:4қ:wʌ: |:#�^:%B:��%:L�	:�M�9���9�z_9Cw�8��27Wź�O�D�����v�ȹ�����h��1/�N�G�l6`��{x�?M��5L��\:�����W췺ʱú0kϺ6ۺ
��;]�����W���|
��8��������T!�2'���,��Q2��7�2�=��9C���H�dxN�<T�Q�Y��T_���d���j� 2p���u��q{�.����Y���*��q���2͋�����:q��AD��.���왻�  �  ��=�-=��=bw=�=K�=xd=p=2� =�O =��<T,�<r�<|��<_��<�@�<���<���<�
�<�L�<��<K��<��<kL�<��<���<��<3<�<%u�<Ԭ�<'��<�<�K�<�}�<	��<���<�	�<�4�<-^�<E��<1��<���<���<I
�<�$�<�<�<`Q�<�b�<q�<�{�<���<O��<҅�<A��<�x�<�k�<	Z�<�C�<�(�<��<���<L��<U��<�S�<_�< ��<���<�B�<9��<���<�5�<��<�c�<���<�y�<���<#x�<��<�_�<$˺<Z1�<M��<A�<EE�<���<+�<g.�<`s�<3��<2�<�*�<S`�<В�<+¢<��<^�<�?�<ld�<��<���<5ƕ<�<2��<��<�/�<�F�<$\�<zp�<˃�<��<{��<"��<[�}<W�y<��u<(�q<�n<�%j<	Cf<�`b<�~^<ŝZ<��V<u�R<� O<$K< IG<�oC<��?<��;<��7<� 4<�S0<�,<o�(<� %<NB!<-�<��<�"<�w<b�<,3<!�<�<3| <y��;y��;�;�0�;�g�;���;�	�;
w�;���;׌�;�6�;���;�̪;���;���;�٘;��;NZ�;+��;�<�;]�y;o;��d;-RZ;BP;�`F;¯<;-3;w�);Ӱ ;�;��;u>;��:Z��:0|�:2i�:���:��:Nқ:�ˌ:��{:��^:�B::�%:�	:�O�9&��9_9��8�527Ӻ��D�F����ȹ����.l��2/���G�18`�c}x��M���K���9������뷺��ú�lϺwۺ����\�����<��2|
�T8��������S!�� '�q�,�_Q2�
�7�s�=��9C���H�)yN��T�׵Y��T_�Y�d���j��1p���u�@r{�����Z���*�����b͋�4����q��yD��S���왻�  �  v�=�-=��=_w=�=X�=�d=w=?� =�O =1��<u,�<7r�<���<s��<�@�<���<��<�
�<�L�<���<]��<��<~L�<��<���<��<<�<u�<���<
��<�<yK�<�}�<��<���<�	�<�4�<^�<0��<��<���<���<2
�<�$�<�<�<iQ�<
c�<8q�<�{�<��<b��<��<b��<�x�<�k�< Z�<�C�<�(�<	�<���<g��<b��<�S�<��<&��<��<�B�<!��<���<�5�<���<�c�<���<�y�<���<x�<��<�_�<˺<=1�<2��<!�<&E�<q��<�<Y.�<^s�<?��<Y�<�*�<d`�<璤<@¢<��<|�<�?�<}d�<&��<���<Uƕ<(�<F��<��<�/�<�F�<A\�<�p�<Ń�<���<j��<��<,�}<�y<b�u<��q<Bn<�%j<�Bf<�`b<�~^<��Z<t�V<:�R<f O<�#K<�HG<�oC<��?<��;<	�7<2!4<�S0<�,<��(<%<�B!<e�<�<�"<�w<��<t3<X�<�<b| <���;.��;X�;1�;�g�;]��;�	�;�v�;t��;k��;�6�;*��;`̪;G��;X��;�٘;I�;�Y�;ᾇ;b<�;��y;o;�d;�QZ;�AP;QaF;�<;7.3;��);�� ;��;��;�?;���:���:�}�:�j�:͟�:��:�ӛ:�͌:�|:��^:vB:P�%:��	:VK�9߱�9�r_9�k�8z617庸��D�iÕ���ȹg���o�6/�}�G��;`�u�x�aO��fM��;������췺��úlϺ�ۺF�溔[�s������"{
�_7���)���R!� '�p�,�~P2�k�7���=�_9C���H�IxN��T��Y�8U_���d�w�j��2p���u��r{�
����Z��7+��y����͋�����!r���D�����M홻�  �  m�=�-=��=Xw=�=\�=�d=�=N� =�O =e��<�,�<|r�<׷�<���<$A�< ��<C��<�
�<�L�<��<}��<��<�L�<��<���<��<<�<�t�<���<���<��<QK�<@}�<���<s��<k	�<�4�<�]�<��<��<���<���<5
�<�$�<�<�<Q�< c�<@q�<|�<-��<���<��<���<�x�<�k�<[Z�<8D�<7)�<+	�<��<���<���<�S�<v�<<��<��<�B�<&��<r��<�5�<���<�c�<���<�y�<~��<�w�<K�<>_�<�ʺ<�0�<	��<��<E�<Y��<�<V.�<Ts�<O��<K�<�*�<�`�<��<v¢<��<��<�?�<�d�<b��<�<�ƕ<Y�<���<
�<$0�<�F�<C\�<�p�<���<��<`��<���<�}<ͮy<��u<��q<�n<�$j<]Bf<�_b<E~^<)�Z<��V<��R< O<�#K<�HG<�oC<��?<��;<�7<%!4<1T0<\�,<	�(<n%<�B!<�<��<P#<kx<'�<�3<˚<Q<�| <Z��;��;��;&1�;�g�;���;w	�;av�;��;ዽ;�5�;���;[˪;/��;���;Pؘ;��;�X�;5��;�;�;��y;�o;9�d;�QZ;�AP;bF;��<;�.3;^�);�� ;��;3�;�A;g��:���:���:jo�:��:x�:Vכ:�ό:&|:��^:�B:M�%:H�	:M�9���9�h_9�L�8�J07���;E��˕�<�ȹ�����w��?/�1�G��C`��x�\Q���N��J<��M���췺�ú�jϺ�ۺ���;Y����ǹ��y
�^5������Q!���&�˧,��N2���7���=��7C���H�;xN�T�s�Y�U_�4�d��j��3p�$�u��t{�Ԋ��N[��z,��`����΋�}����r���E��d���홻�  �  \�=�-=��=Tw=�=h�=�d=�=b� =�O =���<�,�<�r�<��<��<aA�<H��<���<.�<M�<C��<���<�<�L�<��<��<��<�;�<�t�<Z��<���<��<K�<}�<d��<0��<"	�<r4�<�]�<΄�<���<]��<���<
�<�$�<�<�<�Q�<c�<aq�<?|�<Y��<܆�<W��<ށ�<-y�<&l�<�Z�<sD�<t)�<g	�<I��<���<���<T�<��<L��<ݏ�<�B�<���<I��<{5�<|��<{c�<;��<My�<3��<|w�<�<�^�<�ʺ<�0�<Ց�<��<�D�<(��<��<C.�<Ps�<a��<a�<�*�<�`�<:��<�¢</�<��<0@�<e�<���<3��<�ƕ<��<���<3�<U0�<�F�<\\�<�p�<���<땄<2��<з�<z�}<w�y<��u<��q<kn<a$j<�Af<`_b<�}^<��Z<|�V<��R<��N<]#K<HG<�oC<��?<��;<J�7<V!4<�T0<��,<v�(<�%<~C!<��< �<�#<�x<��<Z4<W�<�<
} <"��;���;�;91�;dg�;��;��;�u�;��;M��;�4�;���;�ʪ;0��;���;=ט;��;�W�;o��;;�;L�y;�o;�d;eQZ;�AP;�bF;u�<;�/3;��);� ;��;*�;�C;:��:��:/��:<s�:��:a �:�ۛ:�Ҍ:�|:Z�^:� B:��%:�	:�H�9Z��9�V_92!�8Pl.7�C���;E��ڕ���ȹ��,��-G/�R�G�LL`�Ҋx�mU��IQ��?�����h��úoiϺ�ۺѻ溒V���������w
�63�	�����O!���&���,�M2���7�i�=�x6C���H�uwN��T���Y��U_���d�%�j�y5p�{�u��v{����D\���-��g���Ћ�u���t���F������  �  H�=w-=|�=Xw=�=p�=�d=�=�� =P =���<=-�<s�<u��<Z��<�A�<���<���<p�<]M�<z��<���<=�<�L�<��<���<��<�;�<�t�<��<j��<M�<�J�<�|�<
��<���<��<4�<I]�<���<p��<+��<c��<�	�<�$�<�<�<�Q�<Cc�<�q�<V|�<���<��<���<1��<�y�<�l�<�Z�<�D�<�)�<�	�<x��<��<׉�<"T�<��<<��<��<lB�<���<&��<F5�<1��<-c�<���<�x�<���<w�<��<�^�<!ʺ<m0�<��<r�<�D�<	��<��<8.�<Us�<W��<��<�*�<�`�<~��<�¢<��<N�<�@�<be�<���<���<!Ǖ<��<���<w�<h0�<G�<x\�<�p�<���<ו�<!��<���<�}<ԭy<�u<d�q<�n<�#j<Af<�^b<�|^<��Z<�V<��R<0�N<
#K<[HG<loC<��?<��;<k�7<�!4<�T0<6�,<��(<�%<.D!<1�<��<�$<�y<l�<5<�<W	<�} <���;c��;=�;o1�;g�;ݮ�;��;Gu�;:��;$��;�3�;-�;-ɪ;ߵ�;'��;֘;G
�;�V�;o��;:�;ءy;� o;f�d;�PZ;
BP;obF;��<;�03;��);_� ;D�;��;5F;���:��:��:�x�:H��:�%�:�ޛ:�֌:�|:V�^:�&B:q�%:v�	:�D�9���9�G_9���8#A,7����XE�����>�ȹb#������Q/�s�G�`S`���x�QY��
T���@��$����F�ú�iϺ�ۺ��溏S�q���ҵ�)u
��0�<���� L!���&��,��J2��7�I�=��5C���H��vN��T�U�Y�_V_�0�d�U�j�%7p��u�vx{�����]���.������Nы� ���.u���G��H����  �  +�=j-=n�=Tw==v�=�d=�=�� =5P =;��<�-�<ls�<ո�<���<$B�<��<-��<��<�M�<Î�<���<b�<�L�<.��<n��<��<�;�<mt�<��<��<��<\J�<U|�<���<n��<��<�3�<�\�<(��<B��< ��<,��<�	�<�$�<�<�<�Q�<Wc�<�q�<�|�<��<O��<���<}��<�y�<�l�<U[�<.E�<*�<
�<���<6��<��<HT�<��<D��<��<QB�<���<��<5�<��<�b�<���<zx�<���<�v�<;�<E^�<�ɺ<0�<��<P�<oD�<ݖ�<��<.�<`s�<\��<��<+�<a�<���<2â<��<��<�@�<�e�<\��<娗<oǕ<4�<1��<��<�0�<BG�<�\�<�p�<���<���<��<r��<Ɏ}<R�y<H�u<��q<�n<#j<D@f<
^b<B|^<W�Z<K�V<Y�R<��N<�"K<"HG<3oC<~�?<��;<��7<"4<-U0<Ƌ,<p�(<$%<�D!<�<��<V%<�z<�<�5<~�<�	< ~ <f��;��;�;�1�;Qg�;���;.�;�t�;���;;�2�;�;�Ǫ;���;���;�Ԙ;��;�U�;���;[9�;��y;"�n;�d;CPZ;�BP;�bF;��<;@23;��);и ;b�;��;�H;M��:���:���:F�:N��:+�:��:zی:�|:��^:*B:�%:��	:B?�9���9�._9��8��*7W컸~E������ȹ�;��A��K\/���G��\`�ßx��Z��cW���B��2��ﷺ0�úiϺ�ۺ���O��������r
�!.����!��2I!�&�&���,�H2��7���=��3C�0�H�/vN�T�T�Y�9W_���d��j�>8p��u�Z{{�U���Z_��*0������ҋ�p���iv��I��p��$��  �  �=V-=i�=Lw==��=�d=�=�� =\P =���<�-�<�s�<.��<��<yB�<G��<z��<�<�M�<��<'��<v�<�L�<*��<c��<��<};�<-t�<���<���<��<J�<�{�<T��<��<�<Z3�<�\�<��<��<���<���<�	�<�$�<�<�<�Q�<ec�<�q�<�|�<��<���<H��<Ђ�<;z�<8m�<�[�<~E�<e*�<S
�<��<X��<F��<sT�<��<V��<ُ�<?B�<���<���<�4�<���<}b�<O��<"x�<��<Ov�<��<�]�<rɺ<�/�<א�<��<&D�<���<��<.�<Qs�<n��<��<D+�<Ba�<瓤<�â<�<��<=A�<f�<���<;��<�Ǖ<��<���<��<�0�<bG�<�\�<�p�<���<���<概<?��<7�}<߬y<��u<�q<:n<I"j<�?f<E]b<�{^<��Z<��V<��R<_�N<)"K<�GG<oC<]�?<��;<��7<;"4<�U0<�,<�(<�%<{E!<��<c�<2&<6{<��<d6<E�<Y
<u~ <]��;w��;��;�1�;<g�;~��;��;�s�;���;��;�1�;��;�ƪ;3��;[��;bӘ;��;�T�;��;j8�;��y;��n;1�d;PZ;BP;�cF;D�<;�33;��);ʹ ;H�;��;ZK;���:���:З�:���:���:�/�:��:�݌:h |:��^:�+B:��%:w�	:9<�9��9�_9�~�8��(7�.��֧E������ȹ�Q��x��ih/�n�G�zg`��x��_���[��E��a ���ﷺʰú�gϺ�ۺ�溚L�u������,p
�E+�t����iF!�q�&��,�}E2���7� �=�N2C�6�H�yuN�T��Y��W_��d���j��:p���u��}{������`���1�����5ԋ�å���w��;J��W��=��  �  �=?-=c�=Kw==��=�d=�=Ӭ =�P =���</.�<'t�<��<y��<�B�<���<���<U�<#N�<��<M��<��<�L�<��<k��<s�<U;�<t�<r��<���<Z�<�I�<�{�<���<���<��<	3�<T\�<���<���<���<���<�	�<�$�<�<�<�Q�<zc�<�q�<�|�<E��<���<���<;��<�z�<�m�<\�<�E�<�*�<�
�<\��<���<p��<�T�<��<`��<ɏ�<EB�<o��<���<�4�<j��<Db�<���<�w�<���<�u�<t�<z]�<ɺ<c/�<���<��<
D�<���<s�<.�<@s�<��<��<b+�<ra�<1��<�â<X�<`�<�A�<{f�<��<���<ȕ<��<���<�<	1�<xG�<�\�<�p�<���<���<���<-��<ō}<T�y<,�u<t�q<�n<�!j<�>f<�\b<�z^<��Z<�V<[�R<��N<�!K<oGG<oC<V�?<��;<��7<^"4<�U0<z�,<��(<O%< F!<f�<�<�&<�{<��<�6<Ν<<�~ <
��;���;k�;�1�;tg�;��;�;ts�;���;B��;q0�;��;@Ū;˱�;��;Ҙ;��;\S�;4��;[7�;Y�y;H�n;ɍd;`PZ;�AP;�cF; �<;w43;-�);ڻ ;��;��;�N;��:���:���:���:���:r3�:��:�:&&|:�^:�.B:��%:�	:�>�9ٌ�9�_9�[�8@�&7a����E�4��2	ɹ�h��c���s/�	H��q`�v�x�7d���\���G���"��ﷺ��úCfϺ�ۺ��iI�������;n
��'������C!���&�?�,��C2�	�7�4�=��0C���H��tN�T��Y��W_���d�K�j�Q<p� �u��{������a��03��,���Ջ����y��bK��^��A��  �  �=3-=W�=Hw==��=�d=
	=� =�P =	��<x.�<et�<ǹ�<���<C�<��<
��<��<PN�<O��<q��<��<�L�<%��<]��<[�<:;�<�s�<I��<e��<�<vI�<_{�<���<o��<��<�2�<\�<g��<���<`��<���<y	�<�$�<�<�<�Q�<�c�<r�<!}�<���<'��<ć�<y��<�z�<�m�<O\�<F�<+�<�
�<���<Ժ�<���<�T�<�<m��<Ǐ�<+B�<T��<p��<f4�<4��<�a�<���<�w�<u��<�u�<+�<7]�<�Ⱥ< /�<X��<~�<�C�<\��<Y�<�-�<?s�<���<��<�+�<�a�<`��<Ģ<��<��<�A�<�f�<O��<ҩ�<`ȕ< �<���<Y�<-1�<�G�<�\�<�p�<���<���<���<���<w�}<�y<��u<��q<n<!j<N>f<\b<^z^<y�Z<��V<��R<��N<�!K<>GG<�nC<I�?<��;<�7<�"4<9V0<�,<�(<�%<�F!<�<��<}'<m|<5�<�7<D�<g<X <���;���;��;�1�;Qg�;ͭ�;��;�r�;J��;p��;�/�;��;VĪ;ڰ�;촞;-ј;��;hR�;.��;�6�;	�y;�n;�d;�OZ;�AP;�dF;i�<;�53;��);� ;a�;�;�P;է�:���:ˡ�:ʍ�:rº:�7�:��:��:�+|:��^:E4B:��%:>�	:�9�9��9��^9-)�8�%7������E�iD���ɹ�{�����v{/��H��y`�8�x��f���_���I��R$���U�ú�dϺ�ۺί�xF�x������k
�&�������A!���&��,��A2���7�I�=��/C�+�H��sN��T��Y�gX_�Y�d���j��=p���u�ǁ{�����c��'4��`���֋�'���z��_L��/�����  �  ܇=7-=Q�=Ew==��=�d=	=� =�P =I��<�.�<�t�<��<���<]C�<��<@��<��<wN�<s��<���<��<�L�<3��<K��<[�<8;�<�s�<*��<*��<��<?I�<{�<x��<,��<@�<�2�<�[�<-��<e��<:��<���<�	�<z$�<�<�<�Q�<�c�<.r�<:}�<���<J��<��<���<{�<n�<�\�<^F�<++�<�<���<��<���<�T�<�<e��<Ώ�<B�<]��<Z��<:4�<��<�a�<���<<w�<(��<Xu�<��<�\�<�Ⱥ<�.�<��<\�<�C�<R��<Z�<�-�<Ks�<���<��<�+�<�a�<���</Ģ<��<��< B�<�f�<���<��<�ȕ<A�<# �<{�<?1�<�G�<�\�<�p�<���<���<���<ݶ�<1�}<��y<?�u<��q<~n<� j<�=f<�[b<�y^<�Z<1�V<��R<F�N<O!K<MGG<�nC<<�?< �;<�7<�"4<\V0<;�,<T�(<M%<G!<Y�<B�<�'<}<��<	8<��<�<� <��;���;��;:2�;g�;߭�;��;r�;���;���;�.�;��;@ê;���;�;&И;��;�Q�;S��;$6�;�y;_�n;��d;-OZ;=BP;�dF;1�<;�63;Y�);�� ;��;"�;�Q;٬�:	�:Х�:��:�ĺ:-<�:m�:��:F/|:��^:)3B:�%:��	:�3�9:��9��^9h �8�1$7�Ἰ�F�dU���*ɹI���!����/��H�=`�|�x��h���b��4J���#��a�S�ú|eϺ�ۺ���DD�<���f���i
��$�?��-��-?!���&���,��?2���7�>�=�D/C���H�tN��T�/�Y��X_��d�˜j��>p��u�q�{�����d��5�����׋�9����z��-M�����^��  �  Շ=!-=E�=Bw==��= e="	=� =�P =`��<�.�<�t�<*��<��<tC�<7��<\��<��<�N�<���<���<��<M�<7��<B��<=�<;�<�s�<��<��<��<I�<�z�<]��<��<&�<c2�<�[�<��<K��<)��<���<\	�<p$�<�<�<�Q�<�c�<Er�<T}�<Ä�<a��<!��<���<0{�<-n�<�\�<tF�<M+�<-�<���<��<ˊ�<�T�<�<s��<Џ�<B�<2��<<��<(4�<���<�a�<_��<w�<��<@u�<��<�\�<lȺ<�.�<��<?�<�C�<+��<5�<�-�<Ls�<���<��<�+�<�a�<���<DĢ<��<��<5B�<g�<���</��<�ȕ<W�<A �<��<^1�<�G�<�\�<�p�<���<t��<|��<Ͷ�<�}<d�y<	�u<P�q<Cn<T j<�=f<K[b<�y^<ԘZ<��V<Y�R<�N<0!K<�FG<�nC</�?<�;</�7<�"4<�V0<i�,<��(<}%<OG!<��<n�<-(<D}<��<C8<�<�<� <|��; ��;+�;U2�;g�;p��;2�;�q�;��;O��;x.�;i�;�ª;���;���;�Ϙ;!�;UQ�;	��;�5�;q�y;��n;G�d;�NZ;QBP;�dF;ʶ<;T73;2�);�� ;H�;��;�R;y��:��:z��:o��:�ƺ:�=�:���:��:�2|:��^:�5B:�%:�	:�1�9��9��^9=��8*Z#7�����F��]���0ɹ����a����/��H���`�տx�lj���c��wL��&����'�ú/dϺuۺԬ溩B�S������i
��#����O��w>!���&�͖,�?2���7�v�=�P.C���H�jsN�LT�V�Y��Y_�h�d�Q�j�W?p���u�E�{�7���d���5�����؋�����V{���M��T �����  �  ׇ=!-=S�=Hw=
=��=�d=!	=� =�P =n��<�.�<�t�<8��<6��<{C�<I��<u��<��<�N�<���<���<��< M�<(��<X��<V�<;�<�s�<���<��<��<I�<�z�<>��<���<�<W2�<�[�<��<8��<#��<���<a	�<�$�<�<�<�Q�<�c�<9r�<I}�<Ʉ�<l��<0��<փ�<6{�<Nn�<�\�<xF�<f+�<<�<���<��<���<�T�<�<j��<���<!B�<;��<F��<&4�<���<�a�<N��<
w�<���<u�<��<�\�<YȺ<�.�<���<$�<�C�<1��<K�<�-�<:s�<���<��<�+�<�a�<���<TĢ<�<��<9B�<6g�<É�<8��<�ȕ<e�<M �<��<\1�<�G�<�\�<�p�<���<���<��<Ӷ�<�}<X�y<�u<0�q<,n<" j<e=f<[b<�y^<��Z<�V<U�R<��N<8!K<�FG<�nC<D�?<��;<'�7<�"4<�V0<e�,<��(<�%<�G!<��<��<|(<T}<��<x8<�<<� <l��;���;�;2�;^g�;֭�;C�;r�;��;N��;W.�;(�;�ª;��;3��;xϘ;��;Q�;���;{5�;I�y;��n;u�d;�OZ;BP;�dF;�<;�63;��);*� ;��;z�;�S;Ԯ�:��:ʩ�:���:bȺ:�>�:l��:��:�0|:t�^:76B:�%:P�	:�8�9���9F�^9=��8��"7+���{F��`���4ɹ5������c�/��H�S�`�I�x�l��ec��
L���$��X�;�ú�dϺ�ۺc��zC�����2��nh
�8#�l�����=!�|�&��,��>2�B�7�t�=�c.C�W�H�lsN��T� �Y��X_�W�d��j��?p���u�\�{�x����d���5��-���؋�ԩ���{���M��] ������  �  Շ=!-=E�=Bw==��= e="	=� =�P =`��<�.�<�t�<*��<��<tC�<7��<\��<��<�N�<���<���<��<M�<7��<B��<=�<;�<�s�<��<��<��<I�<�z�<]��<��<&�<c2�<�[�<��<K��<)��<���<\	�<p$�<�<�<�Q�<�c�<Er�<T}�<Ä�<a��<!��<���<0{�<-n�<�\�<tF�<M+�<-�<���<��<ˊ�<�T�<�<s��<Џ�<B�<2��<<��<(4�<���<�a�<_��<w�<��<@u�<��<�\�<lȺ<�.�<��<?�<�C�<+��<5�<�-�<Ls�<���<��<�+�<�a�<���<DĢ<��<��<5B�<g�<���</��<�ȕ<W�<A �<��<^1�<�G�<�\�<�p�<���<t��<|��<Ͷ�<�}<d�y<	�u<P�q<Cn<T j<�=f<K[b<�y^<ԘZ<��V<Y�R<�N<0!K<�FG<�nC</�?<�;</�7<�"4<�V0<i�,<��(<}%<OG!<��<n�<-(<D}<��<C8<�<�<� <|��; ��;+�;U2�;g�;p��;2�;�q�;��;O��;x.�;i�;�ª;���;���;�Ϙ;!�;UQ�;	��;�5�;q�y;��n;G�d;�NZ;QBP;�dF;ʶ<;T73;2�);�� ;H�;��;�R;y��:��:z��:o��:�ƺ:�=�:���:��:�2|:��^:�5B:�%:�	:�1�9��9��^9=��8*Z#7�����F��]���0ɹ����a����/��H���`�տx�lj���c��wL��&����'�ú/dϺuۺԬ溩B�S������i
��#����O��w>!���&�͖,�?2���7�v�=�P.C���H�jsN�LT�V�Y��Y_�h�d�Q�j�W?p���u�E�{�7���d���5�����؋�����V{���M��T �����  �  ܇=7-=Q�=Ew==��=�d=	=� =�P =I��<�.�<�t�<��<���<]C�<��<@��<��<wN�<s��<���<��<�L�<3��<K��<[�<8;�<�s�<*��<*��<��<?I�<{�<x��<,��<@�<�2�<�[�<-��<e��<:��<���<�	�<z$�<�<�<�Q�<�c�<.r�<:}�<���<J��<��<���<{�<n�<�\�<^F�<++�<�<���<��<���<�T�<�<e��<Ώ�<B�<]��<Z��<:4�<��<�a�<���<<w�<(��<Xu�<��<�\�<�Ⱥ<�.�<��<\�<�C�<R��<Z�<�-�<Ks�<���<��<�+�<�a�<���</Ģ<��<��< B�<�f�<���<��<�ȕ<A�<# �<{�<?1�<�G�<�\�<�p�<���<���<���<ݶ�<1�}<��y<?�u<��q<~n<� j<�=f<�[b<�y^<�Z<1�V<��R<F�N<O!K<MGG<�nC<<�?< �;<�7<�"4<\V0<;�,<T�(<M%<G!<Y�<B�<�'<}<��<	8<��<�<� <��;���;��;:2�;g�;߭�;��;r�;���;���;�.�;��;@ê;���;�;&И;��;�Q�;S��;$6�;�y;_�n;��d;-OZ;=BP;�dF;1�<;�63;Y�);�� ;��;"�;�Q;٬�:	�:Х�:��:�ĺ:-<�:m�:��:F/|:��^:)3B:�%:��	:�3�9:��9��^9h �8�1$7�Ἰ�F�dU���*ɹI���!����/��H�=`�|�x��h���b��4J���#��a�S�ú|eϺ�ۺ���DD�<���f���i
��$�?��-��-?!���&���,��?2���7�>�=�D/C���H�tN��T�/�Y��X_��d�˜j��>p��u�q�{�����d��5�����׋�9����z��-M�����^��  �  �=3-=W�=Hw==��=�d=
	=� =�P =	��<x.�<et�<ǹ�<���<C�<��<
��<��<PN�<O��<q��<��<�L�<%��<]��<[�<:;�<�s�<I��<e��<�<vI�<_{�<���<o��<��<�2�<\�<g��<���<`��<���<y	�<�$�<�<�<�Q�<�c�<r�<!}�<���<'��<ć�<y��<�z�<�m�<O\�<F�<+�<�
�<���<Ժ�<���<�T�<�<m��<Ǐ�<+B�<T��<p��<f4�<4��<�a�<���<�w�<u��<�u�<+�<7]�<�Ⱥ< /�<X��<~�<�C�<\��<Y�<�-�<?s�<���<��<�+�<�a�<`��<Ģ<��<��<�A�<�f�<O��<ҩ�<`ȕ< �<���<Y�<-1�<�G�<�\�<�p�<���<���<���<���<w�}<�y<��u<��q<n<!j<N>f<\b<^z^<y�Z<��V<��R<��N<�!K<>GG<�nC<I�?<��;<�7<�"4<9V0<�,<�(<�%<�F!<�<��<}'<m|<5�<�7<D�<g<X <���;���;��;�1�;Qg�;ͭ�;��;�r�;I��;o��;�/�;��;VĪ;ڰ�;촞;-ј;��;hR�;.��;�6�;	�y;�n;�d;�OZ;�AP;�dF;i�<;�53;��);� ;a�;�;�P;է�:���:ˡ�:ʍ�:rº:�7�:��:��:�+|:��^:E4B:��%:>�	:�9�9��9��^9-)�8�%7������E�iD���ɹ�{�����v{/��H��y`�8�x��f���_���I��R$���U�ú�dϺ�ۺί�xF�x������k
�&�������A!���&��,��A2���7�I�=��/C�+�H��sN��T��Y�gX_�Y�d���j��=p���u�ǁ{�����c��'4��`���֋�'���z��_L��/�����  �  �=?-=c�=Kw==��=�d=�=Ӭ =�P =���</.�<'t�<��<y��<�B�<���<���<U�<#N�<��<M��<��<�L�<��<k��<s�<U;�<t�<r��<���<Z�<�I�<�{�<���<���<��<	3�<T\�<���<���<���<���<�	�<�$�<�<�<�Q�<zc�<�q�<�|�<E��<���<���<;��<�z�<�m�<\�<�E�<�*�<�
�<\��<���<p��<�T�<��<`��<ɏ�<EB�<o��<���<�4�<j��<Db�<���<�w�<���<�u�<t�<z]�<ɺ<c/�<���<��<
D�<���<s�<.�<@s�<��<��<b+�<ra�<1��<�â<X�<`�<�A�<{f�<��<���<ȕ<��<���<�<1�<xG�<�\�<�p�<���<���<���<-��<ō}<T�y<,�u<t�q<�n<�!j<�>f<�\b<�z^<��Z<�V<[�R<��N<�!K<oGG<oC<V�?<��;<��7<^"4<�U0<z�,<��(<O%< F!<f�<�<�&<�{<��<�6<Ν<<�~ <
��;���;k�;�1�;tg�;��;�;ts�;���;B��;q0�;��;@Ū;˱�;��;Ҙ;��;[S�;4��;[7�;Y�y;H�n;ɍd;`PZ;�AP;�cF; �<;w43;-�);ڻ ;��;��;�N;��:���:���:���:���:r3�:��:�:&&|:�^:�.B:��%:�	:�>�9ٌ�9�_9�[�8@�&7a����E�4��2	ɹ�h��c���s/�	H��q`�v�x�7d���\���G���"��ﷺ��úCfϺ�ۺ��iI�������;n
��'������C!���&�?�,��C2�	�7�4�=��0C���H��tN�T��Y��W_���d�K�j�Q<p� �u��{������a��03��,���Ջ����y��bK��^��A��  �  �=V-=i�=Lw==��=�d=�=�� =\P =���<�-�<�s�<.��<��<yB�<G��<z��<�<�M�<��<'��<v�<�L�<*��<c��<��<};�<-t�<���<���<��<J�<�{�<T��<��<�<Z3�<�\�<��<��<���<���<�	�<�$�<�<�<�Q�<ec�<�q�<�|�<��<���<H��<Ђ�<;z�<8m�<�[�<~E�<e*�<S
�<��<X��<F��<sT�<��<V��<ُ�<?B�<���<���<�4�<���<}b�<O��<"x�<��<Ov�<��<�]�<rɺ<�/�<א�<��<&D�<���<��<.�<Qs�<n��<��<D+�<Ba�<瓤<�â<�<��<=A�<f�<���<;��<�Ǖ<��<���<��<�0�<bG�<�\�<�p�<���<���<概<?��<7�}<߬y<��u<�q<:n<I"j<�?f<E]b<�{^<��Z<��V<��R<_�N<)"K<�GG<oC<]�?<��;<��7<;"4<�U0<�,<�(<�%<{E!<��<c�<2&<6{<��<d6<E�<Y
<u~ <]��;w��;��;�1�;<g�;~��;��;�s�;���;��;�1�;��;�ƪ;3��;[��;bӘ;��;�T�;��;i8�;��y;��n;1�d;PZ;BP;�cF;D�<;�33;��);ʹ ;H�;��;ZK;���:���:З�:���:���:�/�:��:�݌:h |:��^:�+B:��%:w�	:9<�9��9�_9�~�8��(7�.��֧E������ȹ�Q��x��ih/�n�G�zg`��x��_���[��E��a ���ﷺʰú�gϺ�ۺ�溚L�u������,p
�E+�t����iF!�q�&��,�}E2���7� �=�N2C�6�H�yuN�T��Y��W_��d���j��:p���u��}{������`���1�����5ԋ�å���w��;J��W��=��  �  +�=j-=n�=Tw==v�=�d=�=�� =5P =;��<�-�<ls�<ո�<���<$B�<��<-��<��<�M�<Î�<���<b�<�L�<.��<n��<��<�;�<mt�<��<��<��<\J�<U|�<���<n��<��<�3�<�\�<(��<B��< ��<,��<�	�<�$�<�<�<�Q�<Wc�<�q�<�|�<��<O��<���<}��<�y�<�l�<U[�<.E�<*�<
�<���<6��<��<HT�<��<D��<��<QB�<���<��<5�<��<�b�<���<zx�<���<�v�<;�<E^�<�ɺ<0�<��<P�<oD�<ޖ�<��<.�<`s�<\��<��<+�<a�<���<2â<��<��<�@�<�e�<\��<娗<oǕ<4�<0��<��<�0�<BG�<�\�<�p�<���<���<��<r��<Ɏ}<R�y<H�u<��q<�n<#j<D@f<
^b<B|^<W�Z<K�V<Y�R<��N<�"K<"HG<3oC<~�?<��;<��7<"4<-U0<Ƌ,<p�(<$%<�D!<�<��<V%<�z<�<�5<~�<�	< ~ <f��;��;�;�1�;Qg�;���;-�;�t�;���;;�2�;�;�Ǫ;���;���;�Ԙ;��;�U�;���;Z9�;��y;"�n;�d;CPZ;�BP;�bF;��<;@23;��);ϸ ;b�;��;�H;M��:���:���:F�:N��:+�:��:zی:�|:��^:*B:�%:��	:B?�9���9�._9��8��*7X컸~E������ȹ�;��A��K\/���G��\`�ßx��Z��cW���B��2��ﷺ0�úiϺ�ۺ���O��������r
�!.����!��2I!�&�&���,�H2��7���=��3C�0�H�/vN�T�T�Y�9W_���d��j�>8p��u�Z{{�U���Z_��*0������ҋ�p���iv��I��p��$��  �  H�=w-=|�=Xw=�=p�=�d=�=�� =P =���<=-�<s�<u��<Z��<�A�<���<���<p�<]M�<z��<���<=�<�L�<��<���<��<�;�<�t�<��<j��<M�<�J�<�|�<
��<���<��<4�<I]�<���<p��<+��<c��<�	�<�$�<�<�<�Q�<Cc�<�q�<V|�<���<��<���<1��<�y�<�l�<�Z�<�D�<�)�<�	�<x��<��<׉�<"T�<��<<��<��<lB�<���<&��<F5�<1��<-c�<���<�x�<���<w�<��<�^�<!ʺ<m0�<��<r�<�D�<	��<��<8.�<Us�<W��<��<�*�<�`�<~��<�¢<��<N�<�@�<be�<���<���<!Ǖ<��<���<w�<h0�<G�<x\�<�p�<���<ו�<!��<���<�}<ԭy<�u<d�q<�n<�#j<Af<�^b<�|^<��Z<�V<��R<0�N<
#K<[HG<loC<��?<��;<k�7<�!4<�T0<6�,<��(<�%<.D!<1�<��<�$<�y<l�<5<�<W	<�} <���;c��;=�;o1�;g�;ݮ�;��;Gu�;:��;$��;�3�;-�;-ɪ;ߵ�;'��;֘;G
�;�V�;o��;:�;ءy;� o;f�d;�PZ;
BP;obF;��<;�03;��);_� ;D�;��;5F;���:��:��:�x�:H��:�%�:�ޛ:�֌:�|:V�^:�&B:q�%:v�	:�D�9���9�G_9���8#A,7����XE�����>�ȹb#������Q/�s�G�`S`���x�QY��
T���@��$����F�ú�iϺ�ۺ��溏S�q���ҵ�)u
��0�<���� L!���&��,��J2��7�I�=��5C���H��vN��T�U�Y�_V_�0�d�U�j�%7p��u�vx{�����]���.������Nы� ���.u���G��H����  �  \�=�-=��=Tw=�=h�=�d=�=b� =�O =���<�,�<�r�<��<��<aA�<H��<���<.�<M�<C��<���<�<�L�<��<��<��<�;�<�t�<Z��<���<��<K�<}�<d��<0��<"	�<r4�<�]�<΄�<���<]��<���<
�<�$�<�<�<�Q�<c�<aq�<?|�<Y��<܆�<W��<ށ�<-y�<&l�<�Z�<sD�<t)�<g	�<I��<���<���<T�<��<L��<ݏ�<�B�<���<I��<{5�<|��<{c�<;��<My�<3��<|w�<�<�^�<�ʺ<�0�<Ց�<��<�D�<(��<��<C.�<Ps�<a��<a�<�*�<�`�<:��<�¢</�<��<0@�<e�<���<3��<�ƕ<��<���<3�<U0�<�F�<\\�<�p�<���<땄<2��<з�<z�}<w�y<�u<��q<kn<a$j<�Af<`_b<�}^<��Z<}�V<��R<��N<]#K<HG<�oC<��?<��;<J�7<V!4<�T0<��,<v�(<�%<~C!<��< �<�#<�x<��<Z4<W�<�<
} <"��;���;�;91�;dg�;��;��;�u�;��;M��;�4�;���;�ʪ;0��;���;=ט;��;�W�;o��;;�;L�y;�o;�d;eQZ;�AP;�bF;u�<;�/3;��);� ;��;*�;�C;:��:��:/��:<s�:��:a �:�ۛ:�Ҍ:�|:Z�^:� B:��%:�	:�H�9Z��9�V_92!�8Ol.7�C���;E��ڕ���ȹ��,��-G/�R�G�LL`�Ҋx�mU��IQ��?�����h��úoiϺ�ۺѻ溒V���������w
�63�	�����O!���&���,�M2���7�i�=�x6C���H�uwN��T���Y��U_���d�%�j�y5p�{�u��v{����D\���-��g���Ћ�u���t���F������  �  m�=�-=��=Xw=�=\�=�d=�=N� =�O =e��<�,�<|r�<׷�<���<$A�< ��<C��<�
�<�L�<��<}��<��<�L�<��<���<��<<�<�t�<���<���<��<QK�<@}�<���<s��<k	�<�4�<�]�<��<��<���<���<5
�<�$�<�<�<Q�< c�<@q�<|�<-��<���<��<���<�x�<�k�<[Z�<8D�<7)�<+	�<��<���<���<�S�<v�<<��<��<�B�<&��<r��<�5�<���<�c�<���<�y�<~��<�w�<K�<>_�<�ʺ<�0�<	��<��<E�<Y��<�<V.�<Ts�<O��<K�<�*�<�`�<��<v¢<��<��<�?�<�d�<b��<�<�ƕ<Y�<���<
�<$0�<�F�<C\�<�p�<���<��<`��<���<�}<ͮy<��u<��q<�n<�$j<]Bf<�_b<E~^<)�Z<��V<��R< O<�#K<�HG<�oC<��?<��;<�7<%!4<1T0<\�,<	�(<n%<�B!<�<��<P#<kx<'�<�3<˚<Q<�| <Z��;��;��;&1�;�g�;���;w	�;av�;��;ዽ;�5�;���;[˪;/��;���;Pؘ;��;�X�;5��;�;�;��y;�o;9�d;�QZ;�AP;bF;��<;�.3;^�);�� ;��;3�;�A;g��:���:���:jo�:��:x�:Vכ:�ό:&|:��^:�B:M�%:H�	:M�9���9�h_9�L�8�J07���;E��˕�<�ȹ�����w��?/�1�G��C`��x�\Q���N��J<��M���췺�ú�jϺ�ۺ���;Y����ǹ��y
�^5������Q!���&�˧,��N2���7���=��7C���H�;xN�T�s�Y�U_�4�d��j��3p�$�u��t{�Ԋ��N[��z,��`����΋�}����r���E��d���홻�  �  v�=�-=��=_w=�=X�=�d=w=?� =�O =1��<u,�<7r�<���<s��<�@�<���<��<�
�<�L�<���<]��<��<~L�<��<���<��<<�<u�<���<
��<�<yK�<�}�<��<���<�	�<�4�<^�<0��<��<���<���<2
�<�$�<�<�<iQ�<
c�<8q�<�{�<��<b��<��<b��<�x�<�k�< Z�<�C�<�(�<	�<���<g��<b��<�S�<��<&��<��<�B�<!��<���<�5�<���<�c�<���<�y�<���<x�<��<�_�<˺<=1�<2��<"�<&E�<q��<�<Y.�<^s�<?��<Y�<�*�<d`�<璤<@¢<��<|�<�?�<}d�<&��<���<Uƕ<(�<F��<��<�/�<�F�<A\�<�p�<Ń�<���<j��<��<,�}<�y<b�u<��q<Bn<�%j<�Bf<�`b<�~^<��Z<t�V<:�R<f O<�#K<�HG<�oC<��?<��;<	�7<2!4<�S0<�,<��(<%<�B!<e�<�<�"<�w<��<t3<X�<�<b| <���;-��;X�;1�;�g�;]��;�	�;�v�;t��;k��;�6�;*��;`̪;G��;X��;�٘;I�;�Y�;ᾇ;b<�;��y;o;�d;�QZ;�AP;QaF;�<;7.3;��);�� ;��;��;�?;���:���:�}�:�j�:͟�:��:�ӛ:�͌:�|:��^:vB:P�%:��	:VK�9߱�9�r_9�k�8z617庸��D�iÕ���ȹg���o�6/�}�G��;`�u�x�aO��fM��;������췺��úlϺ�ۺF�溔[�s������"{
�_7���)���R!� '�p�,�~P2�k�7���=�_9C���H�IxN��T��Y�8U_���d�w�j��2p���u��r{�
����Z��7+��y����͋�����!r���D�����M홻�  �  ��=�-=��=bw=�=K�=xd=p=2� =�O =��<T,�<r�<|��<_��<�@�<���<���<�
�<�L�<��<K��<��<kL�<��<���<��<3<�<%u�<Ԭ�<'��<�<�K�<�}�<	��<���<�	�<�4�<-^�<E��<1��<���<���<I
�<�$�<�<�<`Q�<�b�<q�<�{�<���<O��<҅�<A��<�x�<�k�<	Z�<�C�<�(�<��<���<L��<U��<�S�<_�< ��<���<�B�<9��<���<�5�<��<�c�<���<�y�<���<#x�<��<�_�<$˺<Z1�<M��<A�<EE�<���<+�<g.�<`s�<3��<2�<�*�<S`�<В�<+¢<��<^�<�?�<ld�<��<���<5ƕ<�<2��<��<�/�<�F�<$\�<zp�<˃�<��<{��<"��<[�}<W�y<��u<(�q<�n<�%j<	Cf<�`b<�~^<ŝZ<��V<u�R<� O<$K< IG<�oC<��?<��;<��7<� 4<�S0<�,<o�(<� %<NB!<-�<��<�"<�w<b�<,3<!�<�<3| <y��;y��;�;�0�;�g�;���;�	�;
w�;���;׌�;�6�;���;�̪;���;���;�٘;��;NZ�;+��;�<�;]�y;o;��d;-RZ;BP;�`F;¯<;-3;w�);Ӱ ;�;��;u>;��:Z��:0|�:2i�:���:��:Nқ:�ˌ:��{:��^:�B::�%:�	:�O�9&��9_9��8�527Ӻ��D�F����ȹ����.l��2/���G�18`�c}x��M���K���9������뷺��ú�lϺwۺ����\�����<��2|
�T8��������S!�� '�q�,�_Q2�
�7�s�=��9C���H�)yN��T�׵Y��T_�Y�d���j��1p���u�@r{�����Z���*�����b͋�4����q��yD��S���왻�  �  ݊=d0=��=�z=�=��=Qi=�=ұ =�U =$��<N:�<��<|��<z�<S�<8��<���<� �<Td�<��<
��<!*�<nj�<���<���<�$�<�`�<B��<���<��<�C�<�x�<��<G��<�<3?�<�l�<���<\��<���<v�<�/�<�O�<�l�<��<'��<���<���<���<���<���<t��<6��<���<���<���<���<���<�r�<cO�<�&�<I��<"��<��<�I�<M�<���<�c�<

�< ��<�C�<B��<\d�<I��<l�<��<�[�<�ʼ<�4�<���<Q��<�P�<c��<��<�?�<N��<Qȭ<Q�<@�<?v�<ɨ�<ؤ<6�<h-�<�S�<�w�<���<��<�֗<9�<�<b$�<;�<YP�<>d�<�v�<t��<Ę�<C��<Ͷ�<�Ā<��}<�y<Y�u<_�q<�n<cj<4f<Lb<�d^<�}Z< �V<8�R<��N<u�J<�G<�-C<wP?<�u;<�7<��3<a�/<#,<{V(<u�$<�� <E<�L<$�<.�<�9<��
<��<�]<A��;X��;'�;"��;���;S��;��;�]�;v��;�8�;�Ļ;yf�;��;O�;�Ӣ;BҜ;B�;�;�b�;BŅ;yA�;�u;^k;`;`V;�TL;�{B;�8;YX/;5&;��;$;�A;r�;y~�:]��:��:���:~3�:Pפ:l��:��:��p:�S:JW7:�X:�a�9T��9ܒ9j;9�+�8�/��;���qd�0褹�(׹\{�p/���5��N��3f�F9~����i햺G���6���X;��K�ź��Ѻ�"ݺf���9������Y��M�I��z��MX���!�֡'�B-���2�z8�
>�R�C��BI�Y�N��nT�/Z���_�=4e���j�vdp���u�v�{������e���3��B��oϋ������l��Q<������ݙ��  �  ؊=k0=��=�z=�=��=Si=�=� =�U =5��<e:�<#��<���<��<2S�<A��<���<� �<ed�< ��<��<!*�<Hj�<���<���<�$�<�`�<8��<���<��<�C�<�x�<Ѭ�<1��<��<,?�<vl�<��<G��<���<p�<�/�<�O�<�l�<���<��<��<���<���<��<���<���<I��<���<��<���<���<���<�r�<iO�<�&�<[��<+��<���<�I�<\�<���<�c�<
�<��<�C�<-��<Fd�<&��<�k�<��<�[�<�ʼ<e4�<���<B��<�P�<[��<
��<�?�<X��<Wȭ<*�<@�<Jv�<ߨ�<#ؤ<@�<�-�<�S�<
x�<���<8��<�֗<Q�<*�<i$�<!;�<hP�<Fd�<�v�<i��<֘�<J��<ٶ�<�Ā<��}<̼y<=�u<'�q<�n<Nj<�3f<�Kb<zd^<�}Z<�V<�R<��N<^�J<�G<�-C<�P?<�u;<��7<��3<|�/<K#,<�V(<��$<�� <\<�L<g�<`�<�9<ϔ
<��<�]<���;���;)�;���;���;���;�;7^�;R��;�8�;�Ļ;Cf�;�;�;ZӢ;�ќ;*�;�;Lb�;�ą;8A�;ǭu;Hk;�`;^`V;UL;�zB;��8;�X/;�&;��;S;}B;�;��:���:0��:��:�4�:�ؤ:ؾ�:��:�p:2�S:�U7:U:�e�9'��9�ݒ96;9�'�8cx���N���|d����*׹�~�m2�D�5��N��5f��:~�����햺����򂮺�:����ź݊Ѻ"#ݺ���q8��=�����QL����Ь�/W���!�p�'�IA-���2��y8�	>�ݪC�FBI�'�N�<oT��Z�i�_��3e���j��dp��u��{����Tf���3������ϋ����m���<������ݙ��  �  Ǌ=\0=��=�z=�=��=gi=�=� =�U =^��<�:�<R��<���<��<YS�<q��<��<!�<�d�<4��<%��<K*�<\j�<���<���<�$�<|`�<��<���<��<fC�<�x�<���<��<��<?�<El�<Ǘ�<)��<c��<W�<�/�<�O�<�l�< ��<��<��<���<���<1��<���<���<x��<���<*��<ѽ�<ϩ�<��<�r�<�O�<�&�<f��<D��<��<�I�<b�<���<jc�<�	�<���<�C�<	��<&d�<���<�k�<��<�[�<�ʼ<:4�<h��<��<�P�<;��<���<�?�<E��<dȭ<;�<>@�<[v�<�<Aؤ<^�<�-�<(T�<2x�<љ�<]��<�֗<��<U�<�$�<>;�<pP�<ld�<�v�<x��<Ԙ�<)��<���<�Ā<\�}<��y<�u<��q<cn<�j<�3f<�Kb<d^<o}Z<��V<ϲR<\�N<�J<�G<v-C<�P?<�u;<�7<��3<��/<}#,<�V(<�$<:� <�<:M<��<��<X:<;�
<*�<�]<��;ӄ�;��;��;��;c��;��;�]�;���;88�;Ļ;�e�;z�;o�;�Ң;Iќ;��;N�;�a�;�ą;�@�;�u;Rk;c�`;�_V;AUL;�{B;��8;�Y/;&;��;8;�C;��;E��:���:"��:���:�7�:�ۤ:���:��:��p:��S:�Z7:'W:�g�9���9�ג9~;9��8����o����d������4׹a���6�~�5��N�J9f�H?~���������܄���;����ź��Ѻ� ݺv��27��C���	���J�������NV���!��'��?-���2��x8�'>���C�AI�G�N��nT��Z�n�_��4e��j��ep�,�u�Ø{�����g��l4��S��MЋ�̞���m���<��c��Wޙ��  �  ��=P0=��=�z=�=��=hi=�=� =V =���<�:�<���<��<�<�S�<���<W��<_!�<�d�<e��<E��<G*�<mj�<���<���<�$�<]`�<���<M��<X�<C�<ux�<P��<���<��<�>�<
l�<x��<���<(��<$�<�/�<�O�<�l�<��<+��<��<���<���<d��<+��<���<���<M��<���</��<��<��<s�<�O�<'�<���<X��<��<�I�<N�<���<ac�<�	�<ɩ�<mC�<���<�c�<���<fk�<A�<*[�<Sʼ<�3�<��<���<uP�<��<���<�?�<9��<Pȭ<J�<3@�<tv�<"��<~ؤ<��<�-�<rT�<�x�<3��<���<'ח<��<��<�$�<l;�<�P�<rd�<w�<|��<˘�<7��<���<fĀ<�}<�y<z�u<P�q<�n</j< 3f<�Jb<�c^<�|Z<�V<X�R<��N<��J<TG<�-C<vP?<�u;<�7<��3<��/<�#,<hW(<p�$<�� <b	<�M<n�<_�<�:<��
<��<�^<��;h��;��;E��;���;Z��;��;f]�;s��;l7�;9û;�d�;��;)�;�Ѣ;(М;��;r�;�`�;�Å;�?�;��u;}
k;6�`;�_V;�TL;|B;��8;EZ/;�&;��;�;�E;��;j��:;�:��:���:�;�:Dߤ:�ŕ:��:�p:��S:�Z7:WY:�c�9[��9�֒9��:9�ݢ8G�X�����d��	��ZN׹��qA�8�5��N��Cf�G~������¢�~���<����źv�Ѻ� ݺ����3��H�������H�)����7S� �!�y�'��=-���2��v8��>�T�C��@I��N��nT�Z�	�_�J5e���j�>gp�v��{�����'h��6��q���ы������n��>��K��4ߙ��  �  ��=40=��=�z= =��=i=�= � =(V =���<1;�<��<j��<~�<�S�<��<���<�!�<�d�<���<���<p*�<�j�<���<���<|$�<*`�<͚�<��<"�<�B�<x�<���<U��<3�<?>�<�k�<��<���<���<��</�<gO�<�l�<���<<��<5��<���< ��<���<p��<D��<��<���<���<���<r��<���<js�<P�<3'�<���<���<9��<�I�<J�<s��<*c�<�	�<���<*C�<���<_c�<\��<k�<��<�Z�<�ɼ<�3�<���<���</P�<ޤ�<���<�?�<)��<Qȭ<a�<W@�<�v�<U��<�ؤ<��<;.�<�T�<�x�<���<��<�ח<�<��<%�<�;�<�P�<�d�<-w�<���<Ę�<��<u��<:Ā<z�}<��y<��u<|�q<.n<qj<O2f<Jb<�b^<|Z<i�V<�R<k�N<��J<�G<M-C<eP?<�u;<N�7<[�3<~�/<J$,<�W(<�$<u� <'
<�N<?�<�<�;<l�
<n�<�^<��;���;���;��;��;J��;j�;�\�;޿�;�6�;|»;Rc�;*�;��;Т;�Μ;��;G�;!_�;�;?�;$�u;.	k;��`;W_V;�TL;�|B;�8;\/;�&;�;
;�H;��;-��:c�:?��:2��:"B�:��:{ʕ:��: �p:��S:_7:
\:d�9���9*ʒ9�:9-��8<۸�����-�d���:e׹d��?M��5�w#N�6Pf��M~��������Ţ�܆���<��l�ź��ѺiݺH��v0��N���-��JF�'��n��(P�>�!���'��:-���2��t8�>��C�^?I���N�:nT�DZ���_�	7e�I�j�ip��v�Y�{�Y���si��y7�����DӋ�O���Lp��l?��!��,����  �  ��=*0=��=�z= =��=�i==K� =WV =W��<�;�<v��<���<��<T�<���<��<"�<ae�<��<���<�*�<�j�<���<���<_$�<`�<���<���<��<dB�<�w�<���<���<��<�=�<@k�<���<E��<���<��<O/�<QO�<�l�<���<7��<_��<��<N��<���<���<���<���<��<W��< ��<��<���<�s�<mP�<�'�<��<���<e��<�I�<O�<a��<
c�<^	�<I��<�B�<��<c�<���<�j�<R�<;Z�<}ɼ<!3�<L��<,��<�O�<���<`��<�?�<��<Vȭ<[�<�@�<�v�<���<٤<L�<�.�<GU�<Oy�<��<���<�ח<��<P�<o%�<�;�<Q�<�d�<Iw�<���<̘�<��<a��<Ā<�}<ͺy<�u<��q<@n<�j<51f<(Ib<�a^<W{Z<��V<�R<��N<�J<�G<-C<hP?<�u;<s�7<��3<��/<�$,<�X(<�$<L� <<�O<,�<�<�<<Q�
<<�<�_<)��;=��;���;��;J��;W��;�;X\�;���;U5�;���;)b�;��;<�;D΢;�̜;��;x�;�]�;+��;�=�;+�u;�k;�`;�^V;oUL;�|B;v�8;L]/;o&;Q�;�;�K;D�;Ɣ�:��:���:���:�I�:��:�ϕ:j�:��p:��S:7e7:�[:�f�9���9�Ò9y�:9�k�8;^��+M���e�-=��ۀ׹��T]���5�&1N� Zf��Z~���������Ǣ�����'=����ź��Ѻ.ݺ��>,�����N���B�V��q���L�Q�!��'��7-���2��q8�;>�ʥC�>I��N�>nT�Z���_��7e��j�Kkp�
v�U�{�����Lk��M9����� Ջ�#����q���@�����Xᙻ�  �  [�=0=��=�z=	 =��=�i=$=y� =�V =���<<�<��<k��<l�<�T�<��<���<p"�<�e�<A��<���<�*�<�j�<���<r��<@$�<�_�<7��<��<Y�<�A�</w�<��<i��<5�<]=�<�j�<O��<տ�<H��<e�</�<7O�<ul�<��<C��<���<C��<���<Q��<!��<��<���<���<���<{��<e��<Z��<At�<�P�<�'�<H��<���<���<�I�<F�<1��<�b�<	�<���<B�<���<�b�<S��<j�<��<�Y�<�ȼ<�2�<ٖ�<���<�O�<6��<��<Y?�<�<Rȭ<j�<�@�<�v�<䩦<_٤<��</�<�U�<�y�<���<��<nؗ<��<��<�%�<Z<�<KQ�<e�<hw�<���<���<ৄ<B��<�À<m�}<8�y<B�u<��q<9n<�j<?0f<MHb<�`^<_zZ<ДV<h�R<T�N<]�J<bG<�,C<DP?<�u;<��7<%�3<.�/<�%,<QY(<��$<0� <<�P<1�<#�<�=<B�
<�<�`<���;#��;y��;���;z��;��;��;�[�;ɽ�;�4�;���;�`�;��;X�;�̢;˜;R�;��;X\�;���;�<�;�u;�k;f�`;�]V;eUL;*}B;��8;�^/;�&;;�;�;�O;��;���:��:���:���:+P�:��:֕:.��:�p:9�S:j7:y]:f�9��9���9"�:9��8�G��8���Ee��\����׹���k���5�"AN�&gf��g~� �����]ˢ�����:?����źN�Ѻ+ݺl���&��s���F��k?����~���H�K�!�6�'�&4-�d�2��n8�Z	>��C�f<I��N��mT�pZ�џ_��8e���j�Kmp�]v���{�����Tm���:������֋�+����s���B����G♻�  �  ?�=�/=��=�z= =�=�i=O=�� =�V =*��<�<�<k��<���<��<jU�<���< ��<�"�<�e�<���</��<�*�<�j�<���<f��< $�<�_�<���<#��<�
�<�A�<�v�<���<���<��<�<�<Tj�<ݕ�<t��<���<�<�.�<	O�<al�<��<g��<���<���<���<���<���<���<n��<��<C��<��<٫�<ג�<�t�<6Q�<#(�<���<��<���<J�<A�<��<�b�<��<���<B�<5��<b�<���<�i�<I�<8Y�<rȼ<#2�<a��<T��<)O�<룴<��</?�<݅�<Qȭ<��<�@�<@w�<%��<�٤<�<}/�<0V�<7z�<���<p��<�ؗ<s��<%�<(&�<�<�<�Q�<6e�<�w�<���<���<ʧ�<��<|À<��}<��y<{�u< �q<Y n<�j<?/f<IGb<�_^<{yZ< �V<��R<��N<��J<�
G<�,C<4P?<�u;<�7<u�3<��/<+&,< Z(<��$</� <<�Q<0�<�<�><8�
<��<$a<О�;���;��;O��;ť�;��;[�;[�;��;?3�;L��;_�;>�;��;�ʢ;2ɜ;p��;��;�Z�;��;L;�;��u;=k;�`;X]V;sUL;m~B;��8;�`/;V&;�;H;�R;��;a��:"�:��:P��:;X�:R��:�ܕ:���:�p:��S:�m7:�b:�f�9���9g��9��:93ҡ8a�������}e�bw��i�׹���={���5��NN��tf�Cs~��%��<��w΢������?���źɂѺ�ݺ��躊"��G���ц��;�������D���!�6�'�20-�
�2�l8��>�@�C��:I��N�*mT��Z���_�Y:e�B�j�pp�v�٦{�F���o���<���
���؋�즎�Vu�� D��v���㙻�  �  2�=�/=�=�z= =�=�i=m=�� =�V =���<�<�<ރ�<O��<q�<�U�<���<S��<?#�<if�<ɨ�<g��<	+�<�j�<���<h��< $�<}_�<ә�<���<�
�<&A�<Yv�<��<m��<C�<_<�<�i�<q��<��<���<��<�.�<�N�<cl�<��<o��<���<���<'��<���<���<���<���<{��<���<r��<D��<K��<�t�<�Q�<}(�<���<<��<���<J�<0�<��<b�<��<a��<�A�<���<�a�<_��<i�<��<�X�<�Ǽ<�1�<<���<�N�<���<��< ?�<څ�<@ȭ<��<�@�<nw�<d��< ڤ<r�<�/�<�V�<�z�<��<껙<`ٗ<���<y�<�&�<�<�<�Q�<Se�<�w�<���<���<ħ�<ܵ�<dÀ<!�}<��y<��u<%�q<i�m<�j<X.f<BFb<_^<�xZ<5�V<�R<��N<��J<�
G<x,C<+P?<�u;<�7<��3<T�/<�&,<�Z(<O�$<�� <�<�R<O�<��<�?<�
<��<b<��;���;���;ƌ�;ť�;'��;��;~Z�;w��;�1�;	��;�]�;��;��;�Ȣ;�ǜ;�ޖ;*�;Y�;ɼ�;�9�;ءu;tk;��`;�]V;4UL;�~B;��8;@b/;�&;�;{;SU;O�;U��:h&�:i��:>�:�_�:>��:�:��:��p:-�S:�p7:�c:�c�9���9���9�}:9���84P��St����e�q���[�׹��I���6�
\N�8�f��}~��+������Т�/����?����ź��Ѻ=ݺe��J��Ȗ�����^9���s���@��!���'�*--�o�2��h8�>�H�C�:I�:�N�mT��Z���_��;e��j�}rp�4v��{������p���>������ڋ����� w���E�����噻�  �  �=�/=l�=�z= =#�=�i=�=ܲ =�V =���<F=�<6��<���<��<;V�<N��<���<�#�<�f�< ��<���<@+�<�j�<���<Z��<�#�<I_�<���<���<d
�<�@�<�u�<���<��<��<<�<yi�<��<˾�<Z��<��<p.�<�N�<Hl�<���<x��<��<���<Q��<��<$��<6��<7��<���<!��<���<���<���<Yu�<�Q�<�(�<���<b��<ۊ�<J�<)�<���<Ub�<m�<��<xA�<���<Ia�<���<�h�<d�<OX�<�Ǽ<E1�<���<���<�N�<h��<x�<�>�<Å�<=ȭ<��<A�<�w�<���<5ڤ<��<30�<�V�<{�<Ԝ�<H��<�ٗ<7��<��<�&�<'=�<R�<�e�<�w�<���<���<���<���<À<��}<[�y<�u<s�q<��m<�j<�-f<�Eb<H^^<�wZ<��V<~�R<|�N<�J<2
G<,,C<P?<�u;<Z�7<�3<��/<G',<F[(<�$<�� <�<ES<�<��<^@<ƚ
<h�<b<���;O��;x��;?��;���;
��;��;�Y�;_��;11�;��;G\�;K�;��;�Ǣ;Ɯ;eݖ;��;�W�;���;9�;3�u;�k;��`;�\V;/UL;7B;�8;�c/;&;�;D;�X;:�;��:j,�:;��:��:@e�:��:��:��:C�p:y�S:�v7:5e:pc�9��9���9<`:9�]�8d	������w�e�N���)�׹:��F��&6�2hN��f�{�~��.��q	��CԢ�]����@����źu�Ѻ�ݺ�����F������
6��������=��!��'�*-�x�2�g8�>��C�a8I�(�N��lT�3Z�ۡ_�7=e���j�Ctp��v�a�{�Z���fr��I@��2��&܋�A���qx���F������噻�  �  ��=�/=e�=�z= =�=�i=�=�� =W =&��<�=�<���<
��<�<�V�<���<	��<�#�<�f�<6��<���<O+�<�j�<���<T��<�#�<B_�<]��<d��<
�<�@�<�u�<j��<���<�<�;�</i�<��<}��<��<d�<U.�<�N�<4l�<���<~��<߲�<���<x��<U��<b��<���<l��<2��<r��<��< ��<Փ�<�u�<R�<�(�<'��<���<ۊ�<J�<6�<��<Tb�<P�<��<<A�<.��<a�<���<Ph�<��<�W�<7Ǽ<�0�<O��<R��<NN�<5��<f�<�>�<���<Eȭ<��<A�<�w�<Ū�<mڤ<��<0�<.W�<j{�<��<���<	ڗ<v��<&�<'�<`=�<,R�<�e�<�w�<ǈ�<���<���<���<�<N�}<ͷy<��u<�q<
�m<Vj<�,f<�Db<�]^<qwZ<�V<�R<�N<��J<-
G<,C<P?<v;<C�7<F�3<��/<�',<�[(<��$<H� <R<T<��<��<�@<h�
<��< c<��;΋�;Ȅ�;+��;9��;	��;��;�Y�;κ�;�0�;ﺻ;l[�;j�;F�;SƢ;�Ĝ;+ܖ;��;W�;v��;78�;��u;� k;Ε`;Q\V;�UL;xB;�8;�d/;O&;�;E;D[;��;��:�1�:+��:P�:�h�:
�:��:!
�:�p:��S:w7:�e:�g�9N��9k��9T:9�)�8|濷&��;�e�龥��عG��Z��d!6�.pN�v�f���~�2��I��բ�����uA����ź܀Ѻ�ݺØ躾���������3����J���;�7�!�M�'�(-��2�6e8�B>��C�u7I�{�N��lT��Z�R�_� =e���j��up�v���{�6����s���A�����f݋�����Ty��H������晻�  �  �=�/=[�=�z= =-�=j=�=� =-W =@��<�=�<���<2��<7�<�V�<�<'��<�#�<�f�<O��<���<k+�<k�<���<E��<�#�<_�<T��<F��<�	�<g@�<�u�<@��<���<b�<�;�< i�<���<^��<���<Q�<?.�<�N�<"l�<��<���<���<��<���<w��<���<���<���<[��<���<;��<'��<���<�u�<)R�<)�<?��<���<��<0J�<)�<ҵ�<*b�<3�<ӧ�<A�<��<�`�<y��<#h�<��<�W�<Ǽ<�0�<��<3��<-N�<(��<A�<�>�<���<@ȭ<��<$A�<�w�<۪�<�ڤ<�<�0�<^W�<�{�<C��<ȼ�<3ڗ<���<@�<&'�<|=�<MR�<�e�<�w�<҈�<���<~��<���<�<$�}<��y<=�u<��q<��m<j<�,f<�Db<E]^<wZ<��V<��R<��N<��J<�	G<�+C<�O?<v;<��7<��3<'�/<�',<\(<ԓ$<�� <�<XT<�<��<QA<��
<3�<Kc<V��;g��;D��;���;I��;���;�;:Y�;���;$0�;���;�Z�;��;�ߨ;�Ţ;9Ĝ;�ۖ;��;FV�;��;�7�; �u;% k;��`;�[V;[UL;�B;�8;�e/;5&;�;a;#\;>�;���:�3�:l��:��:fk�:��:��:b�:H�p:��S:Iz7:�h:�d�9/��9z��9?G:9Q�8�c���-��f��ʥ��ع��P���&6�;vN���f�&�~��3�����*ע�����iB����źѺ]ݺ���:��U����~��2�6����]:�
�!���'��&-�8�2�d8�_ >��C��6I���N�1lT�YZ���_�r>e���j�qvp��v�Ư{����bt��-B��*��ދ�=���&z���H��l���晻�  �  �=�/=l�=�z= =*�=j=�=� =5W =P��<�=�<ń�<C��<T�<�V�<ݛ�<B��<�#�<g�<W��<���<_+�<k�<���<U��<�#�<_�<E��<'��<�	�<R@�<su�<1��<v��<>�<~;�<�h�<���<U��<���<=�<5.�<�N�<Fl�<؆�<���<���<
��<���<���<���<���<���<f��<���<W��<0��<!��<�u�<:R�< )�<D��<���<��<%J�<�<��<2b�<*�<���<�@�<��<�`�<g��<h�<��<�W�<�Ƽ<�0�<	��<,��<N�<��<6�<�>�<���<-ȭ<��<A�<�w�<⪦<�ڤ< �<�0�<|W�<�{�<`��<ܼ�<Fڗ<���<O�<2'�<�=�<YR�<�e�<�w�<ň�<���<���<���<�<�}<p�y<$�u<n�q<��m<�j<J,f<fDb</]^<�vZ<��V<��R<��N<��J<�	G<&,C<�O?<�u;<v�7<h�3<?�/<	(,<#\(<��$<�� <�<{T<)�<��<�A<�
<T�<gc<{��;���;��;���;��;��;v�;Y�;��;�/�;v��;yZ�;[�;sߨ;HŢ;�Ü;?ۖ;��;�U�;久;i7�;��u;��j;Ô`;�\V;UL;�B;��8;�e/;w&;p;�;�\;Y�;t��:o5�:0��:v�:�m�:�:�:}�:��p:s�S:uy7:Bg:{a�90��9疒9C:9��8H����5���f�ϥ�!عO��ȩ��(6��xN���f��~��5������ע�����A����ź�Ѻݺ=�����e���~��1�A��Ə�s9�l�!�e�'��%-���2��c8���=���C�7I���N��lT�aZ�ԡ_�p>e�[�j�^wp�rv�'�{�_����t���B�����}ދ�f����z���H�����t登�  �  �=�/=[�=�z= =-�=j=�=� =-W =@��<�=�<���<2��<7�<�V�<�<'��<�#�<�f�<O��<���<k+�<k�<���<E��<�#�<_�<T��<F��<�	�<g@�<�u�<@��<���<b�<�;�< i�<���<^��<���<Q�<?.�<�N�<"l�<��<���<���<��<���<w��<���<���<���<[��<���<;��<'��<���<�u�<)R�<)�<?��<���<��<0J�<)�<ҵ�<*b�<3�<ӧ�<A�<��<�`�<y��<#h�<��<�W�<Ǽ<�0�<��<3��<-N�<(��<A�<�>�<���<@ȭ<��<$A�<�w�<۪�<�ڤ<�<�0�<^W�<�{�<C��<ȼ�<3ڗ<���<@�<&'�<|=�<MR�<�e�<�w�<҈�<���<~��<���<�<$�}<��y<=�u<��q<��m<j<�,f<�Db<E]^<wZ<��V<��R<��N<��J<�	G<�+C<�O?<v;<��7<��3<'�/<�',<\(<ԓ$<�� <�<XT<�<��<QA<��
<3�<Kc<V��;g��;D��;���;I��;���;�;:Y�;���;$0�;���;�Z�;��;�ߨ;�Ţ;9Ĝ;�ۖ;��;FV�;��;�7�; �u;% k;��`;�[V;[UL;�B;�8;�e/;5&;�;a;#\;>�;���:�3�:l��:��:fk�:��:��:b�:H�p:��S:Iz7:�h:�d�9/��9z��9?G:9Q�8�c���-��f��ʥ��ع��P���&6�;vN���f�&�~��3�����*ע�����iB����źѺ]ݺ���:��U����~��2�6����]:�
�!���'��&-�8�2�d8�_ >��C��6I���N�1lT�YZ���_�r>e���j�qvp��v�Ư{����bt��-B��*��ދ�=���&z���H��l���晻�  �  ��=�/=e�=�z= =�=�i=�=�� =W =&��<�=�<���<
��<�<�V�<���<	��<�#�<�f�<6��<���<O+�<�j�<���<T��<�#�<B_�<]��<d��<
�<�@�<�u�<j��<���<�<�;�</i�<��<}��<��<d�<U.�<�N�<4l�<���<~��<߲�<���<x��<U��<b��<���<l��<2��<r��<��< ��<Փ�<�u�<R�<�(�<'��<���<ۊ�<J�<6�<��<Tb�<P�<��<<A�<.��<a�<���<Ph�<��<�W�<7Ǽ<�0�<O��<R��<NN�<5��<f�<�>�<���<Eȭ<��<A�<�w�<Ū�<mڤ<��<0�<.W�<j{�<��<���<	ڗ<v��<&�<'�<`=�<,R�<�e�<�w�<ǈ�<���<���<���<�<N�}<ͷy<��u<�q<
�m<Vj<�,f<�Db<�]^<qwZ<�V<�R<�N<��J<-
G<,C<P?<v;<C�7<F�3<��/<�',<�[(<��$<H� <R<T<��<��<�@<h�
<��< c<��;΋�;Ǆ�;+��;9��;	��;��;�Y�;κ�;�0�;ﺻ;l[�;j�;F�;SƢ;�Ĝ;+ܖ;��;W�;v��;78�;��u;� k;Ε`;Q\V;�UL;xB;�8;�d/;O&;�;E;D[;��;��:�1�:+��:P�:�h�:
�:��:!
�:�p:��S:w7:�e:�g�9N��9k��9T:9�)�8|濷&��;�e�龥��عG��Z��d!6�.pN�v�f���~�2��I��բ�����uA����ź܀Ѻ�ݺØ躾���������3����J���;�7�!�M�'�(-��2�6e8�B>��C�u7I�{�N��lT��Z�R�_� =e���j��up�v���{�6����s���A�����f݋�����Ty��H������晻�  �  �=�/=l�=�z= =#�=�i=�=ܲ =�V =���<F=�<6��<���<��<;V�<N��<���<�#�<�f�< ��<���<@+�<�j�<���<Z��<�#�<I_�<���<���<d
�<�@�<�u�<���<��<��<<�<yi�<��<˾�<Z��<��<p.�<�N�<Hl�<���<x��<��<���<Q��<��<$��<6��<7��<���<!��<���<���<���<Yu�<�Q�<�(�<���<b��<ۊ�<J�<)�<���<Ub�<m�<��<xA�<���<Ia�<���<�h�<d�<OX�<�Ǽ<E1�<���<���<�N�<h��<x�<�>�<Å�<=ȭ<��<A�<�w�<���<5ڤ<��<30�<�V�<{�<Ԝ�<H��<�ٗ<7��<��<�&�<'=�<R�<�e�<�w�<���<���<���<���<À<��}<[�y<�u<s�q<��m<�j<�-f<�Eb<H^^<�wZ<��V<~�R<|�N<�J<2
G<,,C<P?<�u;<Z�7<�3<��/<G',<F[(<�$<�� <�<ES<�<��<^@<ƚ
<h�<b<���;O��;x��;?��;���;
��;��;�Y�;_��;01�;��;G\�;K�;��;�Ǣ;Ɯ;eݖ;��;�W�;���;9�;3�u;�k;��`;�\V;/UL;7B;�8;�c/;&;�;D;�X;:�;��:j,�:;��:��:@e�:��:��:��:C�p:y�S:�v7:5e:pc�9��9���9<`:9�]�8d	������w�e�N���)�׹:��F��&6�2hN��f�{�~��.��q	��CԢ�]����@����źu�Ѻ�ݺ�����F������
6��������=��!��'�*-�x�2�g8�>��C�a8I�(�N��lT�3Z�ۡ_�7=e���j�Ctp��v�a�{�Z���fr��I@��2��&܋�A���qx���F������噻�  �  2�=�/=�=�z= =�=�i=m=�� =�V =���<�<�<ރ�<O��<q�<�U�<���<S��<?#�<if�<ɨ�<g��<	+�<�j�<���<h��< $�<}_�<ә�<���<�
�<&A�<Yv�<��<m��<C�<_<�<�i�<q��<��<���<��<�.�<�N�<cl�<��<o��<���<���<'��<���<���<���<���<{��<���<r��<D��<K��<�t�<�Q�<}(�<���<<��<���<J�<0�<��<b�<��<a��<�A�<���<�a�<_��<i�<��<�X�<�Ǽ<�1�<<���<�N�<���<��< ?�<څ�<@ȭ<��<�@�<nw�<d��< ڤ<r�<�/�<�V�<�z�<��<껙<`ٗ<���<y�<�&�<�<�<�Q�<Se�<�w�<���<���<ħ�<ܵ�<dÀ<!�}<��y<��u<%�q<i�m<�j<X.f<BFb<_^<�xZ<5�V<�R<��N<��J<�
G<x,C<+P?<�u;<�7<��3<T�/<�&,<�Z(<O�$<�� <�<�R<O�<��<�?<�
<��<b<��;���;���;Ō�;ť�;'��;��;~Z�;w��;�1�;	��;�]�;��;��;�Ȣ;�ǜ;�ޖ;*�;Y�;ɼ�;�9�;ءu;tk;��`;�]V;4UL;�~B;��8;@b/;�&;�;{;SU;O�;U��:h&�:i��:>�:�_�:>��:�:��:��p:-�S:�p7:�c:�c�9���9���9�}:9���84P��St����e�q���[�׹��I���6�
\N�8�f��}~��+������Т�/����?����ź��Ѻ=ݺe��J��Ȗ�����^9���s���@��!���'�*--�o�2��h8�>�H�C�:I�:�N�mT��Z���_��;e��j�}rp�4v��{������p���>������ڋ����� w���E�����噻�  �  ?�=�/=��=�z= =�=�i=O=�� =�V =*��<�<�<k��<���<��<jU�<���< ��<�"�<�e�<���</��<�*�<�j�<���<f��< $�<�_�<���<#��<�
�<�A�<�v�<���<���<��<�<�<Tj�<ݕ�<t��<���<�<�.�<	O�<al�<��<g��<���<���<���<���<���<���<n��<��<C��<��<٫�<ג�<�t�<6Q�<#(�<���<��<���<J�<A�<��<�b�<��<���<B�<5��<b�<���<�i�<I�<8Y�<rȼ<#2�<a��<T��<)O�<룴<��</?�<ޅ�<Qȭ<��<�@�<@w�<%��<�٤<�<}/�<0V�<7z�<���<p��<�ؗ<s��<%�<(&�<�<�<�Q�<6e�<�w�<���<���<ʧ�<��<|À<��}<��y<{�u< �q<Y n<�j<?/f<IGb<�_^<{yZ< �V<��R<��N<��J<�
G<�,C<4P?<�u;<�7<u�3<��/<+&,< Z(<��$</� <<�Q<0�<�<�><8�
<��<$a<О�;���;��;O��;ť�;��;[�;[�;��;?3�;L��;_�;>�;��;�ʢ;2ɜ;p��;��;�Z�;��;K;�;��u;=k;�`;X]V;sUL;m~B;��8;�`/;V&;�;H;�R;��;a��:"�:��:P��:;X�:R��:�ܕ:���:�p:��S:�m7:�b:�f�9���9g��9��:93ҡ8a�������}e�bw��i�׹���={���5��NN��tf�Cs~��%��<��w΢������?���źɂѺ�ݺ��躊"��G���ц��;�������D���!�6�'�20-�
�2�l8��>�@�C��:I��N�*mT��Z���_�Y:e�B�j�pp�v�٦{�F���o���<���
���؋�즎�Vu�� D��v���㙻�  �  [�=0=��=�z=	 =��=�i=$=y� =�V =���<<�<��<k��<l�<�T�<��<���<p"�<�e�<A��<���<�*�<�j�<���<r��<@$�<�_�<7��<��<Y�<�A�</w�<��<i��<5�<]=�<�j�<O��<տ�<H��<e�</�<7O�<ul�<��<C��<���<C��<���<Q��<!��<��<���<���<���<{��<e��<Z��<At�<�P�<�'�<H��<���<���<�I�<F�<1��<�b�<	�<���<B�<���<�b�<S��<j�<��<�Y�<�ȼ<�2�<ٖ�<���<�O�<6��<��<Y?�<�<Rȭ<j�<�@�<�v�<䩦<_٤<��</�<�U�<�y�<���<��<nؗ<��<��<�%�<Z<�<KQ�<e�<hw�<���<���<ৄ<B��<�À<m�}<8�y<B�u<��q<9n<�j<?0f<MHb<�`^<_zZ<ДV<h�R<T�N<]�J<cG<�,C<DP?<�u;<��7<%�3<.�/<�%,<QY(<��$<0� <<�P<1�<#�<�=<B�
<�<�`<���;#��;y��;���;z��;��;��;�[�;ɽ�;�4�;���;�`�;��;X�;�̢;˜;R�;��;X\�;���;�<�;�u;�k;f�`;�]V;eUL;*}B;��8;�^/;�&;;�;�;�O;��;���:��:���:���:+P�:��:֕:.��:�p:9�S:j7:y]:f�9��9���9"�:9��8�G��8���Ee��\����׹���k���5�"AN�&gf��g~� �����]ˢ�����:?����źN�Ѻ+ݺl���&��s���F��k?����~���H�K�!�6�'�&4-�d�2��n8�Z	>��C�f<I��N��mT�pZ�џ_��8e���j�Kmp�]v���{�����Tm���:������֋�+����s���B����G♻�  �  ��=*0=��=�z= =��=�i==K� =WV =W��<�;�<v��<���<��<T�<���<��<"�<ae�<��<���<�*�<�j�<���<���<_$�<`�<���<���<��<dB�<�w�<���<���<��<�=�<@k�<���<E��<���<��<O/�<QO�<�l�<���<7��<_��<��<N��<���<���<���<���<��<W��< ��<��<���<�s�<mP�<�'�<��<���<e��<�I�<O�<a��<
c�<^	�<I��<�B�<��<c�<���<�j�<R�<;Z�<}ɼ<!3�<L��<,��<�O�<���<`��<�?�<��<Vȭ<[�<�@�<�v�<���<٤<L�<�.�<GU�<Oy�<��<���<�ח<��<P�<o%�<�;�<Q�<�d�<Iw�<���<̘�<��<a��<Ā<�}<ͺy<�u<��q<@n<�j<51f<(Ib<�a^<W{Z<��V<�R<��N<�J<�G<-C<hP?<�u;<s�7<��3<��/<�$,<�X(<�$<L� <<�O<,�<�<�<<Q�
<<�<�_<(��;=��;���;��;I��;W��;�;X\�;���;T5�;���;)b�;��;<�;D΢;�̜;��;x�;�]�;+��;�=�;+�u;�k;�`;�^V;nUL;�|B;v�8;L]/;o&;Q�;�;�K;D�;Ɣ�:��:���:���:�I�:��:�ϕ:j�:��p:��S:7e7:�[:�f�9���9�Ò9y�:9�k�8;^��+M���e�-=��ۀ׹��T]���5�&1N� Zf��Z~���������Ǣ�����'=����ź��Ѻ.ݺ��>,�����N���B�V��q���L�Q�!��'��7-���2��q8�;>�ʥC�>I��N�>nT�Z���_��7e��j�Kkp�
v�U�{�����Lk��M9����� Ջ�#����q���@�����Xᙻ�  �  ��=40=��=�z= =��=i=�= � =(V =���<1;�<��<j��<~�<�S�<��<���<�!�<�d�<���<���<p*�<�j�<���<���<|$�<*`�<͚�<��<"�<�B�<x�<���<U��<3�<?>�<�k�<��<���<���<��</�<gO�<�l�<���<<��<5��<���< ��<���<p��<D��<��<���<���<���<r��<���<js�<P�<3'�<���<���<9��<�I�<J�<s��<*c�<�	�<���<*C�<���<_c�<\��<k�<��<�Z�<�ɼ<�3�<���<���</P�<ޤ�<���<�?�<)��<Qȭ<a�<W@�<�v�<U��<�ؤ<��<;.�<�T�<�x�<���<��<�ח<�<��<%�<�;�<�P�<�d�<-w�<���<Ę�<��<u��<:Ā<z�}<��y<��u<|�q<.n<qj<O2f<Jb<�b^<|Z<i�V<�R<k�N<��J<�G<M-C<eP?<�u;<N�7<[�3<~�/<J$,<�W(<�$<u� <'
<�N<?�<�<�;<l�
<n�<�^<��;���;���;��;��;I��;j�;�\�;޿�;�6�;{»;Rc�;*�;��;Т;�Μ;��;G�;!_�;�;?�;$�u;-	k;��`;V_V;�TL;�|B;�8;\/;�&;�;
;�H;��;-��:c�:?��:2��:"B�:��:{ʕ:��: �p:��S:_7:
\:d�9���9*ʒ9�:9-��8<۸�����-�d���:e׹d��?M��5�w#N�6Pf��M~��������Ţ�܆���<��l�ź��ѺiݺH��v0��N���-��JF�'��n��(P�>�!���'��:-���2��t8�>��C�^?I���N�:nT�DZ���_�	7e�I�j�ip��v�Y�{�Y���si��y7�����DӋ�O���Lp��l?��!��,����  �  ��=P0=��=�z=�=��=hi=�=� =V =���<�:�<���<��<�<�S�<���<W��<_!�<�d�<e��<E��<G*�<mj�<���<���<�$�<]`�<���<M��<X�<C�<ux�<P��<���<��<�>�<
l�<x��<���<(��<$�<�/�<�O�<�l�<��<+��<��<���<���<d��<+��<���<���<M��<���</��<��<��<s�<�O�<'�<���<X��<��<�I�<N�<���<ac�<�	�<ɩ�<mC�<���<�c�<���<fk�<A�<*[�<Sʼ<�3�<��<���<uP�<��<���<�?�<9��<Pȭ<J�<3@�<tv�<"��<~ؤ<��<�-�<rT�<�x�<3��<���<'ח<��<��<�$�<l;�<�P�<qd�<w�<|��<˘�<7��<���<fĀ<�}<�y<z�u<P�q<�n</j< 3f<�Jb<�c^<�|Z<�V<X�R<��N<��J<TG<�-C<vP?<�u;<�7<��3<��/<�#,<hW(<p�$<�� <b	<�M<n�<_�<�:<��
<��<�^<��;h��;��;E��;���;Z��;��;f]�;s��;l7�;9û;�d�;��;)�;�Ѣ;(М;��;r�;�`�;�Å;�?�;��u;}
k;6�`;�_V;�TL;|B;��8;EZ/;�&;��;�;�E;��;j��:;�:��:���:�;�:Dߤ:�ŕ:��:�p:��S:�Z7:WY:�c�9[��9�֒9��:9�ݢ8G�X�����d��	��ZN׹��qA�8�5��N��Cf�G~������¢�~���<����źv�Ѻ� ݺ����3��H�������H�)����7S� �!�y�'��=-���2��v8��>�T�C��@I��N��nT�Z�	�_�J5e���j�>gp�v��{�����'h��6��q���ы������n��>��K��4ߙ��  �  Ǌ=\0=��=�z=�=��=gi=�=� =�U =^��<�:�<R��<���<��<YS�<q��<��<!�<�d�<4��<%��<K*�<\j�<���<���<�$�<|`�<��<���<��<fC�<�x�<���<��<��<?�<El�<Ǘ�<)��<c��<W�<�/�<�O�<�l�< ��<��<��<���<���<1��<���<���<x��<���<*��<ѽ�<ϩ�<��<�r�<�O�<�&�<f��<D��<��<�I�<b�<���<jc�<�	�<���<�C�<	��<&d�<���<�k�<��<�[�<�ʼ<:4�<h��<��<�P�<;��<���<�?�<E��<dȭ<;�<>@�<[v�<�<Aؤ<^�<�-�<(T�<2x�<љ�<]��<�֗<��<U�<�$�<>;�<pP�<ld�<�v�<x��<Ԙ�<)��<���<�Ā<\�}<��y<�u<��q<cn<�j<�3f<�Kb<d^<o}Z<��V<ϲR<\�N<�J<�G<v-C<�P?<�u;<�7<��3<��/<}#,<�V(<�$<:� <�<:M<��<��<X:<;�
<*�<�]<��;҄�;��;��;��;c��;��;�]�;���;88�;Ļ;�e�;z�;o�;�Ң;Iќ;��;N�;�a�;�ą;�@�;�u;Rk;c�`;�_V;AUL;�{B;��8;�Y/;&;��;8;�C;��;E��:���:"��:���:�7�:�ۤ:���:��:��p:��S:�Z7:'W:�g�9���9�ג9~;9��8����o����d������4׹a���6�~�5��N�J9f�H?~���������܄���;����ź��Ѻ� ݺv��27��C���	���J�������NV���!��'��?-���2��x8�'>���C�AI�G�N��nT��Z�n�_��4e��j��ep�,�u�Ø{�����g��l4��S��MЋ�̞���m���<��c��Wޙ��  �  ؊=k0=��=�z=�=��=Si=�=� =�U =5��<e:�<#��<���<��<2S�<A��<���<� �<ed�< ��<��<!*�<Hj�<���<���<�$�<�`�<8��<���<��<�C�<�x�<Ѭ�<1��<��<,?�<vl�<��<G��<���<p�<�/�<�O�<�l�<���<��<��<���<���<��<���<���<I��<���<��<���<���<���<�r�<iO�<�&�<[��<+��<���<�I�<\�<���<�c�<
�<��<�C�<-��<Fd�<&��<�k�<��<�[�<�ʼ<e4�<���<B��<�P�<[��<
��<�?�<X��<Wȭ<*�<@�<Jv�<ߨ�<#ؤ<@�<�-�<�S�<
x�<���<8��<�֗<Q�<*�<i$�<!;�<hP�<Fd�<�v�<i��<֘�<J��<ٶ�<�Ā<��}<̼y<=�u<'�q<�n<Nj<�3f<�Kb<zd^<�}Z<�V<�R<��N<^�J<�G<�-C<�P?<�u;<��7<��3<|�/<K#,<�V(<��$<�� <\<�L<g�<`�<�9<ϔ
<��<�]<���;���;)�;���;���;���;�;7^�;R��;�8�;�Ļ;Cf�;�;�;ZӢ;�ќ;*�;�;Lb�;�ą;8A�;ǭu;Hk;�`;^`V;UL;�zB;��8;�X/;�&;��;S;}B;�;��:���:0��:��:�4�:�ؤ:ؾ�:��:�p:2�S:�U7:U:�e�9'��9�ݒ96;9�'�8cx���N���|d����*׹�~�m2�D�5��N��5f��:~�����햺����򂮺�:����ź݊Ѻ"#ݺ���q8��=�����QL����Ь�/W���!�p�'�IA-���2��y8�	>�ݪC�FBI�'�N�<oT��Z�i�_��3e���j��dp��u��{����Tf���3������ϋ����m���<������ݙ��  �  K�=;3=�=�~=$=N�=@n=
=�� =�[ =)  =~H�<D��<���<��<�e�<��<��<�7�<�|�<���<[�<G�<���<���<�	�<XH�<��<q��<���<�7�<-p�<���<h��<��<�D�<&v�<Υ�<���<W��<)�<hP�<bu�<���<S��<���<���<��<��<o&�<U2�<�:�<�>�<�>�<�:�<Y2�<Z%�<��<��<��<��<��<gl�<�9�<�<��<o|�<t0�<���<U��<F$�<���<BP�<d��<:b�<���<�Z�<ξ<V;�<ࢻ<��<a�<��<
�<�V�<���<9�<!�<�[�<H��<Ũ<1��< �<�H�<�n�<���<;��<�Л<��<5�<��<r6�<�K�<h_�<�q�<͂�<���< ��<���<1��<�Ƃ<�р<��}<�y<��u<n�q<$n<�j<�$f<�6b<`I^<�\Z<:qV<ÆR<<�N<7�J<Z�F<��B<F?<�$;<
F7<[i3<��/<��+<��'<�$<�J <��<K�<@<�L<h�<��	<�J<��<*�;S
�;K��;���;_�;d(�;�Z�;���;���;�e�;q�;ǀ�;R0�;Q��;�֠;�Ϛ;�;�;�R�;��;�[|;�q;��f;�v\;5?R;�8H;hf>;z�4;V+;�";�;�';�t;���:�)�:���:��:%��: ��:V�:;l�:x��:C�d:�4H:@/,:+�:���9m��9��~9~�9��58G�f�s��Ez��'���O7���#$��`<��nT��Wl�a��ݍ�����hR������땼��*Ⱥ��Ӻ�5ߺ��꺙!��4� �Cv�
#�Q���p�}�3�"�<G(�3�-�Zq3��9��>�}D�'�I�9:O�7�T�GVZ���_��ue�Nk�C�p�,)v�̼{�K���>r���<������ы�}����g���3��0 ��Ι��  �  <�=C3=�=�~=$=K�=Bn==�� =\ =7  =�H�<E��<���<��<�e�<��<!��<�7�<�|�<���<e�<G�<��<���<�	�<aH�<���<L��<���<z7�< p�<p��<[��<��<�D�<v�<���<{��<D��<�(�<?P�<Eu�<���<J��<���<���<��<��<�&�<o2�<�:�<�>�<�>�<�:�<r2�<q%�<��<���<#��<��<#��<�l�<�9�<�<
��<r|�<i0�<���<;��<$�<v��<,P�<[��< b�<���<�Z�<ξ<I;�<ɢ�<��<�`�<��<�	�<�V�<͞�<2�<
!�<�[�<J��< Ũ<M��<' �<�H�<�n�<���<Y��<�Л<��<;�<��<�6�<�K�<�_�<�q�<т�<���<(��<���<0��<�Ƃ<�р<p�}<��y<b�u<]�q< n<�j<V$f<�6b<CI^<�\Z<qV<��R<�N<��J<{�F<��B<B?<�$;<�E7<bi3<��/<��+<��'<$<�J <��<��<�<M<e�<��	<�J<��<�*�;
�;Z��;h��;��;U(�;�Z�;���;M��;�e�;�;���;0�; ��;�֠;�Κ;���;��;�R�;Ҳ�;[|;��q;�f;�w\;�>R;�8H;tf>;��4;gV+;�";�;?(;}u;{��:�*�:H��:`��:���:���:�W�: m�:
:��d:�6H:�/,:k�:���9���9�~99�9058g����(|�����c:���i&$��a<��qT�VYl����zލ�=����R�����H���2*Ⱥ��Ӻ�5ߺ�����z� ��u�n"�j���o���@�"�G(��-�|p3�K9��>�*D��I�`:O���T�2VZ���_��te�(k�3�p�*v�H�{�m����r���<��<���ы�����h���3��� ��nΙ��  �  /�=83=�=�~= $=T�=Tn==�� =\ =S  =�H�<���<��<�<f�<Y��<b��<�7�<�|�<���<y�<8G�<���<���<�	�<BH�<߅�<6��<w��<D7�<�o�<(��<��<��<|D�<�u�<o��<I��<
��<�(�<7P�<*u�<���<(��<���<���<�<�<�&�<�2�<�:�<?�<#?�<$;�<�2�<�%�<��<7��<g��<��<E��<�l�<�9�<3�<��<�|�<H0�<���<��<$�<]��<�O�<&��<�a�<Q��<�Z�<�;<;�<x��<g�<�`�<ﷶ<�	�<�V�<���<�<!�<�[�<l��<0Ũ<f��<G �<�H�<�n�<鑟<���<�Л<<�<��<��<�6�<�K�<�_�<�q�<�<���<4��<���<��<�Ƃ<xр<`�}<��y<��u<��q<r n<"j<�#f<6b<�H^<=\Z<�pV<)�R<�N<ĴJ<M�F<9�B<-?<%;< F7<�i3<��/<E�+<��'<�$<#K <�<�<�<�M<�<��	<QK<��<#+�;�
�;��;���;��;(�;UZ�;���;��;ge�;D�;��;�.�;+��;�ՠ;�͚;	��;��;�Q�;���;8Z|;{�q;W�f;	w\;�=R;Y9H;�f>;M�4;#W+;j";�	;o);�w;W��:�/�:6��:��:� �:���:�[�:Vo�:QĀ:ɧd:�8H:!3,:��:̍�9���9��~9�t9�58Eg����]���x����H�����.$��i<��zT��_l�I��]ߍ�T���T�����������(Ⱥ��Ӻ>3ߺ����k� �Lt�_ ����nm���0�"��D(��-��n3�@ 9���>�kD���I��9O���T�NVZ��_��ue��k�q�p�o+v��{�Z����s���=��^���ҋ�ʝ��
i���4��\���Ι��  �  �="3=�=�~=$=]�=gn=9=׷ =D\ =z  =I�<��<p��<��<bf�<¬�<���<"8�<}�<<��<��<XG�<��<���<�	�<5H�<���<��<��<�6�<�o�<Ԧ�<���<*�<D�<uu�<��<���<���<t(�<�O�< u�<o��<)��<���<���<!�<D�<�&�<�2�<;�<P?�<�?�<~;�<3�<&�<T�<���<���<j��<���<�l�<+:�<M�<��<x|�<B0�<j��<��<�#�<���<�O�<���<ta�<���<Z�<N;<�:�<��<�<j`�<���<�	�<uV�<���<�<!�<�[�<���<bŨ<���<� �<KI�<*o�<O��<���<Vћ<��<��<Y �<7�<NL�<�_�<4r�<��<���<3��<���<��<�Ƃ<Lр<Ŷ}<��y<P�u<1�q<��m<Kj<#f<35b<�G^<�[Z<	pV<��R<D�N<e�J<��F<3�B<*?<%;<EF7<�i3<_�/<չ+<��'<"$<�K <��<��<�<zN<Ŝ<8�	<L<��<M,�;��;���;��;��;7(�;;Z�;��;T��;d�; �;�~�;�-�;���;Ԡ;�̚;rޔ;M
�;�P�;Ű�;iW|;��q;*�f; v\;>R;f9H;�f>;Q�4;�X+;�";Y;L,;1z;k��:�5�:��:*��:=�::�`�: u�:wɀ:W�d:g?H:�6,:b�:��9n��9]�~98`9֟48'h�v! �����!���Pc����2;$�:v<���T��il�W��^卺�����V������ϗ��h)Ⱥ�Ӻe1ߺ�������� ��q���=���j�j��"��A(�B�-�/l3�s�8�_�>�oD���I�9O���T�WVZ���_��ve�dk�ޚp�.v���{������t��S?���	��iԋ�:���ij��6������ϙ��  �  ��=3=��=�~=%$=q�=|n=^=�� =u\ =�  =�I�<w��<���<  �<�f�<M��<6��<�8�<f}�<���<��<zG�<5��<���<�	�<H�<z��<���<���<�6�<o�<R��<4��<��<�C�<�t�<���<e��<\��<(�<�O�<�t�<C��<��<���<���<I�<|�<('�<)3�<v;�<�?�<@�< <�<�3�<�&�<��<'��<(��<���<ڙ�<m�<c:�<o�<,��<g|�<'0�<7��<���<v#�<���<6O�<8��<�`�<N��<�Y�<�̾<:�<���<��<`�<(��<8	�<4V�<h��<��<
!�<�[�<���<�Ũ<���<� �<�I�<�o�<ے�<w��<�ћ<�<i�<� �<�7�<�L�<@`�<�r�<L��<钊<J��<���<�<WƂ<р<�}<9�y<}�u<#�q<��m<6j<"f<4b<�F^<~ZZ<#oV<фR<��N<�J<��F<��B<?<,%;<�F7<Ij3<��/<b�+<u�'<$<�L <
�<��<<{O<�<E�	<M<l�<�-�;$�;J��;���;D�;(�;�Y�;:��;��;�b�;��;�|�;�+�;��;Ҡ;�ʚ;nܔ;w�;wN�;j��;�T|;I�q;��f;�t\;�=R;9H;
h>;��4;�Z+;�";�;�/;�};���:�=�:Y��:���:L�:'��:sh�:�{�:!΀:��d:GH:�;,:��:���9`��9̤~9�C9�48��h��L �����hڴ�7�湷���K$�C�<���T�,zl�x���ꍺ֨��oZ�����
���)Ⱥ��ӺE/ߺ ����9� ��m�������f����"��=(���-��h3�Q�8�8�>�D�F�I��7O���T��VZ���_��xe� 
k���p��0v���{�٬���v��yA������֋�)���wl���7�����?љ��  �  ό=�2=��=�~=,$=}�=�n=�=0� =�\ =�  =&J�<��<���<� �<g�<ۭ�<���<9�<�}�<���<D�<�G�<F��<���<p	�<�G�<@��<o��<i��<6�<�n�<Х�<���<�<�B�<Ut�<��<���<���<�'�<RO�<yt�<��<���<���<���<j�<��<�'�<�3�<�;�<H@�<�@�<�<�<14�<2'�<o�<���<���<O��<K��<~m�<�:�<��<9��<k|�<0�<��<[��<#�<��<�N�<���<W`�<���<�X�<̾<h9�<��<��<~_�<���<��<�U�<6��<��<!�<�[�<͒�<�Ũ<N��<O!�<6J�<p�<b��<��<wқ<��<	�<e!�<8�<(M�<�`�<�r�<���<��<[��<���<Ϻ�<'Ƃ<�Ѐ<v�}<I�y<r�u<�q<��m<�j<� f<�2b<�E^<sYZ<nV<ӃR<�N<8�J<�F<��B<�?<G%;<�F7<�j3<��/<>�+<[�'<'$<�M <>�<4�<;<�P<�<Z�	<N<[�<W/�;p�;Y��;/��;��;�'�;cY�;}��;L��;�a�;�;�z�;�)�;��;�Ϡ;EȚ;.ڔ;T�;�L�;t��;�Q|;�}q;S�f;�s\;�<R;�9H;�h>;��4;�\+; ";s;�3;2�;���:�G�:
��:A��:�:_��:�p�:���:�Հ:\�d:�OH:�@,:��:���9���9��~9�9S\38��i�"� ��߂�G���ª����k_$�љ<��T�g�l��#������\���@^�����Y���](Ⱥ��Ӻ�+ߺ��꺔���� ��i���u���a�B��"��8(���-�Ld3���8���>�sD�K�I� 7O��T��VZ��_�ze��k��p��4v���{�߮��Gy���C��X���؋�����n���9������ҙ��  �  ��=�2=��=�~=5$=��=�n=�=g� =�\ =A =�J�<���<<��<\!�<+h�<q��<R��<�9�<K~�<T��<��<�G�<c��<���<b	�<�G�<��<��<���<�5�<n�<-��<���<g�<PB�<�s�<\��<U��<T��<7'�<�N�<*t�<��<ζ�<���<���<��<�<�'�<4�<c<�<�@�<%A�<:=�<�4�<�'�<�<6��<=��<���<���<�m�<�:�<��<C��<f|�<�/�<���<
��<�"�<���<N�<��<�_�<���<2X�<i˾<�8�<O��<`�<�^�<B��<i�<�U�<��<��<	!�<�[�<��<ƨ<���<�!�<�J�<�p�<�<���< ӛ<g�<�	�<�!�<�8�<�M�<a�<s�<ԃ�<5��<m��<���<���<�ł<fЀ<��}<V�y<h�u<��q<;�m<�j<[f<�1b<qD^<6XZ<mV<ԂR<�N<z�J<��F<N�B<�?<e%;<G7<Sk3<�/<�+<I�'<M$<0O <|�<��<�	<5R<N�<��	<7O<[�<1�;��;���;���;��;�'�;�X�;���;���;�_�;.�; y�;�'�;(�;r͠;�Ś;�ה;��;wJ�;���;/N|;{q;�f;]r\;�;R;�9H;�i>;��4;_+;�"";�;j7;�;r�:R�:Z��:p��:�"�:���:jz�:{��:<܀:+�d:AXH:KH,:<�:h��9���9�y~9��9�28*sj�:� �|���(�����	��s$�]�<���T���l�(,������Z���Db��5��_����'Ⱥ�Ӻ�'ߺל꺋��&� ��e����h\������"��3(��-��_3��8�V�>�WD��I�{5O���T��VZ�B�_�{{e��k�K�p�L8v��{�:����{��RF����cۋ�.����p���;�����.ԙ��  �  ��=�2=��=�~=9$=��=�n=�=�� =&] =� =]K�<P��<���<
"�<�h�<��<���<&:�<�~�<���<��<(H�<���<���<R	�<�G�<���<���<���<(5�<m�<���<[��<��<�A�<s�<͢�<���<���<�&�<�N�<�s�<���<���<���<���<��<A�<3(�<v4�<�<�<gA�<�A�<�=�<�5�<�(�<��<���<���<C��<��<%n�<;�<��<X��<Z|�<�/�<���<���<H"�<,��<�M�<m��< _�<O��<wW�<�ʾ<	8�<���<��<k^�<˵�<�<OU�<���<��<!�<\�<0��<cƨ<��<,"�<4K�<Cq�<���<Y��<�ӛ<�<D
�<�"�<.9�<N�<�a�<}s�<��<`��<{��<���<���<�ł<)Ѐ<ٳ}<g�y<N�u<��q<
�m<cj<�f<E0b<9C^<�VZ<�kV<�R<-�N<��J<�F<��B<�?<u%;<fG7<�k3<ђ/<��+<J�'<[$<sP <ډ<��<<}S<��<��	<QP<`�<�2�;�;���;���;-	�;�'�;GX�;ɛ�;��;z^�;�߹;�v�;U%�;��;�ʠ;)Ú;`Ք;��;)H�;���;�J|;Kxq;U�f;�p\;O;R;�9H;Kj>;C�4;Ha+;�%";�;�;;s�;?�:�\�:���:���:-�:���:^��:瓏:Z�:��d:�`H:�M,:�:���9	��9(\~9��9��18RIk��!��)��M��1������$���<���T�_�l�f3��h�������f�����s����'Ⱥ��Ӻ�$ߺ���K��m� ��a�t���iW�x��Ĕ"��.(��-��[3�
�8��>�ID�S�I�/4O���T�YWZ�L�_��}e��k���p�<v�~�{�����Q~��I�����ދ�����Us��5>���	���ՙ��  �  [�=�2=��=�~==$=��=�n= =Ƹ =f] =� =�K�<��<s��<�"�<ai�<���<h��<�:�<9�<��<-�<VH�<���<���<A	�<wG�<���<p��<��<�4�<�l�<��<���<�<A�<kr�<D��<8��<O��<U&�<*N�<�s�<w��<���<���<��<��<��<�(�<�4�<n=�<�A�<QB�<o>�<6�< )�<B�<e �<C��<���<���<zn�<^;�<�<k��<H|�<�/�<W��<p��<�!�<���<M�<���<q^�<���<�V�<ʾ<b7�<��<*�<�]�<J��<��<U�<���<��<� �<4\�<Q��<�ƨ<Q��<�"�<�K�<�q�<(��<ﵝ<oԛ<��<�
�<!#�<�9�<�N�<�a�<�s�<H��<���<���<|��<x��<ył<�π<�}<��y<O�u<��q<��m<j<�f<�.b<B^<�UZ<�jV<��R<P�N<V�J<��F<��B<�?<�%;<�G7<&l3<��/<��+<M�'<m$<�Q <�<!�<c<�T<�<��	<kQ<\�<G4�;��;^��;O��;C	�;�'�;X�;���;���;�\�;�ݹ;�t�;m#�;��;�Ƞ;���;�Ҕ;���;@F�;���;�G|;Euq;R�f;8o\;�:R;�9H;!k>;��4;mc+;�(";�;@;��;��:�e�:��:��:�6�:>��:t��:��:3�:K�d:�iH:S,:#�:ي�9���9�F~9ɸ94#18�3l��O!�J���m���$��1��$��<�b�T�U�l�;����������j���	������O(Ⱥ��Ӻ5"ߺ������ܯ ��]������R�Q���"��)(���-�]W3���8�-~>��D���I��2O�,�T��WZ���_��e��k��p�x?v�w�{����������K���������㪎�au��C@��p���י��  �  6�=2=��=�~=F$=��=o==� =�] =� =bL�<d��<���<-#�<�i�<.��<���<;�<��<`��<e�<�H�<ɉ�<��<(	�<MG�<O��<%��<���<L4�<�l�<���<;��<��<�@�<�q�<���<���<���<&�<�M�<`s�<T��<���<���<��<�<��<�(�</5�<�=�<iB�<�B�<�>�<�6�<�)�<��<� �<���<��<՛�<�n�<�;�<1�<y��<G|�<|/�<)��<)��<�!�<Y��<�L�<`��<�]�<��<BV�<yɾ<�6�<���<� �<s]�<���<V�<�T�<f��<]�<� �<D\�<w��<�ƨ<���<�"�<L�<Fr�<���<w��<�ԛ<%�<Z�<�#�</:�<�N�<=b�<t�<~��<���<���<o��<Q��<Xł<�π<u�}<��y<^�u<��q<��m<!
j<�f<.b<�@^<�TZ<�iV<8�R<��N<��J<G�F<u�B<?<�%;<�G7<�l3<��/<N�+<��'<Y$<�R <�<<�<g<�U<��<	�	<GR<�<�5�;��;F �;���;�	�;s'�;�W�;X��;���;�[�;aܹ;)s�;`!�;��;�Ơ;ؾ�;є;v��;yD�;��;SE|;sq;Y�f;En\;:R;�9H;�k>;�4;Ie+;�*";�;�B;ȓ;��:�n�:��:6�:?�:+ƭ:�:ʡ�:��:_�d:�pH:~X,:��:���92�9�3~9)�9��08g�l��!�2h������vD��B�H�$���<�'�T���l��A��
���Ù��m�� ��v���Z'Ⱥ3�Ӻhߺ,�����0� ��Z�&���PN�p����"��%(��-��S3�_�8�v{>��D��I��1O���T�6XZ��_���e�%k�$�p�>Bv�4�{���������{M��C���⋻���nw��#B������ؙ��  �  �=m2=��=�~=F$=��=$o=5=� =�] =% =�L�<���<f��<�#�<Vj�<���<I��<_;�<��<���<��<�H�<ɉ�<��<*	�<2G�<#��<��<���<�3�<8l�<*��<���<5�<@�<�q�<L��<l��<���<�%�<�M�<+s�<6��<u��<���<��<0�<��<)�<�5�<>�<�B�<#C�<Y?�<�6�<�)�<-�<3�<��<e��<3��<�n�<�;�<L�<v��<F|�<o/�<��<��<<!�< ��<,L�<��<i]�<���<�U�<ɾ<o6�<��<Z �<]�<���<�<�T�<B��<V�<� �<>\�<���<Ǩ<���<B#�<[L�<�r�<���<ඝ<E՛<��<��<�#�<z:�<EO�<�b�<Dt�<���<���<���<y��<B��<7ł<]π<�}<%�y<��u<�q<��m<b	j<�f<>-b<!@^<5TZ<:iV<�R<0�N<?�J<��F<Q�B<�?<�%;<�G7<�l3<W�/<�+<��'<�$<=S <Ԍ<�<$<�V<��<��	<�R<ѳ<�6�;W�;�;���;�	�;�'�;7W�;ę�;���;�Z�;۹;r�;
 �;2�;(Š;#��;�ϔ;���;AC�;���;�B|;qq;��f;xm\;�9R;�9H;l>;��4;�f+;�,";�";LE;^�;B%�:u�:�:J�:�E�:�˭:8��:規:���:��d:WvH:[\,:�:���9>}�9�$~99608Kom��!��|�������Z��P���$�&�<���T�'�l�+G������Ǚ��p���������S'Ⱥ?�Ӻ�ߺ�������Q� �X�^�R���J����h�"��"(�I�-�,Q3���8��x>�+D�m�I��1O���T��WZ���_���e��k�E�p�Ev���{����_����N����䋻�����x��bC��U���ٙ��  �  �=Z2=��=�~=M$=��=/o=A="� =�] =A =�L�<��<���<�#�<�j�<˰�<���<�;�<��<���<��<�H�<��<��<	�< G�<��<̿�<c��<�3�<�k�<��<���<��<�?�<Eq�<��<)��<]��<�%�<~M�<s�<��<j��<���<1��<E�<��<)�<�5�<F>�<�B�<nC�<�?�<B7�<D*�<h�<}�<H��<���<C��<�n�<�;�<Z�<���<1|�<b/�<���<ف�<!�<ٹ�<L�<���<)]�<d��<�U�<�Ⱦ<6�<ܝ�< �<�\�<z��<��<tT�<+��<I�<� �<]\�<���<Ǩ<���<`#�<�L�<�r�<<��<��<�՛<��<��<>$�<�:�<zO�<�b�<\t�<Ǆ�<֓�<���<f��<4��<ł<Iπ<��}<��y<W�u<��q<z�m<�j<bf<�,b<�?^<�SZ<�hV<AR<�N<�J<��F<-�B<d?<�%;<7H7<m3<��/<�+<�'<i$<�S <`�<��<�<3W<@�<@�	<kS<,�<%7�;��;e�;���;�	�;z'�;�V�;X��;���;@Z�;�ڹ;q�;�;�;4Ġ;d��;�Δ;��;@B�;!��;�A|;Upq;N�f;ql\;n9R;[9H;�l>;��4;�g+;=-";)#;G;�;*�:y�:y�:��:zI�:ZЭ:X��:���:���:i�d:�yH:|^,:o�:��9�z�9n~9�u9��/8ʹm���!�����ź���n�X�[�$���<��U��l�pI��y��,ə�}r��'������'Ⱥ�Ӻ�ߺي�[���N� �;V������CI�^��g�"�� (��-�mO3�8�8�>x>�sD���I��0O��T��XZ��_���e��k�[�p��Ev�N�{����_���P�����+勻�����y��3D�����Xڙ��  �  	�=X2=��=|~=N$=��='o=Q=.� =�] =H =	M�<��<���<�#�<�j�<��<���<�;�<+��<���<��<�H�<��< ��<	�<"G�<��<���<G��<�3�<�k�<��<���<��<�?�<)q�<��<��<K��<x%�<bM�<s�<��<x��<���<9��<6�<�<@)�<�5�<\>�<�B�<�C�<�?�<]7�<b*�<r�<��<O��<���<U��<*o�<�;�<H�<���<*|�<i/�<���<ˁ�<!�<���<�K�<���<+]�<J��<sU�<�Ⱦ<6�<ޝ�<���<�\�<^��<��<iT�<(��<D�<� �<b\�<���<8Ǩ<��<w#�<�L�<�r�<S��<$��<�՛<��<�<N$�<�:�<�O�<�b�<�t�<���<Г�<���<Y��<>��<ł<?π<e�}<��y<#�u<a�q<��m<�j<f<l,b<�?^<�SZ<�hV<R<��N<��J<��F<9�B<K?<�%;<2H7<�l3<Ȕ/<F�+<8�'<�$<�S <}�<��<<RW<l�<S�	<�S<g�<�7�;G�;�;���;�	�;d'�;W�;O��;]��;�Y�;nڹ;�p�;�;��;�à;���;+Δ;��;�A�;ݣ�;A|;{oq;�f;el\;�9R;9H;%m>;�4;�g+;�.";�#;�G;V�;w+�:�y�:/�:��:$J�:�ѭ:؜�:ګ�:	��:��d:|H:g\,:æ:���9}�9�~9�o9,�/8t�m���!����������t�[���$���<�-U�O�l�1J����gʙ�s��C��K����'Ⱥ��Ӻ%ߺ��������� ��U�~��^���H�.����"�{ (���-�O3�l�8��w>�R
D��I��0O���T��XZ���_��e��k�f�p��Fv��{�B���S����P��h���勻�����y���D�����ڙ��  �  �=Z2=��=�~=M$=��=/o=A="� =�] =A =�L�<��<���<�#�<�j�<˰�<���<�;�<��<���<��<�H�<��<��<	�< G�<��<̿�<c��<�3�<�k�<��<���<��<�?�<Eq�<��<)��<]��<�%�<~M�<s�<��<j��<���<1��<E�<��<)�<�5�<F>�<�B�<nC�<�?�<B7�<D*�<h�<}�<H��<���<C��<�n�<�;�<Z�<���<1|�<b/�<���<ف�<!�<ٹ�<L�<���<)]�<d��<�U�<�Ⱦ<6�<ܝ�< �<�\�<z��<��<tT�<+��<I�<� �<]\�<���<Ǩ<���<`#�<�L�<�r�<<��<��<�՛<��<��<>$�<�:�<zO�<�b�<\t�<Ǆ�<֓�<���<f��<4��<ł<Iπ<��}<��y<W�u<��q<z�m<�j<bf<�,b<�?^<�SZ<�hV<AR<�N<�J<��F<-�B<d?<�%;<7H7<m3<��/<�+<�'<i$<�S <`�<��<�<3W<@�<@�	<kS<+�<$7�;��;e�;���;�	�;z'�;�V�;X��;���;@Z�;�ڹ;q�;�;�;4Ġ;d��;�Δ;��;@B�;!��;�A|;Upq;N�f;ql\;n9R;[9H;�l>;��4;�g+;=-";)#;G;�;*�:y�:y�:��:zI�:ZЭ:X��:���:���:i�d:�yH:|^,:o�:��9�z�9n~9�u9��/8ʹm���!�����ź���n�X�[�$���<��U��l�pI��y��,ə�}r��'������'Ⱥ�Ӻ�ߺي�[���N� �;V������CI�^��g�"�� (��-�mO3�8�8�>x>�sD���I��0O��T��XZ��_���e��k�[�p��Ev�N�{����_���P�����+勻�����y��3D�����Xڙ��  �  �=m2=��=�~=F$=��=$o=5=� =�] =% =�L�<���<f��<�#�<Vj�<���<I��<_;�<��<���<��<�H�<ɉ�<��<*	�<2G�<#��<��<���<�3�<8l�<*��<���<5�<@�<�q�<L��<l��<���<�%�<�M�<+s�<6��<u��<���<��<0�<��<)�<�5�<>�<�B�<#C�<Y?�<�6�<�)�<-�<3�<��<e��<3��<�n�<�;�<L�<v��<F|�<o/�<��<��<<!�< ��<,L�<��<i]�<���<�U�<ɾ<o6�<��<Z �<]�<���<�<�T�<B��<V�<� �<>\�<���<Ǩ<���<B#�<[L�<�r�<���<ඝ<E՛<��<��<�#�<z:�<EO�<�b�<Dt�<���<���<���<y��<B��<7ł<]π<�}<%�y<��u<�q<��m<b	j<�f<>-b<!@^<5TZ<:iV<�R<0�N<?�J<��F<Q�B<�?<�%;<�G7<�l3<W�/<�+<��'<�$<=S <Ԍ<�<$<�V<��<��	<�R<ѳ<�6�;W�;�;���;�	�;�'�;7W�;ę�;���;�Z�;۹;r�;
 �;2�;(Š;#��;�ϔ;���;AC�;���;�B|;qq;��f;xm\;�9R;�9H;l>;��4;�f+;�,";�";LE;^�;B%�:u�:�:J�:�E�:�˭:8��:規:���:��d:WvH:[\,:�:���9>}�9�$~99608Kom��!��|�������Z��P���$�&�<���T�'�l�+G������Ǚ��p���������S'Ⱥ?�Ӻ�ߺ�������Q� �X�^�R���J����h�"��"(�I�-�,Q3���8��x>�+D�m�I��1O���T��WZ���_���e��k�E�p�Ev���{����_����N����䋻�����x��bC��U���ٙ��  �  6�=2=��=�~=F$=��=o==� =�] =� =bL�<d��<���<-#�<�i�<.��<���<;�<��<`��<e�<�H�<ɉ�<��<(	�<MG�<O��<%��<���<L4�<�l�<���<;��<��<�@�<�q�<���<���<���<&�<�M�<`s�<T��<���<���<��<�<��<�(�</5�<�=�<iB�<�B�<�>�<�6�<�)�<��<� �<���<��<՛�<�n�<�;�<1�<y��<H|�<|/�<)��<)��<�!�<Y��<�L�<`��<�]�<��<BV�<yɾ<�6�<���<� �<s]�<���<V�<�T�<f��<]�<� �<D\�<w��<�ƨ<���<�"�<L�<Fr�<���<w��<�ԛ<%�<Z�<�#�</:�<�N�<=b�<t�<~��<���<���<o��<Q��<Xł<�π<u�}<��y<^�u<��q<��m<!
j<�f<.b<�@^<�TZ<�iV<8�R<��N<��J<G�F<u�B<?<�%;<�G7<�l3<��/<N�+<��'<Y$<�R <�<<�<g<�U<��<	�	<GR<�<�5�;��;F �;���;�	�;s'�;�W�;X��;���;�[�;aܹ;)s�;`!�;��;�Ơ;ؾ�;є;v��;yD�;��;SE|;sq;Y�f;En\;:R;�9H;�k>;�4;Ie+;�*";�;�B;ȓ;��:�n�:��:6�:?�:+ƭ:�:ʡ�:��:_�d:�pH:~X,:��:���92�9�3~9)�9��08h�l��!�2h������vD��B�H�$���<�'�T���l��A��
���Ù��m�� ��v���Z'Ⱥ3�Ӻhߺ,�����0� ��Z�&���PN�p����"��%(��-��S3�_�8�v{>��D��I��1O���T�6XZ��_���e�%k�$�p�>Bv�4�{���������{M��C���⋻���nw��#B������ؙ��  �  [�=�2=��=�~==$=��=�n= =Ƹ =f] =� =�K�<��<s��<�"�<ai�<���<h��<�:�<9�<��<-�<VH�<���<���<A	�<wG�<���<p��<��<�4�<�l�<��<���<�<A�<kr�<D��<8��<O��<U&�<*N�<�s�<w��<���<���<��<��<��<�(�<�4�<n=�<�A�<QB�<o>�<6�< )�<B�<e �<C��<���<���<zn�<^;�<�<k��<H|�<�/�<W��<q��<�!�<���<M�<���<q^�<���<�V�<ʾ<b7�<��<*�<�]�<J��<��<U�<���<��<� �<5\�<Q��<�ƨ<Q��<�"�<�K�<�q�<(��<ﵝ<oԛ<��<�
�<!#�<�9�<�N�<�a�<�s�<H��<���<���<|��<x��<ył<�π<�}<��y<O�u<��q<��m<j<�f<�.b<B^<�UZ<�jV<��R<Q�N<V�J<��F<��B<�?<�%;<�G7<&l3<��/<��+<M�'<m$<�Q <�<!�<c<�T<�<��	<kQ<\�<G4�;��;^��;O��;C	�;�'�;X�;���;���;�\�;�ݹ;�t�;m#�;��;�Ƞ;���;�Ҕ;���;@F�;���;�G|;Euq;R�f;8o\;�:R;�9H;!k>;��4;mc+;�(";�;@;��;��:�e�:��:��:�6�:>��:t��:��:3�:K�d:�iH:S,:#�:ي�9���9�F~9ɸ94#18�3l��O!�J���m���$��1��$��<�b�T�U�l�;����������j���	������O(Ⱥ��Ӻ5"ߺ������ܯ ��]������R�Q���"��)(���-�]W3���8�-~>��D���I��2O�,�T��WZ���_��e��k��p�x?v�w�{����������K���������㪎�au��C@��p���י��  �  ��=�2=��=�~=9$=��=�n=�=�� =&] =� =]K�<P��<���<
"�<�h�<��<���<&:�<�~�<���<��<(H�<���<���<R	�<�G�<���<���<���<(5�<m�<���<[��<��<�A�<s�<͢�<���<���<�&�<�N�<�s�<���<���<���<���<��<A�<3(�<v4�<�<�<gA�<�A�<�=�<�5�<�(�<��<���<���<C��<��<%n�<;�<��<X��<Z|�<�/�<���<���<H"�<,��<�M�<m��< _�<O��<wW�<�ʾ<
8�<���<��<k^�<˵�<�<PU�<���<��<!�<\�<0��<cƨ<��<,"�<4K�<Cq�<���<Y��<�ӛ<�<D
�<�"�<.9�<N�<�a�<}s�<��<`��<{��<���<���<�ł<)Ѐ<ٳ}<g�y<N�u<��q<
�m<cj<�f<E0b<9C^<�VZ<�kV<�R<-�N<��J< �F<��B<�?<u%;<fG7<�k3<Ғ/<��+<J�'<[$<sP <ډ<��<<}S<��<��	<QP<`�<�2�;�;���;���;-	�;�'�;GX�;ț�;��;z^�;�߹;�v�;U%�;��;�ʠ;)Ú;`Ք;��;)H�;���;�J|;Kxq;U�f;�p\;O;R;�9H;Kj>;C�4;Ha+;�%";�;�;;s�;?�:�\�:���:���:-�:���:^��:瓏:Z�:��d:�`H:�M,:�:���9	��9(\~9��9��18RIk��!��)��M��1������$���<���T�_�l�f3��h�������f�����s����'Ⱥ��Ӻ�$ߺ���K��m� ��a�t���iW�x��Ĕ"��.(��-��[3�
�8��>�ID�S�I�/4O���T�YWZ�L�_��}e��k���p�<v�~�{�����Q~��I�����ދ�����Us��5>���	���ՙ��  �  ��=�2=��=�~=5$=��=�n=�=g� =�\ =A =�J�<���<<��<\!�<+h�<q��<R��<�9�<K~�<T��<��<�G�<c��<���<b	�<�G�<��<��<���<�5�<n�<-��<���<g�<PB�<�s�<\��<U��<T��<7'�<�N�<*t�<��<ζ�<���<���<��<�<�'�<4�<c<�<�@�<%A�<:=�<�4�<�'�<�<6��<=��<���<���<�m�<�:�<��<C��<f|�<�/�<���<
��<�"�<���<N�<��<�_�<���<2X�<i˾<�8�<O��<`�<�^�<B��<i�<�U�<��<��<
!�<�[�<��<ƨ<���<�!�<�J�<�p�<�<���< ӛ<g�<�	�<�!�<�8�<�M�<a�<s�<ԃ�<5��<m��<���<���<�ł<fЀ<��}<U�y<h�u<��q<;�m<�j<[f<�1b<qD^<6XZ<mV<ԂR<�N<z�J<��F<N�B<�?<e%;<G7<Sk3<�/<�+<I�'<M$<0O <|�<��<�	<5R<N�<��	<7O<[�<1�;��;���;���;��;�'�;�X�;���;���;�_�;.�; y�;�'�;(�;r͠;�Ś;�ה;��;wJ�;���;.N|;{q;�f;]r\;�;R;�9H;�i>;��4;_+;�"";�;j7;�;r�:R�:Z��:p��:�"�:���:jz�:{��:<܀:+�d:AXH:KH,:<�:h��9���9�y~9��9�28*sj�:� �|���(�����	��s$�]�<���T���l�(,������Z���Db��5��_����'Ⱥ�Ӻ�'ߺל꺋��&� ��e����h\������"��3(��-��_3��8�V�>�WD��I�{5O���T��VZ�B�_�{{e��k�K�p�L8v��{�:����{��RF����cۋ�.����p���;�����.ԙ��  �  ό=�2=��=�~=,$=}�=�n=�=0� =�\ =�  =&J�<��<���<� �<g�<ۭ�<���<9�<�}�<���<D�<�G�<F��<���<p	�<�G�<@��<o��<i��<6�<�n�<Х�<���<�<�B�<Ut�<��<���<���<�'�<RO�<yt�<��<���<���<���<j�<��<�'�<�3�<�;�<H@�<�@�<�<�<14�<2'�<o�<���<���<O��<K��<~m�<�:�<��<9��<k|�<0�<��<[��<#�<��<�N�<���<W`�<���<�X�<̾<h9�<��<��<~_�<���<��<�U�<6��<��<!�<�[�<͒�<�Ũ<N��<O!�<6J�<p�<b��<��<wқ<��<	�<e!�<8�<(M�<�`�<�r�<���<��<[��<���<Ϻ�<'Ƃ<�Ѐ<v�}<I�y<r�u<�q<��m<�j<� f<�2b<�E^<sYZ<nV<ӃR<�N<8�J<�F<��B<�?<G%;<�F7<�j3<��/<>�+<[�'<'$<�M <>�<4�<;<�P<�<Z�	<N<[�<W/�;p�;Y��;.��;��;�'�;cY�;}��;L��;�a�;�;�z�;�)�;��;�Ϡ;EȚ;.ڔ;T�;�L�;t��;�Q|;�}q;S�f;�s\;�<R;�9H;�h>;��4;�\+; ";s;�3;2�;���:�G�:
��:A��:�:_��:�p�:���:�Հ:\�d:�OH:�@,:��:���9���9��~9�9S\38��i�"� ��߂�G���ª����k_$�љ<��T�g�l��#������\���@^�����Y���](Ⱥ��Ӻ�+ߺ��꺔���� ��i���u���a�B��"��8(���-�Ld3���8���>�sD�K�I� 7O��T��VZ��_�ze��k��p��4v���{�߮��Gy���C��X���؋�����n���9������ҙ��  �  ��=3=��=�~=%$=q�=|n=^=�� =u\ =�  =�I�<w��<���<  �<�f�<M��<6��<�8�<f}�<���<��<zG�<5��<���<�	�<H�<z��<���<���<�6�<o�<R��<4��<��<�C�<�t�<���<e��<\��<(�<�O�<�t�<C��<��<���<���<I�<|�<('�<)3�<v;�<�?�<@�< <�<�3�<�&�<��<'��<(��<���<ڙ�<m�<c:�<o�<,��<g|�<'0�<7��<���<v#�<���<6O�<8��<�`�<N��<�Y�<�̾<:�<���<��<`�<(��<8	�<4V�<h��<��<
!�<�[�<���<�Ũ<���<� �<�I�<�o�<ے�<w��<�ћ<�<i�<� �<�7�<�L�<@`�<�r�<L��<钊<J��<���<�<WƂ<р<�}<9�y<}�u<#�q<��m<6j<"f<4b<�F^<~ZZ<#oV<фR<��N<�J<��F<��B<?<,%;<�F7<Jj3<��/<b�+<u�'<$<�L <
�<��<<{O<�<E�	<M<l�<�-�;$�;J��;���;D�;(�;�Y�;:��;��;�b�;��;�|�;�+�;��;Ҡ;�ʚ;nܔ;w�;wN�;j��;�T|;I�q;��f;�t\;�=R;9H;
h>;��4;�Z+;�";�;�/;�};���:�=�:Y��:���:L�:'��:sh�:�{�:!΀:��d:GH:�;,:��:���9`��9̤~9�C9�48��h��L �����hڴ�7�湷���K$�C�<���T�,zl�x���ꍺ֨��oZ�����
���)Ⱥ��ӺE/ߺ ����9� ��m�������f����"��=(���-��h3�Q�8�8�>�D�F�I��7O���T��VZ���_��xe� 
k���p��0v���{�٬���v��yA������֋�)���wl���7�����?љ��  �  �="3=�=�~=$=]�=gn=9=׷ =D\ =z  =I�<��<p��<��<bf�<¬�<���<"8�<}�<<��<��<XG�<��<���<�	�<5H�<���<��<��<�6�<�o�<Ԧ�<���<*�<D�<uu�<��<���<���<t(�<�O�< u�<o��<)��<���<���<!�<D�<�&�<�2�<;�<P?�<�?�<~;�<3�<&�<T�<���<���<j��<���<�l�<+:�<M�<��<x|�<B0�<j��<��<�#�<���<�O�<���<ta�<���<Z�<N;<�:�<��<�<j`�<���<�	�<uV�<���<�<!�<�[�<���<bŨ<���<� �<KI�<*o�<O��<���<Vћ<��<��<Y �<7�<NL�<�_�<4r�<��<���<3��<���<��<�Ƃ<Lр<Ŷ}<��y<P�u<1�q<��m<Kj<#f<35b<�G^<�[Z<	pV<��R<D�N<e�J<��F<3�B<*?<%;<FF7<�i3<_�/<չ+<��'<"$<�K <��<��<�<zN<Ŝ<8�	<L<��<M,�;��;���;��;��;7(�;;Z�;��;T��;d�; �;�~�;�-�;���;Ԡ;�̚;rޔ;M
�;�P�;Ű�;iW|;��q;*�f; v\;>R;f9H;�f>;Q�4;�X+;�";Y;L,;1z;k��:�5�:��:*��:=�::�`�: u�:wɀ:W�d:g?H:�6,:b�:��9n��9]�~98`9֟48'h�v! �����!���Pc����2;$�:v<���T��il�W��^卺�����V������ϗ��h)Ⱥ�Ӻe1ߺ�������� ��q���=���j�j��"��A(�B�-�/l3�s�8�_�>�oD���I�9O���T�WVZ���_��ve�dk�ޚp�.v���{������t��S?���	��iԋ�:���ij��6������ϙ��  �  /�=83=�=�~= $=T�=Tn==�� =\ =S  =�H�<���<��<�<f�<Y��<b��<�7�<�|�<���<y�<8G�<���<���<�	�<BH�<߅�<6��<w��<D7�<�o�<(��<��<��<|D�<�u�<o��<I��<
��<�(�<7P�<*u�<���<(��<���<���<�<�<�&�<�2�<�:�<?�<#?�<$;�<�2�<�%�<��<7��<g��<��<E��<�l�<�9�<3�<��<�|�<H0�<���<��<$�<]��<�O�<&��<�a�<Q��<�Z�<�;<;�<y��<g�<�`�<ﷶ<�	�<�V�<���<�<!�<�[�<l��<0Ũ<f��<G �<�H�<�n�<鑟<���<�Л<<�<��<��<�6�<�K�<�_�<�q�<�<���<4��<���<��<�Ƃ<xр<`�}<��y<��u<��q<r n<"j<�#f<6b<�H^<=\Z<�pV<)�R<�N<ĴJ<M�F<9�B<-?<%;< F7<�i3<��/<E�+<��'<�$<#K <�<�<�<�M<�<��	<QK<��<#+�;�
�;��;���;��;(�;UZ�;���;��;ge�;D�;��;�.�;+��;�ՠ;�͚;	��;��;�Q�;���;8Z|;{�q;W�f;	w\;�=R;Y9H;�f>;M�4;#W+;j";�	;o);�w;W��:�/�:6��:��:� �:���:�[�:Vo�:QĀ:ɧd:�8H:!3,:��:̍�9���9��~9�t9�58Eg����]���x����H�����.$��i<��zT��_l�I��]ߍ�T���T�����������(Ⱥ��Ӻ>3ߺ����k� �Lt�_ ����nm���0�"��D(��-��n3�@ 9���>�kD���I��9O���T�NVZ��_��ue��k�q�p�o+v��{�Z����s���=��^���ҋ�ʝ��
i���4��\���Ι��  �  <�=C3=�=�~=$=K�=Bn==�� =\ =7  =�H�<E��<���<��<�e�<��<!��<�7�<�|�<���<e�<G�<��<���<�	�<aH�<���<L��<���<z7�< p�<p��<[��<��<�D�<v�<���<{��<D��<�(�<?P�<Eu�<���<J��<���<���<��<��<�&�<o2�<�:�<�>�<�>�<�:�<r2�<q%�<��<���<#��<��<#��<�l�<�9�<�<
��<r|�<i0�<���<;��<$�<v��<,P�<[��< b�<���<�Z�<ξ<I;�<ɢ�<��<�`�<��<�	�<�V�<͞�<2�<
!�<�[�<J��< Ũ<M��<' �<�H�<�n�<���<Y��<�Л<��<;�<��<�6�<�K�<�_�<�q�<т�<���<(��<���<0��<�Ƃ<�р<p�}<��y<b�u<]�q< n<�j<V$f<�6b<CI^<�\Z<qV<��R<�N<��J<{�F<��B<B?<�$;<�E7<bi3<��/<��+<��'<$<�J <��<��<�<M<e�<��	<�J<��<�*�;
�;Z��;h��;��;U(�;�Z�;���;M��;�e�;�;���;0�; ��;�֠;�Κ;���;��;�R�;Ҳ�;[|;��q;�f;�w\;�>R;�8H;tf>;��4;gV+;�";�;?(;}u;{��:�*�:H��:`��:���:���:�W�: m�:
:��d:�6H:�/,:k�:���9���9�~99�9058g����(|�����c:���i&$��a<��qT�VYl����zލ�=����R�����H���2*Ⱥ��Ӻ�5ߺ�����z� ��u�n"�j���o���@�"�G(��-�|p3�K9��>�*D��I�`:O���T�2VZ���_��te�(k�3�p�*v�H�{�m����r���<��<���ы�����h���3��� ��nΙ��  �  ߏ=76=z�=��=R(=��=Bs=t=Z� =.b =� =�V�<Q��<���</0�<%x�<��<j�<bN�<���<���<; �<�d�<?��<���<�,�<�l�<b��<���<�'�<�c�<���<L��<I�<�E�<"{�<���<���<��<B?�<zk�<���<&��<���<X�<�#�<�?�<�X�<kn�<~��<��<���<U��<.��<���<���<<��<��<�m�<1T�<@5�<��<���<#��<�}�<@�<���<E��<�]�<��<���<J=�<R��<kZ�<��<�\�<���<�E�<��<e�<�u�<�ϸ<$�<<s�<��<��< B�<�}�<δ�<��<�<wB�<�j�<���<ʱ�<Yџ<R�<L	�<"�<9�<tN�<�a�<6t�<ۄ�<J��<E��<��<���<Dņ<�΄<Eׂ<J߀<��}<��y<	�u<��q<o�m<�j<�f<� b<z-^<�:Z<UIV<�XR<iN<�{J<w�F<G�B<ٹ><��:<g�6<	3<�(/<�J+<�p'<љ#<��<��<s0<�l<t�<h�<aD	<ј<T�<@��;]��;�c�;�V�;�Y�;o�;%��;��;'�;�~�;.��;d��;�+�;��;�;���;���; �;)*�;(��;�x;>,m;�b;& X;��M;��C;<!:;)�0;�$';��;��;\;�{;��:B��:�J�:�g�:�ӵ:c��:.��:Bو:��t:-KX:F<:9� :`h:��9��9�V9���8�-7k[��oB�j)��^�Ĺ����#��D+��7C�\�Z�@�r��������^[����~��g���Xwʺ�պ,T��������r\����L��6:�R���c#���(��}.��4���9��?��D��J���O�"U��Z��-`���e�+>k���p�LUv�5�{�����C~��GE��	��uӋ������b���*��p�s����  �  ď=;6=y�=��=V(=��=Js=x=i� =8b =� =�V�<Z��<���<?0�<Jx�<��<�<�N�<��<���<A �<�d�<M��<���<r,�<�l�<Z��<���<�'�<bc�<���<N��<;�<�E�<{�<���<���<��<.?�<ak�<W��<��<��<B�<�#�<�?�<�X�<yn�<���<��<���<u��<"��<���<ƛ�<N��<��<�m�<NT�<[5�<��<��<0��<�}�<%@�<���<+��<�]�<��<L��<.=�<4��<mZ�<���<�\�<���<�E�<��<b�<�u�<�ϸ<�#�<�r�<���<��<B�<�}�<۴�<��<�<�B�<�j�<���<㱡<Xџ<w�<Z	�<3"�<%9�<rN�<b�<Kt�<���<T��<T��<'��<���<5ņ<�΄<Rׂ<߀<O�}<��y<��u<��q<B�m<�j<mf<� b<R-^<�:Z<KIV<�XR<7iN<4{J<��F<C�B<��><�:<��6<'	3<�(/<�J+<�p'<�#<��<��<�0<�l<®<p�<�D	<�<��<­�;x��;d�;W�;Z�;�n�;K��;��;4�;u~�;���;x��;�+�;t�;j;E��;w��;��;=*�;߇�;�x;�*m;�b;� X;8�M;a�C;�!:;�0;%';3�;l�; ;�|;��:΂�:>L�: i�:�յ:���:��:�ڈ:�t:�NX:�G<:s� :7j:�9{�9��V9���8�R 7Su���|B�^(���Ĺd���&'��F+�&9C�|�Z�ʟr����?���b_����G}�����Ewʺ�պ�Rẅ�����)���[����I��9�����b#�U�(��}.��4��9�?���D��J��O��!U�h�Z�.`��e��?k���p�;Vv���{������~���E������Ӌ�
����b���*���� ����  �  ��=16=p�=��=X(=��=[s=�=�� =Ob =� = W�<���<V��<�0�<�x�<]��<��<�N�<C��<3��<] �<�d�<N��<���<f,�<�l�<@��<W��<t'�<c�<���<���<��<�E�<�z�<S��<@��<��<�>�<:k�<>��<ټ�<���<*�<�#�<�?�<�X�<�n�<���<=��<��<נ�<u��<��<��<���<x��<n�<�T�<�5�<��<0��<D��< ~�<!@�<���<��<�]�<q�<*��<
=�<���<Z�<���<�\�<��<vE�<���<��<yu�<Kϸ<�#�<�r�<Ѽ�<��<�A�<�}�<մ�<��<+�<�B�<�j�<��<A��<�џ<��<�	�<�"�<�9�<�N�<yb�<|t�<3��<z��<v��<2��<���<:ņ<�΄<Cׂ<�ހ<*�}<!�y<F�u<�q<u�m<!j<�f<�b<�,^<(:Z<�HV<3XR<iN<�zJ<]�F<�B<��><�:<��6<k	3<�(/<hK+<q'<Ě#<\�<m�<�1<�m<��<+�<SE	<��<��<���;���;�d�;-W�;KZ�;�n�;��;���;��;F~�;���;<��;d*�;�;,��;ܲ�;[��;@�;�(�;|��;� x;�)m;ǉb;� X;��M;��C;�!:;��0;�%';��;B�;� ;�;L�:��:�Q�:Hn�:ݵ:ٔ�:X��:�ވ:"�t:�TX:�J<:�� :$j:��9Fߟ9�V9���8���6����U�B�;>���Ĺ�����2�CR+�+DC��[�S�r����a����a������]~��C���qvʺ;�պ�P���n�����<Y��������5�����_#���(�{.��4�\�9�2?���D�zJ���O��!U�C�Z��.`���e�Ak�x�p��Wv�>�{�-���2����F�����ԋ�����d��;,������B����  �  ��=6=`�=��=](=	�={s=�=�� =�b =4 =yW�<;��<���<1�<+y�<���<K�<7O�<���<���<� �<e�<h��<���<m,�<�l�<��<��<'�<�b�<@��<o��<l�<�D�<z�<ԭ�<���< �<w>�<�j�<��<���<���<"�<�#�<�?�<Y�<�n�<��<���<V��<;��<���<��<���<(��<��<�n�<U�<�5�<F�<��<���<2~�<%@�<���<��<�]�<*�<̣�<�<�<q��<�Y�<��<\�<���<�D�<3��<o�<u�<�θ<^#�<}r�<���<��<�A�<�}�<ߴ�<+�<u�<C�<Yk�<j��<���<,ҟ<T�<6
�<#�<:�<HO�<�b�<�t�<���<Δ�<���<[��<ʺ�<@ņ<�΄<ׂ<�ހ<^�}<W�y<��u<1�q<��m<j<�f<�b<�+^<=9Z<�GV<gWR<9hN<KzJ<ӍF<٢B<��>< �:<��6<�	3<�)/< L+<�q'<��#<U�<o�<�2<�n<��<:�<<F	<��<��<8��;\��;�e�;�W�;�Z�;�n�;���;���;��;�|�;7��;ɂ�;�(�;k�;!��;ɰ�;{��;��;Q'�;+��;l�w;A'm;�b;�X;u�M;B�C;F":;M�0;C(';`�;��;E$;�;��:��:MZ�:w�:��:v��:П�:Z�:��t:#_X:�S<:�� :vk:�
�98ߟ9A�V9�U�8�y�6���-�B�	X����Ĺ����wD�uc+�YRC��[�Ͷr�����Ɛ�=f������H�������7vʺ"�պ M���'
��/���U�r�����2�����[#�K�(�$w.�p 4���9�9?� �D��J�c�O�A!U�#�Z�}/`���e�1Ck���p�[v�:�{�캀������H��?��׋�Z����e���-��t���꿙��  �  h�=�5=P�=w�=i(=%�=�s=�=� =�b =~ = X�<��<���<�1�<�y�<���<��<�O�<;��<���<� �<.e�<���<���<O,�<�l�<ë�<���<�&�<9b�<���<���<��<=D�<cy�<��<!��<x�<�=�<Sj�<x��<V��<���<�<�#�<@�<JY�<o�<b��<��<��<͡�<���<.��<]��<��<���<Mo�<�U�<�6�<��<���<���<V~�<M@�<t��<߯�<W]�<��<^��<<�<���<�X�<P��<A[�<���<D�<k��<��<Yt�<Zθ<�"�<r�<=��<]�<�A�<�}�<��<K�<��<lC�<�k�<���<A��<�ҟ<��<�
�<�#�<�:�<�O�<vc�<�u�<���<��<䢌<���<꺈<'ņ<p΄<�ւ<gހ<}�}<^�y<^�u<��q<1�m<j<)f<Pb<<*^<�7Z<�FV<iVR<IgN<�yJ<d�F<��B<y�><N�:<G�6<>
3<*/<�L+<'s'<˜#<��<��<�3<_p<�<��<�G	<��<�<ձ�;���;�f�;�X�;�Z�;�n�;/��;��;��;�z�;m�;r��;4&�;��;X��;��;���;�;�$�;2��;��w;/$m;�b;�X;��M;��C;�#:;ݍ0;*';�;'�;H);Շ;V*�:G��:Lf�:V��:�:��:*��:4�:�t:�iX:[<:� :zq:?�9�ן9�V9��8�E�6�}��dC������ŹE��C[��z+��iC�l/[�m�r��!��Hΐ��k����������� ��Fvʺ��պrJ�@�캃��
��&Q��������,����V#���(��q.���3�"�9�
?���D�J���O�K U���Z�l0`�+�e�OEk�/�p��^v���{����������K����ڋ����h��!0��`��������  �  -�=�5=:�=p�=s(=5�=�s==/� =c =� =�X�<���<V��<�2�<�z�<[��<�	�<}P�<Ŗ�<u��<d!�<|e�<���<���<5,�<bl�<f��<I��<&�<�a�<��<��<��<wC�<�x�<K��<g��<��<<=�<�i�<��<��<J��<��<�#�<.@�<sY�<qo�<��<���<���<~��<]��<��<%��<���<j��<�o�<RV�<47�<1�<M��<��<~~�<f@�<p��<���<]�<e�<��<�;�<"��<&X�<���<gZ�<���<FC�<���<��<�s�<�͸<W"�<�q�<ϻ�<�<�A�<�}�<&��<��<�<�C�<Vl�<���<ﳡ<�ӟ<��<��<�$�<�;�<�P�<%d�<v�<���<���<H��<���<��< ņ<E΄<�ւ<�݀<��}<3�y<��u<h�q<��m<�j<�f<�b<�(^<i6Z<1EV<)UR<ffN<�xJ<��F<3�B<Z�><r�:<��6<�
3<+/<N+<Mt'<.�#<�<��<�5<�q<ų<Y�<I	<K�<-�<A��;���;�g�;uY�;5[�;Nn�;���;���;��;Zy�;�;�}�;z#�;��;m��;#��;���;Cߌ;"�;���;��w;!m;΂b;�X;��M;��C;�$:;]�0;l-';b�;z�;~.;��;�5�:+��:'s�:��:��:9��:���:���:��t:�zX:Yh<:� :�u:��9I͟9�jV9���8}�6����rC�
���W0Ź�B��rt���+��C�]F[�6�r�:,��gՐ��r������������yuʺv�պ"F�������צ��K����ԋ��%�����O#��(�$l.�n�3�s~9��?���D�J���O��U�8�Z��1`���e��Hk���p��cv�V�{�s���ȇ���N����(݋�B���ek���2������qÙ��  �  ��=�5=!�=l�=|(=N�=�s=G=t� =fc =; =�Y�<���<<��<�3�<�{�<.��<y
�<=Q�<]��<���<�!�<�e�<��<��<$,�<,l�<��<���<z%�<�`�<?��<=��<�<�B�<�w�<u��<���<�<�<�<i�<���<���<��<��<�#�<A@�<�Y�<�o�<T��<.��<7��<R��<0��<ڤ�<��<���<?��<�p�<(W�<�7�<��<���<x��<�~�<s@�<o��<���<�\�<�<W��<�:�<n��<cW�<���<�Y�<���<SB�<���<�<�r�<�̸<�!�<q�<s��<� �<uA�<�}�<8��<��<j�<gD�<�l�<S��<Ĵ�<lԟ<��<��<{%�<`<�<|Q�<�d�<�v�<��<��<���<���<��<ņ<΄<Gւ<�݀<��}<��y<��u<��q<��m<=j<�f<b<�&^<�4Z<�CV<�SR<7eN<�wJ<)�F<ȡB<C�><��:<��6<�3<�+/<)O+<�u'<џ#<��<> <�7<�s<��<�<�J	<�<v�<{��;U��;�i�;BZ�;�[�;Cn�;��;���;_�;w�;��;S{�;h �;{ޤ;��;���;w��;�ی;_�;~�;��w;3m;+�b;X;��M;I�C;�%:;��0;�0';� ;l;�3;Z�;0C�:���:u��:���:�
�:���:K:m�:3u:��X:�t<:�� :�x:G
�9Rǟ9gKV9�P�8�q�6&����C��ܓ�YgŹ�x��V����+���C�3a[��r��6���ߐ�tz��|��v�������tʺ��պ�@���������#F���!�������cH#�k�(��e.���3�ry9�
?�_�D�J���O�U�c�Z�,3`���e�'Lk��p�iv���{�wÀ�;���aR�������������zn���5�������ř��  �  ǎ=|5=
�=d�=�(=g�=t=}=�� =�c =� =qZ�<l��<��<p4�<q|�<��<8�<�Q�<��<���<*"�<f�<��<��<,�<�k�<���<o��<�$�<H`�<l��<j��<:�<�A�<�v�<���<���<+�<�;�<�h�<	��<&��<���<��<�#�<U@�<�Y�<"p�<͂�<ב�<ۜ�<���<��<���<��<j��<��<�q�<�W�<v8�<p�<3��<¶�<�~�<�@�<Z��<c��<f\�<��<ҡ�<:�<���<xV�<���<�X�<
��<_A�<���<+�<�q�<7̸<� �<�p�< ��<~ �<TA�<{}�<M��<�<��<�D�<�m�<�<z��<F՟<��<�<[&�<9=�<IR�<�e�<iw�<���<y��<���<,��<(��<ņ<�̈́<�Ղ<.݀<��}<��y<!�u</�q<<�m<l j<�f<0b<6%^<3Z<9BV<�RR<dN<wJ<f�F<g�B<�><��:<L�6<@3<�,/<WP+<�v'<-�#<n�< <Q9<�u<j�<��<lL	<K�<��<߸�;��;�j�;[�;�[�;,n�;;��;���;��;�t�;E�;=x�;N�;Zۤ;���;k��;��;�،;�;q{�;@�w;�m;d}b;�X;<�M;)�C;�&:;��0;b3';�;�;9;�;�P�:;��:��:���:C�:�Ϧ:w͗:��:h#u:��X:T<:\� :�{:��95��9{!V9���8���6�E��D������Ź�������s�+�g�C��{[��s��@��P鐺+������������tʺ��պ�<���\�������@�3��,~���Y��UA#���(�_.���3�t9�0�>�݄D��J��O��U�ߨZ�j4`�}�e�)Ok�#�p��mv���{��ƀ������U��E��1䋻�����q���8�������Ǚ��  �  ��=P5=��=[�=�(=~�=;t=�=�� =d =� =+[�<8��<���<75�<2}�<���<��<�R�<���<���<�"�<`f�<7��<��<�+�<�k�<V��<���<[$�<�_�<���<���<d
�<�@�<v�<���<���<x�<9;�<�g�<��<���<s��<v�<t#�<x@�<-Z�<�p�<<��<H��<���<���<���<|��<���<0��<ۆ�<Ur�<�X�<!9�<��<���<%��<.�<�@�<I��<5��<&\�<�<=��<�9�<���<�U�<���<�W�<4��<�@�<׫�<k�<1q�<�˸<c �<p�<���<I �<,A�<q}�<m��<C�<)�<HE�<n�<���<-��<�՟<J�<D�<'�<>�<S�<Wf�<x�<+��<�<S��<_��<@��<ņ<�̈́<�Ղ<�܀<b�}<��y<��u<��q<��m<��i<q
f<~b<�#^<�1Z<�@V<_QR<�bN<vJ<��F<"�B<�><��:<��6<�3<�-/<7Q+</x'<��#<��<�<�:<Dw<��<~ <�M	<ġ<)�<���;��;2l�;�[�;:\�;n�;ڑ�;.��;�;�r�;�;�u�;��;2ؤ;���;���;Э�;֌;x�;�x�;X�w;�m;%zb;�X;L�M;�C;�':;ӕ0;�6';�;�;�>;��;�\�:���:���:7��:I%�:ۦ:�ؗ:��:a2u:[�X:��<:�� :؀:��9l��94V9U��8�x�6{ɾ�;oD��@��n�ŹC�������+�n�C��[��(s��J�������'����������tʺ��պX8���캣���D��K;�t��Fx�����3;#�1�(�HY.���3�o9���>�+�D��	J���O��U�b�Z�l5`��e�Sk���p�=rv�|��ɀ�����[Y��E ���狻����t��e;��/��ʙ��  �  c�=;5=��=P�=�(=��=Vt=�=1� =Jd =5	 =�[�<��<���<�5�<�}�<z��<��<%S�<��<^��<�"�<�f�<V��</��<�+�<�k�<)��<���<�#�<_�<*��<��<�	�<+@�<Hu�<	��<<��<��<�:�<|g�<%��<z��<J��<A�<x#�<�@�<SZ�<�p�<���<���<��<Y��<^��<7��<`��<��<���<�r�<+Y�<�9�<T�<���<a��<N�<�@�<N��<���<�[�<��<ݠ�<	9�<U��<U�<1��<�V�<b��<�?�<��<��<�p�<�ʸ<��<�o�<O��< �<�@�<�}�<���<e�<b�<�E�<�n�<%��<Ѷ�<�֟<��<��<�'�<�>�<�S�<�f�<�x�<���<E��<���<���<`��<�Ć<�̈́<sՂ<r܀<��}<p�y<��u<}�q<8�m<V�i<�f<b<$"^<_0Z<�?V<5PR<+bN<zuJ<T�F<��B<Ÿ><��:<��6<S3<E./<'R+<,y'<ϣ#<F�<<v<<�x<��<�<VO	<��<6�<���;R��;m�;�\�;�\�;�m�;:��;���;�;�q�;��;�s�;�;�դ;�;���;F��;=ӌ;&�;�v�;��w;�m;�xb;�X;��M;U�C;�(:;3�0;�8';�;�;�B;�;g�:���:9��:���:l1�:��:��:B"�:�Au:��X:�<:z� :s�:V	�9F��9 �U9I�8��6]?��A�D��f����Ź���T��K�+���C���[�%;s��T��l���z���I��v���a	�� sʺ��պ�5�Ќ�����p��7�4���r���~��<5#���(�T.���3�'k9���>��~D�J�}�O��U���Z�7`�S�e�Uk���p��vv��|�3̀�{���\��}#��Eꋻ����9w���=��u���˙��  �  <�=5=��=L�=�(=��=wt=�=g� ={d =g	 =H\�<Z��<+��<s6�<}~�<���<	�<�S�<���<���<"#�<�f�<h��<)��<�+�<ik�<��<K��<�#�<�^�<���<���<=	�<�?�<�t�<���<���<r�<5:�<g�<ґ�<-��<��<2�<t#�<�@�<�Z�<q�<��<4��<^��<���<ը�<���<��<n��<��<ms�<�Y�<�9�<��<C��<���<��<�@�<B��<��<�[�<��<���<�8�<���<�T�<���<vV�<���<.?�<���<�< p�<kʸ<{�<Jo�<��<���<�@�<q}�<���<��<��<F�<�n�<|��<9��<ן<���<��<d(�<+?�<#T�<Zg�<�x�<��<���<Ѥ�<���<[��<�Ć<�̈́<4Ղ<"܀<��}<��y<��u<��q<3�m<j�i<�f<"b<#!^<l/Z<�>V<UOR<saN<�tJ<щF<h�B<��><��:<*�6<�3<�./< S+<�y'<��#<7�<�<�=<�y<��<�<AP	<��<�<Z��;}��;@n�;]�;�\�;�m�;���;���;��;!p�;>�;r�;<�;�Ӥ;	��;c��;���;Jь;��;u�;k�w;�m;Fvb;�X;��M;^�C;�(:;ޘ0;�:';;D;�E;@�;�n�:���:��:���:�8�:3�:�:�'�:6Pu:�X:�<:�� :D�:��9���9��U9P �8��6���	�D�g���zƹ*.������,���C��[��Gs�M[�������������z����	���sʺ*�պ�1ẵ��������%4����Ro���!���0#���(�PP.���3�3h9�r�>��|D�J�K�O�U��Z�8`�T�e��Wk�I�p�zv�|��̀�����]���%��+싻����y��a?��+��͙��  �  ,�=
5=��=I�=�(=��=�t==o� =�d =�	 =�\�<���<x��<�6�<�~�<T��<g�<�S�<���<���<N#�<�f�<���<"��<�+�<]k�<ɩ�<$��<X#�<v^�<d��<1��<��<F?�<jt�<(��<d��<�<�9�<�f�<���<��<���<4�<f#�<�@�<�Z�<#q�<��<H��<���<��<?��<���<C��<ʗ�<Y��<�s�<�Y�<M:�<��<_��<���<��<�@�<0��<��<�[�<j�<L��<X8�<���<;T�<H��<�U�<t��<�>�<'��<��<�o�<1ʸ<=�<o�<๳<���<�@�<`}�<���<��<��<F�<o�<Ք�<���<~ן<���<��<�(�<�?�<�T�<�g�<6y�<'��<���<뤌<���<e��<�Ć<�̈́<Ղ<܀<��}<4�y<&�u<��q<y�m<��i<f<Ob<[ ^<�.Z< >V<�NR<�`N<�tJ<��F<\�B<��><��:<L�6<3<%//<!S+<{z'<L�#<�<�<7><�z<Q�<�<Q	<{�<��<���;@��;�n�;�]�;�\�;�m�;���;]��;_�;To�;��;�p�;��;8Ҥ;���;A��;�;
Ќ;*�;t�;��w;m;�ub;X;��M;�C;�):;{�0;�;';>;�;gH;�;yu�:'��:ö�:���:�=�:��:{�:�-�:�Su:��X:C�<:�� :]�:��9��9��U9���8���6�⿸�E����2/ƹ�J����e,��D���[�Ts��^��t��h���C������
��Xtʺ��պ�0��캒������G1����l�D�!��c.#�
�(� M.�4�3��e9���>�9{D�RJ���O��U�7�Z�8`�T�e�~Xk�$�p��{v��|�gπ�𗃻�_���&���틻~����z���@������͙��  �  )�=5=��=F�=�(=��=t=2=� =�d =�	 =�\�<ͥ�<���<�6�<�~�<j��<d�<�S�<Й�<��<|#�<�f�<���<0��<�+�<Hk�<���<��<;#�<`^�<E��<6��<��<+?�<[t�<��<g��<�
�<�9�<�f�<{��<	��<���<%�<e#�<�@�<�Z�<7q�<C��<b��<՞�<��<C��<	��<X��<��<h��<�s�<�Y�<l:�<��<���<Է�<y�<�@�<2��<׮�<w[�<[�<,��<<8�<���<T�<P��<�U�<`��<�>�<��<��<�o�<ʸ< �<o�<ѹ�<���<�@�<h}�<���<��<��<JF�</o�<唣<���<�ן<���< �<�(�<�?�<�T�<�g�<Wy�<E��<�<奈<���<|��<�Ć<v̈́<Ղ< ܀<G�}<�y<��u<��q<q�m<F�i<�f<b<L ^<�.Z<�=V<�NR<�`N<�tJ<g�F<;�B<��><�:<K�6<�3<�//<eS+<�z'<R�#<�<�<X><�z<z�<�<Q	<��<��<s��;��;an�;�]�;]�;�m�;K��;+��;8�;�n�;<�;6p�;�;�Ѥ;(��;
��;f��;Ќ;��;�s�;�w;�m;Hub;qX;C�M;�C;�*:;�0;�<';?;�;zI;֪;�u�:��: ��:��:�>�:���:?�:~/�:�Vu:z�X:��<:E� :��:F�9s��9w�U9���8��6����E�d����,ƹ�R��F��M,��	D�G�[�Xs�`����������󙳺���sʺl�պ�1ẝ��~������0���ck������-#���(�3M.�?�3��d9��>�QyD�2J��O�U�U�Z��8`���e��Xk��p�4|v��|��π�����&`��&'��L�����z��9A��5��{Ι��  �  ,�=
5=��=I�=�(=��=�t==o� =�d =�	 =�\�<���<x��<�6�<�~�<T��<g�<�S�<���<���<N#�<�f�<���<"��<�+�<]k�<ɩ�<$��<X#�<v^�<d��<1��<��<F?�<jt�<(��<d��<�<�9�<�f�<���<��<���<4�<f#�<�@�<�Z�<#q�<��<H��<���<��<?��<���<C��<ʗ�<Y��<�s�<�Y�<M:�<��<_��<���<��<�@�<0��<��<�[�<j�<L��<X8�<���<;T�<H��<�U�<t��<�>�<'��<��<�o�<1ʸ<=�<o�<๳<���<�@�<`}�<���<��<��<F�<o�<Ք�<���<~ן<���<��<�(�<�?�<�T�<�g�<6y�<'��<���<뤌<���<e��<�Ć<�̈́<Ղ<܀<��}<4�y<&�u<��q<y�m<��i<f<Ob<[ ^<�.Z< >V<�NR<�`N<�tJ<��F<\�B<��><��:<L�6<3<&//<!S+<{z'<L�#<�<�<7><�z<Q�<�<Q	<{�<��<���;@��;�n�;�]�;�\�;�m�;���;]��;_�;So�;��;�p�;��;8Ҥ;���;A��;�;	Ќ;*�;t�;��w;m;�ub;X;��M;�C;�):;{�0;�;';>;�;gH;�;yu�:'��:ö�:���:�=�:��:{�:�-�:�Su:��X:C�<:�� :]�:��9��9��U9���8���6�⿸�E����2/ƹ�J����e,��D���[�Ts��^��t��h���C������
��Xtʺ��պ�0��캒������G1����l�D�!��c.#�
�(� M.�4�3��e9���>�9{D�RJ���O��U�7�Z�8`�T�e�~Xk�$�p��{v��|�gπ�𗃻�_���&���틻~����z���@������͙��  �  <�=5=��=L�=�(=��=wt=�=g� ={d =g	 =H\�<Z��<+��<s6�<}~�<���<	�<�S�<���<���<"#�<�f�<h��<)��<�+�<ik�<��<K��<�#�<�^�<���<���<=	�<�?�<�t�<���<���<r�<5:�<g�<ґ�<-��<��<2�<t#�<�@�<�Z�<q�<��<4��<^��<���<ը�<���<��<n��<��<ms�<�Y�<�9�<��<C��<���<��<�@�<B��<��<�[�<��<���<�8�<���<�T�<���<vV�<���<.?�<���<�< p�<kʸ<{�<Jo�<��<���<�@�<q}�<���<��<��<F�<�n�<|��<9��<ן<���<��<d(�<+?�<#T�<Zg�<�x�<��<���<Ѥ�<���<[��<�Ć<�̈́<4Ղ<"܀<��}<��y<��u<��q<3�m<j�i<�f<"b<#!^<l/Z<�>V<UOR<saN<�tJ<щF<h�B<��><��:<*�6<�3<�./< S+<�y'<��#<7�<�<�=<�y<��<�<AP	<��<�<Z��;}��;@n�;]�;�\�;�m�;���;���;��;!p�;>�;r�;<�;�Ӥ;	��;c��;���;Jь;��;u�;k�w;�m;Fvb;�X;��M;^�C;�(:;ޘ0;�:';;D;�E;@�;�n�:���:��:���:�8�:3�:�:�'�:6Pu:�X:�<:�� :D�:��9���9��U9P �8��6���	�D�g���zƹ*.������,���C��[��Gs�M[�������������z����	���sʺ*�պ�1ẵ��������%4����Ro���!���0#���(�PP.���3�3h9�r�>��|D�J�K�O�U��Z�8`�T�e��Wk�I�p�zv�|��̀�����]���%��+싻����y��a?��+��͙��  �  c�=;5=��=P�=�(=��=Vt=�=1� =Jd =5	 =�[�<��<���<�5�<�}�<z��<��<%S�<��<^��<�"�<�f�<V��</��<�+�<�k�<)��<���<�#�<_�<*��<��<�	�<+@�<Hu�<	��<<��<��<�:�<|g�<%��<z��<J��<A�<x#�<�@�<SZ�<�p�<���<���<��<Y��<^��<7��<`��<��<���<�r�<+Y�<�9�<T�<���<a��<N�<�@�<N��<���<�[�<��<ݠ�<	9�<U��<U�<1��<�V�<b��<�?�<��<��<�p�<�ʸ<��<�o�<O��< �<�@�<�}�<���<e�<b�<�E�<�n�<%��<Ѷ�<�֟<��<��<�'�<�>�<�S�<�f�<�x�<���<E��<���<���<`��<�Ć<�̈́<sՂ<r܀<��}<p�y<��u<}�q<8�m<V�i<�f<b<$"^<_0Z<�?V<5PR<+bN<zuJ<T�F<��B<Ÿ><��:<��6<S3<E./<'R+<,y'<ϣ#<F�<<w<<�x<��<�<UO	<��<6�<���;R��;m�;�\�;�\�;�m�;:��;���;�;�q�;��;�s�;�;�դ;�;���;F��;=ӌ;&�;�v�;��w;�m;�xb;�X;��M;U�C;�(:;3�0;�8';�;�;�B;�;g�:���:9��:���:l1�:��:��:B"�:�Au:��X:�<:z� :s�:V	�9F��9 �U9I�8��6]?��A�D��f����Ź���T��K�+���C���[�%;s��T��l���z���I��v���a	�� sʺ��պ�5�Ќ�����p��7�4���r���~��<5#���(�T.���3�'k9���>��~D�J�}�O��U���Z�7`�S�e�Uk���p��vv��|�3̀�{���\��}#��Eꋻ����9w���=��u���˙��  �  ��=P5=��=[�=�(=~�=;t=�=�� =d =� =+[�<8��<���<75�<2}�<���<��<�R�<���<���<�"�<`f�<7��<��<�+�<�k�<V��<���<[$�<�_�<���<���<d
�<�@�<v�<���<���<x�<9;�<�g�<��<���<s��<v�<t#�<x@�<-Z�<�p�<<��<H��<���<���<���<|��<���<0��<ۆ�<Ur�<�X�<!9�<��<���<%��<.�<�@�<I��<5��<&\�<�<=��<�9�<���<�U�<���<�W�<4��<�@�<׫�<k�<1q�<�˸<c �<p�<���<I �<,A�<q}�<m��<C�<)�<HE�<n�<���<-��<�՟<J�<D�<'�<>�<S�<Wf�<x�<+��<�<S��<_��<@��<ņ<�̈́<�Ղ<�܀<b�}<��y<��u<��q<��m<��i<p
f<~b<�#^<�1Z<�@V<_QR<�bN<vJ<��F<"�B<�><��:<��6<�3<�-/<7Q+</x'<��#<��<�<�:<Dw<��<~ <�M	<ġ<)�<���;��;1l�;�[�;:\�;n�;ڑ�;-��;�;�r�;�;�u�;��;2ؤ;���;���;Э�;֌;x�;�x�;X�w;�m;%zb;�X;K�M;�C;�':;ӕ0;�6';�;�;�>;��;�\�:���:���:7��:I%�:ۦ:�ؗ:��:a2u:[�X:��<:�� :؀:��9l��94V9U��8�x�6{ɾ�;oD��@��n�ŹC�������+�n�C��[��(s��J�������'����������tʺ��պX8���캣���D��K;�t��Fx�����3;#�1�(�HY.���3�o9���>�+�D��	J���O��U�b�Z�l5`��e�Sk���p�=rv�|��ɀ�����[Y��E ���狻����t��e;��/��ʙ��  �  ǎ=|5=
�=d�=�(=g�=t=}=�� =�c =� =qZ�<l��<��<p4�<q|�<��<8�<�Q�<��<���<*"�<f�<��<��<,�<�k�<���<o��<�$�<H`�<l��<j��<:�<�A�<�v�<���<���<+�<�;�<�h�<	��<&��<���<��<�#�<U@�<�Y�<"p�<͂�<ב�<ۜ�<���<��<���<��<j��<��<�q�<�W�<v8�<p�<3��<¶�<�~�<�@�<Z��<c��<f\�<��<ҡ�<:�<���<yV�<���<�X�<
��<_A�<���<+�<�q�<7̸<� �<�p�< ��<~ �<TA�<{}�<M��<�<��<�D�<�m�<�<{��<F՟<��<�<[&�<9=�<IR�<�e�<iw�<���<y��<���<,��<(��<ņ<�̈́<�Ղ<.݀<��}<��y<!�u</�q<<�m<l j<�f<0b<6%^<3Z<9BV<�RR<dN<wJ<f�F<g�B<�><��:<L�6<@3<�,/<WP+<�v'<-�#<n�< <Q9<�u<j�<��<kL	<K�<��<߸�;��;�j�;[�;�[�;,n�;;��;���;��;�t�;E�;=x�;N�;Zۤ;���;k��;��;�،;�;q{�;@�w;�m;d}b;�X;;�M;)�C;�&:;��0;b3';�;�;9;�;�P�:;��:��:���:C�:�Ϧ:w͗:��:h#u:��X:T<:\� :�{:��95��9{!V9���8���6�E��D������Ź�������s�+�g�C��{[��s��@��P鐺+������������tʺ��պ�<���\�������@�3��,~���Y��UA#���(�_.���3�t9�0�>�݄D��J��O��U�ߨZ�j4`�}�e�)Ok�#�p��mv���{��ƀ������U��E��1䋻�����q���8�������Ǚ��  �  ��=�5=!�=l�=|(=N�=�s=G=t� =fc =; =�Y�<���<<��<�3�<�{�<.��<y
�<=Q�<]��<���<�!�<�e�<��<��<$,�<,l�<��<���<z%�<�`�<?��<=��<�<�B�<�w�<u��<���<�<�<�<i�<���<���<��<��<�#�<A@�<�Y�<�o�<T��<.��<7��<R��<0��<ڤ�<��<���<?��<�p�<(W�<�7�<��<���<x��<�~�<s@�<o��<���<�\�<�<W��<�:�<n��<cW�<���<�Y�<���<SB�<���<�<�r�<�̸<�!�<q�<s��<� �<uA�<�}�<8��<��<j�<gD�<�l�<S��<Ĵ�<lԟ<��<��<{%�<`<�<|Q�<�d�<�v�<��<��<���<���<��<ņ<΄<Gւ<�݀<��}<��y<��u<��q<��m<=j<�f<b<�&^<�4Z<�CV<�SR<7eN<�wJ<)�F<ȡB<C�><��:<��6<�3<�+/<)O+<�u'<џ#<��<> <�7<�s<��<�<�J	<�<v�<{��;T��;�i�;BZ�;�[�;Cn�;��;���;^�;w�;��;S{�;h �;zޤ;��;���;w��;�ی;_�;~�;��w;3m;+�b;X;��M;I�C;�%:;��0;�0';� ;l;�3;Z�;0C�:���:u��:���:�
�:���:K:m�:3u:��X:�t<:�� :�x:G
�9Rǟ9gKV9�P�8�q�6&����C��ܓ�YgŹ�x��V����+���C�3a[��r��6���ߐ�tz��|��v�������tʺ��պ�@���������#F���!�������cH#�k�(��e.���3�ry9�
?�_�D�J���O�U�c�Z�,3`���e�'Lk��p�iv���{�wÀ�;���aR�������������zn���5�������ř��  �  -�=�5=:�=p�=s(=5�=�s==/� =c =� =�X�<���<V��<�2�<�z�<[��<�	�<}P�<Ŗ�<u��<d!�<|e�<���<���<5,�<bl�<f��<I��<&�<�a�<��<��<��<wC�<�x�<K��<g��<��<<=�<�i�<��<��<J��<��<�#�<.@�<sY�<qo�<��<���<���<~��<]��<��<%��<���<j��<�o�<RV�<47�<1�<M��<��<~~�<f@�<p��<���<]�<e�<��<�;�<"��<&X�<���<gZ�<���<FC�<���<��<�s�<�͸<W"�<�q�<ϻ�<�<�A�<�}�<&��<��<�<�C�<Vl�<���<ﳡ<�ӟ<��<��<�$�<�;�<�P�<%d�<v�<���<���<H��<���<��< ņ<E΄<�ւ<�݀<��}<3�y<��u<h�q<��m<�j<�f<�b<�(^<i6Z<1EV<)UR<ffN<�xJ<��F<3�B<Z�><r�:<��6<�
3<+/<N+<Mt'<.�#<�<��<�5<�q<ų<Y�<I	<K�<-�<A��;���;�g�;uY�;5[�;Nn�;���;���;��;Zy�;�;�}�;y#�;��;m��;#��;���;Cߌ;"�;���;��w;!m;͂b;�X;��M;��C;�$:;]�0;l-';b�;z�;~.;��;�5�:+��:'s�:��:��:9��:���:���:��t:�zX:Yh<:� :�u:��9I͟9�jV9���8}�6����rC�
���W0Ź�B��rt���+��C�]F[�6�r�:,��gՐ��r������������yuʺv�պ"F�������צ��K����ԋ��%�����O#��(�$l.�n�3�s~9��?���D�J���O��U�8�Z��1`���e��Hk���p��cv�V�{�s���ȇ���N����(݋�B���ek���2������qÙ��  �  h�=�5=P�=w�=i(=%�=�s=�=� =�b =~ = X�<��<���<�1�<�y�<���<��<�O�<;��<���<� �<.e�<���<���<O,�<�l�<ë�<���<�&�<9b�<���<���<��<=D�<cy�<��<!��<x�<�=�<Sj�<x��<V��<���<�<�#�<@�<JY�<o�<b��<��<��<͡�<���<.��<]��<��<���<Mo�<�U�<�6�<��<���<���<V~�<M@�<t��<߯�<W]�<��<^��<<�<���<�X�<P��<A[�<���<D�<k��<��<Yt�<Zθ<�"�<r�<=��<]�<�A�<�}�<��<K�<��<lC�<�k�< ��<A��<�ҟ<��<�
�<�#�<�:�<�O�<vc�<�u�<���<��<䢌<���<꺈<'ņ<p΄<�ւ<gހ<}�}<^�y<^�u<��q<1�m<j<)f<Pb<<*^<�7Z<�FV<iVR<IgN<�yJ<d�F<��B<y�><O�:<G�6<>
3<*/<�L+<'s'<˜#<��<��<�3<_p<�<��<�G	<��<�<ձ�;���;�f�;�X�;�Z�;�n�;/��;��;��;�z�;l�;r��;3&�;��;X��;��;���;�;�$�;2��;��w;/$m;�b;�X;��M;��C;�#:;ݍ0;*';�;'�;H);Շ;V*�:G��:Lf�:V��:�:��:*��:4�:�t:�iX:[<:� :zq:?�9�ן9�V9��8�E�6�}��dC������ŹE��C[��z+��iC�l/[�m�r��!��Hΐ��k����������� ��Fvʺ��պrJ�@�캃��
��&Q��������,����V#���(��q.���3�"�9�
?���D�J���O�K U���Z�l0`�+�e�OEk�/�p��^v���{����������K����ڋ����h��!0��`��������  �  ��=6=`�=��=](=	�={s=�=�� =�b =4 =yW�<;��<���<1�<+y�<���<K�<7O�<���<���<� �<e�<h��<���<m,�<�l�<��<��<'�<�b�<@��<o��<l�<�D�<z�<ԭ�<���< �<w>�<�j�<��<���<���<"�<�#�<�?�<Y�<�n�<��<���<V��<;��<���<��<���<(��<��<�n�<U�<�5�<F�<��<���<2~�<%@�<���<��<�]�<*�<̣�<�<�<q��<�Y�<��<\�<���<�D�<3��<p�<u�<�θ<^#�<}r�<���<��<�A�<�}�<ߴ�<+�<u�<C�<Yk�<j��<���<,ҟ<T�<6
�<#�<:�<HO�<�b�<�t�<���<͔�<���<[��<ʺ�<@ņ<�΄<ׂ<�ހ<^�}<W�y<��u<1�q<��m<j<�f<�b<�+^<=9Z<�GV<gWR<9hN<KzJ<ӍF<٢B<��>< �:<��6<�	3<�)/< L+<�q'<��#<U�<o�<�2<�n<��<:�<<F	<��<��<8��;\��;�e�;�W�;�Z�;�n�;���;���;��;�|�;7��;ɂ�;�(�;k�;!��;ɰ�;{��;��;Q'�;+��;l�w;A'm;�b;�X;u�M;B�C;E":;M�0;C(';`�;��;E$;�;��:��:MZ�:w�:��:v��:П�:Z�:��t:#_X:�S<:�� :vk:�
�98ߟ9A�V9�U�8�y�6���-�B�	X����Ĺ����wD�uc+�YRC��[�Ͷr�����Ɛ�=f������H�������7vʺ"�պ M���'
��/���U�r�����2�����[#�K�(�$w.�p 4���9�9?� �D��J�c�O�A!U�#�Z�}/`���e�1Ck���p�[v�:�{�캀������H��?��׋�Z����e���-��t���꿙��  �  ��=16=p�=��=X(=��=[s=�=�� =Ob =� = W�<���<V��<�0�<�x�<]��<��<�N�<C��<3��<] �<�d�<N��<���<f,�<�l�<@��<W��<t'�<c�<���<���<��<�E�<�z�<S��<@��<��<�>�<:k�<>��<ټ�<���<*�<�#�<�?�<�X�<�n�<���<=��<��<נ�<u��<��<��<���<x��<n�<�T�<�5�<��<0��<D��< ~�<!@�<���<��<�]�<q�<*��<
=�<���<Z�<���<�\�<��<vE�<���<��<yu�<Kϸ<�#�<�r�<Ѽ�<��<�A�<�}�<մ�<��<,�<�B�<�j�<��<A��<�џ<��<�	�<�"�<�9�<�N�<yb�<|t�<3��<z��<v��<2��<���<:ņ<�΄<Cׂ<�ހ<*�}<!�y<F�u<�q<u�m<!j<�f<�b<�,^<(:Z<�HV<3XR<iN<�zJ<]�F<�B<��><�:<��6<k	3<�(/<hK+<q'<Ě#<\�<m�<�1<�m<��<+�<SE	<��<��<���;���;�d�;-W�;KZ�;�n�;��;���;��;F~�;���;<��;d*�;�;,��;ܲ�;[��;?�;�(�;|��;� x;�)m;ǉb;� X;��M;��C;�!:;��0;�%';��;B�;� ;�;L�:��:�Q�:Hn�:ݵ:ٔ�:X��:�ވ:"�t:�TX:�J<:�� :$j:��9Fߟ9�V9���8���6����U�B�;>���Ĺ�����2�CR+�+DC��[�S�r����a����a������]~��C���qvʺ;�պ�P���n�����<Y��������5�����_#���(�{.��4�\�9�2?���D�zJ���O��!U�C�Z��.`���e�Ak�x�p��Wv�>�{�-���2����F�����ԋ�����d��;,������B����  �  ď=;6=y�=��=V(=��=Js=x=i� =8b =� =�V�<Z��<���<?0�<Jx�<��<�<�N�<��<���<A �<�d�<M��<���<r,�<�l�<Z��<���<�'�<bc�<���<N��<;�<�E�<{�<���<���<��<.?�<ak�<W��<��<��<B�<�#�<�?�<�X�<yn�<���<��<���<u��<"��<���<ƛ�<N��<��<�m�<NT�<[5�<��<��<0��<�}�<%@�<���<+��<�]�<��<L��<.=�<4��<mZ�<���<�\�<���<�E�<��<b�<�u�<�ϸ<�#�<�r�<���<��<B�<�}�<۴�<��<�<�B�<�j�<���<㱡<Xџ<w�<Z	�<3"�<%9�<rN�<b�<Kt�<���<T��<T��<'��<���<5ņ<�΄<Rׂ<߀<O�}<��y<��u<��q<B�m<�j<mf<� b<R-^<�:Z<KIV<�XR<7iN<4{J<��F<C�B<��><�:<��6<'	3<�(/<�J+<�p'<�#<��<��<�0<�l<®<p�<�D	<�<��<���;x��;d�;W�;Z�;�n�;K��;��;4�;u~�;���;x��;�+�;t�;j;E��;w��;��;=*�;߇�;�x;�*m;�b;� X;8�M;a�C;�!:;�0;%';3�;l�; ;�|;��:΂�:>L�: i�:�յ:���:��:�ڈ:�t:�NX:�G<:s� :7j:�9{�9��V9���8�R 7Su���|B�^(���Ĺd���&'��F+�&9C�|�Z�ʟr����?���b_����G}�����Ewʺ�պ�Rẅ�����)���[����I��9�����b#�U�(��}.��4��9�?���D��J��O��!U�h�Z�.`��e��?k���p�;Vv���{������~���E������Ӌ�
����b���*���� ����  �  }�=[9=�=��=�,=��=Ux=�=&� =Yh =U =�d�<:��<���<OA�<���<���<��<oe�<���<R��<}<�<���<2��<��<7P�<���<���<��<�R�<���<��<j�<�B�<W{�<ز�<���<`�<P�<��<��<���<�<�.�<�S�<�u�<��<���<���<���<���<��<q�<�
�<�<��<�<���<	��<��<���<]��<�d�<6�<� �<;��<Ӏ�<[6�<~��<m��<+�<l��<�T�<���<b�<t��<4T�<�ÿ<�,�<r��<O�<�C�<���<�<�'�<Si�<��<�ݮ<�<�@�<l�<���<<�أ<-��<��<,�<gC�<�X�<@l�<=~�<���<���<B��<���<�<s̊<Ո<�܆<�<��<H�<h�}<E�y<(�u<��q<��m<��i<�f<_
b<^<JZ<� V<"*R<z4N<C@J<MF<~[B<Kk><�|:<,�6<��2<�.<��*<v�&<S#<�?<Bj<�<�<�	<�J<�<�<�4<�!�;���;k��;դ�;���;��;���;X��;-�;n��;��;^t�;�;!Ǣ;���;���;ه�;��;6�;^�~;Svs;��h;�];j�S;hI;An?;�5;,;S�";��;�;c�;ܩ�:���:��:�v�:X½:y`�:�O�:���: �:��g:f�K:��/:�:���9�۾9~��9%�-9�[�8E������e�=B���չ��p��#�2�I0J��a��y����e����'��ܝ��.
���m���̺�&غ�{㺓��8����RH����"x�N
�Ζ��$��)��$/���4�N:�l�?��E�ЈJ��P�|U��Z��u`�b�e��wk���p�t�v��|��ƀ�׉���M�����ԋ�*����\��� ���喻����  �  i�=U9=�=z�=�,=��=hx=�=8� =dh =d =�d�<[��<���<cA�<�<���<��<�e�<̭�<s��<�<�<ڂ�<K��<��<#P�<���<���<��<�R�<p��<���<T�<iB�<:{�<���<���<?�<P�<��<��<���<�<�.�<�S�<�u�<��<���<���<���<���<-��<��<�
�<.�<��<<�<���<��<;��<ï�<s��<�d�<"6�<� �<F��<Ԁ�<F6�<|��<Z��<�*�<S��<�T�<���<�a�<F��<T�<cÿ<k,�<X��<K�<iC�<䔷<��<�'�<Oi�< ��<�ݮ<��<�@�<.l�<���<���<
٣<L��<��<J,�<C�<�X�<bl�<R~�<���<ʝ�<h��<���<�<�̊< Ո<�܆<�<��<"�<<�}<�y<�u<t�q<��m<��i<.f<
b<�^<*Z<� V<�)R<O4N<�?J<�LF<U[B<-k><�|:<b�6<�2<=�.<8�*<��&<�#<�?<�j<<�<H�<'
<K<V�<5�<#5<"�;��;(��;D��;���;���;��;-��;�,�;;��;"�;Vt�;��;aƢ;=��;��;H��;���;@�;��~;�us;��h;X�];b�S;\gI;*n?;2�5;�,;�";��;�;B�;]��:���:���:�x�:�Ľ:Kc�:�P�:4��:��:��g:��K:*�/:��:��9�ܾ9���9g�-9�K�8��*����e�A���չ]�������2�m6J�	�a��y���V����)������J
��,o����̺Z%غ7y�p�� ������G�����w������$��)��#/���4�~:�9�?��E���J�P��{U�|�Z��v`���e�yk�m�p�X�v�$|��ƀ�����#N�����KՋ������\�� !��<斻U����  �  M�=I9=��=~�=�,=��=zx==b� =�h =� =e�<Ѯ�<s��<�A�<I��<]��<[�<�e�<��<���<�<�<���<Q��<��< P�<g��<���<��<yR�<��<���<��<�A�<�z�<9��<M��<��<�O�<���<���<t��<��<�.�<�S�<�u�<���<���<��<���<'��<���<	�<b�<��<o	�<��<7��<���<���<��<���<:e�<F6�<� �<G��<���</6�<Z��<(��<�*�<��<T�<B��<^a�<���<�S�<�¿<�+�<؎�<��<�B�<���<��<}'�<-i�<�<ޮ<��<�@�<Kl�<��<J��<m٣<���<[�<�,�<�C�<NY�<�l�<�~�<0��<��<���<뷎<�<�̊<+Ո<�܆<��<m�<��<��}<U�y<:�u<��q<��m<��i<.f<?	b<�^<MZ<�V<)R<�3N<?J<�LF<"[B<;k><�|:<u�6<I�2<��.<��*<I�&<v#<�@<xk<J�<-�<?<�K<J�<�<�5<l#�;���;���;w��; ��;���;���;���;�+�;v��;��;�r�;�;Ģ;���;-�;���;���;��;f�~;Uss;�h; �];��S;�fI;�n?;t�5;�,;r�";��;��;��;���:���:Ό�:U��:�˽:�k�:JW�:���:5�:��g:�K:&�/:7�:`��9��9���9�-9 �8��򷘸��6f�^[��4չ��������2��EJ��a�:y�%������-��𠪺����o����̺%غ�w�W��G�����D����5t�������$�6�)�o /��4��:���?�pE���J�� P��{U��Z�Bw`�h�e��zk��p�2�v�p
|��Ȁ�|����O������֋�󚎻x^���"���疻)����  �  $�=#9=��=y�=�,=��=�x=8=�� =�h =� =�e�<y��<"��<�B�<��<��<��<�f�<���<0��<=�<<��<{��<��<P�<)��<J��<+�<�Q�<���< ��<;�<GA�<z�<���<���<�<O�<��<#��<��<��<v.�<�S�<�u�<��<���<r��<\��<���<��<��<�<P�<-
�<n�<���<0��<:��<���<4��<�e�<�6�<� �<Z��<р�<6�<��<Ҋ�<>*�<~��<�S�<���<�`�<��<�R�<$¿<5+�<$��<4�<nB�<��<7�<&'�<�h�<ץ�<ޮ<��<,A�<�l�<l��<���<�٣<T��<�<u-�<�D�<Z�<�m�<h�<Ï�<���<,��<[��<9Ì<�̊<=Ո<�܆<��<#�<��<��}<]�y<�u<X�q<J�m<t�i<�f<�b<h^<Z<�V<(R<�2N<�>J<'LF<�ZB<#k><�|:<Ԑ6<�2<m�.<��*<Z�&<�#<�A<�l<��<��<�<eM<��<T�<�6<F%�;���;���;J��;F��;���;Լ�;���;o*�;���;��;�p�;��;¢;ؑ�;}|�;��;T��;Y�;�~;�os;Șh;��];��S;2fI;�n?;Q�5;�,;E�";�;��;��;��:���:*��:���:ؽ:�u�:�b�:���:q�:��g:<�K:��/:4�:F��9A߾9}�9�]-9Iԍ8 P�����tf�����A]չ�����9�2��ZJ���a��&y�},��9����3������$���p��a�̺�"غIs����-���?�#���n�r��X��$� �)�./�z�4��:�2�?��	E��J���O�"{U�_�Z��x`���e�}k��q��v��|�ˀ�
����R��m���ً�y����`��%���閻����  �  �=�8=��=o�=�,=��=�x=y=�� =.i =I =�f�<o��<
��<�C�<Ռ�<��<��<Ig�<R��<���<�=�<���<���<��<�O�<���<���<��<XQ�<ގ�<,��<c�<Y@�<!y�<���<���<@�<,N�<O�<z��<{��<0�<2.�<�S�<�u�<8��<=��<���<���<;��<���<h�<��<6�<!�<d�<���< ��<��<m��<Ԏ�<#f�<�6�<)�<���<���<�5�<���<m��<�)�<���<�R�<���<�_�<��<�Q�<&��<3*�<<��<L�<�A�<`��<�ߵ<�&�<�h�<���<�ݮ<��<jA�<m�<�<k��<�ڣ<&��< �<S.�<�E�<�Z�<sn�<S��<���<k��<Ĭ�<㸎<�Ì<͊<XՈ<�܆<��<��<<�<��}<�y<��u<��q<��m<}�i< f<�b<�^<AZ<�V<�&R<�1N<�=J<{KF<nZB<�j><}:<P�6<��2<q�.<��*<��&<;#<�C<�n<��<��<{<nO<c�<��<k8<�'�;���;m��;k��;���;���;a��;���;�(�;V~�;U�;�m�;t	�;���;F��;!y�;]�;	��;�;�y~;�js;ߔh;J�];ĒS;�eI;�n?;ܭ5;!",;��";��;��;�;6��:�:��:%��:��:_��:�q�:��:-#�:�g:�K:�0:��:���9oݾ9)w�9�?-9�|�8P���L�n�f����!�չ��?���2��xJ���a��Ay��7��S���;��ݪ��,��r����̺Gغ�n�ܷ���������9�c���f�f��w���$�o�)��/�4�4��:�}�?��E�9�J���O�^zU���Z��y`�3�e�?�k�~q�H�v�C|��΀������V������݋����od��=(��Q얻~����  �  ��=�8=��=h�=�,=
�=�x=�==� =�i =� =�g�<}��<)��<�D�<���<��<��<*h�<��<o��<>�<��<���<��<�O�<���<��<!�<�P�<��<F��<h�<K?�<x�<���<���<7�<9M�<h~�<ĭ�<���<��<�-�<cS�<�u�<X��<���<Q��<���<���<���<U�<��<R�<0�<o�<���<��<���<8��<���<�f�<s7�<k�<���<���<�5�<c��<щ�<)�<��<�Q�<���<�^�<���<�P�< ��<)�<,��<P�<�@�<���<ߵ<1&�<Lh�<���<�ݮ<��<�A�<�m�<���<%��<�ۣ<��<��<p/�<�F�<\�<�o�<J��<{��<8��<|��<s��<Č<Z͊<yՈ<�܆<w�<t�<��<~�}<~�y<��u<��q<n�m<S�i<��e<�b<y
^<FZ<	V<%R<Z0N<�<J<�JF<�YB<�j><K}:<��6<_�2<��.<[�*<x�&<#<�E<�p<�<�<�<�Q<l�<��<:<�*�;���;"��;f��;0��;z��;���;��;�&�;�{�;#�;*j�;��;���;B��;�t�;C{�;��;~݄;�r~;ees;E�h;�];R�S;�dI;�n?;"�5;�$,;��";��;��;��;p��:��:��:{��:���:���:���:S��:[0�:��g:��K:0:g�:x��9�߾9vl�9�-9r�8������*Gg�]�����չ $�\&��2���J�Ob�_y��E���ʓ��D��粪�a���s��y�̺�غ<i㺢���������2�����^�X���{��$�؉)�/�ȋ4�;	:�Ѕ?�hE��}J���O�hyU�:�Z�5{`�S�e��k�qq���v�l|�dҀ������Z��{���ዻ1���Qh���+��������  �  X�=�8=��=Y�=�,=+�=:y= =�� = j =B =�h�<���<Z��<�E�<%��<��<� �<&i�<��<��<�>�<U��<��<��<�O�<p��<��<��<�O�<$��<T��<H�<+>�<�v�<K��<v��<�<:L�<�}�<��<+��<�<�-�<#S�<�u�<x��<ڱ�<���<��<���<���<e	�<�<q�<[�<��<���<��< ��<��<S��<Ig�<�7�<��<���<���<k5�<��<D��<C(�<!��<�P�<���<r]�<���<\O�<���<�'�<�<F�<�?�<đ�<J޵<�%�<�g�<=��<�ݮ<�<B�<�m�<.��<�<{ܣ<!��<�<�0�<�G�<8]�<�p�<[��<���<��<D��< ��<�Č<�͊<�Ո<p܆<4�<�<�<�}<��y<��u<��q<�m<�i<8�e<Rb<"^<Z<'V<J#R<�.N<�;J<�IF<[YB<�j><r}:<>�6<H�2<��.<��*<.�&<2!#<H<>s<\�<w�<L<�S<��<��<�;<�-�;>��; ��;���;���;��;���;���;�$�;'y�;��;�f�;��;[��;ą�;=p�;w�;Ù�;�ل;=l~;_s;�h;g�];�S;�bI;�n?;n�5;�',;��";`�;K�;;���:.,�:~��:���:��:Q��:咟:�ǐ:?�:F�g:I�K:�+0:��:���9߾9�]�9J�,9�r�8��4�H�g�4��uֹ�G�jM��3���J��3b��}y��S���ד�SO�����P��Vw����̺�غ�b㺪����ܐ�1+���FV�����r�#�#��)��/�g�4�c:��?��D�zJ���O��xU���Z�g}`�@f�k�k�Rq�r�v��#|��ր�P���b_��a#���拻˩���l��/��������  �  �=[8=r�=P�=�,=P�=my=M=�� =oj =� =�i�<���<���<	G�<I��<G��<�!�<j�<Ǳ�<���<&?�<���<]��<�<�O�<(��<���<��<!O�<F��<F��<7�<=�<�u�<#��<G��<�<'K�<�|�<��<���<��<-�<�R�<�u�<���<)��<8��<���<���<d �<Y
�<%�<��<��<��<��<=��<���<��<��<�g�<O8�<�<���<���<45�<���<���<�'�<;��<�O�<y��<L\�<v��<N�<q��<�&�<͉�<�<�>�<ᐷ<�ݵ<%%�<�g�<��<�ݮ<J�<XB�<qn�<֖�<���<Vݣ<��<%�<�1�<I�<b^�<�q�<x��<{��<���<��<���<�Č<�͊<�Ո<c܆<��<��<��<��}<�y<��u<c�q<��m<��i<��e<��a<�^<�Z<V<�!R<N-N<q:J<�HF<�XB<`j><�}:<Β6<�2<��.<b�*<��&<##<<J<�u<¥<��<�<<V<�<��<�=<�0�;���;���;��;G��;ܢ�;޹�; ��;�"�;Fv�;��;�b�;���; ��;1��;�k�;�r�;���;�Մ;e~;�Xs;[�h;��];�S;�aI;�n?;q�5;X*,;o�";�;��;
;���:�>�:���:G��:��:i��:K��:Zא:3M�:�	h:�K:x;0:��:}�9�޾9�S�9q�,9l��8�����w�w-h��x���bֹAm��r��C3���J��Ub�ݟy��a���䓺X��D���d!��Py����̺�غ@]�y��P�����$���M�����h���#��w)���.��{4�p�9�|y?�*�D��vJ�Y�O�5wU�d�Z�"`��f�{�k��q��v��+|��ڀ�����d���'��V닻*����p���3��[���幙��  �  Ӑ=(8=V�=A�=�,=m�=�y=�=M� =�j =+ =�j�<Ǵ�<���<.H�<\��<N��<�"�<�j�<���<w��<�?�<��<���<
�<zO�<��<*��<e�<kN�<z��<X��<@�<�;�<�t�<��<%��<�<0J�<�{�<W��<���<�<�,�<�R�<�u�<ϕ�<m��<���<U��<5��<C�<B�< �<��<��<��<��<;��<���<δ�<���<�h�<�8�<G�<���<���<5�<0��<*��<�&�<m��<�N�<s��<@[�<A��<�L�<I��<v%�<�<�<�=�<��< ݵ<�$�<0g�<ݤ�<�ݮ<j�<�B�<�n�<k��<n��<4ޣ<	��<(�<�2�<2J�<o_�<�r�<t��<`��<Т�<���<=��<dŌ<4Ί<�Ո<I܆<��<M�<�<<�}<��y<�u<r�q<��m<R�i<��e<��a<�^<�Z<7V<�R<�+N<[9J<HF<`XB<j><�}:<?�6<�2<��.<��*<�'<�$#<=L<�w<��<^�<�<eX<�<��<\?<�3�;I��;���;���;���;���;��;���;� �;�s�;�ݵ;5_�;���;��;}�;�g�;2n�;���;�ф;�^~;#Ss;j�h;�];ÈS;�`I;�n?;��5;�,,;��";	�;i�;K;�	�:�N�:���:���:=1�:�̮:���:k�:v[�:Dh:�K:�L0::�:��9�ܾ9gK�9��,9�x�8(< ���[�h�����:�ֹ{�����Bf3�+K��tb���y��n����a���Ȫ��%��E{���̺�غ�W�H��b���N����l���D�D���_�J�#�|o)���.��t4���9�Qt?�Y�D�'sJ�j�O��vU�E�Z���`��f���k��q�D�v��2|��ހ������h��A,���_����t��07�����������  �  ��=�7=7�=:�=-=�=�y=�=�� =.k =� =�k�<���<���<I�<T��</��<�#�<�k�<2��<��<@�<]��<���<�<]O�<���<���<��<�M�<���<���<S�<;�<�s�<��<C��<�<YI�<�z�<���<P��<��<�,�<�R�<�u�<��<���<��<���<���<��<�<��<��<��<��<��<��<���<���<c��<�h�<9�<x�<
��<���<�4�<���<���<I&�<���<N�<���<:Z�<M��<�K�<C��<y$�<�<@�<=�<j��<dܵ<($�<�f�<���<�ݮ<x�<�B�<Jo�<ꗧ<��<�ޣ<���<�<�3�<K�<a`�<�s�<L��<4��<���<R��<���<�Ō<_Ί<�Ո<G܆<��<��<��< �}<"�y<��u<��q<��m<��i<��e<��a<�^<
Z<�V<vR<�*N<U8J<]GF<�WB<�i><�}:<��6<��2<��.<��*<�'<�&#<�M<�y<�</�<�<=Z<��<q�<�@<6�;��;��;���;��;h��;L��;\��;��;�q�;�ڵ;A\�;f��;t��;~y�;d�;�j�;C��;�΄;�X~;�Ms;K}h;��];ՆS;`_I;o?;��5;�.,;��";�;��;1;c�:~\�:B��:���:�?�:ܮ:dß:
��:~g�:�4h:�L:�W0:�:�9r޾9�>�92u,9��8|U��*�Z�h��ꥹ��ֹ�����3��#K�Βb�O�y�{������fj��	Ϫ��)���}��S�̺	غS㺍�������������=�����X���#�h)��.�$n4�'�9�mo?���D��pJ�!�O��uU�h�Z���`�:f�k�k�� q��v��8|�7※����.l��20��l�9���Tx��B:��l��������  �  ^�=�7= �=5�=-=��=�y=�=�� =jk =� =7l�<P��<A �<�I�<��<���<W$�<Hl�<���<~��<i@�<���<���<#�<KO�<o��<|��<p�<aM�<)��<���<� �<`:�<�r�<M��<���<V�<�H�<_z�<)��<���<G�<<,�<sR�<�u�<���<��<Y��<-��<Y��<p�<��<��<.�<=�<w	�<���<���<K��<���<ޒ�<\i�<e9�<��<��<~��<�4�<���<J��<�%�<-��<{M�<���<zY�<���<K�<x��<�#�<��<��<w<�<鎷<�۵<�#�<�f�<���<�ݮ<��<#C�<�o�<W��<���<uߣ<y��<��<f4�<�K�<a�<[t�<<ϕ�<���<հ�<��<ƌ<�Ί<ֈ<A܆<l�<��<3�<G�}<�y<c�u<u�q<~�m<-�i<�e<i�a<q ^<�Z<rV<bR<�)N<u7J<�FF<zWB<�i><~:<�6<#�2<z�.<��*<�'<�'#<KO<�z<k�<��<g<�[<	�<��<�A<8�;h��;]��;h��;m��;L��;���;C��;3�;�o�;�ص;Z�;��;��;�v�;a�;[h�;���;�̄;hT~;EJs;.zh;��];�S;m^I;Co?;_�5;�0,;�";!�;��;;~!�: g�:��:O �:�K�:��:�͟:��:'o�:�Dh:)L:}a0:�:>"�9�߾97�9�T,9S��8)��h�}Ei�m���׹k�������3�8K���b���y�-���+��q��DԪ��-�� ����̺غ�N㺳����4{�x�����8�
��?S���#�c)���.�Pi4�i�9�]k?�"�D�4nJ�J�O��uU���Z��`�wf���k�_$q��v��=|��䀻`����n��`3��%���㸎��z���<�����������  �  J�=�7=�=/�=-=��=�y= =�� =�k = =�l�<϶�<� �<;J�<s��<P��<�$�<�l�<��<���<�@�<���<���<�<CO�<\��<U��<?�<M�<؉�<���<; �<�9�<sr�<ߩ�<��<��<LH�<�y�<۩�<���<%�<!,�<nR�<�u�< ��<���<��<i��<���<��<�<�<��<��<�	�<'��<,��<���<j��<��<�i�<�9�<��<!��<h��<�4�<t��<��<�%�<ؼ�<M�<s��<Y�<��<�J�<���<A#�<���<&�<<�<���<�۵<�#�<zf�<}��<�ݮ<��<5C�<�o�<���<ѽ�<�ߣ<���<�<�4�<>L�<�a�<�t�<b��<2��<a��<��<E��<&ƌ<�Ί<ֈ<3܆<g�<��<�<��}<w�y<��u<��q<��m<�i<;�e<[�a<��]<�Z<�V<�R<)N< 7J<vFF<dWB<�i><�}:<�6<V�2<��.<O�*<�'<�(#<,P<�{<L�<��<G<�\<�<~�<�B<9�;T��;���;׭�;S��;H��;u��;���;��;�n�;�׵;xX�;J�;1��;�t�;p_�;Yf�;���;�ʄ;vQ~;�Gs;�wh;��];1�S;h^I;�n?;̵5;�1,;c�";�;��;�;�'�:�n�:~�:o�:�R�:!�:�՟:z�:<v�:�Lh:�#L:�f0:0:&�9j۾9�5�9�F,9̊�8������ti��,��q&׹������3�HK�<�b���y�^���"��qt���֪�%/��O����̺�غM㺠��	����x��J���4����WO�z�#�_)�h�.�:f4�4�9��i?�D�D�CmJ���O�|uU�!�Z��`�df��k��&q���v��@|�~总$����p��5��9��������|��V>��������  �  @�=�7=�=,�=-=��=z=) =�� =�k = =�l�<��<� �<dJ�<���<y��<�$�<�l�< ��<���<�@�<ǅ�<���< �<?O�<@��<3��<'�<�L�<���<d��<& �<�9�<Mr�<ĩ�<���<��<*H�<�y�<ɩ�<z��<�<�+�<YR�<�u�<��<���<���<���<���<�<�<+�<��<��<
�<U��<G��<���<���<0��<�i�<�9�<��<2��<a��<�4�<T��<	��<j%�<���<�L�<K��<�X�<���<�J�<ҹ�<#�<~��<��<�;�<k��<�۵<{#�<]f�<u��<�ݮ<��<9C�<�o�<���<꽥<�ߣ<���<A�<�4�<bL�<�a�<u�<v��<9��<���<��<l��<3ƌ<�Ί<ֈ<0܆<M�<n�<��<`�}<V�y<Z�u<[�q<k�m<��i<�e<�a<F�]<�Z<UV<�R<�(N<�6J<(FF<1WB<�i><~:<<�6<o�2<<�.<v�*<'<�(#<QP<W|<��<��<�<�\<��<��<�B<t9�;���;���;7��;���;@��;��;F��;5�;0n�;\׵;�W�;��;���;`t�;_�;�e�;���;Nʄ;�P~;xGs;
wh;}�];�S;�]I;�n?;~�5;�1,;��";+�;j�;�;�'�:`p�:��:�	�:U�:�:]ן:E�:=x�:�Oh:b'L:�h0:,:�*�9)ھ9,2�9�7,9�x�8�����Ui�
6��p*׹�������3�	MK�R�b���y�-���\���u���ت��0�����C�̺Xغ�L������w�v�;���3�}��2N���#�}])���.�f4��9�*i?��D��lJ�5�O��tU�=�Z��`��f���k��'q��v��A|��总�����q��f5������/����|���>�� �����  �  J�=�7=�=/�=-=��=�y= =�� =�k = =�l�<϶�<� �<;J�<s��<P��<�$�<�l�<��<���<�@�<���<���<�<CO�<\��<U��<?�<M�<؉�<���<; �<�9�<sr�<ߩ�<��<��<LH�<�y�<۩�<���<%�<!,�<nR�<�u�< ��<���<��<i��<���<��<�<�<��<��<�	�<'��<,��<���<j��<��<�i�<�9�<��<!��<h��<�4�<t��<��<�%�<ؼ�<M�<s��<Y�<��<�J�<���<A#�<���<&�<<�<���<�۵<�#�<zf�<}��<�ݮ<��<5C�<�o�<���<ѽ�<�ߣ<���<�<�4�<>L�<�a�<�t�<b��<2��<a��<��<E��<&ƌ<�Ί<ֈ<3܆<g�<��<�<��}<w�y<��u<��q<��m<�i<;�e<[�a<��]<�Z<�V<�R<)N< 7J<wFF<dWB<�i><�}:<�6<V�2<��.<O�*<�'<�(#<,P<�{<L�<��<G<�\<�<~�<�B<9�;T��;���;׭�;S��;H��;u��;���;��;�n�;�׵;xX�;J�;1��;�t�;p_�;Yf�;���;�ʄ;vQ~;�Gs;�wh;��];1�S;h^I;�n?;̵5;�1,;c�";�;��;�;�'�:�n�:~�:o�:�R�:!�:�՟:z�:<v�:�Lh:�#L:�f0:0:&�9j۾9�5�9�F,9̊�8������ti��,��q&׹������3�HK�<�b���y�^���"��qt���֪�%/��O����̺�غM㺠��	����x��J���4����WO�z�#�_)�h�.�:f4�4�9��i?�D�D�CmJ���O�|uU�!�Z��`�df��k��&q���v��@|�~总$����p��5��9��������|��V>��������  �  ^�=�7= �=5�=-=��=�y=�=�� =jk =� =7l�<P��<A �<�I�<��<���<W$�<Hl�<���<~��<i@�<���<���<#�<KO�<o��<|��<p�<aM�<)��<���<� �<`:�<�r�<M��<���<V�<�H�<_z�<)��<���<G�<<,�<sR�<�u�<���<��<Y��<-��<Y��<p�<��<��<.�<=�<w	�<���<���<K��<���<ޒ�<\i�<e9�<��<��<~��<�4�<���<J��<�%�<-��<{M�<���<zY�<���<K�<x��<�#�<��<��<w<�<鎷<�۵<�#�<�f�<���<�ݮ<��<#C�<�o�<W��<���<uߣ<y��<��<f4�<�K�<a�<[t�<<ϕ�<���<հ�<��<ƌ<�Ί<ֈ<A܆<l�<��<3�<G�}<�y<c�u<u�q<~�m<-�i<�e<i�a<q ^<�Z<rV<bR<�)N<u7J<�FF<zWB<�i><~:<�6<#�2<z�.<��*<�'<�'#<KO<�z<k�<��<g<�[<	�<��<�A<8�;h��;]��;h��;m��;L��;���;B��;2�;�o�;�ص;Z�;��;��;�v�;a�;Zh�;���;�̄;hT~;DJs;.zh;��];�S;m^I;Co?;_�5;�0,;�";!�;��;;~!�: g�:��:O �:�K�:��:�͟:��:'o�:�Dh:)L:}a0:�:>"�9�߾97�9�T,9S��8)��h�}Ei�m���׹k�������3�8K���b���y�-���+��q��DԪ��-�� ����̺غ�N㺳����4{�x�����8�
��?S���#�c)���.�Pi4�i�9�]k?�"�D�4nJ�J�O��uU���Z��`�wf���k�_$q��v��=|��䀻`����n��`3��%���㸎��z���<�����������  �  ��=�7=7�=:�=-=�=�y=�=�� =.k =� =�k�<���<���<I�<T��</��<�#�<�k�<2��<��<@�<]��<���<�<]O�<���<���<��<�M�<���<���<S�<;�<�s�<��<C��<�<YI�<�z�<���<P��<��<�,�<�R�<�u�<��<���<��<���<���<��<�<��<��<��<��<��<��<���<���<c��<�h�<9�<x�<
��<���<�4�<���<���<I&�<���<N�<���<:Z�<M��<�K�<C��<y$�<�<@�<=�<k��<dܵ<($�<�f�<���<�ݮ<x�<�B�<Jo�<ꗧ<��<�ޣ<���<�<�3�<K�<a`�<�s�<L��<4��<���<R��<���<�Ō<_Ί<�Ո<G܆<��<��<��<�}<"�y<��u<��q<��m<��i<��e<��a<�^<
Z<�V<vR<�*N<U8J<]GF<�WB<�i><�}:<��6<��2<��.<��*<�'<�&#<�M<�y<�</�<�<=Z<��<q�<�@<6�;��;��;���;��;g��;L��;\��;��;�q�;�ڵ;A\�;f��;t��;}y�;d�;�j�;B��;�΄;�X~;�Ms;K}h;��];ՆS;`_I;o?;��5;�.,;��";�;��;1;c�:~\�:B��:���:�?�:ܮ:dß:
��:~g�:�4h:�L:�W0:�:�9r޾9�>�92u,9��8|U��*�Z�h��ꥹ��ֹ�����3��#K�Βb�O�y�{������fj��	Ϫ��)���}��S�̺	غS㺍�������������=�����X���#�h)��.�$n4�'�9�mo?���D��pJ�!�O��uU�h�Z���`�:f�k�k�� q��v��8|�7※����.l��20��l�9���Tx��B:��l��������  �  Ӑ=(8=V�=A�=�,=m�=�y=�=M� =�j =+ =�j�<Ǵ�<���<.H�<\��<N��<�"�<�j�<���<w��<�?�<��<���<
�<zO�<��<*��<e�<kN�<z��<X��<@�<�;�<�t�<��<%��<�<0J�<�{�<W��<���<�<�,�<�R�<�u�<ϕ�<m��<���<U��<5��<C�<B�< �<��<��<��<��<;��<���<δ�<���<�h�<�8�<G�<���<���<5�<0��<*��<�&�<m��<�N�<s��<@[�<A��<�L�<I��<v%�<�<�<�=�<��< ݵ<�$�<0g�<ݤ�<�ݮ<j�<�B�<�n�<k��<n��<4ޣ<	��<(�<�2�<2J�<o_�<�r�<t��<`��<Т�<���<=��<dŌ<4Ί<�Ո<I܆<��<M�<�<<�}<��y<�u<r�q<��m<R�i<��e<��a<�^<�Z<7V<�R<�+N<[9J<HF<`XB<j><�}:<?�6<�2<��.<��*<�'<�$#<=L<�w<��<^�<�<eX<�<��<\?<�3�;I��;���;���;���;���;��;���;� �;�s�;�ݵ;5_�;���;��;}�;�g�;2n�;���;�ф;�^~;#Ss;j�h;�];ÈS;�`I;�n?;��5;�,,;��";	�;i�;K;�	�:�N�:���:���:=1�:�̮:���:k�:v[�:Dh:�K:�L0::�:��9�ܾ9gK�9��,9�x�8(< ���[�h�����:�ֹ{�����Bf3�+K��tb���y��n����a���Ȫ��%��E{���̺�غ�W�H��b���N����l���D�D���_�J�#�|o)���.��t4���9�Qt?�Y�D�'sJ�j�O��vU�E�Z���`��f���k��q�D�v��2|��ހ������h��A,���_����t��07�����������  �  �=[8=r�=P�=�,=P�=my=M=�� =oj =� =�i�<���<���<	G�<I��<G��<�!�<j�<Ǳ�<���<&?�<���<]��<�<�O�<(��<���<��<!O�<F��<F��<7�<=�<�u�<#��<G��<�<'K�<�|�<��<���<��<-�<�R�<�u�<���<)��<8��<���<���<d �<Y
�<%�<��<��<��<��<=��<���<��<��<�g�<O8�<�<���<���<45�<���<���<�'�<;��<�O�<y��<L\�<v��<N�<q��<�&�<͉�<�<�>�<␷<�ݵ<%%�<�g�<��<�ݮ<J�<XB�<rn�<֖�<���<Vݣ<��<%�<�1�<I�<b^�<�q�<x��<{��<���<��<���<�Č<�͊<�Ո<c܆<��<��<��<��}<�y<��u<c�q<��m<��i<��e<��a<�^<�Z<V<�!R<N-N<q:J<�HF<�XB<`j><�}:<Β6<�2<��.<b�*<��&<##<<J<�u<å<��<�<<V<�<��<�=<�0�;���;���;��;G��;ܢ�;޹�; ��;�"�;Fv�;��;�b�;���; ��;1��;�k�;�r�;���;�Մ;e~;�Xs;[�h;��];�S;�aI;�n?;q�5;X*,;o�";�;��;
;���:�>�:���:G��:��:i��:K��:Zא:3M�:�	h:�K:x;0:��:}�9�޾9�S�9q�,9l��8�����w�w-h��x���bֹAm��r��C3���J��Ub�ݟy��a���䓺X��D���d!��Py����̺�غ@]�y��P�����$���M�����h���#��w)���.��{4�p�9�|y?�*�D��vJ�Y�O�5wU�d�Z�"`��f�{�k��q��v��+|��ڀ�����d���'��V닻*����p���3��[���幙��  �  X�=�8=��=Y�=�,=+�=:y= =�� = j =B =�h�<���<Z��<�E�<%��<��<� �<&i�<��<��<�>�<U��<��<��<�O�<p��<��<��<�O�<$��<T��<H�<+>�<�v�<K��<v��<�<:L�<�}�<��<+��<�<�-�<#S�<�u�<x��<ڱ�<���<��<���<���<e	�<�<q�<[�<��<���<��< ��<��<S��<Ig�<�7�<��<���<���<k5�<��<D��<C(�<!��<�P�<���<r]�<���<\O�<���<�'�<���<F�<�?�<đ�<K޵<�%�<�g�<=��<�ݮ<�<B�<�m�<.��<�<{ܣ<!��<�<�0�<�G�<8]�<�p�<[��<���<��<D��< ��<�Č<�͊<�Ո<p܆<3�<�<�<�}<��y<��u<��q<�m<�i<8�e<Rb<"^<Z<'V<J#R<�.N<�;J<�IF<[YB<�j><r}:<>�6<H�2<��.<��*<.�&<2!#<H<>s<\�<w�<L<�S<��<��<�;<�-�;>��; ��;���;���;��;���;���;�$�;&y�;��;�f�;��;[��;ą�;<p�;w�;Ù�;�ل;=l~;_s;�h;g�];�S;�bI;�n?;m�5;�',;��";`�;K�;;���:.,�:~��:���:��:Q��:咟:�ǐ:?�:F�g:I�K:�+0:��:���9߾9�]�9J�,9�r�8��4�H�g�4��uֹ�G�jM��3���J��3b��}y��S���ד�SO�����P��Vw����̺�غ�b㺪����ܐ�1+���FV�����r�#�#��)��/�g�4�c:��?��D�zJ���O��xU���Z�g}`�@f�k�k�Rq�r�v��#|��ր�P���b_��a#���拻˩���l��/��������  �  ��=�8=��=h�=�,=
�=�x=�==� =�i =� =�g�<}��<)��<�D�<���<��<��<*h�<��<o��<>�<��<���<��<�O�<���<��<!�<�P�<��<F��<h�<K?�<x�<���<���<7�<9M�<h~�<ĭ�<���<��<�-�<cS�<�u�<X��<���<Q��<���<���<���<U�<��<R�<0�<o�<���<��<���<8��<���<�f�<s7�<k�<���<���<�5�<c��<щ�<)�<��<�Q�<���<�^�<���<�P�< ��<)�<,��<P�<�@�<���<ߵ<1&�<Lh�<���<�ݮ<��<�A�<�m�<���<%��<�ۣ<��<��<p/�<�F�<\�<�o�<J��<{��<8��<|��<s��<Č<Z͊<yՈ<�܆<w�<t�<��<~�}<~�y<��u<��q<n�m<S�i<��e<�b<y
^<FZ<
V<%R<Z0N<�<J<�JF<�YB<�j><K}:<��6<_�2<��.<[�*<x�&<#<�E<�p<�<�<�<�Q<l�<��<:<�*�;���;"��;f��;0��;y��;���;��;�&�;�{�;"�;)j�;��;���;A��;�t�;C{�;��;~݄;�r~;ees;D�h;�];R�S;�dI;�n?;"�5;�$,;��";��;��;��;p��:��:��:{��:���:���:���:S��:[0�:��g:��K:0:g�:x��9�߾9vl�9�-9r�8������*Gg�]�����չ $�\&��2���J�Ob�_y��E���ʓ��D��粪�a���s��y�̺�غ<i㺢���������2�����^�X���{��$�؉)�/�ȋ4�;	:�Ѕ?�hE��}J���O�hyU�:�Z�5{`�S�e��k�qq���v�l|�dҀ������Z��{���ዻ1���Qh���+��������  �  �=�8=��=o�=�,=��=�x=y=�� =.i =I =�f�<o��<
��<�C�<Ռ�<��<��<Ig�<R��<���<�=�<���<���<��<�O�<���<���<��<XQ�<ގ�<,��<c�<Y@�<!y�<���<���<@�<,N�<O�<z��<{��<0�<2.�<�S�<�u�<8��<=��<���<���<;��<���<h�<��<6�<!�<d�<���< ��<��<m��<Ԏ�<#f�<�6�<)�<���<���<�5�<���<m��<�)�<���<�R�<���<�_�<��<�Q�<&��<3*�<<��<L�<�A�<`��<�ߵ<�&�<�h�<���<�ݮ<��<jA�<m�<�<k��<�ڣ<&��<�<S.�<�E�<�Z�<sn�<S��<���<k��<Ĭ�<㸎<�Ì<͊<XՈ<�܆<��<��<<�<��}<�y<��u<��q<��m<}�i< f<�b<�^<AZ<�V<�&R<�1N<�=J<{KF<nZB<�j><}:<P�6<��2<q�.<��*<��&<;#<�C<�n<��<��<{<nO<c�<��<k8<�'�;���;m��;k��;���;���;a��;���;�(�;V~�;U�;�m�;t	�;���;F��;!y�;]�;	��;�;�y~;�js;ߔh;I�];ĒS;�eI;�n?;ܭ5;!",;��";��;��;�;6��:�:��:%��:��:_��:�q�:��:-#�:�g:�K:�0:��:���9oݾ9)w�9�?-9�|�8P���L�n�f����!�չ��?���2��xJ���a��Ay��7��S���;��ݪ��,��r����̺Gغ�n�ܷ���������9�c���f�f��w���$�o�)��/�4�4��:�}�?��E�9�J���O�^zU���Z��y`�3�e�?�k�~q�H�v�C|��΀������V������݋����od��=(��Q얻~����  �  $�=#9=��=y�=�,=��=�x=8=�� =�h =� =�e�<y��<"��<�B�<��<��<��<�f�<���<0��<=�<<��<{��<��<P�<)��<J��<+�<�Q�<���< ��<;�<GA�<z�<���<���<�<O�<��<#��<��<��<v.�<�S�<�u�<��<���<r��<\��<���<��<��<�<P�<-
�<n�<���<0��<:��<���<4��<�e�<�6�<� �<Z��<р�<6�<��<ӊ�<>*�<~��<�S�<���<�`�<��<�R�<$¿<5+�<$��<4�<nB�<��<7�<''�<�h�<ץ�<ޮ<��<,A�<�l�<l��<���<�٣<T��<�<u-�<�D�<Z�<�m�<h�<Ï�<���<,��<[��<9Ì<�̊<=Ո<�܆<��<#�<��<��}<]�y<�u<X�q<J�m<t�i<�f<�b<h^<Z<�V<(R<�2N<�>J<'LF<�ZB<#k><�|:<Ր6<�2<m�.<��*<Z�&<�#<�A<�l<��<��<�<eM<��<T�<�6<F%�;���;���;J��;F��;���;Լ�;���;o*�;���;��;�p�;��;¢;ؑ�;}|�;��;T��;Y�;�~;�os;Șh;��];��S;2fI;�n?;Q�5;�,;E�";�;��;��;��:���:*��:���:ؽ:�u�:�b�:���:q�:��g:<�K:��/:4�:F��9A߾9}�9�]-9Iԍ8 P�����tf�����A]չ�����9�2��ZJ���a��&y�},��9����3������$���p��a�̺�"غIs����-���?�#���n�r��X��$� �)�./�z�4��:�2�?��	E��J���O�"{U�_�Z��x`���e�}k��q��v��|�ˀ�
����R��m���ً�y����`��%���閻����  �  M�=I9=��=~�=�,=��=zx==b� =�h =� =e�<Ѯ�<s��<�A�<I��<]��<[�<�e�<��<���<�<�<���<Q��<��< P�<g��<���<��<yR�<��<���<��<�A�<�z�<9��<M��<��<�O�<���<���<t��<��<�.�<�S�<�u�<���<���<��<���<'��<���<	�<b�<��<o	�<��<7��<���<���<��<���<:e�<F6�<� �<G��<���</6�<Z��<(��<�*�<��<T�<B��<^a�<���<�S�<�¿<�+�<؎�<��<�B�<���<��<}'�<-i�<�<ޮ<��<�@�<Kl�<��<J��<m٣<���<[�<�,�<�C�<NY�<�l�<�~�<0��<��<���<뷎<�<�̊<+Ո<�܆<��<m�<��<��}<U�y<:�u<��q<��m<��i<.f<?	b<�^<MZ<�V<)R<�3N<?J<�LF<"[B<;k><�|:<u�6<I�2<��.<��*<I�&<v#<�@<xk<J�<-�<?<�K<J�<�<�5<l#�;���;���;w��; ��;���;���;���;�+�;v��;��;�r�;�;Ģ;���;,�;���;���;��;f�~;Uss;�h; �];��S;�fI;�n?;t�5;�,;r�";��;��;��;���:���:Ό�:U��:�˽:�k�:JW�:���:5�:��g:�K:&�/:7�:`��9��9���9�-9 �8��򷘸��6f�^[��4չ��������2��EJ��a�:y�%������-��𠪺����o����̺%غ�w�W��G�����D����5t�������$�6�)�o /��4��:���?�pE���J�� P��{U��Z�Bw`�h�e��zk��p�2�v�p
|��Ȁ�|����O������֋�󚎻x^���"���疻)����  �  i�=U9=�=z�=�,=��=hx=�=8� =dh =d =�d�<[��<���<cA�<�<���<��<�e�<̭�<s��<�<�<ڂ�<K��<��<#P�<���<���<��<�R�<p��<���<T�<iB�<:{�<���<���<?�<P�<��<��<���<�<�.�<�S�<�u�<��<���<���<���<���<-��<��<�
�<.�<��<<�<���<��<;��<ï�<s��<�d�<"6�<� �<G��<Ԁ�<F6�<|��<Z��<�*�<S��<�T�<���<�a�<F��<T�<cÿ<k,�<X��<K�<iC�<䔷<��<�'�<Oi�< ��<�ݮ<��<�@�<.l�<���<���<
٣<L��<��<J,�<C�<�X�<bl�<R~�<���<ʝ�<h��<���<�<�̊< Ո<�܆<�<��<"�<<�}<�y<�u<t�q<��m<��i<.f<
b<�^<*Z<� V<�)R<O4N<�?J<�LF<U[B<.k><�|:<b�6<�2<=�.<8�*<��&<�#<�?<�j<<�<H�<'
<K<V�<5�<#5<"�;��;(��;D��;���;���;��;-��;�,�;;��;"�;Vt�;��;aƢ;=��;��;H��;���;@�;��~;�us;��h;X�];b�S;[gI;*n?;2�5;�,;�";��;�;B�;]��:���:���:�x�:�Ľ:Kc�:�P�:4��:��:��g:��K:*�/:��:��9�ܾ9���9g�-9�K�8��*����e�A���չ]�������2�m6J�	�a��y���V����)������J
��,o����̺Z%غ7y�p�� ������G�����w������$��)��#/���4�~:�9�?��E���J�P��{U�|�Z��v`���e�yk�m�p�X�v�$|��ƀ�����#N�����KՋ������\�� !��<斻U����  �  G�=�<=��=��=31=�=�}=X#=�� =qn =� =+r�<ļ�<a�<R�<���<e��<�1�<m|�<���<�<*Y�<_��<���<V/�<�t�<��<2��<->�<�<Ⱦ�<]��<�:�<w�<,��<��<�$�<�[�<'��<���<���<B&�<�S�<J~�< ��<��<���<T�<\&�<�=�<�Q�<�a�<�m�<v�<z�<�y�<�t�<`k�<�\�<�H�<)/�<y�<���<��<f��<�N�<��<��<�q�<��<n��<GP�<���<�i�<w��<%f�<��<%G�<ڭ�<4�<ah�<���<�<�S�<4��<Xղ<G�<uB�<r�<��<Nĩ<��<��<�$�<�>�<V�<gk�<�~�<c��<i��<�<)��<Ȓ<�Ґ<�ێ<��<��<`��<��<*��<���<���<;�}<��y<	�u<��q<��m<�i<=�e<��a<�]<�Y<9�U<K�Q<Y�M<�J<9
F<�B<�><e%:<�16<�?2<QP.<�c*<z&<,�"<g�<\�<m�<+<�^<T�<��<�<n <׆�;�@�;_	�;���;H��; ��;���;���;R)�;hs�;�Գ;YM�;1ߦ;?��;$R�;s5�;5�;HR�;���;��y;F�n;J�c;0>Y;��N;��D;�:;U1;�|';.;�;=/;~;���:�a�:9'�:�J�:2ȵ:���:���:V4�:^�u:�Y:�I>:$+#:~q:G)�9�9�-i9j\9���7ܴ��lE(�� ��2��� ��q�
�-{"�2�9�xOQ�1|h����Z8��&��������Q��b�����ú�+Ϻ�lں*��l�����3��j;	�3��Z�d���e���$��\*���/�'C5���:�T@�n�E���J�UfP�*�U��H[���`�;5f��k��,q�f�v��)|�Հ������U��U���Ջ�A����U�����ז�o����  �  ?�=�<=��=��=21=��=�}=e#=� =}n =� =gr�<���<��<AR�<���<���<42�<�|�<���<<�<CY�<���<���<W/�<�t�<���<��<#>�<�~�<���<,��<�:�<�v�<���<���<^$�<u[�<���<���<���<?&�<sS�<(~�<��<��<���<c�<u&�<�=�<�Q�<�a�<n�<Mv�<Vz�<z�<:u�<�k�<�\�<�H�<=/�<��<���<���<z��<�N�<��<��<�q�<��<f��<1P�<���<xi�</��<�e�<���<�F�<���<��</h�<r��<�
�<�S�<��<9ղ<>�<qB�<�q�<@��<cĩ<��<��<�$�<�>�<IV�<�k�<�<���<���</��<U��<'Ȓ<�Ґ<܎<�<��<[��<��<��<i��<���<;�}<T�y<��u<d�q<�m<��i<��e<?�a<��]<��Y<��U<��Q<V�M<�J<
F<�B<�><`%:<�16<�?2<�P.<�c*<Nz&<~�"<�<��<��<{+<_<˘<�<! <Qn <W��;A�; 
�;���;Z��;&��;3��;n��;6)�;Zs�;�ӳ;�L�;(ަ;>��;hQ�;�4�;?4�;?Q�;֋�;��y;��n;D�c;�=Y;��N;��D;d�:;)1;Q}';�.;c;g0;�~;- �:Se�:+�:�N�:7̵:ş�:aŗ:�7�:�u::�Y:�L>:�-#:Ct:D'�9��9,(i9iK9���7_���5O(�+��쿵�����
���"��:��WQ�>�h�X���:��¡��F���S�����G�ú�+Ϻ�lں��������K���:	�v��^X�q���c���$�[*��/��A5��:�2@���E���J��eP�U�U��H[�0�`�6f�|�k��,q�x�v��*|��Հ����PV��<��a֋�Q���rV������ז�p����  �  �=�<=��=��=<1=��=�}=�#=;� =�n =  =�r�<���<8�<�R�<���<)��<�2�<}�<��<��<�Y�<á�< ��<f/�<�t�<ٸ�<���<�=�<�~�<��<���<:�<Uv�<j��<;��<�#�<�Z�<|��<A��<��<�%�<+S�<~�<���<��<���<��<�&�<L>�<HR�<Zb�<�n�<�v�<�z�<�z�<�u�<)l�<~]�<yI�<�/�<�<���<A��<���<�N�<��<���<�q�<��<���<�O�<���<�h�<���<Te�<��<OF�<��<_�<�g�<껹<|
�<cS�<ݖ�<ղ<-�<sB�<
r�<p��<�ĩ<*�<<�<%�<A?�<�V�<9l�<��<:��</��<���<ڼ�<�Ȓ<)Ӑ<M܎<K�<��<p��<��<���<C��<���<q�}<W�y<��u<j�q<��m<��i<p�e<&�a<p�]<��Y<��U<��Q<��M<�J<�	F<�B<�><�%:<�16<n@2<Q.<�d*<E{&<��"<��<��<(�<�,<J`<�<H�<4!<[o <"��;9B�;�;c��;���;0��;���;���;�'�;�q�;ҳ;�J�;Uܦ;E��;EO�;,2�;42�;8O�;��;��y;��n;O�c;�;Y;z�N;)�D;ּ:;1;�~'; 1;E;K4;��;��:Dn�:'4�:X�:xյ:㨦:7Η:Q@�:��u:��Y:�X>:�6#:�z:U-�9��9:!i9�79��7����(��J�� ߵ�c���
� �"�,:�vhQ��h����B������5���V��p�����ú.+Ϻ�kں�庽����\���6	���T�����^���$��V*���/��=5��:��@�Z�E���J��dP���U��H[��`�F7f���k��/q�i�v��.|��׀�6���yX������؋�o���eX������ٖ�����  �  ݔ=]<=��=��=I1=��=�}=�#=�� =o =� =�s�<���<4	�<�S�<���<#��<�3�<�}�<���</�<Z�<	��<K��<q/�<�t�<���<���<N=�<�}�<|��<���</9�<cu�<k��<F��<�"�<Z�<���<���<}��<M%�<�R�<�}�<إ�<��< ��<��<'�<�>�<�R�<(c�<mo�<�w�<�{�<�{�<�v�<%m�<l^�<BJ�<�0�<��<t��<���<ۉ�<�N�<��<���<Qq�<+�<b��<O�<8��<�g�<���<Ed�<��<AE�<���<q�<�f�<2��<�	�<�R�<s��<�Բ< �<iB�<Gr�<���<ũ<��<��<�%�<@�<�W�<1m�<���<6��</��<���<���<fɒ<�Ӑ<�܎<��<A�<���<��<���<���<$��<H�}<%�y<&�u<��q<�m<��i<��e<�a<��]<��Y<5�U<��Q<F�M<�J<	F<B<�><�%:<z26<A2<R.<�e*<�|&<4�"<ε<��<0<�.<Rb<��<�<�"<�p <}��;jD�;q�;���;!��;���;+��;���;>&�;�o�;�ϳ;�G�;٦;���;|K�;�.�;a.�;�K�;���;F�y;��n;1�c;�8Y;��N;:�D;n�:;�1;�';f4;�;�8;M�;��:_}�:MD�:Th�:��: ��:�ݗ:IM�:�v:��Y:�i>:0D#:U�:=�9��9�i9�90 �7]���v�(�x��[���C湵��"��4:�G�Q���h�(��OM��M���&��2\�������ú�*Ϻ�fں��9����H���/	����AL�����V���$��N*�|�/�075���:�@�&�E���J��bP���U�rI[�{�`��9f�>�k�v4q�-�v�!5|�Zۀ�⛃�~\������܋�%����[�����ܖ�q����  �  ��=<={�=��=Q1=��=~=&$=�� =�o = =�t�<ƿ�<l
�<"U�<���<_��<�4�<�~�<���<��<�Z�<q��<���<w/�<t�<W��<��<�<�<!}�<���<���<8�<%t�<+��<��<�!�<�X�<���<���<���<�$�<?R�<F}�<���<���<F��<#�<�'�<�?�<�S�<!d�<�p�<�x�<}�<�|�<x�<Sn�<�_�<TK�<|1�<q�<(��<(��<(��<O�<��<���<�p�<��<���<N�<.��<�f�<w��<�b�<���<�C�<���<:�<�e�<1��<��<R�<ו�<XԲ<��<\B�<tr�<���<�ũ<^�<�	�<�&�<"A�<�X�<_n�<ځ�<p��<h��<α�<���<_ʒ<�Ԑ<�ݎ<!�<��<���<��<���<x��<���<��}<^�y<�u<i�q<��m<�i< �e<��a<�]<��Y<�U<��Q<��M<� J<�F<�B<{><�%:<�26<�A2<�S.<ag*<�~&<\�"<,�<��<�<s1<�d<��<l�<.%<�r <ӎ�;aG�;[�;	��;���;���;F��;���;
$�;�l�;a̳;�C�;�Ԧ;��;�F�;*�;�)�;vG�;���;��y;�n;��c;�4Y;A�N;i�D;��:;l1;�';�8;�";�?;V�;�'�:Ԑ�:�W�:P|�:���:`̦:�:�^�:�,v:�Z:��>:eV#:~�:I�9��9� i9��9��7�V��MD)�̵��m\��\��o-���"��\:�4�Q���h�k��\��ڿ������d������J�ú�*Ϻcں�������� ���'	����xB�H���L�
�$��D*�(�/��.5�G�:��@�U~E�$�J�V`P���U��I[���`��=f�κk��:q�K�v�E=|��߀������a��c!���ዻ�]`������ߖ������  �  :�=�;=N�=�=h1=	�=]~=y$=^� =p =� =Vv�<*��<��<�V�<:��<���<6�<��<���<��<K[�<���<���<�/�<[t�<���<���<�;�<6|�<o��<���<�6�<�r�<���<���<0 �<xW�<J��<d��<���<�#�<�Q�<�|�<q��<��<r��<��<2(�<I@�<�T�<2e�<�q�<Nz�<�~�<T~�<�y�<�o�<�`�<�L�<�2�<t�<���<���<���<=O�<��<G��<Up�<��<���<M�<���<�e�<���<va�<,��<YB�<*��<�	�<Ld�<�<��<AQ�<7��<�Ӳ<��<kB�<�r�<o��<2Ʃ<&�<�
�<�'�<uB�<OZ�<�o�<X��<ꔚ<Ф�<*��<��<s˒<�Ր<Cގ<��<��<���<��<U��<��<���<�}<?�y<��u<��q<��m<(�i<��e<��a<D�]<��Y<��U<��Q<��M<X�I<�F<�B<G><!&:<�36<C2<�T.<Ii*<ۀ&<�"<�<f�<�<�4<�g<o�<G�<�'<u <���;(J�;��;~��;u��;���;��;$��;l!�;=i�;(ȳ;M?�;�Ϧ;�z�;,A�;$�;V$�;B�;�}�;"�y;a�n;��c;I0Y;D�N;��D; �:;#1;�';�=;�(;UH;�;�<�:���:No�:���:/�:�:��:bt�:BOv:�:Z:��>:ii#:s�:�T�9��9��h9��9���7'��M�)���������a���Y��#���:���Q�� i�q��Xn���Ζ��"��Am��ӱ����ú�(Ϻk_ں���9���������	�����7�V���@�(�$��9*�M�/��$5���:��@��xE���J�$]P�^�U�	J[�{�`�ZAf�!�k��Aq���v��F|��䀻.���/g���'��W狻�����e���$���㖻����  �  ԓ=�;=$�=q�=u1=1�=�~=�$=�� =�p =S =�w�<���<��<2X�<٢�<6��<u7�<\��<���<��<\�<���<��<�/�<-t�<���<���<;�<G{�<>��<F��<95�<<q�<-��<���<��<�U�<��<��<���<�"�<�P�<n|�<"��<��<���<�<�(�<&A�<�U�<cf�<#s�<�{�<��<��<{�<Wq�<Pb�<�M�<�3�<��<���<[��<���<`O�<x�<���<�o�< �<���<�K�<���<d�<U��<�_�<���<�@�<���<%�<�b�<���<��<LP�<|��<mӲ<I�<bB�<�r�<鞫<�Ʃ<�<��<1)�<�C�<�[�<oq�<ᄜ<���<X��<���<S��<�̒<�֐<ߎ<e�<S�<
�<��<��<���<(��<9�}<
�y<&�u<��q<��m<�i<��e<��a<!�]<��Y< �U<R�Q<��M<��I<�F<1B<><P&:<M46<ZD2<uV.<fk*<.�&<��"<ʽ<��<
<�7<Lk<��<1�<`*<ow <��;�M�;��;���;��;a��;��;��;g�;�e�;�ó;K:�; ʦ;�t�;_;�;*�;��;5<�;�x�;A�y;��n;��c;�*Y;a�N;��D;y�:;�1;��';�C;,0;BQ;��;�R�:���:҈�:J��:�+�:���:|�:b��:�vv:^Z:5�>:A�#:6�:�a�9�9,�h9�{9��7%��7B*��P�����GH���6>#��:�R��0i�C��􁋺�ݖ�K0��mw��f���\�ú�'Ϻ�[ں���b���������	����,�p��24�M�$�E-*�+�/�	5���:�^�?�`rE�C�J�_ZP�a�U��J[��`�Ef�O�k��Hq���v�Q|��ꀻZ���8m���-��f틻����^k���)���薻�����  �  o�=O;=��=d�=�1=[�=�~=G%=Z� =>q =� =0y�<6��<�<�Y�<Z��<���<�8�<���<���<��<�\�<��<a��<�/�<
t�<@��<C��<D:�<6z�<��<���<�3�<�o�<���<k��<�<�T�<��<׾�<s��<�!�<+P�<�{�<��<���<���<\�<�)�<B�<�V�<�g�<{t�<.}�<���<i��<�|�<�r�<�c�<MO�<�4�<p�<���<���<P��<�O�<`�<���<Qo�<T�<ų�<�J�<?��<�b�<���<&^�<���<?�<ॾ<��<ga�<T��<��<VO�<���<�Ҳ<�<RB�< s�<E��<�ǩ<��<��<s*�<-E�<<]�<�r�<m��<��<ݧ�<��<�<�͒<�א<�ߎ<��<��<7�<��<���<���<b��<<�}<��y<��u<+�q<��m<��i<��e<D�a<�]<�Y<]�U<��Q<��M<�I<�F<�B<�><�&:<�46<`E2<X.<Em*<��&<;�"<��<��<><;<on<��<0�<%-<�y <��;�P�;��;���;���;6��;���;���;n�;�a�;n��;W5�;�Ħ;o�;E5�;@�;y�;�6�;Cs�;ěy;6�n;ۻc;�%Y;��N;P�D;��:;01;ʎ';I;W7;Y;�;�h�:��:L��:��:�D�:�:6�:���:��v:b}Z:��>:`�#:9�:�s�9��9=�h9�>9��7A�����*�����sZ��'��"���p#���:�>R�b]i��*������N>�����������ú�'Ϻ�Vں�庇�����Y{�#
	�d����m���'��$�!*�R�/�a5��:���?��kE���J��WP��U�]K[�-�`��If���k��Pq���v�@[|�"���A����s��4���󋻫����p���.��햻߫���  �  �=;=��=O�=�1=��=/=�%=�� =�q =� =z�<���<{�<O[�<å�<(��<%:�<҃�<��<��<x]�<v��<���<�/�<�s�<ն�<���<�9�<5y�<��<���<x2�<En�<��<���<��<$S�<%��<���<d��<!�<�O�<b{�<���<���<��<��<*�<�B�<�W�<�h�<�u�<�~�<��<��<~�<.t�</e�<zP�<6�<b�<S��<���<���<�O�<9�<b��<�n�<��<��<�I�<��<(a�<`��<�\�<=��<j=�<U��</�<�_�<(��<��<�N�<	��<eҲ<��<=B�<4s�<���<ȩ<��<��<�+�<aF�<�^�<Lt�<���<y��<B��<a��<�Ô<�Β<vؐ<���<~�<�<]�<f�<{��<p��<���<u�}<��y<0�u<s�q<�m<��i<��e<=�a<A�]<V�Y<��U<��Q<��M<��I<kF<�B<f><�&:<�56<WF2<�Y.<	o*<��&<��"<x�<��<6<@><`q<��<��<�/<| <���;�S�;��;��;.��;���;���;���;�;F^�;v��;�0�;ÿ�;�i�;�/�;��;��;�1�;n�;W�y;9�n;��c;!Y;��N;��D;޼:;�1;=�';�M;�=;�`;|�;R|�:���:ŷ�:3��:&]�:s,�:�L�:���:��v:+�Z:Y�>:�#:S�:ˀ�9��9��h9S�9���7����U+�冹���
��i���#��;�BlR�
�i��?����������I������Ÿ���ú�'Ϻ]Rں}庇�����Cs�	����j�2��E�x�$��*���/�5�{:���?��eE���J��TP��U��L[���`�NNf�s�k��Wq��v��d|�����ŷ���y��:������4���Qv���3��T񖻐����  �  =�:=��=H�=�1=��=q=�%=0� =?r = =�{�<���<��<~\�<��<T��<>;�<ք�<���<S�<^�<��<���<�/�<�s�<���<7��<�8�<jx�<��<���<L1�<m�<٧�<���<b�<�Q�<��<���<���<U �<�N�<{�<v��<���<��<�<�*�<kC�<�X�<�i�<�v�<��<)��<��<E�<gu�<Kf�<�Q�<�6�<;�<���<��<��<�O�<*�< ��<Sn�<�<��<�H�<���<�_�<��<J[�<���<<�<	��<��<�^�<��<��<�M�<s��<Ҳ<��<1B�<Js�<
��<�ȩ<]�<��<�,�<pG�<�_�<�u�<#��<���<}��<���<�Ĕ<�ϒ<Gِ<Q�<�<\�<p�<a�<@��<	��<��<��}<��y<�u<*�q<��m<_�i<�e<��a<��]<��Y<��U<��Q<P�M<@�I<~F<EB<E><�&:<66<^G2<�Z.<�p*<��&<��"<��<�<�<�@<�s<�<.�<�1<�} <���;sV�;�;��;���;���;���;4��;_�;a[�;ⷳ;�,�;U��;e�;�*�;��;9�;�,�;�i�;��y;�n;�c;wY;4�N;r�D;�:;�1;y�';BR;2C;
h;�;���:���:���: ��:�p�:�@�:�^�:ŉ:0�v:�Z:?:��#:��:���9��9|th9Q�9Q�7�x����+�6%�������F�����#�SG;��R��i��P��Ƶ�����{U��͓��ʸ���úQ'ϺPں�u�ٙ�ú��!l����σ�%�B����o�$�*���/���4��s:�C�?��`E���J�vRP���U��L[���`��Qf���k�
^q��v�$m|��������y~��)?������(����z��8����������  �  ��=�:=��==�=�1=��=�=%&=}� =�r =� =}|�<���<��<p]�<��<<��<<�<���<|��<��<p^�<B��<��<�/�<�s�<F��<���<Q8�<�w�<C��<���<d0�<l�<ۦ�<���<e�<�P�<9��<߻�<���<��<zN�<�z�<.��<���<?��<X�<�*�<�C�<Y�<Uj�<�w�<���< ��<��<;��<av�<&g�<bR�<�7�<��<t��<V��<>��<�O�<,�<���<n�<��<���<	H�<��<_�<��<;Z�<���<;�<���<��<�]�<:��<��<M�<��<�Ѳ<Q�<:B�<fs�<H��<�ȩ<��<"�<<-�<MH�<�`�<�v�<��<���<m��<_��<�Ŕ<|В<�ِ<��<b�<��<��<T�<���<���<���<��}<s�y<l�u<r�q<��m<e�i<��e<��a<��]<6�Y<�U<d�Q<1�M<4�I<�F<�B<><�&:<w66<H2<�[.<�q*<Պ&<l�"<��<��<�<�B<v<�<�<c3<8 <y��;KX�;��;���;/��;D��;���;��;x�;WY�;���;�)�;跦;Ka�;%'�;�	�;v
�;>)�;�f�;F�y;�zn;2�c;Y;~�N;p�D;d�:;.1;�';GU;bG;�l;��;��:��:���:�:��:�P�:m�:{Ӊ:��v:E�Z:�?:��#:��:��9��9�Sh9<�9>��7����,�XZ���)��.�蹽2���#�Tg;�вR���i��]��������]��ș��(θ�"�ú�%ϺzMں
q庐��ձ��tg����|���@��2
�s�$��*��~/���4��n:�`�?�A]E���J��PP���U�KM[���`��Sf���k�Obq���v��s|�{�������b���@C�����!���f~��V;������ִ���  �  _�=�:=}�=4�=�1=��=�=P&=�� =�r =� =�|�<F��<J�<^�<���<���<�<�<��<���<J�<�^�<h��< ��<�/�<�s�<��<���<8�<cw�<ʵ�<F��<�/�<k�<D��<��<��<hP�<���<\��<e��<g�<5N�<�z�<��<���<G��<~�</+�<KD�<�Y�<�j�<x�<��<���<���<Ҁ�<�v�<�g�<�R�<"8�<7�<���<���<`��<�O�<�<���<�m�<9�<��<�G�<���<�^�<y��<�Y�<5��<h:�<`��<S�<g]�<���<x�<�L�<���<|Ѳ<2�<)B�<ss�<h��<8ɩ<B�<��<�-�<�H�<&a�<
w�<���<E��<���<ܹ�<;Ɣ<�В<Sڐ<%�<��<��<��<E�<���<���<X��<�}<|�y<g�u<W�q<q�m<1�i<��e<��a<��]<�Y<��U<i�Q<J�M<��I<bF<dB<�><�&:<�66<ZH2<B\.<�r*<Ջ&<h�"<��<�<<D<3w<'�<�<m4<B� <,��;�Y�;G�;��;;��;��;t��;2��;g�;�W�;5��;�'�;ϵ�;4_�;�$�;��;>�;.'�;�d�;`�y;*wn;$�c;Y;��N;��D;<�:;�1;͘';8W;�J;�p;��;���:�:1��:k�:(��:Y�:Mu�:Jۉ:�	w:��Z:� ?:��#:��:��9�9aHh9D�9��7Ya���M,�Zz���L�����D�d�#��y;���R�]�i�f��/ʋ�]��>c��띭��и���ú|&Ϻ6Lں�n��𺎫���c� ���x���������$�S *��z/��4��j:��?�~ZE�^�J��OP�~�U��M[���`��Uf���k��eq���v��w|������������E�����MÎ�����h=�����������  �  R�=v:=y�=3�=�1=��=�=W&=�� =�r =� =7}�<���<w�<S^�<���<��<�<�<C��<��<K�<�^�<���<4��<�/�<�s�<��<~��<�7�<>w�<���<��<�/�<Ek�<��<���<��<1P�<u��<E��<G��<L�<N�<gz�<��<���<O��<��<A+�<SD�<�Y�<�j�<;x�<L��<��<܅�<��<#w�<�g�<S�<H8�<H�<���<���<��<�O�<�<���<�m�< �<���<aG�<y��<O^�<<��<_Y�<���<":�<!��<�<2]�<���<O�<�L�<���<kѲ<6�<B�<�s�<���<Jɩ<B�<��<�-�<�H�<la�<<w�<�<t��<7��<��<mƔ<'ђ<Xڐ<1�<��<��<��<D�<���<^��<?��<��}<F�y<*�u<��q<��m<��i<P�e<�a<#�]<��Y<��U<6�Q<�M<l�I<F<TB<�><�&:<�66<�H2<]\.<�r*<$�&<ƨ"<
�<��<a<D<�w<��<��<�4<�� <;��;�Y�;��;���;3��;@��;S��;���;�;W�;겳;�&�;촦;W^�;�#�;��;P�;Z&�;�c�;��y;Mvn;^�c;tY;ؾN;/�D;I�:;�1;ę';�W;�J;�p;��;���:��:W��:��:׍�:�\�:�y�:�݉:�w:��Z:k!?:5�#:��:���9#�9XLh9�9�)�7)z���],����Z��p�蹀L�b$�1�;�)�R���i� i���ˋ�����d�������Ѹ��ú'Ϻ+Kں�l庯��l����b����Fw����\��9�{�$�:�)��x/�u�4��i:���?�"ZE���J��NP�~�U��M[���`�Wf���k��fq���v��x|�� ���Ã�����F�����7Ď������=��=�������  �  _�=�:=}�=4�=�1=��=�=P&=�� =�r =� =�|�<F��<J�<^�<���<���<�<�<��<���<J�<�^�<h��< ��<�/�<�s�<��<���<8�<cw�<ʵ�<F��<�/�<k�<D��<��<��<hP�<���<\��<e��<g�<5N�<�z�<��<���<G��<~�</+�<KD�<�Y�<�j�<x�<��<���<���<Ҁ�<�v�<�g�<�R�<"8�<7�<���<���<`��<�O�<�<���<�m�<9�<��<�G�<���<�^�<y��<�Y�<5��<h:�<`��<S�<g]�<���<x�<�L�<���<|Ѳ<2�<)B�<ss�<h��<8ɩ<B�<��<�-�<�H�<&a�<
w�<���<E��<���<ܹ�<;Ɣ<�В<Sڐ<%�<��<��<��<E�<���<���<X��<�}<|�y<g�u<W�q<q�m<1�i<��e<��a<��]<�Y<��U<i�Q<J�M<��I<bF<dB<�><�&:<�66<ZH2<B\.<�r*<Ջ&<h�"<��<�<<D<3w<'�<�<m4<B� <,��;�Y�;F�;��;;��;��;t��;2��;g�;�W�;5��;�'�;ϵ�;4_�;�$�;��;>�;.'�;�d�;_�y;*wn;$�c;Y;��N;��D;<�:;�1;͘';8W;�J;�p;��;���:�:1��:k�:(��:Y�:Mu�:Jۉ:�	w:��Z:� ?:��#:��:��9�9aHh9D�9��7Ya���M,�Zz���L�����D�d�#��y;���R�]�i�f��/ʋ�]��>c��띭��и���ú|&Ϻ6Lں�n��𺎫���c� ���x���������$�S *��z/��4��j:��?�~ZE�^�J��OP�~�U��M[���`��Uf���k��eq���v��w|������������E�����MÎ�����h=�����������  �  ��=�:=��==�=�1=��=�=%&=}� =�r =� =}|�<���<��<p]�<��<<��<<�<���<|��<��<p^�<B��<��<�/�<�s�<F��<���<Q8�<�w�<C��<���<d0�<l�<ۦ�<���<e�<�P�<9��<߻�<���<��<zN�<�z�<.��<���<?��<X�<�*�<�C�<Y�<Uj�<�w�<���< ��<��<;��<av�<&g�<bR�<�7�<��<t��<V��<>��<�O�<,�<���<n�<��<���<	H�<��<_�<��<;Z�<���<;�<���<��<�]�<:��<��<M�<��<�Ѳ<Q�<:B�<fs�<H��<�ȩ<��<"�<<-�<MH�<�`�<�v�<��<���<m��<_��<�Ŕ<|В<�ِ<��<b�<��<��<T�<���<���<���<��}<s�y<l�u<r�q<��m<e�i<��e<��a<��]<6�Y<�U<d�Q<1�M<4�I<�F<�B<><�&:<w66<H2<�[.<�q*<Պ&<l�"<��<��<�<�B<v<�<�<c3<8 <x��;KX�;��;���;/��;D��;���;��;x�;WY�;���;�)�;跦;Ka�;$'�;�	�;v
�;>)�;�f�;F�y;�zn;1�c;Y;~�N;p�D;d�:;.1;�';GU;bG;�l;��;��:��:���:�:��:�P�:m�:{Ӊ:��v:E�Z:�?:��#:��:��9��9�Sh9<�9>��7����,�XZ���)��.�蹽2���#�Tg;�вR���i��]��������]��ș��(θ�"�ú�%ϺzMں
q庐��ձ��tg����|���@��2
�s�$��*��~/���4��n:�`�?�A]E���J��PP���U�KM[���`��Sf���k�Obq���v��s|�{�������b���@C�����!���f~��V;������ִ���  �  =�:=��=H�=�1=��=q=�%=0� =?r = =�{�<���<��<~\�<��<T��<>;�<ք�<���<S�<^�<��<���<�/�<�s�<���<7��<�8�<jx�<��<���<L1�<m�<٧�<���<b�<�Q�<��<���<���<U �<�N�<{�<v��<���<��<�<�*�<kC�<�X�<�i�<�v�<��<)��<��<E�<gu�<Kf�<�Q�<�6�<;�<���<��<��<�O�<*�< ��<Sn�<�<��<�H�<���<�_�<��<J[�<���<<�<	��<��<�^�<��<��<�M�<s��<Ҳ<��<1B�<Js�<
��<�ȩ<]�<��<�,�<pG�<�_�<�u�<#��<���<}��<���<�Ĕ<�ϒ<Gِ<Q�<�<\�<p�<a�<@��<	��<��<��}<��y<�u<*�q<��m<_�i<�e<��a<��]<��Y<��U<��Q<P�M<@�I<~F<EB<E><�&:<66<^G2<�Z.<�p*<��&<��"<��<�<�<�@<�s<�<.�<�1<�} <���;sV�;�;��;���;���;���;4��;^�;a[�;ⷳ;�,�;U��;e�;�*�;��;9�;�,�;�i�;��y;�n;�c;wY;4�N;r�D;�:;�1;y�';BR;2C;
h;�;���:���:���: ��:�p�:�@�:�^�:ŉ:0�v:�Z:?:��#:��:���9��9|th9Q�9Q�7�x����+�6%�������F�����#�SG;��R��i��P��Ƶ�����{U��͓��ʸ���úQ'ϺPں�u�ٙ�ú��!l����σ�%�B����o�$�*���/���4��s:�C�?��`E���J�vRP���U��L[���`��Qf���k�
^q��v�$m|��������y~��)?������(����z��8����������  �  �=;=��=O�=�1=��=/=�%=�� =�q =� =z�<���<{�<O[�<å�<(��<%:�<҃�<��<��<x]�<v��<���<�/�<�s�<ն�<���<�9�<5y�<��<���<x2�<En�<��<���<��<$S�<%��<���<d��<!�<�O�<b{�<���<���<��<��<*�<�B�<�W�<�h�<�u�<�~�<��<��<~�<.t�</e�<zP�<6�<b�<S��<���<���<�O�<9�<b��<�n�<��<��<�I�<��<(a�<`��<�\�<=��<j=�<U��</�<�_�<(��<��<�N�<	��<eҲ<��<=B�<4s�<���<ȩ<��<��<�+�<aF�<�^�<Lt�<���<y��<B��<a��<�Ô<�Β<vؐ<���<~�<�<]�<f�<{��<p��<���<u�}<��y<0�u<s�q<�m<��i<��e<=�a<A�]<V�Y<��U<��Q<��M<��I<kF<�B<g><�&:<�56<WF2<�Y.<	o*<��&<��"<x�<��<6<@><`q<��<��<�/<| <���;�S�;��;��;.��;���;���;���;�;F^�;v��;�0�;¿�;�i�;�/�;��;��;�1�;n�;V�y;9�n;��c;!Y;��N;��D;޼:;�1;=�';�M;�=;�`;|�;R|�:���:ŷ�:3��:&]�:s,�:�L�:���:��v:+�Z:Y�>:�#:S�:ˀ�9��9��h9S�9���7����U+�冹���
��i���#��;�BlR�
�i��?����������I������Ÿ���ú�'Ϻ]Rں}庇�����Cs�	����j�2��E�x�$��*���/�5�{:���?��eE���J��TP��U��L[���`�NNf�s�k��Wq��v��d|�����ŷ���y��:������4���Qv���3��T񖻐����  �  o�=O;=��=d�=�1=[�=�~=G%=Z� =>q =� =0y�<6��<�<�Y�<Z��<���<�8�<���<���<��<�\�<��<a��<�/�<
t�<@��<C��<D:�<6z�<��<���<�3�<�o�<���<k��<�<�T�<��<׾�<s��<�!�<+P�<�{�<��<���<���<\�<�)�<B�<�V�<�g�<{t�<.}�<���<i��<�|�<�r�<�c�<MO�<�4�<p�<���<���<P��<�O�<`�<���<Qo�<T�<ų�<�J�<?��<�b�<���<&^�<���<?�<ॾ<��<ga�<T��<��<VO�<���<�Ҳ<�<RB�< s�<E��<�ǩ<��<��<s*�<-E�<<]�<�r�<m��<��<ݧ�<��<�<�͒<�א<�ߎ<��<��<7�<��<���<���<b��<<�}<��y<��u<+�q<��m<��i<��e<D�a<�]<�Y<]�U<��Q<��M<�I<�F<�B<�><�&:<�46<aE2<X.<Em*<��&<;�"<��<��<><;<on<��<0�<%-<�y <��;�P�;��;���;���;5��;���;���;n�;�a�;m��;W5�;�Ħ;o�;D5�;@�;y�;�6�;Cs�;ěy;6�n;ۻc;�%Y;��N;O�D;��:;01;ʎ';I;W7;Y;�;�h�:��:L��:��:�D�:�:6�:���:��v:b}Z:��>:`�#:9�:�s�9��9=�h9�>9��7A�����*�����sZ��'��"���p#���:�>R�b]i��*������N>�����������ú�'Ϻ�Vں�庇�����Y{�#
	�d����m���'��$�!*�R�/�a5��:���?��kE���J��WP��U�]K[�-�`��If���k��Pq���v�@[|�"���A����s��4���󋻫����p���.��햻߫���  �  ԓ=�;=$�=q�=u1=1�=�~=�$=�� =�p =S =�w�<���<��<2X�<٢�<6��<u7�<\��<���<��<\�<���<��<�/�<-t�<���<���<;�<G{�<>��<F��<95�<<q�<-��<���<��<�U�<��<��<���<�"�<�P�<n|�<"��<��<���<�<�(�<&A�<�U�<cf�<#s�<�{�<��<��<{�<Wq�<Pb�<�M�<�3�<��<���<[��<���<`O�<x�<���<�o�< �<���<�K�<���<d�<U��<�_�<���<�@�<���<%�<�b�<���<��<LP�<|��<mӲ<I�<bB�<�r�<鞫<�Ʃ<�<��<1)�<�C�<�[�<oq�<ᄜ<���<X��<���<S��<�̒<�֐<ߎ<e�<R�<
�<��<��<���<'��<9�}<	�y<&�u<��q<��m<�i<��e<��a<!�]<��Y< �U<R�Q<��M<��I<�F<1B<><P&:<M46<ZD2<uV.<gk*<.�&<��"<ʽ<��<
<�7<Lk<��<1�<`*<ow <��;�M�;��;���;��;a��;��;��;g�;�e�;�ó;J:�; ʦ;�t�;_;�;*�;��;5<�;�x�;@�y;��n;��c;�*Y;a�N;��D;y�:;�1;��';�C;,0;BQ;��;�R�:���:҈�:J��:�+�:���:{�:b��:�vv:^Z:5�>:A�#:6�:�a�9�9,�h9�{9��7%��7B*��P�����GH���6>#��:�R��0i�C��􁋺�ݖ�K0��mw��f���\�ú�'Ϻ�[ں���b���������	����,�p��24�M�$�E-*�+�/�	5���:�^�?�`rE�C�J�_ZP�a�U��J[��`�Ef�O�k��Hq���v�Q|��ꀻZ���8m���-��f틻����^k���)���薻�����  �  :�=�;=N�=�=h1=	�=]~=y$=^� =p =� =Vv�<*��<��<�V�<:��<���<6�<��<���<��<K[�<���<���<�/�<[t�<���<���<�;�<6|�<o��<���<�6�<�r�<���<���<0 �<xW�<J��<d��<���<�#�<�Q�<�|�<q��<��<r��<��<2(�<I@�<�T�<2e�<�q�<Nz�<�~�<T~�<�y�<�o�<�`�<�L�<�2�<t�<���<���<���<=O�<��<G��<Up�<��<���<M�<���<�e�<���<va�<,��<YB�<*��<�	�<Ld�<�<��<AQ�<7��<�Ӳ<��<kB�<�r�<o��<2Ʃ<&�<�
�<�'�<uB�<OZ�<�o�<X��<ꔚ<Ф�<*��<��<s˒<�Ր<Cގ<��<��<���<��<U��<��<���<�}<?�y<��u<��q<��m<(�i<��e<��a<D�]<��Y<��U<��Q<��M<X�I<�F<�B<G><!&:<�36<C2<�T.<Ii*<܀&<�"<�<f�<�<�4<�g<o�<G�<�'<u <���;(J�;��;~��;u��;���;��;#��;l!�;=i�;(ȳ;M?�;�Ϧ;�z�;+A�;$�;V$�;B�;�}�;"�y;a�n;��c;I0Y;D�N;��D; �:;#1;�';�=;�(;UH;�;�<�:���:No�:���:/�:�:��:bt�:BOv:�:Z:��>:ii#:s�:�T�9��9��h9��9���7'��M�)���������a���Y��#���:���Q�� i�q��Xn���Ζ��"��Am��ӱ����ú�(Ϻk_ں���9���������	�����7�V���@�(�$��9*�M�/��$5���:��@��xE���J�$]P�^�U�	J[�{�`�ZAf�!�k��Aq���v��F|��䀻.���/g���'��W狻�����e���$���㖻����  �  ��=<={�=��=Q1=��=~=&$=�� =�o = =�t�<ƿ�<l
�<"U�<���<_��<�4�<�~�<���<��<�Z�<q��<���<w/�<t�<W��<��<�<�<!}�<���<���<8�<%t�<+��<��<�!�<�X�<���<���<���<�$�<?R�<F}�<���<���<F��<#�<�'�<�?�<�S�<!d�<�p�<�x�<}�<�|�<x�<Sn�<�_�<TK�<|1�<q�<(��<(��<(��<O�<��<���<�p�<��<���<N�<.��<�f�<w��<�b�<���<�C�<���<:�<�e�<1��<��<R�<ו�<XԲ<��<\B�<tr�<���<�ũ<^�<�	�<�&�<"A�<�X�<_n�<ځ�<p��<h��<α�<���<_ʒ<�Ԑ<�ݎ<!�<��<���<��<���<x��<���<��}<]�y<�u<i�q<��m<�i< �e<��a<�]<��Y<�U<��Q<��M<� J<�F<�B<{><�%:<�26<�A2<�S.<ag*<�~&<\�"<,�<��<�<s1<�d<��<l�<.%<�r <Ҏ�;aG�;Z�;	��;���;���;F��;���;
$�;�l�;a̳;�C�;�Ԧ;��;�F�;*�;�)�;vG�;���;��y;�n;��c;�4Y;A�N;i�D;��:;k1;�';�8;�";�?;V�;�'�:Ԑ�:�W�:P|�:���:`̦:�:�^�:�,v:�Z:��>:eV#:~�:I�9��9� i9��9��7�V��MD)�̵��m\��\��o-���"��\:�4�Q���h�k��\��ڿ������d������J�ú�*Ϻcں�������� ���'	����xB�H���L�
�$��D*�(�/��.5�G�:��@�U~E�$�J�V`P���U��I[���`��=f�κk��:q�K�v�E=|��߀������a��c!���ዻ�]`������ߖ������  �  ݔ=]<=��=��=I1=��=�}=�#=�� =o =� =�s�<���<4	�<�S�<���<#��<�3�<�}�<���</�<Z�<	��<K��<q/�<�t�<���<���<N=�<�}�<|��<���</9�<cu�<k��<F��<�"�<Z�<���<���<}��<M%�<�R�<�}�<إ�<��< ��<��<'�<�>�<�R�<(c�<mo�<�w�<�{�<�{�<�v�<%m�<l^�<BJ�<�0�<��<t��<���<ۉ�<�N�<��<���<Qq�<+�<b��<O�<8��<�g�<���<Ed�<��<AE�<���<q�<�f�<2��<�	�<�R�<s��<�Բ< �<iB�<Gr�<���<ũ<��<��<�%�<@�<�W�<1m�<���<6��</��<���<���<fɒ<�Ӑ<�܎<��<A�<���<��<���<���<$��<G�}<%�y<&�u<��q<�m<��i<��e<�a<��]<��Y<5�U<��Q<F�M<�J<	F<B<�><�%:<z26<A2<R.<�e*<�|&<4�"<ε<��<0<�.<Rb<��<�<�"<�p <}��;jD�;q�;���;!��;���;*��;���;>&�;�o�;�ϳ;�G�;٦;���;|K�;�.�;a.�;�K�;���;E�y;��n;1�c;�8Y;��N;:�D;n�:;�1;�';f4;�;�8;M�;��:_}�:MD�:Th�:��: ��:�ݗ:IM�:�v:��Y:�i>:0D#:U�:=�9��9�i9�9/ �7]���v�(�x��[���C湵��"��4:�G�Q���h�(��OM��M���&��2\�������ú�*Ϻ�fں��9����H���/	����AL�����V���$��N*�|�/�075���:�@�&�E���J��bP���U�rI[�{�`��9f�>�k�v4q�-�v�!5|�Zۀ�⛃�~\������܋�%����[�����ܖ�q����  �  �=�<=��=��=<1=��=�}=�#=;� =�n =  =�r�<���<8�<�R�<���<)��<�2�<}�<��<��<�Y�<á�< ��<f/�<�t�<ٸ�<���<�=�<�~�<��<���<:�<Uv�<j��<;��<�#�<�Z�<|��<A��<��<�%�<+S�<~�<���<��<���<��<�&�<L>�<HR�<Zb�<�n�<�v�<�z�<�z�<�u�<)l�<~]�<yI�<�/�<�<���<A��<���<�N�<��<���<�q�<��<���<�O�<���<�h�<���<Te�<��<OF�<��<_�<�g�<껹<|
�<cS�<ݖ�<ղ<-�<sB�<
r�<p��<�ĩ<*�<<�<%�<A?�<�V�<9l�<��<:��</��<���<ڼ�<�Ȓ<)Ӑ<M܎<K�<��<p��<��<���<C��<���<q�}<W�y<��u<j�q<��m<��i<p�e<&�a<p�]<��Y<��U<��Q<��M<�J<�	F<�B<�><�%:<�16<o@2<Q.<�d*<E{&<��"<��<��<(�<�,<J`<�<H�<4!<Zo <"��;9B�;�;b��;���;0��;���;���;�'�;�q�;ҳ;�J�;Uܦ;E��;EO�;,2�;42�;8O�;��;��y;��n;O�c;�;Y;y�N;)�D;ּ:;1;�~'; 1;E;K4;��;��:Dn�:'4�:X�:xյ:㨦:7Η:Q@�:��u:��Y:�X>:�6#:�z:U-�9��9:!i9�79��7����(��J�� ߵ�c���
� �"�,:�vhQ��h����B������5���V��p�����ú.+Ϻ�kں�庽����\���6	���T�����^���$��V*���/��=5��:��@�Z�E���J��dP���U��H[��`�F7f���k��/q�i�v��.|��׀�6���yX������؋�o���eX������ٖ�����  �  ?�=�<=��=��=21=��=�}=e#=� =}n =� =gr�<���<��<AR�<���<���<42�<�|�<���<<�<CY�<���<���<W/�<�t�<���<��<#>�<�~�<���<,��<�:�<�v�<���<���<^$�<u[�<���<���<���<?&�<sS�<(~�<��<��<���<c�<u&�<�=�<�Q�<�a�<n�<Mv�<Vz�<z�<:u�<�k�<�\�<�H�<=/�<��<���<���<z��<�N�<��<��<�q�<��<f��<1P�<���<xi�</��<�e�<���<�F�<���<��</h�<r��<�
�<�S�<��<9ղ<>�<qB�<�q�<@��<cĩ<��<��<�$�<�>�<IV�<�k�<�<���<���</��<U��<'Ȓ<�Ґ<܎<�<��<[��<��<��<i��<���<;�}<T�y<��u<d�q<�m<��i<��e<?�a<��]<��Y<��U<��Q<V�M<�J<
F<�B<�><`%:<�16<�?2<�P.<�c*<Nz&<~�"<�<��<��<{+<_<˘<�<! <Pn <W��;A�; 
�;���;Z��;&��;3��;n��;6)�;Zs�;�ӳ;�L�;'ަ;=��;hQ�;�4�;?4�;?Q�;֋�;��y;��n;D�c;�=Y;��N;��D;d�:;)1;Q}';�.;c;g0;�~;- �:Se�:+�:�N�:7̵:ş�:aŗ:�7�:�u::�Y:�L>:�-#:Ct:D'�9��9,(i9iK9���7_���5O(�+��쿵�����
���"��:��WQ�>�h�X���:��¡��F���S�����G�ú�+Ϻ�lں��������K���:	�v��^X�q���c���$�[*��/��A5��:�2@���E���J��eP�U�U��H[�0�`�6f�|�k��,q�x�v��*|��Հ����PV��<��a֋�Q���rV������ז�p����  �  Q�='@=��=�=�5=z�=��=�(=�� =at = =Q�<���<a�<4b�<I��<���<�F�<6��<?��<+�<;v�<���<C
�<�R�<-��<���<�%�<�i�<o��<*��<�.�<un�<��<Z��<�&�<�a�<ƛ�<��<�
�<a?�<r�<\��<$��<���<�"�<�G�<�h�<Ά�<.��<���<���<���<���<���<j��<���<_��<���<&��<���<��<�s�<�I�<��<���<U��<�V�<]�<���<�L�<D��<�s�<���<�{�<l��<@f�<��<(5�<撽<+�<H;�<q��<�˶<��<�E�<�z�<���<S֭<��<��<�>�<�Y�<+r�<���<К�<���<I��<ɚ<h՘<x��<b�<�<���<� �<�<�	�<{�<��<�<3�<]�<d~<�
z<�v<��q<��m<=�i<��e<��a<��]<^�Y<�U<��Q<s�M<W�I<+�E<��A<��=<�9<��5<��1<]�-<X�)<Y�%<
"<�<�:<�Z<Y�<I�<��
<�<,X<�>�;���;��;gD�;B�;���;���;���;��;��;�N�;���;K�;���;�6�;D��;iϑ;�ǋ;�߅;��;��t;��i;��^;[GT;��I;��?;U�5;#,;��";pe;�Y;��;���:���:�x�:�l�:+��:�t�:���:��:���:J'g:>�K:=�0::`��9��9寐9�1<9T:�8��1�w�ڸ��N�즗� �ǹ1����	��_*�d�A��X�eo����F^�����;ڤ�&���9���fƺ��Ѻk�ܺ��續
�>/�����5
����D�����< �5�%��+�}�0���5�{K;��@��	F�jK�G�P��/V��[�va�urf�,�k��Zq�g�v��J|�l※J����\������Ջ�L���rM���	��ǖ�����  �  H�=@=��=�=�5=x�=͂=�(=�� =xt =) =��<��<��<�b�<���<���<0G�<r��<v��<*+�<Ev�<���<5
�<�R�<9��<s��<�%�<�i�<Y��<���<�.�<n�<���<��<t&�<�a�<a��<���<k
�<;?�<�q�<E��<��<���<�"�<�G�<
i�<��<<��<޷�<���<���<���<���<���<��<���<C��<u��<��<5��<t�<�I�<��<���<_��<�V�<7�<���<�L�<��<~s�<#��<Q{�<)��<�e�<���<�4�<|��<��<;�<P��<�˶<~�<�E�<�z�<
��<B֭<#��<��<�>�<Z�<_r�<���<'��<K��<���<_ɚ<�՘<���<��<H�<���<�<�<�	�<��<��<��<�<J�<S~<�
z<v<��q<��m<��i<;�e<�a<�]<��Y<��U<R�Q<\�M<.�I<��E<��A<��=<�9<��5<�1<y�-<��)<��%<�
"<� <H;<P[<�<��<W�
<�<�X<�?�;��;&��;�D�;�;5��;6��;,��;���;��;YN�;ס�;#�;6��;�5�;2�;-Α;�Ƌ;;ޅ;c�;��t;޼i;��^;�FT;�I;��?;��5;�",;5�";Bf;uZ;e�;i��:���:�~�:�q�:�Ƽ:z�:���:�:���:�,g:٨K:1�0:�:�9D��9D��9�1<9O�8�=2���ڸ�N�1����ǹb��L��i*���A�E�X��qo�����a��Ѣ��Uۤ�����;��kfƺ��ѺA�ܺ����	�.��\��54
�R���A����W: ���%�F+���0�_�5�4J;�ҩ@�1	F�0iK�(�P��/V���[��a�Lsf���k�9[q���v�M|��〻�����]��2���֋������N���
���ǖ�G����  �  	�=�?=��=�=�5=��=��=)=� =�t =} =e��<���<|�<Zc�<_��<���<�G�<��<��<�+�<�v�<��<\
�<�R�<$��<H��<I%�<i�<ë�<c��<�-�<gm�<��<I��<�%�<�`�<���<��<�	�<�>�<rq�<��<���<���<�"�<�G�<Li�<J��<���<~��<`��<���<���<���<���<���<d��<���<%��<|��<ӗ�<�t�<TJ�<��<���<T��<�V�<��<.��<TL�<x��<�r�<|��<�z�<l��<e�<���<!4�<���</�<k:�<���<0˶<"�<�E�<�z�<	��<]֭<s��<& �<"?�<�Z�<�r�<���<ܛ�<��<j��<*ʚ<p֘<��<T�<��<d��<��<��<&
�<��<��<��<��<�
�<5~<e	z<�v<��q<m�m<D�i<��e<��a<��]<Q�Y<Z�U<!�Q</�M<-�I<m�E<}�A<��=<%�9<��5<��1<d�-<��)<��%<�"<"<�<<�\<��<��<��
<<�Y<oB�;f��;��;}F�;��;���;��;���;���;��;/L�;���;��;���;3�;5�;ˑ;.ċ;�ۅ;�;��t;R�i;��^;�CT;��I;ҿ?;��5;�#,;t�";�i;]^;��;���:���:/��:&}�:�Ӽ:@��:O��:���:��:�@g:a�K:v�0:�:ª�9���9���9�#<9J�8�5�}Q۸$O��ڗ���ǹ:<��='���*�j�A���X��o�!���j��C���[㤺����>���gƺ�Ѻ��ܺY���%��A��N/
����8<�����3 �1�%��+��}0� �5�1E;� �@�tF�fK�v�P�C/V��[�a�,uf�{�k��_q���v��Q|�`总�����`������ً�����wQ��-��ʖ������  �  Ɨ=�?=z�=܎=�5=��=1�=k)=h� =Fu = =���<'��<��<�d�<���<���<I�<+��< ��<s,�<Yw�<o��<�
�<�R�<��<��<�$�<�h�<��<u��<�,�<4l�<���<���<c$�<}_�<x��<���<��<�=�<�p�<^��<x��<���<�"�<H�<�i�<Ӈ�<l��<F��<q��<���<���<��<���<-��<���<;��<?��<���<���<3u�<�J�<;�<:��<?��<lV�<��<���<�K�<���<�q�<9��<Ly�<���<�c�<���<�2�<w��<��<^9�<Մ�<�ʶ<�
�<CE�<�z�<���<�֭<���<� �<�?�<t[�<t�<ʉ�<)��<\��<���<{˚<�ט<��<t�<���<)��<:�<��<�
�<��<��<��<y�<O
�<�~<�z<��u<J�q<��m<��i<�e<��a<��]<��Y<�U<]�Q<��M<�I<�E<�A<��=<r�9<��5<��1<��-<K�)<��%<1"<�$<�?<�_<r�<T�<��
<�<R\<VF�;���;��;6H�;��;"��;���;��;��;��;vI�;J��;��;��;.�;H�;OƑ;�;�օ;��;��t;U�i;��^;@T;=�I;ľ?;��5;�&,;1�";n;bd;�;��:'�:���:s��:�:���:p��:g
�:(��:�cg:N�K:�0:	#:ν�93��9Ⱀ9u<9��8*9���۸�O�E���
ȹ5��� S���*�r�A���X��o�1��~z��]���r줺����B��	jƺ��Ѻ�ܺ5�������X���&
�n���1�1��=) ���%��
+�
t0��5�=;��@���E��bK���P��-V���[��a�jxf���k�Leq�$�v�sZ|�(뀻����f���"��
ߋ�����?V������͖�q����  �  d�=p?=U�=׎=
6=��=��=�)=�� =�u =� =��<���<��<jf�<f��<z��<�J�<���<A��<|-�<7x�<���<�<�R�<��<���<$�<�g�<��<9��<i+�<�j�<��<\��<�"�<�]�<��<o��<�<�<�<�o�<���<���<��<�"�<9H�<j�<���<f��<g��<���<	��<o��<���<���<���<]��<���<���<ڶ�<���<&v�<�K�<��<e��<,��<6V�< �<ǫ�<�J�<a��<fp�<���<�w�<=��<�a�<���< 1�<���<e�<8�<���<�ɶ<�	�<�D�<kz�<�<�֭<+��<!�<�@�<�\�<^u�</��<���<��<r��<+͚<g٘<@�<��<B��<B��<2�<��<�
�<��<��<o�<��<�	�<�~<Oz<�u<^�q<��m<8�i<��e<��a<��]<��Y<F�U<��Q<��M<x�I<)�E<b�A<`�=<��9<y�5<��1<��-<q�)<��%<"<�'<�B<'c<�<״<��
<�<C_<�K�;%��;�;�J�;e�;���;���;���;���;�
�;fE�;���;W�;���;(�;�;���;���;#х;�;νt;��i;��^;�:T;!�I;Ͻ?;��5;�(,;A�";ot;�l;a�;���:�#�:>��:��:��:4��:�Þ:�"�:�ρ:ǎg:�K:8�0:|<:	��9U��9���9�;9��8m�>���ܸ�P�n���gȹi�����R�*�mB��
Y��o��G��Z���Pʙ�����&���I��qkƺ,�ѺU�ܺ��纠��	�����n
����%�Ԣ�X ��%���*�Mh0���5��2;�P�@�d�E�/]K�P�P�a,V���[��a�Q}f���k��mq���v�1e|�����®���l��$)���勻Ϡ��\����jҖ������  �  �=$?=�=Î=!6=,�=�=U*=�� =�v =� =��<���<z�<ah�<X��<Z �<dL�< ��<���<�.�<y�<���<r�<S�<���<&��<~#�<�f�<���<���<�)�<�h�<&��<h��<� �<\�<��<���<��<O;�<�n�<؟�<Y��<��<�"�<tH�<�j�<O��<^��<»�<3��<���<M��<���<���<���<B��<���<m��<H��<��<w�<KL�<G�<���<��<�U�<]�<���<eI�<���<�n�<���<�u�<E��<�_�<���<�.�<܌�<��<n6�<3��<eȶ<��<D�<z�<�<"׭<���<:"�<�A�<�]�<�v�<��<���<�<g��<$Ϛ<Pۘ<&�<��<���<���<&�<t�<�<1�<��<�<M�<��<n
~<�z<��u<��q<��m<l�i<��e<��a<��]<9�Y<�U<��Q<�M<v�I<��E<`�A<�=<��9<`�5<\�1<k�-<��)<q&<m"<k+<�F<7g<#�<�<��
<�#<�b<�Q�;L��;���;<N�;]�;���;f��;F��;���;H�;�@�;[��;f��;���;� �;�ݗ;/��;���;�Ʌ;��;=�t;H�i;4�^;�4T;@�I;=�?;D�5;�*,;��";�z;�t;��;��:QA�:���:���:%�:�ح:��:*A�:��:M�g:�)L: 1:�T:t	�9"�9���9��;9 ��8v�D���ݸh�P�,Θ���ȹ1d�����!+�LB�rFY��p�Na�������ޙ�0��e0��6R��pƺ��Ѻߧܺ�级��q���S��<
����$�C��� �/%�|�*�)Y0�=�5�R';�׋@���E�WK�$�P��*V�ݙ[�7a���f���k��vq���v��q|����}���4t��K1��:틻����Cc��S��ؖ�v����  �  ^�=�>=��=��=76=a�=H�=�*=?� =aw =p =ֆ�<���<��<wj�<���<Z�<?N�<Ι�<"��<�/�<z�<r��<��<?S�<���<���<�"�<�e�<j��<!��<(�<�f�<��<R��<��<�Y�<��<���<4�<�9�<�m�<מ�<���<���<�"�<�H�<7k�<4��<���<&��<���<���<2��<���<���<���<\��<w��<2��<׹�<p��<Cx�<(M�<��<���<��<WU�<��<��<!H�<y��<�l�< ��<�s�<��<�]�<m��<�,�<ˊ�<��<�4�<ʀ�<!Ƕ<�<rC�<�y�<���<[׭<c��<#�<
C�<`_�<lx�<͎�<x��<��<uÜ<Bњ<dݘ<�<V�<@��<���<9�<N	�<��<j�<��<��<�
�<��<~<��y<f�u<&�q<��m<D�i<1�e<x�a<��]<w�Y<o�U<½Q<��M<;�I<^�E<a�A<��=<L�9</�5<��1<x�-<��)<�&<�"<H/<�J<�k<u�<^�<�
<g'<+f<X�;���;��;�Q�;<�;���;��;���;���;I�;Q<�;4��;���;cy�;�;�՗;��;ة�;(;��;ɤt;Ҕi;{�^;~-T;��I;��?;��5;C-,;V�";U�;J~;�;W*�:^�:���:/��:�F�:���:b�:c`�:�
�:��g:�WL:�.1:�r: .�9z �9+��9Z�;9�8�rL�<#߸_pQ��=��Bɹ������Qe+�
�B�F�Y�EWp��}������B�T��)>���Z���sƺ��Ѻ¢ܺj�纁��#����z�
�L��T������(n%���*�J0�8�5��;�Հ@���E�ePK�u�P�.)V�H�[��a�x�f�kl�b�q���v��|�L�������k|���9����������j��p$��Aޖ�B����  �  ݕ=c>=��=��=G6=��=��=c+=�� =*x =T =���<���<� �<�l�<���<]�<P�<���<���<$1�<{�<��<5�<GS�<I��<*��<�!�<qd�<��<���<I&�<e�<��<3��<|�<�W�<��<!��<��<v8�<Fl�<��<��<l��<�"�<�H�<�k�<��<���<o��<v��<\��<��<���<���<���<b��<e��<���<���<���<[y�<N�<E�<��<��<�T�<��<٨�<�F�<���<-k�<��<rq�<���<W[�<0��<�*�<���<��<�2�<D�<�Ŷ<��<�B�<Sy�<ת�<�׭<���<$�<"D�<�`�<#z�<���<o��<��<�Ŝ<VӚ<kߘ<��<!�<���<:�<Z�<
�<~�<��<��<?�<�	�<��<u~<��y<��u<f�q<��m<��i<��e<�a<��]<��Y<�U<��Q<ȺM< �I<��E<��A<c�=<�9<�5<m�1<��-<-�)<�&<�"<3<O<�o<�<��<@�
<;+<�i<_^�;��;���;�T�;a�;f��;���;L��;���;r��;?7�;m��;�;Dr�;*�;�͗;*��;���;���;��;s�t;͉i;�^;�&T;L�I;Ѷ?;��5;�/,;�";ȉ;ɇ;Ǻ;9F�:;{�:E�:��:�h�:��:�&�:��:'�:�)h:e�L:1T1:А:�R�9�5�9)��9"�;9�Y�8��S�J\��'R�ߤ����ɹ_��\H�|�+�A�B���Y��p�����َ��	��~/��bL���b���wƺˊѺ��ܺY��2��b���?o���	��v�T���q����v]%���*�;0���5��;�w@���E�JK���P��'V�q�[��a�R�f�Gl��q��w�T�|�����ƃ����,B���������!r��Y+��T䖻�����  �  k�=>=r�=��=]6=��=��=�+=u� =�x = =���<���<�"�<�n�<k��<L�<�Q�<��<���<M2�<�{�<���<��<^S�<��<���<!�<~c�<���<&��<�$�<4c�<��<4��<��<�U�<-��<B��<�<7�<)k�<��<\��<��<�"�<@I�<Il�<���<���<���<���<���<���<���<���<���<4��<E��<���<���<���<^z�<�N�<��<E��<͞�<�T�<5�<���<�E�<k��<�i�<��<so�<���<6Y�<��<�(�<���<�޻<T1�<�}�<�Ķ<"�<B�<�x�<Ǫ�<�׭<e �<�$�<0E�<b�<�{�<7��<S��<淞<�ǜ<B՚<S�<��<���<W��<{�<c�<�
�<�<��<a�<��<-	�<��<~<��y<��u<��q<��m<��i<��e<�a<��]<ºY<��U<ɷQ<9�M<E�I<(�E<��A<��=<��9<�5<��1<��-<��)<�
&<�"<�6<S<�s<�<��<J�
<�.<5m<Nd�;)��;���;nW�;��;3��;W��;���;U��;��;[2�;'��;��;k�;�	�;Ɨ;���;.��;���;]�;�t;.i;��^;� T;�I;��?;X�5;�2,;��";~�;t�;m�;O^�:���:3�:�.�:8��:�<�:gD�:۞�:{A�:�Yh:߬L:�v1:��:�u�9�J�98��9=`;9'��8�Y��h�D�R�����-ʹ
�������+�dC��Z�]�p���������?���>��KX��|l��E{ƺ'�Ѻ"�ܺq��=��l���\d���	�Fi�����b����N%�X�*�=,0�Q�5�t;�"m@���E�-EK��P�&V���[��a�\�f� l�z�q�w��|�N��΃�،��	J�����T����y���1���閻�����  �  ��=�==C�=}�=d6=�=H�=F,=�� =}y =� =���<5��<>$�<Mp�<��<��<@S�<t��</��<Q3�<�|�<J��<��<eS�<��<3��<a �<�b�<���<���<'#�<�a�<|��<���<��<1T�<���<���<���<�5�<%j�<D��<���<���<�"�<XI�<�l�<v��<���<���<)��<`��<y��<��<B��<���<���<���<���<3��<��<A{�<[O�<2�<U��<���<IT�<��<��<�D�<"��<!h�<���<�m�<���<aW�<=��<�&�< ��<jݻ<�/�<�|�<�ö<L�<�A�<�x�<���<ح<� �<o%�<F�<%c�<�|�<���<է�<���<>ɜ<�֚<��<=�<��<���<��<<�<u�<g�<��<O�<��<��<��<� ~<:�y<��u<��q<��m<��i<j�e<��a<y�]<зY<��U<$�Q<
�M<c�I<�E<��A<��=<��9<��5<��1<7�-<��)< &<�!"<�9<EV<>w<��<��<��
<�1<	p<xi�;� �;ܥ�;9Z�;��;���;��;D��;���;���;\.�;I|�;Y�;�e�;��;���;���;ד�;���;}�;��t;�ui; �^;�T;H�I;ز?;��5;�3,;��";��;�;��;�r�:¬�:<K�:�H�:���:XW�:l^�::��:�X�:��h:h�L:��1:K�:���9S�9��9�@;9k'�8?m`�i�orS�0Z��3�ʹ�8��Ϻ��,��HC�=Z�y q�̓�%��"1��N��d���s��E~ƺ�Ѻ�ܺ��c�򺛮���Z�7�	��]�����U�?���@%�Ա*�� 0�>�5���:�\d@���E��?K���P��%V�G�[�wa��f�/l�ܜq�%!w�1�|���xԃ�����Q������Ǝ�y��z7��Ϧ���  �  ��=�==�=k�=t6=!�=��=�,=[� =�y =]  ='��<{��<�%�<�q�<i��<	�<sT�<���<��<4�<7}�<���<�<{S�<���<���<��<�a�<٢�<���<	"�<y`�<��</��<r�<�R�<O��<���<���<�4�<ji�<���<���<t��<�"�<|I�<�l�<��<)��<���<#��<���<���<w��<���<���<$��<���<��</��<Ѡ�<�{�<�O�<q�<p��<���<�S�<C�<q��<�C�<>��<�f�<[��<ql�<���<�U�<���<O%�<ǃ�<6ܻ<�.�<�{�<�¶<��<&A�<\x�<���<,ح<6�<�%�<�F�<�c�<�}�<ʔ�<��<ݺ�<{ʜ<.ؚ<1�<q�<G��<���<Y�<��<��<��<�<<�<+�<A�<I�<��}<`�y<��u<X�q<�m<��i<��e<��a<��]<\�Y<k�U<(�Q<~�M< �I<
�E<��A<f�=<�9<�5<��1<G�-<C�)<�&<�#"<9<<�X<�y<�<��<�
<{4<Xr<m�;��;=��;\�;��;W��;t��;%��;Z��;)��;�+�;hx�;'ߪ;�`�;���;���;�;���;���;��;,zt;�oi;��^;�T;+�I;S�?;��5;E5,;	�";��;͜;��;҂�:���:i^�:}^�:��:�k�:yt�:Dʐ:�k�:*�h:g�L:��1:~�:z��92]�9�9;9�ܫ8l"e��#��S����F�ʹ��������H,�sC�iZ��(q��ރ�6���=���Y��gl���x��ÂƺވѺR�ܺS����֣��zT���	�(T�����J�B���6%�]�*��0���5�Y�:�h^@���E��;K�ȮP��$V���[��a��f�bl�ɢq��(w���|�����ك�����MV����̎�G����;����ͩ���  �  h�=S==��=e�={6=3�=��=�,=�� =7z =�  =э�<5��<P&�<`r�<"��<�	�<U�<��<���<�4�<�}�<���<2�<�S�<���<���<��<_a�<=��<.��<Z!�<�_�<g��<a��<��<R�<���<���<���<Z4�<�h�<;��<0��<O��<�"�<�I�</m�<C��<���<.��<���<"��<U��<'��<P��<���<���<���<���<���<e��<V|�<!P�<��<���<���<�S�<� �<���<7C�<���<Lf�<���<�k�<���<U�<���<�$�<��<wۻ<.�<{�<b¶<C�<�@�<7x�<���<Dح<a�<F&�<AG�<{d�<v~�<c��<���<���<J˜<�ؚ<��<�<���<��<��<I	�<:�<��<*�<3�<�<��<��<f�}<�y<��u<��q<��m<I�i<�e<f�a<B�]<ݳY<�U<߱Q<O�M<�I<J�E<��A<I�=<4�9<^�5<T�1<B�-<n�)<&<%"<�=<bZ<�{<ס<C�<��
<�5<�s<�o�;�;3��;$]�;��;���;Q��;m��;���;o��;Q)�;v�;�ܪ;^�;���;w��;ӑ�;Ջ�;ѥ�;b�;�ut;�ji;ҟ^;�T;��I;c�?;��5;!6,;��";h�;��;��;<��:���:�i�:�i�:%Ž:�x�:��:�Ր:�u�:��h:��L:Z�1:d�:S��9�c�9ð�9�;9a��8�^h����,T��ǚ���ʹ۹�����c,��C��Z��?q�
ꃺ$!���G���a���r���|��Z�ƺ9�Ѻ7�ܺ�纜��=����O�"�	�7O�A��%E����W0%���*��0�T5���:��Y@���E��9K���P��#V�Z�[��a�ǝf��!l�8�q��-w�	�|�����܃�����Y�����Ύ�6���z>��b�������  �  a�=E==��=b�=s6==�=��=�,=�� =Oz =�  =+��<���<�&�<�r�<`��<(
�<nU�<`��<���<�4�<�}�<��<@�<tS�<���<���<k�<Ra�<��<��<!�<i_�<��<��<N�<�Q�<=��<���<���<#4�<�h�<.��<��<\��<�"�<�I�<Qm�<]��<���<L��<���<w��<���<f��<���<���<��<��<��<���<���<_|�<6P�<��<}��<���<�S�<� �<��<"C�<T��<f�<D��<Mk�<m��<�T�<���<7$�<���<&ۻ<�-�<�z�<P¶<&�<�@�<7x�<���<Hح<~�<Z&�<FG�<�d�<�~�<���<��<ͻ�<�˜<8ٚ<3�<|�<)��<H��<�<]	�<Y�<��<�<)�<�<��<��<2�}<��y<�u<'�q<��m<��i<j�e<��a<��]<%�Y<��U<z�Q<�M<��I<�E<��A<=�=<�9<��5<��1<j�-<��)<v&<�%"<M><
[<|<{�<��<]�
<�6<t<Kp�;8�;���;�]�;��;z��;\��;W��;���;L��;�(�;�u�;�۪;�\�;���;5��;���;���;x��;ʽ;tt;ii;P�^;�T;��I;ٯ?;\�5;�5,;��";F�;��;��;��:��:Jp�:�m�:�ɽ:�}�:o��:,ܐ:{�:�h:�M:ʺ1:O�:;��9c�9n��9�	;9ur�8O�h�r���GT��Қ��˹�����m,�ΗC�щZ��Jq���#��J��fb��9t���}���ƺF�Ѻܺ��+�򺳚��~N��	�^L�$��.C�)��%.%�R�*��0��|5�$�:�-Y@��E��8K���P�S$V���[�ja���f�<"l��q�H/w���|���	ރ�T����Z��r��CЎ�����}?��%��������  �  h�=S==��=e�={6=3�=��=�,=�� =7z =�  =э�<5��<P&�<`r�<"��<�	�<U�<��<���<�4�<�}�<���<2�<�S�<���<���<��<_a�<=��<.��<Z!�<�_�<g��<a��<��<R�<���<���<���<Z4�<�h�<;��<0��<O��<�"�<�I�</m�<C��<���<.��<���<"��<U��<'��<P��<���<���<���<���<���<e��<V|�<!P�<��<���<���<�S�<� �<���<7C�<���<Lf�<���<�k�<���<U�<���<�$�<��<wۻ<.�<{�<b¶<C�<�@�<7x�<���<Dح<a�<F&�<AG�<{d�<v~�<c��<���<���<J˜<�ؚ<��<�<���<��<��<I	�<:�<��<*�<2�<�<��<��<f�}<�y<��u<��q<��m<I�i<�e<f�a<B�]<ݳY<�U<߱Q<O�M<�I<J�E<��A<I�=<4�9<^�5<T�1<C�-<n�)<&<%"<�=<bZ<�{<ס<C�<��
<�5<�s<�o�;�;3��;$]�;��;���;P��;m��;���;o��;Q)�;v�;�ܪ;^�;���;w��;ӑ�;Ջ�;ѥ�;b�;�ut;�ji;ҟ^;�T;��I;c�?;��5;!6,;��";h�;��;��;<��:���:�i�:�i�:%Ž:�x�:��:�Ր:�u�:��h:��L:Z�1:d�:S��9�c�9ð�9�;9a��8�^h����,T��ǚ���ʹ۹�����c,��C��Z��?q�
ꃺ$!���G���a���r���|��Z�ƺ9�Ѻ7�ܺ�纜��=����O�"�	�7O�A��%E����W0%���*��0�T5���:��Y@���E��9K���P��#V�Z�[��a�ǝf��!l�8�q��-w�	�|�����܃�����Y�����Ύ�6���z>��b�������  �  ��=�==�=k�=t6=!�=��=�,=[� =�y =]  ='��<{��<�%�<�q�<i��<	�<sT�<���<��<4�<7}�<���<�<{S�<���<���<��<�a�<٢�<���<	"�<y`�<��</��<r�<�R�<O��<���<���<�4�<ji�<���<���<t��<�"�<|I�<�l�<��<)��<���<#��<���<���<w��<���<���<$��<���<��</��<Ѡ�<�{�<�O�<q�<p��<���<�S�<C�<q��<�C�<>��<�f�<[��<ql�<���<�U�<���<O%�<ǃ�<6ܻ<�.�<�{�<�¶<��<&A�<\x�<���<,ح<6�<�%�<�F�<�c�<�}�<ʔ�<��<ݺ�<{ʜ<.ؚ<1�<q�<G��<���<Y�<��<��<��<�<<�<+�<A�<I�<��}<`�y<��u<X�q<�m<��i<��e<��a<��]<\�Y<k�U<(�Q<~�M< �I<�E<��A<f�=<�9<�5<��1<G�-<C�)<�&<�#"<9<<�X<�y<�<��<�
<{4<Xr<m�;��;=��;\�;��;V��;t��;%��;Y��;)��;�+�;hx�;'ߪ;�`�;���;���;�;���;���;��;,zt;�oi;��^;�T;+�I;S�?;��5;E5,;	�";��;͜;��;т�:���:i^�:}^�:��:�k�:yt�:Dʐ:�k�:*�h:g�L:��1:~�:z��92]�9�9;9�ܫ8l"e��#��S����F�ʹ��������H,�sC�iZ��(q��ރ�6���=���Y��gl���x��ÂƺވѺR�ܺS����֣��zT���	�(T�����J�B���6%�]�*��0���5�Y�:�h^@���E��;K�ȮP��$V���[��a��f�bl�ɢq��(w���|�����ك�����MV����̎�G����;����ͩ���  �  ��=�==C�=}�=d6=�=H�=F,=�� =}y =� =���<5��<>$�<Mp�<��<��<@S�<t��</��<Q3�<�|�<J��<��<eS�<��<3��<a �<�b�<���<���<'#�<�a�<|��<���<��<1T�<���<���<���<�5�<%j�<D��<���<���<�"�<XI�<�l�<v��<���<���<)��<`��<y��<��<B��<���<���<���<���<3��<��<A{�<[O�<2�<U��<���<IT�<��<��<�D�<"��<!h�<���<�m�<���<aW�<=��<�&�< ��<jݻ<�/�<�|�<�ö<L�<�A�<�x�<���<ح<� �<o%�<F�<%c�<�|�<���<է�<���<>ɜ<�֚<��<=�<��<���<��<<�<u�<g�<��<O�<��<��<��<� ~<:�y<��u<��q<��m<��i<j�e<��a<y�]<зY<��U<$�Q<
�M<c�I<�E<��A<��=<��9<��5<��1<7�-<��)< &<�!"<�9<EV<>w<��<��<��
<�1<	p<xi�;� �;ܥ�;9Z�;��;���;��;D��;���;���;\.�;H|�;Y�;�e�;��;���;���;ד�;���;|�;��t;�ui; �^;�T;H�I;ز?;��5;�3,;��";��;�;��;�r�:¬�:<K�:�H�:���:XW�:l^�::��:�X�:��h:h�L:��1:K�:���9S�9��9�@;9k'�8?m`�i�orS�0Z��3�ʹ�8��Ϻ��,��HC�=Z�y q�̓�%��"1��N��d���s��E~ƺ�Ѻ�ܺ��c�򺛮���Z�7�	��]�����U�?���@%�Ա*�� 0�>�5���:�\d@���E��?K���P��%V�G�[�wa��f�/l�ܜq�%!w�1�|���xԃ�����Q������Ǝ�y��z7��Ϧ���  �  k�=>=r�=��=]6=��=��=�+=u� =�x = =���<���<�"�<�n�<k��<L�<�Q�<��<���<M2�<�{�<���<��<^S�<��<���<!�<~c�<���<&��<�$�<4c�<��<4��<��<�U�<-��<B��<�<7�<)k�<��<\��<��<�"�<@I�<Il�<���<���<���<���<���<���<���<���<���<4��<E��<���<���<���<^z�<�N�<��<E��<͞�<�T�<5�<���<�E�<k��<�i�<��<so�<���<6Y�<��<�(�<���<�޻<T1�<�}�<�Ķ<"�<B�<�x�<Ȫ�<�׭<e �<�$�<0E�<b�<�{�<7��<S��<淞<�ǜ<B՚<S�<��<���<W��<z�<c�<�
�<�<��<a�<��<-	�<��<~<��y<��u<��q<��m<��i<��e<�a<��]<ºY<��U<ɷQ<9�M<F�I<)�E<��A<��=<��9<�5<��1<��-<��)<�
&<�"<�6<S<�s<�<��<J�
<�.<5m<Md�;)��;���;nW�;��;2��;W��;���;U��;��;Z2�;'��;��;k�;�	�;Ɨ;���;.��;���;\�;�t;-i;��^;� T;�I;��?;X�5;�2,;��";~�;t�;m�;O^�:���:3�:�.�:8��:�<�:gD�:۞�:{A�:�Yh:߬L:�v1:��:�u�9�J�98��9=`;9'��8�Y��h�D�R�����-ʹ
�������+�dC��Z�]�p���������?���>��KX��|l��E{ƺ'�Ѻ"�ܺq��=��l���\d���	�Fi�����b����N%�X�*�=,0�Q�5�t;�"m@���E�-EK��P�&V���[��a�\�f� l�z�q�w��|�N��΃�،��	J�����T����y���1���閻�����  �  ݕ=c>=��=��=G6=��=��=c+=�� =*x =T =���<���<� �<�l�<���<]�<P�<���<���<$1�<{�<��<5�<GS�<I��<*��<�!�<qd�<��<���<I&�<e�<��<3��<|�<�W�<��<!��<��<v8�<Fl�<��<��<l��<�"�<�H�<�k�<��<���<o��<v��<\��<��<���<���<���<b��<e��<���<���<���<[y�<N�<E�<��<��<�T�<��<٨�<�F�<���<.k�<��<rq�<���<W[�<0��<�*�<���<��<�2�<D�<�Ŷ<��<�B�<Sy�<ת�<�׭<���<$�<"D�<�`�<#z�<���<o��<��<�Ŝ<VӚ<kߘ<��<!�<���<:�<Z�<
�<~�<��<��<>�<�	�<��<u~<��y<��u<f�q<��m<��i<��e<�a<��]<��Y<�U<��Q<ɺM< �I<��E<��A<c�=<�9<�5<m�1<��-<-�)<�&<�"<3<O<�o<�<��<@�
<;+<�i<^^�;��;���;�T�;`�;f��;���;K��;���;r��;?7�;m��;�;Cr�;)�;�͗;)��;���;���;��;s�t;̉i;�^;�&T;L�I;Ѷ?;��5;�/,;�";ȉ;ȇ;Ǻ;9F�:;{�:E�:��:�h�:��:�&�:��:'�:�)h:e�L:1T1:А:�R�9�5�9)��9"�;9�Y�8��S�J\��'R�ߤ����ɹ_��\H�|�+�A�B���Y��p�����َ��	��~/��bL���b���wƺˊѺ��ܺY��2��b���?o���	��v�T���q����v]%���*�;0���5��;�w@���E�JK���P��'V�q�[��a�R�f�Gl��q��w�T�|�����ƃ����,B���������!r��Y+��T䖻�����  �  ^�=�>=��=��=76=a�=H�=�*=?� =aw =p =ֆ�<���<��<wj�<���<Z�<?N�<Ι�<"��<�/�<z�<r��<��<?S�<���<���<�"�<�e�<j��<!��<(�<�f�<��<R��<��<�Y�<��<���<4�<�9�<�m�<מ�<���<���<�"�<�H�<7k�<4��<���<&��<���<���<2��<���<���<���<\��<w��<2��<׹�<p��<Cx�<(M�<��<���<��<WU�<��<��<!H�<z��<�l�< ��<�s�<��<�]�<m��<�,�<ˊ�<��<�4�<ʀ�<"Ƕ<�<rC�<�y�<���<[׭<c��<#�<
C�<`_�<lx�<͎�<x��<��<uÜ<Bњ<dݘ<�<V�<?��<���<9�<N	�<��<j�<��<��<�
�<��<~<��y<f�u<%�q<��m<D�i<1�e<x�a<��]<w�Y<o�U<½Q<��M<;�I<_�E<b�A<��=<L�9</�5<��1<x�-<��)<�&<�"<H/<�J<�k<u�<^�<�
<g'<+f<X�;���;��;�Q�;;�;���;��;���;���;H�;P<�;3��;���;by�;�;�՗;��;ة�;(;��;Ȥt;єi;{�^;}-T;��I;��?;��5;C-,;U�";U�;J~;�;V*�:^�:���:/��:�F�:���:b�:c`�:�
�:��g:�WL:�.1:�r: .�9z �9+��9Z�;9�8�rL�<#߸_pQ��=��Bɹ������Qe+�
�B�F�Y�EWp��}������B�T��)>���Z���sƺ��Ѻ¢ܺj�纁��#����z�
�L��T������(n%���*�J0�8�5��;�Հ@���E�ePK�u�P�.)V�H�[��a�x�f�kl�b�q���v��|�L�������k|���9����������j��p$��Aޖ�B����  �  �=$?=�=Î=!6=,�=�=U*=�� =�v =� =��<���<z�<ah�<X��<Z �<dL�< ��<���<�.�<y�<���<r�<S�<���<&��<~#�<�f�<���<���<�)�<�h�<&��<h��<� �<\�<��<���<��<O;�<�n�<؟�<Y��<��<�"�<tH�<�j�<O��<^��<»�<3��<���<M��<���<���<���<B��<���<m��<H��<��<w�<KL�<G�<���<��<�U�<]�<���<eI�<���<�n�<���<�u�<E��<�_�<���<�.�<܌�<��<n6�<3��<eȶ<��<D�<z�<�<"׭<���<;"�<�A�<�]�<�v�<��<���<�<g��<$Ϛ<Pۘ<&�<��<���<���<%�<t�<�<1�<��<�<M�<��<n
~<�z<��u<��q<��m<l�i<��e<��a<��]<:�Y<�U<��Q<	�M<v�I<��E<a�A<�=<��9<`�5<\�1<k�-<��)<q&<m"<k+<�F<7g<#�<�<��
<�#<�b<�Q�;L��;���;;N�;]�;���;f��;F��;���;H�;�@�;[��;e��;���;� �;�ݗ;/��;���;�Ʌ;��;<�t;G�i;3�^;�4T;?�I;=�?;D�5;�*,;��";�z;�t;��;��:QA�:���:���:%�:�ح:��:*A�:��:M�g:�)L: 1:�T:t	�9"�9���9��;9 ��8w�D���ݸh�P�,Θ���ȹ1d�����!+�LB�rFY��p�Na�������ޙ�0��e0��6R��pƺ��Ѻߧܺ�级��q���S��<
����$�C��� �/%�|�*�)Y0�=�5�R';�׋@���E�WK�$�P��*V�ݙ[�7a���f���k��vq���v��q|����}���4t��K1��:틻����Cc��S��ؖ�v����  �  d�=p?=U�=׎=
6=��=��=�)=�� =�u =� =��<���<��<jf�<f��<z��<�J�<���<A��<|-�<7x�<���<�<�R�<��<���<$�<�g�<��<9��<i+�<�j�<��<\��<�"�<�]�<��<o��<�<�<�<�o�<���<���<��<�"�<9H�<j�<���<f��<g��<���<	��<o��<���<���<���<]��<���<���<ڶ�<���<&v�<�K�<��<e��<,��<6V�< �<ǫ�<�J�<a��<fp�<���<�w�<=��<�a�<���< 1�<Ꮍ<e�<8�<���<�ɶ<�	�<�D�<kz�<�<�֭<+��<!�<�@�<�\�<^u�</��<���<��<r��<+͚<g٘<@�<��<A��<B��<2�<��<�
�<��<��<o�<��<�	�<�~<Oz<�u<^�q<��m<8�i<��e<��a<��]<��Y<F�U<��Q<��M<y�I<)�E<b�A<`�=<��9<z�5<��1<��-<q�)<��%<"<�'<�B<'c<�<״<��
<�<C_<�K�;$��;�;�J�;d�;���;���;���;���;�
�;eE�;���;W�;���;(�;�;���;���;#х;�;νt;��i;��^;�:T;!�I;Ͻ?;��5;�(,;A�";ot;�l;a�;���:�#�:>��:��:��:4��:�Þ:�"�:�ρ:ǎg:�K:8�0:|<:	��9U��9���9�;9��8m�>���ܸ�P�n���gȹi�����R�*�mB��
Y��o��G��Z���Pʙ�����&���I��qkƺ,�ѺU�ܺ��纠��	�����n
����%�Ԣ�X ��%���*�Mh0���5��2;�P�@�d�E�/]K�P�P�a,V���[��a�Q}f���k��mq���v�1e|�����®���l��$)���勻Ϡ��\����jҖ������  �  Ɨ=�?=z�=܎=�5=��=1�=k)=h� =Fu = =���<'��<��<�d�<���<���<I�<+��< ��<s,�<Yw�<o��<�
�<�R�<��<��<�$�<�h�<��<u��<�,�<4l�<���<���<c$�<}_�<x��<���<��<�=�<�p�<^��<x��<���<�"�<H�<�i�<Ӈ�<l��<F��<q��<���<���<��<���<-��<���<;��<?��<���<���<3u�<�J�<;�<:��<?��<lV�<��<���<�K�<���<�q�<9��<Ly�<���<�c�<���<�2�<w��<��<^9�<Մ�<�ʶ<�
�<CE�<�z�<���<�֭<���<� �<�?�<t[�<t�<ʉ�<)��<\��<���<{˚<�ט<��<t�<���<)��<:�<��<�
�<��<��<��<y�<O
�<�~<�z<��u<J�q<��m<��i<�e<��a<��]<��Y<�U<]�Q<��M<�I<�E<�A<��=<r�9<��5<��1<��-<K�)<��%<1"<�$<�?<�_<r�<T�<��
<�<R\<VF�;���;��;6H�;��;"��;���;��;��;��;vI�;I��;��;��; .�;H�;OƑ;�;�օ;��;��t;U�i;��^;@T;<�I;ľ?;��5;�&,;1�";n;bd;�;��:'�:���:s��:�:���:p��:g
�:(��:�cg:N�K:�0:	#:ν�93��9Ⱀ9u<9��8*9���۸�O�E���
ȹ5��� S���*�r�A���X��o�1��~z��]���r줺����B��	jƺ��Ѻ�ܺ5�������X���&
�n���1�1��=) ���%��
+�
t0��5�=;��@���E��bK���P��-V���[��a�jxf���k�Leq�$�v�sZ|�(뀻����f���"��
ߋ�����?V������͖�q����  �  	�=�?=��=�=�5=��=��=)=� =�t =} =e��<���<|�<Zc�<_��<���<�G�<��<��<�+�<�v�<��<\
�<�R�<$��<H��<I%�<i�<ë�<c��<�-�<gm�<��<I��<�%�<�`�<���<��<�	�<�>�<rq�<��<���<���<�"�<�G�<Li�<J��<���<~��<`��<���<���<���<���<���<d��<���<%��<|��<ӗ�<�t�<TJ�<��<���<T��<�V�<��<.��<TL�<x��<�r�<|��<�z�<l��<e�<���<!4�<���</�<k:�<���<0˶<"�<�E�<�z�<	��<]֭<s��<& �<"?�<�Z�<�r�<���<ܛ�<��<j��<*ʚ<p֘<��<T�<��<d��<��<��<&
�<��<��<��<��<�
�<5~<e	z<�v<��q<m�m<D�i<��e<��a<��]<Q�Y<Z�U<!�Q</�M<.�I<m�E<}�A<��=<%�9<��5<��1<d�-<��)<��%<�"<"<�<<�\<��<��<��
<<�Y<oB�;f��;��;|F�;��;���;��;���;���;��;/L�;���;��;���;3�;5�;ˑ;.ċ;�ۅ;�;��t;R�i;��^;�CT;��I;ҿ?;��5;�#,;t�";�i;]^;��;���:���:/��:&}�:�Ӽ:@��:O��:���:��:�@g:a�K:v�0:�:ª�9���9���9�#<9J�8�5�}Q۸$O��ڗ���ǹ:<��='���*�j�A���X��o�!���j��C���[㤺����>���gƺ�Ѻ��ܺY���%��A��N/
����8<�����3 �1�%��+��}0� �5�1E;� �@�tF�fK�v�P�C/V��[�a�,uf�{�k��_q���v��Q|�`总�����`������ً�����wQ��-��ʖ������  �  H�=@=��=�=�5=x�=͂=�(=�� =xt =) =��<��<��<�b�<���<���<0G�<r��<v��<*+�<Ev�<���<5
�<�R�<9��<s��<�%�<�i�<Y��<���<�.�<n�<���<��<t&�<�a�<a��<���<k
�<;?�<�q�<E��<��<���<�"�<�G�<
i�<��<<��<޷�<���<���<���<���<���<��<���<C��<u��<��<5��<t�<�I�<��<���<_��<�V�<7�<���<�L�<��<~s�<#��<Q{�<)��<�e�<���<�4�<|��<��<;�<P��<�˶<~�<�E�<�z�<
��<B֭<#��<��<�>�<Z�<_r�<���<'��<K��<���<_ɚ<�՘<���<��<H�<���<�<�<�	�<��<��<��<�<J�<S~<�
z<v<��q<��m<��i<;�e<�a<�]<��Y<��U<R�Q<\�M<.�I<��E<��A<��=<�9<��5<�1<y�-<��)<��%<�
"<� <H;<P[<�<��<W�
<�<�X<�?�;��;&��;�D�;�;5��;6��;,��;���;��;YN�;ס�;#�;6��;�5�;1�;-Α;�Ƌ;;ޅ;c�;��t;޼i;��^;�FT;�I;��?;��5;�",;5�";Bf;uZ;e�;i��:���:�~�:�q�:�Ƽ:z�:���:�:���:�,g:٨K:1�0:�:�9D��9D��9�1<9O�8�=2���ڸ�N�1����ǹb��L��i*���A�E�X��qo�����a��Ѣ��Uۤ�����;��kfƺ��ѺA�ܺ����	�.��\��54
�R���A����W: ���%�F+���0�_�5�4J;�ҩ@�1	F�0iK�(�P��/V���[��a�Lsf���k�9[q���v�M|��〻�����]��2���֋������N���
���ǖ�G����  �  ��=�C=��=x�=�:=��=�=G.=?� =z =� =Ƌ�<���<w$�<�q�<���<��<[�<���<���<�E�<���<I��<0,�<�v�<���<	�<AP�<3��<��<��<�a�<D��<��<�#�<�b�<���<f��<��<jR�<L��<��<���<�$�<�R�<�}�<C��<���<8��<e�<� �<m6�<;H�<_V�<{`�<�f�<Hh�<Re�<�]�<CP�<n=�<$�<[�<3��<���<x�<(9�<��<P��<�I�<��<��<F�<���<�<É�<I��<�a�<�¿<��<�q�<ƿ�<s�<0I�<��<l��<>�<��<>�<�`�<@~�<��<`��<���<]Ң<��<|�<���<U�<�
�<��<�<��<B#�<�&�<�(�<�)�<p)�<�'�<�$�<� �<��<
+~<�z<:v< r<�m<��i<��e<��a< �]<�Y<w�U<͘Q<�M<�I<-�E<�zA<gu=<�p9<_m5<@k1<)k-<"m)<$r%<�z!<��<��<�<��<��<y
<6O<��<��;"�;��;o�;�,�;c��;���;m��;1��;h�;��;�Z�;͹�;�3�;Qɛ;�|�;�N�;z?�;*Q�;{;��o;ڎd;�Y;�O;'�D;�:;S�0;';,�;�f;�h;��;�"�:an�:�(�:cK�:Iֳ:�ä:f�:Ƴ�:�Ts:��W:�<:7{":�n:��9@٪9hnq9�=9�/8
V��"�0�u��~���ٹ�1�ae��c2��8I���_�hv�g��M���'�������ʲ�jؽ�i�Ⱥ��Ӻ+ߺa"�u9���' �����8�t���8�	���!�r�&���+��C1���6�|�;��;A�ƊF���K�O0Q�ʈV��[��Ea���f��l���q���v��i|�ɨ���b������ԋ�H���tD��:���Ǵ���n���  �  ��=�C=��=}�=�:=��=�=P.=Z� =Ez =&  =(��<Z��<�$�<�q�<a��<Y�<�[�<��<-��<(F�<���<l��<A,�<w�<���<��<)P�<��<���<��<.a�<��<���<�#�<b�<S��<��<B�<R�<��<���<���<~$�<�R�<�}�<U��<���<]��<��<� �<�6�<�H�<�V�<�`�<�f�<�h�<�e�<�]�<�P�<�=�<j$�<{�<R��<���<x�<B9�<���<2��<�I�<���<��<��<!��<��<q��<���<-a�<�¿<G�<yq�<l��<?�<I�<���<N��<6�<��<�>�<�`�<S~�<D��<���<¤<�Ң<O�<��<���<��<Y�<��<w�<	�<}#�<�&�<
)�<�)�<�)�<�'�<�$�<� �<p�<�*~<z<�v<X�q<D�m</�i<��e<��a<A�]<Y�Y<ġU<-�Q<��M<͇I<�E<�zA<xu=<�p9<�m5<�k1<Mk-<�m)<�r%<�{!<��<��<ױ<L�<Z�<E
<P<;�<?��;�"�;l��;�o�;2-�;��;���;��;���;��;B�;�Y�;���;2�;!ț;:{�;M�;L>�;�O�;M{;f�o;�d;)�Y;�O;p�D;��:;0�0;�';y�;.h;�i;ݢ;�'�:�t�:�.�:BR�:k۳:�Ȥ:2�:	��:�as:K�W:��<:�":+s:��9�ܪ90}q9K;9ߢ/8�BV�93��v�����Ծٹ�>��n��o2�jDI��_��sv�yl������������I̲�ڽ���Ⱥ��ӺRߺF �8���& ���Y6�8���5�����!���&�o�+��@1���6���;��9A��F�y�K�c/Q�އV���[��Fa�[�f��l��q�	�v�wl|�����E���d�����Ջ������E������ ���Uo���  �  @�=�C=��=t�=�:=��=V�=�.=�� =�z =�  =��<[��<&�<s�<���<O�<u\�<���<���<�F�<.��<���<w,�<$w�<���<��<�O�<|��</��<��<a`�<��<���<~"�<ba�<G��<���<p�<NQ�<P��<Z��<��<:$�<fR�<�}�<s��<��<���<"�<�!�<�7�<�I�<�W�<�a�<
h�<�i�<�f�<�^�<�Q�<{>�<2%�<�<���<��<$x�<?9�<���<��<RI�<C��<�~�<�<D��<��<T��<���<`�<~��<8�<�p�<���<y�<_H�<���<��<�<��<�>�<�`�<�~�<혨<q��<�¤<�Ӣ<<�< �<��<��<`�<��<]�<��<H$�<{'�<�)�<F*�<�)�<�'�<�$�<e �<��<t)~<�z<�v<��q<-�m<
�i<}�e<��a<!�]<��Y<%�U<��Q<B�M<��I<H�E<KzA<Lu=<!q9<n5<|l1<�l-<o)<ht%<R}!<t�<��<?�<��<��<I 
<R<��<���;&�;���;�q�;H.�;���;t��;���;���;��;��;�V�;���;{.�;+ě;w�;�H�;K:�;�K�;�z;��o;k�d;M�Y;~O;��D;��:;k�0;�';I�;fl;	o;��;�4�:%��:">�:�c�:Y�:�ۤ:�&�:ɇ:8�s:yX:�=:�":�:���9��9E�q9�%9�!/8�$W�M��#pv��Ū�
�ٹ$_�P����2��gI�G`���v�y��꜑�T����Ƨ�ZҲ�lݽ���Ⱥ��Ӻ[ߺ��/��! �����/����C.����3!�Y{&�9�+�791�|�6���;��3A� �F���K�B-Q��V���[�fHa���f��l�\�q�%�v��r|���h���Xh���!��ڋ�둎�qI��� �����r���  �  �=cC=��=i�=�:=��=��=/=@� =O{ =V! =͎�<��<�'�<�t�<:��<�<#^�<7��<3��<�G�<��<c��<�,�<?w�<c��<b�<O�<���<"��<z�<�^�<`��<��<� �<�_�<���<c��<��<�O�<*��<x��<Z��<�#�<(R�<�}�<ť�<p��<���<	�<�"�<�8�<K�<gY�<�c�<�i�<sk�<h�<�`�<)S�<�?�<J&�<�<���<l��<ox�<49�<w��<K��<�H�<S��<�}�<��<���<��<{��<���<9^�<���<��<o�<,��<J�<{G�<Ã�<}��<��<��<�>�<ia�<��<ܙ�<���<FĤ<Nբ<��<��<���<��<�<��<��<)!�<Z%�<h(�<2*�<�*�<�)�<�'�<^$�<��<9�<�'~<1z<
v<r�q<��m<��i<2�e<R�a<Ĳ]<S�Y<$�U<�Q<4�M<0�I<�~E<�yA<u=<wq9<�n5<�m1<Qn-<0q)< w%<b�!<��<)�<ȷ<Q�<F�<�#
<�U<�<��;g*�;���;"t�;<0�;n��;?��;N��;V��;9�;��;R�;���;�(�;���;�p�;�B�;�3�;�E�;>�z;ږo;�~d;��Y;jO;��D;�:;ʸ0;�';�;fr;�v;��;�J�:���:<Z�:_�:+
�:g��:XB�:)�:׳s:�/X:v4=:�":��:y��9q��9��q9�9L.8�X����5 w����bSڹԑ����Z�2�-�I�GF`���v����������Ɯ�`ӧ�nݲ��佺��Ⱥy�Ӻߺ�� "�� ���=$�]��2 ���G!��m&�d�+�n+1�`�6�!�;�+A��}F���K��)Q�/�V�b�[��Ja�g�f�{"l��q��w�`~|�A���ﴃ�4o��(�����������O�����񽖻v���  �  _�=�B=`�=]�=�:=2�=�=�/=�� =/| =E" =А�<I��<*�<w�<���<;�<`�<��<���<=I�<(��<0��<V-�<`w�<D��<��<DN�<���<���<��<
]�<m��<���<��<t]�<Z��<a��<��<1N�<���<0��<f��<#�<�Q�<�}�<��<��<���<O
�<Z$�<�:�<�L�<z[�<�e�<
l�<�m�<�j�<�b�<U�<�A�<�'�<:�<~��<��<�x�< 9�<,��<���<�G�<���<�{�<�	�<���<��<)��<���<�[�<]��<o�<�l�<_��<��<4F�<���<ֹ�<}�<��<Q?�<b�<���<��<(��<Ƥ<-ע<�<��<��<��<Q�<��<��<�"�<�&�<�)�<$+�<U+�<4*�<�'�<$�<�<:�<�$~<z<�v<��q<��m<�i<��e<��a<��]<^�Y<t�U<ϐQ<X�M<�I<F}E<�xA<�t=<�q9<�o5<eo1<�p-<t)<�z%<2�!<�<��<��<%�<�<w(
<�Y<�<��;J0�;���;�w�;�2�;s��;D��;���;m��;Nݼ;~�;L�;���;7!�;���;h�;�9�;J+�;>�;��z;�o;:sd;&�Y;fO;�D;��:;�0;�';��;�z;/�;�;ch�:P��:#|�:ţ�:�/�:��:�f�:U�:��s:7jX:�f=:N�":�:���9��9��q9��9x�,8[Z�l��q�w�����ڹg�����3���I�*�`�yw����H̑�ޜ��姺v벺���Ⱥ��Ӻ�޺��>��l � ��������σ��� �%[&���+�1�^t6���;�cA�!tF�(�K�+%Q�-�V���[��Ma���f��*l�Ǟq�;w�z�|����$���%x��M1���鋻Ӡ��nW�����OĖ��{���  �  ��=�B=�=G�=;=}�=��=L0=�� = } =a# =H��<���<�,�<�y�<'��<��<�b�<0��<���<�J�<^��<!��<�-�<�w�<��<P�<cM�<C��<��<��<�Z�<��<P��<��<�Z�<֘�<���<��<&L�<��<���<E��<M"�<xQ�<�}�<j��<���<���<��<&�<�<�<OO�<�]�<ph�<�n�<^p�<Im�<
e�<WW�<�C�<�)�<��<���<���< y�<
9�<���<ȟ�<SF�<[��<z�<��<'��< �<}��<���<Y�<���<��<�j�<J��<��<�D�<���<��<	�<��<�?�<�b�<���<���<賦<Ȥ<�٢<��<���<� �<�
�<��<�< �<�$�<�(�<+�<4,�< ,�<{*�<�'�<�#�<T�<�<�!~<rz<Lv<��q<��m<��i<(�e<��a<E�]<e�Y<�U<�Q<'�M<T�I<�{E<�wA<mt=<6r9<q5<dq1<Fs-<uw)<]~%<��!<�<�<�<��<�<�-
<�^<��<���;C7�;,��;.|�;25�;���;���;��;y��;^ؼ;��;E�;���;��;׫�;C^�;�/�;�!�;4�;��z;_zo;fd;��Y; O;�D;��:;��0;';�;��;�;��;���:D��:3��:R��:�Z�:�G�:���:,/�:Y=t:��X:��=:�#:��:�&�9�,�9S�q9ؼ9��+8Y|\�K�ܚx��	��S`۹�#�^�e3�*8J���`�<Uw��҆��ꑺ���i���{���������Ⱥ��Ӻ��޺�麃���� �`����}�����n�a� ��E&�@�+�a1�?b6���;��A��iF���K� Q�.�V���[�PQa���f�j4l��q��#w�9�|����ǃ�;����;���(���,a��K���˖������  �  �=B=��=9�=8;=��=�=�0=�� =&~ =�$ =ԕ�<���<�/�<�|�<���<k�<e�<u��<���<�L�<���<��<[.�<�w�<Ŀ�<��<HL�<ɐ�<Z��<��<�X�<j��<���<(�<�W�<��<#��<G�<�I�<���<&��<���<k!�<�P�<�}�<Ȧ�<���<���<8�<�'�<�>�<�Q�<�`�<2k�<|q�<+s�<p�<�g�<�Y�<�E�<_+�<
�<���<m��<Ly�<9�< ��<ў�<�D�<���<x�<0�<���<4�<�~�<���<V�<���<�<h�<䶺<���<�B�<^��<(��<��<��<�?�<�c�<Ȃ�<)��<͵�<;ʤ<ܢ<"�<S��<��<U�<��<��<s"�<�&�<o*�<n,�<C-�<�,�<�*�<�'�<#�<c�<��<�~<ez<��u<��q<�m<M�i<C�e<�a<ģ]<b�Y<U�U<ǈQ<��M<j}I<�yE<@vA<"t=<�r9<@r5<\s1<�u-<{)<��%<{�!<R�<w�<��<v�<c	<N3
<d<X�<���;�>�;���;`��;�7�; �;y��;���;���;Ӽ;O��;�<�;���;=�;}��;|S�;�$�;�;�)�;�z;�ho;�Wd;e�Y;�N;��D;��:;��0;�';��;B�;z�;�;��:�	�:���:Z��:���:zu�:���:zY�:M�t:��X:��=:>#:^	:MX�9�F�9Ӗq9��9��)8��^���X�y�������۹�w�P��D�3�%�J�	4a���w�3���������L���������Ⱥ��Ӻ!�޺h��A�������t���
�em����8X��� �/&�g�+���0�<O6�*�;�A�`^F���K��Q��~V�C�[�Va�F�f�e?l��q��3w�ү|�;��=҃�b����G��<��������j������Ӗ�R����  �  _�=�A=��=�=J;= �=��=�1=�� =3 =�% =L��<@��<S2�<u�<���<�<xg�<ƴ�<��<+N�<���<���<�.�<�w�<p��<��<>K�<]��<���<��<V�<Ӗ�<���<S�<U�<?��<|��<��<�G�<��<}��<���<� �<�P�<r}�<��<O��<���<��<�)�<�@�<T�<c�<�m�<Nt�<v�<�r�</j�<\�<�G�<)-�<��<���<(��<�y�<�8�<���<��<�C�<���<�u�<��< ��<f�<�{�<���<S�<ȴ�<:�<we�<���<���<SA�<�<I��<�<��<_@�<ad�<���<���<���<w̤<Tޢ<��<��<j�<#�<P�<*�<�$�<%)�<.,�<�-�<a.�<l-�<+�<m'�<|"�<~�<f�<$~<a
z<�u<��q<��m<��i<��e<)�a<@�]<1�Y<��U<��Q<M<�zI<wwE<�tA<�s=<�r9<�s5<ku1<�x-<z~)<͆%<<�!<`�<�<��<v�<+<�8
<-i<B�<��;�E�;���;���;�:�;� �;���;���;��;�ͼ;��; 5�;���;l�;
��;�H�;��;N�;��;Ȫz;�Wo;�Hd;�zY;��N;��D;��:;��0;�';F�;��;�;��;���:0�:L��:�&�:���:ʣ�: �:���:#�t:T9Y:�>:�n#:#-	:4��9h_�9�q9�S9-I(8Ca�H��8�z��'����ܹ���8��4���J�Ҍa�.�w���E0���2���+��������^�Ⱥ��Ӻ�޺��,������e���
�fZ����	B��� ��&��}+���0��<6��;�N�@��RF��K�DQ��|V�/�[�|Za���f�~Il���q��Cw��|�Y���܃������R���
������$u���(��ܖ�v����  �  ��=A=9�=��=c;=d�=��=U2=Q� =� =�& =���<���<�4�<��<I��<��<�i�<ܶ�<�<�O�<,��<���<b/�<�w�<*��<B�<2J�<��<���<��<�S�<[��<J��<��<sR�<���< ��<Y
�<�E�<0�<���<���<��<P�<_}�<n��<���<���<"�<i+�<�B�<GV�<�e�<kp�<�v�<�x�<<u�<�l�<D^�<�I�<�.�<��<���<���<�y�<�8�<��<��<iB�<S��<	t�<� �<s��<��<�x�<���<1P�<��<��<�b�<~��<���<�?�<�}�<l��<��<��<�@�<�d�<��<��<V��<uΤ<��<L�<���<	�<��<��<�!�<�&�<+�<�-�<N/�<C/�<.�<V+�<J'�< "�<��<.�<�~<�z<��u<��q<��m<8�i<.�e<Ĥa<�]<'�Y<�U<��Q<�{M<xI<buE<�sA<s=<Hs9<�t5<�v1<o{-<��)<��%<��!<d�<T�<��<��<j<O>
<+n<��<���;YL�;-��;H��;A=�;��;E��;���;���;"ɼ;/�;.�;R��;��;U��;w>�;��;K�;V�;4�z;/Ho;�:d;ioY;2�N;1�D;��:;ù0;�"';��;*�;ɱ;��;\��:�T�:U!�:�O�:=�:�ͥ:��:���:Q!u:'yY:�O>:��#:}N	:Y��9%x�9[�q9%!9�&8c�����f{������-ݹ�Uc��p4�ICK���a�EIx�1D��jO���N��UB��/�����ɺ=�Ӻ��޺��麴���)����V��
��G�����-��� �,&��h+���0�++6��;���@��GF�8�K��Q�{V��[��^a�P�f�YSl���q��Rw�K�|�/)��烻K���b]��0���ʎ����1���㖻%����  �  '�=�@=��=�=p;=��=d�=�2=� =� =�' =���<���<7�<g��<���<��<�k�<���<�<Q�<)��<s��<�/�<�w�<��<��<@I�<Ȍ�<L��<��<�Q�<L��<��<V�< P�<Y��<���<p�<�C�<�}�<���<���<��<�O�<K}�<���<z��<���<K�<�,�<�D�<)X�<�g�<�r�<y�<�z�<`w�<�n�<"`�<pK�<80�<�<��<?��<�y�<�8�<���<$��<?A�<���<Ur�<���<k��< �<fv�<b��<�M�<���<\�<�`�<���<R��<`>�<�|�<���<6�<��<�@�<�e�<셪<?��<κ�<Ф<{�<F�<���<P�<��< �<�#�<�(�<�,�<>/�<i0�< 0�<�.�<{+�<+'�<�!�<��<�<,~<Iz<�u<��q<5�m<��i<r�e<�a<��]<�Y<C�U</}Q<�xM<�uI<�sE<�rA<�r=<ss9<au5<�x1<�}-<s�)<͍%<L�!<\�<��<�<��<<�B
<7r<b�<{��;#R�;���;Ƌ�;?�;��;���;ż�;3��;�ļ;��;I'�;F�;H�;ۄ�;�5�;��;���;"�;��z;L:o;�.d;�eY;�N;�D;ۈ:;��0;�$';��;��;}�;�;�
�:[s�:.A�:�r�:�:��:�5�:�̈:�^u:9�Y:�>:��#:�k	:���9у�9�q9.�999%8?�e��<�l1|������ݹ6_����4�z�K��&b��x�7b��Wl���f��\V���>���#��Oɺ��Ӻ��޺t��?���m����J�\�
�U8����>�0� ��%�!X+�[�0�o6��|;�5�@�6?F���K��Q�*zV���[��ba���f��\l���q�A`w��|�
1���q����f��^���ӎ�����9��yꖻ�����  �  ��=f@=��=В=|;=��=��=93=�� =�� =m( =?��<���<�8�<��<;��<Y �<Um�<��<<�<�Q�<ޜ�<	��<�/�<�w�<���<:�<�H�<ߋ�<<��<��<oP�<���<V��<��<bN�<���<��<��<HB�<a|�<���<���<y�<EO�<:}�<§�<���<j��<�<�-�<�E�<�Y�<i�<Et�<�z�<u|�<y�<1p�<�a�<�L�<K1�<��<"��<���< z�<m8�<(��<���<a@�<���<q�<8��<���<���<�t�<���<�K�<խ�<�	�<K_�<��<!��<Z=�<�{�<%��<��<w�<	A�<f�<���<��<黦<|Ѥ<�<��<n�<��<��<��<,%�<U*�<�-�<K0�<,1�<�0�<�.�<�+�<'�<$!�<:�<4�<(~<� z<�u<y�q<��m< �i<�e<��a<�]<��Y<0�U<�zQ<�vM<�sI<drE<�qA<;r=<�s9<v5<�y1<-<|�)<G�%<L�!<��<
�< �<�<�<�E
<�u<p�<���;CV�;���;���;�@�;�;
��;n��;��;m��;��;d"�;�y�;��;F~�;/�;B �;�;d�;}z;B/o;�%d;^Y;�N;y�D;$�:;��0;o&';��;�;8�;�; �:���:�Z�:���:��:7�:�Q�:�:��u:��Y:�>:��#:��	:���9I��9{q9)�9Q$8)g�#����|�;x��޹>�����s�4���K��]b�L�x�{��򁒺Ox��e�� J���*��-ɺn�Ӻ��޺���������hA��
��+����s�*{ ���%��J+�ޮ0��6��r;���@�K9F�)�K��	Q�yV���[��ea��f�Scl���q�5jw��|��7������L����m��;%���ڎ�ȍ��?���ڟ���  �  h�=)@=��==�;=��=ߋ=3=�� =� =�( =(��<���<�9�<'��<I��<a!�<0n�<Ժ�<��<�R�<b��<Q��</0�<�w�<���<��<H�<>��<q��<��<�O�<���<L��<s�<3M�<���<)��<��<|A�<�{�<���<,��<�<O�<)}�<��<(��<���<��<�.�<�F�<lZ�<j�<Mu�<�{�<�}�<z�<1q�<bb�<�M�<�1�<z�<���<��<?z�<X8�<���<1��<�?�<'��<8p�<`��<���<���<is�<K��<�J�<���<��<K^�<9��<@��<�<�<m{�<ƴ�<��<m�<-A�<Jf�<���<���<���<=Ҥ<��<���<w�<�<��<��<&�<"+�<�.�<1�<�1�<.1�</�<�+�<�&�<� �<��<��<�~<5�y<Z�u<��q<��m<ζi<��e<?�a<�]<��Y<o~U<�xQ<uM<�rI<cqE<=qA<�q=<�s9<gv5<�z1<�-<߇)<ܑ%<�!<k�<0�<6�<c�<�< H
<Rw<�<���;&Y�;��;ڏ�;�A�;r�;���;���;B��;$��;��;k�;v�;6�;Tz�;�*�;���;��;��;�uz;:)o;�d;�XY;��N;��D;�:;C�0;�'';��;Я;D�;f;�,�:���:�j�:h��:�1�:3�:�b�:j��:�u:��Y:�>:��#:��	:.�9ʜ�9vq94�9�#8l8h���,}�J���(L޹����-5��K�nb��x�񉇺����G���o��R���/���ɺ5�Ӻ��޺D��]�������];�ư
�1%����
�Br ���%�DB+�S�0�;
6��l;�W�@��4F�_�K�iQ�3xV��[��ga���f�hl���q��pw���|��;������ⷆ�^r���)���ގ������B����ߢ���  �  `�=@=��=��=�;=��=�=�3=�� =� =�( =���<���<9:�<���<���<�!�<�n�<,��<E�<�R�<~��<i��<E0�<�w�<o��<��<�G�<'��<3��<��<!O�<@��<���<�<�L�<��<���<n�<*A�<D{�<ͳ�<��<��<O�<
}�<��<A��<���<��<�.�<�F�<�Z�<tj�<�u�<6|�<�}�<fz�<�q�<�b�<�M�<22�<��<���<���<@z�<78�<���<��<�?�<���<�o�<��<@��<;��<�r�<���<OJ�<@��<�<�]�<歺<���<�<�<B{�<���<��<Q�<7A�<_f�<��<ң�<޼�<�Ҥ<(�<<��<��<n�<�< �<|&�<z+�</�<(1�<�1�<H1�<;/�<�+�<�&�<� �<��<��<U~<��y<��u<��q<��m<�i<��e<z�a<?�]<�Y<�}U<HxQ<�tM<frI<qE<qA<�q=<�s9<�v5<�z1<[�-<)�)<}�%<��!<%�<��<��<8�<y<�H
<x<ح<���;�Y�;���;Q��;B�;;�;���;!��;ʱ�;ܾ�;��;7�;�t�;��;�x�;W)�;���;'�;R�;�rz;�&o;#d;�WY;G�N;��D;��:;^�0;(';z�;��;P�;�;-2�:��:q�:��:�7�:B%�:8g�:���:c�u:��Y:	�>:��#:W�	:w�99hgq9�9�H#8;vh����S}�齮�f޹������!5�_�K�A�b���x�[���t��������p��XT��J2��5ɺ��Ӻ��޺���k�������d9��
�c"������o ��%��?+�g�0��6�-j;�%�@��3F���K��Q�9xV���[�#ha���f��hl�D�q�
sw�f�|�=��-���q����s��i+��4�������C����������  �  h�=)@=��==�;=��=ߋ=3=�� =� =�( =(��<���<�9�<'��<I��<a!�<0n�<Ժ�<��<�R�<b��<Q��</0�<�w�<���<��<H�<>��<q��<��<�O�<���<L��<s�<3M�<���<)��<��<|A�<�{�<���<,��<�<O�<)}�<��<(��<���<��<�.�<�F�<lZ�<j�<Mu�<�{�<�}�<z�<1q�<bb�<�M�<�1�<z�<���<��<?z�<X8�<���<1��<�?�<'��<8p�<`��<���<���<is�<K��<�J�<���<��<K^�<9��<@��<�<�<m{�<ƴ�<��<m�<-A�<Jf�<���<���<���<=Ҥ<��<���<w�<�<��<��<&�<"+�<�.�<1�<�1�<.1�</�<�+�<�&�<� �<��<��<�~<5�y<Z�u<��q<��m<ζi<��e<?�a<�]<��Y<o~U<�xQ<uM<�rI<cqE<=qA<�q=<�s9<gv5<�z1<�-<��)<ܑ%<�!<k�<0�<6�<c�<�< H
<Rw<�<���;%Y�;��;ڏ�;�A�;q�;���;���;B��;#��;��;j�;v�;6�;Tz�;�*�;���;��;��;�uz;:)o;�d;�XY;��N;��D;�:;C�0;�'';��;Я;D�;f;�,�:���:�j�:h��:�1�:3�:�b�:j��:�u:��Y:�>:��#:��	:.�9ʜ�9vq94�9�#8l8h���,}�J���(L޹����-5��K�nb��x�񉇺����G���o��R���/���ɺ5�Ӻ��޺D��]�������];�ư
�1%����
�Br ���%�DB+�S�0�;
6��l;�W�@��4F�_�K�iQ�3xV��[��ga���f�hl���q��pw���|��;������ⷆ�^r���)���ގ������B����ߢ���  �  ��=f@=��=В=|;=��=��=93=�� =�� =m( =?��<���<�8�<��<;��<Y �<Um�<��<<�<�Q�<ޜ�<	��<�/�<�w�<���<:�<�H�<ߋ�<<��<��<oP�<���<V��<��<bN�<���<��<��<HB�<a|�<���<���<y�<EO�<:}�<§�<���<j��<�<�-�<�E�<�Y�<i�<Et�<�z�<u|�<y�<1p�<�a�<�L�<K1�<��<"��<���< z�<m8�<(��<���<a@�<���<q�<8��<���<���<�t�<���<�K�<խ�<�	�<K_�<��<!��<Z=�<�{�<%��<��<x�<	A�<f�<���<��<黦<|Ѥ<�<��<n�<��<��<��<,%�<T*�<�-�<K0�<,1�<�0�<�.�<�+�<'�<$!�<:�<4�<(~<� z<�u<y�q<��m< �i<�e<��a<�]<��Y<0�U<�zQ<�vM<�sI<drE<�qA<;r=<�s9<v5<�y1<-<|�)<G�%<L�!<��<
�< �<�<�<�E
<�u<p�<���;CV�;���;��;�@�;�;
��;n��;��;l��;��;d"�;�y�;��;F~�;/�;A �;�;c�;}z;B/o;�%d;^Y;�N;y�D;$�:;��0;o&';��;�;8�;�; �:���:�Z�:���:��:7�:�Q�:�:��u:��Y:�>:��#:��	:���9I��9{q9)�9Q$8)g�#����|�;x��޹>�����s�4���K��]b�L�x�{��򁒺Ox��e�� J���*��-ɺn�Ӻ��޺���������hA��
��+����s�*{ ���%��J+�ޮ0��6��r;���@�K9F�)�K��	Q�yV���[��ea��f�Scl���q�5jw��|��7������L����m��;%���ڎ�ȍ��?���ڟ���  �  '�=�@=��=�=p;=��=d�=�2=� =� =�' =���<���<7�<g��<���<��<�k�<���<�<Q�<)��<s��<�/�<�w�<��<��<@I�<Ȍ�<L��<��<�Q�<L��<��<V�< P�<Y��<���<p�<�C�<�}�<���<���<��<�O�<K}�<���<z��<���<K�<�,�<�D�<)X�<�g�<�r�<y�<�z�<`w�<�n�<"`�<pK�<80�<�<��<?��<�y�<�8�<���<$��<?A�<���<Ur�<���<k��< �<fv�<b��<�M�<���<\�<�`�<���<R��<`>�<�|�<���<6�<��<�@�<�e�<셪<@��<κ�<Ф<{�<F�<���<P�<��< �<�#�<�(�<�,�<>/�<i0�< 0�<�.�<{+�<+'�<�!�<��<�<,~<Iz<�u<��q<5�m<��i<r�e<�a<��]<�Y<C�U</}Q<�xM<�uI<�sE<�rA<�r=<ts9<bu5<�x1<�}-<t�)<͍%<L�!<\�<��<�<��<<�B
<6r<b�<z��;"R�;���;Ƌ�;?�;�;���;ļ�;3��;�ļ;��;I'�;F�;H�;ڄ�;�5�;��;���;"�;��z;L:o;�.d;�eY;�N;�D;ۈ:;��0;�$';��;��;}�;�;�
�:[s�:.A�:�r�:�:��:�5�:�̈:�^u:9�Y:�>:��#:�k	:���9у�9�q9.�999%8?�e��<�l1|������ݹ6_����4�z�K��&b��x�7b��Wl���f��\V���>���#��Oɺ��Ӻ��޺t��?���m����J�\�
�U8����>�0� ��%�!X+�[�0�o6��|;�5�@�6?F���K��Q�*zV���[��ba���f��\l���q�A`w��|�
1���q����f��^���ӎ�����9��yꖻ�����  �  ��=A=9�=��=c;=d�=��=U2=Q� =� =�& =���<���<�4�<��<I��<��<�i�<ܶ�<�<�O�<,��<���<b/�<�w�<*��<B�<2J�<��<���<��<�S�<[��<J��<��<sR�<���< ��<Y
�<�E�<0�<���<���<��<P�<_}�<n��<���<���<"�<i+�<�B�<GV�<�e�<kp�<�v�<�x�<<u�<�l�<D^�<�I�<�.�<��<���<���<�y�<�8�<��<��<iB�<S��<	t�<� �<s��<��<�x�<���<1P�<��<��<�b�<~��<���<�?�<�}�<l��<��<��<�@�<�d�<��<��<W��<uΤ<��<L�<���<	�<��<��<�!�<�&�<+�<�-�<N/�<C/�<.�<V+�<J'�< "�<��<.�<�~<�z<��u<��q<��m<8�i<.�e<Ĥa<�]<'�Y<�U<��Q<�{M<xI<buE<�sA<	s=<Is9<�t5< w1<o{-<��)<��%<��!<d�<T�<��<��<j<O>
<+n<��<���;YL�;,��;H��;@=�;��;D��;���;��;!ɼ;.�;.�;R��;��;U��;v>�;��;J�;V�;3�z;.Ho;�:d;hoY;2�N;0�D;��:;¹0;�"';��;*�;ɱ;��;\��:�T�:U!�:�O�:=�:�ͥ:��:���:Q!u:'yY:�O>:��#:}N	:Y��9%x�9[�q9%!9�&8c�����f{������-ݹ�Uc��p4�ICK���a�EIx�1D��jO���N��UB��/�����ɺ=�Ӻ��޺��麴���)����V��
��G�����-��� �,&��h+���0�++6��;���@��GF�8�K��Q�{V��[��^a�P�f�YSl���q��Rw�K�|�/)��烻K���b]��0���ʎ����1���㖻%����  �  _�=�A=��=�=J;= �=��=�1=�� =3 =�% =L��<@��<S2�<u�<���<�<xg�<ƴ�<��<+N�<���<���<�.�<�w�<p��<��<>K�<]��<���<��<V�<Ӗ�<���<S�<U�<?��<|��<��<�G�<��<}��<���<� �<�P�<r}�<��<O��<���<��<�)�<�@�<T�<c�<�m�<Nt�<v�<�r�</j�<\�<�G�<)-�<��<���<(��<�y�<�8�<���<��<�C�<���<�u�<��< ��<f�<�{�<���<S�<ȴ�<:�<we�<���<���<SA�<�<I��<�<��<_@�<ad�<���<���<���<w̤<Tޢ<��<��<j�<#�<P�<*�<�$�<%)�<.,�<�-�<a.�<k-�<+�<m'�<|"�<}�<f�<#~<a
z<�u<��q<��m<��i<��e<)�a<@�]<1�Y<��U<��Q<M<�zI<wwE<�tA<�s=<�r9<�s5<ku1<�x-<{~)<͆%<<�!<`�<�<��<v�<+<�8
<,i<A�<��;�E�;���;���;�:�;� �;���;���;��;�ͼ;��; 5�;;l�;	��;�H�;��;M�;��;Ȫz;�Wo;�Hd;�zY;��N;��D;��:;��0;�';F�;��;�;��;���:0�:L��:�&�:���:ʣ�: �:���:#�t:T9Y:�>:�n#:#-	:4��9h_�9�q9�S9-I(8Ca�H��8�z��'����ܹ���8��4���J�Ҍa�.�w���E0���2���+��������^�Ⱥ��Ӻ�޺��,������e���
�fZ����	B��� ��&��}+���0��<6��;�N�@��RF��K�DQ��|V�/�[�|Za���f�~Il���q��Cw��|�Y���܃������R���
������$u���(��ܖ�v����  �  �=B=��=9�=8;=��=�=�0=�� =&~ =�$ =ԕ�<���<�/�<�|�<���<k�<e�<u��<���<�L�<���<��<[.�<�w�<Ŀ�<��<HL�<ɐ�<Z��<��<�X�<j��<���<(�<�W�<��<#��<G�<�I�<���<&��<���<k!�<�P�<�}�<Ȧ�<���<���<8�<�'�<�>�<�Q�<�`�<2k�<|q�<+s�<p�<�g�<�Y�<�E�<_+�<
�<���<n��<Ly�<9�< ��<ў�<�D�<���<x�<0�<���<4�<�~�<���<V�<���<�<h�<䶺<���<�B�<^��<(��<��<��<�?�<�c�<Ȃ�<)��<͵�<;ʤ<ܢ<"�<S��<��<U�<��<��<s"�<�&�<o*�<n,�<C-�<�,�<�*�<�'�<#�<c�<��<�~<ez<��u<��q<�m<M�i<C�e<�a<ģ]<b�Y<U�U<ǈQ<��M<j}I<�yE<AvA<"t=<�r9<Ar5<\s1<�u-<{)<��%<{�!<R�<w�<��<v�<c	<N3
<d<X�<���;�>�;���;_��;�7�; �;x��;���;���;Ӽ;O��;�<�;���;=�;|��;|S�;�$�;�;�)�;߽z;�ho;�Wd;e�Y;~�N;��D;��:;��0;�';��;B�;z�;�;��:�	�:���:Z��:���:zu�:���:zY�:L�t:��X:��=:>#:^	:MX�9�F�9Ӗq9��9��)8��^���X�y�������۹�w�P��D�3�%�J�	4a���w�3���������L���������Ⱥ��Ӻ!�޺h��A�������t���
�em����8X��� �/&�g�+���0�<O6�*�;�A�`^F���K��Q��~V�C�[�Va�F�f�e?l��q��3w�ү|�;��=҃�b����G��<��������j������Ӗ�R����  �  ��=�B=�=G�=;=}�=��=L0=�� = } =a# =H��<���<�,�<�y�<'��<��<�b�<0��<���<�J�<^��<!��<�-�<�w�<��<P�<cM�<C��<��<��<�Z�<��<P��<��<�Z�<֘�<���<��<&L�<��<���<E��<M"�<xQ�<�}�<j��<���<���<��<&�<�<�<OO�<�]�<ph�<�n�<^p�<Im�<
e�<WW�<�C�<�)�<��<���<���< y�<
9�<���<ȟ�<SF�<[��<z�<��<'��< �<}��<���<Y�<���<��<�j�<J��<��<�D�<���<��<	�<��<�?�<�b�<���<���<賦<Ȥ<�٢<��<���<� �<�
�<��<�< �<�$�<�(�<+�<4,�<�+�<{*�<�'�<�#�<T�<�<�!~<rz<Lv<��q<��m<��i<(�e<��a<E�]<e�Y<�U<�Q<'�M<T�I<�{E<�wA<mt=<6r9<q5<dq1<Fs-<uw)<]~%<��!<�<�<�<��<�<�-
<�^<��<���;C7�;+��;-|�;15�;���;���;��;y��;]ؼ;��;E�;���;��;׫�;B^�;�/�;�!�;4�;��z;^zo;fd;��Y; O;�D;��:;��0;';�;��;�;��;���:D��:3��:Q��:�Z�:�G�:���:+/�:Y=t:��X:��=:�#:��:�&�9�,�9S�q9ؼ9��+8Y|\�K�ܚx��	��S`۹�#�^�e3�*8J���`�<Uw��҆��ꑺ���i���{���������Ⱥ��Ӻ��޺�麃���� �`����}�����n�a� ��E&�@�+�a1�?b6���;��A��iF���K� Q�.�V���[�PQa���f�j4l��q��#w�9�|����ǃ�;����;���(���,a��K���˖������  �  _�=�B=`�=]�=�:=2�=�=�/=�� =/| =E" =А�<I��<*�<w�<���<;�<`�<��<���<=I�<(��<0��<V-�<`w�<D��<��<DN�<���<���<��<
]�<m��<���<��<t]�<Z��<a��<��<1N�<���<0��<f��<#�<�Q�<�}�<��<��<���<O
�<Z$�<�:�<�L�<z[�<�e�<
l�<�m�<�j�<�b�<U�<�A�<�'�<:�<~��<��<�x�< 9�<,��<���<�G�<���<�{�<�	�<���<��<)��<���<�[�<]��<o�<�l�<_��<��<4F�<���<ֹ�<}�<��<Q?�<b�<���<��<)��<Ƥ<-ע<�<��<��<��<Q�<��<��<�"�<�&�<�)�<$+�<U+�<3*�<�'�<$�<�<:�<�$~<z<�v<��q<��m<�i<��e<��a<��]<_�Y<t�U<АQ<Y�M<�I<G}E<�xA<�t=<�q9<�o5<eo1<�p-<t)<�z%<3�!<�<��<��<%�<�<w(
<�Y<�<��;J0�;���;�w�;�2�;s��;D��;���;m��;Mݼ;}�;L�;���;7!�;���;h�;�9�;J+�;>�;��z;�o;9sd;%�Y;fO;�D;��:;�0;�';��;�z;/�;�;ch�:P��:#|�:ţ�:�/�:��:�f�:U�:��s:7jX:�f=:N�":�:���9��9��q9��9x�,8[Z�l��q�w�����ڹg�����3���I�*�`�yw����H̑�ޜ��姺v벺���Ⱥ��Ӻ�޺��>��l � ��������σ��� �%[&���+�1�^t6���;�cA�!tF�(�K�+%Q�-�V���[��Ma���f��*l�Ǟq�;w�z�|����$���%x��M1���鋻Ӡ��nW�����OĖ��{���  �  �=cC=��=i�=�:=��=��=/=@� =O{ =V! =͎�<��<�'�<�t�<:��<�<#^�<7��<3��<�G�<��<c��<�,�<?w�<c��<b�<O�<���<"��<z�<�^�<`��<��<� �<�_�<���<c��<��<�O�<*��<x��<Z��<�#�<(R�<�}�<ť�<p��<���<	�<�"�<�8�<K�<gY�<�c�<�i�<sk�<h�<�`�<)S�<�?�<J&�<�<���<l��<ox�<49�<w��<K��<�H�<S��<�}�<��<���<��<|��<���<9^�<���<��<o�<,��<J�<{G�<Ã�<}��<��<��<�>�<ia�<��<ܙ�<���<FĤ<Nբ<��<��<���<��<�<��<��<)!�<Z%�<h(�<1*�<�*�<�)�<�'�<^$�<��<9�<�'~<0z<

v<r�q<��m<��i<2�e<R�a<Ĳ]<S�Y<$�U<�Q<5�M<0�I<�~E<�yA<u=<wq9<�n5<�m1<Qn-<0q)< w%<b�!<�<)�<ȷ<Q�<F�<�#
<�U<�<��;g*�;���;"t�;;0�;m��;?��;M��;U��;9�;��;R�;�;�(�;���;�p�;�B�;�3�;�E�;>�z;ږo;�~d;��Y;jO;��D;�:;ʸ0;�';�;fr;�v;��;�J�:���:<Z�:_�:+
�:g��:XB�:)�:׳s:�/X:v4=:�":��:y��9q��9��q9�9L.8�X����5 w����bSڹԑ����Z�2�-�I�GF`���v����������Ɯ�`ӧ�nݲ��佺��Ⱥy�Ӻߺ�� "�� ���=$�]��2 ���G!��m&�d�+�n+1�`�6�!�;�+A��}F���K��)Q�/�V�b�[��Ja�g�f�{"l��q��w�`~|�A���ﴃ�4o��(�����������O�����񽖻v���  �  @�=�C=��=t�=�:=��=V�=�.=�� =�z =�  =��<[��<&�<s�<���<O�<u\�<���<���<�F�<.��<���<w,�<$w�<���<��<�O�<|��</��<��<a`�<��<���<~"�<ba�<G��<���<p�<NQ�<P��<Z��<��<:$�<fR�<�}�<s��<��<���<"�<�!�<�7�<�I�<�W�<�a�<
h�<�i�<�f�<�^�<�Q�<{>�<2%�<�<���<��<$x�<?9�<���<��<RI�<C��<�~�<�<D��<��<T��<���<`�<~��<8�<�p�<���<y�<_H�<���<��<�<��<�>�<�`�<�~�<혨<q��<�¤<�Ӣ<<�< �<��<��<_�<��<]�<��<H$�<{'�<�)�<F*�<�)�<�'�<�$�<e �<��<t)~<�z<�v<��q<-�m<
�i<}�e<��a<!�]<��Y<%�U<��Q<B�M<��I<H�E<KzA<Lu=<!q9<n5<}l1<�l-<o)<it%<R}!<t�<��<?�<��<��<I 
<R<��<���;&�;���;�q�;G.�;���;t��;���;���;��;��;�V�;���;{.�;+ě;w�;�H�;K:�;�K�;�z;��o;j�d;L�Y;~O;��D;��:;k�0;�';I�;fl;	o;��;�4�:%��:">�:�c�:Y�:�ۤ:�&�:ɇ:8�s:yX:�=:�":�:���9��9E�q9�%9�!/8�$W�M��#pv��Ū�
�ٹ$_�P����2��gI�G`���v�y��꜑�T����Ƨ�ZҲ�lݽ���Ⱥ��Ӻ[ߺ��/��! �����/����C.����3!�Y{&�9�+�791�|�6���;��3A� �F���K�B-Q��V���[�fHa���f��l�\�q�%�v��r|���h���Xh���!��ڋ�둎�qI��� �����r���  �  ��=�C=��=}�=�:=��=�=P.=Z� =Ez =&  =(��<Z��<�$�<�q�<a��<Y�<�[�<��<-��<(F�<���<l��<A,�<w�<���<��<)P�<��<���<��<.a�<��<���<�#�<b�<S��<��<B�<R�<��<���<���<~$�<�R�<�}�<U��<���<]��<��<� �<�6�<�H�<�V�<�`�<�f�<�h�<�e�<�]�<�P�<�=�<j$�<{�<R��<���<x�<B9�<���<2��<�I�<���<��<��<!��<��<q��<���<-a�<�¿<G�<yq�<l��<?�<I�<���<N��<6�<��<�>�<�`�<S~�<D��<���<¤<�Ң<O�<��<���<��<Y�<��<w�<�<}#�<�&�<
)�<�)�<�)�<�'�<�$�<� �<p�<�*~<z<�v<X�q<D�m</�i<��e<��a<A�]<Y�Y<ġU<-�Q<��M<͇I<�E<�zA<xu=<�p9<�m5<�k1<Mk-<�m)<�r%<�{!<��<��<ױ<L�<Z�<E
<P<;�<>��;�"�;l��;�o�;2-�;��;���;��;���;��;B�;�Y�;���;2�;!ț;:{�;M�;L>�;�O�;M{;f�o;�d;)�Y;�O;p�D;��:;0�0;�';y�;.h;�i;ݢ;�'�:�t�:�.�:BR�:k۳:�Ȥ:2�:	��:�as:K�W:��<:�":+s:��9�ܪ90}q9K;9ߢ/8�BV�93��v�����Ծٹ�>��n��o2�jDI��_��sv�yl������������I̲�ڽ���Ⱥ��ӺRߺF �8���& ���Y6�8���5�����!���&�o�+��@1���6���;��9A��F�y�K�c/Q�އV���[��Fa�[�f��l��q�	�v�wl|�����E���d�����Ջ������E������ ���Uo���  �  A�=H=f�=V�=�?=��=V�=�3=�� =� =w% =��<���<>1�<��<^��<6�<}n�<;��<�<�`�<���<U �<�N�<��<1��<�2�<|�<!��<�
�<�P�<���<s��<��<�^�<v��<��<� �<)_�<>��<^��<��<�G�<�{�<!��<"��<��<-�<�P�<mp�<}��<��<���<���<-��<���<A��<���<H��<��<3��<��<ƚ�<w�<�K�<��<���<6��<SF�<j��<b��<S#�<���<g5�<��<�&�<y��<��<{W�<
��<���<hJ�<N��<C̷<�<6�<bb�<��<ƪ�<�Ǭ<�ߪ<J��<*�<�<j�<�'�<�/�<_6�<�;�<z@�<�D�<�G�<�J�<GL�<M�<{L�<�J�<yG�<�B�<�<�<h5�<�,�<wF~<�1z<"v<�r<=�m<��i<��e<��a<R�]<�Y<�wU<ygQ<!XM<�II<�;E<'.A<	!=<39<;5<
�0<��,<��(<B�$<
� <S�<��< <Y<�0<�S	<>~<p�<d��;�V�;���;��;L9�;���;!��;d��;���;g��;�ų;���;*M�;��;WB�;.�;]��;?��;5��;�u;�Dj;�%_;�JT;رI;�X?;f?5;�a+;��!;�[;<0;�>;��:�:���:i�:a��:Ԁ�:ì�:|8�:XR~:��b:  H:ʰ-:��:���9��9�G�9��@9�ܾ8T x�'(����?�{⎹ƚ��칅�G�#���:�;�P�Mg�y}���˻��������������u��.g˺�aֺ�`�xg캲p���>����F���-:�r��@"�]l'��,�T2�7R7���<���A�G�WPL���Q�_�V�.\���a���f�wDl�u�q��w�{�|���������^g������ы�����'9��i쓻�����U���  �  !�=�G=R�=O�=�?=��=r�=�3=�� =� =�% =���<]��<�1�<��<���<��<�n�<���<s�<a�<3��<� �<�N�<+��<��<�2�<�{�<���<�
�<UP�<#��<��<!�<y^�<��<���<[ �<�^�<Û�<��<f�<OG�<�{�<���<.��<��<2-�<�P�<�p�<׌�<q��<>��<l��<���<,��<���<���<���<���<���<<��<
��<Sw�<�K�<��<���<��<(F�<(��<��<#�<>��<�4�<���<&�<��<���<W�<���<���<�I�<	��<�˷<��<�5�<5b�< ��<ߪ�<�Ǭ<(�<���<��<�<��<_(�<0�<�6�<0<�<A�<E�<qH�<K�<�L�<MM�<�L�<�J�<�G�<�B�<�<�<@5�<�,�<�E~<1z<;v<�r<]�m< �i<��e<�a<p�]<�Y<�vU<�fQ<�WM<)II<S;E<�-A<� =<b9<�5<z�0<�,<��(<�$<�� <O�<��<� <�<�1<�T	<F<g�<���;RX�;���;��;�9�;��;���;ש�;��;���;ų;?��;�K�;~��;�@�;��;���;ř�;���;�u;Aj;*#_;!IT;�I;�W?;5>5;ib+;g�!;H];2;
A;��:��:҉�:=p�:�Ĺ:��:o��:�A�:�`~:(�b:�H:[�-:��:���9d��9�N�9��@9�83\���c���?�*������� ���H�#���:��
Q�L[g���}�ɉ�PÔ�곟�������x���i˺�`ֺ�^��c��l��<����{B���[6���*"�-i'���,��2�`N7�}�<���A�WG��NL�6�Q���V�9.\�օa��f��Fl�_�q��w��|�I���R����h�����wӋ�\����:��&/����V���  �  Ǟ=�G=6�=J�=�?=�=��=4=D� =F� =S& =��<���<N3�<x��<���< �<Np�<���<~�<�a�<��<�<=O�<J��<���<e2�<o{�<"��<�	�<BO�<���<���<��<]�<���<>��<��<�]�<���<%��<��<�F�<O{�<Ǭ�<>��<!�<�-�<cQ�<�q�<ލ�<���<���<���<O��<���<��<��<���<���<���<?��<ܛ�<�w�<L�<��<���<Δ�<�E�<���<=��<"�<��<�3�<��<�$�<j��< ��<~U�<(��<>��<�H�<��<˷<C�<�5�<b�<)��<��<+Ȭ<��<r��<��<��<4 �<�)�<�1�<48�<�=�<�B�<hF�<�I�<L�<�M�<N�<VM�<@K�<�G�<�B�<y<�<�4�<�+�<gD~</z<�v<Qr<��m<9�i<}�e<�a<��]<r�Y<�tU<�dQ<�UM<�GI<x:E<V-A<� =<�9<&	5<��0<��,<��(<4�$<�� <��<��<V<<�4<�W	<�<�<u��;`\�;���;���;3;�;���;���;G��;���;ӣ�;³;>��;NG�;y��;D;�;�;ު�;?��;I��;��u;�8j;a_;(CT;��I;�U?;=5;=c+;�!;�`;p7;�G;�"�:s'�:��:��:޹:��:I˛:i[�:|�~:�c:L1H:��-:F:j#�9���9�Z�9��@9���8rϕ�O����@�y,��� ��m�i@�!$���:��9Q�ӈg�b�}��ۉ��Ԕ�8���$���.����{��Wk˺_ֺ.[Ẍ[�b���4����"9�^���+���u�!�1\'���,�9�1�-D7��<���A�:G��IL�K�Q�f�V�8.\�x�a��f��Kl���q�F"w��|�H ����n���$��*ً�򌎻�?����%���Z���  �  E�=[G=�=C�=@=P�=0�=�4=� =%� =O' =%��<��<�5�<؃�<���<T"�<yr�<���<5�<hc�<��<��<�O�<y��<���<�1�<�z�<��<f�<�M�<��<���<��<�Z�<J��<��<��<�[�<��<���<Y�<�E�<�z�<���<C��<��<W.�<dR�<�r�<x��<N��<���<���<y��<��<s��<B��<9��<���<y��<ֹ�<��<�x�<�L�<�<���<��<E�<���<��<j �<5��<�1�<ȭ�<?"�<��<���<8S�<骾<$��<�F�<��<�ɷ<K�<�4�<�a�<1��<i��<�Ȭ<��<���<%�<y�<M"�<�+�<�3�<�:�<@�<�D�<�H�<�K�<�M�<1O�<YO�<KN�<�K�<H�<�B�<%<�<-4�<�*�<�A~<�+z<Sv<(�q<0�m<��i<�e<{�a<1�]<4�Y<�pU<caQ<SM<�EI<�8E<|,A<� =<9<L
5<k 1<��,<��(<��$<�� <��<Y�<	<<�9<c\	<��<�<���;�b�;���;d��;�=�;��;���;ҧ�;���;�;���;V�;
@�;���; 3�;�ڒ;i��;Ջ�;��;�u;;+j;�_;�9T;ˤI;�P?;�;5;�c+;��!;.g;�?;�R;=�:�D�:x��:ة�:j�:�Ū:3�:�~�:e�~:�Tc:LlH:�.:�.:�f�9D'�9-v�9̝@9�R�8Es����¸��@����bn�����Ą�Y]$��;�ĀQ���g���}�C�����؟�5������������m˺�\ֺOSẠN캞P���)����)�4����D����!��I'���,�5�1�347��x<���A�X�F�EBL�3�Q��V�o.\�B�a���f��Sl���q��.w���|���������w���-��#⋻����;H��!���f����_���  �  ��=�F=��=/�=*@=��=��=|5=�� =M� =�( =��<��<�8�<���<���<T%�<'u�<C��<l�<2e�<}��<��<pP�<���<���<<1�<�y�<���<{�<�K�<���<���<��<�W�<:��<��<�<�X�<���<���<��<�D�<�y�<��<8��<��<)/�<�S�<ft�<y��<���<��<���<���<1��<���<I��<��<_��<���<Ի�<���< z�<�M�<��<���<��<!D�<5��<.��<C�<˪�<�.�<��<�<ˋ�<Z��<P�<	��<q��<�D�<`��<6ȷ<�<�3�<Qa�<2��<竮<�ɬ<�<g��<:
�<��<�$�<�.�<�6�<�=�<3C�<�G�<K�<AN�<FP�<(Q�<�P�<|O�<�L�<|H�<�B�<�;�<;3�<�)�<3>~<�'z<�v<��q<{�m<��i<Ӵe<>�a<Z�]<�{Y<�kU<]Q<WOM<�BI<�6E<A+A<; =<�9<�5<�1<�,<[�(<p�$<�� <7�<� <m<y$<@<�b	<:�<3�<>��;Pj�;\��;$��;$A�;���;c��;ȥ�;��;Қ�;���;U�;�6�;f��;�'�;�Β;���;F��;���;^vu;�j;s_;X-T;�I;�J?;�85;<d+;�!;Vn;VJ;`; ^�:Cl�:���:���:�2�:]��:�#�:)��:�1:{�c:h�H:	U.:�c:,��9�^�9l��9ݡ@9���8do�ĸ�kA����G���ԑ������$�)j;���Q�,h��J~��#���������ժ�ᱵ�j���Kr˺XZֺ<I�1?��9�������a�%�����n���!��0'���,���1�8 7��e<�.�A���F�9L�	�Q���V�p/\�W�a���f�%^l���q�=?w���|����˃�̓���9��k
����R�����Ŵ���f���  �  Ĝ=HF=f�=�=S@=�=j�=_6=� =�� =* =��<p��<C<�<���<j��<�(�<Rx�<.��<��<Lg�<*��<(�<Q�<��<K��<z0�<Ex�<վ�<`�<�H�<���<���<?�<JT�<Õ�<���<��<�U�<֓�<B��<�
�<C�<�x�<���</��<y�<0�<U�<Uv�<���<k��<*��<��<���<���<��<���<O��<i��<���<��<���<�{�<tN�<��<���<]��<C�<���<��<��<ߧ�<�+�<b��<j�<#��<���<mL�<���<?��<�A�<��<-Ʒ<��<�2�<�`�<-��<a��<�ʬ<��<Y��<��<��<�'�<2�<r:�<3A�<�F�<3K�<�N�<KQ�<�R�<iS�<�R�<�P�<�M�<�H�<�B�<;�<12�<(�<9:~<�"z<�
v<��q<��m<��i<­e<T�a<��]<huY<�eU<�WQ<#KM<L?I<S4E<�)A<�=<=9<I5<E1<��,<��(<��$<�� <��<�<�<�+<sG<�i	<��<^�<���;ps�;���;���;�D�;$��;���;|��;���;r��;ﭳ;�߬;�+�;Q��; �;���;r��;-s�;��;	_u;�j;��^;�T;��I;�C?;V55;�d+;��!;�v;�V;p;σ�:���:��:F�:Zk�:�1�:]�:��:��:Qd:I:��.:[�:��9���9���9W�@9|w�8����{Ÿ�`B�Ꝑ�Ŭ��%S�6E�Q+%�7�;�
QR�A�h�ݱ~�S��`<��\��󪺊ǵ�7���Qx˺�Wֺ?�-캵��;���]���u�R��$R���!�G'�Mk,�(�1�7��P<�q�A�1�F��-L�1~Q���V��0\�S�a�.�f�kl���q��Rw�T�|�|��5ك�f����G�����o���P_��L��׾��o���  �  ޛ=�E=�=��=z@=}�=�=L7==� =�� =�+ =���<��<@�<X��<1��<I,�<�{�<6��<��<�i�<��<o�<�Q�<��<���<�/�<�v�<���<�<F�<���<P��<��<P�<��<���<+�<�R�<ސ�<���<��<lA�<�w�<���<+��<��<!1�<�V�<Xx�<D��<=��<m��<���<���<}��<���<q��<���<���<^��<���<���<}�<qO�<Y�<���<���<�A�<���<߄�<�<���</(�<���<��<��<���<�H�<⠾<��<�>�<a��<	ķ<���<�1�<.`�<"��<٬�<�ˬ<#�<p��<�<��<E+�<�5�<,>�<�D�<�J�<�N�<=R�<�T�<�U�<�U�<�T�<bR�<�N�<LI�<�B�<a:�<�0�<`&�<�5~<�z<�v<��q<i�m<�i<�e<��a<]<�nY<�_U<ARQ<vFM<�;I<�1E<(A<9=<�9<�5<�1<M-<��(<$�$<� <�<<�<�3<LO<*q	<�<��<6�;P}�;��;���;7H�;���;d��;���;��;���;I��;լ;��;H��;�;:��;�z�;e�;4r�;>Fu;�i;?�^;T;��I;�;?;�15;qe+;��!;�;�c;ـ;E��:��:&Q�:�F�:t��:[o�:���:%�:��:�vd:�pI:��.:��:U��9���9ݑ9��@9 ��8�8��
ǸNdC��?���h��t ﹘����%�qS<��R��i�� �'���&j���@������޵������~˺�Uֺ�4�i������ �=q�����Z�n�� 4���!���&��M,��1�~�6��:<�݅A���F��"L�	wQ�5�V��1\�2�a�g��xl�@�q�jhw���|��,���烻T���*W��������l��}���ɖ�x���  �  ��=�D=��=ؗ=�@=��=��=58=a� =R� =%- =���<���<�C�<5��<���<�/�<�<8��<6�<�k�<���<��<�R�<,��<���<�.�<mu�<��<���<PC�<J��<���<�
�<�L�<��<)��<��<?O�<��<��<x�<�?�<wv�<Y��<��<T�<2�<X�<Hz�<���<��<���<	��<J��<G��<���<��<L��<���<6��<���<���<x~�<^P�<��<R��<���<�@�<��<���<S�<���<�$�<ϟ�<��<��<���<�D�<��<c�<�;�<���<���<��<�0�<�_�<���<N��<�̬<��<m��<��<h!�<v.�<+9�<�A�<�H�<UN�<�R�<�U�<�W�<�X�<DX�<�V�<�S�<|O�<�I�<dB�<�9�<�/�<�$�<F1~<Iz<��u<��q<�m<s�i<?�e<��a<�w]<lgY<:YU<�LQ<�AM<�7I<�.E<e&A<�=<9<n5<�
1<�-<1)<�%<V!<�<�<^&<�;<W<�x	<�<,�<��;Ć�;3�;>��;�K�;� �;���;���;��;���;%��;�ʬ;��;�y�;���;���;l�;�V�;cd�;V,u;��i;��^;��S;qxI;3?;y-5;Pe+;�!;*�;4p; �;Z��:��:S��:v�:��:��:�؜:`�:�?�:L�d:��I::C/:�':E��9H*�9:��9s�@9ej�8[)]�D�ȸtsD�䑹�"����`)�X&���<�)ES�W�i����i���3���/i���1����������O�˺Uֺ�*��_����� �_\�����@����u��y!���&�s0,���1���6��$<�<sA��F��L�pQ���V�z3\��a�g��l��r��}w��|��:��F���w���Qf��6���ˎ��z���'��Ԗ�|����  �  �=PD=;�=��=�@=?�=X�=9=g� =�� =�. = ��< ��<;G�<���<Q��<=3�<%��<��<��<�m�<3��<��<S�<K��<2��<�-�<t�<(��<Q��<�@�<B��<���<s�<I�<���<���<E�<L�<��<���<k�<$>�<[u�<���<���<��<�2�<zY�<|�<ښ�<���<���<B��<���<���<��<p��<���<���<���< ��<Q��<��<#Q�<�<"��<H��<T?�<Q��<]��<��<���<M!�<V��<��<;|�<���<�@�<���<�<�8�<(�<���<r��<�/�<�^�<∰<���<�ͬ<�<D �<��<$�<t1�<o<�<2E�<@L�<�Q�<�U�<�X�<�Z�<*[�<dZ�<uX�<U�<FP�<�I�<4B�<9�<�.�<�"�<-~<=z<��u<��q<P�m<4�i<��e<��a<�p]<�`Y<"SU<zGQ<=M< 4I<,E<�$A<�=<�9<�5<�1<S	-<T)<�%<:!<8<s<a-<�B<^<�	<��<-�<�;m��;E�;&��;O�;,�;���;���;���;��;퓳;���;I�;�m�;��;���;i^�;I�;�W�;Pu;��i;M�^;/�S;[lI;+?;^)5;e+;��!;a�;�{;Z�;	��:�!�:Ҵ�:	��:�::�:��:R��:pt�:>e:�%J:�/:e:�C�98c�9��9��@9ڻ8�m~��5ʸ%vE�C{��r���S��ݑ�|�&�m?=��S�n�i����IꊺW�����kP��c������˺/Tֺ�!�I�������� �xI�X�� (� �� ���]!�F�&�l,�3k1�v�6��<��bA��F��L�jQ���V�J5\���a�Ug���l��r�w��}�9G�����̽���t���(��,َ�b����3���ޖ�(����  �  S�=�C=��=��=�@=��=ۑ=�9=R� =�� =�/ =ƭ�<��<NJ�<���<Z��<6�<Ä�<f��<�!�<wo�<}��<��<�S�<g��<���<�,�<�r�<���<[��<G>�<���<���<e�<�E�<f��<���<L	�<~I�<���<���<��<�<�<kt�<��<���<	�<�3�<�Z�<�}�<˜�<��<��<���<���<���< �<g �</��<;��<��<��<ʧ�<݀�<�Q�<H�<���<���<R>�<���<�~�<��<��<��<6��<��<�x�<���<�=�<���<d�<6�<�|�<뽷<��<�.�<N^�<͈�<��<bά<,�<��<��<W&�<�3�<'?�<.H�<IO�<�T�<�X�<�[�<]�<R]�<P\�<�Y�<.V�<�P�<;J�<B�<Z8�<{-�<z!�<o)~<�z<��u<+�q<>�m<��i<��e<r|a<�j]<M[Y<NU<�BQ<A9M<�0I<�)E<2#A<9=<�9<�5<�1<-<)<.%<1!<�<_#<�3<4I<fd<��	<�<'�<��;��;�;���;�Q�;D�;���;y��;�~�;Wz�;���;ݷ�;���;�b�;.�;��;oR�;8=�;eL�;[ u; �i;��^;$�S;bI;K$?;6%5;�d+;�!;�;�;��;!�:�E�:���:���:EJ�:H�:�A�:�ǎ:��:Ïe:�mJ:��/:�:^��9o��9�0�9�@9�M�82����˸�LF�� ��Tr¹(c�!����&���=�VT�TVj�+������蕺����j���!�������˺(Sֺ�������� �>9���^��|����sE!���&��+��U1���6���;�mSA���F�:L��dQ���V�&7\�2�a��"g���l�(!r���w�,%}�	R�����ʆ�/����4��K去h����=���疻�����  �  ��=TC=��=o�=�@=��=?�=@:=� =n� =�0 =گ�<+��<�L�<��<���<18�<ц�<3��<>#�<�p�<p��<X	�<�S�<k��<x��<P,�<�q�<R��<���<�<�<�~�<x��<1�<�C�<
��<Q��<�<\G�<���<���<S�<�;�<�s�<���<���<0	�<@4�<g[�<�~�<G��<���<���<��<���<���<C�<��<G��<4��<���<���<��<���<eR�<f�<���<��<o=�<���<}�<��<��<Q�<ϖ�<6
�<kv�<��<N;�<+��<4�<#4�<A{�<���<���<�-�<�]�<���<0��<�ά<�<�<;�<(�<�5�<AA�<]J�<zQ�<W�<[�<�]�<�^�<�^�<�]�<[�<W�<pQ�<ZJ�<�A�<�7�<�,�<V �<�&~<Sz<��u<��q<��m<i�i<ϋe<�wa<f]<�VY<JU<5?Q<<6M<�.I<�'E<�!A<�=<�9<�5<�1<$-<�)<a%<!<�<�'<U8<�M<
i<
�	<X�<��<~&�;Ȝ�;X �;��;^S�;��;��;P��;�{�;�u�;��;9��;7��;KZ�;�ݘ;6��;fI�;�4�;�C�;�t;Ġi;#�^;��S; ZI;s?;�!5;Kd+;��!;��;C�;I�;�1�:{`�:���:��:�l�::�:be�:Y�:b:��e:D�J:��/:>�:���97��9�=�9��@9ݺ8ް���̸��F��j��}�¹���8�2'���=��eT�`�j�ZO���3������Ơ��~���1��������˺LSֺr����5���I� ��,�Ę���k�C���3!���&���+�#E1�S�6��;��GA�8�F���K�PaQ���V��8\���a�~)g�Ʃl��,r�i�w��4}��Z�����$ӆ�����>��3?����E���y����  �  ^�=
C=n�=]�=�@=��=t�=�:=n� =� =R1 =%��<���<�M�<y��<��<�9�<��<Q��<0$�<�q�<��<�	�< T�<e��<P��<�+�<Bq�<���<���<o;�<s}�<-��<� �<B�<q��<���<��<F�<���<���<n �<�:�<s�<p��<���<O	�<w4�<�[�<��<��<���<)��<b��<*��<b��<��<��<���<`��<���<R��<���<4��<�R�<��<���<ӏ�<�<�<���<&|�<��<՘�<��<n��<��<�t�<Y��<�9�<ʒ�<��<�2�<#z�<���<9��<7-�<�]�<���<Q��<>Ϭ<��<��<�< )�<,7�<�B�<�K�<�R�<vX�<h\�<�^�<'`�<�_�<�^�<�[�<~W�<�Q�<tJ�<�A�<�7�<,�<��<�$~<8	z<�u<�q<�m<�i<��e<zta<(c]<TY<�GU<=Q<<4M<�,I<�&E<T!A<\=<�9<!5<S1<�-<�)<l%<Y!<�<�*<F;<�P<l<��	<�<Y�<�*�;F��;P#�;���;�T�;�;���;��;gy�;�r�;D��;:��;]�;eU�;ؘ;�{�;BC�;�.�;�>�;��t;��i;E�^;'�S;�TI;�?;� 5;�c+;	�!;��;ǐ;ʼ;d?�:�r�:<�:'�:ԃ�:�Q�:}�:g�:�؀:�e:�J:�0:��:���9���9�G�9k�@9���8e2��#@͸�eG�����A0ù�>��a�te'�@">���T���j��c��vH�����aנ������;��b�����˺/Tֺ[�������� ��%�ۏ�G���`�����'!�-�&���+��:1��6���;�bAA�E�F��K��_Q�O�V��9\���a��-g�c�l�>4r�Թw�]>}�`��6���ن������D���󎻄����J���Y����  �  B�=�B=\�=Q�=�@=��=��=�:=�� =$� =�1 =���<���<`N�<��<i��<:�<w��<���<�$�<�q�<Z��<�	�<IT�<e��<8��<�+�<q�<R��<t��<	;�<�|�<���< �<�A�<+��<"��<>�<�E�<!��<l��< �<�:�<�r�<Q��<~��<v	�<�4�<'\�<��<\��<'��<���<���<���<���<,�<W�<��<���<9��<���<��<k��<�R�<��<���<���<�<�<���<�{�<>�<`��<\�<��<��<jt�<���<9�<P��<H�<�2�<�y�<U��<���<-�<v]�<���<t��<^Ϭ<��<�<l�<�)�<�7�<C�<,L�<oS�<�X�<�\�<__�<�`�<l`�<�^�<\�<�W�<�Q�<�J�<�A�<x7�<�+�<n�<$~<vz<��u<�q<�m<�i<%�e<�sa<b]<SY<�FU<9<Q<�3M<�,I<<&E<!A<(=<9<r5<�1<-<�)<B%<8!<c<�+<<<�Q<�l<�	<Ѵ<O�<,�;U��;k$�;`��;?U�;*�;}��;���;�x�;/r�;�;���;��;�S�;�՘;�z�;@B�;a,�;�<�;��t;��i;w�^;��S;-SI;(?;�5;Nc+;`�!;_�;��;ݾ;�C�:Wz�:[�:��:؊�:�X�:���:�:�ހ:)f:��J:�0:�:i��9���9uR�9�z@9���8�l��8{͸ފG��ē��Kù�_�p��w'�E+>�t�T�z�j�k��mP��`��ݠ�����m?��.����˺�Tֺ��q��N����� ��"���	��M]���� $!��&� �+�F71�ӎ6�4�;��?A�T�F���K�E^Q�x�V��:\���a��/g��l��6r�ܼw�B}�b��@ ���ۆ�葉�SF�� ���z���cL�����������  �  ^�=
C=n�=]�=�@=��=t�=�:=n� =� =R1 =%��<���<�M�<y��<��<�9�<��<Q��<0$�<�q�<��<�	�< T�<e��<P��<�+�<Bq�<���<���<o;�<s}�<-��<� �<B�<q��<���<��<F�<���<���<n �<�:�<s�<p��<���<O	�<w4�<�[�<��<��<���<)��<b��<*��<b��<��<��<���<`��<���<R��<���<4��<�R�<��<���<ӏ�<�<�<���<&|�<��<՘�<��<n��<��<�t�<Y��<�9�<ʒ�<��<�2�<#z�<���<9��<7-�<�]�<���<Q��<>Ϭ<��<��<�< )�<,7�<�B�<�K�<�R�<vX�<h\�<�^�<'`�<�_�<�^�<�[�<~W�<�Q�<tJ�<�A�<�7�<,�<��<�$~<8	z<�u<�q<�m<�i<��e<zta<(c]<TY<�GU<=Q<<4M<�,I<�&E<T!A<\=<�9<!5<S1<�-<�)<l%<Y!<�<�*<F;<�P<l<��	<�<Y�<�*�;F��;P#�;���;�T�;�;���;��;gy�;�r�;C��;:��;]�;eU�;ؘ;�{�;BC�;�.�;�>�;��t;��i;E�^;&�S;�TI;�?;� 5;�c+;	�!;��;ǐ;ʼ;d?�:�r�:<�:'�:ԃ�:�Q�:}�:g�:�؀:�e:�J:�0:��:���9���9�G�9k�@9���8e2��#@͸�eG�����A0ù�>��a�te'�@">���T���j��c��vH�����aנ������;��b�����˺/Tֺ[�������� ��%�ۏ�G���`�����'!�-�&���+��:1��6���;�bAA�E�F��K��_Q�O�V��9\���a��-g�c�l�>4r�Թw�]>}�`��6���ن������D���󎻄����J���Y����  �  ��=TC=��=o�=�@=��=?�=@:=� =n� =�0 =گ�<+��<�L�<��<���<18�<ц�<3��<>#�<�p�<p��<X	�<�S�<k��<x��<P,�<�q�<R��<���<�<�<�~�<x��<1�<�C�<
��<Q��<�<\G�<���<���<S�<�;�<�s�<���<���<0	�<@4�<g[�<�~�<G��<���<���<��<���<���<C�<��<G��<4��<���<���<��<���<eR�<f�<���<��<o=�<���<}�<��<	��<R�<ϖ�<6
�<kv�<��<N;�<+��<4�<#4�<A{�<���<���<�-�<�]�<���<0��<�ά<�<�<;�<(�<�5�<AA�<]J�<zQ�<W�<[�<�]�<�^�<�^�<�]�<[�<W�<pQ�<ZJ�<�A�<�7�<�,�<U �<�&~<Sz<��u<��q<��m<i�i<ϋe<�wa<f]<�VY<JU<5?Q<<6M<�.I<�'E<�!A<�=<�9<�5<�1<$-<�)<a%<!<�<�'<U8<�M<
i<
�	<X�<��<~&�;Ȝ�;X �;��;]S�;��;��;P��;�{�;�u�;��;8��;7��;KZ�;�ݘ;5��;eI�;�4�;�C�;�t;ài;#�^;��S;�YI;r?;�!5;Kd+;��!;��;B�;H�;�1�:z`�:���:��:�l�::�:be�:Y�:b:��e:D�J:��/:>�:���97��9�=�9��@9ݺ8ް���̸��F��j��}�¹���8�2'���=��eT�`�j�ZO���3������Ơ��~���1��������˺LSֺr����5���I� ��,�Ę���k�C���3!���&���+�#E1�S�6��;��GA�8�F���K�PaQ���V��8\���a�~)g�Ʃl��,r�i�w��4}��Z�����$ӆ�����>��3?����E���y����  �  S�=�C=��=��=�@=��=ۑ=�9=R� =�� =�/ =ƭ�<��<NJ�<���<Z��<6�<Ä�<f��<�!�<wo�<}��<��<�S�<g��<���<�,�<�r�<���<[��<G>�<���<���<e�<�E�<f��<���<L	�<~I�<���<���<��<�<�<kt�<��<���<	�<�3�<�Z�<�}�<˜�<��<��<���<���<���< �<g �</��<;��<��<��<ʧ�<݀�<�Q�<H�<���<���<R>�<���<�~�<��<��<��<6��<��<�x�<���<�=�<���<e�<6�<�|�<콷<��<�.�<N^�<͈�<��<bά<,�<��<��<W&�<�3�<'?�<.H�<IO�<�T�<�X�<�[�<]�<R]�<O\�<�Y�<.V�<�P�<;J�<B�<Z8�<{-�<z!�<n)~<�z<��u<+�q<>�m<��i<��e<r|a<�j]<N[Y<NU<�BQ<A9M<�0I<�)E<2#A<9=<�9<�5<�1<-<)<.%<1!<�<_#<�3<4I<fd<��	<�<'�<��;��;�;���;�Q�;C�;���;y��;�~�;Vz�;���;ݷ�;���;�b�;.�;��;nR�;8=�;eL�;Z u;�i;��^;$�S;bI;K$?;6%5;�d+;�!;�;�;��;!�:�E�:���:���:EJ�:H�:�A�:�ǎ:��:Ïe:�mJ:��/:�:^��9o��9�0�9�@9�M�82����˸�LF�� ��Tr¹(c�!����&���=�VT�TVj�+������蕺����j���!�������˺(Sֺ�������� �>9���^��|����sE!���&��+��U1���6���;�mSA���F�:L��dQ���V�&7\�2�a��"g���l�(!r���w�,%}�	R�����ʆ�/����4��K去h����=���疻�����  �  �=PD=;�=��=�@=?�=X�=9=g� =�� =�. = ��< ��<;G�<���<Q��<=3�<%��<��<��<�m�<3��<��<S�<K��<2��<�-�<t�<(��<Q��<�@�<B��<���<s�<I�<���<���<E�<L�<��<���<k�<$>�<[u�<���<���<��<�2�<zY�<|�<ښ�<���<���<B��<���<���<��<p��<���<���<���< ��<Q��<��<#Q�<�<"��<H��<T?�<Q��<]��<��<���<M!�<V��<��<;|�<���<�@�<���<�<�8�<)�<���<s��<�/�<�^�<∰<���<�ͬ<�<D �<��<$�<t1�<o<�<2E�<@L�<�Q�<�U�<�X�<�Z�<)[�<cZ�<uX�<U�<EP�<�I�<4B�<9�<�.�<�"�<-~<<z<��u<��q<P�m<4�i<��e<��a<�p]<�`Y<"SU<zGQ<=M<!4I<,E<�$A<�=<�9<�5<�1<S	-<T)<�%<:!<9<s<a-<�B<^<�	<��<,�<�;l��;E�;%��;O�;+�;���;���;���;��;쓳;���;H�;�m�;��;���;i^�;I�;�W�;Pu;��i;M�^;/�S;[lI;+?;])5;e+;��!;a�;�{;Z�;	��:�!�:Ҵ�:	��:�::�:��:R��:pt�:>e:�%J:�/:e:�C�98c�9��9��@9ڻ8�m~��5ʸ%vE�C{��r���S��ݑ�|�&�m?=��S�n�i����IꊺW�����kP��c������˺/Tֺ�!�I�������� �xI�X�� (� �� ���]!�F�&�l,�3k1�v�6��<��bA��F��L�jQ���V�J5\���a�Ug���l��r�w��}�9G�����̽���t���(��,َ�b����3���ޖ�(����  �  ��=�D=��=ؗ=�@=��=��=58=a� =R� =%- =���<���<�C�<5��<���<�/�<�<8��<6�<�k�<���<��<�R�<,��<���<�.�<mu�<��<���<PC�<J��<���<�
�<�L�<��<)��<��<?O�<��<��<x�<�?�<wv�<Y��<��<T�<2�<X�<Hz�<���<��<���<	��<J��<G��<���<��<L��<���<6��<���<���<x~�<^P�<��<R��<���<�@�<��<���<T�<���<�$�<ϟ�<��<��<���<�D�<��<c�<�;�<���<���<��<�0�<�_�<���<N��<�̬<��<m��<��<h!�<v.�<+9�<�A�<�H�<UN�<�R�<�U�<�W�<�X�<DX�<�V�<�S�<|O�<�I�<dB�<�9�<�/�<�$�<F1~<Iz<��u<��q<�m<s�i<?�e<��a<�w]<lgY<:YU<�LQ<�AM<�7I<�.E<e&A<�=<9<o5<�
1<�-<2)<�%<V!<�<�<^&<�;<W<�x	<�<,�<��;Æ�;2�;=��;�K�;� �;���;���;��;���;$��;�ʬ;��;�y�;���;���;l�;�V�;bd�;U,u;��i;��^;��S;qxI;3?;y-5;Pe+;�!;)�;4p; �;Z��:��:S��:v�:��:��:�؜:`�:�?�:L�d:��I::C/:�':E��9H*�9:��9s�@9ej�8\)]�D�ȸtsD�䑹�"����`)�X&���<�)ES�W�i����i���3���/i���1����������O�˺Uֺ�*��_����� �_\�����@����u��y!���&�s0,���1���6��$<�<sA��F��L�pQ���V�z3\��a�g��l��r��}w��|��:��F���w���Qf��6���ˎ��z���'��Ԗ�|����  �  ޛ=�E=�=��=z@=}�=�=L7==� =�� =�+ =���<��<@�<X��<1��<I,�<�{�<6��<��<�i�<��<o�<�Q�<��<���<�/�<�v�<���<�<F�<���<P��<��<P�<��<���<+�<�R�<ސ�<���<��<lA�<�w�<���<+��<��<!1�<�V�<Xx�<D��<=��<m��<���<���<}��<���<q��<���<���<^��<���<���<}�<qO�<Y�<���<���<�A�<���<߄�<�<���</(�<���<��<��<���<�H�<⠾<��<�>�<a��<	ķ<���<�1�<.`�<"��<ڬ�<�ˬ<#�<p��<�<��<F+�<�5�<,>�<�D�<�J�<�N�<=R�<�T�<�U�<�U�<�T�<bR�<�N�<LI�<�B�<a:�<�0�<`&�<�5~<�z<�v<��q<i�m<�i<�e<��a<]<�nY<�_U<ARQ<vFM<�;I<�1E<(A<9=<�9<�5<�1<M-<��(<%�$<� <�<<�<�3<LO<*q	<�<��<6�;O}�;��;���;6H�;���;c��;���;��;���;H��;լ;��;G��;�;:��;�z�;e�;3r�;=Fu;�i;>�^;T;��I;�;?;�15;pe+;��!;�;�c;ـ;D��:��:&Q�:�F�:t��:[o�:���:%�:��:�vd:�pI:��.:��:U��9���9ݑ9��@9 ��8�8��
ǸNdC��?���h��t ﹘����%�qS<��R��i�� �'���&j���@������޵������~˺�Uֺ�4�i������ �=q�����Z�n�� 4���!���&��M,��1�~�6��:<�݅A���F��"L�	wQ�5�V��1\�2�a�g��xl�@�q�jhw���|��,���烻T���*W��������l��}���ɖ�x���  �  Ĝ=HF=f�=�=S@=�=j�=_6=� =�� =* =��<p��<C<�<���<j��<�(�<Rx�<.��<��<Lg�<*��<(�<Q�<��<K��<z0�<Ex�<վ�<`�<�H�<���<���<?�<JT�<Õ�<���<��<�U�<֓�<B��<�
�<C�<�x�<���</��<y�<0�<U�<Uv�<���<k��<*��<��<���<���<��<���<O��<i��<���<��<���<�{�<tN�<��<���<]��<C�<���<��<��<ߧ�<�+�<b��<k�<#��<���<mL�<���<@��<�A�<��<-Ʒ<��<�2�<�`�<-��<a��<�ʬ<��<Y��<��<��<�'�<2�<r:�<3A�<�F�<3K�<�N�<KQ�<�R�<iS�<�R�<�P�<�M�<�H�<�B�<;�<02�<(�<8:~<�"z<�
v<��q<��m<��i<­e<T�a<��]<huY<�eU<�WQ<#KM<L?I<S4E<�)A<�=<=9<I5<F1<��,<��(<��$<�� <��<�<�<�+<sG<�i	<��<^�<���;os�;���;���;�D�;#��;���;{��;���;r��;;�߬;�+�;P��;��;���;r��;-s�;��;_u;�j;��^;�T;��I;�C?;V55;�d+;��!;�v;�V;p;΃�:���:��:F�:Zk�:�1�:]�:��:��:Qd:I:��.:[�:��9���9���9W�@9|w�8����{Ÿ�`B�Ꝑ�Ŭ��%S�6E�Q+%�7�;�
QR�A�h�ݱ~�S��`<��\��󪺊ǵ�7���Qx˺�Wֺ?�-캵��;���]���u�R��$R���!�G'�Mk,�(�1�7��P<�q�A�1�F��-L�1~Q���V��0\�S�a�.�f�kl���q��Rw�T�|�|��5ك�f����G�����o���P_��L��׾��o���  �  ��=�F=��=/�=*@=��=��=|5=�� =M� =�( =��<��<�8�<���<���<T%�<'u�<C��<l�<2e�<}��<��<pP�<���<���<<1�<�y�<���<{�<�K�<���<���<��<�W�<:��<��<�<�X�<���<���<��<�D�<�y�<��<8��<��<)/�<�S�<ft�<y��<���<��<���<���<1��<���<I��<��<_��<���<Ի�<���< z�<�M�<��<���<��<!D�<5��<.��<C�<˪�<�.�<��<�<ˋ�<Z��<P�<	��<q��<�D�<`��<6ȷ<�<�3�<Qa�<3��<竮<�ɬ<�<g��<:
�<��<�$�<�.�<�6�<�=�<3C�<�G�<K�<AN�<FP�<(Q�<�P�<|O�<�L�<|H�<�B�<�;�<;3�<�)�<3>~<�'z<�v<��q<{�m<��i<Ӵe<>�a<Z�]<�{Y<�kU<]Q<WOM<�BI<�6E<A+A<; =<�9<�5<�1<�,<[�(<p�$<�� <8�<� <m<y$<@<�b	<:�<2�<>��;Pj�;[��;#��;#A�;���;c��;ǥ�;��;њ�;���;T�;�6�;f��;�'�;�Β;���;E��;���;]vu;�j;r_;X-T;�I;�J?;�85;<d+;�!;Vn;VJ;`; ^�:Cl�:���:���:�2�:]��:�#�:)��:�1:{�c:h�H:	U.:�c:,��9�^�9l��9ݡ@9���8eo�ĸ�kA����G���ԑ������$�)j;���Q�,h��J~��#���������ժ�ᱵ�j���Kr˺XZֺ<I�1?��9�������a�%�����n���!��0'���,���1�8 7��e<�.�A���F�9L�	�Q���V�p/\�W�a���f�%^l���q�=?w���|����˃�̓���9��k
����R�����Ŵ���f���  �  E�=[G=�=C�=@=P�=0�=�4=� =%� =O' =%��<��<�5�<؃�<���<T"�<yr�<���<5�<hc�<��<��<�O�<y��<���<�1�<�z�<��<f�<�M�<��<���<��<�Z�<J��<��<��<�[�<��<���<Y�<�E�<�z�<���<C��<��<W.�<dR�<�r�<x��<N��<���<���<y��<��<s��<B��<9��<���<y��<ֹ�<��<�x�<�L�<�<���<��<E�<���<��<k �<5��<�1�<ȭ�<@"�<��<���<8S�<骾<%��<�F�<���<�ɷ<L�<�4�<�a�<1��<i��<�Ȭ<��<���<&�<y�<M"�<�+�<�3�<�:�<@�<�D�<�H�<�K�<�M�<1O�<YO�<KN�<�K�<H�<�B�<%<�<,4�<�*�<�A~<�+z<Sv<(�q<0�m<��i<�e<{�a<1�]<4�Y<�pU<caQ<SM<�EI<�8E<|,A<� =<9<M
5<k 1<��,<��(<��$<�� <��<Y�<	<<�9<c\	<��<�<���;�b�;���;c��;�=�;��;���;ҧ�;���;�;���;U�;	@�;���;3�;�ڒ;i��;ԋ�;��;�u;;+j;�_;�9T;ˤI;�P?;�;5;�c+;��!;.g;�?;�R;=�:�D�:x��:ש�:j�:�Ū:3�:�~�:e�~:�Tc:KlH:�.:�.:�f�9D'�9-v�9̝@9�R�8Fs����¸��@����bn�����Ą�Y]$��;�ĀQ���g���}�C�����؟�5������������m˺�\ֺOSẠN캞P���)����)�4����D����!��I'���,�5�1�347��x<���A�X�F�EBL�3�Q��V�o.\�B�a���f��Sl���q��.w���|���������w���-��#⋻����;H��!���f����_���  �  Ǟ=�G=6�=J�=�?=�=��=4=D� =F� =S& =��<���<N3�<x��<���< �<Np�<���<~�<�a�<��<�<=O�<J��<���<e2�<o{�<"��<�	�<BO�<���<���<��<]�<���<>��<��<�]�<���<%��<��<�F�<O{�<Ǭ�<>��<!�<�-�<cQ�<�q�<ލ�<���<���<���<O��<���<��<��<���<���<���<?��<ܛ�<�w�<L�<��<���<Δ�<�E�<���<=��<"�<��<�3�<��<�$�<j��<��<~U�<(��<?��<�H�<��<˷<C�<�5�<b�<)��<��<+Ȭ<��<s��<��<��<4 �<�)�<�1�<48�<�=�<�B�<hF�<�I�<L�<�M�<N�<UM�<@K�<�G�<�B�<y<�<�4�<�+�<fD~</z<�v<Pr<��m<9�i<}�e<�a<��]<r�Y<�tU<�dQ<�UM<�GI<x:E<V-A<� =<�9<&	5<��0<��,<��(<4�$<�� <��<��<V<<�4<�W	<�<�<u��;`\�;���;���;3;�;���;���;G��;���;ӣ�;³;>��;MG�;y��;C;�;�;ު�;?��;I��;��u;�8j;`_;(CT;��I;�U?;=5;<c+;�!;�`;p7;�G;�"�:s'�:��:��:޹:��:I˛:i[�:|�~:�c:L1H:��-:F:j#�9���9�Z�9��@9���8rϕ�O����@�y,��� ��m�i@�!$���:��9Q�ӈg�b�}��ۉ��Ԕ�8���$���.����{��Wk˺_ֺ.[Ẍ[�b���4����"9�^���+���u�!�1\'���,�9�1�-D7��<���A�:G��IL�K�Q�f�V�8.\�x�a��f��Kl���q�F"w��|�H ����n���$��*ً�򌎻�?����%���Z���  �  !�=�G=R�=O�=�?=��=r�=�3=�� =� =�% =���<]��<�1�<��<���<��<�n�<���<s�<a�<3��<� �<�N�<+��<��<�2�<�{�<���<�
�<UP�<#��<��<!�<y^�<��<���<[ �<�^�<Û�<��<f�<OG�<�{�<���<.��<��<2-�<�P�<�p�<׌�<q��<>��<l��<���<,��<���<���<���<���<���<<��<
��<Sw�<�K�<��<���<��<(F�<(��<��<#�<>��<�4�<���<&�<��<���<W�<���<���<�I�<	��<�˷<��<�5�<5b�< ��<ߪ�<�Ǭ<(�<���<��<�<��<_(�<0�<�6�<0<�<A�<E�<qH�<K�<�L�<MM�<�L�<�J�<�G�<�B�<�<�<@5�<�,�<�E~<1z<;v<�r<]�m< �i<��e<�a<p�]<�Y<�vU<�fQ<�WM<)II<S;E<�-A<� =<b9<�5<z�0<�,<��(<�$<�� <O�<��<� <�<�1<�T	<F<g�<���;QX�;���;��;�9�;��;���;ש�;��;���;ų;?��;�K�;~��;�@�;��;���;ř�;���;�u;Aj;*#_;!IT;�I;�W?;5>5;ib+;g�!;H];2;
A;��:��:҉�:=p�:�Ĺ:��:o��:�A�:�`~:(�b:�H:[�-:��:���9d��9�N�9��@9�83\���c���?�*������� ���H�#���:��
Q�L[g���}�ɉ�PÔ�곟�������x���i˺�`ֺ�^��c��l��<����{B���[6���*"�-i'���,��2�`N7�}�<���A�WG��NL�6�Q���V�9.\�օa��f��Fl�_�q��w��|�I���R����h�����wӋ�\����:��&/����V���  �  P�=�L=P�=��=%E=8�=��=�8=�� =�� =Y* =���<��<<�<���< ��<�-�<x��<���<�'�<3{�<���<� �<Er�<0��<��<�]�<<��<d��<,<�<��<���<�<�V�<a��<���<;#�< f�<���<#��<�&�<�c�<��<���<}
�<�;�<yi�<{��<���<4��<��<+�<�-�<�A�<�R�<�_�<
i�<n�<�n�<.j�<`�<[O�<}7�<��<���<��<���<�@�<���<���<K:�<���<�[�<���<Y�<;��<d5�<��<F��<bG�<���<hۻ<j�<=U�<���<��<wݲ<���<9�<<2�<�D�<S�<�]�<�e�<Xk�<@o�<�q�<�s�<�t�<�u�<^v�<�v�<�v�<�u�<�s�<�p�<wl�<�f�<_�<�U�<,K�<:?�<�c~<�Gz<�*v<�r<��m<��i<F�e<��a<0~]<�dY<MU<[6Q<S M<"I<��D<��@<��<<��8<s�4<x�0<�x,<�f(<]W$<DK <D<2B<�F<�R<�e<�<�<d� <w�;�z�;���;��;w5�;L��;l��;�x�;�\�;�T�;!b�;���;�ȣ;�%�;���; =�;s��;�ڃ;��{;}p;��d;��Y;�N;�D;4�9;��/;!�%;�;;��;?�	;�� ;`�:��:�:�/�:��:���:�#�:���:%wl:ЦQ:��7:U�:k�:4-�9be�9�Qn9#�9�B?8�(:�x=�*fi�]���!�й��������f,�-�B�j�X�#�n�)H���!���헺G����y���@��dú��ͺ��غ���c��ǯ���[�����^�����K�a��#�7c(���-�Y�2��8��B=�zmB�]�G���L���Q�f0W�kr\�h�a�[g��kl�(�q�Z2w�Z�|����嵃��i������̋�E|��|+��ړ�1����9���  �  #�=rL=B�=��=.E=L�=ߒ=9=�� =�� =�* =���<���<�<�<!��<���<o.�<��<j��<(�<�{�<���<&!�<lr�<D��<��<�]�< ��<��<�;�<���<h��<}�<�U�<Ӛ�<��<�"�<de�<"��<���<f&�<Dc�<Ý�<���<L
�<�;�<�i�<���<��<���<s��<��<N.�<�B�<6S�<J`�<�i�<�n�<]o�<�j�<�`�<�O�<�7�<=�<��<��<���<�@�<���<1��<�9�<��<[�<��<pX�<���<�4�<\��<���<�F�<#��<�ڻ<�<�T�<h��<յ�<Kݲ<��<[�<2�<E�<}S�<a^�<Uf�<�k�<�o�<jr�<2t�<ku�<]v�<�v�<'w�<�v�<v�<0t�<q�<�l�<�f�<_�<�U�<K�<�>�<@c~<�Fz<�)v<�r<j�m<��i<�e<X�a<�|]<�cY<LU<^5Q<�M<d
I<��D<��@<��<<��8<��4<�0<�y,<�g(<=X$<jL <@E<�C<H<�S<�f<1�<^�<�� <Q�;�|�;z�;F��;36�;���;+��;Vx�;�[�;;S�;�`�;���;ǣ;�#�;��;�:�;J��;H؃;�{;�p;d�d;m~Y;ףN;�D;9�9;9�/;W�%;�<;��;�	;r� ;dg�:��:�%�:|8�:R��:`��:�,�:F�:ǈl:�Q:ɒ7:��:W�:�C�9�t�9ddn9��9?�>8ww:��a���i�1��ѹ���h�D{,��B���X�x�n�=Q��&)�������������D���ú3�ͺ��غe��˪�����W����hZ����3G�ί��#�^(�Q�-���2�"8�/?=��iB��G���L��Q��/W��r\�z�a��g�]nl���q�6w�t�|����u����k����ϋ��~���-��ܓ����Z;���  �  ��=,L=�=��=OE=��=?�=�9=�� =z� =�+ =h��<���<�>�<*��<���<W0�<��<��<{)�<�|�<���<�!�<�r�<|��<��<=]�<b��<��<�:�<"��<���<��<T�<ܘ�<��<� �<�c�<���<��<4%�<Ib�< ��<)��<
�<�;�<�i�<C��<ܺ�<���<���</�< 0�<ZD�<DU�<\b�<�k�<�p�<.q�<�l�<b�<Q�<�8�<��<���<P��<���<I@�<P��<b��<�8�<���<sY�<Z��<�V�<���<�2�<C��<���<�D�<v��<@ٻ<��<�S�<���<_��<ݲ<%��<��<3�<�E�<�T�<�_�<�g�<�m�<�q�<�t�<8v�<�w�<[x�<�x�<�x�<ox�<Tw�</u�<�q�<.m�<�f�<_�<�U�<�J�<>�<Ca~<aDz<�&v<$r<��m<��i<�e<h�a<y]<T`Y<�HU<�2Q<yM<�I<b�D<�@<��<<%�8<��4<��0<|{,< j(<)[$<�O < I<�G<hL<�W<]k<+�<7�<� <G�;	��;W�;���;-8�;��;N��;^w�;�Y�;�O�;�\�;]��;5��;-�;ߗ�;`3�;}��; у;��{;_�o;�d;huY;��N;D;h�9;ĥ/;��%;k?;p�;��	;� ;�|�:���:1C�:-V�:��:�:N�:(�:�l: �Q:4�7:�#:��:�w�9��90�n9Q�9{>8�9;�w��Vj�"a���sѹ= ���=�p�,��C�RY�go�sm��B�����Y͢�r���`O���ú��ͺT�غ�����~����N�y��GM���8�����"�3M(�a�-��2��8�i3=�J_B�)�G��L��Q��-W�Ir\���a��g�ul���q�b@w���|��
���s��1&���֋�j���w4��6⓻w���m?���  �  	�=�K=��=x�=yE=��=�=^:=�� =�� =�, =L��<���<B�<k��<���<_3�<���<���<�+�<�~�<P��<#�<�s�<���<s�<�\�<V��<���<�8�<��<R��<��<.Q�<ԕ�<��<��<�`�<��<���<'#�<�`�<ɛ�<H��<�	�<�;�<[j�<B��<;��<n��<���<��<�2�<WG�<AX�<�e�<�n�<�s�<*t�<Eo�<td�<2S�<�:�<U�<���<���<���<�?�<Y��<��<7�<���<W�<���<�S�<x��<m/�<��<���<�A�<���<�ֻ<��<!R�<d��<{��<�ܲ<)��<)�<4�<JG�<dV�<�a�<[j�<xp�<�t�<�w�<ry�<�z�<^{�<�{�<�{�<�z�<ly�<�v�<;s�<n�<Yg�<_�<U�<�I�<�<�<�]~<1@z<�!v<�r<��m<��i<˨e<S�a<Gs]<�ZY<�CU<@.Q<�M<�I<O�D<��@<o�<<��8<P�4<�0<�~,<0n(<�_$<EU <�N<�M<�R<�^<�q<{�<�<w� <�;a��;6�;���;�;�;���;@��;Vu�;*V�;�J�;�U�;_y�;���;��;��;�'�;��;�Ń;��{;1�o;��d;�eY;��N;�C;�9;��/;W�%;�C;��;Q�	;�� ;)��:���:�n�:߆�:j�:��:ʁ�:�X�:�%m:�MR:|8:�j:�7:��9ߧ9�n98�9��=8�<��S�5�j�:⣹-ҹ�������-�eC��Y��lo����ak���/���좺A����`��E"ú	�ͺ��غ��㺃��1���v?�W��>9�����d����"��3(�J{-���2���7� =��NB��~G�^�L���Q��*W��r\���a�%g�Sl�+�q�$Qw�˽|�o��"˃�`��Q2���⋻����F?���듻ꘖ��F���  �  *�=K=��=e�=�E=o�=��=l;=�� =0� =~. =��<���<*F�<���<��<p7�<u��<���<�.�<E��<L��<`$�<ft�<���<.�<�[�<���<���<`6�<$}�<���<V�<AM�<ё�<��<��<�\�<^��<���<~ �<x^�<3��<-��<A	�<�;�< k�<]��<��<���<��<��<B6�<=K�<M\�<�i�<�r�<�w�<x�<�r�<�g�<�U�<�<�<�<���<Q��<���<P?�<#��<Z��<�4�<���<�S�<���<�O�<6��<6+�<ȍ�<L��<�=�<��<�ӻ<��<�O�<���<d��<7ܲ<-��<��<:5�<I�<�X�<�d�<�m�<t�<�x�<�{�<�}�<�~�<t�<��<�<�}�<|�< y�<�t�<,o�<�g�<_�<�T�<wH�< ;�<6Y~<�:z<Mv<��q<@�m<Ľi<Ġe<#�a<fk]<sSY<D=U<�(Q<�M<%I<��D<d�@<�<<��8<'�4<�0<��,<Ls(<%f$<"\ <�V<V<\[<gg<Lz<�<�<� <�#�;���;��;��;@�;���;��;�r�;�Q�;.D�;�L�;�n�;��;��;	~�;o�;�Չ;O��;�w{;T�o;�jd;�QY;�N;n�C;<�9;�/;t�%;�I;��;�	;u;<��:���:c��:kƿ:IU�:SW�:�Œ:r��:?�m:~�R:�|8:5�:s�:�E�9�*�9`.o9��9�=8��>�J���k����g�ҹ�R ���B�-�@�C�� Z�q�o��Ԃ�7���V^����Uŭ��w��U0úF�ͺ}�غ��Iy�}e��5,�n�����������e���"��(��Z-�ؙ2��7�u=�6:B�PmG��L���Q��&W��s\�*�a��'g�Ռl�Z�q��fw�V�|��#��wڃ�����$B����!����M������񣖻P���  �  �=DJ=�=K�=�E=��=|�=�<=Q� =�� =�0 =_��<R��<�J�<o��<���<�;�<���<���<2�<��<���<�%�<bu�<Y��<��<�Z�<9��<s��<�3�<�y�<��<%�<�H�<&��<W��<(�<�X�<W��<��<f�<�[�<.��<���<��<�;�<�k�<���<߿�<=��<��<w!�<\:�<�O�<�`�<nn�<�w�<�|�<`|�<�v�<Jk�<�X�<k?�<��<���<���<���<�>�<���<1��<2�<���<�O�<���<K�<U��<<&�<Ԉ�<x��<~9�<䇽<�ϻ<��<LM�<���<��<�۲<@��<��<�6�<K�<D[�<�g�<Sq�<)x�<}�<L��<f��<���<��<ꃗ<$��<���<�<�{�<�v�<fp�<�h�<�^�<�S�<�F�<�8�<�S~<@4z<�v<S�q<U�m<_�i<+�e<�{a<Qb]<KY<y5U<�!Q<2M<��H<P�D<y�@<z�<<c�8<H�4<w�0<��,</y(<@m$<Td <e_<�_<4e<Fq<-�<L�<��<�� <2�;'��;��;a��;�D�;���;���;�o�;yK�;�;�;_B�;�a�;n��;���;�l�;��;�É;���;pV{;��o;�Nd;H:Y;�lN;p�C;ԟ9;�/;��%;;P;�;��	;�;���:<�:e��:��:_��:���:��:��:�1n:ES:��8:U(:��:���9���9m�o9��9��;8k]A���%m�gK����ӹ�� ����(.��zD�N�Z��|p�d���ߍ�2���yC���뭺����HAú��ͺָغ^��Ca��B��5��������p�����?�m�"�_�'��5-�qw2���7���<�p"B��YG���L���Q�"W��t\���a��3g��l��r��w�o�|�4��$샻%���U��{������,^�� ��L����Z���  �  �=rI=��= �=F=��=h�=�==�� =�� =�2 =���<:�<P�<���<���<�@�<8��<���<�5�<��<���<�'�<Pv�<���<P�<�Y�<l��<���<]0�<�u�<��<x��<�C�<��<+��<3�<�S�<��<��<��<Y�<��<k��<��<�;�<Cl�<��<���<���<��<=%�<�>�<=T�<�e�<}s�<�|�<|��<��<${�<	o�<3\�<B�<��<-��<n��<P��<�=�<&��<��</�<���<�K�<���<�E�<��<� �<f��<>��<w4�<Z��<�˻<8�<qJ�<���<���<�ڲ<$��<!�<�7�<M�<�]�<+k�<-u�<�|�<Ɓ�<S��<|��<���<��<���<k��<Y��<T��<0~�<�x�<�q�<i�<�^�<�R�<vE�<�6�<N~<&-z<�v<@�q<��m<;�i<��e<nqa<hX]<�AY<$-U<EQ<�M<��H<��D<K�@<��<< �8<r�4<�0<��,<(<�t$<�l <�h<�i<�o<�{<��<j�<J�<X� <)A�;��;#)�;F��;�I�;���;���;[l�;NE�;�2�;�6�;�S�;���;"�;Z�;�;���;���;�1{;��o;�0d; Y;mWN;��C;��9;@�/;��%;�U;�;�
;�2;x5�:�y�:51�:2Y�:�:���:,e�:�7�:p�n:��S:6q9:˕:*.:�N�9��9{�o9s�9?}:8�D���"�n��#����Թu]��0�}�.��E�E:[�Sq��c���#��TӘ�Ow�����Ĳ���Tú� κҶغ�x�G�.�����o���M�P����tq"�u�'�-�AR2��7�X�<��B��EG�J�L���Q��W��v\�6�a�J@g�.�l�]%r�X�w��}�F������2����i�����eƎ�ip��_������g���  �  ��=�H=�=��=NF=�=?�=?=i� =�� =�4 =���<�<U�<���<���<�E�<���<���<'9�<���<��<2)�<4w�<���<��<\X�<��<j��<-�<<r�<���<���<�>�<���<��<"�<O�<v��<%��<y�<=V�<ݓ�<���<��<�;�<�l�<G��<���<x��<7�<�(�<�B�<�X�<�j�<�x�<��<Y��<�<^�<�r�<o_�<�D�<�!�<[��<���< ��<�<�<g��<���<,�<B��<�G�<J��<�@�<ı�<Y�<�}�<���<u/�<�~�<�ǻ<�
�<�G�<A~�<���<�ٲ<
��<��<>9�<O�<�`�<�n�<y�<倣<���<<��<���<Í�<퍙<@��<���<��<���<���<~z�<�r�<�i�<�^�<�Q�<�C�<q4�<H~<&z<zv<�q<��m<�i<H�e<ga<pN]<I8Y<�$U<�Q<�M<��H<�D<��@<��<<��8<t�4<q�0<`�,<��(<�{$<1u <3r<�s<z<��<�<��<��<�� <@P�;���;3�;q��;WN�;���;ʤ�;]h�;�>�;�)�;�*�;�E�;|�;jќ;/G�;vߏ;��;&~�;�{;�io;�d;�Y;�AN;x�C;׉9;�/;-�%;�[;�;
;%H;(k�:q��:Vv�:ѥ�:�A�:�I�:O��::�do:�]T:6�9:l :H�:���9�7�9eAp9��9�98�$G��#�"�o�����$�չ&������g/���E���[���q�&����h�����h����>���Ҹ�fjú9	κ��غ�k㺎/�����I��-T�s���)����H"�Ԛ'���,�-2��o7�ѯ<���A�%2G�6yL���Q��W��x\���a�:Ng���l�x=r�۹w�P6}�]X�����ʆ�F~��.���َ�҂��
)��%Ζ�us���  �  ��=�G=~�=��=nF=��=�=#@=�� =C� =�6 =���<�
�<�Y�<v��<��<J�<ƚ�<���<_<�<���<.��<�*�< x�<���<>�<(W�<���<���<*�<�n�<���<~��<;:�<'~�<E��<a�<�J�<E��<L��<2�<�S�<���<W��<�<q;�<Ym�<Z��<���<���<!�<�,�<�F�<&]�<Uo�<8}�<���<���<���<E��<Qv�<Sb�<�F�<�#�<_��<[��<ʃ�<�;�<���<J��<7)�<պ�<�C�<���<5<�<���<I�<�x�<���<�*�<Qz�<�û<I�<�D�<|�<z��<ٲ<���<@�<k:�<�P�<c�<�q�<�|�<؄�<ˊ�<Ύ�<P��<j��<n��<r��<��<���<`��<��<C|�<�s�<�i�<8^�<�P�<,B�<52�<eB~<6z<��u<��q<��m<J�i<�xe<U]a<$E]<�/Y<gU<�Q<��L<��H<p�D<��@<��<<
�8<5�4<��0<�,<;�(<Ԃ$<�| <�z<�|<��<S�<��<��<A�<�<^�;E��;�<�;H��;�R�;��;V��;�d�;!8�;� �;��;h8�;m�;��;b5�;!͏;É�;�k�;��z;lIo;p�c;��X;m-N;��C;=9;�/;�%;b`;($;�#
;1\;A��:���:B��:���:B��:h��:��:�Ѕ:g�o:��T:ua::�a :��:,K�9K��9��p9��9uy789�I�G,�g9q��ʧ���ֹip�dV�L�/��\F�w\��Or�u�˪��TJ��-ݣ�/g���񸺯~ú�κ��غ0`㺻��������!;�͢�8	��k�(��H""�u'���,��2��P7�@�<�>�A��G��kL�&�Q�KW��{\�'�a�=[g�	�l�Tr��w��U}�Ii��%���݆�b���.A��9쎻Փ��9��	ܖ��~���  �  z�=�F=�=��=�F=��=��=A=�� =�� =/8 =U��<r�<�]�<k��<���<�M�<T��<���<?�<؎�<���<�+�<�x�<���<��<"V�<��<���<�'�<�k�<)��<���<%6�<�y�<��<G�<�F�<���< ��<]�<Q�<Տ�<��<I�<B;�<�m�<E��<��<���<��<x/�<3J�<�`�<Fs�<*��<u��<Վ�<���<���<>y�<�d�<�H�<�$�<B��<���<���<�:�<t��<I��<�&�<ڷ�<@�<��<�7�<m��<��<zt�<���<�&�<�v�<v��<d�<EB�<0z�<.��<3ز<���<��<b;�<kR�<'e�<t�<��<J��<���<ђ�<A��<k��<W��<��<Ԓ�<n��<܊�<���<�}�<�t�<7j�<�]�<%P�<�@�<70�<y=~<Oz<��u<�q<f�m<��i< pe<�Ta<�<]<�'Y<�U<�Q<_�L<s�H<o�D<��@<��<<L�8<��4<.�0<r�,<�(<v�$<�� <�<��<��<��<"�<��<��<o<�i�;	��;D�;���;�U�;'��;��;>a�;�2�;��; �;�,�;`�;A��;�%�;%��;{y�;$\�;��z;�-o;?�c;9�X;aN;p�C;>v9;��/;��%;�c;?,;�/
;�l;*��:�!�:N��:D&�:w˱:�բ:D�:Q�:,fp:cLU:�::_� :S:��9`é9e�p9��9�68�HL��[er�U|��g_׹�������0���F��\�X�r��2��3⎺}�����"������ú�κ��غyX㺫����;���%�ۉ� ���M�����"�ZU'���,���1��67��}<���A��G��`L��Q�lW�O~\�/�a�fg�*�l��gr���w��p}�?x��[5��W����Q����������{F��薻����  �  ��=YF=��=b�=�F='�=2�=�A=�� =�� =k9 =��<E�<�`�<t��<� �<�P�<��<4��<'A�<���<��<�,�<�x�<���<M�<6U�<���<��<p%�<i�<���<���<"3�<�v�<˺�<9��<�C�<އ�<���<�<@O�<V��<���<��< ;�<�m�<��<+��<Z��<��<�1�<�L�<�c�<v�<1��<y��<���<a��<3��<`{�<�f�<iJ�<�%�<���<���<W��<:�<;��<���<�$�<y��<|=�<(��<�4�<7��<k�<q�<u��<�#�<�s�<׽�<�<W@�<�x�<��<�ײ<���<��<'<�<�S�<�f�<v�<܁�<ኣ<E��<���<E��<o��<0��<ڗ�<]��<���<Ɍ�<e��<�~�<bu�<jj�<�]�<iO�<�?�<�.�<�9~<�z<��u<Q�q<K�m<��i<iie<�Na<�6]< "Y<3U<� Q<?�L<�H<��D<��@<7�<<�8<��4<&�0<#�,<��(<Ì$<�� <��<z�<-�<Ȟ<G�<��<X�<v<�r�;���;�I�;*��;�W�;���;��;2^�;�-�;u�;H�;�#�;V�;��;D�;���;m�;pP�;u�z;]o;3�c;�X;<N;C�C;�m9;%�/;�%;2f;�2;89
;'y;w��:E�:W�:rS�:���:��:4u�:�?�:�p:W�U:�;:�� :sI:h��9f��9V�p9�9��48MwN�4���Ns�M
����׹R:��6��0��JG��b]��2s��b����� ����)��0����!����ú�$κd�غuR�j��������G�Xw����C7�J��C�!�*='��,���1�d"7��l<���A��G��XL���Q�"W�?�\�N�a��og���l��wr�_�w�
�}�����uA�����Z���+^�����s����P��������  �  5�=�E=c�=B�=�F=O�=z�=$B=j� =c� =/: =���<)�<�b�<~��<g�<}R�<���<���<mB�<���<���<=-�<By�<���<�<�T�<��<��<#$�<�g�<���<���<1�<�t�<���<��<�A�<��<���<��<N�<���<N��<M�<�:�<n�<`��<���<H��<��<3�<TN�<Xe�< x�<*��<w��<���<(��<�<�|�<�g�<RK�<�&�<I��<���<��<�9�<���<͉�<}#�<��<�;�<6��<�2�<���<=�<�n�<I��<�!�<�q�<4��<� �<3?�<�w�<e��<5ײ<O��<��<�<�<?T�<�g�<2w�<Q��<x��<��<���<J��<a��<��<���<ꖕ<��<ۍ�<T��<W�<�u�<}j�<�]�<O�<�>�<�-�<*7~<�z<W�u<��q<n�m<h�i<Iee<LJa<�2]<@Y<�U<��P<��L<*�H<B�D<��@<��<<z�8<8�4<C�0<�,<ҕ(<��$<Ë < �<Z�<-�<��<9�<e�<��<�<x�;	��;fM�;���;tY�;"��;[��;�\�;=+�;��;y	�;�;7O�;��;��;䨏;1e�;KH�;��z;<
o;ļc;��X;|N;�C;i9;�/;��%;�g;6;�>
;�;���:]�:�0�:9p�:��:'�:���:b^�:4�p:��U:^8;:`!:=h:g#�9r�9��p9�9:48��O��5���s��`���bعu�hr�}&1���G�!�]�Xts�%���#*��V����>�������.��o�ú�)κ�غ�N㺊����������Kk����z(�����!��-'��},���1�7�ca<�2�A�v�F��SL�D�Q��W��\���a��ug���l�>�r��
x���}�늁�I�����~����f��e��˵���W��?�������  �   �=�E=Q�=9�=�F=]�=��=SB=�� =�� =m: =P��<��<Pc�<��<��<S�</��<>��<�B�<��<E��<c-�<hy�<���<��<T�<���<���<�#�<(g�<��<E��<r0�<t�<6��<h��<A�<h��<Z��<O�<�M�<%��<��<"�<�:�<-n�<���<��<���<�<�3�<�N�<�e�<�x�<���<��<1��<���<5��<^}�<;h�<�K�<�&�<m��<
��<��<�9�<B��<k��<#�<���<@;�<���<72�<>��<��<Bn�<���<� �<*q�<���<+ �<�>�<bw�<%��<ײ<I��< �<�<�<�T�<h�<�w�<ڃ�<���<���<)��<ܚ�<�<���<)��<b��<���<7��<���<��<�u�<�j�<v]�<�N�<�>�<g-�<06~<�z<8�u<`�q<+�m<�i<0de<�Ha<g1]<Y<�U<��P<��L<O�H<��D<��@<��<<��8<q�4<��0<��,<��(<��$<�� <@�<��<]�<4�<k�<��<��<�<�y�;���;�N�;7��;/Z�;^��;)��;�[�;*�;N�;��;i�; M�;㝜;��;���;*c�;�E�;��z;}o;��c;f�X;N;b�C;g9;�~/;}�%;�h;r7;A
;�;v��:�e�:*8�:}y�:9#�:�/�:���:�h�:�q:R�U:FJ;:w&!:zs:5�9��9�q9��9O�38o-P��b��t��{����ع��0��.=1�F�G��]�_�s�݈���3���Ù�
F��u����3��ݫúf+κ�غ�K�<��Ҝ������f�����#�t~�g�!�)'�xx,�@�1�a7�O]<�a�A�y�F�RL�-�Q�!W���\���a�xg���l�)�r�x��}�e����K���������\i�����7����Y�����������  �  5�=�E=c�=B�=�F=O�=z�=$B=j� =c� =/: =���<)�<�b�<~��<g�<}R�<���<���<mB�<���<���<=-�<By�<���<�<�T�<��<��<#$�<�g�<���<���<1�<�t�<���<��<�A�<��<���<��<N�<���<N��<M�<�:�<n�<`��<���<H��<��<3�<TN�<Xe�< x�<*��<w��<���<(��<�<�|�<�g�<RK�<�&�<I��<���<��<�9�<���<͉�<}#�<��<�;�<6��<�2�<���<=�<�n�<I��<�!�<�q�<4��<� �<4?�<�w�<e��<5ײ<O��<��<�<�<@T�<�g�<2w�<Q��<x��<��<���<J��<a��<��<���<ꖕ<��<ۍ�<T��<W�<�u�<}j�<�]�<O�<�>�<�-�<*7~<�z<W�u<��q<n�m<h�i<Iee<LJa<�2]<@Y<�U<��P<��L<+�H<C�D<��@<��<<z�8<8�4<C�0<�,<ҕ(<��$<Ë < �<Z�<-�<��<9�<e�<��<�<x�;	��;fM�;��;tY�;!��;[��;�\�;<+�;��;y	�;�;7O�;��;��;䨏;1e�;JH�;��z;<
o;ļc;��X;|N;�C;i9;�/;��%;�g;6;�>
;�;���:]�:�0�:9p�:��:'�:���:b^�:4�p:��U:^8;:`!:=h:g#�9r�9��p9�9:48��O��5���s��`���bعu�hr�}&1���G�!�]�Xts�%���#*��V����>�������.��o�ú�)κ�غ�N㺊����������Kk����z(�����!��-'��},���1�7�ca<�2�A�v�F��SL�D�Q��W��\���a��ug���l�>�r��
x���}�늁�I�����~����f��e��˵���W��?�������  �  ��=YF=��=b�=�F='�=2�=�A=�� =�� =k9 =��<E�<�`�<t��<� �<�P�<��<4��<'A�<���<��<�,�<�x�<���<M�<6U�<���<��<p%�<i�<���<���<"3�<�v�<˺�<9��<�C�<އ�<���<�<@O�<V��<���<��< ;�<�m�<��<+��<Z��<��<�1�<�L�<�c�<v�<1��<y��<���<a��<3��<`{�<�f�<iJ�<�%�<���<���<W��<:�<;��<���<�$�<y��<|=�<(��<�4�<7��<k�<q�<u��<�#�<�s�<ؽ�<�<W@�<�x�<��<�ײ<���<��<'<�<�S�<�f�<v�<܁�<ኣ<E��<���<E��<o��</��<ڗ�<]��<���<Ɍ�<e��<�~�<au�<jj�<�]�<hO�<�?�<�.�<�9~<�z<��u<Q�q<K�m<��i<iie<�Na<�6]< "Y<3U<� Q<?�L<�H<��D<��@<7�<<�8<��4<&�0<$�,<��(<Ì$<�� <��<z�<-�<Ȟ<G�<��<X�<v<�r�;���;�I�;)��;�W�;���;��;2^�;�-�;u�;H�;�#�;V�;��;D�;���;m�;pP�;t�z;\o;2�c;�X;<N;C�C;�m9;%�/;�%;1f;�2;89
;'y;w��:E�:W�:rS�:���:��:4u�:�?�:�p:W�U:�;:�� :sI:h��9f��9V�p9�9��48MwN�4���Ns�M
����׹R:��6��0��JG��b]��2s��b����� ����)��0����!����ú�$κd�غuR�j��������G�Xw����C7�J��C�!�*='��,���1�d"7��l<���A��G��XL���Q�"W�?�\�N�a��og���l��wr�_�w�
�}�����uA�����Z���+^�����s����P��������  �  z�=�F=�=��=�F=��=��=A=�� =�� =/8 =U��<r�<�]�<k��<���<�M�<T��<���<?�<؎�<���<�+�<�x�<���<��<"V�<��<���<�'�<�k�<)��<���<%6�<�y�<��<G�<�F�<���< ��<]�<Q�<Տ�<��<I�<B;�<�m�<E��<��<���<��<x/�<3J�<�`�<Fs�<*��<u��<Վ�<���<���<>y�<�d�<�H�<�$�<B��<���<���<�:�<t��<I��<�&�<ڷ�<@�<��<�7�<m��<��<zt�<���<�&�<�v�<v��<d�<EB�<0z�<.��<3ز<���<��<c;�<kR�<'e�<t�<��<J��<���<ђ�<A��<k��<W��<��<Ԓ�<n��<܊�<���<�}�<�t�<7j�<�]�<$P�<�@�<70�<y=~<Nz<��u<�q<f�m<��i< pe<�Ta<�<]<�'Y<�U<�Q<`�L<s�H<p�D<��@<��<<L�8<��4<.�0<r�,<�(<v�$<�� <�<��<��<��<"�<��<��<n<�i�;��;D�;���;�U�;'��;��;=a�;�2�;��;��;�,�;`�;@��;�%�;$��;zy�;#\�;��z;�-o;?�c;9�X;`N;p�C;=v9;��/;��%;�c;?,;�/
;�l;*��:�!�:N��:D&�:v˱:�բ:D�:Q�:,fp:cLU:�::_� :S:��9`é9e�p9��9�68�HL��[er�U|��g_׹�������0���F��\�X�r��2��3⎺}�����"������ú�κ��غyX㺫����;���%�ۉ� ���M�����"�ZU'���,���1��67��}<���A��G��`L��Q�lW�O~\�/�a�fg�*�l��gr���w��p}�?x��[5��W����Q����������{F��薻����  �  ��=�G=~�=��=nF=��=�=#@=�� =C� =�6 =���<�
�<�Y�<v��<��<J�<ƚ�<���<_<�<���<.��<�*�< x�<���<>�<(W�<���<���<*�<�n�<���<~��<;:�<'~�<E��<a�<�J�<E��<L��<2�<�S�<���<W��<�<q;�<Ym�<Z��<���<���<!�<�,�<�F�<&]�<Uo�<8}�<���<���<���<E��<Qv�<Sb�<�F�<�#�<_��<[��<ʃ�<�;�<���<J��<7)�<պ�<�C�<���<5<�<���<I�<�x�<���<�*�<Qz�<�û<J�<�D�<|�<z��<ٲ<���<@�<k:�<�P�<c�<�q�<�|�<؄�<ˊ�<Ύ�<Q��<j��<n��<r��<��<���<`��<��<C|�<�s�<�i�<7^�<�P�<,B�<52�<eB~<6z<��u<��q<��m<J�i<�xe<U]a<$E]<�/Y<gU<�Q<��L<��H<q�D<��@<��<<�8<5�4<��0<�,<;�(<Ղ$<�| <�z<�|<��<S�<��<��<A�<�<^�;D��;�<�;G��;�R�;��;U��;�d�; 8�;� �;��;g8�;m�;��;b5�; ͏;É�;�k�;��z;kIo;o�c;��X;l-N;��C;<9;�/;�%;a`;'$;�#
;0\;A��:���:B��:���:B��:h��:��:�Ѕ:g�o:��T:ua::�a :��:,K�9K��9��p9��9uy789�I�G,�g9q��ʧ���ֹip�dV�L�/��\F�w\��Or�u�˪��TJ��-ݣ�/g���񸺯~ú�κ��غ0`㺻��������!;�͢�8	��k�(��H""�u'���,��2��P7�@�<�>�A��G��kL�&�Q�KW��{\�'�a�=[g�	�l�Tr��w��U}�Ii��%���݆�b���.A��9쎻Փ��9��	ܖ��~���  �  ��=�H=�=��=NF=�=?�=?=i� =�� =�4 =���<�<U�<���<���<�E�<���<���<'9�<���<��<2)�<4w�<���<��<\X�<��<j��<-�<<r�<���<���<�>�<���<��<"�<O�<v��<%��<y�<=V�<ݓ�<���<��<�;�<�l�<G��<���<x��<7�<�(�<�B�<�X�<�j�<�x�<��<Y��<�<^�<�r�<o_�<�D�<�!�<[��<���< ��<�<�<g��<���<,�<C��<�G�<J��<�@�<ı�<Y�<�}�<���<u/�<�~�<�ǻ<�
�<�G�<A~�<���<�ٲ<��<��<>9�<O�<�`�<�n�<y�<倣<���<<��<���<Í�<썙<@��<���<��<���<���<~z�<�r�<�i�<�^�<�Q�<�C�<q4�<H~<&z<yv<�q<��m<�i<H�e<ga<pN]<I8Y<�$U<�Q<�M<��H<�D<��@<��<<��8<u�4<q�0<`�,<��(<�{$<1u <3r<�s<z<��<�<��<��<�� <?P�;���;3�;p��;VN�;���;ɤ�;\h�;�>�;�)�;�*�;�E�;~|�;iќ;.G�;vߏ;��;%~�;�{;�io;�d;�Y;�AN;w�C;։9;�/;,�%;�[;�;
;%H;(k�:q��:Vv�:ѥ�:�A�:�I�:O��::�do:�]T:6�9:l :H�:���9�7�9eAp9��9�98�$G��#�"�o�����$�չ&������g/���E���[���q�&����h�����h����>���Ҹ�fjú9	κ��غ�k㺎/�����I��-T�s���)����H"�Ԛ'���,�-2��o7�ѯ<���A�%2G�6yL���Q��W��x\���a�:Ng���l�x=r�۹w�P6}�]X�����ʆ�F~��.���َ�҂��
)��%Ζ�us���  �  �=rI=��= �=F=��=h�=�==�� =�� =�2 =���<:�<P�<���<���<�@�<8��<���<�5�<��<���<�'�<Pv�<���<P�<�Y�<l��<���<]0�<�u�<��<x��<�C�<��<+��<3�<�S�<��<��<��<Y�<��<k��<��<�;�<Cl�<��<���<���<��<=%�<�>�<=T�<�e�<}s�<�|�<|��<��<${�<	o�<3\�<B�<��<-��<n��<P��<�=�<&��<��</�<���<�K�<���<�E�<��<� �<f��<>��<x4�<Z��<�˻<8�<qJ�<���<���<�ڲ<$��<!�<�7�<M�<�]�<+k�<-u�<�|�<Ɓ�<S��<|��<���<��<���<j��<Y��<S��<0~�<�x�<�q�<i�<�^�<�R�<vE�<�6�<N~<&-z<�v<@�q<��m<;�i<��e<nqa<hX]<�AY<$-U<FQ<�M<��H<��D<L�@<��<<�8<r�4<�0<��,<(<�t$<�l <�h<�i<�o<�{<��<i�<J�<W� <(A�;��;")�;E��;�I�;���;���;Yl�;ME�;�2�;�6�;�S�;���;!�;Z�;�;���;���;�1{;��o;�0d; Y;lWN;��C;��9;@�/;��%;�U;�;�
;�2;x5�:�y�:51�:2Y�:�:���:,e�:�7�:p�n:��S:6q9:˕:*.:�N�9��9{�o9s�9?}:8�D���"�n��#����Թu]��0�}�.��E�E:[�Sq��c���#��TӘ�Ow�����Ĳ���Tú� κҶغ�x�G�.�����o���M�P����tq"�u�'�-�AR2��7�X�<��B��EG�J�L���Q��W��v\�6�a�J@g�.�l�]%r�X�w��}�F������2����i�����eƎ�ip��_������g���  �  �=DJ=�=K�=�E=��=|�=�<=Q� =�� =�0 =_��<R��<�J�<o��<���<�;�<���<���<2�<��<���<�%�<bu�<Y��<��<�Z�<9��<s��<�3�<�y�<��<%�<�H�<&��<W��<(�<�X�<W��<��<f�<�[�<.��<���<��<�;�<�k�<���<߿�<=��<��<w!�<\:�<�O�<�`�<nn�<�w�<�|�<`|�<�v�<Jk�<�X�<k?�<��<���<���<���<�>�<���<2��<2�<���<�O�<���<K�<U��<<&�<Ԉ�<x��<~9�<䇽<�ϻ<��<LM�<���<��<�۲<@��<��<�6�<K�<D[�<�g�<Tq�<*x�<}�<L��<f��<���<��<ꃗ<$��<���<�<�{�<�v�<fp�<�h�<�^�<�S�<�F�<�8�<�S~<?4z<�v<S�q<U�m<_�i<+�e<�{a<Qb]<KY<z5U<�!Q<2M<��H<P�D<y�@<{�<<d�8<H�4<x�0<��,</y(<@m$<Td <e_<�_<4e<Fq<,�<L�<��<�� <2�;&��;��;`��;�D�;���;���;�o�;xK�;�;�;^B�;�a�;m��;���;�l�;��;�É;���;oV{;��o;�Nd;G:Y;�lN;o�C;ӟ9;�/;��%;;P;�;��	;�;���:<�:e��:��:_��:���:��:��:�1n:ES:��8:U(:��:���9���9m�o9��9��;8k]A���%m�gK����ӹ�� ����(.��zD�N�Z��|p�d���ߍ�2���yC���뭺����HAú��ͺָغ^��Ca��B��5��������p�����?�m�"�_�'��5-�qw2���7���<�p"B��YG���L���Q�"W��t\���a��3g��l��r��w�o�|�4��$샻%���U��{������,^�� ��L����Z���  �  *�=K=��=e�=�E=o�=��=l;=�� =0� =~. =��<���<*F�<���<��<p7�<u��<���<�.�<E��<L��<`$�<ft�<���<.�<�[�<���<���<`6�<$}�<���<V�<AM�<ё�<��<��<�\�<^��<���<~ �<x^�<3��<-��<A	�<�;�< k�<]��<��<���<��<��<B6�<=K�<M\�<�i�<�r�<�w�<x�<�r�<�g�<�U�<�<�<�<���<Q��<���<P?�<#��<Z��<�4�<���<�S�<���<�O�<6��<6+�<ȍ�<M��<�=�<��<�ӻ<��<�O�<���<e��<7ܲ<.��<��<:5�<I�<�X�<�d�<�m�<t�<�x�<�{�<�}�<�~�<t�<��<�<�}�<
|�< y�<�t�<,o�<�g�<_�<�T�<wH�<;�<5Y~<�:z<Mv<��q<@�m<Ľi<Ġe<#�a<fk]<sSY<D=U<�(Q<�M<%I<��D<e�@<�<<��8<'�4<�0<��,<Ms(<%f$<"\ <�V<V<\[<gg<Lz<�<�<~� <�#�;���;��;��;@�;���;��;�r�;�Q�;-D�;�L�;�n�;��;��;~�;n�;�Չ;N��;�w{;S�o;�jd;�QY;�N;m�C;<�9;�/;t�%;�I;��;�	;u;;��:���:c��:kƿ:IU�:SW�:�Œ:r��:?�m:~�R:�|8:5�:s�:�E�9�*�9`.o9��9�=8��>�J���k����g�ҹ�R ���B�-�@�C�� Z�q�o��Ԃ�7���V^����Uŭ��w��U0úF�ͺ}�غ��Iy�}e��5,�n�����������e���"��(��Z-�ؙ2��7�u=�6:B�PmG��L���Q��&W��s\�*�a��'g�Ռl�Z�q��fw�V�|��#��wڃ�����$B����!����M������񣖻P���  �  	�=�K=��=x�=yE=��=�=^:=�� =�� =�, =L��<���<B�<k��<���<_3�<���<���<�+�<�~�<P��<#�<�s�<���<s�<�\�<V��<���<�8�<��<R��<��<.Q�<ԕ�<��<��<�`�<��<���<'#�<�`�<ɛ�<H��<�	�<�;�<[j�<B��<;��<n��<���<��<�2�<WG�<AX�<�e�<�n�<�s�<*t�<Eo�<td�<2S�<�:�<U�<���<���<���<�?�<Y��<��<7�<���<W�<���<�S�<x��<n/�<��<���<�A�<���<�ֻ<��<!R�<e��<|��<�ܲ<)��<)�< 4�<JG�<dV�<�a�<[j�<xp�<�t�<�w�<ry�<�z�<^{�<�{�<�{�<�z�<ly�<�v�<;s�<n�<Xg�<_�<U�<�I�<�<�<�]~<1@z<�!v<�r<��m<��i<˨e<S�a<Gs]<�ZY<�CU<@.Q<�M<�I<O�D<��@<o�<<��8<P�4<�0<�~,<0n(< `$<EU <�N<�M<�R<�^<�q<{�<�<w� <�;`��;5�;��;�;�;���;?��;Vu�;*V�;�J�;�U�;_y�;���;��;��;�'�;��;�Ń;��{;1�o;��d;�eY;��N;�C;�9;��/;W�%;�C;��;Q�	;�� ;)��:���:�n�:߆�:j�:��:ʁ�:�X�:�%m:�MR:|8:�j:�7:��9ߧ9�n98�9��=8�<��S�5�j�:⣹-ҹ�������-�eC��Y��lo����ak���/���좺A����`��E"ú	�ͺ��غ��㺃��1���v?�W��>9�����d����"��3(�J{-���2���7� =��NB��~G�^�L���Q��*W��r\���a�%g�Sl�+�q�$Qw�˽|�o��"˃�`��Q2���⋻����F?���듻ꘖ��F���  �  ��=,L=�=��=OE=��=?�=�9=�� =z� =�+ =h��<���<�>�<*��<���<W0�<��<��<{)�<�|�<���<�!�<�r�<|��<��<=]�<b��<��<�:�<"��<���<��<T�<ܘ�<��<� �<�c�<���<��<4%�<Ib�< ��<)��<
�<�;�<�i�<C��<ܺ�<���<���</�< 0�<ZD�<DU�<\b�<�k�<�p�<.q�<�l�<b�<Q�<�8�<��<���<P��<���<I@�<P��<b��<�8�<���<sY�<Z��<�V�<���<�2�<C��<���<�D�<v��<@ٻ<��<�S�<���<_��<ݲ<%��<��<3�<�E�<�T�<�_�<�g�<�m�<�q�<�t�<8v�<�w�<[x�<�x�<�x�<ox�<Tw�<.u�<�q�<.m�<�f�<_�<�U�<�J�<>�<Ca~<aDz<�&v<$r<��m<��i<�e<h�a<y]<T`Y<�HU<�2Q<zM<�I<b�D<�@<��<<&�8<��4<��0<|{,< j(<)[$<�O < I<�G<hL<�W<]k<+�<7�<� <G�;��;W�;���;-8�;��;N��;]w�;�Y�;�O�;�\�;]��;5��;,�;ޗ�;`3�;|��; у;��{;_�o;�d;huY;��N;D;g�9;ĥ/;��%;k?;p�;��	;� ;�|�:���:1C�:-V�:��:�:N�:(�:�l: �Q:4�7:�#:��:�w�9��90�n9Q�9{>8�9;�w��Vj�"a���sѹ= ���=�p�,��C�RY�go�sm��B�����Y͢�r���`O���ú��ͺT�غ�����~����N�y��GM���8�����"�3M(�a�-��2��8�i3=�J_B�)�G��L��Q��-W�Ir\���a��g�ul���q�b@w���|��
���s��1&���֋�j���w4��6⓻w���m?���  �  #�=rL=B�=��=.E=L�=ߒ=9=�� =�� =�* =���<���<�<�<!��<���<o.�<��<j��<(�<�{�<���<&!�<lr�<D��<��<�]�< ��<��<�;�<���<h��<}�<�U�<Ӛ�<��<�"�<de�<"��<���<f&�<Dc�<Ý�<���<L
�<�;�<�i�<���<��<���<s��<��<N.�<�B�<6S�<J`�<�i�<�n�<]o�<�j�<�`�<�O�<�7�<=�<��<��<���<�@�<���<1��<�9�<��<[�<��<pX�<���<�4�<\��<���<�F�<#��<�ڻ<�<�T�<h��<յ�<Kݲ<	��<[�<2�<E�<}S�<a^�<Uf�<�k�<�o�<jr�<2t�<ku�<]v�<�v�<'w�<�v�<v�<0t�<q�<�l�<�f�<_�<�U�<K�<�>�<@c~<�Fz<�)v<�r<j�m<��i<�e<X�a<�|]<�cY<LU<^5Q<�M<d
I<��D<��@<��<<��8<��4<�0<�y,<�g(<=X$<jL <@E<�C<H<�S<�f<1�<^�<�� <Q�;�|�;z�;E��;36�;���;+��;Vx�;�[�;;S�;�`�;���;ǣ;�#�;��;�:�;J��;G؃;�{;�p;d�d;m~Y;ףN;�D;9�9;9�/;W�%;�<;��;�	;r� ;dg�:��:�%�:|8�:R��:`��:�,�:F�:ǈl:�Q:ɒ7:��:W�:�C�9�t�9ddn9��9?�>8ww:��a���i�1��ѹ���h�D{,��B���X�x�n�=Q��&)�������������D���ú3�ͺ��غe��˪�����W����hZ����3G�ί��#�^(�Q�-���2�"8�/?=��iB��G���L��Q��/W��r\�z�a��g�]nl���q�6w�t�|����u����k����ϋ��~���-��ܓ����Z;���  �  �=�Q=��=7�=�J=��=(�=�==h� =ڈ =]. =���<���<cD�<���<��<;�<���<���<>�<&��<���<�A�<u��<b��<�:�<��<���<6$�<o�<��<��<>J�<��<}��<� �</g�<A��<<��<B6�<�x�<F��<v��<�2�<�j�<^��<(��<���<�%�<�J�<�k�<n��<���<ú�<���<���<��<��<���<y��<���<O��<���<Ϳ�<��<�n�<+7�<b��<��<R�<���<��<��<Ɛ�<	�<ax�<���<�>�<���<.�<�0�<@s�</��<��<J�<�;�<�]�<�y�<��<Ǡ�<���<:��<^��<���<���<\��<B��<˯�<���<���<���<b��<̡�<���<���<���<��<���<�|�<up�<ob�<S�<*�~<|`z</;v<kr<��m<o�i<7�e<%�a<�a]<�AY<#U<�Q<3�L<!�H<��D<�@<�v<<=X8<?94<�0<��+<��'<��#<��<Ŗ<ĉ<��<x�<7�<��<��<���;P#�;���;��;���;�!�; ��;Vu�;$6�;m�;��;�;m��;)-�; z�;~�;ut�;U&�;���;'�u;5j;��^;)�S;��H;i2>;��3;��);	 ;|z;�';f;&m�:�2�:�t�:X2�:�o�:-�:�f�:x�:��t:*�Y:�?:�X&:�:�y�9R��9]�9�99��8�ܴ=)��mE8��̉��:���f�V������4���J� �`�p5v��х�|����'���9N����i�ź�Wкm&ۺr��������
	�T��h�=r�o��S,$��p)���.���3���8�$�=��C�$#H�9M�0VR��}W�)�\��a�8g��l�S�q�$Ew�1�|����淃��h��o���ċ��o��I��ē��m������  �  ��=�Q=��=4�=�J=��=_�=9>=�� =+� =�. =q��<���<iE�<ԕ�<��<�;�<K��<���<�>�<̕�<~��<7B�<���<}��<�:�<��<���<�#�<�n�<N��<,�<qI�<=��<���<��<Rf�<`��<���<�5�<4x�<Ǹ�<��<�2�<�j�<f��<I��<7��<-&�<'K�<il�<��<p��<���<���<���<��<���<u��<@��<L��<���<+��<@��<Q��<�n�<17�<E��<���<�Q�<��<~��<�<��<�<ww�<���<�=�<���<H�<�/�<�r�<���<�<��<�;�<�]�<�y�<3��<��<$��<Ҵ�<���<.��<f��<��<1��<߰�<���<���<ħ�<)��<n��<F��<J��<��<`��<ᆉ<�|�<Yp�<Lb�<�R�<+�~<N_z<�9v<	r<�m<��i<p�e<t�a<`]<8@Y<�!U<�Q<"�L<7�H<H�D<Г@<v<<qX8<�94<�0<��+<<�'<��#<?�<_�<i�<ǅ<��<;�<6�<X�<���;�%�;l��;��;\��;�"�;���;ju�;�5�;��;��;.�;��;�*�;w�;:�;Pq�;�"�;_��;d�u;0j;��^;�S;+�H;�/>;��3;��);�	 ;�{;i*;;;w�:�=�:�~�:?�:�|�:F;�:�w�:�-�:��t:�Y:s�?:�m&:&�:t��9���9�r�9�+99�(�8ص�*E��p8�쉹	]�����m��*��L5��K�R�`�Qv�!߅������#������@V��������ź�Xк�$ۺ��2��U���{���ڀ� ��l�����#$��h)�!�.�Q�3�j�8�$�=�C��H�n5M�TR��|W�>�\���a�>9g�t�l�W�q��Iw��|�r	��Y���l�����ȋ�5s��,���Ɠ�#p������  �  .�=/Q=��=7�=(K=V�=�=�>=�� =+� =�/ =���<<��<H�<{��<���<�>�<ɓ�<���<�@�<v��<���<,C�<@��<���<�:�<���<���<�"�<m�<q��<��<"G�<ˎ�<(��<)�<�c�<��<h��<�3�<�v�<���<��<�1�<�j�<���<���<��<K'�<�L�<>n�<'��<Ѧ�<��<K��<:��<���<���< �<� �<e��<���<���<[��<��<:o�<U7�<���<��<�P�<���<���<��<ȍ�<��<�t�<���<J;�<$��<��<�-�<�p�<���<��<�<�:�<w]�<�y�<���<�<E��<^��<Ӻ�<W��<ӻ�<���<޶�<���<S��<0��<Q��<���<{��<��<���<1��<"��<Y��<�|�<�o�<�a�<�Q�<��~<�[z<�5v<�r<#�m<��i<<�e<f|a<[]<�;Y<�U<� Q<T�L<��H<ƮD<ޒ@<yv<<,Y8<;4<�0<u�+<��'<	�#<�<��<א<R�<2�<З<��<��<N��;<.�;���;o�;���;�%�;g��;�u�;|4�;(�;��;��;��;�"�;In�;�ٓ;�g�; �;��;��u;pj;��^;[�S;��H;o(>;��3;5�);� ;�;`1;�;O��:�[�:5��:�e�:%��:[f�:Ţ�:�X�:�u::.Z:@:ղ&:A�:��9"�9���9`l99�d�8�l�۹���8�j;���ķ�	�
���K��f5�ASK��a��v�Y�����:B���ԥ�i�����2�ź8[к� ۺ���������n����o�Y��W�C��\$��R)�Љ.���3���8���=��B��H�-M�CNR�&yW���\��a��>g���l���q��Ww�S�|�a��8Ń� v��4%���ы�}��5&���Γ�Ww��� ���  �  L�=�P=3�=0�=eK=��=��=�?=�� =ċ =�1 =ӯ�<s��<jL�<��<��<�B�<���<g��<�C�<��<���<�D�<?��<(��<^:�<���<���<� �<�j�<���<���<C�<܊�<	��<�<�_�</��<���<�0�<�s�<`��<���<�0�<j�<���<x��<I��<)�<�N�<q�<���<a��<��<���<���<��<���<�</�<���<���<���< ��<N��<�o�<X7�<h��<ݦ�<�N�<x��<��<�	�<��<��<�p�<���<�6�<��<�߿<�)�<\m�</��<��<e�<�9�<
]�<z�<h��<9��<$��<���<���<���<s��<½�<��<㷝<���<m��<>��<��<ȧ�<ѣ�<���<���<X��<���<�|�<to�<x`�<�O�<|~<LVz<�/v<br<n�m<t�i<іe<ta<3S]<F4Y<�U<&�P<u�L<E�H<�D<t�@<=v<<Z8<-=4<�0<�,<�'<��#<�<e�<x�<-�<E�<��<V�<j�<��;Q;�;���;��;���;T*�;���;�u�;2�;l �;�;�ٮ;H�;e�;y`�;�ʓ;�W�;9	�;t��;�u;�j;3�^;'|S;��H;�>;��3;��);( ;u�;3<;�-;ӵ�:���:���:��:�:���::�:��:��u:��Z:��@:�':;:���9���9��9k�99V��82>E��ߺ���9��hl��b�幡k	����G�5���K�K�a��w��>���ݐ�Gq��?���0������G�ź�^к�ۺ���'�𺂻��Z����\S����'6�$��4�#�X0)��g.���3�g�8���=�`�B��H�bM�ER��tW���\���a�NHg�l�l�+r��mw���|�� ��|ԃ�O����5��Y⋻v����4���ۓ�����Y*���  �  "�=�O=��=�=�K=��=��=eA=�� =ɍ =�3 =��<��<�Q�<���<���<H�<���<���<�G�<H��<x��<�F�<p��<���<:�<���<���<;�<ig�<���<^��<�>�<���<���<��<�Z�<0��<C��<�,�<fp�<���<t��</�<yi�<���<Q��<� �<c+�<�Q�<�t�<���< ��<H��<���<��<���<!�<2	�<��<��<��<���<^��<˟�<�p�<K7�<���<b��<�L�<w��<>|�<c�<7��<S��<k�<���<I1�<e��<�ڿ<3%�<0i�<���<�ݸ<<�<s8�<p\�<*z�<L��<ͤ�<���<ɻ�<`��<ĥ<Kģ<�¡<��<���<,��<Ͷ�<j��<Я�<�<X��<�<#��<ڒ�<���<�|�<�n�<�^�<�M�<v~<Oz<'v<��q<7�m<��i<
�e<>ia<�H]<}*Y<3U<��P<�L<g�H<��D<��@<�u<<[8<�?4<�#0<�,<��'<��#<��<̯<q�<��<�<�<j�<��<��;�K�;���;O"�;,��;00�;W��;�u�;6/�;I��;;ٵ;�ͮ;ܧ;��;N�;��;�C�;��;̀;��u;�i;&{^;�aS;^�H;}>;�3;	�);� ;E�;�I;�@;5��:���:K�:P��:�;�::�:�C�:��::=v:Z[:$-A:(�':2�:e�9��9i�9�L:9��8�c��� ����:��n��fF����湧�	��a �M�6���L�0=b���w�G����%������1��1����6��W�źYdк�ۺ��庍�𺍒��[@� ���/�#����wk���#�)��<.��j3��8��=���B���G�yM��9R�2oW�L�\���a��Tg�T�l�r���w�_�|��3���胻����K������ࠎ��G���쓻/����6���  �  ��=�N=5�=��=L=M�=�=�B=�� =� =�6 =���<	�<iX�<��<���<%N�<?��<��<$L�<��<o��<�H�<���<��<�9�<h��<���<7�<�c�<3��<;��<�8�<��<^��<W�<]T�<R��<���<�'�<Kl�<-��<���<�-�<�h�<П�<5��<��<�-�<aU�<�x�<���<���<.��<1��<���<�<q
�<�<f�<��<D��<J��<���<~��<uq�<F7�<���<���<�I�<���<�w�<M �<��<*��<�d�<5��<�*�<��<�Կ<��<2d�<l��<;ڸ<��<�6�<�[�<Ez�<5��<���<*��<J��<�ŧ<�ȥ<�ɣ<�ȡ<�Ɵ<ĝ<���<��<K��<:��<���<|��<B��<���<���<���<�|�<�m�<!]�<�J�<o~<�Fz< v<��q<.�m<�i<!e<|\a<�<]<Y<�U<��P<��L<l�H<_�D<�@<u<<>\8<�B4<�(0<�,<��'<�#<G�<��<:�<լ<r�<_�<4�<��<^ <_�;2��;n/�;)��;�6�;���;u�;)+�;��;dε;&��;˧;M�;a8�;ܟ�;-+�;e܆;i��;�hu;�i;OV^;�BS;zH;N�=;Կ3;L�);� ;��;�X;�V;� �:�	�:9l�:�F�:���:�h�:d��:�b�:�
w:o\:��A:�H(:M;:�F�9�ʼ9�9��:9�8�q��U���]�;��?��>F�����"�
��!�]T7��MM�	c���x��膺�x������n���ⰺ>[���ź�mк�ۺ���4��d���"����Q��t���
8���#��(��
.��;3��d8�-�=��B���G��L��,R�`iW�E�\�b��cg�u�l�%:r���w�!}��I��� �������d�����与��]��� �������D���  �  "�=�M=��=Ȣ=FL=	�=�=�D=�� =�� =j9 =���<��<N_�<��<��<�T�<K��<���<�P�<��<~��<�J�<���<^��<�8�<��<��<��<|_�<A��<���<�2�<y�<���<��<�M�<��<���<e"�<�g�<r��<��<�+�<�g�<���<��<j�<�0�<�X�<:}�<���<d��<e��<���<l��<��<!�<Q�<-�<��<���<���<���<8��<$r�<7�<x��<u��<�F�<���<*s�<���<Zy�<`��<�]�<��<`#�<�{�<�Ϳ<��<�^�<ȝ�<eָ<��<�4�<{Z�<5z�<	��<���<緫<�©<'ʧ<-Υ<�ϣ<Pϡ<�͟<�ʝ<�Ǜ<�Ù<~��<�<Ƶ�<ί�<���<G��<-��<8��<d|�<�l�<[�<�G�<Rg~<(=z<=v<��q<�m<��i<Cqe<�Na<M/]<�Y<��T<��P<c�L<ܴH<ǟD<>�@<t<<]8<zE4<c-0<J,<L�'<�#<��<&�<��<�<��<��<��<��<� <xs�;G��;=�;���;�<�;A��;�s�;{&�;~�;+µ;���;���;�ܠ;} �;ц�;L�;*;Ӛ�;7u;��i;�-^;A S;�]H;�=;Z�3;a�);L ;M�;�h;Zm;�Z�:JR�:���:��:� �:�զ:��:"҉:��w:��\:R�B:��(:K�:X0�9O�9�]�9�A;9��8|�𵴂���E=��'���a��OJ鹾c���!��(8��'N���c�Zy�N��Eԑ�pI�������������ź�yк�ۺ*���k��4���p�9���D����T�ER#�Θ(���-�m
3��78�Sa=�,�B���G���L�R R��dW���\��b�Ytg���l�gYr���w�pL}��a�����Eφ�����+���Ҏ�rv�����ҵ���T���  �  ��=rL=��=��=�L=��=:�=/F=�� =�� =/< =��<'�<f�<ٶ�<��<[�<T��<��<�U�<��<��<�L�<!��<���<S8�<C��<���<s�<3[�<=��<���<�,�<gr�<���<���<�F�<z��<���<�<c�<���<��<�)�<xf�<���<���<
�<73�<a\�<���<���<��<���<h��<$�<��<��<��<��<��<��<3��<��<¤�<�r�<�6�<D��<4��<�C�<���<?n�<#��<s�<���<WV�<���<�<�t�<=ǿ<W�<PY�<��<�Ҹ<��<�2�<cY�<z�<ה�<.��<���<wƩ<�Χ<Vӥ<�գ<�ա<9ԟ<�ѝ<DΛ<Iʙ<�ŗ<���<���<��<��<���<���<劉<|�<fk�<�X�<�D�<__~<�3z<5v<[�q<��m<��i<6ce<�@a<�!]<Y<2�T<��P<��L<0�H<��D<2�@<�r<<�]8<H4<�10<�,<l(<��#<��<��<�<��<��<t�<4�<+�<M <\��;��;dJ�;��;C�;���;�r�;D!�;t�;뵵;ڠ�;���;BǠ;��;Sm�;���;���;���;�u;�\i;^;��R;qAH;8�=;(�3;S�); ;�;�v;�;Ĕ�:֘�:�:��:�g�:�?�:2��:�?�:��x:n�]:�XC:��):�Z:	�9,�9�͍9�;9�ݸ8tv��z���>����7�����&!��"��9��O��d��0z������0��Қ��N����Q��D����ƺޅк�
ۺ���4M�������K����	��s����#��b(�U�-���2��
8�:=�.iB�b�G��L��R��_W�۶\�-b���g���l�byr���w�ox}�z���4���ꆻ����!G��*펻鎑�-��Sɖ�ae���  �  ��=KK="�=>�=�L=O�=@�=�G=�� =/� =�> =���<-�<Ql�<7��<��<a�<ʳ�<��<�Y�<\��<7��<�N�<&��<���<�7�<���<��<,�<W�<}��<u��<�&�<l�<4��<��<u@�<h��<X��<�<�^�<��<<��<�'�<Ve�<+��<l��<~�<�5�<~_�<\��<T��<M��<h��<t��<w�<�<��<R!�<�<�<��<G��<O��<#��<^s�<G6�<���<��<�@�<��<�i�<���<$m�<J��<�O�<յ�<2�<$n�<���<~�<"T�<x��<�θ<��<�0�<;X�<�y�<���<���<���<�ɩ<�ҧ<إ<�ڣ<wۡ<Wڟ<؝<�ԛ<ZЙ<q˗<�ŕ<O��<˷�<'��<<��<c��<�{�<#j�<�V�<�A�<�W~<{*z<��u<��q<��m<�{i<Ve<�3a<A]<K�X<t�T<6�P<��L<��H<ܕD<�@<�q<<]^8<[J4<�50<�!,<�(<��#<7�<,�<m�<��< �<W�<��<�	<�' <���;4��;�V�;���;`H�;/��;�p�;�;�ؼ;��;���;ٓ�;���;��;(U�;�݌;���;�g�;/�t;T1i;��];0�R;�%H;�=;K�3;��);x ;�;|�;��;���:K��:^�:6W�:�Ķ:R��:�:o��:�~y:�m^:^D:�.*:��:7��9=ɾ9(2�9+<9 ��8��7�7hø`@�����~���!�����?t#���9���O��e���z�c�������眺R<������׻�F.ƺ}�к2ۺ��41�i������Z*�Њ�����D������"�I0(��p-�I�2���7�=�wKB���G���L�q
R�}\W���\��#b���g��m�)�r�Ox���}� ���9M���������a��������B���ۖ�%u���  �  ��=NJ=z�=��=�L=��=�=�H=� =� =�@ =i��<L!�<�q�<���<�<f�<���<�<_]�<M��<h �<UP�<מ�<���<�6�<,��<���<9�<�S�<U��<���<u!�<�f�<���<f��<;�<��<l��<��<�Z�<Ѡ�<���<&�<@d�<��<���<��<p7�<b�<���<3��<���<J��<���<��<B�<�"�<1&�<�#�<Z�<
�<���<&��<1��<�s�<�5�<���<��<>�<���<�e�<:��<�g�<���<�I�<گ�<K�<nh�<j��<m�<�O�<���<�˸<K �<�.�<(W�<py�<㕯<ᬭ<澫<^̩<�է<ܥ<eߣ<f�<�ߟ<Gݝ<�ٛ<�ՙ<MЗ</ʕ< Ó<��<���<æ�<��<���<D{�<�h�<�T�<B?�<(Q~<�"z<��u<��q<Ùm<{pi<vJe<�(a<Y
]<��X<�T<��P<ɲL<��H<��D<P�@<Np<<�^8<L4<!90<9&,<�(<C$<�<��<��<��<��<d�<�<�<�0 <ب�;��;d`�;���;<L�;u��;�n�;>�;@Ѽ;F��;���;9��;堠;�ޙ;�@�;�Ȍ;�x�;�R�;v�t;�i;¼];z�R;�H;G�=;|�3;�);c ; �;A�;��;���:l�:���:[��:&�:���:�E�:���:I(z:�_:#�D:�*:8F:y��9�H�9B��9_R<9�q�8RW�bŸ�EA�����h���[�칍o��$�q|:�$�P��Af�S�{��c���Ԓ�z+��hu���������Fƺ��к�ۺ�庼𺣺��ȳ�J��i������p�?�"��(��G-���2�Ծ7���<�2B�6pG�شL��R��ZW�}�\��-b���g�W*m���r��<x�"�}�����b�����p̉�	w��t��G����T���떻�����  �  ��=�I=��=��=�L=�=��=�I=D� =q� =}B =��<+%�<�u�<���<#�<�i�<��<#�<`�<���<�<�Q�<c��<���<:6�<�~�<*��<��<�P�<
��<6��<��<zb�<Q��<��<�6�<�<���<'�<�W�<V��<���<�$�<Wc�<���<��<�	�<�8�<d�<.��<#��<'��<���<���<��<]�<�&�<�)�<�&�<G�<��<���<���<��<�s�<�5�<���<���<�;�<��<�b�<���<d�<j��<ZE�<:��<�
�<�c�</��<��<L�<���<�ȸ<H��<\-�<IV�<.y�<1��<ح�<[��<jΩ<pا<ߥ<��<�<��<f�<�ݛ<oٙ<�ӗ<�͕<
Ɠ<���<���<-��<<勉<�z�<�g�<WS�<+=�<	L~<mz<��u<�q<V�m<�gi<�Ae<�a<�]<�X<��T<y�P<Z�L<m�H<T�D<	@<Ko<<�^8<NM4<�;0<�),<�(<�$<��<T�<��<-�<��<��<	<�<<7 <���;��;�g�;P��;FO�;C��;gm�;P�;˼;���;qz�;�w�;|��;�ϙ;T0�;׷�;�g�;�B�;�t;=�h;S�];ԧR;��G;f�=;�|3;��);  ;�;G�;�;p�:H8�:���:t��:�O�:S7�:f��:�>�:��z:�_:�E:f+:ϙ:��9M��9ӿ�9�}<9�C�8:�q�kpƸ�9B��Z���B�����"��G�$��;�}Q��f�R0|��������a��֡��!ݱ�����Zƺ@�к�ۺg�庺�����^�����CQ�w������O��"���'�R(-��g2�p�7���<�{B�?aG���L���Q�kYW���\��5b��g�E;m�(�r��Ux�#�}�7���Ds���+��މ�>���D,���ɑ��b��n�������  �  ܛ=�H=��=��=�L=N�=�=BJ=�� =[� =�C =G��<�'�<;x�<=��<��<Zl�<C��<)�<�a�<۲�<�<+R�<���<���<�5�<>~�<��<�
�<O�<���<���<��<�_�<���<W��<
4�<d|�<G��<��<V�<���<���<�#�<�b�<_��<:��<
�<�9�<;e�<���<��<?��<D��<�<U�<� �<J)�<.,�<)�<1�<�<���<]��<���<�s�<>5�<0��<���<�:�<k��<�`�<M��<�a�<���<�B�<i��<��<a�<w��<�<�I�<���<aǸ<
��<p,�<�U�<�x�<c��<[��<B��<�ϩ<ڧ<��<��<��<�<��<}��<�ۙ<@֗<�ϕ<�Ǔ<���<���<���<p��<���<�z�<dg�<dR�<�;�<�H~<�z<)�u<�q<�m<\bi<,<e<Ja<f�\<��X<�T<c�P<թL<H<6�D<�}@<vn<<�^8<)N4<=0< ,,<�(<�$<��<��<��<J�<��<��<.
<�<�; <���;��;�l�;k��;<Q�;Q��;!l�;��;_Ǽ;���;�s�; p�;���;	ƙ;&�;w��;�]�;!8�;�zt;U�h;g�];-�R;��G;U�=;\v3;�);� ;ߴ;�;��;A(�:�Q�:��:���:�u�:�^�:��:�g�:	�z:��_:_HE:}M+:1�:�e�9e�9$�9�<9�8����"OǸv�B�G���G���>S��1�B�$�Z;��kQ�&#g���|��̈��3��g�������1���^)��zgƺ�к|ۺ�}�������.��a��0A�������<���"���'��-�EU2��7�'�<�=B�LXG��L���Q��XW�D�\��:b�ۻg�JEm���r�2ex�>�}�7����}��6���艻	����6���ӑ��k��a ��쓙��  �  ��=�H=�=��=�L=^�=0�={J=5� =�� =�C =��<{(�<y�<��<w�<8m�<��<��<ib�<Z��<��<NR�<۟�<���<�5�<�}�<���<�	�<fN�<`��<��<0�<�^�<���<D��<3�<�{�<~��<D�<jU�<��<
��<S#�<�b�<J��<G��< 
�<�9�<�e�<=��<���<���<��<��<'�<�!�<%*�<-�<�)�<��<��<n��<���<���<t�<%5�<��<9��<:�<���<�_�<���<�`�<���<�A�<K��<��<2`�<���<?�<I�<抺<�Ƹ<���<,�<�U�<�x�<s��<s��<���<Щ<�ڧ<��<��<a�<��<��<Q�<�ܙ<ח<=Е<�ȓ<}��<4��<.��<���<	��<�z�<1g�<�Q�<l;�<bG~<Iz<��u<��q<t�m<^`i<�9e<<a<��\<\�X<��T<�P<w�L<��H<U�D<}@<7n<<�^8<dN4<{=0<�,,<�(<�$< <z�<��<��<��<��<�<!<�< <u��;��;Xn�;&��;�Q�;���;�k�;��;�ż;ҏ�;Lq�;�m�;���;
Ù;�"�;r��;fY�;�4�;�tt;M�h;:�];d�R;��G;��=;�s3;ϟ); ;m�;ߚ;0�;~0�:KZ�:���:R�:p��:�l�:y��:u�:�{:��_:r]E:a+:��:���9d��9��9��<9/��8M4����ǸC��䐹9俹~�K��
%��w;�׍Q��Dg�T�|�Cو�5@��l����ɧ������0��dlƺ��к�ۺ�{����ފ��;�����R<�������(5�y�"�&�'��-�O2�؎7�%�<�B�~TG�L�L��Q��XW�%�\�o<b��g�fIm���r�'jx���}�\���ꀄ�r:��퉻���:���֑��n����������  �  ܛ=�H=��=��=�L=N�=�=BJ=�� =[� =�C =G��<�'�<;x�<=��<��<Zl�<C��<)�<�a�<۲�<�<+R�<���<���<�5�<>~�<��<�
�<O�<���<���<��<�_�<���<W��<
4�<d|�<G��<��<V�<���<���<�#�<�b�<_��<:��<
�<�9�<;e�<���<��<?��<D��<�<U�<� �<J)�<.,�<)�<1�<�<���<]��<���<�s�<>5�<1��<���<�:�<k��<�`�<M��<�a�<���<�B�<i��<��<a�<w��<�<�I�<���<aǸ<
��<p,�<�U�<�x�<c��<[��<B��<�ϩ<ڧ<��<��<��<�<��<}��<�ۙ<@֗<�ϕ<�Ǔ<���<���<���<p��<���<�z�<dg�<dR�<�;�<�H~<�z<)�u<�q<�m<\bi<,<e<Ja<g�\<��X<�T<c�P<թL<H<6�D<�}@<vn<<�^8<)N4<=0< ,,<�(<�$<��<��<��<J�<��<��<-
<�<�; <���;��;�l�;k��;<Q�;Q��;!l�;��;_Ǽ;���;�s�; p�;���;	ƙ;&�;w��;�]�; 8�;�zt;U�h;g�];-�R;��G;U�=;\v3;�);� ;ߴ;�;��;A(�:�Q�:��:���:�u�:�^�:��:�g�:	�z:��_:_HE:}M+:1�:�e�9e�9$�9�<9�8����"OǸv�B�G���G���>S��1�B�$�Z;��kQ�&#g���|��̈��3��g�������1���^)��zgƺ�к|ۺ�}�������.��a��0A�������<���"���'��-�EU2��7�'�<�=B�LXG��L���Q��XW�D�\��:b�ۻg�JEm���r�2ex�>�}�7����}��6���艻	����6���ӑ��k��a ��쓙��  �  ��=�I=��=��=�L=�=��=�I=D� =q� =}B =��<+%�<�u�<���<#�<�i�<��<#�<`�<���<�<�Q�<c��<���<:6�<�~�<*��<��<�P�<
��<6��<��<zb�<Q��<��<�6�<�<���<'�<�W�<V��<���<�$�<Wc�<���<��<�	�<�8�<d�<.��<#��<'��<���<���<��<]�<�&�<�)�<�&�<G�<��<���<���<��<�s�<�5�<���<���<�;�<��<�b�<���<d�<j��<ZE�<:��<�
�<�c�</��<��<L�<���<�ȸ<H��<]-�<IV�</y�<1��<ح�<[��<jΩ<pا<ߥ<��<�<��<f�<�ݛ<oٙ<�ӗ<�͕<
Ɠ<���<���<-��<<勉<�z�<�g�<WS�<*=�<	L~<mz<��u<�q<V�m<�gi<�Ae<�a<�]<�X<��T<y�P<Z�L<m�H<T�D<	@<Ko<<�^8<NM4<�;0<�),<�(<�$<��<T�<��<-�<��<��<	<�<<7 <���;��;�g�;O��;FO�;C��;fm�;O�;˼;���;qz�;�w�;|��;�ϙ;S0�;׷�;�g�;�B�;�t;<�h;R�];ӧR;��G;e�=;�|3;��);  ;�;G�;�;p�:H8�:���:t��:�O�:S7�:f��:�>�:��z:�_:�E:f+:ϙ:��9M��9ӿ�9�}<9�C�8:�q�kpƸ�9B��Z���B�����"��G�$��;�}Q��f�R0|��������a��֡��!ݱ�����Zƺ@�к�ۺg�庺�����^�����CQ�w������O��"���'�R(-��g2�p�7���<�{B�?aG���L���Q�kYW���\��5b��g�E;m�(�r��Ux�#�}�7���Ds���+��މ�>���D,���ɑ��b��n�������  �  ��=NJ=z�=��=�L=��=�=�H=� =� =�@ =i��<L!�<�q�<���<�<f�<���<�<_]�<M��<h �<UP�<מ�<���<�6�<,��<���<9�<�S�<U��<���<u!�<�f�<���<f��<;�<��<l��<��<�Z�<Ѡ�<���<&�<@d�<��<���<��<p7�<b�<���<3��<���<J��<���<��<B�<�"�<1&�<�#�<Z�<
�<���<&��<1��<�s�<�5�<���<��<>�<���<�e�<;��<�g�<���<�I�<گ�<K�<nh�<k��<m�<�O�<���<�˸<K �<�.�<)W�<qy�<㕯<ᬭ<澫<^̩<�է<ܥ<eߣ<f�<�ߟ<Gݝ<�ٛ<�ՙ<MЗ<.ʕ< Ó<��<���<¦�<��<���<D{�<�h�<�T�<A?�<(Q~<�"z<��u<��q<Ùm<{pi<uJe<�(a<Y
]<��X<�T<��P<ʲL<��H<��D<Q�@<Op<<�^8<L4<!90<9&,< (<C$<�<��<��<��<��<c�<�<�<�0 <ب�;��;c`�;���;;L�;t��;�n�;=�;?Ѽ;E��;���;8��;䠠;�ޙ;�@�;�Ȍ;�x�;�R�;t�t;�i;��];y�R;�H;F�=;{�3;�);c ; �;@�;��;���:k�:���:[��:&�:���:�E�:���:I(z:�_:#�D:�*:8F:y��9�H�9B��9_R<9�q�8RW�bŸ�EA�����h���[�칍o��$�q|:�$�P��Af�S�{��c���Ԓ�z+��hu���������Fƺ��к�ۺ�庼𺣺��ȳ�J��i������p�?�"��(��G-���2�Ծ7���<�2B�6pG�شL��R��ZW�}�\��-b���g�W*m���r��<x�"�}�����b�����p̉�	w��t��G����T���떻�����  �  ��=KK="�=>�=�L=O�=@�=�G=�� =/� =�> =���<-�<Ql�<7��<��<a�<ʳ�<��<�Y�<\��<7��<�N�<&��<���<�7�<���<��<,�<W�<}��<u��<�&�<l�<4��<��<u@�<h��<X��<�<�^�<��<<��<�'�<Ve�<+��<l��<~�<�5�<~_�<\��<T��<M��<h��<t��<w�<�<��<R!�<�<�<��<G��<O��<#��<^s�<G6�<���<��<�@�<��<�i�<���<%m�<K��<�O�<յ�<2�<$n�<���<~�<"T�<x��<�θ<��<�0�<;X�<�y�<���<���<���<�ɩ<�ҧ<إ<�ڣ<wۡ<Wڟ<؝<�ԛ<ZЙ<q˗<�ŕ<N��<ʷ�<'��<<��<c��<�{�<"j�<�V�<�A�<�W~<z*z<��u<��q<��m<�{i<Ve<�3a<A]<K�X<t�T<6�P<��L<��H<ݕD<�@<�q<<^^8<\J4<�50<�!,<�(<��#<7�<,�<m�<��< �<W�<��<�	<�' <���;3��;�V�;���;_H�;-��;�p�;�;�ؼ;��;���;ؓ�;���;��;'U�;�݌;���;�g�;.�t;S1i;��];/�R;�%H;�=;J�3;��);w ;�;|�;��;���:K��:^�:6W�:�Ķ:R��:�:o��:�~y:�m^:^D:�.*:��:6��9=ɾ9(2�9+<9 ��8��7�7hø`@�����~���!�����?t#���9���O��e���z�c�������眺R<������׻�F.ƺ}�к2ۺ��41�i������Z*�Њ�����D������"�I0(��p-�I�2���7�=�wKB���G���L�q
R�}\W���\��#b���g��m�)�r�Ox���}� ���9M���������a��������B���ۖ�%u���  �  ��=rL=��=��=�L=��=:�=/F=�� =�� =/< =��<'�<f�<ٶ�<��<[�<T��<��<�U�<��<��<�L�<!��<���<S8�<C��<���<s�<3[�<=��<���<�,�<gr�<���<���<�F�<z��<���<�<c�<���<��<�)�<xf�<���<���<
�<73�<a\�<���<���<��<���<h��<$�<��<��<��<��<��<��<3��<��<ä�<�r�<�6�<D��<4��<�C�<���<?n�<#��<s�<���<WV�<���<�<�t�<=ǿ<X�<PY�<��<�Ҹ<��<�2�<cY�<z�<ؔ�<.��<���<xƩ<�Χ<Vӥ<�գ<�ա<9ԟ<�ѝ<DΛ<Iʙ<�ŗ<���<���<��<��<���<���<劉<|�<fk�<�X�<�D�<__~<�3z<4v<Z�q<��m<��i<6ce<�@a<�!]<Y<2�T<��P<��L<1�H<��D<2�@<�r<<�]8<H4<�10<�,<l(<��#<��<��<�<��<��<t�<3�<*�<M <[��;��;cJ�;��; C�;���;�r�;B!�;r�;굵;٠�;���;AǠ;��;Rm�;���;���;���;�u;�\i;^;��R;pAH;7�=;'�3;S�); ;�;�v;�;Ĕ�:֘�:�:��:�g�:�?�:2��:�?�:��x:n�]:�XC:��):�Z:	�9,�9�͍9�;9�ݸ8uv��z���>����7�����&!��"��9��O��d��0z������0��Қ��N����Q��D����ƺޅк�
ۺ���4M�������K����	��s����#��b(�U�-���2��
8�:=�.iB�b�G��L��R��_W�۶\�-b���g���l�byr���w�ox}�z���4���ꆻ����!G��*펻鎑�-��Sɖ�ae���  �  "�=�M=��=Ȣ=FL=	�=�=�D=�� =�� =j9 =���<��<N_�<��<��<�T�<K��<���<�P�<��<~��<�J�<���<^��<�8�<��<��<��<|_�<A��<���<�2�<y�<���<��<�M�<��<���<e"�<�g�<r��<��<�+�<�g�<���<��<j�<�0�<�X�<:}�<���<d��<e��<���<l��<��<!�<Q�<-�<��<���<���<���<8��<$r�<7�<y��<u��<�F�<���<*s�<���<Zy�<`��<�]�<��<`#�<�{�<�Ϳ<��<�^�<ȝ�<fָ<��<�4�<{Z�<5z�<
��<���<緫<�©<'ʧ<-Υ<�ϣ<Pϡ<�͟<�ʝ<�Ǜ<�Ù<}��<�<Ƶ�<ͯ�<���<F��<-��<8��<d|�<�l�<[�<�G�<Rg~<(=z<<v<��q<�m<��i<Cqe<�Na<M/]<�Y<��T<��P<d�L<ݴH<ȟD<?�@<t<< ]8<{E4<c-0<K,<M�'<�#<��<'�<��<�<��<��<��<��<� <ws�;F��;=�;���;�<�;?��;�s�;y&�;|�;*µ;���;���;�ܠ;| �;І�;K�;);Қ�;�6u;��i;�-^;@ S;�]H;�=;Y�3;a�);L ;M�;�h;Zm;�Z�:IR�:���:��:� �:�զ:��:"҉:��w:��\:Q�B:��(:K�:X0�9O�9�]�9�A;9��8}�𵴂���E=��'���a��OJ鹾c���!��(8��'N���c�Zy�N��Eԑ�pI�������������ź�yк�ۺ*���k��4���p�9���D����T�ER#�Θ(���-�m
3��78�Sa=�,�B���G���L�R R��dW���\��b�Ytg���l�gYr���w�pL}��a�����Eφ�����+���Ҏ�rv�����ҵ���T���  �  ��=�N=5�=��=L=M�=�=�B=�� =� =�6 =���<	�<iX�<��<���<%N�<?��<��<$L�<��<o��<�H�<���<��<�9�<h��<���<7�<�c�<3��<;��<�8�<��<^��<W�<]T�<R��<���<�'�<Kl�<-��<���<�-�<�h�<П�<5��<��<�-�<aU�<�x�<���<���<.��<1��<���<�<q
�<�<f�<��<D��<J��<���<~��<uq�<F7�<���<���<�I�<���<�w�<M �<��<*��<�d�<6��<�*�<���<�Կ<��<3d�<m��<<ڸ<��<�6�<�[�<Ez�<6��<���<*��<J��<�ŧ<�ȥ<�ɣ<�ȡ<�Ɵ<ĝ<���<��<K��<:��<���<|��<B��<���<���<���<�|�<�m�<!]�<�J�<o~<�Fz< v<��q<.�m<�i<!e<|\a<�<]<Y<�U<��P<��L<l�H<`�D<�@<u<<>\8<�B4<�(0<�,<��'<�#<G�<��<:�<լ<r�<_�<3�<��<^ <_�;1��;m/�;(��;�6�;���;u�;(+�;��;bε;%��;˧;L�;`8�;۟�;,+�;d܆;i��;hu;	�i;NV^;�BS;zH;M�=;Կ3;L�);� ;��;�X;�V;� �:�	�:9l�:�F�:���:�h�:d��:�b�:�
w:o\:��A:�H(:M;:�F�9�ʼ9�9��:9�8�q��U���]�;��?��>F�����"�
��!�]T7��MM�	c���x��膺�x������n���ⰺ>[���ź�mк�ۺ���4��d���"����Q��t���
8���#��(��
.��;3��d8�-�=��B���G��L��,R�`iW�E�\�b��cg�u�l�%:r���w�!}��I��� �������d�����与��]��� �������D���  �  "�=�O=��=�=�K=��=��=eA=�� =ɍ =�3 =��<��<�Q�<���<���<H�<���<���<�G�<H��<x��<�F�<p��<���<:�<���<���<;�<ig�<���<^��<�>�<���<���<��<�Z�<0��<C��<�,�<fp�<���<t��</�<yi�<���<Q��<� �<c+�<�Q�<�t�<���< ��<H��<���<��<���<!�<2	�<��<��<��<���<^��<˟�<�p�<L7�<���<b��<�L�<w��<>|�<c�<7��<S��<k�<���<I1�<e��<�ڿ<3%�<0i�<���<�ݸ<=�<s8�<p\�<*z�<M��<Τ�<���<ɻ�<`��<ĥ<Lģ<�¡<��<���<,��<Ͷ�<j��<Я�<�<X��<�<#��<ڒ�<���<�|�<�n�<�^�<�M�<v~<Oz<'v<��q<7�m<��i<
�e<>ia<�H]<}*Y<3U<��P<�L<h�H<��D<��@<�u<<[8<�?4<�#0<�,<��'<��#<��<̯<q�<��<�<�<j�<��<��;�K�;���;N"�;+��;/0�;U��;�u�;5/�;H��;:ٵ;�ͮ;ܧ;��; N�;��;�C�;��;̀;��u;�i;%{^;�aS;^�H;}>;
�3;	�);� ;D�;�I;�@;5��:���:K�:P��:�;�::�:�C�:��::=v:Z[:$-A:(�':2�:e�9��9i�9�L:9��8�c��� ����:��n��fF����湧�	��a �M�6���L�0=b���w�G����%������1��1����6��W�źYdк�ۺ��庍�𺍒��[@� ���/�#����wk���#�)��<.��j3��8��=���B���G�yM��9R�2oW�L�\���a��Tg�T�l�r���w�_�|��3���胻����K������ࠎ��G���쓻/����6���  �  L�=�P=3�=0�=eK=��=��=�?=�� =ċ =�1 =ӯ�<s��<jL�<��<��<�B�<���<g��<�C�<��<���<�D�<?��<(��<^:�<���<���<� �<�j�<���<���<C�<܊�<	��<�<�_�</��<���<�0�<�s�<`��<���<�0�<j�<���<x��<I��<)�<�N�<q�<���<a��<��<���<���<��<���<�</�<���<���<���< ��<N��<�o�<X7�<h��<ݦ�<�N�<x��<��<�	�<��<��<�p�<���<�6�<��<�߿<�)�<\m�<0��<��<f�<�9�<
]�<z�<h��<:��<%��<���<���<���<s��<½�<��<㷝<���<m��<>��<��<ȧ�<ѣ�<���<�<X��<���<�|�<to�<x`�<�O�<|~<LVz<�/v<br<n�m<t�i<іe<ta<3S]<G4Y<�U<&�P<u�L<E�H<�D<t�@<>v<<Z8<.=4<�0<�,<�'<��#<�<e�<x�<-�<E�<��<V�<j�<��;P;�;���;��;���;S*�;���;�u�;2�;k �;
�;�ٮ;G�;d�;x`�;�ʓ;�W�;8	�;s��;�u;�j;2�^;&|S;��H;�>;��3;��);( ;u�;3<;�-;ӵ�:���:���:��:�:���::�:��:��u:��Z:��@:�':;:���9���9��9k�99V��84>E��ߺ���9��hl��b�幡k	����G�5���K�K�a��w��>���ݐ�Gq��?���0������G�ź�^к�ۺ���'�𺂻��Z����\S����'6�$��4�#�X0)��g.���3�g�8���=�`�B��H�bM�ER��tW���\���a�NHg�l�l�+r��mw���|�� ��|ԃ�O����5��Y⋻v����4���ۓ�����Y*���  �  .�=/Q=��=7�=(K=V�=�=�>=�� =+� =�/ =���<<��<H�<{��<���<�>�<ɓ�<���<�@�<v��<���<,C�<@��<���<�:�<���<���<�"�<m�<q��<��<"G�<ˎ�<(��<)�<�c�<��<h��<�3�<�v�<���<��<�1�<�j�<���<���<��<K'�<�L�<>n�<'��<Ѧ�<��<K��<:��<���<���< �<� �<e��<���<���<[��<��<:o�<U7�<���<��<�P�<���<���<��<ȍ�<��<�t�<���<J;�<$��<��<�-�<�p�<���<��<�<�:�<x]�<�y�<���<�<E��<^��<Ӻ�<W��<ӻ�<���<޶�<���<S��<0��<Q��<���<z��<��<���<1��<!��<Y��<�|�<�o�<�a�<�Q�<��~<�[z<�5v<�r<#�m<��i<<�e<f|a<[]<�;Y<�U<� Q<T�L<��H<ƮD<ޒ@<zv<<,Y8<;4<�0<u�+<��'<	�#<�<��<א<R�<2�<З<��<��<M��;;.�;���;n�;���;�%�;f��;�u�;{4�;'�;��;��;��;�"�;Hn�;�ٓ;�g�;�;��;��u;pj;��^;Z�S;��H;o(>;��3;5�);� ;�;`1;�;O��:�[�:5��:�e�:%��:[f�:Ţ�:�X�:�u::.Z:@:ղ&:A�:��9"�9���9`l99�d�8�l�۹���8�j;���ķ�	�
���K��f5�ASK��a��v�Y�����:B���ԥ�i�����2�ź8[к� ۺ���������n����o�Y��W�C��\$��R)�Љ.���3���8���=��B��H�-M�CNR�&yW���\��a��>g���l���q��Ww�S�|�a��8Ń� v��4%���ы�}��5&���Γ�Ww��� ���  �  ��=�Q=��=4�=�J=��=_�=9>=�� =+� =�. =q��<���<iE�<ԕ�<��<�;�<K��<���<�>�<̕�<~��<7B�<���<}��<�:�<��<���<�#�<�n�<N��<,�<qI�<=��<���<��<Rf�<`��<���<�5�<4x�<Ǹ�<��<�2�<�j�<f��<I��<7��<-&�<'K�<il�<��<p��<���<���<���<��<���<u��<@��<L��<���<+��<@��<Q��<�n�<17�<E��<���<�Q�<��<~��<�<��<�<ww�<���<�=�<���<H�<�/�<�r�<���<�<��<�;�<�]�<�y�<3��<��<$��<Ҵ�<���<.��<f��<��<1��<߰�<���<���<ħ�<)��<n��<F��<J��<��<`��<ᆉ<�|�<Yp�<Lb�<�R�<+�~<N_z<�9v<	r<�m<��i<p�e<t�a<`]<8@Y<�!U<�Q<"�L<7�H<I�D<Г@<v<<qX8<�94<�0<��+<<�'<��#<?�<_�<i�<ǅ<��<;�<6�<X�<���;�%�;l��;��;\��;�"�;���;ju�;�5�;��;��;-�;��;�*�;w�;9�;Pq�;�"�;_��;c�u;0j;��^;�S;+�H;�/>;��3;��);�	 ;�{;i*;;;w�:�=�:�~�:?�:�|�:F;�:�w�:�-�:��t:�Y:s�?:�m&:&�:t��9���9�r�9�+99�(�8ڵ�*E��p8�쉹	]�����m��*��L5��K�R�`�Qv�!߅������#������@V��������ź�Xк�$ۺ��2��U���{���ڀ� ��l�����#$��h)�!�.�Q�3�j�8�$�=�C��H�n5M�TR��|W�>�\���a�>9g�t�l�W�q��Iw��|�r	��Y���l�����ȋ�5s��,���Ɠ�#p������  �  D�=mW=� =��=/Q=��=��=�B=�� =G� =/1 =j��<(��< I�<l��<���<E�<ĝ�<���<S�<g��<i	�<0c�<���<��<)f�<C��<_�<�V�<���<z��<�:�<*��<]��<��<�c�<��<~��<-?�<��<P��<��<�S�<��<���<j�<&:�<Yi�<���<y��<���<?��<��<�4�<�K�<�`�<�r�<��<?��<E��<̕�<֐�<c��<@o�<hP�<s'�<N��<��<�h�<��<!��<�D�<���<�L�<M��<�.�<Ò�<x��<IB�<ߎ�<%Ծ<h�<�I�<�z�<l��<yǵ<��<���<u	�<!�<��<��<�<��<v�<G��<�<�<K�<|ۙ<�՗<�Е<�˓<,Ǒ<���<��<���<_��<���<���<z{�<�h�<��~<�{z<�Nv<� r<�m<��i<-�e<oa<�F]<�Y<o�T<d�P<1�L<S�H<lD<H@<�!<<�7<+�3<"�/<�y+<�N'<�%#<Z <K�<��<n�<Ƭ<��
<�<��<���;`,�;��;���;�u�;J��;Ӓ�;"4�;���;y��;Tv�;�]�;h^�;�z�;���;1�;�;�5�;|;��o;x!d;�X;H�M;��B;�8;��-;��#;�;�};>2;`I�:J��:C~�:,��:P��:'�:��:K��:;{:�$`:'F:)�,:Qs:�*�9&h�9�W�9�|]99,�#8g2D���
��ud�C�ׅ˹x��������'�c�=��S�~lh�m�}�YT��O̓�h;�������������Ⱥ�Һ�wݺ{N��@�D��J��8
�����@�C��r ��d%�ћ*��/�l�4���9��>�ѾC�_�H�3�M�űR���W��\�b�iSg�M�l���q�qNw���|���������c��}�����5_��S��먓��M�����  �  ��=KW=� =��=BQ=��=�=(C= � =�� =�1 =���<I��<~J�<���<���<>F�<��<���<�S�<&��<�	�<�c�<Ի�<�<)f�<��<
�<;V�<���<���<�9�<��<B��<A�<*b�<��<b��<@>�<!��<���<0�<rS�<���<���<w�<K:�<�i�<���<��<j��<%��<��<�5�<)M�<b�<-t�<��<i��<^��<���<���< ��<�o�<�P�<�'�<T��<ӳ�<�h�<>�<w��<�C�<���<�K�<��<�-�<T��<��<A�<���<&Ӿ<��<&I�<�y�<���<Gǵ<��<���<�	�<��<>�<e�<��<��<��<f��<T��<��<��<�ܙ<�֗<�ѕ<�̓<ȑ<j<���<��<���<���<���<>{�<h�<_�~<�zz<Mv<�r<��m<x�i<c�e<ma<xD]<�Y<��T<��P<αL<$�H<�kD<�G@<�!<<J�7<��3<�/<�z+<CP'<�'#<�<��<#�<;�<�<S�
<]�<��<���;;0�;H��;��;x�;���;���;`4�;\��;a��;"t�;r[�;�[�;Ow�;|��;��;���;�0�;Y�{;H�o;hd;��X;�|M;�B;s8;x�-;��#;�;";�5;nQ�:v��:���:���:Hȸ:`/�:8"�:E��:�F{:�K`: @F:�-:�:nd�9?��9w�9��]9�!9��#8�?D�+�
�M�d�x����˹���{���'�X�=��=S��h���}�f��#ۓ�uG��򰨺���l����Ⱥ��Һ�uݺ�J�(9�0<������0
�����7�(��A �aX%���*��/�'�4�F�9���>��C�­H�+�M��R�q�W���\�b�`Ug���l��q�PTw�f�|��
��Z���\h���������c��^��Y����P��r����  �  I�=�V=� =��=�Q=|�=��=D=)� =� ==3 =���<���<N�<���<���<�I�<=��<���<�V�<]��<��<e�<���<v�<f�<���<�<�T�<��<R��<�6�<��<
��<��<�^�<���<7��<T;�<���<w��<��<3R�<��<9��<��<�:�<�j�<���<��<���<��<�<G9�<�P�<�e�<�w�<���<��<���<x��<&��<���<Eq�<�Q�<'(�<w��<h��<�g�<��<���<�A�<��<�H�<ǽ�<*�<ʍ�<���<�=�<a��< о<��<G�<;x�<���<qƵ<��<��<N
�<��<��<r�<c�<k�<�	�<� �<���<"�<=�<8��<Dڗ<�ԕ<�ϓ<qʑ<_ď</��<&��<!��<ћ�<-��<lz�<�f�<�~<vz<�Gv<�r<e�m<�i<��e<\fa<�=]<�Y<�T<"�P<�L<8�H< jD<�F@<�!<<2�7<��3<�/<�~+<�T'<	-#<�<��<{�<��<=�<��
<��<��<x��;N;�;Ϙ�;��;M~�;��;ו�;�4�;���;���;�n�;�T�;�R�;�l�;���;� �;J�;�#�;��{;��o; d;�X;�lM;ԖB;O8;��-;��#;�;��;�?;l�:���:ִ�:;�:v��:h�:�[�:jً:�{:��`:��F:�u-:��:��9J�9���9�S^9�z9�($8��D�S��De�񀟹�6̹y����r�ia(��>���S��i�k*~�����U��tn��Ш�6��å��q'Ⱥ��ҺDpݺ�=躎#�5 ��E��T
����j��������;%�/t*�S�/���4���9��>�"�C�z�H�ٜM���R� �W��\��b�2\g�^�l��r�=fw���|����!ǃ�[u��[!��ʋ�mp�����9����Y�������  �  '�=V=M =��=�Q=9�=��=�E=�� =8� =�5 =#��<��<�S�<���<q��<wO�<J��<� �<�Z�<Դ�<��<g�<
��<�<�e�<���<^�<PR�<���<���<�2�<'|�<���<o�<OY�<<��<+��<�6�<}�<��<��<4P�<���<���<��<�;�<�l�<��<O��<���<t�<�#�<�>�<}V�<�k�<�}�<q��<@��<]��<���<���<'��<�s�<�S�<)�<���<ز�<�f�<��<ȫ�<>�<���<�C�<~��<T$�<���<���<�7�<,��<`˾<�
�<�C�<mu�<���<Bŵ<�<W��<\�<t�<q�<��<B�<��<��<h�<���<��<+�<�<�ߗ<�ٕ<ԓ<(Α<�Ǐ<���<ŵ�<��<���<���<y�<�d�<�~<�nz<]?v<hr<��m<��i<k�e<#[a<B3]<�Y<i�T<��P<ۧL<s�H<�fD<$E@<�!<<��7<��3<_�/<��+<+\'<�5#<c<�<6�<��<��<��
<��<y�<N�;�L�;���;]�;Q��;:
�;Q��;G5�;`��;f��;&f�;�H�;�D�;<\�;=��;(�;%j�;��;Z�{;(�o;}�c;JqX;�RM;	�B;��7;|�-;A�#;�	;�;�M;���:��:B��:=^�:�J�:���:���:�9�:Nz|:�za:`G:<.:N�:��9��9%��9�4_9-9e�$8��E����8f��+��5͹h���+�)��>��XT�}�i���~�)扺RO��뫞�e��&^�������5Ⱥ��ҺhݺN)�g����z�.�	�|�N��b�����%��D*�k/���4�"�9��>��C���H���M�A�R�g�W�(�\�(b�\gg���l�Kr���w��|��)���ۃ�a���n7��#���]����'��ȓ�+h���	���  �  ��=U=��=}�=SR=3�=$�=vG=A� =�� =�8 =���<��<n[�<-��<� �<�V�<���<��<�_�<@��<�<�i�<ſ�<��<�e�<Y��<�<O�<Ù�<���<�,�<�u�<ݾ�<U�<&R�<?��<���<�0�<z�<w��<	�<vM�<��< ��<�</=�<�n�< ��<T��<y��<.�<`*�<�E�<�]�<s�<(��<���</��<ǣ�<���<���<#��<�v�<�U�<B*�<���<��<�d�<��<٧�<19�<*��<R=�<���<��<j��<2��<�0�<F~�<ž<C�<�>�<�q�<靷<võ<H�<���<��<��<��<�!�<D �<��<9�<j�<��<���<���<?�<r�<��<�ٓ<�ґ<vˏ<�<뷋<&��<��<���<#w�<�a�<]�~<eez< 4v<�r<u�m<��i<�ve<�La<�%]<� Y<��T<��P<��L<�H<QbD<�B@<5!<<+�7<Z�3<�/<�+<me'<�@#<+<<��<�<f�<5�
<W�<z�<�;Cc�;Ϻ�;� �;*��;��;H��;?5�;i��;z��;|Z�;{9�;�1�;�E�;�z�;Ґ;�N�;'�;��{;ioo;�c;�GX;0M;fB;`�7;�-;��#;�;=�;�`;���:5I�:B�:���:o��:�/�:/�:���:in}:�eb:�AH:��.:[<:�<�9Y��92T�9�_`9��9�q%8��F�g����g�r��|+ι������)���?��=U�B�j�9���M���������H�����_轺MȺ�Һ�_ݺ��=��~���NW���	��K�0��6)������$��*�J1/��J4�EX9�j^>�nbC�gH��sM�։R�S�W���\�E%b�^wg� �l��<r�ݨw��}��B����������T��i���J����@���ޓ��{������  �  ѧ=�S= �=`�=�R=*�=��=�I=�� =� =J< =���<:�<*d�<��<�	�<�^�<���<��<�e�<Z��< �<�l�<f��<O�<e�<���<J �<'K�<���<x��<�%�<n�<���<���<�I�<���<���<Z)�<�s�<��<��<.J�<���<���<?�<O>�</q�<���<���<(��<��<�1�<�M�<6f�<�{�<ҍ�<,��<>��<��<��<^��<���<z�<�W�<@+�<���<���<+b�<L�<4��<`3�<j��<�5�<3��<G�<aw�</��<(�<v�<���<���<19�<2m�<���</��<7�<���<��</�<#�<�&�<&�<c"�<��<��<��<g�<c��<���<l�<E�<��<�ؑ<�Ϗ<�ō<��<0��<��<|��<�t�<9^�<,�~<�Yz<�&v<��q<>�m<��i<�ee<�;a<]<��X<�T<��P<��L<vyH<]D<d?@<� <<��7<�3<�/<`�+<9p'<MM#<z-<<*�<��<j�<6�
<��<�<�7�;�|�;���;2�;���;��;k��;�4�;��;	��;hL�;�&�;��;1,�;�]�;���;B.�;,҃;�@{;D2o;!zc;�X;�M;*EB;�7;V�-;��#;�;ȣ;[u;��:ӓ�:b��:$�:�*�:4��:��:�@�:�~:�zc:nHI:��/:x:���9��9\9�9��a9C]9I&8��H���Gi�
#��̅Ϲ������A�*��@��OV�F�k� \��8Ɋ����^`������Գ�����jȺ��Һ�Wݺ���>�������/��	�$������C?�Ɉ$���)���.�G4�(9�q,>��6C��DH�tYM�(yR��W�M�\��/b�Z�g�[�l��ar���w��L}�`�����Ɇ�bv��
�������^������
����,���  �  ��=ZR=$�=&�="S= �=S�=�K=�� =S� =@ =��<�<lm�<<��<��<�g�<׽�<��<Jl�<���<�<�o�<��<��<Qd�<���<!��<�F�<I��<���<[�<�e�<��<���<e@�<���<��<�!�<�l�<���<���<hF�<K��<���<?�<u?�<�s�<+��<~��<���<o�<9�<�U�<3o�<���<��<(��<���<��<���<"��<@��<�}�<;Z�<C,�<���< ��<�_�<N�<��< -�<��<�-�</��<�
�<�m�<���<��<1m�<���<p��<3�<%h�<Ж�<���<�߳<���<��<��<�&�<R+�<�+�<p)�<�$�<�<��<��<��<���<���<�<��<7ޑ<aԏ<aɍ<R��<;��<ۛ�<���<)r�<3Z�<��~<�Mz<zv<��q<��m<D�i<�Re<;)a<>]<�X<�T<~�P<ՊL<�pH<�VD<�;@<Q<<� 8<��3<v�/<�+<6{'<�Z#<�<<�"<@<��<��<C�
<�<�<�V�;��;l��;D�;��;'#�;k��;�3�;��;}�;J<�;��;9�;��;>�;��;F�;ٮ�;��z;%�n;>c;�W;��L;. B;�7;��-;��#;Z;��;��;"?�: ��:���:q��:ש�::�:
K�:�֍:��:՞d:XJ:��0:�:r/�9�U�9*�9?�b9k9Sg&8�K�����j��T����й�V��"���+�'�A�WtW���l�Zꀺ0O��Õ���˟��󩺕���K��|�Ⱥ�Һ�Pݺp��|��A����Sq	�!��|B�C�����7>$�ix)�7�.���3���8���=��	C��!H��>M��hR���W���\��<b�^�g��m���r�`x�*�}�����9��9톻:���SB���㎻�����`����A���  �  ��=�P=7�=ɨ=gS=�=Υ=�M=P� =�� =�C =@��<�%�<�v�<r��<��<Fp�<���<�<kr�<���<�<1r�<���<�<Tc�<���<���<:B�<���<#��<��<t]�<��<o��<7�<с�<y��<{�<pe�<۰�<���<~B�<���<��<��<j@�<�u�<���<��<���<) �<A�<L^�<x�<��<��<��<��<y��<���<���<ƛ�<��<8\�<-�<��<t��<�\�< �<���<�&�<���<-%�<:��<2�<�c�<���<�<Jd�<@��<�<�,�<c�<ʒ�<���<^޳<a��<�<��<I*�< 0�<�1�<I0�<R,�<�&�<��<��<��<��<��<���<s�<��<�؏<�̍<U��<��<Z��<\��<9o�<$V�<�w~<�@z<�	v<n�q<�m<�mi<�?e<ra<S�\<>�X<��T<$�P<�L<�gH<5PD<�7@<�<<�8<'�3<M�/<~�+<߅'<�g#<�K<�3<? <�<�<�<�<^#<.u�;(��;l��;�U�;���;"+�;��;h1�;B��;q�;,�;���;��;��;�;�n�;��;�;$�z;i�n;? c;��W;��L;$�A;ږ7;�|-;��#;;�;؛;�w�:;-�:�Z�:z�:-%�:«:�ڜ:�i�:bm�:�e:iK:�1:��:�P :R��9��9id9��9��%8��M�h*�t�l������yҹ� ���.�,���B���X���m��z��bՋ����_9��P��Rg�������Ⱥ��Һ�Oݺ���%[���>��JA	������M]�Э���#��/)��_.���3�h�8���=���B�w�G��%M�zYR��W���\��Jb���g��2m���r�W;x�\�}�����\\��������Lg���������4��OƖ�W���  �  ��=<O=J�=e�=�S=��=�=�O=�� =y� =G =���<�-�<�~�<��<$�<Jx�<��<�"�<x�<0��<�!�<�t�<���<�<Yb�<^��<d��<�=�<��<���<r�<~U�<s��<���<R.�<'y�<6��<��<�^�<��<���<�>�<̈́�<���<c�<&A�<�w�<y��<&��<� �<P&�<�G�<f�<,��<{��<���<#��<���<[��<ͽ�<��<˟�<˃�<^�<�-�<]��<ի�<�Y�<&��<���<r �<���<9�<���<��<�Z�<��<�<�[�<x��<;�<�&�<$^�<�<;��<�ܳ<���<��<�!�<V-�<,4�<7�<�6�<a3�<e.�<�'�<X �<3�<��<��<V��<��<��<�܏<fύ<��<���<ɚ�<���<Rl�<>R�<;m~<�4z<��u<��q<;�m<\i<7.e<�a<2�\<?�X<\�T<}�P<�tL<U_H<�ID<�3@<�<<>8<�3<Y�/<�+<��'<ws#<bY<�B<�0<�#<U<I<|$<�2<ې�;w��;J�;ce�;���;�1�;ө�;/�;9��;ve�;>�;�;.Ѥ;Dם;���;N�;�ŉ;Ci�;`rz;�nn;��b;wW;�|L;�A;�z7;�h-;؛#;�;Q�;��;���:�p�:L��:3g�:j��:s?�:�^�:p�:%��:V�f:AeL:\�2:��:�� :���9�ӡ9�e9�9B%8kgP��x���n������ӹY� �^��|�-�QD�ԶY��o�F��V��w���G�������Ǯ�����,�Ⱥ,Ӻ_QݺL�纞7����λ��	��o������hk��#���(��.�KJ3�Rp8�Ē=��B���G�^M�.LR���W���\�'Xb�Q�g��Rm��r��kx�q�}�Ϳ���}���4��u㉻9���`(��[����P���ޖ�Ml���  �  ��=�M=W�=��=�S=`�=*�=6Q=�� =� =�I =��<�4�<��<.��<&+�<�~�<^��<(�<�|�<��<i$�<tv�<���<�<Ha�<F��<x��<:�<Z�<=��<	�<�N�<7��<)��<�&�<�q�<��<F�<�X�<ĥ�<���<e;�<U��<��<��<�A�<�x�<��<���<�<w+�<�M�<vl�<��<���<���<���<!��<T��<���<3��<0��<2��<h_�< .�<���<)��<�V�<���<��<�<E��<K�<"��<c��<�R�<���<i�<dT�<���< �<�!�<�Y�<���<���<]۳<w��<Y�<F#�<�/�<�7�<�;�<�;�<t9�<�4�<�.�<v'�<H�<q�<%�<<�<���<�<"��<�э<��<���<,��<��<�i�<�N�<\d~<*z<s�u<F�q<�m<Mi<�e<��`<��\<`�X<��T<P�P<JkL<�WH<�CD<�/@<�<<|8<V�3<��/<�+<��'<m}#<e<�O<�><�2<,<�+<d2<�?<\��;���;"�;Qr�;���;*7�;B��;F,�;=��;$[�;�;}׫;��;�;K�;_2�;降;�K�;�9z; 8n;��b;�HW;SUL;n�A;�a7;{V-;�#;�;��;��;)��:���:}��:���:���:���:Ν:Xf�:'j�:j�g:�7M:�p3:�>:u�:_x�9�y�9��e9�V9I�$8$4S�y���<p�pɦ��2չ2���b��.���D���Z�J�o�kw��`Ō����������y뾺,�Ⱥ,Ӻ5Sݺ���k����������JD�;����e3��v#��(�d�-��3��A8��j=�֕B�)�G�:�L��AR��W���\��fb���g�om��s���x��)~��ځ�d����R��������E���ڑ��i�������~���  �  :�=�L=��=��=�S=��=�=^R=C� =�� =L =���<�9�<���<���<�0�<��<��<=,�<Y��<���<�&�<�w�<Z��<��<d`�<���< ��<�6�<�{�<Ͽ�<7�<OI�<i��<7��<� �<�k�<���<G�<T�<̡�<-��<�8�<}��<���<t�<�A�<�y�<���<��<K�<S/�<[R�<Xq�<f��< ��<��<e��<��<���<���<f��<���<��<O`�<F.�<5��<Ȩ�<�T�<���<}��<��<Z��<�<`��<8��<TL�<?��<C��<�N�<l��<K޼<w�<DV�<ш�<ô�<ڳ<���<��<Q$�<�1�<[:�<�>�<�?�<>�<�9�<34�<�,�<�$�<��<�<��<c��<0�<��<vӍ<X<!��<���<���<�g�<�K�<j]~<�!z<��u<�q<mtm<Ai<�e<��`<��\<�X<ύT<�wP<�cL<|QH<w?D<~,@<V<<U8<��3<��/<��+<ݝ'<ӄ#<�m<�Y<jI<�=<�7<E7<=<�I<ֹ�;���;�.�;�{�;;��;d:�;ī�;�)�; ��;�R�;��;�ɫ;G��;���;і;�;��;�4�;cz;�n;�lb;%W;7L;ϚA;OM7;�H-;,�#;�;s�;�;:��:���:�,�:���:I?�:��:�%�:׾�:�:kVh:\�M:
4:�:��:!�94�9,cf9�9��#8!�U�9��&�q����k*ֹ�0�N���/�(�E�j[�v�p��Ԃ�����<���B���3���!������ɺ(Ӻ�Vݺ{��`�~���:�����#��r���T��J#��(�ͽ-�4�2��8�M=��|B���G�J�L��;R���W���\��qb���g�K�m��s�Էx��O~����(j��-�������[���|����������  �  M�=L=$�=c�=�S=��=d�=S=*� =� =sM =���<$=�<͎�<
��<�3�<I��<��<�.�<���<���<�'�<�x�<���<��<�_�<���<���<�4�<Hy�<��<�<�E�<׋�<���< �<Yh�<��<�<7Q�<@��<��<�6�<(�<��<�<B�<�z�<Ϯ�<���<B
�<�1�<-U�<rt�<���<P��<n��<���<��<���<A��<_��<2��<��<�`�<m.�<���<��<�S�<���<A��<9�<S��<��<�}�<t��<�H�<���<���<K�<��<Tۼ<��<T�<��<u��<Yٳ<���<��<�$�<�2�<�;�<�@�<ZB�<�@�<=�<a7�<E0�<(�<��<�<g
�<���<�<�<}ԍ<�<@��<9��<ڀ�<]f�<J�<�X~<vz<��u<M�q<,mm<�9i<Me<X�`<��\<��X<��T< rP<1_L<�MH<i<D<z*@<J<<A8<��3<l�/<��+<�'<��#<Os<�_<�O<�D<g><�=<�C<�O<#��;]��;;6�;؁�;C��;�<�;���;:(�;d��;BM�;z��;���;���;Ƞ�;�Ö;]�;q��;'�;��y;�m;fSb;�W;�#L;��A;T@7;?-;��#;�;��;!�;�:��:�L�:�"�:Jm�:�*�:hY�:��:���:C�h:D<N:_4:�:]7:���9�=�9�f9�9I#8�V��,��br��"����ֹ���xh��/�`F���[��-q�z��}R���n��"o���Z���A��,���$ɺ�1Ӻ�Yݺ���~��6m���y������l[�w������/#��l(��-���2��8� :=�$nB�W�G�t�L�
7R���W��\��xb�h�Ĕm��/s���x��g~�w���g���rx��a(���͌�Dj������Έ��=����  �  �=�K=��=Q�=�S=�=��=]S=� =H� =�M =���<?>�<��<i��<5�<b��<��<�/�<L��<I��<`(�<�x�<���<��<�_�<A��<��<Y4�<ox�<(��< �<�D�<���<=��<��<g�<��<��<?P�<W��<X��<m6�<�~�<���<�<B�<�z�</��<<��<�
�<�2�<V�<�u�<���<���<ȹ�<���<:��<���<���<��<ɧ�<d��<
a�<g.�<���<���<S�<\��<���<D�<S��<w�<h|�<(��<�F�<���<B��<�I�<딾<[ڼ<��<lS�<���<��<$ٳ<���<��<$%�<N3�<<�<�A�<C�<�A�<$>�<�8�<�1�<X)�< �<*�<M�<���<��<��<�ԍ<$Ë<D��<��<���<�e�<�I�<oW~<�z<��u<�q<�jm<57i<4e<��`<]�\<��X<v�T<ApP<�]L<|LH<_;D<�)@<�<<78<��3<��/<��+<آ'<�#<u<�a<AR<(G<:A<t@<F<�Q<���;���;9�;3��;r��;q=�;��;�'�;"��;}K�;X��;���;���;���;r��;�	�;�~�;!�;"�y;/�m;�Jb;tW;�L;M�A;d<7;�;-;(�#;\;��;b�;�
�:Y��:+X�: /�:d|�:�<�:^k�:]
�:|�:f�h:�`N:}4:':UM:X��9�W�9/�f9��9*$#8�WW�
f�_�r�M��[׹���_���0��EF�d\�]q�q ��~e��l����}���h��_K���3���*ɺ
4Ӻ_Zݺp��U��e���t���e��S����a��%#�xb(�;�-�*�2��8�4=��hB���G���L��5R���W��\��zb�h��m��5s��x��o~� ���Ä��}���.��Lӌ��n��6�������� ����  �  M�=L=$�=c�=�S=��=d�=S=*� =� =sM =���<$=�<͎�<
��<�3�<I��<��<�.�<���<���<�'�<�x�<���<��<�_�<���<���<�4�<Hy�<��<�<�E�<׋�<���< �<Yh�<��<�<7Q�<@��<��<�6�<(�<��<�<B�<�z�<Ϯ�<���<B
�<�1�<-U�<rt�<���<P��<n��<���<��<���<A��<_��<2��<��<�`�<m.�<���<��<�S�<���<A��<9�<S��<��<�}�<u��<�H�<���<���<K�<��<Tۼ<��<T�<��<u��<Yٳ<���<��<�$�<�2�<�;�<�@�<ZB�<�@�<=�<a7�<E0�<(�<��<�<g
�<���<�<�<}ԍ<�<@��<9��<ڀ�<]f�<J�<�X~<uz<��u<M�q<,mm<�9i<Me<X�`<��\<��X<��T< rP<1_L<�MH<j<D<{*@<J<<B8<��3<m�/<��+<�'<��#<Os<�_<�O<�D<g><�=<�C<�O<#��;]��;;6�;؁�;B��;�<�;���;9(�;c��;AM�;z��;���;���;Ƞ�;�Ö;]�;p��;'�;��y;�m;fSb;�W;�#L;��A;T@7;?-;��#;�;��;!�;�:��:�L�:�"�:Jm�:�*�:hY�:��:���:C�h:D<N:_4:�:]7:���9�=�9�f9�9I#8�V��,��br��"����ֹ���xh��/�`F���[��-q�z��}R���n��"o���Z���A��,���$ɺ�1Ӻ�Yݺ���~��6m���y������l[�w������/#��l(��-���2��8� :=�$nB�W�G�t�L�
7R���W��\��xb�h�Ĕm��/s���x��g~�w���g���rx��a(���͌�Dj������Έ��=����  �  :�=�L=��=��=�S=��=�=^R=C� =�� =L =���<�9�<���<���<�0�<��<��<=,�<Y��<���<�&�<�w�<Z��<��<d`�<���< ��<�6�<�{�<Ͽ�<7�<OI�<i��<7��<� �<�k�<���<G�<T�<̡�<-��<�8�<}��<���<t�<�A�<�y�<���<��<K�<S/�<[R�<Xq�<f��< ��<��<e��<��<���<���<f��<���<��<O`�<F.�<5��<Ȩ�<�T�<���<}��<��<Z��<�<`��<8��<TL�<?��<C��<�N�<m��<K޼<w�<DV�<ш�<ô�<ڳ<���<��<Q$�<�1�<[:�<�>�<�?�<>�<�9�<34�<�,�<�$�<��<�<��<c��<0�<��<vӍ<X< ��<���<���<�g�<�K�<j]~<�!z<��u<�q<mtm<Ai<�e<��`<��\<�X<ύT<�wP<�cL<|QH<x?D<~,@<V<<U8<��3<��/<��+<ݝ'<ӄ#<�m<�Y<jI<�=<�7<E7<=<�I<ֹ�;���;�.�;�{�;:��;c:�;ë�;�)�;���;�R�;��;�ɫ;F��;���;і;�;��;�4�;az;�n;�lb;%W; 7L;ϚA;NM7;�H-;,�#;�;s�;�;:��:���:�,�:���:I?�:��:�%�:׾�:�:kVh:\�M:
4:�:��:!�94�9,cf9�9��#8!�U�9��&�q����k*ֹ�0�N���/�(�E�j[�v�p��Ԃ�����<���B���3���!������ɺ(Ӻ�Vݺ{��`�~���:�����#��r���T��J#��(�ͽ-�4�2��8�M=��|B���G�J�L��;R���W���\��qb���g�K�m��s�Էx��O~����(j��-�������[���|����������  �  ��=�M=W�=��=�S=`�=*�=6Q=�� =� =�I =��<�4�<��<.��<&+�<�~�<^��<(�<�|�<��<i$�<tv�<���<�<Ha�<F��<x��<:�<Z�<=��<	�<�N�<7��<)��<�&�<�q�<��<F�<�X�<ĥ�<���<e;�<U��<��<��<�A�<�x�<��<���<�<w+�<�M�<vl�<��<���<���<���<!��<T��<���<3��<0��<2��<h_�< .�<���<)��<�V�<���<��<�<E��<K�<"��<d��<�R�<���<i�<dT�<���< �<�!�<�Y�<���<���<]۳<w��<Z�<G#�<�/�<�7�<�;�<�;�<t9�<�4�<�.�<v'�<H�<p�<%�<;�<���<�<"��<�э<~��<���<,��<��<�i�<�N�<[d~<*z<r�u<E�q<�m<Mi<�e<��`<��\<`�X<��T<Q�P<KkL<�WH<�CD<�/@<�<<}8<V�3<��/<�+<��'<m}#<e<�O<�><�2<,<�+<d2<�?<[��;���;"�;Pr�;���;)7�;A��;D,�;<��;#[�;�;|׫;��;�;J�;^2�;;�K�;�9z;8n;��b;�HW;SUL;m�A;�a7;zV-;�#;�;��;��;)��:���:}��:���:���:���:Ν:Xf�:'j�:j�g:�7M:�p3:�>:u�:_x�9�y�9��e9�V9I�$8$4S�y���<p�pɦ��2չ2���b��.���D���Z�J�o�kw��`Ō����������y뾺,�Ⱥ,Ӻ5Sݺ���k����������JD�;����e3��v#��(�d�-��3��A8��j=�֕B�)�G�:�L��AR��W���\��fb���g�om��s���x��)~��ځ�d����R��������E���ڑ��i�������~���  �  ��=<O=J�=e�=�S=��=�=�O=�� =y� =G =���<�-�<�~�<��<$�<Jx�<��<�"�<x�<0��<�!�<�t�<���<�<Yb�<^��<d��<�=�<��<���<r�<~U�<s��<���<R.�<'y�<6��<��<�^�<��<���<�>�<̈́�<���<c�<&A�<�w�<y��<&��<� �<P&�<�G�<f�<,��<{��<���<#��<���<[��<ͽ�<��<˟�<˃�<^�<�-�<]��<ի�<�Y�<&��<���<r �<���<9�<���<��<�Z�<��<�<�[�<x��<<�<�&�<$^�<�<;��<�ܳ<���<��<�!�<V-�<-4�<7�<�6�<a3�<e.�<�'�<X �<3�<��<��<U��<��<��<�܏<fύ<��<���<ɚ�<���<Ql�<>R�<;m~<�4z<��u<��q<;�m<\i<7.e<�a<2�\<?�X<\�T<~�P<�tL<U_H<�ID<�3@<�<<?8<�3<Z�/<�+<��'<ws#<cY<�B<�0<�#<U<I<{$<�2<ڐ�;u��;I�;ae�;���;�1�;ѩ�;/�;7��;te�;=�;�;-Ѥ;Bם;���;N�;�ŉ;Ai�;^rz;�nn;��b;wW;�|L;�A;�z7;�h-;כ#;�;Q�;��;���:�p�:L��:3g�:j��:s?�:�^�:p�:%��:V�f:@eL:\�2:��:�� :���9�ӡ9�e9�9B%8kgP��x���n������ӹY� �^��|�-�QD�ԶY��o�F��V��w���G�������Ǯ�����,�Ⱥ,Ӻ_QݺL�纞7����λ��	��o������hk��#���(��.�KJ3�Rp8�Ē=��B���G�^M�.LR���W���\�'Xb�Q�g��Rm��r��kx�q�}�Ϳ���}���4��u㉻9���`(��[����P���ޖ�Ml���  �  ��=�P=7�=ɨ=gS=�=Υ=�M=P� =�� =�C =@��<�%�<�v�<r��<��<Fp�<���<�<kr�<���<�<1r�<���<�<Tc�<���<���<:B�<���<#��<��<t]�<��<o��<7�<с�<y��<{�<pe�<۰�<���<~B�<���<��<��<j@�<�u�<���<��<���<) �<A�<L^�<x�<��<��<��<��<y��<���<���<ƛ�<��<8\�<-�<��<t��<�\�< �<���<�&�<���<-%�<:��<2�<�c�<���<�<Jd�<@��<�<�,�<c�<ʒ�<���<^޳<a��<�<��<I*�<0�<�1�<I0�<S,�<�&�<��<��<��<��<��<���<r�<��<�؏<�̍<T��<��<Z��<[��<9o�<$V�<�w~<�@z<�	v<n�q<�m<�mi<�?e<ra<S�\<?�X<��T<%�P<�L<�gH<6PD<�7@<�<<�8<(�3<N�/<�+<��'<�g#<�K<�3<? <�<�<�<�<^#<-u�;&��;k��;�U�;���; +�;��;f1�;@��;q�;,�;���;��;��;�;�n�;��;�;"�z;g�n;= c;��W;��L;#�A;ٖ7;�|-;��#;;�;؛;�w�:;-�:�Z�:y�:-%�:«:�ڜ:�i�:bm�:�e:iK:�1:��:�P :R��9��9id9��9��%8��M�h*�t�l������yҹ� ���.�,���B���X���m��z��bՋ����_9��P��Rg�������Ⱥ��Һ�Oݺ���%[���>��JA	������M]�Э���#��/)��_.���3�h�8���=���B�w�G��%M�zYR��W���\��Jb���g��2m���r�W;x�\�}�����\\��������Lg���������4��OƖ�W���  �  ��=ZR=$�=&�="S= �=S�=�K=�� =S� =@ =��<�<lm�<<��<��<�g�<׽�<��<Jl�<���<�<�o�<��<��<Qd�<���<!��<�F�<I��<���<[�<�e�<��<���<e@�<���<��<�!�<�l�<���<���<hF�<K��<���<?�<u?�<�s�<+��<~��<���<o�<9�<�U�<3o�<���<��<)��<���<��<���<"��<@��<�}�<;Z�<C,�<���< ��<�_�<N�<��<!-�<��<�-�<0��<�
�<�m�<���<��<2m�<���<q��<3�<%h�<і�<���<�߳<���<��<��<�&�<R+�<�+�<p)�<�$�<�<��<��<��<���<���<�<��<6ޑ<aԏ<`ɍ<R��<:��<ۛ�<���<)r�<3Z�<��~<�Mz<yv<��q<��m<D�i<�Re<;)a<>]<�X<�T<�P<֊L<�pH<�VD<�;@<R<<� 8<��3<w�/<��+<7{'<�Z#<�<<�"<A<��<��<B�
<�<�<�V�;��;j��;D�;��;%#�;i��;�3�;��;}�;H<�;��;7�;��;>�;	��;E�;خ�;��z;#�n;>c;�W;��L;- B;�7;��-;��#;Y;��;��;"?�: ��:���:q��:֩�::�:
K�:�֍:��:՞d:XJ:��0:�:r/�9�U�9*�9?�b9k9Sg&8�K�����j��T����й�V��"���+�'�A�WtW���l�Zꀺ0O��Õ���˟��󩺕���K��|�Ⱥ�Һ�Pݺp��|��A����Sq	�!��|B�C�����7>$�ix)�7�.���3���8���=��	C��!H��>M��hR���W���\��<b�^�g��m���r�`x�*�}�����9��9톻:���SB���㎻�����`����A���  �  ѧ=�S= �=`�=�R=*�=��=�I=�� =� =J< =���<:�<*d�<��<�	�<�^�<���<��<�e�<Z��< �<�l�<f��<O�<e�<���<J �<'K�<���<x��<�%�<n�<���<���<�I�<���<���<Z)�<�s�<��<��<.J�<���<���<?�<O>�</q�<���<���<(��<��<�1�<�M�<6f�<�{�<ҍ�<,��<>��<��<��<^��<���<z�<�W�<@+�<���<���<+b�<L�<4��<`3�<j��<�5�<3��<H�<aw�</��<(�<v�<���<���<29�<2m�<���<0��<8�<���<��<0�<#�<�&�<&�<c"�<��<��<��<g�<c��<���<l�<E�<��<�ؑ<�Ϗ<�ō<��<0��<��<|��<�t�<8^�<,�~<�Yz<�&v<��q<>�m<��i<�ee<�;a<]<��X<�T<��P<��L<vyH<]D<e?@<� <<��7<�3<�/<a�+<9p'<NM#<{-<<*�<��<j�<6�
<��<�<�7�;�|�;���;2�;���;��;i��;�4�;��;��;fL�;�&�;��;/,�;�]�;���;A.�;+҃;�@{;B2o;zc;�X;�M;)EB;�7;U�-;��#;�;ǣ;[u;��:ғ�:a��:$�:�*�:3��:��:�@�:�~:�zc:nHI:��/:x:���9��9\9�9��a9C]9I&8��H���Gi�
#��̅Ϲ������A�*��@��OV�F�k� \��8Ɋ����^`������Գ�����jȺ��Һ�Wݺ���>�������/��	�$������C?�Ɉ$���)���.�G4�(9�q,>��6C��DH�tYM�(yR��W�M�\��/b�Z�g�[�l��ar���w��L}�`�����Ɇ�bv��
�������^������
����,���  �  ��=U=��=}�=SR=3�=$�=vG=A� =�� =�8 =���<��<n[�<-��<� �<�V�<���<��<�_�<@��<�<�i�<ſ�<��<�e�<Y��<�<O�<Ù�<���<�,�<�u�<ݾ�<U�<&R�<?��<���<�0�<z�<w��<	�<vM�<��< ��<�</=�<�n�< ��<T��<y��<.�<`*�<�E�<�]�<s�<(��<���</��<ǣ�<���<���<#��<�v�<�U�<B*�<���<��<�d�<��<٧�<19�<+��<R=�<���<��<j��<3��<�0�<G~�<ž<D�<�>�<�q�<靷<võ<I�<���<��<��<��<�!�<D �<��<9�<k�<��<���<���<?�<r�<��<�ٓ<�ґ<vˏ<�<뷋<&��<��<���<"w�<�a�<]�~<dez< 4v<�r<u�m<��i<�ve<�La<�%]<� Y<��T<��P<��L<�H<QbD<�B@<6!<<+�7<Z�3<�/<�+<me'<�@#<+<<��<�<f�<5�
<V�<z�<�;Bc�;κ�;� �;(��;��;F��;=5�;g��;x��;zZ�;y9�;�1�;�E�;�z�;Ґ;�N�;&�;��{;hoo;�c;�GX;0M;fB;_�7;�-;��#;�;=�;�`;���:5I�:B�:���:o��:�/�:/�:���:in}:�eb:�AH:��.:[<:�<�9Y��92T�9�_`9��9�q%8��F�g����g�r��|+ι������)���?��=U�B�j�9���M���������H�����_轺MȺ�Һ�_ݺ��=��~���NW���	��K�0��6)������$��*�J1/��J4�EX9�j^>�nbC�gH��sM�։R�S�W���\�E%b�^wg� �l��<r�ݨw��}��B����������T��i���J����@���ޓ��{������  �  '�=V=M =��=�Q=9�=��=�E=�� =8� =�5 =#��<��<�S�<���<q��<wO�<J��<� �<�Z�<Դ�<��<g�<
��<�<�e�<���<^�<PR�<���<���<�2�<'|�<���<o�<OY�<<��<+��<�6�<}�<��<��<4P�<���<���<��<�;�<�l�<��<O��<���<t�<�#�<�>�<}V�<�k�<�}�<q��<@��<]��<���<���<'��<�s�<�S�<)�<���<ز�<�f�<��<ȫ�<>�<���<�C�<~��<T$�<���<���<�7�<,��<`˾<�
�<�C�<mu�<���<Cŵ<�<X��<\�<u�<q�<��<B�<��<��<h�<���<��<+�<�<�ߗ<�ٕ<ԓ<(Α<�Ǐ<���<ĵ�<��<���<���<y�<�d�<�~<�nz<\?v<hr<��m<��i<k�e<#[a<B3]<�Y<i�T<��P<ۧL<s�H<�fD<$E@<�!<<��7<��3<_�/<��+<+\'<�5#<c<�<6�<��<��<��
<��<y�<N�;�L�;���;\�;O��;9
�;P��;F5�;^��;d��;$f�;�H�;�D�;;\�;<��;'�;$j�;��;X�{;'�o;|�c;IqX;�RM;�B;��7;|�-;A�#;�	;�;�M;���:��:B��:=^�:�J�:���:���:�9�:Nz|:�za:`G:<.:N�:��9��9%��9�4_9-9d�$8��E����8f��+��5͹h���+�)��>��XT�}�i���~�)扺RO��뫞�e��&^�������5Ⱥ��ҺhݺN)�g����z�.�	�|�N��b�����%��D*�k/���4�"�9��>��C���H���M�A�R�g�W�(�\�(b�\gg���l�Kr���w��|��)���ۃ�a���n7��#���]����'��ȓ�+h���	���  �  I�=�V=� =��=�Q=|�=��=D=)� =� ==3 =���<���<N�<���<���<�I�<=��<���<�V�<]��<��<e�<���<v�<f�<���<�<�T�<��<R��<�6�<��<
��<��<�^�<���<7��<T;�<���<w��<��<3R�<��<9��<��<�:�<�j�<���<��<���<��<�<G9�<�P�<�e�<�w�<���<��<���<x��<&��<���<Eq�<�Q�<'(�<w��<h��<�g�<��<���<�A�<��<�H�<Ƚ�<*�<ʍ�<���<�=�<a��<!о<��<G�<;x�<���<qƵ<��<��<N
�<��<��<r�<c�<k�<�	�<� �<���<"�<=�<8��<Dڗ<�ԕ<�ϓ<pʑ<_ď</��<&��<!��<Л�<-��<kz�<�f�<�~<vz<�Gv<�r<e�m<�i<��e<\fa<�=]<�Y<�T<"�P<�L<8�H<jD<�F@<�!<<3�7<��3<�/<�~+<�T'<	-#<�<��<{�<��<=�<��
<��<��<w��;N;�;Θ�;��;L~�;��;֕�;�4�;���;���;�n�;�T�;�R�;�l�;���;� �;I�;�#�;��{;��o; d;�X;�lM;ԖB;O8;��-;��#;�;��;�?;l�:���:մ�::�:v��:h�:�[�:jً:�{:��`:��F:�u-:��:��9J�9���9�S^9�z9�($8��D�S��De�񀟹�6̹y����r�ia(��>���S��i�k*~�����U��tn��Ш�6��å��q'Ⱥ��ҺDpݺ�=躎#�5 ��E��T
����j��������;%�/t*�S�/���4���9��>�"�C�z�H�ٜM���R� �W��\��b�2\g�^�l��r�=fw���|����!ǃ�[u��[!��ʋ�mp�����9����Y�������  �  ��=KW=� =��=BQ=��=�=(C= � =�� =�1 =���<I��<~J�<���<���<>F�<��<���<�S�<&��<�	�<�c�<Ի�<�<)f�<��<
�<;V�<���<���<�9�<��<B��<A�<*b�<��<b��<@>�<!��<���<0�<rS�<���<���<w�<K:�<�i�<���<��<j��<%��<��<�5�<)M�<b�<-t�<��<i��<^��<���<���< ��<�o�<�P�<�'�<T��<ӳ�<�h�<>�<w��<�C�<���<�K�<��<�-�<T��<��<A�<���<&Ӿ<��<&I�<�y�<���<Gǵ<��<���<�	�<��<>�<e�<��<��<��<f��<T��<��<��<�ܙ<�֗<�ѕ<�̓<ȑ<j<���<��<���<���<���<>{�<h�<^�~<�zz<Mv<�r<��m<x�i<c�e<ma<xD]<�Y<��T<��P<αL<$�H<�kD<�G@<�!<<J�7<��3<�/<�z+<CP'<�'#<�<��<#�<;�<�<S�
<]�<��<���;:0�;G��;��;x�;���;���;_4�;\��;`��;!t�;r[�;�[�;Ow�;{��;��;���;�0�;Y�{;G�o;gd;��X;�|M;�B;s8;x�-;��#;�;";�5;nQ�:v��:���:���:Hȸ:`/�:8"�:E��:�F{:�K`: @F:�-:�:nd�9?��9w�9��]9�!9��#8�?D�+�
�M�d�x����˹���{���'�X�=��=S��h���}�f��#ۓ�uG��򰨺���l����Ⱥ��Һ�uݺ�J�(9�0<������0
�����7�(��A �aX%���*��/�'�4�F�9���>��C�­H�+�M��R�q�W���\�b�`Ug���l��q�PTw�f�|��
��Z���\h���������c��^��Y����P��r����  �  v�=*^=�=��=
X=:�=C�=rG=� =�� =c2 =0��<���<�H�<?��<c��<�J�<0��<��<�e�<^��<x&�<��<���<�;�<u��<p��<�:�<}��<l��<.(�<=u�<��<��<�[�<���<a��<5B�<���<[��<�$�<~m�<���<���<�5�<�p�<d��<���<��<V.�<�R�<�s�<Q��<���<���<���<���<��<��<�-�<7�<�9�<�4�<f&�<��<���<���<2}�<4�<���<�|�<I�<���<H�<���<*��<�O�<H��<���<?�<��<���<<�<��<j<�<�Y�<p�<H�<���<���<υ�<}�<~p�<fa�<�P�<@�<�/�<!�<c�<�	�<=�<7��<X��<��<��<���<l׋<eˉ<���<��<���<-��<N�~<��z<�ev<�/r<��m<P�i<v�e<>^a<�-]<��X<��T<�P<%L<PUH<X*D<��?<^�;<@�7<�f3<�./<D�*<�&<��"<�M<�<Y�<V�<��<f�	<U�<��<d��;��;�v�;?��;O�;F��;
S�;���;{��;�.�;]�;��;��;N��;ؔ;;"�;ő�;�(�;4�u;Τi;s�];�OR;�$G;K<;I�1;[|';�~;�;RB
;�� ;���:KQ�:5�:1��:���:�"�:�F�:��:ֳd:q�J:Fa1:�):��:9��9�B�9��z9}6#9���8	x+���ø�9�EI���	��z�߹���@��0�*F�-[� "p��w��"Ɍ�v���G������õ�����~ʺ 	պ[�ߺΊ�ӄ��M �����}���V����{!�C�&���+���0���5�J�:�h�?�kyD�FHI�� N��S��W�3]�,b��_g���l�L�q��Iw���|�� ��ŭ��hX��S ������pH���萻����a&��ǘ��  �  (�=^=�=��=-X=p�=��=�G=�� =/� =3 =���<���<�J�<��<%��<mL�<���<9�<'g�<g��</'�<���<%��<(<�<���<O��<�:�<׊�<���</'�<t�<���<H�<�Y�<Ħ�<���<�@�<a��<B��<�#�<�l�<.��<r��<�5�<q�<���<y��<��<//�<�S�<Iu�<ѓ�<"��<���<��<���<U�<C!�<X/�<P8�<�:�<z5�<	'�</�<	��<ȹ�<"}�<�3�<���<�{�<H�<h��<��<u��<���<�M�<��<f��<�=�<�~�<o��<E�<�<�;�<�Y�<p�<o�<���<��<r��<�}�<�q�<�b�<_R�<�A�<�1�<�"�<7�<v�<��<���<���<��<S�<��<�׋<�ˉ<���<���<v��<��<��~<��z<�cv<-r<��m<�i<�e<�Za<�*]< �X<T�T<�P<w}L<TH<�)D<��?<��;<��7<�g3<"0/<��*<I�&<M�"<�P<�!<��<�<��<�	<��<��<A��;$�;{�;k��;�Q�;��;IT�;@��;D��;w-�;�;廩;]��;��;MӔ;��;N��;�!�;v�u;��i;��];[GR;�G;hE<;��1;�z';;�;,E
;S;���:S_�:�H�:���:��:9<�:ga�:�!�:��d: �J:9�1:�Z:?�:3�9�|�9�z9p�#9��8V�)��øL99�Tg��l7����߹˿��h���0��=F��d[�cXp�����ߌ� ��dX������ε�[����ʺպ˳ߺ?��Q{���G ����Zs���ے�*��m!�]�&�I�+���0�1�5���:��?�2pD�BI�zN� S���W��
]��,b��ag�A�l���q�bQw���|��������^��e��+���ON���퐻���;*��=ʘ��  �  J�=r]=�=��=�X='�=��=I=#� =�� =*5 =K��<x �<�O�<��<��<1Q�<5��<8�<�j�<h��<�)�<���<n��<�<�<���<���<O9�<���<��<$�<zp�<���<��<|U�<H��<w��<�<�<���<���<#!�<�j�<���<|��<�5�<q�<���<$��<��<�1�<JW�<y�<��<ô�<w��<i��<r��<-�<�%�<�3�<<�<*>�<38�<3)�<��<���<��<�|�<�2�<O��<�y�<X�<ܑ�<��<��<���<�H�<ɠ�<���<A9�<�z�<���<q�<��<W:�<�X�<�o�<��<���<ǋ�<���<ŀ�<u�<�f�<�V�<LF�<{6�<�'�<'�<U�<m�<���<_��<�<�<��<|ً<�̉< ��<���<k��<�}�<B�~<ȓz<�\v<0%r<�m<*�i<ǃe<�Qa<9"]<�X<�T<ʠP<�xL<[PH<:'D<C�?<��;<8�7<�j3<=4/<��*<��&<��"<Y<7+<�<,�<�<0�	<��<:�<��;3�; ��;��;�Z�;��;�W�;"��;O��;&)�;~�;���;���;I��;�Ô;&�;9z�;��;��u;0yi;>�];�-R;�G;�5<;O�1;4t';"};
�;�M
;o;��:��:�:�:t��:]��: ��:Aq�:�e:CYK:�*2:��:�c:��92�9|9aa$9���8A�%���øɪ9��ň�,���0��*�R���p1���F���[���p��ӂ�� ���Z��񋡺Ӹ��~쵺�0���ʺ�	պ�ߺ�q�3]���4 �/��VW�)��{o�>���F!���&���+���0�w�5�=�:���?�~VD�-I�q
N��R���W��]��0b��jg���l��
r��hw�d�|�����ă�jp��W��꽋�__������=���I6���Ә��  �  ް=�\=B=Ͱ=!Y=, =�=!K=�� =ߓ =o8 =a��<�<�W�<5��<���<�X�<-��<��<<p�<��<v-�<M��<B��<�=�<w��<���<B7�<��<���<�<�j�<6��<��< N�<��<$��<�5�<w��<���<��<
g�<��<��<#5�<�q�<��<f��<�<E6�<]\�<�<ƞ�<��<;��<`��<m�<��<,-�<M:�<B�<:C�<�<�<{,�<��<E��<h��<|�<1�<���<�u�<��<C��<��<y�<G��<5A�<��<8��<Y2�<`t�<���<��<V�<�7�<%W�<@o�<H��<m��<��<&��<*��<Yz�<�l�<~]�<�M�<N>�<�/�< #�<�<��<��<O��<��<F��<��<�ۋ<�͉<R��<�<Ɠ�<L{�<��~<`�z<�Qv<�r<1�m<F�i<�te<�Ba<]<&�X<��T<ݖP<zpL<^JH<E#D<j�?<��;<B�7<}n3<:/<�+<Z�&<C�"<Wf<�9<7<z�<��<��	<D�<��<��;�J�;#��;���;�f�;���;�\�;2��;�}�;L"�;~ذ;���;���;W��;`��;���;�]�;>�;<ju;�Ei;|y];�R;I�F;�<;ڝ1;j';�z;��;�Z
;�#;�Q�:%��:@��:hU�:Qa�:8��:.�:h�:�f:�UL:�3:�:�):�Z�9:P�9�}99�%9���8*m!��7ĸ�T:��_��ŗ��0�ṟ��ܡ��D2��G��\�M�q��F�����������ܡ���� ���S����ʺ�պ��ߺ3V��3��� �G���+����:8�/��_!��L&��x+��0�H�5�at:��S?�/D��I� �M��R�(�W�%]��5b�Zxg�f�l� )r���w���|��.��
���܍���6��Uۋ�{���������~I��+㘻�  �  �=5[=�=̰=�Y=z=��=�M=�� =�� =�< =���<��<�a�<|��<
�<b�<;��<��<Nw�<
��<62�<֍�<���<�>�<'��<���<Z4�<���<���<~�<�b�<���<���<�D�<O��<���<�,�<A{�<r��<��<Tb�<���<���<?4�<Tr�<ݫ�<g��<A�<�;�<�b�<���<j��<n��<��<���<��<�%�<�6�<�B�<�I�<�I�<�A�<�0�<��<���<���<�z�<�.�<���<�p�<X �<Ԅ�<���<�o�<u��<7�<��<z��<&)�<�k�<G��<�ݻ<��<D4�<�T�<^n�<���<A��<'��<r��<���<	��<�t�<Hf�<AW�<@H�<1:�<R-�<�!�<��<&�<��<���<���<
�<�ދ<�ω<���<ݨ�<V��<�w�<ҷ~<~z<�Bv<�r<�m<"�i<Xae<�/a<�]<��X<�T<ЉP<�eL</BH<�D<n�?<~�;<��7<�s3<�A/<+<��&<�"<Zw<wL<Y(<S<��<[�	<~�<��<Q+�;�h�;���;��;�v�; ��;�b�;���;�x�;o�;�ɰ;���;Ko�;�k�;���;�͍;9�;)π;&"u;�i;l:];��Q;2�F;D�;;�1;=Z';�u;��;.j
;N=;���:9-�:{=�:�ҽ:��:���:`Ώ:ʗ�:��g:H�M:J4:��:%:a�9���9��9u''9�q�8���b�ĸ�_;��4��\���G*�Q��'���]3���H�0^�ws��ك�.���6���G���T���d��w����ʺ�պ/�ߺ�2�,��������p�t�
�(v�����\�� �|�%�>'+��<0��>5�j0:�2?���C�y�H���M�%�R�x�W�]�X?b���g�s�l��Pr��w��1}�3P���������>]��W��@����8���Γ��b�������  �  ��=�Y=�=��=[Z=�=�=nP=9� =�� =]A ='��<I�<�m�<_��<��<�m�<���< #�<]�<���<t7�<ő�<���<�?�<���<���<�0�<�|�<��<��<�Y�<g��<���<<9�<݅�<���<g"�<�q�<���<w�<�\�<]��<��<3�<�r�<l��<���<��<�A�<|j�<`��<:��<8��<���<\�<d�<N1�<eA�<�L�<eR�<EQ�<�G�< 5�<��<M��<���<�y�<�+�<V��<�j�<���<�{�<���<�d�<���<+�<��<���<2�<%b�<���<xֻ<��<�/�<R�<1m�<��<⍰<��<%��<���<���<p}�<Kp�<0b�<�S�<F�<(9�<b-�<�"�<��<j�<��<t��<��<��<�Љ<���<j��<j��<s�<�~< oz<e1v<�q<m�m<�i<Je<�a<��\<{�X<��T<�yP<�XL<-8H<�D<��?<��;<��7<�x3<�I/<&+<+�&<�"<��<�a<~?<�$<Y<�	
<�
<D<*R�;���;
��;�'�;���;U��;gh�;���;�r�;L�;<��;mw�;QQ�;{I�;�c�; ��;��;��;��t;�h;�\;��Q;<�F;��;;�d1;�F';-n;`�;�x
;�X;~��:��:���:e_�:���:3E�:I��:�V�:�Zi:PO:��5:P:@:T��9�E�9C,�9w�(9�0�8b ���Ÿ��<��8��������������,�4��=J�r�_��pt����e����ɘ��ɢ�;�������ؿ����ʺ:պ�ߺ�����l����;�δ
�j-�����XY �i�%�v�*���/���4���9���>��C���H�f�M���R�/�W�]��Kb���g�Fm��r�-�w�Fw}�dw���.��k������<.��tʎ��`��	�l���~���  �  ͩ=�W=�=i�=�Z==4�=HS=�� =� =nF =E��<#)�<z�<���<*"�<[y�<���<�,�<Ň�<���<�<�<���<��<S@�<���<W��<�,�<�v�<Ϳ�<��<�O�<S��<���<�,�<vy�<���<��<?g�<���<��<,V�<o��<���<D1�<�r�<���<���<��<�G�<3r�<���<���<���<���<��<�)�<`=�<�L�<>W�<�[�<�X�<	N�<�9�<��<���<���<�w�<.(�<��<d�<y��<&r�<��<�X�<��<��<�u�<?��<V�<iW�<��<sλ< �<+�<�N�<pk�<��<z��<���<�<f��<���<݆�<�z�<�m�<`�<�R�<�E�<Z9�<�-�<9#�<q�<��<��<'�<�<f҉<v��<y��<���<�m�<t�~<�^z<1v<��q<Ѡm<�fi<�0e<��`<��\<S�X<�T<�hP<�JL<�,H<�D<��?<>�;<��7<�}3<2R/<�$+<��&<��"<4�<�x<�W<(><@,<>#
<#<2,<�{�;Ү�;'��;�?�;~��;���;�m�;9��;�j�;���;��;�\�;o0�;�#�;,9�;7v�;5ކ;As�;Wot;QWh;��\;2FQ;�EF;��;;�?1;�/';�b;Q�;C�
;ss;I4�:���:V8�:E��:18�:���:�K�:� �:��j:��P:�7:�p:Xm:n��9+�9�e�9P�*9X��8\��_�Ǹ�(>�Bg������\�湒�	�/ �
6��K��a�?�u��H��Xk���j���W��,6��~�� ��?˺}1պ�{ߺL�����$?�����r
�����G�������6%��d*�M�/���4�d�9���>���C���H�c�M���R�(�W�\	]��\b��g��7m�%�r�->x���}�C����]��*��˼��_����������������",���  �  ��=�U=[=�=?[=>=�=V=\� =N� =NK =+��<�4�<G��<[��<U.�<��<,��<Y6�<���<z��<B�<��<��<�@�<S��<}��<5(�<�p�<E��<���<�E�<��<���<s �<�l�<H��<N�<i\�<��<e��<tO�<N��<B��<D/�<%r�<E��<v��<�<�M�<�y�<z��<���<���<��<�<6�<LI�<�W�<Va�<~d�<``�<	T�<>�<��<���<��<Ou�<Q$�<���<�\�<���<h�<���<tL�<5��<��<�h�<��<U�<FL�<7��< ƻ<Q��<�%�<9K�<di�<���<Ӑ�<���<���<���<P��<���<F��<y�<l�<�^�<�Q�<FE�<9�<3-�<9!�<��<i�<\��<$�<vӉ<̼�<H��<"��<|h�<v�~<�Mz<P
v<^�q<"�m<�Mi<me<��`<��\<��X<ltT<�VP<�;L<� H<D<8�?<��;<��7<��3<�Y/<�/+<�'<��"<�<ێ<�o<HW<�E<o<
<F;<�B<Σ�;���;.�;�V�;���;��;%q�;.��;�a�;V�;[��;�@�;��;d��; �;.H�;%��;�B�;wt;�g;IM\;j�P;�F;�h;;�1;�';�T;
�;��
;��;h~�:\�:D��:��:Eܯ:v��:R�:u�:�|l:R:��8:��:��:t��9�t�9䏃9,9t�8Ҫ�AXɸ+�?�X���cR��@���@t!���7�SGM���b�f�w��	��� ��d��꣺����z��SO���;˺qIպ�yߺ��麩Q������3���2
�������J������$�~*�-#/��74�bB9�hH>�rMC��WH�lM���R���W��]�"ob���g�>cm�{�r��x�.~�E΁������B��ϐ���(��F���A���Ŗ��H���  �  >�=�S==^�=_[='=ï=}X= =-� =�O =-��<�?�<���<���<}9�<���<���<?�<a��<h��<�F�<��<���<�@�<���<���<�#�<
k�<��<Q��<�;�<^��<z��<��<a�<���<@ �<@R�<��<}��<�H�<N��<���<C-�<sq�<��<���<�!�<>S�<c��<���<���<��<p�<T*�<gA�<2T�<>b�<�j�<�l�<%g�<=Y�<�A�<��<n��<���<s�<c �<T��<,V�<���<�^�<��<�@�<���<>�<;\�<_��<���<�A�<���<���<��<� �<�G�<ag�<��<���<�<���<��<Q��<F��<���<���<w�<Fj�<)]�<.P�<CC�<Q6�<>)�<m�<��<���<M�<ԉ<���<��<8��<<c�<ǂ~<X=z<��u<�q<�rm<6i<X�d<��`<��\<?�X<aT<�EP<-L<�H<N�C<��?<Z�;<ڧ7<m�3<2`/<V9+<�'<m�"< �<H�<�<dn<z]<�S
<�Q<�V<k��;���;(�;�j�;���;�;s�;���;X�;}޷;w�;%�;��;�ך;"�;?�;z��;��;/�s;˨g;�[;"�P;J�E;@7;;�0;��&;)G;��;{�
;��;��:���:�!�:��:r�:-Z�:E��:���:��m:AyS:W�9:�� :��:ޠ�9�Ҳ9,��9�A-9�e�8����&˸ڙA��ڎ�*缹���A,���"��8���N��d�y�����u͐�/����s���)���ڷ�/���|m˺gaպr}ߺ-���$��e���(����	��P�Ħ�����<��w$��)�%�.���3�8�8�8	>��C��/H�mPM��R���W��]��b�� h�׍m��&s��x�o]~�����p����q���������U��:⑻�f���斻,e���  �  ġ=�Q=� =��=j[=�=�=wZ==\� =�S =���<�H�<��<s��<�B�<���<>��<PF�<���<S��<;J�<|��<���<Z@�<n��<���<��<�e�<���<���<X3�<y�<���<^
�<�V�<���<���<XI�<���<���</C�<���<7��<+�<�p�<���<���<�$�<�W�<���<S��<���<���<��<�3�<�J�<^]�<�j�<xr�<Zs�<�l�<�]�<�D�<�!�<���<	��<�p�<��<���<!P�<g��<QV�<���<�6�<u��<p��<oQ�<��<���<�8�<�z�<���<��<�<(D�<>e�<#�<?��<瞮<å�<��<��<;��<Ŗ�<G��<e��<�s�<�f�<VY�<�K�<>�<�/�<� �<��<���<��<fԉ<��<���<��<{^�<�v~</z<1�u<1�q<�^m<�!i<��d<�`<��\<|mX<PT<�6P<_ L<6H<}�C<V�?<��;<˧7<
�3<�e/<=A+<'<V�"<��<��<��<��<Wq<g
<*d<gh<Y��;��;�=�;�{�;J��;W�;t�;���;�N�;Mз;�c�;I�;#ҡ;���;R��;)��;Y�;��;�hs;\^g;l�[;�yP;��E;�;;��0;��&;�7;��;.�
;�;���:���:T}�:�y�:��:��:
S�:\9�:�!o:��T:{�::��!:Rz	:D�9n�9La�9�E.9��8�"��"͸Y6C��􏹌N���}칈(�V�#�j:�!�O�yce�aOz��`��-d���9�� ȑ��k0�� �����˺}|պ�ߺڮ����tp���|���	�<��d��������*$��[)��.��3���8�D�=��B��H��9M�fsR�ǿW�; ]�M�b��h�`�m��Vs�'�x�M�~�/������?����G���茻<}������������}���  �  Ɵ=KP=��=;�=c[=F=�=�[==ɭ =]V = ��<�O�<f��<���<HJ�<w��<p��<�K�<*��<��<�L�<"��<N��<@�<%��<���<��<�a�<���<���<�,�<�q�<ظ�<_�<�N�<���< ��<vB�<���<>��<�>�<��<���<m)�<�o�<���<���<'�<�Z�<4��<f��<���<& �<��<+;�<:R�<�d�<`q�<Xx�<lx�<�p�<�`�<�F�<�"�<���<2��<�n�<�<���<OK�<���<�O�<���</�<2��<���<I�<���<E��<�1�<it�<���</�<h�<�A�<�c�<n~�<u��<$��<��<說<o��<t��<Ĝ�<뒢<���<({�<n�<g`�<NR�<�C�<�4�<%�<��<�<�<�ԉ</��<�<}�<�Z�<pm~<�#z<R�u<�q<�Om<�i<�d<��`<	�\<_X<�BT<'+P<sL<�H<v�C<�?<I�;<��7<��3<<i/<G+<�#'<)#<�<��<��<�<��<Uv
<_r<iu<���;��;�M�;���;R��;@�;\t�;���;nG�;0ŷ;dT�;���;Ȼ�;���;ͥ�;k،;5:�;�;�+s;�$g;f�[;NIP;�mE;��:;&�0;�&;�+;��;H�
;��;x�:M2�:��:���:�R�:5P�:XǓ:�:?p:1�U:{�;:̪":!
:�)�9�δ9���9T�.9qg�8��'���θ�kD�{֐�n����������$�c	;���P��ef��O{�U݇�Pؑ�����:N���⮺�u��º`�˺��պ�ߺ������G���_�$�	�,���3��x� ��4�#�� )��J.�o3���8�í=���B���G��)M��kR�s�W��']�G�b��3h�i�m�s|s��(y���~�38������幇�;h��r��ě��8#��	������ꐙ��  �  ��=EO= �=٭=T[=�=��=�\=D=P� =%X =�  =T�<ئ�<H��<�N�<���<T��<=O�<��<K��<�N�</��<���<�?�<C��<��<w�<�^�<J��<1��<�(�<;m�<���<n��<�I�<ʘ�<f��<>�<ϒ�<���<�;�<���<���<?(�<[o�<ݱ�<���<x(�<�\�<Ό�<���<m��<@�<$�<�?�<�V�<�h�<}u�<|�<�{�<�s�<�b�<RH�<\#�<��<���<�m�<"�<3��<@H�<+��<�K�<���<*�<��<���<�C�<���<^��<-�<fp�<���<:�<��<�?�<\b�<�}�<���<���<~��<<"��<���<���<��<��<��<r�<�d�<^V�<�G�<8�<�'�<��<b�<��<�ԉ<���<���<{�<3X�<fg~<�z<<�u<�q<�Em<�i<��d<�`<:w\<�UX<Y:T<�#P<L<��G</�C<$�?<��;<*�7<��3<�k/<�J+<�('<Y#<D�<��<��<7�<ŉ<y
<4{<�}<-�;>,�;�W�;��;q��;�;7t�;4��;B�;k��;�J�;��;ǭ�;���;��;�Ō;)'�;�u;s; g;rc[;G+P;�RE;y�:;b�0;4�&;h#;��;&�
;��;�/�:_R�:���:��:[��:뒢:v�:���:�p:�V:�J<:�"#:�
:w��9�O�9sU�9�X/9���8ћ+�l�ϸlNE�Ai���$������i�
5%���;�F�Q�g��{�_+���"���蛺L���x������f2º��˺١պ��ߺe�����Y.���N���	�������V����X�#�6�(�E(.��N3��q8�Ŕ=��B��G��M�^fR�˿W�G-]��b��Ch�B�m���s�qEy���~�&J�� ���͇�"|��4��
���U5��p����(��\����  �  !�=�N=��=��=@[=�=ϲ=]=�=̯ =�X =� =�U�<}��<��<AP�<,��<���<[P�<���<��<O�<p��<���<�?�<���<���<��<%^�<��<���<	'�<�k�<P��<���<�G�<��<���<�<�<q��<{��<�:�<��<=��<�'�<"o�<Ա�<���<�(�<s]�<���<���<���<��<�%�<GA�<^X�<Sj�<�v�<;}�<�|�<jt�<\c�<�H�<�#�<���<D��<Fm�<|�<u��<>G�<���<EJ�<[��<b(�<I��<���<�A�<Д�<���<w+�<�n�<���<P�<:�<?�<�a�<�}�<���<"��<���<���<��<Ѩ�<Ρ�<���<���<_��<)t�<.f�<�W�<�H�<	9�<m(�<w�<��<��<wԉ<P��<M��<yz�<|W�<Qe~<@z<m�u<��q<�Bm<i<5�d<M�`<�s\<�RX<r7T<(!P<�L<�G<��C<C�?<�;<Ц7<�3<'l/<�K+<l*'<P	#<��<r�<��<��<f�<��
<E~<\�<��;L0�;[�;���;���;��;�s�;Y��;q@�;$��;�G�;(�;ب�;��;��;K��; �;3g;��r;��f;tW[;� P;IE;�:;B�0;Ѽ&;� ;u�;%�
;G�;7�:�]�:~��:��:���:^��:�$�:#�:��p:�HV:2x<:�J#:��
:n�9�|�9�r�9�r/9J��8�c-�g"иO�E�v���y`��N���!f%���;���Q��?g��)|��E���;��� ��m����*��N����<ºA�˺ݦպ��ߺ۟�2��&���H��	�*���
�9K����=�#���(��.��C3��h8��=�8�B���G��M�}eR���W�9/]��b�tHh��m�"�s��Oy�#�~�XP��s���ԇ�����^#�������;�����	.�������  �  ��=EO= �=٭=T[=�=��=�\=D=P� =%X =�  =T�<ئ�<H��<�N�<���<T��<=O�<��<K��<�N�</��<���<�?�<C��<��<w�<�^�<J��<1��<�(�<;m�<���<n��<�I�<ʘ�<f��<>�<ϒ�<���<�;�<���<���<?(�<[o�<ݱ�<���<x(�<�\�<Ό�<���<m��<@�<$�<�?�<�V�<�h�<}u�<|�<�{�<�s�<�b�<RH�<\#�<��<���<�m�<"�<3��<@H�<+��<�K�<���<*�<��<���<�C�<���<^��<-�<gp�<���<:�<��<�?�<\b�<�}�<���<���<~��<<"��<���<���<��<��<��<r�<�d�<^V�<�G�<8�<�'�<��<a�<��<�ԉ<���<���<{�<3X�<fg~<�z<<�u<�q<�Em<�i<��d<�`<:w\<�UX<Z:T<�#P<L<��G<0�C<$�?<��;<*�7<��3<�k/<�J+<�('<Y#<D�<��<��<7�<ŉ<y
<4{<�}<-�;=,�;�W�;��;p��;�;6t�;3��;B�;k��;�J�;��;ǭ�;���;��;�Ō;)'�;�u;s; g;qc[;F+P;�RE;y�:;a�0;4�&;h#;��;&�
;��;�/�:_R�:���:��:[��:뒢:v�:���:�p:�V:�J<:�"#:�
:w��9�O�9sU�9�X/9���8ћ+�l�ϸlNE�Ai���$������i�
5%���;�F�Q�g��{�_+���"���蛺L���x������f2º��˺١պ��ߺe�����Y.���N���	�������V����X�#�6�(�E(.��N3��q8�Ŕ=��B��G��M�^fR�˿W�G-]��b��Ch�B�m���s�qEy���~�&J�� ���͇�"|��4��
���U5��p����(��\����  �  Ɵ=KP=��=;�=c[=F=�=�[==ɭ =]V = ��<�O�<f��<���<HJ�<w��<p��<�K�<*��<��<�L�<"��<N��<@�<%��<���<��<�a�<���<���<�,�<�q�<ظ�<_�<�N�<���< ��<vB�<���<>��<�>�<��<���<m)�<�o�<���<���<'�<�Z�<4��<f��<���<& �<��<+;�<:R�<�d�<`q�<Xx�<lx�<�p�<�`�<�F�<�"�<���<2��<�n�<�<���<OK�<���<�O�<���</�<2��<���<I�<���<E��<�1�<it�<���<0�<h�<�A�<�c�<n~�<u��<%��<��<說<o��<t��<Ĝ�<뒢<���<({�<n�<g`�<NR�<�C�<�4�<%�<��<�<�<�ԉ</��<�<}�<�Z�<pm~<�#z<R�u<�q<�Om<�i<�d<��`<	�\<_X<�BT<(+P<sL<�H<v�C<�?<J�;<��7<��3<=i/<G+<�#'<*#<�<��<��<�<��<Uv
<_r<hu<���;��;�M�;���;Q��;>�;Zt�;���;lG�;/ŷ;bT�;���;ǻ�;���;̥�;j،;4:�;�;�+s;�$g;e�[;MIP;�mE;��:;%�0;�&;�+;��;G�
;��;w�:M2�:��:���:�R�:5P�:XǓ:�:?p:1�U:{�;:̪":!
:�)�9�δ9���9T�.9qg�8��'���θ�kD�{֐�n����������$�c	;���P��ef��O{�U݇�Pؑ�����:N���⮺�u��º`�˺��պ�ߺ������G���_�$�	�,���3��x� ��4�#�� )��J.�o3���8�í=���B���G��)M��kR�s�W��']�G�b��3h�i�m�s|s��(y���~�38������幇�;h��r��ě��8#��	������ꐙ��  �  ġ=�Q=� =��=j[=�=�=wZ==\� =�S =���<�H�<��<s��<�B�<���<>��<PF�<���<S��<;J�<|��<���<Z@�<n��<���<��<�e�<���<���<X3�<y�<���<^
�<�V�<���<���<XI�<���<���</C�<���<7��<+�<�p�<���<���<�$�<�W�<���<S��<���<���<��<�3�<�J�<^]�<�j�<xr�<Zs�<�l�<�]�<�D�<�!�<���<	��<�p�<��<���<!P�<h��<QV�<���<�6�<u��<q��<oQ�<��<���<�8�<�z�<���<��<�<)D�<?e�<#�<?��<螮<ĥ�<���<��<<��<Ŗ�<H��<f��<�s�<�f�<VY�<�K�<>�<�/�<� �<��<���<��<fԉ<��<���<��<{^�<�v~</z<1�u<0�q<�^m<�!i<��d<�`<��\<}mX<PT<�6P<` L<7H<~�C<W�?<��;<̧7<�3<�e/<>A+<'<V�"<��<��<��<��<Wq<g
<*d<fh<X��;��;�=�;�{�;I��;U�;t�;���;�N�;Kз;�c�;G�;!ҡ;���;Q��;(��;
Y�;��;�hs;Z^g;j�[;�yP;��E;�;;��0;��&;�7;��;.�
;�;���:���:T}�:�y�:��:��:	S�:\9�:�!o:��T:z�::��!:Rz	:D�9n�9La�9�E.9��8�"��"͸Y6C��􏹌N���}칈(�V�#�j:�!�O�yce�aOz��`��-d���9�� ȑ��k0�� �����˺}|պ�ߺڮ����tp���|���	�<��d��������*$��[)��.��3���8�D�=��B��H��9M�fsR�ǿW�; ]�M�b��h�`�m��Vs�'�x�M�~�/������?����G���茻<}������������}���  �  >�=�S==^�=_[='=ï=}X= =-� =�O =-��<�?�<���<���<}9�<���<���<?�<a��<h��<�F�<��<���<�@�<���<���<�#�<
k�<��<Q��<�;�<^��<z��<��<a�<���<@ �<@R�<��<}��<�H�<N��<���<C-�<sq�<��<���<�!�<>S�<c��<���<���<��<p�<T*�<gA�<2T�<>b�<�j�<�l�<%g�<=Y�<�A�<��<n��<���<s�<c �<T��<,V�<���<�^�<��<�@�<���<?�<<\�<_��<���<�A�<���<���<��<� �<�G�<ag�<��<���<���<���<��<R��<F��<���<���<w�<Fj�<)]�<.P�<BC�<P6�<>)�<l�<��<���<L�<ԉ<���<��<8��<<c�<Ƃ~<X=z<��u<�q<�rm<6i<X�d<��`<��\<@�X<aT<�EP<-L<�H<N�C<��?<[�;<ۧ7<n�3<3`/<V9+<�'<n�"<!�<H�<�<dn<z]<�S
<�Q<�V<i��;���;(�;�j�;���;�;s�;���;X�;{޷;w�;%�;��;�ך;!�;>�;y��;��;-�s;ɨg;
�[; �P;I�E;?7;;�0;��&;(G;��;z�
;��;��:���:�!�:��:r�:-Z�:E��:���:��m:AyS:W�9:�� :��:ޠ�9�Ҳ9,��9�A-9�e�8����&˸ڙA��ڎ�*缹���A,���"��8���N��d�y�����u͐�/����s���)���ڷ�/���|m˺gaպr}ߺ-���$��e���(����	��P�Ħ�����<��w$��)�%�.���3�8�8�8	>��C��/H�mPM��R���W��]��b�� h�׍m��&s��x�o]~�����p����q���������U��:⑻�f���斻,e���  �  ��=�U=[=�=?[=>=�=V=\� =N� =NK =+��<�4�<G��<[��<U.�<��<,��<Y6�<���<z��<B�<��<��<�@�<S��<}��<5(�<�p�<E��<���<�E�<��<���<s �<�l�<H��<N�<i\�<��<e��<tO�<N��<B��<D/�<%r�<E��<v��<�<�M�<�y�<z��<���<���<��<�<6�<LI�<�W�<Va�<~d�<``�<	T�<>�<��<���<��<Ou�<Q$�<���<�\�<���<h�<���<uL�<5��<��<�h�<��<U�<GL�<7��<!ƻ<R��<�%�<:K�<di�<���<Ӑ�<���<���<���<P��<���<F��<y�<l�<�^�<�Q�<FE�<9�<3-�<9!�<��<i�<[��<$�<vӉ<̼�<G��<!��<|h�<v�~<�Mz<O
v<]�q<"�m<�Mi<me<��`<��\<��X<ltT<�VP<�;L<� H<D<9�?<��;<��7<��3<�Y/<�/+<�'<��"<�<ێ<�o<HW<�E<n<
<F;<�B<̣�;���;,�;�V�;���;��;#q�;,��;�a�;S�;X��;�@�;��;b��;�;,H�;#��;�B�;tt;�g;GM\;i�P;�F;�h;;�1;�';�T;
�;��
;��;g~�:\�:C��:��:Dܯ:v��:R�:u�:�|l:R:��8:��:��:t��9�t�9䏃9,9t�8Ҫ�AXɸ+�?�X���cR��@���@t!���7�SGM���b�f�w��	��� ��d��꣺����z��SO���;˺qIպ�yߺ��麩Q������3���2
�������J������$�~*�-#/��74�bB9�hH>�rMC��WH�lM���R���W��]�"ob���g�>cm�{�r��x�.~�E΁������B��ϐ���(��F���A���Ŗ��H���  �  ͩ=�W=�=i�=�Z==4�=HS=�� =� =nF =E��<#)�<z�<���<*"�<[y�<���<�,�<Ň�<���<�<�<���<��<S@�<���<W��<�,�<�v�<Ϳ�<��<�O�<S��<���<�,�<vy�<���<��<?g�<���<��<,V�<o��<���<D1�<�r�<���<���<��<�G�<3r�<���<���<���<���<��<�)�<`=�<�L�<>W�<�[�<�X�<	N�<�9�<��<���<���<�w�<.(�<��<d�<y��<&r�<��<�X�<��<��<�u�<@��<V�<jW�<��<tλ< �<+�<�N�<qk�<��<z��<���<�<g��<���<݆�<�z�<�m�<`�<�R�<�E�<Z9�<�-�<9#�<p�<��<��<&�<~�<e҉<u��<x��<���<�m�<s�~<�^z<0v<��q<Рm<�fi<�0e<��`<��\<T�X<�T<�hP<�JL<�,H<�D<��?<?�;<��7<�}3<3R/<�$+<��&<��"<5�<�x<�W<(><@,<>#
<#<1,<�{�;Ю�;%��;�?�;|��;���;�m�;7��;�j�;���;��;�\�;m0�;�#�;*9�;5v�;3ކ;?s�;Tot;NWh;��\;0FQ;�EF;��;;�?1;�/';�b;Q�;B�
;ss;H4�:���:V8�:D��:18�:���:�K�:� �:��j:��P:�7:�p:Xm:n��9+�9�e�9P�*9X��8]��_�Ǹ�(>�Bg������\�湒�	�/ �
6��K��a�?�u��H��Xk���j���W��,6��~�� ��?˺}1պ�{ߺL�����$?�����r
�����G�������6%��d*�M�/���4�d�9���>���C���H�c�M���R�(�W�\	]��\b��g��7m�%�r�->x���}�C����]��*��˼��_����������������",���  �  ��=�Y=�=��=[Z=�=�=nP=9� =�� =]A ='��<I�<�m�<_��<��<�m�<���< #�<]�<���<t7�<ő�<���<�?�<���<���<�0�<�|�<��<��<�Y�<g��<���<<9�<݅�<���<g"�<�q�<���<w�<�\�<]��<��<3�<�r�<l��<���<��<�A�<|j�<`��<:��<8��<���<\�<d�<N1�<eA�<�L�<eR�<EQ�<�G�< 5�<��<M��<���<�y�<�+�<V��<�j�<���<�{�<���<�d�<���<+�<��<���<2�<&b�<���<xֻ<��<�/�<R�<2m�<��<㍰<���<%��<���<���<p}�<Lp�<1b�<�S�<F�<(9�<a-�<�"�<��<j�<��<t��<��<��<�Љ<���<j��<i��<s�<߫~<�nz<d1v<�q<m�m<�i<Je<�a<��\<|�X<��T<�yP<�XL<.8H<�D<��?<��;<��7<�x3<�I/<'+<,�&<�"<��<�a<~?<�$<Y<�	
<�
<D<(R�;���;��;�'�;���;S��;eh�;���;�r�;I�;:��;jw�;OQ�;yI�;�c�;���;��;��;��t;�h;	�\;��Q;;�F;��;;�d1;�F';-n;_�;�x
;�X;~��:��:���:e_�:���:3E�:I��:�V�:�Zi:OO:��5:P:@:T��9�E�9C,�9w�(9�0�8b ���Ÿ��<��8��������������,�4��=J�r�_��pt����e����ɘ��ɢ�;�������ؿ����ʺ:պ�ߺ�����l����;�δ
�j-�����XY �i�%�v�*���/���4���9���>��C���H�f�M���R�/�W�]��Kb���g�Fm��r�-�w�Fw}�dw���.��k������<.��tʎ��`��	�l���~���  �  �=5[=�=̰=�Y=z=��=�M=�� =�� =�< =���<��<�a�<|��<
�<b�<;��<��<Nw�<
��<62�<֍�<���<�>�<'��<���<Z4�<���<���<~�<�b�<���<���<�D�<O��<���<�,�<A{�<r��<��<Tb�<���<���<?4�<Tr�<ݫ�<g��<A�<�;�<�b�<���<j��<n��<��<���<��<�%�<�6�<�B�<�I�<�I�<�A�<�0�<��<���<���<�z�<�.�<���<�p�<X �<Մ�<���<�o�<u��<7�<��<z��<')�<�k�<H��<�ݻ<��<D4�<�T�<^n�<���<B��<'��<s��<���<
��<�t�<Hf�<AW�<@H�<1:�<R-�<�!�<��<%�<��<���<���<	�<�ދ<�ω<���<ݨ�<V��<�w�<ѷ~<~z<�Bv<�r<�m<"�i<Xae<�/a<�]<��X<�T<щP<�eL<0BH<�D<o�?<�;<��7<�s3<�A/<+<��&<�"<[w<wL<Y(<S<��<[�	<~�<��<P+�;�h�;���;��;�v�;��;�b�;���;�x�;m�;�ɰ;���;Io�;�k�;���;�͍;9�;(π;#"u;�i;j:];��Q;1�F;C�;;�1;<Z';�u;��;.j
;N=;���:8-�:{=�:�ҽ:��:���:`Ώ:ʗ�:��g:H�M:J4:��:%:a�9���9��9u''9�q�8���b�ĸ�_;��4��\���G*�Q��'���]3���H�0^�ws��ك�.���6���G���T���d��w����ʺ�պ/�ߺ�2�,��������p�t�
�(v�����\�� �|�%�>'+��<0��>5�j0:�2?���C�y�H���M�%�R�x�W�]�X?b���g�s�l��Pr��w��1}�3P���������>]��W��@����8���Γ��b�������  �  ް=�\=B=Ͱ=!Y=, =�=!K=�� =ߓ =o8 =a��<�<�W�<5��<���<�X�<-��<��<<p�<��<v-�<M��<B��<�=�<w��<���<B7�<��<���<�<�j�<6��<��< N�<��<$��<�5�<w��<���<��<
g�<��<��<#5�<�q�<��<f��<�<E6�<]\�<�<ƞ�<��<;��<`��<m�<��<,-�<M:�<B�<:C�<�<�<{,�<��<E��<i��<|�<1�<���<�u�<��<C��<��<y�<H��<5A�<��<8��<Z2�<at�<���<��<W�<�7�<&W�<Ao�<H��<n��<��<&��<*��<Yz�<�l�<~]�<�M�<N>�<�/�< #�<�<��<��<O��<��<E��<��<�ۋ<�͉<R��<海<œ�<K{�<��~<_�z<�Qv<�r<0�m<F�i<�te<�Ba<]<&�X<��T<ݖP<{pL<^JH<F#D<k�?<��;<C�7<~n3<:/<�+<[�&<C�"<Xf<�9<8<{�<��<��	<C�<��<��;�J�;!��;���;�f�;���;�\�;0��;�}�;J"�;|ذ;���;އ�;V��;^��;���;�]�;=�;:ju;�Ei;{y];�R;H�F;�<;ٝ1;j';�z;��;�Z
;�#;�Q�:%��:@��:hU�:Qa�:7��:.�:h�:�f:�UL:�3:�:�):�Z�9:P�9�}99�%9���8*m!��7ĸ�T:��_��ŗ��0�ṟ��ܡ��D2��G��\�M�q��F�����������ܡ���� ���S����ʺ�պ��ߺ3V��3��� �G���+����:8�/��_!��L&��x+��0�H�5�at:��S?�/D��I� �M��R�(�W�%]��5b�Zxg�f�l� )r���w���|��.��
���܍���6��Uۋ�{���������~I��+㘻�  �  J�=r]=�=��=�X='�=��=I=#� =�� =*5 =K��<x �<�O�<��<��<1Q�<5��<8�<�j�<h��<�)�<���<n��<�<�<���<���<O9�<���<��<$�<zp�<���<��<|U�<H��<w��<�<�<���<���<#!�<�j�<���<|��<�5�<q�<���<$��<��<�1�<JW�<y�<��<ô�<w��<i��<r��<-�<�%�<�3�<<�<*>�<38�<3)�<��<���<��<�|�<�2�<O��<�y�<X�<ܑ�<��<��<���<�H�<ʠ�<���<A9�<�z�<���<q�<��<W:�<�X�<�o�<��<���<ȋ�<���<ŀ�<u�<�f�<�V�<LF�<{6�<�'�<'�<U�<l�<���<_��<�<�<��<|ً<�̉< ��<���<j��<�}�<B�~<Ǔz<�\v<0%r<�m<*�i<ǃe<�Qa<:"]<�X<�T<ʠP<�xL<\PH<:'D<C�?<��;<9�7<�j3<=4/<��*<��&<��"<Y<7+<�<,�<�<0�	<��<:�<��;3�;���;��;�Z�;��;�W�; ��;N��;$)�;|�;���;���;H��;�Ô;%�;8z�;��;��u;/yi;=�];�-R;�G;5<;O�1;3t';"};	�;�M
;o;��:��:�:�:t��:]��: ��:Aq�:�e:CYK:�*2:��:�c:��92�9|9aa$9���8A�%���øɪ9��ň�,���0��*�R���p1���F���[���p��ӂ�� ���Z��񋡺Ӹ��~쵺�0���ʺ�	պ�ߺ�q�3]���4 �/��VW�)��{o�>���F!���&���+���0�w�5�=�:���?�~VD�-I�q
N��R���W��]��0b��jg���l��
r��hw�d�|�����ă�jp��W��꽋�__������=���I6���Ә��  �  (�=^=�=��=-X=p�=��=�G=�� =/� =3 =���<���<�J�<��<%��<mL�<���<9�<'g�<g��</'�<���<%��<(<�<���<O��<�:�<׊�<���</'�<t�<���<H�<�Y�<Ħ�<���<�@�<a��<B��<�#�<�l�<.��<r��<�5�<q�<���<y��<��<//�<�S�<Iu�<ѓ�<"��<���<��<���<U�<C!�<X/�<P8�<�:�<z5�<	'�</�<	��<ȹ�<#}�<�3�<���<�{�<I�<h��<��<u��<���<�M�<��<f��<�=�<�~�<p��<E�<�<�;�<�Y�<p�<o�<���<��<s��<�}�<�q�<�b�<`R�<�A�<�1�<�"�<7�<v�<��<���<���<��<S�<��<�׋<�ˉ<���<���<v��<��<��~<��z<�cv<-r<��m<�i<�e<�Za<�*]< �X<U�T<�P<w}L<TH<�)D<��?<��;<��7<�g3<"0/<��*<I�&<N�"<�P<�!<��<�<��<�	<��<��<A��;$�;{�;k��;�Q�;��;HT�;@��;C��;v-�;�;廩;\��;��;LӔ;��;M��;�!�;u�u;��i;��];ZGR;�G;hE<;��1;�z';;�;,E
;S;���:S_�:�H�:���:��:8<�:ga�:�!�:��d: �J:9�1:�Z:?�:3�9�|�9�z9p�#9��8W�)��øL99�Tg��l7����߹˿��h���0��=F��d[�cXp�����ߌ� ��dX������ε�[����ʺպ˳ߺ?��Q{���G ����Zs���ے�*��m!�]�&�I�+���0�1�5���:��?�2pD�BI�zN� S���W��
]��,b��ag�A�l���q�bQw���|��������^��e��+���ON���퐻���;*��=ʘ��  �  ɺ=	f= =ĸ=�_='=�=�K=i� =8� =p1 =���<���<B�<^��<j��<{J�<���<��<�u�<���<�B�<k��<V	�<�g�<-��<�<p�<���<��<Mc�<h��<��<�P�<,��<��<V@�<̐�<��<�0�<��<���<+�<D^�<]��<x��<n�<�K�<�y�<��<���<���<��<'�<D�<�`�<J}�<���<���<?��<���<��<h��<���<^��<���<N��<QR�<8�<���<�T�<���<ck�<���<(U�<���<��<bj�<���<���<�4�<2i�<���<伺<�۸<3�<��<�
�<�<�<���<��<!ͨ<泦<���<��<�g�<�R�<A�<�2�<1(�< �<��<D�<��<�<X��<Z��<�߇<�˅<���<l��<�~<�z<�v<,Cr<|n<��i<`�e<DPa<�]<�X<��T<^~P<�ML<!H<��C<;�?<�};<V@7</�2<B�.<Nm*<�!&<A�!<L�<�O<l<U�<��<�<9�<�� <޴�;N��;�J�;ά�;��;���;��; ��;��;b��;�R�;�;�;�Ҙ;��;��;�w�;y�{;co;!#c;s>W;��K;)�@;Ǯ5;(+;�� ;��;�B;��;��:� �:Rf�:J�:��:B��:"h�:^��:�ug:B�L:�3:sd:�N:q<�9�'�9M�9��:9�'�8�Q�7Ey��W�g�$����ȹ��*��e$�6y9�dN��c���w�Q���!���2���8��8@��4R���yº��̺y4׺���j�캧����|�](�������%�Z���#��Y(�)w-�n2�TB7���;��@��DE���I���N��SS�{-X�m"]��1b�!Zg���l�#�q�4w��|���@����E��wꈻ����c)��kĐ�^�����������  �  n�=�e==ܸ=�_=o=e�=0L=3� =� =d2 =���<���<`D�<���<���<�L�<���<��<�w�<&��<D�<=��<�	�<<h�<C��<��<�o�<���<w�<�a�<ݰ�<���<�N�<)��<��<_>�<��<f��<d/�<o~�<���<��<^�<R��<���<��<rL�<�z�<=��<t��<l��<�
�<)�<aF�<4c�<��<���<���<@��<X��<��<���<���<��<��<���<9R�<�
�<��<�S�<���<�i�<���<,S�<���<��<<h�<q��<���<�2�<�g�<b��<���<C۸<��<��<�<��<��<���<?�<�Ψ<���<���<��<@j�<,U�<oC�<55�<B*�< "�<��<��<��<�<���<���<��<�˅<F��<Ǚ�<�~<y�z<�~v<�?r<� n<��i<7�e<9La<�]<v�X<��T<�{P<�KL<�H<F�C<��?<�};<A7<G�2<�.<�o*<�$&<��!<(�<T<
<!�< �<��<ս<�� <���;T��;XQ�;̱�;8�;���;��;ډ�;��;+��;�O�;
�;�ܟ;�̘;�ݑ;�;�o�;��{;�So;hc;�1W;=�K;�}@;��5;�#+;�� ;��;pE;r�;��:��:�|�:�d�:�ׯ:oߟ:���:D݁:+�g:QM:<�3:��:�:���9���9}_�9�g;9b��8\�7ѣx�hZ��2g��G��oɹk��Y��$�F�9�}�N��`c���w��$���?���K��8O��LR��\_��<�º!�̺�3׺��Ẵ�������s������mw�r�כ��#��G(��d-��[2��17�4�;�:�@��7E���I�ʋN��NS�f*X�� ]�j2b�F\g�ۚl�!�q�Y>w���|��������lM���򈻕���&1��~ː�d�����ϕ���  �  Y�=5e=�=	�=�`=o=̪=�M=T� =�� =75 =ұ�<���<DK�<���<���<+S�<���<�<U|�<:��<gG�<��<��<Di�<m��<;�< n�<���<W�<�]�<$��<B��<�H�<��<���<h8�<?��<c��<+�<�z�<��<��< ]�<��<j��<C�<�N�<�}�<��<���<���<��<^/�<M�<j�<m��<���<��<��<x��<���<r��<���<@��<X��<!��<�Q�<�	�<ٳ�<�P�<��<Je�<���<AM�<b��<[�<�a�<5��<��<�-�<?c�<ؑ�<<��<Yٸ<��<��<��<��<$�<���<�<BӨ<뺦<���<n��<q�<\�<WJ�<�;�<�0�<�'�<� �<O�<l�<�<* �<"�<���<w˅<��<���<m�~<�z<�uv<=5r<��m<}�i<�ye<�?a<�]<��X<5�T<�sP<~EL<	H<Y�C<��?<r~;<9C7<)3<��.<�v*<H-&<��!<��<�`<{*<?�<N�<�<;�<�� <���;��;�b�;*��;�'�;k��;��;���;O�;*��;�G�;���;�͟; ��;ɑ;���;�X�;}�{;�%o;�b;
W;E�K;Yc@;��5;�+;u� ;��;�K;��;C�:�C�:e��:��:+�:�=�:$�:fJ�:R�h:U�M:�4:bs:�M:���9��9QS�9A�<9�A�8�$�7~w��j�x�g�庞���ɹ����5��&8%�vh:��`O��#d�ŭx�)���񗐺j��������������º�̺�2׺?��2�����Z����>��XL�K���h�'�"�_(�<--��&2�: 7�Z�;�Wn@�5E�F�I��tN�>S�/ X��]��5b�8fg�s�l���q�\w�ȼ|�<������qe��������AH������Uv��U�������  �  ��=d=o=?�=fa=�=۬=�P=�� =m� =�9 =���<��<�U�<s��<K�<c]�<+��<��<��<���<�L�<���<L�<�j�<���<�<�k�<���<
�<uW�<w��<���<�?�<Q��< ��<�.�<[��<C��<$�<u�<���<��<C[�<���<6��<Z�<R�<R��<���<���<���<��<G9�<�W�<�t�<2��<(��<���<*��<���<���<5��<���<{��<M��<Ì�<RQ�<��<���<L�<���<�]�<	��<�C�<\��<	�<~W�<P��<���<i%�< \�<���<���<9ָ<.�<L�<��<�<�
�<l��<��<vڨ<5æ<ɪ�<w��<�{�<�f�<U�<IF�<Z:�<�0�<�(�</!�<�<r�<^�<�<R�<�ʅ<#��<u��<��~<�z<Lgv<�$r<��m<�i<�ee<2,a<�\<{�X<��T<�fP<5;L<�H<��C<Ͳ?<�~;<XF7<�3<��.<s�*<�:&<_�!<~�<Wt<�?<2<��<�<k�<i� <���;�2�;�}�;���;I9�;٣�;P�;��;��;蜵;:�;N�;���;᝘;_��;�؊; 3�;s{;	�n;��b;��V;�SK;�6@;Pr5;|�*;�� ;��;�S;1�;P{�:̎�:��:� �:��:_Ѡ:ˏ�:�:�i:GZO:+�5:��:�u:�9灴9�щ9�L?9���8��7�0u����qh��u����ʹ�;��~���8&��;���P��\e�y�y�����!��*��,���ܮ��Ÿ�A�ºf�̺92׺���%h�9P��$2�����j�a�ߙ�A�_x"��'�K�,���1��6�x;�/@�:�D�ӒI��RN��%S��X��]��:b��vg�O�l�(%r�Ōw��|�n/��-���4���?2���ҋ��l��&������6$��D����  �  (�=�b=�=\�=\b=�	=r�=T=�� =`� =:? =���<>�<�c�<y��<�<�j�<]��<�*�<p��<���<S�<���<��<3l�<s��<K�<h�<y��<�<�N�<L��<K��<;3�<j��</��<,"�<|t�<q��<��<Wm�<���<P�<�X�<˟�<���<��<V�<��<��<���< �<|%�<F�<e�<���<��<���<���<���<���<T��<t��<���<h��<���<U��<(P�<��<��<�E�<���<6T�<���<�7�<��<g��<�I�</��<���<_�<�R�<��<���<�Ѹ<��<f�<Y�<��<��<J�<r��<~�<�ͦ<���<v��<,��<�t�<�b�<�S�<G�<B<�<�2�<�)�<Q �<�<J�<d��<��<�Ʌ<G��<ߏ�<�~<ϙz<�Sv<@r<`�m<
�i<�Ke<a<Q�\<��X<�T<�UP<Q-L<NH<��C<|�?<;<�I7<�3<��.<�*<WK&<_"<?�<��<�Z<�1<�<�	<��<�<�%�;[�;d��;���;�N�;+��;��;��;�
�;���;2'�;IѦ;~��;Gw�;�|�;���;K�;5{;czn;Ib;qyV;|K;��?;�D5;�*;E� ;��;`\;O;^��:!��:V��:���:�W�:��:�^�:�̓:ʻk:}Q:��7:�U:�:���9�Ķ9���9�EB9o�8D�7 ;s���6�i��{��zM̹0!�����F�'�|�<��#R��f�%�{��߇�Tڑ�����l����O������ ú�ͺk7׺ݜ�.7캄���� �N����Ʊ�V9�����
"��H'�Eh,��g1�9M6�6;�s�?��D��ZI��'N��S�� X�g]��Db�_�g���l��Xr�D�w�5D}��[��m��M���f�����k����.��<���E���Ϙ��  �  �=z`=�=H�=;c=�=B�=�W=�� =�� =�E =+��<v#�<�s�<���<��<�y�<@��<07�<@��<���<Z�<���<��<�m�<���<��<�c�<��<���<fD�<7��<���<�$�<Ar�<���<@�<of�<���<��<�c�<��<��<@U�<V��<w��<2!�<fZ�<F��<��<���<��<�2�<�T�<~t�<���<��<%��< ��<��<� �<L�<�<���<���<̾�<���<nN�<5�<��<�=�<���<wH�<i��<�(�<u��<J��<�9�<���<#��<R�<3G�<�z�< ��<X̸<�<���<��<�<�<��<���<��<�٦< Ĥ<)��<ۘ�<�<�r�</c�<mU�<mI�<|>�<�3�<*(�<�<f�<���<)�<ȅ<���<��<��~<*�z<�<v<��q<��m<�ji<�,e<y�`<�\<��X<�gT<AP<�L<l�G<��C<��?<>~;<�L7<�3<�.<�*<=^&<"<\�<��<z<QR<�4<M"	<<�<|Z�;��;&��;��;�f�;���;�%�;i��;P�;x��;��;�;n�;[I�;�H�;�q�;�ƃ;��z;=n;��a;lV;��J;s�?;�5;\�*;6� ;.�;c;�;�	�:V�:[�:.T�:'�:~e�:�I�:kȄ:[�m:;"S:��9:�,!:�	:P��9�U�9�ˍ9ʄE9���8�]�7��q�8|�i;k��ˡ��ιyj��B�� )�C�>���S���h��k}�Xʈ�2����~��=1���گ�����Mú�1ͺ�C׺G��N�۶���� ��E�����N�a���6�$�!���&�#�+�$�0���5���:�2�?�:ND��I��M���R��W��]�-Tb�1�g�m���r��x��}�����I��[�������&B���֎��c��MꓻQm����  �  ��=^=A=�=�c=7=�=�[=[=�� =`L ='��<�3�<���<���<�/�<���<���<1D�<f��<��<'a�<н�<��<dn�<���<��<6^�<o��<��<�8�<��<���<��<�a�<��<��<�V�<���<$�<{Y�<���<��<Q�<4��<a��<1#�<�^�<`��<`��<��<��<�@�<�c�<ʄ�<y��<ڿ�<y��<~��<�<��<��<��<���<���<���<?��<�K�<���<\��<�4�<��<�;�<���<��<mz�<���<N(�<�u�<B��<���<�:�<�o�<���<�Ÿ<��<���<��<*�<`�<��<Y�<G��<F�<^Ҥ<���<[��<ו�<҃�<os�<�d�<2W�<jJ�<�=�<80�<!�<I�<X��<��<�Ņ<��<b��<�~<[pz<*#v<
�q<��m<�Ii<�
e<�`<՟\<�sX<
MT<*P<�	L<��G<��C<��?<C|;<;O7<I3<��.<�*<�q&<_6"<��<"�<��<�t<�W<�D	<<<�=<I��;���;��;F1�;�}�;���;�,�;{��;&��;
o�;j��;���;fB�;��;�;4�;ކ�;cz;��m;�ea;7�U;_WJ;�d?;g�4;h�*;C� ;9�;?e;J*;^P�:[��:Ҟ�:��:�ܲ:(H�:�B�:�Ѕ:t�o:xBU:��;:C #:�h:���9��9(�9��H9���8�h�7kq��m��1m�(O��Y$й���
��L�*���@��V�x�j� ��ˉ�8����V�����v�������ú�iͺ1[׺������?i��� ����Js�r��DW����!�@&�)a+��k0��a5��G:�3%?���C� �H�X�M�z�R���W��]��hb���g�NQm��r�Xsx��~��Ɂ�6����<���扻������띑���噖�K���  �  ܪ=_[=�
=M�=Sd=�={�= _=�=a� =�R =���<jC�<��<S��<@�<$��<8��<�P�<4��<��<�g�<L��<&�<�n�<���<��<eX�<|��<	��<�,�<+s�<���<p�<�P�<��<d��<DG�<5��<s��<�N�<ץ�<���<WL�<���<���<�$�<b�<
��<2��<���<�&�<7N�<�r�<ǔ�<��<r��<v��<���<��<��<_�<s�<U�<���<���<s��<I�<���<<��<�+�<���<A.�<���<D�<i�<���<��<�d�<��<(�<�-�<�d�<���</��<�<*��<P�<��<�<��<^�<t�<l�<:�<͢<���<���<_��<j��<�s�<�d�<V�<gG�<�7�<u&�<��<���<�<�<��<G|�<}�~<�Yz<�v<X�q<�mm<�'i<�d<�`<\<UUX<�1T<}P<��K<�G<8�C<W�?<Qy;<�P7<�"3<��.<M�*<-�&<$M"<<��<b�<��<Ez<�f	<�\<o[<���;���;��;�N�;ܒ�;���;"1�;Ê�;��;�Z�;k׭;8i�;��;W�;�Ր;���;�E�;Y�y;i	m;%�`;�;U;��I;�?;�4;V*;�m ;p�;�c;T9;ю�:��:@ �:��:ޝ�:O$�:�5�:�ӆ:�q:�\W:��=:]	%:g#:P��9;��9C��9��K9e��8_��7
�q��lpo�}��Lҹ����W�٤,�;�B�HX�9m��΀��Њ�����K5��ɮ�����ㇺ��ĺ��ͺ�y׺�}���%���^ � �������1���<��� ��%���*��/���4� �9�o�>���C��H�šM�Q�R���W�� ]�Z�b�d�g��m��(s�b�x��o~����Ȅ�����*��/ǌ�RV���ّ�US���ǖ��:���  �  0�=�X=�=}�=ud=�=��=<b=
=u� =�X =�  =�Q�<5��<���< O�<\��<6�<Y\�<��<>�<�m�<��<��<�n�<��<�	�<sR�<���<T��<v!�<f�<V��<��<�@�<���<���<o8�<���<)��<D�<#��<���<uG�<���<���<�%�<�d�<��<	��<��<i1�<{Z�<���<h��</��<���<��<<�<��<d#�<%$�<=�<"
�<���<���<-��<�E�<a��<��<y"�<���<s!�<i��<���<�X�<���<��<5T�<���<�<&!�<4Z�<Ռ�<K��</ܶ<<��<G�<��<�<��<u�<��<i��<��<�ڢ<TȠ<ӵ�<���<���<��<�p�<�`�<�O�<x>�<+�<P�<[��<�߇<���<ꛃ<<u�<l�~<Dz<��u<E�q<nOm<�i<u�d<~�`<9`\<�8X<�T<��O<��K<��G<��C<��?<�u;<�P7<'3<��.<��*<��&<�a"<.0<<��<��<��<��	<z<�v<N��;D�;�6�;i�;���;���;23�;V��;�߼;�E�;��;�D�;�;R��;���;4��;��;�y;i�l;�y`;��T;h�I; �>;�G4;#*;�I ;,�;E^;�B;���:�m�:���:7.�:�L�:��:��:��:t�s:FHY:��?:+�&:��:���9���9ü�9�FN97��8�7P�s����2�q�����PjԹ�k��|U.��kD�]Z��o��ρ��ȋ�����F	���i��6������hiĺ�ͺ��׺G�������2 ��}���
�*������# �?%��c*��w/��4�~9�rv>��pC��pH�e~M��R� �W�:,]��b��%h�.�m��qs��$y���~�g<��?������k�����������z�������_���  �  ѣ=V==��=cd=�=9�=�d=d=�� =�] =' =^�<��<��<�[�<a��<:�<�e�<��<��<2r�<���<�<n�<���<��<�L�<���<���<N�<�Z�<���<���<�2�<���<���<Q+�<���<f��<�:�<`��<���<�B�<���<���<&�<g�<���<���<��<8:�<�d�<��<ͯ�<��<q��<��<��<O%�<7,�<j+�<�!�<��<���<���<���<�B�<���<���<U�<ܝ�<:�<��<��<BJ�<H��<��<�E�<B��<�տ<$�<�P�<턺<��<�׶<?��<�<>�<@ �<� �<?�<�<��<w��<��<�Ԡ<�<a��<P��<���<�z�<?i�<W�<�C�<�.�<:�<���<^އ<���<%��<�n�<W�~<�0z<t�u<��q<�4m<��h<�d<hs`<E\<3X<� T<s�O<��K<żG<�C<H�?<�q;<P7<�)3<F�.<��*<-�&<�r"<PD<�<��<�<��<�	<�<��<��;�2�;pR�;�}�;���;���;�3�;�~�;�Ҽ;�1�;ᠭ;�$�;�Þ;���;	n�;6��;"҂;S�x;{%l;+`;�uT;�DI;z>;�4;G�);#( ;ɟ;wV;>H;`��:p��:]��:ѥ�:�ܴ:Ŕ�:)ϖ:)��:�u:��Z:7,A:B?(:�:v��9_��9�.�9JP9<�8��7�u�SU���s�_���Oֹ�=��-�V�/�PF�˿[���p����w����N��������E���{����ĺ-κa�׺
��(������  ��L���
�"���(�el������$�x�)��/�%4��-9��2>�29C�GH��bM�$�R���W�d9]�a�b�Mh���m�y�s��qy�-�om��^9���������P>��lȏ��C�����\��ۀ���  �  "�=
T=�=õ=5d=�=Z�=�f=�=�� =�a =_
 =8g�<ͺ�<q�<ge�<b��<{�<m�<���<N�<|u�<���<��<�m�<й�<��<�H�<��<���<U�<�Q�<ڕ�<#��<(�<w�<W��<.!�<&{�<���<r3�<8��<���<D?�<C��<^��<&�<Zh�<h��<���<T�<�@�<�l�<���<"��<���<'��<��<o �<&-�<�2�<�0�<�%�<{�<���<���<d��<@�<���<c��<��<)��<n�<#{�<���<2?�<���<���<�:�<ͅ�<7̿<��<II�<�~�<��<�Ӷ<��<�	�<E�<�!�<�#�< �<��<f�<w��<��<mޠ<r̞<&��<���<��<���<�o�<_\�<�G�<R1�<e�<}��<݇<鹅<N��<�i�<�{~<�!z<�u<^qq<�m<�h<��d<�]`<0\<wX<��S<��O<�K<��G<h�C<9�?<�m;<O7<W+3<�/<��*<C�&<B"<�S<5*<�<�<��<�	<�<�<]>�;oL�;g�;Ì�;X��;���;3�;y�;ȼ;k"�;��;�;[��;ib�;FH�;%^�;���;�Vx;��k;��_;r-T;�I;fA>;��3;'�);� ;$�;�N;J;���:j��:�0�:d��:aI�:�:[�:�!�:��v:�#\:�\B:�X):�:0��9U�9�>�9L�Q9���8U�7��w��z���u�=B����׹�%�*8���0�>NG�]��9r��[���H���햺�S��P���ﴲ��׻�BźMaκ��׺ԚẀ��֤������:(��d
�X��0���$��Z�M�$�A�)�y�.���3���8�>�=��C�%)H�MOM���R���W� E]��b�~lh�m"n���s���y�Gr�����]b��R!���Ί�i����Cj��"֔�W:������  �  n�=�R=�=0�=d=A=�=�g=b=�� =�c = =m�<���<��<gk�<��<��<�q�<���<!�<�w�<��<�<m�<��<� �<�E�<p��<���<O
�<�K�<���<r��<&!�<(p�<��<��<&u�<���<�.�<G��<���<�<�<���<r��< &�<!i�<��<	��<��<�D�<|q�<-��<��<���<1��<��<�%�<�1�<�6�<4�<*(�<�<���<���<_��<=>�<���<��<��<J��<��<�t�<���<8�<���<i��<�3�<2�<ƿ<�<�D�<�z�<ǩ�<SѶ<�<		�<R�<�"�<�%�<#�<"�<��<i�<��<Z�<�Ҟ<0��<s��<���<W��<�s�<�_�<J�<�2�< �<]��<܇<��<���<Rf�<js~<
z<�u<eq<�m<6�h<�d<�O`<�"\<��W<?�S<��O<_�K<��G<��C<�?<�k;<XN7<Z,3<g/<)�*<B�&<�"<�\<5<�<v�<r�<��	<Ʊ<ש<0Q�;/\�;ys�;��;S��;���;@2�;�t�;���;��;�~�;���;H��;WL�;S0�;XD�;͍�;e!x;��k;k�_;�S;a�H;�>;ʿ3;�);��;�;�H;�J;�:��:|Y�:�4�:���:mb�:���:뀉:V�w:��\:�C:]*:��:4��9��9���9v�R96��8���7Qy�*A�{�v�
����عĸ����!�1��H�_�]��s��ʃ������Q��ܰ���᩺�������:ź�κ�׺���ȃ�P���������`H
����ž�����*�jX$��})�֜.�ǵ3�$�8���=�M�B��H�rCM�ڃR�6�W��M]��b��h�=n��t�&�y�X�����T|���<���ꊻ�������ł���씻�M��⫙��  �  ՞=5R=j=�=�c=M=7�=�g=�=Y� =�d =� =�n�<���<��<`m�<
��<Y�<s�<���<"�<&x�<R��<�<�l�<��< �<�D�<'��<���<��<�I�<���<-��<��<�m�<"��<��<s�<���<&-�<ԉ�<���<�;�< ��< ��<�%�<Li�<���<���<��<bF�<s�<��<���<���<9��<��<�'�<�3�<i8�<A5�<)�<��<���<���<���<�=�<.��<׀�<F�<���<��<�r�<���<�5�<<��< ��<�1�<}�<�ÿ<=�<�B�<<y�<���<�ж<��<��<H�<�"�<&�<�#�<U�<�<�<���<M�<�Ԟ<1<f��<[��<䈖<)u�<�`�<�J�<M3�<C�<I��<�ۇ<���<܏�<+e�<Vp~<�z<V�u<�`q<em<m�h<_�d<�J`<"\<��W<_�S<�O<(�K<�G<��C<�?<�j;<�M7<�,3</<��*<Z�&<Ɖ"<�_<�8<�<��<��<��	<Ե<|�<�W�;�a�;�w�;���;���;��;�1�;�s�;���;I�;z�;���;ŋ�;�D�;p(�;�;�;ل�;�x;S�k;��_;R�S;~�H;>;��3;��);�;�~;vF;K;{�:� �:�g�:�G�:ң�:|�:�җ:���:��w:�)]:7ZC:AH*:u�:� �9F6�9b�9K�R9u��8��7��y��z��Ew��O��H!ٹ����p�1�E]H�6^�`s�Lٍ��r��JР���������'��QKźi�κ�غ
����ŏ�������
�[>
��w�#��I��2��G$��m)�O�.�3�3��8���=���B��H�v@M���R��W�CP]��b���h�lFn�t���y�<��a���I���MF��s��������������T��#����  �  n�=�R=�=0�=d=A=�=�g=b=�� =�c = =m�<���<��<gk�<��<��<�q�<���<!�<�w�<��<�<m�<��<� �<�E�<p��<���<O
�<�K�<���<r��<&!�<(p�<��<��<&u�<���<�.�<G��<���<�<�<���<r��< &�<!i�<��<	��<��<�D�<|q�<-��<��<���<1��<��<�%�<�1�<�6�<4�<*(�<�<���<���<_��<=>�<���<��<��<J��<��<�t�<���<8�<���<i��<�3�<2�<ƿ<�<�D�<�z�<ǩ�<TѶ<�<
	�<R�<�"�<�%�<#�<"�<��<i�<��<Z�<�Ҟ<0��<s��<���<W��<�s�<�_�<J�<�2�<�<]��<܇<��<���<Rf�<js~<
z<�u<eq<�m<6�h<�d<�O`<�"\<��W<?�S<��O<_�K<��G<��C<�?<�k;<XN7<Z,3<g/<)�*<B�&<�"<�\<5<�<v�<r�<��	<Ʊ<ש<0Q�;.\�;ys�;��;R��;���;?2�;�t�;���;��;�~�;���;G��;VL�;S0�;WD�;̍�;d!x;��k;j�_;�S;`�H;�>;ʿ3;�);��;�;�H;�J;�:��:|Y�:�4�:���:mb�:���:뀉:V�w:��\:�C:]*:��:4��9��9���9v�R96��8���7Qy�*A�{�v�
����عĸ����!�1��H�_�]��s��ʃ������Q��ܰ���᩺�������:ź�κ�׺���ȃ�P���������`H
����ž�����*�jX$��})�֜.�ǵ3�$�8���=�M�B��H�rCM�ڃR�6�W��M]��b��h�=n��t�&�y�X�����T|���<���ꊻ�������ł���씻�M��⫙��  �  "�=
T=�=õ=5d=�=Z�=�f=�=�� =�a =_
 =8g�<ͺ�<q�<ge�<b��<{�<m�<���<N�<|u�<���<��<�m�<й�<��<�H�<��<���<U�<�Q�<ڕ�<#��<(�<w�<W��<.!�<&{�<���<r3�<8��<���<D?�<C��<^��<&�<Zh�<h��<���<T�<�@�<�l�<���<"��<���<'��<��<o �<&-�<�2�<�0�<�%�<{�<���<���<d��<@�<���<c��<��<)��<o�<#{�<���<2?�<���<���<�:�<΅�<8̿<��<II�<�~�<��<�Ӷ<��<�	�<E�<�!�<�#�< �<��<f�<w��<��<mޠ<r̞<&��<���<��<���<�o�<_\�<�G�<R1�<d�<|��<݇<鹅<M��<�i�<�{~<�!z<�u<]qq<�m<�h<��d<�]`<0\<xX<��S<��O<�K<��G<h�C<:�?<�m;< O7<X+3<�/<��*<D�&<C"<�S<5*<�<�<��<�	<�<�<\>�;nL�;g�;�;W��;���;3�;y�;ȼ;i"�;��;�;Y��;gb�;DH�;$^�;���;�Vx;��k;��_;q-T;�I;eA>;��3;'�);� ;#�;�N;J;���:i��:�0�:d��:aI�:�:[�:�!�:��v:�#\:�\B:�X):�:0��9U�9�>�9L�Q9���8U�7��w��z���u�=B����׹�%�*8���0�>NG�]��9r��[���H���햺�S��P���ﴲ��׻�BźMaκ��׺ԚẀ��֤������:(��d
�X��0���$��Z�M�$�A�)�y�.���3���8�>�=��C�%)H�MOM���R���W� E]��b�~lh�m"n���s���y�Gr�����]b��R!���Ί�i����Cj��"֔�W:������  �  ѣ=V==��=cd=�=9�=�d=d=�� =�] =' =^�<��<��<�[�<a��<:�<�e�<��<��<2r�<���<�<n�<���<��<�L�<���<���<N�<�Z�<���<���<�2�<���<���<Q+�<���<f��<�:�<`��<���<�B�<���<���<&�<g�<���<���<��<8:�<�d�<��<ͯ�<��<q��<��<��<O%�<8,�<j+�<�!�<��<���<���<���<�B�<���<���<U�<ݝ�<:�<��<��<BJ�<I��<��<�E�<B��<�տ<%�<�P�<턺<��<�׶<@��<�<>�<@ �<� �<?�<�<��<w��<��<�Ԡ<�<a��<O��<���<�z�<>i�<W�<�C�<�.�<9�<���<^އ<���<%��<�n�<V�~<�0z<s�u<��q<�4m<��h<�d<hs`<E\<3X<� T<t�O<��K<ƼG<�C<I�?<�q;<P7<�)3<H�.<��*<.�&<�r"<QD<�<��<�<��<�	<�<��<��;�2�;nR�;�}�;���;���;�3�;�~�;�Ҽ;�1�;ޠ�;�$�;�Þ;���;n�;4��;!҂;P�x;y%l;)`;�uT;�DI;z>;�4;F�);"( ;ȟ;vV;=H;_��:o��:]��:Х�:�ܴ:Ŕ�:)ϖ:)��:�u:��Z:7,A:B?(:�:v��9_��9�.�9JP9<�8��7�u�SU���s�_���Oֹ�=��-�V�/�PF�˿[���p����w����N��������E���{����ĺ-κa�׺
��(������  ��L���
�"���(�el������$�x�)��/�%4��-9��2>�29C�GH��bM�$�R���W�d9]�a�b�Mh���m�y�s��qy�-�om��^9���������P>��lȏ��C�����\��ۀ���  �  0�=�X=�=}�=ud=�=��=<b=
=u� =�X =�  =�Q�<5��<���< O�<\��<6�<Y\�<��<>�<�m�<��<��<�n�<��<�	�<sR�<���<T��<v!�<f�<V��<��<�@�<���<���<o8�<���<)��<D�<#��<���<uG�<���<���<�%�<�d�<��<	��<��<i1�<{Z�<���<h��</��<���<��<<�<��<d#�<%$�<=�<"
�<���<���<-��<�E�<a��<��<y"�<���<s!�<i��<���<�X�<���<��<6T�<���<�<&!�<4Z�<֌�<L��<0ܶ<=��<H�<��<�<��<v�<��<j��<��<�ڢ<TȠ<ӵ�<���<���<��<�p�<�`�<�O�<w>�<+�<P�<Z��<�߇<���<ꛃ<<u�<k�~<Dz<��u<D�q<mOm<�i<u�d<~�`<9`\<�8X<�T<��O<��K<��G<��C<��?<�u;<�P7<'3<��.<��*<��&<�a"<.0<<��<��<��<��	<z<�v<L��;B�;�6�;i�;���;���;/3�;S��;�߼;�E�;��;�D�;�;O��;���;1��;��;�y;f�l;�y`;�T;f�I;�>;�G4;#*;�I ;+�;D^;�B;���:�m�:���:7.�:�L�:��:��:��:t�s:FHY:��?:+�&:��:���9���9ü�9�FN97��8�7P�s����2�q�����PjԹ�k��|U.��kD�]Z��o��ρ��ȋ�����F	���i��6������hiĺ�ͺ��׺G�������2 ��}���
�*������# �?%��c*��w/��4�~9�rv>��pC��pH�e~M��R� �W�:,]��b��%h�.�m��qs��$y���~�g<��?������k�����������z�������_���  �  ܪ=_[=�
=M�=Sd=�={�= _=�=a� =�R =���<jC�<��<S��<@�<$��<8��<�P�<4��<��<�g�<L��<&�<�n�<���<��<eX�<|��<	��<�,�<+s�<���<p�<�P�<��<d��<DG�<5��<s��<�N�<ץ�<���<WL�<���<���<�$�<b�<
��<2��<���<�&�<7N�<�r�<ǔ�<��<r��<v��<���<��<��<_�<s�<U�<���<���<s��<I�<���<=��<�+�<���<B.�<���<D�<i�<���<��<�d�<��<(�<�-�<�d�<���<0��<�<+��<Q�<��<�<��<_�<u�<l�<;�<͢<���<���<_��<j��<�s�<�d�<V�<fG�<�7�<t&�<��<���<�<�<��<G|�<{�~<�Yz<�v<W�q<�mm<�'i<�d<�`<\<UUX<�1T<~P<��K< �G<:�C<X�?<Sy;<�P7<�"3<��.<N�*</�&<%M"<<��<c�<��<Ez<�f	<\<n[<���;���;��;�N�;ْ�;���;1�;���;��;�Z�;h׭;5i�;��;T�;�Ր;���;�E�;U�y;f	m;"�`;�;U;��I;�?;�4;V*;�m ;o�;�c;T9;Ў�:��:? �:��:ݝ�:O$�:�5�:�ӆ:�q:�\W:��=:]	%:f#:P��9;��9C��9��K9e��8^��7
�q��lpo�}��Lҹ����W�٤,�;�B�HX�9m��΀��Њ�����K5��ɮ�����ㇺ��ĺ��ͺ�y׺�}���%���^ � �������1���<��� ��%���*��/���4� �9�o�>���C��H�šM�Q�R���W�� ]�Z�b�d�g��m��(s�b�x��o~����Ȅ�����*��/ǌ�RV���ّ�US���ǖ��:���  �  ��=^=A=�=�c=7=�=�[=[=�� =`L ='��<�3�<���<���<�/�<���<���<1D�<f��<��<'a�<н�<��<dn�<���<��<6^�<o��<��<�8�<��<���<��<�a�<��<��<�V�<���<$�<{Y�<���<��<Q�<4��<a��<1#�<�^�<`��<`��<��<��<�@�<�c�<ʄ�<y��<ڿ�<y��<~��<�<��<��<��<���<���<���<?��<�K�<���<\��<�4�<��<�;�<���<��<nz�<���<N(�<�u�<C��<���<�:�<�o�<���<�Ÿ<��<���<��<+�<a�< �<Y�<H��<G�<^Ҥ<���<\��<ו�<҃�<os�<�d�<1W�<iJ�<�=�<70�<!�<H�<X��<��<�Ņ<��<a��<�~<Zpz<)#v<	�q<��m<�Ii<�
e<�`<֟\<�sX<MT<*P<�	L<��G<��C<��?<E|;<=O7<K3<��.<�*<�q&<`6"<��<#�<��<�t<�W<�D	<<<�=<G��;���;��;C1�;�}�;���;|,�;w��;"��;o�;g��;���;cB�;��;��;4�;܆�;_z;��m;�ea;4�U;\WJ;�d?;e�4;f�*;A� ;9�;>e;I*;]P�:[��:Ҟ�:��:�ܲ:'H�:�B�:�Ѕ:t�o:xBU:��;:C #:�h:���9��9(�9��H9���8�h�7kq��m��1m�(O��Y$й���
��L�*���@��V�x�j� ��ˉ�8����V�����v�������ú�iͺ1[׺������?i��� ����Js�r��DW����!�@&�)a+��k0��a5��G:�3%?���C� �H�X�M�z�R���W��]��hb���g�NQm��r�Xsx��~��Ɂ�6����<���扻������띑���噖�K���  �  �=z`=�=H�=;c=�=B�=�W=�� =�� =�E =+��<v#�<�s�<���<��<�y�<@��<07�<@��<���<Z�<���<��<�m�<���<��<�c�<��<���<fD�<7��<���<�$�<Ar�<���<@�<of�<���<��<�c�<��<��<@U�<V��<w��<2!�<fZ�<F��<��<���<��<�2�<�T�<~t�<���<��<%��< ��<��<� �<L�<��<���<���<̾�<���<nN�<5�<��<�=�<���<wH�<j��<�(�<u��<J��<�9�<���<$��<R�<4G�<�z�<!��<Y̸<�<���<��<�<�<��<���<��<�٦<!Ĥ<)��<ۘ�<�<�r�</c�<mU�<lI�<{>�<�3�<)(�<�<e�<���<)�<ȅ<���<��<��~<)�z<�<v<��q<��m<�ji<�,e<y�`<�\<��X<�gT<AP<�L<n�G<��C<��?<?~;<�L7<�3<�.<�*<>^&<"<]�<��<z<QR<�4<M"	<<�<{Z�;��;$��;��;�f�;���;�%�;f��;L�;u��;��;�;n�;XI�;�H�;�q�;�ƃ;��z;:n;��a;jV;�J;q�?;�5;Z�*;5� ;-�;c;�;�	�:V�:Z�:.T�:&�:}e�:�I�:kȄ:[�m:;"S:��9:�,!:�	:P��9�U�9�ˍ9ʄE9���8�]�7��q�8|�i;k��ˡ��ιyj��B�� )�C�>���S���h��k}�Xʈ�2����~��=1���گ�����Mú�1ͺ�C׺G��N�۶���� ��E�����N�a���6�$�!���&�#�+�$�0���5���:�2�?�:ND��I��M���R��W��]�-Tb�1�g�m���r��x��}�����I��[�������&B���֎��c��MꓻQm����  �  (�=�b=�=\�=\b=�	=r�=T=�� =`� =:? =���<>�<�c�<y��<�<�j�<]��<�*�<p��<���<S�<���<��<3l�<s��<K�<h�<y��<�<�N�<L��<K��<;3�<j��</��<,"�<|t�<q��<��<Wm�<���<P�<�X�<˟�<���<��<V�<��<��<���< �<|%�<F�<e�<���<��<���<���<���<���<T��<t��<���<h��<���<U��<(P�<��<��<�E�<���<7T�<���<�7�<��<g��<�I�</��<���<`�<�R�<��<���<�Ѹ<��<g�<Z�<��<��<K�<s��<�<�ͦ<���<v��<,��<�t�<�b�<�S�<G�<B<�<�2�<�)�<P �<�<I�<d��<��<�Ʌ<G��<ޏ�<�~<Ιz<�Sv<?r<`�m<
�i<�Ke<a<R�\<��X<�T<�UP<R-L<OH<��C<}�?<;<�I7<�3<��.<�*<XK&<`"<@�<��<�Z<�1<�<�	<��<�<�%�;[�;b��;���;�N�;(��;��;��;�
�;�;/'�;FѦ;|��;Ew�;�|�;���;I�;2{;`zn;Ib;oyV;zK;��?;�D5;�*;E� ;��;_\;O;]��: ��:U��:���:�W�:��:�^�:�̓:ʻk:}Q:��7:�U:�:���9�Ķ9���9�EB9o�8D�7 ;s���6�i��{��zM̹0!�����F�'�|�<��#R��f�%�{��߇�Tڑ�����l����O������ ú�ͺk7׺ݜ�.7캄���� �N����Ʊ�V9�����
"��H'�Eh,��g1�9M6�6;�s�?��D��ZI��'N��S�� X�g]��Db�_�g���l��Xr�D�w�5D}��[��m��M���f�����k����.��<���E���Ϙ��  �  ��=d=o=?�=fa=�=۬=�P=�� =m� =�9 =���<��<�U�<s��<K�<c]�<+��<��<��<���<�L�<���<L�<�j�<���<�<�k�<���<
�<uW�<w��<���<�?�<Q��< ��<�.�<[��<C��<$�<u�<���<��<C[�<���<6��<Z�<R�<R��<���<���<���<��<G9�<�W�<�t�<2��<(��<���<*��<���<���<5��<���<{��<M��<Č�<SQ�<��<���<L�<���<�]�<	��<�C�<\��<	�<W�<P��<���<i%�< \�<���<���<:ָ</�<M�<��<�<�
�<m��<��<vڨ<6æ<ɪ�<w��<�{�<�f�<U�<IF�<Z:�<�0�<�(�<.!�<�<r�<]�<�<Q�<�ʅ<#��<t��<��~<�z<Lgv<�$r<��m<�i<�ee<2,a<�\<{�X<��T<�fP<6;L<�H<��C<β?<�~;<YF7<�3<��.<s�*<�:&<`�!<�<Xt<�?<2<��<�<k�<i� <���;�2�;�}�;���;G9�;ף�;N�;��;��;朵;:�;L�;���;ޝ�;]��;�؊;�2�;s{;�n;��b;��V;~SK;�6@;Nr5;{�*;�� ;��;�S;1�;O{�:ˎ�:��:� �:��:_Ѡ:ˏ�:�:�i:GZO:+�5:��:�u:�9灴9�щ9�L?9���8��7�0u����qh��u����ʹ�;��~���8&��;���P��\e�y�y�����!��*��,���ܮ��Ÿ�A�ºf�̺92׺���%h�9P��$2�����j�a�ߙ�A�_x"��'�K�,���1��6�x;�/@�:�D�ӒI��RN��%S��X��]��:b��vg�O�l�(%r�Ōw��|�n/��-���4���?2���ҋ��l��&������6$��D����  �  Y�=5e=�=	�=�`=o=̪=�M=T� =�� =75 =ұ�<���<DK�<���<���<+S�<���<�<U|�<:��<gG�<��<��<Di�<m��<;�< n�<���<W�<�]�<$��<B��<�H�<��<���<h8�<?��<c��<+�<�z�<��<��< ]�<��<j��<C�<�N�<�}�<��<���<���<��<^/�<M�<j�<m��<���<��<��<x��<���<r��<���<@��<X��<!��<�Q�<�	�<ٳ�<�P�<��<Je�<���<AM�<b��<\�<�a�<5��<��<�-�<?c�<ّ�<=��<Yٸ<��<��<��< �<$�<���<�<CӨ<캦<���<n��<q�<\�<WJ�<�;�<�0�<�'�<� �<N�<l�<�<* �<!�<���<v˅<��<���<l�~<�z<�uv<<5r<��m<}�i<�ye<�?a<�]<��X<5�T<�sP<EL<
H<Z�C<��?<s~;<9C7<)3<��.<�v*<I-&<��!<��<�`<{*<?�<N�<�<;�<�� <���;��;�b�;)��;�'�;j��;��;���;N�;(��;�G�;���;�͟;���;�ȑ;���;�X�;{�{;�%o; �b;W;D�K;Xc@;��5;�+;t� ;��;�K;��;C�:�C�:e��:��:+�:�=�:#�:fJ�:R�h:U�M:�4:bs:�M:���9��9QS�9A�<9�A�8�$�7~w��j�x�g�庞���ɹ����5��&8%�vh:��`O��#d�ŭx�)���񗐺j��������������º�̺�2׺?��2�����Z����>��XL�K���h�'�"�_(�<--��&2�: 7�Z�;�Wn@�5E�F�I��tN�>S�/ X��]��5b�8fg�s�l���q�\w�ȼ|�<������qe��������AH������Uv��U�������  �  n�=�e==ܸ=�_=o=e�=0L=3� =� =d2 =���<���<`D�<���<���<�L�<���<��<�w�<&��<D�<=��<�	�<<h�<C��<��<�o�<���<w�<�a�<ݰ�<���<�N�<)��<��<_>�<��<f��<d/�<o~�<���<��<^�<R��<���<��<rL�<�z�<=��<t��<l��<�
�<)�<aF�<4c�<��<���<���<@��<X��<��<���<���<��<��<���<9R�<�
�<��<�S�<���<�i�<���<,S�<���<��<<h�<q��<���<�2�<�g�<c��<���<D۸<��<��<�<��<��<���<@�<�Ψ<���<���<��<@j�<,U�<oC�<55�<B*�< "�<��<��<��<�<���<���<��<�˅<E��<Ǚ�<�~<y�z<�~v<�?r<� n<��i<7�e<9La<�]<w�X<��T<�{P<�KL<�H<F�C<��?<�};<A7<G�2<�.<�o*<�$&<��!<(�<T<
<!�< �<��<ս<�� <���;T��;XQ�;˱�;8�;���;��;ى�;��;*��;�O�;
�;�ܟ;�̘;�ݑ;�;�o�;��{;�So;gc;�1W;<�K;�}@;��5;�#+;�� ;��;pE;r�;��:��:�|�:�d�:�ׯ:nߟ:���:D݁:+�g:QM:<�3:��:�:���9���9}_�9�g;9b��8\�7ѣx�hZ��2g��G��oɹk��Y��$�F�9�}�N��`c���w��$���?���K��8O��LR��\_��<�º!�̺�3׺��Ẵ�������s������mw�r�כ��#��G(��d-��[2��17�4�;�:�@��7E���I�ʋN��NS�f*X�� ]�j2b�F\g�ۚl�!�q�Y>w���|��������lM���򈻕���&1��~ː�d�����ϕ���  �  ��=Xo=�=?�=�h=�=î=8O=�� =�� =- =���<���<2�<��<���<�A�<Ȩ�<�<��<���<�^�<`��<w2�<.��<���<�P�<*��<���<�O�<[��<���<�C�<���<1��<>;�<���<���<�6�<���<#��<�/�<�~�<<��<3�<\R�<e��<���<��<��<�<�<�]�<}�<ܛ�<"��<���<��<� �<�C�<�d�<v��<ޙ�<��<E��<7��<���<gi�<y4�<���<��<�9�<���<oM�<���<1�<Β�<���<=9�<�<��<��<"�<�I�<fj�<V��<J��<��<ʜ�<��<���<pj�<�K�<�(�<��<�ݤ<׹�<ۘ�<�|�<�e�<wT�<AH�<2@�<7;�<f7�<k3�<v-�<�$�<v�<��<��<�Ճ<���<%/<��z<�v<�\r<Mn<��i<��e<�Ga<�]<�X<ۏT<�WP<< L< �G<��C<�r?<0;<�6<��2<�>.<��)<��%<�!!<��<�o<�%<��<n�<U�<�<C�;�n�;��;!�;�h�;V��;@�;���;)#�;К�;��;��;M�;6�;W��;ێ;���;|E�;�vu;��h;Ye\;�nP;��D;@�9;��.;
R$;�;~5;y�;1$�:ɢ�:l��:��:U��:x�:��:�ǂ:}h:%	M:�)3: �:��:�J�9�ֲ9l̊9KMG9L��8��08��KE��WB��0�������Yݹ������N-���A�XrV�[�j���~��m��cV���1��*���ְ�õ���ĺ��κY5ٺ&�������w��d|�lQ�:#����с�P�$�9*�+H/��!4���8�OS=�`�A��$F�|�J�O���S��JX��#]� b�q<g��pl�ѷq��w�\^|��ـ�Ձ���&���ǈ��e��l��������)������oQ���  �  �=(o=�=_�=�h=5=r�=P=�� =� =�. ={��<���<'5�<��<���<�D�<���<��<?��<���<q`�<���<W3�<ǖ�<���<P�<���<���<9N�<{��<o��<�A�<1��<���<�8�<+��<R��<�4�<��<���<�.�<#~�< ��<'�<�R�<��<���<���<��<?�<W`�<��<���<E��<���<	�<�#�<�F�<�g�<ׄ�<��<ê�<���<1��<���<�i�<_4�<h��<H��<�8�<T��<[K�<���<�.�<��<���<n6�<\|�<`��<���< �<:H�<7i�<���<���<���<>��<ϔ�<��<�k�<�M�<+�<�<��<���<��<��<�h�<�W�<"K�<�B�<�=�<�9�<;5�<�.�<�%�<,�<N�<��<LՃ<-��<�,<\�z<�v<Xr<>n<��i<�e<{Ba<�]<��X<��T<�SP<�L<#�G<ͮC<|r?<�0;<Q�6<�2<�A.<n�)<Յ%<1&!<M�<�u<,<+�<��<�<��<�N�;gy�;X��;��;p�;���;D�;���;3$�;���;l�;���;�G�;'�;]ؕ;Ҏ;��;S;�;�au;��h;kR\;^P;]�D;*�9;!�.;�L$;y;�5;k�;�0�:}��: ��:���:�Ѳ:�6�:�<�:���:w�h:�jM:s�3:)1:`=:��9>r�9�T�9�CH9��8�38���⸣XB��<���Ƴ��ݹ���-����-��CB��V�k��6�����t|��8S��� ��{��ƺ��ĺ��κ4ٺ�㺳��8���Y��Nl�@�����4j���$�!*�C//�	4���8��==��A��F�Q}J���N�*�S��EX�!]�� b�/?g�wwl���q�aw��n|��※ڋ��V1���҈�$p���	��۞���1���Õ��V���  �  ��=xn=�=��=�i=�=\�=lR=~� =:� =�2 =��<���<�>�<���< ��<�M�<��<%�<���<Z��<�d�<;��<�5�<h��<K��<�O�< ��<��<UJ�<f��<U��<�:�<f��<Q��<30�<*��<���<-.�<i��<!��<G+�<�{�<��<-�<�S�<C��<%��<���<��<#E�<[g�<�<K��<k��<e��<r
�</-�<JO�<�o�<��<���<���<ǲ�<F��<���<�j�<>4�<D��<���<5�<���<�E�<���<�&�<���<��<�-�<t�<���<%��<i�<�C�<�e�<o��< ��<���<k��<���<F��<p�<�R�<?1�<K�<��<hŢ<Y��<N��<mr�<�`�<�S�<�J�<oD�<�?�<&:�<�2�<�(�<;�<R�<��<$ԃ<���<�%<�z<j�v<bJr<� n<V�i<�se<�1a<��\<��X<�T<�IP<�L<��G<��C<�q?<52;<��6<�2<.I.<��)<g�%<�3!<��<Æ<j><�<��<I�<�<Sq�;Ә�;���;S'�;���;���;�O�;���;�'�;��;/�;v��;�9�;$�;<��;���;�Ӈ;��;K!u;�kh;�\;}+P;��D;�z9;��.;�<$;[;_7;��;�U�:x��:��:�M�:F4�:먢:l��:䀃:�
j:ΛN:�4:�Z:�R:��9�=�9�ߌ9x�J9�M�8�98�~�J���EB��r��IL���o޹�U�m��b.��/C���W� l������yڶ���s��w-��t�����ĺ]�κ�-ٺط�J�� ���)��'A�6�������1$���$���)�`�.���3�r8�C�<��wA���E��VJ�P�N��vS�6X��]�a"b�Ig�j�l��q��;w��|�����G����Q��K􈻶���5(��t���cI���֕�-e���  �  ��=3m=2=?�=k=�=C�=V=� =�� =�8 =��<��<:M�<_��<���<�[�<���<�)�<��< �<�k�<���<�9�<���<���<�N�<��<b��<�C�<��<D��</�<�<T��<#�<}w�<��<r#�<Kz�<���<�%�<4x�<��<�<gU�<W��<���<��<�'�<�N�<Ur�<	��<ʴ�<���<��<&�<Y;�<�\�<�{�<ٖ�<���<���<���<��<���<l�<�3�<��<ݔ�<</�<��<�;�<s��<Y�<pz�<U��<��<�f�<���<4��<1�<T<�<O`�<�|�<��<蜵<埳<��<!��<�v�<[�<;�<v�<A��<Ӣ<���<��<��<�n�<a�<�V�<UO�<�H�<�A�<'9�<:-�<)�<��<o�<�у<İ�<�<�z<R�v<04r<��m<j�i<lYe<�a<1�\<͠X<�kT<Z9P<�L<j�G<�C<�o?<�3;<��6<�2<�T.<��)<��%<
I!<��<��<)[<p!<p�<(�<��<&��;b��;5�;PL�;,��;  �;�a�;���;�,�;��;��;��;�!�;�Μ; ��;]��;���;��;,�t;
h;��[;��O;�[D;�B9;a�.;�!$;(;^9;�;#��:�8�:uK�:���:�г:~[�:���:�[�:��k:�vP:��6:�%:�	:S#�9�	�9�V�9|�N9n��8�C8t���D�߸�3B�u㊹�+����߹V<�h����/���D�;VY�W�m�1���hڊ�~����Z��g���h���D��[	ź��κ7&ٺ���6S�S��]I�_����qx�~$�]��U $��^)�n.�xO3�\8��<��!A��E�mJ���N��SS�/ X��]��%b��[g���l��r�zw��|��)��dڃ������(��;ċ��X��琻8p�������}���  �  ��=Wk=u=��=�l=)=ŷ=�Z=�� =6� =3@ =���<9�<'`�<���<e�<�m�<T��<�8�<��<��<�t�<6��<8>�<���<#��<�L�<��<���<�:�<چ�<���<��<�n�<��<��<vf�<1��<;�<'n�<���<�<s�<��<]�<�V�<ߖ�<l��<��<~1�<�Z�<J��<���<$��<���<	
�<%,�<�M�<8n�<���<Ϥ�<r��<h��<���<F��<ԗ�<5m�<�2�<���<D��<$'�<a��<J/�<���<�	�<�h�<��<��<WU�<C��<���<��<+2�<�X�<qw�<��<"��<R��<���<Ǒ�<�~�<#e�<OG�<�&�<I�<��<=Ơ<;��<��<1��<Br�<|f�<!]�<�T�<�K�<�@�<�2�< �<�	�<f�<�΃<0��<�	<��z<hv<�r<�m<�|i<26e<��`<��\<��X<QT<$#P<5�K<��G<��C<7l?<~4;<��6<��2<wb.<�*<�%<d!<�<��<K�<0H<�<�<	�<���;k�;�8�;�z�;^��;S�;�v�;p��;�0�;2��;���;�u�;G �;Ǥ�;.h�;1Q�;�d�;���;�5t;��g;~C[;�kO;��C;v�8;�M.;�#;��;�6;�;#��:��:���:�q�: ��:�>�:4��:�t�:�(n:d�R:��8:�z :A>	:�#�9���9�b�9V�S9��9#O8Π�D1޸,rB�#���gg��řṮt��u1�0�F��t[���o����拺\����3��u����.�������Pź�Ϻ�&ٺ�u������5�ڨ��V������~&���#�$�(�H�-��2��~7�%$<���@�?E���I�\oN��*S��X�u	]��/b��wg���l�qOr���w�N}�=d������Ɇ�)n��0	��ՙ��:"�������!��ҟ���  �  Ը=�h=@=��=�m=�=��=�_=�=�� =�H =,��<�%�<�u�<c��<�#�<��</��<sI�<^��<��</~�<��<�B�<
��<���<�I�<A��<���<�/�<6y�<���<��<�Z�<���< ��<cR�<i��<?�<]_�<���<��<&l�<���<��<�W�<R��<5��<�<L<�<�g�<!��<���<���<���<��<�A�<�b�<ہ�<���<���<���<'��<���<ݸ�<��<�m�<�0�<5��<��<�<���<��<��<9��<�S�<u��<4��<�@�<���<m��<���<�%�<O�<�p�<�<|��<I��<5��<���<��<Cp�<�T�<�6�<��<���<o۠<���<���<	��<���<Kx�<�l�<�a�<2V�<�H�<38�<�#�<p
�<|�<ʃ<棁<��~< �z<XIv<��q<q�m<�Si<Ze<a�`<��\<s^X<1T<+P<��K<v�G<.�C<�f?<4;<��6<C�2<%q.<�#*</�%<p�!<
4<�<j�<ht<�J<'.<9<M <�N�;2v�;��;���;�<�;o��;U��;'2�;㊺;��;�W�;�ף;bq�;F+�;�;J�;�W�;��s;T�f;��Z;��N;��C;�8;
.;a�#;��;-;�;��:g��:�V�:�#�:�k�:l@�: ��:���:��p:��U:��;:�"#:��:Z��9v��9Tʕ9�Y9�D9�S[85�ٷC�ܸ�C�Q���:
�����8�������3��H���]��r�UM���!�������7��p����Ⲻ-;��ЯźYQϺ!3ٺ	Y㺍�� ������^K����!~�������"��(�')-��2���6�2�;�_:@�B�D�s|I�`1N�l S�0�W�B]�Ab�8�g�m��r��3x�w�}�𩁻�g���������lZ��玻�h���ᓻ�U��Tɘ��  �  S�=�e=�=D�=�n=�=!�=�d=J	=j� =�Q =I��<�;�<���<c��<x:�<���<���<�Z�<7��<�#�<���<���<�F�<R��<X��<�E�<t��<���<O#�<�i�<��<���<zE�<'��<y��<r<�<���<z��<�N�<̬�<�	�<d�<���<4�<�W�<���<���<,�<;G�<�u�<@��<H��<f��<
�<q6�<�X�<�x�<���<Z��<���<`��<	��<���<#��<p��<�m�<�-�<l��<c�<��<G��<��<W|�<���<�<�<���<���<�)�<�m�<A��<-�<
�<D�<mh�<���<���<i��<���<R��<p��<�{�<c�<�G�<�*�<��<��<�מ<���<��<;��<���<�|�<o�<�`�<�P�<a=�<&�<H
�<��<dă<\��<��~<g�z<P'v<"�q<wm<�&i<Z�d<4�`<�f\<�6X<�T<��O<�K<��G<ۅC<�^?<�1;<��6<��2<l.<�7*<��%<~�!<GX<<��<�<	z<�\<�K<UF <{��;h��;���;I�;I[�;��;_��;�0�;`~�;KӲ;	5�;a��;�7�;y�;ÿ�;�Ɔ;6�;��r;�Af;�Z;XN;/C;�08;�-;g�#;��;�;��;U8�:*V�:1��:9��:L�:G�:�Ֆ:�:Ӛs:�yX:�>:}�%:K]:�v�9H��9�O�9�:_9��9��f8P�ͷ�ܸ25D������������V�	������5��~K�W�`�hSu�?����z������X��苪�Y����ټ�c!ƺ��Ϻ�Lٺ�H�����Zs����p����dq�M��k+"��^'�\r,�(g1�9A6�
;�C�?�pD��)I���M���R�h�W��	]�Zb���g��Zm���r�
�x�FP~�����z���-s�����W����;�������&�����������  �  e�=,b=V=m�=+o=�=Q�=Ri=E=ִ =�Z =�  =�P�<̢�<��<�P�<i��<�
�<�k�<s��<J/�<��<���<�I�<���<��<�@�<���<l��<��<"Z�<Ԟ�<���<r/�<G}�<|��<�%�<}��<1��<>�<U��<���<0[�<e��<��<�V�<���<.��<c�<=Q�<t��<��<_��<��<�(�<�L�<�n�<t��<Ū�<~��<���<L��<���<���<{��<��<il�<*�<���<�u�<U�<&��<��<Fh�<���<3%�<�y�<���<��<�W�<���<Ծ<X	�</8�<j_�<D~�<}��<���<ѥ�<��<���<�<qp�<�W�<4=�<@"�<��<r�<�֜<���<)��<��<���<�{�<�j�<�W�<�A�<�'�<(	�<��<ƽ�<���<B�~<�ez<\v<c�q<�Km<&�h<��d<�o`<<:\<�X<J�S<i�O<��K<�G<�vC<oU?<�-;<��6<��2<�.<J*<&<��!<�{<�;<\<��<��<��<Cw<Hn <���;'��;	�;dA�;Xv�;ݯ�;|��;�+�;n�;-��;��;�w�;���;���;4q�;�q�;�Q;�5r;��e;snY;N�M;c�B;8�7;�Z-;�J#;х;[;t�;�Z�:Ȥ�:�W�:�}�:Y�:�F�:���:+G�:�Sv:�N[:ArA:J�(:��:��9���9���9_nd9IL9F�p8�Fŷ�ݸ(�E��=�����ue� c���!�r>8�� N�zc��2x��#��9ݏ�"M��*��������������1�ƺ��Ϻ5uٺ�H㺙f�d����1���f�Jq�`��O4��{!�p�&�e�+�+�0���5��x:�D?��D��H���M�=�R��W�]��zb�,h�Ϧm��^s��y���~��E������͇��w��U����������m���͖�L+���  �  x�=�^=�=-�=1o==��=Am=�=p� =Yb =�	 =Cd�<#��<��<�d�<w��<@�<�z�<
��<99�<_��<��<�K�<��<
��<v;�<ق�< ��<	�<�J�<��<��<��<�g�<���<��<`l�<���<u-�<P��<f��< R�<��<��<NU�<���<���<s!�<�Y�<ˍ�<��<���<��<;<�<4a�<a��<0��<��<���<���<���<���<���<���<���<pj�<�%�<���<gl�<<��<�x�<���<�T�<���<��<�b�<���<}��<EC�<���<7þ<&��<~,�<AV�<�w�<I��<石<Ѧ�<���<U��<��<;|�<6f�<�M�<�4�<��<��<R�<՚<9��<���<���<���<s�<a]�<�D�<6(�<6�<`�<�<���<=�~<WHz<$�u<Iq<q"m<��h<��d<8D`<a\<��W<��S<��O<�K<WG<WgC<�J?<A(;<a�6<j�2<��.<�Y*<6&<6�!<b�<`<�)<��<5�<M�<�<�� <��;(�;k?�;9b�;@��;���;���;#�;�[�;��;M�;EG�;3��;�]�;�&�;H!�;��~;Ɍq;v�d;��X;�3M;�B;�V7;�-;�#;�U;��;��;�o�:!��:��:��:uٷ:]+�:��:�n�:7�x:��]:�D:C++:�>:V@�9#j�9/��9'�h9-�9&x8�\���i޸ڳG�:ʐ�O��36�����#�!�:���P�� f���z�[���,������?���ۈ���[�� 2��x$Ǻ�Gк��ٺ�U�fJ�p����� ��F�(�����Q�O���� ��&�'+� 0��5���9��>�1�C���H��M���R�n�W��&]�͟b�x;h�x�m���s���y�Ud�����lc���#���Ί��d���䏻�R��򲔻%	���\���  �  �=[=z=Ͽ=�n=�=��=Np=�=�� =�h =: =�t�<g��<�<�u�<���<�*�<C��<h��<RA�<��<q��<�L�<��<���<A6�<t{�<k��<���<�<�<�}�<���<<�<�T�<|��<���<�Z�<d��<��<ǃ�<���<�I�<ŧ�<o �<JS�<���<���< &�<�`�<)��<s��<H��<$�<�L�<sr�<���<��<{��<���<2��<��<���<Y��<���<{��<*h�<!�<L��<�c�<I��<�k�<���<D�<��<u��<�N�<ǝ�<��<1�<u�<j��<{�<�!�<�M�<yq�<��<읳<��<��<��<_��<<r�<�[�<�D�<,�<H�<���<��<nϘ<���<��<Ꮢ<�y�<�a�<�F�<#(�<��<�܅<v��<��<��~<Y.z<T�u<�]q<�l<��h<�\d<�`<u�[<}�W<��S<o�O<~K<_lG<�XC<�@?<<";<��6<J�2<}�.<�e*<�+&<*�!<Ե<a~<rK<�<�<��<J�<� <�S�;�T�;�b�;�{�;Ԝ�;I��; ��;S�;J�;f��;�Ī;��;%��;�"�;v�;_څ;�~;�p;�]d;�HX;h�L;�A;��6;��,;��";G(;��;�;'w�:
�:��:��:ns�:8�:�:!h�:��z:M`:'5F:�J-:.4:k��9_�9���9Πl9��9�?}8�ʾ��'�ئI�&A���W��������%���<���R�pth��P}����LT���������\g������ξ�͞Ǻi�кv�ٺ\j㺐<�R��!� �U�,N���#���R ��y%���*���/�К4���9�i>�
pC��iH�sM���R��W��:]���b��ph�~:n��t���y�T��Ԃ�����o�����&���`-��$���A;>��9����  �  A�=5X=o=��=zn=5= �=|r=�=�� =�m =� =ʀ�<O��<.+�<���<���<�5�<���<��<'G�<��<���<M�<ѝ�<��<�1�<du�<õ�<2��<%2�<�q�<���<��<�E�<���<���<�L�<���<��<�y�<���<�B�<���<���<ZQ�<R��<<��<*)�<�e�<
��<
��<��<�/�<LY�<g�<���<W��<���<���<���<���<���<v��<"��<��<f�<M�<���<\�<���<a�<���<�6�<���<w��<:?�<U��<2��<�"�<h�<Ȩ�<H�<\�<�F�<,l�<���<���<���<���<x��<���<��<{�<�f�<IP�<9�<U!�<�	�<��<�ژ<Ė<f��<���<w~�<�d�<H�<�'�<��<<م<��<�x�<;�~<�z<��u<�Cq<��l<^�h<�>d<B `<��[<��W<ˎS<�zO<�kK</]G<�LC<�7?<�;<��6<��2<��.<�n*<08&<z "<��<C�<^d<w8<<;�<?�<�� <�{�;�u�;�|�;
��;I��;��;~��;c�;o:�;ik�;t��;���; d�;W��;ذ�;���;3�};�p;2�c;��W;-TL;;FA;�6;�r,;��";� ;ϯ;I�;�t�:�$�:�A�:"��:��:�s�:d��:�"�:e|:�a:X�G:'�.:��:�_�9ו�9-ȣ9�8o9$�9�N�8I������*UK���������������b*'�>�ɊT�n>j��*�����7��2t���^��������#L���Ⱥ��к�ں���Q:�1��ϰ �f��+�5N������]���%�**��9/�@4��?9�}=>�:<C�AEH��\M��R���W�M]���b��h��sn��\t��Nz�I����yㅻ)����V��uꍻ�e���ʒ�r��Fh��묙��  �  �=RV==��=n=`=��=�s=�=U� =�p =O =~��<z��<�3�<���<��<p<�<n��<���<�J�<W��<���<6M�<ٜ�<��<�.�<hq�<��<E��<J+�<�i�<��<���<l<�<3��<5��<D�<{��<=�<ds�<6��<�>�<��<x��<�O�<���<���<	+�<�h�<��<I��<��<�6�<a�<���<թ�<3��<?��<1��<��<���<���<M��<���<{��<pd�<��<��<�W�<���<rZ�<P��<W.�<���<���<T5�<h��<���<��<�_�<_��<�ݼ<��<uB�<�h�<��<���<]��<h��<~��<���<d��<���<m�<�W�<A�<�)�<��<���<��<7ʖ<���<|��<j��<uf�<�H�<)'�<E�<�օ<r��<Dt�<(|~<�z<ԝu<3q<�l<Nwh<q+d<�_<��[<��W<"S<:mO<�_K<�SG<EC<.2?<;<�6<�2<`�.<�s*<�?&<b
"<��<q�<$t<<I<P#<�	<�<� <��;���;��;H��;���;��;'��;�	�;�/�;�\�;t��;X�;�I�;"֓;)��;���;�[};�;p;��c;g�W;�L;�A;�x6;J,;�r";��;�;
�;Kr�:�1�:b�:��:C'�:Tɩ:@�:���:%}}:�b:,�H:A�/:}�:���9���9P֤9��p9f�9K�8c��D8�V{L�-[���ù}�l��U(�8!?���U�!hk��,���3��7ʓ�����Pޥ�5���\��{����CȺHѺ*3ں#���9� ���� ����H�
�!��S���)����$�W�)���.��4��9�Q>��C��.H��OM���R�W�W�}Z]���b�M�h�ޗn�k�t��z��:��Y)������Έ��|��K��L���6쒻=��Â���Ù��  �  �=�U=�
=]�=n=r=�=It=~=;� =�q =w =��<��<E6�<V��<���<�>�<r��<e��<�K�<$��<.��<OM�<���<U��<�-�<�o�<��<,��<�(�<�f�<2��<���<S9�<5��<��<A�<���<�	�<<q�<9��<�<�<��<���<WO�<��<��<�+�<�i�<���</��<�
�</9�<�c�<K��<}��<���<���<J��< ��<l �<���<���<���<d��<�c�<��<��<?V�<���<0X�<���<q+�<���<e��</2�<4��<O��<��<�\�<ើ<�ۼ<��<�@�<�g�<<��<	��<R��<���<&��<ٟ�<�<y��<7o�<Z�<�C�<V,�<m�<W��<Q�<U̖<h��<ߛ�<i��<�f�<�H�<
'�<� �<�Յ<1��<�r�<x~<2z<��u<^-q<�l<�ph<n%d<��_<~�[<ɒW<�yS<�hO<�[K<PG<;BC<:0?<�;<��6<T�2<*�.<�u*<MB&<"<	�<*�<Uy<�N<�(<S	<6�<�� <w��;��;���;��;M��;��;K��;��;�,�;�W�;���;lڢ;A�;�˓;"��;�t�;�C};�$p;��c;��W;�K;>�@;�g6;�:,;=f";U�;�;#�;-r�:@5�:l�:��:�>�:]�:v�:J��:k�}:�c:=;I:q/0:U�:^B :m�9K6�9�^q9��9H�8/k��4��&�L������pùǚ����_(��y?���U�X�k��\���d��b���++���	������3��$���o[Ⱥ�*Ѻ�>ں����8�k���� �
��D�
��/B�Lo����W�$�D�)�N�.��3���8�|>��C�'H�BLM�P�R���W�j_]� c���h�S�n�ϙt���z��D���4������ۈ��������~��������G��ǋ��̙��  �  �=RV==��=n=`=��=�s=�=U� =�p =O =~��<z��<�3�<���<��<p<�<n��<���<�J�<W��<���<6M�<ٜ�<��<�.�<hq�<��<E��<J+�<�i�<��<���<l<�<3��<5��<D�<{��<=�<ds�<6��<�>�<��<x��<�O�<���<���<	+�<�h�<��<I��<��<�6�<a�<���<թ�<3��<?��<1��<��<���<���<M��<���<{��<pd�<��<��<�W�<���<rZ�<P��<W.�<���<���<T5�<h��<���<��<�_�<_��<�ݼ<��<uB�<�h�<��<���<^��<i��<~��<���<d��<���<m�<�W�<A�<�)�<��<���<��<7ʖ<���<{��<j��<tf�<�H�<('�<E�<�օ<r��<Dt�<'|~<�z<ԝu<3q<�l<Nwh<q+d<�_<��[<��W<"S<:mO<�_K<�SG<EC<.2?<;<�6<�2<a�.<�s*<�?&<b
"<��<r�<%t<=I<P#<�	<�<� <��;���;��;G��;���;��;%��;�	�;�/�;�\�;s��;W�;�I�;!֓;(��;���;�[};�;p;��c;f�W;�L;�A;�x6;J,;�r";��;�;
�;Jr�:�1�:b�:��:C'�:Tɩ:@�:���:%}}:�b:,�H:A�/:}�:���9���9P֤9��p9f�9K�8c��D8�V{L�-[���ù}�l��U(�8!?���U�!hk��,���3��7ʓ�����Pޥ�5���\��{����CȺHѺ*3ں#���9� ���� ����H�
�!��S���)����$�W�)���.��4��9�Q>��C��.H��OM���R�W�W�}Z]���b�M�h�ޗn�k�t��z��:��Y)������Έ��|��K��L���6쒻=��Â���Ù��  �  A�=5X=o=��=zn=5= �=|r=�=�� =�m =� =ʀ�<O��<.+�<���<���<�5�<���<��<'G�<��<���<M�<ѝ�<��<�1�<du�<õ�<2��<%2�<�q�<���<��<�E�<���<���<�L�<���<��<�y�<���<�B�<���<���<ZQ�<R��<<��<*)�<�e�<
��<
��<��<�/�<LY�<g�<���<W��<���<���<���<���<���<v��<"��<��<f�<M�<���<\�<���<a�<���<�6�<���<x��<;?�<U��<3��<�"�<h�<Ȩ�<H�<\�<�F�<,l�<���<���<���<���<y��<���<��<{�<�f�<JP�<9�<U!�<�	�<��<�ژ<Ė<f��<���<w~�<�d�<H�<�'�<��<<م<��<�x�<:�~<�z<��u<�Cq<��l<^�h<�>d<B `<��[<��W<̎S<�zO<�kK<0]G<�LC<�7?<�;<��6<��2<��.<�n*<08&<{ "<��<C�<^d<w8<<;�<?�<�� <{�;�u�;�|�;��;G��;��;{��;a�;m:�;gk�;q��;���;�c�;U��;ְ�;���;0�};�p;/�c;��W;+TL;:FA;�6;�r,;��";� ;ί;H�;�t�:�$�:�A�:"��:��:�s�:d��:�"�:e|:�a:X�G:&�.:��:�_�9ו�9-ȣ9�8o9$�9�N�8I������*UK���������������b*'�>�ɊT�n>j��*�����7��2t���^��������#L���Ⱥ��к�ں���Q:�1��ϰ �f��+�5N������]���%�**��9/�@4��?9�}=>�:<C�AEH��\M��R���W�M]���b��h��sn��\t��Nz�I����yㅻ)����V��uꍻ�e���ʒ�r��Fh��묙��  �  �=[=z=Ͽ=�n=�=��=Np=�=�� =�h =: =�t�<g��<�<�u�<���<�*�<C��<h��<RA�<��<q��<�L�<��<���<A6�<t{�<k��<���<�<�<�}�<���<<�<�T�<|��<���<�Z�<d��<��<ǃ�<���<�I�<ŧ�<o �<JS�<���<���< &�<�`�<)��<s��<H��<$�<�L�<sr�<���<��<{��<���<2��<��<���<Y��<���<{��<*h�<!�<L��<�c�<J��<�k�<���<D�<��<v��<�N�<ȝ�<��<1�<u�<k��<|�<�!�<�M�<zq�<��<읳<��<��<��<`��<<r�<�[�<�D�<,�<H�<���<��<nϘ<���<��<���<�y�<�a�<�F�<"(�<��<�܅<u��<��<��~<W.z<S�u<�]q<�l<��h<�\d<�`<u�[<}�W<��S<p�O<~K<`lG<�XC<�@?<=";<��6<K�2<~�.<�e*<�+&<+�!<յ<a~<sK<�<�<��<J�<� <�S�;�T�;�b�;�{�;ќ�;F��;���;O�;J�;b��;�Ī;��;"��;�"�;t�;\څ;�~;�p;�]d;�HX;e�L;�A;��6;��,;��";F(;��;~�;&w�:
�:��:��:ms�:8�:�:!h�:��z:M`:'5F:�J-:.4:k��9_�9���9Πl9��9�?}8�ʾ��'�ئI�&A���W��������%���<���R�pth��P}����LT���������\g������ξ�͞Ǻi�кv�ٺ\j㺐<�R��!� �U�,N���#���R ��y%���*���/�К4���9�i>�
pC��iH�sM���R��W��:]���b��ph�~:n��t���y�T��Ԃ�����o�����&���`-��$���A;>��9����  �  x�=�^=�=-�=1o==��=Am=�=p� =Yb =�	 =Cd�<#��<��<�d�<w��<@�<�z�<
��<99�<_��<��<�K�<��<
��<v;�<ق�< ��<	�<�J�<��<��<��<�g�<���<��<`l�<���<u-�<P��<f��< R�<��<��<NU�<���<���<s!�<�Y�<ˍ�<��<���<��<;<�<4a�<a��<0��<��<���<���<���<���<���<���<���<pj�<�%�<���<gl�<<��<�x�<���<�T�<���<��<�b�<���<~��<FC�<���<8þ<'��<,�<BV�<�w�<J��<蟳<Ҧ�<���<U��<��<<|�<7f�<�M�<�4�<��<��<R�<՚<8��<���<���<���<s�<`]�<�D�<5(�<5�<_�<�<���<;�~<VHz<#�u<Hq<q"m<��h<��d<8D`<b\<��W<��S<��O<�K<YG<YgC<�J?<C(;<c�6<l�2<�.<�Y*<7&<8�!<c�<`<�)<��<5�<M�<�<�� <��;(�;h?�;6b�;<��;���;���;#�;�[�;���;I�;AG�;/��;�]�;~&�;F!�;��~;Ōq;r�d;��X;�3M;�B;�V7;�-;�#;�U;��;��;�o�: ��:��:��:uٷ:]+�:��:�n�:7�x:��]:�D:C++:�>:V@�9#j�9/��9&�h9-�9&x8�\���i޸ڳG�:ʐ�O��36�����#�!�:���P�� f���z�[���,������?���ۈ���[�� 2��x$Ǻ�Gк��ٺ�U�fJ�p����� ��F�(�����Q�O���� ��&�'+� 0��5���9��>�1�C���H��M���R�n�W��&]�͟b�x;h�x�m���s���y�Ud�����lc���#���Ί��d���䏻�R��򲔻%	���\���  �  e�=,b=V=m�=+o=�=Q�=Ri=E=ִ =�Z =�  =�P�<̢�<��<�P�<i��<�
�<�k�<s��<J/�<��<���<�I�<���<��<�@�<���<l��<��<"Z�<Ԟ�<���<r/�<G}�<|��<�%�<}��<1��<>�<U��<���<0[�<e��<��<�V�<���<.��<c�<=Q�<t��<��<_��<��<�(�<�L�<�n�<t��<Ū�<~��<���<L��<���<���<{��<��<il�<*�<���<�u�<U�<&��<��<Fh�<���<4%�<�y�<���<��<�W�<���<Ծ<Y	�<08�<k_�<E~�<~��<���<ҥ�<��<���<���<rp�<�W�<5=�<@"�<��<r�<�֜<���<(��<~��<���<�{�<�j�<�W�<�A�<�'�<'	�<��<Ž�<���<@�~<~ez<[v<c�q<�Km<&�h<��d<�o`<<:\<�X<K�S<j�O<��K<�G<�vC<qU?<�-;<��6<��2<�.<J*<&<��!<�{<�;<]<��<��<��<Bw<Gn <���;$��;�;`A�;Tv�;ٯ�;x��;�+�;n�;(��;��;�w�;���;���;0q�;�q�;�Q;�5r;��e;pnY;J�M;a�B;5�7;�Z-;�J#;υ;Z;s�;�Z�:Ǥ�:�W�:�}�:Y�:�F�:���:+G�:�Sv:�N[:ArA:J�(:��:��9���9���9_nd9IL9F�p8�Fŷ�ݸ(�E��=�����ue� c���!�r>8�� N�zc��2x��#��9ݏ�"M��*��������������1�ƺ��Ϻ5uٺ�H㺙f�d����1���f�Jq�`��O4��{!�p�&�e�+�+�0���5��x:�D?��D��H���M�=�R��W�]��zb�,h�Ϧm��^s��y���~��E������͇��w��U����������m���͖�L+���  �  S�=�e=�=D�=�n=�=!�=�d=J	=j� =�Q =I��<�;�<���<c��<x:�<���<���<�Z�<7��<�#�<���<���<�F�<R��<X��<�E�<t��<���<O#�<�i�<��<���<zE�<'��<y��<r<�<���<z��<�N�<̬�<�	�<d�<���<4�<�W�<���<���<,�<;G�<�u�<@��<H��<f��<
�<q6�<�X�<�x�<���<Z��<���<`��<	��<���<#��<p��<�m�<�-�<l��<c�<��<H��<��<W|�<���<�<�<���<���<�)�<�m�<B��<.�<�<D�<nh�<���<���<j��<���<S��<q��<�{�<c�<�G�<�*�<��<��<�מ<���<��<;��<���<�|�<o�<�`�<�P�<`=�<&�<G
�<��<că<[��<��~<f�z<N'v<!�q<wm<�&i<Z�d<4�`<�f\<�6X<�T<��O<�K<��G<݅C<�^?<�1;<��6<��2<n.<�7*<�%<��!<HX<<��<�<	z<�\<�K<TF <x��;e��;���;E�;E[�;��;Z��;�0�;\~�;FӲ;5�;\��;�7�;u�;���;�Ɔ;3�;}�r;�Af;�Z;XN;,C;�08;�-;e�#;��;�;��;T8�:)V�:0��:8��:L�:G�:�Ֆ:�:Ӛs:�yX:�>:}�%:K]:�v�9H��9�O�9�:_9��9��f8P�ͷ�ܸ25D������������V�	������5��~K�W�`�hSu�?����z������X��苪�Y����ټ�c!ƺ��Ϻ�Lٺ�H�����Zs����p����dq�M��k+"��^'�\r,�(g1�9A6�
;�C�?�pD��)I���M���R�h�W��	]�Zb���g��Zm���r�
�x�FP~�����z���-s�����W����;�������&�����������  �  Ը=�h=@=��=�m=�=��=�_=�=�� =�H =,��<�%�<�u�<c��<�#�<��</��<sI�<^��<��</~�<��<�B�<
��<���<�I�<A��<���<�/�<6y�<���<��<�Z�<���< ��<cR�<i��<?�<]_�<���<��<&l�<���<��<�W�<R��<5��<�<L<�<�g�<!��<���<���<���<��<�A�<�b�<ہ�<���<���<���<'��<���<ݸ�<��<�m�<�0�<5��<��<�<���<��<��<:��<�S�<v��<5��<�@�<���<n��<���<�%�<O�<�p�<���<}��<J��<6��<���<��<Cp�<�T�<�6�<��<���<o۠<���<���<	��<���<Jx�<�l�<�a�<2V�<�H�<28�<�#�<o
�<{�<ʃ<壁<��~<�z<WIv<��q<p�m<�Si<Ze<a�`<��\<t^X<1T<,P<��K<x�G<0�C<�f?<4;<��6<E�2<'q.<�#*<0�%<r�!<4<�<j�<it<�J<&.<8<L <�N�;/v�;��;���;�<�;k��;Q��;#2�;ފ�;��;�W�;�ף;^q�;B+�;�;G�;�W�;��s;O�f;�Z;��N;��C;�8;.;_�#;��;-;�;��:f��:�V�:�#�:�k�:k@�: ��:���:��p:��U:��;:�"#:��:Z��9v��9Tʕ9�Y9�D9�S[85�ٷC�ܸ�C�Q���:
�����8�������3��H���]��r�UM���!�������7��p����Ⲻ-;��ЯźYQϺ!3ٺ	Y㺍�� ������^K����!~�������"��(�')-��2���6�2�;�_:@�B�D�s|I�`1N�l S�0�W�B]�Ab�8�g�m��r��3x�w�}�𩁻�g���������lZ��玻�h���ᓻ�U��Tɘ��  �  ��=Wk=u=��=�l=)=ŷ=�Z=�� =6� =3@ =���<9�<'`�<���<e�<�m�<T��<�8�<��<��<�t�<6��<8>�<���<#��<�L�<��<���<�:�<چ�<���<��<�n�<��<��<vf�<1��<;�<'n�<���<�<s�<��<]�<�V�<ߖ�<l��<��<~1�<�Z�<J��<���<$��<���<	
�<%,�<�M�<8n�<���<Ϥ�<r��<h��<���<F��<ԗ�<5m�<�2�<���<D��<$'�<b��<J/�<���<�	�<�h�<��<��<WU�<D��<���<��<,2�<�X�<rw�<��<#��<S��<���<ȑ�<�~�<$e�<OG�<�&�<J�<��<=Ơ<;��<��<1��<Ar�<{f�< ]�<�T�<�K�<�@�<�2�<~ �<�	�<e�<�΃<0��<�	<��z<hv<�r<�m<�|i<26e<��`<��\<��X<QT<%#P<6�K<��G<��C<9l?<�4;<��6<��2<xb.<�*<�%<d!<�<��<L�<0H<�<�<	�<���;i�;�8�;�z�;[��;O�;�v�;l��;�0�;.��;���;�u�;C �;ä�;+h�;-Q�;�d�;���;�5t;}�g;zC[;�kO;��C;t�8;�M.;�#;��;�6;�;"��:��:���:�q�:���:�>�:4��:�t�:�(n:c�R:��8:�z :@>	:�#�9���9�b�9V�S9��9#O8Ϡ�D1޸,rB�#���gg��řṮt��u1�0�F��t[���o����拺\����3��u����.�������Pź�Ϻ�&ٺ�u������5�ڨ��V������~&���#�$�(�H�-��2��~7�%$<���@�?E���I�\oN��*S��X�u	]��/b��wg���l�qOr���w�N}�=d������Ɇ�)n��0	��ՙ��:"�������!��ҟ���  �  ��=3m=2=?�=k=�=C�=V=� =�� =�8 =��<��<:M�<_��<���<�[�<���<�)�<��< �<�k�<���<�9�<���<���<�N�<��<b��<�C�<��<D��</�<�<T��<#�<}w�<��<r#�<Kz�<���<�%�<4x�<��<�<gU�<W��<���<��<�'�<�N�<Ur�<	��<ʴ�<���<��<&�<Y;�<�\�<�{�<ٖ�<���<���<���<��<���<l�<�3�<��<ݔ�<</�<��<�;�<s��<Z�<pz�<V��<  �<�f�<���<5��<2�<U<�<P`�<�|�<��<霵<柳<��<"��<�v�<[�<;�<v�<A��<Ӣ<���<��<��<�n�<a�<�V�<TO�<�H�<�A�<'9�<9-�<)�<��<n�<�у<ð�<�<~�z<Q�v<04r<��m<j�i<lYe<�a<1�\<͠X<�kT<[9P<�L<k�G<�C<�o?<�3;<��6<�2<�T.<��)<��%<I!<��<��<)[<p!<p�<(�<��<%��;`��;3�;ML�;)��; �;�a�;���;�,�;��;��;��;�!�;�Μ;���;[��;��;��;)�t;
h;��[;��O;�[D;�B9;`�.;�!$;';]9;�;"��:�8�:tK�:���:�г:}[�:���:�[�:��k:�vP:��6:�%:�	:R#�9�	�9�V�9|�N9n��8�C8t���D�߸�3B�u㊹�+����߹V<�h����/���D�;VY�W�m�1���hڊ�~����Z��g���h���D��[	ź��κ7&ٺ���6S�S��]I�_����qx�~$�]��U $��^)�n.�xO3�\8��<��!A��E�mJ���N��SS�/ X��]��%b��[g���l��r�zw��|��)��dڃ������(��;ċ��X��琻8p�������}���  �  ��=xn=�=��=�i=�=\�=lR=~� =:� =�2 =��<���<�>�<���< ��<�M�<��<%�<���<Z��<�d�<;��<�5�<h��<K��<�O�< ��<��<UJ�<f��<U��<�:�<f��<Q��<30�<*��<���<-.�<i��<!��<G+�<�{�<��<-�<�S�<C��<%��<���<��<#E�<[g�<�<K��<k��<e��<r
�</-�<JO�<�o�<��<���<���<ǲ�<F��<���<�j�<>4�<D��<���<5�<���<�E�<���<�&�<���<��<�-�<t�<���<%��<i�<�C�<�e�<p��<��<���<l��<���<F��<p�<�R�<@1�<L�<��<hŢ<Y��<N��<mr�<�`�<�S�<�J�<oD�<�?�<%:�<�2�<�(�<;�<R�<��<$ԃ<���<�%<�z<i�v<bJr<� n<V�i<�se<�1a<��\<��X<�T<�IP<�L<��G<��C<�q?<62;<��6<��2</I.<��)<h�%<�3!<��<Ć<j><�<��<I�<�<Rq�;Ҙ�;���;Q'�;���;���;�O�;���;�'�;��;-�;t��;�9�;"�;:��;���;�Ӈ;��;H!u;�kh;�\;{+P;��D;�z9;��.;�<$;Z;_7;��;�U�:x��:��:�M�:E4�:먢:l��:䀃:�
j:ΛN:�4:�Z:�R:��9�=�9�ߌ9x�J9�M�8�98�~�J���EB��r��IL���o޹�U�m��b.��/C���W� l������yڶ���s��w-��t�����ĺ]�κ�-ٺط�J�� ���)��'A�6�������1$���$���)�`�.���3�r8�C�<��wA���E��VJ�P�N��vS�6X��]�a"b�Ig�j�l��q��;w��|�����G����Q��K􈻶���5(��t���cI���֕�-e���  �  �=(o=�=_�=�h=5=r�=P=�� =� =�. ={��<���<'5�<��<���<�D�<���<��<?��<���<q`�<���<W3�<ǖ�<���<P�<���<���<9N�<{��<o��<�A�<1��<���<�8�<+��<R��<�4�<��<���<�.�<#~�< ��<'�<�R�<��<���<���<��<?�<W`�<��<���<E��<���<	�<�#�<�F�<�g�<ׄ�<��<ê�<���<1��<���<�i�<_4�<h��<H��<�8�<T��<\K�<���<�.�<��<���<n6�<\|�<`��<���< �<:H�<7i�<���<���<���<?��<ϔ�<��<�k�<�M�<+�<�<��<���<��<��<�h�<�W�<"K�<�B�<�=�<�9�<;5�<�.�<�%�<+�<M�<��<LՃ<-��<�,<\�z<
�v<Xr<>n<��i<�e<{Ba<�]<��X<��T<�SP<�L<#�G<ήC<|r?<�0;<Q�6<��2<�A.<o�)<օ%<2&!<M�<�u<,<+�<��<�<��<�N�;gy�;W��;��;p�;���;
D�;���;2$�;���;j�;���;�G�;&�;\ؕ;Ҏ;��;R;�;�au;��h;jR\;^P;\�D;)�9; �.;�L$;x;�5;k�;�0�:|��: ��:���:�Ѳ:�6�:�<�:���:w�h:�jM:s�3:)1:`=:��9>r�9�T�9�CH9��8�38���⸣XB��<���Ƴ��ݹ���-����-��CB��V�k��6�����t|��8S��� ��{��ƺ��ĺ��κ4ٺ�㺳��8���Y��Nl�@�����4j���$�!*�C//�	4���8��==��A��F�Q}J���N�*�S��EX�!]�� b�/?g�wwl���q�aw��n|��※ڋ��V1���҈�$p���	��۞���1���Õ��V���  �  ��=Tz=%=J�=�r=B=ߴ=/R=�� =i� =�% =���<���<z�<�i�<O��<'.�<���<��<��<��<�y�<3��<�]�<i��<X+�<ω�<���<G:�<Ύ�<���<G6�<P��<%��<�4�<ۊ�<���<A9�<���<$��<�@�<��<���<;�<��<��<��<�;�<�h�<��<��<1��<B��<W
�<�*�<&O�<hw�<��<���<���<.*�<�O�<�l�<�}�<���<�s�<U�<�$�<���</��<�-�<���<>�<���<��<Jy�<R��<l�<ZU�<Ì�<n��< �<@�<� �<G3�<�=�<�>�<�5�<*#�<��<�<e��<̂�<�N�<5�<��<h��<]��<�<"k�<�^�<hX�<�V�<�V�<�V�<T�<mM�<6A�<J/�<��<k��<-ف<ti<�{<�v<!~r<�.n<��i<��e<Ga<I�\<�X<VuT<M5P<��K<P�G<HyC<�4?<,�:<!�6<�12<��-<S)<��$<a_ <K�<9z<<4�<��
<�m<*`< ��;x��;$I�;���;��;�}�;���;P�;���;��;���;<��;�|�;��;Cܒ;���;�Ȅ;�{;�n;/�a;pU;bI;��=;*�2;Z�';�9;&;n5	;��:8�:���:3w�:)��:K�:}��:�e�:�*h:�JK:�N0:�=:� :W��9A̬9��9�E9��8$]]8�̀�`n���M$�}oq�J��_�ȹ�M��b�!�9�5��J��^���q�xЂ�����)Q�����g����<��鼺d�ƺڶкۺ���˫������+�	�$����F����!��9'��~,��|1��06���:���>��C�L!G��<K�tpO�b�S�FRX��
]���a�Mg�B2l�vvq���v��|�+���8V������Q���q/��Lō�qX���璻�u�����  �  i�=z=%=��=Is=�=׵=WS=_� =�� =h' =���<���<��<n�<���<E2�<a��<s�<���<��<�{�<
��<"_�<s��<�+�<���<��<=9�<I��<j��<�3�<7��<���<1�<8��<6��<�5�< ��<���<�>�<���<��<�:�<��<���<�<_=�<�j�<���<ҳ�<z��<���<[�<9/�<�S�<�{�<_��<���<��<{-�<�R�<Ao�<��<���<�t�<�U�<�$�<���<S��<W,�<���<v;�<���<;�<�u�<���<��<�Q�<j��<r��<l�<t�<W�<�2�<c=�<�>�<�6�<d$�<5�<&�<���<�<>R�<��<��<�à<���<o��<io�<�b�<#\�<�Y�<�Y�<Y�<V�<O�<sB�< 0�<��<��<K؁<�f<�{<��v<%xr<(n<��i<9�e<�?a<X�\<˱X<�oT<�0P<��K<@�G<HxC<�4?<5�:<G�6<�42<��-<�W)<c�$<�e <��<?�<�"<4�<~�
<�v<�h<6��;D�;V�;��;`�;���;2��;�T�;(��;L�;��;��;Zw�;	�;�ђ;Ȳ�;���;U�{;�n;�a;�VU;LI;B�=;-x2;G�';J4;�;P7	;-�:xM�:���:]��:�ε:�z�:Ϸ�:ա�:��h:��K:��0:��:n� :��9���9���93�F9��8��a8q4t�"��j�#��Rq��U��>�ȹ��{S���!�O76�pJ��}^��^r�
���ό������'������FV��������ƺl�к�ںɖ���,���/����	�����������!��'�`\,��Y1��6���:�a�>���B��
G��)K��`O�+�S��HX��]���a�Dg��9l�2�q�f�v��)|�����c��
��룈��=���ҍ��d��{�[~���
���  �  ��=�y=&%=Z�=�t=�=��=�V=^� =�� =�, =��<��<�&�<{�<���<S>�<���<��<��<U�<H��<��<�b�<���<-�<���<���<�5�<t��<���<�+�<�}�<V��< &�<2|�<���<,�<���<k��<&9�<���<���<:�<���<���<C�<�A�<�p�<��<1��<��<���<�<�;�<j`�<���<ݳ�<���<V�<7�<[�<Dv�<���<��<�w�<�W�<b%�<���<ƌ�<(�<Ǵ�<�3�<æ�<��<j�<���<"�<�F�<_�<Ȱ�<)ۿ<���<Y�<E0�<�<�<�?�<�8�<�'�<��<��<+��<H��<\�<�)�<���<qР<���<e��<�{�<Gn�<�f�<Kc�<�a�<�_�<�[�<SS�<�E�<�1�< �<7��<�Ձ<M^<�{<ιv<Rfr<�n<�i<�te<�)a<��\<U�X<`T<
$P<��K<�G<uC<�4?<��:<��6<p<2<�-<�d)<o�$<=x <�<}�<�;<��<&�
<�<��<��;�6�;�{�;���;�5�;ƛ�; �;a�;���;��;�{�;O�;�e�;���;���;��;ϓ�;N�{;�Nn;�wa;4
U;
I;Dv=;�M2;Ί';�#;�;>	;GP�:N��:��:��:�A�:�:�S�:�P�:�%j:�hM:�|2:mj:�#:���9!{�9�0�9��J9��9njm8hO�]���J�"���p��v���Gɹ~��� ���"�xD7��K�|�_��s�Ҹ��w����.����*�������1����ƺ3�кG�ںLp�i\��������	�n�����Mq�)-!���&�}�+���0�L�5�x*:��w>�\�B���F���J��4O��S�"1X��\���a�g�UOl���q�
w��e|�}ျ����0��Ј��h�������������얕�����  �  z�=9x=%=Q�=�v==��=�[=~� =Ė =�4 =$��<_��<�:�<^��<e��<jQ�<Q��<u.�<Т�<�<���<���<sh�<���<�.�<ӈ�<j��<l0�<B��<4��<��<�n�<���<��<�j�<���<@�<�w�<���<�/�<��<���<18�<3��<n��<��<�H�<wy�<ԣ�<��<��<��<{,�<#O�<�t�<���<\��<.��<7�<F�<�g�<��<O��<v��<c|�<Z�<�%�<w��<=��< !�<���<�'�<"��<s��<�X�<}��<���<5�<(o�<���<SϿ<���<��<,�<�:�<@�<Y;�<I,�<��<��<<ɫ<���<Rk�<-;�<l�<�<���<z��<8��<���<pw�<r�<�n�<�j�<\d�<�Y�<J�<94�<U�< ��<с<�O<@�z</�v<,Ir<�m<<�i<Qe<�a<S�\<5�X<+FT<�P<��K<C�G<�oC<Q3?<4�:<(�6<;H2<�-<y)<%<=� <�%<,�<�b<�<��
<��<�<~U�;y�;j��;��;y_�;���;��;Qr�;�ƿ;��;&r�;Ԩ;�G�;�ԙ;���;6U�; T�;�{;��m;?�`;?�T;�H;�=;I2; Y';C;�;EE	;��:���:��:Y��:-�:�ե:iF�:$a�:{l:��O:�5:��:U�:���9�ô9f��9�oQ9�{9�q8[���ب��^!�ƍp��ݠ�y?ʹ�%��#"��#$�,�8�{�M���a�t�u�qЄ�f������D~���٪�{.������oǺ]�к�ںl;庁��0��aY�R7	�%���p��g� �4&�LR+�=Q0�H5���9�A�=��2B��eF���J�3�N��iS�MX���\��a�2!g��tl���q��Rw���|�o���̃��u�����歋��<��]Ð�/C��r����:���  �  ��=%v=x$=(�=�x=�=]�=�a==ɟ =? =��<�<�T�<���<�<�i�<���<�B�<A��<�&�<ӗ�<��<�n�<E��<�/�<��<���<�(�<u�<���<��<�Z�<���<p��<%S�<ɫ�<7�<�d�<���< #�<���<z��<5�<��<���<!�<XP�<��<*��<3��<���<� �<D�<:h�<h��<���<~��<�
�<�3�<�X�<x�<H��<���<��<T��<4\�<%�<���<���<�<���<�<���<���<�@�<��<;��<��<�Y�<���<\��<��<U�<�%�<�7�<�?�<�=�<�1�<|�<���<�֫< ��<�~�<�P�<`%�<w��<�ڞ<d��<4��<���<���<���<a~�<�w�<�n�<�a�<O�<�6�<��<j�<wʁ<�;<|�z<�v<k"r<��m<�qi<w!e<��`<�\<2YX<e#T<p�O<��K<�G<GfC<C0?<��:<5�6<�U2<�-<�)<k&%<�� <|O<��<F�<YL<�<��<��<ܲ�;;��;* �;7D�;���;���;U7�;P��;JϿ;a�;�b�;5��;c�;@��;V?�;X�;���;�Pz;1m;D`;��S;�H;Ţ<;Ħ1;�';��; �;VH	;��:�.�:��:7�:η:>ܦ:
y�:���:6uo:�	S:_K8:!;:��:���9!0�9�ђ9��Y9V9ީ�8�p���J�����sp����|�˹f����&�]L;�6P�V�d���x��E��f揺�T�������ƫ�贺����cǺ��кY�ںW庸�ﺃ������C�����^q�4�����E%�Ӏ*� �/�$J4�f�8� M=��A���E��:J���N�~/S� �W��\�$�a��?g�4�l�%/r�<�w�NL}�|h���"���ц�t��^
������}������~����d���  �  �=4s=3#=w�=�z=�!=i�=�h=t	=ѩ =�J =��<0#�<r�<[��<A#�<w��<3��<#Y�<���<�6�<���<�<u�<Z��<}/�<փ�<���<�<�f�<��<���<�B�<]��<���<h7�<Ґ�<���<;N�<y��<��<�u�<��<V0�<���<���<��<AX�<)��<���<��<�<9�<�^�<���<��<2��<��<}%�<�K�<5n�<��<���<ģ�<Ü�<ԅ�<s]�<#�<���<�x�<]
�<Q��<��<%m�<G��<�$�<�t�<3��<��<�?�<�x�<꫿<ٽ<5��<��<�2�<P>�<�?�<q6�<�#�<2�<��<m��<l��<�i�<~@�<\�<���<�ۜ<�Ě<c��<w��<��<叒<텐<�y�<-i�<�S�<�7�<��<1�<u��<]"<��z<�Wv<��q<��m<�:i<0�d<.�`<3`\<)X<m�S<��O<ݨK<��G<gYC<3*?<0�:<�6<�b2<�.<��)<H%<$� <�~<�!<��<��<�Q<+<�<��;,�;R�;���;���;�;�T�;`��;~ӿ;��;UL�;���;r�;�[�;��;���;l��;�{y;x:l;Rs_;�*S;`G;�<;�/1;,�&;)�;��;�@	;���:���:��:g��:���:���:�З:VC�:��r:��V:C<:��":�d:-c�9�\�9�:�9/�b9��9�A�8M���������q�ȣ���͹BN��_���q(��>��TS�eh�U|�$ ��]���qۚ����[謺�ε�v�����Ǻh(Ѻ�ںy�亁F�R��f��SH�s�9���j�,��:]$���)���.��g3�y8��<�U�@��`E��I�ON���R�7�W�c�\��b��kg���l�Εr��Ax���}�FŁ�R����>���㉻�w��?����o��Yؓ��9��♘��  �  Y�=Po=!=�=|=�$=�=*o=�=� =�V =��<�@�<���<���<�A�<s��<��<Xp�<K��<�F�<���<��<7z�<'��<�-�<�~�<Q��<��<�V�<���<0��<�'�<rs�<���<��<*s�</��<,5�<�<��<�g�<���<�)�<h��<���<��<P_�<���<���<��<�(�<R�<vz�<���<���<7��<�<lA�<�d�<݃�<��<��<-��<���<��<Y]�<n�<i��<�m�<���<�z�<b��<S�<T��<��<�T�<W��< ��<d#�</_�<<�ƽ<�<2�<1,�<-;�<�?�<!:�<�*�<�<���<ѩ<���<l��<�\�<�8�<��<���<d�<�͘<��<���<���<Ǔ�<ʃ�<�o�<�V�<�7�<l�<�<���<�<#�z<�*v<��q<�Zm<�h<�d<c`<&\<��W<Z�S<̧O<�K<WjG<�HC<� ?<��:<Q�6<En2<_.<��)<�i%<�!<T�<�X<�
<��<��<Vj<�P<D��;Í�;���;'��;� �;�7�;�n�;���;Aҿ;���;�.�;f�;*��;��;c��; E�;�)�;i�x;RMk;��^;�SR;��F;�g;;��0;�M&;P;�;�,	;���:���:��:���:���:&�:�/�:�؉:*Xv:�kZ:��?:\�&:0:[w�9���9���9�!l9I094J�8I�!6I��p���ar�R1��8#йS�������+��)A��V��k�+�� 扺F`��F����s���0��ٶ�"����eȺnѺ��ں���o�����<�}���i������6��h#�M�(���-�kz2�z27�=�;�0U@���D��`I�� N��R�#�W���\��%b���g�`Mm��s�H�x��~�:,��q���r���2^���>m���ב�4��؆��&ט��  �  ��=�j=3=��=�|=*'=�=u=�=ѽ ==b =� =>]�<��<O�<�_�<���<7!�<���<���<[U�<���<��<�}�<[��<�*�<Ex�<L��<'�<QE�<��<���<d�<�U�<���<���<�T�<���<2�<��<a��<X�<?��<�!�<�}�<���<��<�d�<��<���<��<A=�<(j�<}��<���<(��<��<<8�<�\�<2}�<���<߬�<Ƿ�<4��<��<Ҋ�<�[�<X�<���<sa�<|��<�f�<���<8�<���<��<4�<�}�<���<�<�D�<�<���<��<s�<$�<�6�<�>�<Y<�<�0�<��<�<��<��<2��<~x�<8V�<Q6�<1�<R��<��<�Ԗ< Ô<�<N��<���<<u�<�X�<<6�<m�<�ރ<m��<��~<_pz<��u<��q<> m<��h<�kd<j$`<_�[<ȼW<��S<�}O<lfK<�OG<5C<?<	�:<��6<�v2<�-.<��)< �%<�2!<3�<�<#E<�<�< �<f�<��;���;~��; �;(1�;�Y�;���;���;�ʿ;{�;c�;84�;�l�;���;�6�;0ۉ;���;��w;�Zj;�];�uQ;��E;D�:;�0;��%;�;�c;�	;��:*��:�f�:;�:�{�:\9�:D��:a_�:��y:�^:�C:е*:��:oX�9���9�9��t9��$9x�8~Ʊ6L�������ut����-�ҹ�8 �q�_�-�R]D�RQZ���o�-��(؋��?��HH��A��&���d���Km��(ɺ��Ѻ�&ۺ]�����-$�����sY�4��IY�����2��z"�E�'�ݫ,��1�F^6��;��?��VD���H�w�M�>�R�/�W�y�\��Pb�a�g�u�m���s��wy�"\������n��x1��dۊ�lk���⏻iC��(���"ؖ�����  �  Q�=�e=�=�=J|=�(=(�=�y=\ =S� =�l =� =Hw�<���<!�<�z�<4��<@8�<���<!��<�a�<���<<$�<��<;��<�&�<�p�<���<(��<�3�<?q�<ׯ�<��<G9�<���<���<�7�<=��<%�<n�<���<�H�<��<��<x�<��<> �<�h�</��<���<h�<|O�<��<��</��<��<-�<�R�<u�<��<���<u��<���<h��<x��<&��<�X�< �<W��<�T�<Y��<S�<��<�</v�<���<��<�^�<���<��<K+�<�h�<���<һ<3��<�<�0�<�;�<=�<�4�<d$�<��<��<�ҧ<y��<���<q�<�Q�<�4�<��<� �<�<�Ԕ<%��<���<���<�x�<�X�<X3�<]�<=Ճ<���<��~<tIz<�u<Wq<E�l<Ƅh<M/d<��_<g�[<�W<%jS<�TO<DK<�3G<% C<�?<��:<��6<�{2<�9.<e�)<#�%<bU!<<[�<]z<�=<%
< �<��<�V�;�?�;;�;RE�;�Y�;�s�;���;Ѩ�;|��;eѷ;J�;� �;�+�;4q�;Hې;�u�;	I�;ӻv;�si;�\;+�P;E;�:;��/;Cc%;w�;J";i�;���:��::��:���:B2�:(�:v��:O��:��|:�pa:�<G:�0.:�;:���9l�9���9�V|9��*9��8���6��� ��#w�9��W�չ��h�Z�0��uG��]��1s��⃺;�������񟺠����ذ�V���R��H�ɺ�iҺqۺ��亊������������Y�I��	�h���!�S�&���+��0�a�5��i:�U*?�#�C��H�l�M�ӃR�ϧW���\���b��9h��n�Lt��z�)	������݅������R��
፻�R��窒���'��\���  �  )�= a=k= �=�{=$)=P�=�}=�%=K� =u =V =��<���<�8�<��<���<aK�<��<^�<�k�<3��<�'�<���<��<�!�<pi�<���<;��<[$�<�^�<њ�<���<M �<m�<���<)�<��<��<SZ�<���<�:�<���<1�<r�<���<��<�j�<t��<-��<#(�<g^�<���<D��<i��<��<HD�<i�<���<���<���<@��<$��<���<���<5��<�T�<��<?��<�H�<���<lA�<x��<?�<"]�<P��<���<�C�<c��<d��<��<�T�<���<�û<��<V�<�*�<�8�<|<�</7�<�)�<u�<��<��<�ĥ<e��<���<Wi�<�K�<�/�<��<���<Y�<�˒< ��<���<�z�<X�<�/�<�<L̃<瑁<N�~<W&z<��u<�)q<�l<�Ph<=�c<g�_<>[<iYW<9@S<)0O<%K<8G<BC<�><��:<D�6<�}2<-B.<��)<��%<�q!<�*<r�<�<Vm<w:<�<��<���;V��; t�;Jq�;�x�;���;"��;i��;L��;���;���;�Ч;��;�*�;���;��;e�;��u;��h;/�[;�O;liD;�v9;K/;Z�$;�F;�;��;E��:
��:���:�:^��:��:㜜:��:o:�@d:,J:� 1:W:p�:Q�9Ș�9�7�9�/9^d�8f7\Ӗ�8�!�V�y�|K����ع\���|�|3�.J���`��]v�����+R��暘�3j���ة�"�����~&º�bʺ\�Һ��ۺ��������q��������<�$������ ��	&��+�40��4���9��>���C�fpH�[dM�wR���W��]��b�7�h��wn��t�i�z��Y��=W���?��Z��b���'H��������A��+o������  �  %�=]=p=�=�z=X)=��="�=�)=n� =f{ =�$ =k��<���<'J�<��<���<�Y�<��<�<s�<���<%*�<i��<���<o�<c�<"��<���<��<P�<C��<p��<��<�X�<M��<d
�<2o�<���<�J�<��<"/�<X��<��<�l�<���<h�<l�<��<��<�0�<mi�<��<���<�<M-�<�U�<�y�<���<q��<��<���<��<���<���<Ո�<�Q�<%�<���<�>�<���<Z3�<a��<;��<~I�<���<���<p.�<�v�<��<,�<�D�<ׁ�<��<B�<�
�<c%�<v5�<p;�<�8�<�-�<��<�<�<�ҥ<��<���<�z�<Z]�<L@�<$�<��<�<�Ӓ<���<Λ�<�{�<�V�<],�<���<�ă<8��<��~<U
z<��u<�q<[�l<�(h<3�c<�_<X[<�4W<.S<�O<K<jG<��B<��><��:<,�6<	~2<wG.<
*<2�%<`�!<sD<�<`�<��<�^<'3<g<��;��;���;��;��;Ȓ�;Θ�;|��;��;��;�;m��;��;��;K�;5Ո;5��;�Vu;Uh;�`[;=TO;��C;�8;Ҙ.;��$;��;ժ;ޑ;�[�:���:���:M�:5!�:7v�:�P�:��:
��:C]f:w_L:�U3:K.:A�:^r�9�p�9Wt�9C429�(�8�k70���#�mx|����~�ڹe:��&���4��SL��
c���x��Ȇ����/ә�����7媺d�fߺ�6�º?�ʺBOӺxܺ^*�V������eO�2t���������?�Hc ��|%�ˊ*�@�/���4�gw9��c>�YOC�ZEH�kLM��qR�v�W��8]���b�6�h��n��t��{�����Z���s����\��x��������M�����?����ș��  �  �=cZ=z=��=�y=H)=Q�=��=�+=�� =? =F) =���<���<2U�<˭�<��<�b�<{��<��<Ow�<\��<	+�<��<��<h�<�^�<���<���<��<�F�<��<߼�<� �<�K�<R��<���<Bc�<���<�@�<[��<�'�<F��<�<Pi�<7��<n�<`l�<���<���<�5�<0p�<3��<��<��<,8�<�`�<D��<���<���<���<	��<���<���<Я�<���<�N�<`�<���<�8�<���<J*�<��<���<=�<���<��<� �<�i�<ʱ�<���<�:�<�x�<���<�<�<�!�<3�<~:�<�8�<�/�<� �<��<$��<Pۥ<俣<7��<⅟<7h�<�J�<l-�<��<���<�ؒ<��<o��<�{�<�U�<�)�<���<���<<C�~<a�y<#qu<E�p<�wl<�h<�c<�q_<S?[<�W<�	S< O<��J<��F<��B<K�><��:<�6<�}2<�I.<*<_�%<�!<T<*<P�<�<�u<JI<W#<� <`��;g��;��;���;a��;/��;u��;ٖ�;��;���;��;��;�Η;7"�;���;Wm�;	�t;��g;��Z;��N;r�C;Ա8;�U.;�f$;x�;l�;�w;:�:���:x��:%m�:?\�:Rʬ:d��:Y?�:J�:��g:}�M:2�4:��:):���9�/�9ʄ949�6�8�7⇘�<$$�"-~��9���eܹ�#�^9��+6���M���d��gz�M����d��R���L��^���4����d���Aú>H˺1�Ӻ>ܺ�H�ܴ�)u���;��S��y�������3�� ��$%��3*��;/�=4��89�G0>�|)C��+H��@M��qR��W��M]�c��h��n�*#u��X{����˃�ؼ��n���z@���ˎ��2���{�������̗�7虻�  �  ��=mY=�=!�=�y=M)=��= �=�,=�� =�� =�* =��<[�<�X�<T��<�<|e�<��<��<�x�<A��<`+�<��<d��<2�<D]�<���<���<��<nC�<�{�<۸�<8��<�G�<��<H��<5_�<���<a=�<Q��<%�<��<M�<�g�<@��<�<zl�<Y��<���<y7�<�r�<���<@��<��<�;�</d�<���<���<p��<L��<���<���<^��<��<a��<�M�<��<���<W6�<7��<!'�<w��<���<�8�<���<x��<N�<ee�<���<���<X7�<�u�<���<�ݹ<M�<X �<02�<<:�<9�<�0�<�!�<Z�<���<#ޥ<,ã<���<���<�k�<N�<�0�<��< ��<=ڒ<��<���<�{�<0U�<�(�<���<⽃<��<�z~<8�y< ju<u�p<�ol<�h<2�c<�h_<�6[<�W<�S<��N<�J<*�F<��B<=�><X�:<��6<�}2<�J.<�*<=�%<r�!<�Y<f<L�<d�<}<�P<W*</
 <u��;��;۩�;Ԟ�;m��;���;Y��;���;��;2��;��;3��;z;��;��;�\�;��t;�g;��Z;$�N;�nC;�8;*>.;4R$;��;,y;Tm;�+�:F��:,��:�w�:�n�:n�:��:�l�:b}�::h:E3N:!*5:��:Dt:�?�9�Ͱ9C9�9�495�8�N 7ɘ�.�$�w�~�%���[�ܹ�v�J��q�6�h,N��e���z��݇�ت���ߚ������̫�����S����hú.i˺ĮӺRܺ;U�ö�|p��15��I�Rj�Q�����������b%�>*�. /�h$4��"9�>��C��#H��<M�qR���W�CV]�|c��h�o��8u�Mq{��Ѐ�ۃ�f͆������Q��<ݎ��C��?������5ٗ�;��  �  �=cZ=z=��=�y=H)=Q�=��=�+=�� =? =F) =���<���<2U�<˭�<��<�b�<{��<��<Ow�<\��<	+�<��<��<h�<�^�<���<���<��<�F�<��<߼�<� �<�K�<R��<���<Bc�<���<�@�<[��<�'�<F��<�<Pi�<7��<n�<`l�<���<���<�5�<0p�<3��<��<��<,8�<�`�<D��<���<���<���<	��<���<���<Я�<���<�N�<`�<���<�8�<���<J*�<��<���<=�<���<��<� �<�i�<ʱ�<���<�:�<�x�<���<�<�<�!�<3�<~:�<�8�<�/�<� �<��<$��<Pۥ<忣<7��<⅟<7h�<�J�<l-�<��<���<�ؒ<��<o��<�{�<�U�<�)�<���<���<<B�~<`�y<#qu<E�p<�wl<�h<�c<�q_<S?[<�W<�	S< O<��J<��F<��B<L�><��:<�6<�}2<�I.<*<`�%<�!<T<*<Q�<�<�u<JI<W#<� <_��;f��;��;���;_��;.��;s��;ז�;��;���;��;��;�Η;6"�;���;Vm�;�t;~�g;��Z;��N;p�C;ӱ8;�U.;�f$;w�;l�;�w;:�:���:w��:%m�:?\�:Rʬ:d��:Y?�:J�:��g:}�M:1�4:��:):���9�/�9ʄ949�6�8�7⇘�<$$�"-~��9���eܹ�#�^9��+6���M���d��gz�M����d��R���L��^���4����d���Aú>H˺1�Ӻ>ܺ�H�ܴ�)u���;��S��y�������3�� ��$%��3*��;/�=4��89�G0>�|)C��+H��@M��qR��W��M]�c��h��n�*#u��X{����˃�ؼ��n���z@���ˎ��2���{�������̗�7虻�  �  %�=]=p=�=�z=X)=��="�=�)=n� =f{ =�$ =k��<���<'J�<��<���<�Y�<��<�<s�<���<%*�<i��<���<o�<c�<"��<���<��<P�<C��<p��<��<�X�<M��<d
�<2o�<���<�J�<��<"/�<X��<��<�l�<���<h�<l�<��<��<�0�<mi�<��<���<�<M-�<�U�<�y�<���<q��<��<���<��<���<���<Ո�<�Q�<%�<���<�>�<���<Z3�<a��<;��<I�<���<���<p.�<�v�<��<,�<�D�<؁�<��<B�<�
�<c%�<w5�<q;�<�8�<�-�<��<�<�<�ҥ<��<���<�z�<Z]�<L@�<$�<��<�<�Ӓ<���<Λ�<�{�<�V�<\,�<���<�ă<8��<��~<T
z<��u<�q<Z�l<�(h<3�c<�_<X[<�4W</S<�O<K<kG<��B<��><��:<-�6<~2<xG.<
*<3�%<a�!<tD<�<`�<��<�^<'3<g<��;��;���;��;��;ƒ�;˘�;y��;��;��;�;j��;��;��;	K�;3Ո;3��;�Vu;Rh;�`[;:TO;��C;�8;И.;��$;��;Ԫ;ݑ;�[�:���:���:
M�:4!�:7v�:�P�:��:
��:C]f:v_L:�U3:K.:@�:^r�9�p�9Wt�9C429�(�8�k70���#�mx|����~�ڹe:��&���4��SL��
c���x��Ȇ����/ә�����7媺d�fߺ�6�º?�ʺBOӺxܺ^*�V������eO�2t���������?�Hc ��|%�ˊ*�@�/���4�gw9��c>�YOC�ZEH�kLM��qR�v�W��8]���b�6�h��n��t��{�����Z���s����\��x��������M�����?����ș��  �  )�= a=k= �=�{=$)=P�=�}=�%=K� =u =V =��<���<�8�<��<���<aK�<��<^�<�k�<3��<�'�<���<��<�!�<pi�<���<;��<[$�<�^�<њ�<���<M �<m�<���<)�<��<��<SZ�<���<�:�<���<1�<r�<���<��<�j�<t��<-��<#(�<g^�<���<D��<i��<��<HD�<i�<���<���<���<@��<$��<���<���<5��<�T�<��<?��<�H�<���<lA�<x��<@�<"]�<Q��<���<�C�<c��<e��<��<�T�<���<�û<��<W�<�*�<�8�<}<�<07�<�)�<u�<��<��<�ĥ<e��<���<Wi�<�K�<�/�<��<���<X�<�˒<���<���<�z�<X�<�/�<�<K̃<摁<M�~<V&z<��u<�)q<�l<�Ph<=�c<g�_<?[<iYW<:@S<+0O<%K<:G<DC<�><��:<E�6<�}2</B.<��)<��%<�q!<�*<s�<�<Vm<w:<�<��<���;T��;�s�;Gq�;�x�;~��;��;d��;H��;���;���;�Ч;��;�*�;���;��;b�;��u;��h;+�[;�O;hiD;�v9;I/;X�$;�F;�;��;D��:	��:���:�:^��:��:✜:��:o:�@d:,J:� 1:W:p�:Q�9Ș�9�7�9�/9^d�8f7\Ӗ�8�!�V�y�|K����ع\���|�|3�.J���`��]v�����+R��暘�3j���ة�"�����~&º�bʺ\�Һ��ۺ��������q��������<�$������ ��	&��+�40��4���9��>���C�fpH�[dM�wR���W��]��b�7�h��wn��t�i�z��Y��=W���?��Z��b���'H��������A��+o������  �  Q�=�e=�=�=J|=�(=(�=�y=\ =S� =�l =� =Hw�<���<!�<�z�<4��<@8�<���<!��<�a�<���<<$�<��<;��<�&�<�p�<���<(��<�3�<?q�<ׯ�<��<G9�<���<���<�7�<=��<%�<n�<���<�H�<��<��<x�<��<> �<�h�</��<���<h�<|O�<��<��</��<��<-�<�R�<u�<��<���<u��<���<h��<x��<&��<�X�< �<W��<�T�<Y��<S�<��<�<0v�<���<��<�^�<���<��<L+�<�h�<���<һ<5��<�<�0�<�;�<=�<�4�<e$�<��<��<�ҧ<z��<���<q�<�Q�<�4�<��<� �<�<�Ԕ<$��<���<���<�x�<�X�<V3�<\�<<Ճ<���<�~<sIz<�u<Wq<E�l<ńh<M/d<��_<g�[<�W<'jS<�TO<DK<�3G<' C<�?<��:<��6<�{2<�9.<g�)<%�%<cU!<<\�<^z<�=<%
<�<��<�V�;�?�; ;�;NE�;�Y�;�s�;���;˨�;v��;`ѷ;E�;� �;�+�;/q�;Dې;�u�;I�;̻v;�si;�\;'�P;E;�:;ރ/;Ac%;u�;I";h�;���:��:9��:���:A2�:(�:u��:N��:��|:�pa:�<G:�0.:�;:���9l�9���9�V|9��*9��8���6��� ��#w�9��W�չ��h�Z�0��uG��]��1s��⃺;�������񟺠����ذ�V���R��H�ɺ�iҺqۺ��亊������������Y�I��	�h���!�S�&���+��0�a�5��i:�U*?�#�C��H�l�M�ӃR�ϧW���\���b��9h��n�Lt��z�)	������݅������R��
፻�R��窒���'��\���  �  ��=�j=3=��=�|=*'=�=u=�=ѽ ==b =� =>]�<��<O�<�_�<���<7!�<���<���<[U�<���<��<�}�<[��<�*�<Ex�<L��<'�<QE�<��<���<d�<�U�<���<���<�T�<���<2�<��<a��<X�<?��<�!�<�}�<���<��<�d�<��<���<��<A=�<(j�<}��<���<(��<��<<8�<�\�<2}�<���<߬�<Ƿ�<4��<��<Ҋ�<�[�<X�<���<sa�<|��<�f�<���<8�<���<��<4�<�}�<���<�<�D�<�<���<��<u�<$�<�6�<�>�<[<�<�0�<��<�<��<��<2��<~x�<8V�<Q6�<1�<Q��<��<�Ԗ<�<ﱒ<M��<���<;u�<�X�<;6�<l�<�ރ<l��<��~<]pz<��u<��q<= m<��h<�kd<j$`<`�[<ɼW<��S<�}O<nfK<�OG<5C<?<�:<��6<�v2<�-.<��)<"�%<�2!<4�<�<$E<�<�< �<e�<��;���;z��;��;#1�;�Y�;���;���;�ʿ;u�;]�;24�;�l�;���;�6�;,ۉ;���;�w;�Zj;�];�uQ;��E;A�:;�0;��%;�;�c;~	;��:(��:�f�:;�:�{�:[9�:D��:a_�:��y:�^:�C:е*:��:oX�9���9�9��t9��$9x�8~Ʊ6L�������ut����-�ҹ�8 �q�_�-�R]D�RQZ���o�-��(؋��?��HH��A��&���d���Km��(ɺ��Ѻ�&ۺ]�����-$�����sY�4��IY�����2��z"�E�'�ݫ,��1�F^6��;��?��VD���H�w�M�>�R�/�W�y�\��Pb�a�g�u�m���s��wy�"\������n��x1��dۊ�lk���⏻iC��(���"ؖ�����  �  Y�=Po=!=�=|=�$=�=*o=�=� =�V =��<�@�<���<���<�A�<s��<��<Xp�<K��<�F�<���<��<7z�<'��<�-�<�~�<Q��<��<�V�<���<0��<�'�<rs�<���<��<*s�</��<,5�<�<��<�g�<���<�)�<h��<���<��<P_�<���<���<��<�(�<R�<vz�<���<���<7��<�<lA�<�d�<݃�<��<��<-��<���<��<Y]�<n�<i��<�m�<���<�z�<b��<S�<U��<��<�T�<X��<!��<e#�<0_�<�<�ƽ<�<4�<3,�<.;�<�?�<#:�<�*�<�<���<ѩ<���<m��<�\�<�8�<��<���<c�<�͘<��<���<���<Ɠ�<Ƀ�<�o�<�V�<�7�<k�<�<���<�<!�z<�*v<��q<�Zm<�h<�d<c`< &\<��W<\�S<ͧO<��K<YjG<�HC<� ?<��:<T�6<Hn2<b.<��)<�i%<�!<V�<�X<�
<��<��<Uj<�P<B��;���;��;"��;� �;�7�;�n�;���;;ҿ;���;�.�;f�;$��;��;^��;E�;�)�;a�x;KMk;��^;�SR;��F;�g;;��0;�M&;P;�;�,	;���:���:��:���:���:&�:�/�:�؉:*Xv:�kZ:��?:\�&: 0:[w�9���9���9�!l9I094J�8I�!6I��p���ar�R1��8#йS�������+��)A��V��k�+�� 扺F`��F����s���0��ٶ�"����eȺnѺ��ں���o�����<�}���i������6��h#�M�(���-�kz2�z27�=�;�0U@���D��`I�� N��R�#�W���\��%b���g�`Mm��s�H�x��~�:,��q���r���2^���>m���ב�4��؆��&ט��  �  �=4s=3#=w�=�z=�!=i�=�h=t	=ѩ =�J =��<0#�<r�<[��<A#�<w��<3��<#Y�<���<�6�<���<�<u�<Z��<}/�<փ�<���<�<�f�<��<���<�B�<]��<���<h7�<Ґ�<���<;N�<y��<��<�u�<��<V0�<���<���<��<AX�<)��<���<��<�<9�<�^�<���<��<2��<��<}%�<�K�<5n�<��<���<ģ�<Ü�<ԅ�<s]�<	#�<���<�x�<]
�<R��<��<&m�<G��<�$�<�t�<4��<��<�?�<�x�<뫿<ٽ<6��<��<�2�<R>�<�?�<r6�<�#�<3�<��<n��<m��<�i�<@�<\�<���<�ۜ<�Ě<b��<v��<~��<䏒<셐<�y�<+i�<�S�<�7�<��<0�<t��<Z"<��z<�Wv<��q<��m<�:i<0�d</�`<4`\<)X<n�S<��O<ߨK<��G<jYC<6*?<3�:<
�6<�b2<�.<��)<H%<&� <�~<�!<��<��<�Q<+<�<��;,�;R�;���;���;�;�T�;Z��;xӿ;��;OL�;���;m�;�[�;��;���;h��;�{y;q:l;Ls_;�*S;�_G;�<;�/1;)�&;'�;��;�@	;���:���:��:f��:���:���:�З:VC�:��r:��V:C<:��":�d:,c�9�\�9�:�9/�b9��9�A�8N���������q�ȣ���͹BN��_���q(��>��TS�eh�U|�$ ��]���qۚ����[謺�ε�v�����Ǻh(Ѻ�ںy�亁F�R��f��SH�s�9���j�,��:]$���)���.��g3�y8��<�U�@��`E��I�ON���R�7�W�c�\��b��kg���l�Εr��Ax���}�FŁ�R����>���㉻�w��?����o��Yؓ��9��♘��  �  ��=%v=x$=(�=�x=�=]�=�a==ɟ =? =��<�<�T�<���<�<�i�<���<�B�<A��<�&�<ӗ�<��<�n�<E��<�/�<��<���<�(�<u�<���<��<�Z�<���<p��<%S�<ɫ�<7�<�d�<���< #�<���<z��<5�<��<���<!�<XP�<��<*��<3��<���<� �<D�<:h�<h��<���<~��<�
�<�3�<�X�<x�<H��<���<��<T��<4\�<%�<���<���<�<���<�<���<���<�@�<��<<��<��<�Y�<���<^��<��<W�<�%�<�7�<�?�<�=�<�1�<}�<���<�֫<!��<�~�<�P�<`%�<w��<�ڞ<d��<3��<�<���<���<`~�<�w�<�n�<�a�<O�<�6�<��<i�<vʁ<�;<{�z<�v<i"r<��m<�qi<w!e<��`<�\<3YX<g#T<r�O<��K<��G<IfC<E0?<��:<8�6<�U2<�-<�)<m&%<�� <~O<��<G�<YL<�<��<��<ڲ�;8��;' �;3D�;���;���;P7�;K��;DϿ;\�;�b�;0��;^�;<��;Q?�;T�;���;�Pz;+m;D`;��S;�H;¢<;��1;�';��;�;UH	;��:�.�:��:7�:η:>ܦ:
y�:���:6uo:�	S:_K8:!;:��:���9!0�9�ђ9��Y9V9ީ�8�p���J�����sp����|�˹f����&�]L;�6P�V�d���x��E��f揺�T�������ƫ�贺����cǺ��кY�ںW庸�ﺃ������C�����^q�4�����E%�Ӏ*� �/�$J4�f�8� M=��A���E��:J���N�~/S� �W��\�$�a��?g�4�l�%/r�<�w�NL}�|h���"���ц�t��^
������}������~����d���  �  z�=9x=%=Q�=�v==��=�[=~� =Ė =�4 =$��<_��<�:�<^��<e��<jQ�<Q��<u.�<Т�<�<���<���<sh�<���<�.�<ӈ�<j��<l0�<B��<4��<��<�n�<���<��<�j�<���<@�<�w�<���<�/�<��<���<18�<3��<n��<��<�H�<wy�<ԣ�<��<��<��<{,�<#O�<�t�<���<\��<.��<7�<F�<�g�<��<O��<v��<c|�<Z�<�%�<w��<>��< !�<���<�'�<"��<s��<�X�<~��<���<5�<)o�<���<TϿ<���<��<,�<�:�<@�<Z;�<J,�<��<��<=ɫ<���<Rk�<-;�<l�<�<���<z��<7��<���<pw�<r�<�n�<�j�<[d�<�Y�<J�<84�<T�<���<с<�O<?�z<.�v<+Ir<�m<<�i<Qe<�a<S�\<6�X<,FT<�P<��K<E�G<�oC<S3?<6�:<*�6<=H2<�-<y)<%<?� <�%<-�<�b<�<��
<��<�<|U�;y�;g��;��;u_�;}��;��;Mr�;�ƿ;��;"r�;Ԩ;�G�;�ԙ;���;2U�;�S�;�{;��m;:�`;;�T;�H;�=;G2;�X';A;�;DE	;��:���: ��:X��:-�:�ե:iF�:$a�:~{l:��O:�5:��:U�:���9�ô9f��9�oQ9�{9�q8[���ب��^!�ƍp��ݠ�y?ʹ�%��#"��#$�,�8�{�M���a�t�u�qЄ�f������D~���٪�{.������oǺ]�к�ںl;庁��0��aY�R7	�%���p��g� �4&�LR+�=Q0�H5���9�A�=��2B��eF���J�3�N��iS�MX���\��a�2!g��tl���q��Rw���|�o���̃��u�����歋��<��]Ð�/C��r����:���  �  ��=�y=&%=Z�=�t=�=��=�V=^� =�� =�, =��<��<�&�<{�<���<S>�<���<��<��<U�<H��<��<�b�<���<-�<���<���<�5�<t��<���<�+�<�}�<V��< &�<2|�<���<,�<���<k��<&9�<���<���<:�<���<���<C�<�A�<�p�<��<1��<��<���<�<�;�<j`�<���<ݳ�<���<V�<7�<[�<Dv�<���<��<�w�<�W�<b%�<���<ƌ�<(�<Ǵ�<�3�<Ħ�<��<j�<���<"�<�F�<`�<ɰ�<)ۿ<���<Z�<F0�<�<�<�?�<�8�<�'�<��<��<,��<H��<\�<�)�<���<qР<���<e��<�{�<Gn�<�f�<Kc�<�a�<�_�<�[�<RS�<�E�<�1�<�<6��<�Ձ<L^<�{<ιv<Rfr<�n<�i<�te<�)a<��\<U�X<`T<$P<��K<�G<�uC<�4?<��:<��6<r<2<�-<�d)<p�$<>x <�<~�<�;<��<&�
<�<��<��;�6�;�{�;���;�5�;Û�; �;a�;���;��;�{�;L�;�e�;���;���;��;͓�;J�{;�Nn;�wa;2
U;
I;Bv=;�M2;̊';�#;�;>	;FP�:M��:��:��:�A�:�:�S�:�P�:�%j:�hM:�|2:mj:�#:���9!{�9�0�9��J9��9njm8hO�]���J�"���p��v���Gɹ~��� ���"�xD7��K�|�_��s�Ҹ��w����.����*�������1����ƺ3�кG�ںLp�i\��������	�n�����Mq�)-!���&�}�+���0�L�5�x*:��w>�\�B���F���J��4O��S�"1X��\���a�g�UOl���q�
w��e|�}ျ����0��Ј��h�������������얕�����  �  i�=z=%=��=Is=�=׵=WS=_� =�� =h' =���<���<��<n�<���<E2�<a��<s�<���<��<�{�<
��<"_�<s��<�+�<���<��<=9�<I��<j��<�3�<7��<���<1�<8��<6��<�5�< ��<���<�>�<���<��<�:�<��<���<�<_=�<�j�<���<ҳ�<z��<���<[�<9/�<�S�<�{�<_��<���<��<{-�<�R�<Ao�<��<���<�t�<�U�<�$�<���<S��<X,�<���<v;�<���<;�<�u�<���<��<�Q�<j��<r��<m�<t�<W�<�2�<c=�<�>�<�6�<d$�<5�<&�<���<�<>R�<��<��<�à<���<o��<io�<�b�<#\�<�Y�<�Y�<Y�<V�<O�<sB�<�/�<��<��<J؁<�f<�{<��v<$xr<(n<��i<9�e<�?a<X�\<˱X<�oT<�0P< �K<@�G<IxC<�4?<6�:<H�6<�42<��-<�W)<d�$<�e <��<?�<�"<4�<~�
<�v<�h<5��;C�;V�;��;_�;���;1��;�T�;&��;J�;��;��;Yw�;�;�ђ;ǲ�;���;S�{;�n;�a;�VU;LI;A�=;,x2;F�';I4;�;P7	;-�:wM�:���:]��:�ε:�z�:η�:ա�:��h:��K:��0:��:n� :��9���9���93�F9��8��a8q4t�"��j�#��Rq��U��>�ȹ��{S���!�O76�pJ��}^��^r�
���ό������'������FV��������ƺl�к�ںɖ���,���/����	�����������!��'�`\,��Y1��6���:�a�>���B��
G��)K��`O�+�S��HX��]���a�Dg��9l�2�q�f�v��)|�����c��
��룈��=���ҍ��d��{�[~���
���  �  !�=L�=c2=b�=�~=�=T�=cT=&� =6� =M =.d�<���<���<<�<8��<�
�<4��<��<Ĉ�<L�<���<�<���<���< e�<���<#�<u{�<���<�'�<d~�<���<0.�<>��<���<�:�<K��<1��<�K�<���<��<�[�<���< �<gG�<���<���<!��<`�<F"�<�:�<eS�<�n�<��<9��<��<��<V�<ٓ�<���<k�<7�<3X�<�h�<�f�<(P�<%�<0��<���<�1�<B��<�>�<'��<��<�p�<���<��<E:�<j�<ő�<���<�̾<I�<`�<��<�<-״<-��<2��<�Z�<��<)٩<-��<jN�<��<�֠<ҩ�<'��<br�<rg�<�e�<�i�<�p�<�w�<�z�<9x�<�n�<�\�<{C�<�#�<���<��<�W{<�w<��r<Tn<5�i<Y�e<�Qa<��\<�X<�aT<�P<�K<F�G<�HC<��><��:<�C6<�1<~O-<��(<�($<E�<v�<4h<��<'�<�>	<�<�<T�;�V�;���;�(�;d��;��;���;���;GA�;���;߭;�6�;ܟ�;L$�;$ɏ;���;���;vKu;&�g;l�Z;8GN;�B;�c6;�+;HK ;}�;�;t�;c��:���:�0�:�̸:T��:��:�:�g:"H:�J+:s�:��9�3�9���9C�r9X�/9�Q�8l�H8��D����w�̴U�땏�����*�ܹKD��;�u*���=��Q���d��Xx�Oх��l��$����������f��\޾�(yȺ�QҺˈܺ2�b�\��#�3g�*��f��R��P$�"�)�xM/��74�;�8�r�<��@�H�D��BH���K�N�O�+�S�a:X�2�\�͢a�/�f�9�k��q��`v�~�{�Jw��[��B����I��mኻ�u�����%��� ��Щ���  �  ��= �=�2=��=�= =��=�U=� =e� =� =�i�<[��<���<(B�<B��<��<���<w�<��<��<���<��<ʍ�<��<f�<!��<�"�<Xz�< ��<-%�<�z�<���<�)�<D��<���<�5�<א�<j��<�H�<_��<]�<[�<հ�<� �<�H�<J��<��<���<�	�<G&�<�?�<�X�<#t�<ה�<M��< ��<� �<�[�<���<A��<k�<D:�<�Z�<+k�<gh�<\Q�<�%�<���<���<10�<��<�;�<6��<\�<�k�<M��<?��<O5�<�e�<��<|��<�ʾ<�޼<��<��<��<tش<���<���<P]�<8 �<:ݩ<ӗ�<�S�<`�<�ܠ<ޯ�<<��<Hx�<m�<�j�<'n�<�t�<�z�<�}�<�z�<Mp�<�]�<�C�<i#�<���<��<;S{<*�v<��r<�Jn<T�i<�e<�Ga<[�\<¥X<�ZT<xP<��K<�G<HC<p�><��:<�F6<_�1<�T-<	�(<>0$<�<��<^s<��<��<:K	<f<�<�-�;�j�;k��;�7�;K��;�&�;���;���;�E�;��;�ݭ;03�;���;=�;ӻ�;���;�t�;�$u;��g;'�Z;�$N;��A;�K6;�+;�A ;��;��;7�;\��:���:�X�:t��:��:�G�:�3�:/�g:��H:8
,:��:a��9��9��9�Su9X29!g�83O8!�-�t�������U��h��Į��~�ܹ�k�}|� �*��^>��R�ݖe�_�x��!��+���Y@��f���y!��*�����e�Ⱥ�OҺ�zܺy�GB����^�3K����o��Y(��"$���)��/�4�<�8��<��@��qD��#H�@�K�
�O���S��,X���\�D�a�b�f���k�r"q��sv���{�����'���ą�^����������������)�������  �  �=Ć=!3=\�=Ɂ=#=��=�Z=�� =�� =�! =by�<0��<���<�S�<���<L!�<���<T�<K��<��<���<�<]��<�<�h�<���<R!�<�v�<1��<�<�p�<j��<��<�s�<(��<�'�<��<G��<�?�<���<���<�X�<ư�<h�<
L�<'��<g��<��<r�<�1�<�L�<7g�<5��<��<���<���<�1�<�k�<���<g��<��<D�<c�<�q�<m�<~T�<'�<���<
��<M+�<ѵ�<(2�<���<��<�\�<��<���<�&�<UX�<���<e��<�þ<eڼ<o�<��<h�<�۴<ؿ�<9��<�e�<B*�<��<:��<�b�<�$�<J�<���<柜<G��<�|�<$y�<#{�<��<t��<���<뀌<u�<.a�<�E�<#�<1��<��<D{<��v<b�r<0n<}�i<=e<�*a<��\<��X<<FT<�P<{�K<L�G<FC<$�><�:<*O6<��1<�c-<v�(<MF$<�<C<=�<�<z�<�o	<WB<!0<�m�;���;��;e�;^��;F�;���;[�;QR�;{��;lۭ;?'�;���;���;ڔ�;�T�;H@�;�t;LMg;QOZ;��M;��A;6;��*;T  ;��;1�;�;�
�:�F�:��:K��:���:�:��:��i:;�J:11.:¹:�
�9,�9��9��|9h�89�)�81Nc8�.ֶ0돸P� BS��쎹����jzݹ	���O�0�+�ػ?���S�Vg��z�d
������&��`��Q���B嵺�-���Ⱥ;GҺVܺ������S~�������
��@���]��؞#��C)���.��y3��8�HB<��;@�hD�z�G�ƕK���O� �S�bX���\���a�;�f��k�$Kq��v��|�Z����\������ꘈ�h.��Ͻ���F���ɒ��H��Gŗ��  �  k�=��=�3=3�=��=�'=*�=�a=�� =w� =- =��<���<>�<�o�<4��<x;�<*��<,�<��<�-�<��<�'�<�<��<�k�<��<��<�p�<l��<��<�_�<~��<��<N\�<k��<��<�n�<���<�0�<&��<���<�T�<���<;�<�P�<^��<��<F��<Q"�<GC�<a�<E~�<~��<���<���<��<�L�<&��<��<���<m)�<�R�<o�<�z�<t�<�X�<�(�<��<Y��<�"�<��<�"�<���<��<�D�<��<4��<)�<�B�<Gp�<{��<x��<�Ҽ<5�<��<;�<O�<ǲ<㡰<�q�<e9�<���<*��<>z�<l>�<~	�<�ݞ<���<��<��<�<K��<V��<$��<���<m��<|�<{e�<G�<�!�<f��<��<H,{<k�v<-er<�n<��i<	Oe<b�`<p�\<�eX<�$T<_�O<o�K<�zG<�@C< ?<~�:<3[6<7�1<Az-<_�(<�g$<��<MI<U�<�P<��<�	<�z<-f<���;)��;aJ�;`��;7�;.u�;9��;s �;�b�;L��;�ӭ;-�;a�;�ɖ;�T�;D�;��;h�s;t�f;�Y;bM;�A;�5;F�*;��;��;��;: ;P[�:&��:�c�:�I�:9�:��:)T�:0l:xN:��1:�8:��9���9o�9ND�9�+C9�9p��8�kڴ� ��>=�Y�P�b���ӵ��o޹���ʭ�m-���A�@V��.j�l�}�p�������]J��5t��n���ۇ�������ȺvHҺ])ܺ��j�$����\��y
�ج�������"��h(�î-��2��17��z;�M�?��lC�CG�4#K��%O�]S�M�W���\�ފa���f��l�ޏq�w�f�|�P��ٲ��rZ�������������7���b
���z��;闻�  �  K�=��=�3=��=H�=�,=��=	j=.=�� =; =A��<}��<�>�<�<J��<�\�<���<WG�<���<`A�<��<P4�<��<��<Zn�<$��<}�<^g�<���<-��<�H�<��<(��<=�<ٕ�<���<�R�<I��<$�<4��<���<�M�<۬�<^�<U�<"��<"��<�	�<j4�<2Y�<�z�<R��<���<��<�<<�<;o�<L��<��<��<e?�<�d�<_}�<���<o{�<�\�<$)�<���<Մ�<
�<1��<4�<�t�<���<9%�<p�<S��<���<}&�<cW�<���<���<�Ǽ<\޺<��<H�<��<�β<��<���<�K�<��<�ԧ<���<_�<7,�<4�<ߜ<9ƚ<ٵ�<���<���<⦒<�<͟�<O��<���<�i�<�G�<,�<��<mv<w
{<@�v<�1r<��m<Xii<�e<o�`<~r\<1X<��S<�O<v�K<�hG<P7C<��><U�:<�g6<�2<p�-<)<�$<C <�<�<��<)9<x�	<�<�<�P�;�q�;^��;���; V�;ɬ�;���;K=�;�r�;i��;�ĭ;��;K.�;V��;p��;Y��;�x�;�s;Ӡe;.�X;�EL;�\@;j�4;`*;��;�{;մ;�.;l��:\F�:G�:�8�:���:���:��:�+p:TR:��5:��:�:N��9���9���9NIP9�A9s{�801�6>�t�y%�ddN�����i���๟:�n����/�.E�H�Y���m��ڀ��x���֓������饺 ����m���2���#ɺY_Һhܺ?,���� ��J����	����(�L���!�.Q'���,�y�1�&"6��~:���>�0�B�0�F���J�N�N��	S�#�W��p\��a���f�Xl��q���w��:}�g��>%���Ն��v��\������o���Yb������j���  �  ��=X�=[2=��=�=O1=��=�r=f=+� =�J =���<��<�f�<z��<B�<w��<8��<�e�<���<�V�<��<A�<���<��<6o�<���<��<�Z�<٠�<C��<�,�<�v�<���<��<2p�<(��<
1�<|��<��<!o�<���<�C�<���<g�<X�<��<
��<��<�G�<q�<��< ��<���<

�<�5�<od�<R��<���<���<-�<ZW�<&x�<'��<Y��<��<<_�<�'�<���<Dz�<W�<:��<��<�U�<î�<U��<�H�<��<o��<	�<@9�<�i�<���<���<�Ժ<��<;�<��<�ղ<0��<��<�_�<$*�<��<���< ��<�S�<�)�<��<��<�٘<�̖<pĔ<Z��<ط�<}��<ퟌ<.��<_l�<FF�<o�<)�<�V<2�z<�hv<�q<D�m< i<r�d<Uq`<�+\<�W<��S<ٗO<�sK<PG<�(C<��><��:<r6<2<M�-<�:)<�$<�> <��<�L<��<z�<F
<T< �<���;���;E�;�Y�;��;'��;�$�;�V�;|�;0��;ܫ�;ť;��;�-�;!��;t&�;X�;��q;�|d;*�W;�?K;�v?;W54;�s);G#;�3;l�;
-;���:1��:e��:�0�:��:�
�:Ŀ�:�Nt:űV:��::�� :љ:�a�9>˺9.��9��^9�9�h�8;�l7&^��u �0�L���������Y�0��
��3��H�4�]��yr�?4���ό�|��\�������+�����������ɺ˚Һ��ۺ���9X��N���[�17	��&�x����w� ��&��J+�J=0�J�4�!a9�5�=�"�A���E��J�^GN�z�R�gjW�(_\�4�a��g���l�Grr�KAx��~�7⁻@����h��a��)������|x��}͓�����^���  �  H�=�{=�/=�=�=$5=��=m{=h=ĺ =�Z =��<�A�<ܐ�<��<�D�<���<��<Ȅ�<���<�k�<���<AL�<n��<@�<�m�<��<?�<K�<���<���<��<�R�<���<���<�F�<���<��<w�<b��<�W�<���<�6�<ğ�<� �<�X�<��<��<c&�<=Z�<ƈ�<ϳ�<���<g�<�2�<�_�<���<��<���<��<J�<o�<���<���<%��<Q��<_�<X#�<,��<�l�<|��<�k�<U��<[3�<��<}��<M�<�`�<��<���<��<�L�<D}�<���<�Ǻ<l޸<��<s�<�ڲ<���<B��<.s�<�B�<{�<"ܥ<���<�|�<BT�<�1�<a�<��<��<���<�Ւ<�ɐ<׻�<���<̎�<�l�<>B�<��<�ց<�0<Y�z<3-v<�q<I8m<��h<&nd<r`<�[<ѩW<g�S<�cO<�JK<c1G<C<A�><6�:<'x6<�&2<=�-<C\)<P�$<ou <�<Ė<.5<w�<j�
<Bk<1J<(u�;�s�;��;
��;��;��;.F�;%h�;:|�;���;���;P��;��;]ʕ;��;М�;��~;�p;�:c;L`V;�J;�t>;IY3;��(;ś;��;�Y;;3�:��:r�:��:��:G��:̓�:`�x:�q[:{�?:Z&:�:���9�X�9��9�m9�$9E��8���7��J�6����K��ގ�[k���i�z/	�K��Ƃ6���L���b��xw�_˅�Uc������fF��L����ٱ�t깺V	º)Yʺ�Ӻ�ܺ��庨��<���4��Д�&[�!����d���$�e�)��.���3��98���<���@��-E�zI�{�M�fxR�JW��_\�;�a��Sg�Gm�s�6y���~��k���G��(��ͳ��]>��έ�����WF��|��z����  �  ��=�u=),=��=Q�=�7=��=Ԃ=f%=v� =j = =bh�<���<��<vm�<���<�6�</��<�<u~�<���<�T�<���<�<di�<���<B��<V9�<u�<��<���<�-�<@u�<o��<�<�|�<���<T�<��<�>�<ڴ�<�'�<W��<���<�V�<.��<���<�1�<�j�<z��<���<���<�+�<Z�<ň�<̷�<���<�<�>�<Je�<��<��<��<{��<)��<�\�<��<���<�\�<���<�Q�<��<�<�_�<t��<���<�4�<vv�<p��<#��<n.�<�c�<���<w��<�Ӹ<T�<W�<ݲ<�Ȱ<1��<]��<hY�<�+�<,��<�ϣ<��<�}�<�Z�<�<�<�"�<g�<0��<��<�ِ<�Ǝ<���<���<pj�<�;�<��<�Ɓ<�<�zz<Z�u<�fq<��l<zxh<�d<A�_<'�[<�_W<�@S<i,O<mK<lG<��B<��><6�:<�x6<502<H�-<�y)<o%<�� <�@<$�<%�</5<��
<־<��<��;���;f��;��;�#�;OC�;�]�;!n�;�q�;�i�;�Y�;FK�;EI�;�_�;1��;��;y};|fo;�a;�U;�H;$f=;�o2;� (;�;�c;�;&�;���:GH�:���:gս:o%�:��:�L�:��|:�`:��D:�L+: :��9���9���9�j{9R�/9þ�8c��7
G<����ҵL�D��!仹��/��w�"�$::�\Q�VMg���|�`s������������
ī������a��>.ú.1˺��Ӻ�iܺ������ ��tx�����:�����7�u�#��(���-��s2��7���;��@�%�D��H��M��JR��?W�>w\���a��g�0�m�D�s���y�������y养J���^��/捻�L������Ŕ��疻g���  �  &�=�n=z'=�=��=
9=�=��=�-=� =�w =� =R��<���<Z6�<"��< ��<�U�<&��<�$�<2��<8��<�Z�<[��<��<c�<H��<���<�&�<�]�<H��<���<�	�<�N�<���<g��<�T�<���<>2�<���<l%�<0��<��<<��<���<�R�<���<���<*:�<x�<��<���<�<gL�<�}�<��<"��<`
�<�4�<�[�<&}�<���<}��<9��<��<���<#X�<��<)��<�K�<��<�7�<H��<��<9�<:��<o��<L
�<�M�<]��<���<��<�J�<�}�<��<�Ǹ<#۶<�<ݲ<�̰<;��<���<�l�<SD�<��<U�<:ɡ<D��<��<�_�<"C�<_)�<G�<���<��<�Ύ<���<*��<�e�<J3�<)��<ѵ�<��~<�Fz<	�u<!q<��l<�'h<t�c<�w_<q>[<�W<1S<}�N<u�J<��F<&�B<��>< �:<�t6<�42<��-<�)<K4%<V� <�w<K<��<�<e@<�
<M�<b��;R]�;2L�;8K�;�T�;a�;�j�;�j�;�^�;QF�;&�;x�;��;���;�!�;��;�L|;[,n;ų`;W�S;��G;�_<;R�1;�>';�e;5�;k�
;5�;��:LO�:�.�:pd�:�:� �:$Ύ:��:O+d:oI:A0:*�:�� :���9R�9΃9�99v��8��8�k3�rh���N�'��Y˾����S!��
&�'�=��FU���k��ƀ� ���Ǒ�����@㥺�̭�%e��{ݼ��_ĺ�̺";Ժ-�ܺS����T���r'��������n�����'��`"��|'�z,��Y1��6���:��f?���C�O�H��SM��2R�>HW���\�/:b�h�b)n��at�q�z��t��􅃻}��{R����񆎻o吻�!��SB��jR��&]���  �  ˪=Vh=�"=��=�=19=?�=��=\4=^� =�� =�* =[��<���<�U�<ذ�<r�<�n�<q��<�5�<7��<���<E^�<ʹ�<��<�[�<���<��<5�<�H�<({�<��<G��<k,�<zx�<���<2�<Ğ�<2�<���<Y�<���<2�<3}�<��<KM�<Ѧ�<K��<�?�<��<���<���<�1�<bg�<e��<F��<f��<6(�<P�<Ms�<���<L��<y��<̲�<���<	��<FR�<�
�<r��<s;�<
��<��<�{�<���<�<
]�<2��<-��<�)�<�n�<K��<���<G3�<oj�<g��<T��<FҶ<�ܴ<�ڲ<�ΰ<b��<?��<e|�<�X�<3�< �<��<�<>��<f}�<�]�<]@�<�$�<�
�<>�<Ԏ<ҳ�<���<?`�<7*�<��<���<4�~<�z<�yu<c�p<LYl<��g<�|c<0_<�Z<��V<�R<��N<1�J<��F<��B<�><5�:<jm6<�42<��-<�)<�N%<=� <��<FS<�<��<u�<J<t<<��;���;H��;���;Bx�;Kt�;n�;*`�;�F�;!�;~�;#Ť;5��;���;��;��;�D{;�m;��_;B�R;�F;�v;;H�0;�&;��;Vs;�X
;�r;�i�:#6�:AQ�:�ƾ:���:�:��:���:R�g:�/M:r�3:=�:��:/��9��92ƈ9�-A9^�8�^8�/�i��\Q�<��U���7���y���(��'A�~�X�,�o�v�r9���ʖ������⧺Z��������9���~ź:ͺ��Ժ�Nݺ>>�n���������-�-z�P�����F�_l!��&���+�+o0��J5��:���>���C�nTH��-M��,R�X_W�=�\�ʅb��|h�˫n��u��h{��※� �����߉�G���	���k������᱕����������  �  ۣ=�b=,=��=*�=�8=c�=��=�8=�� =֊ =�4 =F��<(�<�m�<���<�#�<���<���<�A�<���<��<�_�<l��<�
�<U�<o��<F��<��<u7�<!g�<X��<:��<��<�\�<���<��<��<f��<{z�<��<]}�<:��<�r�<	��<�G�<)��<���<C�<ƈ�<���<��<�B�<�{�<б�<���<��<�>�<�d�<ބ�<���<���<C��< ��<���<!��<�L�<9�<���<�-�<ɥ�<��<�e�<N��<I��<�@�<��<+��<��<bT�<��<�<� �<�Z�<G��<ϰ�<8ʶ<C״<dز<"ϰ<��<���<c��<0g�<,E�<"�<W��<oڟ<���<���<�q�<PQ�<d2�<��<���<׎<ʳ�<ۊ�<�Z�<�!�<�<Z��<�~<��y<,Nu<��p<b$l<	�g<IDc<"�^<8�Z<��V<ٚR<śN<-�J<�F<d�B<��><�:<�e6<�22<�-<��)<a%<!<��<�z<�3<��<b�<�y<H<H<�;���;&��;x��;���;�~�;�l�;�S�;�/�;���;CȬ;�;x`�;�I�;�\�;٧�;�tz;�@l;�^;�R; F;�:;�0;o�%;�Z;J;�

;7;��:��:[�:?�:D�:��:u�:5��:�%j:�P:��6:��:�z:��9���9�^�9q�F9���8�8�-�oj��˒S�T&���7Ĺ���;d��+�i�C�N�[�p4s�ۤ��|�������V��w��1��QC���O��&kƺ)�ͺ��պ!�ݺ��Q�ﺦ�����������MO��z�V���� ���%��*��/���4���9��k>�cDC��$H�|M��/R�_yW���\�	�b���h�ho�U�u�� |�<:���a���k��'M��K ��r����Ց�����V
��	�����  �  F�=�^=A=��=ʇ=M8=��=V�=�;=�� =͏ =�: =���<�#�<q|�<%��<1�<��<q��<�H�<���<1�<B`�<���<��<xP�<<��<b��<4��<-,�<>Z�<݊�<N��<� �<K�<��<O�<st�<:��<�l�<���<s�<���<�k�<���<'D�<��<��<�D�<���<��<"�<wM�<��<���<A��<r"�<�L�<q�<���<,��<��<2��<���< ��<��<�H�<���<V��<�$�<��<3 �<}W�<���<B��<�.�<�q�<���<���<�C�<���<:ҿ<��<%P�<���<ǩ�<�Ķ<fӴ<6ֲ<�ΰ< ��<ꨬ<
��<'p�</P�<�.�<X�<�<*ŝ<S��<�}�<�[�<�:�<p�<@��<W؎<0��<���<�V�<�<�ك<���<�~~<>�y<<2u<x�p<�l<��g<F c<z�^<�Z<��V<�}R<�N<��J<(�F<��B<o�><��:<�_6<S02<��-<@�)<�k%<�"!<�<D�<LO<<��<:�<~c<tl�;"�;���;��;ڜ�;��;�i�;�I�;��;��;��;!k�;�5�;��;�$�;>j�;��y;��k;�9^;�Q;�E;8H:;[�/;��%;1;K�;��	;;���:���:�W�:\�:C]�:��:�t�:�_�:��k:E�Q:ſ8:� :�9	:,-�9�?�9���9��I9 ��8��8fh.��k��zaU��n����Ź<��S���,��sE���]��>u�E������)���2h��x������N������ǺNDκ��պ�޺��溑��N���z�������C�� �5��C �GL%��Q*�,Q/��K4��>9��+>��C�)	H��M��6R��W�{ ]�X�b��i�#`o�'�u��c|�r��럄�V���8���|G���ȏ����]>���B��,3������  �  ��=�]=-=��=@�=&8=��=ّ=x<=�� =�� =�< =`��<r(�<���<��<�5�<���<���<K�<���<�<`�<���<L�<�N�<��<���<��<G(�<�U�<΅�<���<���<�D�<Л�<L��<�n�<���<*h�<���<�o�<���<Oi�<���<�B�<��<���<UE�<ڍ�<���<��<Q�<b��<G��<B��<x'�<CQ�<iu�<"��<��<ظ�<S��<5��<��<�~�<G�<���<���<�!�<���<���<�R�<)��<R��<m(�<:k�<^��<���<�=�<]��<rͿ<`�<�L�<}�<0��<�¶<�Ѵ<uղ<�ΰ<���<��<��<7s�<�S�<L3�<%�<!�<ʝ<���<��<(_�<J=�<6�<j��<�؎<��<���<HU�<y�<E׃<���<�w~<��y<�(u<��p<�k<zyg<c<2�^<B�Z<�{V<�sR<'yN<�J<ɐF<�B<�><�~:<�]6<�/2<N�-<G�)</o%<�'!<�<��<�X<0<�<M�<�l<�|�;�/�;���;p��;h��;���;�h�;�E�;��;)�;���;#_�;�&�;��;P�;�T�;.�y;:�k;|
^;�PQ;d[E;:;͉/;|�%;��;ŷ;��	;T ;S��:���:X�:�)�:
q�:�>�:,��:(��:dDl:sZR:�a9:�;!:.�	:�E�9�+�9�O�9Q�J9��8A�8)W.��+���V�+痹�ƹ=���Q�0-��F��t^�
�u�1��6v������Ƣ��Ѫ�kH���\���F���:Ǻtqκ�ֺ)޺��溴�ﺛ������Z��R�����N�4� ��#%��)*�,/��*4��"9�t>�P	C�} H�KM�I8R�ՕW��,]�c�+$i�Pxo�=�u�م|�p��������Ň�a����_��ᏻ@0��HT���V���D��f+���  �  F�=�^=A=��=ʇ=M8=��=V�=�;=�� =͏ =�: =���<�#�<q|�<%��<1�<��<q��<�H�<���<1�<B`�<���<��<xP�<<��<b��<4��<-,�<>Z�<݊�<N��<� �<K�<��<O�<st�<:��<�l�<���<s�<���<�k�<���<'D�<��<��<�D�<���<��<"�<wM�<��<���<A��<r"�<�L�<q�<���<,��<��<2��<���< ��<��<�H�<���<V��<�$�<��<3 �<}W�<���<C��<�.�<�q�<���<���<�C�<���<:ҿ<��<&P�<���<ǩ�<�Ķ<gӴ<7ֲ<�ΰ<��<ꨬ<��<(p�</P�<�.�<X�<�<*ŝ<S��<�}�<�[�<�:�<p�<@��<V؎<0��<���<�V�<�<�ك<��<�~~<=�y<<2u<x�p<�l<��g<F c<z�^<�Z<��V<�}R<�N<��J<)�F<��B<p�><��:<�_6<T02<��-<A�)<�k%<�"!<�<E�<MO<<��<:�<~c<sl�;"�;���;��;ٜ�;��;�i�;�I�;��;��;��;k�;�5�;��;�$�;=j�;��y;��k;�9^;�Q;�E;6H:;Z�/;��%;1;J�;��	;;���:���:�W�:\�:C]�:��:�t�:�_�:��k:E�Q:ſ8:� :�9	:,-�9�?�9���9��I9 ��8��8fh.��k��zaU��n����Ź<��S���,��sE���]��>u�E������)���2h��x������N������ǺNDκ��պ�޺��溑��N���z�������C�� �5��C �GL%��Q*�,Q/��K4��>9��+>��C�)	H��M��6R��W�{ ]�X�b��i�#`o�'�u��c|�r��럄�V���8���|G���ȏ����]>���B��,3������  �  ۣ=�b=,=��=*�=�8=c�=��=�8=�� =֊ =�4 =F��<(�<�m�<���<�#�<���<���<�A�<���<��<�_�<l��<�
�<U�<o��<F��<��<u7�<!g�<X��<:��<��<�\�<���<��<��<f��<{z�<��<]}�<:��<�r�<	��<�G�<)��<���<C�<ƈ�<���<��<�B�<�{�<б�<���<��<�>�<�d�<ބ�<���<���<C��< ��<���<!��<�L�<:�<���<�-�<ɥ�<��<�e�<O��<J��<�@�<��<+��<��<cT�< ��<�<� �<�Z�<H��<а�<9ʶ<D״<eز<#ϰ<��<���<c��<1g�<,E�<"�<W��<oڟ<���<���<�q�<PQ�<c2�<��<���<׎<ɳ�<ڊ�<�Z�<�!�<�<Y��<
�~<��y<+Nu<��p<a$l<	�g<IDc<"�^<9�Z<��V<ښR<ƛN</�J<�F<f�B<��><	�:<�e6<�22<�-<��)<a%<!<��< {<�3<��<b�<�y< H<F<�;���;#��;u��;���;�~�;�l�;�S�;�/�;���;?Ȭ;펤;t`�;�I�;�\�;֧�;�tz;�@l;�^;�R;�F;�:;�0;m�%;�Z;I;�

;7;��:��:[�:>�:D�:��:u�:4��:�%j:�P:��6:��:�z:��9���9�^�9q�F9���8�8�-�oj��˒S�T&���7Ĺ���;d��+�i�C�N�[�p4s�ۤ��|�������V��w��1��QC���O��&kƺ)�ͺ��պ!�ݺ��Q�ﺦ�����������MO��z�V���� ���%��*��/���4���9��k>�cDC��$H�|M��/R�_yW���\�	�b���h�ho�U�u�� |�<:���a���k��'M��K ��r����Ց�����V
��	�����  �  ˪=Vh=�"=��=�=19=?�=��=\4=^� =�� =�* =[��<���<�U�<ذ�<r�<�n�<q��<�5�<7��<���<E^�<ʹ�<��<�[�<���<��<5�<�H�<({�<��<G��<k,�<zx�<���<2�<Ğ�<2�<���<Y�<���<2�<3}�<��<KM�<Ѧ�<K��<�?�<��<���<���<�1�<bg�<e��<F��<f��<6(�<P�<Ms�<���<L��<y��<̲�<���<	��<FR�<�
�<r��<s;�<��<��<�{�<���<�<]�<3��<.��<�)�<�n�<L��<���<H3�<pj�<h��<V��<HҶ<�ܴ<�ڲ<�ΰ<d��<@��<f|�<�X�<3�<!�<��<�<>��<f}�<�]�<\@�<�$�<�
�<=�<Ԏ<ѳ�<���<>`�<6*�<��<���<2�~<�z<�yu<b�p<KYl<��g<�|c<0_<�Z<��V<�R<��N<3�J<��F<��B<�><8�:<lm6<�42<��-<�)<�N%<?� <��<GS<�<��<u�<J<s<:��;���;D��;���;=x�;Ft�;n�;$`�;�F�;� �;x�;Ť;0��;���;���;��;�D{;�m;��_;=�R;�F;�v;;E�0;�&;��;Ts;�X
;�r;�i�:"6�:@Q�:�ƾ:���:�:��:���:R�g:�/M:r�3:=�:��:/��9��92ƈ9�-A9^�8�^8�/�i��\Q�<��U���7���y���(��'A�~�X�,�o�v�r9���ʖ������⧺Z��������9���~ź:ͺ��Ժ�Nݺ>>�n���������-�-z�P�����F�_l!��&���+�+o0��J5��:���>���C�nTH��-M��,R�X_W�=�\�ʅb��|h�˫n��u��h{��※� �����߉�G���	���k������᱕����������  �  &�=�n=z'=�=��=
9=�=��=�-=� =�w =� =R��<���<Z6�<"��< ��<�U�<&��<�$�<2��<8��<�Z�<[��<��<c�<H��<���<�&�<�]�<H��<���<�	�<�N�<���<g��<�T�<���<>2�<���<l%�<0��<��<<��<���<�R�<���<���<*:�<x�<��<���<�<gL�<�}�<��<"��<`
�<�4�<�[�<&}�<���<}��<:��<��<���<#X�<��<)��<�K�<��<�7�<H��<��<9�<;��<p��<M
�<�M�<^��<���<��<�J�<�}�<��<�Ǹ<%۶<�<ݲ<�̰<<��<���<�l�<TD�<��<V�<;ɡ<E��<��<�_�<!C�<^)�<F�<���<��<�Ύ<���<)��<�e�<H3�<'��<ϵ�<��~<�Fz<�u<!q<��l<�'h<t�c<�w_<r>[<�W<3S<�N<w�J<��F<)�B<��><#�:<�t6<�42<��-<�)<M4%<Y� <�w<L<��<�<e@<�
<L�<_��;N]�;.L�;3K�;�T�;a�;�j�;�j�;{^�;IF�;&�;q�;��;���;�!�;��;�L|;S,n;��`;P�S;z�G;�_<;N�1;�>';�e;3�;j�
;3�;��:JO�:�.�:od�:�:� �:$Ύ:��:O+d:oI:A0:*�:�� :���9Q�9΃9�99v��8��8�k3�rh���N�'��Y˾����S!��
&�'�=��FU���k��ƀ� ���Ǒ�����@㥺�̭�%e��{ݼ��_ĺ�̺";Ժ-�ܺS����T���r'��������n�����'��`"��|'�z,��Y1��6���:��f?���C�O�H��SM��2R�>HW���\�/:b�h�b)n��at�q�z��t��􅃻}��{R����񆎻o吻�!��SB��jR��&]���  �  ��=�u=),=��=Q�=�7=��=Ԃ=f%=v� =j = =bh�<���<��<vm�<���<�6�</��<�<u~�<���<�T�<���<�<di�<���<B��<V9�<u�<��<���<�-�<@u�<o��<�<�|�<���<T�<��<�>�<ڴ�<�'�<W��<���<�V�<.��<���<�1�<�j�<z��<���<���<�+�<Z�<ň�<̷�<���<�<�>�<Je�<��<��<��<{��<)��<�\�<��<���<�\�<���<�Q�<��<�<�_�<u��<���<�4�<wv�<q��<$��<p.�<�c�<���<y��<�Ӹ<V�<Y�<!ݲ<�Ȱ<2��<^��<jY�<�+�<-��<�ϣ<��<�}�<�Z�<�<�<�"�<f�</��<��<�ِ<�Ǝ<���<���<nj�<�;�<��<�Ɓ<�<�zz<X�u<�fq<��l<zxh<�d<B�_<(�[<�_W<�@S<k,O<oK<oG<��B<��><9�:<�x6<902<L�-<�y)<r%<�� <�@<%�<&�<05<��
<վ<��<��;���;a��;��;~#�;HC�;�]�;n�;�q�;�i�;�Y�;?K�;>I�;�_�;+��;��;y};rfo;�a;�U;�H;f=;�o2;� (;�;�c;�;$�;���:EH�:���:fս:o%�:��:�L�:��|:�`:��D:�L+: :��9���9���9�j{9R�/9þ�8c��7
G<����ҵL�D��!仹��/��w�"�$::�\Q�VMg���|�`s������������
ī������a��>.ú.1˺��Ӻ�iܺ������ ��tx�����:�����7�u�#��(���-��s2��7���;��@�%�D��H��M��JR��?W�>w\���a��g�0�m�D�s���y�������y养J���^��/捻�L������Ŕ��疻g���  �  H�=�{=�/=�=�=$5=��=m{=h=ĺ =�Z =��<�A�<ܐ�<��<�D�<���<��<Ȅ�<���<�k�<���<AL�<n��<@�<�m�<��<?�<K�<���<���<��<�R�<���<���<�F�<���<��<w�<b��<�W�<���<�6�<ğ�<� �<�X�<��<��<c&�<=Z�<ƈ�<ϳ�<���<g�<�2�<�_�<���<��<���<��<J�<o�<���<���<%��<Q��<_�<X#�<-��<�l�<|��<�k�<V��<\3�<��<~��<N�<�`�<��<���<��<�L�<F}�<���<�Ǻ<n޸<��<u�<�ڲ<���<D��</s�<�B�<|�<"ܥ<���<�|�<BT�<�1�<a�<��<��<���<Ւ<�ɐ<ջ�<���<ʎ�<�l�<<B�<��<�ց<�0<V�z<1-v<�q<H8m<��h<%nd<s`<�[<ҩW<i�S<�cO<�JK<f1G<C<E�><:�:<*x6<�&2<@�-<F\)<S�$<ru <�<Ŗ<05<x�<j�
<Bk<0J<%u�;�s�;	��;��;��;��;'F�;h�;2|�;���;���;H��; ��;Vʕ;�;ʜ�;��~;�p;|:c;D`V;�J;�t>;EY3;��(;;��;�Y;;0�:��:r�:��:��:F��:˓�:_�x:�q[:z�?:Z&:�:���9�X�9��9�m9�$9E��8���7�J�6����K��ގ�[k���i�z/	�K��Ƃ6���L���b��xw�_˅�Uc������fF��L����ٱ�t깺V	º)Yʺ�Ӻ�ܺ��庨��<���4��Д�&[�!����d���$�e�)��.���3��98���<���@��-E�zI�{�M�fxR�JW��_\�;�a��Sg�Gm�s�6y���~��k���G��(��ͳ��]>��έ�����WF��|��z����  �  ��=X�=[2=��=�=O1=��=�r=f=+� =�J =���<��<�f�<z��<B�<w��<8��<�e�<���<�V�<��<A�<���<��<6o�<���<��<�Z�<٠�<C��<�,�<�v�<���<��<2p�<(��<
1�<|��<��<!o�<���<�C�<���<g�<X�<��<
��<��<�G�<q�<��< ��<���<

�<�5�<od�<R��<���<���<-�<ZW�<&x�<'��<Y��<��<<_�<�'�<���<Dz�<W�<:��<��<�U�<Į�<V��<�H�<��<p��<
�<B9�<�i�<���<���<�Ժ<��<=�<��<�ղ<2��<��<�_�<%*�<��<���<!��<�S�<�)�<��<��<�٘<�̖<oĔ<Y��<׷�<|��<럌<,��<^l�<EF�<m�<(�<�V<0�z<�hv<�q<B�m< i<r�d<Vq`<�+\<�W<��S<ܗO<�sK<PG<�(C<��><��:<r6<2<P�-<�:)<"�$<�> <��<�L<��<{�<F
<S<��<���;���;@�;�Y�;��; ��;�$�;�V�;�{�;)��;ԫ�;�ĥ;��;�-�;��;n&�;N�;��q;�|d;#�W;�?K;�v?;S54;�s);D#;�3;j�;-;���:/��:d��:�0�:��:�
�:Ŀ�:�Nt:űV:��::�� :љ:�a�9>˺9.��9��^9�9�h�8;�l7&^��u �0�L���������Y�0��
��3��H�4�]��yr�?4���ό�|��\�������+�����������ɺ˚Һ��ۺ���9X��N���[�17	��&�x����w� ��&��J+�J=0�J�4�!a9�5�=�"�A���E��J�^GN�z�R�gjW�(_\�4�a��g���l�Grr�KAx��~�7⁻@����h��a��)������|x��}͓�����^���  �  K�=��=�3=��=H�=�,=��=	j=.=�� =; =A��<}��<�>�<�<J��<�\�<���<WG�<���<`A�<��<P4�<��<��<Zn�<$��<}�<^g�<���<-��<�H�<��<(��<=�<ٕ�<���<�R�<I��<$�<4��<���<�M�<۬�<^�<U�<"��<"��<�	�<j4�<2Y�<�z�<R��<���<��<�<<�<;o�<L��<��<��<e?�<�d�<_}�<���<o{�<�\�<$)�<���<ք�<
�<2��<5�<�t�<���<:%�<p�<T��<���<~&�<dW�<��<���<�Ǽ<^޺<��<J�<��<�β<��<���<�K�<��<�ԧ<���<_�<8,�<4�<ߜ<9ƚ<ص�<���<���<঒<�<̟�<M��<���<�i�<�G�<+�<��<kv<u
{<>�v<�1r<��m<Wii<�e<p�`<r\<1X<��S<�O<x�K<�hG<S7C<��><Y�:<�g6<�2<s�-<)<�$<E <�<�<��<*9<x�	<�<�<�P�;�q�;Z��;���;�U�;ì�;���;D=�;�r�;b��;�ĭ;��;E.�;P��;j��;S��;�x�;�s;̠e;'�X;�EL;�\@;f�4;]*;��;�{;Ӵ;�.;j��:[F�:E�:�8�:���:���:��:�+p:TR:��5:��:�:N��9���9���9NIP9�A9s{�801�6>�t�y%�ddN�����i���๟:�n����/�.E�H�Y���m��ڀ��x���֓������饺 ����m���2���#ɺY_Һhܺ?,���� ��J����	����(�L���!�.Q'���,�y�1�&"6��~:���>�0�B�0�F���J�N�N��	S�#�W��p\��a���f�Xl��q���w��:}�g��>%���Ն��v��\������o���Yb������j���  �  k�=��=�3=3�=��=�'=*�=�a=�� =w� =- =��<���<>�<�o�<4��<x;�<*��<,�<��<�-�<��<�'�<�<��<�k�<��<��<�p�<l��<��<�_�<~��<��<N\�<k��<��<�n�<���<�0�<&��<���<�T�<���<;�<�P�<^��<��<F��<Q"�<GC�<a�<E~�<~��<���<���<��<�L�<&��<��<���<m)�<�R�<o�<�z�<t�<�X�<�(�<��<Z��<�"�<��<�"�<���<��<�D�<��<5��<*�<�B�<Hp�<|��<y��<�Ҽ<7�<��<=�<P�<ǲ<塰<�q�<f9�<���<+��<>z�<l>�<~	�<�ݞ<���<��<��<���<J��<U��<#��<���<l��<|�<ze�<�F�<�!�<e��<��<F,{<i�v<,er<�n<��i<	Oe<c�`<q�\<�eX<�$T<`�O<q�K<�zG<�@C< ?<��:<5[6<9�1<Cz-<a�(<�g$<��<OI<V�<�P<��<�	<�z<,f<���;&��;]J�;\��;3�;)u�;3��;m �;�b�;F��;�ӭ;(�;a�;�ɖ;�T�;@�;�;b�s;n�f;�Y;]M;�A;�5;C�*;��;��;��;9 ;N[�:%��:�c�:�I�:8�:��:(T�:/l:wN:��1:�8:��9���9o�9ND�9�+C9�9p��8�kڴ� ��>=�Y�P�b���ӵ��o޹���ʭ�m-���A�@V��.j�l�}�p�������]J��5t��n���ۇ�������ȺvHҺ])ܺ��j�$����\��y
�ج�������"��h(�î-��2��17��z;�M�?��lC�CG�4#K��%O�]S�M�W���\�ފa���f��l�ޏq�w�f�|�P��ٲ��rZ�������������7���b
���z��;闻�  �  �=Ć=!3=\�=Ɂ=#=��=�Z=�� =�� =�! =by�<0��<���<�S�<���<L!�<���<T�<K��<��<���<�<]��<�<�h�<���<R!�<�v�<1��<�<�p�<j��<��<�s�<(��<�'�<��<G��<�?�<���<���<�X�<ư�<h�<
L�<'��<g��<��<r�<�1�<�L�<7g�<5��<��<���<���<�1�<�k�<���<g��<��<D�<c�<�q�<m�<~T�<'�<���<
��<M+�<ѵ�<)2�<���<��<�\�<��<���<�&�<VX�<���<f��<�þ<fڼ<p�<��<i�<�۴<ٿ�<:��<�e�<B*�<��<:��<�b�<�$�<J�<���<柜<F��<�|�<#y�<"{�<��<t��<���<ꀌ<u�<-a�<E�<#�<0��<��<}D{<��v<b�r<0n<|�i<=e<�*a<��\<��X<=FT<�P<|�K<N�G<FC<&�><�:<,O6<��1<�c-<x�(<NF$<��<D<>�<�<{�<�o	<WB< 0<�m�;���;	��;e�;Z��;F�;���;W�;MR�;w��;hۭ;;'�;���;���;ה�;�T�;F@�;�t;HMg;MOZ;��M;��A;6;��*;S  ;��;0�;�;�
�:�F�:��:K��:���:�:��:�i::�J:11.:¹:�
�9,�9��9��|9g�89�)�81Nc8�.ֶ0돸P� BS��쎹����jzݹ	���O�0�+�ػ?���S�Vg��z�d
������&��`��Q���B嵺�-���Ⱥ;GҺVܺ������S~�������
��@���]��؞#��C)���.��y3��8�HB<��;@�hD�z�G�ƕK���O� �S�bX���\���a�;�f��k�$Kq��v��|�Z����\������ꘈ�h.��Ͻ���F���ɒ��H��Gŗ��  �  ��= �=�2=��=�= =��=�U=� =e� =� =�i�<[��<���<(B�<B��<��<���<w�<��<��<���<��<ʍ�<��<f�<!��<�"�<Xz�< ��<-%�<�z�<���<�)�<D��<���<�5�<א�<j��<�H�<_��<]�<[�<հ�<� �<�H�<J��<��<���<�	�<G&�<�?�<�X�<#t�<ה�<M��< ��<� �<�[�<���<A��<k�<D:�<�Z�<+k�<gh�<\Q�<�%�<���<���<10�<��<�;�<6��<]�<�k�<M��<?��<O5�<�e�<��<}��<�ʾ<�޼<��<��<��<uش<���<���<P]�<9 �<:ݩ<ԗ�<�S�<a�<�ܠ<ޯ�<<��<Gx�<m�<�j�<'n�<�t�<�z�<�}�<�z�<Mp�<�]�<�C�<i#�<���<��<:S{<*�v<��r<�Jn<T�i<�e<�Ga<[�\<¥X<�ZT<yP<��K<�G<HC<q�><��:<�F6<`�1<�T-<
�(<?0$<�<��<^s<��<��<:K	<f<�<�-�;�j�;i��;�7�;J��;�&�;���;���;�E�;��;�ݭ;.3�;���;;�;ѻ�;���;�t�;�$u;��g;%�Z;�$N;��A;�K6;�+;�A ;��;��;7�;[��:���:�X�:s��:��:�G�:�3�:.�g:��H:8
,:��:a��9��9��9�Su9X29!g�83O8!�-�t�������U��h��Į��~�ܹ�k�}|� �*��^>��R�ݖe�_�x��!��+���Y@��f���y!��*�����e�Ⱥ�OҺ�zܺy�GB����^�3K����o��Y(��"$���)��/�4�<�8��<��@��qD��#H�@�K�
�O���S��,X���\�D�a�b�f���k�r"q��sv���{�����'���ą�^����������������)�������  �  �=;�=�A=��=��=d*=U�=U=R� =�s =� =-.�<�`�<͢�<?��<�[�<���< X�<���<I�<v�<+��<�9�<I��<�5�<���<U�< f�<��<}�<}q�<���<�'�<��<t��<�?�<0��<���<�U�<��<�<�r�<6��<,�<��<���<�	�<�;�<�a�<R|�<��<@��< ��<'��<!��<t
�<\@�<R��<���<��<s�<���<��<W<�<�]�< i�<�[�<�6�<���<���<�F�<u��<�Q�<|��<�%�<�{�<���<� �<�0�<�V�<�t�<���<;��<��<K��<�<m��<��<�V�<��<�֮<��<�)�<Cͧ<�r�<; �<k٠<���<kz�<3d�<Z]�<c�<\q�<���<��<j��<���<���<Î�<%t�<TQ�<�(�<��<g�{<jAw<u�r<q�n<,j<��e<Cma<Y]<��X<VT<tP<u�K<�iG<�C<k�><zm:<�5<�v1<��,<�*(<l#<	�<^�<�0<�<�<��<�<_��;��;k�;m��;���;e�;L��;)%�;���;k˺;��;�3�;�k�;���;��;���;2_�;�y|;Ӌn;�`;A�S;��F;��:;�.;�m#;|�;(6;+5;���:���:,��:N1�:��:z��:���:0(f:�lD:��$:��:^��9 i�9���9�-@9��9�8ǯ7��F������D�����ߌ��b?ʹ�M���h��.2��AE�!X�6�j���}��J�����8��������N�����z�ɺ �ӺͿݺsp� ������c��������ZD!�)�'�ay-�	�2�U�7�K�;�j�?��:C�LrF�L�I�(�L�
6P���S��W�.n\��-a��-f�Yk��p�8�u��{�#������8I���ۇ��q����6���.��/����?���  �  ��=W�=�B=��=?�=,=N�=�W=�� =�v = =�5�<�h�<9��<���<Dd�<���<�_�<8��<"��<s�<t��<y=�<e��<U8�<_��<;	�<f�<��<s�<Cn�<���<x"�<�~�<���<�8�<���<���<�P�<%��<��<aq�<���<�,�<���<���<��<t?�<�e�<��<���<���<<��<���<E��<��<�H�<}��<���<'�<iy�<{��<{�<Q@�<wa�<�k�<�]�<�7�<���<6��<"E�<���<�M�<o��<��<'u�<���<|��<*�<�P�<�o�<��<���<ç�<孻<q��<❷<#��<�Y�<,!�<�ڮ<ˈ�<�/�<�ӧ<7z�<$(�<��<��<���<Zl�<e�<j�<�w�<��<���<���<��<\��<␈<xu�<�Q�<(�<��<ݗ{<a9w<(�r<E}n<�j<�e<�_a<� ]<��X<�MT<L�O<��K<5hG<�C<r�><+q:<�6<.}1<P�,<T3(<�v#<1�< �<"@<��<%<"�<�<d
�;^-�;���;��;ՙ�;�0�;��;�2�;b��;�Ӻ;��;�4�;�h�;Y��;��;��;
J�;�I|;Xn;l�`;R�S;(�F;�v:;�.;xZ#;�;@4;t:;t�:&�:�*�:Il�:O©:B�:N�:h�f:�RE:��%:h�:Z�9ъ�9�9�D9��9v�8�5�73oԷ}*����� C�P.���(��sʹ�`�f��]8�1�2���E�s�X�'�k���~�����o'�����8��rq��z����ɺe�Ӻ,�ݺ�J�*��F����A����Ҫ��n�_	!�KV'��6-�ە2��i7�Y�;�D�?�mC�bAF��jI�c�L�P���S�E�W��]\��#a�Y+f��]k���p��u��5{��7���΂�`c�����%���� ��6����>���Ĕ��F���  �  �=��=D=v�=ӑ=�0=��=4^=�� =� =� =pK�<1��<|��<`�<X|�<���<�t�<h�<-��<7+�<���<�G�<���<?�<(��<��< f�<ֻ�<��<@d�<U��<��<�l�<Q��<%�<���<���<tB�<���<g�<�l�<T��<�-�<N��<���<_�<"I�<6q�<���<���<���<���< ��<� �<H+�<8a�<��<��<m;�<���<���<2�<�K�<�j�<Es�<�c�<d;�<���<d��<@�<2��<�A�<k��<%�<�a�<��<���<��<�?�<:a�<�|�<ђ�<@��<���<Ϭ�<���<���<Pa�<�*�<S�<̖�<�?�<;�<���<�>�<���<�<?��<ڃ�<{�<5~�<���<Ԙ�<4��<��<���<��<���<�x�<�R�<&�<��<&�{<� w<ռr<Zn<G�i<��e<�8a<��\<(�X<�3T<��O<�K<QbG<�C<��><�z:<�6<ю1<��,<=M(<�#<u�<�<l<��<�V<x�<��<�h�;n��;{��;kM�;?��;<f�;K��;zX�;���;�;��;I7�;�^�;���;z�;h�;��;��{;s�m;/)`;��R;�CF;�:;�O.;�#;/l;,;�H;tQ�:�g�:y��:7�:���:,"�:A�:&?i:��G:��(:�:�>�9ް�9��9�`O9��9��8��8*7���H��1��O!?�դ��W%���ɹ���5��0 � 4��G�@�Z�Mn�r���!�J������0ȥ� ߮��᷺P���LʺEtӺq[ݺ���!���`���p�B$�&��	a ��&�w,�)�1���6�#�:�7�>�@dB�t�E���H�H=L���O��S�g�W�&2\��	a�)%f�Cok�p�p��8v�`�{��s���������\F���؊�"g����p���锻�]���  �  ��=G�=�E=��=�=7=��=�g=�� =� =,  ==m�<���<���<>�<J��<��<��<$ �<��<WA�<���<KW�<~��<vH�<>��<;�<yd�<���<��<�S�<���<Y��<O�<���<�<-d�<��<�*�<ȑ�<���<3d�<���<�.�<ԉ�<���<��<W�<`��<C��<���<���<��<��<&�<�Q�<���<^��<��<[�<���<���<�-�<�\�<�x�<~�<k�<b?�<2��<K��<�6�< ��<R.�<���<:��<�A�<}��<���<L��<}#�<aI�<j�<���<��<2��<���<��<Ɛ�<el�<�8�<���<���<�X�<��<@��<b�<"�</�<���<Ҩ�<~��<o��<*��<���<���<���<���<��<P��<!}�<�R�<�!�<�<�h{<��v<��r<@ n<:�i<�Ve<�`<��\<EQX<�T<��O<p�K<�VG<>C<#�><��:<#6<U�1<�-<t(<��#<N<�X<��<3<��<�K<|<���;��;|R�;��;6�;���;�,�;ŏ�;\��;��;�#�;�5�;�J�;do�;߯�;`�;`��;\�z;S�l;1_;R;�kE;�O9;h�-;�";�.;�;TT;:��:��:h�:��:���:�r�:��:��l:��K:��,:�i:���9�_�9v�9��`9>�9^{�8��48���4����c���X9�� }��颹�_ɹ.h�1�l�!�dP6�މJ�4c^���q�<���<닺�*��v@��>-����
����M��c%ʺSRӺH ݺ�Q�^�'*��HL����Y�}���Z�4�%��H+�y�0�rt5���9��=�)mA���D�4H���K�L9O��S�p[W�a�[���`�P&f�x�k��q�,�v��7|�׀� ���^,��{ƈ�PV��ۍ��T��#Ò�'��b����  �  ��=��=�F=�=�=V>=�=�s=	=�� =D3 =��<��<I�<Zo�<���<HC�<���<<E�<��<P\�<���<�h�<��<�Q�<ҵ�<8�<)`�<~��<���<�<�<��<��<k'�<�~�<���<:;�<���<Q
�<�w�<S��<6W�<���<O-�<u��<|��<5+�<�f�<i��<���<^��<���<��<�/�<U�<y��<���<���<;�<��<���<b�<bF�<�p�< ��<D��<r�<TB�<#��<���<-)�<���<'�<9t�<~��<��<
[�<r��<?��<���<)�<-P�<Hr�<_��<x��<M��<���<M��<x�<�H�<7�<Ŭ<-w�<�&�<�ץ<쎣<�N�<M�<n�<�ך<�Ș<�Ė<~ǔ<�͒<�Ӑ<�Վ<Ќ<t��<̥�<C��<�P�<��<��<?{<��v<�Gr<��m<aei<S e<E�`<wR\<]X<��S<~�O<?nK<KCG<WC<��><%�:<�66<W�1<5<-<O�(<G�#<8O<̥<\<�{<�<��<�w<�\ <
��;��;%A�;��;v�;�z�;���;'�;y$�;.�; +�;8(�;�2�;�X�;v��;� �;�y;�k;�];t�P;�JD;BW8;8�,;0$";6�;�;�P;���:Ex�:4.�:��:��:��:5��:<4q:��P:�2:aX:�7�9n��9���9@Ew9u49Q�8h�q8Tl6mX����?3�4y�]ߡ�E�ɹ���p���'$��}9�C}N�Q�b��v��)������C����}�����gp��߳������?tʺ�KӺo�ܺl��*�����0��]�
�J]�����$���)��/�G�3�`_8��q<�{7@���C�'OG�&�J���N���R��W�3�[���`�Q:f���k�5�q�FVw�}� ]��i ��5҆��p�����9v��,ݐ�4��~��×��  �   �=`�=F=�=h�=E=Q�=o=�=�� =oH =���<u�<�Q�<T��<H	�<�v�<���<&n�<���<�x�<g��<@z�<W��<�Y�<���<��<X�<ߜ�<*��</�<|b�<(��<���<L�<q��<
�<\s�<���<W�<!��<uE�<��<m(�<��<��<Y5�<�u�<���<���<I��<~�<�<�<Fa�<i��<���<	��<,�<�l�<���<���<j-�<`�<���<���<ђ�<�v�<B�<X��<ҏ�<j�<G��<_��<bK�<���<���<�%�<lb�<֚�<���<��<�/�<bY�<�|�<���<>��<䩷<���<"��<�W�<� �<�߬<'��<N�<��<���<��< R�<�)�<��<��<'�<��<#�<!�<}�<�ތ<_ʊ<�<*��<1K�<��<n�<m	{<!}v<R�q<{um<� i<��d<�>`<�[<:�W<��S<�aO<�CK< 'G<�C<[�><^�:<�F6<�1<a`-<u�(</7$<�<��<�h<8�<�x<O#	<A�<�� <�;��;
��;(#�;�x�;���;4�;�+�;g7�;�+�;�;���;h�;�;0�;z{�;6x;X�i;�Y\;�RO;j�B;�&7;8�+;�d!;�J;֘;r2;K�:���:���:T��:h1�:۫�:/��:{v:AyV:��8:H:7�:���9�x�9�7�9{�J97�	9;��8ۏ�7�.��wո��-���u�������ʹ�}�����!3'��u=�TS�+�h��}��Y��๑�&����6��Le��bR��~��8�º1 ˺�|Ӻ��ܺ>N�F���
��F���
��L�E��D��"��(�R-��22�6�6���:�1�>�ǥB�gZF�#J��N�%7R���V�q�[�?�`�kf��7l��+r�K-x�U%~�� ���ل�?����=��;Ō�u1��v���ݿ���앻����  �  �==eC=�=�=J=4�=l�=c&=�� =�] =<��<�=�<���<���<=B�<��<��<���<!�<��<��<���<'��<�]�<b��<�<vK�<r��<���<���<�8�<z�<���</�<�n�<��<�@�<N��<x1�<��<�.�<l��<6�<C��<���<�;�<���<=��<���<Y�<�A�<j�<��<���<���<�)�<�c�<���<���<��<�L�<%x�<��<��<Ę�<�w�<q=�<(��<'�<���<l�<k��<I�<:g�<:��<���<�'�<�b�<���<���<7
�<�;�<If�<��<՝�< ��<��<���<�c�<3�<���<���<�u�<4�<���<a��<<��<�c�<�C�<G,�<z�<G�<x�<��<���<1�<�Њ<5��< |�</A�<2��<�e<?�z<�.v<ߘq<{m<L�h<�%d<��_<�[<�VW<�4S<�O<�K<� G<L�B<��><��:<8O6<��1<;-<�(<�p$<r�<�R<	�<�T<�<ܚ	<�]<�5<�F�;1G�;f�;��;���;�
�;-2�;�C�;�:�;@�;g�;ˮ�;��;Uh�;,z�;1;�v;Lh;ƢZ;��M;ucA;��5;��*;� ;��;w%;��;���:n	�:�U�:I��:%Y�:<8�:3��:��z:�-\:,?:�$:��
:ED�9��9|&�9ѥa9#�9��8�p�7Dw	��ȸK*���t�[��t�̹�4��
���*�nB��X�J�n��끺<����;������A��
�������Լ�35ĺ�˺��Ӻ�ܺm�DL�s.��hQ�V=	��@��@��#��� �)O&�,�+�pe0��5��]9��=��A��mE��gI��M�~�Q�I�V�:�[��a�h�f���l���r��*y��^�p���&����u������������9>���_��o��[w���  �  >�=	�=�>=��=�=�L=��=��=3=� =r =" =r�<���<&�<Ey�<_��<4L�<i��<d4�<���<�!�<��<���<�\�<���<7��<�:�<br�<���<���<��<�G�<Ƌ�<o��<�4�<���<h�<T��<!	�<���<��<��<��<D��<���<>�<)��<���<<�<5�<,e�<���<���<?��<�+�<�a�<l��<(��<��<E;�<�h�<���<���<%��<M��<�s�<~4�<���<�j�<|��<�I�<���<���<�0�<�p�<5��<_��<�(�<Ig�<c��<���<p�<)L�<Pt�<'��<���<���<���<�k�<�A�<R�<�ժ<ؚ�<3`�<�'�<��<�ğ<���<�x�<i\�<)F�<�4�<c&�<��<��<[�<nҊ<���<�s�<�2�<��<�.<��z<��u<�7q<��l<�h<�c<�Y_<�[<��V<�R<%�N<~�J<w�F<F�B<D�><a�:<{N6<G�1<��-<d!)<ģ$<�" <i�<�,<��<�_<�
<��<��<Q�;���;���;� �;��;8<�;�L�;NI�;�+�;���;1��;8Z�;.�;�ڑ;�Љ;y �;�t;H�f;��X;�K;*�?;�a4;~�);J�;��; �;f�;�j�:|��:��:�E�:@�:&��:�N�:_:x�a:sVE:��*:�:�f�9�9'��9Jmw9.�/9�p�8'� 8��ط����(�\v��5���Ϲ��������.�x G�&�^�-Pu�ln��]���#ژ��y��Km��.ذ��㷺�����źc�̺
�Ժ�ݺj.�X����]��ۅ� M������1C�;�$�!�)��.�]3�@�7�"8<�4q@���D�;�H��"M�گQ�҇V�ƺ[�~Ka��5g��gm���s��@z��V���y��~��NZ��%	��U����ِ����$
��.����蘻�  �  ��=�z= 8=y�=B�=�M=��=K�=U==,� =Ã =) =��<���<^M�<��<x�<�t�<,��<�N�<���<�-�<���<��<�W�<%��<��<f'�<�Y�<���<���<s��<�<�V�<��<���<�d�<��<SY�<?��<<m�<Z��<P��<B�<�v�<���<<�<w��<���<��<L�<���<��<���<N'�<'^�<���<���<?��<�-�<Z�<��<~��<���<��<ʗ�<Pl�<%(�<=��<�S�<���<�&�<xw�<:��<S��<F8�<t�<[��<:��<3�<w�<���<���<�0�<[^�<a�<���<���<ψ�<ko�<XK�<4�<L�<亨<L��<�T�<�$�<���<�͝<h��<e��<�j�<UR�<<�<�'�<g�<P�<Њ<���<�g�<�!�<Jҁ<��~<	?z<�u<��p<i9l<�g<�>c<��^<ѰZ<;�V<�R<��N<H�J<��F<�B<A�><�y:<�E6<m�1< �-<<)<	�$<�[ <�<�<�<w�<"x
<V5<��<خ�;�y�;�]�;�T�;�W�;�[�;�V�;U>�;�;�Ĳ;rf�;���;Y��;oM�;�)�;OC�;�Us;^�d;�*W;�KJ;U@>;��2; p(;�};};��;';���:҇�:�s�:.��:�۰:��:6Ȑ:㞁:BOf:��J:k�0:O:�:�C�9^��9�S�9��?9�s�8��A8�V��G���9�)�m<y�I𦹁�ӹܓ���	3� �K�	Bd� �{�Sψ������T��:Ϥ�N�������t?��[���OHǺ!+κ;�պ��ݺ>�溂�@C��Ew����=����~�����#��"(��-�b�1���6�|;�ډ?�y�C�^]H��L�y�Q�r�V�!�[��a�>�g�	n���t�Y{�����m6��M���5��錻�d��z������������_���  �  �=�q=�0=d�="�=�L=5�=��=E=:� =� =J: =��<��<�w�<8��<�3�<��<]��<~c�<���<�5�<ߚ�<.��<�P�<��<���<�<�A�<�i�<���<x��<���<�'�<r�<���<�4�<k��<F0�<���<N�<3��<�k�<E��<�i�<���<$7�<M��<(��<�<�]�<؛�<���<��<XO�<B��<���<���<!�<�L�<�r�<ȑ�<���<���<���<j��<�b�<��<l��<�=�<���<j�<�Q�<Ғ�<���<��<�@�<[~�<��<��<�M�<$��< پ<8�<�H�<n�<���<���<���<�o�<FQ�<v+�<D�<�Ԩ<>��<z�<�M�<"�<��<Л<���<���<�i�<`M�<2�<�<��<�ʊ<c��<SZ�<f�<.��<��~<~�y<?=u<��p<�k<�Mg<��b<M�^<�RZ<�:V<b9R<�GN<�]J<�rF<�~B<B{><Dd:<C86<��1<Y�-<0N)<=�$<�� <1&<$�<>o<<��
<��<�N<�9�;��;I��;��;P~�;�k�;OR�;�(�;��;ˎ�;u�;¤�;�,�;�ʐ;���;J��;S�q;,_c;H�U;��H;��<;�1;W';��;�?;�L;��;0�:b�:�0�:)��:�8�:7L�:��:D*�:@-j:chO:~�5:�:rj:*n�9��9x+�9�L9�y 9��Y8����7����+�8p}�G	��zع�.��C�-�6�]P�Ti�ę��6ɋ�q��dd�������A������i��W�ºb�ȺnhϺ�ֺ�c޺����F�)��>�������4�wy�ũ�5�!�Z�&��+��0��s5�>-:���>�WoC��H��L���Q���V��G\�Eb�aQh���n���u��[|�_���oބ�j��8�������&��&c���j���I�����bΙ��  �  e�=�i=j*=l�=Κ=,K=��=��=IJ=� =�� =
G =4��<�=�<���<M��<P�<��<�<�q�<��<�9�<Ț�<9��<uI�<p��<X��<o�<�-�<CR�<5u�<d��<Z��<�<�K�<��<��<׈�<��<ҟ�<�4�<���<�Y�<v��<�]�<���<�1�<]��<`��<$�<�i�<0��<��<W/�<\m�<��<c��<"�<|<�<lc�<B��<���<Ю�<ʳ�<���<���<wY�<��<��<�*�<O��<c��<�3�<7q�<��<���<��<UV�<`��<t��<�,�<�w�<ſ�<N �<U6�<�^�<Zx�<���<~�<n�<T�<V3�<Z�<,�<⾦<ؕ�<=l�<B�<��<��<�ę<T��<[z�<�X�<e8�<��<~�<(Ŋ<J��<N�<>�<u��<^�~<|�y<Nu<�Ap<H�k<� g<��b<�9^<�Z<�U<d�Q<vN</J<�JF<�]B<-`><]O:<*6<��1<��-<�X)<%<� <�P<&�<֪<�\<�<��<�<H��;UA�;C��;���;��;�p�;�G�;��;1ú;�]�;��;Y�;LӘ;�a�;��;Q�;&�p;`4b;�}T;ڰG;��;;��0;u&;P�;n�;�
;�";L�:v��:`��:]x�:�c�:x¡:���:rE�:�m:��R:ŵ9:ŝ!:�j
:N�9¼9+��9c%U9u�9�i8����a���L.�ր�w�����۹�g�����9���S�%Zm�΂�W"���|���ˡ�����k�����'��tĺʺ�xк�k׺^ߺx�V��Y2�� �BD�yr���������� �]�%�{�*��/��4�q�9�fQ>��C���G���L���Q�W�U�\�n�b�M�h�Hio�#=v�o,}�	���c�����H���I����������h� Ö��y��)���  �  �=od=�%=��==�=�I=u�=�=NM=�� =٢ =�N =���<0Q�<ʫ�<N�<[a�<g��<�<�z�<O��<�;�<ܙ�<���<�C�<���<���<&��</ �<�B�<Zc�<`��<^��<���<K3�<W��<��<"r�<���<���<'$�<4��<�M�<A��<�U�<r��<0-�<J��<���<�'�<�p�<���<���<�?�<��<c��<���<"�<�L�<6q�<���<K��<���<^��<Y��<��<�R�<7�<D��<��<e��<!��<~ �<�[�<���<���<5��<�<�<ʀ�<M��<S�<�d�<﮾<��<�)�<�T�<�o�<	|�<$z�<Al�<'U�<�7�<6�<p�<.ͦ<¦�<�~�<�U�<+�<���<�ԙ<���<s��<�_�<�;�</�<7�<���<���<�E�<���<���<�u~<<�y<��t<�p<�ek<�f<�Zb<�^<��Y<�U<y�Q<��M<�J<10F<GB<�M><�@:<K6<��1<��-<�])<@%<M� <�j<�<(�<�<f:<O�<(�<��;�t�;q�;=��;\��;�p�;�=�;|��;���;J;�;ͷ�;�&�;���;7�;P·;!�;�p;lva;)�S;a�F;�;;0;��%;�H;I*;2c
;��;C��:N!�:��:D\�:�q�:
�:}'�:s�:��n:��T:/<:$:u�:���9���9xy�9ТZ9)�
9dhq8�����j��}`0��d��%����%޹����!�[�;�3EV� �o��6��i���.��S��,����β��K���H��ź]�ʺ�0Ѻغ)�ߺ������|E�������/�\>��C�@�28 �0%�V,*�f*/��%4�Z9��>���B�"�G��L�]�Q�P(W�-�\�&�b�B"i���o�:�v���}�OV����� ��x���g ���Q���G��!��b����e���  �  ě=yb=Q$=��=F�=2I=_�=H�=5N=?� =� =uQ =��<�W�<���<��<[g�<v��<�<Q}�<���<T<�<���<���<�A�<X��<���<$��<��<>=�<2]�<l��<���<s��<�*�<҃�<���<,j�<o��<���<n�<e��<SI�<~��<�R�<��<}+�<���<��<�(�<!s�<#��<B�<ME�<��<��<���<�(�<�R�<�u�<x��<���<���<~��<���<$��<BP�<.�<\��<��<q��<7��<��<T�<R��<J��<_��<4�<Ox�<7��<��<-^�<%��<��<�%�<�P�<�l�<�y�<�x�<�k�<fU�<�8�<��<(��<Ҧ<���<`��<�\�<�1�<�<eڙ<�<���<�a�<�<�<>�<]�<Ͼ�<V��<�B�<�<���<�k~<w�y<N�t<�p<�Uk<3�f<�Ib<��]<f�Y<��U<��Q<}�M<>J<*'F<�>B<�F><P;:<>6<��1<<�-<�_)<�%<c� <s<�&<��<��<dH<��<��<R��;���;�(�;{��;ȣ�;Xp�;�9�;c��;7��;�.�;Ҩ�;��;��;��;n��;�F;l�o;�4a;�{S;��F;��:;��/;��%;�;6;�B
;�;x��:��:߆�:R�:�u�:��:gL�:c)�:�Uo:�U:��<:�$:(�:dM�9�a�92��9�o\9O�9�s8������6.1���y����߹�j�DF"�˰<�GW���p�Q���2#��R����ڣ�����J����������gźE;˺vqѺ�=غK�ߺ���$���L��>�������0���r ���$��)���.��3���8���=���B���G�~�L��Q�97W��\�v�b�NAi�
�o���v���}��p���օ�C��I���͎�B���q���e��-,��dט�Vz���  �  �=od=�%=��==�=�I=u�=�=NM=�� =٢ =�N =���<0Q�<ʫ�<N�<[a�<g��<�<�z�<O��<�;�<ܙ�<���<�C�<���<���<&��</ �<�B�<Zc�<`��<^��<���<K3�<W��<��<"r�<���<���<'$�<4��<�M�<A��<�U�<r��<0-�<J��<���<�'�<�p�<���<���<�?�<��<c��<���<"�<�L�<6q�<���<K��<���<^��<Y��<��<�R�<7�<E��<��<e��<!��< �<�[�<���<���<6��<�<�<ˀ�<N��<T�<�d�<﮾<��<�)�<�T�<�o�<
|�<%z�<Bl�<(U�<�7�<7�<p�<.ͦ<¦�<�~�<�U�<+�<���<�ԙ<���<s��<�_�<�;�<.�<6�<���<���<�E�<���<���<�u~<;�y<��t<�p<�ek<�f<�Zb<�^<��Y<�U<z�Q<��M<�J<20F<GB<�M><�@:<M6<��1<��-<�])<A%<M� <�j<�<)�<�<f:<O�<(�<��;�t�;o�;;��;Y��;�p�;�=�;y��;���;G;�;ʷ�;�&�;���;4�;N·;�;�p;iva;&�S;^�F;�;;0;��%;�H;H*;1c
;��;B��:M!�:��:C\�:�q�:	�:}'�:s�:��n:��T:/<:$:u�:���9���9xy�9ТZ9)�
9dhq8�����j��}`0��d��%����%޹����!�[�;�3EV� �o��6��i���.��S��,����β��K���H��ź]�ʺ�0Ѻغ)�ߺ������|E�������/�\>��C�@�28 �0%�V,*�f*/��%4�Z9��>���B�"�G��L�]�Q�P(W�-�\�&�b�B"i���o�:�v���}�OV����� ��x���g ���Q���G��!��b����e���  �  e�=�i=j*=l�=Κ=,K=��=��=IJ=� =�� =
G =4��<�=�<���<M��<P�<��<�<�q�<��<�9�<Ț�<9��<uI�<p��<X��<o�<�-�<CR�<5u�<d��<Z��<�<�K�<��<��<׈�<��<ҟ�<�4�<���<�Y�<v��<�]�<���<�1�<]��<`��<$�<�i�<0��<��<W/�<\m�<��<c��<"�<|<�<lc�<B��<���<Ю�<ʳ�<���<���<wY�<��<��<�*�<P��<c��<�3�<7q�<��<���<��<VV�<`��<u��<�,�<�w�<ƿ�<P �<W6�<�^�<[x�<���<�~�<n�<T�<W3�<[�<-�<⾦<ؕ�<=l�<B�<��<��<�ę<S��<[z�<�X�<d8�<��<|�<'Ŋ<H��<N�<<�<t��<\�~<z�y<Lu<�Ap<G�k<� g<��b<�9^<�Z<�U<f�Q<xN</J<�JF<�]B</`><_O:<*6<��1<��-<�X)<%<!� <�P<'�<֪<�\<�<��<�<F��;SA�;@��;���;��;�p�;�G�;�;,ú;�]�;��;Y�;GӘ;�a�;��;M�;�p;Y4b;�}T;հG;��;;��0;u&;N�;l�;�
;�";L�:u��:_��:\x�:�c�:w¡:���:rE�:�m:��R:ŵ9:ŝ!:�j
:N�9¼9+��9c%U9u�9�i8����a���L.�ր�w�����۹�g�����9���S�%Zm�΂�W"���|���ˡ�����k�����'��tĺʺ�xк�k׺^ߺx�V��Y2�� �BD�yr���������� �]�%�{�*��/��4�q�9�fQ>��C���G���L���Q�W�U�\�n�b�M�h�Hio�#=v�o,}�	���c�����H���I����������h� Ö��y��)���  �  �=�q=�0=d�="�=�L=5�=��=E=:� =� =J: =��<��<�w�<8��<�3�<��<]��<~c�<���<�5�<ߚ�<.��<�P�<��<���<�<�A�<�i�<���<x��<���<�'�<r�<���<�4�<k��<F0�<���<N�<3��<�k�<E��<�i�<���<$7�<M��<(��<�<�]�<؛�<���<��<XO�<B��<���<���<!�<�L�<�r�<ȑ�<���<���<���<j��<�b�<��<m��<�=�<���<j�<�Q�<Ӓ�<���<��<�@�<\~�<��<��<�M�<&��<"پ<:�<�H�<n�<���<���<���<�o�<HQ�<x+�<E�<�Ԩ<?��<z�<�M�<"�<��<Л<���<���<�i�<_M�< 2�<�<��<�ʊ<a��<QZ�<e�<,��<��~<|�y<==u<��p<�k<�Mg<��b<N�^<�RZ<�:V<d9R<�GN<�]J<�rF<�~B<E{><Gd:<F86<��1<\�-<3N)<@�$<�� <3&<&�<?o<<��
<��<�N<�9�;��;D��;��;I~�;�k�;GR�;�(�;��;Î�;m�;���;�,�;�ʐ;���;D��;I�q;#_c;@�U;��H;��<;�1;W';��;�?;�L;��;-�:`�:�0�:(��:�8�:6L�:��:C*�:@-j:chO:~�5:�:rj:*n�9��9x+�9�L9�y 9��Y8����7����+�8p}�G	��zع�.��C�-�6�]P�Ti�ę��6ɋ�q��dd�������A������i��W�ºb�ȺnhϺ�ֺ�c޺����F�)��>�������4�wy�ũ�5�!�Z�&��+��0��s5�>-:���>�WoC��H��L���Q���V��G\�Eb�aQh���n���u��[|�_���oބ�j��8�������&��&c���j���I�����bΙ��  �  ��=�z= 8=y�=B�=�M=��=K�=U==,� =Ã =) =��<���<^M�<��<x�<�t�<,��<�N�<���<�-�<���<��<�W�<%��<��<f'�<�Y�<���<���<s��<�<�V�<��<���<�d�<��<SY�<?��<<m�<Z��<P��<B�<�v�<���<<�<w��<���<��<L�<���<��<���<N'�<'^�<���<���<?��<�-�<Z�<��<~��<���<��<ʗ�<Pl�<%(�<>��<�S�<���<�&�<yw�<;��<T��<G8�<	t�<\��<<��<�3�<w�<ù�<���<�0�<]^�<d�<Ñ�<���<ш�<mo�<ZK�<6�<M�<庨<M��<�T�<�$�<���<�͝<g��<d��<�j�<TR�<}<�<'�<e�<M�<Њ<���<�g�<�!�<Hҁ<��~<?z<�u<��p<g9l<�g<�>c<��^<ҰZ<=�V<�R<��N<K�J<��F<
�B<E�><�y:<�E6<q�1<$�-<<)<�$<�[ < �<�<�<x�<"x
<U5<��<ծ�;�y�;�]�;�T�;�W�;�[�;�V�;L>�;	�;�Ĳ;if�;���;Q��;gM�;�)�;HC�;�Us;S�d;�*W;�KJ;N@>;��2;p(;�};y;��;%;���:χ�:�s�:,��:�۰:��:6Ȑ:㞁:AOf:��J:k�0:O:�:�C�9^��9�S�9��?9�s�8��A8�V��G���9�)�m<y�I𦹁�ӹܓ���	3� �K�	Bd� �{�Sψ������T��:Ϥ�N�������t?��[���OHǺ!+κ;�պ��ݺ>�溂�@C��Ew����=����~�����#��"(��-�b�1���6�|;�ډ?�y�C�^]H��L�y�Q�r�V�!�[��a�>�g�	n���t�Y{�����m6��M���5��錻�d��z������������_���  �  >�=	�=�>=��=�=�L=��=��=3=� =r =" =r�<���<&�<Ey�<_��<4L�<i��<d4�<���<�!�<��<���<�\�<���<7��<�:�<br�<���<���<��<�G�<Ƌ�<o��<�4�<���<h�<T��<!	�<���<��<��<��<D��<���<>�<)��<���<<�<5�<,e�<���<���<?��<�+�<�a�<l��<(��<��<E;�<�h�<���<���<%��<M��<�s�<~4�<���<�j�<|��<�I�<���<���<�0�<�p�<6��<`��<�(�<Kg�<e��<���<s�<,L�<Rt�<*��<���<ě�<���<�k�<�A�<T�<�ժ<ٚ�<5`�<�'�<��<�ğ<���<�x�<h\�<'F�<�4�<a&�<�<��<Y�<lҊ<���<�s�<�2�<��<�.<�z<��u<�7q<��l<�h<�c<�Y_<�[<��V<�R<(�N<��J<{�F<J�B<I�><f�:<�N6<L�1<��-<i!)<ȣ$<# <l�<�,<��<�_<�
<��<��<M�;���;���;� �;��;/<�;�L�;DI�;�+�;���;'��;.Z�;%�;�ڑ;�Љ;r �;�t;<�f;��X;�K;"�?;�a4;y�);F�;��;�;c�;�j�:y��: ��:�E�:@�:%��:�N�:_:w�a:sVE:��*:�:�f�9�9'��9Jmw9.�/9�p�8'� 8��ط����(�\v��5���Ϲ��������.�x G�&�^�-Pu�ln��]���#ژ��y��Km��.ذ��㷺�����źc�̺
�Ժ�ݺj.�X����]��ۅ� M������1C�;�$�!�)��.�]3�@�7�"8<�4q@���D�;�H��"M�گQ�҇V�ƺ[�~Ka��5g��gm���s��@z��V���y��~��NZ��%	��U����ِ����$
��.����蘻�  �  �==eC=�=�=J=4�=l�=c&=�� =�] =<��<�=�<���<���<=B�<��<��<���<!�<��<��<���<'��<�]�<b��<�<vK�<r��<���<���<�8�<z�<���</�<�n�<��<�@�<N��<x1�<��<�.�<l��<6�<C��<���<�;�<���<=��<���<Y�<�A�<j�<��<���<���<�)�<�c�<���<���<��<�L�<%x�<��<��<Ę�<�w�<q=�<(��<'�<���<l�<l��<J�<;g�<;��<���<�'�<�b�<���<���<9
�<�;�<Lf�<��<ם�<��<��<���<�c�<3�<���<���<�u�<4�<���<a��<<��<�c�<�C�<F,�<y�<E�<v�<��<���</�<�Њ<2��<�{�<-A�<0��<�e<<�z<�.v<ܘq<ym<K�h<�%d<��_<�[<�VW<�4S<�O<�K<� G<P�B<��><��:<=O6<��1<?-<#�(<�p$<u�<�R<�<�T<�<ܚ	<�]<�5<�F�;+G�;�e�;ܘ�;���;�
�;#2�;�C�;�:�;5�;\�;���;��;Kh�;$z�;);��v;Lh;��Z;��M;mcA;��5;��*; ;��;t%;��;���:k	�:�U�:G��:#Y�:;8�:3��:��z:�-\:,?:�$:��
:DD�9��9|&�9ѥa9#�9��8�p�7Dw	��ȸK*���t�[��t�̹�4��
���*�nB��X�J�n��끺<����;������A��
�������Լ�35ĺ�˺��Ӻ�ܺm�DL�s.��hQ�V=	��@��@��#��� �)O&�,�+�pe0��5��]9��=��A��mE��gI��M�~�Q�I�V�:�[��a�h�f���l���r��*y��^�p���&����u������������9>���_��o��[w���  �   �=`�=F=�=h�=E=Q�=o=�=�� =oH =���<u�<�Q�<T��<H	�<�v�<���<&n�<���<�x�<g��<@z�<W��<�Y�<���<��<X�<ߜ�<*��</�<|b�<(��<���<L�<q��<
�<\s�<���<W�<!��<uE�<��<m(�<��<��<Y5�<�u�<���<���<I��<~�<�<�<Fa�<i��<���<	��<,�<�l�<���<���<j-�<`�<���<���<ђ�<�v�<B�<X��<ӏ�<k�<G��<`��<cK�<���<���<�%�<mb�<ؚ�<���<��<�/�<eY�<�|�<���<A��<穷<���<$��<�W�<� �<�߬<)��<N�<��<���<��< R�<�)�<��<��<%�<��<!�<�<{�<�ތ<\ʊ<�<'��</K�<��<j�<j	{<}v<P�q<yum<� i<��d<�>`<�[<<�W<��S<�aO<�CK<'G<�C<`�><c�:<�F6<�1<f`-<y�(<37$<�<��<�h<:�<�x<O#	<@�<�� <�~�;��;��; #�;�x�;���;*�;�+�;\7�;�+�;�;���;_�;�;(�;r{�;6x;L�i;�Y\;�RO;b�B;&7;2�+;�d!;�J;Ә;p2;H�:���:���:S��:g1�:ګ�:.��:zv:@yV:��8:H:7�:���9�x�9�7�9{�J97�	9;��8ۏ�7�.��wո��-���u�������ʹ�}�����!3'��u=�TS�+�h��}��Y��๑�&����6��Le��bR��~��8�º1 ˺�|Ӻ��ܺ>N�F���
��F���
��L�E��D��"��(�R-��22�6�6���:�1�>�ǥB�gZF�#J��N�%7R���V�q�[�?�`�kf��7l��+r�K-x�U%~�� ���ل�?����=��;Ō�u1��v���ݿ���앻����  �  ��=��=�F=�=�=V>=�=�s=	=�� =D3 =��<��<I�<Zo�<���<HC�<���<<E�<��<P\�<���<�h�<��<�Q�<ҵ�<8�<)`�<~��<���<�<�<��<��<k'�<�~�<���<:;�<���<Q
�<�w�<S��<6W�<���<O-�<u��<|��<5+�<�f�<i��<���<^��<���<��<�/�<U�<y��<���<���<;�<��<���<b�<bF�<�p�< ��<D��<r�<TB�<$��<���<-)�<���<(�<:t�<��<��<[�<s��<@��<���<)�</P�<Jr�<a��<z��<O��<���<P��<x�<�H�<9�<Ŭ<.w�<�&�<�ץ<펣<�N�<M�<m�<�ך<�Ș<�Ė<|ǔ<�͒<�Ӑ<�Վ<Ќ<r��<ɥ�<@��<�P�<��<��<�>{<��v<�Gr<��m<aei<S e<F�`<xR\<_X<��S<��O<BnK<NCG<[C<��><*�:<�66<[�1<9<-<S�(<J�#<;O<Υ<^<�{<�<��<�w<�\ <��;z��;A�;���;n�;�z�;���;�;p$�;.�;�*�;/(�;�2�;�X�;o��;� �;צy;�k;�];l�P;�JD;<W8;3�,;,$";3�;�;�P;���:Bx�:2.�:��:��:��:4��:;4q:��P:�2:aX:�7�9n��9���9@Ew9u49Q�8h�q8Tl6mX����?3�4y�]ߡ�E�ɹ���p���'$��}9�C}N�Q�b��v��)������C����}�����gp��߳������?tʺ�KӺo�ܺl��*�����0��]�
�J]�����$���)��/�G�3�`_8��q<�{7@���C�'OG�&�J���N���R��W�3�[���`�Q:f���k�5�q�FVw�}� ]��i ��5҆��p�����9v��,ݐ�4��~��×��  �  ��=G�=�E=��=�=7=��=�g=�� =� =,  ==m�<���<���<>�<J��<��<��<$ �<��<WA�<���<KW�<~��<vH�<>��<;�<yd�<���<��<�S�<���<Y��<O�<���<�<-d�<��<�*�<ȑ�<���<3d�<���<�.�<ԉ�<���<��<W�<`��<C��<���<���<��<��<&�<�Q�<���<^��<��<[�<���<���<�-�<�\�<�x�<~�<k�<b?�<2��<K��<�6�<��<S.�<���<;��<�A�<~��<���<M��<#�<cI�<j�<���<��<3��<���<��<Ȑ�<fl�<�8�<���<���<�X�<��<A��<b�<"�</�<���<Ѩ�<}��<n��<)��<���<���<���<���< ��<N��<}�<�R�<�!�<�<�h{<��v<ފr<? n<9�i<�Ve<�`<��\<FQX<�T<��O<s�K<�VG<AC<&�><��:<#6<Y�1<�-<"t(<��#<P<�X<��<4<��<�K<|<���;��;xR�;
��;6�;���;�,�;���;U��;~�;�#�;�5�;�J�;]o�;ٯ�;Z�;Z��;R�z;J�l;1_;R;�kE;�O9;d�-;�";�.;�;ST;7��:��:h�:��:���:�r�:��:��l:��K:��,:�i:���9�_�9u�9��`9>�9^{�8��48���3����c���X9�� }��颹�_ɹ.h�1�l�!�dP6�މJ�4c^���q�<���<닺�*��v@��>-����
����M��c%ʺSRӺH ݺ�Q�^�'*��HL����Y�}���Z�4�%��H+�y�0�rt5���9��=�)mA���D�4H���K�L9O��S�p[W�a�[���`�P&f�x�k��q�,�v��7|�׀� ���^,��{ƈ�PV��ۍ��T��#Ò�'��b����  �  �=��=D=v�=ӑ=�0=��=4^=�� =� =� =pK�<1��<|��<`�<X|�<���<�t�<h�<-��<7+�<���<�G�<���<?�<(��<��< f�<ֻ�<��<@d�<U��<��<�l�<Q��<%�<���<���<tB�<���<g�<�l�<T��<�-�<N��<���<_�<"I�<6q�<���<���<���<���< ��<� �<H+�<8a�<��<��<m;�<���<���<2�<�K�<�j�<Es�<�c�<d;�<���<d��<	@�<2��<�A�<l��<%�<�a�<��<���<��<�?�<;a�<�|�<Ғ�<A��<���<Ь�<���<�<Ra�<�*�<T�<͖�<�?�<<�<���<�>�<���<�<?��<ك�<{�<4~�<���<Ә�<3��<��<���<��<���<�x�<�R�<&�<��<%�{<� w<Լr<
Zn<F�i<��e<�8a<��\<)�X<�3T<��O<�K<SbG<�C<��><�z:<�6<ӎ1<��,<?M(<!�#<w�<�<l<��<�V<x�<��<�h�;k��;x��;hM�;;��;7f�;F��;uX�;���;�;��;D7�;�^�;���;v�;h�;��;��{;l�m;*)`;��R;�CF;�:;�O.;�#;-l;,;�H;rQ�:�g�:x��:6�:���:+"�:A�:&?i:��G:��(:�:�>�9ް�9��9�`O9��9��8��8*7���H��1��O!?�դ��W%���ɹ���5��0 � 4��G�@�Z�Mn�r���!�J������0ȥ� ߮��᷺P���LʺEtӺq[ݺ���!���`���p�B$�&��	a ��&�w,�)�1���6�#�:�7�>�@dB�t�E���H�H=L���O��S�g�W�&2\��	a�)%f�Cok�p�p��8v�`�{��s���������\F���؊�"g����p���锻�]���  �  ��=W�=�B=��=?�=,=N�=�W=�� =�v = =�5�<�h�<9��<���<Dd�<���<�_�<8��<"��<s�<t��<y=�<e��<U8�<_��<;	�<f�<��<s�<Cn�<���<x"�<�~�<���<�8�<���<���<�P�<%��<��<aq�<���<�,�<���<���<��<t?�<�e�<��<���<���<<��<���<E��<��<�H�<}��<���<'�<iy�<{��<{�<Q@�<wa�<�k�<�]�<�7�<���<6��<"E�<���<�M�<p��<��<'u�<���<|��<*�<�P�<�o�<��<���<ħ�<死<r��<㝷<$��<�Y�<-!�<�ڮ<ˈ�<�/�<�ӧ<7z�<$(�<��<��<���<Zl�<e�<j�<�w�<��<���<���<��<[��<␈<wu�<�Q�<(�<��<ܗ{<`9w<(�r<D}n<�j<߿e<�_a<� ]<��X<�MT<M�O<��K<6hG<�C<t�><,q:<�6<0}1<Q�,<U3(<�v#<2�<!�<"@<��<%<"�<�<c
�;]-�;���;��;ә�;�0�;��;�2�;_��;�Ӻ;��;�4�;�h�;V��;��;��;J�;�I|;Xn;i�`;O�S;&�F;�v:;�.;vZ#;�;?4;s:;s�:%�:�*�:Hl�:N©:B�:N�:h�f:�RE:��%:h�:Z�9ъ�9�9�D9��9v�8�5�73oԷ}*����� C�P.���(��sʹ�`�f��]8�1�2���E�s�X�'�k���~�����o'�����8��rq��z����ɺe�Ӻ,�ݺ�J�*��F����A����Ҫ��n�_	!�KV'��6-�ە2��i7�Y�;�D�?�mC�bAF��jI�c�L�P���S�E�W��]\��#a�Y+f��]k���p��u��5{��7���΂�`c�����%���� ��6����>���Ĕ��F���  �  ��=��=�S=�=��=�7=!�=ZU=�� =�_ =W��<���<{�<(=�<&��<s��<�}�<��<��<Yi�<��<��<Nb�<N��<�t�<;��<�M�<~��<g�<Cb�<s��<��<��<��<0J�<��<�	�<�f�<!��<�!�<т�<h��<pJ�<«�<!�<�T�<ٔ�<���<Y��<^��<���<���<���<� �<��<�B�<-��<���<v1�<8��<��<_z�<��<$+�<�a�<�|�<(z�<�Z�<
!�<���<Rm�<���<Zx�<R��<gL�<��<���<k�<�<�<�U�<f�<�p�<fw�<nz�<�x�<�n�<VY�<m4�<7��<���<aU�< �<�r�<���<Â�<��<ؽ�<My�<�L�<8�<�8�<gK�<�i�<���</��<Ȏ<�Ռ<xՊ<'ƈ<���<6��<mV�<�&�<��{<U�w<"3s<+�n<uj<f<k�a<�0]<N�X<�TT<5�O<��K<BHG<��B<q�><A>:<��5<%%1<�i,<��'<A�"<ئ<��<��<��<-]
<o�<Ʊ<dQ�;v��;�&�;t��;���;���;[3�;��;��;�U�;@p�;�~�;���;S��;��;؄�;�)�;[�u;1�g;Z;P�L;��?;��2;K�&;�f;�;5;ܢ�:t�:-��:u��:3��:_��:xV�:+�f:v{A:�:y��9��99ފ9�<9���8��V8�߆6 0�F=����޸����C�9�w��}���r��'޹>���m��0'��9���K�W�]�6eo����������\���ݜ��`��4¯�����Gº4D˺�ԺG�޺P麵����� �����lH�ȵ���$���+���1��l7��$<��@�\oC��>F�;�H��(K�^�M���P�$�S�!�W���[�Ԑ`���e���j�[ p��3u��Rz�}[�&-�������:��OЉ��n�����Ʈ��QA���Ȗ��  �  ��=��=U=��=�=n:=�=�X=F� =�c =���<4��<��<�H�<��<�<���<�<(��<qq�< �<P��<�g�<��<�x�<l��<P�<���<�<=`�<���<a�<�{�<���<cA�<1��<�<�^�<��<�<��<>��<�J�<���<��<�X�<B��<���<X��<��<���<���<] �<u�<D$�<N�<���<+��<!<�<��<5�<��<���<1�<-g�<-��<�}�<f]�<�"�<���<l�<���<�s�<���<_D�<��<Q��<(�<�3�<1N�<`�<_l�<�t�<|y�<y�<�p�<\�<8�<��<ķ�<X[�<��<]z�<��<���<�"�<\ɠ<-��<yX�<MC�<�C�<U�<r�<L��<޴�<Ύ<1ی<�ي<�Ɉ<g��<̄�<�V�<[%�<I�{<��w<�%s<��n<�cj<�e<��a<@ ]<M�X<#JT<�O<��K<�GG<E�B<��><�D:<��5<�.1<�t,<Y�'< �"<��<��<�<I<u
<�<��<�~�;���;�L�;M�;���;l��;RK�;���;�/�;�c�;�z�;��;Ԓ�;z��;���;op�;X�;�u;��g;�Y;�VL;MK?;ͻ2;S�&;�Q;]�;{:;��:N��:���:l��:�
�:\�:�Æ:όg:��B:7X:~2�9���9�ԍ9�}B9�=�8�xl8��7��"o��O�׸���,,A�ruu�����A����ݹ�~����R�'�J,:��uL�}|^�up��L��!���1㓺LS�����-��} ��%º>5˺-�Ժ�i޺W麤���4� �"w����j��m���$�;c+�E�1�\7���;���?�~C���E��{H���J�}M��YP�U�S�JuW���[�d|`�	�e���j��p��Mu��yz�[��;M��^҄��^��+�K���,�����N���ϖ��  �  �=&�=IX=n=��=JA=��=�a=�� =�o =���<C�<�.�<�j�<H��<�'�<n��<{<�<���<���<�4�</��<[w�<T�<ă�< ��<�U�<¯�<�<�Y�<���<�	�<�f�<��<'�<���<���<2H�<[��<+�<w�<8��<UK�<���<N�<�b�<���<<��<��<n
�<��<��<��<@*�<E�<|p�<���<��<[�<X��<k/�<I��<��<�A�<Pu�<��<j��<dd�<o&�<���<�g�<���<Be�<���<�,�<�|�<y��<{��<�<�7�<�M�<�^�<Ll�<�u�<�y�<�t�<qc�<�A�<��<Ʊ<'l�<q�<��<W�<���< B�<��<W��<mz�<d�<b�<�p�<���<P��<Ȑ<�ގ<��<�<�ӈ<���<���<WV�<g �<T�{<�gw<|�r<��n<�/j<��e<�Za<��\<�X<�)T<��O<=�K<�DG</ C<ҳ><OV:<@�5<�I1<`�,<�'<��"<7�<��<�<�U<�
<�K<j<��;{<�;)��;�g�;�)�;Q��;x��;��;�`�;犸;{��;���;���;W��;�Ӑ;�1�;ὁ;m�t;0�f;�X;��K;��>;-2;�P&;�;Df;�B;Y�:#"�:u�:���:���:���:���:l]j:5�E:��":pz:�:�9c�9�S9��9�o�8'ֻ7#���m�W*ĸ]��9��0o��򕹓ʷ�$cܹ�a�%���(�D�;�޷N��Ba�L�s������+��dl������F˧��Ű�y����Lº�˺85Ժ��ݺ�b�"��/ ����U��N�A��e�#�2f*���0���5���:�w�>��(B�;E���G�@J���L�x�O��7S��W�/u[�/F`��le���j�>5p���u�r�z�b��h���>9��Rɇ��Z���팻-|��� ��Dy���喻�  �  {�=��=Y\=�=խ=K=��=wo=�� =l� =t =�5�<~a�<���<���<&\�<G��<%j�<��<���<VS�<���<���<>�<��<���<�\�<V��<> �<iM�<��<*��<�D�<��<p��<f\�<���<T#�<���<���<�g�<:��</J�<r��<��<]p�<ݶ�<���<~�<'�<4�<$=�< H�<>Z�<ux�<���<*��<�0�<S��<��<%V�<���<��<�Y�<���<��<k��<Wm�<t*�<��<�^�<>��<�L�<��<��<�Q�<l��<���< ��<��<S/�<!H�<j]�<`n�<�x�<�y�<�l�<UO�<��<�ڱ<ބ�<� �<4��<�B�<֥<
s�<��<�ܞ<���<��<���<ޛ�<���<5˒<��<��<Q��<R��< �<���<|��<T�<��<�{<35w<��r<DJn<��i<-ne<	a<5�\<xEX<�S<X�O<frK< <G<)C<m�><�m:<c�5<"p1<"�,<j�'<#<n2<\M<�w<��<�%<P�<z<��;~��;Ge�;���;/��;�W�;���;�_�;��;o��;�;9��;W��;�u�;���;�Ȉ;�9�;B�s;}e;�W;�QJ;B=;&@1;�%;��;m.;0A;Uh�:���:6[�:y��:N�:ǐ�:Sщ:�n:ܝJ:�a(:~�:�'�9���9�en9��"9$�8�M68�I ���)�u�.���r;/�)Lf�Cm���@���۹p�A��9f*�{�>�1xR��e�´x�����َ�>헺٠�������d��~�ºI
˺��Ӻ�2ݺ"t纍��, ��;�%��5��Y�K"�h�(���.��N4�<9��(=���@�B�C�$�F��=I��L��O�\�R��V��[�� `�[Pe��j�6�p�"(v���{�K���xB��ᅻAv�������������h����������  �  ��=��=�_=�=8�=�U=��=r=�=� =�& =�p�<s��<���<)7�<ў�<8�<{��<6:�<X��<"x�<@�<��<�,�<ܢ�<�	�<b�<���<w��<j:�<x�<��<��<�i�<X��<�"�<"��<���<�a�<���<;P�<d��<	E�<���<{"�<�}�<+��<��<�,�<�H�<�\�<�l�<P~�<Ɩ�<���<<��<�&�<�q�<,��<�%�<��<C��<d4�<�u�<��<���<-��<�t�<�+�<��<P�<���<�*�<r��<W��<��<-U�<���<���<��<��<�'�<�F�<5a�<t�<�{�< u�<�\�<�0�<��<Z��<5C�<�ܪ<�s�<��<ణ<�`�<� �<�<�ך<z͘<qі<�ߔ<�<�<��<#�<{	�<}�<�Ć<ٍ�<�M�<h�<`~{<�v<Her<��m<ii<��d<(�`<'7\<w�W<��S<�vO<NK<�)G<�C<��><ʃ:<Z6<��1<�,<�7(<�f#<s�<ٶ<��<�><׮<�D<�<���;%��;�8�;,��;�G�;���;�[�;��;���;��;?հ;���;b�;11�;��;F7�;���;�$r;��c;��U;��H;�;;��/;a�$;��;`�;";��:�c�:�D�:�:iʰ:�^�:���:(�s:%�P:�</:w':N��9�ɴ9�B�9��C9��9�p�8gŽ7�έ�,5��j��s#���\��ᎹQ�9GڹS��&{�|,-�^�B��W���k����RB��0n���J��У�e���쳺󤻺Rú;2˺�Ӻ|�ܺ����w�Vv���*�d��������� �+�&���,�--2�W�6�-%;�.�>��B�E�"H��K��CN��Q��V�H�Z���_�Je��k�4q�@�v���|��F����������]���勻�W��H�������+��eS���  �  w�=ӧ=}`=�=�=<_=6�=U�=� =B� =2C =��<E��<�.�<S��<"��<�_�<E��<�q�<��<%��<\2�<g��<9>�<��<"�<Mb�<^��<=��<2 �<iZ�<q��<���<_)�<�~�<���<�D�<ڴ�<l-�<���<>1�<ڶ�<�9�<���<9&�<���<K��<��<�G�<Bk�<*��<��<V��<\��<��<�5�<ys�<���<,�<>b�<���<$�<�V�<`��<F��<ٽ�<��<�w�<�'�<���<K:�<���<���<�N�<���<���<��<�A�<�s�<m��<���<���<�(�<M�<i�<�x�<�x�<�e�<�?�<m�<Լ�<�f�<	�<��<�K�<��</��<�m�<�?�<� �<H�<o�<�<��<�'�<�-�<�)�<t�<���<�ǆ<܉�<A�<��<�;{<��v<k�q<mem<��h<jkd<�`<ٶ[<�xW<LS<�.O<aK<�
G<�B<_�><^�:<;76<��1<�&-<w(<��#<�<�*<ys<��<�I<��<��<���;��;f �;�y�;U��;_�;���;�
�;�'�;�;�߰;͊�;A*�;*ї;�;9��;�T;�2p;v�a;��S;��F;]&:;�h.;>a#;�;�2;��;���:��:���::�:�%�:�:�+�:�#y:�W:"�6:��:�9�
�9���9�h9$9N��8� H8��/4��A�YŸ�����T��G��Ա�!�ڹb;����}�0�_�G�l�]�nfs�%ꃺŚ��þ��Y��Lp�����HQ��Z[���fĺ%�˺��Ӻ�.ܺ���h�'	��;@���
��q�6�����$�Xz*�2�/���4���8�%�<�|H@�i�C�_�F���I��vM�LLQ��U�!fZ���_�koe��{k��q�_�w��3~����Z��Ї�u�������S��Ï��H������鲗��  �  ��=��=�]=	=S�=�e=2=P�={3=�� =�_ =���<P3�<�}�<h��<:8�<Z��<�#�<Ȩ�<�3�<H��<sL�<���<�I�<���<��<�[�<��<���<���<.�<oa�<I��<P��<>2�<���<%��<�p�<���<�{�<
�<$��<�'�<ѫ�<#�<���<��<�&�<^�<��<���<~��<���<v�<�N�<���<���<��<�Q�<E��<���<�5�<�u�<���<���<���<ū�<Gs�<p�<4��<+�<�|�<���<V�<)N�<��<U��<���<�'�<�^�<q��<���<��<�1�<�V�<\n�<�t�<(h�<"H�<��<ԯ<���<l3�<�ݨ<���<3=�<k��<̽�<͎�<�k�<dT�<�G�<mC�<ED�<�E�<�C�<�8�<!�<���<2Ć<�~�<]-�<ۦ<��z<s/v<�|q<��l<oHh<��c<Qn_<�&[<o�V<��R<��N<&�J<B�F<8�B< �><ې:< C6<��1<�M-<��(<[$<zN<�<��<�g<��<��<W><� <2��;(�;o9�;y��;��;��;�D�;�H�;0!�;ϰ;�[�;�֟;+U�;
�;9��;}a};bn;eY_;�rQ;�ZD;�8;��,;�!;p�;:b;�O;���:���:�5�:��:�)�:��:1'�:�K~:g�]:�t>:Od!:��:w�9��9ꎇ9]IG9�9��8}�7^������ܨ��0P�b`���m��ݹ�`��;��5�[�M��Fe���{�d����k��i���I䣺񉫺咲�0)��f�����źɩ̺�Ժ�?ܺy�ѹﺦ����v��	����f� ���y"�(��C-��2���6���:��t>�B�L�E�RI�v�L�,�P��[U��YZ�=�_�E�e�4l���r�OCy�������������G����$��+n��B���񀔻�]��"/���  �  �=Η=�W=�=	�=�h=�
=.�=KC=!� =�z =� =Nz�<}��<�!�<I��<���< a�<���<�[�<���<&`�<���< N�<���<��<fM�<܄�<t��<���<"��<g&�<OX�<:��<���<�?�<���<#)�<Ų�<UF�<���<�y�<��<���<��<��<l��<�.�<�m�< ��<���<q �<P/�<Sa�<Y��<{��<��<�P�<B��<q��<9�<fY�<���<��<5��<M��<��<�g�<�	�<��<)��<P�<���<)��<u�<e6�<9i�<ߞ�<���<e�<W�<���<�׿<2�<�=�<�\�<�i�<c�<@I�<��<��<x��<�X�<?�<�Ŧ<,��<�B�<�
�< ۝<³�<"��<�~�<p�<f�<�]�<R�<@�<6"�<���<$��<�l�<]�<4`<��z<ɿu<��p<�El<M�g<�,c<��^<��Z<TqV<�jR<nwN<��J<B�F<7�B<-�><v�:<�?6<Z�1<�f-<��(<�@$</�<�
<{<~�<	�<�%	<��<נ <���;���;���;��;�-�;�Q�;�`�;kL�;��;��;�;�j�;Ö;o0�;+˅;nS{;�k;��\;+O;��A;$�5;A�*;�I ;ő;Gc;��; �:��: �:E��:���:���:MÑ:8c�:�\c:�E:	�):�:yK�9I��9[ �9��h9ܹ#9#V�8~$8�˚�gМ�kM�`!O�Y��*ᴹ�.��Z��J!�[�:��AT��m��S��V���i������+����ׯ�AT��K���º��Ǻ�
κ��Ժ]�ܺ���)���J��3����@����4���S �0�%�$�*�"�/�AN4�פ8��<���@���D��`H��aL�	�P�c[U���Z��7`�pbf���l���s�
�z��ƀ�����C��U6���ꌻ2_��씑�ƒ��ld��c�� ��  �  n�=��=BN==	=B�=�g=�=��=�O=�� =v� =�5 =���<��<�g�<���<�+�<���<>�<�|�<���<�l�<0��<CK�<ө�<���<�9�<�j�<h��<���<.��<���<��<�M�<���<���<b�<���<Dt�<d�<���<�T�<��<��<��<�z�<���<�/�<Vv�<���<���<0'�<`�<���<P��<^�<�T�<3��<"��<N
�<�B�<�u�<���<���<���<	��<ș�<�U�<��<�p�<��<W!�<�]�<̏�<���<)��<6�<+O�<6��<���<_�<�b�<���<w�<| �<�E�<IX�<AW�<�C�<Y�<|�<ⴭ<�v�<w7�<F��<���<��<yP�<��<��<FΙ<���<_��<���<on�<oZ�<�@�<V�<�<��<�U�<\��<�<12z<�Ou<�xp<ζk<�g<��b<�4^<��Y<��U<�Q<�N<�;J<�aF<mzB<�}><5e:<�.6<Y�1<�q-<��(<�q$<`�<h<K�<�y<�<ϴ	<�c<!<P��;s��;�r�;+g�;�j�;�m�;�`�;3�;�ݸ;�[�;���;��;�&�;Sq�;��;�Ny;��i;r�Z;��L;�?;��3;��(;�;�5;�J; �;p��:��:/^�:���:�ֳ:25�:��:;-�:�Ih:��K:
1:7�:=T :GG�9��9�P�9�=9
��8w�W8`������`�фQ�)��\帹&�������%�Q@���Z� �t�.���1���99���K��4��Q�����Vz���ĺO�ɺ�Ϻ�;ֺ(�ݺx9������y��v,�������<��k�4�#�.�(���-��N2�,�6��H;��?���C�:�G��*L���P���U�?�Z���`�J!g���m���t�R(|�h���f��5_��Ud��g����������ꖔ��G��Vؗ��_���  �  ��=~~=�C=� =a�=�d=�=��=;X=;� =�� =^L =���<WF�<]��<���<�^�<��<�)�<���<-�<9s�<��<�C�<���<��<n#�<�O�<ro�<2��<Ĝ�<P��<���<��<�R�<t��<��<t��<�;�<���<��</1�<A��<�k�<.��<�k�<���<i+�<5y�<��<�<OE�<���<L��<;�<�O�<���<}��<\��<e2�<Ia�<���<���<m��<+��<H��<���<�@�<���<�Q�<��<���<�*�<�U�<�|�<ä�<��<��<�H�<��<���<�0�<��<gǽ<E�<�,�<D�<�G�<~9�<��<w�<���<h��<�W�<�"�<%�<I��<*��<�X�<P)�<���<�ԗ<0��<��<�x�<�\�<�;�<��<�ڈ< ��<�<�<�ց<.�~<[�y<��t<�p<�7k<�f<vb<׬]<~Y<�uU<��Q<��M<��I<	 F<DB<RQ><VB:<�6<��1<�q-<�)<ה$<�! <^�<�H<j�<��<�+
<V�<ي<���;I*�;l��;��;@��;Vr�;nK�;*	�;L��;��;�M�;�s�;���;/��;��;w;u�g;U�X;ЕJ;��=;J�1;�';�';��;�7;?�;?�:��:�~�:q
�:���:Vo�:ǩ�:h�:8 l:��P:7:5�:g�:3��9�3�9���9�aQ9Qu9ɘ�8�m�	@��[��@V��������W��I��"*�&�E�Q�`�U�{�4z������z������E���Է��p��Kmº�*Ǻ�̺tѺ7�׺~�޺W纫<�&3���W�ƹ�=!�Qz�������!���&���+��0��n5� :���>�5%C��G�$!L�c�P�T�U�Pl[�$la��g���n�� v���}��r��(��
\���o��y0������ױ��{����������T����  �  �= s=�9=��=I�=�`=�=��=�]=�=�� =] =Y
 =�p�<���<h(�<N��<���<sB�<k��<a�<mu�<.��<�:�<���<H��<3�<�7�<pS�<�f�<w�<���<���<���<��<�x�<���<-t�<�<Ҷ�<;e�<E�<���<�U�<���<�\�<���<0%�<�x�<���<k�<rZ�<���<x��<[6�<Az�<���<���<�"�<�O�<�v�<o��<)��<���<���<���<�z�<�-�<���<7�<��<���<��<�'�<�I�<�n�<
��<w��<"�< _�<c��<��<�\�<��<1�<W�<;1�<�8�<�.�<��<��<ɭ<q��<�n�<A�<��<}�<=��<���<�P�<F�<��<;ƕ<i��<�}�<g[�<N5�<��<�ˈ<���<�&�<���<͌~<��y<O�t<��o<��j<� f<�a<�A]<�Y<�U<N7Q<qmM<ԬI<�E<SB<�(><� :<j�5< �1<l-<)<��$<�G <�<n�<�3<`�<��
<�-<\�<��;��;�)�;��;T��;9j�;�.�;��;�c�;"��;���;
�;��;.�;0u�;�v;f;��V;��H;)<;�e0;)�%;��;��;�P
;�;���:��:���:\h�:eG�:�n�:��:a\�:��n:/zT:�;:7�#:1�:���9j�9��9>`9ʎ9*�8���@��L���l[��,��s%¹��񹷩�<�-���I���e�-��������V��,ң��ܬ��z���Һ��%��T�ĺ�<ɺ�ͺ��Һ��غj�ߺ$��E��@z���K��v�U��@�����հ��� �W�%�gu*�fl/��^4�%B9��>���B�auG�n0L��Q�1JV���[��b���h���o�Lw���~���ֹ��$$��B����!n��L{��-:���������u���  �  �=k=$3=?�=��=�]=&= �=�`=�=׸ =$g =@ =���<D��<B�<l��<C��<%Q�<*��<3�<�u�<���<�3�<F��<Z��<�<w'�<�@�<�P�<V^�<�o�<��</��<���<�V�<D��<�T�<��<М�<)N�<#��<"��<�F�<���<&R�<���<��<w�<���<��<�f�<���<��<�N�<���<��<�	�<�8�<6a�<���<'��<���<5��<a��<r��<do�<` �<>��<�$�<A{�<͹�<���<�	�<q)�<oL�<�w�<!��<���<�>�<��<t��<�E�<���<~ֻ<��<$�<�-�<r&�<��<��<�̭<��<�|�<�S�<R*�<���<�Ϡ<���<$i�<=4�<E�<ҕ<=��<��<uY�<�/�<���<��<�t�<�<���<�c~<5cy<�at<mo<m�j<�e<�Ta<{�\<J�X<�T< Q<0<M<n�I<L�E<��A<�><!	:<a�5<�1<f-<K)<��$<�] <<<ȵ<nd<�<|�
<�b<�	<�i�;=��;lU�;���;���;;`�;��;���;p8�;;���;>;b��;�΋;�	�;�!u;se;��U;��G;�;;p/;/�$;�&;�,;�	;B�;�	�:��:7��:���:���:r[�:B�:�؅:}kp:��V:X@>:R�&:�>:�/�9g��9��9/i9u9\�8d<�5�3���D�r^_��͘��NŹޛ�����2I0���L�i�Di���{���i���������H���z��������bƺ,�ʺ�Ϻ�Ժ��ٺ٫�ͅ�iG񺈺��~M�]T��W�J�}(���������$�Σ)�l�.�#�3���8�M�=�1�B��gG��CL�NFQ��V��B\��ob�i��Bp��w�Tf�����J0������ȍ����� ���,���ֱ���)��~���ɚ��  �  ��=;h=�0=2�=�=�\=�
=2�=~a=�=f� =�j =X =s��<0��<�J�<b��<���<�U�<J��<��<yu�<���<61�<���<��<���<�!�<�9�<[I�<�U�<7f�<~��<��<��<�J�<���<�I�<��<ݓ�<6F�<"��<��<dA�<@��<CN�<���<��<$v�<3��<<�<�j�<���<_�<^W�<i��<���< �<A@�<g�<ԇ�<���<���<X��<B��<O��<[k�<��<���<��<t�<���<���<i��<@�<�@�<Lk�<��<;��<�3�<��<t��<�=�<���<%л<V�<S�<�)�<i#�<�<�<�ͭ<���<��<Z�<2�<@�<�ؠ<���<wq�<h;�<��<�Օ<P��<[��<xX�<�-�<m��<6��<�o�<��<w��<3U~<�Ry<jOt<{Xo<7|j<��e<�<a<��\<��X<�T<�P<N+M<erI<�E<��A<]><� :<��5<�1<bc-<�)<�$<�d <�<��<*u<�#<��
<�t<<r��;���;pc�;A��;���;�[�;��;��;�(�;�y�;[��;6��;���;?��;��;�t;��d;��U;��G;��:;8/;��$;��;>�;�~	;p[;��:���:���:T��:ܲ:�O�:&N�:���:��p:�bW:@/?:��':L[:Zi�9@��9��9W#l9�99ޒ�8���5�搸�;���`�����rƹ��������%1�Z�M��6j����/(��� ��󲦺i����=��Uh��Z�º��ƺ1˺sϺaԺ�)ں�����s�����P�WJ�h@�}%����!��Ј��g$��])�5i.�r�3�X�8��=���B�feG��LL��XQ�ުV�c\�u�b�RKi��up�2�w�l������LY��:Њ�+��������#���(��-ۖ� O��
����暻�  �  �=k=$3=?�=��=�]=&= �=�`=�=׸ =$g =@ =���<D��<B�<l��<C��<%Q�<*��<3�<�u�<���<�3�<F��<Z��<�<w'�<�@�<�P�<V^�<�o�<��</��<���<�V�<D��<�T�<��<М�<)N�<#��<"��<�F�<���<&R�<���<��<w�<���<��<�f�<���<��<�N�<���<��<�	�<�8�<6a�<���<'��<���<5��<a��<r��<do�<` �<>��<�$�<A{�<͹�<���<�	�<r)�<pL�<�w�<"��< ��<�>�<��<u��<�E�<���<ֻ<��<$�<�-�<s&�<��<��<�̭<��<�|�<�S�<S*�<���<�Ϡ<���<#i�<=4�<E�<ҕ<<��<��<tY�<�/�<���<��<�t�<~�<���<�c~<4cy<�at<mo<l�j<�e<�Ta<{�\<J�X<�T< Q<1<M<p�I<M�E<��A<�><#	:<c�5<�1<f-<M)<��$<�] <=<ȵ<od<�<|�
<�b<�	<�i�;;��;iU�;���;���;7`�;��;���;l8�;댯;���;:;_��;�΋;�	�;�!u;ne;��U;��G;�;;p/;-�$;�&;�,;�	;A�;�	�:��:6��:���:���:r[�:B�:�؅:|kp:��V:X@>:R�&:�>:�/�9g��9��9/i9u9\�8e<�5�3���D�r^_��͘��NŹޛ�����2I0���L�i�Di���{���i���������H���z��������bƺ,�ʺ�Ϻ�Ժ��ٺ٫�ͅ�iG񺈺��~M�]T��W�J�}(���������$�Σ)�l�.�#�3���8�M�=�1�B��gG��CL�NFQ��V��B\��ob�i��Bp��w�Tf�����J0������ȍ����� ���,���ֱ���)��~���ɚ��  �  �= s=�9=��=I�=�`=�=��=�]=�=�� =] =Y
 =�p�<���<h(�<N��<���<sB�<k��<a�<mu�<.��<�:�<���<H��<3�<�7�<pS�<�f�<w�<���<���<���<��<�x�<���<-t�<�<Ҷ�<;e�<E�<���<�U�<���<�\�<���<0%�<�x�<���<k�<rZ�<���<x��<[6�<Az�<���<���<�"�<�O�<�v�<o��<)��<���<���<���<�z�<�-�<���<7�<��<���<��<�'�<�I�<�n�<��<x��<#�<_�<d��<��<�\�<��<2�<Y�<=1�<�8�<�.�<��<��<ɭ<r��<�n�<A�<��<~�<=��<���<�P�<E�<��<:ƕ<g��<�}�<e[�<M5�<��<�ˈ<���<�&�<���<ʌ~<��y<M�t<��o<��j<� f<�a<�A]<�Y< U<O7Q<smM<֬I<�E<VB<�(><� :<m�5<�1<l-<)<��$<�G < �<o�<�3<a�<��
<�-<[�<��;��;�)�;��;N��;3j�;�.�;��;�c�;��;���;
�;��;.�;*u�;�v;�f;��V;��H;#<;�e0;%�%;��;��;�P
;�;���:��:���:[h�:eG�:�n�:��:a\�:��n:.zT:�;:7�#:1�:���9j�9��9>`9ʎ9*�8���@��L���l[��,��s%¹��񹷩�<�-���I���e�-��������V��,ң��ܬ��z���Һ��%��T�ĺ�<ɺ�ͺ��Һ��غj�ߺ$��E��@z���K��v�U��@�����հ��� �W�%�gu*�fl/��^4�%B9��>���B�auG�n0L��Q�1JV���[��b���h���o�Lw���~���ֹ��$$��B����!n��L{��-:���������u���  �  ��=~~=�C=� =a�=�d=�=��=;X=;� =�� =^L =���<WF�<]��<���<�^�<��<�)�<���<-�<9s�<��<�C�<���<��<n#�<�O�<ro�<2��<Ĝ�<P��<���<��<�R�<t��<��<t��<�;�<���<��</1�<A��<�k�<.��<�k�<���<i+�<5y�<��<�<OE�<���<L��<;�<�O�<���<}��<\��<e2�<Ia�<���<���<m��<+��<H��<���<�@�<���<�Q�<��<���<�*�<�U�<�|�<Ĥ�<���<��<�H�<��<���<�0�<��<iǽ<G�<�,�<D�<�G�<�9�<��<y�<���<i��<�W�<�"�<&�<J��<*��<�X�<O)�<���<�ԗ</��<
��<�x�<�\�<�;�<��<�ڈ<��<�<�<�ց<+�~<W�y<��t<�p<�7k<
�f<vb<׬]<~Y<�uU<��Q<��M<��I< F<DB<VQ><[B:<�6<��1<�q-<�)<۔$< " <a�<�H<k�<��<�+
<V�<؊<���;D*�;f��;���;8��;Mr�;dK�; 	�;B��;|�;�M�;�s�;쐕;&��;��;�~w;h�g;I�X;ƕJ;��=;C�1;�';�';��;�7;=�;?�:��:�~�:o
�:���:Uo�:ǩ�:g�:7 l:��P:7:4�:g�:3��9�3�9���9�aQ9Qu9ɘ�8�m�	@��[��@V��������W��I��"*�&�E�Q�`�U�{�4z������z������E���Է��p��Kmº�*Ǻ�̺tѺ7�׺~�޺W纫<�&3���W�ƹ�=!�Qz�������!���&���+��0��n5� :���>�5%C��G�$!L�c�P�T�U�Pl[�$la��g���n�� v���}��r��(��
\���o��y0������ױ��{����������T����  �  n�=��=BN==	=B�=�g=�=��=�O=�� =v� =�5 =���<��<�g�<���<�+�<���<>�<�|�<���<�l�<0��<CK�<ө�<���<�9�<�j�<h��<���<.��<���<��<�M�<���<���<b�<���<Dt�<d�<���<�T�<��<��<��<�z�<���<�/�<Vv�<���<���<0'�<`�<���<P��<^�<�T�<3��<"��<N
�<�B�<�u�<���<���<���<	��<ș�<�U�<��<�p�<��<W!�<�]�<͏�<���<+��<7�<,O�<8��<���<b�<�b�<���<z�< �<�E�<LX�<DW�<�C�<\�<~�<崭<�v�<y7�<H��<���<��<yP�<��<��<EΙ<���<]��<���<ln�<mZ�<�@�<T�<�<��<�U�<Y��<�<-2z<�Ou<�xp<̶k<�g<��b<�4^<��Y<��U<��Q<�N<�;J<�aF<szB<�}><;e:</6<_�1<�q-<��(<�q$<c�<h<N�<�y<�<ϴ	<�c<!<K��;m��;�r�;"g�;�j�;�m�;�`�;s3�;�ݸ;�[�;���;��;�&�;Hq�;��;�Ny;��i;d�Z;�L;�?;��3;��(;�;�5;�J;��;k��:��:,^�:���:�ֳ:15�:��::-�:�Ih:��K:	1:7�:=T :GG�9��9�P�9�=9
��8w�W8_������`�фQ�)��\帹&�������%�Q@���Z� �t�.���1���99���K��4��Q�����Vz���ĺO�ɺ�Ϻ�;ֺ(�ݺx9������y��v,�������<��k�4�#�.�(���-��N2�,�6��H;��?���C�:�G��*L���P���U�?�Z���`�J!g���m���t�R(|�h���f��5_��Ud��g����������ꖔ��G��Vؗ��_���  �  �=Η=�W=�=	�=�h=�
=.�=KC=!� =�z =� =Nz�<}��<�!�<I��<���< a�<���<�[�<���<&`�<���< N�<���<��<fM�<܄�<t��<���<"��<g&�<OX�<:��<���<�?�<���<#)�<Ų�<UF�<���<�y�<��<���<��<��<l��<�.�<�m�< ��<���<q �<P/�<Sa�<Y��<{��<��<�P�<B��<q��<9�<fY�<���<��<5��<M��<��<�g�<�	�<	��<*��<P�<���<+��<v�<f6�<:i�<��<���<h�<W�<���<�׿<5�<�=�<�\�<�i�<c�<CI�<��<��<{��<�X�<A�<�Ŧ<-��<�B�<�
�<۝<���< ��<�~�<
p�<f�<�]�<|R�<@�<3"�<���<!��<�l�<[�</`<��z<ſu<��p<�El<L�g<�,c<��^<��Z<VqV<�jR<rwN<��J<H�F<=�B<3�><}�:<�?6<`�1<�f-<��(<�@$<3�<<"{<��<
�<�%	<��<ՠ <���;���;���;��;�-�;�Q�;�`�;]L�;��;��;�;�j�;�;c0�; ˅;[S{;��k;��\;O;��A;�5;9�*;�I ;��;Cc;��;�:��: �:B��:���:���:LÑ:8c�:�\c:�E:	�):�:yK�9I��9[ �9��h9ܹ#9#V�8~$8�˚�gМ�kM�`!O�Y��*ᴹ�.��Z��J!�[�:��AT��m��S��V���i������+����ׯ�AT��K���º��Ǻ�
κ��Ժ]�ܺ���)���J��3����@����4���S �0�%�$�*�"�/�AN4�פ8��<���@���D��`H��aL�	�P�c[U���Z��7`�pbf���l���s�
�z��ƀ�����C��U6���ꌻ2_��씑�ƒ��ld��c�� ��  �  ��=��=�]=	=S�=�e=2=P�={3=�� =�_ =���<P3�<�}�<h��<:8�<Z��<�#�<Ȩ�<�3�<H��<sL�<���<�I�<���<��<�[�<��<���<���<.�<oa�<I��<P��<>2�<���<%��<�p�<���<�{�<
�<$��<�'�<ѫ�<#�<���<��<�&�<^�<��<���<~��<���<v�<�N�<���<���<��<�Q�<E��<���<�5�<�u�<���<���<���<ū�<Gs�<p�<4��<+�<�|�<���<W�<*N�<���<V��<���<�'�<�^�<t��<���<��<�1�<�V�<`n�<�t�<,h�<%H�<��<ԯ<���<n3�<�ݨ<���<4=�<l��<̽�<͎�<�k�<cT�<�G�<kC�<BD�<�E�<�C�<�8�<!�<|��</Ć<�~�<Z-�<զ<��z<o/v<�|q<��l<nHh<��c<Rn_<�&[<r�V<��R<��N<+�J<H�F<>�B<&�><�:<C6<��1<�M-<��(<`$<~N<�<��<�g<��<��<V><� <,��;!�;f9�;n��;��;��;�D�;�H�;!!�;ϰ;�[�;�֟;U�;��;.��;ha};Pn;UY_;�rQ;�ZD;�8;��,;�!;j�;5b;�O;���:���:�5�:��:�)�:��:0'�:�K~:f�]:�t>:Nd!:��:w�9��9ꎇ9]IG9�9��8}�7]������ۨ��0P�b`���m��ݹ�`��;��5�[�M��Fe���{�d����k��i���I䣺񉫺咲�0)��f�����źɩ̺�Ժ�?ܺy�ѹﺦ����v��	����f� ���y"�(��C-��2���6���:��t>�B�L�E�RI�v�L�,�P��[U��YZ�=�_�E�e�4l���r�OCy�������������G����$��+n��B���񀔻�]��"/���  �  w�=ӧ=}`=�=�=<_=6�=U�=� =B� =2C =��<E��<�.�<S��<"��<�_�<E��<�q�<��<%��<\2�<g��<9>�<��<"�<Mb�<^��<=��<2 �<iZ�<q��<���<_)�<�~�<���<�D�<ڴ�<l-�<���<>1�<ڶ�<�9�<���<9&�<���<K��<��<�G�<Bk�<*��<��<V��<\��<��<�5�<ys�<���<,�<>b�<���<$�<�V�<`��<G��<ڽ�<��<�w�<�'�<���<K:�<���<���<�N�<���<���<��<�A�<�s�<p��<���<���<�(�< M�<i�<�x�<�x�<�e�<�?�<p�<׼�<�f�<	�<��<�K�<��<0��<�m�<�?�<� �<F�<n�<�<��<�'�<�-�<�)�<q�<���<�ǆ<ى�<A�<��<�;{<��v<h�q<jem<��h<ikd<�`<۶[<�xW<LS<�.O<fK<�
G<�B<e�><d�:<A76<��1<�&-<!w(<��#<#�<�*<{s<��<�I<��<��<���;���;_ �;�y�;K��;_�;t��;�
�;}'�;��;�߰;���;3*�;ї;蒏;.��;�T;�2p;f�a;t�S;��F;S&:;�h.;7a#;�;~2;��;���:��:���:7�:�%�:�:�+�:�#y:�W:!�6:��:�9�
�9���9�h9$9N��8� H8��/4��A�YŸ�����T��G��Ա�!�ڹb;����}�0�_�G�l�]�nfs�%ꃺŚ��þ��Y��Lp�����HQ��Z[���fĺ%�˺��Ӻ�.ܺ���h�'	��;@���
��q�6�����$�Xz*�2�/���4���8�%�<�|H@�i�C�_�F���I��vM�LLQ��U�!fZ���_�koe��{k��q�_�w��3~����Z��Ї�u�������S��Ï��H������鲗��  �  ��=��=�_=�=8�=�U=��=r=�=� =�& =�p�<s��<���<)7�<ў�<8�<{��<6:�<X��<"x�<@�<��<�,�<ܢ�<�	�<b�<���<w��<j:�<x�<��<��<�i�<X��<�"�<"��<���<�a�<���<;P�<d��<	E�<���<{"�<�}�<+��<��<�,�<�H�<�\�<�l�<P~�<Ɩ�<���<<��<�&�<�q�<,��<�%�<��<C��<d4�<�u�<��<���<-��<�t�<�+�<��<P�<���<�*�<s��<X��<��<.U�<���<���<���<��<�'�<�F�<7a�<t�<�{�<#u�<�\�<�0�<��<\��<8C�<�ܪ<�s�<��<ᰣ<�`�<� �<�<�ך<y͘<oі<�ߔ<�<�<��<!�<x	�<z�<�Ć<֍�<�M�<f�<\~{<�v<Eer<��m<ii<��d<)�`<(7\<y�W<��S<�vO<NK<�)G<�C<��><Ѓ:<_6<��1<�,<�7(<�f#<w�<ܶ<��<�><خ<�D<�<���; ��;�8�;$��;�G�;���;�[�;��;���;��;3հ;���;�a�;&1�;��;=7�;���;�$r;��c;��U;��H;�;;��/;[�$;��;\�;
";	��:�c�:�D�:�:gʰ:�^�:���:'�s:$�P:�</:v':M��9�ɴ9�B�9��C9��9�p�8gŽ7�έ�,5��j��s#���\��ᎹQ�9GڹS��&{�|,-�^�B��W���k����RB��0n���J��У�e���쳺󤻺Rú;2˺�Ӻ|�ܺ����w�Vv���*�d��������� �+�&���,�--2�W�6�-%;�.�>��B�E�"H��K��CN��Q��V�H�Z���_�Je��k�4q�@�v���|��F����������]���勻�W��H�������+��eS���  �  {�=��=Y\=�=խ=K=��=wo=�� =l� =t =�5�<~a�<���<���<&\�<G��<%j�<��<���<VS�<���<���<>�<��<���<�\�<V��<> �<iM�<��<*��<�D�<��<p��<f\�<���<T#�<���<���<�g�<:��</J�<r��<��<]p�<ݶ�<���<~�<'�<4�<$=�< H�<>Z�<ux�<���<*��<�0�<S��<��<%V�<���<��<�Y�<���<��<k��<Xm�<t*�<��<�^�<?��<�L�<��<��<�Q�<n��<���<��<��<U/�<#H�<l]�<bn�<�x�<�y�<�l�<WO�<��<�ڱ<���<� �<6��<�B�<֥<s�<��<�ܞ<���<��<���<ݛ�<���<3˒<��<���<O��<O��<�<���<z��<T�<��<�{<15w<��r<BJn<��i<-ne<	a<6�\<zEX<�S<[�O<jrK<$<G<.C<q�><�m:<h�5<'p1<&�,<n�'<#<q2<_M<�w<��<�%<P�<z<��;z��;Ae�;���;'��;�W�;���;{_�;ؤ�;e��;鷰;/��;M��;�u�;���;}Ȉ;�9�;5�s;}e;�W;�QJ;;=; @1;�%;ܛ;j.;.A;Qh�:���:4[�:w��:N�:Ɛ�:Sщ:�n:ܝJ:�a(:~�:�'�9���9�en9��"9$�8�M68�I ���)�u�.���r;/�)Lf�Cm���@���۹p�A��9f*�{�>�1xR��e�´x�����َ�>헺٠�������d��~�ºI
˺��Ӻ�2ݺ"t纍��, ��;�%��5��Y�K"�h�(���.��N4�<9��(=���@�B�C�$�F��=I��L��O�\�R��V��[�� `�[Pe��j�6�p�"(v���{�K���xB��ᅻAv�������������h����������  �  �=&�=IX=n=��=JA=��=�a=�� =�o =���<C�<�.�<�j�<H��<�'�<n��<{<�<���<���<�4�</��<[w�<T�<ă�< ��<�U�<¯�<�<�Y�<���<�	�<�f�<��<'�<���<���<2H�<[��<+�<w�<8��<UK�<���<N�<�b�<���<<��<��<n
�<��<��<��<@*�<E�<|p�<���<��<[�<X��<k/�<I��<��<�A�<Pu�<��<j��<dd�<o&�<���<�g�<���<Be�<���<�,�<�|�<z��<|��<�<�7�<�M�<�^�<Ml�<�u�<�y�<�t�<sc�<�A�<��<Ʊ<(l�<r�<��<X�<���< B�<��<W��<mz�<d�<b�<�p�<���<O��<Ȑ<�ގ<��<�<�ӈ<���<���<VV�<f �<Q�{<�gw<z�r<��n<�/j<��e<�Za<��\<�X<�)T<��O<@�K<�DG<2 C<ճ><RV:<C�5<�I1<d�,<�'<��"<9�<��<�<�U<�
<�K<i<��;x<�;%��;�g�;�)�;K��;q��;��;�`�;���;t��;���;���;Q��;�Ӑ;�1�;۽�;d�t;(�f;�X;��K;��>;-2;�P&;�;Af;�B;V�:!"�:u�:���:���:���:���:k]j:4�E:��":pz:�:�9c�9�S9��9�o�8&ֻ7#���m�W*ĸ]��9��0o��򕹓ʷ�$cܹ�a�%���(�D�;�޷N��Ba�L�s������+��dl������F˧��Ű�y����Lº�˺85Ժ��ݺ�b�"��/ ����U��N�A��e�#�2f*���0���5���:�w�>��(B�;E���G�@J���L�x�O��7S��W�/u[�/F`��le���j�>5p���u�r�z�b��h���>9��Rɇ��Z���팻-|��� ��Dy���喻�  �  ��=��=U=��=�=n:=�=�X=F� =�c =���<4��<��<�H�<��<�<���<�<(��<qq�< �<P��<�g�<��<�x�<l��<P�<���<�<=`�<���<a�<�{�<���<cA�<1��<�<�^�<��<�<��<>��<�J�<���<��<�X�<B��<���<X��<��<���<���<] �<u�<D$�<N�<���<+��<!<�<��<5�<��<���<1�<-g�<-��<�}�<g]�<�"�<���<l�<���<�s�<���<_D�<��<Q��<(�<�3�<2N�<`�<`l�<�t�<}y�<y�<�p�<\�<8�<��<ŷ�<Y[�<��<^z�<��<���<�"�<\ɠ<-��<yX�<MC�<�C�<U�<r�<K��<ݴ�<Ύ<0ی<�ي<�Ɉ<g��<˄�<�V�<Z%�<H�{<��w<�%s<��n<�cj< �e<��a<A ]<N�X<$JT<�O<��K<�GG<F�B<��><�D:<��5<�.1<�t,<Z�'<�"<��<��<	�<I<u
<�<��<�~�;���;�L�;J�;���;h��;OK�;���;�/�;�c�;�z�;��;В�;w��;���;lp�;U�;�u;��g;�Y;�VL;KK?;ʻ2;Q�&;�Q;\�;z:;��:L��:���:k��:�
�:[�:�Æ:όg:��B:7X:~2�9���9�ԍ9�}B9�=�8�xl8��7��"o��O�׸���,,A�ruu�����A����ݹ�~����R�'�J,:��uL�}|^�up��L��!���1㓺LS�����-��} ��%º>5˺-�Ժ�i޺W麤���4� �"w����j��m���$�;c+�E�1�\7���;���?�~C���E��{H���J�}M��YP�U�S�JuW���[�d|`�	�e���j��p��Mu��yz�[��;M��^҄��^��+�K���,�����N���ϖ��  �  N=R�=5h=�=U�=eH=�=�S=�� =FB =r�<�l�<�|�<{��<��<�l�<q �<��<�s�<�B�<��<��<��<m/�<K��<�0�<���<���<�P�<���<��<�|�<���<XY�<���<*�<ވ�<���<�;�<a��<���<�\�<���<�/�<���<
��<�'�<�Q�<�c�<Ua�<9P�<�8�<�$�<�<?*�<^R�<��<>��<v�<��<��<d.�<���<t%�<�v�<���<c��<g��<�Z�<
�<Z��<%4�<���<d*�<��<���<M#�<xM�<[d�<l�<�i�<�b�<�Z�<\S�<EJ�<6;�<Y �<��<
��<O�<0ׯ<5J�<8��<i�<+u�<��</x�<u$�<A�<��<��<4�<jL�<���<���<��<u
�<a�<��<��<E��<͇�<1U�<9J|<��w<��s<pDo<��j<Xwf<��a<�r]<y�X<5aT<b�O<_�K< (G<E�B<s�><�:<��5<!�0<��+<��&<��!<��<�C<�<5<�K<��<��;��;E��;Bm�;ل�;1��;���;۲�;t]�;E��;��;�٭;���;���;˶�;��;�a�;c~;�o;r^a;�\S;P�E;@8;z+;;�;R ;o;��:�'�:�c�:���:{�:�:O�:pzi:Z�@:Y:X8�9dk�97E9�%�8/�6��h���ҸzZ
��0!�[A3���E�y`]��s}�^��I����ι���
���r/��?@��P��"a���q��d��]m���哺�����w������p��ntúyV̺hպߺ̴麙������������}1���!���)��1�\�7��i=�B�?�E��/H�$ J�*�K��M�ձN�t�P���S��V�[���_���d��j��So�Pht��Oy�~��e���̃�GJ���䈻�����S�����j����G���  �  �=�=�j=�=ʵ=>L=R�=sX=� =)H =Z�<�z�<d��<���<w
�<�|�<��<G��<��<N�<�<J��<X��<�6�<���<�6�<;��<}��<�Q�<��<P�<�u�<���<uN�<۸�<�<g}�<���<�3�<��<���<K\�<���<�3�<���<V��<./�<�Y�<~l�<#k�<"[�<E�<(2�<�+�<:�<�b�<$��<$
�<τ�<N�<_��<Q9�<Q��<7.�<�~�<���<}��<O��<�^�<��<ѥ�<"1�<���<="�<�<��<��<A�<�X�<b�<b�<�]�<ZX�<PS�<{L�< ?�<e%�<��<��<�V�<�߯<T�<Q��<��<"��<���<;��<�4�<��<��<���<�#�<�X�<���<fː<���<r�<��<�	�<��<���<t��<_T�<NC|<��w<��s<a/o<)�j<�^f<��a<*]]<��X< TT<A�O<�}K<	*G<��B<��><N&:<+�5<<�0<�,<�'<��!<��<w^<6<�5<�l<_�<�G�;aM�;��;��;´�;h��;S��;���;^}�;�ܽ;8��;��;x˥;Q��;���;��;(H�;L�};�>o;�a;��R;@:E;��7;��*;,�;��;�;x��:wj�:��:�6�:�|�:�D�:���:��j:�@B:�:���9&!�9��L9k{�8ot7��H���ø�n�#���-���@��X��ly��.�����{�̹���9l
�?�AY/�<�@���Q�\]b�!s��$��1+�� ���n<���觺�e��`����lú+̺�!պ�޺eK��3���I����=������!!��')��0�h?7���<� �A�PE�y�G��I��EK�\�L��eN�7�P��DS��V���Z���_��d�nj��Zo�5�t��y�vU~�����Y����z���������zv��'���œ�8L���  �  ;
=&�=q=�=F�=�V=4�=�e=�� =Y =P��<��<���<��<M:�<���<6<�<`��<��<�n�<.9�<"��<z��<�K�<p��<$F�<6��<���<�R�<p��<	�<%a�<D��<�-�<6��<���<[�<��<��<O��<���<�Z�<E��<�=�<���<���<�B�<�o�<��<���<?z�<h�<vY�<�V�<h�<$��<���<R8�<���<�8�<���<rX�<���<�F�<��<þ�<:��<֥�<�g�<��<���<�'�<���<�	�<�f�<���<���<��<6�<bD�<�J�<�M�<YP�<=R�<Q�<9I�<P3�<�	�<Tȴ<�l�<���<�o�<�٪<�?�<R��<�%�<޶�<�d�<2�<G�<?)�<�J�<.{�<p��<��<.�<�(�<\,�<!�<i��<7Ƅ<���<UQ�<-.|<'�w<�Ws<��n<��j<�f<V�a<�]< �X<g,T<��O<�sK<�-G<��B<У><�E:<�5<�1<�>,<]:'<�"<o�<�<�<c�<��< G<E <U�;�s�;`<�;�=�;�T�;~\�;<8�;���;*,�;�?�;�"�;��;���;͟�;��;���;��|;vBn;��_;t�Q;�/D;��6;�%*;?
;	�;I;��:S�:���:ZU�:p��:⫞:@�:7n:0F:s:��9c�95$d9sM�8x�8�׷�w���޸�'	����>�2��lL��Ln��0�������"ɹ�<�U�	�:�m\0�#�B�ǪT�3f�kKw�th��i��S���`���p@���G��h����eúx�˺�iԺ�ݺ�(躨��t� �n����i�����,�'��:/���5��g;�6@�%�C�iF���H�Q4J���K���M���O��R�\"V�@`Z�i7_�yd���i�sto�_�t��z����������d������@?��tގ�Is����C\���  �  �
=�=iy=�'=C�=�e=;�=y=6� =�r =D��<���<���<�3�<��<���<S��<�&�<S��<���<:d�<� �<���<�h�<���<	[�<���<��<�Q�<���<���<D>�<��<���<u[�<"��<�#�<؉�<��<�c�<���<�T�<|��<!J�<]��<��<^�<���<���<��<Ũ�<`��<���<a��<k��<H��<�!�<��<���<cu�<.��<��<�<�i�<ò�<E��<���<���<es�<S�</��<��<G��<���<U4�< {�<߳�<���<���<��<9$�<�2�<�@�<�M�<VV�<�U�<�E�<� �<�<���<��<���<�	�<�v�<�<�i�<:��<5��</|�<Af�<'k�< ��<ͯ�<x��<�<�3�<�G�<�G�<R2�<�	�<ф<���<�I�<�|<ׁw<�s<W�n<Cj<�e<\'a<=�\<�GX<!�S<��O<�^K<<-G<��B<�><vo:<V�5<,S1<ʁ,<T�'<�n"</F< <�<�<�b	<��<� <� �;y�;�&�;;�;/
�;��;���;�R�;a��;���;sh�;�;N��;x�;3\�;Zu�;�{;ݦl;�,^;�P;�B;�i5;��(;u1;!/;�;j�:H��:r��:l��:Ԃ�:}��:?V�:�Xs:�L:��%:�]:*��9��9�r!9�"�8T�7H�)�nҡ��ܸR3��5��c:��m^�A��j���yPĹ��鹍	����O2��EF��{Y��l��+~�����	�����pࢺ����Fѳ�(Ȼ��ú�P˺�Ӻ>{ܺ�溣#�������$\��L��?���%�-�+�3�<9�h�=��oA��]D���F���H�M`J�^TL�ưN��Q�
OU�_�Y���^��#d��i���o��tu�H
{��7���ւ�i��4�����������������@F��U����  �  �=A�=��=D2=��=�u=�='�=Z=p� =b =r6�<VX�<F��<'��<~Q�<m��<�u�<�#�<��<���<UK�<���<N��<&�<�n�<���<��<�J�<t��<6��<7�<[�<���<��<]p�<���<G�<��<�:�<]��<TH�<��<tS�<d��<-�<xz�<D��<��<���< ��<=��<'��<���<�	�<t:�<M��<���<G�<}��<�@�<���<�1�<���<���<���<���<e��<�{�<��<n��<K��<�V�<%��<j��<m-�<�a�<c��<���<���<?��<;�<�'�<KB�<pV�<�^�<
V�<7�<���<Ϭ�<�C�<�ȭ<�B�<���<�5�<"��<[�<�<5ڜ<���<���<mϖ<��<��<Q=�<[�<ni�<)d�<LI�<�<�ل<Z��<n:�<��{<%)w<�r<]�m<zi<��d<@�`<�$\<��W<�S<�YO<9K<�!G<XC<��><`�:<�*6<C�1<��,<(�'<.�"<n�<��<ѱ<��<|!
<�<�W</��;���;�G�;]�;���;���;Ib�;��;�;���;��;K0�;۪�;�0�;bی;U��;&�y;�zj;F�[;E�M;+8@;c3;�J';T�;Ei;��;}�:���:^�:�_�:Y[�:֢:�ݏ:�Jy:S:��-:
�
:	��99^�P9��84[8Sy��s�+�Nޙ���Ӹ/W��3&�fHM�5~�<͜��ۿ�7b繵	��+��l5�72K��.`��Bt�C���
���땺Q����Ԧ�%������$��;ĺ�˺��ҺSGۺ���A�7���.e�����x���#��c*�/�0�66�x�:���>��A��fD��F��H��J��M���P��tT�7�X�0^���c�#�i�<1p�Ibv�kl|�N��wꃻ����2��D���%���w��=����Ô��Ŗ��  �  �=O�=s�=�9=�=(�=�=}�=�+=�� =9: =ݏ�<^��<e��<	O�<���<�9�<z��<�n�<f�<I��<�s�<��<��<��<"|�<#��<��<�:�<�h�<֘�<	��<��<�Y�<ׯ�<0�<�}�<���<Ex�<?�<��<�1�<���<�T�<T��<�=�<F��<B��<���<��<��<h#�<�1�<�I�<o�<X��<]��<o@�<s��<��<U��<���<�_�<��<���<Y
�<���<���<|{�<��<�w�<`��<��<ha�<��<���<��<+�<UU�<X�<s��<2��<��<�,�<lM�<`�<7_�<�F�<��<�ɲ<�h�<���<�}�<v�<e��<h�<*¡<�x�<�C�<e$�<�<z�<]3�<�N�<|j�<N�<u��<{�<�Y�<j#�<�ل<���<P!�<�z{<��v<��q<;Vm<˿h<�<d<��_<;w[<�7W<�S< O<��J<�G<��B<�><��:<�Q6<!�1<-<�3(<�A#<�E<�M<)g<<�<��
<z|<�-<��;5(�;ۀ�;��;���;�b�;$��;
M�;Vf�;B8�;�ɮ;H+�;?u�;K;�,�;Ỹ;�ew;;�g;=�X;��J;!u=;��0;7%;�];�N;z�;u�:\��:���:��:*޶:���:8�:�&:cLZ:��6:�:I�9�>�9-�9�l19N�8<8t���&������yݸ[d��Z>�_7r��o��e'��׽�)
���!�"�9�V�Q�(�h�ZH~�Z��p蒺ZЛ����ޭ����������'���(ź�v˺3tҺ�ں���Q�������(��D�ː����a� �tb'�8d-���2�+y7�*�;�9�>���A��D��G��I�iL�?�O���S�Z�X���]���c��Yj���p�,�w�]4~��>��:���
��r���*��My�����(����n��m2���  �  ��=ο=}�=J;=��=��=m$=�=�C=�� =�` =7��<� �< g�<���<%�<��<�#�<���<U�<��<���<*�<��<"�<~�<`��<I��<)�<?�<�_�<���<���<���<�F�<��<��<��<")�<L��<�i�<~�<@��<K�<���<EC�<C��<���<��<�2�<!M�<
f�<��<ϧ�< ��<��<X�<��<��<e�<���<�,�<��<���<i�<,�<	�<���< p�<���<tT�<S��<���<�<O<�<tf�<ܐ�<���<���<�"�<\�<c��<���<�<9�<�U�<�\�<=K�< �<�ܲ<셰<
!�<´�<�G�<'ߦ<��<`,�<�<:��<s��<�u�<�n�<,t�<g��<���<随<���<��<f_�<�!�<�΄<�k�<x�<�{<
0v<Yq<��l<L�g<fec<��^<��Z<�V<��R<�N<:�J<��F<�B<��><W�:<�b6<��1<�>-<�y(<]�#<;�<��<�<�k<f�<�^<h
<ܱ�;��;���;?�;{�;!��;z\�;���;j��;�M�;8��;���;b�;�(�;)U�;#��;��t;��d;��U;t�G;r[:;_.;��";-q;��;��;���:�O�:/��:"��:���:G�:��:��:W�`:&!?:FQ:��:�s�9��9Z�h9t�9M �80!8�1綒�F��ȴ�����&4���k�Pؖ�kF����蹴f���%�ѳ?�}pY�mBr��ք����i����d��pD���3���K��i��� ���+�ƺ�̺��Һ�oں<e�/��s���9,�j�	�������� ��P$�**��O/�^4�R8�<�q|?�ÎB�xE��iH�ʘK��8O�tS�_bX�^��Md��k�a"r��Gy��'��懃����������Y���Ɏ������쒻p���dD��˗��  �  p�=��=Hz=�6=v�=��=7+=��=RW=� =� =q =y��<"��<�'�<���<4��<�u�<y��<��<��<��<`5�<���<��<s�<B��<���<���<f�<��<7�<�[�<���<���<�8�<���<w7�<���<T~�<L1�<���<<��<h5�<���<�;�<���<���<�!�<@P�<�x�<m��<���<� �<x:�<�z�<e��<"�<]]�<���<9�<NY�<���<���<��<K�<��<%��<pX�<���<�'�<g�<��<`��<���<���<]�<�K�<���<���<4�<BR�<���<��<��<?�<�M�<�B�<��<R�<e��<�@�<��<���<�-�<�ۤ<���<#Q�<�<��<�̙<���<���<z��<���<=��<���<K��<�W�<+�<f��<K�<R�<d�z<o�u<ȧp<��k<�g<��b<, ^<�Y<��U<��Q<�N<�KJ<q�F<�B<6�><>�:<2Z6<m�1<�X-<y�(<y�#<�/<\v<��<�0<�<�8<�<8�;#��;���;���;�;"^�;
��;ݱ�;ᒿ;�/�;J��;���;7��;�l�;�_�;l��;��q;��a;oR;Q7D;(7;"+;�: ;�L;b.;m�;h�:��:q�:���:z��:댦:�1�:���:K�f:�F:��(:\:2y�9-�9Oَ9�5Q9�Y9Y�8;�7J�ַ����l����0��k�1���A�����!��*���F�^b���|��܊�5D���k��@���ð�����V�����%ź�^ɺ�9κ�Ժ*ۺ%�������������� ?�D��\��2h!���&���+�%�0��D5��j9��?=���@� 3D���G��"K�~O�/�S���X���^�)
e�`l��s��#{�rP���脻FE���V��3��={��x���?S���ڕ��8��T����  �  ^�=ˢ=�l=L,=O�=E�=s,=��=Qe=�=K� =vD =��<:,�<F��<���<�N�<���<�2�< ��<�2�<s��<�5�<���<��<=]�<M��<z��<���<W��<a��<���<W �<4,�<�o�<���<=F�<���<�~�<�5�< ��<ݴ�<,m�<d�<U��<W)�<z��<���<�'�<�b�<��<Z��<J�<�N�<ݒ�<��<��<1f�<F��<���<68�<{�<���<���<-�<>�<=��<��<�7�<��<��<�(�<J�<�`�<�u�<'��<ү�<w��<w�<H`�<&��<�	�<�`�<���<��<�<�3�<D/�<R�<��<���<�U�<N�<���<r�<-�<��<9��<�w�<�D�<��<���<0ܕ<}ʓ<Ľ�<_��<�<z�<nE�<d��<���<�"�<�:<�z<	u<��o<)	k<Cf<n�a<�K]<�Y<�U<"IQ<	�M<��I<b,F<�fB<ɀ><Ts:<&;6<��1<0\-<8�(<�'$<�<I�<Aa<+�<ih<-�<G�<�H <l�;��;8��;���;��;���;��;�a�;��;,"�;��;��;қ�;^�;aQ�;�3o;�^;�5O;_�@;@�3;88(;ۤ;_;^];�4;y��:�?�:f��:ۉ�:��:n^�:���:�6�:9�j:"�L:v�0:0�: ��9Q��9%��9�~9�549��8�	D8����u��&n��1�]Iq�񜹯�ƹʦ�����C�0�Z�M��k�x����Ő�W������U᯺��+ּ�Yh���*źf�ȺE5̺(|к��պA�ܺW���I�����u3�f�f�,��8u�q���$��)��-��2��7�U;��b?��EC��G��K��>O���S�FGY�(R_�\f�9fm�g)u��}��~��'G���ˉ�k���ؿ���������������F:��~Y���  �  z�==�=4]==��=$�=�)=2�=?n=�=�� =tb =� =Ey�<0��<�3�<��<���<^�<���<~A�<���<�-�<��<���<�A�<�u�<���<2��<���<��<���< ��<���<��<�n�<;��<��<b1�<���<��<߃�<�C�<1��<���<��<�}�<���<4%�<�k�<h��<5��<}A�<_��<���<'�<�m�<���<���<�&�<	^�<R��<���<���<��<y��<^��<���<��<�{�<]��<��<e�<��<<�<U/�<�M�<�{�<���<�	�<�d�<���<�&�<�<�Ǽ<���<�<��<,��<�ղ<<ga�<�!�<��<ʨ�<�o�<�7�<���<�Ş<���<�V�<
'�<���<ߓ<,ő<ܬ�<ˏ�<g�<�,�<a܆<u�<C��<��~<ڧy<xt<iXo<Yj<��e<+�`<m�\<�jX<�{T<�P<UM<tI<��E<=B<�>><�;:<>6<z�1<dO-<V�(<wK$<#�<N<l�<�n<<4�	<�7<�� <��;�u�;�;���;���;���;ji�;��;Ă�;���;���;H;�;�Α;5j�;�l~;S�l;��[;WL;">;/'1;f�%;eJ; 
;n�	;�;�A�:�%�:'��:t�:0��:�:#��:'Ӆ:��m:S�Q:�g7:� :o:m�9�P�9Ӕ�9��T9�k
9���8��/6��m����z�6��Zz�b���͹bI��Y��I�6�yU��Ys��^������e������Ƶ������
º�
ƺ2ɺn̺�Ϻ��Һx�׺OT޺�,溳Tﺟ���3+�����1����������Ѩ!�N�&�r+��T0�;$5���9��T>���B���F��+K�*�O���T�>Z�J`��2g�A�n�
�v���~�q��������)��l��C<������x������*��/���(���  �  E�=T=dN=/=�=�z=�$=��=1s=�=� =<x =�( =}��<��<l�<<��<-�<|�<���<�H�<��<�"�<N��<��<'�<W�<4q�<�x�<
s�<�h�<�c�<@l�<���<���<1$�<���<�=�<7��<x��<���<�Y�<��<���<q�<!��<ii�<���<w�<9n�<��<Z�<f�<��<��<�`�<��<��<%�<<L�<x�<���<���<T��<v��<���<���<,f�<4��<�U�<��<3��<���<���<��<���<n �<�.�<�p�<���<&�<q��<��<{T�<��<�ٺ<���<���<��<�ǲ<���<#f�<:2�< �<:Ч<���<�n�<m9�<J��<���<��<�I�<g�<!�<�Ƒ<N��<��<�R�<*�<ￆ<OT�<�ҁ<�~<-Dy<\t<��n<f�i<��d<V`<v�[<��W<��S<jBP<b�L<bI<N�E<A�A<i><:<`�5<c�1<�;-<��(<\_$<a�<>�<?4<��<?{<�
<P�<{?<ү�;��;�e�;���;S��;�q�;�+�;#þ;� �;{8�;�
�;ܤ�;- �;���;�|;��j;��Y;�J;�;;J�.;�#;�e;�[;$;}u ;u	�:�1�:��:ܛ�:�Ǵ:�ܤ:@*�:�:wyo:p�T:�<:F�$:��:��9���9�L�95�l9Rq9WZ�8�0$7�!f��p����=�������Թ�"�,���<���Z��+z�K5���Q���禺㪱�_k���/��R1ƺk�ɺ�̺M�κ9�Ѻ�#պ��ٺkຟ�红z��A���H�9�� ��H���t��0�a��_�$�E�)���.��3���8��=�aQB��F�pK�
(P��=U��Z��3a��=h��o�5x�*F���y��5���<?������lg��P���E���c����������ٚ��  �  �=�s=�C=�=��=�t=� =��=gu=�"=�� =i� =�8 =���<>5�<֎�<���<8�<V��<���<�K�<n��<r�<�z�<6��<��<pA�<Y�<�]�<{T�<^F�<�<�<�A�<�]�<:��<\��<�r�<��<���<1��<Uj�<>=�<��<��<�\�<��<TZ�<U��<E�<n�<���<��<�{�<1��<�2�<̄�<���<��<�8�<�b�<
��<ק�<��<6��<	��<>��<^��<Q�<���<y;�<y�<��<F��<&��<��<���<���<v��<A�<���<L��<�i�<�տ<�7�<.��<Hº<��<H�<�۴<��<U��<Vg�<�:�<|�<��<\��<7��<�]�<�"�<>�<~��<�^�<�#�<��<�ő<���<nu�<�C�<�<���<f=�<+��<EE~<=y<Իs<��n<ysi<�d<_�_<��[<1�W<�S<m�O<�cL<Q�H<LE<��A<��=<��9<�5<R�1<D+-<�(<Bh$<� <�<j<<{�<�a
<�<�<��;�E�;l��;S�;��;WS�;���;���;2ٵ;y�;��;�=�;Ȫ�;��;�u{;�hi;aX;=�H;�P:;��-;R,";�);�@;�);�/�:���:,��:���:���:�߳:�0�:�Δ:��:_p:!�V:�>:�s(:�:��9��9���9�M{9��(9Ͳ8m�a7x�d�������B�7���V`��d�ٹ�����!���?���^�u�~�𵎺S��Щ�����oe���ĺ3�Ⱥ�;̺��κ��к�SӺ?�ֺ=ۺ{>��躤X������j�Wq�[�	�Q��/?������#��(��-���2��8�99=��'B�
�F�E�K���P�;�U��u[�P�a�E�h�2�p�y�aʀ����q(����oM���&��ow��dD��B����������P���  �  i�=Jo=@=T=�=?r=/=4�=
v=�$=� =͉ =�= =u��<bA�<t��<S��<e@�<1��<6��<|L�<���<��<�u�<��<��<�9�<PP�<�S�<�I�<]:�<a/�<(3�<ON�<���<���<�b�<��<���<|��<	_�<3�<m��<��<eU�<���<�T�<��<��<�m�<���<�#�<��<���<�=�<���<���<��<�B�<j�<���<��<���<���<���<���<���<wI�<L��<2�<o�<t��<D��<���<e��<��<��<���<�0�<���<#��<B]�<$ʿ<M-�<�~�<Ṻ<V۸<��<[ִ<Ḳ<��<�g�<�=�<��<��<`ȥ<���<�i�<�.�<�<���<|e�<%(�<��<ő<���<
q�<'>�<���<-��<.5�<��<�0~<(�x<��s<in<�Ti<>td<O�_<�x[<�aW<ʆS<��O<�KL<��H<�8E<&�A<,�=<~�9<�5<�w1<�$-<��(<�j$<� <��<�{<�/<��<�z
<<�<<�;_�;���;b�;k��;�F�;���;�n�;Ծ�;�ɬ;���;��;���;`�;A{;��h;��W;!H;��9;�-;��!;ͻ;��;�;��:���:]T�:Nm�:� �:닳:J�:���:�	�:�p:HAW:��?:̥):Cn::	�9��9���9��9#�,9�߷8cau7%�d��H��pE����������۹�����"���@��Z`����^���]���SЪ�
����i��yź��ɺyͺirϺF�Ѻ�ӺK8׺�ۺ���麗��{��/z�km��B�p��s����z��4#��*(�rU-���2�}�7�=�?B�'�F���K�y�P���U�ī[��b�;i�:q�Yy������B���a��C/��5���5h��_�������٘�mܙ������y���  �  �=�s=�C=�=��=�t=� =��=gu=�"=�� =i� =�8 =���<>5�<֎�<���<8�<V��<���<�K�<n��<r�<�z�<6��<��<pA�<Y�<�]�<{T�<^F�<�<�<�A�<�]�<:��<\��<�r�<��<���<1��<Uj�<>=�<��<��<�\�<��<TZ�<U��<E�<n�<���<��<�{�<1��<�2�<̄�<���<��<�8�<�b�<
��<ק�<��<6��<	��<>��<^��<Q�<���<y;�<�y�<��<F��<&��<��<���<���<v��<A�<���<M��<�i�<�տ<�7�</��<Iº<��<I�<�۴<��<V��<Vg�<�:�<|�<��<]��<8��<�]�<�"�<>�<}��<�^�<�#�<��<�ő<���<mu�<�C�<�<���<e=�<*��<CE~<;y<ӻs<��n<ysi<�d<_�_<��[<1�W<�S<n�O<�cL<S�H<LE<��A<��=<��9<�5<T�1<F+-<�(<Dh$<� <�<j<<{�<�a
<�<�<��;�E�;h��;O�;��;RS�;���;|��;-ٵ;t�;��;�=�;Ī�;��;�u{;�hi;	aX;8�H;�P:;��-;O,";�);�@;�);�/�:���:*��:���:���:�߳:�0�:�Δ:��:_p:!�V:�>:�s(:�:��9��9���9�M{9��(9Ͳ8n�a7x�d�������B�7���V`��d�ٹ�����!���?���^�u�~�𵎺S��Щ�����oe���ĺ3�Ⱥ�;̺��κ��к�SӺ?�ֺ=ۺ{>��躤X������j�Wq�[�	�Q��/?������#��(��-���2��8�99=��'B�
�F�E�K���P�;�U��u[�P�a�E�h�2�p�y�aʀ����q(����oM���&��ow��dD��B����������P���  �  E�=T=dN=/=�=�z=�$=��=1s=�=� =<x =�( =}��<��<l�<<��<-�<|�<���<�H�<��<�"�<N��<��<'�<W�<4q�<�x�<
s�<�h�<�c�<@l�<���<���<1$�<���<�=�<7��<x��<���<�Y�<��<���<q�<!��<ii�<���<w�<9n�<��<Z�<f�<��<��<�`�<��<��<%�<<L�<x�<���<���<U��<v��<���<���<,f�<4��<�U�<��<4��<���<���<��<���<o �<�.�<�p�<���<&�<s��<��<~T�<"��<�ٺ<���<���<��<�ǲ<���<$f�<<2�< �<;Ч<���<�n�<m9�<I��<���<��<�I�<f�<�<�Ƒ<L��<��<�R�<(�<�<MT�<�ҁ<�~<*Dy<Yt<��n<d�i<��d<V`<w�[<��W<��S<mBP<e�L<eI<Q�E<E�A<m><�:<e�5<g�1<�;-<��(<__$<d�<A�<A4<��<@{<�
<O�<z?<ί�;z��;�e�;���;K��;�q�;�+�;þ;� �;r8�;�
�;Ӥ�;% �;���;�|;v�j;��Y;�J;��;;C�.;��#;�e;�[;$;zu ;p	�:�1�:��:ڛ�:�Ǵ:�ܤ:?*�:�:vyo:o�T:�<:F�$:��:��9���9�L�95�l9Rq9WZ�8�0$7�!f��p����=�������Թ�"�,���<���Z��+z�K5���Q���禺㪱�_k���/��R1ƺk�ɺ�̺M�κ9�Ѻ�#պ��ٺkຟ�红z��A���H�9�� ��H���t��0�a��_�$�E�)���.��3���8��=�aQB��F�pK�
(P��=U��Z��3a��=h��o�5x�*F���y��5���<?������lg��P���E���c����������ٚ��  �  z�==�=4]==��=$�=�)=2�=?n=�=�� =tb =� =Ey�<0��<�3�<��<���<^�<���<~A�<���<�-�<��<���<�A�<�u�<���<2��<���<��<���< ��<���<��<�n�<;��<��<b1�<���<��<߃�<�C�<1��<���<��<�}�<���<4%�<�k�<h��<5��<}A�<_��<���<'�<�m�<���<���<�&�<	^�<S��<���<���<��<y��<^��<���<��<�{�<]��<��<f�<��<=�<V/�<�M�<�{�<���<�	�<�d�<��<�&�<�<�Ǽ<���<�<��</��<�ղ<�<ja�< "�< �<̨�<�o�<�7�<���<�Ş<���<�V�<'�<���<ߓ<)ő<٬�<ȏ�<g�<�,�<^܆<u�<@��<��~<էy<xt<gXo<Yj<��e<+�`<n�\<�jX<�{T<�P<YM<tI<��E<CB<�>><�;:<D6<��1<jO-<[�(<|K$<(�<"N<n�<�n<<4�	<�7<�� <��;�u�;�;���;}��;���;]i�;s�;���;驭;u��;;;�;�Α;*j�;�l~;A�l;��[;�VL;>;$'1;]�%;]J;
;i�	;�;�A�:�%�:#��:q�:.��:�:"��:&Ӆ:��m:R�Q:�g7:� :n:m�9�P�9Ӕ�9��T9�k
9���8��/6��m����z�6��Zz�b���͹bI��Y��I�6�yU��Ys��^������e������Ƶ������
º�
ƺ2ɺn̺�Ϻ��Һx�׺OT޺�,溳Tﺟ���3+�����1����������Ѩ!�N�&�r+��T0�;$5���9��T>���B���F��+K�*�O���T�>Z�J`��2g�A�n�
�v���~�q��������)��l��C<������x������*��/���(���  �  ^�=ˢ=�l=L,=O�=E�=s,=��=Qe=�=K� =vD =��<:,�<F��<���<�N�<���<�2�< ��<�2�<s��<�5�<���<��<=]�<M��<z��<���<W��<a��<���<W �<4,�<�o�<���<=F�<���<�~�<�5�< ��<ݴ�<,m�<d�<U��<W)�<z��<���<�'�<�b�<��<Z��<J�<�N�<ݒ�<��<��<1f�<F��<���<68�<{�<���<���<-�<>�<=��<��<�7�<��<��<�(�<J�<�`�<�u�<)��<ԯ�<y��<y�<K`�<)��<�	�<�`�<���<��<�<�3�<H/�<U�<��<��<�U�<Q�<���<r�<-�<��<9��<�w�<�D�<��<���<.ܕ<zʓ<���<\��<<z�<jE�<`��<���<�"�<�:<�z<u<��o<'	k<Cf<n�a<�K]<�Y<�U<&IQ<�M<�I<i,F<�fB<Ѐ><[s:<.;6<��1<7\-<>�(<�'$<�<M�<Ea<-�<jh<-�<F�<�H <f�;ٻ�;.��;��;��;��;��;�a�;��;"�;��;��;ě�;^�;TQ�;�3o;��^;�5O;P�@;3�3;-8(;Ҥ;W;X];�4;q��:�?�:b��:؉�:��:l^�:���:�6�:7�j:!�L:v�0:0�: ��9P��9%��9�~9�549��8�	D8����u��%n��1�\Iq�񜹯�ƹʦ�����C�0�Z�M��k�x����Ő�W������U᯺��+ּ�Yh���*źf�ȺE5̺(|к��պA�ܺW���I�����u3�f�f�,��8u�q���$��)��-��2��7�U;��b?��EC��G��K��>O���S�FGY�(R_�\f�9fm�g)u��}��~��'G���ˉ�k���ؿ���������������F:��~Y���  �  p�=��=Hz=�6=v�=��=7+=��=RW=� =� =q =y��<"��<�'�<���<4��<�u�<y��<��<��<��<`5�<���<��<s�<B��<���<���<f�<��<7�<�[�<���<���<�8�<���<w7�<���<T~�<L1�<���<<��<h5�<���<�;�<���<���<�!�<@P�<�x�<m��<���<� �<x:�<�z�<e��<"�<]]�<���<9�<NY�<���<���<��<K�<��<&��<pX�<���<�'�<g�<��<a��<���<���<_�<�K�<���<���<7�<FR�<���<��<��<?�<�M�<�B�<��<V�<h��<�@�<��<���<�-�<�ۤ< ��<#Q�<�<��<�̙<���<}��<w��<���<9��<���<G��<�W�<&�<b��<K�<K�<^�z<j�u<ħp<��k<�g<��b<- ^<!�Y<��U<��Q<�N<�KJ<x�F<!�B<?�><F�:<;Z6<u�1<�X-<��(<��#<�/<av<��<�0<�<�8<�<8�;��;���;���;r�;^�;���;˱�;ϒ�;�/�;8��;���;&��;}l�;�_�;^��;��q;�a;�nR;@7D;7;�!+;�: ;�L;[.;h�;`�:��:l�:���:w��:錦:�1�:���:I�f:�F:��(:[:1y�9-�9Oَ9�5Q9�Y9Y�8;�7I�ַ����l����0��k�1���A�����!��*���F�^b���|��܊�5D���k��@���ð�����V�����%ź�^ɺ�9κ�Ժ*ۺ%�������������� ?�D��\��2h!���&���+�%�0��D5��j9��?=���@� 3D���G��"K�~O�/�S���X���^�)
e�`l��s��#{�rP���脻FE���V��3��={��x���?S���ڕ��8��T����  �  ��=ο=}�=J;=��=��=m$=�=�C=�� =�` =7��<� �< g�<���<%�<��<�#�<���<U�<��<���<*�<��<"�<~�<`��<I��<)�<?�<�_�<���<���<���<�F�<��<��<��<")�<L��<�i�<~�<@��<K�<���<EC�<C��<���<��<�2�<!M�<
f�<��<ϧ�< ��<��<X�<��<��<e�<���<�,�<��<���<j�<,�<	�<���< p�<���<tT�<T��<���<�<P<�<vf�<ސ�<���<���<�"�< \�<g��<���<�<9�<�U�<�\�<BK�< �<�ܲ<���<!�<Ŵ�<�G�<*ߦ<��<a,�<�<:��<q��<�u�<�n�<)t�<d��<���<嚏<���<��<a_�<�!�<�΄<�k�<q�<�{<0v<
Yq<�l<K�g<fec<��^<��Z<�V<��R<�N<A�J<��F<�B<��><`�:<�b6<��1<�>-<�y(<d�#<A�<��<�<�k<h�<�^<f
<ױ�;��;��;3�;{�;��;i\�;���;W��;�M�;%��;���;P�;�(�;U�;��;��t;��d;��U;b�G;c[:;R.;��";%q;��;��;���:�O�:*��:��:���:E�:��:��:V�`:%!?:EQ:�:�s�9��9Y�h9s�9M �80!8�1綑�F��ȴ�����&4���k�Pؖ�kF����蹴f���%�ѳ?�}pY�mBr��ք����i����d��pD���3���K��i��� ���+�ƺ�̺��Һ�oں<e�/��s���9,�j�	�������� ��P$�**��O/�^4�R8�<�q|?�ÎB�xE��iH�ʘK��8O�tS�_bX�^��Md��k�a"r��Gy��'��懃����������Y���Ɏ������쒻p���dD��˗��  �  �=O�=s�=�9=�=(�=�=}�=�+=�� =9: =ݏ�<^��<e��<	O�<���<�9�<z��<�n�<f�<I��<�s�<��<��<��<"|�<#��<��<�:�<�h�<֘�<	��<��<�Y�<ׯ�<0�<�}�<���<Ex�<?�<��<�1�<���<�T�<T��<�=�<F��<B��<���<��<��<h#�<�1�<�I�<o�<X��<]��<o@�<s��<��<U��<���<�_�<��<���<Y
�<���<���<|{�<��<�w�<a��<��<ia�<���<���<��<+�<XU�<[�<w��<6��<��<�,�<pM�<`�<<_�<�F�<��<�ɲ<�h�<���<�}�<y�<g��<j�<+¡<�x�<�C�<d$�<
�<x�<Z3�<�N�<xj�<K�<q��<{�<�Y�<f#�<�ل<���<M!�<�z{<�v<��q<8Vm<ʿh<�<d<��_<=w[<�7W<�S< O<��J<�G<��B<�><ű:<�Q6<*�1<-<�3(<�A#<�E<�M<-g<?�<��
<z|<�-<��;.(�;Ҁ�;�;~��;�b�;��;�L�;Df�;/8�;�ɮ;6+�;.u�;:;�,�;K̃;ew;$�g;)�X;t�J;u=;��0;�6%;�];�N;u�;m�:V��:���:��:(޶:���:8�:�&:bLZ:��6:�:H�9�>�9,�9�l19N�8<8m���&������yݸ[d��Z>�_7r��o��e'��׽�)
���!�"�9�V�Q�(�h�ZH~�Z��p蒺ZЛ����ޭ����������'���(ź�v˺3tҺ�ں���Q�������(��D�ː����a� �tb'�8d-���2�+y7�*�;�9�>���A��D��G��I�iL�?�O���S�Z�X���]���c��Yj���p�,�w�]4~��>��:���
��r���*��My�����(����n��m2���  �  �=A�=��=D2=��=�u=�='�=Z=p� =b =r6�<VX�<F��<'��<~Q�<m��<�u�<�#�<��<���<UK�<���<N��<&�<�n�<���<��<�J�<t��<6��<7�<[�<���<��<]p�<���<G�<��<�:�<]��<TH�<��<tS�<d��<-�<xz�<D��<��<���< ��<=��<'��<���<�	�<t:�<M��<���<G�<}��<�@�<���<�1�<���<���<���<���<e��<�{�<��<o��<L��<�V�<&��<k��<o-�<�a�<e��<���<���<B��<?�<�'�<OB�<tV�<�^�<V�<7�<���<Ӭ�<�C�<�ȭ<�B�<���<�5�<#��<[�<�<5ڜ<���<���<kϖ<��<��<N=�<	[�<ji�<%d�<HI�< �<�ل<W��<k:�<��{< )w<��r<Z�m<zi<��d<A�`<�$\<��W<�S<�YO<9K<�!G<_C<��><h�:<�*6<J�1<��,</�'<4�"<s�<��<Ա<��<}!
<�<�W<*��;���;�G�;R�;���;z��;:b�;��;�;���; ��;;0�;˪�;�0�;Tی;H��;�y;ozj;4�[;5�M;8@;�b3;�J';L�;?i;��;}�:���:Z�:�_�:W[�: ֢:�ݏ:�Jy:S:��-:	�
:��99]�P9��84[8�y��s�+�Mޙ���Ӹ/W��3&�fHM�5~�<͜��ۿ�7b繵	��+��l5�72K��.`��Bt�C���
���땺Q����Ԧ�%������$��;ĺ�˺��ҺSGۺ���A�7���.e�����x���#��c*�/�0�66�x�:���>��A��fD��F��H��J��M���P��tT�7�X�0^���c�#�i�<1p�Ibv�kl|�N��wꃻ����2��D���%���w��=����Ô��Ŗ��  �  �
=�=iy=�'=C�=�e=;�=y=6� =�r =D��<���<���<�3�<��<���<S��<�&�<S��<���<:d�<� �<���<�h�<���<	[�<���<��<�Q�<���<���<D>�<��<���<u[�<"��<�#�<؉�<��<�c�<���<�T�<|��<!J�<]��<��<^�<���<���<��<Ũ�<`��<���<a��<k��<H��<�!�<��<���<cu�<.��<��<�<�i�<ò�<E��<���<���<fs�<S�<0��< �<H��<���<V4�<{�<��<���<���<��<;$�<�2�<�@�<�M�<ZV�<�U�<�E�<� �<�<���<�<���<�	�<�v�<�<�i�<;��<5��<.|�<@f�<%k�<���<˯�<u��<�<�3�<�G�<�G�<O2�<�	�<|ф<���<�I�<�|<Ӂw<~s<U�n<Bj<�e<]'a<?�\<�GX<%�S<��O<�^K<A-G<��B<#�><|o:<]�5<2S1<Ё,<Y�'<�n"<3F< <�<�< c	<��<� <� �;y�;�&�;3�;%
�;���;���;�R�;S��;曶;eh�;��;A��;x�;(\�;Pu�;��{;̦l;�,^;�P;�B;�i5;��(;o1;/;�;j�:C��:n��:i��:҂�:{��:>V�:�Xs:�L:��%:�]:)��9��9�r!9�"�8R�7H�)�nҡ��ܸR3��5��c:��m^�A��j���yPĹ��鹍	����O2��EF��{Y��l��+~�����	�����pࢺ����Fѳ�(Ȼ��ú�P˺�Ӻ>{ܺ�溣#�������$\��L��?���%�-�+�3�<9�h�=��oA��]D���F���H�M`J�^TL�ưN��Q�
OU�_�Y���^��#d��i���o��tu�H
{��7���ւ�i��4�����������������@F��U����  �  ;
=&�=q=�=F�=�V=4�=�e=�� =Y =P��<��<���<��<M:�<���<6<�<`��<��<�n�<.9�<"��<z��<�K�<p��<$F�<6��<���<�R�<p��<	�<%a�<D��<�-�<6��<���<[�<��<��<O��<���<�Z�<E��<�=�<���<���<�B�<�o�<��<���<?z�<h�<vY�<�V�<h�<$��<���<R8�<���<�8�<���<rX�<���<�F�<��<þ�<:��<֥�< h�<��<���<�'�<���<�	�<�f�<���<���<��<	6�<dD�<�J�<�M�<[P�<?R�<�Q�<;I�<R3�<�	�<Wȴ<�l�<���<p�<�٪<�?�<S��<�%�<߶�<�d�<2�<G�<>)�<�J�<-{�<n��<��<,�<~(�<Y,�<�<g��<5Ƅ<���<TQ�<*.|<$�w<�Ws<��n<��j<�f<V�a<�]<"�X<i,T<��O<�sK<�-G<��B<ԣ><�E:<�5<�1<�>,<a:'<�"<r�<�<�<e�<��< G<D <R�;�s�;[<�;�=�;�T�;v\�;48�;���; ,�;�?�;�"�;��;���;ş�;��;���;��|;jBn;��_;k�Q;�/D;��6;�%*;;
;�;F;��:O�:���:XU�:n��:᫞:?�:7n: 0F:s:��9b�94$d9rM�8w�8�׷�w���޸�'	����>�2��lL��Ln��0�������"ɹ�<�U�	�:�m\0�#�B�ǪT�3f�kKw�th��i��S���`���p@���G��h����eúx�˺�iԺ�ݺ�(躨��t� �n����i�����,�'��:/���5��g;�6@�%�C�iF���H�Q4J���K���M���O��R�\"V�@`Z�i7_�yd���i�sto�_�t��z����������d������@?��tގ�Is����C\���  �  �=�=�j=�=ʵ=>L=R�=sX=� =)H =Z�<�z�<d��<���<w
�<�|�<��<G��<��<N�<�<J��<X��<�6�<���<�6�<;��<}��<�Q�<��<P�<�u�<���<uN�<۸�<�<g}�<���<�3�<��<���<K\�<���<�3�<���<V��<./�<�Y�<~l�<#k�<"[�<E�<(2�<�+�<:�<�b�<$��<$
�<τ�<N�<_��<Q9�<Q��<7.�<�~�<���<}��<O��<�^�<��<ѥ�<"1�<���<>"�<�<��<��<A�<�X�<b�<b�<�]�<[X�<QS�<|L�<!?�<g%�<��<��<�V�<�߯<T�<R��<��<#��<���<;��<�4�<��<��<���<�#�<�X�<���<eː<���<q�<��<�	�<��<���<s��<^T�<LC|<��w<��s<a/o<)�j<�^f<��a<*]]<��X<!TT<C�O<�}K<*G<��B<��><P&:<-�5<>�0<�,<�'<��!<��<x^<6<�5<�l<_�<�G�;`M�;��;��;���;d��;O��;���;Y}�;�ܽ;3��;��;s˥;L��;���;��;$H�;E�};�>o;�a;��R;=:E;��7;��*;*�;��;�;u��:uj�:߸�:�6�:�|�:�D�:���:��j:�@B:�:���9&!�9��L9k{�8
ot7��H���ø�n�#���-���@��X��ly��.�����{�̹���9l
�?�AY/�<�@���Q�\]b�!s��$��1+�� ���n<���觺�e��`����lú+̺�!պ�޺eK��3���I����=������!!��')��0�h?7���<� �A�PE�y�G��I��EK�\�L��eN�7�P��DS��V���Z���_��d�nj��Zo�5�t��y�vU~�����Y����z���������zv��'���œ�8L���  �  /=�=�x=_&=��=\=u�=Q=�� =b =���<���<��<���<G$�<���<�K�<D�<i
�<��<s �<���<,��<uq�<z�<dw�<=��<;0�<<��<���<_�<m��<�`�<��<r^�<���<$�<%r�<ѻ�<��<�_�<��<�3�<��<��<�z�<R��<g��<���<��<^��<xb�<�,�<_	�<=�<�&�<�t�<���<��<�G�<0�<z��<���<'.�<۞�<���<���<��<]��<�E�<���<�t�<�<���<���<�R�<��<���<H��<қ�<7z�<gV�<�7�<�!�<��<��<��<Y��<�h�<���<^�<$��<�۪<	�<{>�<<9��<<��<�X�<Q�<t�<r��<_�<t�<>ϐ<'�<pC�<@P�<�?�<��<��<1��<=w�<n�|<pVx<.t<��o<גk<$g<%�b<�]<z$Y<ulT<Y�O<MGK<��F<&�B<P><��9<�l5<ɩ0<��+<�T&<8� <�3<j�<�<��
<��<�<���;!��;o��;c�;s��;m�;���;�2�;���;�W�;}Q�;|
�;\��;l�;�`�;���;�)�;��w;��i;t~[;�CM;��>;)�0;�#;��;l�	;�#�:���:���:;��:�+�:nϟ:.k�:՛o:�LD:o�:\��9�
�9���8���+7 ���P��b��#L�����������ܒ����s���x*����T�ùt�F�R��ħ'��@8�EEG��U��nb�Bep�����ڈ�	ɒ� j���=���ò������źeEκR�ֺ��ߺB������*��.
�g0�|��Y\&��/�8�5x?��fE�d�I�g�L�XwN�60O�.YO��dO�K�O�g�P�d�R�!+V�hQZ��5_���d�q�i��o�b�s�*Mx�r|�gH��Br���Մ��~���c���f��hi��9L��d����  �  =��=y}=�+=��=/b=��=�W=D� =�  =t�</��<���<���<C;�<I��<a�<.1�<��<�<A�<O��<���<�}�<
�<ԁ�<Y��<:7�<��<��<9[�<���<QU�<���<8N�<��<��<Le�<X��<�<Y^�<h��<�9�<S��<�#�<���<-��<���<���<5��<���<�s�<�?�<�<��<�=�<���<�<���<�Z�<�"�<��<ơ�<;�< ��<`��<���<���<p��<0K�<��<is�<M��<�y�<M��<C�<���<��<ܡ�<@��<5q�<bQ�<�6�<�$�<��<<
�<>�<A·<<t�<��<k�<a��<o�<��<R�< ��<��<-��<�o�<g�<���<}˕<�#�<���<qݐ<c$�<�O�<@\�<K�<{"�<��<O��<�x�<��|<`Ix<�	t<K�o<sk<Bg<�pb<��]<kY<�]T<��O<�HK<K�F<��B<4b><�:<��5<��0<(�+<5p&<�� <AU<�<�5<��
<1�<�E<��;�9�;t�;�c�;c��;Ѫ�;}2�;3h�;�1�;���;�}�;,1�;�͢;�}�;�c�;1��;��;��w;25i;= [;��L;�>;�f0;��";��;Ӳ	;�O�:'%�:�v�:
��:��:��:34�:�Dq:�F:(�:!6�9eވ9��8 ��Zt�[AE��{����!ݒ��G��:莹�o���N��I������ ���u���4�2��1O'��`8�4�G�T0V� d�Jr�����߉�����f'��$¨����������ź��ͺ$ֺ�ߺ�3�C1��6����	�^��X8��%��/�@u7�V�>�
�D�KI�wL���M�t�N� �N� �N��WO��}P���R�A�U���Y�c�^��Id���i�Uo���s�Q�x�G�|�l~��)���k��u���ޚ��<���C����W�������  �  �=��=G�=�:=��= s=��=>k=�� =v8 =�<�<��<>�<F2�<�~�<n��<���<�j�<kP�<&D�<�8�<& �<Q��<	��<�-�<���<���<�I�<��<���<"O�<���<v2�<+��<��<q��<���<]>�<c��<���<�X�<��<wH�<u��<�>�<(��<���<=�<l�<��<���<���<�v�<?Z�<[�<���<���<�D�<D��<��<	T�<�<L��<S_�<���<S�<o�<���<��<zY�<4��<�m�<c��<B\�<X��<h�<=M�<�l�<vs�<-i�<�U�<�A�<d3�<z+�<�'�<k �<��<�<���<�#�<A��<Jݭ<��<)M�<6��<vܢ<YO�<n�<���<B��<Dė<��<JT�<b��<#�<aI�<�r�<_}�<�i�<;=�<� �<���<�|�<Є|<%!x<J�s<�so<�k<��f<�b<Co]<0�X<�0T<��O<KK<'G<x�B<�><B:<��5<Q1<1,<ϼ&<qF!<x�<�"<V�<sj<�q<�<;�;:�;��;":�;8��;pX�;b��;g��;��;~�;���;���;a�;���; i�;�h�;@��;�wv;�g;��Y;�@K;�=;9/;��!;�=;w�	;l��:�"�:���:[_�:
״:ا�:Zf�:g�u:dK:�l:���9Y��9�9�[�7�5���#�L�Z���{��|ͅ��ă��c����B]�������5����ٹ����0���u&�p�8��I� �Y�ʾh�'�w�J���팺�w��If���U���߳�d���`�ĺ��̺r�ԺBݺ�<纁󺓎 �R���r����3$�&>-���5�q�<���B�G��J���K���L�QM�l�M�� N�b\O��Q�y�T�*Y�m^�ͣc��Zi���n�+7t��!y�w�}��!��n��
߅�8}��B������ڐ�l}�����  �  O =��=��=�N=��=��=/=	�=�� =\ =6��<s�<Bt�<���<}��<�_�< �<���<���<Z��<�u�<xV�<!�<���<*Y�<#��<��<�`�<���<U��<�7�<:��<g��<c�<���<�6�<��<��<Id�<m��<�K�<���<uZ�<���<�c�<���<��<fF�<xP�<x>�<�<&��<o��<,��<���<���<�6�<?��<�;�<���<���<aW�<��<Ȓ�<"��<A7�<�A�<��<���<�j�<��<}_�<=��<�)�<O�<���<���<|�<�'�<*�<'�<R%�<�(�<-1�<�:�<�=�<0�<��<���<�R�<�°<��<�Z�<S��<U�<p;�<ƴ�<'S�<g�<u
�<2 �<zT�<���<��<�>�<�}�<���<��<���<�a�<��<p͂<}�<�b|<j�w<`s<t�n<�wj<��e<\qa<K�\<�ZX<��S<ĄO<�CK<�G<��B<��><m�:<�6<�`1<De,<T+'<��!<�C<��<�b<K1<�C<��<���;J��;�i�;��;���;�W�;���;q��;P��;`Ǽ;p��;�(�;��;Yߚ;4\�;��;��;��t;�e;vW;��H;	�:;�E-;*c ;�R; 4	;��:�[�:���:H��:w��:���:ay�:W�|:�jR:��':�O�9˫9��F9���8mo��Of޸�x(���L��M_���e��jf���g���o�&5���[������3йs.��3���%�O:���M�P�_�<�p��������x瑺�����!������s��+5��hĺ�_˺#�Һ��ںϋ�=:���x��������F�!��*�^�2�9��M?���C��G�� I�g]J�VK�%�K��^L�t�M�P��fS�8�W�H�\�8�b���h���n��t�N<z��e�A.������F"������T���펻9p��;ʓ�����  �  5$=	�=&�=�b=[=��=�+=9�=�=�� =	��<��<���<�<Gl�<*��<(y�<0�<���<���<���<��<�V�<+��<^��<���<�9�<�t�<p��<���<p�<#W�<���<�<�c�<���<�4�<c��<��<֢�<j2�<F��<�g�<���<W��<���<�I�<~y�<q��<��<of�<�H�<�1�<+�<�<�<!l�<���<�'�<���<�N�<���<:��<�C�<��<.�<wd�<5j�<z@�<���<Rv�<b��<E�<a��<���<c$�<\�<���<`��<���<���<(��<��<u�<�.�<�H�<�W�<mR�<�0�<��<���<���<�Y�<S��<���<�J�<y��<�4�<�מ<���<m��<���<��<���<C;�<��<��<c׍<dڋ<�<�<�5�<�ׂ<�t�<'|<%qw<��r<�2n<�i<�e<�`<�#\<��W<pS<+?O<,)K<�%G<v%C<�?<�:<p6<��1<f�,<C�'<^T"<��<H�<�E<�+<NM<�<���;W��;]-�;?�;�7�;t�;C��;&��; V�;߆�;@I�;>��;��;���;�)�;��;1�;#Jr;��b;��S;�zE;D�7;N�*;�H;i�;�|;���:�P�:M��:��:DA�:e��:q��:��:Y�Z:�S1:��:v��99)[9rX8d�3���Ѹ?��3�*�_28��b?��<F���R���j�f�������ǹE�T���&��'=�;7S��g��r{�����Z珺&����$���N������.�UU��@Jĺ�>ʺ/�к�tغI��47�!������l� $����K&'���.��5�?(;�ձ?��"C�f�E��:G��YH�nII��cJ��L�N���Q��}V��[��b���h�Y6o���u���{��ۀ�ڞ��(E���ֈ��Z��Bˍ����vL��;L��?$���  �  e!=�=ն=Wq=�=^�=C=��=�;=�� =	- =U^�<y�<���<Y�<r�<���<���<�d�<�/�<f��<���<���<�$�<���<u�<#M�<z{�<���<'��<��<_�<eB�<��<���<6F�<��<v7�<P��<fa�<y	�<���<�g�<�<���<��<�m�<G��<`��<6��<��<���<h��<H��<���<���<�N�<l��<�1�<���<�W�<^��<l��<���<�V�<Ć�<-��<�V�<���<|t�<7��<��<:U�<@��<���<���< �<�!�<�B�<f�<���<Һ�<���<d�<�I�<pe�<&i�<�M�<��<v��<6.�<=��<��<�W�<��<�6�<Yġ<l�<1�<��<��<y'�<PQ�<%��<J��<��<��<>��<Z݉<ל�<,B�<6Ղ<@^�<
�{<Y�v<Wr<4Mm<��h<Bd<��_<8[<��V<�R<��N<��J<�G<m4C<-:?<!;<��6<}2<\--<�(<��"<�<�c<�?<�B<nw	<]�<Ό <���;��;��;M��;B��;���;�|�;��;��;�ȵ;�;��;��;[��;|��;��;�:o;�,_;��O;5vA;n�3;>';ɖ;��;7K;*��:�w�:ȝ�:��:�O�:��:%v�:��:J�b:;:�:���94ݠ9')O9�8��7	*�2#���g�& ����&��29�L1U�~�~��������4a칍y�A(��A�\[��r��v�����*���ɠ�e����Ư������5f��{ź��ɺp�Ϻ��ֺ#�ߺ��꺚����`�[�B��Դ��w#���*���0���6��;���>��A�/�C��E�G�i�H���J��;M���P��U��9[�u�a��h���o��#w�~��T��f��
A��"犻�Z��ٙ�����=r��"��y����  �  r=��=ķ=�u=�#=��=R=s�=�Y=!� =o` =���<-�<]E�<��<-�<���<��<���<�{�<�7�<j��<r��< 8�<��<�<	M�<�o�<���<,��<̔�<3��<���<�<]P�<���<F+�<b��<�[�<v�<r��<w��<<U�<d�<��<�!�<~�<ٺ�<"��<���<���<w��< �<�,�<�Y�<��<"��<�F�<���<�.�<E��<a5�<c��<��<m�<g��<ҏ�<�X�<���<�_�<��<���<&�<C�<f2�<�J�<Mg�<��<��<���<W&�<�k�<δ�<��<]7�<�_�<�k�<"V�<v�<cĳ<Q�<�̮<t@�<2��<02�<���<�W�<��<�ȝ<V��<^��<4��<m��<�Ɠ<S�<U
�<��<l�<��<?��<J<�<5��<(6�<5M{<�4v<�/q<�Gl<=�g<��b<Ts^<',Z<�V<�R<�NN<ӔJ</�F<�C<9?<� ;<��6<�52<�g-<Gn(<Q\#<C<u3<�9<�_<�
<�<ɾ<T�;Z�;�R�;��;V��;�X�;��;cb�;�e�;���;��;��;҄�;�;ӱ�;�+};�k;�[;NxK;��<;<�/;�g#;�d;�};��;���:�{�:|z�:�,�:��:��:j
�:ZR�:�h:$�C:��:��9h�9�֋9�%:9ri�83	8F�k���e�������긌S�k�'��H��v�[0���p��c;���VZ,���H���d�C���7���f��sQ���ꩺz6���B���'���$��B�ú=�ƺپʺ�Ϻ�WֺZ�޺��麔J��?/��	��B����7���e&��^,��1��\6�\_:���=�j�@�E�B��
E��&G���I� �L��gP��BU��#[�]�a�lbi��5q��y��h��'��om��A|��7��ܙ��9���Pe���ٔ�����6���  �  O =��=w�=�n=�=,�=�V=��=p=�� =� =�% =���<���</�<w��<�	�<��<��<ٹ�<�_�<��< ��<�4�<��<� �<�6�<�O�<S�<SJ�<D@�<�>�<bN�<�u�<s��<�<���<'3�<��<1��<���<�^�<�/�<C��<ȑ�<9�<�w�<z��<��<x�<l)�<�I�<�q�<��<���<�)�<�y�<���<�.�<���<��<1j�<���<�+�<�m�<$��< ��<D�<,��<8�<t�<���<���<���<���<��<y��<��<s�<�b�<��<0�<�m�<�ƿ<D�<�C�<�V�<EG�<e�<�ų<�`�<�<y�<A�<+��<T:�<L�<���<NZ�<@(�<��<��<�<���<7�<Z�<i�<v
�<݉<��<]!�<���<��<��z<nu<>p<P2k<WUf<Ѯa<CB]<�Y<U<NQ<h�M<J<)�F<��B<?<' ;<�6<02<Ox-<�(<�#<��<B�<Y!<hm<�<ZM<)�<2,�;t��;���;���;	J�;?��;)-�;�h�;VP�;!͵;7ج;�~�;�ݙ;e�;�n�;G�y;��g;ֺV;�F;�C8;�+;2P;|�;��;(d;���:�O�:l �:$-�:�x�:�ī:�?�:"J�:Y�l:A%J:2w):)O:���9[I�9uȁ9��39��8�;8߳ж��N��Y������J���gG���x�"����ù[�j
���2�~�Q�op��}�����P檺{r���3��NK��e�ºl�źͭǺ��ɺ��̺�(ѺZ׺��ߺ���%���ٔ��{�Sh����{�tm"��'��-���1�E.6�W:���=�f�@�ߔC��PF��6I�b�L�s�P���U��[���b��j��s�ֈ{�����A����Ҍ�����󑻜Փ��N��1p���V��S%���  �  ��=��=ę=�]='=��=)R=-�=w}=�=m� =�V =)��<V�<��<��<zz�<���<b�<���<�u�<E	�<��<��<��<U��<��<��<��<d �<J��<���<p��<B��<"%�<5��<�<���<?s�<-N�<Y5�<��<���<n��<8l�<���<�\�<���<���<G�<�K�<��<|��<g�<�[�<J��<?��<�J�<ʘ�<��<F:�<؍�<P��<8'�<m[�<q�<�^�<!�<Ӧ�<� �<T0�<�?�<�:�<-�<� �<V�<�.�<�R�<���<���<�?�</��<��<��<3۽<��<�.�<�$�<���<���<�^�<���<䠬<�F�<��<��<�`�<4�<�۞<8��<j�<s@�<�$�<��<��<��<�	�<T��<-��<�i�<#��<Gb�<�r<c	z<؟t<Lo<�!j<=0e<f�`<V\<��W<�T<wP<3�L<�I<�F<&|B<�><۷:<Yy6<�2< d-<d�(<��#<g0<�<5�<�Z<|�<�[<Q�<���;�W�;
��;��;��;��;o�;��;��;Q�;�E�;�̢;I��;f�;n�;��v;� d;�zR;�TB;�3;�&;eE;�Q;�;�� ;���:)�:�h�:���: ��:O8�:"A�:n�:�n:;�N:A�0:&�:��9��9��9[�u9E�*9x��8j�8����F��*[��� ��vO�₹4���	͹�=�������:�ʚ[���|�5�������w��V/��C���}�ºSEǺ�ɺ�b˺�h̺��ͺZ�Ϻ��Ӻ��ٺ��zn�;���Ӎ����/��������
$���(��-�[|2�Z�6�6;��?�ުB�qF�tI�p.M���Q���V��\��:d�bl�g'u�\1~�,��� ч�ⱋ�������;������8��P�������>���  �  	�=}�=�="G=I�=}�=EG=��=��=�&=�� =�} =b. =���<# �<|�<���<2�<]��<��<0}�<���<g��<���<
c�<[��<���<���<���<���<Ӎ�<�l�<P^�<cm�<ɡ�<���<���<L7�<"�<���<2��<X��<���<ȍ�<><�<<��<[7�<���<D��<Y�<�^�<��<�<�`�<���<��<5h�<���<���<�)�<e�<O��<=��<��<m=�<DJ�<`1�<��<�o�<<��<���<���<��<U��<���<d��<��<���<T�<�e�<���<�O�<���<!@�<���<߻<���<���<]ӵ<(��<�O�<��<&��<�u�<9�<� �<fǣ<
��<�F�< �<���<�|�<�J�<�&�<��<��<��<�ʋ<5��<I:�<]��<1&�<��~<�cy<��s<@on<�,i<�*d<	u_<v[<�W<�:S<��O<�HL<�H<��E<�
B<ZQ><�Z:<'6<��1<7-<��(<1$<�t<��<!�<�<�<�;	<�<s= <0��;���;�4�;��;7��;���;��;U�;姴;D��;���; �;��;���;�s;_�`;ߪN;Q>;w�/;_�";�;;,�;��:��:���:�>�:��:��:<��:*��:<�:(�n:�Q:\#6:��:��:���9��9a �90�\9�i9��8��}5�+s�2��(�$�]����kͮ���ع�����"��%C��pe�����������p���u��@�ĺ��ʺ9}κ�Nк��к�%ѺۺѺtӺ��ֺe~ܺ�&�ȡ��j�����ײ��B�(���p��)�s� ��%�Qt*��z/��4�y_9�+�=��6B�z2F��J��*N��R�� X�l^���e�vIn��[w��d��^��܈������������E���㗻��������x��^���  �  h�=D�=�i=(1='�=R�=�:=X�=�=�0=�� =<� =�P = =�p�<���<<�<�e�<���<��<E|�<���<�e�<���<�9�<���<��<8��<B��<!v�<E�<B�<��<N
�<�9�<ʖ�<&"�< ��<���<���<���<���<<��<�\�<@�<X��<��<�m�<���<I�<g�<$��<J0�<U��<Y�<lg�<��<R��<�+�<>W�<���<٫�<���<� �<t�<�"�< �<k��<�<�<��<_��<��</��<�f�<�D�<3�<�9�<_�< ��<��<~�<��<���<��<�g�<.��<͹<>˷<F��<Jy�<<�<D��<�Ŭ<Ԕ�<oj�<�@�<��<�ڡ<���<G�<���<ܥ�<�a�<�,�<��<p�<�ˍ<s��<�g�<��<4��<5��<�l~<��x<?@s<0�m<�ih<�[c<$�^<�AZ<^;V<,�R<�
O<�K<prH<�E<��A<��=< :<_�5<=z1<w-<ł(<�$<��<�D<=�<�<"P<t�	<L\<�� <9f�;=X�;4��;��;}��;\�;�"�;軼;� �;�֪;�7�;�4�;��;���;�q;�];)�K;�#;;�s,;�;V�;xi;ut;,��:X�:U]�:�D�: L�:PZ�:��:֖�:�ͅ:�m:�5R:�|9:�d#:S3:���9T��9��9�9�.9MI�8k�r7 7^��:���2��l�:����i���M� ���e)�!�J���m�Dň������������ ú'n˺�Ѻ�GԺ��պ��պ�1պ�Oպ��ֺ�ٺ�Mߺa��e�ﺵ3���z�������_�����g!�s��	#���'��F-�g�2�u8��D=��B���F���J��6O��S��}Y�t�_��yg���o�Fy��{���O���늻F�����a���Tᗻ�j��p\��Aݚ�M��xV���  �  =�=^=�X="!=v�=��=�0=��=�=�5=�� =ҩ =f = =���<���<�@�<���<
��<D�<Fx�<f��<�P�<G��<��<Cb�<���<��<)x�<�J�<��<:��<(��<5��<��<~S�<r��<W��<�x�<�p�<Ft�<�t�<�d�<�9�<	��<�<|��<'V�<���<��<&i�<,��<J�<���<�3�<>��<��<Q%�<�P�<�q�<���<���<���<���<z�<��<���<&��<��<De�<S��<�y�<X�<�,�<��<���<r��<��<ia�<���<8E�<���<[�<5ھ<<A�<���<���<)��<׏�<b�<\,�<���<�ʬ<��<N��<�g�<A�<�<hƟ<ir�<w�<Ͻ�<�m�<-�<
��<֏<���<>��<�H�<��</l�<�ʁ<�~<L|x<�r<RIm<��g<F�b<!^<S�Y<Q�U<�R<q�N<�WK<�H<�D<cYA<"�=<[�9<C�5<vF1<��,<Vk(<�$<��<�q<�:<q�<?�<kG
<P�<�<���;���;���; ��;�d�;��;���;�J�;��;�T�;p��;Ӟ�;GL�;e�;�to;��[;��I;�9;d*;�;��;b�	;�;�(�:��: �:Q#�:DG�:Pr�:�:�%�:ń:b�l:n�R:�K;:��&:��:��:���9bt�9!\�9%RA9�u�8;M�7U<W�����:��_x�����)��u�����.���O��\s��狺֎���ƭ�ֻ��3ǺR�ϺPպnغ1�غL�غ��׺��׺��غ�ܺ2X���4�񺐐�������,�������-�����B}!�{&�D�+� �1��a7�9�<�?B���F�4mK�$�O��T�-|Z�a�Q�h��.q��z�5�� ���ҋ�����ƶ��F똻"g���E��/����ۛ�a����  �  `�=�x=�R=L= �=��=%-=[�=��=s7=b� =B� =m =' =8��<]�<�M�<���<V��<p�<}v�<>��<�H�<���<��<V�<�}�<��<,j�<�;�<��<I��<���< ��<)��<�<�<���<2��<Ne�<�^�<6d�<Of�<W�<�,�<��<�s�<@��<MM�<��<��<xi�<���<�R�<���<�B�<���<���<E4�<�\�<�z�<o��<V��<���<B��<���<���<T��<�<��<�W�<Zs�<�h�<�E�<��<���<b��<���<G�<lJ�<<��<_1�<ý�<�J�<k˾<�3�< {�<C��<���<���<TY�<g&�<X��<̬<���<���<�t�<gP�<��<�֟<Ӏ�<�"�<�Ř<�q�<�,�<I��<�Ϗ<ɪ�<�}�<S=�<�߆<�_�<.��<M�}<r[x<H�r<3!m<��g<m�b<��]<"�Y<P�U<��Q<�yN<�5K<�G<�D<?A<:�=<w�9<s�5<f31<s�,<Zb(<�$<�<t�<2Q<<�<�i
<��<�7<{�;c��;��;���;�R�;Z��;Ȝ�;�!�;yY�;&�;�{�;i�;��;��;��n;�K[;�I;�d8;9�);A�;.;�	;�[;V.�:���:pH�:e_�:ϋ�:B��:oH�:���:�_�:.Kl:ƖR:��;:��':4M:�q:x�9���9@!�9ԅG9va�8wG�7(�U��t����=�K�|����S�ù������/��XQ�gYu���nƞ�����=����Ⱥ�ѺF�ֺRٺ!"ں*�ٺ��غz�غu�ٺ��ܺ�iX�G5�������������2~���J� ���%��{+��I1��$7�_�<�aB�#G�i�K��FP�H:U��Z� ba�@�h�5�q�){��v��~i���"���l��������F��𽚻Q���g���1���;���  �  =�=^=�X="!=v�=��=�0=��=�=�5=�� =ҩ =f = =���<���<�@�<���<
��<D�<Fx�<f��<�P�<G��<��<Cb�<���<��<)x�<�J�<��<:��<(��<5��<��<~S�<r��<W��<�x�<�p�<Ft�<�t�<�d�<�9�<	��<�<|��<'V�<���<��<&i�<,��<J�<���<�3�<>��<��<Q%�<�P�<�q�<���<���<���<���<z�<��<���<&��<��<De�<S��<�y�<X�<�,�<��<���<s��<��<ja�<���<9E�<���<[�<6ھ<>A�<�<���<+��<ُ�<b�<^,�<���<�ʬ<��<O��<�g�<A�<�<hƟ<ir�<v�<ν�<�m�<-�<	��<~֏<���<<��<�H�<��<-l�<�ʁ<�~<J|x<��r<QIm<��g<F�b<!^<S�Y<R�U<�R<s�N<�WK<�H<�D<fYA<%�=<^�9<F�5<yF1<��,<Yk(<�$<��<�q<�:<r�<@�<kG
<P�<�<���;���;���;��;�d�;��;���;�J�;��;�T�;j��;͞�;AL�;_�;wto;��[;��I;�9;d*;�;��;^�	; �;�(�:��:�:O#�:CG�:Or�:�:�%�:ń:b�l:n�R:�K;:��&:��:��:���9bt�9!\�9%RA9�u�8<M�7U<W�����:��_x�����)��u�����.���O��\s��狺֎���ƭ�ֻ��3ǺR�ϺPպnغ1�غL�غ��׺��׺��غ�ܺ2X���4�񺐐�������,�������-�����B}!�{&�D�+� �1��a7�9�<�?B���F�4mK�$�O��T�-|Z�a�Q�h��.q��z�5�� ���ҋ�����ƶ��F똻"g���E��/����ۛ�a����  �  h�=D�=�i=(1='�=R�=�:=X�=�=�0=�� =<� =�P = =�p�<���<<�<�e�<���<��<E|�<���<�e�<���<�9�<���<��<8��<B��<!v�<E�<B�<��<N
�<�9�<ʖ�<&"�< ��<���<���<���<���<<��<�\�<@�<X��<��<�m�<���<I�<g�<$��<J0�<U��<Y�<lg�<��<R��<�+�<>W�<���<٫�<���<� �<t�<�"�< �<k��<�<�<��<_��<��</��<�f�<�D�<3�<�9�< _�<!��<��<~�<��<��<��<�g�<1��<͹<A˷<I��<My�<<�<F��<�Ŭ<֔�<pj�<�@�<��<�ڡ<���<G�<���<ڥ�<�a�<�,�<��<n�<�ˍ<p��<�g�<��<1��<2��<�l~<��x<;@s<-�m<�ih<�[c<$�^<�AZ<`;V<.�R<�
O<�K<urH<�E<��A<��=< :<e�5<Cz1<}-<˂(<�$<�<�D<?�<�<#P<t�	<K\<�� <4f�;6X�;,��;��;r��;\�;t"�;ܻ�;� �;u֪;�7�;�4�;��;���;�q;ٻ];�K;�#;;{s,;�;N�;qi;ot;$��:Q�:P]�:�D�:L�:NZ�:��:Ֆ�:�ͅ:�m:�5R:�|9:�d#:R3:���9T��9��9�9�.9MI�8l�r7�6^��:���2��l�:����i���M� ���e)�!�J���m�Dň������������ ú'n˺�Ѻ�GԺ��պ��պ�1պ�Oպ��ֺ�ٺ�Mߺa��e�ﺵ3���z�������_�����g!�s��	#���'��F-�g�2�u8��D=��B���F���J��6O��S��}Y�t�_��yg���o�Fy��{���O���늻F�����a���Tᗻ�j��p\��Aݚ�M��xV���  �  	�=}�=�="G=I�=}�=EG=��=��=�&=�� =�} =b. =���<# �<|�<���<2�<]��<��<0}�<���<g��<���<
c�<[��<���<���<���<���<Ӎ�<�l�<P^�<cm�<ɡ�<���<���<L7�<"�<���<2��<X��<���<ȍ�<><�<<��<[7�<���<D��<Y�<�^�<��<�<�`�<���<��<5h�<���<���<�)�<e�<P��<=��<��<m=�<DJ�<`1�<��<�o�<<��<���<���<��<V��<���<f��<��<���<W�<�e�<���<�O�<���<&@�<���<#߻<���<���<aӵ<,��<�O�<��<)��< v�<�9�<� �<gǣ<
��<�F�< �<���<�|�<J�<�&�<��<��<��<�ʋ<1��<E:�<Y��<-&�<��~<�cy<��s<<on<�,i<�*d<	u_<w[<�W<�:S<��O<�HL<�H<��E<B<bQ><�Z:<'6<��1<7-<�(<8$<�t<��<%�<�<�<�;	<�<q= <)��;���;�4�;��;(��;���;ҥ�;�T�;ӧ�;2��;���;��;v�;濃;��s;G�`;ɪN;�P>;g�/;Q�";�;;%�;��:֢�:���:�>�:��:��::��:(��:;�:'�n:�Q:[#6:��:��:���9��9a �90�\9�i9��8	�}5�+s�1��(�$�]����kͮ���ع�����"��%C��pe�����������p���u��@�ĺ��ʺ9}κ�Nк��к�%ѺۺѺtӺ��ֺe~ܺ�&�ȡ��j�����ײ��B�(���p��)�s� ��%�Qt*��z/��4�y_9�+�=��6B�z2F��J��*N��R�� X�l^���e�vIn��[w��d��^��܈������������E���㗻��������x��^���  �  ��=��=ę=�]='=��=)R=-�=w}=�=m� =�V =)��<V�<��<��<zz�<���<b�<���<�u�<E	�<��<��<��<U��<��<��<��<d �<J��<���<p��<B��<"%�<5��<�<���<?s�<-N�<Y5�<��<���<n��<8l�<���<�\�<���<���<G�<�K�<��<|��<g�<�[�<J��<?��<�J�<ʘ�<��<F:�<؍�<P��<8'�<m[�<q�<�^�<!�<Ӧ�<� �<U0�<�?�<�:�<-�<� �<X�<�.�<S�<���<���<�?�<4��<��< ��<8۽<��<�.�<�$�<���<���<�^�<���<蠬<�F�<��<��<�`�<4�<�۞<7��<j�<p@�<�$�<��<��<��<�	�<O��<'��<�i�<��<Bb�<�r<[	z<ҟt<Lo<�!j<;0e<e�`<W\<��W<�T<
wP<:�L<�I<�F</|B<�><�:<cy6<�2<*d-<m�(<��#<n0<�<:�<�Z<~�<�[<O�<���;�W�;���;��;ִ�;��;[�;l�;��;�P�;vE�;�̢;4��;S�;\�;��v;� d;}zR;�TB;��3;�&;WE;�Q;�;�� ;���:)�:�h�:���:���:L8�: A�:m�:�n::�N:@�0:%�:��9��9��9[�u9E�*9x��8k�8����F��*[��� ��vO�₹4���	͹�=�������:�ʚ[���|�5�������w��V/��C���}�ºSEǺ�ɺ�b˺�h̺��ͺZ�Ϻ��Ӻ��ٺ��zn�;���Ӎ����/��������
$���(��-�[|2�Z�6�6;��?�ުB�qF�tI�p.M���Q���V��\��:d�bl�g'u�\1~�,��� ч�ⱋ�������;������8��P�������>���  �  O =��=w�=�n=�=,�=�V=��=p=�� =� =�% =���<���</�<w��<�	�<��<��<ٹ�<�_�<��< ��<�4�<��<� �<�6�<�O�<S�<SJ�<D@�<�>�<bN�<�u�<s��<�<���<'3�<��<1��<���<�^�<�/�<C��<ȑ�<9�<�w�<z��<��<x�<l)�<�I�<�q�<��<���<�)�<�y�<���<�.�<���<��<1j�<���<�+�<�m�<%��<!��<D�<-��<8�<t�<���<���<ä�<���<��<|��<��<w�<�b�<��<5�<�m�<�ƿ<J�<�C�<�V�<KG�<k�<�ų<�`�<�<y�<D�<.��<V:�<M�<���<NZ�<>(�<��<��<�<���<2�<U�<c�<q
�<݉<��<X!�<���<��<�z<nu<>p<L2k<UUf<Ѯa<DB]<�Y<U<$NQ<o�M<J<3�F<��B<%?<2 ;<#�6<'02<Zx-<�(<�#<��<H�<^!<km<�<ZM<'�<,,�;j��;��;z��;�I�;+��;-�;�h�;>P�;͵;ج;�~�;�ݙ;P�;�n�;"�y;��g;��V;��F;�C8;�+;#P;o�;��; d;���:�O�:d �:-�:�x�:�ī:�?�:!J�:W�l:?%J:1w):(O:���9[I�9uȁ9��39��8�;8سж��N��Y������J���gG���x�"����ù[�j
���2�~�Q�op��}�����P檺{r���3��NK��e�ºl�źͭǺ��ɺ��̺�(ѺZ׺��ߺ���%���ٔ��{�Sh����{�tm"��'��-���1�E.6�W:���=�f�@�ߔC��PF��6I�b�L�s�P���U��[���b��j��s�ֈ{�����A����Ҍ�����󑻜Փ��N��1p���V��S%���  �  r=��=ķ=�u=�#=��=R=s�=�Y=!� =o` =���<-�<]E�<��<-�<���<��<���<�{�<�7�<j��<r��< 8�<��<�<	M�<�o�<���<,��<̔�<3��<���<�<]P�<���<F+�<b��<�[�<v�<r��<w��<<U�<d�<��<�!�<~�<ٺ�<"��<���<���<w��< �<�,�<�Y�<��<"��<�F�<���<�.�<E��<a5�<c��<��<m�<g��<ҏ�<�X�<���<�_�<��<���<'�<D�<g2�<�J�<Pg�<��<��<���<[&�<�k�<Ӵ�<���<c7�<�_�<�k�<(V�<|�<iĳ<Q�<�̮<x@�<6��<22�<���<�W�<��<�ȝ<U��<[��<1��<i��<�Ɠ<N�<P
�<��<f�<��<9��<D<�<0��<#6�<-M{<�4v<{/q<�Gl<;�g<��b<Vs^<*,Z<�V<�R<�NN<ܔJ<9�F<�C<"9?<� ;<�6<�52<�g-<Rn(<Z\#<C<|3<�9<�_<�
<�<Ⱦ<M�;O�;�R�;���;C��;�X�;��;Kb�;ke�;���;��;��;���;��;���;�+};«k;r[;3xK;s�<;)�/;zg#;xd;�};��;���:�{�:tz�:�,�:��:��:h
�:XR�:�h:#�C:��:��9h�9�֋9�%:9ri�83	8D�k���e�������긋S�k�'��H��v�[0���p��c;���VZ,���H���d�C���7���f��sQ���ꩺz6���B���'���$��B�ú=�ƺپʺ�Ϻ�WֺZ�޺��麔J��?/��	��B����7���e&��^,��1��\6�\_:���=�j�@�E�B��
E��&G���I� �L��gP��BU��#[�]�a�lbi��5q��y��h��'��om��A|��7��ܙ��9���Pe���ٔ�����6���  �  e!=�=ն=Wq=�=^�=C=��=�;=�� =	- =U^�<y�<���<Y�<r�<���<���<�d�<�/�<f��<���<���<�$�<���<u�<#M�<z{�<���<'��<��<_�<eB�<��<���<6F�<��<v7�<P��<fa�<y	�<���<�g�<�<���<��<�m�<G��<`��<6��<��<���<h��<H��<���<���<�N�<l��<�1�<���<�W�<^��<l��<���<�V�<Ć�<-��<�V�<���<}t�<8��<��<;U�<B��<���<���< �<�!�<�B�<f�<���<׺�<���<j�<�I�<ve�<,i�<�M�<��<{��<;.�<A��<#��<�W�<��<�6�<Zġ<l�<1�<��<��<v'�<LQ�< ��<E��<��<��<8��<T݉<ќ�<&B�<0Ղ<;^�<�{<R�v<Rr<0Mm<��h<Bd<��_<8[<��V<�R<��N<��J<�G<w4C<8:?<,;<��6<�2<g--<�(<��"<��<�c<�?<�B<pw	<]�<̌ <���;��;��;=��;/��;���;}|�;��;��;lȵ;��;��;��;F��;h��;��;�:o;�,_;��O;vA;\�3;�=';��;��;/K;��:�w�:���:��:�O�:��:#v�:��:G�b:~;:~�:���93ݠ9&)O9�8��7*�2#���g�% ����&��29�K1U�}�~��������4a칍y�A(��A�\[��r��v�����*���ɠ�e����Ư������5f��{ź��ɺp�Ϻ��ֺ#�ߺ��꺚����`�[�B��Դ��w#���*���0���6��;���>��A�/�C��E�G�i�H���J��;M���P��U��9[�u�a��h���o��#w�~��T��f��
A��"犻�Z��ٙ�����=r��"��y����  �  5$=	�=&�=�b=[=��=�+=9�=�=�� =	��<��<���<�<Gl�<*��<(y�<0�<���<���<���<��<�V�<+��<^��<���<�9�<�t�<p��<���<p�<#W�<���<�<�c�<���<�4�<c��<��<֢�<j2�<F��<�g�<���<W��<���<�I�<~y�<q��<��<of�<�H�<�1�<+�<�<�<!l�<���<�'�<���<�N�<���<:��<�C�<��<.�<xd�<5j�<{@�<���<Sv�<c��<E�<b��<���<e$�<\�<���<c��<���<���<,��<��<z�<�.�<�H�<�W�<rR�<�0�<��<���<���<�Y�<W��<���<�J�<z��<�4�<�מ<���<l��<���< ��<���<?;�<��<��<^׍<_ڋ<轉<섇<�5�<�ׂ<�t�<'|<qw<��r<�2n<�i<�e<�`<�#\<��W<pS<1?O<3)K<�%G<%C<?<�:<p6<��1<o�,<L�'<fT"<��<N�<�E<�+<OM<�<���;P��;T-�;3�;�7�;d�;1��;��;V�;ʆ�;*I�;(��;��;���;�)�;	��;1�;Jr;��b;��S;�zE;4�7;@�*;�H;`�;�|;���:�P�:F��:��:@A�:b��:o��:��:W�Z:�S1:��:t��99([9pX8e�3���Ѹ?��3�*�_28��b?��<F���R���j�f�������ǹE�T���&��'=�;7S��g��r{�����Z珺&����$���N������.�UU��@Jĺ�>ʺ/�к�tغI��47�!������l� $����K&'���.��5�?(;�ձ?��"C�f�E��:G��YH�nII��cJ��L�N���Q��}V��[��b���h�Y6o���u���{��ۀ�ڞ��(E���ֈ��Z��Bˍ����vL��;L��?$���  �  O =��=��=�N=��=��=/=	�=�� =\ =6��<s�<Bt�<���<}��<�_�< �<���<���<Z��<�u�<xV�<!�<���<*Y�<#��<��<�`�<���<U��<�7�<:��<g��<c�<���<�6�<��<��<Id�<m��<�K�<���<uZ�<���<�c�<���<��<fF�<xP�<x>�<�<&��<o��<,��<���<���<�6�<?��<�;�<���<���<aW�<��<Ȓ�<"��<A7�<�A�<��<���<�j�<��<}_�<>��<�)�<P�<���<���<~�<�'�<*�<!'�<V%�<�(�<11�<�:�<�=�<0�<��<���<�R�<�°<��<�Z�<U��<W�<q;�<Ǵ�<'S�<f�<t
�<0 �<xT�<���<��<�>�<�}�<���<��<���<�a�<��<l͂<}�<�b|<e�w<`s<q�n<�wj<��e<]qa<M�\<�ZX<��S<ʄO<�CK<�G<��B<��><u�:<�6<�`1<Le,<[+'<��!<�C<��<�b<M1<�C<��<���;E��;�i�;��;���;�W�;���;`��;?��;NǼ;_��;q(�;�;Hߚ;%\�;��;��;�t;һe;cW;{�H;��:;�E-;!c ;�R;�3	;��:�[�:���:D��:s��:���:_y�:U�|:�jR:��':�O�9~˫9��F9���8po��Of޸�x(���L��M_���e��jf���g���o�&5���[������3йs.��3���%�O:���M�P�_�<�p��������x瑺�����!������s��+5��hĺ�_˺#�Һ��ںϋ�=:���x��������F�!��*�^�2�9��M?���C��G�� I�g]J�VK�%�K��^L�t�M�P��fS�8�W�H�\�8�b���h���n��t�N<z��e�A.������F"������T���펻9p��;ʓ�����  �  �=��=G�=�:=��= s=��=>k=�� =v8 =�<�<��<>�<F2�<�~�<n��<���<�j�<kP�<&D�<�8�<& �<Q��<	��<�-�<���<���<�I�<��<���<"O�<���<v2�<+��<��<q��<���<]>�<c��<���<�X�<��<wH�<u��<�>�<(��<���<=�<l�<��<���<���<�v�<?Z�<[�<���<���<�D�<D��<��<	T�<�<L��<S_�<���<S�<o�<���<��<{Y�<5��<�m�<d��<C\�<Y��<i�<>M�<�l�<xs�</i�<�U�<�A�<g3�<}+�<�'�<n �<��<�<��<�#�<D��<Mݭ<��<*M�<8��<wܢ<ZO�<n�<���<B��<Cė<��<HT�<_��<!�<^I�<�r�<\}�<�i�<8=�<� �<���<�|�<̄|<!!x<H�s<�so<�k<��f<�b<Do]<2�X<�0T<��O<KK<,G<~�B<��>< B:<��5<V1<6,<Լ&<vF!<|�<�"<Y�<tj<�q<�<9�;:�;��;:�;0��;gX�;W��;\��;ݾ�;q�;���;;T�;���;�h�;�h�;6��;�wv;��g;��Y;�@K;�=;�8/;��!;�=;s�	;e��:�"�:���:X_�:״:֧�:Yf�:e�u:cK:�l:���9X��9�9�[�7�5���#�L�Z���{��|ͅ��ă��c����B]�������5����ٹ����0���u&�p�8��I� �Y�ʾh�'�w�J���팺�w��If���U���߳�d���`�ĺ��̺r�ԺBݺ�<纁󺓎 �R���r����3$�&>-���5�q�<���B�G��J���K���L�QM�l�M�� N�b\O��Q�y�T�*Y�m^�ͣc��Zi���n�+7t��!y�w�}��!��n��
߅�8}��B������ڐ�l}�����  �  =��=y}=�+=��=/b=��=�W=D� =�  =t�</��<���<���<C;�<I��<a�<.1�<��<�<A�<O��<���<�}�<
�<ԁ�<Y��<:7�<��<��<9[�<���<QU�<���<8N�<��<��<Le�<X��<�<Y^�<h��<�9�<S��<�#�<���<-��<���<���<5��<���<�s�<�?�<�<��<�=�<���<�<���<�Z�<�"�<��<ơ�<;�< ��<`��<���<���<p��<0K�<��<is�<M��<�y�<M��<C�<���<���<ݡ�<A��<6q�<dQ�<�6�<�$�<��<=
�<?�<B·<=t�<��<k�<b��<p�<��<R�<��<��<.��<�o�<g�<���<|˕<�#�<���<pݐ<a$�<�O�<?\�<�J�<y"�<��<M��<�x�<��|<^Ix<~	t<J�o<sk<Bg<�pb<��]<mY<�]T<��O<�HK<M�F<��B<7b><�:<��5<��0<+�+<8p&<�� <CU<�<�5<��
<2�<�E<��;�9�;q�;�c�;^��;̪�;w2�;-h�;�1�;���;�}�;%1�;|͢;�}�;�c�;,��;��;��w;*5i;6 [;��L;�>;�f0;��";��;в	;�O�:$%�:�v�:��:��:��:34�:�Dq:�F:'�: 6�9eވ9��8��Zt�[AE��{����!ݒ��G��:莹�o���N��I������ ���u���4�2��1O'��`8�4�G�T0V� d�Jr�����߉�����f'��$¨����������ź��ͺ$ֺ�ߺ�3�C1��6����	�^��X8��%��/�@u7�V�>�
�D�KI�wL���M�t�N� �N� �N��WO��}P���R�A�U���Y�c�^��Id���i�Uo���s�Q�x�G�|�l~��)���k��u���ޚ��<���C����W�������  �  ��=ӯ=m=�%=��=�f=��=_H=� =ͼ�<�E�<K��<���<��<���<�}�<I�<�J�<�r�<���<���<���<���<ߞ�<[*�<I��<@��<�&�<�|�<��<_v�<��<x��<�x�<-�<B��<���<a�<=%�<N�<:��<<��<�[�<���<>m�<:��<QB�<yn�<wg�<�0�<���<�h�<���<��<܎�<��<���<��<Ka�<�Y�<�i�<Dx�<�n�<�7�<���<:�<��<*��<ӭ�<(O�<t��<ҋ�<�1�<��<Sm�<���<�(�<9�<��<���<.u�<e�< ��<���<-��<㏼<j��<�]�<��<풳<%ް<���<��<�ۧ<|Τ<�<�"�<���<df�<�m�<#��<�#�<���<2G�<E̐<)0�<h�<bq�<�Q�<��<�̈́<k��<�W�<L{|<urx<�t<y�p<�kl<nh<RQc<�[^<�@Y<^(T<W7O<ƂJ<mF<��A<��=<�u9<�5<�Q0<m.+<ԣ%<��<�<u�<K<��<"|<ie�;i��;+q�;���;���;�d�;���;���;If�;8�;Z�;d�;":�;�|�;���;��;�^�;�~;5q;ɬc;�U;�zG;wc8;��(;�;�&;���:���:2m�:O��:�B�:�$�:�:E}t:YVJ:�:Ԥ�9��c9E8�e	�����@�Ź����������G���6�ۖҹ:��s���삹���ǹ'��U�m��$^)��:��*I��T�UZ\�8�c��&m��y�(Ʌ�nߐ�I����ܪ�"���d�ºXY̺KmԺ��ۺ>�<-����������S��-!���,�9�7�؆A���I�3P��iT���V�*�V�x�U�T��UR�n=Q��[Q��S��<V�d�Z�nZ`��<f��k�H�p��*u���x�H\{�@.~��ɀ�3���hƅ�T������|[��j������  �  ��=ط={v=�/=��=�p=1�=S=S� =���<#`�<� �<���<b��<}�<��<�g�<g�<���<C��<,��<�
�<���<w��<?�<^��<���<6�<���<F��<uu�<{�<��<�f�<��<�k�<��<���<�<MJ�<ӎ�<���<�h�<���<���<���<�V�<#��<m|�<;F�<k��<`��<��<T��<Y��<���<��<���<�~�<)u�<J��<"��<&��<�L�<��<z&�<�3�<?�<���<L\�<���<[��<�-�<���<>]�<b��<]�<�"�<'�<��<l�<��<���<���<��<%��<���<�q�<�%�<��<��<|�<��<���<�<��<�B�<nÜ<��<���<NΖ<�>�<6˓<,^�<)�<xE�<}�<t��<lf�<)�<Eބ<Ζ�<J_�<�}|<�gx<�lt<�kp<�Bl<r�g<m'c<&8^<�'Y<cT<T7O<ӎJ<�&F<��A<��=<��9<u65< z0<�W+<n�%<��<6�<]�<>�<1<�<���;�i�;���;>T�;b�;���;�*�;N<�;���;���;��;�D�;���;���;�*�;?�;�]�;Tb~;y�p; c;�CU;`�F;��7;�v(;�Y;g;�"�:�7�:H�:㴿:��:s�:�i�:�w:��L:�:�k�9aBp9ćF8�7��@Ņ�8���ɰ�j���ڑ���l���}�̹ߠ��Q[��kT��d�¹(�ܹQ���ص���'�c�9���H�GuT��]���e���o�G�|�������_v��$_��$���i�ºR�˺��Ӻ}�ںU�ẓ���8��\O�u��C�u[ ��+�1�6�]�@���H��,O�eS�b�U���U��U�2VS���Q�X�P�]�P��\R�$�U�2Z���_�/�e���k���p�!u���x�5�{�`�~�����R�����fZ��L医fs��S���ħ���  �  �=��=�=�K=��=�=\=�p=�� =� =���<�S�<?%�<<-�<�s�<��<���<d��<���<`�<22�<�E�<�1�<b��<px�<O��<q!�<�_�<���<���<�p�<���<��<�/�<s��<�+�<��<���<i��<:=�<^��<D�<D��<�"�<���<P5�<���<,��<��<���<�,�<���<�h�<u#�<V	�<
%�<|�<�<|��<���<6��<���<.��<b��<%�<_�<Vk�<<@�<k��<(��<�	�<���<p �<���<e,�<���<���<���<q��<?��<�O�<>�<���<���<�̾<�ϼ<�ɺ<���<�]�<q߳< ,�<�J�<�I�<�<�<�9�<�T�<鞟<j"�<a�<\�<�"�<ߋ�<[�<���<�<�<:��</��<e��<�]�<��<��<�r�<%�|<�Dx<%t<p<��k<�Vg<`�b<=�]<��X<]�S<3O<R�J<)dF<�DB<�2><�
:<��5<��0<]�+<�D&<�l <�b<fP<�`<"�<�|<n�;���;�V�;s��;���;��;�,�;�2�;���;�~�;���;>)�;@V�;�j�;}��;�@�;R�;|�};�ro; xa;W\S;��D;B�5;�';�h;��
;A��:v��:o��:��:0�:��:u�:�v~:�dT:m_&:o��9��9���8E���/�]�6	��(�˹��แ
�2�޹�Ϲ|���i�������ʥ��P��%�ι�]������"���6�k�G���U��@a�	�k���v�sU�����D��� $��'�����&���S�ɺT�к%�׺^�޺�N�ښ��} ��@	�$W��G��t)�`04���=���E�A4L��sP���R��ZS�i�R��,Q���O�ǲN�X�N�y�P���S�rX��"^��Rd�{j��'p�Uu�I?y���|�d%��X��BT��U�� +��%{��~������b���  �  "=��=˳=0r='=^�=%3=Y�=�� =�> =�< ��<���<A��<��<݋�<H�<h4�<E�<Bh�<c��<��<7��<A<�<��<�&�<�f�<��<}��<H�<nb�<y��<�O�<���<�R�<���<:�<�q�<���<G"�<��<� �<��<�b�<���<-��<��<��<>�<���<	��<s0�<���<���<�<��<E�<)��<�X�<S:�<_2�<�,�<��<���<V`�<��<7��<E��<d+�<��<�$�<���<��<�s�<��<-�<�a�<t�<g�<E�<��<o��<���<���<���<^�<��<��<z��<�+�<�z�<���<J��<��<沥<Iۢ<�.�<E��<0x�<�s�<D��< �<�x�<c��<gt�<�ҏ<��<��<N�<^��<bJ�<��<���<hx|<x<<�s<Zo<��j<Zf<��a<\]<�TX<�S<�O<T�J<W�F<�B<F�><�:<�A6<��1<�h,<��&<� !<�,<%5<�a<L�	</�<7��;�5�;��;	��;%\�;5t�;8��;��;���;/��;Y�;Eh�;qy�;�Y�;6K�;!��;�$�;�o|;sYm;�^;35P;<�A;03;?�$;ݾ;��	;?��:^��:m��:���:f��:{�:��:�<�:r�^:1:F�:�;�9^9��]����� ����������Ĺ���������㤹3���)|��w�� ���c��c�߹������2��<G���X��g��Su�jn���ٕ��V�����⯺�+��?$����Ǻa�ͺ�?Ӻ�ٺmg����	��д�y��uB��&�-\0���9��sA���G���K�adN��UO�	O���M�B�L��L��bL��N��SQ�V��[�1gb�'i�-vo��:u��Jz���~�Yx��;�������ݤ��҆���|���T���ᓻ����  �  �5=R	=��=ژ=tF=��=�[=��="=�x =`��<�n�<*]�<�w�<���<XB�<���<���<���<g��<���<'��<V��<��<��<'s�<���<���<���<
�<D�<���<��<�V�<���<�0�<���<�<�q�<���<ϊ�<5�<���<3��<�I�</��<!.�<[�<�Y�<�1�<|��<��<�l�<�H�<H�<2r�<���<�N�<	��<���<1��<���<�n�<�&�<}��<��<��<���<�i�<���<q8�<���<���<m �<�g�<���<���<G��<���<��<e��<m��<���<��<0�<P�<nY�<>�<��<�w�<�˱<���<��<R&�<_F�<��<Q�<r�<�1�<o#�<�C�<_��<��<�a�<�Α<&�<Z�<cb�<�=�<��<숅<A�<\��<�S|<�w<O�r<Rkn<��i<�Xe<�`<$\<�W<5(S<;�N<c�J<��F<�(C<�G?<�6;<�6<="2<*-<ߖ'<��!<<
F<�<q3<�<�c<��;?�;4�;�z�;HE�;0�;���;�P�;�;n4�;㬳;*��;�H�;T��;��;;#zz; Xj;��Z;�K;27=;m�.;�,!;|G;"�;�M�:��:���:��:�d�:n�:w �:HJ�:Si:��<:�:���9d�[9|�8��v�5�$��.p��5��޲��Ƙ��P���A�������pu��d|��錹������̹����wo���/�$'H�|^�8�q�����������������r]���!���J��kQ���!����ź�9ʺ��κպ%�ݺ��躎��t�M������"�b�+��_4��;�G�A��F�I�H�-eJ���J��RJ��I�BUI���I�P�K���N��S���Y��~`���g�>o�M�u���{�)ƀ��Q���ǅ��C��ӊ�k������A>��2<��Fꕻ�  �  �?=�=��=!�=.c=��=�z=�=�N=�� =0 =X�<��<�E�<A��<��<۫�<�m�<�M�<�B�<?�<�2�<j�<���<�N�<$��<���<u��<7��<���<��<2�<gk�<Ÿ�<��<	~�<@��<r�<��<B��<cj�<Z7�<��<���<��<9
�<�g�<2��<^��<�~�<R�<�#�<��<��<��<�B�<՚�<��<���<ya�<�(�<���<ǻ�<{f�<���<�.�<S8�<��<
��<���<�8�<�f�<w��<���<���<��<��<*(�<�9�<�L�<�i�<A��<���</�<�L�<x{�<���<Xr�<�(�<���<��<�I�<>x�<���<�<78�<���<=D�<l�<'�<k�<��<f�<��<a�<�g�<3��<b��<y�<�(�<���<�)�<9��< |<{�v<�	r<h>m<c�h<�c<�a_<z�Z<k�V<bzR<4�N<��J<}G<[sC<}�?<��;<\I7<�2<`�-<Z&(<��"<H�<�`<)�<"�<�<4<�`�;�;�;b��;���;�
�;ޜ�;"�;�\�;p�;o0�;F��;��;f�;�-�;�s�;���;1�w;@uf;�V;��F;n�7;�);m�;��;�x;Q�:[_�:���:��:��:Ľ�:�ڟ:��:�`q:�eF:=�:���9i�9G�9A38|p�|5���<�v^�7�l�>�l�yFc�O~X�bT�P�^��}��8��K��4���!H/��K��df�k�~�;��e��y��T����d��h��FM��.뾺9eºz.ź�Ⱥ9�˺�Ѻ��ٺ6%��C���������*��(�&���.��w5�n";�V�?���B��E�$CF��F���F�\G�V�G��I��M���Q�!�W�,_��g�w.o�bw�Mw~�����妅�`s�����L���"̏��ԑ�싓��	���  �  �:=�!=k�=|�=�m=a=��=- =Vp=A� ={Y =��<U��<��<�m�<���<�e�<4
�<r��<=��<8|�<�Z�<*�<��<d�<y��<���<b��<t��<���<���<I��<C��<{�<�M�<Բ�<�1�<���<j�<~M�</0�<��<��<���<̒�<,�<�|�<���<ڻ�<���<��<ʎ�<v��<T��<��<2�<p�<���<n]�<���<Y��<YD�<	��<,��<���<�@�<�I�<�<���<���<��<�*�<�+�<�)�<�*�<r2�<A�<�W�<Uy�<ʨ�<h��<;:�<F��<��<�I�<{��<ڙ�<<�9�<�Ŵ<�-�<i��<�ʬ<��<�y�<��<�x�<�<�ԝ<���<��<���<�̕<��<�L�<ω�<`��<O��<W��<�<�<d��<�#�<it�<�{< &v<��p<��k<�g<�Qb<��]<ƅY<�rU<A�Q<�M<�vJ<�G<�|C<��?<;�;<�n7<��2<�-<@}(<h#<ʹ<�h<�;<�;<Jj	<��<#X <�:�;�9�;���;ӊ�;ݫ�;#��;���;8��;
��;�
�;�ի;��;_�;�ڍ;CЃ;>t;a�a;��P;�l@;�1;�#;6�;��;��;��:q��:���:2��:�O�:�7�:ZV�:(Î:[�u:��L:��$:ؼ�9��9�s9��94B;8�5��B���t���#���4���;���=�}�B���Q�H<r���lp��գ�׵��22�zR���q�Ko��z{��0柺����j����6�������ĺXRź�Fƺ��Ǻ%�ʺ^к��غ�㺋��a� �3?	�m���:�'�!�V�(��/��j4��9���<���?� B���C���D�
�E���F��I�oiL�w-Q�idW���^��Kg��4p�('y�$܀��τ��]��)����>�����������X=�����~����  �  Q%="=�=�=pc=��=�=�=A�=n=�� =�& =p��<[��<+9�<6��<��<~��<w.�<J��<Y��<a�<��<���<:O�<>��<C��<���<��<*��<Z�<5�<�)�<�>�<z�<��<je�<*�<7��<��<���<���<]��<N��<�|�<
�<�h�<���<���<h��<���<���<=
�<�C�<���<%��<�9�<{��<���<�o�<Q��<w�<��<u��<D��<"*�<�0�<M��<�~�<���<���<���<B��<���<�q�<2a�<�c�<�{�<1��<���<7V�<���<�E�<���<p"�<Df�<�~�<ng�<�!�<#��<O-�<_��<z�<�y�<���<��<�8�<C�<���<�^�<�0�<��<��<�4�<�\�<���<棎<���<�}�<�(�<"��<	��<�6�<�z<E,u<ïo<#gj<_e<��`<�)\<�X<'(T<��P<1M<��I<(�F<8;C<�?<-�;<�@7<�2<��-<��(<j#<�K<�H<g<ץ<��
<i<��<��;��;[`�;u��;	C�;��;���;{X�;�a�;=ʹ;�;찡;�^�;nь;L�;!"p;v�\;��J;��9;�*;Ƕ;�0;�\;E ;��:���:h��:Z��:}!�:��:�=�:���:��u:"�O:��*:�&	:Q�9�d�9�=f9��9���8���6ϚP��ȸ^�v9!���2���B�m�X���{��3��oտ����c1��9��\����V�����������%��bg��Pź��Ⱥ�ʺ��ʺ��ɺnaɺ�ɺ�s̺�Ѻ�ٺ����P�� ��_�l��+�h��{�#��	)�N.���2�,/7�>!;��z>�9.A��QC��'E�2G���I�M���Q�RX���_��h�)r�� |�ς�:I��eK���������ޓ�ꇕ�k����?��烗�*����  �  z=�=��=-�=9G=
�=
r=%�=��=�=z� =d =� =���< ��<MI�<���<��<�{�<��<���<�H�<���<���<^�<�p�<���<>��<?q�</�<���<5��<�}�<4}�<Q��<�	�<��<�^�<�J�<)W�<�t�<���<���<���<9C�<���<e1�<o�<���<Q��<���<@�<=l�<���<.�<z��<���<�;�<���<_��<-�<���< ��<�b�<J��<)��<>��<غ�<k>�<���<P��<�i�<0�<;��<M��<��<��<���<���<N@�<���<�J�<���<k�<�۾<�%�<�?�<9)�<�<�<F�<k��<�"�<���<�k�<&$�<�ߣ<ʘ�<�K�<"��<M��<�u�<SQ�<�E�<�O�<�c�<�s�<
o�<�F�<���<j�<��<��<b�y<2t<)hn<~�h<C�c<$�^<щZ<2�V<��R<�uO<�JL<�4I<�F<��B<�?<�;<L�6<I,2<�W-<sj(<*#<N�<��<2a< �<d_<��<|E<=f�;&c�;Ĭ�;Y�;7i�;���;�A�;���;U��;[��;R��;�Ơ;�F�;�o�;>��;��k;$wW;أD;�3;ۉ$;`�;��;�;�N�:���:���:+��:��:���:d��:O�:��:��q:	sN:��-:��:���9>"�9ӳ�9ʀl9�b"9��8�7-�B���ϸ��2"6��R��pp���������7ιy �*���C�N.i�����KK���ު����Bĺ�o̺�ѺG�Ӻ��Ӻ�8ҺW�Ϻ)κ��ͺs#кtJպhwݺ�N����s�a�o�����A�%���#��y(��T-�K2�+7�O�;���?���B��E�iEH��'K�R�N�-�S���Y���a�	�j���t��f��섻�Չ�8��{�~攻0���}���9���i��	B������  �  .�=��=��=�p=� =[�=�T=i�=
�=,)=�� =q� =�P =o =�}�<���<��<8`�<��<��<��<��<���<�J�<���<"�<�M�<�H�<��<��<En�<p�<���<���<���<N�<9��<���<ٶ�<���<C�<:4�<�H�<E6�<s��<&��<|��<+�<c�<���<*��<wC�<���<&2�<G��<��<}z�<ܾ�<���<� �<VT�<���<���<x.�<yu�<I��< ��<�h�<8��<5)�<�)�<o��<ڭ�<+X�<��<���<���<e��<�*�<F��<�(�<}��<�s�<�<ф�<Ѽ<d�<�ָ<혶<w@�<4ݱ< ~�<�,�<��<׽�<蔦<�f�<�)�<�ٟ<�y�<��<ʷ�<�o�<yB�<I/�<�-�<�/�<$�<+��<<��<�b�<�<�y<Ms<�5m<&�g<sRb<Oy]<�Y<�$U<��Q<�cN<�`K<4kH<�[E<�B<�t><G|:<#-6<��1<��,<f(<6m#<p�<�q<C"<��<~<�	<x`<�L�;���;_��;߱�;?@�;�1�;R_�;��;3r�;�ղ;���;_��;k��;N�;�~};��g;��R;�E?;��-;��;;)�;d�:��:wH�:��:��:'�:Y�:eި:1K�:��:�]k:PK:%.:�j:>� :$�9�:�9.<�9��j9k}9j �8�}%��;��Z;�;�B�!�k�j؈�����������Ag
���)�ЊN��xv�鱏�Pf��w1���=ĺB�Ϻ�غڝܺQ�ݺ��ܺ��ٺ�^ֺ[�Ӻ�Ӻ�պT5ں�V���캤��A��J������b������������#���(��c.��4�Ȩ9�V�>�C���F��	J��ZM��4Q��V�g]\��-d�ptm���w�t��7���{8���␻f̔��֗����.��Ĥ��T����
�������  �  Ӭ=�=%�=�I=2�=ۛ=L7=��=	{=�-=�� =X� =�| =�> =���<m6�<In�<C��<���<��<]w�<'��<�x�<��<{�<\��<���<���<���<~n�<��<���<b]�<bA�<�]�< ��<mW�<1�<=�<�k�<8��<N��<B��<3��<���<�3�<���<`��<X-�<a{�<���<fV�<y��<�{�<��<���<g��<��<�>�<=S�<�i�<���<+��<5��<P1�<iU�<�R�<`�<h��<&��<#��<ܗ�<"?�<���<݂�<&F�<�1�<�L�<��<�<��<>`�<��<\��<�0�<�~�<���<���<6L�<���<���<Za�<�*�<8�<��<7�<�Ȥ<ړ�<)A�<�ԝ<�Z�<��<�}�<"5�< 
�<;��<��<�ً<#��<zV�<�̈́<T�<�S~<IMx<�6r<\;l<��f<�-a<ON\<��W<UT<��P<~M<}�J<��G<#�D<�nA<F�=<i�9<n�5<4
1<�h,<��'<0I#<+�<��<��<i�<O<�	<�.<�T <W��;�"�;���;���;���;�v�;�x�;�K�;���;{a�;/`�;Բ�;���;cz;�d;�N;k�:;�i);@;�;�b;Ѩ�:���:�o�:���:���:�V�:%�:��:���:�ł:��d:��F:l-:S�:�: �9e��9d��9���9a]J9��8�t7�䐸�>�7�R�9Ȃ�{p��<��ɜι;����D�x4�hMY��)��$^���ꪺ�����-ͺ�4ٺ�F�yq庋��些Aມ(ܺ�ٺغ�ں�!ߺ3���b��]�C�	�����~������v��� �ï%���+���1��Z8�?L>���C���G�d�K���O���S���X�]�^�v�f��p�
�z�*���)����+�������C'���:���W��M���KE�����8��  �  �=�='f=�,=s�=q�=�!= �=�r=�.=0� =�� =)� =c] = =�r�<]��<��<��<Y�<Uc�<���<?K�<���<�B�<���<���<Z��<���<�.�<&��<�X�<?	�<��<���<[�<���<���<���<�"�<
f�<��<]��< ��<�k�<���<�c�<���<��<�`�<a��<7^�<��<���<#E�<��<�"�<W�<�k�<{o�<s�<^��<@��<���<T �<Y�<-�<���<r]�<d��<���<�S�<���<��<�)�<h��<���<Z��<(;�<M��<�^�<4�<���<�t�<��<tB�<�]�<�J�<e�<�ͳ<(��<�I�<�$�<*�<9�<*�<��<�Ӣ<��<@�<a��<b��<���<�'�<R�<N͏<Ϻ�<���<�t�<m�<��<�ց<$�}<��w<�q<~�k<��e<�q`<T�[<V1W<�WS<7�O<-�L<c	J<:3G<8D<p�@<�\=</f9<�5<�0<�,<b�'<�(#<�<��<9�<|�<��<C`
<_�<z� <�i�;cn�;���;p��;��;#��;��;�t�;̰;I��;�;7˒;���;Fx;�a;�L;�68;��&;BV;E�
;� ;���:���:
f�:M�:��:)ȼ:���:"��:�U�:T�:��_:j�C:��+:a�:'
: !�9>��9�b�9E��9F6g9�#9��7 ׆��y��_�Ta���g��̭��b�ܹ����v`;�8�`��B��ܚ��ޯ���º�Һ�"ߺ�/纀��j�a�躈��.ຏ�ܺF�ۺ��ݺ����S���~���{�wy
�$�������(~�������#���)�Y�0�ϥ7�h.>���C���H�>%M��Q��QU�WZ��`��zh���q��|����-≻Xr���h��]�����������ໞ�$螻�q������'휻�  �  k�=s|=�[=h"=P�=y=�=P�=�o=�.=[� =�� =� =�g =� =׆�<��<
��<���<��<�[�<N��<�:�<u��<{.�<��<��<l��<,s�<�<˩�<;>�<,��<���<	��<S:�<��<��<>��<�	�<�N�<��<<��<5��<W�<���<�O�<���<��<�V�<��<,`�<��<ص�<�W�<]��<<8�<%j�<�z�<{x�<�u�<�<���<x��<Z��<9
�<�<���<H�<���<cz�<�;�<���<}m�<�<���<1��<���<��<���<�B�<���<.��<�]�<�ݽ<�,�<|H�<�5�<O�<��<�w�<RA�<�!�<��<f�<�$�<��<��<���<`�<���<��<���<�"�<��<E��<���<�<[`�<'	�<r�<���<߫}<`�w<]nq<�^k<T�e<1`<L[<��V<}S<8�O<��L<��I<rG<�D<��@<�2=<<9<p�4<}0<��+<rt'<#<��<��<�<R<�<ό
<�<� <���;���;���;��;���;9��;�h�;&�;y|�;�2�;W.�;�w�;�;�;|�w;Z�`;d3K;�A7;��%;�T;��	;f��:(�:���:���:��:\��:���:.N�:cL�:�:�Z}:�!^:ckB:Y+:�2:+*:��9���9ƿ�9��9��p9W�9p+	8���-I���c��㏹ Ω�ܙù��ṙ��� ��>���c�v���1m��������ĺ��Ժm/Ắ:���@�m��0�����,޺�
ݺ1�޺��L�o��|� ����c�
�!��
����(��������#�S)�YJ0�6m7�*>�o#D�k;I���M�ܯQ���U���Z��Ha��!i�/�r�/F}��j���I��{㏻�┻C���&��3��7��\Z��ڞ�S
���F���  �  �=�='f=�,=s�=q�=�!= �=�r=�.=0� =�� =)� =c] = =�r�<]��<��<��<Y�<Uc�<���<?K�<���<�B�<���<���<Z��<���<�.�<&��<�X�<?	�<��<���<[�<���<���<���<�"�<
f�<��<]��< ��<�k�<���<�c�<���<��<�`�<a��<7^�<��<���<#E�<��<�"�<W�<�k�<{o�<s�<^��<@��<���<T �<Y�<-�<���<r]�<d��<���<�S�<���<��<�)�<h��<���<[��<);�<O��<�^�<6�<���<�t�<��<vB�<�]�<�J�<g�<�ͳ<*��<�I�<�$�<+�<:�<+�<��<�Ӣ<��<@�<`��<a��<���<�'�<Q�<L͏<ͺ�<���<�t�<k�<��<�ց<!�}<��w<�q<|�k<��e<�q`<T�[<W1W<�WS<8�O</�L<f	J<=3G<�8D<s�@<�\=<3f9<�5<�0<�,<f�'<�(#<�<��<;�<}�<��<C`
<_�<y� <�i�;^n�;|��;i��;��;��;��;�t�;̰;@��;�;/˒;���;�Ex;ݫa;�L;�68;��&;:V;?�
;� ;���:��:f�:I�:��:'ȼ:���: ��:�U�:S�:��_:j�C:��+:a�:'
: !�9>��9�b�9E��9F6g9�#9��7 ׆��y��_�Ta���g��̭��b�ܹ����v`;�8�`��B��ܚ��ޯ���º�Һ�"ߺ�/纀��j�a�躈��.ຏ�ܺF�ۺ��ݺ����S���~���{�wy
�$�������(~�������#���)�Y�0�ϥ7�h.>���C���H�>%M��Q��QU�WZ��`��zh���q��|����-≻Xr���h��]�����������ໞ�$螻�q������'휻�  �  Ӭ=�=%�=�I=2�=ۛ=L7=��=	{=�-=�� =X� =�| =�> =���<m6�<In�<C��<���<��<]w�<'��<�x�<��<{�<\��<���<���<���<~n�<��<���<b]�<bA�<�]�< ��<mW�<1�<=�<�k�<8��<N��<B��<3��<���<�3�<���<`��<X-�<a{�<���<fV�<y��<�{�<��<���<g��<��<�>�<=S�<�i�<���<+��<5��<Q1�<iU�<�R�<`�<h��<'��<$��<ݗ�<"?�<���<ނ�<(F�<�1�<�L�<��<�<��<A`�<��<`��<�0�<�~�<��<���<:L�<���<���<^a�<�*�<:�<���<8�<�Ȥ<ړ�<(A�<�ԝ<�Z�<��<�}�<5�<
�<8��<��<�ً<��<vV�<�̈́<Q�<�S~<CMx<�6r<Y;l<��f<�-a<ON\<��W<WT<��P<~M<��J<��G<*�D<�nA<M�=<q�9<v�5<<
1<�h,<��'<6I#<1�<��<��<l�<O<�	<�.<�T <P��;�"�;���;���;���;�v�;�x�;tK�;���;ja�;`�;Ų�;���;�bz;�d;�N;X�:;�i);@;��;�b;���:{��:�o�:���:���:�V�:"�:��:�:�ł:��d:��F:k-:R�:�: �9e��9d��9���9a]J9��8�t7�䐸�>�7�R�9Ȃ�{p��<��Ȝι;����D�x4�hMY��)��$^���ꪺ�����-ͺ�4ٺ�F�yq庋��些Aມ(ܺ�ٺغ�ں�!ߺ3���b��]�C�	�����~������v��� �ï%���+���1��Z8�?L>���C���G�d�K���O���S���X�]�^�v�f��p�
�z�*���)����+�������C'���:���W��M���KE�����8��  �  .�=��=��=�p=� =[�=�T=i�=
�=,)=�� =q� =�P =o =�}�<���<��<8`�<��<��<��<��<���<�J�<���<"�<�M�<�H�<��<��<En�<p�<���<���<���<N�<9��<���<ٶ�<���<C�<:4�<�H�<E6�<s��<&��<|��<+�<c�<���<*��<wC�<���<&2�<G��<��<}z�<ܾ�<���<� �<VT�<���<���<x.�<yu�<I��< ��<�h�<8��<5)�<�)�<p��<ۭ�<,X�<��<���<���<h��<�*�<J��<�(�<���<�s�<�<ׄ�<�Ѽ<j�<�ָ<�<|@�<9ݱ<%~�<�,�<��<ٽ�<ꔦ<�f�<�)�<�ٟ<�y�<��<ȷ�<�o�<uB�<D/�<�-�<�/�<z$�<%��<飇<��<�b�<�<�y<Fs<�5m<#�g<qRb<Oy]<�Y<�$U<��Q<�cN<�`K<=kH<\E<�B<�t><R|:<.-6<��1<��,<o(<?m#<x�<�q<H"<��<~<�	<w`<�L�;���;S��;б�;.@�;�1�;<_�;i��;r�;�ղ;}��;H��;U��;9�;�~};q�g;m�R;gE?;��-;�;�;�;M�:��:iH�:��:��:'�:U�:aި:.K�:��:�]k:NK:%.:�j:>� :$�9�:�9.<�9��j9k}9k �8�}%��;��Z;�;�B� �k�j؈�����������Ag
���)�ЊN��xv�豏�Pf��w1���=ĺB�Ϻ�غڝܺQ�ݺ��ܺ��ٺ�^ֺ[�Ӻ�Ӻ�պT5ں�V���캤��A��J������b������������#���(��c.��4�Ȩ9�V�>�C���F��	J��ZM��4Q��V�g]\��-d�ptm���w�t��7���{8���␻f̔��֗����.��Ĥ��T����
�������  �  z=�=��=-�=9G=
�=
r=%�=��=�=z� =d =� =���< ��<MI�<���<��<�{�<��<���<�H�<���<���<^�<�p�<���<>��<?q�</�<���<5��<�}�<4}�<Q��<�	�<��<�^�<�J�<)W�<�t�<���<���<���<9C�<���<e1�<o�<���<Q��<���<@�<=l�<���<.�<z��<���<�;�<���<_��<-�<���< ��<�b�<J��<)��<>��<ٺ�<l>�<���<Q��<�i�<0�<=��<O��<���<��<���<���<R@�<���<�J�<���<k�<ܾ<�%�<�?�<@)�<�<���<M�<p��<�"�<���<�k�<)$�<�ߣ<ʘ�<�K�< ��<J��<�u�<NQ�<�E�<�O�<�c�<�s�<o�<�F�<���<yj�<��<��<X�y<*t<#hn<z�h<@�c<$�^<ӉZ<6�V<��R<�uO<KL<�4I<F<��B<�?<
;<Z�6<W,2<�W-<j(<5#<W�<��<8a<�<f_<��<zE<5f�;c�;���;Y�;!i�;o��;�A�;l��;9��;>��;5��;�Ơ;�F�;�o�;'��;z�k;�vW;��D;��3;$;K�;��;�;�N�:���:���:!��:��:�:`��:M�:��:��q:sN:��-:��:���9>"�9ӳ�9ʀl9�b"9��8�7+�B���ϸ��2"6��R��pp���������7ιy �*���C�N.i�����KK���ު����Bĺ�o̺�ѺG�Ӻ��Ӻ�8ҺW�Ϻ)κ��ͺs#кtJպhwݺ�N����s�a�o�����A�%���#��y(��T-�K2�+7�O�;���?���B��E�iEH��'K�R�N�-�S���Y���a�	�j���t��f��섻�Չ�8��{�~攻0���}���9���i��	B������  �  Q%="=�=�=pc=��=�=�=A�=n=�� =�& =p��<[��<+9�<6��<��<~��<w.�<J��<Y��<a�<��<���<:O�<>��<C��<���<��<*��<Z�<5�<�)�<�>�<z�<��<je�<*�<7��<��<���<���<]��<N��<�|�<
�<�h�<���<���<h��<���<���<=
�<�C�<���<%��<�9�<{��<���<�o�<Q��<w�<��<u��<D��<#*�<�0�<N��<�~�<���<���<���<D��<���<�q�<5a�<�c�<�{�<6��<���<=V�<���<�E�<½�<x"�<Lf�<�~�<vg�<�!�<*��<V-�<e��<�<�y�<���< ��<�8�<C�<���<�^�<�0�<��<��<�4�<�\�<�<ޣ�<���<�}�<�(�<��<��<�6�<�z<<,u<��o<gj<_e<��`<�)\<�X<-(T<��P<1M<��I<5�F<F;C<��?<=�;<�@7<�2<��-<��(< j#<�K<�H<g<ۥ<��
<i<��<��;��;J`�;`��;�B�;��;���;\X�;�a�;ʹ;ԍ�;Ͱ�;~^�;Qь;�K�;�!p;L�\;x�J;w�9;��*;��;�0;�\;9 ;��:���:]��:Q��:v!�:��:�=�:���:��u:�O:��*:�&	:P�9�d�9�=f9��9���8���6͚P��ȸ^�v9!���2���B�m�X���{��3��oտ����c1��9��\����V�����������%��bg��Pź��Ⱥ�ʺ��ʺ��ɺnaɺ�ɺ�s̺�Ѻ�ٺ����P�� ��_�l��+�h��{�#��	)�N.���2�,/7�>!;��z>�9.A��QC��'E�2G���I�M���Q�RX���_��h�)r�� |�ς�:I��eK���������ޓ�ꇕ�k����?��烗�*����  �  �:=�!=k�=|�=�m=a=��=- =Vp=A� ={Y =��<U��<��<�m�<���<�e�<4
�<r��<=��<8|�<�Z�<*�<��<d�<y��<���<b��<t��<���<���<I��<C��<{�<�M�<Բ�<�1�<���<j�<~M�</0�<��<��<���<̒�<,�<�|�<���<ڻ�<���<��<ʎ�<v��<T��<��<2�<p�<���<n]�<���<Y��<YD�<	��<,��<���<�@�<�I�<�<���<���<��<�*�<�+�<�)�<�*�<u2�<A�<�W�<Zy�<Ϩ�<n��<A:�<M��<��<�I�<���<♻<���<�9�<�Ŵ<�-�<o��<�ʬ<��<�y�<��<�x�<�<�ԝ<���<��<���<�̕<��<�L�<ǉ�<Y��<G��<O��<�<�<\��<�#�<ct�<�{<�%v<��p<��k<�g<�Qb<��]<˅Y<�rU<J�Q<�M<�vJ<�G<�|C<��?<K�;<�n7<�2<'�-<N}(<u#<չ<�h<�;<�;<Lj	<��<!X <y:�;�9�;|��;���;ë�;��;���;��;霽;�
�;�ի;m�;@�;�ڍ;'Ѓ;�=t;5�a;��P;�l@;Ό1;�#;"�;��;��;��:a��:���:)��:�O�:�7�:VV�:&Î:W�u:��L:��$:ּ�9��9�s9��94B;8�5��B���t���#���4���;���=�}�B���Q�H<r���lp��գ�׵��22�zR���q�Ko��z{��0柺����j����6�������ĺXRź�Fƺ��Ǻ%�ʺ^к��غ�㺋��a� �3?	�m���:�'�!�V�(��/��j4��9���<���?� B���C���D�
�E���F��I�oiL�w-Q�idW���^��Kg��4p�('y�$܀��τ��]��)����>�����������X=�����~����  �  �?=�=��=!�=.c=��=�z=�=�N=�� =0 =X�<��<�E�<A��<��<۫�<�m�<�M�<�B�<?�<�2�<j�<���<�N�<$��<���<u��<7��<���<��<2�<gk�<Ÿ�<��<	~�<@��<r�<��<B��<cj�<Z7�<��<���<��<9
�<�g�<2��<^��<�~�<R�<�#�<��<��<��<�B�<՚�<��<���<ya�<�(�<���<ǻ�<{f�<���<�.�<S8�<��<��<���<�8�<�f�<y��<���<���<
��<��<.(�<�9�<�L�<�i�<G��<���<6�<�L�<�{�<���<`r�<)�<���<��<�I�<Dx�<���<�<:8�<���<=D�<k�<%�<h�<|�<f�<��<[�<�g�<,��<[��<�x�<�(�<�<�)�<3��<�|<r�v<�	r<c>m<`�h<�c<�a_<~�Z<q�V<jzR<>�N<��J<�G<isC<��?<��;<lI7<*�2<n�-<h&(<��"<S�<�`<0�<&�< �<4<�`�;�;�;T��;��;�
�;Ŝ�;�!�;�\�;P�;O0�;&��;e�;G�;�-�;~s�;���;�w;uf;[V;߇F;R�7;��);Z�;��;�x;=�:L_�:���:x�:��:���:�ڟ:��:�`q:�eF:;�:���9i�9F�9?38|p�|5���<�v^�6�l�=�l�xFc�N~X�bT�P�^��}��8��K��4���!H/��K��df�k�~�;��e��y��T����d��h��FM��.뾺9eºz.ź�Ⱥ9�˺�Ѻ��ٺ6%��C���������*��(�&���.��w5�n";�V�?���B��E�$CF��F���F�\G�V�G��I��M���Q�!�W�,_��g�w.o�bw�Mw~�����妅�`s�����L���"̏��ԑ�싓��	���  �  �5=R	=��=ژ=tF=��=�[=��="=�x =`��<�n�<*]�<�w�<���<XB�<���<���<���<g��<���<'��<V��<��<��<'s�<���<���<���<
�<D�<���<��<�V�<���<�0�<���<�<�q�<���<ϊ�<5�<���<3��<�I�</��<!.�<[�<�Y�<�1�<|��<��<�l�<�H�<H�<2r�<���<�N�<	��<���<1��<���<�n�<�&�<~��<��<��<���<�i�<���<r8�<���<���<o �<�g�<���<���<J��<���< ��<j��<r��<���<��<	0�<P�<vY�<>�<��<�w�<�˱<���<��<V&�<bF�<��<R�<r�<�1�<m#�<�C�<[��<��<�a�<�Α<&�<�Y�<\b�<�=�<��<戅<;�<V��<�S|<�w<I�r<Nkn<��i<�Xe<�`<$\< �W<<(S<D�N<m�J<��F<�(C<�G?<7;<#�6<K"2<7-<�'<��!<<F<�<u3<�<�c<��;�>�;)�;�z�;5E�;�/�;���;�P�;��;R4�;Ƭ�;��;�H�;9��;���;ֺ�;�yz;�Wj;��Z;��K;7=;X�.;�,!;nG;�;sM�:��:���:��:�d�:j�:t �:FJ�:Pi:��<: �:���9c�[9z�8��v�5�$��.p��5��޲��Ƙ��P���A�������pu��d|��錹������̹����wo���/�$'H�|^�8�q�����������������r]���!���J��kQ���!����ź�9ʺ��κպ%�ݺ��躎��t�M������"�b�+��_4��;�G�A��F�I�H�-eJ���J��RJ��I�BUI���I�P�K���N��S���Y��~`���g�>o�M�u���{�)ƀ��Q���ǅ��C��ӊ�k������A>��2<��Fꕻ�  �  "=��=˳=0r='=^�=%3=Y�=�� =�> =�< ��<���<A��<��<݋�<H�<h4�<E�<Bh�<c��<��<7��<A<�<��<�&�<�f�<��<}��<H�<nb�<y��<�O�<���<�R�<���<:�<�q�<���<G"�<��<� �<��<�b�<���<-��<��<��<>�<���<	��<s0�<���<���<�<��<E�<)��<�X�<S:�<_2�<�,�<��<���<W`�<��<7��<E��<e+�<��<�$�<���<��<�s�<���<-�<�a�<"t�<g�<E�<��<t��<���< ��<���<c�<�<��<���<�+�<�z�<���<N��<!��<鲥<Kۢ<�.�<E��</x�<�s�<B��< �<�x�<_��<bt�<�ҏ<��<��<H�<Y��<]J�<��<���<`x|<�x<7�s<Zo<��j<Zf<��a<_]<�TX<�S<�O<\�J<a�F<��B<Q�>< �:<�A6<��1<�h,<��&<� !<�,<+5<�a<O�	<1�<7��;�5�; ��;���;\�;&t�;&��;��;���;��;A�;-h�;Zy�;�Y�; K�;��;�$�;�o|;TYm;׵^;5P;'�A;3;1�$;Ҿ;��	;1��:S��:e��:���:b��:x�:��:�<�:p�^:1:E�:�;�9\9��]����� ����������Ĺ���������㤹3���)|��w������b��c�߹������2��<G���X��g��Su�jn���ٕ��V�����⯺�+��?$����Ǻa�ͺ�?Ӻ�ٺmg����	��д�y��uB��&�-\0���9��sA���G���K�adN��UO�	O���M�B�L��L��bL��N��SQ�V��[�1gb�'i�-vo��:u��Jz���~�Yx��;�������ݤ��҆���|���T���ᓻ����  �  �=��=�=�K=��=�=\=�p=�� =� =���<�S�<?%�<<-�<�s�<��<���<d��<���<`�<22�<�E�<�1�<b��<px�<O��<q!�<�_�<���<���<�p�<���<��<�/�<s��<�+�<��<���<i��<:=�<^��<D�<D��<�"�<���<P5�<���<,��<��<���<�,�<���<�h�<u#�<V	�<
%�<|�<�<|��<���<6��<���<.��<b��<%�<_�<Vk�<<@�<k��<)��<�	�<���<p �<���<f,�<���<���<���<t��<A��<�O�<A�<���<���<�̾<�ϼ<�ɺ<��<�]�<u߳<,�<�J�<�I�<�<�<�9�<�T�<ꞟ<j"�<`�<[�<�"�<݋�<X�<���<�<�<6��<+��<a��<�]�<��<
��<�r�< �|<�Dx<%t<	p<��k<�Vg<a�b<?�]<��X<a�S<3O<X�J</dF<�DB<�2><�
:<��5<��0<e�+<�D&<�l <�b<jP<�`<$�<�|<n�;���;�V�;l��;���;��;�,�;�2�;���;�~�;���;-)�;/V�;�j�;n��;@�;R�;c�};�ro;xa;F\S;��D;6�5;�';}h;��
;7��:n��:i��:��:-�:��:s�:�v~:�dT:l_&:m��9��9���8F���/�]�6	��(�˹��แ
�2�޹�Ϲ|���i�������ʥ��P��%�ι�]������"���6�k�G���U��@a�	�k���v�sU�����D��� $��'�����&���S�ɺT�к%�׺^�޺�N�ښ��} ��@	�$W��G��t)�`04���=���E�A4L��sP���R��ZS�i�R��,Q���O�ǲN�X�N�y�P���S�rX��"^��Rd�{j��'p�Uu�I?y���|�d%��X��BT��U�� +��%{��~������b���  �  ��=ط={v=�/=��=�p=1�=S=S� =���<#`�<� �<���<b��<}�<��<�g�<g�<���<C��<,��<�
�<���<w��<?�<^��<���<6�<���<F��<uu�<{�<��<�f�<��<�k�<��<���<�<MJ�<ӎ�<���<�h�<���<���<���<�V�<#��<m|�<;F�<k��<`��<��<T��<Y��<���<��<���<�~�<)u�<J��<"��<&��<�L�<��<z&�<�3�<?�<���<L\�<���<[��<�-�<���<>]�<c��<^�<�"�<)�<��<l�<��<���<���<��<'��<���<�q�<�%�<��<��<}�<��<���<�<��<�B�<nÜ<��<���<NΖ<�>�<5˓<+^�<'�<vE�<}�<r��<jf�<)�<Cބ<̖�<H_�<�}|<�gx<�lt<�kp<�Bl<q�g<m'c<'8^<�'Y<eT<W7O<֎J<�&F<�A<��=<��9<y65<$z0<�W+<q�%<��<9�<_�<@�<2<�<���;�i�;���;;T�; b�;���;�*�;G<�;���;���;��;�D�;���;���;�*�;7�;�]�;Gb~;m�p;�c;�CU;X�F;��7;�v(;�Y;d;�"�:�7�:H�:ി:��:s�:�i�:�w:��L:�:�k�9`Bp9F8�7��@Ņ�8���ɰ�j���ڑ���l���}�̹ޠ��Q[��kT��c�¹(�ܹQ���ص���'�c�9���H�GuT��]���e���o�G�|�������_v��$_��$���i�ºR�˺��Ӻ}�ںU�ẓ���8��\O�u��C�u[ ��+�1�6�]�@���H��,O�eS�b�U���U��U�2VS���Q�X�P�]�P��\R�$�U�2Z���_�/�e���k���p�!u���x�5�{�`�~�����R�����fZ��L医fs��S���ħ���  �  ��=�M=I=��=׬=�O=��=2(=b =��<�M�<���<u-�<r�<�B�<W��<���<� �<��<��<v��<���<&��<��<��<1�<U�<��<P��<�O�<��<���<��<���<3��<��<�>�<G�<�1�<��<))�<�h�<��<s��<)@�<���<�s�<��<F��<�d�<*��<m2�<T��<���<c��<ɪ�<�
�<	��<}��<�"�<���<^��<w&�<��<���<P�<n��<_��<IB�<���<�j�<x'�<1 �<x��< ��<�H�<���<���<J�<Ҿ�<�<�n�<���<A��<���<ꑼ< ��<���<tv�<���<�3�<;!�<$ת<�p�<��<�Р<�ם<Z6�<p��<C�<���<�?�<0�<H�<&��<��<H�<�:�<��<���<� �<Gʁ<	><	Q{<շw<�Bt<�p<k�l<�}h<��c<�L^<j�X<sS<�M<ŀH</�C<��?<��;<8<�4<x/<�X*<Ϝ$<hW<�<R�<@
<��<��;���;Q1�;�A�;���;6��;��;T�;$��;��;�<�;�ѳ;���;�"�;×;0�;��;�;`s;�tg;�I[;@N;�|?;�^/;�4;��;�#�:'�:���:��:���:�V�:|��:��h:�F:�4:P��9YQX9�~;�vk��p۹S���R6��H��%M���F���7��$�L������	깇�繝M�������"���:���P��b��/l��o�sho���n�;rq�U�z��"��Jᒺo�������.ĺ�LҺ��ܺi�ܛ�QG��W��Ĕ��C�����G,��'�A�4��)B�s4N� X�]�^���b���c�'5b���^���Z���V��$T��kS��U���X� �^�.�e��l���r��w�B�z��?|�Z�|��}��������>󄻕ֈ�7V��y����U������  �  ��=�]=N/=)�=I�=S`=b�=�7=(r =1�<�s�<3��<WZ�<$7�<�q�<��<�<�I�<��<�;�<Q��<���<���<[��<i�<�U�<fx�<��<���<�_�<��<���<���<���<�l�<���<O(�<q6�<�)�<N�<�4�<�}�<m��<@��<�d�<��<��<\��<r��<��<���<�U�<S��<�#�<���<���<�9�<���<��<KJ�<O��<�<�E�<[<�<l��<�(�<��<C��<�c�<���<��<;3�<��<��<1��<�1�<F��<��<4�<k��<z�<�r�<p��<���<��<߳�<�˺<E˸<���<��<�Q�<C@�<��<���<�5�<���<��<te�<Z%�<�D�<��<wf�<N5�<%�<ڴ�<q0�<Ii�<^�<��<���<�A�<b�<�d<#d{<3�w<�-t<=�p<�l<�Ih<oc<&&^<b�X<"S< �M<��H<�$D<@<�7<<�^8<\F4<�/<*�*<��$<��<��<56<�
<�Q<3G�;4X�;1��;L��;�4�;�@�;r��;��;�s�;%�;�ż;ec�;�;�;!��;!C�;hX�;IA�;[�;Es;�g;�Z;1`M;��>;?�.;s�;T�;�E�:2��:�C�:G��:�:���:�ׄ:�&m:�J:$!:���9��h9S�6��W�n�й��go0��5B��iG��fA��2�H��z��,��~@��߹���^9�XH���6�VM�8G_�	�j�J�o��Sp�9�p��-t�K�}������,���|�����T�ú{^Ѻ�ۺ?��lk���뺧�}�����b��}.�V&��3���@���L�o�V�e�]��ka�hb���`���]�-�Y���U��+S��pR�<T���W�5�]���d�P�k��r��)w��tz�9F|�ZR}��~�Cf���`��ER���!������L��Z4�������  �  ʼ=��='_=�/=�=�=	=b=$� =Y��<��<!A�<���<���<���<���<B��<��<�!�<��<'�<B�<�D�<v �<w�<���<��<'��<')�<���<��<���<}��<<z�<L#�<��<p��<J�<R�<O �<�R�<��<�L�<x�<K��<�r�<8��<1�<)'�<7��<�V�<��<|�<��<�W�<qa�<���<!x�<�{�<J��<1�<g�<4��<ԏ�<W5�<���<�|�<3�<���<�7�<��<�Q�<��<���<i�<���<j1�<�1�<0��<��<���<�y�<F�<C��<a�<��<�)�<r'�<��<�o�<0��<���<�R�<��<���<�w�<���<F�<���<Tŗ<.�<SҔ<떓<,^�<+�<(��<oÍ<���<�{�<��<̛�<|0�<_�<g�{<1�w<5�s<�p<kl<'�g<�b<��]<�LX<��R<!�M<� I<�D<��@<v�<<19<��4<�h0<w@+<�%<XG< �<�
<%�<�R<yh�;,��;E�;.��;l
�;���;$�;g@�;���;>��;�:�;��;,ˬ;�9�;2��;Ip�;��;W�;��r;�e;��X;k&K;k<;��,;,;ǽ;�s�:���:'��:{��:Y��:4Ǘ:��:��x:q�U:3�+:�F�9��9�^8n� �t�����h�.$1�P7��)2��%��)��Q �q���͹��ɹ��ع���.�:+��PC���W�of���n�W]s���v�{|�N���NR�����%;���)��96ú�κ�u׺Hݺ�������.�Q������w1��{�Q/#�x0��]=�>�H�ylR�b9Y��3]��f^�,3]��LZ���V�S��P���O�6<Q���T�z�Z�υa���h�l�o�Ջu��y�\r|�|Z~�!"��������Rp��%�����O*���ᕻh蘻�  �  ��=3�=��=Zp=C+=��=iA=Ϛ=}� =} =Vv�<0��<L��<-��<}��<a�<�A�<Re�<��<	�<�x�<ֲ�</��<Sw�<���<�8�<�V�<�g�<P��<q��<3+�<M��<�f�<��<���<��<2q�<E��<D��<��<}w�<��<Ѷ�<3��<gG�<���<l�<0��<G��<8L�<a��<uD�<l��<�P�<��<3�<��<z@�<[2�<�Y�<���<���<y�<8��<إ�<q��<���<!��</7�<j��<.�<]v�<���<���<N�<u�<$��<1��<J�<4,�<���<z�<wJ�<�D�<�_�<ވ�<6��<t��<hb�<Uݴ<&�<��<lѫ<���<OK�<M2�<�T�<���<�}�<���<�ߖ<�o�<�!�<[ڒ<��<���<c:�<�:�<���<\��<<�<W��<,�<��{<g�w<\ps<1^o<!&k<�f<��a<��\<9�W<_�R< �M<{I<�mE<8�A<"�=<N:<%�5<P1<,<{d&<l8 </�<j?<��<>�<eY<���;�Q�;���;6��;�Q�;�D�;*/�;Z��;Gc�;�)�;��;�;�J�;��;8�;��;��;T�q;��c;=�U;OdG;�8;�");s};6
;��:pa�:��:`W�:���:k�:z�:W#�:Lwd:d
::\�	:�{�9�r�8�%������ѹ����]���<����Q�e��ù��?��뛺���ع����i���5��M�KEa��jo��Ky�v���N������k ��4���-��$�����º�˺��Ѻ�1ֺ��ٺ��ݺ�G��Y�!���f��p�� %�v�+�/%8�C��L�-�R�?�V��HX��W��oU��QR��6O�s�L�\DL�ƗM�Q���V�y]��e���l��gs���x��}�	!��ɡ���\�������S��񔋻(�����������旻�  �  h=� ='�=4�=wg=��=�w=�=C=ZU ='�<���<y��<��<��<�^�<v)�<�.�<�`�<��<���<�!�<�"�<S��< o�<���<���<���<���<��<�&�<���<���<�z�<=��<=l�<c��<�'�<&��<c��<���<IK�<��<���<���<rp�<���<��<�<��<1W�<��<ou�<@+�< �<�6�<���<
7�<��<{�<^=�<�h�<��<i�<��<�j�<�r�<\/�<s��<�<�K�<��<��<�3�<���<���<���<���<���<e��<���<�h�<nm�<��<�ɿ<k�<-"�<��<�Ϸ<eE�<�z�<{�<LY�<:-�<��<L�<�O�<�ǝ<[��<{�<���</&�<�<�\�<��<�i�<2��<<���<��<��<���<�k�<��{<r2w<^�r<�En<��i<YBe<ь`<��[<��V<�MR<��M<��I<�$F<r�B<��><@;<q�6<o,2<��,<�C'<33!<��<У<4�<ֻ<�b<��;W]�;V��;��;��;��;�1�;���;�0�;@�;���;� �;�`�;lc�;d�;}��;���;6p;fU`;�Q;EB; $3;/$;4�;ص;u��:^/�:>��:4 �:;��:,T�:�:���:��r:t�G:UX:c��9[6M9XlX7R�F1��v�ȹ""�c���d�����ŒڹBt��bu��[��������p��>Z���i�W���=(��;D�Fm]�fNr�g���Q���N������t��}���Y�������uú�ɺ �̺*$Ϻ<�Ѻ�պ��ܺ�+纘����;��������&���1�p�;��.D�pkJ�S�N��P�>Q��O�:�M�3:K��iI�
�H�1J��ZM�%�R��oY��Ua�ېi��sq�)tx�CU~�y����̓�\����X������Ѝ�C���mH��El��
 ���  �  �>=N-=u= �=�=q&=��=!�=�M=�� =���<��<���<ʥ�<6��<yr�<[!�<���<t�<�*�<�U�<s�<�n�<8�<Y��<��<�6�<V0�<v�<��<P�<N"�<�`�<p��<Q�<o��<G��<�{�<��<ȼ�<0��<�v�<�k�<�X�<L)�<s��<�3�<z^�<HQ�<s�< ��<�u�<d3�<��<�<�R�<%��<B�<l��<4��<���<&��<��<Y��<tY�<*��<���<���<�<�O�<�t�<���<���<޹�<R��<\��<,�<��<��<N�<��<6�<r�<���<z�<�Y�<�z�<yh�<�<��<�Ų<�֯<�Ѭ<�˩<�ئ<z�<``�<g�<���<c�<���<�ݖ<lJ�<̓<�M�<���<���<m�<���<o}�<�<�B�<ӎ�<��{<��v<��q<��l<v#h<_yc<��^<�BZ<��U<k�Q<,�M<�J<�F<�3C<k�?<�;<N�7</�2<:�-<��'<W"< <�<c?<��
<��<�� <���;���;�d�;���;���;K��;���;I~�;d�;to�;(��;z��;ZӞ;�k�;��;!�;kpm;m�[;!5K;�i;;VG,;��;�S;
;���:{3�:���:9#�:'��:ѓ�:��:��:@V|:��Q:'�#:��9Y�9Zg�8N ��F#�߹����������2�ùH���]?�����Tx���!��ڒ}��#���̢�EV˹o �Jd��E>�37]��-y������(��9����䬺ݴ�(��>º�ƺ�HȺ�4ɺ�ɺn�˺ҿϺ�׺]4�;,�ƺ�)	������!�Q�+��Q4�ޡ;�QuA���E�6�H��J��(J�R9I�0�G���F��}F�E�G���J��O�ujV���^��_g��dp�n�x��U��Ĳ��A���rQ��ߋ��Z��#����ג������Ǖ�d����  �  6H=�?=S%=y�=�=1=;�=�=%n=V� =>9 =^h�<���<���<��<���<��<_��<w��<J��<M��<��<p��<TN�<a��<?�<�`�<�R�<%�<-��<���<s��<ԥ�<��<��<̄�<��<��<Wp�<�X�<�^�<qt�<Z��<���<+R�<���<�L�<.s�<�k�<,F�<B�<���<���<*��<� �<�l�<<��<J�<,��<;��<R�<�+�<g�< ��<�j�<r��<��<��<�*�<�e�<�o�<-Z�<�8�<T�<��<���<���<��<3�<�@�<��<���<�K�<h��<�-�<"{�<K��<^��<*)�<2��<�޲<��<>(�<UR�<���<�<�m�<��<��<�~�<�l�<ǁ�<���<��<y�<�Ր<��<(+�<�<��<��<YZ�<���<W{<O�u<WPp<�k<�(f<bda<R�\<`|X<�kT<I�P<�0M<��I<a�F<utC<�?<
<<��7<{�2<ǳ-< 2(<$�"<�<�A<��<j�<�<�<�%�;���;i��;�.�;�Z�;���;n��;'��;���;��;YP�;@��;6x�;޸�;Љ;~;��i;�$V;�)D;m�3;�?$;�W;�	;ɱ�:�	�:��:F��:��:NV�:�^�:�Q�:鱒:�C:�cU:ݢ):�x�9�ժ9�+D9��8�؄��;���p�����?*��q������y���Pv�vs����9~���5����������>�1b�+q�����:����B������)���ú�*Ⱥէʺ�#˺�ʺ7�Ⱥ?�ǺDɺGKͺ2պ�����ﺑ� �SW
�9��I�r�%���,�I-3���8�g=��@�X{C�bE�b�E��E�F~E��E�G���I�n�N��U�;N]��f�.�p�߽z�m��(X������=�������P���3������j�������ǖ��  �  36=z4=�=:�=R�=4=��==�v=� =\v =Y =�b�<1��<D�<k}�<���<�i�<��<���<���<}�<�]�<�$�<���<�$�<�K�<:�<2��<��<G�<B��<~��<L��<�<�g�<���<���<K��<V��<I�<�?�<)h�<�k�<�:�<���<�$�<�I�<�K�<�>�<�5�<�B�<�l�<d��<]�<=p�<���<�9�<
��<��<ê�<�N�<
 �<b��<F>�<"��<���<���<��<�B�<�6�<q��<���<V\�<]�<���<0��<��<(�<�[�<���<�[�<���<C��<��<[^�<y�<�V�<>��<)l�<���<��<�S�<���<�0�<3å<�c�<a
�<���<�e�<\'�<m�<��<�.�<�n�<���<���<��<	�<��<L�<t:�<�K�<�z<P�t<I�n<�5i<��c<x"_<z�Z<�V<��R<�mO<�XL<|eI<gjF<q=C<Z�?<Q�;<;b7<��2<g-<�(<3�"<�Y<�9<KL<m�<_�	<|2<,� </�;oL�;��;�T�;�+�;S�;�}�;�X�;�;n�;���;�1�;n0�;�͈;��z;��d;c�O;�Z<;��*;Z�;�;�;LX�:���:[w�:���:�w�:�E�:�'�:f��:jh�:qkz:��Q:��(:Zo:"=�9q��9D�)9*U�8_�I7'�`�u���31��B^��{��5��\c�����^Ń�������1ǹ���I^��3D�دl�����Js�����建��ƺ-�κ��Ӻ��պxFպȐҺ!�κY˺\~ɺ*fʺ4�κqH׺�W��P򺬌��6
������;� ��R&��u+��R0�[5���9�e�=�4A���C��E���E���F�YH��K��{O��U�@�]���g���r��}�d���p���ڍ�}���t������=���Ø��̘�.^��eė��  �  }=�=��=i�=U^=��=�j=y�=�i=� =�� =XT =[ =*��<���<�Q�<˝�<���<hL�<���<Ns�<b5�<S�<2��<jd�<���<���<���<j��<�6�<���<4C�<U��<���<���<#I�<D��<���<���<�1�<Z��<���<��< �<���<u�</��<X��<7��<��<�+�<�o�<��<�Q�<���<�M�<z��<�<KG�<'��<���<4H�<���<�Y�<y��</<�<�a�<�:�<���< ��<4��<��<��<���<� �<$��<���<i��<P��<xm�<"	�<���<�~�<�-�<߶�<�
�<m�<@��<E��<�	�<qo�<�د<�V�<��<ʩ�<�o�<4�<H�<B��<{'�<b��<uc�<Z+�<��<5�<�c�<<��<���<���<�K�<��<M�<��<l�y<]Cs<�m<?g<��a<Q�\<�mX<_�T<Q<�	N<�BK<��H<a�E<�B<�?<�;<+�6<��1<ײ,<(�'<'s"<"�<��<�m<�<��<� <�I<m��;=s�;E�;���;���;U�;�0�;���;@D�;�ұ;Rq�;��;��;51�;�v;	_;��H;�b4;�M";��;e�;7��:P�::;�:*�:�::��:U˷:c�:.6�:D��:��n:J�G:]q":{Y:G��9S�9n�y9��:9+�8L5_8�v��B����&��a� N��W͐������_��w�����s[۹@�f/(��O���{��B��D˩��$�̺v�غ�w�AF�R;�:Ẻ�ۺ��պ��кOκ�)Ϻ�Ժn ݺ�`�����F~��P�g	�W��� ���$��I)�J6.���3�V9��?>�Q�B�+�E���G���I�r[K�=	N�61R�AX��\`��Rj�{�u�$񀻆��*�������nە���m������$��т��bw���a���  �  |�=I�=M�=�{=W=��=�/=��=�M=�� =P� =� =�W =� =��<2��<�&�<DH�<:s�<��<p2�<���<���<�B�<���<Z�<���<��<g3�<3��<p �<3��<��<���<���<�B�<���<���<�&�<���<0�<i�<���<β�<�w�<\��<�C�<�k�<v��<��<�<}�<H�<F��<�o�<���<Fc�<ޡ�<���<d��<R��<�$�<�{�<���<\�<���<>��<c��<L�<;{�<jW�<���<9c�<��<�9�<��<g��<ޱ�<� �<���<H�<��<���<c��<tC�<���<J��<[p�<Q�<m��<�<�<�<�<-�<:��<h�<%פ<�<^=�<g��<�+�<k��<�/�<��<ޑ<�<f�<+0�<�#�<q܇<iO�<�|�<z�~<�rx<��q<ׁk<~je<��_<�Z<�gV<�R<emO<-�L<J<]�G<��D<~�A<X.><�:<�5<B�0<��+<��&<k"<(�<P<A<�.<7�<�n<ס<�7�;b �;r��;��;k��;D��;/f�;�
�;c�;��;�˦;2~�;r<�;�C�;R�q;C�Y;p@B;8 -;^;^�
;l%�:��:��:92�:i��:���:H �:�-�:�_�:ͧ�:���::H_:��9:wV:,2�9���9���9~��9#��9��S9�<9�t8����� �0{W������U��,ͱ�6����gŹ�+عZd�������5�`�^�RF���]���Ե��ʺ�IܺM��\����h��Q��po��޺�غ�պ�ֺ�mۺU���w�A���-���4���
�������L�#�\�(���.�r�5�t<�:xB��?G��J�X+M�\O�8R�+ V���[�:�c���m���y��.������돻�e��ՙ����[���/����^���>��y����S���  �  ۛ=�=w�=�==s�=*k=��=��=�.=� =:� =ũ =-� =�[ =@ =rn�<ބ�<��<%��<���<���<�j�<�<'��<�d�<���<f�<��</��<�;�<ۖ�<z��<g�<��<��<�o�<C%�<11�<���<���<���<���<6:�<�@�<���<�z�<���<��<�<�_�<{��<�x�<B�<��<���<�y�<��<�<��<� �<9��<���<�'�< z�<P��<�2�<�^�<BF�<���<��<���<*n�<d��<�<�{�<��<���<4��<�4�<���<P��<���<Ss�<C;�<ξ<�<:$�<`�<��<\
�<��<A�<��<��<�2�<�K�<�J�< �<�<@&�<+u�<��<�#�<���<���<,��<���<��<M��<�g�<��<�<*�}<�kw<ȿp<�+j<�c</1^<(!Y<A�T<�Q<
N<�mK<�I<��F<�C<W�@<�==<� 9<\�4</�/<��*<M
&<��!<{a<�<��<U�<��<hu	<��<���;& �;�Q�;�(�;���;K]�;`��;��;;s�;x6�;+�;�Κ;���;�i�;��m;��T;V�<;�&;��;�3;��:��:���:!M�:���:�Ż:H�:\:�:��:ތ:Ou: �O: ,:M�:Z�9���9*�9�ʮ9���9�o�9_�O9�&�8�g7�aԸ��V�Ԓ���޸��E͹�ڹ(��m��(K��#���C��m�4���W�����/uֺ@��|(��P���������D���R(����aCߺ$ܺ�Mݺ�����w�������e
�����L��WX�v��}&������$�~�+�6y3�~;�#�B��I���M�+�P��^S��V���Y���_�jJg��Sq��E}�g>��'�������`�����Z���;��'���V������>מ�V4���  �  �q=u=�S=�=�=q;=��=d=3=�� =h� =b� =u� =� =>< =B��<S��<���<��<p��<���<h�<q��<�`�<0�<���<��<���<Hl�<���<6�<��<>��<9��<���<���<b��<���<{�<{��<�$�<ҝ�<���<9��<���<]�<�`�<x��<M��<0 �<���<�o�<(V�<�D�<��<���<�+�<aR�<�C�<��<���</��<���<�'�<;~�<$��<���<���<�|�<���<��<��<�f�<\��<���<�|�<o>�<�N�<U��<EW�<3�<?'�<6�<��<�u�<¼<�ĺ<V��<�!�<��<�F�<�<(��<��<�M�<0�<���<�g�<6�<`c�<��<�Θ<j�<#��<�@�<�,�<G<�<Q�<TK�<L�<��<]��<D}<u�v<k�o<�Di<o�b<�$]<�X<2�S<�P<�!M<]�J<CH<��E<=C<y&@<��<<�a8<�3<B�.<�$*<�{%<5)!<-<<�<1<�u<�~<
<(<��;���;Wo�;���;G�;�=�;k<�;̤�;��;Ϭ;G��;���;�;�;��;�j;#sQ;,/9;�#;#�;  ;��:v��:��:��:4E�:���:T�:��:q�:� �:nVi:kD:Q�!:�:��9,��9��9�-�9��97�9%u9V�9!!8yu����Y��A��''ȹ���1I�0��;�����-��uN���w�e瓺ܙ��Ǻ�޺��x����&�X ��E��V���F��
`�=���k�p�������̠��]�� ��������q���r�JB�*�Bb�ܱ"���)��92��;�UgC��mJ���O�~S�VV��%Y���\�tPb��i��s����絆�ɬ��$b���W��^"��Q~��+T������㣻GC���R������  �  b=^e=OC=(�=Ě=�)=�=0W=k=�� =�� =N� =� =ċ =�H =`��<��<w��<I��<t|�<��<6�<X��<w<�<���<t_�<i��<<��<M�<4��<1�<�^�<���<i�<�_�<ҷ�<Cs�<ʉ�<T��<Cq�<:�<'~�<���<R��<)��<���<�;�<�l�<!��<��</��<yk�<�[�<@S�<�1�<���<�D�<�g�<�R�<��<V��<���<���<
�<P[�<��<��<S��<�[�<���<�e�<���<B�<z��<,��<�M�<�<x�<���<\+�<�
�<��<U��<M¿<�U�<���<���<2c�<a��<���<*�<��<l�<9�<lV�<ߏ�<.��<<��<��<gw�<4��<�Ҙ<Q�<0|�<r(�<�<D�<-�<�(�<��<�k�<���<�}<�lv<Q�o<��h<�b<�\<��W<XS<P�O<��L<LJ<G�G<S�E<��B<B�?<�D<<�8<6�3<ʹ.<�)<�G%<!<�,<��<�0<�<�<�F
<1X<��;���;u�;׭�;���;��;���;��;.q�;I�;�8�;0�;�;b��;j�i;�FP;��7;��!;�[;��:���:�?�:��:�:�9�:ْ�:6�:\��:�`�:�̈́:��d:)�?:B$:�:��9V��9ڑ�9�ڽ9�S�9�`�9K�9P� 9�"8!���0T[�����޹͹�������Ѫ�Jl�H����1�YR���{�����Wׯ�g|ɺ��ມ��#� �����k�Ț�����y��k�T��[_�������w.��O� � ������a��P�����+�p��"M����F�!�\3)�d�1���:��C���J�O�P��yT��rW�JZ���]��Yc��j�|�t��~���=���@��/���	��ܟ��:�����i��S���J٢��۠�S���  �  �q=u=�S=�=�=q;=��=d=3=�� =h� =b� =u� =� =>< =B��<S��<���<��<p��<���<h�<q��<�`�<0�<���<��<���<Hl�<���<6�<��<>��<9��<���<���<b��<���<{�<{��<�$�<ҝ�<���<9��<���<]�<�`�<x��<M��<0 �<���<�o�<(V�<�D�<��<���<�+�<aR�<�C�<��<���</��<���<�'�<;~�<$��<���<���<�|�<���<��<��<�f�<]��<���<�|�<p>�<�N�<V��<GW�<3�<A'�<8�<��<�u�<	¼<�ĺ<Y��<�!�<��<�F�<�<*��<��<�M�<1�<���<�g�<6�<_c�<��<�Θ<h�<!��<�@�<�,�<D<�<Q�<QK�<J�<��<[��<D}<q�v<h�o<�Di<m�b<�$]<�X<2�S<�P<�!M<`�J<CH<��E<	=C<~&@<��<<b8<�3<H�.<�$*<�{%<:)!<1<<
�<4<�u<�~<
<(<��;���;Qo�;���;>�;�=�;a<�;���;��;Ϭ;<��;���;�;�;��;��j;sQ;/9;�#;�;���:Ғ�:j��:��:��:.E�:���:P�:��:q�:� �:lVi:iD:Q�!:�:��9+��9��9�-�9��97�9%u9V�9"!8yu����Y��A��''ȹ���1I�0��;�����-��uN���w�e瓺ܙ��Ǻ�޺��x����&�X ��E��V���F��
`�=���k�p�������̠��]�� ��������q���r�JB�*�Bb�ܱ"���)��92��;�UgC��mJ���O�~S�VV��%Y���\�tPb��i��s����絆�ɬ��$b���W��^"��Q~��+T������㣻GC���R������  �  ۛ=�=w�=�==s�=*k=��=��=�.=� =:� =ũ =-� =�[ =@ =rn�<ބ�<��<%��<���<���<�j�<�<'��<�d�<���<f�<��</��<�;�<ۖ�<z��<g�<��<��<�o�<C%�<11�<���<���<���<���<6:�<�@�<���<�z�<���<��<�<�_�<{��<�x�<B�<��<���<�y�<��<�<��<� �<9��<���<�'�< z�<P��<�2�<�^�<BF�<���<��<���<+n�<e��<�<�{�<��<���<7��<�4�<���<T��<���<Xs�<H;�<ξ<�<@$�<e�<��<a
�<���<	A�<��<��<�2�<�K�<�J�< �<�<>&�<)u�<��<�#�<���<���<'��<���<z��<H��<�g�<��<�<"�}<�kw<¿p<�+j<�c<-1^<(!Y<C�T<�Q<N<�mK<�I<�F<�C<a�@<�==<� 9<f�4<9�/<��*<V
&<��!<�a<��<��<X�<��<hu	<��<���; �;�Q�;r(�;���;8]�;L��;��;%s�;b6�;�;}Κ;z��;�i�;k�m;s�T;9�<;��&;��;�3;ʫ�:ӄ�:���:M�:���:�Ż:H�:W:�:��:�݌:Ou:�O:,:L�: Z�9���9*�9�ʮ9���9�o�9_�O9�&�8�g7�aԸ��V�Ԓ���޸��E͹�ڹ(��m��(K��#���C��m�4���W�����/uֺ@��|(��P���������D���R(����aCߺ$ܺ�Mݺ�����w�������e
�����L��WX�v��}&������$�~�+�6y3�~;�#�B��I���M�+�P��^S��V���Y���_�jJg��Sq��E}�g>��'�������`�����Z���;��'���V������>מ�V4���  �  |�=I�=M�=�{=W=��=�/=��=�M=�� =P� =� =�W =� =��<2��<�&�<DH�<:s�<��<p2�<���<���<�B�<���<Z�<���<��<g3�<3��<p �<3��<��<���<���<�B�<���<���<�&�<���<0�<i�<���<β�<�w�<\��<�C�<�k�<v��<��<�<}�<H�<F��<�o�<���<Fc�<ޡ�<���<d��<R��<�$�<�{�<���<\�<���<>��<c��<L�<<{�<kW�<���<;c�<��<�9�<"��<k��<��<� �<���<H�<��<���<j��<{C�<���<R��<bp�<X�<t��<�<���<�<�<1�<=��<j�<'פ<�<]=�<e��<�+�<g��<�/�<��<�ݑ<
�<_�<$0�<#�<j܇<bO�<�|�<n�~<�rx<��q<Ёk<yje<��_<�Z<�gV<�R<kmO<5�L<J<h�G<��D<��A<g.><�:<�5<P�0<��+<��&<w"<2�<P<#A<�.<:�<�n<ԡ<�7�;U �;b��;��;S��;)��;f�;�
�;�b�;��;x˦;~�;T<�;�C�; �q;�Y;G@B; -;�];E�
;B%�:���:��:#2�:X��:���:> �:�-�:�_�:ɧ�:���:7H_:��9:vV:*2�9���9���9}��9#��9��S9�<9�t8����� �/{W������U��,ͱ�6����gŹ�+عZd�������5�`�^�RF���]���Ե��ʺ�IܺM��\����h��Q��po��޺�غ�պ�ֺ�mۺU���w�A���-���4���
�������L�#�\�(���.�r�5�t<�:xB��?G��J�X+M�\O�8R�+ V���[�:�c���m���y��.������돻�e��ՙ����[���/����^���>��y����S���  �  }=�=��=i�=U^=��=�j=y�=�i=� =�� =XT =[ =*��<���<�Q�<˝�<���<hL�<���<Ns�<b5�<S�<2��<jd�<���<���<���<j��<�6�<���<4C�<U��<���<���<#I�<D��<���<���<�1�<Z��<���<��< �<���<u�</��<X��<7��<��<�+�<�o�<��<�Q�<���<�M�<z��<�<KG�<'��<���<4H�<���<�Y�<y��</<�<�a�<�:�<���<��<5��<��<��<���<� �<'��<���<n��<U��<~m�<)	�<���<�~�<�-�<趿<�
�<w�<I��<N��<�	�<yo�<�د<�V�<��<ϩ�<�o�<4�<H�<A��<x'�<_��<pc�<U+�<��<�4�<�c�<3��<���<���<�K�<���<E�<��<_�y<RCs<zm<?g<��a<P�\<�mX<c�T<Q<�	N<�BK<��H<q�E<'�B<�?<�;<=�6<��1<�,<8�'<5s"<.�<��<�m<�<��<� <�I<b��;-s�;�D�;���;ػ�;�T�;�0�;���;D�;�ұ;,q�;��;s�;1�;��v;�_;y�H;�b4;�M";��;K�;��:.�: ;�:�:�:.��:M˷:c�:*6�:A��:|�n:G�G:\q":zY:F��9S�9n�y9��:9,�8N5_8�v��A����&��a� N��W͐������_��w�����s[۹@�f/(��O���{��B��D˩��$�̺v�غ�w�AF�R;�:Ẻ�ۺ��պ��кOκ�)Ϻ�Ժn ݺ�`�����F~��P�g	�W��� ���$��I)�J6.���3�V9��?>�Q�B�+�E���G���I�r[K�=	N�61R�AX��\`��Rj�{�u�$񀻆��*�������nە���m������$��т��bw���a���  �  36=z4=�=:�=R�=4=��==�v=� =\v =Y =�b�<1��<D�<k}�<���<�i�<��<���<���<}�<�]�<�$�<���<�$�<�K�<:�<2��<��<G�<B��<~��<L��<�<�g�<���<���<K��<V��<I�<�?�<)h�<�k�<�:�<���<�$�<�I�<�K�<�>�<�5�<�B�<�l�<d��<]�<=p�<���<�9�<
��<��<ê�<�N�<
 �<b��<F>�<"��<���<���<��<�B�<�6�<s��<���<Y\�<`�<���<4��<��<.�<�[�<���<�[�<���<M��<��<f^�<y�<�V�<I��<3l�<���<��<�S�<���<�0�<6å<�c�<a
�<���<�e�<X'�<h�<��<{.�<�n�<���<���<��<��<��<B�<k:�<�K�<��z<D�t<@�n<�5i<��c<w"_<|�Z<�V<��R<nO<�XL<�eI<xjF<�=C<n�?<e�;<Pb7<��2<g-<�(<B�"<�Y<�9<TL<s�<b�	<|2<)� <#�;^L�;��;oT�;�+�;�R�;�}�;�X�;ȗ�;C�;f��;q1�;F0�;�͈;��z;��d;+�O;�Z<;��*;7�;�;�;&X�:q��:Dw�:o��:�w�:�E�:�'�:a��:gh�:lkz:��Q:��(:Yo:!=�9p��9C�)9+U�8g�I7$�`�s���31��B^��{��5��\c�����^Ń����줢��1ǹ���I^��3D�دl�����Js�����建��ƺ-�κ��Ӻ��պxFպȐҺ!�κY˺\~ɺ*fʺ4�κqH׺�W��P򺬌��6
������;� ��R&��u+��R0�[5���9�e�=�4A���C��E���E���F�YH��K��{O��U�@�]���g���r��}�d���p���ڍ�}���t������=���Ø��̘�.^��eė��  �  6H=�?=S%=y�=�=1=;�=�=%n=V� =>9 =^h�<���<���<��<���<��<_��<w��<J��<M��<��<p��<TN�<a��<?�<�`�<�R�<%�<-��<���<s��<ԥ�<��<��<̄�<��<��<Wp�<�X�<�^�<qt�<Z��<���<+R�<���<�L�<.s�<�k�<,F�<B�<���<���<*��<� �<�l�<<��<J�<,��<;��<R�<�+�<g�< ��<�j�<r��<��<��<�*�<�e�<�o�</Z�<�8�<W�<��<���<���<��<9�<�@�<��<���<�K�<s��<�-�<-{�<V��<i��<5)�<<��<�޲<��<E(�<[R�<���<�<�m�<��<��<�~�<�l�<���<���<��<y�<�Ր<��<+�<�<���<��<PZ�<���<W{<B�u<NPp<�k<�(f<ada<U�\<f|X<�kT<T�P<1M<��I<s�F<�tC<+�?<&
<<��7<��2<۳-<22(<4�"<�<�A<��<p�<�<�<�%�;���;W��;�.�;�Z�;l��;I��;���;���;��;-P�;��;x�;���;�ω;�~;��i;I$V;�)D;B�3;v?$;�W;�	;���:�	�:ˮ�:4��:��:DV�:�^�:�Q�:汒:�C:�cU:ۢ):�x�9�ժ9�+D9��8�ׄ��;���p�����?*��q������y���Pv�us����9~���5����������>�1b�+q�����:����B������)���ú�*Ⱥէʺ�#˺�ʺ7�Ⱥ?�ǺDɺGKͺ2պ�����ﺑ� �SW
�9��I�r�%���,�I-3���8�g=��@�X{C�bE�b�E��E�F~E��E�G���I�n�N��U�;N]��f�.�p�߽z�m��(X������=�������P���3������j�������ǖ��  �  �>=N-=u= �=�=q&=��=!�=�M=�� =���<��<���<ʥ�<6��<yr�<[!�<���<t�<�*�<�U�<s�<�n�<8�<Y��<��<�6�<V0�<v�<��<P�<N"�<�`�<p��<Q�<o��<G��<�{�<��<ȼ�<0��<�v�<�k�<�X�<L)�<s��<�3�<z^�<HQ�<s�< ��<�u�<d3�<��<�<�R�<%��<B�<l��<4��<���<&��<��<Y��<uY�<+��<���<���<�<�O�<�t�<���<���<��<U��<`��<0�<��<��<T�<��<6�<#r�<���<��<�Y�<�z�<�h�<�<'��<�Ų<�֯<�Ѭ<�˩<�ئ<}�<b`�<h�<���<`�<���<�ݖ<fJ�<̓<�M�<���<���<c�<���<e}�<�<�B�<ˎ�<��{<��v<��q<��l<r#h<^yc<��^<�BZ<��U<v�Q<9�M<J<#�F<�3C<�?<�;<c�7<C�2<M�-< �'<g"< <�<l?<��
<��<�� <���;���;�d�;���;j��;+��;���;"~�;�c�;Jo�;���;P��;1Ӟ;�k�;v�;� �;-pm;6�[;�4K;i;;3G,;��;�S;�;c��:d3�:���:,#�:��:˓�:��:��:;V|:��Q:%�#:��9X�9Xg�8P ��F#�߹����������1�ùH���]?�����Tx���!��ڒ}��#���̢�EV˹o �Jd��E>�37]��-y������(��9����䬺ݴ�(��>º�ƺ�HȺ�4ɺ�ɺn�˺ҿϺ�׺]4�;,�ƺ�)	������!�Q�+��Q4�ޡ;�QuA���E�6�H��J��(J�R9I�0�G���F��}F�E�G���J��O�ujV���^��_g��dp�n�x��U��Ĳ��A���rQ��ߋ��Z��#����ג������Ǖ�d����  �  h=� ='�=4�=wg=��=�w=�=C=ZU ='�<���<y��<��<��<�^�<v)�<�.�<�`�<��<���<�!�<�"�<S��< o�<���<���<���<���<��<�&�<���<���<�z�<=��<=l�<c��<�'�<&��<c��<���<IK�<��<���<���<rp�<���<��<�<��<1W�<��<ou�<@+�< �<�6�<���<
7�<��<{�<^=�<�h�<��<i�<��<�j�<�r�<]/�<t��<�<�K�<��<��<�3�<���<���<���<���<���<k��<���<�h�<vm�<��<�ɿ<u�<7"�<��<�Ϸ<nE�<�z�<!{�<RY�<?-�<��<O�<�O�<�ǝ<Z��<{�<���<*&�<纔<�\�<	��<�i�<)��<䴌<���<��<��<���<�k�<��{<h2w<V�r<�En<��i<XBe<ӌ`<��[<��V<�MR<��M<�I<�$F<��B<��><R;<��6<�,2<
�,<�C'<A3!<��<ڣ<<�<ۻ<�b<��;Q]�;L��;��;��;ɗ�;�1�;���;�0�;�;���;o �;�`�;Gc�;�c�;\��;c��;�5p;5U`;nQ;B;�#3;�.$;�;ǵ;Z��:I/�:.��:( �:3��:&T�:�:���:��r:q�G:SX:a��9X6M9ElX7R�F1��v�ȹ!"�c���c�����ŒڹBt��bu��[��������p��>Z���i�W���=(��;D�Fm]�fNr�g���Q���N������t��}���Y�������uú�ɺ �̺*$Ϻ<�Ѻ�պ��ܺ�+纘����;��������&���1�p�;��.D�pkJ�S�N��P�>Q��O�:�M�3:K��iI�
�H�1J��ZM�%�R��oY��Ua�ېi��sq�)tx�CU~�y����̓�\����X������Ѝ�C���mH��El��
 ���  �  ��=3�=��=Zp=C+=��=iA=Ϛ=}� =} =Vv�<0��<L��<-��<}��<a�<�A�<Re�<��<	�<�x�<ֲ�</��<Sw�<���<�8�<�V�<�g�<P��<q��<3+�<M��<�f�<��<���<��<2q�<E��<D��<��<}w�<��<Ѷ�<3��<gG�<���<l�<0��<G��<8L�<a��<uD�<l��<�P�<��<3�<��<z@�<[2�<�Y�<���<���<y�<8��<إ�<q��<���<!��<07�<j��</�<^v�<���<���<P�<u�<'��<5��<O�<9,�<���<�z�<~J�<�D�<�_�<戽<>��<|��<ob�<\ݴ<-�<�<qѫ<���<RK�<P2�<�T�<���<�}�<���<�ߖ<�o�<�!�<Uڒ<|�<���<\:�<}:�<���<U��<5�<Q��<,�<��{<^�w<Vps<-^o<&k<�f<��a<��\<?�W<g�R<)�M<!{I<�mE<E�A<0�=<]:<4�5<P1<&,<�d&<x8 <9�<r?<��<B�<gY<���;�Q�;���;)��;sQ�;zD�;/�;@��;+c�;�)�;��;��;�J�;瀛;�;f�;���;'�q;Z�c;�U;0dG;��8;�");b};6
;j�:_a�:���:VW�:���:f�:w�:U#�:Iwd:b
::[�	:�{�9�r�8�%������ѹ����]���<����Q�e��ù��?��뛺���ع����i���5��M�KEa��jo��Ky�v���N������k ��4���-��$�����º�˺��Ѻ�1ֺ��ٺ��ݺ�G��Y�!���f��p�� %�v�+�/%8�C��L�-�R�?�V��HX��W��oU��QR��6O�s�L�\DL�ƗM�Q���V�y]��e���l��gs���x��}�	!��ɡ���\�������S��񔋻(�����������旻�  �  ʼ=��='_=�/=�=�=	=b=$� =Y��<��<!A�<���<���<���<���<B��<��<�!�<��<'�<B�<�D�<v �<w�<���<��<'��<')�<���<��<���<}��<<z�<L#�<��<p��<J�<R�<O �<�R�<��<�L�<x�<K��<�r�<8��<1�<)'�<7��<�V�<��<|�<��<�W�<qa�<���<"x�<�{�<J��<1�<g�<4��<ԏ�<X5�<���<�|�<3�<���<�7�<��<�Q�<��<���<i�<���<l1�<�1�<3��<��<���<�y�<K�<H��<f�<��<�)�<x'�<��<�o�<4��<���<�R�<��<���< x�<���<F�<���<Sŗ<.�<PҔ<薓<(^�<'�<$��<jÍ<���<�{�<��<Ǜ�<w0�<V�<_�{<+�w<0�s<�p<il<'�g<�b<��]<�LX<��R<(�M<� I<�D<�@<��<<;9<��4<�h0<�@+<�%<`G<�<�
<)�<S<|h�;,��;A�;'��;c
�;���;�#�;W@�;���;*��;�:�;��;ˬ;u9�;��;5p�;��;�V�;��r;��e;��X;V&K;�j<;��,;,;��;{s�:���:��:t��:T��:0Ǘ:��:��x:n�U:2�+:�F�9��9�^8o� �t�����h�.$1�P7��)2��%��)��Q �q���͹��ɹ��ع���.�:+��PC���W�of���n�W]s���v�{|�N���NR�����%;���)��96ú�κ�u׺Hݺ�������.�Q������w1��{�Q/#�x0��]=�>�H�ylR�b9Y��3]��f^�,3]��LZ���V�S��P���O�6<Q���T�z�Z�υa���h�l�o�Ջu��y�\r|�|Z~�!"��������Rp��%�����O*���ᕻh蘻�  �  ��=�]=N/=)�=I�=S`=b�=�7=(r =1�<�s�<3��<WZ�<$7�<�q�<��<�<�I�<��<�;�<Q��<���<���<[��<i�<�U�<fx�<��<���<�_�<��<���<���<���<�l�<���<O(�<q6�<�)�<N�<�4�<�}�<m��<@��<�d�<��<��<\��<r��<��<���<�U�<S��<�#�<���<���<�9�<���<��<KJ�<O��<�<�E�<[<�<l��<�(�<��<C��<�c�<���<��<<3�<��<��<2��<�1�<G��<��<4�<m��<|�<�r�<r��<���<��<⳼<�˺<H˸<��<��<�Q�<E@�<��<���<�5�<���<��<te�<Z%�<�D�<��<vf�<L5�<"�<״�<o0�<Gi�<^�<��<���<�A�<_�<�d<d{<0�w<�-t<;�p<�l<�Ih<oc<(&^<d�X<%S<#�M<��H<�$D<#@<�7<<�^8<bF4<��/</�*<��$<��<��<86<!�
<�Q<5G�;4X�;/��;H��;�4�;�@�;k��;���;�s�;�$�;�ż;Zc�;�;�;��;C�;]X�;@A�;R�;�Ds;�g;�Z;&`M;��>;7�.;m�;N�;�E�:,��:�C�:D��:�:���:�ׄ:�&m:�J:$!:���9��h9;�6��W�n�й��go0��5B��iG��fA��2�H��z��,��~@��߹���^9�XH���6�VM�8G_�	�j�J�o��Sp�9�p��-t�K�}������,���|�����T�ú{^Ѻ�ۺ?��lk���뺧�}�����b��}.�V&��3���@���L�o�V�e�]��ka�hb���`���]�-�Y���U��+S��pR�<T���W�5�]���d�P�k��r��)w��tz�9F|�ZR}��~�Cf���`��ER���!������L��Z4�������  �  (w=�G=�9=�4=�=*�=�p=�� =y��<#��<��<���<s�<��<���<|��<&��<�f�<_4�<�
�<���<�#�<W$�<��<���<���<a��<��<~��<�l�<o�<B��<��<P:�<$&�<b��<���<���<�3�<��<Z��<̛�<��<���<���<M�<���<�`�<Au�<��<Ah�<}�<ф�<���<� �<��<�l�<�\�<���<rh�<�3�<���<�l�<~��<W)�<#K�<W��<Yf�<[��<��<���<қ�<;��<*��<��<���<�M�<�7�<ɪ�<���<��<���<ؽ�<�?�<�'�<�b�<qù<��<c%�<ҳ<�
�</ԭ<SG�<��<�Ţ<D,�<K�<�<�ז<��<9Г<!Β<��<c��<׏<�[�<�x�<1�<雇<�<;1�<!v<={<ܾw<��t< r<�o<e�k<HUg<�?b<	l\<�V<ѤO<�tI<��C<�'?<�=;<��7<*�4<pO1<_H-<Ci(<��"<�<�<O<��<���;km�;��;d��;Y��;8��;^)�;��;���;R��;c�;<M�;���;�"�;9�;�ɋ;Ǌ�;��u;�ii;8)_;�U;�\K;+?;Z0;��;xL;���:c%�:���:忆:le:�UK:�;:�-:�}:P�:0)�9z.9��v��	�� ��f�L�?�}�s���d���Ǘ� ���VT����d�,�E��;-��N�P����,�d�E��	f�h���_?������X���ZD�������ˋ�����㊺_���9ꢺ#����ͺ���n��ZZ����5U���@K�H��?�?��z?"��1�� A�,)Q���_��ek�	Es���v��v��r��l�68e��_�[���Y��X\��b�Qwj�It��C}�SI��lt�����wy���`��ˊ��h���8A���}��9������������O���  �  ��=�c=�U=�N=6=��=Z�=4� =%��<�
�<Y��<C�<�J�<;��<�#�<���<-�<��<)a�<�1�<���<�F�<�I�<��<m�<���<)��<���<���<��<��<��<���<�(�<��<ו�<ͻ�<��<�4�<1��<��<���<�K�<�%�</�<�6�<a�<6��</��<?�<��<&��<y��<���<u_�<�F�<��<��<6��<���<*^�<��<%��<ë�<�O�<Jv�<,/�<���<D��<	H�<���<���<���<I��<|�<���<�2�<<�<���<׸�<��<��<���<5n�<�\�<G��<���<�C�<�N�<���<�,�<-��<dm�<~��<s��<*f�<�'�<�]�<��<�Z�<��<���<;�<"�<��<耎<���<�_�<�χ<��<Pi�<D�<�{<��w<L�t<��q<b�n<|ek<� g<6b<4K\<`V<��O<��I<t3D<��?<�;<�R8<| 5<�1<�-<��(<��"<�J<�<(�<�Q<���;Ty�;�;���;���;���;L��;+S�;U]�;�e�;��;��;	�;���;'�;E��;(T�;��v;u*j;�n_;�sU;H�J;q>;)�/;~8;��
;c��:F3�:��:
��:��k:�eR:��A:��3:�":*�:�=�9	a@9�+�pv����
�*�E�ev��狺�-��;Г�o"��v~�!�_��)A���(����o ��'���?�oA_�	��N荺̪���{���'���֑��x��)x���;��;������fOͺ�P⺺�����������g\�V��bF������� !���/���?���O���]�!`i�('q���t�[.t�mp��j���c���]���Y���X��[��`�/�h��Rr��{��z���Ƀ�2����F���i���Ă����D����ڇ�|w���
���ꗻ=W��P����  �  !�=3�=d�=��=�u=�.=��=�	=j2 =g|�<<��<G��<���<���<M��<ϑ�<��</�<���<w��<�D�<{��<��<KR�<ԓ�<���<�l�<aY�<��<M��<%��<���<���<���<���<�G�<z�<gh�<\2�<� �<`��<�@�<��<��<0��<���<��<
��<��<ڠ�<���<o�<�?�<Ʉ�<r�<^�<8m�<dO�<��<&�<���<�}�<1��<��<���<b��<T��<9-�<�<
��<DW�<��<2��<���<R��<܌�<���<���<W�<�<��<���<o=�<��<��<�-�<q��<ĸ<��<�[�<���<�W�<"ت<�/�<���<��<ޜ<��<[֗<'
�<���<y��<Ŋ�<֊�<�^�<|�<��<�ފ<+^�<y��<��<�{�<�v|<��x<� u<��q<�n<��j<~�f<G}a<�[<��U<x�O<v/J<$E<�@<��<<}9<�76<�2<$v.<�y)<��#<t<:<�<��<]� <�l�;��;���;�2�;d�;5��;��;���;��;���;rط;e��;�M�;��;&�;cq�;<z;},l;E`;~�T;�0I;#5<;,<-;�?;�	;��:���:�n�:<�:f�}:Y�e:��T:=?E:�1:59:3B�9w�q9C�!7��n�)��E�1�j�_����WQ�����
���[�l�`P�j�3��|�y��(����`�.�Z�L��l�9Մ�%������A��N�������l捺�L����������X����̺��޺7��8���p}������@���`O��ן�������I�&g,���;�uK�A�X�0�c�!5k�)�n���n���k�*^f�HS`�'�Z�@�V�ƦU���W���\��yd���m���v�n�~���o��{ȃ�v���K~�����ⅻN���;>��:I��I����<��S����  �  �1==�=��=;�=�z=��=�L=�y =� �<D�<ҁ�<���<b��<���<5��<ǰ�<E�<?��<?�<f��<.�<�<�<���<F�<�U�<L=�<}$�<N1�<�}�<�<x��<���<���<�A�<���<o�<��<��<�.�<h�<���<f��<8��<��<{�<�*�<��<ǂ�<(�<X��<��<��<�s�<��<s�<��<�[�<��<���<|��<M�<gw�<���<!F�<���<�i�<���<K�<���<���<"~�<\)�<h��<>��<��<�R�<�A�<*��<�U�<��<��<���<y��<J��<I��<�F�<�r�<dY�<��<��<�ݮ<vp�<��<�_�<��<��<,8�<5�<�<؍�<�N�<5�<��<)�<-s�<嫍<ь�<
!�<Z��<{Ӄ<|9�<�}<&Py<'`u<ʥq<��m<F�i<ke<�{`<�$[<|�U<^P<�J<� F<� B<!g><�;<ϴ7<��3<e�/<ψ*<�$<$2<�J<�=<%T	<��<9��;`��;�!�;[=�;k��; ��;��;I�;�.�;2��;Td�;(z�;�|�;��;xO�;/M�;��~;��n;�`;jQS;o/F;J8;�$);`�;��;��:��:�t�:Jw�:PZ�:��:�n:\]:��F:z�':�`�9�9D0�8�t�<#������H>���\��(m��oo�9�e�2�R�06:��� �	u��w��z���ɩ���rj3��R��q�ު��t���됺Ej������������Q0��sP��n���%g̺ՎںZ��M�캌��J��!���� S���*������?�'��6��5D���P�'[��Rb��f�0�f��Od�)`��[��;V�>�R��dQ���R� qW�uz^�n)g��Rp���x��[������I�����؄�������%m����咻���Oٚ�y����  �  e�=y~=�q=�W=)!=��=<=&�=x� =e��<-#�<���<�.�<�<�U�<n��<?��<&�<Aq�<P��<�^�<c��<
��<���<���<B�<��<<��<g��<|��<5G�<���<�T�<���<��<=��<X�<]��<���<	F�<���<�}�<�a�<�a�<^�<y5�<>��<��<��<J��<�'�<K��</��<���<=Z�<�p�<&��<���<���<5��<K�<��<���<��<���<I'�<�<˺�<��<mV�<���<���<�@�<I��<�<:b�<Ņ�<�w�<�<�<(��<���<�B�<�"�<�4�<ar�<�ý<��<��<��<�c�<���<zd�<	�<��<�Z�<5*�<N5�<���<�@�<�J�<��<6�<��<鸒<Cp�<���<@�<�7�<p�<]V�<=��<E��<��~<��y<�lu<�q<��l<�oh<��c<k_<��Y<�T<��O<$_K<�*G<�hC<�?<��<<=09<�E5<r�0<g�+<��%<X<k�<��<s<}A<!&�;��;f�;@�;3��;�p�;j��;��;�W�;.�;��;�X�;���;�Q�;⢕;-�;LZ�;��p;�`;�P;E�A;ۋ2;�/#;k~;6�;F��:U��:;з:Α�:�:���:]m�:u�t:K[:ȇ9:��:[)�9*#$9�0X�@6��)��S��:2��|B�!G�q�A��4�f!�V��x���6۹�ӹW�߹ � �'��l8��$X�P
u��;���펺$B���\��臟�X饺�/��kE��Uú�-κ��׺E޺h��D*��W���交�躖�����i�	��R��L"� �/��F<���G�X�P��W��[�\�\�~�[�TY��VU��Q��N��RM��qN�09R�{}X��`�V�i�h�r�G�z������1��I1�����%ۈ�����΍��搻���)��ʳ�������  �  ��=��=u�=2�=k\=*�=he=�=v� =�9 =���<u��<�o�<�x�<���<�K�<w�<��<�:�<�}�<��<@�<�<��<<r�<L��<��<��<Vh�<!M�<�Q�<z�<���<�<��<���<o�<q��<H��<y-�<���<���<H��<�<���<��<�9�<�j�<�U�<|�<j��<\=�<���<˯�<��<���<�D�<��<���<��<���<�2�<[�<�]�<��<���<��<0Q�<g��<���< �<�<�'�<iC�<�^�< s�<jy�<�n�<mW�<e>�<c0�<�9�<fb�<P��<&�<`�<��<���<dI�<L��<PԲ<=ů<���<�o�<iT�<�Y�<N��<���<���<���<���<��<���<�3�<
ϑ<Q�<���<.��<�v�<��<�P�<��<K�<>z<�u<6 p<�Jk<��f<��a<d]<�cX<�S<�O<�K<�G<NyD<;A<��=<�G:<*6< v1<n*,<s^&<M; <a�<|�<�<��<�b<���;p��;��;�	�;��;���;�y�;���;}��;���;lp�;�2�;:	�;K�;�d�;"��;/<q;�'^;�/L;�*;;��*;1S;�j;���:���:���:�k�:��:�ơ:�@�:c��:t'�:�?i:�E:<4:�Q�95�d9ӳ8����z����ع�#��<����E��=��Ό
�������ܹ��ƹ@����Ĺ��߹wB��#���D�g.f�偂��珺0M��i���˭���������ź�ͺ�ӺEb׺��ٺ��ٺ ,ٺ"�غ�ۺ���V^�B�������@���z)��\4��>��F�oBL��lP��R�.S�% R�v3P�D�M���K�`�J�H�K�ΜN�hT���[���d�f;n�c�w�����ۃ���*���ڟ���&��ܡ��<���,������E������  �  *�=/�=S�=��=sm=��=g=!�=�=�o =��<���<D��<���<<!�<���<S6�<S��<���<5��<"��<��<��<���<M��<���<y
�<���<���<�Z�<��<k��<V��<�<�W�<_��<�O�<N�<s��<���<��<��<�G�<_�<�H�<���<lS�<|q�<�Z�<�%�<J��<ɾ�<ɫ�<���<T��<@2�<���<�.�<���<H��<���<{�<u�<
`�<I!�<C��<<��<B��<��<J1�<�&�<���<��<��<]o�<hL�<�5�<�.�<L:�<�\�<���<:��<m]�<���<�P�<_��<GҼ<m��<�R�<*��<ֲ<��<|�<�<�-�<�r�<�ա<�X�<���<�ǚ<���<�і<��<�r�<\�<.Z�<ܰ�<^Ԍ<���</P�<ë�<�؂<��<}z<�Ft<�n<LUi<C2d<+O_<ůZ<[ZV<SR<��N<�/K<'H<��D<��A<N�><%�:<"e6<ׅ1<�+,<~{&<� <Q�<�<��<�1
<�<�> <�S�;��;���;�l�;M��;nO�;�.�;���;���;%9�;c�;���;�;!~�;��;�o;�SZ;kF;�3;�!;��; �;��:l��: �:Y�:�:G��:{�:���:���:c�l:,UF:3:cK�9��9�M�8E|3�7B*�1_���F���ӹ5鹋[���P������I8չG�Ĺ�������(iӹ�	�����n�:��)`��􂺉ה�:���U��w���oɺ�AѺ�ֺmhں��ۺEۺ30ٺ�Rֺ��ӺY�Ӻ�ֺ#3޺ ?�sX��W��9��L��$��r-��'5���;�6JA���E�(I�<@K��gL���L�"L�+K���J��=K���M�O<R�`Y���a���k���v�����+~���򉻙ߍ�a>������N��% ���"�����Gܙ�ߠ���  �  ��=�=�=ܬ=LN=��=�;=y�==`� =B =9S�<T��<���<�Z�<2��<�+�<���<?�<��<r��<��<7��<���<�a�<��<s�<���<���<�<,��<~<�<p��<���<���<�b�<��<���<��<qA�<���<|��<K?�<[�<q5�<;��<�<C�<��<;��<���<� �<�:�<��<���<Vf�<Q��<�E�<��<�:�<&��<|�<W?�<_�< ��<YQ�<���<�w�<���<�!�<J��<���<Y6�<ɾ�<Q�<���<���<���<'��<MK�<���<e�<}�<���<dA�<s��<}��<pw�<���<\M�<��<���<���<�Y�<�ҧ<�^�<���<���<�.�<(қ<���<XT�<3H�<g�<+��<
�<Db�<`��<���<�E�<���<5ς<��<�By<��r<��l<�g<p�a<��\<� X<��S<5gP<Z7M<�PJ<f�G<��D<��A<�[><�e:<��5<��0<�y+<��%</t <X!<?<�<�?<g~<<�<��;���;k��;5+�;&:�;���;�5�;/��;��;��;V�;���;�֙;O�;~G�;�Zl;"�T;�S>;�);�;=;OI�:1��:=��:Pǿ:1�:�D�:�Ӧ:��:[ʒ:A+�:�d:]�;:�7:��9�Ń9ݲ9i��7��t�>��a�K��C���֢�n&��3ҹv�߹S�����,ٹ$Oѹ,Eѹ�L߹�l���Y��;��d��ׇ�}���Z1���xĺz�ӺJߺZ��F�꺌������%�ySݺ��׺=ԺԺ\jغ����p����	�	0�����!��*(��-��2�w�7�,7<�]�@��D��uH��K���L�(M�%PM�6�M�F�O��pS��Y���a�^l�Rx����u�������r���{��B����������F᜻1j���~��g���  �  B�=�= �=�p=1=�}=��=,Z=� =�x =C+ =���<�i�<M��<&^�<r��<��<?�<e�<H��<�g�<2�<Z�<��<���<�d�<���<��<�6�<��<���<U\�<���<���<X��<���<#��<1��<��<g��<��<���<���<f�<J��<D�<ds�<�t�<�h�<{o�<���<��<΍�<�/�<���<d�<���<C&�<M`�<*��<R��<-:�<���<@k�<A�<Ȱ�<��<��<�<��<���<��<{r�<o��<n�<+��<eV�<U�<6��<� �<���<~��<��<�N�<;�<�5�<�4�<��<�T�<$��<��<�?�<Ĭ<�q�<�<�<:�<\ߣ< ��<s)�<7��<��<p��<�=�<��<*�<�l�<w<`�<	�<}�<|[�<E|�<��~<x<qeq<��j<?�d<��^<P�Y< 6U<�qQ<BN<��K<�I<��F<gD<A<ݐ=<�k9<��4<5�/<�,*<��$<��<4�<Nw<�'<7�<Uw	<��<���;l��;5��;6��;���;�|�;�;�A�;���;as�;�o�;T6�;���;��;{��;5^g;��M;B�5;d�;}*;��:>�:�:2s�:S1�:D��:�M�:4��:��:-��:(�x:`�Q:"�':�g�9��9fe9��9�΋8��7��ϷsT���
���T�N������ݹn���� �/% �����j,��%' � ���4$�'�E��\p�a>��dA��Ol���׺���@���	X���U�������`�������^�ݺ]ٺ1�ٺ�]ߺ+꺑��K����£��	��� ���$�I�'��`+�6l/�;k4��@:��t@�mF�K�K��:O��iQ��dR�S��RT�TIW�I�\�r�d�8
o��m{��s��v@�������Y�����=�����!���l��޶�� '���  �  �=I�=|l=0=��=�=́=i� =6� =V =�. =� =r��<���<#�<�a�<4n�<a�<�Z�<y�<���<�r�<�I�<8�<��<Q��<��<�<H��<-�<bC�<�u�<r��<�[�<�H�<b��<�i�<��<{�<���<�h�<�<�j�<�}�<�3�<A��<���<��<���<X��<)-�<!��<5��<Z��<-t�<X$�<���<��<���<���<v��<��<\�<Ο�<�C�<���<�M�<�d�<t�<;?�<W�<�m�<��<���<���<�O�<��<���<�S�<���<���<���<���<���<[�<���<��<?!�<�~�</ų<��<ӟ�<�a�<]Z�<;s�<X��<W��<�X�<��<s>�<�u�<���<��<��<E{�<���<��<�F�<�r�<5U�<�ل<���<Ԗ}<B�v<m�o<.�h<�/b<0\<|�V< �R<O<�#L<F�I<՞G<�uE<	C<�@<�`<<�8<�$3<��-</�(<d#<f�<�j<t�<��<y	<"�
</n<�k<O�;-��;S��;0��;�Q�;9�;|�;�s�;���;���;$�;�Ɩ;��;��|;��a;��F;'[-;�;��;'��:�9�:7�:��:I��:���::�:37�:��:8�:��b:9:dv:YN�9]�9*M,9F<�8ͭ�8��8�f]8��7�"�~���m�Ԯ��g湺������.����ш����&� ��T5��V�ཀ�YY���̵�|�к8麦.������C	���	�d�8���������e��gr�W�⺛��z������j�����kt������!���"��
$��%��E)���.���5�t�=���E�mM�DS�yW���X�*�Y��Z���\��Ha���h�ps�$���(��o���ĕ����>!������DR���n���=���(��ɳ��3o���  �  AA=_J=�=��=B=�=3=Ѣ =;R =N+ =S$ =�+ =�, =T =���<���<&��<s~�<d7�<�<;�<մ�<�z�<�j�<�W�<��<��<2��<�+�<�|�<`��<���<h��<�T�<0�<1��<>Y�<���<�4�<���<���<D|�<3��<��<���<i��<��<��<}��<��<���<���<ή�<n��<��<g��<��<�:�<�<���<x�<AT�<:r�<9��<Hp�<��<���<6��<.y�<ճ�<�s�<���<=��<���<���<�9�<���<+��<�B�<��<��<�/�<�H�<�1�<0;<	�<�ܺ<�^�<���<�<�T�<���<w��<l,�<���<	ۦ<��<1�<sh�<���<���<ϡ�<o��<2�<>ˏ<=ڍ<'�<5��<�Ĉ<���<�P�<0y�<��|<��u<�;n<�g<�0`<�Z<^�T<BaP<��L<�VJ<27H<�PF<�QD<v�A<)�><4';< �6<!�1<#=,<w�&<��!<ێ<��<�a<�*<��<��<�<j<�w�;�w�;�z�;�*�;`�;]_�;Y��;XX�;���;�l�;Iޞ;u��;v�;�%x;��\;M�@;�2&;��;�`�:�h�:H~�:?ܩ:1�:���:gY�:N��:��:B�:��r:
RL:M :nB�9	��9�79ą�8o�8�h�8# �8"��8OG�8 ��7�{��*�K�����K�����)�d�1�p2��.��-���4�1BG���f��G��0ܣ������޺y����	�~�F����C������W����Lj�����A���� ��^	�3�����a�S="���"�K:"��!�4"��%�R�*��q2��<��\F���O���W�	�\��8_�T`���`��Bb�$f�hm��Cw��%��Ȩ��𓑻*@�� ��ir��������s���Ȩ�-��H?��Ǧ���  �  �=�=s�=�=��=�`=�� =�^ =� =+	 =D =�4 =SF =s8 =���<��<���<s��<a�<���<[��<�(�<���<D��<C��<n��<��<3%�<n��<a�<�%�<�%�<�A�<R��<%t�<��<1��<<��<O��<(��<ta�<9�<O��<>��<��<tU�<�N�<?7�<�A�<��<}Q�<�_�<O��<k��<��<)��<hi�<ex�<�3�<���<cF�<e��<I��<�C�<���<>~�<��<CD�<%�<2N�<��<�_�<�h�<S�<�L�<x��<�<��<N��<�d�<_�<ô�<���<�˿<�e�<L��<(^�<�з<O�<GT�<oï<���<ٟ�<D�<`��<�<�D�<*.�<���<�ٝ<��<g��<�{�<��<9H�<�F�<Ր�<W��<(E�<�K�<��<��<��{<��t<�:m<Q�e<��^<��X<:5S<��N<��K<D"I<�,G<]iE<��C<x%A<�><�@:<&�5<ax0<m
+<��%<�� <ٷ<�8<�2<+Q<�5<�<+<��<;�;���;7�;g�;�U�;�@�;i��;��;G��;���;�5�;T=�;Ӕ�;[u;�Y;��<;4g!;��;+��: ��:bN�:3��:Z�:��:[��:���:y!�:@؁:(bd:��;:�0:�c�9If9zO�8��~8��c8m��8���8�i9*��8�k�8��'��:������= ��"�@%9�5D��E�V3A�4�>���C�/�T��s�Lo�������Ⱥ���&]�����k�w���k�|��>�H���������W�y�z���*(�=�/��]��#���$��$�""��K �� �W�"��2(�|�0��m;�R�F���Q��Z�P�`���c���d��'e�?Of���i��Hp�IOz�����ef��]�����������2U��������A#���'��38��|���;���  �  ��==��=�l=��=(E=,� =�E =B =���<) =�6 =gN =1D =�	 =�5�<���<߈�<��<R��<��<���<��</��<(��<l�<���<� �<��<:��<���<<��<�<�g�<x1�<k��<�b�<g��<�q�<nU�<�:�<_��<�_�<a�<���<�$�<��<^��<��</j�<�-�<kK�<>��<&��<�-�<��<u��<6��<}=�<���<x3�<���<3��<k�<:��<~G�<���<��<{��<^)�<���<U8�<<�<��<��<?�<���<���<;L�<�+�<iM�<V��<���<���<�?�<Mm�<0�<��<Q۴<Q�<���<<W�<��<H�<���<T�<�Y�<�G�<�ʠ<W�<�ƚ<���<�d�<�<Y�<]�<�Y�<UÉ<e�<�"�<�ƃ<��<�q{<�St<U�l<Sqe<$d^<X<s�R<�dN<�$K<Y�H<��F<\E<�6C<�@<�=<��9<)F5<�0<W�*<xK%<H} <gf<z<�<�Z<�W<��<�`<�)<x�;f��;\��;��;(��;\w�;�ո;�9�;�֫;gۤ;ܚ�;��;T�;��s;�W;�H;;��;��; ��:,��:Y�:�$�:V��:\W�:�d�:Ac�:���:�:�_:�5:p�:ω�9b9K9��8c78�;82͡8ٗ�8/9��	9뮛8����#�5�0������O&���>���J�iL���G�Q�D�I5I�UY��w������qO˺�꺋%������i��^�P8����Y�\q ������Y�����q��G��N����� �Jv$�&�%���$�""�����q�]�!�s'��50�E>;�X:G�a�R���[��Xb��e�s�f���f���g��k�/sq��i{��H�����K��=g��'���Z[������������n����層٣���͢��  �  �=�=s�=�=��=�`=�� =�^ =� =+	 =D =�4 =SF =s8 =���<��<���<s��<a�<���<[��<�(�<���<D��<C��<n��<��<3%�<n��<a�<�%�<�%�<�A�<R��<%t�<��<1��<<��<O��<(��<ta�<9�<O��<>��<��<tU�<�N�<?7�<�A�<��<}Q�<�_�<O��<k��<��<)��<hi�<ex�<�3�<���<cF�<e��<I��<�C�<���<>~�<��<CD�<&�<2N�<��<�_�<�h�<S�<�L�<y��<�<��<P��<�d�<b�<ƴ�<���<�˿<�e�<P��<,^�<�з<S�<KT�<rï<���<۟�<F�<b��<�<�D�<*.�<���<�ٝ<��<e��<�{�<��<6H�<~F�<Ґ�<S��<$E�<�K�<��<��<��{<��t<�:m<N�e<��^<�X<:5S<��N<��K<G"I<�,G<aiE<āC<%A<�><�@:<.�5<hx0<t
+<��%<�� <߷<�8<�2</Q<�5<�<+<��<;�;���;/�;]�;�U�;�@�;[��;��;8��;u��;�5�;E=�;Ŕ�;Au;{Y;x�<;!g!;x�;��:��:ON�:$��:N�:��:T��:���:u!�:>؁:%bd:��;:�0:�c�9Ff9wO�8�~8��c8m��8���8�i9+��8�k�8��'��:������= ��"�@%9�5D��E�V3A�4�>���C�/�T��s�Lo�������Ⱥ���&]�����k�w���k�|��>�H���������W�y�z���*(�=�/��]��#���$��$�""��K �� �W�"��2(�|�0��m;�R�F���Q��Z�P�`���c���d��'e�?Of���i��Hp�IOz�����ef��]�����������2U��������A#���'��38��|���;���  �  AA=_J=�=��=B=�=3=Ѣ =;R =N+ =S$ =�+ =�, =T =���<���<&��<s~�<d7�<�<;�<մ�<�z�<�j�<�W�<��<��<2��<�+�<�|�<`��<���<h��<�T�<0�<1��<>Y�<���<�4�<���<���<D|�<3��<��<���<i��<��<��<}��<��<���<���<ή�<n��<��<g��<��<�:�<�<���<x�<AT�<:r�<9��<Hp�<��<���<6��<.y�<ֳ�<�s�<���<>��<���<���<�9�<���</��<�B�<��<��<0�<�H�<�1�<6;<�<�ܺ<�^�<���<�<�T�<���<|��<p,�<���<ۦ<��<1�<rh�<���<���<ˡ�<j��<,�<8ˏ<7ڍ<'�<.��<�Ĉ<���<�P�<)y�<��|<��u<�;n<�g<�0`<�Z<]�T<DaP<��L<�VJ<:7H<�PF<�QD<��A<6�><B';<�6</�1<0=,<��&<��!<�<��<�a<+<��<��<�<j<�w�;�w�;�z�;w*�;J�;D_�;>��;<X�;i��;�l�;,ޞ;Y��;[�;p%x;[�\;#�@;�2&;��;�`�:�h�:"~�:!ܩ:�:䙜:ZY�:D��:��:B�:��r:RL:M :jB�9��9�79���8n�8�h�8$ �8#��8PG�8%��7�{��*�K�����K�����)�d�1�p2��.��-���4�1BG���f��G��0ܣ������޺y����	�~�F����C������W����Lj�����A���� ��^	�3�����a�S="���"�K:"��!�4"��%�R�*��q2��<��\F���O���W�	�\��8_�T`���`��Bb�$f�hm��Cw��%��Ȩ��𓑻*@�� ��ir��������s���Ȩ�-��H?��Ǧ���  �  �=I�=|l=0=��=�=́=i� =6� =V =�. =� =r��<���<#�<�a�<4n�<a�<�Z�<y�<���<�r�<�I�<8�<��<Q��<��<�<H��<-�<bC�<�u�<r��<�[�<�H�<b��<�i�<��<{�<���<�h�<�<�j�<�}�<�3�<A��<���<��<���<X��<)-�<!��<5��<Z��<-t�<X$�<���<��<���<���<v��<��<\�<Ο�<�C�<���<�M�<�d�<u�<<?�<X�<�m�<��<���<���<�O�<��<���<�S�<��<���<���<���<��<#[�<���<(��<I!�<�~�<9ų<��<۟�<�a�<cZ�<?s�<[��<Y��<�X�<��<p>�<�u�<���<��<��<={�<���<��<�F�<�r�<+U�<�ل<���<Ė}<4�v<a�o<$�h<�/b<0\<{�V<"�R<!O<�#L<Q�I<�G<�uE<C<�@<�`<<�8<�$3<��-<A�(<d#<u�<�j<�<��<~	<%�
</n<�k<D�;��;<��;��;�Q�;�8�;V�;�s�;y��;���;��;rƖ;l�;x�|;[�a;u�F;�Z-;�;��;���:n9�:�:��:/��:u��:+�:)7�:��:8�:��b:9:av:UN�9[�9(M,9D<�8έ�8��8�f]8��7�"�~���m�Ӯ��g湺������.����Ј����&� ��T5��V�ཀ�YY���̵�|�к8麦.������C	���	�d�8���������e��gr�W�⺛��z������j�����kt������!���"��
$��%��E)���.���5�t�=���E�mM�DS�yW���X�*�Y��Z���\��Ha���h�ps�$���(��o���ĕ����>!������DR���n���=���(��ɳ��3o���  �  B�=�= �=�p=1=�}=��=,Z=� =�x =C+ =���<�i�<M��<&^�<r��<��<?�<e�<H��<�g�<2�<Z�<��<���<�d�<���<��<�6�<��<���<U\�<���<���<X��<���<#��<1��<��<g��<��<���<���<f�<J��<D�<ds�<�t�<�h�<{o�<���<��<΍�<�/�<���<d�<���<C&�<M`�<*��<R��<-:�<���<@k�<A�<Ȱ�<��<��<Ü�<��<���<��<}r�<r��<q�</��<jV�<U�<=��<� �<���<���<��<�N�<G�<�5�<5�<��<�T�<0��<��<�?�<Ĭ<�q�<�<�<>�<^ߣ< ��<q)�<4��<��<j��<�=�<��<
*�<�l�<k<T�<��<q�<q[�<:|�<�~<x<beq<��j<7�d<��^<O�Y<#6U<�qQ<BN<̄K<�I<äF<{D<"A<��=<�k9<ղ4<M�/<�,*<��$<��<D�<[w<�'<>�<Yw	<��<���;^��; ��;��;���;c|�;��;hA�;Ɛ�;/s�;�o�;!6�;Q��;R�;P��;�]g;[�M;�5;,�;N*;���:�=�:��:
s�:31�:,��:�M�:(��:��:'��:�x:Z�Q:�':�g�9��9de9�9�΋8	��7��ϷpT���
���T�M������ݹn���� �/% �����j,��$' � ���4$�'�E��\p�a>��dA��Ol���׺���@���	X���U�������`�������^�ݺ]ٺ1�ٺ�]ߺ+꺑��K����£��	��� ���$�I�'��`+�6l/�;k4��@:��t@�mF�K�K��:O��iQ��dR�S��RT�TIW�I�\�r�d�8
o��m{��s��v@�������Y�����=�����!���l��޶�� '���  �  ��=�=�=ܬ=LN=��=�;=y�==`� =B =9S�<T��<���<�Z�<2��<�+�<���<?�<��<r��<��<7��<���<�a�<��<s�<���<���<�<,��<~<�<p��<���<���<�b�<��<���<��<qA�<���<|��<K?�<[�<q5�<;��<�<C�<��<;��<���<� �<�:�<��<���<Vf�<Q��<�E�<��<�:�<&��<|�<W?�<_�< ��<YQ�<���<�w�<���<�!�<K��<���<[6�<̾�<�Q�<���<���<���<.��<VK�<���<e�<��<���<qA�<���<���<}w�<���<iM�<*��<���<���<�Y�<�ҧ<�^�<���<���<�.�<%қ<���<QT�<*H�<g�< ��<
�<7b�<S��<���<�E�<���<)ς<��<�By<��r<��l<�g<k�a<��\<� X<��S<@gP<h7M<�PJ<{�G<��D<��A<�[><�e:<��5<��0<�y+<��%<Dt <j!<N<�<�?<k~<<�<��;���;S��;+�;:�;���;�5�;���;��;��;�;���;�֙;�N�;NG�;�Zl;ѼT;�S>;�);l;;I�:���:��:-ǿ:�:�D�:�Ӧ:��:Tʒ:<+�:x�d:Y�;:�7:��9�Ń9۲9i��7��t�=��`�K��C���֢�m&��3ҹv�߹S�����,ٹ$Oѹ,Eѹ�L߹�l���Y��;��d��ׇ�}���Z1���xĺz�ӺJߺZ��F�꺌������%�ySݺ��׺=ԺԺ\jغ����p����	�	0�����!��*(��-��2�w�7�,7<�]�@��D��uH��K���L�(M�%PM�6�M�F�O��pS��Y���a�^l�Rx����u�������r���{��B����������F᜻1j���~��g���  �  *�=/�=S�=��=sm=��=g=!�=�=�o =��<���<D��<���<<!�<���<S6�<S��<���<5��<"��<��<��<���<M��<���<y
�<���<���<�Z�<��<k��<V��<�<�W�<_��<�O�<N�<s��<���<��<��<�G�<_�<�H�<���<lS�<|q�<�Z�<�%�<J��<ɾ�<ɫ�<���<T��<@2�<���<�.�<���<H��<���<{�<u�<`�<I!�<C��<=��<B��<��<K1�<�&�<���<��<��<`o�<mL�<�5�<�.�<T:�<�\�<Ș�<E��<y]�<���<�P�<m��<VҼ<{��<�R�<8��<ֲ<��<��<�<�-�<�r�<�ա<�X�<���<�ǚ<���<�і<��<{r�<Q�<!Z�<ΰ�<PԌ<���<!P�<���<�؂<��<iz<�Ft<s�n<CUi<>2d<*O_<ȯZ<cZV<"SR<ЛN<�/K<<H<��D<�A<i�><A�:<>e6<�1<,,<�{&<�� <d�<�<��<�1
<�<�> <�S�;ܾ�;���;nl�;&��;BO�;k.�;���;���;�8�;�b�;^��;�;�}�;P�;��o;`SZ;"F;�3;͝!;��;۩;ұ�:<��:���:=�:��:8��:q�:���:���:\�l:(UF:3:`K�9��9�M�8E|3�6B*�1_���F���ӹ5鹊[���P������I8չG�Ĺ�������'iӹ�	�����n�:��)`��􂺉ה�:���U��w���oɺ�AѺ�ֺmhں��ۺEۺ30ٺ�Rֺ��ӺY�Ӻ�ֺ#3޺ ?�sX��W��9��L��$��r-��'5���;�6JA���E�(I�<@K��gL���L�"L�+K���J��=K���M�O<R�`Y���a���k���v�����+~���򉻙ߍ�a>������N��% ���"�����Gܙ�ߠ���  �  ��=��=u�=2�=k\=*�=he=�=v� =�9 =���<u��<�o�<�x�<���<�K�<w�<��<�:�<�}�<��<@�<�<��<<r�<L��<��<��<Vh�<!M�<�Q�<z�<���<�<��<���<o�<q��<H��<y-�<���<���<H��<�<���<��<�9�<�j�<�U�<|�<j��<\=�<���<˯�<��<���<�D�<��<���<��<���<�2�<[�<�]�<��<���<��<1Q�<g��<���< �<�<�'�<lC�<�^�<s�<py�<�n�<uW�<m>�<l0�<�9�<rb�<\��<3�<`�<"��<���<rI�<Y��<\Բ<Hů<Û�<�o�<oT�<�Y�<Q��<���<���<���<���<��<���<�3�<�Α<�P�<���< ��<�v�<���<�P�<��<5�<�=z<�u<* p<xJk<��f<��a<g]<dX<�S<��O<��K<�G<dyD<;A<��=<H:<2*6<v1<�*,<�^&<b; <s�<��<��<��<�b<���;h��;��;}	�;��;[��;�y�;W��;J��;Ǖ�;4p�;u2�;	�;�J�;�d�;�;�;q;�'^;p/L;�*;;��*;S;�j;���:[��:���:sk�:��:xơ:�@�:[��:o'�:�?i:�E:94:�Q�92�d9γ8����z����ع�#��<����D��<��Ό
�������ܹ��ƹ@����Ĺ��߹wB��#���D�g.f�偂��珺0M��i���˭���������ź�ͺ�ӺEb׺��ٺ��ٺ ,ٺ"�غ�ۺ���V^�B�������@���z)��\4��>��F�oBL��lP��R�.S�% R�v3P�D�M���K�`�J�H�K�ΜN�hT���[���d�f;n�c�w�����ۃ���*���ڟ���&��ܡ��<���,������E������  �  e�=y~=�q=�W=)!=��=<=&�=x� =e��<-#�<���<�.�<�<�U�<n��<?��<&�<Aq�<P��<�^�<c��<
��<���<���<B�<��<<��<g��<|��<5G�<���<�T�<���<��<=��<X�<]��<���<	F�<���<�}�<�a�<�a�<^�<y5�<>��<��<��<J��<�'�<K��</��<���<=Z�<�p�<&��<���<���<5��<K�<��<���<��<���<I'�<�<˺�<��<nV�<���<���<�@�<L��<�<>b�<ʅ�<�w�<�<�</��<���<�B�<�"�<�4�<mr�<�ý<��<��<��<�c�<���<�d�<�<#��<�Z�<9*�<Q5�<���<�@�<�J�<��<�5�<��<ฒ<9p�<���<@�<�7�<d�<QV�<1��<:��<��~<��y<�lu<�q<��l<�oh<��c<n_<��Y<&�T<��O<4_K<�*G<iC<*�?<��<<V09<�E5<��0<}�+<ұ%</X<|�<��<�s<�A<(&�;��;xf�;2�;��;�p�;I��;ǥ�;pW�;�-�;f�;sX�;q��;xQ�;���;�,�; Z�;��p;\`;��P;�A;��2;\/#;J~;�;��:5��:#з:���:��:���:Wm�:l�t:E[:ć9:��:X)�9'#$9�0X�@6��)��S��:2��|B�!G�p�A��4�f!�V��w���6۹�ӹW�߹ � �'��l8��$X�P
u��;���펺$B���\��臟�X饺�/��kE��Uú�-κ��׺E޺h��D*��W���交�躖�����i�	��R��L"� �/��F<���G�X�P��W��[�\�\�~�[�TY��VU��Q��N��RM��qN�09R�{}X��`�V�i�h�r�G�z������1��I1�����%ۈ�����΍��搻���)��ʳ�������  �  �1==�=��=;�=�z=��=�L=�y =� �<D�<ҁ�<���<b��<���<5��<ǰ�<E�<?��<?�<f��<.�<�<�<���<F�<�U�<L=�<}$�<N1�<�}�<�<x��<���<���<�A�<���<o�<��<��<�.�<h�<���<f��<8��<��<{�<�*�<��<ǂ�<(�<X��<��<��<�s�<��<s�<��<�[�<��<���<|��<M�<gw�<���<!F�<���<�i�<���<K�<���<���<#~�<])�<j��<@��<��<�R�<�A�<0��<�U�<��<��<���<���<T��<S��<�F�<�r�<nY�<��<��<�ݮ<}p�<��<�_�<��<��<-8�<4�<	�<ԍ�<�N�<5�<��<!�<$s�<ܫ�<ǌ�< !�<P��<qӃ<s9�<�}<Py<`u<��q<��m<B�i<ke<�{`<�$[<��U<hP<�J<� F<B<3g><�;<�7<��3<x�/<�*<��$<42<�J<�=<.T	<��<?��;`��;�!�;O=�;Z��;	��;Ѵ�;�H�;n.�;��;,d�;�y�;�|�;��;QO�;	M�;T�~;C�n;��`;6QS;B/F;�I8;�$);E�;��;���:��:�t�:;w�:FZ�:��:�n:T]:��F:w�':�`�9�9?0�8�t�<#������H>���\��(m��oo�9�e�2�R�06:��� �	u��w��z���ɩ���rj3��R��q�ު��t���됺Ej������������Q0��sP��n���%g̺ՎںZ��M�캌��J��!���� S���*������?�'��6��5D���P�'[��Rb��f�0�f��Od�)`��[��;V�>�R��dQ���R� qW�uz^�n)g��Rp���x��[������I�����؄�������%m����咻���Oٚ�y����  �  !�=3�=d�=��=�u=�.=��=�	=j2 =g|�<<��<G��<���<���<M��<ϑ�<��</�<���<w��<�D�<{��<��<KR�<ԓ�<���<�l�<aY�<��<M��<%��<���<���<���<���<�G�<z�<gh�<\2�<� �<`��<�@�<��<��<0��<���<��<
��<��<ڠ�<���<o�<�?�<Ʉ�<r�<^�<8m�<dO�<��<&�<���<�}�<1��<��<���<b��<T��<9-�<�<
��<EW�< �<3��<���<T��<ތ�<���<���<W�<Ǘ�<��<���<u=�<��<��<�-�<y��<ĸ< ��<�[�<���<�W�<'ت<�/�<�<��<ޜ<��<Z֗<%
�<���<u��<���<ъ�<�^�<u�<��<�ފ<$^�<r��<}�<{{�<xv|<z�x<� u<}�q<�n<��j<~�f<H}a<�[<��U<�O</J</E<��@<��<<#}9<�76<��2<2v.<�y)<��#<<C<��<��<a� <�l�;��;���;�2�;X�;&��;��;���; ��;���;Vط;H��;eM�;�;
�;Hq�;�;z;O,l;`;Z�T;�0I;5<;<-;?;�	;���:���:�n�:<�:W�}:N�e:��T:8?E:�1:39:0B�9t�q9'�!7��n�)��E�1�j�_����WQ�����
���Z�l�`P�j�3��|�y��(����`�.�Z�L��l�9Մ�%������A��N�������l捺�L����������X����̺��޺7��8���p}������@���`O��ן�������I�&g,���;�uK�A�X�0�c�!5k�)�n���n���k�*^f�HS`�'�Z�@�V�ƦU���W���\��yd���m���v�n�~���o��{ȃ�v���K~�����ⅻN���;>��:I��I����<��S����  �  ��=�c=�U=�N=6=��=Z�=4� =%��<�
�<Y��<C�<�J�<;��<�#�<���<-�<��<)a�<�1�<���<�F�<�I�<��<m�<���<)��<���<���<��<��<��<���<�(�<��<ו�<ͻ�<��<�4�<1��<��<���<�K�<�%�</�<�6�<a�<6��</��<?�<��<&��<y��<���<u_�<�F�<��<��<6��<���<*^�<��<%��<ë�<�O�<Jv�<,/�<���<D��<	H�<���< ��<���<I��<}�<���<�2�<>�<���<ٸ�< ��<��<���<8n�<�\�<K��<���<�C�<�N�<���<�,�<0��<gm�<���<u��<+f�<�'�<�]�<��<�Z�<��<���<8�<"�<��<䀎<���<�_�<�χ<��<Li�<>�<�{<��w<H�t<��q<`�n<{ek<� g<6b<6K\<cV<��O<�I<y3D<��?<�;<�R8<� 5<��1<�-< �(<��"<�J<�<,�<�Q<���;Vy�;�;���;��;���;D��;!S�;I]�;�e�;��;��;�~�;���;�;7��;T�;��v;]*j;�n_;�sU;7�J;q>;�/;t8;��
;W��:=3�:��:��:z�k:�eR:��A:��3:�":(�:�=�9a@9�+�pv����
�*�E�ev��狺�-��;Г�o"��v~�!�_��)A���(����o ��'���?�oA_�	��N荺̪���{���'���֑��x��)x���;��;������fOͺ�P⺺�����������g\�V��bF������� !���/���?���O���]�!`i�('q���t�[.t�mp��j���c���]���Y���X��[��`�/�h��Rr��{��z���Ƀ�2����F���i���Ă����D����ڇ�|w���
���ꗻ=W��P����  �  z =q��<� =�M =� =_� =`K =�s�<���<���<�2�<=��<���<ZV�<�u�<hC�<��<��<���<��<.��<��<c��<r�<��<+��<�H�<���<��<��<�3�<���<P��<Ē�<��<s�<Z`�<$��<h��<7��<;�<��<��<���<�-�<`��<�G�<�M�<v��<ۆ�<���<N��<�h�<�K�<���<"W�<���<���<,��<���<���<���<�w�<֋�<���<K��<���<յ�<��<���<}b�<n��<��<,��<O\�<���<�,�<���<3�<��<��<N.�<��<{/�<��<���<�o�<QR�<�<��<�~�<�N�<ۖ�<���<Lj�<x�<�<���<⭓<�<���<�7�<���<�׎<���<��<,؉<g�<��<#��<]1{<��u<u�q<)�n<��l<k<'i<yef<�bb<�\<�HV<��N<�0G<�	@<#�9<Q�4<yI1<��.<'�,<�l*<�{'<e#<��<�L<Ӫ<��<q��;�;L+�;vI�;6�;�o�;��;��;R��;��;��;���;��;-�;�ލ;�Ԁ;' j;2V;c�G;˶=;��6;�1;=N*;�( ;'N;#�:#�:�ٙ:Q�R:[8�9I�}9�^�8S��7��7'8��Y8��7}f��z���U���lB��������@bú�պ�sݺK#ں��ͺ�������ې��6��nCx�b7�����,x��C^��9�Ӻ��3>�ƪ�\����ҺR�ú�縺f��~�Ӻ��ﺨ���Z�jE"��)�\q,�E�*�4m&��!�����!�Pn(��N4�^1D��jV���h���y�*����ㇻjy���x���e��Y����x� 
q�X�l�C�l���q��{�tp���j��䖑�y敻S͗�aP�����𯑻���d4���$��������������B�������l���  �  �0 = =5 =Gq =E� =�� =�` =x��<=��<|��<�h�<]#�<�&�<Χ�<���<��<���<���<���<^��<��<�:�<��<=7�<���<&@�<��<o<�<b�<# �<Zj�<��<&��<̍�<���<�a�<�U�<l��<6��<c�<�z�<�f�<���<���<z�<��<̀�<u}�<D��<'��<���<���<��<���<���<���<o�<45�<v��<$��<��<���<���<���<��<��<]�<g �<o��<��<��<?��<�4�<���<�`�<5��<��<.��<��<o��<J��<�`�<A)�<K|�<�k�<��<���<�<J#�<�4�<⤯<Zt�<`��<���<"��<-��<�<�<�J�<���<�X�<�8�<�o�<HǏ<� �<9�<�@�<�
�<�L�<�0�<2��<��{<o�v<=xr<Mgo<�%m<�?k<)'i<�Jf<c=b<��\<NCV<��N<�}G<|@<�g:<D�5<M�1<@N/<�,-<&�*<��'<^�#<KF<b�<�<G�< ��;ƺ�;Yu�;&��;Fc�;���;��;p��;Y7�;��;���;�B�;���;W�;Y	�;V�;�l;�Y;�J;�v?;(�7;��1;01*;߶;�;؋�:[y�:w�:��X:T3:�,�9�+9oz8H,^8kٗ8dԦ8��2869r��m��n<�@���V��s����кhFغ�7պ]ɺѶ�l衺�E����I9s��z�ʖ��qQ�������κ��ߺzl�@���޺jHѺDEú}�����q��GGԺ�ﺕ~�۶��  �qW'���)��<(�9$�8��+�G$ ��2'��3���B�I�T�og��w�nZ��o����1���G���X���0���kw���o��Wk��ak��kp���y��X���1���L��L�������@_��NP��2`�������g���l�����!�����������Ю��I���  �  �� =Q� =w� =\� =�� =�� =l� =| =0O�<�<�<��<=��<'��<-��<Ĵ�<�x�<]��<!��<�|�<�x�<C�<���<��<���<K��<(�<�y�<#�<�=�<���<X��<�o�<��<�x�<7��<g(�<u0�<{��<I$�<���<(�<8�<���<G��<FP�<���<E�<� �<lT�<�<�`�<�^�<I�<�U�<���<���<�<��<���<~�<Q�<�j�<Y�<� �<D��<;w�<���<���<���<~��<�}�<�n�<{��<2�<f�<�d�<a��<���<{��<��<
>�<Y��<L޾<�O�<aL�<�¸<}��<�>�<���<�<}�<�۬<X5�<�K�<�V�<���<�<�6�<'�<�2�<���<��<&L�<s�<zO�<p��<���< ��<n��<Yԁ<%�}<ax<^t<خp<  n<��k<,i<@�e<�a<�t\<�%V<�?O<�BH<,�A<��;<�A7</�3<R1<@�.<0,<��(<��$<�<+v<�<�-	<
c<��;B�;�Z�;Z�;V��;�;+K�;�7�;)��;�b�;�>�;'�;���;-M�;>��;��s;�`;4P;F(D;.�:;u�2;��);?:;�;�m�:���:&��:�Hh:I8:
7�9omy9H29��#9�@+9(�#9�?�8�Uq�� 8�%<ѹMQ+�lSo���a���_º�ɺ�?Ǻ����2���2������Vr�]e���j��›.����f��y���ѺR(ۺXsܺ��ֺ��̺��ºr���M����\ĺg�պ����\V��G��� ���"�b/!�V���W��]��F��#�ɿ/��?�&FP��a��q�Ϝ}��炻�����䃻�_���f{��Ys��Pl�#h���g��%l���t��L���Ɔ�U������0z��Yӓ�����꜐�7Ȏ�����T��_Ғ��O��v	��b
���Z���,���  �  F>=�,= A=�`=�l=~J=�� =�J =N��<���<���<���<m;�<���<J�<���<� �<9��<�W�<)�<4��<:8�<�%�<,��<��<h.�</��<Fk�<Br�<��<U��<0��<�<�B�<�.�<��<���<M��<`h�<q!�<"�<�Z�<r�<�)�<ȁ�<D��<��<y��<���<���<8�<q%�<�>�<ny�<��<���<f�<_�<���<�w�<nI�<��<]��<B��<�G�<K�<	��<w��<�<�1�<m��<�W�<VL�<�Z�<�V�<:�<�e�<0<�<���<���<P��<���<�ӿ<2w�<�<+��<ӟ�<�2�<Wz�< M�<㙰<j�<�ܩ<��<�Y�<���<�o�<���<�D�<�v�<�<, �<��<9�<b�<X�<�V�<���<�<M�<_�<.�z<2Dv<�cr<�o<�l<��h<O9e<��`<Ʊ[<��U<�O<X4I<EC<�><��9<#86<�m3<]�0<� .<zk*<F�%<6 <�<�u<�
<�<D%�;���;���;Vt�;���;���;@��;��;���;ͼ;0��;5�;j��;1��;Eъ;�v~;c�i;��X;n]J;�b>;Rr3;_+(;�E;x�;���:�]�:K�:�Q|:M�::��:^}�9�Ы9�7�9�'�9��9��I9��8ݸ�r��<P��vP�������#��{����z��B���{��t��vay��&`�Z�R���T��f�^��V����!��CX����Ⱥ kͺA�̺�Ⱥ�úG,��Bºa�ʺ��ٺ���x� �[�
�1Q����n�T��v��x����N�9��"+���9���I��PY�l�g�Ms�c�z��K~���}�,�y�Qt��om�psg��c�3�b��Jf���m���w��偻����i$������m��H{���ُ��E��:{������G��옻�l��L�����㬻�  �  !�=��=��=��=��=�=�3=l� =���<���<��<�4�<#��<~~�<���<�]�<l�<��<&L�<4��<�i�<���<���<�V�<��<�a�<)�<���< ��<���<<q�<�+�<'�<A��<̈�<8
�<	V�<�x�<���<˪�<���<-��<Sh�<ވ�<���< ��<���<"]�<!v�<�/�<"��<T��<)V�<���<��<���<S�<,��<��<2��<*'�<��<+�<`8�<���<U�<���<f4�<^]�<m��<���<�=�<=��<:}�<b�<S��<��<���<��<�{�<���<�0�<���<*��<�ݼ<�L�<�͹<T,�<�;�<�<Y�<��<��<��<d��<��<0��<�6�<�ޗ<��<�a�<Z�<ߑ<x��<rp�<q�<��<�ω<26�<�b�<���<x�}<}�x<�t</�o<+l<�-h<kd<s_<DmZ<SU< uO<��I<��D<q*@<�8<<��8<�6< 3<��/<M�+<�&<=!<��<< <�<�;`
�;3��;���;���;p��;*��;y5�;�u�;��;J��;�r�;VЦ;��;WW�;�݄;�Qt;j+a;�IP; *A;73;@�$;�U;��;G��:H��:秦:�&�:��X:	/:��:�v:���9���9���9R4�9�9^�%��S}�����N-���^�wɃ�IJ��ٱ��p���R��*���\�|�Nd���N���A�S�?�4�K��d��j��@������8d��|k���>ú�Dź.\ƺ�xȺI5ͺmmպẳ���u��-K�"E
�	�.}��E���
�`_
�j���"���լ&��4��*B�+�O�\\���f���m��q�)�q���o�C�k��g�L�b�vT_� m^�'�`��Of�d�n��Zy����bކ��������ꯎ������ؑ�ړ�Ǻ��]���k���q���糧�}���  �  �q=Mr=�u=jh=�8=��=OW=)� =7��<�W�<���<#j�<�'�<d�<c�<#��<���<���<T"�<�o�<w��<P��<��<���<;<�<cU�<�1�<���<���<��<���<q8�<ޣ�<��<O��<�<�}�<���<�f�<~��<t��<��<���<��<@��<���<�k�<~��<+��<�w�<^�<��<�W�<�<?�<^4�<���<q�<�r�<$��<$��<�)�<�c�<!t�<e<�<���<k��<�1�<�{�<	��<���<#��<�<yX�<b��<ѡ�<E��<'�<hH�<�<i��<{��<~��<���<��<c�<��<�޸<=��<�'�<VN�<�;�<J	�<Nͧ<ș�<M�<�<<�<A��<ws�<-��<*�<Ɉ�<�!�<���<9�<�<)w�<�<�{�<�<C�<�bz<?u<�Zp<M�k<��f<�3b<�f]<V�X<٪S<8�N<�,J<��E<R�A<�Y><�0;<�$8<��4<m1<>�,<,}'<�!<��<P<<:�<K�<�<h��;q�;�q�;���;ɪ�;�i�;X��;#�;eF�;f�;ˉ�;ک;3�;�;a��;G!};Dh;OT;��A;�a0;5�;�;���:ȕ�:��:�:O/�:
�n:f�N:�<8:�j(:�:$�
:���9���9��19!��gC�,i��!��<�4��pV�9fo� ~��"��s~��s�Ne��U�AyE�`�9��4��l:��JK��)f��ǃ�kS���~����x����ƺ�Pκ��պ�ݺ���$�����j�����l���53��1�����r����Ü����$���/�R�;�lG��DQ���Y��g`�\dd���e�J�e��<d���a�b_�d:]�G\��n]�_Ha�E�g�n�p�|�z��j������KÊ��덻F���6	��lk��ߗ�gc��t�������Zݡ����������  �  ~�=q�=�=9�=WL=�=C==�� =���<K��<�s�<.e�<�q�<��<���<.n�<V�<���<���<v��<���<���<��<���<Gr�<���<j��<���<cn�<-�<���<L��<m��<)�<R�<���<1T�<�<M��<��<���<��<�C�<i�<&c�<h�<o}�<���<��<OR�<y)�<s�<��<1�<�f�<Z��<�5�<9��<���<�d�<4J�<@�< ?�<V8�<�<F��<;��<��<F&�<N�<�H�<�,�<J�< ��<���<co�<�B�<(�<T#�<_1�<XR�<���<���<�;�<J��<q�<�-�<�<*��<l�<�<	�<=+�<�F�<�q�<í�<���<p�<�<GȘ<���<h��<�ݒ<I+�<w��<�
�<�m�<���<8��<��<�r�<휀<Sp{<Ҭu<� p<�qj<�e<w�_<ܽZ<
V<�Q<�M<��I<�F<��B<X�?<%�<<=W9<�5<�\1<�u,<�'<MX!<n�<��<�<5�
<�!<���;"��;�x�;���;��;��;n��;��;!��;�h�;-��;m�;���;9ؗ;iҌ;�[�;r�k;�TU;��?;+;�l;�9;���:���:�M�:a��:�S�:�*y:c4b:`6P:],@:��-:�:@r�9�,�90'9����o9�mr�����>��b*�{K>���L�~U��Y�0�Z��W���Q��I��a@���9�X9�Q�A���T�Iq�T�������]뭺���d�ͺ'�ۺl��	��tN���m��h� �k��ޖ�S� ��?���������������Ԭ�D�|����$���.�˽7��@� �G��cN�v�S�~RX�2s[�T�]���^��}_�gM_�[�^���]��1^�cH`���d���k�;�t�r=��߄��퉻����:�Ӗ��@����8M��+頻}
������������  �  ��=�=��=��=�=a�=�� =�? =�c�<Sv�<p��<+�<�q�<���<�?�<���<_��<�`�<0��<h�<�'�<�<�!�<�.�<s�<t��<G��<���<��<�&�<ʪ�<�9�<���< ��<5��<'1�<���<��<+�<b�<���<�+�<�y�<%��<�a�<��<���<���<���<̱�<��<x�<w�<���<m~�<��<<�<Y��<�`�<���<
M�<���<c��<�x�<�X�<��<��<.��<�C�<�y�<�Z�<@�<���<���<Eo�<%��<���<��<ζ�<��<��<�<ɺ�<<T�<5Ѿ<��<\�<h��<��<S-�<�M�<^��<�ު<�[�<i�<v��<Q*�<ӽ�<�J�<*ԙ<Bb�<��<�Ȓ<F��<��<XU�<5͋<�0�<)Y�<�-�<J��<bӀ<h�{<�Au<X�n<�h<��b<��\<k�W<ZS<�O<�K<cH<�E<v�B<��?<u�<<ch9<�A5<<v0<%+<�%<��<��<j}<��<��<�.<%n<�3�;�r�;Z��;���;��;���;�;e�;T��;�r�;ڟ�;���;�s�;�ٍ;�3�;��k;�S;Ғ:;�	#;;��:*d�:�F�:��:��:.5�:|�u:�hf:L�W:�rF:T�.:{�:KR�9��l9�-p8�;ǸI8h�+R��>�й���S2��$��4#�y1���?���L�W�@�\���\���W�3�O���I��J�
�U��l�HD�����ο���ź<�ںS�LF���9�C���
�Pf	��\�R}��K�����}1��D����:���B��K�]��Oo ��B)�}�0���6���;�I�@�0�D�W�I�qHN��.S�\X�?�\��X`�c�b���c���c�tpc�:�c�pbf�	�k�Kns���}�+����Ɋ�ߐ�7���Λ�I"���R��P@�����㥻/(������䢻�  �  g�=��=��=�1=��=d� =gI =@h�<��<$��<h��<8X�<��<���<�@�<u��<I��<)��<0��<���<�:�<g��<��<��<m6�<�<@��<,��<�T�<X��<�<�D�<���<_:�<)�<���<�Q�<���<5��<ט�<�D�<p��<`:�<{A�<��<��<���<���<��<2��<.�<p��<�{�<ke�<�C�<���<z�<���<��<F��<^��<U(�<C��<�M�<�,�<�<r��<��<���<�/�<��<�z�<���<v��<��<�X�<L��<E��<"�<[��<�{�<I]�< >�<���<��<証<�h�<�ʷ<��<��<�"�<W��<�0�<n�<��<��<��<~��<�=�<U��<]��<2��<�R�<��<��<�1�<Q��<mF�<W��<6��<Na�<G��<��z<�#t<�-m<<Cf<¢_<��Y<n2T<��O<�L<I<�F<@D<�A<�d?<�L<<zy8<��3<:�.<��(<�/#<��<��<�p<�e<(�<C�<�V<^�;�&�;�;�;��;�;&��;e��;ٸ;�D�;�`�;�]�;�q�;��;���;M�;�h;&N;6;3;/N;�f;A�:�1�:C��:E��:jh:Zp:�\f:qY]:��P:��<:+�:9,�9mB�9��87����e��i��?��	Ϲ�kչ��ܹ��빜������h0�_�J��Ob�t�k}��|���t�Kj�,�c��f�c�v�?���枺�r����Ѻ���<��+����j�A�L��?K���	���`� �;P��͌��3Q����� �~~)�r�0�E�5���8�\�:�<��!>��A���F���M��OU��5]�j:d���i�a}l�L0m��]l��nk���k�E6o��u����������>I���C��E���R���	�������Ы�����f���`q��n[���  �  �~=�{=�8=j�=<=�K =�2�<��<Qp�<�*�<�1�<�]�<�~�<�f�<���<�<���<��<�$�<?��<-�<"��<���<���<��<�,�<	��<2�<S��<��<�3�<T7�<`W�<~��<��<��< ��<Y�<���<���<��<N�<t��<���<��<��<���<2i�<�=�<�l�<��<I�<�<�<���<ü�<K��<#'�<�?�<�<��<AT�<B1�<�`�<:��<���<&��<���<\7�<�8�<n��<�m�</��<���<֮�<���<���<�A�<1�<|��<�V�<mZ�<�z�<���<l�<��<��<S~�<���<-��<���<�í<�T�<�G�<È�<��<�Z�<���<�n�<��<���<�ӗ<�<W��<��<���<�׊<�e�<��<��<A �<7΂<��<��y<�r<%>k<��c<��\<�]V<�P<_�L<N I<ȋF<�D<t�B<��@<K><P;<��6<��1<�6,<9&<zi <�*<Э<��<�<��<�]	<ʢ<h$<���;ɠ�;2��;U�;Q��;tB�;k��;N��;�]�;��;��;�p�;��;��~;�Nd;��G;b+;P9;���:@��:���:�M�:��k:�4[:�T:Q:�L:?�@:�):�:���9�9����߁�����2�J�p޹1�˹����p�����۹�}��K*���P�x�u�G����������,��2��g�������Ϟ�����䕧�I:º'�ߺ������������K�"�wK"�[;���������	�%��$��'��O���X��+�24��>:�� =��=�*�;���9��9��<�u�A�;J���T�Q�_��j���q�I�v�1.x�w��t���s�qCu��z��聻�X�������(��� ���:��ݬ����F����������8���,}�������  �  h6=�+=��=�@=q} =�Z�<���<���<#a�<�]�<ŷ�<;�<m��<��<}a�<�m�<�<wO�<n��<��<U��<�c�<O�<&��<e�<PH�<�&�<�{�<!>�<���< t�<�I�<i:�<�y�<�3�<0��<�t�<z��<v��<f��<���<��<2 �<2��<,A�<�<���<�%�<���<^>�<@�<xO�<���<���<5��<x�<[��<��<G	�<V�<&��<;�<$4�<��<���<
��<���<�\�<p��<��<���<��<���<x��<�i�<{k�<N��<��<�A�<f*�<]�<(��<��<&Ҿ<AI�<�3�<���<|��<Y_�<�B�<�{�<Q.�<]�<W�<���<�k�<��<bܠ<�F�<�,�<н�<�8�<gސ<��<5u�<b��<+�< �<�ǅ<=�<|.�<�<A�x<\Iq<�i<E�a<�NZ<V�S<N!N<9�I<Z�F<�[D<��B<�2A<|?<�=<��9<f5<�0<��)<�#<q�<R�<0�<zO<��<�V<�	<�k<U<:�;�0�;:?�;>G�;�D�;���;��;+��;5��;�;ґ�;���;���;kz;l�_;!-B;��#;�;���:��:� �:cZa:��F:l�;:qf::�}<:��::�/:>:���9�"^9�W�?�o���ҹC[����,�(L��͹Rխ�򀦹�����T����)��B[�eW��K���k����Q��w��Iݛ�B璺����qp���
��B���C�̺��캦��:	�[T"���*��-�m�,�(J'���\�����\	�����
��J��$���)��G5�?>��?C�O*D���A��=�:W9��7�Y�8�B�>���H���U��hc��.p��7z��4���8��������}��f{�tz{�t��J-��	���Gɒ�����gW��"���2������q��莶��곻|=���W������  �  	=��= �=�� =� =�|�<X�<9�<ě�<	��<�T�<�<q��<���<g��<���<h�<V�<\'�<5p�<�.�<��<6i�<}��<�C�<ä�<x��<��<	��<��<T��<���<�z�<���<tJ�<f��<���<"�<��<MK�<�q�<$P�<��<O|�<ê�<�\�<���<qC�<��<f�<4S�<K��<Ӑ�<�o�<��<AC�<|��<?��<���<�</%�<k��<�\�<Ͼ�<.��<���<���<��<-�<��<�d�<���<�_�<���<��<��<���<���<U_�<�`�<��<*�<m�<b�<lҼ<���<�<+ϴ< ��<�X�<��<�Z�<���<�s�<ps�<�g�<��<��<�y�<A�</��<�ޓ<RL�<+(�<���<���<WN�<Q8�<��<]��<5��<c9~<��w<�Sp<�Uh<�I`<��X<��Q<EL<��G<��D<��B<}sA<W/@<�><�A<<��8<3E4<�.<*c(<)�!<�<��<�<o<��<�<��	<��<G�<l��;[T�;���;��;���;��;�w�;�z�;�W�;f��;��;Ȣ�;��;\@w;�D\;�3>;��;� ;�T�:�^�:rIs:h�E:#�-:I6&:��(:�.:��-:��!:4�:��9 9j�����E��<!���'�"3�Gi��ѹ�Ǧ�k���A˲�bS��ޭ+��?d�>���̣��ﱺꤶ�s���E��Ha�������d�����Y��}�Ӻ'���b?��T��V)���1�F/5�1f3�gc-��$�+��a�Ԭ��O�5��L�#��I0�=q<��XE�@�I���I�f{E�-b?�i9�6�5���6�c�<��H�ؚV��Kf��t��!��ۧ���ӄ�p���#��fj����������څ��b��d��������.���d��ȵ��������`⹻�϶�󥲻P��C̪��  �  ��=8�=fw=� =���<o-�<���<���<�S�<���<.�<��<��<H�<B��<B��<�<.�<Y��<3�<A��<e0�<��<�r�<���<�i�<Sn�<8��<���<���<��<.p�<�6�<S�<g��<iF�<C�<���<���<�<EG�<�)�<v��<�N�<ht�<�<V��<u��<��<��<`�<Ԓ�<�q�<=f�<��<�S�<]��<���<-��<E��<���<�B�<��<�k�<K�<�y�<��<Ն�<u��<|f�<�<�<n�<�,�<x��<�P�<�3�<���<���<��<��<(v�<��<fB�<�9�<M��<�w�<b��<9��<{4�<.�<�@�<��<�n�<�E�<[�<�c�<��<]'�<)��<�E�<���<g��<��<t�<�L�<_�<\��<���<_߄<�{�<��<��}<�vw<��o<��g<��_<�X<>Q<d�K<�UG<�VD<�]B<�A<��?<�H><��;<-�8<��3<N-.<]�'< Y!<{\<BS<r<�<ƣ<Q�<m�	<��<İ<+�;wV�;:�;���;�ۿ;pĳ;f:�;A9�;0(�;��;L4�;2�;�B�;6v;}[;�<;�C;�.�:���:QT�:i:��;:��$:G�:u�":��(:E):�:ko :?��9�T�8#;��Ĺ�T�-�*��;0�k�"��D��<Թ\ �������)#�W�,���g�Ø��狀Nȶ��̻��������O~��$���J���n��Z����ֺ����"�܌�C�+�ts4�7�7�C�5���/�}x&��|�V��~��٘��u�m��7%���2��?���G�L��wK�e�F��@���9���5�,<6�;}<�,�G��
W�ng���v��<��o焻����E��	F��.d���΀�X^���v������f��"͞��0���������
���Q��h���շ��|������i���  �  	=��= �=�� =� =�|�<X�<9�<ě�<	��<�T�<�<q��<���<g��<���<h�<V�<\'�<5p�<�.�<��<6i�<}��<�C�<ä�<x��<��<	��<��<T��<���<�z�<���<tJ�<f��<���<"�<��<MK�<�q�<$P�<��<O|�<ê�<�\�<���<qC�<��<f�<4S�<K��<Ӑ�<�o�<��<AC�<|��<?��<���<�</%�<k��<�\�<Ͼ�<.��<���<���<��<-�<��<�d�<���<�_�<���<��<��<���<���<W_�<�`�<��<.�<m�<b�<pҼ<���<�<0ϴ<%��<�X�<��<�Z�<���<�s�<rs�<�g�<��<��<�y�<A�<-��<�ޓ<OL�<'(�<���<���<RN�<L8�<��<X��<0��<Z9~<��w<�Sp<�Uh<�I`<��X<��Q<EL<��G<��D<��B<�sA<]/@<�><�A<<��8<<E4<��.<3c(<2�!<<�<�<v<��<�<��	<��<G�<i��;UT�;}��;���;~��;��;�w�;|z�;�W�;S��;��;���;��;8@w;yD\;�3>;��;�� ;�T�:�^�:7Is:9�E:��-:,6&:x�(:�.:��-:��!:.�:��9�9w�� ���F��<!���'�"3�Gi��ѹ�Ǧ�j���@˲�bS��ޭ+��?d�>���̣��ﱺꤶ�s���E��Ha�������d�����Y��}�Ӻ'���b?��T��V)���1�F/5�1f3�gc-��$�+��a�Ԭ��O�5��L�#��I0�=q<��XE�@�I���I�f{E�-b?�i9�6�5���6�c�<��H�ؚV��Kf��t��!��ۧ���ӄ�p���#��fj����������څ��b��d��������.���d��ȵ��������`⹻�϶�󥲻P��C̪��  �  h6=�+=��=�@=q} =�Z�<���<���<#a�<�]�<ŷ�<;�<m��<��<}a�<�m�<�<wO�<n��<��<U��<�c�<O�<&��<e�<PH�<�&�<�{�<!>�<���< t�<�I�<i:�<�y�<�3�<0��<�t�<z��<v��<f��<���<��<2 �<2��<,A�<�<���<�%�<���<^>�<@�<xO�<���<���<5��<x�<[��<��<G	�<V�<&��<;�<$4�<��<���<
��<���<�\�<p��<��<���<��<���<z��<�i�<~k�<R��<��<�A�<l*�<]�<0��<��</Ҿ<II�<�3�<���<���<b_�<�B�<�{�<X.�<
]�<\�<���<�k�<��<cܠ<�F�<�,�<̽�<�8�<aސ<��<-u�<Z��<�*�< �<�ǅ<=�<t.�<�<2�x<OIq<�i<=�a<�NZ<R�S<M!N<<�I<_�F<�[D<��B<�2A<+|?<�=<��9<f5<�0<��)<.�#<��<b�<?�<�O<�<�V<	�	<�k<U<4�;�0�;*?�;)G�;�D�;���;��;��;��;��;���;���;���;�jz;*�_;�,B;��#;�;O��:ڮ�:� �:Za:c�F:4�;:Hf::�}<:��::�/:
>:���9�"^9[W�F�o���ҹD[����,�(L��͹Rխ�񀦹�����T����)��B[�eW��K���k����Q��w��Iݛ�B璺����qp���
��B���C�̺��캦��:	�[T"���*��-�m�,�(J'���\�����\	�����
��J��$���)��G5�?>��?C�O*D���A��=�:W9��7�Y�8�B�>���H���U��hc��.p��7z��4���8��������}��f{�tz{�t��J-��	���Gɒ�����gW��"���2������q��莶��곻|=���W������  �  �~=�{=�8=j�=<=�K =�2�<��<Qp�<�*�<�1�<�]�<�~�<�f�<���<�<���<��<�$�<?��<-�<"��<���<���<��<�,�<	��<2�<S��<��<�3�<T7�<`W�<~��<��<��< ��<Y�<���<���<��<N�<t��<���<��<��<���<2i�<�=�<�l�<��<I�<�<�<���<ü�<K��<#'�<�?�<�<��<AT�<B1�<�`�<:��<���<'��<���<]7�<�8�<o��<�m�<0��<���<خ�<���<���<�A�<1�<���<�V�<vZ�<�z�<���<l�<��<��<`~�<���<:��<Ð�<�í<�T�<�G�<ˈ�<��<�Z�<���<�n�<��<���<�ӗ<ꤔ<O��<��<���<�׊<�e�<��<���<4 �<+΂<��<��y<�r<>k<��c<��\<�]V<�P<b�L<U I<ӋF<�D<��B<Ϸ@<%K><g;<��6<��1<�6,</9&<�i <�*<�<��<�<��<�]	<΢<h$<���;���;��;�T�;.��;KB�;=��;��;�]�;��;��;�p�;n�;&�~;@Nd;|�G;+;9;5��:���:1��:�M�:D�k:74[:mT:�Q:ҍL:)�@:�):�:{��9�9����߁�����2�J�p޹0�˹����p�����۹�}��K*���P�x�u�G����������,��2��g�������Ϟ�����䕧�I:º'�ߺ������������K�"�wK"�[;���������	�%��$��'��O���X��+�24��>:�� =��=�*�;���9��9��<�u�A�;J���T�Q�_��j���q�I�v�1.x�w��t���s�qCu��z��聻�X�������(��� ���:��ݬ����F����������8���,}�������  �  g�=��=��=�1=��=d� =gI =@h�<��<$��<h��<8X�<��<���<�@�<u��<I��<)��<0��<���<�:�<g��<��<��<m6�<�<@��<,��<�T�<X��<�<�D�<���<_:�<)�<���<�Q�<���<5��<ט�<�D�<p��<`:�<{A�<��<��<���<���<��<2��<.�<p��<�{�<ke�<�C�<���<z�<���<��<F��<^��<V(�<C��<�M�<�,�<�<r��<��<���<�/�<��<�z�<���<y��<��<�X�<R��<L��<#"�<e��<�{�<U]�<>�<���<��<���<�h�<�ʷ<��<*��<�"�<d��<�0�<x�<��<��<��<��<�=�<Q��<W��<)��<�R�<��<��<�1�<A��<]F�<G��<&��<?a�<8��<��z<#t<�-m<.Cf<��_<��Y<m2T<��O<�L<&I<��F<@D<'�A<�d?<�L<<�y8<��3<Z�.<
�(<0#<�<��<�p<�e<5�<L�<�V<^�;�&�;q;�;��;��;���;2��;�ظ;oD�;|`�;~]�;Yq�;G�;���;�L�;��h;�%N;�:3;�M;Ff;��:�1�:�:��:	h:�Yp:�\f:JY]:��P:o�<:�:(,�9bB�9��8D����e��i��?��	Ϲ�kչ��ܹ��빜������h0�^�J��Ob�t�k}��|���t�Kj�+�c��f�c�v�?���枺�r����Ѻ���<��+����j�A�L��?K���	���`� �;P��͌��3Q����� �~~)�r�0�E�5���8�\�:�<��!>��A���F���M��OU��5]�j:d���i�a}l�L0m��]l��nk���k�E6o��u����������>I���C��E���R���	�������Ы�����f���`q��n[���  �  ��=�=��=��=�=a�=�� =�? =�c�<Sv�<p��<+�<�q�<���<�?�<���<_��<�`�<0��<h�<�'�<�<�!�<�.�<s�<t��<G��<���<��<�&�<ʪ�<�9�<���< ��<5��<'1�<���<��<+�<b�<���<�+�<�y�<%��<�a�<��<���<���<���<̱�<��<x�<w�<���<m~�<��<<�<Y��<�`�<���<
M�<���<c��<�x�<�X�<��<��</��<�C�<�y�<�Z�<A�<���<���<Jo�<*��<���<��<ض�<��<��<�<غ�<MT�<FѾ<��<o�<z��<��<d-�<N�<m��<�ު<�[�<r�<|��<T*�<ӽ�<�J�<%ԙ<;b�<��<�Ȓ<9��<��<HU�<$͋<�0�<Y�<�-�<9��<RӀ<L�{<�Au<C�n<�h<��b<��\<i�W<^S<�O<�K<cH<�E<��B<��?<��<<�h9<B5<`v0<A%+<	�%<��<ܗ<�}<�<�<�.<*n<�3�;�r�;E��;���;ݧ�;}��;G�;&�;��;hr�;���;M��;�s�;Tٍ;m3�;v�k;2S;j�:;_	#;�;���:�c�:0F�:��:٤�:5�:?�u:ahf:-�W:�rF:F�.:q�:?R�9��l9�-p8�;ǸJ8h�*R��=�й���R2��$��4#�y1���?���L�W�@�\���\���W�3�O���I��J�
�U�l�HD�����ο���ź<�ںS�LF���9�C���
�Pf	��\�R}��K�����}1��D����:���B��K�]��Oo ��B)�}�0���6���;�I�@�0�D�W�I�qHN��.S�\X�?�\��X`�c�b���c���c�tpc�:�c�pbf�	�k�Kns���}�+����Ɋ�ߐ�7���Λ�I"���R��P@�����㥻/(������䢻�  �  ~�=q�=�=9�=WL=�=C==�� =���<K��<�s�<.e�<�q�<��<���<.n�<V�<���<���<v��<���<���<��<���<Gr�<���<j��<���<cn�<-�<���<L��<m��<)�<R�<���<1T�<�<M��<��<���<��<�C�<i�<&c�<h�<o}�<���<��<OR�<y)�<s�<��<1�<�f�<Z��<�5�<9��<���<�d�<4J�<@�< ?�<V8�<�<F��<;��<��<F&�<N�<�H�<�,�<L�<$��<���<ho�<�B�<(�<^#�<k1�<eR�<Ȉ�<���<�;�<\��<��<�-�<'�<<��<}�</�<�<J+�<�F�<�q�<ʭ�<���<p�<�<CȘ<���<_��<�ݒ<;+�<h��<�
�<�m�<睊<&��<��<�r�<ݜ�<5p{<��u<� p<�qj<�e<p�_<۽Z<
V<�Q<+�M<ШI<�F<��B<w�?<G�<<`W9<�5<�\1<v,<�'<lX!<��<��<�<E�
<�!<	��;"��;�x�;޷�;��;���;<��;���;᱿;�h�;㠲;"�;���;�ח; Ҍ;�[�;��k;]TU;P�?;�+;zl;_9;<��:$��:�M�:)��:�S�:�*y:54b:?6P:F,@:��-:�:3r�9�,�9('9���o9�mr�����=��b*�zK>���L�~U��Y�0�Z��W���Q��I��a@���9�X9�Q�A���T�Iq�T�������]뭺���d�ͺ'�ۺl��	��tN���m��h� �k��ޖ�S� ��?���������������Ԭ�D�|����$���.�˽7��@� �G��cN�v�S�~RX�2s[�T�]���^��}_�gM_�[�^���]��1^�cH`���d���k�;�t�r=��߄��퉻����:�Ӗ��@����8M��+頻}
������������  �  �q=Mr=�u=jh=�8=��=OW=)� =7��<�W�<���<#j�<�'�<d�<c�<#��<���<���<T"�<�o�<w��<P��<��<���<;<�<cU�<�1�<���<���<��<���<q8�<ޣ�<��<O��<�<�}�<���<�f�<~��<t��<��<���<��<@��<���<�k�<~��<+��<�w�<^�<��<�W�<�<?�<^4�<���<q�<�r�<$��<$��<�)�<�c�<!t�<e<�<���<k��<�1�<�{�<
��<���<%��<�<}X�<g��<ס�<L��</�<rH�<�<v��<���<���<ħ�<��<c�<-��<�޸<O��<�'�<fN�<�;�<W	�<Xͧ<Й�<S�<Ő�<=�<?��<ss�<&��< �<���<�!�<|��<9�<�~�<w�<m�<�{�<Ⲃ<$�<ebz<�>u<�Zp<=�k<��f<�3b<�f]<Z�X<�S<F�N<�,J<�E<m�A<�Y><�0;<�$8<��4<�1<`�,<M}'<��!<��<h<<N�<[�<��<s��;q�;�q�;���;���;�i�;(��;��;'F�;#�;���;�٩;��;� �;��;� };�h;�NT;��A;pa0;�;�;���:n��:���:��:&/�:��n:9�N:�<8:�j(:�:�
:x��9���9��19��gC�,i�� ��;�4��pV�9fo� ~��"��r~��s�Ne��U�AyE�`�9��4��l:��JK��)f��ǃ�kS���~����x����ƺ�Pκ��պ�ݺ���$�����j�����l���53��1�����r����Ü����$���/�R�;�lG��DQ���Y��g`�\dd���e�J�e��<d���a�b_�d:]�G\��n]�_Ha�E�g�n�p�|�z��j������KÊ��덻F���6	��lk��ߗ�gc��t�������Zݡ����������  �  !�=��=��=��=��=�=�3=l� =���<���<��<�4�<#��<~~�<���<�]�<l�<��<&L�<4��<�i�<���<���<�V�<��<�a�<)�<���< ��<���<<q�<�+�<'�<A��<̈�<8
�<	V�<�x�<���<˪�<���<-��<Sh�<ވ�<���< ��<���<"]�<!v�<�/�<"��<T��<)V�<���<��<���<S�<,��<��<2��<*'�<��<+�<`8�<���<U�<���<g4�<_]�<n��<���<�=�<?��<=}�<f�<W��<!��<���<��<|�< ��<�0�<���<8��<�ݼ<M�<ι<e,�<�;�<#�<h�<��< ��<��<k��<��<3��<�6�<�ޗ<��<�a�<R�<�ޑ<l��<dp�<c�<��<�ω<"6�<�b�<q��<\�}<d�x<�t<�o<l<�-h<fd<s_<HmZ<[U<,uO<��I<��D<�*@<9<<��8<�6<< 3<�/<l�+<$�&<=!<��<1<<�</�;j
�;3��;���;���;T��;��;M5�;zu�;��;��;�r�;Ц;j�;W�;I݄;7Qt;�*a;FIP;�)A;�3;��$;�U;f�;���:	��:���:z&�:W�X:�/:��:�v:���9���9���9K4�9�9l�%��S}�����N-���^�wɃ�HJ��ٱ��p���
R��*���\�|�Nd���N���A�S�?�3�K��d��j��@������8d��|k���>ú�Dź.\ƺ�xȺI5ͺmmպẳ���u��-K�"E
�	�.}��E���
�`_
�j���"���լ&��4��*B�+�O�\\���f���m��q�)�q���o�C�k��g�L�b�vT_� m^�'�`��Of�d�n��Zy����bކ��������ꯎ������ؑ�ړ�Ǻ��]���k���q���糧�}���  �  F>=�,= A=�`=�l=~J=�� =�J =N��<���<���<���<m;�<���<J�<���<� �<9��<�W�<)�<4��<:8�<�%�<,��<��<h.�</��<Fk�<Br�<��<U��<0��<�<�B�<�.�<��<���<M��<`h�<q!�<"�<�Z�<r�<�)�<ȁ�<D��<��<y��<���<���<8�<q%�<�>�<ny�<��<���<f�<_�<���<�w�<nI�<��<]��<B��<�G�<K�<
��<w��<�<�1�<n��<�W�<XL�<�Z�<�V�<>�<�e�<6<�<���<���<Y��<���<�ӿ<>w�< ��<8��<៸<�2�<dz�<M�<<j�<�ܩ<��<�Y�<���<�o�<���<�D�<�v�<	�<% �<�</�<W�<X�<�V�<���<�<A�<R�<�z<Dv<�cr<�o<�l<��h<K9e<��`<ɱ[<��U< �O<f4I<-EC<�><��9<;86<�m3<w�0<� .<�k*<^�%<"6 <��<
v<�
<�<S%�;���;���;Nt�;���;���;#��;��;k��;�̼;��;�4�;4��;���;ъ;�v~; �i;a�X;]J;eb>;r3;%+(;�E;O�;G��:�]�:#�:�Q|: �::��:/}�9�Ы9�7�9s'�9��9��I9	��8�ݸ�r��<P��vP�������#��z����z��B���{��t��vay��&`�Y�R���T��f�^��V����!��CX����Ⱥ kͺA�̺�Ⱥ�úG,��Bºa�ʺ��ٺ���x� �[�
�1Q����n�T��v��x����N�9��"+���9���I��PY�l�g�Ms�c�z��K~���}�,�y�Qt��om�psg��c�3�b��Jf���m���w��偻����i$������m��H{���ُ��E��:{������G��옻�l��L�����㬻�  �  �� =Q� =w� =\� =�� =�� =l� =| =0O�<�<�<��<=��<'��<-��<Ĵ�<�x�<]��<!��<�|�<�x�<C�<���<��<���<K��<(�<�y�<#�<�=�<���<X��<�o�<��<�x�<7��<g(�<u0�<{��<I$�<���<(�<8�<���<G��<FP�<���<E�<� �<lT�<�<�`�<�^�<I�<�U�<���<���<�<��<���<~�<Q�<�j�<Y�<� �<E��<;w�<���<���<���<��<�}�<�n�<}��<3�<f�<�d�<d��<���<���<	��<>�<`��<T޾<�O�<jL�<�¸<���<�>�<���<���<��<ܬ<^5�<�K�<�V�<���<�<�6�<&�<�2�<���<��< L�< s�<sO�<h��<���<��<d��<Pԁ<�}<ax<Pt<ˮp<��m<�k<&i<=�e<�a<�t\<&V<�?O<�BH<8�A<��;<�A7<@�3<d1<R�.<'0,<��(<��$<�<9v<�<�-	<c<�;H�;�Z�;T�;K��;���;K�;�7�;��;`b�;�>�;�;���;M�;��;_�s;w`;�3P;
(D;��:;F�2;˦);:;�;qm�:{��:
��:uHh:(8:�6�9,my9�G29��#9�@+9�#9�?�8�Vq�� 8�%<ѹMQ+�lSo���a���_º�ɺ�?Ǻ����2���2������Vr�]e���j��›.����f��y���ѺR(ۺXsܺ��ֺ��̺��ºr���M����\ĺg�պ����\V��G��� ���"�b/!�V���W��]��F��#�ɿ/��?�&FP��a��q�Ϝ}��炻�����䃻�_���f{��Ys��Pl�#h���g��%l���t��L���Ɔ�U������0z��Yӓ�����꜐�7Ȏ�����T��_Ғ��O��v	��b
���Z���,���  �  �0 = =5 =Gq =E� =�� =�` =x��<=��<|��<�h�<]#�<�&�<Χ�<���<��<���<���<���<^��<��<�:�<��<=7�<���<&@�<��<o<�<b�<# �<Zj�<��<&��<̍�<���<�a�<�U�<l��<6��<c�<�z�<�f�<���<���<z�<��<̀�<u}�<D��<'��<���<���<��<���<���<���<o�<45�<v��<$��<��<���<���<���<��<��<]�<g �<o��<��<��<?��<�4�<���<�`�<6��<��<0��<��<r��<M��<�`�<E)�<O|�<�k�<��<���<ǐ�<O#�<�4�<椯<^t�<d��<���<$��</��<�<�<�J�<���<�X�<�8�<�o�<EǏ<� �<5�<�@�<�
�<�L�<�0�<-��<��{<f�v<6xr<Fgo<�%m<�?k<&'i<�Jf<b=b<��\<PCV<��N<�}G<|@<�g:<M�5<V�1<IN/<--<0�*<��'<f�#<SF<i�<�<L�<(��;̺�;\u�;&��;Dc�;���;ߴ�;e��;L7�;���;x��;�B�;���;D�;F	�;C�;�l;�Y;|J;xv?;�7;i�1;1*;Ͷ;��;���:Hy�:�v�:��X:C3:�,�9�+9�nz8,^8Uٗ8VԦ8��28?9r���m��n<�?���V��s����кhFغ�7պ]ɺѶ�l衺�E����I9s��z�ʖ��qQ�������κ��ߺzl�@���޺jHѺDEú}�����q��GGԺ�ﺕ~�۶��  �qW'���)��<(�9$�8��+�G$ ��2'��3���B�I�T�og��w�nZ��o����1���G���X���0���kw���o��Wk��ak��kp���y��X���1���L��L�������@_��NP��2`�������g���l�����!�����������Ю��I���  �  T�<��<z��<�.�<U��<a��<��<�k�<V�<���<�q�<���<��<{�<�&�<�</��<���<��<d<�<���<f �<�#�<�m�<��<`r�<��<</�<�9�<�;�<� �<'��<�f�<��<Ƥ�<$]�<Z��<3��<���<�;�<���<�}�<���<�d�<���<��<���<���<��<�$�<���<}��<�4�<���<�<��<�G�<���<�l�<z��<T#�<E�<���<x�<�2�<��<�L�<�S�<H��<�p�<��<K��<~��<�*�<k��<n�<�L�<���<*�<�.�<���<���<��<��<~��<�֮<�c�<l4�<�έ<^ˬ<��<Y#�<���<[e�<��<�З<��<5�<���<y�<�<lw�<��<~�<���<�|�<Nu�<�x<Aw<so<��g<fCb<�k^<�V\<Ǜ[<ـ[<z[<7mY<��U<��O< �G<
�><u5<g�,<\�%<Vc <+<Z�<�I<�<�(<��<��<�<�<k�;���;�z�;�Q�;���;鶷;�R�;�"�;	�;֪�;���;��;;Е;�y�;=Kq;��O;�;/;|�;��:��:_'�:�D�:��:�:�:��:'�o:���9�Y��Vz�/ej��̚�����]����𲕺�"��6�n�Z�m�����Wٜ�O���?���]�����| �������
�g*��A��ٺ�ںV%��)����;$)��:�)OE��NI�*�E�Y�;���-�0��>��>���i"�J6�{UL��Ta�y�q��.{��	}�h�w�]�m��za�15W���Q��LS�O�[�m�j�25}�K����ߑ��*��/����(��ӫ��)Ι����*k����������Kތ���������q���SL��-���S���{��l=��o��,t��S?��$d��we��-ܫ�]L���I���ʻ�Dջ��ܻ�  �  ��<	��<rT�<���<���<c��<�0�<H��<�4�<M$�<z��<w8�< 
�<Lk�</��<_�<Z��<���<E�<�q�<�,�<|3�<a�<V��<�p�<���<�}�<4��<���<���<���<v��<��<���<R��<�c�<M�<G��<�7�<��<c�<��<Hx�<	��<��<���<��<���<��<U�<~��<,��<�y�<�:�<p`�<�$�<|��<���<���<��<�^�<%w�<��<$��<�s�<`�<R��<���<�<���<��<B��<�<Ck�<���<Z~�<�P�<B��<���<�Z�<Jǽ<mX�<W|�< |�<s�<kO�<FѮ<w��<d�<v�<�<�Q�<Խ�<N��<�P�<'#�<�f�<OP�<3��<\�<�[�<U��<�(�<�N�<"�<���<㽃<2�<~x<:p<��h<AAc<H[_<~(]<�B\<��[<Z[<�Y<��U<��O<�5H<�D?<�6<[�-<{�&<K[!<�$<C�<W<�<��<i6<��<9�<�f<N�;���;���;l��;=y�;�*�;-��;jU�;��;���;�q�;7��;�ϖ;*��;�Nt;S;�3;S�;9�;�?�:�b�:��:K�:���:&��:V�::�q:��9�+7����\��$��-���z��񝠺*H����{�ff��f���� ���1N��`���8����S.�ڔ�e��� �����k����⺽�ֺe�׺��� ����I�%�h$6��WA��|E��HB�T�8�ы+��������Z��1�!�@�4�HJ��X^�8%n�Pw�xy�xt��j��y^�M�T��O�`�Q��TZ���h�zD{��y����������<��[���$P��3�������͈���劻�ɉ�M���ט�����P��Iq���ƶ��	��U���	���3Ƕ�A���긪��-���M������ѳ��k��&�ɻʫӻ��ڻ�  �  ��<���<դ�<}��<���<m��<���<��<��<���<�e�<��<���<�q�<��<Bb�<N��<���<���<��<J��<���<�<m��<}s�<��<Y��<��< �<a��< ��<4��<��<N;�<M��<pl�<�4�<�@�<J��<h��<o��<+L�<u��<]B�<�H�<���<��<���<=��<9��<
]�<�g�<�7�<x�<[�<.�<���<>��<��<���<���<2��<#v�<k6�<��<<�<=��<f�<�j�<O�<e��<#�<2��<��<��<o��<S�<��<N��< ��<|��<�W�<y��<�ѳ<�ұ<��<��<���<L�<Z��<W��<Jʨ<�C�<�E�<)�<�<g�<�[�<� �<}S�<7�<�t�<���<�Ҋ<bg�<�P�<��<�
�<fz<2�r<��k<�f<D�a<On_<�
^<�*]<��[<�Y<w�U<> P<x�H<�_@<�7< �/<�)<j$<S� <B3<eh<ұ<�8<�c<��<U�<|�<���;EV�;��;���;��;�N�;�y�;v��;Uٰ;�٭;���;��;kp�;�	�;ŗ|;t�\;�>;�#;��;*��:T��:�+�:w��:���:�*�:�ަ:�^w:��:���8e���>�6�o1{��r���@��� ���{���^�eXO�Z�T�Baq�{h�����O�Ժ,h��p��&��5=�
�o�����r�y}ں�*Ϻ��κ�ۺ�9��	���2+�3"6�A�:���8�1�&�%����$C�ܵ�6R�����0� �C�XV��<d��el���m��6i��\`��7V��"N���J�U{M�ilV���d�kv��Q���댻ݺ��J��m���fy���3������i3��s㈻�̇�X���0���s[�����Z>���7��Rx��if�����9�����.k��붦�X/��F��M���n"���9ƻ�=ϻ �ջ�  �  ���<e��<��<�f�<89�<.��<���<���<�O�<Fs�<�X�<M=�<wa�<���<|!�<���<o2�<���<2��<e��<�B�<�U�<���<���<:��<���<l��<6�<��<Ͼ�<��<���<���<"y�<���<^�<�P�<ϱ�<u��<e��<�=�<E:�<���<�A�<��<)%�<��<u�<�A�<�h�<� �<�4�<�>�<�\�<���<���<�<�<�R�<���<;��<���<	��<�	�<q��<��<�a�<�8�<���<�^�<�Q�<]��<N��<�G�<���<���<E��<y:�<��<���<{R�<Iy�<c��<�k�<���<�ҳ<'��<���<���<f��<"o�<�9�<kZ�<��<��<b/�<�\�<��<��<�<���<Dq�<>s�<E��<5w�<�<*�<B{�<X�<i�}<�uv<��o<�$j<N�e<}�b<�w`<��^<۲\<��Y<�U<�%P<�ZI<�A<�:<��2<�,<�(<f�$<��"<��!<H <1+<j�<�<�<[	<�Z<� �;FR�;z%�;!�;:y�;��;^�;`��;+ְ;��;���;v��;�r�;o�;I�j;]�M;��3;�/;;;��;���:JF�:�W�:���:�q�:��{:�:��T9��3��& ���<�~�^�f�g��]��}I���7��L2���>��@^����i���2;ĺ�*����Dj�����M�!��ø�/@�	к'�ź�IĺAͺd�������8�@S�]�%�#+��+�+9&������i$�a�����G��&,���;�y�J�,V�.�\�N�]���Y���R�`�J�&aE��ED� rH��Q��_�xo����(���X�Eʑ��r���Ӓ�[��hΌ��+��k��fk��IɆ�͊��?���U���š�B#���Y���ڰ������a����������|���p��%$��
[��@�������Ȼbλ�  �  ;;�<�;�<b��< �<݄�<C��<��<i#�<���<��<+K�<��<���<Z��<"��<���<S��<� �<���<�I�<���<���<0j�<
��<<�<՗�<���<f�<�O�<��<ě�<���<5;�<#��<���<��<�5�<���<;��</*�<��<^�<�0�<�x�<�<ź�<N.�<s7�<)��<I��<��<2��<}M�<���<<v�<��<��<��<S�<��<z��<�#�<p�<�Q�<���<�u�<���<��<C��<D��<���<��<���<���<���<G��<���<���<~��<$��<Sb�<�+�<�K�<'�<1�<c��<`��<�\�<h�<��<{��<뽩<bv�<��<V�<�֛<���<�Õ<�Y�<�_�<�ȏ<�u�<m>�<���<�x�<���<�Y�<О�<Ӈ�<d�z<St<R�n<��i<f</�b</`<�]<�xY<6U<P�O<��I<��B<�@<<�6<��0<]�,<`W)<9�&<o%<��"<��<$�<H�<��<�R
<kD<gT�;ѿ�;�g�;>��;e��;�X�;�o�;�\�;zv�;m�;ǎ�;y�;L��;b͉;�y;�-_;@F;�^0;UA;��;�	;� �:���:f�:-j�:��y:��%:(v�9����򀊹�s�/���( �R����-Y��x��m.��P���}�)����,����˺��ߺ���3����E�캗$���ӺƙǺ���O���������κ`8������	�Ʉ����o-�����������W�n���<�ɕ(�� 4�,�>��F���J�@K�3`H�+�C��F?�uJ=��	?�^�D��JN�R�Z�PYh�fv�����Sֆ�hn��DB���a��q��'ވ�t��ވ������🄻s��#C������=���p&��~H�������Щ�����nV��@���'�������꫻ϰ�0Ƕ�V�T»�/ƻ�  �  �E�<yB�<�d�<��<�f�<���<-�<M�<���<�f�<}��<N��<~u�<`�<���<?W�<�#�<�&�<�M�<���<��<���<��<7�<�:�<>�<���<�r�<S�<sx�<���<��<�d�<A4�<���<�i�<i��<U��<�<T8�<���<�I�<f@�<}q�<s��<h��<��<���<'��<��<ۜ�<a]�<"�<:�<��<�T�<���<��<���<��<��<4B�<Mc�<�L�<u��<@�<���<'@�<:n�<s��<u��<z+�<k��<$>�<���<N�<�&�<��<Lj�<`��<���<tU�<��<�Թ<�	�<�x�<n��<w[�<�q�<�+�<t��<ٯ�<���<}t�<cI�<�3�<�G�<S��<J�<��<���<�9�<���<d�<�v�<+��<<B{�<�<�"~<�dx<�r<�m<[
i<X�d<�`<$�\<�\X<I�S<��N<
I<bhC<~�=<a�8<�M4<��0<XO-<�*<_�'<�$<g� <�<��<K
<��
<L�<���;���;���;��;��;�E�;���;��;V��;7Z�;���;cP�;T֗;�;���;�n;�W;��@;ߦ,;Џ;DS
;�j�:���:�l�:��:��k:$%:���9�i9�����@b�]ǣ������ι�ܹ�I�����OC-��~Q�s�y� ���ڼ��e����Lƺ�к�a׺J�ٺ\�׺�Ӻ;o̺pźH�����������pBĺE�к^���T��'�X9
�3@��$�4m�Q�9�������!��'��.���4���8��:�X�:�\=9�j7�2�6��8�.�=��E��cN��X�$�c���n�J7x�Z���.���8���B��*j��!셻|���M��C�_������􈻣R��_�����������c���P˥�_񦻏��L���U���*������Y����z��7����⾻�  �  ���<Ϋ�<х�<�-�<��</��< ��<�^�<�7�<,&�<�2�<^�<���<d��<�T�<��<�8�<5��<�h�<M-�<�<>�<9��<���<�~�<d��<]��<9��<��<,��<ű�<B��<
�<�l�<��<L�<b��<�_�<��<��<C��<���<���<���<̺�<�r�<���<��<��<��<��<�A�<Ȅ�<z��<
V�<��<+_�<-��<l��<P5�<���<���<���<m��<yb�<��<UC�<�&�<,��<���<�!�<2�<�8�<M:�<�2�<��<���<S��<���<�D�<��<|��<��<0�<rl�<]��<*��<���<'5�<���<h˫<���<P2�<�x�<;Ѡ<�7�<�<��<���<�%�<�Ƒ<W��<r�<���<>ȉ<��<�m�<���<���<O/�<R9{<��u<*_p<|�j<��e<�x`<�a[<�WV<!YQ<�iL<��G<��B<}�><�|:<j�6<IW3<b0<[�,<��(<��$<U�<��<V<��<n
<<;��;��;c��;|y�;ʎ�;���;'��;꾻;��;��;��;G�;2�;NY�;�a�;�x;?c;Z�L;��6;Q!;��;�I�:��:�C�:zy�:�O:Tq:o�9%gT9_o�8��6�����P��>��$������!^��B�-�g�����D���f��?Y������bø�����;]ĺD�ȺB�˺Kͺ�̺�ʺ �ǺPwźpź߂ɺ�jҺ�Yߺ}�`'������4�������b��o �4$���'��*�!+-��.�uy/�s/��&/��F/�t�0��C4��8:�V
B���J���S��\���c��j�v�o��0u��z���~��l��K��Ԅ��ꅻ͉���І�����do�������ي��F�������1��ԛ�U*��p���v�����$C���ԯ�<��Ws���f��������������  �  O; =_% =���<K �<��<�}�<l�<���<%��<8G�<i��<���<�V�<���<�s�<��<F��<���<���<%4�<���<
��< ��<���<���<<��<�X�<?��<�|�<C:�<��<��<XF�<G2�<~Y�<��<fp�<�\�<�}�<���<.�<NS�<�p�<lQ�<���<
�<��<b��<w��<H��<	��<��<B]�<I�<6,�<j��<�w�< ��<���<��<�J�<���<vA�<��<��<�	�<���<=5�<�$�<���<���<��<E.�<B��<�(�<���<�Z�<<+�<�(�<�R�<���<n	�<�u�<Tһ<��<��<���<R�<�!�<(�<�D�<"��<�!�<Z�<\Ӡ<�<N��<�:�<��<��<N�<�G�<橌<'X�<x^�<���<�F�<��<�U�<�w�<�v|<.Sw<��q<h�k<�ce<�-_<&Y<�uS<w5N<$tI<6E<�sA<
><)�:<c�7<˲4<�21<\2-<\�(<�I#<�<C�<�b<O<��<�u<k <T��;>��;c+�;��;��;�;�;�/�;K�;��;`��;�;�6�;�A�;�a�;�<|;��h;�S;=�;;)5#;��
;0=�:��:mQ�:�u_:�t%:�:�9(�9�'W98��8vF48� �_a����Ϲ�t�)E��p��I���閺�a��鴡��٢�!��3K��|N���G���q���Gͺ9�׺�޺Q��@ߺ�/ں�!Ժ{кg�к�Q׺\+㺴7� �1�����6��z'�ަ,�h90���1��1��
0�L�-�b+���)��)�=�+�k�0�$�8��]B�*�L�l�V��^��/d�i�g���i��kk���m�fq�!6v�l�|��)����//���w��V�������1�����1ˋ�yC��s*��ZK���S���㞻����	���ꮻ�󲻩 �����{
���1������ ��Y���  �  �@ =� =b�<�<^q�<���<��<���<�$�<_��<D�<�U�<ܕ�<��<( �<|?�<���<D|�<���<}��<9��<}�<���<��<v��<���<{��<)��<��<�(�<"��<K��<b�<��<��<���<���<\ �<��<�9�<:��<�W�<�u�<0 �<wK�<��<Jt�<��<��<_��<�F�<>W�<���<5�<���<��<��<9�<���<҆�<�!�<� �<G�<8 �<��<0g�<��<��<M��<&��<=��<�[�<H��<Դ�<2��<���<�y�<(O�<��<4�<���<���<�J�<�ʻ<��<���<3�<���<�b�<"�<�(�<`��<ь�<O١<�Z�<�՞<1�<��<9E�<;;�<��<Պ�<_�<���<�b�<���<�w�<qv�<f�<��<�@|<�ow<%�q<�"k<I(d<.]<~?V<��O<ކJ<�E<7/B<{.?<B�<<�I:<ż7<�4<�0<4=,<�&<k <��<��<�J<1�	<��<��<���;��;�@�;��;��;q�;���;���;�[�;��;���;R�;���;hP�;�l�;M�y;��h;��S;ux;;� ;	;�:�!�:�m:':GK�9��9-T9�39I��8�hR8���.�b���v	�>�F�Ľ���#��B˩�<���厱��ȫ����������ܢ�v���x���kֺ��麽���P: �U ��"��#��H�vۺ!�ں�㺽��0�y��2���5*�Q04�/;�ny>��r>�w;���6�h�0��!,��r)�/�)��L.�Ķ6�BxB�^�O�ٺ\��g���m�R�p���o��_m���j�l�i�Y�k�;mq��qz�������r|��s���	����ꔻ"����r��ө��A7��%����%��u]���ߟ�7���9������u͹��D�����򾻘����f��!���t���  �  [
 =���<�{�<��<Q��<k��<>��<���<q�<�A�<I��<��<�x�<���<�l�<�f�<]��<e��<2��<���<f��<�7�<A[�<��<���<���<!.�<���<��<���<d��<u��<���<�<H��<f�<g�<���<�b�<�f�<S�<���<� �<it�<�B�<��<���<ٷ�<�G�<x�<c[�<���<���<���<ُ�<���<Wb�<@E�< ��<á�<���<P�<��<̲�<q��<w�<��<wi�<J�<��<�A�<H��<��<t��<�B�<8�<���<m�<���<���<ʣ�<�Ľ<g��<_Q�<�^�<�Ͷ<���<��<�Y�<�٨<�֥<�u�<���<��<��<��<�-�<�0�<y��<x-�<jg�<��<�Љ<���<t.�<�v�<�b�<���<z�<�,~<o{<ǚv<��p<��i<�_b<]�Z<)'S<�sL<n�F<�RB<%�><`�<<�:<[�8<��6<K�3<�/<�^*<��#<x�<��<�6<�	<L�<ب<9� <H��;�Z�;�5�;�j�;��;��;�h�;{�;z��;�;㿎;���;Ƶ�;��;7~};x�s;�e;�P;S8;h�;��: [�:Ո:�Q5:AI�9�o9��8�*�8��R8o"8�N6k���/m�t��7��逺���o���̺�2к�ɺպ�����i����ɘ��d�������tǺg���V �`����c����.�;���K캆>溼�꺑l��:{��*��&��5���A�P�I���L���K�!vF���>���6��0�ڿ,�5�-�T�4�m@��UO���_��n��Iy���~��~��ez�݀s��l��h��ji�!�o�~�z����$J���Ԕ�<�������������$����#���������ᕻ���)O������8$��Ժ�����ĻKƻ9Ż��»���V���NA���  �  �y�<i��<py�<�o�<�
�<]��<���<c��<EC�<���<���<��<t,�<��<�|�<�T�<|e�<��< ��<UZ�<���</�<\W�<�+�<�]�<l��<�<�<�E�<��<��<��<���<4��<M��<w<�<���<��<�4�<wJ�<���<#��<�T�<�]�<���<�%�<��<T��<���<<�<~�<���<�q�<���<�;�<_�<���<=l�<[�<��<��< R�<�`�<"�<��<"��<d��<���<x<�<C=�<�b�<Ơ�</�<Z��<�i�<6��<���<���<���<�I�<sD�<���<��<N�<��<���<Vٵ<&b�<.y�<�{�<�Ϧ<�ã<G��<�
�<�4�<"��<��<8�<N?�<P��<��<�Ő</n�<�U�<�ل<�3�<Gs�<�~<~<�i}<� |<�y<gu<¡o<��h<,�`<�OX<jP<�gI<�C<?<?<�+<<.:<��8<�l7<�}5<��2<�!.<3M(<�?!<p�<��<N<�<��<�$�;���;$��;�<�;9�;M��;��;�~�;�l�;�)�;�a�;2_�;fІ;컀;��z;�}w;�s;��l;r�_;�}L;�R3;��;���:OT�:�Je:�
:�qr9!zV82J)�݄��jU�9�'�U9���T"�ȩ�Ǧ�I<e�훜�N@º��ݺ�B�\=�a�ߺ��ʺ�U�������D��毝�����Ϻ���jQ�1�bO!��"����b�F	�b���c�����j����]��Eu/��@�O�M�}7V��dY��*W�ssP���F�t=��+5��w1�px3�O�;���I���[�Bhn���~�x̄�����	��S���?z�zp��}i���h�8�o�X}����]���Cؚ��Ρ�񪥻*������Q\�����S)���2��8U���j%���E������PG���ƻ2�ʻ�$̻��ʻTǻQ�»w���i����  �  ���<�B�<���<�u�<���<<`�<ke�< 9�<���<@��<��<i~�<���<���<�t�<�4�<V�<;]�<���<�5�<{��<%��<g��<��<E<�<���<��<(��<m�<2��<�v�<3�<���<A��<"4�<Q��<���<�L�<e��<���<P�<��<N��<��<{O�<p�<G��<g�<��<�!�<�]�<:m�<��<���<�)�<���<�`�<[��<��<~��<�S�<y)�<���<�:�<7��<�i�<��<�[�<��<��<t�<���<�=�<���<5��<��<���<��<�G�<�]�<�ͼ<�J�<X��<�(�<��<,�<5s�<�V�<N.�<4h�<bX�<�)�<f۞<�A�<��<���<��<�6�<�o�<ﭔ<�B�<ա�<�G�<Й�<7׀<."~<aV|<��{<dq{<��z<pYx<�et<(�n<�lg<�6_<�V<��N<�[G<��A<E*=<%A:<w~8<�a7<�A6<�v4<xt1<��,<�&<�C<B&<�;<�O<]�<
��;���;�C�;?��;�%�;���;q��;3N�;:?�;��; ��;Q�;@�;�\�;��v;��p;5�n;;�l;��f;�Q[;��H;pw/;�,;�x�:��:;G:�\�9v��81��������#��9���׸� �*�c���ҹ`	0����C��]�׺�F���� ��������׈ֺ����M飺r��k]��
��kֺ���9�5�"�e,���-�h�(�gU���	6�}�������=Q����"���5��GG�]U��^���a�I�^�'eW��L�k�A��B9�,e5��7�fA�2 Q�*�d�H�x��˄��c���^��*������uy�hs�s�j��5i�
=p��"�����n唻U���ަ��,��*ë���X ������V��Z����a��zz��]������W���;Ļ��ʻ�ϻ�;л��λ��ʻ�Żp���z����  �  ���<7�<�i�<c�<{r�<���<���<���<Ņ�<9�<���<=H�<J��<4��<�n�<Z&�<J��<P!�<fD�<7��<��<�K�<�v�<�j�<���<?�<�;�<�y�<���<M\�<�=�<���<;]�<�K�<���<>$�<b6�<���<�9�<��<���<��<���<^��<���<X��<�*�<���<
V�<Z��</��<��<z��<֗�<Q�<���<(Y�<9��<�{�<ű�<B��<	��<vF�<���<5	�<���<��<��< I�<ڛ�<@��<,M�<���<T�<��<�O�<���<�a�<w�<G�<(��<��<M�<d��<�ѷ<մ<f�<��<F��<��<�ס<��<n�<t�<�ȝ<��<yܜ<a0�<�e�<���<0�<OV�<��<q'�<�[�<1'}<�e{<�z<J�z<*�y<��w<�t< Jn<g<Z�^<�V<��M</�F<��@<�p<<M�9<Y�7<H�6<��5<�4<C1<i,<6"&<e�<�K<�H<Q<q�<U��;/�;#�;"��;���;���;���;l�;��;,�;�f�;YV�;�l�;��~;��r;G9m;gzk;��i;
�d;)�Y;�CG;� .;�s;�a�:$?�:�n<:]��9���8f_�PCD��3G�i#��������^}�CK�6�9�� ����rߺ�-��{���j�\�����ں[~���G������_Ξ�G��5ٺ��D�(S&�r�/���1�Ǧ,�d�!�u������X��~ ������_�$�b�7��I��KX�lva�.�d�5�a��Y�,�N�߮C�w�:���6�[�9��C���S���g� F|�]���8^���A��Va��j�������=t��%k�hi�c�p��������?��,���筨�c ������J򪻈֥���Ѕ��Z���V,���:���3��9���%���SŻi_̻Îл-�ѻ�ϻ	�˻,�ƻ����oh���  �  ���<�B�<���<�u�<���<<`�<ke�< 9�<���<@��<��<i~�<���<���<�t�<�4�<V�<;]�<���<�5�<{��<%��<g��<��<E<�<���<��<(��<m�<2��<�v�<3�<���<A��<"4�<Q��<���<�L�<e��<���<P�<��<N��<��<{O�<p�<G��<g�<��<�!�<�]�<:m�<��<���<�)�<���<�`�<[��<��<~��<�S�<y)�<���<�:�<7��<�i�<��<�[�<��<��<u�<���<�=�< ��<7��<��<���<��<�G�<�]�<�ͼ<�J�<]��<�(�<��<2�<<s�<�V�<T.�<:h�<hX�<�)�<k۞<�A�<��<���<��<�6�<�o�<�<�B�<ѡ�<�G�<̙�<2׀<#"~<UV|<��{<Xq{<��z<eYx<�et<�n<�lg<�6_<�V<��N<�[G<��A<G*=<(A:<|~8<�a7<�A6<�v4<�t1<��,<�&<�C<N&<�;<�O<h�<��;���;�C�;I��;�%�;���;q��;/N�;3?�;��;�;@�;@�;�\�;X�v;��p;�n;�l;_�f;�Q[;e�H;Ew/;�,;�x�:e�:�G:5\�9*��8������w�#��9�!�׸2� �L�c���ҹd	0����D��]�׺�F���� ��������׈ֺ����L飺r��k]��
��kֺ���9�5�"�e,���-�h�(�gU���	6�}�������=Q����"���5��GG�]U��^���a�I�^�'eW��L�k�A��B9�,e5��7�fA�2 Q�*�d�H�x��˄��c���^��*������uy�hs�s�j��5i�
=p��"�����n唻U���ަ��,��*ë���X ������V��Z����a��zz��]������W���;Ļ��ʻ�ϻ�;л��λ��ʻ�Żp���z����  �  �y�<i��<py�<�o�<�
�<]��<���<c��<EC�<���<���<��<t,�<��<�|�<�T�<|e�<��< ��<UZ�<���</�<\W�<�+�<�]�<l��<�<�<�E�<��<��<��<���<4��<M��<w<�<���<��<�4�<wJ�<���<#��<�T�<�]�<���<�%�<��<T��<���<<�<~�<���<�q�<���<�;�<_�<���<=l�<[�<��<��< R�<�`�<"�<��<"��<d��<���<x<�<C=�<�b�<Ǡ�<0�<\��<�i�<8��<���<���<���<�I�<zD�<���<��<X�<��<���<aٵ<2b�<:y�<�{�<�Ϧ<�ã<P��<�
�<�4�<(��<��<:�<N?�<O��<��<�Ő<(n�<�U�<�ل<�3�<<s�<�~<�~<�i}<� |<ˑy<jgu<��o<��h<�`<�OX<jP<�gI<�C<B<?<�+<<
.:<��8<�l7<�}5<��2<�!.<JM(<�?!<��<��<d<�<��<%�;���;9��;�<�;$9�;M��;���;�~�;�l�;�)�;�a�;_�;<І;���;i�z;P}w;��s;W�l;�_;�}L;@R3;E�;"��:�S�:-Je:�	:�or9sV8�O)�߄��mU�Y�'�:��U"�ȩ�Φ�M<e��O@º��ݺ�B�\=�a�ߺ��ʺ�U�������D��毝�����Ϻ���jQ�1�bO!��"����b�F	�b���c�����j����]��Eu/��@�O�M�}7V��dY��*W�ssP���F�t=��+5��w1�px3�O�;���I���[�Bhn���~�x̄�����	��S���?z�zp��}i���h�8�o�X}����]���Cؚ��Ρ�񪥻*������Q\�����S)���2��8U���j%���E������PG���ƻ2�ʻ�$̻��ʻTǻQ�»w���i����  �  [
 =���<�{�<��<Q��<k��<>��<���<q�<�A�<I��<��<�x�<���<�l�<�f�<]��<e��<2��<���<f��<�7�<A[�<��<���<���<!.�<���<��<���<d��<u��<���<�<H��<f�<g�<���<�b�<�f�<S�<���<� �<it�<�B�<��<���<ٷ�<�G�<x�<c[�<���<���<���<ُ�<���<Wb�<@E�< ��<á�<���<P�<��<̲�<q��<w�<��<xi�<J�<��<�A�<J��<��<w��<�B�<8�<���<#m�<���<ȑ�<֣�<Ž<v��<nQ�<�^�<�Ͷ<ɥ�<��<Z�<�٨<�֥<�u�<���<��<��<��<�-�<�0�<w��<t-�<dg�<��<�Љ<���<e.�<�v�<�b�<���<i�<�,~<O{<��v<��p<��i<�_b<M�Z<'S<�sL<l�F<�RB<.�><n�<<'�:<q�8<��6<g�3<�/<�^*<��#<��<ݼ<�6< �	<g�<�<L� <f��;�Z�;�5�;�j�;��; ��;�h�;U�;L��;�;���;p��;���;q�;�}};��s;Te;��P;�8;��;O��:UZ�:�Ԉ:Q5:�G�9��o9���8�'�8B�R8l"8��M6$���C/m�3t��7��逺���o���̺�2к�ɺպ�����i����ɘ��d�������tǺg���V �`����c����.�:���K캅>溼�꺑l��:{��*��&��5���A�P�I���L���K�!vF���>���6��0�ڿ,�5�-�T�4�m@��UO���_��n��Iy���~��~��ez�݀s��l��h��ji�!�o�~�z����$J���Ԕ�<�������������$����#���������ᕻ���)O������8$��Ժ�����ĻKƻ9Ż��»���V���NA���  �  �@ =� =b�<�<^q�<���<��<���<�$�<_��<D�<�U�<ܕ�<��<( �<|?�<���<D|�<���<}��<9��<}�<���<��<v��<���<{��<)��<��<�(�<"��<K��<b�<��<��<���<���<\ �<��<�9�<:��<�W�<�u�<0 �<wK�<��<Jt�<��<��<_��<�F�<>W�<���<5�<���<��<��<9�<���<҆�<�!�<� �<G�<8 �<��<0g�<��<��<M��<'��<>��<�[�<J��<״�<7��<���<�y�<1O�<��<A�<���<���<�J�<�ʻ<��<Σ�<H�<¹�<�b�<5�<�(�<p��<ߌ�<[١<�Z�<�՞<5�<��<7E�<6;�<��<ʊ�<_�<���<�b�<{��<�w�<]v�<�e�<��<�@|<�ow<�q<�"k<1(d<]<p?V<��O<܆J<�E<B/B<�.?<X�<<�I:<�7<�4<+�0<\=,<F�&<Hk <��<��<�J<Q�	<�<��<���;��;�@�;��;��;�p�;���;T��;i[�;��;���;�Q�;H��;P�;4l�;��y;�h;�S;�w;;�� ;�;L�:� �:ߧm:�':�I�9x�9B+T9�29c��8�eR8����.�{���v	�C�F�Ž���#��B˩�;���厱��ȫ����������ܢ�v���x���kֺ��麽���P: �U ��"��#��H�vۺ!�ں�㺽��0�y��2���5*�Q04�/;�ny>��r>�w;���6�h�0��!,��r)�/�)��L.�Ķ6�BxB�^�O�ٺ\��g���m�R�p���o��_m���j�l�i�Y�k�;mq��qz�������r|��s���	����ꔻ"����r��ө��A7��%����%��u]���ߟ�7���9������u͹��D�����򾻘����f��!���t���  �  O; =_% =���<K �<��<�}�<l�<���<%��<8G�<i��<���<�V�<���<�s�<��<F��<���<���<%4�<���<
��< ��<���<���<<��<�X�<?��<�|�<C:�<��<��<XF�<G2�<~Y�<��<fp�<�\�<�}�<���<.�<NS�<�p�<lQ�<���<
�<��<b��<w��<H��<	��<��<B]�<I�<6,�<j��<�w�< ��<���<��<�J�<���<vA�<��<��<�	�<���<>5�<�$�<���<���<��<H.�<F��<�(�<���<�Z�<F+�<�(�<S�<���<�	�<�u�<iһ<��<��<خ�<i�<�!�<(�<�D�<5��<"�<h�<gӠ<�<R��<�:�< ��<��<E�<�G�<ש�<X�<e^�<���<xF�<��<�U�<�w�<xv|<Sw<��q<H�k<�ce<~-_< &Y<�uS<u5N<*tI<6E<�sA<#><H�:<��7<�4<�21<�2-<��(<�I#<�<n�< c<*O<��<�u<k <p��;L��;c+�;���;Ԙ�;�;�;�/�;�;j�;��;��;96�;4A�;�a�;/<|;��h;S;��;;�4#;+�
;G<�:��:�P�:vt_:t%:89�9'�9v&W9��8sC48$�i �{a����Ϲ�t�+E��p��I���閺�a��贡��٢�!��3K��{N���G���q���Gͺ9�׺�޺Q��@ߺ�/ں�!Ժ{кg�к�Q׺\+㺴7� �1�����6��z'�ަ,�h90���1��1��
0�L�-�b+���)��)�=�+�k�0�$�8��]B�*�L�l�V��^��/d�i�g���i��kk���m�fq�!6v�l�|��)����//���w��V�������1�����1ˋ�yC��s*��ZK���S���㞻����	���ꮻ�󲻩 �����{
���1������ ��Y���  �  ���<Ϋ�<х�<�-�<��</��< ��<�^�<�7�<,&�<�2�<^�<���<d��<�T�<��<�8�<5��<�h�<M-�<�<>�<9��<���<�~�<d��<]��<9��<��<,��<ű�<B��<
�<�l�<��<L�<b��<�_�<��<��<C��<���<���<���<̺�<�r�<���<��<��<��<��<�A�<Ȅ�<z��<
V�<��<+_�<-��<l��<P5�<���<���<���<n��<zb�<��<UC�<�&�<,��<���<�!�<2�<�8�<Q:�<�2�<��<���<]��<���<�D�<��<���<��<+0�<�l�<u��<B��<��<>5�<ʐ�<}˫<���<a2�<�x�<FѠ<�7�<���<��<���<�%�<�Ƒ<J��<r�<퉋<*ȉ<t�<nm�<���<���<8/�<%9{<��u<_p<Z�j<��e<�x`<va[<�WV<YQ<�iL<��G<��B<��><}:<��6<rW3<�0<��,<*�(<�$<��<��<8V<��<;n
<3<d��;��;r��;}y�;���;���;���;���;ٚ�;9�;{�;�F�;�1�;�X�;�a�;)�x;�c;��L;W�6;�P!;�;�H�:?��:C�:�x�:)�O:�p:a�9�eT9m�8׭6�P��LP��>��6�����$^��B�-�g�����D���f��?Y������bø�����;]ĺD�ȺA�˺Kͺ�̺�ʺ �ǺOwźpź߂ɺ�jҺ�Yߺ}�`'������4�������b��o �4$���'��*�!+-��.�uy/�s/��&/��F/�t�0��C4��8:�V
B���J���S��\���c��j�v�o��0u��z���~��l��K��Ԅ��ꅻ͉���І�����do�������ي��F�������1��ԛ�U*��p���v�����$C���ԯ�<��Ws���f��������������  �  �E�<yB�<�d�<��<�f�<���<-�<M�<���<�f�<}��<N��<~u�<`�<���<?W�<�#�<�&�<�M�<���<��<���<��<7�<�:�<>�<���<�r�<S�<sx�<���<��<�d�<A4�<���<�i�<i��<U��<�<T8�<���<�I�<f@�<}q�<s��<h��<��<���<'��<��<ۜ�<a]�<"�<:�<��<�T�<���<��<���<��<��<4B�<Mc�<�L�<u��<A�<���<'@�<:n�<t��<v��<}+�<n��<)>�<���<T�<�&�<��<Xj�<n��<��<�U�< �<�Թ<�	�<�x�<���<�[�<�q�<�+�<���<쯩<���<�t�<mI�<�3�<�G�<T��<H�<��<~��<x9�<���<S�<�v�<��<���<,{�<��<�"~<fdx<��r<�m<;
i<<�d<ν`<�\<�\X<H�S<��N<�
I<uhC<��=<�8<�M4<��0<�O-<�*<��'<K�$<�� < <��<o
<�
<f�<���;��;���;��;���;�E�;���;��;��;�Y�;N��;P�;�՗;��;g��;Pn;@W;,�@;>�,;=�;�R
;�i�:��:�k�:���:��k:`#%:���95h9�����Ab��ǣ����ι�ܹ�I�����PC-��~Q�r�y�����ڼ��e����Lƺ�к�a׺I�ٺ[�׺�Ӻ:o̺pźH�����������pBĺE�к^���T��'�X9
�3@��$�4m�Q�9�������!��'��.���4���8��:�X�:�\=9�j7�2�6��8�.�=��E��cN��X�$�c���n�J7x�Z���.���8���B��*j��!셻|���M��C�_������􈻣R��_�����������c���P˥�_񦻏��L���U���*������Y����z��7����⾻�  �  ;;�<�;�<b��< �<݄�<C��<��<i#�<���<��<+K�<��<���<Z��<"��<���<S��<� �<���<�I�<���<���<0j�<
��<<�<՗�<���<f�<�O�<��<ě�<���<5;�<#��<���<��<�5�<���<;��</*�<��<^�<�0�<�x�<�<ź�<N.�<s7�<)��<I��<��<2��<}M�<���<<v�<��<��<��<S�<��<z��<�#�<p�<�Q�<���<�u�<���<��<D��<E��<���<��<���<���<���<M��<���<���<���<1��<bb�<�+�<�K�<:�<E�<w��<u��<�\�<}�<��<���<���<pv�<��<
V�<�֛<���<�Õ<�Y�<�_�<�ȏ<�u�<_>�<���<�x�<���<�Y�<���<���<<�z<�Rt<.�n<v�i<�f<�b<`<�]<�xY<5U<U�O<��I<��B<�@<<6<��0<��,<�W)<a�&<�%<��"<�<J�<l�<��<�R
<�D<�T�;��;�g�;>��;Y��;�X�;go�;h\�;Bv�;,�;���;�x�;���;͉;6�y;�,_;`?F;^0;�@;I�;
	;���:%��:oe�:�i�:ĕy:��%:<u�9�ї�q���t�N���( �_���2Y��x��m.��P���}�)����,����˺��ߺ���3����E�캗$���ӺƙǺ���O���������κ`8������	�Ʉ����o-�����������W�n���<�ɕ(�� 4�,�>��F���J�@K�3`H�+�C��F?�uJ=��	?�^�D��JN�R�Z�PYh�fv�����Sֆ�hn��DB���a��q��'ވ�t��ވ������🄻s��#C������=���p&��~H�������Щ�����nV��@���'�������꫻ϰ�0Ƕ�V�T»�/ƻ�  �  ���<e��<��<�f�<89�<.��<���<���<�O�<Fs�<�X�<M=�<wa�<���<|!�<���<o2�<���<2��<e��<�B�<�U�<���<���<:��<���<l��<6�<��<Ͼ�<��<���<���<"y�<���<^�<�P�<ϱ�<u��<e��<�=�<E:�<���<�A�<��<)%�<��<u�<�A�<�h�<� �<�4�<�>�<�\�<���<���<�<�<�R�<���<;��<���<	��<�	�<q��<��<�a�<�8�<���<�^�<�Q�<^��<P��<�G�<���<���<J��<:�<��<���<�R�<Uy�<p��<�k�<���<�ҳ<8��<��<���<w��<2o�<�9�<xZ�<��<��<j/�<�\�<��<��<�<���<>q�<6s�<:��<(w�<�<�<2{�<�W�<G�}<suv<��o<�$j<2�e<e�b<�w`<�^<в\<��Y<�U<�%P<�ZI<#�A<�:<��2<�,<�(<��$<�"<ɢ!<>H <R+<��<�<�<r	<�Z<� �;ZR�;�%�;!�;0y�;��;�]�;:��;�հ;K�;d��;7��;rr�;*�;��j;��M;,�3;B/;�;v�;2��:�E�:W�:��:�q�:�{:k�:x�T9��3��& ��<���^�w�g�#�]��}I���7��L2���>��@^����i���2;ĺ�*����Cj�����M�!��ø�/@�	к'�ź�IĺAͺd�������8�@S�]�%�#+��+�+9&������i$�a�����G��&,���;�y�J�,V�.�\�N�]���Y���R�`�J�&aE��ED� rH��Q��_�xo����(���X�Eʑ��r���Ӓ�[��hΌ��+��k��fk��IɆ�͊��?���U���š�B#���Y���ڰ������a����������|���p��%$��
[��@�������Ȼbλ�  �  ��<���<դ�<}��<���<m��<���<��<��<���<�e�<��<���<�q�<��<Bb�<N��<���<���<��<J��<���<�<m��<}s�<��<Y��<��< �<a��< ��<4��<��<N;�<M��<pl�<�4�<�@�<J��<h��<o��<+L�<u��<]B�<�H�<���<��<���<=��<9��<
]�<�g�<�7�<x�<[�<.�<���<>��<��<���<���<2��<#v�<k6�<��<<�<=��<g�<�j�<O�<f��<#�<4��<��<��<r��<#S�<��<T��<'��<���<�W�<���<�ѳ<�ұ<(��<��<���<X�<e��<a��<Tʨ<�C�<�E�</�<�<g�<�[�<� �<zS�<7�<�t�<���<�Ҋ<Xg�<�P�<��<�
�<�ez<�r<޶k<�f<1�a<>n_<y
^<�*]<��[<ܾY<v�U<A P<~�H<�_@<��7<�/<)<~$<i� <Y3<}h<�<�8<�c<��<g�<��<���;ZV�;��;���;��;�N�;�y�;a��;:ٰ;`٭;k��;��;?p�;�	�;d�|;�\;B>;L#;~�;���:���:K+�:���:��:U*�:Pަ:^w:M�:���8����c�6��1{��r���@��� ���{���^�fXO�Z�T�Baq�{h�����O�Ժ,h��p��&��5=�
�o�����r�y}ں�*Ϻ��κ�ۺ�9��	���2+�3"6�A�:���8�1�&�%����$C�ܵ�6R�����0� �C�XV��<d��el���m��6i��\`��7V��"N���J�U{M�ilV���d�kv��Q���댻ݺ��J��m���fy���3������i3��s㈻�̇�X���0���s[�����Z>���7��Rx��if�����9�����.k��붦�X/��F��M���n"���9ƻ�=ϻ �ջ�  �  ��<	��<rT�<���<���<c��<�0�<H��<�4�<M$�<z��<w8�< 
�<Lk�</��<_�<Z��<���<E�<�q�<�,�<|3�<a�<V��<�p�<���<�}�<4��<���<���<���<v��<��<���<R��<�c�<M�<G��<�7�<��<c�<��<Hx�<	��<��<���<��<���<��<U�<~��<,��<�y�<�:�<p`�<�$�<|��<���<���<��<�^�<%w�<��<$��<�s�<`�<R��<���<�<���<��<B��<�<Dk�<»�<[~�<�P�<E��<���<�Z�<Nǽ<rX�<]|�<|�<s�<qO�<LѮ<}��<j�<|�<�<�Q�<ٽ�<R��<�P�<)#�<�f�<OP�<2��<\�<�[�<R��<�(�<�N�<�<���<ݽ�<,�<rx<-p<��h<6Ac<>[_<u(]<�B\<��[<Z[<�Y<��U<��O<�5H<�D?< 6<c�-<��&<U[!<�$<O�<c<�<��<t6<��<C�<�f<\�;���;���;p��;=y�;�*�;%��;_U�;��;~��;�q�;"��;�ϖ;��;vNt;�S;�3;"�;
�;|?�:�b�:��:�J�:o��:���:1�:��q:���9�+77��Դ\��$��1���z��󝠺+H��{�ff��f���� ���0N��`���8����S.�ڔ�e��� �����k����⺽�ֺe�׺��� ����I�%�h$6��WA��|E��HB�T�8�ы+��������Z��1�!�@�4�HJ��X^�8%n�Pw�xy�xt��j��y^�M�T��O�`�Q��TZ���h�zD{��y����������<��[���$P��3�������͈���劻�ɉ�M���ט�����P��Iq���ƶ��	��U���	���3Ƕ�A���긪��-���M������ѳ��k��&�ɻʫӻ��ڻ�  �  ��<��<���<!��<H��<'��<���<T:�<-��<�,�<1��<x�<�/�<^v�<��<Aq�<"�<QD�<���<?o�<���<ڟ�<�m�<��<?��<���<Q��<]2�<��<Y�<�t�<Wf�<#��<M�<��<���<���<���<Dw�<H�<f��<�<\�<�
�<Tb�<l��<���<���</L�<��<a�<
��<�Z�<Y�<P/�<���<�v�<���<���<aG�<1��<�g�<6F�<���<�I�<'��<H�<ȏ�<���<��<瘻<M��<~�<g�<���<U��<���<�m�<3,�<$��<�Z�<}J�<�'�<3�<���<�*�<���<tt�<�נ<4��<=�<�<�<�G�<�p�<� �<j̏<Z݋<���<�6�<���<Ҥ�<7��<6)�<�ˀ<�	}<d4v<ym<�-b<�V<(�K<�_B<w�;<S�8</=8<�":<��<<�?<?<w<<�j5<9�+<��<�|<	<���;)�;�@�;�J�;~e�;,�;�b�;/� <Z��;36�;�C�;h=�;9��;��;9�;�i�;���;a��;�E�;���;7ǃ;�Lz;o�d;�E;�;�[�:y�:;��9�M��O�T�7��-2����x
¹t���h�����&s�E&ź����8�CJ]���u�#E��@$}�Cn��(X�7)@��+��������!�'t.���?��CQ�Y9`�*�i�r�l�� i���_� �S��$H��|@��@���H���[��~w�c��������!��ZP��H6��1���ĵ���ʗ�ꊻ]&���y���k؈��8��{��6;����Ļ"�˻��˻�ƻ۽������¢�a����������ro���f��Q���)f��I�������»�F��V����������찻V2���]��Smƻ�Bֻ���K���/A�o��*
�%)�����Tﻄ�㻆gܻ+ۻޔ��b컖v��������I���  �  i��<k��<ŧ�<�R�<�S�<��<���<Wx�<%��<Wg�<�5�<M��<B��<���<���<��<}t�<���<���<���<0��<��<��<҈�<V��<�]�<U��<+
�<-��<"D�<}�<��<��<��<�<��<��<���<���<H��<���<�d�<Z��<��<�#�<+�<�Q�<���<��<��<HU�<K��<U��<|n�<V��<�N�<���<�5�<'6�<���<���<��<��<5�<o��<%�<ڭ�<�L�<�}�<f��<g�<�y�<Z��<J�<�"�<@��<�"�<K��<|t�<L��<K߮<X�<w�<gO�<�^�<~��<P��<��<KN�<�١<IF�<�s�<�~�<���<�j�<�"�<�=�<N�<	��<n��<���<�=�<Af�<*�<s�}<P�v<+�m<Hc<'�W<1"M<�D<ړ=<�&:<�9<P;<��=<S�?<W�?<�k<<��5<�[,<J� <�<�f	<� <&z�;Ԓ�;Wf�;��;�?�;a� <=(<��;�;�.�;�M�;O&�;�|�;q̨;��;Ԇ�;��;���;���;�;�*|;�g;нH;a�!;{��:���:;o�9<�����蹝��ӄ���q����Rh� ׈��2���Fj�f'���
�C4�SkW�=vo��y�}v��+h���R�� <�T�(�0��)����o�,�Q=���N�kF]�еf���i�}&f��O]�i�Q�c2F�B�>�34>��F���X�|s��m��5����٥��ﭻ��G����2��>Ǖ��d��h	���x��G}����󘕻糧A�������AUȻ�ȻK�»_ٸ�2����ߠ�T������jۓ�I���xe��ѩ��	�����;)��f����־��Ժ��㵻�����K?���$����Ļ�Իz�������� �*�Qs����ԁ���|����cۻ�+ڻH�߻p����`��-y�����  �  ���<�C�<���<63�<
��<T!�<���<d�<*u�<���<���<ך�<��<)��<�
�<���<Sf�<�[�<am�<�4�<~R�<���<���<l��<D �<�P�<b��<�f�<�1�<�o�<� �<�w�<z.�<Mo�<���<�s�<|��<*��<�O�<$��<T��<Z��<�9�<�+�<�9�<���<ް�<���<L�<��<���<QW�<t[�<O�<ґ�<�h�<���<�<�<l�<:L�<�r�<�$�<=	�<���<���<`Q�<_`�<�T�<���<�<���<w��<�m�<I��<m"�<���<���<P1�<�4�<��<�O�<���<8�<S��<���<�,�<���<��<���<ķ�<��<��<��<TM�<�-�<��<�J�<�"�<Գ�<h��<�ф<��<g��<Ꮑ<�~<gx<Op<�=f<��[<xtQ<�H<UUB<o�><�=<Q�><Zd@<O�A<f�@<��=<�%7<.<5#<��<�A<��<J��;���;� �;���;�<.�<��<�� <�)�;6p�;��;�}�;'r�;S6�;j��;R�;E�;ӎ;de�;��;�V�;�Ol;��O;v�+;U�;d?�:�G9:�zQ9.J"�����Ᾱx���?6�>D����@�v�׹,�R��Ԯ�����&���F��]�
�f���c�aW���D�O�0��� �b���Q��{�o�'��~7���G��U�X�]�v�`���]��#V���K��VA��|:���9�g2A��5Q���h�U����Ɛ�b���tr��㿦�(W��*#���/���@���.z��s���x��z���%����C>��'/��g��3��鹻�谻����曻Rh���鐻����xb���ݝ������R���I��ز���-��Nົ�t������n��w��������ot��r<λ}�ݻ�:�W�����������r���-��Ld���޻`�ػ��׻Aݻ5�˾��_�� �	�*~��  �  �]�<6��<��<%��<���<���<���<���</��<i��<u��<I��<���<}�<?��<@i�<x��<�`�<�,�<Y��<���<�&�<���<�>�<U>�<6�<��<���<Ξ�<���<s��<��<V��<���<f�<�&�<c��<F�<�7�<k�<���<v�<8��<:x�<�%�<�N�<�v�<=&�<��<O�<f^�<���<�?�<�|�<� �<���<Џ�<J��<�N�<�6�<��<���<܌�<��<{��<���<7��<+�<���<݁�<P �<T��<���<��<8y�<�s�<�O�<�ݿ<�*�<&�<fY�<=Y�<b�<y��<�<R�<`�<+ʣ<P�<'��<7��<�p�<���<���<�$�<�O�<&Ɏ<���<RG�<�`�<��<(΄<r��<�<[�<�+z<��r<fj<G�`<��W<�O<�EI<&EE<tyC<�[C<X�C<�D<Z�B<}�><��8<�a0<��&<�N<�<T<9<֛<�<��<u<x<C|<y�<2$�;��;�C�;��;o��;%��;�6�;f+�;�O�; �;���;T��;���;?�q;;X;118;:J;v9�:��:+#:��9�?m8�ʷD=[����7���7�)���H����4��՘��ߺ9��d�.�xB�L�J�mTI�w�?�$�1��"���������S�z�"��M0�!>�T�I�2Q���S�N2R�qL��<D�?�;��U6�c�5��M;��H��4[��r��K��v���`����B��a��s搻�K��S��r���m�l�r��\���������X�������H^��^�����*ॻ~a��P���A���9�������9��j���`Ģ�X<���G���?��o絻V��#����˯�����󫻡������%-����ƻ�ӻ�"�7l�]������Gq黣J�Y�ٻLaջ�-ջ�ٻ���y������Q���  �  {D�<�f�<d7�<Rm�<���<N��<3�<���<�	�<>��<HD�<>��<K�<�1�<s�<��<]	�<uI�<��<}��<��<�^�<>�<���<�I�<m��<.�<���<ā�<?�<@��<���<�^�<��<�<���<���<���<<�<z��<���<N��<��<��<'C�<d��<��<��<�o�<�:�<�y�<�Q�<���<7��<���<��<T�<A�<8��<���<�w�<r��<p��<���<��<�{�<��<�*�<��<�T�<���<���<���<��<��<+4�<��<X^�<��<��<��<rD�<֔�<]��<Uا<4��<4�<�ܥ<�W�<\Y�<û�<�x�<(��<Wh�<���< ��<�g�<$��<r�< ۈ<T
�<8v�<��<�8�<�&�<{-{<��t<%�m<��e<�^<oW<�Q<��L<iJ<�H<�G<�VF<��C<�?<�9<|�2<D�)<�@!<(7<�<^�<R<�	<h	<ت<�<�w<��<�m�;R��;E��;��;���;���;���;�	�;��;��;��;���;�3�;�Et;��];�B;,$;�;	��:7��:?�D:��:L�9���9�o9��9�I���5��$��*��"��ݟ������=#�^+���+���&��0��������������^�K��1�*���4�/G=���B��E��E�Q�B��>�g�8��W5��4��8�+�A�O�T%`��?r�g?���$���쉻�=��X�������Jt���k�Wji�^�m�iCy�j�,���݀���M��ࡻ����$��QN���ؔ�96�������7��o^������x0��>S������©�v��� ������î��M��~񫻎������Ѱ����-|���Lɻ�ӻM�ۻ+P������߻{�ٻV3ջ@�һ�ӻ}׻^޻�经��-����� ��  �  ���<0��<P�<h��<���<
��<���<+�<�X�<H[�<O�<nO�<�o�<��<�<R��<��<���<r��<1n�<b1�<���<-�<��<5��<��<��<?)�<�)�<ԧ�<���<��<[��<��<�3�<��<��<���<r��<,d�<�+�<m�<p2�<�h�<���<���<���<�!�<���<���<���<%�<�0�< p�<���<jR�<��<3��<�Z�<8@�<"6�<"�<V��<�b�<݃�<z>�<y��<x��<<��<���<BR�<C�<t9�<��<��<l��<g��<ln�<ro�<���<�d�<S�<�د<SO�<�Q�<>ǩ<��<�I�<`�<�*�<��<���<��<�:�<�\�<щ�<D͑<�$�<@��<s�<ܿ�<֚�<|��<◁<;<=�z<
�u<
p<�j<5�c< �]<u|X<+�S<�4P<�>M<�J<��G<trD<)�?<�f:<p�3<'�,<9�%<�<[�<� <��<�N<0<�
<N><+�<� <i��;Z��;G��;���;ky�;��;[F�;��;Tc�;�X�;@�;�߈;*��;&p;`
];�G;�/;ۇ;ȱ�:u�:��:��s:D�::v�:���9	m9c6�7��m�����f�e&���ͺ���������5��!�r��Y7����8 ��j�jV�K"�K�(��^.���2��_6�+	9�:�:��;���;�b�:�5:���:�D�<�VRA��H��R���]��h�1eq�O�v��|x�=Kv�͋q��Cl�w�h��eh��l�u�0L������|��1ݐ��H��t�6����Đ�&ڎ�ƍ�<���}����8���ŕ�a���k����%�����m���t਻�������;㬻?���rO���¯�o@��T��a��DM����ǻ��ͻb�һ��ջ�ֻ��ջ��ӻ�һ{gѻU�һJֻb�ۻ�%�������!��  �  W��<+h�<��<��<���<0�<3O�<�o�<��<o	�<��<�K�<b
�<���<�1�<�t�<ʍ�<ܚ�<%��<� �<Yv�<��<���<�o�<� �<	f�<!��<��<'�<qP�<���<Gs�<�<�<��<	��<�Q�<���<���<���<�7�<5��<<�<&��<���<���<bA�<!��<��<Vk�<I��<�<�<���<H��<^��<@��<g�<��<]c�<ܟ�<4��<' �<Y��<��<���</c�<F��<z0�<4�<N��<��<��<���<O�<p��<���<�<�<�9�<��<�=�<Bm�<ޘ�<��<�\�<��<��<߫<vϩ<|��<�O�<�ܢ<^�<��<��<)@�<Q�<��<`��<�D�<D��<���<�ׇ<��<�^�<��<��{<`�w<@�s<:p<�l<1�g<"�b< 0^<XxY<�T<}�P<�aL<<.H<g�C<��><~�9<��3<�/.<ʢ(<�}#<��<��<��<*<2<<<b�<V�<�F�;���;P��;��;T��;�
�;���;�;�,�;���;��;��;d��;}jt;Jbc;eS;8�C;�-3;�d!;FF;c��:���:���:0��:.�<:5��9ϣr9-���񑹜���[��p��i���V�ɺQ|޺���I����m�3	�h������M��U#��(�;+��\,��,�F�,��-��-0�cd4���9��>��yC�ȱF�,�H��vI�iJ�&K��\M�Q�kV��T[�9S`�xXd�g�|vh��4i��j�g6l�{p�ŷu��I|�_g��H<���f���釻n�������\?��h$���ŏ��蒻U,���2������$t��s����{��L���@(������f��'Ы��m��ދ������ὶ�i��^t������n���r��,�û�fǻO�ʻ0ͻvϻ�\лWhѻa�һ��Ի��׻|ۻ��޻_�����63��  �  �|�<l��<���<sp�<���<�4�<ֹ�<ʘ�<���<��<��<���<o��<��<���<���<�Z�<G��<H�<!��<���<�A�<�H�<e��<��<Ms�<s��<
N�<��<���<��<�<�#�<Y^�<���<�2�<2��<�n�<EA�<�/�<�!�<���<���<���<+	�<���<�R�<��<u��<���<֤�<���<p�<�#�<��<D��<px�<h��<�1�<��<�)�<`��<�B�<���< �<yT�<ٌ�<!��<2	�<��<f��<��<���<��<֎�<�J�<=�<b��<'c�<%�<��<��<��<E��<�]�<�ì<��<���<i��<�_�<%��<G	�<~�<�j�<�	�<]��<��<�<�<�Ɗ<:7�<���<r>�<:�z<�v<T�r<��o<�m<<�k<��h<�e<��a<��\<��W<<R<�L<� G<��A<N�<<Ά7<ȯ2<{-.<�*<L&<� "<o�<�y<�m<a�<��<Ǘ<7g�;���;R��;ѿ�;T��;��;{��;	��;�Q�;���; 4�;aÕ;�{�;�t;�_;a�M;9T@;z�5;��,;�s";�;��;���:O.�:ʞ�:{1R:z6�9��#9J���aչ��+�O9e�.ꊺ�0���ذ�ߤ��VdӺÐ�o��������a(���2�h�9�>�<�=;��l6��0���+���)�Nd,�h3�#�<��^H��
S�l[��2_�bf_��[\�*YW�)R��GN���L�fcN��FR��X�/�^���e�j�k�E�p�u��x���{���}� �~������)〻�ւ�G��y���._��/���s���[���d��9i��瘤������w���.��>�����lt���4��_=�������»y�»����I���}���㽻���̕��˴û,�ǻ��˻=�ϻuӻ-�ֻ�-ٻMۻ$iݻt�޻��߻�g�d��  �  �!�<��<�d�<2�<Z��<F�<�A�<��<�v�<h��<���<O,�< K�<���<��<�r�<5��<["�<8��<��<�"�<`��</��<���<]#�<�h�<�R�<K��<�p�<j��<�c�<g��<1n�<J&�<�0�<ȗ�<�\�<{�<{��<�X�<J��<w��<0�<,�<>a�<9�<���<]��<c"�<zH�<O�<�$�<���<��<$0�<ΰ�<cT�<d�<m$�<���<���<���<2��<B\�<~��<l��<���<���<��<>��<�b�<���<��<�d�<(��<���<LP�<��<p�<�D�<�<�)�<�m�<R�<C��<9��<�ۨ<8Ӥ<���<��</͙<�e�<�Е<4�<O[�<ܶ�<���<��<�Ӎ<3.�<��<���<�z<�s<q�n<%�k<{j<�]i<M�h<�h<�*f<��b<�h^<>�X<WR<�K<_�D<3�><vK9<�v4<C[0<�,<g�)<z�&<�f#<�+<!�<h�<@><Nd<�R�;m�;0 �;r��;���;�9�;\G�;�Y�;���;�%�;���;4C�;��;��|;�];-cC;�01;�&;�W ;��;I�;��;V�
;��:���:���:UP:�.�9��7Gʥ�M���EV��߀�k7��곛��񦺍c��ϵɺ���h����� .���@��9O�9�V��1W�3�P��E�T~9�3�/�'0+��p-�S�6�OE���V�dh�B@u��1|�x1|�"v� �k�"K_��ET�F�L�n<J�u�L�r?S�Y]��*h���r��{��쀻����䂻�ꁻ���ڑ|��z��3|����b���2g��Ǘ��j��|੻�读`���u	��7o��u5��s ��ޠ�֟��<죻򎪻r���������ƻ�iͻ��л��л�ͻ��Ȼr�û�ȿ�J���%������L�ŻA�˻��ѻ��׻<_ܻt�߻vộ�ỉ�;�߻{�޻{�޻�  �  9��<F��<}?�<I�<��<���<6{�<[	�<���<E��<}d�<r�<�7�<1�<��<C��<�T�<7>�<X�<�8�<�_�<��<�3�<ʡ�<���<���<�T�<L@�<O�<2��<��<�C�<`Y�<���<qt�<���<s��<6�<p�<��<���<y��<��<�[�<P��<��</��<�:�<�G�<�j�< ��<6-�<J�<`��<DG�<l�<5��<�:�<��<���<���<�.�<��<bw�<�9�<]��<��<�-�<�&�<s2�<�:�<OR�<���<K��<"D�<�,�<4s�<�0�<ji�<��<��<dµ<c>�<s �<�>�<،�<%�<�R�<ɉ�<nA�<�ٕ<�<2c�<�#�<sY�<-k�<�ˑ<��<�5�<�.�<:V�<^~<��t<|�l<�)g<" d<�Ec<j�c<ye<V�e<�e<=�b<[J^<$dX<dSQ<x�I<,=B<�q;<��5<�1<z-<L�*<��(<-M&<K%#<�<b�<�-<�W<���;���;�:�;^w�;2�;�9�;�V�;s�;�+�;�~�;|;�;�;���;]��;~;h;�$C;��%;Ѥ;�	;�/;��	;�g;ۀ;�;���:w�:9�:XN=:hɋ9M�%���LS����IV���Ŝ��ġ����s���vRͺ�`�	@�.*��=E���\���m�`�u�K}s��\h��pW��^E� �6���/�q�1��l=���P�rh��,�����y��!���2L���Ɓ��eq��`��"S��L��KM��LT�) `�`wn�Ѧ|�1+�����o�����Zo���セ����{�t}������J�������������舸��|�����_���7Z��4��87��~��Ǣ��m���5��22ǻ�.ӻ%�ۻ�R໤�߻�^ۻEԻ=�˻��Ļ����[/���dƻF�ͻ�ջW$ݻo㻺��#=�-z�=����;{߻�޻�  �  �X�<V��<���<WE�<�g�<���<��<��<���<���<��<���<%�<4e�<�]�<s��<��<oo�<^��<�I�<1�<A�<��<���<Z"�<���<l
�<rk�<\��<i	�<�}�<k�<�7�<�E�<#��<�2�<�A�<U��<��<6�<�<�<&;�<�K�<b�<��<�,�<N�<f��<��<8��<*��<7�<�<�D�<�_�<�<�B�<I�<M��<t�<U�<?Z�<=�<���<��<�<�<Rx�<A��<an�<��<I��<W��<B��<-��<~��<Cǻ<؈�<H�<2Ѷ<���<��<)��<|��<ce�<�C�<~H�<�ڟ<!��<��<Z�<G,�<�]�<g��<'s�<��<��<Hi�<&r�<E�<Ѿ�<kz<�3o<�`f<�\`<�`]<[]<"�^<��`<h�b<0#c<}Xa<`O]<IW<��O<2�G<_�?<�Z8<�a2<��-<�*<��(<'<[%<�"<�n<v�<9I<A<�V�;�X�;��;?��;>3�;r�;�G�;S��;���;	q�;��;Q�;��;���;k�U;]3,;/;%�:Ë�:�P�:��:5��:ܕ;
A;�d�:q'�:�:��#:�9n`��Z�9�����L��ʧ�ݬ���r���������F�׺�s �����;��_[���v�W���ri���3���}���g�i;Q�~�>���5���7�gE�%\��x��񉻙딻@��Z��|M��:%��-Ձ��pm�\��pR�jyQ��{X���e�$�u�;�����
s������r������Tf��W�� �������Յ�Q6��7��S0��tй���ŻTLͻ6:ϻW~˻27û�����u��	{��ď�����p��8����л�B޻X�軫�0��=���޻�4Ի�ʻ��û�s���1û��Ȼ��лj�ٻ�g�,黓F��l�컔Q�Q����O���  �  ��<���<��<���<X��</��<j��<�<�<�R�<F��<��<6��<'1�<-��<���<�1�<�!�<$�<���<oH�<��<���<���<���<-Q�<x\�<k��<���<�+�<g��<���<��<S]�<HF�<���<5�<�4�<��<�J�<ە�<dy�<ې�<��<�b�<i�<-�<!,�<���<�y�<ư�<ހ�< ��<���<���< }�<���<�v�<ʁ�<#:�<�7�<�9�<���<��<:��<ة�<���<��<�#�<��<0��<��<�,�<�D�<���<��<K��<���<�c�<�ܶ<d�<�8�<um�<��<�<��<�5�<�ڣ<g�<oh�<_��<��<?ߍ<�M�<A�<��<��<1�<َ<�Ջ<?D�<_��<��v<wqk<�b<��[<˳X<r�X<N�Z<��]<dx`<�ya<� `<AE\<%1V<؁N<�	F<	�=<%26<�0<+�+<?�(<��&<+�%<�#<l� <�.<�*<?�< *<���;Ë�;�)�;00�;+X�;W-�;���;^��;�9�;���;���;uP�;PP�;OOy;A�H;%;æ�:��:9��:�ӽ:!��:�#�:���:t��:>��:�=�:!�:[9:��8j�[�[�����������8������������ź���ܑ��%�D�H��Ik��C����ڬ��0��������s�,�Y��*E�cJ:��5<��K�Fsd� �������Q���<��_֤��g���I��
�����w��c��W���U�ٽ\��{j���{��؆��3���䒻�^��𲒻����3C��Cs���ၻP�������[J���ʡ��K���6»+	ϻ��ֻ�Rػ�ӻh
ʻw�aa���E���ϧ�7����d���YŻ�1ֻr��6��2q������V�����Q{ڻGQϻIXǻ/�ûMŻ�ʻ8Iӻ�ܻ97滀t��������컍��A�.��  �  3��<1z�<�B�<-�<���<6��<p��<�f�<���<�6�<��<��<��<ׄ�<��<���<���<(��<�W�<���<��<P�<s��<B��<]��<���<	��<�]�<w��<�K�<ĭ�<zr�<�<���<�d�<���<6��<1��<���<!V�<�@�<�W�<O�<s�<ţ�<a��<�q�<��<���<���<ѿ�<A�<�:�<���<22�<��<#>�<"9�<���<���<	��<�<�<�6�<��<X��<��<���<���<��<�p�< ��<���<�<�p�<	��<,�<7�<Z��<�{�<��<+�<�,�<1�<���<mT�<�ͨ<�Q�<&a�<���<���<?�<��<ג�<�L�<қ�<��<u�<���<}��<��<{*�<��u<�j<L�`<Z<9W<�W<ecY<V�\<��_<��`<͡_<��[<��U<1�M<�nE<9�<<?l5<QQ/<��*<�(<�U&<�%<no#<H� <��<;�<�<� <��;�^�;���;յ;�5�;�n�;b��;�<�;H�;��;��;@T�;��;�u;��C;�;��:T��:�ث:��:�:���:wa�:�K�:[�:��:މ�:$�:/���������g�=M��u���A]����O湺���A4ɺ�溣]
��)�?�M��q��~���p��~������k�����w�-#]�xG�%<���=�;^M��g��ƃ�T����J��9���7������?��\����{��f�@Z���W��^�nql��E~�]-��n����y��-�j)���ۏ��^���f��:���0샻�牻ޔ��⣻_鴻mBŻ�Yһ�'ڻ��ۻ�ֻ�x̻�߿�?ӳ��U������������ǻ�gػ�� ������� S�����S�_�ܻ
ѻ(�ȻP�Ļ�.ƻ��˻QԻB4޻��/���U�bJ���"�7����}�����  �  ��<���<��<���<X��</��<j��<�<�<�R�<F��<��<6��<'1�<-��<���<�1�<�!�<$�<���<oH�<��<���<���<���<-Q�<x\�<k��<���<�+�<g��<���<��<S]�<HF�<���<5�<�4�<��<�J�<ە�<dy�<ې�<��<�b�<i�<-�<!,�<���<�y�<ư�<ހ�< ��<���<���< }�<���<�v�<ʁ�<#:�<�7�<�9�<���<��<:��<ة�<���<��<�#�<��<1��<��<�,�<�D�<���<��<M��<���<�c�<ݶ<h�<�8�<{m�<��<�<&��<�5�<�ڣ<o�<wh�<g��<��<Eߍ<�M�<F�<��<��<1�<َ<�Ջ<=D�<\��<��v<mqk<�b<��[<��X<b�X<?�Z<��]<Tx`<�ya<� `<5E\<1V<ρN<�	F<�=<"26<�0<-�+<C�(<��&<3�%<!�#<x� <�.<�*<N�<*<ǰ�;��;�)�;L0�;DX�;m-�;���;l��;�9�;���;���;pP�;FP�;3Oy;�H;�~;_��:���:���:1ӽ:���:f#�:y��:���:ɰ�:=�:� �:�8:��8!k�˴[���������K������ǳ����ź���ݑ��%�D�H��Ik��C����ڬ��0������ߟs�,�Y��*E�cJ:��5<��K�Fsd� �������Q���<��_֤��g���I��
�����w��c��W���U�ٽ\��{j���{��؆��3���䒻�^��𲒻����3C��Cs���ၻP�������[J���ʡ��K���6»+	ϻ��ֻ�Rػ�ӻh
ʻw�aa���E���ϧ�7����d���YŻ�1ֻr��6��2q������V�����Q{ڻGQϻIXǻ/�ûMŻ�ʻ8Iӻ�ܻ97滀t��������컍��A�.��  �  �X�<V��<���<WE�<�g�<���<��<��<���<���<��<���<%�<4e�<�]�<s��<��<oo�<^��<�I�<1�<A�<��<���<Z"�<���<l
�<rk�<\��<i	�<�}�<k�<�7�<�E�<#��<�2�<�A�<U��<��<6�<�<�<&;�<�K�<b�<��<�,�<N�<f��<��<8��<*��<7�<�<�D�<�_�<�<�B�<I�<M��<t�<U�<?Z�<=�<���<��<�<�<Sx�<B��<bn�<��<J��<Y��<D��<1��<���<Hǻ<ވ�<P�<;Ѷ<���<��<6��<���<re�<�C�<�H�<�ڟ<0��<��< Z�<S,�<�]�<p��<.s�<��<��<Hi�<%r�<A�<˾�<[z<�3o<�`f<�\`<m`]<>]<�^<|�`<J�b<#c<bXa<HO]<�HW<��O<$�G<U�?<�Z8<�a2<��-<��*<Ȥ(<,'<o%<�"<�n<��<VI<4A<�V�;�X�;D��;t��;n3�;��;�G�;n��;���;q�;��;H�;��;���;%�U;
3,;�;P�:ފ�:P�:��:=��:b�;�@;�c�:�&�:@�:R�#:S�9ub��2�9�g���M��9ʧ�����r��'�������M�׺�s �����;��_[���v�W���ri���3���}���g�h;Q�~�>���5���7�gE�%\��x��񉻙딻@��Z��|M��:%��-Ձ��pm�\��pR�jyQ��{X���e�$�u�;�����
s������r������Tf��W�� �������Յ�Q6��7��S0��tй���ŻTLͻ6:ϻW~˻27û�����u��	{��ď�����p��8����л�B޻X�軫�0��=���޻�4Ի�ʻ��û�s���1û��Ȼ��лj�ٻ�g�,黓F��l�컔Q�Q����O���  �  9��<F��<}?�<I�<��<���<6{�<[	�<���<E��<}d�<r�<�7�<1�<��<C��<�T�<7>�<X�<�8�<�_�<��<�3�<ʡ�<���<���<�T�<L@�<O�<2��<��<�C�<`Y�<���<qt�<���<s��<6�<p�<��<���<y��<��<�[�<P��<��</��<�:�<�G�<�j�< ��<6-�<J�<`��<DG�<l�<5��<�:�<��<���<���<�.�<��<bw�<�9�<]��<��<�-�<�&�<t2�<�:�<QR�<���<O��<&D�<�,�<<s�<�0�<ui�<��<��<tµ<v>�<� �<�>�<팫<!%�<�R�<މ�<�A�<�ٕ<Ԍ�<Bc�<$�<~Y�<5k�<�ˑ<��<�5�<�.�<2V�<�]~<��t<\�l<e)g<�d<bEc<@�c<Oe<+�e<�e<�b<8J^<dX<KSQ<d�I<=B<~q;<��5<�1<%z-<^�*<�(<IM&<k%#<&�<��<�-<(X< ��;���;3;�;�w�;I2�;�9�;�V�;*s�;�+�;�~�;|;�;��;���;8��;;h;8$C;)�%;:�;	;#/;��	;g;.�;e�;���:�u�:( �:oL=:Ƌ9�%�O���LS�)���V���Ŝ��ġ�9��������Rͺ�`�@�/*��=E���\���m�_�u�K}s��\h��pW��^E��6���/�p�1��l=���P�rh��,�����y��!���2L���Ɓ��eq��`��"S��L��KM��LT�) `�`wn�Ѧ|�1+�����o�����Zo���セ����{�t}������J�������������舸��|�����_���7Z��4��87��~��Ǣ��m���5��22ǻ�.ӻ%�ۻ�R໤�߻�^ۻEԻ=�˻��Ļ����[/���dƻF�ͻ�ջW$ݻo㻺��#=�-z�=����;{߻�޻�  �  �!�<��<�d�<2�<Z��<F�<�A�<��<�v�<h��<���<O,�< K�<���<��<�r�<5��<["�<8��<��<�"�<`��</��<���<]#�<�h�<�R�<K��<�p�<j��<�c�<g��<1n�<J&�<�0�<ȗ�<�\�<{�<{��<�X�<J��<w��<0�<,�<>a�<9�<���<]��<c"�<zH�<O�<�$�<���<��<$0�<ΰ�<cT�<d�<m$�<���<���<���<2��<B\�<~��<l��<���<���<��<?��<�b�<��<��<�d�<.��<���<UP�<��<}�<E�<��<�)�<�m�<4R�<\��<S��<ܨ<SӤ<���<(��<F͙<�e�<�Е<D�<[[�<嶓<���<��<�Ӎ<,.�<��<狁<��z<��s<E�n<��k<Hj<O]i<�h<�h<�*f<��b<�h^<�X<�VR<�K<N�D<)�><tK9<�v4<Q[0<1�,<��)<��&<g#<�+<Q�<��<t><�d<BS�;qm�;� �;���; ��;:�;�G�;Z�;���;�%�;��;C�;��;/�|;4];�bC;A01;�&;�V ;!�;q�;!�;��
;���:?��:6��:�P:�*�9�ـ74ͥ�}���FV��߀��7������񦺣c��ݵɺ���h����� .���@��9O�9�V��1W�2�P��E�S~9�3�/�&0+��p-�S�6�OE���V�dh�B@u��1|�x1|�"v� �k�"K_��ET�F�L�n<J�u�L�r?S�Y]��*h���r��{��쀻����䂻�ꁻ���ڑ|��z��3|����b���2g��Ǘ��j��|੻�读`���u	��7o��u5��s ��ޠ�֟��<죻򎪻r���������ƻ�iͻ��л��л�ͻ��Ȼr�û�ȿ�J���%������L�ŻA�˻��ѻ��׻<_ܻt�߻vộ�ỉ�;�߻{�޻{�޻�  �  �|�<l��<���<sp�<���<�4�<ֹ�<ʘ�<���<��<��<���<o��<��<���<���<�Z�<G��<H�<!��<���<�A�<�H�<e��<��<Ms�<s��<
N�<��<���<��<�<�#�<Y^�<���<�2�<2��<�n�<EA�<�/�<�!�<���<���<���<+	�<���<�R�<��<u��<���<֤�<���<p�<�#�<��<D��<px�<h��<�1�<��<�)�<`��<�B�<���< �<yT�<ڌ�<"��<3	�<��<h��<��<���<��<܎�<�J�<H�<n��<6c�<0%�<��<��<��<`��<�]�<�ì<��<���<���<�_�<?��<^	�<��<�j�<�	�<g��<��<�<�<�Ɗ</7�<���<_>�<�z<�v<�r<O�o<��m<�k<k�h<��e<{�a<��\<w�W<�;R<֡L<� G<��A<L�<<Ն7<ׯ2<�-.<*<s&<� "<��<�y<.n<��<�< �<�g�;��;���;"��;���;#��;���;��;�Q�;���;�3�;.Õ;_{�;s�t;_;��M;\S@;��5;��,;�r";�;��;���:�,�:U��:�.R:�1�9�#9Ў�odչ��+�:e�{ꊺ�0���ذ�����fdӺ͐�u��������a(���2�g�9�>�<�=;��l6��0���+���)�Md,�h3�#�<��^H��
S�l[��2_�bf_��[\�*YW�)R��GN���L�fcN��FR��X�/�^���e�j�k�E�p�u��x���{���}� �~������)〻�ւ�G��y���._��/���s���[���d��9i��瘤������w���.��>�����lt���4��_=�������»y�»����I���}���㽻���̕��˴û,�ǻ��˻=�ϻuӻ-�ֻ�-ٻMۻ$iݻt�޻��߻�g�d��  �  W��<+h�<��<��<���<0�<3O�<�o�<��<o	�<��<�K�<b
�<���<�1�<�t�<ʍ�<ܚ�<%��<� �<Yv�<��<���<�o�<� �<	f�<!��<��<'�<qP�<���<Gs�<�<�<��<	��<�Q�<���<���<���<�7�<5��<<�<&��<���<���<bA�<!��<��<Vk�<I��<�<�<���<H��<^��<@��<g�<��<]c�<ܟ�<4��<' �<Y��<��<���</c�<G��<z0�<4�<O��<���<��<���<S�<u��<���<�<�<:�<��<�=�<Tm�<�<��<�\�<��<��<%߫<�ϩ<���<�O�<ݢ<7^�<��<#��<;@�<_�<��<f��<�D�<A��<���<�ׇ<��<�^�<��<i�{<(�w<�s<�p<Rl<��g<��b<�/^<'xY<��T<Y�P<�aL<(.H<\�C<��><��9<��3<�/.<�(<~#<��<��<(�<d<o<<J<��<��<G�;B��;���;��;���;�
�;���;�;�,�;`��;g�;��;��;�it;vac;0dS;G�C;�,3;�c!;PE;���:9��:9��:���:z�<:z��9��r99G����������[�q������~�ɺl|޺���T����m�3	�i������M��U#��(�:+��\,��,�F�,��-��-0�cd4���9��>��yC�ȱF�,�H��vI�iJ�&K��\M�Q�kV��T[�9S`�xXd�g�|vh��4i��j�g6l�{p�ŷu��I|�_g��H<���f���釻n�������\?��h$���ŏ��蒻U,���2������$t��s����{��L���@(������f��'Ы��m��ދ������ὶ�i��^t������n���r��,�û�fǻO�ʻ0ͻvϻ�\лWhѻa�һ��Ի��׻|ۻ��޻_�����63��  �  ���<0��<P�<h��<���<
��<���<+�<�X�<H[�<O�<nO�<�o�<��<�<R��<��<���<r��<1n�<b1�<���<-�<��<5��<��<��<?)�<�)�<ԧ�<���<��<[��<��<�3�<��<��<���<r��<,d�<�+�<m�<p2�<�h�<���<���<���<�!�<���<���<���<%�<�0�< p�<���<jR�<��<2��<�Z�<8@�<"6�<"�<V��<�b�<݃�<z>�<y��<y��<<��<���<CR�<F�<w9�<��<��<u��<q��<yn�<�o�<���<�d�<j�<ٯ<nO�<�Q�<[ǩ<#��<J�<}�<�*�<��<��<��<;�<�\�<ۉ�<J͑<�$�<=��<k�<ѿ�<ƚ�<i��<̗�<
<�z<ёu<�p<�j<��c<��]<A|X<��S<�4P<�>M<��J<��G<irD<'�?<�f:<��3<?�,<Y�%<�<��<� <*�<�N<J0<;�
<�><b�<$� <Š�;���;���;ǈ�;�y�;���;\F�;��;1c�;jX�;��;P߈;κ�;8%p;�	];/�G;+�/;�;��:��:;�:f�s:Y�::٥:��95m9"�7.�m�����f��&��E�ͺ�� ����6��!�t��Z7����7 ��j�jV�K"�K�(��^.���2��_6�*	9�:�:� �;���;�a�:�5:���:�D�<�VRA��H��R���]��h�1eq�O�v��|x�=Kv�͋q��Cl�w�h��eh��l�u�0L������|��1ݐ��H��t�6����Đ�&ڎ�ƍ�<���}����8���ŕ�a���k����%�����m���t਻�������;㬻?���rO���¯�o@��T��a��DM����ǻ��ͻb�һ��ջ�ֻ��ջ��ӻ�һ{gѻU�һJֻb�ۻ�%�������!��  �  {D�<�f�<d7�<Rm�<���<N��<3�<���<�	�<>��<HD�<>��<K�<�1�<s�<��<]	�<uI�<��<}��<��<�^�<>�<���<�I�<m��<.�<���<ā�<?�<@��<���<�^�<��<�<���<���<���<<�<z��<���<N��<��<��<'C�<d��<��<��<�o�<�:�<�y�<�Q�<���<7��<���<��<T�<A�<8��<���<�w�<r��<p��<���<��<�{�<��<�*�<��<�T�<���<���<���<��<���<34�<%��<d^�<��<��<-��<�D�<씬<u��<nا<O��<"4�<�ܥ<�W�<uY�<ڻ�<y�<;��<gh�<���<	��<�g�<%��<o�<ۈ<J
�<*v�<��<�8�<�&�<K-{<y�t<��m<��e<g^<=W<YQ<��L<DJ<єH<�G<�VF<��C<�?<�9<��2<Z�)<�@!<K7<.�<��<�<�	<�	<�<$�<�w<��<�m�;���;���;:��;���;��;���;�	�;h�;s�;r�;���;�3�;Et;��];C�B;E+$;E�;]��:���:+�D:�:��9܄�9W o9��9k��Z8����c*��g�����	���=#�!^+���+���&��0��������������^�J��1�*���4�/G=���B��E��E�Q�B��>�g�8��W5��4��8�+�A�O�T%`��?r�g?���$���쉻�=��X�������Jt���k�Wji�^�m�iCy�j�,���݀���M��ࡻ����$��QN���ؔ�96�������7��o^������x0��>S������©�v��� ������î��M��~񫻎������Ѱ����-|���Lɻ�ӻM�ۻ+P������߻{�ٻV3ջ@�һ�ӻ}׻^޻�经��-����� ��  �  �]�<6��<��<%��<���<���<���<���</��<i��<u��<I��<���<}�<?��<@i�<x��<�`�<�,�<Y��<���<�&�<���<�>�<U>�<6�<��<���<Ξ�<���<s��<��<V��<���<f�<�&�<c��<F�<�7�<k�<���<v�<8��<:x�<�%�<�N�<�v�<=&�<��<O�<f^�<���<�?�<�|�<� �<���<Џ�<J��<�N�<�6�<��<���<܌�<��<{��<���<8��<+�<���<ށ�<R �<V��<���<��<<y�<�s�<�O�<�ݿ<�*�<3�<tY�<NY�<t�<���<-�<R�<2`�<@ʣ<e�<;��<J��<�p�<Ɔ�<���<�$�<�O�<*Ɏ<���<PG�<�`�<��<΄<d��<�<7�<`+z<��r<;j<�`<q�W<�O<�EI<EE<UyC<�[C<D�C<�D<R�B<{�><µ8<�a0<��&<�N<7�<)T<29<��<'<��<�<=x<k|<��<u$�;L��;D�;@��;���;2��;�6�;Y+�;�O�;��;Y��;��;O��;��q;u:X;�08;�I;8�:t�:�#:��9�m8uGʷP�[�К�7�[�7w3���J��|�4�&֘�ߺN��s�.��B�R�J�qTI�z�?�%�1��"���������S�z�"��M0�!>�T�I�2Q���S�M2R�qL��<D�?�;��U6�c�5��M;��H��4[��r��K��v���`����B��a��s搻�K��S��r���m�l�r��\���������X�������H^��^�����*ॻ~a��P���A���9�������9��j���`Ģ�X<���G���?��o絻V��#����˯�����󫻡������%-����ƻ�ӻ�"�7l�]������Gq黣J�Y�ٻLaջ�-ջ�ٻ���y������Q���  �  ���<�C�<���<63�<
��<T!�<���<d�<*u�<���<���<ך�<��<)��<�
�<���<Sf�<�[�<am�<�4�<~R�<���<���<l��<D �<�P�<b��<�f�<�1�<�o�<� �<�w�<z.�<Mo�<���<�s�<|��<*��<�O�<$��<T��<Z��<�9�<�+�<�9�<���<ް�<���<L�<��<���<QW�<t[�<O�<ґ�<�h�<���<�<�<l�<:L�<�r�<�$�<=	�<���<���<`Q�<_`�<�T�<���<�<���<x��<�m�<K��<p"�<���<���<V1�<�4�< �<�O�<���<E�<a��<���<�,�<���<��<���<ҷ�<��<��<��<]M�<�-�<�<�J�<�"�<ҳ�<d��<�ф<��<]��<֏�<��~<�fx<2p<�=f<��[<ZtQ<�H<:UB<W�><ӣ=<?�><Ld@<E�A<`�@<��=<�%7<.<5#<	�<�A<�<~��;7��;� �;;��;�<K�<��<�� <*�;_p�;��;�}�;:r�;\6�;j��;I�;3�;�Ҏ;Ae�;��;�V�;WOl;Y�O;��+;��;k>�:�E9:esQ9NQ"�.���侹2���6�dL���@�ׅ׹��R� ծ�����&���F��]��f���c�aW���D�O�0��� �b���Q��{�n�'��~7���G��U�X�]�u�`���]��#V���K��VA��|:���9�g2A��5Q���h�U����Ɛ�b���tr��㿦�(W��*#���/���@���.z��s���x��z���%����C>��'/��g��3��鹻�谻����曻Rh���鐻����xb���ݝ������R���I��ز���-��Nົ�t������n��w��������ot��r<λ}�ݻ�:�W�����������r���-��Ld���޻`�ػ��׻Aݻ5�˾��_�� �	�*~��  �  i��<k��<ŧ�<�R�<�S�<��<���<Wx�<%��<Wg�<�5�<M��<B��<���<���<��<}t�<���<���<���<0��<��<��<҈�<V��<�]�<U��<+
�<-��<"D�<}�<��<��<��<�<��<��<���<���<H��<���<�d�<Z��<��<�#�<+�<�Q�<���<��<��<HU�<K��<U��<|n�<V��<�N�<���<�5�<'6�<���<���<��<��<5�<p��<%�<ڭ�<�L�<�}�<f��<g�<�y�<[��<K�<�"�<B��<�"�<N��<�t�<Q��<Q߮<^�<~�<nO�<�^�<���<X��<��<SN�<�١<PF�<�s�<�~�<���<�j�<�"�<�=�<N�<��<l��<���<�=�<<f�<$�<e�}<A�v<�m<oHc<�W<""M<�D<̓=<�&:<٦9<�O;<��=<N�?<T�?<�k<<��5<�[,<P� <��<�f	<� <Az�;��;vf�;	�;@�;q� <L(<,��;&�;�.�;�M�;]&�;�|�;v̨;��;І�;���;���;w��;ݸ�;q*|;vg;��H;#�!;���:��:=m�9�������z�������������Th��׈�[3��CGj��'���
�K4�XkW�Avo��y�}v��+h���R�� <�T�(�0��(����n�,�Q=���N�kF]�еf���i�}&f��O]�i�Q�c2F�B�>�34>��F���X�|s��m��5����٥��ﭻ��G����2��>Ǖ��d��h	���x��G}����󘕻糧A�������AUȻ�ȻK�»_ٸ�2����ߠ�T������jۓ�I���xe��ѩ��	�����;)��f����־��Ժ��㵻�����K?���$����Ļ�Իz�������� �*�Qs����ԁ���|����cۻ�+ڻH�߻p����`��-y�����  �  g8�<
A�<��<�;�<]r�<�v�<�_�<��<`��<��<P�<�P�<eE�<���<��<���<H-�<��<-��<>��<���<���<,��<QU�<��<���<�z�<�<�<J��<��<��<�h�<[O�<?F�<g,�<�Q�<���<�k�<Ƹ<#�<�/�<4��<�<��<Ɇ�<��<	��<���<���<J^�<ig�<
��<h��<���<��<���<�s�<���<}��<}��<^��<�~�<e��<�Y�<��<�,�<���<_\�<VX�<hq�<�0�<���<K�<v��<��<�Ī<@�<�D�<Y��<䱚<é�<�݈<[��<��y<�.v<�Ax<.�~<ƿ�<�X�<�<<S�<y��<�%�<:�<�n�<�U�<�|<�8v<�.q<�m<�k<u�h<�ie<�(`<�W<jGL<�V=<�(,<�s<�1
<_��;q��;P��;6��;���;�<��<��<< <C8<�D�;���;��;��;��a;|�E;�QA;�R;R�q;R�;TA�;��;�ɲ;ٱ;��;]�;?\�;o?z;�r\;�D;�32;��%;�3;n�;[�;Xx�:�:1��9�@�ﺨ�>���}�����̣�縥�W����b�����f���^���k�����U|����»]��1������
�����i��5��k�ϻb���x��D�����Ϙ��J��.M��.ϫ�41��Bo��t}��CO��5~�����J���X��I����˻}Y廓�������q% �� ��.�P��K�@���-��0eܻ�{߻{��Wp�*'�Uj���'��-�O�,�K�&��������P�����ڻ:Iٻ�hݻ�们����󻺒����� Y��8 �����e��������A���/!��0�ޘ=���G�<�L�2L��F�!<�wj0���%���@��xf ��)��[6��D�WJQ��XZ��  �  ���<��<?,�<�]�<^W�<��<���<���<�*�<���<C�<��<ȓ�<2��<��<���<�w�<H�<6��<{��<^��<��<�7�<��<���<�<�׵<���<M$�<Uc�<��<�i�<�<~��<���<���<�1�<'�<\��<�
�<�}�<S�<f�<x�<̯<���<�ǻ<s~�<���<���<t��<N�<|��<���<}W�<�6�<��<�/�<��<��<���<��<V�<u��<���<��<w��<��<���<K�<���<��<>�<홤<<(^�<��<6Ш<A:�<�v�<韒<��<��<h�|<\y<��z<�<ݶ�<a�<֜�<��<Vَ<�N�<�d�<c��<p��<�}<��v<g�q<cIn<��k<�i<$�e<׋`<"�X<� M<��><.�-<��<��<Z0 <�|�;x�;ͫ�;=�;5Y<8�<6<<�\<@��;$(�;U�;��;�l;�YQ;V�L;K�\;ۄz;Uv�;Ԡ;�­;5�;���;���;
̝;�T�;¾|;e_;�.G;5;7(;�;um;� ;B�:�+�:�2�9��)��ߺ�)5��r�N����䝻01���ޘ��R����x��ya�Z�*Vg��#��փ������d{޻\���0�3�����fN�����J�̻JH��M�LF���e���#���|��@��V��L����ﯻq'��^;��a����c��/���ki���%����Ȼ�7� �� B�k��2�����?��O"���T�[+ڻ�;ݻ5A��� �?1�����$��%*�F�)�f$��z���2��P�sn��ٻs�ػ,�ܻ���α�O�����{��Q�����i��[��k��@���'�m���s�P�-��:��D���I�V_I���C���9��.�^$�oh�I{��=��)(�8�4�gB���N���W��  �  ���<���<4��<�x�<���<r��<���<���<W��<�<�<���<4)�<�a�<!��<��<���<%;�<V��<�[�<wM�<.�<Κ�<qq�<���<j��<p%�<���<gɵ<�@�<�@�<���<d@�<�c�<���<_I�<�^�<���<�3�<E�<L4�<-,�<��<ɇ�<�j�<�M�<q�<3��<��<���<y,�<���<6z�<�5�<���<C4�<�2�<���<��<��<מ�<�3�<��<���<v��<���<E�<Iq�<t�<���< �<M��<r��<ml�<.3�<�Ǫ<��<��<�I�<��<��<X�<QS�<���<�[�<ƚ�<�G�<G̃<�T�<���<qߍ<4h�<|M�<s��<�Ê<,�<X�<p]<�x<��s<��o<��l<�j<A�f<ea<%�Y<8CO<n�A<��2<��"<�<@<Ɗ <�i�;D�;��<*A<��<�I<�<~	<�u�;x��;�Һ;��;z�;�#r;9�l;��y;��;^
�;/��; �;���;VD�;�
�;؋�;�͐;ǩ�;+=g;FuO;z�<;'�.;y�";s;�+;���:���:e(�9��ٹU���f��i(T��*���O��ė�����£��f��R��]M��[���|�?2��������ѻ������I3��o����4���ػe�ûNE���(�������ݔ�ͩ��(���������� �����������Jq������栻�!���H��>����:ûi�ٻ��
^����������|
�p����B뻱�ۻ�&Ի]׻h)以���ߤ�.[��U���!��!��s�a���X	��m���'�yF޻��׻23׻'ۻ��6�����G󻨛��������ﻋT5������g`����P�'�?�3�Y�<���A�~lA��n<�&�3�o�)�Wx ��.�����6\$�S�/��v<�(�G��O��  �  "��<d��<�<���<���<{��<�<��<���<�b�<kE�<���<Jb�<�0�<�h�<��<�)�<*o�<S��<�o�<�i�<�@�<Z��<^?�<���<���<���<��<-?�<��<ň�<�l�<���<EN�<�g�<Rg�<.0�<�$�<0�<�ݺ<Ș�<��<��<��<u:�<�_�<3��<L��<���<݌�<��<��<���<wm�<�L�<�{�<}�<�/�<h��<��<mg�<%�<]��<�j�<G��<i��<"8�<*ή<�)�<��<���<��<a�<	 �<G��<Q�<���<�J�<�Z�<���<�T�<4.�<�B�<�C�<4u�<Z��<�Z�<�؊<(c�<L�<M�<?��<:��<���<#��<R8�<�ـ<N�{<�gv<r<�Xn<��j<�f<C�a<X�Z<�Q<��E<��8<i2+<�g<^�<�<�f	<�
<�<h<�b<~�<<��<�<�X�;;�;�}�;<�;��;4��;���;��;k��;l��;E̶;ܗ�;S��;g��;��;���;�ǅ;�}q;cdZ;��F;��6;�<(;=�;v�;%��: 5�:g�&:�Y���{�P��j�(��P�A8j�nJs�C�m���]��DK���=�e�;�(iJ��i��<���>���羻�@ԻJ-�+�TB��cػ�ɻ
g�����\���o���@���ە�����c��Ꞣ�;���񽦻���!'��W���R��ѕ��o𤻊.������ϻ@��6o����� 	�� 
���� �2�r)߻oһ��˻�λ*ڻ-�n ��z
�s�������,����
��4�<��%D��kۻ��ֻc�ֻ�ڻdl߻W&廔2�D������.�����)��;�������^
�����z�'�)��F1��5�l�5��1���*�U�"������4w�h��q����(�O�3�]=��D��  �  ٩�<�<���<.(�<-��<��<���<j��<w�<��<"�<��<�-�<�V�<r��<�.�<���<ۚ�<+P�<Z��<���<��<���<*�<K�<�Y�<w��<�F�<*�<�x�<�T�<�1�<�[�<��<1��<�u�<2��<3_�<aR�<�:�<pڼ<�Ǻ<�J�<PN�<z�<�P�<AN�<��<���<��<�h�<*�<��<l��<M;�<��<RV�<)(�<��<��< ��<eq�<v\�<9v�< ��<0	�<S��<�ݳ<�@�<h��<|<�<�I�<��<YN�<���<̶�<D�<�N�<K�<�-�<�ݝ<�×<R��<���<�<[��<��<G>�<Ub�<e�<T�<dގ<��<���<Ň<�Ԅ<��<,~<m�x<��s<�o<ݏj<��e<ݍ`<�.Z<�_R<�I<��><�3<�~)<̴ <�M<q�<>I<L�<�w<Vg<9G<�<m8<�M<��;���;c3�;2[�;���;�(�;ͧ;p��;���;#Q�;>��;#C�;�F�;k;�;��;eɔ;:�;�{;�d;8P;~�<;�X*;\;Er;�k�:��:��?:�� 9^"�ze����d�3�2�a>���>��7�yA-��*'��*�1h9�ĩU��"|��㓻�8�� ��>�ƻ\�˻Nʻ�=û;7���/��h#�������I���񖻥җ����@}��Sڞ�����̡��-���
�����v塻'Q������㭻$9���ŻggԻ���.ﻌ��2������'C��޻��ѻL�ǻ��û�;ƻ݆ϻ��ݻGg��.��7#�gW��d�æ��� �Ȇ���I��Ở�ۻ�ٻ�Sٻ��ۻ �޻�����廸�軺�껨F�H�K����"@�Z���"�Gh��������~��w$��'��`(���%�� ���������d�O-��!�y�)�`1�w�6��  �  �7�<��< ��<���<���<���<"��<k��<��<���<��<��<._�<��<~�<���<q��<���<z��<m��<ٹ�<Hh�<8��< ��<��<&.�<��<Zy�<+��<~��<e��<��<���<�g�<�I�<�<��<�A�<tW�<�h�<C��<�W�<ʼ�<��<���<%A�<k��<V��<B��<��<*[�<�z�<��<Ġ�<N��<v�<V�<��<���< �<*J�< d�<�W�<��<F�<G�<,��<#�<�ʵ<*�<4��<�]�<.��<�X�<س<K��<�l�<.گ<�<qJ�<�&�<�)�<�Ҙ<y�<7/�<�ˑ<��<m��<V�<[�<�>�<)��<���<�<q��<4Ƅ<m�<R�<x<z<�at<wXn<�Mh<`b<Ӈ\<I�V<bGP<�jI<�B<�~:<�23<��,<1m'<��#<�,"<8�!<��!<�!< �<�<��<6J<�~< ��;Z8�;<��;���;B��;�W�;2��;լ�;@�;$u�;��;S�;�Ӣ;��;�ؒ;�;�~�;�*l;��U;�>;��%;0�;���:jI�:��:�f+:�j[9�㊹�RC�����;Һ	$����
�)�����E��X������+���D��td�!���.<���^��rm���ұ������`J��~֨��Ƥ�)Ρ�I����-�����������F��;��������b�������{��y^���o��  ����������N_ɻƢѻX�ػmvݻ?�޻r$ܻ�ֻ��ͻ/�Żc����1��I����zƻ�л"�ܻ��Z�sQ��h�������������.軂q仙.��E��8����	�Ȳ�G��0��G軫;����.�)��$���aG �l[��,�-��ba�}��"��1���]�������ǉ��X�A=���6�����e �ȵ%��)��  �  ���<1��<.�<�s�<���<`<�<ǯ�<�N�<�>�<���<9�<�<B��<���<Ֆ�<Օ�<*�<S�<�#�<�Z�<?��<���<z�<���<��<a�<��<�]�<8�<*�<���<vd�<�A�<���<�7�<���<���<Q�<�}�<��<#
�<���<?��<�\�<}��<�{�<�<��<�i�<�Z�<(��<�Y�<�Q�<�W�<5&�<{�<�*�<2�<���<��<;�<=��<���<���<���<;Y�<�<�Һ<B�<��<��<Tk�<S�<��<3�<�ִ<�<��<bW�<��<$��<m��<���<�˚<�<ʙ�<(N�<��<C�<��<$��<ވ<^X�<��<���<���<u'�<��<�,z<�3s<�sk<�c<s�[<X%U<!YO<XhJ<YF</�A<��=<,�9<�5<�$2<��.<p,<��)<2�'<�X%<�"<֓<V�<~�<��<O<J�;-�;��;6q�;9��;��;���;զ�;X��;C�;���;�[�;2�;둌;�f�;�c�;V�m;2�T;d�7;#>;�)�:$�:��:'	):1��9��8�?P����]�?��r���Ԣ��ξ�.rպ���N7��
���|���$��y:�oNS�l8m���������;V��u���	w���"���1��w˪��������������̭�k󪻥馻�������u���b��#롻�u��|��`���������O����~»��ûd>Ż�ƻ�ǻw�Ȼ��ȻP�ǻ7�Ļ�������s��gṻM�������m6ǻa�λ��ջ��ۻ����㻘0�R軖k�Â��� |��r�y��ع黺������&�V0�g������	����(�HK����]	���
�����#��T��q�LE����������:�E���-�ǩ�t|�T��H�zJ�6����  �  �2�<���<���<�N�<A��<w��<���<���<���<A��<�c�<�K�<��<���<m��<+x�<`�<&�<O�<�`�<\|�<?��<��<�P�<j�<���<J��<�l�<���<9��<���<���<��<��<->�<��<�#�<�X�<�w�<���<���<���<g^�<���<=��<X��<��<㵿<�b�<u�<{h�<pտ<��<���<��<���<�Q�<3��<uy�<���<�ͼ<��<��<ډ�<�Ӹ<��<x��<<��<�"�<�6�<�Ȼ<��<]ѹ<�v�<a�<�<��<�q�<��<���<?��<���<L��<�i�<��<�~�<��<h��<�ǋ<,C�<_�<�T�<�7�<ځ<7ف<5��<��<�Q~<kMx<�p<R\f<�/\<��R<��J<��D<0�@<��><��=< I=<0�<<k;<�V9<�z6<�3<�J/<�G+<�&<p["<#K<��<J<.<<�F <0 �;;'�;>x�;B��;տ;�Ű;[�;��;���;� �;! �;���;�ց;XӀ;�Ny;B�g;��L;m�);�;��:��P:Jj�9S�i7`�H�B根�¹�ݹ0w�4  �#�K�:W���ꟺ~���c��������$�1}7�$cJ�y�\�Jn��;~�Pކ��̎�'q������b������˼�J�»��Ļ�»��T���k�ɷ���렻+���;���_��"_��!'ƻ|�λ��ӻ�+ջ�ӻ�λ��ȻBaûͷ������Ĺ�����������a���p���"��X��x��������pŻk&ɻ�ͻ*�ѻ!׻%*޻��V������
 ��}��%����{���C�����}�黳Z���뻎��FO��F���������{������#�Z������
�h&	�����	��Z	���	��*
�^�
�{���A����w�����5�r}��  �  ���<
��<�<�<�_�<�[�<���<���<d\�<�j�<���<t��<v��<Tx�<#�<\8�<��<Lg�<VS�<^�<bh�<~��<�<<��<o��<4�<7�<^��<��<��<M��<̥�<���<i�<�<�<A��<y��<��<	i�<~F�<v�<��<���<���<,[�<e�<�C�<���<2H�<��<�N�<� �<]�<��<��<8��<{��<��<'��<g�<Sc�<n�<�D�<|o�<}#�<p<�<NU�<T�<�t�<�w�<���<>��<�ݼ<PL�<Q>�<��<�t�<8��<@��< 4�<_�<l��<P5�<}�<J;�<$A�<l��<�$�<��<��<�d�<��}<pgy<�-x<)Xy<�{<��}<��}<�#{<�t<nRk<��_<S<�_G<��=<��7<y�4<��4<�l6<�(9<��;<i=<��<<o�:<��6<c2<�,<�&<]!<��<�d<�<5<_�<K�<8��;t��;���;���;G޷;�K�;z�;H[z;U�b;Q�V;��U;�^];�gg;��m;�yk;7�[;�?>;
�;t��:w,H:֝�8��!�H���j��Dd�B�D����q���Q�����=��(��E���ٺ�����n�*��;��?I�z�U��]a���m��|��X�����73������j�Ļ|aһ��ۻ��޻h�ۻ��һ6ƻ|������?����:��򾯻�����;̻ �ۻ���zI�Ӣ6���߻Ԣӻ��ǻ�������g����氻�Q�� ���#��zﺻ\V���
����������4�� L»(�Ļ��ɻ�
һŴݻ&������q�4���m��?�w���	���B���jn���D��P�����+���������!_�bh�1��p����%f�ؼ����}8����o��V
�v����	���P�<��Zx��v��V��  �  �@�<��<z��<�L�<+��<� �<4\�<���<���<=	�<l��<���<1��<���<..�<c8�<xT�<;�<o��<�F�<�?�<�C�<�Z�<�%�<��<(K�<<�<�F�<��<֩�<�3�<u�<D��<�^�<|S�<з�<���<���<v1�<�y�<�H�<G7�<$��<y�<���<���<��<UF�<2g�<=|�<뮱<���<&�<HL�<���<Y��<���<�*�<P �<��<��<��<���<d�<��<\>�<b(�<�<�c�<h}�<�)�<�u�<�<-�<FA�<Y�<R��<�:�<V,�<�[�<Ҙ�<���<�<���<r�<V$�<nt�<�l�<���<�x<I�o<t�k<8�k<x�n<,s<Lw<1y<c	w<�p<a�e<F,X<�|I<��;<��0<�*<��'<)<zF-<��2<8<��;<L=<��;<�;8<��2<�$,<U%<h�<�<�<��<Cb<K�<n�<;_�;���;r��;a��;�`�;}8�;�ln;�F;9�+;f|!;�b&;V�5;Z�H;�EW;�Z;(L;�0,;���:�҇:��9;�*��{��)�Ϻ�ٺҬǺWƣ��}s��d*����$���zW%��p�����+�ݺv	�� �n�3���B���M�5�U�\�]���g�H�w�[击|Y��D���=�»�@ػ�K껍@���-���x��G黤aػ��ƻw�����w����幻�*ʻ�޻'��e� �6������� ����w�ҳл���nǵ�p����-��l�����(?��(J»��ûa�ûAl»�����6��»R Ȼ2�һ1��1������q��+��������_����$a��T����+���ղ��,n�������"�'�)��Q-���,�}�'�3� ���A]���	��P�M���������������K�	�w����ld�|���<���  �  3��<B��<�]�<
�<ϊ�<��<���<˄�<t�<���<�^�<�q�<���<R��<t(�<���<T��<���<�\�<���<5f�<�B�<���<N�<���<�G�<�I�<8�<A��<��<��<g��<���<�Q�<{�<�g�<�h�<d��<��<�:�<�&�<|��<�:�<G��<�\�<H�<v�< ˮ<Jw�<���<F�<�ӯ<��<�#�<`j�<E��<Ǉ�<���<.�<!��<O�<V�<ͤ�<?h�<ل�<�o�<^�<�h�<M��<]��<>Ƚ<B�<�Z�<挸<V�<��<�;�<H۬<^ �<���<�<cZ�<أ<��<��<�<�<��<�^�<#_y<�l<z�c<��_<:�`<MOe<��k<�rq<�st<f�r<X?l<p�`<�Q<�A<Ƕ1<"�%<n%<��<�<�p$<�,<f�3<L9<s<<,�;<��7< 2<:�*<�i#<�W<'H<C�<��<� <�0<B�<:f�;�l�;�|�;��;�/�;�s};h<D;�8;n��:���:�I�:�R;~u-;M'B;5	I;xg<;\�;���::��й�*��g����5�l����rr��=�f�}d�&�	���(��s�'������,���9*���=�%�K�b+T���Y�7>_���h���y������F�����g$ѻO��g �������6��c����q��8ӻ�����D��HƸ��û�mֻ���&r���{��������Wj��x��HۻҞǻp��Ѱ�^���pp�����К���}û�ǻgɻ�Ȼ�yŻ�»�����»��ɻ��ֻ &���z������#���(���)��&%���T���!	���3��x��	����*.!���,��T5��Q9��A8���2�i�)�II�v��V���,���8����
��������cQ������	������j��  �  ?�<I��<f��<���<af�<a�<
z�<qd�<G�<1c�<�n�<H�<�
�<�(�<`��<�W�<$��<)�<�K�<�[�<�h�< �<q��<�{�<��<I��<d��<�3�<)	�<��<��<�<�<�U�<�{�<T�<�g�<���<�1�<� �<���<���<�q�<�j�<��<�b�<�d�<5��<��<L[�<am�<EJ�<L��<�$�<��<⨼<�6�<v�<�<�ʶ<aL�< ϩ<���<���<�E�<u��<� �<&��<eS�<SJ�<���<!9�<�ټ<��<���<!��<U.�</�<�ѫ<D�<�ɨ<<��<�i�<f}�<W�<	��<T>�<}h�<�7r<�d<)w[<c�W<_Y<	�^<e�f<�^m<? q<h�o<�%i<��\<h�L<Qh;<��*<~�<�<��<;
<s<�'<e�/<<�6<\�:<A�:<�I7<�F1<G�)<~�!<#r<G=<&�<�?<"�	<I<�<��;���;���;��;fG�;�'d;�s&;�]�:�ȴ:tѧ:z_�:��:�;H3;��<;W�0;��;gŮ:�N�9�H�����Z�P�7�ӫ9��1(���	�lͺ�\����>�>R�b4�<�}����N-�`���1���E���R���Y�0�]�8b��1k��^}�׍��t�� ^��<�ۻA(�� ���(��'�{�L�d���ۻ��Ȼ�Y���ξ�cʻ��޻x��u���� ��0������=
�����X���+ͻ<~���ⲻC*��z�P��3o���ǻ�~˻@�̻({˻ ȻYoĻ�c»�4Ļ�˻;�ڻA�|����!��t+�9B1�l�1��v,��5#�`���-�#m��~��:�L�gF���&�=�3�Q=���A�h@�+:�j40��Z$�<��u�����>��=���i�3��8������"8��i�y��8w�:��D��  �  ��<�,�<���<��<A�<��<��<��<䷻<�&�<|e�<�>�<^�<f��<K�<<��<3��<�<�<�6�<x�<���<��<�/�<�.�<"Խ<�!�<>�<���<���<��<��<|�<��<�*�<���<8�<�(�<���<���<��<���<�9�<��<��<⤽<g�<�]�<���<��<���<p�<LV�<�,�<�,�<��<@��<qu�<�h�<��<�Y�<&��<_=�<��<5˟<�4�<���<���<鋲<,��<�X�<���<r��<���<"ķ<�I�<�Ӱ<Sʭ<n�<���<&��<�W�<N¥<�7�<'9�<(~�<��<�g�<0S�<@�o<��a<�|X<��T<��V<U�\<p�d<C�k<n�o<@�n<6h<��[<�[K<�d9<�y(<�<=<F�<�X<K�<�/%<��.<6<�:<�L:<��6<5�0<P)<)B!<U�<y<^�<p�<E	<�<Yz<F��;�b�;��;�S�;���;w�Z;�;��:�.�:j��:y��:j-�:��;��-;�8;�s,;�a	;I��:�R9i�j�
���*�ދC��E��x2��~�spں�ꕺ�dK�k^$���9��W��ӓ��D���b����4��H�CU�S�[��T_��]c��sl�
��%��5x���M��E�߻. ��k�
���V�Z+�^��B��r߻�e˻����,	����̻����@��A����?�������
��N ���YPϻ"轻.ͳ�ٰ�ʝ��������fȻ��̻�iλ��̻(ɻ.9Ż?ûq�Ļ�̻�0ܻݗ��"������#�gN.�g64� k4�g/��k%�������i��ܙ��^�5��	����(�6���?��|D��SC���<�r�2�:&����������<�a@����������M�q�i�����X�`��э�����  �  ?�<I��<f��<���<af�<a�<
z�<qd�<G�<1c�<�n�<H�<�
�<�(�<`��<�W�<$��<)�<�K�<�[�<�h�< �<q��<�{�<��<I��<d��<�3�<)	�<��<��<�<�<�U�<�{�<T�<�g�<���<�1�<� �<���<���<�q�<�j�<��<�b�<�d�<5��<��<L[�<am�<EJ�<L��<�$�<��<⨼<�6�<v�<�<�ʶ<aL�< ϩ<���<���<�E�<u��<� �<&��<eS�<SJ�<���<!9�<�ټ<��<���<#��<W.�</�<�ѫ<I�<�ɨ<�<��<�i�<o}�<a�<��<^>�<�h�<�7r<�d<;w[<s�W<_Y<�^<n�f<�^m<C q<i�o<�%i<��\<`�L<Gh;<��*<o�<��<��<(
<`<�'<R�/<*�6<J�:<2�:<�I7<�F1<>�)<x�!<r<G=<(�<�?<*�	<I<�<��;��;���;�;�G�;�'d;�s&;�^�:�ɴ:�ѧ:�_�:C��:*�;H3;��<;X�0;��;7Ů:�M�9��H�^��[���7��9��1(���	�ͺ@]����>�cS�s4�5�}�~����-��`�Ҷ1�ưE��R���Y�<�]�@b��1k��^}�׍��t�� ^��<�ۻA(�� ���(��'�{�L�d���ۻ��Ȼ�Y���ξ�cʻ��޻x��u���� ��0������=
�����X���+ͻ<~���ⲻC*��z�P��3o���ǻ�~˻@�̻({˻ ȻYoĻ�c»�4Ļ�˻;�ڻA�|����!��t+�9B1�l�1��v,��5#�`���-�#m��~��:�L�gF���&�=�3�Q=���A�h@�+:�j40��Z$�<��u�����>��=���i�3��8������"8��i�y��8w�:��D��  �  3��<B��<�]�<
�<ϊ�<��<���<˄�<t�<���<�^�<�q�<���<R��<t(�<���<T��<���<�\�<���<5f�<�B�<���<N�<���<�G�<�I�<8�<A��<��<��<g��<���<�Q�<{�<�g�<�h�<d��<��<�:�<�&�<|��<�:�<G��<�\�<H�<v�< ˮ<Jw�<���<F�<�ӯ<��<�#�<`j�<E��<Ǉ�<���<.�<!��<N�<V�<ͤ�<?h�<ل�<�o�<^�<�h�<N��<]��<?Ƚ<B�<�Z�<錸<V�<��<�;�<P۬<h �<���<�<qZ�<أ<��<��<�<�<��<�^�<H_y<*�l<��c<�_<U�`<dOe<��k<�rq<�st<h�r<T?l<f�`<ٌQ<�A<��1<�%<N%<��<��<�p$<�,<A�3<[L9<Q<<�;<��7<�2<(�*<�i#<�W<&H<H�<��<� <�0<[�<tf�;�l�;}�;��;�/�;6t};�<D;9;y��:���:tJ�:S;�u-;|'B;M	I;yg<;E�;8��:�:��йz+��Y���t6�������s�O򨺤�f��f�\�	�ɡ(�Ȟs�����=��{��:*���=�N�K��+T���Y�F>_���h���y������F�����g$ѻO��g �������6��c����q��8ӻ�����D��HƸ��û�mֻ���%r���{��������Wj��x��HۻҞǻp��Ѱ�^���pp�����К���}û�ǻgɻ�Ȼ�yŻ�»�����»��ɻ��ֻ &���z������#���(���)��&%���T���!	���3��x��	����*.!���,��T5��Q9��A8���2�i�)�II�v��V���,���8����
��������cQ������	������j��  �  �@�<��<z��<�L�<+��<� �<4\�<���<���<=	�<l��<���<1��<���<..�<c8�<xT�<;�<o��<�F�<�?�<�C�<�Z�<�%�<��<(K�<<�<�F�<��<֩�<�3�<u�<D��<�^�<|S�<з�<���<���<v1�<�y�<�H�<G7�<$��<y�<���<���<��<UF�<2g�<=|�<뮱<���<&�<HL�<���<Y��<���<�*�<P �<��<��<��<���<d�<��<\>�<b(�<�<�c�<i}�<�)�<�u�<���<1�<KA�<"Y�<[��<�:�<c,�<�[�<䘨<���<�<���<��<q$�<�t�<m�<���<x<y�o<��k<^�k<��n<3,s<'Lw<<y<f	w<�p<S�e<0,X<�|I<��;<a�0<�*<��'<�)<DF-<L�2<�8<{�;<�K=<l�;<�;8<f�2<�$,<U%<^�<�<�<��<Yb<h�<��<�_�;D��;֗�;���;a�;�8�;�mn;PF;��+;}!;Jc&;��5;��H;�EW;�Z;(L;�0,;%��:�ч:8�9�+�<}����Ϻ��ٺ~�Ǻȣ��s�h*�����f���dZ%�=p�篨�3�ݺ�	�E� ���3�׿B�'�M�U�U�q�]���g�P�w�^击~Y��D���=�»�@ػ�K껍@���-���x��G黤aػ��ƻw�����v����幻�*ʻ�޻'��d� �6������� ����w�ҳл���nǵ�p����-��l�����(?��(J»��ûa�ûAl»�����6��»R Ȼ2�һ1��1������q��+��������_����$a��T����+���ղ��,n�������"�'�)��Q-���,�}�'�3� ���A]���	��P�M���������������K�	�w����ld�|���<���  �  ���<
��<�<�<�_�<�[�<���<���<d\�<�j�<���<t��<v��<Tx�<#�<\8�<��<Lg�<VS�<^�<bh�<~��<�<<��<o��<4�<7�<^��<��<��<M��<̥�<���<i�<�<�<A��<y��<��<	i�<~F�<v�<��<���<���<,[�<e�<�C�<���<2H�<��<�N�<� �<]�<��<��<8��<{��<��<'��<g�<Sc�<n�<�D�<|o�<}#�<p<�<NU�<T�<�t�<�w�<���<?��<�ݼ<SL�<V>�<��<�t�<D��<N��<04�<s�<���<i5�<'}�<h;�<DA�<���<�$�<$��<��<�d�<��}<�gy<�-x<QXy<<�{<ɵ}<��}<�#{<�t<]Rk<��_<�S<�_G<��=<L�7<<�4<V�4<ul6<P(9<h�;<*=<��<<:�:<e�6<<2<Ì,<�&<Q!<��<�d<&�<P<��<v�<���;���;P��; ��;�޷;L�;��;@\z;<�b;#�V;Q�U;_];(hg;�m;�yk;9�[;�?>;��;���:*H:&��8#���H���j�Id�x�D�&��͏��h����u�=�7*���F��ٺ���a��ʋ*�E;�@I���U��]a���m�'�|��X�����83������j�Ļ{aһ��ۻ��޻h�ۻ��һ6ƻ|������?����:��򾯻�����;̻ �ۻ���zI�Ӣ6���߻Ԣӻ��ǻ�������g����氻�Q�� ���#��zﺻ\V���
����������4�� L»(�Ļ��ɻ�
һŴݻ&������q�4���m��?�w���	���B���jn���D��P�����+���������!_�bh�1��p����%f�ؼ����}8����o��V
�v����	���P�<��Zx��v��V��  �  �2�<���<���<�N�<A��<w��<���<���<���<A��<�c�<�K�<��<���<m��<+x�<`�<&�<O�<�`�<\|�<?��<��<�P�<j�<���<J��<�l�<���<9��<���<���<��<��<->�<��<�#�<�X�<�w�<���<���<���<g^�<���<=��<X��<��<㵿<�b�<u�<{h�<pտ<��<���<��<���<�Q�<3��<uy�<���<�ͼ<��<��<ډ�<�Ӹ<��<x��<<��<�"�<�6�<�Ȼ<��<aѹ<w�<h�<�<��<�q�<0��<���<X��<���<k��<�i�<�<�<2��<���<ȋ<OC�<1_�<U�<�7�<5ځ<Hف<B��<�<�Q~<cMx<qp<4\f<�/\<\�R<y�J<��D<��@<��><��=<�H=<�<<�j;<�V9<]z6<�3<�J/<aG+<�&<c["< K<��<^<L<E<�F <� �;�'�;�x�;Ѣ�;�տ;[ư;�[�;���; ��;!�;� �;�;2ׁ;�Ӏ;�Ny;C�g;��L;�);q�;|�:��P:c�9��h7��H�jM�¹�ݹ�{�� �l�K�8Y���쟺���ͬ�l�s���$��}7�acJ���\�in��;~�Vކ��̎�)q������b������˼�I�»��Ļ�»��S���k�ɷ���렻+���;���_��"_��!'ƻ|�λ��ӻ�+ջ�ӻ�λ��ȻBaûͷ������Ĺ�����������a���p���"��X��x��������pŻk&ɻ�ͻ*�ѻ!׻%*޻��V������
 ��}��%����{���C�����}�黳Z���뻎��FO��F���������{������#�Z������
�h&	�����	��Z	���	��*
�^�
�{���A����w�����5�r}��  �  ���<1��<.�<�s�<���<`<�<ǯ�<�N�<�>�<���<9�<�<B��<���<Ֆ�<Օ�<*�<S�<�#�<�Z�<?��<���<z�<���<��<a�<��<�]�<8�<*�<���<vd�<�A�<���<�7�<���<���<Q�<�}�<��<#
�<���<?��<�\�<}��<�{�<�<��<�i�<�Z�<(��<�Y�<�Q�<�W�<5&�<{�<�*�<2�<���<��<;�<=��<���<���<���<;Y�<�<�Һ<C�<	��<��<Wk�<W�<���<;�<�ִ<"�<'��<uW�<3��<>��<���<���<�˚<:�<<ON�<�<h�<<��<E��<#ވ<yX�<��<���<���<}'�<��<�,z<�3s<�sk<�c<A�[<%U<�XO<hJ<F<��A<m�=<��9<��5<u$2<G�.<:,<��)<�'<�X%<�"<ԓ<_�<��<��<y<lJ�;�-�;7�;�q�;���;���;.��;j��;罨;�C�;���;e\�;��;.��;$g�;d�;X�m;�T;�7;�=;a(�:��:�}�:�):-�9�8�RP�R��4�?�/u��ע��о�tպ����8�����P}�\�$��y:��NS��8m���������BV��y���w���"���1��w˪��������������̭�k󪻥馻������u���b��#롻�u��|��`���������O����~»��ûd>Ż�ƻ�ǻw�Ȼ��ȻP�ǻ7�Ļ�������s��gṻM�������m6ǻa�λ��ջ��ۻ����㻘0�R軖k�Â��� |��r�y��ع黺������&�V0�g������	����(�HK����]	���
�����#��T��q�LE����������:�E���-�ǩ�t|�T��H�zJ�6����  �  �7�<��< ��<���<���<���<"��<k��<��<���<��<��<._�<��<~�<���<q��<���<z��<m��<ٹ�<Hh�<8��< ��<��<&.�<��<Zy�<+��<~��<e��<��<���<�g�<�I�<�<��<�A�<tW�<�h�<C��<�W�<ʼ�<��<���<%A�<k��<V��<B��<��<*[�<�z�<��<Ġ�<N��<v�<V�<��<���< �<*J�< d�<�W�<��<F�<G�<,��<#�<�ʵ<+�<6��<�]�<2��<�X�<�س<U��<�l�<>گ<#�<�J�<�&�<�)�<Ә<%y�<Z/�<�ˑ<��<���<{�<5[�<?�<G��<���<%�<���<@Ƅ<"m�<V�<p<z<�at<ZXn<tMh<�_b<��\<
�V<GP<VjI<�B<9~:<n23<:�,<�l'<��#<�,"<�!<��!<��!<��<�<�<JJ<<O��;�8�;���;G��;���;X�;Ũ�;h��;�@�;�u�;e�;��;�Ӣ;��;#ْ;L�;�~�;�*l;r�U;�>;�%;��;���:�G�:��:9b+:aX[9>특�WC�󡝺Y=Һ/&����
�����������|��}�+�D�D�ud�8���><���^��ym���ұ������aJ��~֨��Ƥ�)Ρ�I����,�����������F��;��������b�������{��y^���o��  ����������N_ɻƢѻX�ػmvݻ?�޻r$ܻ�ֻ��ͻ/�Żc����1��I����zƻ�л"�ܻ��Z�sQ��h�������������.軂q仙.��E��8����	�Ȳ�G��0��G軫;����.�)��$���aG �l[��,�-��ba�}��"��1���]�������ǉ��X�A=���6�����e �ȵ%��)��  �  ٩�<�<���<.(�<-��<��<���<j��<w�<��<"�<��<�-�<�V�<r��<�.�<���<ۚ�<+P�<Z��<���<��<���<*�<K�<�Y�<w��<�F�<*�<�x�<�T�<�1�<�[�<��<1��<�u�<2��<3_�<aR�<�:�<pڼ<�Ǻ<�J�<PN�<z�<�P�<AN�<��<���<��<�h�<*�<��<l��<M;�<��<RV�<)(�<��<��< ��<eq�<v\�<9v�<��<0	�<S��<�ݳ<�@�<i��<~<�<�I�<��<^N�<���<Զ�<O�<�N�<\�<�-�<�ݝ<ė<n��<���<=�<|��<��<i>�<vb�<��<q�<ގ<��<���< Ň<�Ԅ<��</~<f�x<��s<�o<��j<a�e<��`<�.Z<i_R<�I<��><��3<F~)<�� <�M<;�<I<$�<�w<@g<-G<�<t8<�M<J��;���;�3�;�[�;F��;r)�;�ͧ;���;	��;�Q�;���;�C�;	G�;�;�;C�;�ɔ;a�;#{;�d;�7P;1�<;SX*;�;�q;�i�:��:��?:3� 9�&��g��&��e�*�2��a>�y�>��7�B-��+'�G*��h9��U��"|��㓻�8��
��D�ƻ`�˻Pʻ�=û<7���/��h#�������I���񖻤җ����@}��Rڞ�����̡��-���
�����v塻'Q������㭻$9���ŻggԻ���.ﻌ��2������'C��޻��ѻL�ǻ��û�;ƻ݆ϻ��ݻGg��.��7#�gW��d�æ��� �Ȇ���I��Ở�ۻ�ٻ�Sٻ��ۻ �޻�����廸�軺�껨F�H�K����"@�Z���"�Gh��������~��w$��'��`(���%�� ���������d�O-��!�y�)�`1�w�6��  �  "��<d��<�<���<���<{��<�<��<���<�b�<kE�<���<Jb�<�0�<�h�<��<�)�<*o�<S��<�o�<�i�<�@�<Z��<^?�<���<���<���<��<-?�<��<ň�<�l�<���<EN�<�g�<Rg�<.0�<�$�<0�<�ݺ<Ș�<��<��<��<u:�<�_�<3��<L��<���<݌�<��<��<���<wm�<�L�<�{�<}�<�/�<h��<��<mg�<%�<]��<�j�<G��<i��<#8�<*ή<�)�<��<���<��<d�< �<L��<Q�<���<�J�<[�<ѻ�<�T�<I.�<�B�<�C�<Nu�<u��<[�<�؊<Bc�<&L�<e�<U��<M��<���</��<[8�<�ـ<Q�{<�gv<r<�Xn<��j<��f<�a<*�Z<ډQ<L�E<��8<32+<�g<+�<�<Yf	<�
<�<�g<}b<t�< <��< �<�X�;v�;<~�;��;�;���;&��;x��;ֵ�;���;�̶;9��;���;���;8�;���;�ǅ;!~q;ddZ;o�F;^�6;p<(;��;��;���:�3�:;�&:Qt��a�{���E�(���P�9j�*Ks��m�,�]�JEK�o�=���;�tiJ�M�i�=���>���羻�@ԻO-�.�VB��cػ�ɻ
g�����\���o���@���ە�����c��Ꞣ�;���𽦻���!'��W���R��ѕ��o𤻊.������ϻ@��6o����� 	�� 
���� �2�r)߻oһ��˻�λ*ڻ-�n ��z
�s�������,����
��4�<��%D��kۻ��ֻc�ֻ�ڻdl߻W&廔2�D������.�����)��;�������^
�����z�'�)��F1��5�l�5��1���*�U�"������4w�h��q����(�O�3�]=��D��  �  ���<���<4��<�x�<���<r��<���<���<W��<�<�<���<4)�<�a�<!��<��<���<%;�<V��<�[�<wM�<.�<Κ�<qq�<���<j��<p%�<���<gɵ<�@�<�@�<���<d@�<�c�<���<_I�<�^�<���<�3�<E�<L4�<-,�<��<ɇ�<�j�<�M�<q�<3��<��<���<y,�<���<6z�<�5�<���<C4�<�2�<���<��<��<מ�<�3�<��<���<v��<���<E�<Iq�<t�<���< �<N��<s��<ol�<13�<�Ǫ<��<��<�I�<��<&��<X�<`S�<���< \�<ٚ�<�G�<[̃<U�<���<�ߍ<Eh�<�M�<���<�Ê<,�<X�<w]<
�x<��s<��o<��l<�j<(�f<�da<�Y<CO<I�A<��2<_�"<�<�?<�� <�i�;�;��<A<��<�I<�<!~	<�u�;���;�Һ;��;��;$r;��l;c�y;]��;�
�;y��;J �;щ�;�D�;�
�;��;�͐;ݩ�;C=g;GuO;d�<;��.;7�";;�+;���:���:�#�9��ٹ������)T�H+���O�����)��/��f�1�R��]M��[�Ҭ|�O2��ʆ���ѻ������L3��p����4���ػe�ûNE���(������ݔ�ͩ��(���������� �����������Iq������栻�!���H��>����:ûi�ٻ��
^����������|
�p����B뻱�ۻ�&Ի]׻h)以���ߤ�.[��U���!��!��s�a���X	��m���'�yF޻��׻23׻'ۻ��6�����G󻨛��������ﻋT5������g`����P�'�?�3�Y�<���A�~lA��n<�&�3�o�)�Wx ��.�����6\$�S�/��v<�(�G��O��  �  ���<��<?,�<�]�<^W�<��<���<���<�*�<���<C�<��<ȓ�<2��<��<���<�w�<H�<6��<{��<^��<��<�7�<��<���<�<�׵<���<M$�<Uc�<��<�i�<�<~��<���<���<�1�<'�<\��<�
�<�}�<S�<f�<x�<̯<���<�ǻ<s~�<���<���<t��<N�<|��<���<}W�<�6�<��<�/�<��<��<���<��<V�<u��<���<��<w��<��<���<K�<���<��<>�<<�<+^�<��<:Ш<G:�<�v�<�<��<��<z�|<oy<��z<���<綄<j�<ߜ�<��<^َ<�N�<�d�<g��<t��<�}<��v<e�q<^In<}�k<�i<�e<ȋ`<�X<� M<��><�-<��<��<G0 <�|�;�w�;���;�<�;,Y<1�<2<<�\<K��;4(�;k�;��;D�l;(ZQ;��L;��\;)�z;}v�;:Ԡ;�­;X�;ʜ�;͢�; ̝;U�;پ|;&e_;�.G;5;�6(;�;Hm;� ;� �:+�:0�9��)���ߺ)*5�B�r�t����䝻R1���ޘ�
S��"�x�za�4Z�FVg��#��߃�����h{޻_���1�3�����gN�����K�̻JH��M�LF���e���#���|��@��V��L����ﯻq'��^;��a����c��/���ki���%����Ȼ�7� �� B�k��2�����?��O"���T�[+ڻ�;ݻ5A��� �?1�����$��%*�F�)�f$��z���2��P�sn��ٻs�ػ,�ܻ���α�O�����{��Q�����i��[��k��@���'�m���s�P�-��:��D���I�V_I���C���9��.�^$�oh�I{��=��)(�8�4�gB���N���W��  �  �<2�<P��<O�<k
�<b��<ַ�<��<���<(��<�E�<�q�<�'�<���<w+�<<��<k��<��<�o�<D~�<�a�<͒�<@�<�N�<y�<1��<��t<�-g<�b<�dh<��v<�I�<���<cΘ<+(�<�Ǟ<wv�<}�<�ن<]�v<чc<��W<4�U<
�]<� n<�ށ<�Ѝ<UC�<���<��<@t�<�_�<V��<�ɯ<�ɮ<��<A��<�ܭ<%H�<��<�ݭ<���<�ͦ<�@�<		�< ��<��w<^�_<1L<�x@<�3><oQE<��S<*'f<�w<(�<��<~�<̿q<��Y<HD><�[#<��<�� <��;��<�?<b&<�:<�M<$[<��c<9�f<"�d<}�_<{Y<�+R<��K<=PF<X�A<�=<��8<Q�1<~'<	=<�<���;�ߜ;��H;���: L�9���q���9ߵ�:F;�I;Gn;��n;ױG;V�:Q��99��;��]��}��9����z��x6��ʺdĝ�neH:���:�'�:��;6��:	d�:���:�m/:G��9�^��B���S�&Gb���������L���%pȻ��5�-u5���F�1�N��L���B���2�l�!�87�Д��6��w�D�0���I��vc���x�&#���ل��n���cs�2+^�[�F���/�8u��� F�/F��� � ����B�����;��@����X��O	����j|!�Ρ5���M���f�Bi~��q������)���y���
����l�7X�x4H�3W@�SB���M�
a�x��&��H���*��t����������]s�2�[��#F���4��(��"�� �(!�NV#�C�%�"�'��}(��(��@(��(�"�+�a42��=�ZZO�Øe���~��F��m���f���D壼]͢���T瓼�\��4y�0Cr���m�d�s�$2��6͋�����&4������  �  �M�<�b�<�ь<�b�<���<۞�<�b�<*ݽ<���< ��<O�<U��<�L�<\&�<�_�<��<��<l�<x�<��<>��<(��<|Ǫ<�q�<�	�<��<ٗy<�-l<]�g<�7m<C {<E�<H`�<��<�E�<`ߟ<T��<US�<x��<q�z<B'h<�\<��Z<��b<�Er<���<�#�<*-�<�<2`�<m��<�h�<���<��<��<�5�<��<��<�c�<���<��<���<��<ş<f�<�$�<R{<q�c<n�P<߁E<�2C<(�I<��W<&�i<v�z<^D�< �<��<�)t<s�\<1�A<'�'<q<��<��<�I	<�@<
�)<+�<<~�N<�\<d<еf<�d<��_<-WY<��R</L<��F<�
B<a�=<Q�8<� 2<��'<��<�<�;�;�ZW;	I�:1�%:�Wh�D�w�D�9�ĩ:�;��S;�-w;��w;��P;wS;�:�͏��i)��7q�y]���F���h�'o'�������6�%�]:���:�� ;4;�K�:
��:�h�:��5:7y�9\857㈹8�
��`�tî��C��I�g����û����:��0�H�A���I�`H�YL>��3/���@��[Q����s�O.���F�Li_��+t�i����M���~�Yo��Z�D�C�j�-�vV�ދ� ��2��� � ��8��p��O�}��~�������	�7��q ���3�K��pc��7z�I���$������"����}��i�NhU�'�E�'&>��@�zK��&^��|t�x���P������𐼮���A�$p�iY�C�D���3�>(��!�V ��� �3#�4s%��9'�X(�4(��(�w�(��y+���1�@Q=�N���c�|�_n���v��ć���Y���T��L˚��������|�p�o���k� Wq����<��׬��n���.���  �  s�<TL�<z�<q��<E|�<�\�<��<���<���<H��<@�<2��<��<��<��<~�<�U�<��<pd�<��<��<��<X��<#t�<K�<�h�<%7�<�0z<�v<��z<,��<TH�<��<���<�d�<Z�<o�<�7�<BE�<��<2u<��j<7(i<�	p<T~<�m�< ��<���<Y֤<��<Q��<.S�<���<M�<�P�<ﱮ<1d�<�i�<��<5��<�ͭ<٭�< ��<��<B�<��<�M�<_o<�1^<�S<�>Q<�W<�`c<ws<,,�<���< �<
�<��z<��d<��K<\i3<��<��<�<_4<�Q"<K2<�6C<8xR<W^<8�d<B�f<�d<��_<��Y<�XS<k0M<��G<ϺB<�><��8<�1<�,(<�b<�<���;l	�;l�;��%;���:Ad:3�O: y�:=� ;�b<;ejq;�f�;�Շ;.�i;N^#;�2�:�L���F:�(�[�ĉY�q17�{����f�5
&9&�:��:�o;G�;�w�:ũ�:㵕:9xE:��9�Ɛ8si����]a��C��Yb��	A��f��{���6��>�*�#���3��E;��e:��2�x�$�I�X�
��������a��$&��<���S�g� s��Ov��p��8c�' Q���<��?)�X��lk�����Y�@� ����u�����Q�p�e��|��B��[	��b��4n/�,D�Z�{�n���~��
��Vn��*����cr���_�jtM��?��8���9�݋D���U�j]j��~�����kj���剼y<����z�Zg�S�l�@�w�1�1�'���!�d. �+� �#�"�P�$�H8&��)'�ʊ'�W�'��(��+�W�1���;�SK�`^��at�9\��{T���Y5���_��Po���y��e8��(\u�K�i���e���j�gyx��˅�K������pE���  �  N�<,K�<]�<͢<0Ī<Ҵ�<���<���<�e�<� �<p��<�Z�<���<��<a�<���<�`�<s��<ϳ�<c̽<��<���<S��<s7�<+�<d�<�c�<�?�<i|�<	h�<	��<��<��<J��<��<yH�<D��<��<�M�<?�<m6�<d�<��}<<9l�<=�<�Q�<kD�<���<y�<��<$��<�
�<��<�<~(�<�ݮ<���<�{�<��<{�<� �<yk�<��<���<��<`��<��<}:q<�'h<s�e<bVj<�Zt<c��<g��<�R�<c�<i_�<k�<�q<֎Z<e�D<�j3<m(<I�$<~�(<��1<
><�K<ȰV<�T_<�d<ye<�c<��^<x�Y<��S<=.N<�H<�C<�=<F�7<�z0<6'<��<<�M�;2t�;�?�;��k;��/;,�;��;�;��A;5-r;���;��;�;�+�;��M;���:�n:��7��'ӺC���

�;M��n����|���:��:���:.�:�S�:�v�:��:I�:b1T:���9> 9K�Y����@�t�����=g���;�&(���I���pӻ�����m��"��G&�$A&�t���M��	�| ����+�����	�ۈ���.���B�x�S�c^�v~a�"]��kR���C��x3�A�#��T��a�K��������R�L���Y�������ɉ��f�	S
��L�c���W*�\;�S\M�f:^�ͥk��ns��$t�7�m��<a��Q���A��Y5��B/��1��m:��I��\[�aXl�Uy�w ���Z���w�J!k�:z[�|+K��@<�tI0�(�i#��!���!�x�"�h�#�L:%�}K&�R5'��G(��*�$-��2�(};��H�X��Aj��|�����Č�=ʏ��(������Y��f�x�`j��7`�]���a��m��o~�mR���r������  �  �ˡ<3~�<��<�:�<o��<�'�<p��<5��<�F�<h��<���<��<�*�<$��<�o�<��<+��<<Y�<�<��<S��<Y��<M`�<�2�<G��<v��<o�<n��<�o�<F��<��<���<_0�<���<�߫<�<^%�<ǐ�<i�<�T�<rb�<	��<Ÿ�<Yy�<`�<[��<�e�<��<Z��<BL�<ǫ<�[�<-U�<��<6,�<�'�<��<sZ�<ω�<�f�<�۪<���<��<6r�<��<���<��<x�<U#�<�g<Bz}<-Z�<"�<#�<铍<c��<��<�(�<��<��~<��k<�NY<z$J<p@<��;<,�<<
B<	hI<�bQ<�xX<y�]<$`<�c`<��^<��[<{X<�S<�GN<yH<*B<�[;<�4<�,<��"<C?<pp<DO�;w?�;��;4ʛ;�p�;�l;Wqd;�xq;~�;�_�;6��;���;��;�w�;̡~;_J7;��:a:C�E��)�CD����j��b�9��`:b�:�A�:��:J��:��:��:7�:4TS:X��9ӈ�8����qF9�)͘�a|ۺ�i�H�B��y�����y��&�ݻ�R��:��2�����
��;�����=�h]�%8��S��2%��>�)/�;?=�F{F�B�I��lG�{k@��v6�&=+��J ���������
��:�����������K�52������s�
�}�����*���t'�j�3��@�J�L�tsV��\��L\�*W��:M���@��,4��T*�
�%��&'�"�.�	X;���I���W��Xb��h�(Gh��]c�k�Z�J�O�l�D��P:���1��+��(���%���$��+$�^$�4 %��f&��6(���*���-�ɪ1���6��G>��G���S��`��cn��jz�W����胼�\��a!���u��Ui���]�_�U�bnS�ЇW��ka��&o�N	~�h���*b���  �  s\�<� �<��<��<W��<�L�<%��<oֹ<I��<�M�<R�<�O�<�d�<?��<��<��<���<�P�<���<�߶<��<��<��<��<{�<�}�<x�<��<��<�z�<���<Kƥ<7U�<�8�<X�<%��<y:�<���<6��<�%�<���<`�<#�<Xj�<P�<틚<�d�<>�<Ӣ<��<��<q��<�Ԫ<Qx�<?��<�:�<���<9�<�4�<���<��< �<�N�<�X�<.��<GH�< p�<^͏<�ǌ<1ӊ<-W�<�v�<��<l�<��<��<�c�<��<,M�<'E�<H�|<��m<��`<m.W<ÇQ<}BO<�pO<�Q<�GS<NCU<*�V<�W<,�V<*mV<��U<Q�S<R�P<�L<��F<��><Z6<��,<�>#<;�<�h<�<q�;��;���;Y�;E��;�0�;��;Qd�;+ͬ; B�;|�;���;x�;^S�;;��;k�r; T5;M��:m�:�E:h%	:e�9��:��9:1~c:��:�Ռ:Ǳ�:4�:@�:k݃:9�h:7�3:�9�Տ��3��L�ֺʏ�E�7�+^�^B��߀��g-��"û�ջ�l仳Q��fﻔ뻪k�ڏػ\ѻYiл�	ػ$��^ ����fZ�6�&���.�z	3�aj3���0�R�,��('���!�O��7 ������������X����������N
�ܑ��L�~:��g�#��k)�hf0��~7���=���B���E���D�m�@�[A9��0���&����b��F�b$�o-��s8�6C���K�k�P�UR�7�P�M�H���B�\S=�s�8�3�4�P1��-��*��Z(���&�;�&�8h(���+�-�/�3#5�w�:�tO@�GF���L�tT���[��@c���i���n�S�p��jo��{j�.�b���Y�_�Q��L�P�J�n�M�P�U��`�|k���u��}��  �  ��<QW�<>�<I;�<꠲<�N�<V�<<�<%(�<�4�<iڸ<m��<��<���<O��<� �<A�<�]�<DX�<D��<>��<�E�< ��<��<Bʦ<J�<��<*?�<��<�s�<���<�~�<c�<�Ʋ<��<��<0E�<�Q�<%��<���<�7�<�k�<�j�<[�<5/�<���<�V�<@]�<,˜<oӝ<���<2�<�?�<�N�<�ª<��<�ث<!�<J0�<3��<�؟<��<���<D�<ʖ<bԕ<�<���<��<M�<~>�<m�<���<��<�\�<���<x��<��<���<��< ǅ<�K<�-t<��j<c<��\<sW<p�R<}�N<��K<	6I<��G<1H<cI<�)K<�XL<��K<�lH<>�A<d�8<IJ-</!<�d<<u<Q<�;�-�;���;f�;�C�;���;f��;�\�;���;���; ��;���;o,�;?��;u�;���;޺�;�u;i5G;+;��:Nh�:�۝:�t:�{6:)�:��9p�g9��C9�s9�v�9�<�9�5:<�9d�9������r��׺q���JJ�K�q��=��$j��}m�����ch��Ժ�����XŻ�ǻj ƻ�
û�׿�䢾�ɏ��U�ɻ��׻^n��L��
��=�����% ���#�H�&��@(��+)�%P)�z�(�kp&�E�"��z��5����;��	� Q	�t���O�Bi�� ��'�:
,�5}/�.�1��-3�~4�\f4��)4�H3�H�0��-�4�'���!�^��C��R�����G.���!��_)�#1��7���<�S�@�	C���D�	 F���F�ײF���E���C���?���:��5���/�I,�Y�*���,���1���8���@���H��JO��gT��
X���Z�Vp\�+�]��o^�v^��]�>O[�NuW�SR�	�L���G��`D�i�C�|F���K�'>S�<V[��c��wi��  �  ���<c��<��<K�<eW�</ �<)�< �<1!�<�ܬ<�ݰ<�Y�<�S�<QԻ<�)�<��<�<_��<;�<��<�~�<���<��<���<t1�<�Ԧ<J��<>��<3�<=�<ϧ�<�L�<�Ǵ<ߵ<fV�<3�<��<��<(ɰ<�8�<��<�Ҩ<��<��<�<l�<�	�<W�<j̓<�ܓ<|��<�>�<�̝<���<h�<k��<�b�<��<4��<vG�<�<e��<��<�<�s�<�#�<wv�<���<1J�<�#�<.y�<�c�<^��<fH�<X �<�I�<_��<��<uP�<:�<@�<T�</d�<��x<ˡn<t�c<��X<�!N< +D<J�;<�6<��3<ߑ4<<8<?=<��A<ٹC<��A<��:< z/<�!<:�<�<�o�;��;
�;��;*��;�Q�;���;n/�;��;^h�;��;q��;�)�;,��;���;S��;�H�;�ж;�1�;C��;�|;z<Z;��4;$�;���:�l:��9拹��8����Y���en�{k'�(©�J���n	��䄹M!I�^�Ⱥx< ���]�a���󄠻fѮ�/ٵ�X+���Ҵ������?����j��ך��o����Q��ĭ�����������$�̻=�ڻ�"껸���R]����r�ű�]�"�z�*�,�1��F7�r:�GO:�ay6�jV/�_&�yu�^����T5������'��D2�d�:�|@�y�A�M@��n<��$7�I1��+���&�:""��8���������������;��7�`��O#���(�co.���4���;�	C�J��2Q�MBV�s�X�t�W�GS�G�K���B��I:�w4�2�1��74�'";��3E���P�t[��Gc��h�5Qi���g��c�S�^�RaY��aT�sP�d]L�I� �E���B�1�@��r?���?�R�A��.E�`�I��#O�
�T��}Z��  �  ��<J��<n��<���<4L�<4x�<�L�<퇝<���<-�<��<��<�<�<���<3�<�߯<�֨<"w�<�<2Ӗ<�A�<�n�<�ޙ<�Ȟ<�Z�<@Щ<��<9%�<���<��<:��<pd�</�<Q�<��<3�<v?�<���<�a�<;�<dC�<�7�<��<]ݝ<P�<w�<-�<!<)�<�]�<[�<�0�<��<��<H�<t�<럠<W�<=ړ<��<�d�<o,�<��<7ȅ<�Љ<K�<_�<�O�<!0�<w��<�<��<Ew�<�;�<h|�<�F�<ۨ�<ӫ�<xS�<��<i��<-�<�r�<��s<I�d<8fT<��C<,@4<�'<$%<�	<	><��$<�-<+�4<��9<��8<�|1<.1$<Ҽ<���;H_�;���;k��;8X�;VL�;.��;P��;��;(��;A��;���;��;���;��;�u�;4T�;���;�[�;Ͻ;C�;!��;;HW~;�\R;��;���:�X:���M\��oU�)��=!�:"��h�KР�_�N����OL��m���w�N�]�ه���嵻��λ
ܻN8޻L׻��ɻ+,��,�������׾��[���e��j1���ע��Ū�����`=���PǻS�ѻd�ܻŢ軙�����T<����w�$�W�2�4�?���I�suP��Q�-M���C��B7�I)*��H���y+�щ���*���8��gF�wFQ��wW��X�M�S���J��@��R4�kX)��3 �i����Z�@m����/d�D��˴�W+��:����9��4`��&��/�/l:��XG�?�T���`�tXj��vo�t,o��ji�|P_�%�R�N�F�>�e�:���=�a}F�G�S���b�h-p�ATz�N^���~�]y��gp��e��Z�ӠP�z�H�=C�I�?�?�=���<�T�<�F)=�o>�&�?�N�A��D��bG�n�K�&FQ��  �  ���<mU�<��<2�<%��<;��<�	�<2��<ؒ<$w�<�x�<m]�<�j�<���<{��<�<��<��<}�<��< �<�e�<�p�<���<×<�ڟ<K��<爮<���<;̶<H]�<Ǹ<υ�<���<�Z�<�ն<�p�<��<Ƅ�<|�<f��<�#�<?�<��<�y�<gf�<���<��<{Xz<Hlx<=�}<���<[��<K��<�Q�<��<V�<��<��<�]�<�ӂ<�x<mp<T�o<�tv<�+�<���<-��<~�<#��<�g�<{�<B"�<��<x��<���<:�<K��<��<�:�<�<�<���<:�<]�<�t<la<O�K<=6<��!< �<�V<�<��<��<J�<g�'<��.<�)/<�x'<G_<�<ǰ�;5`�;Pp�;�+�;10z;Ǉ;̓�;^��;�K�;���;�8�;x<>�<��;��; �;!��;U}�;���;���;�!�;6 �;w�;�:�;�Q[;J;N��:ʝ�E��as%�a�]���|���~���f���<�����Ǻ�?���������΅F�����hG��%H�xO��y�����������]�˻ղ�[�������_Y���������Ꝼ�{��������/�Ż68λ�yֻ��߻ @�8����
������+��[>�CP���^�;�g���i�6d��>X�;�H�|08�3�*��"���"�ɩ*���8�ΰI���Z���g��To�Huo��h��#\�_fL�C�;�M�+�������L�&���:����+��x������Z�' �{w�����m�"�3�.�1>���O�`*b��s�������u����h�r�@#c��S���H�8D�W�G��^R�mb���t�֦��ʈ�]���[ˊ�W�������Np��A`���Q�!�F��-?��5;���9�0>:�,k;���<��7>�NU?�/S@���A���C�iG��M��  �  p��<G��<"��<6��<�k�<?Ȑ<���<6+�<(��<tD�<ړ�<�ܟ<��<fo�<��<)A�<��<]�<���<嫆<f��<%�}<J��<��<ܐ<��<ж�<�&�<�q�<-Z�<� �<]�<���<�Ƿ<;�<�W�<��<_�<��< 5�<�:�<�\�<�+�<=��<�d�<�Z�<Ӏ<&vp<��e<U�c<:j<L�w<��<@��<BN�<ا�<!��<��<C�<��<�Tt<�{d<w�[<*P[<o]c<Mr<�b�<�F�<�c�<:��<�v�<���<�ȣ<�Q�<��<o=�<���<o�<���<#G�<���<�M�<I��<
<�nq<�*[<[ B<;{(<��<�
�;���;���;�7�;�) <��<�r<T%<�q&<�w<��<R��;y�;�M�;��T;�N-;֧);�"G;�@};[K�;/��;��;�B�;��<�-<�� <���;L��;'4�;�[�;{��;2Z�;�;��;�A�;�È;��W;�;3gC:koK�7���Om�"��_��4姻/8��%�{�rh@�_$��j������&�i7r�Yʨ���ڻ�P�O��X��Z�\���p ��C߻�����٣��摻&ى�����M葻Wɜ��꨻I���ѱ��,�ƻ'�ͻԻ��ܻ2黊f���@A��3��^J���_��Iq�*|��F~�O�w��i�bW��QD��4���+���+��4�knD�8X��k�={�m
��2��ٕ{��Sl���X��>D���0�� �e��Q���H�/I����c���������j���]�ڎ�����#�,1���C��?Y�P�o����7É� 썼���Ja��&��q��W_��MR�V�L�w�P���\�{#o����񷋼�Ԓ�����锼#���������{��g���U�ͮG��m>�I�9��8���9�%�;�6�=��8?�L#@���@�3�@��4B��E��4L��  �  ���<L�<<ӭ<�t�<�'�<G��<��<b�</؁<
�<�?�<�x�<dx�<#E�<���<��<p,�<%��<�&�<*E�<ʍs<��o<�u<�܁<�ڋ<#�<+�<U��<>Ȳ<�5�<�3�<!g�<���<�p�<�o�<z׵<���<�۵<V�<}J�<08�<W��<0�<��<=.�<��<�`v<�^c<I�W<�fU<��\<�l<,�<dr�<*ޒ<Q��<2��<��<��<�[~<͞h<U2W<VpM<bM<�V<�f<:�{<�<�-�<�o�<���<a��<�У<�?�<��<�Ɯ<��<fd�<')�<��<��<�Q�<&\�<��<��n<�:V<~�:<��<E�<z��;�&�;2��;W �;W��;PS<|�<8�<Q[ <d6<��<S��;�!�;��k;�;/��:��:�a;PVR;��;g�;���;u��;;A<�B<C� <-��;���;\b�;tB�;���;�	�;���;��;�P�;ɳ�;@�P;@�:iK�9�ۦ��'@��܏�&���s�Ļ]tû�"��\8���fc���*����w��zS@������溻������ �@;(���%��	��X
�"���Ȼ6����`���=���/������o'������F��݁��pȻ:�λtԻ�Hܻo�����c-�JH"�|:��>S�Mk�YX~�+���;��y�����u�rca�K�L�]�;���1��1��A;��wL��b�S�w�ba��`������j��g�w�) b�6�J��85�G#��x��� �{N�K�C.����{��?���!�@Q��e����q9$�!�3�*�H�c�`��Jy�����o�������Ŕ��܏��f���oz��g�D�X�S�F�V�P�c�D�w�S=���ڑ�Q���3���囼����	�}tm�NY��}I���>�/�9��e8�-�9�H<��>�%;@�pA��"A�%!A��B�UiE���L��  �  �`�<\:�<���<:��<U>�<�>�<��<~�z<@�~<iՅ<�]�<C�<�/�<#�<}�<�ۦ<מ<`�<%1�<%|<��n<i�j<��p<�X<5�<r��<�0�<��<�u�<��<)�<�\�<X�<`I�<�=�<X��<���<��<Fܵ<MB�<�#�<���<���<ϝ<���<	A�<�Mr<E�^<ЯR<�XP<V�W<:�g<��|<(��< ��<nv�<�q�<F��<N��<��z<bzd<?|R<�dH<;	H<_PQ<+Yb<�x<��< P�<O�<A��<d��<jã<�,�<���<|��<���<r+�<7��<U�<��<�B�<�8�<�ˀ<�bm<ZST<j8<�<yu <��;��;�y�;���;���;V�<��<�d<�,<��<d<c��;�ɠ;�tZ;%O;;|�:(W�:�';(�B;т�;���;���;�;�� <:$<�� <�G�;��;V��;�i�;
�;p�;@�;�m�;s�;A��;R�M;��:�d�9Q㾺ŁO�O꘻�㼻1�λ�<ͻ���߽��z�o��*5�������qI�!;���K��5M��Kx��%�F-���*��`�r��s���̻����h�������J��L���rt�����������A���ɻ�ϻ$�ԻV\ܻ�\黴���$�-�#�Rl<�?�V��"o�B�����������:��y���d��kO�x�=��%4�
4��=��MO��{e��{�k����������ʆ���{�~e��rM��6�*I$�w���4��-��i�M�w��g6�������JT��g��x��&���$�5��kJ��2c�_�|����"���BD���(���e��ӿ}���i��5[�S2U�!Y�tof���z���������S��� d���c��?䎼�}��5�o�L�Z��NJ��[?���9�@v8�u�9��^<�v�>��@�lA��jA��HA��%B�̄E�i�L��  �  ���<L�<<ӭ<�t�<�'�<G��<��<b�</؁<
�<�?�<�x�<dx�<#E�<���<��<p,�<%��<�&�<*E�<ʍs<��o<�u<�܁<�ڋ<#�<+�<U��<>Ȳ<�5�<�3�<!g�<���<�p�<�o�<z׵<���<�۵<V�<}J�<08�<W��<0�<��<=.�<��<�`v<�^c<I�W<�fU<��\<�l<,�<dr�<*ޒ<Q��<2��<��<��<�[~<͞h<U2W<VpM<bM<�V<�f<:�{<�<�-�<�o�<���<a��<�У<�?�<��<�Ɯ<��<kd�<-)�<��<��<�Q�<0\�<��<�n<;V<��:<ʣ<^�<���;�&�;Z��;z �;u��;\S<��<=�<R[ <a6<��<?��;�!�;��k;̚;���:�:-a;�UR;䤏;6�;x��;J��;'A<xB<4� <��;���;Sb�;sB�;���;�	�;ƚ�; ��;�P�;;��P;�@�:bN�96ۦ�9'@�[܏���H�Ļ6tûo"��@8���fc���*�|��w���S@������溻1��"���� �U;(���%��	��X
�9"�'�Ȼf����`��!>���/�������'�����F�����pȻD�λ
tԻ�Hܻr�����c-�JH"�|:��>S�Mk�YX~�*���;��x�����u�rca�K�L�]�;���1��1��A;��wL��b�S�w�ba��`������j��g�w�) b�6�J��85�G#��x��� �{N�K�C.����{��?���!�@Q��e����q9$�!�3�*�H�c�`��Jy�����o�������Ŕ��܏��f���oz��g�D�X�S�F�V�P�c�D�w�S=���ڑ�Q���3���囼����	�}tm�NY��}I���>�/�9��e8�-�9�H<��>�%;@�pA��"A�%!A��B�UiE���L��  �  p��<G��<"��<6��<�k�<?Ȑ<���<6+�<(��<tD�<ړ�<�ܟ<��<fo�<��<)A�<��<]�<���<嫆<f��<%�}<J��<��<ܐ<��<ж�<�&�<�q�<-Z�<� �<]�<���<�Ƿ<;�<�W�<��<_�<��< 5�<�:�<�\�<�+�<=��<�d�<�Z�<Ӏ<&vp<��e<U�c<:j<L�w<��<@��<BN�<ا�<!��<��<C�<��<�Tt<�{d<w�[<*P[<o]c<Mr<�b�<�F�<�c�<;��<�v�<���<�ȣ<�Q�<��<u=�<���<x�<���<1G�<��<�M�<\��<<�nq<+[<� B<j{(<��<�
�;A��;���;�7�;�) <��<s<T%<�q&<�w<��<+��;F�;DM�;,�T;BN-;'�);"G;�?};�J�;���;'�;�B�;y�<�-<o� <���;.��;4�;�[�;���;JZ�;9�;��;
B�;Ĉ;b�W;��;jC:wlK�z��Om��!�����䧻�7����{�h@�%$�kj�����*�&��7r��ʨ���ڻ�P�t�����Z����+q �QD߻鰾�0ڣ��摻wى�֩���葻�ɜ�먻q���𱾻D�ƻ9�ͻԻ��ܻ2黍f���@A��3��^J���_��Iq�*|��F~�O�w��i�bW��QD��4���+���+��4�knD�8X��k�={�m
��2��ٕ{��Sl���X��>D���0�� �e��Q���H�/I����c���������j���]�ڎ�����#�,1���C��?Y�P�o����7É� 썼���Ja��&��q��W_��MR�V�L�w�P���\�{#o����񷋼�Ԓ�����锼#���������{��g���U�ͮG��m>�I�9��8���9�%�;�6�=��8?�L#@���@�3�@��4B��E��4L��  �  ���<mU�<��<2�<%��<;��<�	�<2��<ؒ<$w�<�x�<m]�<�j�<���<{��<�<��<��<}�<��< �<�e�<�p�<���<×<�ڟ<K��<爮<���<;̶<H]�<Ǹ<υ�<���<�Z�<�ն<�p�<��<Ƅ�<|�<f��<�#�<?�<��<�y�<gf�<���<��<{Xz<Hlx<=�}<���<[��<K��<�Q�<��<V�<��<��<�]�<�ӂ<�x<mp<T�o<�tv<�+�<���<-��<�<$��<�g�<}�<E"�<��<~��<���<E�<X��<��<�:�<�<�<���<V�<|�<$t<�a<��K<�6<��!<@�<W<�<)�<��<j�<~�'<��.<�)/<�x'<5_<�<���;�_�;�o�;�+�;9/z;�Ƈ;F��;ד�;K�;��;X8�;B<�<���;ހ�;��;	��;P}�;���;��;�!�;~ �;pw�;*;�;�R[;B ;V��:[|�,	��Zr%�e�]���|���~���f��<�z��S�Ǻ�?������#���F������G���H��O��Fy�!��!���B����˻�ղ�ݘ��z����Y��[��]���띻|��%�� ��R�ŻP8λ zֻ��߻(@�<����
������+��[>�CP���^�:�g���i�5d��>X�;�H�{08�3�*��"���"�ɩ*���8�ΰI���Z���g��To�Huo��h��#\�_fL�C�;�M�+�������L�&���:����+��x������Z�' �{w�����m�"�3�.�1>���O�`*b��s�������u����h�r�@#c��S���H�8D�W�G��^R�mb���t�֦��ʈ�]���[ˊ�W�������Np��A`���Q�!�F��-?��5;���9�0>:�,k;���<��7>�NU?�/S@���A���C�iG��M��  �  ��<J��<n��<���<4L�<4x�<�L�<퇝<���<-�<��<��<�<�<���<3�<�߯<�֨<"w�<�<2Ӗ<�A�<�n�<�ޙ<�Ȟ<�Z�<@Щ<��<9%�<���<��<:��<pd�</�<Q�<��<3�<v?�<���<�a�<;�<dC�<�7�<��<]ݝ<P�<w�<-�<!<)�<�]�<[�<�0�<��<��<H�<t�<럠<W�<=ړ<��<�d�<o,�<��<7ȅ<�Љ<K�<_�<�O�<"0�<x��<�<��<Kw�<�;�<r|�<�F�<먘<竕<�S�<8��<���<O�<	s�<>�s<��d<�fT<�C<~@4<;�'<m%<�	<D><ҝ$< -<G�4<�9<��8<�|1<1$<��<Y��;�^�;���;߬�;�W�;�K�;���;���;�;���;���;-��;I�;K��;H�;�u�;T�;���;�[�;<Ͻ;VC�;y��;[��;DX~;�]R;��;,��:�]:����Y��:T�	��9!�W!�Ug�'Ϡ�РN�4���OL�&n��)x�ݣ]�6���浻!�λ�ܻ�8޻�׻��ɻ�,������m���o������ f���1���ע��Ū�ڪ���=��Qǻt�ѻ{�ܻԢ転�����U<����w�$�W�2�3�?���I�suP��Q�-M���C��B7�H)*��H���y+�щ���*���8��gF�wFQ��wW��X�M�S���J��@��R4�kX)��3 �i����Z�@m����/d�D��˴�W+��:����9��4`��&��/�/l:��XG�?�T���`�tXj��vo�t,o��ji�|P_�%�R�N�F�>�e�:���=�a}F�G�S���b�h-p�ATz�N^���~�]y��gp��e��Z�ӠP�z�H�=C�I�?�?�=���<�T�<�F)=�o>�&�?�N�A��D��bG�n�K�&FQ��  �  ���<c��<��<K�<eW�</ �<)�< �<1!�<�ܬ<�ݰ<�Y�<�S�<QԻ<�)�<��<�<_��<;�<��<�~�<���<��<���<t1�<�Ԧ<J��<>��<3�<=�<ϧ�<�L�<�Ǵ<ߵ<fV�<3�<��<��<(ɰ<�8�<��<�Ҩ<��<��<�<l�<�	�<W�<j̓<�ܓ<|��<�>�<�̝<���<h�<k��<�b�<��<4��<vG�<�<e��<��<�<�s�<�#�<wv�<���<2J�<�#�</y�<�c�<b��<mH�<a �<J�<n��<��<�P�<U�<'@�<(T�<Vd�<D�x<"�n<��c<�X<1"N<[+D<��;<�6<ߢ3< �4<G<8<>?=<лA<�C<��A<��:<�y/<�!<	�<�<<o�;f��;e	�;A��;r��;Q�;��;�.�;5�;�g�;���;��;�)�;���;���;M��;�H�;�ж;=2�;���;�};�=Z;�4;w�;���:��l:R�9�ڋ���8��z��W���an�3h'����r����_	��䄹!"I�4�Ⱥ= ���]�߻������Ү��ٵ�,���Ӵ�����Ԓ��򢩻sk��u�������VR���ĭ����������U�̻a�ڻ�"�ʤ��W]�Ų�t�Ʊ�]�"�z�*�,�1��F7�r:�FO:�ay6�jV/�_&�yu�^����T5������'��D2�d�:�|@�y�A�M@��n<��$7�I1��+���&�:""��8���������������;��7�`��O#���(�co.���4���;�	C�J��2Q�MBV�s�X�t�W�GS�G�K���B��I:�w4�2�1��74�'";��3E���P�t[��Gc��h�5Qi���g��c�S�^�RaY��aT�sP�d]L�I� �E���B�1�@��r?���?�R�A��.E�`�I��#O�
�T��}Z��  �  ��<QW�<>�<I;�<꠲<�N�<V�<<�<%(�<�4�<iڸ<m��<��<���<O��<� �<A�<�]�<DX�<D��<>��<�E�< ��<��<Bʦ<J�<��<*?�<��<�s�<���<�~�<c�<�Ʋ<��<��<0E�<�Q�<%��<���<�7�<�k�<�j�<[�<5/�<���<�V�<@]�<,˜<oӝ<���<2�<�?�<�N�<�ª<��<�ث<!�<J0�<3��<�؟<��<���<D�<ʖ<bԕ< �<���<��<N�<>�<p�<���<��<�\�<
��<���<��<���<��< ǅ<FL<�-t<�j<cc<+�\<osW<��R<��N<�K<]6I<��G<tH<>cI<�)K<�XL<�K<�lH<4�A<L�8<#J-<�!<�d<�<�t<�;�;�,�;	��;��;�B�;��;���;�[�;��;��;ǰ�;i��;L,�;9��;��;.��;+��;�u;d6G;1,;���:k�:�ޝ:�t:��6:��:*ɭ91 h9o�C9's9�}�9�A�9�7:��9��9S�����r�2�׺G���KJ�v�q�*>���j��9n������&i���Ժ�n��XYŻ6ǻ� ƻxû/ؿ�E��������ɻ��׻�n��L��#
��=����% ���#�I�&��@(��+)�%P)�y�(�kp&�D�"��z��5����;��	� Q	�t���O�Bi�� ��'�:
,�5}/�.�1��-3�~4�\f4��)4�H3�H�0��-�4�'���!�^��C��R�����G.���!��_)�#1��7���<�S�@�	C���D�	 F���F�ײF���E���C���?���:��5���/�I,�Y�*���,���1���8���@���H��JO��gT��
X���Z�Vp\�+�]��o^�v^��]�>O[�NuW�SR�	�L���G��`D�i�C�|F���K�'>S�<V[��c��wi��  �  s\�<� �<��<��<W��<�L�<%��<oֹ<I��<�M�<R�<�O�<�d�<?��<��<��<���<�P�<���<�߶<��<��<��<��<{�<�}�<x�<��<��<�z�<���<Kƥ<7U�<�8�<X�<%��<y:�<���<6��<�%�<���<`�<#�<Xj�<P�<틚<�d�<>�<Ӣ<��<��<q��<�Ԫ<Qx�<?��<�:�<���<9�<�4�<���<��< �<�N�<�X�<.��<GH�< p�<_͏<�ǌ<2ӊ</W�<�v�<�<r�<��<*��<�c�<��<CM�<BE�<��|<ʜm<D�`<�.W<�Q<�BO<�pO<@Q<HS<�CU<{�V<W<m�V<amV<ʂU<o�S<c�P<�L<��F<��><66<Q�,<r>#<��<Ch<��<��;��;@��;��;���;0�;y��;�c�;�̬;�A�;?�;���;x�;tS�;l��;�r;�T5;3��:5o�:��E:�*	:��9��:`�9:Ѓc:���:،:
��:+�:��:�ރ:�h:�3:+�9�t5�>���ֺĐ�e�7�M,^�C������".���û��ջZm�]R�~g�$�*l�I�ػ�\ѻ�iл�	ػU��p ����oZ�<�&���.�|	3�bj3���0�R�,��('���!�O��6 ������������W����������N
�ܑ��L�~:��g�#��k)�hf0��~7���=���B���E���D�m�@�[A9��0���&����b��F�b$�o-��s8�6C���K�k�P�UR�7�P�M�H���B�\S=�s�8�3�4�P1��-��*��Z(���&�;�&�8h(���+�-�/�3#5�w�:�tO@�GF���L�tT���[��@c���i���n�S�p��jo��{j�.�b���Y�_�Q��L�P�J�n�M�P�U��`�|k���u��}��  �  �ˡ<3~�<��<�:�<o��<�'�<p��<5��<�F�<h��<���<��<�*�<$��<�o�<��<+��<<Y�<�<��<S��<Y��<M`�<�2�<G��<v��<o�<n��<�o�<F��<��<���<_0�<���<�߫<�<^%�<ǐ�<i�<�T�<rb�<	��<Ÿ�<Yy�<`�<[��<�e�<��<Z��<BL�<ǫ<�[�<-U�<��<6,�<�'�<��<sZ�<Ή�<�f�<�۪<���<��<6r�<��<���<��<x�<V#�<�g<Fz}<0Z�<&�<)�<�<m��<��<�(�<��<�~<�k<OY<�$J<�@<�;<~�<<q
B<\hI<�bQ< yX<]<D$`<d`<��^<��[<�X<��S<�GN<wyH<�)B<�[;<�4<�,<��"<�><$p<�N�;�>�;�;�ɛ;&p�;kl;Lpd;�wq;�;b_�;���;���;��;�w�;$�~;�J7;k��:�d:q�E�7)�]>D���uV��l�9��`:��:	D�:��:��:*�:�:��:�TS:f��9���8�����H9��Θ� ~ۺ�j�g�B�K�y�%��� ��ϒݻ�S�����2���#�
��;�G���>軮]�]8� T��B%��>�%)/�A?=�J{F�D�I��lG�|k@��v6�&=+��J ���������
��:�����������K�52������s�
�}�����*���t'�j�3��@�J�L�tsV��\��L\�*W��:M���@��,4��T*�
�%��&'�"�.�	X;���I���W��Xb��h�(Gh��]c�k�Z�J�O�l�D��P:���1��+��(���%���$��+$�^$�4 %��f&��6(���*���-�ɪ1���6��G>��G���S��`��cn��jz�W����胼�\��a!���u��Ui���]�_�U�bnS�ЇW��ka��&o�N	~�h���*b���  �  N�<,K�<]�<͢<0Ī<Ҵ�<���<���<�e�<� �<p��<�Z�<���<��<a�<���<�`�<s��<ϳ�<c̽<��<���<S��<s7�<+�<d�<�c�<�?�<i|�<	h�<	��<��<��<J��<��<yH�<D��<��<�M�<?�<m6�<d�<��}<<9l�<=�<�Q�<kD�<���<y�<��<$��<�
�<��<�<~(�<�ݮ<���<�{�<��<{�<� �<yk�<��<���<��<`��<��<~:q<�'h<v�e<gVj<�Zt<h��<m��<�R�<)c�<w_�<0k�<$q<�Z<��D<�j3<Em(<��$<��(<��1<P
><K<�V<�T_<d<�e<�c<��^<��Y<��S<?.N<�H<�C<ǜ=<#�7<�z0<�5'<x�<�<cM�;�s�;W?�;��k;��/;<�;��;V�;��A;�,r;���;��; �;�+�;>�M;���:q:	�7��%Ӻ]���	
�1KẴl���|��:���:|��:�/�:GU�:�w�:���:�I�:2T:���9� 9�Y�����t�-���h���;��(��J��sqӻU����m�#��G&�^A&�����M��	�� �;���Y���̦	�����.���B�|�S�!c^�x~a�#]��kR���C��x3�A�#��T��a�J��������R�L���Y�������ɉ��f�	S
��L�c���W*�\;�S\M�f:^�ͥk��ns��$t�7�m��<a��Q���A��Y5��B/��1��m:��I��\[�aXl�Uy�w ���Z���w�J!k�:z[�|+K��@<�tI0�(�i#��!���!�x�"�h�#�L:%�}K&�R5'��G(��*�$-��2�(};��H�X��Aj��|�����Č�=ʏ��(������Y��f�x�`j��7`�]���a��m��o~�mR���r������  �  s�<TL�<z�<q��<E|�<�\�<��<���<���<H��<@�<2��<��<��<��<~�<�U�<��<pd�<��<��<��<X��<#t�<K�<�h�<%7�<�0z<�v<��z<,��<TH�<��<���<�d�<Z�<o�<�7�<BE�<��<2u<��j<7(i<�	p<S~<�m�< ��<���<Y֤<��<Q��<.S�<���<M�<�P�<ﱮ<1d�<�i�<��<5��<�ͭ<٭�< ��<��<B�<��<�M�<_o<�1^<	�S<�>Q<�W<�`c<~s<1,�<���<(�<"
�<��z<��d<�K<�i3<��<�<2�<�4<�Q"<2K2<7C<exR<�^<^�d<c�f<"�d<��_<
�Y<�XS<m0M<��G<ĺB<�><��8<��1<�,(<�b<�<3��;	�;�;�%;{��:j>d:ɑO:�w�:�� ;?b<;%jq;�f�;�Շ;E�i;�^#;J3�:�I���rE:���[��Y��07�����f��&9��:^��:Up;ɿ;�x�:j��:S��:�xE:�9QÐ8vvi����&_a��D���b��
A�g��٠�����F>�Z�#��3��E;��e:��2���$�8I�q�
�������a��$&��<���S�
g�"s��Ov��p��8c�' Q���<��?)�X��kk�����Y�?� ����u�����Q�p�e��|��B��[	��b��4n/�,D�Z�{�n���~��
��Vn��*����cr���_�jtM��?��8���9�݋D���U�j]j��~�����kj���剼y<����z�Zg�S�l�@�w�1�1�'���!�d. �+� �#�"�P�$�H8&��)'�ʊ'�W�'��(��+�W�1���;�SK�`^��at�9\��{T���Y5���_��Po���y��e8��(\u�K�i���e���j�gyx��˅�K������pE���  �  �M�<�b�<�ь<�b�<���<۞�<�b�<*ݽ<���< ��<O�<U��<�L�<\&�<�_�<��<��<l�<x�<��<>��<(��<|Ǫ<�q�<�	�<��<ٗy<�-l<]�g<�7m<C {<E�<H`�<��<�E�<`ߟ<T��<US�<x��<q�z<B'h<�\<��Z<��b<�Er<���<�#�<*-�<�<2`�<m��<�h�<���<��<��<�5�<��<��<�c�<���<��<���<��<ş<f�<�$�<R{<r�c<o�P<��E<�2C<)�I<��W<)�i<{�z<aD�<	 �<��<�)t<��\<B�A<:�'<*q<ɩ<��<J	<A<#�)<C�<<��N<�\<3d<�f<#�d<��_<5WY<��R</L<��F<�
B<W�=<D�8<� 2<��'<��<�<��;���;�ZW;FH�:��%:,�i�@x��A�9�ĩ:�;��S;�-w;��w;��P;�S;��:�͏�i)�V7q�O]��zF����h��n'�������6���]:���:�� ;X4;=L�:_��:�h�:��5:;y�9�*57�㈹ߘ
�˩`��î�3D��I������û8����:��0�`�A���I�uH�lL>��3/���L��eQ����z�T.���F�Ni_��+t�j����M���~�Yo��Z�D�C�j�-�vV�ދ� ��2��� � ��8��p��O�}��~�������	�7��q ���3�K��pc��7z�I���$������"����}��i�NhU�'�E�'&>��@�zK��&^��|t�x���P������𐼮���A�$p�iY�C�D���3�>(��!�V ��� �3#�4s%��9'�X(�4(��(�w�(��y+���1�@Q=�N���c�|�_n���v��ć���Y���T��L˚��������|�p�o���k� Wq����<��׬��n���.���  �  &`Z;Ҵz;;��;���;[#<q\M<;fs<�3�<�}�<���<.��<��<�Q�<1��<�l�<���<�؞<?�<��<f�<-%�<�x{<�bX<��.<�.<�;�N;qd�:��:��;�Aj;rB�;x�<�!<��4<e�7<��)<~^<,�;Y��;�;��P:�:+��:E
S;ݞ�;�<+�/<�9T<�q<w��<2�<�]�<���<4 �<��<���<�^�<��<�<6��<4�<�m<J�P<��+<�� <���;�A-;&;1:a��`��[�9g;V��;�d�;)��;d�<'��;���;wr�;e9�:�R����\�Π��B���rs��� ��`�9� 0;:��;ҍ�;�k<7�<T�<L<��<�<g�
<r�<��;`W�;'V�;���;"J�;��B;�#P:���������77$��wB��Q��wO�d�=�5� �`^���»���.���w�����\��b.G�B�n�޴�������}��~��F]��`6�3��8׻���`yp�-�D�545�;�9��I��1_��v�^��������Y��ͭ����ػ���!�4}G��1t����:���Ee��Z�ɼ��μ�g˼���&t���4��1ܓ������>��v3���"���P��ϼ�e༏�IQ��漺�ؼ:�żOV���|���&��:u���`���S���L�>�I���H���H��*I���I�p�J�>,N�F"U�e�a��sv�ʸ��=+��oe���sǼM�ۼZv뼶���I���
+ݼֹʼ裸�򨪼'����������ʜ����Ѽ�传<�ف��=7�����z߼;V˼���e���3���i����w�f�m��Fi��h�wh��di���j��%l�"�n���s��2}�T��������ע����~�̼���vK��$��.�1��Js���4�)�ڼ7�ɼ ����!Z��·ʼi7ܼ��� �<,��  �  �d};)K�;5J�;zN <CK(<|�P<Xtu<䫉<B��<㓛<Z`�< �<^)�<-ؠ<`O�<z��<1��<�
�<��<L�<�K�<��|<z�Z<E�2<`u<E��;�An;ф;l��:kS%;�@�;zE�;�<G{&<�8<k�;<;.<-a<�2�;庐;m)#;$��:#��:�K;�-p;���;u{
<��2<��U<B�q<ϸ�<��<�&�<ހ�<�ڍ<,ύ<��<n:�<B�<@׊<�\�<��<:n<["R<Ud.<�1<nz�;��I;۾�:�8���V:��;�ґ;k��;,( <+�	<�O<y�;���;4��:�M^�	�;�HE��놻��S���ʺ�!:u�?;��;1�;��<@�<�o<��<k<�l<$�
<-�<	M�;���;D��;�k�;���;��E;0*o:vhҺ�!��dv�l���:���H�=�F���5������/��fΓ��f���K��t޻���v@��!g�#z��o����E���av���V�gu1�Ո��!ӻ�'��;�o�,�E���6�;;�� K��`��mw�I��bQ������f���ٻ[c����GE�fp��L��˙���p���Fż,Yʼ�3Ǽ��.���x�����������B��e�������J���y˼d[ܼ���@��
��ռ��¼)������R��J�t�-�`�e�S��-M�j6J�	EI�'I��fI�m J��[K�h�N��U��b�#�u�"���vŚ�vC����ļ.ؼ�`缢�＀��)���ټ~�Ǽ����}����������[������μ	
Ἑ��$�����e�뼈ܼa�ȼ����Ԡ�d���79���w��(n�;�i��ph���h��i�e�j�>tl��o�2%t��}�����-��j⡼����lʼ��߼u��|������"�����C��:�׼�^Ǽ����L���4L���*ȼ`cټ��X �����  �  ���;X��;���;H�<�5<~�Y<�Pz<��<XT�<�Ú<`i�<0�<*��<]�<��<��<��<�%�<��<��<�?�<��~<�j`<a<<��<[��;���;5�u;D�^;��;w�;��;Q<Jc3<�ZD<��F<�:<E� <wC�;���;$<~;m>8;��,;\�];�`�;���;�<<�:<��Y<��r<<�<F��<�3�<c��<E�<�[�<R'�<��<���<�<�m�<��<"�n<nU<�W5<�f<���;:�;j�';#�:�B�:�8;�q;9C�;��;�B<h�<�n<x�;ۻ�;�p6;���9μ���$��-��X���%ѹ�:ϋh;r��;�*�;��<-O<Px<��<��<|Z<��	<ް<��;3[�;$��;�)�;�Z�;��K;�ԛ:��k�+ǻ���=z"��0�
�.� ��nA��һdԝ��x�1�l��%��o�û���{u-��BQ��k��v��r��3a�?\E��D$�ʼ�Wyɻ�י���q�4[L��>���A���O��c�r�z������ݗ�[g��_����ۻXZ�Sz�AP?��f�#���P��	o���2��L����S��2��ꤼ����p���ń�������v��`���2_����мޏڼ�ܼx׼'�ʼ����h7��D���u����s�s�a���U�bO��K��mJ�J�%GJ��K�e�L�TxP�6XW��'c�EPu�xK��F�����.���xNμ7�ۼ��ӷ�1~ܼ�Tϼ����`ٮ��Y�����&[������j��ѻż�ּ�]㼕�鼒�輢�༒�ҼP@�����ŝ�?���)��:+y��p�f�k�
�i�|�i��|j�E�k���m���p��v��1�r߆�<|������谼5ļ7׼-�F6������B����c�P�'�ϼ��������u��z���y���_Ѽ�㼘����  �  �%�;�-<��<�&*<D�F<ed<ؤ~<�I�<���<�C�<zܛ<��<Z�<z+�<�Ҟ<Mٝ<�>�<�ߙ<�\�<�*�<���<i<�f<�WH<ţ(<�%
<���;���;H��;c��;�g�;��<xY.<v�F<�9U<FCW<	L<��5<)o<J��;�w�;ۣ;���;��;n�;�u<WF%<�gB<N#\<7�p<C!�<
f�<W��<���<�ϋ<3>�<�<�?�<�ʉ<�w�<0҃<@�|<P�l<�bW<A�<<��<��;�q�;8�;x\t;Vn;�>�;���;�c�;�F<�+<��$<x�<�	<��;N�;'�; ,:g��}Z��RS8���:�T1;�r�;�о;���;��<��<�-<�<oI<u�<N�<Pe<��;��;���;J=�;>�;��H;U�:�t �9:(��ۗ��Ի<n ������<����һz���%�j��'3�+�K�Y�z`��M�ܻ�C���0���G���R���P��$C��5-�;��F�������К���V\`���R��S�̟\���l�~3�������p������ǻ����&������9�X`Z��,}��e������Z���֫�\ʩ��B��&&��1��`���xx���z�����Nؑ������a��W���ȼY�ʼ�nƼü����!���z��'��Yu���e��Z��S�/�O�*SM�UAL��sL���M��P�YLU���\�܉g��Yw�pI���x��f�����~q��ך˼	�ѼӺѼ>|˼�,��2������@��jғ�����朜�O9��R����ƼNҼ��׼�5׼��мreż�c��H���#�����P�����}�m@u�)p��zm��gl��l�(n�!�p�'�t�{��!��fĈ�A쑼�ʝ�o
��O����s˼Fټ�:�Ĭ�/���ݼW�Ѽ7rüDm���`��GF��$ݭ������wż��Լؾ��k��  �  �^%<��'<^2<.C<SW<jlk<T~<�D�<�Ѝ<��<�Ɩ<���<J��<���<R��<�8�<>ɘ<�j�<�'�<�ۋ<�I�<0sz<�>g<�Q<'�:<��$<�<��<bA<�q<�L<�1<)+I<��\<�h<�Yj<E�`<tMN<�'6<�O<�<���;_b�;���;��
<��<`2<�G<�Y<�qi<w"v<�<��<ц<�ڈ<��<��<�`�<���<ڱ�<��|<�=r<F�d<�-T<x�@<w�*<y�<1$�;�C�;���;��;�
�;�3�;�<  %<R3<ܗ7<i�0<�N<�V<���;�y�;�K;"�;���:�.;X�<;�|;�e�;@��;\��;�s�;}�<8�<)�<�	<C<�&<�;[K�;��;8�;�;޾y;�D/;�C�:���?�ֺ�-O��Ǔ�®���Ż�û���]���S�P�3���ĺ���G4
��{\�����]�]�^�M�)�Mu*��"��e���H=⻦���������Ʂ�td{�ͳt�T*v�����㉻ש���«��Z»p#ܻҒ������~!�X8�;�P�J�j�1ၼ�{���ߓ�G���8c����������VM{�l���d�CJg�j�t��c��j���ɠ��K���ĳ�M��yﳼ���k����������Z��H�|���o�ؗe���]�|�W��6S�W�P��Q�ӤS�
OX���^��/g���q�)3��ه������q�����Ӱ���x��툽�����9���^g���袼��������;���E��ꡑ�k������\���;罼�üUü�'��݆��ح����ٟ��I󐼕ω�U1������Hy�ѝt�r�q�*,q���r��w�=}�$�����������0���Q��Tר��4��Gs���Fɼ�=м\Ӽ91Ѽ��ʼ\����,��Ó��4:��2Ơ�Oף����|��/=ļٸϼ^�׼�  �  Q�M<,�K<]zO<H�V<��`<�3k<z�u<��<K�<׻�<�f�<Გ<�.�<oE�<�z�<��<�<��<���<ڣ�<�:y<��l<MR`<nnS<�F<&
;<�1<u-<�-<��4<U�A<̀R<B;d<�Bs<�F|<�9}<"�u<�g<d;T<o�@<p�/<xM$<��<E�<�#%<?.<ݥ8<��C<��N<zqY<��c<n<J�w<�_�<Eσ<���<r��<t�<=i<��u<�
k<��_<DST<�zH<�3<<��/<5#<<:�<!�<K�<��<3!<e0<><��G<�J<q�C<��4<=_<��<W��;�;�;u��;J?�;�;0#�;�#�;�զ;]��;r�;���;Y�;P��;���;2�;���;u��;���; 6�;�;�v�;�q;�2;?-�:�S:�U#�d	���r��D6���Z�U	k���c�$�D������!�4�6?��fP��_m�Y ��Z�q��p�ɻ��f�����Ǡ�+� ������⻜ ӻ�bĻ�ζ��T��y"��������MS�������n���;»��޻U���Y������.���>���N���^�Upm�5�y����}���W���vy��m�X�_�VpU�z�P��T�i�_�B�q��܃�����|��D6��U���z͢��X�����PᖼR��ŋ��V�����ܐw�,|m��`d�gF]�WY�>bY��u]���d�8an��y����ʇ�8���l���'ݙ�m؟�f��wʨ�B$��R���)ˣ��o��i���'Ԋ����ƿ����������َ����
��uǩ������g��BG��	����J��������Ah���W���i��~���D��N>��g+{�[y��{�p����f��ϊ�
���\���پ������v����J��@0��|���+��Rü��S��L������k����#��Gb���㙼�G��n\��"c�������ü�  �  >]o<��h<0d<V�a<�n`<&�`<��b<@g<��n<K�x<�y�<ˈ<t=�<��<�H�<�ҏ<���<��<;mx<>j<`R^<AU<� O<QK<?�H<`H<��H<z:K<�XP<h]X<bc<y�o<�[|<]w�<���<>ʆ<��<M}<M+o<f`<��R<f�G<ff?<��9< �6<�5<��4<�(6<O�9<�?<�H<T<<Pa<cPn<�x<y�~<}�~<�fx<�gm<��_<RUQ<�sD<~:<}2<~-<x*<��(<�K(<#)<=�+<�i0<{�7<�@<�K<�,T<��Y<Z<L�S<��G<�w6<��"<�Q<�%�;�u�;).�;s��;�ʧ;N�;P��;��;�;b��; ��;NY�;���;L��;.��;��;'��;�f�;-��;��S;�;�}�:Z�9L�˹
_�������8�ͺ-VԺ��ɺ8����l��K͹�y9�:.GP:�{,:^9��:��캇C��f�������j���Ի�F�%����sL���T��N����L��߻v�λ+|��U/��"R��.��LŻ!�⻤���2�o)�dI9�0�E���O���V��+\�L,`��b�(�c�iOb�$G^���W�[�O�yG�InA���?�	pC��
M��h[�ޅl�B~�R���4o��ZE������ă��3���������V���=��Ƨ��a�������v��l��f���e�^�k�K�v��?��X�������┼	��������Y���񜼐᜼%
��)%���ꖼ/B��k]��rЅ��$�ƚu��q�Εr�8z�����M������&���C������q���䤼	���٥��ݤ���������J���������{ˈ�����;䂼�P��&���������ݝ��C��0M���欼�A��쩰�Z���Z���{���r��� ���$���/���י�?-��Y���?��x:�����+����G��݉��b����  �  ��<�'{<&1n<�Ba<�8U<�qK<n�E<9E<SK<��V<��f<��x<��<��<%�<���<�
�<�fm<FtY<�G<�:<4<Ye3<�7<R@<J<�T<�^_<��i<�s<s}<�p�<,��<� �<�	�<��<F��<�7�<�M�<F�y<n<�>b<7:V<��I<DX=<B1<� &<�<"j<$�<6%<�Q3<��D<B�V<X�e<��m<�n<[�e<8�V<��C<;�0<�:!<��<�<3O<}x<Xs#<͢-<��7<��A<�sJ<q�R<< Z<��`<e<V�g<�&f<f4`<V<��H<�>9<��(<�<�<�6�;�E�;��;�u�;Nf;I�<;r ';f4);bC;�p;�;��;z��;`f�;��;�֋;��?;9ӽ:[�R8�����s����2���p)ź�D���y
��-��>��9��C:��:U��:Q��:��:T;�:Jw:5�9`%�o�ǺЫ"�ņa�����P���λ	�� J����Y����E?����(Q�@ﻵ�ػ�Uͻ�һ/��$Z�>�i�5��K��\\���f�0�j�C�i� �d�i�]��lV�VHO���H�ԭB�-=��8��4���1�(b2�i�6�`�>���I���V���d��or�������s��n��Vp��������Fܥ�'���UH��e���)�����/�n�v�pv���~�_Ɇ��"�� ���`Q��1q��0t��턧��E��~�����������	��C���K����:� �u��cm��Fg���d���e�sk��ws��}������m���j������@✼3H��2j��w���#B���Y��Uf���^��-ؤ��	��2���~���|���Ό�Y����F��^=������A���{���ѻ�y^���۶�R!���䬼=���;z��с��������������������>��є������f����@���$��*0���  �  �<Ӭ�<��m<#W<��@<�-<[%!<�<�b"<��0<ՕE<��\<�q<__~<���<5�y<h<~=P<?�6<r� <��<�N<�7<�9<m�-<(B<�V<e(i<�y<o߂<�Ӈ<���<rn�<H_�<S�<��<���<<�<�ى<��<�9�<�&s<��b<v|O<��9<�f#<�w<���;֞�;,��;d'�;�<�[%<��<<e�O<�Z<��Z<�OP<k�<<w�$<\�<���;���;��;=o�;�<�t<��(<vN<<�9M<ϽZ<��d<��k<��o<�{q<��p<��m<�5h<��_<]@U<��H<S�:<�V*<�|<��<d&�;�Z�;�hW;*�:2�F:�9�!�8~:�V�:Xp.;�Vu;L/�;���;��;E�=;1�:���$���>h�׌�٦���u���S�������U2�� vL:�:���:��;Sm;��;ݵ;�m�:�q�:�?q:J��9���)������g��V����ϻ9�"���8/�z>�VpE�C���7��&���Z3�S���)�����a��H:���W��r��l������Ն�`z��p�v�łe�fhT��;E�\9��T0���*��w'��T&���&��~)�*&.���4�n=��wG��R���_�F�n�Q^��}������4��cɫ�9!��߸�����R���p���~���i���䄼.����������j���>���I@���ຼ�����������h��Q-�����cw��%�v��vm��Of��a�̒]��@\�P^]���`��kf���m�?w�)R��܅��pJ��ₛ���������	��aü�	Ǽ��ż����h���쪼��ݗ��x�����cޝ�|�������Px��LIʼֹμ
XμЙɼ����oҷ���V����Ĕ��s��f���_��3>����������#��gm�������Ϗ�S���0U���  �  ���<���<Tf<nF<�Z'<��<���;i-�;���;\�
<M�$<��@<=Z< rj<.|n<q(e<�P<�g3<߻<0K�;�Q�;���;�;nB�;{I<�3<"�P<��j<e�<�ɇ<�1�<���<z��<�w�<羓<6h�<�r�<�ې<�v�<�ي<@w�<�{<�f<�M<10/<u�<Ў�;��;v��;Y��;ک;���;"$<�"<�2:<�oG<&�G<��:<t#<�<���;�բ;]��;@N�; R�;6��;�m�;�< �8<DtP<ߋb<m�n<l�u<l�x<|�x<UGv<�9r<��l<ioe<s�\<�IR<�E<`4<\k<k�<R��;��;�l�:�#���Ǻ����"��C���#�p�`:87;�4Q;�&a;)�;;0a�:��ƹ��$�=����,Ż1j߻l�߻d�ǻ�S��#_U���Ӻ?����Ȑ:�;_�%;pe6;�8;&�0;,";n�;���:�(�:[�I:Z"�8�"@����!Q��˟�g�߻��.n3��}P�lMe���n�R�k���]�6�G�/�����`��,��5�c�V�ƻy�y4���㖼 k��ֈ��x!��I놼�s��Z�U�C��2��E&�G���E�?��P� �d$�!Q)��5/�6�	>��H�� U��_f��~|���������謁�ӹ�P�ż��̼��ͼ�_ȼ̗����������I������PV��4���0S���﮼�����)ɼ��ϼ��ϼ��ɼ�'��}=���7��Kԓ��V����z�'|l���b�J�\�֌Y���W�ϢW��X�t�Z�^���c�ySl�Y�x�鄼�:�����{��<��m˼�ּ sۼ�ڼ��Ӽ�Ǽ����(��;������ o���'��g���_�żD$Լ��޼�t�4��G�ڼ��μ���3ﱼzZ������p<��) ���7�������ւ��v��������� !���`���������������  �  ��<^�~<�D[<��4<��<�}�;;�;��;ze�;ZC�;:~<�m)<�jF<QY<#^<ϛS<g�;<3�<�D�;\	�;��;�;};js�;���;�C�;�I#<�.G<p%g<)n�<༉<���<��<���<d �<��<"z�<�Ǔ<���<�ϐ<rr�<KƇ<X~<٭e<NqF<"<�e�;�;{j;�M$;��;��I;���;�!�;H�<؋'<��6<{&7<�(<��<��;|�;��<;� ; R ;_>:;ؑ;�j�;��<g`1<��N<�d<�s<��z<}X}<�%|<3�x<�t<��n<Ah<ǌ`<��V<��I<]�7<0�<X� <1Զ;.�H;�N:���2j��Q��+�~����2���}:Q�	;w;c��:�\�9	��ES��.4ӻ�{�
���w���� �л������I<�HR�:��;�?9;�K;`�J;�d>;��+;�;�s�:<��:�Ά:��9n$�,�Ӻ��P�P���p����#��#L��	o�샼Ԃ��
���~��c���F�|�-������a�-�/�I�Jo�LH����������\D��5M��i����d��񁼄Rc���F���0��2"��`���g���>���!�8�&��Z,��,2�F*9��B��^P���c���}���5����𴼣%Ǽ�ռ�l޼��߼&�ټ
ͼѼ��+������X喼�����֝�N-��������̼@ڼJ�Ἴ���<ڼ��̼L����'��[u��I6��%�x�wh���]�wX���U��,U�9xU��_V�m�W�iwZ�u_�3.g�(�t�+�������\��S6��pȼ��ټ#��^�v켃K伓�ּ�)Ƽ����^ ���4���証�ϲ��¼��Ӽ8�4&�����O�꼸xۼO�ɼE���������𨎼ɱ������ก�� ���7��l����f���z���/���!��������  �  *�<Еy<�0R<I)'<���;���;%J�;YW[;h+y;r��;" �;s�</(9</�M<YS<d�G<u�-<RS
<�	�;D�;4=3;��;�CE;�8�;�{�;��<�?<��b<��<��<y��<��<Sg�<坕<%[�<��<�P�<�k�<պ�<�d�<l�<��}<��b<@<��<.t�;Dڈ;�{;�m�:��Z:
��:�NY;yX�;�k�;��<j|+<��+<B&<)1�;I�;IvV;�j�:<�9���9���:`BU;iW�;��<�*<�DK<��c<%t<V�|<�<�~}<�y<��t<�Ao<�i<��a<��X<�K<>�8<ߏ<�/�;�:�;V;,O�&eG�����Eǻj�ɻ�㬻�	p�}����8d�:��:�$�:�;�@�2�\��� ���"�D,�;`*�����/��V}��T>��%I���|:��;�R?;�R;�Q;��C;{�/;�L;�b;���:��:VH	:{1��M5Ѻ�jX�ܖ�����`1��^��A��ُ��ٕ�9�������v��nV�+�:��*�>�)��A9�S�W�bv�2������j����|��������Vƚ��!��NYk��K���1��X!������c��F���� ���%��)+�R�0�^97�+�@�P�N�l�c��'����������d���м9��ߊ�O��A�1�׼O�ż�����㤼����Z5������{����ļ�׼���������Ǒ���ּ�hüʩ��'ؚ��ɉ�p#y���f�n�[�=V��AT�<T�1�T��wU�e�V�p�X�Z#]�/fe��s�3������3���6����м0��\����u�����B���μP����"��P«�����~R���ɼ��ܼ ������ ��M��B�������мY������o%��ԏ����,���oր��q��궀��<���遼�т�FR���*���T��{����  �  :��<�uw<�N<�#"<0��;=3�;��^;AS8;(PW;�(�;���;�<�y4<"�I<�O<�C<H)<3~<�,�;�j;��;3��:-�#;D�;+�;r<�;<�a<V�~<�<�Ð<C�<���<�ĕ<Kz�<��<�s�<:��<H�<���<?~�<Fv}<�a<I�=<�<�e�;Z�u;L��:"�:�I�9q��:��;;㳦;��;�<��'<;�'<��<���;���;{K9;��}:����BD��Z8{:��8;R�;�Y�;�'<��I<Lrc<�2t<��|<�n<1�}<K�y<t�t<�oo<zXi<yJb<Y<��K<e�8<��<���;_�;w;�Zb��d��^���ػ�/ۻ*���/���&�ǗL�ic�:��:ݧg:�{>��H�s��M��~�%�{�4���2�_ ��8��յ���L��?m��qk:C�;'<@;vT;`=S;E;d�0;/(;�P;( �:P �::��9�Һ�}\��㷻lf��j6���d��������;��Wԗ��ύ��U}��\��?��.�lp-��e=��Y\�˞��q��h���%ٸ��Խ�M��⫮�e؝��t����n���L��2��_!�R/�Ώ�?a����� �K�%���*�U60�[�6�&G@�R�N��:d��΀��X�����q%��%ԼM���i�b�b<ۼ��ȼgA�����܃��/���5�������Ǽ`�ڼ����?��'򼽡�k*ڼ�AƼ���4��y�����y��f�vf[�&�U�"�S���S�,\T�Z:U�'nV�D}X�]�\��e���s� ��zt�������x����Ӽ	�缼���������� ������ѼH���A�����@�������@�̼Y8��� �����������I|ӼjX���ܪ�g���б��dՆ��x��c����G��ѕ��o��gɁ�������a���4��Yٔ��  �  *�<Еy<�0R<I)'<���;���;%J�;YW[;h+y;r��;" �;s�</(9</�M<YS<d�G<u�-<RS
<�	�;D�;4=3;��;�CE;�8�;�{�;��<�?<��b<��<��<y��<��<Sg�<坕<%[�<��<�P�<�k�<պ�<�d�<l�<��}<��b<@<��<.t�;Dڈ;�{;�m�:��Z:
��:�NY;yX�;�k�;��<j|+<��+<B&<)1�;I�;IvV;�j�:�;�9���9���:_BU;iW�;��<�*<�DK<��c<%t<Y�|<�<�~}<�y<�t<�Ao<i<��a<ϴX<#�K<W�8<��<�/�;;�;zV;EM��dG�ֲ���Eǻ9�ɻ�㬻L	p��|���8�d�:��:�$�:�<�p�2�-\��� ���"�)D,�W`*����0���}���>�Q'I�+�|:O�;WR?;��R;�Q;��C;f�/;�L;c;ӡ�:;�:TI	:/���4Ѻ]jX�������� `1��^��A��ُ��ٕ�-����󉼮�v��nV�"�:��*�=�)��A9�\�W�ov�;������v����|�������eƚ�"��lYk�K���1��X!�����t��T���� ���%��)+�W�0�b97�.�@�R�N�m�c��'����������d���м9��ߊ�O��A�1�׼O�ż�����㤼����Z5������{����ļ�׼���������Ǒ���ּ�hüʩ��'ؚ��ɉ�p#y���f�n�[�=V��AT�<T�1�T��wU�e�V�p�X�Z#]�/fe��s�3������3���6����м0��\����u�����B���μP����"��P«�����~R���ɼ��ܼ ������ ��M��B�������мY������o%��ԏ����,���oր��q��궀��<���遼�т�FR���*���T��{����  �  ��<^�~<�D[<��4<��<�}�;;�;��;ze�;ZC�;:~<�m)<�jF<QY<#^<ϛS<g�;<3�<�D�;\	�;��;�;};js�;���;�C�;�I#<�.G<p%g<)n�<༉<���<��<���<d �<��<"z�<�Ǔ<���<�ϐ<rr�<KƇ<X~<٭e<NqF<"<�e�;�;{j;�M$;��;��I;���;�!�;H�<؋'<��6<{&7<�(<��<��;|�;��<;� ;�Q ;^>:;ؑ;�j�;��<g`1<��N<�d<s<��z<�X}<�%|<A�x<�t<��n<]h<�`<��V<	�I<��7<d�<�� <�Զ;�H;�R:��2j�+� ����~����2���}:~�	;!w;2��:�Z�9ÿ麃S��{4ӻ|�<��-x����v�л0�����:C乪P�:	�;�>9;KK;��J;�d>;��+;�;�s�:���:�φ:���9��ʣӺ#�P��O��:p��Z�#��#L��	o��냼����󡇼�~�ɼc���F�j�-������j�-�@�I�co�]H��͡�����vD��QM������e��)񁼿Rc���F���0��2"��`������>���!�K�&��Z,��,2�N*9��B��^P���c���}���5����𴼣%Ǽ�ռ�l޼��߼&�ټ	ͼѼ��+������X喼�����֝�N-��������̼@ڼJ�Ἴ���<ڼ��̼L����'��[u��I6��%�x�wh���]�wX���U��,U�9xU��_V�m�W�iwZ�u_�3.g�(�t�+�������\��S6��pȼ��ټ#��^�v켃K伓�ּ�)Ƽ����^ ���4���証�ϲ��¼��Ӽ8�4&�����O�꼸xۼO�ɼE���������𨎼ɱ������ก�� ���7��l����f���z���/���!��������  �  ���<���<Tf<nF<�Z'<��<���;i-�;���;\�
<M�$<��@<=Z< rj<.|n<q(e<�P<�g3<߻<0K�;�Q�;���;�;nB�;{I<�3<"�P<��j<e�<�ɇ<�1�<���<z��<�w�<羓<6h�<�r�<�ې<�v�<�ي<@w�<�{<�f<�M<10/<u�<Ў�;��;v��;Y��;ک;���;"$<�"<�2:<�oG<&�G<��:<t#<�<���;�բ;]��;?N�;R�;6��;�m�;�< �8<EtP<�b<q�n<s�u<w�x<��x<iGv<:r<��l<�oe<��\<�IR<*E<�4<�k<��<��;%��;-o�:��x�Ǻ����"��A�½#�ޟ`:�7;>5Q;�&a;�;;�`�:��ƹ_�$�����-Ż�j߻�߻�ǻfT��p`U�3�Ӻ�
��]Ɛ:�;w�%;�d6;K�8;��0;�+";c�;@��:�)�:f�I:.8�8_@���� Q�Z˟�Ǌ߻����m3�<}P�Me�f�n��k�Ļ]��G��/������`��,�#�5���V���y��4���㖼Dk�������!��s놼q�s�  Z���C�(2��E&����F�o��x� �0d$�;Q)��5/�6�>��H�� U��_f��~|���������謁�ӹ�P�ż��̼��ͼ�_ȼ̗����������I�����PV��4���0S���﮼�����)ɼ��ϼ��ϼ��ɼ�'��}=���7��Kԓ��V����z�'|l���b�J�\�֌Y���W�ϢW��X�t�Z�^���c�ySl�Y�x�鄼�:�����{��<��m˼�ּ sۼ�ڼ��Ӽ�Ǽ����(��;������ o���'��g���_�żD$Լ��޼�t�4��G�ڼ��μ���3ﱼzZ������p<��) ���7�������ւ��v��������� !���`���������������  �  �<Ӭ�<��m<#W<��@<�-<[%!<�<�b"<��0<ՕE<��\<�q<__~<���<5�y<h<~=P<?�6<r� <��<�N<�7<�9<m�-<(B<�V<e(i<�y<o߂<�Ӈ<���<rn�<H_�<S�<��<���<<�<�ى<��<�9�<�&s<��b<v|O<��9<�f#<�w<���;֞�;,��;d'�;�<�[%<��<<e�O<�Z<��Z<�OP<j�<<w�$<\�<���;���;��;<o�;�<�t<��(<vN<<�9M<ҽZ<��d<��k<��o<�{q<��p<��m<%6h<��_<�@U<1�H<��:<PW*<)}<�<+'�;�[�;kjW;I�:.�F:*9mJ�8��:�X�:q.;.Wu;s/�;��;��;߬=;�/�:��,���?h��׌�����cv����S����� ��zb��apL:��:���:��;�l;g�;��;pm�:Rr�:<Aq:S��9���s'�������g��U��Ūϻ�8����N8/�>��oE�� C���7���&���;3�3���)�������H:��W�r�"m����.ֆ��z��ؔv�,�e��hT�<E��9��T0��*�:x'��T&���&�)�K&.���4��=�xG�%�R���_�I�n�Q^��}������4��bɫ�9!��߸�����R���p���~���i���䄼.����������j���>���I@���ຼ�����������h��Q-�����cw��%�v��vm��Of��a�̒]��@\�P^]���`��kf���m�?w�)R��܅��pJ��ₛ���������	��aü�	Ǽ��ż����h���쪼��ݗ��x�����cޝ�|�������Px��LIʼֹμ
XμЙɼ����oҷ���V����Ĕ��s��f���_��3>����������#��gm�������Ϗ�S���0U���  �  ��<�'{<&1n<�Ba<�8U<�qK<n�E<9E<SK<��V<��f<��x<��<��<%�<���<�
�<�fm<FtY<�G<�:<4<Ye3<�7<R@<J<�T<�^_<��i<�s<s}<�p�<,��<� �<�	�<��<F��<�7�<�M�<F�y<n<�>b<7:V<��I<DX=<B1<� &<�<"j<$�<6%<�Q3<��D<B�V<X�e<��m<�n<[�e<8�V<��C<;�0<�:!<��<�<2O<|x<Xs#<͢-<��7<��A<�sJ<w�R<F Z<��`<ցe<r�g<�&f<�4`<GV<ݤH<?9<��(<$�<"<w7�;�F�;���;dv�;f;��<;"';�5);�C;
p;n�;7�;���;jf�;��;�֋;��?;]ѽ:cR8�����"���������� -źEH����
��_��ْ�9�C:	~�:��:-��:}��:6;�:�Jw:��9�"���Ǻ��"�m�a�����O��4�λ'��I�J��������>�?���P��?�r�ػ�Uͻ�һO��DZ�n���5�X�K��\\��f���j���i���d���]�jmV��HO�\�H�4�B��=�8��4���1�Vb2���6�|�>���I���V���d��or�������s��n��Vp��������Fܥ�'���UH��e���)�����/�m�v�pv���~�_Ɇ��"�� ���`Q��1q��0t��턧��E��~�����������	��C���K����:� �u��cm��Fg���d���e�sk��ws��}������m���j������@✼3H��2j��w���#B���Y��Uf���^��-ؤ��	��2���~���|���Ό�Y����F��^=������A���{���ѻ�y^���۶�R!���䬼=���;z��с��������������������>��є������f����@���$��*0���  �  >]o<��h<0d<V�a<�n`<&�`<��b<@g<��n<K�x<�y�<ˈ<t=�<��<�H�<�ҏ<���<��<;mx<>j<`R^<AU<� O<QK<?�H<`H<��H<z:K<�XP<h]X<bc<y�o<�[|<]w�<���<>ʆ<��<M}<M+o<f`<��R<f�G<ff?<��9< �6<�5<��4<�(6<O�9<�?<�H<T<<Pa<bPn<�x<y�~<}�~<�fx<�gm<��_<QUQ<�sD<~:<}2<~-<x*<��(<�K(<$)<?�+<�i0<��7<�@<�K<-T<��Y<&Z<z�S<.�G<1x6<5�"<$R<�&�;yv�;/�;Y��;�˧;�N�;6;���;«�;��;Ŏ�;�Y�;e��;���;Z��;��;��;�f�;Ҁ�;��S;Q�;�z�:��9Ï˹'	_�H��M����ͺ�YԺ�ɺ-��*�l��T͹�k9��:�EP:D{,:oa9��:�r캌C�Sf������i��� Ի�E�<��+��K���S������L��߻��λ�{��/���Q��-��mŻd������2��)��I9���E��O�(�V�j,\��,`���b���c��Ob��G^�'�W���O�HyG��nA�ܡ?�/pC��
M��h[��l�L~�U���6o��[E������ă��2���치�����V���=��Ƨ��a�������v��l��f���e�^�k�J�v��?��X�������┼	��������Y���񜼐᜼%
��)%���ꖼ/B��k]��rЅ��$�ƚu��q�Εr�8z�����M������&���C������q���䤼	���٥��ݤ���������J���������{ˈ�����;䂼�P��&���������ݝ��C��0M���欼�A��쩰�Z���Z���{���r��� ���$���/���י�?-��Y���?��x:�����+����G��݉��b����  �  Q�M<,�K<]zO<H�V<��`<�3k<z�u<��<K�<׻�<�f�<Გ<�.�<oE�<�z�<��<�<��<���<ڣ�<�:y<��l<MR`<nnS<�F<&
;<�1<u-<�-<��4<U�A<̀R<B;d<�Bs<�F|<�9}<"�u<�g<d;T<o�@<p�/<xM$<��<E�<�#%<?.<ݥ8<��C<��N<zqY<��c<n<J�w<�_�<Eσ<���<r��<t�<=i<��u<�
k<��_<DST<�zH<�3<<��/<5#<<;�<$�<O�<��<3!<t0<'><��G<�J<��C<��4<~_<�<���;�<�;?��;!@�;��;$�;�$�;�֦;3��;�r�;���;�Y�;ֿ�;��;_2�;Ȱ�;~��;���;�5�;��;Sv�;��q;v~2;B*�:\S:*q#�����t�|F6���Z��
k��c�f�D���d��q�4��A���P���m�� �0Z��p����ɻ���#��Y���� ��������ӻ�aĻ*ζ�AT���!��I��د��*S�������n��.<»1�޻�������v���.�^�>�N�N���^��pm���y����������wy�!m���_��pU���P��T���_�W�q�݃�����|��F6��V���z͢��X�����PᖼR�� ŋ��V�����ܐw�,|m��`d�gF]�WY�=bY��u]���d�8an��y����ʇ�8���l���'ݙ�m؟�f��wʨ�B$��R���)ˣ��o��i���'Ԋ����ƿ����������َ����
��uǩ������g��BG��	����J��������Ah���W���i��~���D��N>��g+{�[y��{�p����f��ϊ�
���\���پ������v����J��@0��|���+��Rü��S��L������k����#��Gb���㙼�G��n\��"c�������ü�  �  �^%<��'<^2<.C<SW<jlk<T~<�D�<�Ѝ<��<�Ɩ<���<J��<���<R��<�8�<>ɘ<�j�<�'�<�ۋ<�I�<0sz<�>g<�Q<'�:<��$<�<��<bA<�q<�L<�1<)+I<��\<�h<�Yj<E�`<tMN<�'6<�O<�<���;_b�;���;��
<��<`2<�G<�Y<�qi<w"v<�<��<ц<�ڈ<��<��<�`�<���<ڱ�<��|<�=r<F�d<�-T<x�@<v�*<y�<1$�;�C�;���;��;�
�;�3�;�<3 %<k3<��7<��0<�N<�V<:��;�z�;8K;��;���:0;��<;��|;f�; ��;��;Et�;��<t�<X�<�	</C<�&<�;)K�;���;��;��;��y;�C/;�@�:�P��k�ֺ~/O��ȓ�������Ż��û���������P��3�/�ĺ��4
��{\�w��s]�����)��t*���"�Xe�!��<����O��G��a����c{��t��)v�����㉻󩘻2ë�#[»�#ܻ[�����'!��8���P���j�eၼ�{���ߓ�v���dc��̖�������M{�;l���d�eJg���t��c��q���ɠ��K���ĳ�M��yﳼ���k����������Z��H�|���o�ؗe���]�|�W��6S�W�P��Q�ӤS�	OX���^��/g���q�)3��ه������q�����Ӱ���x��툽�����9���^g���袼��������;���E��ꡑ�k������\���;罼�üUü�'��݆��ح����ٟ��I󐼕ω�U1������Hy�ѝt�r�q�*,q���r��w�=}�$�����������0���Q��Tר��4��Gs���Fɼ�=м\Ӽ91Ѽ��ʼ\����,��Ó��4:��2Ơ�Oף����|��/=ļٸϼ^�׼�  �  �%�;�-<��<�&*<D�F<ed<ؤ~<�I�<���<�C�<zܛ<��<Z�<z+�<�Ҟ<Mٝ<�>�<�ߙ<�\�<�*�<���<i<�f<�WH<ţ(<�%
<���;���;H��;c��;�g�;��<xY.<v�F<�9U<FCW<	L<��5<)o<J��;�w�;ۣ;���;��;n�;�u<WF%<�gB<N#\<7�p<C!�<
f�<W��<���<�ϋ<3>�<�<�?�<�ʉ<�w�<0҃<?�|<P�l<�bW<A�<<��<��;�q�;9�;\t;Vn;�>�;��;�c�;�F<�+<��$<��</�	<r��;�N�;�;F�,:�]���U���S8U��:�U1;gs�;cѾ;r��;
�<�<�-<<�I<��<R�<Ge<���;��;E��;�<�;� �;��H;�|�:�y ��;(��ܗ��Ի�n ��������)�һȇ����j��'3�͕+�$�Y�N`��
�ܻ�C���0���G�`�R�b�P��$C��5-�������`���4К����v[`��R�,S�l�\�o�l�}3��ћ���p�����q�ǻ��9'�'��>�9��`Z��,}��e��ʷ������<֫�ʩ��B��B&��.1��`���xx���z�����Vؑ������a��Y���ȼZ�ʼ�nƼü����!���z��'��Yu���e��Z��S�/�O�*SM�TAL��sL���M��P�YLU���\�܉g��Yw�pI���x��f�����~q��ך˼	�ѼӺѼ>|˼�,��2������@��jғ�����朜�O9��R����ƼNҼ��׼�5׼��мreż�c��H���#�����P�����}�m@u�)p��zm��gl��l�(n�!�p�'�t�{��!��fĈ�A쑼�ʝ�o
��O����s˼Fټ�:�Ĭ�/���ݼW�Ѽ7rüDm���`��GF��$ݭ������wż��Լؾ��k��  �  ���;X��;���;H�<�5<~�Y<�Pz<��<XT�<�Ú<`i�<0�<*��<]�<��<��<��<�%�<��<��<�?�<��~<�j`<a<<��<[��;���;5�u;D�^;��;w�;��;Q<Jc3<�ZD<��F<�:<E� <wC�;���;$<~;m>8;��,;\�];�`�;���;�<<�:<��Y<��r<<�<F��<�3�<c��<E�<�[�<R'�<��<���<�<�m�<��<"�n<nU<�W5<�f<���;:�;l�';#�:�B�:�8;�q;HC�;��;�B<{�<o<Ux�;��;Nq6;7��9�̼��$�-��V��nѹ�	�:��h;���;+�;�<VO<rx<��<��<�Z<��	<ٰ<���;[�;���;�)�;-Z�;��K;/ӛ:��k��ǻ��uz"��0�9�.�I���A�+һ�ԝ�-�x�9�l�s%��P�û���[u-�hBQ��k�Ϸv���r��3a�\E�OD$�����xɻrי�$�q��ZL���>���A�G�O���c�p�z������ݗ��g������[�ۻ�Z��z�xP?�J�f�&#���P��'o���2��g���T���2��ꤼ÷��~���ń�������v��d���5_����мߏڼ�ܼx׼'�ʼ����h7��D���u����s�s�a���U�bO��K��mJ�J�$GJ��K�e�L�TxP�6XW��'c�EPu�xK��F�����.���xNμ7�ۼ��ӷ�1~ܼ�Tϼ����`ٮ��Y�����&[������j��ѻż�ּ�]㼕�鼒�輢�༒�ҼP@�����ŝ�?���)��:+y��p�f�k�
�i�|�i��|j�E�k���m���p��v��1�r߆�<|������谼5ļ7׼-�F6������B����c�P�'�ϼ��������u��z���y���_Ѽ�㼘����  �  �d};)K�;5J�;zN <CK(<|�P<Xtu<䫉<B��<㓛<Z`�< �<^)�<-ؠ<`O�<z��<1��<�
�<��<L�<�K�<��|<z�Z<E�2<`u<E��;�An;ф;l��:kS%;�@�;zE�;�<G{&<�8<k�;<;.<-a<�2�;庐;m)#;$��:#��:�K;�-p;���;u{
<��2<��U<B�q<ϸ�<��<�&�<ހ�<�ڍ<,ύ<��<n:�<B�<?׊<�\�<��<:n<["R<Ud.<�1<nz�;��I;ݾ�:w�8M��V:��;�ґ;v��;3( <5�	<P</y�;���;���:�L^���;�E���ꆻ3�S���ʺ��!:�?;N��;f�;��<U�<�o<��<k<�l<&�
<*�<�L�;���;%��;ak�;a��;r�E;s(o:aiҺ�!���v黊���:��H�U�F���5�����C��rΓ��f���K���s޻���v@��!g�z��b����E��gav���V�Iu1����Y!ӻ�'����o���E�m�6��:;�] K�u`��mw�Q��rQ������f���ٻrc���cE�4fp�M��ۙ���p��Gż:Yʼ�3Ǽ
�!.���x�����������B��h�������J���y˼d[ܼ���@��
��ռ��¼)������R��J�t�-�`�e�S��-M�j6J�	EI�'I��fI�m J��[K�h�N��U��b�#�u�"���vŚ�vC����ļ.ؼ�`缢�＀��)���ټ~�Ǽ����}����������[������μ	
Ἑ��$�����e�뼈ܼa�ȼ����Ԡ�d���79���w��(n�;�i��ph���h��i�e�j�>tl��o�2%t��}�����-��j⡼����lʼ��߼u��|������"�����C��:�׼�^Ǽ����L���4L���*ȼ`cټ��X �����  �  ��������"�]�� ������V���Z;pH�;�B<i�9<��M<]fY<X_<�a<��`<"E^<,FY<tP<"�@<�1(<di<��;�V�:�{K��^����H�p���������������:Mu���8����5a����!�ۺaGL��Qƻ�("��c��B���坼f^���'����v���3���һ����K;���;$d�;�@<�+<%�5<{;<��<<"�<<�y:<575<� +<��<a��;�b�;h\;=���ϻ[(4���y�*ܗ� Ŧ��V��̙��7��1�E�c�ξ���ړ�q���Y�񻈟4��{��A��Q[���ʼ<�ɼ<]���-��=����7�����g�LP��4�:&?;�3=;�MH;��@;��-;�/;~�:�n:�l;�A��b���e��,-�fNu�^���ȼ��Y���6����G*��C�߼���9]��蓼�������خ���μ[F�1	�c��=>��e�ķ�������ؼ\���,��~.r�#�I���.���(z��r�'k���m&�x0��>�D�R��No�`���N���RdƼ�켢�	�����,�K7���:�)
7�v-�X%��n��������N����4���!�(2��c@��!I�2�J���D��8���'�W,�m��I����ɼ՞��;���񨞼Ll��t���k���i�������-U���_��U��-����4ȼɏ�ɖ����'��i8�ĶE���L���L���E���8���(�9Z��1������v����I.�X�=��J��/P���N�f�F���8�o '��p�?������μ�#���x��Pf����������줼���z����~�����!����̼��⼖���17��C$�%7���G��.S��1X��U��L���>�`�.�%��������	^����͍.�+?�P7N��X��  �  iB����x�\�P��M�.Ȟ�r���$�f;�[�;�<p�8<�UL<��W<�]<j�_<�_<�]<��W<��N<�?<0&'<#N<�ȩ;���:�23����}�=�٨w��G���,��#ʉ�Hh�~�-�G�޻��j��Ѻ!3��6V.�Ľ����XUW�mX��j���w혼%��7sj�2�)�1Ļ.�ٺX�;N��;;��;v�<>C*<�r4<��9<��;<��;<,19<q�3<ϑ)<�y<v�;>
�;J�;��ͺ&»O�*���m�m�]_����;֒��v��P;��'�����D���8��U⻸`+��p�Pߙ� F��I�¼��¼ߞ���l���v�\�1�Il�3@a�M<P�#9�:�Z;��6;��B;�;;6&);��;���:��V:�獹m�}J����޻�\*�2p�����ü�c�x ��;y�����e���ټ���9$���F��M,���q��F���w�ɼjs켣�����������^}	�-�����ԼS9�������'q�!J���/��, �|��5��q�����l�'�K�1���?�T��Lp�g������ļ����R1���)�K�3��7�q3���)�bO�
����S�����;��oR��r��	/���<��mE��F�DA��l5��Z%��Z�)��fp�g�ɼK����L���n��`*���b���;���<��X_��Y��]&����������S	ȼ���$� �PT���$�"g5�>?B�o7I��'I�m%B�c�5��A&���'K��=��?��%��Y��;+���:���F�	uL��NK��IC��5�;�$�D��d�����s�μ�����1���,���]�����W|���V���g��(A���Ѳ��@����̼�T��P�����zL"���4��`D��O�9uT�%R�a6I���;�H ,����$��^������B,��><��J��U��  �  �r\��[P��,�~�ﻧ�e����9=ρ;�^�;Ou<�%4<��F<u�R<DY<��[<�[<��X<1 S<�$I<J�9<��"<��<z�;av;-�B���N����R�j�s��C|��k��_C��|�(樻����
Ĺ�G��P���xۂ����Y�4���e��������C0s�ȁH����\k��R|w�D�#;S��;*E�;#�<��$<3J/<c=5<D�7<�7<��4<�.<�$<I<���;��;�M&;��l��A���h�J�L�RX{�*���w���G~���R�:.�,�ѻ����>?�Lb�絻�'��JQ�PƇ�5>��紭�J��Iޡ������^��� �S�ͻf�T���f���Q:v�:�� ;R�.;ڿ*;��;�*�:�2�:�2:N��U�	�"�����ܻ]�#���b��n���4����Ҽ��7����9���ȼgF�� (���������D������|�����ۼ����<�������ȉ ����
�ɼ�"�� �� �o�ՊL��d4���%�J�zp�����#���+���6�;DE��GY��qt��O������5��H�����h�B9 �_)�ҁ,�GD)��� ��B��?������<�켕�����}��&M&�3���:��{<�Zy7���,�r��U��EE��D��ɼ�����Ҫ�7.������-���]1��:.������󛜼h桼M���ɶ�0Eȼ#J߼Y���T����]-�D�8�{�>�Ұ>�}B8���,�������L��eY �tJ����2��b]#�z�1��s<�*�A��A�V�9�N�-����X��C���X��Fϼի��cܴ��筼 ֩��ק�"i��#X��h����䮼8���@����"μ������,��]��Z-�`�;�v�E���I���G�$�?��3���$���2���9�0v�ڭ�	%���3��hA���J��  �  ����f��&�����lG�:};�;���;�m<�!)<�;<!�G<ÏO<ƠS<$�S<)pP<-.I<��=<��-<FG<g+�;`��;�9(;/���X~������AL8��>�/�͆��|��I�0���L@�:���:_:0�����a� ���+���E�p(K��:������ӻc$W�03��P0;���;X��;�^<�#<��$<�<,<m�/<�/<��+<�K$<<��<WV�;n��;Sq.;P�:�/�\�o�ٻ�F	D���X���X���C�cz�	��۲����5n���2ں�+h��)Իn�"�9�Y�u�������UO������j�?=��'�亻�bT�B���*9qі:�B�:N\;�];� �::[lD: f �⪫��5��\��Mc���A�R�̏��_��V����%˼-ӼT}м��ü>ʯ���G���m�:f��"v�o����%��ePü��ܼ3��_���z�����e|Ӽ�b��C���`��2r�o�T�	i?�X1��,)� �%�k�&��V+��3��$@�A;P���d�r�~�r����գ��⻼V׼���z�����g~�O�9�F���B�[>����%ݼ�QݼW��.b�����KK���$�Y�+��9-��c)��� �2P�ZA�[����K߼ż˼�E������������������(����������ġ�S����������w�ʼ�<޼-���3���1��e!�L�*���/��L/���)���0_�)E�������>��/> ���
�̣�G$�k�-��2�2��m,�#�"��z�n	�����19��~Ҽo�ļ��������Ԯ�Y��-O��Ye���_��8K��zl��CAż�aҼfa�ځ����-��v#��/��87�ě:�r�8��k1�i�&�+�:����������w��x����'�1[3�j�;��  �  S���V7���$�����	1���;B=�;fi�;��;!H<�w&<�5<��?<��E<��F<@B<,�8<L�*<�<��<�+�;�I�;((-;r��9�=������ƻ�r�:�\һ6$���z�_�Y94�;�l;?�y;R<;Ld|:��Ⱥ�'��M/ϻ̈�����w{��M!ʻ":����eY�9�';��;ٻ;��;><�<� <5u"<]s"<�<��<�<y�;c��;l^�;�4;�e$9�\�i����Kػݒ�����(���*����m��S�����9�s:
=�9�6����o�Ϋ׻��U3@��3W��+]�n�R��	<�J:���������w�Jh�%���0k�V�:���:�0�:���:�H:��P�7`��z0'�ޅ���$���/��G(!�T[H���q�I�]j��[ê�����g��i���%��_a�9A^�,�H���C�g+R�ӧq����{J����T̼�4Լ��Ӽ��˼pi���뭼hϜ��ό���}���f�{CT���E��;��5��D4��E8�i�A��SP��	c��Qy�yw��b��"���+ ���eϼZ伄9��tV�,�	��6���(��N+���C�etӼ3C˼w�˼j�ռ3:�GM����	����!��6��W����>��	��.�(�ἣ�Ҽ=�ż�������Ϊ�
���5ܢ��Ţ�_g��4v������(����}ż�^Ҽ?x� ����OG�I��-M��k�u����7)���M�����$��63�{��3g��n�	�d�C4�t� �!���M���j�/:�!���W�輱�ڼ_�μa5żlE���9���Q���籼;��o0���p��l�ż��ϼ֪ۼ���g���X����+K�x!�&'��	)���&�� ��������8��g��q���`���*��h6�����"���)��  �  �b��1�������S[(��p:g�	;�X;;V�;ٟ�;Oi�;=�<�4<�(<�51<Z3<*$-<1 <�
<I��;[�;���;>OT;	��:EJ:~�J����@:��(U��xG��@�p�,��I�:t�P;��;X��;�x�;i�;�Ls;V.�:�!�����\a��������
�`��a!�����^򑸁Ś:#�;s�s;��;S��;�q�;z�<�k<�<q�<���;`��;�ڢ;�Wn;�G;�:�����պs�<��[���h���ڣ��ȗ�<vm��a	�,�����:�*;�6H;{\*;���:AGK�MO����4�����������Ź��%���Z̻���}ш�GWN�~����4��G��O���)���Һi\?�2ב�[ ǻ�����N�n�1��J���b���y��3��~G��]���~ɉ�A���E�g�H�K�{�2��N#��� �p-��\G���j�����j֚����籼������}���ʥ��@��Ő��t򋼒f����u�!�e��bW�wM�[�H��K�ДV��rh��`�ϛ��B
��_\��a���*��-�ͼDڼp/����6�%n�^C��G�M5׼бɼj�����������P¼��м�T⼼���ea�<���
���/����� �����:�����jּ�˼�@������pذ��ܬ������m���f��!���X(˼Mּ��뼜���Z� �S��I
�u�������(L��l ���� "�nռ�ϼwDмu�ؼ�漋L������
��>����(����6������������߼�ռ�˼c�ü7���»�k����¼�˼Sռ}�)��s#��	'���F+�3B��g�x�����lD��������� �������7�^�"�󼱋�t*
��4��e��  �  0�;���:!��:#{:q�h:zԀ::#�:>��:Һ:;��;�˶;r�;Ra<�<��<��<s��;�]�;�}�;^xI;��:�y>:f@G8-"�����(�ы�Kz����:���:7-?;p��;i�;���;V <��<��;P��;ϕ�;UJ;>$�:l��9p�'��5���uϺ���7�ߺ~1ƺ���3���M:�;��s;ʏ�;�K�;��;;��;���;)P�;�v;��;�
7:�x��c��7���V�����r�#%�ٺ��v��%�8���:o0;
z;��;�i�;�M�;��b;&��:���'@�ϩx��"�� лJ�4\��������6	�ˉ��]��7�ǻVѠ�o�o��'�������x��Ee�n꨻��j���-� �C���S���^��Me�|i��Kj��'h�j�a���U��WE��E1����(v��Q�������� ��<���[�cz��q��:ᔼ1c��\���p���!��	}������w��1?������*z����|�B�l�6d��e�q~r��n��㒼���R���Ǥ��t�ȼX�ϼ��Լk�׼l�ټ�Uڼdټn{ռ�Nϼ��Ƽ輼qE��qͫ��A���ɩ�#����ʻ�D�ɼ��ؼ/<漬������<���#��������� ��������� i���⼯ ּ�ɼ�ٿ��G���
���2��O�ȼpռ�#��!�r���_������2��U3�r����e �6m�����y�6�׼q/̼<Kü�徼�뿼T=Ƽ��м��ݼ���T���x; �������5��n`��.��.�l��� �������m�߼)oԼ?[̼~�ȼf˼YUҼ<ݼ��a������N�	���&��S1�������,�	�k���� �A��;����޼��׼a9ռaFؼ�U༘�.m���M�&	��  �  v�;jjl;τ;bHr:�}��$㣺[:�7�ۺ�zn���9��;T�;���;f<�;(m�;��;�ٮ;
�^;<<�:B�D���z5�R;�=/�����i����Z:"�;tW;�E�;Fq�;��;��<�;<x�<qX<�b<;�<�X�;���;	�;R�L;��:�$�9ԙd��a��U��Ą�@��<�����A�ύ��$Q :�(;�W�;7�;��;( �;�C/;�.6:�߭�P8G��i��H�����O|��m:��ݺ���`X2:�M�:��C;_��;�-�;���;���;�h�;��;���;˂;:� ;�O:Kj���&�Vg��(@�����/�H�#� �1���6���0�� ��a�}�ػ ����肻�2s�����R㽻��\�'�kM��$k���~��w��	R��bxz��k��Z�O/I�P�7���&�I��S��Pe��ջ��ʻ[�ͻ���0 �\:�0��0K�ɯe���e��˘�	Ԥ��篼"޸��D��Rݾ�����Q��!+���1���l��{�������6��,��z_��ڽ���ϼ�ݼZ"強��8'�Rh߼\�׼4�ϼ�jǼ�D��I-��#��u��ՠ�1-���q���T�������)���*����μ4+ڼ���A�\���r���y<�F[�J�
�ʇ�5���Ar６:߼�Ҽ�ʼ6ʼ� Ѽ,�ݼ�����[�$���Kg��	��o��� ��������t��	ؼ�ͼs�ü�������������q�����"پ�Ʊȼ�Ӽ[�޼��.&��O �M����
� �����
2����� ����+�����,�ݼvټ��ۼ#6������:�
��H��Q�Փ��P��'����s	����<��j/��� �u�߼�ּ�μ�ɼ�	ȼeʼ?]м�ټG����aA���  �  o�;���;��;e��i(��@��鱶��"��'7��_pi�Ƨ����: _;JǞ;�5�;Eϑ;Z�.;�Ee9��ۚ���λ���/ֻ�v����]�����~�:�~L;F�;�i�;�. <��<� <d<*<�/<�0<��*<�� <��<� <i��;��;#�N;P��:�B����i��ͻ����h��u�B�뻒s���B8�1���{�:��<;��?;w0�:�'��/��J��r��p�������ӻ-L���[�#�+6�~ ;A�m;���;���;�;!��;O>�;^��;O�;���;��;֌;uK7;=8�:�_�Z!G�ꮲ��E���,�G�Q�l�l��nz��w��#e��SF��!��7���cϻ�����sֻ;5��&2�a�a��5���q�����C���K��3�����~�Cs\���;��%��3�e���ɻ#d�����頻RϦ�ͷ��ӻ�����g�)��$F��7f�#-��"���"���N}���CҼu�ݼ)y�G6ݼ]}Ѽ���~=���k��k┼K��s؜�-׭�5ļ��ۼ��� ��y�ӷ�������m޼��ͼ�����n������};������\��y��\���B��������Ȧ�#;���;����ʼ��ڼ�켠#���>	������Ϧ��V�i��������$�����iܼ��ۼ��h�� ���,�`��w��%��E���0����D~�������ӼibǼ���谴��$��ǰ������d���ʫ����U����¼vμ��ۼ�뼴����g���j��z ��#��!�p��[�"0	�������)���������B����#�z�"�g�&��p&��["�6_�'��Z�	��� �(����5ټh�ϼt>ȼ!�¼� ��*6���	��brļ�˼�Ӽ+޼�Y��  �  �w�;7�;�L�:���K֥�S���VE��I'��������<���4�麚�i:�-;��L;x\;QWg8|�=��sƻ~i��K.�E�7��/+�w���|����/���9?Z;M�;���;�-<�[&<_82<��9<Ze=<5N=<r9<0�1<�#&<�<�K�;��;po;�;a:���������z5�L�]�N�w";��x���ɻ9�M�l.�̪C:+�R:y)���?�`mû{��g�;��WR���S���?�q�LNֻ��\�{���L�;��;���;�;`�<��<�<u�<�<UN�;&��;9`�;��;�i;�K��h�5�û�T�.BS�V���8���6�����<��������U�tT+�7��w�}����0��b��-��Ӈ���]���bż�Sļ���i٥�"'��F�j��F<���2�뻏p��՟��g��@턻l愻.����K���J����ѻ����O���4��7[��ۄ��h��(����׼K��p���p��7 �L��ݼj�Ƽr�����q-��K��4ü�|ݼ����-	���l��@�����J�����fҼ����˪��1��I����Z��}ۉ����]!��q{��ߏ��qR��_���8���d����¼O\ּ���x��K{�<�c�'��-�&.��()�����s�������x��S�F�����O����U�(��s.���.���)�8� ��x�+T��-��̗޼��˼�o�������ͪ�����HS���	��`���j-��៨��9��Sq����ļCռ�h��� ���_��S{'��H0��~4�BS3���,��"�$-��p
��������T���d�H��:��Y+�OL4�
n8�7�+�0�ύ&���� �7� ���켬�ۼ��μ�cżƽ��k����t���o���k������?LɼުӼGn��  �  �C�;貇;���9�}o�y���f�2���W���d�X�9�3�����UR�������PQ:z�:�j�9���������I�ek���t��yd�e=��)��̍�QJ���G;|4�;�4<Et <�2<��<<W�B<;tE<IE<�B<�;<Å1<�M!<�M	<YO�;�Rl;38y9�m��|��8�:�Ƿk�RB��,)���rv�N<K�?u�����Z�/�����:��V#�����_��H�c�v�������Lw�J\I�,Q�7w��o脺�I;L��;��;}�<�<R�<cR<�G<�<H�<R�;���;�!�;ܺ5;�\[9^E�K3߻)4��y�pl�������۾��N��e~��Qj��{���EP�խ,�Փ���,��R��O��1��\ü]ټ�%�O��o+Ӽ���}����|}�`D����	ݻi����N���An��c��h���z�����o��O�����
���,��yY��N���I��j�ʼ9��6&�0������[������;iۼ$Jļ�ڵ�d��������Լ���d	��`�>� ��"$�Z� �����
�������ټ�⾼/���&���U֍��c��t^���΃����r������*�����ϧ��ݭ�[����ּ&��>L	����'H)�=}5�أ<�օ=���7�-�v��� 
�`���������)v�ٷ�;,��7���=�b�=���7��,��9�O�^����g߼3ɼ̃���Ƭ� ���f���𝼃��-������/W��Lh��5����L����Ҽ�3�H:����$�ۖ3��n>���C���B�{];��`/��)!�f���	��1�cP�'���q�E+��&9�ZVC���G��E�Y�=��81���!�D����=K켵:ؼ	�ɼ�����*�������峼������������6��klü�5μ��ݼ�  �  ���;�6q;�������=��.W��"��{}��{���xY�x� �(�Ļg-.�փ�d�19�s}���m�S��k�7��p��l��dk�����W`�0r"�$��w����B/;���;� 	<�U%<��7<u1B<?�G<�pI<��H<�ZF<�@<��6<ə&<7J<��;�<^;�м�瘻E1�J�Z�)Έ��꘼�*��TD���co�y�2��c�0 ���W�yH��nz���߻�.��Jl�@*��~����ڜ��Î��Tj�6(�����vںh3;�à;�N�;~�<fc<	�<u<,�<��<�"<� �;���;I��;K�A;��A9�u[�]���OH��]��棬��_Ƽ��ӼS3Ӽ
ż_����̏��	i���A�O	3��@��i��蒼P����ռЫ�L%���"��L���jʼ1���u���ML�!��:&ٻ2%����z�o�X���O��$X���k�y�����������׻���*��Y[� ��S���E�ռ�����6�	��b�\�����q:�|J���ϼ�����:���ȼ��༩� ������ �R$+�o�.��*�X� ���T��B����tC��5���S��Ꮔ�5���!o���䂼`o��t爼
����E��M��Ы�y��zXؼǐ�����g �;N1���>�-�F�^H�w�A�c6�M�&�!K�`�
�D�!��Y�	�����^%�}�4��nA��UH�6?H�h*A��M4�s�#����\ �yzἣ�ȼȣ��+���P��Q����Û��+��I����c��7���ܦ��6;������ӼA��E��p�s�+�)<�-CH��8N��M��E��8�M�(�:�����
��V�IV�AB#�Z3�`pB�+�M��_R�0P�(G���8��'�t�����Pv��F׼ZǼ�μ��v���#���ұ��Ա�=鲼D������ӱ���˼�gܼ�  �  �q�;r�d;��]����� %��:d��^���������f��H,���ػ7O��f��b��X��n���ݜ�8�C���}��Ñ��▼w8����l���,�ӄƻG$̺j�$;�;�;��	<3�&<9<M�C< �H<��J<�J<S�G<OPB<9�8<p(<�7<�T�;�?W;w��糧~c�5�f�;���EI������Z���#|���=�����1����!0���*�ʌ��U�f�8�t�x��0���m��!D��R���VGv�T�1���λ����S�:'�;~��;�@
<��<v�<+�<:�<k�<�^	<3��;n��;�?�;�8D;�9t`e�ս �ƌO�Wk��ݲ��rͼ�Vۼ'�ڼ�˼޲�(����q�EI���9�`�G�9�q�볗�U���=ܼ����YM ��g��b"�r�ϼX|��j��S�O��K�P�ػ[���w�t���R�|JJ��ZS��Bg����Tl�������%Ի+��y*�ك\�A���rz����ټ�( ��z���p  �=������/Լ�üƝ��}̼_7弤&�=���V$��.��J2�|V.�C�#�6�����6�⼍2ü;���ꖼ�����ă��ြ���nH��:؄��@���ی�)y���5��vU������3ټ~����1�a"��74�#YB�}�J���K���E��N9�C�)�ޙ�σ�e �t���z�J%�t(��8�F�D��L���K���D��H7��&��E�.!�.v���ȼ8��x��͉��4%��!��
������p�������᥼�����]��cӼ�#�zv�cK�#O.�PB?�$�K�o�Q���P��H�D;�b!+�E �������n��Z�F�%�36�J�E��Q��V���S�cJ���;��)��6����} 0׼��ƼN��\���Jp���7��dE��xP��q���5ĸ���Y˼�@ܼ�  �  ���;�6q;�������=��.W��"��{}��{���xY�x� �(�Ļg-.�փ�d�19�s}���m�S��k�7��p��l��dk�����W`�0r"�$��w����B/;���;� 	<�U%<��7<u1B<?�G<�pI<��H<�ZF<�@<��6<ə&<7J<��;�<^;�м�瘻E1�J�Z�)Έ��꘼�*��TD���co�y�2��c�0 ���W�zH��nz���߻�.��Jl�@*��~����ڜ��Î��Tj�6(�����vںi3;�à;�N�;��<kc<�<
u<7�<��<�"<� �;��;~��;��A;��A9:u[����*H�u]��ԣ���_Ƽ��ӼD3Ӽ
żT����̏��	i���A�M	3��@��i��蒼%P����ռޫ�\%���"��^���jʼ.1���u��NL�A��u&ٻd%��P�z���X���O��$X�ƨk�q�����������׻���*�uY[����A���3�ռ�����6� �xb�T�����k:�tJ���ϼ�����:���ȼ��༬� ������ �Y$+�w�.��*�a� ���^�C�,����C��5���S��폄�?���*o���䂼eo��y爼����E��O��Ы�y��zXؼƐ�����g �;N1���>�-�F�^H�w�A�c6�M�&�!K�`�
�D�!��Y�	�����^%�}�4��nA��UH�6?H�h*A��M4�s�#����\ �yzἣ�ȼȣ��+���P��Q����Û��+��I����c��7���ܦ��6;������ӼA��E��p�s�+�)<�-CH��8N��M��E��8�M�(�:�����
��V�IV�AB#�Z3�`pB�+�M��_R�0P�(G���8��'�t�����Pv��F׼ZǼ�μ��v���#���ұ��Ա�=鲼D������ӱ���˼�gܼ�  �  �C�;貇;���9�}o�y���f�2���W���d�X�9�3�����UR�������PQ:z�:�j�9���������I�ek���t��yd�e=��)��̍�QJ���G;|4�;�4<Et <�2<��<<W�B<;tE<IE<�B<�;<Å1<�M!<�M	<YO�;�Rl;38y9�m��|��8�:�Ƿk�RB��,)���rv�N<K�?u�����[�/�����;��V#�����_��H�d�v�������Lw�J\I�,Q�8w��q脺�I;P��;��;��<�<^�<sR<�G<�<h�<��;��;7"�;��5;Ll[9SE��2߻�(4��y�Ml��c����۾�dN��L~��<j��j��yEP�ǭ,�ғ���,���R��O��1��sü7]ټ�%�p�ἒ+Ӽ �������|}��D�ϯ�zݻ����PO�� Bn��c��h���z�����o������ỵ�
�V�,�yyY��N���I��F�ʼ��%&������r[������,iۼJļ�ڵ�c��������Լ���d	��`�L� ��"$�k� ����!�
�#�����ټ�⾼P���D���p֍��c���^���΃�"���%r�����+�����ҧ��ݭ�\����ּ&��>L	����'H)�=}5�ף<�օ=���7�-�v��� 
�`���������)v�ٷ�;,��7���=�b�=���7��,��9�O�^����g߼3ɼ̃���Ƭ� ���f���𝼃��-������/W��Lh��5����L����Ҽ�3�H:����$�ۖ3��n>���C���B�{];��`/��)!�f���	��1�cP�'���q�E+��&9�ZVC���G��E�Y�=��81���!�D����=K켵:ؼ	�ɼ�����*�������峼������������6��klü�5μ��ݼ�  �  �w�;7�;�L�:���K֥�S���VE��I'��������<���4�麚�i:�-;��L;x\;QWg8|�=��sƻ~i��K.�E�7��/+�w���|����/���9?Z;M�;���;�-<�[&<_82<��9<Ze=<5N=<r9<0�1<�#&<�<�K�;��;po;�;a:���������z5�L�]�N�w";��x���ɻ9�M�l.�˪C:)�R:{)���?�`mû|��g�;��WR���S���?�q�MNֻ��\�����O�;��;���;)�;l�<��<�<��<�<�N�;���;�`�;$�;�j;P����5�KûWT��AS�%���8���6��އ���������k�U�ST+�$��w����ԍ0�b��-��􇧼�]���bż�Sļ����٥�U'����j��F<�r��Ү�q���՟�Oh��~턻�愻4����K���J����ѻ$����N�@�4�T7[��ۄ��h�������׼��A����o��7 ��K���ݼT�Ƽc�����q-��R��Cü}ݼ���.-	�������X��7��K���	gҼ˭��/˪��1��n��� [���ۉ����q!���{��돏�yR��e���<���f����¼O\ּ���w��K{�<�c�'��-�&.��()�����s�������x��S�F�����O����U�(��s.���.���)�8� ��x�+T��-��̗޼��˼�o�������ͪ�����HS���	��`���j-��៨��9��Sq����ļCռ�h��� ���_��S{'��H0��~4�BS3���,��"�$-��p
��������T���d�H��:��Y+�OL4�
n8�7�+�0�ύ&���� �7� ���켬�ۼ��μ�cżƽ��k����t���o���k������?LɼުӼGn��  �  o�;���;��;e��i(��@��鱶��"��'7��_pi�Ƨ����: _;JǞ;�5�;Eϑ;Z�.;�Ee9��ۚ���λ���/ֻ�v����]�����~�:�~L;F�;�i�;�. <��<� <d<*<�/<�0<��*<�� <��<� <i��;��;#�N;P��:�B����i��ͻ����h��u�B�뻒s���B8�3���{�:��<;��?;v0�:�'��/��J��s��q�������ӻ.L���[���+6�~ ;M�m;��;���;7�;L��;�>�;���;��;0��;+�;�֌;�L7;V;�:M�_��G�����E�Q�,�͛Q���l�Knz���w�,#e�RSF���!�B7���cϻ�����sֻY5�'2���a��5���q�����|���K��q���Y�~��s\�S�;�8&�a4���|�ɻ�d��Q���A頻YϦ��̷�\ӻ��������)�J$F�E7f��,������䢭�}���CҼ<�ݼ�x�6ݼ3}Ѽ���c=���k��b┼J��|؜�?׭�25ļ��ۼ�� �z���ǫ������m޼��ͼ4����n��Ѻ���;��۶��~��;y��t���B��������Ȧ�(;���;����ʼ��ڼ�켟#���>	������Ϧ��V�i��������$�����iܼ��ۼ��h�� ���,�`��w��%��E���0����D~�������ӼibǼ���谴��$��ǰ������d���ʫ����U����¼vμ��ۼ�뼴����g���j��z ��#��!�p��[�"0	�������)���������B����#�z�"�g�&��p&��["�6_�'��Z�	��� �(����5ټh�ϼt>ȼ!�¼� ��*6���	��brļ�˼�Ӽ+޼�Y��  �  v�;jjl;τ;bHr:�}��$㣺[:�7�ۺ�zn���9��;T�;���;f<�;(m�;��;�ٮ;
�^;<<�:B�D���z5�R;�=/�����i����Z:"�;tW;�E�;Fq�;��;��<�;<x�<qX<�b<;�<�X�;���;	�;R�L;��:�$�9ՙd��a��U��Ą�@��<�����A�Ѝ��#Q :�(;�W�;7�;��;( �;�C/;�.6:�߭�R8G��i��H�����R|��m:��ݺ���wX2:�M�:��C;v��;�-�;��;̇�;i�;���;=��;�˂;�� ;0�O:Dj���&�Sf��?������.��#�~�1��6���0��� ��a���ػ�����肻�2s������㽻����'��M�]%k��~�x��LR���xz���k���Z��/I���7��&��������e�m�ջ'�ʻd�ͻk�� �&:�y�0�>0K�a�e�����d���ʘ��Ӥ��篼�ݸ�|D��ݾ�J��vQ���*���1���l��q�������6��",���_��@ڽ��ϼݼ�"����|'弘h߼��׼y�ϼ
kǼ�D���-��I#���u��)ՠ�R-���q���T�������2���0����μ5+ڼ���A�\���r���x<�E[�J�
�ʇ�5���Ar５:߼�Ҽ�ʼ6ʼ� Ѽ,�ݼ�����[�$���Kg��	��o��� ��������t��	ؼ�ͼs�ü�������������q�����"پ�Ʊȼ�Ӽ[�޼��.&��O �M����
� �����
2����� ����+�����,�ݼvټ��ۼ#6������:�
��H��Q�Փ��P��'����s	����<��j/��� �u�߼�ּ�μ�ɼ�	ȼeʼ?]м�ټG����aA���  �  0�;���:!��:#{:q�h:zԀ::#�:>��:Һ:;��;�˶;r�;Ra<�<��<��<s��;�]�;�}�;^xI;��:�y>:f@G8-"�����(�ы�Kz����:���:7-?;p��;i�;���;V <��<��;P��;ϕ�;UJ;>$�:l��9q�'��5���uϺ���7�ߺ~1ƺ���3���M:�;��s;ʏ�;�K�;��;:��;���;(P�;�v;��;�
7:�x��h��=���Y�����r�"%�ٺ��v��)�8��:�0;mz;��;j�;N�;��b;���:�臸�>��x��!���л3�[�����/����Ј��z��p�ǻ�Р�j�o�]�'�A���u��Sx�)Fe��꨻F�zj�U�-���C�Q�S��^�INe�i�GLj�w(h��a�@�U�XE�@F1�յ�Vv��Q������b� ���<���[��bz��q�������b��:\���p���!���|��}���w���>��Ğ��z��m�|��l�!d��e��~r��n��$㒼F�������������ȼ��ϼ��Լ��׼��ټVڼ�ټ�{ռ'Oϼ��Ƽ@輼�E���ͫ�B���ɩ�4����ʻ�L�ɼ��ؼ2<漮������<���#��������� ��������� i���⼯ ּ�ɼ�ٿ��G���
���2��O�ȼpռ�#��!�r���_������2��U3�r����e �6m�����y�6�׼q/̼<Kü�徼�뿼T=Ƽ��м��ݼ���T���x; �������5��n`��.��.�l��� �������m�߼)oԼ?[̼~�ȼf˼YUҼ<ݼ��a������N�	���&��S1�������,�	�k���� �A��;����޼��׼a9ռaFؼ�U༘�.m���M�&	��  �  �b��1�������S[(��p:g�	;�X;;V�;ٟ�;Oi�;=�<�4<�(<�51<Z3<*$-<1 <�
<I��;[�;���;>OT;	��:EJ:~�J����@:��(U��xG��@�p�,��I�:t�P;��;X��;�x�;i�;�Ls;V.�:�!�����\a��������
�`��a!�����`򑸀Ś:#�;s�s;��;R��;�q�;z�<�k<�<p�<���;`��;�ڢ;�Wn;�G;�:ȑ���պu�<��[���h���ڣ��ȗ�vm��a	�	�����:*;n7H;M]*;���:{BK��KO�L���3��@������;��[%���Y̻'����Ј��UN��|����n���������)���Һ;]?��ב�
!ǻ���� O��1���J�e�b�?�y��3���G�������ɉ�q�����g���K���2��N#��� �p-��\G�\�j�f���=֚�����籼�������}��?ʥ�W@������9�\f����u�ԗe�hbW�OM�F�H��K��V��rh��`�����p
���\���a��+��p�ͼ�ڼ�/��7�dn�C�H�{5׼��ɼ������������P¼��мU�º��ga�=���
���/����� �����:�����jּ�˼�@������pذ��ܬ������m���f��!���X(˼Mּ��뼜���Z� �S��I
�u�������(L��l ���� "�nռ�ϼwDмu�ؼ�漋L������
��>����(����6������������߼�ռ�˼c�ü7���»�k����¼�˼Sռ}�)��s#��	'���F+�3B��g�x�����lD��������� �������7�^�"�󼱋�t*
��4��e��  �  S���V7���$�����	1���;B=�;fi�;��;!H<�w&<�5<��?<��E<��F<@B<,�8<L�*<�<��<�+�;�I�;((-;r��9�=������ƻ�r�:�\һ6$���z�_�Y94�;�l;?�y;R<;Ld|:��Ⱥ�'��M/ϻ̈�����w{��M!ʻ":����eY�9�';��;ٻ;��;><�<� <5u"<]s"<�<��<�<y�;b��;k^�;�4;�e$9�\�j����Kػݒ������������m�S��K��9M�s:�B�9�4��~�o�.�׻����2@�G3W�+]���R�p	<��9����� ��,�w��f�z���dY���:Ф�:L1�:���:�G:T�P��a��v1'�z����%���0���(!��[H���q��􌼚j���ê��������Fi���%���a�aA^�C�H���C�Y+R���q�쁎�ZJ��� ��%̼X4Լ��Ӽ��˼2i��r뭼+Ϝ�Rό�R�}���f�(CT�r�E�Ҭ;���5��D4��E8�y�A��SP�
c��Qy��w�����W���e ��fϼ]Z��9���V�J�	��6���?��w+���C⼃tӼKC˼��˼y�ռ?:�OM����	����"��7��W����=��	��.�'�ἣ�Ҽ<�ż�������Ϊ�
���5ܢ��Ţ�^g��4v������(����}ż�^Ҽ?x� ����OG�I��-M��k�u����7)���M�����$��63�{��3g��n�	�d�C4�t� �!���M���j�/:�!���W�輱�ڼ_�μa5żlE���9���Q���籼;��o0���p��l�ż��ϼ֪ۼ���g���X����+K�x!�&'��	)���&�� ��������8��g��q���`���*��h6�����"���)��  �  ����f��&�����lG�:};�;���;�m<�!)<�;<!�G<ÏO<ƠS<$�S<)pP<-.I<��=<��-<FG<g+�;`��;�9(;/���X~������AL8��>�/�͆��|��I�0���L@�:���:_:0�����a� ���+���E�p(K��:������ӻc$W�13��P0;���;X��;�^<�#<��$<�<,<m�/<�/<��+<�K$<<��<WV�;n��;Qq.;h�:�0�\�p�ٻ�E	D���X���X���C�Zz��໷������<m���1ں�*h�_)Ի,�"���Y�L�������%O��p����j�?=�2'�Q㺻�aT����*9?Ӗ:D�:�\;,^;� �:���:�jD:�o �y����5�%]���c�p����R�����M_������&˼�-Ӽ|}м��ü[ʯ���G���m�=f��"v�b���z%��JPü��ܼ�2��_��wz��̤�3|Ӽ�b�����1���r�!�T��h?��W1�f,)���%�\�&��V+�+�3��$@�j;P���d���~������գ��⻼�׼3�󼔌���~�f�%9�Y���B�x>�����3%ݼ�Qݼd��7b�����MK���$�Z�+��9-��c)��� �2P�ZA�[����K߼ż˼�E������������������(����������ġ�S����������w�ʼ�<޼-���3���1��e!�L�*���/��L/���)���0_�)E�������>��/> ���
�̣�G$�k�-��2�2��m,�#�"��z�n	�����19��~Ҽo�ļ��������Ԯ�Y��-O��Ye���_��8K��zl��CAż�aҼfa�ځ����-��v#��/��87�ě:�r�8��k1�i�&�+�:����������w��x����'�1[3�j�;��  �  �r\��[P��,�~�ﻧ�e����9=ρ;�^�;Ou<�%4<��F<u�R<DY<��[<�[<��X<1 S<�$I<J�9<��"<��<z�;av;-�B���N����R�j�s��C|��k��_C��|�(樻����
Ĺ�G��P���xۂ����Y�4���e��������C0s�ȁH����\k��R|w�D�#;S��;*E�;"�<��$<3J/<c=5<D�7<�7<��4<�.<�$<I<���;��;�M&;�l��A���h�J�L�QX{�)���v���G~���R�1.��ѻ����P>?��b��浻�'��JQ�6Ƈ�>��Ǵ��(��&ޡ�}����^�_� ���ͻm�T�v�f���Q:cw�:� ;��.;�*;��;�*�:S2�:81:����	�������ܻ��#�Ȝb��n���4��߸Ҽ��W���(9���ȼwF��,(����������D������m���q�ۼ����/��������� ������ɼ�"�����ío���L��d4�h�%��I�ep������#���+���6�XDE��GY��qt��O��-����5��k�����h�T9 �_)��,�VD)��� ��B��?������<�*켞��������'M&�3���:��{<�Zy7���,�r��U��EE��D��ɼ�����Ҫ�7.������-���]1��:.������󛜼h桼M���ɶ�0Eȼ#J߼Y���T����]-�D�8�{�>�Ұ>�}B8���,�������L��eY �tJ����2��b]#�z�1��s<�*�A��A�V�9�N�-����X��C���X��Fϼի��cܴ��筼 ֩��ק�"i��#X��h����䮼8���@����"μ������,��]��Z-�`�;�v�E���I���G�$�?��3���$���2���9�0v�ڭ�	%���3��hA���J��  �  iB����x�\�P��M�.Ȟ�r���$�f;�[�;�<p�8<�UL<��W<�]<j�_<�_<�]<��W<��N<�?<0&'<#N<�ȩ;���:�23����}�=�٨w��G���,��#ʉ�Hh�~�-�G�޻��j��Ѻ!3��6V.�Ľ����XUW�mX��j���w혼%��7sj�2�)�1Ļ.�ٺX�;N��;;��;v�<>C*<�r4<��9<��;<��;<,19<p�3<ϑ)<�y<v�;>
�;J�;��ͺ&»O�*���m�m�\_����:֒��v��P;��'����{D��{8��2⻣`+���p�Cߙ�F��9�¼��¼̞��}l��Z�v�8�1�l໲?a�}:P��9�:A[;��6;��B;.�;;<&);�;Q��:ԷV:ꍹ�m�J����޻�\*�Vp���
�ü�c伉 ��Cy�����e���ټ���?$���F��M,���q��A���o�ɼ`s켝�����������U}	������ԼA9�������'q�J���/��, �m��+��k�����q�'�U�1���?�*T��Lp�u������ļ��&��[1���)�T�3��7�q3��)�hO�
����S�����=��qR��r��	/���<��mE��F�DA��l5��Z%��Z�)��fp�g�ɼK����L���n��`*���b���;���<��X_��Y��]&����������S	ȼ���$� �PT���$�"g5�>?B�o7I��'I�m%B�c�5��A&���'K��=��?��%��Y��;+���:���F�	uL��NK��IC��5�;�$�D��d�����s�μ�����1���,���]�����W|���V���g��(A���Ѳ��@����̼�T��P�����zL"���4��`D��O�9uT�%R�a6I���;�H ,����$��^������B,��><��J��U��  �  �H��^B��0�5l�9Ｆ���?�i�����v]���9��&;�A�;��;�ٰ;;n�;^ש;i��;�];��:Ұ���[����*�h����ȼ�o�t8#��r<��]L�`P���G��4�$�����;�Ѽ�ݴ�򿯼�SüS���X���+���B��P�9�R���H��y3���T���꯼��n�:�8?��������`:�;�,D;�Z;�rZ;t�E;��;5K:�L��𛈻�u
��5f��ꪼ�����*2���H���T��T�s�H��3�YS��b��Yؼż��ʼ�������)�^F�]�[�1�g�Z�f�ݐY���B��%��l�.SѼ����[�h���+�K����һ�������1���Z�ƻ�6��Z���%��iR��������dw��11��vQ�?�m�[������"F���{w��Z`�F�
.���^$�/���1�!�K���h�7���YǊ�]��	���.���l�S$N��.��-�_���μ_���^��t�	���g��c����������h���f��b׼������}.�;�M���n��@���C�����,2������^���s��[s� S]��NP���N�+�Y�Wo��,���F�����E���m��*N�� ̗����cs�B�S�|7����<���� ��X（��)sݼٔڼvnڼ��ܼ��h�����E�����4�B�P��p����o���&᡽�䧽󼧽����������/�w��c�ZX���Y���g�oT~�v挽�8���z��s��������s������.���mNm���N�m24�϶�����I�2�����|��
�#�#��q�����*�<�-���F��Bd�N9������㟽`���z���V���x���0���
�����z�0Ji���b���h���y�R]���P��&𳬽�  �  �EB��O<��A+����R輰)���e����cab�mB��;�R~;�#�;�-�;��;��;�%�;=�N;�K�: 麺8ݫ�S�(�1凼�ü� �ׇ���6�n6F��J���A�wN/��N����`�ʼrܮ��䩼;����<���W�&�=���J��L�ЬB��[.��������3���dk���P����|º�':��;��7;p�N;O; �9;�	;#�E:�����-l
�_$c�Yr��h��l��)-���B��N���N���B�j>.���������Ѽ�<���żS�u��	(%�1�@���U��Ma�Y�`��S��=�3�!�����Rμwm��Ei�e+.����ڻ[w������$���m̻�����	��;)�
LU�&ψ����%h�[\���-��M��/h��o{���*����q��L[���A��*��z��;�!��.���G�_�c��b}�����5������^d��*h���J��,�!�[#��μK|��E������Y���XΒ����&���.��1v�����ܝؼ��������-��iK��ak�V焽)x���������}���ޏ����	o���Y��HM�QL�0�V��Gk���騐��!��6!���H��d\��u<������hp��R�ǜ6����k3�<d�B"���a�޼�ۼ=�ۼ�u޼i�伧��@5 �Љ������3���N��/m�=���/������ä�����0���s퓽Mچ��s�I�_�]iU��V�Z-d�az�ԋ���}��Pt��}r���s��"������8���F�j�tPM�2�3�����1�k ��v��kV𼣓�%$�q�|��������0h��w��|-�ߢE��)b���������;������!����k�����d��tՇ�Xw�}0f���_�@xe�-v�vD���Ԕ����ߜ���  �  ā0�l[+��6�$���ּ���/�Y�X��gx���%�'�:��P;lN�;�^�;2�;ِ;��q;� ;&U :!���<���b%�����@�����v���P'���4��B8�&�0���������fo�����6��	ժ�9ϼ����,���n,���8�;��>2��& �	����ؼޡ����c����g��k����ǒ�:��;�/*;2�*;�;ķ:��:8�8 �8��g�Y�\�M���]�Լo��F��2�2=�G�<��32��C�/���`⼋_�������7����ϼVw�����P,1��D�h�O�i5O��(D�q�0��������Ƽ7��3�l���6��?� V�k%ջsdʻ Iλ�߻H�������4��>_�nы��@���Jݼ���4%�_!A��dY�o�j��'r�r�n��qa���L��5�)R �������n�$�P�;���U�nWm�)~��W���"��R�q���[�ʴA�R�&��-�ta�+pѼ�Y��_ר�oe���ޘ��u��E��� ���=o��:#����żC
ݼ��������)��D�n�a��|�,���F�������ޏ�3���kz�ȅc��1P�ڬD�`�C�(�M��`�e4y�7=���͓�AI���u���"������恽�dh��6M�4�4�U � �������F;�o 伟�༒]�k��.꼣V�����x���'62�zrJ�.�e����^;���ۖ�����?����*��Bi��*i���#i���V�h	M��|N���Z�%o�A܃�&����꘽����Ɯ�����z���C�z�c���I�{{2����Y�����?�������l�t�����F����j����:���T-�0C���\��{x�����ؕ�84��9�������8���ꍽ����H&m��\]��wW��\�$+l�8N��ȍ�����栽�  �  9��u�������&ֽ�!c��D�O����=U������"�9�F�:�&B;��h;c<p;e�X;�b!;�U�:��C���P�$�λ�T'�%@t����nӼ����U
�,���:��B�Z���較���I}�����.-��%���U��g�ؼ��������Db!�v��`�pa�z�ü�����_�%���Cǻ��a�u{��(wb8�s�:	b�:�i�:��:��9�'��ǺW�΅���o�_�Y��Ŕ�	��R1��!U�o�#�{�"��z����K�鼘A¼n���Õ�����L���ڼ?�N�:�+��5��6��-�|���	�2����V���!�x�VJ�̍'����5���^M�1"��I�Q��+T*�~�J��t�屓�xH��,2ټ�O�����{0�bRD��TR��>X�U�UI���7�*o#����r��� �c���M�)���@�)�U��kd�<�j���g��W\��J���5�{��G������2�ؼW�ü������Ϟ���Z���������!T��뾼��м|��(.�u��&���<��2T���j��
}�Qp��S���(��ϩx�%f�ZIR�ܠA� �7�7���?�ƳP�V@f��d|��}��dL������/H��+
��'At�h�]��G���3��H"��X�l	�D�Я���{�{Y鼑 �(��4���9 �N\�^��� ���1�o�E���[��Ir�9e��p.���8������ŉ�i<��n�m���X���H�@w@���A��sL��T^��s�tD��S�����,-���f���!��kq��[�/�E���2���"�,�,s������������c�����k���f���z,�_����.�NA��+V���l�_���9S�������dȒ�����<���Sq�Z�]�rP���J���O��,]���p��F��2!�����  �  ސ�c�i޼2Tż���5|��}�R����/�ڻO��� ���P��N4�:�k�:��;!�:]�:Ӊ��.H�3���l���8���r�G�����[ؼ���b��~G ��|�ڼ٭��+�����o���J���D��q^�@����諼~�ϼ�=� � �g ��켒�м�����ۑ�V�h���3�>������q�"����Q��D6����@�����Vh�F÷��s�1�qe��A��&��[:м� �2`�Ĝ���<��O�ݼ&J��2���p���4p��z�ݰ���b��ټ����~�����]���� #
�ݵ��ےڼ+��6V��3��9�n��M���2��`������T��v0��L��p�����	���L����ۼ�������sJ��Y-�}7�}�:�M7��-�[��������\��^�5��N����
(��9���F��M�:L���D���8��>*�t�����1��P�pUּ3�Ƽt�����rg��[���7�������zмHK�A���Û�L���%��66��GG�TW�jd�|�l��n�׶h��8]�X�M�@�=�??0��R(�(�'��/�O�=��O�eXb�b.r�\�|�W��g|��Kr��zd���T���D���5���(����y��A:
��9��}��98�����p���#��DZ	�u�����;'��e4�A:C�]7S��Bc�֨q�,X|�R���3t�C�v��#h��V��E��Z8��x1�J�2�~z;�QJ�[ \�/�m��K{�ډ���⁽��}��hr�+�c�	T��D��p6���)��8�K��������̎���������V�����6(�r4��eB���Q� Ab�&r�"��Bp���ꅽ�׃���|�@m�g�[���K�#T@�� <��@��KK�[�8�m�nO~��/���  �  &_��s��Ah�������A��>���Km���I�k�$��+��񻲻U�Z�f_׺�&�����˻q�����a��\mֻIw��V;��b�^��媖�����}��5Cļ_ɼS�ż�a��݉���d��V0W��i(����p��A>���D��{�V���7V����ƼnϼT�μ��Ƽ���4���������Ze�֋?���d��#?����^�ߣ&�N$���W�#k���&໡%�oc=�/�c�㘄�P�������/����ȼܦҼ|>ռ�μ�0���0��l�����h��gC���2���;���]�-g��J騼�Gȼ߫��������g��,��?�ּ��Ƽ�O��4���H���b���7�g��M�P�=��S:��D��\�G8~��œ�������8oռ�꼈&�����������L�s���Q�������"Ｆؼ}�ȼ��ļdpͼλ�|����ڃ��)�{0��&2�R�/���*��e#��f�`)�k�
�p�k���⼎�ӼH/ȼ
¼У¼�	ʼ��׼�7�������
�j��d� �P�*�d�4���>�kQG���M�oQ�T�P��K�5^A�z5��(��9��T��^�����*��8� �G�(&U��^�nc��Wc�\L_���X�VFP��]G��6>���4�K+�aw!�����S�����M��YO��{�9��6b ��<*���3�xM=��F��O��/X��p_��8d�9Ie���a�bqY��SM��J?�9�1��N'�4�!���"�#�)��5�q�C�)R���]���e��ah�/�f��a�nZ�pR�JII��Y@��;7���-�hO$��@�����Q�S"�1^�����'�3D"�1=,��I6�f@�C�I��	S��0\���d�vZk�61o�C�n���i�_Y`��zS��vE��8���/���,�H�/�3�8�p�E��OT��b�f�l��  �  �ⅼ����8��X0��8����З�/����m���zv���P��!%����㨻�xr��}Y��6���Q��

�k�8���e���V-��՚��|��Ä��2���S&��,X���.��`����`�T�4�(T	���˻����l��n��p�����&�KU�P���Ź��"?m����� 쮼0a��W0���v���9��s���i���;�q���ݻ�����ƴ�X<ػ�;�o8���e�i�����7������W���D鱼�������9����m��M|��ѭo�&�E�>��{�����*��6�AG���y�� ������7����ϼ-ټС޼)fἕ��V%߼$�ؼ��ͼ<*������H疼�:���r�q9k��v��=��՟����yҼ��7��������N�	���
�׍
��� *�Q\�����:)ڼ�Ƽ���oL��+���v������.�ռ�S＞/��
��l�b@��� ���"���#�`;#��;!��7�g���J�{Y��������Qiۼ��ڼ��� +��p.���j���)�l�1�͊7�;���<���=��Y=�:T;��=7��0��7(�vo�����t��m	���	�o��%���E#�ɡ/�d1;���D�`�K�<P�d|R�hS�US��aQ���M��"H���?�̓5�&*�T3�2������m�����q�(��J4���>�tmG���M��RQ��SS���S�*}S�=�Q���M�{�G��w?�S5���)��U�Us��}��8�����"�E�-��C9�ǽC�iL�P�Q�$�U�XhW�hX�pW�nU��~Q��1K�uB���7��,�A�"�k{�[���� ���)���4���@�u�J�(�R�{?X���[��M]�U�]�S]�7�Z�e�V���O���F�� <�p�0�eS'�� ��f��� �ז'��1��#=���H�ЃR��  �  �(C��Ni�1o��6���
��C���`7��S1��`����������bTI������n߻Sg ��A'���\�͔��Z9��!�� �ļ�ż�񾼦V��~����E����-[���5�(���{Ի�i���7��2��ẩ����}�k���V��#�.��U�.|��ϐ�f.��妴���üdμ��Ѽ�[̼�2���奼����[}\�Ss/�����]�e,�^�W�t{��\أ�����̼ixӼ�>Ѽ_�Ǽዹ�m����������h���D� � �����i.Ż�x��ᒻah���eͻ�����0�A ^�=Յ��曼4����ż� ڼF�켁<��6�ym�� ���� �ڼc��nB���a���Y�����������ƼW�aL����zb�RE�ѳ�X��o�����AX��&�漕�ռ*�ļޜ������ѧ��3���:ӏ�\��7���?k��Cgɼd�߼�����Z����h���/#���+�B�2���6�J!6��	1���'��[�ps�6l�[6���T��>������c*���8��C�"J�b�K��H��MC��#<�R4�LV,��N$��&�5�����V��Њ��U}�������y��m����k���x&���0�~�:��/D��xM��8V�0�]��b���d���a�O�Y�|0N��@�%2���&�(E ������%���0�v�>���L���X�c)a���d���c�4�^�۽W��]O�/�F��x=�VG4���*��/!�r�����I
�t3�!��"�����M�l!%��$/��8�lrB���K��T���]���d�Y�h�Hmi��.e��C\��O�"�A�+�4��+�̸&���(�>�0��4=�O�K��Y���d���k��n���k�Rf��^��lV�}�M��D��;��52���(�����������5��	�j��� ��*��"4�b*>��  �  r	��P�r��j:��&�Ǽq��(��d�������\Ӽ`�������b�:�8�~X-�EB��Xs��L��=|����߼ɞ���E����������̼ͭ��?���`���+�����Lt���:K�����rg��:G�!:,u�8���j�-��ᙻ�軕�!���U�����짼9Mȼ���������������|ܼ���}9��0?u�yJT�9�R���p�o��RԶ�N�ټŕ����h��� �A����μ�t���Y����g���5�`K���λ͓�leO����<���,���r��n��E���/$��S�6ʃ��;��ģ��z��$�����?��!����a��������Tм�ι�^=��X߸���ϼ�i������,���3�b4���-��F"����ܥ����NrѼ�����M�����*��,	����x�*�y�k4���x��V��Q��jb¼�ڼ���hV	�X����*���:��)H�~�P��YS���N���C�Y�4�r$����ߟ�8�
�`w����v1��KD�aiU��~a�E�f���d���\��TP�4�A��2�ع$�hf�1��L��w��e�Z�輭��y���J���5�Z�}���#���0�2�?���O��_�U�n��*z�����B��Qw��wi��)X���F�=8���/�sz/���6���D�@0V��g��v��~�aJ���n{��p�Yfb���R���B�0N4�Gv'�P�`��`|
�7 ��2��'�������nM������ �;�,�gZ:���I���Y��i���w��a���xy��Ty�j�ĜX�
H�&�;�c)6���8�/�B��xR�>�d���u��F��ǟ���h��(逽��u���f�'5W���G�_":��.�Ɉ#����r��C�h�	�����
�"�������Jq%��\0��  �  H5�/N�R	��˾���뼒��0�����R/�|� P������s����v�&�h�k뀼 l��C�Ƽ-P���ĺ�����r�"
��5�Oe¼/����Z�������Ae>���Y�'Y7:u��:�-;�];x�:ԕ|:�,비)�����/�lG�������0�,����H=!���!��;�E	�~���߾�OM���g��"i��e���������o�X`�"���"�6V� �
�8o�ӿ��m���m[�`��b�лxɃ�O������0���
�.�|�0���%Z��Ŭ������X1�2�o��.��RYȼ�%��m��y�'��7���>���<�$�2�D�!�B�����ڼKϼ�׼�k�hB� $�D�9���I�l�Q��P�q�E�:5�Sa �s�
�y�HUȼ�F���ݔ��=���q��gb��P\��Z^�,h�M�y�޿�������ﯼ�lʼ���������W[6� �L���_�K�l��2q�F{l�ۙ_��3M�G9��g'�u�>���A!�Q>1�c�F�&�]��q�G�g������Ks�C
a���K�s�6��#�T���y����ԫ輲�޼cټ�f׼U�ټ�I߼��輤7��������j��5-��A��$W��m�Vw�������g�����5H��C'���o�|pZ��I��?��>�\�G�@DX�w7m�q�����hp��Ǝ�y��� Ă�#q��Z���D��*1� � �-u�1	��d������m��]�q0����5����Y�R��P�՟&�<8���L�Xac���y������H��F���
w���݊�rY�n���Z�6�K�)E�dH��?T�Jg���|�܉�����ܔ���y��b���\��}s��2]�(H�r�5��\&�'T�f��#
��T�������������G����d'��t(��  �  � ��{ Y�}���ݗؼ�]��2�r-�5�2���,��.�\���Lݼ�+��@����`������oA��B�뼒��tU$�f�2�ɉ6�0�/����Ns���ؼZ���Z�a�����f��+CӺ�:��;��=;':Z;�%\;��D;P�;MUk:Ŋ��iu����fG�i��%�ȼ{9 ���Q�.��:���;�T2����bD��-༪���(ơ�����%Z��\�ۼ<����ZJ1�*<��*<���1�����=Ӽ�᝼��]����wE��b+1�����7�B8��:��:�L�8*iF���D�|�ӻ1� ���g������Ӽ}Y���"�3<���N�8WX���V�I+K�L�7�l� ���
�c��4��W�����I�8�r�P�[ c�z~k���h���[���F��X-�mv��e��Ƽg��eԊ��(r�&A[���N��9J�xM��JV�JDf�o~�����v̥�^5ü��}���[&���B��Z^�-�u�ظ��{���Z	��gMw�=b��J��;6�y)�40&�7�.�c�@�3�X���r�߄�l}�������닽����Oq��W��<���$�"���U�*d켍Vݼa�ӼDϼIYμ�м��ռ{޼�뼈k��t�	��t��B-��+E�;`�t�{�슽!���
��P����Җ�1�������nk�B.W���K��K��pU��h�YQ���\��
��}q�����34��j{������<d�xI��1��\��9��o����9�3����\�va��4񼷉��_������$� �9���R��n��߄�s*��3��k����i������݌�^Ā��zj��JY��Q���T��b�%cx�z���(?��vʜ�����w랽���T���=��*e�wEK�(�4���"��Q��}�p��X ������������*�������Z	�2�$��  �  \���d���*뼉���_-�oy>�_D�E#>�!+-�������Ƽrަ�J����S��{�ѼW�w#�~�4�D�	@H�H@�l�-�>���86���Yk�/�|����ҁ�\��:e�/;��f;`;�>�;�k;�<;<_�:����S� ��ZtL�������ּR�
��'���>�}�K��M��UC�LH/�|��Mm��P_˼7���]l����Ǽ/�����-��(B�#�M�*�M�'�A���+�;��⼹�����c�Ј�3������u��k�7:���:��:�S%:Ic%��M��Q�T��1������)g��J����ݼ����G.���J��|_��j�Ηh���[��eF��-��������A�s��j*��FF��`��;t�r@}� z�a]k���S�4�6�������mȼ����5����f���O�Z�C�'�@��D��L�#�[���r�p艼��������m��c,�)L���j��m��5>��=~������4����p�V�� @���1��t.�U7���J�<+e���������;���ɗ�I>��O��w}���_��B�%%'����Pc��7��v׼Bμʼ �ɼ�˼��м��ؼ+�����H�����Q.��I��*g�r+��R���������	���bR��=��UM��4v��`�.T��S��^��s��ц��x��lO���A���C��2\��K?��T�k�o�M�H23�~r����/� ���񼵽缺'⼞�Ϳ�RT伈�뼂����>O� i$��;�t�W�Fv�����|W��Dv���\��w:���]���5�������t��Jb���Y���]���l�����}���#��l��[|��!���oџ�к��S��Urk��N��5���!�)�ڨ�D��~b��{L��ed��72�������L
����#��  �  $���i�vG��o�[��2�T�D���J�LD��2�����7���̼�����ԣ�q���ټUi��;"��{:�0TJ��N�"BF�R�2���bd�vI���oo����|���T���:��=;ngs;�D�;ի�;��w;ȔI;~�:/�$�_�J�""�u�N����Z;ܼBf��j,�t6D��&R���S�{[I�O�4��.� @����Ѽ����6R���hμJ-��oy�)t2��!H�?T���S��zG�4�0�����缒䩼��f�R�?���'��7Ѫ���l:��:��:x P:[�7�9���F�a5��w1�2�g�4)�����^���u2�ɱO��je��Zp�J�n�5�a�C�K�[{1�����������D�����'.�:K��;f�lWz��ȁ�H��X�p��fX�b�:��6������Pɼ����R脼cc�S0L���@�:�=�"iA�YJ�Q�X�M9o��/��I���K"��}�� ��*�.��O�^^o�N(���I��x����Ύ�>x���t��Z��C�ڽ4�\1�`o:�fN�~wi�9��揽`V��.�8��������b��D�f'(����E���I��f�ռ!x̼xpȼ�*ȼ��ʼyaϼD>׼�W�!��H6�����/�e�J���i�K������럽�צ�⫧� U����1���z���c�U%W��sV���a�Uw����Ț��#t���u���`��m'��Hו�#5���xn��mO�k�3��l��T�U- ���	漤�༡�޼�]߼���J�鼀���mM����f�$�E�<�AnY��Oy�ۭ���욽bk�������[���J���̖��:���x�0te��\�ړ`�Rp� ��鑽bힽM{��M������p������"׆�_�m���O�� 6���!��]����s� �n��������
��)���Uy��� �g@	����9#��  �  \���d���*뼉���_-�oy>�_D�E#>�!+-�������Ƽrަ�J����S��{�ѼW�w#�~�4�D�	@H�H@�l�-�>���86���Yk�/�|����ҁ�\��:e�/;��f;`;�>�;�k;�<;<_�:����S� ��ZtL�������ּR�
��'���>�}�K��M��UC�LH/�|��Mm��P_˼7���]l����Ǽ0�����-��(B�#�M�*�M�'�A���+�;��⼹�����c�ψ�/���t�����ސ7:�:��:�T%:�^%�M���T�[1�����p)g��J��u�ݼ���G.��J�w|_��j�ŗh���[��eF��-��������A�v��n*��FF��`��;t�{@}�
z�l]k�	�S�?�6����.���mȼ����5����f���O�h�C�/�@��D��L��[�}�r�e艼��������c��c,�L���j��m��0>��8~������0����p�V�� @���1��t.�U7���J�A+e���������;���ɗ�N>��"O���}���_��B�0%'����ac��7��v׼$Bμʼ(�ɼ
�˼��м��ؼ+�����H�����Q.��I��*g�r+��R���������	���bR��=��UM��4v��`�.T��S��^��s��ц��x��lO���A���C��2\��K?��T�k�o�M�H23�~r����/� ���񼵽缺'⼞�Ϳ�RT伈�뼂����>O� i$��;�t�W�Fv�����|W��Dv���\��w:���]���5�������t��Jb���Y���]���l�����}���#��l��[|��!���oџ�к��S��Urk��N��5���!�)�ڨ�D��~b��{L��ed��72�������L
����#��  �  � ��{ Y�}���ݗؼ�]��2�r-�5�2���,��.�\���Lݼ�+��@����`������oA��B�뼒��tU$�f�2�ɉ6�0�/����Ns���ؼZ���Z�a�����f��+CӺ�:��;��=;':Z;�%\;��D;P�;MUk:Ŋ��iu����fG�i��%�ȼ{9 ���Q�.��:���;�T2����bD��-༪���(ơ�����%Z��\�ۼ<����ZJ1�*<��*<���1�����=Ӽ�᝼��]����oE��G+1�F���(�B8(�:S�:\�8�fF�U�����ӻ� �B�g����y�ӼgY���"�<���N�%WX�o�V�:+K�@�7�b� ���
�\��2��W�����U�8���P�k c��~k���h���[���F��X-��v��e�9�Ƽ>g���Ԋ�*)r�KA[���N��9J�{M��JV�5Df�O~�����[̥�>5ü��j���[&���B��Z^��u�θ��q���Q	��YMw�1b��J��;6�v)�40&�:�.�i�@�<�X���r� ߄�t}�������닽����Oq��W�(�<��$�4���U�Id켨Vݼx�Ӽ'DϼYYμ�м�ռ"{޼�뼋k��u�	��t��B-��+E�:`�t�{�슽!���
��P����Җ�1�������nk�B.W���K��K��pU��h�YQ���\��
��}q�����34��j{������<d�xI��1��\��9��o����9�3����\�va��4񼷉��_������$� �9���R��n��߄�s*��3��k����i������݌�^Ā��zj��JY��Q���T��b�%cx�z���(?��vʜ�����w랽���T���=��*e�wEK�(�4���"��Q��}�p��X ������������*�������Z	�2�$��  �  H5�/N�R	��˾���뼒��0�����R/�|� P������s����v�&�h�k뀼 l��C�Ƽ-P���ĺ�����r�"
��5�Oe¼/����Z�������Ae>���Y�'Y7:u��:�-;�];x�:ԕ|:�,비)�����/�lG�������0�,����H=!���!��;�E	�~���߾�OM���g��"i��e���������o�X`�"���"�6V� �
�9o�ӿ��m���m[�]��W�лeɃ��X���</���
�~�|�s.���$Z�0Ŭ�K���wX1�ʂo��.��Yȼ�%��O��[�'��7���>���<��2�3�!�4��ͤ��ڼHϼ�׼�k�sB�# $�X�9���I���Q��P���E�X5�qa ���
���}UȼG���ݔ��=���q��gb��P\��Z^�,h�0�y�ȿ�������ﯼ�lʼ[�꼪��j��8[6��L���_�.�l��2q�.{l�ƙ_��3M�:9��g'�q�>���A!�Y>1�o�F�7�]��q�G�t�����Ls�b
a���K���6��#�o���y� �������޼ټ�f׼g�ټ�I߼�輬7��������j��5-��A��$W��m�Uw�������g�����5H��C'���o�|pZ��I��?��>�\�G�@DX�w7m�q�����hp��Ǝ�y��� Ă�#q��Z���D��*1� � �-u�1	��d������m��]�q0����5����Y�R��P�՟&�<8���L�Xac���y������H��F���
w���݊�rY�n���Z�6�K�)E�dH��?T�Jg���|�܉�����ܔ���y��b���\��}s��2]�(H�r�5��\&�'T�f��#
��T�������������G����d'��t(��  �  r	��P�r��j:��&�Ǽq��(��d�������\Ӽ`�������b�:�8�~X-�EB��Xs��L��=|����߼ɞ���E����������̼ͭ��?���`���+�����Lt���:K�����rg��:G�!:,u�8���j�-��ᙻ�軕�!���U�����짼9Mȼ���������������|ܼ���}9��0?u�yJT�9�R���p�o��RԶ�N�ټŕ����h��� �B����μ�t���Y����g���5�YK�s�λ�̓�eO�0�����,���r�)n�������.$�S��Ƀ�v;��|���0���������>�w!����G��o�����<м�ι�Z=��_߸���ϼj������,���3��4���-��F"���� ����뼏rѼ����	N��:���*��B	����x�.�y�c4���x��:���P��;b¼Oڼ����FV	�4��э*���:�`)H�\�P��YS�|�N�r�C�D�4�c$����ڟ�8�
�ew�����1��KD�ziU��~a�e�f���d��\�#UP�Z�A���2���$��f�P��g��w����{��Ƞ�y�"��J���5�Z����#���0�2�?���O��_�T�n��*z�����B��Qw��wi��)X���F�=8���/�sz/���6���D�@0V��g��v��~�aJ���n{��p�Yfb���R���B�0N4�Gv'�P�`��`|
�7 ��2��'�������nM������ �;�,�gZ:���I���Y��i���w��a���xy��Ty�j�ĜX�
H�&�;�c)6���8�/�B��xR�>�d���u��F��ǟ���h��(逽��u���f�'5W���G�_":��.�Ɉ#����r��C�h�	�����
�"�������Jq%��\0��  �  �(C��Ni�1o��6���
��C���`7��S1��`����������bTI������n߻Sg ��A'���\�͔��Z9��!�� �ļ�ż�񾼦V��~����E����-[���5�(���{Ի�i���7��2��ẩ����}�k���V��#�.��U�.|��ϐ�f.��妴���üdμ��Ѽ�[̼�2���奼����[}\�Ss/�����]�e,�_�W�u{��\أ�����̼ixӼ�>Ѽ`�Ǽ⋹�n����������h���D�� �m���4.ŻZx�������g��	eͻ���^�0��^��ԅ�A曼�3��c�ż� ڼ��0<���5�Um�a �O����ڼ>��TB���a���Y�����ĭ����Ƽ=W�|L���b�xE��������������X��o����ռc�ļ������꧗�A���<ӏ�S��#���k��gɼ/�߼V����Z�t��@��b/#���+��2�ф6�&!6��	1�w�'��[�^s�*l�O6���T��D�
���z*���8�+�C�?"J���K�C�H��MC��#<�:R4�sV,�O$��&�T�����m������t}�������y��m����n���x&���0�~�:��/D��xM��8V�0�]��b���d���a�O�Y�|0N��@�%2���&�(E ������%���0�v�>���L���X�c)a���d���c�4�^�۽W��]O�/�F��x=�VG4���*��/!�r�����I
�t3�!��"�����M�l!%��$/��8�lrB���K��T���]���d�Y�h�Hmi��.e��C\��O�"�A�+�4��+�̸&���(�>�0��4=�O�K��Y���d���k��n���k�Rf��^��lV�}�M��D��;��52���(�����������5��	�j��� ��*��"4�b*>��  �  �ⅼ����8��X0��8����З�/����m���zv���P��!%����㨻�xr��}Y��6���Q��

�k�8���e���V-��՚��|��Ä��2���S&��,X���.��`����`�T�4�(T	���˻����l��n��p�����&�KU�P���Ź��"?m����� 쮼0a��W0���v���9��s���i���;�q���ݻ�����ƴ�X<ػ�;�p8���e�i�����7������W���E鱼�������8����m��I|��ĭo��E�"��U��>��i*�b6��G���y�u ��R���������ϼ�ټz�޼�e�A��%߼��ؼD�ͼ*������!疼�:���r�j9k��v��=��'՟�;���yҼO��������+��y�	���
��
�4��E*��\�����k)ڼ Ƽ��~L��.���v�������ռ�S＂/��
��l�;@��� ��"�q�#�6;#��;!��7�F���J�cY��������Diۼ��ڼ���7+���.�/��j���)���1��7�:;���<���=�Z=�cT;��=7�>�0��7(��o����
u��m	���	�x��-���E#�͡/�f1;���D�`�K�<P�d|R�hS�US��aQ���M��"H���?�̓5�&*�T3�2������m�����q�(��J4���>�tmG���M��RQ��SS���S�*}S�=�Q���M�{�G��w?�S5���)��U�Us��}��8�����"�E�-��C9�ǽC�iL�P�Q�$�U�XhW�hX�pW�nU��~Q��1K�uB���7��,�A�"�k{�[���� ���)���4���@�u�J�(�R�{?X���[��M]�U�]�S]�7�Z�e�V���O���F�� <�p�0�eS'�� ��f��� �ז'��1��#=���H�ЃR��  �  &_��s��Ah�������A��>���Km���I�k�$��+��񻲻U�Z�f_׺�&�����˻q�����a��\mֻIw��V;��b�^��媖�����}��5Cļ_ɼS�ż�a��݉���d��V0W��i(����p��A>���D��{�V���7V����ƼnϼT�μ��Ƽ���4���������Ze�֋?���d��#?����^��&�N$���W�#k���&໢%�pc=�0�c�㘄�P�������/����ȼܦҼ|>ռ�μ�0���0��b�����h��gC���2�t�;���]� g��騼[Gȼ��⼨���T����f�������ּ@�ƼBO��󷥼���3����g���M�3�=��S:��D�\��8~�Ɠ�����@��}oռ���&�����?�����L�����Q�/��ב��"��ؼ��ȼ��ļ[pͼ���\��������|)�X0��&2�)�/�u�*��e#��f�:)�H�
��o�4��[��k�Ӽ0/ȼ�¼ϣ¼�	ʼ��׼�7�!�����
������ �w�*���4�ؠ>��QG���M�.oQ�y�P�!K�T^A��5�0�(��9��T��^�����*���8��G�)&U��^�nc��Wc�[L_���X�VFP��]G��6>���4�K+�aw!�����S�����M��YO��{�9��6b ��<*���3�xM=��F��O��/X��p_��8d�9Ie���a�bqY��SM��J?�9�1��N'�4�!���"�#�)��5�q�C�)R���]���e��ah�/�f��a�nZ�pR�JII��Y@��;7���-�hO$��@�����Q�S"�1^�����'�3D"�1=,��I6�f@�C�I��	S��0\���d�vZk�61o�C�n���i�_Y`��zS��vE��8���/���,�H�/�3�8�p�E��OT��b�f�l��  �  ސ�c�i޼2Tż���5|��}�R����/�ڻO��� ���P��N4�:�k�:��;!�:]�:Ӊ��.H�3���l���8���r�G�����[ؼ���b��~G ��|�ڼ٭��+�����o���J���D��q^�@����諼~�ϼ�=� � �g ��켒�м�����ۑ�V�h���3�>������q�"����Q��D6����@�����Vh�G÷��s�1�qe��A��&��[:м� �2`�Ĝ���<��I�ݼJ��&���p���4p��z������b���ټ���`�����:������"
�������ڼ����U�������n�ˠM���2�s`�������T��v0�U�L��p�Ӻ��@��M��:�ۼ��������J��Y-��7���:�k7��-�)[����&����\��^�-��N�����(���9��F�mM��9L�j�D���8��>*�O�����1���?Uּ�Ƽ�s�����hg��[���A������{мpK�r���ߛ�!L�ؙ%�#76��GG�?TW�'jd���l�n���h�9]�p�M�T�=�Q?0��R(�3�'��/�U�=��O�hXb�d.r�]�|�W��g|��Kr��zd���T���D���5���(����y��A:
��9��}��98�����p���#��DZ	�u�����;'��e4�A:C�]7S��Bc�֨q�,X|�R���3t�C�v��#h��V��E��Z8��x1�J�2�~z;�QJ�[ \�/�m��K{�ډ���⁽��}��hr�+�c�	T��D��p6���)��8�K��������̎���������V�����6(�r4��eB���Q� Ab�&r�"��Bp���ꅽ�׃���|�@m�g�[���K�#T@�� <��@��KK�[�8�m�nO~��/���  �  9��u�������&ֽ�!c��D�O����=U������"�9�F�:�&B;��h;c<p;e�X;�b!;�U�:��C���P�$�λ�T'�%@t����nӼ����U
�,���:��B�Z���較���I}�����.-��%���U��g�ؼ��������Db!�v��`�pa�z�ü�����_�%���Cǻ��a�u{��wb8�s�:b�:�i�:��:��9�'��ȺW�υ���o�_�Y��Ŕ�	��R1��!U�n�#�z�"��z����D�鼎A¼`���Õ�����L���ڼ,�N�"�+�֝5�}6�ˏ-�]����	�������"�����x��UJ���'��������3M�'"�J�m��WT*���J�= t�����H��c2ټ�O�ܚ�|0��RD�UR��>X�)U� UI���7�7o#���r��� �c�{�A�)���@��U��kd�"�j�n�g�pW\���J�ݘ5�^��+�������ؼ/�ü���v�������Z��������1T��뾼Йм���?.���&���<��2T���j��
}�`p��`���(���x�9f�kIR��A�+�7�7���?�˳P�Y@f��d|��}��dL������/H��*
��'At�h�]��G���3��H"��X�l	�D�ϯ���{�{Y鼑 �(��4���9 �N\�^��� ���1�o�E���[��Ir�9e��p.���8������ŉ�i<��n�m���X���H�@w@���A��sL��T^��s�tD��S�����,-���f���!��kq��[�/�E���2���"�,�,s������������c�����k���f���z,�_����.�NA��+V���l�_���9S�������dȒ�����<���Sq�Z�]�rP���J���O��,]���p��F��2!�����  �  ā0�l[+��6�$���ּ���/�Y�X��gx���%�'�:��P;lN�;�^�;2�;ِ;��q;� ;&U :!���<���b%�����@�����v���P'���4��B8�&�0���������fo�����6��	ժ�9ϼ����,���n,���8�;��>2��& �	����ؼޡ����c����g��k����ǒ�:��;�/*;2�*;�;ķ:i�:8�8 �8��g�Z�\�N���]�Լo��F��2�1=�F�<��32��C�-���`⼁_�������7��v�ϼ?w�����A,1���D�V�O�U5O�|(D�\�0�ͭ�����x�Ƽ�6���l���6�X?��U�6%ջUdʻIλ�߻o�������4��>_��ы�A��!Kݼ���4%�u!A��dY���j��'r���n��qa���L��5�0R �������n�$�G�;���U�`Wm�~��W���"��=�q���[���A�=�&��-�Pa�
pѼ�Y��Hר�^e���ޘ��u��E������Ho��K#����ż^
ݼ��������)��D���a��|�7���P�������ޏ�;���kz�ԅc��1P��D�g�C�-�M��`�h4y�8=���͓�BI���u���"������恽�dh��6M�4�4�U � �������F;�o 伟�༒]�k��.꼣V�����x���'62�zrJ�.�e����^;���ۖ�����?����*��Bi��*i���#i���V�h	M��|N���Z�%o�A܃�&����꘽����Ɯ�����z���C�z�c���I�{{2����Y�����?�������l�t�����F����j����:���T-�0C���\��{x�����ؕ�84��9�������8���ꍽ����H&m��\]��wW��\�$+l�8N��ȍ�����栽�  �  �EB��O<��A+����R輰)���e����cab�mB��;�R~;�#�;�-�;��;��;�%�;=�N;�K�: 麺8ݫ�S�(�1凼�ü� �ׇ���6�n6F��J���A�wN/��N����`�ʼrܮ��䩼;����<���W�&�=���J��L�ЬB��[.��������3���dk���P����|º�':��;��7;p�N;O; �9;�	;"�E:����.l
�_$c�Yr��h��l��)-���B��N���N���B�i>.���������Ѽ�<���żS�o��(%�)�@���U��Ma�N�`� �S���=�(�!�����Rμdm��#i�G+.����ڻ@w���󶻋$���m̻�����	��;)�%LU�6ψ����9h�f\���-��M��/h��o{���*����q��L[��A��*��z��;�!��.���G�Y�c��b}�򱇽5������Yd��h���J�տ,��H#�
�μ<|��9������R���TΒ����)���.��:v������ؼ�������-��iK��ak�[焽.x��	�������}���ޏ����	o���Y�IM�TL�3�V��Gk���騐��!��6!���H��d\��u<������hp��R�ǜ6����k3�<d�B"���a�޼�ۼ=�ۼ�u޼i�伧��@5 �Љ������3���N��/m�=���/������ä�����0���s퓽Mچ��s�I�_�]iU��V�Z-d�az�ԋ���}��Pt��}r���s��"������8���F�j�tPM�2�3�����1�k ��v��kV𼣓�%$�q�|��������0h��w��|-�ߢE��)b���������;������!����k�����d��tՇ�Xw�}0f���_�@xe�-v�vD���Ԕ����ߜ���  �  ��ʽ�dŽ�Z�����`���V��k%����򞳼�n���<�����/7û���-�̻T���q�S��"���ȼ��=�4�2�g�厽)����彽�9˽�wνi*ǽ\ⶽ����5艽k�l���T��P���`�I��K��!���<	½@�ͽ��ϽI�ƽ�紽�뜽=7���O�4s ����20���ˆ��N�� %�_�&� �� ���
���!�%I��Â�����]�W���XJ���~�7��ǲ�ڟŽ��Ͻ*�ϽEŽ���y-���8����j�~6Z��"^��v��莽�ᦽ@���eнX�ٽ:�ؽ�!ͽj_��4���V��w�Y���-�Z�	���ݼq뷼Q�����V����=���A��c���z��=�ļ�꼥��9�0�g[�֘��x������)�ӽ�X�Bc�2��M�ڽr�ƽ�����j��X6��C��x����m������@ʽj�߽t/�N�����ｃ:� @˽/d��Y����#}�ʱS�6�2�w���
����T�4�&�Q���?����� ���/��-L�uq�"������lĽ��޽�'���� ������<}�JRڽ�	Ľ�T��S�������'���k���ս���4 ��4�}����/�󽳜۽���Pk�������u�n�V���?�L�/�.9%�������0���Q��!$�$.�3/=�{%S��2q�/��P��̊��vؽP
���_������x��J�kkٽ�ý&�������A���20���5ȽyQ߽������l��O ��� �\�� �Խ�������ݽ��o��$S�?�ԃ1���(�$�j"�Yq#�EV'���.�Iq:�|�K���d�b���֗��p���J˽������g��~
�6 �Y�9� 
׽'������K����L���y��Zcս%����|��  �  :]Ž�F���ɱ�|Y���1��z�R�zo#����J���#烼�_B�������L�λ�aȻmػ�} �R�#��0Y��]����ȼ�D��)2�$xc��؋�����=/��TƽhɽP½�2��n윽ȉ��W?g���O���K��O[���{�܎���������ȽDʽ��������7t��Mi���L������`ӵ�����F�T�ކ+�c_�L^�P�����(�m�O�;���MN���\꼀u�zkG�D�y��ږ�d�������|ʽ�1ʽ,��3:��6a�����Yte�'bU��>Y�[�p�����[ܤ��EJ˽�tԽgӽ[Ƚ�Q���c��݃��W�s�,�A
�i�߼:꺼�^���������{��������������Ǽ�켪���0�?�Y��҄�����6Ӹ�*XϽ�E߽D�(���ս0h½�g���o��ॊ��څ��������t����Ž�۽���ܓ�j�꽷�ܽ�{ǽ��������({��)S�)w3����"��4+��b�������S���Ho�3��?�_�0���L��@p�b�}�u_���ڽp�+����0 ��������5Eֽ����Z��������������N��SUѽ�;轆m�����w�rA �iN�D$ؽ�R��	ڤ�mꍽ�uu�`VW��A�$O1�W�&��l ��W��%������%�p�/�?�>��T�1q�,M���١��#���ս{�콅����S�~�������ћսeۿ������P�������k��C�Ľ�Z۽�5��b<��b�g-����齂_ѽ����ٞ��@���=o�1T���@�^#3��x*���%�a�#��$�>�(��J0��<�\CM��ge��Â������Ƚ":�Ǌ��T�f`��z���0��tӽ)ﾽ؎���&��>ï�P���0�ѽV�轋^��A���  �  X���������Ow��9I�0������a���Ry��ַV��"(���	��*�.��E���,��58�A"m��P��?�̼���jj,�#�X�k����ʙ�j	���u������v��v���Qz����y��4W�Y�A�)�=��GL��Cj���������������~]��:泽�����4�q�˪D�������2��~���g�i�'�?�fQ%��[�u��Q#�?<��Md�$��x!��}:켪��q@��m�����*΢��������=��'豽v���𛍽�9t�KKV�ܝG��NK���`��M��ȿ������伽�tŽ2�ĽQ�����/ϔ�,|�0�P��*�D��á�	�ļ�Ĭ�Q���V���a����)������ⷼS�Ѽbs��3��U0�aaU�<��:���j���v�½ѽ�׽�ӽVȽJT���9������W���}�wჽ_6��*������{�ͽ�A۽ ���ܽ��Ͻ���Z馽m8���zv���R��5�8A �J���K�l �Ա��P������N�z���.!��4�;VN��n�*��7q�� ��k�ϽG�b(�*R�T�/�ݽS�ʽ����p���q���'����et��v�ƽ1�۽�\�m'��P��t��uJ㽺�ν�����ڠ��O��<v�#�Z�ѫE�y6���+�(%�^�!�|�!�ā$���*�8�4��\C�sW�	r������$�������˽��V=����+C��Һ��!߽��ʽ۶��Y��#a��J������ň��н#'�՜�3q�����.���u޽��Ƚ��������#X���p�H�W��E��Q8�n/�C9*� J(�(h)���-��h5�'%A�b�Q��h������ה�-��.8��� ؽ�콂������"/��e�E�ݽFɽt��>���E������J;����ǽ|�ܽ��ｓ���  �  [i��4���8�����b�1�=�a�� ��!�Ƽ�l����}�5HN��6-���� O�� ��78�U�^�������Jؼ���B�&���J���p��v���6��S�������b���u��pQ]��"?��x,��)�n�5���O�jTr�l$��7M�����������៽����悽��`�5�;���|����T˼q���Sd��@e���G�f�8��28���E��Ea�K���&.����Ƽ������K�7���\�����:��QM������U��f��mێ�F#{��iY���?���2�Z6�IsI�p�h�����`��1���	����|���觽�^���7����m��xJ�&9+���	u��7ؼ<<���ѯ��Ӧ��$��͑��O��.�ʼ���+�����3��*R�ߪu��鍽F����������(���	��hƳ�/g�����P@��g�p��Ri�zr��Ą�0���ao��O���s�Ž�ʽ��ǽ�ڽ�ᰮ��Ŝ��d����r��T�)z<��:)�Ї�������ڏ�q����	��=�1@�=�*�T7=�MT�~�o�IA�����r�.L���nϽI�ؽ�K۽H�ս��ɽ��������LW��պ��+�������1���޶�F2ɽ��ؽ
<�	L�6�޽�Fҽr����㮽�\���u��A�y��b��O�8B@� 35�e�-�W�)���)��-�C�3�v�>���L�N_�r�v��s���������Q���sнݽ�:�5Q㽬�ڽ�Z̽벺�ha���㛽>������؂���h����н�_޽�r�����ܽ�ν+���w��r���ш���&v��[`�&0O��B�\�8�e�2�i^0�`�1��p6�$�>���J�|�Z�Oo�W���A��x���-���&ʽ�Hڽ�����~q�1�۽��˽J��w���?��T홽����$������3˽�۽�_��  �  mW��%�^~��-i���O��m5��4��H��ἊA���I��q{���5d��#M�hG��bS��vp�[T��#���t�˼��D�~R&��@�_v[�Q�t������~���ފ�;D����t�6�X�kL;�g["�����(�	��V0���L��j��-���y���������KP��`�k�SSQ���6�=�o��q�輎ƼgE����h}� �j�\�i��Jz�f����f���¼������/��W4��N��-i�,����o��্����>ʄ���q�1U��{9�|J$����;� ^-�T�G���f��ӂ����O��Pv���ڒ�������{�%b���H���1�\v�Ͳ�����%�߼T̼���������üR:ҼԵ�b�������&���<��tT�q�n�����Y���ĝ�����,���㤽����L��m��;*h�HdV��P�X���k��������������2��������"��Rȟ��R���Z��;�s�Ѭ]��J��$9�T�*�P��Z��A!������2�>�+���:�ٳL���`��
w�@����a���0��o.��ϼ���!��K	½�
��
첽r���&����ދ�1���	)��4��`������i��u��K�ȽƗ˽FȽ����Yf��C?������샍�'I����p�U?_��/P�]�C�;��b6�6��;:�̉B�dgN�/]�;n��ွ��7E��6����Ʋ�f���9�ǽX�˽�ʽ��½�N������~S��,��5n��yF��,����Ӝ�V����2����Ž�0̽��̽��ǽ[��ٱ���������>Ջ��8����o��u_���Q��F�|�?�
�<�%+>��	D���M��[���j�Q}��Ј�pm���9��o���,ͻ��ǽՑν��н�Oͽ3Ľ�޶��������!���������Zڙ��T���o���GĽ�Tν�  �  ��]�6 `��C[�+VQ��lD��6��<'�����/���u#ϼO�������/T���K��8��ɟ�_麼�ۼ�����I�����B/�@�>��GM��@Z���c���g�^wd�kY���F��/�#�}d�4v��,�3������=t&���>�H�S�� c�Y{j�d�i��c�i�W�,J�4W;��',�b��@Y�`t���ּ����˓��V[����������-����Ӽ��m�
�����*���9�x�H�S�V�u�b� �j�oll���f��X��#E�R>.��h����|) �p��!�EI%��>���W�[%m��G{����x�&�w��\l��_�E�P�)sB���3�0R$�?��L`������伿`߼y�<"����	��z�|z,�yt>� �O��j`�0�p�l ��J���Ì�������������6���s�L�\�V�H�s�:�Ǣ6� �<���L�۫c�`)}�҇���֓�dX��zĚ������䓽
���Y������cp�UTa��Q�ޚB�_�4�I�)��o#�-�"�{(� �2��A��S��1e�qw����Z���b�����I䢽�����Y���?������쐽�녽t�y���n�Vn��w�����$ϐ�-@���1��t ���ϳ�졳�.��(�������L&���u�������[����w��xg���X���M��fG��G���L�n%W�7ve���u�<��n���X��Q��ɍ��E���J���cq���<���*���"�� 럽�����������v�_x��ρ�А���o���D������r��wε�wk��e&�����������;���@���&��|�w�+h���Z��vQ�!|M�OiO��W��[c���r��́�LE���}���p��#2��~����������'��6���{g���A��2]�����o̊��O����������[������=��ǣ���u���  �  ��4�qM=�\DB�i�D�B�D�6�B��r>��Y6�*����q�����ɼ�4��+����๼��Ҽ=*��.��� �t�0�ǜ<��kD���H���J�?�J�^H�AC�r:�Iz-������	�&���м�,�������ǼCN����o���(�m�7�PC�ZJ���M��\O�T�N�h�K��$F�Ҁ<�]�.�}X�H2
�v����Ҽ <¼�\���7м-)�'�xa�g-��];�8�E��K�UO��P�EO���K���E�ݾ;�L�-���ed
��1�Ղڼ�~ϼ �Լ�p鼒l�%��~�.�N�A��Q���[��b�X�f�yh�( h�#e�T�^���T�
�F���5�p�#�:����J��<��@� �%���9��fN��|`�ڧn���x�`�~�5倽Ce��n߀�?-~��Ew�ihl�:�]�%TL���:��++�!�68�>m#��0���A���V�\�j��7|��ф�f��}(������[፽�,���&��Ve������t�	xb��P�FB�K9���7��]>��L���^��ps�����C(��
����ݖ�}r��8���
���I��a,���H���c��۴����{�e�j�%L]���U��NU���\�&Ak���}����̐���\���	����������AH���@p��zo���������������s�� e�;�\��W\�P�c��q�x遽�����o��@���� �<���8����!��z���H���Ԡ�����z��r������Wr�a�d�2^�_���g��w�݄�����cN��{A��� �����)������0}�������B��PӜ�)[��)Z��Xۂ���t�;h�Y�b�6(e��Bo�5�'��/Β��S��?�������VE��0����檽(+��E'���m�������疽j���QR��x�d�l���h��tl�U�w��3������ m�������  �  ���Ԗ&�6���D�	MR���\�ȸa�3�_�C�U��MD���-�nD�q��-輯��N�����8��5���K��*\���d���e�&�_�~XU��H���9���*�:��J������<ռ����a}��}ے�娐�B<���b���nʼ����Y����'���6�	�E��T�`��"i���k�7g��2Z�*�F��/�|��f�������0�Rc��},��7D�l|X��<f�Fl�g%j�a/b�HV��XH���9���*� E�z���:����ؼ�ᾼӬ�2u�����(�����Լ���B���x1���B�fS���b�m�q��}��͂��j��(!����q�p�]��IG��`2��W#�nc��!�t�0�plF���_��Dx�����g2��K�������P���B����v��qh�P�Y��J�HZ;�Z�+�������
�@+	�3u��P���%�ؙ6�X�H��|Z��k��*|���ƽ��������=Μ�A���q���*��8w��Ucr���^�ȱR�j0P�DX��i�x���\������ǡ�e����~���m���,����ْ�͋�����xz��Yk�^\��,O��E�1�?��?�7�E�k"Q�d`�q��L���Ӊ������ڙ��u��d����î�e��QI��Ǳ��B��]��k����̉��J����u��u���~�������'���\!��v��1�������(��*:���?���Ԛ�+7���a��>D���u���e��W���M��H�k�I�>P��[���j��e{��'���d���Z��c�����Ǡ��a���嵽�&���v���᪽IR��^u���e��l<��R-{�<h~��Ʌ����� ��pȧ�� ��Pල������������˫����9O��Ƕ��ލ�⾅�P{�W�k�,�^�:vV�zS�oiV���^�B�k�	�{�=Q��-Î��  �  �g���/�5�/�P�:�j��"���ꆽ�M�������]s���W�h:��c �/)��;
������&�[�B�X�`���{�����0����-�������&k�rcQ��7���v���>�RAļ����O���u���`���]���l������<���ſۼ�!�Y���H/�f�I�
\d���|�c���s���O������+t��3W��9��"��e����r ���6���S�CKq�k��������d��������h��M���3��v�h	����ifƼrR��QV���ሼ����l������E��{�Ǽ�r鼹���V��95�MhO� 	k����������aW��5���0��H���؁m���R�j?�vm7���<��N�*�i�����;d��L�������m������>5�������w�)�^��$H��4���"����7x�����v|�i��#��=�"������/��C��dY���q�h���Г��젽oܫ�GᲽ}���[L��೦����@���}�ϯm�5j�2�s������8���좽�ܰ����㥾���������Ӫ�QO��ׅ����xu��b�"yR��D�ɱ9�i2�jR.���.���3���<��FI�τX��j���}��ꉽC-���]��W��������gƽ]V˽��ʽC�ýG'�� ����嚽(뎽;��Ҧ��Xэ��L���ͧ�A}��T�½��ɽ�Y˽cǽ������aۤ�X����������4n��f]��O�߀C�~�;��7�q�8�Ɯ=���F��\S�+�b��bt�VB�������8��Q���|ض��x½��ʽ�ν b˽Ný�G�����;����@��皊�o����䔽�ѡ�?ذ�9����ɽ�sϽ�Ͻɽ��������V������d挽����l�r���b�s�U��LK���D��B�8�D�2�K��V�԰c���s��<���  �  �����#��>��d�������V��'k����������K����l]���=��)��#��,-�hoE�^g���������%+��Aw���������f���y{b��p=��K����u�ʼ���Nׅ��M^�Sg?�7�.��,�P�8�d�R�j{�on���'���,꼿���\1��U�7�{�]e��\K��3��ה���B��ۓ��JX~��Z�_&>���-���,�ī;�FiW�@nz�#ڎ����4G���ϥ����\z���G���%[���6�b'�0:����ȼ�'�� ��<~s��^�Z�W��_�F�v��������lɼ�����1�L�T���z�����l���q5���'���d���C��)���"T���r�"OZ�!SP��iV�g�k�����ʘ��g�������⽽�V���r��!����Y���怽��^��c@��'�Z��~��+���� ټ�gؼ>�޼/��s� �<���7 �h/6�LQ���p��v�����',��yݿ��Pʽj�ͽMɽ���������� ���zÃ�kf��G������=T��9��-�Ƚ��ӽ�w׽iӽ�Ƚ�Ҹ�Ϧ�������K�k��lT��GB��4�c�*�YY$�˪!��w"�]�&�^.�f�9��%H�S�Z���q��ǆ�g/���s��1S���ͽu�۽ł�z�㽙fܽ��ν�)���j��&��������2��9���ʁ������̽��ڽ�-�j��k�ܽj|Ͻ�L�������R��x刽��u�&_�D%M��=?�i
5��w.�L�+�x,��:0�g�7��`C���R�#�e��!~��ƍ�Gޞ�=���+LĽJ�Խ"0��潷��A۽��˽����1��خ������p��8h��x����Ž�"ֽ��L�轉�潄�ݽ
�ν��C������k	���x��c���R��.F�pQ=�f8��j6��H8�¹=���F�D}S��d��y��  �  b	��oz�F�J�nZy��K���n��//��w_���E��|�P����z�v�V�t�>���7�SNC��_�z߂�����'���:����M��K`��^C��`���Tu���G���Mc�����󫑼wd���8��w��,�b_���?I.���T��)��=�����߼���(8���d�D����^��I���蔺����}k���ã�����־v�۞U�ĴB���A���R�-�r�[y��kơ�>���@���Y��K\���䡽����E$k�!|>�V��M�B���"@���q�')O�;�<�^�7�V�?�T��:w���������wo伏���3��I^��y����粽\g½l�ɽ�MȽ/뽽����y���(��p�p��e�6�k����}��O墳�����̽)�ӽg[ѽ�ƽ1���8��tm���d��?�!��>
��|�T�ܼ��μG`ȼUȼDiμ��ڼ�8��ib���/��O��;u�R�������پ��0ҽ�,߽L���޽t�ѽ6����{��d왽/���j���=��6���Ԛ���ʽi�ܽ*h�$>����	ڽ?�ƽ�1���͙��j��rh��CM���8�T�*��!�ہ�d\��E�^!�t#%��/��n>�RR�~ql�ú������H밽W(Ƚk�ݽ)��T������������ͽ%L��q����0�����3/������G˽�߽��Q$���F���Q���߽I�ʽՊ��&&���5��G>q��'W�'�C��{5�|�+�3�%�^g#���#�!�'�K�.��9��-I��{^��~z�<͎�����;{��d�ѽ�/�bV������ix��
�ｪ6޽V�ɽsG��f姽rl���#������r���EֽF���;��<�������^+���ݽ��ǽ�Ͱ��*��^���r�[mZ���H�w�<�Y4�]�/�:Y.���/���4��8=��I��+[���r��  �  A���-n$��T� ~���ӝ��B�������fƽ�����q��fӝ�*T���#g�0M�d�E��R��;p�(��*�>Ϸ�(�ĽYGȽ���}����S��ہ�˛P��"�%W��F��v���|�O�9%$� P	��-������)��a�D�?�^�x�v?���ݼӶ�Z�>���p�>h������@
��TLɽX�ʽ'���t���iܚ������@e���P��O�n'b�j��Vd��^���|`���@ʽ�(ʽ� ���������"�w�_�E��a�e�G���Ɖ��"]�Po;�*��6&��$.���A�BCc�/���歼�j޼�.�QA7�Z�f��`������"��=gн��ؽ?=׽4�˽cc������莽޴���r�z��	���%���w���b˽o�۽}��&�߽�ӽ�྽�V��п����i��0@��/��t��ҼA-żh8���t��Tż�&Ѽ
��&���P4�k�-���O�*6z�4����ۯ��cɽ�߽���L����	y߽�R˽?Y��|'��䶕������q���-���ؾ�U9ֽ����4��-�������`��sнm\��56���\��ah��bJ�>s4��o%�������C������i�� ��t*��9���N��j������ԝ�=ٶ���н=*�^h��P��bf����������ؽ��½���0��;���m߮�R5���1ֽ�_��9��R��	�G���|�뽖�ӽ�˹�{����t���&p��S���>�M0���&�MD!�p���m�n�"�ތ)�k4�>�D��i[��z�Q��������[��@<۽�P�Z��������������a1Խp���[���Q���A��C����˽���.*���i�
��"#��6�� ��Z�Ͻh"���睽��p��^V��C��c7�(r/��%+��)�o+���/�N8�u�D�)�V�`cp��  �  ������&�W�X�0a��~����ݷ��ƽ�˽�,ƽ�9������Ί�<�l�|R�1^J��2W��@v�~ǐ��:��-����ʽ�ͽƽc�������-T��#�m���R��������I�Գ�?>����-�� ����Qd9�7�r��8��s�ܼ3���]A��/u�E���\ծ���½j�νr�Ͻq�ƽ�P��Fɞ�t뇽ͽj���U�J{T�čg������=��\���nŽ�Ͻ�oϽ��Ľ纱�����d|�H������鼊=��������V�G35�K$�έ ���(��<�v�\��b���9��'�ܼqe���8���i�q��(��`pýWhս�=޽��ܽ��н�Ž��9��!����y��U�w�G�T������?����н���c4轊�2�׽/�½�T���Ǝ��k�0�@�ѥ�	��d漄[ϼ�¼S��c����t¼yμq��C���-�?�P��K|�م���*6ͽ��Ʒ�����A��yϽ�Ҹ�����:��`���p��(-��lt½Ղڽ�ｦv��� �M������CԽS���럽�6���h���I��3���#�'H�p�nQ��M�E������(��8�r�M���j�gA��#%�����tԽwC�� �}j���]���]�i�ܽD�Ž>��Z������a���hýGڽ���ģ�w�����j����~�ֽ%��,!��o���p���R�Y=��.��;%����t��Q� P!�^�'�3�2�7C�֢Z��Kz�WK��7S��3�ý'�޽�����&�(b��U��H������׽z½B�����������{��W�ν���"���� ���	����� �x����ҽ�)��D	��'T��0�o�?9U�1gB�Z�5���-��)��{(�c�)�n.�Us6��C�.�U�i�o��  �  A���-n$��T� ~���ӝ��B�������fƽ�����q��fӝ�*T���#g�0M�d�E��R��;p�(��*�>Ϸ�(�ĽYGȽ���}����S��ہ�˛P��"�%W��F��v���|�O�9%$� P	��-������)��a�D�?�^�x�v?���ݼӶ�Z�>���p�>h������@
��TLɽX�ʽ'���t���iܚ������@e���P��O�n'b�j��Vd��_���|`���@ʽ�(ʽ� ���������"�w�_�E��a�e�F���Ɖ��"]�Ho;�*��6&��$.���A�(Cc� ���	歼�j޼�.�EA7�N�f��`��������6gн��ؽ:=׽0�˽`c������莽۴���r�z��	���%���w���b˽t�۽���,�߽�ӽ�྽�V��׿����i�1@� �/��t��ҼI-żm8���t��Tż�&Ѽ �����H4�b�-���O�6z�.����ۯ��cɽ�߽���G����y߽�R˽<Y��z'��㶕������q���-���ؾ�X9ֽ����4��-�������`��sнt\��;6���\��#ah��bJ�Gs4��o%� �����H������i�� ��t*��9���N��j������ԝ�=ٶ���н=*�^h��O��bf����������ؽ��½���0��;���m߮�R5���1ֽ�_��9��R��	�G���|�뽖�ӽ�˹�{����t���&p��S���>�M0���&�MD!�p���m�n�"�ތ)�k4�>�D��i[��z�Q��������[��@<۽�P�Z��������������a1Խp���[���Q���A��C����˽���.*���i�
��"#��6�� ��Z�Ͻh"���睽��p��^V��C��c7�(r/��%+��)�o+���/�N8�u�D�)�V�`cp��  �  b	��oz�F�J�nZy��K���n��//��w_���E��|�P����z�v�V�t�>���7�SNC��_�z߂�����'���:����M��K`��^C��`���Tu���G���Mc�����󫑼wd���8��w��,�b_���?I.���T��)��=�����߼���(8���d�D����^��I���蔺����}k���ã�����־v�۞U�ĴB���A���R�-�r�[y��kơ�>���@���Y��K\���䡽����E$k�!|>�V��L�?���@���q�)O�&�<�C�7�4�?���T�T:w�߲������Po�y���3��I^��y��󝽵粽Pg½a�ɽ�MȽ&뽽����t���(��l�p��e�8�k���~��U墳�����̽4�ӽs[ѽ�ƽ>���8���m���d�?�,!��>
��|�i�ܼ��μO`ȼUȼ?iμt�ڼ�8��Yb���/��O�;u�F�������پ�|0ҽ�,߽@����޽l�ѽ/����{��a왽-���j���?��:���ٚ���ʽq�ܽ4h�/>����	ڽL�ƽ2���͙��j��#rh��CM���8�c�*��!���m\��E�d!�x#%��/��n>�RR�~ql�ú������H밽V(Ƚk�ݽ)��T������~������ͽ%L��q����0�����3/������G˽�߽��Q$���F���Q���߽I�ʽՊ��&&���5��G>q��'W�'�C��{5�|�+�3�%�^g#���#�!�'�K�.��9��-I��{^��~z�<͎�����;{��d�ѽ�/�bV������ix��
�ｪ6޽V�ɽsG��f姽rl���#������r���EֽF���;��<�������^+���ݽ��ǽ�Ͱ��*��^���r�[mZ���H�w�<�Y4�]�/�:Y.���/���4��8=��I��+[���r��  �  �����#��>��d�������V��'k����������K����l]���=��)��#��,-�hoE�^g���������%+��Aw���������f���y{b��p=��K����u�ʼ���Nׅ��M^�Sg?�7�.��,�P�8�d�R�j{�on���'���,꼿���\1��U�7�{�]e��\K��3��ה���B��ۓ��JX~��Z�_&>���-���,�ū;�FiW�@nz�#ڎ����4G���ϥ����\z���G���%[���6�b'�.:����ȼ�'�����&~s��^�4�W���_��v��������lɼ���c�1�*�T���z�w���[���`5���'���d���C�����T��|r�OZ� SP��iV�p�k�����ʘ��g�������⽽�V���r��3����Y���怽�^��c@��'�r��~��+���� ټ�gؼ7�޼��f� �*���7 �N/6�.Q���p��v�����,��gݿ��PʽZ�ͽMɽ������������xÃ�jf��I������ET��C��9�Ƚ��ӽ�w׽)iӽ�Ƚ�Ҹ�,Ϧ�#������k�k�mT�HB�1�4�u�*�hY$�ت!��w"�e�&�^.�j�9��%H�U�Z���q��ǆ�g/���s��1S���ͽu�۽ł�z�㽙fܽ��ν�)���j��&��������2��9���ʁ������̽��ڽ�-�j��k�ܽj|Ͻ�L�������R��x刽��u�&_�D%M��=?�i
5��w.�L�+�x,��:0�g�7��`C���R�#�e��!~��ƍ�Gޞ�=���+LĽJ�Խ"0��潷��A۽��˽����1��خ������p��8h��x����Ž�"ֽ��L�轉�潄�ݽ
�ν��C������k	���x��c���R��.F�pQ=�f8��j6��H8�¹=���F�D}S��d��y��  �  �g���/�5�/�P�:�j��"���ꆽ�M�������]s���W�h:��c �/)��;
������&�[�B�X�`���{�����0����-�������&k�rcQ��7���v���>�RAļ����O���u���`���]���l������<���ſۼ�!�Y���H/�f�I�
\d���|�c���s���O������+t��3W��9��"��e����r ���6���S�CKq�k��������d��������h��M���3��v�g	�}��cfƼhR��DV���ሼ����l��귕��E��G�Ǽ�r鼗���V�|95�#hO��k����������NW��$���0��<���ām���R�j?�um7���<�'�N�;�i�����Id��]��������������T5��-���'�w�R�^��$H�4��"����Jx� ����|�l��#��3���Ь���/��C��dY�ѷq�S���Г��젽Yܫ�3Ჽj���JL��ѳ�����@���}�ȯm�5j�8�s������8���좽�ܰ�����������#����Ӫ�gO��텑�-��:xu�7�b�AyR�1�D��9�|2�zR.���.���3���<��FI�҄X��j���}��ꉽC-���]��V��������gƽ]V˽��ʽC�ýG'�� ����嚽(뎽;��Ҧ��Xэ��L���ͧ�A}��T�½��ɽ�Y˽cǽ������aۤ�X����������4n��f]��O�߀C�~�;��7�q�8�Ɯ=���F��\S�+�b��bt�VB�������8��Q���|ض��x½��ʽ�ν b˽Ný�G�����;����@��皊�o����䔽�ѡ�?ذ�9����ɽ�sϽ�Ͻɽ��������V������d挽����l�r���b�s�U��LK���D��B�8�D�2�K��V�԰c���s��<���  �  ���Ԗ&�6���D�	MR���\�ȸa�3�_�C�U��MD���-�nD�q��-輯��N�����8��5���K��*\���d���e�&�_�~XU��H���9���*�:��J������<ռ����a}��}ے�娐�B<���b���nʼ����Y����'���6�	�E��T�`��"i���k�7g��2Z�*�F��/�|��f�������0�Rc��},��7D�l|X��<f�Gl�h%j�b/b�HV��XH���9��*�E�x���:����ؼ�ᾼ�Ҭ�u�����������ԼN���A�����w1�|�B�7S���b�<�q���}�x͂�tj��!��t�q�T�]�zIG��`2��W#�lc��!��0��lF���_�Ex� ��|2��*K��ɯ���P���B����v��qh�{�Y�D�J�iZ;�v�+�.������
�A+	�.u��P�y�%���6�9�H�j|Z�Ũk�Y*|�������� ������&Μ�,���q���*��*w��Acr���^���R�j0P�DX��i�����'\������ǡ�z����~��7�����E����ْ�.͋�����)xz�Zk�}\��,O��E�C�?� �?�A�E�s"Q�i`��q��L���Ӊ������ڙ��u��d����î�e��QI��Ǳ��B��]��k����̉��J����u��u���~�������'���\!��v��1�������(��*:���?���Ԛ�+7���a��>D���u���e��W���M��H�k�I�>P��[���j��e{��'���d���Z��c�����Ǡ��a���嵽�&���v���᪽IR��^u���e��l<��R-{�<h~��Ʌ����� ��pȧ�� ��Pල������������˫����9O��Ƕ��ލ�⾅�P{�W�k�,�^�:vV�zS�oiV���^�B�k�	�{�=Q��-Î��  �  ��4�qM=�\DB�i�D�B�D�6�B��r>��Y6�*����q�����ɼ�4��+����๼��Ҽ=*��.��� �t�0�ǜ<��kD���H���J�?�J�^H�AC�r:�Iz-������	�&���м�,�������ǼCN����o���(�m�7�PC�ZJ���M��\O�T�N�h�K��$F�Ҁ<�]�.�}X�H2
�v����Ҽ<¼�\���7м-)�'�xa�g-��];�8�E��K�UO��P�EO���K���E�ܾ;�J�-���_d
��1󼿂ڼ�~ϼ��Լ�p�wl���[�.�'�A��Q�S�[���b�&�f��xh���g��e�)�^���T���F���5�Y�#�*����H��A��@��%��9��fN��|`��n�΅x���~�N倽]e���߀�o-~�'Fw��hl�]�]�BTL��:��++�!�88�8m#��0���A���V�;�j��7|��ф�f��d(��⋍�B፽�,��h&��@e������at��wb���P��EB�K9���7��]>��L���^��ps�Ѱ��W(������ݖ��r��R���3
���I��y,���H���c�����{���j�;L]���U��NU���\�.Ak���}� ��͐���\���	����������AH���@p��zo���������������s�� e�;�\��W\�P�c��q�x遽�����o��@���� �<���8����!��z���H���Ԡ�����z��r������Wr�a�d�2^�_���g��w�݄�����cN��{A��� �����)������0}�������B��PӜ�)[��)Z��Xۂ���t�;h�Y�b�6(e��Bo�5�'��/Β��S��?�������VE��0����檽(+��E'���m�������疽j���QR��x�d�l���h��tl�U�w��3������ m�������  �  ��]�6 `��C[�+VQ��lD��6��<'�����/���u#ϼO�������/T���K��8��ɟ�_麼�ۼ�����I�����B/�@�>��GM��@Z���c���g�^wd�kY���F��/�#�}d�4v��,�3������=t&���>�H�S�� c�Y{j�d�i��c�i�W�,J�4W;��',�b��@Y�`t���ּ����˓��V[����������-����Ӽ��m�
�����*���9�x�H�S�V�u�b�!�j�oll���f��X��#E�M>.��h����o) �_��!�,I%�˲>���W�4%m��G{�����w���w��\l��_��P��rB�Z�3�R$�#��7`�����ފ伻`߼��R"����	��z��z,��t>�(�O�k`�_�p�� ��c���Ì������������6���s�b�\�e�H�|�:�ɢ6��<���L�ȫc�G)}�Ç���֓�PX��dĚ�w���䓽񦍽A������cp�/Ta���Q�ĚB�K�4�;�)��o#�-�"��(��2���A��S��1e��w����!Z���b�����a䢽,�����-Y���?������쐽�녽��y���n�dn��w�����'ϐ�/@���1��t ���ϳ�롳�.��'�������L&���u�������[����w��xg���X���M��fG��G���L�n%W�7ve���u�<��n���X��Q��ɍ��E���J���cq���<���*���"�� 럽�����������v�_x��ρ�А���o���D������r��wε�wk��e&�����������;���@���&��|�w�+h���Z��vQ�!|M�OiO��W��[c���r��́�LE���}���p��#2��~����������'��6���{g���A��2]�����o̊��O����������[������=��ǣ���u���  �  mW��%�^~��-i���O��m5��4��H��ἊA���I��q{���5d��#M�hG��bS��vp�[T��#���t�˼��D�~R&��@�_v[�Q�t������~���ފ�;D����t�6�X�kL;�g["�����(�	��V0���L��j��-���y���������KP��`�k�SSQ���6�=�o��q�輎ƼgE����h}� �j�\�i��Jz�f����f���¼������/��W4��N��-i�,����o��্����=ʄ���q�1U��{9�rJ$����;��]-�=�G���f��ӂ�����O��;v��pڒ�������{��$b���H���1�:v����������߼T̼���������üf:Ҽ��w�������&��<��tT���n�����Y��ŝ�0����,���㤽����L��w��I*h�PdV��P�X���k����������������������"��<ȟ��R��vZ���s���]��J��$9�<�*�>��N��;!������2�O�+���:���L���`��
w�T����a���0���.��强��!��^	½�
��첽����2����ދ�:���)��9��`������i���u��L�ȽƗ˽FȽ����Yf��B?������샍�'I����p�T?_��/P�]�C�;��b6�6��;:�ˉB�dgN�/]�;n��ွ��7E��6����Ʋ�f���9�ǽX�˽�ʽ��½�N������~S��,��5n��yF��,����Ӝ�V����2����Ž�0̽��̽��ǽ[��ٱ���������>Ջ��8����o��u_���Q��F�|�?�
�<�%+>��	D���M��[���j�Q}��Ј�pm���9��o���,ͻ��ǽՑν��н�Oͽ3Ľ�޶��������!���������Zڙ��T���o���GĽ�Tν�  �  [i��4���8�����b�1�=�a�� ��!�Ƽ�l����}�5HN��6-���� O�� ��78�U�^�������Jؼ���B�&���J���p��v���6��S�������b���u��pQ]��"?��x,��)�n�5���O�jTr�l$��7M�����������៽����悽��`�5�;���|����T˼q���Sd��@e���G�f�8��28���E��Ea�L���&.����Ƽ������K�7���\�����:��QM������U��e��lێ�B#{��iY�y�?���2� Z6�9sI�]�h�����`��"��������|���觽�^���7����m��xJ�9+����t��W7ؼ<���ѯ��Ӧ��$��ԑ��_��G�ʼʃ�A�����3�	+R��u��鍽X����������(��
��tƳ�:g�����V@��n�p��Ri�vr��Ą�)���Xo��C���f�Ž �ʽ��ǽ�ڽ�ϰ���Ŝ�~d��ύr���T�z<��:)���������Տ�p����	��=�?@�P�*�k7=�hT���o�YA�������@L��oϽZ�ؽ�K۽V�ս��ɽ��������TW��ܺ��0�������"1���޶�G2ɽ��ؽ
<�	L�6�޽�Fҽq����㮽�\���u��@�y��b��O�8B@� 35�e�-�W�)���)��-�C�3�v�>���L�N_�r�v��s���������Q���sнݽ�:�5Q㽬�ڽ�Z̽벺�ha���㛽>������؂���h����н�_޽�r�����ܽ�ν+���w��r���ш���&v��[`�&0O��B�\�8�e�2�i^0�`�1��p6�$�>���J�|�Z�Oo�W���A��x���-���&ʽ�Hڽ�����~q�1�۽��˽J��w���?��T홽����$������3˽�۽�_��  �  X���������Ow��9I�0������a���Ry��ַV��"(���	��*�.��E���,��58�A"m��P��?�̼���jj,�#�X�k����ʙ�j	���u������v��v���Qz����y��4W�Y�A�)�=��GL��Cj���������������~]��:泽�����4�q�˪D�������2��~���g�i�'�?�fQ%��[�u��Q#�?<��Md�$��x!��}:켪��q@��m�����*΢��������=��&豽u�����9t�FKV�՝G��NK���`�M����������伽�tŽ'�ĽE�����"ϔ��+|��P��*�1�������ļ�Ĭ�B���N���_����)������ⷼk�Ѽ�s��3��U0�xaU�<��G���w�����½+ѽ�׽�ӽ_ȽQT���9������W���}�vჽ\6��%������r�ͽ�A۽���ܽ��Ͻ���M馽a8��kzv��R��5�(A �=���K�e �ͱ��O������N�����.!��4�NVN�+�n�6��Dq����w�Ͻ#G�n(�6R�T�8�ݽ\�ʽ����p��r���'����gt��x�ƽ2�۽�\�m'��P��t��uJ㽺�ν�����ڠ��O��<v�#�Z�ѫE�y6���+�(%�^�!�|�!�ā$���*�8�4��\C�sW�	r������$�������˽��V=����+C��Һ��!߽��ʽ۶��Y��#a��J������ň��н#'�՜�3q�����.���u޽��Ƚ��������#X���p�H�W��E��Q8�n/�C9*� J(�(h)���-��h5�'%A�b�Q��h������ה�-��.8��� ؽ�콂������"/��e�E�ݽFɽt��>���E������J;����ǽ|�ܽ��ｓ���  �  :]Ž�F���ɱ�|Y���1��z�R�zo#����J���#烼�_B�������L�λ�aȻmػ�} �R�#��0Y��]����ȼ�D��)2�$xc��؋�����=/��TƽhɽP½�2��n윽ȉ��W?g���O���K��O[���{�܎���������ȽDʽ��������7t��Mi���L������`ӵ�����F�T�ކ+�c_�L^�P�����(�m�O�;���MN���\꼀u�zkG�D�y��ږ�d�������|ʽ�1ʽ,��3:��5a�����Vte�#bU��>Y�U�p�����Wפ��@J˽�tԽgӽ[Ƚ�Q���c��݃�{W�h�,�7
�X�߼,꺼�^���������z�������������Ǽ�켳���0�K�Y�ӄ�����=Ӹ�1XϽ�E߽J�.���ս4h½�g���o��᥊��څ��������t����Ž�۽���֓�d�꽰�ܽ�{ǽ��������({��)S�w3�}����/+��b�������W���Lo�8���?�g�0�ŀL��@p�h󍽃�|_���ڽ$p�1����0 ��������9Eֽ����]��������������N��SUѽ�;轆m�����w�rA �iN�D$ؽ�R��	ڤ�mꍽ�uu�`VW��A�$O1�W�&��l ��W��%������%�p�/�?�>��T�1q�,M���١��#���ս{�콅����S�~�������ћսeۿ������P�������k��C�Ľ�Z۽�5��b<��b�g-����齂_ѽ����ٞ��@���=o�1T���@�^#3��x*���%�a�#��$�>�(��J0��<�\CM��ge��Â������Ƚ":�Ǌ��T�f`��z���0��tӽ)ﾽ؎���&��>ï�P���0�ѽV�轋^��A���  �  �4��0�UH#�k���F����Ƚ-����z���C�Ç�������Ѽ2ʸ�<`��
��L���
���=�ܼ���%�%�LvR�c���+���f!ս��֨�Ns(�٣3��M6�0��""�Ɖ��.���s׽~Hý������̽X�轸���X7+��?5��6��A/�0 ����\뽒���e����p�i>�V��UG��(+ټ>�ü�$��V��������ռM)�������8��i�r���������t	�.�H�-��Y6��6��-��D��
�I���Dҽ2�ý0�ƽ@ڽ� ���b���$��4�(�;��:�5�0����H�
�>)齲��	���Rz�%M���,�S'�c�	�e���� �R�"[�)A��I/�6�M�I0w��
��G~���<�z����q>1�3?�9�D�D�A�616��%����, ��9G߽��罬
 ������%��58�DE�V�I��^E�}�8�$&��X�-q��X�˽י��uy���ut���W�A9E��:���4�X�4���9�˥C�	�S�ٍk�ɭ��ˠ��zk���$�7N����~�1��C�YO��R��!L�ѣ>�x,��t�"�	�Ť��E���M���'l&�+:���J�.�T�3mV�x�N���?���+�zK�7�����׽�������)؊�[{�^i�G^��"Y�L�X�&j]�bvg��*x�����3ۚ��i��+
ӽ�r���p�2�(�k�=��WM�\�U�AkU��WL�Dy<�)��D�����. �2�F�
��s���-���@�S�O���V�mZU�))K�:���$������i�ͽ�ޯ����KK����y���j��:b�h�^��`�Bg�P�s�����%���o��?q��m��H�JE�/z2�&�E���S�z2Y�w�U��AJ�{�8��>%��v���IN��9�����#��J7�lJI���U��  �  ��/���+�e��Q�Zu�u�Ž�]���z���D�"��/����(׼	��$x���,��ڳ�(�ļ�0⼝e��^'���R�兽����|�ѽ�����H�Rp$��9/���1�(�+��2�)�����ҽ�D�����E�Ƚ��㽀��-��E'��0��62��+����\	�������Yf��Up�RU?���e� ��s޼ �ȼ�6������|�ƼP(ۼ�\��j��U:���i��Y��JE���⽚��7p�H�)���1�1���(�փ����į�7�ͽ�����½"�ս�����: !�ƶ/��A7�&&6�,�,�d��&��r��漽Ե��xiz���N��F/����3T�]3��i�E��I��,����1�ޕO��4x����m����;߽z(�w���k-�t�:��A@�&=�42��o!�կ��r����㽱f۽ݪ�7J������j"�m+4���@�/E��A���4���"�W��wD�d5ʽ�%��鎽ov�uZ�X�G��<��c7��H7�x-<�f@F��RV���m�����|㝽}����$޽8���[�?R.���?�ƯJ���M���G�r�:�N)�Ѧ�<2�:�������%�� �nM#��v6���F��nP�#�Q���J��5<�Ӻ(�E)����\ֽ����8[��5򋽗�}��l��a���[�.P[���_��j���z�@㉽�����e���ѽp���vf�]&���9��*I�$RQ�=�P�0H���8��%�=����
r��:j��G����*���<��<K��^R�t�P�nG���6��9"�H��*s�/�̽Y���̙��{���<|��gm�+�d�xta��c���i� Mv�&ꄽ\-��0�k������<��6Z/��B�U=O�}�T��hQ�")F��E5��B"����\] ��+����� ���3��>E��iQ��  �  I#��������;��\t���r���y���H���#�C��	9��lμy0��k�����ü'�ռxL󼪎��-�dV������)��#^Ƚ���y
��J���"�%�k�t���̾⽤�Ž�ӳ�����g���Hս�^�� ��66��'$���%��A��T�'���۽xJ�������Nq���D�B]"��7	�s]�Zټ��ͼ�'ͼ]׼��e������?�^k�e��V���8׽����|����O%���$�������E����ڽ�����봽]~����Ƚ�潷��b���#���*�x�)��M!�_���� ���۽	����8��#}��U��Y7��["�:���*�)�'x����a%��/:���V���|�����.u��݆׽J���`�2�"���.��3���0��&��W��;����ؽYн�׽����~����(�`/4��{8���4� *��%��z����Kƽ����N�r}�w�b��`P��D��7?���>��D�oN�@�^��v�Gˊ�=m������xQٽ�����[��
%���4�uT>�$�@���;��/�]������� �𽊁����	��x�/,���:���C�=KE�p�>��2��� ��}�b���ӽAx������u�����yut�F(i��tc�gc�"h��r�����ƍ�I`��.,����ϽE���
�?�E�/��=�|�D��CD��+<��.���T:�����KE����&���-!��2��?�`�E��zD���;�o"-�.��_��M.��n˽Z\���ꜽ%���4e���u���l�G4i���j�r��~�r���˖�n/��=�����޽Y� �]��x�&��w7�14C���G���D��:��.+�b��:
����>������b��'[���)�"�9���D��  �  ���� ��S�=��!ҽc����/���|�3�S��U2�� ����+���ۼ�׼��߼���D�	�ɨ�X<�H�_�ܡ������
��0IܽU8���j	���P���n���h�� $˽���埢�Ɵ��������2ܽ�@����	���GE�]�x���83ͽ�Ү�j]����w��Q�<�1����AO���q7�)|�Q��v��[��,�.���L�i�r��R���X���}ɽ{��!���n����e��X������A�=�Ľ����6������õ��Ͻ������N��p
����o+�����P�ޙϽu^�����������b��dG���2���#��Y����G���%�105��jJ�r�e�����嘽Uұ���ν?���R�-��U�!��T�H��7j�V�\�ؽy@ƽ����mƽ�Fٽ0���A�	�K ��!�)�%��d#����������V߽�ý����7\��!��	s��K`�.�S��M�y�L��R�1�]�1�n�Q	��M֑��)���d����ԽZz�l	�"�U�$�)y,��9.�)��+��U�����x���޽x�ܽJ������[�َ��d)��X1���2�(.�+�#�%��4����ZOҽ)���J7�������7���	����w��(q�׽p��iv����Ɖ�s���ܤ��Է�/�ν1� �N����!�'�,���2���1��*�Xm����;%����2u�O�b�h�M�j�!��:-�/3��}2�ޟ+����|7���D��g�˽ɵ�.ң� ����{��~�����z���v���x��b��T��?@��YV���殽�UýU�۽�Y�����C��}(���1�S�5���2��)�KB��>�c?��62�J�8�9����'5��	)���2��  �  �w��������-�׽T�½ܬ��A������W�i�qYL���2��/�M�����AR �<��@��W#�[a:�Y�U�Qtt��������@���Uʽ�>߽�(�������S��F߽�ǽ�2��Y��������������ȥ�Y��g(ֽ�\���+���V���c�Uֽ�e��ɪ�w���������h�nL�"�3���� #��>	� ��������<&1��?I�xGe�k���U\��A;��g�����ӽ�S罼%��, ��`u��Dڽ����ᝪ��٘��#��	9���ܞ��ݳ�fVͽ7d潃V����̓������`��\۽��Ž����������6'|�
.b�jL��;���0�O1-�a1��^<�PN���d�9��`������������Ƚ�޽��������
���0B	��������ս:´�谽����8_��������׽}k�{��	����#���L
�Ӂ���]�ؽ� Ľ����q���"��І�]fy�.|j���a���`��@g���t��$��YT��!����}���O���Խ ��� ��
�XF��s�y
�1��9��� �L��>�ս(ʽsvȽԌѽ��㽉����z
��6��'��:� \��_�W�
�D�������ս�cýw#���Ť�&]���:��o↽�䂽�����'������ٖ��򢽥��������ҽ����v��+	��1��������K���j���K���ս,?̽��ͽVٽEn�����L�� ��4H����t�����4���@~�Yѽʿ��c��Uޢ��`��gN���5��|��� І����>Ɠ�����r��.J���˽"�ݽ�u�T9��	T������ �������m�
������q�'�ֽ0�н�ս���)���
��}�����  �  ��ν�xн�1̽��ýP���a:��+%��������?�t��Y���@��,�����*��v"���1�`�G���a���}�:q������/���}��/a��!ɽ!ѽgԽ7�ѽk4Ƚf丽�⥽Lq���7����p�=m��Tz����aɝ�����K(ý��Ͻ2�ս7�Խ-�ν�~Ž91���5���<��������t�@�Y���A�b�/�p%���$�K�-�iy?�T�V��Yq��O������Z��㦬����G#Ľ!�ͽ��Խ�ֽ�ѽo�Ž���-䡽��������v���y����iΗ��5�������~ѽ6�ܽ��a߽�&ؽ�Iν�
ý�S��(Y����
��@��Zcq�Ε\��gN��I�a�M���[�:q�;Ʌ�����g��g.��zN����ɽ�HֽS�ὸ�꽚D������A�۽~[ʽ�;��k/���������CR��Χ�K���ӌν�������m���V���P��]�$w���ؽ�ͽ���D���>��~T���|��%	��p�~�	�|�r,�������L��r��>n�����V5ν�4۽8���
����P������ �c��i߽��̽�d��C���1��(����ɽB&ܽ�`���e��l
��%
�.)�la�q\��B���Խ��ƽڸ�Ld��TZ��� ��
��������9��L���ǲ��������Ľ	ҽ�޽G�[c��gt�)f��	�7b
�������5�ŝ߽X�̽N_���������W��A7ѽز佝'�����P	�/���	�KF�+�����	�꽩t޽��ѽ|NĽ6����ө��Þ�������W��8M���Z���屽ڒ���[ͽ!�ڽ�u�������ɘ�U$
�M���l����I����e޽W�̽[|���黽Lڿ���˽~&ݽq�����	��  �  '𬽱���&q������3������"�������m��&��Zֆ���n���T�U�C���>��5G�7[�*Jw�߃��Κ�_���KT������غ�2������D���.�����IJ����������o��V�1�G�,�D�(O���d��̀�p���ӡ��������ω���o��fs������Uϻ��-��R������뻕����r�m��(V�½H���G�[T���j�]0��
쓽�d������M��c@��ݫ��IX��������	���������ۓ�A�����l���W�!N��XQ��Qa���{��������������ù��6½!^ǽ�ʽ��ʽmUʽ��ǽP�½�	��F,��-ޟ�Zѐ�xT��2�s��k�YZq������6��Oq��5ǯ��/��Sgɽ-ѽp�ս��׽.4ؽ�5׽�3Խ�aν�1Ž�ʸ��/��2��/���z�������w��f>��f|���஽������̽m�׽��޽���r���dr㽒	�ɱٽ~�Ͻ�ý�Q��6�������M��:���x��N$��Wﭽgw���\ν1�۽���Ws�$����J��	���� E�6ܽ�.Ͻkt��A���b�����������ä����y���UϽ�޽#��5��\���t���-����!�����V��x�-�⽍EԽ vĽAY��0b��\����:��=�������r½%9ҽi��"��8��������X��'���Y��o�������.J�/o���ѽ(½R����v���ڢ�٬���Ϊ�#��'Nƽeֽ�^�a���~��g"���_��2�������2��������`��ѽ����~ĳ����J��q���o��h���˽Q۽I/齥���;���p��ñ �+� �mI ��_���N��������u�ѽ�\½�����]���秽�󪽚�������Wѽk�བྷN��  �  �b������s��Mv��"sĽ�ͽ_Nѽ��Ͻ�Xǽ]츽3[����Bʁ��`m�kg�A�q��Å�3뗽)⫽u��7�˽�ҽ�%ӽν|ŽC��~-�������dg��\�u���Z��B�f]/���#�i�!�B�)��;:��Q���k�錃����3��u���a¶�u½��̽��ӽ�\ֽqiҽ��ǽ���W.��쐽1t��Saq�'hp�����掽`䡽�t���#ƽlѽ�ֽTaԽL�ͽs�ý���Z��؟��9��# ���q��+X��*B�Aq2�3e+��D.���:�ގO�ɸi�sB���ؑ�����`d���R����ƽv�ҽ�~ܽ"�����1�ݽ��ѽ����Ğ������xM���
���F������b��Nx���9ҽ⽱�뽮�����S�ٽ�Gνso½}T��ǩ�mǜ�]ď������Ss�Vqf�^�b�E�h��"x��T���̔�\#��@`��3���	̽��ؽ}�����ߺ��	:��������彥�ӽ����>{����y���n���}A���ʽ۸޽u�P���3��/�<��C�����ａp�ʺؽF�̽�@���k��sͦ�9k��p��������f��b����Κ������X��m½Y-нPGݽs������� �&���	�m�
�˔��8��!������GϽW�����.n��\K��� ͽ:$����>�����K
��y	����&�������Bt޽�ѽ�ZĽ���r����������T������k��ᠽ�������|cȽ
�ս"���ｲ*��IK�r���)>�W0����[Q�M�޽�d̽r��������"'ƽ��ֽj��o����� :����`�
����(��ת������E߽/fҽ��Ľ�~��ͪ��3�������!ؘ�G̟��_���4����Ľ�ҽ�  �  ���;������4�ý�ؽ%��u��(_��ګ�{�߽�ɽX���К��������qT������w����Ͻ�����������ܝ��a��(W׽}���AB���엽����pj��}M��b4����P�rx������!� ,���C�`_���~����M����)���&н��佟i�����c���'��-Sݽ�*ŽY߬�B�����"������0U��Q½?�ڽ��������
����z��~ҽ*���{B������� ���d���I��2�7� �g�����+L�+y��X-�̸C�{�^��}�Ǟ�������t��,�ͽ���bu��S��X�����L������̽0t��$��2)�����J$���ǽ���-���+��c`
�Z
�U5�����*{Ͻ�ͺ�0��c��@����x�{c�hS��bI���F��L�&aX�6�j�3B�����y����5�� �ýi�ؽ~��F��D���}I����r��~��Qc޽<zɽ����$�������ѽ���,�����o������d��_j�����Ix⽐�ν뾼�����h7���j��(ى������~���~��	���$�����lW��?���vp��O:н#��rc�����
��ڱ�|���5��������D9뽬�׽O\̽��˽
�ս��GG �<���\�����'�1��R���T������ ҽe��؞�������і�>B�������S��؃����K����7��	���n^Ž{�׽��C� �Y������d���*������I��������ս�,ν�VѽԿ޽'��9d�4�s'�ձ��>�$3�]��@X�$����� ѽ���l����ţ�0����������3���}k���ߏ�v������$ఽ����  �  Y}��𗽄%Խ$��*�E���C�OE��e�� �T$ͽ�벽_��������Ԥ�������Խ����������H�-q�����Fн����^����A{�H_S��-3�w��P��i��9[�8�2���[�@���(�
lF�6k�>	�����FpĽʥ㽵u �	�a�������_�y�彁�ǽc��,���Gġ� ��g�Ľ��̠��&�������~�\������ǽ����D��*_q���L��S/���L
	�fT��:���e���z�����)�1<D���e��<������� ��}۽Gv���J���-|����s ��t����8н�@��$ŷ���Ƚ�3�� �ݐ�yi��~�p��X�
�τ����׽u캽����Ό�	�w��\]��I�"�;��14���2��7�k}A���Q���g��0���ޓ�Fc����½�/�q���|��
��$�Y_'���#�X��DM��,��Y����н �̽0sսU꽀G����k^ ��z)��j,���(��s�*�P����O̽����h��������]�z�/Jo���i��j�_Np�b|�k��6쒽K���e����)˽������e�����+�a!2�g2��2,�Ǡ �q��p*��e�X�པ�߽�4����%&������*�$�1��>2�3N,�1!�+��N������ͽW��8X���d��[ɉ�B��5\w�H$r��s���y�	a��A��C��0��Q뼽��Խ���}��Z%��%�=/���3��2���)�2��=��, �	��C�潓j���('��h%���/�P�4�-#3��Y+�����ė ��&���ʽ�s���$��k��Q�u������|�R��~d��֋�G����*���  �  nz�����Z����彧��ޚ��L ���#��n���~���n&ǽ=!��K���Ŷ��ͽ3���}�����!�ȷ$���˺���7G��� ��v� �G���#�Q�	�\7�Sּ��ɼ��Ǽ�м/�W����Z�8���b�����k7��8�н�������]���$�w�%�x���g�� ���޽�<ýX���������6P۽���}���n�]%%�&4%������������Yս>e���̏�Q�i�]s?�������c��⼏�ۼ��%/����j���4�X�Y�mA��h����ý!��j�6����&���,�N+�^Q"�)����Z��U'νI�ý�ɽa�ܽ���ZB�� �&q,��2��/�u&���wb�y���+��m���ڇ��ui�57M�+y9�&�,�41&��%��")��2���A���W���u�ࠎ�Ƨ���ƽZ�5}��d��|+��G6���9�w�5���*�g��;�	����b`�g0ݽcT罧��}��^�!��l1�{�;��>���9�*=.������
�Dg��ν��������V����{���j��w`��[�&C\�t�a���l���}�l犽	���P���˽�a���zV��m-���;��,D���D�4�=���0�Ҵ������ ������� �����_��׽.�4�<��SD��jD���<��.�/2���	���Bν�(�������~������s�|i��d��Ee��]k�iw�Z���7���#��K㹽tsֽzp��/�O"�Έ3�q>@��DF�ED��H;�,�,�G2���
�h�������b��!�=�Am%�u�5��B��aG�?�D�;���+�2���pi�;�ɽl��������X��僽'�y���q��/o�W�q��y��׃�_,��Y���[ٯ��  �  N{����Ƈǽ��
��{ ���,���0���+��m����o���X�Խ'þ�G^��q�½$�۽I��ѫ�qy#�kx.��e1���+�S7��m�4콎����G���v���B�ԡ�|.��7ݼc	Ƽ� ���Y��Y����YӼ��
��2��\`�ħ������ڽ+�<����'��<1�lI2���*��D�k�	�/3���Ͻeɾ�0׽��Uͽ�S�O���O��m)�I�1�}�1�7))���֏�]�߽Rd��8䑽��g���9����dt �i��\0Ҽ��̼R=Ѽ�3༐W����g}-�ڃT���L����ʽ�������R$���2�t�9�L�7�.��(��~����Jڽ�Ͻ6�Խo��Ԃ�����2+��8�W�>�J<��1����T>�^��Y�ýi����*����b��E�.�0�ޏ$�[M��J��I!��g*�ST9��O�|�n�x���@h��]�ʽ����bP$��]6��|B���F��B��5�l�$����������;�<�8��#r���+�-=��IH�`wK�5�E���8�&����V�����ѽt���%��}����Is��Ab�	=X�C�S��kT�u�Y��~d��8u�����i�������̽+��E���"�C7�n9G�;�P���Q��J��;���(��D�.#�������/���C�˷&�Zp9�Y�H���P���P�LfH�N�8�2�$��>������Sн�>���ݚ�s���(�z�K�j�#a�,�\�Yy]��Cc�֚n�\`��kȍ�B���{���<Pٽ�b������y*���=��L�Z�R�WQ��G� �6�*�#����������q������/��A��TN��T��4Q�$F���4�- ��
���콚�ʽ�Ү�⤙��=��=�=�q���i��qg�k�i�n�q��$�p��-%���ﭽ�  �  �U|�8m����ʽ����o���f$�Z�0�f
5��70�Dr#�Ue�C���Ckٽ7�½�@����ƽ���ً��F�j�'�B�2���5���/�� "�ǂ���𽋢Ľe���F�v���A����E��)�׼J�����cK���k��μ�{����1��`�ӌ��������޽h����`�+���5��6��/�& ������zԽ5�½������ѽD����
�1�ѯ-�lT6��96�2P-��&�
b�S��͸��풽�g��E8�"�������ݼ�ͼ~�ǼF>̼ۼ/ ���~��X+��KS�v!��来�Ԝͽt��ƙ�y�'�-�6�a>�vd<��B2��!�ޔ� ����޽�ҽ��ؽ�|�LU��J��(/�<=�	DC��m@��5��D#�������Ž14���څ���`���B��J.���!�������~����'��6�%M�y�l��W��_��}̽���r���'��I:���F��(K�X�F���9�1"(������7��j������s�?�/��A��L��O�C5J��|<��-)��8�/����Eӽ�W��X���^�����p�;�_�&�U�qCQ���Q��IW���a�
�r�����^;��:�����ͽ[����br%��:��QK��U�A'V��^N�y]?�'A,�����`	��} �9���������>�)��:=��L��U�jnU���L�Kj<���'�/=��U��p[ѽ�5��(��5k���.x��h�"p^�q4Z�#�Z�9�`�P�k��.~�����ꟽ������ڽ0�~��x-�O�A��UP��kW���U��3K��:� '������2� �v�R����y2��	E��R�{�X��U�pJ�-.8��"��C�����1˽����������|��n�f\g���d��hg�o�ǀ|��Ȉ�:.��~����  �  N{����Ƈǽ��
��{ ���,���0���+��m����o���X�Խ'þ�G^��q�½$�۽I��ѫ�qy#�kx.��e1���+�S7��m�4콎����G���v���B�ԡ�|.��7ݼc	Ƽ� ���Y��Y����YӼ��
��2��\`�ħ������ڽ+�<����'��<1�lI2���*��D�k�	�/3���Ͻeɾ�0׽��Uͽ�S�O���O��m)�I�1�}�1�7))���֏�]�߽Rd��8䑽��g���9����ct �d��V0Ҽ��̼H=Ѽ}3༂W����]}-�σT���
L����ʽ�������N$���2�q�9�I�7�.��(��~����Jڽ�Ͻ7�Խq��Ղ�����2+�
�8�[�>�N<��1����X>�e��`�ýp����*����b��E�4�0��$�]M��J��I!��g*�NT9���O�s�n�r���:h��V�ʽ����^P$��]6��|B���F��B��5�j�$����������;�<�9��%r��+�0=��IH�cwK�8�E���8�&����]����ѽ{���%�������Is��Ab�=X�H�S��kT�x�Y��~d��8u�����i�������̽+��E���"�C7�n9G�;�P���Q��J��;���(��D�.#�������/���C�˷&�Zp9�Y�H���P���P�LfH�N�8�2�$��>������Sн�>���ݚ�s���(�z�K�j�#a�,�\�Yy]��Cc�֚n�\`��kȍ�B���{���<Pٽ�b������y*���=��L�Z�R�WQ��G� �6�*�#����������q������/��A��TN��T��4Q�$F���4�- ��
���콚�ʽ�Ү�⤙��=��=�=�q���i��qg�k�i�n�q��$�p��-%���ﭽ�  �  nz�����Z����彧��ޚ��L ���#��n���~���n&ǽ=!��K���Ŷ��ͽ3���}�����!�ȷ$���˺���7G��� ��v� �G���#�Q�	�\7�Sּ��ɼ��Ǽ�м/�W����Z�8���b�����k7��8�н�������]���$�w�%�x���g�� ���޽�<ýX���������6P۽���}���n�]%%�&4%������������Yս>e���̏�Q�i�\s?�������[��⼁�ۼϜ�/����j���4�C�Y�aA��h��{�ý��j�/��y�&���,�N+�XQ"�%��
��U��S'νH�ý�ɽe�ܽ���^B�� �+q,��2���/�|&�&��b����	,��y���*ڇ��ui�E7M�7y9�.�,�91&��%��")��2���A���W���u�ՠ���ŧ���ƽ�Y�.}��d��|+��G6���9�q�5���*�c��8�	����``�g0ݽeT罫�����b�!��l1���;��>���9�1=.������
�Sg��ν��������V����{���j��w`���[�.C\�z�a���l��}�m犽
���P���˽�a���zV��m-���;��,D���D�4�=���0�Ҵ������ ������� �����_��׽.�4�<��SD��jD���<��.�/2���	���Bν�(�������~������s�|i��d��Ee��]k�iw�Z���7���#��K㹽tsֽzp��/�O"�Έ3�q>@��DF�ED��H;�,�,�G2���
�h�������b��!�=�Am%�u�5��B��aG�?�D�;���+�2���pi�;�ɽl��������X��僽'�y���q��/o�W�q��y��׃�_,��Y���[ٯ��  �  Y}��𗽄%Խ$��*�E���C�OE��e�� �T$ͽ�벽_��������Ԥ�������Խ����������H�-q�����Fн����^����A{�H_S��-3�w��P��i��9[�8�2���[�@���(�
lF�6k�>	�����FpĽʥ㽵u �	�a�������_�y�彁�ǽc��,���Gġ� ��g�Ľ��̠��'�������~�]������ǽ����D��*_q���L��S/�}�F
	�VT��%���K���z�����)�<D�|�e��<������� ��h۽2v��{J����$|����l ��t����1н���@��&ŷ���Ƚ�3�� ����i��~�y��X�
������׽�캽����"Ό�$�w��\]�'�I�.�;��14���2��7�b}A���Q���g��0���ޓ�5c����½�/�\���r��
��$�P_'���#�Q��>M��,��S����н �̽3sս[꽄G����r^ ��z)��j,���(��s�*�[����O̽(����h��-������q�z�@Jo���i��j�hNp�!b|�n��7쒽K���f����)˽������e�����+�a!2�g2��2,�Ǡ �q��p*��e�X�པ�߽�4����%&������*�$�1��>2�3N,�1!�+��N������ͽW��8X���d��[ɉ�B��5\w�H$r��s���y�	a��A��C��0��Q뼽��Խ���}��Z%��%�=/���3��2���)�2��=��, �	��C�潓j���('��h%���/�P�4�-#3��Y+�����ė ��&���ʽ�s���$��k��Q�u������|�R��~d��֋�G����*���  �  ���;������4�ý�ؽ%��u��(_��ګ�{�߽�ɽX���К��������qT������w����Ͻ�����������ܝ��a��(W׽}���AB���엽����pj��}M��b4����P�rx������!� ,���C�`_���~����M����)���&н��佟i�����c���'��-Sݽ�*ŽY߬�B�����"������0U��Q½?�ڽ������������z��~ҽ*���|B������� ���d���I���2�/� �]��z��L�y��X-���C�Z�^��}����������t���ͽ���Ju��G��M����:������̽(t�� ��1)�����P$���ǽƇ�=���4��n`
�f
�a5�4���'�C{Ͻ�ͺ�F��(c��Q����x��c�wS��bI���F��L�aX�#�j�'B�����f����5���ýP�ؽd��F��D���rI�����r��~��Fc޽5zɽ����#�������ѽŲ�,�����o�ɐ���q��lj����bx⽨�ν�������y7���j��5ى������~���~��	���$�����mW��@���vp��O:н#��rc�����	��ڱ�|���5��������D9뽬�׽O\̽��˽
�ս��GG �<���\�����'�1��R���T������ ҽe��؞�������і�>B�������S��؃����K����7��	���n^Ž{�׽��C� �Y������d���*������I��������ս�,ν�VѽԿ޽'��9d�4�s'�ձ��>�$3�]��@X�$����� ѽ���l����ţ�0����������3���}k���ߏ�v������$ఽ����  �  �b������s��Mv��"sĽ�ͽ_Nѽ��Ͻ�Xǽ]츽3[����Bʁ��`m�kg�A�q��Å�3뗽)⫽u��7�˽�ҽ�%ӽν|ŽC��~-�������dg��\�u���Z��B�f]/���#�i�!�B�)��;:��Q���k�錃����3��u���a¶�u½��̽��ӽ�\ֽqiҽ��ǽ���W.��쐽1t��Saq�'hp�����掽`䡽�t���#ƽlѽ�ֽTaԽM�ͽs�ý���Z��؟��9��" ���q��+X��*B�6q2�$e+��D.�u�:�ÎO���i�_B���ؑ�����Fd���R����ƽY�ҽ�~ܽ�⽨���ݽs�ѽ������������tM���
���F������m��\x���9ҽ����������o�ٽ�Gν�o½�T��ǩ��ǜ�mď������Ss�`qf�`�b�?�h��"x��T���̔�J#��+`�����	̽��ؽ`�����ú���9����������彖�ӽ����6{�� ��y���r����A���ʽ�޽��f���?��<�J��`�����｝p��ؽ_�̽�@���k���ͦ�Hk��|��������f��h����Κ������X��m½Y-нPGݽs������� �&���	�m�
�˔��8��!������GϽW�����.n��\K��� ͽ:$����>�����K
��y	����&�������Bt޽�ѽ�ZĽ���r����������T������k��ᠽ�������|cȽ
�ս"���ｲ*��IK�r���)>�W0����[Q�M�޽�d̽r��������"'ƽ��ֽj��o����� :����`�
����(��ת������E߽/fҽ��Ľ�~��ͪ��3�������!ؘ�G̟��_���4����Ľ�ҽ�  �  '𬽱���&q������3������"�������m��&��Zֆ���n���T�U�C���>��5G�7[�*Jw�߃��Κ�_���KT������غ�2������D���.�����IJ����������o��V�1�G�,�D�(O���d��̀�p���ӡ��������ω���o��fs������Uϻ��-��R������뻕����r�m��(V�½H���G�[T���j�]0��
쓽�d������M��c@��ޫ��JX��������	���������ۓ�>�����l���W�� N��XQ��Qa�~�{��������������ù��6½^ǽ�ʽ��ʽPUʽ��ǽ7�½�	��3,��ޟ�Nѐ�oT��(�s��k�_Zq������6��]q��Gǯ��/��lgɽGѽ��ս�׽L4ؽ�5׽�3Խbν�1Ž�ʸ��/��,2��/���z�������w��_>��[|���஽������̽U�׽�޽ߙ��q����Gr�w	཰�ٽh�Ͻ�ý�Q��*�������M��:���x��V$��cﭽvw���\νG�۽���rs�6$���h��&����E�#6ܽ�.Ͻ}t��P���b����������ä����|���UϽ�޽#��5��\���t���-����!�����V��x�-�⽍EԽ vĽAY��0b��\����:��=�������r½%9ҽi��"��8��������X��'���Y��o�������.J�/o���ѽ(½R����v���ڢ�٬���Ϊ�#��'Nƽeֽ�^�a���~��g"���_��2�������2��������`��ѽ����~ĳ����J��q���o��h���˽Q۽I/齥���;���p��ñ �+� �mI ��_���N��������u�ѽ�\½�����]���秽�󪽚�������Wѽk�བྷN��  �  ��ν�xн�1̽��ýP���a:��+%��������?�t��Y���@��,�����*��v"���1�`�G���a���}�:q������/���}��/a��!ɽ!ѽgԽ7�ѽk4Ƚf丽�⥽Lq���7����p�=m��Tz����aɝ�����K(ý��Ͻ2�ս7�Խ-�ν�~Ž91���5���<��������t�@�Y���A�b�/�p%���$�K�-�iy?�T�V��Yq��O������Z��㦬����G#Ľ"�ͽ��Խ�ֽ�ѽn�Ž���*䡽���������v���y����[Η��5�����o~ѽ�ܽ��F߽�&ؽ�Iν�
ý�S��Y����
��0��Bcq���\��gN��I�f�M��[�Nq�IɅ�����g��.���N���ɽ�Hֽp����꽵D�	����U�۽�[ʽ�;��t/��
�������@R��Χ�@���Ōν�������m���V���P��@�w���ؽmͽ�����C���>��oT��|��	��h�~�	�|�v,�������L�����Pn������n5ν�4۽T����4��^��)���� �x��i߽�̽�d��C���1��.����ɽE&ܽ�`���e��l
��%
�.)�la�q\��B���Խ��ƽڸ�Ld��TZ��� ��
��������9��L���ǲ��������Ľ	ҽ�޽G�[c��gt�)f��	�7b
�������5�ŝ߽X�̽N_���������W��A7ѽز佝'�����P	�/���	�KF�+�����	�꽩t޽��ѽ|NĽ6����ө��Þ�������W��8M���Z���屽ڒ���[ͽ!�ڽ�u�������ɘ�U$
�M���l����I����e޽W�̽[|���黽Lڿ���˽~&ݽq�����	��  �  �w��������-�׽T�½ܬ��A������W�i�qYL���2��/�M�����AR �<��@��W#�[a:�Y�U�Qtt��������@���Uʽ�>߽�(�������S��F߽�ǽ�2��Y��������������ȥ�Y��g(ֽ�\���+���V���c�Uֽ�e��ɪ�w���������h�nL�"�3���� #��>	� ��������<&1��?I�xGe�k���U\��A;��g�����ӽ�S罼%��, ��_u��Cڽ����ޝ���٘��#�� 9���ܞ��ݳ�WVͽ&d�oV�������j���~`��\۽��Ž����������'|��-b��iL�ӝ;���0�M1-�f1��^<�bN���d�X��#`������آ��ʛȽ!�޽��������
���:B	��������սB´�谽����5_��������׽pk�{��	�������L
�Ɓ���D�ؽ� Ľ����q���"��І�Ify�!|j���a���`��@g���t��$��fT��1����}���O���Խ��� ��
�eF��s��
�;��B��� �Y��I�ս1ʽzvȽٌѽ��㽌����z
��6��'��:� \��_�W�
�D�������ս�cýw#���Ť�&]���:��o↽�䂽�����'������ٖ��򢽥��������ҽ����v��+	��1��������K���j���K���ս,?̽��ͽVٽEn�����L�� ��4H����t�����4���@~�Yѽʿ��c��Uޢ��`��gN���5��|��� І����>Ɠ�����r��.J���˽"�ݽ�u�T9��	T������ �������m�
������q�'�ֽ0�н�ս���)���
��}�����  �  ���� ��S�=��!ҽc����/���|�3�S��U2�� ����+���ۼ�׼��߼���D�	�ɨ�X<�H�_�ܡ������
��0IܽU8���j	���P���n���h�� $˽���埢�Ɵ��������2ܽ�@����	���GE�]�x���83ͽ�Ү�j]����w��Q�<�1����AO���q7�)|�Q��v��\��,�.���L�i�r��R���X���}ɽ{��!���n����e��X������A�:�Ľ����6������õ��Ͻ������E��g
����e+�����P�əϽb^��
���������b�wdG��2���#��Y���H���%�?05��jJ���e�����嘽hұ���νS���R�7��(U�!��T�O��=j�V�c�ؽ|@ƽ����mƽ�Fٽ(���;�	�D ��!� �%��d#����������V߽�ý햪�(\��	!���s��K`�#�S��M�x�L��R�<�]�A�n�\	��Z֑��)���d����Խnz�v	�*"�_�$�3y,��9.�
)��+��U����y���޽}�ܽO������[�ڎ��d)��X1���2�(.�+�#�%��4����ZOҽ)���J7�������7���	����w��(q�׽p��iv����Ɖ�s���ܤ��Է�/�ν1� �N����!�'�,���2���1��*�Xm����;%����2u�O�b�h�M�j�!��:-�/3��}2�ޟ+����|7���D��g�˽ɵ�.ң� ����{��~�����z���v���x��b��T��?@��YV���殽�UýU�۽�Y�����C��}(���1�S�5���2��)�KB��>�c?��62�J�8�9����'5��	)���2��  �  I#��������;��\t���r���y���H���#�C��	9��lμy0��k�����ü'�ռxL󼪎��-�dV������)��#^Ƚ���y
��J���"�%�k�t���̾⽤�Ž�ӳ�����g���Hս�^�� ��66��'$���%��A��T�'���۽xJ�������Nq���D�B]"��7	�s]�Zټ��ͼ�'ͼ]׼��e������?�^k�e��V���8׽����|����O%���$�������D����ڽ�����봽X~����Ƚ�潳��]�z�#���*�q�)��M!�W���� ���۽�����8��}��U��Y7��["�1���*�)�)x����a%� 0:���V���|�����;u���׽Y���g�:�"���.��3���0��&��W��;����ؽYн �׽����{���(�[/4��{8���4��*�~%��z�x��Kƽ겨�C�r}�h�b��`P��D��7?���>��D�wN�K�^��v�Pˊ�Gm�������Qٽ�����[��
%���4�|T>�+�@���;��/�a������� �!𽏁����	��x�/,���:���C�=KE�p�>��2��� ��}�b���ӽAx������u�����yut�F(i��tc�gc�"h��r�����ƍ�I`��.,����ϽE���
�?�E�/��=�|�D��CD��+<��.���T:�����KE����&���-!��2��?�`�E��zD���;�o"-�.��_��M.��n˽Z\���ꜽ%���4e���u���l�G4i���j�r��~�r���˖�n/��=�����޽Y� �]��x�&��w7�14C���G���D��:��.+�b��:
����>������b��'[���)�"�9���D��  �  ��/���+�e��Q�Zu�u�Ž�]���z���D�"��/����(׼	��$x���,��ڳ�(�ļ�0⼝e��^'���R�兽����|�ѽ�����H�Rp$��9/���1�(�+��2�)�����ҽ�D�����E�Ƚ��㽀��-��E'��0��62��+����\	�������Yf��Up�RU?���e� ��s޼ �ȼ�6������|�ƼP(ۼ�\��j��U:���i��Y��JE���⽚��7p�H�)���1�1���(�փ����ï�5�ͽ�����½�ս�����7 !�ö/��A7�"&6�(�,�d��&��r��漽ε��miz���N��F/����/T�[3��i�F��L��1����1��O��4x����s����;߽}(�{���k-�w�:��A@�&=�72��o!�֯��r����㽲f۽ܪ�5J������j"�k+4���@�/E��A���4���"�S��pD�]5ʽ�%��鎽�nv�
uZ�R�G��<��c7��H7�y-<�i@F��RV��m�����㝽�����$޽<���[�CR.���?�ɯJ���M���G�u�:�P)�Ӧ�>2�=�������%�� �oM#��v6���F��nP�#�Q���J��5<�Ӻ(�E)����\ֽ����8[��5򋽗�}��l��a���[�.P[���_��j���z�@㉽�����e���ѽp���vf�]&���9��*I�$RQ�=�P�0H���8��%�=����
r��:j��G����*���<��<K��^R�t�P�nG���6��9"�H��*s�/�̽Y���̙��{���<|��gm�+�d�xta��c���i� Mv�&ꄽ\-��0�k������<��6Z/��B�U=O�}�T��hQ�")F��E5��B"����\] ��+����� ���3��>E��iQ��  �  < ���$���V��=q���L��(�I����ս橽���c��C�%�.���#��� �&�ʏ3�o�J�azn���g���8����D1�KXV�}Oz����j����͗�d�������m���L��1�c� �qy���(��@��2_����*�������嗾*���B΄���g���B�q��}��Ɖʽ�Y��˲���y_��\C�2�Ț)��)���0�ߡ@�FD[�3���t.���ŽM������OI>��ac�l肾�@��/l��k��DP���ށ�Ec���C���+�~�,�!�ޜ1�(�L�|�m��%��D哾g���H���Đ��z����a��<��>��)��3�ɽ䶥�*֋��Dt�d�]��wQ�r�M�)�Q��^��[s�P��J���|½r�YE��=3���W���|�����3@������<��Zh��������f��JI�8�4�"-���3��H��e���������T���"���Kݝ�+ ��c��^_b�z�=����� ��Xֽ����������.<�����!���a��eꋽ�O��[ت�u+Ž$�0�q�)��#L�Vq� ���ę�KZ�����҆���唾�i��i�j�o�O�N@?�|r<��G���_���~����P������������[Ԕ��ヾ�b���>�V�������z�ý����qz����My��'2���薽����OV���p��3ݽ��V�o:���]�"����͒��)���U�������.������y_���%c�L�J��&>���?��iO�<�i��;���?��̼��J��|���
	������{�{���V��#4��T�����/fؽ���ݞ������ᴘ������5���}���[��*��̽������@'�H�l�l�ʾ��*������Q��Ng��My�����@iz�c�\���G���?�WSF��Z��Cw�/��ac������  �  t"��xm�������k���H��b%��g��ս"�������Pg�I2G���2���'�\%��0*���7��N��Ir��[��wӴ���)F��S.���Q��t�~����͑�*�k����;���h��aH���-�~v�eb��3%�]�;��Z�b�y�释�/Ғ�����̭����b��-?����r��Vʽd��o���c�݌G��26�;�-��"-�"�4���D�"\_�xt��IS��K Ž0��������:���^�ֱ�ݰ��m���Q=��^����v}�=^�0�?�@(��f�j���-��<H�>h�烾z?��񌖾b}���L����1]�ǰ9��v�����T�ɽ��������ix���a��U�-�Q��U�K*b���w�����D(����½��콯�5�0���S��{w��j��N����5��w��n����ƀ�	�a��PE��l1�*���0�+D�T�`�k����z����ĝ��&��yя�$����V^��2;��P�� ��	׽���x���休�gN��w��������h�������`��������ƽ������(��1I��l��܇��X��8����ࡾU֜�V�������4f���K�<�]X9��{D�g[���y�V쌾z����ڢ�������������f���_�̅<����}���vrŽ���*���6ҙ��}���5����������a���9½�/޽���to��_8���Z��N~�񽏾���������"��ƚ������}}��^�%;G�k;�V�<��K���e��|���������\(���碾ɐ��X����Vw��S�,[2�0�����ҹٽ�ֿ�����3����������L<������Us����6tνb��k����%���E���h��������ݠ�t��á�����F����u�d�X��nD��<�7C��*V�wr��C�������P���  �  NU��/����w���\���=����b3Խ�����!��c(t�ĽT���?��a4�Q\1�#�6���D���\��%�%{���<����P@	���&��CF���d�}~�;N��/$�� \��$�s��5X��o;��G#�Xa�U��o�	0���K�*�h�P����"��UR��'��'r�GMU�q�5���f����˽e���n��+�p��U�RC�C:�E�9�A��;R�1�l�H�������%ƽo������1��Q�V�n�|҂�{鈾̄��}���5�k�]9O�#�3��W�����x�L�#�x�;���X�A�u���7Ƌ�튾����
o��Q�֌1���;����˽�����G����Go�+Hb�G^�WYb�
1o�)���򚒽g֨��bƽ׉�5�jQ*�ĕI�=i�Yt���V��Mk��㍾4C����p�!T��
:�-�'�^Q!��h'�4)9�JES���p�텾�r�������ԏ�~����r�K�S�k[4����$ �1ڽ�
������q���َ�։��$��R���"���} ���#����˽����
�)�#��{A�T@a�a
��X匾���"��z{���I���`u��Y��eA�N�2�Z�0�֮:��O�WFk�8��(����)���\������/��!Iu���U���6�����(�	��}p˽o^���K��EF��<����h���b���ŧ���?YȽ���>������.3��Q�"<q�&T��Ṓ�ј�mh��f�������!�n�5�R��H=�C22��3�`mA���X��u�ڈ��ԓ�%_���U�����������(k��K���-��[�����޽�-ƽ@v���c�����k+���|��X��P6��i����%Խ�$�:m��#�H1?�la^��}�oˌ�E����������9U��fW����g��]M�.�:�"�3���9��$K���d��
���l��6ϗ��  �  �xq�_�l�.^�D�H�p}/�:O�l�����ֽ�2���ț��䆽{n���W�(�J�1G�3HM�!]�
v��E�����	���1!ήF����6��MO�2�c�a�p�ps���j�*�X��@�$=(�q������[�V��у�U6��N� #d��;q���s�pk��Z���B��y)�����P����Ͻ8J��,����Y��k�m��8Z��O�gPO��mX���j�oI������~歽�˽>H����rR&���?�DhW���i��s�e�q�Rf�y�Q��^9�]�!���^_����P���(�1B���Z��#n��Vx���w�P>l���X�T�@��['�����l��%�ҽӶ�˲���Ϗ�uɃ���x�	�s�_x��R�����n��殴�VJϽ��ｚ����"�-�;�G^U���k��|{��ڀ�  }�#n�0X�0y?�@)�J���,�1v���(�9?���X�b�o��*���c����3�s�n0^�9>E�9",��*��~�_��?�Ƚ�\��� ��j����㔽��◽�����ԭ��ɿ�*�ֽO�|���@�7���Q�elj��R��o��kb���Ju�V	^���E�v�1�t<%��:#��,���=��U���n���������鉾h����z���b��aI�r�0��d���	o��׽<Ľ#���oӫ�,���GK���ت�<������ֺԽ9���Y�l���s-���E�{�_��,w�"����s���׈�����cq���X�u�@�g.�B�$��+&���1�pF��^���v�=߄�N���m,���`���s��Z�%]A�dg)��q�����w齩�ҽ�C������g�����􁪽rӰ�sǻ��j˽��^��s)�	� �(�7�2�P�Cj��4�����/��֬���$��sl�5S��<���,��&��+���:���P��i�nj��̃���  �  �ZN�`L��cB�&�3�W"�jd������7�ǽ�P���国S֊�E�{�z�k�"bg��o�3����2��qY��7�����ν�O�[���[�'�˹8�w�F�4O�ۺO�H��#9���%����� ���콸�������	�����O1�|�B�`�M�*Q�1L�`y@��m0�G���%��*��<�ݽ�Ľ.���<��*��
;}��p�y�o��{�#���ꗽ�������[ڽCL��L�
��V�\+.��>���J���P���N��eD���3���������.�����b�� u'���;���K�`	U���U�T�N�YsA��0�	��'���\���ʽEе��.��Yu���y���������)��p����T���Wɽ�5���������op/�24A���P��D[���^���Y��lM�Xe;��^'�tY����f�b��DI���'��n<�*�O�Xv]��c���a�� X��:I���7�w9&����l
�����8ݽ�[ɽ��²���|���������v򲽰���7�Խ=�������W:�mg0�f{B���S��b�Q�j�&�k��8d�A�U�-�B��'/����P���I�~�.)�â<�,!Q���b�`�m�7q��=l�t~`��dP�ɉ>���,�^���h�������ؽ��ȽGS�����������-��E$ǽG�ֽ˼齦���1��<����*�
�;��M��J^�Z�j�p�p��\n��d�(<S�2 ?�%�+� ��}�����ɕ�Q�/�JD���W��xg��)p�A�p��)i���[���J�C9�(�'������
�N�����Y�ս�+ǽ�l��7���	����½�kϽZ�m���>�U%���!��w2�mAD���U�pae���o�v<s�Ln���a��OO�� ;��(�����	����5'�E<9�īM���`�� n��  �  ��,���-���)���"�[��#l�����#��P���Iн�ͺ��}Җ����۫��~����������*���n�ֽ���J ��#
����-f��.&�=�,�C�/�^�-�~;&����LE
�����i�ڽإʽ��ǽ�\ҽ���v������!���+�5k0�ע/��w*�n�"��C�_������l0㽉~ͽ�/���,��-���M������S��	'��������ʽ~t�l�����dV���c6!�f)�� /�9j0��,��7#����T��N���ֽ��˽>ν�޽����r��]��|U*�3�o26��4�	.�o�%�Do�����u	��(��Kw�_cս\��Oo��`Ĥ�Q���1���­�R]����ҽ�G�����Ht
�V���p�#+(��d1��
9�
�=�]g=���7��-�������� �,s��j��,����� �_�/�q;��-B�%TC���?��8���/�VC&������	��1���A�=ս�Žv����������~u̽
�޽����D�L����r�$��.��Y8�gGA��*H�SeK�=�I��^B�M6�bB'�%���B����H���>�^���#�{R3�%�A�X�K�<rP�˪O��xJ�uB�p&9��}/��%�C���'�n=�u��a��W\ս�9ͽ&�̽��ӽ;���b�����O��I,��3$���-�^�7���@�N I���N��$P��3L�}�B�L5�%����C3
��;�P�Á�lH��)�	�8���E�5&N��P���N�6MH��?��h6�P�,��&#���`��q�����o�òԽO:Ͻ��ѽ%Q۽z&�
���X
��9�*����)��Y3�c�<�q)F�U�M�J.R���Q�+L�G-A��p2� q"�z"��3
��w���	��Q'!��B1�Pl@��L��  �  ,�g��������������D��*��-	�����L�܁˽|������W�����GK��j�ѽ�뽬�����d5�����|�x]�/��+{����Y������hʽo��,P�����\0���<���bؽH��|��и������q��X��dE���ND�O+��)��p��/%�RȽ9��)]��~����T���zŽ�!ݽ^l��a�����~��/����-R����L���#�Ơ��G�,i��G�ܽ�Ž8���xG��e_���sϽue�v]�S6����'��B� �[I"���"�eK"��_ �M��w�����& �����ѽ�½����6X����̽�S⽠����
�i6���Ƞ$�V�'��7)��|)���(��s&���!�s���}�������t۽&ͽ�GȽ��ͽ��ܽ!+󽞃��D��6��e&�4�+�#y.�|�/���/�'�.�[4,�<:'��h�����������O�ivؽSսE�ܽ��u�~+�����I&�m .�~�2��a5��j6�&q6��Z5�\�2�<-�%�n�lZ���������a��*�@�����Q����$�:�.�M�5�4�9���;�r�<��$<�I�:�z�6���0���'�5�΀�i������`轻����T����i;&���/�� 6�F�9�˂;��;��};���9�K�5��C/�V�%�/��q��������	꽞N��7b�7���?�c�(�J�1�M�7�e�:��<�	�<��><��0:�-�5�b�.��%��b���-�`����U������L��� �ř �;�+�d4���9���<�->�#D>��q=�L;��q6�	�.�Ы$��~����0���L{�>�)M ������U $�m�.��  �  U6����ͻ��X�X#��*�pD.�� -�qq&�`��-��OA��3�۽6�ɽ��Ľ�ͽ���L������h��G)�y�.���.�yw*���"�T��qK�F�������(�Ͻ���ү��.d��}@�������������vα�W�ƽ��ܽ5��J�������� �t�(��.���0���-��N%�]��T��x��}ؽbWʽ��ɽ�<ֽ�&�]o�yR�|�#�`�,��0�,�.�Y)�� ��`������O��"x߽Lʽ!��������喽�㐽4����/�����W��_�ֽ{r��� ��������s<)��P1�݃6�F7�)�2�̧(����q�
�����?��۽	�߽ ��)��N����&�yp3�v;�=-=��/:���3�M�*���!�B�xi��l����;�޽v8˽����\���묽�N������^ν\㽤���L��������f&��0��#9�^a@�g5D�V1C�ܭ<�c&1�jF"�ӧ��=��1��ŷ��������	�U��49)��E8�7mC�]BI��I��7E�I�=���4�,�+�#"�������/�%��F�c�ҽ)�ʽV�ɽ��нV,޽@��`�O$���}#�^�,�?�6�D�?��^H��vN�&�P��yM���D���7���'���I���}�2�l
��b�a�%���5�dGC�RlL��P��tN���H�rg@��7��u-���#����A8��`����i�m�ӽ�,ͽ�#νɲֽa������3���I��\�&��Y0��:��KC��<K��KP���P��L�5�A�n�3��#�M��f�	�����Y��>��-��<��H��[P��>R�7!O�weH���?�w>6�I�,�o�"�����-��d�Y��%�ὦEֽ�ҽ��ս���oK�S���������  �  �⽜W ��"��#��4�PC���L���N��rH���:���'��x����Uz�е�g�����U�
�,���>�XoK��P��hL���A��82�^� ����a���@�7lƽ臯�-���$#��0�}��o�%&m�%�v�g���c����/��E ���ս���e�a��h�+��b<���I�v�P��O���F���6�@#�R0�<S���j뽘s����ʲ �6�4�<E�� O��P�d�J�3�=�`F-�rc�3
�4���$�ؽ\���y�����f����~�M�u��*y�./�����RA��7����νZ�;X�D����%�4�7�#�G��hS�7X��T�׋I�_=8�-H$�w��9��P�����W�����2�&QF�sKU���\��#\�w�S�
�E���4���"�����I뽕Խ������� ���o������	�����(��(eĽ��ٽ�-�گ�g��j�&���8�UJ�Y-Y�m�b���d�h�^��Q��s>�p~*��/������
����j��v1��@F�y�X�L�e��aj�*�f��h\��M��;�!2*���+��!s��IM�|1սΗŽ?�����������
��t�ý�Yӽ�r潕���^�
�����[(���9��tK�,:\�'ei��jp�i�o��ef�egV�B���.���<^�L��x�Nd,��@��T���d��n��Rp��j��l]�M�L��
;�b�)�����������l�Hֽ��ƽM��"��Jַ�i���lʽ*�ڽx�b���~����]8.��?���Q�.�a�'m���q��<n���b�� Q�p�<��)��ڹ��D�W-#��n4��H�\��j��+r�:q���h�5}Z��PI���7�ǵ&�y���$
��w��݋���սt/ȽgR��8��������ǽս����x����	��  �  !�׽t �s��0���I�Y_���m���q�)Ck��Z��C�h�*�@$�������a	���l�0�(�I���_�t�n��r��cl�b\�i�E�B�,�1��/S����ӽ�<��Ě�Q����.o�fJZ�ūN�ĲL��T��e�"������O���Lƽ��r.
��^"���;�("T��g���r�!Ds�f i���U�|=�%��b�*�C�����P�"�?�:��S�/g��yr�Bs�O�h��\V�.�>���$�J���-�< ʽ�լ�ω�������(m�á\���U���X��{e���{������1�������۽s>������0���J�}�a�1�r�>�z��x�f�j���U�Y.=�p:&�Hi�� ��y��?�w�4��N�b f��w����j\}��]p���[�K+C���)�mr��[����ڽۿ�ϙ������f<��梈��ӆ��ё��H��Ai��Q|Ž��ud�.���$-� �F�*�_�8u��ȁ�N��D���f3q��fZ�9�A�z,�������!�ex2���I�}"c��y�,I������-p���w�
�`���G�9�.�{��ؗ��2��tӽ4���M[��rd���3���ԧ����z׾�Lѽ������ *��LB��[���s����*��o��]D��U>u���\��tD�\�0��z%�#�$���.���A���Y�wr�>�����D���A����u�: ^�1�D�0<,�������̟�B�ӽ����]������Kͦ�^p��;�)����Ž��ٽ������f42��K��d���{�FS��?���������V�n�o�U�%x>�:R-�_�%�ʯ(�6��HK�,d���{�����	����;��R�����p���W��>�p'�@������>轹zҽ����Wֵ������VC���_������ѽ`	�{	��  �  !�ս�9��  �sw?�#�^�rPy�`�����������T�v�$�[�/�>��f%���������*�2pE�Q�b�bh|�r���g������Ju��YY���9�T��{���н����ˎ�Ųs�
 V���B�?�8��7���=�]M�"�f�����#����ÿ��%�-�&�,�ϜL�9�j��u�������>��e��]hp��T���7�K� �`���������4�˺P�]Vm�vO���ӈ�kۈ��l���m���O�q50�4�9l�DĽ�����*����m���T�4F��*@��C�{�N�?�b�Ì�3������lo׽�������=��X]��)z�Ї�����^�������9o��kR�ߚ7�5�#�C4��,��(/�8/H�f�e�򵀾���8���h���Gi��Pq��yR��3��"������(ӽ󒴽�ݝ�gȍ��A����z��x�ٳ}�0���U�������{�����ؽ�A �=���5�o<U�lt�r���+��� �����o����cr�v�U�m�<�_,���'�!�/�MfC��s^�]�{�C
�����&��쑾`����'t���T�,6�˞�C�����7mǽ�E��T��𒜽�N��D���h��Ѥ���Ľ�޽�q������.���L��|l��C���T���`���
���(����~s�iW�g@�N�2��,2���=�I�S��p��V��<���z���K����-��/����~o���O�T�1�8H����G὿�ǽ���j���-���Lq~���S��C������nͽG�ʚ�l�n�8���W�yQw�����ᥔ�鹙�"8���i��o�
�j���O���;�[�2�e6��F�0�^��{�'����ٕ��W���4��'現� ���Kg���G��*���������ܽ��Ž����٩�uS������&��j|��p���Ľ��۽�����  �  ��ֽ����'�9�J�4�m�yޅ�����b���X��QǄ�,�k�yL�EN0�V��I���-!�}!6��wS���s������M��%ɓ�ߎ�G���r�g�RD��9!����нmm��[���df���H���5��3,�$�*�81�W@��Y��~�fؙ����5	�P��jD5�9Y���z�(!��>%��5�������F��Rec�8%D���*�E��g��d�(���@��_�S0�j��7���M���{<���4~���\��9�������½���#���@`�J�G�OS9�t�3�?�6�M�A���U��St��>��٥���
׽]D�U$��AG�k��ȅ�⑾O���>���č��-����`��HC���-�I�#�ON(���9��DU��xu���Vt���|��s���ǎ�9F����]��:����J���c�н�W���e������Py�eTn��k�_(q�7�~��㊽!������G�ս�� �RN���<�wK`����ϐ������m���y������V��pc�X�G�ќ5�y�0�mz9��N��rl�n��
ǔ��D���ᠾ����Ґ��&���_�B_<��\����N߽`�������6������u�����������L#��uW��UCٽ����i�Ɖ3��,U�F�x�$b��T��������У��\��N��bg����c�TCJ���;�_;�J�G�,.`�5	�XC��]���G��Y?������q����X|���X� �6�

�� �ʿܽ�X�����$��\9��񼕽�E���ښ�r⣽�O��ҁǽ���c�����>�<`a�����S������>y���ᢾ�J������
Ky��|[���E��;���?�v�P��k�@ԅ�<��� =���%�����WF��������r�UO�Ф.�4���\���׽�F��G���>�����_�,ݜ��颽`����9�� ֽ�����  �  ��׽�$���)�f�N�}s��4������u@�����'����q���P�W&4��9!����>�$�B':�}oX���y�3n��$��h���*�������ѷl���G�)�#�o2���нƍ��m^��Cdb�bnD�&�1��'(�ݝ&�}�,���;���T���z�����/ý����&x��p8�*�]��p���������ޗ��;��K���u�h�c�H���.������H9,��2E�}	e��Â����j���X��cǏ�)"��j�a��[<�<�1���
�½�㜽�=���/\��fC�8D5�!�/�)�2���=�kzQ��Rp�%���ᬭ��W׽Z�a�&��J�F'p�1�v�������V���I��x>����e��gG��1��'���+�_�=�;�Y�A!{�,c��w'��mY��zۛ��+��#��?b�}p=�[��M����н孽�y��I턽�'u�xCj�ٸg��m�F�z��Έ�/�����'DսB����T}?�id��x���%������K��.5���d��Q:��n�g��wK��8��3���<��R�0gq��m���=���������f����	��������b�?�>�������l޽K�󏪽Wj���퓽���������ꓽ�������ez����׽�g���$��b5�tXX��w}��W���}��9Ȧ�J��������;��\����g�6�M�W?�h+>��K��~d��,���n��#���+�����(����瑾+�����[�c�8����� ��۽����髽�,��P���@���ʘ��ʡ�J��U�ŽE����� ��@�Qe�����ו�\U��bS������UΝ�,���`~���_��H�L�>�E�B�uT��mp����
R����>���l������֊��Vw��2R��90�c_�q���Jֽ�Z��e2���)�������혽 ՚��ՠ�B���F����ԽZD���  �  ��ֽ����'�9�J�4�m�yޅ�����b���X��QǄ�,�k�yL�EN0�V��I���-!�}!6��wS���s������M��%ɓ�ߎ�G���r�g�RD��9!����нmm��[���df���H���5��3,�$�*�81�W@��Y��~�fؙ����5	�P��jD5�9Y���z�(!��>%��5�������F��Rec�8%D���*�E��g��d�(���@��_�S0�j��7���M���{<���4~���\��9�������½���"���@`�H�G�LS9�p�3�9�6�G�A�|�U��St�z>��ӥ���
׽ZD�U$��AG�k��ȅ�⑾M���>���č��-����`��HC���-�I�#�ON(���9��DU��xu���Xt���|��u���ǎ�;F����]�
�:����R���j�н�W���e�����Qy�hTn��k�](q�3�~��㊽!������A�ս�� �NN���<�sK`����ϐ������m���y������V��nc�W�G�М5�y�0�nz9��N��rl�n��ǔ��D���ᠾ����Ґ��&���_�F_<��\����N߽f�������;������x�����������L#��vW��VCٽ����i�Ɖ3��,U�F�x�$b��T��������У��\��N��bg����c�TCJ���;�_;�J�G�,.`�5	�XC��]���G��Y?������q����X|���X� �6�

�� �ʿܽ�X�����$��\9��񼕽�E���ښ�r⣽�O��ҁǽ���c�����>�<`a�����S������>y���ᢾ�J������
Ky��|[���E��;���?�v�P��k�@ԅ�<��� =���%�����WF��������r�UO�Ф.�4���\���׽�F��G���>�����_�,ݜ��颽`����9�� ֽ�����  �  !�ս�9��  �sw?�#�^�rPy�`�����������T�v�$�[�/�>��f%���������*�2pE�Q�b�bh|�r���g������Ju��YY���9�T��{���н����ˎ�Ųs�
 V���B�?�8��7���=�]M�"�f�����#����ÿ��%�-�&�,�ϜL�9�j��u�������>��e��]hp��T���7�K� �`����������4�˺P�]Vm�vO���ӈ�lۈ��l���m���O�q50�4�9l�DĽ�����*����m���T�.F��*@�|C�n�N�0�b�@̀�)��璲�^o׽������ۉ=��X]�y)z�Ї�����[�������4o��kR�ܚ7�3�#�B4��,��(/�;/H�j�e��������<���l���Ki��Xq��yR��3��"�����)ӽ�����ݝ�nȍ��A����z��x�ֳ}�,���O�������q�����ؽ�A �6���5�g<U�lt�n���'��������l����cr�r�U�j�<�~_,���'�"�/�OfC��s^�b�{�F
�����)��쑾e����'t���T�,6�Ҟ�J�����BmǽF��
T�������N��D���h��!Ѥ���Ľ�޽�q������.���L��|l��C���T���`���
���(����~s�iW�g@�N�2��,2���=�I�S��p��V��<���z���K����-��/����~o���O�T�1�8H����G὿�ǽ���j���-���Lq~���S��C������nͽG�ʚ�l�n�8���W�yQw�����ᥔ�鹙�"8���i��o�
�j���O���;�[�2�e6��F�0�^��{�'����ٕ��W���4��'現� ���Kg���G��*���������ܽ��Ž����٩�uS������&��j|��p���Ľ��۽�����  �  !�׽t �s��0���I�Y_���m���q�)Ck��Z��C�h�*�@$�������a	���l�0�(�I���_�t�n��r��cl�b\�i�E�B�,�1��/S����ӽ�<��Ě�Q����.o�fJZ�ūN�ĲL��T��e�"������O���Lƽ��r.
��^"���;�("T��g���r�!Ds�f i���U�|=�%��b�*�C�����P�"�?�:��S�/g��yr�Bs�O�h��\V�.�>���$�J���-�< ʽ�լ�͉�������(m���\���U���X��{e���{������1�������۽h>������0��J�q�a�&�r�4�z��x�^�j���U�T.=�l:&�Fi�� ��y��?�|�4��N�j f��w����u\}��]p���[�W+C���)�xr��[����ڽ#ۿ�ۙ������l<��颈��ӆ��ё��H��6i��C|Ž��ld�#���$-���F��_�8u��ȁ�I��?���^3q��fZ�5�A�z,��������!�hx2���I��"c��y�1I������3p���w��`���G�E�.�������2��tӽ4��&�V[��yd���3���ԧ����|׾�Lѽ������ *��LB��[���s����*��o��]D��U>u���\��tD�\�0��z%�#�$���.���A���Y�wr�>�����D���A����u�: ^�1�D�0<,�������̟�B�ӽ����]������Kͦ�^p��;�)����Ž��ٽ������f42��K��d���{�FS��?���������V�n�o�U�%x>�:R-�_�%�ʯ(�6��HK�,d���{�����	����;��R�����p���W��>�p'�@������>轹zҽ����Wֵ������VC���_������ѽ`	�{	��  �  �⽜W ��"��#��4�PC���L���N��rH���:���'��x����Uz�е�g�����U�
�,���>�XoK��P��hL���A��82�^� ����a���@�7lƽ臯�-���$#��0�}��o�%&m�%�v�g���c����/��E ���ս���e�a��h�+��b<���I�v�P��O���F���6�@#�R0�<S���k뽘s����ʲ �6�4�<E�� O��P�e�J�3�=�`F-�sc�3
�4���#�ؽ[���y�����f����~�?�u��*y�#/�����BA��%�����νB�.X�6����%�%�7��G��hS�7X���T�͋I�V=8�'H$�s��6��P�����W������2�/QF�}KU���\��#\���S��E���4���"�����_뽨Խ����(������o�����������(��eĽt�ٽ�-�ί�Z��\�&���8��TJ�J-Y�_�b���d�]�^��Q��s>�j~*�/������
����j��v1��@F���X�W�e��aj�8�f��h\�M��;�02*���7��8s��]M轍1սܗŽ?�����������
��x�ý�Yӽ�r潖���^�
�����[(���9��tK�,:\�'ei��jp�h�o��ef�egV�B���.���<^�L��x�Nd,��@��T���d��n��Rp��j��l]�M�L��
;�b�)�����������l�Hֽ��ƽM��"��Jַ�i���lʽ*�ڽx�b���~����]8.��?���Q�.�a�'m���q��<n���b�� Q�p�<��)��ڹ��D�W-#��n4��H�\��j��+r�:q���h�5}Z��PI���7�ǵ&�y���$
��w��݋���սt/ȽgR��8��������ǽս����x����	��  �  U6����ͻ��X�X#��*�pD.�� -�qq&�`��-��OA��3�۽6�ɽ��Ľ�ͽ���L������h��G)�y�.���.�yw*���"�T��qK�F�������(�Ͻ���ү��.d��}@�������������vα�W�ƽ��ܽ5��J�������� �t�(��.���0���-��N%�]��T��x��}ؽbWʽ��ɽ�<ֽ�&�]o�yR�|�#�`�,��0�,�.�Y)�� ��`������O��!x߽Jʽ��������喽�㐽*����/�����vW��J�ֽcr�����������c<)��P1�΃6�F7��2���(����j�
�����:��۽�߽��/��U����&��p3��;�L-=�0:���3�]�*���!�Q��i��l����M�޽�8˽����\���묽�N������^ν�[㽐���@��ل����~f&��0��#9�Na@�X5D�H1C�Э<�X&1�bF"�̧��=��1��ŷ��������	�[��<9)��E8�CmC�kBI���I��7E�Y�=���4�<�+�!#"��������/�8��F�p�ҽ4�ʽ^�ɽ��нZ,޽D��a�P$���}#�^�,�?�6�D�?��^H��vN�&�P��yM���D���7���'���I���}�2�l
��b�a�%���5�dGC�RlL��P��tN���H�rg@��7��u-���#����A8��`����i�m�ӽ�,ͽ�#νɲֽa������3���I��\�&��Y0��:��KC��<K��KP���P��L�5�A�n�3��#�M��f�	�����Y��>��-��<��H��[P��>R�7!O�weH���?�w>6�I�,�o�"�����-��d�Y��%�ὦEֽ�ҽ��ս���oK�S���������  �  ,�g��������������D��*��-	�����L�܁˽|������W�����GK��j�ѽ�뽬�����d5�����|�x]�/��+{����Y������hʽo��,P�����\0���<���bؽH��|��и������q��X��dE���ND�O+��)��p��/%�RȽ9��)]��~����T���zŽ�!ݽ^l��a�����~��/����-R����L���#�Ơ��G�*i��D�ܽ�Ž2���pG��Z_��ᗺ�cϽbe�j]�G6������2� �KI"���"�UK"��_ �M��w�����& �����ѽ�½����9X����̽�S⽰����
�u6�$��נ$�f�'��7)��|)���(��s&���!�����}�������t۽&ͽ�GȽ��ͽ��ܽ+󽖃��D��6�ue&�$�+�y.�k�/���/��.�L4,�-:'��h�������ؓ���O�dvؽSսI�ܽ��|��+�����I&�{ .���2��a5��j6�7q6��Z5�l�2�"<-�%�*n�vZ��������� b��*�D�����R����$�:�.�M�5�4�9���;�q�<��$<�I�:�z�6���0���'�5�΀�i������`轻����T����i;&���/�� 6�F�9�˂;��;��};���9�K�5��C/�V�%�/��q��������	꽞N��7b�7���?�c�(�J�1�M�7�e�:��<�	�<��><��0:�-�5�b�.��%��b���-�`����U������L��� �ř �;�+�d4���9���<�->�#D>��q=�L;��q6�	�.�Ы$��~����0���L{�>�)M ������U $�m�.��  �  ��,���-���)���"�[��#l�����#��P���Iн�ͺ��}Җ����۫��~����������*���n�ֽ���J ��#
����-f��.&�=�,�C�/�^�-�~;&����LE
�����i�ڽإʽ��ǽ�\ҽ���v������!���+�5k0�ע/��w*�n�"��C�_������l0㽉~ͽ�/���,��-���M������S��	'��������ʽ~t�l�����eV���c6!�f)�� /�9j0��,��7#����R��I���ֽ��˽u>ν�޽|���h��R��oU*��3�`26��4��.�^�%�4o�z���u	��(��6w�Ncս	\��Fo��[Ĥ�P���1���­�]]����ҽH����Ut
�e���p�3+(��d1��
9��=�kg=���7��-�������� �1s��f��,�|��� �U�/��p;��-B�TC��?�ބ8���/�GC&������	��1���A�0ս��Žq�����������u̽�޽����D�!L������$��.��Y8�xGA��*H�ceK�K�I��^B�&M6�lB'�-���B����M���>�`���#�|R3�&�A�Y�K�<rP�˪O��xJ�~uB�p&9��}/��%�C���'�n=�u��a��W\ս�9ͽ&�̽��ӽ;���b�����O��I,��3$���-�^�7���@�N I���N��$P��3L�}�B�L5�%����C3
��;�P�Á�lH��)�	�8���E�5&N��P���N�6MH��?��h6�P�,��&#���`��q�����o�òԽO:Ͻ��ѽ%Q۽z&�
���X
��9�*����)��Y3�c�<�q)F�U�M�J.R���Q�+L�G-A��p2� q"�z"��3
��w���	��Q'!��B1�Pl@��L��  �  �ZN�`L��cB�&�3�W"�jd������7�ǽ�P���国S֊�E�{�z�k�"bg��o�3����2��qY��7�����ν�O�[���[�'�˹8�w�F�4O�ۺO�H��#9���%����� ���콸�������	�����O1�|�B�`�M�*Q�1L�`y@��m0�G���%��*��<�ݽ�Ľ.���<��*��
;}��p�y�o��{�$���ꗽ�������[ڽCL��L�
��V�\+.��>���J���P���N��eD���3���������&��ｿ�[��u'���;���K�S	U���U�F�N�KsA��0�	�����F��ٲʽ6е�y.��Pu���y�����!����)��z����T���Wɽ	6ὗ������-��}p/�A4A���P��D[�˸^���Y��lM�`e;��^'�yY����f�`��@I���'��n<� �O�Mv]��c���a�� X��:I���7�h9&����`
����z8ݽ�[ɽ�𸽻����|�����ô��~򲽻���E�ԽO��������e:�{g0�t{B���S��b�_�j�3�k��8d�L�U�6�B��'/����U���I�~�.)�Ģ<�-!Q���b�`�m�7q��=l�t~`��dP�ɉ>���,�]���h�������ؽ��ȽGS�����������-��E$ǽG�ֽ˼齦���1��<����*�
�;��M��J^�Z�j�p�p��\n��d�(<S�2 ?�%�+� ��}�����ɕ�Q�/�JD���W��xg��)p�A�p��)i���[���J�C9�(�'������
�N�����Y�ս�+ǽ�l��7���	����½�kϽZ�m���>�U%���!��w2�mAD���U�pae���o�v<s�Ln���a��OO�� ;��(�����	����5'�E<9�īM���`�� n��  �  �xq�_�l�.^�D�H�p}/�:O�l�����ֽ�2���ț��䆽{n���W�(�J�1G�3HM�!]�
v��E�����	���1!ήF����6��MO�2�c�a�p�ps���j�*�X��@�$=(�q������[�V��у�U6��N� #d��;q���s�pk��Z���B��y)�����P����Ͻ8J��,����Y��k�m��8Z��O�gPO��mX���j�oI������~歽�˽?H����rR&���?�DhW���i��s�e�q�Rf�x�Q��^9�[�!���[_�~��P���(�*B���Z��#n��Vx���w�D>l���X�H�@��['�����l���ҽӶ������Ϗ�nɃ���x��s�_x��R�����"n������gJϽ��､��̷"�9�;�S^U��k��|{��ڀ�
 }�#n�7X�5y?�"@)�L���,�/v���(�9?���X�[�o��*���c����(�s�b0^�->E�-",��*��~�N��0�Ƚ�\��� ��d����㔽��◽�����ԭ��ɿ�9�ֽ'O����K�7�	�Q�qlj��W��#o��pb���Ju�^	^���E�{�1�x<%��:#��,���=��U���n���������鉾h����z���b��aI�r�0��d���	o��׽<Ľ#���oӫ�,���GK���ت�<������ֺԽ9���Y�l���s-���E�{�_��,w�"����s���׈�����cq���X�u�@�g.�B�$��+&���1�pF��^���v�=߄�N���m,���`���s��Z�%]A�dg)��q�����w齩�ҽ�C������g�����􁪽rӰ�sǻ��j˽��^��s)�	� �(�7�2�P�Cj��4�����/��֬���$��sl�5S��<���,��&��+���:���P��i�nj��̃���  �  NU��/����w���\���=����b3Խ�����!��c(t�ĽT���?��a4�Q\1�#�6���D���\��%�%{���<����P@	���&��CF���d�}~�;N��/$�� \��$�s��5X��o;��G#�Xa�U��o�	0���K�*�h�P����"��UR��'��'r�GMU�q�5���f����˽e���n��+�p��U�RC�C:�E�9�A��;R�1�l�H�������%ƽo������1��Q�V�n�|҂�{鈾̄��}���5�k�\9O�"�3��W�����x�I�#�t�;���X�;�u���4Ƌ�튾����o��Q�Ό1����:��x�˽�������A����Go�&Hb�E^�ZYb�1o�.�������q֨��bƽ��=�rQ*�͕I�Fi�^t���V��Qk��㍾7C����p�$T��
:�.�'�_Q!��h'�2)9�FES���p�텾�r�������ԏ�z����r�B�S�c[4����$ ��0ڽ�
������k���{َ�}։��$��T���&���� ���#����˽����
�0�#��{A�\@a�f
��]匾���&��~{���I���`u��Y��eA�Q�2�\�0�خ:��O�XFk�8��(����)���\������/��!Iu���U���6�����(�	��}p˽o^���K��EF��<����h���b���ŧ���?YȽ���>������.3��Q�"<q�&T��Ṓ�ј�mh��f�������!�n�5�R��H=�C22��3�`mA���X��u�ڈ��ԓ�%_���U�����������(k��K���-��[�����޽�-ƽ@v���c�����k+���|��X��P6��i����%Խ�$�:m��#�H1?�la^��}�oˌ�E����������9U��fW����g��]M�.�:�"�3���9��$K���d��
���l��6ϗ��  �  t"��xm�������k���H��b%��g��ս"�������Pg�I2G���2���'�\%��0*���7��N��Ir��[��wӴ���)F��S.���Q��t�~����͑�*�k����;���h��aH���-�~v�eb��3%�]�;��Z�b�y�释�/Ғ�����̭����b��-?����r��Vʽd��o���c�݌G��26�;�-��"-�"�4���D�"\_�xt��IS��K Ž0��������:���^�ױ�ݰ��m���Q=��^����v}�<^�/�?�@(��f�j���-��<H�>h�烾x?������`}���L����1]�ð9��v�����N�ɽ��������ix���a��U�,�Q��U�O*b���w�����I(����½��콳�9�0���S��{w��j��P����5��w��o����ƀ��a��PE��l1�*���0�+D�R�`�i����z����ĝ��&��wя�"����V^��2;��P�� �}	׽���t���ἑ�eN��v��������h�������`��������ƽ������(�2I�"�l��܇��X��:����ࡾW֜�W�������7f���K�<�^X9��{D�g[���y�V쌾{����ڢ�������������f���_�̅<����}���vrŽ���*���6ҙ��}���5����������a���9½�/޽���to��_8���Z��N~�񽏾���������"��ƚ������}}��^�%;G�k;�V�<��K���e��|���������\(���碾ɐ��X����Vw��S�,[2�0�����ҹٽ�ֿ�����3����������L<������Us����6tνb��k����%���E���h��������ݠ�t��á�����F����u�d�X��nD��<�7C��*V�wr��C�������P���  �  R)����۾�M��D𡾶���R�٨&��k��4ֽQG��Ι��<���߁��p�G}��@����I��>W��d�ὠ���0�^�^����0~��?�Ǿ��c�����3n�B׾Q��ՠ�f ���x���r�������:���˾���B���������oԾ<��������w�OGE�?x�h����ͽH(��̻������'��{ǃ��a��ե�����sȽ&���.���?�6q��V��"���a�оɏ����L-�F�徹�ξ���"���ϒ��W�t���w���__�����l־��4��#*���q� ξ$���Y���Sl�(&=���������Ͻ�������F������1���is���E��˴ɽ5-��n���0��;\�=n��4����ľ�8���K)��C'��$�;~T�������s�����������#����˾�徇������LF�����5*˾�Ҭ��쎾}�h��<������u�߽��ǽ�'��r����Y��^ ��� ���yҽ�C�?�&��XK���y�7���z	��0վ�����Ch����G���˾௾�M��^����#��Gw�������"���ܾ��b��{����E侂�Ǿ���M틾�Ge�=^<����A��s�i�ֽ��ɽ2ýt�½cdȽ��Խ$�������i�7�ڟ_�ߋ��RR��)�þJ��M���z��������S�޾þ]���vO��N��J���!��5���zɾť侮	���n�N����4C۾���%%�� +��A	W��1�rj�.�?a潩Խ�lɽ�BŽ�ǽu�ν}�ݽj����0�p�$��F��,q��ْ�1���3,Ͼ#��UG���8��� �:=�׾O(��5>��$����j��U�������]��V>Ծ��(8 ��  �  �}�P�"Zվ��������Ձ�0kP�&����v�ؽoM�����|g��_섽縂� ���Ґ��}��SD�����B]�ޡ/�R@\�ë�� ڥ�1�¾��ھԅ�()��zѾ驷����Z���s��n�n�����˫�Ŭƾ�ݾ����z��I�ξ�o������t�n�C��@�����ϽII�����񭍽F-��Dˆ���ݘ���� /˽������XT>���m�ނ���篾��˾�q��=�E��E�߾�hɾ.ʮ��H��Fс���o���r�N#��_�>i��y�о���Đ���S��ɾ�������8ei�<�������ҽtӷ�G��"]����������/���P}����̽9��K�0{0��&Z��_�������W���ھ���~��ګ�GྠȾ"O���b���ׄ�M[}�O����链8���H�ƾ��߾8���+�����-�H�ƾ�t��þ���Pf�V<���5�����(˽^Q������QX�����/ý/�ս`.����&�_J�#w��*��me��.CоJ��BV��'��:U�W�߾�kƾ{%��dV�����ȹ�����P���'绾@�־e��r4���S��\���޾�þu������c��&<�-��������j"ڽ��̽i7ƽ�Ž��˽��׽�3�N.�+��&�7� ^��ن�a~��u��۾���4V��������>pپڿ���$������v����ӈ�5>����9�ľI)߾���8��|��-��L־չ�����˳����U�?�1��i��� ���A׽�̽�CȽ�ʽҽ/'�Ч��bl�qW%�ڔE�Io��ː��]����ʾ��4���/���F���Aa꾁Ҿ=#��4��[�����Q,���霾�r��u`Ͼ�W����  �  $�ھ�nվ��ž�7��򁕾�Ex���J��%�-����oH���V��Ga��p������*��r暽jЬ�ǽ�O뽝	���-���U�q@������m��P�ʾ��ؾ7�۾v�Ӿ����X�������[}�n�d��R`��ap��"���蟾�%���̾;�پ��۾ĄҾ�$���������j���?�0����3�ؽq~���3���}��ݖ���.��aA��1���]���qԽJZ������;��,e�����0ꤾ�`���оZ�ھ�=ھ��ξ����𠢾n���/t��6b�ce�g�{���������y����rԾ�޾��ܾ�о����
�������
b��9�N^�k� �mܽ�%½�i��2���W���(��T����ƾ�R�ֽ�0�������/��1U�k���J��5��m˾�ܾ� �]�޾k�Ͼ�������2d����z���o�9qy��&��𛠾����Ͼ�߾S���4ྈ�о��`e��c����`�O;�+^�����콡wս�Gƽ�+��T���.����;ͽ`�߽(���+��g�(��H�fp�M���=����þ��ؾ8Y�X�� ���Oо|U��D����P���������!��� ���OȾsݾK��B��ͼ�sUо76��j4���s��*�_�Xp<�B� �������]a���ֽ[�Ͻ�0Ͻ9Cս��st��5�	����wz8�n�Z���������﴾kn;�����S�}�޾��ʾ���Iq������@����ҁ����_��y*��t�Ͼ]Y����e���fݾ��Ⱦߛ��S˕��|�ߕS��3����j����b��)ֽ�ѽY�ӽ�ܽt��\�����'�AE��$j�,s��_���������վq��I�����پ�ľ�ӫ�����9��{ㅾ�#��
k�������3ؾI��  �  Ɍ��j��������^��� kj���E��&��s�3x򽌰ҽ;w��!W��?O������<���$������?ڽW��3{��+.�6�N�q}t�ᎾY/���B������2�����~'������3����d�u�O�~�K��Y��Rv�}z������v����y��U����h��]ӫ�a����ڃ��`��'=�I ��i��K�Q�ͽ����"���=���Ǡ�٭��˼����ʽ�2罧�����>69��o[�ON����������Ҹ����������\���ϐ���z���\�ìM�B!P���c�Q�������P��^O��:�þ	�¾t�������ɔ�[/���:Z�Za9��]����8��'�ս��½5���ݲ��ﵽ�P����ѽ2@����/��C2�e�P�*>u�<䎾❣��$���\þ��Ⱦ�ľX&��	ť�I`��]'~���d�a[���c��T|�)j��I,���Y����ž@˾�2Ǿ�躾���l�������[���<���#�ͨ�� �Ĕ轁8ؽNϽ-"ͽz�ҽ�k߽/5��	�L���-���H���i�ݼ��l��^ɰ�J���F�̾�+ϾTKȾ����63��,��=|��m�n��!k��(y�� ������Z"���ľ#�Ͼ*�Ѿ7�ʾ���¨�`����� &]�b�?�:5(�]\����)��"�F���߽���C�������.�1t%��y<�X�X�+N{��G�����X���Q�Ⱦ��о� о�ƾ7��u������l|�˥l�Ȭn�&ꀾ�Q��|�� y��y/ɾ�OѾj<оdƾV(䡾�<��;t�'AS��8�X;"����������W�N$��U���My��8�ծ�І.��aG���e�����J��� ��4���:�;��Ҿ��ξ�B¾����W6������c�w�n��v�d#��{4��Rɭ�y���Kξ�  �  �2��!���ޘ����%�|�#J`�u2F�G/�:���	�f�򽙞ؽ4�Ľ�����'���ݺ�Y&ɽ��޽.���؅�� ���4���L�H�g��A��fM��{����	��.���z���E��Dx��rbb��+G��m6��H3��T>�2�U���t�缊�,��������:���b��(��F�u���Y��@��[*���������\<սt�ýT��Շ��#����ҽXJ�߸�&��¹'� �=��FV� �q�fM����������&��˂��c��}o���^x��$Y�|7A��!5�;67�	'G��b�_���1ޑ�7�6��.���XU��=8���t���Jr�}cW�Dh?�@l*��	�X��:���9'߽Uѽ�z˽{Ͻ�g۽����������&��L;��[R�=al��c���Ò�5����_���^���|��d-���b��c|��^�C~J���B���I�<�]��!{�XC��&��������魾�ܫ�����si���9�� v�;\��!E�\1�q���0\���;�X���9��Y������"�F�'�V|:�ïO��g��[���ˏ�睾'����ְ�����������9!��|����e�N?U���R���]�cu��O���ܚ����6O���Ǵ�Yo������bL��Lڊ�)�y�р`�->J�;�6�Um%�st��3
�yY�k��|���* ����خ��L#�94��lG�G]��"v�%����N��"ˤ�*'���6������!���e������x��q`�3�S��U�Ze��t�$鏾V���0Ǭ�	ҳ�h��������c��Ɏ���1��aq�eDY�zD�P~1�J!����
��� ������o���{�p*���%�*�S<�wnP��Tg�ݟ��sˎ�o'���᩾c���쪵�^���}K���_��j懾-r���]��U�d\��o�uU���ږ��-���I���  �  �����������\}�[�n���_��	Q��	B��d2�m�!��O��������ڽ�dֽ�ݽ�F�V��K���b&���6�mF��}U��d���s�G󀾜���ED��X܇�������o�W�U�=���(�s�d���2"��	4���K���e��C|�5��E���ß��;-���5{�\_l��X]�DnN�5?�E7/������ߡ���8�H�۽:۽a*潈������p�b-�5#=�W^L�
<[��2j�;y� A�����wo��灆�1~�%Ih�=O�P7�t�$����B�D�)�\y>�	X�q�q�M���`J���p���W���#���|� �m���^��P���@�	�0�~m ����no�r��o����Zv �=������-���>���N�@^�,]m��|�Ѫ����Oя��a�������gn�w,U���>�o4/��)�^�.�lT>�8U�^o��ă��+��YR���ⒾĈ��!����Z����u�;�f��X��H��^8�i(����!���G��j����0�*�_/��@��?Q��a�%Qp�}��[������$>�����SΕ���8C��?t�o�[�3G���:���8��A���S�X�k��Ⴞ�I��E��ř��ј�Y��k����F���m}��hn��_� O�{:>�Z�-�i��G���d����B�O�+�<�m�L��\�k"l�f{�k������DG�����z��	����������n�tV�|�C�@G:���;�joG��[�¹t��iW���ߗ�Lי�񚗾�M��?X���܃���x���i�}Z�$FJ��9�)�l���E�~�����B�Kr#��2���C�K)T�)d�Z<s�R����������U���*���;��zƕ�l ��A2����h��R�)4B�i.<�t&A��1P���f�e���,���p���  �  Ub�O�i�!dm���n�B�n�W{m�ϭi�"b���U�1E�@�1��A� ����q���@��Y���"��6�7�I���Y�/e���k�?o�{cp��6p�}�n�(j���a���T��{C���/�"������Y��������@��\'��Q;�]N�N@]�^�g���m���p�Bzq��q���n��i���`�\�R�;A�0-��K��g����΂�
�G�	�*���>�y�P�V5_�e�h�A#n��pp�_�p��Gp�=�m��1h�T^��O��=�5�)�¾�S)
�@s�`���5�����1��F��HX��ef���o���t��w���w���v��)t��n�̡c���T��B���.������76�����s���(���<���P��[b��o���w�]N|��~��`~�zQ}��z��Ks���g�i3X��OE�6�1�5!�ƣ������5J!�N�2���F�iZ�2Fk���w� >�����L��lU��ܩ��P���x�.l�(�[��tH��J5��2%����(����V*��B<�K�P�d�"<t�����_�����n���w���턾܂�J�}�� q��%`���L��;:��
+���!�c� ��L'�5�4�OG�.t[�UWn�I�}����|��y���݈�b���փ�������Z��%�r���`�L�L���9���*�{"�� "�)���7�YJ�\@^�Rp�r�~�H������,���y���&��t醾����U~�b�o��V]�sI��7�()�g"��#�D�+��;��)N��b�S�s�����?<��h���M���舾�{������􃾭@}�x�m��&[�SG���5��(� �"�]2%��E/�Z?�T�R�C�f��w��V���r��y���)w��4���9
��Dc��:�6v|�{ul�rOY��E��r4���(��+$���'�D3�Q�C���W��.k�C�{��  �  �^B��~Q�|�`���o��1~�W��JZ�����y���'r�|�Y�k�@�H�*�78�� �T���B/�	vF��&`���w�cv��m�������ߐ��;�|�m�m���^�hP�i�@�1�ߏ ����7� �+��ܽ�rٽE��\���BY	�֐�/_*��:�)J��Y�h h��)w�}��������ˉ�c����݀��l�}lS���:�6�&�_p�#����$���7��fP���i� u��솾����g����eOx��Qi�LZ��bK��<�7,����A{�����[Gݽ=�߽i��7��2Q�zl#�i�4��
E�,�T��c�?/s����䱇����팾HS��zR��3l� �R���;�#�*�dJ#���&���4���J�g@d��W}�����
����菾�!������i���q�wc�0T�X�D�̲4��F$���?�p_��-���������V����%�77�o�G�P�W�b%g�Bv������ �����tO��µ�������J����p���W�]�A�2�3��#0�nK7�.H���_���y�kֈ�W�������ߕ�����ǋ�(���U3z���k�p�\��LM�a(=�g-�w�Q�K�����Ƴ�g��8)�ƣ9���J��Z��pj��ny��6�� ���癒���Aƙ�0���-����*��bs��/Z�/FF�L�:�MJ:��nD�qyW���o�먄�B���l�Lv���֗�7풾� �����*Pz��dk�k\���K�2A;�n�*�v��Z�1�����f����*�.�Ca?��P��`�Z_o�k\~�����-�����j���Ι��������������k�T�ƺB���:�>���K�B�`��Sz�����Xe���1���j��ؕ��*둾CЊ��Q���w�P�h��KY���H�H8�g�(��q����5f��&�Ʉ�AZ'��
7���G��gX��  �  ��/��3G���a�N1~�TT�����������`��rD��v�����9f�E�I���6�O|1��B:���O���m�Os���C���m��[��Ԡ�ɗ�S���Py�B4]��C�^�,��%�ũ�!��x�׽��Ľb�����'E����ν3��U
���~$��9��HR�q�m�k/���������������6��~0���~���]��D��j5�Y�4�P�A��Z��@z��d��⚾��91���Ğ�(�����j:p��T��<�΁&������Kv齱�ҽ3ý����/!ɽ0Fܽ�"���
��v���0�Z>G���`��}�8��@C��h���q���\���
���э��{�Q�\�B�F���<��FA��5S��`o�9F��t1���U��De��9|���>���y��Ls��,\t���Y�|\B���-�a��5�����"X�яܽ�pؽ�vݽ 3�8C ���a7��0��TE���\�fYw����(=���~��b����d���^��a&��8㎾�A}�a���N�b�I���R�h�h�B���W>��
:��늭�CP��Z,��R6���y��/9��/�x��_�"�H�dH5�C3$��g��>	�] �N�������������8���!���1�E�D�8Z�9�r��憾1K��j
�����������������܎��}���c���T��T�Ha�Vz��⌾v+�������Ʋ����Ϫ�����g�������t�{\��jF��_3�b�"�g$�׀�` �q�������.���	��r�=�&��7�.�K���a�[{�����u���B���尾�촾�������R��)����#u���^�xT�x�X�,j�~�T����������� ��/���^栾�ڒ�'�����n�.�V��JB��0�� �W�����>�����_� ��[���� ���.�t	A��  �  8�'��RG�4`l�����g4�����������F0��`_���<��ą�Ch�½P�v�I�N�T��bo��p�����Be��ԥ���@��枻�����z��v͆�Jme���A�ӗ#�
+��j���нr޹�⩽����x���P��}]��8xƽ��὾~�j��SP4�_�U�(I|��ߒ��֦�l��Y|����,���{���e���]����`�1XN��TM��]��|����kG��x궾�j��"���nI����6��� 0��f\Y�0k7��O�a���彏Cʽ"���.������e\������
��z�ֽG\���1��&��bD���g�S��~�������_���ž<�¾6����᥾����Z>}�Z�a�ARU��Z���p��䉾���:?��~����ǾvQžnA��������.8�� [�X#;��!��>������߽�ͽ�ý�忽m(Ľ%�Ͻ�F⽸������Xh#��^=�+]�R��������y����Ⱦ �˾�KƾV���D��� H��}g��qh�S�a��,m����	���̫�EQ��V�ʾvξ��Ⱦd���w���
[��Z���']�9[?�D'��2�Oc�@���u�形�ݽ�ܽ�㽹L�>��B����"��8�n�T��u��E��F���涾�Ǿpsо8�о}`Ⱦ�Q���4���%��j��|�m�_�l��2}�%��Iơ�=���ƾ�=о"�оO-Ⱦg���餾�(��oQy��ZW�6.;�xx$��v�>y��9��M����>὆D����0����'�)�ڃA�C_�8+��"���멾<��PI˾��Ѿ�sϾ�!ľ[���۝��Ǌ���y���l���q�Vރ�T'��\���&����˾fuҾF�Ͼ�ľ�r���������[�o��O���5�� ����=�k.��������Yp�s)�|����I5���3��  �  �s&�	�L�i�z�o떾⠰�oǾ�6־�7۾��Ծw�ľ�����Ǖ�u߀�Zf�"P^�Ek��*���A������Jɾ�׾e�۾�5Ծ<+þ�ȫ�鑾c�q��zE��� �IV��Oݽ�t���禽�!��3D��!���韽����ν����;��I5���]������ᠾ�Ṿ�@ξ�Kھ�۾��Ѿ����ަ��;����x�r7c�@b��Fu�0Ō������:�Ͼf�ھp�ھ5�Ͼ�=��j��������b�i�8�������mӽ�붽���{�������є�� ���Q��[)ý��P��_#��gG��0s�!���͠��q�ľ��־ld߾��ܾ�ϾUݺ��Ȣ�#q���Jx���i�1p�����׀��;α��ɾ��ھK�S�޾��о�������i󇾛wa��l:��b������佛�˽�U��o���j���D�������"Ͻ��C��>X�B<��b��C���ҡ������Ѿn-ᾼ=�P �v�Ͼ-T��L������/	~��Uv���������˧�RQ���-־���;��k�ᾂ�оT?��Vs���z����`�a�<�h ���8�����n�ӽ��̽qN̽�:ҽ�޽5x�2N���+4��DU��D~�������@�ɾ�B޾TA��i�7j�Vtξ%���n����[�������`������#Գ���˾ ~߾����]�߾(̾8��L���`I��!�X���6����{
	����0�ό4սɄϽ(Sн��׽��j����M�le"�U>��b�<ˆ���������{�Ѿ���Z3쾡��@WܾsPǾ�������- ��z���A����m��Ǥ��弾�Ծ<M�n��=�۾�kž����W���1v�vO�:�/���P�X6�f���׽7Խx�׽�!���B��~��-��  �  ��'��R�+B��
-��Q��x�־��羿��|�澈�Ծ y������r�����t���k���y��E�� ���U���T�پ���8�|�徵AҾ����Xe���|�|%J��I!�ˬ��ԽIX��t����<��φ�>����f��MÕ��è��:Ž���u���7���e�`�;L��դǾ�޾hw������6�;�}���P���f���'q���o���������f��M�ʾ���-,�D�o��Zʾ�[�����j��;��D��M���ɽ˶������,N��)Ή��z���^���!������-ڽ�,��K#�Y�K�s�|�ͬ���4���cӾZ�����h&�B���Cɾ3���Eʕ�����tw�E~�km��������ؾ�:쾣���R������	Ⱦ�2���/��'�g�&<���������ڽp���zI��fz����������#�Ľi�޽s��;;�P+=��`h�"%������;Ⱦ�����������F�߾��ƾ0��*7���=�������(������:���cξ/�������8�����[�߾;.ž_����p�e��=�����E�:׽�ɽi@ý"�½�{ȽE�Խ�软�������2�(�W��������c��h�׾���>l��=�������ݾ�Kþq��)��%S��/����J�� W��'���ھ$���������o��sCھrL���栾�r����[��6��V�m]��9뽾q׽�y˽�$ƽ3�ƽ��ͽ�۽�|�}���|�"<>��)f�o����ħ��8ž�V�����ɟ������Ȳվ�Ӻ�-졾纏�l����Ɗ�i䘾rd��ʾ>��e����n��F'��	�^yҾ����������|��P��
.�8��g�k��o�׽[]ν�'˽f�ͽ� ׽z��K ��l��+��  �  �T(��U�X�����������#gܾ�f�#g���$�Xھ[I��މ��u�����y�6�p�k?���>Ȫ��ƾc�߾�L�E���7���׾@��O������: L�
�!��	�BҽCC���d�����Hƃ������N��펒�����d½)�뽏����8�(�h������$����̾�����_�����
HӾ�����䜾�A���v�O�t�Y��,���ɴ��Rо�����󾧳󾫶�~�Ͼ�W��괓�)@n��\=�4K�����ƽX����[���9���҆��{��wC��������׽�t�q�#�MSM��N������u����ؾ~ ��{������c~澿fξK������p���A|�줁��j���ߧ��þ�|޾Y��u��W���k�g�̾4Ů�N���4~j���<�9�]s����׽VK�����j��H��T���4���������۽� ������=���j��c��������̾�U��]���m��B����d�˾I�� H��RɈ��Z��Xɋ�oԝ�PJ���gӾ���O��	� ��/��v���ɾ���آ����g��o=���Ny���齎�ӽF�ƽz1��Cؿ��]Ž^Nѽ��佖�� ���2��Y��|������?;���ܾ\���2~��>�w�������Ǿ���T���Ɗ�Z�����'ө�L�ľ5྿���������B���mi߾�G¾�������@]�h6�fs�@����|;ԽC^Ƚ�!ý��ý]�ʽxXؽl_�Ї����>�t�g��~��U̪�yyɾk�從������N1���4�ھX ��;���i�����;I���⛾>)����ξ�j��W��n��� �A��+@׾;/��O�79�ƋQ���-�) ��������Խ!L˽d'ȽA�ʽ�ӽ�B�9���~E��1+��  �  ��'��R�+B��
-��Q��x�־��羿��|�澈�Ծ y������r�����t���k���y��E�� ���U���T�پ���8�|�徵AҾ����Xe���|�|%J��I!�ˬ��ԽIX��t����<��φ�>����f��MÕ��è��:Ž���u���7���e�`�;L��դǾ�޾hw������6�;�}���P���f���'q���o���������f��M�ʾ���-,�D�o��Zʾ�[�����j��;��D��M���ɽʶ������+N��'Ή��z���^���!������-ڽ�,��K#�T�K�o�|�ˬ���4���cӾW�����f&�@���Cɾ2���Dʕ�����tw�E~�lm��������ؾ�:쾥���T��Ý��	Ⱦ�2���/��+�g�*<���������ڽt���|I��gz����
���	����Ľe�޽p��7;�L+=��`h� %������;Ⱦ����������D�߾��ƾ
0��*7���=�������(������:���cξ1�������8�����]�߾>.žb����t�e��=�����K�:׽ �ɽl@ý%�½�{ȽF�Խ�软�������2�(�W��������c��h�׾���>l��=�������ݾ�Kþq��)��%S��/����J�� W��'���ھ$���������o��sCھrL���栾�r����[��6��V�m]��9뽾q׽�y˽�$ƽ3�ƽ��ͽ�۽�|�}���|�"<>��)f�o����ħ��8ž�V�����ɟ������Ȳվ�Ӻ�-졾纏�l����Ɗ�i䘾rd��ʾ>��e����n��F'��	�^yҾ����������|��P��
.�8��g�k��o�׽[]ν�'˽f�ͽ� ׽z��K ��l��+��  �  �s&�	�L�i�z�o떾⠰�oǾ�6־�7۾��Ծw�ľ�����Ǖ�u߀�Zf�"P^�Ek��*���A������Jɾ�׾e�۾�5Ծ<+þ�ȫ�鑾c�q��zE��� �IV��Oݽ�t���禽�!��3D��!���韽����ν����;��I5���]������ᠾ�Ṿ�@ξ�Kھ�۾��Ѿ����ަ��;����x�r7c�@b��Fu�0Ō������:�Ͼf�ھp�ھ5�Ͼ�=��j��������b�i�8�������lӽ�붽���x�������є�� ���Q��Q)ý��J��_#��gG��0s����ɠ��m�ľ��־hd߾��ܾ�ϾSݺ��Ȣ�"q���Jx���i�2p�����؀��>α�ɾ��ھK�X�޾��о	�����n󇾣wa�m:��b������佢�˽�U��r���j���D�������"Ͻ��=��7X�:<�݋b��C���ҡ������Ѿi-Ᾰ=�L �s�Ͼ*T��	L������-	~��Uv���������˧�TQ���-־���?��o�ᾇ�оY?��[s���z���`�i�<�h ���8�����u�ӽ�̽uN̽�:ҽ�޽7x�2N���+4��DU��D~�������@�ɾ�B޾TA��i�7j�Vtξ%���n����[�������`������#Գ���˾ ~߾����]�߾(̾8��L���`I��!�X���6����{
	����0�ό4սɄϽ(Sн��׽��j����M�le"�U>��b�<ˆ���������{�Ѿ���Z3쾡��@WܾsPǾ�������- ��z���A����m��Ǥ��弾�Ծ<M�n��=�۾�kž����W���1v�vO�:�/���P�X6�f���׽7Խx�׽�!���B��~��-��  �  8�'��RG�4`l�����g4�����������F0��`_���<��ą�Ch�½P�v�I�N�T��bo��p�����Be��ԥ���@��枻�����z��v͆�Jme���A�ӗ#�
+��j���нr޹�⩽����x���P��}]��8xƽ��὾~�j��SP4�_�U�(I|��ߒ��֦�l��Y|����,���{���e���]����`�1XN��TM��]��|����kG��x궾�j��"���nI����6��� 0��f\Y�0k7��O�`��	�彍Cʽ"���.������^\������
��l�ֽ6\���1��&��bD���g�L��w�������_���ž7�¾2����᥾����V>}�X�a�@RU��Z���p��䉾	���>?�������Ǿ}QžuA��%�����48��,[�c#;��!��>������߽�ͽ�ý�忽j(Ľ�Ͻ�F⽬������Oh#��^=�]�K�� ������r����Ⱦ�˾�KƾQ���@����G��yg��qh�S�a��,m�������̫�JQ��[�ʾvξ��Ⱦk���~���[��Z���']�D[?�D'��2�Wc�L����彪�ݽ�ܽ��㽽L�?��C����"��8�n�T��u��E��F���涾�Ǿosо8�о}`Ⱦ�Q���4���%��j��|�m�_�l��2}�%��Iơ�=���ƾ�=о"�оO-Ⱦg���餾�(��oQy��ZW�6.;�xx$��v�>y��9��M����>὆D����0����'�)�ڃA�C_�8+��"���멾<��PI˾��Ѿ�sϾ�!ľ[���۝��Ǌ���y���l���q�Vރ�T'��\���&����˾fuҾF�Ͼ�ľ�r���������[�o��O���5�� ����=�k.��������Yp�s)�|����I5���3��  �  ��/��3G���a�N1~�TT�����������`��rD��v�����9f�E�I���6�O|1��B:���O���m�Os���C���m��[��Ԡ�ɗ�S���Py�B4]��C�^�,��%�ũ�!��x�׽��Ľb�����'E����ν3��U
���~$��9��HR�q�m�k/���������������6��~0���~���]��D��j5�Y�4�P�A��Z��@z��d��⚾��91���Ğ�(�����k:p��T��<�΁&������Hv齭�ҽ�2ý�����#!ɽ!Fܽt"��ڧ
��v���0�L>G���`��}�0��8C��`���j���\���
���э��{�L�\�?�F���<��FA��5S��`o�=F��y1���U��Je��@|���>���y��Us��;\t���Y��\B���-�k��=�����+X�Տܽ�pؽ�vݽ�2�3C ���W7��0��TE���\�WYw�	��� =���~��[����d���^��[&��4㎾�A}�a���N�b�I���R�m�h�E���[>��:��񊭾JP��a,��Z6���y��79��?�x�_�/�H�pH5�N3$��g��>	�] �X�������������:���!���1�E�D�8Z�9�r��憾1K��j
�����������������܎��}���c���T��T�Ha�Vz��⌾v+�������Ʋ����Ϫ�����g�������t�{\��jF��_3�b�"�g$�׀�` �q�������.���	��r�=�&��7�.�K���a�[{�����u���B���尾�촾�������R��)����#u���^�xT�x�X�,j�~�T����������� ��/���^栾�ڒ�'�����n�.�V��JB��0�� �W�����>�����_� ��[���� ���.�t	A��  �  �^B��~Q�|�`���o��1~�W��JZ�����y���'r�|�Y�k�@�H�*�78�� �T���B/�	vF��&`���w�cv��m�������ߐ��;�|�m�m���^�hP�i�@�1�ߏ ����7� �+��ܽ�rٽE��\���BY	�֐�/_*��:�)J��Y�h h��)w�}��������ˉ�c����݀��l�}lS���:�6�&�_p�#����$���7��fP���i� u��솾����g����eOx��Qi�LZ��bK��<�6,����?{������RGݽ3�߽\��/��(Q�nl#�\�4��
E��T��c�-/s����۱�����팾AS��tR��)l���R���;� �*�cJ#���&���4���J�p@d��W}���������菾�!������i���q��c�0T�e�D�ײ4��F$���D�v_��.���������P����%�-7�b�G�A�W�R%g�	Bv������ �����kO�����������J��{�p���W�X�A�0�3��#0�pK7�$.H���_���y�qֈ�^�������ߕ����ȋ�1���g3z���k��\��LM�m(=�q-�w�X�Q�����ɳ�i��8)�ǣ9���J��Z��pj��ny��6�� ���癒���Aƙ�0���-����*��bs��/Z�/FF�L�:�MJ:��nD�qyW���o�먄�B���l�Lv���֗�7풾� �����*Pz��dk�k\���K�2A;�n�*�v��Z�1�����f����*�.�Ca?��P��`�Z_o�k\~�����-�����j���Ι��������������k�T�ƺB���:�>���K�B�`��Sz�����Xe���1���j��ؕ��*둾CЊ��Q���w�P�h��KY���H�H8�g�(��q����5f��&�Ʉ�AZ'��
7���G��gX��  �  Ub�O�i�!dm���n�B�n�W{m�ϭi�"b���U�1E�@�1��A� ����q���@��Y���"��6�7�I���Y�/e���k�?o�{cp��6p�}�n�(j���a���T��{C���/�"������Y��������@��\'��Q;�]N�N@]�^�g���m���p�Bzq��q���n��i���`�\�R�;A�0-��K��g����΂�
�G�	�*���>�z�P�V5_�e�h�A#n��pp�_�p��Gp�>�m��1h�T^��O��=�3�)����P)
�<s�Z���5������1��F��HX��ef���o���t��w���w���v��)t��n���c�t�T��B���.�|����76�����s���(��<���P��[b��o���w�oN|��~��`~��Q}��z��Ks���g�u3X��OE�=�1�;!�ɣ������1J!�G�2��F�iZ�$Fk���w�>�����	L��cU��ө��?���x� l��[��tH��J5��2%����(����V*��B<�U�P�d�0<t����`�����w�������턾!܂�Z�}�� q��%`���L��;:��
+���!�h� ��L'�8�4�OG�/t[�VWn�I�}����|��y���݈�b���փ�������Z��$�r���`�L�L���9���*�{"�� "�)���7�YJ�\@^�Rp�r�~�H������,���y���&��t醾����U~�b�o��V]�sI��7�()�g"��#�D�+��;��)N��b�S�s�����?<��h���M���舾�{������􃾭@}�x�m��&[�SG���5��(� �"�]2%��E/�Z?�T�R�C�f��w��V���r��y���)w��4���9
��Dc��:�6v|�{ul�rOY��E��r4���(��+$���'�D3�Q�C���W��.k�C�{��  �  �����������\}�[�n���_��	Q��	B��d2�m�!��O��������ڽ�dֽ�ݽ�F�V��K���b&���6�mF��}U��d���s�G󀾜���ED��X܇�������o�W�U�=���(�s�d���2"��	4���K���e��C|�5��E���ß��;-���5{�\_l��X]�DnN�5?�E7/������ߡ���8�H�۽:۽a*潈������p�b-�5#=�W^L�
<[��2j�;y� A�����wo��灆�1~�$Ih�;O�M7�q�$�
���B�=�)�Ty>�	X�e�q�G���YJ���p���W���#���|��m���^�}P���@���0�um ����io�r��n���^v �C������-���>���N� @^�=]m��|�ڪ����Wя��h�������'gn�,U���>�q4/��)�\�.�hT>�2U�Uo�ă��+��QR���Ⓘ��������Z���u�+�f��X�r�H��^8�`(������~G��j����0�1�_/��@��?Q��a�5Qp�#}��[�����->�����[Ε����>C��%?t�x�[� 3G���:���8��A���S�Y�k��Ⴞ�I��E��ř��ј�Y��k����F���m}��hn��_� O�{:>�Z�-�i��G���d����B�O�+�<�m�L��\�k"l�f{�k������DG�����z��	����������n�tV�|�C�@G:���;�joG��[�¹t��iW���ߗ�Lי�񚗾�M��?X���܃���x���i�}Z�$FJ��9�)�l���E�~�����B�Kr#��2���C�K)T�)d�Z<s�R����������U���*���;��zƕ�l ��A2����h��R�)4B�i.<�t&A��1P���f�e���,���p���  �  �2��!���ޘ����%�|�#J`�u2F�G/�:���	�f�򽙞ؽ4�Ľ�����'���ݺ�Y&ɽ��޽.���؅�� ���4���L�H�g��A��fM��{����	��.���z���E��Dx��rbb��+G��m6��H3��T>�2�U���t�缊�,��������:���b��(��F�u���Y��@��[*���������\<սt�ýT��Շ��#����ҽXJ�߸�&��¹'� �=��FV�!�q�fM����������&��˂��b��}o���^x��$Y�y7A��!5�667�'G��b�[���+ޑ�1�6��&���PU��58���t���Jr�ocW�6h?�5l*��	�P��.���0'߽Pѽ�z˽}Ͻ�g۽����������&��L;�\R�Mal��c���Ò�=����_���^���|��i-���b��j|��^�E~J�  C���I�8�]��!{�TC��!��������魾�ܫ�����ki��{9���v�-\�s!E�Q1�q���*\����;�X���9��Y������"�O�'�b|:�ЯO�&�g��[���ˏ�睾/����ְ�������ì��=!������e�S?U���R���]�cu��O���ܚ����6O���Ǵ�Yo������bL��Lڊ�)�y�р`�->J�;�6�Um%�st��3
�yY�k��|���* ����خ��L#�94��lG�G]��"v�%����N��"ˤ�*'���6������!���e������x��q`�3�S��U�Ze��t�$鏾V���0Ǭ�	ҳ�h��������c��Ɏ���1��aq�eDY�zD�P~1�J!����
��� ������o���{�p*���%�*�S<�wnP��Tg�ݟ��sˎ�o'���᩾c���쪵�^���}K���_��j懾-r���]��U�d\��o�uU���ږ��-���I���  �  Ɍ��j��������^��� kj���E��&��s�3x򽌰ҽ;w��!W��?O������<���$������?ڽW��3{��+.�6�N�q}t�ᎾY/���B������2�����~'������3����d�u�O�~�K��Y��Rv�}z������v����y��U����h��]ӫ�a����ڃ��`��'=�I ��i��K�R�ͽ����"���=���Ǡ�٭��˼����ʽ�2罧�����>69��o[�ON����������Ҹ����������[���ϐ���z���\���M�>!P���c�M�������P��YO��4�þ�¾n�������ɔ�U/���:Z�Oa9��]����+���ս��½�4���ݲ��ﵽ�P����ѽ>@����/��C2�q�P�6>u�B䎾靣��$���\þ�Ⱦ��ľ]&��ť�L`��a'~���d�a[���c��T|�&j��E,��|Y����ž@˾�2Ǿ�躾�𨾻l�������[���<��#�Ũ�} ����z8ؽJϽ-"ͽ}�ҽ�k߽95��	�L���-���H��i�伇�l��eɰ�Q���L�̾�+ϾYKȾ����:3��,��?|��q�n��!k��(y�� ������Z"���ľ#�Ͼ*�Ѿ7�ʾ���¨�`����� &]�a�?�:5(�]\����)��"�F���߽���C�������.�1t%��y<�X�X�+N{��G�����X���Q�Ⱦ��о� о�ƾ7��u������l|�˥l�Ȭn�&ꀾ�Q��|�� y��y/ɾ�OѾj<оdƾV(䡾�<��;t�'AS��8�X;"����������W�N$��U���My��8�ծ�І.��aG���e�����J��� ��4���:�;��Ҿ��ξ�B¾����W6������c�w�n��v�d#��{4��Rɭ�y���Kξ�  �  $�ھ�nվ��ž�7��򁕾�Ex���J��%�-����oH���V��Ga��p������*��r暽jЬ�ǽ�O뽝	���-���U�q@������m��P�ʾ��ؾ7�۾v�Ӿ����X�������[}�n�d��R`��ap��"���蟾�%���̾;�پ��۾ĄҾ�$���������j���?�0����3�ؽq~���3���}��ݖ���.��aA��1���]���qԽJZ������;��,e�����0ꤾ�`���оZ�ھ�=ھ��ξ�����m���.t��6b�ae�d�{���������u����rԾ�޾��ܾ�о�����������
b���9�H^�f� �mܽ�%½�i��0���W���(��X����ƾ�Z�ֽ�0���� �/��1U�o���J��"5��m˾�ܾ� �`�޾n�Ͼ�������3d����z���o�8qy��&�������Ͼ�߾N���4྄�о��[e��_����`�H;�$^�����콚wս�Gƽ�+��T���0����;ͽf�߽1���1��m�(�
�H�fp�Q���A����þ��ؾ=Y�\�����OоU��F���!�Q���������!��� ���OȾsݾK��B��ͼ�sUо76��j4���s��*�_�Xp<�B� �������]a���ֽ[�Ͻ�0Ͻ9Cս��st��5�	����wz8�n�Z���������﴾kn;�����S�}�޾��ʾ���Iq������@����ҁ����_��y*��t�Ͼ]Y����e���fݾ��Ⱦߛ��S˕��|�ߕS��3����j����b��)ֽ�ѽY�ӽ�ܽt��\�����'�AE��$j�,s��_���������վq��I�����پ�ľ�ӫ�����9��{ㅾ�#��
k�������3ؾI��  �  �}�P�"Zվ��������Ձ�0kP�&����v�ؽoM�����|g��_섽縂� ���Ґ��}��SD�����B]�ޡ/�R@\�ë�� ڥ�1�¾��ھԅ�()��zѾ驷����Z���s��n�n�����˫�Ŭƾ�ݾ����z��I�ξ�o������t�n�C��@�����ϽII�����񭍽F-��Dˆ���ݘ���� /˽������XT>���m�ނ���篾��˾�q��=�E��E�߾�hɾ.ʮ��H��Fс���o���r�M#��^�=i��w�о������Q��ɾ�������3ei�<��������ҽpӷ�G��!]����������1���S}����̽>��N�4{0��&Z��_�������W���ھ���~��ܫ�GྡȾ#O���b���ׄ�N[}�O����链7���F�ƾ��߾7���+�����-�E�ƾ�t�������Pf�R<���2�����(˽\Q������QX�����!/ý2�սd.����&�_J�#w��*��oe��1CоM��EV��'��<U�Y�߾�kƾ|%��eV�����ɹ�����P���'绾@�־e��r4���S��\���޾�þu������c��&<�-��������j"ڽ��̽h7ƽ�Ž��˽��׽�3�N.�+��&�7� ^��ن�a~��u��۾���4V��������>pپڿ���$������v����ӈ�5>����9�ľI)߾���8��|��-��L־չ�����˳����U�?�1��i��� ���A׽�̽�CȽ�ʽҽ/'�Ч��bl�qW%�ڔE�Io��ː��]����ʾ��4���/���F���Aa꾁Ҿ=#��4��[�����Q,���霾�r��u`Ͼ�W����  �  $�A��;���+��.�����Ǿ����JFu�	DA�X�m� ��ݽT�ƽ���H~��\弽��˽�I彼l��j#�~bL�����+	��*Ҿ���m��P�0���>���A���9��(��)���kξl%��Zٲ�����U�ᾞ��RW�a�2�+�?���A��68�ʁ%�'u��=�lH��˗���wd�N^5�rx�@���ǮؽwŽ�+��������ý�ս�R����0��^�Ii���%���a⾩o
�s�"��N6�^�@��\@�.�4�e� ��3	�]	�פľٳ�>����˾�d��M�^�&��V9���B��A��B4��]�ʀ�>۾uQ��v����Y��/�v��Ɉ������ҽ��ͽ*'ѽՉݽ�2�����;�%�ɲJ��a}����?�ɾ�����L��-��>��E�$<A��f2����@�����ľ�:��}þ�ݾU���,B1�l<A��G�WRA��W1���T���Ѿ����ġ��mW�_�1� z�/��h���΅꽍B�Z��6���`�y� �&�=�g��r��;���\�߾Ӭ��!�,x7�ŎE�:�H���@��\/�:����h�ݾ�ƾE�¾��Ѿu����f�&�(;��H���I�=j@�į-�x��U}��xɾ\����K�� bU�.c3�������t����U���x��4�
�`d���/�ltP���}�m��q6ľ ��A����*��n>��I���H�G�<���(�HM�I&����Ծ)�þx�ž��ھ�r�����w�-��X@�y�I�Z�G���:��%���8'��a���y����s�!^I��P+����$a	�`��������m���k�H�!��M;��_�7��v����Ӿ��w��2���C�P�J��ZF��v7���!��*
���IIξj�þT<̾
����GO�6}5��bE��  �  ��;�CY6��	'�AI�b�mþ֚��t�m�A������i��˽���ջ��[��^Eн���͍��$�(�L�3%��_ȣ��ξ��������+�_�8�b<��:4�(J#��I���fɾSP���+��ʖ��7bܾ]7�����-��:��;���2�i� ���	�tJ�LF���+���c�e6�[`�����hݽ�ʽd���m���2PȽ�cڽ"���#�M�1�{�]�$���U��_�ݾ���X�=1��6;�n�:�S^/��=����ׇ�KX��(���y����ƾ���i���"�w�3�k%=�Gd;�a/����Q���־!⫾�y����Y��1��
�� ��>�j^׽<ҽ�ս�#�=��� ��'��qK��l|�qE��5'ƾ�f��p����(��
9�t�?���;�I_-������`ܾ���������[
پq$ ����Q,�3�;��BA���;��x,��������Wξǥ����PX�2k3�<��:F����H����j�[o�ѹ�>�"�;Z?��[g�Ԙ��_L��=�۾�������i2���?�H"C�Tb;���*����4��m�ؾ�þ�'����;z���c��*"���5�	JB��"D��	;�I)������uƾXK���
���hV��J5����y��������X�����������1���Q�N�}��'��wf��W��6��s&�D!9�"ZC� �B�߁7�j]$����u��USо����w¾W־����n���/)�a�:���C��B�I�5���!���	���㾉�K}����s���J��e-���*�����+� ��������%�#�/=�n�`�%���h���ɐо������"�-��:>��E�`�@��o2���������5@ʾ\�FȾ⾽���;�:�0���?��  �  ��+�p'�I���������ﹾ�.���r���D���"�\>
�;t��ڽ��̽"lɽ�QϽ��޽c��ע��[*�|�N�O�~�T&��}Sþp������h)�,�(%����y�@ݾL��Uv��⽤�޲��zV;y����p]�L*�y�+�$��s��M ��־���������c��:�������W�'Jؽ�:ν��ͽ.�ֽ[D�6t�A��RP6��A^��E��� ���Ѿ�y��)�w"�V[+���*��� �����K���Ѿ�6��n����ͧ�D���1ھ]����$��--���+��!�����l��v˾����h��x�[��H6�~���]����g�.�߽qR�n�����S��-�{�N�!{�����?��L���=�:��]�)���/��	,�zl�������;�S���9���泾:˾k��_���:,��<1��z,�4$�� ����e�ľ ��s��~[��\9�� �c����p���%(��P} ����J<�F�)���D��ui��猾�����оR����l�>�$��T0��3��>,�%\���	��H쾤�˾)6��2�������F�ݾ�������'�z�2��44��I,�z���t��M澷��� ������Z���;���%���������=�I�
��S��.#���8�)V��/~�I��1���0�����C�d�*��}3���2���(�r�����z&ᾘ)ľ�x��j^��ޑɾ�1龞Y��6��+�94�er2�c�'�H&��G�q�ؾ�Ͳ��k���gu�)�O�	^4�g� �T���
�څ������[K��@+�O9C�)d������ɩǾ�A��p��� �~/���4�#)1��}$�E���]��vw׾�׾�����D��(8Ծ�9�������"��^0��  �  �O�W���;��q��ξ�[�� ����t���M���/�`x�/���5����{὏,����!�
����g�6��V��~��F������[׾�e��fy
����<��O�������epľ����'Q���/����AL��l�־���m�
����1��7���:������ľ��Ks��e�h��@E�)~)�������C��}潨�彣�｝;����&��nA���c�.x��W`���}�Pa��6����^���|���+[ھ�t��SG������ꗾB~���M¾���1{���;��Q��]o�Z��1j޾�+�����ƅ���b�:B�H
)������Lm��2�������=����ّ#�?�:��zX�R�}�>W������N�Ҿ�����	����yP����b���e��f�־�踾g��Nǜ��H��?춾jԾ�]��\��\���������RX���پ�F��e�������d��AF�@+/����ܐ��
�`	�F�����P$���7�
Q��0q�Xь��ɥ�0�þ��R��T������Ⱦ��f
�-�����Ӿ9p��l������,��`�ǾO��s����4�X��7���g�����:.վ����ꑚ��Z���Be�igI�p�3�Y�#��������k����!��m1�UHF�jFa�'ف��z�������Ѿ���{	��T��;���&�j�~�>~ʾ�-���ѥ��k�������=Ѿ�5�B�	���_}�{����E�M��vEʾ�,���ɒ�s|���[��`B��.�c| �D^��������,(���9��`P��m�S����̠�����x2ݾ�������?��3{�Y�����3����¾�ꭾ����p���俾Y2ݾ+����;��~��  �  �l��|�����1.Ӿ�1���ǥ�����"��8�a�'xG��]0�����5��.�B������T��[!�6�5���M��5i��O��^t���>��t¾��ؾa:�h;��>���L���۾-9¾2���j���/��6����a���������Ѿ��������"�|���̾����F�������M�w���Z��A��z+�Mk�j_�JZ�e���/�����)�͓>��W�rt��j��e]���Ჾ��ɾ��߾�;�������� ��©Ӿ�[���I��.5���������*���f���U���L۾�b�����!
���H�d�޾�4Ⱦ�]��gf��Z����t��Y�Q%A���,����A�J���-�B���'��T;���R��m�ͨ��������LL���mؾ�c��J��D� �?h��@��b~Ҿ��������l���h��ڣ��)C������>MѾLJ�x��B��) ��y��޾�Ǿɲ��f���F!��Mx��]��G�:4���%�����3���*���:���O��(h�ak��������̸�q�Ͼ�~澊�����������T�dѾ�-���ˡ�Xє������g���譾��ƾgi�,������;���������(ݾ+�ž�"��[ɜ�����z��ga�[NK��.9��,��	%��$���*��:7�S�H��X^��aw� ����k��Gk��/�¾�ھ�!�A� �����&��0���sɾME������9��
���Q���!���=�Ͼׄ�M����m��y���t��Xվ�w��@v������2����r�xvZ���E�7M5��@*��}%��m'���/�06>��JQ�*(h�,4��3���|���i��9�˾��F���wV�������?���S�ܾ�����O�������uǘ��5���R��Y�پ��7[��  �  o̾Q̾�Pƾ�W����������љ�����n����[m��kT�5=��`*��a����I� ��Y.��B�<}Z��s�V��u����ߜ�TI��;������
�Ⱦ~�;�̾�¾���h����ǋ�L�v���b�_�	El�������iڪ�߻��$ɾKEξu2̾ޒľ�̹�����z��C���싾Q���g��dN�'B8�U_'�����r�N�%�K�5���K�5d�k�|�@h�������蠾�a��"���þu/˾S�;Ҽɾ%���Ҭ�p���=���Ho���`��2c�C/v��3����q3���þO4ξ�
Ѿ;�0ľ���#?��R塾ɖ��h����~�"(f�TlN�^7:��,��&�8&)���4�ܗG��^��]x�����P���!
���c��x����¾�,;��Ӿ5Ծ��;M$��l����������w��n�E�v�fH��B옾/1��.j��YϾ��־g+׾U5Ѿ�@Ǿ"���� ��ä�"����
��|����k�!AT�H�A��;6�<33��;9���G�r\�*ut�w���
Y������^��.ֵ�����2;,�־�۾�ھ��оH���tC���Ϛ�#���9���X�~����!��	��)���;<�پ�޾_�ܾ��Ծ�ʾ�D��򦲾�_��n����������7n��X��G�1�=��=�)�E�A�U� ?k�U䁾5b��t\��]���6����z��*FȾ�EӾSd۾o6޾b�پLTξ��d먾�핾�h�� �������*�����������\����Ѿ9�۾)x޾fQھ�bѾ[ƾ%X����ȣ�7Q��39���p�\g���R��?D��=��h@�©K�e�]���t������h���4��J����е�����>;�׾q7޾�޾qؾ{Mʾ�������������`��U���J���`4���������H�ȾvQ׾�  �  '槾�:������Ȇ������5����4��z§����V瑾�����h��N�0U>�=�9��7A��T�-�n�2���X��0g���ǩ�*���⪰�[O���6���0���?��i6��j���7��a ��m�d���L���=�>;�C�D��^Y�Ru��։�Z+��N���T^�����-_���ױ�����[T���쬾bB���ϛ�M#��4�}���`�J�=�z_<���G� �]�"6z��V���>�����<���Ư��2��P|��.��\���Ȣ���^��\��6^���jx��x\��sG�E�<���>�f�L�v�d��S���ؐ�I����-���ۯ�GH�� ���%派�v��n���7c������}���ڌ���{���`��EM�%�D���H�p�X�T�q��釾3���t���:���7���!��r+���L��z������֯��q=��	-��o����Y}��Zc���Q��K��$Q�=�b���|������Ӝ��������r�������o��@u��B����%�������������rW�����8f��(V���Q�x�Y�I+m�n5��-����w�� ���,�����5���徾{ھ�!罾~���0��X���ܣ���Џ��X��J(k���\�ǨZ�^�d��|y��������؀������������������¾����=��:���N���ͫ�����Ў�	M����i���\�I	\���g��s}�����U7���'�����l���п�I��}���kA������7ջ�8��������s���2��1|�?�f���[��]]�!�j�s��乏�y�v��� Ƕ��E��������+¾	�������^���z��ݧ�by��CB���/y�Ece�'y\��
`��vo��	��U풾5��3"��Yɸ�P�������u�¾��¾�¾V뿾���u����W����������\�v���d�A�]�pXc��t�k)���A���+��Wű��  �  R����A����]��������ƾ �̾̾�ľ�T���2��0>��[<z���c�3]���g�娀��ǒ����w����ƾa;;q̾S�žJ4������L裾�����m�����%�j�ֽQ�;��0)����W���#�ߘ2��G���_�C�x�������IK��5������������ʾ\oξj˾\���GT���w�����"s�Yya��|`�Dp�h���,�����/���dʾ�4ξL ˾�¾偷������/��&���_���'K{��rb��9J��5�T�%�<?�e��Y/*��<���R��cl��삾��&�������W�������CȾ.�Ͼd�Ѿ�&̾Ԍ��㦭�ෙ��r��uRt���h���m�����sx��6����7����ɾ��Ҿ�fԾ�XϾt�ž_l��0����h��%F��!ˌ�5���u�h�NVQ�(�=�h1�B�,�1��
>���Q���i�7�������"˙� ������#G��L�Ǿj�Ѿ��׾�׾�3Ͼ���3���/ę�1ӈ��{��du�I"��L)���{���س���ƾn5Ծ@�ھ��پ\ Ӿ�Ⱦ�$������~���c��Џ�����o���X���G�kV=��;�@C�ÛR���g�,��ʌ���n��'������V�ƾ�Ҿ��ھ�޾�t۾��о�E���_���显�`��������^����ϖ�>���[󽾞Ͼ'VھJ1޾c۾��Ҿ��Ǿ(׻�F[���)��oÙ����C���j�U�T���D�I=��">�cH�6GY�+�o�~?��.���ߝ�������9���׾���ʾ6Wվ��ܾp�޾;پ�I̾�=���#��o����4��d�������������s���?ž?�Ծ�uݾ<�޾��پ�Kо��ľ���g̭�`���	��Hኾ�|�	e��WQ��D�?�=8C���O��c���z�.܉�
0���  �  ɀ�����ݦ��q���tԾJ��[-�������g��޾�ž����-۔����.���E����������q#̾4&�����'O�������E�*о���G���FA��X|���^���D�7<.����D��i���-��k	������%���:�;KS��Ko�Ѷ���G��{w���pƾ|�ܾBNﾮ����@��eX�,ؾ���T��͏��6��͑������c��� ��QIվ6�ID���������޾l�Ⱦ����[*��ST��[r�u�U��1=��
(��Qd�����6��#�I���/���F���`�,�~��^���������j9Ѿ��澃���-��i���g��Z�Ӿ�2���堾�<��qf���Ê��˘������ɾ�@������@ ������%��޾��Ǿ�����������hv�I�[��#D�(e0�;(!�.��vG�}���!�CK1�qE�95]��Nx�X����_���ű��[ȾY^߾��+� �cH��}���*�WѾ`��.���[葾Ͼ���є�F����*��,�ؾj-�;� ����B� �M���ݾ��ƾ�����������z�Dxa��iK��59���+��T$�	X#�|�(�h�4���E��*[�q�s��������A����Ŀ�f�־2�Wu��������T��T���;�3��Ԧ������e���͝�x��T�ʾ6(�u�������jT ����v�ؾ�����Q��y{��R0��
v�n1]���G�x�6�n�*���$�6m%���,��4:���L���b�Qy|��⌾�����9���-ǾBU޾���	�����d�|s��aྺ�žq��FE���>���j���@���W��n�Ծ� �� �Q�����������辐,Ҿ@����즾:����{����o��7X��%D�F�4�
*�\�&���)�>k3��B�:bV���m�YT���  �  ��u����D����о@K�?��2��i����4�˫�ɾ�@���������
�������о�m�p����������W���뾿�ɾ�����,��|n���I�*�,�b��]���󽚾潮v佄��H�����;�"�۝<��]�彃��r���һ��=ݾ��������I�M��� �1X�����K	��^;���T���3��itܾx���X��>��b	���ߛ ���ྦྷ���F�����sa�(�?��.%�m�������轭[� e��,��Q��x�.���K� �o�������9�ɾ'��n�����u��v���R���پ@%���ţ�{ٙ���������˾Et�(�DN����f��R5�����2ܾ�D���띾@g��GYc�fBD��,����Ŵ�1��qf��I�������a�-�q�E��d��Ņ�}Ꝿ&Ế��۾!5���y����Y���M���
�y	����Ծ*����i������慨V���q)ݾT9������=��D�pu����:��g�׾`�������,��Ef�1�I�c�3�5#�o��L���L������S�.��C�1]�mX~� ���í��̾8~�K)����	���M�������>�xϾDx���ަ����C(���̾M�A�����M�������1����\8Ͼuj��p0��Հ�ȶ_�pE�4�0��`!��[�<���F��D�c�$���4�5�J�fg��s���盾pA���־����%'�1��������b����l�VƾHʯ�F�������P��i׾����s�����5����m�����׬ž�O��������w���X�i2@�&�-�� ����P��Ih�3�j8,��p>�$QV���t��  �  :~t�*ї�����Y:�"����g�'�3�+��&������6��@P���	������Fʭ��>Ǿ����+
�B��O�(� ,��%�C4�)���ܾ�F������$k�w�?����Y@�.����ٽXνN\̽��ӽc�~ �ַ�.�0�yW�娄�pv��Гʾ����*��k �#�*�{�+�qD#�Z/�Et��L8׾�;��H榾��˄��_-Ӿ��������!��4+��;+���!�M,�.���ξ������5�[��S4��i�r����9�׽;н�9ҽ��ݽl��L
��x!�A6A�ák��L��!u���d۾�
�`�pl&���-���+��m �~�������ϾU4���^��-A��S(þɿ�Ȉ�����(��z/��T,�!A �����9/Ⱦ�l��Z7���C[���7�E��r��1���~��r�����fe �����V���8���[��������)�ƾm%�;M�g$ �"%-�b{1�[,�B��8��C�`̾:絾񐯾����Ӿ�;��֋���"�^U/�ʽ2�wm,�N��tU
�B)�����w[���|���\��?<��M%��N�b�
�-���,��N	�KK�� �65�wVQ�עw������Ĵ���ھ�~��C�v}(���2���3��A+��&�'-����Ⱦw����ŵ��Wž�c�������)��*3�#73���)��2�.��b�޾g7�������{��aT�uI7��Y"�����
�������q����}�&�L]=���\��T��"���N������	�k��/�,��R4�C2���&����H� �Sܾ�5���5��^칾V�ξa�H�!��
C.�F�4�%�1�z%��'�H ��~�Ҿ�Э�-��� �o��(L��2��t�0���v����c�E�P7�y<0�V�I�=4l��  �  K�v�������ž/���m��Y&(��7��<�v�5�w=&����S\���;�$���歾�O���վ�S��E��"�*��f8�d<���4��$�����꾴㼾�����l��D<��e��� �چ�o{˽(�������(�ŽGֽ�����I�+���U�솾8ު�O6־�%�	����.��z:��;��#2�" ��	��c�j�ľ�����}������%������9f0�&;�};��D0�&6����3۾���F?��'�Z�w�/����s���VGڽ��ɽ��½�Ľ��Ͻ������N6=���k�tє����e�����O�#�;G5��=�4v;���.�T�����޾����"Ƴ�%.���lо����Pz��r'�f8� ?��;�s�-��	��� ���ҾsΨ�߸���X�?92�k���-�T��㽙3߽���B�Co�c ��)3�IY��9��˘��ӱо��������-���<�0�A�Jt;���+�,s������پ� ���빾�~ž��:n�:N��1���>�ʹB��r;���*��p�Q]����ʾlN�������mX���5�8��:�����N���s����:�w�
�V�H.�3IL��Bv��8��#+���}澎D�r�"���6���B���C�� :���'�Ǔ�)B��.�Ծ�a���P��l�Ѿ���f��t�%�X8�1C�l	C�E8��;%�u��.�c'��t[����z�N�O��0�����h�C��0}���E ��J�}O��I�B�6�0�X������)���Ⱦ���[�f9*���;��GD���A��5��� ��:
�p���̾ۜ����ľl�۾� ��	���,�!y=�]�D�HA��33��?��*���ܾ�2������ym�~�F���*����e��N���!�"(���
���T)��C��ei��  �  vx� ����ɾ9���ȑ��-�X�<���A�zv;� #+�B��h�����ҾI������:c����ھD�<,���/��>���A��@:���(�[g��+3���0����l��r;�p���B��Q�۽��ƽ�2��+g���;���ѽ�I�H���*�ʸU�(���1e��R�ھ�c��0���3�4@�B�A���7���$�FZ�Q'�kQɾ�N��Y6��d0ƾ�{�w�
��"��5���@� �@�ʈ5���!��	�I�߾�����r����Z�o.������Q�ս	Ž,E���G��]+˽+�Ǧ ��1��B<���l��Q��v���=�Wn��X(�[�:���C��)A���3���Ё�}	�J$žxq��,
���"վn���Zf��@,�a�=��OE�8wA�3�2������C�־n���ꁇ�b�X�w�0�װ�F�������޽r�ڽ�߽&��;�y���1��X��↾~���klԾq���1�2�HB��UG�~A���0��y����޾��ľ������ɾ9#�A��ǆ ��6�ʖD���H���@�̏/�Y(�֨��E�;����a��=�W�(4�գ�/d�o�6&��/E��������Ũ�k,���J� Cv�6F������c��u��)I'���;��=H��I�d�?��,�M����*پ�#žF	ľ!־DP��P��U*��=�z�H���H��=��)�/���ﾷ���	����#{�wsN��.����
��c��!��V*����.��F�-5�x�W��σ�v�����˾�(�����1�.��'A�|J���G�s,:�AM%�����/��"ѾHþ��ȾX��O��W��+�1���B�;�J���F��68��Q"��+	���ྮ\���ۑ��m��	E�(�(����4	�kF�y�������y�"T���&�dB���h��  �  K�v�������ž/���m��Y&(��7��<�v�5�w=&����S\���;�$���歾�O���վ�S��E��"�*��f8�d<���4��$�����꾴㼾�����l��D<��e��� �چ�o{˽(�������(�ŽGֽ�����I�+���U�솾8ު�O6־�%�	����.��z:��;��#2�" ��	��c�j�ľ�����}������%������9f0�&;�};��D0�&6����3۾���F?��'�Z�w�/����r���TGڽ��ɽ��½ �Ľ��Ͻ�������K6=���k�rє����b�����M�#�:G5��=�3v;���.�S�����޾����"Ƴ�&.���lо����Qz��r'�g8�?��;�t�-��	��� ��ҾvΨ�Ḇ��X�B92�m���-�T��㽙3߽���B�Ao�a ��)3�EY��9��ɘ��ѱо��������-���<�/�A�It;���+�+s������پ� ���빾�~ž��;n�;N��1���>�˹B��r;���*��p�S]����ʾnN�������mX���5�;��<�����Q���u����:�x�
�V�I.�3IL��Bv��8��#+���}澎D�r�"���6���B���C�� :���'�Ǔ�)B��.�Ծ�a���P��l�Ѿ���f��t�%�X8�1C�l	C�E8��;%�u��.�c'��t[����z�N�O��0�����h�C��0}���E ��J�}O��I�B�6�0�X������)���Ⱦ���[�f9*���;��GD���A��5��� ��:
�p���̾ۜ����ľl�۾� ��	���,�!y=�]�D�HA��33��?��*���ܾ�2������ym�~�F���*����e��N���!�"(���
���T)��C��ei��  �  :~t�*ї�����Y:�"����g�'�3�+��&������6��@P���	������Fʭ��>Ǿ����+
�B��O�(� ,��%�C4�)���ܾ�F������$k�w�?����Y@�.����ٽXνN\̽��ӽc�~ �ַ�.�0�yW�娄�pv��Гʾ����*��k �#�*�{�+�qD#�Z/�Et��L8׾�;��H榾��˄��_-Ӿ��������!��4+��;+���!�M,�.���ξ������5�[��S4��i�q����6�׽7н�9ҽ�ݽd��L
��x!�:6A���k��L��u���d۾�
�]�ml&���-���+��m �}��
�����ϾU4���^��.A��T(þʿ�Ɉ�����(��z/��T,�$A �����>/Ⱦ�l��_7���C[���7�J��v��6������r�콾��de �����V���8���[��������$�ƾh%�8M�d$ �%-�_{1�Y,�B��8��C�^̾9絾񐯾����Ӿ�;��׋���"�`U/�ͽ2�ym,�Q��vU
�G)�����{[���|���\�@<��M%��N�e�
�0���,��N	�LK�� �75�xVQ�עw������Ĵ���ھ�~��C�v}(���2���3��A+��&�'-����Ⱦw����ŵ��Wž�c�������)��*3�#73���)��2�.��b�޾g7�������{��aT�uI7��Y"�����
�������q����}�&�L]=���\��T��"���N������	�k��/�,��R4�C2���&����H� �Sܾ�5���5��^칾V�ξa�H�!��
C.�F�4�%�1�z%��'�H ��~�Ҿ�Э�-��� �o��(L��2��t�0���v����c�E�P7�y<0�V�I�=4l��  �  ��u����D����о@K�?��2��i����4�˫�ɾ�@���������
�������о�m�p����������W���뾿�ɾ�����,��|n���I�*�,�b��]���󽚾潮v佄��H�����;�"�۝<��]�彃��r���һ��=ݾ��������I�M��� �1X�����K	��^;���T���3��itܾx���X��>��b	���ߛ ���ྦྷ���F�����sa�(�?��.%�l�������轥[�e��&��J��o�.���K��o�鉎���2�ɾ ��j�����u��v���N���پ>%���ţ�{ٙ����	�����˾Ht�*�GN����i��U5�����!2ܾ�D���띾Fg��RYc�nBD��,����ɴ�3��qf��I�������Z�-�i�E�ۘd��Ņ�vꝾẾ��۾5���y�}��V���M���
�u	����Ծ)����i������慨X���t)ݾX9������=��D�su����:��n�׾g�������,��Of�:�I�k�3�5#�t��P���L������T�.��C�1]�mX~� ���í��̾7~�K)����	���M�������>�xϾDx���ަ����C(���̾M�A�����M�������1����\8Ͼuj��p0��Հ�ȶ_�pE�4�0��`!��[�<���F��D�c�$���4�5�J�fg��s���盾pA���־����%'�1��������b����l�VƾHʯ�F�������P��i׾����s�����5����m�����׬ž�O��������w���X�i2@�&�-�� ����P��Ih�3�j8,��p>�$QV���t��  �  ɀ�����ݦ��q���tԾJ��[-�������g��޾�ž����-۔����.���E����������q#̾4&�����'O�������E�*о���G���FA��X|���^���D�7<.����D��i���-��k	������%���:�;KS��Ko�Ѷ���G��{w���pƾ|�ܾBNﾮ����@��eX�,ؾ���T��͏��6��͑������c��� ��QIվ6�ID���������޾l�Ⱦ����[*��ST��[r�u�U��1=��
(��Nd�����6��#�B���/���F���`��~��^���������a9Ѿ���{��-��b���b��U�Ӿ�2���堾�<��qf���Ê��˘� ���ɾ�@������@ ������%��޾�Ǿ�����������hv�T�[��#D�.e0�?(!�0��vG�{���!�=K1�qE�/5]��Nx�Q����_���ű��[ȾP^߾��&� �_H��}���*��VѾ]��,���Z葾Ͼ���є�H����*��0�ؾp-�?� ����F� �V���ݾ��ƾ�����������z�Oxa��iK��59���+��T$�X#��(�j�4���E��*[�r�s��������A����Ŀ�f�־2�Wu��������T��T���;�3��Ԧ������e���͝�x��T�ʾ6(�u�������jT ����v�ؾ�����Q��y{��R0��
v�n1]���G�x�6�n�*���$�6m%���,��4:���L���b�Qy|��⌾�����9���-ǾBU޾���	�����d�|s��aྺ�žq��FE���>���j���@���W��n�Ծ� �� �Q�����������辐,Ҿ@����즾:����{����o��7X��%D�F�4�
*�\�&���)�>k3��B�:bV���m�YT���  �  R����A����]��������ƾ �̾̾�ľ�T���2��0>��[<z���c�3]���g�娀��ǒ����w����ƾa;;q̾S�žJ4������L裾�����m�����%�j�ֽQ�;��0)����W���#�ߘ2��G���_�C�x�������IK��5������������ʾ\oξj˾\���GT���w�����"s�Yya��|`�Dp�h���,�����/���dʾ�4ξL ˾�¾偷������/��&���_���&K{��rb��9J��5�Q�%�8?�`��R/*��<���R��cl��삾	���������M������}CȾ%�Ͼ\�Ѿ�&̾͌��ަ��ܷ���r��rRt���h���m�����vx��;���8����ɾ��Ҿ�fԾ�XϾ}�žil��:����h��-F��(ˌ�;����h�VVQ�-�=�k1�C�,�
1��
>���Q�~�i�1�������˙� ��󃰾G��B�Ǿ`�Ѿ��׾�׾�3Ͼ���.���+ę�/ӈ��{��du�J"��N)���{���س���ƾv5ԾH�ھ��پe Ӿ"�Ⱦ�$�� ����~���c��Џ������o���X���G�pV=��;�@C�śR���g�,��ʌ���n��'������U�ƾ�Ҿ��ھ�޾�t۾��о�E���_���显�`��������^����ϖ�>���[󽾞Ͼ'VھJ1޾c۾��Ҿ��Ǿ(׻�F[���)��oÙ����C���j�U�T���D�I=��">�cH�6GY�+�o�~?��.���ߝ�������9���׾���ʾ6Wվ��ܾp�޾;پ�I̾�=���#��o����4��d�������������s���?ž?�Ծ�uݾ<�޾��پ�Kо��ľ���g̭�`���	��Hኾ�|�	e��WQ��D�?�=8C���O��c���z�.܉�
0���  �  '槾�:������Ȇ������5����4��z§����V瑾�����h��N�0U>�=�9��7A��T�-�n�2���X��0g���ǩ�*���⪰�[O���6���0���?��i6��j���7��a ��m�d���L���=�>;�C�D��^Y�Ru��։�Z+��N���T^�����-_���ױ�����[T���쬾bB���ϛ�M#��4�}���`�J�=�z_<���G� �]�"6z��V���>�����<���Ư��2��P|��.��\���Ȣ���^��\��6^���jx��x\��sG�@�<���>�_�L�m�d�S���ؐ�B����-���ۯ�=H������派�v��e���.c��햦�w���ڌ���{���`��EM�$�D���H�t�X�[�q��釾$3���t���:���7���!��|+���L���������߯��y=��-��t����Y}��Zc���Q��K��$Q�8�b���|������Ӝ�����򰲾i�������o��6u��8����%����������}��mW�����8f��(V���Q�{�Y�N+m�r5��2����w�����%,�����"5���徾�ھ�+罾����0��`���⣞��Џ�Y��Q(k���\�̨Z�b�d��|y��������ـ������������������¾����=��:���N���ͫ�����Ў�	M����i���\�I	\���g��s}�����U7���'�����l���п�I��}���kA������7ջ�8��������s���2��1|�?�f���[��]]�!�j�s��乏�y�v��� Ƕ��E��������+¾	�������^���z��ݧ�by��CB���/y�Ece�'y\��
`��vo��	��U풾5��3"��Yɸ�P�������u�¾��¾�¾V뿾���u����W����������\�v���d�A�]�pXc��t�k)���A���+��Wű��  �  o̾Q̾�Pƾ�W����������љ�����n����[m��kT�5=��`*��a����I� ��Y.��B�<}Z��s�V��u����ߜ�TI��;������
�Ⱦ~�;�̾�¾���h����ǋ�L�v���b�_�	El�������iڪ�߻��$ɾKEξu2̾ޒľ�̹�����z��C���싾Q���g��dN�'B8�U_'�����r�N�%�L�5���K�5d�k�|�@h�������蠾�a��"���þu/˾S�;Ѽɾ%���Ҭ�o���<���Ho���`��2c�=/v��3����j3���þG4ξ�
Ѿ;�0ľ���?��J塾ɖ��h����~�(f�LlN�Y7:��,��&�:&)���4��G�#�^��]x�����W���)
���c�������¾�,;��Ӿ>Ծ��;T$��q���񸙾�����w��n�C�v�dH��>옾*1��(j��RϾ��־^+׾K5Ѿ~@Ǿ���� ��ä�����
��v����k�AT�C�A��;6�<33��;9���G�y\�3ut�}���Y������^��7ֵ�����2;6�־�۾�ھ��оN���yC���Ϛ�&���;���]�~����!��
��)���;<�پ�޾_�ܾ��Ծ�ʾ�D��򦲾�_��m����������7n��X��G�1�=��=�)�E�A�U� ?k�U䁾5b��t\��]���6����z��*FȾ�EӾSd۾o6޾b�پLTξ��d먾�핾�h�� �������*�����������\����Ѿ9�۾)x޾fQھ�bѾ[ƾ%X����ȣ�7Q��39���p�\g���R��?D��=��h@�©K�e�]���t������h���4��J����е�����>;�׾q7޾�޾qؾ{Mʾ�������������`��U���J���`4���������H�ȾvQ׾�  �  �l��|�����1.Ӿ�1���ǥ�����"��8�a�'xG��]0�����5��.�B������T��[!�6�5���M��5i��O��^t���>��t¾��ؾa:�h;��>���L���۾-9¾2���j���/��6����a���������Ѿ��������"�|���̾����F�������M�w���Z��A��z+�Mk�j_�JZ�e���/�����)�͓>��W�rt��j��e]���Ჾ��ɾ��߾�;�������� ��©Ӿ�[���I��-5���������'���b���P���L۾�b�����
���H�[�޾4Ⱦ�]��_f��S����t��Y�I%A���,����>�J���-�F���'��T;���R��m�Ԩ��������UL���mؾ�c��J��H� �Fh��F��g~Ҿ��������l���h��٣��&C������:MѾFJ�x��>��) ��y��޾�Ǿ����^���?!��Ax��]��G�44��%�����5���*���:���O��(h�gr�������̸�z�Ͼ�~澓����������$T�iѾ�-���ˡ�[є������g���譾��ƾhi�-������;���������(ݾ+�ž�"��[ɜ�����z��ga�[NK��.9��,��	%��$���*��:7�S�H��X^��aw� ����k��Gk��/�¾�ھ�!�A� �����&��0���sɾME������9��
���Q���!���=�Ͼׄ�M����m��y���t��Xվ�w��@v������2����r�xvZ���E�7M5��@*��}%��m'���/�06>��JQ�*(h�,4��3���|���i��9�˾��F���wV�������?���S�ܾ�����O�������uǘ��5���R��Y�پ��7[��  �  �O�W���;��q��ξ�[�� ����t���M���/�`x�/���5����{὏,����!�
����g�6��V��~��F������[׾�e��fy
����<��O�������epľ����'Q���/����AL��l�־���m�
����1��7���:������ľ��Ks��e�h��@E�)~)�������C��}潨�彣�｝;����&��nA���c�.x��W`���}�Pa��6����^���|���*[ھ�t��RG������ꗾ@~���M¾���/{�߻�7��N��Zo�Z��*j޾�+�����ƅ���b��9B�A
)�������Hm��1��������=����ߑ#�G�:��zX�]�}�DW������U�Ҿ#�����	����|P����d���e��i�־�踾g��Nǜ��H��>춾jԾ�]��Z��\���������JX���پ�F��_�������d��AF�9+/����ؐ��
�`	�G�����P$���7�Q��0q�^ь��ɥ�7�þ��U��T������ʾ��f
�1�����Ӿ<p��n������,��a�ǾO��s����4�X��7���g�����:.վ����ꑚ��Z���Be�igI�p�3�Y�#��������k����!��m1�UHF�jFa�'ف��z�������Ѿ���{	��T��;���&�j�~�>~ʾ�-���ѥ��k�������=Ѿ�5�B�	���_}�{����E�M��vEʾ�,���ɒ�s|���[��`B��.�c| �D^��������,(���9��`P��m�S����̠�����x2ݾ�������?��3{�Y�����3����¾�ꭾ����p���俾Y2ݾ+����;��~��  �  ��+�p'�I���������ﹾ�.���r���D���"�\>
�;t��ڽ��̽"lɽ�QϽ��޽c��ע��[*�|�N�O�~�T&��}Sþp������h)�,�(%����y�@ݾL��Uv��⽤�޲��zV;y����p]�L*�y�+�$��s��M ��־���������c��:�������W�'Jؽ�:ν��ͽ.�ֽ[D�6t�A��RP6��A^��E��� ���Ѿ�y��)�w"�V[+���*��� �����K���Ѿ�6��m����ͧ�D���1ھ[����$��--���+��!�����l���u˾����h��q�[��H6�y�	��X����g�.�߽rR�r�����S��-���N�#!{�����?��Q���=�=��`�)���/��	,�|l�������;�S���9���泾:˾k��]���:,��<1��z,�2$�� ����`�ľ ��o��w[��\9�� �`����n���%(��Q} ����M<�J�)���D��ui��猾�����оW����l�A�$��T0��3��>,�'\���	��H쾦�˾*6��3�������G�ݾ�������'�z�2��44��I,�z���t��M澷��� ������Z���;���%���������=�I�
��S��.#���8�)V��/~�I��1���0�����C�d�*��}3���2���(�r�����z&ᾘ)ľ�x��j^��ޑɾ�1龞Y��6��+�94�er2�c�'�H&��G�q�ؾ�Ͳ��k���gu�)�O�	^4�g� �T���
�څ������[K��@+�O9C�)d������ɩǾ�A��p��� �~/���4�#)1��}$�E���]��vw׾�׾�����D��(8Ծ�9�������"��^0��  �  ��;�CY6��	'�AI�b�mþ֚��t�m�A������i��˽���ջ��[��^Eн���͍��$�(�L�3%��_ȣ��ξ��������+�_�8�b<��:4�(J#��I���fɾSP���+��ʖ��7bܾ]7�����-��:��;���2�i� ���	�tJ�LF���+���c�e6�[`�����hݽ�ʽd���m���2PȽ�cڽ"���#�M�1�{�]�$���U��_�ݾ���X�=1��6;�n�:�S^/��=����ׇ�KX��(���y����ƾ��i���"�v�3�j%=�Ed;�`/����Q���־⫾�y����Y��1��
�� ��>�h^׽<ҽ��ս�#�@��� ��'��qK��l|�tE��7'ƾ�f��r����(��
9�u�?���;�J_-������`ܾ���������Z
پp$ �~���Q,�2�;��BA���;��x,��������Wξǥ����LX�/k3�9��9F����G����k�\o�ҹ�A�"�>Z?��[g�֘��aL��@�۾�������i2���?�J"C�Ub;��*�	���4��n�ؾ�þ�'����;z���c��*"���5�	JB��"D��	;�I)������uƾXK���
���hV��J5����y��������X�����������1���Q�N�}��'��wf��W��6��s&�D!9�"ZC� �B�߁7�j]$����u��USо����w¾W־����n���/)�a�:���C��B�I�5���!���	���㾉�K}����s���J��e-���*�����+� ��������%�#�/=�n�`�%���h���ɐо������"�-��:>��E�`�@��o2���������5@ʾ\�FȾ⾽���;�:�0���?��  �  dF��y��&��&c��8�wr���L���3B�� �U�1�/��.��;��H�������F���c	��X��M7��`�H4��������P��|B�O�l����[���B���򐿿o��_e[�GV4����h�b���q	�].%���I�9�q��슿�J��U��Ț��ގ~���U�0�+�t3���ξ�����!z��>I���'�����h��������?����|�$�@vD��Ms�욾n�Ⱦ�8�w'�9�P��y������i���ؖ�.r���v���M�2�(��4�g��%a����V�0��W����%��1�����X���V�r���H�&! �g������ ����n�}�C��'���;H
��u�"��*�k� ���9��o^�����H3�����8��8��Cb� ���듿�5��=�������l�U�D�'("���
��d��v	��S�
�@�d�h�1����ʕ�z����֕��ˇ���h��G>����N��o����R����k��2F��@-�e��M��{������"�175���Q��p{�)���žGA���� ��LI��s�;r���Ҙ��ɛ�Ѝ��"����b�O<����Bt
�d��@��r-���Q��Az�k��rs���*��W����h����]�'�3�[��߾�ϯ��+���Xi�5�G���1�AK$����"]�f#���/��|D��kd�����P�����ؾ�O
��1/�8�X����@��L�����������J~� V���0�iU����tT	�	e��~8��	_��u����������P���ꎿ!�y���O�V�&�|C�	�;a$��B��[]��8@��l-���"�`8�>����'�y#7��lO���s�~��������l��A=��xg�E���Q���=͜�DΘ�����ɦq��I�O�&���_�c�J�#�fE�ALm��ډ��ۗ��  �  ����2���π��c\��4�^s��pݾ����H�����W�"�2��y�eu	�� �����nA����;���<:���b�~A��(����X���R=�Q�e�B����U��S��H"��Z�z�q�T�}{/��o�����T��Q���� �N�C�|j�?d���:���ޒ�+݊��v��O���'����|y̾���f{�}�K��+�� ������ �]� ��h����'�(G���t������lƾh����##�$�J�	Dr��N���J������Dև��in�+�G�C$���	�||�������(,�KQ�$�w�ee���y���⑿h���k���C����`�����
��"�p���F��Y*����Bj�Ҁ	�?��[_�Q$��<�,�`�RL��yN���޾�e���3���[��ဿ�����9B��}�����e��@?��.�����P���v��{�e�;��b��u��ݐ�̕�fꐿ�����a���9�����_��������<"n��@I�'�0��� � �����0�K&�F|8�g�T�Cg}������þf�������"D�
el�����͓�Ƞ������6���}\�O<7��X����WM�5�3)�I&L���r������c�������$�~���W���/�,��7�ܾ�C��΍�,�k�9K�{5��x'�K� ��j �?&���2���G�Og��f��֚��ދ־c���B+��R�(rz��h��bg���ޕ����v�EP�p,������W{����9�3��X��~�V쎿Gꖿ�A���f��6r�*J�e'#��@�(+̾V���)���7`��{C��0�]�%��C!��#�'+�o:�i�R��Vv��锾и��)��@�8�a��|�����e����ӓ��H��]�j��*D�'#�L���U������s5@��mf�����풿�  �  ���G̀�U�j��TJ�b_'�8��ٳվ*���7{��U�_�7�<� $�����a
���������-))��"D�GFj��z��c���ᾦ���r/�YSR�Hq�V���7	����}�}d�c�B��!�^O����� �����O�3���U���s��h��݄��{��a�P?��������ƾ���G�����T�cm5�������
��
��M��p��F2��}P�b�z�������������Q';�3M]�\9y�PY���ك��lv�s]Y��7�d�۞ ����`�F���k�?�S�a�G�|�is��C���u�V�W��5��5�t9뾮u���▾��w��tP���4��H"��3�,��_��n��.�)�F��Vi������謾�׾��nc'�2WJ��*k�Sρ�����n�����q��R�GX0���g���R����e��G_-��&O�go�$e������4�����o���O���,���������e���&Yv�jS��;��+��U"��U �H�$��G0��C��c^��o��BꜾ�����5�q���C6��'Y���w��#�����E���:vk��J���)��1��������,���T��B<��@^��?|�T������N��P\i���G���$��x�L&׾�ծ������u�?oU�m�?��k1�*\*���)��#0��K=��+R�Orp�x��y���o�Ѿv��� ��MC��ze�����qu������~�E�a���?�h0 ����������X���&��XG�
�h��끿�∿�{���B|��b^���;����AZ���ȾD棾}���c�i��N���:�mr/�B�*���,��85��D���\��~��%��$k��|-�B�l�,��O��ap�j������e9��D�v��W��C5����-
��6��̙��9���1��uS�9�s��t���  �  �c�7�\�� K�2�z������"ξ㢪�_Ȏ��Lr���P���7�$�%���u��i_���)��&=�1X���{�Yє�5R���׾���"�Q8�.P�(�_�91c�*EY� dD��)����^�־{�Ѿ�������E���8�q8Q�ۄ`��!c���X���C���)��v��뾭�¾�������?h���I�B�2�@s#��q����"�џ0�9F�?d�vN���3������J��U�ZE&���@��tV��Lb��2a��1S��;��% �NU����ҾEfվ���G�a.'���B�`�X��d��Xb�QT�s�<���!��h��"�๾N����A��8dd�;�H��'5���(���#�Eq&�K�0��8B��"[��|�_B�������CѾ�h��A����2�bL�gG_�{g�s�a�P�O�u}6�X������"�X�ؾZ������wG4��rN��_a�Ʉh�CBb�wP�zz7��4���fپl���<ؙ��U��2�g�;�N�q=�P}3�H1�3D6���B�w�V��jr�=$��%?��zٿ��U�L�	���#�o&?�DW�@�f�;j�s`�h�K�f
1�N0��_ �B����ᾠ<�N"�)�%��>A���Y��h�0nk�^�`��L�D�1���v�����ҾZױ�����+��!�i��R��TC�kJ;���:���A�MzP��cf�����QR��D���<ξ�w��.t�k.�dI�k�^���j�^ki��i[���C��S(��w��-��"�⾱&��\��y��1�.��I�e�_���j�.i�j�Z���C��(�^��D��ƾ����&���}�Vb�*�M���@��;�ݸ=��oG���X�"q�Ɉ��᝾�����۾�h�����8�z�Q�t}d��Bl���f��U��;�z��L�����TR�F���@�k�8�g�R��|e��  �  8�9�V96�Z�*�Q���U�����'; P���P���@��Zhs�X�W�t{B�{5�x�1���7��F��]���z������[���0���Ծ��.��,�%.��C8�<�9���1�z�!��5���k�ξGd��ˉ����þ<�����@��+���7�zL:�-�3�a�%��A�m���%�"0žԵ�������}���~k���Q���>��4�YL4�0G=�gO��
h�cm���X��4奄���SJ޾�n�������#�@:2���9� 8��-�@����X�sƾl��s����̾���!��f� ���1��:��n:��71�S�!����3��-۾"ſ�Į��~Ԕ�i���L�i��R��ZC���<��+@�
�L�8�a�}b}�8��68���	��
�Ѿ����$	������,��69���=��9��j+����S������pǾy����ž�#޾iS�����*�,9�K6?���;�Q�/��7�������&ؾ6J���`���o�����J�n��Y��fM��-J���P�9(`�ڄw����2曾Ư��ƾ=�᾿� ������$�)�4�q2?���@�'�8�{)�Z��a �؈޾�Bʾ,�ƾK8Ծ4����(P!�,�3�
�?���B��<��0.��z�b
�,s�fkվ�߼�Q֧����������q�R�^��T�, T��]���n�����f���[��d���Ҿv����Z�V,��j:�S�A��B@�HF5�H#��.�������־�NǾ�Dɾ�ܾ]������n�'�׌8�ЛA��)A��7�df(��/��-�5��̾���G����U��e���+zk�i�[�H�T�5vW�4�c�4x� ������٬�&�¾��۾���6Y��� �o�1��l>��C�->�΁0�"�S���t���о�ZǾ�Ͼ�������.��E=��  �  ������K��������龊8پ��Ⱦ����D������-��0�j�~=Y��%T�$J\��}p�����e��W����c��s;Kkݾ>^C ��o	��7����������R��I�H�žq�������V���ݢ���ʹ���־��������Q��{���g���������`�F�Ծ%�ľ�U���7���:��,~�.}e���W�o�V�LBc���z�+��@ ��"���l¾E�Ҿ �^c���^��?�h�������K�	�u�����پp���꒦�~���1��[r���þ0���� �>��ty��@���������Q��U�Ҿ}C¾�հ��˞�qn���,}�eZh��]_���c��vt�
ԇ��ɘ�@(���R��-}ξ)�޾юﾫ� ���	�kb�S������x	�v���)׾��3D���W���Q���C��"8վax��7	��o��8�T��������aQ�&���7&�`�Ӿ-.þ=t���t�������#���#q��~l��u��߄��ϓ�ot��K跾u�ɾ�ھ��꾦�����FG�>��w�����9��-��Ծ?���N��`����Ӵ��!ʾ��Z%���8��K��(����~�����P���~/�ܻԾ�nþ�B��:����k����w�X�v�Պ��.Q��'������1!���zҾ���?J�%N�b���i��C�(����	���V ��̾A���qG������Z�����Ҿ��p������N�����3�̺��	��� ���\�߾�AϾ|���D�������=銾H��+!w�6�z� ���[��5ǣ����Z�Ǿ&پ�X�T������u#�ș��O�d@�.<����� �H�Ϡž�Ʋ�Ш���o���-þm�ݾ����H�׆��  �  �$��l��gZ�����N��ja��<W������u⾖�Ͼ�"�������������;���䢓����ω��i|Ծ�c澑|�>���[O�������������7+����Zྼ�̾����7ܟ�/ڍ�;낾Sހ�����C�������¾gؾ�e�wx���������Z���1���������(�:�ݾUQɾew������ϴ���������-���x���ʯ���ƾwy۾�v��x���:��������e������������t�&$ھU&ž�W���S��卉�����D��K��9���9���`̾���iF𾙗������;+��,a���
��z
��K��8쾈�ھ2~ž�Ԯ�W���������=j�����%����4��F	Ծ���p����=���� �_��i��%������4�����F�ھ�ž_�����������������
������Xľ��ھv������*�Ť�� �O�P��
"�������2�ھ;|ľE5���}��Ao����������9��|���]�˾3��>��@���<��v����y��YH����7���	���&۾�ľJ���rC��N����Ȑ��(������[l��3nӾ=��{���͂��J��<��c�,G����ee�EP�����P[پ!v¾��������
���~��2���d�������־Uz�#���v��a1�I����
����T������@y��lվ<����b���r���U��.e��Ft���ڭ�a�þ �ھ�������E�����2��G�4����-�������羇-Ҿ%U��٦�N��us�����兟�%豾8Ⱦ)�޾d��@ ��X�p���d��
]���"��(;��O��Ͼ4d���������Y���8(����4��H�̾�+�"����  �  N�ɾ1�پ?�꾤�����������������QJ�'���ɾn���󗞾�����}�������о
�g������1T�rq�����b��}��n;׾B�ƾ�赾�죾ב��I��	qh��X���U��&`�gv��W������C��iϿ��cо)������d��u�q���������0���[߾�[��詩��Z�����/���6;����۾���˨
�SC�������������7T�⾖�ѾVA��k䯾Sɝ�r��3;y�ޕb��oW��uY��nh��"��tÑ�� �������Ǿ0�ؾ#'龮���ī��f����͝�����	�������ؾS����W���T��D+���F���;��H1��G������J��j�{?�Rs��Ƣ�]qӾ5�¾n5��A(�����f����l�h�e��#l�D�~�^�������{����þ}Ծ��侗��������1�!?�TD��I�����0���{վ3c�����A����ҭ������ݾ������|�FD����>�����~����5�Ծyľ�c��ѕ��VS��h�����w�'�u����nA�����(v��þ�pVоh���6�G&�QE
��K�!������
����Y�9QѾ����	E�������w��&ξ(�뾺X�����H����������^�
�����b�"�J�Ѿ�.������7���������m�v�%x��F���㏾�3��OB��h^ľ��վ���t����YB�����I��"��!��P�KH��c�5�Ⱦl���5��i׮� ����EؾP���Y�
���W�7��~�����t����� ���ݾ�;k��M9��s������l��Sx�K~��R��le��Ʉ��9Ĺ��˾�  �  �a����ξ�n�U�P���b+���6�>�9��c3�$��k�����Ӿ���P���Lھ3 ��C�B�(�(�5��<:��#5�<X(�@�#����澰@ɾ����������D�o���T�DA�8�5��j3�w�:�DgK�apc�y����P��~���齾��پK����F!��0��b9��O9�a�/����b�	�����ʾr���-���J�Ǿ_�� ^�ye�4.��8�ְ9�O�1���"�����o���wܾPN��j������zZ��\f�r�M�f=�E�4���6�M�A�ƐU��_p��b������t���\ɾ0��
c�����g(�g�5��<�9�8��,���r��z�]_Ǿ�!���3��q�վ�����V�_�%��5�3C=�SH;���0�4� ��?�����{�پ��������(���V��8Ol�QV��EH��lC�C;H��NV��tl������v���⨾�=��uپ	^�����; �"�0�M6<��W?�%�8��*�%�/���޾K�Ǿ�j���9̾,���e����/�=|<���@�$�;��"/������������׾���(ר��o��K�����r���_���T��R�&�Z���k�|���"���Ƣ�G����lξ���=�P��r)���8�_}A�6bA���7���&����y���=�ھp�Ⱦ�ǾO�׾����[U�%`$�Q6���@��A�3�9��+��������쾾�о{θ�nW��Y���w>����m��{\��T��!U�5�_�s�r�ˎ���v���ߨ�3����־�	��0�
��c���.�sv<���B��J?���2�c! �@�
�oC�oӾ�Ǿ��˾�W�������M+���:�4�B�M�@���5���%��t�Ű�5�/rɾ_ᲾW_���h����2�i�YE[��U��ZZ�	�g�׷}�x���2�������  �  �#���+о����r:���3�uHL��]��5c�?p[�H�Z�-�ho�$�����ؾ�Nо��ݾ"����o�x4�n^M�6�^�B]c�g�Z�đG�w�-���E��ZȾn5��|���m��M��5�?
%����;�G) �Е-�YB���^��ށ�	ϙ����DY߾XD��!�u�<�{�S�}|a�B�b�6�V��W@�]%��
�J�뾚uԾ>2Ӿy������!��\=��wT���a��b�h�U���?�>�$�9�	����L����z��������a�E���/��"�����B��A&�X�6���N�K,n�ʋ��4Υ�PHǾ��&j��,���F�"[��e���a���Q��i9����������7־g�ܾ�i������-��H�8T]��f��b�nuR�JR:�P����L�ܾ\��������I��� f��K��?9�T.�-V*�p8.��9�UiL��f��q��򗚾� ��۾���Q��C�8�ƻQ��c���h�e�`�)�M�i�3��6��0�p��EbܾD,�o'�D���:�(�S�e�~j�4�a��XN���4�x�jT �l/־A/������!#��M�j�`xS��jC���:�˟9���?���M���b�=b�M��!I��ɾH�ﾕ}��$*��E���[�E�i���j�2�^�[H��-��y�	s��)_侼��������)��VE�v\���i��)j�1�]�,�G���,��� ��UH̾�����(������e�ėO�nA�]�:�%�;��D�@�S�m-k�p��T���_����Ծ+^�����13��QM��a��k�W-h�KHX�
�?�$���
�z��KV�����Z�'�3�GEN��b���k���g���W�?��R$�"-
����x¾e�������%z�x�_���L��A���<��Q@��IK���]�gw�沌������  �  ����@Mؾ�D��F)�WDL�x'l�rK������W����h�[H�(�&���
�֦�T8�%����U��!.��P�*<o�v4��!��+�}�e���D�j"�1���Jξ�8�������Z�`R9�2"�P��_�
�Mk	����¤�A9.�s�J�9s�pG��b���)�qs�Њ5��$X���u�:�p����z��_��r=�������d�����:��k�9��d[�=�w��3��b5��8x�X�[��<9����s�����c�����w�/`N��0�s���}�z�f��^��g#��Y:�m[��=��2%���2̾\\ �����B�Kmd���~��܅������at�QV��74����( ��8� ���Q1�v&���G���h����ņ������s��S��1�ˠ�#��X��D*����v���Q�4�7���&����r����3'��8��bR�]�v�Ɔ��4���9�¼���.�׸Q���q�F��·�g��+^n��N��,�2�������F� ��܇��k4��qV���u��~��hi��1߂��l�i�K���(����`ܾ�/������ \w�[�V���?��11�}�)��(��T.���:�}�N��zk����������˾D��������=�O`�f�}��·�ֹ���R��6g�~pE�n%�h��H����p����	�۽!�"�A��^c�=��5�� :�����ѭc�GYA����L� ��:Ͼ-ͨ�h%��e�n�g�P��}<�i�/�2�)�H�*��2���@�O�V��w�R ��g�����پ{����&��^I�!�j�X���s���-���z��V\�d:�n��c+����/N ����B!,��_M��Kn�#ƃ��j��ә��];x��Y�-76����AG�;j¾�{�������	f���K�:��/��,��/���8�G�I��5c�ۣ��N����  �  �ӭ��lྨY�=E6���^������Î�v'��Ծ�����[��5��]��3�8���D��Ӡ��F=���c�����ޏ��&���DO|�-V�2�-�V	�/�Ծ�]���(��2�Q��/��������;�9������R�A�#�&0A�Cl�,���|��ġ���hND�Bl��+������|����7����t���N���)�@��f���P��P0��<&��;J���p������$����	���5Gp��H��!��-����þ'U��ώq�M�D���&��������v���s
�d �'0��!R�
���"ѣ�0Ҿ����E+�9`S�6;z��\���擿��������`j���C�Ou!��	��������sw�[14�<�Y����V���ٔ�S���o����f�̖>��7�}�ĺ����:o���G�^g-��l����H�4\���.��JH�I�n�0ǒ�y���&Y����P�;�'d�@{��k~��f敿˄��Ղ��`�V�:��<�E&�;^�m�
���!���C�N.j�K��%���x��V�������\��4����4��lR��0K����n��1L�YL5��'�����*��w$�{a0��D�g�a�2���Y����ξ��rM%��L��kt��<��Ѡ������U<����|�v�V�W�1�Ҙ�������#�U1.�H2R�H�x�u���D&��s"������]x�ѵP�))�\9���Ӿ����Z�[#e��hF�2���%��b ��!�G(��6���L��n�T���[���}߾ȟ���1���Y�Na��>���� ���
�����p��J�M�'�g��O�����<���9�ʎ_�捂����9���3���	��il���C��m��1��T'žQ���Ӂ��\�x4A�L�/���%��"��n%��.�	J?�Y�U<��㚾�  �  � ����㾓o�];�bhe�w�������R��襒�jC����a�F#:��&��,��+��=��Ī�u�B���j�_"��qޔ��P��u����D��?k\�LL2����S�׾b+��⮁� �O�.�+�L�ȩ�VQ������)��y�t �m]>���j��ʔ�I������V� ���I���s�5���P����ԗ�le�|���T�W�.�w�W� ��������y�*��<P��sx�K[���@���9��'D��f�w��MN���$�MU ���ž落�gp��?B�(J#�KF�n���D��*����H�۹�p�,�0�O�
��5s��
�ԾV�	�_�/�q�Y�+"��z#�����̖�a����q��I��%��K�!�D���!�L 9��`������.��@�������҉�I�m�˥C��{�k[�$��ä���/m�I�D�{*��-����i�D�L����*��DE�B�l�숒��߹�������@��j� Ȉ��q�����l�������g�u�?���.
���`��s�%���H��Uq�]��I%������;ܔ�����(4c�9�����|�F��;Џ�3l��I���1��#������!O!��-���@���^�⧅��;���о
"�}�(���Q�g�{��ʏ�k����ܛ��󒿦h����\���6������i����2�3X��6��Z��2B��>���K��	��XiV���,�ww���վ&ਾ�-��!fb�k.C��.�)�"��U��
�m�$�|�2�_[I��k�꾎����� ��0��6�`�he��xb��3G��"����,����w�ħO���+�M����r�����>�~"f�����ߕ�'���h3���m��s���H��� �s���Y�ƾ2����΀�]Y�}�=���,�-�"�j���U"�Kr+���;�%V��}�M����  �  �ӭ��lྨY�=E6���^������Î�v'��Ծ�����[��5��]��3�8���D��Ӡ��F=���c�����ޏ��&���DO|�-V�2�-�V	�/�Ծ�]���(��2�Q��/��������;�9������R�A�#�&0A�Cl�,���|��ġ���hND�Bl��+������|����7����t���N���)�@��f���P��P0��<&��;J���p������$����	���5Gp��H��!��-����þ'U��ώq�L�D���&��������t���s
�b �$0��!R���� ѣ�.Ҿ����E+�8`S�4;z��\���擿��������`j���C�Nu!��	��������sw�[14�=�Y����V���ٔ�T���o����f�Ζ>��7��ĺ����:o���G�`g-��l����H�3\���.��JH�F�n�.ǒ�w���$Y����N�;�&d�?{��j~��f敿ʄ��Ղ��`�V�:��<�E&�;^�n�
���!���C�O.j�K��%���x��W�������\��4����6��oR��2K����n��1L�\L5��'�����*��w$�{a0��D�g�a�3���Y����ξ��rM%��L��kt��<��Ѡ������U<����|�v�V�W�1�Ҙ�������#�U1.�H2R�H�x�u���D&��s"������]x�ѵP�))�\9���Ӿ����Z�[#e��hF�2���%��b ��!�G(��6���L��n�T���[���}߾ȟ���1���Y�Na��>���� ���
�����p��J�M�'�g��O�����<���9�ʎ_�捂����9���3���	��il���C��m��1��T'žQ���Ӂ��\�x4A�L�/���%��"��n%��.�	J?�Y�U<��㚾�  �  ����@Mؾ�D��F)�WDL�x'l�rK������W����h�[H�(�&���
�֦�T8�%����U��!.��P�*<o�v4��!��+�}�e���D�j"�1���Jξ�8�������Z�`R9�2"�P��_�
�Mk	����¤�A9.�s�J�9s�pG��b���)�qs�Њ5��$X���u�:�p����z��_��r=�������d�����:��k�9��d[�=�w��3��b5��8x�X�[��<9����s�����c�����w�/`N��0�r���}�x�f��^��g#��Y:�g[��=��.%���2̾Y\ �����B�Hmd���~��܅������at�OV��74����( ��8� ���Q1�v&���G���h����ņ������s��S��1�͠�(��\��H*����v���Q�7�7���&����r����3'��8��bR�W�v���/����8㾿����.�ԸQ���q�D��~·�f��)^n��N��,�1�������F�!��݇��k4��qV���u��~��ii��3߂��l�l�K���(����dܾ�/������&\w�`�V���?��11���)��(��T.���:�~�N��zk����������˾D��������=�O`�f�}��·�ֹ���R��6g�~pE�n%�h��H����p����	�۽!�"�A��^c�=��5�� :�����ѭc�GYA����L� ��:Ͼ-ͨ�h%��e�n�g�P��}<�i�/�2�)�H�*��2���@�O�V��w�R ��g�����پ{����&��^I�!�j�X���s���-���z��V\�d:�n��c+����/N ����B!,��_M��Kn�#ƃ��j��ә��];x��Y�-76����AG�;j¾�{�������	f���K�:��/��,��/���8�G�I��5c�ۣ��N����  �  �#���+о����r:���3�uHL��]��5c�?p[�H�Z�-�ho�$�����ؾ�Nо��ݾ"����o�x4�n^M�6�^�B]c�g�Z�đG�w�-���E��ZȾn5��|���m��M��5�?
%����;�G) �Е-�YB���^��ށ�	ϙ����DY߾XD��!�u�<�{�S�}|a�B�b�6�V��W@�]%��
�J�뾚uԾ>2Ӿy������!��\=��wT���a��b�h�U���?�>�$�9�	����L����z��������a�E���/��"�����B��A&�R�6���N�C,n�ŋ��/Υ�IHǾ��"j���,���F�"[��e���a��Q��i9����������7־h�ܾ�i��	����-��H�;T]��f���b�quR�NR:�T���S�ܾb�������J��� f��K��?9�V.�-V*�n8.��9�PiL��f��q��헚�� ��۾���M��?�8�ûQ��c���h�b�`�'�M�g�3��6��0�o��EbܾE,�o'�E���:�*�S�e��j�8�a��XN���4�x�mT �r/־G/������%#��U�j�fxS��jC���:�Ο9���?���M���b�=b�M��!I��ɾH�ﾔ}��$*��E���[�E�i���j�2�^�[H��-��y�	s��)_侼��������)��VE�v\���i��)j�1�]�,�G���,��� ��UH̾�����(������e�ėO�nA�]�:�%�;��D�@�S�m-k�p��T���_����Ծ+^�����13��QM��a��k�W-h�KHX�
�?�$���
�z��KV�����Z�'�3�GEN��b���k���g���W�?��R$�"-
����x¾e�������%z�x�_���L��A���<��Q@��IK���]�gw�沌������  �  �a����ξ�n�U�P���b+���6�>�9��c3�$��k�����Ӿ���P���Lھ3 ��C�B�(�(�5��<:��#5�<X(�@�#����澰@ɾ����������D�o���T�DA�8�5��j3�w�:�DgK�apc�y����P��~���齾��پK����F!��0��b9��O9�a�/����b�	�����ʾr���-���J�Ǿ_�� ^�ye�4.��8�ְ9�O�1���"�����o���wܾPN��i������yZ��\f�p�M�d=�B�4���6�G�A���U��_p��b������t���\ɾ(��c�����g(�c�5��<�5�8��,���p��w�[_Ǿ�!���3��s�վ�����V�b�%��5�6C=�WH;���0�8� ��?�������پ��������(���V��?Ol�QV��EH��lC�A;H��NV��tl������v���⨾�=���tپ^�����; ��0�I6<��W?�!�8��*�#�	/���޾I�Ǿ�j���9̾.���e����/�A|<���@�(�;��"/������������׾���.ר��o��O�����r���_���T��R�(�Z���k�}���"���Ƣ�G����lξ���=�P��r)���8�_}A�6bA���7���&����y���=�ھp�Ⱦ�ǾO�׾����[U�%`$�Q6���@��A�3�9��+��������쾾�о{θ�nW��Y���w>����m��{\��T��!U�5�_�s�r�ˎ���v���ߨ�3����־�	��0�
��c���.�sv<���B��J?���2�c! �@�
�oC�oӾ�Ǿ��˾�W�������M+���:�4�B�M�@���5���%��t�Ű�5�/rɾ_ᲾW_���h����2�i�YE[��U��ZZ�	�g�׷}�x���2�������  �  N�ɾ1�پ?�꾤�����������������QJ�'���ɾn���󗞾�����}�������о
�g������1T�rq�����b��}��n;׾B�ƾ�赾�죾ב��I��	qh��X���U��&`�gv��W������C��iϿ��cо)������d��u�q���������0���[߾�[��詩��Z�����/���6;����۾���˨
�SC�������������7T�⾖�ѾVA��j䯾Sɝ�q��1;y�ەb��oW��uY��nh��"��oÑ�� ��ل���Ǿ(�ؾ'龤�������f����ɝ�����	�������ؾP����W���T��E+���F���;
��K1��G������!J��j��?�\s��Т�fqӾ<�¾t5��F(�����k����l�i�e��#l�?�~�[�������{����þ}Ծ��侍������	��1�?�PD��I�����0���{վ0c�����A����ҭ������ݾ������|�JD����>���!��"~����=�Ծ�ľ�c��֕��ZS��l�����w�+�u����oA������)v��þ�pVоh���6�G&�QE
��K�!������
����Y�8QѾ����E�������w��&ξ(�뾺X�����H����������^�
�����b�"�J�Ѿ�.������7���������m�v�%x��F���㏾�3��OB��h^ľ��վ���t����YB�����I��"��!��P�KH��c�5�Ⱦl���5��i׮� ����EؾP���Y�
���W�7��~�����t����� ���ݾ�;k��M9��s������l��Sx�K~��R��le��Ʉ��9Ĺ��˾�  �  �$��l��gZ�����N��ja��<W������u⾖�Ͼ�"�������������;���䢓����ω��i|Ծ�c澑|�>���[O�������������7+����Zྼ�̾����7ܟ�/ڍ�;낾Sހ�����C�������¾gؾ�e�wx���������Z���1���������(�:�ݾUQɾew������ϴ���������-���x���ʯ���ƾwy۾�v��x���:��������e������������t�&$ھU&ž�W���S��㍉�����A��K��5���9��z`̾���aF𾏗������1+��"a���
��q
��K��0쾁�ھ-~ž�Ԯ�T���������>j�����(����4��L	Ծ��x���>���� �_��i� &������4�����M�ھ�žc�����������������
������Xľ��ھn������*����� �J�K��"�����م�,�ھ6|ľA5���}��@o����������9������b�˾9��E��I���<��v������^H����@������&۾�ľN���vC��Q����Ȑ��(������[l��3nӾ>��{���͂��J��<��c�,G����ee�EP�����P[پ!v¾��������
���~��2���d�������־Uz�#���v��a1�I����
����T������@y��lվ<����b���r���U��.e��Ft���ڭ�a�þ �ھ�������E�����2��G�4����-�������羇-Ҿ%U��٦�N��us�����兟�%豾8Ⱦ)�޾d��@ ��X�p���d��
]���"��(;��O��Ͼ4d���������Y���8(����4��H�̾�+�"����  �  ������K��������龊8پ��Ⱦ����D������-��0�j�~=Y��%T�$J\��}p�����e��W����c��s;Kkݾ>^C ��o	��7����������R��I�H�žq�������V���ݢ���ʹ���־��������Q��{���g���������`�F�Ծ%�ľ�U���7���:��,~�.}e���W�o�V�MBc���z�+��@ ��"���l¾E�Ҿ �^c���^��?�h�������K�	�u�����پo���蒦�~���1��Xr���þ+�⾽� �:��py��@���������H��M�ҾuC¾�հ��˞�mn���,}�bZh��]_��c��vt�ԇ��ɘ�E(��S��5}ξ2�޾ێﾱ� ���	�pb�W������x	�{��*׾��5D���W���Q���C��8վ\x��4	��o��8�O��������\Q����.&�X�Ӿ%.þ7t���t�������#���#q��~l��u��߄��ϓ�tt��Q跾}�ɾ#�ھ��꾰�����KG�C��w�����<��-��Ծ?���N��b����Ӵ��!ʾ��Z%���8��K��(����~�����O���~/�ܻԾ�nþ�B��:����k����w�X�v�Պ��.Q��'������1!���zҾ���?J�%N�b���i��C�(����	���V ��̾A���qG������Z�����Ҿ��p������N�����3�̺��	��� ���\�߾�AϾ|���D�������=銾H��+!w�6�z� ���[��5ǣ����Z�Ǿ&پ�X�T������u#�ș��O�d@�.<����� �H�Ϡž�Ʋ�Ш���o���-þm�ݾ����H�׆��  �  8�9�V96�Z�*�Q���U�����'; P���P���@��Zhs�X�W�t{B�{5�x�1���7��F��]���z������[���0���Ծ��.��,�%.��C8�<�9���1�z�!��5���k�ξGd��ˉ����þ<�����@��+���7�zL:�-�3�a�%��A�m���%�"0žԵ�������}���~k���Q���>��4�YL4�0G=�gO��
h�cm���X��4奄���SJ޾�n�������#�@:2���9� 8��-�@����X�sƾl��p����̾�����c� ��1��:��n:��71�N�!����3��$۾ſ�����yԔ�d���E�i�
�R��ZC���<��+@��L�>�a��b}�$8��<8���	���Ѿ����$	������,��69��=��9��j+����U������pǾy����ž�#޾hS�����*�,9�G6?���;�L�/��7�������ؾ/J��`���o�����D�n��Y��fM��-J���P�=(`��w����8曾 Ư���ƾE��ĳ ������$�.�4�v2?���@�*�8�~)�\��c �ۈ޾�Bʾ.�ƾM8Ծ5����(P!�,�3�
�?���B��<��0.��z�b
�,s�fkվ�߼�Q֧����������q�R�^��T�, T��]���n�����f���[��d���Ҿv����Z�V,��j:�S�A��B@�HF5�H#��.�������־�NǾ�Dɾ�ܾ]������n�'�׌8�ЛA��)A��7�df(��/��-�5��̾���G����U��e���+zk�i�[�H�T�5vW�4�c�4x� ������٬�&�¾��۾���6Y��� �o�1��l>��C�->�΁0�"�S���t���о�ZǾ�Ͼ�������.��E=��  �  �c�7�\�� K�2�z������"ξ㢪�_Ȏ��Lr���P���7�$�%���u��i_���)��&=�1X���{�Yє�5R���׾���"�Q8�.P�(�_�91c�*EY� dD��)����^�־{�Ѿ�������E���8�q8Q�ۄ`��!c���X���C���)��v��뾭�¾�������?h���I�B�2�@s#��q����"�џ0�9F�@d�vN���3������J��U�ZE&���@��tV��Lb��2a��1S��;��% �MU����ҾCfվ���G�_.'���B�]�X��d��Xb�MT�o�<���!��h�{"�๾H����A��1dd�5�H��'5���(���#�Gq&�N�0��8B��"[��|�dB�������CѾ�h��D����2�"bL�kG_�~g�v�a�S�O�w}6�Y������"�X�ؾY������uG4��rN��_a�Ƅh�@Bb�wP�vz7��4���`پf���7ؙ��U��+�g�6�N�q=�N}3�H1�5D6���B�|�V��jr�A$��*?���ٿ��U�P�	���#�s&?�HW�D�f�;j�
s`�k�K�h
1�P0��_ �D����ᾡ<�N"�)�%��>A���Y��h�0nk�^�`��L�D�1���v�����ҾZױ�����+��!�i��R��TC�kJ;���:���A�MzP��cf�����QR��D���<ξ�w��.t�k.�dI�k�^���j�^ki��i[���C��S(��w��-��"�⾱&��\��y��1�.��I�e�_���j�.i�j�Z���C��(�^��D��ƾ����&���}�Vb�*�M���@��;�ݸ=��oG���X�"q�Ɉ��᝾�����۾�h�����8�z�Q�t}d��Bl���f��U��;�z��L�����TR�F���@�k�8�g�R��|e��  �  ���G̀�U�j��TJ�b_'�8��ٳվ*���7{��U�_�7�<� $�����a
���������-))��"D�GFj��z��c���ᾦ���r/�YSR�Hq�V���7	����}�}d�c�B��!�^O����� �����O�3���U���s��h��݄��{��a�P?��������ƾ���G�����T�cm5�������
��
��M��p��F2��}P�b�z�������������Q';�3M]�\9y�PY���ك��lv�s]Y��7�d�ڞ ����^�F���i�?�Q�a�E�|�gs��A���u�T�W��5��5�o9뾪u���▾z�w��tP���4��H"��3�,��_��n��.�-�F��Vi�����鬾�׾��pc'�5WJ��*k�Uρ�����o�����q��R�HX0���g���R����e��F_-��&O�go�#e������3�����o���O���,���������b��� Yv�jS��;��+��U"��U �J�$��G0��C��c^��o��EꜾ�����5�s���C6��'Y���w��#�����F���<vk��J���)��1��������,���T��B<��@^��?|�T������N��P\i���G���$��x�L&׾�ծ������u�?oU�m�?��k1�*\*���)��#0��K=��+R�Orp�x��y���o�Ѿv��� ��MC��ze�����qu������~�E�a���?�h0 ����������X���&��XG�
�h��끿�∿�{���B|��b^���;����AZ���ȾD棾}���c�i��N���:�mr/�B�*���,��85��D���\��~��%��$k��|-�B�l�,��O��ap�j������e9��D�v��W��C5����-
��6��̙��9���1��uS�9�s��t���  �  ����2���π��c\��4�^s��pݾ����H�����W�"�2��y�eu	�� �����nA����;���<:���b�~A��(����X���R=�Q�e�B����U��S��H"��Z�z�q�T�}{/��o�����T��Q���� �N�C�|j�?d���:���ޒ�+݊��v��O���'����|y̾���f{�}�K��+�� ������ �]� ��h����'�(G���t������lƾh����##�%�J�	Dr��N���J������Dև��in�*�G�C$���	�||�������(,�KQ�#�w�ee���y���⑿g��
�k���C�
���`�� ���
���p���F��Y*����Aj�р	�@��\_�R$��<�/�`�TL��{N���޾�e���3���[��ဿ�����9B��~�����e��@?��.�����P���v��{�e�;��b��u��ݐ�̕�eꐿ~�����a���9�����_��������9"n��@I�&�0��� � �����0�L&�H|8�j�T�Fg}������þi�������"D�el�����͓�Ƞ������6���}\�P<7��X����XM�5�3)�I&L���r������c�������$�~���W���/�,��7�ܾ�C��΍�,�k�9K�{5��x'�K� ��j �?&���2���G�Og��f��֚��ދ־c���B+��R�(rz��h��bg���ޕ����v�EP�p,������W{����9�3��X��~�V쎿Gꖿ�A���f��6r�*J�e'#��@�(+̾V���)���7`��{C��0�]�%��C!��#�'+�o:�i�R��Vv��锾и��)��@�8�a��|�����e����ӓ��H��]�j��*D�'#�L���U������s5@��mf�����풿�  �  O�=�3�˿"��t솿z�N����xT꾕沾PQ��ZBd�?�A�-P,�\� �6��ֺ"�<r0���H��n�
���������F4&�U\� ����*��KcҿI��~�Q3࿻ſ���xO���Q���3��(.�UjA��k�J����]��b�տ���%�쿟�ݿm��)����<x��<����־ot��]i����X�N6;��2)�x �;���'�vs8��T�a'��%����оAr	�:�6���p�Zu��U����ۿ>��F�꿵MؿJ���ԏ��UQq���D�Y�.�<�1��4M�me~��������^R޿#1� 5��Dֿ�嶿x�����d��b-�����Ǿ���Ĕ|��(U��7<��.�,�(���+���6���K�m��Տ�C��p��?���9L��������1ʿ@$俦/ￄ&迎ѿ!��������Ud��?��J1�q<��w_��V������Pοo�濱����kjοM߬�m���K0T�'!�"L��W�~����z���X���C���8��56�F�;���I���b�$���m��x�˾I��|-���b��*������q�տvw������k�ȿ��DD�� �Y���;�zu6���I��t�h5��ϔ����ٿ���m��[�w�ſ�����>��,E�A?���F�������(y��L[�*:I�v@���?���G��tX���t�w6���Ѱ�1�Y����>�o�x�Ő�����.0߿)�￥�xܿq"��ֹ��k�y�M�'7���9�T-U� ���W����ſ��ῷ��E��t�ٿC3���Ж�'Ck���3�g	���Ծ: �����(jn��U��fF���@���B���M���a�zx������j���������mQ�������?�̿m��G����V�ӿ���_
���&i���C��5��A���c�ڎ���=���mпf���  �  t3�)�ۿ2CĿ~k������j�I�]#��|辘'��ƍ�kOh��+F���0��$�0�!�\�&���4���L�1�r��J���彾x��3#���V��j�����̤ʿ�(߿V�R�׿S���4���s�|���K�}k/��*�J�<���d��J�������Ϳ@����,�տ]����r��iq�3�8��#���վ2������8]�+�?��q-��$��$�8�+���<���X�[큾1���I@Ͼ���	3��Qj������඿��ҿR����Eп{o��D���fj���?�#�*�b�-�R�G�O�v��P��1 ���ֿ$��L῏^οG�������G�^��#*��m��>ǾV)���.��Y�#�@��C2���,���/��;��P�.q�a��K|����辻9�ӤG��O��:����¿B�ۿ	�fi߿�ɿ����{9���)^��o:�oI-���7���Y�:#��I��5�ƿAD޿a�濵O޿� ǿ�(������APO���(t�;4���򘾼�~�_>]��"H��<��J:���?��MN���f�����c���Vk˾���j*�Du]�TՍ��y��ο��⿕��@hۿ���ᆡ�w^���T���7�h2��D��dm�r���h;��!�ѿ��7��ۯٿƶ��#���©y�MA��O�� ��c���?���b}�I�_�(yM���D��D���K�t�\���x�Z��������h߾��~.;�6r�ݥ��n ��a ׿���忧oԿ0����ؖ���r� H�W3���5���O���~���������ٿ4����C�ѿ峿�I��se�Q�0�D��VԾ�#��� ���r��aY���J���D��G�z�Q�p^f�ԇ��O!�����}�8p�v�L�}ꃿ~4��ſ�3޿ڮ�F��I̿�������j�b��.?���1�ۖ<�4^��Z��`s���ɿ�S��  �  ��˿�/Ŀ�G�������p�i'=�O��k��r��-C��|v��[T�26>���1�(w.�(�3��B�2[�w��$A��m(���I�Ԭ��9H�U�}����������Eǿ�i˿������S׎�)]g���<��o#����3/���R��_��Ƴ���@��T�ȿ�˿�����%���zV_�͂.�ە�k�Ծ�ͩ��:��]Ik�ɥM���:�Z1���0�^&9�>�J�gg�|5�����̴ξG���q)��2Y��b���ि�ü��2ʿ_ɿ�s��¡���M��)@W���1��q��!�k9��Hb�c����<���}��7�˿�6ɿ���ѣ���炿(�O���!�����B�ǾHӡ�����7�g�hkN�A`?�R�9�u�<� �H�1^�������>���O�����;�o�n��Γ�>r���yĿ;pͿ�ǿ�괿:���j|��M���-��"�1~+��I�$w��w�������ƿo?ο��ƿl��gԗ��[v�@�B��U�������o��=Z���mk�E�U��I���F�{�L��\�{+u��-��������̾������"�O�%G��>���1��Ǿʿ%�ο �Ŀ�x������:o���D��+�_'��`7���Z�����x颿zv����̿�8Ͽ�9ÿ3���叿�g�θ6�t�����)����\��������m���Z�~WQ���P�� Y���j�G���2D��5�����޾"��U�1�H`a�~��  ������5Yο~�Ϳ1���&˥��u���_�c#:�ؚ'���)�o�@��j��y嫿
ÿ!Ͽo�̿�b�� �74���*V���(����վ^ͮ�����iz���9g�K�W��^Q��S�$b_�u�t��u��١���¾u������@���s�Uk��+��$ǿ�
п�Jʿ�t��M���~�����Q�v_2��&�0��M�N�{�5���Oٴ�M�ȿ�  �  ���r���u��O���C�U���-����b徚彾�ӟ�Q㈾�Zo��W�B�H���D��WK�0�[��v�𾍾W0��q1ƾ;�-��"R6���_�ʅ�ի��A󦿆���4����<���Yt���H�i&������b��18�x�`�3����ߚ�˯��ȩ������A��\s��>H�c"�3���ؾ1��,|��熃��h�!�R�XH�3sG�p#Q��d��`�������I���:Ӿz� ��`��rC��$n�2ь�;���[ ��O�������	���%e���;�x�������b�#�^E��o��_��,����C�������_���	���)f��g<�����a��{0ξ.d���m��1���th�?�V��P�W�S�r9a���x��f���飾YR��H��!�dk-���T�c8��hI��5B��C���hc������X�����Z�&v4����L��{C��Q1���V�.����
���զ�����!L��3���{��~[��3�		�CY�w�Ⱦ�����9��_6��z�n�R�`�o]�|Rd�ju�O>���S���U�Ӿ���sg��)=��df�~6����Wl���~��oF���򓿶�{���P��d.�m�M��#�_�@���h�,􊿉��k㫿����!�
l����{��~P���*�����Y�P3ľ�����������ys�<h��kg�q��x��ef��װ��dc��b����&���K�bZv�,�����E��lv�������0��qom�:D���%�b����j{+�*�L��{w�����6�����L���!����X��1�l�mC��|��F�ZH۾z]��>��\9���n���Ho�t�g�A�j�Hx�Ψ��[��ମ�o�˾�M��Q�G�2���Y��Ԃ�|痿৿�������+��<��	�_�iK9�Ӵ��+�]����5���Z�᥃�D#��U⨿�  �  m��N<��$�t�ŤY�{�<�3�!��0��:�mOҾ�̷�|ᠾ����!#~��l�#�f��/o�=���ԑ�����_����.پ�_���!���'��JC��o`�o�z��х�1P����H6h�1�G�zJ'��4��1���Y��;�������8�$FZ�:�w��~�������灿�l�=�P��3�_��%��l�ʾ�ǰ����0���x��j���i�L3v�`��̧��������ƾ���7����D�0��L���i�������F�6Rz�<�]��W<����ɞ��W�����:5��~$�˦D���e��a��q���?!���~�ILe��CH�m,��[�a� ��^��ľE���n��a��2{�r��ev��ك�9���;�����X־K�����3�"�lB=��BZ�rv��c��	q��ɫ��y~u�S�V��p5�t���q����V7����'�2�϶S�z|s��l��$������rbz� _�_	B�`G'�M���0���Zݾ(�¾p8���=��[Ҋ�s��nc�������KǞ�����˾����}�J��^�.��#J�3Jg������J��%׊�	���O�o��:O�\/�"!�̨�J����� #��JA�U�b�w%��n�������^��YNu�O�X��<���"��P�����Iھ�������:��GD���@���؄����_��謨�����־@��G�
�r��x�8��)U�3�q�aք�Z>��	���N����e���D�:�%����;�+�����,�hL��l�i惿���8���7����k���N��3�4����u�B�Ѿm���	��Ĕ���������s݆�8F��6i��R3����ƾ��྅b������(��wB��{_��?{����O��DA��d�z�l�[�f_:�ޡ�:2
�X�������4�6�F�W�<�w��w���  �  ~�R��Q���H���;�0-�9������q��C��N�Fgƾ�m��+񚾅���񊾏����䞾����XY̾)�f��}<�o����"���0��?�d�K�wOS�%rR���G��P5��.�1!���-GҾQξH�ܾ�9�����tm+�w�@�[O��DT�R0P��ZE�X7�>+)��J�����!�
򾘂ؾn���7��hȖ�; ��!���<9��٥�E,���jվD�ʨ�!"�����f'�&r5�0�C�I�N���S���O��SB�#�-�� ��" ��`߾��ξ5IѾ>��V�LQ��3��qG� $S�M4U�\�N��VB��4��8&�v���_����'��Ӿ�޺�Vɥ�5���T���&q���<��9[��UCʾ�)�C���=�
��S�?"��w/�[�=��kK�hU�!JW��P���?���)��N�����W�߾^�վP3޾����~��(���>���O�nlX�KLW��[N��A�<�2��J%��N�1���'��F뾥�Ѿ
���ر��r���&�����7�������hzپ|�H�	�ŋ���)���7�`�E���R��AZ�w}Y��"O���<��%��������G��J޾�,�e�����3��I�{W�ˣ\��X���M�9�?��j1�x$�:���B�W"�����!ϾA���ʦ��������5���׵��0̾_w���|���<���"��/���=�:�K��/W��/\�aX�L�J��5��Y��N����Y�޾��=�������#��;�:sN���Y�U�[��@U���H�{�:���,�Vp ����\	����uM�ytǾ�'���#���|��/��w�������S@վ����)�z�h��yr'�A�4��C�,�P�7OZ�)�\��2U��D���.�@����+U���޾JQ��� ����X,���B�bT��  �  &���*��W,�vu,�!{,�[^,���*�b�%��Y����Q���r۾�迾�0�����(0��Awž��������W�'���+�k�,�7�,�g�,�u�,��*�B�$���I��`���׾׼�]�����Gk���rʾ���#�2��r!�k�(��>,��-�-��-��,�%*��#�m����	����XҾɛ���Ы�J���i���Ͼ�0����v���"��s)�M,�4�,�4�,���,��,�_
)��!������쾨G;6U���ݪ�����Lg����ԾR����
|��n%���+��$.�6�.���.�2�.���-��*�06"��������;;�������ն��FnþW^޾�2��hE�Q��S�(�G,.��0��S0�P0�-F0��/�F�*�b$"�k
�������(V̾��kɱ�@����ʾ���"�����8"�u�+�,Q0���1�l�1�L�1���1��90�vP+���!��%�o��;���˾�(��7��C���=Ҿ���������%�BX.��w2�t�3�e�3�,�3��3��1�"�+�W�!����D)�M澚o̾���=����ľ4�ھ@S��yz��/�sx)��%1�-�4��b5�'V5��V5��4��N2�<�+��� �V�����a⾂�ɾ�ͻ�7��:eǾ�߾14���������*���1��n4�L 5�?�4�� 5�8\4��L1�?%*�e\����yf��$�ݾlƾQ����A��'�ʾN��<�����ov!��E,��o2���4��05�,5�-25��K4��0�|�(��@��v��v����پ�.ľ�����f����ξ��}�t��+�#�x�-�%c3��L5�Z�5�i�5��5��H4�b0��Q'�h(�9
�y��־�r¾������ |Ӿ%��N�����G&��  �  ���f�6| ���-�:[<���I��6R���R���I���8���!�p
��|�)Ծ��̾%iؾ�^������:'��+=�M�)�S�*Q�s9G��9��9+����K����y���d~ܾ�¾kw������k�b勾X��"����6���:Ѿ�������h�f��bn%��S3�z�A��M��T�n�Q��E�E�1��Z������mkо�UϾ���1g����4/�#�C���P�bT�p�N�j�B�{�4�+�&�"��_�;��dI�W�Ӿ�������f��������]��4���u���}�۾�����6���a�Jd+�O�9�]�G��/R�b�U��7P�/aA��,��v��h��ྕ�Ҿ�%ؾ���}%��v"���9�G�K�nV��{V��N�$�A��d3�Y�%�����2���B�q�Ҿ�f���+��落�z����!��VG���`����Ѿs��K���f�V����%��l3�T�A��O�שW�waX�]�O��>���'�"8�a?��C྆�ؾ���=� �z��Ҽ-�G�C���S���Z�c�W�7N��]@�2�s%�p=�"��{�J뾬�Ѿ�����x������꛾�V�����;�Ⱦ�ᾟ����+
�,���E!�[�-�j�;���I�+�U�.\�ݬY���M�d�9��c"��������g��O߾����e	�a��a97�ǍK�+�X�\�,�V�8K���<�<�.�41"�̝���Ⱦ�� ���ʾ�ȴ�2���w`��p�������c���uо��I��Y���K�H%�D2�}C@�h5N���X��j\���V���G��b2�"��\�� 쾨�޾N��c��J��b�'��?��RQ��R[�ݲ[�3�S��F�"�8�++�Y���i�Ϸ�7�����ܾ}Pľ�⯾�&������3��� ���¾�9ھ���8���  �  ���d>��&#��!>�(F[�/Mv�'���hp��'X���l�L�L�,�������9�������33��{T�;s�K?������{/��q�6&U�<8�@�`0�4h��QξTm����������{��k��h��s�Gt���0E���¾��޾	�����c\,��`H�}be��h~�h���↿d�~��;c��5B��~"�|�	�Ϗ��$����ND��k>�_�_��{��S������:���8h�jZK�Y/�T9����ږ�<ž�n���h�������ku��j��*l��v{�5K����������;���ގ�����6��S��o��.���s������Hx��aZ�)9�Ia�T;�����	� ���S�+�\uL��l�|��/��$5����|��Rb�0E�a�)�c�����`�޾Y�þ�z���ј������y�1�x�;�i/���d�����oþ;_޾���5��ޡ(�g�C�^�`���{�}`��t-��.���kr���R���1��w�� �\���\�tJ�m�9��Z��y�M���P������6�w���[��?���$�c!�q���ܾ��¾$ᬾ�����3��{���C��D���ZC�������׺��@Ӿvg�@F��Z���4��P���m��M���Ɋ�k񊿯Q���Jk�2>J�h�*�����E� �����B'��lF�/�g����)\��~��jJ��p`p�B�S�o=7��r��	��
�1zվ5Ƽ�
���X���c���!����|���֌�N��S(��-%¾R�۾sK��!H�s�#�z=��@Z�ٖv� y������\@��<�~�v�`��c?���!�"F����ǈ����Ll1�lR��er�MÅ�2����Љ�V����g��eJ�g/�_�����=龕ξ�������E��>�����ؓ��K��� ���y���˾v��  �  D��f ���/���W��������y2��2�����lm����{�vlO�a�*�����0�U���$2���X�*Ⴟ��O������Ϣ�1t��oz���N�>�'�T"��޾� ��a?��aT��+�k��_U���H�זF���N���`�f+}���������<�̾������=��g��{������'V���p���`���Ҍ���l�y�B�3"�(�3/�&9�
E>�"�g��a�������Ũ�"6��a���n�k��0A��u������о|^��U'���L��,�c��P��H�s�I���U��l��,��Ǜ������ܾ���$�%��L�=Uw�7'��lM��#̪����vԚ���,&`��o8����?��%���*�-�M�M�y��撿G���⿫��&��l���R��S�`���7�i�����!�˾�*���N���b���Ek��[���V��[�nk�$?�����V���{Lʾ���L���#5��r]�鲄�<���맿xҬ�L^��{<�������9U�Z�0�����>�D��E^8�C_�$��M���i���u��o3���ܕ�C�����U���.�;����7Ǿ�������p��;t��h��Kf�[�n����E ��3~������ݾ���n!�fYE�[o�/���$����i�����[k��ڐ���t���J�>*��%��+��5'�%CF���o�d��7���Yͬ�r���`E���Ǐ���s�dI�1�$��@�85ᾂ���pr���y��1ԁ��_p��<g��mh�L�s����N����੾��ž�~�5Q��b,�R�R���}�_r��~������uV��0��`���hYf�g�>�v�"�v2�H��j0���S��Y�4���Ϊ���b�� ê����눿V�e��<����5��}�վ�j���h���N��ж~���n�_&i��m��|��֊��j��$ȳ�LaҾ�  �  �����G�?�V�s�����Z���ſK�˿�lÿ�׮�o���o�GJB�P�%�����*��!K�Z{��ؙ�T��Րƿ��˿$���	F���t��wh���5��*���ܾn���M��{�p��FQ���<���1�f0�t�6�7(G�W�a�W���'��y%Ǿ���0�"�0�P������s�������ɿ߾ʿ�����c���,��}Y_��-7�!G!�� �;3�RZ�� ��O��������ɿQ�ɿi���-h��b͆��IV�>'������˾�w��8����e�>�I���8��1��#3���=�͵Q�j�p��������e�پ<�
��e2���c����I������O̿�ȿv����"��恿WR�Q�/�h� ���&��.A�8�l��ߑ�n����nÿ09Ϳ�Oȿz3��c͛�~��I�%�6��ľ���l���R�i�� R���D��!@��D�R�Tli�p.���&���0¾���#W�+9E�Foy�Bl���a��A�ǿ�RοK2ƿ;���QK���Ou��/H�.�+���#�Ƿ0�TQ�Ҁ��
��/���D�ɿh�ο?0ſ����ߓ���n���<�p�����ѽ�
��� ��;o�[[��
Q�ߤO�r
W�;�g��.��yՔ������׾Q����*��#Y�@އ����������'Ϳh�ο¿�j���0���\g��-?��D)�(�i�;�0b�� ��Q�����W�Ϳ;�Ϳ/˿��z���㊿�{^��:/���	��;ܾг��������i�~X���P���Q�@�[�	o�����׷���廾vk�P���9��gj��j��0����Ŀ_Ͽs̿^"��D��O����nX���5���&��,�3�F�l�r����Xq���ƿ�ϿG�ʿ|̸�;f��r���0<N�XF"��P �"wξ�O������AY}�8qe�5�W���R���V�O�c���z����s\��Dʾ�  �  *��io���L�Ä��L��D�ſ��ܿL=係�ڿ��¿������R��H2��)� �7���\�鉿�j��H%ɿ�_޿�#�m�ؿW���^���<�{��@A�����޾\���z����b�T%C��[/��%�VX#�M�)�cF9�vkS�B�{�Ѧ��Ϳƾi��T1+��`�f�������ϿJB�;8��XԿ��fG��+�s���E���,���+���A�֙m������\��<�ѿMH�O>���ѿ<&��������f�PB0�<��|̾
R���[��\�V���;���+���$��k&�o[0�"�C���b�?���g����i۾ƪ�y=�Zv�<�����
~׿<�俍���3Ϳ�6��ɘ���wd��D=��2,���2�Y�P�ic���򠿫.��Frڿ������ʿD򫿼U����V��@$����P�¾����J���I[��GD�j�7�]u3�@�7��{D��<[�D�~�ʙ�	%�������� ��VR��������ȿ�B߿/�濿�ݿ*�ſॿ���iX�vA8�/�Y�=�f�b��������a̿G���y�`#ܿD�¿Ca���;���!H��z�����Һ��㗾[$��ra���M�a#D�p�B���I�S�Y�]t�zP���5��C[׾O
��3���h��7��tǵ��&ӿ0U忄F�cؿN���@K��J�{�A�M�R�4��3�:�I���u�Ġ���^��n�տoO��H�r�տ�8��eƗ��"o��v8�����tܾ����`����!w��[�TEK���C��D��8N�:�`�lW�A���Z}���辸_�G�C���|��b��tW����ڿ���A��]п�U������ʋj�qGC��$2�f�8�Y�V�9>������1�ÿ�"ݿr}近��+wͿ*���)���3\��y)�ϯ��̾)5��Qቾ�"o�Q�W��J�|�E�G�I��V�cl�_��������7Ⱦ�  �  ����U�Q��ψ�����_Ϳg>�lX�%S�lʿ*����;��sXX�6�6�?-��6<���b�;\���|����п�'�{<�D��ƿbb���}����E���Fk�!���ㇾL�^�v�>�v+��� �A�*�%���4��O���w�풚�z0ǾE���.�!�f��������$׿�2��@��ܿ����m����z�K�3 1�|�/�t�F���t���������&�ٿE�a=�C�ٿ����]����Am���3��5�/�̾{`���}�o�R�Xy7��'�a� � U"��,�T?��}^�!���)	��X�ܾ����EA��[}��O���Ŀ;�߿/�����*տDy��8���k��
B��:0�l<7�IsV��Z��?u���Vȿ��⿄������ҿ��������bP\�$'��@���¾\�����{�R�V���?�OW3�*`/���3��,@��V�ݹz��a��k���{����#�`]W������֮�Uп���m���̿����%��?^�֩<��3��OB�w
i��|��.���F	Կq꿋��6��\ʿ�ʧ��鄿X�L�v��Dj�sO���K��6|�ã\��I���?�U�>��E�kFU�=�o�aq�� ����׾�����6���n�ט�i.���ۿ�E�O�>��b�ÿ�p���~���S��9�ٶ7���N�A�|�����k���H�ݿL��Gￛ�ݿ�п�����ru��<��i�9ݾj���MɎ���r�PSW��G��?��@�w�I�ʑ\��"{�i���ҷ��%�2h�1�G�t���䙤��Oǿ#㿵 �{��1.ؿ����K���q�<H�U,6��=�6A\��5��$C���˿b��T���}�'!տ�-����a�],�����̾�棾eꇾ4�j�dS�zUF���A�ŒE��Q��h�����M���
Ⱦ�  �  *��io���L�Ä��L��D�ſ��ܿL=係�ڿ��¿������R��H2��)� �7���\�鉿�j��H%ɿ�_޿�#�m�ؿW���^���<�{��@A�����޾\���z����b�T%C��[/��%�VX#�M�)�cF9�vkS�B�{�Ѧ��Ϳƾi��T1+��`�f�������ϿJB�;8��XԿ��fG��+�s���E���,���+���A�֙m������\��<�ѿMH�O>���ѿ<&��������f�PB0�<��|̾
R���[��\�V���;���+���$��k&�n[0� �C��b�=���f����i۾Ū�x=�Zv�;�����
~׿;�俌���3Ϳ�6��ɘ���wd��D=��2,���2�Y�P�ic���򠿬.��Grڿ������ʿD򫿼U����V��@$����R�¾����L���I[��GD�k�7�]u3�?�7��{D��<[�A�~� ʙ�%�������� ��VR��������ȿ�B߿.�濾�ݿ)�ſॿ���iX�vA8�/�Z�=�g�b������� b̿G���y�`#ܿE�¿Da���;���!H��z�����Һ��㗾]$��ta���M�c#D�q�B���I�S�Y�]t�zP���5��C[׾O
��3���h��7��tǵ��&ӿ0U忄F�cؿN���@K��J�{�A�M�R�4��3�:�I���u�Ġ���^��n�տoO��H�r�տ�8��eƗ��"o��v8�����tܾ����`����!w��[�TEK���C��D��8N�:�`�lW�A���Z}���辸_�G�C���|��b��tW����ڿ���A��]п�U������ʋj�qGC��$2�f�8�Y�V�9>������1�ÿ�"ݿr}近��+wͿ*���)���3\��y)�ϯ��̾)5��Qቾ�"o�Q�W��J�|�E�G�I��V�cl�_��������7Ⱦ�  �  �����G�?�V�s�����Z���ſK�˿�lÿ�׮�o���o�GJB�P�%�����*��!K�Z{��ؙ�T��Րƿ��˿$���	F���t��wh���5��*���ܾn���M��{�p��FQ���<���1�f0�t�6�7(G�W�a�W���'��y%Ǿ���0�"�0�P������s�������ɿ߾ʿ�����c���,��}Y_��-7�!G!�� �;3�RZ�� ��O��������ɿQ�ɿi���-h��b͆��IV�>'������˾�w��8����e�=�I���8��1��#3���=�ɵQ�e�p��������a�پ:�
��e2���c����I������N̿�ȿu����"��恿WR�Q�/�h� ���&��.A�9�l��ߑ�o����nÿ19Ϳ�Oȿ|3��e͛�~��I�(�6��ľ���n���V�i�� R���D��!@��D�R�Pli�n.���&���0¾��� W�)9E�Coy�@l���a��@�ǿ�RοJ2ƿ:���QK���Ou��/H�.�+���#�ȷ0�TQ�Ҁ��
��0���E�ɿi�οA0ſ����ߓ���n���<�s�����ѽ���� ���;o�	[[��
Q��O�t
W�<�g��.��yՔ������׾Q����*��#Y�@އ����������'Ϳh�ο¿�j���0���\g��-?��D)�(�i�;�0b�� ��Q�����W�Ϳ;�Ϳ/˿��z���㊿�{^��:/���	��;ܾг��������i�~X���P���Q�@�[�	o�����׷���廾vk�P���9��gj��j��0����Ŀ_Ͽs̿^"��D��O����nX���5���&��,�3�F�l�r����Xq���ƿ�ϿG�ʿ|̸�;f��r���0<N�XF"��P �"wξ�O������AY}�8qe�5�W���R���V�O�c���z����s\��Dʾ�  �  D��f ���/���W��������y2��2�����lm����{�vlO�a�*�����0�U���$2���X�*Ⴟ��O������Ϣ�1t��oz���N�>�'�T"��޾� ��a?��aT��+�k��_U���H�זF���N���`�f+}���������<�̾������=��g��{������'V���p���`���Ҍ���l�y�B�3"�(�3/�&9�
E>�"�g��a�������Ũ�"6��a���n�k��0A��u������о|^��T'���L��+�c���P��H�o�I���U��l��,��Ǜ������ܾ���!�%��L�9Uw�5'��jM��"̪����uԚ���*&`��o8����?��%���*�/�M�O�y��撿H���㿫��&��l���R��V�`���7�
i�����&�˾+���N���b���Ek��[���V��[�kk�"?�����R���vLʾ���I���#5��r]�粄�<���맿vҬ�K^��y<�������9U�Y�0�����>�D��F^8��C_�%��O���i���u��q3���ܕ�E�����U���.�>�$���7Ǿ������s��@t��h��Kf�]�n����E ��4~������ݾ���n!�fYE�[o�/���$����i�����[k��ڐ���t���J�>*��%��+��5'�%CF���o�d��7���Yͬ�r���`E���Ǐ���s�dI�1�$��@�85ᾂ���pr���y��1ԁ��_p��<g��mh�L�s����N����੾��ž�~�5Q��b,�R�R���}�_r��~������uV��0��`���hYf�g�>�v�"�v2�H��j0���S��Y�4���Ϊ���b�� ê����눿V�e��<����5��}�վ�j���h���N��ж~���n�_&i��m��|��֊��j��$ȳ�LaҾ�  �  ���d>��&#��!>�(F[�/Mv�'���hp��'X���l�L�L�,�������9�������33��{T�;s�K?������{/��q�6&U�<8�@�`0�4h��QξTm����������{��k��h��s�Gt���0E���¾��޾	�����c\,��`H�}be��h~�h���↿d�~��;c��5B��~"�|�	�Ϗ��$����ND��k>�_�_��{��S������:���8h�jZK�Y/�T9����ږ�<ž�n���h�������ku��j��*l��v{�1K����������;��ێ�����6���S��o��.���s������Hx��aZ� )9�Ha�S;�����	� � �U�+�^uL�	�l�~��1��&5��ú|��Rb�#0E�e�)�g�����f�޾^�þ�z���ј������y�1�x�9�g/���d�����oþ5_޾���0��ڡ(�b�C�Y�`���{�z`��r-��,���kr���R���1�w�� �\���\�uJ�n�9��Z��y�O���R������:�w���[��?���$�g!�q����ܾ��¾)ᬾ�����3��
{���C��E���[C�������׺��@Ӿvg�@F��Z���4��P���m��M���Ɋ�k񊿯Q���Jk�2>J�h�*�����E� �����B'��lF�/�g����)\��~��jJ��p`p�B�S�o=7��r��	��
�1zվ5Ƽ�
���X���c���!����|���֌�N��S(��-%¾R�۾sK��!H�s�#�z=��@Z�ٖv� y������\@��<�~�v�`��c?���!�"F����ǈ����Ll1�lR��er�MÅ�2����Љ�V����g��eJ�g/�_�����=龕ξ�������E��>�����ؓ��K��� ���y���˾v��  �  ���f�6| ���-�:[<���I��6R���R���I���8���!�p
��|�)Ծ��̾%iؾ�^������:'��+=�M�)�S�*Q�s9G��9��9+����K����y���d~ܾ�¾kw������k�b勾X��"����6���:Ѿ�������h�f��bn%��S3�z�A��M��T�n�Q��E�E�1��Z������mkо�UϾ���1g����4/�$�C���P�bT�p�N�j�B�{�4�+�&�"��_�;��dI�W�Ӿ�������d��������]��0���p���w�۾�����2���a�Ed+�J�9�X�G��/R�^�U��7P�,aA��,��v��h��ྕ�Ҿ�%ؾ���~%��v"���9�K�K�rV��{V��N�*�A��d3�^�%�����2���B�v�Ҿ�f���+��𤘾z����!��TG���`����Ѿn��H���f�R����%��l3�O�A��O�ҩW�raX�Y�O��>���'� 8�_?��B྆�ؾ���?� �|��ռ-�K�C�ŶS�ĕZ�h�W�<N��]@�!2�x%�u=�&���P뾱�Ѿ�����x�������꛾�V�����<�Ⱦ�ᾟ����+
�,���E!�[�-�j�;���I�+�U�.\�ݬY���M�d�9��c"��������g��O߾����e	�a��a97�ǍK�+�X�\�,�V�8K���<�<�.�41"�̝���Ⱦ�� ���ʾ�ȴ�2���w`��p�������c���uо��I��Y���K�H%�D2�}C@�h5N���X��j\���V���G��b2�"��\�� 쾨�޾N��c��J��b�'��?��RQ��R[�ݲ[�3�S��F�"�8�++�Y���i�Ϸ�7�����ܾ}Pľ�⯾�&������3��� ���¾�9ھ���8���  �  &���*��W,�vu,�!{,�[^,���*�b�%��Y����Q���r۾�迾�0�����(0��Awž��������W�'���+�k�,�7�,�g�,�u�,��*�B�$���I��`���׾׼�]�����Gk���rʾ���#�2��r!�k�(��>,��-�-��-��,�%*��#�m����	����XҾɛ���Ы�J���i���Ͼ�0����v���"��s)�M,�4�,�4�,���,��,�_
)��!������쾧G;5U���ݪ�����Ig����ԾR����|��n%���+��$.�1�.���.�-�.���-��*�,6"�����{���;;�������ֶ��HnþZ^޾�2��kE�T��W�(�L,.��0��S0�P0�2F0��/�J�*�f$"�n
�������*V̾��kɱ�?����ʾ��� �����8"�q�+�(Q0���1�g�1�F�1���1��90�rP+���!��%�l��8��
�˾�(��7��D���@ҾŎ�������%�FX.��w2�z�3�j�3�2�3��3�!�1�&�+�[�!����G)�M澞o̾���=����ľ5�ھAS��yz��/�sx)��%1�-�4��b5�'V5��V5��4��N2�<�+��� �V�����a⾂�ɾ�ͻ�7��:eǾ�߾14���������*���1��n4�L 5�?�4�� 5�8\4��L1�?%*�e\����yf��$�ݾlƾQ����A��'�ʾN��<�����ov!��E,��o2���4��05�,5�-25��K4��0�|�(��@��v��v����پ�.ľ�����f����ξ��}�t��+�#�x�-�%c3��L5�Z�5�i�5��5��H4�b0��Q'�h(�9
�y��־�r¾������ |Ӿ%��N�����G&��  �  ~�R��Q���H���;�0-�9������q��C��N�Fgƾ�m��+񚾅���񊾏����䞾����XY̾)�f��}<�o����"���0��?�d�K�wOS�%rR���G��P5��.�1!���-GҾQξH�ܾ�9�����tm+�w�@�[O��DT�R0P��ZE�X7�>+)��J�����!�
򾘂ؾn���7��hȖ�; ��!���<9��٥�E,���jվD�ʨ�!"�����f'�&r5�1�C�I�N���S���O��SB�#�-�� ��" ��`߾��ξ2IѾ>��V�IQ��3��qG��#S�I4U�W�N��VB��4��8&�q���_����!��Ӿ�޺�Sɥ�4���S���'q���<��<[��ZCʾ�)�J���A�
��S�?"��w/�`�=��kK�mU�&JW��P���?���)��N�����X�߾^�վO3޾����~��(���>���O�jlX�FLW��[N��A�7�2��J%��N�-���'��F뾠�Ѿ���ֱ��q���&�����:�������lzپ|�H� 	�ʋ���)��7�e�E���R��AZ�{}Y��"O���<��%��������G��J޾�,�e�����3��I�{W�ˣ\��X���M�9�?��j1�x$�:���B�W"�����!ϾA���ʦ��������5���׵��0̾_w���|���<���"��/���=�:�K��/W��/\�aX�L�J��5��Y��N����Y�޾��=�������#��;�:sN���Y�U�[��@U���H�{�:���,�Vp ����\	����uM�ytǾ�'���#���|��/��w�������S@վ����)�z�h��yr'�A�4��C�,�P�7OZ�)�\��2U��D���.�@����+U���޾JQ��� ����X,���B�bT��  �  m��N<��$�t�ŤY�{�<�3�!��0��:�mOҾ�̷�|ᠾ����!#~��l�#�f��/o�=���ԑ�����_����.پ�_���!���'��JC��o`�o�z��х�1P����H6h�1�G�zJ'��4��1���Y��;�������8�$FZ�:�w��~�������灿�l�=�P��3�_��%��l�ʾ�ǰ����0���x��j���i�L3v�`��̧��������ƾ���7����D�0��L���i�������F�6Rz�;�]��W<����Ȟ��W�����85��~$�ȦD���e��a��o���=!���~�ELe��CH�m,��[�]� ��^��ľ@���n��a��|2{�r��ev��ك�"9���;�����X־R�����7�"�qB=��BZ�wv��c��q��ʫ��|~u�U�V��p5�u���q����V7����%�2�ͶS�w|s��l��$������mbz��_�[	B�[G'�I���0���Zݾ#�¾l8���=��YҊ�r��nc�������NǞ�����˾����}�N��b�.��#J�7Jg������J��'׊����R�o��:O�^/�$!�Ψ�K����� #��JA�U�b�w%��n�������^��YNu�O�X��<���"��P�����Iھ�������:��GD���@���؄����_��謨�����־@��G�
�r��x�8��)U�3�q�aք�Z>��	���N����e���D�:�%����;�+�����,�hL��l�i惿���8���7����k���N��3�4����u�B�Ѿm���	��Ĕ���������s݆�8F��6i��R3����ƾ��྅b������(��wB��{_��?{����O��DA��d�z�l�[�f_:�ޡ�:2
�X�������4�6�F�W�<�w��w���  �  ���r���u��O���C�U���-����b徚彾�ӟ�Q㈾�Zo��W�B�H���D��WK�0�[��v�𾍾W0��q1ƾ;�-��"R6���_�ʅ�ի��A󦿆���4����<���Yt���H�i&������b��18�x�`�3����ߚ�˯��ȩ������A��\s��>H�c"�3���ؾ1��,|��熃��h�!�R�XH�3sG�p#Q��d��`�������I���:Ӿz� ��`��rC��$n�2ь�;���[ ��O�������	���%e���;�x�������a�#�\E���o��_��*����C��ޙ���_���	���)f��g<�����a��v0ξ*d���m��.���ph�=�V��P�X�S�u9a���x��f���飾^R��N��$�gk-���T�e8��jI��7B��E���ic������Y�����Z�'v4����L��{C��Q1���V�-����
���զ�����L��3���{��{[��3�	�=Y�r�Ⱦ�����9��]6��w�n�P�`�o]�~Rd�ju�Q>���W���Z�Ӿ$���vg��)=��df��6����Yl���~��qF���򓿸�{���P��d.�n�M��#�_�@���h�,􊿉��k㫿����!�
l����{��~P���*�����Y�P3ľ�����������ys�<h��kg�q��x��ef��װ��dc��b����&���K�bZv�,�����E��lv�������0��qom�:D���%�b����j{+�*�L��{w�����6�����L���!����X��1�l�mC��|��F�ZH۾z]��>��\9���n���Ho�t�g�A�j�Hx�Ψ��[��ମ�o�˾�M��Q�G�2���Y��Ԃ�|痿৿�������+��<��	�_�iK9�Ӵ��+�]����5���Z�᥃�D#��U⨿�  �  ��˿�/Ŀ�G�������p�i'=�O��k��r��-C��|v��[T�26>���1�(w.�(�3��B�2[�w��$A��m(���I�Ԭ��9H�U�}����������Eǿ�i˿������S׎�)]g���<��o#����3/���R��_��Ƴ���@��T�ȿ�˿�����%���zV_�͂.�ە�k�Ծ�ͩ��:��]Ik�ɥM���:�Z1���0�^&9�>�J�gg�|5�����̴ξG���q)��2Y��b���ि�ü��2ʿ_ɿ�s��¡���M��)@W���1��q��!�j9��Hb�c����<���}��5�˿�6ɿ���ϣ���炿&�O���!�����>�ǾEӡ�����3�g�ekN�@`?�R�9�v�<�"�H�1^�������>���O澂����;�r�n��Γ�?r���yĿ<pͿ	�ǿ�괿:���j|��M���-��"�0~+�I�$w��w�������ƿm?ο��ƿj��eԗ��[v�>�B��U�������o��;Z���mk�C�U��I���F�|�L��\�~+u�.��������̾������"�O�&G��@���1��ɾʿ&�ο�Ŀ�x������:o���D��+�_'��`7���Z�����x颿zv����̿�8Ͽ�9ÿ3���叿�g�θ6�t�����)����\��������m���Z�~WQ���P�� Y���j�G���2D��5�����޾"��U�1�H`a�~��  ������5Yο~�Ϳ1���&˥��u���_�c#:�ؚ'���)�o�@��j��y嫿
ÿ!Ͽo�̿�b�� �74���*V���(����վ^ͮ�����iz���9g�K�W��^Q��S�$b_�u�t��u��١���¾u������@���s�Uk��+��$ǿ�
п�Jʿ�t��M���~�����Q�v_2��&�0��M�N�{�5���Oٴ�M�ȿ�  �  t3�)�ۿ2CĿ~k������j�I�]#��|辘'��ƍ�kOh��+F���0��$�0�!�\�&���4���L�1�r��J���彾x��3#���V��j�����̤ʿ�(߿V�R�׿S���4���s�|���K�}k/��*�J�<���d��J�������Ϳ@����,�տ]����r��iq�3�8��#���վ2������8]�+�?��q-��$��$�8�+���<���X�\큾1���I@Ͼ���	3��Qj������඿��ҿR����Eп{o��D���fj���?�#�*�b�-�Q�G�N�v��P��1 ���ֿ$��L῎^οF�������F�^��#*��m��>ǾU)���.��
Y�!�@��C2���,���/��;��P�.q�a��M|����込9�դG��O��;����¿C�ۿ	�gi߿�ɿ����{9���)^��o:�oI-���7���Y�:#��I��5�ƿAD޿`�濴O޿� ǿ�(������@PO���&t�94���򘾹�~�]>]��"H��<��J:���?��MN���f�����d���Xk˾���k*�Eu]�UՍ��y��ο��⿖��Ahۿ���↡�w^���T���7�h2��D��dm�r���h;��!�ѿ��7��ۯٿƶ��"���©y�MA��O�� ��c���?���b}�I�_�(yM���D��D���K�t�\���x�Z��������h߾��~.;�6r�ݥ��n ��a ׿���忧oԿ0����ؖ���r� H�W3���5���O���~���������ٿ4����C�ѿ峿�I��se�Q�0�D��VԾ�#��� ���r��aY���J���D��G�z�Q�p^f�ԇ��O!�����}�8p�v�L�}ꃿ~4��ſ�3޿ڮ�F��I̿�������j�b��.?���1�ۖ<�4^��Z��`s���ɿ�S��  �  �3�wp,��4��R��fS��.Ɏ�7�P��@�1J�P��5\��K�o�.�S��E��A��G�5Y�ix�S'���G��l��18$��1`������̿�,�k���t/���3��)�
���7�÷���.bo�L�f��S��Ȱ��wԿ�s��7 ���0��63��'�(��+D�v���9��?�<��C�E�Ҿyؤ�إ����f��PO��D��|C��\M�.�b�3Ճ������.̾͜��
6��x��,����߿���
�$�cs2���1���"��t	�}Wڿ?�������h��_l��q������h#�@���C'���3�g1�>� ������ӿS,����i��+�Q	 ��ľ�ݜ��*ge��S�L�c�O�G�]���x�����n�������iM��ڋ��?�������Z��+���4���.�]����yʿq�����~�O�i�Y�z�/���ſ�%��7z���-��A5���-�������ÿ�����CV�ú��S�~9��屙��]��yik�y]���Y�ޙ`�}�r��B���m��{�Ⱦ���+��g��w��2пn���b��11�Im5���*����#&�Vλ����]�w�So��������,�ؿ��Y"�u�2��T5��()����mq��!���"����D��p�$��X���̖��_��txo��;d��c�.wm�a����쓾ٲ��.\ܾ���1>�B���?J����;����&�W�4�L�3���$�f���޿'u���,��\p�ܢt�x���������a��W)�B=5�h�2��B"�{n��4׿r|��M�p��]2�����Ѿ���������N~��zk���c���f���t��{��1����,���1�B$�~�R��t�� ۾�?h������-��6�G0��7��L��̿_��}����-n��?����N=ǿ�S�������.��  �  �f,�GK%������I蹿>튿[�L����0j��Ⲿ����Du�CaY�)VJ��KF��L���^�$�}�£���Ҽ����CI"� �[�����ƴſBE��vC�+(�H+,�D"�P��Xm俛����Њ��Ai��a���}�(�����̿,B�߹��`)�Ŀ+��- ���	���ݿ1{����{� �9�Ee
��]Ӿ)��n\��%l���T��bI�ݾH�q�R�-�h�В���Ԣ��4;���R3�is�����ȝ׿h�}�j+��<*���a��~ҿ㢿�M��8b��cf��z��̶��W�޿�)
��n ��,�0�)���0��ԁ̿�����d�7�)�VY����ž�H��`�����j�sX�<]Q�N�T��Qc��C~������a�����9����I�=���$��ӷ�^�.�$�YM-���'�����^��J�ÿ���rx�X�c��/t�o;��(X�����@b���&���-��&�ks�Ȩ��������LR��A�es�����J���,��Z�p��ab�v�^�%�e�sGx�G���餾RHʾ�� ��!)��ab����H"ɿJ������x�)���-���#�7���Y�H���w��q���i�����Ң�I0ѿ:d�����+���-��I"�D�⿔���������A����T���7��+���N.��!�t��i���h���r��]��
���b����aݾ[
��y;��={����ۿ		�d! �L-�'V,�� ��6�h�ֿP����o�j�]�n�Q���鯰�������:"�;�-�`+����9���ϿU؝�o�k��.0�wB��Ҿ�+��ih��񁾅�p�$=i�=l��#z�qK���������S��m���N��֊�)����U����%�>�.��)�b��������ſ�j���|��h���x�r���	�������4q�=�'��  �  ���������ֿ騿e怿C����6��6��ߙ��փ���j�Y�Z�"�V���]�up�D:���P���%þ���j�6�O�7=��%���oE����s�0���A�e����̿�꠿��~�O*X��Q�8�i�ww��>]���O�k���C��a��m���{ǿh����{k���2�R	� �׾0�����_Z~�x�e���Y��Y��c�s�z��M����(Ҿ[$�U�,�<d�_H���&¿7W� ������;�*�	��*�` ���/��]<n��R��U�(y�����ǿ������k�����u�J<�gܸ�}_���X�j�$�������˾�Χ����|��Qi�(�a�vge�۾t��M��۰��:��� 1�K��@���}�� ���zӿ�C �������G����ݿ'������h�e�a�S��=b�)Շ��'��8ٿ����Y�\m��X����RٿY���8����H��R��� ž�5���`��G=��W�r��o��v�g���E��>�����о<T�E�$���V�l���c��۲�T���0���������zlп;��z���}`��xY��Vr�i��������P=
�Ң�H��C��ܟ���˿�%��Ⱦs���:��K����!��-����H�������y��/y������l��ٟ�����U�yB� 5��6l��e���HƿB~�����n���T�Y��_�&U��b��>�v�ZQZ���]�����ǧ��{˿�V��ʮ����~�X 
�	�꿿+�� ���p�^��L+�a���ؾn���e���d劾�ۀ�p�y���|��Ʌ��x������%Ǿ���`���F��y��뛨��ֿ���6��!I������\�5��cz��%Yj��X���f���`���Eۿ���[`��  �  ��G�￹׿��������`i���8�Nr�����ʾ�,��5���=���w�x���s���{�_Έ��3���|����Ҿ����%��%�B�N.v�в������J�ݿ���e����O뿥Ͽ-���T����H^��k?�w�9�Z�M��ay�����Ŀ��@࿍��3R���`��̿�3��X����gX��$,�4����m���ʤ��p�������w��Kv�+����u������ֳ���'ྼ����'�X�R� ���$��%�ȿ��濟O��? ��}�&ÿP����5�?Q�i|:�!w=��Y�=e������˿
V�6����������"M¿�\���i~�e�I���!�����۾B߹�b
���4��H�Э~�7����k���ޙ�� ����;����.��P"8�,g�SV��&���ږտ&�����_���ۿ����R��J�q�k K���<�YH���l�h�0����ؿ�6�{���ݞ�F�ٿ`���Ε� �n�.q>����+�����վ������^w���f��k��G}��B����;��뽿�KMྃ��T�"�R�I��}�r!������I῜&��8N��1����ҿ���<����if���G��B�`V��퀿�C��	Ŀ\��8J��č��\��ѿa���Ì���`�\4��7��Z��%�о(�!����ǒ������1��Ӎ������n����̾�T����/�O�Z�m���F���Ϳ��&~��uQ��?E��ǿ�䣿)Ƀ�iY�-�B�țE��a��N��Ы��nϿ����G���G���忒�ſ
���E���mP�&(�):
�m辇�ƾ�������P$��DG��:3��%ؕ����x���Qlؾq�������W=��_l���[A��j7ؿ�]�e���I��R޿y���Ř�Awv���O�{A�s�L�q�2'��&-��+�ڿ�A���  �  ���}F��V��=����k~�!�V��6�:��=�Z��:_̾Ҳ�}Y��LW���揾�`��;���=���Ӿ�����J�!��<��"_��<���䚿�ů�h���_x��A����d��n#���a��:�O%#���W�-�hN�T�{����,���袽�����8=��ʤ�ZZ����p�F|K�Y-��R�y��o;�@4ľ�|��!L��G���%y��Wƙ����1��U�ݾz�������-*�уG��$l�騋�=7��w[����/e��d������Ox��UR�(S0��y���!���6�:v\�t����,���M�����Pm��퓲�]<��0���&e��'B��H&���̔����ھQv��r
��0��������E��𰣾̶��K�ϾUH��=a�#�6�neV��~}��
���
��l廿��¿���ū������yt�mI��,��8"�<�*�,�E���o�u/���⩿�5���tÿ������{g��n򁿿\���;�β!����� ���׾�]������Y���(���⡾�����>ž,Hྍ ���y�(�%�C�f������S���7��;��uĿH,�����K���~�h��*B��V+��*'�G"6�Y�V����"����岿U�����Ŀ t������1����Fy���S��5��~�Ϋ	�o��YԾ^���_����ń���ҩ�M(��8/Ѿã�+u����S2�I�O��]t�`ʏ�G]�������Ŀ¿�ʹ��L��������Z��8�}�'��)�d�>��3d�@[���ӣ�ظ�DĿ��¿�鵿Ѝ��G㊿d�k���H���,�V������p�V̾�x��oҧ�#q������!������ �ھ6��Z��"�k�;�[�{Z��⨗�D���D����Uſ����LS������ey��AN���1��&�zw/��UJ�v-t��R�����r>���  �  �V��ꏿ�����{�X0f��R��B�M�2�Ħ"�ˆ������߾)yľ񝳾߼���u����ɾ�.�y�������&�NM6��E�J,W�^<k������������䐿D7���v��1T�a2��E�0�(�n���B%���D���g�ߵ���u�������K��8���*u���_���M��t=���-����O%��r�� 8־!z��c������_��:Ӿ2��4
�2����+��;�8kK�4}]�br��'�� T�����\��+��o>k�4MH�|*(��f�H���3�-)�6m/��P��s�)�������(�����𮂿Yo���Z��I���9��8*�/����QEdѾ�1���h���2��Ⱦ��-[��	��d$���4�VD���T�b�g�V}��\���I������V��OC��ՠc���@��%#���E������ �b�=���`�l*�����P��k���wA��0���B�k�qAX���G�w8��*(���Ξ�@���?о,���H�����¾�־%󾊏
�_L��L-��%=���L��^��r�����0��܉��m��9ӌ��}���[��,:��=��7�P������-�q5M��=p�,�r���b5���Ӱ��փ}�`Ih���U�a�E��6���%��>����8R澀�ξgp��:����k̾L��� �����#��4���C���S���e�=�z��L���|���ᕿ�5���2����s�	�P�Po0�G�����,0�����7�,sX�#{��
��Ƈ��숕�u֏����]�u�ʥa��'P�px@���0�u ��w����p�ݾ_ɾ�X����þ��ӾHO�4��-n��)���9�:SI�0�Y���l��H������c꓿="��9�҄�S�h���E���'�����N�9a�_E%��VB�p�d��<������  �  �.^��d��5e���d���d��Ee���c���]���P��@=�:�%��������ݾ'�־��5N��V���g+�~8B�0}T�d�_���d�шe�fe��<e�Ğe���c�ny\�MBN�L�9�%I"��d����۾��׾�6�j�����v�/���E��-W��xa��oe���e��Ae���e���e�%c�O�Z�gK�r96��r�:
�Lb�**ھ�پV������w�3�Q"I��;Y�Qb��ge�tTe���d�-Le�~8e���a��MX�|�G���1��2��w���� �ؾ�ھ�z�R�	�.j ��Y8��wM�1�\��d�3g���f�_�f�-:g���f�0�b�kX���F�C40�p��,���x��iܾ���k���g���&�<=>�EvR�Yc`�'Vg��i�D�h�'�h��i�Ah��c��KW���D���-�my�O�|i��]߾���d� ����A,�F�C�L�V�{�c�[�i���j��:j��?j���j�>ii��Cc��GV���B���+�@q�.����%��<h�2}��/�	�1�Q�H�XB[���f���k�-ll���k� l�)�l���j���c�sU��<A��)�z�� �w쾇6�ؾ����
�>C ��8�lfN���_���i���m�hn�}�m�Y�m��n�[k�w�b�m�S�mR>���&��t���6�%�7a��%����#�E�;�.7Q��Wa��uj���m���m�,m���m�·m��#j�ɣ`�]%P�fI:��x"�H��;������&�������4���'�|�?�]zT� ~c��}k���m���m�jcm�$�m���m��Di��^��M���6������	�����Y�_��F�z�k,�C�C���W�#�e���l�9Fn�@�m���m�JLn�l�m�#Vh�a}\��I���2�Cm�~)�s��M�辕��~V�9�vz0��G���Z��  �  �Y3�h�B��S�\Ug��4}����/8��GD��ъ���{��Y��[7����-���O�ޞ��q ���>���a�"3������ʑ�D6�����\�x�Sc�+8P�q�?��`0��8 ����'���8�ھ����𕲾�˯�)�����ξE$��0�s���})�\$9���H�~�Z�wo�q���p?��񢑿�8��QY���Bq�wxN�F_-�v����������*��~J�	hm�o������B���B�������P-q��Z\�waJ�-~:�\�*��]�n��X��BѾ`Q���y���+��9��$�ؾ|���������	0��?�K�O���b���w�|І�"l��yƒ�Uގ��Ѓ��g�[�D���%�K��1I�2
��.���6��Y�sr{�!p���Ò�ޏ��(�������m���Y�~�H�9�MB)��_�,���i�1�о�A��Z���;b���&Ͼ,|�j����Y�(�=�8��bH��>Y��l��T��Ƌ�c�	 ����������n_�k(=�A� ���uh	������&��9E�Q9h�ㅄ�~^���3�����H������j��!W�z�F�ml7��c'��@�����꾢6Ѿ��¾����A�ɾ2߾,���@��4!�q�1���A�NQ�[�b��hw�?����_������'N���i��[y�,�V��k5���޿���W���2���R�Kvu��ꉿˍ��2Ε���������ky�%�d���R�o�B�`<3�"�"��%�������ᾛy˾Ai�������Ͼ�����J*�͑&���6��cF���V��2i��~��#��:������(%��v��3n��'K��	,���@����� ���<�m�^��o������c���)��D��� Z����r���^���M��A>��t.�f��Z��8V��ppھA�Ǿ���sƾ:�׾��
�����,��  �  �c�s�7�ًX�#g���s��p﻿�����ظ�����G���ah�6F?�e%�d��)�)�AUG��%s�U��`���Ļ�r����l��)��	����w�C�P�ɱ1�����o��8�lȾmɯ� t���͒��֐��]㦾����ؾ���xq��&��bB�+�e����Q���MԲ��+���Ŀ��޳��t��<ꄿW�Y�,5��*!�� ��2���T���V����̱�U�
���h���?���i��m�i�$�E�͘(��i��f���v۾d��Xר�����~���Ȓ��ܜ��ʮ�{0Ǿ�����A��-0�o�N�V�t�W[������θ�����V��m��5��:�z�GN��.��� ��v&���>��Uf�����;��
���P¿��xy��%a��Ä���`���>���#�ZX��^���$پJ⾾X����c������𜾏����׽�x�׾��h��v�"�W=��	^��#��J����*��?����vÿ���樿�#���2n�g/E��d+���#�-�/���M�k�y��U���`�����&EĿGټ�8���jz����~��W�e�8�*�����z���pN׾P�����������FW��tc����;�U�s��\���.���J�1.n�M<���⢿�󶿻Eÿl�ÿ�������q�a�R4=��0)�K(��:�	�\����0���wֵ���¿{�ÿF����&�������#r���M�Y�0����{���!�Ͼ���-'���P���T��e��������վ*�f�
������6�huU�%^{����O
��5���Ŀ�3������6������77T���4�P�&�W,��QD�0l�ю�b���ȭ����Ŀ����(������`^����e��
D��4)�����R��C㾐�Ⱦ�=���妾w������������oƾ�\�4J��]���  �  F��A;��bl��甿ʖ����ؿ��Q��0��$VԿ�������`e���B��8��?H�8Hp��)��9���eKۿ���Z����쿸ҿ��΍�4�`�%{2������h�žJ���!�� Y��Cx��Iu�Q��#݋�MZ��i۷���پ�t�8�!�V�J�������(yÿv��3������n���ɿKХ�������W���<��N;�+]S��Y��Rӡ��ſǮ俫���<����B忱ǿ39���H����O�d�%��:�ݾu���F����|�������v���x�	3��>�������ľ7��=����/���\�[���嬿�dϿh뿿r���,��{�߿�ľ��#����x��)N�ʾ;�O�B�AOc�����*���mҿ2�������*�ݿh�������v�� D�j���8��KؾP������H����
���G䅾{���/g�������־���G��6�@�a�q�;���P����ۿƛ����qW�\'׿�n�������Lk�ˉH�v�>��dN���v�hS��G༿��޿�����V���F𿿄տ�a���?��B�g��o9����:3���Ծ�g��xB���ɓ��݋�����,��QJ��3��Ⱦ�꾅��LN*�=S��G��˰��ѝǿ�������u����뿤�Ϳ�ة�}�����_���D�6SC��a[��\���ץ���ɿ*�迌���, ��=X�i7˿W��@j���X���-��]��(˾�ذ������	��j
��ы�W���q���/���GҾ������K\6��Qc�{j��7���ҿ������k���������Q=���~�2T���A�V�H�%i����������*տ-���B��_)�����P ���+����{��=I�"�"�"k�/�⾔�¾����5�������ދ��쎾��������{���޾���  �  k����E�����X���Yٿ߳�������a�%t ��Կ|��ヿ* \�r�O��<c�0����밿{޿w�����������u���$Ͽ�㡿wv���:�&����߾r���C������>�h�Q�Z��7X��+a�v��9��ޥ��ʾT���x�%���Y�Rȏ�]������	�l��P�=����,�ĿU����Rv��T��	S�Dq�x_���п����g�
����i��K�
�3��𙿿y���o`�hC*��*��NϾ)�	^��ty��Hc��Y�{[�p�h��X��sr��_ǲ��ܾKP�a�6�:�p�
����ʿ���#��}'�v{�ې���信���ܯ���i�lS�k�[��1���}����п���U��}���������q��6��鈿�P�7\�Y���ZȾ�o��������qn�8h���m��%�(����l��qeƾ����_��{K�3���{��7ܿc����#t��������ֿ`i���چ�� b��U��[i��ٍ��������������ܦ�~����ҿIT���^}���A�:��}	�	�¾�	�����������
z�Fx������d��G���ރ��4�۾�I��-��Ib������ξ��+�*&���Z��������u�ȿ���bZ~���\�M[��y�pb��3�ÿN�����ů�������n�1�ÿ(��<�h��2�'o�i�߾�U������U���������x�A<z�Q���H��᣾������� �4N=��?w�\��d"ο����V~�{�����'	���翖������n p���X���a�5���[��cVӿsX �e)�+�R����	��Ѵ�m����[U���$�����Ҿi������䅉�K���\�z�^���\���/���ǭ���ξ�����  �  �#��@P��>���ż����Te� &��i,���$�����G��N��
����m���_���u�����GĿNf�����'�)J,���"�� ���g����E��-C�}���Bܾ>�7����p��_W�x9J�u�G��@P�pd�G��dn���)ž2�����*�.?g��P��!�ο�����<�)��{+�'7����Q�ۿv8��h�Yne��ac��肿�g��g�տ���-���*���*�����B�ԿQT��6�n��?0����jʾ�����2��sg��UR��`I��%K���W��p��\�����B�ؾu���&>�ٳ���﬿v��#��&�!�mj,��F)����F �#˿�}���]}��c��Em�1ڍ�����n��b��L�#�&-��b(����n�����Ŀ�����\[��:#��������<���vⅾT�m��L]���W�j:]��m�'k��ΐ�������\�!����U�I���1���*�������l'�c�-�~�%�Q8�b*��=�������s�o�e��|�R��;gǿ˓����1)� �-�T�$�2���W����!����J�}��m~�?f��*��������v�'{i�E�g�&�p��`��	������Z�վ�_��.3�՞o��}���ҿ	��+����+�i�-��>!�N�
���߿'>��B����sm��ek�놿�j����ٿǬ�����,�ƺ,�P���(�ؿbt��P)w���8������ھ���sp������Vr��h�N�i���u�`����Ú����y澪��h�D�S	���@�����	p�	0#��
.���*�͙�L���4ο����}�����h�4-s��Ő�Wr��˫�nN�(%�x.���)��0�Δ���ǿN�����`�u(�>��̾ҧ��ӏ�����"Np�=~j��Do���B���yꤾ��ǾAg���  �  G���cT�r:���Yÿ������@-�`�3�|�+�=������Lտ�4r���3t��Ke���|��Ɯ��_˿���'S�w�.�j�3���)�#
�k�￴���BŇ�S�F�>��۾몾����~Ok���Q���D���B���J��^��;��r��;�þ;p �w-���l�����Lֿ���&t!�<1�|�2�]�%��+�B��
󯿏։��_k�W:i�?���㪿v�ݿM��#�� 2��2�V�#�~�[�ܿ�c��u�t���2�T�ɾcl��!u��a~a��L�I'D�2�E��QR���j�����稾��׾����OA�����ݕ���>꿌���x(���3���0�Is��d��ҿ����+����h��ws���@ѻ����}��վ*���4�"�/��:�6s�%k˿w7����_�Z%�����J7��-�����Lh��W��R�R�W��h�v�������[���:^�1!���Y�=���ƿ�G��9���.�(H5�w	-��>�p���¿�k���4z�	Yk��k��۟��~ο�=�����j0��t5� �+�b���>�����<8���yM��"����zb��tJ��S����p��*d�irb��k��%�ɸ������C�Ծ����}5���t��D��nuڿ}
�J�#�tH3�I�4��(�M1�h�翵���cڍ��ds�>q�f����宿���g�V�%��&4� %4���%���#��σ���|�;����xwپ�Ȯ�ᯒ��̀���l�,Zc�<�d��Zp�@*����������`���H��M��t浿[��	3��*�΄5�6-2��!����l�տ�����+���n��_y�������������/��,���5���0����p��ο�Ԛ�Ne�_E*��(��~ʾ�M�������{�D�j�#Ae���i��y�+��X��*�ž�h���  �  �#��@P��>���ż����Te� &��i,���$�����G��N��
����m���_���u�����GĿNf�����'�)J,���"�� ���g����E��-C�}���Bܾ>�7����p��_W�x9J�u�G��@P�pd�G��dn���)ž2�����*�.?g��P��!�ο�����<�)��{+�'7����Q�ۿv8��h�Yne��ac��肿�g��g�տ���-���*���*�����B�ԿQT��6�n��?0����jʾ�����2��rg��UR��`I��%K���W� �p��\�����@�ؾt���&>�س���﬿u��#��%�!�mj,��F)����F �#˿�}���]}��c��Em�1ڍ�����o��b��M�#�&-��b(����n�����Ŀ�����\[��:#��������=���vⅾU�m��L]���W�j:]��m�&k��͐�������\� ����U�I���1���*�������l'�b�-�~�%�Q8�b*��=�������s�o�e��|�S��<gǿ̓����1)� �-�T�$�3���W����"����J�~��o~�@f��+��������v�({i�F�g�'�p��`��	������Z�վ�_��.3�՞o��}���ҿ	��+����+�i�-��>!�N�
���߿'>��B����sm��ek�놿�j����ٿǬ�����,�ƺ,�P���(�ؿbt��P)w���8������ھ���sp������Vr��h�N�i���u�`����Ú����y澪��h�D�S	���@�����	p�	0#��
.���*�͙�L���4ο����}�����h�4-s��Ő�Wr��˫�nN�(%�x.���)��0�Δ���ǿN�����`�u(�>��̾ҧ��ӏ�����"Np�=~j��Do���B���yꤾ��ǾAg���  �  k����E�����X���Yٿ߳�������a�%t ��Կ|��ヿ* \�r�O��<c�0����밿{޿w�����������u���$Ͽ�㡿wv���:�&����߾r���C������>�h�Q�Z��7X��+a�v��9��ޥ��ʾT���x�%���Y�Rȏ�]������	�l��P�=����,�ĿU����Rv��T��	S�Dq�x_���п����g�
����i��K�
�3��𙿿y���o`�hC*��*��NϾ)�^��sy��Hc��Y�{[�m�h��X��qr��\ǲ��ܾIP�_�6�8�p�
����ʿ���"��|'�v{�ڐ���信���ܯ���i�lS�l�[��1���}����п���V��~���������q��6��鈿�P�9\�\���ZȾ�o��������sn�8h���m��%�&����l��oeƾ�����_��{K�2���z��5ܿc����"t��������ֿ`i���چ�� b��U��[i��ٍ��������������ݦ������ҿJT���^}���A�<���	��¾�	�����������
z�Hx������d��G���ރ��5�۾�I��-��Ib������ξ��+�*&���Z��������u�ȿ���bZ~���\�M[��y�pb��3�ÿN�����ů�������n�1�ÿ(��<�h��2�'o�i�߾�U������U���������x�A<z�Q���H��᣾������� �4N=��?w�\��d"ο����V~�{�����'	���翖������n p���X���a�5���[��cVӿsX �e)�+�R����	��Ѵ�m����[U���$�����Ҿi������䅉�K���\�z�^���\���/���ǭ���ξ�����  �  F��A;��bl��甿ʖ����ؿ��Q��0��$VԿ�������`e���B��8��?H�8Hp��)��9���eKۿ���Z����쿸ҿ��΍�4�`�%{2������h�žJ���!�� Y��Cx��Iu�Q��#݋�MZ��i۷���پ�t�8�!�V�J�������(yÿv��3������n���ɿKХ�������W���<��N;�+]S��Y��Rӡ��ſǮ俫���<����B忱ǿ39���H����O�d�%��:�ݾt���F����|�������v���x�3��<�������ľ2��:����/���\�Y���嬿�dϿh뿽r���,��z�߿�ľ��#����x��)N�ʾ;�O�B�BOc�����*���mҿ3�������,�ݿ	h�������v�� D�m���8��KؾS������H�� ��
���F䅾y���-g�������־���D��3�@�]�q�9���P����ۿě����oW�Z'׿�n�������Lk�ˉH�v�>��dN���v�iS��H༿��޿�����V���F���տ�a���?��E�g��o9����?3���Ծ�g��{B���ɓ��݋�����,��QJ��4��Ⱦ�꾅��LN*�=S��G��˰��ѝǿ�������u����뿤�Ϳ�ة�}�����_���D�6SC��a[��\���ץ���ɿ*�迌���, ��=X�i7˿W��@j���X���-��]��(˾�ذ������	��j
��ы�W���q���/���GҾ������K\6��Qc�{j��7���ҿ������k���������Q=���~�2T���A�V�H�%i����������*տ-���B��_)�����P ���+����{��=I�"�"�"k�/�⾔�¾����5�������ދ��쎾��������{���޾���  �  �c�s�7�ًX�#g���s��p﻿�����ظ�����G���ah�6F?�e%�d��)�)�AUG��%s�U��`���Ļ�r����l��)��	����w�C�P�ɱ1�����o��8�lȾmɯ� t���͒��֐��]㦾����ؾ���xq��&��bB�+�e����Q���MԲ��+���Ŀ��޳��t��<ꄿW�Y�,5��*!�� ��2���T���V����̱�U�
���h���?���i��m�i�$�E�͘(��i��f���v۾d��Wר�����~���Ȓ��ܜ��ʮ�w0Ǿ�����>�� -0�k�N�R�t�U[������θ�����T��m��4��8�z�FN��.��� ��v&���>��Uf�����;�����P¿��zy��(a��Ä���`���>���#�]X��^���$پM⾾Z����c������𜾍����׽�u�׾���f��r�"�S=��	^��#��H����*��=����vÿ�����樿�#���2n�f/E��d+���#�-�/���M�m�y��U���`�����'EĿIټ�:���lz����~��W�i�8�.��Õ����uN׾S�����������HX��uc����;�U�s��\���.���J�1.n�M<���⢿�󶿻Eÿl�ÿ�������q�a�R4=��0)�K(��:�	�\����0���wֵ���¿{�ÿF����&�������#r���M�Y�0����{���!�Ͼ���-'���P���T��e��������վ*�f�
������6�huU�%^{����O
��5���Ŀ�3������6������77T���4�P�&�W,��QD�0l�ю�b���ȭ����Ŀ����(������`^����e��
D��4)�����R��C㾐�Ⱦ�=���妾w������������oƾ�\�4J��]���  �  �Y3�h�B��S�\Ug��4}����/8��GD��ъ���{��Y��[7����-���O�ޞ��q ���>���a�"3������ʑ�D6�����\�x�Sc�+8P�q�?��`0��8 ����'���8�ھ����𕲾�˯�)�����ξE$��0�s���})�\$9���H�~�Z�wo�q���p?��񢑿�8��QY���Bq�wxN�F_-�v����������*��~J�	hm�o������B���B�������P-q��Z\�waJ�-~:�\�*��]�n��X��BѾ_Q���y���+��9�� �ؾx��������	0��?�G�O���b���w�zІ� l��wƒ�Sގ��Ѓ��g�Y�D���%�K��1I�2
��.���6��Y�vr{�"p���Ò�Ꮢ�*�������Ǌm���Y���H�	9�QB)��_�.���i�3�о�A��Z���:b���&Ͼ)|�h����V�(�9�8��bH��>Y���l��T��Ƌ�a� ������	����n_�i(=�?� ���uh	������&��9E�S9h�兄��^���3�����K������j��!W��F�ql7��c'��@�����꾥6Ѿ��¾����B�ɾ2߾,���@��4!�q�1���A�NQ�Z�b��hw�?����_������'N���i��[y�,�V��k5���޿���W���2���R�Kvu��ꉿˍ��2Ε���������ky�%�d���R�o�B�`<3�"�"��%�������ᾛy˾Ai�������Ͼ�����J*�͑&���6��cF���V��2i��~��#��:������(%��v��3n��'K��	,���@����� ���<�m�^��o������c���)��D��� Z����r���^���M��A>��t.�f��Z��8V��ppھA�Ǿ���sƾ:�׾��
�����,��  �  �.^��d��5e���d���d��Ee���c���]���P��@=�:�%��������ݾ'�־��5N��V���g+�~8B�0}T�d�_���d�шe�fe��<e�Ğe���c�ny\�MBN�L�9�%I"��d����۾��׾�6�j�����v�/���E��-W��xa��oe���e��Ae���e���e�%c�O�Z�gK�r96��r�:
�Lb�**ھ�پV������x�3�Q"I��;Y�Qb��ge�uTe���d�-Le�~8e���a��MX�|�G���1��2��w������ؾ��ھ�z�P�	�+j ��Y8��wM�-�\��d�3g���f�Z�f�(:g���f�,�b�gX���F�A40�n��+���x��iܾ���m���g��&�?=>�IvR�]c`�+Vg��i�I�h�,�h��i�Ah��c��KW���D���-�oy�O�}i��]߾���c� ����A,�C�C�I�V�w�c�V�i���j��:j��?j�}�j�9ii��Cc��GV���B���+�>q�
.����%��>h�3}��/��1�T�H�[B[���f���k�2ll���k� l�.�l���j���c�sU��<A�	�)�|�� �y쾉6�ھ����
�?C ��8�lfN���_���i���m�hn�}�m�Y�m��n�[k�w�b�m�S�mR>���&��t���6�%�6a��%����#�E�;�.7Q��Wa��uj���m���m�,m���m�·m��#j�ɣ`�]%P�fI:��x"�H��;������&�������4���'�|�?�]zT� ~c��}k���m���m�jcm�$�m���m��Di��^��M���6������	�����Y�_��F�z�k,�C�C���W�#�e���l�9Fn�@�m���m�JLn�l�m�#Vh�a}\��I���2�Cm�~)�s��M�辕��~V�9�vz0��G���Z��  �  �V��ꏿ�����{�X0f��R��B�M�2�Ħ"�ˆ������߾)yľ񝳾߼���u����ɾ�.�y�������&�NM6��E�J,W�^<k������������䐿D7���v��1T�a2��E�0�(�n���B%���D���g�ߵ���u�������K��8���*u���_���M��t=���-����O%��r�� 8־!z��c������_��:Ӿ2��4
�2����+��;�9kK�4}]�br��'�� T�����\��+��o>k�4MH�|*(��f�G���3�+)�4m/���P��s�(�������(�������Xo���Z��I���9��8*�,����MEdѾ�1���h���2��Ⱦ��/[��	��d$���4�ZD���T�g�g�V}��\���I������V��QC��נc���@��%#���E������ �`�=���`�j*�����N��i���uA��-���=�k�lAX���G�s8��*(���˞�=���?о+���H�����¾�־�%󾌏
�aL��L-��%=���L��^��r�����0��މ��m��;ӌ� �}���[��,:��=��7�P������-�q5M��=p�,�r���b5���Ӱ��փ}�`Ih���U�a�E��6���%��>����8R澀�ξgp��:����k̾L��� �����#��4���C���S���e�=�z��L���|���ᕿ�5���2����s�	�P�Po0�G�����,0�����7�,sX�#{��
��Ƈ��숕�u֏����]�u�ʥa��'P�px@���0�u ��w����p�ݾ_ɾ�X����þ��ӾHO�4��-n��)���9�:SI�0�Y���l��H������c꓿="��9�҄�S�h���E���'�����N�9a�_E%��VB�p�d��<������  �  ���}F��V��=����k~�!�V��6�:��=�Z��:_̾Ҳ�}Y��LW���揾�`��;���=���Ӿ�����J�!��<��"_��<���䚿�ů�h���_x��A����d��n#���a��:�O%#���W�-�hN�T�{����,���袽�����8=��ʤ�ZZ����p�F|K�Y-��R�y��o;�@4ľ�|��!L��G���%y��Wƙ����1��U�ݾ{�������-*�уG��$l�騋�>7��w[����/e��d������Ox��UR�(S0��y���!���6�8v\�s����,���M�����Nm��ꓲ�[<��.���&e��'B��H&�
��ǔ����ھNv��p
��/��������E��񰣾϶��O�ϾYH��Aa�'�6�seV��~}��
���
��n廿��¿���ū������yt�mI��,��8"�;�*�+�E���o�t/���⩿�5���tÿ������yg��l򁿻\���;�˲!����� ��{�׾�]������Y���(���⡾�����>ž0Hྏ ���}�(�)�C�f������S���7��;��wĿJ,�����L�����h��*B��V+��*'�H"6�Y�V����"����岿U�����Ŀ t������1����Fy���S��5��~�Ϋ	�o��YԾ^���_����ń���ҩ�M(��8/Ѿã�+u����S2�I�O��]t�`ʏ�G]�������Ŀ¿�ʹ��L��������Z��8�}�'��)�d�>��3d�@[���ӣ�ظ�DĿ��¿�鵿Ѝ��G㊿d�k���H���,�V������p�V̾�x��oҧ�#q������!������ �ھ6��Z��"�k�;�[�{Z��⨗�D���D����Uſ����LS������ey��AN���1��&�zw/��UJ�v-t��R�����r>���  �  ��G�￹׿��������`i���8�Nr�����ʾ�,��5���=���w�x���s���{�_Έ��3���|����Ҿ����%��%�B�N.v�в������J�ݿ���e����O뿥Ͽ-���T����H^��k?�w�9�Z�M��ay�����Ŀ��@࿍��3R���`��̿�3��X����gX��$,�4����m���ʤ��p�������w��Kv�+����u������׳���'ྼ����'�X�R� ���$��%�ȿ��濟O��? ��}�&ÿP����5�?Q�i|:� w=��Y�<e������˿V�5���������� M¿�\���i~�a�I���!�����۾?߹�`
���4��G�Э~�8����k���ޙ�� ����;����1��S"8�,g�UV��'���ܖտ(�����a���ۿ����R��K�q�k K���<�YH���l�g�/����ؿ�6�y���ܞ�D�ٿ`���Ε��n�*q>����'�����վ�������]w���f��k��G}��D����;���OM྅��W�"�U�I��}�t!������I῞&��9N��2����ҿ���=����if���G��B�aV��퀿�C��	Ŀ\��8J��č��\��ѿa���Ì���`�\4��7��Z��%�о(�!����ǒ������1��Ӎ������n����̾�T����/�O�Z�m���F���Ϳ��&~��uQ��?E��ǿ�䣿)Ƀ�iY�-�B�țE��a��N��Ы��nϿ����G���G���忒�ſ
���E���mP�&(�):
�m辇�ƾ�������P$��DG��:3��%ؕ����x���Qlؾq�������W=��_l���[A��j7ؿ�]�e���I��R޿y���Ř�Awv���O�{A�s�L�q�2'��&-��+�ڿ�A���  �  ���������ֿ騿e怿C����6��6��ߙ��փ���j�Y�Z�"�V���]�up�D:���P���%þ���j�6�O�7=��%���oE����s�0���A�e����̿�꠿��~�O*X��Q�8�i�ww��>]���O�k���C��a��m���{ǿh����{k���2�R	� �׾0�����_Z~�x�e���Y��Y��c�s�z��M����(Ҿ[$�V�,�<d�_H���&¿7W� ������;�*�	��*�` ���/��]<n��R��U�'y�����ǿ������j�����u�I<�eܸ�|_���X�h�$�������˾�Χ����|��Qi�'�a�wge�ݾt��M��ݰ��<���1�K��@��}�� ���zӿ�C �������G����ݿ'������i�e�a�S��=b�)Շ��'��8ٿ����Y�\m��X����QٿW���7����H��R���ž�5���`��F=��V�r��o��v�h���E��@�����о=T�G�$���V�m���c��ݲ�T���0���������{lп<��z���}`��xY��Vr�i��������P=
�Ң�H��C��ܟ���˿�%��Ⱦs���:��K����!��-����H�������y��/y������l��ٟ�����U�yB� 5��6l��e���HƿB~�����n���T�Y��_�&U��b��>�v�ZQZ���]�����ǧ��{˿�V��ʮ����~�X 
�	�꿿+�� ���p�^��L+�a���ؾn���e���d劾�ۀ�p�y���|��Ʌ��x������%Ǿ���`���F��y��뛨��ֿ���6��!I������\�5��cz��%Yj��X���f���`���Eۿ���[`��  �  �f,�GK%������I蹿>튿[�L����0j��Ⲿ����Du�CaY�)VJ��KF��L���^�$�}�£���Ҽ����CI"� �[�����ƴſBE��vC�+(�H+,�D"�P��Xm俛����Њ��Ai��a���}�(�����̿,B�߹��`)�Ŀ+��- ���	���ݿ1{����{� �9�Ee
��]Ӿ)��n\��%l���T��bI�ݾH�q�R�-�h�В���Ԣ��4;���R3�is�����ȝ׿h�}�j+��<*���a��~ҿ㢿�M��8b��cf��z��̶��V�޿�)
��n ��,�0�)���/��ԁ̿�����d�6�)�TY����ž�H��_�����j�sX�;]Q�O�T��Qc��C~������a�����:����I�=���$��Է�^�.�$�YM-���'�����^��J�ÿ���rx�X�c��/t�n;��(X�����@b���&���-��&�js�Ȩ��������LR��A�cs�����J���,��Y�p��ab�v�^�&�e�tGx�H���餾THʾ�� ��!)��ab����H"ɿK������x�)���-���#�7���Y�H���w��q���i�����Ң�I0ѿ:d�����+���-��I"�D�⿔���������A����T���7��+���N.��!�t��i���h���r��]��
���b����aݾ[
��y;��={����ۿ		�d! �L-�'V,�� ��6�h�ֿP����o�j�]�n�Q���鯰�������:"�;�-�`+����9���ϿU؝�o�k��.0�wB��Ҿ�+��ih��񁾅�p�$=i�=l��#z�qK���������S��m���N��֊�)����U����%�>�.��)�b��������ſ�j���|��h���x�r���	�������4q�=�'��  �  �ր�B�v���X��9/��=�6���� ��Q�@�6M���־����ip��iz��"h�BAc�6#k�h���ד�4&�����>7�k�O��㑿-�Ϳ֑�k�8��`�/{�ޞ��}q��P��%�VJ��^m�������N��;v��O�ۿ�����=� cd���|��J��b�n��K��� �IF��8��zq���-��� �B�ƾ��������$]t��f�B�e�\�q��[���6���t��9��� �'�XQh�*���Ʀ����G�Lk��~��@~���g��MB��x�J��t���'���Y������>�$!���K�пn�1n���1}���d�.>�����Iֿ�x���eY��H�(��b�����׆���v��Qn�wr�#끾�v��ݐ����׾ c��=�1Ճ�W��� ��Q+�RU�qu��C��d�y���]�+$5�i�
�6=п!���J�������ʿ��V�0�@�Y�:�w�1����x� �Y�z�0���E�������cF�`��������������������{�a'��hB�����{��jN�R�{�V�bW���ѿ�J���:�lbb�5�|�����Xs���Q���'�fm��~����坿J���Bɭ�$��!�'�?���f����[��J�p���M�h�"��s��_��~�y��6�&	��׾�밾�����O���j�����:��z��b\����ѾA����/�v�p�[ʧ�k��/��a&I��em�À�/����i��nD�{��翘���#f��܏���8���P���#�\�M�ۑp�N����~�x|f�q�?�,a���ٿ�Λ�_`���$�������Ⱦ	ԧ�`U��շ������넾�V�����4������6��PC��o��������,���V�mv����W6{���^��^6����ҿ�l������G���`̿����1�T�Z���x��  �  ��v�u	l��^O�(�]������������>�C@��ؾ�ޭ�l葾.���ɦn���i���q�Dԃ��K���7��-�徬���L�5i��Yǿ1��Z1��W��?p��/v��2g�XG�!+��*�t��#c���b���q���5ԿUM���5��Z�Ur�"�u�.Zd�w'C��c�Q��C~��?m�q},��I�ǀɾ:�������{�m��Kl�ݣx��Љ������;ľ�����&�Md��G��׿ݿU����>��5a�~t�$Xs��^�0G:�9����ڿ;��0���:��_��I��]���BC�w�d�/�u��Or�>[��N6����AϿ�����*V�m��Z ����0����F��n�}�#�t���x�CK����԰�.3ھ�����;��%��:泿?���m$�7SL���j��pw�DFo�gKT�B�-����:\ɿ�l���k���x��S�ÿI��hj)�٦P��jm���w��hm�9�P��u)�� �Ot���ʆ��.D�Y��,��3���s���a���]���%���o�����Sf��.�þ�!�ן�M�S��ܑ��tʿ��	��3�I�X���q���w�Xi�HFI��+!�K��������.����è�ӈؿev��8�l�\� -t���w�zf�~DE��}���0����Iu�F�4�	u	�P�پ�F��d(��7���{����?��jl��*���skԾ(p�C�.�}l�(e��v��n����@�/Oc���v��uu� !`��g<�t��t߿5|���l���n��e���h����(E��kf�\�w�=t�й\�4�7�t����ҿ�	����\��D$��>��C�˾D���Ė�,��:U���*���������Ļ������/A�㿃� ������^�%��M���k�<�x���p���U�;
/�j����˿�ơ�X���ɞ�	�ſ��K�*�S�Q��rn��  �  UX��+O�P6�2�������`�y��#:�d��5������]��z��N����}�2��=ގ��ˢ����(P��ÈF���������.����� =���R��X��K�x�/�'.��Sؿ��q���	y��:����������-� ��[@��sT��mW��H�,�oW	�6�ϿBV��BYb�AA*�����RӾ+x��eP���)��e���m3�������������Zξ�? ��%���Z�����ȿ)Z�bA(��E���V�}�U�v,C�m$�����/ſ	ڙ��(���ˇ�7�����ѿ�a	�M1,���H���W�V�T�Ԛ@��$!�C>���ڼ��%���N��X��D��gSɾ���4e��72���`��0�������X������L㾴@��!8� u�Х��߿���!4�N��1Y��0R���:������Ό��h���������W����*�o!���7���P�M�Y���P�P�7�UT�1�翁X����|�?�H�L��qSľ�騾�B��j����#���ŏ�񵛾�䯾�[ξU������{kM�~��V0���B������>�=�T���Y�[�L�}�1�+��kܿ�A���䍿S��� 뚿=�ÿ ���"��B��V�+�Y��J�,.�Yq��Կ/}����j�	w2��� ��w����y���J��/����L�� ����0���3����޾6^�=)-���b�<%��>Ϳ3n� X*�J�G��X�حW�@KE�׌&�ɦ��oɿ��`�������إ�Q�տ&V�?.���J���Y�E]V�AFB���"�w����/��F|���tU���#��1�\E־&Ķ��⡾Im��TW��ZV��	���s����Ǿ�
�,���]=��Iz��i��!#�~L�KW5�NcO��Z��zS�4<�:��q�S︿�픿�����Z��[߳��f꿄8���8���Q��  �  ��.���'�n��m����ÿ>9���Lj��8��,�_���� оw�����������ɐ�]������l��~ؾˏ ��R���B���w�1a����ο���}%�c�*�d�.�ɔ$��D��-��(��#$��ҳq��i��������q�ѿر��9���+��C.���"�A1�Z�
�������{X��,�W(�=z�t�ƾw���K����˒��J��iC��J���{þs��;	�2�'�r�R�����Qͮ�8��I
��� �އ-�B�,��c�����$׿,O��+���'�j�n�n�$ȋ��2���e���~�"��.��;,�������iտ�勵d��'�I���!�M3�R/�����]��3���[��n��!���i��j4ӾA���M}���7�7�g��Ҕ�#���p�Hm��I'���/�EK*��5�I1���!ȿ)g���L��[=l�|�|�ƚ���¿:���E��3*)��C0�ZH)��t�I.���]ƿ�󙿩�o��8>�0��_� ��v۾*1������>���������rl���ƾhV�R�C)#���I���~�Qգ��Uҿ?i�����z,�Hr0��j&�T+���M5���G��Nz��r�hT��lF����տO���_��.��e0��%�6N�A�v7��p&��%�`�CP4�tS�7���f�־� ��⫾碾
d��_]�����E5Ӿ�����"���/�7�Z�����ﲿ-�b`���"��/��.�܁ �x���aۿ:����ǉ�w�r�-w�Xڏ��-���B�c~�=�$��H0�J�-���j��J�ؿ�E��	����0P�Dy(���� �j�;:ٶ�&m��_R��.�������{�¾Z(޾��;��!=���l��l��P�¿f�������(�(1���+��z�����ʿq̞������p�裀�	ޚ��#ſ������v/*��  �  �R�0 �e��-�ƿ�������De��B��6'��a�+�����ؾ���~Ȱ��f��Z���ľt�߾��U�-�W�I��Pn�Y���wج���ο�A�I����2���yۿ���/���Bl�:�K���E�:�Z��`���i���=˿���]��������|ݿƿ���������Y�;V9����
���оT����ծ��,������Ç;�����`���6�C�T��|��=���Ϸ�R�ٿ����������.ϿVK��pn��a^���F�F�I���g����������׿[b����V����a/ӿU���ْ��t�p%O�t�1���m9�ص�RL̾�㹾���Ty����þ�ܾxN������(���B���d�[������Ŀj"�=����K�����s�ĿL���5��L�W���H�OU�{�P�������{忖d �˰��c�%\꿵�ɿ�L������d�j��H�p�,�����x��x��˾hѼ�c���=忾C�Ѿ��쾜������3�,�P�;u�Tk��qK�� ҿ>��k��\��t0��==߿繿a��Vpt��3T��PN��Bc�M���������Ͽ��'��7�����7��S󿿴ן��C���]a���A�e�'��"����\�ྻ�ʾ�wE����Ⱦ�ݾ���I��P%��+>��]�V����_��������ݿV�� ���������gӿ����O���r�f��N�^�Q���o�́��⵿�ۿ;������s��s��)�ֿ�����0��Uo{��U�.n8��M �4��,k��K�ؾ�ƾ�����.���`Ͼ^P羝��B���b-��(H��i��������ÍǿN���F�ɛ�f�X ��ǿǿ�����ې\�%�M���Y�^���읿=�¿ڐ�fh��  �  �n��Ŭ��!���)��qF�������!u���`�9L��5�g��V+	���ﾨ�پ�5Ӿ/=ݾ�q�������#�4;�/Q�Ĩe�pz����lҖ�����h���h������9�'㡿7G����b��0=�'�&�)�"�s:1��P��|�[=��%����b��u¿"绿yP��B���տ��i����n��Z��rE�9�.�h���8�8n�=f־�tվ��#�*��+���B�?=X�H`l�p��������Y���v��@����=��2�Ù��ـ���T�ۮ3��d#��%��:�to^�oц�����K�������ν������~����e�������4~��i��cU���?�)�(�bb������n���ؾ��ݾ)k�'
�%����6�iM�rib�:�v��K�������?��*Z�����!�ÿʁ��$�����m�u�� L��r0��8&�c�.��H��Nq�,��O�����e+Ŀ~n��zյ�t饿����t��t�z��jf���Q�*m;��j$���9U��b�� {߾���w���O�J�*�$�A��X�m�l�f���!���F���w��cݹ�5�ÿ TĿ*����������N�j� DE�92/�D,+�è9��Y�Ø�������D��*����HƿD%��u���i2���쒿�:��Iw�"�b�T�M���6�M���L����Հ������s1	��;���3�b�J��b`�,�t��Ȅ��,���*��L��������ſes¿�$��\������&�\�M�;���+�&�-��B��.f�~���[`���5���@Ŀ�ſC�����̻���M���r��,Wp��\�/+F��/�c������Y��s~��������U
%�|"<�\�R��g���{��䈿(���ޥ�~���^S¿�Aƿ���᳭�J����z�W�P�]05���*��,3��+M�f�u��K���`��?����  �  �;������Ò�����0���Ԓ����������V��Ur�0%R�&y2�m\�*��Z����
����AP9�,�Y�a�x��ψ�O�����ђ�����P�����}���������Qm�~M�	�-��.��r�J��NE���!���>��J_���}������1��WA���˒��*�����lG��G+��V�������A?h���G�])��
��0�:|���qF&��D�@�d��������%��}��1���*������h��W��v4���b�B��$���������H�8J+��#J��j�QЃ�������E���:;���撿a�������ҷ���֊���}�%Q_��	?���"�������}	�K��\2���Q�$r��ۆ�����O��Zϔ�o��Bړ�ؚ�������Α������z���[�j�;��Z ����S�<���I�u�8���X��x�y���Z����i��D�������=���猕��V��K�������w�+�W�oF8�rE�����	�C���#���?�X*`�J���7��"���[|���G��$���Yŕ���������o���y1����t�*�T��5��)�F��p������b*��LG�8�g��)��mҎ�Br��P~�����D]�������m��XK���
��}���"`p�{�O��p1�~��=�����uT.�W!L���l��#��F��*ʕ��A��B���e�������A������M����g���j�\J�g�,���_<�Ҡ�����2��Q�r��U��`e��p\���O�������=��떿gP�����C%��g>���e��ZE���(��������[��� 8�kUW��w�����.����薿�g������Ax��;<��:]���o������
���`���@��3%����Z������"��M=�z,]���|������  �  ��a�S2v�_c��������糿L$���S���O������K��/�i��+B��")��!�!E-���I�Yat��񒿣p���_�������n���Ű�����v��U郿�r���]���H��T2�TM��>�*��4ؾ.cԾ�ᾏ���˞��(��0?��T�nCi���}����-����ܩ�미�S��Vֿ�>8�����/.��N�[��f8�v%���#�/[5��W��`��1H��� ��ݾ������广
���o!���A������k��V��NA��Z*�ܹ������=�_վW/׾xb�ŷ����0�Q�G�K]��Oq� j���>��g���+鯿8���¿��������m˖�E�{�ԊP��92��$�-B*��A�~h��#��_���Wn��c�¿�����a�� ا�赗�6���;k|��h�@�S���=�q�&�������V�便�۾&�㾻����%��%��C<�Q�R�mg�g�{�'$���֖��Ц�➶�(����Ŀ���~S��0'����o�lH��'/��(�o{3��IP�9�z�9���ǭ��ľ��Xſ�����<�� ���w��F`��ky�;e�%P�p�9�F�"�����T��� ����X����#��0���G��w]���q��3��A-���������ռ��rſ7�ÿ�L������:����c��u@�2-�t
,�g=�m-_�Gi��S���.�� �¿\�ſ)�������F��[k���*��'ss�?_�	�I���2���#7�0��<'徶 �����eI�\� �o�7���N���c��x�Ć�G���)���B��x���V)ƿ�����������l"����V��L8�_�*��#0��VG� �m�Fꎿ�m��&���Yſ�aĿ����_q���R���U��~׀�Y\m���X�5�B�2�+�Λ�?V�&QA�,�쾕��3t�26)�"]@��V��  �  �"D�v)g�a��#O����ȿH鿎� �Q�����ῄ6���n��o�s��)O�z�D��%U�;2� >����Ŀov�E� �zZ����}���L������'����_���=��~#��?��Y��u�Ծnx��믾#j��E4���uɾ��^~��N�ް1��xO���u�ᨓ��n��GSԿ���������m�����տ�ï�?����4e��I�ƎG��`��F������Olѿ@q�>���m������׿.�������.z���R�|L4��u�mW���辍�˾Yŷ�9	�������U��Ӿ�2�r��"�� <��p\�|��	��g[��J�*���v������ʿ]i��{ヿ�3[���G���O�:hq��;��������޿9k���eS��k�pοˬ��9����o��K��@/����������˾�8��T2�������ʾsM�������g�-��I�Ȫl�H!��H���q˿[��������6����������[����y�@0U���J��T[�5����n��ȿ��/[�O�8B �5!���ĿJ��tv��� f���D�ժ*��������+�9!;e㿾6����ƾ�ھ�g������!�',:�C�W�"~�ߗ�����~ؿ7����a��������ٿг��Ő��Cm�1Q��O���h��M�������vտ ����x�������ۿ���Qƚ��B��2[��<���#�_��a?���@ܾ��Ǿ�����F����˾u�ok �6,�O)��B�'3c��x��z`��β��3Y㿶���3F����,�FͿ#��������Aa�8�M��eU��6w����a��;�ῐ��<a�����ѿ8g��sّ��t���P�Pw4�N����O���վ��ľy����þ�{Ӿ�쾻�����1��  �  �:��wm��e��2[ƿ c��S]�x�(�Y�.�'��I���ܽ�Gd���Ov��h�Z�~��\����ȿ7=��N���*���.�ې%��9���!��� ���8a�U2�����ik˾Xj��y���œ��´���U���D��S{����޾���]$"���J�Eu������5�׿��j��h,�j�-�1�!�Z��A࿒����=���m�l�k�1���٩�LHڿ����78-�98-����x���!ݿ$K������ƞO���%�(a�SH�-��?6��F���:T�������Q���T��D�ɾ�����)m/�ɻ\�Ʋ���U��,��<��6$�c�.���+�H�����Ͽ�᡿Egik�ɸu�X0��������h�F&���/���*�X��3���Ϳ ՟�zx��C�.������ݾ.��ު����񙙾V������ƾ�ܾ���	"��s@���r�h%��ɿ���R���*�PG0�Ww(�9��L��������_���W|��n��S���y��̿Ժ ��)�]�+�0��H'����b6��3��w��{1h�Ia9����أ��]Qھ����Kn��8p���ס�����Iַ��3Ͼ�zﾓX��*��S�?���Eͫ���ۿ	1�ʽ�bw.��0�'�#�(��M�󺲿;E��D�u�{�s��6��T୿UP޿+!
�P�!��@/�C/��!� �
�vE��r��F&��u�W�R�-��������Ѿ�������"-���$��{���a<��HPؾu������D6��|c�n��C���"�����%��0�Nb-����C�[�ҿ錄G��aq�~�{�s��0����o������'�k�0��D,���Le��pпt���P}���H�'d#��#����1�ɾ⛴����ߢ������岾VǾ�e侶���$ ��  �  �<���}���� {����08�(P�HWX�fVN�V�4�����T��ڬ�O���e����ё�O��Ǔ�K��ٛ;�0 R��&X�#L�(f1�v(�>ڿ�N����m��2�	� oھ-F���p��L���7@���h�V>���/�������Ǿ}����u�P�$ǌ�EN���R��8�"���A��T��!W��kG�f6*�e�O�οFʟ�3���兿�囿�lȿ��Pm&���D��-V�V���D��h&��l�k�ſ�y��W��h"����O�˾�F������Me���Y��'q������k���~����׾���.�"rg���sԿC���A.�0J��'X��/T�gM?�qI�� ��}ٽ�G)��`Y���ۋ�9����ݿ
���42��M�@	Y�U�R��h<�H�����n���*����F�U��F�� �ƾ�e���A���O���������Q����k����ľ ����oB�����C��8뿀G�1�9�j�Q���Y���O�MM6�si�2I��د�6��������ᔿ�-��$��j��<=���S�o�Y���M�<3������ݿ�Ĥ�}�t��9�;A���辠þ���p������Ï�΋��-���LN��+�ؾ3��n~&��Y����тÿ>��^�$���C�9W��-Y�SuI�>,� k	���ҿ�ѣ�9��뉿�럿Gs̿֌�^r(��F�96X��X���F��w(�M~�`�ɿJ����n_��*�����Hܾ9����0���i������쐾�ݘ�By���3�����ۭ���4��1n�����h׿*T���/���K���Y�?�U���@�� �B3�������*��U���ю�Ԉ����߿�@���3��eN��ZZ�],T�4�=�{�Mm����<ˇ�!7L�2���(��#�о�Z�������є��쐾���N��������H;'�������  �  ��A��~���%��߂��d*��VQ�P,m�ؖv��j��iM�.�%�B����d���ۘ�wY���䞿}Uʿ���/�t8U��Wo��_v��sh��gI�r@!��'�}宿^;z��_5�S%��"Ѿ~���t
���g~�^5n�V`k�P�u����y%��5a���0𾠣�|X�}����Iҿ?��08��l\���r��%u���b���@��h�Y�忘��^���/�����L�޿��ؗ<�?�_�+t��s���_�"�<�n�.�ٿJ��?`�B�#�h���W����֞��ǈ�w�w�Z�l���n�<#~��T���]��Uξ)]���0���r�O������@�E��/f�Rv�-�q�rnY�44�ڬ�Wҿi���D6��,����X��Zf���$"��)J��Qi�~=w�*p��V���/�$���$ſ����7�L���@��fѻ��松�A��t ��_V{�׀��Ԋ����	湾�@澦���qG�3?���徿�����+��R���n���w�AZl��N�Yb'�b����d��᛿�b����iͿ!T�~�0�k�V���p�ox�W'j�BK���"����[�����oi<��H���߾ͷ��)��@���;׆�����Z������Ƭ�"ξ4� �!'���`������}ֿ��E:��~^���t��1w���d��C�tn�����&��P�������������a��Ԝ>���a�qv��	v�w�a�b�>�����ݿ�r��Kdh���+����XҾ�2�������䋾���҆��0��. ��>յ��-ܾHN��7�|y���������!RG���g��w�&Fs��[�*�5��3�hտƻ���1��g���J���M��K�#���K��j�ɏx�uwq��dW�>1�+(���ǿ/,��� R�~9�_0����žܧ�����>���E�ډ�
���:~���:¾�g���  �  9SD�����m(¿���I�1�ۢZ���w�Jր��pu�jV�H�,�T��Ŀ,G��J:��蠣�-`ѿ����6���^��z�Q���f�r�sKR��(��5��^'���\��!7�����ξ���������w���g���d���n����������q��k�b�'�[�J���B�ٿ���-@�fEf���}�:����l�[I�W��d_�峴�ɟ���	��Hﯿu�濬���D�<�i���~���~��i���D��o�]}�(�����c���$��h��ŷ���r���W���:q��Pf��Vh�Zvw�����
���p˾t��*2��hw��6��#N�R�#��WN�|~p�
���2v|��c���;�];�blٿ"������	���t��E�����(���R�߬s�K'����z�!�_� t7��l�˿S␿\�O�X��羟���/q��_ׇ�5s{���t��'{��n��(}������q#侘����I�}P����Ŀ���*3�Q�[�k2y�Յ��i�v���W�\.�+����ǿ�L��rC������VrԿT���8��9`�i�{����[�t�~T���)�m��������)��+>����5ݾ���W����@��Y���y��O���K��;V���/˾?���O�'�Xd�O��� �ݿ����BB�TWh����F���o��bK�=� ��h��������0��������꿊����F���k���������ۺk���F�����念���&4l���,�J��82Ͼ9˫�フ������܂�y���H֊������~��G�پ��
�B�8��&~�b��������<%���O��#r�����7~�u�d��o=�p��0pܿǦ������ ���fÿzQ�@M*�#YT��u��Ё��:|� �`���8�7i��,οĂ����T����C���¾�f��L���Q;��˸�����o3��������IJ�x���  �  ��A��~���%��߂��d*��VQ�P,m�ؖv��j��iM�.�%�B����d���ۘ�wY���䞿}Uʿ���/�t8U��Wo��_v��sh��gI�r@!��'�}宿^;z��_5�S%��"Ѿ~���t
���g~�^5n�V`k�P�u����y%��5a���0𾠣�|X�}����Iҿ?��08��l\���r��%u���b���@��h�Y�忘��^���/�����L�޿��ؗ<�?�_�+t��s���_�"�<�n�.�ٿJ��?`�B�#�h���W����֞��ǈ�v�w�Z�l���n�;#~��T���]��Tξ(]���0���r�~O������@�E��/f�Rv�,�q�rnY�44�ڬ�Wҿi���D6��,����X��Zf���$"��)J��Qi�~=w�*p��V���/�%���$ſ����8�L���B��gѻ��松�A��t ��_V{�׀��Ԋ����湾�@澥���qG�2?���徿�����+��R���n���w�@Zl��N�Yb'�b����d��᛿�b����iͿ!T�~�0�l�V���p�px�W'j�BK���"����[�����pi<��H���߾ͷ��)��A���;׆�����Z������Ƭ�"ξ4� �!'���`������}ֿ��E:��~^���t��1w���d��C�tn�����&��P�������������a��Ԝ>���a�qv��	v�w�a�b�>�����ݿ�r��Kdh���+����XҾ�2�������䋾���҆��0��. ��>յ��-ܾHN��7�|y���������!RG���g��w�&Fs��[�*�5��3�hտƻ���1��g���J���M��K�#���K��j�ɏx�uwq��dW�>1�+(���ǿ/,��� R�~9�_0����žܧ�����>���E�ډ�
���:~���:¾�g���  �  �<���}���� {����08�(P�HWX�fVN�V�4�����T��ڬ�O���e����ё�O��Ǔ�K��ٛ;�0 R��&X�#L�(f1�v(�>ڿ�N����m��2�	� oھ-F���p��L���7@���h�V>���/�������Ǿ}����u�P�$ǌ�EN���R��8�"���A��T��!W��kG�f6*�e�O�οFʟ�3���兿�囿�lȿ��Pm&���D��-V�V���D��h&��l�k�ſ�y��W��h"����O�˾�F������Me���Y��%q������i���|����׾���.� rg�쮜�rԿC���A.� 0J��'X��/T�gM?�qI�� ��|ٽ�G)��`Y���ۋ�9����ݿ
���42��M�A	Y�U�R��h<�I�����n���*����F�V��H��"�ƾ�e���A���O���������P����k����ľ����oB�����C��8�G�0�9�j�Q���Y���O�LM6�si�1I��د�6��������ᔿ�-��$��j��<=���S�o�Y���M�<3������ݿ�Ĥ��t��9�=A���辣þ���p������Ï�ϋ��.���MN��,�ؾ3��n~&��Y����тÿ>��^�$���C�9W��-Y�SuI�>,� k	���ҿ�ѣ�9��뉿�럿Gs̿֌�^r(��F�96X��X���F��w(�M~�`�ɿJ����n_��*�����Hܾ9����0���i������쐾�ݘ�By���3�����ۭ���4��1n�����h׿*T���/���K���Y�?�U���@�� �B3�������*��U���ю�Ԉ����߿�@���3��eN��ZZ�],T�4�=�{�Mm����<ˇ�!7L�2���(��#�о�Z�������є��쐾���N��������H;'�������  �  �:��wm��e��2[ƿ c��S]�x�(�Y�.�'��I���ܽ�Gd���Ov��h�Z�~��\����ȿ7=��N���*���.�ې%��9���!��� ���8a�U2�����ik˾Xj��y���œ��´���U���D��S{����޾���]$"���J�Eu������5�׿��j��h,�j�-�1�!�Z��A࿒����=���m�l�k�1���٩�LHڿ����78-�98-����x���!ݿ$K������ƞO���%�(a�SH�-��?6��F���9T�������Q���T��A�ɾ�����&m/�ƻ\�Ų���U��+��;��6$�b�.���+�G����߽Ͽ�᡿Dgik�ɸu�X0��������h�F&���/���*�Y��4���Ϳ՟�}x��C�.������ݾ1��ު����񙙾V���~���ƾ�ܾ���"��s@���r�g%��ɿ���Q���*�OG0�Vw(�8��K��������_���W|��n��S���y��̿Ժ ��)�]�+�0��H'����d6��3��	w��~1h�Ka9����ۣ��`Qھ����Mn��:p���ס�����Jַ��3Ͼ�zﾓX��*��S�?���Eͫ���ۿ	1�ʽ�bw.��0�'�#�(��M�󺲿;E��D�u�{�s��6��T୿UP޿+!
�P�!��@/�C/��!� �
�vE��r��F&��u�W�R�-��������Ѿ�������"-���$��{���a<��HPؾu������D6��|c�n��C���"�����%��0�Nb-����C�[�ҿ錄G��aq�~�{�s��0����o������'�k�0��D,���Le��pпt���P}���H�'d#��#����1�ɾ⛴����ߢ������岾VǾ�e侶���$ ��  �  �"D�v)g�a��#O����ȿH鿎� �Q�����ῄ6���n��o�s��)O�z�D��%U�;2� >����Ŀov�E� �zZ����}���L������'����_���=��~#��?��Y��u�Ծnx��믾#j��E4���uɾ��^~��N�ް1��xO���u�ᨓ��n��GSԿ���������m�����տ�ï�?����4e��I�ƎG��`��F������Olѿ@q�>���m������׿.�������.z���R�|L4��u�mW���辌�˾Xŷ�7	�������U�� Ӿ}2�p��"�� <��p\�z��	��e[��H�(���u������ʿ\i��{ヿ�3[���G���O�;hq��;��������޿:k���fS��k�pο!ˬ��9����o��K��@/����������˾�8��T2�������ʾpM�������e�-��I�Īl�F!��F���q˿Y��������5����������[����y�?0U���J��T[�5����n��ȿ��0[�P�9B �7!���ĿL��vv��� f���D�ت*��������+�<!;g㿾7����ƾ�ھ h������!�',:�C�W�"~�ߗ�����~ؿ7����a��������ٿг��Ő��Cm�1Q��O���h��M�������vտ ����x�������ۿ���Qƚ��B��2[��<���#�_��a?���@ܾ��Ǿ�����F����˾u�ok �6,�O)��B�'3c��x��z`��β��3Y㿶���3F����,�FͿ#��������Aa�8�M��eU��6w����a��;�ῐ��<a�����ѿ8g��sّ��t���P�Pw4�N����O���վ��ľy����þ�{Ӿ�쾻�����1��  �  ��a�S2v�_c��������糿L$���S���O������K��/�i��+B��")��!�!E-���I�Yat��񒿣p���_�������n���Ű�����v��U郿�r���]���H��T2�TM��>�*��4ؾ.cԾ�ᾏ���˞��(��0?��T�nCi���}����-����ܩ�미�S��Vֿ�>8�����/.��N�[��f8�v%���#�/[5��W��`��1H��� ��ݾ������广
���p!���A������k��V��NA��Z*�ܹ������=�^վU/׾vb�ķ����0�N�G�H]��Oq�j���>��e���(鯿8���¿��������k˖�C�{�ӊP��92��$�-B*��A�h��#��`���Yn��e�¿�����a��#ا�굗�8���?k|��h�C�S���=�s�&�������W�便�۾%�㾹����%��%��C<�N�R�mg�c�{�%$���֖��Ц�����&����Ŀ���}S��/'����o�kH��'/��(�p{3��IP�;�z�9���ǭ��ľ��Xſ�����<��"���w��H`��oy�>e��%P�s�9�H�"�����T��� ����Y����#��0���G��w]���q��3��A-���������ռ��rſ7�ÿ�L������:����c��u@�2-�t
,�g=�m-_�Gi��S���.�� �¿\�ſ)�������F��[k���*��'ss�?_�	�I���2���#7�0��<'徶 �����eI�\� �o�7���N���c��x�Ć�G���)���B��x���V)ƿ�����������l"����V��L8�_�*��#0��VG� �m�Fꎿ�m��&���Yſ�aĿ����_q���R���U��~׀�Y\m���X�5�B�2�+�Λ�?V�&QA�,�쾕��3t�26)�"]@��V��  �  �;������Ò�����0���Ԓ����������V��Ur�0%R�&y2�m\�*��Z����
����AP9�,�Y�a�x��ψ�O�����ђ�����P�����}���������Qm�~M�	�-��.��r�J��NE���!���>��J_���}������1��WA���˒��*�����lG��G+��V�������A?h���G�])��
��0�;|���qF&��D�@�d��������%��}��1���*������h��W��v4���b�B��$���������H�7J+��#J��j�PЃ�������C���8;���撿_�������з���֊���}�#Q_��	?���"�������}	�L��\2���Q�$r��ۆ�����O��\ϔ�q��Dړ�ښ�������Α������z���[�k�;��Z ����S�;���I�t�8���X��x�x���X����i��B�������;���䌕��V��I�������w�)�W�nF8�qE�����	�C���#���?�Z*`�M���7��$���^|���G��'���[ŕ���������q���{1����t�-�T��5��)�G��q������b*��LG�8�g��)��mҎ�Br��P~�����D]�������m��XK���
��}���"`p�{�O��p1�~��=�����uT.�W!L���l��#��F��*ʕ��A��B���e�������A������M����g���j�\J�g�,���_<�Ҡ�����2��Q�r��U��`e��p\���O�������=��떿gP�����C%��g>���e��ZE���(��������[��� 8�kUW��w�����.����薿�g������Ax��;<��:]���o������
���`���@��3%����Z������"��M=�z,]���|������  �  �n��Ŭ��!���)��qF�������!u���`�9L��5�g��V+	���ﾨ�پ�5Ӿ/=ݾ�q�������#�4;�/Q�Ĩe�pz����lҖ�����h���h������9�'㡿7G����b��0=�'�&�)�"�s:1��P��|�[=��%����b��u¿"绿yP��B���տ��i����n��Z��rE�9�.�h���8�8n�=f־�tվ��#�*��+���B�?=X�H`l�p��������Y���v��@����=��2�Ù��ـ���T�ڮ3��d#��%��:�so^�nц�����I�������̽������|����e�������4~��i��cU���?�'�(�ab������n���ؾ��ݾ+k�'
�'����6�iM�uib�>�v��K�������?��-Z�����#�ÿ́��	$�����o�u�� L��r0��8&�c�.��H��Nq�
,��O�����d+Ŀ|n��xյ�q饿����t��p�z��jf��Q�'m;��j$���7U��a�� {߾���x���O�L�*�&�A��X�q�l�h���!���F���w��fݹ�7�ÿ"TĿ,����������P�j�"DE�:2/�E,+�è9��Y�Ø�������D��*����HƿD%��u���i2���쒿�:��Iw�"�b�T�M���6�M���L����Հ������s1	��;���3�b�J��b`�,�t��Ȅ��,���*��L��������ſes¿�$��\������&�\�M�;���+�&�-��B��.f�~���[`���5���@Ŀ�ſC�����̻���M���r��,Wp��\�/+F��/�c������Y��s~��������U
%�|"<�\�R��g���{��䈿(���ޥ�~���^S¿�Aƿ���᳭�J����z�W�P�]05���*��,3��+M�f�u��K���`��?����  �  �R�0 �e��-�ƿ�������De��B��6'��a�+�����ؾ���~Ȱ��f��Z���ľt�߾��U�-�W�I��Pn�Y���wج���ο�A�I����2���yۿ���/���Bl�:�K���E�:�Z��`���i���=˿���]��������|ݿƿ���������Y�;V9����
���оT����ծ��,������Ç;�����`���6�C�T��|��=���Ϸ�R�ٿ����������.ϿVK��pn��a^���F�E�I���g����������׿Zb����U����_/ӿU���ْ�߿t�m%O�r�1���k9�յ�PL̾�㹾���Ty����þ�ܾ{N������(���B���d�]������Ŀl"�?����K�����t�ĿL���5��M�W���H�NU�{�P�������{忕d �ʰ��c�#\꿳�ɿ�L������a�j��H�m�,�����x��x��˾gѼ�c���>忾E�Ѿ��쾞������3�/�P�;u�Vk��sK��ҿ@��l��\��u0��?=߿�繿b��Wpt��3T��PN��Bc�M���������Ͽ��'��7�����7��S󿿴ן��C���]a���A�e�'��"����\�ྺ�ʾ�wE����Ⱦ�ݾ���I��P%��+>��]�V����_��������ݿV�� ���������gӿ����O���r�f��N�^�Q���o�́��⵿�ۿ;������s��s��)�ֿ�����0��Uo{��U�.n8��M �4��,k��K�ؾ�ƾ�����.���`Ͼ^P羝��B���b-��(H��i��������ÍǿN���F�ɛ�f�X ��ǿǿ�����ې\�%�M���Y�^���읿=�¿ڐ�fh��  �  ��.���'�n��m����ÿ>9���Lj��8��,�_���� оw�����������ɐ�]������l��~ؾˏ ��R���B���w�1a����ο���}%�c�*�d�.�ɔ$��D��-��(��#$��ҳq��i��������q�ѿر��9���+��C.���"�A1�Z�
�������{X��,�W(�=z�t�ƾw���K����˒��J��iC��K���{þs��;	�2�'�r�R�����Qͮ�8��I
��� �އ-�B�,��c�����$׿,O��+���&�j�m�n�#ȋ��2���e���~�"��.��;,�������iտ�勵d��%�I���!�K3�P/�����]��3���[��o��#���i��l4ӾD���O}���7�:�g��Ҕ�#���p�Im��I'���/�EK*��5�J1���!ȿ)g���L��\=l�{�|�ƚ���¿9���D��2*)��C0�YH)��t�G.���]ƿ�󙿦�o��8>�.��]� ��v۾(1������=���������tl���ƾkV�R�E)#���I���~�Sգ��Uҿ@i�����z,�Hr0��j&�T+���N5���G��Oz��r�hT��mF����տO���_��.��e0��%�6N�A�v7��p&��%�`�CP4�tS�6���f�־� ��⫾碾
d��_]�����E5Ӿ�����"���/�7�Z�����ﲿ-�b`���"��/��.�܁ �x���aۿ:����ǉ�w�r�-w�Xڏ��-���B�c~�=�$��H0�J�-���j��J�ؿ�E��	����0P�Dy(���� �j�;:ٶ�&m��_R��.�������{�¾Z(޾��;��!=���l��l��P�¿f�������(�(1���+��z�����ʿq̞������p�裀�	ޚ��#ſ������v/*��  �  UX��+O�P6�2�������`�y��#:�d��5������]��z��N����}�2��=ގ��ˢ����(P��ÈF���������.����� =���R��X��K�x�/�'.��Sؿ��q���	y��:����������-� ��[@��sT��mW��H�,�oW	�6�ϿBV��BYb�AA*�����RӾ+x��eP���)��e���m3�������������Zξ�? ��%���Z�����ȿ)Z�bA(��E���V�}�U�v,C�m$�����/ſ	ڙ��(���ˇ�6�����ѿ�a	�L1,���H���W�U�T�Ӛ@��$!�B>���ڼ��%���N��X��D��eSɾ���3e��72���`��0�������X����� M㾵@��!8�"u�Х�!�߿���!4�	N��1Y��0R���:������ό��h���������W����*�n!���7���P�M�Y���P�O�7�UT�0�翀X����z�?�F�I��oSľ�騾�B��i����#���ŏ�򵛾�䯾�[ξW������|kM���W0���B������>�=�T���Y�\�L�}�1�+��kܿ�A���䍿T��� 뚿=�ÿ ���"��B��V�+�Y��J�,.�Yq��Կ/}����j�	w2��� ��w����y���J��/����L�� ����0���3����޾6^�=)-���b�<%��>Ϳ3n� X*�J�G��X�حW�@KE�׌&�ɦ��oɿ��`�������إ�Q�տ&V�?.���J���Y�E]V�AFB���"�w����/��F|���tU���#��1�\E־&Ķ��⡾Im��TW��ZV��	���s����Ǿ�
�,���]=��Iz��i��!#�~L�KW5�NcO��Z��zS�4<�:��q�S︿�픿�����Z��[߳��f꿄8���8���Q��  �  ��v�u	l��^O�(�]������������>�C@��ؾ�ޭ�l葾.���ɦn���i���q�Dԃ��K���7��-�徬���L�5i��Yǿ1��Z1��W��?p��/v��2g�XG�!+��*�t��#c���b���q���5ԿUM���5��Z�Ur�"�u�.Zd�w'C��c�Q��C~��?m�q},��I�ǀɾ:�������{�m��Kl�ݣx��Љ������;ľ�����&�Md��G��׿ݿU����>��5a�~t�$Xs��^�/G:�9����ڿ;��0���:��_��I��]���BC�w�d�/�u��Or�>[��N6����AϿ�����*V�l��X ����/����F��n�}�#�t���x�CK����԰�/3ھ�����;��%��;泿?���m$�7SL���j��pw�DFo�gKT�B�-����:\ɿ�l���k���x��S�ÿH��hj)�٦P��jm���w��hm�9�P��u)�� �Ot���ʆ��.D�X��+��3���s���a���]���%���o�����Sf��/�þ�!�؟�N�S��ܑ��tʿ��	��3�J�X���q���w�Xi�IFI��+!�K��������.����è�Ԉؿev��8�l�\� -t���w�zf�~DE��}���0����Iu�F�4�	u	�P�پ�F��d(��7���z����?��jl��*���skԾ(p�C�.�}l�(e��v��n����@�/Oc���v��uu� !`��g<�t��t߿5|���l���n��e���h����(E��kf�\�w�=t�й\�4�7�t����ҿ�	����\��D$��>��C�˾D���Ė�,��:U���*���������Ļ������/A�㿃� ������^�%��M���k�<�x���p���U�;
/�j����˿�ơ�X���ɞ�	�ſ��K�*�S�Q��rn��  �  ^ߪ�����ׁ��8g�HY,����1���h�D'��0����ľ��~��G���b܀�az��-A��RV����ξ}�ށ3��{��ʵ�����'9�ot����Ww��b�����,����Z�s�!���ϼ�[ ����ҿ��Z/@��z�Z����U��w-���چ�mvS��9���ֿz���P��w��澧���Ƽ��9Ê������=��v^��e-���h��1�h�RFH� ����Ϳ\M��L�P���{ ��{j������ެ���r���kF���c�ؿV3��ʡ����N���S����8���@���ѧ�[����M{��@�|�	��]��B���Y�;��,�gQؾ�����������8e���ƈ�}�7����ƾ ����%�?�c��P���꿻'�h�a�~*��Ga���F����Ш���n�>�4��:���ʿx���.<ƿ�����.��Gh����s3������P?���1��o�h��-�C���驿�>n�$�,�ǫ��о�}��#J��$ɏ��1��:��E$��
|���@ܾ��	`:�u���C��#w�E�:�+*v�ŕ�QX���w��O
��ɰ��\�k$�����+��lb���U׿���t^B��|��o��/���M2��?�������U��R���ڿ*:���ZX���5�����Ⱦ��[(֒��a�������V��C�ľ�L����sP��+��ҿ�`�L�N��Ǆ�����y��g���Q��������H������ܿ1���C뽿�1�c���U�����%���"��]����q��Q�|���A��4�\����S��f�B����{P�S޽��~���Ɨ�t`���z��va�������Ѿ/Z��Z*���h��ꤿ���cf(���b��ҍ��	������4��GH����o���5��g���̿趿H�ȿ	���/��di�ؑ��^����  �  0����}���P��bs]�%�e�������e���&�|���ρȾ���q�������c����V���L���n��8�Ҿ���2�#x��󰿀7����1�;j�ax��BG��S;���@��ރ��	Q����|g�@���殿<̿i}��k8��#p����Gw��aʢ�EW�����J�*f�>5пA���1N�)��,��M���ן�s���0y�����KJ��E��jn��xU�p����F��G���ǿ����GD�)|��A�����EZ�����tv��X>���&�ѿ����<��;@޿U���J�G���w�������������p��D8�@�����3���#�:�����۾�+����-f���(������'������ʾи��%�� a�����P㿊� �YX����Ya��]���}��+p��߽d��-�V���tĿ����vK������a�'���^�����2���1���-��� ����^���&��]��ե�+k��h,������Ӿ�����K��Ĝ��x���;�V/�� �����߾d��m�9�X�~�cl��� �;o3��k�[V�� (��N"��?1���ل��S������� ����F����п��	���:��Pr��������^ݣ��h��x����L�A��`Կ�%���nV�@ �:����̾ ����������	)��Uo��4n���Ⱦ��W"��N��c��)�˿��#^F�xB~��O��+���j��I/���4x��~@��F���տ7U�������z⿳g�y�L�z���c���ӣ�p������Dr�y�9��K�y�����j�A�Ϩ����r���Ď��]���G$���J���]��˵� �վ����]*�V<f��0��G��[�!��kY�V��	�������!����\�e��.�j� ���ƿ#Ɀ۝¿�!��%�(���_�#y��A����  �  �S���&����p�P#C�����|տ��$_�(�3y�6�վ����!f������e��r����f���"���`߾!�
�n�2�� o�~���0	�!����M���y���������q��;�g�,m8�8�
�+GϿ맿�ʠ�Fҹ�~���@#�IIS�_~�ɶ��f���u����b�f3���?4������f�J�;��IT���$ʾ�L��]K��}\��ݑ��Ǚ�`���,ƾ�Y�L��*D���������A ��-�ӈ]��ׂ�a��Cy������eX�T(������V��z���QX��F1ɿA��3���b����b���Ì��s~��S�T{#��xￄƫ��y�H:�#2�]y�0�¾�;��6����򕾠��������4���ؾ̺���&��[�`��R�Ͽ*}���>��<m�R=�����������v�׌I�T��q�Oz������c��t޿�5�TD��lr����1���։��Rr�}�D���86ؿ����a�d���-��	���@���1������ع��.)��TG��FȾ��쾓[��9�A�u�32�����B����O�ܠ{��x������a��,�i��s:����ӿ=��a$��?/������n%��uU��D��ˍ�d������d��75����_ÿ������R�B�"�����eھ����>w��̂��w���쩾ZϺ��F־$����p�EXL�G����0�� U�}�/�!�_�����"�������+����Z�y*�������¿�����bͿ��5�x�d�ԅ�����֝������PU��'%����"��G��+�@�f��]x���Ͼ��������@�I���(��cþ}㾚	��&,���`�5���A2ҿV���@���n�N���c������8�w�x�J�~>���;ҵ������B�����hV��mE�*}s��x���  �  s�f�E
]�c*C�;  �����ƨ���*��n\���/�������nϾ����2���譥��쫾U(���T־�(�����=�8���h�u��<ȿ��](��J���`��Uf��X��t;����v�ʛ���4�����������˿g9�~+��:M���b���e��V��<8�����⿲���x��RL�t�$������p;Ǿ@����ꧾ�Q��dٰ�pKľ��Ὰ=�� ���F�O}�y�����ۿ���#B4��:S��d���c��8P�.t/��
���ѿ�����f���6����;}߿���K�7��NV��f���b�t�M�X�,�K[��LϿ¦��@4q�a?������G޾xKþ�K��dC���d������-�Ҿ���/���i/�J\Z��勿D����������@�f�[�Z�g��`��gG�$�����¿�����̍�a瘿'ͼ��I��� ��D�Uu^�*h��k^�[�D�܀!��C���b��s㐿��a�4`5�����	���ھz]þ����b ������ɾRt�AC��J�$�?�^�o�������˿����*���K�.�b��h��Z��a=�+��g���Ѵ�{�������e��Bп�e���-�eO�ٷd�g�g��9X��\:�s$�*�=��@����T�X�,��6��7���o׾��¾���Tu������tԾ���5[���(��$O�Â�sͩ�i�߿���M[6�^VU�O�f���e��ZR��1�6B��5ֿ�ǧ�����i��n����㿹|���9�{X�R�g��}d�@fO��z.�H
�Z�ҿ�����w��E��K"������a�Ͼ ���:?������	Ǿ��ݾ����	�.�4���_����WW��u����N�T�A�']���h��ga���H�wW%�<� �#�Ŀh���� ��"5����ل��21!��'E��z_��  �  H?,��&����E��.Aοr���r��;h��DF��A*��T�/���e޾8�˾K�ƾ�ϾCn侀���w��F0�!iM�21q�����jv��5ؿ͂�k��V�(���+��!��A�i�濇�������:t��Ml�� ��)�пC�l���)��+�C�!�������v��� ���MJ���\��<��X"����]򾀺׾=dɾ$�Ⱦ�gվ;��wG	�s}���9�i}X��M��m��? ���_翗>�ǡ��#+�f�)�`������eտ(���l��Rm�Rfq�av��F���BI�r�
�f[ �V�+�i*��&�?��o޿ab��Sᓿ w���R��45� ����H�*�վ�D̾)cоt�ᾶ?���>��*�1�F���g�'��#���j˿�������%��0-���'�E��J��l�ƿ�����f��lo�������������������v&���-��|'�e�D��%�п�9������J�m�b�K���/���*��N���׾L�Ҿy�۾HD��	��#��7��GT��x��s���ﲿx�ۿ�<�Z�\j*��-�<�#��(���h���=ޓ���|�^�t��M���@��oYԿ7�y��wC+�z�-��#�������Ŀ\"���n����d��E���*� ���H����։پc�ؾ��_���:_���'�ݲA�Y�`�-������&���뿀W�@�!�AA-��,��	����u�ٿDZ��������u�r�y�a��������%�a���&"���-���+�D���7��g�ѽ��->���4~�|Y���;�N�"�\?�����O��@ؾ�ܾ}U�;�ƻ��E0���K���l������G���ο�������&��.�,�(�j8�A���Geɿ���q�T�s�*́�w7��I$Ŀ ����&z'��  �  D���`h�d�࿲Lʿ=n���t��+>��h���:�u�Q�Y���<���!��6��$���B��'� �%���'��lC�d`��{�V���P��<��G0��ߝϿDc� ����ʑ�cf˿@#��]>��Y�b���E�ޔ@��AS��?|�`o��������ۿӈ�Z��H;���ٿ� ÿf=�����bE���σ�g2m���P�B�3��]�����������c����C�0�HM��i��H������2替#���R��A"׿};뿸���1���w޿�k���֞��π��rV��DA�1D��^�H7��4����Hȿ������h|��yI�r ӿ�b������#����ٌ��L��~e���H�\�,��!�خ�1	���| �tD��V"��=��Z��\v��0��U�������� �� �ɿ�L����������N׿�F��c9���Au�Q���C���N�<�p��������ŝԿ���ߛ���+��D}�`ͿZ*��-�������s��LD{��l_���B�c�'�� �S���� ������U2.��J�)g��]��E���ʚ�s�����ӿy���[��`���x7�.)Ͽ���L<��k�wEN��I���[��i��G���6E��������9������޿�9ǿCo��*ա��i��
�cu�\�X�
<��w"�
(�������u������8��dU��r�_���ْ����F(��Z~ĿRSۿVq￉��������x�Ŀk������^���I�hBL���f��!���|����˿�1��J��������@Xֿ^���]R����85�������l�{2O��,3��]���
�l���[�J�q�'�j�B��|_���{�mΊ��K���8�������I̿m��x���ʵ���e���ٿqɹ�Ю���z�r�U��lH��+S��u��L��.��H�ֿ���  �  =߰�<���,���d_���p��l��B���≰������U��;��V�ۣ4����bp�V	#�:7;���^�SV�������è�_�����س�sj���Բ���������d���L���.��=Rx�h*P�L0�����E�0l&��@�=�e�����盿W���y!��}������}s��1��ش��4�����H���\ٍ��kq��@J�>x,��%�.A���)�JOF�C�l��w��c���c�������1̴��2���;��A��Vô��`��9��������#���j�b!D�<u(�#��[����-��L�QLt��`��8��������x��г��.���y��kǵ�:���O��Z���򿇿�e��A���'��n�q� ��4�pU���}�ړ�ť������X��!+���}���0��m������������٩�ʄ�����`���=�c&����I�$�]�:�q]��5��#����
��j���lg���������+���˶��V���C��q`���"���b��B�[���:���%�����I)�V�A��\e�᥇����0��ޕ��i��T���㵿pK��L�������ﲿ�Z蔿R��
X��8�M�%���"���.�:KI�/qn��O��K3���?��<i���O���跿����yb������X�����Ϥ��쑿�y�!ZR�B�4��7$�ER#�8�1��bN�F�t��Ӣ�VͰ��η�X츿RX���f��*q����������+5��ޡ��\���vr�SL���0���"��$�}�5�aFT�p�{�������'���h���Ӹ�v)�����׷�&������g��c��������k��NG���-�
l"�+�&�(`:�׮Z����O���m��"%����ø�w��ж��Q��nL��^2��v����1�����e�:�B�!+��m"��o)�0X?�,ea��Q��3�����  �  �Y���딿�P��w�����˿2�ῗ򿙺�����cп\������Ii�{�H�sy?��4N���s����4���׿���Z��0�ￌ`ݿa�ƿAO��'���G��҅�q�$\U���8��+���	�������B%��5��],�ڋH��ge�y>���̌������5�� ޼�܏ӿҙ迋3��w���⿈$ƿ����Q����\�CnC�,B�ȞX�y���۠��p¿@���ƫ��vc���տ���+���,
�����r��h��`K�9/�T�lt��C��a����*�B��$6��S�n�o��������#,������H�Ŀ��ۿ����0�� ��j"ۿ��������{���S�p�B�IsI�]�g�A���x��2�ο]�$������	�пfù����%R��B����~���b��E��9*�������x���������)(��C�.�`�q�|���D������J��OPο2��O����t��Q��3ӿ�y��a�Wro�M�N��E�,nT��
z��,��i~��kaڿ�O�������|�࿂#ʿ`Ǵ����� ƕ�P\����x���\�'@���%�u�����؊�Z�����f�4�Q�J�m�*���c�������r��n����׿��RW�����$���7ʿ)���љ����d�>�K��"J��`������椿t~ƿ�俥���5���"��ڿDÿ/'��=��\)��ߩ���p�"�S��a7��������������#���=�'UZ�V�v�ތ��1��g���X��rRȿO&߿'����,��jf޿�:��Wɝ��ဿ�Y��H��XO�׍m�t�� B��AfѿW�	��������迖�ҿca��ﮩ�����R������!�g���J�0/��e�HD	�"��G/��]��w,���G���d�<C���  �  <j�f��ra���п
���x.�{�&�<,��b$�R&��w����̔�۰x���j��P�������ǿ>��O9�[L'�9,�z�#�Շ������Yǿ�#�����n]b�ڛA�XY&�E�[���2۾̾ʾ۴Ǿ�[Ҿu��d	�
��E5��S�Xx���������߿�}����+*�a7+�>)�z+	�Z<޿ F��=����|p��|n�������5sؿR�L��q*�5�*����m�	�}��͹����:�|��_V���7����'��Z���*ԾCOȾ.%ʾЇپ4)������$�J�?���_�:��\b���ÿ��J}���"�Ca,���(�>���IEο䡿�ꃿj1n��3x�򶒿�]���8��[���#�p�,�^�(��d����x׿�5��o=���r�FO�1�2���D}��-뾄�־�gϾ��վ[[�B�͗��0�o@M���o�(���"���eӿ�� ���/&(�s�-���%�a���Z�a俿	ʗ�O�~���p�oi�����0�ʿ(�������(���-��%�SE����<�ʿ5���W����oi���H��-�6��؉����]�ھ�ؾ���0����v"$��=��[��o���������Y�ߕ	�����<,��E-�5!��4��K�RR��o��Y�x��v�{�����D~ܿ�X���|,�/�,�� ������ ���|雿.�����^��$@��E&�_A��%��My�@aؾ}�پ5��!������+��F�[�f�F���������ƿ�u�,�x$��.��*�>������cѿ����w��,t�C~������;����ߺ���$��@.��C*���1]�ڿױ�������w��T�A�7����v
�&����D�ƭؾ��޾L)򾀋�(����4� AQ��  �  eF_��B�����L��,,"�W�D�^�H�f��\�VA�����2��᷿�c�������¿M; �3%�E.H�`�c{f���Y�M�=������l.���-���6T��-*�����뾟l˾
5���㨾a���Ӑ��Xn��0Iܾ��}���?��s��T��_�ѿ��	�-s.���N��'c�_ee�g�T���5�h��ܿ�ߩ�W���B1������Shտ�E��1��Q�
cd��Jd���Q��S2�l���Wؿ����y�GD�9��8��l�߾�¾���3=������B��#�ɾku龆V
��'��+P�-���r���-��k���:���W��pf��<b��L���)������ɿ|}��1���dz���J��a뿒e��>���Z��^g�,�`��OI�5'���[�ƿ�����Ti��:���,> �&�ܾ�<þ ܳ�}���J��8¾E�ھ*������=7���d�e���^��
����#�	JF��m_�`h�{]��pB�+@��)���⺿�k��*Ď�I���ſ���(�&���I���a�y1h�#�[�r�?������|��������F[��Z1�uf�<���G�ھ��ľ�۸��涾����Ѿ����	��=$�T`H��{�����pֿ���0�.Q�T9e��sg��V���7��o��$��魿���c9��ཀྵ��qٿ2K���3�_�S�bmf�xWf��S��e4������ܿ#B�������L��,'���D��Ӿc.��l0��;W����þ�ؾi��Az�3�.��W��h��ϱ�Ç���.<�BoY�+h���c���M�_~+�MN��Ϳ΀��Z����q���:���E���~?�c\���h��.b��J�u�(��@�2JɿZ>��ȗn�CR?�����R�Z����̾V^�������P����ʾf��,�S���=;��  �  ��b�"����tٿx
��E��;s�~ω�vT�����+�n��m@���y�ؿ���ї��V?�����T��d:K��w��*���/��j����i�*#;�*+�	ʿ�����T�XC!�h����Ͼ���^x���$���N��Hݗ��:������)��{u��\;�:�{��=��t$���%���U����~��������VE`�k0����m�ƿ���ͼ���"������+��[�����ߍ�ȍ����.[���*�{���]����<��$�@���h:�M�þH�����lꑾ(��	㜾�ǯ���;F#�����^EO�����8}ÿ4���)6�m�e�Z������v��)�|��%Q�-8!��������n���y{��r�ӿ���p�;�7�j�Ɯ��^����y��v�x�^&L�����Xz���n���3�����w��6�������%8���9���ѩ�A�����Q
�F�/�BGh��y��6ܿqi��1G�͖t�5}�����U��7Hp�d�A�L���ۿ��������O����F���L�ۗy�# �����\��ߵk���<�"��5�Ϳu���d�[�7m(��P�#�޾cP��c	������x���F��Vط���Ѿ�h��<����C�*9���{���^��c�'���W�/������������Nb��r2����_�ʿ�����Ħ�
+ſ����-�N"]�������KΎ�U����]��-�I �D͸�m��GI��f����xmԾ����==��Pǡ�6����"��}���d8ܾn/��$�_V������ƿRk	�M�7��5g�e�������E��^~��R���"�L�����������t����ֿ��==�3Kl�3J���M��v ��<�y�'sM�am�6����i�s���8��������n˾\_��/���{���=��Ӗ����Ⱦ+p��c���3��  �  ��i�Ua���Y￈�(��`������>��.����ƛ�����FUZ���#�!��y%��������Ŀ� ��i/�N�f��8��J����[��=��8I��OT�f��*ݿ4ə��Y��2��B�¾o���m���K-�����!�����������۾���͠<�0���:(�����M;�Is��
��]������b���!��G�V���"ۿ�E���-��M�Կy��|�A��-y��C��Nϡ�š��8���8y��'A�	�N�ÿ�����C�g����HL��/�������#��]L��gL���S���#�����?i��0S�����'տs���2N�v����~��M=���%�����ٙm�3�5�y��^�ʿ�����	���P�S�"�T�z���d���<ˣ�e�����C�g�6�/�����~+����v��f3�/���׾�ĳ������j��es���!��w���Y����Ծ,\�� /�,mo�;#��+���)�z�a�oP�����#3��Dz��y���.�[�`%�'��0��ƒ����ǿ�'�o�0��hh���߃���3�����J%����U����e��IF��X�`��Z&�i� ��`Ѿ޴���>����Ϟ�������~�þ��b��cE�>���{e������=�y`u�������������g��_���J�I�M��s,߿wN���5��g�ؿ���ŎC�W4{��G��MԢ�Dˢ�@��J{�~;C��'�z�ǿ�����]K�i��e���ƾgE��̜�P��Ж��~��:0��ǩξl���x_"�X	Z�v��ؿ�<�3�O�?����R�������d����$o��}7��@���ͿŐ�����#H�� �
IV�$V���6���t��]���?P���i�O�0����α��&|���8��[��Q���ER��횾E����$��棥��຾�Bݾ�m	���2��  �  V9m�Y�������#}/�ԅj�����X���ݪ����i����c�^�*�zI����������U�ʿvo�/�6���p����B˥����F���H��H^]�+#��q�X���\���/2�]����f�����._������;���g镾_	����׾}��Ŀ=�`߅��������A�B�N%~�C���/���ө���� 2���FP�E���⿄����f�� ܿK���I�������X������|0��.qI��n��ɿ�&��<oD������ܾ}E��뗾)ֈ�Ob�������\��<��1����v��JU�G˗�� ܿ���'W�ی���`��*���gP���Z��U�w�R�=���
�]ѿ馴�B���`�� u%�^�+���Lk��]"��v=���	���
r�U�6�����ϳ�Ԣz�-�3�g����Ӿ����H���u���Ѱ���L���ܘ�K=���-Ѿ�$��S/��r�Of��X�����0�t�k������������(r��V���sJe�x,��R��jſϚ����Ϳ!���B8��~r��M��$���S���s���$���_���$�p���Ԡ�c�0<&������u;����A���.���Ց������w���¿�h达*�t<F�����ſ���E�W��V����7���ڪ�0���6��JNR�9��������n��"�zO���K�5��
��O��-��|��29���K�<���Ϳ�U����L��5�3R�}�¾u/���☾6-�����׊������ʾ�����"��"\�g,���Z߿�8���X�;a��4��If������#���y��?��O��YԿܢ��ĩ¿�����&��s_�H=�����I̫��������`Xs��8��I��r�����(29�3��V$޾���I�����x��N������7Ķ��~پ6�:S3��  �  ��i�Ua���Y￈�(��`������>��.����ƛ�����FUZ���#�!��y%��������Ŀ� ��i/�N�f��8��J����[��=��8I��OT�f��*ݿ4ə��Y��2��B�¾o���m���K-�����!�����������۾���͠<�0���:(�����M;�Is��
��]������b���!��G�V���"ۿ�E���-��M�Կy��|�A��-y��C��Nϡ�š��8���8y��'A�	�N�ÿ�����C�g����GL��/�������#��\L��fL���S���#�����>i��0S�����'տs���2N�v����~��M=���%�����ٙm�3�5�y��^�ʿ�����	���P�S�"�T�z���d���<ˣ�e�����D�g�6�/�����~+����v��f3�0���׾�ĳ������j��es���!��w���Y����Ծ+\� /�,mo�;#��*���)�y�a�nP�����#3��Dz��y���.�[�`%�'��0��ƒ����ǿ�'�o�0��hh��������3�����J%����U����f��IF��Y�`��Z&�j� ��`Ѿߴ���>����О��������þ��b��cE�>���{e������=�y`u�������������g��_���J�I�M��s,߿wN���5��g�ؿ���ŎC�W4{��G��MԢ�Dˢ�@��J{�~;C��'�z�ǿ�����]K�i��e���ƾgE��̜�P��Ж��~��:0��ǩξl���x_"�X	Z�v��ؿ�<�3�O�?����R�������d����$o��}7��@���ͿŐ�����#H�� �
IV�$V���6���t��]���?P���i�O�0����α��&|���8��[��Q���ER��횾E����$��棥��຾�Bݾ�m	���2��  �  ��b�"����tٿx
��E��;s�~ω�vT�����+�n��m@���y�ؿ���ї��V?�����T��d:K��w��*���/��j����i�*#;�*+�	ʿ�����T�XC!�h����Ͼ���^x���$���N��Hݗ��:������)��{u��\;�:�{��=��t$���%���U����~��������VE`�k0����m�ƿ���ͼ���"������+��[�����ߍ�ȍ����.[���*�{���^����<��$�@���h:�M�þH�����kꑾ(��㜾�ǯ���;D#�����]EO�����7}ÿ3���)6�l�e�Y������v��)�|��%Q�-8!��������n���z{��r�ӿ���p�;�7�j�Ɯ��^����y��v�x�_&L�����Yz���n���3�����w��7�������%8���9���ѩ�@�����Q
�E�/�@Gh��y��6ܿpi��1G�̖t�5}�����U��7Hp�d�A�L���ۿ��������O����F���L�ۗy�$ �����\��ߵk���<�#��6�Ϳv���e�[�9m(��P�%�޾dP��d	������x���F��Wط���Ѿ�h��=����C�*9���{���^��c�'���W�/������������Nb��r2����_�ʿ�����Ħ�
+ſ����-�N"]�������KΎ�U����]��-�I �D͸�m��GI��f����xmԾ����==��Pǡ�6����"��}���d8ܾn/��$�_V������ƿRk	�M�7��5g�e�������E��^~��R���"�L�����������t����ֿ��==�3Kl�3J���M��v ��<�y�'sM�am�6����i�s���8��������n˾\_��/���{���=��Ӗ����Ⱦ+p��c���3��  �  eF_��B�����L��,,"�W�D�^�H�f��\�VA�����2��᷿�c�������¿M; �3%�E.H�`�c{f���Y�M�=������l.���-���6T��-*�����뾟l˾
5���㨾a���Ӑ��Xn��0Iܾ��}���?��s��T��_�ѿ��	�-s.���N��'c�_ee�g�T���5�h��ܿ�ߩ�W���B1������Shտ�E��1��Q�
cd��Jd���Q��S2�l���Wؿ����y�GD�9��8��k�߾�¾���2=������B��!�ɾhu龄V
���'��+P�+���r���-��k���:���W��pf��<b��L���)������ɿ|}��1���dz���J��a뿓e��>���Z��^g�,�`��OI�5'���]�ƿ�����Ti��:���-> �(�ܾ�<þ!ܳ�}���J��7¾D�ھ'������=7���d�d���^��
����#�JF��m_�`h�{]��pB�+@��)���⺿�k��*Ď�I���ſ���(�&���I���a�z1h�$�[�r�?������~��������F[��Z1�vf�?���I�ھ��ľ�۸��涾����Ѿ����	��=$�T`H��{�����pֿ���0�.Q�T9e��sg��V���7��o��$��魿���c9��ཀྵ��qٿ2K���3�_�S�bmf�xWf��S��e4������ܿ#B�������L��,'���D��Ӿc.��l0��;W����þ�ؾi��Az�3�.��W��h��ϱ�Ç���.<�BoY�+h���c���M�_~+�MN��Ϳ΀��Z����q���:���E���~?�c\���h��.b��J�u�(��@�2JɿZ>��ȗn�CR?�����R�Z����̾V^�������P����ʾf��,�S���=;��  �  <j�f��ra���п
���x.�{�&�<,��b$�R&��w����̔�۰x���j��P�������ǿ>��O9�[L'�9,�z�#�Շ������Yǿ�#�����n]b�ڛA�XY&�E�[���2۾̾ʾ۴Ǿ�[Ҿu��d	�
��E5��S�Xx���������߿�}����+*�a7+�>)�z+	�Z<޿ F��=����|p��|n�������5sؿR�L��q*�5�*����m�	�}��͹����:�|��_V���7����'��Y���*ԾBOȾ,%ʾ·پ1)������$�H�?���_�:��[b���ÿ��I}���"�Ca,���(�>���IEο
䡿�ꃿj1n��3x�򶒿�]���8��[���#�q�,�_�(��d����x׿�5��q=���r�FO�3�2���F}��-뾅�־�gϾ��վZ[�B�˗��0�m@M���o�
(���"���eӿ�� ���.&(�s�-���%�a���Z�`俿	ʗ�N�~���p�oi�����1�ʿ)�������(���-��%�TE����=�ʿ7���X����oi���H��-�7��ى����_�ھ�ؾ���1����w"$��=��[��o���������Y�ߕ	�����<,��E-�5!��4��K�RR��o��Y�x��v�{�����D~ܿ�X���|,�/�,�� ������ ���|雿.�����^��$@��E&�_A��%��My�@aؾ}�پ5��!������+��F�[�f�F���������ƿ�u�,�x$��.��*�>������cѿ����w��,t�C~������;����ߺ���$��@.��C*���1]�ڿױ�������w��T�A�7����v
�&����D�ƭؾ��޾L)򾀋�(����4� AQ��  �  �Y���딿�P��w�����˿2�ῗ򿙺�����cп\������Ii�{�H�sy?��4N���s����4���׿���Z��0�ￌ`ݿa�ƿAO��'���G��҅�q�$\U���8��+���	�������B%��5��],�ڋH��ge�y>���̌������5�� ޼�܏ӿҙ迋3��w���⿈$ƿ����Q����\�CnC�,B�ȞX�y���۠��p¿@���ƫ��vc���տ���+���,
�����r��h��`K�9/�T�lt��C��_����*�@��$6��S�k�o��������!,������F�Ŀ��ۿ����0�����i"ۿ��������{���S�p�B�JsI�^�g�A���x��3�ο	]�%������	�пhù����'R��D����~���b��E��9*�������x���������)(��C�+�`�n�|���C���}���J��MPο0��N����t��P��3ӿ�y��a�Vro�M�N��E�,nT��
z��,��j~��laڿ�O�������~�࿃#ʿbǴ�򄣿ƕ�Q\����x���\�)@���%�w�����ي�Z�����g�4�Q�J�m�*���c�������r��n����׿��RW�����#���7ʿ)���љ����d�>�K��"J��`������椿t~ƿ�俥���5���"��ڿDÿ/'��=��\)��ߩ���p�"�S��a7��������������#���=�'UZ�V�v�ތ��1��g���X��rRȿO&߿'����,��jf޿�:��Wɝ��ဿ�Y��H��XO�׍m�t�� B��AfѿW�	��������迖�ҿca��ﮩ�����R������!�g���J�0/��e�HD	�"��G/��]��w,���G���d�<C���  �  =߰�<���,���d_���p��l��B���≰������U��;��V�ۣ4����bp�V	#�:7;���^�SV�������è�_�����س�sj���Բ���������d���L���.��=Rx�h*P�L0�����E�0l&��@�=�e�����盿W���y!��}������}s��1��ش��4�����H���\ٍ��kq��@J�>x,��%�.A���)�JOF�C�l��w��c���c�������1̴��2���;��A��Vô��`��9��������#���j�b!D�<u(�"��Z����-�~�L�OLt��`��7��������x��г��.���y��iǵ�9���N��Y���񿇿�e��A���'��n�q� ��4�qU���}�ړ�ť������X��#+���}���0��o������������٩�˄�� ���`���=�c&����H�$�\�:�o]��5��!����
��i���jg���������+���˶��V���C��o`���"���b��A�[���:���%�����I)�W�A��\e�⥇����0������i��T���㵿rK��N�������ﲿ�[蔿T��
X��8�N�%���"���.�:KI�/qn��O��K3���?��<i���O���跿����yb������X�����Ϥ��쑿�y�!ZR�B�4��7$�ER#�8�1��bN�F�t��Ӣ�VͰ��η�X츿RX���f��*q����������+5��ޡ��\���vr�SL���0���"��$�}�5�aFT�p�{�������'���h���Ӹ�v)�����׷�&������g��c��������k��NG���-�
l"�+�&�(`:�׮Z����O���m��"%����ø�w��ж��Q��nL��^2��v����1�����e�:�B�!+��m"��o)�0X?�,ea��Q��3�����  �  D���`h�d�࿲Lʿ=n���t��+>��h���:�u�Q�Y���<���!��6��$���B��'� �%���'��lC�d`��{�V���P��<��G0��ߝϿDc� ����ʑ�cf˿@#��]>��Y�b���E�ޔ@��AS��?|�`o��������ۿӈ�Z��H;���ٿ� ÿf=�����bE���σ�g2m���P�B�3��]�����������c����C�0�HM��i��H������2替#���R��B"׿};뿸���1���w޿�k���֞��π��rV��DA�0D��^�G7��3���Hȿ���	���g|��wI�p ӿ�b������!����ٌ��L��~e���H�[�,��!�خ�1	���| �tD��V"��=��Z��\v��0��W�������� ��!�ɿ�L����!������N׿�F��c9���Au�Q���C���N�;�p��������ÝԿ���ݛ���+��B}�^ͿX*��-�������s��ID{��l_���B�a�'�� �R���� ������W2.��J�)g��]��G���ʚ�t����ӿz���[��b���z7�/)Ͽ���M<��k�xEN��I���[��i��G���6E��������9������޿�9ǿCo��*ա��i��
�cu�\�X�
<��w"�
(�������u������8��dU��r�_���ْ����F(��Z~ĿRSۿVq￉��������x�Ŀk������^���I�hBL���f��!���|����˿�1��J��������@Xֿ^���]R����85�������l�{2O��,3��]���
�l���[�J�q�'�j�B��|_���{�mΊ��K���8�������I̿m��x���ʵ���e���ٿqɹ�Ю���z�r�U��lH��+S��u��L��.��H�ֿ���  �  H?,��&����E��.Aοr���r��;h��DF��A*��T�/���e޾8�˾K�ƾ�ϾCn侀���w��F0�!iM�21q�����jv��5ؿ͂�k��V�(���+��!��A�i�濇�������:t��Ml�� ��)�пC�l���)��+�C�!�������v��� ���MJ���\��<��X"����]򾀺׾=dɾ$�Ⱦ�gվ;��wG	�s}���9�i}X��M��m��? ���_翗>�ǡ��#+�f�)�`������eտ(���l��Rm�Qfq�av��E���BI�q�
�e[ �V�+�i*��&�>��m޿_b��Qᓿ�~w���R��45������	H�)�վ�D̾*cоu�Ᾰ?���>��*�4�F���g�'��%���j˿�������%��0-���'�E��J��m�ƿ�����f��lo�������������������v&���-��|'�e�C��$�п�9������G�m�`�K���/���*��N���׾L�Ҿy�۾JD��	��#��7��GT��x��s���ﲿz�ۿ�<�Z�]j*��-�=�#��(���h���>ޓ���|�^�t��M���@��oYԿ7�y��wC+�z�-��#�������Ŀ\"���n����d��E���*� ���H����։پc�ؾ��_���:_���'�ݲA�Y�`�-������&���뿀W�@�!�AA-��,��	����u�ٿDZ��������u�r�y�a��������%�a���&"���-���+�D���7��g�ѽ��->���4~�|Y���;�N�"�\?�����O��@ؾ�ܾ}U�;�ƻ��E0���K���l������G���ο�������&��.�,�(�j8�A���Geɿ���q�T�s�*́�w7��I$Ŀ ����&z'��  �  s�f�E
]�c*C�;  �����ƨ���*��n\���/�������nϾ����2���譥��쫾U(���T־�(�����=�8���h�u��<ȿ��](��J���`��Uf��X��t;����v�ʛ���4�����������˿g9�~+��:M���b���e��V��<8�����⿲���x��RL�t�$������p;Ǿ@����ꧾ�Q��dٰ�pKľ��Ὰ=�� ���F�O}�y�����ۿ���#B4��:S��d���c��8P�.t/��
���ѿ�����f���6����:}߿���K�7��NV��f���b�s�M�X�,�J[��LϿ����>4q�_?����
��G޾wKþ�K��dC���d������/�Ҿ���1���i/�L\Z��勿F����������@�g�[�[�g��`��gG�$�����¿�����̍�`瘿&ͼ��I��� ��D�Uu^�*h��k^�[�D�ۀ!��C���b��q㐿��a�2`5�����	���ھy]þ����b ������ɾTt�BC��J�%�?�`�o�������˿����*���K�.�b��h��Z��a=�+��g���Ѵ�{�������e��Bп�e���-�eO�ٷd�g�g��9X��\:�s$�*�=��?����T�X�,��6��7���o׾��¾���Tu������tԾ���5[���(��$O�Â�sͩ�i�߿���M[6�^VU�O�f���e��ZR��1�6B��5ֿ�ǧ�����i��n����㿹|���9�{X�R�g��}d�@fO��z.�H
�Z�ҿ�����w��E��K"������a�Ͼ ���:?������	Ǿ��ݾ����	�.�4���_����WW��u����N�T�A�']���h��ga���H�wW%�<� �#�Ŀh���� ��"5����ل��21!��'E��z_��  �  �S���&����p�P#C�����|տ��$_�(�3y�6�վ����!f������e��r����f���"���`߾!�
�n�2�� o�~���0	�!����M���y���������q��;�g�,m8�8�
�+GϿ맿�ʠ�Fҹ�~���@#�IIS�_~�ɶ��f���u����b�f3���?4������f�J�;��IT���$ʾ�L��]K��}\��ݑ��Ǚ�`���,ƾ�Y�L��*D���������A ��-�ӈ]��ׂ�a��Cy������eX�T(������V��y���QX��F1ɿA��3���b����b���Ì��s~��S�S{#��xￄƫ��y�G:�"2�\y�/�¾�;��6����򕾠��������4���ؾͺ���&��[�`��S�Ͽ*}���>��<m�S=�����������v�׌I�T��q�Oz������c��t޿�5�TD��lr����0���։��Rr�|�D���76ؿ����_�d���-��	���@���1������ع��/)��UG��FȾ��쾔[��9�C�u�42�����C����O�ܠ{��x������a��,�i��s:����ӿ=��a$��?/������n%��uU��D��ˍ�d������d��75����_ÿ������R�B�"�����eھ����>w��̂��w���쩾ZϺ��F־$����p�EXL�G����0�� U�}�/�!�_�����"�������+����Z�y*�������¿�����bͿ��5�x�d�ԅ�����֝������PU��'%����"��G��+�@�f��]x���Ͼ��������@�I���(��cþ}㾚	��&,���`�5���A2ҿV���@���n�N���c������8�w�x�J�~>���;ҵ������B�����hV��mE�*}s��x���  �  0����}���P��bs]�%�e�������e���&�|���ρȾ���q�������c����V���L���n��8�Ҿ���2�#x��󰿀7����1�;j�ax��BG��S;���@��ރ��	Q����|g�@���殿<̿i}��k8��#p����Gw��aʢ�EW�����J�*f�>5пA���1N�)��,��M���ן�s���0y�����KJ��E��jn��xU�p����F��G���ǿ����GD�)|��A�����EZ�����tv��X>���&�ѿ����<��;@޿U���J�G���w�������������p��D8�@�����3���"�:�����۾�+����-f���(������(������ʾѸ��%�� a������P㿊� �YX����Ya��]���}��+p��߽d��-�V���tĿ����vK������`�'���^�����2���1���-��� ����^���&��]��ե�+k��h,������Ӿ�����K��Ĝ��x���<�W/��!�����߾d��m�9�X�~�cl��� �<o3��k�[V�� (��O"��?1���ل��S�����������F����п��	���:��Pr��������^ݣ��h��x����L�A��`Կ�%���nV�@ �:����̾�����������	)��Uo��4n���Ⱦ��W"��N��c��)�˿��#^F�xB~��O��+���j��I/���4x��~@��F���տ7U�������z⿳g�y�L�z���c���ӣ�p������Dr�y�9��K�y�����j�A�Ϩ����r���Ď��]���G$���J���]��˵� �վ����]*�V<f��0��G��[�!��kY�V��	�������!����\�e��.�j� ���ƿ#Ɀ۝¿�!��%�(���_�#y��A����  �  ������`����]����Q����Ŀ+兿_	=� ����پ#j��3E��k$��P쌾���T��H���V����h�K�q����ֿd��	�a��y�����l���g������[��5���5D�Do�|�ܿ�1ѿt����Q)��j�e5�����������bW��N��)���:�+ �󶬿��m�k�*��X ���˾O���_ގ�M_��4b���<��*Ǿ7���$��yd��L�����?�3�Xz�"��ɴ��������*ٻ�z���q�͉/� �
�ҿ�oؿ
��A=�[��l����V��I�������L��#���M&j�=�%��=����rRU�$������¾�r���>���u�������������2^۾����9�g�����]��T�J��ĉ�_���]��.��:���1�����S~[�5X�[��:[ѿ�� ����S�����>�������w��5����1������S����=ǿ����<�B��[��8��������w6���E�������h����Ǿ��� ���R����9ڿ�y �Imc�|Y��Q��iO���Q������\���'���^F�&��v��U�տ7W���+�pHl��M���������D���j��T��C8���=�d+��ް�v�k�2�Å��+ܾl\��&�������������m��c׾���~�,���l�k���&��7�5�k|��/���ÿ���h�����E���t���1��@�׿�ܿE�
�D0?�6��|���ZG��1��������&���z���k��'�d�俟���\��k"�߾��f�Ͼ�������u���Ϡ��������N�Lw�@A?�����������8L�l��d5����L�������Zϳ�AU����\����Z�®ӿ�Y����yU�CR���~�����  �  �����J��A���R���.I�����O���냿8�<��0�2޾����ʠ�8q��=$��Aq��i��\J����R �r�J����T�п9��WX�����5��G����|���X���=�����a<�K^��տG�ʿ\���"��r`�����:*������������ԝ�1dw�P�3�"��� Ȩ��[k��*���dо�ï�xc�����o����̚��ݬ��˾k���*%�eb�!���k-��,�jyo��0���z��u���5�����Li����g���(�Kh���q̿E�ѿ���S�5�'[w�lƝ��"������5���P��T
���i`�ū��ڿ�ҕ���S�%��8���tǾ{
������Ǯ��{`��� ��`@����߾���Y�9�Я��	:��E����B�4��S ���ս�!:��]�����������R��t��
濣;˿5��U.�	kK�ׇ�$��������������*���"���J�����¿S���(B����a�龴�þo���D����}�����k���lw̾��c��7�Q� ���Q	Կ9���Z���������f��M��b>��l�����>��
��ڿ4gϿf����%��b�Nړ�9A���4�����l�������y�'�5������﬿)�s�3�-D
����� ��V����L��,Ȣ����������۾L���S-�m�j�iݥ�WQ񿇬.��q��>��쉷��.��7G��n��}��j�K�*����j�пu'ֿ,���7�:hy�8�(��������*��{���b�@\!���ݿM0��<�Z�"`#�"\ ��CԾ�����㨾 �������q��Dnƾܱ���$?��M���ӻ����D�Ñ���ȥ��}������ZD��J>���;��X�S�����]� �Ϳe�|W�ڐL��f���������  �  D��в��RC��'�m��f2�l���F���C�w�=�<���B��Ǿ�b������f��}:��=糾k�ξv9��M��J��2��N���@o	��V?��S{������������p��ˣ���`�X'�q��*�¿�й��ٿ$��F����E�������s���1���y���Y� �M��!4��]�f�J�-�Ϋ���߾���������������,騾	���=۾�>�9�(�7�^��1���	ٿ� �p!S�VN��@���q����������.��"xL��&�s�߿�����O�z4!�d�Y�����@���_���U��	}��/#���LF�OC�bpɿ�#���{R�	S!����׾����q��������妾�w����ʾi��-����;�^0z��h��
&��_-�r1h��ߐ��y��Z�������Ö���u�|>:�Kg�0ѿ�Y��q�̿>��$4��(o����P��� ��c������Po���3��c �����D\��(-C�I������Ӿ�0����������ڰ�h����ܾ���f�!��Q�v���.]Ŀ�-��A��}�����������gb��&���Ӫb��#)�on��wHǿ�8��#޿�R�EH����4���s*��I����D��ኋ��\��5"��$濾[����n�96����&"�DϾiѺ�����j ������9̾Sv뾹`���0��g��O��w-ݿ�5��9U��[��G���Ǯ�z��?���B����N��P�����^��-�ÿ+��J#���[�-���"u��я�����0U��������G�O����̿����,Y�h�'�[������Ǿ+Ƕ���������龾��վ9���&���@��k��������d.���i�刑��"���M��<���Ec��
�v��n;�u�	��lӿᬼ�^�οL�<5��Dp�E�������  �  ��������R�m�(	B����z�ܿ*P��v{��bF��s!�T���~�ʾ6�|��l���Xо���]�S�(�r�P���Q��Kq����XL�vtv��Z��Č��]����d��[6�G�	�3�ο����{���F������!���P���z�u��Z������!0`���2�8'�Hȿ���g��)9��.���Ûܾ,žu긾T=��gþ�Dپ ������4���a�T��-^��n���-��=[�������"0��S~�u�U��&�F���g���z��^ ��\ɿQ0�y,1�!�_�_��$����}����z���Q���#��V�� 𵿱Љ���W�?�.����e��Շ׾ľ�������ڕξd��ʃ��!�+=E�n�w�O���׿D�"�=�{Sj����=b��mۈ��*s�rG�÷�)���ܳ��r��hk��v�ݿ���B��n��̇�ѩ��y����;o��iC�4���߿���H����K�='�YW�I�񾑫־�ǾG�¾�2ʾ��ܾ���4���/��W����β�����V �vN��0x�8;��N����L��xxf��b8�Q���;ӿ<ڬ��쥿}c��������#�#�R�\�|�����_n��y���FRb�h�4�B	��>̿i��tp��`A��> ���L�쾋Lվɾ�hȾ�BӾNu�+�����*�<���i�Qr��	�ſ]���/��X]�v��Pь�wA���;��E�W���(�
���u�¿!æ�@��75ͿE=�g)3�-�a�I˃��o�� X����|�*{S��%�T����P��'/��ڋ^��5��f�����來cоcȾ!T˾�ھ�����;�&���J��(}�d���ڿ�b�+?�r�k�YȆ��
������mt��RH�C����L4���Ť�4�����!��C�p��O���  �  �hQ�/�I��3��������¿]����M��̳`��@��[$�>��z���⾌�۾��徬O��n��I*�DG�si�P���	����̿ �����9�"�L��Q���D�U�*�,&
���տ�|������&���eݗ�T���{n�����v:��M�Y�P���C��*�V��3�8����&��пz���U�6�6�*��R'������޾�޾1�쾞
����e�3���Q���u����ZV��3oܿ3�	��'�m[A�#�O���N��=� ��B���ÿ�嚿�P��҉��`����Ͽ���n'���B���P��mN��<�Jw!���K�ҿ�Q��*��yo��tL��O/����P���쾏���M澅k��?-��$��G@��c`�����M��q��"i￿��K�1�ǴH�cSR��fK�c5�}*�g��+���&���ꇿ(Ƒ���������2�L�I��R���J��R5�gP��>����ſ�D��x���4f���E��	*�m	���$"B��6�%��ݜ�
�0���M�;�o�����>���/п���.v�zz;��N���R��{F���,��#�ڿ䯪�܏�` ���4��=�¿m������M�<���O���R���E�-��-�ji濷ٹ��N�����O�]��?���$�\E�����-�h@�����"���!��;���Y��+~����z�������)��xC�R���P��=?�&5"��E��!ȿ�(��[�������%�ӿz���O)��`D�=�R�� P��>� $#�7M��ֿ���Z���H�u��S�L�5�/�ג	�W���i��/�l��u��O`*��E�+�e�]M�����h�¿������83��J��S�7�L�u�6�Lh�D�����퀖��=�����(Ƴ��G�����3���J��  �  N�9��c���}$ҿ�ػ��ʪ�y������y�>�V��6�lM�UF�������qS"���=��|^�Ld������q���g���o���ؿ"����_��������	�6��ȿ�f�� с�	U`�C�Y�-�p�i��Cµ���߿�#����|�xr�<� �!��xPʿ����2��"w���쇿�n�� L���-��.�N�
��
��5�B�*��cH��j����O����I���೿j�ǿB(�9`���,�H��������	�M��Ӿ���ot�r�Z��^�Xa~�Z���:�ÿW��7��Λ����<!
�k�����ۿٔÿ}�� 顿�2���7��`\d��OC��Y'�,��w����D�6��ZV���x����ES��=���'���Eѿ��쿷��L��i�T�� ��ؿ�Ү�������l�m�\�)�i�A���-ު��ӿ����,�������_��4��u�Կ[�������Ҟ��ŏ�H�~�2z\��<�L:#�3Q�����7�N�(�<0D�
)e��Ƀ�y
���좿h汿��ÿx�ۿU)���
����������J���G̿an����N�h�	Wb�� y�}������] 俥N�~6�7��K���	������οS(���7�������Gv� ET���5��G�����.��K���2��P��?r���ə��g����Ż˿�W忑J��I�|>����m��fM迏J��X�����|���b�;Df�	=��������ǿ�p�b
��W�Ou�A���&���E߿��ƿ�h��I��Ë��u�����j��I� �-���9�����#��m<�Y�[��~�������k���G<����ӿt5��(������4��e�'�ڿAF��R����q�fya�݄n�[���>��W�տ|������  �  �dϿL[ӿ�ѿ(EϿ=^Ͽ��ѿ�^ӿ��ο����⬿(r���u���L�73�85,��7�ѣT����UL���2���ſ�п��ӿ|sѿ�=Ͽ��Ͽ&�ҿ�UӿѡͿ��������K����m�u�G��O1��#-�g�;��E[����ĝ�����Yȿ'�ѿS�ӿOѿ<Ͽ�[п�ӿFӿ��˿��
䤿���{�f���B��\/��L.���?��a��2����������vʿ7�ҿLӿ3tп��οd�п�ӿk+ҿ��ɿ <��?c�������R_�>��-���/�G�D��Vi�������������!Ϳ/�ӿ�ӿ��п��Ͽ3�ѿ�HԿnRҿ�Qȿ����5:�������7[�?�<�R@/�]�4�YL�[s��4��t竿9���-�Ͽ�"տ $Կr|ѿbѿAWӿ�Kտ�.ҿ��ƿɲ�ʙ�����Z�V���:���0� 9��TS� |�xb���ǰ�B�ſ/%ҿ�ֿԿҿ�ҿ\�Կ)ֿ4�ѿn�Ŀ#���[N���z�f�R���9��\2���=��[����'���r����.ɿFԿ�	׿��Կ�ҿ�Vӿ
ֿ��ֿO/ѿſ¿*���A'����u���O���9���5�5(D�4�c�T`������g���̿63ֿ��׿�Zտxӿ��Կ�;׿j/׿1п��������%����n���J��r7��a6��G�mj�0@��������s�οɠֿk?׿�ԿH-ӿX�ԿuX׿�gֿ��Ϳ�{��ݡ���ي�۽g��mF�X�5��8��L��q������Q�����пN;׿�ֿ�HԿ`Uӿ�TտB�׿��տҩ˿���� v��6؆��oa��B��?5��}:���Q���x�%��������kĿ0wҿv�׿�ֿ�ԿȨӿ9�տ]�׿��Կ�Iɿ�[��$P������[�$�?��.5���=���W�Oj���~���ղ���ǿ�  �  �֜�]����漿\�ӿ�ￋ$���s9�������d Ͽ�^���ꅿ��c�I�X��qj�80�������~ؿe- �yp�\��x��4��:鿺-ο ḿ�q��֙�y�����s���Q� d2��:�� �[	�����&��#C��d�@T���H��a����;���Ŀ~�ܿ����hp
��������)�h0��͓��_�{�+C]�t�[��w�ǖ�������.��&E�4���6�����߿�Iƿ�ڲ�0^��O���R���q�g��KF��#)���8�	�i3��b���/�"�N�5�p��U������ň�������P̿;�濉��V�(�� ����2@޿텴�����:�p�)�[�
d�6���ˣ�h�˿B{��<k�/���U�o������\ؿ	��sD�� h�������P��kq`���?��.%������zr��6#�L^=�!�]��������b���^��3����KֿVN�(�~�W���N�����o�ѿfN��:爿��i�}�^���p�[���1���ۿ��\'�7I�T��"�����ѿ\[��f��a���(���{��%Y�!8:�#?"�0/���o�%/��K��m�򡇿����2I������#Tȿ��࿅���4��n��8���	�;?�BſS���{ ���Xe��c��'��Қ�X��������1Q���`��A{ ���㿒|ʿ��[�������+���Up���N�r}1��^�L��n9�<> �wr7��V��x��܌��S��������Ͽ81�!������֞�^A�bvῸ����ד�1�v���a�w�i��i��०���ο�5������#�����	�d����ڿ��ÿ걿����(��:僿6�e���D�	*��@�G����ɡ'�R�A�C�a���������  �  H���B9���&ſ����4��Kj5�nJ��dQ�A�G���/�b���g߿�㬿e���υ��Q��7���L��*��5�ANK��TQ���F�w�/������,��4Ù��̀��4[�s�;�� �k<
�����ݾ�Z�C/�i��/��L�b�o�	ԍ�����[�Կ�����"���=��N�<"P��$A���%�?��n�̿�����C�����ۜ���ƿN
���!��>�H1O���O��4@�v�%�F�#�ٿD>���q���s��O���1�~A�G��Jc�X�ݾR�߾lq�ԩ�����K9�3�X�A~��W��?}��_��1���,��7E�~cQ��BM�Su9�	=���������z��x���l���橿oxڿ����$-�X�F�xR���L��99�������S�˿�����
��~�j�;I���,�)��j�:�N����EG��G���*���F�q�g��@��F�����ǿxJ�������6���K�`�R��I�!	1�,��]�寿�n��Wሿk��������r���7�{M�S��H�-A1�^���6����C��uX���jb�<�B��(����׵����6����7�
�d����7�+U��2x�����̯���ؿ-����$�r�?�/�P�02R��1C�/�'�����п�����N�����j堿%�ʿ����#���@�=Q�ܤQ��EB�I(��
���ݿ�s��ѩ��K�{��*X��!:�d� �t$��������ﾨ} �c?�N�%�~~@��_�ґ��켚�ܻ��!���}.���F��S�-�N�n;�(���������������7����Ӭ�>Zݿ���.���G��_S�:N�6�:��:�� ��ο�T��������o��:N���1����{G��������|��������=�.��K�S�k��  �  c�~��妿��)8���D�-p� �������~���vk�C+>�Kx�`:ؿ�����b��ʕ��/�� �0�H��Zt�����֌������,g��k:�����;ҿ��=q���?����I�eo�iȾW�����4���(�Ծ!��������.��Y�����5��`���&�y�S��n|�8��0������y?]�O�.�t��jƿ#5��Su��&�����xT)�45X��$��5���ax��=��-�X�z+��~ � #����Z^��l2�R�(c��o׾�¾.������v�ƾcN߾ƿ�#���h<��(l�蘿8̿ݽ	��5���b�����T���M5��%
y��|N�&��������Q��	��[Fӿ:����9��g������M���@���Au���J�=��=�*C���焿V�Q�.�*����
���־kož(J����ľ��վG��:��D`(��N���������b�1��R�E��fq�tM������0����l���?�����@ۿ򟯿s������;鿍��RJ�� v��̉�;���zՅ���h�*)<����3�տn���Px�t�F��$�W�
����!�׾9ʾ;�ǾѾV��C����v`7� �a�7c���y������8(�V���~��ˋ��8��V����I_��0����vʿ�?��W��<0ſ�� ��Z+��<Z�N)�����m�������Z��"-���&W¿�H����f���:�T{�z��L��FTҾ\Ⱦ�fɾ�5־�Y�m	�N�!�iC�_s��L���yϿ8l��`7���d�%}��=������ĥz�P�o>!���y����O������9ֿ �%;�Hi��0������
��W�v���K�{T�(�쿇簿����i�V���/�F������[�྅�ξZ�Ⱦ8�;X޾�O���(��q,��R��  �  �ׁ�����A���5��Iq�ת������MD����������j���/��� ��=ȿCU���bѿ��	�\Z<�tx�����4�����` ��,�����c��!)���kq����r���5�L����[þe��5l���X��R���)���8վj� ��!��[T�y
���̿B���@I�}���G���jq��tA��Gc��	��K�V�9w�������I����e����O�fم�W"���~���Y���ޞ�׽����O�Q;���Կ�G���Z�n#&��t�2�ؾ!t������퟾ K���B������Ț��H��1���k��墿�(翹s#���]�|/���g����������>�=bC�I/��ؿr��	�ſwQ����*�ߤd�����@ƥ�}����n��>ܗ��x�j�<�=��@㾿օ����J����� ����Ծa����2���8��������Ӿ����
�T�E�4����|��f����6��r��X���.��f���ӧ�����xl��c1��$�KL˿zd���rԿ�6���=���y��q��N
�����J���׏�u�e�v�*�� �L�Ĭy�6�<���m|��c�Ҿn���Z`��򖯾�?��%�Ⱦ��;9	��q*���\�7O����пv��	]K�-���H����z��3I���i��P��ɝX�=~ �����¿uS��������Q�4݆��&�������`�����xǆ�{�Q�9S�~�ؿ�{���ec���.����?Y龯�ʾM���ܯ��
�����оs6�k���8�s�r��I����!%��U_�$���=��*���މ��(Q���e����D�h���
ۿ#o��U�ȿ�J��V,��f��4���t��F6����������1z�<E>���������(��}�O���!�զ���޾i�ľj����{��ѹ��ײ¾a�۾� �p�&�I��  �  ����dÿ��Z�L��B��7���c4������xm��rG��gQ��/�F������ۿ)@ɿ�����1U��������|��������Z��7�������D>�)��&���R!y�l�3� ��6<׾���ͳ��HR��AИ��&����ž�M󾕖��XV�J+��ˋ޿��"�)�c�S���R�������H����ط������s��i2����ːпv�Ϳb��� �+�C�k��P���D�����q���7��&c����k��,)����X���^��O"��#��bHɾtb�����B����퓾b���a���<Ծ����.�7q��������7�Y�{�SƟ�^���p������H����#���B]�y ��b��˿��ؿ�Q��p@��с��P���м����U��i!��z���ffU�Z����Ϳ󍿣�J�ؐ�9afž6���u��r������I����þ����z�FE�@���'ƿo���HN����9�����ކ���"��=�����O<H��
��߿�N̿���f����V��э��|������{��,6���ݣ��d��C�?�P��d+������:�����&�&6þ�G���ԣ�>���@���͹�)y־@��&���^��n��n��k�$�v	f��ɕ�<����������	߸� ���r�u��p4�t��=�ԿO�ѿb����.���m�{T��~I������F���:?���l��I�m�lD+��H�1���ff�U�*������پۼ���?��׉������H��AK����4��"�5�q�w��f��� �:/9��U}������2���B���}��E������e�^�x�!��]�|ο�ۿ@����A������������t�������^ȭ��<���V�2��N�пЕ��\�O���������`Ͼ��������':��x��M���̾�I�݊��CI��  �  훈���ȿ����U��e���0���������S�������%���O����3�cϿ~�' ��F^��8���Q��ƙ��>���j���9Z��AI���7F�����8��Q|�	~3�����Ҿ#O��=8��r����ԍ�bo���������Hf�����W��1��"��A)�w�m�%l��⚺�J�������d���Z֢��~���9�����׿_EԿ�>�l�2��v����+M�����6���Vb��o>����u�)�/��ￌ���#�_��!��e��.�ľ�Ǧ�ѹ��Ir������J��������Ͼi&�Ґ.�7�s�q%���@��?��e��N��������`��\e������Ɓ���f�}�&������ѿ��߿���spH��v��t���,.��S��f���������^��H���ӿVX����K��^��8�|���Φ��� �������Ù�����f뾾��C$���E�>\��,�˿J>��W�{���߱����Ty��2���i[������P�j��D�RqҿM���!�7�_�� �����rl���m�����06���%����G�{h
�����R���ר:�V<����E����ǩ����u���dۤ�8/����Ѿ�) �:%�``�4u��}��#+���o��x��å��{���?������}ۣ�-����;����&ۿ3Oؿ�C���4��	x�W	���Q���������|j���G��xx��2����u륿!Hh�� *�4�*;վ���.إ�N��:@���Ө�Z����Q޾aD
�\�5��z�J������t�@��:��'̧�~���2���2������(E��v7h��M(�̆����Կ����U�I�42���7������r���s������������_���+sֿ���h�P����Qf����ʾ�g��ƣ��z��Ţ�i����pǾ@�4�W�I��  �  ����dÿ��Z�L��B��7���c4������xm��rG��gQ��/�F������ۿ)@ɿ�����1U��������|��������Z��7�������D>�)��&���R!y�l�3� ��6<׾���ͳ��HR��AИ��&����ž�M󾕖��XV�J+��ˋ޿��"�)�c�S���R�������H����ط������s��i2����ːпv�Ϳb��� �+�C�k��P���D�����q���7��&c����k��,)����X���^��O"��#��bHɾtb�����B����퓾a���a���<Ծ����.�6q��������7�Y�{�RƟ�^���p������G����#���B]�y ��b��˿��ؿ�Q��p@��с��P���м����U��i!��z���ffU�Z����Ϳ󍿣�J�ؐ�:afž6���u��r������I���þ����z�FE�@���'ƿo���HN����9�����ކ���"��=�����O<H��
��߿�N̿���f����V��э��|������{��,6���ݣ��d��C�?�P��d+������:�����&�&6þ�G���ԣ�>���@���͹�)y־@��&���^��n��n��k�$�v	f��ɕ�<����������	߸� ���r�u��p4�t��=�ԿO�ѿb����.���m�{T��~I������F���:?���l��I�m�lD+��H�1���ff�U�*������پۼ���?��׉������H��AK����4��"�5�q�w��f��� �:/9��U}������2���B���}��E������e�^�x�!��]�|ο�ۿ@����A������������t�������^ȭ��<���V�2��N�пЕ��\�O���������`Ͼ��������':��x��M���̾�I�݊��CI��  �  �ׁ�����A���5��Iq�ת������MD����������j���/��� ��=ȿCU���bѿ��	�\Z<�tx�����4�����` ��,�����c��!)���kq����r���5�L����[þe��5l���X��R���)���8վj� ��!��[T�y
���̿B���@I�}���G���jq��tA��Gc��	��K�V�9w�������I����e����O�fم�W"���~���Y���ޞ�׽����O�Q;���Կ�G���Z�n#&��t�1�ؾ!t������퟾K���B������ǚ��H��1���k��墿�(翹s#���]�{/���g����������>�=bC�I/��ؿr��	�ſwQ����*�ߤd�����Aƥ�}����n��>ܗ��x�j�<�=��A㾿ׅ����J����� ����Ծb����2���8��������Ӿ����
�S�E�4����|��e����6��r��X���.��e���ӧ�����xl��c1��$�KL˿zd���rԿ�6���=���y��q��N
�����J���׏�v�e�v�*�� �M�Ŭy�8�<���o|��d�Ҿo���[`��󖯾�?��%�Ⱦ��;9	��q*���\�7O����пv��	]K�-���H����z��3I���i��P��ɝX�=~ �����¿uS��������Q�4݆��&�������`�����xǆ�{�Q�9S�~�ؿ�{���ec���.����?Y龯�ʾM���ܯ��
�����оs6�k���8�s�r��I����!%��U_�$���=��*���މ��(Q���e����D�h���
ۿ#o��U�ȿ�J��V,��f��4���t��F6����������1z�<E>���������(��}�O���!�զ���޾i�ľj����{��ѹ��ײ¾a�۾� �p�&�I��  �  c�~��妿��)8���D�-p� �������~���vk�C+>�Kx�`:ؿ�����b��ʕ��/�� �0�H��Zt�����֌������,g��k:�����;ҿ��=q���?����I�eo�iȾW�����4���(�Ծ!��������.��Y�����5��`���&�y�S��n|�8��0������y?]�O�.�t��jƿ#5��Su��&�����xT)�45X��$��5���ax��=��-�X�z+��~ � #����Z^��l2�Q�'c��o׾�¾-������t�ƾaN߾Ŀ�"���h<��(l�蘿7̿ܽ	��5���b�����T���M5��%
y��|N�&��������Q��	��[Fӿ:����9��g������M���@���Au���J�>��=�+C���焿X�Q�0�*�������־kož(J����ľ��վF��9��B`(��N���������b�1��Q�E��fq�tM������0����l���?�����@ۿ򟯿s������;鿍��RJ�� v��̉�;���{Յ���h�+)<����5�տn���Px�u�F��$�X�
����#�׾:ʾ<�ǾѾV��D����w`7� �a�7c���y������8(�V���~��ˋ��8��V����I_��0����vʿ�?��W��<0ſ�� ��Z+��<Z�N)�����m�������Z��"-���&W¿�H����f���:�T{�z��L��FTҾ\Ⱦ�fɾ�5־�Y�m	�N�!�iC�_s��L���yϿ8l��`7���d�%}��=������ĥz�P�o>!���y����O������9ֿ �%;�Hi��0������
��W�v���K�{T�(�쿇簿����i�V���/�F������[�྅�ξZ�Ⱦ8�;X޾�O���(��q,��R��  �  H���B9���&ſ����4��Kj5�nJ��dQ�A�G���/�b���g߿�㬿e���υ��Q��7���L��*��5�ANK��TQ���F�w�/������,��4Ù��̀��4[�s�;�� �k<
�����ݾ�Z�C/�i��/��L�b�o�	ԍ�����[�Կ�����"���=��N�<"P��$A���%�?��n�̿�����C�����ۜ���ƿN
���!��>�H1O���O��4@�v�%�F�#�ٿD>���q���s��O���1�~A�G��Ic�W�ݾP�߾jq�ө�����K9�1�X�A~��W��>}��^��0���,��7E�~cQ��BM�Ru9�=���������z��x���l���橿oxڿ����$-�Y�F�yR���L��99�������T�˿�����
����j�<I���,�*��j�:�N����DG��G���*���F�o�g��@��E�����ǿwJ�������6���K�`�R��I�!	1�+��]�
寿�n��Wሿk��������s���7�|M�S��H�.A1�_���6����C��wX���jb�=�B��(����ص����7����7�
�d����7�+U��2x�����̯���ؿ-����$�r�?�/�P�02R��1C�/�'�����п�����N�����j堿%�ʿ����#���@�=Q�ܤQ��EB�I(��
���ݿ�s��ѩ��K�{��*X��!:�d� �t$��������ﾨ} �c?�N�%�~~@��_�ґ��켚�ܻ��!���}.���F��S�-�N�n;�(���������������7����Ӭ�>Zݿ���.���G��_S�:N�6�:��:�� ��ο�T��������o��:N���1����{G��������|��������=�.��K�S�k��  �  �֜�]����漿\�ӿ�ￋ$���s9�������d Ͽ�^���ꅿ��c�I�X��qj�80�������~ؿe- �yp�\��x��4��:鿺-ο ḿ�q��֙�y�����s���Q� d2��:�� �[	�����&��#C��d�@T���H��a����;���Ŀ~�ܿ����hp
��������)�h0��͓��_�{�+C]�t�[��w�ǖ�������.��&E�4���6�����߿�Iƿ�ڲ�0^��O���R���q�g��KF��#)���7�	�h3��b���/�!�N�3�p��U������Ĉ�������P̿9�濈��V�'�� ����1@޿셴�����:�p�)�[�
d�6���ˣ�i�˿C{��=k�0���U�p������\ؿ	��tD��!h�������P��mq`���?��.%������zr��6#�K^=��]��������a���^��1����KֿUN�'�}�V���N�����n�ѿfN��:爿��i�}�^���p�[���1���ۿ��\'�8I�U��#�����ѿ][��h��a���(���{��%Y�"8:�$?"�1/���p�%/��K��m�򡇿����2I������#Tȿ��࿅���4��n��8���	�;?�BſS���{ ���Xe��c��'��Қ�X��������1Q���`��A{ ���㿒|ʿ��[�������+���Up���N�r}1��^�L��n9�<> �wr7��V��x��܌��S��������Ͽ81�!������֞�^A�bvῸ����ד�1�v���a�w�i��i��०���ο�5������#�����	�d����ڿ��ÿ걿����(��:僿6�e���D�	*��@�G����ɡ'�R�A�C�a���������  �  �dϿL[ӿ�ѿ(EϿ=^Ͽ��ѿ�^ӿ��ο����⬿(r���u���L�73�85,��7�ѣT����UL���2���ſ�п��ӿ|sѿ�=Ͽ��Ͽ&�ҿ�UӿѡͿ��������K����m�u�G��O1��#-�g�;��E[����ĝ�����Yȿ'�ѿS�ӿOѿ<Ͽ�[п�ӿFӿ��˿��
䤿���{�f���B��\/��L.���?��a��2����������vʿ7�ҿLӿ3tп��οd�п�ӿl+ҿ��ɿ <��?c�������R_�>��-���/�F�D��Vi�������������!Ϳ.�ӿ�ӿ��п��Ͽ1�ѿ�HԿlRҿ�Qȿ����4:�������7[�>�<�R@/�]�4�ZL�\s��4��u竿:���.�Ͽ�"տ!$Կs|ѿcѿCWӿ�Kտ�.ҿ��ƿɲ��ʙ�����Z�V���:���0� 9��TS��~|�wb���ǰ�A�ſ-%ҿ�ֿ��Կҿ�ҿZ�Կ(ֿ3�ѿm�Ŀ"���ZN��~�z�e�R���9��\2���=��[����(���s����.ɿFԿ�	׿��Կ	�ҿ�Vӿֿ��ֿP/ѿǿ¿+���B'����u���O���9���5�5(D�5�c�T`������g���̿63ֿ��׿�Zտxӿ��Կ�;׿j/׿1п��������%����n���J��r7��a6��G�mj�0@��������s�οɠֿk?׿�ԿH-ӿX�ԿuX׿�gֿ��Ϳ�{��ݡ���ي�۽g��mF�X�5��8��L��q������Q�����пN;׿�ֿ�HԿ`Uӿ�TտB�׿��տҩ˿���� v��6؆��oa��B��?5��}:���Q���x�%��������kĿ0wҿv�׿�ֿ�ԿȨӿ9�տ]�׿��Կ�Iɿ�[��$P������[�$�?��.5���=���W�Oj���~���ղ���ǿ�  �  N�9��c���}$ҿ�ػ��ʪ�y������y�>�V��6�lM�UF�������qS"���=��|^�Ld������q���g���o���ؿ"����_��������	�6��ȿ�f�� с�	U`�C�Y�-�p�i��Cµ���߿�#����|�xr�<� �!��xPʿ����2��"w���쇿�n�� L���-��.�N�
��
��5�B�*��cH��j����O����I���೿j�ǿB(�9`���,�H��������	�M��Ӿ���ot�q�Z��^�Wa~�Z���9�ÿV��6��͛����;!
�i�����ۿהÿ|���衿�2���7��^\d��OC�Y'�+��w����E�6� [V���x����FS��?���(���Eѿ��쿸��L��i�T�� ��ؿ�Ү�������l�m�\�)�i�@���,ު��ӿ����+�������_��2��s�ԿZ�������Ҟ��ŏ�F�~�0z\��<�L:#�3Q�����7�O�(�=0D�)e��Ƀ�z
���좿j汿��ÿy�ۿV)���
����������K���H̿an����O�h�
Wb�� y�}������] 俥N�~6�7��K���	������οS(���7�������Gv� ET���5��G�����.��K���2��P��?r���ə��g����Ż˿�W忑J��I�|>����m��fM迏J��X�����|���b�;Df�	=��������ǿ�p�b
��W�Ou�A���&���E߿��ƿ�h��I��Ë��u�����j��I� �-���9�����#��m<�Y�[��~�������k���G<����ӿt5��(������4��e�'�ڿAF��R����q�fya�݄n�[���>��W�տ|������  �  �hQ�/�I��3��������¿]����M��̳`��@��[$�>��z���⾌�۾��徬O��n��I*�DG�si�P���	����̿ �����9�"�L��Q���D�U�*�,&
���տ�|������&���eݗ�T���{n�����v:��M�Y�P���C��*�V��3�8����&��пz���U�6�6�*��R'������޾�޾1�쾞
����e�3���Q���u����ZV��3oܿ3�	��'�m[A�#�O���N��=� ��B���ÿ�嚿�P��҉��`����Ͽ���n'���B���P��mN��<�Iw!���I�ҿ�Q��*��wo��tL��O/����P���쾏���M澇k��@-��$��G@��c`�����N��r��$i����L�1�ǴH�dSR��fK�c5�}*�h��+���&���ꇿ(Ƒ���������2�K�I��R���J��R5�gP��>����ſ�D��w���4f���E��	*�l	���#"B��6�&��ޜ��0���M�=�o�����>���/п���/v�zz;��N���R��{F���,��#�ڿ䯪�܏�` ���4��=�¿m������M�<���O���R���E�-��-�ji濷ٹ��N�����O�]��?���$�\E�����-�h@�����"���!��;���Y��+~����z�������)��xC�R���P��=?�&5"��E��!ȿ�(��[�������%�ӿz���O)��`D�=�R�� P��>� $#�7M��ֿ���Z���H�u��S�L�5�/�ג	�W���i��/�l��u��O`*��E�+�e�]M�����h�¿������83��J��S�7�L�u�6�Lh�D�����퀖��=�����(Ƴ��G�����3���J��  �  ��������R�m�(	B����z�ܿ*P��v{��bF��s!�T���~�ʾ6�|��l���Xо���]�S�(�r�P���Q��Kq����XL�vtv��Z��Č��]����d��[6�G�	�3�ο����{���F������!���P���z�u��Z������!0`���2�8'�Hȿ���g��)9��.���Ûܾ,žu긾T=��gþ�Dپ ������4���a�T��-^��n���-��=[�������"0��S~�u�U��&�F���g���z��^ ��\ɿQ0�y,1�!�_�_��$����}����z���Q���#��V��𵿰Љ���W�>�.����e��Ӈ׾ľ�������ەξf��˃��!�,=E�p�w�P���׿E�#�=�|Sj����>b��nۈ��*s�rG�÷�)���ܳ��r��gk��u�ݿ���B��n��̇�ѩ��x����;o��iC�4���߿���H����K�<'�XW�H�񾐫־�ǾG�¾�2ʾ��ܾ���5���/��W����β�����V �wN��0x�8;��N����L��yxf��b8�R���;ӿ<ڬ��쥿}c��������#�#�R�\�|�����_n��y���FRb�h�4�B	��>̿i��tp��`A��> ���L�쾋Lվɾ�hȾ�BӾNu�+�����*�<���i�Qr��	�ſ]���/��X]�v��Pь�wA���;��E�W���(�
���u�¿!æ�@��75ͿE=�g)3�-�a�I˃��o�� X����|�*{S��%�T����P��'/��ڋ^��5��f�����來cоcȾ!T˾�ھ�����;�&���J��(}�d���ڿ�b�+?�r�k�YȆ��
������mt��RH�C����L4���Ť�4�����!��C�p��O���  �  D��в��RC��'�m��f2�l���F���C�w�=�<���B��Ǿ�b������f��}:��=糾k�ξv9��M��J��2��N���@o	��V?��S{������������p��ˣ���`�X'�q��*�¿�й��ٿ$��F����E�������s���1���y���Y� �M��!4��]�f�J�-�Ϋ���߾���������������,騾	���=۾�>�9�(�7�^��1���	ٿ� �p!S�VN��@���q����������.��"xL��&�r�߿�����O�z4!�d�Y�����@���_���U��}��.#���LF�OC�apɿ�#���{R�	S!����׾����q��������妾�w����ʾj��.����;�_0z��h��&��`-�r1h��ߐ��y��Z�������Ö���u�|>:�Kg�0ѿ�Y��q�̿>��$4��(o����P��� ��c������Po���3��c �����C\��'-C�H������Ӿ�0����������ڰ�i����ܾ���g�!��Q�w���.]Ŀ�-��A��}�����������gb��&���Ӫb��#)�on��wHǿ�8��#޿�R�EH����4���s*��I����D��ኋ��\��5"��$濾[����n�96����&"�DϾiѺ�����j ������9̾Sv뾹`���0��g��O��w-ݿ�5��9U��[��G���Ǯ�z��?���B����N��P�����^��-�ÿ+��J#���[�-���"u��я�����0U��������G�O����̿����,Y�h�'�[������Ǿ+Ƕ���������龾��վ9���&���@��k��������d.���i�刑��"���M��<���Ec��
�v��n;�u�	��lӿᬼ�^�οL�<5��Dp�E�������  �  �����J��A���R���.I�����O���냿8�<��0�2޾����ʠ�8q��=$��Aq��i��\J����R �r�J����T�п9��WX�����5��G����|���X���=�����a<�K^��տG�ʿ\���"��r`�����:*������������ԝ�1dw�P�3�"��� Ȩ��[k��*���dо�ï�xc�����o����̚��ݬ��˾k���*%�eb�!���k-��,�jyo��0���z��u���5�����Li����g���(�Kh���q̿E�ѿ���S�5�'[w�lƝ��"������5���P��T
���i`�ū��ڿ�ҕ���S�$��8���tǾ{
������Ǯ��|`��� ��`@����߾���Z�9�Я��	:��E����B�4��S ���ս�!:��]�����������R��t��
濣;˿5��U.�	kK�ׇ�$��������������)���"���J�����¿S���(B����`�龳�þo���C����}�����k���mw̾��d��8�Q� ���R	Կ9���Z���������f��M��b>��l�����>��
��ڿ4gϿf����%��b�Nړ�9A���4�����l�������y�'�5������﬿)�s�3�-D
����� ��V����L��,Ȣ����������۾L���S-�m�j�iݥ�WQ񿇬.��q��>��쉷��.��7G��n��}��j�K�*����j�пu'ֿ,���7�:hy�8�(��������*��{���b�@\!���ݿM0��<�Z�"`#�"\ ��CԾ�����㨾 �������q��Dnƾܱ���$?��M���ӻ����D�Ñ���ȥ��}������ZD��J>���;��X�S�����]� �Ϳe�|W�ڐL��f���������  �  ~i��5_������넟��_l�C/#�r`ٿ6��Z�K���Z�羭��+��"�����|:��d���z�ž�c�����=)\��>��.=�A2��~������H���U����������ѽ�q����\�-��9�򿵰��	���=�����Ĭ���������Y������f�������nR��������(���L7�����ؾ)���r�������,��kƞ�+���iӾ���0�0���w�󩵿����I��	���µ�����e���A��-������3Q����D�-�ω��$�urT��{�����������t��:�������J��h���@:��)���.��V�f���&����seξ�Ѱ��q��N8��Q��|C���
��V�辎v�HH��ݍ��ѿ���}d��f��]�������������������J��w��1��G�l��O�����*��rn�#ɟ��I��y���;�����Ś��t3����m���$��ܿ<Ŕ��aQ�����9�ɾ����6��;
���ߦ�䢶��Ӿp� �{&�c���������3�!��S����+���;�� �������׾��(���^�G��r]��<,�1�:@�	���ޭ�����`
���n������j˒���T���D¿uK���?��+����/[ž�����禾Q]������5¾��G�m�8����ɹ��
�yL�p���ж�a���v��	T������~)��%g��%G��]�h����Z:��V��������������\�����������%���߄��;�����\���d]m�:�-�Z�9۾�b��8����9��󾨾
����8̾������^M��{���8Կa�w�e�����1���:���n��Q���������6;x��-2�(o�.���#�f�+�@�o� [������ۀ���  �  �L��G���?c�������b��2�Rӿ[���Y[K�
��l�3%þ4	�������3��^䞾����I�ʾ6����� �^�Z��G��.翧Q+��s�g��o���s��t����6��ֵ��ӏ���S�����K�޿ 0�Xb6���|�l���f������{D��ב��d��������I��
���`���7���
��_ݾ���:���C������녣������Sؾ��$Y1�k\u�·�����w�A�[����޻��Y���T������@���?���U/=��-	�B`�i�濼��4�K�\m��*��o���m���(������ڥ���|��3��_�Eڣ��e��'�}��	bӾ`ĵ��"����������v��.ƾP���T�G�d܋��̿y�[*[�LƔ�c,��%������L=���w���m��W�l�J*�r���Ǜ޿���H.$���d�1 �������d��R���"V������]��}�c�I��:	ֿ_w����P�ɜ�m����ξRص��Ө�����H�������-ؾ�#�'�W�a��ß�_���-���u�6H��Q���X������Y.��~ڶ�v����U�v���� �5k��8�w�؞��W���X/���Y��E�����^����L���G���8Ӄ���?�~	����\ʾ�r���v���誾@���[2Ǿ��辸�[�9���}�����n	�\D����+���x����i���f�����Ϲ�����N]?��]�F��� ����N��w����� ����S��������)���e�~���4������:����k���.�$9��5�ZU¾�l�������V������$?Ѿ.|���u�'M�	z����ο����w\��m��QԺ�����Q��-���V������!n�r+�4 ���࿉���Y%�(�e�G�������j����  �  Z���a������$��eH����9#Ŀ����6L�/�7�����Ӿ�ù�La��ot������ߠ��½۾sK�Y$&���Y��q��a�ԿK��DW�ȶ���B���o���N���x���̟��(}�AU;�7���տ�@˿�Q��"���^����y�����1���`��i.���u�΄3�_���.[����y���:�3���ʾ׌������@��e����ZǾ�龉6��5��q�B���Y��:�,���m�h���=e����������"��\��k;f�=�'�,��S�̿n ҿق���4��u��b��AN��	��������P��R����$_�  ��~޿>��c��,��m	��5侚�ž���D��0(�����ڶ־����`����I�a���?P����GB�҂��W����������ۡ�����ހ��zAQ����^�心�˿��࿶���/J�#Ć�k���q��N��Uǽ�HȦ�LԆ���I������ƿi��ٶQ���"�V��o߾��ž�u���ϳ�}]���˾�辁��,��`��혿6Qؿ�?��Y�����#���R��N8��m���̠�5?�+|=�m8
��<ڿ�Ͽ�����V$�xa�E�������;$��M�������&@����w�à5��������������B����a��h�ھ@�ľ#ݹ�eA����¾}�׾W��[�B=�	>y��������!�.���o������t�������-��/6���3��fh��*��k���ѿWֿ��ſ6���w�5^��u=��<��������*��u����`��!�e��i����i�3a3�1����uҾ}_��.��R⻾#ɾ��ᾦx���!���N�9��>����(
��C�z��� ���P������LE��.������oR���M�3�Ϳ����bTK�BS������l����  �  (
���<��+��;:Z��m&������ó��	��j�U�� -�l�����w׾U>ƾ�i��ɾ]ݾ
�������5�2�`��d��G��2�̢1���e�`������̞��Y���ڀ�M�����x俘�����t<̿=@��^5��k�]���5���N��T��$�|���H����b�ܿWn��+�z�;�F���"�qb�<��s'Ѿ��þ?þ��ξ������4��B�U�s��:����Կ���/�B�a�v��V��^����	��@z���p�%;�$�
��VѿS�����L�ݿ`��G�DT|�M���9����+���_��7"l�-�7��>�f�ǿ����s�h��;����#�c��O�Ͼ�Ǿ��ʾ5�ھ�}���o�@�,���S��
��{ܯ�Q�!��OU�����+1��om���[������`���*�}@����Ŀ����H����V��xx%��<Z�L��� %��������C�����[���'�E��6{��sÊ��
[��2��{��K �<I�nSҾ�;˶վ��hY��d���;�0�g�lᓿF�ÿ���Ra3�ڷg�Eɋ�Fʛ�����J��^ց��O�������d���a���пnt��7�[6m��t��TL���c���g����~�b�J������࿽���ec��	)O�L�*���������_�,Ծ�nӾ],߾�9��i��Y'�}?J�v�{��Z��uٿd��<�D��y��f��H������I�����r�9=������տ�]���d�����L���I�sA~������m�����8��e�m�Ti9�8�	�˿���XQo�{�A�A@!�K�	�7U�ܾ�Ӿ*�־�u�wY�Z���%2�13Y�N����v�����uF#�ޠV������ڗ����� ��\���'Ma��,����\(ǿ����"ÿ>�����&��U[�]>��U����  �  ��k�[�b�-J���(�����տຬ��Y���r���N��m0�t �'������龑u�����_�Q�6�loV��{��8��@ڴ��Oῢ>��|0�o�P���f� rk��h]�J�?�'q���n���������Ѥ��p%ҿ�	��/���Q�`�g��k��,\���?�^D�8����ƿ��������wf�M�D���'��k��3���*��+�K������$��A�%8b���������¿�i�Y���;��jY�&j���h���T���3����]>ؿj"��7���g���N�����;M��<��[��k��Wh��(T���4��Q�/�翲繿�����k&\��3<��>!�������|��5���O�C���0�ŭN���q��v��%٪���ҿj����%�_�G�&�a�j�l�f�d�'�K�}(�t���-ȿ'������\����¿['��>$���H�;Lc��@m�8d�kK��*�Ab�H�ؿ�q�����x�|gT��6����_�	�˪��L<���� �p&���"���=��A]�<T�������Z��f�俔���82��jR�JCh�*=m��C_�}�A�Vr�K;�9���d䛿�T�����9�ֿ����1��S�Ѯi��=m��S^��A�d�%@��d˿(H��bǋ���n���L���/�2������\��i[���=�#8��,��*I��cj���m���V'ƿ����r���=�t�[�vGl��j���V���5�K��"�ܿ�j��8���zƙ�ֵ���4D���=�8�\�3�l��j���U��f6���a�L��7y���m����b�T�B���'�L����ŗ��p7 ���tv��-6�T�e4w�=���r���/տP��u'�=�H��	c�tn��Ff��)M�I[)�>���ʿ�r��
m�������ſ�/ �&%���I��Od��  �  �$��!��f����a�v�Ϳxo���4��r���nD��qh�yE�E�(������k���E.���L���p��������0⭿
o��q�ҿ���܇����5�"��/$�t�՞�%sݿ���n���9r�)�j��D���֞�?dȿDu��^�[!���$�����'�ZC����ݿ�ƿ{+��U���⓿�&��Q�\� ;���!�};�:{����7�`jX�*�}�đ����n8����Ŀ��ڿ�a��+�_N�`y$���!��Q�Ѐ��jOͿ����N|��C�k���o����䋫��Sؿ�D�.��(�#�<�#�o����	��(�l0ֿx?������$F�������Ew�^�R�c�3��+�K��ئ��.)�-�D���g��↿�f���D���r��4Ϳ�����H���� ���%�
�����P��1.���*�������m���|�cЕ�n���ˋ���||�D$&�cp"����_��.���Bп�%����5O��o��V$n�L�J�(�.�\����? ���4��S���w�$������_�������;ֿI`�1D	�4��D�$���%�������nb�2���@����z��rs�̖��W.��پ̿b������D#��'�����J�7A �q7�_˿�T���4��F���l>����d�U%C�*�)T������'���?�`�`�u���ٕ��8���W�� �ȿ4߿=����F��l���&��$�ku�%� ���ѿ�ꦿ]���c1t���w�S*��;���r.ܿ/!�w\�5�%���%�-��܆�v���:�ٿ�Ŀ�㳿����_ᑿo�}�_�X�r�9��K$�?��1��)�.�1<J�m�Y�������⬿���u�Ͽ�\�Z�����0M"�=2'�� �g��򿆠¿���i^���dr�����,��eʽ�ح���8~��  �  8忺�ѷ�͋���6��/�a�俽
ֿ2��M\��7��� ]�F�@�i�8��E���e�f1�����85ĿzGڿ �濦*鿠G�7v��?�~�翁!�H���ҿ����𣜿����rW�h>���9�Q�I� \m�����G���ȿ�/ݿ,��A�#���k�����[����i+�g8Ͽ����ۗ��)z��R�K9<�O
;���N���t������ѱ�؋̿X�߿�T������*�.(忺�迖��h�޿�˿$��%֒���q�3�L��S:���<���S�}��������6�п?q⿋��?��(^�[&俭��6����ݿWȿ"J��^��P
m�A�J���;���A�@	\�ꃿ!���Xڼ�M�տ�W���*B鿄��D�y6�j��>���ۿ��ĿlH�������g���H��=�0F���c����a}��^E¿��ٿ?�����3|��K�De�+��E��~P���ؿ� ���9��M#��sc���F���>���K� Wl�
s��KN��ҙǿ�ݿ#�^�쿹��k����E2뿇�����4sֿ낽�v������_���F��5B��~R�s�u�)D���[����̿��῀쿕V�i�m��5�Ӌ���M��Tӿ�0����$���Z��QD�z!C�>�V�R�|�|���7㵿=�пR��)t��쿹-鿊[�z^�����9�F�⿁NϿKF��\��/`z��U�t�B�W�D�]�[��s��}~�������Կ�����=��迡���&;�z뿈g࿔Q˿:���d���*Cs���P�6�A�o�G���a�z���Ă��)����>ؿ���k��*��+r�N�翋��Y���꿴�ݿI2ǿ�ͪ�w*��1�l��OM�{�A��
K��_h��A��ș��$SĿ��ۿ�  �  0���V��8�οȫ迺���F���!�f�$�fl��=
��^忇Ͷ��Ǒ��Uv�9|i�ɰ}�$阿Ģ��A�C��wG�S%�������x� �!t�<+ʿYз�A���˖��D����b��@�L%����<�����43��R���w�ʎ��t����������ֿ�8�s
�$C�"�#��S#�7j�-���}տ�J������q�n�+�l����������%п	- �m��{"�RX$���?@�"����iٿhÿ6���������l{��V��5�2�������3#�>=��(_�ל��c��Đ��X���&�ȿs/�w����j�����X%��� �M�������ƿ���B����l�Av�@�������̕�@��f��@@%��]#����fq�9��2,ӿT1���®��Z��4]��P�r��N�7�0��u��G��B���.��K���o�抿�*��Bɭ�3��W�ѿvj�>��#����"�8
&�������A�N���qƔ��h|�ϣo����r��f�ÿ�������� �ڿ&�IM!�9��A�����h�Ϳ�P��?��k������5j�m�G�Y-�����gN%���;�~-[�!��s���Ť������ſ�ۿ�v��v���Z�n&��d%�=x����y�ٿuZ��Ì���v�
�t�3��K��^4Կ�5��w���$��g&�I��bU�����ݿ��ǿs���M���Ք� 󁿈�^�q)>���&��=���B+�7�D���f�%?���똿�������̿��㿌����t �2
'���"��X�������ɿ���^M��`�r�� |�Ⓙ:}���b�7 
�A�Ə&���$�45��������տ!���dg��B������w�m�S���5��3"����[� ��.3�GP���s��,*���  �  ���]�����ؿB�� �*�չK��c�D�k���`�pE�̸ �H���8ѽ��Қ�����t����ȿ���2>)���L��d���k�\�_���D���"����Hο�O��<s���l���I��,,������� ��&�z��I�
�޷ ��<�Qy\�u���왿�b��RO�����E6�MNU���h�vqj�XmY�|�9�S'�"��/����픿�����]���ۿ��$�5�wV�Kci���i�/X���9�Ow�E<�E���Mޜ���� �_��	?�w%#��������Ұ���ə �^���)��7G�K�i�⃉���ʿ���*����A���]�3�k�$g�C�P�.��Q�
(пG	���Ӓ�>���'����$D�|B�[r_�{�l�r�f�#�O��n/�,M��.࿋������}��CX�$9�{
���
�����i��}���\�	�}E��7�F�U��z��p���b��pۿJ$
�K�+�M�R-e��:m�Kb���F�$."�r���G����ޝ��������̿MW���*�V^N���f��m�2{a�)�F�{�$�A��q�ѿ\Ъ�������s��%Q���3������	�+)��*���Ǟ�w�yA)�z�D�Se��̅��8������P��p���`8��eW���j�=�l�.{[���;��0���激�������ԏ��di����߿D����7�j�X��ok���k�')Z��<�ݎ�Kp��<�ÿ����䇿fh�+xG���+��!�8��h������Ae�ɝ��^1�RnN���p�b���G姿JkͿi� �s7!��sC�x_�om���h�;R�O�/���	�&8ӿ����ҕ�`؜����K���Ů���C���`�	�m���g��@Q�Ի0����m��u0���'��n)���o]�~8>�5$�-����]���d�����:�!��2;���Y��~��  �  ������������+)��(]�%J��H���I��.����̄�KV�d�!�6ￄ���`���u�ĿEE��i�,�Qb��Չ�����Sޞ�M���?��+�Q�Pp��A迫[��r���bN�+�'������{eԾ�6ž�t¾�0̾�>⾪b���͙;��(j�%6��7kʿPF
�m>:���n�LL��o���'��N���Apy�D�����ڿ�0��,���}Կ�5�E%>���s�Ӕ���x���N���[���/t���?�7�M9ѿ˱���p���?��R��d����;�þ�ľ'�Ҿ_o�[X
��Q%�&cJ�/�x�������qL�K��Kk��d������s���h��3�����ʿ笰�i���@鿑����P�ב��ܗ���Y��Լ���-����c�w�/�����Ӿ�c����a���6��
�s�������о)7ʾaо�F⾘j ��@��4���]�[����y������*���^�����٢��ں���t��A���\�W�X#��@�˿����o�ǿ<0��D.���c�ݨ��O_��o����Ж�����AS��- �k���ۮ�����NU��+/�ӡ��M��M+�Qվo�Ҿ��ܾ�g�
��#�,D�7�r������ο?g�v\<�O�p��W��U����/�����t{{�@'F��!�á޿�<��;7����ؿ�;�U,@��u�癑���_V���d��_Dv�(B����oտAꟿ�ux�I�G�ķ%���f���o)޾QӾO�Ծ�[����F��c~,��fQ����;��uz�/G���M�ץ���C��9���*����A���#j�b�4��P�Ϳ#��������6�Zn��5R��D���E�����oc���ӊ�@e�[ 1���Hy��e���j�f�y�;�:!����/���cھ{Ӿ�پ�����i�*(8���a��  �  �-���ȿum�' L��	����������~���t}���¤��D���E�F�Xܿk�ɿ��濇���S�����)�����g���0��kA��+{��Q�=�A��㸿.���W=C��u��X��SFϾB�������k��Qf��u,þ���:L	�'�-��Re�#J���^�a�"���b��E�����l���}���	�����S�q��1�~��A�пWο�#��*+��#j�e ��U���f���4s��w&���ז��	j�CY)�����>��k�l�!;2��D��o��žӱ�<����o��2;���H;���F����>��\��v���O �@M7��y���]9���/��p���TI����#�[�$���0�Z�˿e ٿ��
�Y?��Ҁ�G١����]���z���4��G���lT�UR�YHҿNs��kZ�'�������o�žަ��iE��I��~eľ �߾u��`|$��T��B�ʿ��]�M����Z��9���BQ���2��Z}�� ��OG����P߿>�̿������]U�����D�������A��z�����]Y����?�)��Sc�����mJ����G*��޾��ƾ����Ķ��������Ӿ"~���i 6���m��������%�8�d�#S��s���Wv������i�����u�s�h�3�����Կe*ҿ�.��/0-��*l����S���x����z��./��	��� l�Kr+���￺u��Q*u��:�h��8��3־0¾�������o�ž�Gܾ�Q �P��ԞE�J���۵�:��K�8�1k{����:��L���p��T��ϲ��(I]�N!��-���ο��ۿ�p�d�@�%�������$���ۍ��
����۫�z��^�U�����Կ-���N_���,������_Ͼ�)������$���(;�����(���X��  �  G���� ؿJ� ���f��ޚ��1��[���dJ�����������[���_�� �j�� �ܿ���^,��p����H���x������tW��f׷��"��%V��[���ſ�n��0A����J��������n'���"���d������P�Ѿ����(���g�"������{6�����&˧��P����������UE������E��-KH��<��'���J����@�����ȫ�-_������B����N����{ڄ�'>��A���Awp�6.�L��ޮվ(_���������c��f榾+ϼ�c� ����;��Ղ�yC��7n�`^N�4���.��P��'���e����^������G-y���3�����߿h���'��CX�TX��n��Z���{������)�����Gbp���(��㿎њ���Z��"�Q����оL����ަ�Q���i��w�����ξr�����jXT�8i��z�ڿc�!��;h�u���1���]��o����g��z?�����a���!�����7�߿S	�e�-�q��ٟ������������3��#�������S�W�B��zɿ�����]H�K�4����;Z�����B^���᱾\�þg�⾩%
�5�1��np��檿k^��̛8�i���Hب�\��O�������L��3���J���RJ�TC�53���ޓ���B�"��
ͬ�d����������W�������� @�>%� ᱿[�x���6��0��@���ž��������0����˾���]����B�0E��������P�-Î�r��P���Š��wb��'���m���z�5�cR�b����ݨ���Y�����ո�����W,����������LV���q�X�)��_�mu���_�&6'���!�ھ�q���a���H��2k��]���M׾�� �Ǘ"�UX��  �  L��^T޿a�&���p�ϡ������q��{e��C8��&������6i��^&�������h���D3��_z���:I���g��/,��������̧��Z@_�����D˿'L��"CA�b��ྍ���V颾鑗�����W���g��\�̾Z��8(�4�i��%��B4����=�)(���U���b��G�������Go�������;����P������7F������H�è���P���e����������*�������!�����E��j�ꗱ�0�r��-����z�о{h��/	���4��|���P ��fз�\�ܾ���j�;��n��ÿ�}�B
W�M<���I��'���e����f�����gҪ����`�:�/���
���!�^a������/��':�����(�������lҦ���z�q)/���!�����[��� �Z�����˾1ǰ�8��,����ɡ�7���S�ɾ�������U�Hߗ��ῳ,(�58r�:��,���!���������~��3���Z�j���'��������}���4��{��ͦ�m���9�������������\�����`����(�ο�Ԍ�pH� l�T���Ⱦ����C}��pѥ�{(��[�����ݾ�]�0�L:r��k��#����?��6���b��&n����������u������@��1�R����z��.Q�����J�6����T���j������������������fŋ���G���M͵�U{��5�A-��P�����c2��������e����ƾ�%�����B��݇�tuƿB,�r�X�������Q]������3��/�����������S<�R�	�E�q����"�C�b�r��T���K���XB��Q�������{��/!|��|0�D�@��_�`�!�%�R��r�վ����+����æ��ʪ�H{���GҾ)���-!�qY��  �  G���� ؿJ� ���f��ޚ��1��[���dJ�����������[���_�� �j�� �ܿ���^,��p����H���x������tW��f׷��"��%V��[���ſ�n��0A����J��������n'���"���d������P�Ѿ����(���g�"������{6�����&˧��P����������UE������E��-KH��<��'���J����@�����ȫ�-_������B����N����{ڄ�'>��A���Awp�6.�L��ޮվ(_���������c��f榾*ϼ�c� ����;��Ղ�xC��7n�`^N�4���.��P��'���e����^������G-y���3�����߿h���'��CX�TX��n��Z���|������)�����Gbp���(��㿏њ���Z� 	"�Q����оM����ަ�Q���i��w�����ξr�����iXT�7i��y�ڿc�!��;h�u���1���]��o����g��y?�����a���!�����7�߿S	�e�-�q��ٟ������������3��#�������T�W�B��zɿ�����]H�K�5����;Z�����C^���᱾\�þg�⾪%
�5�1��np��檿k^��̛8�i���Hب�\��O�������L��3���J���RJ�TC�53���ޓ���B�"��
ͬ�d����������W�������� @�>%� ᱿[�x���6��0��@���ž��������0����˾���]����B�0E��������P�-Î�r��P���Š��wb��'���m���z�5�cR�b����ݨ���Y�����ո�����W,����������LV���q�X�)��_�mu���_�&6'���!�ھ�q���a���H��2k��]���M׾�� �Ǘ"�UX��  �  �-���ȿum�' L��	����������~���t}���¤��D���E�F�Xܿk�ɿ��濇���S�����)�����g���0��kA��+{��Q�=�A��㸿.���W=C��u��X��SFϾB�������k��Qf��u,þ���:L	�'�-��Re�#J���^�a�"���b��E�����l���}���	�����S�q��1�~��A�пWο�#��*+��#j�e ��U���f���4s��w&���ז��	j�CY)�����>��k�l�!;2��D��o��žӱ�;����o��1;���H;���E���>��\��v���O �@M7��y���]9���/��p���TI����#�[�$���0�Z�˿e ٿ��
�Y?��Ҁ�G١����]���z���4��G���lT�UR�YHҿOs��lZ�Ó'�������p�žަ��iE��H��~eľ��߾u��_|$��T��B�ʿ��]�M����Z��9���BQ���2��Z}�� ��OG����P߿>�̿������]U�����D�������A��z�����]Y����?�)��Tc�����mJ����H*��޾��ƾ����Ķ��������Ӿ#~���i 6���m��������%�8�d�#S��s���Wv������i�����u�s�h�3�����Կe*ҿ�.��/0-��*l����S���x����z��./��	��� l�Kr+���￺u��Q*u��:�h��8��3־0¾�������o�ž�Gܾ�Q �P��ԞE�J���۵�:��K�8�1k{����:��L���p��T��ϲ��(I]�N!��-���ο��ۿ�p�d�@�%�������$���ۍ��
����۫�z��^�U�����Կ-���N_���,������_Ͼ�)������$���(;�����(���X��  �  ������������+)��(]�%J��H���I��.����̄�KV�d�!�6ￄ���`���u�ĿEE��i�,�Qb��Չ�����Sޞ�M���?��+�Q�Pp��A迫[��r���bN�+�'������{eԾ�6ž�t¾�0̾�>⾪b���͙;��(j�%6��7kʿPF
�m>:���n�LL��o���'��N���Apy�D�����ڿ�0��,���}Կ�5�E%>���s�Ӕ���x���N���[���/t���?�7�M9ѿ˱���p���?��R��d����;�þ�ľ&�Ҿ]o�ZX
��Q%�%cJ� /�w�������pL�J��Kk��c������s���h��3�����ʿ笰�i���@鿑����P�ב��ݗ���Y��Լ���-����c�x�/�����Ӿ�d����a���6��
�t�������о)7ʾaо�F⾗j ��@��4���]�Z����y������*���^�����٢��ٺ���t��A���[�W�X#��@�˿����o�ǿ<0��D.���c�ݨ��O_��o����Ж�����AS��- �l���ۮ�����NU��+/�ԡ��M��N+�Qվp�Ҿ��ܾ�h�
��#�,D�7�r������ο?g�v\<�O�p��W��U����/�����t{{�@'F��!�á޿�<��;7����ؿ�;�U,@��u�癑���_V���d��_Dv�(B����oտAꟿ�ux�I�G�ķ%���f���o)޾QӾO�Ծ�[����F��c~,��fQ����;��uz�/G���M�ץ���C��9���*����A���#j�b�4��P�Ϳ#��������6�Zn��5R��D���E�����oc���ӊ�@e�[ 1���Hy��e���j�f�y�;�:!����/���cھ{Ӿ�پ�����i�*(8���a��  �  ���]�����ؿB�� �*�չK��c�D�k���`�pE�̸ �H���8ѽ��Қ�����t����ȿ���2>)���L��d���k�\�_���D���"����Hο�O��<s���l���I��,,������� ��&�z��I�
�޷ ��<�Qy\�u���왿�b��RO�����E6�MNU���h�vqj�XmY�|�9�S'�"��/����픿�����]���ۿ��$�5�wV�Kci���i�/X���9�Ow�E<�E���Mޜ���� �_��	?�w%#��������Ѱ���ə �]���)��7G�I�i�჉���ʿ���*����A���]�2�k�$g�B�P�.��Q�
(пG	���Ӓ�>���'����%D�|B�\r_�{�l�s�f�#�O��n/�,M��.࿍�������}��CX�$9�|
���
�����i��|���[�	�|E��7�D�U��z��p���b��pۿI$
�J�+�M�R-e��:m�Kb���F�$."�r���F����ޝ��������̿MW���*�W^N���f��m�3{a�*�F�{�$�A��r�ѿ^Ъ�������s��%Q���3������	�-)��+���Ȟ�w�zA)�z�D�Se��̅��8������P��o���`8��eW���j�=�l�.{[���;��0���激�������ԏ��di����߿D����7�j�X��ok���k�')Z��<�ݎ�Kp��<�ÿ����䇿fh�+xG���+��!�8��h������Ae�ɝ��^1�RnN���p�b���G姿JkͿi� �s7!��sC�x_�om���h�;R�O�/���	�&8ӿ����ҕ�`؜����K���Ů���C���`�	�m���g��@Q�Ի0����m��u0���'��n)���o]�~8>�5$�-����]���d�����:�!��2;���Y��~��  �  0���V��8�οȫ迺���F���!�f�$�fl��=
��^忇Ͷ��Ǒ��Uv�9|i�ɰ}�$阿Ģ��A�C��wG�S%�������x� �!t�<+ʿYз�A���˖��D����b��@�L%����<�����43��R���w�ʎ��t����������ֿ�8�s
�$C�"�#��S#�7j�-���}տ�J������q�n�+�l����������%п	- �m��{"�RX$���?@�"����iٿhÿ6���������l{��V��5�1�������3#�==��(_�֜��c��Ð��V���$�ȿq/�v����j�����X%��� �M�������ƿ���B����l�Bv�@�������̕�@��f��A@%��]#����gq�:��4,ӿU1���®��Z��5]��Q�r��N�8�0��u��G��B���.��K���o�抿�*��Aɭ�2��U�ѿuj�=��"����"�8
&�������A�N���qƔ��h|�ϣo����r��f�ÿ�������� �ۿ&�JM!�9��A�����j�Ϳ�P��?��k����� 6j�n�G�Y-�����gN%���;�~-[�!��s���Ť������ſ�ۿ�v��v���Z�n&��d%�=x����y�ٿuZ��Ì���v�
�t�3��K��^4Կ�5��w���$��g&�I��bU�����ݿ��ǿs���M���Ք� 󁿈�^�q)>���&��=���B+�7�D���f�%?���똿�������̿��㿌����t �2
'���"��X�������ɿ���^M��`�r�� |�Ⓙ:}���b�7 
�A�Ə&���$�45��������տ!���dg��B������w�m�S���5��3"����[� ��.3�GP���s��,*���  �  8忺�ѷ�͋���6��/�a�俽
ֿ2��M\��7��� ]�F�@�i�8��E���e�f1�����85ĿzGڿ �濦*鿠G�7v��?�~�翁!�H���ҿ����𣜿����rW�h>���9�Q�I� \m�����G���ȿ�/ݿ,��A�#���k�����[����i+�g8Ͽ����ۗ��)z��R�K9<�O
;���N���t������ѱ�؋̿X�߿�T������*�.(忺�迖��h�޿�˿$��%֒���q�2�L��S:���<���S�}��������5�п>q⿊��=��&^�Y&俬��5����ݿVȿ!J��
^��O
m�A�J���;���A�A	\�ꃿ"���Yڼ�N�տ�W���+B鿅��D�z6�k��?���ۿ��ĿmH�������g���H��=�0F���c����`}��]E¿��ٿ>�����1|��K�Be�*��D��}P���ؿ� ���9��M#��sc���F���>���K�!Wl�
s��LN��әǿ�ݿ$�_�쿻��l����F2뿈�����5sֿ삽�v��� ���_���F��5B��~R�t�u�)D���[����̿��῀쿕V�i�m��5�Ӌ���M��Tӿ�0����$���Z��QD�z!C�>�V�R�|�|���7㵿=�пR��)t��쿹-鿊[�z^�����9�F�⿁NϿKF��\��/`z��U�t�B�W�D�]�[��s��}~�������Կ�����=��迡���&;�z뿈g࿔Q˿:���d���*Cs���P�6�A�o�G���a�z���Ă��)����>ؿ���k��*��+r�N�翋��Y���꿴�ݿI2ǿ�ͪ�w*��1�l��OM�{�A��
K��_h��A��ș��$SĿ��ۿ�  �  �$��!��f����a�v�Ϳxo���4��r���nD��qh�yE�E�(������k���E.���L���p��������0⭿
o��q�ҿ���܇����5�"��/$�t�՞�%sݿ���n���9r�)�j��D���֞�?dȿDu��^�[!���$�����'�ZC����ݿ�ƿ{+��U���⓿�&��Q�\� ;���!�};�:{����7�`jX�*�}�đ����n8����Ŀ��ڿ�a��+�_N�`y$���!��Q�Ѐ��jOͿ����N|��B�k���o����㋫��Sؿ�D�-��'�#�;�#�o����	��(�k0ֿw?������#F�������Ew�]�R�b�3��+�K��ئ��.)�.�D���g��↿�f���D���r��5Ϳ�����I���� ���%�
�����Q��1.���*�������m���|�cЕ�n���ʋ���{|�C$&�cp"����^��-���Bп�%����4O��o��U$n�K�J�'�.�[����? ���4��S���w�%������_�������;ֿK`�1D	�4��E�$���%�������nb�3���@����z��rs�͖��W.��پ̿b������D#��'�����J�7A �q7�_˿�T���4��F���l>����d�U%C�*�)T������'���?�`�`�u���ٕ��8���W�� �ȿ4߿=����F��l���&��$�ku�%� ���ѿ�ꦿ]���c1t���w�S*��;���r.ܿ/!�w\�5�%���%�-��܆�v���:�ٿ�Ŀ�㳿����_ᑿo�}�_�X�r�9��K$�?��1��)�.�1<J�m�Y�������⬿���u�Ͽ�\�Z�����0M"�=2'�� �g��򿆠¿���i^���dr�����,��eʽ�ح���8~��  �  ��k�[�b�-J���(�����տຬ��Y���r���N��m0�t �'������龑u�����_�Q�6�loV��{��8��@ڴ��Oῢ>��|0�o�P���f� rk��h]�J�?�'q���n���������Ѥ��p%ҿ�	��/���Q�`�g��k��,\���?�^D�8����ƿ��������wf�M�D���'��k��3���*��+�K������$��A�%8b���������¿�i�Y���;��jY�&j���h���T���3����]>ؿj"��6���g���N�����;M��<��[��k��Wh��(T���4��Q�.�翱繿�����j&\��3<��>!�������|��6���O�D���0�ƭN���q��v��&٪���ҿj����%�`�G�'�a�j�l�f�d�'�K�}(�u���-ȿ'������\����¿['��=$���H�;Lc��@m�8d�kK��*�@b�G�ؿ�q�����x�{gT��6����^�	�˪��L<���� �q&���"���=��A]�=T�������Z��h�俔���82��jR�JCh�*=m��C_�}�A�Vr�L;�9���d䛿�T�����9�ֿ����1��S�Ѯi��=m��S^��A�d�%@��d˿(H��bǋ���n���L���/�2������\��i[���=�#8��,��*I��cj���m���V'ƿ����r���=�t�[�vGl��j���V���5�K��"�ܿ�j��8���zƙ�ֵ���4D���=�8�\�3�l��j���U��f6���a�L��7y���m����b�T�B���'�L����ŗ��p7 ���tv��-6�T�e4w�=���r���/տP��u'�=�H��	c�tn��Ff��)M�I[)�>���ʿ�r��
m�������ſ�/ �&%���I��Od��  �  (
���<��+��;:Z��m&������ó��	��j�U�� -�l�����w׾U>ƾ�i��ɾ]ݾ
�������5�2�`��d��G��2�̢1���e�`������̞��Y���ڀ�M�����x俘�����t<̿=@��^5��k�]���5���N��T��$�|���H����b�ܿWn��+�z�;�F���"�qb�<��s'Ѿ��þ?þ��ξ������4��B�U�s��:����Կ���/�B�a�v��V��^����	��@z���p�%;�$�
��VѿR�����L�ݿ`��G�CT|�M���8����+���_��7"l�,�7��>�e�ǿ����r�h��;����#�b��N�Ͼ�Ǿ��ʾ6�ھ�}���o�A�,���S��
��|ܯ�R�!��OU�����+1��om���[������`���*�}@����Ŀ����H����V��xx%��<Z�K���%��������C�����[���'�E��5{��rÊ��
[��2��{��K �;I�mSҾ�;˶վ��iY��d���;�1�g�mᓿG�ÿ���Sa3�ڷg�Eɋ�Fʛ�����J��^ց��O�������d���a���пnt��7�[6m��t��TL���c���g����~�b�J������࿽���ec��	)O�L�*���������_�,Ծ�nӾ],߾�9��i��Y'�}?J�v�{��Z��uٿd��<�D��y��f��H������I�����r�9=������տ�]���d�����L���I�sA~������m�����8��e�m�Ti9�8�	�˿���XQo�{�A�A@!�K�	�7U�ܾ�Ӿ*�־�u�wY�Z���%2�13Y�N����v�����uF#�ޠV������ڗ����� ��\���'Ma��,����\(ǿ����"ÿ>�����&��U[�]>��U����  �  Z���a������$��eH����9#Ŀ����6L�/�7�����Ӿ�ù�La��ot������ߠ��½۾sK�Y$&���Y��q��a�ԿK��DW�ȶ���B���o���N���x���̟��(}�AU;�7���տ�@˿�Q��"���^����y�����1���`��i.���u�΄3�_���.[����y���:�3���ʾ׌������@��e����ZǾ�龉6��5��q�B���Y��:�,���m�h���=e����������"��\��k;f�<�'�+��S�̿n ҿق���4��u��b��AN��	��������P��R����$_�  ��~޿=��
c��,��m	��5侚�ž���D��0(�����۶־����`����I�b���@P����GB�҂��W����������ۡ�����ހ��zAQ����^�心�˿��࿶���/J�#Ć�k���q��N��Uǽ�HȦ�LԆ���I������ƿi��ضQ���"�V��o߾��ž�u���ϳ�}]���˾�辁��,��`��혿6Qؿ�?��Y�����#���R��N8��m���̠�5?�+|=�m8
��<ڿ�Ͽ�����V$�xa�E�������;$��M�������&@����w�à5��������������B����a��h�ھ@�ľ#ݹ�eA����¾}�׾W��[�B=�	>y��������!�.���o������t�������-��/6���3��fh��*��k���ѿWֿ��ſ6���w�5^��u=��<��������*��u����`��!�e��i����i�3a3�1����uҾ}_��.��R⻾#ɾ��ᾦx���!���N�9��>����(
��C�z��� ���P������LE��.������oR���M�3�Ϳ����bTK�BS������l����  �  �L��G���?c�������b��2�Rӿ[���Y[K�
��l�3%þ4	�������3��^䞾����I�ʾ6����� �^�Z��G��.翧Q+��s�g��o���s��t����6��ֵ��ӏ���S�����K�޿ 0�Xb6���|�l���f������{D��ב��d��������I��
���`���7���
��_ݾ���:���C������녣������Sؾ��$Y1�k\u�·�����w�A�[����޻��Y���T������@���?���U/=��-	�B`�i�濼��4�K�\m��*��n���m���(������ڥ���|��3��_�Eڣ��e��'�}��bӾ`ĵ��"����������v��/ƾQ���T�G�d܋��̿y�[*[�MƔ�c,��&������L=���w���m��W�l�J*�r���Ǜ޿���H.$���d�0 �������d��R���"V������]��}�c�H��9	ֿ_w����P�ɜ�l����ξRص��Ө�����H�������.ؾ�$�'�X�a��ß�`���-���u�6H��Q���X������Y.��~ڶ�v����U�v���� �5k��8�w�؞��W���X/���Y��E�����^����L���G���8Ӄ���?�~	����\ʾ�r���v���誾@���[2Ǿ��辸�[�9���}�����n	�\D����+���x����i���f�����Ϲ�����N]?��]�F��� ����N��w����� ����S��������)���e�~���4������:����k���.�$9��5�ZU¾�l�������V������$?Ѿ.|���u�'M�	z����ο����w\��m��QԺ�����Q��-���V������!n�r+�4 ���࿉���Y%�(�e�G�������j����  