H   E���}H@                        m��b�@                        �%�J6;@H      �      �         �  Hu������g���z����t�d(���޿���ޑL�Yl����ʸ�~=���둾�k���"�����| ������	�]�J���٠���8����J�����,��%�����-��|���rd��"�.�����o���7D�̽���J�����l����l��~W������4��:�Y��G�,^¿Dǂ�u�7����-�Ծ�W���&���$��M����S��q����5Ͼ����0��az��c���~�@�P�nC�������0��\��*��n���Բ���E����K�j������v���[��ۖ�����'W��Ţ���,���������A�b� �(��aj��x(������!ξ���X����~��p�������-¾aI�	���3L������`ؿ��"��m�e����_������OY���(��V �����������7��������G��1�&x��G��Y��T6������/U�������զ�
�w��+��[���#�W�����%���Ͼ����������K�������D۾�����,��kk���ϝ��g�;�*���kȰ�|������������������֝���h���&��� �H���O��H�i���}��}������ ����}��N@���S���$^��v�ޭʿ�	���+H��E�mH����оY�������b鰾�����`;P�����k!A�f��ģ��ä��(U��\��d����P��_~���N�������ܹ��q����O��y��i���^���� �`�����e���@��ur��u�������ۻ��!ʊ�BaD��V��ر��w�M�5����9���Ⱦ]����T�����:��`ؾ̀ ��j!�$�V��Ö��ݿ/�%��*p������������7����f���T��V �������:�
��s�A���d3�7_z�o���w��jI���  �  �����������\��_�j�a"�Hؿu����K�����O辠��:���������M阾���Z#ƾIO���3 ��Z\����u�W�0�o�|��y�������������I��s���-���%[�/o�����㿯���v<���Oë��^������2�������CǸ�ܾ��?Q��&�>����9���8�O�	��پz�����Xϕ�~7���0��x��#AԾ8���W1���w�F
�����%�H�����w��Ƈ��t�������rz��&����b��TjC�4��&�b��=���R�,���>���߾���-���������;K��<Q��>|9�����覧�g�h��v)��+��?Ӿ�!��]_��d ��c^��Qu��nRǾ� �l���K��v���ҿ���c��Ś�����-�������d��,J��Hѣ�W~v�/�0�67����e���MW*�d�m��\��`����;��=��}4��'���m����bm���$��ݿ!����V��!�����m�Ծ-����������_����¾/f�	���-��j��ҥ����Ax4�� ��y<��]���2����c��u;���ľ��O���_�� �������P��@�kF��<�������7��������������ݒ��LU��U��ſ�|���yH�b.�F����վ�s��3,��u��������~Ҿ_�����=�A�&��@J�����m�L�$ ��2���v���������������"������b�G�y>���������{-W�c���j���v�������A���ub������J��V�<��> �rW��S�u�A�6�������ξQļ�����ť��'0žG�ݾl��:#��mV������׿����kf������+���U��O��T���`����x��3����y8�uC���,��Bp�?�������EM���  �  ��f3���I��2���]O�����LȿSW��G�L��:����wϾ�[�����˦��\���{��e׾L��w�%�::[�����E�ٿ E���^�����ٿ��:���r�������(ѥ��8���A����ڿ�tϿ�q���G'���f������!���s���/���ҽ�����~���9�a� ��ȱ��x|��-;���z�꾎aƾk���㐤��ꣾ6ĭ�Y�¾ox徹��!5��'s���������M2�|^v�WF���)��QA��	y��/Ӹ�����`n��6-�I6����пBֿ�N�:��u~��M��iZ�����N�����P:����g���%�����g��"yf��e.�z
�\�例�ž���� ���DB���l���dؾ� ���ܒM�����HĿײ���I�5��g���/��1���x]����������Y���]�ׯѿF�翊�S6R�8E���խ�����|n��֐��>����h���R�*d�t�Ϳ	ɑ���W��X'�<��&���˾�����;��1A���.Ӿ3�� !��:3���h�盞�����!�^`b�V���z���}���R���tm��ԧ��Q��� F��J��r㿪^ؿY����+��Pk�@+���Q��T���NY�������/��`e��E�=�r����.��țK��r!�/������(оe�ľ$Cľ�ξ�H㾛��W^�+yE�Ɂ��Ĳ��%��by6�O�z��b��mI���c�����8����̜���r�'�1����aٿ��޿*S���>�H���D��&8���Y���7��]η�s��r�j���(���뿄����s���;�[�[���4�޾G̾�ľ�Ǿ�,վU�_�7�)��X�Y%���4ɿ�E��bL�5Z���4���}���?�����&��R���[�����&�*Zֿ8�쿤h�9�T�ff��[�������  �  �����ݝ����K�a��+�f�������y���RV�ց,�y�,.��Ҿ�1��]E���.ľQ�ؾ ��7���4��Cb�$G��=Ŀ���j|7�M2n����D����Ĥ����&����HT���0�c���	����п�
�#�;��s�x���5���C��<Ԙ�����O�M�T�ῼ;���}���G��\"��C��N�;j����þ���ʾ�i�l}�j��{B��u�����]�ٿ���fI����鰖��}��2��nǔ��Zy��NA�����տ�E9�������N��݂��K��3���s3��?Β�u��E>�݋��̿ş��
l�u!=����n��de徹оfǾ�˾�|ܾ����n�*�/��2X�-9��˴������'���]�z=���@���ץ�����G���i�P~1�"���ʿd���:�ƿ������+��c��B���w���P��>��dL��8�d��f.�6! ��s��X뎿3Ma�8�7������_�;پ��ԾyJݾ�p�m*
��"���B�{	p��9��7˿S
�_�:���q�rȑ�(v��ؒ��&՜�`���2dX���"�X��+HĿ�廿��ٿ�����?�q�w��֔�	F���m���������s�S�ă��V�Ջ���ʆ��#X���2���������\�߾�߾{ �W��k����.��R������訿�E��<�M�z��|И�E����������}���E����Qy޿����z���>뿄3�R�ʄ�� ���i��[���z��^x�:�A������ӿ�P��{_y�=EJ���(�}�uO���q�D@߾����E�8)�<S�=e:���b�wi��K��	��h�*��>`���������$���ߡ�C��$k�F�3��i�,�Ͽ�j��wZ˿p>�W.�(Me�uU�������  �  Kt���j���P���-���
�W�ڿ���������dt��xO�%0����]�f�������5F�R����6�F~W��~��0������濽V��<6�o�W�M�n�S�s�nXe�'mF�mT� j�p��j̙�i�Ʌ���-׿/����5��EY�W�o�ܗs�� d�_F�%"�~R ��˿����HA���Sh�)hE���'�А��q��^�龿��sW����}$�)�A�{�c��g��7꠿e�ſۀ��K����A���`�{r�%q��H\�4�9���nLݿ]�Jy��v����	��R ����B�ic�8�s��q���[�C;���v;��}��f=���U_�l~>��"�F��?��)��������X����3�o�R��8w�A䑿�d��f�ؿ�����+��6O�J�j��-v��n���S�ɏ.��~�*�ο۬��r���ۢ�Bɿޮ��z*��P���l�w�ɔm���S�P�0�_h��	�:�m���_���Z�1x;�Ȟ!��$�)[�2\����u�;�(��KD��e��兿>$��C���������9�if[�$Dr�L�w�}i��IJ�tX#�|�����¿/k�������E��.�߿bQ���9�	�]�@t�0�w��Mh�KaJ��c&�P��Bzӿ$��$�����x���U�S8����l�E�x������K��4���Q��t������)���οg� ��"�H8F�;e���v��Ju���`���=�{:�-��u��5���(�V�����6���gF�(�f��lw�(qt��P_�j>��]�8)����Ŀ�Ǣ�r㉿�xl�TlK���/�����
�Or����"�[%��>��t]�ހ�������޿��^s.���Q��6m���x���p��xV��1���	�WZӿD`��ⴛ��x���Ϳ����,���R�`�n��  �  ~�)�� &����
�+H�͚ѿֿ��9����Û�'Ԉ�"1j���E��?(����ձ����.�*cM��.s�oX���q䰿
¿H+׿5��?�;n�W(�wv)����b�
��㿮z�����wit���l�Ã�ך��	ͿOn������H&��6*�K�"��P��j�㿸�ʿi���<꧿-!��&����L^�6�;�%�!�Pi���/G��7�,�Y��W��/ԓ��ĥ�4c��WRȿʚ߿����}!�ˠ)��	'���M8���ѿ[��ޅ�}em�yq�7狿������ݿ:N����<�)�֌)����Q�&���ݟۿ=�ſbz��ѻ��vs��^�{���U�)�5�����b�hq�x�+��*H�9�l�h!���^��ݮ�󞿿z�ҿ���������y�&��,��y%�������Lƿ�rQ��{�s������2���������'��$��,���(��u���	�����׿�*ÿ�i��sB��h����u�BQ��4�F�!������%���:�gZ�[<��G��xӦ��ط�dɿ�%޿���&�����N�+�^-���"�	_���.����^��������}�[j���L�� �տ��>���*���.���&�������4Mӿ|����,���W���㊿*�n���K���1�m�#�+�"��s/�k0H��j��z����������H���6�п��^v��R��B%���-��N+���S��)�ڿ�᭿�X��M3~����
���綿�����-!���,���,��?"��l������S⿓�̿�.���a����\V��Ճb��PB��,��Q"��$&�X!7��bS���w�������������Ŀ�ؿ ��g�	��e��{)���.�#(�c�������.˿[U���	����|��*��U���U,ƿnG��)�˶&��  �  ���� ��4����+>�ί��!꿎
ۿ 0¿���Kǆ��p^�lA���8���E�$�g�7�����"�ȿ�߿�=쿛�������,y�??���l����׿᷽��X��h����X��>�:��J�իo��$��{��?Ϳ&�������2:����5�(	�}��濇+Կ`븿�h���}��BS���<�5a;���O��cw�a����i��TGѿ�
������3꿶0运Q�%�����㿖�ϿBY��_픿t��ZM��m:�:!=�P<U�<,������U��HzֿB���=�fJ�0~�I,�����Z𿇹�Y��}Ϳo���;���oq���M�ϊ>���D�4`������ ��8t¿�OܿҺ�ao������`2��_�i��b�w,���ʿ�E��������m�4EM��mA��MK���i�����Ȫ�D�ȿ,l�B� ���~��	�x"�ϩ�9��_����X�ǿ�Щ�J����Gj�[)M���D�lR�)[t�T��������IϿ�j�^1����A�򿇓��f��+����������߿�7ſ���n���3i��O���J���[�Lt���̚��'��G�տ9[�j/��b�����(�Т�@g��8�����aܿm������Ɵ���tc���L���K�i�_�ʃ����0����qٿh>�?L���Q��������z��b���l�nؿO޻�>l��u��k^�K�rM��7e�����&$��ʢ¿��ݿ������t���@%�Z��Ǚ�{��zn��a��yԿ@��Ҙ��}�KZ�8zJ��P���k�疌�Q�����ǿ(���񿅖������$��Zi񿛠�����O���k_��Ͽ�J��$q���Nw��V�(�J�kT��r�Zw������ Ϳ�q��  �  �í�9����ҿ�������k�&�d�)��J!��G�\=�}���ȓ�`cx�k����D����ĿD���fI��R$�F*���$���=���翭Aο�4������&���ⅿ�kd�l�@�%�������GO�;?3��S��Xz�א�+"��賿�gſ�ۿ�U��$^�N �/)���(��,�Р���ڿ�����~����p�
�n�q��������)տb��<�T�'�	�)�` �z*������޿�ǿ�;��r����t��x�}�D-W�c�5���������r#��>�^�a�K����8����-ܺ��Ϳ����� �=$�d+�:�&�M��p����s̿򹡿�ބ�q���z��O������[�迧j��j!�(b+��_)��R�����Y���RٿY�Ŀ���Ԛ�������x��tS���4��� ��x�����3��Q�/]v����#
��KD���+Ŀ�YؿGx���
��T��A)�c�,��$�������X������9���:w��;�����S<˿6@��΢�޽'���-���'�m�����$��
1տ�.¿I���UM���O��v�s�N_P�G5�9%��|"�+=-�iUD��#e�#ͅ�jz���ë�������Ϳ���� �&��/#��V-�Լ,��G ���
���̩��S���C�����������EݿI������+�Ѭ-���$��T���t�؃Ͽn��������0a��-h�"�F��c.��n"�P�#�B�2��fM���p�����<��o�����0Կ��u��\��s'�i.���)����r�#�ҿݧ��ꊿ�}�#R��p��9Y���h#�N$�h�-���+����������-�޿b�ɿʸ�{ϧ�%&���j���X]�U�>��D*�'�"�.�(�&�;�j�Y���~��)������  �  �O��Do���eݿ�����/���R���k�Ot���h�u<L���%�D����������bĒ����aͿ�}�B�.���S��7m�*@t�Ҩg�&�K�v(�Hp�W�ҿ������Ksn�ʓJ��,�6���r ����I���x���	�uY �r�<���]��タa2��^��d(�G>��X<�{�\�q���r��9a�H@�8��mj�����o��r���P����?ΏV�/�;�I^�B�q�Rr�T�_��@����$��'=ÿ����ᄿ7a��1?��}"�\��Aj���@����
�����1�*���H�u�l��ԋ�>⧿�Ͽ�����$�޺H�q	f�׬t� �o��sX��P4�R���,ֿ���E����a��;��K���_�"���I��<h�&�u��o�`X���5��1�s�E}��6;��n{��[]��=�<9"�w���e ��p��u���t��� !��;�Z�[����tЗ�������$A���2�u`U�C�n��	w��k�'O���(�nM�ӭǿI���ܘ�.��1�ӿh�
��2�|-W��p���w��%k�N O��+�����ٿ-���.����|�/SY�R8;��"��Z�O	��]�P�����fn1���M��2o��~���ɤ��ǿ�����z�9�@�� a�@;u�ww�!Te��]D����7��G��'��!�������-W�xd��@��)b�<�u��<v�P�c��CD�g$ �I���ŭ˿�w��DY���r��P�B3�F-�$��P��S���Q� ��X9�USW���z�$���V�����տ��W8(�L�sei��x��8s��[��w7����Aܿ����/L���ſ/�����%��L���j�?}x��9r��Z��8�����\�ƾ��9z��v���Qg�$G�s$,�G���	����������ܶ)�>+D���c������  �  �i�����,I����.�=�d��9������X���i��T���ߍ]���&��O���O�����M�ȿ��PY2�g(j�A���P��Ҥ���������X��c#���j���惿��N�'�[�
�Ռ�1Tо
������r�Ǿ�޾o�D��.�;��l��~��I�οlO�ǋ@��Hw�n���Na�����@��>P����J����}�߿�����`���hٿ�f��D���|�@���xa��N0�������|��`F�,��տ8흿�q�+�?�}f�F�����wɾ���v�����Ͼ5R�
� &�zjL������T��Tq�߻�q�S�f���|'�����+���Q��0�q�7�9����(vп����ǎ��h𿅌"���X�����ޞ�������l�����l��J6�m6�2lĿ�����f��Y:�c�����s���Ծ��;�/Ծ	)��h�U����8���c��ꐿL���Og��H1�ܡg����������Y���Ϟ�����`���)��Z���aƿ������ο�,�w5�Wm���������
���mA�������J\���&�����d�������V]��+6���ì�R�ﾗ��z�޾�>�y( ��� +��#M��E}�S���׿��g�D�[}{�L����t���.��R+���Z��O����������u���}�^r�h�H�zV��;���m��-?���×�}����J�S_�{G޿�^���L���P��/-��~��
���̻޾}3�ks����ԫ��@4��QZ� j�������j"�~�V�!X��"ӛ�2���K�������\�t�-�<����pֿ�뺿z�ſ�Q���x%�N�[�C%����������;��������o���8�@��+�ɿ������p��D���$����GD�����Gu�6=澹���0��xR"�|�@���k��  �  K����b̿���D'S������&��X��g����������CL�b4�y�࿐�Ϳ7%�,4��9[����i���<��`���d:���L��0��MXD�e	�۴��]��h�C�C���
˾#l��~���A��_t��G�����޾�-�*�-��?g�����1过<(��j��Ș��7��S�����������k��@�z�$f7�a�gEտzҿ�� ��0��r�R����M��#������,���s��'lr���.�>�������~n���1���
�b�U����Ѭ����0ޥ��U���aʾ�{�9���[@�ˁ�2ƶ��O�s�=�X����9��i��m����;��L%������+d�l%�\��5-ѿT߿���I{F�����J��c������������b��տ\�9����ؿ�[��&�^��*�;���K�ƹȾ7����V��a����Ⱦ����
�q�(�o�Z�va���ѿyr���U��c��nM�������|��H��e�������JO�?@��翓�ӿ5��=!�uK^�D����������(�������i�����6�G�̉�~�ÿ�&��(+R��I%�������ѾS�ž��þ�̾�<�ph ��4�s�>�W`x������9},��n����8N��g���c����}v��Y�~�>t;�V%	��ZݿP�ڿ$��U�4�@�v�W���wW��(��E�������������v�03�0��l��Y�5�B�����������>;��þH$ž��оd:�f���#��:N�6���h|��r��*7A�L�����������7���$�����g,g� f(�BM���!׿�
忊���qI��U��@���[����#��-��x^���2��K]_�u�H0޿����5Ii�}5����,���,ܾ��˾��žڐʾ�ھ����]�^�0��b��  �  穔�]#ݿ��%�o�D����h������^������۔��	��_ng�!
%�/j���n�+����1���x�b����������Ur��;�N���k�]����y~ʿ4��h�A�m�� $���������Ʃ��=������2 ����;�U ��(�Ej��˩�������<�CA��r%��X ���;�����F3�������\��K7O��u����;�O��%|G�jʉ�C��k(�����j����3_��Ǽ�� }D�ܣ�:�΀r���-��F�R;Ѿ(E���l��v��Z4��,���S����y߾���6�=��%��,4ÿL��V�Vo��5:���R������OL��B1������l�� :�� ��B�����{ ��{`����l���O��W�������m���{����y���.�cI�a���~_��%�� �Ծ�b���r��࿤�����S���oӾm���c�"�fZ�Q+�����fp(���q��������BO���N���L������q���|j��(�����$��K����4���{�㎦��������`��P%�����eN��30a�aY��uѿ@��8P�q����f�ؾo�������������!�Ͼ�uﾎS���9�� {��X��D���@��^��l?������N������@��c���e��OES�g��0��P￞����K�ы��J��2�������x��X$��Gs��wӋ���H����Y��������>����+Z�{Ѿ׼���D���Z���#���E׾�|�����FrK�O���ɿ�k�f\Y���-߼�J���RM��%���:���9���l���=���
�J6뿖����|#��yc���������R�������= ��vL���h��h�|�ȓ1�|��@R��j�i��d/�y�
����_�˾�o���@��ʅ����ɾ~�j�$�*�0ab��  �  �A������&,�݆y��ܧ��`��=��
u������=&������}Vq�P�+��} ���eu�T9�v���4?��(��q/���@���k���j��6b��IDg�{��}п�+��c�A��s@ܾfִ�.���C���"���A��g
���Ⱦ�_��S(�s�k�p����A��qD�0'�������r���������������������W����I�W��<��[�O�sȏ����ʌ��e����������bk���܏��L��<	����v�t�x<-�;:�L2̾~2��>���,䐾��͝�m��ˊھ��am=��Ն�tBȿj�!_����H����/���9������H����U��w�A�z��n��������&��i�'�������S����������g���l����5���
��@�`��#����l�ξgZ������
 ��QǤ��S���Iξ����=!�%[���IS�-�.�iK|�Q>��a����~�������;��ɡ���E���gt�ե.����;�!x
��<��9��iǭ�����x������������3��γj��	!�K׿M7��-9P����A���SӾ����3ʱ�Ke��40��ehʾ5T�`*�>9�}���������H�_D��k������������������������[�_"��^��b��������S�	ϑ����n���0���Y�������c��V��Z�P�q� z��ق�>�m���I��˾r㸾G�������r:���!Ҿ�����#�FK�ҡ����ο����mb������M��F���"���������S��i{����D�^�������)���l��2���?�������l��e���n��jخ����ix8�e����B��Ek��.�s�������ƾ]�������ȶ���ľ�V߾Y���^)�> c��  �  穔�]#ݿ��%�o�D����h������^������۔��	��_ng�!
%�/j���n�+����1���x�b����������Ur��;�N���k�]����y~ʿ4��h�A�m�� $���������Ʃ��=������2 ����;�U ��(�Ej��˩�������<�CA��r%��X ���;�����F3�������\��K7O��u����;�O��%|G�jʉ�C��l(�����j����4_��ȼ��}D�ݣ�=�рr���-�F�:;Ѿ�D���l�����3�����������x߾����=�C%���3ÿ�OV�5o��:���R������7L��.1������l���:�� ��B�����{ �|`����l���O��s���������������y���.��I�����_�D%�^� ��ԾMc��=s��忤�؂��KS��-oӾv��ȭ"�ReZ��*����%p(���q����]���!O���N���L�����uq���|j��(����%��S����4���{���.�������8`��r%������N��y0a��Y�0vѿ�@���P��q�5���Q�ؾ,�������%����_�Ͼ�uﾝS���9�� {��X��D���@��^��l?������N������@��c���e��OES�g��0��P￞����K�ы��J��2�������x��X$��Gs��wӋ���H����Y��������>����+Z�{Ѿ׼���D���Z���#���E׾�|�����FrK�O���ɿ�k�f\Y���-߼�J���RM��%���:���9���l���=���
�J6뿖����|#��yc���������R�������= ��vL���h��h�|�ȓ1�|��@R��j�i��d/�y�
����_�˾�o���@��ʅ����ɾ~�j�$�*�0ab��  �  K����b̿���D'S������&��X��g����������CL�b4�y�࿐�Ϳ7%�,4��9[����i���<��`���d:���L��0��MXD�e	�۴��]��h�C�C���
˾#l��~���A��_t��H�����޾�-�*�-��?g�����1过<(��j��Ș��7��S������� ��� l��@�z�%f7�a�hEտzҿ�� ��0��r�S����M��$������.���s��+lr���.�E������~n���1���
��a����~Ѭ�8��Kݥ�VT��k`ʾz���bZ@�Pʁ�^Ŷ�O���=����D9���h��7����;��&%��璕��+d��k%��[��--ѿg߿ى�o{F�����=J��7c��8������������U�\������ؿ\\����^�N�*�0��;M徿�Ⱦ�����V��󉸾��ȾQ�� 
�F�(�
�Z��`��"�ѿ�q�-�U��c��,M�����R|�����d�������JO�#@��翕�ӿ25�>!��K^�c����������b���4����������G�K��i�ÿk'���,R��J%���E��J�Ѿp�ž��þ��̾[=ྙh �5���>�b`x������9},��n����8N��g���c����}v��Y�~�>t;�V%	��ZݿP�ڿ$��U�4�@�v�W���wW��(��E�������������v�03�0��l��Y�5�B�����������>;��þH$ž��оd:�f���#��:N�6���h|��r��*7A�L�����������7���$�����g,g� f(�BM���!׿�
忊���qI��U��@���[����#��-��x^���2��K]_�u�H0޿����5Ii�}5����,���,ܾ��˾��žڐʾ�ھ����]�^�0��b��  �  �i�����,I����.�=�d��9������X���i��T���ߍ]���&��O���O�����M�ȿ��PY2�g(j�A���P��Ҥ���������X��c#���j���惿��N�'�[�
�Ռ�1Tо
������r�Ǿ�޾o�D��.�;��l��~��I�οlO�ǋ@��Hw�n���Na�����@��?P����J����~�߿�����`���hٿ�f��D���|�B���za��P0��
�����|��`F�$,��տ@흿�q�,�?�qf�)����-wɾ���8����ϾP��

�� &��hL�s���kS��p�4��ÇS����*'�����������ۆq���9�����uп����㎿�ah𿻌"�5�X�ￇ����e���X��ò��:�l�QK6�7�qmĿ����ܕf�\[:����������͆Ծ��;M/Ծ�'��g���?�8���c��鐿	����f�%H1�"�g�����+���TY���Ϟ�W��;`�t�)��Z���aƿ������ο�,�Cw5�kWm�Д������Z����A�����OK\�S�&�(��>f�������X]��-6�S����L��#�ྦྷ�޾�?��( �I�"+��#M��E}�V���׿��f�D�Z}{�L����t���.��Q+���Z��O����������u���}�^r�h�H�zV��;���m��-?���×�}����J�S_�{G޿�^���L���P��/-��~��
���̻޾}3�ks����ԫ��@4��QZ� j�������j"�~�V�!X��"ӛ�2���K�������\�t�-�<����pֿ�뺿z�ſ�Q���x%�N�[�C%����������;��������o���8�@��+�ɿ������p��D���$����GD�����Gu�6=澹���0��xR"�|�@���k��  �  �O��Do���eݿ�����/���R���k�Ot���h�u<L���%�D����������bĒ����aͿ�}�B�.���S��7m�*@t�Ҩg�&�K�v(�Hp�W�ҿ������Ksn�ʓJ��,�6���r ����I���x���	�uY �r�<���]��タa2��^��d(�G>��X<�{�\�q���r��9a�H@�9��nj�����q��t���R����?´V�2�;�M^�F�q�Wr�Z�_�@����$��4=ÿ����ᄿ;a��1?��}"�!���i���?�v����z����*���H�7�l�\Ӌ��৿4Ͽ�����$��H��f�%�t�c�o�1sX�]P4���-,ֿ���8����a��r;��������"�^�I�k=h���u�ӥo�1X�z�5�^2�!��~���<���|��g
]�c=�|:"�N��7f ��p���������^!�k�;�T�[�ؚ��ϗ�|�����H@���2��_U�w�n�C	w�b�k��O�A�(�!M�p�ǿ���ܘ�e����ӿ��
�L2�.W���p���w��&k�-!O�Վ+������ٿ���g0���|�\UY�%:;���"� \�;
��^�Ӂ�:���n1�%�M��2o��~���ɤ��ǿ�����z�8�@�� a�?;u�ww�!Te��]D����7��G��'��!�������-W�xd��@��)b�<�u��<v�P�c��CD�g$ �I���ŭ˿�w��DY���r��P�B3�F-�$��P��S���Q� ��X9�USW���z�$���V�����տ��W8(�L�sei��x��8s��[��w7����Aܿ����/L���ſ/�����%��L���j�?}x��9r��Z��8�����\�ƾ��9z��v���Qg�$G�s$,�G���	����������ܶ)�>+D���c������  �  �í�9����ҿ�������k�&�d�)��J!��G�\=�}���ȓ�`cx�k����D����ĿD���fI��R$�F*���$���=���翭Aο�4������&���ⅿ�kd�l�@�%�������GO�;?3��S��Xz�א�+"��賿�gſ�ۿ�U��$^�O �/)���(��,�Р���ڿ�����~����p��n�t��������)տe��?�Y�'��)�` ��*������޿�ǿ�;��|����t��q�}�&-W�(�5�����(��c#��>���a�?����7������ں�=�Ϳ������g$��+���&��������Js̿v����ބ��q�2�z�P��4���/��.k��k!��b+��`)��S�� ��[���Tٿ
�Ŀ����.��������x�'vS�x�4�B� ��x�K���3�1Q�c[v��������B��*ĿXؿ_v���
��S��@)���,�$� ����EX������t9���:w��;��{���	=˿*A��g����'�T�-�� (�a��������2տ0¿⡱��N���P��x�s��`P��5�:%�~}"��=-��UD��#e�6ͅ�uz���ë�񃼿��Ϳ���� �$��/#��V-�Լ,��G ���
���̩��S���C�����������EݿI������+�Ѭ-���$��T���t�؃Ͽn��������0a��-h�"�F��c.��n"�P�#�B�2��fM���p�����<��o�����0Կ��u��\��s'�i.���)����r�#�ҿݧ��ꊿ�}�#R��p��9Y���h#�N$�h�-���+����������-�޿b�ɿʸ�{ϧ�%&���j���X]�U�>��D*�'�"�.�(�&�;�j�Y���~��)������  �  ���� ��4����+>�ί��!꿎
ۿ 0¿���Kǆ��p^�lA���8���E�$�g�7�����"�ȿ�߿�=쿛�������,y�??���l����׿᷽��X��h����X��>�:��J�իo��$��{��?Ϳ&�������2:����5�(	�~��濇+Կa븿�h���}��BS� �<�9a;���O��cw�f����i��\Gѿ�
������3��0迡Q�6�����㿝�ϿBY��S픿�t��ZM�Wm:�t =�C;U��+��@����T��yֿ���1<�H�X|�m*�'��"Y���W㿞|Ϳz�������nq�f�M���>��D��4`�z񆿯��Qu¿Qܿ[��q������K4쿹a��j�hd��-��ʿ�F��L�����m��EM��mA�MK���i�����Ǫ��ȿ�jῥ�����|�� ���p��ￅ��)�ǿ�ϩ�����Gj��(M���D��lR�'\t����񰱿
KϿ$l�
3����6�򿋕��h��-��Z������\߿#9ſ���@���a4i�
�O�T�J�B�[�xt���̚��'��O�տ;[�h/��b�����(�͢�>g��6�����aܿm������Ɵ���tc���L���K�i�_�ʃ����0����qٿh>�?L���Q��������z��b���l�nؿO޻�>l��u��k^�K�rM��7e�����&$��ʢ¿��ݿ������t���@%�Z��Ǚ�{��zn��a��yԿ@��Ҙ��}�KZ�8zJ��P���k�疌�Q�����ǿ(���񿅖������$��Zi񿛠�����O���k_��Ͽ�J��$q���Nw��V�(�J�kT��r�Zw������ Ϳ�q��  �  ~�)�� &����
�+H�͚ѿֿ��9����Û�'Ԉ�"1j���E��?(����ձ����.�*cM��.s�oX���q䰿
¿H+׿5��?�;n�W(�wv)����b�
��㿮z�����wit���l�Ã�ך��	ͿPn������H&��6*�K�"��P��j�㿸�ʿi���<꧿.!��'����L^�8�;�(�!�Ti���5G��7�5�Y��W��6ԓ��ĥ�@c��dRȿٚ߿&�����!�Ӡ)��	'���N8���ѿ�Z���݅�em�lxq��拿6�����ݿ�M�����)�
�)����l�Z����ۿ��ſ�x��{���Sr����{�|�U�.�5�<���b��q�<�+��+H��l�w"��;`���ޮ�����?�ҿ������t��U�&�|,�Jz%���������Mƿe����Q����s�f���K2��$�������3�$�%�,��(��t���	����׿=)ÿHh��A���f��̊u��Q��4���!����w�%���:�{hZ�O=��w���Ԧ�0ڷ�(ɿ�'޿��� �����1�+�+-�C�"��_����򙻿�_��p���p�}��j��M��7�տ��>���*���.���&�������1Mӿz����,���W���㊿)�n���K���1�m�#�+�"��s/�k0H��j��z����������H���6�п��^v��R��B%���-��N+���S��)�ڿ�᭿�X��M3~����
���綿�����-!���,���,��?"��l������S⿓�̿�.���a����\V��Ճb��PB��,��Q"��$&�X!7��bS���w�������������Ŀ�ؿ ��g�	��e��{)���.�#(�c�������.˿[U���	����|��*��U���U,ƿnG��)�˶&��  �  Kt���j���P���-���
�W�ڿ���������dt��xO�%0����]�f�������5F�R����6�F~W��~��0������濽V��<6�o�W�M�n�S�s�nXe�'mF�mT� j�p��j̙�i�Ʌ���-׿/����5��EY�W�o�ܗs�� d�_F�%"�~R ��˿����HA���Sh�*hE���'�Ґ��q��d�����}W�����}$�4�A���c��g��B꠿q�ſ���S����A���`�{r�,q��H\�7�9���_Lݿ?�y��,���o	����뿵���B��c���s�q�1�[�s;�L�u�5:��"��4<���S_��|>�:�"�e�?���񾕏��_��p���3�U�R�
;w��呿;f����ؿY����+��7O��j�J.v��n�{�S�2�.�"���ο���w���ۢ��ɿ���#z*�p�P��l�Yw���m���S�q�0��g�࿰촿�l���]���Z��v;���!��#��Z�B\�����R���(�@MD��e�8煿�%�����̘������9�Fg[��Dr��w�i��JJ��X#�$���|�¿�k��Ȥ���E��K�߿jQ���9�	�]�@t�-�w��Mh�GaJ��c&�N��?zӿ"��#�����x���U�R8����l�E�x������K��4���Q��t������)���οg� ��"�H8F�;e���v��Ju���`���=�{:�-��u��5���(�V�����6���gF�(�f��lw�(qt��P_�j>��]�8)����Ŀ�Ǣ�r㉿�xl�TlK���/�����
�Or����"�[%��>��t]�ހ�������޿��^s.���Q��6m���x���p��xV��1���	�WZӿD`��ⴛ��x���Ϳ����,���R�`�n��  �  �����ݝ����K�a��+�f�������y���RV�ց,�y�,.��Ҿ�1��]E���.ľQ�ؾ ��7���4��Cb�$G��=Ŀ���j|7�M2n����D����Ĥ����&����HT���0�c���	����п�
�#�;��s�x���5���C��<Ԙ�����O�M�T�ῼ;���}���G��\"��C��N�;p����þ���ʾ�i�s}�s��#{B��u�¨��g�ٿ���fI������~��5��qǔ��Zy��NA������տ`9��^����tN�݂�TK����'3���͒�Uu��D>�7����̿����l��=�O��d���c��о�eǾ��˾~ܾz��.p���/��4X�B:��A̴�S���m�'�^�]��=��A���ץ�㘠�}���ki��~1�L���ʿh����ƿ\�����+�Jc��B���w��jP���=��	L���d��e.��  ��r��5ꎿ8Ka���7�������^�{:پ �Ծ4Kݾ�q�{+
�	"���B��p��:��l8˿�S
��:���q��ȑ�v��%���f՜������dX��"����sHĿ�廿ۖٿ�����?�r�w��֔�F���m���������p�S���V�Ӌ���ʆ��#X���2���������\�߾�߾{ �W��k����.��R������訿�E��<�M�z��|И�E����������}���E����Qy޿����z���>뿄3�R�ʄ�� ���i��[���z��^x�:�A������ӿ�P��{_y�=EJ���(�}�uO���q�D@߾����E�8)�<S�=e:���b�wi��K��	��h�*��>`���������$���ߡ�C��$k�F�3��i�,�Ͽ�j��wZ˿p>�W.�(Me�uU�������  �  ��f3���I��2���]O�����LȿSW��G�L��:����wϾ�[�����˦��\���{��e׾L��w�%�::[�����E�ٿ E���^�����ٿ��:���r�������(ѥ��8���A����ڿ�tϿ�q���G'���f������!���s���/���ҽ�����~���9�a� ��ȱ��x|��-;���{�꾐aƾn���琤��ꣾ<ĭ�a�¾yx����!5��'s�������� M2��^v�ZF���)��TA��y��2Ӹ������`n��6-�=6����п�Aֿ��*�:��u~��M��AZ��ؒ��������:��B�g�J�%����*g���wf�Sd.��
��來�ž���㽬��B���m��>fؾ� ���/�M�b���#ĿO��j�I�v�����$0��i����]��������͒Y����|�ٯѿ-��o�)6R�E��`խ�v���Dn�����������h��R��c���Ϳ;ȑ�t�W��W'�J���$��˾2����;���A���/Ӿ���"�<3�4i�������_�!��`b������������������m��Cԧ�R��� F�K��r��^ؿ*Y����+��Pk�@+���Q��R���LY�������/��_e��D�=�q����-��ǛK��r!�/������(оe�ľ$Cľ�ξ�H㾛��W^�+yE�Ɂ��Ĳ��%��by6�O�z��b��mI���c�����8����̜���r�'�1����aٿ��޿*S���>�H���D��&8���Y���7��]η�s��r�j���(���뿄����s���;�[�[���4�޾G̾�ľ�Ǿ�,վU�_�7�)��X�Y%���4ɿ�E��bL�5Z���4���}���?�����&��R���[�����&�*Zֿ8�쿤h�9�T�ff��[�������  �  �����������\��_�j�a"�Hؿu����K�����O辠��:���������M阾���Z#ƾIO���3 ��Z\����u�W�0�o�|��y�������������I��s���-���%[�/o�����㿯���v<���Oë��^������2�������CǸ�ܾ��?Q��&�>����9���8�O�	��پz�����Zϕ��7���0��|��(AԾ;���W1���w�I
�����'�H�����w��ȇ��v�������tz��'����b��TjC�1��&�P��0���R� ���.���˾���-������ȭ��K��Q�� |9�E���������h�v)�~+��>Ӿj!��_��U ���^���u��SǾ�!�m���K�Ew��c�ҿ�^�c��Ś�ߩ��N������}��@J��Wѣ�m~v�>�0�>7����X���?W*�O�m��\��M����;���<��[4�����J���bm���$�y�ݿ� ����V�!�������Ծ��������#������j�¾�f྆	�S�-�� j��ҥ����x4�� ���<������T����c���;���ľ��O��)�_�� ���������P�
�@�kF��;�������6��������������ݒ��LU��U��ſ�|���yH�b.�F����վ�s��3,��u��������~Ҿ_�����=�A�&��@J�����m�L�$ ��2���v���������������"������b�G�y>���������{-W�c���j���v�������A���ub������J��V�<��> �rW��S�u�A�6�������ξQļ�����ť��'0žG�ݾl��:#��mV������׿����kf������+���U��O��T���`����x��3����y8�uC���,��Bp�?�������EM���  �  `��������U�����6k��"�+׿E��� NG�Q��b�޾���f)��e)��a����S��uנ�K��K�뾜E�}�W����s��1�Il}�p��<�������o���
��K������s�[�ڙ��������s�<�`���@������p�������t������9���iQ�������
=~��73�l���Pо㬾�6���p��|ߍ��m������S�ʾ_� �|,�uys��w���d��H��x���/��dm��2���9����,��M|��������C�����������JS�b���5��z��3��Ǿ�������������@�9�����p�66d�Ə$�ח���ʾ|Ѭ�+����і�F{��ꍾ�L��{�S4G��w���?ѿ����Qd�eQ��#u��;��[�����������D��w�`1�"B��|忡���;�*�nn��ɟ�rO����=&��?"��a���K���m�G�$�!~ܿ1���HR�@��L��|̾p���J2���T���z��{���uW׾�+���(�Y�e����7�7�4�iw���ީ��������I��l���dW��س����_�K!�Z�������c�U7A�����s��o:��z���g���s���ܧ���W��>�U�+�^_Ŀ`���C��=�W��Y;*���kʮ�w5���ƶ���ɾeh뾍����<�����϶��F���M�����L������:�������_S������u��<H��W�'����6�f�W�2���6��E`�����E{��m@������)a��J�<�r���ӛ��Xzq�D�1��;
�ҋ���ž ��W���54��!3����Ծ�Q���!��Q�q����eֿ�x�Y�f���|���.�����������"���r���]y�(Q3�ߓ�)��J���,���p�Y���l��f���  �  ޵�����Qͼ�����ra�k
��ѿjq���F��{��X�e������Ɠ��C�������å�¾� �p���V����s��M=*���r��ݠ�h��������\������5O��xM��٬R�i���鿜�ܿ�&��Y5���{�����<���������������������H����~���L{���3���w.վ�䱾��������k��z-�����)�Ͼ�� -�6q��U��i����@��|��\��v'��h������8����������;�����ݿ08俆Z���J����1k��AB����������������FN|�m2���%�����b�x�%������Ͼ�ı��m��4X������O��-�þ�R�����F��u����˿�K���Z�I�������������$.��m��)g���l�D*�����n�޿t����'$���d��!��*���Cq��1���k���)���u���)d�L��:pֿp㒿;�Q����6���� Ѿމ���ϫ��٨�R#���x���Wܾ�_�:*�CXd������뿺�-�Gv�����������_4��J���$X���l��<W��=������������9� !���3���k������[����4�����$��a+M��,��̿��煿��C�:�����ZҾ8b��dY������\�����ξS�����a=�U������������D����kx���F��y��������^���5��[;��xV@�TW�����ױ�XO�P����h��l%����������@��Y5������5�q���\G����o��2�Q^�I�辘�ʾ�й�%-��6̵��	¾$�پ� �A��(xQ�ۤ����пD��k�]������a��5*�������n��P���z���Do���,��7�X:��8��Y�&��g��F����������  �  <	��ۀ�����`����UG��c�����c����G�l��?�� �ʾ�����h��Ą��7Ӥ��µ���Ҿ_���]�!��U��D����ҿ�j��1V��-�� ����������{���E���|�$I:������ӿE-ɿ�?�@!���]�a������}���9.���`��«��Ջt��2�����UQ����u�ͥ6�����得^¾�P���f���à�_�������ཱྀ�	���0���l�7Y���N�ǌ+���l�w	���г�aH������h���#����	e���&�n���{Oʿ��Ͽ:Z� �3��xt�$�������������C���_I��]�^�;|�H9ݿ>ǚ�ٙ`�b*��*�A�߾����`��7�����c⺾b5Ծ������H�l4��1�Э�rB�.����@��C�������ݐ�����Xx��)6Q������忰~˿��۱��/J��ǆ�Z��"���a��_޽����V��J���&BǿDՍ���R��#� ����EȾ�p��������� sϾA#��B�YX/��]c��5����ٿ�����Y�����y������M���Jٺ�BF���$����>��^���ܿ�ҿ� ����%�bKb�4���$������WW��t���Ν� �x���6��� ��������G��1��8���⾱�̾���{����ʾX߾D� �b9�pA��}��������t�/�-�p��%��6��tj��t������¯���^i��+�n_���ӿMؿ���=�7���x�8ݝ�Ἰ�U���T��N���I�����a�b�"���㿅u����m�<�7�_��[����ھP�Ⱦ�r���Wľ�Ѿ�n꾣��A&��#S��c��]ÿ�@���D���g����޼��4������(6��o���l�S��6�#��*п�S�c��}L��������*���  �  
s��2���=u���Y�TD%��;�u������0�P��q(�pE�
��Suξ�E��z��S/��n=Ծڰ��mG���0�q�\�/8�������r�0�1�d��a���`��E���Ҕ��S��L�u���a�v�f譿%*ʿ�7�W4���i��ٌ������˝�Rђ�ֈ{���G������ڿ�d���lv��B�#���I�Ik�A�Ⱦ񵻾
򺾈�ƾ��޾ŕ������=�m+o�	����ҿ"d���A���u������s������o�Q�9�i�	���ο���β��Uۿ�x�F��i{�>���-���ԛ����Ek��7����pƿ~e���'f��8��v�����J̾��þҮǾ�+ؾ���tO�m�+�zS�����{������!�= U����c��VW���H���
���_���*��*����Ŀ �������`V���}%��IZ�����*6���Ο�-��ֆ���[�f�'�����'㶿�/��u�[���3�%��������LվYѾ�Hپv���p�����:>�$Jj�)���ſ̙�L	4��_h�����!��K��ϲ��uJ��bP�O����i���g�ҿq�	�\�8�1_n�R���ޝ�����T�������K�������W���;x��#FS��.�a��ip��N��ܾ�F۾`��Q����Y7+��N�f���G��/�ڿ�����E�z�����.��D��� 	����s��1>�����׿�R���Z����ę�J�z?�,�����-���������n��l:�}�
��#Ϳ_��Kns���E�oe%����u����g�Hs۾l�޾������X3�)r6�A�]� ӊ��������W_$��W�$2��,i������ ���VJ��Jnb��?-�� ��qɿcP��qſ�����'���\�Oԇ��>���  �  G�j�O�a�Q�H�H�'�|��\�ӿ�l������	n��CJ���+�������q��$��Ύ� G����2�pR�]`w��������B'߿H+�gj/��O�re��bj�7Z\���>�8d�F �X������c鏿����oп����.���P�|f��j�'[�4�>�H?�T���#�Ŀ��������bb�ʉ@���#��P�����Z��8��p���	��� ��<���]��ׂ��i���ɿ�+�K7�R�:��BX���h���g���S�s2�җ���տ�Ϧ�k��iR������?�㿫W�8%;��9Z�cgj�Ŭg�%�S�;4���l��Ң���՗�ܰ���Y��9���

����>)�S����{���/�5�M�7q�\���w��v7ҿR�e�%��YG��a�7�l���d���K��(�����ȿ�������Y����¿�;���#$���H�&rc��nm�*kd�5�K��B*�k��@ٿ�ٯ�?���y�fU�x67�E%�A�Ԣ���{���M����%�_�?�ݝ_�(���G���K����濣��e�2�yS�_�h���m��`��B�^e�]D�&μ�7��ۗ��KM����ؿQ+�A�2�L%U�W�j�`n��r_��B��| �15 �K@Ϳ�c��G܍���r�R�P��4�,��V�������2%
�����0��M�.@n����j���ȿ�����h�0�>�&�\�m>m�T�k���W���6����v|޿j^���똿�����ͷ��	�pA���>��]���m�sk�9�V� i7�e�qj�V������n|����f���F��+��y��/�#�r��L���!��u:�]X�u�{�?��	���D_׿1���.(�u�I��%d�6o��eg��IN�l|*��'���̿b���ݸ������]ǿaY��P&���J��|e��  �  ѕ#�y�� ;�s�e���:˿1!���觿�D��"����c�~@�m9$�/���r�
����)�'H�}�l��Z���P��f���PD����п��|u�~����!�O #�����GYۿ�ۭ�����n�̹f�c2���Ŝ�uTƿ�f��<W� ���#����:"�/9����ۿH�Ŀ�!��C��ؑ�^7~��uX�L�6������U�u���w3��0T��y����,����T¿�ؿ�����&��O#��� ��&��*����ʿY���5��Tg��@k����(���C}ֿ�l����=#��J#�\4��7	����;�Կ�����>��0��d���u�isP�^�1�S�"����'� HC�alf�=^�����۩�}����̿�`�^{�zf�/� �s�%��^����I�e�����0��Z�m���|�Lޕ�!��������2���S&�r�"�Y���3��/�h�п􌽿�Y���Ü���Ao�]L��0�������!�R�6��U���y����t0������>ÿ��׿���y�	��@�kR%���&����#\	�b4㿇����O����~��w�4Ո��s���Ͽ���ů�jh$��0(�!��f��Y��a�X6Ϳwp���I�����+G��m�h�,$G���-�\E ��~�d�+���C�id����Ǘ�m&���D����ʿ������$=�`c��'�E%�m�F�� �ӿݨ�ܬ���x��{��!��,~���(޿6�P[��&�-�&����<�����Üۿ��ƿ0�%�����O����]� >�k}(����"�513��N�eq�����56��p��9����ѿ]��f�-��i#��O(���!�Y/��E��.�Ŀ؝�ק����v��܂��^��e��<���N� ��  �  ��⿢��`�u6��W῕�����pK� �ӿ�껿O��c��X��e<��H4��A�ȅa�����ǥ�:¿�ؿVZ�����係O�⿫�忐 �.�࿜�п�������%~��ES��=:���5���E��9i�፿����r�ƿ#ۿM�� 翊���a���
R���Z!߿�-ͿK���ϕ�v���M��8�J�6�FhJ��p�0��ʰ��"fʿ"cݿ�#��H�o��s��u��{@�����Hܿ�ȿ��������bm�4H���5��8�(�O�#Ly���h��fpϿ��T�Ә�\�}�⿔e�������ۿ4�ƿ"/���S��kk���H��:��,@��Z��<��� ��IQ��2տf��d��G��;x�H��T��_��(����ڿ4TĿd
�����$�g��iH�=�`�F��d�E:��򱥿�¿ڿ�)迳@쿦��=�������8쿓�翛Bٿ����wˤ�RĈ��td��mH���@��M�0n�(r���a���ȿ1�޿�K뿬��G뿸C���Ё쿋���	�I�׿�#���D��������c���J�F���V�joz�ǅ��꠳��2Ͽm��TD���F쿜��\9뿷�ￅb�$cտc9��g�&$��*^��BH�GG���Z��i��ʚ��Mҷ�a�ҿŕ�#a��[�EH�vK�U�'�����=ѿ�6������D~���X��F�|�H�O�_�ul���x�������~ֿ?���￞@��A�鿡쿡E� ��v�bͿљ������pw��U�vF��K��f�:∿æ��j���vgڿ� 꿊�ￚ	���g���$�￭��9�߿.rɿ���o��G<q���Q� OF�U�O� m�����,奔�ƿ޿�  �  ���������f̿oV�<i�s��f �m�#��G��	���ӊ��{�����q�ce�g=y�����xm�������0���#�av�P��<���bO�iȿh���'���ĭ�� )���[^��;��!�Ml�߂�8��2�.�`vN�>�s�u���<h��.�������'�Կ�.�&n	�D>�<�"��N"��d����tqӿc=�������j�Z�h�ヿ�ܢ��	ο�9��bZ�nf!��?#�����!��Q��L"׿��� 诿濟�I����v���Q�Q1��%�k����wN�a9��[�A���瓿.��Hh��fǿ��޿��������^�$��S �'!����_�ſ]����Z��k��tt��4��A첿�࿙Z�3z��	%��,#�Ժ�{B�����ҿ�ξ��c��������:r�~>N���0�'J��9��R�{�.�;L�]�o��/��@����+�����^�ѿ9�뿽"����!#��@&��
�������e��fy����}�s8q��͂�����%�Ŀ����1<��!��a'���!��@�>F��>�)�ο�������盿������m�R�K��21��!�3�[�)���?���_�\`��%]��T���;���ȿ�Vݿ1���^��Dl�*'��n&�O�����ۿ�Y��������z���x���������$ֿ@-��n�\%�9^'�����K�Ѱ���߿�ɿ�`��?<��Ŗ�Bヿmb�B��*�:'�E� �4/��H���j�3;���隿^��� ���οu����."��y!�m(��#��`�����?̿���Sf��� w��������������W��"�/�'���%��L�t�	���Nؿ�Ŀ�����6���1���P|��"X�g:���&�~���f%��7�G�T�Whx��H��X����  �  �S��EE���Uֿ����s)���J��b�K�j��_�wLD�M������̐��[����Ǝ�G;��b�ƿ����$(��K���c�O�j���^���C�d�!��� ��%̿�.��"T��INh���E�&�'�e���F��z��m���0�H��L����7�^X���~�ᗿ�W���D�����@5�oIT���g�sli�hX���8�I!�ڄ�g���ݒ��q��}H����ٿ���4��dU�!Nh���h��V���8��V���W������N]���][��:�o���j�M�Ob����p����l�J�&��D�=�f�^#���.����ȿ����_���A�+#]�� k��f��
P�{-�
��U9Ͽ�$��_�������\���T���H0B�'1_�^Il�_[f���O��?/����߿�(���$��,e|���W� �8�M��z�
�����Ӓ�1�����	�����7�plV�\�z�
ԓ��˱���ۿ%Y
��,,��FM��`e�Drm�(�b�]#G�}"���������ٞ���ݔ� `��!�̿L���_+���N�LJg�en�P b�sVG��_%��V��ӿ�(���d����v�kGT��7�� ������6��x�������-��#I�(�i�a��v��9���1��r	�nu9��vX�<�k�Y�m��\���<�Q2�Ϡ�����񚿥��� ]��G��f��3�8�zxY��fl�V�l��[��<�:��G]����ſ���Ӊ��Dl��XK�sj/�]�6v	�2�����3T����pS5�mfR��t�����i橿6nϿɱ��:"�&xD�C}`��un�3�i�_CS���0���
��Nտ�(������e6���������D���a�r�n�<�h�:XR���1�˶���Ai��c���f���a�
�B���(�BO��P�S���o�+��:4&���?�P�^�e���  �  ���\���|��� (�T�[������a��Mx���.�� ;����T�
s ���Z~��uk��ě¿���Ö+���`�dI������ S���f��ϵ���oP��]�濺:��Xb����I��#�:�����
̾^⼾0&��p�þ��پ1����j��~7� f�G*��`ȿA	�Z99���m��ɍ�����-�������jx� C�C�܅ؿm ��Z��Whҿo)�[=���r����c��Ü�aΏ�7s���>����;�ο^h��sk�=;��������"Uܾ�bžyٺ�J伾'w˾�g�k�s:"��|G�Sq|��a��T�߿��9kK�5�~�����m��]����.���h�<�2��"��ɿЯ�鹿%n���VjP�Zi��Eu��F<��袚�+��W�c��/����r������`� 6����A��S㾫�оs#ʾ�>о��q� ���Ͳ4��<^�����⹿i��F�*��^�s��H���|ן�7���������W�ro#����ԍ��<��K�ȿ���X�.�$d�K��槛�(	���!��.r����S�`� ��84���p���;X�dD2�����#�K��N
ݾ��ھZ$�����:�u|'�J�H��4w�ﺝ���п���#t=���q�b�����紟��&��o|��(G�!�2��5��-���|ڿ�4�u$A���v�n��b����ў��ߑ��:w���B�-�#]׿-ء�S|��K�G�)����T��j��M�ھ�Xܾ�9�W4�5��~v0��aU���]��`}濏I��N��'���ƕ�V���=���ō��,k���5�k%�E�ϿCƵ�ڿ�V�:��GS�a΃��ϗ��������o_���Xf�h2��8��ÿ�甿uZk�Cf@�ƥ!��/�Z������\�ܾ�L�P���U	�����<�:f��  �  Zъ���ſ�A�{�J�u��v��0k��������0��W����eD���/�ٿ�Rǿ�o��m�]�R�-T��ꃪ��g������7���>��������<��/��¶�p���?��>���i�ƾ�箾T������t躾�Uھ�.��x)�]9a�F>���S��!�u�a�rÒ����!���9���������O�p�,y0�%� �´ο�̿S���*��i�|x��H�����q���8���=I����h�;7(��P�=����0h���-����G�ݾ����w��;�����㮾�Xƾly�����;�\�|�#(��[���6�ey�<ǝ�$�������Y�����	����Q[��^�T�.�ʿz$ؿ��
�t�>���������ƺ�4���2 ��}��
.���:T�� �|�ѿ8��ObY�=�&������B	ž�Q���4��0K��_�ľWH�kN�L%�<zU�dR���B˿?�¶M��ӈ��u���Ⱦ�Ko��(U����80���jG������߿�cͿ�~꿟w��U����������͌��]��7p��媁�t@@����޺���|���VM���!�fk�@~徕2ξaG¾���9*ɾy`ܾT ���1���:��Ur��ˤ�����0&���e�;ݔ���������
������� ����t�܆4����?�ֿ# Կ)� �).��"m�J�������%������[���1]���m��h,�W��c��~y���>���2�����ݾ+�ɾ����0���Rr;j+�zF�k��8�I����ݷ�� ���9��n|��n��ْ��i�������u���u7���S^�oY"�yF���п޿���D�A�%��L��F%�����RN���g���z��k�V�ݿ��&׿TR���c��@1�w;�����|ؾ`OȾͷ¾ RǾik־�[�̠��;-�5v]��  �  �K��j�տnp��e��I��֝�����h���'�����@ʕ��l^����@B�mڿB���^B+���n����*��� ��������9M��֘��U�oJ���ÿ�O��h�<�j���hܾG��oa���ғ��ӑ�r������.�ɾ�����$�3�c�E������Yv5�K���H��J���32��Pk�������a�����DG��5�&�H�߿��
���?��_��A��/����g���S������}X���J��n�<�����d��I�k���)�+c ���̾�Ѭ�3s��c����g��-����쵾��ھ�
�O�8�y��q������y�M�����9��[��������P�����Yp��F�x�+3��h��2޿���ܸ���W�h%�����F����_��f���Q��*���I/p�Ed(��W㿚s����Y��l!�uG���о���׊��O������A���ϾRt��U&��U�͕�n.ۿ5"�2sh�?�������z���������i��!K��3xa�"��Z���|��i��E.�s r������������0��0������O����X�����ʿ&[���EK�.��:����ԾE���8����?������̾97�����5���t�R��������9� ��Kb��`����D���z��?���l��Bˊ�.RK��@��+뿚迣����C�0f���H������'s���a������@l���`��bA����γ���|�gy:�����;����w��]��������Ӿ����x���F��D��ۨÿL�Q��D�������j���#�����2������[�{��6��^��&�M�󿠸���Z�ם���_��������8���]�����)�r��+���迕���Hd��+��D����ˍȾ����4x�������ƾ��ྛ��XG'�[	]��  �  ����G�ۿ��%��o�G:��b;��@������ܥ��S/���Z����g��>%��u���_ῐ���(2��Dy�:z��������������Y^���������-^�w���#ɿ-���=�B�
�?�׾�A������d=��CL��!g��e¥�;�ľ����� $�Քe����)����<�����Ӯ�[����,��En�������������	�O�/��t�꿟3�n��|�G��!���Ȳ������\��[�������P*��a�D�&H��Q��7*n��
)����CȾ�ߧ����v9�������ܚ�Q�I־���~�8�7������~���lV�-������'?��K����#��^������ ����k:���4志���� �c�`��R��7��Gt��߾������/���}�z�
�.��;�Z>����Z�F, �[���b˾�1���䡾�r������8��%�ʾ����\��K�U�C��v�ῄc(��or�T���~���?��.8�����(���ݝ���j��N(�����vn�����)5��I|�����O���z���J������H��ԙ�\�a��*��пJ8���WK��z�4p���Ͼ>������#����M��xǾ�6��f��5�P�v��������A�g����_���V?���}��&����"��:�����S����Ę��F�S��j�K�E(��iд�^���>h��-i������'���@���H��{�9�����~���9���y��Ⱦ^ ����V����C��w�ξq�����F�V݉��vȿ�-�ҸY�u�����������+<��%���Pf��@���5��j^=���e(�¬����#�#�c�����q��mv���������#��x��;;}���1��|�+{��jOe��t*����޾�þ�ാ�򯾪��������۾L?�=�%�ȸ]��  �  �K��j�տnp��e��I��֝�����h���'�����@ʕ��l^����@B�mڿB���^B+���n����*��� ��������9M��֘��U�oJ���ÿ�O��h�<�j���hܾG��oa���ғ��ӑ�r������.�ɾ�����$�3�c�E������Yv5�K���H��J���32��Pk�������a�����DG��5�'�I�߿��
���?��_��A��0����g���S������~X���J��p�<�����d��L�k���)�%c ���̾�Ѭ��r�����5g������쵾��ھF�
���8��x������P��4�M�t�����7���υ��jP�����Hp��-�x�+3��h��2޿�������W�w%�����`����_������w��O����/p��d(�:X�
t����Y��m!�~H���о'�����T���Ҡ�����A�ϾOs���%�1U��̕��-ۿ�4"��rh���������z����������h��K��xa�"��Z���|��i��E.�� r����+�������0��V������O����X�\��&�ʿ�[���FK��.��;����Ծ
���ӧ��g@�����̾g7�&����5���t�S��������9� ��Kb��`����D���z��?���l��Bˊ�.RK��@��+뿚迣����C�0f���H������'s���a������@l���`��bA����γ���|�gy:�����;����w��]��������Ӿ����x���F��D��ۨÿL�Q��D�������j���#�����2������[�{��6��^��&�M�󿠸���Z�ם���_��������8���]�����)�r��+���迕���Hd��+��D����ˍȾ����4x�������ƾ��ྛ��XG'�[	]��  �  Zъ���ſ�A�{�J�u��v��0k��������0��W����eD���/�ٿ�Rǿ�o��m�]�R�-T��ꃪ��g������7���>��������<��/��¶�p���?��>���i�ƾ�箾T������t躾�Uھ�.��x)�]9a�F>���S��!�u�a�rÒ����!���9���������P�p�-y0�&� �ôο�̿U���*��i�}x��I�����r���:���?I����h�?7(��P�C����0h���-�����ݾB��w���젾���a⮾RWƾ{w���0�;�ȟ|�A'��(Z��c�6��y��Ɲ����r���~Y��}��诏��Q[�n^��S�&�ʿ�$ؿ�
���>�.���!����ƺ�n���t �����P.��C;T�"!�m�ѿ���cY�{�&�����F
ž{R���4���J��m�ľ�F�qM�%��xU��Q���A˿��6�M��ӈ�ku���Ⱦ�o���T��Ȥ��0��UjG������߿�cͿ��w�K�U����$��$�����J]���p��/���A@�D��ػ���}��xXM�6�!��l���4ξ�H¾Ǩ���*ɾ�`ܾ� ���1���:��Ur��ˤ�����0&���e�;ݔ���������
������� ����t�܆4����?�ֿ# Կ)� �).��"m�J�������%������[���1]���m��h,�W��c��~y���>���2�����ݾ+�ɾ����0���Rr;j+�zF�k��8�I����ݷ�� ���9��n|��n��ْ��i�������u���u7���S^�oY"�yF���п޿���D�A�%��L��F%�����RN���g���z��k�V�ݿ��&׿TR���c��@1�w;�����|ؾ`OȾͷ¾ RǾik־�[�̠��;-�5v]��  �  ���\���|��� (�T�[������a��Mx���.�� ;����T�
s ���Z~��uk��ě¿���Ö+���`�dI������ S���f��ϵ���oP��]�濺:��Xb����I��#�:�����
̾^⼾0&��p�þ��پ1����j��~7� f�H*��`ȿA	�Z99���m��ɍ�����-�������jx� C�C�݅ؿn ��[��Yhҿq)�]=���r����e��Ü�cΏ�<s���>����F�οgh��sk�>;����`����Tܾ�až�غ��⼾pu˾ce�
��8"��zG�o|�t`����߿U��}jK�z�~�����m������.��+h���2�e"���ɿsЯ�<鹿on�!���jP��i���u���<��A�������c���/�F��fs��M���0�`��6�[��-B��T�j�о�#ʾ->о���j� �����4��:^����Sṿ� ����*�F�^���꼙�(ן��K���`�W�.o#���򿪍��?��{�ȿř���.�t$d����2����	�� "���r��T�S�(� ���5���q��>X�FF2�5���$�\���ݾ��ھE%徯����:��|'�c�H��4w�󺝿��п���"t=���q�a�����洟��&��n|��(G�!�2��5��-���|ڿ�4�u$A���v�n��b����ў��ߑ��:w���B�-�#]׿-ء�S|��K�G�)����T��j��M�ھ�Xܾ�9�W4�5��~v0��aU���]��`}濏I��N��'���ƕ�V���=���ō��,k���5�k%�E�ϿCƵ�ڿ�V�:��GS�a΃��ϗ��������o_���Xf�h2��8��ÿ�甿uZk�Cf@�ƥ!��/�Z������\�ܾ�L�P���U	�����<�:f��  �  �S��EE���Uֿ����s)���J��b�K�j��_�wLD�M������̐��[����Ǝ�G;��b�ƿ����$(��K���c�O�j���^���C�d�!��� ��%̿�.��"T��INh���E�&�'�e���F��z��m���0�H��L����7�^X���~�ᗿ�W���D�����@5�oIT���g�sli�hX���8�I!�ۄ�i���ݒ��q���H����ٿ���4��dU�%Nh���h�$�V��8��V�&��W������U]���][��:�M���j���0a�H��a����k���&��D�ޞf�"���,��B�ȿ���~���A�V"]� k�q�f�h
P��z-�����8ϿK$��Q������\��#U�{���0B��1_�Jl�2\f���O��@/���e�߿S*��V&���g|���W�ݡ8����\�
�������i�����	�m��H~7�MjV���z��ғ�Fʱ� �ۿ9X
��+,��EM�`e�|qm�{�b��"G��|"�	���S��������ݔ�;`����̿���`+�@�N�Kg�4 n�4!b�dWG��`%��W��ӿ�*��f��\�v��IT��7�M"���������?���-�$I�C�i�h��v��:���0��q	�mu9��vX�<�k�Y�m��\���<�Q2�Ϡ�����񚿥��� ]��G��f��3�8�zxY��fl�V�l��[��<�:��G]����ſ���Ӊ��Dl��XK�sj/�]�6v	�2�����3T����pS5�mfR��t�����i橿6nϿɱ��:"�&xD�C}`��un�3�i�_CS���0���
��Nտ�(������e6���������D���a�r�n�<�h�:XR���1�˶���Ai��c���f���a�
�B���(�BO��P�S���o�+��:4&���?�P�^�e���  �  ���������f̿oV�<i�s��f �m�#��G��	���ӊ��{�����q�ce�g=y�����xm�������0���#�av�P��<���bO�iȿh���'���ĭ�� )���[^��;��!�Ml�߂�8��2�.�`vN�>�s�u���<h��.�������'�Կ�.�&n	�D>�<�"��N"��d����uqӿd=��¦���j�_�h�ヿ�ܢ��	ο�9��fZ�sf!�@#�����!��Q��]"׿���诿𿟿I����v�m�Q��P1��%����H��YM��_9�>�[�$���擿�,���f��Gdǿ��޿	���������$��R �� ������ſ����AZ���k�Aut��4���첿���*[��z��
%��-#�˻�zC�����ҿ�о�$e��8��
���;r��?N���0��J��9��R���.��L�w�o��.��Ҁ��*��K���g�ѿ/�뿶!����0#��?&�
�������Md���x���}�|8q�΂�>�����Ŀ�����<�˚!��b'���!��A�KG��@�+�ο𪼿Ч��Z雿䕉�ϡm��K��31�%�!��3��)�D�?���_�r`��1]��Z���;���ȿ�Vݿ/���]��Cl�)'��n&�O�����ۿ�Y��������z���x���������$ֿ@-��n�\%�9^'�����K�Ѱ���߿�ɿ�`��?<��Ŗ�Bヿmb�B��*�:'�E� �4/��H���j�3;���隿^��� ���οu����."��y!�m(��#��`�����?̿���Sf��� w��������������W��"�/�'���%��L�t�	���Nؿ�Ŀ�����6���1���P|��"X�g:���&�~���f%��7�G�T�Whx��H��X����  �  ��⿢��`�u6��W῕�����pK� �ӿ�껿O��c��X��e<��H4��A�ȅa�����ǥ�:¿�ؿVZ�����係O�⿫�忐 �.�࿜�п�������%~��ES��=:���5���E��9i�፿����r�ƿ#ۿM�� 翊���a���
R���Z!߿�-ͿL���ϕ�
v���M��8�O�6�LhJ���p�5��Ѱ��*fʿ,cݿ�#��H��⿄�࿇�⿌@�	���Hܿ�ȿ��������bm��3H��5��8�
�O��Jy��헿�g��	oϿ�	�%S���b�~�⿠c�!��Y�濘�ۿ��ƿ.��S��Yk�B�H�m:��,@��Z�e=���!��tR���տ
��9��?��Gz�W��U��B��ބ�d�ڿxUĿg��΃��*�g�ujH�%=��F��d��9������ԉ¿�ڿ�'��>쿜�� �������$6�غ�Aٿr���wʤ��È�td�;mH���@�{�M�1n��r���b��i�ȿ��޿�M뿥��`��E��	��������׿
%��F�������c���J��F�0�V��oz�慖������2Ͽp��SD���F쿙��X9뿵�ￄb�#cտc9��g�&$��*^��BH�GG���Z��i��ʚ��Mҷ�a�ҿŕ�#a��[�EH�vK�V�'�����=ѿ�6������D~���X��F�|�H�O�_�ul���x�������~ֿ?���￞@��A�鿡쿡E� ��v�bͿљ������pw��U�vF��K��f�:∿æ��j���vgڿ� 꿊�ￚ	���g���$�￭��9�߿.rɿ���o��G<q���Q� OF�U�O� m�����,奔�ƿ޿�  �  ѕ#�y�� ;�s�e���:˿1!���觿�D��"����c�~@�m9$�/���r�
����)�'H�}�l��Z���P��f���PD����п��|u�~����!�O #�����GYۿ�ۭ�����n�̹f�c2���Ŝ�uTƿ�f��<W� ���#����:"�/9����ۿH�Ŀ�!��C��ؑ�_7~��uX�N�6������U�{���w3� 1T��y����6����T¿�ؿ��� ��&��O#��� ��&��*����ʿ�X��k5��Sg�"@k�a��y���b|ֿ0l�-��R<#��I#�o3��6	����[�Կ����<���
���b���u��qP�V�1�{R��!�L�߻'�HIC�$nf�]_���kݩ�>��ܲ̿�b�^|�tg�� �K�%�M_�����J�"��!�����e�m�N�|��ݕ�m������w��v��S&���"�Y���2��-�q�п���X��W������?o��L��0����#���!�U�6�mU���y�����1��5����@ÿ��׿����	��A�`S%���&�B���\	�l5�Z���}P����~���w�sՈ��s���Ͽ���ȯ�jh$��0(�!��f��Y��a�U6Ϳup���I�����+G��m�h�,$G���-�\E ��~�d�+���C�id����Ǘ�m&���D����ʿ������$=�`c��'�E%�m�F�� �ӿݨ�ܬ���x��{��!��,~���(޿6�P[��&�-�&����<�����Üۿ��ƿ0�%�����O����]� >�k}(����"�513��N�eq�����56��p��9����ѿ]��f�-��i#��O(���!�Y/��E��.�Ŀ؝�ק����v��܂��^��e��<���N� ��  �  G�j�O�a�Q�H�H�'�|��\�ӿ�l������	n��CJ���+�������q��$��Ύ� G����2�pR�]`w��������B'߿H+�gj/��O�re��bj�7Z\���>�8d�F �X������c鏿����oп����.���P�|f��j�'[�4�>�H?�T���#�Ŀ��������bb�ˉ@���#��P�����`��@��z���	�� �%�<���]��ׂ��i���ɿ�+�R7�Z�:��BX���h���g���S�s2�ϗ���տ�Ϧ��j��R��K������HW��$;�9Z��fj���g�M�S�[4�&�����=���ԗ�S����Y�U�9�d�	
����	)���Y�������/�6�M��q�����y��)9ҿ�R�N�%��ZG��a���l�m�d�i�K�G(���\ȿ�������Y��s�¿�:��D#$�-�H�zqc�nm�Njd�K�K�B*���|ٿد��}��%y��cU��47��#�-@�����{���M���O%�-�?��_�}������������ 濕��Z�2�hS�@�h���m�|`���B��e�E�μ����&���~M����ؿZ+�E�2�M%U�U�j�`n��r_��B��| �/5 �H@Ϳ�c��E܍���r�Q�P��4�+��V�������2%
�����0��M�.@n����j���ȿ�����h�0�>�&�\�m>m�T�k���W���6����v|޿j^���똿�����ͷ��	�pA���>��]���m�sk�9�V� i7�e�qj�V������n|����f���F��+��y��/�#�r��L���!��u:�]X�u�{�?��	���D_׿1���.(�u�I��%d�6o��eg��IN�l|*��'���̿b���ݸ������]ǿaY��P&���J��|e��  �  
s��2���=u���Y�TD%��;�u������0�P��q(�pE�
��Suξ�E��z��S/��n=Ծڰ��mG���0�q�\�/8�������r�0�1�d��a���`��E���Ҕ��S��L�u���a�v�f譿%*ʿ�7�W4���i��ٌ������˝�Rђ�ֈ{���G������ڿ�d���lv��B�$���I�Lk�E�Ⱦ����򺾑�ƾ��޾̕������=�z+o�	����ҿ(d���A���u������ s������o�P�9�d�	�p�ο쵮��Ͳ�iUۿhx��F�1i{��=���-���ԛ�����~k��7�O��WoƿQd���%f�!�8�ku�� ����t̾s�þS�Ǿ)-ؾ�����P��+�sS�2���}�����!�� U�,������W��I��/��f�_���*�2+����Ŀ�������V��o}%�`IZ������5��\Ο�����Ն���[���'�#����ᶿ�.��]�[�֏3���������-LվfѾRIپ���r����<>�PLj�Z*��Yſ���
4��`h�c��]"���������J���P������>���������ҿ|�	�b�8�2_n�R���ޝ�����R�������K�������U���9x��"FS��.�`��ip��N��ܾ�F۾`��Q����Y7+��N�f���G��/�ڿ�����E�z�����.��D��� 	����s��1>�����׿�R���Z����ę�J�z?�,�����-���������n��l:�}�
��#Ϳ_��Kns���E�oe%����u����g�Hs۾l�޾������X3�)r6�A�]� ӊ��������W_$��W�$2��,i������ ���VJ��Jnb��?-�� ��qɿcP��qſ�����'���\�Oԇ��>���  �  <	��ۀ�����`����UG��c�����c����G�l��?�� �ʾ�����h��Ą��7Ӥ��µ���Ҿ_���]�!��U��D����ҿ�j��1V��-�� ����������{���E���|�$I:������ӿE-ɿ�?�@!���]�a������}���9.���`��«��Ջt��2�����UQ����u�Υ6�����徙^¾�P���f�� Ġ�#_�������྇�	���0���l�=Y��O�ˌ+��l�z	���г�dH������k���$����	e���&�`���aOʿg�ϿZ���3��xt������y���e��� ���I���^��{�\8ݿiƚ�c�`��`*��)���߾���`�����f��:㺾�6Ծ������i�H�;5���P���B�t���8A������3������@���yx��Z6Q������忳~˿Ԧ࿽���/J��ǆ�0������a��޽������xJ��2Aǿjԍ�;�R�ƽ#�����'DȾp��������tϾ�$��C��Y/�(_c�f6��~�ٿ��L�Y�:���y���������~ٺ�kF���$����>�_�,�ܿҿ� ����%�eKb�4���$������UW��r���Ν��x���6��� � �������G��1��8���⾱�̾���{����ʾX߾D� �b9�pA��}��������t�/�-�p��%��6��tj��t������¯���^i��+�n_���ӿMؿ���=�7���x�8ݝ�Ἰ�U���T��N���I�����a�b�"���㿅u����m�<�7�_��[����ھP�Ⱦ�r���Wľ�Ѿ�n꾣��A&��#S��c��]ÿ�@���D���g����޼��4������(6��o���l�S��6�#��*п�S�c��}L��������*���  �  ޵�����Qͼ�����ra�k
��ѿjq���F��{��X�e������Ɠ��C�������å�¾� �p���V����s��M=*���r��ݠ�h��������\������5O��xM��٬R�i���鿜�ܿ�&��Y5���{�����<���������������������H����~���L{���3���x.վ�䱾��������k��~-�� ���.�Ͼ��-�;q��U��k����@��|��\��w'��i������8����������;�����ݿ8�xZ���J����k��*B�����{���ˍ��^��� N|��l2�񿶘���b�Ԋ%�����Ͼ�ñ��m��$X��L���JP��ݒþ�S뾓���F�Xv���˿�K�%�Z�o������:������@.��)m��:g��5�l�!D*�����p�޿f����'$���d��!�����'q����ok���)���u��C)d����oֿ�Ⓙw�Q���1����Ѿ^���Cϫ��٨��#���y��fXܾI`��*�Yd�"�����-��Gv�@�������
����4��e���9X��m��UW��=����������9�!!���3���k������Z����4��줳��$��`+M��,��̿��煿��C�:�����ZҾ8b��dY������\�����ξS�����a=�U������������D����kx���F��y��������^���5��[;��xV@�TW�����ױ�XO�P����h��l%����������@��Y5������5�q���\G����o��2�Q^�I�辘�ʾ�й�%-��6̵��	¾$�پ� �A��(xQ�ۤ����пD��k�]������a��5*�������n��P���z���Do���,��7�X:��8��Y�&��g��F����������  �  �3���P��s���Ȍ�4�P�����7¿>���-v8�r:���оl_���C���+�������2������:ѱ��ܾ���UG��f��@�Կ����`����9�����������Z"��<ԧ�Ô��u)C��c�rmڿYϿB���}I(�(i�ñ��X~���X��Z�������m������-�9����^�����i��k&�����<�þ�ꢾ����T���4��R��;ڟ�����P���J ��#`�������zt2�U�x�r���� ���n���k���A��ep��Y�p��V.�K����[п�ֿ�m�b�;�����8<��3���1�����������O��4�i��E%�l�߿q����R��u�d7�Ҕ���v��5�������������*���)پg
��9����8����Z��J�����ox���H�����+���&������5t[�YP�u��cKѿ:������S�hÍ�}�������������H���$���GS�	G�a�ǿB���rC�9Y��g羙c���ª��0������HS��_P���̾�i��w0��U�S���ۿM"!��d�\����H��0���
�������ש�r���}|G����,K� ؿ����ʳ,��qm�A���������������a����Â�b,>��;����oDz���6�I��\7�cWþ����즾�`��\���3���"߾*��+�0�H�p��W��	��k�6��}�˪��?����������g��L���|u�Ǯ2�7:��ٿ�޿����,@�Α��{5������`��2b��K�������L�l�0�(�Ԩ�
���`��&�����׾�Z���鬾pᦾ�D���p���Lʾ������G�C��/���¿���{QM�!��� í�B���c���k��S_������]�9� ��K��տʧ�=��CV������������  �  �@������SY��m���bH�sb����ޟ��8�[��.վ��8ɗ��x���4�������3��Nu�����i���XF�ی��aο����CW�����#���#������sѺ�����~��U;�S��ӿ��ȿ)|��!��j_�^>��ۦ��ћ���m���~��R��5_v�z�2���������Hg���&�i��T5Ⱦq����(���܊�aQ��w��\{���Gþ�_���� �^�B���U���x+�kWn�m������8���e����I��Qѕ�+�f�t�'�?���ʿ�qϿ��y4��Lv��J��K�����������E�������8�_��	�%Fٿ󔔿o�Q�j�1�n4þ����꘾GJ��\J���8���ø���ݾK����8�#J���۸�Z����B��ԃ��
������0'������g������ҋR�8l�_��,˿���7(��hK�\ه�?������ߖ��r������}����J�d��o¿���C�m����뾹ƾ�H���|���Ġ�a����ൾ�о���NN��T�,Ǔ��Uտ{A�_�Z�aD��fl�����l�������뷢�r��z�?�����nܿJ�ѿV��M4&�-�c��m��~Ӳ��������������r����z���6����[	����w��/7��S�]����Ǿჴ��,�������Ʋ���ľ����p
�=/1��qn� ʧ��=󿼢/���r�Ĺ��:��@�������<o������ k�f�+�����ҿoؿ���W�8�kez�7A�������|��В��Ǫ���c��c�~`"���߿�<���^��'�=��"�ܾ����~G��d�������︾.�ξ�A�K�uC�Qx�����
��+E����>V��&���o������Cά�ǩ���T�������Ͽ�P���Z�M�$������ ���  �  ����J��d���|�l�=1�Ͻ������ƫz�F9��]��.�/���a����gw���S��m	��]ƾm�e���E�%�������Z��C>�*Az�k6���$���s��B�����	�_�F�%���!���C����׿���
E��}���	�����������4����X�6���߿�*����b���)����׾XӶ�Mc���A��𩗾����������Ҿ�� �6s$�X�Z�� ����ֿ*���Q�һ��Oe��F"���m���R�������GK����$ݿ����$H��R�J ���X�|)�����xM�������)���р��E���/ȿ.捿P����څ����Ҿ���yΦ�����ͣ����f+Ⱦ��f���:��cy��	��������,��h�wɐ��c��������]���G�u��0:�]�Hѿ�J���̿���54�D1o�����������y��o��I�o���3��� �qg��Iɂ�)D�}�=����վ�ཾ��*���m����ľ�5�5�KK$��yS�/��ſI����A��}�d��>���B��K̥�7��a�c�f7*�^���۔ɿ{����w࿵|�vmI������6������U��Kӣ����&]��I#�\E迁u��]s��3:�U���-��k?׾�¾̑��-���������Ӿ6�:>�A�4���j��<���߿,��/V�׈�����9C�����x�����0�O��I�#��pS��'�ſ����F$���\�,���������	k���՜��{��:�H����%�ο����H]�^,�v��$(�<�Ͼ�*��pa������gǾ{b޾>��W��2E������/��M���c}/���j��������ܰ��+��>��-x�ܐ<���
�W�տ�����/ѿ�;��e6��oq�75��/����  �  �c��f��w�l�}�@�E��ݗڿ�����v���A�&��c!�Qݾ�����������Ʈ���5Ǿ�"�+��jm$��SL�_ۂ�W&���H꿗��tFK�cu�l҈�N<��vփ��wc��N5�5����̿�p���{��𷿯��A� ���O�>�y����+׋��%���*_���1�c"��ƿ:蓿{�c�E5�,��Ȑ���gԾ�޼�������������оI����0o0��-]�j#��K'��Њ�r,��Z��Q��,��9����%}�w`T��s%�\���7��^(��������ƿ�!��/0���^�ky���1���'���4z��,Q�TV#����E������(mU�6),����'򾗍Ӿ�k������\}����˾�^�d�ω ��YD�fw�l����%׿`����=��$j�����L���Ȉ�2s�wG�ܦ�8��/ʳ��d��1c���ݿY�B�^o��݇�����Ň��no�ΝC��g����p��"�����L�_(��o�J��[پ�ɾ�ƾ�;=�ྣH��� ��1��Z��ǉ�q��u;�� �#�N��x�\����������\g�i[9����ViտV��r4��1���H��t%��S���}��������KJ���lc���5��U
��_οQ3��1<t�"{E�^N$��
�����8ݾ0�оA>о�۾�:�|	�V� �Ѿ@��m�_���nǿ���(�0�O^��o���L���������T�X�f�)�@���קĿŷ��6���,Ͽ�9��&4�*�b��J�����d؋���}��}T�Z�&�Ѿ��[���;����b��@9������m�<�ؾǀоH�Ӿ�������F��5+���N�>���᥿�Kܿ�{�E@���l��V��\���"����u��sI����K鿺}�����k��}p⿄J�PED��7q�Q���  �  �:P�%cH�,�2����/�3}��?������ \�:�;����#���x�	پ��Ҿ�ܾ�q������%�\�B�ǥd��k��Y���a�ʿi��������8���K�E�O�!�C���)�G	���ӿ`f��w�������3˕�q����^��Ҏ�0p9���L�~�O��B���)�\
�*࿳���j��;�v�A�Q�h�2��w�F��L�Q�־'�վ&���� �����K/���M���q�!я����J2ڿ����g&�U4@���N��kM���;�����������{������ ���h=���Ϳ���F�&��A��P���M��2<�q� �_��saѿ���D싿��l��J�+-�N��xT�'�0޾B+�̑�����~�#�[D?�~}_��G������@����RY��1��H�:&R�t>K�wA5��ZW뿄��e���އ�|�����V%�e���2��J�`�R�%K��5����ӧ���ſŭ���t��g���F��#+�A���8�}�y����~����/3�]6P�!^r��W������}ѿ�j�� ��!<��4O�A�S��CG��y-�l��ܿ%ʬ��	���:��`w��|6ſ���#���=���P��	T�z	G��.�EE�a�迧����h��n����b�=C�=�(��B����������i�j�i�%�_�?�}�]�	��j���f��J��S��K�*��oD� S���Q��5@�5-#�>�&ʿ���������mv����տ��	��M*��_E��S�`!Q�q�?�y&$��P�v
ؿ����ŕ��'�y��2W�h�9�~?!�f���� ����W���k2���B�.�\�I�2 j�+x��0ߡ���ĿF8������S4�%K���T���M�g�7�o���1�պ�[ʘ������_�����Қ鿡����4��&L��  �  ���8���뿄�Ͽ�����|���̙�T���X�t�L>R��V2�������-�3|����,;9��Z��f|�1i��E���<���F��D�տq��tN�������������ƿ�N���t��*\��U��cl�3X������,�ݿ����v��l����-}��Fȿ{𳿥��[m���ⅿ"j�[	H���)�����������§&�:,D�Q�e��܃�����B����Uſ��޿@��{����B�����\�������s��y�o�55V�׸Y��Az�����*���Z��������	����U�ڿ�S¿.ů����z������7#b��6A�a%��&���	��o�����{5�8/U�U�w�����=꛿.����E����п44�����\;�l��V���M�׿r������Q�l���\���i��̉������Կ$���i���%�����C�Iտ&���Gꭿ?���:��g����]�]�=���$�D��{h������*��6F�@Vg���:C��P1���1���:ſ��ܿ�t����
��:��F�	y�7��*�Ϳ�Z������a�l���f���}�N���[��^E�q�X���ô��$������пUI���Q��{���H��eVz��JX���9��=#�������1!���6�P_T� v����2���]T��|�+�ͿD��@��@�]5����	���=꿬;���Vc����f�/0j�k4�������ɿ�l��`��W��u�����+���L�6�ȿes��sU��2���𕈿	 o�=�M���1��N�k��� �(�K�@�L&`�6��ݑ�����ï��k��pֿ�i�D�M��D���2�ƅ�l�ܿ芳�\X��\Kv�f�K!s��L��?a���Kؿ#� ���  �  ^Ϳ6ѿ5gϿ��̿DͿL�ϿEѿڳ̿ꬿ�͚��0-����p��@H��/�q�'��63��4P�F{�<�����,�ÿR�ο1_ѿ�JϿ4Ϳ��Ϳbkп�4ѿǂ˿H���fᦿ2����i�W�C�|%-���(��7��#W��������@��;Mƿs�ϿV{ѿ�Ͽ2Ϳ�Qοѿ��п��ɿ�蹿0٢�����b���>�=<+��'*���;��]�����ݟ�^n���LȿeSп{�п`8ο�̿�Hο��п�Ͽ�Jǿ4쵿����U��t�Z�3�9��Y)��+�ɏ@���e���������	����˿�ҿ�Yҿ��Ͽ��ο��пDӿѿǿ[��� !��w����DY�C�:�l�-���2��J�v�q�u����^��K���nϿQ�Կ��ӿ ѿ�п	�ҿ��ԿL�ѿ�Vƿ~��E���DT���V�.�:�dx0�	9�T{S�]�|���������ſمҿ�ֿ4�Կ�oҿ��ҿ�տt|ֿr&ҿ�.ſ�2��-ߖ��'|��T��;���3�Ӡ?���\���䮝������dʿ�տhTؿ�@ֿVԿ �Կ
V׿x,ؿf�ҿ�?Ŀ�X��M䔿l|y�P�S�l�=���9�O�H��Ch������U�������ο[qؿ�ڿ��׿��տ��ֿ�\ٿgIٿ ҿ�¿n��O(����r�j�N��b;�:L:�\�K�#�m�0������є���|п{�ؿ�+ٿ{�ֿ�տ!�ֿ�Eٿ�Uؿ�Ͽk������ˌ�E�k��TJ���9�{�;��rP�@u�瀒��M���ÿS�ҿ`<ٿ��ؿMMֿ�[տ]׿��ٿ,�׿B�Ϳ4
�������숿c�e���F��u9�'�>��"V�\}����ð��ƿ��Կ��ٿ{�ؿqIֿ��տ�2ؿ&+ڿ	׿l�˿����i����A��*`� &D�v�9�(B��g\�O���ԛ��-����ɿ�  �  z��H@��׎��8ѿ!B�<����}���
�����k�̿%��]����r_��T���e������¬��Kֿ�)��Y��u� �����	̿\����P�����<m���{o�RM��3.�������3��p�V�"��?��b`��F���;�����0��=¿��ڿX����k	�H��.�����鿮$��膘���w��"Y��xW���r�2����j���i���W0����k�
����VYݿ4Ŀ����M���k��ݤ���Sc���A�Ĳ$�
����o$���� ,��"K���m�<܇�����9��a��1˿����j�ɶ�N�z[�M��,ݿ\���qˏ�|�n�@Z�=jb����Z��TH˿;����,�����$��[��l����׿P����㮿�
��4����q�_���?�"�$�RU����ȁ��e#���=�7 ^��W���ߐ�y����Ʈ������ֿ¶򿗲��5�]�����g��svҿ�񩿹����wk��A`�mWr��>���&��g�ܿ�j�������W������}�ҿT���/I��Ȟ�-����H~���\���=�&��,�)��D��~3��P�O�q�x߉��ә�p���z���)�ʿ�"㿏 ����R����i�
��F�Dǿ����V����Hi���g�䆁��Ü�6�¿@������G�!����sq�J��[i̿5�������⚿��6t�ՖR��a5�iE ����a%��,$�+d;�~�Y��|�hڎ�S��������ѿ�7�_��������I����_����{���e�.n�����Ǩ���п,\����	9������
�͕���/ݿ!�ſ�"��$G��,f��%���j��pI�1�.�����>����C,�TRF��f�q���┿�  �  �#��,ߝ��¿U7���t��A4��FI��>P�t�F��y.��v�%ݿ�����&��	�������X���꿞����4��6J�_>P���E�$m.�i��4��g���S����]}�f�V�zL7�`M�"��5��Aؾ��Ծ�������z�*�}H�Q�k�Vȋ��|����ҿ���þ!�*�<�F�M�^O�x@�!�$�f����ʿG|���3������Rƚ��Ŀd���]� ��w=��N�N�C?�E�$�m���g׿����x(��-�n��-K��4-���������⾨kվ��׾~�龎��9��-6���U���{�j	���8���}俼q�6-,��D��P�'�L�|�8��������i�������d댿���^�ٿ+^�2�,�"EF��Q���L��
9�?���J��ʐ˿kO��m�����i�[uH�w&,�l�/����R��E-��|�7��|J+� �G�W�h�����ce��TȿE����.�G�6��K�M�R��SI��N1��Z�Y����,�� ���:���������%��-8���M��S��?I�t�1�wd�Ѓ�X���՚��{���nZe�BF��a+�[���n����������6�����"��<�:�Y�~�|��V��C����ڿ���%���@���Q��;S��7D���(����ҿ�����F�� ���آ�t�̿��3�$�s�A��3R�3�R��;C�{�(����߿�`������&��S	\��>��$������`���gw��kl�1��)�svD���c�%��������޽���j��1�/��G�T�e�O��<�o���&���%¿n���$����Ӓ�C��{߿�.�3�/��H�-uT��PO��;��S����v�пK���"鎿�Ht�úR�6B6�-W����t����)��XG��/O
��6��3�U�O���p��  �  u�y�����<I޿~�>qC���n�o���h�����OSj��=��V���տ�U���&��!\�����D���G�Bs��h���K��Pl��If�:X9�����п�͚���l�q;���t,���پ-���4���_1��n7����̾r쾷q�ι*�x�T����*������%%���R��i{��?��b���[n��:\�y�-�	�n\Ŀ%��0c��g�������F(��%W�g7�
�����u�~�V�W��)����ݻ��ˌ�%�Y��-������ξ�������౾-f���Oؾ�����w���9��ni�������ʿ�	�95��Mb��W��|t�����w�x���M��:����C���t��16���uҿ�/��S9��Rg�a��Q0���&�� u��|J�1������⭿�����Q�*���, ��g־�ž�5���ľ�־}�Q|��(���N�ii����������],F�`�q�=h���Ǎ�"Q���.m��?��N�I�ۿ^^��L6��Ks��3꿎#��J���v���u���%����i���<�cH��׿�š��{�A�I�}('�������߾�Ѿ��Ͼ�Uپi!��t�y�;��f�{��������4��mO)�v!W�����Q��C���fz��jM`���1���bq̿{7���t��L#ǿB���R,�E4[�����I������������[��.�G��XDĿ�6��Ϣj��>��[��d����!ھ��Ͼ�>ѾZ޾c=��2�B�%�UdG�w��M��x|ѿ�n�Dd8�Ӟe�����X��\����{�ZQ��H"�F��f���j���$��pYؿ��".<�gj�����M���Qr���w�mM��n���P ���ŉ�ql[��Y4��)�~����=ؾ��Ѿ�־���������2!1�/�V��  �  �~��_��g\ �Hh4�) p���� ��R���p����v��5yi�M�.������ſ_��)ϿՐ��?;���v�B��Ѩ��q�������o��Y�b�T(�>��P��{]n�=[1�R�	�� ޾����*¤���R
���x��x対�̾�>�����BP�������ʿ���;H����	��
��������n���y�U��p�������z7���࿪��Q�N��Q����������/ά��Q���/����N�>��vҿ#���uV���!����о�㱾�ʟ�Z痾�����󤾿����ݾS<���.��i�K������4�"�A]������ ���s���D����~���B�v��q.׿�����ĿPz��`2*�7Ed�	V�������m���S��
×���x�z�<�dw�킾�)����I��&�����"Ծ�g���ݫ�@'���꫾�h��X�Ӿ����Ϧ���F����v渿��F)7�h�r��s��_J��<������K��yll��1���̿�%��6տ���R>��z�����JN��L7���J���&��RUf���+��n��G��1s|�۪?��������پ��þt�`z���i��;AѾ���S��s�.�Ra���.ӿ3��<sL��+��(��� ���ͯ��������ҞY�G}!����A�Ŀ�H¿�
鿈�� �R��X��m��������ۮ��a���B����R��I���ڿ�i���Bg�)d2����񾂣Ҿ���_���gƸ��oþ�}ؾ����c��}<��v��J����_#&�!Y`�C���g���EA��z��G՛�R���E�̻��#ݿ<�����ʿ2j��3#-��(g�D�����������'���n���J{�G_?��
�d�ÿ�c���FT�zm&�_+�� 辒�;"۾������G�˾d�侳���"���N��  �  S#���
��W���K�������Ҡ���B��۽�����)���ؕE��b�^�ٿEǿ��e�7T��{��`"���k��X��2л�w������G2=����D���@�t��F/�O��ξt����Y��$������|���k㠾i���뾣{��?R����рܿR�!�2�b��:�����#)�����5V��It��3�r�sc1�t� �ۀοp�˿�r��p�*���j�ɗ�,���8��(��E����ԗ��wj�(����y��|Y�E���D�ΐ���ޢ�
ّ�����M��bǖ�K���t�;N����+��en���������6�.{�{������)���l��x��������\��
 ���1�ʿ�ؿ��
�S@�
���9$��j���b����8��Q��=|���4U�e�DͿx���5J�f���Y��ľ����!��-虾xI��<ƫ��Tľ��뾇���E�'���0�ƿJ�*�N�����U������ĥ���E��*���<��ڙH��j���߿yͿ��2�0!W�]������ ������,����+��@����@��_�����f{���=����l��ʾ�r��QX����`]��s&¾<߾�u��{*��Ic���������%�zg�iS��!���:��\.���a���}��p�v��o5�����ֿt�ӿ5� �6�.�x�n�%Й��Ķ��B��q5��V��������n��:,�6��y��ZCj�Č.����h�ᾮ�þ��h\��Z��	&���.ɾ���(��a�9��{��g������1:�Y~����F�������}��dC���l����_��#��v󿹗пN ޿ ��p�B��������
��'I�����9T��[Ɏ���W�i��ҿ�В�crT��<!��� �usؾ���V��pi��TM���M���dվ_���q:��M��  �  v?���|ƿ˰�d{T�@ю�ɜ��TG��5���Q��2��y�����M�������)'Ϳ�X���K,]�����ų������K��Щ�����s%E�3�����x��C/�����hʾ�ޑ�OU��F����&��'I��:͸�6,������S�4&��(|��'���l�����������0����|���S��!}�C�8��z��տ]3ҿ[4���1�-�t��}��uļ�������ռ�J���8�t���.�i^�wt���_[�'���I��H���z�����}���[���馾�Rɾ� �x�+��q��ٯ�����v>�b�������x�����9#������G���Gf�2c&����N�п"�޿���H�RD�� T��=��o�������hд�oΓ��W^���!nӿ������J����72龚￾T���͙�b���J����>�����������H�F�8���j̿8u�k>W�w1������Ϧ����������؃��s����P���}翢0ӿ\�"�#3`��5���X��U���{������U��� u��E�H����������=��H��&��Tžb	���ϥ�r�都�_ھ�Û)���d��������q;,��q�,���-������������]��������<�̈́	��ݿVDڿ=��5��y����-;����.�����
à���x�3����5٧��$l� �-�p����ܾ�澾����� �� ��E���ľk;�U<���9���~�\�������A�����FN����3���>����	���ɘ��Ai�HY)�������ֿ����2�J�2���k����h��%7���@���������`�(����ؿ96��pFU�w
 �do����Ӿ߃��~ɬ��1�������ĸ���о�\������~N��  �  S#���
��W���K�������Ҡ���B��۽�����)���ؕE��b�^�ٿEǿ��e�7T��{��`"���k��X��2л�w������G2=����D���@�t��F/�O��ξt����Y��$������|���k㠾i���뾣{��?R����рܿR�!�2�b��:�����#)�����5V��It��3�r�sc1�t� �ۀοp�˿�r��p�*���j�ɗ�-���8��(��F����ԗ��wj�	(����|��|Y�D���D𾱐��pޢ��ؑ�����M���Ɩ�b���R�;���$�+��dn�e��������6��{��z��f���)��ml��Z��������\��
 ����+�ʿؿ��
�o@����S$����������9��~��j|���4U�je��Ϳ����J� ��[���ľ����M"��3虾6I���ū��Sľ�������E�������ƿ���N����RU��v��������E���)���<����H��j���߿zͿ��G�Q!W�t������F������\����+��o���g�@�`�����{��˓=�������0ʾ�s���X������]���&¾q߾�u��{*��Ic���������%�zg�iS��!���:��\.���a���}��p�v��o5�����ֿt�ӿ5� �6�.�x�n�%Й��Ķ��B��q5��V��������n��:,�6��y��ZCj�Č.����h�ᾮ�þ��h\��Z��	&���.ɾ���(��a�9��{��g������1:�Y~����F�������}��dC���l����_��#��v󿹗пN ޿ ��p�B��������
��'I�����9T��[Ɏ���W�i��ҿ�В�crT��<!��� �usؾ���V��pi��TM���M���dվ_���q:��M��  �  �~��_��g\ �Hh4�) p���� ��R���p����v��5yi�M�.������ſ_��)ϿՐ��?;���v�B��Ѩ��q�������o��Y�b�T(�>��P��{]n�=[1�R�	�� ޾����*¤���R
���x��x対�̾�>�����BP�������ʿ���;H����	��
��������n���y�U��p�������{7���࿫��R�N��Q����������1ά��Q���/����N�B��vҿ)���uV���!�� ��uоF㱾Fʟ��旾�����������ݾ ;�"�.��i�F�����忙�"��]�N�����v����s��YD����~���B�L��C.׿�����Ŀ�z���2*��Ed�:V�������m��T��_×���x��<��w����*��[�I�Z(�!��>$Ծ�h��Dޫ�K'��R꫾�g����Ӿ����l��ڜF�!���\帿>��(7���r�`s��
J�����r�����&ll���1����̿�%��?6տ��MR>�%z����N���7���J���&��Vf�K�+��o��(H��7u|���?��l���&�پ|�þ��`{���j���AѾ��u����.� Ra�󅗿�.ӿ3��<sL��+��(��� ���ͯ��������ҞY�G}!����A�Ŀ�H¿�
鿈�� �R��X��m��������ۮ��a���B����R��I���ڿ�i���Bg�)d2����񾂣Ҿ���_���gƸ��oþ�}ؾ����c��}<��v��J����_#&�!Y`�C���g���EA��z��G՛�R���E�̻��#ݿ<�����ʿ2j��3#-��(g�D�����������'���n���J{�G_?��
�d�ÿ�c���FT�zm&�_+�� 辒�;"۾������G�˾d�侳���"���N��  �  u�y�����<I޿~�>qC���n�o���h�����OSj��=��V���տ�U���&��!\�����D���G�Bs��h���K��Pl��If�:X9�����п�͚���l�q;���t,���پ-���4���_1��n7����̾�r쾷q�ι*�x�T����*������%%���R��i{��?��b���[n��:\�z�-�	�o\Ŀ%��1c��i�������F(��%W�k7�
�����{�~�\�W��)����'ݻ��ˌ�/�Y��-����ώﾕ�ξޣ��w𯾄߱�?d��Mؾ�����u�v�9�li����>�ʿ	�Y5��Lb�RW��t��i���x�8�M��:������t��V6��vҿ�/�aT9�pSg�ha���0��'��u��}J���o�鿇䭿���P
Q�*�:��"�hi־�ž�5��P�ľf־�z��z�%�(�C�N�h��q����+��n+F�r�q��g��iǍ��P��9.m���?�AN���ۿ+^��O6���s�����#���J�=�v�f�������%��y�i��<�OI�~׿ǡ��{���I��*'�|�����p߾��ѾT�Ͼ�Vپ,��!��t���;��f����������4��mO)�v!W�����Q��C���fz��jM`���1���bq̿{7���t��L#ǿB���R,�E4[�����I������������[��.�G��XDĿ�6��Ϣj��>��[��d����!ھ��Ͼ�>ѾZ޾c=��2�B�%�UdG�w��M��x|ѿ�n�Dd8�Ӟe�����X��\����{�ZQ��H"�F��f���j���$��pYؿ��".<�gj�����M���Qr���w�mM��n���P ���ŉ�ql[��Y4��)�~����=ؾ��Ѿ�־���������2!1�/�V��  �  �#��,ߝ��¿U7���t��A4��FI��>P�t�F��y.��v�%ݿ�����&��	�������X���꿞����4��6J�_>P���E�$m.�i��4��g���S����]}�f�V�zL7�`M�"��5��Aؾ��Ծ�������z�*�}H�Q�k�Vȋ��|����ҿ���þ!�*�<�F�M�^O�x@�!�$�g����ʿI|���3������Uƚ��Ŀi���`� ��w=��N�!N�I?�M�$�u���g׿�����(��;�n��-K��4-����r������ajվ�׾(����7��+6��U�s�{�����6��y{俰p�+,,��D�%�P�X�L���8����?������������댿����ٿ�^���,��EF���Q���L��9�S���L��Ӓ˿NQ�������i��wH�r(,��m�/ ����g��e,�|�ʝ��H+���G�g�h�ѡ��|c���Qȿ����-�.�6���K�[�R��RI�N1�Z��㿐����+�����Q:��A������%�7.8�y�M��S��@I���1��e�
��v���ʜ��=����]e��F��c+�#��`p����a���a7����H�"�	<�\�Y���|��V��E����ڿ���%���@���Q��;S��7D���(����ҿ�����F�� ���آ�t�̿��3�$�s�A��3R�3�R��;C�{�(����߿�`������&��S	\��>��$������`���gw��kl�1��)�svD���c�%��������޽���j��1�/��G�T�e�O��<�o���&���%¿n���$����Ӓ�C��{߿�.�3�/��H�-uT��PO��;��S����v�пK���"鎿�Ht�úR�6B6�-W����t����)��XG��/O
��6��3�U�O���p��  �  z��H@��׎��8ѿ!B�<����}���
�����k�̿%��]����r_��T���e������¬��Kֿ�)��Y��u� �����	̿\����P�����<m���{o�RM��3.�������3��p�V�"��?��b`��F���;�����0��=¿��ڿX����k	�H��.�����鿯$��醘���w��"Y��xW���r�6����j���i���\0����r�
�)���hYݿFĿ����[���k��ं��Sc�`�A�x�$����1��z#����,�� K��m��ڇ��}���7���^���˿����i�����M��Z����+ݿy����ʏ���n�Z��jb�������`I˿�����-�����%��\�Ko����׿�����宿����5������_�b�?�B�$��U����J���d#� �=�	^�IV��5ސ������Į�H��(�ֿT��g��~4�Z����^f��Muҿ��,���wk��A`�Xr�?���'����ܿek�q����
Y������ҿ����`K��ʞ�饏��K~��\���=��&�0.����D�u3�P���q��߉��ә�t���{���'�ʿ�"㿎 ����Q����i�
��F�Dǿ����V����Hi���g�䆁��Ü�6�¿@������G�!����sq�J��[i̿5�������⚿��6t�ՖR��a5�iE ����a%��,$�+d;�~�Y��|�hڎ�S��������ѿ�7�_��������I����_����{���e�.n�����Ǩ���п,\����	9������
�͕���/ݿ!�ſ�"��$G��,f��%���j��pI�1�.�����>����C,�TRF��f�q���┿�  �  ^Ϳ6ѿ5gϿ��̿DͿL�ϿEѿڳ̿ꬿ�͚��0-����p��@H��/�q�'��63��4P�F{�<�����,�ÿR�ο1_ѿ�JϿ4Ϳ��Ϳbkп�4ѿǂ˿H���fᦿ2����i�W�C�|%-���(��7��#W��������@��;Mƿs�ϿV{ѿ�Ͽ2Ϳ�Qοѿ��п��ɿ�蹿1٢�����b���>�A<+��'*���;��]�����ݟ�fn���LȿrSп��пq8ο.�̿�Hο��п�Ͽ�Jǿ9쵿���|U��+�Z���9�/Y)��+�{�@��e��������#��ʻ˿�ҿIWҿi�Ͽ$�οH�пӿѿZǿℴ���������CY���:�G�-�G�2�ߠJ���q������_���L��ppϿy�Կ��ӿ�!ѿ��пf�ҿ��ԿP�ѿ�Xƿ���r���%U���V�ʪ:�qx0��9�=zS���|�~�������ſ҃ҿЅֿ��Կ�mҿ(ҿ4	տ3zֿi$ҿ�,ſK1��ޖ��%|�iT�;��3�q�?�-�\�������8���gfʿ�տ�VؿCֿ�	Կ��Կ�X׿�.ؿ{�ҿ�AĿLZ���唿v~y���S���=���9���H�ADh�˜���U��&�����ο]qؿ�ڿ��׿��տ��ֿ�\ٿfIٿ~ ҿ�¿m��O(����r�j�N��b;�:L:�\�K�#�m�0������є���|п{�ؿ�+ٿ{�ֿ�տ!�ֿ�Eٿ�Uؿ�Ͽk������ˌ�E�k��TJ���9�{�;��rP�@u�瀒��M���ÿS�ҿ`<ٿ��ؿMMֿ�[տ]׿��ٿ,�׿B�Ϳ4
�������숿c�e���F��u9�'�>��"V�\}����ð��ƿ��Կ��ٿ{�ؿqIֿ��տ�2ؿ&+ڿ	׿l�˿����i����A��*`� &D�v�9�(B��g\�O���ԛ��-����ɿ�  �  ���8���뿄�Ͽ�����|���̙�T���X�t�L>R��V2�������-�3|����,;9��Z��f|�1i��E���<���F��D�տq��tN�������������ƿ�N���t��*\��U��cl�3X������,�ݿ����v��l����-}��Fȿ{𳿥��[m���ⅿ#j�]	H���)�����������ʧ&�D,D�^�e��܃��������Q���Vſ��޿T�������H�����Y��混��s���o��4V��Y��@z�ڟ������K�������~	�Ί���ڿ~Q¿ï�!����������� b��4A��_%��%���	�&p����}5�>1U��w�C���웿;����G����п�6�6����]<�M������w�׿P���������l�	�\��i�Ỉ�����jԿ������
���������FGտ����"譿-=��H9�����f�]���=���$�����h�����*��8F��Xg�Y��D��O3���3��`=ſw�ܿew����
��;�H��y��8��f�Ϳ�[��������l���f�!�}�����6[��rE�q�X�������$������пRI���Q��z���G��eVz��JX���9��=#�������1!���6�P_T� v����2���]T��|�,�ͿD��@��@�]5����	���=꿬;���Vc����f�/0j�k4�������ɿ�l��`��W��u�����+���L�6�ȿes��sU��2���𕈿	 o�=�M���1��N�k��� �(�K�@�L&`�6��ݑ�����ï��k��pֿ�i�D�M��D���2�ƅ�l�ܿ芳�\X��\Kv�f�K!s��L��?a���Kؿ#� ���  �  �:P�%cH�,�2����/�3}��?������ \�:�;����#���x�	پ��Ҿ�ܾ�q������%�\�B�ǥd��k��Y���a�ʿi��������8���K�E�O�!�C���)�G	���ӿ`f��w�������3˕�q����^��Ҏ�0p9���L�~�O��B���)�\
�*࿳���j��;�v�B�Q�i�2��w�H��L�W�־/�վ0���� �����K/���M���q�,я����Y2ڿ����g&�^4@���N��kM���;������������P���r�������<��e�Ϳ����&�N�A��P���M�|1<�f� �U��v_ѿ	���ꋿҐl�J�,-�ɓ�lS�����/޾�+�o���9��I�#��F?�E�_�fI������=���"�gZ�(�1�	�H�)'R�E?K�%B5���&X�������އ�B�����$���X�2��J�o�R��#K�g�5�k������m�ſݫ���r�� g�!�F��!+��?�*��O�}뾆�����o���13��8P�4ar��Y��󋪿%ѿl� ��"<��5O�7�S��DG��z-����ܿ�ʬ�
��;;���w���6ſ���*���=���P��	T�w	G��.�CE�]�迥����h��m����b�<C�=�(��B����������i�j�i�%�_�?�}�]�	��j���f��J��S��K�*��oD� S���Q��5@�5-#�>�&ʿ���������mv����տ��	��M*��_E��S�`!Q�q�?�y&$��P�v
ؿ����ŕ��'�y��2W�h�9�~?!�f���� ����W���k2���B�.�\�I�2 j�+x��0ߡ���ĿF8������S4�%K���T���M�g�7�o���1�պ�[ʘ������_�����Қ鿡����4��&L��  �  �c��f��w�l�}�@�E��ݗڿ�����v���A�&��c!�Qݾ�����������Ʈ���5Ǿ�"�+��jm$��SL�_ۂ�W&���H꿗��tFK�cu�l҈�N<��vփ��wc��N5�5����̿�p���{��𷿯��A� ���O�>�y����+׋��%���*_���1�c"��ƿ:蓿|�c�F5�,��ʐ���gԾ�޼������������оW����<o0��-]�s#��V'��֊� r,��Z��Q��,��<����%}�y`T��s%�K�����*(��Q���X�ƿ�!�4/0�s�^�y��>1��K'���3z�,Q�xU#����­�������jU�6',�����$��Ӿ�j��z����}���˾�`�ue��� ��[D�"w�軠�1'׿?����=�n%j����M���Ȉ��s��G�0�����iʳ��d��c����ݿ��B��o�Q݇�����CŇ��mo���C�g�8�jo������d�L�a(�n����}YپN�ɾ�ƾ��;���K��z�(�1�DZ��ȉ���7=�� ��N��x�ђ����볅��\g��[9�����iտ����4��b���/H��}%��S���}��������JJ���lc���5��U
��_οP3��/<t�!{E�]N$��
�����8ݾ/�оA>о�۾�:�|	�V� �Ѿ@��m�_���nǿ���(�0�O^��o���L���������T�X�f�)�@���קĿŷ��6���,Ͽ�9��&4�*�b��J�����d؋���}��}T�Z�&�Ѿ��[���;����b��@9������m�<�ؾǀоH�Ӿ�������F��5+���N�>���᥿�Kܿ�{�E@���l��V��\���"����u��sI����K鿺}�����k��}p⿄J�PED��7q�Q���  �  ����J��d���|�l�=1�Ͻ������ƫz�F9��]��.�/���a����gw���S��m	��]ƾm�e���E�%�������Z��C>�*Az�k6���$���s��B�����	�_�F�%���!���C����׿���
E��}���	�����������4����X�6���߿�*����b���)����׾ZӶ�Oc���A����������æ����Ҿ�� �?s$�b�Z�� ����ֿ.���Q�ջ��Re��I"���m���R�������GK����$ݿm����G��� �=�X�N)�����3M��U���o)��bр�R�E�Q��.ȿ8卿�P����������Ҿ`���ͦ�����jͣ�����,Ⱦ��쾴����:��ey��
�����(�,�6h��ɐ�.d��^���.��������u�1:�3]�qѿ�J����̿z���4��0o��������\���y������o���3�� �Wf��OȂ�zD��{����n�վ�߽����4��mn���ľp7�`��L$�a{S�3�:�ſ���Q�A�̹}�������?C���̥�m����c��7*����� �ɿ�����w࿿|�|mI������6������T��Iӣ����&]��I#�ZE�u��\s��3:�U���-��k?׾�¾̑��-���������Ӿ6�:>�A�4���j��<���߿,��/V�׈�����9C�����x�����0�O��I�#��pS��'�ſ����F$���\�,���������	k���՜��{��:�H����%�ο����H]�^,�v��$(�<�Ͼ�*��pa������gǾ{b޾>��W��2E������/��M���c}/���j��������ܰ��+��>��-x�ܐ<���
�W�տ�����/ѿ�;��e6��oq�75��/����  �  �@������SY��m���bH�sb����ޟ��8�[��.վ��8ɗ��x���4�������3��Nu�����i���XF�ی��aο����CW�����#���#������sѺ�����~��U;�S��ӿ��ȿ)|��!��j_�^>��ۦ��ћ���m���~��R��5_v�z�2���������Hg���&�j��U5Ⱦr����(���܊�cQ��w��`{���Gþ�_���� �^�F���Y���x+�nWn�n������:���f����I��Rѕ�*�f�r�'�4���ʿ�qϿ����x4��Lv��J��,�������d������������_�<	��Eٿs�����Q�[i��/ﾉ3þ;���꘾6J���J��89��gĸ���ݾ�����8��J��Hܸ�����B��ԃ���	���Z'��ϑ����������R�Ml�t��,˿��$(��hK�Gه�"����������D��k���O��i�J��o¿����C����]���ƾH���|���Ġ�����"ᵾիо���O�uT��Ǔ��Vտ�A���Z��D���l��N�������ʹ����������?�����nܿb�ѿV��Q4&�/�c��m��~Ӳ��������������r����z���6����Z	����w��/7��S�]����Ǿჴ��,�������Ʋ���ľ����p
�=/1��qn� ʧ��=󿼢/���r�Ĺ��:��@�������<o������ k�f�+�����ҿoؿ���W�8�kez�7A�������|��В��Ǫ���c��c�~`"���߿�<���^��'�=��"�ܾ����~G��d�������︾.�ξ�A�K�uC�Qx�����
��+E����>V��&���o������Cά�ǩ���T�������Ͽ�P���Z�M�$������ ���  �  AH��,������lf��/+�du��⤿F0d�!�"���ǟ��s晾s}��̃u� �o��'y��c��|���qƾ�� �S$/���w�]���t��E8��\s�3^��&�����̑��U-��( Y�r� ��j�%����챿��п����'?�ަy��֖��$��y���ʪ��,X���qR��4�n�ԿX���
L�Nd��i޾�c��3���ԋ���t���s�����ϐ�d���r�׾, ���C�&ዿ	�˿�/�.�K�p)��2m���ը�i��w��1��V<E�#`��3ֿ�ֲ�0L������5��R��I��f̝�!���y��FG��	�z��m?�B��Z!��<����9�`����Ӿ}߬����/؇����}����.�����e�ľ���2$���b�8������m�&��da����jM��e4��4���Y���R�n�(�4��/���ʿ����+ƿ�����.�gLh����?�����5T��I����h���-������R���o��-����7Ҿ�谾5���뿒�+u��U���%��E����ྐ0�j�<�R����������;�a�v�X����%׫��s��:&���]��"%�.
���pÿ����ٿ;���C���}�����K������,̟��v��ΧV�ed��ݿQ��a|\�)�#�	���f�о:糾ע�����3��0M��T��IV̾b��yg�MT�����ӿ�V�`�O�C��ǉ��.����"��:����q�I������޿�v��῿)�w_���V��9��s���m����,��S����}��B�29���ÿ�_��#�F�l��v��0ƾ�٭��*���̚��Mߦ��4���Vھ�����.�t<m�������@)���c�v`��ܗ��x|��Ħ�?ؓ��q�7�.�� AϿ�3���ʿa1�>1�B�j��'���N���  �  ��h�������H\�He$��S迲Π��a��S"����n��M���~��7+}�`w�np��7o������ɾ���p.�Ȫs�5ɮ����m�0���h�����������\���CW���O����Q� +���Ӭ�*ʿu�d7��o�Gc��5����G���Ԗ�����O�I��a�,ο����J�������[_��~���}��Pu|�a{{�����I甾_����ھ���:^B���7�ſ$��'C�g{�w���?����Ġ�������t�*=���
�`1ϿC���^걿�ۿ�>��I�����n��F���>�����|�o�e�7�_��z᷿p���4�8���	��d׾4���1������Ȇ�!��� )���#��b�ȾP���5$�O7`��9����⿺v ��W����M���أ��m��/c��3�d�z-�����`Ŀ"{��s;������e�'�̬^�w����?���C��-C��q��3_�'�#���>���l�
S-�5���־�������
����6�������������T�98�#<�����t���2~�4��jl�I���/���$������GN��BT��������۽�M���4�ҿ��
�|�;� ss�L�������k��
���_�����M����}ֿ�<��g�Z��($�����Ծk��2Ȧ��{������8���0��\о�I�����L�R��O��2�Ϳ!��7TG��8�˖�j���<������,y�^wA� @��׿�I��Sy���q�d���M�q������{S��K��yg��Gs���:��O�s����"��'�E����� ��Dʾ�鱾���|�������r۪��Q���6޾#�ۮ.��j��]����9#��Z��O�����O!��@�������~g�r�/����jɿ�-���Ŀwr���(*�Z�`����M���  �  ڼ�������o���A�G[��+ӿi���C�Z��#�i���u�̾����d������Sv������$����M��˔־X/��M.�0�j�⎢�������4�L�X�x�Y�����������f�X`7�7�	��0Ϳ/֥�E���B���ͭ�@9"�"BR�cX}��3���,���'���a��2��� +��؂����F�ɣ��*�����b������o����v���H��]���a��\���?��q��	۵�tH����,�@e\��D������������8W�s&'��E�������j�������ƿ���72�#�a�逄����qm���}�<S���"�4<�ʊ����v�|�7�6��	����G��"��[����~��8�����վ۾�Z�%��Z�4���>ϿiQ��>�:m�(���������E�v��vI�����W� e�� ���6寿ln޿�7��]D��r����m��k��ۃr��D�J���ؿ2���ve�q�.�i
��I�+�¾߭�-���u���5���W"��\m̾�0� ����;�Eqx��z�����;7 �RP�QI|�Ќ�k]��ȇ��j�xl;�5����տ�v���f��uu���b���&���V�Հ�}Z���P��[I����e�M6��.��|ſ�Ǐ�M!W���&���Hk��vž�^���^��eө�Y�����¾�޾Ҧ�WK"��1P��������"K���0�[�`�a�����"��������[��q+��n ��Ŀ{���ی��AYϿ�	�$6�e�e�nS���A����O����RV��*&�����o,������D�<��X���l�׾���}Y��uZ������������˾?��f��w0�2e�J'���aԿ3���A���o�t��h��B��(y���K��`�"꿨���E��������;�F��t�&���  �  9e�<�[���A�����3��.X���܋�F�W��K+�L��ٞ�bdƾ'���ѡ������l���J���;w\�0��Q4���d�������ſP���J'��	I�B�_�Fe�d�W�7g:�Ѝ�^�a��� ��2��������ɿ�1��v*�[4L���a�ױd�HU��77����࿔��ro��m?H�� �����ݾ
��h��T����
��L���=W`پ�� ����ߥB���x��w����ٿ*���3��R�ڔc���b��O�vH.�`��o�Ͽ�3����������Ʃ��lݿ�����6�	�U�yUe�= b�3M��0,�����ο^k��9�n���<�c�"���ھ�W��𝮾�ާ��J��7Ǹ��&о���u���.���Y������b�������Y@�է[�T]g�T�_�~HG�I$�����h¿7�������:ޘ��̼��U���( �:1D�o�^��4h�%�^�)�D�ܴ!�#���	˾��M����b�.K6����;:��;iݾ�	ƾ]���9;������̾��zw�͟�1�A�M`r�����̿�c�<�*��|L�HNc�5�h��K[�V?>���g���������6��&�����ҿN�	���.�q�P���e���h��TY��t;��9�>C鿗Z��f����X���0��B��<��e߾T�ʾc쿾/G��l�Ⱦ�6ܾ¸��q7�>�,�D�R�W���{���k������Q7��LV��g���f�RS��2��:��'ؿ��������z_�����j���y���:�<Y���h�D~e��gP��|/��
�¯Կ#���|���I��l&�����]�I*ؾ��ƾo���ސ¾c�Ͼ�d�X��vU�%9���c��������0����h���B�tC^�D�i���b���I��x&����-�ƿ�>��Zl��Z����c�������["��SF�ӧ`��  �  +���$�
������:�˿�/��5���N�c���A�n�%�	������}վ��¾鮽�e"ƾ��۾)B������+��I���l�ύ��M���ֿ�p����'��*�r� ��3���俆h������=p��&h��xޠ�J�Ϳ�����(�O�*�� ����E��.���0A��H�X���8�D����s,꾃�Ͼ3&���Q��1;~V���?��G5��+T���z�~9���Ź�]忪
�]|��)�u�(������-ӿZͤ��%��g�h�~
m�#]��X���3m߿��	�B���+�sc)�?��@����ܿ�&�����u��mP���2�B������V込.Ҿ0�Ⱦ�B;k߾\���a��)�3�E���f�Aǈ�QR��$˿����k�t%�;-�f'�w����a�ƿ���kO���n�n�~�I���'¿�������?�&�=�-�C�'�R��_q���gѿ����*��>�n���L�Z�0�/�	a�%��+�ھ_"־K߾!���!��R ��_9�%�V��z�����9��X�ܿ���� �n+�4n.�r�$������I���"ꕿ5u�� 2y�;��� }����ֿ8W�@�:b,��/���$����*���ƿ@��)�����h�1I���.����^C����~e�#��nU��N��=��v+�^�E���d�h����z���¿	x�M���"��7.��-�q����\�ۿFL��0���x�y��}�����������N���%#���.��,�����9	�`n�9ƹ��H���&����]���?�L�&��h�^� ��}�����T���	���@�4�� P�Sq�Rw���8п#�����o(���/���)�ZX��
���˿M������Ox�b�����KwƿhU�����>�(��  �  р�N￳a޿a�ǿI��$����m��/q��GU��[8��b�F��t,��OS�����X�2A#��?�V\���w��m��y%������	��EyͿ�@�9����t�Kɿ�	��\&����^�	�A�n<��O�~x��_��[线G�ٿ�|�;O���0뿾�׿\��� 4�����H<���Ɓ�i�!�L���/�JE�V��#��n�ﾩ;����5�,��
I�~�e�h ������J���Tȩ���q�Կ���{�h�(ܿ"������W}�[�Q���<���?�8�Z�JK���㤿ƠƿI��n��,���翮�ѿ�'��7����n�������6~��0c���F��*��+����/�������P��!�b�;��Y�ru��Ǉ��Q��.C���ĳ�/Lɿ��߿6��k����x�d׿Z��
����t��P�V�C��N�i�p��9���$��U�Կ������ʑ����㿜xͿ����x���`��2⊿�0|�\n`�ѰC�$�(��v���U]�^��r��:30�f:L� si����+Q�����I ����2]Կ�&������������r�п�ǯ�����o�0gR��GM�>!`�����F����ÿW�3���������KG�?dɿ���������
����yy��\�i@��q&���������=Z�Ǽ#��<�	AY�]�u��K��Ɣ���G���jƿ�?ݿ;^� ��� �����\�ƿR�� ���?�b�}xM�	.P�k�j�o���v��h�Ϳ/�J�����h���\ؿ�����Z��`���A��𯅿�3p�yWS�$V7�?��q������
�5C��:,�K�F�Z�c����4����x��%h��S�}ο�'�=�������m��ܿ���u�ء~�M^Z�<M��W��y������m��ٿ���  �  ɂ��*J��|���
������ñ�R���=��U��r��[�z�c�Q�"#0��������l�6�5tZ�I#�����������Cò������C�����c���f��1E���/��j���t�e�K�zR,�9���*H"���<�U�a�����cڙ�騿�����t����i���'���β��+���뫿����ϋ�tUm�N(F��\(���D�ۼ%��!B��wh�uY��s���J������ʘ���������v����{��3��,��� X���ڇ���e��?�$��y����#�)�s�H���p��č�a���!��������6��"�����v>��Ì��_b��*䩿y��������c�\'?���%�w���U�� 3�îS�\l|�?Q���L��������ε��!���ӳ��O��\I���4�������:���؄��J`��e=�*4&�F����$��;��U]�Qi��bA��E^�������η�V#������畵��4�� �������ר�'���7�F#]���;�'��$!���*��eC��Pg������1��La��YӶ�Ӯ�������-��O���rK���\���V��\j�����w���A�[�/i<�~*�q�&�#3�	�M�%�r�����m��*z������Ƅ������ո������ ��/p���#���ڦ���:�}�\TV���8�~%(�;'���5��CR���x�t��G�����������\غ�RD���R���]���亿+���T#��ͣ��L���Xv�WcP�B�4���&���(���9��7X����� �����]���i���ֺ�.��?���๿i0����qu�����%���p�g|K���1�%�&��+��>�9�^�������������O�����}�1J����-���4����m�������V��t߉�)j�MG��/�+'�'.�i�C�0f�����b��Ig���  �  D�����������%7���Cɿ��߿Y�￳n�i���οlV��7Ì���d�J]D��;���I��Go�^�������ԿC��-.���W��7ۿςĿ�*��{靿�&��)����`m�i%Q��N4�����y�����B�w��P��>(�AoD�FMa�dd|�I���֪���+���Ժ���ѿ���w*�5��q��JĿ����!����yX��O?�u�=�(wT�cb��p����R����ݿiZ�~�0运�ӿܼ�ߵ��BĘ�y���TT~���c���F�{�*�Y��.' ����0��V��t���2���O���l�����R���ꝿ�����ÿ��ڿُ�����^�dڿ����~�����y��R���@�|�G��<f�k����׬��ο7��R���m����忲�Ͽf��N����� U���]}�D�a��,E�8�)��?�oV�������� �"y(���C��'a�@1}�ez�����5~��������οq��2��p���%� �ӿ`������g�p��VP��%G��V�I�{�N������yۿ*z����@���$�wm˿����Ӥ����J�����{���_��pC�N�)��^�y�	��������� ��:9�_~U�er�󽆿I��Q+��b���?ÿ��ٿ���Un���������\=̿���Ֆ���h��mO��N�z�d�0s���զ��lȿ��A���l���%o��ۿ-0ſ���*�����	����bt��W�[C;��"���������w��Q�'�x�A��L^�Y�z����(��+����\���Xʿ�.�z1��g��������v�M���ݟ������$^�0�L��S���q�%;���e��u�ӿ�/�����2�����P�Կu���Z嫿�.������ރ��/l�-BO�j�3���#���<��������1�R\L�7^i�l����  �  �e�����	���Rο���,�\�%�+�,>#����2�X��������4t�"[f�j.|�N���hſu��� ��4&��"+�,�"��s�b�(5ſ2������^��a=��""���
�WH�l�ҾLk¾9g���ʾ�~�}��r����0���N�8At�V���򵳿=�ݿy�C���&)��2*�n$�^&�N1ܿ�9���ꈿ7^l�Zj�`7~��YYֿ(C�7��])���)�t�����Ő�����s���!x���Q�93��k�|��F��=�˾���]I¾�Ҿ�3
��!���<�]�n�!��'W¿.���'/"���+�<f(�T��� �YIͿ��b��xwl�ǌv��A���U�����^#���,���(�`5�C��L׿T׮�Xߏ���q�՛N���1�މ�u�^�꾆i־�LϾ�վ��龥��p�bs1�@�M��p�;���������ӿI� ���[(��-��&�������n���Ey�����ur��5��j�����˿�y��j���)�(�.�Z&�����J���̿�릿�6l�,�K��0�������Q�ʉ�M྿8�������(��B�u`�j���,���*���?濫�
�J��H-�'N.�V:"��7�eL�;O�� ����{|��uz���������lm޿�O	�a �er-�J�-��!�����r翿_֝��w�� �b��D�l%*�-#��v�F�3྾����l�!��E�/��J�Țj�=�������v�ȿ0|��C0�2}%�&/�L�+�t�����jxӿT��X
��cx��+�����c]���+�����
&��U/�Z+����v�!Jܿ���Y���=|���X�.<�x�#� �K���j��ᾪ辿k���1��o!��9���U��  �  }�Z��荿F��Q����!��C���\�U�e���Z���?�����y����%��<z��o������cA���$��G��_�ee�P�X��<���Fp���������O�i�%����"|㾛þh۬�>����X���H���+��cԾ������{�;���n��I��N�Ͽ���n-��M�f#b��`d���S���4��b��ڿbҧ�/��� ������Qӿ�8�N�0�1�P��Oc��4c��P�=81����ֿ�Ϡ�gu���?�dO�;���/�־$!��B����.������ꬾ^�¾8�⾓H�e�$�DwM�ӻ��{3����1��A�9�I+W��e���a���K��k)��H��ɿ���é��Z���u|�����{�o�=�gZ��#g��`�4I��'����uJƿ�=���h��n9�W	��w��ξ۾��¾����Og���x���¾<�۾�����g��7���e�1n��p���w����#��F���_�?Gh���]�÷B�^��w������%��Q���?̞�?�ƿ�=��E'��TJ�9Tb�?�h��!\�V/@�Rt�-U�Q��� ���^��A4��v�~� �2��(̾�o��ʾ�s6ǾY~پ�����S���(� �L�N��Ť�VCؿ2)���1��R�zDf��{h�(�W���8��o��!�i㯿�����-�����bۿ�B���4���T��cg��Mg��T��[5�����p޿/��t肿W�P��
+�N��������ھ-�ǾK��|.���u˾��k����q�7�2�U[��i���ѳ�^��)�:2=�ptZ�X i�(�d�-�N���,��X��Ͽ����g���Ύ���Y��qg�����@��]��i�BEc�ǲK�R�)��Z���˿w��s�E�C�}K"�&�	���־�ƾ������ž,)Ծ�쾦�����?��  �  �^�^��I׿�����D�Xr��;��|��������m�KK?��}��ֿ�ԩ��[�������俹h�� J���v�!���j���Ã��y�h��:���]�ǿ玿#pP�	����J�Ǿʳ�����ъ�,��<�����������J߾[�D7�d�w��2��d��$�J�T�s�:�������|q��?@_��e/�����yĿ�w������d��� ���*�-Z�A���SV��+=���e����Y���)������\�����#g<�b��b��<���Ǡ��ݐ��󉾉���!���}쨾�5Ǿ����%�˓L�vd��r?¿*$�(�5�8�d��g��(Ҏ�y1���D|�2�P�� ���U෿����1����ҿ�6�r;���j��x�������^���kx��K�����5�'��d�m���2����p��.���Y���B��.&��m��mJ��k�����%�
�-�0�5i�<䞿��ܿ����hG�y�t�����!���u����p�V6B� t��ܿ֯�aa���������{�*BM�<z��B���P��6��~Rl��}=�$����ο�ڕ��^�gQ+��[	�OM��Ǿ�/��Ѓ���F���Y��/&��@ھ� ��L��>H��j����������(��Y�J����������|��	Qc��r3���Ί̿H������;ǿ:��n.�S^�����`��XI��Ut���^��.���&����Z��c#M��D ��K�1ܾ�c��
��/���w���u���S�ƾf!�"'�	�(��Z����G�ȿ�m
���8�:h�����o��oɍ�Ff�1�S���#�
���ٽ�	�������ؿ�!��O>�M^m�RԈ�6ؐ������ {��N�j��~l迣U���=x��Q=��)�����e�Ծ�{���?�������v��Gٻ���Ѿ���^�;�8��  �  �5e�D�� ��]'��n_�f�����5��4��!h���2Y�w�"��P�`繿�J��T¿���O.�ɻe�L����$��Т��������S���~�ڿm���B\U������꾢��k#���`����}��hz�<��ܸ���ܪ���Ҿ�k�B�8��u����������9�lDr�����k��c���ߕ�}~�l�F�O��)ٿ�6��~���ҿc���|@�]x�{����E��Q:��x����x�K
@���
��z���A��A�>���UC׾7���؈�������v|��t�{��h�������ĳ辥��րP��F��E�ӿ���Q�M��e���6������[������."m�'�5�P���ɿǶ��%-��-x�g���wT�Bw��c��d�������x����g��U/�˜��=ͮ�</v���2�NA�Y�־��������/���c��	X���\��q��k�վW���/��5p�܍��Z��*�)-b�Hl��2	���Q������B؈�="\���%�WP���꿿�M���Wȿ ��[1���h��A��ğ�y���:��+r���mV�_9����)���.jc�h=)�����׾�t���X��r��v_���磾�в�rJ̾�y���V��}I��B�¿�
��0>��qv�����@{����� �������J�����%�E���)����ڿ4��U�D�[+|�Õ�rO��QF�����@|��1D�	�\�ɿ5���7:O�Z���g��:�ξn��䘤�/ŝ�����[����ɒ־jo�{Z&��^�n�݄ڿ?�q�P�Y��cՙ�����w��B��.p��8�YL���Ͽҫ���!���g��!�[W��߆����������F��܎�r2j�W�1��������}N���=�ł�f����ƾjn������埾l]��Y殾�,ľv��#�G�7��  �  o�h�GJ�� i��zR.�Z\i��O��0ţ��J���+���p��5�b�r)�	������!S����ȿ�S���5��o�����?���*�����������J\��"��N�G7����W������羽2�����_g��\v��r�_�~������˦�{UϾ��9�9��Ӄ�K�����
�w�A�� }�� ��Ȭ���Q�� �������qAO�>�����t����U����ٿ�?�׷H������W��䇨�K����^������SH�yO��bǿ 房��?�al���Ӿ���z��8�����t�E�w�:.���q���ʵ���YC�ۚR����d�ڿ��<�V��C��e��QP�����[��
�w�^$=�5`
�.п�ȳ��о�c��4%�V�]�a]��|E��)��]!�����d�q�Ȟ6�����q���y��P3�)��Ҿ>ܮ�(����=�����������Y��X����.Ҿ���@	0�	�s��Э�����|1�Zl������#��X���'���z��?�e��m,��
��v�ſ/U����οbV�ߥ8���r�����Vݦ��ѫ��/���p����_�V�%��3��)��l�e��)��i���ӾpQ���W��a���m������������2Ⱦ������%�J��N���ȿ���$F���X4��޼���^������᷆�}NS����G�迠����b��N�ΌG�S�L�����V_��u���9���|m��1���{L�tz��Ͽ�B���P������zʾ{���ů�����ݚ��g�������Ҿ� ��	&�!`�_-��M]��: �$�Y�U������_��|�������-�z��#@��Z�grֿ齹��Ŀ������'��`��ƌ�����V���o���;��=qt��89��d�V����-��*�=��i�b-羯�¾*e���8���"������)⪾?��%�⾙���8��  �  �5e�D�� ��]'��n_�f�����5��4��!h���2Y�w�"��P�`繿�J��T¿���O.�ɻe�L����$��Т��������S���~�ڿm���B\U������꾢��k#���`����}��hz�<��ܸ���ܪ���Ҿ�k�B�8��u����������9�lDr�����k��c���ߕ�}~�l�F�O��*ٿ�6��~���ҿc���|@�^x�|����E��R:��y����x�N
@���
��z���A��D�>���DC׾�������a����u|��s����\���U���-�辳���P�"F����ӿ0���M��e���6��~���/�������!m���5��O���ɿ����6-��Wx鿉���wT�dw��8c����������������g�*V/������ͮ�k0v���2�&B���־������������c���W���[��{���վ����/�d4p�0������2*��,b�l�����OQ��͛��؈�"\�p�%�%P��o꿿�M���Wȿ��6[1���h��A��4ğ�=y���:��er��<nV��9����ڛ��hkc�x>)����D�׾
v���Y���r��`��b裾	Ѳ��J̾�y���V��}I�"�C�¿�
��0>��qv�����@{����� �������J�����%�E���)����ڿ4��U�D�[+|�Õ�rO��QF�����@|��1D�	�\�ɿ5���7:O�Z���g��:�ξn��䘤�/ŝ�����[����ɒ־jo�{Z&��^�n�݄ڿ?�q�P�Y��cՙ�����w��B��.p��8�YL���Ͽҫ���!���g��!�[W��߆����������F��܎�r2j�W�1��������}N���=�ł�f����ƾjn������埾l]��Y殾�,ľv��#�G�7��  �  �^�^��I׿�����D�Xr��;��|��������m�KK?��}��ֿ�ԩ��[�������俹h�� J���v�!���j���Ã��y�h��:���]�ǿ玿#pP�	����J�Ǿʳ�����ъ�,��<�����������J߾[�D7�d�w��2��d��$�J�T�s�:�������|q��?@_��e/�����yĿ�w������f��� ���*�/Z�C���TV��-=���e���Y���)�����]����)g<�_���a㾌<��7Ǡ�-ݐ���T�������v꨾3Ǿ����#���L�Bc��>¿q#�d�5�p�d�>g���ю�'1��wD|�ǩP��� ���෿����R���e�ҿ�6�fr;�p�j�y��ꅏ�0_��Plx���K����	7�q����m���2�]����!������NC��<&���l��7I������㾈�
�8�0��i��➿8�ܿן��gG���t�����L!���u��4�p��5B��s�*ܿ�կ�da��&����5|��BM��z�&C��Q��o6��WSl��~=���+�ο5ܕ�|�^�wS+��]	�;P�3Ǿ�1��P����G���Z���&���ھA� ��L��>H��j����������(��Y�I����������|��	Qc��r3���Ί̿H������;ǿ:��n.�S^�����`��XI��Ut���^��.���&����Z��c#M��D ��K�1ܾ�c��
��/���w���u���S�ƾf!�"'�	�(��Z����G�ȿ�m
���8�:h�����o��oɍ�Ff�1�S���#�
���ٽ�	�������ؿ�!��O>�M^m�RԈ�6ؐ������ {��N�j��~l迣U���=x��Q=��)�����e�Ծ�{���?�������v��Gٻ���Ѿ���^�;�8��  �  }�Z��荿F��Q����!��C���\�U�e���Z���?�����y����%��<z��o������cA���$��G��_�ee�P�X��<���Fp���������O�i�%����"|㾛þh۬�>����X���H���+��cԾ������{�;���n��I��N�Ͽ���n-��M�f#b��`d���S���4��b��ڿcҧ�0��� ������Qӿ�8�P�0�5�P��Oc��4c���P�D81�����ֿ�Ϡ�{u���?�aO����ֿ־� ��a���O-��F��笾��¾���cF�˲$�@tM�����1����#��0�9�?*W��e���a���K��j)��H�lɿʙ�����������|��F�����=��gZ�q$g��`�J I��'����sLƿm?��E�h�zq9���?{����۾ݨ¾����bg���w��8�¾��۾����He�F�7�l�e�Zl��j����t��m�#�~F�p�_�AFh��]��B�ҍ����������$��V����̞���ƿ>�^F'�JUJ�Ub�G�h��"\�|0@�wu�aW�b�����U^��D4�@y��� �����̾�q���˾��7Ǿ@پa���4T��(��L�]��Ť�WCؿ2)���1��R�zDf��{h�(�W���8��o��!�h㯿�����-�����bۿ�B���4���T��cg��Mg��T��[5�����p޿/��t肿W�P��
+�N��������ھ-�ǾK��|.���u˾��k����q�7�2�U[��i���ѳ�^��)�:2=�ptZ�X i�(�d�-�N���,��X��Ͽ����g���Ύ���Y��qg�����@��]��i�BEc�ǲK�R�)��Z���˿w��s�E�C�}K"�&�	���־�ƾ������ž,)Ծ�쾦�����?��  �  �e�����	���Rο���,�\�%�+�,>#����2�X��������4t�"[f�j.|�N���hſu��� ��4&��"+�,�"��s�b�(5ſ2������^��a=��""���
�WH�l�ҾLk¾9g���ʾ�~�}��r����0���N�9At�V���򵳿=�ݿy�C���&)��2*�o$�_&�N1ܿ�9���ꈿ:^l�Zj�b;~��^Yֿ+C�;��])���)�|�����ؐ�#����s���!x���Q�}93��k�G�����/�˾��LG¾�	ҾC1
�]~!�ê<�\]�V삿]���T¿���Q���-"���+�@e(����l� �\HͿ/���Pwl�5�v�E�����꿠�x_#�¸,���(��6�����׿�ٮ��᏿��q�N�N���1�.��0���꾹j־�LϾ�վ������/��p1���M��{p�����@����ӿ������Z(���-��&������}����x�����vr��5�������˿J{���j���)�Y�.�c[&�+��rM��p̿jZ�&;l�μK�(�0�����T�`��G�9:�~��p��Ҁ(�B��`�q���",���*���?濫�
�J��H-�'N.�V:"��7�eL�;O�� ����{|��uz���������lm޿�O	�a �er-�J�-��!�����r翿_֝��w�� �b��D�l%*�-#��v�F�3྾����l�!��E�/��J�Țj�=�������v�ȿ0|��C0�2}%�&/�L�+�t�����jxӿT��X
��cx��+�����c]���+�����
&��U/�Z+����v�!Jܿ���Y���=|���X�.<�x�#� �K���j��ᾪ辿k���1��o!��9���U��  �  D�����������%7���Cɿ��߿Y�￳n�i���οlV��7Ì���d�J]D��;���I��Go�^�������ԿC��-.���W��7ۿςĿ�*��{靿�&��)����`m�i%Q��N4�����y�����B�w��Q��>(�BoD�FMa�dd|�I���֪���+���Ժ���ѿ���x*�5��q��KĿ����"����yX��O?�z�=�.wT�gb��v����R����ݿtZ�~�0迣�ӿ,ܼ�󵨿UĘ�����eT~���c���F�E�*�����& ������U��r�1�2���O�N�l�����P��0蝿񾮿!�ÿ��ڿ?��Q����\￠ڿx�m���1�y�R���@���G�>f�R���٬�, ο3�迡���������忈�Ͽ�h�����y���fW���a}���a�o/E�/�)�6A�W�9�����V�Aw(�3�C��$a�R-}�x��6��s{��������ο��50�������^�ӿ�
�������p��UP��%G�LV���{�a��z���u{ۿ_|�w���B���'�vp˿���֤�����Ê���{��_��sC���)�r`��	�������q� �e;9��~U�?er����I��T+��b���~?ÿ��ٿ���Tn���������\=̿���Ֆ���h��mO��N�z�d�0s���զ��lȿ��A���l���%o��ۿ-0ſ���*�����	����bt��W�[C;��"���������w��Q�'�x�A��L^�Y�z����(��+����\���Xʿ�.�z1��g��������v�M���ݟ������$^�0�L��S���q�%;���e��u�ӿ�/�����2�����P�Կu���Z嫿�.������ރ��/l�-BO�j�3���#���<��������1�R\L�7^i�l����  �  ɂ��*J��|���
������ñ�R���=��U��r��[�z�c�Q�"#0��������l�6�5tZ�I#�����������Cò������C�����c���f��1E���/��j���t�e�K�zR,�9���*H"���<�U�a�����cڙ�騿�����t����i���'���β��+���뫿����ϋ�uUm�P(F��\(���H��%��!B��wh�{Y��|���V������ۘ��������������{��C��6���"X���ڇ�_�e���?��$��x������)�g�H��p�'Í�u���箭�+���E4��R����𱿯;��%����_��⩿����P���ބc��%?���%�L��[V��!3���S��n|��R���N��=�������е��$��oֳ��R��L��S7������V<��#ڄ��L`�g=��4&�V���$�L;��S]��g���?��-\��{���7̷�t ������꒵��1��m���P���cը�g�������=!]�v�;��'�%!�P�*��fC�Sg�n����3��c���ն���������1��`���hN��q_��Y���l��󂖿������[�k<��*���&��#3���M���r�4����m��6z������Ƅ������ո������ ��.p���#���ڦ���:�}�\TV���8�~%(�;'���5��CR���x�t��H�����������\غ�RD���R���]���亿+���T#��ͣ��L���Xv�WcP�B�4���&���(���9��7X����� �����]���i���ֺ�.��?���๿i0����qu�����%���p�g|K���1�%�&��+��>�9�^�������������O�����}�1J����-���4����m�������V��t߉�)j�MG��/�+'�'.�i�C�0f�����b��Ig���  �  р�N￳a޿a�ǿI��$����m��/q��GU��[8��b�F��t,��OS�����X�2A#��?�V\���w��m��y%������	��EyͿ�@�9����t�Kɿ�	��\&����^�	�A�n<��O�~x��_��[线G�ٿ�|�;O���0뿾�׿\��� 4�����H<���Ɓ�i�"�L���/�LE�X��*��w�ﾯ;����?�,��
I���e�s ������Z���gȩ�)����Կ/���{�h�(ܿ������}���Q��<���?���Z�KJ���⤿/�ƿ_㿙l�c*�����ѿ-%������jl��^���	3~�F-c���F��*�E*�$��ߝ������c���	!���;��Y��uu��ɇ�T���E���ǳ�Oɿ��߿ܠ�ֻ���z�(	׿������M�t���P�e�C�w�N�#�p��8���#����Կ�����������㿲uͿ��������y]���ߊ��,|�k`�8�C�9�(��u���`]������B50�"=L��vi� ����S��`��#������2`Կ�)꿿���������J�пɯ����io��hR��HM�"`�����t����ÿ(W�<���������HG�<dɿ���������	����yy� �\�i@��q&���������=Z�Ǽ#��<�	AY�]�u��K��Ɣ���G���jƿ�?ݿ;^� ��� �����\�ƿR�� ���?�b�}xM�	.P�k�j�o���v��h�Ϳ/�J�����h���\ؿ�����Z��`���A��𯅿�3p�yWS�$V7�?��q������
�5C��:,�K�F�Z�c����4����x��%h��S�}ο�'�=�������m��ܿ���u�ء~�M^Z�<M��W��y������m��ٿ���  �  +���$�
������:�˿�/��5���N�c���A�n�%�	������}վ��¾鮽�e"ƾ��۾)B������+��I���l�ύ��M���ֿ�p����'��*�r� ��3���俆h������=p��&h��xޠ�J�Ϳ�����(�O�*�� ����E��/���1A��H�X���8�D����v,꾈�Ͼ9&���Q��<;�V���?��G5�,T���z��9���Ź�o忴
�g|�!�)�|�(������ӿ8ͤ��%����h��	m�w\��r���l߿��	�^��|+�Kb)������0�ܿ�$��ѣ��#
u�BjP���2�������cT�c-Ҿ��Ⱦ�C;P߾b���x���)�x�E���f�kɈ��T���˿�����l�Tu%�^-�g'�K��^��Y�ƿ�����O�� �n���~�����<¿�������B�&��-��'����n��2eѿ�����'��5�n�E�L�x�0���Z_�����ھs"־�߾����#�U ��b9�ŸV�3�z�h���<��	�ܿ����+�`o.�x�$�c �J��`����ꕿ�u���2y�����[}��ޘֿCW�F�<b,��/���$����*���ƿ@��'�����h�1I���.����^C����~e�#��nU��N��=��v+�^�E���d�h����z���¿	x�M���"��7.��-�q����\�ۿFL��0���x�y��}�����������N���%#���.��,�����9	�`n�9ƹ��H���&����]���?�L�&��h�^� ��}�����T���	���@�4�� P�Sq�Rw���8п#�����o(���/���)�ZX��
���˿M������Ox�b�����KwƿhU�����>�(��  �  9e�<�[���A�����3��.X���܋�F�W��K+�L��ٞ�bdƾ'���ѡ������l���J���;w\�0��Q4���d�������ſP���J'��	I�B�_�Fe�d�W�7g:�Ѝ�^�a��� ��2��������ɿ�1��v*�[4L���a�ױd�HU��77����࿔��so��m?H�	� �����ݾ
��h��Y����
��U���If`پ�� �Ą��B���x��w���ٿ1���3��R��c���b��O�vH.�[��V�Ͽ�3��O��H���jƩ�lݿ+��Y�6�F�U��Te�?b�'M��/,�|���ο�i���n��<��`�^���(ھ�U��ڜ��{ާ�eK���ȸ�F)о��񾞬���.���Y�����}d��3��1���Z@��[�P^g�0�_�5IG��$�i����¿~������� ޘ�v̼�$U��[( ��0D���^��3h��^�
�D���!�����ɾ��K��c�b�aH6�I���6���fݾ�ƾ����I;����s�̾��gy�;��B��cr�i⛿+�̿�d�d�*��}L�dOc�8�h�sL[�@>����N�쿤3���7��h���քҿ\�	���.�u�P���e���h��TY��t;��9�<C鿕Z��e����X���0��B��<��e߾T�ʾc쿾/G��l�Ⱦ�6ܾ¸��q7�>�,�D�R�W���{���k������Q7��LV��g���f�RS��2��:��'ؿ��������z_�����j���y���:�<Y���h�D~e��gP��|/��
�¯Կ#���|���I��l&�����]�I*ؾ��ƾo���ސ¾c�Ͼ�d�X��vU�%9���c��������0����h���B�tC^�D�i���b���I��x&����-�ƿ�>��Zl��Z����c�������["��SF�ӧ`��  �  ڼ�������o���A�G[��+ӿi���C�Z��#�i���u�̾����d������Sv������$����M��˔־X/��M.�0�j�⎢�������4�L�X�x�Y�����������f�X`7�7�	��0Ϳ/֥�E���B���ͭ�@9"�"BR�cX}��3���,���'���a��2��� +��؂����F�ʣ��*�����d������t����v���H��g���n��e���?��q��۵�}H����,�Fe\��D��	����������8W�p&'��E�������j��:��-�ƿw���2���a���������m��R�}�vS��"��:���Y�v���7����e�����E��_��3���!��J𠾽�����վ^��3�%�M�Z�r��X@Ͽ)R��>�	m�l(��m�������͝v�KwI�����W�3e�����寿n޿�7�)]D�r�5�������r�?�D���7�ؿ���Wte�z�.��	
�CG�F�¾�ݭ���������嶥��#��_o̾N3񾳴���;��sx�|��M��	8 ��RP�,J|��Ќ��]��Yȇ���j��l;����
�տw���f���u��c����&�ƗV� Հ�}Z���P��ZI����e�M6��.��|ſ�Ǐ�L!W���&���Gk��vž�^���^��eө�Y�����¾�޾Ҧ�WK"��1P��������"K���0�[�`�a�����"��������[��q+��n ��Ŀ{���ی��AYϿ�	�$6�e�e�nS���A����O����RV��*&�����o,������D�<��X���l�׾���}Y��uZ������������˾?��f��w0�2e�J'���aԿ3���A���o�t��h��B��(y���K��`�"꿨���E��������;�F��t�&���  �  ��h�������H\�He$��S迲Π��a��S"����n��M���~��7+}�`w�np��7o������ɾ���p.�Ȫs�5ɮ����m�0���h�����������\���CW���O����Q� +���Ӭ�*ʿu�d7��o�Gc��5����G���Ԗ�����O�I��a�,ο ����J�������[_�����}��Tu|�f{{�����M甾d����ھ���?^B���;�ſ&��'C�j{�y���@����Ġ�������t�*=���
�Q1Ͽ+���:걿��ۿp>���I�~���G������=��Ѽ���o��7����෿ڃ��1�8��	�Uc׾-�|��0���
Ȇ�]����)���$����Ⱦ���� 6$�o8`�6:��B��w �|�W���9M���أ��m��Tc��l�d�<z-�����)`Ŀ${��];������>�'���^�S����?��C���B��9���_��'�c��9>���l�R-�_��Y־�����������6��\���O������	V�9�2 <�<���(����~�{4�kl�����h���Y���J���lN��{T�������ܽ�o���K�ҿ��
���;�"ss�M�������k��
���_�����M�
���}ֿ�<��g�Z��($�����Ծk��2Ȧ��{������8���0��\о�I�����L�R��O��2�Ϳ!��7TG��8�˖�j���<������,y�^wA� @��׿�I��Sy���q�d���M�q������{S��K��yg��Gs���:��O�s����"��'�E����� ��Dʾ�鱾���|�������r۪��Q���6޾#�ۮ.��j��]����9#��Z��O�����O!��@�������~g�r�/����jɿ�-���Ŀwr���(*�Z�`����M���  �  }?��<yu��eW�.�)��:�������S<�(���;���f���fh�Z2V��bQ��VY�ro�;��^Z��t۾���CpK�@����u˿�~�.�7���_���y�,���np���N�û$��2��*W��鉗��;��xd���ٿ����<��\c��{�͏�>�m�!�J�����=�l0��im�o�)������������Z���c�h*V�yVU�da��|�3Ҕ�w ������Y#�P�c�i{��o�@����E��'j�X~��}���f��"A�MM��f�����ؑ����ܴ��!� ���J���m����Ԅ|�z-d���=����տNB����V���:��U��*떾�ꂾԬo��g�!Yl��Q~������_����վ��t=�z��h���� �/)+�*U���t�M1����y��|]��5�|�
��п����.5��s䠿�
ʿ�����0���Y��x�r���/x� Z�1�0���-���_$���@G�-������-���e���������.��"���a�����N�ľu����y ��*Y�����7Zҿ���\Z;��
c��{}�d���$t�9�R�Q�(�: �+�¿]��qә����U�;?��A�3�g�m��8���q���N�{�#�L����x����}��':����+߾S踾i����0��A���ӊ�!ݐ�u8������Yپ9��ƥ3��Xt�ʵ������`J��[n��H������H�j�ofE�ɒ���迈���]Z��r���0��>I���	$�3�N���q��́�����}g���@�[d���ۿٝ��&d�i)����=�о&���������M`��&ԕ��'�����8*����YG�����! ����	�-��W�{�w�yy��U|���_��7�?���Կf���Z옿K���:�ο	����2�;�[��*z��  �  Hhu�o�j��2N�s�&�qb��gi�����:�5��3�Ͼˤ�ވ��/o�~�\�C�W�0�_���u�%w��l����ܾPl��H��>����Ŀ���H0��V��/o�i u�$f��JF�e��}^��{N���O��+`���%ҿ�E���4�r�Y�_q���t�
Uc��"B�j_���㿶u��:�h�%l(�ho���Z���盾�Ѓ���j���\��[��h��y��#6��\ǻ���[A"�	�_�C��3�ۿ����=�~`�pWs��/r���\�]9�g�(zؿy西|㍿����u-��Hr翢���[B���c�u�m�q�skZ�Ͱ5��z�y
οu}���S�mJ�H��iQ���[���Z���Ev�+n��r�����Zu�����D@ؾ���E;��ɀ�Џ�������D$��*L�uj�lKw��$o�3/T�R�-�$���=ɿ*S���V��h���~ÿǧ�-r)���P�a�m��x�b�m��P�I�)��� ��ۻ��4���E������dd��(ޟ����O��9b������*���5�����Ǿ���J ��KV�"��׼˿p�
�A�3�uY�Ҭr���x�Y�i�2%J��"��N���ż�<қ��㕿������ڿr��/59���]�?Gu�T�x���g�'YF���l7�*���py�~�8����G�ᾃC��;��6���}{��F��M1��p���Zy��� ܾI	��2�FTp��P�����A����A�jEd�A�w��lv�Pa�l_=����/�%o���`��}d��j{���￢���%F�Ojg��x��u� �]�r�8����A�Կ����`�ra(�$����Ӿ"������jg��/��������4�����CTľ�����rE��셿^�������c�&�7�N��	m���y�N�q���V�[+0����οJ��*��T���"ȿ��� �+�:�R�֟o��  �  �&W���M�{S5����/�⿅M����t�Ƌ5�V�	�e�ؾt꯾�S���x��R(q���k�֗t�� ��:���<����;���/B��{��B������m��~<�`�Q�L�V�$J�ߝ.�j!��;ֿ����ɑ���e��w����������.��WU?��mS�=hV��G�H
+��R�s�Ϳ�M��?H^��/&�i����,˾�N���"��{����p�i�o��*}�����s���q�žs����� ��pV��֑�8�ƿ};��'���D�OZU�shT�2B�)C#��\ ���¿���6₿֐��q���H�Ͽk��N+�hH��W�I T���?�=� ����룻�)���!eL�k������ľbݥ�cy������U�������N���۞��ٹ�CV�a�=X7��[t�[x���1߿����3���M��
Y��R���:�G�����l���x��[���+���㒱��0�,���7�2�P��Y��P��8�Ά�#���������>z@�
��k��#�ƾ�S���왾���]���J��P���� ����Ҿ�v���N ���O��^���w�����|8�+�?�U@U�"�Z��M��q2����f޿�T��z�������ƿp'���#��C���W��Z� �K��@/�����5ֿN���E�n�\�6������0�Ǿ�g���+��$����������$מּ(�þ?�+7�1���f�����Ͽd�N+���H���Y���X��BF���'���aa˿
��JT��f�ϧ���׿.S�/�P�K�)�Z��]W��GC��#��� �48¿����)�Y��(��R��޾<��3=���Н�IØ�˚�� ����a�Ͼp�����q�A��~�U����T促f�}r6��P�}�[���T�T=�[:�}��[6���6��vF��%����/��˹�9c��:���R��  �  ��-�պ&����W���M���蔿0�e�a)4�w���w�Ǿ���\������^ڇ�,��[��������9Ͼ\\�����xJ>���s��8���̿�� �8��)� �-�N�#�7�+�,�������m��`e�����X꠿G�Ͽڪ�~3���*�>-���!�p,�:�]������jT�W	(�f�&T�4d��ʤ�z���,���S	��D����)�������Wܾ�����#�2N�K���#���M�ݿ�(	���(b,���+��;�vb��Կ���vJ��Xf�Vmj�6���V1��i��8��z'"���-�^�+��C�Jj�3Կ����j]~�� G��~����E�۾���|r������~���T�M���崾��оd������7�\�f�y���˿����A�$'�ƣ/�D&*���+����ǿ]E���2���l���|�����3�¿.�������J)��l0��v)�ʦ�ŕ����ƿ"]��ǖp�?�T�������ݾf����-��?��pI��l���5����ʾذ�0�	�ߐ%�KL���� ���ӿ��k���&-��(1�#0'�����q$���O��'Q~��Tv�=���8z���ؿ����z�3/��~1��&�3c��e쿣V���?����d��k8�,d�� ��޾ež�³������0��*"��o\¾f�ھ����q��y�3�`�^����*۴���`V���#���0���/�-y!�A�	�gRݿ�{��Һ����v�Z�z�\ё�&���<�:|��%�H1���.�f�������ڿ�M��JŅ�MIT�ѕ,�m���i���վ�3��dа�T����-�����
 ˾��S��}vA�Fq������ĿpD�������)��92�C�,����� ���̿y����P~u� 򂿧.���vǿ������\+��  �  �$�T����A��zĿ(=��N����r`�U�=�ϣ"�s������Ͼ[��XЧ��w���s�������־1D�������(�/fE���i��͌����	q̿ ��� �M�<m���]ٿ볿_Ph��G�D�A���V�P��wZ���/ɿЭ�g� �U�����sۿ����¡���(~��U��D5��������8aȾ�u������r륾3q���1že�⾣l�����1�]�P�kx����6����f׿����t��u��k�<�̿��)����Y�_IB���E��gc�â��e@��`=ֿr���aa�WM�[����ѿ������Ur���L��t/�Bx�A
�'��"cȾ1<������[�������پ�������0'��B��c�ɻ��թ���Ŀ������n!�� �O�ndĿ��P����W���H�0U�+{�
ϛ����!��m� ����m��3��V�ɿ(���4���Yk���H�	�-�b����������ξ����ܻ�jXþ�վ����	�^��D6��S��w���������FOӿ���G�<��������࿄���(痿�ex��PX��R��g��Ԋ�_嫿��ѿu9��"B��P�L �g��\¿���>]��ۄe�&�E��+��)����פ�g�Ҿ��ƾ�ƾ6�о\c�e�ŗ�?�(��B���`��n��=K���⽿��߿����������m���zWտ\t��
���S�j���R���U��ys�Pz��&ܷ���ݿ������ݦ��u����ؿ�����8��׃���Y���<�^n$���B�����.ξyiƾI�ɾR�׾���f���6���1�y~L��n�aߌ�[Ш���ɿ���Fc�X��ބ�6`�*`ɿk��儿�#a��7R�=^�����?���Fſ��鿀���  �  ���R��v���GԠ��� k��N�p��\\��G��H1��2�'��澃�оiFʾ�VԾp��c	������6���L��Oa�m�u���������\िF��8H��"���CԳ��ǟ��-��5�^�A9���"�ѭ��-�gL���x�^/��=��V��k����ܹ��F��$�����������j��V��`A�D�*���_D���;߾E-ξ�3;�jܾ��������'� �>���S�
h���|��Ԋ��ș���T2��V����w����{��t+}�/P��G/���?q!�6�r�Z�[�����*��j��6p���o��Nu��(0��z�����{�7Hg�iS�"[=��y&�JR��������:�վҟھG�ﾊ��L_�δ5��}L�іa���u�����2��~墿V���V��{Jÿ�1���ܪ�[C��Fhu��K��?0�{&��.��H�^�q��X������d����Ŀv����>���T���m���߈�2k{�JKg�\�R�	o<���%�*������y辒�⾏%�p�pI�{�,��D��`Z�8o�;��f��ȍ��=���*���;ſ�ſ���9���֎��en��I�M73� R/�k�=�4V]�Ǆ�����_x����ÿUzȿ�S¿����~W��0��zT��YF{��g�߭Q�A�:�Z�#��C��n��hV�LY������L!�S�7�L�N��:d�Pfx�W���?�����Hq��|����ǿ0aĿ����蟿(�����`�.�?�*�/�R�1���E��j�����\��W3���?ƿw ǿ�	����*��U��}���ot�3 `��KJ��=3�n��d�	�(��NP�2��1�	�R)��n@�?W���k�l��2���Y������2���Ŀ�|ȿ1Y���󯿊E���@�g�U�7�9�Ow/�`�7���Q�nPz����u���r���  �  mߌ�N�� l������D���Q����P������6���m�h�M���-����K����t�����4�A+U��lt������"��ܐ�����+�,�����{\�� �x���i���H�k�)�4�8I�����!	������:��.[�ʲy������&��7����!��Y����>���"���犿����X,d���C��F%�������[ ����"��?��Y`��}�^ʉ�l��������G������A��А��"�������{�q�]��=�r& �]�
���������i�A�'��F���g��V��U����������X�������]��SĒ�C���ϭ���{��+]�B�<�>� �!��	3��������1�U�P�mq��b��뱏�^퓿{r������-��2?���_��w������^z��![��7;�) ���)=�����m�u=9��YY�,dy�T承8W���ϕ���&���,��>���*Õ�$������'�x�i�X�}9�V���9�J�
��o�+�%��A��;b�7݀�1b��R���(���[����Ӗ����ߗ��O��I ��!���N�w�e�W�#P9�*� �����o���.�a�K��*l��Z��+��΢�� ����-��0����ژ�����^��/�������ft�S�S�Pg5��
��(�4n�$���32���O��p���-����*-������	������.��ц��x��NV��7�n�==N�ܿ0����$��������6�@�U�av�S��od��C]��(R��$���MD��j󘿨Z������3���N����i��I�"-�d��������"�VC<�3�[�D�{�����政���閙�kϘ�L����r����������:莿�I���/e��E���)��f�����-['���A�N�a��Հ�)��  �  �8]�:~q�����Ñ��á�U���ּ����Q���=����� oe�6�=���$��n�	�(���E��o���?��E1�� ���eD��f����s���ݎ��Ɓ�h�m�<�Y�ƹD��.�a���[0㾖�Ͼ~̾��ؾ�F��y���$�1;�2�P�[-e�R�y�h숿����ӧ�h����J���ͽ�X/��'����#���W��M4�F� �����61���R��H��H,��Z ������k��&���]K���瘿����x{�ԍf��WR��<�G�%�M�^@��g�ھ�̾�CϾj�ᾬ&�7D�f�-�2�D�ZZ�Żn�3,�����:k��d���f�������u��@���^�����y���N�Qi0�,=#��(��@���f�h���(��)񷿰K¿�d�����i|��DZ��!Y��l�{��jg���R�(=�S&��>��\��q�<�۾$�������s��r%�M�<��XS�z-h��|�ُ���C���<���
��<H¿�Ŀ!���lר�S���U q��jI�Ғ0�L�)��5��R��|��9��Zڮ��迿�ƿC ¿���U��[���f�����{���g�rS���<��"&�,v�Y�|�ﾩ��z�����
�/W���4�L���a�[v��`���V���៿�'����ǿ��ſ�T������9�� �g��eD��1�y�/�BIA�qc��W��H@�����Ŀ�ǿ�쿿���z2��UW��&��IMw��c�J�M�В6������X��$����_ �k:�~�$���;�h�R���g�}|��ƈ���������\J����¿�5ȿ�¿Q��~���6���Z�\~<�Z%/�,^4�y�K�Hr�*������@��[�ǿ�ƿ[(�����ކ������>����q�~U]��:G��!0�%�O���v���p�����X�;��-��E�pg[��  �  �i?�]ub�t	�������eƿ������+�#���y�޿��=,���:o���J��8@�ƲP���z����͓¿�E��'��0D�����࿆&��@n���܂���Z��9��D�5		����8z̾������t��=�F4��^`ݾeb ��4�	�-��bK��q�B����e���Jҿo����_���w�I�ӿ��������a���D��nC���\�
2���s���PϿ{Q���Y��_�#�տ����a��F�u�mUN�5�/��������߾xJþ�h����`֧���9̾Q�����]7�n9���Y��ၿfӜ�u)����޿�p���	��x����fɿ�m����fY�	.F���M�Q�o�����V�]޿������� �O�dο�n��qݎ�v�n���J��.�:F��W�Q=��e˾Nݺ�E�������˾z���J��K�S�.��aJ��|m�Ӎ���y����˿�j쿾���K& ��j�ƨ������� {�ϘV�WGL���\�둃�S��<�ȿ���������� �`�\ƿ�O��!É���h���G�:�-���s���	�b\Ծ�tǾ�ža�ξ�p�1���=��&�<�>��M\��;�����'ĸ�e�ڿ&�����a���k�ۿ�ε������3q��	U��S���l�=��+���d׿nk�����n�����c�ݿh��K���O/��4_���@��'����� �k侽�Ͼ��ž�Ǿ�Ӿ��龑_��#��-�:�F��4g�9{���d��,�ÿ~a��~ �SL�5��Q=�jXϿ����/��@se�2R�	�Y��u{��7���d��� ��v�n��2�G:ӿC�������>y��@U�K�8��!�@n����,�޾P�;`�Ǿ��̾r�ܾ.������}�,�6��  �  @?6���h�����Ŀ��5�^�'�j�-�J�%�R&��ￆ����#����q��c�Bz�R%����ƿA
���l�6�(�S�-��{$��%���쿧���~ݎ�C�\�u.��g��羃þ������(A��h���������>���n־� �����F��~�Y����տJ�*���c+�#�,�ó ��
�g7޿q���s1��$�i���g�	��ŧ��0ؿX���:&,��#,���������ڿ���佂�z!K��(!�7���xپ̀�������Z��A\��:�����u���Kþz�羡����,��-Z��w��5"����迾[���#�DW.�p5+�[���0�g�οy���|
���i�t�Od���Z�������&�5k/��*����.� ��wͿ!x���Ww��	C���3g��ܾ4$���I�����܂��j֝�����{���ݾ?J����9A�%�s�ƒ��d�ɿ������U=*���0�S�(�2��͋���n����¾}���o�����F��q�̿50�¨��@,�U1���'�q���v�ry����b�j�#<�L��{[�$��kƾu����檾����t��������׾��������.�VmW�Eه�L���O�ݿ;@	�� ���/�K1���$�z�)L�ᵴ�=����y�Y�w��'���ϯ��>�����"��60��80���"����1��^�������[���1�5������{bپ�G��g~��	���1����l��lƾ�8�������B:�q~g���������5����&�"�1�ri.��!�M���Կ�����×u�����:�������������(��2�[-�^1�%~���ҿ����6ဿpM�!�'���������Ҿ�������N���꯾(���о���Tv
��$��  �  8;8�i y�t+���%�|���7�� O�Z1W��1M���3�W��D࿑���F`���R�������޴��^�и�q�:��Q�jW�� K��Q0�<��ؿ&,��dli�b�-�2��[ҾG૾j��~���3�q�t�n���y�Arg��ꩿ�����e�L�Ἂ��D���I��ܬ!�V�@���S�<V�gF��1)��_�5�̿꽝�(%���Ճ��ә�SXƿ}��_%���C�
U���T�-mC�6O%�%Q��hÿ&=���R������þ����_���Jr|���p���s������ؒ��N����Ѿ����i+���d�mu����ҿ��Ů-���I�\�W�r�S���>� ���1��I�bF��!{����-ɨ��;ܿ{�1�1���L���X��R��6<����vs����΄�~GF�������_�žƘ����������>����G��5��o&��%�ž�ﾐ��#7C������p�����9��Q��Y��O��6�r���������V���P��%���[�Ԇ������=��LT�dZ�`N�L�3�����޿P���Lw���;�� ����|ɾ�P��)��Tl�� u��=���^ા���O+��>�E�*�c]�F)��G�ſ���e�%���D�RX�4Z��xJ�T?-�3j
�i�ԿUɥ�8.���݋��ܡ��bο���h)�E�G�*,Y�yY���G��m)�t�Z�˿����	Ic�|�.�Ȕ
�侢m¾�����5���Ø�����M[��ɾ�������8�Z3r�b
��1mٿYW��0���L���Z�b�V���A�P�!��G����¿gC��p��;���4��R���4�zO�Dp[��BU���>�T.�W���xC�����]�P�,>"����$�پKm������������S���ǧ��C����־2 �=���  �  ==��$���͹�9X �d;)�E.P�5l��pu�O�i�8FL���$�����g$���������r���)ȿ�����-� T��@n��Iu�_^g�dSH�8- �b��¬��u�\"1�g����Ⱦ����8����m�#�]���Z�@
e�]�}��蓾F)�����̋��eT�:���G@п����+7��h[�c�q�`!t�f�a�F�?�}c�D��B��~|��t���$����}ܿ���a�;�ԭ^���r��r� �^�u;��R�9�׿4��&�[�/�����ϸ�!D���h���g��]��_���o�ڕ�����-Ⱦ���r.� 4p�/�����'}��E�^�e���u�&q���X���3�}7�:#ѿ�ڢ��W��S䖿o�������!�"�I��i�w�v���o�0�U�P�/�ƪ�7�Ŀ�/��z1L��^��辶Һ����⯊�����*6{�����N��6���[亾
y�R{��9H�詉�2T������+���R�!�n��1x���l��O���'��A ��¿�������o���")ο��i1�^KW��}q�^�x���j�
�K�%�#�`���f���F쁿�(?��&�U��W$���פ�٧���/���Y��0������L��Z�־D���e+�>Be�b���ؿ"��S;�ӊ_���u��7x���e��D��m�P�뿌��o���q ��������w��j�?��b�a
w�Q�v�+�b��?�]u���߿X_��k>l���/��z���پ������������卾a������9���������H�;�;��}}�*������GVH���h�7�x�IMt� \�_�6�	>�$׿�Ԩ��L���Ӝ��i��ko��=�$�ŠL�+�k�(�y���r�O|X��V2�1B	�X�ɿ�d����V�y�!��/��� Ͼ����񧓾�������ܜ�Jʮ�R�˾9����|��  �  Z�?��5���п�SZ��~0��zY���v�SC��$Lt�xFU���+��2�ϋ¿#	������\g���(Ͽ�
�o5�y�]�F�x�,/��%�q�77Q���&�>������{�f�2�%���Cƾ�K���2����f�VW��YT��m^� �v�U{���9���}��J��W�����~׿���V)?�(Ae���|�/ ��k�qVH�K��PT쿒���쑔����^ݭ�������r�C�ܘh�]�}���}���h���C�WT��C߿�J��Tj_��* �-�� ��㒾*�y�sa���V��`Y��:i�.%������[xžo3�?�/���t�������� #���M�"�o�m��9�{�u�b�%k;����U�ؿǧ�?���-������p���y�(�%�R�(cs����G�z�Fc_��C7�����/˿����2�N�������ݷ��?���5F���z���t�X�{��釾<��a����[� ����J���� Wſ��A=3��6\��ky�����w� X���.��#�#{ȿo�������(f��y0տ�	�|�8�+�`�/|��ԁ��&u���T��W*�E����帿�|����@����:�"պ�xY���B��Wꊾt��£���-�������Ӿ��e#,�9�h��	���߿>���QC�Bci�B`��J���
p��cL�b�!�Nc��в��Қ�����嵿$�쿟��l�G�٤l�����������l���G��v����)���Fp�Y�0����|�־�����J��|^�������l��X�������1g����ᾒ��`�<�C���������?&��Q��(s����[���e��x>����؆޿�����3�������ſLb�2_+�7lU��v�A[��Q}���a�[�9�<���bп�����HY��"��B����˾:y��l���a��茾�Ϗ��u���R��{bȾ�������  �  ==��$���͹�9X �d;)�E.P�5l��pu�O�i�8FL���$�����g$���������r���)ȿ�����-� T��@n��Iu�_^g�dSH�8- �b��¬��u�\"1�g����Ⱦ����8����m�#�]���Z�@
e�]�}��蓾F)�����̋��eT�:���G@п����+7��h[�c�q�`!t�f�a�F�?�}c�D��C��|��t���%����}ܿ���b�;�֭^���r��r��^�u;��R�?�׿9��-�[�"/�����ϸ��C��vh��@�g��]���_���o�������[	Ⱦ���/.��2p�b��̇鿱|�E��e�v�u��%q��X�\�3�L7��"ѿ�ڢ��W��g䖿����j���L�!�o�I� 	i���v�'�o���U���/�;���Ŀ�0���2L��_����>Ժ�����������:6{����DN������⺾%w�*z�I8H�!���US���+�+�|�R���n�r1x�9�l��O�b�'�pA �k¿�����������c)ο3���1��KW�P~q�חx�+�j���K���#�S���G���큿*?�)(�g��&��٤������0��ZZ������䥟������־W���e+�FBe�d���ؿ"��S;�ӊ_���u��7x���e��D��m�P�뿌��o���q ��������w��j�?��b�a
w�Q�v�+�b��?�]u���߿X_��k>l���/��z���پ������������卾a������9���������H�;�;��}}�*������GVH���h�7�x�IMt� \�_�6�	>�$׿�Ԩ��L���Ӝ��i��ko��=�$�ŠL�+�k�(�y���r�O|X��V2�1B	�X�ɿ�d����V�y�!��/��� Ͼ����񧓾�������ܜ�Jʮ�R�˾9����|��  �  8;8�i y�t+���%�|���7�� O�Z1W��1M���3�W��D࿑���F`���R�������޴��^�и�q�:��Q�jW�� K��Q0�<��ؿ&,��dli�b�-�2��[ҾG૾j��~���3�q�t�n���y�Arg��ꩿ�����e�L�Ἂ��D���I��ܬ!�V�@���S�<V�gF��1)��_�6�̿뽝�)%���Ճ��ә�UXƿ}��_%� �C�U���T�2mC�<O%�+Q��hÿ0=����R�!�����þ���������p|���p���s�%���t֒�	L���Ѿ���[g+�(�d��s����ҿ��߭-��I���W���S���>�����0����F��{��5���ɨ�|<ܿt{���1�n�L���X���R��7<�l��6u�Y��YЄ�JF�������Z�ž ��� �������M����F���3��O$��?�žR��R���4C����v������~���9���Q�?�Y�W�O�V�6����?��O����U���P��c����󺿐�������=��MT��dZ�aN�D�3������޿���Ow�k�;�9#��	�-�ɾpS��Z���n��Vv��A���!᪾�����+�?�]�*�c]�J)��I�ſ���e�%���D�RX�4Z��xJ�T?-�3j
�i�ԿUɥ�8.���݋��ܡ��bο���h)�E�G�*,Y�yY���G��m)�t�Z�˿����	Ic�|�.�Ȕ
�侢m¾�����5���Ø�����M[��ɾ�������8�Z3r�b
��1mٿYW��0���L���Z�b�V���A�P�!��G����¿gC��p��;���4��R���4�zO�Dp[��BU���>�T.�W���xC�����]�P�,>"����$�پKm������������S���ǧ��C����־2 �=���  �  @?6���h�����Ŀ��5�^�'�j�-�J�%�R&��ￆ����#����q��c�Bz�R%����ƿA
���l�6�(�S�-��{$��%���쿧���~ݎ�C�\�u.��g��羃þ������(A��h���������>���n־� �����F��~�Y����տJ�*���c+�#�,�ó ��
�g7޿r���t1��&�i���g���"ŧ��0ؿ[���?&,��#,���������ڿ���򽂿�!K��(!�0��bxپa���ܸ���Y���Z��CK
���r���Gþr�羢��5�,��)Z�qu����� �迃Z�z�#�'V.�s4+����0�k�ο����
���i��t��d��}[��J�쿥��&�Il/�O�*�̞�o� �AzͿmz��/\w�XC�:���i�c�ܾd'���K��4���򂙾{՝�艪�
x��[�ܾ�G�����5A���s�p����ɿ ������<*���0�T�(�_�������m��x
��/�}���o�	���G��q�̿�0�����A,��1���'�ő�<y��{��ŕ���j��&<����Y^�����nƾ����K骾����㽰�����׾h��ʩ��.�jmW�Jه�O���P�ݿ:@	�� ���/�K1���$�z�)L�ᵴ�=����y�Y�w��'���ϯ��>�����"��60��80���"����1��^�������[���1�5������{bپ�G��g~��	���1����l��lƾ�8�������B:�q~g���������5����&�"�1�ri.��!�M���Կ�����×u�����:�������������(��2�[-�^1�%~���ҿ����6ဿpM�!�'���������Ҿ�������N���꯾(���о���Tv
��$��  �  �i?�]ub�t	�������eƿ������+�#���y�޿��=,���:o���J��8@�ƲP���z����͓¿�E��'��0D�����࿆&��@n���܂���Z��9��D�5		����8z̾������t��=�F4��^`ݾeb ��4�	�-��bK��q�C����e���Jҿo����_���w�J�ӿ��������a���D��nC���\�2���s���PϿ�Q���Y��_�6�տ����%a��i�u��UN�A�/��������߾�Iþ�g����ӧ��%̾6�뾣���3��i9��Y�߁��М��&����޿�m�����w�����ɿll���񂿡eY��-F�*�M���o������︿�_޿������y!�B�eο�q��@�����n�h�J��.��I��Z�JA徦h˾�޺�a��x���˾���<H��H�Y�.�$]J�Rwm������v����˿�g�I����#% ��h�C���{�����z�!�V�cGL���\������T����ȿ����V��M� �0c翆	ƿ�R��Ɖ�W�h���G�k�-�w��j��s�:`Ծ�wǾ7�ž �ξ	r� ���U=�2&�a�>��M\��;�����'ĸ�e�ڿ%�����a���k�ۿ�ε������3q��	U��S���l�=��+���d׿nk�����n�����c�ݿh��K���O/��4_���@��'����� �k侽�Ͼ��ž�Ǿ�Ӿ��龑_��#��-�:�F��4g�9{���d��,�ÿ~a��~ �SL�5��Q=�jXϿ����/��@se�2R�	�Y��u{��7���d��� ��v�n��2�G:ӿC�������>y��@U�K�8��!�@n����,�޾P�;`�Ǿ��̾r�ܾ.������}�,�6��  �  �8]�:~q�����Ñ��á�U���ּ����Q���=����� oe�6�=���$��n�	�(���E��o���?��E1�� ���eD��f����s���ݎ��Ɓ�h�m�<�Y�ƹD��.�a���[0㾖�Ͼ~̾��ؾ�F��y���$�1;�2�P�[-e�R�y�i숿����ӧ�h����J���ͽ�X/��(����#���W��M4�I� �����61���R��H��O,��c ������k��9���sK���瘿����x{��f��WR��<�'�%��L�v?���ھ�̾�@Ͼ���`$�TA�ۢ-���D�,UZ�K�n�7)�����h��7���`�������s��1�������Z�y��N�bh0��<#�y�(�-@�ճf�߄��*��w�^N¿�g���������]��E\��D�{�-pg�aS��=�]&��@�`���r�]�۾ҝ�%���`q��o%���<�TS�5(h��}|�����P@��e9��F��E¿@}Ŀ����aը�������p�kiI��0�Y�)��5�aR���|�9;��~ܮ�D뿿؍ƿ}#¿����\Y���Õ�����Ź{�2�g�9S��<�F&&��x�7[����<��h�����
��W��4�ZL�$�a�pv��`���V���៿�'����ǿ��ſ�T������9�� �g��eD��1�y�/�BIA�qc��W��H@�����Ŀ�ǿ�쿿���z2��UW��&��IMw��c�J�M�В6������X��$����_ �k:�~�$���;�h�R���g�}|��ƈ���������\J����¿�5ȿ�¿Q��~���6���Z�\~<�Z%/�,^4�y�K�Hr�*������@��[�ǿ�ƿ[(�����ކ������>����q�~U]��:G��!0�%�O���v���p�����X�;��-��E�pg[��  �  mߌ�N�� l������D���Q����P������6���m�h�M���-����K����t�����4�A+U��lt������"��ܐ�����+�,�����{\�� �x���i���H�k�)�4�8I�����!	������:��.[�ʲy������&��7����!��Y����>���"���犿����Y,d���C��F%������ \ ����"�!�?��Y`�.�}�jʉ�|��������G������A��А��"�������{�S�]���=��% ���
�����F���g�؞'�ӳF��g��T������4���l��� ��4����Z��H���}���a���̲{�d(]���<��� �0���2�p�����1�A�P�0q�.e������\𓿵u��ޫ������|B���b���y�������bz�)%[�6:;�� ����:=�7��l�&;9��VY�(`y��㉿jT���̕��앿S#��y)������	���0!��1����x�4�X��z9�͕��8�W�
�Xp�ӭ%���A�J?b�X߀��d��@���e���Џ���ז�����◿�R��1��������w��X�S9�o� �C��c�l����.��K�J+l��Z��<��ע��$����-��/����ژ�����^��/�������ft�S�S�Pg5��
��(�4n�%���32���O��p���-����*-������	������.��ц��x��NV��7�n�==N�ܿ0����$��������6�@�U�av�S��od��C]��(R��$���MD��j󘿨Z������3���N����i��I�"-�d��������"�VC<�3�[�D�{�����政���閙�kϘ�L����r����������:莿�I���/e��E���)��f�����-['���A�N�a��Հ�)��  �  ���R��v���GԠ��� k��N�p��\\��G��H1��2�'��澃�оiFʾ�VԾp��c	������6���L��Oa�m�u���������\िF��8H��"���CԳ��ǟ��-��5�^�A9���"�ѭ��-�gL���x�^/��=��V��k����ܹ��F��$�����������j��V� aA�E�*���cD���;߾L-ξ�3;�jܾ�������#�'�2�>���S�6
h���|�Պ��ș�.��j2���V�����x����{��6+}��P�,G/����o!�@6��Z����@���(���g��Tm���l��r���,��e�����{� Cg��S�MW=�}v&��O�m������݅վݠھ��ﾄ��
b�S�5�E�L�՛a���u���5���袿���Y��IMÿ4��ߪ��D���ju���K��@0��&�]�.���H��q��V��~������/�Ŀ[���f;��1Q��\j���܈�Ie{� Fg�ʥR�>k<���%��'������x辫��%'�q��K���,�zD��eZ��o�LŁ��i��;����ë�v-���>ſ�ſ"��>;���؎��hn��!I� 93�gS/�\�=��V]�ZǄ�����xx����ÿ[zȿ�S¿����|W��.��yT��XF{��g�߭Q�A�:�Z�#��C��n��hV�LY������L!�S�7�L�N��:d�Pfx�W���?�����Hq��|����ǿ0aĿ����蟿(�����`�.�?�*�/�R�1���E��j�����\��W3���?ƿw ǿ�	����*��U��}���ot�3 `��KJ��=3�n��d�	�(��NP�2��1�	�R)��n@�?W���k�l��2���Y������2���Ŀ�|ȿ1Y���󯿊E���@�g�U�7�9�Ow/�`�7���Q�nPz����u���r���  �  �$�T����A��zĿ(=��N����r`�U�=�ϣ"�s������Ͼ[��XЧ��w���s�������־1D�������(�/fE���i��͌����	q̿ ��� �M�<m���]ٿ볿_Ph��G�D�A���V�P��wZ���/ɿЭ�g� �U�����sۿ����¡���(~��U��D5��������<aȾ�u��Ĝ��z륾=q���1žw�⾯l� ����1�v�P�!kx���J����f׿����t��u��k�3�̿� ���(��@�Y��HB���E�fc����� ?���;ֿ[���+`��K������ѿ��S����Pr�^�L��p/��t�����U`Ⱦ�:��ˢ���\�����-�پ���̈��4'�"B��c����������Ŀ��Ҕ���"�G� �Q��eĿ'����u�W���H�� U��){��͛�����;��G� �������'��A�ɿ%���[��FTk�J�H��-�������zξY���5ܻ��Yþ��վ7���	��a��H6�� S���w�u�������vRӿ��sI����������*���w藿�gx�RX�B�R��g�!Պ��嫿ݼѿ�9��'B��P�L �f��Z¿���=]��ڄe�&�E��+��)����פ�g�Ҿ��ƾ�ƾ6�о\c�e�ŗ�?�(��B���`��n��=K���⽿��߿����������m���zWտ\t��
���S�j���R���U��ys�Pz��&ܷ���ݿ������ݦ��u����ؿ�����8��׃���Y���<�^n$���B�����.ξyiƾI�ɾR�׾���f���6���1�y~L��n�aߌ�[Ш���ɿ���Fc�X��ބ�6`�*`ɿk��儿�#a��7R�=^�����?���Fſ��鿀���  �  ��-�պ&����W���M���蔿0�e�a)4�w���w�Ǿ���\������^ڇ�,��[��������9Ͼ\\�����xJ>���s��8���̿�� �8��)� �-�N�#�7�+�,�������m��`e�����X꠿G�Ͽڪ�~3���*�>-���!�p,�:�]������jT�X	(�g�(T�6d��ʤ�}���1���Z	��M����)�������Wܾ�����#�2N�W���2���]�ݿ�(	���0b,��+��;�sb�
�Կ���;J���f�[lj�����o0��<��{���&"���-�9�+��B�i��0Կr���@Y~�G��{�>����۾����=p��{���=���𕾷O���贾��оX������_7�k�f��{��Tο�&�C�] '��/�B'*�c�z����ǿ F��3���l��|�j���H�¿�������I)�dk0��u)����2����ƿ�Z����p�S?������w�ݾM����+��G���I������7��їʾC����	�;�%�4L�M���m����ӿ�����(-�*1�*1'���I�%��cP��iR~��Uv�����tz��ؿ����z�6/��~1��&�2c��e쿡V���?����d��k8�,d�� ��޾ež�³������0��*"��o\¾f�ھ����r��y�3�`�^����*۴���`V���#���0���/�-y!�A�	�gRݿ�{��Һ����v�Z�z�\ё�&���<�:|��%�H1���.�f�������ڿ�M��JŅ�MIT�ѕ,�m���i���վ�3��dа�T����-�����
 ˾��S��}vA�Fq������ĿpD�������)��92�C�,����� ���̿y����P~u� 򂿧.���vǿ������\+��  �  �&W���M�{S5����/�⿅M����t�Ƌ5�V�	�e�ؾt꯾�S���x��R(q���k�֗t�� ��:���<����;���/B��{��B������m��~<�`�Q�L�V�$J�ߝ.�j!��;ֿ����ɑ���e��w����������.��WU?��mS�=hV��G�H
+��R�s�Ϳ�M��?H^��/&�j����,˾�N���"�������p�r�o��*}�����}����ž������ ��pV��֑�B�ƿ�;��'���D�TZU�whT�4B�'C#��\ ���¿틗��Ⴟ}���������Ͽ�j�N+��H��
W�q�S��?�Z� ���N�����bL�*�����ľۥ��w��ˊ��'������O���ݞ�xܹ��Y�%c��Z7��^t��y���3߿p���3���M��Y��R�P�:�������im���x��`�������w����/进+��7�v�P�A�Y��P��8����[��L�������w@�������4�ƾpQ��Z뙾o���]��`K��ֈ������Ҿ�z��FQ �B�O��`��gy�����t9�%�?�GAU��Z���M��r2�e��g޿mU���������ƿ}'���#���C���W��Z���K��@/�����5ֿM���D�n�\�6������0�Ǿ�g���+��$����������$מּ(�þ?�+7�1���f�����Ͽd�N+���H���Y���X��BF���'���aa˿
��JT��f�ϧ���׿.S�/�P�K�)�Z��]W��GC��#��� �48¿����)�Y��(��R��޾<��3=���Н�IØ�˚�� ����a�Ͼp�����q�A��~�U����T促f�}r6��P�}�[���T�T=�[:�}��[6���6��vF��%����/��˹�9c��:���R��  �  Hhu�o�j��2N�s�&�qb��gi�����:�5��3�Ͼˤ�ވ��/o�~�\�C�W�0�_���u�%w��l����ܾPl��H��>����Ŀ���H0��V��/o�i u�$f��JF�e��}^��{N���O��+`���%ҿ�E���4�r�Y�_q���t�
Uc��"B�j_���㿶u��:�h�%l(�ho���Z���盾�Ѓ���j���\��[��h��y��(6��cǻ���aA"��_�G��8�ۿ����=��`�sWs��/r���\�]9�
g�zؿe西\㍿����5-���q�i��`[B�k�c��u���q��jZ�U�5�&z��	ο�|����S�CI�W���O���Z��Z���Dv��n���r�'���Zv��x���Bؾ����;��ʀ���������GE$�+L��uj��Kw�M%o��/T���-�T��)>ɿJS���V���g���~ÿ����q)�T�P���m�x��m���P�˦)�C� ��ڻ�54��yE�������b��ݟ�[���O��?b��$���󄔾c���Z�Ǿ���� ��LV��"����˿�
�ø3��uY�T�r�1�x���i��%J�-"�O��/Ƽ�xқ��㕿�����ڿy��359���]�@Gu�T�x���g�&YF���k7�*���py�~�8����G�ᾃC��;��6���~{��F��M1��p���Zy��� ܾI	��2�FTp��P�����A����A�jEd�A�w��lv�Pa�l_=����/�%o���`��}d��j{���￢���%F�Ojg��x��u� �]�r�8����A�Կ����`�ra(�$����Ӿ"������jg��/��������4�����CTľ�����rE��셿^�������c�&�7�N��	m���y�N�q���V�[+0����οJ��*��T���"ȿ��� �+�:�R�֟o��  �  �2�tC+�	������ ���x���1L���J$ܾ���H���]�I�A��3�1/��5�MaG���f��[��؄��ñ�I��=�[�����\�ʿ��<��Fd.�s�2���'�����﫵�
ތ�o9k���b��B������Dhҿ�l��1�ƭ/�e12�&�����;�^���}�Ϝ8�j4�kʾf����}�X6V���>���3��3�v�<��aR���v�(���þ V�1�1���t������sݿ�j���#��O1��w0�c\!��M�
ؿ��9����c�w�g�,Q��򇰿�;�}��Ew&�}�2��[0�9��*�5�ҿ����y�g��b)�Ap���
��*�����}���]�$�K��sE�c�I��UX��s�eۏ�8~�����K!���L�Z����m{���3� �+���4�O�.����� �mUʿ�����~�VQi�T~z�����ſ�6��%����-�)d5���-�G���r���tÿV둿W�C��#/�<;��;㛾Rǅ��p��b��`���g��Tz��X��
Ȧ��S;�f�>�-�{�i������xѿև��	 ��1��$6� �+��W����ֺ������{���s�/�����;�ڿ��	��n#�f�3��h6�|;*�m���쿢:��s6��� I���l��	������D���)���s�7"s��|�wI��ޠ���c�� 
�%��zB��y��5��������'���5���4���%����࿇f��3���Ct�t�x�7z��@���������*��<6���3��C#��p	�;ٿ������t��u6�I�
���پ�	��f򗾱���c@|�#�t���w��Ђ�G��������ƾe����y!���V�٣�����A������F$.�K87��e1��W�n��2Ͽfe�������r�+�R��U�ɿ�T ������/��  �  �8+�D$�������f�������;H��/�IDܾ=Ʃ��ᇾ�0c�^_G�wf8�Zn4�`;���L��Vl�W؎�����E�[��A/W�k���x�ÿ� ��G2��'��+��!�ӽ�T��������?e�!�\��ly�����ʿ`; �����Z(�}�*�)�R��Z�ۿs���w���5��U�V=˾ើ�7����[�~fD�H�8��H8�M?B���W�,o|��j���ľ|��</��n��š�eտo������)��)������2п�����~�D�]�[b��\�������ܿ@J	�%���S+�%)�$o��� ��M˿�U��B�b��4'�B����m��q���d����7c�7Q�аJ�C�N���]��Sy�e}��4o���?�@���I��燿ӵ��g뿅6�u�$�s(-��'�����+��~`ÿ�ᗿQ�w�S�c��t��3��\��a��.t���&��-���&�����
�u
��"��?#S��!�3P����|��@���d=v��;h��He���l����2!���A��_�ξ�/�c�+���d��\��Phʿ8} �m��'�*���.��$�J���&�f���]𐿔�u�p�m��+�������Zӿ�y������,���.��\#�+&��)�m��������E�0����뾥9��,u�����0M��+y�dx��/�����d^�������f��hO?�4�� ���ݿ�
�Y!��.��L-����H.���ؿ�	���q��Eun���r����+���a�俦�9#���.�m`,�F��<� �ѿ|�����o�7G4��^
��;۾ u�����LK���π�fz��%}�1����ђ��.��9�Ⱦ�2���6 �WS�1���񺿝��G��v'�ʸ/�W4*�O�+��3?ȿ�������Zm�j}�Ҙ��¿W;����Z�(��  �  �������g ��jԿ�����+}��q>�TA�P�޾�԰��̐��u��X���H���D���K�4�^�?�~�8����b��~T쾂��xoK�����ΰ�!߿���Hc����/3�k���olʿӞ���z��T���L�X�e�cg��sN��KB�-�_}�������
d�HsſQ���?lg�%r.�����Ͼ*˦��[��5	n���U��_I��H�EUS�tj�g��ŏ����ɾ�� �٥(�"�_�_��9���
���������A��Tֺ��葿{�i���M�#[Q���t������ſ������,$���������-����U��R"�����VǾ�{���Պ�%"u�Fb�9�Z��I_�5o��х�Lz��mɺ��q����0@��}����x(ӿ  �,j�����$�����ݿ�e��#�be��S��!b��Ї��/���2ٿ6���v�s����Q#�u�ٿP��^
��.[I��3�����1Ǿ`g���ɑ�'䃾�x���u�$�}�M͈�sT���籾*վ6��Ac'�#Y����g���M�忮a�����`�B��
���3ҿ*Ѧ��u����d���]���v��ޖ��ɾ�Ƚ��R���s����������Ϳ�>����w�s�>�=_�!�m#Ǿ���-��e抾d����]��k����%��X���{�¾�꾂���8��p�DP���3ȿ�i��������VK�q��N�`Eÿ~S��v}z�/9^�M�a�S���	����tͿR��[��Y��%��!�Z���1��F�����b��d/�P}
��#ᾩ�������?���>���-���Ԇ�G��!���I1���оei������xJ�1����ͪ��Lؿ'������f�����2�4���G��i�����n��2]�Luk��i��	���;�ݿ��w���  �  ����A���ԿhK�������d�1`4������}f���������by���f���a�( j�����_��'����ʾ�%��=��f�>���q�����5u���ۿ���ϣ��*3鿫�̿�Č���Z��B;���5�z{I�~Au�����R���N4޿ �G��'W��ʿk+��B���AXT�_(������ܾ�K��D���jH��xu�ӳf�	�e�{r�j'��O����J��Z�׾�y�oi#��?N��͂��죿A�ƿ�L俽
���������6��?m����z�v�L�96�P69��U�cs��F0��ʿ��翑h��ƕ��^~�b��Y*���|�jG�v,��T�ڊ־�����휾�S���R��-�w���|�����\��cí�+�˾@#�M��Eg7��{f�� ���N���Bտ�j�	���97��Cۿ<f��$��g[q���J�g�<�2DH���l�� ��*$����ؿ�v���x��;ڿ�Ƹ��7��Ӫo��J?�������`�׾\���2���x��{L���7���MT���@���ľ;��k��1%��ML�ғ�>f���N¿��⿔}�������v�ltԿ(V��`y��Oj�ҹK��6F��FZ�3��9k���/ƿ ��ft��T���E���%ӿ���܎���d��y8�K�7n����ؾ�⼾Qp��P����i�������L���>���ʹ���Ծo�������3���^�/���1��.ϿԤ쿶j���>��p3�F�ɿ"ե�����UN]��F�`�I���e��F���ɭ�jѿ����F���H��/��ǿA���k���C�T�R>,�yV�MU��	Ͼ���^ ��5���沓�����zU���˃þ���I�αA�v�p�i#��]u���mڿ����}����S��,P࿶_���
��M{�nPT��F��Q�V�u�9z�������ݿ/����  �  �^��w츿b����R����y��Q�wt1�c���������Kþ�ǩ��X��s_�������z��^��ei��:Aʾ��mn�bb�[�8�4�Z����9���`��������Y��o���I��0
����\���5����]��w�)�A�I���w�r������r���g���y3��p����Q��o�l��lG��I)�C������پ���<T�����̉��>������ʡ�A���վ�E���z�T�%��)C�\�g��q��F���n��W��� ���W���ؗ��n|��M���+�%.�����2�-�X�Iф�5���rʳ�/B�����4U��u��8`��<�b���?���#������@E־�\���*��m��"���+��rݠ�*����;�A����Ñ���5�ӱU�&�|�t����������� f¿����ց��1b��Pt�� I��,��"���*�@�E���o��T������{����ÿd���{��9И��\����\��_<�ٕ"�����$����پ���������9��UK��(K��~���H6ɾ�便W�M���+�\NF�U�h�������������
�¿=iſ4���P���Q���Έl�:�E�;O/��A+�P:�{�Z��9��8板���*
Ŀ8�ƿ*���?��t����y}��W�ۭ9�0�!�l��pp���Kܾ`{ľO7��n۩��J��U���=���w�ؾZT��L���d)6���S�g3x�`����H��tq��q
ƿ�Ŀ����;��ꕆ�T�^�O{<�S�+���-��B�/$h�U��/ϥ��պ�!ƿj�Ŀ6췿!���~錿��o���L��1����M�� ��qԾ�Ҿ�U5���ܩ�Kj��o���#oʾSz�P� �"W�N�&�l6@�j�_�%����ܙ��᯿������ǿ:���&����`��.�}���R�~6��y+��4��N���x������O�������  �  ?������o)��WJw���a�-N�i~=��.�����Y����־6x�����Υ�������kZݾ�!��Y7��&"�f�1�M�A���R���f�T�|�(����Ǝ�����\r���O��1.���r�������t
�j"!�Z�@���c�d���Ij��O�B��)v�� q���[�^�I�te9�f�)����i�?N��ξ,M��%0���m�����ʾ�0龌��iK��'�i37�`G�+Y���m��쁿����t���Ō� Â�+�f�_�C�h�#���9W ��!� D��+���M���p�	�������ܐ�hB���y��o�l���X�5&G�h�7���'�/P�[��@1�%�;ߐ�����=��
>ž�|߾�0 � �{x#���3�U\C���S��g��|���	�d0���������'c��@���"������7��6� �e3>��`��f���F���i��6��'����#���l�&Y��iH�a�8��)������;��Ҿ�w¾���+Jƾ-$ھ
�����1��Y�/���?�'GO�	�`���t�4W��u|��ߕ��ѕ��L������G&_��=�C�"����V�+���1��wQ�F�t�o��tڔ��]��ԧ��_Ӌ�;���F|l�f�Y�/�I��1:��)�E?�����5d־�>ɾ�xȾO*Ծ)��۩�����s'���7�}G�SoW��i�<z~�98���h��pΗ�)#��!���tw�{~T�R4�~������P� �h;��f\�g�������������ؑ�����	z��e�<T���D�%�4��,$�q��ٜ��'���Ѿ��Ⱦ�Y̾�ܾ�����!�b���.�(>�<�M��4^�"Qq��|��G3��#��U]���,��w���-m�,pJ���,��i���������)���F�J�i�z���\���  �  vY��X_���`�`��#`���`�Z[_�J4Y�0L���8��f!��"
�����ԾW�;8پ@q��DQ�6'��=� P�|�[��`�-8a���`��`�Za��t_�C<X��J�Y�5����5���3�Ӿ:�Ͼ	�ݾ����!��H�+���A��S��c]�g\a���a��0a��a�%�a��_�عV�WG��(2��`�6���5徎�Ѿ��о�⾷��v��]Q/�8�D���T�I^�%a���`��`��`��`�R]���S�ETC�x�-�x��9  �P6�udо
Ӿi��H	���65�o�J�%�Y��*b���d�P�d��\d���d���d�<T`���U�ZZD�a.����Ů�I��پ�޾�"����ab%�Y+=�?�Q�*�_��f��Zh���g���g��[h�9�g��ob�{�V�|<D��v-������,߾�����c����,�ND�4�W�%]d�8Tj��k��k�:k���k��Fj��(d��9W���C�y�,�֣��z�V�� ��ٮ��@�J��4��K��]��0i��.n���n��vn���n�Yo��Tm��Lf�\^X�wUD��-����������o#�����}$�a_<��R�m�c��7n��$r�
\r���q�r�Q,r��xo��g���W��RB�g}*�����������������'��k?�U��-e�AKn�kq�.aq�q�vkq��_q���m�m~d��T��'>�8Y&���Uc ����V��qk�H%�M�+�e�C��tX��{g��~o�y�q���q��oq�q�q�ѕq��\m�2�b�n-Q��:��#�������A�����=���K�a0�x�G�w\���i���p��r��Er��/r��r���q�S�l�R�`��lN�.�7�������#�����y,����	�F��P%5��fL�C�_��  �  �.�\0>��O�תb�)�x�j���ꍿw�������V�v�G2U���2�GI�A�X����+�M��d:��J]��~��Њ�n�������脿�Rt���^�o�K���;�}#,�l����
�0p��eҾ�9��tD��?���kH��D[ƾ�㾡���� g%�E5�~�D�d}V�~k�a����7��G���81��\Q���1m�WfJ�XK)�5�����P� �/{�2�%�&SF��5i�EÃ�z^��򕏿ъ��j����l�U�W�i�E�$6��r&����Ms�y�澥�Ⱦ	���x_��Ra��h˸���ѾT#�L�
���kV-��=��tM��$`�[�u������B��r���濍�r���%�e�l�B���#�#!�ϒ���f��̎5���W��Vz�n��S���*��x����e��9�l��X�'�G��Z8���(�����\����}о�߽�!\��Sx���|Ͼ���U�y.�?x)�R�9��/I��Z�F�m�R��3���_��Es�����(��Ê`��[>���!������
��i��u(��G��1j�p���3|��3_���ړ�𾋿����l�2�Y��vI��.:��H*��O�$����Kjؾʾ��Ǿ�Ҿ�n�؞�:���{%��86���E��U�)3g���{�h͈��s��!̗�~W��n��[}�e�Z�C]9�������������H�5��bV��Ny��Ջ��x����W���A����A}��wh�ʅV���F�7���&������v]�	DӾ�8Ⱦ�ɾ�o׾ѷﾾ��3!��*���:�*eJ�i�Z�r;m��H���+��YȔ�� ��P3������Ar��PO��60��2�av��I�q0%���@��b�ȕ��GB��i����V������ʋ���*w��Pc�,BR��B���2�"��l��h�������оe�ɾ��Ͼ�@�g������n �(�1��  �  ��g�2���S��#|������"��G����n��N����У�
����c���:�*� ��q�=8%���B���n�z䐿�⨿$�������7B��� ���⏿Ses���L��p-�a��M6 ��ݾ��/k��a��|�����Q|�����^����aо���Z��"�7O>��a�_	��C����̰��#��켽��ֱ�el��4Ⴟ~�U��1�����1�-���P����c�������CѼ�O����a��ݞ��6���qe�p'A�9$$������`�Ҿ.����`��jܐ�ㆉ��"��z����槾.�����޾E� �����-��SL�1Tr�D/��i�������as��E׼��]��i���y��1L���,��E�[�$�� =���d�jc��-�����������������x���g����_�K>�dM#���$;��#)ؾd���쩾D�� ��������}��~�ؾo:��q<���#�Y�=���^����������k����ÿ���k��&���Gho�hzF���,�it%��c1�<@O��I{��H��$e��#5���iſ�	��Ҭ�E���W����}Z�N;�Ӕ"�v�7����ݾ�ž����������8��������վ���h5	�$�,�2��O��pr��Y��b������Tſ{�ſ�򹿃����̼e��A�{-���+���=�W�`�����J���������Ŀ4�ſ팺�P���s����u���Q�u�4�L��eW
�����׾u�����Z ���)��a�����ž�ݾ�������F�"��:�QzY��f�S���v��T)��*�ƿ�AÿR����H���WdX�[�8�!++�>�0���H�VFp�����}��,ֽ��ǿ��ÿ|@��m+��b���l5j�:|H��-�������L��Ѿ�Y��6���*���5��ǻ���ϾB���T��K��  �  sZ�x�6���g������C��}ֿ�����H��ҿ�K��=����`��>��4���C���k�����_u���ٿn_��������f�Ͽ<˭�����x�\�<:.��v��{㾃��S1�����x�(�g���d��To�؜��%�������Ѿ����$����F�T!|��~��q���}࿎��f�����忖{ǿJǣ�����~~S��8�`27��<O�D�~�㽟�;�ÿe���������D�Ŀ���-���_K��!�`����Ծ����������&�q��f�_�i��z�N׋�QP��*���侌5�G-��4Z��艿����H@οH꿋X�����޿�Ľ�U-��,�v�w^L�:��VA���a�3���~���ѿ���)��<$����ݿ�	���4��_�u��MC����s� �	(׾.���#=��P���6�������0���M���������-�׾�� �0O���A�*�r�^��x���>�ۿ��G=��y��$�׿b ���I����l�m�I�g
@���O��x�Q,��ɽ� �߿����qs���p�ظֿ2��������Dj��<�y�{���5ھ󽽾慨�̚�F2���D������a��(2��A�о���6�.���W��h���ͦ�R�ɿ�����0������>�Ͽ�ԫ���� �c�D�H��5G��@_��J���ħ���˿��꿆��������B�&"ͿB���U����[���1�p8�G���M�Ҿq���l��JԘ�ڒ�3���2���R������5ھ&~������]:��Vg��n��;=��-�Կ��������y�����"�ÿ�Q��p��zcX�~�E��M��[m�%�������P׿���m��`V�����1¿�_�����p�M�RT'��
���뾈�˾��N��R�������%��|F��.eɾ\R辋���  �  �.��IA�܈�����׿����|����=�$����ѿ�9��Ȣ��>�W�
:K���^�󉈿����2Hܿ��>���������L��r�̿z���_2r�a6���
��W׾/���ލ���r��X�ZJ��G�`�P���e���������3�¾����dz!�M�U�G���㜸���������7L�H�����/�¿y}���<r�G�P���N��l��L������z��^�	�r������	�[��h���ґ�g\���%���� �ƾ�H���܅��qh�%S��J���L��Z��Au�;��Ԭ��&׾��	��4��'n��ݜ���ɿ�z���K�s��c��A�[����� Ŏ�23h�HQ��PZ�.d��p����Ͽ�Q��1��
��?��Ϡ�M�ڱ�|���dkO�ͯ������7Ǿ�u���S��`r~��[m�h�19n����YW��d����Ǿr���F%��OL�\��v�����ܿ�G��8����x�/"�;�׿��������zc��(W�\�j�����gി��⿑�[��4��8�� �S�ӿ=�������8D�������ȾU��S��y���J��&���𓈾�o��F����྾>�g��	92�Ǝf�.��m����C￫/����A^�������4�ʿ�����"���`���^���|��P��,�ſc����B����	��+��.�ſc���l�*c6��I�)��S��fd���h��U��wF��Q�Mc��O���Rȫ���Ⱦq���zOA�tD{�n`���(п���f��������/
����"��!є��1t�`/]� f��:��}��8zտ�k��=�j@��&�j6��;����ʼ��$�Y��)��9�~�۾^���k ����������w���,�� ���|�������׾n���  �  k���K��抿op����=���$��C+��m#�K����e���ɍ�
\i�2$[��q�����¿s3��)���s&��3+�t�!�]����x���#��D�>�R����ӾY���҄�2`�k�F���9��V7��?�۔S�@�u�8������`�����&��+c�zG����̿����k�(��w*�33�w��X�ٿ�.��p惿�Ua�cE_��؀�7U��=�ӿ���?�ʪ)���)�����|��jҿ���8yj���+�k����b�����2uy��V��HB���9��S<�b�I��)c�`������Ӿ�5���;�m�~�-ū�C�࿽;�� !���+���(�}��n���{4ʿ����S�{��Ga���k��	��$ʹ��#�ϛ��{#�f�,�x+(���S����'Ŀ2�����Z�ߎ"�{e��ϳ��u������Z�l���\�w�W�ؠ]�-zn��%��?�������;����b ��V��k����$�������'�Q.�o6&�d}�5��Nܼ�򨓿D1u��g���}�5Λ��1ȿ�l����l�)�p~.��*%�k����WJ��7 ���L�y��m0�B^���;��������w���v����pc��,����d���O޾��ys7��s������տ
�����W�,���.�~@"����,�῝6���ꋿ9Zq�/Ho��ڈ��X����ۿѢ�V �S�-�!�-�� �r��%�ڿ�_��{��]<�d��iN�)Ӹ�W1�� `���р�E:x��{y�d�gڎ���������m�d����H����EE����t�5$��/�	�+���t��IпF���7ȃ�]/m�mgw��䒿ꓺ����|a�Z0&�t�/�!�*�6H�x����Sɿ�͘�e�?�,�/��Cվ�ڰ�m显�É��L����|�0ۀ��ψ�[E��-@��Ѿh��  �  t �ЯO��⎿>��0;��Xp��,�x�2���*�����G��ƒ���1����o�r�`��Jx�o����*ɿ.� ��:�/�-�0�2���(������ck��䢅�jFB���RӾ5���(���Z�i6A��L4��2�YS:�q�M�
p�֒�W�������d)�%nh����&DԿ���Dp �E80���1�i�$�~'�K��4魿�ˇ��Fg�Ae�2����Ш�W�ۿ.
��"��1��
1��"���	�Oڿ�/���$p��i.�����H���Ε�o�s���P���<���4��7��=D���]��c�� ����XҾP-���>�Ă�ek��鿞����'�^3��0����S����ѿ����pH����f�Y�q��A��5����Q|��v*��c4�sl/���,C��˿�ۗ��(_��_$�4������D5��xO���/g��SW��R��QX��h�Y����������������!�ѵZ��g��_�ƿV����,���.��5�}I-�6��I���cÿ���{�{��l�E"��W���^GϿ���d��0��5��-,��S��s���<��N��P���Ʊ��Y�����rE��d^~�%�r�-yq���z�*����蘾����^ ݾh�)�9��$y��d���ܿt���$�O4�V�5��)��0���'�Џ�iKw�� u�왌�԰����p��&�M5�[5�޺&�D���0o���U��"�>�"p�80ᾐ����p��z����;|���r��5t�w��H��e����������4
L�>P���귿���7� !+�ފ6�J43��"����ح׿N����D����r��}�f���������C�/,-�?
7�]2�O��E��:п7����i���.�ޣ��}Ӿ�V���������B}���w�nd|����$w��ǭ��vMϾ�h��  �  k���K��抿op����=���$��C+��m#�K����e���ɍ�
\i�2$[��q�����¿s3��)���s&��3+�t�!�]����x���#��D�>�R����ӾY���҄�2`�k�F���9��V7��?�۔S�@�u�8������`�����&��+c�zG����̿����k�(��w*�33�x��X�ٿ�.��q惿�Ua�dE_��؀�8U��?�ӿ���@�̪)���)�����|��jҿ���Cyj���+�q����b������ty���V�HB�O�9�UR<�H�I�'c����{��TӾ�4��;���~�9ī�B��:;�f !�>�+���(�"��ݖ��4ʿ�����{�}Ga�Ôk��	��ʹ�g$�#���{#���,��+(�i��\����(Ŀ ���F�Z�^�"�h�����'���%���l���\���W��]��xn��$��������������a �R�V��j����#�����'��.�6&�
}�����ۼ�����1u��g��}�}Λ�g2ȿRm��U�ݯ)��~.�E+%��k�̎�`K��-��ԥL���3�`���=��K��)��w�L�v�T���c������e��P޾���s7��s������տ
�����W�,���.�~@"����,�῝6���ꋿ9Zq�/Ho��ڈ��X����ۿѢ�V �S�-�!�-�� �r��%�ڿ�_��{��]<�d��iN�)Ӹ�W1�� `���р�E:x��{y�d�gڎ���������m�d����H����EE����t�5$��/�	�+���t��IпF���7ȃ�]/m�mgw��䒿ꓺ����|a�Z0&�t�/�!�*�6H�x����Sɿ�͘�e�?�,�/��Cվ�ڰ�m显�É��L����|�0ۀ��ψ�[E��-@��Ѿh��  �  �.��IA�܈�����׿����|����=�$����ѿ�9��Ȣ��>�W�
:K���^�󉈿����2Hܿ��>���������L��r�̿z���_2r�a6���
��W׾/���ލ���r��X�ZJ��G�`�P���e���������3�¾����dz!�M�U�G���㜸���������7L�H�����0�¿y}���<r�H�P���N��l��L������~��a�	�u������	�h��$h���ґ�|\���%�����ƾfH��]܅�zph�g#S�K
J���L�ִZ��<u���1Ь�"׾A�	��4�Y$n��ۜ��ɿ
y���J���������I������Ď��2h��GQ��PZ��d������Ͽ�R�������1��ˡ�G��۱�G����nO���������;Ǿ�x��
V���u~�~]m�:h��7n�Z�� U���`���Ǿ����`"�6LL����������ܿ�F��7�������!�0�׿������:zc��(W���j����6ᴿ���C�0��5��9�� �e�ӿ:���f��-<D�����j�Ⱦ�X��V��춊��K���������}p������ι�侃��92�Ўf�0��n����C￫/����A^�������4�ʿ�����"���`���^���|��P��,�ſc����B����	��+��.�ſc���l�*c6��I�)��S��fd���h��U��wF��Q�Mc��O���Rȫ���Ⱦq���zOA�tD{�n`���(п���f��������/
����"��!є��1t�`/]� f��:��}��8zտ�k��=�j@��&�j6��;����ʼ��$�Y��)��9�~�۾^���k ����������w���,�� ���|�������׾n���  �  sZ�x�6���g������C��}ֿ�����H��ҿ�K��=����`��>��4���C���k�����_u���ٿn_��������f�Ͽ<˭�����x�\�<:.��v��{㾃��S1�����x�(�g���d��To�؜��%�������Ѿ����$����F�T!|��~��q���}࿎��g�����志{ǿJǣ������~S��8�c27��<O�J�~�罟�A�ÿl��!���#��� �W�Ŀ���?���_K��!�i����Ծ���
��������q�7�f��i��z��Ӌ��K������㾳1��-�0Z�承�����=οsE� V������޿^ý�<,����v��]L��:�FWA�˽a� �������ѿ����+���&��n�ݿ����7��l�u�@RC���� ��-׾簷��@������p�؀��(���K��B�����Y�׾� �K�یA�
�r��������n�ۿR
���:��N��U�׿�����H����l���I�s
@�w�O�"x�l-���ʽ��߿&���v��fs񿺻ֿ���|����Ij��<�N}������ھFý�n�К�5���F��(��c��3����о�� �N�.���W��h���ͦ�R�ɿ�����0������>�Ͽ�ԫ����!�c�D�H��5G��@_��J���ħ���˿��꿆��������B�&"ͿB���U����[���1�p8�G���M�Ҿq���l��JԘ�ڒ�3���2���R������5ھ&~������]:��Vg��n��;=��-�Կ��������y�����"�ÿ�Q��p��zcX�~�E��M��[m�%�������P׿���m��`V�����1¿�_�����p�M�RT'��
���뾈�˾��N��R�������%��|F��.eɾ\R辋���  �  ��g�2���S��#|������"��G����n��N����У�
����c���:�*� ��q�=8%���B���n�z䐿�⨿$�������7B��� ���⏿Ses���L��p-�a��M6 ��ݾ��/k��a��|�����Q|�����^����aо���Z��"�7O>��a�_	��C����̰��#�����ֱ�el��5Ⴟ��U��1�����7�-��P����j������OѼ�_����a��,ݞ��6���qe��'A�T$$�������Ҿ�����_���ڐ��������珕�F⧾y�����޾%� �(�Y�-�NL��Mr�,��6��������p���Լ��[�����-�x��/L���,��E���$�
=���d��d��"���⁸�D�������1�����k����_�  >��R#�U���B��/ؾ����奄���@������S���y����ؾ+3��8�o�#���=�C�^�����R��ŕ��<���ÿ���ti��z����eo��xF�)�,�vt%��d1��AO�]L{�gJ��[g���7���lſ���|լ���������E�Z��S;�$�"��z�'�����ݾo�ž?��f��2���9	��{�����վd��5	�;$�H�2��O��pr��Y��b������Tſ{�ſ�򹿃����ͼe��A�{-���+���=�W�`�����J���������Ŀ4�ſ팺�P���s����u���Q�u�4�L��eW
�����׾u�����Z ���)��a�����ž�ݾ�������F�"��:�QzY��f�S���v��T)��*�ƿ�AÿR����H���WdX�[�8�!++�>�0���H�VFp�����}��,ֽ��ǿ��ÿ|@��m+��b���l5j�:|H��-�������L��Ѿ�Y��6���*���5��ǻ���ϾB���T��K��  �  �.�\0>��O�תb�)�x�j���ꍿw�������V�v�G2U���2�GI�A�X����+�M��d:��J]��~��Њ�n�������脿�Rt���^�o�K���;�}#,�l����
�0p��eҾ�9��tD��?���kH��D[ƾ�㾡���� g%�E5�~�D�e}V�~k�a����7��G���81��]Q���1m�YfJ�ZK)�7�����T� �5{�:�%�0SF��5i�NÃ��^�����&ъ��j����l���W���E�E6��r&����$s�ҝ澔�Ⱦr�9]��D^��bǸ���Ѿ��Y�
�[��Q-��=��mM��`�Gzu�����?��d���4���+���{�e���B���#� �������۰�"�5���W��Zz����V���-������i��h�l���X���G�j`8���(����7`�����"о�὾F\���v���yϾ뾡R�R*�;s)���9�)I��Z��m�����)0��H\��)p��9�����0�`�MY>�%�!�-����
��j�rw(��G��5j�͕����nb��Oޓ��������l�i�Y�N}I��4:�$N*�ZT��'����1oؾ�ʾu�Ǿ�ҾLp�r�����1|%��86���E�-�U�/3g���{�g͈��s��!̗�~W��n��[}�e�Z�D]9�������������H�5��bV��Ny��Ջ��x����W���A����A}��wh�ʅV���F�7���&������v]�	DӾ�8Ⱦ�ɾ�o׾ѷﾾ��3!��*���:�*eJ�i�Z�r;m��H���+��YȔ�� ��P3������Ar��PO��60��2�av��I�q0%���@��b�ȕ��GB��i����V������ʋ���*w��Pc�,BR��B���2�"��l��h�������оe�ɾ��Ͼ�@�g������n �(�1��  �  vY��X_���`�`��#`���`�Z[_�J4Y�0L���8��f!��"
�����ԾW�;8پ@q��DQ�6'��=� P�|�[��`�-8a���`��`�Za��t_�C<X��J�Y�5����5���3�Ӿ:�Ͼ	�ݾ����!��H�+���A��S��c]�h\a���a��0a��a�&�a��_�ٹV�WG��(2��`�8���5徕�Ѿ��о�⾿�����kQ/�K�D���T�j^�La��`�!�`�O�`��`�9R]���S�>TC�P�-�$��� ��4�"bо�Ӿ1�羏�"��15�s�J�g�Y�0$b���d��d��Ud���d��|d�N`�Q�U��UD��.�-����1�徖پV�޾�%��R��e%��/=�P�Q��_���f��ah�ch��g��bh��g�vb�߱V� AD��z-�������-߾J��7����6�,��D�كW��Vd�ZMj���k�k��k�M�k��?j�U"d�-4W�7�C��,�7��(y�����徺��B��C4�BK���]�Q7i�
6n�y�n�e~n���n��%o��[m�dSf�dX�JZD��!-�ޜ�*�����&��������}$��_<�7�R���c��7n��$r�\r���q�r�Q,r��xo��g���W��RB�h}*�����������������'��k?�U��-e�AKn�kq�.aq�q�vkq��_q���m�m~d��T��'>�8Y&���Uc ����V��qk�H%�M�+�e�C��tX��{g��~o�y�q���q��oq�q�q�ѕq��\m�2�b�n-Q��:��#�������A�����=���K�a0�x�G�w\���i���p��r��Er��/r��r���q�S�l�R�`��lN�.�7�������#�����y,����	�F��P%5��fL�C�_��  �  ?������o)��WJw���a�-N�i~=��.�����Y����־6x�����Υ�������kZݾ�!��Y7��&"�f�1�M�A���R���f�T�|�(����Ǝ�����\r���O��1.���r�������t
�j"!�Z�@���c�d���Ij��O� B��)v�� q���[�^�I�te9�g�)����j�BN��ξ1M��+0���m��)��-�ʾ1龙��{K�-�'��37��G�VY���m��쁿����t���Ō�Â��f��C���#��V �Z ��A�k�+�:�M�k�p����ɳ���ِ� ?��@v��e�l�֙X��G��|7���'��K����,꾗�;玹�5��e���@ž�߾�3 ���:}#�=�3��bC���S��g�F�|����j���z3�����`���i+c���@�p�"�������p���� ��0>���`�]d���C���f��������� ��.xl�Y�GcH���8��)�M�^��S�쾄�Ҿ1v¾����Kƾ�'ھ4��!�������/���?��MO�P�`�.�t�[��1����╿�ԕ��O��푀�E*_��=���"���MX�G���1�xQ���t�����ڔ��]��ا��`Ӌ�;���E|l�e�Y�/�I��1:��)�E?�����5d־�>ɾ�xȾP*Ծ*��۩�����s'���7�}G�SoW��i�<z~�98���h��pΗ�)#��!���tw�{~T�R4�~������P� �h;��f\�g�������������ؑ�����	z��e�<T���D�%�4��,$�q��ٜ��'���Ѿ��Ⱦ�Y̾�ܾ�����!�b���.�(>�<�M��4^�"Qq��|��G3��#��U]���,��w���-m�,pJ���,��i���������)���F�J�i�z���\���  �  �^��w츿b����R����y��Q�wt1�c���������Kþ�ǩ��X��s_�������z��^��ei��:Aʾ��mn�bb�[�8�4�Z����9���`��������Y��o���I��0
����\���5����]��w�)�A�I���w�r������r���g���z3��p����Q��o�l��lG��I)�C������پ���?T�����#̉��>�����ˡ�S���,վ�E��{�n�%�*C���g��q��\������h��� ���W���ؗ��n|���M��+�$-������2���X��τ�D���"ȳ��?�����R��?��
]��&�b�H�?���#����}��E?־$X���'�������!���,���ߠ��-��	�;\H�������J�5�ݷU���|��������������h¿��������c���t�W"I��,��"��*���E�I�o��R�����#y����ÿ�`���x���̘�rY��b�\��Y<���"���q����پw�������S8��mK���L�������:ɾ.�侗[�����+�ZTF�׎h�X����$���P�¿=lſڬ������,���ǋl���E�Q/��B+�Q:�1�Z��9��b板���9
Ŀ?�ƿ-���?��s����y}��W�ۭ9�0�!�m��qp���Kܾa{ľP7��n۩��J��U���=���w�ؾZT��L���d)6���S�g3x�`����H��tq��q
ƿ�Ŀ����;��ꕆ�T�^�O{<�S�+���-��B�/$h�U��/ϥ��պ�!ƿj�Ŀ6췿!���~錿��o���L��1����M�� ��qԾ�Ҿ�U5���ܩ�Kj��o���#oʾSz�P� �"W�N�&�l6@�j�_�%����ܙ��᯿������ǿ:���&����`��.�}���R�~6��y+��4��N���x������O�������  �  ����A���ԿhK�������d�1`4������}f���������by���f���a�( j�����_��'����ʾ�%��=��f�>���q�����5u���ۿ���ϣ��*3鿫�̿�Č���Z��B;���5�z{I�~Au�����R���N4޿ �G��'W��ʿk+��C���AXT�`(������ܾ�K��F���mH��u�ݳf��e�${r�u'��^����J��t�׾�y��i#��?N��͂��죿S�ƿ�L��
���������6��&m��%�z��L�g6�*59�~�U�[r���.��^ʿ��Nf��H����{࿵���'���|�{eG�[(�fQ��־+���ꜾTQ��!Q����w�K�|�����#_���ǭ���˾�)�;���k7�f�����Q���EտPm�|���b9�Eۿ�g��%%���\q���J�w�<��CH�b�l������"����ؿ�t�	�����8ڿ�ø��4����o�!F?�������~�׾�����}��:��gK��	8��J򍾸V���D���ľe��"�B6%��RL�%��i���Q¿���[������-y�VvԿ�W���z���Pj�K�K��7F��GZ�|��kk���/ƿ��qt��Y���F���%ӿ���܎���d��y8�K�8n����ؾ�⼾Rp��P����i�������L���>���ʹ���Ծo�������3���^�/���1��.ϿԤ쿶j���>��p3�F�ɿ"ե�����UN]��F�`�I���e��F���ɭ�jѿ����F���H��/��ǿA���k���C�T�R>,�yV�MU��	Ͼ���^ ��5���沓�����zU���˃þ���I�αA�v�p�i#��]u���mڿ����}����S��,P࿶_���
��M{�nPT��F��Q�V�u�9z�������ݿ/����  �  �������g ��jԿ�����+}��q>�TA�P�޾�԰��̐��u��X���H���D���K�4�^�?�~�8����b��~T쾂��xoK�����ΰ�!߿���Hc����/3�k���olʿӞ���z��T���L�X�e�cg��sN��KB�-�_}�������
d�HsſQ���?lg�&r.�����Ͼ+˦��[��9	n���U��_I��H�QUS��j�g��ӏ��îɾ�� ��(�4�_�i��E���
���������;��Cֺ��葿�i��M�QZQ���t�N�����ſ�������C#�����(���,��H�U��O"�����RǾ0x��[ӊ��u�Yb���Z��J_��7o��Ӆ�F}��@ͺ�cv�΄�4@�r}�����p*ӿ �$k����h%������ݿ�f���Ice�%�S�6!b��Ї�4/���1ٿ���v������M"�p�ٿ_������WI�1�����Ǿ"d��1Ǒ��⃾��x���u�ݫ}��Έ��V��^뱾\.վϷ�Jf'�q&Y���m���g�忼b�����a���q����4ҿҦ��v����d���]���v�ߖ��ɾ�޽��R���t����������Ϳ�>����w�s�>�>_�!�m#Ǿ ���-��e抾d����]��k����%��X���{�¾�꾂���8��p�DP���3ȿ�i��������VK�q��N�`Eÿ~S��v}z�/9^�M�a�S���	����tͿR��[��Y��%��!�Z���1��F�����b��d/�P}
��#ᾩ�������?���>���-���Ԇ�G��!���I1���оei������xJ�1����ͪ��Lؿ'������f�����2�4���G��i�����n��2]�Luk��i��	���;�ݿ��w���  �  �8+�D$�������f�������;H��/�IDܾ=Ʃ��ᇾ�0c�^_G�wf8�Zn4�`;���L��Vl�W؎�����E�[��A/W�k���x�ÿ� ��G2��'��+��!�ӽ�T��������?e�!�\��ly�����ʿ`; �����Z(�}�*�)�R��Z�ۿs���w���5��U�V=˾ើ�7����[��fD�L�8��H8�S?B���W�6o|��j���ľ���D/��n��š�eտr��"���)��)������2п옠��~���]��b��\������=�ܿ�I	�â�S+��)��n�I� ��L˿�T����b�\3'������k��������5c�6Q���J���N�_�]��Uy��~��+q��*B侬��^I��臿Ե��h�7���$��(-��'���,���`ÿ◿��w�Y�c��t�x3���[������s�9�&���-��&�+���	�q	��1���!S�Z ��M�g���z������;v��:h��He���l�y���"���C����ξ1���+�g�d��]��^iʿ�} ������*��.���$�����'�ߘ���� �u���m�,�����[ӿ�y������,���.��\#�+&��)�l��������E�0����뾦9��-u�����0M��+y�dx��/�����d^�������f��hO?�4�� ���ݿ�
�Y!��.��L-����H.���ؿ�	���q��Eun���r����+���a�俦�9#���.�m`,�F��<� �ѿ|�����o�7G4��^
��;۾ u�����LK���π�fz��%}�1����ђ��.��9�Ⱦ�2���6 �WS�1���񺿝��G��v'�ʸ/�W4*�O�+��3?ȿ�������Zm�j}�Ҙ��¿W;����Z�(��  �  ��꿕�ῘUɿ�̧������J�M�r%������4��LR���/��N�e��^�����7��R�6�I#]��G���K���<���!�	�W����p��"Aп��%���޿�¿����68���WM���/��*�=H=���g��𑿣P��k�ӿ���0�꿄�ۿ�d��f���d.t�&�8�
��ξ�X��~�v���H���*����D����2���'��D���o�J���Ǿ-*�kx2��pl��B���Y����ؿ_�{Y�{
ֿ���6N����l��`@��*��-��I��}z�r����0��:�ܿn��~�迫տ����`R���Lb��	+��� �
þ�����t�EM�[�4���&��%"�.�%�KO1�c�F�4�h��㍾�T���龶����K��ń�Χ�9�ɿ������v����п�R��vi��~d��>�Q1�CO<�j_��[��o&���tο翣F�rH�+�οG?�������T�@�!�P���ҿ�܂���U�
�]��!I�b�>��<�<�B�bzQ���j��ۈ�Y񥾵@о�2�
�/��ue��n���ܶ��׿���A�iX��mʿ����-���k]�;�?�&�:�g�M�B=x�$P��걼�6�ۿ������1俾�ǿ�ˤ��P���.I��Q���/����~��cy����j���X��P�QoO�`W���g�����ᗾ�z������a�u�B�E�|��z����ÿn���f��8f޿������P�}���P�+;�v�=�*Y���:Q��ߌǿ���W�򿯕￳�ۿa7���֘�So��8����ܾ�@��Le�����e��+W�plQ���S���^��s�����-���IȾE���� $���U��ቿ�묿�Ͽ��X�����+�տH���N���m�XTH���:��E�ʠh��᏿�����ҿ�R��  �  ��+;ٿ����F��㤀�x9E�$���M߾�������])V�=4�~����X�����#��S;�^a�w����+��K���9OR��D��mꩿ��ȿTݿ���Щտ�㻿>����x�[�G�nC+���%�3q8�4�`�}<������ɣ˿W�޿��xӿ�����j��xZm�O�4�t��;f��z���L��R/��#�$;�Ҭ�m�!J,��IH�# s��,����ƾk�#�.���e��W��]���L�пYZ�yd߿Xο�,��xn��u�e��g;��&�k)���C�h	s�r}���N��!wԿ���W�߿AͿ�_��-̍�s}\���'��8��n�¾X�����w�^Q��8��+�8;&��)�y�5��K� �l��l��g���ip�ȃ�D�F����lI����¿yJۿ8��]%߿{HɿvW���
����]�4/:�5-���7�1|Y��)��t^���ǿ�z޿�,翜�޿�[ǿ܉�����!P�8r�!9��7��m��������b�:nM���B�d�@���F��U��o��Ɋ�%/��о���Ā,���_����_����`ϿI�����~�ܿ�Xÿ4@���1��e�W�z�;��u6��I�S�q�ؚ��ZX��WԿw�������ۿ!���*�����}��)E�rb��f��3��Ӗ���`o��]�<T�ۈS��M[��9l��)��ŧ���\��C羗��?�Sv����뼿��ؿ��ֻ�P]ֿۈ��nȘ�o�v���K�m�6���9���S��R��Y��ɧ���ۿԖ�]�濂�ӿ3鵿�O�� �i�:�4�3���ܾ�c��}I��C���3j��\[�&�U���W�u�b�djw����r����Ⱦ�'���!�7Q���vh���ǿAl���꿸9�OοN��)�r�g�h�C�M�6�O3A�w�b�ɭ���ȫ��[˿����  �  E.ɿ����&𭿧����=l�w�8�C�d�۾(M���&��n�c��GB��4,����O��L&"���0���I��_n��~���n��q��iX�^�C�ly�x�������q%ſaKɿ�̾�d���^����.c�Sn8��G�ԛ��*�HkN�*Q�������4��k�ƿ��ȿ���` ��c����G[��t*�V��si̾��������
[��`=��{*�v!��j �|�(�?H:��lV����)���7ƾ���� %���T�o0������������ǿ�ǿ/2���`��}����R�:�-��"�@��n5�r^�/���������3ʿ�ǿ�ͷ�{m�����5M�ߛ�� ���eþh��	}���_��F��48�!�2�'~6��C��9Y��z�O��j}����"���;���m�f~���"���+Ŀ�%Ϳ%qǿ5���N��N|�J�L��`-�-�!��b+�I��8w�*���1貿ǿ+�οD?ǿ�b��I7���(w�DpC��/����Ua¾�u��d����=p��[���O�]JM��S�c�,*}�bo��"���[Ѿ�]�7�$��Q�����BV��Z}��f̿�Zп�ƿ-��;b��z�r�WkH���/��+��{;�5_�����������=�οrVѿ�Uſ�L��������k���:�W�����¾�O��힍��m}��mj���`�F`�6�h�7z��:���[Y��p�澤���i5�4e�Fh���꪿��¿'Eп?tϿڊ��ѹ��Je���ic��>��+���-�E�D���m������୿�ſ�ѿؖο�d�����>:���:Z���,�~	�(@ݾ���8ٛ��ˈ�,�w�>xh�5b�8�d� \p��Ȃ����0q��
z˾�w���,TE��.x�M���~F���Oɿ�Eҿ�̿���������gV�L�6��K+��4�*+R��������'1���<˿�  �  R���s6��v��.�|���P�	)�����3ܾ󿴾s������gG]��E�K�6��3��9�+8J���d��n���w������=��2�`A[���������Ӥ�,ا������!���'p��D��="�����	��@�[4��e\����Ԙ�⤥�#���ڵ���9���Lo��/D�3U�ca����Ͼ�櫾(_��4�v���W���B��7��7��@��iT��"r�2F��Yާ�a�ʾs����;?���i�욊�3���e㦿H���R���ˆ���`���7�F_�xj
�
�����z<A�Csl�@����)��dܨ��I��z ���ԇ��c��:��������Өɾ����C.��{��g`��O��gI��cM�7�[��s�d(��z꡾d���65澑_���,��T��������I�H���I��^���[��45Z�x&4�^��7V��.� U1���V�	����9��������Y���/���$ჿ�[�9�3�����"���ʾo��+l��}���1�s��f�o�c��$k���|�4���&��X��,\ؾQS����Ƨ?�E�h��{��Ig�������䮿����}���xX��WT��!2�
���K�C�'�ðD��m����L2���������	��ׅ�������T���.����n�26̾ɐ�������䋾�P��w�w���v�EF���+�����8\���Ⱦ�	뾄��qX*�fsO��.z��ڒ����1��,c����������Nq��H���)�x�����@h/��P��n{������3����������`����\��?�p�`G���#�s^�e��͝¾І�������Ȉ�����x�h�{�"����.��
꠾E����Ծ/���ȫ���6�,T^����������(Ѱ�m5���j��uX��Ed�q�=��G$�3���u"��q:���_�R���{���<���  �  ���Oⁿ�6p�T�T���7�A1�z�����)ɾv���tΗ�⪄��!l��'Z�JU��d]�uSr�A���*��!����tоX��F���q#�o�>�S'\�Iv�E����1��ת}�� d�GvC��#��		�����$� �j��;�4��+V�L�s�t�����T��I�h��rL�{�/�@Q�H��Q߾����骨��㒾z���5h�$-Z��TY���e��8~�Y��皥�<h���۾A��A��5,���H��?e���|��ބ�������u�� Y���7�<&�T�@��l�R�p� ��0A���b���}�[I���Ӆ��)|� �b���E�*�`��u����۾�C��Z}���b������vt��ik�1:p����8���7����ЇԾ.A����0"��<�|�Y�S\u�����!���a����t�=V��5��z��6�k9��e*�q����2�� T��s�+����u��rT���({���_�}�B��(�������{?߾��ľ�i��q���4n��V���t˂�gm��6_�����J��V}Ͼ�K����Qi�Z1�}�L�R�i�v��Q����:�������r���R��2����+}	�n���"��'�vE���f��B���ϋ��؍��1��H�y�u�\�?@�Ұ&��c����EL⾮�Ⱦ����������������͒���`[��u�ž��޾�c������#�K�<�=�X���u�����L*������<��S�i�1yH��)�z���"���W���0�}	P�v�p�JㅿJ������v�����o���R��7�
��4������پ%���HZ�����#��/b���Q��6×�0量Y¸��cϾЖ龆��A��v,���F�p�c�-��R:��`G���~����`���>��/"������>f�'��G�;�(�\��W|��щ��  �  �CN�M��0D���6�b�(�G5��=�>��;���־?T���c����
������!� ��ݪ�o�þ�fݾ�[�����b�s��gd,���:��G��O�r5N��C�N1��������y��ɾN�ž|Ծ ��՟�;S'���<��K��0P�L�JA��H3��%��<�)��v���龽eоXﶾH�������	c��]���ꕝ�I޳��;������e�
�h��#��1��+?��J�ewO��`K���=�mL)����)���N�־.�ƾZVɾ�޾\�������0�ځD�qfP��R�L��?�~�1�r�#�"��y�Г �ڷ��OϾض������e��6��AS���`���¯���Ǿ5�K���S
����Ƈ!�e�.�� =���J��kT�F�V��nO��N?�U)�)������c߾�Aվ�)޾w�������n(�24?�<�P� Y��
X��'O���A��~3�%&��-������M�d�ӾY���H���S���3���f��#��onľ�ݾ.���6��f�>���P,��:�u{H��CU��\�CA\��R���?���(�WG�%������D��.���z
�<7 ���7��9M�I�[�+�`���\���Q�v�C���5�ƛ(�N���L��#�S��׾���嘮�*㤾mN���쬾U����Ӿ�"�b�O���2�&��e3�zA���O�[�d`���[��uN�d�9�B9"��0��[�����t��������̤'�!	?��lR���]�)�_�EY���L���>���0�@�$���x�$$�-�辯�Ͼ����j����社B���u*���ƾZ�ݾ�����z��m�N���+�~9��mG��U���^�K�`�٭Y��tI�)Z3�A���:��z� �0��<q��c1�l�G�߸X��  �  H`!��#&���'��'�r�'�i�'��)&��>!������	��>��hҾ+趾c9��S���J��������پ�N�������5#�6O'�w(���(�)�(�#Y(�kU&��� �r���&��Ĩξ����@����ӡ�'��4¾��ྈ	�F������$�d,(�;)���(�
)��(��&�������T����龷6ʾ�u��n����ڢ��0���ƾl��'�����X�1/%�q�'��(��f(��a(�p�'�H�$�t�B���[�\���ľ� ��/Ǣ�r֤�����C�;���%t����D�"�x#)�/�+�5,,�?5,�PC,�xe+�:�'�3��n��� ����jmɾ�s��[�����ӄ��
�۾�����2������'��c-��^/�؟/��/���/�c.��)*��!�,~�ȃ�w!辻�˾����(���'�����ʾ']��s�?�5�"�S=,��1�ǣ2��2�V�2�>�2��1��8,��"��)����/^�P;ξe＾�6�������վ_K󾡖
����(��0���4��6��*6��@6��6�5.4���.�B�$�����a���ӾGcľ������̾���� ����7d!���-��_5�Y�8�6�9�-�9��{9�@�8��a6���/���$�a����:�kѾ�þ��¾�Ͼ��F��r��J�"��z.�a5�bB8��8���8���8��28��$5���-��7"�������K��4ξ|�¾�ľҕҾ��Q����1p%��B0�ip6�<�8�;99�89� B9��_8���4���,��` �#��/�������̾�þ��ƾ�a׾� � c	�����7(��G2��7�i�9���9�X�9���9�E�8��{4���+�����������'߾?�˾Fľ�Gʾ��ܾJ������_W�@�*��  �  T;������iI)���7���D�\�M�PN��kE�g�3�tG�'��|�.2˾8�þ��Ͼ0�쾱'�R�"���8�0�H��wO���L�'�B��65���&�=��'�ۣ�rl�Ծ6���a�����N���_���+׊��X������Rɾ���x��U	�5���]!�8D/���=��I���O��M�YvA���-�gK�>U����۾[@ȾE$Ǿ��ؾ�����|��+��O?��GL���O�%AJ���>��J0�%:"����k�	�����\���ʾ���v3���V��٧��zH���������j����վ���wR�������)�Q7�|LE�a�O���S��N��>?�X�)�/|�)���hkܾ�2Ͼ�Ծ���!�	�:!��}8�K�U.U�w�U���M�3A��2�c%�E�������"'뾧�Ѿ�9���kB��n���5������󹾶�Ҿ����,�Q������&��F4�ŬB�X�O� �X��JY��zP�3 ?���(��f�v������2�۾��羱��^��{�/���E�y�U���\�3ZZ��P���B�
�4���'�������:����nؾQX�����F������.������о�(����b�����|%�K�1���?�bN��Z��@`��]�4�Q�"�=��U&���������,辐����?��{#��;�GbO��g\���_���Z��N�Y�@���2��&��u�8���������Ҿ\���R���.���C��Pm��bC��\ؾ<��������L��)��6��OD�[ER���\���`���Z���K�:�6������	�I������bM�	��G��D,��QC�g�U��_��`��3X�L]K�=��q/��H#�����2��������b;����_L��34���l��uc���N˾_��^c���K��  �  <i�g���w��w9�y�V�<�q�
Y���$������Ah��`H�+�'���=����꾱��Q���.�RP�`�n����4r��E����l���P���3������������ž�������;���j���Z�{X���b�Qay�K�����4m���־A���_���K(�QD��Sa��Zz�����qۄ��z��-_�G&>��m����e�+��ܦ��#��E:��p[���w��6��r䄿V*|���c���F�ا*��������%�ؾX���ͣ��莾H[|��6e��mZ��]��m�����L�������.Ⱦ�Y��g���}4��TQ���m�|��iY���턿�/v�]ZX��47����-o��_�����*���\*�".K�7�k����������ˆ�v�{�Иa�{D��()����>R���ݾ��¾���9	��������~��Mx�J�P���	��t�E�ľq�߾�;��#���x)��vD���a�՞|�g҇���������rs�öS�;3�I��Z�]l�$�	����QP;���\���{��������S����Rz�wt^��A���'���������B⾒�ȾB-���O��e&��ܻ���ˋ��v��,=��� ���þ�۾����
}��� ���8���T���q�[��wҌ������Q���Bo��/N�7n.����N(��d�����+��CJ��vk�F���F��9���&4��=4t��]W��;�RI"��������0ݾ߀ľc�� Z��6d��L����P���������|���ʾע��� ��H���'�J�A��L^�ͦz�����ō�_N��3i����d�"�C���%�^w�����
�/�I�5��HV���v��뇿�䍿�����%��C�k���N��3��*����3��׾��ϫ��a���c��Q����̑��E���L��|Ͻ�g	վ
���  �  �6޾il	�s�*�PS�zL�+3��]䢿pɧ�P��X&��sw���J�w&��e�y���A�P�-�؆T�p��������飿Q�T���L��23v���J��#�����B־}����ԓ��{�>[���D��68��6�@#>��nP���l����T����ľM���
���8��c�lt������uO��+j���Y���ˊ�M�h��x>�k������+��$:�վc�gL��������zͦ�W�������_g�b�<�_�4M���Ⱦ���������o�4!S��@�u�8���:�Q�G�ެ^����Y֕�k��I�׾���P#�X�I�%u�����2������{���̙�����8^�L�6�̹�������)�ЇL�nvx��N��v���G���������p�-�_�<7�9��&y�DJʾb�� Z��I���##j�v"[�hV�H\���k��ꂾ�񔾐���x�˾����i���5��P^�1#�����t^���H���ڦ�����1���hV�a2��/����T���9�F�`�e������>r��t��� X������ⁿKGX��n1����.2�n�̾��O��'����‾agv�P9u��?~�N������ ���trľ�澄	�Ƣ%���I�K�s�檏�k���fr��Ń��+k��֒�>�x��xN���-�'��
��+�;J�ӻs��N��s���<���+㮿/��i���J�w�_9M���(���4��#uƾ-���8������{��%�v�7x��ρ�蠌�vy���ͱ��;yy�	R�9g0���V�����Xz��s������wd��E�������j�M�B���&�h�R=�B�4���W��Ё�<Ǘ�"Ө�u����﬿K4��d��FAj��^A�����F�޾�i���q��Ya��yw��������{��!��	����"�������'��E�۾�  �  :l޾)�;��Lo��_���X���¿�IɿF#��ϐ��J*����j���=��q!��F�8'&�\�F�,�v�ۥ���#��jbĿ`Xɿ�����N��9�c�d1�A��M8Ծh-��C↾�`�܌@��&,�ZU!�bx�u&���6��*Q�MEx��������:�����}�L�����Wl������ǿ9�ȿ�󻿱\��%���H[�+3��1�`����/�D�U�H�9��0�����ǿ2�ǿ,����?������6�Q�٥"������ þVԚ��R|�DT�,W9�&)�B="��n$���/�IoD� d�R��� ���דԾ{V���/��wa�W���
.��gÿ��˿��ǿ�򶿖'�����~P�O".��$�?+%���?�<nk�2�������¿�̿��ǿ;ε��m��M[}��OH��]�T�����¾5���������g���P�)�C���?�^�D��R�$�j�����Q��y�þ�J���(�1F�QOz�Sݙ�vӴ��.ȿ5�οȯƿ�-��ږ� v��pI�Z7-�~*%�^+2���R�آ��\ꝿ'���4�ʿ~�ϿxOƿvװ�h��(iq��0?���\!�zþ���W���G|��i�qP_��y^��_f�.\w�v>��!	�����:#���A,/�$T]����������I0Ͽ,�п�Ŀ�f��F)��EHk�?C��&-���+���?�?�e�v쌿�;��S���9�Ͽ��Ͽ����d���͌�%Qb�(3������㾷�������$d��5.y��h�@`��Pa��Nk���~�Ք������&�þ�e�$��`=��on��p��*���)ƿkѿu!οs2��KV�������\�!":�]+��0��7K�i�v��Ζ�`���0Fȿ�ҿ:Ϳ����ٗ��j؃�רR���&����l׾�N���������Z�w���i�I	e�gi�[;v�#����嗾һ���Ӿ�  �  �O�m��|,H��m������ˏÿ�;ڿ���rؿǁ��འ��ـ��N�
�-�u�$�I!3��&X�5���$8����ƿ�1ܿx��8�ֿ1a��?Ҝ��Vw���<��L�a�־V1��C��>)R�Bk2���W�R���O�)�(���B�jFk��v��3���m��''�\�\����n����Ϳ�;߿�1�Rҿy涿�?��s�o�߻A���(���'��=��yi�R����G���Ͽl,࿉� �Ͽf���J���P�b�R�+�0��aþF���1�o��9F��+�5��f����m"�}6��7V�Cǂ�F)���,־�,���:��
t�h���_����jֿڢ���߿e4̿�>������J�b��{;��v*�M@1��;O�����B��:�����ٿ�[��߿�wʿ��������:FV�T�#�֤���[��ܙ��}�z�Y�0/C���6�\S3��8�;dE�Ѩ\��R������<����0��ɻ!�m2S�j�w���
ɿ�߿�r���ݿm ƿHo�����éY�H�9�jj0��?��Bd�׍��s���LͿ��Z���>ݿAĿ����_w��$�J����k��x���̝��V��n��p[�DZR�|�Q��Y��^i�t��������9�߾�L���7��m��L���ط�g3տ>]�J�}bڿ��C�������Q���8��z7���M��py�L����I����׿P9迣2�-�׿w"������M�r�M<�����'�<\��R���O���9k���Z�'�S���T�S�]�ҳp�ޑ�������p�����`���G����h��n_¿��ܿ���C&��mҿ�g��������n��xG��Z6�o=���Z��_���㥿:ƿ�J߿�꿄��r�Ͽɼ�� $����`��-��%���վ}4��5꒾ʣ��r�i�C�\�[X�+\���h�b�~�!��'^��ڠѾ�  �  kM��d� 3M�dz���ɩ��˿K�⿪뿼	�X�ǿhp��C���%�S�x52�	�(��7��p^�P'���I��@�ο~��.��߿�ĿC<����~�TlA������׾���X�~��N�e.��h��_�����_m$��>� �g�c�����xb��e}*�o~b�<���|
��Bտ/,�0:�Q�ڿ����~e���v�f�F�-�e�+���B���p�:���繿�׿:)鿼鿈�׿����?W����h�Z�/�-��1ľ�ĕ��!l���A��1'����������7��%2�qR����ʀ���U׾�5�?�>��{�C0����¿��޿ķ�-���Կ����G��D-i��A@�~.���5��T������å�~�ǿ^_��r�*q迬!ҿ͔��6��A�[�Nu&������c��䎘���y�'iU��>��2�C@/��3�NA��JX�z�|�폙�uZ��.���d$��8X������G��X�п�k��𿥗�]uͿC"�����&_���=��j4� �C�A�j�mG�������Կ;k뿴�񿣼忦;˿����?%���O�oT�������H4���@����i�7!W�x0N���M���T���d�K�����;i���%ྚ��1;�Ss�0욿�?���,ݿ�M�R򿩟�'�ſvi���t��*�V���<�g�;�j�R�%@�� ���/�����߿�5�1�U�߿ƺ��K����Gy�3�?��A�5��i������*����f�+�V�pmO��hP�ΪY�bQl�ww��&���^ƿ�D �i���K�����럦��Wɿ-忭�}�F>ڿ&���U_���Au�y=L��a:��WA��`�uW���f���;Ϳ��������nP׿����a��2�e�r�0�.L���վ款I�&�|�6�e�ѠX�BET��X�(Hd�ܚz�}������wѾ�  �  �O�m��|,H��m������ˏÿ�;ڿ���rؿǁ��འ��ـ��N�
�-�u�$�I!3��&X�5���$8����ƿ�1ܿx��8�ֿ1a��?Ҝ��Vw���<��L�a�־V1��C��>)R�Bk2���W�R���O�)�(���B�jFk��v��3���m��''�\�\����n����Ϳ�;߿�1�Rҿy涿�?��s�o�߻A���(���'��=��yi�T����G���Ͽp,࿎�&�Ͽm���R���^�b�]�+�&0��aþ=�����o�9F�M�+�C����Y���j"��z6�4V�ł��&���)־+�ܷ:��t�_���S����iֿ���߿�3̿=>��1�����b�t{;��v*�@1�<O�ᣀ��B�����|�ٿ�\��߿�xʿ�������*HV��#�����d^��]ޙ���}�+�Y��0C���6�pS3��8��bE�A�\�.Q����������o-���!�v0S�]�v���	ɿ�߿r���ݿ�ƿ�n������7�Y��9�oj0�	?�xCd�z׍��t��IMͿ��]���?ݿ`Ŀ����rx��'�J�p�	o��{���Ν��X��ln�s[�p\R�0�Q�:Y��_i����������[�߾�L���7��m��L���ط�g3տ>]�J�}bڿ��C�������Q���8��z7���M��py�L����I����׿P9迣2�-�׿w"������M�r�M<�����'�<\��R���O���9k���Z�'�S���T�S�]�ҳp�ޑ�������p�����`���G����h��n_¿��ܿ���C&��mҿ�g��������n��xG��Z6�o=���Z��_���㥿:ƿ�J߿�꿄��r�Ͽɼ�� $����`��-��%���վ}4��5꒾ʣ��r�i�C�\�[X�+\���h�b�~�!��'^��ڠѾ�  �  :l޾)�;��Lo��_���X���¿�IɿF#��ϐ��J*����j���=��q!��F�8'&�\�F�,�v�ۥ���#��jbĿ`Xɿ�����N��9�c�d1�A��M8Ծh-��C↾�`�܌@��&,�ZU!�bx�u&���6��*Q�MEx��������;�����}�L�����Wl������ǿ9�ȿ�󻿱\��%���H[�,3��1�b���/�H�U�K�9��5�����ǿ<�ǿ8���@������Q�Q��"������ þFԚ�R|�DCT��U9�R)��:"�k$�!�/��iD�1d�#�������ԾBS�p�/�ta�\���,��w����˿R�ǿS�z&���񀿞}P��!.�w$��+%���?��ok�3��A��;�¿ѿ̿��ǿ>е��o��A_}�fSH�Aa�l�����¾����x�����g�#�P���C���?���D���R�%�j�r��PM��@�þ�D��&%�hF�GKz�<ۙ�_Ѵ��,ȿ\�ο&�ƿw,���ؖ��}v��oI��6-��*%��+2���R������띿������ʿi�Ͽ�Qƿ�ٰ����Hmq��4?�����'�þܫ��[��|N|�i��T_�}^�9bf�^w�.?���	��E	��z#���N,/�*T]����������I0Ͽ,�п�Ŀ�f��F)��EHk�@C��&-���+���?�?�e�v쌿�;��S���9�Ͽ��Ͽ����d���͌�%Qb�(3������㾷�������$d��5.y��h�@`��Pa��Nk���~�Ք������&�þ�e�$��`=��on��p��*���)ƿkѿu!οs2��KV�������\�!":�]+��0��7K�i�v��Ζ�`���0Fȿ�ҿ:Ϳ����ٗ��j؃�רR���&����l׾�N���������Z�w���i�I	e�gi�[;v�#����嗾һ���Ӿ�  �  �6޾il	�s�*�PS�zL�+3��]䢿pɧ�P��X&��sw���J�w&��e�y���A�P�-�؆T�p��������飿Q�T���L��23v���J��#�����B־}����ԓ��{�>[���D��68��6�@#>��nP���l����T����ľM���
���8��c�lt������uO��+j���Y���ˊ�O�h��x>�l������0��$:�ݾc�lL���������ͦ�h�������_g���<���bM���Ⱦ���K����o�pS���@�ݐ8�	�:��G��^����`Е��c��%�׾-��K#� �I��u�����/�����E
��˙�T~��}6^���6���m��p��.)�ÉL�"yx�DP��3x��7J������J��D�����_��7���ԁ��Qʾ���_�����.(j�%[�QhV�
\�K�k�炾�씾d����˾���e���5�PK^�H ��1����[��iF���ئ�2���0���fV��2��.�����T�T�9���`�� �����t������Z������偿MX�qt1����;;�]�̾����GU��ח���怾bmv� >u�TC~�������������rľ4澠	�ע%���I�N�s�窏�k���fr��Ń��+k��֒�>�x��xN���-�'��
��+�;J�Իs��N��s���<���+㮿/��i���K�w�_9M���(���4��#uƾ-���8������{��%�v�7x��ρ�蠌�vy���ͱ��;yy�	R�9g0���V�����Xz��s������wd��E�������j�M�B���&�h�R=�B�4���W��Ё�<Ǘ�"Ө�u����﬿K4��d��FAj��^A�����F�޾�i���q��Ya��yw��������{��!��	����"�������'��E�۾�  �  <i�g���w��w9�y�V�<�q�
Y���$������Ah��`H�+�'���=����꾱��Q���.�RP�`�n����4r��E����l���P���3������������ž�������;���j���Z�{X���b�Qay�K�����4m���־A���_���K(�QD��Sa� [z�����qۄ��z��-_�I&>��m����	e�3�����#��E:��p[�ȯw�7���䄿|*|��c� G��*���֔��;�ؾ�W��:ͣ�莾 Y|��3e��iZ��]��m��{���E��W����%Ⱦ�O�p�@��Cw4�LNQ��m�K��vV��넿:+v��VX��17��~�%n�U_�������<_*�T1K�N�k�1���y����Ά�#�{���a�сD�/)�����\��@�ݾX�¾M����������,�~��Mx�NG�i������b쬾��ľ+�߾�0���Mr)��oD��a��|�χ�������<ns�A�S��3����BY�kl��	����S;���\�m�{�_�������Ç��Yz��{^�.�A�W�'���������L��ȾY4���U��+�������΋�)y���>���!���þ��۾����+}��� ���8���T���q�[��wҌ������Q���Bo��/N�8n.����N(��d�����+��CJ��vk�F���F��9���&4��=4t��]W��;�RI"��������0ݾ߀ľc�� Z��6d��L����P���������|���ʾע��� ��H���'�J�A��L^�ͦz�����ō�_N��3i����d�"�C���%�^w�����
�/�I�5��HV���v��뇿�䍿�����%��C�k���N��3��*����3��׾��ϫ��a���c��Q����̑��E���L��|Ͻ�g	վ
���  �  T;������iI)���7���D�\�M�PN��kE�g�3�tG�'��|�.2˾8�þ��Ͼ0�쾱'�R�"���8�0�H��wO���L�'�B��65���&�=��'�ۣ�rl�Ծ6���a�����N���_���+׊��X������Rɾ���x��U	�5���]!�8D/���=��I���O��M�ZvA���-�iK�AU����۾b@ȾN$Ǿ��ؾ�����|��+�P?��GL���O�NAJ�ؑ>�,K0�Y:"������	�����B�侥�ʾ� ��C2���T��^���"E���������c���վ����L���������(��I7�3EE�p�O�`�S�F N�(:?�z�)�@y�"���.iܾ&2ϾS�Ծ��쾛�	��=!�]�8��K�{4U�J�U���M��A���2��"%���Ӓ�q��0�ͼѾK���Җ��ID�������3��Ŗ���ǗҾ+�쾦'�6����=�&�?4�	�B���O�ބX�mDY��tP�u?�ĕ(�*d�����'��P�۾��羥��P��p�/���E�`�U�w�\��aZ�L�P���B��4��'���������'�&ؾ�^��o���w��T���e1���	��g�о�)�)��b����}%�T�1���?�cN��Z��@`��]�5�Q�#�=��U&���������,辐����?��{#��;�GbO��g\���_���Z��N�Y�@���2��&��u�8���������Ҿ\���R���.���C��Pm��bC��\ؾ<��������L��)��6��OD�[ER���\���`���Z���K�:�6������	�I������bM�	��G��D,��QC�g�U��_��`��3X�L]K�=��q/��H#�����2��������b;����_L��34���l��uc���N˾_��^c���K��  �  H`!��#&���'��'�r�'�i�'��)&��>!������	��>��hҾ+趾c9��S���J��������پ�N�������5#�6O'�w(���(�)�(�#Y(�kU&��� �r���&��Ĩξ����@����ӡ�'��4¾��ྈ	�F������$�d,(�<)���(�
)��(��&�������U����龻6ʾ�u��u����ڢ��0���ƾ���5������X�R/%���'��(��f(�b(���'�l�$�t�8��{[�W[㾜�ľ�����Ģ��Ҥ�_�_�;��o����7�"��)��+��$,��-,��;,�p^+���'�������
��
��aiɾaq���Z��m�������۾����A7�ӥ���'��j-�)f/���/��/��/�;j.�H0*���!������.'辐�˾����R������ �ʾ�W�p������"��6,�z1��2�,�2�d�2���2�c1� 2,���"�@%����X龭7ξ���6�������վCQ󾕚
�����(���0�P�4��6��26��H6��6��54�V�.�:�$����7f� ��Ӿ�gľS����̾�
�y� ����d!��-��_5�i�8�=�9�0�9��{9�@�8��a6���/���$�b����:꾀kѾ�þ��¾�Ͼ��F��r��J�"��z.�a5�bB8��8���8���8��28��$5���-��7"�������K��4ξ|�¾�ľҕҾ��Q����1p%��B0�ip6�<�8�;99�89� B9��_8���4���,��` �#��/�������̾�þ��ƾ�a׾� � c	�����7(��G2��7�i�9���9�X�9���9�E�8��{4���+�����������'߾?�˾Fľ�Gʾ��ܾJ������_W�@�*��  �  �CN�M��0D���6�b�(�G5��=�>��;���־?T���c����
������!� ��ݪ�o�þ�fݾ�[�����b�s��gd,���:��G��O�r5N��C�N1��������y��ɾN�ž|Ծ ��՟�;S'���<��K��0P�L�JA��H3��%��<�)��w�����eо[ﶾL�������c��i�������^޳�;��������
�:h��#��1�,?��J��wO�aK���=�BL)�F��������־��ƾ�Rɾ��޾t��,����0��|D�o`P�m�R��L���?�"�1�R�#�r~�h�~� �ݮ辯HϾҶ�!�wc���5��|T���c��Uǯ�F�Ǿs�L���%
���܎!���.�(=�J�J��rT���V�9tO��S?��X)�������e߾'Bվ(޾����@���j(��/?��P��Y��X��O��A��v3��&��&����X��D�X�Ӿ�S��E��<R���3���h���&���sľQ�ݾw���Ô�jl�T  �PX,��:�o�H�TKU���\��G\��R���?���(��J�����?�龓�b1���{
��7 ���7��9M�y�[�E�`���\���Q�x�C���5�Ǜ(�O���L��#�U��׾���昮�+㤾nN���쬾U����Ӿ�"�b�O���2�&��e3�zA���O�[�d`���[��uN�d�9�B9"��0��[�����t��������̤'�!	?��lR���]�)�_�EY���L���>���0�@�$���x�$$�-�辯�Ͼ����j����社B���u*���ƾZ�ݾ�����z��m�N���+�~9��mG��U���^�K�`�٭Y��tI�)Z3�A���:��z� �0��<q��c1�l�G�߸X��  �  ���Oⁿ�6p�T�T���7�A1�z�����)ɾv���tΗ�⪄��!l��'Z�JU��d]�uSr�A���*��!����tоX��F���q#�o�>�S'\�Iv�E����1��ת}�� d�GvC��#��		�����$� �j��;�4��+V�L�s�t�����T��I�h��rL�{�/�@Q�H��Q߾����모��㒾}���5h�/-Z��TY�ľe��8~�%Y������\h���۾w��$A�6,�̒H�@e���|��ބ�������u�� Y���7��%�CS�����h�P��� �--A���b��}��F���Ѕ�#|�R�b�S�E��*�q�Ek��d�۾ <���v���]��4�����s�6ik�Z<p�e��O�������@����ԾpK�P��7"���<�T�Y�cu�����$��'d���t��V�75��|��7��9���)�Е�C�2�V�S�#�s������r��.Q���!{���_���B��(��}�:���%6߾�ľ�c��✛�8k���ބ��˂�o��mb��۳���P��x�Ͼ|U�a���o�&1���L���i�������>�����Z�r���R��2�Z��"	�����#�y'��vE�6�f��B���ϋ��؍��1��L�y�w�\�?@�Ӱ&��c����HL⾰�Ⱦ����������������͒���`[��u�ž��޾�c������#�K�<�=�X���u�����L*������<��S�i�1yH��)�z���"���W���0�}	P�v�p�JㅿJ������v�����o���R��7�
��4������پ%���HZ�����#��/b���Q��6×�0量Y¸��cϾЖ龆��A��v,���F�p�c�-��R:��`G���~����`���>��/"������>f�'��G�;�(�\��W|��щ��  �  R���s6��v��.�|���P�	)�����3ܾ󿴾s������gG]��E�K�6��3��9�+8J���d��n���w������=��2�`A[���������Ӥ�,ا������!���'p��D��="�����	��@�[4��e\����Ԙ�⤥�#���ڵ���9���Lo��/D�3U�da����Ͼ�櫾)_��9�v���W���B�&�7��7�(�@��iT��"r�FF��sާ���ʾ����6�Z?���i�����D���t㦿Q���R���ˆ�O�`�+�7��^��i
�Ó����>:A�ppl������'��ڨ�NG������ч���c��:���E���K�ɾK���*)��P{�Ab`��O�gI��eM�U�[���s��,��G�u���|=�Ad���,�mT�\���������̰������_��n]��t7Z��'4�%��HV�.��S1�h�V�����8�����������O���=ރ�q�[���3������V�ʾ3 ��;g��֘��i�s���f���c�E'k��|��7���+���	��dؾ�W����S�?�$�h� ��Dj���ī�,箿9Ħ�~����[�BZT��#2�����L�,�'�k�D�m����d2���������	��م�������T���.����n�56̾ː�������䋾�P��x�w���v�EF���+�����8\���Ⱦ�	뾄��qX*�fsO��.z��ڒ����1��,c����������Nq��H���)�x�����@h/��P��n{������3����������`����\��?�p�`G���#�s^�e��͝¾І�������Ȉ�����x�h�{�"����.��
꠾E����Ծ/���ȫ���6�,T^����������(Ѱ�m5���j��uX��Ed�q�=��G$�3���u"��q:���_�R���{���<���  �  E.ɿ����&𭿧����=l�w�8�C�d�۾(M���&��n�c��GB��4,����O��L&"���0���I��_n��~���n��q��iX�^�C�ly�x�������q%ſaKɿ�̾�d���^����.c�Sn8��G�ԛ��*�HkN�*Q�������4��k�ƿ��ȿ���` ��c����G[��t*�V��si̾ �������
[��`=��{*�|!��j ���(�OH:��lV�(��
*���7ƾ:���� %���T�{0��ɩ��������ǿ�ǿ/2���`��h��L�R�Ȃ-�K"�V��35��p^�.��R���1�2ʿ:�ǿ�˷�~k������2M�y�����u`þ�c��yy����_�U�F��28���2�^6��C�{>Y�A�z�]#��]������o��7;�p�m�m����$���-ĿY'Ϳ�rǿ����g���|�b�L�Fa-�:�!�9b+� I�#7w�����沿uǿU�οF=ǿ�`��55���$w�|lC�(,����\¾uq��򉈾�8p�t�Z��O�zJM���S���c��/}�s���#��<aѾ�`���$��Q����kX�����y̿�\пr	ƿ���qc��k�r��lH�͇/��+��|;��_�=���������G�οwVѿ�Uſ�L��������k���:�X�����¾�O����m}��mj���`�F`�7�h�7z��:���[Y��p�澤���i5�4e�Fh���꪿��¿'Eп?tϿڊ��ѹ��Je���ic��>��+���-�E�D���m������୿�ſ�ѿؖο�d�����>:���:Z���,�~	�(@ݾ���8ٛ��ˈ�,�w�>xh�5b�8�d� \p��Ȃ����0q��
z˾�w���,TE��.x�M���~F���Oɿ�Eҿ�̿���������gV�L�6��K+��4�*+R��������'1���<˿�  �  ��+;ٿ����F��㤀�x9E�$���M߾�������])V�=4�~����X�����#��S;�^a�w����+��K���9OR��D��mꩿ��ȿTݿ���Щտ�㻿>����x�[�G�nC+���%�3q8�4�`�}<������ɣ˿W�޿��xӿ�����j��xZm�O�4�t��;g��z���L��R/��#�(;�֬�m�)J,��IH�1 s��,����ƾk�-�.���e��W��d���S�п^Z�|d߿Xο�,��nn��P�e�Gg;�ǉ&��j)� �C��s��|��BN��XvԿִ�[�߿9Ϳ�^��*ˍ��{\��'��5����¾���	�w�L[Q���8��+� ;&���)��5� K�`�l�o������gs�}��'�F� ��|J����¿�Kۿ0��9&߿5IɿX��)����]��/:�;-���7��{Y��)���]��.ǿ�y޿�+翏�޿mZǿƈ�����P�pp��5�����0��������b��lM�ܹB�s�@���F���U��o��ˊ�}1��� о�����,���_���������aϿa�����e�ܿ�Yÿ�@��&2��1�W��;�v6�5I���q�횕�hX��_Կ|�������ۿ"���*�����}��)E�rb��f��3��Ӗ���`o��]�<T�ۈS��M[��9l��)��Ƨ���\��C羗��?�Sv����뼿��ؿ��ֻ�P]ֿۈ��nȘ�o�v���K�m�6���9���S��R��Y��ɧ���ۿԖ�]�濂�ӿ3鵿�O�� �i�:�4�3���ܾ�c��}I��C���3j��\[�&�U���W�u�b�djw����r����Ⱦ�'���!�7Q���vh���ǿAl���꿸9�OοN��)�r�g�h�C�M�6�O3A�w�b�ɭ���ȫ��[˿����  �  
ꕿ�Ő������f^�o,4�����a׾�����9z�"KC��\���Pv轲l׽�ӽ˲ڽWｅ�	��%��OO�G{��ܮ���k��1>��dh��ᆿ;���$���֎���~�4W�w(0�K��#������D��!�xE��m��ሿ@@�����l����z�֋Q���'��'�;�ƾ\�����i��9�t��X���S��=۽�gڽ��彏�����<�3���b�j���Y�������"�DGL��u��Ƌ�o3��Ԡ���9��#�q�A`I��F$��������0�����-�(T��Z|�ۜ��h2������\T��H~p���F��������64�������e�Dt;�u�#��1�������������!5�g�Z�8"������a2�@��n7��a�����;������������9l�S=D���!���
�[2��W	�J��	A��%i��ㇿ�����:���%���#���Di�?����+:�j���_6����o�;�J�C2�}#�ab�6"����}5*�E&=�^Z��(��(F��c�ɾp� �UX#�B�K��v�r���])���/���������0Nf���?�K� �]?��
��:�R|1�U�U�P^~�A'������=��#ѕ��x���a��8��i��&��η�y���y�N�W�_A�,�3�8-�n�,��t2�Q�>�b�S�g�s�PO������S�/!��3�ޘ\�� �������q��㜿~��j����Y���4��8��w��=�Q�n<��b��p��8���J��Q���쐿�}���S���*�W�/־�[��ˁ��J�m�5�P�K>�xK3��/���0���8��.H��`�������^¾���r����A���k��܉�����F�����p獿2+v�N�S�+��R���ج��x(�/J�+�q��2��(6���  �  _����؋���|���W�n/���	��8Ծ<|����z���E��j ��f����ݽٽ���������(�cGQ�~����a���H�sb��9��Ia�Ws��6��@������tv�0�P��M+�E�#�����%��m����?�cf��X��q0���Ր��Ԉ��r� �K��#�qW���bľ���Q9k���;������ï�h]὘�པ콌��<G�G�6��
d�6����\?�����dxF�f�m�X��������o�����i�zC�������������/%��h(�f�M�UYt��މ�K��l���;х�i.i��5A��=����'���ő���g��S>�W"��h�pS����������-��78�8�\�R���7����JݾU����2�O1[�K���Î�)Ô�c�������'e���>���D������X�7t���;�8Kb������������:���ヿ�b�zR:���(��n������q4r���M��\5��:&�=w�)��"��p-�vf@���\��!��iP��B_Ⱦdh��8�� �F���n�RO���#������5��������_�*�:�����V�a1�"���;-�z:P�M�v�X����u��������N���f�[��3����O���B������F�{�E�Z���D���6��G0�&�/���5�K=B�_W�hv�*
���=��C.޾����/���V��E~�:S���R���ʗ��፿M�z���S��P0�q�����jd
����g�7�X�\�hm���萿�蘿�A���h���=v��5N��6'�T�MZԾ�E��ni����p��T�ncA�Rm6�02��3�� <�IzK�äc�Ã�늝�Rz��o��3��b=��je�F�������nݙ���x����o�޳H�+�'�A�u�����ϟ$���D��k��釿?H���  �  ������|�4�e���E�͹"�d���{̾i�����~�W�M�ڔ*�.��O�����(��g���*�����2��X������Z����ؾ��	�'+��N�r�l�]���$낿;�y���_�"�>�4���$�%j�9x��>�������/���Q���o��^���ӂ�L�w�c]�AB;�b��\��8Ӿ�┖���p���D�1;%�zY�[K�<v��d��
��������!���?�j/j��#��i���\�'c�9�6�o�X��t�;$�������q���T�, 3�C������x����E`��d��k<��S^���y�Z���˂�Xs��\U���2�j��$�澆趾7l����n��H���,�%��n��h�OR���c�)�qB��^e������P���H־�`�ݾ&�׷I��j�=�������3b��Rq�ХQ���/�I�����&�ﾁ���)���w-�r\O�ƻo�����?����׃��p���P�>�-���lY�����q��\lz���W�%�?��U0�l(�"�&�,�+��7��J�(�f�-؆�W����Sžx��&!�L�8��[���z��x���򉿡��(�n�`�M�F*-����#��] ���
�[!�oU@�]\b��0���������T/��}m���K�y�(���	��4߾ ն�y���kg��(e�VO���@�k�9��Z9���?���L��{a� �����!B���Jپ�����$�j G�sNi������`��㉿�@��tre�l�C�L$����� ��[�i��ç*�2KK���l�\胿.኿|��q#���jb�L�?�H���@ �@�о���-򐾟�z�?�^�q�K�b6@�͖;� �=��1F�G�U�0�m�����Ɵ�d����y����0���S���t�â���ȋ��v���{�-�[���9�u� ���2�B6�4���m6�� X��Lx�Cχ��  �  f^�MX��QF��X-������T�ľ"t������`���>���%����ʞ	���������]�+�`�F�H1j�Y�������Ͼ/ ��>��D	4�E�K�5�[��^��U�5/@��S%�>Q
�����Tξ/hɾ��ھ����9*���4��!M�Tp\�_�͌T���?�2�%��i
�a��m��ږ�����|X��|9���"��4�A*�'�
�ڱ�t. �;�5�BpS�[�y��ɕ�?�����ݾ�X�!�iy<��R�@�]���\���N�pL7����r�"�ݾRfʾ�c;2�4��I�#�\?���U�oSa���_��Q�h�:�ϕ�e�	�۾�V���>��d��\���@��-�O�!�+/�[ �5+��3=���V�L�w��u���鬾��ϾZ�����<2�o�K�q�^�"|f���`�-kO��	6�Ԕ�����侙�ؾ���0����4���N�-�a��i���b��2Q��A8����Y���ھ�j��⿛�G_���	l��S�b�B�|19�N7�� =�`7J�D�^�*�z�i���*Ц���ľ�,꾿��r&�2�A���Y�j`i���l��\c���N��M4�+��Z������N���$�h�)��XE�v�]���l�ғo��	e�%;P�r�5�������ھ�ֹ�`������]y��nb�8�R���J��:J�GQ���_���u�H��������浾��վZ��F��=2��L�_|b�Zn��Cm�D_�-�G�J2,��X������p���쾄�������2���M���c�^�n�{m�i�^�p�G��,���k���%Ͼs찾�f��)8����r���^�ǶQ��cL�&�N��hX�֛i�����`����������h�0���.!��}<�V���h�иp��+k�b�Y�@��n$�PN�?�������~��</
�Y�!�V==�"UW�1j��  �  �5�l�1�:�%�����r⾒�þ_!���+���$���Ba���E�	{0� �#������%�5��L�Ui�\߅���������o˾A(�_z�c��P�)��4��5���-����J	����x�ƾ���~A��a����Xؾ�v��'��J�'�us3��96�x�/�B�!�4������ھ�������t�����z�#M[��uA���.�	�$� �#�$�,���>�ǆW�W@v�R���2���2r���վ5������{�b�-��W5�y�3�N�(��������۾E�� D�������-ž��澳B�w�L�.��8���7��.�%d��?������~־�@��h@�� �����~���a��;K��;<�,N6��	:��,G�"�\�D�x��+���b���b���о|?x����R,�Ԗ8�D=�u8���*�*��8��p"�)�ƾ�����ž6@޾�~�1��&�*���9���?�-^<��0�� �ܞ��O��U�پ;��bI��Fy��+>���zs�%_�PS�rPP��@W��Rg��3�z���w8���K��me˾�}�A'�{��{'�@�7���A�b�C���;�9,�1����H��:�ѾrBξ�ܾ=����#�Ah%��8�(�C�+�F�|&@�6R2��� �|/������yݾ��ľ�Ư��k��3��������]n��.d��c��zl�]4~�֞�����F������d�پ����������/��?>���E��D�] 9�D$'�j�aO��xK޾ϾѾ"��]a���*�+��<���E�!*E��;�*n,�k;�{=�&\�>
վ`罾��������
ԉ��,|�_Yl�ӊe�~]h�`�t�3����8��혢��z��f8˾Z��jg�X���5%�_6�N�B��G���B�l5���!��d����fھԉо�Wؾ�X�7Y
��y�Om3�p�A��  �  �(��|�
��g�pk�D��Y о�̿�7����(���	��It���X�aOG��IB�B�J���^��E|�G����衾�����mľ6�Ծt�徲���(����+I�qQ�GP	�$<���۾�k��~h��:��
e���`��&���yWξ���߮�s=��������X	��� �y��GIݾ��̾}���?��� ���!��V�m��?U�QG���F��R��Zj��鄾����
ƨ�@��6Zʾ�ھ���N��������g�fg����'-ѾK&���O���u��?q������漾��۾�Z����
�	�����{�#�	��� �Uﾱf޾CξAܽ�������du��ѝu�e8a���X�$d]�j�n��<��vs�����%r����̾�Yݾ)������B	� ��v��q�������i-���a־�O���Ө�����G��cr���վ� ��~�	�"����������Y��'����?����վOž�}��p����������v��r��{�d������y��;)���>ξ�B߾���pn �ܐ	����ʨ���<Q�Y��q��ɍ��ϱ۾�Eþ?���=��ޗ���Ҿ�ﾚ:��+�c��Ip"�!M �k�����Ư�����=��ܾ�^˾)%��s��qؖ�bq���������N:��R����ä�՝����Ⱦ`ھ>������ �U�F=�����!�D����4g�>��{Ծ5U����� ���|�¾��ھU ��,����SK ��!��7�������/���<�����x׾,�žbʳ�DF���B��z���[����兾�$�������U��ތ��\�оf��C�Z�C
�L��Y��!�v�"���6�E����ּξf컾ش�����yp̾�:��(����a;��  �  ��#�'��/��$�����զ澀Pپ�gƾ��������u���m��jy��Ɗ��ើ}���ͺ˾��ݾ��)?𾑯�:?�9��H�O��uD���׾&9ľv�������;���u9u�,q����K��WУ�S����9оx<�sS���y��>��g��s��w{����վM:���^������2����s�]�r������A��a���l\���!Ӿ������l �A�f��1���O��LwѾ�����إ����g��^zs���v�3��%��^����CƾH1۾���|�������l��.���?w�����y��֨��־Ia��7᪾mƖ��h��6��H���/���	���Ϻ��Ѿ���P<������o' �� �X� ��{ �������������پ=ľθ��;W���.���z��,��K�����Mž��۾��V������p�,�����
��������zq��ܾ��ƾ+�������.�����`*��䨣�*2��{{Ͼ+�徐"���D�����5�^>� ���%����N��P%��˾����i4���ә�jD��Mܟ��k���sľ��۾�&�s�$���n	��]
��
�%]
���	�Tl�?��6���+=�!LʾI����f���ř�Q3���š�����bǾ/D޾��ڒ�����	�$�	�3�	���	�����o��@�i-�,%ݾ$Dƾ�$��t9��K"��T7��hL�����0�˾x}������������	�F:
��S
��(
�?(	�/E�� �;�ﾥuھʥþE2��Hu��;ޙ�V���{���m����о�r���������w
�2�
�<���
���	�3B�j �� ؾ�v������u?���+��#a��i0��L���*־H��7U���  �  �1��^�о�Y��^�K����-�V0��.
��x��y�߾����9���堕�ɫ��똘�"��e Ⱦ�A����w�n2�' ��!
�Š�c���6߾��ξ�y���w�������t��p�q�#�W� /H�SE�ҡO��e�� ���ԓ�}��a����>ȾŒؾ۵�r�����i�;�����������EC׾�@�������7���t���`�����/~Ӿq�}�e�7��	��o�����x�꾂`پ5ɾ����E��(?��^���˸h��}R�y�G��wJ�PZ�I�t��[������ܰ���¾BxӾ"K侴���]��!���@j�<�����8�� վ4򸾱Ĥ�)�����S���Oʾ�|�k�I��,�l��u����э���R�}.Ҿ����}"��|8��J���u~���k��ie�Gl�1���L��#ܟ�v���ѻľA�վ�c�@H��ɨ�l�����#�'0��@���	�B_��\�׾w罾B9��a���P�	�ľ�(�Tj �u���ς�*m�����0��������U�Ydھ��ɾ�U��զ�\▾�h���$��q0�������������񑴾��ƾ%�ؾ�1�F}���F�-a�Aa�u���"�z �$���h/���پ.[������:��'���վ�T�N+	�Pz����!�F��_��������c���龟Eپ�Ǿ𺵾����S[������ ���䃾�������w���-���P̾�ݾ]��|��{	��M���W] �\:"��=�mp�Zl�N��ySѾμ�I���K���9Ǿ%������A��f��2�!��`"�V����w�����������H־@jľB�����%���]��X��{^��P��������ڰ��#þվ�  �  Q��"žF�=��� ���&�}$2��C5�C�.��������lʾ����b���	��pѾIG�����s2$��}1�H�5���0�W$�q��Zc ��v޾���������6���4�B�^�mCD�^a0�7�$��"��i*���:��S��q�3#��U���ĵ��pѾ��V�(:�[w,�{W5�E5�`�+����(�����ґ¾����j��� ����a޾�>�A���)�(a4��x5��p-�o��3������~�Ӿɥ���������A�s�r�U�b�=�.-���%��'�H�3�t/H�U�c��p��w��2+���Uľ��ᾤ�C��)&�̶3���9���6��x*�!��3��CH߾�þ����/���7�Ҿ����B���$���4��W<�}r:���/����B�����jGؾ|ɽ�r_��s���g���j��,U���G��*C��tH��W��m�Hb��=���)��P���4۾���D���!��1�=�"E@���9��+�:2�WY�^W�j�ʾ�Aľ'BϾy��!�P���1��>��#C��.>�I1�-Q ���������Sܾf�þ�{��X���Ì�O��m$m���b��a��	j��C{��􉾰6�����9��+�־7U�]	�fk���-�k�<�]�E�j`E���;�U�*�����F��`�8aо�[Ͼ|t߾�,��&)��2(�
�9�hD��E���=�_�.�H��}�
�lp���Kؾ�~������?��^���@N}��	l�b�c���d�yno��S���s���a��Ұ��ƾz�޾������o!�=3���@��F�JfC��7�rE$��������۾�lϾzVԾB���?�'��/�_P?�T�F��D�,W:��1*�Y��W����R^Ҿ׻��^���q��p ��@�{���m��[h���l�'�z�(��MN�����m���  �  2���#�ƾeQ���%�.���G���X�"�^���V��C�I)�������Ͼ�`Ǿ�վ$����O�/���H��#Z�_�\�V��AC���)�R[��e�%ڿ�"���9��y�\���<���$�Y`�@�-�	��������1��HN�;bs����b���7׾B5�U����8���O�Pq]�Y�^�=�R�"L<�/� �Pr�Dg�^S̾�
˾��߾o�����89��MP���]���]�JYQ��@;�d| ����۾�[��`ᓾ��v�CQ�}4�ݪ��V�Х�ܦ��Q�z�)�%B��fb�J���s���bI¾�K�L��[*���D���X���b��_�N�O��m7�_��? ��n��Ҿdپ�Z��\G���,�ۤG�PF\�6�e��a���Q���9��g��E��<۾�q��ꐙ��6��%d��^J��#8�bY-��"*��.�Om:���M��Uh�*���~曾�x��\�ܾ)��]���9�r�R�Y�c� �i�<�a��N���4�`��l��{�m*߾� �q���n �S<��U�O%g�Y2l��c���P�77����5��Xf۾�����D�����31w�j``���P���H��9H��O�C]���r� ����s��ր���EѾ���̜��?.��#I�'�_���m�_�n���b�)KL���0�_��������~��P����-�G)I��G`��m���m��ya�oK�Y�0�/�� ���9�Ӿp���ܛ�׈�]�t�P_���P�0YJ�pFK�9�S���c��z��
��ZF���X��5�ܾ3�U�'=7�ZaQ���e�v�o�Il�#h\��C�_/(��#�un��؁����G4����~�7�/�R�b g��Cp�|+l��\���C�ͺ(����@�ﾛ˾	��������M�q���^�FNS�0AO���R���]�=p�]	��\�� ���  �  �3��m�ξ���L�$���G���g���}�Ă��|��2d���C�rQ"��C�ǯ�]J޾4�����X�)���K�\�j�6��邿!�z���a���@�����d����ž����[5x���I�^�(��]�j=��l��o���'��s+
����p:�b�b�k��ei�����\d�}1�RT��q����������v��[�]f9�J�������0b⾑X��ٮ��z5�WAW�+�s����`��5�s��SW�W�4���辒W������u�f��=�Bv ������ ����������zK���-�_O�zs}�f읾�9Ǿ*������@�;b��|�r΄�	񂿠]r�T��O2���������龄���	�y%�ezF���g�대�8J����� 9r�|(S�J0����a���������P�t�P��s6�!�%�y�^i�[[��(��9��6T�?y��ڕ�����;�����<�/��R��r��z��:F��M����eo�F%O�i�-���� ����2^���X6�N1X�;�w��}���w�������o��N��K+�	X��P�撷��K��k�����b���L��>�/�7��>7��V=�.J��j^���{����*��FӾ���-����A�cd�|ဿщ�j����M�� k��ZI���(�Z�����b���A�%��cE�>1g�xみ����"��4����g��+E�Y�"�<U���־�}���ٓ�~�3``�L�OI?�9��O:�+�A�xGP��f��t����ǫ��H��z�[�*�gjM��o����<$���;����~��z`�j�>� �a\
��� ���H3�d0�D�Q�o�r�dl����ƈ�Ι|��]��:�pC��)��^V˾�q��橎�qx�Z�]�DL�.�A�tz>���A��ZK��j\���u�Q��c���  �  0b��׾����1���Y�b�~�{u���ې�}u��i}{���V�ԃ0�����p��A��� ��2���8�Zk_�F���ǯ������遊�_�w�^�Q�i�)����Hi̾�圾ps�A��=�v���g�=��޽���m����E���0�+�[�(y��W��h�����@@�o5h�"&��	���
���G2��e�p���J�`�%�Z�	�w���)���""�KF�i�l�E������r��烆�?l�cQD�B��Y��u��Ə�ݘ`�T=4���X��9��F��轌i�����>�#��|F�[+x�%���(;|���(��$Q��x�+K���ڒ�غ��X����nh���A�,���S�ZO����U�� �2�ɡX��i~�nʍ�^\���$������f���=����n�}�����m�F�U�+�n[��`��������9w/�T%J�?q�����0����ܪ���<���d��턿�X^������X����a�L�;��t�o�����P#�P&E�^�k�R߇�� ��l�����������8_�
 7��o����,����䕾IVz�nX��B�H}4���-���-��n3��?�W�S���q�ѥ���F���0׾�+��k)���P�Fx��B���������G7��/i���Z���5��y���	����C���2�V�́|�M��������P����.|�o�T���,�L
��w۾�A�������t���U���A��k5���/���0���7�Z�E��O\���}�mF��U���~�ǣ���5�&�]�i�����W,��� ��������t�
.N��+�dO�
�����6{��!>� �c�ڳ���.��ʩ���`��79���rp�c3H�-�!�
�vξ�	��ӊ�x"n�MYS�ZB��D8�v�4���7�!3A�m�Q���k������L���  �  ,����Qھs��t6���`�����h��B���\��j���)L]���5����b���=��5��<��P>�Ĕf���1���l$��pX�����qX��.����k,Ͼ���|r���>�,�Д����V۽��ؽ�@�V&�����-�%.Z�����$��'��A���E�_�o�W�������.ϕ��錿�x�ʼP��*���ʊ������u
�I�&�8L��Pt�G���)��;��(&����s�pJ��� �5����������_���1�2��f������>C߽��⽱�̲�� ���C��w��>����Ͼ0��5-�wHW�Q��u�����AǕ�L����o��G�8�#�ނ
�����}�������7�)3_��Z�����ʅ���#��Pk���m�
�B�������޺�+v���k�� C���(�r��F����ף�1���/,�p G���n�1ߓ��]��AB�u��^tA�[�k��:�� 斿�����蕿����3�h��A��= ��f�`s�$+�6W'��J�B
s��F��&����������Ȇ�בe���;��+��꾚���j����w�fIU�v�>�CB1���*��*�C0�=x<�ϋP�w�n��ƍ�\m��,�ؾ�A	��-��V�����Б�����۝��r`����`�m:�������{���V�J}6��\�����B���*���&��R4���灿�;Z�v�0�gL��~ݾx����᏾��q�8�R��Y>�D2���,�>�-���4�3�B��$Y�	g{�>���2���� ��4��:��d�-m��<l���R������<���|��S���/�~�)E�l��`&#��C��ij��ڈ�R���Ӟ�K`��ǜ��@rw�nBM��%����|sϾ�릾�͉��*k�RP��>�{(5���1���4�h�=�E�N�Ͽh�=懾a���  �  0b��׾����1���Y�b�~�{u���ې�}u��i}{���V�ԃ0�����p��A��� ��2���8�Zk_�F���ǯ������遊�_�w�^�Q�i�)����Hi̾�圾ps�A��=�v���g�=��޽���m����E���0�+�[�(y��W��h�����@@�o5h�"&��	������G2��e�p���J�a�%�[�	�y���)���""�NF�l�l�G������w��탆�Nl�rQD�P��q����Ə�ɘ`�=4�w��~��7�3D�i���d�������#��xF�)&x�)����$;����(��"Q��
x�-J���ْ���������mh��A����`S�5O�������޺2�ϢX�&k~�7ˍ�D]���%������f���=�Ն�"r�Հ��ʕ���m��F��+�I]��a����"��Y���t/��!J��q�����-���������<���d��섿��f]����HX��s�a�v�;�ct��n�"��R�{Q#�2'E���k�����!��g����������.;_�*"7��q����|����畾J[z�=rX�wB� �4�8�-���-�p3��?�#�S��q�����F���0׾�+��k)���P�Gx��B���������G7��/i���Z���5��y���	����C���2�V�́|�M��������P����.|�o�T���,�L
��w۾�A�������t���U���A��k5���/���0���7�Z�E��O\���}�mF��U���~�ǣ���5�&�]�i�����W,��� ��������t�
.N��+�dO�
�����6{��!>� �c�ڳ���.��ʩ���`��79���rp�c3H�-�!�
�vξ�	��ӊ�x"n�MYS�ZB��D8�v�4���7�!3A�m�Q���k������L���  �  �3��m�ξ���L�$���G���g���}�Ă��|��2d���C�rQ"��C�ǯ�]J޾4�����X�)���K�\�j�6��邿!�z���a���@�����d����ž����[5x���I�^�(��]�j=��l��o���'��s+
����p:�b�b�k��ei�����\d�}1�RT��q����������v��[�]f9�K�������4b⾗X��ݮ��z5�_AW�6�s����j��M�s��SW�t�4����農W������O�f���=�iu ������ �\��t���P���E�p�-�|VO�ei}��松q3Ǿ���F��,�@�7b�B�|��̄�u�Zr��T�%N2��������q��C���	��%�X|F��g�i����K��􍃿�<r�z,S�N0�I��;��6ƶ����<�t�4P��x6���%�Y��i��Y�3(���9��/T�zy�KՕ�p���T��5��=�/���R��{r��x��mD�������bo�!#O���-� ��l �����^���6��3X�	�w�W��by�������o�N��O+��[��W�R����Q��H����b�S�L���>���7�fB7��Y=�0J�Bl^��{�^��p�$GӾ���4����A�cd�|ဿщ�j����M�� k��ZI���(�Z�����b���B�%��cE�?1g�xみ����"��4����g��+E�Y�"�<U���־�}���ٓ�~�3``�L�OI?�9��O:�+�A�xGP��f��t����ǫ��H��z�[�*�gjM��o����<$���;����~��z`�j�>� �a\
��� ���H3�d0�D�Q�o�r�dl����ƈ�Ι|��]��:�pC��)��^V˾�q��橎�qx�Z�]�DL�.�A�tz>���A��ZK��j\���u�Q��c���  �  2���#�ƾeQ���%�.���G���X�"�^���V��C�I)�������Ͼ�`Ǿ�վ$����O�/���H��#Z�_�\�V��AC���)�R[��e�%ڿ�"���9��y�\���<���$�Z`�@�.�	��������1��HN�;bs����b���7׾B5�U����8���O�Pq]�Y�^�=�R�#L<�0� �Rr�Gg�cS̾�
˾¹߾t�����89�NP��]���]�jYQ��@;��| ����۾�[��pᓾs�v��Q��{4����8T���͡�UK�8y)��B��Zb����5���+@¾�A���$V*�H�D���X���b���_���O�{j7�������l⾺�Ҿeپ=]��QI�p�,�I�G�oJ\��e�L�a��Q���9�m�'K��F۾Uz������5=��X/d��fJ��(8�\-��"*���.��h:�e�M��Kh�懅��ޛ��o����ܾՠ����U�9�řR���c��i���a�.�N���4��]��k� z羅*߾�"�����p �*V<�^�U��)g��7l���c�^�P�7�������{p۾Ϟ���L���
���<w� j`���P���H��>H�TO��E]���r�龇�It��6���
FѾ��֜��?.�$I�'�_���m�`�n���b�*KL���0�_��������~��P����-�G)I��G`��m���m��ya�oK�Y�0�/�� ���9�Ӿp���ܛ�׈�]�t�P_���P�0YJ�pFK�9�S���c��z��
��ZF���X��5�ܾ3�U�'=7�ZaQ���e�v�o�Il�#h\��C�_/(��#�un��؁����G4����~�7�/�R�b g��Cp�|+l��\���C�ͺ(����@�ﾛ˾	��������M�q���^�FNS�0AO���R���]�=p�]	��\�� ���  �  Q��"žF�=��� ���&�}$2��C5�C�.��������lʾ����b���	��pѾIG�����s2$��}1�H�5���0�W$�q��Zc ��v޾���������6���4�B�^�mCD�^a0�7�$��"��i*���:��S��q�3#��U���ĵ��pѾ��W�(:�\w,�{W5�E5�a�+����)�����֑¾ ���r���+����a޾�>�A���)�?a4��x5�q-����c��K�����Ӿ�������􃋾{�s���U��=��-�P�%���'�-�3�7%H���c�?i��4n�� !��\Jľ���%����"&�|�3���9�Y�6��t*����s��yD߾�þ����h���!�ҾZ���w�ҽ$���4�P]<��x:��0�����������gSؾLԽ��h��a���m����j�\3U���G��*C��qH�� W�Ѣm�\��r����������ھ����k���!�B�1�=�1?@���9�!+��.��V��S�ŞʾBľDϾ&꾰$����1���>��)C��5>�R�1�SX ���C���w`ܾ��þ󅮾�`���ʌ�`��7.m�g�b�#�a��j�^G{������7����\:��s�־aU��]	�kk���-�l�<�^�E�l`E���;�V�*�����F��`�9aо�[Ͼ}t߾�,��&)��2(�
�9�hD��E���=�_�.�H��}�
�lp���Kؾ�~������?��^���@N}��	l�b�c���d�yno��S���s���a��Ұ��ƾz�޾������o!�=3���@��F�JfC��7�rE$��������۾�lϾzVԾB���?�'��/�_P?�T�F��D�,W:��1*�Y��W����R^Ҿ׻��^���q��p ��@�{���m��[h���l�'�z�(��MN�����m���  �  �1��^�о�Y��^�K����-�V0��.
��x��y�߾����9���堕�ɫ��똘�"��e Ⱦ�A����w�n2�' ��!
�Š�c���6߾��ξ�y���w�������t��q�q�#�W� /H�SE�ҡO��e�� ���ԓ�}��a����>Ⱦƒؾ۵�r�����i�;�����������HC׾�@�������7��u���`�����C~Ӿ+q��}��X��2����������`پyɾ�����D���>������7�h�-zR�6�G��pJ�(Z���t��T�����Ұ���¾okӾK=�6��zV���y��c��{� ��k���Ծk¤���Z ��!W���Tʾ~����`N��2�3�������F��k'�_⾽:ҾF����+���?���O��#}~�]�k�je��Cl�m��}G��՟��y��.�ľ �վ�U澜9��*�����;
����)�;��	��W����׾�㽾{7�����W��ľ�.�On �m�����|t�t���8���ӧ���c�1qھ��ɾ�_��Xݦ�6閾jn��)���3��kÇ�������������ƾ��ؾ2�o}���F�2a�Ca�w���"�| �%���i/���پ.[������:��'���վ�T�N+	�Pz����!�F��_��������c���龟Eپ�Ǿ𺵾����S[������ ���䃾�������w���-���P̾�ݾ]��|��{	��M���W] �\:"��=�mp�Zl�N��ySѾμ�I���K���9Ǿ%������A��f��2�!��`"�V����w�����������H־@jľB�����%���]��X��{^��P��������ڰ��#þվ�  �  ��#�'��/��$�����զ澀Pپ�gƾ��������u���m��jy��Ɗ��ើ}���ͺ˾��ݾ��)?𾑯�:?�9��H�O��uD���׾&9ľv�������;���u9u�,q����K��WУ�S����9оx<�sS���y��>��h��t��x{����վO:���^������7���+�s�o�r�����B��v����\���!Ӿ��>�U��� �B�����1�>�p��1wѾ����ץ�����e���ts�&�v�d���
��Ю���:ƾ�&۾��꾔n��W����]������fh���w�����x��`�־sY��=۪�N�pf���5��sI��3������ֺ���Ѿ��徭H��^����. ��� �� �� ���������뾠�پ� ľ����$[���0���z��{��}G��`����ž5�۾T���I�����4i�F�����a{�������fﾌ�ܾ�ƾ����<���,�����j,��ᬣ�%8��y�Ͼ$��j.���K�R����-=��F����:-�g#��Z���/��#˾Т��B:��tؙ�H��ߟ��m��;uľɒ۾D'��H���n	��]
� �
�(]
���	�Vl�A��9���.=�#LʾJ����f���ř�R3���š�����bǾ/D޾��ڒ�����	�$�	�3�	���	�����o��@�i-�,%ݾ$Dƾ�$��t9��K"��T7��hL�����0�˾x}������������	�F:
��S
��(
�?(	�/E�� �;�ﾥuھʥþE2��Hu��;ޙ�V���{���m����о�r���������w
�2�
�<���
���	�3B�j �� ؾ�v������u?���+��#a��i0��L���*־H��7U���  �  �(��|�
��g�pk�D��Y о�̿�7����(���	��It���X�aOG��IB�B�J���^��E|�G����衾�����mľ6�Ծt�徲���(����+I�qQ�GP	�$<���۾�k��~h��:��
e���`��&���yWξ���߮�s=��������X	��� �y��HIݾ��̾ }���?��� ���!��^�m��?U�]G�ϬF�2�R��Zj� ꄾ���.ƨ�p��sZʾN�ھ��뾰�������+g�xg��p�`,Ѿ%���M���r���m�����༾V�۾�Q��=�
�����f�ѳ	�,� ��F�LY޾�6ξ�ѽ����������o���u�4a���X��f]�f�n�A��z�����<|��i�̾�fݾO+�� �J	�}��}�5x�f��q��5��ag־tS���ը�����E���n��h�վ(��͋	�������������SR� �q����得�վ�ž�t��H������=�����v�B�r���{��g����������2���Iξ`O߾"��v ���	�������F#��W�V�����������۾EKþɢ���@�������Ҿ�;�M,����hp"�2M �t�����ɯ�����=��ܾ�^˾+%��u��rؖ�cq���������N:��R����ä�՝����Ⱦaھ>������ �U�F=�����!�D����4g�>��{Ծ5U����� ���|�¾��ھU ��,����SK ��!��7�������/���<�����x׾,�žbʳ�DF���B��z���[����兾�$�������U��ތ��\�оf��C�Z�C
�L��Y��!�v�"���6�E����ּξf컾ش�����yp̾�:��(����a;��  �  �5�l�1�:�%�����r⾒�þ_!���+���$���Ba���E�	{0� �#������%�5��L�Ui�\߅���������o˾A(�_z�c��P�)��4��5���-����J	����x�ƾ���~A��a����Xؾ�v��'��J�'�us3��96�x�/�B�!�4������ھ�����u�����z�(M[�vA���.��$��#�8�,��>��W��@v�q���[���gr��U�վ����9���{���-��W5���3�H�(�Y�������۾����A��F���k)ž2��C?��r�m�.�-�7���7���.��]�.9������r־�5���6��|����~���a��4K�.8<�bM6��:�B2G��\���x��2��zk���l���оL�S�S��,�9�8��I=��z8��*������	&��ƾ;��� �ž�<޾|������*�ҫ9���?��W<��0�������B��9�پ]���?��eq���7��[qs��_�\	S��PP��CW�-Yg��=�����@���U���p˾R��	.����'�O�7�c�A���C�<�;�#,�7��:�����]�Ѿ�Eξ�ܾ���7$��h%�18�U�C�E�F��&@�=R2��� �/������yݾ��ľ�Ư��k��5��������]n��.d��c��zl�^4~�֞�����F������d�پ����������/��?>���E��D�] 9�D$'�j�aO��xK޾ϾѾ"��]a���*�+��<���E�!*E��;�*n,�k;�{=�&\�>
վ`罾��������
ԉ��,|�_Yl�ӊe�~]h�`�t�3����8��혢��z��f8˾Z��jg�X���5%�_6�N�B��G���B�l5���!��d����fھԉо�Wؾ�X�7Y
��y�Om3�p�A��  �  f^�MX��QF��X-������T�ľ"t������`���>���%����ʞ	���������]�+�`�F�H1j�Y�������Ͼ/ ��>��D	4�E�K�5�[��^��U�5/@��S%�>Q
�����Tξ/hɾ��ھ����9*���4��!M�Tp\�_�͌T���?�2�%��i
�a��m��ۖ�����X��|9��"��4�K*�3�
����. �X�5�hpS���y��ɕ�i���Ŀݾ+�z�!��y<��R�\�]���\���N�PL7��������ݾWdʾ�`;x.���j�#��X?��U��Na���_���Q��:�e��4�a۾�M��_7�������[��@���-�E�!��.�G] �n+��:=���V�x��|��G���Ͼ���~��MB2���K�ư^��f�a��nO��6������T�侼�ؾy���������4�
�N���a��i���b�8-Q��;8�a��cT���ھ(b��J����X����k�x�S�z�B�/9�4N7�9=��<J�-�^���z����ئ���ľ 7�G�^x&�!�A���Y�fi��m��ac���N��P4������P��D���%��)�)YE���]���l��o��	e�+;P�v�5������ھ�ֹ�d������]y��nb�:�R���J��:J�GQ���_���u�H��������浾��վZ��F��=2��L�_|b�Zn��Cm�D_�-�G�J2,��X������p���쾄�������2���M���c�^�n�{m�i�^�p�G��,���k���%Ͼs찾�f��)8����r���^�ǶQ��cL�&�N��hX�֛i�����`����������h�0���.!��}<�V���h�иp��+k�b�Y�@��n$�PN�?�������~��</
�Y�!�V==�"UW�1j��  �  ������|�4�e���E�͹"�d���{̾i�����~�W�M�ڔ*�.��O�����(��g���*�����2��X������Z����ؾ��	�'+��N�r�l�]���$낿;�y���_�"�>�4���$�%j�9x��>�������/���Q���o��^���ӂ�L�w�d]�AB;�b��\��8Ӿ�┖���p���D�4;%�~Y�`K�Iv��u��!��������!���?��/j��#������\�<c�Q�6���X�.�t�F$�����~�q�o�T��3������Zw�����^��b��i<�8Q^���y��	���ɂ�s��XU�̻2����V��fⶾ�f���n�sH�@�,�T��O�;h��S�	���)��wB��fe��Ɗ��V��uO־Rd���&�ջI��j�)���d����c��q���Q�P�/�b����?�ﾎ���(��'v-�XZO�!�o����v����Ճ�p�p���P�B�-�C���R�򀶾yl���cz���W���?�.R0��(�?�&��+���7���J���f��܆�䈡��Yž���%�p�8��[���z�{����O���n���M�C,-�����$��^ �n�
��[!��U@��\b��0���������W/��}m���K�{�(���	��4߾ն�{���mg��+e�WO���@�l�9��Z9���?���L��{a� �����!B���Jپ�����$�j G�sNi������`��㉿�@��tre�l�C�L$����� ��[�i��ç*�2KK���l�\胿.኿|��q#���jb�L�?�H���@ �@�о���-򐾟�z�?�^�q�K�b6@�͖;� �=��1F�G�U�0�m�����Ɵ�d����y����0���S���t�â���ȋ��v���{�-�[���9�u� ���2�B6�4���m6�� X��Lx�Cχ��  �  _����؋���|���W�n/���	��8Ծ<|����z���E��j ��f����ݽٽ���������(�cGQ�~����a���H�sb��9��Ia�Ws��6��@������tv�0�P��M+�E�#�����%��m����?�cf��X��q0���Ր��Ԉ��r� �K��#�qW���bľ���R9k���;������ȯ�o]ὡ�འ코��GG�U�6��
d�B����n?�����qxF�s�m�_����� ���o�����i��yC�b��B���������$��g(�Q�M�Xt��݉�j��w���9Ѕ�^,i��3A�<����������c�g��O>�,T"��f�YR�������h��J0�;8�v�\�獈�<��� Nݾ6����2�d3[�V���Ď�Ĕ�8���Á���(e���>�����������X��s���;�Jb�����������9���⃿ėb�hP:�����꾸k������/r�Y�M�EZ5�69&�ev�)��"��r-�Ki@���\��#��ES���bȾl��@��(�F���n�mP���$������6��b����_�4�:�� �aW��1�~���;-��:P�m�v�b����u��������O���h�[��3����Q���B������H�{�F�Z���D���6��G0�&�/���5�K=B�_W�hv�*
���=��C.޾����/���V��E~�:S���R���ʗ��፿M�z���S��P0�q�����jd
����g�7�X�\�hm���萿�蘿�A���h���=v��5N��6'�T�MZԾ�E��ni����p��T�ncA�Rm6�02��3�� <�IzK�äc�Ã�늝�Rz��o��3��b=��je�F�������nݙ���x����o�޳H�+�'�A�u�����ϟ$���D��k��釿?H���  �  ��<�B67��9'�q��0v�~˽�م��h�b��.�� 	��Aݽ���S좽�Ӗ��ȓ��S��d,�������� ���:���r��a��Muɾ�,��)��	Z,�$c:�r�=��{5���#�@����0�ž�خ����s����پ,���?��.��;�ĥ=��'4�}t!�Yi	��(�W5��.���%VT�U=%��V��׽�^����������#��2�������~ҽ/��� �<UM����6�����پ�&�c�P�1�t�<�?<��I0�b������ݾVI��ҭ���P���þ��I��ds#�ET6� @�r>��1�����!�_f־���u􄾩Q�J%'�f�	�Լ�ҙҽ[�Ľ����^-Ž��ҽ9V��U�U�!��(G�B3z�;����:Ⱦ��������,�.�=��E��@�*�1��Z����?i�N?ľ�ٹ�?�¾��ݾ�i��-���1���A���G�"�A��2��[�����Ӿ�a��,l��*<[���5����!�
��2 ��������<!���e��-���(���F�T0p��%��g^�����*�VV$��:��7H�S�K��C�Hj2�G��a��\�侈:ξ�WʾZ�پ*��������*��.?�OL���M��xD��1����]D ��xѾ-���w4��e��C�P`+������(�[�����q��C�(��?�D�_�Ȗ��.
��h�˾R���U���.�BB���L�ZXL���@���,��*�����ugܾ�w˾��;;��ڧ�1��y�1�GQD���M��K�H�>�\�)���\E���þ秞����	�Y���;��e'�w�3]�Ta�?�����
v!���2��|L�i9q�nᑾ�)��6�ܾ�~�3���,7��-H�NJO���J�*�;� M&������n׾��̾Cuվ�8�.e�<�#��,:�UJ��  �  #-7�o�1��Z"���t��5,��)�����a�e�/���
�����E������?��# ��dʝ��׬��ƽ
��Kf��5;��p�)!��hžu������K'��4���7�
0��q	���l�����^妾�V���'Ծ�9��J��&�)���5�-�7���.������^5۾93��D����S�"D&��>��Eܽn��d���� ������㺧�����] ׽N��Y-!��M������ᨾ�&վM���	�M�,�p�6��D6��+�{���V��ؾ� ��Z�������c��O㾸����C�0��V:���8���,����6� �&#ҾO��6���2Q��(����p��K׽�Xɽ�Ž"�ɽ/4׽�	��	�u�#���G��8y�М���ľ� ����0(�pw8��K?�;���,��,�ؓ��Z۾%7���4��#⾾�پ; �C�ˡ,��<�\�A��^<��'-�&x�C���P�Ͼ<|��#Ն�1�[�/�7���.����mf�����
G ����Z��i�*�PH��mp��H�����!{�z��4 �d�4�z�B��E�G>���-�;�������߾Q_ʾ�ƾ3eվ�r��mX��)&�|�9��UF�/1H��?��+-���c����vξ0@��󉾩!f���D�y�-����*��W����"�*���*�/A���`�p���ģ�nɾ�f������E*�x�<��.G���F��Z;�I8(�8���a��&ؾR�Ǿ��ɾq-޾,� ����$-���>���G�}F���9�Ŀ%�����뾴���������~>[���=�Ž)�}j�Z������������#��5�?N���q�g���l��hMپR�����f2�˫B��xI�&3E��6�  "��j�����eӾ�ɾ�Ѿ�N��3	����<5���D��  �  &'��]"�A���Ӛپ���������_�՘2�����3�BPͽ������_���-���>���}�ս����R=���m�������΁�jT��q�o)%���'�e� �k������=�Ծ�����)���w���r��ž���ʰ	�H��8&���'� ��f�j�����;|p��Oτ���S�'y*����&�%̽�oЭ�j'���뵽W�Ƚ��D�:�%�֓M�ှ������ȾL��!��F$�X'��l&�[t��|�W��Ⱦ�髾=��������Ӿ�=��]��:"�yc*�G)�ׄ�i"�X��%�ƾ4-���끾X�R�X�-����Ѐ����Y^׽��ҽ�I׽R�彂������|�)�\IK���w�+����໾��例����^V)��E/���+�,��%����#;�Ѵ��߫�����.<˾y������C�,�O�1�-����>���a�-�ƾkآ��܅��^��v=��_%�����	����G�B4�����m�1��pM�w|r�|���	t����վ]���F��N#'� �2���5�� /�|d ������Ҿ�t���(���uɾ^很�����+�8�6�(C8��X0�� ��~��Y�ƾ ���P퉾�Uj�]vK�u5��m%��K�/�T���:���#�]o2���G��ce�ٴ��=栾��� �辏�	����i.�zR7���6�;�,�Q��՘����i�˾gC���.��?hѾ��@K��+ ���/�F8�r6�ү+��-��R���ྶ�<���Xꂾk`���D�gB1���#�f��UZ�.�� ��U+�>]<�1hT�Xju��^=��gfо������OW%���3��u9��5�!�(��|�8�r��-�Ǿ����4Lƾ�zݾ�B ������'�>5��  �  #����ی�羜�že��8�����a�{�;�R���S�e>��6н����[Ž�
�Ľ�ֽ\��c*��#%��E��`m�g����U���}ξ���6�,`��M��d������Qݾc������{���錾�ؗ������ξCY���r��A��4x�	[���޾�ڼ��k���a��
vX� 5��\����Xl罎|ѽƽCXŽJϽ��㽈K���+�0�yS��(~�J|��>j����پ�)����	�M���
�E���E��Ѿ:��c������%������3����ܾ�������!���$��
�l�����پ���������N��N�Y�ش9�b� �����l �D^������%h��r���
��6���T�$�z�֔��#���xѾ�C�	�d5�.���s�������վ<E��?ꣾ�t���$��K����Ծ����mc�����A����d������^۾�񺾕n���ӆ���g��[J���3�P�"����O�K<����+�\�+� �?��Y��&z��t��I����_Ⱦ�����/��m/��J����#j������@ھ�`���6��񄬾�ɷ��EϾ���Fq���?@ �	�!�����u���\:ݾ����톢�lC����t��	Y��^C� 3��(��O"���!���&��21�L�@�^�U�1�p�v�����u���إؾ�F���L��'��!��V ����I�	��8�=Ҿ��%����;�������پ���E��g��ky!��z �e�0M
����cҾ�R��"���p���Yl���R�m?��-1�!(�e$�g&�"�,�L79��J���a�e�C2�����a�ž}�循��F�xp�1�"���7���m���˾@��*M��ꩵ��'ɾ�~�&����\3��  �  ���t쾎8޾��ɾ�沾F���2j����m�0�O��@5�9���
� l�����Ὄ꽓;��Ͷ��6$��G<�b�W�@w�(͍���w��-Lоӳ㾰��4B��<��hӾ/ع�0���a����y���t�!������*Q����Ⱦ9�߾���:�����xھx�ľ٬��A◾�����g�0�J�9^1��V��C	��d���K�wi�M����3����R.�>�F��cc�-��)픾�c��~`��H[׾y���U����U�˾m谾����Q���Fw���z��'������d��վ1�꾼���;����T�q�پ�þoƬ�����o���E�k���P�7�8�U�$��A��M5�U
����p�"�u�6��jN�bi������|��󏩾�񿾂 ׾k 쾇���3 ��L���龝�Ѿ�U��d�������4 ��̌���a���趾��Ѿ뾒z�����Z� �q�󾙦߾��Ⱦ�c���S������{���a��wK���8���*���"��!�{#&���1��B���W�=�p��]���W���������ܒԾ�뾧�����)����:P��P׾�Ž�ҭ������왾���˥���ξ5a��F �����	�k�����u>律ξ0$��U���zoR���	q�<�Z�N�H�P�;�ej4���3��(:���F�X�וm�UN��������7	��|�ʾ������t���������� ���?.Ѿ���nФ����QQ�������y���o׾�n��)�� ��+M����Bnݾ��ƾj���1E��{i��Ę��Sk��\V���E��;�eR6��S8��@��@O�ugb�Wy��ԉ��ܘ�0��`&��>zԾ��뾜Q �����k
�nP�`������	˾�k��g���뜾e ��7x���ȾB4�}�����  �  )�¾f�¾��x���s��Yԛ�����Lo��Ԣs�x$[�GB�	#+�a�tt�	��������0���H� b�7�z��򈾬8��w����}��, ��|g���Jž�þY������j#���m���:f�v?R�Z�N���[�V�w�с��Ȫ��,�������n#ƾsľMx�������󥾂g���1��^܃��o�-�V� A>��(��2�����5���u�%�";���S�"bl�����^���z���棾1���3����¾edž�%��Y���0V���}��Ѕ{�*_��Q�GT���g�-Q��H���#��p����Ⱦ
�˾�Ⱦnn���O��宨��f��z]������mv���]�0�F�ڿ2��%�~��"��,/�kB��NZ�_$t��׆��Bw��3�Զ��ԁ����˾��ҾMӾ�̾���s�����it��[�v��<n���v�
w��KU��_խ��G��+оuؾ �ؾ�Ҿ3�Ⱦ[Q��H�������hr�������샾\�o��X���F�A�;��.9���?��qN�H�c��[|�&������������D���ˑƾ%1Ҿ�۾���t߾��־-vǾF��*X��Q����������1���"֛��Ȯ�oþ� վ��ᾠ�����ݾ/,ҾQƾ����T��u⣾����.R��l�}���g���V�|M�sL���T� �d��z�Ȃ������\���|\��#����ľX�ϾN�ھ�
��徱�ᾤ־~�ľ٥��	����-���������>��mء��s���Fɾ��پR�㾏w�DX�qپ�.ξIv¾���j���̇��'x�������w�.uc��U���N�3OQ��\��o�������[	���ާ��5��V���Hʾ־�l������ᾜLӾj���쨬��ݚ�*����܉�:����v��R�����'Ҿ����  �  �t��1ӣ��V��L2���@���z������	���u���ˈ�L�s��U���<�h,�\�'�5o/��^B�:F]��{���������.���楾������L���/���4���_��������χ��~q�iT�C
<�ve-�c�*��o4���H���d�⦁�� ��7~��y<��|���D��F�������dA��nۤ��1��G�������m���P���9���,�%#,�e�7�_qM���i�B�����;���ֺ��'[�����c���t���+󦾢��ћ��ڐ�������g�e&L�C�7��z-���/���>�`IW�>�u��ϊ�����У��ê�.f��⯾"I��[ﯾ9��� ��9K���薾�̈�$�s��6Y�3F�@>���B�p�R�`l�9���	��S����v��t�����������𶾿[���B��y��)���#��"�����{��+b���P�׭J��,Q��9c���}�:t��>�����l ������9)����A%���b��5���������&�������恾\Gk�:�[���W��3`���s�7ׇ�������]���ԧ��/���g�¾m�þ��þ�¾�M��$���<�����7���R҇�v�x��k�#4i��s�i��3���%��N������þ{Ⱦ�ɾ�4ʾ��ɾ�Ⱦt�ľ6��7����奾����
��[&y��(l��^k�9�v��\��&����գ��ı�������þ�nǾ\�Ⱦ�>ɾ��Ⱦ[Ǿ�~þ�;���3���)��'퓾	؅��`v�c�k�o�l��z�*���'���~ݦ�nr�����0Ež��Ⱦ)�ɾiʾ-�ɾ��Ǿc�þ���������C�������&v��Mm�.�p�b7������{�������·�Hs���dǾ=Lʾ{Z˾s�˾��ʾ��Ⱦ��þy��W��<���Q����z����v��p�P�u�����u������G����.���  �  ����ِ��>��	������#���tþ��¾����9��u ��25���<h���Q�<XK�2�U��o����)��߶��NA��`�ľ�þv�������7����a���/������7sr���Y���@�Z*�T��i�������$"�S'7��O��h��q���M-������xv��ﺹ���¾�]ƾ�Yþ3⸾�C��%f��6�F�b��FQ�0AP���_�l�}��ꑾZ٥��궾1¾��ž��¾�+����*�������r�����`j���Q��9��$��������$�=�.��]F�{`���z�����ރ��P������x︾��þ�Q˾27;��Ǿg������֕������<m���a���g��T}�JǏ����>�����Ǿ�Ѿ�Ҿ��;�oľ|	���`��������]���U���f��O���<�R0�,3,��-1�+�>���R�.+k������/���&��
��������W�ɾӎӾ�hپ��ؾ,$Ѿ��¾��������R��.z���&{�
9���x��;��������ʾ#mؾ�%߾>x޾��׾�;�¾���Ǵ��FȠ��l������H{�.�e���T��HK�BJ�z!R���a��iw����vʔ�2 ��X�����;,þ��ξھ�⾀|澎[�F�ؾ�Ⱦ�%�� �������B��`�������rr��o�����ž�־��^��I���Rھ"AϾ�zþ���pӬ��p���s��g���ȍy�N3d�r�T��L�P�M�%�W�� i��p��)��&�������`����@��Y�ƾٸҾZuݾ������9�ˈԾ-�¾�s����c����������������9���%����;�0ݾ��}��<���پ+�;����ڮ��\������i����j���:w�ˏc�$\V��zQ��U��Pb�2�u�磆��;��?����  �  ��n�%�����1���)˾�l߾s��Kc�B�l�վ�輾����mۋ��z�z}q��S���������YþPe۾���{��U����ܾf�Ǿ����p����jk���M�J�3�=z���
�����'��A�>���s�5O�td*���B���^��)��)���\��Y����ԾZ;�K��0�LH�6о;���@��Q����:x���v�ׅ�Jy��|Ѳ�:;@��p��
��-=�x־�2�����?���/р�)a��E�ێ,�^����3���+���j��F����τ#�<;�d�U��$t��[��o(��[��ٯ̾qf���������������ϾpX���0��񰋾7��g����ҕ�TV��Ǿ������ʥ������`��ݾ2[ƾM���d;���h��t�bsY�<TB�S�.�� ��������#c"�Pv2��G��G_��z�����g枾wd��fʾ�ᾖ]���v�7�o��X6쾈�Ӿdh��[��ڋ��Ȑ���՗��.������ܾH��l������:��m��%�⾠�˾-����?��N}�����m!m���W�m�E�x&9�e.2�g�1���7�TD�0mU���j�b聾^���$������i�Ǿ��޾m)������ӗ�5��y��k�վ�𻾽\��6���.���s�����x{Ҿ����\�_����\#������i�bɾ
���%���ݐ�\����l��EW�qF�:��74��5�X<�C�I�(S\���r��-��	۔����t@��z<Ͼ�k����1�Ф	�*��p����e辺�;u������'���$ޞ������¾�6ݾ.���]�H�	�(��!������ھ1Zľ9ϯ�7띾Pq������ Ij�SJV�?�F�K�<��69�aY<�p�E�f4U�i�I�������  �  cc�V���5����]ǾR 龌c����O���/�� ����	��A�����]#���Г��;��+�ǾA���lO��H�to�v���8p��=y��ǭ����]���8���h�����/jҽ��ŽX]ý��˽�߽�����L�H,��rM� 8w��T��v���(&վ
�����?���A�H
��v���Fؾ���]���]���1��}2��3���DԾU������0�������	�����@5ؾ֚���Ɨ�\"{��P�e�.�ܢ�� �.�)�ѽ.8ʽg�ͽ��۽���(�A<#�#�@��ce������;��b(žZ羿n����V�c�8
�����v=վ�s���8��~u���ʚ�����v�Ⱦ�����V@�	������h����s�ھ�幾a����(��g	a�9-B�qQ*�JQ����29��2�����C��,��;/���G�^g��1��Mw������Qݾ_����]�H������F�l���3���־�e������ᢾ6⫾Х��B���f�h���B��d�\���a�X����{ܾ-����#��-����$q��,U���?���/��5%�������\�$�N�.��C>�L�R��m��6���%���ݵ�$6Ծ�����-�x���� �=@!�i�բ����5׾�-��S���9���Rκ���Ӿ+��g�
������ �)� ����r�2f����־���ڝ�P���uo��T�
@���0�>�&�8"�K�"�P�(��A4�)�D�>�Z�V�v��k��*磾MH���޾ib �76�#D���!����b��ʼ�ʼ��ξ�+�������p�þ��߾� ���������"��> ���^�j�ȅξ2�������鄾Țj��CR�ڬ?��M2��%*��Q'�)�)�:�1���>��Q�Di�����  �  ��a��i��w�����۾�2�2�s#��c'���!����� �8�پ�P����E����夾�c��.����� �2l$�J�'�Kk!���������Ծa������5Z�o
/�R�����(ν����i%���B���˲��$Ľ�(ཛX�Ԋ �T�F�"y�yX��Oy¾e��J �Kb�y�&�M�'�q<�6'�c��X%Ͼ�&���͞��՝��b��7˾b��@��E��3'��'�U��e��F��[Qƾ�����5~�Z�J�:�#���^��hɽ{ظ��p������F�½��ٽ!������>6�;a��W�������־�� �d���H$�q�+�Z�)�ik�g��w$�H9̾B�������x��N��1�ᾑ9����w�'�Ƃ.�Ss+��q��/��E���ƾ���������X��5��/��B
�����o��Pr����d4��=�!��+;��s^������D��E�Ⱦ��5.�j	!��.��k2��-��G�M�l��oξix���I���Ἶ�־����K�&�$�jP1���4��.�J5 �O����ƾ����Ո�o3g�y�G��e1�"�!��)�l�Dd�����_!�)�/���D�g@a��ك�����ݼ���⾗���G��{,���6���7��-/�������~�Ͼ�j��	p����̾���j�����Iw-�d�6��7���-�G��r����ݿ�H[��ύ��H�c��F���1��S#��B�c$������8�&�{6�V1M���l��L������+�Ⱦ���/��}�!�D�0�'j8��66�7�*���H���k�b�ɾ����_¾v!׾����k]���#�_�2�=9���5�j�)�����w�op۾-���)}��߀�'^�8D�H�1�(%���4K�C��w�$���0�L�B�vN\����  �  ��c��M���i���o������#��k2�|k7��T1���!��9�US�E�ľ�-��E���Nk���̾d���s���/&��
4���7�s0�<���c	�9�&]���	���-[��e+�c���A�����.���e��B���-���a]��#ѽ�������jE���}�C����ξ�3������*�;r6���7��.���R���P߾ü�t�� a������B�ھ���}�LF,�F�6�B�6��,��dz�p�Ҿ펦�7ʁ���I�5���< ��Fֽqú��ꪽx	���>������]˽�j����G2���a����xĶ��b侃�
�A�!��&3�L�;�uk9���,���?.�۾>l���[���뵾�X;
��D'��=&��7�%�>���:��)-��F�q< ��1ѾX|���y����V��'0���п��A����޽���\����v��H`5�۬[�H����+��~[ҾU� �&��R�.�]j=��sB��m<�g�,������ܾs�þ����XȾ|徔�n�L�2���@�A�D�]�=��-����[4��^�Ͼv���M����c��A���)��`�8��x�J��������.h(�y�=�/\�(���K���Bþ���M�*'���:�p|F���G��>���+�$v������fܾ�ɾ�ǾaLپ(Z��k���V)��&<���F���F�	<��)��������ƾ��K%���_�g�?��Q*�����/�lS�q��Q����)/�L�F� h��x��()����о�&���f�xH.���?��^H�$�E�+%9�u%��b�A�oZվȾ�M;�h侄���P�]51�v�A�U"I��mE� �7�Ǣ"�P�
�v���������d���X�A�<�;*�]�����z�����P��I)�'�;�3zV�>8|��  �  �9e�wK���#���4�Q���p(�d8��==���6�P�&�@�j����ɾ���'����~��P�Ѿ,��j���A+���9�ԕ=�/�5�M�$�
���羞�������\���*�����۽Kc������4 ���M���:��@���v̽����/��lE����<G���}ҾX�}&�`�/�p+<��=��{3��� ��Q	�s�<��\6��������%T�����R�1�߷<� �<�DY1��i����86׾�G������/J���������ѽc��|w�������X��'`ƽ���f��_U1�;@b��`���๾�t�55�--&�T�8�ޓA��?�N�1�0!�l��]ྱ���T���ƹ��Ҿ���H�+�(�<�@TD���@�[,2��X��=�$վd����C��;DV�;�.�����f ����qݽ�ڽ
h�HQ�g�����3�o)[��U���(��\־}���� l3��C�\EH���A���1�Q���;���ྩvǾVA���g̾�'꾦]
��="���7���F��J�rC�o�1�5���?���ҾL�� �����b�Ǹ?�6�'�������q?
�bO
������&��;�1�Z��'��pX����ž���֊��L+���?�Q5L��}M�flC��0�g/�a����/�̾r�˾�ݾ����Sd�t�-�xtA�ߠL�A�L��WA��s-����#m���ɾ�7��?��#�]�_�=���'����3���%����q�������,�7�D�g�g��ǋ�ܨ��p�Ӿ���� �C�2�;E��+N�̢K��K>��p)����h���e�پD�˾ *Ѿx����z=��6��IG�3�N�BK��<���&�>�����!?���ǚ��
��W���:���'��l�����T��b�����&�Y~9���T�,�{��  �  ��c��M���i���o������#��k2�|k7��T1���!��9�US�E�ľ�-��E���Nk���̾d���s���/&��
4���7�s0�<���c	�9�&]���	���-[��e+�c���A�����.���e��B���-���a]��#ѽ��������jE���}�C����ξ�3������*�;r6���7��.���S���P߾ü�t��"a������F�ھ���}�QF,�L�6�L�6�
,��sz���Ҿ���Gʁ���I� ���< ��Eֽº��誽����:��ޓ��e˽lc�A|��B2��a��܏������^侕�
�S�!��$3���;��i9�^�,����h-��۾�k���[��O쵾�Y;v��=(�:?&�S7�Ӆ>���:�o+-��H�`> ��5Ѿ����|���V�D,0������wE��#�޽V�����������[5���[�7���6(���WҾ\� �!��Q.�rh=��qB�[l<��,������ܾ��þ%����YȾ��k�����2�H�@��D�X�=��-����h8��6�Ͼ�y���P��E�c��A�/�)�nd���^z���-����� i(��=�y/\�+(���K���Bþ���	M�*'���:�p|F���G��>���+�$v������fܾ�ɾ�ǾaLپ(Z��k���V)��&<���F���F�	<��)��������ƾ��K%���_�g�?��Q*�����/�lS�q��Q����)/�L�F� h��x��()����о�&���f�xH.���?��^H�$�E�+%9�u%��b�A�oZվȾ�M;�h侄���P�]51�v�A�U"I��mE� �7�Ǣ"�P�
�v���������d���X�A�<�;*�]�����z�����P��I)�'�;�3zV�>8|��  �  ��a��i��w�����۾�2�2�s#��c'���!����� �8�پ�P����E����夾�c��.����� �2l$�J�'�Kk!���������Ծa������5Z�o
/�R�����(ν����i%���B���˲��$Ľ�(ཛX�Ԋ �T�F�"y�zX��Oy¾e��J �Kb�y�&�M�'�q<�7'�c��Z%Ͼ�&���͞��՝��b��?˾l��G��O��@'��'�l��������QƾҚ��+6~�n�J��#������fɽ�Ը�qk��c����½S�ٽ���U���46��/a��Q��>�����־�� �����D$��+�`�)��h�O��A!�7̾�������1�������m;�A��G�'���.��v+�pu��3�KM���ƾj!������%�X���5��6�-H
����'�｟r�ۗ�1��8�>!�c#;��i^��}�� >���Ⱦ���S*��!�.�9h2��-�oE�K�^��mξow���I���⼾C�־>����M���$��S1�k�4�ѡ.�=9 �K����w�ƾ����Xۈ��>g��G�$n1���!�P/��p��g�����a!���/���D�:Aa��ك�����ݼ��⾛���G��{,���6���7��-/��������Ͼ�j��	p����̾���j�����Iw-�d�6��7���-�G��r����ݿ�H[��ύ��H�c��F���1��S#��B�c$������8�&�{6�V1M���l��L������+�Ⱦ���/��}�!�D�0�'j8��66�7�*���H���k�b�ɾ����_¾v!׾����k]���#�_�2�=9���5�j�)�����w�op۾-���)}��߀�'^�8D�H�1�(%���4K�C��w�$���0�L�B�vN\����  �  cc�V���5����]ǾR 龌c����O���/�� ����	��A�����]#���Г��;��+�ǾA���lO��H�to�v���8p��=y��ǭ����]���8���h�����/jҽ��ŽX]ý��˽�߽�����L�H,��rM� 8w��T��v���(&վ
�����?���A�H
��v���Fؾ���`���b���7���2��>���DԾi������B�������	������5ؾ$���#Ǘ��"{�+�P�,�.�1��̟ �$*但�ѽn0ʽ#�ͽ{�۽������,0#�~@��Se����$2��3ž�羑i���^R��^��
�״�� 9վqp��7��!u���˚�霬�<ɾ��Y��@D��������m�K����ھ�ﹾ�����0��1a��9B�|[*��X�����;��2�z��?��%�2/�{�G��g��)���m��b{��hFݾ{���5X�*��?���B�����-����־�b������ᢾ�㫾Ϩ������i����F��i����Yg������ܾ����T-�����h4q��:U���?���/��=%������G�$�L�.��E>���R��m�;7���%���ݵ�86Ծ�����-�y���� �>@!�j�֢����5׾�-��T���:���Rκ���Ӿ+��g�
������ �)� ����r�2f����־���ڝ�P���uo��T�
@���0�>�&�8"�K�"�P�(��A4�)�D�>�Z�V�v��k��*磾MH���޾ib �76�#D���!����b��ʼ�ʼ��ξ�+�������p�þ��߾� ���������"��> ���^�j�ȅξ2�������鄾Țj��CR�ڬ?��M2��%*��Q'�)�)�:�1���>��Q�Di�����  �  ��n�%�����1���)˾�l߾s��Kc�B�l�վ�輾����mۋ��z�z}q��S���������YþPe۾���{��U����ܾf�Ǿ����p����jk���M�J�3�=z���
�����'��A�>���s�5O�td*���B���^��)��)���\��Y����Ծ[;�L��0�NH�8о=���@��U����:x���v�'ׅ�Wy���Ѳ�Q;`�⾛��C��v=��x־�2��7������iр�E)a�oE��,�ܪ�o�C������'^�>����Gx#�E�:���U�t��P������N��)�̾�Y��������%�������ϾS���,��⮋���������Օ��Z��PǾ� �m��������������$ݾ�gƾ�ʯ��F��	s��p,t�݂Y��`B���.�' �`������G]"�Um2��G�o8_�Բz���ڞ��W��U�ɾNᾝP���p�i1�	e���-��{ӾUc����>���㐐�kח�;2��o���5�ܾ������ �+A�M{��Ð��˾����K��O���l��n2m�2�W�yF�Q09�L62���1���7� D��oU���j�遾����$�������Ǿ��޾s)������ԗ�6��{��l�վ�𻾾\��6���.���s�����x{Ҿ����\�_����\#������i�bɾ
���%���ݐ�\����l��EW�qF�:��74��5�X<�C�I�(S\���r��-��	۔����t@��z<Ͼ�k����1�Ф	�*��p����e辺�;u������'���$ޞ������¾�6ݾ.���]�H�	�(��!������ھ1Zľ9ϯ�7띾Pq������ Ij�SJV�?�F�K�<��69�aY<�p�E�f4U�i�I�������  �  ����ِ��>��	������#���tþ��¾����9��u ��25���<h���Q�<XK�2�U��o����)��߶��NA��`�ľ�þv�������7����a���/������7sr���Y���@�Z*�T��i�������$"�S'7��O��h��q���M-������yv��𺹾��¾�]ƾ�Yþ5⸾�C��(f��:�O�b��FQ�AAP���_���}��ꑾt٥��궾a¾!�ž��¾�+��{��s*������s������_j���Q�ӹ9�a�$�������������.��OF�j`��z�~���{w�� ���ꬾdḾ%�þeD˾+;��Ǿ�]��z����Е�����08m���a�X�g��Z}�1̏�� �������Ǿ�Ѿ�Ҿ��;
~ľ����n���+���������f��f���O���<��U0�~3,�p*1���>�y�R�ik��}���%������������	⽾��ɾ��ӾT[پ��ؾOѾ�¾9�����5O��px���&{�;���|��������)�ʾoxؾ�2߾7�޾��׾ �;�$¾ ���e«��Ԡ��w��đ��Y{���e� �T��QK�
IJ��&R���a��lw����7˔�� ���������S,þ��ξھ�⾅|澒[�I�ؾ�Ⱦ�%��!�������B��`�������sr��o�����ž�־��_��I���Rھ"AϾ�zþ���pӬ��p���s��g���ȍy�N3d�r�T��L�P�M�%�W�� i��p��)��&�������`����@��Y�ƾٸҾZuݾ������9�ˈԾ-�¾�s����c����������������9���%����;�0ݾ��}��<���پ+�;����ڮ��\������i����j���:w�ˏc�$\V��zQ��U��Pb�2�u�磆��;��?����  �  �t��1ӣ��V��L2���@���z������	���u���ˈ�L�s��U���<�h,�\�'�5o/��^B�:F]��{���������.���楾������L���/���4���_��������χ��~q�iT�C
<�ve-�c�*��o4���H���d�⦁�� ��7~��z<��|���D��F�������eA��oۤ��1��I�������m���P���9���,�6#,�|�7�|qM��i�]��8���j������t[��^�������݋��������ћ��ڐ�����g��#L�5�7�:u-�t�/��>�1=W�J�u��Ɗ���ţ�����JX���ӯ��:��"᯾�+��t���>@��Mߖ�2ň�o�s��.Y��.F�M>�=�B���R� jl�������������������3���M϶�r���'j��hP��s���!%���,�������{�-3b���P�.�J�l)Q��2c��}��l�����Ψ����B}��������&��BT��p๾6�������J�����2ၾ@k���[��W��7`���s�݇�F����������Ӵ��r����þ�þ#�þ=þ�[��A����G��D�������ه�2�x�k�~;i���s�-k����@��������^�þ�Ⱦ.�ɾ�4ʾ��ɾ�Ⱦ{�ľ6��;����奾����
��]&y��(l��^k�:�v��\��&����գ��ı�������þ�nǾ\�Ⱦ�>ɾ��Ⱦ[Ǿ�~þ�;���3���)��'퓾	؅��`v�c�k�o�l��z�*���'���~ݦ�nr�����0Ež��Ⱦ)�ɾiʾ-�ɾ��Ǿc�þ���������C�������&v��Mm�.�p�b7������{�������·�Hs���dǾ=Lʾ{Z˾s�˾��ʾ��Ⱦ��þy��W��<���Q����z����v��p�P�u�����u������G����.���  �  )�¾f�¾��x���s��Yԛ�����Lo��Ԣs�x$[�GB�	#+�a�tt�	��������0���H� b�7�z��򈾬8��w����}��, ��|g���Jž�þY������j#���m���:f�v?R�Z�N���[�V�w�с��Ȫ��,�������n#ƾtľNx�������󥾂g���1��`܃��o�1�V�A>��(��2�����5�����%�E";�ʌS�ebl���6_��F{��E磾��������i�¾�dž�%��B����U��*}��'�{�&_�ZQ��T��g�/K��ꎘ�R��-��^�ȾO�˾Ⱦm`���A��=���Z���Q��f	��\v�X�]�!�F�2�2�P
%�:}��#��2/�`tB��[Z��4t��ᆾ?���ك�������ĵ�&�����˾K�ҾEYӾ¼̾&���¬�����6x��Q�v�E=n�?�v��s���O��%έ��>��� о5ؾ��ؾ��Ҿ��Ⱦ�B��=���dz���f��-䃾]so���X���F���;��.9�U�?�yN�P�c��j|�8/���×�R���w��α��ڠƾI@Ҿ��۾����߾T�־D�Ǿه��F_�����d��G���񣍾0؛�cʮ�{þ>!վ�����;��ݾ=,ҾQƾ����T��{⣾����1R��q�}���g� �V�~M�sL���T� �d��z�Ȃ������\���|\��$����ľX�ϾN�ھ�
��徱�ᾤ־~�ľ٥��	����-���������>��mء��s���Fɾ��پR�㾏w�DX�qپ�.ξIv¾���j���̇��'x�������w�.uc��U���N�3OQ��\��o�������[	���ާ��5��V���Hʾ־�l������ᾜLӾj���쨬��ݚ�*����܉�:����v��R�����'Ҿ����  �  ���t쾎8޾��ɾ�沾F���2j����m�0�O��@5�9���
� l�����Ὄ꽓;��Ͷ��6$��G<�b�W�@w�(͍���w��-Lоӳ㾰��4B��<��hӾ/ع�0���a����y���t�!������*Q����Ⱦ9�߾���:�����xھx�ľ٬��A◾ ���	�g�3�J�<^1��V��C	��d���K꽔i�s����3����.�z�F�dc�`��h픾d���`���[׾̞�V�����Uι˾�簾��������Aw�,�z�<#������^��վ̅�"w������GH���پt{þ;���>՗������k���P���8���$�;�S��4��
�!����"���6�ByN�Xsi����ć���������l-׾%-쾬���9 ��V��[��{�Ѿ�Z�����g���\ ��H���e^���㶾S�Ѿ�뾳p����:� ����g�߾��Ⱦ�V��H��jꌾ��{�[�a�nkK�c�8���*��"�	!��&&�{�1���B���W�N�p�1g���b��'�������c�Ծ�����Y����d���Y��X׾̽����5����~�������j�ξb�G �'���	�|������>徕ξ8$��\����tR���	q�A�Z�Q�H�R�;�fj4���3��(:���F�X�ؕm�UN��������7	��|�ʾ������t���������� ���?.Ѿ���nФ����QQ�������y���o׾�n��)�� ��+M����Bnݾ��ƾj���1E��{i��Ę��Sk��\V���E��;�eR6��S8��@��@O�ugb�Wy��ԉ��ܘ�0��`&��>zԾ��뾜Q �����k
�nP�`������	˾�k��g���뜾e ��7x���ȾB4�}�����  �  #����ی�羜�že��8�����a�{�;�R���S�e>��6н����[Ž�
�Ľ�ֽ\��c*��#%��E��`m�g����U���}ξ���6�,`��M��d������Qݾc������{���錾�ؗ������ξCY���r��A��4x�	[���޾�ڼ��k���a��vX� 5��\����bl罜|ѽ$ƽ[XŽ!JϽ��㽣K��[�0��S� )~�||��xj����پ�)����	�h���
�>��JE��ѾD���	�����#������.��;�ܾ������������
���V�پ����Y���F��y�Y�B�9�(� ����Kg �;X𽝞�s��p������x�6���T�M�z�(ߔ��-��%�Ѿ=N��	�n:�����w�������:־,H���룾u���#�������Ծ����_����=�����^����T۾~纾!e��Tˆ�.�g��OJ�Ō3��"�.���M�t<����$1�&,�`�?��Y��5z��}�����mjȾ��龧������4�uO�i��n�����0FھYe��b:�������˷�GϾ��q���f@ � �!�����u���e:ݾ����󆢾qC����t��	Y��^C�#3��(��O"���!���&��21�L�@�^�U�1�p�v�����u���إؾ�F���L��'��!��V ����I�	��8�=Ҿ��%����;�������پ���E��g��ky!��z �e�0M
����cҾ�R��"���p���Yl���R�m?��-1�!(�e$�g&�"�,�L79��J���a�e�C2�����a�ž}�循��F�xp�1�"���7���m���˾@��*M��ꩵ��'ɾ�~�&����\3��  �  &'��]"�A���Ӛپ���������_�՘2�����3�BPͽ������_���-���>���}�ս����R=���m�������΁�jT��q�o)%���'�e� �k������=�Ծ�����)���w���r��ž���ʰ	�H��8&���'� ��f�j�����;|p��Pτ���S�)y*����&�,̽﷽{Э�z'���뵽t�Ƚ��5D�\�%��M�,ှ����ڑȾy��9��]$�j'��l&�Vt��|�����Ⱦ�諾̕���񟾊�����Ҿ�9�����l�!�O`*��)�3�������ƾ�&��恾�R���-�̾��u��B�"Z׽��ҽmL׽)�����1����)�"SK���w������绾��T��{!��Y)��H/���+����6��
��%;�Ҵ��߫�����=:˾����?��M�,���1�r-����`���Y��xƾ�Ѣ��օ���^��m=��X%������	�;��G� 6����t����1�zM�F�r������z��]�վ=���K��H''���2��5��#/�Dg �o!�k����Ҿiw���*��wɾ_���R��D�+�T�6�9C8��X0�� ��~��Y�ƾ���T퉾�Uj�avK�x5��m%��K�/�T���:���#�]o2���G��ce�ٴ��=栾��� �辏�	����i.�zR7���6�;�,�Q��՘����i�˾gC���.��?hѾ��@K��+ ���/�F8�r6�ү+��-��R���ྶ�<���Xꂾk`���D�gB1���#�f��UZ�.�� ��U+�>]<�1hT�Xju��^=��gfо������OW%���3��u9��5�!�(��|�8�r��-�Ǿ����4Lƾ�zݾ�B ������'�>5��  �  #-7�o�1��Z"���t��5,��)�����a�e�/���
�����E������?��# ��dʝ��׬��ƽ
��Kf��5;��p�)!��hžu������K'��4���7�
0��q	���l�����^妾�V���'Ծ�9��J��&�)���5�-�7���.������^5۾93��D����S�#D&��>��Eܽr��i���� ��ƀ���˱��q ׽[��j-!��M������ᨾ�&վY���	�Y�,�z�6��D6��+�n��vV�fؾ1 ��� ������Hb��fM㾫�x����0�7U:�Ľ8��,����N� ��Ҿ�K��%����Q���(�R��Rk�H׽^VɽHŽf�ɽ.7׽_�S�	���#���G��>y�cӜ��ľ�$����2(�Ty8�IM?��;��,��-�����[۾�7���4���ι�پP: �7�|�,�!<���A��\<��%-�"v�S�����Ͼ�x��҆���[��7�<������d������G ����'��%�*��H�<sp�L��j��྆��6 �x 5�y�B���E��H>�1�-�w�������߾�`ʾ�ƾ�eվZs���X��)&���9��UF�71H��?��+-� �f����vξ3@��󉾬!f���D�z�-����*��W����"�*���*�0A���`�p���ģ�nɾ�f������E*�x�<��.G���F��Z;�I8(�8���a��&ؾR�Ǿ��ɾq-޾,� ����$-���>���G�}F���9�Ŀ%�����뾴���������~>[���=�Ž)�}j�Z������������#��5�?N���q�g���l��hMپR�����f2�˫B��xI�&3E��6�  "��j�����eӾ�ɾ�Ѿ�N��3	����<5���D��  �  5�꾦�ƣѾ��������5�u��D@��L�E�ȱ������Wk�>L�;<��	8���?��lT��x��3������M��>=��M�"}���蠾���Oؾ���X\�/ 㾱�ξ���|������~g�ZJb�a�t�����ԧ���þX�۾le꾙�쾒����˾���V鐾�g�0/5��b��jڽ�쬽���?o���T�N�G���F�i�Q��Vj��]������6Iӽ���8/��`�3񌾷���waȾ�߾]U�K��Aݾ�>ƾ����{u����x�^�d�~�h��4S���C���о0�L�����Uf�39ɾ�ƫ��v���?c�&@4�+'����ꩿ����Q��-i�������������`��a����(彿����-��EY����뤾��þv߾����� ���/徱/̾����헾2�e����^����i���2�˾9?����P����u��(�q�̾)[��ۊ��Pl��G@��s� �������ѽ0�ý���0����\½]ν������[��t�/�]�T�����|r������J!ھt�����$��Z��}�뾬SѾUf�����5���`������鄭�v�Ǿ�㾶����U��r�� ��8��Ͼ�����Г�t�t���K�L�,����������L轶��K�_��,󽓶�����(��G���n��$���쬾Җ˾����G��~���w�ڀ��#l���ʾMR�����|���(��<���_���\Ѿ+�쾐� �9j�M�-���~P�4�ž;B��MP��dg�x�A���%�g��+���n����� ��������  �Z���^�� 6�hW�JI��Q����^��k�׾�m�̔����Z(�=<��3ྗ:ľ%Z��������J���LG��ک��W�ݾt|������  �  ��شݾI�˾Ud��rG��)q��=���A彘$������q��R��(B� >�>F�Q�Z��m~�� ��;������^D���J�����D�����8uҾp⾇�従�ܾNɾ�J���Ĕ�t}���b�7z]��@o��_��Ǚ�����h�վ�㾱��;�۾éƾ�\��*��d�Q3��+�.�۽񒯽 ���u���Z���M���L��7X���p�΅���x��B�ԽF����-� ]�����w��!-þ��ؾ��f侉(׾����1n���	��Mss�@"`�:�c�h�}�躔�(�����ʾ��߾���Z�w۾�Dľ���芾�U`� 3�9U����a�½)F��߆��8��z�������������ý���zf��5-�<+W�����f������
|پ�v�f����ﾮQ߾5Ǿ%���񾔾(W��:�|��Ѓ�듾�ԫ�5&Ǿ�Ą�4��l󾔄��Ⱦ( ��_��׽i���?������ڤ��Խ�ƽ;��a���!fŽ��ѽ���*� ������/�`�S��L��� ��[R���Gվ�������� ������徻�̾������%���*(��|(��X�þ�޾����I�e!�����T�澴�˾e	��] ��`Ls�X�K��i-���U7������l���佝N佀��O��?J�v\�O�)���F��Nm��r������ǾkT�w)��~�}+��e��#ᾔwƾ�ᬾ%N���M���������p����̾��<�����E�����_Y޾+���ѱ���؉��?f��%B���&�n*��g�ܡ���G����뽆	������o�m����6��V�?�� ����#��ˇӾ���i ��Y����D`�$۾�5��$+�������5��Fe���,��Ӿ��v�ؾ@�񾵵��  �  �Ѿ̾�p��F㥾H7��j�e��t8�������o�����4����f�0U��P�?7Y�%�n�a����ࣽ�OȽ�5��qo�&8D�=Es�sn��HାX¾$о�3Ӿr˾/s��:���I���l�2VT���O���_��ꀾĶ������w�ľg�Ѿ.�Ӿ�jʾ6��m����	��1�Z�w�/��u���4���mU�����D�n���`�Q�_���k�Ě���Ȗ�伳��۽|A�Lk*��{T�ᖂ�{{��A鴾�ȾKmҾ��Ѿy"ƾ2��mK��Oc����c�ҀR��U��Zm�������,]����ξ��ؾ�D׾�˾���͝�b#��xY�-�0�H��RT��1̽񛲽婡�$���e���0������~̴���ͽ"���\�,��,R�A�@���W����8ʾ��ھ��ᾲ�ݾ��ξ�?���;��������y�	o�� y�9/���ؠ�{���#gоn��:���o�� ҾT�����������<d��>��9!���
�Ɯ��o߽��нҁɽ��Ƚ��νLz۽Y+�q��g�'k1��Q���y�ː��x��&	Ⱦ,�ݾo����a�?־�����!��c���|􈾺���q������*���lо���|��l��h��oIؾ '�����AW���so��L��o0����YQ�����;���1�����B ��j
�U����,�ӧG�3�i�9��&��������վ>J�������X�|SҾ�I��9.��
y��ok��ߠ��_唾�9����ٴ׾�H꾧��s��pl���о����i蝾+����c�	�C�8�*����W�
�Ia����zD�V��f���^���x�'�"�r 9�ifV���{�~/�� v���eǾ^�޾^Sﾺ5��D����.";�崾-��~��Sh��p��nf��]����˾>�ᾡ��  �  ��������������=����W��\3��g��T��Uν.i��-U��/Z��`�v���q�/Z{������ל���ٽx����U=��Ac��K����������n���򼸾��������f ���u���S�9#?�2G;��I���e�FH��К��d���V���c��fN��ڼ��/�����w���O��-�������4%˽�ѭ�ϗ��Ո�����x��EL���D���B���ƽ����C���(���J���q�񞍾���7X��/f���t��ֈ���������mJj�'�L�>�A�JU�,Qw�4z���!��w|���0��ݘ��t!��G���4w�];Q��0�q���^ ��Z߽�ƽ���0N���ॽ�穽-D����ǽw"�p� ��z���.�
�M�Ger�E����V��괾.¾�}ǾH�þ +���㤾������|�@�c�.�Z��uc��{|�d����������~�ƾb\̾�wȾ�N���q��,��}Ɂ�a-_��p@���'�X���y*�Ϛ⽉Dڽ>PٽJ�߽���#���.� ���6�}�Q���r�����|P���Ƶ��Ǿ�Ҿ�Ծ^�;�~��Ea�� ���4��ޑ|��y�b�.���p5���庾�̾>�׾��پ-�ҾH�þA����ߛ�������l���O�r�7���$�[�L�
��c�1���4I�����?�	�&��\"�G�4��K�.h��?��a☾�����<��φо��ؾ��׾��;ż�/q��y۔��υ�(6|�%I~������,���]��ea���Ѿ�Fپw:ؾjξ����G����Y���B���c�}H���2��!�F?�>�
�im�p�� ����F��2���+�]�?��X��Nw�Gɍ�����϶��[ɾ|�־z�۾Z�׾�A˾3ɸ��H���ܑ�L��T5��k:��f��̀��S��',ʾk�׾�  �  ������������4���j���M�J�3������t���ν�|��A �����Ot���N��z���ώ���b׽b��$��~�#�R�;���V��Ws����-v��[����C����Q߈��1r��Q��6�v�%�c�"���-�UE��%d� ����ʐ�J���Hr��� ��/L������be�ړI�l0�]F�3���I�JyͽE���h���֙��9��䞡��7����ɽ���/-�n;���,�:�E��a�]�}��P������ԯ�����M������u�g��H�'Y1�V�%�,K(���8�fkT��v�N����+���Ġ�2`���a���o���̂��,i�pN�7�6���!� ���������fн."ý-o���½@н�g�*z �����1#�7�7�k9O��xi���xu��A��+��R8��h��f/��^���g�z���]��I��uB�N�I���]�R�{�Fӎ�C�������7��*-���'�����֊��~y�	�_�e�H���4��#�[�������� `󽙳�y3��ܣ��[����
0��/C�3�X�q�V ��L���wߢ�B���_�����wD��Ō���E��܇��p�r�8c�=�`���l��3�������������4��$���yc��+����=���Œ�Ǆ�B5p��Y��;F�i�4���%�����������^����*�#��z2�)fC�F�V��ul�멂��z���랾}j���ɶ��ܻ��9��Rϱ�����Ǔ�v��~�o���c�|?e�/�t�3����ʗ��㧾�����Ȼ�v���V���q��補��N���Հ�)�i��T���A���1�R�#����KY�&4�	���r��3�|1,�0�;���M���a�j�x�/\��3�������������������Ū���J��hh������2����o��h�O�n�-��ȡ���0��l�������  �   M|�6Z}�~�v�'�j�S\��fM�d�>���/�� �����W��a�߽��ƽ������O����̽��罊������b%��5�1D�NLS��zb���p��|��ƀ�p�~���r���^��EF��.-�bR�8��)	�����#�L�;��7U�}�k���{��r������|-x�Vk��>\��<M�[V>��/��#�ws�����Ru޽�Ƚ|���Q�����Ž<۽����^����ا,���;�̕J��wY��Fh��u�W'�����.|�sm�ӱW���>���&�e��F���������0�BK���e���{�愾�O��Km���c���>s���d���U��QG�jK8���(��b�9 	�����{��߽$��M������+��)���:��dK�[�Zcj���y�+U���������PÎ�t�������l�:�S��=�0].�)���.� �>���U�#Dp�V����5��!���L?��Q��"��*����)y�=}j���[�yL��}<��l,�Χ�����
��Y	�����	��S&� $7�ջH��Y�bj��y��y��3���~��IO���D���1��������:��>\h�yT�\�H�$G� OP���b��7{�����|���)��񳡾�Š�|M������42������~�޵n��^���M�.=�~C.�z�"�����D���!�v,���:��0K�j�[�Ql�Q{��"��ͩ��G%���暾����� ���2��<Ė��ċ�h!~���e�W\S���I��)K�?W��ok�j>��jَ��F��l֟�Zա�����8[��^m�����������<z���j�f�Z�UJ�N):�b�,�v#������ ��9(��{4���C���T��ie�Q^u�Q���ۉ�Xw���ޘ�H.��#���'��Ở�o����:��h{��Kd�^T���N�_�S���b�7%y�fi��=���ڞ��  �  =O�^�V�o�Z�h)\��F\� �Z��>W���O���C���2�����0�M����W�
Bܽ~}�:H��o=�F3%�r8��mH���S�S�Z�a^�m8_�9_��w]�9-Y�r�P���C�ٮ2����������R���⽊��������:�*��=���L���W��]��r`��Sa�b�`��^�E�Y���P���B�L�0�N��5
�9�������,������l[.�z|@�Y�N��BX��]��_�n6`��v_�.�\��^W�ŏM��$?��-�I����H5��Ӷ�ݚ�{B �ë��$�;:��M�Ϸ[���e�Pk���m��sn�U�m�Vk��re�s([��KL�:���&�]��T�	�����������#���7��|L��i^�\�k��t��By�`<{� �{��z���w���p�"�e�M0V�_�C��p0�$��(���-����}�!��p3�h�G��4\��um��"z�������K惾� �� d�������{���o�f�_���L�M�9��=*��L �G��:�#��1�wnC��$X�l�P�|��L���Hǉ����O����������4���&|��k�FY��F�::8�Z�/�*�.���5���C��V���j�z�}�7��������
��m���ΐ�J����f��Sӌ��*��%��P<p��<\��<I��B:�S�1�s@1���8���F�9�Y�=nm�A��U��kߋ�w���{Ə�����ŏ������ċ��Ԇ���K�l��X���F��8�Þ1��2��;���J���]���q�ځ�����L:���������>���˘��!3��P"��ֆ��l~�ݳk���W��4F�mc9�i�3��6��<@�^cP���c�O�w�ԁ��f ���%���U���<��me���⑾�E������0���s~��`k�y�W���F���:�l�6��S:���E���V��Yj���}��L���  �  ]|/�ѯ>���M�<]�e�k�v�w�iE~��}���r�]�_���G�cr.�Ξ�0L
��&����S����4�ڔN�_*f�~w�������w�-^k���\���M��?�( 0�C ����+����w���Ƚ�ݺ��a��������ս���M7	����_*���9�s�H�{�W�sg�~�t�f[�
����#�n�q�N�\��XC�߇*����Q��
�g���'��"@��pY��o�Me}��S��A��Iu�W�g���X���I�|�:��l+����(�ΰ���z۽"Ƚ�k��^�½ 0ҽ����	��x)��u:��J��3Z���i�y�9<��˶��]�������sz�/d�<*K�C4��#����{� ���.�o&E�HZ_�<�x�������:��5���<	���~�@7o�P`���Q���B�)�2��"�/a����t���s���  �ZM	�����w'��9�)7J�Z� 	j�6\y�K[��X�������K��]��������X����t��2\���F�QP9���5��n=���N�)�f�����Ȍ�=ĕ�Y���_����������i��K����u�Zog�OfX���H�K9�x+�47 ���@��32���)��d8�II��4Z�K�j�3Jz������)��4����������ڞ��Y�������獾z;����i���U��8J���I�d�S��f����?�����Y�����o����������sG���ʄ���z�Hhk�3T[�ϦJ��h:�T>,�Y�!����s��$���/�<�>�2O���_��	p�t[��3���Ɏ�:B��"Ӝ��0��"���qR���;��iՊ�1|���d�R|S��K�4�N�ˈ\���q������ �����Wۡ����*R��밚�|����*�������z��6k���Z�OYJ���:�Ʃ-���$���!���$�
-���9���I�ۗZ�D:k��  �  p���d4���N�шk��	���P��*T��j2�����>Ӊ���t��(T�˾7��%���� {(�9�=�,\��T}�p���Q����c���-��>+���d��T5h��)L�R�2���I�G���YϽ�2��Ė������#���M�����c�Ľ�a��U�j8�r�)�qB��Y]��8z��芾����@	��*���-��1'��en�p�M��4��L%��s$���1�>ZJ�S�i��<��;���C���y�y��Bԋ��d|�L|_��D�ie+���N��T�\gɽ�a��9����|������C᭽3P½�~ݽ�����i�5	&��;=��KW�b�s�䈈��ו�ˠ��6ѣ��3������y߉�_ms��pU�Ý?�*6���:��SM���i�ƅ�%ꕾD��6���/ħ�����-����	����q�KW�	�?��+�s��6R
�l����1�W4۽y�׽��ݽ͂�=a�j���3 �b�2�kH� �_�$�z�쥋����A��1Q��DD��xR��P3������f���S�3O���X���n�񆾂㗾=��͝����������Ω�m4�����%@��#fi�?mS��V@��/�eh!�F���e����q��F������!��r0��hA�1�T�Bj��=��1َ�r:�����鵾j廾Q���ܳ�~Ħ������q����r�2d��Sc���p�n���~z��T¤�E��V]��A���aC��4��� ��R��� ���`k�f�U�J�B���1�ؓ#����Y�����F��������5'�Z6���G��{[���q����C����2���_���
��A��@U���찾Ø��o/���邾Ieo�^Ke��li�a{�-s���⛾����%�������ǳ���p�����#����i��,����h��5T��B��%2��$�z<�+���'�JV����d;$�"�1�T�A�$�S��  �  ����4���Y�\S���镾�ʧ��س�������)D��+��$wy��V���>��8���B�V�]������C��.���v쑸��������D咾7�|��bT�*�0���������ͽ�o���}��ќ�������|�Y���}��k���u��_��p��$��E�Fl��̊��ƞ������p���	���v���q��a\��s�p�|P��:>��0=��M�,Sl�3䉾A ��໮�4��t���� ��	[��̝����o�#�H�7�&���
�����UŽ�b��s���;݊�h4���$������>P��A��86޽9����p:�1^^�(g���c��Z���Q����������C~��p���1�����u�U�Z���N�jYT���j�/ �������믾�𾾨�ž�þ9��������H��W�}��tX�j�8�����:
��i��nBܽ�i˽�����~��,�Ľ�"ѽX�佼-������%��@�_`�P����:���ث�������ɾ��;�?Ⱦ����m§�a����"��o�m��yg�Ls��8��Q\���]��R¾1�ξF�Ҿ�Q;���˦��M0��	T���kg�7�I��I2�r��aX����g���Ț�����, �ij���7 �22�ȫH��ld��/7���窾@ξ���ξJؾe�ؾ�$о���M髾ԗ�ȵ��}}�J|��5��ڜ��7^�����qLξ*�׾jIؾ��Ͼ�2������-ȗ�0K����f��J���3���!������	� ���8��� �K�?�BV�nP&�
p9�-qQ�^
o��0��f/��� ��Rž}nӾ"ھZ�׾`̾����(+������*����}��m���Y�����/$��
�ž�lԾ�۾4�ؾ�t;�8����t��pĀ���a�YrG���2��"��a�O�(��~�����0���!���1�n�F��  �  ���:��h�1���8V��S���"�̾�	ҾX�˾@�� 夾e���q�o�	nT�nvL��DY���x�p��+Ѫ������ξ��Ҿ�˾j���B3���[��ǩ`��4������g���c���ʆ����m��3^��[�9f�R~�&H����WHԽ�����$�A�M�7�}��Θ�gѱ�13ƾ�?ҾxuӾ3�ɾ񔶾_՞�*1��L�h�LS���Q��e������⳾��ǾݒҾs�Ҿ��Ǿ��8��o?����Q�=(�J���1ٽ���c-��q���G�s�D�k��q��L��+��⪽�̽)K��� �w�=�*�i�4���+���@��5hҾ�6۾%�ؾt�˾����= ��Ȉ��?q��c�Ԟi�(������c8��/�ƾFeؾYX�K�ܾ4Ͼdu����x���5�^�w�7��#����&��ɽ�L���ְ����ݳ�&;���ѽG��H������>���e��ቾ����1H��ԷӾ� �_�m����Ѿc{��뒣�y���E����{�C���0��������þm�پ��Q��'��'վ�轾�B���p���0k��SG�>h+�	��$��Rp�����罊 轥���5���L����*�@�C�fe�����
��績o�Ѿ�!��h6��-��/־�a��O���U���x����`������+��	l���dӾ^羍0�FD��Z�u�Ӿ����-���눾&h��@F��,�p�6/
�uK �k>�������c������G��z�ND2�aBN��r��Ў�޷�������پ�뾼`��U��a���Ͼ�d����󀐾�����P阾�K��isž��ܾ���������l�㾣1ξFǴ��0��)����`�	�A���)�La����9�A���T<��Mi����~����5>)���@��  �  Ƿ�"�?���s��ؖ�o��]q;�޾���ژݾQ�˾Ig��/���6�����b��Z�4h��j��>䝾t鸾@ѾR�xa�@�ܾ�ɾ%���ב��k��*9��^�������!ۑ�Uyv��Y�%IK�YI���R�=�i�/�������-,ͽ��rR'�[wU��܅�%9������U�־�k�v���ھ�žYt��zF��ߴx�
a���_�Y�t��~��G��J�¾ݭؾ{��h��=]ؾ¾������=NZ�GU+������ҽ>y������=u�u�`���Y��_��Jq�����5ܠ��<ý�����E�A�cs�W���³��Ͼݤ㾆���A�ܾ'bž,Ī��"���;���p�&�w�f��`H��'f��Vy־��j����޾0�ƾɿ���ό�Je��9��P����K\׽޽��I��O���Υ��e��M���[ǽ��x��`��`�?��mk�aď��Ŭ���ɾ�i�n�������.����ᾒ�Ⱦkt��E����Ȉ�������樝�:y���ѾV����U���1���^�ɾ��������7�o���G���(�,�Ep���i��1޽��޽� 彏��g����l�&�ªB��g�抾���Pþ�߾���� ��������wi���ʾ2ư�?ћ�{����I���晾��`�Ǿ�W�;���I�E��������ž���'���#k�oiE�6�(���Q�xe��g��EE��潑!����n��H���[/�u)N�&v����;ү�N;�s������f�^�#P��o�ݾ�"þ)D������!9��`�� 鷾�ҾC`쾫���-���[��?۾�k��Jm���1���b�W�?�>&�*y�E��.d��������;��+���U�����+%��u>��  �  ur��BB��Dx�hH��Q���&Ӿ)/�9�- ��<Ѿ�7��Z���8�����g���^��wm�b���|����O�־<�羅
��D�G"Ͼ���������n�q%;�����[� ��Ǝ��p��S��7E�C���L�}^c�H̄������?˽�e��(�ЂX�~�������ľ2�ܾ����)��>˾v�2ڔ��k~���e�5�d�;�z��������,Ⱦ��޾r��7w��q޾
4Ǿ��+_���]��,������н���>���9�n��iZ���S��+Y��"k��~���ɝ�����~(�>�[sC�^#w��!��e���pԾ���'T����2�⾰�ʾ��rr��cꂾ�~u���|� b���
������ܾ�f�W}���L�����JG˾�R��f/���g��{:�3��+v���lԽ����d���B���Ӣ�]���%���(Ľ
߽���2H�;�@�O�m�#���4��Ğξk龀0��� ��4��g����;KQ������R���
��ᣎ��ݠ�n���k�־8𾶙 ����|��C�龵4ξ㯾���q��H�+(������ ���콭m཯۽&�۽���ͷ�9��i�x�%���B���h�#k��Q����'Ǿ9��:����h��$�^^ ����}Ͼ�Y��o���>j�����������l��+"̾���`��������/����b�ɾ I��(����l�BnE���'��`�9w�6/��g�bB�q�����������X��.�UrN���w�n����ٲ���Ѿ���e��F��(L��L���㾞OǾ���Oʚ��Y��һ��$^��쭻��^׾����8a�S*�������t���	̣��~��icc���?�/�$�4������4����ａ����������w��$��>��  �  Ƿ�"�?���s��ؖ�o��]q;�޾���ژݾQ�˾Ig��/���6�����b��Z�4h��j��>䝾t鸾@ѾR�xa�@�ܾ�ɾ%���ב��k��*9��^�������!ۑ�Uyv��Y�%IK�YI���R�=�i�/�������-,ͽ��rR'�[wU��܅�%9������U�־�k�v���ھ�žZt��{F���x�a���_�^�t��~��G��Q�¾�ؾ���y��S]ؾ-¾���8���kNZ�fU+������ҽ�x������:u�a~`�Y�t_��Aq�줈�+ՠ�[4ýE�����.�A��\s����1���
Ͼw��\��4�ܾ͂"`ž�ª��!�� ;����p���w��f���I���g���{־��y�����޾ʃƾXé�Vӌ�uPe���9��U�����-c׽þ��L���P��%ϥ�]d���I���Vǽ�I��a����?��gk�����I¬� �ɾf�����V���Q��S�ᾚ�Ⱦ�r��J���Ȉ�
���v��󩝾�z���Ѿ�X����\X���5����,�ɾw���E�����o���G��(��0�Ot�q���㽶޽��޽�#彼��8�H��ك&��B��g�$抾���	Pþ�߾���� �������xi���ʾ3ư�?ћ�{����I���晾��`�Ǿ�W�;���I�E��������ž���'���#k�oiE�6�(���Q�xe��g��EE��潑!����n��H���[/�u)N�&v����;ү�N;�s������f�^�#P��o�ݾ�"þ)D������!9��`�� 鷾�ҾC`쾫���-���[��?۾�k��Jm���1���b�W�?�>&�*y�E��.d��������;��+���U�����+%��u>��  �  ���:��h�1���8V��S���"�̾�	ҾX�˾@�� 夾e���q�o�	nT�nvL��DY���x�p��+Ѫ������ξ��Ҿ�˾j���B3���[��ǩ`��4������g���c���ʆ����m��3^��[�9f�R~�&H����WHԽ�����$�A�M�8�}��Θ�gѱ�23ƾ�?ҾxuӾ4�ɾ򔶾a՞�,1��Q�h�RS���Q��e������⳾��Ǿ��Ҿ��ҾșǾ+ﳾ�8���?��3�Q�W=(�]���1ٽ,����+������c�s��k��q��C��춒�>ժ���˽\8������u=�t�i���@$���9���aҾ�0۾��ؾ��˾���@���kƈ��=q�}c�.�i����������;����ƾnjؾ6^ྵ�ܾ�ϾQ|���#�������^��8�|-�-��:4�ɽ�S��Dڰ�f���ڳ��4��F�ѽO��)��e����>�'�e��ډ��{��A��ѰӾ7��3����2�Ѿ�w�������[���5�{�L���3������u�þJ�پͯ辴����`վE�J���w���=k��_G��r+�3�����{}��٧��罇'���:��/N����*���C��e�����
��績r�Ѿ�!��j6��-� 0־�a��O���V���y����`������+��	l���dӾ^美0�FD��Z�u�Ӿ����-���눾&h��@F��,�p�6/
�uK �k>�������c������G��z�ND2�aBN��r��Ў�޷�������پ�뾼`��U��a���Ͼ�d����󀐾�����P阾�K��isž��ܾ���������l�㾣1ξFǴ��0��)����`�	�A���)�La����9�A���T<��Mi����~����5>)���@��  �  ����4���Y�\S���镾�ʧ��س�������)D��+��$wy��V���>��8���B�V�]������C��.���v쑸��������D咾7�|��bT�*�0���������ͽ�o���}��ќ�������|�Y���}��k���u��_��p��$��E�Gl��̊��ƞ������p���	���v���q��c\��x�p�|P��:>��0=�(�M�@Sl�A䉾S ������54������� ��M[�����4�o���H���&��
�"��kTŽ/`���򖽣׊��,�����؍��5@�����!޽�+����_:�2L^��]��BZ��֚��.��A��������w��	������u��Z��N�L[T��j��#������������ž�þ����u���QR����}�`�X�>�8�z��zF
�}���Pܽhs˽�������Ľ�ѽ���:�������%��@���_�ݡ���0���Ϋ�Ƶ��{�ɾZ�;8Ⱦ����*���m���\ ���m�!zg�-s��;��{`��Jc��!¾#�ξ3�Ҿ�[;�����y:���]��0~g��
J��X2�����c�'��ߝ��L�������/ �cm�N��9 �;32���H�md��C7���窾Eξ���ξJؾh�ؾ�$о���O髾ԗ�ȵ��~}�K|��5��ڜ��7^�����qLξ*�׾jIؾ��Ͼ�2������-ȗ�0K����f��J���3���!������	� ���8��� �K�?�BV�nP&�
p9�-qQ�^
o��0��f/��� ��Rž}nӾ"ھZ�׾`̾����(+������*����}��m���Y�����/$��
�ž�lԾ�۾4�ؾ�t;�8����t��pĀ���a�YrG���2��"��a�O�(��~�����0���!���1�n�F��  �  p���d4���N�шk��	���P��*T��j2�����>Ӊ���t��(T�˾7��%���� {(�9�=�,\��T}�p���Q����c���-��>+���d��T5h��)L�R�2���I�G���YϽ�2��Ė������#���M�����c�Ľ�a��U�j8�r�)�rB��Y]��8z��芾����@	��+���-��3'��in�v�M��4��L%��s$���1�VZJ�s�i��<��X���j�����y���ԋ�De|� }_�)D��e+�5����R�Xdɽ0]��T���Xs�����Tѭ�\<½�fݽ�����X���%�5'=��5W�O�s�-}���˕������ƣ�c*�����؉�[cs��iU�ޙ?�.)6��:�/YM�\�i��˅�o��L�����ϧ�&����������q��`W��@�Q�+���^
�c���>署:۽�׽f�ݽ�w콲X����% �O�2���G�`�_��jz�ݙ���百�5���E���9��?I��y+��a���ꀾ�f�}�S�G3O�
�X�{�n���� ꗾg��`���m�������Tک��@��1"��&L���|i��S�wi@�3�/�Dv!�����o��������J����>�!��t0�&jA��T��j��=��Iَ�~:�����鵾o廾Q���ܳ��Ħ������q����r�2d��Sc���p�o���~z��T¤�E��V]��A���aC��4��� ��R��� ���`k�f�U�J�B���1�ؓ#����Y�����F��������5'�Z6���G��{[���q����C����2���_���
��A��@U���찾Ø��o/���邾Ieo�^Ke��li�a{�-s���⛾����%�������ǳ���p�����#����i��,����h��5T��B��%2��$�z<�+���'�JV����d;$�"�1�T�A�$�S��  �  ]|/�ѯ>���M�<]�e�k�v�w�iE~��}���r�]�_���G�cr.�Ξ�0L
��&����S����4�ڔN�_*f�~w�������w�-^k���\���M��?�( 0�C ����+����w���Ƚ�ݺ��a��������ս���M7	����_*���9�s�H�|�W�tg��t�g[�����#�q�q�R�\��XC��*����	R��
�{��3�'� #@��pY� o��e}��S���A�|Ju��g�{�X�f�I� �:��l+�����'�u����u۽EȽ�`��S�½ҽ�i�j����be)��`:��uJ�Z��i�u�x�m/������������fbz��d�KK�r;4���#����� ���.��/E��f_�-�x�>����͌�F��󟋾b��G&~��Po�p�`���Q���B���2���"�`k������� �� �G	�����j'�M�8��#J�iZ���i�ABy��M��դ��Ǯ�����񇔾�{��/P����t��(\���F�M9��5�rr=��N��f�F����ь��Ε��d���l������횐�gw���,��`�u���g�<{X�J�H� .9��+�
B �W%�.���7��)��g8�wI�w6Z�I�j��Jz�ک���)��C��� �����������Y�������獾};����i���U��8J���I�e�S��f����?�����Y�����o����������sG���ʄ���z�Hhk�3T[�ϦJ��h:�T>,�Y�!����s��$���/�<�>�2O���_��	p�t[��3���Ɏ�:B��"Ӝ��0��"���qR���;��iՊ�1|���d�R|S��K�4�N�ˈ\���q������ �����Wۡ����*R��밚�|����*�������z��6k���Z�OYJ���:�Ʃ-���$���!���$�
-���9���I�ۗZ�D:k��  �  =O�^�V�o�Z�h)\��F\� �Z��>W���O���C���2�����0�M����W�
Bܽ~}�:H��o=�F3%�r8��mH���S�S�Z�a^�m8_�9_��w]�9-Y�r�P���C�ٮ2����������R���⽊��������:�*��=���L���W� �]��r`��Sa�c�`��^�G�Y���P���B�P�0�S��5
�K������&��V��)�����[.��|@���N�^CX���]�Ƽ_�-7`��w_���\��_W��M�I$?��-����V��8-�����*��9 ������$�A:���L���[��oe���j�	�m��Xn� �m�=k��[e��[�V:L���9���&�����	����w������#��8�)�L�4}^��l��t��\y��W{�h�{���z�٪w��q���e��AV���C��{0�o�����.�W��̼!�ff3���G��#\��am��z����t��]؃���uV��E���\�{��o��_���L���9��6*�HI ����	�#�71��yC�T3X�,(l���|��X�����IՉ�o����������L��7A���<|�p�k��$Y���F��E8���/�j�.�j�5���C�-�V��j���}����������
��6m���ΐ�V����f��[ӌ��*��"%��W<p��<\��<I��B:�U�1�u@1���8���F�9�Y�=nm�A��U��kߋ�w���{Ə�����ŏ������ċ��Ԇ���K�l��X���F��8�Þ1��2��;���J���]���q�ځ�����L:���������>���˘��!3��P"��ֆ��l~�ݳk���W��4F�mc9�i�3��6��<@�^cP���c�O�w�ԁ��f ���%���U���<��me���⑾�E������0���s~��`k�y�W���F���:�l�6��S:���E���V��Yj���}��L���  �   M|�6Z}�~�v�'�j�S\��fM�d�>���/�� �����W��a�߽��ƽ������O����̽��罊������b%��5�1D�NLS��zb���p��|��ƀ�p�~���r���^��EF��.-�bR�8��)	�����#�L�;��7U�~�k���{��r������}-x�Wk��>\��<M�]V>��/��#�{s�����`u޽�Ƚ����p�����Žq۽����� ��*�,��;�P�J��xY�\Gh�Ǩu�(�D���E.|��rm� �W��>�D�&�|���A��~�[x�E�0��3K���e�w�{�4ۄ��C���`���V���$s�\{d���U��;G��78��x(�1U�������s�4�߽��位���h��R�]�)�# ;��yK�z"[�||j���y�ab����������Ύ�+~��2遾�l�ڷS�;�=��`.�^)���.���>���U��6p�㒄��+���}���2��,�������񃾤y��dj���[��eL�>m<�C_,�������
��Y	�4����e^&��17� �H�b�Y�gj�M�y�N���A�������\���Q���=��𨕾F$��>B���ih�L�T�Y�H�8G�sTP��b��:{�����1��*��9����Š��M��Ю��A2������~��n��^���M�3=��C.�}�"� ���D���!�v,���:��0K�j�[�Rl�Q{��"��ͩ��G%���暾����� ���2��<Ė��ċ�h!~���e�W\S���I��)K�?W��ok�j>��jَ��F��l֟�Zա�����8[��^m�����������<z���j�f�Z�UJ�N):�b�,�v#������ ��9(��{4���C���T��ie�Q^u�Q���ۉ�Xw���ޘ�H.��#���'��Ở�o����:��h{��Kd�^T���N�_�S���b�7%y�fi��=���ڞ��  �  ������������4���j���M�J�3������t���ν�|��A �����Ot���N��z���ώ���b׽b��$��~�#�R�;���V��Ws����-v��[����C����Q߈��1r��Q��6�v�%�c�"���-�UE��%d� ����ʐ�J���Hr��� ��/L������be�ۓI�l0�_F�6���I�SyͽQ���h���֙��9������7��Źɽ+��f-��;�0�,���E�ua���}��P������������7���2���g���H��U1�s�%��D(�o�8��`T�)v�����#������xU��XV��%d��E����i��ZN���6���!�a��������
Zн�ý�m��B�½�Iн�w�� �O���A#���7�;NO��i����]����L��@6���B��@q��D7��ņ��#�z�L�]�d�I�vB�p�I���]��{�͎����������!������显�ʊ�Lgy�Z�_���H���4�|�#��}�4�r����Z�����9����e���0��AC���X��$q�],��ʶ��좾�̮�,���"��[N��w���6M�������r�d"c���`���l��5��Y�����������?5��c����c��D����=���Œ�Ǆ�S5p��Y�<F�p�4���%�����������_����+�#��z2�*fC�F�V��ul�멂��z���랾}j���ɶ��ܻ��9��Sϱ�����Ǔ�w��~�o���c�|?e�/�t�3����ʗ��㧾�����Ȼ�v���V���q��補��N���Հ�)�i��T���A���1�R�#����KY�&4�	���r��3�|1,�0�;���M���a�j�x�/\��3�������������������Ū���J��hh������2����o��h�O�n�-��ȡ���0��l�������  �  ��������������=����W��\3��g��T��Uν.i��-U��/Z��`�v���q�/Z{������ל���ٽx����U=��Ac��K����������n���򼸾��������f ���u���S�9#?�2G;��I���e�FH��К��d���V���c��fN��ڼ��/�����w���O��-�������9%˽�ѭ�ϗ��Ո�.����x��bL���D��C��)�ƽ���(D�D�(���J�O�q�.������tX��`f���t��Ĉ��s�������|Hj�G�L�>��A�CU�vHw��t�����1u���(��������裾|���!w�*Q�C~0�{���R �UG߽��Ž:��fH��uߥ�멽+L��)�ǽ�3�^� �ׇ��.���M��wr�ܖ���`����G7¾�Ǿ�þ�1��餾����T�|�!�c�n�Z�1sc��v|�����ҧ������ƾ�S̾dnȾE���g��P���	����_��`@��t'�����u�j򽉑�@ڽ�Pٽh�߽����*���g� �9�6�R���r�q����Z��ѵ��ǾSҾ�Ծ��;���ug��菱�9����|��y�e��������6��q溾��̾��׾ëپN�Ҿ]�þP����ߛ�������l���O�z�7���$�`�O�
��c�4���6I�����@�	�&��\"�G�4��K�.h��?��a☾�����<��φо��ؾ��׾��;ż�/q��y۔��υ�(6|�%I~������,���]��ea���Ѿ�Fپw:ؾjξ����G����Y���B���c�}H���2��!�F?�>�
�im�p�� ����F��2���+�]�?��X��Nw�Gɍ�����϶��[ɾ|�־z�۾Z�׾�A˾3ɸ��H���ܑ�L��T5��k:��f��̀��S��',ʾk�׾�  �  �Ѿ̾�p��F㥾H7��j�e��t8�������o�����4����f�0U��P�?7Y�%�n�a����ࣽ�OȽ�5��qo�&8D�=Es�sn��HାX¾$о�3Ӿr˾/s��:���I���l�2VT���O���_��ꀾĶ������w�ľg�Ѿ.�Ӿ�jʾ6��n����	��2�Z�x�/��u���8���rU�����V�n���`�p�_���k�ߚ���Ȗ�����۽�A�k*�;|T�����{��m鴾ȾlmҾ�Ѿk"ƾ�1�� K���b����c��}R�C�U��Um�����'	���X����ξՌؾp>׾�˾E���HƝ����=�X��0�y���C�"$̽}�����������d��?3������Xմ���ͽw!�G���,��8R�	N���H���g?ʾ�ھ	��(�ݾ��ξpC��s>���Ë���y�7o�y�j-��0֠�Ȇ���bо����i���Ѿ<����f����0d�ׯ>�0!�_�
������߽'�н�~ɽ��Ƚ9�νD�۽�5�W���o�Ru1���Q���y���������Ⱦr�ݾh�뾕ﾺg�4D־���c%��i����������js������﬷��о�侷���󾀰�~Iؾ+'�����HW���so��L��o0����\Q�����;���1� ����B ��j
�U����,�ӧG�3�i�9��&��������վ>J�������X�|SҾ�I��9.��
y��ok��ߠ��_唾�9����ٴ׾�H꾧��s��pl���о����i蝾+����c�	�C�8�*����W�
�Ia����zD�V��f���^���x�'�"�r 9�ifV���{�~/�� v���eǾ^�޾^Sﾺ5��D����.";�崾-��~��Sh��p��nf��]����˾>�ᾡ��  �  ��شݾI�˾Ud��rG��)q��=���A彘$������q��R��(B� >�>F�Q�Z��m~�� ��;������^D���J�����D�����8uҾp⾇�従�ܾNɾ�J���Ĕ�t}���b�7z]��@o��_��Ǚ�����h�վ�㾱��;�۾éƾ�\��*��d�R3��+�0�۽󒯽 ���u���Z���M���L��7X���p������x��b�Խ[����-�& ]�����w��8-þ��ؾ(��n侂(׾�����m��R	��=rs�� `�=�c�Ԋ}�I���-���c�ʾ��߾��꾹V龠s۾PAľ�����劾eO`�X3�*P�*��\�½�@��$���$}��
���Ï�f�������&�ý��;k�j;-�c1W�'����V���پ+z�=i��[��T߾7Ǿ���������W��R�|��Ѓ�*꓾qӫ�G$Ǿ�|����j1������Ⱦ����
\��n�i���?���������Խ��ƽ���}����gŽ��ѽ�佷� �a����/�b�S��O��0�� V���KվW��Q���w� ��	������̾񪲾.��f��	����(��
)����þM�޾$���X�n!�����\�澺�˾i	��a ��fLs�]�K��i-���V7������l���佝N佀��O��?J�v\�O�)���F��Nm��r������ǾkT�w)��~�}+��e��#ᾔwƾ�ᬾ%N���M���������p����̾��<�����E�����_Y޾+���ѱ���؉��?f��%B���&�n*��g�ܡ���G����뽆	������o�m����6��V�?�� ����#��ˇӾ���i ��Y����D`�$۾�5��$+�������5��Fe���,��Ӿ��v�ؾ@�񾵵��  �  N���d�����}�Ht^��:�������	��GU��FI�)��8�����ͼ�4���8��J	���ټ�H�!:(� �[�y���ҁ���C��p ��/E�b7i�����|���Y������nH|���\��I<��� �������,�V�/���N�R�o��셾r���Fˏ�w��dxy���W�-�2�����d޽&y��vN��$UI�wj�;J�~���Ҽz�Ѽ�\༴# ����{B��G{��\���ֽV
�'�-���R��(u��臾B����������Gs���R�r�3���(�Ա�M#���>��`���������ޔ���������?{�EX���3��?��罝���*���w���U���@�q6��4�k:��>H��}_������f��澺�����:�o0��8U��Fz��{��L�����L9��[x��%肾�Oe��H���3��z,���3�.H�6
f������������΢��D���m���΄�Bje�ZA�= �)��6޽u@�����M������ጽS;��!�������`���˺�(�ս����Q?���2�B�U�{�����Pݞ�����l'��c$��&���逋��Vw���\�-�L�stJ��JV��=n��;���,����a������a��Ƞ�������;r��CN�f{.�^��# ��a�R5ͽ]���0��Yױ����]1���;����ʽ��޽�G��� �y*���I��"m��'���h��ȧ���������I٦�Q_��2���r��:Z�=�M�hhO�_��y�%��6&������^������<������ ��fg��kD�f�&����[��N߽��̽���$5�����������i��lȽt(ؽJ/ｙ��v1�	�8�y�Y�S-~������١��n���<���\��.x�������F��'�n��Z�c/R�N�X�Z�l�U'���/ä�Ty���  �  ����5���Tw��Y��6������Y��J��!cL��x�������ռ�R���C���0ƼY��cp��	,���^�����[������(���@�Ԁc��-���Q��}��H��ǭu��GW���7�X8������	� ���q+�$�I��i��c���������ۅ�y7s��R�2/�+���ZܽfE���X����L��y#�Ez��.�v�ڼC�ټ���S�]��F�>�}��T����Խ�G�LV*���M��
o��Y��N@���ꊾ%t���m���M�m�/�Ƌ�}����$����:�A=[��{{��k������=��~F���ju�(�S�9�0��{�h>�Jϸ�9p���e{�$�Y�#�D��!:��8�~>��WL���c����������!/�L��t�-��RQ���t��8��m������q�������e`�D��x0��k)�xh0�b<D�,Ea�j	�����ǚ�ɞ��S���!��q���fa�Dr>�	��m6���޽�ѿ��ꩽ�c��w���~䎽47��s�����`i�������K׽������=Q1���R�o�v��Ռ��o��eϤ��G���q���m��篈�p�r�H#Y���I�|WG���R��j�+\���|��4.��ِ��|ګ��ť�-���W3��S�n�L�v-��C�p� ��佪<Ͻ ��/?���۳�ه��;?��XS����̽�u�3l��g���)���G�ͺi�����X���7���"��4ɪ��E���:��ys��aVn���V�ܖJ�@L��i[�O4u��\��晾���q��;䪾����Q���*�����c�U�B���%�R���������l�νýU@������,���{���ʽ�%ڽr��������b7�zW��Lz�uꎾ����	����_������������:҃�(�j�
�V��O�.U�6�h�&�������\��\����  �  ��}��ew�Qe��8J��0+���(a߽�|���-���mW���+��}�`�lټw�Ӽl�߼,R�����{�8���h�!c��^����=e�5���S�,um���}����H�w��c��zG�\�*�c�������Y�
����).;��:X��p�H���7���w��b�y0E� �%���m�׽�5v����X���0����1����T�� %����e2,�KSR�91���{���$ѽ��R!�>�@�F<^���t�Ȕ���4����r�``[���>�<�#�>��-Z�X���{��
.���K��Ji��5���G���Hf}��he��G��e(�@����޺��a�����[Yg��*R���F�{_D���J��GY�q�򂉽㚠��ﾽ�����
��t'���F�Ȏf��>���.��#R��ی�P���o�8�R��8��'�� ��%'��F9���S�^�q������O�����t������su���V���7�]}�}����XŽ3z��"�� D�����XO���Ι��������½�Nܽ�O����P@-��J�C�j�= ��U���L��v��J��$�����@�e��N�}@��z>��I��8^�T.z��ǋ��<���ߟ����5ś��吾:q���0e�wF��6+���j��@꽹�ս}�ǽ�����k���ꪽ��ƽ�\ӽ,�潠h ����Ԧ'��TB�)�`��5���X��s�����*9��La���~�xCb�G�L���A��BC��Q�M�h�����������:T��TR����������DP{���[��;>�9�$�]������D� �ս��ɽ�½XϿ��D��qǽ�Fѽ���.���$�	����u4�B�P�S�o�v���룕�P���=������T���_��\�y�W�_�UFM��[F��.L��]�X�w�a��P̗��8���  �  "�^���Y��\K�O�5���������ٽ�.������ػn�?E���%�.�����6A���/�V;�e�/�AKR��D�f˛�Dj�����>��or%��5>�Y�R���_�Mb�ȴY���G�,00�������]콫��N���s�ǽ%�ת>���S�w�`���c��C[�m�I���2��c��� ��8ս*ܯ�.?���Dq��J���-�f�c��B���Eg*�K�E�:k��`�����Ͻ�����f8/�B�F���X�J|b�UXa��U��xA��5)�e������ct���j7�t�s75��N���b��lm�>(m��Hb�20O�W7��>����B�������K��⽐�*����tj��d]��Y�gr`�+�p�5����>��[��T�ǽ��������\A9���R�
Ci��#y��z���z��8l��dV���=�x(�p������B���(���?���Y�9Hq�����x���R��Dmv��$a�?bH��q/�����*�n�t�нaD��y���h��g��� ���ޤ�Vz������{Ͻ�D罱F����5)��dA��A[�}Ot������<���Ό�����/r��j��iR�w�>��2��)1�P:��L�<�d���}�����Y��«�������܄�\~r���X��@���)�����MU�����V1Խ�?ʽ��ĽɜĽ!ɽ�Xҽn8཮���}��y���&���<��'U��n�*1��\Q������}��Պ���a��,h��QP���=��r4���5�=�A��U�2kn�U���̌�c����(���d��@�����j���Q���9�c�$�:]�l6����e}⽟�ս_�ͽz�ʽ�I̽��ҽ�ݽ��p/��H��{�)2�"I�Tb�)�{�����������#���~��>e���N��?��39�7>��:M��mc�A�|�<ʉ�K푾�  �  �x;��>9�H�/�2� ����������ڽAD��^���勽�@o��lM���3�>$$��  �.�'�� ;�
�W��r|�����$$����ǽ|�jW��Z���'���5�Y$>���>�T27�Z(����� �cP�Q�˽��ǽ��ս��"���� ��s2��=�"�@��<�LU0��P ����*���ڽ�v���������#t��CT��!=��~0�C�/�(�:��P�#7o�B���Ù��&|����ս�����9����-��L:�"4@��>�S�3�Lp#����ό��(�ܽd�ν�ҽ�轇��L���/���@��5J�f~K�=�D�=�7��t'�/���;�YB�(�ѽ	;��`楽�甽�函�g��Fz�g���
���x����D����ٽK�����	������,�k�>��,N�L�X��u\���W�R~K���9�a�%��,�	�\��^�����!Z(�~�=��Q��]_�z�e�Ad�
�Z�e>L��;���)��D�t�
�����Z��<ҽ�z½����ǒ��%��m���������н1N�r���U
�����`(�@�9��L�s�]�h*l���t�7Av�2To��Ja��N�9�;���+�CK"��,!���(���7�ƁK��:`�=�q��g}��]���{�yp���_��N��<��M,�m��,����7���/p�F�۽ Yս��Խ�uڽ�e彠���D���ަ�h�)�d�9�)K��]�T�m���y����K�}�\^s�Y�b���N�g;��',��$���%�J:/� �?���S�ɘg�yTw��	��0G��2y���k��[�?I�P@8�[�(�#:�x!�{�:��������޽��ڽ��ܽ���8|�G�T���B��w$��U3���C�T�U�ϓg�fw�OԀ�݉��C��t�s��`a�7%M���:��+.�~h)���-�@�9��K��W`�=Bs��y���  �  ���x ��?��&��Q�$�����mսx���ޫ�!���͂���e��zQ� �K��V�XTn�����������1:ɽ��ݽ&�񽜞��=���c��h��:���b������ӽ�z��q������)o����ǽ/�?9�9y�E��C6 ��v��S��d��-	��=����뽝ؽ�%ý7w��[)���$���8m�#�\���[��Sj��킽i��ri��������Խ�������[k��������n�����
����kc�J��q\ν�X�� ��}���v½�;޽`  ����P	��U(���+��C*�(�$�rv��l�*.
�p� �N��ڽ��Ž����ߡ�L�������������+���}ɽz��v������P��h�8T%�;�.��|6��;��;�>�5�M+�����[�Y�����v��v���Ai��F!��&1�r=�<�D�&�E��}B���;���2��)��P ����}�������|޽�Ͻ�ǽ��Ž/U̽��ٽ��٩�YS�`��w�#���-���7�v�A��K��6R��U�.LT��nM�f�A��;3��e$�4����e�cw�XQ"�+�1��gB���P�N0[���_��=_�nZ��R��H�T?��95�	!+� ������
�(8����e��뽣9� �P	����{���K)�!V3�>=�m�F��P��UX��]��h_�e�[�$R�|jD���4��T%�ܲ�m����E&��(�,�8�>�H�g�U�^^�=�`��^�'eX���O���F�y=�c3�()����	>�H�	�,=�3��<��dS�>=�����+����Hy&���0��;���D�J�N�X�W�Kq_�a�c��c�~^�	+S���D���4�>Z&��B����c�%��3���C��+S���^��  �  �@���L�i��E�=e�Lq����.���S��{�ؽs���a��Г��h$���c������b㗽�t��}�ǽ���kP���4����^	�VT
�]E
�V	�D�� �pL�"Oڽdh����b2���.�����C���g�������0ѽ�=�����z���	�i���{�7/�`�
��8�[#�lI��iٽC������`K��F���-���C��;ؼ��ֽ�/�Ţ���$���	�l����/B�q	�_��aj�����-սü��w���%��=̎�fꑽ�E��gЎϽ�&뽀����������������AY������4�o�����ؽj)ý5;��	z����������׽9G�|��8�B�+I!���$�XQ&�X�&��&���#�ӕ��g����l��j��?ٽ��˽p�ǽ��ͽ��ݽd���*��z���P ���(��].�[l1���2�<3��:2���/���*��R#�a��E�}��bｩF��ཿ�轲`���5	�ͯ���#���.�Q�6���;�ݠ>�|�?��/@�}[?���<���7��0���%� E�=��d���� ��x �B��m�v����'��4��>�&1E��rI���K�!L�_�K��J�(vF�?:@��7���+������6	����BX���b.���ɰ)��Y5�B�>�#E���H�֬J�n-K�)�J��H�fE�6�>��&5�_w)���/��_����D���K
���xP ��-��8�szA�m�G��K�ҟL��
M��vL��xJ��NF��Y?�9�5���)�S!�.��R�	�p)����@����[%���1���<��qE��K��4N��O�	�O��"O�b�L��HH���@���6���*�/��B����3	�6���������X*���6�l�A��  �  �rԽ@h�*����F�������_��)��{����`!ӽ�Ƿ����۠������h��p�۽8;��Q�������f�� >���9��/����p�?�׽�Uý��J���W���Nl�0>Z��+W���c��}�c���#�����euѽ����o���h����Rm�l��:� ����I������qѽ�s���F���q������ͽ�콏$������AB �;������F����2���V�4�ӽ����	�������Є���q��[g�Ym��&��0>���ç��n���G׽� ���IA�#o�z$ �p(���-���.�"P*��� �����`�Xo�v,ֽ��ͽyuӽ��K���O"�<]/�+d7� �9��7���0�A(� �����/��A��<�۽jȽ�۸�r����P���������Vн�/�j��)
�	�6]�Ej)�sG3��z<�V�C�r�G���F���@��F5��&��P��8
����� �V��C�����0��@�v�K���Q�nR��`N��7G���>��z5�d,�2(#�
��?��r��=������_(��/�(�콊#���*���_b��I(�H�2�zp<��F���O�5�W���]�_`�7�\��9T�P�F�	7�8['�W�����=<����D�%���4�Y�D�ueR���[��8_�3�]���W�ɖO�uCF��<��3�)�ō���LI	�) ����C�1S��������3�G ��!�r�,�|�6�b@��J�isS�}t[�#�`�B>a�
x\��UR�!D��24��w%����������f� ��.�K">�=�M��*Z��a��c�1�`�^�Y��KQ�n�G�`q>���4���*�L+ �v��d�������������������>��z�Bv ��]+��  �  M���+۽%����_�4�!���0�_U:��h<�/*6�g(����h���߽��Ƚ½0ͽ��(���6��y-��:��>��;�fy0�9!�C������Wq۽Pp��ɺ����It���S��[;�R`-�N+�x�4�h�I���g�C���9o��S6���ѽr�e{	��p��L,�@�9�ڮ@�L�?���6�o�&���sZ��zI޽1
̽��ʽ9O۽�������"�$��5���>���@��(:��k-�k��@�
�ZC�m�ӽ')��Ο�"���Pq��fU�yC�x�;�^RA�"�R���n��牽֟����#(ԽH���8
��_�^�.���>�=�J���O��L�z�A��l0����e
�YB���ｐ���*������-���A� #Q��Y��X��{P���B�!�1�� �ބ�O� �<#置,н�J���֫�K���W ��)~��O����,���I��!bǽ]�ݽ�����E	����$�)�`<�ܵM��\��Tf�c�h�ћb��0U�O�B��/��=/�������@�$��F8��|M�Mj`���m�}�r���o�{e��qV��@E��4��S$��_�Z*
����P�콗.޽��ӽ�yν�ν�6ս"�����>���"�51(���7�X'I�G
[���k�^�x�0��x�~���u�P�e���Q���=�ȵ-�ً$�% $��),���;��#O�k1c���s���}��t�N6y���l��\�@J���8�:)�v<�������'���o��LL۽ )ֽ�׽j�ݽe�齭*��D	��}��h���-��@>���O�M�a��q�?o}�7��q�~�.s���a�a|M�v�:�8�,�Ћ&��()�c#4��vE���Y�1Im��|�����O���!z�l���Z��6I��y8��i)�l��9�����*����콵��S�ཇ��c�콵8�����|��u��  �  i��ݍڽ̷�#/�2S7�{�L�0/[���_���X���H�d�1�p���&�3��C���5�!�~�*8�;\N�� ]���a�3[��(K���4�&��W��zcؽ���M����ar�RJ�B},�����h��
�W���$�&�>�G�b�����Х�<uɽ����:�.�+�D��rW�!�b�o<c���X���E��y-�>�^�E����[���k�lw*�g�B���V��8b���b�)�X���E��.����xb��!vͽ{���U���X�k�<�H�0��5!� &�?=!�FS0���H���j�9��s@��&ǽk��K���'��A�0	Y��cj�H�r���o�7�b�W�M�s�5����:s��^��3�]�aP/�`�H��]a���s�.H|���y��m�2�X��L@�s.'�S��L���zֽ���>���ɗ��9��h���n��j��c/��Y��������gɽ��������A0���I�� c���x�B���!䅾���ZOu��^��lF��Y1�Գ#��2 �V�'��8�=pP�=j�V���@���Ê�qŇ�~���j�0GQ���8��"�����D���׽6sʽ ����ɽ�3|��"�ýY�ͽ�Nܽ�J����a�EW$���9���Q��ck������c��e吾�#�����G��*-l�Z�S���?���4���3��>���P�"i�Kʀ�͊������Ր��ԋ�f����Om���S��x;���%���i%����wc���ҽ�ʽ)�Žܟƽ<6̽�uֽL^� 0���.	����!�+��<B��3[���t�=텾Zw���k���5����_Yf��&O�\>�Uc6���9�G�HQ\��Fu�����U��8a��SOg��O��ݘi��SP���8���$�g��'�ڜ��R��Eڽ�ӽ��нD'ӽ�jڽ^M�s���LD�y���  �  iѯ�/��dE��,�gL���f�L�x���~��xw��Zd�q�I�8�,��i�H�����������D�3�AQ��j��{��T���x��d��0H�{�(�{�	�4�ܽV3��d��,qZ�t�0�mn�[m ���켪���������%�6�I�<|��F����ɽ<���4��8�<�0�Z���r�?����:��t�v�ie`�iD��'������������$��@�0-]�Xkt��������t�G/]��~?�������ν�ң�7o����R��o/�� ���
����I��%���}0�܇Q��~�'ל�x�½#�����Y4�mT��vq�]���<Ј�
�����Q[g��J��Y0����G��^��9)�s�B��h`�ӹ|��툾���Eڋ�����3	n�H�O��\0�g�� ����νH�����������K����x��gw���~�Hi��V���Oڥ�@���?�ݽP������8�8�X�I�w�]���p��x�������E���1�v��?Z���A���1�D-���5��I��	e��|������P����;��Z7���l��~d}�Ow^��@�m�$�H(�����޽��ʽ�ɽ�������{}��Ot�������_Ͻy�⽎x���#t$��}>�Dd\�|��	��l����.����֚�,���Eb���?f��:O��B�\TA�M�[c��)�x卾4���5��L'������-$��2�~�`_���@�M�&�������F���ӽ�ƽ\���*��������ʽ�ؽ@	�(d���=e-���H���g���������ɜ�C桾�l��!���<:����{�5�`��L�Q�C��HG���V�y�o�Wf���8��y��%��h砾$���XƋ�o�x���Y��<�
�#�=���y ����XWٽCIν��ǽ��Ž�
Ƚ-�ν��ٽ{�� �_���  �  ������}T�D�7�w
[�a;y�Wˆ��4���4��Yw�z�Y��:��P������g��m$���A���a�m~�*���j���9��6�u��[V�73� 2��⽳E������I�N��y#��� ����Ӽ�,Ѽ w޼���y��,9=�Ŏr�Oz��s�̽Cr�z %���H���j������h��-�����r�*cS��"4�e��6��6��ȟ���0���O��o��P���t���`������m�@^L���(�\���Xҽb���� |�r�F��/"���
�0���}���������M#�@gD��r�����jb½�������a>��3b��r�� �������c/���͉�Ңx�;JY�S<���&�HQ�{�!�0�3���O��Qp�`���K������>K��o���s}��[���7��f����i0̽�v������X���tu��l��+k�]r��瀽H���`������Ǧڽ���@�]�?���c�rp�����ZМ��O���n�����}����g��nL�ɵ:���5�v<?���T���r��剾6t��'��7����Y��D��������h�S2F���'��+�����8ؽĽ����d��gP���7������ۺ���Ƚ�Hܽߣ���)���%��C���d��9��T'��[����������f
��b���2
��ѿr�WwY��	K��4J�fW�2No����Җ�R���Dת�XЪ�a���mu���Å� �g���E�N(�{=��j��4���̽��8���Ӵ�u���#���Eý�ѽ<�dh�$N���/�x�N�-xq�h���?˚�٦�����A������ؔ���+l�BV��^L��kP���a�[�|��a��˔���ܨ�ϭ��\��S��#~��Y5��a��h@�x�$�Ә�j����h��ҽY�ǽ@���z��������ǽ��ҽ��X���oE��  �  �̱�B�꽩�r�;���`���z�������~��_���>�)"��N�%�	�#��Os(���F���g�����_������䉾	@|�5�[���6�O��)u�t���X܄�o�K��x�Ƽ��޼�˼ ɼ�Gּ�b���f���9���o�oF��;νL��L(��}M���p�����ۏ��9����x�U�X�ڍ8�t����v���(��5�u�T��_u��釾�K���4��������s�Q���+���Խ������y��KC�*�����������Ɲ����3�Dn@�H�o�y��F�½K����˼A��Ag�[����F��/r�����RS��d�~�6a^�A'@��*�he ��+%���7�QT���u����y���(`��9��Ł��G���AY_���:�-������Ե˽����-�� H��Sq�yh��/g��Vn���}�+6���p������ڽ���g� ��B���g�_/���镾�����,�� )��o���_���\l�0CP���=�Z9�p�B� �X���w��⌾�蛾4쥾�Ш�����z��7Z��`l�7�H��(��g�`3��Տֽ�½�ش�(M��7D���-��1쯽
����sƽjڽ1W������&�~�D���g�������N=�����^�������㛾 ����*w�*]�c.N��RM�"�Z�Ԟs�һ������A��㭮���������|���"���*k���G��&)��7��9��lH޽�ʽ/׽�I+��.в��o������-����Ͻ�f�'�� s�%�0�o�P�Bu�� ����py�����N䮾����痾�~��Ip�&�Y�CtO�5�S�*ke�"���p6���蠾����l������f��IP��X����c���A��6%��Y��E���|�3{нE�Ž����Ъ�������Ž��нl�὾��,���  �  ������}T�D�7�w
[�a;y�Wˆ��4���4��Yw�z�Y��:��P������g��m$���A���a�m~�*���j���9��6�u��[V�73� 2��⽳E������I�N��y#��� ����Ӽ�,Ѽ w޼���y��,9=�Ŏr�Pz��s�̽Cr�z %���H���j������i��-�����r�+cS��"4�g��9��:��͟���0�əO�o��P���t��
a�����F�m�u^L��(�����Xҽs���r |�~�F��-"���
�W���Ԫ���q������B#�ZD�v�r��UX½�������$>�J-b��o����������,���ˉ�0�x�kGY�\<���&�Q��!���3��O��Tp�g���hM��o���6N��� ��.z}�-[���7�ul������9̽�~����m]��E{u�l��+k�8Zr��䀽C���Z��	�����ڽ���;�"�?�
�c�&m��ې��B͜��L���k��}��@{���g��lL��:���5�p=?���T���r�_牾{v���)��,���]��wG���ą�d�h��8F�Ɉ'��1����JAؽ�ĽD���Vi���T��(;��X��)ݺ�H�Ƚ�Iܽ�����)���%��C���d��9��V'��]���	�������g
��c���3
��ҿr�WwY��	K��4J�fW�2No����Җ�R���Dת�XЪ�a���mu���Å� �g���E�N(�{=��j��4���̽��8���Ӵ�u���#���Eý�ѽ<�dh�$N���/�x�N�-xq�h���?˚�٦�����A������ؔ���+l�BV��^L��kP���a�[�|��a��˔���ܨ�ϭ��\��S��#~��Y5��a��h@�x�$�Ә�j����h��ҽY�ǽ@���z��������ǽ��ҽ��X���oE��  �  iѯ�/��dE��,�gL���f�L�x���~��xw��Zd�q�I�8�,��i�H�����������D�3�AQ��j��{��T���x��d��0H�{�(�{�	�5�ܽV3��d��,qZ�t�0�mn�[m ���켫���������%�7�I�<|��F����ɽ<���4��8�<�1�Z���r�?����:��v�v�ke`�kD��'����$�������ǒ$���@�G-]�wkt�1���6���;�t��/]�b?�g������ν�ң��n����R�Dl/������
�e��������_h0�FnQ��j~��Ŝ��½���=���M4��`T�jq������ʈ�*z��^��VTg���J�	V0����ԋ�����;)��B��n`���|�=�F����ߋ��ǃ��n���O��h0����E.����ν}���锚��!���Q��5�x�!hw��~�mc��g���TΥ�P���ݽ.��߸���8��|X���w��V���j���{�������d�v��:Z�R�A��1�6D-�x�5�ÙI�e����Ď�d���UA��=��%s���q}�D�^�S@�(�$�3�"���޽{�ʽ�ս�c��x���-����y�������bϽ���#z����|t$�&~>�`d\�|��	��o����0����֚�.���Fb���?f��:O��B�]TA�M�[c��)�x卾4���5��L'������-$��2�~�`_���@�M�&�������F���ӽ�ƽ\���*��������ʽ�ؽ@	�(d���=e-���H���g���������ɜ�C桾�l��!���<:����{�5�`��L�Q�C��HG���V�y�o�Wf���8��y��%��h砾$���XƋ�o�x���Y��<�
�#�=���y ����XWٽCIν��ǽ��Ž�
Ƚ-�ν��ٽ{�� �_���  �  i��ݍڽ̷�#/�2S7�{�L�0/[���_���X���H�d�1�p���&�3��C���5�!�~�*8�;\N�� ]���a�3[��(K���4�&��W��zcؽ���M����ar�RJ�B},�����h��
�W���$�'�>�G�b�����Х�<uɽ����:�/�+�D��rW�"�b�q<c���X���E��y-�C�^�$E����w���k��w*���B��V��8b���b���X�&�E�.�%��oc���vͽ����栌���k�s�H��0��*!�m� *!��:0�Q�H�*�j��#���'��I
ǽ�{:���'�ːA�'�X��Sj��r��o�a�b���M��5�|��Bp�/^��5�a��V/�I��ha���s��V|���y��(m���X�)^@�??'������s�ֽI	���P��'ח��B���l��3o��f��'���}��{u��MRɽ��彃�����00��I��c�&�x�瑃�m܅�2����Cu���^��eF��T1���#��2 ���'�/�8��wP��Fj�p���.G���ˊ�·����R(j�|YQ�O�8���"�:.���~7���׽݄ʽ�����ս�������ý�ͽ�Rܽ�M�)���b��W$�Ȭ9���Q��ck������c��i吾�#�����G��--l�]�S���?���4���3��>���P�"i�Kʀ�͊������Ր��ԋ�f����Om���S��x;���%���i%����wc���ҽ�ʽ)�Žܟƽ<6̽�uֽL^� 0���.	����!�+��<B��3[���t�=텾Zw���k���5����_Yf��&O�\>�Uc6���9�G�HQ\��Fu�����U��8a��SOg��O��ݘi��SP���8���$�g��'�ڜ��R��Eڽ�ӽ��нD'ӽ�jڽ^M�s���LD�y���  �  M���+۽%����_�4�!���0�_U:��h<�/*6�g(����h���߽��Ƚ½0ͽ��(���6��y-��:��>��;�fy0�9!�C������Wq۽Pp��ɺ����It���S��[;�R`-�N+�x�4�h�I���g�C���:o��S6���ѽ	r�f{	��p��L,�B�9�ܮ@�M�?���6�s�&���Z���I޽E
̽��ʽ[O۽)���ݐ�I�$��5��>���@�):�-l-�����
��D�G�ӽt)���͟�����:Jq�`]U�.C�V�;��:A��R�P�n� щ����������Խ҉��$
��J�P�.�$�>�c�J���O�y�L�)rA� a0�����_
�/;��Qｵ�����Ֆ�,�-���A��2Q��,Y�b�X�B�P��B�X�1�)/ �H��� ��B�~Gн�`���竽����>&���~��b�g"��&:���Lǽ�ݽs����3	�>��C�)���;��M���\��@f���h�9�b��"U���B�/�J�s,�݃����f�$��O8���M�y`�ˢm���r���o��e�M�V�$WE��04�1h$��r�];
��%��+��qD޽��ӽ��ν��ν�?ս2��(���?�h�� ��1(�K�7��'I�c
[���k�l�x�<����~���u�V�e��Q���=�ʵ-�ۋ$�& $��),���;��#O�l1c���s���}��t�N6y���l��\�@J���8�:)�v<�������'���o��LL۽ )ֽ�׽j�ݽe�齭*��D	��}��h���-��@>���O�M�a��q�?o}�7��q�~�.s���a�a|M�v�:�8�,�Ћ&��()�c#4��vE���Y�1Im��|�����O���!z�l���Z��6I��y8��i)�l��9�����*����콵��S�ཇ��c�콵8�����|��u��  �  �rԽ@h�*����F�������_��)��{����`!ӽ�Ƿ����۠������h��p�۽8;��Q�������f�� >���9��/����p�?�׽�Uý��J���W���Nl�0>Z��+W���c��}�c���#�����euѽ����o���h����Sm�n��<� ����I�
�����qѽ�s���F���q��!��7�ͽ"�콺$�Ө�i���B ����K���G����~���W罔�ӽ_�������d˄��|q�eGg���l����!)��8����P���%׽p�����*��W� �Y(���-�r�.��=*��~ ����V�Wa꽚$ֽ7�ͽzӽ�潗S����]"�sn/��w7���9�p7�%�0��0(������)$�;S�[1��۽�|Ƚ�踽#���iQ������V���Dн��RL��r
���GG��R)�S/3�Ub<���C��G��F�m�@�h75��&�lG�F2
�x��' ���JJ�|����0�� @�j�K�?�Q�@�R�AyN��PG���>�+�5�{,�v=#�;��-�������n��9�==彂��p+���-����c��J(���2��p<��F���O�M�W�
�]�n`�C�\��9T�W�F�	7�;['�Z�����?<����E�%���4�Y�D�veR��[��8_�3�]���W�ɖO�uCF��<��3�)�ō���LI	�) ����C�1S��������3�G ��!�r�,�|�6�b@��J�isS�}t[�#�`�B>a�
x\��UR�!D��24��w%����������f� ��.�K">�=�M��*Z��a��c�1�`�^�Y��KQ�n�G�`q>���4���*�L+ �v��d�������������������>��z�Bv ��]+��  �  �@���L�i��E�=e�Lq����.���S��{�ؽs���a��Г��h$���c������b㗽�t��}�ǽ���kP���4����^	�VT
�]E
�V	�D�� �pL�"Oڽdh����c2���.�����C���g�������0ѽ�=�����z���	�i���{�8/�b�
��8�]#�rI��iٽM������vK��c���B-���C��~ؼ�ֽ_0�`���2%�/�	��l�Y���B��q	����j��
��N+ս����|r��$������cܑ��3��Rش�,tϽn뽃��������������\���A���<����a���h�lؽ*ý83��Wx��#!�������׽�^�̊�pJ�V�>_!��$��i&���&��7&�p$�����z����i��8��Lٽ��˽�ǽ�ͽA�ݽ����������^> ��(�G.�T1�߱2�:�2��"2�߯/���*�@#��	�9�qs�/V�u@㽂����dn���?	�4��0�#�ݭ.�#�6�a�;��>�]@�{I@��t?���<��7��/0�Y�%�{T�6�#��?� �� �fG��q�{����'�_4��>��1E�SsI�ށK�A!L�{�K��J�:vF�M:@��7���+������9	����DX���c.���ʰ)��Y5�C�>�#E���H�֬J�n-K�)�J��H�fE�6�>��&5�_w)���/��_����D���K
���xP ��-��8�szA�m�G��K�ҟL��
M��vL��xJ��NF��Y?�9�5���)�S!�.��R�	�p)����@����[%���1���<��qE��K��4N��O�	�O��"O�b�L��HH���@���6���*�/��B����3	�6���������X*���6�l�A��  �  ���x ��?��&��Q�$�����mսx���ޫ�!���͂���e��zQ� �K��V�XTn�����������1:ɽ��ݽ&�񽜞��=���c��h��:���b������ӽ�z��q������)o����ǽ/�?9�9y�F��C6 ��v��S��d��-	��=����뽡ؽ�%ý>w��e)���$���8m�N�\�%�[��Sj��킽Ti���i��1����ԽA�������k�X��g��lo�6���
�����b���KWνcQ������eo��ce½�%޽����������2B(�o�+�N-*��s$�_�V��
��� ��*�l�ٽ�nŽn	��Iҡ�� ����L������N�ɽ�������&��De�C��k%���.��6�4;�c0;�u�5��+�]���e�Xf������潰��� `�5:!��1�`=��qD���E�hfB���;���2���)��: �������z��K �Uj޽��Ͻ�ǽ#�Ž�[̽�ڽ8"���c����R�#���-�8�tB��,K�lOR�z�U��aT�Y�M���A��J3��r$��>���l��|�LU"��1��iB�%�P�51[�&�_��=_��Z�&R�0�H�l?��95�!+�̈ ������
�-8����j��
뽥9� �P	����{���K)�!V3�>=�m�F��P��UX��]��h_�e�[�$R�|jD���4��T%�ܲ�m����E&��(�,�8�>�H�g�U�^^�=�`��^�'eX���O���F�y=�c3�()����	>�H�	�,=�3��<��dS�>=�����+����Hy&���0��;���D�J�N�X�W�Kq_�a�c��c�~^�	+S���D���4�>Z&��B����c�%��3���C��+S���^��  �  �x;��>9�H�/�2� ����������ڽAD��^���勽�@o��lM���3�>$$��  �.�'�� ;�
�W��r|�����$$����ǽ|�jW��Z���'���5�Y$>���>�T27�Z(����� �cP�Q�˽��ǽ��ս��#���� ��s2��=�#�@��<�MU0��P ����*�� ڽ�v���������#t��CT�"=��~0�u�/�i�:�9�P��7o�����&����|��(�ս���i���1�-�XM:��4@�,>�"�3��o#�9��0���_�ܽ�ν��ҽ轶��r���/�s@�$J�kK�ձD�D�7��_'����h(��콛ѽ���%Х�}֔��ه�tZ�!Dz�K������������(���ǧٽT����	������,���>��AN�P�X�:�\�s�W���K�(�9�B�%��2�>����������Q(�9=��
Q�'M_���e�d�ŹZ��(L� �:��~)�]1���
�a����i彑&ҽ�j½�ﶽ����~��U��������н�d�;;���e
�;��8u(���9�A1L��]��@l�
u��Tv� fo��Za���N�и;�v�+� S"�3!�|�(�K�7�]�K��<`�z�q��h}��]��m�{��p���_��N��<��M,�{��6����A���7p�L�۽Yս��Խ�uڽ�e彡���D���ަ�i�)�d�9�)K��]�T�m���y����K�}�\^s�Y�b���N�g;��',��$���%�J:/� �?���S�ɘg�yTw��	��0G��2y���k��[�?I�P@8�[�(�#:�x!�{�:��������޽��ڽ��ܽ���8|�G�T���B��w$��U3���C�T�U�ϓg�fw�OԀ�݉��C��t�s��`a�7%M���:��+.�~h)���-�@�9��K��W`�=Bs��y���  �  "�^���Y��\K�O�5���������ٽ�.������ػn�?E���%�.�����6A���/�V;�e�/�AKR��D�f˛�Dj�����>��or%��5>�Y�R���_�Mb�ȴY���G�,00�������]콫��N���s�ǽ%�ת>���S�w�`���c��C[�m�I���2��c��� ��8ս-ܯ�2?���Dq��J���-�~����j� ��g*���E��k�a��n��:�Ͻ����|���8/���F�#�X��|b�zXa�ĒU�>xA��4)�������l�N���0��k��-5�d�N�v�b��]m�Vm�'8b��O��E7��-�Ջ�|��c����5���Ru���aj��Y]���Y��x`��p�����N��3o��\�ǽb;�I��\���R9�	�R�ETi�*4y�B����z�aDl��nV�W>�z(���ܜ��@�3�(���?�_�Y��<q����p��EJ���[v��a��PH��`/����m��T���н3��t�������:����x㤽����Ѵ���Ͻ[��S���zF)��vA�LT[�
bt�����KE��׌������x��^*j��sR�`�>�x�2��.1��S:��L�\�d�<�}����[Y����������܄�~r���X��@���)�����ZU�����]1Խ�?ʽ��Ľ˜Ľ !ɽ�Xҽo8཯���}��y���&���<��'U��n�*1��\Q������}��Պ���a��,h��QP���=��r4���5�=�A��U�2kn�U���̌�c����(���d��@�����j���Q���9�c�$�:]�l6����e}⽟�ս_�ͽz�ʽ�I̽��ҽ�ݽ��p/��H��{�)2�"I�Tb�)�{�����������#���~��>e���N��?��39�7>��:M��mc�A�|�<ʉ�K푾�  �  ��}��ew�Qe��8J��0+���(a߽�|���-���mW���+��}�`�lټw�Ӽl�߼,R�����{�8���h�!c��^����=e�5���S�,um���}����H�w��c��zG�\�*�c�������Y�
����).;��:X��p�H���7���w��b�y0E�!�%���n�׽�8v�� �X���0����B��󼍕�F%�ӿ��2,��SR�p1��|�� %ѽ��CR!���@��<^���t�䔀�5����r��_[���>���#�B��qW�����v��.���K��Bi�1���B��E���\Z}��\e���G��Y(�*�����̺��R��W���Eg�2R�>�F��]D��J��QY��q�'������� ��]����g�'��F�1�f��D���4���W���ߌ�5T���o�y�R���8��'�� �'$'��C9���S���q������J��F����������fu�s�V��7� r�O��@���HŽ	n�����>������O���љ���������ýP^ܽ�b������K-��K�Hk��������:R���{������ ��ŀ��e���N���@��~>��I��:^��/z�ȋ��<�������Oś��吾Gq���0e�!wF��6+���q��I���ս��ǽ�����l���쪽��ƽ�\ӽ,�潡h ����Ԧ'��TB�*�`��5���X��s�����*9��La���~�xCb�G�L���A��BC��Q�M�h�����������:T��TR����������DP{���[��;>�9�$�]������D� �ս��ɽ�½XϿ��D��qǽ�Fѽ���.���$�	����u4�B�P�S�o�v���룕�P���=������T���_��\�y�W�_�UFM��[F��.L��]�X�w�a��P̗��8���  �  ����5���Tw��Y��6������Y��J��!cL��x�������ռ�R���C���0ƼY��cp��	,���^�����[������(���@�Ԁc��-���Q��}��H��ǭu��GW���7�X8������	� ���q+�%�I��i��c���������ۅ�z7s��R�2/�+���ZܽgE���X����L��y#�Lz��.켍�ڼ`�ټ>��T�~��HF�w�}�U�� �Խ�G�nV*���M��
o��Y��\@���ꊾt���m��M���/�������������:��9[��w{�"i��@���:��eC��=du���S�|0�/v��3�Ƹ�Mh���X{�&�Y�0�D��:��8��>�U]L��c�����M��\���'9����|�-��XQ�!u�<��&p���"��;t��>����ih`��D��y0��k)��g0��:D��Ba�������'Ś�5ƞ��P�����'��p`a�l>�:��,1���޽ʿ�x䩽�^��]����⎽N7��)���c��Un������S׽u��p��FW1��R�/�v�Vٌ�5s���Ҥ�K��|t���o����� �r�7&Y��I�WYG�A�R��j��\���|��e.�������ګ��ť�6���^3��^�n�L�v-��C�t� ��佭<Ͻ��1?���۳�ڇ��<?��YS����̽�u�4l��g���)���G�ͺi�����X���7���"��4ɪ��E���:��ys��aVn���V�ܖJ�@L��i[�O4u��\��晾���q��;䪾����Q���*�����c�U�B���%�R���������l�νýU@������,���{���ʽ�%ڽr��������b7�zW��Lz�uꎾ����	����_������������:҃�(�j�
�V��O�.U�6�h�&�������\��\����  �  ��!��4�������nн/ӣ��av���1�J���dk����Q�5��������`�u:K��^����Ȼc����z�2I��f����G�Lg��������߽���xn�1�"�i%��0��\����d�ֽ@���0��N�������'Ƚ��e
���,	%�t�&���������PF˽:����Jq��0��W��*x��ory�.E3��E��+��a�� �d�+�{�m�!�����D;)�(h��@���Žl?�,�����F&���%�k���:��{��d�Ͻ����S)���ک�`n���Q�������~(�R�0��0�=�&��'�^p���ֽ�6���#��{4X��[,�PL����w�ټ�ϼ��μIټ�)�L����=��.h��6���=���wܽp��A<���.���<���B�ݗ?��[4��]#��>������F潲޽�B罰% ��X�_�&�;w9��F�ĮK�I�G��X;�,�(��]�����޽ҽ�㰽%@��>���%�i�ՉX���N�"]K�DM�ެS�}_��Pq�m��A���Ʈ�-3ͽ�y���K�%�#�;���M��zY���\�n3W�NJ�=b8��%�P�
�����?���!���4���H���Y�@�c�:�e�:^�0O���:��$�-��3'��\�ս���T2���՛�
쒽q��g���ф���Ќ� ԑ�|-��Zڦ�*����ѽ�3���s�!��8��L� �\��	e���d���[�~�K��8��%��(�ִ����*�-!*�ѕ=��P�,e_�G�f�NPe�.[�.J��5�3��3�	�Op�н�湽�^��������������� ������`⛽.٥�~��A�Ƚ>�*��z���-�}D���W�?Pe�U	k���g�<?\�Q�J�c7�v�%�P�լ����+�$�|%6�R�I�P
\���h��  �  A�x��^���T��-M˽�����s���0��c��#^���[�.d�V���t�����s�|Ֆ�n�ݻ#^*��Y����¼�T�EeF��h���*��ͨڽ�3�{k�EE��� ���m������Gѽ7���J-���������	ý�N罶�����Z� �
"�f��g����ǽx�����n�l0�}����ᵼ�⁼��=����=u��C���)S�M6�Cx��������j5)���e�Ɨ�6m��M��!
��X�{�!��>!�����|	�&*�ʽ�l���M��_�)���r�ڽ�^�N���5$��O,���+��"���������0ӽ^��vW����X�	.�������e+߼|#Լ��Ӽ�޼�H������T ?��#i�q֏�N���(mٽcs�m��+��j8��>��#;�U@0�e��OB�.��F ⽸=ڽW/�7��� s��N#��r5��>B�3.G��UC�o{7���%�-��Ͼ���ѽ0u����������2al��,[���Q��M��O�,V��	b�r�s�����Y��� ���t̽�p�����"��)8�U�I��U��6X���R�d)F��4� #�+��&���	���P@�k�1��2E�m�U��~_�-a�x Z�A�K��8��z"�Y�����Nyս;Ƽ�EL������=�����������ȋ�����%��z�����������ѽ��z�
���,5�kI�2^X���`��/`�CiW��H�T5�h#������������We'�F:���L�q[��Eb�U�`��W�ŹF��^2����X����н����6����T��g���⓽C[��}S��Xז��4��@�������pɽj��+f�]��{~+���@�A�S�� a�X�f��Rc��&X��VG�g4��:#�;������l,"��93�6uF���W�
=d��  �  �g����P�����_���r��z.k���/�g{��"g��,�|�1�/��0��ǒû�Ʒ�G8ֻ5��ؕL�������ϼ~t�+D�����y�Ъ̽h��E����O)�����R���㽭n��-���c��������������C�ս�����
����k���F:�n��Y���-A��;i�
f1� ���ż�ᒼɫ_���2�Rg����L�.��X�5��5E��;��o�*�Hja�+��������ܽg% ���� ���������kJܽ�ӻ�X(��AM���˚��J��2�˽g0�
	
� ����\Q��P��?	����ɽ⥽�冽eW[�~f4�U��r'���8伽g�x��6��I���'��F�}vm��������ѽ�n�����Xd �DZ,�Zb1��.�I�$�a��<��q/�dOֽq=Ͻ��׽��0<�mu��*���5�r�:��<7�K�,�0���
�\��
7ͽ�	��[������4�t�u�c�"�Y��U�(W���]�w%j�8|�������Uv��;9˽͋��F������.�U�>���H��uK���F��;��c+����_�'>�T���
�����(�4�:��I���R�kwT�I8N�eSA�� 0�E����	�1?��սsd��6��q^��tw��HŒ�1⏽5�����-[��'���`૽4}��xNҽ���x�P��c-��?��L��S�Z�S��yK��q=�U,�~������(��	��v�i����0��A���N��U��pT�O�K��7=�=+���������+ҽ�۽���������9��~ݗ�+;��>���욽Bv���P���#���˽<�㽰� ��!��K%��k8�(I���T���Y���V�h�L��?=���+��B��L�+3�����X��*� �<��L�B�W��  �  9���*e���1�}u˽�V������6�d�Lz3�6�
��Ӽ	���Jo���8�/d��8��g#��xL������߲��=�c���E�Q�y�Z���N����ؽ��� ����03������ǽ ԩ�Lܐ�W���;�}�]-��Pʞ�(����ٽn)�q}����s����)�˽���nɎ��f�(�7��9�H1�u��.��I�l��BS���Q�Qh����
ǭ���ܼj��L&2���_��ኽ*񨽬�ǽ	e你:������-�z����޽�����ॽY�I������\H���Ŵ��Խ��a��3��g��:������۽�w��Ŭ���R��~Wd��VB���'��d��8�X) ��u��m}������ ���7��T���x�p⑽�b��D�Ƚ�轥��N_�q�����5I����������bֽy�ĽZ���8ƽO�ٽ�����
�fe��#�j(���%����,�����Mʽ����Q/��1y���p��Ԁs��_h�Uc�1rd�G�k��x� ��5t��
��%����˽���k�������!�i�.���6���8�\4���*��-�&��w�T"�����������T��RH+�kN8�Gh@�"B�:Q=�;�2��%����(A�*���0ٽ]�Ž�ܵ�l���RF�����𻖽<��*P������ާ�ڻ����½�ս��U��>��"�8!1�c<��A�^A�%�9���-����d���q�_���� ������#���1��=��C��sB�4�;���/��\!�3���6�Ns콷�ֽ�Ľr�������ڣ�w�����'��&L��Cb��Ys������Ndѽ��������� 1���,�7.:�#�C�.[G��D���;� S.�8c�X��2d�1�� ��	"������-���;�Q�E��  �   �ѽ�SϽ�Ľnj��'t��Nڇ�g�f���A�Z� �`��<8Լ@驼�����Zm���c���x��խ��Q�͗�k�.�-�Q�E�x�Nӑ��	�� ��@νP&ؽ��ؽx�Ͻ[����I��x⍽��r��Y�.UU�of������������P�ʽףؽ��ܽ�׽�.ɽ��sO��Y���bcm��FI�9)���輷⿼����Y꒼�B⟼�\���"��
	���$�r�D�5h��ʇ��5��-�����ƽ�սC�ܽ�ڽ��ͽ�9��x���؋�ډu���e�i�k�"���k����e��ޤν����=�v��z7�<Kܽ��Ƚdг��f��(Ȍ�%�x�Z�[�V�B�"F.�����0���0�-0&�3�9��-R�p�n�����	m��Z����½"%ٽ�?�X(�1��8�	�s1����d��V�ҽ�����L��Mʪ�@/��w���9*ٽ<��#������(�\�z	��v�9b���,߽7&˽�$���H��Zy������A�����x���x��T��󇽑������'���HB����ѽC��-��ȅ	��_�!E�ں"��#����Ek�Oz�s�yJｗJ��~�O�v ��`�2�S$�7+�g-�1�*�ǫ#����o�[:� *��P�ὦ�ѽ�ýi����v���������Ġ��B��,�������n#Ͻ�߽���Z��O��A"�k�)�\1-��+���%��s��B��k�Ӗ��YK��콮���ed�ֶ�3��%o(���-�>.���)���!��������?�񽲘ཛTѽ��ý𖸽��������?��K�������vԵ�3����ͽ��ܽ���D ��
����\� �x*��`0��g2��t/�O�'�B������p�Ul��I������J����]��o=(��0��  �  "���ܪ�,���5p��"Г��8����x�`�7`F�.�+�i(���Aɼ{%��d����ȶ���ռ�Q�и���7��7S�|�m�8������M���䦽u����}���ۯ�7����X��u��ZBb�&B��i.�`	+�1�8�ëT�2z����ȥ��z,��2��᬴�Wɮ�Z�����,��j�F�j�P��4�g��4���߼P˼�ʼ�6ܼ���<��+1�NML�5�f�����>���3��e����s���������Q۰�
���!t��(�����a���G��<�w�A�~X��{������2��Iǽɗ̽=f˽T0Ž/ỽb��fѥ��@���F���ہ���j�^KS���?�,3��X/���5��.E��t\�˘x�Ig��{z��������_�ýH�н�Eܽ;���r뽑n�}��-ؽ�ǽ�t��B���������DF������*�����нS��<�������Y9 �����������ȣ߽Խ�RȽ'����l4�������6��p>����������\�������G½6ѽvu߽[�Y<���w�p7	�������\�E�w$�Z����4�q�ֽ�jν�'ν�3ֽ�_�w��������t�,���e��t�h�� ��m���c��z~�� 2׽Ŭɽ�����P���"��fˮ��T�����u�ǽ*ս9��(4�a�����9�
������>�����n ��[����c�����Sݽֽ4׽���Ƒ����j���7��$�2��\[�(P����ǧ��!��?w�_?彨�׽
˽��7t��1���ض��6���hǽ�Խ��A�� S��!�*f���6�����x��C�#������)W��-�彩��T�佭��5,��6�������  �  :-����������ȓ�{��۾���F���ψ��}�'zc�<&E�£&�����B��,D�Y# ��Q�d�0���P���o��儽ѡ���3k��6晽 ᙽ�:��`E���1�������i��6K��-�F�Z�Q���P��"�9@�+`��>~�����c����C���:���N���杽bƛ�50��6^������k�EL�7.��g�z��z-�r(�L�*��UH��g��?��:܍�"��ᚽC<���ޝ��������!���қ���>����h�pK��0�n��-��}���+��NH���j��T��{���y�����?೽1����������0j������Gx�����8F���́�|�i�_8X��R��Y�D}l�&���yЕ��������v½?ʽ;Ͻ��ѽ��ҽ�ҽ�PϽZ�ɽ���h��3䦽u�����j�����-���t&���6���j���O½�н�6ܽ���U�ޕ꽡6��A꽍*�{*���׽m˽Y'���*������/���Ӡ�!S��D󻽭Mͽ��ݽ�2�h���!��&1��I�����2�K� ��R��E����b�׽�_ʽ���!����߹�*f���a̽��۽��9[�����<E	��*����6(����c���M
� G�T� �ߛ򽫽⽽�ӽ��ǽ�����Y���Wƽ��ѽ%��6R����R�E}	����J����yX�n�O�	��i�M��j����ལgҽ�jǽ����N�½.ʽ�gֽ\�����S���\����E�'���8���y(����� ������սF˽R�ƽ��Ƚѽ�޽%��M���e��RK�=��/�<�y{����is�*~����|� 
�����*ٽ��Ͻۤ̽��Ͻ�ٽ���Ӱ��1���	��  �  (?]��v�5����'���J��$��s�������ɢ�T�������J]�+�;���%�����*���D��Ui��ň����ű�������Z��������ڗ��#�����jlg�azM�M�2���������ټoü 㿼��ϼXT�4��Y*��F��Ta�.p{�1I������vP����������*_���u��䧽W����L���b��(C�֜1�M�0��K@�N�]��ၽZd�����w:���ֵ����,3��h/��g�������"6�M_f���L���2��}������u伊�f��}��19��EX� �w���C�������*���z��a�ʽumѽl�ҽQͽ%���U+�������������z����\'���m��ܱ���@ɽX�ٽ�T�:���W�p޽&Խ�ɽZ|��p�����������"}������:o�
�c��a�-Di��?z��7��퀗�#��������ý�lѽ�޽U����`����3�S������/�ޟܽy+ʽ�t��S���W���Qɵ��8ĽW�׽0R�r �C��?�����5�
�D����@+�����ὒ�ս��ɽF)���������������6������'��`�ý7�ѽ�/�B����&��K
��#��;����I��v��Mk�|;
�r �|���ݽpս7�Խ�eܽV8뽕;�����DL�����`����N<�:K�ӓ
�8��K����8��⽄lսKXȽ�輽ʄ���`����������;��ˇ̽,-ڽ-�v���rC�P��j��Wp��E��I�������<a�g�	�����M����&�ڽ�Wݽ�������o�Q�����������Q��r�wE�ۅ����y�x:����轧�۽zϽ
�Ľ0���=��)���A�Ľ�Ͻu�ܽ�w꽙\���  �  C�?�1f��&��t_���ӳ�q�Ž:ѽ�ӽ�̽r�������{:����m�2�Q�h�I���W��x�`��������½|(ҽؽ�Խ�|ǽF���ğ��8��`l���G��'��f
�������ӛ�����F�����<���>ռ�{�![�(�=��ma�y��7������sĽ�`Խ��ܽ�۽��н�m���I��- ����r��v\��2[�1o��_���P�������νU�ڽ�ܽ�Wս�!ƽ  ��FN�������f��D���%�c���Q�ɼ�e���Э�����U�ϼ��������0�XQ��{u�󖎽�9��(����ѽG�彤^������v������d�ս%������]�����ൖ�����cH����ֽ���m�[��������M��k߽<$ʽ�͵�
f���#��������q�@�]��O��F��E�<�L�d�Z�,�n�������� ���+��0ɽZ�޽�k�������!��	�-��-�
��=����ZӽY�ƽA�ý��˽N�ݽ�@��~Z�#�f����5[�k�e��ok������éѽ �½������c�����_@�����䌞��X���氽�����<̽��ܽ���98��������!�#�(��-�#o,�s�&��������ֺ�����n��#��GR��R����Q�%�O�+�d�,�I0)���!�������.&�ٗ��޽�:Ͻj��ӗ�����w���	`������`T������6h���ƽ��Խ�+�<�����T�h���%���,�Rv/��T-�=h&�@��1����?K�������T �/�
��}��`#�3f,�U1��0�d�+��D#�����"����������]�Խ��ǽ��܀�����KR���O���괽���]�Ƚ�_ֽ����  �  )�1���d�y��eƮ��[ͽ�S�3���_��������b��ƽ�����ۤ{�c�q�XK��Z���V��"�Ͻ+���Y��^� �zR���e�=�̽��O����g��7��
�-����,���;�]�+�A�E>�J�R�T)�My��6�ϼ#g��[*�\`W��J���;��I�ý���g!��Ϸ�_�3���b�⽊�Ž����=������m߁���������½��߽W���������#����㽛�ƽS���hĉ�'\^�6�1��t��8⼲ķ�����m≼�셼�̎��K����ż�n󼒠�.&:���d�̋�}਽�Ƚ܅�܍�L�n&��� 	����P�ܽ2���A*��p%���_���#���YؽD���!�
�q+�����h��	���8��]ҽO⵽E�������@p�]�V�MD�8���1�_�1��7��D��
V�R�m��녽4N��.r����Ƚ�7����Fg����?L(��#+��{'�+�����1��W��T۽��׽A@ὦ�����	������'��W1���4��]1��X(�P\�i��oi���ཕ�ɽR��c���T���}�������*��������Y���٣��6��f���c�ҽ�s�,�L��� �tH/���:�JaA�p�A�Pc;���/��!��F��I�U������L'�x���1��-��:��@�(SA�Pg;��O0���!��y��~��:�H�սQ�½��2���k��ߡ��O��?���f6������u8��$ָ���Ƚ��ܽr����Q����hJ'��@5�Ԃ?�!>D��zB��w:�8�-����j���������*���@(��6�O:A��&F���D���<�X�0�;�!�3H����h��GٽȽ�����6���䨽 �����1Ǥ�xo����[���rmɽ��ڽ�  �  ��.�{�k�󝙽�7�� �����p�o'������bb��A.��LN��+���Z<��hg��йʽ[��@_�N���^�a����Q���罽�=���.l�&�2��T�N���������Q��
#���
������j�A���櫯���n�!��=W�=񋽗ð�Ci׽j����X�u��ۜ���u�Ὄ����^��>���l����⠽�]��tݽ1��rd����z��*��+�۽����6��ʈ_�~&*�� ��7ü�񗼺�x�{\���V��ch����[����Ӽ���5.�"(_�<���@ְ�Ǯ׽�������/��$��3#��j�1�f���`0׽�^��4ж�8�����н���/
�K[�'(��.�l,���"����|�@ݽ$��T���o�a���F�}L4�
)���#�}]$��**�rX5�#EF���]�9c}��"���嬽�9̽,o�O������.��9���=�ĥ9���.�),��W��z��X��z'轱�� �����(���8�ʑC�y�F�d|B��7���&�\����z�⽄�ƽ���N�������}���0�������Ȉ�Af��@���4����+���Ѹ�Yν&X�����V�i�*�϶<��K��kS�k(T�.)M�_�?���.�c��%������z���)��ڬ,�(�=�V�K��dS�LS���K��>��V,�4%������콘�ѽ�[��/���o��Ye���w��/L��^ȑ�j9䚽��������½��ٽ5_���=�@2�#t2��C�4�P� �V���T�\�K��	=�u�+����J��PL
�
����Y%�Ά6��G��FS�N�X��KV�E�L��:=�b�*�n��W���E�UԽ����=z���-��`\��p���T���Ν�~����	��;��� ½�ս�  �  E�/��t�_��1jͽ����B���2(�%���8�֓����ѽ+���6�X���H.���|����۽������v ��Z�} ������	ʽ⮟���r��q2��P�����Ny���/�4w��
׻٠ѻH���m ���_�����qj㼲��u�Z��q���ƺ��1�^}�I��>!��O"�w��%R�Q���Tν� ���鞽���k��jbʽj;�bL
�cd�E�!��!���{s	���꽭����<����c�Fu(�����0⳼BJ���X���<�b�8��<J��p�喼xü$3 �'Q)��^�����Wٷ�;Y㽀��*m��*�D1���/��3&��|����彔~̽�����Ƚb޽ ����&&�
j4�8�:��e8���-����cV�3�:���O㜽�ꁽ�I[�@�>���+��� �h����g"��;-�`�=��U�j�v��F��9���TgнW����Q��'�p�9�&F�eJ��F��:���(�����w�=����O���'�����;�2�ZD��P���S��fN�X�A�@;/��d�����彠�ƽ����t����Ԑ�//���������.ׄ��X���Z��_V���!������ "ͽo�N���U��2�[SF�Q}V��_���`��BY�q�J��8�n`%��9�4��k�����O#�>�5��|H�v�W��`�7	`�dW���G���3�j���	����y�н�y���A���*���1��Vu��@j�� ⍽�ᐽ淪��֟�[���8���Yٽ�;�������$��:��N��\\��?c��|a��W��dG�X�4���"�K��K��T�ε��
-�9*@��>R�}�_�ele�/�b�]�W��bF�|�1�t;��B�Q<�"�ҽҟ��l_���棽�8��n����u���ޙ��ٝ�bĤ�L_������o�ӽ�  �  ��0�,�w��V���Rҽ�\������p�ٯ"�`���=�o�����׽s��E��ʒ���_��Yq��P��a�����!�m�$����������	�νߘ��.�u�T3�����㮼oo�p[%�*�{�»�f��L�߻;��YuU������+༛?��g\�u������a�뽹�
���-�%���&�b��+�#9��n�ӽ�����ߢ�V⡽[ӱ��Ͻ���6�����D&��#&��4�;�z����ý:�����e��o(����i���6��7�M���2��%/��h@��f�����O���&���(�E _�}ّ�3���Ƕ��
�V&�\S.�K�5�qO4��`*�J)�t$���пн��Ž�̽:�����u/��s*�R�8�pN?���<�-�1�g( ���
���ۚ��Z���靁��zY�R1<�V1)��A�����:������*��=;��9S���t�>㐽���z)ҽ�/��j���*�{�=�:zJ��N�*lJ��
>�r,�Gb����_J�������{��#���!��l6�XsH�otT�MX�3�R��KE��N2�[�����i�+ǽ^&��������ه�����n��ᎃ�����������'괽��̽Z�뽯���;��4���I�'�Z�tUd��]e���]���N��b;�m(�Pw������h���%���8��FL��[�_�d���d���[�K�8�6��h ���
�q�ｸ�н?������Cݚ������+��b&������2����U������E�������ٽa������,'�ϝ=���Q���`���g��e�R�[��K�2�7��P%�@������X�
�4�/�K�C��5V���c���i�:�f���[�l�I�U84�e��8	����OWҽ����X&��w����雽aD���2��l�������Pr��`!�����(1ӽ�  �  E�/��t�_��1jͽ����B���2(�%���8�֓����ѽ+���6�X���H.���|����۽������v ��Z�} ������	ʽ⮟���r��q2��P�����Ny���/�4w��
׻ڠѻI���m ���_�����rj㼳��v�Z��q���ƺ��1�^}�J��>!��O"�x��%R�T���Tν� ���鞽��l��vbʽz;�mL
�qd�W�!��!���s	�>�����6=��
�c�eu(����b೼�F����W�8�<�r�8��"J�Q�p�і�b ü% �A)���^��}���η�CN����g�U*�1?1���/��/&��y��u�彡|̽�����Ƚ޽' ������&�>n4���:��j8�j�-����[��=�f����윽���W[���>�q�+��� ���F���d"�	6-��=���U���v��>���]нc���'L�#�'���9��F�`J�HF�:�x�(�?��u��;�������Ӱ���|�2�^D�^
P�ޙS�lN�+�A�0A/��j�ŭ���彍�ƽ����c��qې�	5���������gڄ�Z[���\���W���"�������"ͽ��g���U��2�`SF�U}V��_���`��BY�s�J��8�o`%��9�5��k�����O#�>�5��|H�v�W��`�7	`�dW���G���3�j���	����y�н�y���A���*���1��Vu��@j�� ⍽�ᐽ淪��֟�[���8���Yٽ�;�������$��:��N��\\��?c��|a��W��dG�X�4���"�K��K��T�ε��
-�9*@��>R�}�_�ele�/�b�]�W��bF�|�1�t;��B�Q<�"�ҽҟ��l_���棽�8��n����u���ޙ��ٝ�bĤ�L_������o�ӽ�  �  ��.�{�k�󝙽�7�� �����p�o'������bb��A.��LN��+���Z<��hg��йʽ[��@_�N���^�a����Q���罽�=���.l�&�2��T�N���������Q��
#���
������k�A���端���n�!��=W�=񋽗ð�Ci׽k����X�v��ܜ���u�ὒ����^��H���y����⠽�]���ݽ*1���d�/�$�Zz�>+��ڃ۽?��&7����_��&*�t� �}4üd뗼ҡx���[�6�V�j1h��凼4���lӼ:m��.�._�$���������׽������%�p�$�%+#�6c��Ֆ���)׽�Z��f϶�b����н��}5
�%b�/(�!.�`),�>�"����}���Tݽ�/�� ��I����b���F�v]4��)���#��]$��%*��M5��4F�C�]�pH}����Ӭ��%̽�Y�R�������.���9�&�=�3�9���.�+&�nS��t��l�콪'��8��Ɗ�%�(�W�8���C�dG��B��7�9�&�wg�� �N���ǽY%��� ��%��S����9��Y����Έ�.k��������.��	Ӹ�Zν�X����V�w�*�ض<��K��kS�p(T�2)M�b�?���.�e��&������z���*��ڬ,�)�=�W�K��dS�LS���K��>��V,�4%������콙�ѽ�[��/���o��Ye���w��/L��^ȑ�j9䚽��������½��ٽ5_���=�@2�#t2��C�4�P� �V���T�\�K��	=�u�+����J��PL
�
����Y%�Ά6��G��FS�N�X��KV�E�L��:=�b�*�n��W���E�UԽ����=z���-��`\��p���T���Ν�~����	��;��� ½�ս�  �  )�1���d�y��eƮ��[ͽ�S�3���_��������b��ƽ�����ۤ{�c�q�XK��Z���V��"�Ͻ+���Y��^� �zR���e�=�̽��O����g��7��
�-����,���<�]�+�A�E>�K�R�U)�My��7�ϼ$g��[*�]`W��J���;��J�ý���i!��з�`�6���g�⽑�Ž����=�������߁��������½߽����ы�1������̀㽋�ƽL���Jŉ�j]^���1��s��3⼫���kr��+Ή�!х�Ũ������ż},�y���9��d������è��xȽ�g��~������	�{n����ܽɠ���$��N$���b��+��,eؽ�����
��6�����v�o������{ҽ8����/��5����gp�W�NeD��8�z�1��1���7��D���U���m��؅��7���X���qȽ�P���W�Ax��=(�D+��o'����,���+�xO��P۽��׽�Dέ�����	�]��t�'�d1��4��l1��h(�zl�~����������ɽ���x���g���������������������7_���ݣ�z9��x���Ƥҽ�t�n�r�� ��H/���:�SaA�x�A�Vc;���/��!��F��I�X������M'�x���1��-��:��@�(SA�Pg;��O0���!��y��~��:�I�սQ�½��2���k��ߡ��O��?���f6������u8��$ָ���Ƚ��ܽr����Q����hJ'��@5�Ԃ?�!>D��zB��w:�8�-����j���������*���@(��6�O:A��&F���D���<�X�0�;�!�3H����h��GٽȽ�����6���䨽 �����1Ǥ�xo����[���rmɽ��ڽ�  �  C�?�1f��&��t_���ӳ�q�Ž:ѽ�ӽ�̽r�������{:����m�2�Q�h�I���W��x�`��������½|(ҽؽ�Խ�|ǽF���ğ��8��`l���G��'��f
�������ӛ�����F�����=���>ռ�{�![�(�=��ma�y��8������sĽ�`Խ��ܽ�۽��н�m���I��7 ����r�
w\��2[�H1o�`���P��T���X�νͦڽ��ܽ}Xս�"ƽ:!��lO��������f�xD���%�`�����rɼ�L������kӶ��dϼm���j��p0�D!Q��>u��u��'������ũѽ���;��9q��K���:��jyս��H	��W��/������t���5V��V�ֽ���z��������z��9�߽vHʽ�ﵽ����@�����¶q�6�]�0O���F���E�N�L���Z���n����💽U���)����Ƚ��޽�E�����H��b������|���
�O)������OӽZ~ƽ��ýn̽K�ݽ�P��!e�0�Bu����m����#���!C��h��t�ѽ��½1ĵ��̪�c��J��
N���������(_���밽����l?̽^�ܽ	�8��������!�3�(��-�-o,�{�&��������ۺ�����q��%��GR��R����R�%�P�+�d�,�I0)���!�������.&�ڗ��޽�:Ͻj��ӗ�����w���	`������`T������6h���ƽ��Խ�+�<�����T�h���%���,�Rv/��T-�=h&�@��1����?K�������T �/�
��}��`#�3f,�U1��0�d�+��D#�����"����������]�Խ��ǽ��܀�����KR���O���괽���]�Ƚ�_ֽ����  �  (?]��v�5����'���J��$��s�������ɢ�T�������J]�+�;���%�����*���D��Ui��ň����ű�������Z��������ڗ��#�����jlg�azM�M�2���������ټoü 㿼��ϼYT�4��Y*��F��Ta�/p{�2I������wP����������-_���u��䧽^����L���b��(C���1���0��K@���]��ၽ�d�����:��J׵�u��44���0������º���7��_f���L�f�2��w���$���O�������ޒ��9��X�sdw�p̊�|��Ц�����Q���ʽ�Fѽ�{ҽ�0ͽ4���3������b������z���1��7}��|ƴ�PZɽ��ٽfw�����C޽�OԽ6*ɽ�����۱�$������G���� ���Qo�)�c�&�a�:i��*z��'��vk������9s����ýFѽ�V޽	�꽰g���q����:��̟��'�o�ܽ�ʽ�i��Ӱ�������ϵ��DĽ3�׽�i�t� �����������
�<����V���6����ֽbʽ�C��/����Ϋ�굧�C��Q�������ý/�ѽr2��C���W'�7L
��#��;����Z�����Vk��;
�#r �����ݽtս;�Խ�eܽX8뽗;�����DL�����`����N<�:K�ӓ
�8��L����8��⽄lսKXȽ�輽ʄ���`����������;��ˇ̽,-ڽ-�v���rC�P��j��Wp��E��I�������<a�g�	�����M����&�ڽ�Wݽ�������o�Q�����������Q��r�wE�ۅ����y�x:����轧�۽zϽ
�Ľ0���=��)���A�Ľ�Ͻu�ܽ�w꽙\���  �  :-����������ȓ�{��۾���F���ψ��}�'zc�<&E�£&�����B��,D�Y# ��Q�d�0���P���o��儽ѡ���3k��6晽 ᙽ�:��`E���1�������i��6K��-�F�Z�Q���P��"�9@�+`��>~�����c����C�� ;���N���杽dƛ�80��:^������k�(EL�,7.��g�����-��(���*�OVH���g�@���܍�����ᚽJ=���ߝ����ץ�����/���>����h�)K�0���Nq�y���+��&H��j�s8��Ed���p���ɭ�;������|��NZ��wB���t��7W������.��]�����i��)X�oR�Y��l��τ��啽����<���&½�eʽ`dϽB�ѽv�ҽ�-ҽ�xϽ>�ɽ������n���Ά��������"��݊��N���%��&T��	4½[�н�ܽЬ�\+�j��
�D�!�U���׽�P˽q��aݮ����0��0��ڠ�x_��~���eͽ�޽U�����J��?G��`�i��:I��� �;z��8"���/ ؽKwʽ׫��E���l칽@p��Ei̽Z�۽+��^�����E	�9+�Ш�a(����{���M
�G�_� ��򽷽�Ɠӽ��ǽ�����Y���Wƽ��ѽ'��7R����R�E}	����J����yX�n�O�	��i�M��j����ལgҽ�jǽ����N�½.ʽ�gֽ\�����S���\����E�'���8���y(����� ������սF˽R�ƽ��Ƚѽ�޽%��M���e��RK�=��/�<�y{����is�*~����|� 
�����*ٽ��Ͻۤ̽��Ͻ�ٽ���Ӱ��1���	��  �  "���ܪ�,���5p��"Г��8����x�`�7`F�.�+�i(���Aɼ{%��d����ȶ���ռ�Q�и���7��7S�|�m�8������M���䦽u����}���ۯ�7����X��u��ZBb�&B��i.�`	+�1�8�ëT�2z����ɥ��{,��2��⬴�Xɮ�Z�����,��m�N�j��P��4�x��4�2�߼OP˼ʼ87ܼ�������+1�NL�3�f�R��O?��u4��y����t�����ʝ���۰������r��$���H�a�o�G�g�;��A�\�W���{�|g��쨽����7&ǽr̽t>˽dŽ���=�2������'��6���l�j�b(S�9�?�j3�V/���5��AE�>�\���x�q���R�������ȶ�+�ý��н*oܽ��彳��~�뽧��Hؽ�#ǽZ���*������ᕽA������y����н��R��������% �}���\�����꽮z߽1�ӽ/Ƚ�����w�����Mꗽ�+��9������)���z��������,���c½�Vѽa�߽�6��f����xM	�-��>���"���4��
��L���ֽHzνa4ν�=ֽPg�����������t�����e� u����!�����"d���~��2׽Ѭɽ�����P���"��iˮ��T�����w�ǽ+ս:��(4�b�����9�
������>�����n ��[����c�����Sݽֽ4׽���Ƒ����j���7��$�2��\[�(P����ǧ��!��?w�_?彨�׽
˽��7t��1���ض��6���hǽ�Խ��A�� S��!�*f���6�����x��C�#������)W��-�彩��T�佭��5,��6�������  �   �ѽ�SϽ�Ľnj��'t��Nڇ�g�f���A�Z� �`��<8Լ@驼�����Zm���c���x��խ��Q�͗�k�.�-�Q�E�x�Nӑ��	�� ��@νP&ؽ��ؽx�Ͻ[����I��x⍽��r��Y�.UU�of������������Q�ʽأؽ��ܽ�׽�.ɽ��tO��[���gcm��FI�B)���<��⿼*����꒼�⟼p]���#�O	�|�$�R�D�Sh�vˇ��6�������ƽҒս��ܽڽ\�ͽ08�������Ӌ�}u���e�x�k���������P���ν(��|�pr��j&ܽ˲Ƚn����D�������Ux��v[�Y�B�*'.�t���������7��@&�o�9��QR�o�0���F����8��\�½Jٽeｱ:����u�	�@�"�����(�ҽj���3R���ʪ��*������0ٽ=�������k�qJ�����c�D<��߽�˽8���,���a�������2��\�~��x�E�x��Y��t���젒�?������k_��x�ѽ1<�T��y�	��s��X�{�"�v�#�j��my�������[��X�Q���W�� �;c��3�� $��7+��g-���*��#������u:�)*��o�ὼ�ѽýu����v��������Ġ��B��,�������o#Ͻ�߽���Z��O��A"�k�)�\1-��+���%��s��B��k�Ӗ��YK��콮���ed�ֶ�3��%o(���-�>.���)���!��������?�񽲘ཛTѽ��ý𖸽��������?��K�������vԵ�3����ͽ��ܽ���D ��
����\� �x*��`0��g2��t/�O�'�B������p�Ul��I������J����]��o=(��0��  �  9���*e���1�}u˽�V������6�d�Lz3�6�
��Ӽ	���Jo���8�/d��8��g#��xL������߲��=�c���E�Q�y�Z���N����ؽ��� ����03������ǽ ԩ�Lܐ�W���;�}�]-��Pʞ�(����ٽo)�r}����s����*�˽���oɎ��f�.�7��9�\1�(u��O����l�CS��Q�h����ǭ���ܼ����&2���_�A⊽��g�ǽ�e�W;������-��y��r�޽����5ݥ�������o���k<�����W�Խ���fU��&��Y��+�u���u�۽�Z�������8���)d�b/B�t�'��K�>'�� ��q����U���!��8��U�v�x������}��P�Ƚ�=����Zn���2��3U���������kֽ&�Ľ°��Vƽ&�ٽG�����
�;[�&�#�(� �%�tw���������ɽ3ܱ�����e��Ha��Ris��Oh��Mc��rd���k��y�i������4���,��O̽����������!�`�.�)�6�K�8�q�4�=�*��7��.��.������/��p�Z���I+�gO8��h@��"B��Q=�n�2��%����?A�M��
1ٽp�Ž�ܵ�u���YF���������>��,P������ާ�ۻ����½�ս��U��>��"�8!1�c<��A�^A�%�9���-����d���q�_���� ������#���1��=��C��sB�4�;���/��\!�3���6�Ns콷�ֽ�Ľr�������ڣ�w�����'��&L��Cb��Ys������Ndѽ��� ����� 1���,�7.:�#�C�.[G��D���;� S.�8c�X��2d�1�� ��	"������-���;�Q�E��  �  �g����P�����_���r��z.k���/�g{��"g��,�|�1�/��0��ǒû�Ʒ�G8ֻ5��ؕL�������ϼ~t�+D�����y�Ъ̽h��E����O)�����R���㽭n��-���c��������������C�ս�����
����k���F:�o��Z���.A��>i�f1�%���ż�ᒼ��_���2��g�b��ԁ.�kX��5���E�������*��ja��������� ݽ�% �Ǽ�6 �����"����Hܽdѻ��$��&H��Ś�B����˽�#�
���|��pG�5F�>5	�v�FlɽfΥ��ӆ�R7[��J4��������z���d�t��?��X��'�2F���m�`���6/���ѽ���΍�o �}d,��k1���.���$�q������5뽶Rֽ�=ϽÎ׽E���7��o��*�t�5��|:�]27�v�,�!����
�+��*#ͽ����i�����M�t���c�6�Y���U��W��]�31j�nI|������+��톰�L˽o���Q� ��M�.���>�f�H��K��F�F;�2k+����d�SB�cW�.�
������(�;�:�ĴI�-�R��wT�8N��SA� 0�[����	�L?��ս�d��@��x^��yw��LŒ�3⏽7�����.[��(���`૽4}��xNҽ����x�P��c-��?��L��S�Z�S��yK��q=�U,�~������(��	��v�i����0��A���N��U��pT�O�K��7=�=+���������+ҽ�۽���������9��~ݗ�+;��>���욽Bv���P���#���˽<�㽰� ��!��K%��k8�(I���T���Y���V�h�L��?=���+��B��L�+3�����X��*� �<��L�B�W��  �  A�x��^���T��-M˽�����s���0��c��#^���[�.d�V���t�����s�|Ֆ�n�ݻ#^*��Y����¼�T�EeF��h���*��ͨڽ�3�{k�EE��� ���m������Gѽ7���J-���������	ý�N罶�����Z� �
"�g��g����ǽy�����n�l0������ᵼ�⁼�=����u������oS�pM6��Cx����,��5)�
�e�IƗ�pm�����C
��X���!��>!�����|	�K)�7�ʽ�j��GK��������ڽ�[�����1$��J,�׭+���"�"�������%ӽ;��)N��	�X��.��������߼iԼ�Ӽ޼�R���}��e?�43i�Zߏ�.����wٽ�x��9+�Cp8�~>�*(;�,D0�����D�x���!��=ڽ�-�4����p��K#��n5��:B�C)G�NPC��u7�9�%�}��ٳ��|ѽ�k��ū�������Ul�$[��}Q�b�M��O�</V��b�f�s�l����������e~̽G{�@����"��/8�6�I�3U�E<X�i�R��-F���4�O#����Q���	���VA�,�1�{3E�ˇU��~_�Wa�� Z�U�K�8��z"�Y�����XyսCƼ�JL������=�����������ȋ�����%��z�����������ѽ��z�
���,5�kI�2^X���`��/`�CiW��H�T5�h#������������We'�F:���L�q[��Eb�U�`��W�ŹF��^2����X����н����6����T��g���⓽C[��}S��Xז��4��@�������pɽj��+f�]��{~+���@�A�S�� a�X�f��Rc��&X��VG�g4��:#�;������l,"��93�6uF���W�
=d��  �  t󤽭ɟ��搽b�u�3�A�ʸ��p��.�G�����f;���;�<�a/<��<<��><��5<6� <%��;�J�;�*��\�6y��s�޼��"��=Y������⛽eW���������_���#��BQ�o�*� �����W����@��Pm�����R����}��XK�����9ǔ�k�y�lqD�����\��7"e�r�ӻ�jw���=;}L�;���;��;�2�;��;��;��T;� ߹c!��3\U����VE
���>�q5t�`�������ʯ�󱯽ۀ���p��Z�z�V�O�mi/��Z ��&���?�z�i�;�h��2����Ľ��ý���i��Ս���g��86�� ���мo+���3s�)�F�Le/�u(�'�-���>���Z�d��蟼�ȼI&���"���N����6,���W��M�ν;�߽{"�m�㽱׽�|ý�A��A0��ы���5���;��=�������=�˽^i⽮h������v���G��нdd���c��o���Tb���B��x+�X�����u������k5��P��)��v9�m�O���m�]����%��}���tn׽1���8=��p��r
�U�ޯ��6ܽ\Pʽ�ӿ�����OȽ�-ڽ]�h��������i��J��[��)���3�޽��ĽiŬ�[䘽�R����{���k��+a���Z�<�W��W�~+Z�V�_���i��y�F�������1 ���h��|�۽Ш��4��u��*���Ծ� v�L#����Ὠ�нO�ǽ�ɽ�eԽ�罹���[�
��h�h��������#��C���ڽ����e���K���~��k�����s��k��g�G�e���f��#k��r���~��R��Yݔ���������]ӽ�]���3��k�����	�<V�$-	�R��1Y��׽`Mҽ�0׽߄彡���>	�M��fP��  �  *��������U�� n�X<�)��^x��ҧE�`	�� E�:dN�;-E<�=)<="7<�%9<@�/<�<b��;J~;}{q����҃��(ڼ���G%S����,���$��G\���^��`����w��J�[�$����G�	�����p:�g�e�k��������/����������@t����r�Dl?�2��p���d���ڻ��c�#;�;ߡ�;1��;���;�;)��;ɯ:;��J��aû�^U�����Y�T�9��m�jq�����녪��d��z��.����s��I�]%*����g0!�z:��;c����ס�&�����������Ma���
��;����lc�j�3� 5
��vѼ�Y���Ky�2pM���5�!�-�jA3�J&D�:�`�χ�����# ˼M' �"z"�`�L���}��i��c���yʽ��ڽ��Ὀ�޽�:ҽN6������G6������ф����8ٙ�l����ǽ�ݽ:9�ހ�c｡��7ͽt���/���bw����a��C���,�J���|�����+�Zv����h��[�*���:�l�P��n�s���vo��RYԽ(�^����.�
���E� �_���ؽ7wǽ
P��������Ž�׽5��T|��F�E�zO�1�z���9���rܽ��½�	��(Ә�Z����}�KOm���b�;T\��7Y�W Y�d�[�c�a�ˀk���z�m������,Z����qHٽ�K�ʇ�(�� ��oZ�;�K8��S����޽�ͽ|QŽ+�ƽ-�ѽA:�!����_����]�U�������ģ���׽m_���詽i����*\��x�u��$m�K�h�*g��dh��l�)bt��3������s/��e������	�ѽ��뽻��@��p���6��h����-����4^��$ս��Ͻb�Խ���x����wo�����  �  ����V���;�4QY���,��r������kC�����D$:���; l�;��< �$<P'<Ջ<�<9^�;z�.;B���%�����ͩμ�����B��Lo�@��"���kR��Pԑ�8r��F+`�9a7�����X��������
���(�~�P�y3z�����A��-������r����_�9�1�x�����_�f�D����}�:^�w;)��;(��;��;n��;.s�;�>�:�'����޻�(Y�@��������,�i%[�S���U��������y��/b��d����]���7��"����Wm�s+���P��}�W锽f@���ү�A	��I���▽�.���W���-��~��Լ�������DQb�J�I��q@��D�V���s�R��������Ӽ7���,"�E^H�qt�� ���z�����s̽r�ҽ��Ͻ�uĽ!���~������ض��<�{�����֜��:����軽})н-�޽h��K%�4ս��½���������(��Va�)�E�j1�g�"���l�����-��&���#�Ę/���?�K�T�$�o�6È�Z���-᳽� ̽�㽼0���O��3��� �@
��'��*Ͻ_���(��ƚ��5���0ν����v���=���
�����=��� �;�콜�ս�����n��%���Q��x݀��xr�*�g�Ua���]�{]�[`�B�f�w�p�0G�������z��� =����ҽH��N��������|#�u������H�սAƽ�a������u�ɽ��ڽU�ｩ��M�	����I����ߙ��3齹ҽ
:��( ���2��5댽�у���z�*r��,m�ȅk���l��xq��y�MÂ��-��艖��O��x���ͽ=K�8Z�����^��Ʒ�U�[
���"���ڽ�ͽɽ�lͽ�Fڽ)�����
�|U��  �  �Nu��1o���Z�xq<�%u���,2��fL��һ�ͺ��;!�;n��;��<�<�.�;h��;�Jl;^��9����;��Q��~�ür#��R,���P�qgn��p��sT��0�x���_��!>����n����Լ�hμ^�_�1�H4U���s�/\��^b���\��f��E��� ����ꬴ�c�v��F�t���
����c�:�gW;kc�;�;�`;ST�:� T��΋�����j�ƭ�>��%��]B��\d�Ν~�:�������0{��{_�`�=�#*������{������)5�Z�\�qɁ��/�������ݚ���D:���Sm���I�~Y'��	�'�߼�����b��� n��b��e��|v��#���,��?7��Zz弼q	�R�$�	 E�<}i��>���j��y���ݷ��ͼ�����$���3��~Q�����m��xg�Нq��C��o喽�o���@���ɽ��ν��̽ý�g��9뢽~�=��S�c�/1L�\�9��u,�	#��x�,��-��10#�"M,���8�� I�	]�H?u�i$��y��X�������G�ӽJ��h�T�.���]ེ�н*����9��|f�����x�������{ ӽ������ë���� ��r��dG��߽�ͽ�~��5������@��p���A|��$q��i�8�e��e���h���o��sz��d��q���E�������1��©ʽ��ݽǵ������O��� ��`�����jٽ�0Ƚj˺��򳽈���꽽��̽��޽�_�a��K��XX�'������Foݽ��ʽ�	���0��{ݛ�e��w���5��m1{��u�2�s��#u�N>z�<|�����=������v���u��e�ǽ<�ڽb_�{���������"������^]޽�,ν&�½i�����½Z�ͽ�4޽i�𽢜 �����  �  �*C��@�4v3����&��N�ּ���;�o�+v�[����b���:\�m;y��;8ݫ;��;�H*;��0��+q�������L��ґ��y¼Fc��'��x0��E�8Q��9R��CG�"�1�����}��������d�������d�ݼ����)�MuC�a:T��jY���R�`B�c+��V��,񼼙�����R�<
��G�����'8��:t�:�\9ծ�c�������J����^᷼���6���)�	A���R�1�[�q�X�u�J��3���[����QӼ¼��˼)��Y�r�5���V�H|q�^뀽�����D~��lm���V�:<>�I&���_����2׼j躼L��ƅ��l֊�7 �������ɿ��߼���+��-��G��Gb���~����������Ҡ�kƣ�ؠ��m����s�|���c��_S���N���W�;m��e���ܕ�����j>��<䵽�j��N{�����c�������� ��X�l��Y���I���<�2��+�(��)���/���9��H���X��=l��Ѐ������������{����rýA�νD{ս׽l�ҽTɽ8¼�����k����~��V���������dX���н��ݽ!c�,G��%��ݽh{ҽe^Ž���>����_���g������������v��@r���q��v��d~�$��$������@垽s���=]��֤ýK�нv�ܽ��� 꽈�轵�b�Խ�]ƽ�"������n��"a���ï��$���˽��ٽM]彰��j�콚��E1޽Sҽ�Ž�A��D}�����YΘ�'ʐ�� �����D������׀��냽�������[×� ����q��a4���&Ľ~�ѽ�߽kc��|���!#����ڽ�X̽����.����@��B����徽>�̽�۽C������  �  �t����-[�2��>���8ؼ����&��qV|��F<�����+��l1��N�=:���:1/�8�$�w۷�#X�ASb�`O���T��fZԼ��󼖻�!��h���
$�� ����e����ټ+��#���X���P�~	s�.`���]ʼ1�����g"���)��)�I�"�2���
�������ؼ���ׂ����p���/�5��H	���vD��C?�Ǔ��m=໣)�ߞi�����Vf��/�ռ2���������"���*���,��z'�m��W�)��Xs���4����2��i���伨�`z)�1�@��P�oyX�JEX�U�Q��G�L;�3.��� �����T���RѼA���q���
d��=����˼�3꼐m�s���e.�WA�H�R�4�c��Nt�Ӝ������\D��/����⇽O����/m��W��~D�8��'5�5�<��lN�'�f�/߀�����⒗�T�����������̙�����Wf��U����I��q�]�b��kT���G��>��89�:���@��UM��]���p��2���Ӌ�����흽�����������»��Ǿ�A��ع��������ޝ�2�������YZ���Ֆ�=�����p�(KŽ�mͽ�}ѽ^�ѽ�-ν=�Ƚ�����E��n���,���:i��X��������[�����#����p�� /�����f����ј�Q7��Zq���e��M%��b�����ǽU�ͽ$�ѽ��ҽ�Ͻ��Ƚ�����̲��~���Ğ�3X��X"�����᪽9ݶ�#�½U�̽�8ӽ4�ս�oԽOJн^Sʽ�pý�-��@����
��N������H��x���+5���[���v���j������{����#����������7��Ž��̽
�ӽ�hٽ`�ܽlܽ;ؽ<н\~Ž�ǹ�z;���姽�D���짽�f��;K���ƽ)$ҽ۽�  �  I�ҼR.伜�����i������~�u�ټ1
¼ r��p�{�*12�����ї�Is���%���	�voP�����ᵼ<7ּ����(
��6�n[��W�v�������jԼ)����T��W�S�=��v��ݻ%���>��e������\�ϼ�p��t�$�	�����?�������`������5޼�����s����a���'����?#���"�6�Z�5R��������ڼ�X����8��o&�:$�GH�-G��_�����G�޼BM��ڥ��#�x�J7M���=��0O��c��{�����ҼY� �L����&�ń3��<�4>A���C��}D��{B�F7=��
4���&���4S��N�4�ۼ�~ּZa�؇�������&��<�/.P��_�%�j���q���u�I�w��Zw�zt�OIn�`2d��ZV�;�E�JG5��"'�(Z����z�#���1��SE�Tn[��q�����YV��{������u���JE���쓽�@��]ߎ�J����_���5t���c��sV���N���N�v�V�a1f�pz��_������J��[\���J���r���J��g���魽Oa��b���룽������a��&Z��{D���넽�p��_?��/��Yȥ�Ϧ���Ƿ�ӵ��i�����ý�ZĽ�
Ľ�½~���=�������.Ǫ�y���ٗ�^����X�����ˏ��ɖ��ٟ�n����j��u���sϾ�.½��ýXTĽ��ýY½�9���&��'���>���Ơ�.����S�����/���`/��tӚ�VJ�����(���q���ý�!ƽ�ǽUȽD�ǽ�7ƽ��½j����G���i�����i���o����WV�����4����W��.$��;Ͻ�]�Ľ�NɽD2̽@�ͽC ν��ͽ~�˽sȽ}½⺽�ᱽf����|�������i���堽"f��:��b��TŽ�  �  @y������Dּ���|��h��}��U�J��� ����ʼ����f���1���#�λ?��v���~���޼���߈����o� �� �G�����A!�.�ͼ�k�����Be_�T�Cʻ��^�r|꺘Fκ�7��̭�����{Q�R芼*}��f�̼W켼z������ �jD)�,��a'������r6߼����WЊ�Kmj��h�����m髼	ڼ�������&��O,��_*�Pb"�1�����P>��n�ּj�� Ϛ��7y��@����ua�I!ֻse���w$���a��;���޾���缏��Q\�q_,�Ք=��kM�ǗZ�F5c�pLe��_�wDR��*?�ԩ)�v��;�����	�����P1��@L��Bf�xp{�2���{F���0���F��?@y�'Bl�}�^���P���B�� 4���%�hp���hG������=Y�%6)���;��HO���b���t�AH��Ë��֓�i���Р���o���V������K�������r�3h�b�f�&�p������@��CЛ��9�������H��>ø�ʶ��h�������d����d��_����䋽B��/�~��Xv���r�_t���{�'��T5���4���^��u;������𴷽.q��J�ƽC�̽�ѽaҽ��ϽlMɽ�`��ꆳ��§�O<���Ƙ�Ut��T���n������꽽xȽ�Ͻ�
ҽ�1ѽSMͽ�lǽ�����'��ܛ���٩�]С����"����ˊ��Ʌ��`���烽vT���8��)Д�&=��Vϥ��*��I?��t ����Ž
�̽�ҽ+lֽ��ֽ�@ӽV�˽�a��맵�ƻ��>����4��Z�������4��oQ��oʽ�ӽn�ٽ�`۽��ٽ�$ս�Ͻ�Ƚr����c������2���Ұ��?%���瓽)я�z���������i'���3���ѫ��j���  �  m�c�����B-ּ6d��� ��D6�r"D��4G�mK>�!�*�|��c���-���̅��;��j��5l�������5�^H��O�#FK�ـ<�&���漍���i���iA����������}�SW�:i�;cd&;"�:M�Ĺ ,T�KA߻��3��р�����u�ݼ/[	�)?$���<�zP��AZ�T�X���K��4�м�����Yż���P����A���!�d����1���I�{]X�$[�6QR�>@��T(����b�vָ��펼��U��q���̻���2�{�&���f�_m��2��m�P��f�������`��B�b�(���E�.,b��{���������܈��c��3Ik���O�?i6��?$�՜��e$�`�7��T��^u��C���T��� ������Vq������D��Vm��U�9?���+�)O�js�e\�h1�������<w���F�'���$���6�c�K�G�b��Q|�f܋�?����t��!���~��{��1�����jJ��ƒ������d���C��*݅�AY�������.���⿽A]ʽ
Ͻ�ͽ�Fǽ�#���1������ߐ���s��t���~���r��=i��4c��a��Cc�!�i�r�s��ŀ�刽����A��O������}V��=�ν۽�佫k齐��|�Ὅ)ֽ��ǽ~۸�)ܬ���������¼��a9����Ž�qԽ[���罋f�A�-)ܽ Bн^ý��B���q,�������T��#:������|dy�k�u���v��|�󳂽����ᐽٙ�M�������<��;�ɽ�׽���B뽹��,�����V׽��ȽC������8���^���˶�W�ý�ӽ8k�eb����������սǵȽ���9���Z���b�����N��~��z�����^���ъ��6���1��2t��$䨽�  �  =�A�3۟�������>��=^���r��oy��Gp�w1Y�̬8��6�o���¼�z���B̼aZ��� �$-E��Be�t�z��ɀ���x���b���B��2����}���i����%Vp��=	�
�/;�ȓ;R�;���;�8�;z?L;V:v,:��q�ovQ��V��5��ޕ�n�;���^���z�zQ��L�����|�!�a� �>��������(�ܼ��ڼ����.���:�9^���z�}��� ��)�}�$Nc� �@�Ʃ���;v���p����h��MG#�����9���9���)>"�����m����]�]y��AӼH�	���.���U��Z}�]4���0������D7�����@P��� u�5�U�?�%k6���=��T�ƛv�H͎�_,��L����� ��Ǭ�2˞�C���lw�[�T�n87�_��a���{��k�>tټ�sԼ��ּ׏�#e�����(��O'�|�>�@�Z�ڛ{��M���٣�h�����ƽ��ѽx6ս"1ѽnQƽ�ض�r���h��76��"���꒽�n��$���4.ƽ�l׽�H����Nc佀ڽ�	˽'���+�����\z���-���n�@]b��Z��tU��cT�ܽV��i\��ie�ƹq������[���/���k��Y���iǽ�\ڽ<�������� �C� �tn��Ԥ�$۽�_ɽ�亽ȗ����n���mnǽ��ؽ
������L� ��� �@�����\ܽ��ɽX���$J��Oi����4��W�|�֨r��Fl���i��Lj�ån�a�v�����̈�V����֞�����X⾽'�ѽn��]b��<� �������������A۽܇ʽ�(��˪���2��OŽ#
ս�J罸x��F�����=��98 ���R(�c�ͽ���@����۟����z��s_������������z��能F������Ç���/���  �  ?:�M���o���v�.��I\��n���U��7����������֞[���2����� ��?����X��E?�Oi����O#��M����Ր�#ۂ��3^��1�V��������\��ػ+��;�L�;���;�t�;S�;L��;�+�;��A;� �t���=�x=��ۅ�q�$��5S���~�F���o���������������`�T7��;��U��R�7e�q=3�:�[��
��S^���z��,���:������@�Y�A�+�c����	��b�^�}���e�M��O9�E��:7�;H�;	z�:Y�6�H��wٻ��9��+���s̼�!��8��h�Q������r���j���-���8�������A����o�݃U�zK�+/S��l������ݟ��ô��iĽ��˽ʽ@[���֭��k�����$Z���5�I��\��d�1�Ҽ�ǼxļpǼRм��߼������
�'���u8�A�X�s���p��<N���uŽSٽ�d�J.�8��4?ڽ�HȽ2���Ȱ��Y阽u���ҝ����;���ؽ��뽣���Rn��X������ؽC�½B(���e���݈�
�w�#1e��iX��}P���L�L��}N���S�
$\���g��w� 0�������\��yb����ν@/潾������(y������M���'���@׽��ƽ���R���?Ž
ս�7齀���~���������4�N�������ѽ�x��������� ��m��t�r��ri�/�c��ha��#b��e�DBm�qnx�!���厽L��������ý%�ڽ���ZJ�\�
���B��MH�F�����|�׽8_ɽV
ý�Žjsѽ�}�Rv��#��[�����D�&�	��| �뽫-Խа���
��Wߜ��0������P���$7}�v�x�e�w�6�y�T�~��΃�Q4��(��� ���  �  �=��o��z�	�a>��Yq��B��纜������h���
��%s�%rF��8�q�oi��'�
�Iy)���S��Ԁ��ڔ�=�������#���B:��sr�Gm?�y��1���F�\��2»����{�l;]!�;���;lP<�<�<���;�f�;�t8:
э�Z7�Q��ɨ���s0�ѳd�����H���j������E ��t���JCv���I�
�%�6V��<��"��oE�,]q�ӎ�H���}��a���7��������k�9R8�����8��>�Z���ۻ��\*�:�p6;q�c;��W;�f;��-:����������'��S��`�˼a����@�d�u�RǕ�����{��hȽx$ǽ�?��l)��ǔ�	����nd���X��Wa��|�pE���Z��B½w�ҽK�ڽ`�ؽC\̽ʞ��!����W���_�� 7�J��h����ݼc�ȼ�������N���bǼ�uּp�켄�����d?6�2�Y� ������f%��3н��������5��Kt�� ��~Խ����૽�������������o�˽�R������%��S�R������^ʽb����S��B҈�u�]�`�_2S��LK���G�~hG�T�I�bO��W��b�#�r�vN���ے��\��5���"�Խ���E���<�)��/l�����c������ཽoν�ĽS�ý`�̽�!޽�!��&*�c�������w����ؽ+	���٨�N���_���|�ļm�pd�I_���\��]�P<a��.h��Es��Ӂ��\���Ҝ�j����ǽ�ὃ����Z	�������E�����c��xYཚ�н��ɽ�ͽ�ٽ�)���������%���������+� �ٽ3n��䠬��ۛ��)�������>Px��Qt�<^s�Y7u�z�o;���������ٝ��  �  Uw?��������g'D�n�x��ݒ�aޡ���������Ғ�Ys{��eM�J%�c|
����&�[~/��[�("�������@��l ��(���AYy�X�D�������]�첼���@��(�;&�;�<�<H�<�j<f��;�`�;fk�:d�����6��m��� �w�4��k�i׎��뢽��������Ǝ�� ~��lP�G[+�|?�O��.(�N�K�y��X������ү�����������e�r�==��a	�����]�Z���Ի�ںh�:��N;j=z;�|m;�%0;�:�ĺ�@��|"��ֆ�U^̼0B���C��{�2N�����|Ľ��ͽ�r̽�5��d����z��5ă�ǩi� �]�	Pf�>������j����ƽpؽ�C��ݽ�	ѽ��������a����a���7��`�����^ڼm�ż����w!�������ļ�oӼgT����Q���5�	cZ����#l��\���ӽ?�꽱������ӧ��O�V'ؽ����?�������=蟽����������Ͻ2\�D/��rk������vI��:+�*�̽�B���/��-����`t��P_��Q�
�I��"F���E��}H�ۏM�DzU���`�-0q�qʃ��Ò��᥽a���A׽�򽅨�J��r�I�@������������-ѽ�ƽ��ŽK}ϽmT�����rl�2�������u�7��2���fڽ�s��u��I����懽�z��l��b���]�Ä[��6\��_�W�f���q��%��0����뜽0��HWɽ�j�����i�+������������k�tӽ�Z̽҂Ͻ�bܽ����z>�O��x��h�D��J*����۽}�½� ������𖎽�T���T~���v��r���q���s���x��k��7冽y`�������  �  �=��o��z�	�a>��Yq��B��纜������h���
��%s�%rF��8�q�oi��'�
�Iy)���S��Ԁ��ڔ�=�������#���B:��sr�Gm?�y��1���F�\��2»����{�l;]!�;���;lP<�<�<���;�f�;�t8:э�Z7� Q��ʨ���s0�ҳd�����H���j������F ��v���NCv���I��%�?V��<�&�"��oE�G]q�-ӎ�`���%}��0a���7��&���&�k��R8�9��t9����Z���ۻTr�[�:P�6;j�c;g/X;4�;	�/:hn���V���'�p7����˼/��Tq@�}�u�ƽ������r���_Ƚ�ǽ�8���#�������<kd���X��Ya���|�I���_��i½��ҽn�ڽ7�ؽ�e̽^�������a����_�7�������,ݼ��ȼ��� ��qO��7^Ǽ�kּ�u켻���u�!16��Y�B����v�����^�Ͻ�彔���t-���l������ӽ����ޫ�I�����A�������˽���X��}��N*�wX�J����⽃ʽ>���]���ڈ�� u�h�`��>S�WK�v�G��oG�5�I�
O��W���b�"�r�*O��Vܒ��\��b���;�Խ���J���<�,��2l�����c�������ཿoν�ĽT�ýa�̽�!޽�!��'*�c�������x����ؽ+	���٨�N���_���|�ļm�pd�I_���\��]�P<a��.h��Es��Ӂ��\���Ҝ�j����ǽ�ὃ����Z	�������E�����c��xYཚ�н��ɽ�ͽ�ٽ�)���������%���������+� �ٽ3n��䠬��ۛ��)�������>Px��Qt�<^s�Y7u�z�o;���������ٝ��  �  ?:�M���o���v�.��I\��n���U��7����������֞[���2����� ��?����X��E?�Oi����O#��M����Ր�#ۂ��3^��1�V��������\��ػ+��;�L�;���;�t�;S�;K��;�+�;��A; �t���=�y=��݅�r�$��5S���~�G���q���������������`�T7��;��U��R�Ve��=3�o�[��
���^���z��y���������d�Y�y�+�����U��[�^�	�����M�d^6���:�8;�.;C�:����G���ػ� 9��􍼮6̼� �]�7��g������o��Ta��SZ������+�������9����o�Q}U�K��2S��l�����$矽�ϴ��wĽ� ̽%%ʽ?m��魽!~�����;0Z���5�,��I��6�-Ӽ��Ǽ4ļUǼ!Iм��߼'|���
�����Y8���X�����^��^;���bŽ�ٽ�R��뽀�潈2ڽ1>Ƚ[��������昽�����ԝ����|����ؽ#������T������$�뽋�ؽ�ýT;���w����x�bLe���X�?�P��L�7L�4�N���S�+\��g���w�{1��p���w]���b����ν_/�������/y����#��T���-���@׽��ƽ���S���AŽ
ս�7齁���~���������4�N�������ѽ�x��������� ��m��t�r��ri�/�c��ha��#b��e�DBm�qnx�!���厽L��������ý%�ڽ���ZJ�\�
���B��MH�F�����|�׽8_ɽV
ý�Žjsѽ�}�Rv��#��[�����D�&�	��| �뽫-Խа���
��Wߜ��0������P���$7}�v�x�e�w�6�y�T�~��΃�Q4��(��� ���  �  =�A�3۟�������>��=^���r��oy��Gp�w1Y�̬8��6�o���¼�z���B̼aZ��� �$-E��Be�t�z��ɀ���x���b���B��2����}���i����&Vp��=	�	�/;�ȓ;Q�;���;�8�;w?L;�U:|,:��q�qvQ��V��7�����p�;���^���z�|Q��O�����|�*�a��>����߄��\�ܼ��ڼL���g���:�r9^��z��}��#��;�}�yOc���@�p����~x����p����V���#�rN�
��9,��9����� �0٫��5��0]��*����Ҽ�	��O.��U��&}����H���w���"��t��=A��o	u�ƝU��?�*i6�L�=���T���v��ڎ�=���#���$��8���ଽN垽g���dCw��*U��d7�
��r������%A�h�ټ1�Լ�ּ��QJ񼩘���T.'�$~>�Z�0k{��3��J�������w�ƽ�lѽZսoѽ�?ƽʶ�f����a���2��^�����v��İ��i=ƽN׽^����*}佦9ڽ�%˽޸��-0���+��F���QY�Y�n�b��2Z�C�U��wT��V�]v\��se�8�q�Q����]���0���l������iǽ]ڽ^�������� �L� ��n��ߤ콇$۽�_ɽ�亽̗����p���nnǽ��ؽ������M� ��� �A�����\ܽ��ɽX���$J��Oi����4��W�|�֨r��Fl���i��Lj�ån�a�v�����̈�V����֞�����X⾽'�ѽn��]b��<� �������������A۽܇ʽ�(��˪���2��OŽ#
ս�J罸x��F�����=��98 ���R(�c�ͽ���@����۟����z��s_������������z��能F������Ç���/���  �  m�c�����B-ּ6d��� ��D6�r"D��4G�mK>�!�*�|��c���-���̅��;��j��5l�������5�^H��O�#FK�ـ<�&���漍���i���iA���������
�}�PW�:g�;`d&;�!�:o�Ĺ,T�OA߻��3��р�����x�ݼ1[	�,?$���<�}P��AZ�Z�X���K��4�޼�����Yż�������B��"����L�1�i�I�D^X�' [��RR��?@��V(����f�5ٸ����U��f�n�̻ق�bf1�>�%��ze�ʣ��!&��TP�x��X\�������"�(���E���a��z��z��<���OÈ��M���$k�u�O�0U6�X4$�j��Pl$���7�F�T�9u�+X���l�����ة��V����5���d����m��BU��:?���+�;y����v��U�����n�eg��6� ����#���6�ߛK���b��|������ܙ��S������S��������8��T������&`���C��#ⅽ�b��� �[A�����bwʽ58Ͻ��ͽ�gǽ�E���S�����t���A���J݆���~�w�r��ai��Rc��8a��Wc��i���s�Iʀ�f舽#��vC��E���o���V��~�ν6۽���k齧�轍�὚)ֽ��ǽ�۸�.ܬ���������ļ��c9����Ž�qԽ\���罌f�A�-)ܽ Bн^ý��C���q,�������T��#:������|dy�k�u���v��|�󳂽����ᐽٙ�M�������<��;�ɽ�׽���B뽹��,�����V׽��ȽC������8���^���˶�W�ý�ӽ8k�eb����������սǵȽ���9���Z���b�����N��~��z�����^���ъ��6���1��2t��$䨽�  �  @y������Dּ���|��h��}��U�J��� ����ʼ����f���1���#�λ?��v���~���޼���߈����o� �� �G�����A!�.�ͼ�k�����Be_�T�Cʻ��^�v|꺝Fκ�7��̭�����{Q�S芼,}��h�̼
W켾z������ �nD)�
,��a'�������6߼田��Њ��mj�kh����	꫼�	ڼ��B���&�Q,�)a*�d"�)��̪�8B��h�ּ���M͚��+y�l@�&a�4��v�ջް��%$��a�镼%��.K缌T�~�,�eN=��$M�DRZ���b��e�b_��R�]?�F�)�B��{.�٪�G�	����`k1�eL��of�@�{� ���g��qS��uj����y�ۇl���^���P���B�?04���%�B��L0�"R�i����{F��)�4�;�fO�Pb�b�t��&������(�������%����ѣ�9{��(:��h��B8������:�r���g�	�f�+�p�3����P���䛽�R���ֱ��h��A渽������Ԭ�������������Ғ������Y����~��zv�k�r��ut���{��-��d:��i8��sa�� =�����������q����ƽ}�̽�ѽ5aҽ��Ͻ�Mɽ�`�������§�V<���Ƙ�Xt��T���n������꽽yȽ�Ͻ�
ҽ�1ѽSMͽ�lǽ�����'��ܛ���٩�]С����"����ˊ��Ʌ��`���烽vT���8��)Д�&=��Vϥ��*��I?��t ����Ž
�̽�ҽ+lֽ��ֽ�@ӽV�˽�a��맵�ƻ��>����4��Z�������4��oQ��oʽ�ӽn�ٽ�`۽��ٽ�$ս�Ͻ�Ƚr����c������2���Ұ��?%���瓽)я�z���������i'���3���ѫ��j���  �  I�ҼR.伜�����i������~�u�ټ1
¼ r��p�{�*12�����ї�Is���%���	�voP�����ᵼ<7ּ����(
��6�n[��W�v�������jԼ)����T��W�S�=��x��ݻ%���>��e������]�ϼ�p��t�%�	�����?�������`�����6޼Ϥ��	t����a�n�'�!���#���"�w�Z�S������ �ڼUZ��<�����&(�-&�TJ�I�8a����k�޼1G��K���a�x�M��j=���N�Y(�����ˣҼgm ��t���&�tA3���;�C�@�Y�C��5D�E7B���<�0�3���&�6���2�a!２�ۼ�yּ2p�ߪ������&���<�tdP�|�_�8�j��r�0v��w��w��t��n��kd�I�V�� F��f5�V8'�pe�����#�ִ1�<6E��F[��p��ၽm6��PX�������g������Ǔ� ��=����j��5G���t���c��_V���N�Z�N���V�&Gf�&�z��t��#4��Uh���}���n��蘫��q���E��S��	����A��5��4���)��?v���k��S�������y��iF��=4��̥�e���Lɷ�󶽽%����ý�ZĽ-Ľ"�½����[�������>Ǫ�����ٗ�d����X�����ˏ��ɖ��ٟ�o����j��v���tϾ�/½��ýXTĽ��ýY½�9���&��'���>���Ơ�.����S�����/���`/��tӚ�VJ�����(���q���ý�!ƽ�ǽUȽD�ǽ�7ƽ��½j����G���i�����i���o����WV�����4����W��.$��;Ͻ�]�Ľ�NɽD2̽@�ͽC ν��ͽ~�˽sȽ}½⺽�ᱽf����|�������i���堽"f��:��b��TŽ�  �  �t����-[�2��>���8ؼ����&��qV|��F<�����+��l1��N�=:���:0/�8�$�w۷�#X�ASb�`O���T��fZԼ��󼖻�!��h���
$�� ����e����ټ+��#���X���P�	s�.`���]ʼ2�����g"���)��)�K�"�4���
�������ؼ*���ꂙ�(�p�3�/�ن�
���xD�yF?������?�3)��i����h��S�ռ���-�������"�q�*�"�,�n{'�+l��T���⼄a�����Eˎ���4/��j�伴���I)�F@�v�P�+8X�� X�ȦQ�L\G��;��-�aP ��k�$%����_Ѽ�
s���^���K���˼�g����%��.�QFA��S��8d���t������Ǉ��e��+�������d����Wm���W���D�'8��(5��<�wYN��f��ˀ��x��Bw��T�������h���{ѓ��B���s�����p�Mob�9ET���G��>��/9��:�KA�GjM���]���p�jK��T����.�����˩��mݮ�n7���绽3뾽ub���������&��'󝽇�������e���ޖ����������MŽIoͽѽ�ѽ;.ν��Ƚ���-F������K���Qi��i��������[�����(����p��/�����h����ј�R7��[q���e��M%��c�����ǽU�ͽ$�ѽ��ҽ�Ͻ��Ƚ�����̲��~���Ğ�3X��X"�����᪽9ݶ�#�½U�̽�8ӽ4�ս�oԽOJн^Sʽ�pý�-��@����
��N������H��x���+5���[���v���j������{����#����������7��Ž��̽
�ӽ�hٽ`�ܽlܽ;ؽ<н\~Ž�ǹ�z;���姽�D���짽�f��;K���ƽ)$ҽ۽�  �  �*C��@�4v3����&��N�ּ���;�o�+v�[����b���:\�m;y��;8ݫ;��;�H*;��0��+q�������L��ґ��y¼Fc��'��x0��E�8Q��9R��CG�"�1�����}��������e�������e�ݼ�����)�MuC�b:T��jY���R�	`B�c+��V��,񼼦����R�g
�&H��&����8�:`�:|\9h���e������J�.��>㷼��輗��"!)��
A�!�R�O�[���X���J�]�3���2���P:Ӽ(����˼���:���5�ޝV��Jq�Ѐ��؂��~�%-m� �V�$�=�(�%����P����ּ����̣�n_�������ꊼ���g�������4�/��UZ��1.�fRG�S�b���~���nؘ���Z⣽$񠽹���	,���|���c��iS���N�D�W���l�hX��˕�mꤽy%��Hȵ��L��d[��Nv���k���،��‽GLl� �Y���I��p<�b�1���*��(�{�)��/�7:��"H��Y�}il� ꀽ����ƙ��ç�a����ý��νa�ս, ׽�ҽ�lɽ�׼�*���¤�x��������������\��%#н�ݽ�d�2H齅&潎�ݽ�{ҽ�^Ž ��g����_���g��"������	��"�v��@r���q��v��d~� $��%������A垽s���=]��פýK�нv�ܽ��� 꽈�轵�b�Խ�]ƽ�"������n��"a���ï��$���˽��ٽM]彰��j�콚��E1޽Sҽ�Ž�A��D}�����YΘ�'ʐ�� �����D������׀��냽�������[×� ����q��a4���&Ľ~�ѽ�߽kc��|���!#����ڽ�X̽����.����@��B����徽>�̽�۽C������  �  �Nu��1o���Z�xq<�%u���,2��fL��һ�ͺ��;!�;n��;��<�<�.�;h��;�Jl;^��9����;��Q��~�ür#��R,���P�qgn��p��sT��0�x���_��!>����n����Լ�hμ_�_�1�H4U���s�/\��^b���\���f��E��� �	���򬴼w�v�	G�����y����a�:�fW;�b�;�;n�`;[M�:�2T��ы����n�j��ǭ���;���B��]d���~��:�������/{��y_�"�=�o#�������X��'���5�I�\�r������*噽�Ś�����U ���m��pI�N)'�*��bo߼'η��晼*���+�m���a�- e�̐v��;��7R���i��¹�N�	��$�/E�`�i��X�����A/��V����伽v���6��mB���\�����:�m��yg�	�q��<���ږ��a���.��Oɽ�ν�o̽��½M���Т��ؐ��$���yc��	L���9�KZ,�E�"�-k�x������7#��[,��9�]=I�X,]��hu��;���.��1������.�ӽ�e�T���l�޵�5rཕѽ~���yF��q��b&�� �������>$ӽp��`���	���[� �]s���G�5�߽�ͽ�~��Y������S��}���(A|��$q�%�i�@�e���e���h���o��sz��d��q���E�������1��©ʽ��ݽȵ������O��� ��`�����jٽ�0Ƚj˺��򳽈���꽽��̽��޽�_�a��K��XX�'������Foݽ��ʽ�	���0��{ݛ�e��w���5��m1{��u�2�s��#u�N>z�<|�����=������v���u��e�ǽ<�ڽb_�{���������"������^]޽�,ν&�½i�����½Z�ͽ�4޽i�𽢜 �����  �  ����V���;�4QY���,��r������kC�����D$:���; l�;��< �$<P'<Ջ<�<9^�;z�.;B���%�����ͩμ�����B��Lo�@��"���kR��Pԑ�8r��F+`�9a7�����X��������
���(��P�y3z�����A��.������r����_�:�1�{�����m�f�k��S��|�:��w;���;���;X��;|��;�q�;�8�:0����޻�*Y�K���[���o�,�>&[�¹������Ѽ���y���a��Dc����]��7��}��Ea�J�*��P��}��ܔ��1���¯�+���]
���Ж����C�W��m-�y_��Լ!ꦼ�s��1b��qI�\Y@���D�9V�0�s����������Ӽ����J"�kH�p�t�/������ ���̽��ҽ��Ͻ��Ľ�+������[ƍ�������{�Q���͗�������޻��н��޽�佩Ὥ
ս��½묽D�������6a�I~E���0��"�c�����њ������"�#��/���?��T�"�o��ӈ�8��%���S̽g!�.D��/Y�}<�ɔ �����%⽺5Ͻ;h��0��Ϡ�����<4ν��⽽x���>�9�
����+>��� �v��ʸս����n��8���Q���݀��xr�4�g�]a���]� {]�[`�D�f�x�p�1G�������z��� =����ҽH��N��������|#�u������H�սAƽ�a������u�ɽ��ڽU�ｩ��M�	����I����ߙ��3齹ҽ
:��( ���2��5댽�у���z�*r��,m�ȅk���l��xq��y�MÂ��-��艖��O��x���ͽ=K�8Z�����^��Ʒ�U�[
���"���ڽ�ͽɽ�lͽ�Fڽ)�����
�|U��  �  *��������U�� n�X<�)��^x��ҧE�`	�� E�:dN�;-E<�=)<="7<�%9<@�/<�<b��;J~;~{q����҃��(ڼ���G%S����,���$��G\���^��`����w��J�[�$����G�	�����p:�g�e�l��������/����������@t����r�El?�3��"p���d���ڻf� �#;�~�;���;��;:��;E��;���;&�:;i�J��bû�_U�E��AZ���9��m��q��6�������d��Q�������s�c�I��!*�ڑ�%*!�-r:�62c�����tС�����M���̔��X��p������4Zc�֫3��$
��YѼ�@���"y�6PM��5���-��>3��-D���`�]���^	��˼�4 ���"���L��}�/s�������ʽ��ڽ��(�޽iAҽ�;��%��� 9�����6ф�Ƿ���֙�t�����ǽd�ݽ�1�hx�lZ���gͽ��������}n��n�a��C�I�,�[��pu����C)��v�c�����E�*�$�:�/Q�� n�䒉������x��ycԽe�h��Ť���
�A��� �����ؽ�{ǽ�S��Ŗ��)�Ž�׽����|��F�UE��O�61�����9��sܽ��½�	��2Ә�a����}�SOm���b�?T\��7Y�Y Y�e�[�d�a�ˀk���z�m������,Z����qHٽ�K�ʇ�(�� ��oZ�;�K8��S����޽�ͽ|QŽ+�ƽ-�ѽA:�!����_����]�U�������ģ���׽m_���詽i����*\��x�u��$m�K�h�*g��dh��l�)bt��3������s/��e������	�ѽ��뽻��@��p���6��h����-����4^��$ս��Ͻb�Խ���x����wo�����  �  8-���U�˼秗�O�4�V]�c	t;h�<��l<l��<�ե<�<���<*j�<�9�<	�<���<���<ީ�<�T�<�2A<��;�S�������������������������@ǰ� �u����\ûu����\ �|�Q��a����ռ++�~V�����P���漾O��u?^�t`»"�t:���;�54<��g<�^�<+m�<$��<eJ�<�K�<���<ˮ�<i��<�j<U�7<k��;/+�:
t����V�����F漏�	�eH�ש��4�-�
t��M���H�H�(�;��S~�����+����H/�a�<��R=�D�1��,��Y ���ļ�!��z�2�֦Ȼ�/�P��,G:1O�: u�:�J:�I����к�lW�x0���Z���Q��|��h=ʼrN���%��F�-�c��Px�gွ��~�Uzp��/Z�1�@�'�)�-}�+F�?���U2���M��dl��	�������1��#��^���}w��Z���;����\��q�K�Լ`ż����Ð��V߽�SüIk˼��ּ���ƺ���R����S5���Q��[r��<��!}�����P���i��
��ߨ�vf��=�����wQ���W��rn��V����Ǡ�#W��l����ý[}Ľ@���a;���%��R�����-�r�U[��(I��<�73�b-��#*��(���(���)���,�n2��;�s�G�;iY�1�p�rM��.���.��/ݴ���G6ƽ�"ƽ����%���ǧ�b���=]��q!����k쒽	q��$J��ƹ���ĽpYɽ�iȽ�p��@���,צ�c��4ꇽxu�,A`��iP��_E��2>�n�9���7�ə7�.�8�P�:��?��F��TP��_�p�r��������J���T��;Bý�ͽ[_ѽZϽ�ǽм���@���塽 ;�����(��M䡽��������.oɽ\ҽ�  �  C���6⼏���o���z'��}9�>s�;e� <I�k<|C�<��<�+�<3�<6��<�߹<�<���<���<;��<4�<�q@<C��;���9�O�Qq�O������r������;��n�ؼ?0��P�e����W��4B��O@�9C��{���a˼	���
�cF�o�7�ܼZ��/ZR�E���*�:խ�;fZ2<Q�d<Z��<���<��<;�<��<�/�<���<;)�<��f<�5<���;��:A���R<K�7���Iܼq�����g�N����w~���Ձ�cB<�W��w/��Sq�����B��ӳ��)�zC6��37�%,��o��Y��t����8����0�� ʻ�9�}�1�'e:�/�:��m:R:�9���K����d�w彻��vS�䓼5�Ǽ�%�/�"�s�B�`V^��Br�	g{���x���j�'U�އ<�~M&��h��c����w�.���I�U~g�|;��ꊽ�������f�� s���V��9����H��ּ�#Ǽ`Y��$���<����ļ��̼�&ؼ �缡L�������l�4�cmP���o��f��7���1��iޭ��尽���u������2��Za����^��m҅����c�������䖸��뿽*X��h�����������ԕ������r�Y>[���I���<���3�/?.�#�*�g)��W)���*���-��S3��;��:H�fY���o��n�������0��d[���6��MýB�½^
����O���W����������㊊�MA��_w���墳�������z0ƽQŽ!����<��5���O���)����t��``��Q�6F�J?���:�C�8�G8��69��;�g@��F�sQ��j_��r����� ������r(��*����ʽ7ν�>̽��Ľ6�� �����&���韔�c����!�� w���.����ƽEϽ�  �  ��ɼ�N��렢��?l����q���$�;�w"<�<f<�e�<�Y�<\x�<�ݱ<fK�<�X�<s?�<��<���<(S�<w<B<<���;�đ:����R�I�����X�Ƽ��ۜ��ڼ�U��1���s�7��˻�M��-�����N��mgx�sŭ�RT׼����L��X伷#�������X2�4=�����:�m�;� +<MZ<׋{<��<'�<�N�<�W�<Z6�<�o�<Ī|<��[<�.<���;x�:&U��0�,�J卼��������-��E����F���ļz	��.Y��B�)b���o�;AL�#����6μ�o�%.�e�$��&��~�fF
�R/��챼�ڀ�0�,�8�ѻ
�]�@���l�;����9xz�9T�9�4���v��^���#Ի̧��X��V����¼�������}6��wO�zba��i�p�f�dZ���F�Rb0�&���P-�����$��
>� �Y��r��H��"D�������{�R�f���M�G�3������z���ڼ\�̼��ļ�8¼o�ü%�ȼOѼ�0ݼ��� �������g�3��L��%i��l������^��w3���󧽆Z��y.�����-j�������v�Hw��?���b��/2��
L���B��_��:����h�����is���ґ�rG��Ip�z�[��jK��p?��6�i1��i-���+� �+�.-��0��:6���>�)J��Y�8n��5��uѐ�ƻ��g�����O���!���������,��S��j&��y��oM�����_ٖ��?��UB��/���M��裼����뗬��ߟ�iF���D���s�F?a��)S���H���A�>�=��";�Ƌ:�j�;��6>���B�B�I��S���`�-�r�0R��C��FO��-��7��Z���YŽt|ýے���
��������`D���x���C��!��…��!��猾�Ďƽ�  �  ����>���ao���'�S��s��9��;��<,W<>�<*�<�<�<�Q�<���<��<���<��<�0�<Oc<e/<���;P�:DSa������l��#��b���V���e���ʊ���F�MZ�W0�:�����9&Ⱥp��Q�,�U����,��N�V��������ڗ�[a�`��,JC�C��:3��;��<=|D<�<e<tM}<N��<}�<���<�̆<e~<af< F<]�<�y�;_
;��4�
��<`�xo���3���_ʼd�ɼ��������d�;���Ļ�q��ι�5��j�?���5�׼o���[�
�g
�"�a���ɼ�ʠ���r��{-�\��[4��~�3�ɺn�j��;R�������b9h���.����/�
�g�v��mM��!��[���%��K:�� I�R�O��!M� AB��g1��;����$��w���H��5��p,�t�D�U�Z��+k���r�H�p�J�f���U�d�A�z�,����67	����MQ�4�׼��ϼ��˼�r̼u?Ѽ�ڼ����z�������#�!�K�3�P.I���`��ey�Bg�� (��`���ݚ�ș��x���ች��q]r���i���j���t��f�������?����������(y��𬗽����󊁽|�n�̰]�8�O�7�D��p<�@6�'2��0�00�c�1�p�5�"�;���C�a�N�`\��_m�~���1䋽�?������cl��.���h#��.@��Ο�8s��:=��HA��`~����}d��3q���E���ţ�O�H��h
���c���>�����鍽_O��M�s��Jd���W�?�N�z|G�'�B�5�?���>���?��C�?+H�K_O���X���d�� t��P����͆��Pޤ�����:����g���������<]�����^������ =������������������;���;����  �  �5���/�Hf�����|��[��:6�;|�<
7<��^<�h�<FT�<�}�<x*�<^�<d��<#��<+E�<Y�f<m�><j�<�b�;�q;������»����R�#�o��Ks�})Z�w6(�Nͻ�A��0�:�Dt;��;Ca;�Z�Ab��P���iY������\���z�V�X��"���ǻ�L��a�:�}�;�i�;��<wh@<n�[<�o<0y<ty<��o<$�\<$�A<* <��;��;@��:�F��QȻ��$��^��w�������H���:}���H�/
��򛻅P�ZP�����b1�����(q�SM���ļ`mڼ���|ڼ8Lȼ2��f��Eo�ޜ=����߻�f��{u��S<�,}(�{,=��{�bn���9��"R$�íS�;����Š��|��L���4��g�5#���-��1�%+/���%�-�ݫ���������V�mb������A,��R?���M�2UU��U�Q\O��HD�֊6�b(��z�Xr��N�L����꼝��ۼ�5ڼ�x޼���Z���I��6�Wz��)�x�7�dyH��2Z��Ql��h}��ǅ�6e��4̋�����r�����{���l�|�`��tZ�o�[��hd�l�s��q��d7��ቕ����z����M��S���<ɏ���������?q�F�c��[X�zFN���E�\�>�x�9��7��6�3K9�8>�+�D��sM� wW��c�~Cp��2��������# ��j���������Mř������	��כ��kv�zao���p���y�Zo���s��GC��=E���G��9���\ڞ��Q��)���c��=˂�T�w�U�k��a�^X�otP�>�J�JG���E�1G�o�J���P��X��5b�O)m�B�y�����ދ�2���J���:��d���e�������si������_$���D�������͂�;ꄽv������x5������(ت��  �  ^j��������t�׋�H��H��:��e;F
�;n��;p$<
�H<~j<NT�<�R�<+Ӌ<T{�<�u<ΓT<Pj-<=<��;��L;�VB:iҺ}�|�	���I����$��H�ǻe���{��J;�;D��;%d <��;x.�;w�:W�F��4˻O�
�:�A��j��J�仏m���>�c?����:�w;�`�;{�	<cE+<!�D<�ZR<[�R<��E<-<޵<X�;��y;*��:5\S���G��}�������'+��1��&��	�J˽�s�6�7L�6�T;9+;��:C)d�Y�����7�X���������i���.��up���Μ�L�������f���H���*�TC�m�C���祻⊪��/˻�1��+��[�����:���X���tμĜ�������d�����<���S�sh	����� �伯)м�Oü���J�ͼ������1�cc#��Q0���8���;�P�:�*6�Z�/���(�9!�����<���
��I�����S������dm��P�������)��6�[�A�3�M���X�${c�y<m�Y�t�b�y��y�ͻu��qm�\�b�r�W���N�MbJ��K�umS�4`��o��������"���Ď���������ω������W��4�y�Gp�G�f���\��AS��J�]ED���@��@���C���I��dR�� \���e�ƫo�Q+y�'C��>ۅ��2��䍽<Z������D���3��x;��Ŝ|��Ko��e���_�-�`�b9h��0t�fS��C���?���׀��/���_�������t��dg��l%���π���x�n�o�{ef�u�]��=V�^>Q�^WO�[�P���U��9]���f�t�p��<{�ͨ������(p���)����������%��ʘ�S&���ݍ����׀��"y��4v�Χy��o�����ρ��˄�������  �  	;tI:��X�0���Ҥ$�֧����8w�:	o7;[��;���;=^'<�"K<F�a<��f<��X<�A:<��<%�;��F;�':ĵ��.��L��(d��i���Y��a/��]ĺD5�9�u+;cq�;�� <1#<~7<K�9<#�)<@	<i��;�):;��8�v���x��ȟ�%���I=���2���{��`��� �R�뽥�\c�:���;�m�;Ş<� <�y!<6�<���;�I�;2�:�=���Y��Ɯ��񺻽˻`ѻ��λ�ûI��F����t��u}8�;b�;�ͻ;E>�;F�;i7D;���Sl��|S.���[��I~�?Q���u��艘���N��Gӕ�*Ì��+~��\��|8�,�J����}`�X;��Ql�Oo���Ʈ�A
ȼNܼ�'�E;�������9��h' ��b��E����H�X�߼��ͼ����f���0���������2�¼MXܼ5����P
�����# ��'��+��.��D0�L�0�G`/�X*,��&���='��q�ޟ��>�[a�.V
�ʅ���!�*�/���=�{�I��"S���Y���^��a�Ćc��3d��Vc��{`��\[��0T��K���C���=�/g;�|>=���C��M�]YZ���g��t�[>~��ڂ�5J��I���=��'&��QX��ٟ��3��H{���p�ze���Z��Q�M���L�#LQ���Y��`d���o�u�z�����ް������������Dꇽ	��H��p\��&n|��&r��g��\�0(U��fQ�WR�'�W�@a��pl��Ex�0~���ą�cψ�����nы�2?��:���7��b��"^��}"����y��o��Ye��g^�*�[�5t]���c���m�VWy�h����އ�.����䎽����O�����%ᑽ�琽�쎽����nZ��!��Ȅy��0p���i���g�+�j�ĭq�q�{��냽�Ή�ꎽ�  �  ���;:�;8��:Y���+���R`�����xk��̗���;bݮ;�<�%<�-<�<�Q�;�t;]��8��S������h��'ﻞ�ջ�[��QP�;M���|:�+K;M��;���;4� <ްA<�2[<z�i<��j<5�^<�F<B$<'L�;RϨ;�^1;�t�9Ȥ�����)ӻ�r�&���%� ��.��󱝻����J�:�c�;��;���;�_�;�;�}��z���� t��S+�j�&��2��T��M��=yW��ߡ�H�P:�9;e�;���;Sz<h�<'�<�5<��;�	v;�-G:��!��)��#����A�.q��<���-��ӵ������3Ƽ�4�����Q,������� b�0�E��>�R��:}�>��I��x�C�������
����3� �������Լ�żKh���b�� ���(�������͍�O�ʓ���X��KӼ(Y��|�XJ�ܢ�n�$�U/��8��6@�{�D�|E�_�@�"\8��-�ZJ!�nw� ��a��D���%���5�� G��W��bc�u�j��m��(l��g���a��[��7T�RpM�,�F�߶?��9�pi3��/��.���0��*6��[>�	�H�p�S��O_�)Hj���t���~�A&��!���Cy��2�������������Ʉ�=�{�A�m��2b���[�xX[��Da��8l��z��,���J���w��$D���Ǐ��y�������څ�~~��>z��q��g��R^�l6U�^ZM�#�G�;E�f�E�`J�fQ��Z��#d�cn�gx�q���慽K����������t���nY���\���	�������Pw�W�m���i��Fl��t�Y���U���,��� ����ƙ�ј��:��z���Ȕ���X���	��/���8)z���p�Wph�*ta���\��[�Q�]�W.c�%k�y�t��$�`����  �  ��<��;���:>O�T�˻���1=���E�'�1�n��|;��(uI8�/v;��;+��;���;�G;����̻��'��T��Gg�BW]���:��6��V��f�I�Eg7;� �;!p<͘6<KX<�0s<�J�<�k�<��<�߃<��t<R;Y<�6<��<|�;�{0;�s�������/�L�I0{���������o�r��<�~(ﻚaH��2�9_�;�$;l�.:�S2�Y#�68���q�F9������]���\��`#�ʻ����$y:Pe};�h�;��<!<uN2<��9<ߕ6<nO(<N<W�;�5�;D��:���Z�»��"��\i��p��P[����ܼtP������2��X5��Ӽ�o���痼���U|�嗈�#K��� Ǽ-p�|��?7�?$��%�j] �����{����oDؼ~{��;n�����%����T��%vs��o�+v�vw��\Ő�Sq�����"�ϼ.�������[�$�P�6���G�r�U��5_�1_b�{�^��|T�R;F�]�6�Z�)���!�Ew!��Z)�uT8���K�l�`�40s��X��J����Y��A����t�\g�EIY�1~L��nA��F8�M�0�o+�<�&���$���$�'��+�h�2�7;��UE���P��]��j��?z�PL����������.�������
O��gX��al���ŉ�^��.�s�uWk���j�Ipr��)��߈�i����昽QO��*9������(f���M���q��QO���p��Ad�]FY���O�X�G�łA�;N=�U|;��+<��X?��D��]L�z�U��`�5:l��z��Ƅ�(���*���S���s��+����>��w������|��8X����~�n^y��3|�{O��CE��Lp�����A����>���-��dԣ�����ݷ������������j�u�|k� �b�ʈ[�� V�7�R�"R���S�X�/j^�f�f�\sp��{��  �  ��*<$C�;���9"9���.�P"z�5��Bt��S3����r�=�&�ui���,�t�;�Q;l��:ƶ���\�K��y��NE���î�VФ�w���$lJ�ȷ���⺎�P;(#�;��0<�9\<�=}<���<���<l�<�_�<�|�<���<�F}<��\<��2<zK�;�kj;�|���Kڻ��H�]Ď��:���hü��ļ�ѳ�F���WU�h�d�q�����U���]�����[IN�� ��0���dƼ��Ǽ���~䗼��^�i�~�A��#�:�e�;��	<��,<DND<�Q<��U<�P<
�B<��+<��<cJ�;ӢS;����8��3Z�4kw�����޼�����ry�?���d��y�m� m��B���כ����E�ļ����<�)'�B�8�S�A��A�|8���(����	����Xؼ�L��4��U���4Mp�ݔ]�W T�M�S��k[�Ek�'���sj���J��3m����ڼ����I��L*�$�B���Y��m�l{�����K|��Bp�y�^���K�*;��1�a0��8��TJ�]Aa���y�󐇽����?�����M��揂� ,q��]���J��;���/�L'�M�!�l!�����z����=$�ZC*�R2�n�;�,�G�J�U�&Ag���{�����s�����Z�����EM�������֟��{��?銽
;��vz��y�+���b≽�b��8ꞽo��%S��˴�������Π�!������ʣ��'�m�Yv]�ukP�>TF���>�cF9���5���4�|65�4�7�:j<�!!C��L���W��f���w��h���͑�p7���Y��Qɮ�M��9<���ū�{���#���z����[���#���Ʌ�������n���}ݪ������3���>������n��t�����������6�|�Cn�nGb��RY�O�R�62N�k�K��HK�{�L��/P���U�IE]�v)g�O�s��  �  ��.<:��;s������Lt�gk����Ǽ\kҼ\Ǽ˨�lz����T��� J�H�9buغ�0���y=����$뼼��ټ�q�Lռ�_���慼�� ��TU�4"4;5��;�A<�jq<�͉<�K�<�8�<�M�<��<���<�ϔ<���<��r<@�E<o�<�h;��6*� ���.���}�ݼx�������R�_���:���D�k���E�������޻�;����Z2������~������Ǣ�ﾼߌ���,�>L����:!=�;(e<V�A<�Y<T�e<9�g<
a<�&S<x�=<M� <w��;ْ;Z3:	����}!������¼�����R��-� `7��6�"�+��p�)M���ܼ�9���������� ��L	�J�$��X>��Q�I�[�JZ��nN�Mw:�H�!�(���޼ⴼ-���5y��Z��H��|@��A���J���Y���o������r��B����Ӽy���w �?�1��O��Qk�����䉽T�������	�s��?]���I�z�=��O<�`�E��uY��Ls�lg������ڛ�]������b��v���lJ|��#c�siL��9���+���!����������i��������%��y,�Y&6���B���R��Jg����&p��}���}���������gN��g���+>���]��Q;���H�������D��Ts������D+��#⳽0T���o��@0����������I�������Ln�k�Z���K�f�@��+9�U4��?1��70�R�0��3�(7�6�=���F�%KS��d��Ny�ND���(���������ֳ��5+��/��� ���譽��v�������c��~;��mP��:���ͪ�ʒ���C���6ý��������e���u��镽�'���E|�#�j�4E]��S��AM��5I��4G���F�R>H�vAK�FP�G�W�lb��p��  �  ��,<���;KU7���+� ���Ƽ��� ���9�$�ȼ����RI�A�ػ�U=�
��7Vz�f����n�n���8�ݼ�����{��;�Ѽy|��#1C����Q�;��;'�G<��{<3��<2�<�U�<`�<㣣<���<<�<�u�<��}<� N<��<�T;�T���-��X����ϼd����g��.�;�g༝�����p�Z����һ�2λl(�"yg������ܼ�S�J�	��\��U�ڼ${��S�J�&,����:�"�;�"<�L< �d<��o<��p<p�i<�[<5_G<�A+<|h<���;8�:����K*�Н��LeӼQ�
��'�U�=�� I���H�Z�<�R0(�����&4ѼPż�ѼQ��;���12��N���b�@Vm�}`k���]�7G��Y+����*��\���鑼p���N�U�<��6��8���A�_�P�e�e�
j���피���'ѼZ����/���7��\X�9�w��C��j�������������ڿ����h�ɳS�vF��zD�x�N��c�uc�����t������l˧��줽>����z���`��s^h�
�N���9���)�aI�������4=���� )�{���H"�\�)�V3��@��R�S�h�Ł�j��������2��¯��yb��^.½t����벽����eʘ������ʇ�1w��J�������������P��2½`0½�?���f���Y����������o��=Z��I�\ >��D6�ea1���.��-�*~.�e0�c\4��:�wD�֍Q���c�cf{�����P@���֪������½[�ǽ��ƽ�E���@��q5��Λ�����e���손�A/��������fw��N�ǽu̽8Fʽ��½W̶�EI������Ί��}�=ti�o�Z��P��aJ�ɎF��D�X�D���E���H��iM��T��_�n�n��  �  �~+<%ׅ;��[�ڡ9�"��;�Ѽ\���,P��m��Լ Ң���Y� ���>n�y�)� !���;����E'���7���>	��7�-ܼg���O��b���@�:V��;dI< �~<v[�<_��<<�<�W�<,��<7�<{�<�A�<h��<�lP<BD<��J;� m��$8���sBټ{����p�C	
����;��[��K�'���)���1!�G�v��8���6缞M	��Q��,�h�����^��4V�Vٷ���u:*�;��$<R1O<xh<j"s<S�s<l<W>^<�EJ<��.<��<�x�;]h�:g=���
.��z�� ټ���!�,��C��nO�<�N��vB�!`-��D�NH��-�׼"˼R�׼�������h7���S��i�Ȧs�f�q�jTc�0�K�v�.�{x�y��KJ�����مm���K��.9���2�v�5�9,?�$�M�0�b��]�;��ܘ���м����Hl�~:�H�[��U|������r��**��[�������q2���m�:&W��vI��XG���Q�/"g��Ӂ����kw���������姽FB��������Igj�u�O���9���)�I��� �J��pp�����v� <��l!�6�(��}2���?�vR��#i�����H��ǌ������p����|Ľ�UŽ���&����Q��Ͼ�����MF��p�������j���⦽qi��L���XŽ�OŽw#���᳽�O��h������p��7Z��JI��P=��^5�[�0�(.��A-�/�-��/��}3���9��OC�NQ�`d��Q|���� Ŝ��묽L��*�Ž�$˽� ʽ�2ý�׷�Xi��(���Q0�����	���噽��L��A����ʽhEϽ.Wͽ��Žv�����K��dz���x}�!<i�QZ�!P��|I���E�JD���C�+E���G�F�L��S�.�^��n��  �  ��,<���;KU7���+� ���Ƽ��� ���9�$�ȼ����RI�A�ػ�U=�
��7Vz�f����n�n���8�ݼ�����{��;�Ѽy|��#1C����Q�;��;'�G<��{<3��<2�<�U�<`�<㣣<���<<�<�u�<��}<� N<��<�T;�T���-��X����ϼf����g��.�=�m༥�����p�t��1�һ�2λ�(�lyg����Ʉܼ�S�|�I������ڼ|��m�J�#0����:"�;�"<�L<��d<"�o<��p<��i<�[<{yG<`a+<*�<��;/:�����*��~��@EӼ1w
�+�'��=�cI��H��<��&(�������U.Ѽ�Nż@�Ѽ?��w��:2�9N��
c��cm�fok���]�:GG�j+�j��H�sx��g���6p��O��<�+(6���8���A�L�P���e�I]���ܔ��خ�lѼ����� ���7�ALX���w�s;��Ub������!���k닽I�����h�+�S��sF��zD��N���c��j�R���A��������ҧ�������������/i��:oh��N���9�)�)��U�]�����E���@.��� L"�χ)��W3�T�@��R�؅h�<Ł����������2��̯���b��d.½y����벽����gʘ������ʇ�2w��J�������������P��2½`0½�?���f���Y����������o��=Z��I�\ >��D6�ea1���.��-�*~.�e0�c\4��:�wD�֍Q���c�cf{�����P@���֪������½[�ǽ��ƽ�E���@��q5��Λ�����e���손�A/��������fw��N�ǽu̽8Fʽ��½W̶�EI������Ί��}�=ti�o�Z��P��aJ�ɎF��D�X�D���E���H��iM��T��_�n�n��  �  ��.<:��;s������Lt�gk����Ǽ\kҼ\Ǽ˨�lz����T��� J�G�9buغ�0���y=����$뼼��ټ�q�Lռ�_���慼�� ��TU�4"4;5��;�A<�jq<�͉<�K�<�8�<�M�<��<���<�ϔ<���<��r<?�E<m�<�h; ��9*����1�����ݼ}�������Z�_���:���D����[F��Y����޻��;�����2���伦��������弓�������,��S��֪�:b;�;(g<*�A<��Y<֡e<��g<�1a<VOS<]&><� <�n�;���;�Q9:𸄻�!��C����¼i���4�{�,��D7�#�6�X�+�n^��>���ܼ�.������(���W��V	���$��l>���Q�ľ[��fZ��N�w�:���!������޼����\��W�y��_Z��8H��@���A�=�J���Y���o�2؆�&R���]���cӼ���D�U�1���N��1k�k����Չ�y��)㊽�냽m�s�T2]���I�!�=�P<�Q�E�Y��Zs��p��>����盽��������r������k|�CDc�o�L��9��+���!�d������������������%��~,��)6� �B���R��Kg�;��Wp��0}��~���������tN��q���3>���]��U;���H�������D��Vs������E+��#⳽1T���o��A0����������I�������Ln�k�Z���K�f�@��+9�U4��?1��70�R�0��3�(7�6�=���F�%KS��d��Ny�ND���(���������ֳ��5+��/��� ���譽��v�������c��~;��mP��:���ͪ�ʒ���C���6ý��������e���u��镽�'���E|�#�j�4E]��S��AM��5I��4G���F�R>H�vAK�FP�G�W�lb��p��  �  ��*<$C�;���9"9���.�P"z�5��Bt��S3����r�=�&�ui���,�t�;�Q;l��:ƶ���\�K��y��NE���î�VФ�w���$lJ�ȷ���⺎�P;(#�;��0<�9\<�=}<���<���<l�<�_�<�|�<���<�F}<��\<��2<uK�;�kj;}���Kڻ��H�aĎ��:���hü��ļ�ѳ�V����WU�Oh�}�q����AY��K�]�j���\JN�Q!�����eƼ�Ǽ�!���旼��^��!��A���:Fc�;��	<��,<@]D<g	R<�V<��P<��B<H,<i#<1�;9�U;���\������v� �����ݼ|��X���R�%��1F�`�N���P��$2��7ԛ�&!����ļ����S��7'�x�8���A���A�צ8���(���- ��ؼ����5Q���ֆ���p���]��RT��S�5n[��.k��o��9G��0���3��kMڼ�A��� �� *�UB�X�Y��jm�G�z�.��q(|��$p���^���K�q;��1��0��8�UbJ�@Ua���y������,��T���̐�8-��^���[q��5]���J�&�;�@�/��m'�ݫ!��:������d
 ��H$�:L*�2�J�;���G���U��Bg���{�_���t�����=Z�����XM�������֟��{��E銽;��$vz�
�y�-���d≽�b��9ꞽo��&S��˴�������Π�!������ʣ��'�m�Zv]�ukP�>TF���>�cF9���5���4�|65�4�7�:j<�!!C��L���W��f���w��h���͑�p7���Y��Qɮ�M��9<���ū�{���#���z����[���#���Ʌ�������n���}ݪ������3���>������n��t�����������6�|�Cn�nGb��RY�O�R�62N�k�K��HK�{�L��/P���U�IE]�v)g�O�s��  �  ��<��;���:>O�T�˻���1=���E�'�1�n��|;��'uI8�/v;��;+��;���;�G;����̻��'��T��Gg�BW]���:��6��V��g�I�Eg7;� �;!p<͘6<KX<�0s<�J�<�k�<��<�߃<��t<P;Y<}�6<��<|�;�{0;s�������9�L�W0{�����ø����r��<��(ﻣbH��'�9��;��$;��.:�W2��%��8���q��:�������_���\��f#��ʻ�����x:/_};o�;��<I1!<k2<��9<�6<Ζ(<R�<��;#6�;�5�:X��,}���"���h�����＼��ܼ0��_\������u��2�Ҽ�>���ė�����M|�+����e��J*Ǽ�����_��F$��%��� �j'�����w��4�ؼ�ؿ�����@O���1������ʹs��o��-v��i�������E��Ef��Cϼ��gW��[���$�0c6�JMG�l�U�,_��/b��d^��WT�F�O�6��)�J�!��w!�|c)��d8��K�	�`��Vs��n������Dt������t��Qg���Y��L�>�A��t8��1��'+���&��$���$��'�(�+�J�2�F?;��[E�ТP��]���j��@z��L��惍�����V�������"O��yX��ol���ŉ�f��:�s�~Wk���j�Npr��)��߈�j����昽RO��+9������)f���M���q��RO���p��Ad�]FY���O�X�G�łA�;N=�U|;��+<��X?��D��]L�z�U��`�5:l��z��Ƅ�(���*���S���s��+����>��w������|��8X����~�n^y��3|�{O��CE��Lp�����A����>���-��dԣ�����ݷ������������j�u�|k� �b�ʈ[�� V�7�R�"R���S�X�/j^�f�f�\sp��{��  �  ���;:�;8��:Y���+���R`�����xk��̗���;bݮ;�<�%<�-<�<�Q�;�t;]��8��S������h��'ﻞ�ջ�[��QP�;M���|:�+K;M��;���;4� <ްA<�2[<z�i<��j<4�^<�F<B$<#L�;MϨ;�^1; t�9ޤ�����)ӻ�r�*&���%�:�'/��J���e�����:�b�;��;���;^�;��;��������!���v�4W+���&�8�Ya�=[��t�W�����P:�9;���;��;1�</�<<�<�u�;~�w;�0P:�_�����& �eA�xEp�HŎ�����f]���{����ż�����ǲ��杼"J����a��VE���>�(R��u}�i��܇�����;!���4�J�!�
����u� �=�6Q�`Bռ�Ƽ���������4��WL��:���Uύ��ᖼDs���'���	ӼL	�,N��'j��`$���.��^8���?�E�D���D��@�338��,��0!�Sf����b�N���%���5��CG�D0W��c�W0k�g�m��fl�
�g���a��D[�'tT�ۨM��F���?��99�Ռ3���/���.���0�h:6��g>� �H� �S�'T_�:Kj���t��~��&��t����y��a�������������Ʉ�T�{�S�m��2b���[��X[��Da��8l��z��,���J���w��$D���Ǐ��y�������څ�~~��>z��q��g��R^�m6U�^ZM�#�G�<E�f�E�`J�fQ��Z��#d�cn�gx�q���慽K����������t���nY���\���	�������Pw�W�m���i��Fl��t�Y���U���,��� ����ƙ�ј��:��z���Ȕ���X���	��/���8)z���p�Wph�*ta���\��[�Q�]�W.c�%k�y�t��$�`����  �  	;tI:��X�/���Ҥ$�ק����8w�:	o7;[��;���;=^'<�"K<F�a<��f<��X<�A:<��<%�;��F;�':ĵ��.��L��(d��i���Y��a/��]ĺ@5�9�u+;bq�;�� <1#<}7<J�9<"�)<?	<f��;�):;���8�v���x��ȟ�3���\=���2��|��������R�����a�:���;cm�;b�<o� <y!<_�<���;G�;���:;P��MY��͜������˻�'ѻ��λ4)ûR�������e�Q�8�2;A��;�,�;n��;Б�;��E;�F��]�i�f"���-���Z�d}��؊�������Xw���ڙ��f��a����}��[��8�s���R�_��;z�@;�y�l��������fȼ�ܼ]�뼳�����������d �{������q���߼�%μ�=������D���¥��쯼 �¼�$ܼKy�� '
�~S������&��+�Gm.�80�*[0�6%/���+�({&�������W�U���5��a��_
����N�!�6"0��>�=�I��[S��'Z�3�^�E�a�0�c��td�4�c���`�ޒ[�baT��L��D��>���;�TS=�-�C���M��bZ�ǲg��t��A~��ۂ��J��ɪ��j=��m&���X�����Q�I{���p�ze���Z�!�Q�$M��L�)LQ���Y��`d���o�v�z�����ް������������Dꇽ	��H��p\��&n|��&r��g��\�0(U��fQ�WR�'�W�@a��pl��Ex�0~���ą�cψ�����nы�2?��:���7��b��"^��}"����y��o��Ye��g^�*�[�5t]���c���m�VWy�h����އ�.����䎽����O�����%ᑽ�琽�쎽����nZ��!��Ȅy��0p���i���g�+�j�ĭq�q�{��냽�Ή�ꎽ�  �  ^j��������t�׋�H��H��:��e;F
�;n��;p$<
�H<~j<NT�<�R�<+Ӌ<T{�<�u<ΓT<Pj-<=<��;��L;�VB:jҺ}�|�	���I����$��I�ǻe���{��J;�;C��;$d <��;v.�;`�:^�F��4˻R�
�:�F��q��\�仦m���>��?���:(w;N`�;B�	<E+<D<8ZR<��R<��E<-<��<�T�;0�y;��:ܓS��H�釬����)��~-+��1�	�&��	�B����F6���^7;�4,;�{�:h�]�����`��W�9,��]��������������W���0������Ie�H�N*�|��k���q�� ����x���`˻�k���+��[�f���W����跼��μ���Q�������`����1����	����� ��Mм�bü����f~ͼk�������:#��"0�Z8�;�[X:���5�ݘ/��k(�, !�����"}
��(�̚�����҄�"����I'���7:��)��H6��2B�>�M���X��c��|m�h>u���y�.z�;�u���m��b�x�W���N�u{J�j�K�t}S�x`�'�o�o��.��:$���Ŏ�>�R���ω�>���2X����y�OGp�u�f��\��AS���J�kED���@�"�@���C���I��dR�� \���e�ǫo�R+y�(C��>ۅ��2��䍽<Z������D���3��x;��Ŝ|��Ko��e���_�-�`�b9h��0t�fS��C���?���׀��/���_�������t��dg��l%���π���x�n�o�{ef�u�]��=V�^>Q�^WO�[�P���U��9]���f�t�p��<{�ͨ������(p���)����������%��ʘ�S&���ݍ����׀��"y��4v�Χy��o�����ρ��˄�������  �  �5���/�Hf�����|��[��:6�;|�<
7<��^<�h�<FT�<�}�<x*�<^�<d��<#��<+E�<Y�f<m�><j�<�b�;�q;������»����R�#�o��Ks�})Z�w6(�Nͻ�A��0�:�Dt;��;@a;�Z�Db��Q���iY������\���z�\�X��"�Эǻ'M�a�:}}�;�i�;\�<Eh@<,�[<Zo<�/y<�sy<�o<6�\<��A<� <��;��;ʓ�:�U��ZȻ��$�9�^��y��K����H��
7}���H���	�G���{������e��~y��~I���p����Bļ0ڼ2 �Gڼ��Ǽ��������{n���<�%r��޻]s��X�s�SI;���'��=��u{�հ�t�����$��4T��I��w������s6㼚j�ٝ�(j#���-�i2��U/��&��K����L������`X�!T���eq��#,�k.?�@�M��%U��mU�t&O�dD��S6���'��G�dC��$�r���U^�.��p�ڼ�'ڼ�y޼ ��28��a��U�ß�v.)�2,8�?�H�`jZ�R�l�x�}��ㅽt����勽Z׉��Ȅ�'�{�"m��a�:�Z�˔[�wd���s��u��b:��������y���^N��ϔ���ɏ����	���?q���c�\X��FN�̡E�m�>���9��7��6�9K9�<>�.�D��sM�wW��c�Cp��2��������# ��j���������Mř������	��כ��kv�zao���p���y�Zo���s��GC��=E���G��9���\ڞ��Q��)���c��=˂�T�w�U�k��a�^X�otP�>�J�JG���E�1G�o�J���P��X��5b�O)m�B�y�����ދ�2���J���:��d���e�������si������_$���D�������͂�;ꄽv������x5������(ت��  �  ����>���ao���'�S��s��9��;��<,W<>�<*�<�<�<�Q�<���<��<���<��<�0�<Oc<e/<���;P�:DSa������l��#��b���V���e���ʊ���F�MZ�X0�������9+Ⱥp��R�,�V����,��O�X��������ڗ�ba�h��XJC�ϔ�:��;o�<|D<�<e<>M}<+��<�|�<i��<�̆<�~<`f<�F<��<�u�;�
;��4����@`�|q���5��aʼ|�ɼ���h���'d�����_Ļ4��YU���l�Ԭi�b���4N׼�J��0�
����O���/�7|ɼ�t����q���,�����F���!2���ƺ�Rg�GVP�s �x��m�h��o���) �Cp/�dh��a��o��� �I;���%�jw:�j*I��O��DM�f_B�À1�?O����'������t�R)�;^,��D�s�Z��k�Ѩr�Y�p�8rf���U�Z�A���,�qw�	�?�����׼
rϼķ˼�f̼I@ѼMڼ���à���4����{�!��"4�fYI�.�`�۔y��~��R?�������#���z���1�.Ѐ��sr��j�ӭj���t�-k�����FB��i�U��Ū�������y��?�������!�����n���]�\�O�Q�D��p<�%@6�'2��0�60�g�1�t�5�$�;���C�b�N�`\��_m�~���1䋽�?������dl��/���h#��.@��Ο�8s��:=��HA��`~����}d��3q���E���ţ�O�H��h
���c���>�����鍽_O��M�s��Jd���W�?�N�z|G�'�B�5�?���>���?��C�?+H�K_O���X���d�� t��P����͆��Pޤ�����:����g���������<]�����^������ =������������������;���;����  �  ��ɼ�N��렢��?l����q���$�;�w"<�<f<�e�<�Y�<\x�<�ݱ<fK�<�X�<s?�<��<���<(S�<w<B<<���;�đ:����R�I�����X�Ƽ��ۜ��ڼ�U��1���s�7��˻�M��-�����O��ngx�sŭ�ST׼����L��Y伹#�������X2�D=�����:�m�;{ +<6Z<��{<��<�<�N�<�W�<%6�<Fo�<�|<��[<�.<߲�;��:JY����,��捼���̯��.��F���aE鼺�ļ����Y�*���� E��L��ԕ��μ�Y�s�S�$���%��`�Z'
�)����������,���л&R\��^��ׅ.�pl�9R$�9�8����j��������Ի����Y�_���r�¼�X������6���O��a���i�Cg��yZ�n�F�p0�y/����-����x�$���=��|Y��vr��<��`6��������{�d�f��M�P�3����������0�ڼ�̼{�ļ�'¼C�ü��ȼ�XѼ�Bݼ�(�:� �4���Y�3�}�L�Fi�`}��O����n��JC�����Bh���:���(���s��������v��Rw��C���e���4���M��D��>��Յ��^i��a����s���ґ��G��|p���[��jK��p?��6�s1��i-���+��+�.-�
�0��:6���>�)J��Y�9n��5��uѐ�ƻ��g�����O���!���������,��S��j&��y��oM�����_ٖ��?��UB��/���M��裼����뗬��ߟ�iF���D���s�F?a��)S���H���A�>�=��";�Ƌ:�j�;��6>���B�B�I��S���`�-�r�0R��C��FO��-��7��Z���YŽt|ýے���
��������`D���x���C��!��…��!��猾�Ďƽ�  �  C���6⼏���o���z'��}9�>s�;e� <I�k<|C�<��<�+�<3�<6��<�߹<�<���<���<;��<4�<�q@<C��;���9�O�Qq�O������r������;��n�ؼ?0��P�e����W��5B��P@�:C��{���a˼
���
�cF�o�7�ܼ[��2ZR�N����)�:ǭ�;]Z2<E�d<R��<���<��<+�<��<�/�<���<)�<L�f<��5<;��;��:_����=K�砣��Iܼ������g��M���⼐{��с��5<��E��a/��7q�꫼yr�l��)�o56��$7�],��_��9��f�����Lv0�w�ɻ�Q9�O/�$!:�˄:�sn:��9	��s��De��$��_8�F7S�����dȼ�5�D�"���B�Tf^�;Rr�Mu{�m�x��j�j'U���<�^R&�k�d���� �.���I�Zug��5���㊽�
������^���s�N�V��9�ϸ�::�0ּ^Ǽ`L��b��W8���ļ��̼(0ؼ��缙^���������4�}P�G�o�Vo���%���:���歽S������������7��e��͝����ԅ����������������� 쿽{X������Ы������ԕ������r�m>[���I���<���3�4?.�'�*�g)��W)���*���-��S3��;��:H�fY���o��n�������0��d[���6��MýB�½^
����O���W����������㊊�MA��_w���墳�������z0ƽQŽ!����<��5���O���)����t��``��Q�6F�J?���:�C�8�G8��69��;�g@��F�sQ��j_��r����� ������r(��*����ʽ7ν�>̽��Ľ6�� �����&���韔�c����!�� w���.����ƽEϽ�  �  	@�:��;"ܛ;�G
<��Q<�=�<:��<���<���<\��<���<,	�<�L�<j��<���<��<6�<���<���<D��<9P�<�F�<"��<�`<G<���;�U*:H�亏��D���ӱ:�p�;�<��E<S�f<�Ck<��R<��!<���;[��:����,h���~�r ��*:1�;�<s�]<e�<�ũ<�v�<��<|��<�}�<���<&��<�v�<�<�<���<f�<I��<o!�<�~�<m�<��Z<�<��;n���d�Rذ��ƶ�K���B���$;�l�;��<��<�<�!�;ݘ:Ѧl�����D�"Ri�@�o��PX�Z)���ֻ�!�~�:<�;�|�;H�<W<��#< !!<�<��<>�<Z��;Vf�;$��;��!;��=��$W����C��銼v����ּ������ ���mu켆�Ӽ���df��o0���A���@������s|Ӽ�����0����7� �9!�.�������r�μ���������S����q���f���d��i�y�q��E}��q��
�����������HƵ�aJ̼*���[���.�'�B���S�+g_�`d�h�a���X��JL�k�>��4��4.�	:/��b7�wE�	W���h��x������΁��/~��Hr�o�a��vO�V2=�$�,���w��x��h'
����$I�y�����hs�����j
�^��޲�z����,�{U=���O�.c�w�t�~��J�������";��E�u�b f�^�V���J���D��F��ZN��&\�[�l���|������͇�)S��.K��T�x��g��"U���C�`�4���(��W �(��_��z���q�,���W�<��m���]�G�"�l/+�ؚ6�aE�
W�gcj��}��$��`���Ï�޸���D���b���w��h�~�^��A[��&_�s�i���x��c���z���  �  ��;�P;���;�<*�Y<��<�3�<u�<۔�<_��<��<bE�<X��<��<MU�<~��<xS�<��<���<a?�<�B�<!��<y�<�f<��<�>�;��:�a_��Rƺ�WṠ�;9�;�<H�M<S�m<2r< HZ<��*<���;_�/;�"�'-�,aC���Ϻ�P�:�;J<�b<u��<��<D�<D[�<���<���<�7�<��<���<���<��<���<� �< ��<���<M%�<�6_<�<�>�;՞:w�-��^���Q��":S�Ju��0<;���;n[
<+|<L	<�N�;�F�:}hA������6�R�Z�za�~K�C��?Ż�����:,�;o?�;�w<F�<U$"<Ш<XK<4�<w� <*X�;1��;'׌;Z�;�\��8�R���=(>�V↼� ��c}м.��9��T�����)�ͼG����/��(���f懼Ĺ��槬�:�μ��q�
��R���֕�_��-�e��p�˼�2��������� "s�9Lh�2f�Ujj�r�r��C~�����O%���@���9���,���7̼1輵�W���,��@�~P�U�[�J`���]���U��mI���<���1��i,�2|-��|5��>C�(gT�m�e���t���}�T����z�35o�ym_���M��<�pH,�%g���|���
����9����$�;���/��
��,����ɇ��b,��><�(4N�ѭ`�̏q�u�~��؂��悽
�~�&�r�@tc���T�d�H��C��ED��cL���Y���i�Ȕy�J؂�
����|��A���x�u��Ke��S��B�j44���(�ԕ ��%����%K������ܢ�l���,����xB#�VN+�^d6���D�e�U�?lh���z������Q��z卽`䌽���m恽t��f���\�~�Y��Z]�w�g�hzv��y�����/���  �  �;�׸;^��;/�2<�o<�<S˳<6��<�\�<��<]�<���<�C�<��<�i�<bi�<9��<�c�<��<��<�f�<N�<�̚<=�u<��2<S�;�Et;���:�^�:1;#P�;�;�5<��d<Mƀ<̂< �o<��C<V=
<��;���:I�ĸ���	�Q:�m\;"�;Ӣ/<qKn<	�<g�<�n�<?��<��<*�<���<�#�<��<�b�<+8�<z��<�d�<�<`�<�S�<�j<��)<�R�;D�*;�>��c�Z���QZ����:���;Z��;|T<�d+<
q<���;�W;օ���j��'_�31��k8���%�:[�����Q�����;���;v�;� <�<@�<��<<<��	<���;��;���;���;P�;�BY��^M��ڻ_0��Qx�蜟� ���Y}ռ!���߼�pҼ�＼�?���A���Y����|�q������9�����㼁���-�d��.���
�����b��+�ļ����0`��b҅�D�w�Էm��dk�:�n���v��܀�
ׇ�@S������	���B	����̼6��y��?��&��A8�B!G�&aQ�S�U�o�S��:L��UA���5��;,��V'���(�50�e�<�z�L�F+]�_�j�cVs��ku���p�Ĵf���X���H��9�.�*�Qe����/�����<	�%��(������	u	��-�(w��������D+�׀9�'�I��Z�@i�y�t�>I{�V{�u���i�)�[��%N��~C�=(>�YP?���F�C4S�tb��zp�o�{������V��M�y���m�b*_� ZO��X@�f3�K#)��!��z��G�7�����m�����3�i~���Vv$�[�+��%6�"C�	dR�"'c���s��$��2T�� ���+����Ƀ��]{� fm��`���W� �T��>X�P�a�/uo�p�~�6�����  �  <<c�<��1<�U[<�R�<X��<c�<έ�<�X�<�<+~�<�!�<���<���<k��< 2�<7��<h��<=�<���<`��<��<��<xʄ<�4R<]p<f��;v��;{ �;���;��;��,<�\]<�@�<{��<�^�<u��<��h<՚6<��<�
�;��o;hW;���;���;�<�H<~{<W��<h��<ƶ<f�<D�<���<.y�<(�<���<&��<t�<&�<��<���<���<�L�<��u<|DA<k<+�;�%H;�M�:50�:B1;9��;	��;�!<ܜ><3�G<	9<n<b��;�R�:_T�ލ��������Ӕớ����Q(��9#9�%4;肢;RP�;$z <�<�<H�<W�<�Q<��;o��;��;u]X;���:1�4��FW��uϻ� ��+\�ȗ��2y��i}���¼�����󵼕ϣ��􎼙�x��'b�0(`��lu��܏��C��=2˼�r�j��b��U@����8�鼺yӼR�����������≼`i��;Uy�qv�nx�	`~��r�������֔��ߟ����r༼%�ϼM���u ��-�(���K-���9�okB��!F���D�6e>�G5�j�+��#����W(!�4(�ɔ3�2�A�D'P��:\�*�c�)f�l�b�;�Z�raO�B�t�5�,4*�*� �\���
�%��Y����	�q	�Q	�
�O	�G��[�r8�@� ��*�6�6���C��4Q�#�]�}g�G#l�6�k��pf���\�БP�M�D�o;���6���7��|>�WI��VV���b��l���q���q�~Xl�~�b�L�V��J���=�	W3�P�*�;/$�Oh����s��r����eq��1�%"��B'��.���6�(�A��vN��>\���i�7�u��@~��������]y���n���b�-�W��P��rM���P���X���d��Mr��^~�;v���  �  �U<�+X<�{i<�ӂ<oܓ<��<�&�<���<�L�<8��<�*�<���</��<J�<���<�<6��<L6�<���<���<kf�<n�<���<�\�<C�p<��J<i7,<�_<�<�[#<�u?<`+e<J|�<@L�<wn�<L��<r�<Wb�<�k<h�?<Q�<%�<-��;�<�<�X:<�u^<�N�<���<=��<��<���<E4�<��<���<�n�<lM�<�<N�<��<z��<R�<a �<w��<,,{<W$U<�U.< �
<c�;�K�;���;Q��;.�<��-<��M<k�c<�i<��Z<:�9<#�	<*��;�_�:6)���Z9���j�Y�iv���)�@�:�'<;��;�|�;Dt�;6y�;"��;���;���;I��;�n�;^{�;Gu;�	;:��9�躺H����ӻ�&�^,B�\�m������$����o�������/��h�k�?�N�/
>��f>��R�-w���������)�Ƽ��ټ�A��0��`�y�Լ:Ƽ�涼T���ϓ��x����Ћ��冼�)������ą�����S������⨼��Ƽ��׼��꼖����+�M��C�!��
+��}1��84�6�2�� .�%'�"{�{�W���f�����z(�ܐ4���@��0K��R���T�3S�I�M�F��=��3�J�+��$�M���K�h���D����d��g�����a�����t'�[�$��[,��5�}�>�lJH��Q�Y�W���Z��&Z�HRU��*M�]6C�Ir9���1�i,.�/���4���=��}H��S��`[�'`���`�}]��W�w�N���E��H=��5���.��B)�~�$��� �9�����!����Y�@�"��,'��,�M�2��:�ozB�5�K���U��_�`2h�n��_p���n��h���_�vV��M�y�F�X�D�x�G���N���X�b�c�G�m��Iu��  �  rJ�<�
�<���< ړ< �<n'�<gt�<"ҷ<J�<{��<bT�<F��<���<F��<��<!��<�}�<���< ��<ü<9ڰ<��<�i�<#Ӎ<���<�p<f"a<�NY<)�[<T9i<D^�<�Y�<�ٞ<�Ϋ<���<f?�<$��<��<xU�<)�}<:E_<+iI<0~><	v><8vG<D�V<�i<Ý|<�F�<'X�<���<��<��<�ݹ<
��<�g�<�U�<�o�<,S�<=��<�`�<_^�<=c�<�}�<�/s<�_]<�1H<5f5<ݳ'<��!<��%<,�3<��I<�&c<�Mz<���<�u�<=}<D`<��7<�d	<���;a�N;�߲:ɠ9`y�ޥ9��-:+�:�j;�A;�:t;'`�;r�;���;Vx�;���;��;U��;;�x;-�
;��q9R�byr��d��z����b�2��M�2c�9�r���x�E0t��e�C
P��8���#�h.�!� �-�oM��Vv��b���8����\Y¼m�Ǽ��Ǽ�:ļ�U��!���o���J����
��9���W����ڑ��6��/���w����P��/������hƼ�ּ[��3?�����},
�=e���`��6R!�n�"��L!�Z���y�� ���@��or������'��21��:��q@�x�C��kD���B���>�&Z:�gi5��T0��*+��%�9� �Qp�5��U��d�n_��K����K��^� �	u&��,��1�Q7�|<�h�A��;F��UI��GJ�̐H��D�\n=���5�"�-�r$(��R%�(&���*���1�WY:�]�B�o�I���N�Q�P��O��4M��AI�ָD�E@��B;��z6���1�X�,�9D(��u$�b�!�:!��,"��&%�ݘ)�r /���4���:���@�E�F�ˇL�KR�"�W�"\�g�^��F_�!�\�w�W���P��0I�=?B��=��<�wW>��C���K�F�T�:8]���c��  �  @x�<*У<���<��<�՛<) �<���<�Y�<uy�<+2�<���<�2�<���< ��<��<�g�<��<�h�<�]�<Tۤ<�T�<��<Xa�<H��<h�<'��<�$�<��<|��<nb�<}��<�q�<N�<g��<v�<!O�<�/�<<t�<���<��<&�<C�<�v<r�k<p�e<M�b<eYb<��d<�k<Ȗw<1��<C��<�(�<�#�<.��<���<��<���<�<�y�<�S�<Y?�<2�p<��b<$�Y<WHT<�Q<!Q<��R<BX<��a<S�o<��<gƉ<Pk�<���<�ϔ<g�<K��<��a<J&;<"�<�`�;+&�;�c;<�;#��:h�z:�: ��9d�9��Z:m�:�� ;;�`;cQ�;���;���;�c;9��:�T������_����ֻsv��"��!*�>�4�3<�,�@�?�A���>��m6�Ԇ)��|��J	������L����z$���'��KI�)n�� ���ژ�����y��u����w��0뾼i���x@���Q��躼�8��G.��G]��V���R��L����ԩ�z跼�Eɼ�ۼ��p�����	�#��E5��<�֜��!�͋�������?���X���'�wC�.��Ǵ�����#��*�Q1�s�5�� 9�S�:��;���;�G;�8�9��i6�f�1�,,��%�������S�b	����É�8�%��a,�6y2��n7��;�gZ=�٦>�`6?��'?�Y>��<��[9�~�4��>/��&)��|#��>��A�����\!���&��-��e4�F�:���?�	MC���E��G��G���G��$G��NE��$B�ɟ=��8��&2���,�f)���'�$)�+�,���2�_�9�g�@���F�ڹK��AO�ƏQ���R�B�S�"�S���R���P� �M�[�H�9CC��o=�Y\8�b 5��4���5�AB:�qh@�ikG�:QN�2ST��  �  8��<�<�7�<���<�(�<���<��<`�<E��<���<��<�W�<ɴ�<�5�<#��<?�<��<���<��<^��<<>u<Q�g<[4e<�l<#�y<�]�<2��<��<ڪ�<6V�<' �<	��<�G�</��<(��<r��<��<�X�<���<���<4�<|z�<�<҃<ARq<e�[<�H<^;<�6<%P;<��K<h�e<��<V��<i�<6��<pŦ<��<���<Ic�<�qc<�&G<��3<��+<`�-<W�8<T;H<�3Z<�ol<~<;v�<�<!��< p�<��<ے�<�X�<�Ě<L�<��<�vc<��@<WR<��;Է;�[q;���:�k�8_���Ո$�AH��BA���y�����9���:ī";J ;;��:�M��.O5����g���(�=�@���M�ٖO�`XI��>���0���"�������Xo�8�ڻƻ�9���7��}9ƻd{���w�$���C�'�c��������Vӟ��>�� ����ȼ�Ӽƈڼ��ܼ5�ټ��Ѽ_�Ƽ����B���vS�����X��/&˼�:������L�����v��v�x����I%��1��W����V��u �=!���R���d���} �����"
���ի�����g%��+���1��7�&y=��BB�^�E�#�F�%sE��7A�:���2��w*�V�#��; �� �/�#�f*�I2�2�:���A���F��H��%H��|E��rA��<��7��2�<�-���(���#�S������'���>��������#���(�J�.��t4��=:�E @���E�)K�ȪO�k�R�zlS�asQ���L�f�E�L<>�F 7�\�1��/��I1��\6�|>���F�q]O��6V�ًZ�\��#[��GX�tGT���O��!K��sF�j�A�?�<�T38���3��90���-�-�K�.�F2��6�u<��pB��rH��  �  ���<lG�<q"�<��<���<G�`<VK<��D<�(O<7�h<br�<�@�<ᡫ<Mض<@]�<�m�<�9�<���<�p<��I<:�.<#�#<W�(<1�<<FhZ<@}<[�<Pܠ</Y�<#��<<��<G?�<E��<cl�<r��<|l�<�g�<���<Q`�<���<ᾶ<���<�P�<�߈<@�k<��D<�n <AH<���;jp�;L<��%<HM<��u<�h�<:Ɣ<���<���<��v<0�M<��#<��<@�;]��;�d�;Q�<�g.<��Q<Ht<�O�<Rܕ<��<���<�ϫ<,�<|ڭ<���<��<k��<Ƌ�</f�<��`<��=<ǒ<�B�;-�;k��:�X庉~���ʻB�컐��u�ѻ�C����7�@2����%9%�9�8��8�y�������RE�X(m����?��W~��хm�[�P��2����Bw����λ�)��Mq���p��bn���O���8��~����h�j	��$���B�nd������瘼����*ż	�ڼ�����js���������E�k�ӼqTƼB�����{�̼9X�����
���K���#��2$��!��H�@���(���W�����X���I��H�-��2�������������7	�!e��8���'&��g/�.K9�z@C��VL��[S��(W�C�V�[�R�ՙJ���@�I6�v�-��()�(�(��w-���5��@��|J�ZS��)X�p6Y��BV�7P���G�¦>�d�5�%�-��w&� ������lw��q�ݥ�X8��#�>��]�=k ��g&��i-�|�5�Q�>�9�H��gR��[�Zpa��Ld��c�t�]��hU�X�K��'B�3O;��{8��_:�G�@��NJ�vZU��_�\�g�M�k�"�k��.h��~a�!Y��FP���G��N@�'�9�\�4�M(0���,��(*�ػ(�4�(���)��P,���/�H�4�:��~@��  �  ��<���<�ˡ<��<2V<�l(<�i	<_�;��<c'<iS<��<
�<�ߤ<,�<��<�؍<�=j<_B5<�<��;_�;���;*�<[�2<�d<b��<_��<�ڵ<��<�Z�<�r�<���<|+�<��<N�<���</h�<<$�<ex�<���<���<d�</�<)�Y<<e#<�,�;&��;��B;�/8;��;���;�\<�G<6�o<�D�<4��<|qq<��I<G�<���;]t;2�;��;�_;X�;V&<�><��n<��<�1�<0@�<a�<�7�<�D�< ��<]��<�8�<1��<�ޖ<��<��t<�"P<
w$<���;�^;J'Ĺ�K������$���<��,?���,��,�SĻVp� �
���躢�:����L9��$K������9���ɥ�S������*ڌ��n��@�d+�c��)!��V熻��a�^�O���R��h��������Ļ���F��^�.��[S���~� Ҙ�#U���bӼx������#q����	�Up ��%���ڼ��м5�Ѽaj޼s ���4	����lx&��Q0���4��3�Y4.��%��/��N�ަ��������'�z��\��˅�{����６��������>��
�"�֯�P$� 00�J�=��xK��?X��Qb��%h�P�h���c�DeZ��>N���A�q�7��1�V�1��7�^A��M�{Z�23d���i�)bj�܊e��f\��{P��|C���6���+�)�"�b���L�z���'�����S���U� ��P��'���!���)��^4�ʰ@��DN��[�-h�C>q�8�u�$�t���n�ϐd�Z�X�M�p�D�;A��DC���J�TV���c��o�1:y��}�G�|��v���l���`���S�&�G���=���5��d/���*�]�'�u&�6%�ZK%�S&�8M(�xB+��Z/���4�0	<��  �  {�<xP�<��<�un<�,<���;Ý;@)�;?~�;*t�;2"<�Z<���<��<{��<�w�<��w<�!?<V�<���;�G+;+� ;%>;��;��<n�I<��<�E�<ɔ�<-_�<���<iK�<AA�<Z��<���<U��<��<�q�<Q��<�O�<���<���<�<��<�XD<��<��;�7�:_75�(\z��Ϸ92	B;ݿ�;w <�N<�h<q�i<��P<�5#<A��;oA;i�	9�����c��7}56;���;
�&<e	c<�u�<Ű�<��<N��<L��<���<���<��<s��<���<<��<jR�<_�<߀X<6�'<�Y�;�%;�J�O�ӻ��+�� ^��Uz���|�n!g��>��L������>���h����`�ﻕe5�'�z�������\ļ�eļ����6 ��Sd����R�~��;8�,z��xc��J3�9�#�y�,�d�G�@�p����������ٻ���$�@L��k}��m��Y��b��� ��--�b� �
,�t�����~Y ����z�߼�߼D��l^�߼��%�q�4�/Y?�6 D�VB��d:�?�.�� ����`�����e�@8�v��3k�۸�k�漶���(�#����T�@�[���=-$�ɮ2��B�3�S�yc���o�� w�0x���r���g���Y��K���?��G9��9��2?�E�J��X��Ug���r�']y��|y�2Os�E�g�<Y��6I���9��-,��>!�p��d���������]�w��Q��#�6g�^M��R�U�(�^D5�?%D�^�T�s\e��Ht�hd�-~�����~#}�smq��}c��BV���L��_H���J��]S��}`� �o���}�"�����������ف��Xw��Kh���X��I�Z{=��3�Z�,�(��#%�d�#�U#��Y#�!C$���%�h�(�k,�_2��:��  �  .�<���<���<zX<��<n�;z�;��:�;v0�;,<f4><f�s<k��<�<m�<T_<#7"<�3�;��;���8,����9''J;��;�*5<�/{<�4�<8�<,��<�n�<��<(��<��<ʎ�<%��<�<���<Ց�<���<���<�B�<AH�<�cz<w'3<	��;@r;�%�R���f��`	�o�E:o]�;FA<��8<�3U<h-V<;<�|	<�n�;�J:Q��!A�����O�ןG:���;+~<S-X<<�<�ޟ<���<��<��<<E�<ه�<�µ<~s�<���<��<ӑ<��<lI[<QO'<���;:�:��Q�O��`N�����Q=��Tn��E'����a���+��l��^�����{�����aP��e��<p��W8˼UBټ��ؼ�Fʼ�<���𑼟b�%�?��M���~�Q����q���P��.8��Db�\犻ʩ�.�ϻ�h ��f ��)J�\z��R��E�ż¦�E*
�����M&��a+�6h)��.!����0=��J����鼆t�G����H	���!u-�7�=���I�T[N�<�K�gC���5���%��$�/��E��Y�꼳���ݼL�ݼ�S�$��c��n��r������ҷ��{�����%�F5��@G��Z��|k��Ly�/����L��S�|�P�p��a��"R��vE�G7>�i�=� �D��Q� �`��=p�|�|��끽-��|�--p�X�_��M�fc<��6-�y!�m$�5��Z�DU�{��d��������~�������(�#�6�0G�T�Y�:l���|�s�������OH��Op��\z���j�qo\���Q�p<M�c�O��Y�?Ng���w�K���9���̋��͊�s����
n��u\�� L��>�G3��+�f�&���#��n"��"�nd"�f=#�|�$�w*'��+��0�υ9��  �  ��<,��<�׎<�O<��<�U�;ڎ�:�,�9+�:�Bq;*�;g4<2�k<���<N��<�d�<��V<o<I:�;M�:�U��kź��ιߪ;!�;nt-<�!v<�ߛ<�ֶ<:�<l�<���<���<���<�#�<+n�<ܻ�<8��<�X�< ��<�^�<5�<�h�<�qv<k�,<| �;���:]���Æ��"��$B��[̷f�v;��;��0<�@N<�EO<�r3<�l <0Ӏ;w�6��N����4���O���7"d�;��<W�S<�2�<V��<��<4��<�ѽ<.�<m�<�>�<��<>�<<e��<̦�<b�[<̥&<"��;_|�:}�o�+����Z�<�\����Қ����t�m��E6��f��+���N����λ��	�Y���������dҼ���K�߼h�мmѶ��A���h���(�ҕ��n��ۜM��I�?��e�ح3�!%^�ﱈ�[4���ͻ�����P���I�TR��顼��ȼ������ ����)�/��-�8{$�����	��U���/�7���I��:`�TR�hi0��XA��2M�9R��lO��)F�))8���'��g����1����꼽�/�ܼc�ܼ�߼� �lI�]EＡC���
��tY�>�6��t%��6���H��V\�\en�J�|����*)������	t��cd�JqT��hG���?���?�l�F�>JS��Jc��as�},���ǃ��ȃ�x-��(s�vb�)nO�8q=���-�#!�������{������)�W�W�����w����ø��[��)�\<7�qaH��w[�Ƚn���o_��p���h ���(��}��um�|�^�b�S���N�ߒQ�C[�E�i��z��,�����Z����������8怽�Ap���]���L��e>��;3��Y+�@H&�(g#�"�R�!��"��"�.a$�@�&�D�*���0�hr9��  �  .�<���<���<zX<��<n�;z�;��:�;v0�;,<f4><f�s<k��<�<m�<T_<#7"<�3�;��;���8,����9''J;��;�*5<�/{<�4�<8�<,��<�n�<��<(��<��<ʎ�<%��<�<���<Ց�<���<���<�B�<AH�<�cz<u'3<��;5r;�9�R���f��`	�ȣE:T]�;5A<~�8<�3U<B-V<�;<�|	<Yn�;˻J:S��dB��U���hS���G:�;�|<�+X<n;�<�ޟ<X��<���<2 �<I�<4��<ʵ<�|�<f��<��<R�<{�<ts[<�}'<��;n��:��P��n�5+N�'ǂ��%���X��a����a���+��I��J����������s��#vP��s�������L˼0YټS�ؼ�`ʼdW�����ELb�FF%�I0������AR�Km���K���O8�yGb��ي�6�����ϻ�K �C �D J��K��9����żR��
�9��A&��U+�v])��%!���Y7��B������t鼢���M	�*��}-��>���I��gN���K�gC�֤5���%�3��<��^����꼖�Ἂ�ݼ?�ݼ#a�j�伔�����'������e��}�o��=%��5��@G��Z��|k��Ly�7����L��]�|�X�p��a��"R��vE�I7>�k�=�"�D��Q�!�`��=p�|�|��끽-��|�--p�X�_��M�fc<��6-�y!�m$�5��Z�DU�{��d��������~�������(�#�6�0G�T�Y�:l���|�s�������OH��Op��\z���j�qo\���Q�p<M�c�O��Y�?Ng���w�K���9���̋��͊�s����
n��u\�� L��>�G3��+�f�&���#��n"��"�nd"�f=#�|�$�w*'��+��0�υ9��  �  {�<xP�<��<�un<�,<���;Ý;@)�;?~�;*t�;2"<�Z<���<��<{��<�w�<��w<�!?<V�<���;�G+;+� ;%>;��;��<n�I<��<�E�<ɔ�<-_�<���<iK�<AA�<Z��<���<U��<��<�q�<Q��<�O�<���<���<�<��<�XD<��<��;h7�:�75��\z��ͷ9�B;���;�v <լN<��h<)�i<v�P< 5#<��;
lA;��	9d����������7k,6;$��;�&<wc<�t�<n��<��<⎶<��<�<��<�%�<Cӭ<ƥ<�ϛ<�q�<��<=�X<�J(<��;ɭ&;LZ����һ�`+�&�]�L�y���|���f��>���4���B��ch�5�����Q�5���z��'��-����ļ��ļ1��4��E���ES��>�,�໻���5d��04�T�$��`-�4(H���p��e��&m��~�ٻ=Q�fb$��K��}��<��~%��-�����X�T� �N������9N �����߼��߼���f����g+%��4��n?�D�.B��:��.��� ���p���2���켸`�,������@�漀���6�*����X�J�z��v�%.$�^�2�j�B�}�S�<yc��o�� w�Kx���r���g���Y��K���?��G9��9��2?�G�J��X��Ug���r�(]y��|y�2Os�F�g�<Y��6I���9��-,��>!�p��d���������]�w��Q��#�6g�^M��R�U�(�^D5�?%D�^�T�s\e��Ht�hd�-~�����~#}�smq��}c��BV���L��_H���J��]S��}`� �o���}�"�����������ف��Xw��Kh���X��I�Z{=��3�Z�,�(��#%�d�#�U#��Y#�!C$���%�h�(�k,�_2��:��  �  ��<���<�ˡ<��<2V<�l(<�i	<_�;��<c'<iS<��<
�<�ߤ<,�<��<�؍<�=j<_B5<�<��;_�;���;*�<[�2<�d<b��<_��<�ڵ<��<�Z�<�r�<���<|+�<��<N�<���</h�<;$�<dx�<���<���<
d�</�<%�Y<6e#<�,�;��;o�B;n/8;��;w��;�\<֋G<��o<�D�<��<�pq<�I<o�<~��;�Wt;^�;f�;{_;��;�"<u><��n<���<d1�<oA�<��<�>�<�N�<���<��<!R�<���<��<��<�Zu<+�P<��$<P��;�a;�ⱹK&��q���r$��D<���>���,���
�{�û��o��.
����//;��g���r�rK�䂼q��/���^���C��]#����n���@����O��^��­��,c�s�P��zS��bh�b���须�jĻ�n��f�ܝ.�1�R�7O~�Ռ��7��Ӽ-�E���^��P����I�	�~[ ��켪�ڼ�м��ѼFv޼[7��ME	�v��Ȓ&�p0�\
5�|4��Z.��/%��V�u����0��s,�A�<��M"���}	�𼮷��B����D��
��ױ��$��00��=��xK�@X�6Rb�&h�v�h���c�ZeZ��>N���A�{�7��1�[�1��7�aA��M�}Z�33d���i�*bj�܊e��f\��{P��|C���6���+�*�"�b���L�z���'�����S���U� ��P��'���!���)��^4�ʰ@��DN��[�-h�C>q�8�u�$�t���n�ϐd�Z�X�M�p�D�;A��DC���J�TV���c��o�1:y��}�G�|��v���l���`���S�&�G���=���5��d/���*�]�'�u&�6%�ZK%�S&�8M(�xB+��Z/���4�0	<��  �  ���<lG�<q"�<��<���<G�`<VK<��D<�(O<7�h<br�<�@�<ᡫ<Mض<@]�<�m�<�9�<���<�p<��I<:�.<#�#<W�(<1�<<FhZ<@}<[�<Pܠ</Y�<#��<;��<G?�<E��<cl�<r��<|l�<�g�<���<P`�<���<ྶ<���<�P�<�߈<:�k<��D<�n <5H<���;@p�;�K<l�%<�GM<��u<�h�<	Ɣ<���<u��<�v<)�M<��#<��<�;4��;D^�;{�<gc.<�Q<rCt<N�<�ە<���<���<�׫<�8�<w�<ç�<7�</��<���<M��<"|a<�><K.<���;AH�;$�:P�ߺ)����Ȼf�뻭��ֱл�p��~z6��]���/.9���9]$:�jF9�.��"^��E��m� ����l��oՁ��8n�:�Q���2�0��"����л���:;�����%ى�쇏��=��jj��G��	��C$�ՅB�C�c�pW������HZ��T�ļ"Uڼ���V����#��~���˼�Y�㼋�Ӽe:Ƽc5������̼7t�����5
��.�j�]�#�I_$�;7!��x�p��H�l�������#���K��~�'��g������4�����>	�Yj�a<�����(&��h/��K9�	AC�WL�?\S��(W�s�V���R��J��@� I6���-��()�/�(�x-���5��@��|J�[S��)X�q6Y��BV�8P���G�¦>�d�5�%�-��w&� ������lw��q�ݥ�X8��#�>��]�=k ��g&��i-�|�5�Q�>�9�H��gR��[�Zpa��Ld��c�t�]��hU�X�K��'B�3O;��{8��_:�G�@��NJ�vZU��_�\�g�M�k�"�k��.h��~a�!Y��FP���G��N@�'�9�\�4�M(0���,��(*�ػ(�4�(���)��P,���/�H�4�:��~@��  �  8��<�<�7�<���<�(�<���<��<`�<E��<���<��<�W�<ɴ�<�5�<#��<?�<��<���<��<^��<<>u<Q�g<Z4e<�l<#�y<�]�<2��<��<ڪ�<6V�<' �<	��<�G�</��<'��<r��<��<�X�<���<���<3�<zz�<�<҃<:Rq<]�[<��H<�];<�6<P;<o�K<A�e<���<6��<�h�<���<*Ŧ<���<"��<�b�<Npc<%G<��3<��+<��-<%}8<�6H<�.Z<7kl<�~<�u�<߀�<�<y�<,�<���<�s�<��<�2�<�+�<n�c<ɆA<B�<�y�;H�;�ft;���:�9�w��7�!���E�D�>�CR��Jx�l]�9ɾ�:�>#;�! ;���:8�����6�}����Ǫ(��pA��PN��XP� J�5�>�1U1��?#�pH�Z������-~ۻ;�ƻ!����v���>ƻZF仾t�2$�tC�ac��V������t���ڭ�ι��Y�ȼ�Ӽ`)ڼ=qܼ�oټ-�ѼʇƼWк�Xy��^E�����Dh��FE˼Th�.����������0�F��������nO��Y��d�]��u���&� �%^������ȏ��� �t���-
� �����Ү�Xj%���+�2���7��y=�UCB���E�m�F�]sE��7A��:���2��w*�d�#��; �� �5�#�j*�I2�4�:���A�F��H��%H��|E��rA��<��7��2�<�-���(���#�S������'���>��������#���(�J�.��t4��=:�E @���E�)K�ȪO�k�R�zlS�asQ���L�f�E�L<>�F 7�\�1��/��I1��\6�|>���F�q]O��6V�ًZ�\��#[��GX�tGT���O��!K��sF�j�A�?�<�T38���3��90���-�-�K�.�F2��6�u<��pB��rH��  �  @x�<*У<���<��<�՛<) �<���<�Y�<uy�<+2�<���<�2�<���< ��<��<�g�<��<�h�<�]�<Tۤ<�T�<��<Xa�<H��<h�<'��<�$�<��<|��<nb�<}��<�q�<N�<g��<v�<!O�<�/�<<t�<���<��<$�<C�<�v<m�k<i�e<D�b<ZYb<��d<	�k<��w<!��<.��<�(�<�#�<��<���<���</��<��<.y�<S�<j>�<��p<�b<��Y<DT<4�Q<Q<�R<�>X<W�a<I�o<D��<�ω<�y�<���<��<�:�<�ށ<y/b<3�;<�q<���;䎣;��f;�;3W�:�ă:r: M�9V��9�.e:G��:�";Db;&׊;Y�;���;z}c;� �:ѐ͸�;�Qj��K.ػ`%������*���5���<��rA��B�	O?��7�x*����.�	�P����ﻋ������i'�u�H�X�m�t���B����]�����/����1������������������������0����������X���;婼q��ttɼ�!ܼ������&?�2
����l�Kt�U��3V�?���������d����O��>��U����������#�U�*�M1���5�-9�S�:���;�T�;��G;���9��i6���1�9,,�*�%��� ��^�j	����ǉ�;�%��a,�8y2��n7��;�hZ=�ڦ>�`6?��'?�Y>��<��[9�~�4��>/��&)��|#��>��A�����\!���&��-��e4�F�:���?�	MC���E��G��G���G��$G��NE��$B�ɟ=��8��&2���,�f)���'�$)�+�,���2�_�9�g�@���F�ڹK��AO�ƏQ���R�B�S�"�S���R���P� �M�[�H�9CC��o=�Y\8�b 5��4���5�AB:�qh@�ikG�:QN�2ST��  �  rJ�<�
�<���< ړ< �<n'�<gt�<"ҷ<J�<{��<bT�<F��<���<F��<��<!��<�}�<���< ��<ü<9ڰ<��<�i�<#Ӎ<���<�p<f"a<�NY<(�[<T9i<D^�<�Y�<�ٞ<�Ϋ<���<f?�<$��<��<wU�<'�}<8E_<(iI<,~><v><1vG<<�V<�i<��|<�F�<X�<���<��<��<�ݹ<��<tg�<�U�<mo�<�R�<���<D`�<y]�< b�<�|�<�,s<�[]<f-H<�a5<ï'<=�!<��%<V�3<��I<9c<djz<'��<n��<*c}<X�`<B8<	�	<�޷;�7Q;�S�:}�9x�Y��39�W::�:�Y;��C;|�v;�u�;�Y�;]��;^��;�2�;z��;mh�;��w;ݥ	;��W9�R�C�t������������
�3�P�M���c��Js��Xy��t�[>f�}P�ut8�($��N���
�-�:7M�Ov��*������/���s¼s\Ǽ�Ǽ��ü�ｼ6$��Z2��D`��»��N��xe��/���Z��[���y����`���M��xö���Ƽ��ּb�漐������l`
����,H�����!�P�"��x!�n��f���?��)�
��!������$��'��81�	:��t@���C�]mD���B�e�>��Z:��i5��T0�++�A�%�[� �jp�H��-U��d�v_��K����N��`� �u&��,��1�Q7�|<�h�A��;F��UI��GJ�̐H��D�\n=���5�"�-�r$(��R%�(&���*���1�WY:�]�B�o�I���N�Q�P��O��4M��AI�ָD�E@��B;��z6���1�X�,�9D(��u$�b�!�:!��,"��&%�ݘ)�r /���4���:���@�E�F�ˇL�KR�"�W�"\�g�^��F_�!�\�w�W���P��0I�=?B��=��<�wW>��C���K�F�T�:8]���c��  �  �U<�+X<�{i<�ӂ<oܓ<��<�&�<���<�L�<8��<�*�<���</��<J�<���<�<6��<L6�<���<���<kf�<n�<���<�\�<C�p<��J<i7,<�_<�<�[#<�u?<`+e<I|�<@L�<wn�<L��<r�<Vb�<�k<g�?<O�<"�<&��;�<�<�X:<�u^<�N�<���<3��<��<���</4�<��<��<�n�<.M�<�~�<�M�<M�<���<��<d�<@�<;){<� U<�Q.<�
<G\�;QG�;:��;f�;��<��-<��M<`�c<f3i<�
[<��9<��	<��;�d�:QX���6��h�cV���T�;��:d�>;V)�;3��;�k�;�G�;���;g��;���;���;�I�;�#�;�5t;��;��j97 �<v����ԻU��c�B�j�n�/_��*E��
��M����˔�/c��j�k�P O�<'>�Zi>�x�Q���v��ғ��W����Ƽ�]ټ��㼩��_༯�ԼQ�ż*���4X��E������%���𳆼��͛����������0a��5����
��$��U�Ƽ�ؼS+�} �IZ�%��[�!�
:+�>�1��c4� 3��D.�('���������v�M��{�(�:�4���@��4K�X R���T��S�?�M��F�P=��3���+��$�x���K����D�%���d��g�����a�����u'�\�$��[,��5�}�>�mJH��Q�Y�W���Z��&Z�HRU��*M�]6C�Ir9���1�i,.�/���4���=��}H��S��`[�'`���`�}]��W�w�N���E��H=��5���.��B)�~�$��� �9�����!����Y�@�"��,'��,�M�2��:�ozB�5�K���U��_�`2h�n��_p���n��h���_�vV��M�y�F�X�D�x�G���N���X�b�c�G�m��Iu��  �  <<c�<��1<�U[<�R�<X��<c�<έ�<�X�<�<+~�<�!�<���<���<k��< 2�<7��<h��<=�<���<`��<��<��<xʄ<�4R<]p<f��;v��;{ �;���;��;��,<�\]<�@�<z��<�^�<u��<��h<Ԛ6<��<�
�;��o;hW;��;���;�<�H<�}{<Q��<`��<	ƶ<X�<�C�<���<y�<�'�<V��<���<"�<��<e��<I��<۵�<�K�<��u<�AA<a	<%�;{H;�A�:�3�:P1;��;˴�;��!<O�><�G<�=9<��<'>�;D2�:���뢨�4��R����v������&�NG9�J6;w��;)7�;�� <ic<S<F�<J�<)W<m��;�v�;���;�2W;�ǿ:j;��1Y���лP� ��\�Vዼs����¸�hO¼�1��&������|���!y�`?b�7*`�Yu��Ǐ��$��3	˼�@�0��i�s�ފ��:c��.ӼDQ��3|���_������8���y�K�u���w�3L~�Vs��񾋼�씼I ��;������м����� ��S�<��1s-�c�9���B��DF��D���>�4a5�+�+�N�#����|5!��(�؜3�B�A��+P��=\�o�c��*f���b�
�Z�bO�7�B���5�n4*�Z� ����8��h����	�x	�W	�
�R	�J��[�t8�A� ��*�7�6���C��4Q�#�]�}g�H#l�6�k��pf���\�БP�M�D�o;���6���7��|>�WI��VV���b��l���q���q�~Xl�~�b�L�V��J���=�	W3�P�*�;/$�Oh����s��r����eq��1�%"��B'��.���6�(�A��vN��>\���i�7�u��@~��������]y���n���b�-�W��P��rM���P���X���d��Mr��^~�;v���  �  �;�׸;^��;/�2<�o<�<S˳<6��<�\�<��<]�<���<�C�<��<�i�<bi�<9��<�c�<��<��<�f�<N�<�̚<=�u<��2<S�;�Et;���:�^�:0;#P�;�;�5<��d<Mƀ<̂< �o<��C<V=
<��;���:�ĸ����Q:�m\;�;͢/<jKn<�<a�<�n�<5��<��<*�<���<�#�<���<�b�<�7�<0��<}d�<��<�_�<@S�<?j<��)<�N�;ކ*;nw��g�����(Z����:�ԙ;���;+j<�+<F�<���;��X;6}���խ���H�0��
8�a|%�*����3���Z���L;*��;<��;~g<xC<.�<��<v&<j�	<{��;<h�;�`�;$�;��
;[pl�0�N�L�ۻ=�0�X�x��П�G徼b�ռ��A�߼��Ҽ����V���Q��Ub��0�|�n����	��'����f�Ł��~��y��h
�ǚ��e�ἆ�ļ�����2������w�8m��9k���n���v��݀�߇��b��7Ț�����g-����̼4������Y���&��]8��<G��{Q�G�U���S��OL�hA���5��I,�!b'��(��#0��<���L�q.]���j�Xs��lu���p�Z�f���X��H��9�^�*�te����+/�����<	�,��.������u	��-�*w��������D+�׀9�'�I��Z�@i�y�t�?I{�V{�u���i�)�[��%N��~C�=(>�YP?���F�C4S�tb��zp�o�{������V��M�y���m�b*_� ZO��X@�f3�K#)��!��z��G�7�����m�����3�i~���Vv$�[�+��%6�"C�	dR�"'c���s��$��2T�� ���+����Ƀ��]{� fm��`���W� �T��>X�P�a�/uo�p�~�6�����  �  ��;�P;���;�<*�Y<��<�3�<u�<۔�<_��<��<bE�<X��<��<MU�<~��<xS�<��<���<a?�<�B�<!��<y�<�f<��<�>�;��:�a_��Rƺ�WṠ�;9�;�<H�M<S�m<2r< HZ<��*<���;]�/;(�"�*-�0aC���Ϻ�P�:�;J<�b<s��<��<@�<?[�<���<��<�7�<��<���<���<���<���<� �<Ÿ�<[��<�$�<�5_<��<�<�;��:�-��_��OQ���4S��E�rE<;��;�f
<C�<`_	<�~�;�,�:��@�g�����6�AzZ�;�`��J������Ļ��I��:l��;���;6�<��<<"<y�<�T<3�<� <w>�;x�;	��;�;&,��f�S���\>�����;���м�������i����弭�ͼI����7�������懼$���P���̖μ���@�
�"H������Q� ��m켴�˼b�������x��Z�r�/h��f��[j�B�r�D~����E-���L��&I��e?���M̼[I����d��,��+@�9�P��[�W`���]�_�U�,wI��<��2��o,��-���5��AC�diT��e��t���}�����z��5o��m_���M��<��H,�7g������� �
����=����$�<���/��
��,����ɇ��b,��><�)4N�ѭ`�̏q�v�~��؂��悽
�~�&�r�@tc���T�d�H��C��ED��cL���Y���i�Ȕy�J؂�
����|��A���x�u��Ke��S��B�j44���(�ԕ ��%����%K������ܢ�l���,����xB#�VN+�^d6���D�e�U�?lh���z������Q��z卽`䌽���m恽t��f���\�~�Y��Z]�w�g�hzv��y�����/���  �  lH�<���<���<��<X5�<���<0�=��=	K='�=�<=Q�=B�=N=�v=��=|=��=�#=��=f=|=t�<���<��<�޳<j��<���<8ő<���<\�<��<}��<?�<C�<��<���<���<ݵ<��<�W�<��<G,�<�Ջ<�Й<��<a��<'G�<�:�<�]�<�# =v,=7�=2@=`L=M)=��=^�=�C=a^=��=�r�< �<C�<���<��<�E�<�1�<�|<��h<��d<��p<ҫ�<?�<JA�<���<r9�<¡�<Jv�<_��<�R<� !<�(�;�;�.�;��;8��;��<��:<��Z<u<�k�<��<f��<O"�<�ׁ<�y<ٝm<�a<~YU<|-H<q�8<S�%<��<},�;Iч;� �:���0F��^Y�������/�E(1���"�_	���׻�u��Ԇ��f��{����D�E�$���U�B_���,��$暼����o���(��pe�E�A��}"��`
�&L���=����q�����r��u0��"'�i�3��'A��{Q��f�"�������1��������ڼ���¸��h���,��v��^,���������3�W𼒤��������)?���&���,��|.��+��%����t���S�׫��m�4Z�}޼��ڼ�ټ/Tټ�xټ2�ټ�=ڼ�ۼ��ܼ&��U9缼���; �Z�	��Z�͈���)���1��]6�9�6�ɵ2�>t+��n"�;��������8m��r�ů�'�'�4=1���8��<�L5<�)�7���/��&� �����s�	����K������u9���3�����������+�������f��J?�����4�������H,!�
�,�.�7�B�A��I�W�L��K���F�V�>���5��-��3(��s&��(��[/���8��B�n�K��R��  �  ��<��<*��<�K�<m��<Q�<�=�/=MU=��=�!=�=m=L�=h==�==��=�	=��=�(=�b=AB�<<��<:��<;;�<|�<�ۙ<7$�<�ɚ<^��<M,�<���<a\�<��<\�<h��<$s�<�޸<��<�^�<6j�<���<E��<�t�<���<���<���<��<O��<�" ==ޘ=I(=�9=�=L�=ޟ=&,=�B=�o=<g�<oC�<�<���<!��<%#�<���<g|�<zjq<�{m<r�x<�8�<H�<��<�<}�<Ɇ�<Q��<�*�<��X<{[(<� <���;C�;4��;v6�;D'<+\><�C]<5v<���<Ƈ<�D�<��<ϧ�<��x<�im<�|a<� U<��G<�8<�}%<��<�,�;S��;+��:�ĺo�����3�8	'��(�f��u��1̻�ޚ��<}����������0|�.JO�1){�z���������J������f�`���>��� �D�	�Q��u�黭����������P�:C'�(�3�vbA���Q�\f�rĀ������림�Ⱦ��ؼ?r𼍵��8
����%��y�	�����������#��U��w����ju�4u��$�1�*��L,�6�)�TK#�l��k��������[�
F޼�ۼ��ټ�xټ�ټ�ټ�aڼ�Aۼ�ݼ���mB�go����u���I����(��/��04� w4�Ӭ0���)� � �Q�=��]���m�T�:[���%�*`/���6��k:�::�L�5�-#.�?�$�q���S��v	�f���_��U���n���_��+�����WK��Я��g���pZ����y.�SL�?s��Z ��R+�BM6���?��G�ORJ� tI�T�D��!=�+q4���,��)'��y%�'�'�{-.��7��A�J�|`P��  �  ���<���<u�<��<�L�<L^ =�;=N�=W6=� =a�=w,=�=��=F1=�=�=br=�=�=�"=�=^�<"��<T��<�x�<-r�<�<8u�<ś�<	^�<�`�<h[�<b��<j��<��<���<���<�b�<��<7��<뙗<�ʕ<�}�<_��<�̷<?��<�y�<��<��<>��<J�==��=R�=��=۬=nV=c�=M�=�� =��<��<���<�V�<��<a�<z��<~ȍ<?΄<nւ<]Ӈ<D�<�c�<���<��<�m�<��<��<�m�<Pj<a�<<x�<L"�;U��;KQ�;�#<&�+<�RH<�c<�x<�|�<M��<Y=�<��<��<��w<��l<��`<�T<�{F<��6<�$<�t<��;���;�;lF7��:_�������H9��=�7����ݻ���������N�0*V��퍻u ͻ/���<��e��?������ 늼=@����p���S�Y6��������>���)�nvﻦ����-�m�����{�'�O�4�зB�#S��vg����隐��ܣ�'�����м�缽K��^!�S����05�N�����	��T�^��^T���*��f����;�$�;'&���#�p>�]�x�J������۩����`*߼;ܼ?�ڼ�ڼ�ڼ�TڼF�ڼ@ܼ�޼���`���#�/
���%��x�*�-#��*�7.�IY.�V�*�7�$�����������֙�(�Ė��{!��*���0�yE4���3�k0��h)�� !�q���3�����c �����W��������Ŋ��G���+P���6 ����Wi��X�s���U�KC��"(�U2��:�� A�[*D�kC�?"?�E8�"Z0��")��7$��"�%���*��3�c=<���D�baJ��  �  ��<���<��<�7�<���<F�=�P	=�~=(S=��=�_=�=�J=�!=��=��=c�=vO=�C=,a=+b
=�= ��<r��<m�<�P�<|�<�Y�<���<��<6�<��<{��<�a�<�@�<F��<M��<S�<�	�<���<���<و�<欧<W�<���<��<�a�<��<)/�<ID�<	��<iW= �=��=13= P=�=��=��=��=�L�<���<s�<���<��<%��< l�<�>�<s��<Zj�<7��<L��<�#�<���<�$�<l��<}J�<�߶<x��<P4�<%(�<Y[<�t9<L�"<��<�X<�*<F�><�T<#�h<#(y<9��<���<1��<���<�0~<�<u<��j<��^<�EQ<�B<e\2<#�<*	<!��;_�;n�-;���9���޺���1����ӻP�ػ�ƻD���Kv�us/�eH
�9�&�X��W��p9��� ��E���a���q�t�+�j�=Y�.�B���+�X��}��)����#���r��Й�/	����v��)�5�7�*�F�}�W���k����L��ᾠ�zi����Ƽ!�ټGl�O������qi��v`��n��t�NM߼��ܼYP�p=��i�����a��������.����� ����g�	�_��@���Ey����̺ἃr޼l�ܼ�~ۼ@#ۼ�jۼTWܼ��ݼ�n�&D�J�p(���?������0��!��.%��Z%�[k"�,��X��S��
�˜�8k��t������{K"�N (��>+��4+�o,(�!�"�c�%��J<�(���6�C2�1�������x���A���s�������A���TD���ӭ�!K	�u+�Wg�@��r�#��#,��Z3��8��);�v�:�W�6��1��F*��$����=���� ���%��"-��&5�[d<���A��  �  ���<�2�<���<���<� =��=�<	==�=�=�2=�=��=�=
�=��=Z�=�=�=,�=��=�'='�=i��<��<'�<��<8�<��< E�<EX�<���<n�<R1�<���<<�<yX�<f,�<=i�<���<"�<=�<B�<=�<���<Q��<���<���<���<8��<��<y��<S�<�v =�=��=� =�=k/=�� =JT�<���<�b�<�s�<K��<���<҂�<]��<�θ<��<`�<��<��<��<���<_L�<��<�_�<��<
�<�ͣ<�b�<x�~<\�`<̖K<y�@<χ?<��E<�/Q<*&^<$ij<�Gt<S�z<}~<AG~<��{<��v<��o<�Kf<q	Z<_fK<��:<��(<�f<= <_�;7!�;��I;b��:��m��k�R�����*��3�s��A����d���lj��g��� �Nur�;˺��` �W| ���9��I��XN���J��@��3�
�$��`�������Y@����i�	�--�����R!��S.�}�=�3�N�a�L-u�߲��)�������m������5̼}�ؼ��O輣�輱��+�߼��ؼ#�ӼE�Ҽ�ּ~�߼��켳���Z�֨���>���J�Y���I��b�Zq������(�I��k��F�ci�{o޼�{ݼ��ݼ�2߼_��q/�5��%���1����O���	���Q���������V��d���@	�K�����3��*��m���S%�D�	� �<D!��n�����L��d�%��M�	��\�>��"��)� �v����������?/ ����U�5���\�.�����ݪ��:��6 �p#&��Z+�j$/�C�0�{:0�&G-��(��##�7&�J��2������ �j%&���,�\�2�H7��  �  ��<�F�<�~�<�Q =�o=��= =�T	=Q�=��=�=P~=��=�=�}=@G=�+=�n==Y
=�=z�=v =+�<��<!�<���<T��<���<���<���<�x�<Q[�<]��<��<�� =6� =P��<���<���<��<M��<���<���<"��<� �<m�<Q�<�N�<�~�<���<�x�<NP�<���<�+�<J1 =E=�� =�n�<��<��<���<�#�<,�<�<ԓ�<h��<yL�<�0�<�S�<y�<.1�<(��<x�<��<x�<r��<�G�<�<v�<Bn�<ü�<�Y�<<��<�Ds<��e<:a^<�I\<\�]<�e`<Y�c<4�f<Oi<E?k<Bzl<�l<Wk<��f<�V^<��Q<�AA<b�-<�<3�<��;PX�;Ë;֋G;  �:9n?:6߇�d��t�º��Ϻ�����:`�����C9q��9��V��x�!g�����B&��5�������!��+�iW.��`-���)�H�%��M!�O�����f���H�)[�q�����(���6�lH��\��q��:��wύ�gF��������-4������b4ɼJ�ϼkuӼ�[Լ��Ҽ�ϼ0˼b|ȼ��ȼ)�̼�
ռ_Z��h�\��3������	�/�	�e��r�.���8��?��������	��2���+v�e�Ἦ�Ἵ伭��M�켇��R��*F���2�G\�f��%�����ۇ�Ba� ��̒������W��1���&��,~���z�-����
����a��y������~�m�
�����;������
�Up�<R��X�������}��X�+�D����	�`��9������e�����q!��O$�~C&�[�&��&�%�#� ���
4���<+���<�;��g$��M)�'-��  �  �U=XT=��=^�=�_=6 =W=�)=�=_�=��	=c�=�=�b=�d=C�=��=�>=�0=V[ =�.�<v�<^e�<B��<)6�<�?�<��<���<���<N�<Y(�<&��<�d=
�=G=��=7U=�h =�g�<E��<]a�<�e�<���<9��<<��<��<)�<��<��<S��<���<|T�<���<���<u��<B��<�k�<*�<z�<d�<��<�h�<:��<)��<�#�<�B�<���<u%�<���<)&�<�n�<J��<���<���<�/�<h��<���<���<�q�<.��<�g�<\:�<�<Ky�<ѭ�<�u<�i<6`<ZX<��R<E�N<pN<p�O<�S<�7W<a�Y<f�X<�'R<�'E<fI2<_:<�b<CT�;���;���;�K;�;ſ�:^�:�:�-::9c:Q�:�,F:3c�:UJ�:N�:���:+Dm:���8x�����&�z��������3޻�� ���Sf��n#�"�*�2�0���4�P�6�Z�5��*3���.���*�}�(�n�+��-4�#+C���W�،o�)?��2������녣��Ȫ�=���ȫ��>鹼�z���7�������S¼���9-��'����e�����F�ļ*�˼l,ռ��߼�^��������� �i�+{��Q����Ж��������V�R����u������Q輍(�cV������W�����������	���	��G
��h
��'
��a	����M��g������������ ��j#���S��H����������%���!������.�nw��W�����M��:����	�L�� !�]�����l�R���������
����p���o�Aq����d�hC���L"����V�dy�����W��If����������� ��4$��  �  �q=r�	=m=��=$�<"��<z�<P�<���<`��<c1=�L=^�	=�=�R=�o
=]�=,�=���<3v�<�o�<8x�<���<�L�<���<�D�<��<���<6y�<���<�*=�E=�+=��=�V==~�=�=�=�,�<���<U��<�J�<*��<��<��</��<m�<Q�<T%�<R$�<|��<߁�<�H�<?l�<X�<q&�<���<��<�t�<@��<���<@U�<w��<�v�<q(�<,�<Z��<m	�<c��<v<�<_��<��<�R�<F��<��<���<���<�J�<�B�<�-�<鬭<e&�<Ȗ<��<���<��k<y�W<J}E<��6<��-<��)<U,<�E3<R<<+D<]�F<B<S�4<��<ly<vc�;�ɒ;�F;�-;���:w!�:vώ:���:���:�=�:��;��;&�;	?$;��%;��;�
;���:��Z:��E��ĳ�x�,��A��ξ��ŀһ2��� �\l$�T�6��;F��R���X���Y���T���L��WC��<��<�[�C�w�S�a�k�Z2����%���1���h������Mƹ�c����{�����"ѵ�:촼hc��`,��pL����|��l�����4�ļnU̼��Լd�ݼ*0��j�MY��%��:��*D��S	�r�� ��x4�N%
�e��(M�����]��P��e𼍭���Z��������i��v� ���D�����=	��c���s]������Z��� ��>�������� ��~���#��l#�hP������
�:L������=��J
�t���'���o��O�'i�e�	������	��(�����<�����s"��j#�E�"�)�!�uz��)��������b�(E�C:��X�Y������v������_��B��k��  �  ==�=�Y=�S =���<\��<���<-�<�I�<t��<K��<���<�=$=7�=M[=
� =���<j��<��<���<+��<� �<s�<@��<}I�<���<w��<��=e=�=I[=�	=�>
=�{
=E%
=�5	=F�=��= {=�� =A%�<1��<h��<�Y�<���<|��<8W�<\C�<ҿ�<��<H��<m��<�,�<���<Y��<���<��<�3�<>��<[��<m��<�α<��<�ֳ<u��<)��<��<E�<��<�-�<��<w{�<	��<8�<mo�<� �<p7�<���<5�<���<�,�<
��<�0�<k�<j��<,1d<�E<*<p�<�<-~ <(�<��<~R<�i+<9M2<@x/<�f!<?�<o�;�;`�;Ԋ:��h���D�ćF�6�!:�@�:��;*�>;f1Z;~�g;�xh;�^;��K;��/;��;�8�:u��9v��ڦغ�B:�T뇻Q���뻜��7/��kK��.d��v�i����*��" {�,�m�H�^��.S��O��}U��-g�LS��r0��Y£�\��������Ƽɼ�%Ǽ�O¼|���ܵ����/������Ԫ�嫼��� ���괼D˹�ϛ��m%Ƽ2ͼ�Լ	�ܼ��弒���#�������	��2���&��`��(�q���0
��^��8������U���X��=����
����������K=���2��OH��+
�89�`� ��q�������x�TK�a���鼍�鼨��׻켁�����h<��v������>�����v�T[�b���"���$�2c$���!�7�N�����*���b�a��
��	���#�Y%��*�@�,��,��*���&�S"�~�����@�?������\��n�����o�����N�_=�����m���  �  .z=�=�g=�[�<J5�<�F�<���<�~�<:��<���</�<���<]��<�(=t�=? =�a�<�r�<���<w��<Z�<��<�%�<5��<G��<���<���<�t�<D={�=g	=��
=��=�=k�=�I=J�
=$�	=F$=�=R8=DZ�<à�<O�<q�<���<3�<���<�J�<���<���<�f�<��<�+�<���<��<���<�]�<r�<<4��<�ƣ<\��<�V�<���<��<~�<��<3�<��<���<~��<�q�<���<$��<���<v��<��<}S�<Ư�<��<��<CU�<�f�<��<l^}<��U<ق.<t�
<Z#�;EC�;7�;�0�;Ʉ�;`� <��<��<M�<-<=a�;>=�;��;�������"LA���T�-�6�)"�cY��:m;q�T;��~;<�;Rʈ;���;\f;��B;{1;jm�:�XT:x9�����h�sm�����W�컰V��<@�}6e��Ђ������W��<����[���I��H7z�a�i�ab�t�g���z�Ҍ�����O���^ƼK�Ӽ?�ڼ7�ۼ��ּ��ͼ�ü���ய��`��M����C��������������P���U������0`¼hsȼyOϼ~׼��Ἀ���C��W0�l|��4��b�O �|� �.��������
���=��e������
��Z�P��g���#�dN#�� ��;��m����������k��p�Ｍ'뼒���R���漌8缊'���D��:���z�����������&�����[&��+�9�.�ļ.�s�+���%�����3��>&�ҧ��N�~F��='���.�N:4���6�$x6��3�"�-�ڸ&� ���2������c ��Z���
��G
��f
���
�W�����\���3��&���  �  w�=�
=��=ex�<���<�
�<�I�<�q�<�1�<n��<~"�<� �<>��<���<c��<��<8)�<,�<���<�<Ն�<,�<�A�<� �<�Z�<���<*K�<���<K�=�=W�
=�=+�=��=LD=��=�>=xy
=�P	=Hk=�_=[��< �<��<�x�<z�<��<���<ɤ�<�<��<�<G˲<�<Q�<ȴ�<հ�<.�<���<���<rf�<F��<v�<S��<c�<�!�<�~�<w��<�`�<���<��<���<���<� �<+�<���<��<���<2q�<�W�<0�<�T�<��<_١<�f�<32t<~�E<��<X��;��;��_;��I;�2m;p�;��;V�;��<�Z<l��;~a�;'�];K�(:j���h������� ��
����*X��@˺��9���:uT;�Ʌ;SÒ;`�;�b�;\�r;w�K;F ;���:��:G�-9�M�s, �,,a�-b��+�����%�BLR��~�.$��v-���k��YB��-y��s=��������|�s�܋w��҅��������Av¼�ּd*��y��켘��r
ټ��ʼ����:��:���X⣼t���O��׈��������#���A��o��� Ƽ`�̼*ռG+�P��w��Ul	��y���_$���(���)���&��� �U���d�ٳ	����G���	��^�t��,e!�~=(��,��.,���(��"������5��2j ��P���\�'�輦0�sn�׎�@#�I�A�o����aM�as���n�}m�s	������$���-��K4���7��7�V�3��J-��_%�\���l��@�����"�3%��#.���6��<���?��)?���:���3�t\+���"�����V��3���
��i	��l	���	�OO
�`�
�a�������������  �  A=�	=��<5��<���<�S�<�a�<�<�=�<��<j��<��<�D�<��<��<2��<?F�<���<J-�<��<Em�<�Ν<w��<���<��<ڢ�<�9�<���<u9=�=�=͓=�=J�=�=0
=E�=	�
=T�	=a�=��=���<��<��<�5�<�p�<��<�y�<́�<��< �<m�<�ة<ʟ�<[�<��<=�<���<�>�<��<��<��<�3}<��|<���<I�<Z��<`_�<P��<�B�< j�<	�<��<���<��<=1�<p��<,�<��<P��<���<��<�X�<�1�<�M�<G;l<�9<��<^ͱ;ZS;��:�z�:��;�k;�.�; ��;���;�Y<���;<��;@S ;�u���T�ʗ�� �ػ��޻(�û�J����Q���q�:��K;�+�;K��;|��;.��;X�w;��N;8�";P��:Ў�:mx�9dE3�{�����`�s����� ���.���_������䜼P�������0���W������咐�����zD~�� ��苋��W������̼�|���o���ݑ��$）W��Ѽ:��dF���:��cp��𣡼��������^���~��J�������񢿼ż�˼'fԼ�;����I����1��!�/�)���.���/�J�,�{�%��/�;��q��|��б���$A�Ћ&�).�#12�>G2�.K.���&�>���L���	�4�H����켋���A�J���;��`����r1���_i�C ��G��0f	����ø�T�(���2�A:�5>���=���9��G2��)�6a!��m�h���d ���(���2�l<���B�!F�)E��G@�Ri8���.�3�$����Lf����2i�v�	����E	���	��
��
�΀�'��lK�]/����  �  ��=�	=�<]6�<��<(x�<�!�<���<\�<��<S�<JE�<���<���<8�<���<���<��<쵺<N�<�#�<9o�<)^�<��<�м<!K�<Q��<��<K=l=�/=�==��=�==��=M�
=�	=N�=ʻ=�L�<2��<���<�3�<U��<D{�<�u�<�.�<iH�<��<۹�<5��<3��<���<��<��<S��<֨�<<��<9l�<�<�|t<��s<$�<ⷐ<ˣ<->�<Iw�<�|�<�<N�<��<���<���<MD�<���<^'�<���<��<`�<z'�< N�<�Ѡ<�k�<�(i<�+5<�� <��;�2;��:Ua�:��:jDO;I�;u�;�r�;���;���;��;��
;9�d�{[r��O���E�
��s{ӻٙ��r�1�i\	����:T�F;B��;��;-Z�;!d�;^�x;u�O;�v#;���:��:��9+�-�B2���a�6������@F2���d�;�������T������c���*��B&S���D�����m��ǒ��B����ݶ�rmϼ|b�!D���������M��j��mӼ��¼�2��D����x��i{��Oբ��o���5��9\��������>r����ļei˼)PԼtm�TO���0�|���X#���+�1�p2�.�.�e�'����n���Ϳ	�L�	�Q��<P�����](��0�/]4��r4�&S0�ϼ(����?X��<
�H������ǹ켏p��弍�a��9�弫u�x��\鼒��5>�)��9����	��������4*�s4�*<��/@��?�$�;��
4��+���"�m}�I����H�!��M*�Pm4���=��E��PH��LG��<B��:��'0���%��s�Ȭ����[�.{	����1 	�v	��	
���
�Ol��v��0�������  �  A=�	=��<5��<���<�S�<�a�<�<�=�<��<j��<��<�D�<��<��<2��<?F�<���<J-�<��<Em�<�Ν<w��<���<��<ڢ�<�9�<���<u9=�=�=͓=�=J�=�=0
=E�=	�
=T�	=a�=��=���<��<��<�5�<�p�<��<�y�<ʁ�<��<��<m�<}ة<�<Q�<��<-�<���<�>�<���<��<��<|3}<��|<0��<�H�<۫�<�^�<���<�B�<j�<�	�< ��<���<V��<�5�<���<!�<���<��<���<w�<^j�<E�<0b�<Sfl<��9<!<$�;� T;�2�:}��:(u;��k;X�;y�;N��;r[<���;w��;� ;Re���T��ڰ�&"ٻ6�޻�-Ļ����%���d��1&�:��J;W�;t�;�s�;ۍ�;Ύw;�N;��";ɯ�:��:��9�1������`�c6��ѓ ��.���_��燼~Μ�:��e������pH�����-������>~�!�������^�����̼Č�2�ɤ��ǧ��!.�o�j0Ѽq���\���O��ۃ������k������yj��k���0���׬��৿��	żԡ˼hԼ�<���"J����1�!�!�F�)���.���/�U�,���%��4�>��s��~��ѱ���%A�Ћ&�*.�$12�>G2�.K.���&�>���L���	�4�H����켋���A�J���;��`����r1���_i�C ��G��0f	����ø�T�(���2�A:�5>���=���9��G2��)�6a!��m�h���d ���(���2�l<���B�!F�)E��G@�Ri8���.�3�$����Lf����2i�v�	����E	���	��
��
�΀�'��lK�]/����  �  w�=�
=��=ex�<���<�
�<�I�<�q�<�1�<n��<~"�<� �<>��<���<c��<��<8)�<,�<���<�<Ն�<,�<�A�<� �<�Z�<���<*K�<���<K�=�=W�
=�=+�=��=LD=��=�>=wy
=�P	=Hk=�_=[��<�<��<�x�<x�<��<���<Ĥ�<z�<���<��<<˲<�<�P�<���<���<�-�<d��<d��<"f�<䣒<��<���<fb�<� �<�}�<m��<�_�<���<���<s��<��<��<�"�<���<��<��<!��<�n�<�J�<us�<�5�<���<���<W�t<�TF<��<ӡ�;�"�;��`;Y�J;�#n;�I�;�[�;)L�;��<o^<���;�5�;�];��%:�����#����������`X���~Y�~�ͺ��9Z[�:��R;�C�;�N�;��;��;t{r;�{K;�A ;���:�́:w69q�J������!`�Dͬ�Q���.%�X�Q�Ⱥ}���������E��D ���[��%��髈�a�|���r�Čw�څ�����X��Ϗ¼�ּ�M���%9����7ټi%˼�<���e���ר���������3�����R&��z��i2��N���x���Ƽ��̼�ռ�-��Q�y���l	�9z�S��0_$�
�(�ҿ)���&�� �a���d�߳	����K���	��^�v��-e!�=(��,��.,���(��"������5��2j ��P���\�'�輦0�sn�׎�@#�I�A�o����aM�as���n�}m�s	������$���-��K4���7��7�V�3��J-��_%�\���l��@�����"�3%��#.���6��<���?��)?���:���3�t\+���"�����V��3���
��i	��l	���	�OO
�`�
�a�������������  �  .z=�=�g=�[�<J5�<�F�<���<�~�<:��<���</�<���<]��<�(=t�=? =�a�<�r�<���<w��<Z�<��<�%�<5��<G��<���<���<�t�<D={�=g	=��
=��=�=k�=�I=J�
=$�	=E$=�=R8=CZ�<���<O�<o�<���<0�<���<�J�<���<���<�f�<��<�+�<s��<��<t��<�]�<�q�<���<ŵ�<nƣ<���<�U�<���<�<*�<��<�1�<��<o��<���<"u�<���<��<t��<k�<:1�<an�<��<�4�<�A�<���<���<>R�<��}<7cV<q�.<�<��;�;���;�ں;��;�� <�<L�<*�<�<b#�;/ݛ;;�;׈�������B�3=V���8����i�gx:��;\�R;�R};�m�;|A�;
J�;^�e;��B;I+;���:�oV:{��_�T���k��%���������?�S�d�|���P���"��s��+2��y'��dz�Ԏi��Ob���g���z�D匼�5���s��x�Ƽ^�Ӽ�ۼ�ۼb�ּ�ͼ>Vü�и��민|����/���s���妼a䩼�ۭ�Sk���k���Ƽ��m¼�}ȼ�Vϼ;�׼u�����E���0��|�5�	c�� ��� �(.�������$�
���E��j������
��Z�R��i���#�eN#�� ��;��m����������k��p�Ｍ'뼒���R���漌8缊'���D��:���z�����������&�����[&��+�9�.�ļ.�s�+���%�����3��>&�ҧ��N�~F��='���.�N:4���6�$x6��3�"�-�ڸ&� ���2������c ��Z���
��G
��f
���
�W�����\���3��&���  �  ==�=�Y=�S =���<\��<���<-�<�I�<t��<K��<���<�=$=7�=M[=
� =���<j��<��<���<+��<� �<s�<@��<}I�<���<w��<��=e=�=H[=�	=�>
=�{
=E%
=�5	=F�=��= {=�� =@%�</��<f��<�Y�<���<x��<2W�<UC�<ȿ�<v�<8��<Y��<�,�<c��</��<_��<��<�3�<���<ө�<Ŀ�<�ͱ<��<gճ<��<���<9�<��<ח�<�-�<��<b�<��<C�<�~�<�5�<+R�<���<�\�<@��<b�<e��<Qq�<��<t؁<��d<�IF<�*<�\<7<�� <J<& <n�<��+<�h2<(~/<�V!<��<���;n�;DY;��:���=q�^�M��Kk�#v:���:��;��<;�^X;5�e;�'g;��];�<K;�4/;/�;�֯:q��93��fֺ�8�����N������{���.���J� �c�0Iv��X���ڙz��zm���^�lS�n�N�!U��Eg��j���R��}����H׿��ǼM`ɼ�rǼ��¼�g���*��	찼�A��$Z��e������0��&+��`���幼����5Ƽ�>ͼ�Լ��ܼ#�弪���%������	�A3�9��N&��`��(�����0
��^��8������c���X��A����
����½����L=���3��OH��+
�89�a� ��q�������x�TK�a���鼍�鼨��׻켁�����h<��v������>�����v�T[�b���"���$�2c$���!�7�N�����*���b�a��
��	���#�Y%��*�@�,��,��*���&�S"�~�����@�?������\��n�����o�����N�_=�����m���  �  �q=r�	=m=��=$�<"��<z�<P�<���<`��<c1=�L=^�	=�=�R=�o
=]�=,�=���<3v�<�o�<8x�<���<�L�<���<�D�<��<���<6y�<���<�*=�E=�+=��=�V==~�=�=�=�,�<���<S��<�J�<(��<��<��<*��<m�<Q�<J%�<D$�<k��<Ɂ�<pH�<l�<�W�<6&�<���<Q�</t�<���<���<ZT�<`��<vu�<�&�<b*�<���<��<T��<�<�<;��<W�<�Z�<���<�-�<Z��<���<�o�<�o�<�a�<�<�h�<S�<!�<��<	}l<B9X<�F<�7<�.<�*<��,<ߦ3<��<<aAD<�F<�B<��4<�<L8<E��;4�;��D;c��:�թ:%�:��:�Ԣ:���:h�:��;Ѯ;;�;K�";��$;��;Ҡ;Z��:��[:�V:�����0+��~������_ѻHl��8|�V�#��5�0�E��yQ��0X�2Y���T��DL�<C�~<���;��C�r�S�2�k�8X��#G��r�q��$Գ�YX�����E���0Ը�gg���$��T;�������n������+$��k��������7���ļ�g̼��Լ��ݼ7�p��\�����!���D�HT	�Ԗ�J���4�x%
����@M�(���^�� P�f𼘭���Z��������k��v�!���D������=	��c���s]������Z��� ��>�������� ��~���#��l#�hP������
�:L������=��J
�t���'���o��O�'i�e�	������	��(�����<�����s"��j#�E�"�)�!�uz��)��������b�(E�C:��X�Y������v������_��B��k��  �  �U=XT=��=^�=�_=6 =W=�)=�=_�=��	=c�=�=�b=�d=C�=��=�>=�0=V[ =�.�<v�<^e�<B��<)6�<�?�<��<���<���<N�<Y(�<&��<�d=
�=G=��=6U=�h =�g�<D��<\a�<�e�<���<7��<9��<��<)�<��<��<H��<���<kT�<���<s��<P��<��<�k�<�)�<�y�<�c�<$�<3h�<O��<��<w"�<_A�<��<�#�<��<;%�< o�<a��<`��<D��<k<�<���<&��<���<n��<���<��<?x�<�R�<AĊ<���<`�u<Y/j<϶`<cY<J+S<P�O<ӋN<-P<�S<ÆW<4Z<��X<w.R<LE<R2<F�<.	<w�;��;-��;�I;C�;#q�:c��:��t:'0: 	:/�:��>:[Q�:o�:>b�:���:�m:��8$w��Mv%��ۃ�.���&ݻ= �v������"��*���/�m�3���5��q5�x�2�)�.�~*�	�(�]u+��/4��FC���W���o��q��hZ��@뚼2ԣ����������D���Խ�V����4¼��¼%����j������<����C��m�ļ��˼�?ռQ�߼�i꼲������� ���'|��R�A��9��������V������u����0��g輝(�oV������W�����������	���	��G
��h
��'
��a	����M��g������������ ��j#���S��H����������%���!������.�nw��W�����M��:����	�L�� !�]�����l�R���������
����p���o�Aq����d�hC���L"����V�dy�����W��If����������� ��4$��  �  ��<�F�<�~�<�Q =�o=��= =�T	=Q�=��=�=P~=��=�=�}=@G=�+=�n==Y
=�=z�=v =+�<��<!�<���<T��<���<���<���<�x�<Q[�<]��<��<�� =6� =P��<���<���< ��<L��<���<���< ��<� �<j�<L�<�N�<�~�<}��<�x�<=P�<���<p+�<81 =.=�� =Zn�<��</�<1��<�"�<:+�< �<���<���<�J�<,/�<:R�<^x�<�1�<V��<4�<��<���<��<�_�<]6�<���<I��<_�<���<�7�<��s<�-f<<_<��\<)^<Ra< Qd<�Ug<{�i<��k<��l<��l<�Dk<�f<]^<,�Q<�A<�-<h�<�q<y��;�A�;���;tE;��:!5:����<���Ǻ�Ժo3���.f�^>��L�69�T�9��X��w�����q��0m���S��w/��0!�we*�O�-���,��I)��$��� ��"1�`����@��i����ݭ(�A�6��FH��Q\�J�q��u��_��ݑ�������]�����N&��^�ɼ>�ϼ��Ӽb�Լ��ҼACϼ*I˼¨ȼ��ȼrͼ�"ռ'm�w�f��������!	���	�d��/�����8�M@��k��a��
�3�D��Gv�z�Ἶ���伵��T�켌��R��-F���2�H\�f��%�����ۇ�Ba���̒������W��2���&��,~���z�-����
����a��y������~�m�
�����;������
�Up�<R��X�������}��X�+�D����	�`��9������e�����q!��O$�~C&�[�&��&�%�#� ���
4���<+���<�;��g$��M)�'-��  �  ���<�2�<���<���<� =��=�<	==�=�=�2=�=��=�=
�=��=Z�=�=�=,�=��=�'='�=i��<��<'�<��<8�<��< E�<EX�<���<n�<R1�<���<;�<yX�<e,�<=i�<���<!�<=�<B�<;�<���<N��<���<���<���<1��<��<m��<S�<�v =�=�=� =��=J/=X� =�S�<	��<�a�<�r�<Z��<���<���<���<�͸<\�<�_�<$�<�<z��<aú<�W�< ��<Iu�<-�<�;�<��<"��<X<@a<�L<�<A<0@<k�F<<�Q<ն^<��j<y�t<�Z{<{�~<q�~<K|<M/w<�p<{Qf<��Y<�AK<H�:<��(<�<dJ�;B�;��;̕G;�#�:�������!U����L���,u�GpB����Ӥ�K�k��w��[�
�I�q�rL��T �% ��9�҅H���M�w#J�B@�#|2��X$�t���N��Y�p���h�C�	���R��DT!��k.��=���N��\a���u���P�����5����潼�̼�MټF�⼛S��!���弾�߼�ټԼ��ҼX�ּL�߼��켓���"�S��]�	��'L�F���J�3c��q�����a)��뼨��F㼄i༔o޼|ݼ��ݼ�2߼g��w/�:��%���2����O���	���Q���������W��d���@	�K�����3��*��m���S%�D�	� �<D!��n�����L��d�%��M�	��\�>��"��)� �v����������?/ ����U�5���\�.�����ݪ��:��6 �p#&��Z+�j$/�C�0�{:0�&G-��(��##�7&�J��2������ �j%&���,�\�2�H7��  �  ��<���<��<�7�<���<F�=�P	=�~=(S=��=�_=�=�J=�!=��=��=c�=vO=�C=,a=+b
=�= ��<r��<m�<�P�<|�<�Y�<���<��<6�<��<{��<�a�<�@�<F��<M��<S�<�	�<���<���<؈�<嬧<U�<���<��<�a�<��<#/�<AD�<���<bW=��=��=$3=P=n=��=^�=o�=|L�<��<xr�<;��<��<��<�j�<�=�<���<�i�<���<��<�'�<�<).�<���<�[�<���<(é<{U�<�N�<��[<��9<�_#<:<x�<vo+<�7?<U<9Zi<őy< &�<���<6��<��<pW~<gRu<^�j<ܐ^<(Q<xzB<�2<�8<��<�;�$�;�,;j��9�h�󧃻����Ի��ٻ6�ǻ%Ф��%w��	0���
��?�|�X�3�����Û �7fE�ea�S#q�u�s��^j�<�X�<5B��d+�U��-������������f�����n�	x�U�)�(�7�W�F��W��k��聼Z<��R�������<Ǽ�1ڼ������BI��~�������B����n߼�ܼ�f�VO��w��%��Q��������^0����n!�=��հ	���������y�*����Ἡr޼��ܼ�~ۼP#ۼ�jۼ\Wܼ��ݼ�n�)D�M�s(���?������0��!��.%��Z%�[k"�,��X��S��
�˜�8k��t������{K"�N (��>+��4+�o,(�!�"�c�%��J<�(���6�C2�1�������x���A���s�������A���TD���ӭ�!K	�u+�Wg�@��r�#��#,��Z3��8��);�v�:�W�6��1��F*��$����=���� ���%��"-��&5�[d<���A��  �  ���<���<u�<��<�L�<L^ =�;=N�=W6=� =a�=w,=�=��=F1=�=�=br=�=�=�"=�=^�<"��<T��<�x�<-r�<�<8u�<ś�<	^�<�`�<h[�<b��<j��<��<���<���<�b�<��<6��<뙗<�ʕ<�}�<^��<�̷<=��<�y�<��<��<7��<E�==��=I�=��=ˬ=ZV=K�=/�=�� =���<���<2��<�U�<f��<��<���<�Ǎ<΄<�ւ<�ԇ<�F�<>h�<,ū<;��<Az�<���<���<1��<ֆj<�&=<��<���;U*�;��;�x<V�+<%�H<�fc<��x<��<��<V�<!�<���<E�w<ܧl<ت`<��S<�ZF<��6<R�#<�4<h�;���;5�;`�<��`��O���_��`���������]޻#ޫ�&��VO��.V�'֍�B�̻b���i<�oce����(\��y�����wp��XS�~�5�+�����{����컫ﻝ������z������'�I�4���B��TS�X�g������������^ܹ�!�м�6��x��%7���8���F�U���5�� �`h�P��a�o��.�vi������$�N(&�Z�#� ?��]�nx����������伄*߼VܼS�ڼ�ڼ�ڼ UڼM�ڼDܼ�޼���b���#�0
���%��x�*�-#��*�7.�IY.�V�*�8�$�����������֙�(�Ė��{!��*���0�yE4���3�k0��h)�� !�q���3�����c �����W��������Ŋ��G���+P���6 ����Wi��X�s���U�KC��"(�U2��:�� A�[*D�kC�?"?�E8�"Z0��")��7$��"�%���*��3�c=<���D�baJ��  �  ��<��<*��<�K�<m��<Q�<�=�/=MU=��=�!=�=m=L�=h==�==��=�	=��=�(=�b=AB�<<��<:��<;;�<|�<�ۙ<7$�<�ɚ<^��<M,�<���<a\�<��<\�<h��<$s�<�޸<��<�^�<6j�<���<D��<�t�<���<���<���<��<M��<�" ==ۘ=E(=�9=�=D�=ԟ=,=�B=�o=g�<4C�<��<n��<���<�"�<C��<|�<Bjq<X|m<��x</:�<��<y��<��<��<��<���<�6�<7�X<�{(<�� <l4�;X�;��;���;_S<a�><Jm]<�[v<z��<OՇ<xQ�<~�<Ю�<��x<�km<Nxa<�U<��G<7�8<�a%<ƥ<;��;���;K�:�pźmǒ�oQ��G�0'��(�.������Y̻E���.Z}�N���p���&��i�;1O��
{���*�����E���>�fz`�v>��c ��b	��������Á����/�����P�0J'���3�vA�^�Q���f��ր��������߾�iؼ��;��>D
�4����y�	����.���Ŧ��-�^�x~�����\w��v���$���*�TM,���)��K#�Il��k�ؕ�5����[�F޼�ۼ�ټ�xټ�ټ�ټ�aڼ�Aۼ�ݼ���nB�ho����u���I����(��/��04� w4�Ӭ0���)� � �Q�=��]���m�T�:[���%�*`/���6��k:�::�L�5�-#.�?�$�q���S��v	�f���_��U���n���_��+�����WK��Я��g���pZ����y.�SL�?s��Z ��R+�BM6���?��G�ORJ� tI�T�D��!=�+q4���,��)'��y%�'�'�{-.��7��A�J�|`P��  �  A]= "=(=��=�E=d�=3$=(=�G*=�++=�+=;W*=re)=�(=9�'=�\'=7'=��&=C&= %=�"=��=��=�=�=�=�=;��<��<z*�<se =d=�&
=�]=��=��=[x=^�	=54=�x�<Qq�<�-�<���<�P�<��<<E =s=��=�H=�=�=��=�u=]�=VM=H�=�=�s=A�=��=�=��=�?=_O=�=�� =��<�?�<���<��<��<e��<���<�	�<���<~��<�<�<�<�>�<�G�<�J�<}��<븝<8'�<"͏<��<
2�<�N�<��<p�<�ݯ<��<A�<fӭ<ۨ<��<8ڜ< �<a�<>C�<!X�<�,�<�,x<̧h<t�T<U|;<|<�%�;��;�;�;��);|��:���:���:��;��U;�S�;��;��;@_I;��:�Ny���� ��_����SϻQֻ� ʻ��������0�^���(�V���-�����M['��oQ�<~��裘�#���&�Ļ��ػ�u�S� ��"�:1�N35��GP��jo�]L��煘��˦�阱�ٷ�B��K{����������������)X��鵱�e����̼�ۼ�R��x４l�K�|?�Jg߼~@Լmjɼ2��7m���Z��3�������&����ȵ�L����1���3�������;ŷ�L��<����Ƽ[Ѽ��ݼӟ�ؿ���, �c���U�6C�F���^�g�:�޼�Yۼ��ܼI�����SY�����N	�B	�������^R��7����Q�ܼ8(׼qԼ��Ӽ&ռ�ּS�ؼ�ڼuۼ&�ۼ�ܼ��ܼ�޼��⼕_�k��`b�����ω�I��� ��C����t�@1��:���������������
��N���� ��& ��  �  �=+^=�F=��=�=!A =��$=�C(=�[*=;2+=7+=�a*=�w)=��(=o�'=t'=�)'=��&=:G&=�%=��"=�-=DI=^V=��=�=m/=d�<�l�<���<\y==��
=��=�Z=~i=I=I�
=�
=r|�<��<��<`L�<���<`/�<�%=��=s=��=Q�=��=+�=`{=I�=�a=��=��=�=��=s�=8=7�=�_=��=Gq=Y=\��<�Q�<��<�z�<t5�<�C�<���<M��<7!�<��<�#�<AD�<�d�<���<d��<���<��<ژ�<�:�<���<c"�<�؝<�8�<���<�C�<O�<M �<�ҭ<��<[�<��<] �<���<rr�<�y�<�C�<'bx<li<�_U<i�<<75 <<<��;�K�;��=;�;Q��:��;2v/;Ĝb;ړ�;|j�;�9�;oR;�i�:iac�F.���x��*���vŻ �̻Vv��;���]��j�V���#�\�!��۬�J'���P�z��뿗�����Ļlػ����� ����ա��.4�_�N��l������x���k��Y���>���ȶ��D���%��p���K��j���d8��؀��L�����ʼ�ټ&��;�� �����;�ݼs�Ҽ�~ȼR���s#��~=��0������y������䄶���������ڶ��඼�����2������_sƼ�{м�]ܼ���#���b���V����� �kr�����_ ��ݼZAڼ��ۼ�἟��&M���I����
�j �K��W���������H ��(ܼO�ּ�]Լ�Ӽ[�Լz�ּ�aؼF�ټ��ڼ��ۼtܼ��ܼ.�޼ɽ⼩	�A�Ib��������o����H��Y��XT��8��m���t(��k���
�������5�����  �  �5=�=�d=BZ=n�=�!=	�%=W�(=Uv*=�*+=�+=o*=��)=��(=)(=��'= L'=[�&=j=&=�%=<�"=�=�8=��=��=�C
=	e=b=%� =�=�=��=�=W�=��={�=V�=��=�i=2=nF�<'��<,k�<4u�<�<��=�=�==Z9==��=I~=�x=7=��=?=L�=l�=��=��=�=�=i�=�(=�=�=FM�<��<G��<�z�<*�<���<�S�<_b�<��<���<� �<�(�<���<���<	��<�|�<t��<���<|�<��<���<
�<�;�<Ԟ�<51�<�Y�<=�<̭�<��<R�<�u�<|��<� �<�܌<.��<�V�<��x<�i<9W<9@<R�%<�<ހ�;�@�;�-u;��?;��,;��8;In[;od�;{V�;���;}��;�j;��;���9�䲺pH��8������%������������u�ŢA�bl�r��qG���,	��k'�ǁO�f�|��~��^#������nOֻ��� ��{�؟���1�#�J�F�f�>��mߐ�xݝ��䧼���4߯�����੼G��J���$V����#������SƼ�FӼp޼g�弎��R��l(�'�ؼ�WϼfƼ�J��L����$�����\���4V��;?��#���~�� �������'඼ҷ�%��
}��@9ż/Aμ��ؼo?�����L���P��M������h����l�YIڼ@2׼O�ؼ�_޼��`=�����P��{��z��h�i{���P�����]�Iۼ[�ּ^Լ�Լ'�Լ�aּY�׼�Xټ}fڼ-ۼ��ۼ��ܼ��޼��gV�g~�����1��	��^��X��k��O�Z&��z��(
��2�k��8��Ӈ��6��M����J��ox��  �  �l=~�=�=��=d�=L#=!x&=m�(=�9*=��*=i�*=�K*=��)=�)=i(=S�'=~Q'=��&=�%=.�$=̼"=��=�6=@�=��=�=I�	=$$=��=�=�	=�o=R*=�U=�(=	=?=|=(�
=�M=�q=| =���<� =K<=j�=��
=�=��=:=�~==c4==��=�Y=5=��=��=�G=��=�z=��=�=c�	=r0=�H =��<�!�<��<3X�<y@�<���< S�<���<���<��<J�<�a�<'i�<��<��<�(�<
��<!	�<O$�<��<�Ч<�<1��<���<��<�5�<��<n�<_M�<�ѝ<�8�<���<�(�<��<�<�^w<�i<��W<�C<)Z,<�s<�0�;���;���;K �;Y�~;/�;8�;�$�;���;q#�;��;3�;c49;��:$Mݹ�����DO��Ҁ�|���}��ȴq�k�L�{�'��������L���3��",��Q�^�z��(��=M���?��ջj3��J��X���Y.0��F��^���x�q��]~��0��� d�����Xꤼ���G���Yg������?���@���ϲ�羼d�ʼ��Լ�ۼ�O޼�(ݼ0�ؼ�0Ҽ�ʼ�Zü���؋��{���r��^+���v��o����������l]��&����]�������ͺ�K���,:ļϵ˼��Լ��ݼ[�����I��<��m�� ���(ۼ�hռ��Ҽ�%Լ�PټD[����S��"���_���S���̀������`���漦�߼Hiڼ��ּ�ռ޾Լ�Rռbּ�׼��ؼc�ټVۼT"ܼ�ݼu�߼l㼝�&％���� ����
�Fe�n6�G4�u�}j
�����s��8�V� �
<�ۆ��
�q���?��d��  �  �a=l=��=r�=�"=��$=��&=�/(=_*)=o�)=��)=ګ)=�f)=_�(=lp(=��'=��&=~&=��$=Ā#=s�!=Lt=��=�6=L�=0= =��=��=�z="C=��=��=uE=g�=M�=��=��==�8=�=a�=�G=��=0�=h%
=��=�s=��=�I=�^==Y=�~=}=�X=9=g�=�%=rr=�=�Q=��=�Z=�q
=b=�a=S��<&��<o&�<�<�F�<d�<�b�<���<e��<���<q��<���<J�<@Y�<���<wC�<=9�<;:�<��<^
�<P�<t�<Z�<s��<�ٯ<�í<��<O�<;�<���<�Y�<;��<`ӌ<9��<�M�<RYs<�1e<�U<'DD<o71<�.<�R	<�;w��;^�;T�;��;��;87�;���;�^�;N�;!��;>=h;Z>;<1:-&1������$�k�=��B��8�@'�ǋ�œ	���\�T!�G�:��Z�ݳ}�⚒�����E���Bxֻ�L�}���%��� ��a1���C���W�bm��Ѐ�3��q㑼b9���뙼�<��S���O;���`��@������U�����@���'����ɼ[�ϼxҼVҼ��ϼ��˼_�Ƽ\����_��g&������졶��ܵ��v���]��n���1���!���k���i���C�������P����ļPDʼF�мL�׼��ݼ� ��G�b�����༃=ڼ�bԼC�ϼ��ͼI6ϼ�ӼF?ڼo�἞c��7＾��3��C�"u�*��T��k�޼�9ۼ��ؼb׼�ּ��ּ�*׼<�׼��ؼڼ��ۼ�Mݼyo߼��YG���C���q��C���l��BO����E	�5N	�b��������M ��:��U����V���s��1��9
����͆��  �  6*"=N�!==�!=�"=��#=!�$=Z�%=C@&=*�&=`'=Y�'=`F(=փ(=lu(=u(=.'=��%=O~$=��"=�0!=�x="�=�=�=ee=oN=v�=6F=5�=l9==�Z=a=�=H�=ܾ=VZ=��=�=*!=�=e�=��
=.�
=��=��=�=�=H7=-=�=��=]�=�E=Z�==�=`�=,�=f�=��=�_=��=�p=`�=	�	=��=�=�r=��=L =(x�<4�<�
�<$* =� =K@ ="��<���<T��<5��<���<n��< ;�<R}�<!͸<��<Z��<C�<�į<���<x�<�)�<u�<rp�<���<�`�<lk�<��<���<�Y�<�=�<	�y<�j<�}\<K;N<��?<x{1<��"<��<'�<D��;'��;���;��;p��;{��;\��;�#�;���;H��;0��;��E;�0�:�P:��ϹL%��yغ"6 �C���y��Tp��&��4�$yE���X�Y=o����������������8�ܻ���!��ft�)�Ϩ7�(�F���U��e�p�s�a���ˆ�cQ���3������܏��揼����bҒ�/��˃��𐥼ec����zL����ü�Ǽ�Qȼ;�ǼF�Ƽ��ļbI¼93���V��U��������W��NⷼB׶�Et��wܶ�U������a��9�������ļB�Ǽ�?˼�ϼ��Ҽb�ּ�eټCۼCۼ�Yټ1ּq�Ѽ�ͼʲʼt~ɼ��ʼ�μ�JӼkHټ=߼����漗:���w����iu��a�Ǥ޼[<ݼ>	ܼ��ڼ��ټ?Bټ�ټ�ټ�ۼy/ݼ�߼�'㼪��%�鼓��`�8����
��Im��:.�������z������ ��
��
����[��LD�����k����m�;���z���
��  �  |'=��%=��$=�,$=��#=#=H�"=)�"=#=��#=��$=��%=��&=�H'=%�&=�%=�0$=�"=T�=�=�=Q===�f=I�={4=��=ʣ=<�=�5=�=�6=�g=�Y=��=r=�_=��=��=Kj=�r=)�=Ġ=��=�=�=�Q=�'=*3=�=L=ml=z�=W0=�F= �=�=Q�=��=W=�=45=Խ	=��=��=�=�_=i�=�=Ћ=3=O�=6�=��=�=o=B =���<[��<G��<���<U�<:��<���<7I�<�s�<E�<���< f�<��<�?�<Y��<#l�<4۟<r�<Ҥ�<<ۙ<���<j��<2h�<P�<r�n<��]<8)N<�@<�U5<�{+<��"<��<'�<b<��<�9<���;���;���;7�;ܶ�;KN�;*X�;ڟ�;.Mv;�*1;?��:�,M:�y���1��ۤ���躒��6/���H�K
_�[�p��~�a%�������[��Y����Ұ��5ʻB"�p���A�
�'���6��D��}O���Y�#�b�ѵk�@�s���{�g/��y����-��eU���;܋����!����S��(���H���D���}��������Ӓ��m�¼Fcļ{}ż�Ƽ�.Ƽ��ż�ļ���R澼���!������`���3ߺ�����e����ż,ɼ��˼��ͼTgϼdsмj8Ѽ4�Ѽ��Ѽ��Ѽ�ѼD�ϼ[ͼ��ʼ�Gȼ�Ƽ�Ƽ�Ǽ!�ɼ�kͼv�Ѽ�ּ��ټ5�ܼ�Q߼w�Y�⼉����伒��0�!��/[�a�Z߼8�ܼV�ۼ$�ۼ�Mݼ�W��r�	�C���l����� ������li���������oE��%o��{���
�������0n������)������������#���n��Ɍ�x������  �  �w*=~(=�W&=�$=��!=� =ܕ=�=�=�'=�� =0�"=Q{$=�n%=iM%=�#=��!=��=O�=��=��=��=�;=n�=�n=�y=��=T�=�J=3�=1�=�=9�=�=��=`}=��=_�=�+=��= =��=��=�=�=�=�+=��	=��=g�=Y	=x�
=R=K=�=c=��= p=�#=�Z=��=GC=��=8�=}=��=Ղ=�i=�%=-�=�=`^=P�=�=J�=�@==5��<E�<��<)��<��< ��<E��<���<�ʾ<�ȶ<��<�Χ<���<抜<.7�<|��<8�<8w�<p[�<'�<�T�<�J�<���<�Gt<�_<��K<T�:<S�-<r�$<�<�<�j<�G<3�<��<sQ<�a<u�	<'�<}z�;���;��;/��;¨;k��;�_;\%;���:�P:;���fx��L��*/��b������ߖ�雠��<������U(��Ć��Ύ��ܼ�-ػ����$�	�&��:�0J��:V���^���c�9qg���i�1ml�:�o�ʤs�p�x�p~��끼�����a����M��͈��O-������z����	��� ���
��l컼	���4�ż;�ɼ�ͼ!ϼ=xϼ<�ͼ��ʼ�SƼ���������m�����+�ü�ɼ�~μ$�Ҽ��ռ�׼*�ּ�ռ{�Ҽ�/м�ͼ+�˼��ɼ)ȼ��Ƽgiż�YļD�ü@�üV�ļ�Ƽ!/ɼ�̼�3ϼ�iҼ��ռ�bټH]ݼ����c��M��G��|�������q�弰9��߼�߼������F��b��(���ak���k��أ��U[��4
��%'�����}6��X����n���_���g�z��s������m���������R ���5 ����  �  �^,=��)=�2&=\�"=e�=έ=�I==�L=��==C=�=��!=�#=^#=�!=ڐ=F�=��= N=��=��=�=�=��=�<=��=��=WR=qI=��=�=��=�=`=��=�V=K�=��=�=t=��=)�=7�=�t=j�
=��=*�=K.=t�=��=��=��=��=�d=P�=>�=_�=�
=R!=��=�� =��<��<�`�<�� =55=ƍ=P�=L	=9�	=��	=��=�=��=5�=�K=&#�<�'�<ݵ�<v��<:��<#��<V��<0�<j�<�J�<��<^��<91�<��<�L�<�O�<�Z�<�]�<��<��<� �<�Ǉ<}<�Ef<>N<6A7<
[$<-< �<h�<��<'�<�m<N�<h<��<��<��<*[
<�<��;��;D
�;��;`��;�a{;��F;�~;�ݟ:IK 9��J~�Ya�pH��2����Ż� ϻz�λ�Ȼ�:��J𹻡Z��Zͻ�,�D	��� �}9���N��v`�o?l��>r�(ys��q�\Mn��Nk���i�k���n���t��#|�F���Ɇ�+���ZM�����e發����c���E��薭������s������ɼ)�м�hּڼ�!ۼ�@ټ��Լ��μ �ȼ�uü!���A����Wļ�Bʼ�vѼ�ؼzF޼��&I⼱N�$Wܼ�3׼J�Ѽ�̼�_ȼ]\ż0{ü&|¼�¼¼n¼aüZ�ü�/ż��Ƽ��ȼ=�ʼ��ͼʘѼ��ּ��ܼ���$����`�������|h��������$���輼�伪��o��]�꼧��s����� ��x���2�B"��2�u���1���V��\�`�����m�p�％�S��� ��X�j����������3����N���  �  t�,=�W)=J�$=" =^=Q�=�=%"=s=�t=�=#M=߆=�� =;� =�=a=��=p�=��=Y�
=��	=ߝ
=c�=�7=��=��=��=�=1b=��=��=\y=F�=�d=��=ju=P
=��=O�=��=�=��=0.=��=�=�= ��<g��<�{�<B��<,� =�o=�W=�=-K==h =uX=��=a��<���<ם�<���<D��<�,�<�	 =W�=L�=�.	=ko
=�
=��	=�'=�=G�=5=���<�,�<c`�<=�<փ�<���<��<��<C�<˯<���<�X�<��<z�<>�<?�<p~�<n2�<�v�<Ә�<�E�<o�<�xq<��W<�p<<ʚ"<~�<�1�;���;��;Ȃ <i�	<n�<��<�?<�<m9<T�<7�<��<��;��;И�;�S�;�ؚ;�]�;%W;�;���:x��8����o<��`��X�����޻h��>���c{���{���ܻ�qѻ˵л)߻s����B���/�OWK�d�RNw�������N���>�n�v��n�0�i���g��j���o�7x������-��ST���8��.�����_���0��g㥼�����ʲ��s���:ż`ϼ��ؼ ��-�弲�v��C߼�׼��ϼ"ɼ$�ż��żV�ɼ-Ѽ8�ټ���o��R��e��v����/eݼ^ռ��ͼ��Ǽ.�ü33��	V��u|���1��	#¼zü��ü<�ļS�żf�Ƽ(�ȼ~�˼м�lּ��޼��缴������ �L���#����Y��2�����꼄X�P����5���n�����H	�3�L�
�+	�t�0z��������������3x�n�C8��l�{���T=��Z������;/��1����6���  �  ��,=�{(=�.#=%O=v=�U=.�=��=d=u�=��=�=��=�<=�=!�=U�=e=��=�	=��=��=��=[�=)�=�=�$=~=��=*�=�I=�%=��=k�=4,=��=L=<=��=�(=�=��=�=�=�
=�=��<�,�<ޅ�<��<` �<՚�<'� =�M=�		==��
=��=@^=�v�<Q<�</��<�0�<��<q-�<���<D��<�j=��=�=�h
=y�
=��	=F=��=�i=?� =N�<���<@�<���<��<�+�<�u�<B��<�ٹ<�۪<7��<+��<Q3�<÷t<r�m<��n<�v<h1�<Ǆ<�݆<��<�|<�Lg<F�K<�K-<�<)��; (�;��;/��;x�;��;��<�<�K<w <�<P�<�<Ԩ<K��;�}�;TV�;�.�;F�;�-�;��[;"!;{�: �"���[�h������߻W��f���������c_�����*������I����<�F[��^v�&�����Y������7��|+��g�t��l�3�g���h�w#n���v�j����C��Ŭ��C�������^ߘ�����e�����ST���������?ɼ]ռ��༹���8l�E��缱�޼G�ռ�"μP�ɼ|)ʼ��μ�
׼�2�K뼏b�S����A��QT����C��%�ټ:Xм׻ȼpüޅ��ؘ����� ���m¼��üfpļt ższż�=Ƽ��Ǽk�ʼ�м�׼�p�i�켭i�������G��I�?a��������������`�$���A���XM�0s
� N��8�f������	�<H�� �����z��v�켞��u��m}�K%�e��S��v��wH��ʈ�����������  �  �\,=�'=��!=KI=�=�1=+=<X	=�	==�=�=��=�=^�=S=��=9�=r=t=��=�Z=�=�F=�=�C
=��=�=�Y=٣=�=S=�*=ҁ=̮=h�=e=P=l�=�=y3=��=]�=Z�=�=�	=:�=}�<��<ov�<P��<PL�<!��<to�<�?=WQ=^�	=a	=��=7Z=͋�<_^�<�R�<��<e~�<���<�,�<��<Le�<�c=��=�
=/�
=�	=2=-�=�!=�` =�[�<� �<���<%_�<���<���<ڻ�<3�<zP�<u�<B��<��<Ʈv<�Jf<�n_<��a<Ͻj<��v<0�<���<���<S�v<^T`<!C<:#<)�<J��;���;�k�;��;[)�;�}�;e<.�<��<��<�<�<�E<X�<���;f�;� �;K��;�s�;^��;�[;�r;wI�:�fù���[���F»��������N� ��m�Og����{)���O�Y�������&��E���e� f���d������6��A��a��Dփ�R�y���n��i���h��m���v�ƀ�����I������Z�����b���xE�����!�����������ej̼_�ټ>\����������z4�������ټ��Ѽ	ͼ�9ͼ�2Ҽ7ۼI漦#�>��5��DX�����O��B�rݼ,�Ҽ\�ɼ1�ü����󂿼4���U���¼�ļ0�ļ�\ż+�żH7Ƽ�Ǽ˼��м�ټ|�㼝[��H������	����
����	�$��6� �%���T򼀾��A�T\�����������޷���jp�������`���Ĭ��~a󼡾�����������&���e������q`��sx������� ���  �  `,,=J'=�>!=&�=v�=�=��	=�=V�=�=�=�=@i=�=�v=vZ=�=J=�#
=F�=m=s��<�=�s=BZ	=-�=�a=�=�z=	�=�M=�%=v=0�=c�=nK=� =�=b�=a/=S�=�=�=G�=��=��=rs�<<H�<���<%q�<���<`��<~��<��=��=��=*�=<=�=V��< K�<s��<��<���<*�<��<+P�<��<��=�=��	=��
="�	=;%=m�=m=I@ =A�<���<R��<�I�<6��<���<�i�<���<�\�<�¥<y��<Ty�<��q<�1a<�nZ<�]<��f<��s<�#<�q�<>�<Z�t<�]<�@<�d<Ep <L0�;�; z�;"��;-V�;}L�;��<�<B�<�{<�<V�<�<��<]��;�-�;�@�;��;T�;ž�;�yZ;I�;��:ط�C�x�����ɻ��t�,�"�U�%������������:��>��G�Q�)���H���i�����rԎ��3��q��:8��<ꌼ�9����{��p���i�-i���m�Z�v��܀�u���GH���C��6����*�������J��/&��!㫼 ����n��B�ͼ!jۼ#c�b���n����������Ｄ�弍Aۼg�Ҽn#μ�Rμ�fӼ@zܼ3��5�?^��k� ��� �uS���������D޼�\Ӽejʼ�#ļ���\�������r����¼pIļ�ż]�żd�żvBƼx�Ǽ	˼b�м��ټ���ٴ�������U
����B��
����>��_���0C���`�f���{�����ƚ���.����������J%� ���f���������K�����k��1F�H������Gt��;���b���#+���  �  �\,=�'=��!=KI=�=�1=+=<X	=�	==�=�=��=�=^�=S=��=9�=r=t=��=�Z=�=�F=�=�C
=��=�=�Y=٣=�=S=�*=ҁ=̮=h�=e=P=k�=�=y3=��=\�=Z�=�=�	=:�=}�<��<nv�<N��<ML�<��<oo�<�?=SQ=Y�	=a	=��=,Z=���<>^�<�R�<^�<+~�<���<{,�<[�<�d�<�c=y�=�
=d�
=��	= 3=��=�#=`c =�b�<0)�<���<�j�<���<��<���<.�<�a�<U1�<*Ж<���<��v<>jf<��_<)�a<D�j<�w<H�<���<O��<F�v<�J`<�
C<��"<��<���;���;�)�;�h�;:��;X6�;f�<�`<Za<��<S�<�<�5<z�<5��;}�;�*�;c��;%��;<#�;t[;��;�D�:G,������d�����)����e�%���� ��T��R�������E�/�����r'���E�N�e�s��ts��0�������}.��s郼�y�uo��5i��i�I�m���v�mр�v���l ����P`����������G��l��E���g���=����j̼��ټ|\�#�����5����4�������ټ�Ѽ$	ͼ�9ͼ�2Ҽ9ۼK漨#�?��6��EX�����P��B�rݼ,�Ҽ\�ɼ1�ü����󂿼4���U���¼�ļ0�ļ�\ż+�żH7Ƽ�Ǽ˼��м�ټ|�㼝[��H������	����
����	�$��6� �%���T򼀾��A�T\�����������޷���jp�������`���Ĭ��~a󼡾�����������&���e������q`��sx������� ���  �  ��,=�{(=�.#=%O=v=�U=.�=��=d=u�=��=�=��=�<=�=!�=U�=e=��=�	=��=��=��=[�=)�=�=�$=~=��=*�=�I=�%=��=k�=4,=��=L=;=��=�(=�=��=�=�=�
=�=��<�,�<ۅ�<��<Z �<͚�<"� =�M=�		==��
=��=,^=�v�<<�<���<c0�<���<�,�<&��<���<Hj=F�=��=�h
=��
=��	=�G=�=Sm=R� =?�<}��<*S�<��<F�<�G�</��<þ�<_��<���<�ڛ<$؍<�S�<��t<%�m<��n<CGv<�A�<�҄<P�<y��<>�|<e:g<<fK<�&-<��<�P�;���;���;OX�;���;�~�;8�<��<><7@ <�<��<Qc<��<$��;*|�;
i�;�U�;���;�z�;�J\;�;�Ч:oZ�����lg��{���D߻d]�`�t��������!���廌⻪�ﻗ�����t=�H[�ʐv������؋�.|���>���\���P��nu�uTl�#h���h��[n�%w�aƀ�zV������0������r瘼:���Pj��/ ���V����������?ɼ�]ռ ��	�H��nl�n�����޼Y�ռ�"μZ�ɼ�)ʼ��μ�
׼�2� K뼐b�T����A��RT����D��%�ټ:Xм׻ȼpüޅ��ؘ����� ���m¼��üfpļu ższż�=Ƽ��Ǽk�ʼ�м�׼�p�i�켭i�������G��I�?a��������������`�$���A���XM�0s
� N��8�f������	�<H�� �����z��v�켞��u��m}�K%�e��S��v��wH��ʈ�����������  �  t�,=�W)=J�$=" =^=Q�=�=%"=s=�t=�=#M=߆=�� =;� =�=a=��=p�=��=Y�
=��	=ߝ
=c�=�7=��=��=��=�=1b=��=��=[y=F�=�d=��=ju=P
=��=O�=��=�=��=0.=��=�=߃=���<a��<�{�<:��<&� =�o=�W=�=K= =Q =YX=��=��<p��<T��<#��<���<%,�<	 =�=��=@.	=~o
=��
=f�	=E*={=��=g=��<}C�<}{�<�\�<§�<���<\��<�?�<%�<���<�ʢ<���<L�<��<pe�<�.�<���<�I�<6��<4��<�G�<�܂<6_q<R�W<<<<�Z"<�L<���;� �;i��;�! <�$	<��<%h</�<Ub<��<n<��<��<���;Q�;k��;��;�+�;˄;�X;Q;��:H��8���:�#������(޻l����4��,����W�ܻ�7ѻR�лl߻����}b��0�\�K�bd�۟w��Ɓ���Eꂼ�t�g5w�odo�	�i�2-h��lj��2p�a~x�����H���j��FK���Д�Q��
��"7���祼�����̲�'u��<ż�`ϼ��ؼ��༒���缱��p߼�׼��ϼ$"ɼ2�ż��ż^�ɼ3Ѽ=�ټ���r��T��f��w����/eݼ^ռ��ͼ��Ǽ.�ü33��
V��u|���1��	#¼zü��ü<�ļS�żf�Ƽ(�ȼ~�˼м�lּ��޼��缴������ �L���#����Y��2�����꼄X�P����5���n�����H	�3�L�
�+	�t�0z��������������3x�n�C8��l�{���T=��Z������;/��1����6���  �  �^,=��)=�2&=\�"=e�=έ=�I==�L=��==C=�=��!=�#=^#=�!=ڐ=F�=��= N=��=��=�=�=��=�<=��=��=WR=qI=��=�=��=�=`=��=�V=J�=��=�=t=��=(�=6�=�t=i�
=��=(�=H.=p�=�=��=��=��=�d=>�='�=C�=��
='!=Y�=z� =z��<-��<�_�<>� =�4=<�=ז=		=_�	=Ŏ	=u�=��=O�=׿=�T=�9�<�C�<*��<@�<K��<"�<f��<sh�<"<�<}��<'٩<K�<�i�<�<�|�<|z�<�~�<�y�<��<��<S�<>��<��|<�f<*�M<��6<��#<;�<�J<K\<�T<tp<��<�d<]�<�/<�L<os<�%
<2�<��;��;
+�;�&�;�"�;an|;�8H;��;w'�:q�<9�Q����%_�Y������k�Ļ
Aλ�*λ�yǻ:Ѿ�V���8��ͻU�mj	��!��M9�MO���`��l��r��s�r��n�g�k�soj��k��8o��u�K{|�Zl���ꆼ�����c���/��t���,����j���K������ݟ���u�������ɼ�м�iּ�ڼ�!ۼ�@ټ��Լ��μ@�ȼ�uü3���N����Wļ�Bʼ�vѼ�ؼ}F޼���(I⼲N�%Wܼ�3׼J�Ѽ�̼�_ȼ]\ż1{ü&|¼�¼¼n¼aüZ�ü�/ż��Ƽ��ȼ=�ʼ��ͼʘѼ��ּ��ܼ���$����`�������|h��������$���輼�伪��o��]�꼧��s����� ��x���2�B"��2�u���1���V��\�`�����m�p�％�S��� ��X�j����������3����N���  �  �w*=~(=�W&=�$=��!=� =ܕ=�=�=�'=�� =0�"=Q{$=�n%=iM%=�#=��!=��=O�=��=��=��=�;=n�=�n=�y=��=T�=�J=3�=1�=�=9�=�=��=`}=��=_�=�+=��==��=��=�=�=�=�+=��	=��=b�=Y	=p�
=H=K=�=O=��=�o=h#=lZ=e�=�B=��=��==
�=@�=Bi=)%=�=!�=\_=]�==��=�G=�={��<l4�<G��<���<K��<���<���<��<b�<��<�G�<Q�<�¡<�Ŝ<�l�<Ͽ�<�_�<���<�q�<���<�W�<hC�<��<t<�9_<~mK<�k:<�E-<j2$<Q�<o�<��<z�<zS<P<�<�<(�	<.U<�'�;��;���;���;]�;�	�;a0`;�&;���:LpW:ei%��p��	��-���_�������.Ɵ�������!���!8���h��#߼��=ػ)����b�M2'��h:�s�J�N�V�� _�;�d�H h�c�j���l�p�i&t��y� o~�����:������+��f�����=�����j���R��U%������������ż:�ɼ�ͼ�!ϼ�xϼ��ͼ;�ʼ�SƼ����5��&���m�����3�ü�ɼ�~μ(�Ҽ��ռ�׼+�ּ�ռ{�Ҽ�/м�ͼ+�˼��ɼ)ȼ��Ƽgiż�YļD�ü@�üV�ļ�Ƽ!/ɼ�̼�3ϼ�iҼ��ռ�bټH]ݼ����c��M��G��|�������q�弰9��߼�߼������F��b��(���ak���k��أ��U[��4
��%'�����}6��X����n���_���g�z��s������m���������R ���5 ����  �  |'=��%=��$=�,$=��#=#=H�"=)�"=#=��#=��$=��%=��&=�H'=%�&=�%=�0$=�"=T�=�=�=Q===�f=I�={4=��=ʣ=<�=�5=�=�6=�g=�Y=��=r=�_=��=ߓ=Kj=�r=(�=à=��=�=ߤ=�Q=�'=&3=�=�K=fl=p�=J0=�F=�=ڌ=1�=��=%=q=�4=z�	=�=%�=i=V_=׼=_=��=�=g�=g�=?�=
$=,"=]L =��<���<��<���<#��<���<f7�<���<��<o��<h�<��<`٩<}�<���<��<J�<q��<���<8�<U��<߹�<|V�<��<�@n<0:]<�M<�K@<F�4<��*<$="<Xh<0M<��<�E<;�<&�;.�;�{�;P��;���;�J�;[~�;8�;#;w;
c2;h��:�T:�2�7�(������T�1���-���F��]��o�l�|�e�������
���Ν��հ��cʻ�y�o�����T(��l7�4�D�P��:Z�J�c��Jl�}t��|��r���;��jf��7!���҉�\���/��b����h���'���U��"N������#�������p���V�¼�dļ�~ż�Ƽ�/ƼT�żļ\����澼���>���(���p���?ߺ�����l���
�ż
,ɼ��˼��ͼUgϼfsмk8Ѽ5�Ѽ��Ѽ��Ѽ�ѼD�ϼ[ͼ��ʼ�Gȼ�Ƽ�Ƽ�Ǽ!�ɼ�kͼv�Ѽ�ּ��ټ5�ܼ�Q߼w�Y�⼉����伒��0�!��/[�a�Z߼8�ܼV�ۼ$�ۼ�Mݼ�W��r�	�C���l����� ������li���������oE��%o��{���
�������0n������)������������#���n��Ɍ�x������  �  6*"=N�!==�!=�"=��#=!�$=Z�%=C@&=*�&=`'=Y�'=`F(=փ(=lu(=u(=.'=��%=O~$=��"=�0!=�x="�=�=�=ee=oN=v�=6F=5�=l9==�Z=a=�=H�=ܾ=VZ=��=�=*!=�=d�=��
=-�
=��=��=�=�=E7=�,=�=}�=T�=�E=K�=*�=G�=�=?�=W�=�_=��=;p=��=��	=?�=c�=-r=��=. =�x�<\6�<��<�- =H� =�G =��<J�<���<���</��<���<�q�<���<;�<�7�<YŲ<G3�<��<�Ү<jK�<�_�<��<��<�ã<w�<�w�<���<cّ<�H�<0#�<=py<�j<t\<��M<�y?<�0<�t"<�f<�o<G��;���;T�;M��;�L�;�\�;�3�;���;K��;\��;5ъ;U�F;���:�!:D¹/v��րԺYB�����.����ps���$�K�2��D���W��Tn��τ��������� »�ݻ���������~)��#8��G�LV���e�R�t�Q'�����h���Yp��1ŏ�����������i񒼨5��;���󠥼�o��
���JS����ü#ǼsTȼ$�Ǽ��Ƽ��ļ.J¼�3��W����������W��sⷼ]׶�Zt���ܶ�a������a��>��"�����ļD�Ǽ�?˼�ϼ��Ҽc�ּ�eټCۼCۼ�Yټ1ּr�Ѽ�ͼʲʼt~ɼ��ʼ�μ�JӼkHټ=߼����漗:���w����iu��a�Ǥ޼[<ݼ>	ܼ��ڼ��ټ?Bټ�ټ�ټ�ۼy/ݼ�߼�'㼪��%�鼓��`�8����
��Im��:.�������z������ ��
��
����[��LD�����k����m�;���z���
��  �  �a=l=��=r�=�"=��$=��&=�/(=_*)=o�)=��)=ګ)=�f)=_�(=lp(=��'=��&=~&=��$=Ā#=s�!=Lt=��=�6=L�=0= =��=��=�z="C=��=��=uE=g�=M�=��=��==�8=�=`�=�G=��=/�=g%
=��=�s=��=�I=�^==Y=�~=}=�X=#=K�=�%=Gr=͉=~Q=7�=QZ=�q
=�=ia=m��<��<N&�<��<�H�<h�<$i�<;��<���<ܝ�<`��<���<<�<m��<Q!�<�t�<�n�<�r�<�I�<cF�<��<A>�<l��<6�<�	�<��<uӪ<&��<꒢<Ь�<U\�<´�<+Č<���<C.�<ss<�d<�9U<D�C<��0<x�<��<�"�;���;;.�;�.�;:�;ۓ�;bʼ;}t�;7�;�;���;7�h;6;ED5:�+�}���##���;�'+@��66��%�P��T��u�����	 �K�9�=Y��(}�y��p����̾���ֻ������|��L!���1�lKD�R|X�|�m�k���r��� ���s��7"��Yn���!��b�����1���ț��͢��'��T�������5�ɼ�ϼi{ҼoXҼc�ϼ�˼Y�Ƽ���e`���&������'����ܵ��v���]������?���+���s���o���H�������P����ļRDʼG�мM�׼��ݼ� ��G�b�����༃=ڼ�bԼC�ϼ��ͼI6ϼ�ӼF?ڼo�἞c��7＾��3��C�"u�*��T��k�޼�9ۼ��ؼb׼�ּ��ּ�*׼<�׼��ؼڼ��ۼ�Mݼyo߼��YG���C���q��C���l��BO����E	�5N	�b��������M ��:��U����V���s��1��9
����͆��  �  �l=~�=�=��=d�=L#=!x&=m�(=�9*=��*=i�*=�K*=��)=�)=i(=S�'=~Q'=��&=�%=.�$=̼"=��=�6=@�=��=�=I�	=$$=��=�=�	=�o=R*=�U=�(=	=?=|='�
=�M=�q={ =���<� =J<=i�=��
=�=��=7=�~==]4==��=�Y=#=��=��=�G=��=�z=p�=��=�	=0=sH =��<<!�<��<�X�<?B�<��<TX�<���<���<v$�<O]�<y�<ʄ�<�"�<9,�<Q�<�ϧ<I7�<ST�<�P�<��<3�<)ʯ<��<��<TX�<���<���<^]�<�ڝ<�:�<M��<A�<ۏ�<�Ё<�w<�h<�W<U4C<��+<e<jm�;���;I��;�S�;��};;��;�ō;�˝;澪;��;v��;�	�;��9;�H�:Xֹy����N�&��:�ú��*&p��LK�2a&�L�	����q����&��E+��YP�rz�g��uO���_��NKջ��ք�������0�DdF�� _�t�x�@��A���b�������o᥼���7��Ξ������Ӝ����O��p۲�4�B�ʼ��Լ܇ۼWR޼�*ݼ��ؼ�1ҼïʼQ[ü��0�������3r���+���v������������u]��-����]�������ͺ�M���-:ļе˼��Լ��ݼ\�����J��<��m�� ���(ۼ�hռ��Ҽ�%Լ�PټD[����S��"���_���S���̀������`���漦�߼Hiڼ��ּ�ռ޾Լ�Rռbּ�׼��ؼc�ټVۼT"ܼ�ݼu�߼l㼝�&％���� ����
�Fe�n6�G4�u�}j
�����s��8�V� �
<�ۆ��
�q���?��d��  �  �5=�=�d=BZ=n�=�!=	�%=W�(=Uv*=�*+=�+=o*=��)=��(=)(=��'= L'=[�&=j=&=�%=<�"=�=�8=��=��=�C
=	e=b=%� =�=�=��=�=W�=��={�=V�=��=�i=2=nF�<'��<+k�<3u�<�<��=�=�==Y9==��=F~=�x=1=��=5=?�=\�=��=��=�=��=>�=�(=��=^=�L�<\�<��<�z�<�*�<���<BV�<'f�<���<`�<*�<6�<$��<X��<���<���<թ�<O��<7�<�6�<6��<�:�<c]�<O��<�O�<Su�<�#�<#­<���<^]�<M|�<ԫ�<�<�ӌ<���<zD�<�Tx<�ui<��V<��?<�n%<n�<���;��;)t;$�>;ҩ+;��7;6�Z;%�;*�;��;���;9�j;A7;z��9p����EG��ʎ�������ؕ���g��*�t�Ə@�f��*������n���&��
O��F|��k���$������zֻ�&뻹� �h�����$(2�|�J��f�c�����$��m���������.��J����/���¡�if��Y(���-��	����Ƽ�KӼ�s޼�弆�����z)���ؼXϼ�Ƽ	K�������$��:���v���GV��J?��.���~���������+඼ҷ�%��}��A9ż0Aμ��ؼo?�����L���P��M������h����l�YIڼ@2׼O�ؼ�_޼��`=�����P��{��z��h�i{���P�����]�Iۼ[�ּ^Լ�Լ'�Լ�aּY�׼�Xټ}fڼ-ۼ��ۼ��ܼ��޼��gV�g~�����1��	��^��X��k��O�Z&��z��(
��2�k��8��Ӈ��6��M����J��ox��  �  �=+^=�F=��=�=!A =��$=�C(=�[*=;2+=7+=�a*=�w)=��(=o�'=t'=�)'=��&=:G&=�%=��"=�-=DI=^V=��=�=m/=d�<�l�<���<\y==��
=��=�Z=~i=I=I�
=�
=r|�<��<��<`L�<���<_/�<�%=��=r=��=P�=��=)�=]{=F�=�a=��=��=��=��=f�=)=$�=�_=q�=(q=�X=��<�Q�<��<�z�<�5�<cD�<˭�<B��<$�<(��<)�<0K�<m�<��<(	�<���<i�<���<�K�<Kђ<I4�<��<mJ�<�ѫ<CS�<�#�<�,�<-ݭ<��<*�<�
�<!�<���<�m�<�r�<�:�<�Jx<b�h<`AU<��<<� <�� <	y�;��;�
=;��;}��:E-;<"/;[b;�|�;U^�;�8�;�1R;O��:m�S�����qx�򩻆7Ż.H̻/��&���"EV�-w#�W���=���J���&�-P��������Ļ�&ػ^��� �a��f���O4���N�4!m�ź��:����~�����RP��+ٶ��S��13���{���U��ݐ��P?��a���������ʼQټ弡���Ｌ��D缣�ݼ��Ҽȼ}����#���=��B���(����������ꄶ���������ڶ��඼�����2������`sƼ�{м�]ܼ���#���b���V����� �kr�����_ ��ݼZAڼ��ۼ�἟��&M���I����
�j �K��W���������H ��(ܼO�ּ�]Լ�Ӽ[�Լz�ּ�aؼF�ټ��ڼ��ۼtܼ��ܼ.�޼ɽ⼩	�A�Ib��������o����G��Y��XT��8��m���t(��k���
�������5�����  �  �+=�J+=��,=l)/=��1=�4=��6=8=O~8=�8=s7=�5=�l4=�M3=��2=�12=6.2=S2=d2=B2=}-1=Rg/=��,=�9)=#H%=	[!=��=�=�=��=f�=�=��!=��#=f2%=�%=i#=�� =�=�_=9G=I=ٴ=�=Ζ=�_=0i=�1=gP!=��"=��"=}"=��!='� =��=��=`k=�u=�=�(=y\=�=�==Z-=_|=Of=6e=�	=�=?H=�M=�E=U�=��	=�
=%�=QQ=�=]o�<kw�<+��<���<��<�Z�<]��<ha�<^�<��<��<��<�"�<[�<*�<��<�F�<�ʱ<)ԫ<잦< &�<,�<_P�<5�<���<��<ki�<!�q<�d\<��F<�2<kT"<l�<ŧ<^�</�<I�<g\<�I<��<5<<O��;�I�;`��;��E;�Y ;��:q�k:�Th:��:�m�:�:�b�:ZL�:.��:��:��9?����[��n���.�+�	�R�4�t�6����a���H��ğ���޻a� �6�0r+�H�A�~�U�.�e���p��Rv�I�v��at�Q#q�.�o�Dr�#z�����}S���C�����^{��`X��@��ݡ��?���'���<=���������ȗ�0��<�������ٛ�HΝ��7���֟����잼���{���ܝ�����Y��
Ө����>M������u_ļ��Ǽ�ȼ��ƼR�¼�������
������HJ���Y�������ļd̼v�ѼT�Լ�Bռ��Ҽ�lμ��ȼü�0��eں��[�������5��9����6����¼ZPļ�=żDoż�0żd�ļ<ż7�Ƽ�ɼlpμ��Լ^�ܼ���b/���x���T��D�򼆃�]L�ۗ�p�ἶ>ἄ���輟�����m�������  �  u�+=H,= q-=~�/=2h2=��4=�7=[@8=�8=�$8=%7=��5=�4=�{3=
�2=�^2=�S2=�o2=�z2=a/2=�G1=[�/=��,=��)=��%=Q�!=&�=�K=�>=O�=0=2�=)-"=mS$=�z%=xL%=��#=P� =�|=��=�=� =�q=�D=i9=�=��=4{=�!=�"=&�"=6�"=r�!=�� =��=��=��=�=�=�B=3q=$+=d+=E=�q=��=��=v= �
=i9=��=*�=/�=j	=�(
=�]
=?	=k�=e=]'�<-`�<z��<��<xK�<D��<)
�<���<�H�<�J�<���<$Z�<<O�<�|�<<<�<Z�<Ҍ�<�"�<	7�<�<\}�<Ut�<ɋ�<jN�<�7�<�Ҋ<�<�r<;<^<�'I<q�5<8L%<<�<8�<�^<��<�e<�<�m<1�<dR<
$�;�z�;؅�;�>O;�;wx�: �:�y�:�R�:��:���:�� ;�X�:�W�:z�:��9D����4������`(��O���q�Y����j���Y��	���]�ܻN��@���j)�3?�%�R���b���m��{s�rit��Jr��ro��Xn�Eq���x���p����U������*��u欼����O4���I��а��l���|��c���%�����7ؗ�쌙�I���3z���؞��v��rS�����Wҝ��P��v���"x��.����F������{E���D��J�¼	�Ƽ�`Ǽ��ż�n��P)������E��
~��H���⵶�Mм���ü��ʼ�_м�xӼ��Ӽ�Ѽ
8ͼ��Ǽ�[¼����C����$���q���	��fa��<;¼��ü��ļż��ļ��ļ/ż�pƼ�Wɼ�μ;`Լ��ۼ3�����Ji𼯎�u��S��:q�m���1	Ἲ��62�RG�g&２����v���:��  �  �-=	.=�G/=H1=C�3=��5=��7=\�8=K�8=�Q8=G\7=C,6=(�4=�3=�;3=��2=$�2= �2=K�2=^\2=H�1=��/=��-=��*='=��#=� =�V=�L=�=��=� !=�O#=�;%=�@&=�&=��$=��!=��=g�=P�=�=��=�==L�=X=9�=�9 =|�!=��"=%*#=��"=�!=Z !=� =�s=J=�=�?=x�=��=�W=Ol=`�=)#=�=UH=�=o�=?
=��=��=o`	=5]
=�$=i%=w�	=�@=�2=�2�<���<P �<�u�<�;�<��<���<E��<���<<�<���<Q�<��<@��<��<%��<bG�<��<@?�<��<0b�<�*�<;�<�Ö<纑<ُ�<�	�<]uv<c<liO<T =<1y-<"<�<�<��<$G<�<��<ȡ<�M	<L�;܍�;��;�Vj;�z);+i�:��:zs�:pQ�:��:dg; <	;�;-��:��:w��9n���R����库~��8G���j�����"*��BL�������ػ����Ѫ�P$�2U8�D�J�5eZ�Wge�	�k��lm�4tl�@�j���j�L�m��u�a=���|��
����ě�gt��(ר��l���;��|¨��ɤ��:��	���������X��� y������蚼�E۝��w��q��f���hQ��y�@R�������ڦ�Pܬ��v���ҹ� ���c¼�Qü����f5��D���@ڴ��^�������2���ﴼ�����2��ЍǼ �̼?`ϼ��ϼ �ͼU�ɼ�0żYk���f��E���R�����|����ּ��0���P��=�¼��ü�Kļ�PļYOļ��ļ�	Ƽo�ȼj�̼��Ҽ�ټ���@��e�Yl�	��zh�Y��&��hl߼�4߼˛ἢ`����e����������  �  ;�0=��0=��1=|l3=�65=��6=�+8=��8=�8=�d8=�7=��6=X{5=M�4=w�3=�o3=b,3=j3=��2=�m2=:�1=�A0=�@.=ή+=T�(=�%==7#=�H!=
L =�^ =h!=�#=_�$=Ѓ&=P'=Y'=K�%=s#=
� =�=�{=D�=O�=�=�p=cO=*Q= !=�o"=�##=<#=��"=#+"=�c!=�� =� =��=d�=��=�=��=�d=A�=�=*�=Z6=`%=X=�M=�*=r�=1m=s�=R4=��=�9=��
=R-=fR='$�<���<��<=��<s��<5h�<��<g �<�3�<*l�<��<���<���<Q��<'��<&�<�(�<�A�<R��<�\�< ��<A �<���<��< �<�3�<%M�<J�z<
�i<�X<�wG<�19< J.<qX'<k/$<��#<�^$<y$<r� <'m<�a<�p�;���;˒�;�$�;x#V;/6+;�Y;��;�9
;^;Ђ;�;V{;I�:_��:s
:z�.�
:g���Ϻ���<�qa�q���
��ZĦ�%��Mpջ�;󻟌
�����.���?�VON�q!Y�E�_�f c�K�c���c�He�^yi�=�q��}�^}��\䎼���%���$墼
e��&����̣�~Ҡ�1_��J,��Η�}���w���D��˛����<��������)���O���!���֜�ź��./������G?��s-��a'������{���qx��k���b��H���s�������ӱ�����_�Z��p��&f�������¼��Ƽ�eɼ��ɼ<:ȼmIż����󽼴�����f��S���ic��WI��^K���"��|����¼�Bü[�ü��ü��ļ�ż>>ȼ��˼̼м�zּ��ܼ#�~��Oj� ���C��Le��)߼�1ݼ�/ݼ|k߼��㼭F�4M�̾��H����  �  �N4=�-4=��4=��5=�6=��7=0h8=ǰ8=ێ8=�8=�j7=��6=�5=n(5=k�4=�3=ބ3=B3=��2=�2=0P1==+0=J�.="�,=cl*=*,(=$&=[�$=	�#=�#=N$=ey%=��&=�'=Ie(=z(=��&=^%=��"=�� =j�=WZ=�=�/=S=�G=� =C�!="=��"=��"=��"=q""=�!=H !=�� =�Z =� =��=��=w==�H==�q=�Y=��=a�=�M=�s=�*=N}=J=�G=\=�U=ط=�	=�}=0=�<��<9�<ق�<���<��<}��<yr�<CH�<f��<9_�<d�<K	�<8M�<�&�<�Ǻ<�U�<2�<_��< ��<4��<A��<���<���<�	�<]߅<%"~<ϗo<��`<��R<>F<o<<��4<�i0<�.<X,<R�)<�.%<�.<��<��<]q�;���;��;��;�_;OQD;vK4;�+;��&;�} ; ';,�;F�:w/�:$�:-N���FI��|������<1�N�Y�f����������`����Ի�Hﻔ.�����%���3���@�K�s�R�<W��Z��^\�ؑ_� �d�lIm�'�x��/������U���e������呞�aA��ր��;֜�Ϛ������H���!��6�����������f����V��+훼6T��G���>ל��0���ݝ����n,��(��\ȧ��ݫ��᯼�Q��ޭ��ϗ��K������=���}���|��Zݫ�J���Jǯ��ֳ��y���뼼�s����¼�ü�E¼�r��K&��i⻼k���������#����ú��,��1�������]��y���j¼�Bü!ļ� ż�Ƽ�ȼl�˼�Aϼn�Ӽ�Cؼ]�ܼ4<���>l� ��f�༝\޼�#ܼ<�ڼ&ۼ�)ݼ����\��I�J����  �  k�7=�17=q+7=]7=С7=��7=��7=��7=�7=F+7=��6=7e6=��5=b5=9�4=zG4=J�3=%�2=��1=�"1=(H0=wU/=�:.=��,=��+=W*=��(=��'=	'=c�&=�'={�'=c{(=m)='A)=��(=��'=��&=&�$=�#=Ψ!=5� = =T =�O = � =�:!=͟!=B�!=7�!=��!=��!=u�!=�|!=�P!=!=� =�O =C�=m<=Ţ=��=�A=�[=;=��=�K=R�=x=�=�X=tt=��=6=�n=�6=$Z=7�	=�o=��=b)�<@8�<^��<���<G��<���<�p�<ۓ�<���<0��<֕�<���<���<��<�R�<ּ�<��<'Ұ<�x�<`�<H�<���<�'�<�Ï<�k�<���<`�~<�Rs<Z�g<Я\<�_R<\I<t�A<�P<<2�7<��3<��.<B�(<��<��<B<��;X��;�H�;�b�;��;�}r;EZ;� F;�$4;[�!;�^;� �:1��:��a:��9:e/�/�=��"����*�B�V��́�U:��&L���$Ļ�-ڻ/���Y�Z�������(�E�3�(�=��qE���K�ѫP��YU�F�Z�jFa�s�i�|st�7��r��y`�������q��H���w��\��י��u����O昼���(��$k�����G㙼�)��,���� ������nǜ��ŝ��Ξ�M埼a��R���p��9������K�������H������ů�ȭ����Q}��e���?���L��9���ۗ��`���e��?$��4���ؼ�`輼^r��F»�������M���W��m����?����z���ׇ������=����'¼	�ühJż�Ƽ��ȼ�zʼ��̼�#ϼ��Ѽ��Լ��׼�Lڼsܼ��ܼ��ܼx�ۼ��ڼ�zټeټ��ټWXۼ�0޼%��>{�%��g���  �  �C:=Ӊ9=w�8=}E8=�7=�7=�v6=m�5=��5=�|5=�5=��5=T�5=�s5=��4=�.4=�3=��1=o�0=c/=[a.=đ-=��,=eP,=�+=�/+=[�*=� *=��)=�|)=�s)=��)=��)=��)=��)="K)=�(=O�'=Zc&=�<%=94$=�\#=ͷ"=�6"=��!=&]!=�� =� =S@ =�	 =  =/ =N =x� =T!=�!=�� =� =�2=&=.=)#=�U=P�=�=�p=g�=��=N=�=C�=�=��=��=5Z=�=��=��	=%�=%�=�% =	f�<���<4��<	`�<�O�<s��<���<X{�<�!�<���<���<R8�<z��<�U�<���<��<X��<H��<�x�<u��<�o�<N�<C�<���<3>�<�{<�us<Rpk<��c<k�[<�1T<��L<�:F<V�?<Vh9<�w2<��*<(!<�O<r9
<���;T�;�y�;yȱ;^�;�;��s;�R;�3;�;���:�ԫ:��c:�d�9 Nq8�z���[N��ĩ�����z�(���Z�.������ި����ѻ���@��M5��$�%���� ���)��I2��l:���A��I�k P��=W��+_�g
h�|�q��|�5����V���鏼Bǒ�0��^����������������Ԝ�V���c㛼�'��᜚�a�������B��V���蟼�ء�ጣ��䤼�㥼_���-_��V���ʨ�6���L$��a���`����R��\Щ��P��1���k��fi����u/������#ղ�޴����cܷ�M���$�����0���<��
,���ؾ��&�����ܾ������Ⱦ�iu�������¼�-ż_�Ǽ7ʼb̼�*μ ϼQ�м� Ҽ�WӼ:�Լ)�ռ��ּ�}׼\�׼��׼k�׼��׼��׼��ؼ�Qڼ�rܼ��޼I��\�C8��  �   <=|�:=ۦ9=�28=$�6=DH5=�4=�F3=�2=�3=1�3=v=4=��4=��4=h�4=ȟ3=�&2=�^0=+�.=�,=i�+=��*=c�*=�*=��*=�N+=�+=K�+=F�+=@\+=�+=e�*=w*=� *=D�)=�@)=��(=:(=A`'=r�&=��%=C%=�m$=�o#=�E"=�� =&�=S�=˼=�O=�b=��=$�=ܩ=�] =�� =�T =�n=�=�v=q�=;�=H�=�=g�=9=j3=)B=v=��=M�=g�=�1=��=-�=ݮ=]=��	=)=�=�=j/�<15�<�=�<3�<| �<���<:U�<4�<̀�<�w�<�J�<�<�s�<D/�<2��<抴<4E�<A��<�
�<��<��<E��<h+�<TӁ<�G{<��t<�o<�k<��f< ua<�~[<��T<2M<4E<��<<��3<��*<%� <�<7<�, <�f�;&��;�ſ;���;37�;��};�!P;wf";ǚ�:�X�:��):
�\9���ѹ{-��Y~��ߵ������9/�o�f��ɑ��R���̻E��j���]�Z��|��o������#�/y*�ڐ2�s!;���C���L���U���^�X�g�Fq��y�$�����Ϋ�����DG�������㕼:���\��������)�����w���U���}��&��c��盼,���q.���=���@������	Z�����J̪�	���������3���̦�zæ�
����S��ͺ���/������{���k��/���ڬ�K<��ҩ���&���ɲ�s�������)���/s��06�����jiü�Lļ�4ļKü���i���e���XB��]���_ļ��Ǽ�u˼��μ=�ѼΔӼ�xԼ�Լu;Լ��ӼI4Ӽ$Ӽ1Ӽ��Ӽ�`Լ�%ռ��ռ;�ּ)�׼T�ؼ=4ڼ��ۼOݼ��޼"��n��  �  �<=?l;="y9=�;7=m�4=J�2=�1=D�/=��/=,10= 81=du2=]�3=�4=`�3=B�2=8�0=�u.=�	,=��)=zf(=ߪ'=�'=VZ(=�`)=߅*=��+=y=,=�,=Ie,=��+=[X+=K�*=�)=�])=f�(=�l(=@(=��'=�r'=��&=�G&=i4%=̵#=E�!=�=�=\�=v�=�=�>=!0=��==�@=��=C�=![=̆=�V=�+=�b=�?=��=� =�=��=ը=�0=\4=�=�x=;�=��=��=nH=��=5>	=m�=�=zs=��<���< ��<�)�<���<� �<]�<}e�<Ɂ�<Qο<��<�Ӹ<	<�<+,�<�<���<#®<��<Hˡ<4[�<6��<r/�<k �<b�v<!fo<�j<M�h<D5g<�e<�Ic<J_<��X<5Q<��G<\�=<a�3<)<j�<�Y</n
<}� <ډ�;�M�;K�;tΰ;��;�\y;�4?;�;�O�:�0�9��'�WF�KY���}�0d��fF����κ�a
��<���y�,�����»�M������	��y����Rw�>���M��e ��V&�T.��H7��]A��K��'V��`��ci�u�q�y�7?���u��䙆��뉼'���E쑼����ज़�e��r��8S������pN��!w���������9���	��T�������=���t��ך���Pﰼ�[��1Y��SI��V��� ��V˦��U��H���1�������[֦����9���H��.��t꫼����9-��?󭼱���ڰ��m��W߶�$��{����ü�iǼg�ɼ��ʼ�BʼviȼL�żü���������~üO�Ƽ�3˼rмk�Լ�ؼx)ڼ��ڼ��ټ��׼D�ռ�ӼM3ҼF|Ѽ�Ѽ?vҼ��Ӽ�Nռx�ּ�_ؼf�ټM�ڼ�ۼi�ܼ9�ݼ��޼�Z��  �  �==�(;=�8= �5=��2=�/=��-=j�,=g,=8-=�.=�0=�2=��2=I�2=�1=�A/=]i,=;q)=�&=�
%=QC$=M�$=�%=�J'=�$)=Y�*=c,=j�,=��,=�=,=&k+=�w*=��)=��(=�8(=��'=,�'=�'=��'=eS'=ޑ&=�;%=�D#=�� =��=�9=S�=�>=*�=�=�]=�I=+P=��=��=�u=�=��=)=qc=�-=��=.v=	=�J=�=,q=ݚ=]=$�=Q�=.�=*�=�A=�=�=C}=m=Բ=�X=B��<�T�<�	�<��<�O�<-�<?��<���<{
�<N۸<���<X�<ر<4�<(��<(9�<�Ƭ<�<f#�<IǕ<<�<��<�>u<ͤi<N�b<��_<�_<��`<�Ob<�)b<��_<�;Z<�QR<zsH<;k=<R�1<��&<�<g�<�<=��;���;���;&��;!�;|*�;�sj;8r%;ҷ�:z��9r����؂�n����(˺��̺	ɺ�Ϻ�J�T��<�L���������Cֻd���5�R��@���(�$Z�Ź����i� �>%��v,���5���@�!WL���W�wGb�R�k�!�s���z�A��*����ۅ�<D��.���˼��Ø��$�� B���i�����t��T�������=��'��5ՠ��$��Ϛ��@��s����꫼p"���P��Ｗ�����s��hU��Xa��dP���ͧ��\���5���G��/L��\ܦ�H����8������c��hԬ���������m���g���e��~���r%��0����ü/ɼ��ͼ��мڙѼ(zм�ͼ�ʼ,�ƼuXļv�ü��ż�ɼ�μf�Լ�uڼ��޼����3�D�߼(�ܼ ټ��ռ��Ҽ&FѼ��мW�Ѽ�wӼ��ռ;�׼�zټ��ڼ ܼ
�ܼݼJlݼ�.޼o�߼�  �  ��<=ۊ:=��7=�4=�0=�N-=��*=w�)=م)=@�*=֔,=��.=�0=2�1=l�1=�_0=��-=�*=�.'=�0$=U"=�B!=o�!=F#=�<%=�'=�)=�+=,=�,=(,=9+=�*=n)=h#(=��'=�R'=�V'=�x'=|�'=�B'=�m&=��$=Ɂ"=y�=�)=��=� =�F=ڝ=�9=��=tF=��=�=��=�l=��=G=M=d�=	f=D�=�t=�:=��=�=�=��=�=��=��=��=qg=μ=��=�C
=��=�f=4=�=�_�<��<q�<&��<M�<-�<ث�<���<;�<���<R��<p�<?+�<�%�<�Ǯ<�<̪<m��<ʣ�<䎒<�̇<�.{<uj<_�]<8!W<�9U<��V<�eZ<u�]<8�_<Zi^<6�Y<CR<��G<�<<��/<�#<��<��<�<<�t�;���;��;d�;�P�;-��;�X;Q�
;�q:F8�6R���<�i�����	�����il��Ѽ��x'���\�Fq��XH���Z�g�@G� "�7�'���(��<'�'u$��f"�\�"�B�%�٘,�F6�uA���M��Y��d��1n� �u�B?|�����-����|���5��E4��>=��?���䩼 ݯ�T᳼�f��YM�������@���L��3K���7��e�������	���W֯�Tﵼ�׺������	��� ��f���!�������m��s.������j��.���R[��1p���\���Ӭ������魼F�������ݜ������B̰�ٝ������
����}ǼFμ�_Ӽ��ּ�|׼��ռBUҼh�ͼ��ɼD�Ƽ��ż'�Ǽn)̼�FҼq ټx�߼�f������d��Cἱjܼ-�׼@+Լ��Ѽ`4ѼZ�Ѽ=�Ӽ�ּG�ؼk�ڼ�Jܼ�;ݼ
�ݼ��ݼ�ݼ�S޼��߼�  �  J{<=��9=�6=t�2=��.=9t+=��(=J�'=Ï'=��(=�+=M�-=��/=s1=�1=x�/=$�,=�Z)=j�%=�c"=� =Y1=��=�L!=)�#=h}&=~)=�+=1,=�u,=��+=��*=�)=y�(=Ԧ'=n'=k�&=�&=�4'=U'=�'=/&=�s$=��!=`�=V�=7=�3=8=��=	S=B=6�=y�=��=�=ê=� =$5=��=�V=ɂ=:�=�`=dC=�"=]�=� =��=Q$=j?=Q=V�=�=fR=2u=�	=�,=��=��=4� =w��<�y�< ��<qx�<���<'��<_��<�&�<+1�<���<�<�R�<��<ɔ�<���<�N�<NV�<�t�<�ݚ<�S�<� �<Hwt<�~b<��U<DO<��M<��P<�iU<GZ<�@]<��\<��X<�KQ<J�F<��:<�=.<��!<5�<!�<y<���;��;f��;0Y�;�E�;�;��I;�
�:�:�%��cϺ����(�M9*�^��2���
���8o2���h�!ř�2�Ż��Q�U���*��s/�U�/�#-���(��u%���$�'��J-���6�IB���N�:[���f��p�"�w�)�}��:�������@������{���a}��>/���d��W7����������y��q���F�������z��������F*���^���ѫ�G���e0��t���.���}(¼�俼%���3浼����Ъ�d
��!��Ǥ�p奼jާ�I%���@���ҭ����YĮ��i���������[﮼�_�� ���k����¼�iʼߛѼW׼��ڼ��ۼ��ټ{vռ�dмȘ˼�Lȼ#kǼ[_ɼ�ͼ�Լ��ۼ6��I輷�&����C�k�޼�ټ�\ռ4�Ҽi�ѼPҼE-Լ��ּMRټl�ۼ�KݼY/޼�g޼B޼�,޼L�޼�Q��  �   V<=��9=ZU6=+b2=].=��*=�!(=��&=��&=�F(=$�*=7-=;y/=��0=W�0=�C/=��,=-�(=�%=_�!=%j=\t=��=z� =�0#=B&=k�(=��*=R,='^,=��+=)�*=�)=�q(=�w'=C�&=��&=��&=D'=+?'=U�&=&=�H$=��!=f%=�R=K�=]�=/|=)�=��=�=k=�?=��=�=c=Ѱ=s�=1M=��=��=�=Т=e�=+�=�=$�=��=��=�=	7=i=D�={*=E=�}	=a�=l�=}�=� =��<
F�<{�<��<H�<��<��<�ܼ<�³<�</�<��<��<���<�	�<L��<�˨<Q�<�8�<x��<"�<�r<l�_<d�R<�5L<�!K<�:N<��S<.�X<MK\<�U\<yX<��P<�F<�`:<��-<�1!<@�<G+<M�<���;���;]-�;���;m�;��;]D;���:;T�9N�O��m��C��3���3�ï'������Q��`�6�C:m��m����Ȼ63������!���,��G2��v2�6/��*���&��P%���'���-�&
7�;�B��SO���[�"Dg���p�.gx��.~��o��)���i���%��tN�������ꝼ`���l�����Gp��b�Mo���q��'���tA��鬥��K��ϸ���������|u���V���쿼�2üܡüK��7¼��궼�Ȱ��Y���d���E���򤼃�����k��ޖ���2�����6��ث��a.��F#�������_������üx{˼��Ҽ��ؼ�Eܼ[�ܼ��ڼv�ּ�KѼR̼z�ȼ��ǼB�ɼ�μTeռZݼ.�֩�d�������Ho��߼Y_ڼ��ռO�ҼC�Ѽ1zҼ�ZԼ�ּ�ټ��ۼ��ݼ��޼��޼I~޼<[޼*�޼����  �  J{<=��9=�6=t�2=��.=9t+=��(=J�'=Ï'=��(=�+=M�-=��/=s1=�1=x�/=$�,=�Z)=j�%=�c"=� =Y1=��=�L!=)�#=h}&=~)=�+=1,=�u,=��+=��*=�)=y�(=Ԧ'=n'=k�&=�&=�4'=U'=�'=/&=�s$=��!=`�=V�=7=�3=8=��=S=B=4�=w�=��=�=��=� =5=��=�V=��=(�=�`=MC=�"=C�=� =��=J$=z?=�Q=ʃ=�=�S=�v=�	=�/=�=�=� =0��<̅�<���<���<���<���<���<�4�<�>�<M��<���<]�<�
�<���<�Ƭ<kQ�<�V�<�r�<�ٚ<�M�<��<Mdt<�hb<��U<�O<9�M<vP<#MU<+Z<#&]<��\<��X<�7Q<��F<��:<�4.<�!<ظ<�<��<S��;O��;��;���;Dx�;(�;PJ;���:��:��#��κ�:�p�'���)��Y��j�*m
�w��p2���h��י�u�Ż�)�f�Z�l4*�|�/�?0��)-��)�B�%��$�)'��d-���6�h^B�@�N�J[���f��)p��w�(�}�I=������;B����>����}���/��Ee���7������<��� z������F�������z��#������J*���^���ѫ�H���f0��t���/���~(¼�俼%���3浼����Ъ�d
��"��Ǥ�p奼jާ�I%���@���ҭ����YĮ��i���������[﮼�_�� ���k����¼�iʼߛѼW׼��ڼ��ۼ��ټ{vռ�dмȘ˼�Lȼ#kǼ[_ɼ�ͼ�Լ��ۼ6��I輷�&����C�k�޼�ټ�\ռ4�Ҽi�ѼPҼE-Լ��ּMRټl�ۼ�KݼY/޼�g޼B޼�,޼L�޼�Q��  �  ��<=ۊ:=��7=�4=�0=�N-=��*=w�)=م)=@�*=֔,=��.=�0=2�1=l�1=�_0=��-=�*=�.'=�0$=U"=�B!=o�!=F#=�<%=�'=�)=�+=,=�,=(,=9+=�*=n)=h#(=��'=�R'=�V'=�x'=|�'=�B'=�m&=��$=Ɂ"=y�=�)=��=� =�F=؝=�9=��=pF=��=�=��=�l=��=G=9=K�=�e="�=et=T:=��=��=a=��=�=��=�=��=�h=�=�=�G
=a�=>m=�;=�=�t�<��<҉�<V��<Oh�<�:�<���<���<8U�</ֲ<�Ǯ<;�<�;�<�2�<eѮ<|��<<ͪ<E�<p��<���<���<�	{<�i<#�]<6�V<�U<��V<�.Z<R�]<Qg_<�8^<&�Y<��Q<��G<� <<��/<��#<��<�<�L<���;/��;��;���;��;��;��X;�n;ku:�s*�J������\�}��g ���������>��p{'��]������|��|�绑���u�TK"�b�'��$)�
x'�Ű$�E�"�:�"�K%&�:�,�TD6�F�A�+�M�
�Y��d�{Gn�nv��L|�)����1�����~��7��`5��>��߻���䩼{ݯ��᳼ g���M�������@���L��@K���7��l����������[֯�Wﵼ�׺������	��� ��g���!�������m��s.������j��.���R[��1p���\���Ӭ������魼F�������ݜ������B̰�ٝ������
����}ǼFμ�_Ӽ��ּ�|׼��ռBUҼh�ͼ��ɼD�Ƽ��ż'�Ǽn)̼�FҼq ټx�߼�f������d��Cἱjܼ-�׼@+Լ��Ѽ`4ѼZ�Ѽ=�Ӽ�ּG�ؼk�ڼ�Jܼ�;ݼ
�ݼ��ݼ�ݼ�S޼��߼�  �  �==�(;=�8= �5=��2=�/=��-=j�,=g,=8-=�.=�0=�2=��2=I�2=�1=�A/=]i,=;q)=�&=�
%=PC$=M�$=�%=�J'=�$)=Y�*=c,=j�,=��,=�=,=&k+=�w*=��)=��(=�8(=��'=+�'=�'=��'=dS'=ޑ&=�;%=�D#=�� =��=�9=R�=�>='�=�=�]=�I=$P=��=��=�u=�=��==Oc=�-=��=�u=�=�J=��=�p=��=S=_�=��=z�=R�=1E=k�=�=�=�=�=�e=���<9u�<�,�<��<{v�<RT�<���<7	�<�/�<��<iδ<N��<��<���<x��<�@�<Ȭ<� �<�<X��<ϋ</l�<�u<�ai<Ub<�Y_<J_<��`<	b<�a<Q_<{�Y<YR<�EH<�G=<��1<߂&<�<H�<-�<���;C�;iK�;0F�;ަ�;վ�;��k;P�&;F7�:(� :�0��=���	����rɺ�}˺.Ⱥ)Ϻ~��@����L��E�����9�ֻ�����O����Y��uz�+��7����!���%��,��-6�YA�e�L��W��lb���k���s�ίz�sH������߅�0G��X���c���IĘ��%���B��Ij��~���ht����������=��$'��Hՠ��$��ښ��@��y����꫼t"���P��񼷼����s��iU��Ya��eP���ͧ��\���5���G��/L��]ܦ�H����8������c��hԬ���������m���g���e��~���r%��0����ü/ɼ��ͼ��мڙѼ(zм�ͼ�ʼ,�ƼuXļv�ü��ż�ɼ�μf�Լ�uڼ��޼����3�D�߼(�ܼ ټ��ռ��Ҽ&FѼ��мW�Ѽ�wӼ��ռ;�׼�zټ��ڼ ܼ
�ܼݼJlݼ�.޼o�߼�  �  �<=?l;="y9=�;7=m�4=J�2=�1=D�/=��/=,10= 81=du2=]�3=�4=`�3=B�2=8�0=�u.=�	,=��)=zf(=ߪ'=�'=VZ(=�`)=߅*=��+=y=,=�,=Ie,=��+=[X+=K�*=�)=�])=f�(=�l(=?(=��'=�r'=��&=�G&=h4%=̵#=D�!=�=�=Z�=t�=�=�>=0=��=v=�@=��=0�=
[=��=�V=�+=�b=N?=}�=� =,�=k�=��=�0=X4=j�=�y=��=��=��=N=�=�G	=�=�=\�=��<8�<�<]W�<��<91�<�<�<ٔ�<@��<���<߹�<��<�X�<�B�<7�<ǡ�<Į<d�<���<�G�<hr�<��<�ۀ<��v<�o<�j<�+h<U�f<�ke<��b<��^<:�X<S�P<ӮG<�=<~n3<U�(<1�<+g<��
<�� <k��;���;`��;hw�;弘;��z;b�@;5*;`O�:���9^�dv�*U�dz�f���a���eκOf
��B<�*lz�Z���E@ûq�㻞$��
�	�>��).�d�������� ���&��o.���7�i�A��L��]V�GG`��i���q�n�y�KH���|��󞆼Dߨ��F(��������e���r���S��쨨��N��Ww��?������49���	��b�������=���t��ܚ���Sﰼ�[��3Y��TI��W���!��W˦��U��H���1�������[֦����9���H��.��t꫼����9-��?󭼱���ڰ��m��W߶�$��{����ü�iǼg�ɼ��ʼ�BʼviȼL�żü���������~üO�Ƽ�3˼rмk�Լ�ؼx)ڼ��ڼ��ټ��׼D�ռ�ӼM3ҼF|Ѽ�Ѽ?vҼ��Ӽ�Nռx�ּ�_ؼf�ټM�ڼ�ۼi�ܼ9�ݼ��޼�Z��  �   <=|�:=ۦ9=�28=$�6=DH5=�4=�F3=�2=�3=1�3=v=4=��4=��4=h�4=ȟ3=�&2=�^0=+�.=�,=i�+=��*=c�*=�*=��*=�N+=�+=K�+=F�+=@\+=�+=e�*=w*=� *=C�)=�@)=��(=:(=@`'=r�&=��%=C%=�m$=�o#=�E"=�� =$�=Q�=ȼ=�O=�b=��=�=ҩ=�] =y� =�T =|n=�=�v=B�=�=�=<=�=�=3=�A=A=��=��=o�=n3=˗=��=�=Ye=	�	==�(=�+=W�<a�<�m�<�e�<S5�<p��<!��<[i�<���<V��<�u�<+�<ۓ�<�H�<*ɷ<��<]G�<P��<��<z��<+ה<��<��<���<9�z< lt<Y?o<ӳj<y(f<-a<� [<BYT<l�L<��D<z�<<y�3<	x*<Ƒ <w%<	V<D[ <���;Pv�;~o�;]t�;��;��;��Q;K$;���: ��:7�/:�r9,{�K ʹ�$*��^|��d��B�����/�/�g��-�� ԰�A�ͻ:��}0��Y��x`��
�-l����#���*�u�2��z;�p>D�M�V��_�I#h�(q���y�R.������������dJ��􍒼N啼R;���]�����"������������U���}��@��.c��盼7���z.���=���@������Z�����L̪� 	���������3���̦�zæ�����S��ͺ���/������{���k��/���ڬ�K<��ҩ���&���ɲ�s�������)���/s��06�����jiü�Lļ�4ļKü���i���e���XB��]���_ļ��Ǽ�u˼��μ=�ѼΔӼ�xԼ�Լu;Լ��ӼI4Ӽ$Ӽ1Ӽ��Ӽ�`Լ�%ռ��ռ;�ּ)�׼T�ؼ=4ڼ��ۼOݼ��޼"��n��  �  �C:=Ӊ9=w�8=}E8=�7=�7=�v6=m�5=��5=�|5=�5=��5=T�5=�s5=��4=�.4=�3=��1=o�0=c/=[a.=đ-=��,=eP,=�+=�/+=[�*=� *=��)=�|)=�s)=��)=��)=��)=��)="K)=�(=O�'=Zc&=�<%=94$=�\#=̷"=�6"=��!=$]!=�� =� =P@ =�	 =� =/ =F =m� =F!=�!=m� =� =�2=X&=�=�"=ZU=�=a=dp=�=3�==�=��=,�=��=�=�^=��=*�=�	
=z=�=�7 =���<�
�<��<���<���<H��<d'�<��<V�<��<��<�_�<���<p�<FϹ<���<���<(��<4j�<:�<7R�<���<��<�͆<$�<�S{<?s<Jk<�$c<�a[<R�S<k�L<`�E<ȓ?<#69<
U2<hp*<�&!<m_<�Y
<�:�;��;b�;�x�;�!�;迋;�\u;&�T;��4;JX;k�:D�:�Qi:=�9�i�8�e��QL��E�������=)��B[��燻�,���I���zһ$��;���\��כ�v�O!�v*�w�2���:�]TB�w`I�.IP�t|W��`_��5h���q��9|��?��,�� \��2�ʒ����/���]����𙼻���������S՜������㛼(������v�������B��_���
蟼�ء�匣��䤼�㥼`���._��W���ʨ�6���L$��a���`����R��\Щ��P��1���k��fi����u/������#ղ�޴����cܷ�M���$�����0���<��
,���ؾ��&�����ܾ������Ⱦ�iu�������¼�-ż_�Ǽ7ʼb̼�*μ ϼQ�м� Ҽ�WӼ:�Լ)�ռ��ּ�}׼\�׼��׼k�׼��׼��׼��ؼ�Qڼ�rܼ��޼I��\�C8��  �  k�7=�17=q+7=]7=С7=��7=��7=��7=�7=F+7=��6=7e6=��5=b5=9�4=zG4=J�3=%�2=��1=�"1=(H0=wU/=�:.=��,=��+=W*=��(=��'=	'=c�&=�'={�'=c{(=m)='A)=��(=��'=��&=&�$=�#=Ψ!=4� = =T =~O =�� =�:!=˟!=>�!=3�!=��!=�!=m�!=�|!=�P!=!=ӽ =�O =$�=G<=��=��=�A=�[=�:=H�=UK=�=N=-�=6Y=�u=��=<9=;s=G==sb=��	=�|=��=�L�<s`�<�"�<���<5��<���<���<���<��<��<8��<��<��<���<�k�<�κ<��<K԰<�r�<�ޥ<�2�<#��<��<��<>�<_΄<�h~<(�r<"fg<zF\<��Q<��H<˩A<�<<��7<�3<M�.<��(<��<��<Aa<$?�;5�;7ܶ;��;�͉;�t;��[;L�G;�5;A#;�;��:]�:�f:���9��#�ͼ;�V�������N*�)W�41�����`箻U�Ļv�ڻY�����m��c�:P)��V4�?�=�i�E��K���P�=�U���Z��ya��j���t��D���|��oh������Vv�����Mz��(���Aٙ��v������昼���O)��ck��5���j㙼�)��@���� ��᛼vǜ��ŝ��Ξ�Q埼d��T���p��;������L�������H������ů�ȭ����Q}��e���?���L��9���ۗ��`���e��?$��4���ؼ�`輼^r��F»�������M���W��m����?����z���ׇ������=����'¼	�ühJż�Ƽ��ȼ�zʼ��̼�#ϼ��Ѽ��Լ��׼�Lڼsܼ��ܼ��ܼx�ۼ��ڼ�zټeټ��ټWXۼ�0޼%��>{�%��g���  �  �N4=�-4=��4=��5=�6=��7=0h8=ǰ8=ێ8=�8=�j7=��6=�5=n(5=k�4=�3=ބ3=B3=��2=�2=0P1==+0=J�.="�,=cl*=*,(=$&=[�$=	�#=�#=N$=ey%=��&=�'=Ie(=z(=��&=^%=��"=�� =j�=VZ=�=�/=R=�G=� =A�!=��"=��"=��"=�"=i""=�!== !=� =nZ =k =e�=׷=�v=�=PH=�=�q=uY=J�="�=�M=�s=O+=X~=�K=�J=w=R[=O�=7	=.�=�==>�<�3�<)�<���<^��<���<���<���<�w�<���<���<F�<G+�<�i�<N=�<�׺<�^�<�<��<�t�<q�<���<B��<
t�<#�<J��<I�}<O8o<�x`<�dR<��E<��;<ʎ4<a&0<k�-<2,,<�)<�%<�-<7�<�</��;x�;w��;�@�;�;a;��E;n�5;�y-;[V(;K�!;e�;��;R��:C�:�:�O�J�G����e���|1��Z��߀�ކ������� ���ջ��В�����%�34�6A�izK�V�R�{�W�ZZ��\�a�_�e�Qom���x��;��(�������ְ�����甞��C��|���uל��Ϛ��	������)"��o�������У��~����V��8훼AT��N���Cל��0���ݝ����p,��*��]ȧ��ݫ��᯼�Q��߭��ϗ��K������=���}���|��Zݫ�J���Jǯ��ֳ��y���뼼�s����¼�ü�E¼�r��K&��i⻼k���������#����ú��,��1�������]��y���j¼�Bü!ļ� ż�Ƽ�ȼl�˼�Aϼn�Ӽ�Cؼ]�ܼ4<���>l� ��f�༝\޼�#ܼ<�ڼ&ۼ�)ݼ����\��I�J����  �  ;�0=��0=��1=|l3=�65=��6=�+8=��8=�8=�d8=�7=��6=X{5=M�4=w�3=�o3=b,3=j3=��2=�m2=:�1=�A0=�@.=ή+=T�(=�%==7#=�H!=
L =�^ =h!=�#=_�$=Ѓ&=P'=Y'=K�%=s#=
� =�=�{=C�=O�=�=�p=bO=(Q=�!=�o"=�##=<#=��"=+"=�c!=w� =� =x�=R�=ަ=�=��=�d=�=�=��=6=#%=&=�M=+=��=n=�=�6=��=S>=��
=5=�[=�:�<���<o��<���<��<w��<��<�G�<[�<���<�8�<L��<~��<��<{��<�*�<�5�<I�<ᝮ<>X�<|�<��<���<0��<?�<M�<9)�<�{z<4@i<r�W<�*G<��8<�.<�'<X�#<}�#<�:$<��#<E� <l<m<؞�;c �;�;J��;bW;TK,;��;5
;y;�Z;��;/H;$�;o<�:>�:b�:�8&��e��xϺ�+:<���a�ǹ�� i���5��T���� ֻm��P�
���kI/�C=@�R�N�pnY�9`�%bc�Md��,d��te���i�>�q���}�E���쎼���� ��袼�g������Σ��Ӡ��_���,��yΗ�ϑ��Jw���D���3��P��������)���O���!���֜�ɺ��1/������I?��t-��b'������{���qx��k���b��H���s�������ӱ�����_�Z��p��&f�������¼��Ƽ�eɼ��ɼ=:ȼmIż����󽼴�����f��S���ic��WI��^K���"��|����¼�Bü[�ü��ü��ļ�ż>>ȼ��˼̼м�zּ��ܼ#�~��Oj� ���C��Le��)߼�1ݼ�/ݼ|k߼��㼭F�4M�̾��H����  �  �-=	.=�G/=H1=C�3=��5=��7=\�8=K�8=�Q8=G\7=C,6=(�4=�3=�;3=��2=$�2= �2=K�2=^\2=H�1=��/=��-=��*='=��#=� =�V=�L=�=��=� !=�O#=�;%=�@&=�&=��$=��!=��=g�=O�=�=��=�==L�=X=8�=�9 =z�!=��"="*#=��"=��!=U !=� =ys=?=�=�?=d�=��=�W=.l=;�= #=��=+H=]�=`�= ?
=��=>�=~a	=�^
=Q'=�(=��	=oF=�9=�B�<P�<<�<���<�T�<E��<���<��<���<i9�<���<�%�<V��<���<m��<!��<�P�<��<Y@�<��<[�<��<}�<۱�<॑<dx�<���<�?v<)�b<&2O<��<<�D-<%�!<�g<m<�<�-<ŀ<��<�<�U	<�l�;���;��;��j;�+*;���:Qa�:�,�:n�:���:�C; 
;]m;�:D?�:���9.����Є�а�I���]G��j�򅻙l��d����j���]ٻE��|���<$��8�M6K�o�Z�ǝe���k��m��l��j�a�j���m��u�;F�����������ț��w���٨�Tn���<��vè�Eʤ�D;��q�������������By������蚼����O۝�x��q��j���kQ��|�BR�������ڦ�Qܬ��v���ҹ� ���c¼�Qü����f5��D���@ڴ��^�������2���ﴼ�����2��ЍǼ �̼?`ϼ��ϼ �ͼU�ɼ�0żYk���f��E���R�����|����ּ��0���P��=�¼��ü�Kļ�PļYOļ��ļ�	Ƽo�ȼj�̼��Ҽ�ټ���@��e�Yl�	��zh�Y��&��hl߼�4߼˛ἢ`����e����������  �  u�+=H,= q-=~�/=2h2=��4=�7=[@8=�8=�$8=%7=��5=�4=�{3=
�2=�^2=�S2=�o2=�z2=a/2=�G1=[�/=��,=��)=��%=Q�!=&�=�K=�>=O�=0=2�=)-"=mS$=�z%=xL%=��#=P� =�|=��=�=� =�q=�D=h9=�=��=3{=�!=�"=%�"=4�"=p�!=}� =��=��=�=�=�=�B=&q=+=S+=E=�q=��=��=e=��
=t9=!�=|�=��=C	=�)
=`_
=MA	=E�=�h=�/�<�i�<R��<���<XX�<���<I�<��<�V�<�X�<���<�f�<�Z�<���<�D�<�<���<�%�<�7�<v��<�y�<�n�<)��<E�<�,�<{Ɗ<�Ԃ<o�r<�^<�
I<Tx5<71%<�<7s<�J<ҭ<�X<͵<�h<��<�V<!5�;��;Ԧ�;=�O;hg;)C�:���:�]�:�;�:���:#��:.N;+#�:#�:��:�9�e���񒺱y��Fb(��O�r�浈����@��������ܻW����F�)�2?���R���b���m��s���t��`r���o�Oin�!q���x�/�������X��M���2,���笼�����4��xJ��1���Jl���|������D���-��Hؗ�����S���;z���؞��v��vS�����Xҝ��P��w���#x��/����F������{E���D��J�¼	�Ƽ�`Ǽ��ż�n��P)������E��
~��H���⵶�Mм���ü��ʼ�_м�xӼ��Ӽ�Ѽ
8ͼ��Ǽ�[¼����C����$���q���	��fa��<;¼��ü��ļż��ļ��ļ/ż�pƼ�Wɼ�μ;`Լ��ۼ3�����Ji𼯎�u��S��:q�m���1	Ἲ��62�RG�g&２����v���:��  �  ��<=ױ<='G==�Y>=��?=³@=�ZA=	hA=��@=��?=�W>=��<=eZ;=0:=k9=9=�9=�c9=��9=o�9=�9=��8=��7=	�5=03=9�0=��.=M�,=3,=,=��,=��-=�R/=yh0=��0=y�0=�h/=��-=<+=�(=��&=�%=%=�\%=�P&=�'=�)=�D*=��*=��*=�q*=nr)=�-(=P�&=Ӷ%=��$=	y$=Tw$=�$=�G%={�%=��%=1�%=�$=�#=6� =�7=d�=�#=8=�=�N=�-=�@=�&==N�=��==��=�q=d =*"�<��<��<,�<X��<#��<���<��<|:�<�-�<��<x��<c�<�I�<�ؾ<c�<#�<Nد<eG�<�
�<K��<��<9T�<\��<���<�r�<���<�wt<�{g<R:]<�V<%�Q<��O<�{N<ZL<��G<�[@<�5<��&<<�<!H�;ʲ�;�¸;Vܪ;."�;᭟;��;���;U�;���;�$o;þC;��;���:)�:�� �cW��o���#��e���C/�P�J�6rk��ቻ�����t��)5߻�x��������#�%�M�,�4�0�y03��4�_�7�zk<��ID��;O�^�\�v"k�Ly�����4F���ቼw����ĉ�釼�����߃�zꂼB��AT��9m��R�������獼{}���;��~!���W��,0�����Z}��8̌��H��	��Yޔ��P��ٷ��;k���᣼iȤ����	���A��J�������G��r坼��������A��$ꮼ&��P����հ�	Ȯ�V(��Q���Tا��2��^Ч�(���������j��(���
J��l8��N[��X趼�9�����,쵼������  ��@����Ƽ�V˼ϼ|Ѽ�<Ҽ
kѼalϼ6�̼k�ʼnɼR�ɼ!�˼�Lϼt�Ӽ��ؼ{�ݼ����  �  �>==$==��==��>=��?=��@=E�A=�A=��@=��?=�y>=@�<=;=�a:=�9= D9=�G9=׉9=R�9=�9=D�9=�9=�7=��5=�{3=C1=!�.=4d-=��,=t,=�-=�A.=��/=ݏ0=�1=)�0=�/=��-=�z+=�5)=�G'=��%=~%=��%=O�&=��'=�Z)=Qv*={+=�+=��*=�)=oQ(=�'=��%=�%=Z�$=��$=��$=�k%=�%=K&=Y�%=o�$=�6#=�!=؆=��=i�=3�=U=��=.z=�|=�R=t�=�=��=z4=�	=Ϯ=�Q =���<ރ�<r��<	��<"/�<N�<z�<BJ�<�s�<�^�<� �<��<�W�<���<�9�<�s�<�s�<
:�<z��<�X�<��<+4�<��<��<�j�<�	�<�`�<�v<9i<��^<�W<�WS<�Q<_iO<#M< vH<��@<N�5<�B'<(�<��<���;1��;��;��;i�;�?�;���;���;Zy�;q�;�p;�}E;?�;/��:J):|�ظW�I�$���Y�����,��H��9i�������8h���ܻ�k���&����2$�rD+��/�a2�o�3���6�j�;���C�٩N���[��!j�Cx�Q���t�����Ɖ�q���A��1��8{��#����؂����S/��U����O�����z��@֏�&�D��L獼J׌�$E�������� ���^����������$����	�������U��Hh���������>��]����ښ�\���񔡼�+������'���R��7谼����������)���~���寮M���^U���ޫ�Qͮ�I���$��u䵼�Զ�b�����������~���N���6ܶ��1��۵��i&��k�ż4�ʼ^Eμ��м2qѼ��м�μ't̼�Tʼ/-ɼ�~ɼ�y˼��μ
Ӽ�]ؼC�ܼL+��  �  m>=/I>=��>=��?=�@=�yA=5�A=�A=�6A=)@=J�>=^==�<=��:=�,:=j�9=��9=4�9=,:=,D:=�:=�T9=8=Y^6="G4=�2=�0=y�.=I�-=k�-=�.=�/=0=��0=�Q1=k�0=�/=y6.=d(,=�*=�N(=�!'=��&=Q�&=�'={�(=l
*=M�*=�n+=�_+=��*=��)=ح(=�v'=�g&=��%=�8%=�)%=qe%=R�%=�$&=C&=��%=%=�#=6�!=�\=��=�=s�=7r=C�=�P=�#=*�=��=P=��=��=%�	=H[=�,=^��<��<�(�<q�<��<��<�.�<E�<O�<���<
��<��<��<Չ�<qI�<���<���<�E�<戭<q�<��<�Т<�G�<n��<"��<<�J�<(�z<en<��c<tI\<�[W<OT<��Q<>�N<ԲI<?�A<�6<��(<�)<x�<�>�;��;���;���;�e�;�i�;���;���;Rw�;���;�t;P�I;�B;.g�:�J:��8�D#������ݺƍ�F�&��C��c�ɞ�����Y"����ջ�5����h*�0Z���&�z�+��.�e�1�F5�I�:���B��.M���Y��^g���t�����&������s��$熼�{��΃��w���恼�G������y��������m��Y������������������X)���;��I�����!Q��{����	�������뚼P��P���Ϊ���?��\���[�����R���'��C��Μ� x��Y���B¨����'���<���Pȭ�����멼]맼%���*J������ʨ��<������°�����ƴ� ����������	D����e.���G��1m��ǡ������,&ļ3kȼX�˼DGμ�2ϼӹμ�0ͼ.˼�gɼR�ȼ�ȼz�ʼ�μ�CҼ��ּ<�ڼ��ݼ�  �  )&@=��?=�J@=��@=��A=�*B=�[B==B=�vA=t@=7?=��=={�<=z�;=��:=�:=wg:=�q:=��:=��:=rH:=B�9=��8=�7=*V5=�p3=�1=�G0=�g/=3"/=_l/=�0=��0=C�1=߲1=�Q1=�Y0=��.=f-=;R+=��)=m�(=sg(=��(=)2)=�*=Z�*=�+=m�+=��+=+=U/*=�)=Y(=�'=�m&=|&=9�%=��%=i=&=�w&=��&=$5&=�v%=8:$="�"=�| =�P=�==Zt=	=:!=��='=�h=�P=ʓ=5=�=�C
=O=yj=���<���<�h�<��<[��<���<g��<!�<+��<5B�<t�<W@�<��<���<^��<0>�<S7�<彲<���<u�<e�<�r�<���<ܙ<E�<r��<�<]a�<q�t<�j<0�b<�6]<CY<PoU<�.Q<�:K<��B<8<�*<�I<�7<��;Ă�;��;��;Z%�;�>�;�7�;)�;i˛;V��;�x;B�N;��;���:]Ix:�`|9{uֹ�6��\ƺV����J=�/[^�@H���\��%i��M�̻���j��K��E�?2 ��&��X*�R@.���2���8��A�HK��W��{c��{o�}�y�&ŀ�%'�����g���� ��2?��}���������Y턼���1>��a��/d�����<C��猼P<��񏋼F8���~��z���k���
U��D������R���7���K��w1��-��b��(��������q�������ƛ�W�:�������ݨ�ߔ��v�����P��Ӽ��vX��Q������[����@��I���'
���|��~���	*��a+��.�������n��/W�����̴������O��uǽ�����"eż��ȼ��ʼ�˼z�˼��ʼ�gɼ!-ȼ��Ǽy?ȼ.ʼ��̼��м�tԼ�ؼ-�ڼ�  �  zB=��A=g�A=�>B=R�B=U�B=��B=L4B=ʀA=k�@=��?=�i>=+h==��<=�;=8c;=j;=�:=k�:=��:=4R:=\�9=��8=��7=�[6=��4=f3=k02=PY1=��0=E�0=
H1=D�1=�2=_2=e�1=��0=6�/=u.=��,=X�+=Ե*=[Y*=�e*=��*=�A+=E�+=*,=^ ,=g�+=�+=�Y*=�z)=K�(==�'=�M'=��&=�&=�&=B�&=�&=P�&=�;&=��%=ʚ$=v?#=8�!=��=��=_S=u�=�=��=?=��=I�=�=�H=iK=��
=�P=��=� =b��<��<�^�<b[�<��<���<���<���<f9�<'�<��<}��<J�<�s�<��<��<O�<��<�ի<�ҧ<��<�K�<.|�<7�<k��<���<޾�<��|<d�r<׈j<T�c<�<^<�Y<cS<rL<`�C<�9<d�,<�s<�<�<���;���;�>�;���;[B�;/�;��;��;3o�;:+y;��P;��$;�:���:��9�0���H��W��O��d�9�=�[�,n����z��ȾûD�ܻ^n��4%�99�����In%�v�*�3�0��7��?�ǗI�cMT�rZ_��i���r�*�y��p~��o�� ̀�V����_��vU��M���Q���3킼6����^�����釉�l���1X��氋����Ex��m0��h�� f���@��黍��Џ��W������r���V�� v�������;��RH��N������u㗼��ך��k��"P������J��U����D����&l������1���4़�]��x��r��M���-��H2��<���D`���q���)������|ϳ����뗴�h������H��� ����y$¼�ļ��Ƽ<)ȼ�ȼ�6ȼ�Ǽ`Ǽ��Ƽt�ǼIZɼ`�˼�μ��Ѽ��Լ��ּ�  �  �C=�C=�eC=HKC=�'C=3�B=�vB=j�A=^(A=�Z@=`�?=Q�>=��==iN==��<= <=�;=F$;=��:=�`:=]�9=�u9=f�8=�8=�7=��5=h�4=��3=X-3=W�2=�`2=O2=T2=�L2=�2=�1=I�0=��/=��.=�-=m-=��,=*,=�,=,=D(,=�,,=�,=��+=BX+=��*=�3*=��)=8)=$�(=�(=Y�'=nR'=�'=��&=��&=$:&=��%=R%=9�$="�#=�d"=2!=8�=,=��=4O=&=/�=3`=U�=��=�9=2j=�V=%'=�=�=C��<V�<N>�<���<���<9�<aC�<���<�a�<��<�k�<�=�<X�<���<Կ�<k��<Q��<nİ<��<���<�6�<�Ϟ<�O�<���<�Ȑ<j��<殆<���<�7z<��q<��i<��b<d�[<��T<��L<�C<�D9<+�-<�!<��<�
<�S <t��;�;�;���; �;�h�;��;�;9��;Q�s;�rM;�%;Zt�:'�:0:�b86������� �y\�P;�	_�﹁�ʚ���k���@����һR�������w�����U!��$(��T/�7�l�?���H��RR���[�+�d��hl���r�zw�	.z��2|���}��~�#4��&��G��Ȋ��hۄ�� ��]D���;����C����Z��Պ�O,���m����q�� ���۵��z���"q��W5��J���Tؖ��y��򤗼����?M��P�����Ę��P���A���Y���Q��������������	�����)c��`���O𥼲.��ã���3������A7��O����į��鰼�����岼ܴ��Lv���D��"=��cx�� ��麼���S��qu��8EüȠļ1zż�ż�Ƽ�8Ƽ�Ƽ�Ǽ�ɼq˼4]ͼ3�ϼ��Ѽ�{Ӽ�  �  �XE=��D=(^D=��C=m5C=<�B=��A=�A=�O@=�?=G+?=`�>=�G>=��==n@==�<=��;=�;=tR:=B�9=�9=P�8=1+8=�7=c77=s�6=��5=G5=��4=��3={r3=?3=G�2=OI2=S�1=zg1=
�0=1'0=�|/=��.=�W.=!�-=S�-=4=-=��,=��,=B,=��+=��*=�v*=� *=��)=sY)=�)=X�(=�(=�:(=��'=�"'=t�&=�%=�l%=��$=�|$=��#=�f#=z�"=�!=�� =X=��=�v=\�=X:=�o=�x=!I=~�=|8=Zt=�=u�=E=�� =��<�+�<ݩ�<*"�<���<7��<~(�<��<���<�h�<���<t�<8��<���<�Ȼ<k�<��<���<���<T��<BC�<��<���<��<?݌<֨�<[�<� �<Lw<��n<�"f<
�]<��T<��K<�VB<�28<��-<d#<�</�<�T<p0�;���;˝�;W��;�F�;_`�;F�;���;W�e;}C;�� ;,��:�7�:i�V:�_f9l�عKF��[�⺴��`1D��lj�GM������>��������̻9T߻�4�-�����+����&��//��7��U@�^I���Q��Y���`��\g�x�l�Bdq�tKu� �x�� |��6��/���������������ԗ��G���t��E�_���n�������o���|��[C��ݍ�QY���͎�,R������Eݐ�㑼<���,��#��������]��S떼h����<��<5��Nf��뷛��	���A���P���7������̡�h�������㤼6:��Ś��"�t��8"��� ���̬�����6����߯��N���ֲ��W��4��������"��Ṽ-麼r��$y������r������}"ü�9ļ(,ż�Ƽ��Ƽoȼ�tɼ8�ʼ��̼μ��ϼR�м�  �  �5F=$�E=��D=M�C=��B=��A=�v@=D�?=]�>=ْ>=Cg>=W>=Y?>=a�==c�==D�<=
�;=��:=�x9=`z8=��7=�47=�6=U�6=M�6=�6=�k6="6=zy5=��4=4=�N3=2=�1=�]1=��0=�^0=9�/=�/=�Z/=h/=��.=�a.=��-=�#-=�J,=[+=o*=Ƣ)=)=Z�(=ҝ(=r�(=-�(=��(=V�(=�t(=k�'=��&=��%=L�$=^!$=b�#=M#=��"=ǖ"=N"=��!=G!=� =��= !=�K=xI=l&=Q�=`�=,=ٲ=�7=��=�W=/�=�=�	�<Y��<��<W�<u��<�@�<N4�<ڐ�<�^�<,��<w��<h,�<��<�<2I�<Y��<�z�<�a�<<��<�B�<9��<ᖖ<1�<,�<���<pj�<�ƅ<�Ł<s�z<}q<S�g<�]<,�S<��I<��?<��5<�,<�"<̤<��<vH<)8�;�b�;���;_�;@�;�	�;�o�;�r;�1P;�r1;(�;���:���:��h:ڡ9�
���䊺Ҟ캙�&�8�T�\'~�,`��sx����������-�˻r�ڻ��뻜����j��r�>���&�y^0� 9��iB�ץJ��0R���X��^�=d��/i�h�m���r�*�w���|������]��o[��ӆ�?��������؇������U���~���*��)]��s�������gq��Ώ�\���1�����\ِ�������������Z���C��dj��������;��}W��*Y���H��i$���㛼�������Ų��v���z���Ѡ�����?|���-���uf����������h물���#���a���%���x��fO�����1ɵ��巼����Ժ�f�����W#��=^��[ռ�Ɵ��S����$��»��güżΑƼ�Ǽ�?ɼ�sʼ"�˼,�̼A_ͼ�-μ�ϼ�  �  �F=J�E=�D=!C=��A=;@=�>=��==j7==�==�N==��==!�==d�==s==�<=VR;=��9=�H8=��6=)�5=�a5=�=5=m5=��5=�"6=�O6=C76=��5="#5=�>4=N=3=�;2=U1=�0=v
0=��/=^|/=&o/=lo/=�_/=P$/=��.=n�-=��,=S�+=�#*=n�(=�'=�8'=<	'=B'=g�'=�N(=��(=W�(=�a(=/�'=�a&=��$=R�#=rx"=Ϫ!=�@!=�*!=�H!=�l!=�e!=)!=�= =D�=�S=L=v=�=�=K�=�@=�=��
=m�=�]=�=��=@:�<ŉ�<�m�<n�<?��<"��<lk�<w��<�<�<�6�<sF�<���<�r�<�,�<a�<FU�<1q�<�ۡ<H�<! �<�?�<�:�<YǍ<D��<��<q�<�r�<�J|<�{r<��g<�\<9pQ<��F<ZB<<*�2<[�)<S!<�4<c<	D	<�� <���;���;���;�0�;��;$�z;&|T;f4;U';��;B��:��:'�f:l
�9����L���v �t7��k���������񭻇���Ļ'2ϻ:"ۻ�b�LG�����{�Z����'�$�2��<��wE�OIM�;�S���Y��p^���b��g�C�l�~r���x�I���b���y���戼q�����;����������KӇ�^����K��'Ή�d��C���E�����Q��{����K��l^��M<��oB����� Ր�K����ђ��{��kT��Y ������O��؛��h��\���z����Ĝ�N���Ý��������^r��7V��WL��/����	��
N�������`��l����������B������d� ʴ��ⷼ�ĺ�}���|��h��s�va�������N���h������o��J=���Zü��ż8�Ǽ	lɼ��ʼ��˼?�̼1ͼQbͼK�ͼ#Zμ�  �  YqF=kE=s�C=�,B=Q:@=�_>=��<=��;=I_;=�;=<=��<=a^==x�==�.==7<=4�:=x�8=�6=.F5=�4=rn3=�c3=�3=܅4=�D5=��5=C�5=��5=�5=�4=��2=��1=ė0=�/=�%/=��.=��.=/=|8/=XL/=�/=4�.=K�-=�,=�m*=��(=�'=��%=�I%=�B%=��%=��&=�'=�>(=�v(=�(=� '=2�%=��#=�*"=b� =��=!J=�X=��=!? =�� =X� =� =8�=v,=G=_�=��=�5=ܧ=�B=�=�
=c===�=^�=��<�l�<I��<�t�<)m�<��<�f�<'��<��<�8�<�4�<��<�	�<B��<��<�"�<Cϭ<�.�<�<�<a�<%��<��<1�<��<��<���<�H�<.|<r<��f<��Z<ӓN<�C<�n8<q�.<fd&<a�<�<n�<�<l��;��;�|�;9��;[�;QA�;�\;Y5;V�;�� ;�I�:Q|�:}�:�W:�9�ٹ.4����k�J��Ł��0����I任"0ƻ�
λyջD�޻���V��������_���)�3n5��?�7�H��dP�aV��"[�6/_�^+c���g��(m���s���{�����G�����������H����������H���� ��k���.7��tڈ�c���k��*���F���w���.)��@���Qޗ��_���������چ���#��.����󒼅ߔ� ���Y��>G�����&����일�ʝ��h��"��D'��᝼�o���ࡼ����Ũ��r��J����:��������ܟ���;���~��̮��L�����o���H���ὼа��a¼��¼W\¼V'������c������DT��`����o����ü�~Ƽ��ȼ�˼��̼2�ͼdμ�μt�ͼ{�ͼ	nμ�  �  �#F=��D=�BC=�*A=T�>=��<=�%;=�:=J�9=+:=B�:=��;=3�<=�'==_�<=��;=�:=�7=��5=��3=Eg2=��1=ҷ1=Q2=-H3=�T4=�+5=֔5=�w5=!�4=��3='~2=� 1=��/=]�.=�W.=.= 9.=��.=��.=/=�.=8..=�,=�O+=�Q)=�G'=�}%=�3$=��#=y�#=Fr$=�%=�&=�'=�(=ϻ'=�&=��$=��"=�� =�&=�=��=8�=J=�=Ĺ=��=V�=B�=�=~�=��=m,=kd=u�=a=�?=�U	=f�=˯=֟=�4=��<��<���<���<]�<!��<C��<j��<��<��<�N�<l��<+�<�N�<V�<��<4J�<C�<�:�<�h�<��<�F�<j�<z��<���<?{�<��<���<B1{<	�p<>#e<~X<<�K<��?<�5<��+<lx#<p<5�<�.<�<���;L��;�t�;�U�;bW�;Q]q;�@;	{;�$�:�2�:�̽:��:"!�:ӚA:�W`9_��zh��f��7K\�i���߭��������Ȼ �ѻ�n׻v�ܻuB�ǐ�OD��������w[�A,��8�,�B��L��HS���X��\��`��$d���h�dqn�>�u��~�&B���	���(���$������̥���E�����򛋼����񈼩���X����׎�/�������������� �����`7��#Ȗ��g�������ۑ��)���y�����������������R��l/���X��p���jI��Ÿ��2���zm��n:�����V榼�0���e�����b�� o���������s��I���Xb��~�����C�����I}������]�ü��ż�IƼ{ż�ü����z�������������%�����ļڇǼzNʼ>�̼�Eμ"/ϼ~jϼ4(ϼW�μ�μ�μ�  �  ��E=��D=��B=dg@=��==ƻ;='�9=M�8=w�8=o 9=`#:=�W;=4[<=��<=ˎ<=Us;=��9=bS7=D�4=�2=�F1=]�0=(�0=v@1=�_2=��3=+�4=y45=D.5= �4= �3=�$2=��0=	e/=d.=*�-=��-=-�-=�%.=ۍ.=*�.=v�.=-�-=��,=&�*=1~(=mG&=�\$=�#=xl"=��"=��#=��$=�C&=�X'=��'=]q'=�B&=�i$=u0"=@�=�=^�=Y=͊=~@=�2=�=�v=\9=�<=߈=_>=��=�=}�=�(=K�=+�
=��=\=zW=PP=y� =m��<G��<�1�<�<Y3�<�+�<Oo�<[;�<ׇ�<$��<m��<w��<�{�<Tſ<�W�<�R�<o,�<r��<8d�<tI�<�Í<��<�<���<��<�S�<gɃ<�<�!z<�o<��c<�V<(�I<x�=<�2<hG)<�d!<��<n<��<{V<��;�l�;���;P�;á�;��_;"�-;ܢ;{��:��:��:ER�:E0�:�/:;�$9d+�����o�#�u�h��N��wB���û��ѻ��ٻ0g޻8��jD�Ma��b��������� �Ŭ-��:��E��4N��TU���Z�6x^��a��(e�k�i���o���w�/����ㅼ����f����������ē�����{��������������#���]��X叼"���T�������ٝ��_��%e��z@���y��5�������*���˴������*��kΘ��z��_ɝ�do���I��\��ӟ�� ���O���/�� ���W���� ��;K��h���T��[B������-�������G��lճ�8�����������ⴼ�8�����¼�Ƽ�(ȼu�ȼ��Ǽ��ż�]ü�0���п�+���ϊ��>�¼�Gż�TȼYB˼Z�ͼ�cϼ�CмZbм��ϼeeϼ<ϼPtϼ�  �  V�E=�dD=�xB=�@=�==�V;=��9=D~8=TA8=��8=��9=a;=�1<=[�<=�s<=cR;=r9=q7==�4=s2=��0=�0=�#0=��0=.
2=�W3=�o4=�5=(5=0x4=d3=�2=ߊ0=�6/=2.=j�-=Uh-=�-=O .=�m.=ݦ.=�v.=,�-=�Z,=�p*=�/(=�%=�#=o�"="=$A"=�5#=��$=�&=O3'=ɯ'=�T'=x&=�7$=��!=g�=��=�o=��=� =�=��=��=�D=2=(=�h=#=�c=�}=��=)�=�=�}
=«=��=6=�1=�� =-��<9��<��<�h�<�n�<qV�<t��<�l�<���<�_�<�z�<FX�<v9�<���<��<��<�ª<0�<���<܅�<W��<�"�<i�<��<�{�<�ބ<�q�<�̀<9�y<�Wo<~=c<�1V<�I<T�<<��1<{w(<~� <<R�<�o<��<��;��;y��;6˨;���;�sY;!)';N ;���:3��:([�:Ь�:��x:"):}p9�X���ƺ�{'�3m�	���Z���ƻ,�Ի��ܻ�ở他������S��&	����;!�O.���:���E���N�!V�B[�X
_��/b���e�j��5p��Ux�����~�����5��(W���͔����ܻ�����p���ʊ�����[�����%H������
���A��0����7��n6������(���4������/ϒ��:���i�����Л�)���ԟ���������%��G��]����g��X8���>������>Ѩ�˞��=B��|������c���LԸ�T㶼�P���ⱼ Y��E���챼3�����𕾼�9ü��Ƽ��ȼ}ɼ��ȼFvƼ��ü�����%��tԿ�<�����¼�ż�ȼO�˼�μ}�ϼ��м~�мHм��ϼ�Oϼd�ϼ�  �  ��E=��D=��B=dg@=��==ƻ;='�9=M�8=w�8=o 9=`#:=�W;=4[<=��<=ˎ<=Us;=��9=bS7=D�4=�2=�F1=]�0=(�0=v@1=�_2=��3=+�4=y45=D.5= �4= �3=�$2=��0=	e/=d.=*�-=��-=-�-=�%.=ۍ.=*�.=v�.=-�-=��,=&�*=1~(=lG&=�\$=�#=wl"=��"=��#=��$=�C&=�X'=��'=Yq'=�B&=�i$=m0"=6�=�=Q�=�X=��=o@=�2=�=�v=f9=�<=�=�>=6�=�=��=�*=��=��
=��=3#=�[=U=�� =7��<{��<"=�<�<�>�<�6�<oy�<�D�< ��<�<���<W��<�}�<�ſ<bV�<�O�<�'�<G��<�\�<�@�<���<��<겇<N��<`�<kH�<Ⱦ�<�<�z<��o<s�c<��V<�I<��=<Ū2<�J)<ak!<��<�z<E�<th<�C�;u��;���;|>�;Ќ;�`;".;��;���:�$�:fz�:Y��:�f�:�0:��$9�i�x����*$��h��o���h��?�û%�ѻx�ٻ�޻P/��t�2�𻓏��ݳ����� ���-��:��E��=N�`\U���Z��|^�n�a�t+e�S�i��o���w�����4䅼-���f��1��������ē����	|������%��������#���]��Z叼"���T�������ٝ��_��%e��{@���y��5�������*���̴������*��kΘ��z��_ɝ�do���I��\��ӟ�� ���O���/�� ���W���� ��;K��h���T��[B������-�������G��lճ�8�����������ⴼ�8�����¼�Ƽ�(ȼu�ȼ��Ǽ��ż�]ü�0���п�+���ϊ��>�¼�Gż�TȼYB˼Z�ͼ�cϼ�CмZbм��ϼeeϼ<ϼPtϼ�  �  �#F=��D=�BC=�*A=T�>=��<=�%;=�:=J�9=+:=B�:=��;=3�<=�'==_�<=��;=�:=�7=��5=��3=Eg2=��1=ҷ1=Q2=-H3=�T4=�+5=֔5=�w5=!�4=��3='~2=� 1=��/=]�.=�W.=.=�8.=��.=��.= /=�.=7..=�,=�O+=�Q)=�G'=�}%=�3$=��#=w�#=Cr$=�%=�&=�'=�(=ƻ'=ݣ&=��$=q�"=p� =�&=�=�=�=�I=l=��=��=j�=�=��=S�=��=Y.=g=��=�e=�D=\	=Ώ= �=��=�>=���<N#�<���<� �<�r�<���<���<B��<ש�</��<Y�<��<A/�<�O�<��<��<AA�<_�<�+�<#X�<���<2�<#҉<�r�<���<�e�<���<���<\{<p�p<�	e<�jX<u�K<v�?< 5<��+<:�#<�<'<(M<Ĩ<��;D9�;���;뮱;䰔;�r;�TA;p;h?�:�(�:E��:�|�:���:c B:$2`9 `�۴����w�\���������n���i�Ȼ3�ѻf�׻f�ܻ��z�����������|��%,�78��C��L�CWS� �X�-]���`��)d�F�h�0tn�Y�u���~��B��e
��?)��%��򫑼󥑼�E������������"񈼰���^����׎�2�������������� �����a7��#Ȗ��g�������ۑ��)���y�����������������R��l/���X��p���jI��Ÿ��2���zm��n:�����V榼�0���e�����b�� o���������s��I���Xb��~�����C�����I}������]�ü��ż�IƼ{ż�ü����z�������������%�����ļڇǼzNʼ>�̼�Eμ"/ϼ~jϼ4(ϼW�μ�μ�μ�  �  YqF=kE=s�C=�,B=Q:@=�_>=��<=��;=I_;=�;=<=��<=a^==x�==�.==7<=4�:=x�8=�6=.F5=�4=rn3=�c3=�3=܅4=�D5=��5=C�5=��5=�5=�4=��2=��1=ė0=�/=�%/=��.=��.=/=|8/=XL/=�/=4�.=K�-=�,=�m*=��(=�'=��%=�I%=�B%=��%=��&=��'=�>(=�v(={(=� '=�%=p�#=�*"=C� =ٸ=�I=�X=z�=�> =�� =S� =� =��=+-=|=A�=~�=�9=Ԭ=I=S=�

=�=#==W�=���<Y��<���<��<܋�<��<B��<[�<A��<KK�<RC�<�	�<��<���<���<��<�­<��<�Ϟ<�i�<�F�<�x�<�Ԍ<L �<�<�ȇ<wl�<�-�<��{<��q<ؐf<��Z<]�N<eC<'n8<3�.<}v&<^�<��<�<J�<�
 <�t�;��;�6�;��;m��;Q�\;X�5;�;7�;�h�:[X�:3}�:ڪW:y�9�۹�գ�^��4K�� ��?���@���~`��o�ƻ<�λ��ջ�
߻��������v���*��5�m�?�KI�yP�qV�/[��8_��2c���g��,m���s�ӣ{����TH��'���
���8I��׉��ޡ��h���	!��}���;7��~ڈ�k���k��/���I���z���0)��B���Rޗ��_���������ۆ���#��.����󒼅ߔ� ���Y��>G�����&����일�ʝ��h��"��D'��᝼�o���ࡼ����Ũ��r��J����:��������ܟ���;���~��̮��L�����o���H���ὼа��a¼��¼W\¼V'������c������DT��`����o����ü�~Ƽ��ȼ�˼��̼2�ͼdμ�μt�ͼ{�ͼ	nμ�  �  �F=J�E=�D=!C=��A=;@=�>=��==j7==�==�N==��==!�==d�==s==�<=VR;=��9=�H8=��6=)�5=�a5=�=5=m5=��5=�"6=�O6=C76=��5="#5=�>4=N=3=�;2=U1=�0=u
0=��/=^|/=&o/=lo/=�_/=O$/=��.=m�-=��,=R�+=�#*=m�(=�'=�8'=9	'=�A'=a�'=�N(=��(=K�(=�a(=�'=�a&=��$=2�#=Mx"=��!=Y@!=Z*!=NH!=�l!=ie!=$!=�= =��=�T=�M=�=k�=5!=c�=�H=s�=ӻ
=;�=l=�/=��=�^�<j��<��<�5�<���<;��<=��<F��<'8�<��<�H�<ES�<���<Ft�<�(�<p�<�E�<�\�<�¡<7�<���<��<��<{��<E^�<[�<��</Q�<|<�Fr<��g<�z\<kXQ<�F<hA<<ߔ2<z�)<V@!<�_<h�<N�	<r� <�Q�;�2�;�n�;H̪;Չ�;��{;y�U;�Y5;C�;�;���:Ǯ:ͨg:��9����_q����,8� �k�l���n�����2���mRŻ�ϻ��ۻB �%���t�-������(��2�5�<���E�4bM��T�Y�Y��|^��c�̨g�F�l�݁r���x�i��Sc���z��B爼`q�����n���<���å��aӇ�o����K��0Ή�k��I���I����� Q��}����K��m^��N<��oB�����!Ր�K����ђ��{��lT��Z ������O��؛��h��\���z����Ĝ�N���Ý��������^r��7V��WL��/����	��
N�������`��l����������B������d� ʴ��ⷼ�ĺ�}���|��h��s�va�������N���h������o��J=���Zü��ż8�Ǽ	lɼ��ʼ��˼?�̼1ͼQbͼK�ͼ#Zμ�  �  �5F=$�E=��D=M�C=��B=��A=�v@=D�?=]�>=ْ>=Cg>=W>=Y?>=a�==c�==D�<=
�;=��:=�x9=`z8=��7=�47=�6=U�6=M�6=�6=�k6="6=zy5=��4=4=�N3=2=�1=�]1=��0=�^0=9�/=�/=�Z/=h/=��.=�a.=��-=�#-=�J,=[+=o*=â)=)=U�(=̝(=k�(=$�(=}�(=I�(=�t(=W�'=��&=��%=(�$=5!$=3�#=#=��"=��"=�M"=��!=E!=� =3�="=�M="L==*=��=.�=�4=N�=�C=��=h=� =2�=2�<e�<���<)G�<k��<�h�<�Y�<&��<�|�<���<���<�:�<�"�<3��<wD�<L��<�i�<�J�<bs�<�"�<x�<�o�<�<붏<���<�@�<��<���<׍z<�Aq<��g<��]<��S<��I<��?<��5<T3,<��"<��< <��<���;��;�w�;*�;h�;R��;��;3s;BAQ;�^2;�;	�:�h�:�^i:���9�׶� ��� ��ޢ'�i�U�]C������!��訰��u��K�̻)�ۻ�<��:��Ÿ�]�������&�o�0�2�9�H�B���J��FR��X�d�^�)Gd�^7i��m��r�^�w� �|������^���[���ӆ���������؇�����U���~���*��4]��{�������lq��
Ώ�^���3�����^ِ�������������Z���C��dj��������;��}W��*Y���H��i$���㛼�������Ų��v���z���Ѡ�����?|���-���uf����������h물���#���a���%���x��fO�����1ɵ��巼����Ժ�f�����W#��=^��[ռ�Ɵ��S����$��»��güżΑƼ�Ǽ�?ɼ�sʼ"�˼,�̼A_ͼ�-μ�ϼ�  �  �XE=��D=(^D=��C=m5C=<�B=��A=�A=�O@=�?=G+?=`�>=�G>=��==n@==�<=��;=�;=tR:=B�9=�9=P�8=1+8=�7=c77=s�6=��5=G5=��4=��3={r3=?3=G�2=OI2=S�1=zg1=
�0=1'0=�|/=��.=�W.=!�-=S�-=3=-=��,=��,=@,=�+=��*=�v*=� *=��)=lY)=�)=M�(= �(=�:(=��'=�"'=U�&=��%=jl%=��$=�|$=��#=�f#=I�"=Ź!=�� =>X=T�=�w=4�="==�s=c~=/P=`�=OC=-�=��=�=xW=�� =���<�W�<=��<N�<a��<��<qO�<k��<	�<Ԃ�<��<Ղ�<���<O��<Ļ<�_�<l�<��<�n�<㝡<��<\��<d͔<1ǐ<N��<�}�<�1�<K�<kw<pnn<��e<@u]<)�T<�K<�UB<�>8<?�-<�(#<��<��<P�<\��;�J�;�L�;�V�;��;��;���;>!�;�	g;D;�a!;�*�:��:�OW:@f9��ڹ�(���Ԏ��0E���k����\���y��Ļ�I�ͻ�������oP�0u��O���&�b/���7��y@�H%I���Q��Y��a��gg���l�Ijq��Ou���x�Z|��8��0��2�����S��6������i���t��Y�n���y�������v������_C��ݍ�SY���͎�-R������Eݐ�㑼<���,��#��������]��S떼h����<��<5��Nf��뷛��	���A���P���7������̡�h�������㤼6:��Ś��"�t��8"��� ���̬�����6����߯��N���ֲ��W��4��������"��Ṽ-麼r��$y������r������}"ü�9ļ(,ż�Ƽ��Ƽoȼ�tɼ8�ʼ��̼μ��ϼR�м�  �  �C=�C=�eC=HKC=�'C=3�B=�vB=j�A=^(A=�Z@=`�?=Q�>=��==iN==��<= <=�;=F$;=��:=�`:=]�9=�u9=f�8=�8=�7=��5=h�4=��3=X-3=W�2=�`2=O2=T2=�L2=�2=�1=I�0=��/=��.=�-=l-=��,= *,=�,=,=C(,=�,,=�,=��+=?X+=��*=�3*=��)=/)=�(=~(=H�'=ZR'=�'=h�&=��&=�9&=d�%=�Q%=�$=�#=Yd"=!==�=j=D�=OP=�=��=d=��=ɱ=~B=�t=(c=t5=�=f-=��<�~�<jh�<y��<X�<�b�<�k�<�!�<���<���<?��<�Q�<��<���<���<���<N��<b��<�<؁�<��<x��<�(�<�|�<���<���<5��<���<3�y<�lq<F�i<?�b<��[<9�T<ҼL<��C<�P9<��-<�"<�<��
<l� <IR�;7��;�D�;0��;!�;��;���;^6�;�t;�]N;�&;���:��:��0:��`8��2_���=�5)��F<�Q-`�W��D��~�������ӻR:�{3��������@���W!��](�݅/��67�ӧ?���H��hR� �[���d�-sl���r�fw�x2z�36|��}���~��4���&��G������ۄ�� ��~D���;��(��Q����Z��Պ�U,��n��񳋼t��"���ݵ��{��𣐼#q��X5��K���Tؖ��y��򤗼����?M��P�����Ę��P���A���Y���Q��������������	�����)c��`���O𥼲.��ã���3������A7��O����į��鰼�����岼ܴ��Lv���D��"=��cx�� ��麼���S��qu��8EüȠļ1zż�ż�Ƽ�8Ƽ�Ƽ�Ǽ�ɼq˼4]ͼ3�ϼ��Ѽ�{Ӽ�  �  zB=��A=g�A=�>B=R�B=U�B=��B=L4B=ʀA=k�@=��?=�i>=+h==��<=�;=8c;=j;=�:=k�:=��:=4R:=\�9=��8=��7=�[6=��4=f3=k02=PY1=��0=E�0=
H1=D�1=�2=_2=e�1=��0=6�/=u.=��,=X�+=Ե*=[Y*=�e*=��*=�A+=C�+=(,=\ ,=d�+=|+=�Y*=�z)=C�(=3�'=�M'=��&=�&=��&=(�&=ͣ&=+�&=�;&=��%=��$=G?#=�!=��=��=�S=�=�=J�=�='=��=4�=ZP=�T=�
=�]=U�=� =ѷ�<,�<���<΁�<A��<>��<}��<@��<X�<B�<���<o��<
!�<�z�<j�<a�<#E�<��<���<Ĺ�<���<�+�<FY�<M�<�b�<�u�<}��<�9|<J�r<�Kj<�c<Y^<��X<KS<heL<l�C<�&9<��,<�<e<B<��;
y�;���;[Z�;�ݽ;-ʴ;���;��;���;�z;D�Q;��%;�:�_�::�9��0���I�����k�E��Wr:���\��������6���bĻiyݻ���Ut����c��O��)�%�q+�6�0�=�7��@��I�zaT�Ej_�P�i��r�Q�y��u~��q���̀�y����`��V��ʸ������y킼k����^����� ���~���>X��𰋼���Jx��q0��k��#f���@��껍��Џ��W������r���V�� v�������;��RH��N������u㗼��ך��k��"P������J��U����D����&l������1���4़�]��x��r��M���-��H2��<���D`���q���)������|ϳ����뗴�h������H��� ����y$¼�ļ��Ƽ<)ȼ�ȼ�6ȼ�Ǽ`Ǽ��Ƽt�ǼIZɼ`�˼�μ��Ѽ��Լ��ּ�  �  )&@=��?=�J@=��@=��A=�*B=�[B==B=�vA=t@=7?=��=={�<=z�;=��:=�:=wg:=�q:=��:=��:=rH:=B�9=��8=�7=*V5=�p3=�1=�G0=�g/=3"/=_l/=�0=��0=C�1=߲1=�Q1=�Y0=��.=f-=;R+=��)=l�(=rg(=��(=(2)=�*=Y�*=�+=k�+=�+=+=Q/*=�)=S(=�'=�m&=p&=*�%=��%=T=&=�w&=�&=5&=�v%=:$=��"=z| =�P=>=�t=}="=6�=(=�k=�T=ɘ=�"=��=�L
=�Y=Uv=��<��<���<�4�<���<���<���<m!�<���<1[�<w+�<�R�<l�<��<H��<o?�<�3�<ѵ�<[��<���<�P�<O[�<j�<���<K�<�}�<ˆ<�B�<פt<>�j<[�b<R]<��X<�RU<�Q<30K<��B<�8<U+<�d<l[<�\�;���;���;Rb�;-��;d��;W��;�l�;JA�;�b�;�ny;FeO;�~ ;���:\ny:F�~9֏ֹ���M�ƺ�V�ޣ���=�.*_�ﺂ�wؘ�뱻�>ͻ�W�	0��V�J���k ��6&�Q�*�j.���2�99��7A��\K��W���c��o�<�y�Ȁ�])��x �����������?��������4���턼��J>��t��=d�����EC��%猼U<������I8���~��{���l���U��E������S���7���K��w1��-��b��(��������q�������ƛ�W�:�������ݨ�ߔ��v�����P��Ӽ��vX��Q������[����@��I���'
���|��~���	*��a+��.�������n��/W�����̴������O��uǽ�����"eż��ȼ��ʼ�˼z�˼��ʼ�gɼ!-ȼ��Ǽy?ȼ.ʼ��̼��м�tԼ�ؼ-�ڼ�  �  m>=/I>=��>=��?=�@=�yA=5�A=�A=�6A=)@=J�>=^==�<=��:=�,:=j�9=��9=4�9=,:=,D:=�:=�T9=8=Y^6="G4=�2=�0=y�.=I�-=k�-=�.=�/=0=��0=�Q1=k�0=�/=y6.=d(,=�*=�N(=�!'=��&=P�&=�'=z�(=k
*=L�*=�n+=�_+=��*=��)=խ(=�v'=�g&=��%=�8%=�)%=de%=C�%=�$&=�B&=��%=f%=ӭ#=�!=�\=��=��=��=�r=ڪ=�Q=%=*�=��=�S=:�=�=��	=�b=5=���<��<�=�<;$�<�%�</��<�D�<�-�<��<���<���</��<"�<7��<�M�<l��<K��<@�<��<��<���<)��<5�<X̘<��<'�<�4�<
[z<��m<Ĥc<)&\<�<W<&5T<��Q<O�N<{�I<��A<M�6<��(<3=<�	<|�;#a�;�<�;�Q�;Z��;é;K�;��;�ʘ;�
�;�Wu;�uJ;��;��:Z�J:#8N#�,O��#q޺��_'�b�C�A�d���b��~���3ֻ������ X����H�&���+���.���1��85�ѱ:�d�B�I=M�~�Y�hg���t����(�������t��膼�|���΃�6x���恼-H��
������������m��f������������������[)���;��K�����"Q��{����	�������뚼P��P���Ϊ���?��\���[�����R���'��C��Μ� x��Y���B¨����'���<���Pȭ�����멼]맼%���*J������ʨ��<������°�����ƴ� ����������	D����e.���G��1m��ǡ������,&ļ3kȼX�˼DGμ�2ϼӹμ�0ͼ.˼�gɼR�ȼ�ȼz�ʼ�μ�CҼ��ּ<�ڼ��ݼ�  �  �>==$==��==��>=��?=��@=E�A=�A=��@=��?=�y>=@�<=;=�a:=�9= D9=�G9=׉9=R�9=�9=D�9=�9=�7=��5=�{3=C1=!�.=4d-=��,=t,=�-=�A.=��/=ݏ0=�1=)�0=�/=��-=�z+=�5)=�G'=��%=~%=��%=N�&=��'=�Z)=Pv*=z+=�+=��*=�)=mQ(=�'=��%=�%=V�$=��$=��$=�k%=�%=@&=L�%=b�$=t6#=�!=̆=��=m�=F�=CU=��=�z=�}=�S=۞=�=��=M7=!	=��=/V =g��<0��<V��<O��<�:�<�(�<��<�T�<�}�<�g�<�(�<��<]�<j��<�;�<Vt�<�r�<7�<䚬<oR�<D��<�+�<���<���<�_�<v��<sU�<kv<�#i<��^<��W<�GS<a�P<�^O<��L<0rH<w�@<��5<kI'<.�<��<H��;���;1�;
0�;�B�;�m�;,�;���;^��;u��;Xq;�E;c�;3��:��):R׸,�I�ۯ�'�(	��-�	�H�F�i��̈�)&��������ܻ1���F?�`(�xI$��Y+�q�/��2��
4��6���;���C�^�N���[��&j��x�����u��{���Ɖ����BB��]1��k{��I����؂����c/��b����O��"�����D֏�)�G��N獼K׌�%E�� ������ ���^����������$����	�������U��Hh���������>��]����ښ�\���񔡼�+������'���R��7谼����������)���~���寮M���^U���ޫ�Qͮ�I���$��u䵼�Զ�b�����������~���N���6ܶ��1��۵��i&��k�ż4�ʼ^Eμ��м2qѼ��м�μ't̼�Tʼ/-ɼ�~ɼ�y˼��μ
Ӽ�]ؼC�ܼL+��  �  `~F=�+F=�BF=ƛF= G=W5G=G=H{F=JxE=nD=�B=0�@=Δ?=Bt>=�==�R==O==ǎ==��==�;>=P>=b>=�L==i'<=�:=29=Õ7=1c6=��5=SZ5=W�5=�6=P�6=�7=�47=2�6=��5=�w4=s�2=�91=g�/=��.=�^.=)X.=�.=�>/=J�/=b	0=��/=5_/=pi.=r'-=V�+=�f*=�>)=g(=��'=��'=1(=Dv(=��(=5)=�.)=x�(=�'=�J&=��$=ߎ"=@� =�=U�=W�=E�=8[=3�=�|=d�=�w=x=�=bl=�=ڏ=��=���<[<�<�X�<���<6�<���<��<v��<��<�7�<,��<���<��<O�<>�<�"�<驴<�<���<sp�<p��<~G�<��<vH�<g%�<�<Ɗ�<>ā<��{<۸u<d�p<��l<��g<|�a<��Y<�SO<��B<S�4<��&<*�<?�<�<��;���;�;[��;V��;:U�;eu�;6Н;��;�cX;Jx#;�3�:�#�:a�9�U_�g2�1���+5���k�ټ�o�1��>X�;c������ƍ���Mͻѱ�3�������������H��-���P$��-�9���D���O��mY�K�`��f���h��i�1[i���h�`�h��4j��m�coq���v�l�|�#��A[��d���\ׅ��酼P��E��$���0���ׁ� O��E����م������r��v���Z؏�ː��̐�B������4d��ʁ��G��9����ď��������Q.������Fy���>���#��{h���r��߸����P]��� ���i��vT���j��"Q��к��At���j������1G��|���0䬼P����䬼����(��Q����4���h��Z$��F����$"���w���o��Ⴜ�},��Vͼ�����PH��b�ļV1ȼrh˼�ͼ�  �  9�F=
kF=�~F=]�F=P-G=�YG=O-G=�F=z�E=9D=��B=%A=ӿ?=+�>=��==a�==2y==�==Z>=OV>=h>=�>=�k==�M<=�:=UM9=��7=��6=��5=ғ5=?�5=D)6=F�6=�$7=�97=g�6=�5=7�4=��2=�e1=�0=�/=�.=��.='�.=xq/={�/=:+0=�0=Mw/=L�.=�D-=��+=��*=�j)=J�(=�(=Y(=d4(=+�(=M)=�M)=F)=z�(=�'=�r&=��$=z�"=n� =�D=��=��=�'=Ty=a�=T�=e�=Hw=��=�"=�==��=��=�P�</��<ƽ�<{�<BT�<���<���<y��<���<`q�<%��<:3�<L�<�u�<`��<Z~�<���<��<�<���<`�<ω�<�g�<���<8��<���<��<9H�<,�|<`�v<�q<"m<�>h<yb<?�Y<�`O<��B<i[5<Lx'<�M<U�<o�<ބ�;
��;�'�;��;���;i&�;�'�;;�׆;okZ;��%;��:�%�:̵�9g.���&��O�������e�l���/���U�����Y��Z����=˻���\������!�c�Wu�!S��j��<$�=�-��8��%D�O���X�D`�e���g���h� �h��h�Oh�{�i�ͷl��
q�wVv�	|�廀�}������Rz��j�������q���6������ާ��Q��+j��R����0�� �����iY���P���^�������u��w:���n��hx��Ə��`���b���;����Θ�}O��i��������������a��Cj���_��i)���Н�R5��_���!������Y`��"������M��t����Q�������^��ճ���ܭ��᯼꠲�q˵��<���&���񚾼˹��|$��X5��Ga�����dǼ�����)���pļ��Ǽ-˼:wͼ�  �  �nG=�G=�&G=fG=ĨG=]�G=�yG=`�F=!�E=8�D=�
C= �A=C9@=^%?=�f>=>=��==�>=�a>=��>=̦>=�a>=+�==Ҵ<=K`;=��9=.~8=�U7=��6=�46=p>6="�6=-�6=�C7=�B7=��6=��5=b�4=-M3=
�1=7�0=�/=#Q/=�F/=��/=�/=�_0=؄0=O0=ص/=��.=��-=�C,=d�*=��)=�)=��(=>(=#�(=!�(=�T)=��)=Q�)=�)=00(=��&=X6%=�a#=��!=~�=��=�}=��=��=\�=ߍ=�=�r=P�=�R=��=�x=7T=��=vO =9��<X��<��<��<���<�@�<^(�<�[�<@�<+��<;�<4	�<c��<3��<�< �<ȩ�<p��<'<�<���<o1�<�7�<���<�ʓ<�<�<ϵ�<�g<.�x<bs<iRn</�h<�0b<�Y<0uO<�pC<�X6<�)<�Y<<x�<F��;x��;U��;Y��;dc�;Db�;��;2q�;�;�`;��,;��:|j�:	:�G	�"O���s��O���޺��q�*�4#P���z�T���X����Żt�ۻ���c���h���U�|\�<���6�M$��z-�7�7�-�B��!M�\.V��S]�QIb��e��;f�Tf��Hf��f��h�R�k� p��u�!�z�
�����	���5o������5���;���@��gx���*����������(�����X����#���򍼹����+������C��Ќ�SB��$n��ဍ�u���������@Ǘ�q��!����X���O������%
����������(����S��M����o���W��$���^��������X��� ��6���?��ޫ��4��LG��$�����J���S����B���1���L�����)A���������.��ο��f��L�����üǼ��ɼ�,̼�  �  }qH=8!H=�H=�7H=QH=>:H=��G=P!G=F=��D=C�C=�'B=�@=��?=K/?=��>=��>=�>=m�>==�>=��>=�>=� >=y<==)<=��:=�u9=-[8=��7=�7=:�6=�7=&H7=�b7=�A7=��6=�6=��4=A�3=�2=�{1=$�0=QV0={F0=w0=8�0=��0=V�0=e�0=0=�/=��-=��,=S�+=\�*=��)=0h)=]9)= H)=8~)=Ȼ)=��)=%�)=�b)=��(=�m'=��%=i>$= �"=r� =i�=?L=�:=v0=�=�=/�=�\='�=��=�M=	=*$=ف=C=߿�<�z�<�`�<E�<�A�<���<��<��<���<*��<�m�<?��<+�<^C�<8��<�.�<M��<yd�<t��<�5�<}�<!F�<3
�<�z�<��<���<Ʌ<\��<�|<,�u<��o<!}i<`0b<��Y<2WO<��C<�7<!+<t;<J�<�W<Z�<���;9��; ��;��;y �;IT�;�Ң;��;c�g;ݡ6;bw;�G�:�?:L.9pA��t�J�|~���?Ѻ����$���H��>q��Ꮋ�>��i��) ӻy�滝M��F��7	����j-�3#�_&$��1-���6��@��xJ���R�1jY�_'^�ca���b�)8c�g�c�>e�Cg���j��n�\}s�sxx�v-}�$�����a߂�}���т��-��Nm���Ѐ����值�݁��}������B����'���狼����u��9S��z׌�T��{��5z������o@���~��l����V���K��/����M���[��b��7���^~��-뙼���W���U���_���<�������਼�z��"}���o꫼ҡ��HT���?��E��������.��i�����'ǵ�_=��$*���i������/���ջ�C�����#м��]�������%üN�ż5VȼSPʼ�  �  T�I=iBI=�!I=nI=��H=ȪH=_ H=,WG=pXF=�3E=��C=R�B= �A=2�@=@=��?=�_?=�F?=�D?=�B?=~*?=,�>=Ap>= �==��<=�;=�:=�~9=��8=�8=��7=g�7=m�7=�h7=i#7=w�6=Z�5=Z5=""4=�03=?c2=�1='z1=b1=�r1=��1=�1=oX1=��0=�50=V/=IW.=N-=�P,=�t+=��*=Q*=�*=��)=A*=�*=$*=��)=��)=��(=X�'=~�&=�*%=��#=�"=^� =�(=2�=ފ={=3p='u=$=�=c�=d�=��	=�=K�=�P=N^ =-�<��<��<���</$�<K�<#|�<���<���<���<oI�<U �<e�<ꪼ<>��<SӴ<�1�<���<(��<��<Z;�<�e�<
B�<��<m�<i�<L��< �<�6x<�q<пi<ϳa<��X<�N<��C<��8<�-<�@"<�R<�<��<{K<S)�;Yk�;pK�;c)�;�߸;��;���;��o;ynA;��;��:[�~:d�9A� ����S����ĺ� ����]CB�k&h������j���`���ɻ�3ݻ2ﻉ��k�����O������$��Q-��X6�<R?�O�G�qO�U���Y�D�\��^���_��}a�I�c��:f�F�i�n�m�7�q�JUv��`z�H�}�A4��8
���j��d��>��Ԧ���I���)��(j���$��c������l������ ۊ�e����?��������0��g�'ȍ�?�����$���ZՔ��[��n��q���4���*���+���{���C��Ɏ��tO��$j����������A���%���������*R��C���¥��h���[Ǫ��1��1��=X���)��/_�����*����巼�T���F��XӺ�c(�����m�����4����h����¼��ļ?�Ƽ�Cȼ�  �  ��J=�EJ=�J=��I=�gI=%�H=�+H=�QG=]F=RZE=�UD=k[C=�uB=5�A=~A=�|@=s@=��?=Ӑ?=�_?=�*?=��>=��>=��==�C==�f<=�s;=�:=>�9=��8=�i8=��7=M�7=u@7=��6=eT6=��5=�5=_4=��3=�+3=��2=
�2=Q^2=^H2=�(2=��1=�|1=D�0=\00=gc/=��.=�-=��,=�?,=i�+=�5+=�*=��*=v*=�S*=,*=J�)=��)=�)=W?(=�4'=W�%=�~$=��"=�o!=1�=&U=��==�=�=7�=�9=И=j�=�F
=��=j=�>=�8=��<Ő�<�[�<g��< �<���<��<g-�<p��<�I�<Y��<*��<0��<�J�<T�<���<ī�<���<eک<��<K��<�X�<���<ٓ<���<�4�<T��<�=�<f
z<ɹq<VFi<�s`<D#W<�SM<� C<��8<��.<7�$<�<Q<��<l�<�.�;��;���;^F�;3��;���;�
�;��u;�K;޲ ;x��:��:�"%:�m�8�t�mVz��6������J�,w?���b�M���Zח�
Z������ޭԻ����s��L2��]�s����t�%�R+.��c6�^H>�v�E���K�$Q��QU�َX�y%[�Z~]��_���b�d%f�ϴi��jm�kq���t��w���z�\�|�sy~������=2���/��='���1��'i��L值����4ꂼ�f�����ʎ��R舼�����Њ��q��� �����%j���h�����:򐼔R��s���Ѧ��+p������]P����������뗼���Ҕ���R��8��,�����ࣼx���Ӧ��`ʨ�2n��@驼�O������==��%���,���-V���������{����ص��x��!и��幼 Ϻ�0�������rɽ�C��ڡ��}>¼F�üHCż�pƼ�  �  2SK=l�J=P�J==J=�zI=��H=��G=��F=�F=:E=}qD=Q�C=C=�fB=��A=�0A=�@=�@=R�?=14?=2�>=M�>=F8>=e�==�e==3�<=�<=�=;=Hf:=�9=��8=(8=Vu7=��6=�M6=��5=�D5=��4=L^4=L�3=��3=Es3=�>3=�	3=~�2=�h2=�1=fC1=׎0=�/=�#/=�~.=�-=oa-=_�,=kk,=��+= �+=)+=�*=�H*=��)=3�)=�3)=��(=�+(=�a'=�Y&=!%=o�#=�"=�Z =Z�=��=b�=�=�\=�=��=�J=��=��
=J<=i=��=�=]1�<k��<W�<�$�<�(�<#$�<7#�<|+�<�<�<~Q�<�c�<�r�<��<��<�Ǻ<�<8��<�W�<H�<"^�<�<���<Lk�<��<yp�<ĺ�<j��<�1�<
�z<�_q<?�g<G^<}�T<�K<boA<,8<��.<�)&<��<)�<�8<đ<ha�;c��;K�; ��;���;�^�;�$�;K�w;h�Q;�+;6;;�s�:��X:��u9���7o��ľ�oq��="��_B���b��-�����r覻4���gλ7J�����<��������)����'�g�/��\7�W2>��SD�r�I��NN��GR�W�U�Y��j\���_�ȷc��yg��k�]_n��Mq�0�s�Xv��x�'�y��k{�n�|�0L~�^��=��[���7‼��� a��\ˁ��x���t������2�������戼�2��(c���|��?���\���}��
m��Q��u#���ܒ�z�����?������}˕��˖�Y�������L������Ꙟ���冡�ע�H���I��nt��ݔ��l���?�������G����������PW���>���m��z簼v���`��(��^ݷ�v��~�S��=���"龼�#��R���o¼�uü�]ļ�'ż�  �  �K=�IK=ȽJ=�J=� I=w#H=�$G=�9F=�oE=��D=�ED=��C=+fC=m�B=�XB=حA=��@=Q%@=�b?=��>=�.>=��==��==T==|==�<=w@<=��;=
�:=��9=��8=~�7=�7=w?6=S�5='5=��4=kJ4=i4=0�3=�3=��3=B�3=5N3= �2=n;2=�v1=��0=��/=�/=��.=�#.=��-=ȓ-=�M-=_�,=K�,=[�+=N+=��*=#�)=�Y)=��(=q(=d(=p�'=!'=�X&=�G%=6�#=�R"=�} =z=pS=G=��=}=.3=��=̾=̗=sz
=>a=�D=�=p�=x�<��<���<���<w��<���<	�<Ε�<6>�<u��<�[�<��<��<�u�<�.�<��<|�<�A�<���</�<	r�<��<�I�<�^�<_�<���<ᝇ<��<I�z<M�o<�e<=[<�SQ<S�G<��><bL6<y-.<�\&<{�<`<5(<��<w0�;u�;N�;��;g��;�N�;3ɋ; �u;�
T;2�1;��;I�:�m~:9��9"����_v��rʺ�-
�k3,��K�ץi��̓�U��������M��&˻�߻�������"H�
,��m"���*�ˊ2��G9��'?�1FD���H���L���P�:�T�r�X�)]��a��/f�LYj�_�m���p�4�r�'!t��=u��Rv� �w�g5y�*{�7a}�����‼����BI��/�������i���a₼�Z��w2��a���Ԇ��u��0+��R܋�s��8܎�A������Q���[-��c���������eL���ӓ�����\͕��S�����S���jƜ�]V��r�������h}���F��"$���+��@g��Ӧ�^���ꩼ1U�����Bi��|������� ���������+���������������������m��V��"t��ѕ���w¼S"ü�ü<ļ�ļ�  �  `�K==K=k�J=�I=#mH=<G=z F=T5E=l�D=�D=#�C=�C=��C=4C=��B=��A=nA=��?=��>=��==�>==��<=�<=~v<=Gt<=�\<=�<=&�;=��:=��9=��8=,�7=v6=`y5=�4=�4=S�3=5�3={�3=��3=�3=��3=��3=�53=��2=�1=��0=[�/=��.=�!.=��-=-=Ђ-=��-=�}-=�E-=��,=G',=�I+=cQ*=�[)=`�(=��'=�b'=�'=��&=��&=B�%=�%=�#=�C"=BV =O&=��=T=��=#|=/4=�=Q=�=5,
=�:=�0= ={�=9�<ӟ�<��<;��<�d�<���<Ok�<��<���<b��<���<1U�<wN�<���<��<�N�<ν�<���<i�<w'�<���<T��<�j�<8��<
	�<z��<���<�D�<�Fy<��m<�{b<��W<TyM<�D<��;<��3<��,<�z%<�V<Z�<ǭ<��<y�;���;]��;�P�;za�;��;�b�;�wo;!�R;̒4;�l;���:���:�]�9֪��톺G�޺�i���:�QZ�Qv��R���2��ٙ�����pʻE�߻����wN����R"�]�%��k.���5���;���@�1;E�lI���L�P�P�%�T���Y��#_�۰d�*�i��kn���q���s��u��au�'_u�?�u��Qv�q�w�Qz��g}��g������[���>�����������P�����_����l���_��F͆���������Ì��Ď�����ّ��Œ��E���h��FN��@!�����A��fۓ�H�'���3����Κ������՞��>��D*��%����.��}�������#Τ���������6��������G��nn������_���u�������#�� ��#���z����ʷ�}6��<���;޾�����E¼tQü��ü�:ļOPļ_ļ�ļ�  �  K=��J=(J=��H=��G=\1F=��D=HD=X�C=�GC=�JC=�hC=(wC=fNC=��B=%B=��@=1�?=�G>=M==Y2<=��;=�h;=t;=w�;=L�;=�;=sH;=��:=�9= _8=�7=��5=Y�4=6�3=K.3=�2=U�2=�3=O3=l�3=ה3=b3=��2=Y2=[�0=��/=)�.=t�-=�-=��,=I�,=	-=vS-=�~-=Ef-=�,=w,,=*+=r�)=��(=��'=&�&=�8&=F�%=�%=r�%=�d%=��$=K�#=�!=��=E�=�%=��=��=/{=�4="=�==x=Y�	=#�=��=̪=�(=���<���<u��<�6�<��<Iz�<D��<`(�<���<9��<��<��<͘�<���<��<uX�<TD�<���<���<���<&��<�ߙ<��<�<�y�<�-�<64�<�<�qw<{Dk<�I_<��S<��I<Z@<�68<�1<Ng*<4�#<%-<J�<J<_�<y�;y>�;�;�;�R�; �;��;�f;��N;�y4;V;���:���:���9g�˹���Z���&�Z�K���j��u��_��V����h��T���b�˻�%�mV���-����E��X)�1 2��9�g�>�.C�V�F��J��~M�rsQ��0V��[�pb�bh�M:n�g�r�D+v�S�w�.x�Bw�.1v�q�u�9�u��Vw�H4z�� ~�:J��7s���;��l��q솼Yˆ�:��J������6!��]؅��7��%��aq���፼+6���2������q����씼�Ȕ��X���ړ�
���c���G]�����������-���ʜ�,3������^��\󢼅���.����p��L���R5������������������>���F��٪���^���|��2@��> ��2��������������f��V���۽�h����¼�ļ�ż}�ż�~żR>żPż%ż�  �  �1K=:�J=�I=8<H=ɹF=�=E=m�C=)C=B=@�B=�B=�C=�PC=�KC=��B=E�A=C�@=�4?=�==�J<=k?;=��:=�f:=��:=g�:=7;={2;=b�:=�F:=�C9=��7=Y�6=�-5=x�3=� 3=�e2=�%2=k62=��2= �2=�/3=XI3=�3=4v2=�|1=�<0=�.=�-=��,=�
,=O�+=�,=̉,=	-=f-=Oi-=�,=R,=��*=�b)=��'=}�&=޿%=�.%=�$=��$=��$=x�$=�=$=�4#=R�!=��=�4=��=��=�#=I�=�\=+X=�=��
=�A	=I�=�=D=�� =Ht�<�<�<t �<s!�<]��<��<��<��<$�<H�<��<3��<h��<��<��<�U�<�ج<� �<#
�<��<�ښ<@�<�Ε<��<式<��<�<���<u<�h<+x\<��P<cQF<�#=<D5<Zy.<�U(<�H"<L�<�S<_�<Ԗ<���;�j�;VH�;��;Y;�;���;��s;^;��I;��2;l�;r��:%��:1L�9�F��� ���w��4�g�Z���y�k���K��:���֫��:����ͻ7f�2��+
��l��"�'[,��5��<��UA��LE�\pH�AZK�ߚN�/�R���W�}�]� �d���k��r� w�Qz�J{���z��9y��Iw�x�u���u��?w���z��#��:��l҄�����Xa������%ň�p ������8������~��g·�Ή�PG�������p���R>��)#���\��f��M\��!���T0��_B��o������a�����A��� 4���&��SJ��뛤��B������ܢ��G&��c���%ܦ������׬�v������(����h��i��=�G_�� ��9�������ؓ��#��+��u�������ļ��ż͝Ƽu�Ƽ�Ƽ�-Ƽ��ż�ż�  �   �J=�EJ=;.I=B�G=�#F=ŔD=�GC=bB=��A=�A=	MB=x�B=�,C=�?C=�B=>�A=��@=�>=Q6==S�;=d�:=A�9=\�9=$�9=�D:=B�:=��:=��:=q:=9=L�7=76=��4=�w3=�|2=?�1=��1=K�1=�2=��2=��2=�
3=��2=n"2=�1=��/=�B.=��,=!�+=}\+=�B+=A�+=�),=��,=K-=b-=I�,=��+=��*=)=�p'=�&=�%=zx$=?A$=�L$=�g$=�U$=��#=��"= `!=�Q=��=�!=T=)�=Z=��=��=J=�{
=��=8=�B=K�=�B =/}�<�<���<��<�z�<�$�<H��</��<�t�<���<���<���<?��<�p�<���<��<Oӫ<ɥ<W��<C��<S��<��<֔<�O�<�!�<��<��<t`�<4t<6<g<�Z<��N<A"D<Y�:<�D3<��,<��&<
!<Ĭ<<7<�R
<W��;���;A��;��;�G�;:��;1��;1.k;Z�W;VlE;��0;�o;�_�:g�:m	�9������(����>�0\e��$���R��Ӕ���������;_��,�ϻmK� q��r�,���#�~a.�s7���=��C���F���I�>`L�a�O�~�S��Y���_�E�f��Bn�B�t���y�=�|���}���|���z�J3x�QHv���u�Uw���z����-�Oυ�+������C^��7"���>��������������:K���T���茼���g��ѩ��>I���,��~V���於���`?��)�����������X��Uٙ��֜�"柼h�������ʝ���ƥ�=1��A2��#;���Ģ��.��������C������:Ѱ��\����� ϵ�w���?!��_��d볼% ��,������������ѿ�[�¼żo�Ƽ{�Ǽ��ǼW~Ǽ�ƼWMƼ�!Ƽ�  �  �J=!(J=C	I=��G=��E=�XD=]C=P#B=�A=}�A=T%B=b�B=�C=:C=
�B=�A=*y@='�>===��;=�[:=�9=jv9=�9=i:=�|:=ϱ:=V�:=�9=��8=��7=h6=l�4=FL3={N2=��1=�x1=��1=j�1=�o2=��2=��2=��2=�2=��0=g�/=�
.= �,=��+=�+=�
+=d+=,=�,=�?-=�]-=z�,=��+=͈*=m�(=B'=��%=��$=	8$=$=*$=�4$=c+$=�#=��"=[E!=r5=��=-�=(=Cj=��=\�=��=��=�V
=.�=H=�(=�= =�%�<���<�6�<�6�<���<���<B�<p��<�6�<���<E��<���<X��<'X�<�j�<�G�<�r�<6W�<�9�<F-�<%�<婖<<x�<��<<�<�ߊ<)�<�'�<�s<P�f<�Y<v�M<�_C<?:<Α2<`,<-N&<�� <�G<��<�	<���;�j�;���;��;V�;�Ɏ;��;�$h;�GU;��C;y0;C;uc�:�t�:�9iL���w��B�p-i����� ��S/��}������@���lл*��U����β�&�$��/���7��>�D�C�=`G��&J�o�L���O��T�G�Y��3`��g��!o���u�A�z���}���~���}�+D{�3�x�tv�L�u�
cw�{�o*��w6��1+������K5��9݊�@���Ұ���v��1f��a膼)>��5{�������$��<�������_��/�����������5��U]���y���䔼z��ӕ�0����.���=���Z�����K������1��T��� q���`���Ԣ��4��H����8���v��H���04���г������M��	8��ˎ��E���07���\���^���A���߹�}�	��üNkż�Ǽ�Ǽz,ȼi�Ǽ Ǽ�Ƽ�QƼ�  �   �J=�EJ=;.I=B�G=�#F=ŔD=�GC=bB=��A=�A=	MB=x�B=�,C=�?C=�B=>�A=��@=�>=Q6==S�;=d�:=A�9=\�9=$�9=�D:=B�:=��:=��:=q:=9=L�7=76=��4=�w3=�|2=?�1=��1=K�1=�2=��2=��2=�
3=��2=n"2=�1=��/=�B.=��,= �+=|\+=�B+=@�+=�),=��,=K-=b-=E�,=��+=��*=)=�p'=�&=�%=px$=6A$=}L$=�g$=�U$=��#=��"='`!=R=)�=�"=�T=K�=�=��=��=�=�~
=�=�;=G=��=G =3��<!�<յ�<���<ق�<�+�<���<���<y�<���<���<T��<C��<5n�<��<:��<nͫ<G¥<���<��<���<��<9͔<�F�<>�<��<��<AZ�<�)t<4g<L�Z<��N<
"D<� ;<J3<��,<�&<Y!<ۺ<�F<�c
<Z <��;���;0�;�i�;�Ӑ;֮�;�_k;Q�W;��E;z�0;�y;�]�:Nڏ:�Q�9�$�uv��s���>���e��H��,x��[����⢻ ���N���|�ϻl廐�����\"�<�#�wj.��#7��>�� C���F���I�}bL��O�έS��Y�W�_���f�Cn���t��y�o�|�ڻ}���|���z�[3x�^Hv���u�Uw���z����/�Qυ�+������C^��7"���>��������������;K���T���茼���g��ѩ��>I���,��~V���於���`?��)�����������X��Uٙ��֜�"柼h�������ʝ���ƥ�=1��A2��#;���Ģ��.��������C������:Ѱ��\����� ϵ�w���?!��_��d볼% ��,������������ѿ�[�¼żo�Ƽ{�Ǽ��ǼW~Ǽ�ƼWMƼ�!Ƽ�  �  �1K=:�J=�I=8<H=ɹF=�=E=m�C=)C=B=@�B=�B=�C=�PC=�KC=��B=E�A=C�@=�4?=�==�J<=k?;=��:=�f:=��:=g�:=7;={2;=b�:=�F:=�C9=��7=Y�6=�-5=x�3=� 3=�e2=�%2=k62=��2= �2=�/3=XI3=�3=4v2=�|1=�<0=�.=�-=��,=�
,=M�+=,=ɉ,=-=�e-=Ji-=x�,=J,=��*=�b)=��'=m�&=Ϳ%=�.%=
�$=��$=��$=w�$=�=$=�4#=��!=A�=k5=َ=)�=�%=&�=�`=�\=@�=|�
=�H	=��=�=KL=J� =���<aN�<��<�1�<���<��<^��<h��<G&�<�M�<N��<���<���<n��<��<�L�<dͬ<��<p��<���<7ʚ<�.�<���<��<Ȭ�<��<I��<��<��u<m�h<Wm\<!�P<�PF<�(=<%N5<`�.<?i(<�`"<��<+r<��< �<�'�;9��;&��;h'�;�x�;�ކ;n$t;k^;��I;��2;ž;���:�|�:��9�K���ǩ�����(5��W[��Qz��������焟�� ��e���;λ���l���(
�D���"�wl,��5�|<��^A��SE�vH��^K�8�N���R���W���]��d�^�k�Wr�~w��z�UJ{���z��9y� Jw���u��u��?w���z��#��:��n҄�����Ya������%ň�p ������8������~��g·�Ή�PG�������p���R>��)#���\��f��M\��!���T0��_B��o������a�����A��� 4���&��SJ��뛤��B������ܢ��G&��c���%ܦ������׬�v������(����h��i��=�G_�� ��9�������ؓ��#��+��u�������ļ��ż͝Ƽu�Ƽ�Ƽ�-Ƽ��ż�ż�  �  K=��J=(J=��H=��G=\1F=��D=HD=X�C=�GC=�JC=�hC=(wC=fNC=��B=%B=��@=1�?=�G>=M==Y2<=��;=�h;=t;=w�;=L�;=�;=sH;=��:=�9= _8=�7=��5=Y�4=6�3=K.3=�2=U�2=�3=O3=l�3=ה3=b3=��2=Y2=Z�0=��/='�.=s�-=�-=��,=E�,=	-=qS-=�~-==f-=�,=k,,=+=a�)=��(=v�'=�&=w8&=-�%=�%=c�%=�d%=Ĵ$=��#=��!=�  =d�=k'=�=��=<=�9=9(=E=h�=��	=c�=��=t�=�4=I��<k��<��<�M�<�<��<���<�6�<��<Z��<x�<���<��<h��<O��<oK�<W4�<��<��<O�<���<�Ǚ<��<2��<&c�<��<� �<��<bUw<o.k<�:_<��S<�I< a@<�D8<�1<�*<�$<�S<�<x<��<%��;ɡ�;Ol�;�z�;m��;P�;�7�;�Mg;��N;f�4;�-;$��:
x�:\��9	�ι®��Pw��O'��^L��nk�f܂�NȎ�A���LѨ�����̻��w����R��1��b�q)��2�/9���>�z8C�s�F�J���M�wQ�|3V�*�[�b�Lch�8;n��r��+v���w�}x�@Bw�\1v���u�S�u��Vw�W4z�� ~�?J��;s���;��l��s솼Zˆ�:��J������6!��]؅��7��%��aq���፼+6���2������q����씼�Ȕ��X���ړ�
���c���G]�����������-���ʜ�,3������^��\󢼅���.����p��L���R5������������������>���F��٪���^���|��2@��> ��2��������������f��V���۽�h����¼�ļ�ż}�ż�~żR>żPż%ż�  �  `�K==K=k�J=�I=#mH=<G=z F=T5E=l�D=�D=#�C=�C=��C=4C=��B=��A=nA=��?=��>=��==�>==��<=�<=~v<=Gt<=�\<=�<=&�;=��:=��9=��8=,�7=v6=`y5=�4=�4=S�3=5�3=z�3=��3=�3=��3=��3=�53=��2=�1=��0=Z�/=��.=�!.=��-=��-=ʂ-=��-=�}-=�E-=��,=9',=�I+=OQ*=�[)=E�(=e�'=db'=�'=��&=��&=A�%=�%=_�#=D"=*W =�'=��=�V=��=�=e:=e=0=�=�7
=�G=P>=d=L�=e6�<���<s#�<���<G�<���<���<��<��<T�<���<_V�<*K�<���<��<?�<G��<ֈ�<��<�<Л�<�u�<�L�<ٔ<�<bz�<��<0�<$y<��m<Mib<��W<�xM<'D<�;<��3<~�,<k�%<ƅ<�<2�<��<ܕ�;��;O�;5º;˧;�y�;W��; p;>S;t�4;s�;��:�O�:���9dR������ຈ1�5�;�
[� w�oӈ�d���������T�ʻ��߻�A��I|���|E�@�%���.�>�5���;��A�>EE�,I�q�L�ԣP���T�`�Y��%_�Z�d�M�i��ln�g�q�=�s�0u�<bu�__u�j�u��Qv���w� Qz��g}��g������[���>�����������P�����_����l���_��G͆���������Ì��Ď�����ّ��Œ��E���h��FN��@!�����A��fۓ�H�'���3����Κ������՞��>��D*��%����.��}�������#Τ���������6��������G��nn������_���u�������#�� ��#���z����ʷ�}6��<���;޾�����E¼tQü��ü�:ļOPļ_ļ�ļ�  �  �K=�IK=ȽJ=�J=� I=w#H=�$G=�9F=�oE=��D=�ED=��C=+fC=m�B=�XB=حA=��@=Q%@=�b?=��>=�.>=��==��==T==|==�<=v@<=��;=
�:=��9=��8=~�7=�7=v?6=S�5='5=��4=kJ4=i4=0�3=�3=��3=B�3=4N3=��2=m;2=�v1=��0=��/=�/=��.=�#.=��-=��-=�M-=T�,=>�,=K�+=�M+=x�*=�)=oY)=��(=�p(=B(=S�'=� '=�X&=�G%=��#=!S"=�~ =�{=�U=~=*�=��=:=�=��=%�=0�
=>o=�S=�+=��=#�<h'�<���<|��<���<���<� �<���<�M�<���<b�<Z��<4��<�l�<Y!�<�<�ٰ<�(�<_ݧ<��<�Q�<�˜<�(�<q>�<0��<ec�<y��<�l�<�hz<U�o<ke<�2[<�RQ<��G<��><)i6<S.<m�&<�<�B<)g<'<Է�;��;ҝ�;o�;��;︝;"%�;�>v;�~T;��1;�;�A�:��}:��9W�����x�f�˺�*-�ܹL�M�j�Y]��-���O��7ط��˻X*��8���%�Hu�2S�َ"��+���2�Z9�%6?��QD���H���L���P��T�b�X�c]���a��0f�EZj��m�C�p���r�z!t�->u��Rv�D�w��5y�%*{�Ga}�����‼����EI��1�������k���b₼�Z��x2��a���Ԇ��u��0+��R܋�s��8܎�A������Q���[-��c���������eL���ӓ�����\͕��S�����S���jƜ�]V��r�������h}���F��"$���+��@g��Ӧ�^���ꩼ1U�����Bi��|������� ���������+���������������������m��V��"t��ѕ���w¼S"ü�ü<ļ�ļ�  �  2SK=l�J=P�J==J=�zI=��H=��G=��F=�F=:E=}qD=Q�C=C=�fB=��A=�0A=�@=�@=R�?=14?=2�>=M�>=F8>=e�==�e==3�<=�<=�=;=Hf:=�9=��8=(8=Vu7=��6=�M6=��5=�D5=��4=K^4=L�3=��3=Es3=�>3=�	3=}�2=�h2=�1=dC1=Վ0=	�/=�#/=�~.=�-=ha-=V�,=`k,=��+=�+=+=�*=�H*=|�)=�)=�3)=l�(=�+(=�a'=�Y&=D%=ǥ#=_"=�[ =�=��=��=x�=�b=�=2�=,U=h�=(�
=�J=	=E�=9�=5T�<3��<`(�<;E�<%G�<�?�<�;�<�?�<)M�<�\�<Tj�<#t�<1~�<��<��<��<���<�=�<�*�<�>�<�_�<�m�<�H�<��<+P�<���<܆<��<(�z<�@q<��g<�;^<��T<oK<T�A<�$8<�/<�X&<z<�%<�y</�<���;�A�;]��;��;I�;̢;��;0�x;~ R;�Q+;b;-l�:��W:0qp9���A�q��T��cW��<#��rC���c�R�����~|�����7�λ��JZ����y�x�����(��0��o7�oA>�z_D���I��UN�)MR�h�U�&Y�9m\���_��c��zg�Gk��_n�%Nq���s��v��x�L�y��k{���|�@L~�j��=��^���:‼���"a��]ˁ��x���t�� ���2�������戼�2��(c���|��?���\���}��
m��Q��u#���ܒ�z�����?������}˕��˖�Y�������L������Ꙟ���冡�ע�H���I��nt��ݔ��l���?�������G����������PW���>���m��z簼v���`��(��^ݷ�v��~�S��=���"龼�#��R���o¼�uü�]ļ�'ż�  �  ��J=�EJ=�J=��I=�gI=%�H=�+H=�QG=]F=RZE=�UD=k[C=�uB=5�A=~A=�|@=s@=��?=Ӑ?=�_?=�*?=��>=��>=��==�C==�f<=�s;=�:=>�9=��8=�i8=��7=M�7=u@7=��6=eT6=��5=�5=_4=��3=�+3=��2=
�2=P^2=]H2=�(2=��1=�|1=B�0=Y00=cc/=��.=�-=��,=�?,=^�+=�5+= �*=��*=v*=jS*=�+*=*�)=x�)=�)=;?(=�4'=Z�%=$=�"=wp!=@�=�V=�=A=#=K=�=�A=��=��=�S
=��=y=�N=5I=���<_��<�|�<���<��<��<���<7A�<��<�T�<��<}��<��<:B�<Թ<ߞ�<��<���<<��<L¥</��<�7�<Ϗ�<븓<�ڎ<��<ބ�<�&�<��y<ӛq<�1i<�h`<{"W<�\M<�3C<F�8<+�.<��$<��<��<��<��<e��;^�;&�;���;��;u#�;�f�;Kv;�wK;� !;��:��:�m$:緓8�W��|�︾��B���@���@�ϙc��!h��)鬻�\��2ջ<�_���\e�����Ź�6�%�B.�4v6�W>���E���K��*Q�1WU�ӒX�|([���]�� `���b�b&f���i�vkm��q��t�S�w�Ěz���|��y~�-�����C2���/��A'���1��)i��N值����5ꂼ�f�����ʎ��R舼�����Њ��q��� �����&j���h�����:򐼔R��s���Ѧ��+p������]P����������뗼���Ҕ���R��8��,�����ࣼx���Ӧ��`ʨ�2n��@驼�O������==��%���,���-V���������{����ص��x��!и��幼 Ϻ�0�������rɽ�C��ڡ��}>¼F�üHCż�pƼ�  �  T�I=iBI=�!I=nI=��H=ȪH=_ H=,WG=pXF=�3E=��C=R�B= �A=2�@=@=��?=�_?=�F?=�D?=�B?=~*?=,�>=Ap>= �==��<=�;=�:=�~9=��8=�8=��7=g�7=m�7=�h7=i#7=w�6=Z�5=Z5=""4=�03=?c2=�1='z1=b1=�r1=��1=�1=nX1=��0=�50=V/=EW.=N-=�P,=�t+=��*=�P*=�*=��)=-*=�*=
*=��)=|�)=��(=?�'=o�&=�*%= �#=0"=� =�)=��=��=d=t=z=P*=��==�=��=1�	=�=ޒ=#_=)m =�K�<)��<��<���<�>�<I�<@��<���<���<���<O�<��<�<,��<E��<kô<%�<�v�<맩<���<��<9H�<F$�<��<`Ȍ<1 �<���<n`<!x<� q<G�i<�a<G�X<p�N<��C<Y�8<�@-<�i"<��<��<30<׆<ˢ�;���;��;���; I�;���;��;�Qp;��A;�";���:�~~:��9���p��s��*�ź�� ��� �N1C�� i�d-���잻ᴻ�ʻE�ݻ4q�`l��@�,�\����}�$�lf-�Ii6�l_?���G��O�EU�J�Y�ޗ\�Б^�� `�ka�y�c��;f���i��m���q��Uv�7az�t�}�Q4��E
���j��#d��D��ئ���I���)��*j���$��c������l������!ۊ�e����?��������0��g�'ȍ�?�����%���ZՔ��[��n��q���4���*���+���{���C��Ɏ��tO��$j����������A���%���������*R��C���¥��h���[Ǫ��1��1��=X���)��/_�����*����巼�T���F��XӺ�c(�����m�����4����h����¼��ļ?�Ƽ�Cȼ�  �  }qH=8!H=�H=�7H=QH=>:H=��G=P!G=F=��D=C�C=�'B=�@=��?=K/?=��>=��>=�>=m�>==�>=��>=�>=� >=y<==)<=��:=�u9=-[8=��7=�7=:�6=�7=&H7=�b7=�A7=��6=�6=��4=A�3=�2=�{1=$�0=PV0=zF0=w0=8�0=��0=U�0=d�0=
0=�/=��-=��,=N�+=U�*=��)=&h)=R9)=H)='~)=��)=o�)=�)=�b)=��(=�m'=��%=l>$=<�"=�� =�=M=<=12=?=/�=>�=�a=G�=Ώ=�U=j&	=z.=�=�N=)��<e��<qy�<Q)�<�X�<h��<���<P�<4��<���<%v�<��<% �<�@�<��<�$�<I��<�T�<��<V!�<3�<�.�<�<�b�<�ʏ<�|�<���<劁<��{<ԯu<��o<�mi<m(b<�Y<^O<��C<�7<�6+<	]<
�<��<��<�3�;s�;F�;Zw�;�|�;��;��;�[�;�Rh;F�6;��;+�:�?:�6,9m:��B8L�j���ZҺ���%��uI�1r� K�����ҽ�!�ӻ���u�������8	� �	J��;��:$�MB-�h7��A��J���R�KoY�F+^�Za���b��9c���c�7e��Cg�6�j���n��}s��xx��-}�6������k߂�����т��-��Qm���Ѐ����值�݁��}������C����'���狼����u��9S��z׌�T��{��5z������o@���~��l����V���K��/����M���[��b��7���^~��-뙼���W���U���_���<�������਼�z��"}���o꫼ҡ��HT���?��E��������.��i�����'ǵ�_=��$*���i������/���ջ�C�����#м��]�������%üN�ż5VȼSPʼ�  �  �nG=�G=�&G=fG=ĨG=]�G=�yG=`�F=!�E=8�D=�
C= �A=C9@=^%?=�f>=>=��==�>=�a>=��>=̦>=�a>=+�==Ҵ<=K`;=��9=.~8=�U7=��6=�46=p>6="�6=-�6=�C7=�B7=��6=��5=b�4=-M3=
�1=6�0=�/=#Q/=�F/=��/=�/=�_0=ׄ0=O0=׵/=��.=��-=�C,=`�*=��)=�)=��(=6(=�(=�(=�T)=��)=A�)=�)= 0(=��&=Q6%=�a#=��!=��=�=�~=��=��=�=�=��=v=��=�W=j�===�[=~�=�W =k��<���<K#�<�%�<ϛ�<�O�<66�<"h�<��<S��<!�<��<��<C��<�z�<ݵ<���<,~�</�<lt�<�!�<�&�<u��<Ź�<!�<�n�<���<L<�x<�Ms<�Bn<z�h<V+b<��Y<zO<�zC<�g6<X)<�q<�(<��<� <#��;���;r��;ӧ�;���;�J�;맠;�N�;�f`;2-;���:���: w	:�3�i�Y�t�\���w�ߺ����s+�w�P�ic{��>��lӭ�q�Ż��ۻ�(�������p��s�y���G��+$���-���7���B��'M�3V�BW]�Lb�� e�A=f�8Uf��If���f���h���k�O p�u�M�z�+��������<o��Ò��9���;���@��ix���*����������)�����Y����#���򍼹����+������C��Ќ�SB��$n��ဍ�u���������@Ǘ�q��!����X���O������%
����������(����S��M����o���W��$���^��������X��� ��6���?��ޫ��4��LG��$�����J���S����B���1���L�����)A���������.��ο��f��L�����üǼ��ɼ�,̼�  �  9�F=
kF=�~F=]�F=P-G=�YG=O-G=�F=z�E=9D=��B=%A=ӿ?=+�>=��==a�==2y==�==Z>=OV>=h>=�>=�k==�M<=�:=UM9=��7=��6=��5=ғ5=?�5=D)6=F�6=�$7=�97=g�6=�5=7�4=��2=�e1=�0=�/=�.=��.='�.=xq/=z�/=9+0=�0=Mw/=K�.=�D-=��+=��*=�j)=G�(=�(=U(=_4(=%�(=F)=�M)=�E)=q�(=�'=�r&=��$=|�"=x� =�D=�=��=�'=�y=A�=|�=��=!y=3�=�%=�=�=��=��=3Y�<��<���<|'�<]�<, �<���<���<���<�v�<`��<?6�<�<Pv�<^��<|�<���<�ޱ<8ݮ<բ�<��<���<]_�<٠�<Q��<���<X�<X@�<ݯ|<܃v<��q<�m<49h<�b<	�Y<(cO<� C<'c5<v�'<Z<��<<�<ئ�;���;L�;74�;Y��;,H�;G�;A��;4��;R�Z;B&;T��:):�:���9@�.��%'�Ԓ��/�h�����'0��<V��'��E���9Ѳ�Md˻���	�����81�%�v���]�ys�0D$�[�-���8��)D�-O�#�X�&`��e���g���h���h�Ch�^Oh���i��l��
q��Vv�&	|���������Uz��m�������r���7������ߧ��R��+j��R����0�� �����iY���P���^�������u��w:���n��hx��Ə��`���b���;����Θ�}O��i��������������a��Cj���_��i)���Н�R5��_���!������Y`��"������M��t����Q�������^��ճ���ܭ��᯼꠲�q˵��<���&���񚾼˹��|$��X5��Ga�����dǼ�����)���pļ��Ǽ-˼:wͼ�  �  �zK=9K=��J=U�J=�J=UkJ=8�I=��H=��G=�hF==�D=JrC=b B=�A=P@=��?=��?=Q�?=�7@=hz@=I�@=́@=�@=�a?=�g>=�F==`%<=B,;=�w:=:=��9=�:=�<:=iS:=�/:=p�9=��8=��7={�6=�b5=P4=T3=�2=>�2=0�2=,�2=��2=�2=�2=G1=�*0=z�.=$�-=09,=�+= D*=��)=��)=��)=��)=�'*=F_*=�`*=�*=oc)=bV(=�&=�l%=��#=�N"=D� =��=��=��=V�=:=�r=N9=��=�=Ԅ=�p=�=#�=R�=J�=Y��<�]�<���<�}�<���<2<�<�=�<i��<�q�<�#�<55�<=��<T�<�	�<&��<�]�<_�<J�<2�<N	�<���<���<���<�A�<}1�<���<J��<�
�<��<��{<��u<��n<�,f<f=\<�Q<��D<t�8<2-<I"<�<��<�	<E�<�'�;���;�7�;���;��;K�;6݀;T O;�6;w{�:���:��:S��8����|5�Za���8��g����TkA���j�Q銻����ܴ��ǻ|�ֻQ{��g�s���{��E
����մ��?$�.��[7��?�*|F�+�K��%O�jQ�US���T�s�V�[ Z��)^��8c�^�h�0�n�Z�s�z]x�֩{���}��~��j}�8�{��"z��x�7�w��w��y���{�cH���������������iz��UX���煼�p��UD�����;���!|��2���%;������॑�"������Z���^���^��'���uu���䖼���� ����b���K�������B��	5�~G���������R�����{ǧ�j����������˭�d)��T������!���������x|���]������&}��m���=��Gּ�8����	¼|ļ�  �  ��K=�6K=K=��J=w�J=��J=��I=I=��G=$F=nE=Z�C=FB=�7A=�y@=�@=��?=B@=�Q@=�@=��@=`�@=�/@=4|?=�>=k==�M<=�U;=x�:=6:=>:=>":=(C:=�P:=�':=��9=��8=��7=�6=z5=�o4=b�3='3=3�2=u�2=� 3=��2=��2=�12=9Z1=�>0=A�.=B�-=�[,=�B+=m*=��)=��)=��)=p�)=�?*=xs*=ds*=?%*=�y)=cq(=�'=`�%=��#=Kv"=�!=%�=��=��=��=52=�f=-=��=D�=��=��=�==A�=Q�=l
 =���<���<���<���<Z]�<�c�<��<ͭ�<:k�<��<y)�<�p�<�Y�<�˹<���<Ò�<xx�<z�<U:�<Iۤ<��<�՚<���<)��<��<�؇<�I�<��<J|<��u<�n<hf<5\<��P<�E<s�8<�i-<��"<dr<�i<tr
<b<�;t��;l��;�p�;���;���;洁;�7Q;=� ; ��:�r�:�:��9O���|-�h!��%:��b�'e�I}?�6Lh�V���J"���s����Ż�ջ<��*�ﻴ]��Ѭ��]
��H��3$���-�o�6��&?�*�E�o�J�vN���P�!R��6T�o~V�_�Y�+�]���b�@uh��n��Ss�:�w�v{���|�Qx}���|��z{��y�/x�gBw�D^w�=�x��E{���~�E[��B���̄��̅� 9��(��I̅�_j���M��M���qʆ������������Bj��Ra��:Ӓ�����	�������Wr��aH��8���Θ�g[��30����T���������X���7���zڨ�l���駼/������ @��g��:P������,ۯ���������״��f�������h��i]������
���C��%?���ļ�ob�������ü�  �  �L=ҩK=stK=�TK=�&K=~�J=E+J=[BI=�H=ھF=XSE=��C=2�B=f�A=��@=7�@=#^@=Sn@=-�@=1�@=��@==�@=�l@=�?=��>=�==ƽ<=��;=V;=��:==\:=�N:=�Q:=TF:=::=�9=�8=/�7=��6=Ͷ5=��4=	4= �3=�d3=�\3=7_3=�H3=~�2=�i2=%�1=x0=(;/=.�-=��,=��+=��*=�\*=�!*=�#*=VM*=R�*=�*=��*=�Z*=��)=��(=�s'=+�%=0g$=y�"=-!=�< =�=��=6�=�=�A=x	=�v=��=��=e�=P�=�t=�6=�:=i =8�<�_�<��<91�<%��<X��<Y��<�Z�<�7�<fi�<*�<D_�<�:�<F��<�E�<�!�<_��<���<Ի�<�q�<��<���<�z�<�w�<~ӌ<.��<�<���<�y|<w�u<>n<�{e<�[<I�P<�CE<H�9<��.<"9$<=<<\<ny<9u�;��;���;;�;�7�; ��;�.�;�:W;��';B��:	�:�;:7w9~�F��\��i|��0��d`�c��TX:�wBb��1��Oc�������"»3�һ��@����� ���
�w���!$��L-��6�y�=��7D�N+I���L�_O�� Q���R��sU�G�X��]���a��bg�l�l���q��v��.y��{��{�ZM{��&z�D�x��Fw��mv�r�v���w�z��P}����A^���烼y���񆅼7��������_��\o��v����@��������Ȍ�2ގ�-��������ɒ�$(��!F���k���ݓ��̔��P���b��O㚼n���U\��u碼������ʲ��x"��@���̧�Pg���"���6���̧����������¬�j ��y��vղ����ô�����7���c��[ص�ɶ��I���J��q�������1��uü�  �  ^�L=NL=L=��K=��K=s*K=�zJ=��I=4dH=>G=4�E=y{D=VPC=�WB=�A=S-A=K�@=��@=�	A=f%A=L0A=A=ھ@=�)@=!Z?==b>=^==m<=��;=�;=;�:=\�:=\:=|+:=��9=o]9=��8=��7=��6=�6=;5=a�4=U:4=�4=A�3=��3=�3=�U3=��2=U�1=��0=H�/=�n.=�O-=�T,=�+=`+=��*=�*=g�*=J�*=;�*=��*=�*=2*=#)=��'=��&=~%=w}#=�	"=C� =�X=H =��=Y�=��=Q�=�I=
�=��=�=�l	=��=}�=��=�� =f�<��<��<���<LC�<Ft�<n�<�[�<�h�<���<[�<8��<K��<꽻<>B�<��<¤�<�/�<�k�<!@�<�<=ɜ<���<K˒<��<�ŉ<�ʅ<A�<��|<tWu<�Rm<N�d<��Z<8LP<:eE<oz:<��/<w-&<3Y<!}<`]<v�<�s <�\�;��;�-�;���;n��;m܇;U4`;%�1;\J;/i�:D�h:���9/vJ�Dd򹢄b��򦺶f�>���33�ĿY��J����W3�� ��=λz�ݻ�`�^I��� ��o��B�����3$���,�|�4�<�;�1�A���F�mJ��L���N��3Q�GT�̔W���[�<�`���e���j��}o��qs��qv�@Vx�! y�w�x��/x�@w�:�u��Ju�Uu��Wv�W_x�	E{�#�~����!����Ѓ�j���a���9��%f������I[��/g���؈�U���g��'��Y���Eɐ������呼����o������$�����8ϗ��6��Ȝ�wV��e�������N��LX��o়����ᦼ���B��������0��?;���é�%���#ȭ�Jӯ�l������t과s����������t1���7��/����q��:s��U}��p`��=����  �  9WM=?�L=�L=muL=�L=
�K=��J=K�I=��H=>~G=sGF=#E=1D=#C=pB=��A=�A=ʍA=��A=v�A=#yA=�VA=NA=��@=��?=��>=
>=�==�I<=n�;=�;=��:='Q:=��9=�9=�9=�f8=��7=	�6=0I6=u�5=�65=@�4=R�4=?�4=ao4=K%4=��3=��2=22=�1=�
0=L�.=u�-=�-=�],=j�+=�+=�b+=�V+=�U+=.N+=�-+=��*=xX*=�)=pq(= '=ߧ%=�$=+�"=9!=̔=.=�a=%�=��=`=��=Nu=��=�P=��	=Z�==j=�k=N|=��<���<�*�<=$�<���<�<�Q�<x��<���<&O�<C'�<ih�<��<��<na�<sյ<�Y�<{ή<��<�
�<���<#��<�<u8�<�t�<�<���<�~�<y�|<y�t<�l<��b<,_Y<�_O<2-E<;<L1<'%(<q�<<~�<Z�	<=.<��;���;"*�;��;��;y�;(�j;5;>;л;�-�:mh�:Ƹ:˭�8�����cF��n��,�պ�	
�� ,�[�P��x�bB���W��������ɻ��ڻ���Vj�����S��ȑ���m�$��g,�$�3�:��}?�?�C�LMG��J��L�CpO��R�xV���Z�sg_��d�/�h�t�l�vhp�&6s�#u�$v�Dv���u��Qu���t�M6t�Ct�*u�5�v��%y�_/|�Ou��H��3���o����n����˛��]=��t
������N�����L"���|��ץ��l���K$��󊐼j琼�l��E��(����7��@��f����ڛ�~)��[O���/������;����e��۹��إ��ݥ��ꥼ� ��j���s���|ڨ�?���z��s���E��-Ա�����������յ��ȶ�n근�C���ͺ�s�����䖿������  �  ��M=ΓM=�FM=��L=�hL=��K='�J=�I=��H='�G=L�F=��E=y�D=��C=�FC=�B=�cB= B=�A=��A=n�A=�vA=�1A=y�@=�3@=�u?=��>=�==��<=�<=R;=��:=":=�9=D9=g�8=��7=�o7=+�6=�m6==6=d�5=�w5=�K5=j5=��4=�n4==�3=3=
?2=`S1=/d0=�z/=R�.=$�-=�0-=d�,=N,=,=��+=�+=��+=0O+=��*=�~*=��)=��(=И'=Q0&=�$=E	#=�a!=��=��=�=�=�=(�=�=i*=	�=ep=�)
= �=Q�=��=��=��<�)�<)a�<UL�<���<x��<��<ޙ�<�/�<���<f��<C�<���<l�<qj�<r��<hڲ<-�<Tr�<���<�c�<9�<TD�<Nq�<q��<�ڋ<�7�<��<�S|<�Es<�j<}�`<HVW<��M<�^D<�;<E"2<_�)<��!<�"<S�<�I<V<{�;���;��;rm�;�=�;uҏ;"�t;��J;�!;��:b[�:��K:�͐9�#V�`:/�E��NϺ�[��'��J�guo�P��E������0ƻ
�ػ�j껥����;�<u��z�Z;�M�%�)�,��2�;�8��}=�b�A�O�D�T�G�N�J�s>N���Q���U��/Z��}^�+�b�H�f��3j�kUm��o�H�q�'�r���s���s��s�D�s�i�s�|�s�	[t�K�u�Ӎw��$z�5&}��"��ם����������#����������
��w������!��b���ݍ�(�����mh��q폼2����ő�q7��b�������t��F��l잼������f��<飼�|���礼:�����]ݥ��\������9��۫��Of��H��)���갼����과7���s�������븼.��Cu��B�����S
�������  �  �;N=��M={�M=�M=�|L=�K=�J=`�I=��H=��G=�
G=B4F=�kE=ٲD=�D=~C= C=��B=94B=�A=��A=�\A=A=��@=�N@=z�?=��>=I>=�%==v<<=�\;=�:=��9=�9=�m8=��7=�e7=��6=�6=Ib6=�(6=>�5=��5=_�5=�e5=z5=�w4=;�3=@�2=B,2=�[1=��0=��/=y*/=�.=��-=q-=8�,=c�,=�;,=��+=b�+=5:+=��*=/e*=��)=��(=��'=Q~&=K�$=�E#=Qz!=,�=k�=��=�q=�E=+=��=s�=ӄ=_=sE
=�8=5=.=�=��<D	�<��<��<��<���<���<q�<Ya�<a_�<at�<���<��<���<�-�<i��<���<7�<iX�<���<ӛ�<�j�</�<A:�<"X�<@d�<�m�<)z�<&{<hCq<��g<��]<ʩT<}�K<:�B<�^:<�22<�[*<��"<^<��<W�<�{<R��;`��;?E�;�]�;�i�;��;�D};�U;X�.;R;t:�:ƾx:�!�9���N�"�g���zϺǁ��&��9G���j�f.��2䛻����$Ļp�׻zd�A���8�a������y �2R'�/�-�3�88�UG<��@�lC���F�ZCJ��N��R�oQV��qZ�5T^���a��e�z h���j��l��n�''p��Vq�Gr���r��s�7�s�@0t�5�t���u���v��y�K�{�j�~����g����%�����������1��OS���N��%���݋�\}��B��y��G܍��>������Ao���q��lǑ�!d���-�����Ә�c���0��8����(��u��+��������w���=���뤼�����	��F���&8�����iI��@ʪ���� v��yf��hJ�����J̵�yf���⸼�:���h���p���Z���)��'߾�}���  �  �SN=�N=��M=LM=�EL=VbK=�nJ=_I=��H=��G='*G=@�F=��E=BQE=�D=ND=$xC=��B=�GB=��A=XA=tA=�@=�w@=M@=C�?=�>=b+>=�:==`9<=u3;=�3:=B9=g8=��7=o7=��6=�h6=�=6=�$6=�6=�6=��5=ݼ5= e5=��4=�64=Kp3= �2=��1=Z+1=i�0=�	0=�/=E/=ݖ.=&.=U�-=��,=�o,=d�+=�_+=&�*=�x*=*=�x)=!�(=��'=��&=�%=�E#=�Z!=�L=^$=.�=E�=�j=l;=�=�=E==�(
=v7=s<=�*=o�=�C�<UW�<�E�<�0�<	3�<*X�<X��<w��<BE�<���<h��<���<�#�<P�<���<��<���<I��<���<T��<�>�<�L�<��<Jx�<Ǔ�<�v�<#6�<��<�)y<��n<Ipd<�Z<ryQ<��H<ƭ@<a�8<�n1<?(*<@�"<.�<Y�<�g</{<�&�;���;�{�;(~�;��;���;K��;<z^;L^9;	�;���:O��:�:q��TL$�K�����׺ �t�)��I���j�,K������#�����û%�ػ�����7�
���� �A#�ƙ)�p$/� �3��88�(<�)�?�=C�e�F�,�J��O��qS�N�W��[�a_��a�{Sd��of��_h��<j�;l�K�m�޳o��kq���r��1t�Bu�Q�u��v���v��w�0y��m{��c~��瀼����T���~d����5���Pފ�oՋ���������6��c������6�������������*ɐ�H[��d���䕼@���D��Fq��׫���՜�����'���W������Ƣ���+���󥼣���"O���ߧ������{������-\��FC���X��t���c����������8[���Ȼ�T弼Y����P���þ�N��qu���  �  3N=D�M=�gM=�L=��K=Y�J=?�I=��H=3H=��G=�G=ǭF=�AF=��E=�5E=0�D=��C=W�B={,B=�vA=y�@=s@=�'@=�?=ʰ?=�T?=��>=�	>=�== <=��:=�9=Z�8=3�7=�6=5B6=��5=5�5=Ա5=)�5=��5=��5=-�5=�5=�#5=�4=&�3=1�2=�2=�W1=<�0=-^0=0=��/=hu/=\/=֑.=��-=�:-=Cv,=^�+=D�*=c*=��)=�k)=�(=QQ(=`v'=O&=�$=�#=�!=x�=��=>+=��=ɀ=�R=�F=X=F}=a�=v�	=� =	=��=�=9O�<�.�<E�<`��<�,�<���<�N�<��<���<�p�<���<G��<��<6��<��<���<�<Җ�<���<���<c�<W��<��<y8�<�[�<@!�<�<��<��v<�k<)a<&W<iN<2�E<)><n�6<� 0<�0)<72"<��<�<=�	<�� <���;��;��;��;d�;qc�;�;\�d;7�A;��;^�:��:��:�ꥸ�G2�M���D�,��0�3�N��}n��q���L�������;Ż�Vۻ�p�q{�A��v��D��U&�E,��@1��y5�)9��<���?���C���G��+L��P�ŮU�Z�ǰ]��`��b�Dd���e���f�JHh�xj��Il���n�_Gq�Y�s�k�u��w�v�w�*Xx��x�Ay�0z�5|���~�M4���6���V���s��Jn���)��z����|��H���9��V4�������������I�������[���4h��YF���������ݽ�����$����F��X ��!'���f��ڠ�<n�����e���ɦ��ŧ��y������[~���.���5����������m������񁵼d᷼��:���+v�������*������ܦ��C���"ӿ��  �  ��M=j�M=�	M=�8L=n;K=�+J=$)I=*NH=5�G=�5G=��F=r�F=�qF=7F=��E=v�D=��C=��B=9�A=|
A=HO@={�?=�w?=�H?=T!?=w�>=�p>=��==��<=ص;=�w:=l29=��7=��6=6=`r5=W5=�5=5=K5=�{5=�5=��5=D5=�4=��3=�3=A02=�]1=!�0=^J0=h0=�/=a�/=��/=g/=��.=�1.=XQ-={Z,=�c+=�*=��)=�-)=j�(=�I(=��'= '=��%=Ն$=�"=�� =([=��=7l=��=�==s=]t=O�=<�=�0={	=��=��=Ǆ=O=�<���<\��<$��<���<��<���<���<��<2�<Z��<(��<d�<��<BU�<��<�<'e�<jY�<U��<�C�<���<��<Ϊ�<vܐ<���<��<��<0Et<o�h<��]<��S<��J<��B<&b;<�4<rG.<��'<9� <�n<c<��<�&�;��;Bj�;���;���;D��;g	�;�U�;�<h;�hG;�0#;��:Y:�:3x:���ՎH�����@����Vg:�V�V���t�!ڊ��1�������tǻ;Z޻�q��������%�r"�%])�[�.�{�3��<7�,{:��=�e�@�0�D�%8I��+N� \S��\X�ܹ\�@$`���b���c�"�d�]>e���e���f���h��Ek�z\n�\�q���t���w�V�y�[�z��{��{�,/{���{��`}���<���Nー3:��F����ˊ�㲌�9(���������B����H���莼엎�o���IՎ�2�������6���\�������"]������矚��7�������������u�����p���]���\���=���֧�����٩�0T������(��/����>��{���D���γ��y�����(���牽�������������Х��6z���i���  �  ��M=rMM=��L=r�K=��J=K�I=ׄH=N�G=� G=C�F=ѬF=3�F=U�F=�FF=��E=��D=w�C=��B=��A=ʛ@=��?=�)?=��>=��>=F�>=1o>=^>=8u=={�<=Mg;=:=��8=Fm7=�F6=^^5=q�4=+v4=�o4=p�4=l�4=�&5=bO5=B5=O�4=�T4=�~3=l�2=v�1=J�0=�!0=��/=ڱ/=��/=��/=�/=њ/=k/=�S.=3Q-=�/,=.+={*=�+)=w�(=�(=�'=<'=��&=t�%=�3$=l"=�K =��=�^=�=�C=d�=k�=1�=��=6Z=��
=@	=;X=�[=Y=s� =��<���<J9�<�B�<��<L��<)&�<���<E+�<�W�<p�<K�<��<���<x��<�A�<���<�>�< �<΃�<O0�<C؜<�3�<N�<HO�<���<�2�<�M~<�r<`:f<�[<��P<�G<x@<9<t�2<޳,</{&<ղ<�<n<l�<Α�;�;�8�;N�;A��;�ٝ;�F�;���;Qj;~�J;X';U��:���:�X:�4�%�`���º�E���&�KeC��^�wo{��{��`��;���u�ɻ�.�P���#��
�c���$%���+��L1�`{5�q�8�{�;���>�t
B��F�i�J�EP�E�U�*�Z�)A_��{b��td�TUe�te�/Ie��Xe��f�o�g��j�Wn�Rr��,v��uy���{��3}��}��m}��5}�.�}��~�/���Q�����o��+���(���Y ��S����u���ΐ�����;��1����7������m��6\��Jڑ�tœ��㕼�염ƞ���Қ�����Λ��ݛ��@������_���>���v���̤�����ߨ�BC���!�������Ϋ�O������᭼�����ڱ�J����W��U&������O߾�Pw���q��`�����������0������  �  !sM=JM=�aL=ElK=�IJ=ZI=�H=�AG=�F=�F=J{F=��F=X�F=�^F=��E=�E=)�C=�B=�qA=�H@=�[?=޸>=�`>=�@>=�7>=j>=��==�;==oX<=R/;=9�9=k8=S7=��5=��4=�L4=4=k	4=�C4=_�4=5�4=�5=}5=ڰ4=w	4=n$3=l2=I1=<G0=��/=�o/=+m/=�/=i�/=��/=y�/=�7/=*c.={I-=�
,=}�*=ȩ)=�(=�(=��'=�B'=��&=�A&=�P%=X�#=D1"=�
 =)�=�=�]=��=�e=A:=�L=�=��=xv
=�==�=��=�O =Z4�<���<�K�<\X�<���< �<ʬ�<�t�<y)�</��<�@�<2O�<��<s��< ��<S��<h@�<�j�<�A�<���<(l�<�/�<���<���<G�<3��<���<w}<�p<�d<2Y<E�N<}F<4G><?�7<�z1<g�+<�%<k�<�<@D< �<�_�;���;z��;�{�;���;���;�Ԏ;���;|�j;��L;X�);n� ;"�:�
:�?c��"s���κ����E-���I���d����s��
�����.`˻'��s���	����3����&���-���2��6�&�9�"�<�d?���B�9G���K��Q��>W��\�/	a��(d���e�ef��f�roe��e�;�e�rtg��wj�*rn���r�c2w�"�z��}�/�~��b�����~�J�~����]���x������@����?�����������r���_��쪑�Cp��J����3��n����}���ޏ�����wz��������� Ҙ����������/��E�������%��`Μ��-���+������[)��ۖ��8��� �����Js��}���ʬ�<N��Z����/G������^)ܺ������Ŀ�gc��eX¼>�¼��¼�"¼���Wo���  �  �_M=��L=aHL=�MK=&J=��H=*�G=�G=�F=(eF=�gF=~�F=��F=�eF=��E=E=}�C=Y�B=\A=b*@=S6?=�>=t7>=�>=�>=��==$�=='==;E<=E;=�9=�N8=m�6=��5=��4=#4=H�3=b�3=%4==�4=�4=�5=��4=�4=H�3=3==�1=��0=�0=O�/=�M/=gS/=K�/=��/=�/=��/=@/=Fg.=�E-=��+=g�*=&�)=��(=��'=�r'=�'=~�&=�$&=08%=�#="=��=A�=�=�7=�=�9=�=$=�p=*�= ]
=.�=�=�=ý=�1 =���<�\�</��<*�<Ԧ�<b��<
��<�]�<'�<���<T�<`�<��<\��<�~�<x��<��<�<u�<�[�<�#�<��<�r�<�k�<���<Ef�<���<O�|<�p<�c<h�X<�JN<�XE<8�=<�7<
1<D+<�8%<%y<�<)�<�<�D�;WK�;�U�;CC�;Zn�;m��;H�;&R�;k;zvM;�M*;Z/;�!�:��:Sjv�?z��Ӻ�J���/��(L�]�f�����5���������� ̻����U���"
�P�3=�o�'�L.��l3��J7��O:�q�<�)�?��)C�ZG�M_L��R���W��<]�D�a���d��jf�)�f�VMf��e��e���e�Rg�Bfj���n��s��w�|b{��~�!��������(�8#�/��i$���Ⴜ�(��nƇ�|������/���Ő�,���n���,�������b���я�:���������D����ǔ���$���Ӛ�G�n��6r��50��H��������������'�������M��iΧ��穼�o��~[��Nì�⬼~����������,��4n��y(���"������Խ�m��������¼@�¼��¼�X¼`��������  �  !sM=JM=�aL=ElK=�IJ=ZI=�H=�AG=�F=�F=J{F=��F=X�F=�^F=��E=�E=)�C=�B=�qA=�H@=�[?=޸>=�`>=�@>=�7>=j>=��==�;==oX<=R/;=9�9=k8=S7=��5=��4=�L4=4=j	4=�C4=_�4=5�4=�5=}5=ڰ4=w	4=n$3=l2=H1=<G0=��/=�o/=*m/=�/=g�/=��/=v�/=�7/='c.=wI-=
,=x�*=©)=��(=�(=��'=�B'=��&=�A&=Q%=q�#=m1"=�
 =��===?^=��=�f=�;=�N=.�=Y='y
=��=D= =J�=S =`;�<���<sR�<�^�<��<�<��<�w�<�+�<v��<'A�<sN�<C��<���<{��<Ա�<*;�<e�<7;�<ۤ�<Ge�<)�<ޠ�<D��<<ߏ<���<İ�<t}<Οp<Ʉd<�/Y<�N<vF<AK><C�7<p�1<�+<�%<��<<�Q<�<)|�;#��;ҳ�;^��;���;���;2�;Џ�;A�j;+�L;��);6� ;ĥ:K�	:cRe�f�s�WϺb�}-�gJ���d�V:������'���6��z˻�>�u�����	���W����&���-���2�,�6���9��<��?��B�G�O�K���Q�D?W�h�\�l	a�)d��e�.ef��f��oe��e�D�e�ytg��wj�.rn���r�e2w�#�z��}�0�~��b�����~�J�~����]���x������@����?�����������r���_��쪑�Cp��J����3��n����}���ޏ�����wz��������� Ҙ����������/��E�������%��`Μ��-���+������[)��ۖ��8��� �����Js��}���ʬ�<N��Z����/G������^)ܺ������Ŀ�gc��eX¼>�¼��¼�"¼���Wo���  �  ��M=rMM=��L=r�K=��J=K�I=ׄH=N�G=� G=C�F=ѬF=3�F=U�F=�FF=��E=��D=w�C=��B=��A=ʛ@=��?=�)?=��>=��>=F�>=1o>=^>=8u=={�<=Mg;=:=��8=Fm7=�F6=^^5=q�4=+v4=�o4=p�4=l�4=�&5=bO5=B5=N�4=�T4=�~3=k�2=u�1=I�0=�!0=�/=ر/=��/=��/=�/=̚/=e/=�S.=+Q-=�/,=$+=p*=�+)=l�(=�(=�'=<'=��&=��%=4$=�l"=4L =h�=�_=j�=�E=��=K�=��=�=�^=��
=�#	=U^=Zb=&==� =�
�<͘�<�E�<oN�<���<���<.�<��<�/�<oZ�<��<��<���<���<m�<69�<l�<n3�<��<�v�<
#�<�ʜ<�&�<��<�C�<7�<�)�<`>~<�r<2f< [<A�P<��G<B@<�"9<��2<-�,<G�&<A�<�'<��<�<<��;@<�;Tk�;{"�;���;���;�d�;��;�1j;K;yV';���:�`�:0�:�8�F�a���ú����&��C� \_�C�{�I���"����ĳ���ɻ�\�-��X6���)��0%�E�+��T1��5�G�8�D�;���>��B�mF���J�J P��U���Z��A_�|b�ud��Ue�Gte�MIe��Xe��f�|�g��j�Wn�Rr��,v��uy���{��3}��}��m}��5}�/�}��~�/���Q�����o��+���(���Y ��S����u���ΐ�����;��1����7������m��6\��Jڑ�tœ��㕼�염ƞ���Қ�����Λ��ݛ��@������_���>���v���̤�����ߨ�BC���!�������Ϋ�O������᭼�����ڱ�J����W��U&������O߾�Pw���q��`�����������0������  �  ��M=j�M=�	M=�8L=n;K=�+J=$)I=*NH=5�G=�5G=��F=r�F=�qF=7F=��E=v�D=��C=��B=9�A=|
A=HO@={�?=�w?=�H?=T!?=w�>=�p>=��==��<=ص;=�w:=l29=��7=��6=6=`r5=W5=�5=5=K5=�{5=�5=��5=D5=�4=��3=�3=@02=�]1=�0=\J0=f0=�/=]�/=��/=g/=��.=�1.=MQ-=oZ,=�c+=�*=u�)=�-)=\�(=�I(=��'='=��%=�$=y�"=R� =.\=]�=+n=�=c�=Kw=?y=�=��=78=
�	=L�=ͼ=5�=�(=+0�<��<J��<��<)�<@��<���<���<!�<��<��<��<R_�<���<LK�<��<��<+U�<H�<��<B1�<��<eߙ<%��<�ː<���<�م<�<94t<��h<n�]<%�S<�J<��B<zr;<T�4<Ia.<[�'<R!<��<�4<K<�s�;�`�;���;d�;���;*�;�3�;v�;%hh;G}G;o.#;Y~�:nڠ:�`:U���DJ�T��GY�����;��W��u��+�����{ϱ�X�ǻ\�޻{�����Ѩ��8�P�"��j)�?/�0�3�dC7���:��=���@���D�:I�q-N�<]S�|]X���\��$`���b�"�c�Z�d��>e���e���f���h��Ek��\n�e�q���t�Íw�Z�y�^�z��{��{�-/{���{��`}�	��<���Nー3:��F����ˊ�㲌�9(���������B����H���莼엎�o���IՎ�2�������6���\�������"]������矚��7�������������u�����p���]���\���=���֧�����٩�0T������(��/����>��{���D���γ��y�����(���牽�������������Х��6z���i���  �  3N=D�M=�gM=�L=��K=Y�J=?�I=��H=3H=��G=�G=ǭF=�AF=��E=�5E=0�D=��C=W�B={,B=�vA=y�@=s@=�'@=�?=ʰ?=�T?=��>=�	>=�== <=��:=�9=Z�8=2�7=�6=5B6=��5=4�5=ӱ5=)�5=��5=��5=-�5=�5=�#5=�4=%�3=/�2=�2=�W1=9�0=)^0=0=��/=bu/=U/=̑.=��-=�:-=4v,=M�+=1�*=�b*=��)=~k)=�(=RQ(=rv'=5O&=g�$=�#=e!=��=��=�-=�=˄=�W=�L=_=F�=T�=F�	=P=7=�=��=�f�<�E�<0�<��<�?�<��<c\�<��<6��<�t�<���<���<2��<��<ъ�<���<�ױ<H��<b��<g�<,L�<W��<���<�"�<�G�<��<���<r��</�v<��k<�a<�%W<�N<��E<$><y�6<� 0<U)<�Z"<o�<��</
<�� <}��;�[�;�d�;�W�;�,�;���;�(�;[�d;��A;��;��:;��:H�:�ȳ��_4��G�����#����1�m�O��Go�WՈ�l�����=�Ż)�ۻ��a����<��X�f&�vR,��K1�[�5��/9�3�<���?���C�Q�G�Q-L�~�P�ѯU��Z�c�]�j�`�J�b�XDd��e���f�hHh��j��Il���n�jGq�a�s�q�u��w�z�w�-Xx��x�By�0z�6|���~�M4���6���V���s��Jn���)��z����|��H���9��V4�������������I�������[���4h��YF���������ݽ�����$����F��X ��!'���f��ڠ�<n�����e���ɦ��ŧ��y������[~���.���5����������m������񁵼d᷼��:���+v�������*������ܦ��C���"ӿ��  �  �SN=�N=��M=LM=�EL=VbK=�nJ=_I=��H=��G='*G=@�F=��E=BQE=�D=ND=$xC=��B=�GB=��A=XA=tA=�@=�w@=M@=C�?=�>=b+>=�:==`9<=u3;=�3:=B9=g8=��7=o7=��6=�h6=�=6=�$6=�6=�6=��5=ܼ5=�d5=��4=�64=Jp3=�2=��1=W+1=f�0=�	0=��/=>/=Ԗ.=.=H�-=��,=�o,=Q�+=�_+=�*=�x*=�*=�x)=#�(=�'=�&=D%=qF#=�[!=2N=[&=��=ʫ=o=�@=W%=�=-=$=�3
=8C=�H=�7=�=�]�<�p�<*^�<cG�<�G�<Xj�<���<x��<�M�<���<i��<	��<I�<�E�<c��<��<��<�y�<��<�<\%�<23�<���<3`�<K}�<-b�<V$�<�ց<�y<�n<�gd<[�Z<��Q<��H<��@<^9<��1<�P*<b#<Թ<i�<I�<��<���;^2�;G��;�ϸ;f4�;��;���;y�^;�z9;�;o��:�y�:N:�誸ѡ&�3P���rٺ��=m*��I��fk�g������a��GHĻ�Uٻ+�W8�,�
����7��S#���)�w0/��4� @8��<���?��C�
�F�0�J�/O��rS�3�W���[��_���a��Sd��of��_h��<j�Ul�_�m��o��kq���r��1t�Gu�U�u��v���v��w�1y��m{��c~��瀼����T���~d����5���Pފ�oՋ���������6��c������6�������������*ɐ�H[��d���䕼@���D��Fq��׫���՜�����'���W������Ƣ���+���󥼣���"O���ߧ������{������-\��FC���X��t���c����������8[���Ȼ�T弼Y����P���þ�N��qu���  �  �;N=��M={�M=�M=�|L=�K=�J=`�I=��H=��G=�
G=B4F=�kE=ٲD=�D=~C= C=��B=94B=�A=��A=�\A=A=��@=�N@=z�?=��>=I>=�%==v<<=�\;=�:=��9=�9=�m8=��7=�e7=��6=�6=Ib6=�(6=>�5=��5=_�5=�e5=y5=�w4=9�3=>�2=?,2=�[1=��0=��/=s*/=�.=��-=q-=+�,=T�,=�;,=��+=M�+=:+=��*=e*=��)=��(=��'=�~&=��$=�F#=U{!=��=~�=��=4u=J=�=s�=}�=�=Si=�P
=(E=�A=g;=m"=���<�#�<-2�<��<���<���<ę�<�}�<(j�<]d�<lu�<���<� �<a}�<��<�<d�<��<	@�<t�<i��<LP�<&ؚ<P!�<�@�<*O�<[�<�j�<]�z<	3q<g<a�]<8�T<ͯK<�B<�|:<W2<��*<W�"<i�<�<{"<%�<2Y�;[O�;��;#��;;'��;Ԡ};��U;٢.;;a��:Эw:�9�F��^%��ʒ�Ѻ�V���&�{ H�a�k������S���o����Ļ9Yػ\�뻌����X�������� ��a'���-��"3�	8�gM<��	@��oC�_�F�uEJ�aN�6R�_RV�irZ��T^�8�a��e�� h���j�&�l��n�<'p��Vq�*Gr���r��s�<�s�D0t�8�t���u���v��y�L�{�k�~����h����%�����������1��OS���N��%���݋�\}��B��y��G܍��>������Ao���q��lǑ�!d���-�����Ә�c���0��8����(��u��+��������w���=���뤼�����	��F���&8�����iI��@ʪ���� v��yf��hJ�����J̵�yf���⸼�:���h���p���Z���)��'߾�}���  �  ��M=ΓM=�FM=��L=�hL=��K='�J=�I=��H='�G=L�F=��E=y�D=��C=�FC=�B=�cB= B=�A=��A=n�A=�vA=�1A=y�@=�3@=�u?=��>=�==��<=�<=R;=��:=":=�9=D9=g�8=��7=�o7=+�6=�m6==6=d�5=�w5=�K5=i5=��4=�n4=;�3=3=?2=]S1=+d0=�z/=L�.=�-=�0-=Y�,=N,=,=��+=��+=��+=O+=��*=�~*=��)=��(=�'=�0&=h�$=�	#=�b!=��=��=z=�==��=��=+2=��=\z=q4
=�=��=i�=�="��<)C�<�y�<c�<_�<���<%$�<��<p8�<���<i��<m�<
��<�a�<�\�<���<�Ʋ<U�<�Z�<&s�<VJ�<�ٞ<*+�<1Y�<���<�Ƌ<&�<4��<�<|<�5s<oj<��`<o]W<��M<�tD<�2;<lE2<��)<��!<pS<j�<~<g�<X��;LG�;jr�;��;F��;��;D3u;�J;��!;��:��:0�J:u͍9��]�R�1�㜔��к�)���'���J�jVp�Z���"����l���ƻ��ػ��껎���{Z��������M�Z�%�H�,��3�Э8�~�=��A���D��G�\�J�@N���Q���U��0Z��~^���b���f�4j��Um���o�b�q�;�r�Йs���s�%�s�J�s�n�s���s�[t�M�u�Սw��$z�6&}��"��ם����������#����������
��w������!��b���ݍ�(�����mh��q폼2����ő�q7��b�������t��F��l잼������f��<飼�|���礼:�����]ݥ��\������9��۫��Of��H��)���갼����과7���s�������븼.��Cu��B�����S
�������  �  9WM=?�L=�L=muL=�L=
�K=��J=K�I=��H=>~G=sGF=#E=1D=#C=pB=��A=�A=ʍA=��A=v�A=#yA=�VA=NA=��@=��?=��>=
>=�==�I<=n�;=�;=��:='Q:=��9=�9=�9=�f8=��7=�6=0I6=t�5=�65=@�4=Q�4=?�4=`o4=J%4=��3=��2=02=�1=�
0=G�.=p�-=�-=�],=a�+=��+=�b+=�V+=�U+=N+=�-+=��*=iX*=�)=sq(=# '=�%=7 $=��"=!=�=�	=cd=Q�=��=�d=�=A|=��=vY=y�	=�=du=Uw=�=#�<���<�@�<�8�<!��<b+�<�_�<K��<}��<S�<,(�<�e�<��<��<+U�<kƵ<H�<���<���<���<���< �<x�<�"�<�`�<�ي<���<^q�<��|<[�t<^�k<�b<�eY<�lO<�@E<(;<l1<�I(<��<�3<\�<P�	<3]<ga�;`M�;e{�;8�;���;�<�;Q�j;�p>;��;(�:)�:��:��8 )���|H�a����׺a�
�c�,���Q���x�O�������-���* ʻۻ�)�ܩ���������������$��r,�ө3��:��?�_�C�xPG�J���L��qO��R��xV�x�Z��g_�d�v�h���l��hp�E6s�;u�6v�"Dv���u��Qu���t�R6t�Ct�,u�7�v��%y�`/|�Pu��H��3���o����n����˛��]=��t
������N�����L"���|��ץ��l���K$��󊐼j琼�l��E��(����7��@��f����ڛ�~)��[O���/������;����e��۹��إ��ݥ��ꥼ� ��j���s���|ڨ�?���z��s���E��-Ա�����������յ��ȶ�n근�C���ͺ�s�����䖿������  �  ^�L=NL=L=��K=��K=s*K=�zJ=��I=4dH=>G=4�E=y{D=VPC=�WB=�A=S-A=K�@=��@=�	A=f%A=L0A=A=ھ@=�)@=!Z?==b>=^==m<=��;=�;=;�:=\�:=\:=|+:=��9=o]9=��8=��7=��6=�6=;5=a�4=U:4=�4=A�3=��3=�3=�U3=��2=S�1=��0=E�/=�n.=�O-=�T,=�+=Y+=��*=�*=[�*=<�*=-�*=��*=ڡ*=&*=#)=��'=��&=�%=�}#=O
"=�� =�Y=�=��=��='=W�=�N=��=`�=�=�t	=9=��=j�=1� =�/�<�*�<���<Y��<zR�<���<Qy�<�d�<o�<$��<��< ��<h��<\��<48�<��<z��<��<=Z�<�-�<:��<k��<S��<���<[	�<���<x��<k�<.�|<�Ku<�Lm<�d<��Z<�VP<XuE<��:<Q0<FK&<^z<�<�<ݭ<@� <ק�;� �;�o�;�ζ;cȟ;S�;v`;$$2;�_;�d�:�Kh:iY�9�%\��=���;d�%狀�~�:����3�tcZ�g����\�������V��كλn#޻=��2}��T7�7���R����>$���,���4���;���A��F�J��L��N��4Q�*T�y�W�!�[���`��e��j�
~o�	rs��qv�TVx�/ y���x��/x�Fw�>�u��Ju�!Uu��Wv�Y_x�E{�$�~����!����Ѓ�j���a���9��%f������I[��/g���؈�U���g��'��Y���Eɐ������呼����o������$�����8ϗ��6��Ȝ�wV��e�������N��LX��o়����ᦼ���B��������0��?;���é�%���#ȭ�Jӯ�l������t과s����������t1���7��/����q��:s��U}��p`��=����  �  �L=ҩK=stK=�TK=�&K=~�J=E+J=[BI=�H=ھF=XSE=��C=2�B=f�A=��@=7�@=#^@=Sn@=-�@=1�@=��@==�@=�l@=�?=��>=�==ƽ<=��;=V;=��:==\:=�N:=�Q:=TF:=::=�9=�8=/�7=��6=Ͷ5=��4=	4= �3=�d3=�\3=7_3=�H3=~�2=�i2=$�1=x0=&;/=,�-=�,=��+=��*=�\*=�!*=�#*=NM*=H�*=�*=��*=Z*=��)=��(=�s'=7�%=Mg$=��"=�!=r= =�=��=��=�=�C=P=_z=��=(�=��=�	={=A==�A=�o =�E�<�l�<��<=�<���<���<O��<a�<U<�<�k�<��<�]�<97�<鎺<�>�<*�<C�<g��<���<�d�<Ŧ�<d��<�m�<Zk�<�ǌ<���<��<O�<�m|<W�u<�n<A{e<��[<��P<OE<@�9<��.<?N$<�(<^1<�)<��<���;���;���;<4�;Ub�;�Ϝ; M�;?iW;�';Z�:��:�::T�t9��I�D_���}�;㲺�&�?f���:�[�b�|l��3����ٯ�/X»K�һ�H�li�u�������
����H��($�S-��6�r�=�;D��-I�e�L��O��Q���R��tU���X�O]���a��bg���l���q��v��.y��{�"�{�aM{��&z�I�x��Fw��mv�t�v���w�z��P}�����A^���烼z���񆅼7��������_��\o��v����@��������Ȍ�2ގ�-��������ɒ�$(��!F���k���ݓ��̔��P���b��O㚼n���U\��u碼������ʲ��x"��@���̧�Pg���"���6���̧����������¬�j ��y��vղ����ô�����7���c��[ص�ɶ��I���J��q�������1��uü�  �  ��K=�6K=K=��J=w�J=��J=��I=I=��G=$F=nE=Z�C=FB=�7A=�y@=�@=��?=B@=�Q@=�@=��@=`�@=�/@=4|?=�>=k==�M<=�U;=x�:=6:=>:=>":=(C:=�P:=�':=��9=��8=��7=�6=z5=�o4=b�3='3=3�2=u�2=� 3=��2=��2=�12=8Z1=�>0=@�.=@�-=�[,=�B+=m*=��)=��)=��)=l�)=�?*=ss*=_s*=:%*=�y)=aq(=�'=g�%=��#=fv"=�!=j�=�=?�=R�=(3=�g=�.=R�=W�=�=N�=ի=?=��=��=� =���<���<���<��<�b�<�h�<��<��<�m�<q��<�)�<�o�<�W�<ɹ</��<?��<;s�<��<4�<�Ԥ<��<Ϛ<᎕<���<��<9Ӈ<�D�<��<)|<̷u<�n<Af<\<��P<�E<39<s-<��"<�~<�v<:�
<z<8�;��;���;+��;���;��;�ā;PQ;~� ;���:�p�:�m:)�9�畹�.��q��������󺀜���?�@�h���K@�������Ż��ջ
�㻘�ﻨp�����d
�s�:��!7$�C�-��6��(?���E���J�l�N�g�P��R��6T��~V���Y�[�]��b�\uh��n��Ss�F�w�{���|�Vx}���|��z{��y�/x�iBw�E^w�>�x��E{���~�E[��B���̄��̅� 9��(��I̅�_j���M��M���qʆ������������Bj��Ra��:Ӓ�����	�������Wr��aH��8���Θ�g[��30����T���������X���7���zڨ�l���駼/������ @��g��:P������,ۯ���������״��f�������h��i]������
���C��%?���ļ�ob�������ü�  �  ��M=PfM=TM=d�L=�JL=G�K=�J=�J=�H=��G=)1F=1�D=s�C=^�B=��A=��A=%VA=&SA=�kA=�A=��A={A=�.A=��@=��?=�?=�;>=Ui==Ͻ<=4E<="�;=��;=x�;=;�;=9;='�:=�:="9=/)8=�.7=K6=1�5=*5=y�4=4z4=�>4=I�3=�k3=[�2= �1=��0=�w/=O:.=�-=�,=�0+=ğ*=�O*=�5*=�=*=-R*=�Y*=�=*= �)=�Q)=�q(=�P'=��%=d�$=�&#=��!=�� =�H=f	=_�=T=�E=�%=�=�!=�f=O�=
=��=TV=�D=�I=���<�]�<��<���<�G�<	x�<.s�<�c�<�x�<1��<���<��<���<]J�<�<.��<�~�<b�<�i�<�]�<���<eM�<}��<˔<�L�<L'�<\[�<̈́<�P�<�g{<��s<��j<ka<�W<FL<-NA<b�6<�,<�k#<� <^t<��<�T<�#�;���;���;m�;F��;_6�;��j;��<;z�;���:��:� :�OA9��_�2��r􂺎Ϻ����l���1B���h�����#����(���/��&�ʻfػ����$�5 ��������'� � ��(�]D0�ס6���;���?�KC�VF�*I�\lL�YiP�9U�?$Z���_���d�O�i�{�m��2q��Is�J<t�9t�#�s�ۄr�Ԋq���p�|q���q�G�s��Lv�\Fy�uN|��~�@����!���l��݉��L��������������:2������s�)܊�Վ��a獼Rݎ�_����������샑�Œ�{x��Ӗ��J��ݠ��:������$���]J��>U��Zۥ�`���ҥ�f����o��������3�kK��L���ɫ�w������F��v��؊��P汼�R������&��au��bF��YY��:���0����T���  �   N= �M=#M=\�L=�aL=��K=�K=LJ=[�H=��G=PHF=��D=��C=q�B=�B=��A=�sA=$mA=,�A=��A=��A=��A=lAA=��@=�@=8?=�W>=��==g�<=YX<=�<=V�;=$�;=b�;=�,;=b�:=i�9=9=�)8=�67=�Z6=��5=�'5=c�4=~�4=�W4=4=H3=O�2=��1=��0=��/=�R.=h(-=�",=_R+=N�*=so*=�Q*=VV*=2g*=�l*=O*=l�)=�d)=ֆ(=�h'=�&=�$=
@#=0�!=�� =�O=�=��=�=�6=X=��=�=]f=��=
=3�=n=S]=1a=���<���<���<6��<Rg�<s��<���<]��<��<��<9��<>U�<�5�<���<!�<��<Z��<�A�<E��<��<y*�<���<
��<h�<˃�<�T�<�y�<�ڄ<xN�<ZI{<8fs<��j<+6a<��V<�5L<"ZA<��6<��,<��#<Q�<-�</]<ȧ<��;s�;�Z�;���;Õ�;l�;ܥl;g�>;��;�M�:��:ȏ(:e*^9MPF����D���*��'N��c6��~@��f���������O��ă��@;ʻ��׻E��_�; �8�����<�N� �N�(�0��E6��^;��f?�P�B�L�E�حH�|L�` P�R�T� �Y�'._��qd�Pi��xm�h�p���r�A�s���s��%s�\/r��>q���p���p���q��ls���u���x���{�7�~�!T��( ��[��Y������K������σ��D������눼�Ɗ�*j��&���򦎼�M��0׏��v��OY�����U���r��iߘ��t�����fi��ts��������
���¥����xl���J���g��7⥼�ʦ�����©�ݑ���X��o箼1��� ~���豼a��8����������U��]��0w���t��5+���  �  �DN=��M=�nM=FM=a�L=�	L=~@K=�CJ=3I=��G=A�F=yHE=$&D=�3C=�|B=�B=�A==�A=��A=	�A=��A=y�A=�tA=B�@=N@=`�?=أ>=v�==c==��<=.'<=��;=�;=�e;=�;=s�:=��9=T9=�(8=fK7=�6=��5=:o5=�5=�4=x�4=R>4=*�3=��2=�
2=&�0=5�/=��.=Bx-=�{,=��+=�+=��*=0�*=�*=�*=��*=�~*=�**=ݗ)=x�(=��'=k`&=��$=��#=="=� =�a==��=a�=	=^�=΍=�=zd=��=�?
=2�=�=��=b�=07�<���<KE�<�5�<���<0�<`�<a$�<�W�<���<O��<7�<p��<�&�<���<�b�<�<x��<��<��<��<^�<d^�<c��<��<�Ȍ<lƈ<0��<\A�<�z<��r<Qj<ߕ`<|V<9 L<�wA<}=7<[�-<��$<e�<��<e<6�<dY�;��;���;o'�;�]�;��;
�q;�D;�;���:�2�:R?:���93����r�������)�@�;��a����������%̹�(ɻy|׻5L�l)��� ��]�?U����� ��[(��T/��P5�E;:��0>�|�A��D���G�bAK�wWO��S��Y��=^��Zc�uh�l��1o�!Gq�Ur�1�r��r�a<q��ip���o���o���p�c|r���t���w�$�z��q}�
��|����,������ׁ��N��V
��7��g��"���߈�����	���5�����Ĵ��WE����}䐼�6��L󓼍��Tr��f���u��������`H��SW��Q祿�&���������#䤼_���}��+\�������6���������3\��K���Φ���^����x����X��`l��Ե������l���\���-�������  �  ��N=y4N=q�M=IsM=�L=�UL= �K=نJ=�cI=*H=��F=��E=��D=�C=C=W�B=vFB=�%B=�B=\#B=�B=< B=غA=�GA=,�@=T�?=?=5>=6q==��<=�L<=��;=�;=3;=��:=�?:=8�9=e�8=28=vb7=m�6=�46=^�5=��5=�E5=/�4=2�4="�3=<3=1N2=S?1=�0=��.=��-=� -=A=,=��+=�N+=�+=�+=��*=�*=��*=Lk*=��)=`)=�(=��&=FZ%=��#=�c"=�� =t=E�=�_=��=>�=n�=�M=�=Z=�=t
=�-=�
=� =}�=���<�y�<`��<��<B�<���<?��<c��<�P�< ��<5��<q4�<:��<7�<���<��<��<MB�<���<���<�h�<��<�6�<A{�<֑<jb�<L'�<��</�<'+z<;�q<Q�h<�_<M�U<�K<ׄA<��7<��.<u&<�<Oq<��<0�<E��;���;���;B\�;]��;F%�;R�x;;�L;,#;R��:���:'ya:�s�9Q�������]��W����]����5���Z������0��Y���&�ǻ�.׻������t���`	� 4�y��� �]�'�s.�P4���8��<�Z�?�;C��dF��J�YEN���R�.�W���\�&�a��-f���i��l�/o��9p���p�gp���o��;o�L�n�)�n�޲o�R5q�,hs�Zv��y���{�=h~�s4��J�������*��꿂�Đ�������腼b\��݈��J������Z���TI���㍼�}���=���E��é���m��9���W֗�g?������ɞ�5���,��"?���飼b>��BV��YQ���S��?�������.ƥ������v���,��[�����D��;G���>����沼�ӳ�����}Q��:㷼����9D��ռ�?-���  �  ��N=ݜN=R?N=W�M=�LM=�L=��K==�J=@�I=ӃH=:[G=#AF=�AE=VfD=j�C=t4C=��B=B�B=7�B=�xB=�eB=�@B=��A=��A=��@=�F@=�u?=�>=��==�==5i<=��;=_;=�:=�g:=��9=�E9=̤8=?8=n7=��6=�6=|26=Y�5=�5=ZW5=��4=�C4=n|3=9�2=T�1=X0=�u/=�|.=��-=b�,=5V,=�+=�+=�{+=�Z+=�7+=�+=,�*=u*=�X)=�W(=0 '=��%=�;$=_�"=�!=y=��=�=*D=�K=G.=��=��=
==��=�
=v=Pc=�]=�U=�: =��<�7�<;�<���<r2�<��<O��<�x�<�2�<�5�<��<=�<�9�<w�<�<,`�<+ذ<�,�<sH�<��<���<<�<�V�<V��<���<|y�<g�<`р<�y<�Fp<�?g<��]<�aT<^�J<9SA<W08<˃/<�V'<��<��<�0<�<5��;���;��;s��;Ь;R��;�؀;zW;�2.;$�;���:�+�:�:|S�8����
LH��x��8�ٺ�x�/��T���y�},����lT��D�ƻTO׻�H�^����(��
�Ł����"!��'���-���2�k7���:��<>���A�HE���H�=M�z�Q�ҙV�IX[���_���c��{g��Qj��cl�w�m�_[n��~n�oLn�3�m���m��m�՞n���o�`�q�K�t�5dw�iYz��#}�H��o׀����T����h��T���^��쇆�����z���������ۋ��}��6��㴍����<���#���쒼:���
/��Oo��˝������{c���ՠ��˱���,��
r��4���[���u���[s��T6���N�����\��o ��s⬼��������8��nZ��kn�����������	���q��⹼�F������H����  �  EO=!�N=�N=�N=8�M=G�L=��K=-�J=>�I='�H=m�G=�F=%�E=RE=�lD=��C=NxC=)C=��B=��B=�B=\kB='B=��A=A=A=��@=g�?=��>=�>=e5==�n<=�;=;=|:=~�9=i\9=�8=UK8=q�7=�a7=�7=��6=�~6=�C6=$�5=��5=�5=Qp4=N�3=4�2=��1=0�0=�/=�/=F.=��-=�	-=Q�,=;,=+�+=ܳ+=�v+=�.+=0�*=ID*=r�)=�(=�f'="&=y$=��"=�&!=zd=�=Y�=��=��=N�=r=�;=�=
�=��
=ܦ=,�=��=��=Gn =N�<vx�<Za�<-�<<��<fK�<\��<2��<F��<K��<���<L��<`�<f�<���<r�<DF�<���<��<i��<Q�<<X�<�3�<�`�<���<��<�O�<�rw<�Hn<�e<k�[<��R<a�I<	�@<�48<"0<�C(<Ū <<�.<��<���;��;��;&n�;�[�;�9�;�L�;|�a;��9;��;�G�:=��:�2:��X9�5����6�!"����Һ	�P�*��N��t�|S��絠�>̳�TSƻ�1ػ^j黨���C���D��U���!���'��1-��1���5��~9���<��x@�|5D�??H�ؑL��Q���U�0�Y�G^�p�a���d��g�t�i��k��l��l���l���l�2m��Gm�_�m�^!o��p��Is��v��"y��5|�!�瀼����=��#M��'U��<\���a���]��&H����9Ȋ��Z���݋�:j��s�����hF��	ΐ�Ԙ��!���נ����������n��"
��	j��D���#l�����$�������GG������-!���٤�'ۥ��(��?����z��2P�����*ү�bc��_ղ�0/���y������k���.9��{e��Kz��)p��C���  �  �gO=�O=ƹN=7;N=?�M=�L=��K=9�J=T J=0	I=H=�BG=�xF=L�E=GE=��D=<	D=Y�C=�>C=��B=�B=qB=P)B=}�A=IQA=�@=��?=C?=�+>=<==�S<=�x;=`�:=��9=�Q9="�8=eA8=��7=}7=
67=d�6=!�6=�6=:o6="6=z�5=I%5=�s4=��3=��2=��1=�1=�L0=��/=��.=AF.=8�-=�5-=��,=W,=��+=�+=s9+=��*=�A*=��)=)�(=R�'=,)&=��$=!�"=0!=&/=8=�3=^%==�=�=(�=T�=a�=E�
=�=2�=��=E�=�v =jH�<rg�<_X�<q/�<0�<���<B��<���<���<��<�^�<���<�k�<{0�<� �<Z9�<�n�<3��<kթ<{ե<���<O�<�g�<܂�<;��<��<@��<K%<�ju<��k<�~b<�ZY<�yP<��G<7�?<��7<i0<�(<I*!<��<ԃ<�	<s��;���;O�;�A�;5!�;��;]S�;��k;YGE;�;�	�: ��:ĒS:�_�9�"E��-�WD���Lкϟ���(���K��p� ����r��?R���ƻ
ڻp컺	���[��.�_s����"#��(�[@-��o1��45���8�QP<�B@���C��(H��L��P��U���X�|s\���_�%`b�+�d���f���h���i���j�u�k��[l�N�l��:m���m�c�n���p�޵r��hu�Ղx�m�{�d/�6������!���g������
���&r��3��cӉ�?V��q���E!��������d׌�����s4���ɐ�~����l��I�����FÙ��R��.������3��D9��o��ޡ������������q���Ϥ�����7j���#�� �������ﯼ̱�Ɗ���'��i���9����)��(8��#���뻼̕��)���  �  (`O=�O=��N=q)N=zM=ΪL=`�K=��J=��I= I=�XH=r�G=��F=�WF=	�E=VE=�D=��C="qC=��B=��B==LB=��A=�A=5A=�@=,�?=C?=O!>=�==0<=";=l/:=�[9=ϥ8=�8=e�7=nI7=D7=��6=�6=r�6=:�6=�l6={6=�5=5=oH4=!~3=Ѱ2=��1=�81=�0=t�/=�l/=��.=iQ.=��-=R/-=�,=�,=��+=_+=֞*=*=�b)=	�(=p'=�&=��$=��"=!� =��=D�=5�=As=�O=�5=>)=+=�:=U=ev
=�=t�=)�=*�=pO =?��<f��<N��<x��<	�<j/�<k�<��<�<�O�<>��<i��<qF�<���<�f�<�=�<�C�<�i�<���<ʥ�<���<j�<Bn�<}�<�Z�<m�<.ڃ<�D}<*
s<Ci<5�_<ҋV<H�M<�E<X><c�6<G{/<�N(<� <gE<�<9j<܄�;?��;6�;1��;߱;t�;蔌;Lt;�jO;�[*;�';(�:�!n:�|�9�&�b�,�^���s�Ӻ�$	�&�)�|�K��Fp�Df���y������Ȼ.�ܻ�8��Z���	�������>�>�$���)�"�-���1�S75�t�8�4j<�8S@�
{D��H��M�$@Q��U�waX�_P[�h�]��6`�7[b��dd��Wf��*h���i�#5k�Tl�.m�Y�m��n���o���p���r��ru���x��|������ ���4������(ꇼBꈼ�����7������JԊ�����8��������I�]������l!���ے�唔��6�����G��7d������
Ҝ����+1���R���_���O��T��Wϣ�s���#�����z���x��$'�����3+���Q���o��s���L�����V��7|���b��������_����Z���  �  �4O=u�N=��N=l�M=�0M=�XL=dtK=D�J=��I=RI=�tH=A�G=%_G=��F=�:F=��E=��D=N/D=�C=��B=KjB=>B=��A=cTA=��@=k@=K�?=:�>=��==��<=��;=�:=��9=�8=$�7=6[7=��6=��6=2�6=��6=K�6=��6=�w6=B6=��5=w^5=&�4=1�3=�.3=Rq2=2�1=d91=M�0=�K0=;�/=#^/=|�.=0.=��-=.�,=�,=u+=�*=QL*=��)=9)='=(=b3'=��%=5[$=W�"=ƒ =�p=�8=��=�=�=8r=�r=��=�=��=�(
=�Y=fu=�q=!J=��<�/�<dB�<S�<�|�<���<HE�<U��<Dj�<���<yY�<H��<���<^��<��<�j�<���<�ΰ<�٬<�<� �<0�<�Ɯ<V#�<&-�< �</��<	�<.({<��p<]Gf<ؠ\<�S<�NK<-�C<�D<<uJ5<n.<lu'<Z) <�a<�
<�,<@��;��;Y��;
��;J��;�&�;�;�1{;��W;�D3;�;��:Չ�:4l�9�)���5�����S6ܺ�L�*+-���N��zr�>b��)��������ʻI�r�������&��*����!���&��+���.�Dd2�o�5��\9��,=��JA���E�J�!TN�7R�&�U�"XX�1�Z�K�\��{^�R\`�wbb���d���f�[i��k�F�l�� n�'o���o���p���q�7�s�� v��5y���|�Fl���|������^������*T��mQ�������V���|������N����������v���a��F���!���Ǒ��r��\���f�����O�����������Bϛ�
��Y`��������^��vs���W������ȥ����������ڨ��z��j��{����簼�<���y��a����N��Oú��ܻ�g���m��@j��;����ʽ��  �  w�N=��N=�9N=ŗM=T�L=��K=VK=�8J=��I=��H=WxH=dH=�G=�/G=h�F=~�E=-%E=oPD=�~C=Q�B=, B=��A=tAA=[�@=r�@=<@=�x?=H�>=��==�<=Kg;=�7:=�9=�8=gJ7=!�6=YN6=�6=�6=�$6=�;6=-G6= 76=[�5=r�5=�5='P4=#�3=
�2=&2=W�1=�"1=K�0=�0=�*0=�/=�0/=K�.=�-=�,=�,=�<+=��*=z�)=sJ)=T�(=�'=��&=f�%= $=GB"=v7 =,=r�=.Z=e=��=/�=��=q�=�3=ށ=x�	=�
=�(=v =`�= /�<�O�<�_�<��<���<Jh�<l,�<Y�<���<E��<|$�<�c�<�i�<N�<s3�<�=�<��<�+�<��<_<�<h�<?s�<:�<���<䯒<>c�<�ׇ<�-�<�y<�n<h�c<��Y<M�P<��H<TA<te:<�3<x$-<M&<P<�<:�<�<8j�;y��;��;�l�;=��;Zf�;*g�;�;�5^;� :;��;u��:dr�:X�9i<E���D�F?�����^��o2�P<S��bv�5*��'z���ҷ�g�ͻa��x����;�mF��?�����#��(�
�,�o 0��m3�{�6��`:��W>�	�B�0G���K�Q�O���S�rV�z�X��aZ�>�[��5]���^���`�[Dc���e��h��ek���m�jo���p�l�q��Rr��^s���t��2w��7z�y�}����UE���v�����MC������k���$6��fo���h���@�������b�����M��\���򚒼�5��q����Ö����Jr��//��4��p
���M��ɝ��h��:����������
��7䥼�����W���>���p��d����물�&��5����� ��ڴ�� ��� ���*���ӽ��)���F���K���\���  �  ��N=�hN=Z�M=�@M=�mL=��K=��J=��I=<I=��H=�mH=�%H=��G=(oG=j�F=,*F=%OE=�^D=ImC=ݎB=��A=�CA=��@=|�@=0@=q�?=j.?=]g>=�n==$M<=�;=^�9=�8=��7=��6="6=�5=��5=��5=��5=7�5=L6= �5=i�5=rG5=��4=��3=�"3=�d2=A�1=�P1=r1=n�0=c�0=�_0=��/=(s/=�.=�-=��,=��+=��*=�0*=�~)=��(=};(=m{'=��&=�N%=z�#=��!=V�=�=T>=M�=Yz=;=�#=�7=bp=E�=�!={	=��=��=��==�=�d�<�v�<���<���<�1�<���<���<k �<�7�<�<߰�<���<���<��<B1�<=��<��<σ�<�Y�<}v�<N��<,ʟ<��<0�<(-�<�׌<x6�<�l�<uFw<l<]a<��W<ͣN<��F<�r?<��8<_2<)�+<�'%<��<��<�,<�<��;�O�;�;�;q>�;X�;1�;�8�;�ȁ;��b;��>;�I;�y�:!��:q��9{�k��OU�ױ��������7�-X�Ԣz�b���j�������7л��滶.��>��m�Rn��) �ճ%�%:*�S�-��K1�vw4���7��s;�ߏ?��D�h�H��LM�9oQ�t�T�BgW�+Y�a]Z�oP[�O]\�)�]���_��db��pe�p�h��k���n��p��1r��&s�i�s���t�>3v�`Qx�}C{���~����$����J���t���Q��Iŋ�t����?��]���4���쌼��������錼Ǖ��g������T����j������;��-���ؗ�9\������􍙼ق���̛�xf��8�����|ꢼ�|��x�������k������屮��q���<q��E���95��vѴ�&^��%���k����6��z@��վ�y�������꾼�  �  �N=�5N=�M=� M=�&L=<K=TZJ=�I=^I=ˢH=�aH=q.H=��G=F�G=�G=�LF=�eE=icD=G\C=hB=��A=��@=܍@=>:@=D�?=J�?=p�>=^5>=�===�<=|�:=��9=�U8=�?7=	`6=��5=k5=�O5=ja5=��5=
�5=��5=+�5=��5=�5=g4=��3=5�2=�2=O�1=W!1=l�0=��0=@�0=n}0=F%0=/�/=��.=j�-=��,=1�+=��*=��)=�3)=N�(=D�'=F5'=�H&=%=1�#=��!=٨=�\=��=�~=�= �=l�=��=�=�x=��
=UA	=Ӈ=�=��=�Q=���<7��<|��</%�<���<���<���<*$�<}a�<�`�<�<x9�<v�<%��<�$�<�¸<Z��< �<%ʪ<��<&!�<�L�<�5�<���<�̑<�r�<�ņ<]�<�v<&�j<��_<��U<� M<�AE<�2><��7<�l1<
+<�V$<��<��<$<w�<���;z��;L �;���;?V�;��;���;ж�;)1e;R�A;��;Q�:���:��9_����b��ݹ��W���T���;���[���}�����ۥ��~����ѻ���p�����	�����s�!�~�&�=U+���.�r2��75�Ά8�@<�=v@��E�N�I��zN�V�R�J�U�-#X���Y��nZ��[���[�-5]�84_���a�,e�W�h��8l�Ko�I�q��Us�Xt�eu���u��!w�L%y��|������ur���؆�(��4������{�������l���Uc����n��`L��S���%�������Q��+��Ԅ��:���)�������W��R���+K���4�����/0��"���/���)��B䤼�C��F��M������Iq���~��񫼯ҭ��������R����]��g�����Z����G��������_���O���  �  TnN=r#N=L�M=5�L=kL=E K=�>J=�I=�H=�H=�\H=�0H=��G=�G=yG=�WF=qlE=dD=UC=wYB=�A=��@=r@=�@=��?=�n?=d�>=1#>=,==�<=��:=x9=7:8=� 7=�>6=$�5=�J5=�25=H5=�u5=��5=־5=i�5=�o5=%�4=�N4=ч3=A�2=��1=ln1=_1=5�0=�0=��0=�0=�10=��/=x�.=A�-=��,=��+=^�*=��)=E)=�s(=f�'=�'=�1&=|%=�#=c�!=�=PE=��=:`=G�=|�=5�=��=y�=�^=��
=r-	=u==�=j=�:=���<��<V��<i��<T��<݄�<���<�$�<�n�<!w�<��<�R�<�"�<o��<~�<㫸<I��<;Ԯ<���<��<J�<��<9�<<��<	��<7M�<:��<>��<��u<�+j<�W_<TpU<\�L<��D</�=<%Q7<51<y�*<5$<��<�<�<{s<���;��;�]�;�;O��;ȟ;���;��;%	f;��B;m�;�(�:4M�:��9T~��H g�E������"���=��]���#��>h������һ�U�p��,
�de�5l��"�:l'���+��E/�Bj2��}5�8�8�ڊ<���@��rE�TEJ�V�N���R��3V�0jX�üY�xZ�� [���[�5]��_���a��e���h��]l���o��r�P�s���t�wyu�C>v��xw��ry�>O|���J7��|����
��4Q���E��tƌ����r/���3��� ����<���'��sp���)���R��Ր������:��t����ݖ��������W�������5��'��k�����0��j8���A��X��iu��}��<��=ᨼ����F���j�������;��3̲�:���'��o��������8��U<�����nٿ���������Tt���  �  �N=�5N=�M=� M=�&L=<K=TZJ=�I=^I=ˢH=�aH=q.H=��G=F�G=�G=�LF=�eE=icD=G\C=hB=��A=��@=܍@=>:@=D�?=J�?=p�>=^5>=�===�<=|�:=��9=�U8=�?7=	`6=��5=k5=�O5=ja5=��5=	�5=��5=+�5=��5=�5=g4=��3=4�2=�2=N�1=V!1=k�0=��0=?�0=m}0=D%0=-�/=��.=g�-=��,=-�+=��*=��)=�3)=L�(=D�'=J5'=�H&=%=K�#=��!=�=�\=�=.=�=��=��=1�=i=ez=��
=�C	=E�=��=��=fT=S��<{��<���<�)�<���<K��<���<�&�<3c�<�a�<5�<�8�<#�<��<�!�<;��<c��<� �<OŪ<�ަ<��<VG�<�0�<���<�Ǒ<�n�<���<Q�<v<�j<��_<��U<s"M<�DE<%7><��7<�s1<e+<�_$<�<2�<�.<<�<���;��;�2�;a��;�d�;p�;|��;¼�;�6e;��A;��;���:+Պ:���9$���u�b�H,����������(<��[��~�����q����#һ˧�i��� �	�������g�!���&��W+��.� 2��85�ԇ8��@<��v@�eE���I��zN���R�u�U�M#X�̔Y��nZ��[���[�65]�?4_���a�,e�Z�h��8l�Ko�J�q��Us�Xt�eu���u��!w�L%y��|������ur���؆�(��4������{�������l���Uc����n��`L��S���%�������Q��+��Ԅ��:���)�������W��R���+K���4�����/0��"���/���)��B䤼�C��F��M������Iq���~��񫼯ҭ��������R����]��g�����Z����G��������_���O���  �  ��N=�hN=Z�M=�@M=�mL=��K=��J=��I=<I=��H=�mH=�%H=��G=(oG=j�F=,*F=%OE=�^D=ImC=ݎB=��A=�CA=��@=|�@=0@=q�?=j.?=]g>=�n==$M<=�;=^�9=�8=��7=��6="6=�5=��5=��5=��5=7�5=K6= �5=i�5=rG5=��4=��3=�"3=�d2=@�1=�P1=q1=m�0=`�0=�_0=��/=$s/=�.=�-=��,=��+=��*=�0*=�~)=��(=~;(=t{'=��&=�N%=��#=��!=��=��=2?=s�=�{=�<=7&=`:=�s=��=�%=�	=��=��=��=v�=�n�<׀�<���<���<+:�<���<��<%�<;�<��<C��<z��<a��<$��<�+�<���<#�<7{�<�P�<�l�<,��<���<��<��<<$�<�ό<i/�<�f�<W=w<��k<�Ya<j�W<��N<f�F<�{?<n�8<�l2<I�+<�9%<2�<��<UA<�<UA�;uv�;�_�;�^�;�s�;�G�;�I�;xԁ;��b;��>;1<;6F�:$O�:q:�9�lo��_V��n���*��EG��?8�oX���z��F��������x[л�滘K���J��x��w��1 ��%�8?*�d.�O1��y4���7�Bu;��?�kD��H�MM��oQ���T��gW�6+Y��]Z��P[�d]\�9�]���_�eb��pe�v�h� �k���n��p��1r��&s�j�s���t�?3v�`Qx�}C{���~����$����J���t���Q��Iŋ�t����?��]���4���쌼��������錼Ǖ��g������T����j������;��-���ؗ�9\������􍙼ق���̛�xf��8�����|ꢼ�|��x�������k������屮��q���<q��E���95��vѴ�&^��%���k����6��z@��վ�y�������꾼�  �  w�N=��N=�9N=ŗM=T�L=��K=VK=�8J=��I=��H=WxH=dH=�G=�/G=h�F=~�E=-%E=oPD=�~C=Q�B=, B=��A=tAA=[�@=r�@=<@=�x?=H�>=��==�<=Kg;=�7:=�9=�8=gJ7=!�6=XN6=�6=�6=�$6=�;6=-G6= 76=[�5=r�5=�5='P4="�3=	�2=%2=U�1=�"1=H�0=
�0=�*0=޽/=�0/=D�.=w�-=�,=�,=�<+=��*=r�)=nJ)=U�(=�'=�&=��%=j$=�B"=8 ==��=�[=~=��=e�=��=��=�8=��=��	=B=�/=�'=��=�=�<1^�<�m�<���<��<kr�<�4�<��<���<��<
%�<9b�< f�<gH�<�+�<�4�<0��<d�<o�<w.�<�Y�<�d�<�+�<��<J��<�W�<�͇<N%�<�y<�n<Ɠc<w�Y<X�P<��H<s`A<�u:<��3<;;-<_f&<�<�:<��<A�<���;��;sK�;F��;{��;���;��;b/�;vE^;:;��;���:1�:���9�qJ��eF�p����b����2�E�S�O�v�Sg�������	����ͻ)��<���XM��U��L�����#�D�(�Ϡ,�%0�Aq3�K�6��b:��Y>�W�B�1G�`�K���O�
�S�erV���X��aZ�f�[��5]���^���`�hDc���e��h��ek�©m�jo���p�n�q��Rr��^s���t��2w��7z�z�}����UE���v�����MC������k���$6��fo���h���@�������b�����M��\���򚒼�5��q����Ö����Jr��//��4��p
���M��ɝ��h��:����������
��7䥼�����W���>���p��d����물�&��5����� ��ڴ�� ��� ���*���ӽ��)���F���K���\���  �  �4O=u�N=��N=l�M=�0M=�XL=dtK=D�J=��I=RI=�tH=A�G=%_G=��F=�:F=��E=��D=N/D=�C=��B=KjB=>B=��A=cTA=��@=k@=K�?=:�>=��==��<=��;=�:=��9=�8=$�7=6[7=��6=��6=1�6=��6=K�6=��6=�w6=B6=��5=v^5=%�4=/�3=�.3=Pq2=/�1=a91=J�0=�K0=6�/=^/=u�.=0.=��-=#�,=�,=u+=�*=GL*=��)=;)=3=(=�3'=��%=�[$=�"=�� =�q=:=��=��=+�=%v=�w=��=L�=��=U0
=�a=�}=�z=(S=� =rA�<+S�<�b�<֊�<=��<�O�<{��<p�<��<&Z�<b��<V��<u��<��<�_�<��<῰<�ɬ<��<3�<��<W��<��<��<�<z�<���<{{<vp<�Af<y�\<�S<YK<P�C<�X<<�b5<ډ.<^�'<�J <ׄ<�.<�P<a�;�"�;K9�;���;cɱ;(N�;
�;�Y{;��W;EB3;\p;���:��:���9�v/��7������Qݺ�����-�IO��s������蠻 鵻�3˻=F�ߣ�������
��l��g�!�c�&��+�5�.��h2���5��_9��.=�\LA�ݥE�J��TN��7R���U�vXX�q�Z�|�\��{^�n\`��bb��d��f�di�k�K�l�� n�+o���o���p���q�8�s�� v��5y���|�Fl���|������^������*T��mQ�������V���|������N����������v���a��F���!���Ǒ��r��\���f�����O�����������Bϛ�
��Y`��������^��vs���W������ȥ����������ڨ��z��j��{����簼�<���y��a����N��Oú��ܻ�g���m��@j��;����ʽ��  �  (`O=�O=��N=q)N=zM=ΪL=`�K=��J=��I= I=�XH=r�G=��F=�WF=	�E=VE=�D=��C="qC=��B=��B==LB=��A=�A=5A=�@=,�?=C?=O!>=�==0<=";=l/:=�[9=ϥ8=�8=e�7=nI7=D7=��6=�6=r�6=:�6=�l6={6=�5=5=nH4=~3=ϰ2=��1=�81=�0=p�/=�l/=��.=aQ.=w�-=G/-=��,=�,=��+=R+=˞*=*=�b)=�(=?p'=<&=��$=K�"=� =��=��=r�= v=S=:=t.=.1=kA=�\=�~
=.�=�=�=9�=uY =���<�<��<H�<��<;�<4t�<[��<��<JP�<��<p��<�>�<���<IZ�<�.�<93�<�W�<���<H��<�o�<1
�<�[�<�k�<LK�<��<�΃<Z3}<,�r<�i<˚_<J�V<�N<S�E<e/><2�6<C�/<
q(<2!<ql<�A<:�<��;���;{�;G)�;��;�J�;}��;�xt;�O;fY*;e;�ÿ:X�l:+��9�0-�/��ۖ�M�Ժ�	��?*���L�Y�p�����fɟ�-L����Ȼy�ܻEp�1s�z
�������J�$�$���)�s�-���1�7;5�y�8��l<�U@�l|D��H��M��@Q�>U��aX��P[���]�7`�W[b��dd��Wf��*h���i�+5k�Tl�.m�]�m��n���o���p���r��ru���x��|������ ���4������(ꇼBꈼ�����7������JԊ�����8��������I�^������l!���ے�唔��6�����G��7d������
Ҝ����+1���R���_���O��T��Wϣ�s���#�����z���x��$'�����3+���Q���o��s���L�����V��7|���b��������_����Z���  �  �gO=�O=ƹN=7;N=?�M=�L=��K=9�J=T J=0	I=H=�BG=�xF=L�E=GE=��D=<	D=Y�C=�>C=��B=�B=qB=P)B=}�A=IQA=�@=��?=C?=�+>=<==�S<=�x;=`�:=��9=�Q9="�8=eA8=��7=}7=
67=c�6=!�6=�6=9o6="6=y�5=H%5=�s4=��3=��2=��1=�1=�L0=��/=��.=:F.=0�-=�5-=��,=W,=��+= �+=f9+=��*=�A*=��)=8�(=u�'=m)&='�$=��"=!=r0=�9=+6=X(=�=��=o�=m�=z�=\�=�
=��=�=��=��=>� =�\�<�z�<mj�<�?�<��<���<���<E��<���<��<�\�<���<�c�<�%�<��<*�<V]�<���<���<J��<���<j�<�T�<q�<*t�<�q�<�v�<E<~^u<]�k<^~b<?`Y<G�P<L�G<��?<W�7<s00<��(<�P!<	�<6�<�,	<�% <�J�;���;���;�X�;�L�;8v�;��k;|]E;_�;���:/U�:qdR:Q�9��L�d5/�s����Ѻ
L�pb)��lL�qjq�/ ���ğ�f���$5ǻlFڻ`���;��Dq�>A�����)�-#�\�(��F-�u1��85�"�8��R<�"@���C��)H�׀L���P�1U�[�X��s\��_�P`b�M�d���f��h���i���j�~�k��[l�S�l��:m���m�e�n���p�ߵr��hu�ւx�n�{�e/�6������!���g������
���&r��3��cӉ�?V��q���E!��������d׌�����s4���ɐ�~����l��I�����FÙ��R��.������3��D9��o��ޡ������������q���Ϥ�����7j���#�� �������ﯼ̱�Ɗ���'��i���9����)��(8��#���뻼̕��)���  �  EO=!�N=�N=�N=8�M=G�L=��K=-�J=>�I='�H=m�G=�F=%�E=RE=�lD=��C=NxC=)C=��B=��B=�B=\kB='B=��A=A=A=��@=g�?=��>=�>=e5==�n<=�;=;=|:=~�9=i\9=�8=UK8=q�7=�a7=�7=��6=�~6=�C6=#�5=��5=�5=Pp4=M�3=2�2=��1=-�0=	�/=�/=�E.=��-=�	-=H�,=;,= �+=ϳ+=�v+=�.+=%�*=DD*=t�)=�(=�f'=a&=�$=|�"=�'!=�e=��=��=��=2�=��=<w=�A=�=��=p�
=�=��=��=˞=Mx =�a�<+��<�r�<)�<��<	W�<���<���<��<��<���<J��<KX�<�[�<A��<�۴<�5�<À�<��<琥<w=�<ή�<��<�"�<RQ�<��<��<�F�<�fw<�Bn<-e<��[<ϱR<�I<��@<UO8</0<f(<�� <4<�V<�	<�$ <Z�;�b�;X��;���;f�;[n�;{�a;Y:;%�;9�:~'�:,x1:��R9<Ȇ���8��F����Ӻ��	�Ł+��KO� �t�����Y������ƻ�oػ���9��� �����S�!b���!���'�S8-��1��5���9� �<�[z@��6D�R@H���L�DQ�	�U���Y��^���a��d��g���i��k��l��l���l���l�7m��Gm�b�m�`!o��p��Is��v��"y��5|�!�瀼����=��#M��'U��<\���a���]��&H����9Ȋ��Z���݋�:j��s�����hF��	ΐ�Ԙ��!���נ����������n��"
��	j��D���#l�����$�������GG������-!���٤�'ۥ��(��?����z��2P�����*ү�bc��_ղ�0/���y������k���.9��{e��Kz��)p��C���  �  ��N=ݜN=R?N=W�M=�LM=�L=��K==�J=@�I=ӃH=:[G=#AF=�AE=VfD=j�C=t4C=��B=B�B=7�B=�xB=�eB=�@B=��A=��A=��@=�F@=�u?=�>=��==�==5i<=��;=_;=�:=�g:=��9=�E9=̤8=?8=n7=��6=�6=|26=X�5=�5=YW5=��4=�C4=m|3=7�2=R�1=V0=|u/=�|.=��-=\�,=.V,=w�+=�+=�{+=�Z+=�7+=�+=#�*=p*=�X)=�W(=O '=޼%=<$=�"=�!=8z=f�=�=�F=O=/2=;�=��=7C=��=��
=3~=�k=�f=�^=�C =��<�H�<�.�<���<�>�<���<���<e~�<�5�<Z6�<.��<�8�<�2�<�m�<�շ<�R�<Cɰ<��<m7�<�<���<��<$F�<�<��<`m�<[�<�ɀ<Q�x<WAp<�?g<��]<�kT<W�J<�fA<IH8<��/<du'<�<�<�T<�2<\��;�(�;�;K��;` �;"�;��;�3W;#F.;Բ;���:�Є:-:)��8�ȳ��$J������ںo��T.0�ѱT�L�z�(w��W^��,�����ƻ��׻z绵��Y;���
�����+!��'�d�-�9�2��7���:�?>�L�A��E���H��=M��Q�A�V��X[��_���c�|g�Rj�dl���m�l[n��~n�vLn�9�m���m��m�מn���o�a�q�L�t�6dw�jYz��#}�H��p׀����U����h��T���^��쇆�����z���������ۋ��}��6��㴍����<���#���쒼:���
/��Oo��˝������{c���ՠ��˱���,��
r��4���[���u���[s��T6���N�����\��o ��s⬼��������8��nZ��kn�����������	���q��⹼�F������H����  �  ��N=y4N=q�M=IsM=�L=�UL= �K=نJ=�cI=*H=��F=��E=��D=�C=C=W�B=vFB=�%B=�B=\#B=�B=< B=غA=�GA=,�@=T�?=?=5>=6q==��<=�L<=��;=�;=3;=��:=�?:=8�9=d�8=28=vb7=m�6=�46=^�5=��5=�E5=.�4=1�4=!�3= <3=/N2=Q?1=�0=��.=��-=� -===,=��+=�N+=�+=�+=��*=�*=��*=Ek*=��)=b)=�(=��&=uZ%=��#=�c"=o� =u=��=�a=ѧ=ݽ=��=�Q=w�=#_=��=<z
=u4=�==�=o��<Q��<��<��<�M�<���<���< �<�U�<���<���<�2�<���<}�<[{�<y�<.��<6�<���<���<�Z�<�ן<�(�<�m�<qɑ<W�<k�<h�<��<w"z<��q<�h<܃_<r�U<��K<ޔA<]�7<<�.<�'&<�0<�<��<��<���;70�;��;��;��;�E�;&y;mM;�;#;���:7l�:��`:��9��ѷB]��>_�l.����{��O6��|[��ڀ��铻^W��ּ��KȻ�[׻�"�C�������m	��>�r��� �C�'��w.�4�|�8�%�<��?��C��eF��J��EN���R���W�:�\�[�a��-f��i�*�l�Ao��9p�Ûp�gp���o��;o�P�n�,�n��o�T5q�-hs�[v��y���{�=h~�s4��J�������*��꿂�Đ�������腼b\��݈��J������Z���TI���㍼�}���=���E��é���m��9���W֗�g?������ɞ�5���,��"?���飼b>��BV��YQ���S��?�������.ƥ������v���,��[�����D��;G���>����沼�ӳ�����}Q��:㷼����9D��ռ�?-���  �  �DN=��M=�nM=FM=a�L=�	L=~@K=�CJ=3I=��G=A�F=yHE=$&D=�3C=�|B=�B=�A==�A=��A=	�A=��A=y�A=�tA=B�@=N@=`�?=أ>=v�==c==��<=.'<=��;=�;=�e;=�;=s�:=��9=T9=�(8=fK7=�6=��5=:o5=�5=�4=w�4=Q>4=*�3=��2=�
2=%�0=3�/=��.=@x-=�{,=��+=�+=��*=*�*=��*=ۢ*=|�*=�~*=�**=ڗ)=y�(=��'=~`&=��$=Ä#=�"=� =kb=�=̍=��=�
=��=|�=�=h=��=6D
=��=ֵ=ŧ=��=�A�<���<O�<�>�<���<j	�<q�<()�<X[�<���<���<�<���<�"�<N��<\�<Y�<֤�<���<���<覣<0�<iT�<֚�<�
�<���<p��<g�<�<�<��z<��r<j<��`<ہV<�L<��A<KK7<\�-<��$<��<�<�y<��<��;��;���;�G�;�y�;��;U�q;��D;!;���:�:��>:���9� �	�)(s�㳱����8��SX<��b�7L���?���B����xKɻ��׻�h�hB�� ��f��\�p��(� �"`(��W/�_S5�T=:�s2>���A�܏D�X�G��AK��WO�g�S�;Y��=^�[c��h�3l��1o�.Gq�Ur�9�r��r�f<q��ip���o���o���p�d|r���t���w�%�z��q}�
��|����,������ׁ��N��V
��7��g��"���߈�����	���5�����Ĵ��WE����}䐼�6��L󓼍��Tr��f���u��������`H��SW��Q祿�&���������#䤼_���}��+\�������6���������3\��K���Φ���^����x����X��`l��Ե������l���\���-�������  �   N= �M=#M=\�L=�aL=��K=�K=LJ=[�H=��G=PHF=��D=��C=q�B=�B=��A=�sA=$mA=,�A=��A=��A=��A=lAA=��@=�@=8?=�W>=��==g�<=YX<=�<=V�;=$�;=b�;=�,;=b�:=i�9=9=�)8=�67=�Z6=��5=�'5=c�4=~�4=�W4=4=H3=N�2=��1=��0=��/=�R.=g(-=�",=]R+=K�*=qo*=�Q*=SV*=.g*=�l*=O*=i�)=�d)=׆(=�h'=�&=$�$=&@#=Z�!=֑ =6P=	=J�=m=�7=�=�=@=4h=��=G
=��=�p=�_=�c=&��<���<���<���<�k�<2��<���<ח�<ʳ�<��<n��<�T�<?4�<߁�<5�<�<Y��<I=�<l��<�<9%�<?��<ݺ�<u�<0�<`P�<�u�<�ׄ<(L�<.F{<�ds<v�j<�7a<�V<	:L<�_A<��6<��,<6�#<N�<��<�g<��< ��;��;�m�;^��;N��;h��;,�l;��>;��;L�:_�:Y(:��\9"�G��W�ۋ���y��D���3c��@�s�f��ǆ�i���	e�������Mʻs�׻��l�"A ��������?��� �x�(�90��F6�`;��g?���B�˥E�:�H��L�� P�~�T�B�Y�@._��qd�Pi��xm�q�p���r�F�s���s��%s�^/r��>q���p���p���q��ls���u���x���{�8�~�!T��( ��[��Y������K������σ��D������눼�Ɗ�*j��&���򦎼�M��0׏��v��OY�����U���r��iߘ��t�����fi��ts��������
���¥����xl���J���g��7⥼�ʦ�����©�ݑ���X��o箼1��� ~���豼a��8����������U��]��0w���t��5+���  �  J�N=�hN=�M=peM=�L=&L=�SK=W\J=hEI=�H=�F=�E=R�D=��C=3#C=g�B=;PB=)$B=B=OB=��A=s�A=tA=�A=�l@=8�?=�?=�M>=ި====f�<=h[<=P<=r�;=dI;=y�:=�:=�R9=C�8=��7=Q�6=�J6=��5=�O5='�4=�y4=8�3=yV3=:�2=d�1=B�0=�/=�c.=�U-=we,=Ɯ+=� +=e�*=H*=r*=��)=��)=2�)=)=.w(=��'=�&=Ak%=�$=_�"=�`!=s =/�=<=��=�=�==C1=�=�=�=��=m3
=��=�=��=�q=E��<�*�<�r�<�m�<��<��<���<uH�<���<|�<��<���<���<��<P�<�ٶ<)i�<w�<,�<�;�<��<���<{4�<^��<�S�<��<a�<�.�<�X�<��|<:�t<��k<�b<]�X<��N<��D<;�:<�r1<�(<�	 </�<(�<�e<�?�;&��;��;M{�;~��;�L�;(S~;�^S;��*;o�;>�:���:�:���8.����;�X����1Ӻ�	�8�+�>�N�C�r�R���1���]��������ɻw�׻[�����b��	����%�������&�Ò,���1��56��0:�L�=���A�Q�E��J��N�?�S�K�X��r]�e�a���e���h�g k�e�l�i=m�X]m��,m�9�l�&�l��Lm��=n���o�E�q��5t���v�� y�&8{�4�|�{'~��,�;��u���􈁼�������}��K��`���t#���^���f��L���)������G�������t���w��W�������B���]��42������QƢ�‣��꣼k��6���X��墤�`+������w��w��E����w���ᬼK�� ��/񯼕���!m��.S��~r��}Ӵ�Ho��02����������B���  �  SO=�xN=�M=�wM=��L=s6L=wcK=�kJ=~UI=-+H=��F=��E=��D=*�C=�:C=��B=ofB=�8B=l"B=:B=��A=��A=��A=hA=z~@=��?=�?=&]>=�==�&==g�<=OY<=�<=b�;=$=;=˲:=�
:=vJ9=}8=v�7=$�6=�T6=��5=e`5=i�4=�4=K	4=�f3=͞2=�1=��0=��/=Nw.=Xk-=,|,=/�+=^+='�*=�]*=�,*=�*=��)=��)=%)=��(=E�'=(�&=�|%=.$=��"=�j!=p =��=�6=�==�.=�"=R�=��=�=i�=F8
=��=Ź=��=m�='��<�G�<���< ��<m;�<��<�<xo�<���<���<���<�(�<���<6�<y�<���<��<\�<4O�<`�<�4�<|ן<�[�<ܖ<q�<�.�<�<�.�<�N�<.�|<�t<��k<��b<��X<'�N<o�D<��:<��1<��(<�A < <=�<T�<O��;���;��;���;��;��;�;'�T;f,;�";�+�:�Ņ:�l:� 9{���/7����к���h*���M�(�q�����V�������b���ɻ�׻���U�����J2	�p��u�����F&��f,�H�1���5�6�9�դ=�lA��mE���I��nN�WS�QX��#]�S�a�)ke���h��j��1l���l�Bm�0�l��l�&�l��m���m���o�_�q���s�Auv���x�l{���|�M"~�T;�'��Pˀ�4���ݷ���
��ڋ���!���������6G��5H��)��N��c���<&������qU���W��Ō��#ؙ�����1�� ���}������S������C���g��h8��������ޥ������R���Щ��V��Ǭ� 
����������@���j�� ���?봼����=��x�������0���  �  d)O=ȤN=�(N=�M=dM=cL=3�K=8�J=y�I=�ZH=�0G=WF=^E=d0D=CC=�B=�B=�qB=�UB=�BB=8)B=9�A=�A=v?A=ƭ@=@=�D?=��>=��==3<==e�<=�Q<=�;=��;=p;=�:=��9=�09=wo8=��7=97=�q6=�5=��5=�)5=�4=R74=l�3=!�2=��1=��0=��/=ͭ.=v�-=�,=��+=.\+=�*=�*=�c*=�7*=D*=(�)=N)=��(=)�'=��&=��%=WY$=��"=��!== =�=#&=�=��=�=�=�=�k=�=ם=F
=�=��=I�=ͬ=��<���<��<u��<ۋ�<��<�t�<���<`i�<�/�<�E�<$��<Nz�<ݒ�<�<�f�<��<�`�<٫�<࿨<嘤<J>�<���<�9�<Ⱦ�<�d�<	5�<�(�<�+�<QF|<��s<$k<��a<�LX<wN<_�D<�
;<��1<�,)<J� <&�<�<�R<Q�;VA�;xM�;�P�;ߗ�;n��;��;��X;��0;W�
;�:�7�::$:JI9Kvp�Z�*�������ʺ�Z�"'�'YJ��Pn���5���}K�����1ʻg�ػ��滻l���"�6�	�yN���L���>&�K�+���0�Y65�V!9�u�<�ް@���D��I��M�A�R���W�#H\��`�Qfd�pg���i��+k���k��0l��l�E�k���k�Fel��Nm�l�n���p��*s���u�[Fx���z�(�|��~��k��W�����~큼���I�������3��Ӣ��<퉼A����ˌ�N���e����ˏ�BA��� �����D0��Fr�����������������w���Ӣ�~J����������ߣ��.��ܶ��z�������#��p�������|��b֭����������ְ�Ƕ��򰲼	س��2������aa��9
��!��������  �  2ZO=a�N=�iN=��M=�RM=��L=}�K=��J=ҽI=&�H=N}G=^iF==oE=/�D=�C=�bC=�C=v�B=n�B=m�B=wdB=�3B=��A=�zA=��@=B@=�?=v�>=^>=�W==;�<=$A<=-�;=X;=��:=bM:=9�9=_9=nU8=��7=x7=ח6=$,6=��5=�j5=��4=<t4=��3="3=	2=�1=�0=��.=�.=5 -=u`,=��+=�L+=��*=��*=�}*=�B*=6�)=�)=h�(=�(= '=��%=S�$=%#=��!=�" =��=k=�b=t�=^�=�=M�=<=��=>�=�V
=�)=l=��=��=&��<��<YC�<=�<��<o��<��<��<Q$�<��<s�<��<�D�<rK�<���<���<rq�<\ݰ<�&�<�>�<��<Ƞ<nJ�<g��<�'�<ɫ�<�P�<q�<��<w|{<��r<rj<z�`<moW<~�M<dYD<�;<�C2<��)<ڵ!<��<Ɲ<�9	<_ <���;��;�/�;��;��;���;�B_;�W7;��;��:�	�:�M;:-�9#:&�V���|��_�º�%�r�"���E���i�)��	���^H���º�uvʻ�ٻot�G����b�
����
!�t����%��P+�0��84�m8���;�L�?��C��3H���L�=�Q�KoV��[�w6_�Z�b���e��
h���i�΃j�n�j�0 k���j��k���k�ril���m�w�o�1&r���t��lw���y��4|�� ~����<����~��l���~��򵄼����Y��K���z�������A����K���!�����T���ϐ�r����������tߘ�������ǳ���!���?���������*���e������wF�����(!���p��C屮턪�"��ّ���⮼�	��������(���W��������������!��N���U����  �  �O=�O=��N=�(N=��M=��L=��K=-K=��I=�H=��G=��F=��E=�E=ZlD=��C=�wC=#+C=f�B=w�B=i�B=kB=B=�A=�)A=s�@=��?=�>=�0>=�o==�<=�"<=��;=�;=�:=��9=�]9=0�8=]+8=��7=�#7=��6=�`6=�	6=m�5=�:5=�4=4=q73=�P2=�W1=W0=�Z/=�n.=*�-=�,=�F,=��+=�b+=�+=��*=�*=b,*=��)=�)=O(=Q'=+#&=��$=WT#=a�!=P* =��=,�=>=[G=iY=�N=J+=��=F�=Ї=�`
=sI=�<=�1=�=[��<�g�<���<*��<Gg�<�<��<�E�<p�<���<?'�<���<_=�<�)�<�N�<؜�<,��<#\�<��<Ѻ�<ᠥ<cQ�<PԜ<8�<���<�<^�<��<6��<Yz<<�q<��h<�u_<V4V<j�L<�C<5	;<��2<�t*<��"<l�<��<�
<�/<���;&��;�$�;?�;�ݜ;;�;wg;��?;�`;��:�ª:� W:.(�9,�����mi|�����f���dW�LA�Rqe�5���j��p\������D˻�5ۻ�������o������� ��j	 ��%�ʸ*��-/�~93�(7���:�)�>���B�.UG���K���P��2U�ǌY��~]���`���c���e�1�g���h�#mi���i���i�-,j��j�t�k���l���n�7#q���s� �v��[y��{�O~��3��+���������-���O���y��c���ʦ��J���Z��d��͋������#Ꮌ�b��>"������#���8���;��������:���=�� ��ơ��;��ɓ��S梼�K���٣�:���������n��(��+���XS��}ծ��3��Hs�������ϳ��	��nU��ѭ��s���Q���}�������  �  x�O=|HO=D�N=�WN=J�M=��L=�"L=F1K=�0J=),I=�-H=�>G=veF=~�E=��D=xkD=��C=ȓC=�HC=�C=��B=��B=�CB=@�A=rUA=�@=��?=�%?=qN>=�x==I�<=��;=JI;=ȫ:=�:=0�9=��8=,m8=�7=,�7=�!7=D�6=��6=-86=��5=0h5=��4=�(4=�]3=v}2=W�1=�0=��/=�.=V.=�o-=��,=�L,=;�+=�q+=x+=U�*=uW*=W�)=�<)=s(=�x'=4M&=�$=t#=��!=�! =(`=��=��=*�=H�=��=��=ț=�|='f=�Z
=VY=�Z=�V=UC== =ۥ�<���<���<���<!��<@�<S�<)��<��<AK�<��<EJ�<��<��<�7�<�x�<��<~��<��<��<���<�>�<<��<�ړ<��<�M�<��<���<�x<��o<w�f<�]<@�T<g�K<�C<��:<h�2<��*<(#<�=<�$<��
<�<���;/�;m��;�@�;���;�z�;�ko;I;��#;P+ ;��:I^t:Z)�9��޶4���$o��`����q��f�=���a�l���~B��kߨ�����̻zlݻ^��46��N$��a��@����z �a�%�?X*���.�#v2��C6��:��>�OPB�޴F��4K�K�O�~T�?X���[���^��a���c�I�e���f�2�g���h��i�%ti�fj���j�	Kl�	n��bp�os���u�B�x���{�
�~�襀�ҁ��낼����*��������m���Ј�:���4"��㾊�wm��mA��tJ���������ґ�R���̦��Ė��o��v!��n���w���1$��-��4砼
���l���z����������\T���U�����n������ o��1��&殼�~��[���W��R����뵼O-���g������#��������h���  �  ϴO=[O=#�N=�iN=H�M=9M=P.L=�CK={QJ=�`I=a{H=��G=m�F=Z/F=ˊE=�D=6lD=|�C=��C=�;C=��B=�B=�NB=e�A=vdA=5�@=�	@=�6?=�T>=�l==�<=��;=��:=8:=�9=� 9={8=�8=r�7=,N7=!7=8�6=ړ6=*L6=�5=2y5=^�4=D34=k3=��2=ö1=��0=�0=�P/=W�.= �-=�a-=��,=HG,=3�+=�S+=��*=Tl*=��)=C)=7z(=��'=�Z&=� %=z#=��!= =�&=�<=�I=�O=kM=�D=m8=�-=+*=B0=-?
=RQ=_=�_=<L=� =���<���<���<W��<��<-��<���<���<V �<Yn�<��<�R�< ��<n��<���<�͵<n��<�"�<?9�<*�<T�<�q�<Ș<���<�	�<�<O(�<sN�<�w<�m<�d<!�[<J�R<4J<��A<O:<�e2<��*<�=#<�q<cS<��
<=�<���;���;���;m��;6F�; �;W�w;IKR;0�-;�m	;�[�:
�:�|:|Z8�e۹�g�mp��W��V�"�;�]`�Զ���ԕ����:���{λ�3�k񻁏 ��#�@�H��;���6!��&�DQ*�<L.��2�]�5���9���=��B�zF���J�O��S�{�V��Y��\��N_�g�a��|c��&e�b�f��g��^h�	i�|�i���j�l���m�p��r��u�a�x�9C|�Px��<������ރ����~��� ���և������!���������E����C��$��[+���z��������}���K��w��6����4��ۗ��ߜ����G������堼�����5��΢��u��V?���:��q���㧼=����Y���;�����Vﰼ����n1��h������*���F���A��-��ӻ��w���  �  ͢O=�OO=a�N=�[N=��M=T�L=L=;;K=ZJ=��I=�H=�G=�RG=��F=pF=�pE=8�D=�HD=k�C=eVC=��B=��B=[;B=��A=�RA=�@=B�?=�*?=N@>=CI==-P<=�_;=��:=5�9=�9=Ir8=q�7=��7=�B7=n
7=��6=�6=��6=�A6=X�5=Pi5=w�4=q4=[3=ȏ2={�1=Q1=V0=�/=B/=d}.=R�-=�F-=e�,=a,= +=��*=^g*=�)=I*)=a(=m'=NH&=�$=�c#=��!=&�=
�=��=�=��=Z�=r�=R�=��=��=��=�
=;/=WF=HJ=�4=� =�o�<{��< ��<<��<���<d%�<1g�<���< �<�z�<9��<�B�<��<0O�<Y�<�<���<��<��<��<&ס<Te�<0��<vؓ<XЎ<N��<��<3<	u<Q�k<�9b<XDY<��P<	xH<l�@<�9<-�1<k*<��"<�(<l <�j
<�n<�A�;�>�;��;-�;�O�;�ؑ;�/;��Z; g6;��;�n�:��:��:SW�8��ҹQg�*N�����=��g<�o`�^؂��=��H���W�����л�h�2���ӱ��P
��M����A?��9"��&��*��}.�2<2�e6�t:�@)>��kB�`�F�Z�J���N�obR�B�U�dX���Z��D]�:}_�r�a���c��We�Z�f�h�8i��j�Qk�Ljl��n�SAp���r��u�[y� �|��=��9����1脼 ���(��g��7����5��{����뉼xD������X���3���M��ݣ��7)��Z̑�y�����W�������a��젚�؛�����9��D[��e���P�����>ܢ�����$i���`����������]���l{��]w��ۀ��<����g���$��ղ������?��r>�����᲻�2:�������  �  yO=�)O=��N=�0N=��M=�L=��K=�K=�LJ=��I=��H=FH=�G=-G=+F=�E=�1E=��D=+�C=(]C=��B=�tB=�B=S�A=z$A=*�@=��?=b?=�>=�==�<=;=�:=�59=�{8=�7==l7=�7=��6=��6=W�6=9�6=�\6=�6=[�5=�<5=��4=��3=�13=�t2="�1=�1=�0=� 0=�y/=��.=,R.=��-=@�,=6G,=ߖ+=�*=�K*=��)=�(=g,(=E;'=�&=J�$=�4#=�t!=.�=^�=9i=�H=�+=�=b==t3=�]=h�=��	=��==
=;=���<|��<�A�<Au�<7��<!��<�`�<@��<8j�<f��<ra�<
��<�<`Y�<h��<�:�</�<dʱ<3ƭ<Oʩ<콥<���<X�<�s�<���<�m�</�<��<%Q}<�s<Ei<�_<��V<��N<Q�F<&?<��7<��0<�)<b9"<�r<>><e�	<� <���;�4�;;��;o��;(¥;�<�;E��;* b;7>;�E;��:�Ɲ:��):�]�8+^չAm�Ғ��ސ����$>���a�Jσ�Od���z�������ӻ���
�������yb�"w�f���m#�ӑ'��b+��/���2�1�6���:�^�>��#C�sRG�/FK� �N��R���T��#W��ZY���[��]��`��Ib�?yd�Upf��h�h~i�Z�j��k�S*m���n���p�|s��v��z���}�<ـ�����q�������<��SD��P����|�+��G\��$�����뤋�J������s������������v��rd��2������dϙ�	����0���y���Ǟ��	���0���4�����,bɤ�����:妼@H���nͫ��ۭ�A��+��t;������Ƿ�0���V���;���廼Z`����� ���  �  AO=w�N=�N=w�M=�EM=��L=ӴK=��J=?1J=i�I=s�H=�yH=b�G=�pG=B�F=T.F=7vE=�D=��C=�TC=\�B=�BB=��A=�`A=�@=�R@=C�?=�>=��==M�<=׼;=�:=�9=P�8=@�7=�_7=��6=�6=�{6=h6=?\6=zJ6=�%6= �5=��5=��4=�_4=^�3=��2=KK2=B�1=,$1=W�0=�;0=��/=�B/=��.=��-=�7-=�k,=&�+=%�*=	"*=9n)=ڴ(=��'=a�&=n�%={�$=!�"=h2!=^?=�)=��=m�=W�=��=�=ɔ={�=��=�:=�}	=��=��=E�=a�=4�<�p�<��<��<z_�<���<@}�<5�<���<���<��<7r�<��<���<���<�G�<�ŵ<�{�<z]�<�T�<G�<�<���</�<q�<��<���<�6�<A�{<:q<�5g<�]<�T<V�L< �D<V�=<|�6<Ƽ/<��(<�G!<�{<:<̍<�(�;N��;/��;��;��;߫�;��;5�;��g;�'D;$;b��: �:�A1:��8�@�~Bw���������_y�.bA�	e��P��� ��nV��9����Tֻ�M���c��Ƃ��M�<3��F ��$�w�(��H,���/��3��7��;�d�?�D��,H���K�)O�.�Q��0T�4V�;"X�K&Z��Z\���^�9Ra���c��Gf��_h��j�X�k���l��,n���o���q�@Wt��nw�� {���~��z��Jx���P��vzB��/H�������p������fƊ�ߊ�U���q�����J����'��⅏�� ���~��m瓼�*���C��>>���.��I+��6E��K���C圼�Z��pП�I/��g��$t��Wc��uI���?��_��׹���Y���<���V�������ֲ�������7Ƹ��6���V���'��R���]���R�������  �  tO=�N=GJN= �M=�M=KAL=�yK=��J=J=��I=\	I=��H=�+H=a�G=G=tiF=S�E=M�D=�D=XFC=�B=�B=�A=�A=��@= @=(g?=�>=͢==�<=x;=�Z:=QL9=�Z8=��7=Q�6=;�6=�G6=�(6=6=6=�6=��5=	�5=�F5=��4=�4=�o3=��2=; 2=�1=�!1=O�0=qc0=#�/=�/=+�.=1.=�`-=�,=W�+=��*=�)= 5)=gs(=u�'="�&=��%=�G$=�"=�� =��=��=�= l=�8=n=n=�)=�Z=��=r�
=�8	=et=)�=^�=�|=D��<q��<�7�<���<�<��<>��<j�<J�<8�<֚�<g��<@�<�<�"�<B�<	��<�'�<N�<Eܨ<�ˤ<}��<�B�<���<v��<?}�<��<��<Rz<�o<��e<?\<�0S<�	K<l~C<�e<<�5<A�.<�'<U <��<4<g�<��;w�;�;�;��;�N�;�*�;�.�;��;�l;��H;5#;k��:���:XM5:"��8�������úDd��#�6�D�
[h�rG���2%��5�û�ػ���r���Im��!�������׊!���%���)�~+-�|�0�9y4�,m8�&�<�5�@�E��	I�H�L��O���Q��S��U� FW�e*Y�b][�	�]���`���c�zEf���h�þj�fl���m�p1o�o�p�^�r��;u�\Ox��{�����
�����@	��1���]�����iƊ��$���I���Q��[�����⋼)����v���������{��}璼�1���L���8������ӗ�����ř�3	��v}��?�������=��Ƞ���У��פ��ɥ�¦��ܧ�O0���ʪ������ͮ�����l��(���oƷ�+���O
���%��m輼8a������vؽ�����  �  &�N=K�N=�N=*�M=I�L=�L=NK=*�J=��I=GyI=�I=(�H=IH=c�G=>G=]�F=��E=�D={D=�9C=�B=��A=BgA=��@=]t@=��?=�:?=fk>=Yx==�h<=�G;=%:=�9=�8=N7=�6=JG6=

6=}�5=y�5=��5=��5=r�5=��5=-5=��4=�3=&A3=�2=L 2=�1=T1=�0=�y0=�0=
�/=R/=}Q.=�w-=��,=��+=R�*=>�)=)=cC(=q'= �&=�i%=L$=c�"=B� =]�=X�=k=S*=��=}�=��=F�=%=�d=#�
=�	=�E=
i=�j=*K=[�<��<���<�B�<��<(��<u��<@��<�~�<)Q�<���<~>�<�X�<YK�<'5�<\7�<n�<�<�<i��<bn�<�E�<�<�I�<r[�<�%�<]��<C4�<Kfy<��n<�wd<��Z<�R<� J<��B<��;<|�4<��-<W '<��<c�<�q<:�<��;���;#�;=<�;��;�d�;�ؗ;q�;s�n;1.K;��%;<��:�&�:%7:�6�8q���3��N�Ⱥ�)���%���G���j��/��o훻�z��tŻ�Tڻ�� ��w	��.�B��@��og"��&��I*�p�-�Rd1��"5�%9�(R=�#�A�z�E�ɬI��M��O�v�Q�B�S��7U�>�V���X���Z�F`]��J`�Yc��Pf��h��8k�m�3�n��o�r�q��rs���u�w�x���|��N���n���������Y;��ܝ�������G����������ڳ������;؋��6��ߌ�Ӎ�5��ph���֑��4���i��Zi��S8��B떼����wr��z��<��� A��M라(���,M���̢�����-���(��#���:��.���� �����$��rt��mԳ�3$��$D�����[�������%g���ս�w��I7��_j���  �  ��N=��N=N=�uM=
�L=��K=>K=U�J=��I=guI=�I=�H=�RH=]�G=�JG=�F=n�E=�D=�D=�4C=�yB=I�A=�VA=v�@=5b@=f�?=�*?=�[>=�h==NX<=86;=�:=��8=8=�67=]�6=:06=�5=i�5=]�5=@�5=�5=�5=�p5=d5=~4=��3=�/3=��2=��1=�z1=%1=��0=�0=U'0=j�/=�/= \.=y-=�,=��+=W�*=��)=��(=�1(= ^'=rp&=�W%=P$=�{"=V� =��=�=�U=7=i�=��=�=R�=�=3P=��
=[�=�5=�X=GZ=�9=���<�Z�<���<z&�<���<>��<��<���<W��<�h�<4�<�W�<Om�<Y�<�9�<�1�<6^�<�ϰ<Ѐ�<�]�<�I�<f"�<Kɛ<�)�<g;�<��<��<��<�y<nQn<^d<��Z<8�Q<ģI<�3B<:;<�{4<��-<��&<�`<��<�,<~r<	�;a2�;_��;���;���;�w�;��;BI�;�do;LL;}z&;�:-�:�`7:4��8�3��NɆ��ʺ�C�F'��H���k�F���<j��������Ż��ڻ�6�$#�j�	���<�q���"���&�|�*��.�Y�1�Ja5�-a9���=�f�A�PF�[�I�j:M�-�O��R�4�S�(U��V��bX�)�Z��4]��+`�<Kc�Wf��i��ek��Bm��n�C<p�!�q���s�*v��6y���|��o������ǲ�����Fi���̉��Њ�iu��eǋ�u݋��֋�[Ջ�����V�����L���`,��판�*����P��f~��qt��89��f▼�����[���`��駚�2-���ޝ������S��@ݢ�q.��M��EL���G��&^��T���W@��!���D��k���y���6M���p���G��x»�Wڼ�铽������5���Y��t����  �  &�N=K�N=�N=*�M=I�L=�L=NK=*�J=��I=GyI=�I=(�H=IH=c�G=>G=]�F=��E=�D={D=�9C=�B=��A=BgA=��@=]t@=��?=�:?=fk>=Yx==�h<=�G;=%:=�9=�8=N7=�6=JG6=

6=|�5=y�5=��5=��5=r�5=��5=-5=��4=�3=&A3=�2=L 2=�1=S1=�0=�y0=�0=	�/=Q/={Q.=�w-=��,=��+=P�*==�)=
)=dC(=q'=&�&=�i%=]$=~�"=h� =��=��=|k=�*=\�=B�=��=^�=i=f=��
=F		=�G=k=�l=9M=s!�<̓�<O��<F�<N��<��<ʆ�<��<��<�Q�<��<>�<�W�<�I�<3�<�4�<k�<��<O��<�}�<mj�<B�<�<.F�<�W�<�"�<���<�1�<�by<��n<�vd<��Z<R<�J<�B<,�;<��4<�.<Z'<�<R�<
z<V�<���;���;1�;�H�;��;�m�;kߗ;���;��n;�-K;��%;��:?	�:�6:�V�8����Tn��t�Ⱥ�K��&��G�k��@���������R�Ż�aڻ��� �|	��2�m������i"�&�K*���-�3e1�M#5��9��R=�v�A���E���I��M�$�O���Q�T�S��7U�H�V�ĔX���Z�K`]��J`�Yc��Pf��h��8k�m�4�n��o�r�q��rs� �u�w�x���|��N���n���������Z;��ܝ�������G����������ڳ������;؋��6��ߌ�Ӎ�5��ph���֑��4���i��Zi��S8��B떼����wr��z��<��� A��M라(���,M���̢�����-���(��#���:��.���� �����$��rt��mԳ�3$��$D�����[�������%g���ս�w��I7��_j���  �  tO=�N=GJN= �M=�M=KAL=�yK=��J=J=��I=\	I=��H=�+H=a�G=G=tiF=S�E=M�D=�D=XFC=�B=�B=�A=�A=��@= @=(g?=�>=͢==�<=x;=�Z:=QL9=�Z8=��7=Q�6=;�6=�G6=�(6=6=6=�6=��5=	�5=�F5=��4=�4=�o3=��2=: 2=�1=�!1=M�0=oc0=!�/=�/=(�.=1.=�`-=��,=S�+=��*=�)=�4)=hs(=y�'=-�&=
�%=�G$=�"=�� =4�=�=§=�l=$:=�=9=�+=8]=F�=��
=�;	= x=��=H�=|�=+��<$��<?�<h��<3�<i��<���<�m�<�L�<��<"��<���<R�<�<��<"=�<G��<c!�<I�<�Ԩ<3Ĥ<ϙ�<1;�<K��<���<'w�<8�<���<�Kz<l�o<I�e<\<�2S<fK<�C<kn<<��5<k�.<��'<�c <M�<�C<�<,6�;�(�;�V�;B	�;cc�;�;�;�;�;���;�l;��H;�*#;Y��:�W�:L�4:�T�8���~���#ĺ���nb#��&E�ڞh�y���ɚ��B���Ļ�ػ��� ����u��(��������!�H�%���)��--�/�0��z4�8n8���<���@��E��	I���L�S�O� �Q�5�S��U�4FW�t*Y�n][��]���`��c�~Ef���h�ƾj�fl���m�q1o�p�p�_�r��;u�\Ox��{�����
�����A	��1���]�����iƊ��$���I���Q��[�����⋼)����v���������{��}璼�1���L���8������ӗ�����ř�3	��v}��?�������=��Ƞ���У��פ��ɥ�¦��ܧ�O0���ʪ������ͮ�����l��(���oƷ�+���O
���%��m輼8a������vؽ�����  �  AO=w�N=�N=w�M=�EM=��L=ӴK=��J=?1J=i�I=s�H=�yH=b�G=�pG=B�F=T.F=7vE=�D=��C=�TC=\�B=�BB=��A=�`A=�@=�R@=C�?=�>=��==M�<=׼;=�:=�9=P�8=@�7=�_7=��6=�6=�{6=h6=?\6=zJ6=�%6= �5=��5=��4=�_4=]�3=��2=IK2=@�1=*$1=U�0=�;0=��/=�B/=��.=��-=�7-=k,=�+=�*="*=6n)=۴(=��'=q�&=��%=��$=i�"=�2!=�?=�*=� =��=
�=��=��=Ɨ=�=��=?=s�	=ƹ=)�=��=��=_�<�{�<}��<=�<7h�<@��<���<:�<{��<��<W�<q�<T��<���<;��<�@�<ս�<�r�<�S�<lJ�<@<�<7�<ੜ<��<��<B�<��<�0�<��{<u3q<h2g<Ѿ]<(�T<��L<T�D<��=<Y�6<��/<��(<�\!<5�<<P<�<�S�;r�;F��;@�;���;Ħ;'�;MA�;b�g;:&D;t;��:���:�q0:��8,�⹉�x�S���<�������A��he�A��`-��k���»xֻ(����p����uV�m:�xL ���$�O�(��K,���/�ȝ3���7�2�;�I�?��D�^-H�0�K�c)O�m�Q�1T�@4V�W"X�`&Z��Z\���^�BRa���c��Gf��_h��j�[�k���l��,n���o���q�AWt��nw�� {���~��z��Jx���P��vzB��/H�������p������fƊ�ߊ�U���q�����J����'��⅏�� ���~��m瓼�*���C��>>���.��I+��6E��K���C圼�Z��pП�I/��g��$t��Wc��uI���?��_��׹���Y���<���V�������ֲ�������7Ƹ��6���V���'��R���]���R�������  �  yO=�)O=��N=�0N=��M=�L=��K=�K=�LJ=��I=��H=FH=�G=-G=+F=�E=�1E=��D=+�C=(]C=��B=�tB=�B=S�A=z$A=*�@=��?=b?=�>=�==�<=;=�:=�59=�{8=�7==l7=�7=��6=��6=V�6=9�6=�\6=�6=Z�5=�<5=��4=��3=�13=�t2= �1=�1=�0=� 0=�y/=��.='R.=��-=9�,=/G,=ؖ+=��*=�K*=��)=�(=o,(=X;'=�&=��$=�4#=<u!=�=U�=�j=�J=�-==z=�=�7=~b=��=��	=��=�=� =	=g��<��<�N�<��<��<�<�h�<e��<�n�<���<�a�<���<�	�<,T�<s��<�1�</�<.��<��<u��<���<V}�<M�<_g�<�~�<c�<�%�<ރ<[E}<�s<�@i<��_<>�V<'�N<��F<�4?<��7<��0<u�)<�R"<P�<_Y<��	<�� <�;�c�;"��;���;�ߥ;�S�;Hς;j.b;[>;�3;���:�c�:K�(:\��8D'ع<�n��i���s���}�b�>�$qb�d������	࿻:�ӻ[����������m�������s#���'��f+��/��2��6�)�:�w�>��$C�SG��FK�d�N��R���T��#W�[Y���[���]��`� Jb�Hyd�\pf��h�l~i�]�j��k�U*m���n���p�|s��v��z���}�<ـ����� q�������<��SD��P����|�+��G\��$�����뤋�J������s������������v��rd��2������dϙ�	����0���y���Ǟ��	���0���4�����,bɤ�����:妼@H���nͫ��ۭ�A��+��t;������Ƿ�0���V���;���廼Z`����� ���  �  ͢O=�OO=a�N=�[N=��M=T�L=L=;;K=ZJ=��I=�H=�G=�RG=��F=pF=�pE=8�D=�HD=k�C=eVC=��B=��B=[;B=��A=�RA=�@=B�?=�*?=N@>=CI==-P<=�_;=��:=5�9=�9=Ir8=q�7=��7=�B7=n
7=��6=�6=��6=�A6=W�5=Oi5=v�4=p4=[3=Ǐ2=y�1=O1=V0=�/=>/=_}.=L�-=�F-=]�,=Y,=�~+=��*=Xg*=�)=J*)=(a(=�m'=vH&=V�$=�c#=Q�!=��=�=
�=��=N�=7�=�=d�=D�=2�=��=A
=-6=�M=�Q=�<=| =�~�<���<V��<2��<�<$.�<n�<���<��<�{�<���<)?�<��<jG�<��<��<E�<j�<Q�<"�<Tȡ<�V�<F��<~˓<�Ď<��<���<�~<u<�k<�9b<yHY<v�P<��H<�@<19<��1<'�*<�
#<wF<�<�
<?�<�y�;s�;�H�;�9�;�p�;��;gQ;��Z;e6;��;#�:���:Bv:Ď�8��չqi��=�����G�C�<�-�`����z��}-��8ս��ѻ����B���^
�~Y�o��YG�@"�^�&�R�*��.��>2�o6�
:�{*>��lB��F���J�.�N��bR���U�7dX���Z��D]�P}_���a���c��We�b�f�$h�=i��j�Tk�Njl��n�TAp���r��u�[y�!�|��=��9����1脼 ���(��g��7����5��{����뉼xD������X���3���M��ݣ��7)��Z̑�y�����W�������a��젚�؛�����9��D[��e���P�����>ܢ�����$i���`����������]���l{��]w��ۀ��<����g���$��ղ������?��r>�����᲻�2:�������  �  ϴO=[O=#�N=�iN=H�M=9M=P.L=�CK={QJ=�`I=a{H=��G=m�F=Z/F=ˊE=�D=6lD=|�C=��C=�;C=��B=�B=�NB=e�A=vdA=5�@=�	@=�6?=�T>=�l==�<=��;=��:=8:=�9=� 9={8=�8=r�7=,N7= 7=8�6=ٓ6=)L6=�5=1y5=]�4=C34=k3=��2=��1=��0=�0=�P/=R�.=�-=�a-=��,=@G,=*�+=�S+=��*=Nl*=��)=C)=Az(=��'=	[&=C%=�z#=-�!=� =�'='>=�K=�Q=aP=:H=�<=�2=�/=e6=�E
=�X=�f=�g=*T=�& =��<���<� �<���<���<A��<��<���<-#�<�n�<o��<O�<���<]��<���<µ<v�<��<g*�<��<�١<�b�<���<'�<���<�
�<��<�G�<�w<'�m<Ðd<d�[<�R<.AJ<�B<5&:<~2<��*<�Z#<��<�r<4�
<��<+"�;���;k �;Z"�;�h�;Q��;*�w;�[R;�-;�X	;"�:���:�T:cD8S�޹�i��h��@�����l<���`���������F���>��Y�λR`໗=񻁠 �n2�_L�~�����T=!�&��U*��O.��2�|�5���9��=�� B��zF�G�J��O�S���V�5�Y�6�\��N_��a��|c��&e�l�f��g�_h�i���i���j�l���m��p��r��u�b�x�9C|�Qx��<������ރ����~��� ���և������!���������E����C��$��[+���z��������}���K��w��6����4��ۗ��ߜ����G������堼�����5��΢��u��V?���:��q���㧼=����Y���;�����Vﰼ����n1��h������*���F���A��-��ӻ��w���  �  x�O=|HO=D�N=�WN=J�M=��L=�"L=F1K=�0J=),I=�-H=�>G=veF=~�E=��D=xkD=��C=ȓC=�HC=�C=��B=��B=�CB=@�A=rUA=�@=��?=�%?=qN>=�x==I�<=��;=JI;=ȫ:=�:=0�9=��8=+m8=�7=,�7=�!7=D�6=��6=,86=��5=0h5=��4=�(4=�]3=t}2=U�1=�0=��/=�.=R.=o-=��,=�L,=3�+=�q+=p+=N�*=oW*=T�)=�<)=s(=�x'=\M&=N�$=ot#=Q�!=�" =>a=��=q�=~�=%�=�=��=y�=4�=l=ba
=D`=b=^=�J=�  =���<���<��<���<���<�H�<9�<	�<��<�K�<{��<�F�<��<	�<�-�<�m�<���<��<Q�<�<���<0�<W��<	Γ<��<�C�<���<@��<$�x<O�o<,�f<'�]<��T<�K<s C<��:<��2<��*<:2#<n[<C<��
<q�<G��;i5�;Y��;$i�;ڟ;��;��o;
I;��#; ;�i�:πs:<��9��E�����p��P��,����x�8>>�4gb�����<��}��OA���̻]�ݻ)��W��Y2��m��J������ ���%�|\*��.��x2��E6�X:�)>�DQB���F�B5K���O��T��X��[���^�&�a���c�Z�e���f�<�g���h��i�)ti�ij���j�Kl�n��bp�ps���u�B�x���{�
�~�襀�ҁ��낼����*��������m���Ј�:���4"��㾊�wm��mA��tJ���������ґ�R���̦��Ė��o��v!��n���w���1$��-��4砼
���l���z����������\T���U�����n������ o��1��&殼�~��[���W��R����뵼O-���g������#��������h���  �  �O=�O=��N=�(N=��M=��L=��K=-K=��I=�H=��G=��F=��E=�E=ZlD=��C=�wC=#+C=f�B=w�B=i�B=kB=B=�A=�)A=s�@=��?=�>=�0>=�o==�<=�"<=��;=�;=�:=��9=�]9=0�8=]+8=��7=�#7=��6=�`6=�	6=l�5=�:5=�4=4=o73=�P2=W1=�V0=�Z/=�n.=&�-=�,=�F,=��+=�b+=�+=��*=�*=\,*=��)=�)=O(=Q'=O#&="�$=�T#=��!=+ =��=u�=�=qI=�[=�Q=�.=��=	�=�=�f
=�O=&C=|8=�$=��<(u�<B��<��<
r�<w�<ӫ�<L�<��<Y��<�'�<B��<�9�<�$�<�G�<7��<��<�P�<J��<�<���<D�<Jǜ<�+�<��<��<bU�<��<^��<
Qz<�q<A�h<y_<�;V<��L<��C<?;<ڪ2<4�*<��"<޵<��<�0
<J<���;��;�N�;�5�;���;��;�$g;�?;�^;���:M~�:�YV:2%�9�α�3E	�0�}�n��v���l��@�A�l�e�(Q����������Iۺ��o˻@\ۻk��m ��4|�A�����k��Y �۸%���*��0/��;3�7�3�:�F�>���B��UG�l�K��P��2U��Y��~]���`���c���e�@�g���h�-mi���i���i�1,j���j�w�k���l���n�8#q���s� �v��[y��{�O~��3��+���������-���O���y��c���ʦ��J���Z��d��͋������#Ꮌ�b��>"������#���8���;��������:���=�� ��ơ��;��ɓ��S梼�K���٣�:���������n��(��+���XS��}ծ��3��Hs�������ϳ��	��nU��ѭ��s���Q���}�������  �  2ZO=a�N=�iN=��M=�RM=��L=}�K=��J=ҽI=&�H=N}G=^iF==oE=/�D=�C=�bC=�C=v�B=n�B=m�B=wdB=�3B=��A=�zA=��@=B@=�?=v�>=^>=�W==;�<=$A<=-�;=X;=��:=bM:=9�9=_9=nU8=��7=w7=ח6=$,6=��5=�j5=��4=<t4=��3=!3=2=�1=�0=��.=�.=1 -=r`,=��+=�L+=��*=��*=�}*=�B*=1�)=�)=i�(=�(=1'=��%=��$=K%#= �!=k# =k�=x=d=)�=w�=��=D�=�?=��=��=q[
=�.=�=�=%�=R��<m�<�M�<�F�<��<$��<>	�<��<�'�< ��<��<���<	B�<%G�<:��<t�<9i�<(԰<��<4�<�<'��<�?�<<��<F�<?��<-I�<G�</�<�u{<R�r<;j<x�`<�uW<��M<weD<[*;<�T2<��)<b�!<)�<�<�O	<�t <A�;?-�;6R�;�կ;Z�;j��;�[_;\c7;��;���:�њ:�::���9�3*�}����p`ú���#�c:F�zKj��K��o+��r���麻v�ʻp�ٻ��_��"��
� � '�N����%��S+�
0��:4��8��;�6�?���C�74H�#�L���Q��oV�[��6_�v�b���e��
h��i�؃j�v�j�6 k���j��k���k�til���m�x�o�2&r���t��lw���y��4|�� ~����<����~��l���~��򵄼����Y��K���z�������A����K���!�����T���ϐ�r����������tߘ�������ǳ���!���?���������*���e������wF�����(!���p��C屮턪�"��ّ���⮼�	��������(���W��������������!��N���U����  �  d)O=ȤN=�(N=�M=dM=cL=3�K=8�J=y�I=�ZH=�0G=WF=^E=d0D=CC=�B=�B=�qB=�UB=�BB=8)B=9�A=�A=v?A=ƭ@=@=�D?=��>=��==3<==e�<=�Q<=�;=��;=p;=�:=��9=�09=wo8=��7=97=�q6=�5=��5=�)5=�4=R74=l�3= �2=��1=��0=��/=˭.=t�-=�,=��+=+\+=�*=��*=�c*=�7*=@*=%�)=N)=��(=.�'=��&=��%=yY$=��"=B�!=� =y�=�&=֕=�=U=��= �==n=y=�=iI
=
=��=0�=İ=n�<D��<r��<T��<��< �<$y�<$��<�k�<1�<�E�<M��<Wx�<я�<�<�a�< �<#Z�<ʤ�<n��<?��<�6�<���<q2�<��<�^�<�/�<�$�<�(�<�A|<p�s<�#k<��a<QX<�}N<�D<O;< �1<E:)<�� <j�<��<pb<�#�;�^�;�h�;�h�;���;ɡ�;:��;tY;�0;?�
;���:��:Ɲ#:'�F9
Gs��+�Z��RI˺|���e'�k�J�-�n��9�������h��,.���'ʻ��ػ+�滳}��*�Z�	��S�L�����JA&���+�p�0��75�i"9�K�<���@��D�I�g�M�|�R��W�FH\�,�`�efd�pg�ưi��+k���k��0l��l�H�k���k�Hel��Nm�m�n���p��*s�¼u�\Fx���z�(�|��~��k��W�����~큼���I�������3��Ӣ��<퉼A����ˌ�N���e����ˏ�BA��� �����D0��Fr�����������������w���Ӣ�~J����������ߣ��.��ܶ��z�������#��p�������|��b֭����������ְ�Ƕ��򰲼	س��2������aa��9
��!��������  �  SO=�xN=�M=�wM=��L=s6L=wcK=�kJ=~UI=-+H=��F=��E=��D=*�C=�:C=��B=ofB=�8B=l"B=:B=��A=��A=��A=hA=z~@=��?=�?=&]>=�==�&==g�<=OY<=�<=b�;=$=;=˲:=�
:=vJ9=}8=v�7=#�6=�T6=��5=e`5=i�4=�4=K	4=�f3=͞2=�1=��0=��/=Mw.=Wk-=*|,=.�+=\+=%�*=�]*=�,*=�*=��)=��)=%)=��(=H�'=.�&=�|%=&.$=��"=�j!=� =A�=#7=��=�=�/=�#=h�=܈=.=��= :
=��=��=��=z�=?��<�K�<m��<���<�>�<���<}�<Uq�<D��<p��<ݺ�<T(�<���<��<�v�<��<
��<� �<�K�<&\�<�0�<�ӟ<X�<Mؖ<�m�<q+�<h�<s,�<�L�<˸|<�~t<��k<ˆb<�X<��N<��D<=�:<�1<��(<_I <�"<Y<s�<1��;�;��;w�;�$�;��;��;F�T;�#,;.";� �:簅:�0::�9�5��^�7��ה�t#Ѻ����*���M�%�q������Л�����p����ɻ�ػ�滧^�����x5	�����������&�"h,�0�1�j�5���9�D�=�qlA��mE���I��nN�!WS�5QX�
$]�a�a�3ke���h�
�j��1l���l�Em�3�l��l�'�l��m���m���o�_�q���s�Auv���x�l{���|�M"~�T;�'��Pˀ�4���ݷ���
��ڋ���!���������6G��5H��)��N��c���<&������qU���W��Ō��#ؙ�����1�� ���}������S������C���g��h8��������ޥ������R���Щ��V��Ǭ� 
����������@���j�� ���?봼����=��x�������0���  �  �`O=��N=3N=��M=E�L=�7L=8cK=kvJ=�uI=�iH=a]G=�[F==oE=��D=��C=YfC=��B=�B=�qB=�>B=�B=��A=�mA=l�@=5u@=�?=�3?=x�>=��==�T==e�<=U<=��;=�m;=8�:=�]:=&�9=�
9=vS8=&�7=��6=�Z6=F�5=I5=��4=k<4=��3=��2=X$2=]@1=�I0=~I/=4J.=�V-=Dx,=�+=u+=��*=�*=)�)='`)=�)='�(=�(=`\'=��&=�%=�a$=�!#=��!=j =�=M�=�=�k=޷=��=w�==�=�=7L=�=��	=*�=W_=6:=&=���<_B�<���<��<��<,D�<���<A��<lz�<�y�<ó�<E0�<$��<f�<��<l�<�Ƴ<��<�N�<0`�<`I�<
�<���<a�<|�<BƎ<P��<'{�<h�<#�|<j-t<Btk<�eb<�Y<G�O<�F<��<<�3<1�*<1]"<��<Pw<��<���;E��;�i�;�!�;H^�;Qp�;���;o�d;>;�#;���:y�:�Y:�0�9񑃸��i�x��ٸ�������G>�'`�������ء�e��G^���λ	Dݻ���)$���`����������{%�}�*�-c/���3���7��+<�u@�a�D�(�I��/N���R�EW��[[���^���a��gd��6f��zg�Ph�'�h��Qi���i���j���k�
Im��)o��Nq���s�0�u��	x�� z���{�D\}���~��K��;?��uY��V�����X��Դ�����z&��j;���D��XR��qw���Ï��A����[Ӕ��і�Aژ��֚�ﰜ��W��ÿ��䠼Rơ�eo��j��T��Z����9��ޤ��������;��C��O���u���.?��$h��w���t��Vr��v���ò��	������/������H���z���  �  �fO=��N=�<N=%�M=��L=�AL=�mK= �J=�I=�uH=�jG=jF=�~E=ԯD=�D=lvC=4C=1�B=g~B=VJB=�B=6�A=xA=�A=�@=�?=�<?=�>=2�==HW==��<=`Q<=��;=�d;=��:=�R:=T�9=�9=bN8=@�7=�6=�^6=��5=�Q5=P�4=�F4=�3=L�2=�.2=/K1=/U0=�U/=�W.=ye-=��,=��+=�+=B�*=5$*=��)=hl)=?)=��(=�(=If'=�&=��%=�j$=�)#=��!=�m =��=��=��=�b=��=J�=�=*�=/�=;F=� =0�	=9�=�d=UA=@=��<�S�<j��<���<���<�Y�<��< ��<��<���<
��<�Q�<��<"�<e9�<���<�߳<0�<]f�<�w�<�`�<
&�<қ<�s�<m�<�Ύ<x��<`v�<�\�<�v|<t<"Fk<+9b<��X<�uO</F<��<<λ3<#�*<�v"<^<'�<��<���;�D�;!��;3w�;뻰;ٛ;A'�;��e;�&?;�:;���:���:��]:f��9v[P��L ��u�M���<������`=��x_�=����{��ݸ���^��s���ϻ��ݻ����t��������A����J���i%���*��?/���3�g�7�^<��J@���D�3UI��N���R�sW�� [���^��a��%d��e�e?g�(h�)�h�Z#i��i��yj�Y�k��m�P o��'q�
us���u���w�4�y��{�?o}�+
��^���T���n��쫃� ���`��t���c���i���,��u2��l>���b�����(-���ޒ�P����������ֺ�������7������à�+���qR���Ң��<������$��ɤ�$���˧���ܧ��0������E�7���f��]|��.����������pȳ����ˑ��U���������nt���  �  �vO=��N=&VN=��M=kM=�^L=׊K=�J=��I=,�H=?�G=n�F=^�E=��D=�1D=��C=?7C=��B=V�B=�kB=�2B=��A=:�A=�$A=@�@=��?=�U?=ۧ>=��==�]==��<=�E<=e�;=I;=[�:=�2:=Г9=��8=�>8=��7=��6=j6=�5=�h5=��4=�b4=��3=J3=
L2=Yi1=ku0=y/=�~.=�-=[�,=��+=�M+=��*=�N*=��)=|�)=/)=/�(=�1(=
�'=�&=E�%=y�$=?#=O�!=�v =[�=�z=}�=�G=ǋ=I�=R�=ٝ=Oo=�4=�=w�	=��=�t=�U=�3=�
�<چ�<���<3��<���<���<^R�<�<��<���<�5�<j��<�m�<�c�<W��<ѷ<�$�<vq�<@��<���<���<�b�<�	�<���<�=�<��<���<�d�<�7�<�|<G�s<P�j<��a<"vX<�O<,�E<a�<<��3<I0+<��"<�g<��<e_	<k <D"�;���;�o�;ϱ;��;R}�;#�h;=B;�b;���:���:��h:��9dxb� ��m�� ��򺦽��n;���]���"𐻊n��5_�����g�ϻPS޻t���j����C���H������8%��B*�V�.��03��]7�s�;���?��ED���H��~M�R�hqV�8uZ���]���`��gc�I?e��f�5{g��h���h�P6i� j�'k���l���n�w�p�s�yu���w��y�
�{���}��f��������߭���ー�,���z��Q����ꈼ� ��K��_������)��9u����ţ������w���w��[j��R;��۝��?��Se��4M����������Y���7f��A裼����e��n��Ϥ������e���̫��$��xe��΍��ģ��統�kӲ����[���Ŷ��=��7���X��%c���  �  ܋O=�O=�yN=��M=�AM=a�L=��K=e�J=��I=l�H=��G=�F=��E=�'E=�{D=h�C=z{C=�!C=��B=՜B=�^B=�B=ټA=LA=��@=�%@=�x?=�>=�>=�d==l�<=�/<=e�;=�;=��:=��9=�b9=��8=�"8=;�7=��6=�w6=x�5=�5=�5=ى4=J�3=�>3=%t2=��1=ߣ0=4�/=j�.=j�-=��,==,=,�+=o	+=m�*=m&*=t�)=�\)=��(=�X(=i�'=��&=��%=��$=^\#=��!=�� =��=�i=��==�U=4v=�{=�h=:D=�=��='�	=آ=ĉ=�q=�S=�N�<��<�<52�<�!�<]��<��<���<�u�<��<	��<�H�<���<��<.�<S>�<���<Ͱ<���<U�<J��<M��<�W�<y�<sm�<���<���<YB�<���<�[{<�r<��i<+�`<A�W<��N<,uE<܎<<��3<�q+<'#<��<��<��	<]� <�Q�;���;���;�e�;�ޞ;䌊;]hm;G;�N";��:8�:E�y:{ :��%8_�չJ,a�Vc���l캇��"�8�t:[�q�}��8��"��:~��EW��Űл�߻^m������Y���u����#����$��)��Y.���2�ؽ6�0�:��3?�"�C�:.H�[�L��?Q�ʃU��lY��\�u�_��?b��!d��e���f��Gg���g���h��bi��j�<l�]�m�O'p�v�r�eu�x�w���y��|��~���_���)���?���@���u������·�P����݉��͊����'���ۍ�[&��ף��ER��`(������
�������J�������ҟ�k���~�����}���-�������>��M��^��pW�������'��������� j��:���D᰼�
���7��s���������-~��ع�*���O���  �  I�O=5!O=˝N=-N=iM=ѭL=�K=��J=��I=I=�H=� G=SGF=�E=��D=�HD=a�C=�mC=�C=g�B=��B=]AB=��A=�sA=��@=�K@=e�?=��>=E!>=�f==;�<=�<=wr;=��:=�I:=M�9=�9=f�8=��7=r7=�6=,�6=�6=9�5=�45=Ӱ4=�4=*f3=7�2=��1=��0=��/=C /=/".=RT-=�,="�+=/b+=��*=�m*= *=�)=R)=�(=d�'=�&=�%=��$=�x#=/"=� =-�=N=��=��=i=�%=�+= ==
�=��=�	=ש=��=ь=�r=W��<��<N]�<t}�<Wx�<�[�<.8�<��<h�<�>�<4��<��<��<@��<g��<��<|��<�.�<�X�<�e�<uL�<��<Ӧ�<�'�<���<��<��<a
�<��<|dz<�q<ڧh<��_<r�V<N�M<��D<�H<<{�3<��+<�#<�`<�<�}
<�<<��;Q6�;�_�;=;�;$�;p�;bs;9$M;Ǒ(;=y;���:�g�:��:���8�p���uT��c����J	���5��X���{������蠻 ر��D»'һ!��_���5���������D!�b����$�?x)��-�~�1��6�H:�	�>���B�_vG�R�K�JP�EeT��&X�;~[� `^�c�`���b��?d�$je�+Of��g�e�g�\�h�%�i��pk��Um�L�o��r�9�t��Zw���y�sc|���~��n��!~������L���5����܅��(�,���Q���1����x��p�������׎�T������:ʓ�ĩ��G����Z����u���𝼜�����࠼񉡼#������<����YǤ��Х��	���k���ꩼlv��� ���|���导�:�������������/L��󕷼%۸�h���5��E���  �  n�O=�5O=ͷN=s)N=υM=��L==�K=%K=�+J=�<I=�RH=�tG=��F=��E=�BE=j�D=_-D=s�C=�^C=
C=$�B='dB=sB=p�A=�A=�g@=}�?=O�>=�(>=�^==��<=��;=!2;=��:=��9=	\9=��8=�B8=5�7=�N7=��6=�6=�#6=ݿ5=�O5=O�4=;44=��3=��2=@�1=�1=&0=�J/=�y.=E�-=�-=,\,=��+=�9+=��*=�<*=��)=�8)=�(=	�'=5'=u	&=��$=��#=p"=� =��=K%=`=}�=ԯ=��=	�=�=�=.�=r�=R�	=j�=T�=�=߆=)��<q;�<��<���<���<���<z��<׺�<���<�
�<ea�<���<�{�<JC�<q/�<v;�<o\�<��<�<l��<p��<�L�<��<vW�<[��<��<4\�<��<�!�<�-y<!(p<\.g<@^<fU<��L<s%D<��;<W�3<v�+<F�#<۱<o<�
<��<�l�;�O�;���;{
�;�R�;�ӏ;R\y;��S;Ǚ/;�V;��:��:�&:��(9FT���gI�Vp�����s��%�3��V��[z��%�����߉����û�Իp�㻻7�� ����|�����������$��8)�Eq-���1�3�5���9��>�UsB���F�s+K��SO��7S�-�V���Y�ż\�'$_�),a�9�b�8d�%Ue��If��4g�8h��ri�q�j�D�l��#o�1�q�Gtt�(Pw�)z���|���.���M#���@���U���a��:a���O���*��_�˳��Nu��`G��g8��7S��ߝ��z������+w��A��n��Ի��tT��b˛����hJ���Q���5������J���K����x���ό��F���Ѧ�7��>���n_����������4��ԯ��G���l����������:.��1T���e���b���M���  �  ��O=�9O=�N=�3N=d�M=c�L=	L=9.K=MJ=�lI=�H=}�G=iG=�SF=v�E=�E=b�D=�D=E�C=�6C=��B=ExB=BB=��A=A=r@=z�?=��>=)!>=�H==2s<=F�;=��:=�2:=��9=n�8=l8=?�7=��7=�7=��6=�u6=a"6=��5=@Y5=��4=�>4=��3=>�2=� 2=�-1=�[0=X�/=�.==.=�k-=X�,=B(,=��+=��*=�r*=_�)=�P)=��(=-�'=	'=x&=�$=��#=�"=cq =�=N�=�=D3=rG=CT=\[=L_=@c=^j=�u=��	=�=��=ћ=��=��<�C�<m��<`��<���<��<�(�<cQ�<���<���<�<�<���<F�<���<D��<ͪ�<�<��<Gͭ<�̩<���<2j�<���<�f�<ޱ�<��<��<�N�<���<�w<�n<$�e<�\<��S<oK<�/C<1);<BN3<��+<��#<;�<*�<��
<�<��;���;L��;Q��;)u�;���;ʲ;#�Z;��6;�X;�M�:ɳ�:G�7:w�_9効&�A�����Yߺ����2�U�U�Z�y��2��?���؟��5GŻ�Tֻ@��g?�����r	����=��\��X �9�$��5)�SQ-�t^1��s5�̞9���=�g+B��mF���J��yN�[R��gU�cX��[�w]�٘_��wa�c�2vd�g�e���f���g�Y@i�4�j� �l���n���q��ut��~w���z���}�?B��4�������_��������!����ȇ��}��1#��Lŉ�$r��?8��W$��>��쇎���������<��딼�����"��_���Q����F��Sw����������[t��)D��9��JĢ������u�����=���%�������f��w&���箼�=���ó�_0��h���ٽ���޸�|幼.Һ�娻��q���  �  �O=+O=%�N=9)N=�M=��L=gL=�3K=�_J=�I=)�H=!H=v_G=ѶF=KF=wE=q�D=aRD=H�C=�VC=J�B=K{B=#B=l�A=�A=�g@=��?=��>=v	>=9%==8@<=#b;=7�:=�9=$9=�8=�8=t�7=�47=N�6=��6=GY6=�6=��5=JN5= �4=�44=O�3=��2=�	2=�E1=B�0=��/=/=�u.=��-=�*-=��,=��+=&>+=��*=��)=GY)=��(=��'=N'=g &=(�$= y#=Q�!=O =�=��=0�=��=��=D�=��=,�==0=�6=�U	=�q=8�=;�=v=[��<i#�<���<���<�<�B�< ��<m��<r4�<���<"�<W��<��<��<F=�<t�<��<�ֱ<�ҭ<�Ʃ<���<p]�<y�<�O�<$��<p��< ��<τ<��<�@v<��l<�c<k�Z<CTR<�J</B<3O:<t�2<�+<wb#<uy<�F<��
<�<��; �;{r�;�ʹ;bH�;@��;?ς;<�a;�=;�;>�:��:�CG:�%�9��{�@�>������]ߺ�����2�	V� ez�Ï��z�����DHǻ��ػk�黙v���#���M�-
�B=�_� ��V%��x)�~-�ւ1��5���9���=�+B��CF��*J�i�M�� Q�(T��V�x|Y�(�[��^�<2`��b���c�Ae���f���g��[i�&�j��l�(o�}�q�E�t���w��7{�-�~��Հ��P������ᄼV�^�������T��[爼�m���������UP���9��S������J��H���� �������.��|���d����=��K{������ڝ�������������ۡ�ݶ��T�����������bѦ�l;���ҩ�ӏ��e���B�����v۲�h�������Z��󎸼,���]����R�����H����  �  8kO=O=�N=N=�iM=�L=��K=1*K=@eJ=r�I=��H=�MH=Q�G=vG=�mF= �E=N*E=�D=��C=1jC=��B=$oB=��A=�wA=7�@=�J@=[�?=3�>=�==��<=�<=�;=^;:=/p9=F�8=�!8=R�7=F97=B�6=��6=�i6=906=��5=��5=h15=a�4=4=�o3=��2=�2=�P1=�0=]�/=�a/=&�.=�'.=͂-=��,=�$,=p+=!�*=�*=�S)=�(=�'=%�&=��%=��$=�U#=�!=i  =tP=�g=�n=ln=l=<m=[u=ֆ=c�=��=��
=B	=�B=�[=�a=R=�V�<x��<�M�<̨�<G �<0_�<���<eC�<��<�F�<���<�6�<���<]�<���<�?�<���<cѱ<嶭<���<#t�<�+�<���<�<�H�<[W�<�P�<
E�<f�~<��t<7k<�b<�3Y<��P<��H<��@<[V9<_�1<'n*<4�"<R�<��<B
<�y<��;C��;���;��;)��;!�;*a�;�`g;��C;��;&��:�:�FS:���9��p�U_?�*�����&��}4��xW�|�GŐ�`ʣ�gȶ��nɻ�oۻ,�����C��=��{���;�=7���!���%�c�)�L�-�Y�1��6��):��S>�MjB��SF���I�RM��YP��S��U�aX��|Z���\��_�9Ga�Bc�%e��f��0h��i��fk�nUm��o�Ar�\Bu��x�� |��}��o��j���r��j����Æ�;����X���舼�_��A͉�uC���ӊ�T���s�����{Ў��4��!���� ��u����啼�,���c��g����Ț�p��A>���x��姟�ZĠ�͡��Ƣ�;��������Υ��
��\u��-��֫�?�����������~���:��4̶�V-��x\���Z��b-��Jݻ�/w������  �  �?O=��N=�pN=3�M=ECM=]�L=Q�K=tK=�`J=��I=I=�|H=~�G=�SG=��F=�F=�dE=��D=�D=�rC=�B=�YB=��A=@SA=V�@=r#@=�k?=p�>=��==*�<=V�;=Y�:=��9=j9=x_8=�7=�F7=��6=8�6=�c6=�36=y6=��5=�r5=�	5=!�4=�3=�M3=��2=8�1=EQ1=�0=b#0=ו/=�/=�n.=N�-=�-=�Y,=*�+=��*=�	*=�D)=�{(=�'=X�&=ô%=�$=Q)#=8�!=��=%=�"==�=�
=�=L=`&=�I=}x=��
=t�=�=�+=�3=�$=���<���<2�<�s�< ��<dg�<��<ϕ�<:7�<B��<tW�<��<�)�<���<�<�d�<���<x��<Ɇ�<_�<r.�<�<�n�<bʗ<`��<���<x߈<���<Q}<2]s<Q�i<7~`<��W<GUO<n`G<��?<�\8<1<<�)<�"<�C<�<��	<�� <
�;K:�;=��;O�;�;
��;8p�;�l;{�H;��$;���:9y�:��[:��9[�p�1�B�8����]废�76��Y�F~����?@��b�����˻��ݻ�:ﻂt��-������c\�m.���"���&���*�X�.��2��6���:��>�G�B���F���I��M�t�O�?FR�@�T�*�V�)[Y���[�2E^�ŭ`���b�� e���f� �h��>j�N�k���m�m8p���r���u�ADy���|��;���������R&���n��+~��:U�������u��@؉��3��)����%��wڋ�����ڍ�h��wt���ב��3��z�������ؖ������X7���s��Z������tg������ӡ��颼������{��aY��.Ĩ�x`���+���������$��F��=嵼/���l鸼`�����3Ȼ�mc��\鼼{m���  �  �O=�N=9IN=ٽM=�M=�lL=ǶK=�K=�WJ=g�I=Y'I=ܝH=|H=��G=��F=�BF=��E=��D=�D= tC=L�B=�BB=��A=�.A=��@=�?=pD?=vt>=ɍ==b�<=�;=y�:=�9=F�8=8=z7=��6=c�6=S_6=�-6=�6= �5=��5=K5=��4=�a4=9�3=�+3=��2=�1=�L1=@�0=5;0=��/=5/=٢.={�-=�F-=S,=ح+=�*=o*=�3)=�_(=��'=z�&=ߊ%=Z$=J�"=�s!=L�=�=+�=��=F�=s�=�=��=��=�=8=t
=��=^�=��=�=�� =:��<�<�<,��<�>�<R��<d�<k�<���<Ј�<C4�<3��<�3�<a��<���<��<�w�<!��<ϖ�<�S�<��<��<���<\#�<w}�<���<W��<�{�<TM�<�P|<[Br<F�h<�I_<X�V<�1N<TF<��><C�7<�J0<��(<�p!<��<q<�<�P <W�;��;�C�;d8�;k�;H��;��;r�o;PLL;��';��;]��:K\a:|��9p}v��G������E麚#��h8�0�[�pG��,=����������?ͻ�߻=^�S� �1O���q��=J�L�=J#�$O'�/7+��!/�+ 3��37��O;�[?��7C���F��J���L��dO��Q�{�S��&V���X��[���]�G`���b��e��g�`�h���j��l�.�n��p��}s���v�g�y�9�}������y���.��O������K��t∼�|��뉼*@���������u��I)������'���c��#���M��9N��������r���r���I���A͙����Qg���ѝ��=��Q���⡼���-���D���g�������ɯ���}��'t��X���0������Kn��Z���}��"���%����F��+Լ�4M��ǽ��  �  ��N=ɞN=:,N=�M=M=tSL=-�K=�J=�OJ=9�I=�1I=�H=�/H=��G=�G=�`F=��E=�D=(D=�rC=H�B=�1B=ݡA=�A=��@=6�?=k'?=AW>=�o==~v<=Ft;=t:=�9=!�8=��7=�J7=��6=�v6=H76=x	6=��5=J�5=�}5=�-5=��4=TE4=�3=�3=�r2=��1=AG1=�0=mH0=J�/='Q/=D�.=.=Nc-=��,=��+=R�*=_ *=
&)=�K(=yj'=y&=�l%=�;$=��"=�S!=�=S�=�=��=��=�=�=�=ƨ=��=�=�M
=L�=9�=��=C�=�� =qk�<;�<���<��<B��<�]�<��<A��<ǹ�<�p�<�<�t�<>��<��<�2�<�~�<Q�<P|�<�,�<{�<a��<\a�<��<"D�<�i�<�`�<}7�<`�<ը{<��q<��g<��^<��U<wM<�E<J1><�6<��/<
{(<{� <� <��<։<���;(l�;��;��;�H�;Oʪ;	e�;mԉ;�q;3�N;�*;8�;���:�Sd:��9&�|���J��&���+����:�9�]��"��J ��񌧻	��jλ��G�򻞒��		�t��_����\��R�#���'�ܩ+��/�$�3�Q�7��;�t�?�O�C�w�F�9J���L�W.O��XQ��tS���U��X�[�Z�dP]�j`�ѯb��e��Ng� Ii�f#k�y�l���n��Iq� �s�& w�bjz�P~��0ɂ�U���E��ma���o��T=��eщ��8��y����Њ�.��I���Wc��TJ��;`������U␼+���c�����ߊ���~���o���o�����zΚ�91��˩��'�������|.��5W��
w�����o᧼�L��ꪼ+���g����Ű�q޲��崼�ƶ��q���ܹ����*껼���8��V�������  �  )�N=V�N=�!N=��M=��L=JL=B�K=[�J=}LJ="�I=�4I=J�H=�8H=�G=�G=�jF=�E=��D=�*D=rC=��B=q+B=��A=6A=Ew@=��?=?=�L>=e==$k<=h;=�f:=�r9=��8=��7=*:7=��6=�g6=i)6=��5=��5=O�5=�r5=�#5=B�4=�:4=�3=�
3=�k2=��1=E1=�0=�L0=j�/=yZ/=��.=�(.=�l-=�,=�+=q�*=F�)=!)=;D(=9a'=�n&=�a%=�0$=��"=�H!=N�=Ͱ=��=��=��=	{=�s=�|=�=�=z�=�@
=>=ܲ=��=��=� =yV�<���<m|�<�
�<-��<�[�<�#�<��<:��<"��<M�<5��<���<��<|:�<��<4�<�q�<h�<ݨ<��<WL�<�՛<�.�<�S�<�I�<��<[�<�m{<�Kq<��g<E?^< yU<�6M<�jE<�=<��6<̖/<mO(<G� <��<��<Gb<���;�0�;���;��;�M�;P�;1��;5"�;�br;>>O;��*;B;l�:{.e:��9$����K�l���P�"Y���:��&^��u��[v���移�|��_�λ��Ỏ=����sK	������Y��S�#���'�K�+�ѻ/���3��7��;���?�ڡC��G�c J�g�L�O��;Q�OS��|U���W��sZ�o2]��_�U�b��$e�"ag�0ei��Fk��%m�@)o��rq�|t�=*w��z��D~�����䂼&���1��4��������\����S������犼�C��>ŋ��w��_���t�����L�8��l��K�������Pt���_��\��xw������A������ ��	������V9���f������@���(����a������xά��Ȯ��ݰ�L�����A嶼摸�t���2$���������X9��B���/���  �  ��N=ɞN=:,N=�M=M=tSL=-�K=�J=�OJ=9�I=�1I=�H=�/H=��G=�G=�`F=��E=�D=(D=�rC=H�B=�1B=ݡA=�A=��@=6�?=k'?=AW>=�o==~v<=Ft;=t:=�9=!�8=��7=�J7=��6=�v6=H76=x	6=��5=J�5=�}5=�-5=��4=TE4=�3=�3=�r2=��1=AG1=�0=mH0=I�/=&Q/=C�.=.=Mc-=��,=��+=Q�*=^ *=
&)=�K(={j'=y&=�l%=�;$=�"=T!=;�=��=[�=�=�=u�=��=��=��=��=�=�N
=��=��=D�=��=D� =�n�<;�<q��<��<���<�_�<F!�<���<���<Wq�<0�<=t�<~��<���<51�<
}�<�<�y�<�)�<��<k��<b^�<�<VA�<�f�<^^�<n5�<���<0�{<��q<��g<��^<W�U<�xM<��E<�4><'�6<��/<J�(<$� <�&<��<�<���;lw�;F%�;�;�P�;�Ъ;j�;�׉;�q;�N;�*;��;ɂ�:d:�_�9~:~���J��V���^�B���+:�Ğ]�w/���,�������%��tλ��3�����	����}�����̐�|�#���'���+���/���3���7�_�;���?�{�C���F�TJ���L�g.O��XQ��tS���U��X�_�Z�gP]�l`�ӯb��e��Ng� Ii�g#k�y�l���n��Iq��s�& w�bjz�P~��0ɂ�U���E��ma���o��T=��eщ��8��y����Њ�.��I���Wc��TJ��;`������U␼+���c�����ߊ���~���o���o�����zΚ�91��˩��'�������|.��5W��
w�����o᧼�L��ꪼ+���g����Ű�q޲��崼�ƶ��q���ܹ����*껼���8��V�������  �  �O=�N=9IN=ٽM=�M=�lL=ǶK=�K=�WJ=g�I=Y'I=ܝH=|H=��G=��F=�BF=��E=��D=�D= tC=L�B=�BB=��A=�.A=��@=�?=pD?=vt>=ɍ==b�<=�;=y�:=�9=F�8=8=z7=��6=c�6=S_6=�-6=�6= �5=��5=K5=��4=�a4=9�3=�+3=��2=�1=�L1=?�0=4;0=��/=5/=ע.=x�-=�F-=P,=խ+=��*=m*=�3)=�_(=��'=��&=�%=�Z$=j�"=t!=��=_�=��=B�=�=k�=4�=0�=o�=k=%:=]v
=4�=�=�=�
=�� =/��<�B�<���<�C�<���<h�<��<���<���<S5�<m��<N3�<��<���<��<�s�<��<���<>N�<#�<A�<���<��<x�<y��<Ț�<�w�<J�<�K|<�>r<r�h<{I_<��V<O5N<YF<�><$�7<�S0<�)<�{!<�<�|<�	</\ </�;��;�U�;H�;�w�;ř;1�;��o;pKL;��';1�;sϺ:J�`:'��9��x�L�G���;�麎V�^�8�y\�w`��.U�������#���Rͻ^�߻�m�� ��T��
����M��}L#��P'��8+��"/�!3�\47�hP;��[?�8C���F��J���L��dO��Q���S��&V�ȇX��[���]�G`� �b��e��g�a�h���j��l�/�n��p��}s���v�g�y�9�}������y���.��O������K��t∼�|��뉼*@���������u��I)������'���c��#���M��9N��������r���r���I���A͙����Qg���ѝ��=��Q���⡼���-���D���g�������ɯ���}��'t��X���0������Kn��Z���}��"���%����F��+Լ�4M��ǽ��  �  �?O=��N=�pN=3�M=ECM=]�L=Q�K=tK=�`J=��I=I=�|H=~�G=�SG=��F=�F=�dE=��D=�D=�rC=�B=�YB=��A=@SA=V�@=r#@=�k?=p�>=��==*�<=V�;=Y�:=��9=j9=x_8=�7=�F7=��6=8�6=�c6=�36=y6=��5=�r5=�	5= �4=�3=�M3=��2=6�1=DQ1=ߵ0=`#0=Օ/=�/=�n.=J�-=�-=�Y,=&�+=��*=�	*=�D)=�{(=�'=b�&=ִ%=2�$=)#={�!=�=�=@#=�=�==l	=J=�(=�L={=��
=�=�=0=/8=�(=g�<���<�<{�<���<$m�<���<���<�9�<���<�W�<2��<�'�<���<��<�_�<���<���<X�<2W�<Z&�<�ڠ<�f�<�<@�<X�<�و<��<�I}<>Xs<��i<~`<��W<�YO<lgG<�?<�g8<�1<��)<?,"<�S<|(<��	<�� <�(�;�V�;ڞ�;p�;ѩ;۩�;dy�;]$l;>�H;�|$;���:z<�:}>[:!g�9�#t�?�C�S���庵J��6���Y��~��'��A`�����ۜ˻1�ݻ�P�e����5�������0a�\2��"�<�&�Ǜ*���.�:�2��6�b�:���>���B�S�F���I��M���O�`FR�Z�T�>�V�8[Y���[�;E^�̭`���b�� e���f��h��>j�P�k���m�n8p���r���u�ADy���|��;���������R&���n��+~��:U�������u��@؉��3��)����%��wڋ�����ڍ�h��wt���ב��3��z�������ؖ������X7���s��Z������tg������ӡ��颼������{��aY��.Ĩ�x`���+���������$��F��=嵼/���l鸼`�����3Ȼ�mc��\鼼{m���  �  8kO=O=�N=N=�iM=�L=��K=1*K=@eJ=r�I=��H=�MH=Q�G=vG=�mF= �E=N*E=�D=��C=1jC=��B=$oB=��A=�wA=7�@=�J@=[�?=3�>=�==��<=�<=�;=^;:=/p9=F�8=�!8=R�7=F97=B�6=��6=�i6=906=��5=��5=g15=a�4=4=�o3=��2=�2=�P1=�0=[�/=�a/=#�.=�'.=ɂ-=��,=�$,=p+=�*=�*=�S)=�(=�'=2�&=��%=��$=�U#=Z�!=�  =Q=�h=�o=�o=�m=Fo=�w=��=��=��=��
=�!	=�G=�`=g=CW=La�<���<*W�<���<V�<<f�<���<H�<H��<�H�<,��<�5�<��<t�<W��<d9�<��<�ȱ<ƭ�<擩<9j�<�!�<쮜<��<@�<xO�<�I�<V?�<��~<��t<�3k<wb<�6Y<��P<��H<��@<�c9<�1<�*<�"</<��<fV
<��<�!�;@��; ��;$��;oͨ;�;jl�;1kg;/�C;�;�`�:��:Q�R:ˑ9Uu���@�2��T�xS��x4���W��\|���񣻿춻��ɻ��ۻ���
���8���������A�<�q�!���%���)�K�-���1��6��*:�YT>��jB�oTF�A�I�GRM��YP��S� �U�yX��|Z���\��_�BGa�Bc�*e���f��0h��i��fk�oUm��o�Ar�\Bu��x�� |��}��o��j���r��j����Æ�;����X���舼�_��A͉�uC���ӊ�T���s�����{Ў��4��!���� ��u����啼�,���c��g����Ț�p��A>���x��姟�ZĠ�͡��Ƣ�;��������Υ��
��\u��-��֫�?�����������~���:��4̶�V-��x\���Z��b-��Jݻ�/w������  �  �O=+O=%�N=9)N=�M=��L=gL=�3K=�_J=�I=)�H=!H=v_G=ѶF=KF=wE=q�D=aRD=H�C=�VC=J�B=K{B=#B=l�A=�A=�g@=��?=��>=v	>=9%==8@<=#b;=7�:=�9=$9=�8=�8=t�7=�47=N�6=��6=FY6=�6=��5=IN5= �4=�44=N�3=��2=�	2=�E1=@�0=��/=	/=�u.=��-=�*-=�,=��+=!>+=��*=�)=EY)=��(=��'=]'=� &=R�$=@y#=��!=�O =��=p�=`�=]�=��=��=��=Y�=�=K=~;=�Z	=w=É=�=�{=ި�<�.�<���<���<�<kJ�<���<���<8�<���<��<$��< �<���<q7�<G��<fڵ<�ͱ<xȭ<<���<RR�<��<WE�<k��<���<Y��<�Ȅ<��<�9v<�l<��c<��Z<�ZR<J<�B<^^:< �2<)+<�w#<��<9]<H�
<)<��;G�;���;�;Ca�;,�;�ۂ;�a;>�=;��;��:�S�:�lF:��9PW��T�?�F����� ��'3�lV���z�Y�&���)<��?mǻ�ػ��^����.��
��U����B��� �WZ%��{)�I�-���1���5���9�Z�=��+B�qDF�+J���M�� Q�K(T�%�V��|Y�=�[��^�I2`��b���c� Ae���f���g��[i�(�j��l�(o�~�q�F�t���w��7{�.�~��Հ��P������ᄼV�^�������T��[爼�m���������UP���9��S������J��H���� �������.��|���d����=��K{������ڝ�������������ۡ�ݶ��T�����������bѦ�l;���ҩ�ӏ��e���B�����v۲�h�������Z��󎸼,���]����R�����H����  �  ��O=�9O=�N=�3N=d�M=c�L=	L=9.K=MJ=�lI=�H=}�G=iG=�SF=v�E=�E=b�D=�D=E�C=�6C=��B=ExB=BB=��A=A=r@=z�?=��>=)!>=�H==2s<=F�;=��:=�2:=��9=n�8=l8=?�7=��7=�7=��6=�u6=a"6=��5=@Y5=��4=�>4=��3=<�2=� 2=�-1=�[0=V�/=�.=9.=�k-=T�,==(,=�+=��*=�r*=[�)=�P)=��(=4�'='=�&=G�$=ċ#="=�q =Ѻ=A�=�=�4=bI=�V=+^=�b=g=�n=vz=�	=~�=i�=��=��=��</O�<���<���<���<�<�/�<�V�<W��<���<�<�<���<*C�<��<8��<[��<B��<U��<�­<e��<��<�^�<��<�[�<Ч�<n��<��<�G�<䊀<�w<e�n<�e<L�\<+�S<�xK<�<C<�8;<f`3<��+<|�#<%�<��<<�/<���;<"�;���;���;���;/��;��;q�Z;��6;�H;7�:�]�:+7:�[9�R��b9C�G>��������2��"V�F1z��b��a����ɳ�smŻ&wֻ���Z������|	������b�.] ���$��8)��S-�G`1�u5��9�l�=�,B�wnF��J�zN��R��gU�0cX�[�#w]��_��wa�'c�9vd�l�e���f���g�\@i�6�j��l���n���q��ut��~w���z� �}�?B��5�������_��������!����ȇ��}��1#��Lŉ�$r��?8��W$��>��쇎���������<��딼�����"��_���Q����F��Sw����������[t��)D��9��JĢ������u�����=���%�������f��w&���箼�=���ó�_0��h���ٽ���޸�|幼.Һ�娻��q���  �  n�O=�5O=ͷN=s)N=υM=��L==�K=%K=�+J=�<I=�RH=�tG=��F=��E=�BE=j�D=_-D=s�C=�^C=
C=$�B='dB=sB=p�A=�A=�g@=}�?=O�>=�(>=�^==��<=��;=!2;=��:=��9=	\9=��8=�B8=4�7=�N7=��6=�6=�#6=ݿ5=�O5=N�4=:44=��3=��2=?�1=�1=}&0=�J/=�y.=B�-=�-='\,=��+=�9+=��*=�<*=��)=�8)=	�(=�'=C'=�	&=��$=�#=�"=�� =��=6&=Ba=��=��=��=��=:�=��=F�=��=@�	=��=ݪ=��=��=���<�F�<���<���<���<���<��<��<Y��<��<�a�<���<#y�<�>�<�)�<B4�<
T�<�z�<���<���<_��<�A�<�ל<M�<���<���<�T�<ò�<��<�&y<�$p<&.g<%C^<nlU<�L<�1D<�;<��3<��+<S�#<��<ą<��
<�<Ֆ�;w�;���;�(�;�k�;��;�uy;�T;�/;�G;�E�:�X�:�0%:��$9ƭ����J�\%��ѝ� ��4��W�F�z�#T��r-��E����û�.Ի�
�yQ� �L�l��|��z��|����$�h;)��s-�Y�1���5���9��>��sB�U�F��+K�TO��7S�[�V���Y��\�<$_�9,a�E�b�"8d�,Ue��If��4g�8h��ri�s�j�E�l��#o�2�q�Gtt�(Pw�)z���|���.���M#���@���U���a��:a���O���*��_�˳��Nu��`G��g8��7S��ߝ��z������+w��A��n��Ի��tT��b˛����hJ���Q���5������J���K����x���ό��F���Ѧ�7��>���n_����������4��ԯ��G���l����������:.��1T���e���b���M���  �  I�O=5!O=˝N=-N=iM=ѭL=�K=��J=��I=I=�H=� G=SGF=�E=��D=�HD=a�C=�mC=�C=g�B=��B=]AB=��A=�sA=��@=�K@=e�?=��>=E!>=�f==;�<=�<=wr;=��:=�I:=M�9=�9=f�8=��7=r7=�6=,�6=�6=9�5=�45=Ұ4=�4=)f3=6�2=��1=�0=��/=@ /=,".=OT-=�,=�+=+b+=��*=�m*= *=��)=P)=�(=j�'='�&=%�%=!�$=�x#=�"=�� =��=�N=��=5�==�'=7.=�"=S=��=��=N�	=��=��=�=x=���<�<�f�<d��<p��<�b�<>�<*#�<� �<�@�<���<��<[��<Q��<%��<���<��<�&�<�O�<�[�<�B�<��<��<J�<呓<��<3~�<��<���<x^z<�q<��h<Z�_<!�V<��M<�D<kV<<&�3<�+<�#<~t<Q&<�
<��<��;qY�;F�;�V�;�#�;~'�;	-s;�.M;?�(;rk;��:��:�#:5��8����C�U����8:级a�D6��Y�<|�䵏����.���f»�Dһ���q��I��d��֙��� &�V����$��z)�"�-� 2��6�I:�ˑ>�@�B��vG���K�RJP�{eT��&X�[~[�`^�v�`���b�@d�,je�1Of��g�i�g�_�h�(�i��pk��Um�L�o��r�9�t��Zw���y�sc|���~��n��"~������L���5����܅��(�,���Q���1����x��p�������׎�T������:ʓ�ĩ��G����Z����u���𝼜�����࠼񉡼#������<����YǤ��Х��	���k���ꩼlv��� ���|���导�:�������������/L��󕷼%۸�h���5��E���  �  ܋O=�O=�yN=��M=�AM=a�L=��K=e�J=��I=l�H=��G=�F=��E=�'E=�{D=h�C=z{C=�!C=��B=՜B=�^B=�B=ټA=LA=��@=�%@=�x?=�>=�>=�d==l�<=�/<=e�;=�;=��:=��9=�b9=��8=�"8=:�7=��6=�w6=w�5=�5=�5=ى4=I�3=�>3=$t2=��1=ޣ0=3�/=h�.=h�-=��,==,=(�+=k	+=i�*=i&*=p�)=�\)=��(=�X(=n�'=��&=��%=��$=�\#=
�!=� =w�=�j=��=(=�V=�w=�}=k=�F=�=��=��	=��=Ѝ=#v=X=NW�<Q��<��<�9�<n(�<'��<���<c��<�x�<v��<[��<�G�<���<T�<���<
9�<k��<ư<q��<t�<0�<+��<�O�<�ݗ<\f�<N��<���<�=�<Z�<�V{<]�r<��i<n�`<�W<��N<?~E<�<<��3<�+<n6#<��<.�<� 
<�<�p�;x��;���;M|�;#�;ך�;�zm;�G;tM";V��:��:�by:��9Ŧ8�@׹�!b��筺��캪6�9�ʂ[��?~��Z���:������<r���л��߻3��	��Ѻ�+���z����^��6�$��)��[.��2�ݾ6���:�Y4?���C��.H���L�5@Q���U�mY�.�\���_��?b��!d�
�e�Ƌf��Gg���g���h��bi��j�>l�^�m�P'p�v�r�eu�y�w���y��|��~���_���)���@���@���u������·�P����݉��͊����'���ۍ�[&��ף��ER��`(������
�������J�������ҟ�k���~�����}���-�������>��M��^��pW�������'��������� j��:���D᰼�
���7��s���������-~��ع�*���O���  �  �vO=��N=&VN=��M=kM=�^L=׊K=�J=��I=,�H=?�G=n�F=^�E=��D=�1D=��C=?7C=��B=V�B=�kB=�2B=��A=:�A=�$A=@�@=��?=�U?=ۧ>=��==�]==��<=�E<=e�;=I;=[�:=�2:=Г9=��8=�>8=��7=��6=j6=�5=�h5=��4=�b4=��3=I3=
L2=Yi1=ju0=y/=�~.=��-=Y�,=��+=�M+=��*=�N*=��)=z�)=/)=.�(=�1(=�'=�&=S�%=��$='?#=�!=4w =��=R{=�=xH=��=v�=��=|�=/q=7=e�=�	=[�=�w=�X=�6=��<���<��<^��<k��<���<�U�<��<���<���<�5�<ɱ�<zl�<�a�<L��<Gͷ<] �<�l�<���<g��<͙�<�\�<Q�<E��<�8�<ߎ<���<oa�<L5�</	|<x�s<4�j<2�a<iyX<�#O<��E</�<<��3<Y:+<~�"<'s<W
<"k	<�v <'8�;ϳ�;���;�ޱ;��;2��;B�h;5CB;�a;���:�ײ:wh:"8�9�+��U𹳸m��~���}����;���]����������t��'�����ϻ�b޻���Av�����`#�������:%��C*���.��13�h^7��;��?�FD���H�M�>R��qV�PuZ���]��`��gc�R?e��f�9{g�h���h�R6i�!j�'k���l���n�x�p�s�yu���w��y�
�{���}��f��������߭���ー�,���z��Q����ꈼ� ��K��_������)��9u����ţ������w���w��[j��R;��۝��?��Se��4M����������Y���7f��A裼����e��n��Ϥ������e���̫��$��xe��΍��ģ��統�kӲ����[���Ŷ��=��7���X��%c���  �  �fO=��N=�<N=%�M=��L=�AL=�mK= �J=�I=�uH=�jG=jF=�~E=ԯD=�D=lvC=4C=1�B=g~B=VJB=�B=6�A=xA=�A=�@=�?=�<?=�>=2�==HW==��<=`Q<=��;=�d;=��:=�R:=T�9=�9=bN8=@�7=�6=�^6=��5=�Q5=P�4=�F4=�3=K�2=�.2=/K1=/U0=�U/=�W.=xe-=��,=��+=�+=@�*=4$*=��)=gl)==)=��(=�(=Kf'=��&=��%=�j$=�)#=�!=�m =��=ԃ="�=�b=7�=��=��=�=(�=SG=0=��	=��=Af=�B=�=��<�V�<H��<5��<��<�[�<��<���<��<��<(��<vQ�<��<�
�<�7�<Ʉ�<�ݳ<�-�<�c�<�t�<�]�<#�<+ϛ<�p�<��<|̎<n��<�t�<V[�<�t|<t<Fk<�9b<L�X<wxO<�	F<�<<z�3<X+<�|"<G<8�<��<� <5P�;���;���;İ;�ߛ;^,�;��e;*?;;:;���:Q�:�t]:&�9*�T��� ���u��}��.p��*��={=���_� ΀�����ġ�|i���|��� ϻ|�ݻ����z��6������\��y���j%�f�*�F@/�6�3���7��<�#K@��D�VUI��N���R��W�� [���^��a��%d��e�h?g�*h�+�h�\#i��i��yj�Y�k��m�P o��'q�us���u���w�4�y��{�?o}�+
��^���T���n��쫃� ���`��t���c���i���,��u2��l>���b�����(-���ޒ�P����������ֺ�������7������à�+���qR���Ң��<������$��ɤ�$���˧���ܧ��0������E�7���f��]|��.����������pȳ����ˑ��U���������nt���  �  �wO=��N=;N=j�M=��L=�'L=6XK=�xJ=��I=��H=��G=�F=<�E=�*E=�D=��C=�qC=�	C=�B=�]B=B=~�A=:KA='�@=�N@=t�?=s?=Jz>=k�==�===�<=�<=�;=J;=Pv:=��9=�A9=G�8=��7=kR7=/�6=�6=��5=��4=�e4=L�3=�#3=rk2=R�1=#�0=,�/=��.=m.=+)-=;T,=�+=b�*=^D*=D�)==4)=t�(=�/(=��'=�&=�2&=HP%=�M$=�,#=��!=�� =r:=��=BD=ұ=�=�Q=~=]�=ˍ=lx=�W=j1=�
	=��=8�=,�=6| =���<��<�q�<���<���< ��<e��<w��<C��<��<$^�<��<���<��<�<���<�<��<F0�<]8�<�%�<S��<J��<�p�<�#�<�ڎ<.��<U`�<�(�<��{<Es<ŋj<Ψa<��X<&�O<�F<O�=<�4<�	,<�u#<s�<�Q<��	<�� <ک�;,��;;"�;_�;`��;{�;�3s;��M;�);�;���:o-�:\:��9d��!�K�!颺�u�p��EV1��GR��8s��艻3登z���9���6�ǻ5.ֻN�仦��s �/X�W��^��\�?��L(%��*�=�.��3��7�b�;��c@���D��UI�	�M�m�Q��U�=&Y�g-\��^���`���b�R�c�e�� f�0g��_h�m�i�<ik��Lm�/co�Z�q�<�s�#v�?x�eLz��F|��;~�����*���I���z��H�������64���f��ꍉ�����nʋ����-��1���X��ա���\���)���������Xl��D���`Q���}���{��6Q��v��$����P��+����ä���������ا�t���d�����������:��!l��ٔ�����벼)���w���ն�;��x�������O���  �  OzO=l�N=�?N=ɛM=y�L=�-L=�^K=�J=9�I=��H=O�G=+�F="�E=P6E=�D="�C=Q|C=�C=2�B=�eB=mB=B�A=�QA=3�@={T@=��?=!?=�}>=V�==�===�<=�<=V�;=�:=3n:=��9=�99=ږ8=7�7=�O7=u�6=�6=ъ5=�4=�j4=��3=�)3=�q2=ۧ1=6�0=��/=O�.=�.=�3-=W_,=��+=��*={O*=��)=�=)=�(=n7(=}�'=P�&=�8&=�U%=�R$="1#=n�!=� =;=_�=�@=F�=?=�H=�t=�=�=q=�Q=�-=a		=2�=�=.�=� =���<2�<5|�<��<���<���<O��<s��<��<M�<tu�<� �<���<؟�<]��<Uɷ<K��<�!�<R?�<�F�<�3�<�<�ƛ<�y�<�)�<eݎ<t��<-Z�<��<@�{<@$s<Thj<D�a<ӅX<yO<�qF<�=<˶4<|,<S�#<��<�b<*�	<�� <z��;���;�[�;d��;�֠;�5�;O�s;�|N;k*;1�;)Q�:C��:W�:�t9&����oI�����I���0���Q��r�Љ�{ݙ�����Ѹ���ǻFbֻ+�仓�x� �p����h�*^�D���%�$�)���.��3�uk7��;��H@�!�D�O6I��M���Q�D�U�a�X�e�[��^���`�
db�w�c���d�� f�Ng�(Eh���i�XQk�:6m�6Oo�C�q�)�s��v�Ax��Vz��X|��T~��,��#;��.Z��R���Ä� ���8��g��p�����������a猼X"��&{������l���ON��t��藼ԫ��W���ޜ�i:��g���e���<������"���4A��>𣼦�������夦�'ͧ����]������0���c=���r�����nʱ�y����9��̇���㶼�E��n���� ���M���  �  S�O=i�N=�LN=��M=��L=�>L=�pK=�J=u�I=��H=��G=w�F=�F=�WE=��D=5D=��C=�0C=�B=�|B=0'B=-�A=LcA=��@=Ud@=�?=H-?=��>=W�==�===��<=�
<=�x;=T�:=�U:=�9=�"9=b�8=��7=�F7=��6=�6=;�5=%5=1x4=�3=�93=ւ2=(�1=�0=��/=�/=a0.=�Q-=�,=ֽ+=+=�o*=��)=%Y)=u�(=
M(=η'=�'=I&=e%=�`$=^=#=�!=�� =T<=�=06=��=i�=/=�X=7l=�k=�[=�A=�#=>	=Y�=��=�=9� =s��<i;�<֚�<���<W��<���<z��<�<�!�<�Z�<��<2E�<���<�ݿ<��<��<A%�<�L�<�g�<�l�<�W�<q(�<��<��<�8�<�<�<�E�<Q��<Lg{<�r<��i<�a<*X<�.O<x=F<Yf=<B�4<�,<̞#<"$<��<{�	<�� <u^�;3f�;=�;&_�;ǯ�;�(�;��u;j�P;��,;t

;���:K��:�&:��59�敹f�C��N��:޺H���/��P�A3r�F���4Ι�ݫ��Z$��k=Ȼ�׻ˈ����� �m��QJ�a��f�-����$�r�)�@W.���2�$(7�Z�;���?�mrD�6�H�})M��?Q�U�OwX��x[�!	^��*`��a��Wc���d�ӧe���f�#�g��ei�sk�r�l�o��\q���s��v�=Ix��vz�a�|���~�AZ��yl���������焼S���E���h��~���q��������ʌ�����Y���Ӑ��n��>%���땼鴗��r��5��˜�����R$��&�����鿡�!m��>��Yɣ�y���nz������<�����PH����������oE����������:󱼰*��gk��}���L��Vf��Լ��(
���K���  �  �O=P�N=�]N=ҾM=�M=zVL=�K=خJ=��I=G�H=0�G=�G=�IF=>�E=%�D=cLD=��C=�\C=[�B=g�B=�EB=V�A=3|A=,A=z@=��?=�=?=��>=��==�:==^�<=�;=�[;=��:=a.:=��9=�8=5c8=.�7=I77=�6=o 6=8�5=�5=��4=��3=P3=�2=$�1=��0=f0=�;/=0Z.=�-=P�,=��+=�A+=��*=*=��)=C�(=m(=��'=�&'=�_&=�y%=�s$=�M#=`
"=�� =�;=��=�#=�=��=&=�+=l?=TB=�8='=�=u�=��=��=��=c� =���<@b�<���<��<�+�<�=�<PJ�<�\�<��<��<~$�<���<gc�<�=�<\8�<�J�<uj�<Պ�<���<ա�<]��<V�<>�<G��<J�<g�<��<�!�<�ǁ<6�z<�r<�Si<�x`<d�W<�N<k�E<<1=<�4<�),<��#<]<��<>,
<S?<Q�;o>�;F��;��;���;���;�1y;�T;�)0;�};�'�:��:8	2:�p]9�+����;�ؗ��{�ںN{��[.�ŶO��@q�FS���͙�F�������;ɻ�ػ��k��hz�6����M��d|������$���)��	.��n2��6�\+;�{�?��C�YH�m�L���P��OT�C�W�V�Z�^7]�a_��-a���b��c�D#e��Mf���g��i�j�j�ףl���n�c q���s�2�u��_x�h�z���|�m�Ȥ��Ӽ���ڂ������"���D��/_��p���x��S~��k�������׍��+��#���*9��3铼����og����������6��E�������Kß�h���n���$���֢����\_���J��X��>���?Ш�^-��q��������V�����J�c6���w��6���\���Q��霸�,⹼[��|M���  �  �O=��N=gnN=��M=;)M=HoL=^�K=�J=��I=�
I=�*H=�RG=~�F=��E=�#E=�D=WD=@�C=@*C=��B=�hB=�B=��A=�A=%�@=(�?=LM?=y�>=��==3==��<=��;=�3;=F�:=��9=/`9=��8=�68=J�7=}7=y�6=86=͡5=�"5=j�4=�	4=�g3=c�2=��1=Y1=�E0=�h/=��.=��-=�,=63,=��+=��*=H*=p�)=�&)=��(=|�'=�A'=\w&=�%=4�$=�\#=�"=� =)6=��==�X=t�=��=@�=8=�
=�=A=q�
=�=��=�=��=� =J��<k��<���<O;�<�j�<R��<r��<���<���<�B�<���<\6�<v��<���<��<q��<c��<�Ѱ<M߬<�ڨ<p��<r��<�1�<�ʗ<jV�< ܎<b�<�<�z�<"z<rCq<�lh<�_<��V<�	N<3dE<��<<�v4<k',<�#<Ǐ<�<m{
<��<���;�1�;!�;�۷;���;t�;�@};�nX;��4;��;�p�:�;�:��?:]{�9��^��2�)}����ֺ�����,�tN��_p��$����,q��z���Dʻg�ٻT�#����@����F-���J��^��3�$�	O)�>�-��2��i6���:�h?��wC���G���K�T�O��eS�y�V�|�Y�.\�b^�B`�f�a�!@c��d���e��g��h��Uj��Nl�ǃn��p��ms���u��x�{��u}�����	��j)��PF��[`���u��=���)�������v��@l��|k�� ~��/�������5m������s����V��$	�� ����A��A����	���9���F���4���	��6Ρ�����Q���'�����X*���]��X������ȉ������t���ޯ��=������y೼^)���n������^鸼;���=���X���  �  5�O=�O=yN=a�M=u:M=$�L=ҼK=��J=�J=�6I=�_H==�G=9�F=�F=nE=��D=�KD=�C=A]C=��B=��B=�B=��A=�.A=֠@=�@=�V?=�>=��==�#==jg<=��;=� ;=�X:=��9=N9=��8=��7=�{7=��6=��6=�6=ʡ5=�)5=��4=\4=�y3=;�2={	2=�=1=�k0=M�/=e�.=��-=E6-=�|,=/�+=�&+=-�*=Y�)=wU)=g�(=((=LY'=(�&=z�%=��$=�e#=."=_� =�(=�=��=4'=�]=�=d�=��=��=��=�=y�
=[�=��=��=��=v� =��<!��<��<i�<\��<���<��<�:�<s}�<$��<IC�<���<�t�<;8�<e�<A
�<��<o�<H�<�
�<|�<d��<�M�<Rڗ<~U�<6Ǝ<�3�<���<��<J.y<�9p<;Vg<a�^<��U<�4M<ƼD<g<<�.4<O,<T�#<��<�I<
�
<��<��;��;�<�;�D�;<M�;y�;7�;M];q�9;>�;���:5��:%N:�/�9x�5�=*��Γ�t�Ӻ�T
�Ɯ+�S�M�G�o��(��cK���.��{�����˻kMۻ�H�c���%2�x�	���������?��M�$�-)�s�-��1�X6�j:��>���B��!G��K�V�N�lcR�ݔU�MuX�E[��D]�@=_���`��b���c�DJe�G�f��Gh�ej�Jl�:Qn���p�@js�/ v� �x�߈{��"~��Q��o���֬���ȃ��؄�݅��Ԇ�W����������g��pY��9c��]����Վ��@��ȑ�Fb�����!���6:��M���5&���t������+���緟�����=t��D��������j�\���?������&
��v���������\%������Y��q_��m����A#���I���b���n��r���  �  B|O=5 O=zN=��M=�AM=��L=��K=B K=�/J=X_I=�H=��G=JG='aF=�E= E=�D=�
D=7�C=�C=¦B=�3B=]�A=l8A=��@=�@=�V?=�>=��==�==�C<=��;=!�:=E:=Co9=}�8=4E8=��7=�F7=��6=�j6=�6=��5=�'5=��4=�4=��3=��2=J2=-V1=�0=$�/=�.=�9.=~-=��,=,=�n+=��*=R%*=Y�)=o�(={((=�h'=Ó&=��%=�$=<d#=�"=� =~=Hm=д=�=�=�:=-U=�i=�z=��=M�=��
=��=m�=<�=>�=�� =�<4��<'�<)��<9��<Y�<�a�<���<Z�<�i�<���<�i�<�<���<J��<�e�<�S�<J�<�>�<�(�<���<z��<�U�</ח<-B�<���<$�<�J�<���<� x<o<�f<1U]<B�T<>L<j�C<��;<�3<��+<н#<�<�L<��
<� <,	�;r��;U2�;%��;��;��;�7�;�Ub;p�>;"�;= �:���:�Q\:!*�9���86#�)���{Ѻ9�	�k�*��.M�J�o��s���ꚻ�.����=�ͻTݻ-{�=���)C�ݩ
�>���4��a�)9 ���$�x0)��y-��1���5��6:�~o>��B�ŘF�mJ�TN��^Q�arT��BW���Y�q \��5^��`��a��^c���d��pf�Kh���i�%�k��Fn���p�k�s�;dv��Hy�d'|���~��̀����
@���Z��ya���T��o6��A
���Ո�k���Bt���Z��N\���~��Î�\&��⡑��+�������E��^ŗ�/5�����ۛ�����.��j:��}4��� ��L��ꢼ�أ��ڤ�0���,6��.���b������}A��;⮼�|��
��/���?hA���~��ئ��ź����������6����  �   gO=}�N=�oN=��M=d=M=�L=��K=�K=
FJ=�I=��H=�H=�TG=?�F=�F=9gE=��D=,AD=,�C=�7C=��B=_>B=��A=�6A=��@=�?=�K?="�>=ٽ==��<=�<=�K;=݆:=�9=M#9=��8=h�7=�}7=7=��6=�F6=��5=Ӆ5=u5=��4=|4=�~3=��2=5!2=re1=��0=��/=\-/=v.=G�-=9-=�a,=��+=v+=�V*=�)=��(=�6(='n'={�&=��%=u�$=uW#=� "=$� =A�=D=��=��=��=[�=� =�=+=�A=!Z=�s
=�=\�=��=�=v� =9��<��<<#�<���<*��<�R�<ȱ�<��<D��<h��<�v�<��<��<�7�<��<ճ�<!��<@m�<R�<0�<��<��<�F�<ƾ�<�</f�<=��<P�<�+�<w<��m<��d<�\<a�S<x5K<0C<�;<73<n[+<fp#<b<�!<ǧ
<"�<$�;r�;���;���;t{�;d�;�k�;�)g;��C;�� ;.�:ܸ�:w�h:ۇ�9�S츿��y؏�G�к�k	��+���M�	�p����nʛ�Rd��X����dϻ&y߻���:��0b����D��������� �J%��^)�֘-���1�" 6�/:��O>� TB��.F��I�>M�(kP�d^S��V���X�=
[��>]��I_��-a���b���d��Pf�jh�4�i��l�qin��q�C�s�Z�v���y���|����<R��.���Xك�T�K�\Ն�9���-a�����"Љ�q����q��ql��:���!ǎ�!������_��s��e򕼪Z��$������@G���}��]���ƞ��֟�۠��֡�VϢ��ͣ��ڤ�+ ���C�������-��̫�{���/���߰�H������׃��,۶���12��5��*"��t ���ؼ��  �  �JO=F�N=\N=��M=/M=��L=��K=�K=mSJ=�I=�H=�7H=ȎG={�F=�FF=o�E= 	E=�oD=��C=NC=��B=�?B=��A=^+A=|�@=m�?=R7?=�q>='�==��<=�;=?;=�G:=]�9=��8=K=8=��7=�;7=��6= u6=�6=L�5=Vk5=�5=��4=+4=Jq3=��2=�2=�k1=��0=�0=uV/=�.=��-=R-=�,=.�+=�9+=��*=E�)=�)=�<(=�j'=��&=>�%=-x$=?A#==�!=�j =I�=�=4J=�m=��=9�=��=��=��=��=y=#>
=d_=b{=��=r�=� =Q��<�}�<��<z��<�<�x�<���<o�<'��<!w�<r��<���<s�< ��<A�<S�<��<�}�<�Q�<]#�<j�<ꔠ<�$�<���<��<I"�<�P�<C|�<�_<��u<L�l<i�c<��Z<2gR<.J<�-B<�W:<~�2<5�*<�#<}<��<7d
<#�<���;�1�;�W�;ր�;��;�;�^�;�zk;�=H;M%;��;Cf�:�ts:3_�9�ȸϛ��ď�GyѺ5�	�r�+���N��q�gՊ�x՜������C���Gѻ��&�v~���y�X��g�T�����!�/u%���)���-�	2��06��M:��T>�7B�4�E��\I���L�@�O�EjR��U���W��Z��h\���^���`���b���d��Uf��0h�b(j�hOl�8�n��Xq��:t��Jw��tz��}��\�� Ձ��1���m�� ����}���T��D��$���Bc������Ɗ�B���@���駍��ގ��.��������/U������8 ��9G������eÚ����� 2���a��3�������L����Ƣ�nգ��3��ue���Ϩ�-[��s�����������F������K���#��Gp��)�������v���2���wW��2���  �  �+O=�N=VCN=,�M=)M=DrL=�K=�K=�YJ=��I=*I=�^H=�G=uG=x}F=�E=�6E=8�D=��C=�\C=e�B=s:B=W�A=2A=�~@=o�?=#?=�U>=9�==��<=Q�;=��:=�:=�I9=��8=��7=js7=��6=�6=XF6=��5=2�5=�M5=.�4=�v4=o�3=u^3=*�2=-2=>k1='�0=0=!v/=��.=�/.=��-=��,=�!,=d+=��*=
�)=;)=�;(=�`'=�w&=Xy%=�_$=K&#=��!=�I =h�=��=%=�3=�F=�V=�g=�|=��=Ϻ=+�=�
=�3=tU=,l=t=/k ==��<�R�<���<Xz�<��<O��<��<9��<�K�<���<�l�<���<t�<���<Ɓ�<��<�ĵ<�<�C�<�	�<�Ť<�l�<v��<la�<���<1܍<���<��<�}~<��t<��k<��b<;�Y<�bQ<�?I<�YA<��9<`�1<�M*<c�"<Õ<�l<�
<�}<���;!�;���;��;ګ�;0R�;���;o;1�K;(;�.;϶�:�c{:���9_Q���v�������Һ��
�3-�\�O�bZs�]���o睻L���*���*�һx�\��� �Xt���l7��^�d#��!�Y�%�!*�:.��[2�x6�_�:��t>�&6B���E�@I�dL�4�N�ޢQ�=T���V�JY���[��^��Z`�"|b�A�d�uf��hh��qj��l�o���q�-�t���w��{��X~�aƀ�@K��k���L��
������zȇ��x��������M������#΋������э�.��bH�����>풼�:���~��O����헼� ��hV��ܑ���ќ�J��_N��ā��̪���ˢ��飼E��;C���� �����a@��>���ׯ�S����h����Ֆ�����w)���5�����D�뫼��f���  �  8O=ɥN=�+N=2�M=M=aL=i�K='K=�ZJ=�I=XI=OzH=��G=�EG=ۥF=� F=�WE=&�D=�D=�dC=��B=�2B=��A=@A=^j@=�?=L?=G<>=�c==Ł<=�;=��:=��9=b9=
d8=��7=�@7=+�6=�q6=�6=��5=]�5=35=��4=�_4=��3=K3=O�2=_2=)g1=D�0=	'0= �/=��.=�S.=;�-=O -=UF,=��+=)�*=L�)=f)=d7(=vU'=�f&=sd%=�H$=#=}�!=, =��=��=^�=�=z=�=�.=LD="b=�=��=��	=0=�4=kN=xX=]Q =zs�<�(�<���<�d�<���<��<�>�<���<���<,�<���<jD�<���<4�<y��<�5�<@ε<sx�<"0�<<�<��<nD�<I˛<!1�<�u�<���<R��<Ƀ<v�}<�&t<G�j<�a<��X<N�P<��H<��@<�9<�p1<��)<�"<i/<�<�	<R5<�1�;���;���;Xm�;LS�;MB�;� �;�q;i�N;�D+;��;i��:�h�:{��97���Z�͑��Ժ@��8.�U!Q���t�Ɖ���՞�7��%û�aԻe�仠�������:�4S�M��N��z��R"�cM&��s*���.�E�2�s�6���:�.�>�!DB��E�G�H�m�K�uN��Q���S��'V���X��?[�ļ]��!`�gb���d�2�f���h���j���l�Lmo�7"r��u��Fx�;�{���~��������f���Z��s��l_�� %��K̈��`���"���o3��*����댼0����&���d��X����|,���^��I��������Ԙ����C��s���ٝ��%���k��/����֢�����/���j������E/��ê�w���C��n��m��������q��o����]������o����x��n=��������  �  �N=�N=�N=,�M=W�L=kTL=��K=b K=ZJ=�I=_ I=�H=��G=�]G=��F=\F=lE=��D=cD=[hC=��B=�+B=�A=�@=R[@=�?=3�>=!*>=`P==)l<=˃;=��:=?�9=V�8=�B8=�7=�7=V�6=zU6=v6=X�5=�r5=N 5=�4=O4=K�3=�<3=k�2=�2=�b1=E�0= .0=�/=�/=j.=��-=�-=�\,=�+=A�*=w�)=x)=�2(=rL'=	Z&=ZU%=�7$=��"=W�!=� =eq=V�=��=h�=O�=m�=i
= =#?=Cg=�=��	=��=�=�9=AE=2? =�Q�<�
�<1��<]T�<���<ߟ�<�O�<��<���<�[�<L��<ev�<��<�X�<JȾ<�C�<oе<qp�<��<�ը<T��<&�<˪�<7�<�O�<�t�<"��<���<sP}<ۤs<�;j<�%a<slX<TP<)H<K=@<��8<1<�)<'�!<��<t�<�y	<Y<,��;���;@��;���;i��;Sӛ;9؊;�Ts;�fP;^�,;p�;(��:}��:5�9몸�g��Ғ��ֺ����/�2R�i�u�%��z���̱�f�û�Iջ"��Ξ����ϻ����N�qW�����_"�ו&�Ƿ*���.���2�#�6���:���>��SB���E�!�H��K�|+N�;�P�:S��U��ZX���Z�\�]��`�`b�)�d���f��h�:�j��7m�H�o��gr�cu�F�x���{��T��S���悼�W��+����������a�����ʑ����������W��� ��T������A���z���������n&���L���i��;���.���0ԙ����]`��˶�����%`������]ᢼ����H������\ݧ��P���檼���Fm���K���*��>��������?��V���ӹ��ֺ�ܲ��)r���!��QϽ��  �  0�N=z�N=�N=V�M= �L=�OL=�K=*�J=�YJ=��I=�#I=U�H=��G=�eG=�F=- F=�rE=��D=�D=riC=�B=9)B=�A=?�@=�U@=�?=�>=�#>=bI==wd<=={;=	�:=��9=K�8='78=t�7=~7=æ6=�K6=�5=P�5=�k5=�5=��4=I4=��3=�73=��2=~�1=:a1=j�0==00='�/=�	/=vq.=��-=� -=d,=�+=��*=��)=�)=91(=I'=[U&=�O%=�1$=v�"=��!=U =�i=��=P�=��=
�=i�=.�=�=O3=D\=ۋ=T�	=��=<=3=�>=9 =TF�<� �<ت�<�N�<���<���<�U�<��<���<�k�<^�<
��<���<fd�<\о<�G�<;е<�l�<��<X̨<�{�<>�<P��<� �<�A�<Re�<�u�<s��<�&}<�ws<j<��`<�<X<�O<'�G<�@<%~8<��0< f)<5�!<E�<�<0e	<�� <<��;���;���;#��;;׬;Y�;�;�s;��P;n-;Qk	;s��:s�:��9ቫ�:���D��Φֺ,��z/�'yR�*=v��S������W��jĻ͛ջ�L�p����@�������u��z�4�|"��&�Y�*�j�.�93�7�;���>��YB���E�ūH��uK�:N�r�P�1S��U��<X���Z�t]���_��^b��d���f�h�h�W	k�UNm�1�o�Ԁr��}u��x��|�_x�Wg������8n������̆�5����u�������+������e���,��)���$��fK���;���F����$���F��`��<x�������Ù����R���������\�����f墼����Q�������觼�\��_󪼙���+|��F\���<��<��Ƶ�uV��T����鹼F캼ǻ�����Y2��b޽��  �  �N=�N=�N=,�M=W�L=kTL=��K=b K=ZJ=�I=_ I=�H=��G=�]G=��F=\F=lE=��D=cD=[hC=��B=�+B=�A=�@=R[@=�?=3�>=!*>=`P==)l<=˃;=��:=?�9=V�8=�B8=�7=�7=V�6=zU6=v6=X�5=�r5=N 5=�4=O4=K�3=�<3=k�2=�2=�b1=E�0= .0=�/=�/=j.=��-=�-=�\,=�+=@�*=w�)=x)=�2(=sL'=Z&=^U%=�7$=��"=f�!=� =�q=�=�=��=��=��=�
=� =�?=h=ߖ=v�	=��=�=;=iF=]@ =T�<@�<W��<]V�<���<s��<$Q�<��<e��<\�<b��<(v�<���<�W�<Ǿ<B�<�ε<�n�<��<eӨ<��<�#�<���< �<N�<)s�<���<f��<yN}<�s<�:j<�%a<mX<�P<H<�?@<ģ8<�1<�)<a�!<��<��<V~	<�<���;ǿ�;C��;��;c��;כ;�ڊ;Ws;?fP;D�,;��;e��:��:i��9|ͬ�ݪ� ���>ֺ����3/�<-R��u��%������ձ��ûxPջI��7����ѽ����YP��X����_`"�x�&�G�*�X�.�G�2�c�6�
�:�&�>��SB���E�4�H���K��+N�C�P�%:S��U��ZX���Z�^�]��`�`b�*�d���f��h�:�j��7m�H�o��gr�cu�F�x���{��T��S���悼�W��+����������a�����ʑ����������W��� ��T������A���z���������n&���L���i��;���.���0ԙ����]`��˶�����%`������]ᢼ����H������\ݧ��P���檼���Fm���K���*��>��������?��V���ӹ��ֺ�ܲ��)r���!��QϽ��  �  8O=ɥN=�+N=2�M=M=aL=i�K='K=�ZJ=�I=XI=OzH=��G=�EG=ۥF=� F=�WE=&�D=�D=�dC=��B=�2B=��A=@A=^j@=�?=L?=G<>=�c==Ł<=�;=��:=��9=b9=
d8=��7=�@7=+�6=�q6=�6=��5=]�5=35=��4=�_4=��3=K3=O�2=_2=(g1=D�0='0=�/=��.=�S.=9�-=M -=SF,=��+=(�*=J�)=e)=d7(=xU'=�f&=|d%=�H$=#=��!=., =�=B�=��=c==� =�/=gE=jc=i�=��=T�	=$=�6=�P=�Z=�S =�w�<3-�<���<�h�<1�<"��<A�<���<i��<L-�<���<�C�<��<]2�<7��<�2�<˵<�t�<3,�<�<8��<"@�<Ǜ<-�<r�<���<Z��<�ƃ<��}<�#t<��j<k�a<��X<ʖP<]�H<|�@<h9<�w1<"�)<""<�7<�<��	<�=<�A�;���;���;y�;�\�;�I�;_%�;��q;��N;�>+;R|;d�:?�:T5�9}ۯ����W��&պ�.��_.�HQ���t�����9瞻H#���ûNoԻH����1���>�{V������V���"��N&��t*�d�.��2���6�_�:�y�>�[DB��E�j�H���K�$uN�Q���S��'V���X��?[�ɼ]��!`�gb���d�4�f���h���j���l�Mmo�7"r��u��Fx�<�{���~��������f���Z��s��l_�� %��K̈��`���"���o3��*����댼0����&���d��X����|,���^��I��������Ԙ����C��s���ٝ��%���k��/����֢�����/���j������E/��ê�w���C��n��m��������q��o����]������o����x��n=��������  �  �+O=�N=VCN=,�M=)M=DrL=�K=�K=�YJ=��I=*I=�^H=�G=uG=x}F=�E=�6E=8�D=��C=�\C=e�B=s:B=W�A=2A=�~@=o�?=#?=�U>=9�==��<=Q�;=��:=�:=�I9=��8=��7=js7=��6=�6=XF6=��5=2�5=�M5=.�4=�v4=o�3=t^3=)�2=,2==k1=&�0=0=v/=��.=�/.=��-=��,=�!,=d+=��*=�)=:)=�;(=�`'=�w&=dy%=�_$=h&#=��!=�I =��=L�=�=o4=�G=�W=�h=~=a�=�={�=P
=�6=cX=>o==w=an =���<Y�<���<��<��<���<�#�<��<�M�<���<(m�<9��<�r�<���<�~�<��<b��<�y�<%>�<��<���<�f�<�<�[�</��<a׍<���<S�<{x~<:�t<��k<��b<��Y<BfQ<�DI<�`A<��9< 2<eX*<�"<�<4y<,
<��<���;{+�;��;�#�;u��;�\�;j��;to;.�K;G�(;�;���:a�z:���9�x��\.�����^Ӻ.�:?-� 
P���s�ԋ������� ���ӻۈ�!�F� ��y����M;��a�&�7�!��%��*�.;.��\2��x6��:��t>�y6B�ɾE�rI��L�R�N���Q�=T���V�)JY���[��^��Z`�%|b�D�d�uf��hh��qj��l�o���q�-�t���w��{��X~�aƀ�@K��l���L��
������zȇ��x��������M������#΋������э�.��bH�����>풼�:���~��O����헼� ��hV��ܑ���ќ�J��_N��ā��̪���ˢ��飼E��;C���� �����a@��>���ׯ�S����h����Ֆ�����w)���5�����D�뫼��f���  �  �JO=F�N=\N=��M=/M=��L=��K=�K=mSJ=�I=�H=�7H=ȎG={�F=�FF=o�E= 	E=�oD=��C=NC=��B=�?B=��A=^+A=|�@=m�?=R7?=�q>='�==��<=�;=?;=�G:=]�9=��8=K=8=��7=�;7=��6= u6=�6=L�5=Vk5=�5=��4=*4=Jq3=��2=�2=�k1=��0=�0=sV/=�.=��-=R-=�,=+�+=�9+=��*=C�)=�)=�<(=�j'=�&=M�%=Ex$=cA#=r�!=�j =��=u=�J=�n=��=��=P�=��=��=(�=N=AA
=�b=�~=~�=Q�=� =��<Z��<��<,��<	�<�}�<���<�r�<���<�x�<���<̓�<��<��</=�<��<q��<Lw�<K�<*�<�<x��<q�<���<W��<d�<jK�<�w�<VY<+�u<�l<G�c<��Z<~kR<�4J<U6B<�a:<F�2<Q�*<#<T<�<gs
<��<�; L�;3o�;'��;-ʪ;��;g�;؂k;M<H;��$;q�;.�:��r:� �9gθ�|��>����Ѻ�@
��#,��N��r���L�XҮ�&]���^ѻ���;�'���������k�D������!�Kw%�a�)��-�
2��16��N:�qU>��7B���E��\I�ٖL�e�O�bjR��U���W��Z��h\���^���`���b���d��Uf��0h�d(j�iOl�8�n��Xq��:t��Jw��tz��}��\�� Ձ��1���m�� ����}���T��D��$���Bc������Ɗ�B���@���駍��ގ��.��������/U������8 ��9G������eÚ����� 2���a��3�������L����Ƣ�nգ��3��ue���Ϩ�-[��s�����������F������K���#��Gp��)�������v���2���wW��2���  �   gO=}�N=�oN=��M=d=M=�L=��K=�K=
FJ=�I=��H=�H=�TG=?�F=�F=9gE=��D=,AD=,�C=�7C=��B=_>B=��A=�6A=��@=�?=�K?="�>=ٽ==��<=�<=�K;=݆:=�9=M#9=��8=h�7=�}7=7=��6=�F6=��5=҅5=t5=��4=|4=�~3=��2=4!2=qe1=��0=��/=Z-/=v.=E�-=6-=�a,=��+=r+=�V*=�)=��(=�6(=+n'=��&=�%=��$=�W#=*"=w� =��=�D=[�=��=��=��=�==�-=uD=H]=w
=я=^�=�=o�=Ԣ =��<U��<E+�<��<���<�X�<���<v�<��<���<w�<4��<Α�<_4�<V�<t��<܄�<;f�<{J�<(�<���<���<�>�<���<��<�_�<���<���<F(�<�v<L�m<��d<\<*�S<�<K<�C<($;<;D3<j+<)�#<�r<�2<��
<�<�C�;�6�;��;P»;��;<r�;Fu�;V2g;D�C;� ;���:z�:]Zh:e �91a����k`���cѺ޵	��g+��M�%�p�
+���뛻J����¾�=~ϻ�߻-��{L���i������g��4���� ��%��`)�V�-���1�6��/:�8P>�rTB��.F�\�I�B>M�QkP��^S��V��X�L
[� ?]��I_��-a���b���d��Pf�lh�5�i��l�rin��q�D�s�Z�v���y���|����<R��.���Xك�T�K�\Ն�9���-a�����"Љ�q����q��ql��:���!ǎ�!������_��s��e򕼪Z��$������@G���}��]���ƞ��֟�۠��֡�VϢ��ͣ��ڤ�+ ���C�������-��̫�{���/���߰�H������׃��,۶���12��5��*"��t ���ؼ��  �  B|O=5 O=zN=��M=�AM=��L=��K=B K=�/J=X_I=�H=��G=JG='aF=�E= E=�D=�
D=7�C=�C=¦B=�3B=]�A=l8A=��@=�@=�V?=�>=��==�==�C<=��;=!�:=E:=Co9=}�8=4E8=��7=�F7=��6=�j6=�6=��5=�'5=��4=�4=��3=��2=J2=+V1=�0="�/=�.=�9.=~-=��,=,=�n+=��*=N%*=W�)=n�(=|((=�h'=͓&=�%=�$=gd#=6"=n� =�=�m=��=�==r<=W=l=Q}=��=��=U�
=m�=��=��=��=*� =�<��<^/�<��<;��<z"�<g�<���<2�<Qk�<@��<�h�<��<(��<���<F`�<uM�<�B�<7�<i �<i��<ᯠ<9M�<ϗ<�:�<ᗎ<9�<�E�<䣀<ex<Ko<�f<�W]<5�T<�EL<�C<L�;<��3<�+<�#<�<>^<H�
<�<�)�;���;�M�;���;b�;���;\A�;�^b;�>;�;O��:嵯:ũ[:i��9�[��:$�յ���Һ�	�@M+�K|M��4p�,���'���N��r3��՛ͻ�kݻ
��Z����J�o�
����69��e�2< �<�$�m2)�}{-�O�1���5�d7:�p>�e�B�!�F�ZmJ��N��^Q��rT��BW��Y�� \��5^��`�!�a��^c���d��pf�Nh���i�&�k��Fn���p�k�s�<dv��Hy�d'|���~��̀����
@���Z��ya���T��o6��A
���Ո�k���Bt���Z��N\���~��Î�\&��⡑��+�������E��^ŗ�/5�����ۛ�����.��j:��}4��� ��L��ꢼ�أ��ڤ�0���,6��.���b������}A��;⮼�|��
��/���?hA���~��ئ��ź����������6����  �  5�O=�O=yN=a�M=u:M=$�L=ҼK=��J=�J=�6I=�_H==�G=9�F=�F=nE=��D=�KD=�C=A]C=��B=��B=�B=��A=�.A=֠@=�@=�V?=�>=��==�#==jg<=��;=� ;=�X:=��9=N9=��8=��7=�{7=��6=��6=�6=ɡ5=�)5=��4=\4=�y3=:�2=z	2=�=1=�k0=K�/=c�.=��-=C6-=�|,=,�+=�&+=*�*=V�)=uU)=f�(=)(=QY'=2�&=��%=Ғ$=�e#=j"=�� =i)=��=��=/(=#_=o�=1�=ʼ=`�=X�=;�=��
=�=��=�=��=ӳ =��<���<��<�p�<"��<x��<�
�<�>�<3��<���<�C�<���<�r�<�4�<�<��<S�<f�<��<��<7ߤ<��<dE�<�җ<=N�<���<�-�<랅<��<B)y<�6p<Vg<��^<��U< <M<�D<]r<<�;4<�,<�#<�<�Z<��
<Z�<q��;�.�;W�;E[�;�_�;D��;��;�U];�9;��;��:LW�:��M:���9�H9��+��V��" Ժ�
���+��M�O%p�L���l���M���ϻ�c�˻Pdۻ�\�����9�һ	���[��`��/����$� /)��-�2�1�H6��j:�|�>���B�?"G� K���N��cR���U�fuX�X[��D]�K=_���`��b���c�HJe�J�f��Gh�gj�Ll�;Qn���p�@js�/ v� �x�߈{��"~��Q��o���֬���ȃ��؄�݅��Ԇ�W����������g��pY��9c��]����Վ��@��ȑ�Fb�����!���6:��M���5&���t������+���緟�����=t��D��������j�\���?������&
��v���������\%������Y��q_��m����A#���I���b���n��r���  �  �O=��N=gnN=��M=;)M=HoL=^�K=�J=��I=�
I=�*H=�RG=~�F=��E=�#E=�D=WD=@�C=@*C=��B=�hB=�B=��A=�A=%�@=(�?=LM?=y�>=��==3==��<=��;=�3;=F�:=��9=/`9=��8=�68=J�7=|7=y�6=86=͡5=�"5=i�4=�	4=�g3=c�2=��1=X1=�E0=�h/=��.=��-=�,=33,=��+=��*=H*=n�)=�&)=��(=}�'=�A'=ew&=�%=M�$=�\#=�"=g� =�6=�=�=�Y=��=��=��= =�=M==��
=x�=0�=��=��=� =�<���<���<B�<�p�<���<��<J��<���<7D�<ݫ�<�5�<���<Ʊ�<"��<���<���<1˰<vج<�Ө<��<}�<�*�<�×<�O�<!֎<�\�<��<�w�<�z<Aq<�lh<%�_<��V</N<�lE<��<<D�4<|4,<*�#<��<�-<��
<��<
�;L�;�5�;��;M��;Ѐ�;�Q};�vX;^�4;�;�I�:}�:�?:B�92)b�Ǚ3�;����J׺:�-��N�g�p�ED��I��ߌ��窺�[ʻ�ٻf�Һ��@G����2��������S�$��P)���-��2��j6�^�:��?�xC��G�<�K���O�fS���V���Y�.\�b^�"B`�n�a�'@c��d���e��g��h��Uj��Nl�ȃn��p��ms���u���x��{��u}�����	��j)��PF��[`���u��=���)�������v��@l��|k�� ~��/�������5m������s����V��$	�� ����A��A����	���9���F���4���	��6Ρ�����Q���'�����X*���]��X������ȉ������t���ޯ��=������y೼^)���n������^鸼;���=���X���  �  �O=P�N=�]N=ҾM=�M=zVL=�K=خJ=��I=G�H=0�G=�G=�IF=>�E=%�D=cLD=��C=�\C=[�B=g�B=�EB=V�A=3|A=,A=z@=��?=�=?=��>=��==�:==^�<=�;=�[;=��:=a.:=��9=�8=5c8=.�7=I77=�6=o 6=8�5=�5=��4=��3=P3=�2=#�1=��0=e0=�;/=/Z.=�-=N�,=��+=�A+=��*=*=�)=B�(=m(=��'=�&'=�_&=�y%=�s$=�M#=�
"=� =�;=�=5$=��=s�=?=-=�@="D=�:=_)=p=4�=��=��=��=�� =���<nh�<���<-�<�0�<UB�<�M�<�_�<��<8��<�$�<���<�a�<>;�<%5�<�F�<�e�<���<���<�<P��<	P�<J�<���<�D�<�ގ<�{�<e�<Ł<��z<
r<�Si<Uz`<�W<?�N<;�E<�9=<��4<64,<U�#<+i<>�<�8
<rK<n5�;�S�;��;���;�	�;i��;�?y;x T;�(0;@u;��:�w�:�1:!1[9Gw��L�<�������ں����.�l�O�Vvq��l��晻�
��J̹� (ɻk$ػ���9�����:�������� ��d�$��)�.��o2���6��+;��?�e�C�EYH���L�ߖP��OT�[�W�h�Z�l7]�a_��-a���b��c�H#e��Mf���g��i�k�j�أl���n�d q���s�2�u��_x�h�z���|�m�Ȥ��Ӽ���ڂ������"���D��/_��p���x��S~��k�������׍��+��#���*9��3铼����og����������6��E�������Kß�h���n���$���֢����\_���J��X��>���?Ш�^-��q��������V�����J�c6���w��6���\���Q��霸�,⹼[��|M���  �  S�O=i�N=�LN=��M=��L=�>L=�pK=�J=u�I=��H=��G=w�F=�F=�WE=��D=5D=��C=�0C=�B=�|B=0'B=-�A=LcA=��@=Ud@=�?=H-?=��>=W�==�===��<=�
<=�x;=T�:=�U:=�9=�"9=b�8=��7=�F7=��6=�6=;�5=%5=0x4=�3=�93=ւ2=(�1=�0=��/=�/=`0.=�Q-=�,=Խ+=+=�o*=��)=#Y)=t�(=	M(=η'=�'=	I&=e%=�`$=s=#=5�!=)� =�<=P�=�6=<�=�=�/=�Y=Pm=�l=.]=�C=n%=/	=j�=��=O�={� =��<�?�< ��<���<���<� �<�<!	�<#�<U[�<��<�D�<���<Gܿ<9߻<P��<�!�<I�<�c�<�h�<hS�<&$�<�ߛ<��<�4�<�ގ<���<tC�<l��<�d{<��r<��i<� a<z,X<�2O<IBF<3l=<�4<7$,<�#<�,<��<@�	<+� <�n�;]u�;��;�j�;y��;�/�;zv;�P;�,;h
; |�:�k�:��&:�;49і��aD�����R޺�B���/��!Q��Xr�i���[ߙ�׻��3���JȻ�׻7������ ����M�����g������$�n�)�	X.�7�2��(7���;�G�?��rD�e�H��)M�@Q�U�`wX��x[�+	^��*`��a� Xc���d�էe���f�$�g��ei�tk�s�l�o��\q���s��v�=Ix��vz�a�|���~�AZ��yl���������焼S���E���h��~���q��������ʌ�����Y���Ӑ��n��>%���땼鴗��r��5��˜�����R$��&�����鿡�!m��>��Yɣ�y���nz������<�����PH����������oE����������:󱼰*��gk��}���L��Vf��Լ��(
���K���  �  OzO=l�N=�?N=ɛM=y�L=�-L=�^K=�J=9�I=��H=O�G=+�F="�E=P6E=�D="�C=Q|C=�C=2�B=�eB=mB=B�A=�QA=3�@={T@=��?=!?=�}>=V�==�===�<=�<=V�;=�:=3n:=��9=�99=ږ8=7�7=�O7=u�6=�6=ъ5=�4=�j4=��3=�)3=�q2=ۧ1=5�0=��/=N�.=�.=�3-=V_,=��+=��*={O*=��)=�=)=�(=m7(=}�'=R�&=�8&=�U%=�R$=-1#=~�!=!� =.;=��=�@=��=�=AI=u=v�=��=�q=�R=�.=b
	=D�=2�=V�= � =ؠ�<u!�<]~�<��<w��<H��<���<��<���<��<�u�<^ �<��<���</��<�Ƿ<���<��<G=�<�D�<`1�<��<pě<�w�<�'�<�ێ<햊<�X�<��<�{<�#s<Jhj<�a<�X<�zO<YtF<�=<K�4<b,<��#<1�<kg<��	<� <���;���;�b�;���;�۠;�9�;a�s;4N;�j*;�;vE�:W��:��:�9�n��&�I����,�ຶ]�� 1���Q�� s�nى�[晻Z���!ٸ���ǻghֻ���B�{� ��q���i�"_���{%���)��.�3��k7�>�;��H@�@�D�g6I���M�ŮQ�O�U�i�X�k�[��^���`�db�y�c���d�� f�Og�)Eh���i�YQk�;6m�6Oo�C�q�)�s��v�Ax��Vz��X|��T~��,��#;��.Z��R���Ä� ���8��g��p�����������a猼X"��&{������l���ON��t��藼ԫ��W���ޜ�i:��g���e���<������"���4A��>𣼦�������夦�'ͧ����]������0���c=���r�����nʱ�y����9��̇���㶼�E��n���� ���M���  �  !lO=f�N=�&N=D}M=\�L=�L=�FK=/uJ=ЛI=
�H=��G=�G=�DF=މE=��D=�GD=�C=�FC=o�B=�mB=�B=3�A=�!A=M�@=�@=N�?=&�>=�F>=D�==X==�h<=+�;=8;=D�:=	:=)n9=�8=�/8=Ȏ7=�6=R6=��5=�5=.�4=��3=uG3=ə2=��1=�1=�H0=�n/=(�.=��-=��,=g
,=\E+=��*=.�)=E;)=��(=��'=�Y'=P�&=��%=�%=�$=�#=��!=� =b=�=��= =i=��=�="8=�W=f=�f=7]=>M
=�9=$=/=��=9��<�F�<a��<�O�<6��<���<�/�<2b�<���<���<Q7�<G��<H�<��<Qܿ<�ϻ<�շ<�<���<��<<��<Gߣ<���<��<$>�<5��<��<�h�<�#�<%߁<�-{<�r<��i<6a<�JX<htO<�F<�=<R15<=�,<�$<t<e�<�
<W0<�6�;��;J��;���;=��;��;�;��Z;	H7;��;X��:��:\P:Ǎ�9�1�ol!����P8ͺPR��^&���F��f��h��n/��ج��ڱ�����`FϻK�ݻ����B��^J�׷	�T�� ���?�$y ��n%��-*�W�.��H3�&�7�7(<��@�#�D���H���L�$�P�FT��%W�p�Y�&6\��@^��
`�S�a�}'c�Ǧd��6f�/�g�,�i�|�k���m��p�Wfr�²t���v��1y��a{�ۍ}�Ͻ�m����!���N��k���ӳ���䆼���:���`��A���l���V���^��ѐ��Y��T�������mD���䘼s���盼�<���o�������v��:V���(��)����Σ�`���t���俦��秼�!��ah��N�������:G��򈯼8ư����pA��$���#ҵ�$���x���̹����yf���  �  �lO=�N=�(N=7�M=��L=�L=:KK=�yJ=�I=��H=>�G=�G=�LF=��E=!�D=�OD=��C=�MC=��B=�sB=�	B=͛A=�%A=�@=@=�?=i�>=6H>=��==�==vf<=��;=u3;=қ:=0:=h9=Q�8=�*8=Պ7=Y�6=�P6=ͷ5=� 5=$�4=��3=�J3=`�2=��1=1=fM0=jt/=@�.=V�-=�,=J,=rM+=��*=�)=�B)=K�(=(=�^'=�&=��%=�%=�"$=�#=��!=�� =�b=Y�=��=��=�d= �=j�=,1=�P=�_=�`=�X=�I
=�7=#=i=��=���<K�<���<uV�<ʵ�<d��<�9�<%n�<��<���<jG�<��<�X�<��<��<o޻<�<(�<���<D�<���<��<q��<��<�B�<���<�<�e�<�<�ց<}{<�wr<��i<�a<93X<Q`O<t�F<��=<�+5<X�,<
$<Rz<�<�!
<*=<�T�;E��; �;�"�;<+�;�S�;l�;�/[;T�7;>�;ޕ�:M�: �Q:���9���l����9�̺�� &�iF�6�f��^���/��;����ﱻ~���umϻ��ݻS�뻆m��]�Y�	�	��Ǽ�S?�9t �#f%��"*��.��93���7�	<�s@���D� �H�2�L�e�P�^�S��W���Y�\� #^���_�p�a�Mc�͒d��$f��g���i���k�N�m�dp��ar���t��v�#<y�	q{���}�x��p���-���Y��ȉ��庅��醼����9��0^��݆��칌�����LW���Ȑ��P��듼�����7���֘��c���כ�#,��i_��r��Qh���H�������ţ���������⸦��᧼����d������� ���J��򎯼�ΰ����M��K����ݵ��.������9ӹ�d ���g���  �  nO=:�N=a/N=a�M=M�L=HL=WK='�J=�I=��H=9�G=�*G=HcF=��E= E=.gD=��C=DbC=f�B=��B=TB=��A=�1A=i�@=T$@=�?=f�>=�K>=6�==�==�_<=n�;=�%;=��:=]�9=�U9=,�8=�8=�~7=�6=$L6=�5=#5=�4=��3==S3=4�2=��1=d*1=$[0=��/=��.=��-=��,=7),=e+=C�*=�)=X)=׶(=c(=6n'=t�&=��%=�%=�+$=f#=��!=u� =�c=1�=�~=��=�V=&�=$�=�=.<=jL=YP=4K=@
=�1=� =/=�=[��<
Y�<���<�i�<G��<��<2X�<+��<���<~�<�v�<���<���<3B�<V�<h�<�<y�<��<[!�<��<���<�џ<���<�M�<Y��<���<X[�<��<���<��z<g.r<�xi<2�`<��W<�%O<7fF<D�=<*5<#�,<�$<x�<��<qB
<\c<v��;R>�;Y��;���;�ƥ;��;g��;4�\;n9;�;���:ߪ:�1W:�m�9�����!2���˺�R��%���E�MXf�L��h9���ᢻ8���9��u�ϻ�A޻�G�j�����]�	���_���@�i �RP%�*��.�	3�|7���;��:@��|D�!�H�ƉL��7P���S�5�V��YY��[���]���_�Ea��b��Zd���e���g���i�s�k�O�m�b�o�lWr���t�Dw��[y�)�{�&�}�&���,��Q���z��ץ��aЅ�����7��19���W��^{�������덼�B�����T7��[Γ�p�� ��󭘼�7������L����/���D��>��g"��s���)Ϣ�/�������5��������Ч�����[��������\U��1����簼,���o������� ��;N������G湼�+���k���  �  �nO=%�N=�7N=Q�M=J�L=2,L=#hK=��J=F�I=T�H=3H=AKG=]�F=��E=o%E=��D=� D=�C=�C=ÜB=�-B=��A=BA=�@=�0@=]�?=�>=�O>=��==��<=1T<=��;=+;=�p:=|�9=�89=e�8=/8=k7=��6=�C6=�5=6%5==�4=��3=�^3=δ2=o�1=<1=Lo0=%�/=N�.=��-=�-=�L,=�+=1�*=�!*=6y)=��(=�/(=�'=�&=e&=�,%=28$=�)#=k "=ؽ =�c=c�=Ht=P�=j@=��=�=��=Y=�-=Q5=25=�/
=T'=�=$=��=/��<�k�<��<���<��<a@�<;��<���<=�<�[�<���<�<�<���<���<]�<�E�<@�<�C�<6I�<3H�<m:�<�<{�<穛<�Z�<=�<���<)H�<�<p��<nz<u�q<
�h<�<`<f}W<m�N<�F<�=<��4<̉,<)$<��<A<lo
<�<�-�;���;�:�;Oz�;Ե�;��;槁;�3_;m�;;��;�_�:-E�:�-_:N��9m�Ҹ�{�;����ȺT���$�?E���e�{<���V���.�����W���(�л�߻Y(��������>
�A=�����H��] ��4%��)��d.�8�2�?7�Ӛ;�Y�?�$D�+0H�$L�]�O��S��V�B�X��([��D]��$_���`�(sb�xd���e�ig�Mi��Zk���m�.�o��Lr���t�l,w�-�y�5�{�j<~�'C��g������t���Ԅ���W��C'��S;���P���l��N����ҍ�G&��b���F������B?��mۖ�jo��.�`�������坼���������砼�ơ����炣�*q���r��B�������B���GQ��V������h��I�������^������`��9��с���Ƹ�����@���t���  �  �lO=U�N=?N=�M=��L=$<L=�zK=��J=j�I=4I=�=H=�sG=��F=D�E=�TE=�D=,D=V�C=K/C=��B=GB=��A=$TA=>�@=�=@=R�?=��>=�Q>=G�==��<=�B<=v�;=-�:=M:=��9=H9=�w8=��7=�O7=@�6=o66=ͭ5=�$5=�4=\4=cj3=��2=22=�O1=��0=��/=��.=.=XB-=�y,=�+= +=�N*=�)=��(=�O(=/�'=��&=&=�;%=�D$=73#=�"=2� =La=m�=(d=��=q!=hi=U�=��=k�=W=�=�=�
=�="=)
=��=K��<}�<��<ޢ�<��<lm�<N��<��<�W�<���<��<G��<6�<O��<��<+��<�<�~�<�{�<�s�<`�<<�<��<켛<�d�<J�<��<}*�<ɾ�<�U�<n�y<Eq<�Th<e�_<��V<�AN<��E<�6=<��4<Xt,<�$<ȷ<�;<��
<��<��;Y��;4�;�v�;"ާ;Jb�;�;Pb;u ?;t�;�Z�:�Ŵ:�i:i
�9�ܖ�^��1Ԇ�FJƺhD���#�0�D���e��?������6���pg��;�»��ѻ�G�tW���tt�2�
����V��]�nZ �v%�x�)�\3.���2�"�6�WI;���?���C���G�syK��O��RR�RU�.X��qZ��\���^�T`� b��c��Ye�h$g�i�B+k�lm���o�KKr�
�t�D^w���y�dW|�ٿ~�n��������ق����O��'���4��=���C��lM���`�����鹍�-���m��l葼�r�����(����!��ۜ������R���������ê�����Ň���l���U��K��tR���o��������I��8������y����쯼�K����������O@��Ȇ���Ƿ�����4���_�������  �  �eO=c�N=�BN=E�M=�L=�IL=ӋK=��J=��I=�.I=�dH=g�G=,�F=�1F=j�E=$�D=�\D=��C=�TC=��B=b`B=�A=AdA=�@=nG@=�?=] ?=�O>=�==r�<=�+<=_x;=�:=y!:=�~9=��8=~J8=�7='-7={�6=�#6=��5=H 5=��4=O4=�r3=S�2=�2=b1=v�0=	�/=!/=�9.=�p-=5�,=��+=�4+=0�*=+�)=�")=4r(=�'=��&=#,&=�H%=5N$=V9#=I	"=6� =�Y=�=N=C�=	�=;<=	q=��=��=��=*�=A�=$�	=�=�=F=�=���<n��<�-�<h��<73�<��<x��<�O�<���<��<.��<
�<���<3P�<]�<��<≠<��<���<|��<K��<�V�<��<ɛ<g�<<��<j~�<a�<���<\�<�/y<�Up<G�g<]�^<�-V<��M<�,E<��<<L�4<�J,<�	$<�<.N<9�
<�<�9�;4(�;o��;.��;�!�;7ږ;���;��e;f�B;oH ;��:޺:��s:Mg�9-2���	��'���ĺ�\�m#�L/D��{e��e���򓻌H��:L���ûVӻ��Ứ��`E����$,�u��2a�����h �8%���)�5.�pk2���6�h�:�_*?��9C�. G�M�J��MN�u�Q��|T�j0W���Y���[��]�J�_�E�a�qJc��e���f���h�Ok�bVm�_�o�N[r���t���w�oHz���|�4`�j瀼����7��PQ���`���f���d��>]��^U���R��\���v�����BN������A���ǔ��M���˗��<��(����盼����@��)P��	P��FE��N6��*��4(���6��sZ��]���{樼�J��K���E5��u����%�����������P�������㶼���/K��?o������*����  �  �YO=��N=�@N=��M=�M=RL=U�K=��J=�J=�MI=�H=��G=�G= hF=��E=�#E=O�D=� D=qyC=�B=�vB={�A=�oA=��@=�K@=٩?={�>=H>=o�==��<=E<=%T;=��:=`�9=;J9=��8=�8=Ȋ7=�7=��6=�6=ܑ5=5=��4=�
4=wu3=H�2=L'2=�o1=�0=�/=V'/=Ab.=v�-=	�,=$,=bk+=&�*=@ *=!K)=K�(=��'=g'=�8&=�P%=)R$=�9#=�"=[� =HL=��=<2=I�=!�=8	=�8=�_=�=�=�=*�=��	=��=��=��=��=��<J��<F4�<k��<�L�<^��<�+�<���<� �<�s�<���<�z�<	�<��<&s�<|;�<��<��<qذ<ü�<㘨<�f�<h"�<�ɛ<$^�<�<�Z�<f͉<�?�<e��<ajx<�}o< �f<z�]<8_U<`�L<��D<�V<<�,4<Y
,<��#<J�<�I<��
<�<-��;	��;5��;��;qb�;�W�;pq�;�ti;�tF;��#;��;�
�:*f~:A�9Ȳ��������rº���"��D��e�۶��'����EY��1Ż2�Ի�D�#a�l���P������j�W��N���� �!&%��)��-��O2�ґ6�&�:�_�>���B���F��/J�B�M�{�P��S�ESV�j�X�k[�~?]�=_�!a���b���d�ǿf��h���j�SWm���o�r�r�W=u��x���z��x}�D��jL���~��8���z���?������Y���b���6r��|c���b���u��]�������Y8��N��������������u���ژ�f1��Fy��t���1ڝ�d���������������+��.%���O��>����騼�V��fӫ��Y��*㮼�h���屼{V��2���
��pK���|�����Q������VǼ��  �  DHO=��N=�8N=8�M=} M=1TL=�K=(�J=b&J=�hI=�H=��G=9GG=2�F=��E=KWE=w�D=V)D=��C=vC=��B=� B=vuA=��@=dI@=b�?=l�>=�:>=�y==��<=�;=�,;=bp:=ݼ9=�9=bu8=a�7=�Y7=��6=c6=`�5=~|5=�5=ω4=�4=�q3=��2=�*2=x1=��0=�0=�D/=~�.=��-=�-=eX,=��+=��*=�,*=�p)=Ұ(=8�'=^'=S@&=�R%=�O$=�3#=)�!=w� =9=�=O=�`=�=��=r�=�"=HC=�`=}=��=�	=�=�=�=�=���<ix�<5.�<���<�[�<���<Y�<���<!O�<���<,X�<8��<�~�<� �<J��<���<�O�<~!�<Q��<�Ѭ<루<�i�<1�<$��<mI�<�<�-�<���<��<w[�<��w<��n<Y�e<�]<��T<�&L<f�C<��;<]�3<J�+<Ţ#<x<*,<�
<<���;��;�C�;kd�;��;��;��;��l;�J;y';n>;Z��:��:�V:.q�6Ƀ��������~����"��fD�vOf�0���.��	 ��s�����ƻ�ֻ����6 �_��Si����'����� ��L%���)��	.��M2�'�6�؜:���>�VtB��F�#�I���L���O���R��~U��X��hZ���\���^�I�`���b���d�1�f���h��k��qm�Ep� �r��u�*px�ZO{�. ~��k������삼���l�������Sᇼ����������u��<�������ߎ�.��=���u󒼐]��ŕ��%��q}��;˙�	���H���x��6���(����͠�[ܡ��ꢼj������'R�����!���n������g���������*>��`����#���x��Ʒ���Ḽ����# ��,���d����  �  13O=߳N=Z+N=��M=V�L=�PL=[�K==�J=a4J=�~I=��H=�H=rG=��F=�&F=7�E=�D=�LD=��C=�$C=�B=bB=�uA=��@=�A@=v�?=r�>=4)>=�c==#�<=~�;=�;=�B:=��9=��8=@8=��7=(*7=[�6=�>6=8�5=d5=��4=Iz4=>�3=qh3=��2=�(2=w{1=��0=O0=G]/=��.=��-=�=-=>�,=��+=�+=�S*=Ȑ)=3�(=]�'=�$'=KB&=RO%=�G$=(#=I�!=� =�"=Q�=��=�8=eq=V�=��=W�=�=�(=XI=�i=X�	=��=O�=��=&�=���<6`�<��<���<m`�<t��<�{�<��<v��<�"�<X��<�H�<���<[{�<T�<˽<ʂ�<�D�<��<�ڬ<��<�`�<n�<���<@+�<��<��<�Q�<ʦ�<G�<��v<��m<��d<�1\<��S<[gK<CC<y=;<>H3<�T+<lS#<�7<��<�
<�<���;L�;m��;W�;�;���;}�;*p;�LM;��*;N(;R��:�B�:.�
:�H�70
���������O���:#�m	E��1g�Ȅ�F�������.����ǻJ�׻/��_����� ��:��n�2���p�%!���%���)�+.�!b2�O�6��:�,t>�&0B���E�.I��=L�9O��R�a�T��SW�C�Y�� \��[^�d`�.�b���d�.�f��h�@,k�_�m��Ap�(	s�E�u��x�"�{���~�.ʀ����oW�� y������cs���R���%��V�(Ɖ�@���j������������莼�.��5���Dܒ�=7������U���Y+��p��ʯ��*뛼�!���R���|��A�������Zۢ������%���_��ۭ����������������]�������������_����㶼� ��ZD���Q��"M���=���*���  �  MO=Q�N=�N=��M=��L=�IL=m�K=��J=O=J=��I=2�H=�:H=4�G=C�F=�MF=4�E=P	E=|iD={�C=�2C=|�B=�B=�qA=��@=o6@=��?=�>=�>=�L==?~<=ͭ;=/�:=�:=�]9=��8=�8=��7=0�6=��6=�6=7�5=�K5=>�4=�h4=N�3=\3=R�2=�"2=z1=)�0=z0=�o/=�.=G.=�a-=�,=w�+=_7+=�s*=s�)=��(=](=�('=@&=9H%=�<$=�#=)�!=� =u=�y=��=`=-G=�p=��=e�= �=�==1@=�d	=�=�=��=��=�g�<�B�<�<���<]�<4��<���<�.�<U��<�e�<� �<)��<�/�<���<}_�<���<��<�\�<k�<�ڬ<ߙ�<vP�<���<;��<��<%q�<�ȍ<M�<p_�< _<Jv<,m<�d<m[<!�R<�J<7�B<�:<�2<�*<�"<��<U�<Ee
<�<��;-_�;�;|��;�M�;<��;���;E�r;k�O;�@-;k�
;��:X��:�x:@8_B��H��Hº�I��#�$�E�98h�Ki��Ҹ��t姻�ø��(ɻ��ػ�绪��˱���4��~��
�v��-^!�F�%��*�CY.��2��6���:�'`>�1B�pE��H��K�^�N��pQ��"T�j�V��FY�}�[�^^��N`�}b�7�d���f�Bi�K\k���m���p��Zs�rOv��Wy�]c|�F`�C��'x��:���Wׄ��ۅ��Ɔ����cf��&+��~�xʊ�ȳ��߳���ˍ�X����7��-����Β�����d�������痼�$���`�������ڜ�i���L���~��H���1բ�� ��Z3���s���ǧ�2��,����H����ę���D��%岼|s��J鵼�B���}������𡺼����z���^���  �  
O=h�N=�N=�}M=�L=\AL=��K=U�J=ABJ=c�I=��H=�PH=1�G=�G=UkF=^�E={"E=+~D=��C=X<C=.�B=*B=lA=��@="+@=Z~?=��>=�>=)9==|g<=��;=��:=��9=k:9=��8=/�7=t\7=�6=�j6=6=��5={65=��4=oX4=�3=�O3=<�2=�2=�v1=p�0=9%0=|/=W�.=q).=�|-=��,=N,=SR+=�*=ռ)=(�(=(=�)'=<&=-@%=�1$="#=G�!=�o =��=�b=�=&�=\%=oK=Xl=��=b�=��=a�=�=�F	=�k==o�=t�=�G�<,'�<��<���<4V�<���<��<�J�<��<���<39�<+��<?k�<��<���< %�<ù<zk�<B�<6լ<&��<�=�<���<�o�<��<�K�<0��<��<\%�<�~<��u<�hl<�}c<+�Z<�dR<�1J<>-B<�H:<et2<S�*<B�"<J�<��<6
<��<��;�]�;�.�;&�;Pܭ;]��;ό�;`�t;.�Q;�3/;�U;�:��:��:ra18:J���<����º���Ќ$�f�F�>-i������a����������`&ʻm ڻl��?��5?�7g�-��m��h�}�פ!�_&�Q*�ʇ.��2���6�J�:�/Y>�r�A�s<E��bH��^K�h9N���P�~�S��QV���X�Qj[��]��0`�Hub���d�k�f�J+i�9�k��n���p��s�7�v�D�y�w�|����b��D���� ���!��0#��	���؇�a���dY������튼�ҋ��Ό��⍼����C��儑��Ȓ�p
���G��J��������옼X&��d��ȥ���蝼U*���g��#����Ԣ�	��C�����᧼5O���Ԫ��n������˯�m}���$��ݸ���2��n����Ǹ�|⹼E⺼�ͻ�}���Ҋ���  �  ��N=��N=5N=ntM=��L=	;L=��K=:�J=wDJ=]�I=k�H=�]H=�G=G=�}F=��E=�1E=��D=��C=tAC=��B=`B=gA=�@=�"@=�t?=�>=y�==�+==5X<={�;=E�:=~�9=�#9=�r8=D�7=E7=�6=\V6=��5=ދ5=1(5="�4=M4=��3=�F3=��2=�2=�s1=Y�0=�(0=R�/=0�.=�7.=�-=��,=-$,=�b+=3�*=��)=j�(=U(=�)'=�8&=�9%=E)$=2#=	�!=jc =��=�R=N�=m�=m=�3=S=�q=z�=۶=��=;	=f3	=0Z=Jz=��=��=:1�<s�<V��<T��<MP�<���<���<C[�<
�<ߵ�<1\�<g��<���<��<���<;�<�ѹ<�r�<��<�Ϭ<��<�/�<Aϟ<�[�<�і<2�<��<��<"��<̆~<�.u<�l<�c<�nZ<�R<��I<��A<� :<-42<Fd*<+�"<�<`\<�
<q�<d�;�V�;,D�;�7�;�1�;+�;?�;��u;>S;�g0;ok;��:�@�:pw:m?8�:��'����púA�9%�+EG���i�&]���ԗ�.���:��j�ʻ��ڻS��2������A��=l����;���V���!�3&�!x*�]�.���2���6���:�fX>���A��E�66H�Z%K�Z�M�r�P��dS��V���X��<[��]�>!`��sb���d���f��Hi���k��;n�5�p�!�s���v���y�}����������0��AQ��+Q���3�� ��B���Zx��8��2���苼�⌼
􍼗��qM��$����ƒ����6��h��Q���|ʘ� ���@��n����͝���[��隡�<֢�z��KO��蘦���d���몼����L6���쯼����N���崼�a��B�������������c��μ������  �  <�N=^�N=c�M= qM=�L=�8L=�K=��J=EJ=T�I=� I=FbH=r�G=[%G=��F=��E=7E=ƎD=��C=CC=��B=�B=�eA=��@=�@=(q?=�>=�==�&==�R<={|;=��:=1�9=�9=�j8=�7=	=7=��6=SO6=��5=8�5=#5=��4= I4=:�3=�C3=��2=�2=Gr1=*�0=�)0=��/=��.=9<.=��-=��,=*,=xh+=��*=n�)=��(=\(=K)'=:7&=�7%=N&$=��"=��!=�^ =��=qM=1�=��=�=�+=tJ=�h=ǉ=k�=�=�=�,	=dT=u=ڋ=̖=�)�<��<��<\��<XN�<%��<���<�`�<>�<C��<h�<��<��<*�<��<B�<?ֹ<Yt�<��<�̬<�}�<�)�<Lȟ<�S�<ɖ<N(�<�t�<ٴ�<r�<�h~<�u<��k<��b<�LZ<��Q<�I<0�A<��9<�2<Q*<p"<�q<�N<�
<٤<&Y�;�T�;^L�;�J�;"O�;fR�;OF�;�=v;��S;�0;`�;�y�:{��:� :KB8vu���ŀ���ú�n�UG%�A�G��!j�U�������^���p���˻w�ڻd껓<��к�4�������t���j���!��B&�w�*��.�M�2�#�6�a�:��X>�o�A��E��'H�4K���M���P��LS�>�U��X��-[��]�b`��sb�1�d�/g�+Si���k�QJn�bq�#�s���v�z�1}�}#��y��������@���a���`���B�����iʈ�4����A��������錼H������JQ�����$ƒ����1��`��.������������4���z���ĝ�e���V��_��� ע�����S������j����k��1��������@��Z�������^\�������q���ͷ������`��� ���ڼ�����  �  ��N=��N=5N=ntM=��L=	;L=��K=:�J=wDJ=]�I=k�H=�]H=�G=G=�}F=��E=�1E=��D=��C=tAC=��B=`B=gA=�@=�"@=�t?=�>=y�==�+==5X<={�;=E�:=~�9=�#9=�r8=D�7=E7=�6=\V6=��5=ދ5=1(5="�4=M4=��3=�F3=��2=�2=�s1=X�0=�(0=R�/=0�.=�7.=�-=��,=-$,=�b+=3�*=��)=j�(=U(=�)'=�8&=�9%=J)$=9#=�!=xc =�=S=p�=��=�=�3=^S=r=�=_�=y�=�	=4	=�Z={=c�=ܛ=�2�<2�<	��<��<�Q�<���<���<B\�<�
�<l��<�\�<x��<ɏ�<��<��<5:�<�й<Wq�<1�<ά<䀨<�-�<�͟< Z�<0Ж<�0�<A~�<࿈<.��<R�~<�-u<	l<�c<RoZ<�R<f�I<��A<>:<�62<4g*<S�"<7�<�_<b
<��<gj�;s\�;lI�;<�;i5�;�-�;�;Q�u;�=S;Pe0;g;_��:�0�:P:�4<8����������úP�i %�OTG���i�Nd���ۗ�f4���@����ʻj�ڻ�������V�����am������wW�Z�!�n3&�xx*���.��2��6���:��X>���A��E�C6H�d%K�b�M�x�P��dS��V���X��<[��]�?!`��sb���d���f��Hi���k��;n�5�p�!�s���v���y�}����������0��AQ��+Q���3�� ��B���Zx��8��2���苼�⌼
􍼗��qM��$����ƒ����6��h��Q���|ʘ� ���@��n����͝���[��隡�<֢�z��KO��蘦���d���몼����L6���쯼����N���崼�a��B�������������c��μ������  �  
O=h�N=�N=�}M=�L=\AL=��K=U�J=ABJ=c�I=��H=�PH=1�G=�G=UkF=^�E={"E=+~D=��C=X<C=.�B=*B=lA=��@="+@=Z~?=��>=�>=)9==|g<=��;=��:=��9=k:9=��8=/�7=t\7=�6=�j6=6=��5={65=��4=oX4=�3=�O3=<�2=�2=�v1=p�0=9%0=|/=V�.=p).=�|-=��,=M,=QR+=�*=Լ)=(�(=(=�)'="<&=3@%=�1$=0#=[�!=
p =�=�b='�={�=�%=�K=�l=j�=?�=��=��= =)H	=m=V�=�=$�=
K�<�*�<���<��<Y�<w �<i��<�L�<���<���<�9�<L��<�j�<M��<���<O#�<���<i�<��<EҬ<��<�:�<�ݟ<�l�<��<I�<���<}��<�#�<?�~<��u<�gl<�}c<�Z<�fR<Q4J<�0B<[M:<|y2<��*<\�"<��<%�<�<
<�<B��;�h�;�8�;�
�;��;ֽ�;n��;��t;��Q;X//;LM;���:���:�a:��+8���}q���ú���(�$���F��Ii�����n��Ѷ��鰹��0ʻ�	ڻ���F��HB��i�b��o�;j�� �ڥ!�0&��Q*�P�.�q�2��6���:�bY>���A��<E��bH��^K�w9N���P���S��QV���X�Uj[��]��0`�Jub���d�l�f�K+i�:�k��n���p��s�7�v�D�y�w�|����b��D���� ���!��0#��	���؇�a���dY������튼�ҋ��Ό��⍼����C��儑��Ȓ�p
���G��J��������옼X&��d��ȥ���蝼U*���g��#����Ԣ�	��C�����᧼5O���Ԫ��n������˯�m}���$��ݸ���2��n����Ǹ�|⹼E⺼�ͻ�}���Ҋ���  �  MO=Q�N=�N=��M=��L=�IL=m�K=��J=O=J=��I=2�H=�:H=4�G=C�F=�MF=4�E=P	E=|iD={�C=�2C=|�B=�B=�qA=��@=o6@=��?=�>=�>=�L==?~<=ͭ;=/�:=�:=�]9=��8=�8=��7=0�6=��6=�6=7�5=�K5==�4=�h4=N�3=\3=R�2=�"2=z1=)�0=y0=�o/=�.=F.=�a-=�,=v�+=]7+=�s*=q�)=��(=](=�('=#@&=AH%=�<$=�#=E�!=2� =�=/z=��=�=�G==q=��=p�=9�=}�=�=�A=�f	=��=(�=S�=�=�l�<�G�<��<���<+a�<���<ɗ�<�1�<x��<lg�<|�<X��<3/�<���<�]�<6��<(��<}Y�<��<V֬<{��<�K�<N�<Ɔ�<x�<+m�<�č<*�<�\�<[<�v<��l<td<Nn[<��R<ҾJ<Y�B<[�:<;�2<�*<�#<��<��<�n
<�< ��;$o�;l�;㱾;�W�;��;��;�r;��O;e:-;t�
;���:�_�:':E8�V��o:��R`º�r��	$��F��`h��|��a˖������Ӹ�7ɻ��ػ��综&��#�����S����9���_!�n�%��*� Z.���2���6��:�p`>�jB�KpE�A�H��K�s�N��pQ��"T�s�V��FY���[�c^��N`�}b�9�d���f�Di�L\k���m���p��Zs�sOv��Wy�^c|�F`�C��'x��:���Wׄ��ۅ��Ɔ����cf��&+��~�xʊ�ȳ��߳���ˍ�X����7��-����Β�����d�������痼�$���`�������ڜ�i���L���~��H���1բ�� ��Z3���s���ǧ�2��,����H����ę���D��%岼|s��J鵼�B���}������𡺼����z���^���  �  13O=߳N=Z+N=��M=V�L=�PL=[�K==�J=a4J=�~I=��H=�H=rG=��F=�&F=7�E=�D=�LD=��C=�$C=�B=bB=�uA=��@=�A@=v�?=r�>=4)>=�c==#�<=~�;=�;=�B:=��9=��8=@8=��7=(*7=[�6=�>6=8�5=d5=��4=Iz4==�3=qh3=��2=�(2=v{1=��0=N0=F]/=��.=��-==-=<�,=��+=�+=�S*=Ɛ)=2�(=^�'=�$'=PB&=[O%=�G$=2(#=k�!=M� =$#=��=�= 9=r=8�=��=��=I
=�*=KK=	l=��	=<�=	�=v�=�=��<f�<E#�<��<ve�<��<��<?
�<��<b$�<d��<�H�< ��<�y�<!�<#Ƚ</�<�@�<�	�<�լ<���<\[�<��<��<&�<&��<���<'N�<���<��<-�v<�m<��d<u3\<�S<)lK<cIC<E;<Q3<p^+<�]#<C<<Z�
<�<���;�_�;��;�+�;m��;b�;P��;p;�KM;ə*;�;���:=�:/1
:E�7�\��U��a���g��m#�<E��cg�����
�����������ǻ@�׻N�滴�����?������՝��r��!� �%���)��+.��b2���6�Y�:��t>�l0B�ۻE�XI��=L��9O�R�p�T��SW�L�Y�� \��[^�i`�1�b���d�0�f��h�A,k�`�m��Ap�)	s�E�u��x�"�{���~�.ʀ����pW�� y������cs���R���%��V�(Ɖ�@���j������������莼�.��5���Dܒ�=7������U���Y+��p��ʯ��*뛼�!���R���|��A�������Zۢ������%���_��ۭ����������������]�������������_����㶼� ��ZD���Q��"M���=���*���  �  DHO=��N=�8N=8�M=} M=1TL=�K=(�J=b&J=�hI=�H=��G=9GG=2�F=��E=KWE=w�D=V)D=��C=vC=��B=� B=vuA=��@=dI@=b�?=l�>=�:>=�y==��<=�;=�,;=bp:=ݼ9=�9=bu8=a�7=�Y7=��6=c6=`�5=~|5=�5=ω4=�4=�q3=��2=�*2=x1=��0=�0=�D/=}�.=��-=~-=cX,=��+=��*=�,*=p)=Ұ(=9�'=a'=Z@&=�R%=�O$=�3#=O�!=�� =�9=x�=�=ka=�=��=��=h$=�D=�b=0=L�=��	=��=�=��=K�=���<�~�<�4�<���<_a�<���<s]�<���<R�<���<WY�<x��<E~�<7�<���<a��<�K�<��<��<�ˬ<Ꝩ<�c�<��<��<�C�<*��<�(�<>��<h��<�X�<4�w<��n<?�e<�]<��T<=,L<f�C<#�;</�3<6�+<��#<p�<�8<��
<^+<m��;q*�;"W�;bu�;���;�ə;��;h�l;�J;<p';.;
��:�׃:��:Ҍ�6�~ �X���º_��6#�G�D�цf��J���G�����H�����ƻ�"ֻ������; �o���m�����*����� �{N%�ض)��
.�ON2�ɀ6�X�:��>��tB��F�S�I���L��O��R��~U��X��hZ���\���^�M�`���b���d�4�f���h��k��qm�Fp�!�r��u�*px�ZO{�. ~��k������삼���l�������Sᇼ����������u��<�������ߎ�.��=���u󒼐]��ŕ��%��q}��;˙�	���H���x��6���(����͠�[ܡ��ꢼj������'R�����!���n������g���������*>��`����#���x��Ʒ���Ḽ����# ��,���d����  �  �YO=��N=�@N=��M=�M=RL=U�K=��J=�J=�MI=�H=��G=�G= hF=��E=�#E=O�D=� D=qyC=�B=�vB={�A=�oA=��@=�K@=٩?={�>=H>=o�==��<=E<=%T;=��:=`�9=;J9=��8=�8=Ȋ7=�7=��6=�6=ܑ5=5=��4=�
4=vu3=H�2=K'2=�o1=�0=�/=T'/=@b.=t�-=�,=$,=_k+=$�*=> *=K)=J�(=��'=j'=�8&=�P%=;R$=�9#="=�� =�L=V�=�2=�=��==
=:=`a=Ł=�=(�=��=��	=��=��=��=��=���<��<�:�<���<uR�<���<E0�<x��<��<�u�<(��<
{�<W�<L��<�p�<8�<��<��< Ӱ<޶�<���<g`�<��<�Û<X�<�ܒ<�U�<�ȉ<<�<���<zfx<�{o<�f<L�]<�bU<��L<��D<a_<<&74<�,<��#<�<�V<��
<c)<���;���;���;���;�p�;�b�;�x�;G{i;�sF;��#;��;���:��}:���9��������m����º����"�[SD�c�e�w҃�[����-���o���EŻ��Ի�T�ao����������kn�d������� ��'%�8�)� .��P2�z�6���:���>���B��F��/J�h�M���P��S�WSV�x�X�v[��?]�=_�!a���b���d�ɿf��h���j�TWm���o�s�r�W=u��x���z��x}�D��jL���~��8���z���@������Y���b���6r��|c���b���u��]�������Y8��N��������������u���ژ�f1��Fy��t���1ڝ�d���������������+��.%���O��>����騼�V��fӫ��Y��*㮼�h���屼{V��2���
��pK���|�����Q������VǼ��  �  �eO=c�N=�BN=E�M=�L=�IL=ӋK=��J=��I=�.I=�dH=g�G=,�F=�1F=j�E=$�D=�\D=��C=�TC=��B=b`B=�A=AdA=�@=nG@=�?=] ?=�O>=�==r�<=�+<=_x;=�:=y!:=�~9=��8=~J8=�7=&-7={�6=�#6=��5=H 5=��4=N4=�r3=S�2=�2=b1=u�0=�/= /=�9.=�p-=3�,=��+=�4+=.�*=)�)=�")=4r(=�'=��&=),&=�H%=FN$=p9#=o	"=l� =�Y=w�=�N=�=��=8==;r= �=O�=t�=V�=��=��	=�=�=r=E�=��<��<H4�<s��<�8�<��<���<ES�<��<��<Y��<Y
�< ��<�N�<��<H�<5ȸ<O��<C��<ʖ�<I{�<�P�<T�<�<2a�<��<�y�<��<���<��<�+y<�Sp<-�g<�^<r1V<��M<�3E<!�<<�4<�U,<�$<f�<�Z<��
<<8Q�;>�;��;,��;�/�;��;�Ȅ;��e;F�B;�? ;���:���:�Is:*@�9|�<��C
����� |ĺe��R#��gD�%�e�s���@��4`��	b����ûӻ<��h��?Q����j0���&d����j ��%�͠)�9.�>l2���6���:��*?��9C�k G�}�J��MN���Q��|T�{0W���Y���[�	�]�P�_�J�a�tJc��e���f���h�Pk�cVm�_�o�O[r���t���w�oHz���|�5`�j瀼����7��PQ���`���f���d��>]��^U���R��\���v�����BN������A���ǔ��M���˗��<��(����盼����@��)P��	P��FE��N6��*��4(���6��sZ��]���{樼�J��K���E5��u����%�����������P�������㶼���/K��?o������*����  �  �lO=U�N=?N=�M=��L=$<L=�zK=��J=j�I=4I=�=H=�sG=��F=D�E=�TE=�D=,D=V�C=K/C=��B=GB=��A=$TA=>�@=�=@=R�?=��>=�Q>=G�==��<=�B<=v�;=-�:=M:=��9=H9=�w8=��7=�O7=@�6=o66=̭5=�$5=�4=\4=bj3=��2=12=�O1=��0=��/=��.=.=WB-=�y,=�+= +=�N*=�)=��(=�O(=0�'=��&=&=�;%=�D$=O3#=�"=b� =�a=��=�d=D�=)"=Kj=g�=��=��==�==?
=%=�==��=1��<��<n"�<I��<��<�q�<L��<�<XZ�<���<��<���<{5�<���<а�<:��<U��<Uz�<�v�<�n�<�Z�<�6�<���<y��<�_�<n��<���<�&�<���<S�<�y<�q<�Th<��_<��V<�FN<�E<I>=<��4<~,<&$<��<#G<�
<��<��;���;��;ꅺ;��;�k�;h$�;�Ub;r?;��;o=�:��:�h:��9נ�����/��3�ƺ�v�z�#���D��e��W��9���i����z����»��ѻ�U��c�e����x��
������_�2\ ��%���)�E4.�<�2���6��I;��?��C�׬G��yK��O��RR�*RU�>X��qZ��\���^�T`�%b��c��Ye�j$g�i�C+k�lm���o�LKr��t�E^w���y�dW|�ٿ~�n��������ق����O��'���4��=���C��lM���`�����鹍�-���m��l葼�r�����(����!��ۜ������R���������ê�����Ň���l���U��K��tR���o��������I��8������y����쯼�K����������O@��Ȇ���Ƿ�����4���_�������  �  �nO=%�N=�7N=Q�M=J�L=2,L=#hK=��J=F�I=T�H=3H=AKG=]�F=��E=o%E=��D=� D=�C=�C=ÜB=�-B=��A=BA=�@=�0@=]�?=�>=�O>=��==��<=1T<=��;=+;=�p:=|�9=�89=e�8=/8=k7=��6=�C6=�5=6%5==�4=��3=�^3=δ2=n�1=<1=Ko0=$�/=M�.=��-=�-=�L,=�+=/�*=�!*=4y)=��(=�/(=�'=�&=j&=�,%=?8$=�)#=� "=�� =3d=��=�t=��= A=d�=��=��=�=/=�6=�6=�1
=l)=4=v=?�=���<lp�<(
�<��<$��<D�<~��<���<b�<=]�<���<�<�<��<g��<6[�<C�<=�<{@�<\E�<D�<6�<��<��<t��<XV�<F��<���<	E�<i�<n��<Qkz<�q<��h<>`<�W<T�N<�F<9�=<�5<Ƒ,<�#$<Ȯ<�$<�x
<��< ?�;���;�H�;Ć�;��;`�;��;U8_;��;;)�;�G�:i"�:��^:���9?�ָ5�/���-ɺ�|��$�VhE�f��O��'i��@���Ĳ�����)�лe)߻j2�j������B
��?����SJ��^ �6%���)��e.���2��?7�1�;���?�]D�X0H�GL�x�O��S��V�N�X��([��D]��$_���`�+sb�{d���e�
ig�Mi��Zk���m�/�o��Lr���t�l,w�-�y�5�{�j<~�'C��g������t���Ԅ���W��C'��S;���P���l��N����ҍ�G&��b���F������B?��mۖ�jo��.�`�������坼���������砼�ơ����炣�*q���r��B�������B���GQ��V������h��I�������^������`��9��с���Ƹ�����@���t���  �  nO=:�N=a/N=a�M=M�L=HL=WK='�J=�I=��H=9�G=�*G=HcF=��E= E=.gD=��C=DbC=f�B=��B=TB=��A=�1A=i�@=T$@=�?=f�>=�K>=6�==�==�_<=n�;=�%;=��:=]�9=�U9=,�8=�8=�~7=�6=$L6=�5=#5=�4=��3==S3=3�2=��1=d*1=$[0=�/=��.=��-=��,=6),=e+=B�*=�)=X)=ֶ(=c(=7n'=v�&=��%=�%=�+$=t#=��!=�� =�c=d�=(=I�=SW=��=��=b=
==hM=xQ=tL={A
=/3=`"=�=��=®�<k\�<���<�l�<0��<<�<�Z�<��<f��<��<w�<���<7��<aA�<�<��< �<
�<��<g�<��<���<pΟ<[��<�J�<���<��<"Y�<�	�<Q��<��z<d-r<�xi<�`<��W<b(O<�iF<��=<;!5<Ǘ,<�$<ܓ<J�<�H
<�i<���;�I�;���;q��;Υ;D�;��;��\;�m9;�;��:nƪ:M�V:�Դ9\-�Ӂ�#g���;˺�o�e�%��F��tf��Y��|F��[C��D����ϻ�I޻�N컐��������	��	�����A�j �%Q%��*�h�.�t3��7���;�;@��|D�@�H�߉L��7P���S�A�V��YY��[���]���_�!Ea��b��Zd���e���g���i�t�k�O�m�b�o�lWr���t�Dw��[y�)�{�&�}�&���,��Q���z��ץ��aЅ�����7��19���W��^{�������덼�B�����T7��[Γ�p�� ��󭘼�7������L����/���D��>��g"��s���)Ϣ�/�������5��������Ч�����[��������\U��1����簼,���o������� ��;N������G湼�+���k���  �  �lO=�N=�(N=7�M=��L=�L=:KK=�yJ=�I=��H=>�G=�G=�LF=��E=!�D=�OD=��C=�MC=��B=�sB=�	B=͛A=�%A=�@=@=�?=i�>=6H>=��==�==vf<=��;=u3;=қ:=0:=h9=Q�8=�*8=Պ7=Y�6=�P6=ͷ5=� 5=$�4=��3=�J3=`�2=��1=1=fM0=jt/=@�.=U�-=�,=J,=qM+=��*=�)=�B)=J�(=(=�^'=�&=��%=�%=�"$=�#=��!=�� =�b=t�=�=��=�d=D�=��=�1=Q=`=�a=6Y=�J
=G8=�#=B=��=\��<�L�<���<X�<L��<� �<;�<%o�<��<8��<�G�<���<�X�<v�<.�<�ݻ<
�<��<9��<��<���<$�<ȼ�<f��<QA�<E��<���<wd�<#�<�Ձ<{{< wr<��i<Ca</4X<�aO<R�F<��=<>.5<C�,<0$<�}<i�<%
<{@<[�;"��;f�;D'�;�.�;�V�;2�;z1[;�7;ޅ;��:���:$�Q:���9=��-0 �i��1�̺��/&�5xF��f��e��K6��������������7rϻ��ݻ�뻴p��_^��	��������?��t ��f%�R#*�_�.�:3��7�+<�"s@�	�D�1�H�?�L�n�P�f�S��W���Y�\�#^���_�r�a�Nc�Βd��$f��g���i���k�O�m�dp��ar���t��v�#<y�	q{���}�x��p���-���Y��ȉ��庅��醼����9��0^��݆��칌�����LW���Ȑ��P��듼�����7���֘��c���כ�#,��i_��r��Qh���H�������ţ���������⸦��᧼����d������� ���J��򎯼�ΰ����M��K����ݵ��.������9ӹ�d ���g���  �  lXO=��N=:N=TcM=��L=��K=8K=SpJ=��I=��H=�H="?G=�~F=3�E=�E=,�D=��C=(lC=\�B=�rB=��A=�|A=��@=,r@=��?=NJ?=�>=�>=�h==�<=�$<=��;=��:=EI:=Q�9=\9=Pl8=u�7=x*7=^�6=��5=�M5=C�4=�4=�m3=��2=a2=�X1=&�0=�/=��.=� .=+J-=v,=�+=U�*=�*=#b)=��(=��'=QA'=��&=�%=��$=��#= #=L�!=}� =I�=)0=��=T=+�=s6=�=
�= =�;=�W=�g=$n=�m	=�g=�]=�O=&<=�C�<���<7��<o9�<H��<�(�<̌�<���<KM�<��<p2�<��<g�<�$�<���<�߻<"Է<�ϳ<�̯<�ī<���<���<�n�<*;�<���<���<�w�<�1�<��<"��<Ÿz<�r<}i<��`<#!X<DoO<[�F<�><%�5<��,<�t$<"�<�R<٤
<\�<���;���;А�;�5�;�٨;���;��;\�e;��B;�� ;
g�:��:�}:{ :��_7(��;du�aS���Z�� ��+�;��A[���z��ጻ`,��0��9湻MOȻ�iֻ�0�D�������ե��j�=���)��-!� &��*�0:/��3�k8�Uc<��@���D�t�H�I-L�ٓO���R�>�U�?X��jZ�	�\�|^�-Z`��0b�Gd���e�yh�~(j�dl��n�*q�ks��u��x�nz���|�'�謀��؁�����8��Wj��<��� ȇ���q"���T�������׍�//��җ��A��B����!�������5��T������Kg��ʟ������͟��ɠ�z���׬��g���������=ʦ������2��'x��Lë�B��?\��ԥ���찼�2��@y��7´�����[�����������C��ꋼ��  �  dXO=7�N=sN=eM=	�L=o�K=�:K=�sJ=R�I=�H=FH=SDG=p�F=�E=�%E=��D=�C=CqC=��B=�vB=��A=�A=��@=�t@=��?=�K?=�>=L>=�h==�<=�"<=E�;=F�:=E:=�9=�9=h8=��7=]'7=�6=4�5=WM5=~�4=�4=Lo3=|�2=�2=�[1=%�0=v�/=��.=%.=	O-=c{,=��+=1�*=�"*=�g)=H�(=|�'=�E'=R�&=I�%=]�$= $=�#=��!=�� =ڃ=0=��=7R=u�=�2=j�=�=�=�6=�R=5c=j=�j	=f=�\=FO=\<=HE�<�<w��<�=�<U��<�.�<���<]��<�V�<���<�=�<0��<=s�<�0�<2�<+�<�ݷ<[س<Kԯ<�˫<<��< ��<�s�<�>�<� �<n��<�v�</�<�<���<Y�z<sr<
ji<�`<X<�_O<�F<�><1�5<��,< u$<��<�V<��
<s�<���;���;���;BV�;��;;o��;��e;�;C;XD!;u ;�=�::0M:!\�7����xt�c븺����o���x;�%-[���z�y䌻�6��[A������mȻ��ֻ�Q�������z��ݭ��o����U(��)!���%�	�*��0/��3�	8��U<�s�@�:�D��qH��L��|O�՛R�rrU�NX�jUZ�(s\�pj^��J`�#b�d���e�q�g�� j�L^l�!�n��q�ms�K�u�#&x�zz���|�&�ȵ���ၼ!�� @���o��,���]ʇ�V����!���R�������Ӎ�~*��F���
��3����������v+��j����
��f[�����~�����������_���ޚ��=�������Ʀ����70���v��+ë����u_������V󰼐:��쁳�#˴�����c��v�������G�������  �  �WO=��N=�N=�iM=ֹL=KL=�BK=�|J=��I=.�H=�H=[SG=��F=��E=�6E=ęD= D=�C=2�B=��B=�B=��A=\A=0{@=h�?=AP?=�>=d>=�g==��<=�<=�y;=��:=�8:=ƙ9=��8=b[8=H�7=7=-�6=��5=TK5=��4=�4=�r3=��2=�2=�b1=w�0=�/=�/=�1.=]-=��,=�+=�*=�3*=!x)=��(=v
(=�Q'=2�&=��%=J�$=�$=�#=:�!=�� =�=T/=��=�L=I�=5(=�~=��=��=�'=�D=�V=�_=�b	=g`=�Y=GN=>==AJ�<��<���<5J�<���<#A�<���<j�<ls�<#��<�_�<���<��<�R�<*$�<��< ��<+�<T�<Bޫ<eʧ<㪣<�~�<G�<��<���<Xr�<N%�< ؅<q��<�wz<\�q<I1i<9�`<<�W<�2O<��F< �=<qr5<f�,<�u$<��<e<c�
<��<�/�;�.�;� �;���;�n�;8?�;�B�;,g;VbD;Lh";h.;;M�:�f�:��:�K�7�(�Or�dܷ�����R��1;�2[���z�X����\��j{��iK��p�Ȼ��ֻ����p��z����������%��!���%���*�9/��3���7�.<�8Y@�D`D��8H���K��:O�LWR��-U���W��Z��9\�N7^�H`���a�
�c�t�e�Z�g�!j��Nl��n�
q��ss���u��@x�/�z�J�|�HK�bЀ�����(���U�����t����ч��������#M��$����ȍ�v�����w����y��b��y���P��Ʉ���隼.9��r���F���~����������������� ���/����ꧼp)��9s���ë����~i����������Q�������崼z0���{��~Ÿ����Q��;����  �  DVO=,�N=�N=�oM=��L=L=�NK=p�J=��I=��H=�.H=�jG=߭F=g�E=�QE=�D=� D=ӖC=�C=o�B="B=ƕA=�A=��@=�?= V?=s�>=/>=Ke==��<=�<=)l;=��:=.%:=q�9=�8=�F8=ة7=�7=ru6=��5=SG5=�4=Q4=�w3=R�2=[$2=m1=��0=d�/==/=�D.=�r-=��,=��+=�+="N*=��)=��(=
 (=e'=��&=q�%=��$=P$=4#=��!=� =�=@-=�=C=��=�=�i=��=k�=@=-=B=�N=UU	=�V=�S=�K=�==QP�<�<���<c\�<>��<�\�<���<04�<���<U�<4��<�&�<���<{��<�U�<�4�<� �<��<X�<��<��<V��<S��<�Q�<�<���<qi�<+�<e��<,i�<�(z<"q<x�h<�,`<+�W<'�N<�UF<��=<vU5<��,<)t$<��<�w<��
<<Ȇ�;��;N�;)N�;O�;g�;��;�h;�/F;31$;~�;~�:kN�:��	:M�C8� ��n�W������%��I�:��Z���z����h���ޫ�Bʺ�U\ɻ��׻�[�'��E��������#��� ��%��!�`�%�Yq*���.��]3�H�7�V�;�W@�D���G��xK��N�3�Q���T��XW�v�Y�s�[���]�3�_�+�a���c��e�¿g���i�z:l�:�n��
q�_�s�V�u��mx�3�z��>}���s����&���P��}x��v���:����އ�n�������F��y��Ĺ���
��"m���ޑ��[��Cߔ�(c��&ᗼPS��>������=��b�� u���y��v���o��Sl��rr�����������ݧ�� ���o��:ƫ�~ ���z���ү�'���w���ų����Z�����m渼'���c�������  �  RRO=*�N=
N=�uM=P�L=�L=�[K=k�J=��I=7I=�HH=�G=��F=F=�sE=[�D=e@D=~�C=�,C=B�B=�(B=�A=!A=֎@=��?=z[?=�>=[>=g`==1�<=�<=Y;=V�:=�
:=�g9=�8=
+8=�7=��6=�d6=R�5=f@5=��4=u4=|3=�2={-2=�x1=��0=M�/=c*/=r\.=΍-=��,=��+=.1+=�o*=�)=��(=;(=u|'=I�&=��%=
%=�$=#=>�!=�� =o�=�(=�=05=��=��=�M=��=��=��=�=z&=T7=�B	=:I= K=>G=�<=~T�<v�<{��<Wp�<E��<M}�<���<=d�<;��<vQ�<��<�k�<�<o��<3��<Lm�<^R�<�>�<�,�< �<5��<ӣ<���<�[�<��<��<MZ�<���<���<�;�<��y<	q<�Zh<��_<TW<�N<�F<��=<�)5<r�,<�j$<�<w�<�
<+D<���;�;��;>�;���;���;�&�;�k;�|H;Uv&;	;��:��:PG:��8`�ع��j�C����i��)H�X~:�ιZ���z��R��*���h���w���%ʻ�hػ9�ʏ�+1 �,U��1�;�����,�h!���%��S*���.��-3�z7���;���?���C��rG�]�J��ON��cQ��9T�!�V��:Y��r[���]�q�_��{a�:tc��{e���g���i�	(l��n�dq��s��&v���x�`,{��}�w��5��-`������진��ą��܆���.��Q!�� B���n����������T��|����7��e���B1����������r��a��������!���9��E��H���H���K��|W��p��P���-ѧ�����n��.ͫ�^0��*�������
S��&��������J��5���ַ�E��"K��6~�������  �  @KO=f�N=�N=�yM=��L=< L=+hK=N�J=��I=t&I=�eH=ƨG=��F=BF=d�E=�D=�cD=c�C=�HC=��B=�;B=-�A=�(A=��@=�?=�^?=+�>=�	>=JX==�<=)�;=LA;=̓:=h�9=�E9=E�8=�	8=�r7=��6=P6=��5=65=��4=�4=�}3=��2=52=Ԃ1=&�0=a0=�?/=v.=��-=s�,=`,=5W+=ו*=��)=G)=�X(=ԕ'="�&=:�%=�%=�#$=,#=g "=�� =́=� =M�=#=݉=��=%,={j=��=�=��==�=A+	=M7=C>=/?=�8=ZS�<�!�<���<���<�<���<��<���<�<��<�"�<���<�`�<��<���<���<��<�k�<R�<6�<��<��<�<a�<r�<��<CD�<Gى<�m�<��<<y<6{p<�g<C"_<E�V<�N<ŝE<�?=<l�4<3�,<�U$<��<"�<	<�d<G�;���;��;�ν;�;��;X�;��m;�K;[);��;,��:y�:�&:`^�81	Ϲ �f�U���2� ��J:���Z�+{� ���儝�i���M���˻�oٻ�D�K���˥ ����V��=�4>��?�!��%�/=*�ʪ.��3��A7�)g;��k?�\IC�&�F��uJ�߻M���P���S��@V��X�-�Z��]��._��4a�v<c��Pe�Pzg���i�	l�\�n��'q���s�Gbv���x�d�{��~��G���z��6���~ǃ��ᄼW���-����u���)���B���h������掼�=��+������ˆ�������i��Ϙ��'��Ar��M���<ٝ�t����
��������+���=���\��Z����ȧ�"���s��Jګ�G�������!��,���X鲼UA������5׶����dJ��nx��Ӡ��vƼ��  �  �@O=*�N=:N=BzM=k�L=�&L='rK=I�J=��I=>I=R�H=�G=�G=oiF=n�E="E=��D=��C==dC=�B=MB=8�A=2A=l�@=�@=�^?=ɳ>=�>=�L==d�<=�;=�%;=zs:=`�9=V9=�~8=��7=tP7=��6=�76=��5=A(5=۞4=�4=O|3=[�2=]92=c�1=P�0=�0=�S/=4�.=��-=�-=A,=�~+=J�*=b�)=�:)=�v(=Ԯ'=��&=�&=� %=4*$=�#= "=�� =�z=K=��==+n=��=D=;A=�r=!�=��=��=��
=�	=�!=�-=q3=1=�J�<��<V��<��<�+�<��<|F�<���<�S�<���<�p�<'�<��<�c�<$!�<(�<���<疴<�s�<xO�<%�<w�<���<o_�<�<���<�&�<l��<�8�<IĀ<��x<q�o<�#g<�^<3�U<��M<�(E<�<<q�4<[m,<2$<��<��<<�y<Ő�;9 �;=Q�;t��;�Ԭ;R&�;���;Np;��M;��+;�
;A��:l�:��:�q�8Qƹ�;c��ӱ��^���"K:�U[�r�{�����#��㭻�A���,̻�ڻ`n�4���k)�5+���jI��q�!`�J!�ٸ%�N4*�^�.���2��7�G';��?�n�B��~F���I��"M�u)P�>�R���U�8$X�q|Z���\�#�^���`��c��0e�;gg�t�i��#l�o�n��Iq���s�-�v��^y�|�W�~�^����ǁ���1���#��{-���0���0���1���8��9J���i�����1ێ�,���������Z���ĕ��)��3���Lڙ�9"��&^��~���ﳞ�GП�6格J���&��)���N��؂��ǧ����0��~e��,ޮ�oU���Ʊ�:/������޵��"���[���������ʻ��弼�  �  �2O=b�N=�N=�vM=!�L=�)L=�xK='�J=WJ=SSI=�H=��G=G:G=^�F=�E=�GE=��D=@D=�}C=�B=�[B=�A=�7A=��@=� @=�Z?=��>=��==�===�<=��;=F;=}Q:=Ԡ9=��8=�V8=ѽ7=�,7=D�6=�6=�5=w5=v�4=U4=w3=�2=:2=C�1=�0= "0=>e/=�.=��-=�%-=Me,=��+=V�*=� *=�[)=�(=��'=��&=�&=�'%=�,$=#=��!=�� =�o=d=?�=e�=;P=��=��=v=�F=�p=��=��=J�
=i�=.	=K=]$=�%=M;�<��<���<��<�9�<j��<jj�<V��<|��<?#�<Q��<�Z�<� �<Z��<�d�<�$�<�<C��<,��<�a�<�/�<f��<{��<DV�<]�<��<��<��< �<��<x<�9o<{f<��]<&XU<c�L<�D<�v<<aO4<U+,<� $<%�<�t<�<��<��;�U�;���;aC�;��;�2�;eÊ;��r;$nP;�H.;�r;���:���:�$:S9s9����`������X��L�:���[��y|�����֞�&��� C���Kͻ�ۻK�黤���n�����E������׍�">!���%�h:*���.���2���6�K�:���>���B��F��dI�яL��O��dR��U�ȝW�kZ��W\�)�^�o�`���b�$e��bg�2�i�f7l�/�n��yq��8t�� w�p�y�w�|��,�Iހ����eA���[��fh���i���b���X��RP���N��Y��ar�������׎��!��Jw��?Ԓ�4������햼�B������ ՚�����F���s��ڙ�������ء�W���<��mH��ł���̧��'������	���������.������/x���ڴ�,.���q��O���$˹��庼d���D
���  �  7#O=�N=�N=vpM=Y�L=�(L=�{K=}�J=�J=�dI=�H=rH=�YG=v�F=�F=CiE=��D=-D=x�C=q�B=�fB=]�A=�9A='�@=p�?=�S?=Ӣ>=��==_-==Cl<=��;=��:=)0:=z|9=x�8= 08=v�7=�	7=�6=�6=r�5=!5=��4=�3=�n3=X�2=572=��1=]�0=�*0=s/=_�.=s�-=�B-=��,=��+=�+=A*=�x)=��(=��'=��&=�&=5+%=-,$=�#=~�!=N� =3b=��=]r=�=H2={=��=Y�==[F=�m=��=B�
=��=�=|=T= =�%�<�<��<Ñ�<AA�<"��<m��<�$�<.��<4`�<���<5��<qG�<!��<נ�<oW�<��<ڴ<��<�l�<�2�<��<��<�F�<Pۖ<b�<�ݍ<S�<�Ƅ<�>�<�w<՛n<��e<K9]<O�T<�gL<�.D<%<<�3<��+<Y�#<�<�S<��
<�y<l��;���;�7�;e׿;�w�;��;(Ӌ;�)u;��R;�0;K�;h��:Kۖ:� ):#{9���_L_��ǰ��#�E��u�:�U&\��Z}�:5��������@���bλ��ܻ������:������S��J��3���g!���%�N*�+�.�;�2�O�6���:��>��5B��E���H��L��O��Q�ގT��&W� �Y�?\��W^�q�`�{�b�ge�zlg�|�i��Wl���n�߱q�D�t��Xw�Q1z���|�>���(���d�����-���ϫ��D�������悈�:r���i���m��=������#ێ�`���k��.�������h��K���u���L��A���b͛����5;���j�����ྡ��碼`�� I������l٧��9��ѩ���'��0����:��Ű�%H�����j&��[{��e����츼.�����a)���1���  �  dO=�N=�M=4hM=x�L=�%L=�{K=��J=G J=lrI=(�H=H=tG=��F=�(F=A�E=�D=�BD=��C=�C=�nB=��A=09A=[�@=�?=�J?=��>=Q�==�==�X<=V�;=;�:=G:='\9=��8=8=\w7=��6=�f6=��5=4n5=?�4=u4=��3=�d3=��2=22=��1=��0=y00=P}/=[�.=.=cZ-=q�,=W�+="+=�[*=v�)=>�(=��'=�'= &=�+%=)$=�#=��!=ϫ =!T=��=C^=l�=�=%\=|�=	�=|�=� =�I=�p=��
=ʹ=��=q�=R=�	=x�<���<S��<��<|C�<���<$��<E�<���<]��<'8�<P��<G��<v(�<���<)��<�4�<��<ȯ�<Bq�<j0�<��<n��<4�<;Ö<�C�<���<�&�<˒�<s�<��v<^n<OIe<o�\<�7T<p�K<5�C<��;<��3<&�+<��#<�g<-<��
<_j<���;-��;���;�I�;��;J�;���;?w;�T;��2;�g;���:�p�:�-:˘!9;ɶ�Y�^��ް�Z��!N�;���\�GB~�ď�u:��Fe���$���[ϻ[�ݻ��������Ɗ�6��C��:������!�q&��i*�&�.���2���6���:��l>���A��WE��H�~�K�p�N�YeQ�!T���V��QY�]�[��+^���`���b�5"e�cg�>�i��}l�L'o��q�K�t�H�w�ǒz��m}����aj�������у�>愼4腼Yۆ��ć����ޓ��o���B���S���w���^㎼R ��f��ذ������;G��Ď��Fӗ�<��pU��l����ќ�	��;E��z��g���Xޢ�%���N��㔦�n駼/N��Kê��F��Wԭ��f�����Ձ��D���:i������ ���,���F���R��0V���W���  �  �O=��N=T�M=7`M=a�L=�!L=�zK=}�J=�%J=�{I=_�H=�,H=y�G=��F=�>F=&�E=��D=�RD=�C=KC='sB=��A=E7A=�@=��?=TB?=��>=f�==�==PH<=x�;=غ:=��9=�B9=�8=@�7=B]7=?�6=iP6=��5=�\5=I�4=;h4=��3=�[3=u�2=�,2=k�1=l�0=k30=�/=��.=g .=�k-=e�,=��+=P7+=�o*=	�)=��(='�'='=�"&=+%=@%$==#=�!=V� =�G=+�=�M=-�=� =�C=�{=��=#�=�=H-=]V=o~
=�=��=��=��=u� =^��<���<���<���<�B�<1��<���<�[�<�
�<���<+b�<{	�<D��<�Q�<���<���<�J�<.��<���<�q�<M+�<�ޣ<���<F"�<���<�)�<ř�<�<�h�<2�<��v<��m<��d<<\<��S<�K<8dC<�Y;<q\3<_+<]W#<Y<<4	<��
<�X<1��;���;=��;��;���;�q�;�\�;��x;DV;=�3;@�;N2�:*O�:�/: �(9;�����^��%��["�r��T<�ρ]�5��;��Ƞ��������� лp�޻M��-���~�����Z�6��t��-��!�%0&�"�*��.�k�2�k�6�s�:��P>�y�A�!E��FH�WNK�":N��Q�R�S��|V�Y��[�G^��s`�j�b�Z-e��g��j�{�l��Qo�ur�u���w���z�l�}��I��N���ނ�����������>뇼̈�V�������ݘ�����������쎼�$���d��t����쓼Y/���o������똼F*���i������라�)���f�������٢����U����������Ja���٪�.a��@�֊��:!������K0��֝��A���J5���^���t��H|���z��w���  �  ��N=�xN=��M=yZM=οL=�L=yK=�J=�(J=)�I=B�H=�6H=`�G=��F=�KF=��E=E=a\D=k�C=+C=�uB=��A=s5A=n�@=��?=]<?=��>=>�==n==l=<=t;=��:=X�9=N29= �8=%�7=�L7=}�6=�A6=��5=>Q5=7�4=�_4=q�3=&U3=�2=�(2=͆1=��0=�40=��/=�.=�(.=�v-=��,=�,=lD+=7|*=ɬ)=3�(=V�'=�'=�#&=�)%=4"$=�	#=��!=� =^?=y�=rB=~�=��=�3=pj=[�=v�=�=C=lE=�n
=�=#�=��=^�=� =
��<���<���<�< A�<z��<��<�i�<R�<r��<�{�<�$�<U��<�j�<��<R��<�W�<��<¹�<�p�<�&�<�֣<}�<y�<O��<��<Ȅ�<��<6M�<�j<�Rv<m\m<�d<��[<s�S<lGK<E*C<&;<�.3<?7+<�4#<�<]�<�
<�K<���;���;���;���;�ʯ;ʞ;9č;�hy;~.W;��4;�; ��:�k�:0u1:R�,9�4��آ^��k��4�����h<�{�]�G�������%���r���P���л�D߻�+�|J��P��	�a���� ��[O���!��H&���*���.���2���6�>�:��@>�̲A���D�%H��K��N�|�P�1�S��PV�I�X���[��]�sm`���b��6e�ѣg��"j�úl��oo��@r��(u�;x�{���}��h�����G ��!)��p:���6���"��A��7∼�É�H���)��������ʍ�
��(���d��*����㓼3!���\��]���\Ҙ�����O��n���S֝����[��G���0آ�t���[��y���?���n��k骼3s���������;��]Ͳ�GP��w�����
W����钺�W���В������  �  �N=�uN=�M=kXM=&�L=�L=xxK=+�J=�)J=�I=��H=Q:H=w�G=Y�F=RPF=G�E=zE=�_D=˺C=�C=IvB=��A=�4A= �@=��?=::?= �>=M�==#==�9<=�o;=.�:=�9=�,9==~8=3�7=�F7=�6=�<6={�5=DM5=��4=j\4=��3=�R3=�2='2=Ņ1=+�0=50=̈/=�.=�+.=Cz-=��,=
,=�H+=a�*={�)=�(=Q�'=�'=$&=j)%=!$=�#=��!=� =P<=�=�>=*�=��=X.=�d=.�=�=��=0=�?=�i
=w�=	�=G�=+�=Q� =a��<���<ί�<N}�<�@�<���<��<Pn�<�#�<w��<Ä�<�-�<\��<Is�<%�<ش�<�[�<�<#��<}o�<8$�<�ӣ<�x�<m�<^��<�<)}�<@�<�C�<]U<Q;v<�Cm<"xd<}�[<1qS<�1K<�C<�;<�3<*+<@)#<�<a�<�
<hG<t��;|��;��;c��;��;��;H�;��y;�|W;�,5;��;��:]Ĝ:|�1:h�-9���$�^� ������$�d�<��$^�z�������G������{��&�л	t߻s[�ux���e�|.	���������n[���!��Q&��*�U�.���2�*�6���:�<>���A�s�D�1H��K��M���P�.�S�UAV�u�X�1y[���]��k`���b��:e���g�]*j���l�izo��Lr��6u��-x��&{��~��s���ʁ�$���4���E��oA��q,������鈼=ʉ�?���i�������΍�����z*��7e��ꢒ���������V�������ɘ�����F��'���=ϝ�b��uW��W����ע����^������H��ys��謁�y��=������"E���ײ�P[�� ˵�d#���b��;���>����������o����  �  ��N=�xN=��M=yZM=οL=�L=yK=�J=�(J=)�I=B�H=�6H=`�G=��F=�KF=��E=E=a\D=k�C=+C=�uB=��A=s5A=n�@=��?=]<?=��>=>�==n==l=<=t;=��:=X�9=N29= �8=%�7=�L7=}�6=�A6=��5=>Q5=7�4=�_4=q�3=%U3=�2=�(2=͆1=��0=�40=��/=�.=�(.=�v-=��,=�,=kD+=6|*=ɬ)=3�(=V�'=�'=�#&=�)%=7"$=�	#=��!=� =j?=��=�B=��=��=�3=�j=��=��=^�=�=�E=\o
=��=��=}�=�=�� =^��<!��<���<R��<AB�<���<��<cj�<��<���<1|�<�$�<3��<pj�<S�<���<�V�<	�<���<ro�<P%�<�գ<�{�<A�<$��<��<̃�<��<L�<�i<�Qv<	\m<�d<Y�[<,�S<�HK<�+C<�';<�03<o9+<>7#<;!<��<��
<	N<���;Q��;���;E��;Jͯ;.̞;�ō;*jy;?.W;��4;��;���:j_�:�W1:�!,9󀴹�^�����®�A� t<��^�&�������*��w���T����л<H߻�.��L��Q�t	�&���������O�?�!�I&�Й*���.���2���6�U�:� A>�ڲA��D�.H��K��N���P�4�S��PV�K�X���[��]�tm`���b��6e�ѣg��"j�ĺl��oo��@r��(u�;x�{���}��h�����G ��!)��p:���6���"��A��7∼�É�H���)��������ʍ�
��(���d��*����㓼3!���\��]���\Ҙ�����O��n���S֝����[��G���0آ�t���[��y���?���n��k骼3s���������;��]Ͳ�GP��w�����
W����钺�W���В������  �  �O=��N=T�M=7`M=a�L=�!L=�zK=}�J=�%J=�{I=_�H=�,H=y�G=��F=�>F=&�E=��D=�RD=�C=KC='sB=��A=E7A=�@=��?=TB?=��>=f�==�==PH<=x�;=غ:=��9=�B9=�8=@�7=B]7=>�6=iP6=��5=�\5=I�4=;h4=��3=�[3=u�2=�,2=k�1=k�0=j30=�/=��.=f .=�k-=e�,=��+=O7+=�o*=	�)=��(='�'='=�"&=+%=F%$=E#=�!=h� =�G=K�=�M=c�=6=�C=�{= �=��=R=.=<W=f
=!�=��=�=,�=�� =���<N��<,��<���<�D�<+��<f��<a]�<��<a��<�b�<�	�<��<�P�<���<q��<GI�<^��<���<�o�<�(�<cܣ< ��<��<M��<�'�<ߗ�<c �<Og�<�<��v<ڡm<��d<�<\<�S<-�K<�fC<1];<@`3<Xc+<�[#<!A<<��
<�]<K��;��;Ҷ�;���;��;v�;]_�;2�x;�CV;��3;ܵ;��:e7�:��/:�'9K���S�^��O���M���p<���]�5 ��E��rѠ��������(л��޻����������G\�s��"u��.���!��0&���*�t�.���2���6���:��P>���A�7E��FH�dNK�,:N��Q�X�S��|V�Y��[�I^� t`�l�b�[-e��g��j�{�l��Qo�ur�u���w���z�l�}��I��N���ނ�����������>뇼̈�V�������ݘ�����������쎼�$���d��t����쓼Y/���o������똼F*���i������라�)���f�������٢����U����������Ja���٪�.a��@�֊��:!������K0��֝��A���J5���^���t��H|���z��w���  �  dO=�N=�M=4hM=x�L=�%L=�{K=��J=G J=lrI=(�H=H=tG=��F=�(F=A�E=�D=�BD=��C=�C=�nB=��A=09A=[�@=�?=�J?=��>=Q�==�==�X<=V�;=;�:=G:='\9=��8=8=\w7=��6=�f6=��5=4n5=?�4=u4=��3=�d3=��2=22=��1=��0=y00=O}/=[�.=.=bZ-=p�,=V�+="+=�[*=u�)=>�(=��'=�'= &=�+%= )$=�#=��!=� =DT=��=�^=��=S=�\=�=��=O�=�!=�J=/r=�
=G�==�="�==�=�<]��<���<7��<�F�<���<���<G�<���<���<�8�<s��<��<�'�<z��<^~�<�2�<g�<鬰<%n�<"-�<,�<
��<�0�<��<�@�<��<3$�<ؐ�<��<��v<Kn<BIe<h�\<�9T<`�K<�C<F�;<�3<"�+<#�#<�n<�3<��
< q<���;��;C��;AS�;v�;�;u��;�w;\�T;��2;�^;���:'O�:��,:�" 9E����_�~�����rm��;�~�\��_~�>ҏ��G���q��!0���eϻY�ݻ���������F��Q��E�<������!�9&�1j*���.���2���6��:��l>���A��WE�)�H���K��N�deQ�$!T���V��QY�a�[��+^���`���b�6"e�dg�?�i��}l�M'o��q�K�t�H�w�ǒz��m}����aj�������у�>愼4腼Yۆ��ć����ޓ��o���B���S���w���^㎼R ��f��ذ������;G��Ď��Fӗ�<��pU��l����ќ�	��;E��z��g���Xޢ�%���N��㔦�n駼/N��Kê��F��Wԭ��f�����Ձ��D���:i������ ���,���F���R��0V���W���  �  7#O=�N=�N=vpM=Y�L=�(L=�{K=}�J=�J=�dI=�H=rH=�YG=v�F=�F=CiE=��D=-D=x�C=q�B=�fB=]�A=�9A='�@=p�?=�S?=Ӣ>=��==_-==Cl<=��;=��:=)0:=z|9=x�8= 08=v�7=�	7=�6=�6=r�5=!5=��4=�3=�n3=X�2=572=��1=\�0=�*0=s/=^�.=r�-=�B-=��,=��+=�+=A*=�x)=��(=��'=��&=�&=;+%=7,$=�#=��!=m� =]b=��=�r=j�=�2=�{=@�=3�==�G=o=6�=�
=��=�=�=|=U=f*�<}�<L��<Օ�<
E�<���<l��<'�<&��<�a�<� �<`��<�F�<��<2��<<U�<��<�ִ<���<�h�<�.�<��<ߞ�<�B�<iז<t^�<`ڍ<-P�<�Ą<=�<a}w<��n<��e<{:]<��T<�kL<o3D<�<<��3<��+<>�#<7�<\<Z�
<8�<0��;X��;�D�;��;���;'�;�׋;.u;�R;�0;7�;p��:��:P�(:"�9���T�_�s��ho���;��K\�C}��F��-���Ȫ��QN��Doλ��ܻK��s���=�� �+��x��������h!���%��N*�ș.���2���6��:�X�>��5B��E���H��L�O�$�Q��T��&W�&�Y�D\��W^�t�`�}�b�ie�{lg�}�i��Wl���n��q�D�t��Xw�R1z���|�?���(���d�����-���ϫ��D�������悈�:r���i���m��=������#ێ�`���k��.�������h��K���u���L��A���b͛����5;���j�����ྡ��碼`�� I������l٧��9��ѩ���'��0����:��Ű�%H�����j&��[{��e����츼.�����a)���1���  �  �2O=b�N=�N=�vM=!�L=�)L=�xK='�J=WJ=SSI=�H=��G=G:G=^�F=�E=�GE=��D=@D=�}C=�B=�[B=�A=�7A=��@=� @=�Z?=��>=��==�===�<=��;=F;=}Q:=Ԡ9=��8=�V8=ѽ7=�,7=D�6=�6=�5=w5=u�4=T4=w3=�2=:2=B�1=�0="0==e/=�.=��-=�%-=Le,=��+=U�*=� *=�[)=�(=��'= �&=�&=�'%=�,$=*#=��!=�� =�o=�=��=��=�P=)�=��=j=�G=&r=	�=N�=&�
=p�=\=�=�&=K(=D@�<q�<���<���<�=�<;��<�m�<"��<���<�$�<2��<)[�<- �<,��<c�<7"�<�<���<?��<�]�<,+�<��<٧�<�Q�<�<t{�< �<L�<[��<�<>x<#8o<�zf<L�]<�ZU<f�L<N�D<1}<<�V4<�3,<z	$<a�<,~<�<��<���;f�;4��;P�;���;u:�;�Ȋ;��r;9mP;B.;�f;���:�r�:�#:�S9�U���ca�b���X� ���:�w�[�5�|�񴎻1螻�Ϯ�PR���YͻW�ۻ�����u��n���H�S�����v��s?!���%�C;*�n�.� �2�G�6���:��>��B�F��dI��L� �O��dR�U�ѝW�sZ��W\�.�^�r�`���b�&e��bg�4�i�g7l�/�n��yq��8t�� w�q�y�x�|��,�Iހ����eA���[��fh���i���b���X��RP���N��Y��ar�������׎��!��Jw��?Ԓ�4������햼�B������ ՚�����F���s��ڙ�������ء�W���<��mH��ł���̧��'������	���������.������/x���ڴ�,.���q��O���$˹��庼d���D
���  �  �@O=*�N=:N=BzM=k�L=�&L='rK=I�J=��I=>I=R�H=�G=�G=oiF=n�E="E=��D=��C==dC=�B=MB=8�A=2A=l�@=�@=�^?=ɳ>=�>=�L==d�<=�;=�%;=zs:=`�9=V9=�~8=��7=tP7=��6=�76=��5=A(5=۞4=�4=N|3=[�2=]92=b�1=O�0=�0=�S/=3�.=��-=�-=A,=�~+=H�*=a�)=�:)=�v(=Ԯ'=��&=�&=� %=@*$= #= "= � =�z=�=�=r=�n==�==7B=!t={�=��=a�=��
=	=�#= 0=�5=�3=P�<�$�<G��<ʒ�<�/�<���<�I�<���<�U�<P��<�q�<Z�<���<\b�<=�<��<߹�<E��<�o�<K�<b �<��<4��<�Z�<���<���<*#�<��<56�<(<ȧx<��o<�#g<m�^<��U< �M<�-E<��<<�4<�u,<-;$<8�<x�<�<`�<���; �;n`�;���;r߬;�.�;��;Sp;�M;í+;��	;Kl�:ȶ�:�r:�N�8�wǹ�c�!(����.��Ww:��2[�e�{�}-���6��Z���iQ��;̻��ڻ�y�����-��.����K��s��a�� !��%�15*��.�t�2��7��';�?���B��~F��I��"M��)P�N�R���U�A$X�x|Z���\�(�^���`��c��0e�=gg�u�i��#l�p�n��Iq���s�-�v��^y�|�W�~�^����ǁ���1���#��{-���0���0���1���8��9J���i�����1ێ�,���������Z���ĕ��)��3���Lڙ�9"��&^��~���ﳞ�GП�6格J���&��)���N��؂��ǧ����0��~e��,ޮ�oU���Ʊ�:/������޵��"���[���������ʻ��弼�  �  @KO=f�N=�N=�yM=��L=< L=+hK=N�J=��I=t&I=�eH=ƨG=��F=BF=d�E=�D=�cD=c�C=�HC=��B=�;B=-�A=�(A=��@=�?=�^?=+�>=�	>=JX==�<=)�;=LA;=̓:=h�9=�E9=E�8=�	8=�r7=��6=P6=��5=65=��4=�4=�}3=��2=52=Ԃ1=%�0=`0=�?/=v.=��-=r�,=_,=3W+=֕*=��)=F)=�X(=Օ'=$�&=>�%=�%=�#$==#= "=�� =��=!=��=m#=c�=_�=�,=nk=�=U�=t�=�=n=I-	={9=�@=�A=:;=PX�<u&�<\��<{��<N�<~��<� �<l��<;�<���<}#�<���<`�<��<��<��<��<Uh�<.N�<�1�<f�<X�<K��<�\�<�<q��<�@�<։<�j�<��<L9y<�yp< �g<�#_<��V<�N<�E<(F=<��4<[�,<l^$<<��<�<n<�X�;֢�;���;q۽;o�;��;H]�;��m;�K;�);Mu;q��:l��:��:)_�8�%й2g��`��Ԇ����t:���Z��S{�h�������)(��(]���'˻ |ٻ�O绫���ҩ �g��8����/@�2A�i!���%�
>*�y�.�y3�?B7��g;�l?��IC�P�F��uJ���M���P���S��@V��X�4�Z��]��._��4a�x<c��Pe�Qzg���i�
l�]�n��'q���s�Gbv���x�d�{��~��G���z��6���~ǃ��ᄼW���-����u���)���B���h������掼�=��+������ˆ�������i��Ϙ��'��Ar��M���<ٝ�t����
��������+���=���\��Z����ȧ�"���s��Jګ�G�������!��,���X鲼UA������5׶����dJ��nx��Ӡ��wƼ��  �  RRO=*�N=
N=�uM=P�L=�L=�[K=k�J=��I=7I=�HH=�G=��F=F=�sE=[�D=e@D=~�C=�,C=B�B=�(B=�A=!A=֎@=��?=z[?=�>=[>=g`==1�<=�<=Y;=V�:=�
:=�g9=�8=
+8=�7=��6=�d6=R�5=f@5=��4=t4=|3=�2={-2=x1=��0=L�/=b*/=q\.=͍-=��,=��+=,1+=�o*=�)=��(=;(=v|'=K�&=��%="
%=�$=##=U�!=�� =��=�(=X�=�5=,�=��=�N=q�=��=�==�'=�8=�D	=.K=M=fI=?=�X�<� �<���<jt�<�<���<���<�f�<4��<�R�<���<#l�<��<_��<���<k�<�O�<c;�<s)�</�</��<�Σ<֙�<�W�<
�<}��<W�<���<J��<�9�<+�y<�q<�Zh<��_<�W<{�N<jF<;�=<#05<��,<�r$<<�<��
<tL<���;�$�;
&�;��;T��; �;�+�;�!k;�{H;Rp&;�;�a�:�:��:�X�8��ٹk�<�Q����n���:�^�Z�&�z��c��b���w������'2ʻ�sػ�B�2���4 �>X�i4�b����_.��!���%�_T*�]�.�^.3�xz7��;�%�?��C��rG�z�J��ON��cQ�:T�,�V��:Y��r[�Ƈ]�u�_��{a�=tc��{e���g���i�
(l��n�dq��s��&v���x�`,{��}�w��5��-`������진��ą��܆���.��Q!�� B���n����������T��|����7��e���B1����������r��a��������!���9��E��H���H���K��|W��p��P���-ѧ�����n��.ͫ�^0��*�������
S��&��������J��5���ַ�E��"K��6~�������  �  DVO=,�N=�N=�oM=��L=L=�NK=p�J=��I=��H=�.H=�jG=߭F=g�E=�QE=�D=� D=ӖC=�C=o�B="B=ƕA=�A=��@=�?= V?=s�>=/>=Ke==��<=�<=)l;=��:=.%:=q�9=�8=�F8=ة7=�7=ru6=��5=SG5=�4=P4=�w3=R�2=Z$2=m1=��0=d�/=</=�D.=�r-=��,=��+=�+=!N*=��)=��(=
 (=e'=��&=u�%=��$=X$=@#=��!=)� =5�=o-=M�=kC=
�=/=rj=E�==�=4=�.=@C=P=�V	=�X=�U=�M=�?=�S�<��<]��<�_�<V��<Z_�<��<=6�<H��<y�<ڔ�<�&�<G��<���<aT�<3�<`�<�<w�<���<;ާ<���<<�N�<��<���<�f�<��<t��<�g�<�&z<~q<k�h<�-`<"�W<�N<�YF<>�=<�Z5<��,<�z$<�<�~<��
<�$<���;��;��;wW�;�#�;6�;��;��h;?/F;J,$;j�;�c�:�,�:��	:��=8q���o�����y
��s����:���Z�2�z��%�������꫻sպ�kfɻ��׻oc���+���i���������&��!�)�%��q*�2�.�K^3���7���;��@�@D���G��xK�0�N�A�Q���T��XW�}�Y�y�[���]�6�_�-�a���c��e�ÿg���i�{:l�:�n��
q�_�s�W�u��mx�3�z��>}���s����&���P��}x��v���:����އ�n�������F��y��Ĺ���
��"m���ޑ��[��Cߔ�(c��&ᗼPS��>������=��b�� u���y��v���o��Sl��rr�����������ݧ�� ���o��:ƫ�~ ���z���ү�'���w���ų����Z�����m渼'���c�������  �  �WO=��N=�N=�iM=ֹL=KL=�BK=�|J=��I=.�H=�H=[SG=��F=��E=�6E=ęD= D=�C=2�B=��B=�B=��A=\A=0{@=h�?=AP?=�>=d>=�g==��<=�<=�y;=��:=�8:=ƙ9=��8=b[8=H�7=7=-�6=��5=TK5=��4=�4=�r3=��2=�2=�b1=v�0=�/=�/=�1.=]-=��,=�+=�*=�3*=!x)=��(=u
(=�Q'=3�&=��%=N�$=�$=�#=G�!=�� =/�=u/=��=�L=��=�(=	=F�=a�=D(=GE=dW=�`=�c	=�a=�Z=�O=�>=�L�<C�<	��<�L�<���<C�<a��<��<�t�<���<`�<��<ڕ�<R�<6#�<X�<���<Y�<K�<ܫ<ȧ<���<�|�<�D�<��<ۻ�<sp�<�#�<�օ<a��<nvz<��q<?1i<�`<��W<�4O<m�F<I�=<<v5<��,<dz$<T�<�i<H�
<��<�8�;\7�;H�;���;Bt�;SC�;AE�;�g;�aD;�d";�';�:�:�N�:e:��7B��ar����y@��i��G;��[���z�Q����e�����RS����Ȼ��ֻV���!���@��%�����%���&�^ !�X�%���*��/�\�3���7�..<�\Y@�``D��8H���K��:O�VWR��-U���W��Z��9\�Q7^�J`���a��c�u�e�Z�g�"j��Nl��n�
q��ss���u��@x�/�z�J�|�HK�bЀ�����(���U�����t����ч��������#M��$����ȍ�v�����w����y��b��y���P��Ʉ���隼.9��r���F���~����������������� ���/����ꧼp)��9s���ë����~i����������Q�������崼z0���{��~Ÿ����Q��;����  �  dXO=7�N=sN=eM=	�L=o�K=�:K=�sJ=R�I=�H=FH=SDG=p�F=�E=�%E=��D=�C=CqC=��B=�vB=��A=�A=��@=�t@=��?=�K?=�>=L>=�h==�<=�"<=E�;=F�:=E:=�9=�9=h8=��7=]'7=�6=4�5=WM5=~�4=�4=Lo3=|�2=�2=�[1=%�0=v�/=��.=%.=	O-=b{,=��+=1�*=�"*=�g)=H�(=|�'=�E'=R�&=J�%=_�$= $=#=��!=�� =�=0=��=SR=��=3=��=Y�=A=7='S=�c=�j=fk	=�f=u]=�O===�F�<S�<���<�>�<w��<�/�<ܔ�<��<�W�<1��<8>�<>��<s�<o0�<��<��<�ܷ<j׳<>ӯ<�ʫ<��<Û�<Cr�<z=�<���<X��<�u�<5.�<c�<���<��z<r<ji<o�`<�X<�`O<l�F<a><(�5<��,<[w$<��<dY<��
<��<C��;E��;���;�Y�;��;>Ė;׻�;��e;�;C;�B!;" ;74�:Q�~:c/:�7���J�t�2��>����O�;�]8[�[�z��錻|;���E�����pȻՌֻ�T�u������e�����pp�T���(��)!�H�%�D�*�1/��3�)	8��U<���@�I�D��qH��L�}O�ڛR�wrU�QX�lUZ�*s\�qj^��J`�#b�d���e�q�g�� j�L^l�!�n��q�ms�K�u�#&x�zz���|�&�ȵ���ၼ!�� @���o��,���]ʇ�V����!���R�������Ӎ�~*��F���
��3����������v+��j����
��f[�����~�����������_���ޚ��=�������Ʀ����70���v��+ë����u_������V󰼐:��쁳�#˴�����c��v�������G�������  �  �EO=@�N=N�M=�LM=�L=��K=B*K=�iJ=@�I=f�H=�H=�]G=�F=��E=�HE=c�D=�D=ӀC=a�B="oB=��A=�`A=6�@=�D@=2�?= ?=�t>=��==P-==�<=.�;=?;=�:=9�9=�V9==�8=[8={n7=��6=P)6=L�5=G�4=fB4=O�3=a�2==F2=��1=��0=�0=(I/=hz.=g�-=#�,=�,=`2+=re*=�)=��(=�(=EK'=/�&=M�%=i�$=:�#=.�"=}�!=�� =��=�d=-=l�=S4=��=�=9v=�==�6=Z]=wy=��
=c�=��=�=��=p� =���<���<$��<#,�<���<�X�<���<�b�<��<�o�<'�<n��<�X�<)�<!�<�ϻ<㹷<�<I��<ȉ�<Sr�< S�<�*�<���<C<5��<�D�<w�<��<�z�<�iz<;�q<LGi<k�`<�X<g�O<��F<�e><;�5<Bd-<��$<g<��<�@<@�<���;��;t�;�5�;=X�;���;�;&o;"�L;�B+;�;
;���:�:�(:�-9�P��6{N������N�"}�^�0�?�O��n�|����ѕ�����8,���g��0Qϻ[�ܻ�����������R�.��������!���&��P+��/��-4�=s8���<���@��pD��H��K���N�ɨQ��eT���V��MY�[��]���_�>�a��d��Ff� �h���j�aDm�6�o� r���t�	�v�ey���{��.~�_I��|������ーp���H��}z��[���G�������X������.����Y���Ƒ��;��4���|0��������p��"���X����(��KF��PX��Nc���k��Pw����������ͦ�y ��(>������ϫ�����l������W��S������c괼7��ǃ��Rи�����e��鮼��  �  qEO=\�N=��M=�MM=T�L=��K=;,K=lJ=ݨI=k�H=>!H=�aG=�F=�E=�LE=��D=�D=��C=��B=rB=>�A=�bA=$�@=wF@=j�?=?=+u>=��==�,==�<=��;=�<;=!�:=�9=qS9=ٰ8="8=�k7=6�6=j'6=�5=��4=3B4=��3=�2=OG2=��1=z�0=�0=pK/=&}.=��-=��,=s,=n6+=�i*=M�)=��(=�(=�N'=F�&=��%=��$=�#=��"=��!=�� =)�=�d=�=q�=�2=^�=�=�r=]�= =�2=�Y=v=��
=
�=:�=�=�=1� =(��<���<��<�.�<N��<]�<���<�h�<��<�w�<q�<��<�a�<�$�<O��<#׻<���<��<���<���<�v�<pV�<f-�<���<5Ö< ��<�C�<���<2��<xu�<L]z<��q<�8i<&�`< X<]vO<��F<0^><��5<�`-<=�$<wg<��<VD<u�<%��;���;!*�;fM�;�s�;¯�;��;�fo;�-M;[�+;p�
;��:�:Z�):?09t꡹h�M��p��Q亙d���0�,�O�)�n���ە�����2?��~��miϻ7�ܻT0�������{��&W�@���4���!�G�&�&K+���/��%4��i8�h�<�7�@�obD��H�rpK���N���Q�jUT���V�_?Y��}[�ͦ]�v�_��a�@d�Af���h���j�)Cm�̰o�y"r�b�t�[w��ny�*�{��;~�(P��ۂ��ܵ���胼���(L���|��d���a������ W��F���/���$V��c�7��q����)������
��Dh�������󜼘 ���>��iQ��1]���f���r������4���rʦ�s����<��σ��BЫ����ro������u��Y��:���1񴼙=��㉷��ո�����h�������  �  0DO=��N=a�M=+PM=�L=�K=�1K=�rJ=�I=-�H=+H=�lG=��F=9F=YE=��D=\ D=-�C=GC=�zB=��A=&iA=e�@=�J@=ʳ?=l?=fv>=��==7+==��<=��;=L6;=)�:=�9=�I9=��8=�8=c7=��6=�!6=�5==�4=tA4=:�3=��2=@J2=ܖ1=N�0=~0=JR/=!�.=��-=��,=�,=)B+=�u*=k�)=��(=�(=�X'=3�&=ϼ%=:�$=��#=C #=�!= � =p�=�d=7=C�=�-=��=�=i=��=��=�'=�N=al=c�
=R�=6�=��=W�=� =��<���<2��<97�<���<j�<���<�z�<��<+��<�$�<��<�z�<=�<c�<k�< Է<4��<���<|��<s��<T_�<E4�<l �<�Ė<���<�>�<D��<鮅<�e�<�8z<q�q<�i<�x`<o�W<�SO<��F<�G><�5<�W-<Z�$<�i</�<�O<C�<���;�(�;�f�;A��;kĬ;2
�;w�;�5p;N;�^,;�N;%��:�o�:K,:�99���r(L�&����{㺮)�o�0���O�L�n�gՆ������ߤ�y������d�ϻ�Fݻow�J=��?��ص��e�X����[���!�u�&��:+�\�/��4��M8��m<�Xi@�O9D��G��@K�KpN�rfQ��%T�޲V�Y�Y[��]�U�_�=�a�b�c�1f�]{h���j��?m�	�o�-+r��t��w�Ԋy���{��`~��c��b���Ȃ�����s(���V�����������������R�������쎼�K������(������������L�KP������ۜ�1	���(���=��sK��*W���e��Zz������æ������9��	���lҫ��$��Vx���ʯ�����j��O������P�������丼},��"r������  �  �AO=M�N=�M=�SM=��L=��K=�9K=`|J=�I=��H=R:H=y}G= �F=RF=xlE=��D=^2D=��C=$C=��B=��A=�rA=�@=Q@={�?=w?=�w>=�==#(==!~<=O�;=k+;=�:=>�9=�99=��8=Y�7=U7=�6=:6=-{5=�4=�?4=��3=>�2=3N2=o�1=E�0=#0=�\/=�.=��-=��,=�",=�T+=؈*=�)=��(=�0(=xh'=��&=��%=!�$=� $=�#=��!=� =��=�c=G= =�%=��==[Y=Q�=��=o=�==�\=�s
=y�=�=�=8�=� =���<c��<(��<NC�<���<�}�<P�<ǖ�<�!�<���<�J�<x��<��<Uc�<O2�<W�<l�<�ڳ<�ů<L��<(��<�k�<f=�<��<#Ɩ<��<�5�<��<���<aL�<F�y<�bq<��h<r5`<G�W<�O<��F<�"><ݲ5<�G-<��$<vk<`�<N`<�<�
�;�t�;���;V�;�B�;闛;��;|q;�PO;+�-;?�;��:���:(�/:r]F9�A��6�I�ׯ��q����`0�!�O��o�;����3���-���ٳ�0»*л��ݻ��껈������S���~�5�����A�!��&��"+��/��3�P#8��<<�m0@�a�C��G���J��"N��Q�s�S�blV���X��[��T]� _���a���c��f��jh���j�a=m��o��:r���t�,>w���y��.|�ޝ~�ƃ��$���悼����>���g��r��������≼����L�����������<���������9��������h���Ϙ�|*��Pw��;���a䝼������B0���?���Q���i�������������5��-����֫��.������ޯ�[4��6���z׳�%��$p������7���A��l��������  �  ==O=��N=�M=�VM=(�L=��K=CK=��J=��I=%I=jMH=ԒG=+�F=�-F=�E=��D=1ID=��C=�$C=��B=,B=�}A=��@=�W@=:�?=A?=*x>=��==#==�u<=��;=�;=or:=k�9=�$9=��8=��7=cB7=�6=&6=fq5=��4=C<4=�3=�2=R2=>�1=�0=	-0=�h/=�.=��-=C-=�8,=l+=�*=��)=^)=�F(= |'='�&=�%=��$=
$=�#=��!=�� =B�=�a=R=��= =��=��=TD=E�=��=s�=�&=�G=�a
=�u=��=ڋ=�=�� =[��<��<H��<�P�<V��<���<�)�<��<J�<���<�z�<�!�<G��<ؓ�<�_�<�6�<��<i��<��<Rī<բ�<Yy�<�F�<Z
�<%Ŗ<�x�<�'�<�Ӊ<m~�<�)�<]�y<�q<@ph<�_<QW<y�N<�ZF<��=<�5<�.-<��$<ti<��<�p<��<�P�;���;
3�;���;��;�K�;�֊;!s;��P;�O/;�!;���:#8�:��4:��V9ZU����F�����A����T50�g�O�f:o�=,������2���|\��g�»�л�b޻���^6���2��
�1�����$�f���!���&��	+��r/�j�3���7� <���?���C�
9G���J�=�M�4�P�{S�"V���X���Z�]�`L_��a��c��f�?Zh�J�j��>m�\�o�dSr�W�t�qw���y�Vx|�4�~�=���`�����e7��]�����Ϡ�����牼:���G������ӎ��+�����Y����f��"Օ��?��N���}���F��v�������t۞�����x��:#���9���V���|��ȭ���ꧼH3������߫��<��
���\����U������� ���O��ՙ��Q߷�P ��W]��*����ϼ��  �  �6O=e�N=u�M=�XM=~�L=� L==LK=֓J=��I=-I=�bH=٪G=[�F=@IF=�E=�D=�bD=�C=&9C=�B=kB=ڈA=��@=�]@=�?=�?=�v>=��==�==�j<=�;=`
;=�\:=��9=�9="h8=K�7=�+7=.�6=��5=�d5=��4=�64=y�3=C�2=�T2=J�1=��0=70=�u/=ϯ.=��-=I-=MQ,=��+=��*=T�)=�))=b_(=�'=ۿ&=��%=C%=S$=7#=�"=I� =�=�]=�=Ǎ=I=y=��=�*=�q=�=��=e=�.=�K
=9c=�t=�=��=@� ==��<@��<���<�]�<��<���<�I�<���<�w�<��<ֱ�<�Z�<W�<���<��<�d�<�=�<M�<C��<�ګ<߳�<c��<�M�<��<���<�m�<��<���<�[�<���<�Ly<!�p<�h<q_<��V<4uN<wF<��=<J\5<�-<��$<�_<��<�|<�<���;�,�;ի�;1�;���;`�;ɵ�;��t;9�R;01;��;�!�:�*�:��9:�h9�#��4�C��`����ຆH��!0���O��o�Ut��얻��������yû��ѻ�&߻"F�0���b~��H�x��% �7���s�!�;w&�_�*�S/�s�3���7���;�G�?�AOC���F��*J�.PM�FP��S�_�U��*X�ڊZ�s�\�P_�Va�c��e��Mh��j�GGm���o�Gur�u���w�0Fz���|��P�Aြ��&>���b��D�������y��� ҈�����G���E�������ǎ����.x���ܒ��D��謕�O��-o���Ù�$��M��􀝼ժ���̟��頼����!���C���n������b槼�3��Ƌ��u뫼NP��붮�����~���۲��2�������˶� ���I��H���߲���㼼�  �  �-O=ǕN=��M=�XM=��L=�L=!TK=ӞJ=Q�I=&/I=xH=x�G=wG=�eF=9�E=�E=�}D=�C=�MC=�B='B="�A=��@=Xb@=�?=	?=�s>=��====�]<=�;=��:=�D:=�9=��8=�K8= �7=w7=�{6=�5=�U5=U�4=�.4=ږ3=i�2=�U2=��1=q�0=�?0=��/=G�.=��-=�2-=�j,=%�+=`�*=*=uE)=�x(=g�'=��&=��%=�%=f$= #=�"=�� =��=]W=R�=`�=�=�c=��=�=LS=Q�=A�=�=�=53
=/N=�c=�s=�|=�~ =���<p��<��<Yg�<�<"��<�h�<��<��<F�<���<���<�H�<��<u��<]��<�e�<R=�<q�<o�<���<���<�P�<	�<·�<�]�<'��<ǘ�<�3�<Ѐ<[�x<e/p<;�g<��^<�{V<=N<��E<�e=<�!5<[�,<1�$<N<��<�<L�<9��;G��;� �;��;�F�;�;k��;��v;��T;�$3;��;��:
-�:�>::y9dT���GA�p���M�(&��-0��*P��p��·��f������*���>CĻu`һ��߻�h������A��+� J�fS�'.�(�!��q&���*�X9/�q3���7��~;�HN?���B��mF��I���L�Q�O�i�R��FU�p�W�6<Z�R�\�R�^��0a���c���e�qIh��j�IXm�^�o�ɠr�ENu��w�Νz��5}�H�����,K���s���������������҇�/戼�������]G��"}������'��Rd���'#��/��� ▼{:��O����Ӛ�[��CJ���x������Ġ�硼�
��e3��(d������姼�8��P�������kh���֮��C������w���i��l���N��9B���x��9���fӻ������  �  �"O=�N=��M=dVM=)�L=[L=�YK=��J=��I=�?I=?�H=��G=�,G=��F=}�E=7E=<�D=��C=GaC=��B=�2B=��A=�A=�d@=��?=!?=)n>=6�==}==�N<=R�;=��:=�+:=�|9=��8=�.8=��7=>�6=hd6=��5=3E5=K�4=1%4=�3=e�2=T2=��1=,�0=�F0=݋/=�.=|.=�G-=�,=��+=,�*=�+*=`)=�(=�'='�&=&&=c%={!$=�#=�"=�� =��=�N=��=9q=#�=M=\�=��=�3=�m=נ=��=�=H
=�7=&Q=~d=q=�u =���<��<x��<�l�<�(�<9��<��<+,�<��<�x�<>"�<���<A��<�:�<���<{��<���<�Z�<�,�<��<#˧<���<�N�<	�<���<�I�<��<�u�<��<>��<rx<ɷo<7g<�^<�V<�M<�UE<=<0�4<�,<�u$<�3<3�<~<V<���;}��;p��;j<�;�;��;�}�;��x;��V;�	5;�;.��:$�:��C:0%�9��z�5?�Ɵ�V�ߺP)��\0��P���p�G7��v헻�[��Rn��Ż�=ӻ������zp��".�}��.J�"{�|w�LF���!�Qu&�v�*�7(/��S3��^7��E;�?�D�B��
F��NI��jL�`O��1R�2�T�:wW�:�Y��\\�g�^��a� qc�	�e�aNh���j��qm��p�Q�r��u�'Ix�_�z�p�}�����S���������_Ƅ�rم��憼������V��)���M���~���������QT��)������2^���������T��e����ۛ�m��EI�� x��+����̡�����'���]��$���ꧼ�A�����������Y����m���ܱ��D�����������<��2x�������Һ�����<���  �  >O=��N=\�M=.RM=W�L=$	L=q]K=��J=C�I=�MI=�H=��G='DG=֚F=�E=�OE=I�D=D=(rC=��B=\<B=��A=�A=�d@=<�?=j?=g>=��==!�<=)?<=ȃ;=��:=k:=b9=�8=�8=�u7=��6=fM6=�5=S45=��4=c4=ه3=��2=�P2=��1=��0=&K0=��/=��.=�.=�Z-=��,=��+=F+=�D*=�w)=��(=�'=#�&=P&=�%=M%$=�#=�"=�� =��=�D=��=a=�=�6=ދ=}�=�=�N=с=�=�= 
=�!=C>=�T=Ld=�k =��<&��<%��<an�<�0�<���<Ĝ�<�K�<��<3��<T�<��<=��<Dl�<�&�<M�<٪�<Is�<+>�<��<Ч<��<DI�<A��<>��<�3�<Iō<`R�<�ބ<�m�<�x<�Do<G�f<�^<�U<�=M<��D<��<<R�4<�v,<�J$<�<0�<�r<�<��;� �;1��;b��;Ά�;b�;�G�;Xyz;}�X;��6;�.;��:�:U�G:�k�9H�q���=�`f����ߺUM���0��Q��Dq�4���-u�������'����ŻcԻ�����5��І�*	����7�����d�"�݀&�Y�*��/��?3��=7�x;���>�QB�S�E���H�[L���N�%�Q�։T�;*W�J�Y��,\��^� a�ic���e�[h���j���m��Fp��s� �u�n�x�U{�N~��L����������W�������z�����G��a��1#���7���W��σ��Ż��t���I�����듼<=��G���ڗ�D#��7h��*����圼����S��@��������颼e���[��8�����tN������D(��ᠭ�e��Ԗ��0���x���ٴ��-���s��a���Eٹ���������6���  �  �O=�{N=?�M=MM=7�L=;L="_K=H�J=J=�XI=4�H=$H=�WG=��F=c	F=�dE=S�D=�D=�C=<�B=eCB=h�A=�A=\c@=��?=�?=�_>=�=="�<=�0<=�r;=]�:=��9=�J9=��8=6�7=�]7=>�6=�86=ɭ5=�$5=v�4=�4=X3=)�2=L2=�1=��0=�M0=6�/=K�.=�&.=�i-=��,=��+=0#+=�Y*=܋)=��(=:�'=�&=�&=�$%=O'$=�#=# "=b� =��=;=��=�R=��=�"=.u=��=j�=�3=�f=Õ=m�=��	=�=�,=F=X=�a =x��<շ�<X��<�l�<X5�<��<��<1e�<�<���<�}�<S/�<���<r��<�K�<��<)ĸ<��<�J�<-�<"ѧ<^��<OA�<��<]��<��<"��<�1�<Q��<;B�<N�w<��n<�3f<+�]<{5U<6�L<L�D<*~<<5_4<�B,<9 $<0�<��<�b<� <��;�%�;��;��;� �;���;U��;��{;��Y;/8;��;a�:ˆ�:+�J:�<�9.�k�Z�<��I��w!�τ��1��Q�k�q����(�2����̷�{�ƻ��Ի�u�_}ﻓ���$��p	�y����_��w���"���&�e�*�`/�43�$&7���:�,�>�B�miE���H�7�K�b�N��~Q�T@T�k�V��Y��\�(�^�;�`�hc�j�e��kh��k���m��pp� <s�1v���x�*�{��[~�{|��Ǽ���킼o���#���,��5/���.���/��7��]G��c��Y���)��������A������5ד��"���l������0����=��-�����������6��co��@����ߢ�e���\���������;\���Ȫ��>��#����<��2���16������0
���^��P����ڸ�����"���;���R���  �  O=�sN=��M="HM=�L=�L=�_K=�J=7J=�`I=��H=�H=;fG=p�F=fF=tE=��D=,D=��C=o�B=HB=��A=�A=aa@=��?=�?=�X>=��==�<=�$<=	e;=Ӧ:=��9=:89=c�8=��7=�J7=s�6=�(6=7�5=!5=��4=�4=�w3=!�2=�G2=N�1=��0=�N0=��/=B�.=N/.=�t-=ѷ,=r�+=�2+=�i*=̚)=��(=f�'=�'=�&=(%=�'$=>#=��!=� =��=~2=b�=�F=��=�=Bc=�=��=:=ZQ="�=�=��	=��==:=�M=ZY =p��<T��<���<Ij�<F7�<N��<ǻ�<�w�<�0�<���<ܜ�<P�</�<<��<\g�<	�<%ָ<ْ�<?R�<7�<Ч<���<�8�<0ߚ<�z�<5�<˓�<4�<���<��<*\w<p�n<D�e<�T]<��T<�L<�eD<ED<<%-4<�,<�#<��<��<sS<�<>!�;�;�;�I�;�R�;�Z�;�c�;�n�;2�|;[;C9;��;���:�:�/M:���9��g��l<�R���d�i��2[1���Q�6zr�Pc��uY������O��� ǻdջ����m��A�T�	����v
�	��q��h1"���&��*�!/��.3�)7���:��r>�3�A�43E��_H�2oK�CdN��AQ��	T���V��]Y�,�[��q^���`��jc���e��|h��k�t�m�'�p�qfs��?v�Uy���{�/�~����iぼ-���4��GF��pL��K���F��]D��H��9U��#n������Î�e���&>������fɓ�����T��o���Jۘ�����_������᝼*!��1_��S����٢����_��M���>���h��ت��Q��sҭ��V�� ڰ�zW���ʳ�40������sʷ�����^%��A��V��Di���  �  ��N=tnN=O�M=�DM=S�L=:L=a_K=J�J=<J=BeI=��H=�H=oG=�F=O#F=�}E=:�D=v3D=��C=��B=�JB=��A=UA=�_@=.�?=�?=T>=�==c�<= <=\;=ќ:=��9=},9=28=��7=�>7=�6=6=͕5=�5=u�4=x 4=�r3=��2=hD2=�1=��0=O0=��/=��.=�4.=�{-=�,=� ,=�<+=Cs*=�)=��(='�'=�'= &=�)%= ($=�#=��!=T� =6�=�,=��=�>=l�=H=�W=��=��=�=�C=t=ɡ=��	=��==22=G=�S =��<��<���<�g�<�7�<v �<���<��<T?�<��<���<Ld�<4�<���<	x�< +�<��<H��<GV�<�<=Χ<W��<�2�<�֚<p�<���<���<��<ą�<�	�<@,w<�]n<��e<v!]<жT<lL<�;D<�<<>4<[�+<��#<.�<�<>H<��<��;�G�;Xd�;�{�;���;��;໏;��};P�[;�9;#;���:E�:,�N:�g�9(ne��G<�ri��R�����3�1��DR���r��������{R��ä���{ǻ�ջ�k�+m�.����=���	�K�7&�s���
A"��&�$�*�g$/��,3��7��:�]>�s�A�E��:H��GK��<N�kQ�"�S��V��GY���[�pi^���`�}nc���e�0�h�-k�s�m��p���s��`v�n=y��|�D�~�޹�������,��6L��u\���`��&]���V��R���S���^���u��똍�)ǎ�����<��~���������E��M���pȘ��	��8L������ѝ�'��]U��啡��֢�$��Db��4������q���⪼T^��V᭼�g��n��l���᳼TH��L����ⷼ(���:���T��~g��gx���  �  v�N=~lN=��M=VCM=[�L=�L=L_K=��J=#J=�fI=�H=OH=/rG=`�F=�&F=ـE=:�D=�5D=��C=&�B=mKB=ѨA=(A=
_@=&�?=�?=TR>=�==#�<=p<=Y;=V�:=��9=m(9=�z8=P�7=�:7=�6=r6=��5=�5=�4=_�3=�p3=��2=<C2=:�1=D�0=#O0=�/=��.=<6.=�}-=��,=�,=�?+=�v*=�)=��(=i�'=�'=)!&=7*%=�'$=Y#=��!=�� =��=�*=/�=�;=J�=�=�S=c�=�=)=Y?=�o=��=��	=Z�==�/=�D=�Q =*��<���<��<cg�<^8�<��<3��<چ�<aD�<"��<���<Ak�<�<[��<�}�<w/�<C�<Z��<>W�<�<Aͧ<g��<0�<�Ӛ<l�<���<]�<j��<�~�<��<Xw<cLn<��e<�]<�T<B\L<�-D<+<<~4<Z�+<��#<��<��<�D<.�<� �;iL�;Rm�;���;���;���;�֏;��};��[;�%:;UX;�F�: /�:%�N:��9D�d��F<��x��A��k�}�1��cR�2�r���������Kn��{ø�I�ǻ��ջ���3�������L���	��"��/��
�+���F"�t�&�O�*��%/�&,3��7�e�:� V>�9�A��E�.H�::K� /N��Q���S�|�V��@Y�%�[�g^�+�`��oc��e���h��2k���m�W�p�"�s��kv�?Jy�u|��~��u��5��\T��6d���g��dc��
\���V���W��Wb���x��	����Ȏ����<���|��v��� ��A��[����������E�������̝����5R����բ�2��:c���������t���檼�b��c歼�m�����Rt���鳼�P��զ��뷼:���B��\[��m���}���  �  ��N=tnN=O�M=�DM=S�L=:L=a_K=J�J=<J=BeI=��H=�H=oG=�F=O#F=�}E=:�D=v3D=��C=��B=�JB=��A=UA=�_@=.�?=�?=T>=�==c�<= <=\;=ќ:=��9=},9=28=��7=�>7=�6=6=͕5=�5=u�4=x 4=�r3=��2=hD2=�1=��0=O0=��/=��.=�4.=�{-=�,=� ,=�<+=Cs*=�)=��(='�'=�'= &=�)%=($=�#=�!=Z� =>�=�,=��=�>=��=e=�W=ٜ=��=�=/D=mt="�=��	=$�=�=�2=�G=%T =��< ��<���<�h�<�8�<:�<7��<~��<�?�<^��<*��<Vd�<�<���<�w�<�*�<^�<���<~U�<=�<Wͧ<j��<�1�<�՚<=o�<���<���<�<;��<Q	�<�+w<�]n<��e<�!]<[�T<�lL<�<D<�<<�4<��+<w�#<�<d�<"J<��<�#�;K�;Gg�;M~�;���;���;꼏;��};�[;��9;� ;���:�ܩ:�yN:y4�9��e��f<��y��V�ຝ��ܢ1�MR���r�����à���U����~ǻ��ջ�m�&o������>�~�	����&���+��GA"�5�&�L�*��$/��,3�7��:�]>�}�A�&E��:H��GK��<N�nQ�$�S��V��GY���[�pi^���`�}nc���e�0�h�-k�s�m��p���s��`v�n=y��|�D�~�޹�������,��6L��u\���`��&]���V��R���S���^���u��똍�)ǎ�����<��~���������E��M���pȘ��	��8L������ѝ�'��]U��啡��֢�$��Db��4������q���⪼T^��V᭼�g��n��l���᳼TH��L����ⷼ(���:���T��~g��gx���  �  O=�sN=��M="HM=�L=�L=�_K=�J=7J=�`I=��H=�H=;fG=p�F=fF=tE=��D=,D=��C=o�B=HB=��A=�A=aa@=��?=�?=�X>=��==�<=�$<=	e;=Ӧ:=��9=:89=c�8=��7=�J7=s�6=�(6=7�5=!5=��4=�4=�w3=!�2=�G2=N�1=��0=�N0=��/=B�.=N/.=�t-=ѷ,=r�+=�2+=�i*=˚)=��(=f�'=�'=�&=(%=�'$=D#=��!=$� =�=�2=~�=�F=մ=�=�c=o�=�=�=�Q=��=��=��	=��=�=�:=�N=QZ =a��<>��<g��<l�<�8�<���<��<�x�<�1�<s��<3��<P�<��<ǳ�<�f�<�<�Ը<~��<�P�<��<GΧ<���<,7�<nݚ<�x�<�	�<_��<��<���<�<[w<ߏn<=�e<U]<�T<��L<�gD<�F<<�/4<�,<��#<b�<��<W<��<(�;*B�;�O�;�W�;�^�;�f�;�p�;�|;�[;z@9;��;���:�:�M:6!�9ah�z�<��q��`��"���k1�uR�*�r��j���`�����V��J&ǻiջ:㻰��p������	����K�������1"�X�&�d�*�>!/��.3�P7��:��r>�F�A�C3E��_H�;oK�JdN��AQ��	T��V��]Y�.�[��q^���`��jc���e��|h��k�u�m�'�p�qfs��?v�Uy���{�/�~����iぼ-���4��GF��pL��K���F��]D��H��9U��#n������Î�e���&>������fɓ�����T��o���Jۘ�����_������᝼*!��1_��S����٢����_��M���>���h��ت��Q��sҭ��V�� ڰ�zW���ʳ�40������sʷ�����^%��A��V��Di���  �  �O=�{N=?�M=MM=7�L=;L="_K=H�J=J=�XI=4�H=$H=�WG=��F=c	F=�dE=S�D=�D=�C=<�B=eCB=h�A=�A=\c@=��?=�?=�_>=�=="�<=�0<=�r;=]�:=��9=�J9=��8=6�7=�]7=>�6=�86=ɭ5=�$5=v�4=�4=X3=)�2=L2=�1=��0=�M0=6�/=K�.=�&.=�i-=��,=��+=/#+=�Y*=܋)=��(=:�'=�&=�&=�$%=U'$=�#=. "=r� =�=";=��=�R=��=#=�u=�=��=24=^g=��=`�=��	=�=*.=gG=]Y=Cc =6��<���<���<}o�<�7�<,��<��<�f�<P�<���<~�<o/�<Q��<̔�<�J�<��<�¸<*��<fH�<��<�Χ<؊�<�>�<g�<���<��<��<�/�<ݶ�<A�<åw<�n<�3f<�]<�6U<j�L<,�D<��<<<c4<#G,<%$<>�<�<h<�<�(�;�.�;�%�;��;o�;��;.�;*�{;:�Y;e+8;�~;���:sm�:�J:���9}�l�*2=��v���O�u��-1�8�Q��r�]��M�������Zշ�O�ƻ��Ի�{�ǂ�?���#���q	����C��Y��C���"�<�&���*��/�[43�[&7��:�N�>� B��iE���H�D�K�l�N��~Q�Z@T�o�V��Y��\�*�^�=�`� hc�k�e��kh��k���m��pp� <s�1v���x�*�{��[~�{|��Ǽ���킼o���#���,��5/���.���/��7��]G��c��Y���)��������A������5ד��"���l������0����=��-�����������6��co��@����ߢ�e���\���������;\���Ȫ��>��#����<��2���16������0
���^��P����ڸ�����"���;���R���  �  >O=��N=\�M=.RM=W�L=$	L=q]K=��J=C�I=�MI=�H=��G='DG=֚F=�E=�OE=I�D=D=(rC=��B=\<B=��A=�A=�d@=<�?=j?=g>=��==!�<=)?<=ȃ;=��:=k:=b9=�8=�8=�u7=��6=fM6=�5=S45=��4=c4=ه3=��2=�P2=��1=��0=%K0=��/=��.=�.=�Z-=��,=��+=F+=�D*=�w)=��(=�'=$�&=S&=�%=T%$=�#=�"=	� =Ә=E=#�=�a=j�=A7=V�=�==�O=��=�=9�=Y
=%#=�?=iV=�e=�m =k��<y��<^��<qq�<�3�<c��<��<�M�<���<?��<�T�<��<��<zk�<�%�<��<Ө�<�p�<�;�<��<ͧ<��<*F�<5��<S��<1�<�<;P�<�܄</l�<�x<�Co<;�f<�^<әU<[@M<S�D<��<<@�4<,|,<tP$<�<��<�x<�<f�;��;��;��;Ǎ�;dg�;{K�;�|z;҆X;�6;I&;��:�a�:z_G:Z��9{s��(>�S����.�Kj���0�h!Q�I`q�e�������)	��12����Ż�Ի"�ỡ���:��C��*,	�a��������e��"���&���*� /�P@3�>7��;���>�:QB�m�E���H�kL���N�/�Q�މT�A*W�N�Y��,\��^� a� ic���e�[h���j���m��Fp��s� �u�n�x�U{�N~��L����������W�������z�����G��a��1#���7���W��σ��Ż��t���I�����듼<=��G���ڗ�D#��7h��*����圼����S��@��������颼e���[��8�����tN������D(��ᠭ�e��Ԗ��0���x���ٴ��-���s��a���Eٹ���������6���  �  �"O=�N=��M=dVM=)�L=[L=�YK=��J=��I=�?I=?�H=��G=�,G=��F=}�E=7E=<�D=��C=GaC=��B=�2B=��A=�A=�d@=��?=!?=)n>=6�==}==�N<=Q�;=��:=�+:=�|9=��8=�.8=��7=>�6=hd6=��5=3E5=K�4=1%4=�3=e�2=T2=��1=,�0=�F0=܋/=�.={.=�G-=�,=��+=+�*=�+*=
`)=�(=��'=(�&=)&=g%=�!$=�#=�"=�� =�=O=��=~q={�=�M=�=J�=�4=�n=ܡ=�=M�=�
=R9=�R=>f=�r=�w =���<���<��<Bp�<�+�<��<���<E.�<���<�y�<�"�<���<��<�9�<t��<���<���<7X�<�)�<���<�ǧ<5��<�K�<���<A��<�F�<"ߍ<^s�<��<���<px<��o<*g<�^<�	V<�M<�YE<�=<��4< �,<@|$<�:<C�<�<<<��;���;f��;�E�;���;���;���;D�x;�V;�5;��;F��:~�:vBC:�d�9!�|���?�e���=ພI�}0��P�S�p��E��P���ch�� z��/ŻvGӻK��_���v���0����L��|��x�dG�l�!�	v&�
�*��(/�1T3�,_7�/F;�2?�i�B�F��NI��jL�#`O��1R�;�T�@wW�?�Y��\\�j�^��a�"qc�
�e�bNh���j��qm��p�R�r��u�'Ix�_�z�p�}�����S���������_Ƅ�rم��憼������V��)���M���~���������QT��)������2^���������T��e����ۛ�m��EI�� x��+����̡�����'���]��$���ꧼ�A�����������Y����m���ܱ��D�����������<��2x�������Һ�����<���  �  �-O=ǕN=��M=�XM=��L=�L=!TK=ӞJ=Q�I=&/I=xH=x�G=wG=�eF=9�E=�E=�}D=�C=�MC=�B='B="�A=��@=Xb@=�?=	?=�s>=��====�]<=�;=��:=�D:=�9=��8=�K8= �7=v7=�{6=�5=�U5=U�4=�.4=ٖ3=i�2=�U2=��1=q�0=�?0=��/=F�.=��-=�2-=�j,=$�+=_�*=*=tE)=�x(=g�'=��&=��%=�%=m$=,#=�"=�� =��=�W=��=��=^�=9d=�=o=T=;�=O�=P�=9=�4
=�O=�e=pu=�~=�� =���<F��<Ѩ�<�j�<X�<��<~k�<�	�<���<MG�<���<��<XH�<��<��<w��<�c�<�:�<g�<$�<6��<O��<M�<��<e��<�Z�<P��<M��<t1�<�΀<-�x<D.p<.�g<��^<�}V<YN<÷E<�j=<H'5<��,< �$<8U<��<S�<q<���;��;+,�;��;O�;%�;t��;n�v;9�T;r3;-�;l�:&	�:��>:��w9 2����A�|�����ບG�EO0��KP��&p�އ�u���Ħ�b���NNĻ[jһ�໽����������.��K��T�H/��!�Gr&���*��9/�wq3��7�8;�xN?���B��mF��I���L�_�O�t�R��FU�v�W�;<Z�W�\�U�^��0a���c���e�rIh��j�JXm�_�o�ɠr�ENu��w�Νz��5}�H�����,K���s���������������҇�/戼�������]G��"}������'��Rd���'#��/��� ▼{:��O����Ӛ�[��CJ���x������Ġ�硼�
��e3��(d������姼�8��P�������kh���֮��C������w���i��l���N��9B���x��9���fӻ������  �  �6O=e�N=u�M=�XM=~�L=� L==LK=֓J=��I=-I=�bH=٪G=[�F=@IF=�E=�D=�bD=�C=&9C=�B=kB=ڈA=��@=�]@=�?=�?=�v>=��==�==�j<=�;=`
;=�\:=��9=�9="h8=K�7=�+7=.�6=��5=�d5=��4=�64=x�3=C�2=�T2=I�1=��0=
70=�u/=ί.=��-=H-=MQ,=��+=��*=S�)=�))=a_(=�'=ܿ&=��%=G%=Z$=B#=�"=`� =$�=�]=H�=�=�=|y=�=�+=~r=Ү=��=�=0=RM
=�d=�v=Ă=��=� =���<���< ��<%a�<��<���<'L�<���</y�<��<���<�Z�<��<���<���<�b�<�;�<��<S��<g׫<���<�<J�<^�<l��<�j�<�<F��<�Y�<	��<�Jy<
�p<�h<r_<��V<4xN<cF<��=<�a5<�-<�$<�f<��<�<��<���;�8�;ζ�;�'�;P��;J�;���;`�t;z�R;+1;=�;��:;�:%`9:єf9����*YD�ٝ��}*��h�&B0�ZP��o��������^+�����g�û&�ѻZ/߻�M컓������J�i���!�k8���W�!��w&���*�{S/�і3�ѻ7��;�u�?�fOC���F��*J�?PM�FP��S�g�U��*X�ߊZ�w�\�S_�Va�Ěc��e��Mh��j�GGm���o�Gur�	u���w�1Fz���|��P�Aြ��'>���b��D�������y��� ҈�����G���E�������ǎ����.x���ܒ��D��謕�O��-o���Ù�$��M��􀝼ժ���̟��頼����!���C���n������b槼�3��Ƌ��u뫼NP��붮�����~���۲��2�������˶� ���I��H���߲���㼼�  �  ==O=��N=�M=�VM=(�L=��K=CK=��J=��I=%I=jMH=ԒG=+�F=�-F=�E=��D=1ID=��C=�$C=��B=,B=�}A=��@=�W@=:�?=A?=*x>=��==#==�u<=��;=�;=or:=k�9=�$9=��8=��7=cB7=�6=&6=fq5=��4=C<4=�3=�2=R2==�1=�0=-0=�h/=�.=��-=B-=�8,=l+=�*=��)=])=�F(= |'=(�&=�%=��$=
$=�#=��!=�� =]�=�a=�=٘=N=�=3�=�D=�=v�=\�=�'=I= c
=�v=	�=m�=��=M� =���<c��<���<T�</��<>��<,�<̻�<�K�<���<{�<�!�<���<��<|^�<�4�<��<��<�ݯ<x��<ӟ�<Bv�<|C�<O�<;<Gv�<6%�<�щ<�|�<k(�<z�y<�
q<5ph<��_<�RW<)�N<O^F<:�=<��5<g4-<��$<�o<5�<�v<!�<Y\�;���;�<�;��;��;�P�;0ڊ;W s;&�P;`K/;I;���:�:�E4:UKU9}���;G�����6����FR0���O��Uo�j9���������g����»��л�j޻+��<��k5������B%�a���!�B�&�J
+�_s/���3���7�7 <���?��C�$9G�J�M�M�@�P� {S�*V��X���Z�]�cL_��a��c��f�@Zh�K�j��>m�]�o�eSr�W�t�qw���y�Vx|�4�~�=���`�����e7��]�����Ϡ�����牼:���G������ӎ��+�����Y����f��"Օ��?��N���}���F��v�������t۞�����x��:#���9���V���|��ȭ���ꧼH3������߫��<��
���\����U������� ���O��ՙ��Q߷�P ��W]��*����ϼ��  �  �AO=M�N=�M=�SM=��L=��K=�9K=`|J=�I=��H=R:H=y}G= �F=RF=xlE=��D=^2D=��C=$C=��B=��A=�rA=�@=Q@={�?=w?=�w>=�==#(==!~<=O�;=k+;=�:=>�9=�99=��8=Y�7=U7=�6=:6=-{5=�4=�?4=��3==�2=3N2=n�1=E�0=#0=�\/=�.=��-=��,=�",=�T+=׈*=~�)=��(=�0(=yh'= �&=��%=%�$=� $=�#=��!=)� =ͩ=d=o=��=�%=�=e=�Y=ޤ=Y�=-=�>=�]=�t
=��=H�=T�=��=Q� =���<��<ʓ�<�E�<��<��<'�<R��<�"�<���<K�<���<ԡ�<�b�<M1�<��<��<�س<�ï<���<���<oi�<�:�<Q�<�Ö<�}�<�3�<��<��<BK�<��y<bq<��h<,6`<��W<�O<��F<x&><�5<QL-<h�$<�p<��<ze<��<R�;�}�;���;J�;{H�;>��;��;q;PO;q�-;d�;O��:?v�:�/:dCE9�ޘ� 
J��ܣ���⺪���w0�`�O�o����>��D7��-⳻�7»1л��ݻB��5��������A��d��������!���&�Y#+�q�/�J�3��#8��<<��0@�|�C���G���J��"N��Q�{�S�ilV���X��[��T]�#_���a���c��f��jh���j�b=m��o��:r���t�,>w���y��.|�ޝ~�ƃ��$���悼����>���g��r��������≼����L�����������<���������9��������h���Ϙ�|*��Pw��;���a䝼������B0���?���Q���i�������������5��-����֫��.������ޯ�[4��6���z׳�%��$p������7���A��l��������  �  0DO=��N=a�M=+PM=�L=�K=�1K=�rJ=�I=-�H=+H=�lG=��F=9F=YE=��D=\ D=-�C=GC=�zB=��A=&iA=e�@=�J@=ʳ?=l?=fv>=��==7+==��<=��;=L6;=)�:=�9=�I9=��8=�8=c7=��6=�!6=�5==�4=tA4=:�3=��2=@J2=ܖ1=M�0=~0=JR/=!�.=��-=��,=�,=)B+=�u*=j�)=��(=�(=�X'=3�&=м%=<�$=��#=I #=�!=� =��=�d=S=g�=�-=ޥ=�=pi=�=O�=(=�O=m= �
=�=�=��=H�=� =��<���<��<�8�<���<�k�<���<�{�<x�<Ǝ�<�$�<)��<�z�<�<�<��<w�<�ҷ<ؿ�<��<֙�<��<�]�<{2�<���<LÖ<&��<,=�<��<⭅<3e�<�7z<�q<�i<Cy`<z�W<~UO<��F<J><��5<�Z-<��$<pm<��<�S<֩<f��;%/�;5l�;,��;tȬ;C�;y�;�7p;�N;"\,;�I;/��:�]�:��+:GQ89�z��~dL��٤�ʜ�e:�$�0�j�O�8�n�݆�$���椻4��h���V�ϻAKݻB{껙@��������f�/��f���o�!�ԧ&�;+���/��4��M8��m<�qi@�b9D��G��@K�TpN�zfQ��%T��V�Y�
Y[��]�W�_�>�a�c�c�1f�^{h���j��?m�	�o�-+r��t��w�Ԋy���{��`~��c��b���Ȃ�����s(���V�����������������R�������쎼�K������(������������L�KP������ۜ�1	���(���=��sK��*W���e��Zz������æ������9��	���lҫ��$��Vx���ʯ�����j��O������P�������丼},��"r������  �  qEO=\�N=��M=�MM=T�L=��K=;,K=lJ=ݨI=k�H=>!H=�aG=�F=�E=�LE=��D=�D=��C=��B=rB=>�A=�bA=$�@=wF@=j�?=?=+u>=��==�,==�<=��;=�<;=!�:=�9=qS9=ٰ8="8=�k7=6�6=j'6=�5=��4=3B4=��3=�2=OG2=��1=z�0=�0=oK/=&}.=��-=��,=s,=m6+=�i*=M�)=��(=�(=�N'=F�&=��%=��$=!�#=��"=��!=�� =2�=�d=�=��=�2=|�==�r=��=\ =3=�Y=\v=�
=u�=��=\�=}�=�� =)��<���<��<�/�<(��<�]�<���<i�<���<�w�<��<��<�a�<s$�<���<�ֻ< ��<^��<П�<ʍ�<�u�<�U�<y,�<��<V<P��<�B�<S��<���<u�<�\z<I�q<�8i<j�`<�X<*wO<��F<v_><Y�5<~b-< �$<Pi<��<;F<O�<���;��;-�;�O�;�u�;X��;��;�go;�-M;��+;�
;Y
�:��:�):��/9�#��}�M�L���V$�@m�=�0���O�g�n��Ɔ��ޕ�"���[B������kϻ{�ܻO2껜���ȭ����W����`�����!�x�&�NK+���/��%4��i8�w�<�D�@�ybD��H�xpK���N���Q�mUT���V�a?Y��}[�Φ]�w�_��a�@d�Af���h���j�)Cm�̰o�y"r�b�t�[w��ny�*�{��;~�(P��ۂ��ܵ���胼���(L���|��d���a������ W��F���/���$V��c�7��q����)������
��Dh�������󜼘 ���>��iQ��1]���f���r������4���rʦ�s����<��σ��BЫ����ro������u��Y��:���1񴼙=��㉷��ո�����h�������  �  �4O=��N=��M=�8M=ȈL=��K=$K=$bJ=ߤI=��H=*H=�oG=H�F=1
F=�`E=i�D=� D=>�C=��B=#eB=�A=DA=��@=�@=?=k�>=l>>=��==�<=iK<=��;=H�:=GU:=��9=y9=tb8=n�7=�7=�p6=(�5=5%5=�~4=��3=[,3=Z~2=��1=�1=�U0=]�/=a�.=��-=;+-=�X,=��+=ղ*=�)=[)=@(=�n'=�&=g�%==�$=��#=�#=N"=3� =j�=��=�V=� =#�=�%=�=�=p=��=O	=�C=rs=a�=��	=��=��=��=��=Y��<���<M��<�d�<''�<)��<���<4,�<���<xk�<��<���<l�<j*�<v��<�ɿ<!��<ō�<�w�<�b�<�K�<1�<��<��<E��</��<�Q�<d�</ى<���<�Z�<�4z</�q<�.i<*�`<'X<�O<�)G<��><y>6<��-<m^%<p�<(n<��<�P<�Y�;���;ԁ�;#�;���;c&�;��;��w;��U;��4;÷;��:䷦:�N:;E�9u�/�k�(�&w����к;M��2&��D�kgc��ŀ�.���i>��ӕ��E���p[ȻI�ջ>�⻳h�ˤ��ҹ��j	�����*�_@��*���"���'�e,�=p0��4��8��<�/�@�uMD���G��	K�cN��Q�̺S�OV�A�X��([�Z]��_�i'b�e�d�7�f��Xi��k�GOn���p�URs���u� Nx�(�z��=}�������K��ȃ��U���.��(��Y`��!���؊����g���������A}���璼�U��VÕ�e-��r����陼x7���x��)����؞��������3���O��Fq������&ʦ�k��yD��-����ث�/(���x��dɯ�����h����������S��样���9������μ��  �  14O=��N=��M=9M=��L=��K=�K=�cJ=��I= �H=�,H=�rG=4�F=9F=�cE=n�D=�#D=�C=e�B=CgB=��A=�EA=ޱ@=�@=�?=��>=�>>=[�==w�<=�J<=d�;=��:=0S:=e�9=�9=�_8=�7=c7=�n6=��5=$$5=
~4=\�3=I,3=�~2=p�1=�1=/W0=Ɠ/=�.=��-=--=>[,=Y�+=ȵ*=�)=_)=�B(=�q'=�&=��%=/�$=*�#=E#=g"=�� =��=��=]V=T =;�=�$=.�=�=nm=�=X=�@=�p==m�	=��=O�=��=�=y��<���<��<�e�<)�<s��<s��<�/�<^��<�p�<0�<���<,r�<�0�<���<rϿ<���<���<|�<�f�<XO�<�3�<��<Y�<@��<c��<Q�<B�<׉<{��<�V�<�+z<��q<�#i<��`<�X<�O<�!G<h�><�96<>�-<M\%<��<o<��<CT<�b�;��;���;*�;���;�<�;��;H�w;9V;߿4;��;��:��:�pO:[i�9��-�(�JF���mк�=�*&���D��ic��ɀ�����I�� �������[mȻ��ջ���	yﻔ���t��qn	�����+�A@��(���"�щ'�Q	,�Zj0�_�4���8���<�ɛ@�BD���G�y�J�N���P�f�S��DV���X�� [��x]�S�_�m"b��d���f��Wi�$�k��Pn�>�p�`Vs���u��Ux���z�aG}�9�����CP�����꾄����*���a�������׊�5��f��������Kz��[䒼�Q������(�������㙼h1���r��J���9Ӟ�������</���L��~n��`���pȦ�>��D��t����٫��)��+{���̯����ym�������
���X��~�����z<������Qм��  �  �2O=/�N=g�M=~:M=ˋL=��K=R"K=RhJ=A�I=p�H=�3H=�zG=��F=F=ulE=,�D=�+D=��C=S�B=gmB=/�A=�IA=~�@=�@=ہ?="�>=�>>===��<=�G<=T�;=d�:=M:=��9=��8=�X8=��7=�7=Wi6=�5=� 5=�{4=:�3=A,3=�2=�1=-1=iZ0=ԗ/=��.=�.=4-=�b,=Y�+=D�*=��)=)=rK(=�y'=L�&=�%=��$=�$=#=W"=� =&�=�=�U=��=L�=s =ך=3=f=�=��=p8=�h=a�=�	=T�=�=��=?�=���<��<��<�i�<�.�<���<�<;�<d��<^�<�$�<���<B��<�B�<G�<-�<��<���<{��<8q�<bX�<K;�<��<f�<|��<���<�N�<��<�ω<͍�<K�<	z<�q<�i<��`<��W<��O<G<�><H,6<'�-< X%<^�<_r<��<t^<�~�;&&�;���;PH�;Nگ;�~�;[B�;bx;P�V;1Y5;�;}'�:|�:�?Q:Q��9+�'�\�&��ʑ�к@�&�w�D�yc��ڀ�ď��m��iЬ�5亻o�Ȼ�ֻ����k���x��{	���_/�n?��$��"�]'���+�xY0�4�4�^�8��<��}@��!D��G���J�r�M��P�ĎS��&V�2�X�5	[��d]���_�b��ud�i�f��Si���k��Tn���p��cs�Q�u�]kx���z�Sc}����,&��^��x���eɄ�Z����0��Pe��.���]׊����6b��Z�������q���ْ�tE��谕����-z��^ҙ����+a��[���`Þ��矼���$��)C���f��E����æ�9����B���[ܫ��.������I֯�,)���z���ʳ�����f��첷�[���MF��/����ռ��  �  �/O= �N=��M=U<M=��L=g�K=�'K=ToJ=��I=2�H=�>H=�G=��F=�#F=vzE=��D=�8D=��C=*
C=�vB=6�A=�PA=ܺ@=�!@=��?=��>=?>=Y�==��<=�B<=��;=��:=C:=p�9= �8=�L8=��7=e7=)`6=��5=5=�w4=�3=�+3=k�2=b�1=�1=1_0=�/=M�.=O.=5>-=
n,=�+=��*=��)=�))=�X(=B�'=��&=�%=G�$=�$=�#=�"=� =��=6�=gT=��=c�=�=.�=��=Z=�=f�=�*=�[=��=��	=��=P�=��=�=���<ŵ�<���<.o�<�6�<��<��<]L�<���<���<J>�<���<���<^_�<(�<i��<ջ<.��<&��<R��<�e�<F�<� �<���<���<Ј�<~J�<Q�<�É<�}�<{7�<%�y<BYq<�h<�N`<�W<�WO<w�F<�{><�6<�-<�O%<h�<iv<m�<n<��;�\�;*��;��;�6�;L�;��;7Oy;�W;�I6;h;u��:꠩:hT:�y�9D��� %�q��ϺR��f�%���D���c�m�����,������47����Ȼ�aֻc�����!�����	���I6�=@�����"��o'�{�+�*@0��y4���8�x�<�-O@�Q�C��_G�ΡJ�T�M��P�l[S���U�txX�l�Z�F]���_�)b�sfd���f�VOi�G�k�p\n���p�sys�^v�\�x�{�ݐ}�t���=��xt�������ڄ���;���k��W���q׊����\��=������yd��'ʒ��2������� ��5`���������sE���|��r����П������4��[��"���C���A���{A������T᫼O7������毼)<��J���	⳼[1��C~���ȷ����jV�������޼��  �  �+O=�N=��M=>M=J�L=j�K=�.K=�wJ=�I=tI=�LH=��G=��F=�5F=]�E=r�D=�ID=��C=�C=��B=�A=�XA=#�@=a&@=��?=	�>=�>>=ה==��<=�;<=d�;=�:=�5:=��9=a�8=�<8=P�7=g�6=�S6=G�5=5=2r4=��3=G*3=��2=��1=�1=�d0=�/=Q�.=:.=�J-=�|,=۬+=��*=B*=;)=�i(="�'=�&=��%=��$=�$=y#=�"=-� =�=ɛ=�Q=��=p�=D=Y�=��=GJ=�=�==�J=�s=��	=��=��=��=I�=w��<u��<ޛ�<u�<M@�<b��<b��<b�<��<M��<_�<��<$��<ԃ�<iK�<��<e�<&ѷ<h��<ה�<�u�<�R�<�)�<B��<�Ú<B��<yC�<k��<���<�g�<3�<}�y<xq<�h<?`<\�W<�O<��F<�R><��5<0�-<eB%<��<Cy<i<�<��;��;zQ�;���;���;�i�;�B�;�~z;��X;�}7;ڏ;P�:��:>�W:�|�9[l�m#��=����κ��A�%���D���c�7&��2�������{������8rɻ�ֻ��ud���S���	��� B�D���O�"��^'���+�"0�NT4��d8�.P<�5@�|�C�NG�'ZJ��mM�WP�MS���U��CX�m�Z�� ]���_��a�Vd���f�8Li���k�9in�$ q�L�s�y.v�пx�IJ{�>�}��#��]��,����Ã��%��nI���u��Τ���؊����1W��Y���W����T��Ŷ����������▼3?������ߚ�"���Z�����������٠�����#��fM���}��>���x��� A��c���髼�C�����������U��㬲�� ���P��8����巼{*��hl��7���n뼼�  �  &O=ÆN=��M=�>M= �L=5�K=v5K=��J= �I=�I=�\H=+�G=��F=�IF=��E=n�D=k\D=@�C='C=��B=��A=.aA=��@=�*@=�?=v�>=�<>=�==��<=�2<=�;=��:=�%:=z9=��8=*8= �7=z�6=�D6=��5= 	5=�j4=��3=�'3={�2=�1="1=)j0=��/=��.="#.=Y-=Č,=�+=�*=T *=�O)=)}(=$�'=.�&=��%=�
%=�$=Z#=D"=�� =��='�=N=��=w�=�=�w=��==7=j�=:�=�="6=�`=��	=��=S�=��=��=`��<ư�<~��<�y�<�I�<4�< ��<�y�<a(�<���<V��<�6�<���<h��<�s�<'A�<a�<��<�˳<���<$��<�^�<2�<N��<WÚ<Z��<N9�<��<q��<M�<f��<�_y</�p<?h<3�_<FW<T�N<yF<!><<�5<$�-<�/%<��<Ox<#<�<P�;H��;R��;�k�;�.�;?��;g�;��{;1Z;[�8;$�;St�:gɭ:.Z[:�9��
��� �kj���Qκ�����%��E��d�?a��Ђ��|b����+����ɻ�i׻<b����;���C�o�	��,��S�FL���k�"�gO'���+��0�k,4��38��<���?��cC�w�F�pJ��M��P�b�R��yU�
X�K�Z���\��e_�.�a�KGd���f�#Mi�)�k��{n��q�B�s��_v�n�x�7�{��~��I�����׵��;䃼\���5���[��Ђ�������܊�d���R�� ���쏼XD��ۡ��6���b���������Bl��%�������4��;g����������硼)��I?���s��&���J���C��}�������S��ܴ�����ct��dϲ��%���v��+¶�g���I��1�����������  �  �O=�N=%�M=�>M=�L=
�K=�;K=.�J="�I=� I=�lH=l�G=�
G=�^F=�E=GE=pD=�C=�6C=��B=AB=iA=�@=.@=t�?=��>=�9>=��==��<=�(<=�u;=��:=�:=pf9=-�8=S8=r7=��6=;46=d�5=Z�4=�a4=P�3=�#3=�~2=��1={$1=�n0=[�/=$�.=�..=cg-=�,=��+=>+=E5*={d)=S�(=ú'=��&=��%= %=�#$=�%#=
"=<� =��=%�=�H=��=�w=#�=�g=�=A"=�n=�=��=�=L=Zr	=��=��=(�=��=[��<q��<Ț�<�|�<Q�<��<-��<���<�E�<.��<���<�`�<��<���<q��<h�<O8�<�<��<���<d��<ui�<:8�<! �<i��<�y�<!,�<�ٍ<Ʉ�<�.�<�ـ<y<�up< �g< f_<�V<E�N<6F</�=<J�5<�\-<�%<��<�r<�<��<�;�;(�;��;���;�;)��;*��;�D};<�[;�L:;d>;f��:b�:�?_:j��9� ���������ͺ {���%�+PE��wd�b�������P՟�<y��#�����ʻ�ػ[��~u��p��|y�h�	�gN��j�Z�� ���"��C'�ɤ+���/� 4�08���;���?��C�CyF�#�I�{�L�u�O���R�5U���W�zVZ�u�\��H_�ʿa�u<d��f�/Si���k�;�n�m?q���s���v�&<y�L�{�ze~��r������H݂�l��(.���P��9q��	���!���㊼p���P��ה��[ᏼ5�������蓼*D��h������B������rϛ����MB��t��Ţ��vС������2���k�����_����G��y������f��Zͮ�r3����������6N��O����궼�.���l��h���ۻ�����  �  �O=|N=n�M=�<M=T�L=��K=t@K=��J= �I=2-I=�{H=��G=8G=sF=��E=�%E=�D=!�C=AEC=¨B=�B=�oA=x�@=80@=`�?=��>=�5>=9�==��<=<=�g;=s�:=I:=@R9=�8= 8=S]7=l�6=�"6==�5=��4=�W4=ļ3=|3=�{2=v�1=�%1=�q0=�/=S�.=�9.=�t-=d�,=��+=�+=�I*=�x)=�(=��'=��&=&= %=R+$=�*#=�"=r� =��=ے=B=��=.l=��=�V=x�=�=�W=�=��=�=�6=�^	=��=��=��=��=��<���<N��<�|�<4V�<A$�<8��<���<fa�<'�<x��<<��<ZD�<�<��<���<�Y�<n)�<���<�ϯ<'��<tq�<�;�<��<�<=o�<��<ō<8j�<��<㴀<	�x<Hp<
�g<�_<��V<a?N<��E<ҫ=<lo5<e5-<�$<��<�g<�<��<@`�;�b�;�W�;wF�;�6�;~/�;87�;��~;�];Ȳ;;�;,k�:�1�:�b:��9J��0&��#����ͺ�{��&�h�E��d����� F��/O�����WX���=˻��ػj��
�)���]��;/
�t�Ն��l��*��"��='�ߕ+���/���3���7���;��L?�,�B�w)F�`I�<sL�_eO��9R���T�:�W��)Z�'�\��0_�R�a��6d�!�f�V^i��l�H�n�Ffq��t�*�v� �y��#|�˷~�~���ց�����-���O��m������W����ŉ��늼#��)Q�����'ُ��'��W{��(ѓ�K'���{��J͗�w��c��g����䜼���U��ƈ��⻡�Q�:(���e��Ϊ��L���~N��謪����{���箼�R����������w���ʵ�����V��ߐ��Lź�����m%���  �  �O=NuN=��M=7:M=��L=��K=�CK=x�J=��I=:8I=[�H=��G=�/G=��F=��E=�7E=0�D=e�C=<RC=6�B=�B=FuA=e�@=1@=-�?=g�>=�0>=~==��<=u<=�Y;=h�:=V�9=�>9=Ԓ8=��7=xI7=ū6=�6=qz5=!�4=hM4=��3=l3=�w2=V�1=u%1=�s0=-�/=�/=�B.=��-=��,=��+=�)+=-\*=b�)=��(=��'=��&=�&=t)%=�1$=I.#=�"=w� =��=��=�:=�=O`=t�=F=��=��=�A=H�=��=��=
"=7L	=1q=y�=��=;�=5��<��<���<�z�<�X�< ,�<p��<Z��<�y�<�6�<_��<��<�j�<z)�<���<N��<w�<:B�<��<(ޯ<���<�v�<m<�<���<Y��<3c�<"�<���<�O�<_�<��<3ox<d�o<!7g<_�^<�KV<[�M<��E<�p=<==5<�-<�$<q�<�X<�<��<xy�;���;"��;���;C��;��;�͐;�;�Y^;��<;��;��:��:�f:ş�9�H޸\���č�Iͺʏ��O&�!�E�ohe��I�������Ơ�"����뽻��˻xHٻY4滫��ny����T_
���$����9���"�d<'���+�i�/���3�J�7�t;��?�ŋB�J�E��I��'L��O�	�Q�/�T�efW��Z���\��_�p�a�16d���f�jmi��l���n���q�7Ot�Hw��y��m|���*ƀ������,��9R��2p��7���j���p���iԉ������ ��T��ݏ���ӏ����,l��ϼ������]��H�������Y=��3�����������j9��$r��r����㢼� ���b��᫦�W���eW��蹪�F#���������jq��Rݱ��B�������=���|�� ���g亼����;���  �  [O=�nN=��M=�6M=�L=�K=FK=��J=�I=AI=v�H=��G=4>G="�F=x�E=9GE=i�D=�C=�\C=��B=�B=yA=�@=�0@=1�?=��>=J+>=w==�<=�<=`M;=�:=��9=�-9=�8=��7=	87=T�6=�6=m5=��4=�C4=�3=e3=;s2=��1=^$1=�t0=��/=�/=+J.=1�-==�,=U,=I8+=�k*=��)=S�(=a�'=E	'=!&=|0%=36$=�0#="=�� =$�=V�=�3=#�=bU={�=7=�=��=X.=do= �=�=�=�;	=gb=��=۞=J�=؀�<F��<Ĉ�<Lw�<�Y�<#1�<[ �<S��<���<O�<u�<���<��<�I�<c	�<*��<w��<HV�<�< �<O��<�x�<;�<���<<1W�<=��<���<�7�<1ӄ<Sq�<�)x<ʀo<��f<�l^<�V<j�M<�nE<�:=<�5<��,<��$<�<�H<��<��<L��;��;w��;���;��;�%�;K�;{�;lo_;]>;�;�k�:ǭ�:�h:6��9S�Ҹ����ۈͺU���&��MF��e�E�������1����n��/a̻G�ٻ�滗�D������
����Y��G���H� �"�J?'��+��/���3�)�7��L;���>� UB�#�E�`�H�d�K��N�޿Q��T��>W�~�Y��~\�;_��a��9d���f�~i�J1l���n��q�{|t�Bw�`�y��|�L��逼3"��8O��0r��)���¢��,���aʈ��≼���t(��QX��Ӑ���Џ�����`����������D��#���uט����b��G���o䝼�"���_��ݜ���ڢ���b��Ů��l���`���ƪ��3���������񌰼
���7d��3ô�n��d`��s���ӹ�J ���(��P���  �  k�N=+iN=r�M=�3M=,�L=��K=3GK=��J=��I=yGI=��H=p�G=)IG=͠F=Y�E=�RE=�D=oD=�dC=��B=�B=o{A=��@=0@="�?=g�>=�&>=;q==��<=B�;=]C;=��:=��9=m 9=4s8=��7=a*7=d�6=��5=lb5=j�4=�;4=f�3=:3=;o2=��1=#1=�t0=��/=C
/=KO.=�-=��,=f,=kC+=Qw*=��)=s�(=o�'=�'=�'&=p5%=N9$=�1#=�"=�� =��=��=�-=��=�L=:�=M+=��=j�===�_=��=t�=�=�.	=�V=~y=�=�=�t�<��<=��<�s�<"Y�<#4�<9�<��<K��<>a�<�#�<#��<Q��<�a�<x �<��<f��<�d�<	*�<P�<;��<�y�<�8�<��<��<�L�<��<Z��<D$�<μ�<6X�<�w<6Go<��f<2^<��U<�{M<�>E<�=<	�4<��,<`�$<�r<O:<9�<;�<���;���;)��;;$�;�M�;�y�;��;���;g@`;��>;5�;���:�Զ:j:�p�9�A˸
k�����U�ͺF��/�&�S�F��Ff�5Ԃ�RQ��*����c���Ծ�0�̻s>ڻ�$绾|�GI���H���
�y���������W���"��C'���+�m�/�g�3��|7�G0;�W�>��+B��wE�إH�ȸK��N�j�Q� eT��!W���Y�[p\��
_��a�,>d���f�^�i�REl�!o���q�v�t��kw�l.z�F�|�������>��-j��u���&�������Ǉ�&و�����/���\�������Ϗ�R���X������锼a2���y��}������J��$����Н����R��I���բ�l��{b�����X	��ai���Ѫ�'A�������,��â��U��{~���޴�o3���{��츸��빼g��Q<���`���  �  ��N=geN=��M=�1M=̑L=3�K=�GK=�J=f�I=[KI=��H=b�G=�OG=��F=� F=�YE=��D=)D=biC=*�B=5!B=�|A=�@=\/@=��?=�>=�#>=Im==�<=��;=�<;=��:=�9=�9=]j8=��7=�!7=+�6=I�5=�[5=h�4=�64=�3=�	3=�l2=
�1=�!1=�t0=c�/=4/=[R.=M�-=�,=�,=AJ+=�~*=��)=F�(=��'='=�+&=g8%=;$=}2#=$"=N� =��=x�=�)=��=�F=��=�#=^~=^�=�=V=�=��=��
=k&	=TO=�r=k�=&�=m�<�|�<�}�<q�<eX�<�5�<X�<���<H��<_l�<�0�<p��<X��<�p�<�.�<���<A��<ym�<s0�<u��<���<�y�<�6�<�<���<�E�<��<{��<��<k��<'H�<Y�w<�"o<J�f<�^<�U<OZM<� E<}�<<C�4<�,<��$<�e<�0<	�<ס<(��;h��;��;�E�;�x�;C��;��;��;��`;T?;0 ;���:���:�k:��9�Ƹ�,�����ͺ!����&��F�|�f�����Ӂ��Y�����������ͻ��ڻQh绻��7����b���
�V��k�����a�}�"�[G'���+���/��3��o7��;�ܩ>��B��[E�z�H�Z�K��N��|Q�lOT�2W���Y��g\�	_�_�a�-Bd���f���i��Rl��o���q��t�w�oLz��}�������O��B{������β��)Ć�Ӈ��∼����x��T4��`��%���\Ϗ�����S���������#'���l��a���R���$<�������ĝ�����J�������Ѣ�Z��Rc������t��
o���ت�J��x���%9�������#��)���:�;E�������ɸ�6����$���H��uk���  �  M�N=dN=s�M=�0M=C�L=�K=�GK=��J=2�I=�LI=H�H=j�G=6RG=s�F=<F=O\E=��D=D=kC=O�B=�!B=7}A=;�@=/@=��?=9�>=i">=�k==K�<=��;=�:;=�:=;�9=�9=Sg8=�7=�7=K�6=��5=CY5=T�4=54=��3=o3=�k2=Q�1=}!1=~t0=��/=�/=IS.=��-=��,=�,=�L+=��*=7�)=��(=��'=�'=g-&=M9%=�;$=�2#="=�� =��=X='(=-�=�D=A�=2!=�{=C�=o=�R=��=��=��
=�#	=�L=�p=��=��={j�<�z�<f|�<ep�<~X�<�6�<��<���<}��<Dp�<B5�<c��<���<�u�<i3�<��<֯�<7p�<:2�<���<p��<Jy�<�5�<n�<|��<�B�<��<�|�<�<H��<mB�<�w<�o<�~f<9 ^<��U<�NM<HE<o�<<��4<%�,<4�$<�a<�-<%�<��<���;���;X�;hQ�;(��;J��;$��;]5�;j�`;	?;d(;���:�÷:�l:���9��Ÿ �ꃍ�"�ͺ��� '���F���f�g�������ҡ����(.��)ͻӛڻ>�绎��.���,l��
���"��߾�[e�3�"��H'���+�M�/���3�l7�;���>��	B�KRE�Y~H�/�K�L�N�$tQ�HT�<
W��Y�ye\��_�M�a��Cd���f�c�i��Wl��o���q�N�t��w��Vz�P}�������U��.���#���귅��Ȇ��և�戼�������6��Ha������1Ϗ����R��◓��ݔ�Q#��yh������C�07���{��g���k��H��狡��Т�����c������ �� q���۪�$M��ĭ�n=������<)������D���JK�������ϸ�� ��u)��0M��-o���  �  ��N=geN=��M=�1M=̑L=3�K=�GK=�J=f�I=[KI=��H=b�G=�OG=��F=� F=�YE=��D=)D=biC=*�B=5!B=�|A=�@=\/@=��?=�>=�#>=Im==�<=��;=�<;=��:=�9=�9=]j8=��7=�!7=+�6=I�5=�[5=h�4=�64=�3=�	3=�l2=
�1=�!1=�t0=c�/=4/=[R.=M�-=�,=�,=AJ+=�~*=��)=F�(=��'='=�+&=h8%=;$=2#=&"=R� =��=�=�)=��=�F=��=�#={~=��=�=EV=�=9�=�
=�&	=�O=Cs=ǐ=��=�m�<�}�<�~�<�q�<Y�<n6�<��<��<���<�l�<�0�<���<_��<�p�<v.�<���<㫼<m�<�/�<��<V��<�x�<6�<a�<��<�D�<P�<��< �<��<�G�<��w<P"o<H�f<%^<M�U<�ZM<e!E<r�<<]�4<��,<�$<Zg<#2<s�<8�<ɗ�;���;��;�G�;xz�;q��;��; �;��`;S?;L�;5��:���:�k:���9ƟǸbD�{�����ͺ����&���F�f�� ����������*�������ͻb�ڻ�i���b���[c�U�
����������a���"�|G'��+�ɣ/�#�3�p7��;��>��B��[E�~�H�]�K��N��|Q�mOT�3W���Y��g\�
_�_�a�-Bd���f���i��Rl��o���q��t�w�oLz��}�������O��B{������β��)Ć�Ӈ��∼����x��T4��`��%���\Ϗ�����S���������#'���l��a���R���$<�������ĝ�����J�������Ѣ�Z��Rc������t��
o���ت�J��x���%9�������#��)���:�;E�������ɸ�6����$���H��uk���  �  k�N=+iN=r�M=�3M=,�L=��K=3GK=��J=��I=yGI=��H=p�G=)IG=͠F=Y�E=�RE=�D=oD=�dC=��B=�B=o{A=��@=0@="�?=g�>=�&>=;q==��<=B�;=]C;=��:=��9=m 9=4s8=��7=a*7=d�6=��5=lb5=j�4=�;4=f�3=:3=;o2=��1=#1=�t0=��/=C
/=KO.=�-=��,=f,=kC+=Pw*=��)=s�(=o�'=�'=�'&=r5%=Q9$=�1#=�"=�� =��=��=�-=��=�L=`�={+=�=��=�=>`=�=��=N=7/	=YW=&z=Ŗ=��=Qv�<[��<���<"u�<wZ�<`5�<W�<���<��<�a�<$�<e��<`��<�a�<! �<���<���<�c�<)�<.�<��<yx�<�7�<o�<š�<�K�<��<K��<W#�<	��<�W�<N�w<�Fo<��f<~2^<W�U<�|M<�@E<{=<*�4<��,<�$<�u<=<��<�<Ŗ�;��;f��;�'�;�P�;�{�;���;��;@`;��>;��;7��:cǶ:8kj:�%�9I�̸:������$�ͺ�����&�ΨF��Rf�ڂ��V��H���:h��Aپ�
�̻�Aڻ�'�[�K��yI���
�'�������X���"��C'�ֆ+���/���3��|7�\0;�h�>��+B��wE��H�θK��N�n�Q�#eT��!W���Y�\p\��
_��a�->d���f�_�i�REl�!o���q�w�t��kw�l.z�F�|�������>��-j��u���&�������Ǉ�&و�����/���\�������Ϗ�R���X������锼a2���y��}������J��$����Н����R��I���բ�l��{b�����X	��ai���Ѫ�'A�������,��â��U��{~���޴�o3���{��츸��빼g��Q<���`���  �  [O=�nN=��M=�6M=�L=�K=FK=��J=�I=AI=v�H=��G=4>G="�F=x�E=9GE=i�D=�C=�\C=��B=�B=yA=�@=�0@=1�?=��>=J+>=w==�<=�<=`M;=�:=��9=�-9=�8=��7=	87=T�6=�6=m5=��4=�C4=�3=e3=;s2=��1=^$1=�t0=��/=�/=+J.=1�-==�,=U,=H8+=�k*=��)=S�(=a�'=F	'=!&=0%=66$=�0#="=�� =3�=j�=�3=E�=�U=��=]7=3�=�=�.=�o=��='�=�=z<	=Ec=��=՟=L�=��<Y��<ϊ�<Gy�<b[�<�2�<��<���<��<�O�<�<E��<"��<oI�<��<j��<v��<U�<��<e�<���<(w�<+9�<���<��<jU�<���<��<A6�<҄<{p�<�(x<1�o<��f<m^<V<�M<qE<�==<�5< �,<J�$<�<�L<�<��<|��;���;u��;��;,�;�(�;=M�;|�;�n_;�>;��;�\�:���:�h:22�9Y�Ը�6������ͺ4����&�h_F�5�e�{�������8���
��$t���f̻�ٻ.��I�r���� ���
����%����yI�p�"��?'�Q�+�$�/��3�N�7��L;���>�UB�2�E�k�H�m�K���N��Q��T��>W���Y��~\�<_��a��9d���f�~i�K1l���n��q�{|t�Bw�`�y��|�L��逼3"��8O��0r��)���¢��,���aʈ��≼���t(��QX��Ӑ���Џ�����`����������D��#���uט����b��G���o䝼�"���_��ݜ���ڢ���b��Ů��l���`���ƪ��3���������񌰼
���7d��3ô�n��d`��s���ӹ�J ���(��P���  �  �O=NuN=��M=7:M=��L=��K=�CK=x�J=��I=:8I=[�H=��G=�/G=��F=��E=�7E=0�D=e�C=<RC=6�B=�B=FuA=e�@=1@=-�?=g�>=�0>=~==��<=u<=�Y;=h�:=V�9=�>9=Ԓ8=��7=xI7=ū6=�6=qz5=!�4=hM4=��3=l3=�w2=V�1=u%1=�s0=-�/=�/=�B.=��-=��,=��+=�)+=-\*=b�)=��(=��'=��&=�&=v)%=�1$=P.#=�"=�� =��=ʍ=�:=D�=�`=��=\F=��=_�=6B=�=��=��=�"=3M	=Br=��=�=x�=���<���<x��<J}�<[�<$.�<`��<��<1{�<�7�<)��<���<�j�<:)�<5��<b��<�u�<�@�<��<1ܯ<���<Qt�<:�<H��<��<a�<
�<���<(N�<
�<��<�mx<��o<7g<�^<3MV<`�M<F�E<�s=<�@5<�-<y�$<�<�]<�<Y�<F��;���;y��;T��;y��;��;DА;r�;TY^;;�<;8�;��:D�:7�e:��9Ɗฦ*�#B�ͺ����e&��	F�m}e��S�����hϠ�J���I󽻁�˻dNٻ�9�2��S}������`
�I��������9�A�"��<'��+���/���3�x�7�Ct;��?�ۋB�\�E��I��'L��O��Q�5�T�ifW��Z���\��_�q�a�36d���f�kmi��l���n���q�7Ot�Iw��y��m|���*ƀ������,��9R��2p��7���j���p���iԉ������ ��T��ݏ���ӏ����,l��ϼ������]��H�������Y=��3�����������j9��$r��r����㢼� ���b��᫦�W���eW��蹪�F#���������jq��Rݱ��B�������=���|�� ���g亼����;���  �  �O=|N=n�M=�<M=T�L=��K=t@K=��J= �I=2-I=�{H=��G=8G=sF=��E=�%E=�D=!�C=AEC=¨B=�B=�oA=x�@=80@=`�?=��>=�5>=9�==��<=<=�g;=s�:=I:=@R9=�8= 8=S]7=l�6=�"6==�5=��4=�W4=ļ3={3=�{2=u�1=�%1=�q0=�/=R�.=�9.=�t-=c�,=��+=�+=�I*=�x)=�(=��'=��&=&=� %=W+$=�*#=�"=�� =��=��=@B=��=hl=�=�V=�=-=[X=��=��=�	=�7=
`	=ւ=�=ܶ=)�=Ԡ�<b��<��<��<�X�<�&�<a��<e��<�b�<e�<Z��<���<wD�<��<h��<���<&X�<�'�<��<^ͯ<ǟ�<�n�<9�<q��<g��<�l�<q�< Í<nh�<0�<���<v�x<xp<�g<�_<0�V<�AN<��E<c�=<�s5<�9-<��$<ٺ<�l<<ϩ<j�;�k�;�_�;�M�;^<�;�3�;:�;5�~;�];�;;݋;�V�:~�:.�b:"��9a�}��Q��{�ͺ+��2&���E��e�"���P��Y������`��HE˻��ػ8������7���0
�Su����m��+���"�>'�C�+���/���3���7���;��L?�E�B��)F�`I�HsL�ieO��9R���T�?�W��)Z�)�\��0_�T�a��6d�"�f�W^i��l�I�n�Ffq��t�*�v� �y��#|�̷~�~���ց�����-���O��m������W����ŉ��늼#��)Q�����'ُ��'��W{��(ѓ�K'���{��J͗�w��c��g����䜼���U��ƈ��⻡�Q�:(���e��Ϊ��L���~N��謪����{���箼�R����������w���ʵ�����V��ߐ��Lź�����m%���  �  �O=�N=%�M=�>M=�L=
�K=�;K=.�J="�I=� I=�lH=l�G=�
G=�^F=�E=GE=pD=�C=�6C=��B=AB=iA=�@=.@=t�?=��>=�9>=��==��<=�(<=�u;=��:=�:=pf9=-�8=S8=r7=��6=;46=d�5=Z�4=�a4=P�3=�#3=�~2=��1={$1=�n0=[�/=$�.=�..=bg-=�,=��+=>+=E5*={d)=S�(=ú'=��&=��%=%=�#$=�%#="=K� =�=@�=�H=��=x=n�=h=}�=�"=~o=��=[�=� =!M=|s	=ϓ=I�=��=T�=F��<_��<���<S�<�S�<F�<i��<���<WG�<w��<��<a�<�<���<�<�f�<�6�<O�<��<k��<<�f�<�5�<t��<ɽ�<w�<�)�<�׍<<3-�<�؀<fy<up<��g<�f_<��V<��N<9F<��=<��5<�a-<�%<��<x<<�<(F�;�1�;f�;���;���;���;+��;WG};��[;�H:;7;a��:W�:��^:_��9�i�h3�l⎺�κE��&�iE��d������됻�ߟ������Ǽ�8�ʻ�ػ^廸z�{u��g{�
��O�l��Z��!�y�"�ZD'�0�+�(�/�B4�e8��;���?��C�WyF�3�I���L��O��R�5U���W�~VZ�w�\��H_�̿a�v<d��f�/Si���k�<�n�m?q���s���v�&<y�L�{�ze~��r������H݂�l��(.���P��9q��	���!���㊼p���P��ה��[ᏼ5�������蓼*D��h������B������rϛ����MB��t��Ţ��vС������2���k�����_����G��y������f��Zͮ�r3����������6N��O����궼�.���l��h���ۻ�����  �  &O=ÆN=��M=�>M= �L=5�K=v5K=��J= �I=�I=�\H=+�G=��F=�IF=��E=n�D=k\D=@�C='C=��B=��A=.aA=��@=�*@=�?=v�>=�<>=�==��<=�2<=�;=��:=�%:=z9=��8=*8=�7=z�6=�D6=��5= 	5=�j4=��3=�'3=z�2=�1="1=(j0=��/=��.=!#.=Y-=Ì,=�+=�*=S *=�O)=)}(=$�'=/�&=��%=�
%=�$=a#=O"=�� =��=B�=3N=��=��=�=Qx=B�=�7=�=��=�=7=�a=�	=�=��= �=H�=2��<���<I��<�|�<&L�<��<I��<�{�<�)�<���<7��<E7�<���<!��<�r�< @�<�<*�<�ɳ<u��<Ã�<p\�<o/�<���<���<�~�<
7�<��<���<�K�<@��<�]y<_�p<�>h<�_<�GW<��N<|F<�$><X�5<��-<l4%<��<�}<j<9�<#�;e��;���;�r�;�4�;��;N�;[�{;u0Z;~�8;�;`�:E��:9[:$}�9���4!�����|�κ��n�%��0E��,d�tl��g���\l������R3��Iʻlp׻
h��������D� �	�K.��T�,M�r��"��O'���+�0��,4��38��<���?� dC���F��J��M��P�i�R��yU�
X�O�Z���\��e_�/�a�LGd���f�$Mi�*�k��{n��q�B�s��_v�n�x�7�{��~��I�����׵��;䃼\���5���[��Ђ�������܊�d���R�� ���쏼XD��ۡ��6���b���������Bl��%�������4��;g����������硼)��I?���s��&���J���C��}�������S��ܴ�����ct��dϲ��%���v��+¶�g���I��1�����������  �  �+O=�N=��M=>M=J�L=j�K=�.K=�wJ=�I=tI=�LH=��G=��F=�5F=]�E=r�D=�ID=��C=�C=��B=�A=�XA=#�@=a&@=��?=	�>=�>>=ה==��<=�;<=d�;=�:=�5:=��9=a�8=�<8=P�7=g�6=�S6=G�5=5=2r4=��3=F*3=��2=��1=�1=�d0=�/=P�.=9.=�J-=�|,=ڬ+=��*=A*=;)=�i(="�'=	�&=��%=��$=�$=�#=�"=:� =+�=�=R=�=��=�=��=�=�J=l�=�=�=TK=�t=��	=�=�=��=��=���<���<_��<tw�<�B�<��<R��<�c�<)�<k��<�_�<"�<=��<���<�J�<��<*�<�Ϸ<���<ߒ�<ys�<WP�<~'�<���<j��<��<qA�<���<!��<�f�<,�<�y<�q<�h<�`<��W<� O<��F<*V><]�5<G�-<�F%<G�<�}<$<7�<���;5��;�X�;,�;ర;�m�;gE�;Q�z;T�X;pz7;��;��:���:�HW:���9����Y#�g���Ϻ���* &�}E���c�C0��~;�����ڃ�� ����xɻ�ֻM���h�v�����%�	���C��D�]���"�H_'�A�+�V"0��T4��d8�RP<�R@���C�_G�5ZJ��mM�WP�TS���U��CX�p�Z�� ]���_��a�Vd���f�9Li���k�9in�$ q�L�s�z.v�ѿx�IJ{�>�}��#��]��,����Ã��%��nI���u��Τ���؊����1W��Y���W����T��Ŷ����������▼3?������ߚ�"���Z�����������٠�����#��fM���}��>���x��� A��c���髼�C�����������U��㬲�� ���P��8����巼{*��hl��7���n뼼�  �  �/O= �N=��M=U<M=��L=g�K=�'K=ToJ=��I=2�H=�>H=�G=��F=�#F=vzE=��D=�8D=��C=*
C=�vB=6�A=�PA=ܺ@=�!@=��?=��>=?>=Y�==��<=�B<=��;=��:=C:=p�9= �8=�L8=��7=e7=)`6=��5=5=�w4=�3=�+3=k�2=a�1=�1=1_0=�/=M�.=O.=5>-=
n,=�+=��*=��)=�))=�X(=B�'=��&=�%=I�$=�$=�#=�"=� =��=J�=�T=��=��=�=o�=�=wZ=��=��=�+=D\=>�=j�	=��==�=��=�=���<ط�<���<)q�<�8�<���<���<�M�<	��<���<�>�<���<Р�<*_�<�'�<���<Ի<�<���<��<d�<JD�<��<��<��<	��<�H�<��<g<�|�<�6�<��y<�Xq<�h<)O`<-�W<sYO<��F<(~><�6<h�-<BS%<.�<Fz<J�<�q<K��;gc�;+�;K��;�:�;��;?��;&Qy;��W;!G6;�b;���:ō�:J�S:��9� ��`%�H3��*�Ϻ/��J&�l�D�ިc����^���f���4 ��B=��`ɻ�fֻCg�u��%�����&�	����7��@�/ �8�"�*p'���+�e@0��y4�Ǒ8���<�DO@�c�C��_G�ڡJ�]�M���P�q[S���U�wxX�o�Z�F]���_�+b�tfd���f�WOi�G�k�p\n���p�sys�_v�\�x�{�ݐ}�t���=��xt�������ڄ���;���k��W���q׊����\��=������yd��'ʒ��2������� ��5`���������sE���|��r����П������4��[��"���C���A���{A������T᫼O7������毼)<��J���	⳼[1��C~���ȷ����jV�������޼��  �  �2O=/�N=g�M=~:M=ˋL=��K=R"K=RhJ=A�I=p�H=�3H=�zG=��F=F=ulE=,�D=�+D=��C=S�B=gmB=/�A=�IA=~�@=�@=ہ?="�>=�>>===��<=�G<=T�;=d�:=M:=��9=��8=�X8=��7=�7=Wi6=�5=� 5=�{4=:�3=@,3=�2=�1=,1=hZ0=ӗ/=��.=�.=4-=�b,=X�+=D�*=��)=)=rK(=�y'=L�&=�%=��$=�$=#=\"=� =0�=�=�U=��=j�=� =�=k=Kf=a�=H�=�8=
i=�=��	=��=��=l�=��=a��<Z��<X��<�j�<�/�<��<��<<�<6��<��<�$�<A��<Q��<�B�<��<�߿<T��<͟�<v��<p�<'W�<�9�<T�<�<,��<c��<�M�<v�<�Ή<��<xJ�<9z<��q<�i<�`<N X<ǃO<�G<��><h.6<��-<�Z%<	�<u<B�< a<��;�*�;ο�;�K�;Rݯ;뀞;�C�;ccx; �V;1W5;|;��:��:+Q::U�9I�(��'��⑺�$к�&��!&���D�,�c������ɏ��r��լ�}躻H�Ȼdֻ�㻁�ﻬ���n���{	�����/��?��$�m�"��'���+��Y0�V�4�x�8�(�<�~@��!D��G���J�x�M��P�ȎS��&V�5�X�7	[��d]���_�b��ud�j�f��Si���k��Tn���p��cs�Q�u�]kx���z�Sc}����,&��^��x���eɄ�Z����0��Pe��.���]׊����6b��Z�������q���ْ�tE��谕����-z��^ҙ����+a��[���`Þ��矼���$��)C���f��E����æ�9����B���[ܫ��.������I֯�,)���z���ʳ�����f��첷�[���MF��/����ռ��  �  14O=��N=��M=9M=��L=��K=�K=�cJ=��I= �H=�,H=�rG=4�F=9F=�cE=n�D=�#D=�C=e�B=CgB=��A=�EA=ޱ@=�@=�?=��>=�>>=[�==w�<=�J<=d�;=��:=0S:=e�9=�9=�_8=�7=c7=�n6=��5=$$5=
~4=\�3=I,3=�~2=p�1=�1=/W0=œ/=�.=��-=--=>[,=Y�+=ȵ*=�)=_)=�B(=�q'=�&=��%=0�$=+�#=G#=j"=�� =��=��=fV=` =K�=�$=F�=�=�m=F�=�=A=�p=�=��	=��=��=!�=s�=;��<V��<���<�f�<�)�<��<��<j0�<���<�p�<l�<���<4r�<�0�<u��<,Ͽ<B��<L��<�{�<�e�<�N�<O3�<K�<��<���<���<hP�<��<�։<��<�V�<;+z<Ƨq<�#i<��`<MX<��O<n"G<\�><;6<w�-<�]%<$�<}p<D�<�U<fe�;
�;+��;�;=��;'>�;���;��w;V;־4;��;}�:��:�_O:{B�9:�-�'(��R���zк�D��0&�o�D��oc��̀�����uL����������XoȻ��ջq��cz﻿������n	�G��&,�~@� )���"��'�l	,�oj0�p�4���8���<�қ@�BD���G�}�J�N���P�h�S��DV���X�� [��x]�S�_�n"b��d���f��Wi�$�k��Pn�>�p�`Vs���u��Ux���z�aG}�9�����CP�����꾄����*���a�������׊�5��f��������Kz��[䒼�Q������(�������㙼h1���r��J���9Ӟ�������</���L��~n��`���pȦ�>��D��t����٫��)��+{���̯����ym�������
���X��~�����z<������Qм��  �  I%O=}N=5�M=�&M=�wL=��K=�K=8YJ=m�I=K�H=�.H=�xG=��F=�F=[lE=��D=�%D=��C=��B=^VB=��A=t&A=��@=;�?=Q?=�>='
>=
c==[�<=�<=zf;=$�:=�:= h9=x�8=8=�k7=��6=O6=�o5=��4=�4=�m3=q�2=�2=U1=��0=�/=8/=^J.=w|-=c�,=��+=�+=�,*=�U)=O~(=Q�'=�&=�%=�%=H$=�&#='"=�!=�  =��=�=JX=x=ś=�'=ܥ=�=�z=q�=�=`=��=��
=��=&
=�!=�2=�==:��<���< p�<S�<�)�<���<���<�t�<�,�<s��<���<aX�< �<���<���<���<�o�<�T�<'<�<�$�<��<O�<SТ<���<4��<�S�<�!�<��<���<}�<_C�<�z<��q<�)i</�`<�DX<�O<:kG<�?<J�6<�<.<��%< t<�<ӓ<�<��;f �;���;���;E��;q�;�x�;ZF;��];U�<;�g;A]�:���:�r:x��97(���~5�V<��F�������(:��4X���u�򙉻���v*���������:�λW�ۻ�,�OL�� ����&��o�X���|�0H���#�hu(���,��1��B5�A9�j=���@��MD�.�G��J���M��P��S��&V���X�qA[��]��>`���b��Be�w�g�cYj�x�l�}o�=r�6�t��,w���y�\=|���~������߁����|Z������?ӆ�y���O������ڋ�y'��{���ԏ�Z4��엒������b��}Ŗ��"��py��\ǚ�����H���}��6����֠�* ��d*���W��8����¦�U���E�� ����ݫ��.������ӯ��%��Cw��lȳ����h������]��HQ�������꼼�  �  �$O=�|N=2�M='M=+xL=@�K=zK=`ZJ=ѡI=��H=�0H=�zG=��F=�F=�nE=��D=�'D=��C=_�B=�WB=�A=�'A=y�@=��?=�Q?=,�>=
>=�b==ֹ<=�<=Re;=ú:=n:=if9=��8=@8=	j7=��6=�6=�n5=��4=�4=am3=O�2=�2=zU1=[�0=L�/=A/=�K.=�}-=�,=��+=�+=�.*=X)=t�(=w�'=�&=��%=o%=�$=�'#=("=�!=Q ==�=֟=X=� =�=�&=\�=�=�x=`�=�=�]=k�=��
=��=�=h =�1=�<=b��<P��<rp�<�S�<'+�<���<ں�<_w�<�/�<��<���<�\�<~�<r��<9��<A��<�s�<)X�<m?�<�'�<a�<P�<�Ѣ<Ϭ�<���<�S�<@!�<��<���<�z�<f@�<�z<��q<�!i<t�`<c=X</�O<�dG<~�><p�6<�9.<�%<s<.<3�<�<T%�;��;b��;A��;퓲;Z��;1��;�k;,^;"#=;2�;��:�ڸ:Cs:��9p9��2��~����U�������':��7X��u���������4�����a���[�λ �ۻ�8軽V��� �N��)��p����9|�PF���#��q(���,��1��<5�c:9��=���@��DD�]�G�J�J���M�ٵP�xS�$ V�ɴX�H<[�ռ]�d;`��b��@e��g��Yj���l�so��r�)�t��2w�1�y�XD|��~�R���"ぼ� ��F]������Ԇ����qP�������ً�z&���y��ӏ�*2��B���{���b_���������u��Ú�9���D���y�������Ӡ�T���(���U����������� ���E��_����ޫ��/�������կ��(���z���˳�D���k��칷�e���S�����_켼�  �  Z#O=O|N=K�M=�'M=�yL=?�K=%K=�]J=ѥI=u�H=�5H=]�G=��F=HF=uE=U�D=�-D=<�C=w�B=^\B=��A=�*A=��@=��?=�R?=ɯ>=
>= b==0�<=h<=b;=ʶ:=�:=9a9=;�8=�8=�d7=�6=�6=k5=�4=�4=4l3=��2=72=uV1=��0=��/=/=O.=�-=̱,=�+=�
+=5*=w^)=؆(=��'=��&=<�%=$%=� $=4+#=�*"=�!=� =��=��=@W=J�=r�=8#=%�=�=s=I�=6=�W=P�=$�
=��=Q==0/=%;=���<��<pq�< V�<�.�<���<���<y�<m9�<���<˫�<�i�<�,�<���<��<n��<�<Pb�<tH�<(/�<��<Y��<�բ<B��<���<pS�<��<��<孉<�r�<P7�<��y<
�q<e
i<=�`<"'X<!�O<ySG<��><:�6<�1.<��%<vq<~	<T�<�<�8�;�!�;�;���;��;P��;��;��;�^;�=;��;Jq�:e��:ϕt:���9�@��~[��D~�hݼ�4]�����):��GX�Xv������(���V��9�������ϻ�ۻ:^��v�� ����0��t�(��Zz��A���#��h(���,�1�d+5��&9���<��@��+D�=�G�3�J���M�#�P�bS��V���X��-[��]�/2`�O�b��<e���g��Zj�+�l��o��r�>�t�YCw���y�uY|��~�>����큼.*��^e��ȟ���ن���/R��뒊��؋�$��v��9Ώ�,��������VU��~������Kh�����D���T8��n������Mʠ�1���M!��oP���������������E��Z����᫼=4������5ݯ�n1�������ֳ�Q'��gv��ķ�e���[��@������  �  � O=�zN=)�M=�(M=�{L=H�K=0K=�bJ=�I=��H=>H=d�G=��F=H)F=$E=E�D=n7D=�C=`�B=RcB=��A=�/A=ѓ@=��?=�T?=��>=�	>=q`==m�<=O	<=�\;=A�:=7:=�X9=��8=�8=5\7= �6=�6=&e5=Z�4=�4=!j3=�2=w2=�W1=C�0=��/=v/=}T.=��-==�,=p�+=�+=�>*=rh)=ѐ(=I�'=��&=��%=r%= '$=Y0#=�."=� != =��=l�=�U=|�=P�=�=V�=�=
j=��="=�M=��=#�
=��=��=r= +=98=~�<�~�<�r�<�Y�<�4�<��<���<1��<TH�<��<���<r}�<OA�<m�<8��<���<���<r�<9V�<�:�<g�<���<*ۢ<s��<���<�Q�<��<���<��<zf�<`(�<M�y<�[q<��h<r`<�X<��O<7G<_�><�}6<�$.<G�%<&n<�
<I�<*<W�;�I�;>2�;m�;��;S��;:�;�C�;h:_;�B>;�;s��:���:P�v:r�9�Q���dC}�z���!�����_2:��eX�wBv�Lۉ�XW��⍦��v��2» Fϻ�!ܻ�����+ ����?<��{�Ў�Ox��;���#�YZ(��,���0��5�Y9���<�w�@�;D��[G�|�J��M��xP��?S��U�4�X��[���]�9$`��b��6e���g��]j���l�Гo��/r�)�t��^w���y�Y{|�2�����J���|9���r������^↼����U������e׋�� ���p���Ə��"��1���䓼�E���������}T��̡��0盼�$���[�����������衼���H��B~��X��������E������6櫼�;��t���}鯼�?��ޔ���糼�8������cԷ���(h��a���m����  �  LO=�xN=��M=�)M=�}L=��K= K=�hJ=��I=��H=eHH=ڔG=��F=16F=>�E=�D=�CD=J�C=jC=lB=�A=|5A=S�@=��?=qV?=�>=�>=^==}�<=�<=}U;=�:=1�9=�M9=�8=6�7=�P7=��6=26=2]5=��4=�4=g3=r�2=c2=Y1=ܠ0=��/=�!/=![.=��-=��,=
�+=y+=)K*=Ku)=��(=��'=��&=&=�%=�.$=�6#=�3"=�#!=� =A�=��=;S=v�=��=6=/�=2�=^=��=��=7@=�x=D�
=H�=h�=�=A%=4=y�<�|�<�s�<h]�<J;�<l�<���<'��<O[�<��<���<��<�[�<&�<��<�˿<僚<���<Hg�<?I�<�)�<��<:�<���<τ�<�N�<��<�֍<���<�U�<|�<��y<^+q<�h<�@`<��W<�oO<:G<��><�d6<.<:�%<�h<L<��<46<={�;uz�;ho�;�a�;�X�;)^�;�y�;ʲ�;`;�$?;�|;&H�:�.�:�7y:���9�?&�$���|����4���ش�KE:���X�ǋv����w����צ�,ɴ�c»
�ϻ*xܻ������I ����qM�������Bw�O5�1�#��I(�t�,�9�0���4���8�w�<��S@�j�C�''G�VJ�'`M��HP�QS�e�U�hX�%�Z��]��`�_�b�+1e�~�g��cj�}m�ѥo�WHr�5�t�փw��z���|�0�؀�����M�����������톼#���Z������֋�S���j��������s���ғ��1��Վ���痼�:������I͛����D���x��^���<١�%
��.>���v����������ZF��������E��ޟ�����-S��V�������iP��̞��근�2��y��$�������  �  |O=�uN=Y�M=�)M=�L=8�K="K=�oJ=�I=�I=
TH=١G=��F=�DF="�E=��D=uQD=�C=�C=�uB=�A=�;A=�@=��?=�W?=�>=+>=�Z==C�<=��;=�L;=�:=�9=�@9=�8=W�7=VC7=��6=��5=�S5=-�4=�	4=�b3=�2=�2=�Y1==�0=��/=A'/=Tb.=d�-=%�,=�+=�,+=QY*=�)=K�(=��'=��&=�&=(%=f7$=�=#=�8"=Z'!== =I�=�=�O=/�=_�==�=e�=�O=i�=�=t0=�i=�
=��=l�=�=�=�.=!r�<Ny�<ks�<�`�<�A�<��<���<̭�<�p�<G1�<���<g��<Az�<uD�<��<��<$��< ��<8z�<�X�<,6�<��<��<��<���<&J�<��<ʍ<#��<A�<���<�ry<"�p<8xh<	`<��W<<O<��F<O�><lE6<��-<B�%<�_<D	<c�<B<6��;��;m��;���;[��;S̢;��;�1�;B"a;T&@;�s;r�:�ѽ:�|:���95������E�z�����ӳ��8��e:���X�t�v��K��W㘻*1�� ,��X�»�л��ܻ>J��H���m ����c�Ǖ�����x��0�M�#��8(��,�D�0�g�4���8�6}<��@���C�n�F�?J�E&M��P���R��U��CX�F�Z��q]�-`��b�-e���g�)lj�_m��o��fr�u�?�w�vKz�3�|�|g���	/��3f������˅�a����-���a������׋�����d������
��Qd��󿓼����u��-̗�����i�������t*���`��씠�ȡ�S����3���o�����������H��	���9����R��G�����`j��	Ĳ�!��,l��#�����%J��s����λ�/���  �  �O=rN=6�M=�)M=�L=/�K=�&K=3vJ=S�I=�I=`H=a�G=� G=`TF=ȪE=E=�_D==�C=QC=�B=�A=�AA=U�@=z�?=�X?==�>=�>=dV==�<=��;=�B;=�:=��9=F29=�8=	�7=�47=�6=c�5=�H5=0�4=�4=�]3=��2=
2=�Y1=�0=.�/=�,/=ii.=_�-=��,=�
,=�:+=/h*=P�)=��(=��'=�'=E&=�2%=@$=AD#=v="=C*!=M	 =��=f�=|K=��==�=�x=<�=/@=��=��=6=�X=��
=~�=�=��=�=n(=/i�<t�<�q�<�b�<�G�<t"�<x��<ο�<���<�J�<}�<1��<!��<^d�<i2�<m�<#ڻ<β�<Z��<1h�<�A�<��<d�<��<��<�C�<_�<q��<'s�<*�<��<�7y<<�p<J7h<��_<_W<5O<��F<�f><�!6<�-<[�%<CS<R<��<�K<���;���;��;�	�;4�;R?�;6p�;���;�3b;�5A;uw ;A��:Ɂ�:*
:��9��6t���C�y�aZ��:������:�RY��Ww�P����9������똵�K>ûB}лOPݻ���h���� ��#��}�t����}}�|.���#�>)(��t,���0�P�4���8�eJ<�D�?�[C���F�n�I�y�L���O�ǯR��oU�LX���Z��[]�!�_��b��+e�1�g��xj��&m�?�o���r��8u���w���z�,}������'L��1���
���(������:���j�����ً�&���_��̬�������T����������[��n���L����J������Ҝ����H�����Զ����)��ni������P���oL��m���J��ha�� î��$�����Q಼8��֊��2ض�� ��3d��]���;⻼����  �  ZO=zmN=X�M=h(M=d�L=k�K=�*K=
|J=�I=�I=�kH=|�G=�G=ocF=�E=�E=nD=�C={)C=��B=g�A=[GA=�@=Q @=�X?=��>=c>=bQ==K�<=��;=8;=Ԅ:=�9=a#9=nv8=c�7=@%7=ŀ6=e�5=X=5=��4=*�3=�W3=��2=�2=NY1=�0=��/=1/=�o.=��-=&�,={,=�G+=�v*=Q�)=��(=�'=�'=!)&=�<%=8H$=QJ#=�A"=s,!=�	 =�=(�=`F=��=v=��=�k=��=!0=��=�=�=�G=�{
= �=`�=��=�=i!=�^�<wm�<�n�<Qc�<GL�<�*�<�<���<���<�c�<F*�<&��<W��<���<jP�<` �<5�<uȷ<'��< v�<L�<B�<N�<_��<�|�<�;�<|��<e��<_�<&�<rƀ<V�x<�rp<�g<
�_<�W<��N<�|F<G9><��5<��-<��%<
D<m�<0�<
S<���;U�;�7�;[�;���;��;:�;\:�;)@c;�=B;[t!;�� ;J#�:��:�5::;R7����x�� �����%����:��wY���w�ߊ����t����	��x�û��л)�ݻ:"����� �H�˚�߽�������/�1�#��(�=a,�ԃ0���4�l`8�a<�g�?� C�goF��I�Z�L���O�~~R�[EU���W�åZ�kH]� �_�҈b�U-e�~�g��j�[=m�(�o�;�r�eu��x�A�z��U}���31��"j������ʄ���������H��8u�����p܋�S���\������v���uF��k����JB�������ᘼ�+���r��G�������+1�� l��ڦ���⢼�!���d��T���L����Q��C�������q��׮�<������l����V��#�������=����'�������"0���  �  �O=�hN=��M=�&M=,�L=��K=�-K=��J=��I=5$I=�uH=S�G=�G="qF=��E=� E=�zD=��C=j3C=��B=��A=�KA=��@=V@=lX?=��>=��==L==K�<=,�;=�-;=�x:=��9=09=�g8=��7=�7=s6=��5=J25=7�4=p�3=�Q3=E�2=�2=�W1=W�0=��/=�4/=Iu.=��-=6�,=8!,=T+=��*=��)=M�(=0�'=�'=�3&=�E%=5O$=qO#=�D"=�-!=C	 =
�=f�=�@=��=*m=�=u_=��=� =]r=h�=��=�7=\l
=�=�=�=�=A=�S�<�e�<�j�<�b�<O�<�1�<��<[��<:��<�y�<�C�<i�<���<ޟ�<�k�<�9�<�	�<�۷<���<	��<%T�<�#�<��<L��<[w�<�2�< �<K��<UK�<���< ��<��x<@5p<.�g<{E_<��V<��N<�IF<><a�5<X�-<m%<?3<f�<�<�V<H��;�8�;o�;f��;ش;^�;~[�;z��;�3d;/C;�Z";��;���:j(�:;:��7���4x���������;�R�Y�NJx��)��D왻v^��!u��V%Ļ�fѻ�4޻*���k��V� ��k�����������a3���#�(��Q,��l0��e4�;8�]�;��|?�y�B��7F�FfI��xL��pO�5RR��U�d�W�ƎZ��8]���_���b��1e�2�g�˘j��Tm�Ap��r���u�hFx�l�z���}�A���N����������ㄼ�
���0��W��:���ȭ��ዼ����Z������됼9:������g۔��+��(z���Ƙ�,���V������ܝ�2���Z������آ����a��h�������)X��Ҷ�����Ӂ���ꮼ�R��O���1��t���ǵ�x���Y������EӺ�l
���@���  �  ��N=�cN=��M=�$M=f�L=f�K=�/K=��J=(�I=-+I=d~H=(�G=�&G=�|F=��E=
,E=��D=�C=�;C=��B=��A=,OA=d�@=�@=\W?=)�>=��==G==ԑ<=[�;=|$;=hn:=0�9=�9=�Z8=k�7=�	7=
g6=��5=r(5=��4=a�3= L3=��2=�2=SV1=��0=��/=J7/=vy.=ʷ-=��,= *,=7^+=ʎ*={�)=��(=7(=%'=�<&=�L%=�T$=YS#=�F"=g.!=X =��=��=�;=�=e=v�=kT=H�=h=&d=ɬ=W�=�)=_
=׎=�=��=��=�=�I�<d^�<�e�<�`�<�P�<r6�<(�<M��<���<R��<�X�<v#�<���<ѷ�<���<�N�<>�<�<��<��<Z�<�&�<y�<\��<�q�<*�<Kݑ<���<�9�<#�<���<��x<m�o<�~g<�_<2�V<o_N<DF<��=<ȴ5<T�-<W%<�"<��<@�<@X<p	�;<V�;y��;+��;� �;�h�;���;X�;e;�C;M#;�h;L��:,�:�:�G�7�H�3�w��������� 2��M;�m-Z�g�x�nm���:��Q���1Զ���Ļv�ѻ��޻�껨����3�����������ϙ��8��#��(�F,�-[0�pM4��8���;�rS?�d�B��F�27I�JKL�CGO�o-R�� U���W�}Z�x-]�T�_�W�b��7e���g�\�j��jm��/p�N�r�^�u��qx�F!{�U�}�_)���h��џ��σ�Z���m���@��Od������~���.拼6���Z��˝���吼�0���}��V˔����e�����������?������ȝ��
��cL�������Т�b���_������q���^�������&������$���g���α��1��ʍ��"⵼?.��yr��ǯ���纼P���O���  �  ��N=�_N=��M=�"M=~L=��K=S1K=+�J=�I=O0I=��H=��G=/G=^�F=��E=�4E=��D=K�C=�AC=v�B=E�A=qQA=��@=�@=:V?=��>=��==�B==��<=�;=#;=!f:=	�9=��8=�P8=G�7= 7=�]6=%�5=� 5=��4=��3=qG3=L�2=6�1=�T1=e�0=|�/=9/=e|.=�-=�,=�0,=�e+=�*=�)=o�(=}(=�,'=1C&=@R%=�X$=V#=hH"=�.!=R =��=n�=~7=��=�^=��=�K=��=�=(Y={�=�=�=�T
=I�=|�=��=_�=U=%A�<X�<�a�<_�<XQ�<�9�<#�<��<��<>��<uh�<�4�<���<���<ғ�<^�<*�<���<ĳ<s��<	^�<2(�<��<Z��<Rl�<�"�<�ӑ<���<>+�<�Մ<J��<�fx<��o<)Tg<^�^<�V<�8N<<�E<c�=<�5<�o-<�D%<<m�<u�<UX<��;k�;��;��;�V�;���;� �;�a�;I�e;�D;7�#;'�;��:3�:v:z�7�1�k�w�����7���-X�c�;�uvZ�Ay������x������s����Ļ�һ��޻1뻽���/�2��{�����8��e��c>�o�#��(�~>,��N0��;4��8���;�M4?���B�Q�E��I�N)L��'O��R�)�T��W�{pZ��%]�O�_�"�b��=e���g�|�j�(}m�=Fp��s���u�J�x��F{���}��=��}��U����ჼ	��P,��mM��o��J�������ꋼ���[��ʛ��Pᐼ�)��Ft��z����
��!U������發b.���t�����������A��녡�~ˢ�e��B_��=�����qd���Ǫ�b0��m���,
���v���౼�D������h���6B���������������*���[���  �  I�N=)]N=��M=2!M=�~L=��K=�1K=��J=M�I=m3I=��H=�G=(4G=ŊF=�E=�9E=��D=��C=cEC=e�B=a�A=�RA=��@=^@=ZU?=z�>=��==@==-�<=��;=p;=�`:=A�9=��8=!J8=ʟ7=��6=�W6=��5=�5=�4=��3=gD3=�2=p�1=�S1=�0=��/=�9/=%~.=��-=w�,=�4,=�j+=?�*=��)=��(=�(=T1'=4G&=�U%=j[$=�W#=&I"=�.!=� =�=I�=�4=6�=]Z=��=2F=s�=M=%R=I�=��=�=N
=7=�=/�=H�=�
=�;�<�S�<_�<�]�<gQ�<�;�<��<s��<��<̢�<nr�<�?�<�
�<���<���<3h�<r2�<���<Yɳ<,��<�_�<�(�<��<��<�h�<��<B͑<�x�<"�</˄<�v�<bMx<��o<�8g<�^<1lV<k N<��E<��=<��5<va-<-9%</<)�<�<�W<�;�w�;y��;�#�;Fx�;�Ϥ;!-�;=��;��e;$�D;�$;�=;~?�:*^�:�:��7���4ww��
�����r�B�;���Z��Py��Ƌ�����
(��N��Ż�Kһk߻m_��.��4C�������'�H�����B��#�w
(�k:,�CG0�14��7���;�!?�f�B�G�E���H�"L��O�/R�+�T�W�W��hZ��!]�a�_���b��Ae�R�g���j��m��Tp�!s���u�S�x��^{��~��J������ǿ��<탼����5���U�� v������{����틼�!���[������ސ��%���n��5������-K������ܙ��#��>j��h���	���j;��0���KȢ����=_�������	��8h���̪��6��/���*��2����뱼�P������h��O��摸�"͹�D���3���c���  �  $�N=4\N=�M=� M=|~L=��K=-2K=)�J=�I=�4I=�H=��G=�5G=��F=��E=�;E=<�D=(�C=�FC=e�B=
�A=3SA=$�@=W@=U?=ߥ>=��==?==��<=��;=�;=�^:=>�9=��8=�G8=��7=��6=�U6=��5=�5=~4=��3=QC3=�2=��1=S1=��0=��/=4:/=�~.=h�-=��,=56,=l+=��*=F�)=��(=X(=�2'=�H&=�V%=5\$=2X#=eI"=�.!=P =��={�=�3=��=�X=E�=PD=b�= =�O=�=z�=S=�K
=2}=C�=��=��=�	=�9�<�R�<(^�<�]�<�Q�<R<�<��<]��<���<���<�u�<C�<��<���<��<_k�<F5�<���<�ʳ<5��<{`�<�(�<-�<嬞<9g�<��<�ʑ<�u�<��<hǄ<pr�<�Dx<�o<�/g<ѿ^<hcV<*N<J�E<�=<�5<�\-<F5%<H	<�<�<2X<��;�|�;,��;�-�;f��;�ݤ;2<�;���;�f;gE;�$$;IX;�n�:D��:I�:74�7��sw����i-��b~�Ǻ;�ǹZ�4gy��Ӌ�ɯ��8��:_���Ż ]һ�%߻�o��=��J�������]�������[D�v�#�#
(�9,��D0��-4�'�7�F�;��?�mB��E���H�!L�O�{�Q�9�T��W��fZ�m ]��_�>�b��Ce�� h�.�j�N�m�Zp�'s�m�u�ѱx��f{��~��N��]���Ă�D񃼙��$9���X��wx��	����&a"���[��Ú��
ސ�{$���l����������G��t���nؙ�����f��R���I�$9�����IǢ�q��,_��
����
���i���Ϊ��8��䦭�@�����ﱼU��񲴼����S�����ѹ�����6���f���  �  I�N=)]N=��M=2!M=�~L=��K=�1K=��J=M�I=m3I=��H=�G=(4G=ŊF=�E=�9E=��D=��C=cEC=e�B=a�A=�RA=��@=^@=ZU?=z�>=��==@==-�<=��;=p;=�`:=A�9=��8=!J8=ʟ7=��6=�W6=��5=�5=�4=��3=gD3=�2=p�1=�S1=�0=��/=�9/=%~.=��-=w�,=�4,=�j+=?�*=��)=��(=�(=U1'=4G&=�U%=k[$=�W#=(I"=�.!=� =�=O�=�4=@�=jZ=�=EF=��=h=ER=o�=�=�=BN
=q=I�=q�=��=1=E<�<�T�<�_�<M^�<�Q�<�;�<-�<���<p��<��<�r�<�?�<�
�<���<l��<�g�<,2�<:��<�ȳ<���<�_�<((�<1�<���<?h�<2�<�̑<gx�<�!�<�ʄ<Rv�<Mx<��o<�8g<7�^<lV<� N<v�E<N�=<p�5<`b-<):%<7<7�<�<�X<�;�y�;��;%�;oy�;�Ф;�-�;��;s�e;[�D;S$;�;;8:�:�W�:G�:N��79���w�����%���w�)�;���Z�&Uy�ɋ�����)���O���	ŻXMһ�߻~`��/���C�T��
��d�{�����B��#��
(�}:,�RG0�!14��7� �;�!?�k�B�J�E���H�$L��O�0R�,�T�X�W��hZ��!]�a�_���b��Ae�R�g���j�	�m��Tp�!s���u�T�x��^{��~��J������ǿ��<탼����5���U�� v������{����틼�!���[������ސ��%���n��5������-K������ܙ��#��>j��h���	���j;��0���KȢ����=_�������	��8h���̪��6��/���*��2����뱼�P������h��O��摸�"͹�D���3���c���  �  ��N=�_N=��M=�"M=~L=��K=S1K=+�J=�I=O0I=��H=��G=/G=^�F=��E=�4E=��D=K�C=�AC=v�B=E�A=qQA=��@=�@=:V?=��>=��==�B==��<=�;=#;=!f:=	�9=��8=�P8=G�7= 7=�]6=%�5=� 5=��4=��3=qG3=L�2=6�1=�T1=e�0=|�/=9/=e|.=�-=�,=�0,=�e+=�*=�)=o�(=}(=�,'=2C&=AR%=�X$=V#=lH"=�.!=X =��=z�=�7=��=�^=��=�K=ʯ=	=fY=á=a�=�=�T
=��=��=�=��=�=?B�<0Y�<�b�<!`�<YR�<�:�<��<���<���<���<�h�<�4�<���<���<���<^�<�)�<���<Só<���<]�<;'�<��<Z��<Wk�<�!�<�ґ<��<�*�<3Մ<؁�<	fx<`�o<&Tg<��^<��V<�9N<`�E<��=<��5<�q-<�F%< <x�<�<SZ<��;�n�;��;��;5Y�;C��;��;ub�;�e;|�D;t�#;1�;���:�ރ:9�:`*�7v񹀲w����R���a�ێ;��Z�y�ۧ���|��a����!����ĻFһW�޻*3뻆���0�ئ������������>���#��(��>,��N0��;4�8���;�Y4?���B�X�E��I�S)L��'O��R�+�T��W�|pZ��%]�P�_�#�b��=e���g�}�j�(}m�=Fp��s���u�J�x��F{���}��=��}��U����ჼ	��P,��mM��o��J�������ꋼ���[��ʛ��Pᐼ�)��Ft��z����
��!U������發b.���t�����������A��녡�~ˢ�e��B_��=�����qd���Ǫ�b0��m���,
���v���౼�D������h���6B���������������*���[���  �  ��N=�cN=��M=�$M=f�L=f�K=�/K=��J=(�I=-+I=d~H=(�G=�&G=�|F=��E=
,E=��D=�C=�;C=��B=��A=,OA=d�@=�@=\W?=)�>=��==G==ԑ<=[�;=|$;=hn:=0�9=�9=�Z8=k�7=�	7=
g6=��5=r(5=��4=`�3= L3=��2=�2=SV1=��0=��/=J7/=vy.=ʷ-=��,= *,=7^+=ʎ*={�)=��(=8(=%'=�<&=�L%=�T$=\S#=�F"=n.!=b =��=��=�;=4�=4e=��=�T=��=�=~d=.�=��=*=�_
=u�=��=<�=��=o=9K�<�_�<yg�<eb�<R�<�7�<X�<W��<���<��<Y�<�#�<���<���<H��<N�<~�<.�<���<䉯<�X�<J%�<�<�<*p�<�(�<ܑ<���<�8�<R�<��<��x<��o<�~g<$_<�V<�`N<�F<��=<	�5<Ԉ-<�Y%<�%<��<"�<[<��;8[�;���;
��;�#�;/k�;D��;�;�e;��C;e#;Nc;��:��:,�:��7K��<�w�=�������?�Y[;�v:Z���x�\s��@��s����ض�ߌĻ<�ѻ �޻���/���*���w�������A��59�5�#��(�NF,�T[0��M4��8���;��S?�q�B��F�:7I�PKL�HGO�s-R�� U���W�}Z�z-]�U�_�X�b��7e���g�\�j��jm��/p�N�r�_�u��qx�F!{�U�}�_)���h��џ��σ�Z���m���@��Od������~���.拼6���Z��˝���吼�0���}��V˔����e�����������?������ȝ��
��cL�������Т�b���_������q���^�������&������$���g���α��1��ʍ��"⵼?.��yr��ǯ���纼O���O���  �  �O=�hN=��M=�&M=,�L=��K=�-K=��J=��I=5$I=�uH=S�G=�G="qF=��E=� E=�zD=��C=j3C=��B=��A=�KA=��@=V@=lX?=��>=��==L==K�<=,�;=�-;=�x:=��9=09=�g8=��7=�7=s6=��5=J25=7�4=p�3=�Q3=E�2=�2=�W1=W�0=��/=�4/=Iu.=��-=6�,=8!,=T+=��*=��)=M�(=0�'=�'=�3&=�E%=8O$=uO#=�D"=�-!=N	 =�=z�=A=��=Tm=C�=�_=��=5!=�r=�=z�=X8=m
=ϛ=��=��=�=1=�U�<�g�<tl�<rd�<�P�<@3�<B�<���<K��<�z�<D�<��<���<���<Mk�<�8�<��<^ڷ<Q��<���<�R�<&"�<��<���<�u�<1�<{�<뙍<#J�<���<;��<s�x<�4p<)�g<�E_<��V<,�N<�KF<�><#�5<g�-<`p%<�6<��<��<[Z<���;�>�;�t�;$��;�۴;P�;m]�;Y��;Z3d;g,C;�U";�;��:*�:%
:�7�7^��7sx��!�����A�A;�I�Y��Yx�1��󙻾d���z���*Ļ�kѻ�8޻����n���� ��l���N��W������3��#�h(��Q,�
m0��e4�;;8�v�;��|?���B��7F�PfI��xL��pO�:RR��U�g�W�ȎZ��8]���_���b��1e�3�g�˘j��Tm�Ap��r���u�hFx�l�z���}�A���N����������ㄼ�
���0��W��:���ȭ��ዼ����Z������됼9:������g۔��+��(z���Ƙ�,���V������ܝ�2���Z������آ����a��h�������)X��Ҷ�����Ӂ���ꮼ�R��O���1��t���ǵ�x���Y������EӺ�l
���@���  �  ZO=zmN=X�M=h(M=d�L=k�K=�*K=
|J=�I=�I=�kH=|�G=�G=ocF=�E=�E=nD=�C={)C=��B=g�A=[GA=�@=Q @=�X?=��>=c>=bQ==K�<=��;=8;=Ԅ:=�9=a#9=nv8=c�7=@%7=ŀ6=e�5=X=5=��4=*�3=�W3=��2=�2=MY1=
�0=��/=1/=�o.=��-=&�,=z,=�G+=�v*=Q�)=��(=�'=�'=")&=�<%=;H$=UJ#=�A"=},!=�	 =.�=?�=~F=�=Ev=��=2l=��=�0=�=��=;=�H=Q|
=ة=H�=��=�=u"=�`�<�o�<�p�<\e�<7N�<�,�<��<��<���<d�<�*�<���<m��<M��<�O�<��</�<3Ƿ<���<|t�<@J�<c�<a�<p��<�z�<�9�<��<ܩ�<�]�<	�<�ŀ<(�x<rp<�g<��_<!!W<d�N<�~F<�;><��5<h�-<`�%<�G<^ <"�<�V<���;#�;�=�;Q`�;��;_��;b�;T;�;�?c;;B;o!;� ;��:�Ԁ:8�:[
C7�����#y��D��������8�:���Y���w�犻����v�����?�û	�л��ݻ6&�A���� �ZI�ڛ�¾�J�����0���#�(��a,��0�߃4��`8�}<�}�?�+ C�uoF��I�b�L���O��~R�_EU���W�ťZ�mH]��_�Ԉb�V-e��g��j�\=m�(�o�<�r�eu��x�A�z��U}���31��"j������ʄ���������H��8u�����p܋�S���\������v���uF��k����JB�������ᘼ�+���r��G�������+1�� l��ڦ���⢼�!���d��T���L����Q��C�������q��׮�<������l����V��#�������=����'�������"0���  �  �O=rN=6�M=�)M=�L=/�K=�&K=3vJ=S�I=�I=`H=a�G=� G=`TF=ȪE=E=�_D==�C=QC=�B=�A=�AA=U�@=z�?=�X?==�>=�>=dV==�<=��;=�B;=�:=��9=F29=�8=	�7=�47=�6=c�5=�H5=0�4=�4=�]3=��2=
2=�Y1=�0=-�/=�,/=ii.=^�-=��,=�
,=�:+=/h*=P�)=��(=��'=�'=F&=�2%="@$=FD#=}="=M*!=Z	 =��=~�=�K=	�=B=�=	y=��=�@=1�=K�=�=�Y=O�
=]�=�=��=�=�)=dk�<Pv�<t�<�d�<�I�<P$�<&��<G��<�<�K�<,�<���<8��<'d�<�1�<��<ٻ<���<Ջ�<~f�<@�<��<f�<��<�<�A�<���<۹�<�q�<�(�<
�<�6y<��p<C7h<i�_<E`W<�O<B�F<�i><%6<��-<)�%<@W<g<԰<�O<5��;���;b��;C�;�#�;�B�;rr�;���;;3b;x2A;�q ;e��:em�:�~:�X�9u�6�T��sz����n���6����:��1Y�]iw������A��������FDû��лUݻ�������o� �%��~�_��ԧ�~� /�*�#��)(�u,��0�}�4�ʊ8��J<�[�?�[C���F�y�I���L���O�̯R��oU�OX���Z��[]�#�_��b��+e�2�g��xj��&m�@�o�r��8u���w���z�,}������'L��1���
���(������:���j�����ً�&���_��̬�������T����������[��n���L����J������Ҝ����H�����Զ����)��ni������P���oL��m���J��ha�� î��$�����Q಼8��֊��2ض�� ��3d��]���;⻼����  �  |O=�uN=Y�M=�)M=�L=8�K="K=�oJ=�I=�I=
TH=١G=��F=�DF="�E=��D=uQD=�C=�C=�uB=�A=�;A=�@=��?=�W?=�>=+>=�Z==C�<=��;=�L;=�:=�9=�@9=�8=W�7=VC7=��6=��5=�S5=-�4=�	4=�b3=�2=�2=�Y1==�0=��/=A'/=Tb.=d�-=%�,=�+=�,+=QY*=�)=K�(=��'=��&=�&=
(%=j7$=�=#=�8"=c'!=K =[�=��=�O=U�=��=T=f�=��=@P=�=��=1=Cj=ܛ
=f�=T�=�==�/=Bt�<q{�<�u�<�b�<�C�<��<5��<7��<�q�<62�<���<ȴ�<Wz�<AD�<
�<��<��<ݚ�<�x�<>W�<f4�<��<��<��<ځ�<UH�<0
�<�ȍ<΄�< @�<���<�qy<��p<2xh<�`<��W<�=O<��F<��><~H6<)�-<�%<�c<5<T�<�E<���;N��;���;��;���;�Ϣ;��;�2�;�!a;d#@;�n;�:㽽:0�{:�b�9�gJ��j�� %{��һ��������ew:���X���v��S���꘻*8��e2���»�л��ܻ;N�=L��o �&��d����@��yy�'1���#��8(�P�,�{�0���4�ڶ8�Q}<��@���C�{�F�JJ�M&M��P���R��U��CX�H�Z��q]�.`��b�-e���g�)lj�_m��o��fr�u�?�w�vKz�3�|�|g���	/��3f������˅�a����-���a������׋�����d������
��Qd��󿓼����u��-̗�����i�������t*���`��씠�ȡ�S����3���o�����������H��	���9����R��G�����`j��	Ĳ�!��,l��#�����%J��s����λ�/���  �  LO=�xN=��M=�)M=�}L=��K= K=�hJ=��I=��H=eHH=ڔG=��F=16F=>�E=�D=�CD=J�C=jC=lB=�A=|5A=S�@=��?=qV?=�>=�>=^==}�<=�<=}U;=�:=1�9=�M9=�8=6�7=�P7=��6=26=2]5=��4=�4=g3=r�2=c2= Y1=ܠ0=��/=�!/= [.=��-=��,=	�+=y+=(K*=Ku)=��(=��'=��&=&=�%=�.$=�6#=�3"=$!=� =Q�=��=VS=��=Î=k=o�=��=v^=�=D�=�@=fy=��
=	�=8�=�=*&=
5=�z�<�~�<tu�<<_�<=�<	�<��<n��<`\�<|�<>��<u��<\�<�%�<���<K˿<��<؄�<�e�<�G�<W(�<�<�ߢ<�<��<"M�<��<TՍ<p��<�T�<��<w�y<�*q<�h<A`<��W<#qO<2G<�><Ug6<�.<��%<l<�<�<�9<ҁ�;���;�t�;of�;�\�;a�;�{�;���;`;�!?;�w;g:�:�:y:��9��3�2���]S|�m5��I��p���U:���X��v����B���ަ��δ�0h»��ϻ@|ܻ������dJ ����dN����Z���w��5���#��I(���,�j�0��4���8���<��S@�y�C�4'G�VJ�/`M��HP�VS�i�U�!hX�'�Z��]��`�`�b�,1e�~�g��cj�}m�ѥo�WHr�5�t�փw��z���|�0�؀�����M�����������톼#���Z������֋�S���j��������s���ғ��1��Վ���痼�:������I͛����D���x��^���<١�%
��.>���v����������ZF��������E��ޟ�����-S��V�������iP��̞��근�2��y��$�������  �  � O=�zN=)�M=�(M=�{L=H�K=0K=�bJ=�I=��H=>H=d�G=��F=H)F=$E=E�D=n7D=�C=`�B=ScB=��A=�/A=ѓ@=��?=�T?=��>=�	>=q`==m�<=O	<=�\;=A�:=7:=�X9=��8=�8=5\7= �6=�6=&e5=Z�4=�4=!j3=�2=v2=�W1=C�0=��/=u/=}T.=��-=<�,=o�+=�+=�>*=rh)=ѐ(=J�'=��&=��%=t%='$=]0#=�."=� !=� =��=}�=�U=��=s�=�=��="=Uj=��=�=N=�=��
=��=+�='=�+=�8=��<u��<:t�<[�<6�<��<��<<��<3I�<��<��<�}�<_A�<G�<���<��<鏻<1q�<&U�<�9�<�<���<�٢<	��<#��<mP�<��<tߍ<��<�e�<�'�<q�y<\[q<��h<�r`<�X<ޛO<�8G<R�>< �6<O'.<��%<�p<�<+�<�,<v\�;�N�;�6�;M�;��;���;��;8D�;:_;�@>;�;:��:��:��v:"�9�ᔷMG�qv}������<��&���?:��rX��Nv�9ቻ�\�����_{��m»�Iϻ�$ܻ���v���), ����=��|�Z���x��;��#��Z(���,���0�5�s9���<���@�GD��[G���J��M��xP��?S��U�6�X��[���]�:$`���b��6e���g��]j���l�Гo��/r�*�t��^w���y�Y{|�2�����J���|9���r������^↼����U������e׋�� ���p���Ə��"��1���䓼�E���������}T��̡��0盼�$���[�����������衼���H��B~��X��������E������6櫼�;��t���}鯼�?��ޔ���糼�8������cԷ���(h��a���m����  �  Z#O=O|N=K�M=�'M=�yL=?�K=%K=�]J=ѥI=u�H=�5H=]�G=��F=HF=uE=U�D=�-D=<�C=w�B=^\B=��A=�*A=��@=��?=�R?=ɯ>=
>= b==0�<=h<=b;=ʶ:=�:=9a9=;�8=�8=�d7=�6=�6=k5=�4=�4=4l3=��2=72=uV1=��0=��/=/=O.=�-=̱,=�+=�
+=5*=w^)=؆(=��'=��&==�%=%%=� $=6+#=�*"=�!=� =��=˟=OW=]�=��=V#=J�==Cs=��=~=�W=��=��
=]�=�=�=�/=�;=���<��<�r�</W�<�/�<���<[��<6��<:�<h��<#��<�i�<�,�<���<���<��<�~�<�a�<�G�<O.�<��<a��<�Ԣ<B��<���<R�<�<��<4��<cr�<�6�<T�y<�q<b
i<��`<�'X< �O<�TG<V�><ё6<�3.<y�%<us<�<^�<�!<�<�;�%�;I�;J��;W��;��;5��;��;Չ^;n�=; �;Yi�:1��:>}t:+��9&0ķ�}��h~�$�Mp��x���2:�QX�0v�溉��,��:Z��m<������Wϻn�ۻJ`軬x��� �@���0�Lu�����z�B�$�#��h(���,�11�{+5��&9��<���@��+D�D�G�9�J���M�'�P�bS��V���X��-[��]�/2`�P�b��<e���g��Zj�+�l��o��r�>�t�YCw���y�uY|��~�>����큼.*��^e��ȟ���ن���/R��뒊��؋�$��v��9Ώ�,��������UU��~������Kh�����D���T8��n������Mʠ�1���M!��oP���������������E��Z����᫼=4������5ݯ�n1�������ֳ�Q'��gv��ķ�e���[��@������  �  �$O=�|N=2�M='M=+xL=@�K=zK=`ZJ=ѡI=��H=�0H=�zG=��F=�F=�nE=��D=�'D=��C=_�B=�WB=�A=�'A=y�@=��?=�Q?=,�>=
>=�b==ֹ<=�<=Re;=ú:=n:=if9=��8=@8=	j7=��6=�6=�n5=��4=�4=am3=O�2=�2=zU1=[�0=L�/=A/=�K.=�}-=�,=��+=�+=�.*=X)=t�(=w�'=�&=��%=p%=�$=�'#=("=�!=U =B�=ܟ=X=� = �=�&=p�=�=�x=��=�=^=��=��
=�=�=� =2="==��<��<q�<aT�<�+�<��<I��<�w�<40�<T��<$��<�\�<��<d��<��<��<�s�<�W�<?�<'�<��<��<uѢ<K��<!��<bS�<� �<:�<d��<4z�<+@�<�z<k�q<�!i<��`<�=X<��O<yeG<4�><C�6<�:.<�%<t<=	<B�<�<L'�;~
�;��;���;��;<��;Ŋ�;yl;
^;Y"=;Ë;̠�:}ո:P6s:�h�9�B�qD���\)��8������u,:�}<X���u�%�������6����������λY�ۻ:軪W�� ����K)�0q����c|�rF��#�r(���,��1��<5�l:9��=���@��DD�`�G�L�J���M�۵P�xS�% V�ʴX�I<[�ռ]�e;`��b��@e��g��Yj���l�so��r�*�t��2w�1�y�XD|��~�R���"ぼ� ��F]������Ԇ����qP�������ً�z&���y��ӏ�*2��B���{���b_���������u��Ú�9���D���y�������Ӡ�T���(���U����������� ���E��_����ޫ��/�������կ��(���z���˳�D���k��칷�e���S�����_켼�  �  �O=rnN=��M=M=EhL=N�K=-K={OJ=��I=��H=S.H=�zG=�F=wF=ioE=��D=)#D=��C=�B=DB=\�A=LA=i@=	�?=�$?=u>=��==l.==��<=��;=+;=6~:=L�9=l$9=�w8=�7=Y7=�q6=��5=25=�h4=8�3=�3=�S2=��1=��0=&#0=	`/=q�.=��-=K�,=�*,=�T+=�|*=��)=9�(=F�'=�'=�$&=<%=�M$=X#=�Y"=Q!=�< =G=<�=s�=�h=�=>�=P8=��=2,=�=t�=&B=��=��=*�	=|*=rP=ao=ه=� =�K�<YW�<�V�<�J�<�3�<P�<{��<c��<���<�R�<e�<��<���<Z��<Ji�<,H�<F+�<��< ��<��<gʪ<��<0��<�p�<wK�<o"�<U��<�Ǎ<疉<�d�<2�<��y<��q<�2i<��`<zmX<�P<{�G< [?<�7<��.<�Z&<<��<�F<��<0��;�;%�;�1�;�Q�;Ӂ�;1ɓ;.�;�ne;��D;�w$;�r;'r�:���:Q:���8����UZ�.F���Ͳ�w�/�4IM��j�G���)���|螭����*Ȼq�Ի 6��=�p�����������c����D��nu �K%�>l)�w�-���1�4�5�j�9��{=��A�k}D���G���J�#�M�/�P���S�#dV�yY�˹[��Z^�i�`�U�c�`;f�v�h��k�o%n���p��gs��v���x��2{�N�}�%)���n��w���\���{7���y������p���H������%㌼�6��o����됼K��y�������i��ė�i��7h�����D��/��,h��j����ѡ�����=��5x��L�������=C������/߫�.1�������د��,��F���5ӳ�/%��wv���Ʒ�T��Xe��%�������  �  SO=BnN=��M=9M=�hL=ƷK=�K=XPJ=��I=��H=�/H=�{G=��F=	F=�pE=�D=�$D=�C=`�B= EB=`�A=!	A=�i@=y�?=%?=�>=��==,.==�<=��;=,*;=)}:=�9=$#9=\v8=��7=7=hp6=��5=55=h4=��3=_3=�S2=��1=*�0=�#0=�`/=0�.=��-=W�,=�+,=7V+=j~*=��)=��(=��'=#
'=&&=g=%=�N$=Y#=�Z"=�Q!=j= =�=\�=Q�=Hh=G=�=\7=U�=�*=��=��=�@=�=5�=��	=#)=3O=an=�=[� =�J�<�V�<�V�<@K�<�4�<��<)��<G��<F��<,U�<B �<0��<���<���<�l�<?K�<8.�<^�<i��<��<+̪<O��<3��<kq�<�K�<Z"�<���<uƍ<J��<�b�<�/�<��y<=�q<�,i</�`<�gX<�	P<��G<�V?<�7<s�.<�X&<<}�<IG<�<���;0�;� �;�:�;_\�;���;֓;�;�;ވe;��D;0�$;�;��:)��:i:���8x���A'Z�q3�����Ư�T�/�)MM�a�j�ă�����q���Χ�����Ȼ��Ի�>ỤE������ʓ����������2���s �%�$�i)���-���1�^�5�޻9��u=��	A�NwD���G���J�D�M���P�#�S��_V��Y���[��X^���`�^�c�c;f���h�=�k��'n���p��ks��v�y�x�8{���}��+��q��ش��w���a9��2{���������I�������⌼#6��A���1ꐼ�H��O���1	��g�����7��:e��孛�1�	-��{e������ϡ����R<��Dw����������YC������ૼm2��=����گ��.��Ȃ���ճ��'��y��Rɷ����eg��굻�����  �  O=�mN=��M=�M=�iL=-�K=�K=�RJ=��I=2�H=�3H=#�G=�F=� F=�uE=��D=)D=�C=!�B=\HB=!�A=aA=zk@=��?=�%?=�>=��==W-==��<=��;=�';=z:=��9=?9=>r8=��7=7=�l6=C�5=i5=�e4=��3=A3=S2=��1=��0=�$0=b/=;�.=4�-=X-=,/,=0Z+=��*=�)=e�(=i�'=�'=E*&=RA%=YR$=\#=�\"=�S!=�> =d=��=�=xg=�=n�=�4=�='=G�=O�=�;=J�=��=h�	=V%=�K=�k=߄=ϗ =I�<V�<NW�<�L�<Z7�<0�<���<��<H��<*]�<�(�<���<E��<S��<�u�<-T�<�6�<��<��<]�<�Ъ<䴦<Õ�<�r�<�K�<�!�<��< Í<���<]�<�(�<��y<7�q<i<��`<#WX<i�O<J�G<�K?<��6<��.<�T&< <��<�I<��<���;+�;�7�;�U�;A|�;ڰ�;8��;Qd�;;�e;9E;8�$;��;�.�:�+�:�B:Î�8�X��+�Y�������֪�3�/�W\M�(�j��ԃ�E�����Zĭ��*��>Ȼ��Ի�Z�>^�d���$����������^��l��o �j�$��`)�?�-�+�1��5���9�xd=��@�1dD���G���J���M�f�P�S��SV�PY�A�[�"R^�[�`�Жc�;f���h�h�k�.n�f�p�pvs��v�=�x�H{�Y�}�4���x����������>��2����������I��G���ጼ�3�������吼�C��󢓼����^��]�������[��h���&眼�$���]��S����ɡ�����b8��Xt�����������C��8����⫼�5���i௼�5��c����ݳ�J0��8����з����Hm������r���  �  �O=MlN=-�M=M=�jL=E�K=�	K=bVJ=�I=}�H=q9H=��G=�F=(F=}E=�D=0D=��C=��B=�MB=u�A=�A=6n@=��?='?=�>=��==�+==N<=��;=w#;=u:=��9=9=�k8=��7=�7=�f6=�5=�5=#b4=8�3=f3=R2=��1=u�0=&0=zd/=]�.=#�-=-=�4,=K`+=^�*=!�)=��(=��'=�'=�0&=[G%=�W$=�`#=�`"=�V!=�@ =�=��=��=�e=b=�=V0=Ů=� =��=�=54=�{=b�=��	=-=�F=Jg=w�=R� =�E�<�T�<�W�<�N�<e;�<��<s��<���<.��<�i�<�6�<�<[��<i��<���<7b�<nC�<k'�<�<��<�ת<4��<]��<�t�<.L�<��<��<a��<<YS�<n�<��y<<fq<6�h<��`<�<X<��O<t�G<9?<��6<��.<SM&<��<ۧ<sM<�<k�;7�;"\�;&��;���;��;[8�;W��;�\f; �E;�^%;)N;i�:�:_�:l��8������X�%Ʃ�k�溝��'�/�3vM�a�j���7��r9����[��DoȻ�)ջ��Ỳ��%���2����K���������5h �6�$�SS)��-�x�1���5���9�I=�Z�@�rFD�ÎG�:�J�r�M�X�P�[}S��?V��X�5�[�H^���`�w�c��:f��h�e�k��8n���p�E�s��*v���x�'a{�~�}�A��W����ǂ����G������Ň�����J��˒��ߌ�0��n����ސ�!;��̘��\���R������j����L�������؜�>���Q����������h���h2���o��򱦼�����C�������櫼�;�������鯼�@��j����과c=�����ݷ��*���v���»�����  �  �O=qjN=p�M=nM=7lL=��K=/K=[J=��I=.�H=AH=.�G=0�F=�1F=��E=w�D=9D=ȕC=O�B=�SB=ٳA=GA=wq@=��?=7(?=4�>=��==�)==|<=.�;=�;=dn:=H�9=�9=c8=E�7=4
7=�^6=ɳ5=�5=!]4=`�3=�3=�P2=G�1=$�0=�'0=5g/=6�.=�-=-=�;,=h+=��*=E�)=�(= (=�'=�9&=O%=~^$=ef#=\e"=Z!=>C =�=)�=��=�c=	=n�=r*=��=�={~=\�=D*=�q=��=��	==�?=_a=�|=� =vA�<�R�<�W�<hQ�<@�<%�<��<H��< ��<�y�<RH�<��<���<��<���<-t�<�S�< 6�<��<���<,�<q��<}��<�v�<�K�<��<��<W��<j~�<yF�<_�<�y<Bq<Q�h<w`<pX<G�O<�nG<� ?<��6<��.<C&<4�<��<YQ<}�<�'�;^[�;��;R��;>�;0�;*��;��;fg;�^F;��%;V�;��:/�:�<:W��8�F���X�;|�����E����/�l�M��k�e��g��4q���/��'����Ȼjջ���{��FS��@E�ױ������)����C` �g�$�C)�v�-��1��5��r9��%=��@� D�DhG�ߏJ��M�K�P��`S�\'V���X��[��<^�&�`�&�c��;f�f�h�>�k�iGn�U�p��s��Fv��x��{�4~�qR������ւ�����R��J���ḋ�[��0M��Ғ���܌��+��.��m֐��0��&����甼�A�������똼�9��ł���Ɯ�,��FB���{������#+���j��ݮ������5E�����G쫼!D��0�������PO�����������N��V���f�w9��߃��nͻ����  �  	O=�gN=<�M={M=�mL=?�K=�K= `J=��I=��H=�IH=ɘG=�F=T<F=��E=0�D=0CD=5�C=��B=0[B=ԹA= A=�t@=,�?=@)?=�>=��==�&==�w<=��;=
;=df:=D�9=9=�X8=��7=* 7=rU6=J�5=a5=W4=��3=\�2=�N2=q�1=��0=�)0=j/=Z�.=l�-=�-=tC,=q+=��*=��)=��(=�
(=$)'=+C&=�W%=:f$=�l#=tj"=�]!=�E =!=�=�= a=�=��=]#=A�= =�s=��=�=f=Y�= �	=t=%7=MZ=w=�� =�;�<�O�<W�<�S�<�D�<�,�<K�<r��<��<���<^\�<[-�< �<,��<O��<���<�f�<�F�<�'�<.	�<=�<�Ʀ<���<x�<iJ�<��<��<p��<�q�<�6�<^��</�y<�q<��h<�K`<��W<��O<LG<�?<m�6<�y.<6&<��<ͤ<�T<'�<�C�;؂�;R��;���;E6�;���;�ޔ;�R�;�g;�G;�&;��;"R�:���::��9m޶�Q7W��2��Aw�ī��/�[�M��dk�JH����������x��4黻��Ȼc�ջ����-����[�w�������G����YX ���$��1)�l-�Ԅ1��z5�N9��<���@�=�C�s<G�OeJ�5qM��cP�S@S�V�S�X��[�[0^���`���c�n>f���h�S�k��Yn��q��s�fhv�/y���{�W@~��f��ʩ��邼�%��`������Շ�L��iP������#ی��'���x��=͐��$���}��ה�/��t���W֘��#��!m��걜��򝼨0���l��O����䢼d#���e��򫦼I���ZG��������6N��﩮�����`������"��ec������� ��K��j���yڻ�|!���  �  �O=�dN=��M=M=qnL=��K=�K=eJ=h�I=bI=�RH=עG=g�F=�GF=�E=��D=�MD=�C=nC=�bB=�A=�A=@x@= �?=�)?=N>=w�==�#==s<=x�;=c;=]:=Q�9=H�8=�M8=��7=1�6=K6=�5=&�4=*P4=-�3=R�2=�K2=-�1=��0=�*0=�l/=a�.=��-=p-=wK,=Cz+=��*=��)=�(=(=4'=`M&=a%=n$=[s#=�o"=~a!=�G =�!=j�=�=�]=��=M�=e=ٕ=x=h=��=�=@Y=��=Z�	=�=�-=bR=�p=�� =�4�<|K�<0V�</U�<pI�<34�<��<��<e��<���<�q�<	D�<y�<���<%��<�<�y�<�W�<]6�<��<)�<%ͦ<֤�<�x�<"H�<z�<;ۑ<��<c�<~%�<��<gZy<��p<r~h<
`<�W<<pO<�%G<��><1�6<wd.<R&&<��<ޠ<QV<�<I_�;���;���;s6�;|��;.ץ;M<�;V��;��h;��G;�v';[C;	��:��:�:� 
9y{��+aV��󨺪c�U���0��N�Q�k��~���ᒻy���Eɮ��=��Uɻ�	ֻ�Y�fD����u������/�������Q ���$�s )�TU-��h1��Y5�@(9��<��]@��C�7G�^8J�GM��=P�BS���U���X��n[��$^���`���c��Bf���h���k��nn��'q�j�s�t�v�+6y���{��m~�i}��Z���9����7��p��P����އ�e���T��0���"ڌ��#��.r��1Đ����eo��Ɣ���� o��Ϳ�����HV������yޝ����]��(���Rڢ�����`��٩������zJ������f����Y��R�������s���β�D&��z���ɶ�����^������+黼H-���  �  �O=FaN=R�M=GM=�nL=P�K=�K=�iJ=c�I=�
I=Y[H=��G=�F=�RF=e�E=��D=dXD=��C=�C=�iB=��A=� A=#{@=��?=
*?=/~>=��==�==�m<=Ѻ;=;=[T:=�9=D�8=8B8=%�7=��6={@6=B�5=��4=�H4=K�3=��2=�H2=p�1=1�0=�+0=o/=��.=��-=�-=BS,=@�+=��*=O�)=1�(=-!(=�>'=LW&=�i%=�u$=�y#=Gt"=�d!=�I =!"=Q�=��=�Y=u�=l�===�=��=%\=ݴ=�=;L=Q�=r�	=�=9$=J=�i==� =�,�<~F�<�S�<�U�<M�<�:�<� �<���<E��</��<,��<.Z�<�.�<��<b��<Ĳ�<Ō�<h�<�C�<��<%��<PҦ<#��<6x�<�D�<@�<ґ<ד�<�S�<��<Ԁ<p-y<[�p<�Mh<��_<C�W<�DO<��F<¿><B�6<[M.<�&<@�<'�<3V<�<\w�;��;�!�;gt�;�ʶ;�*�;���;�;�Si;��H;3(;5�;5��:�&�:��!:��9cU��ͪU��Ĩ�`����30��ON�l�춄��$���I��7��������ɻ�_ֻ������	��M�������^"����>��oM ���$�)�v@-�N1��95�a9�+�<�2@���C���F��J�	M��P��R�5�U�ϞX��_[��^�m�`�Սc�If��i���k�n�9Dq���s���v�L`y�b|���~�T����Ձ����VJ��"���괆��釼b ��"Z������ڌ�B!���l���������ya��w������`Z��ϩ��E����?�������ʝ�����M��܎���Т�,���\������$����N��|������f��MǮ�D(������B䲼�<������඼�+���r��a���h����9���  �  ��N=�]N=ݺM=M=�nL=��K=NK=�mJ=��I=hI=-cH={�G=�G=]F=��E=�	E=�aD=>�C=pC=pB=��A=�$A=i}@=��?=�)?=�|>==�==�==�h<=\�;=��:=}K:=`�9=��8=b78==�7=I�6=k66=��5=j�4=�A4=��3=S�2=E2=Z�1=Y�0=),0=�p/=��.=-�-=y%-=:Z,=X�+=�*=�)=I	)=C+(=tH'=K`&=�q%=�|$=�~#=Zx"=]g!=�J ="=��=ͧ=�U=�=��==݂=�=�P=�=Z�=�?=a�=3�	=��=�=B="c=�} =�$�<�@�<Q�<�U�<�O�<z@�<)�<T�<���<���<��<sn�<�C�<��<���<�ſ<���<�v�<P�<)�<� �<?֦<{��<�v�<�@�<��<�ȑ<χ�<1E�<+�<{��<�y<=�p<�h<��_<gW<IO<��F<��><Ni6<�6.<�&<��<�<�T<�<֊�;���;&M�;���;Z�;�v�;]�;�n�;�j;�\I;��(;�;���:�:-V#:��9����U�����'m溘���b0���N�#ol��f��D����j��缻��ɻq�ֻ��
��I����q��-�".�������J �]�$�")�0.-��61��5�(�8��<�
@�IoC�d�F���I���L�5�O�'�R���U���X��R[��^���`���c��Pf�5i�t�k�G�n��_q�5t�:�v�)�y��-|��~�
���ꁼz%��G\��揅��t􇼖(���_������ڌ���th������P��1U�����������G�������ᙼ�+��s��ĸ������b@������Ȣ�����Y��Z���Z���3S���������+r���ծ�V9����������mR��禵�.���$@�������Ǻ�N��XF���  �  �N=,ZN=v�M=�M=�nL=c�K=:K=�pJ=��I=�I=�iH=�G=�G=�eF=f�E=6E=�iD=}�C=�C=5uB=��A=a'A=@=-�?=@)?={>=��====�c<=��;=��:=�C:=ˏ9=��8=�-8=��7=��6=�-6=چ5=(�4=�;4=F�3=�2=lB2=B�1=T�0=6,0=�q/=9�.=��-=!*-=�_,=�+=��*=]�)=�)=�3(=�P'=�g&=�x%=$�$=w�#=�{"=Pi!=�K =�!=X�=!�=�Q=$�=��=�=�z=��=�F=g�=��=45=�u=O�	=��=�=;= ]=�x =/�<�;�<N�<U�<{Q�<�D�< 0�<��<Q��<���<Ȩ�<��<CU�<�*�<���<�տ<⫻<΂�<�Y�<�0�<��<�ئ<���<u�<�<�<y �<��<�|�<�7�<��<O��<L�x<�dp<�g<i�_<B@W<�N<�F<]�><iP6<�!.<t�%<R�<�<BR<�<s��;;�;�p�;q��;�D�;���;"2�;���;�j;�I;�o);E	;���:�:��$:��9_,��-�T�q���y��S��0�z�N���l�� ��\����ҡ������/��dIʻ(�ֻe<�Fﻃ������9��=�c9�G�����I ���$�N�(��-�O#1�b5�a�8��f<�1�?�NLC�p�F���I�w�L�C�O�w�R�R�U��}X��H[�[^�'�`��c��Xf��i���k���n�/xq��;t�R�v�z�y�S|�`�~���������6���k��Ν���͆�@���<0��:e�����8܌����_e���������K��K���`镼�7������IЙ�3���b�������K5��({��O¢����X�����������W��'���d��}���⮼6H��F����
��?e�����	��IR��q����ֺ����uQ���  �  v�N=OWN=j�M=nM=0nL=��K=�K=�rJ=�I=�I=�nH=��G=�G=lF=��E=�E=�oD=��C=e C=yB=��A=^)A=5�@=X�?=�(?=�y>=d�====�_<=�;=��:=�=:=�9=��8=�&8=9y7=��6=�&6=��5=y�4=�64=�3=��2=�?2=z�1=Z�0=�+0=�r/=ʴ.=�-=�--=5d,=8�+=]�*=~�)=?)=1:(=�V'=�m&=�}%=R�$=#=�}"=�j!=L =!=��=�=�N=4�=�{==�=Gt=��=+?=]�=E�=�,=�m=��	=��=q=t5=dX=u =�<K7�<{K�<T�<�R�<�G�<�4�<��<.��<���<���<|��<�b�<�7�<��<w�<���<���<a�<�5�<[	�<�ڦ<Ө�<As�<U9�<&��<��<&t�<n-�<��<ס�<%�x<JFp<��g<qv_<9"W<��N<l�F<Rj><�<6<h.<]�%<��<Ԇ<�O<<���;�;8��;���;�n�;��;�f�;j�;�k;�fJ;�);�z	;���:�z�:ӑ%:Ѓ9U6���xT������)��0�1
O��m�7H���̓�c���毻�g��e�ʻ�0׻�q�#D������('�IJ�C�������I ���$�n�(�O-�1���4�c�8�yO<��?�2C�"zF�\�I��L�)�O���R��U��sX�!B[��
^���`�z�c�@_f�)i���k�"�n��q�?Rt�gw���y��o|� ��ˀ�+��SD��/x������l׆���x6���i�������݌�}��Oc��ૐ������C������ޕ��+���w��/Ù�=��LV��V����垼-���t��ý�����"W��b���! ���[���������΅��M��S��G�������s���ȵ����U`�������⺼��aZ���  �  $�N=mUN=
�M=�M=�mL=��K=CK=tJ=��I=MI=�qH=�G=�G=3pF=%�E=�E=�sD=V�C=E#C=[{B=D�A=�*A=ˀ@=h�?='(?=�x>=��==
==�]<=�;=�:=�9:=ل9=�8=�!8=t7=�6=@"6=d|5=��4=r34=h�3=��2=>2=D�1=��0=�+0=�r/=��.=��-=�/-=�f,=T�+=��*=`�)=T)=G>(=�Z'=q&=��%=��$=��#=;"=tk!=DL =� =�=h�=�L=��=�x=��=/p=U�=P:=.�=��=�'=�h=գ	=�=p=�1=qU=�r =�<p4�<�I�<�S�<S�<xI�<�7�<��<��<��<'��<���<)k�<U@�<��<��<<(��<Xe�<�8�<N�<aۦ<���<�q�<�6�<���<���<}n�<�&�< ߄<1��<��x<|2p<��g<jb_<2W<��N<�F<�[><06<$.<��%<{�<��<�M<�<|��;s$�;��;��;W��;��;���;(�;t_k;ʮJ;D *;��	;���:�Ԓ:? &:�49�����XT�q���խ�s1���0�\,O��.m��a��Lꓻ�%��l	��y�����ʻ�T׻Z���c�w���,��[1��R��I��^��J �߭$�[�(��-��1� �4���8��@<�2�?�O!C�^iF�e�I�E�L�F�O�߭R���U�:mX�>[�a	^���`� �c��cf��/i�^�k���n�j�q��`t��!w�<�y�B�|���QՀ�S���L��(�������p݆����:��m�������ތ�w��Fb��������?��p����ו�7$���o��к�����N��K����ߞ�(���p��ﺢ�8���V���������V^��`���$��a�����l[�������!��3}��kҵ�!��Ci������3꺼�%��`���  �  J�N=�TN=��M=7M=�mL=�K=wK=�tJ=��I=3I=�rH=*�G=G=�qF=~�E=�E=�tD=q�C=G$C=3|B=��A=�*A=�@=u�?=�'?=Mx>=l�==R==�\<=�;=��:=k8:=j�9={�8== 8= s7=v�6=� 6= {5=��4=^24=i�3=��2=|=2=ې1=V�0=�+0=�r/= �.=�-=C0-=�g,=_�+=�*=��)=�)=�?(=�['=Dr&=Á%=ˉ$=b�#=�"=�k!=FL =� =��=�=�K=��=�w=x�=�n=��=�8=o�=Z�=�%=g=C�	=��=(=�0=mT=�q =��<�3�<8I�<�S�<OS�<1J�<%9�<�!�<��<W��<���<>��<�m�<C�<P�<?�<��<��<�f�<�9�<��<�ۦ<P��<q�<�5�<-��<���<Ml�<`$�<a܄<2��<E�x<�+p<��g<�[_<�W<��N<h�F<5W><�+6<�.<9�%<��<��<�M<<���;�(�;��;��;���;:�;���;�!�;Hwk;��J;h6*;��	;7�:��:�N&:��9đ��0QT����A��t8���0�q:O�B?m��j�����-1�����Ҙ���ʻ�a׻���n�Q���f��?5��U��K���^��J �u�$��(��-��	1��4�V�8��;<���?��C��cF�0�I�f�L���O���R���U��jX��<[�	^���`��c�bef��1i� l�h�n���q��et�/'w��y���|��#�^؀�v���O����������߆����<��n��Q���ߌ�h��b��ר��V�t=��q����Օ��!��Pm��!���e���K�������ݞ�.&��~o����������V��!���n��<_�������%��m������^��kñ��$��_���bյ�F$��Pl��ή���캼�'��(b���  �  $�N=mUN=
�M=�M=�mL=��K=CK=tJ=��I=MI=�qH=�G=�G=3pF=%�E=�E=�sD=V�C=E#C=[{B=D�A=�*A=ˀ@=h�?='(?=�x>=��==
==�]<=�;=�:=�9:=ل9=�8=�!8=t7=�6=@"6=d|5=��4=r34=h�3=��2=>2=D�1=��0=�+0=�r/=��.=��-=�/-=�f,=T�+=��*=`�)=T)=H>(=�Z'=q&=��%=�$=��#=="=vk!=GL =� =�=n�=�L=��=�x=��=?p=h�=f:=G�=�=�'=�h=��	=4�=�=&2=�U=�r =��<�4�<#J�<�S�<|S�<�I�<I8�<= �<��<N��<I��<���<.k�<J@�<��<��<���<琷<e�<�8�<�
�<ۦ<!��<eq�<u6�<2��</��<.n�<z&�<�ބ<��<i�x<\2p<��g<�b_<lW<�N<]�F<u\><�06<�.<��%<A�<|�<�N<J<���;�%�;R��;��;5��;��;���;Y�;Y_k;1�J;0*;/�	;���:В::&:�9A˭��fT�Ğ��P��55���0��/O�72m�ic���듻6'���
������
�ʻ�U׻1�㻤d����q���1��R��I�3�z��J ��$�j�(��-��1��4���8��@<�6�?�R!C�`iF�g�I�F�L�G�O��R���U�;mX�>[�b	^���`� �c��cf��/i�^�k���n�j�q��`t��!w�<�y�B�|���QՀ�S���L��(�������p݆����:��m�������ތ�w��Fb��������?��p����ו�7$���o��к�����N��K����ߞ�(���p��ﺢ�8���V���������V^��`���$��a�����l[�������!��3}��kҵ�!��Ci������3꺼�%��`���  �  v�N=OWN=j�M=nM=0nL=��K=�K=�rJ=�I=�I=�nH=��G=�G=lF=��E=�E=�oD=��C=e C=yB=��A=^)A=5�@=X�?=�(?=�y>=d�====�_<=�;=��:=�=:=�9=��8=�&8=9y7=��6=�&6=��5=y�4=�64=�3=��2=�?2=z�1=Z�0=�+0=�r/=ʴ.=�-=�--=5d,=8�+=\�*=~�)=?)=1:(=�V'=�m&=�}%=S�$=Ć#=�}"=�j!=$L =!!=�=�=�N=D�=�{=V�=et=�=U?=��=~�=+-=/n=��	=��=�=�5=�X=�u =��<!8�<NL�<�T�<WS�<SH�<�5�<G�<���<���<��<���<�b�<�7�<q�<+�<��<B��<�`�<!5�<��<�٦<��<�r�<�8�<r��<i��<�s�<�,�<��<���<��x<Fp<��g<�v_<�"W<\�N<F�F<[k><�=6<�.<��%<4�<Z�<.Q<�<w��;��;���;���;^p�;�;�g�;��;Vk;�eJ;��);�w	;H��:�q�:�|%:�$9�i���T�*���x��l&�M�0�4O�B
m�mK���ϓ�.��鯻)j��z�ʻY2׻6s㻍E�V�������'��J�nC������I ���$���(�g-�(1���4�o�8��O<��?�2C�&zF�`�I�
�L�+�O���R��U��sX�"B[��
^���`�z�c�@_f�)i���k�"�n��q�?Rt�gw���y��o|� ��ˀ�+��SD��/x������l׆���x6���i�������݌�}��Oc��ૐ������C������ޕ��+���w��/Ù�=��LV��V����垼-���t��ý�����"W��b���! ���[���������΅��M��S��G�������s���ȵ����U`�������⺼��aZ���  �  �N=,ZN=v�M=�M=�nL=c�K=:K=�pJ=��I=�I=�iH=�G=�G=�eF=f�E=6E=�iD=}�C=�C=5uB=��A=a'A=@=-�?=@)?={>=��====�c<=��;=��:=�C:=ˏ9=��8=�-8=��7=��6=�-6=چ5=(�4=�;4=F�3=�2=lB2=B�1=T�0=5,0=�q/=9�.=��-=!*-=�_,=�+=��*=\�)=�)=�3(=�P'=�g&=�x%=&�$=z�#=�{"=Ui!=�K =�!=c�=/�=�Q=;�=ˀ==�z=2�=G=��=��=�5=Qv=��	=�=M=�;=�]=�y =^�<�<�<FO�<1V�<�R�<�E�<�0�<��<���<v��<&��<��<OU�<m*�<���<տ<R��<��<Y�<�/�<��<�צ<맢<t�<�;�<{��<,��<|�<B7�<O�<׮�<��x<mdp<�g<��_<�@W<��N<D�F<ӂ><R6<�#.<w�%<m�<�<jT<<v��;�
�;Pt�;U��;"G�;K��;N3�;��;��j;`�I;�l);
	;���:ؑ:��$:�.9u����T�u����溗��0�d�N�@�l�%�������֡�.����2��VLʻ��ֻ�>�F�=��������>��9������I �1�$�x�(��-�j#1�w5�r�8��f<�<�?�WLC�w�F���I�{�L�F�O�z�R�T�U��}X��H[�\^�(�`��c��Xf��i���k���n�/xq��;t�R�v�z�y�S|�`�~���������6���k��Ν���͆�@���<0��:e�����8܌����_e���������K��K���`镼�7������IЙ�3���b�������K5��({��O¢����X�����������W��'���d��}���⮼6H��F����
��?e�����	��IR��q����ֺ����uQ���  �  ��N=�]N=ݺM=M=�nL=��K=NK=�mJ=��I=hI=-cH={�G=�G=]F=��E=�	E=�aD=>�C=pC=pB=��A=�$A=i}@=��?=�)?=�|>==�==�==�h<=\�;=��:=}K:=`�9=��8=b78==�7=I�6=k66=��5=j�4=�A4=��3=S�2=E2=Y�1=Y�0=),0=�p/=��.=-�-=y%-=:Z,=X�+=�*=�)=I	)=C+(=tH'=K`&=�q%=�|$=#=^x"=cg!=�J ="=��=ާ=�U=-�=چ=:=�=Z�=!Q=5�=��=_@=܀=��	=/�=�=�B=�c=�~ =	&�<bB�<�R�<W�<Q�<�A�<8*�<J�<[��<���<f��<�n�<�C�<��<^��<"ſ<��<�u�<
O�<(�<���<�Ԧ<1��<�u�<�?�<��<�Ǒ<Ȇ�<LD�<m�<迀<y<Ջp<�h<��_<�gW<kO<u�F<s�><^k6<�8.<&<��<��<JW<:<���;"��;?Q�;F��;A�;�x�;��;So�;�j;�ZI;<�(;��;���:�:J1#:H*9氹�IU�D���.��+��$o0��N��zl�K�Ok�����`o��"뼻zʻ��ֻ���}��"K��Ϭ�5�y.��.�[����J ���$�U)�Y.-��61�5�=�8�.�<�)
@�ToC�l�F���I���L�9�O�*�R���U���X��R[��^���`���c��Pf�6i�t�k�G�n��_q�5t�:�v�)�y��-|��~�
����ꁼz%��G\��揅��t􇼖(���_������ڌ���th������P��1U�����������G�������ᙼ�+��s��ĸ������b@������Ȣ�����Y��Z���Z���3S���������+r���ծ�V9����������mR��禵�.���$@�������Ǻ�N��XF���  �  �O=FaN=R�M=GM=�nL=P�K=�K=�iJ=c�I=�
I=Y[H=��G=�F=�RF=e�E=��D=dXD=��C=�C=�iB=��A=� A=#{@=��?=
*?=/~>=��==�==�m<=Ѻ;=;=[T:=�9=D�8=8B8=%�7=��6={@6=B�5=��4=�H4=K�3=��2=�H2=p�1=1�0=�+0=o/=��.=��-=�-=AS,=@�+=��*=O�)=1�(=-!(=�>'=MW&=�i%=�u$=�y#=Kt"=�d!=�I =-"=`�=��=�Y=��=��=@=v�=��=w\=;�==�L=ڌ=	�	=��=�$=�J=�j=� =E.�<H�<�U�<XW�<�N�<9<�<�!�<�<*��<��<���<wZ�<�.�<��<��<1��<��<&g�<�B�<�<���<�Ц<���<�v�<tC�<��<�Б<���<�R�<��<oӀ<�,y<�p<�Mh<��_<�W<FO<� G<��><��6<�O.<�&<"�<�<%Y<�<�|�;#��;U&�;Zx�;-ζ;-�;S��;��;:Si;��H;/(;m�;\��:��:o�!:I 9����l�U�P਺�{�����@0�X]N�!"l�����*��O��)!��5�����ɻqcֻ)�⻷�� ��O��������"�: �����M �;�$�T)��@-�8N1��95�y9�>�<�2@���C���F��J�M��P��R�8�U�ўX��_[��^�n�`�֍c�If��i���k�n�9Dq���s���v�L`y�b|���~�T����Ձ����VJ��"���괆��釼b ��"Z������ڌ�B!���l���������ya��w������`Z��ϩ��E����?�������ʝ�����M��܎���Т�,���\������$����N��|������f��MǮ�D(������B䲼�<������඼�+���r��a���h����9���  �  �O=�dN=��M=M=qnL=��K=�K=eJ=h�I=bI=�RH=עG=g�F=�GF=�E=��D=�MD=�C=nC=�bB=�A=�A=@x@= �?=�)?=N>=w�==�#==s<=x�;=c;=]:=Q�9=H�8=�M8=��7=1�6=K6=�5=&�4=*P4=-�3=R�2=�K2=-�1=��0=�*0=�l/=a�.=��-=o-=wK,=Cz+=��*=��)=�(=(=4'=aM&=	a%=n$=^s#=�o"=�a!=�G =�!=y�=�=�]=��=u�=�=�=�=sh=��==�Y=��=��	=�=�.=%S=wq=q� =J6�<(M�<�W�<�V�<�J�<�5�<'�<��<R��<s��<r�<UD�<��<���<���<Y��<$y�<�V�<;5�<��<��<�˦<Y��<$w�<�F�<�<�ّ<<b�<�$�<��<~Yy<��p<n~h<y`<��W<�qO<�'G<��><��6<g.<*)&<��<�<^Y<�<�d�;ۯ�;t��;�:�;ք�;�٥;�=�;��;/�h;��G;�r';^=;���:�:q�:6c	9Mⴹ��V����������0��N���k������璻��cή��B��:Yɻ�ֻ]�:G�����v����U��������IR �B�$�� )��U-��h1��Y5�X(9� �<��]@��C�AG�f8J�GM��=P�ES���U���X��n[��$^���`���c��Bf���h���k��nn��'q�j�s�t�v�+6y���{��m~�i}��Z���9����7��p��P����އ�e���T��0���"ڌ��#��.r��1Đ����eo��Ɣ���� o��Ϳ�����HV������yޝ����]��(���Rڢ�����`��٩������zJ������f����Y��R�������s���β�D&��z���ɶ�����^������+黼H-���  �  	O=�gN=<�M={M=�mL=?�K=�K= `J=��I=��H=�IH=ɘG=�F=T<F=��E=0�D=0CD=5�C=��B=0[B=ԹA= A=�t@=,�?=@)?=�>=��==�&==�w<=��;=
;=cf:=D�9=9=�X8=��7=* 7=rU6=J�5=a5=W4=��3=\�2=�N2=q�1=��0=�)0=j/=Z�.=l�-=�-=sC,=q+=��*=��)=��(=�
(=$)'=,C&=�W%=<f$=�l#=yj"=�]!=�E =!=�=�=a=�=�=�#={�=e=#t=U�=�=�f=�=��	==�7=
[=�w=a� =M=�<2Q�<Y�<9U�<_F�<.�<��<���< ��<t��<�\�<�-�<" �<��<��<���<�e�<�E�<�&�<��<��<�Ŧ<��<�v�<�H�<g�<A�<K��<�p�<6�<���<N�y<q<��h<�K`<��W<�O<�MG<�?<��6<�|.<�8&<w�<��<�W<<[I�;��;���;���;�9�;��;6��;@S�;��g;NG;�&;6�;GC�:	�:��:qB9�A���kW��M��*��ɹ���/���M��qk�{N��Ѧ������}���� ɻ��ջ(⻲�����]�Q�����p����p���X �,�$��1)�;l-���1��z5�1N9��<���@�I�C�|<G�VeJ�;qM��cP�V@S�V�V�X��[�\0^���`���c�o>f���h�T�k��Yn��q��s�fhv�/y���{�W@~��f��ʩ��邼�%��`������Շ�L��iP������#ی��'���x��=͐��$���}��ה�/��t���W֘��#��!m��걜��򝼨0���l��O����䢼d#���e��򫦼I���ZG��������6N��﩮�����`������"��ec������� ��K��j���yڻ�|!���  �  �O=qjN=p�M=nM=7lL=��K=/K=[J=��I=.�H=AH=.�G=0�F=�1F=��E=w�D=9D=ȕC=O�B=�SB=ٳA=GA=wq@=��?=7(?=4�>=��==�)==|<=.�;=�;=dn:=H�9=�9=c8=E�7=4
7=�^6=ɳ5=�5=!]4=`�3=�3=�P2=G�1=$�0=�'0=5g/=6�.=�-=-=�;,=h+=��*=E�)=�(= (=�'=�9&=O%=�^$=hf#=`e"=Z!=FC =�=7�=��=�c=(	=��=�*=��==�~=��=�*=:r=0�=&�	=�=8@=b=�}=�� =�B�<4T�<XY�<�R�<`A�<M&�<��<=��<��<&z�<�H�<"�<���<Ⱦ�<a��<�s�< S�<H5�<��<w��<�ު<0��<3��<Wu�<rJ�<��<f�<P��<�}�<�E�<��<V�y<�Aq<M�h<hw`<4X<i�O<pG<W"?<��6< �.<�E&<��<��<�S<�<�,�;�_�;���;ݻ�;&�;>2�;���;���;
g;�\F;�%;&�;M
�:'Ԍ::�p�8�����KX��������ײ�[�/���M�Q'k����Tl��
v��4��,����ȻLmջp����cU��(F����&��k����_���` ���$�LC)���-�6�1�:�5��r9��%=��@� D�LhG��J� �M�O�P��`S�^'V���X��[��<^�'�`�'�c��;f�g�h�?�k�jGn�V�p��s��Fv��x��{�4~�qR������ւ�����R��J���ḋ�[��0M��Ғ���܌��+��.��m֐��0��&����甼�A�������똼�9��ł���Ɯ�,��FB���{������#+���j��ݮ������5E�����G쫼!D��0�������PO�����������N��V���f�w9��߃��nͻ����  �  �O=MlN=-�M=M=�jL=E�K=�	K=bVJ=�I=}�H=q9H=��G=�F=(F=}E=�D=0D=��C=��B=�MB=u�A=�A=6n@=��?='?=�>=��==�+==N<=��;=w#;=u:=��9=9=�k8=��7=�7=�f6=�5=�5=#b4=7�3=f3=R2=��1=u�0=&0=zd/=]�.=#�-=-=�4,=J`+=^�*=!�)=��(=��'=�'=�0&=\G%=�W$=�`#=�`"=�V!=�@ =�=
�=��=
f=y=,�=y0=�="!=��=U�=�4=|=Ǻ=�	=�=G=�g=�=� =G�<V�<�X�<P�<v<�<��<X��<P��<֜�<j�<�6�<G�<g��<L��<h��<�a�<�B�<�&�<P�< �<�֪<.��<O��<�s�<$K�<��<��<���<3��<�R�<��<!�y<�eq<3�h<K�`<^=X<��O<��G<�:?<l�6<y�.<VO&<��<�<�O<#�<o�;�:�;{_�;��;��;c�;�9�;ݣ�;q\f;]�E;�[%;�I;���:�:<w:z�8bɻ�FY�(ک������O�/��M���j����[;��d=��z���\^��6rȻ),ջ�Ỳ��M'��P3�^�����}�
��	��th �j�$�}S)�	�-���1���5���9�I=�e�@�{FD�ʎG�@�J�v�M�\�P�^}S��?V��X�7�[�H^���`�x�c��:f��h�e�k��8n���p�E�s��*v���x�'a{�~�}�A��W����ǂ����G������Ň�����J��˒��ߌ�0��n����ސ�!;��̘��\���R������j����L�������؜�>���Q����������h���h2���o��򱦼�����C�������櫼�;�������鯼�@��j����과c=�����ݷ��*���v���»�����  �  O=�mN=��M=�M=�iL=-�K=�K=�RJ=��I=2�H=�3H=#�G=�F=� F=�uE=��D=)D=�C=!�B=\HB=!�A=aA=zk@=��?=�%?=�>=��==W-==��<=��;=�';=z:=��9=?9=>r8=��7=7=�l6=C�5=i5=�e4=��3=A3=S2=��1=��0=�$0=b/=;�.=4�-=X-=,/,=0Z+=��*=�)=e�(=i�'=�'=E*&=SA%=ZR$=\#=�\"=�S!=�> =j=��=�=�g=�=��=�4=.�=='=q�=��=�;=��=��=��	=�%=DL=l=E�=9� =�I�<�V�<!X�<�M�<8�<��<���<���<���<�]�<')�<���<N��<?��<�u�<�S�<26�<K�<a�<��<Ъ<+��<��<&r�<=K�<� �<��<�<)��<�\�<w(�<f�y<��q<i<�`<�WX<�O<$�G<�L?<��6<٧.<V&<�<D�<^K<M�<���;��;>:�;�W�;�}�;��;��;�d�;�e;�7E; �$;��;�&�:�"�:u-:���8>���i�Y����_����b�/�XcM��j�3؃�G������ƭ��,��@Ȼ��Ի�\ứ_���W%�*��/��F��������;o ���$��`)�W�-�?�1��5���9��d=��@�7dD���G���J���M�i�P�ēS��SV�QY�B�[�#R^�[�`�Жc�;f���h�i�k�.n�f�p�pvs��v�=�x�H{�Y�}�4���x����������>��2����������I��G���ጼ�3�������吼�C��󢓼����^��]�������[��h���&眼�$���]��S����ɡ�����b8��Xt�����������C��8����⫼�5���i௼�5��c����ݳ�J0��8����з����Hm������r���  �  SO=BnN=��M=9M=�hL=ƷK=�K=XPJ=��I=��H=�/H=�{G=��F=	F=�pE=�D=�$D=�C=`�B= EB=`�A=!	A=�i@=y�?=%?=�>=��==,.==�<=��;=,*;=)}:=�9=$#9=\v8=��7=7=hp6=��5=55=h4=��3=_3=�S2=��1=*�0=�#0=�`/=0�.=��-=W�,=�+,=7V+=j~*=��)=��(=��'=#
'=&&=g=%=�N$=Y#=�Z"=�Q!=l= =�=`�=W�=Oh=P=��=i7=d�=�*=��=�=�@=7�=Y�=��	=O)=cO=�n==�=�� =SK�<RW�<LW�<�K�<5�<��<}��<���<���<\U�<d �<D��<���<���<ol�<K�<.�<�<��<��<�˪<ﰦ<В�<q�<EK�<�!�<a��<&ƍ<��<�b�<�/�<m�y<�q<�,i<L�`<hX<
P<�G<_W?<7<!�.<�Y&<�<G�<H<��<4��;�	�;7"�;�;�;>]�;:��;z֓;�;�;e;b�D;�$;��;��:^��:^:�a�8���[5Z��:��l纇���/��PM�ߡj��Ń���������!���8���Ȼ��Ի�?�`F�=�������,�������N���s �8�$�)i)���-���1�f�5��9��u=��	A�QwD���G���J�F�M���P�$�S��_V��Y���[��X^���`�_�c�c;f���h�=�k��'n���p��ks��v�y�x�8{���}��+��q��ش��w���a9��2{���������I�������⌼#6��A���1ꐼ�H��O���1	��g�����7��:e��孛�1�	-��{e������ϡ����R<��Dw����������YC������ૼm2��=����گ��.��Ȃ���ճ��'��y��Rɷ����fg��굻�����  �  �O=paN=�M=�M=JZL=��K=�J=	EJ='�I=<�H=�)H=UwG=��F=F=�kE=�D=�D=�uC=��B=�.B=u�A=��@=�E@=�?=�>=�Q>=H�=={�<=`N<=G�;=w�:=+B:=��9=�8=@38=k�7=m�6=+#6=hr5=��4=j4=gZ3=u�2=�1=�01=r0=Ư/=v�.=&.=�P-=,=ҩ+=a�*=$�)=)=?7(=dS'=�k&=��%=ҏ$=�#=�"=��!=o� =�i={C==
�=.�=�-=9�=|V=��=2O=��=H=�q=�=�=�>	={r=�=��=��=���<)�<#9�<�G�<oK�<E�<�5�<��<��<M��<��<��<r�<#O�<�.�<��<V��<>޺<1ȶ<���<
��<���<'p�<�U�<;8�<��<?��<4Α<�<|�<�P�<0%�<��y<�q<�Di<��`<��X<NP<� H<��?<�m7<�&/< �&<K�<,K<��<ͪ<e��;.��;7J�;ԝ�;���;�d�;+�;}�;�hl;�L;D	,;
@;ps�:�:v�9:v�x9(�q��\6�������Ӻ)���b%���B�P�_�{|�����䙻*l�����A���9λl�ڻ�w���bX��K#�:p	�������j���-�!�N"&�.r*���.���2�0�6� ^:�r>�ăA���D��#H��FK��ON��BQ�%#T�U�V��Y�d}\�P9_��a�תd��ag��j���l��}o��,r���t�w�P"z�O�|�U\����� D�����DՄ�\���e��ӯ������J�����������H������� ��=^������F��p��NŘ�����a������일	,���i��Φ��䢼�"��Vd��
���C��<��͋��3ݫ��0��D����گ�0��:����ٳ��-��ʀ��ӷ��$��v��@ǻ����  �  lO=HaN=�M=	M=xZL=F�K=��J=�EJ=�I=�H=�*H=]xG=��F=/F=mE=N�D=�D=�vC=��B=�/B=8�A=C�@=[F@=!�?=@�>=�Q>=8�==H�<=�M<=��;=��:=fA:=Ǒ9=�8=>28=b�7=q�6=6"6=�q5=/�4=�4=�Y3=(�2=��1=�01=?r0=��/=��.=�.=�Q-=�,=��+=]�*=+�)=,)=_8(=�T'=m&=��%=͐$=��#=ʛ"=*�!=� =�i=�C==��=��=&-=��=�U=��=6N={�==�p=��=�=�=	=yq=#�=��=B�=���<��<�8�<�G�<�K�<�E�<�6�<��<.�<���<���<��<ft�<lQ�<�0�<H�<���<\�<ʶ<ϴ�<���<1��<q�<OV�<�8�<��<,��<�͑<��<�z�<hO�<q#�<��y<Җq<*@i<��`<l�X<JP<P�G<T�?<Ok7<�$/<��&<��<K<�<��<h��;���;1P�;|��;��;gm�;��;#��;3|l;�*L;�,;PS;��:�:��9:Yy9�Sq��>6�j���}�Ӻ����b%�8�B�;�_��&|����뙻�r��(�������'@λY�ڻ�}�@��\���$�1q	�Ӕ����Zi�����!� &�]o*�V�.�_�2�%�6��Y:���=�'A��D�LH�kBK��KN��>Q��T���V�ǺY��{\�m8_�_�a��d�jbg��j���l�"�o��/r�/�t�؂w�6&z�i�|�e`������E�������ք�}���f��G�������J��j������H������#����\������;���m�������i_������ꝼ*��h��6����⢼�!���c��������<������ݫ��1������,ܯ��1��-����۳��/��ǂ���Է�t&���w���Ȼ����  �  X
O=�`N=��M=2	M=[L=F�K=��J=^GJ=�I=��H=~-H=p{G=�F=�F=wpE=��D=/D=�yC=v�B=62B=B�A=��@=�G@=
�?=��>=�Q>=�==��<=�L<=+�;=��:=	?:=�9=�8=8/8=T7=v�6=e6=o5=�4=4=�X3=5�2=k�1=�01=�r0=��/=��.=(!.=vS-=�,==�+=B�*=F�)=�)=�;(=�W'=tp&=��%=��$=s�#=�"=�!=F� =�j=&D=5=��=0�=�+=��=�S=<�=MK=8�=�=m=!�=L�
=<:	=�n=��=��=��=��<��<�7�<�G�<�L�<jG�<?9�<u#�<z�<	��<���<X��<B{�<mX�<8�<7�<��<��<�϶<���<���<���<�s�<X�<�9�<��<:�<�ˑ<\��<(w�<�J�<!�<��y<1�q<+3i<��`<ՌX<V>P<��G<q�?<.d7<�/<��&<n�<�J<��<ٮ<���;��;a�;}��;��;M��;�	�;आ;��l;�gL;�W,;ӊ;%��:�^�:qf::�}{9σo���5�ߓ��i�ӺT��Ph%���B���_�}A|�E/������B���tǴ�T���lVλl�ڻN��E)�i���)��t	�t������g�v�۪!��&��g*�&�.��2�F�6�0M:�#�=�,qA��D��H��5K��?N�m4Q��T���V���Y�-w\�d5_���a�"�d�Ddg�nj���l��o�8r��t��w�2z���|��l����`K��s����ڄ��!��2i��㱈������I��u���`qE��Y���(����W��S���6���g��������X������㝼a$��c��ߠ��7ߢ����a��a�����m=��P����߫�r4��D����௼�6��録��᳼�5��ˈ���ڷ��+��|��b̻����  �  �O=�_N=9�M=h	M=�[L=��K=�J=JJ=`�I=q�H=�1H=K�G=1�F=�!F=�uE=�D=K$D=[~C=��B= 6B=m�A={�@=�I@=]�?=u�>=�Q>=T�==E�<=�J<=��;=��:=3;:=Ȋ9=u�8=R*8=oz7=��6=�6=�j5=��4=	4=\V3=��2=��1=x01=�r0=��/=��.=g#.=ZV-=��,=E�+=��*=2�)=�!)=A(==]'=�u&=|�%=�$=e�#=N�"=��!=U� =gl=�D=H=	�=�=�)=F�=2P='�=�F=�=-=pg=s�=��
=!5	=�i={�=[�=��=���<@�<�6�<�G�<�M�<,J�<d=�<�(�<]�<��<���<d��<��<�c�<C�<%�<h	�<�<"ض<��<ݩ�<���<Ww�<�Z�<�:�<��<��<�ȑ<���<q�<|C�<��<��y<�uq<[i<��`<�xX<�+P<\�G<*�?<�X7<0/<��&<X�<BJ<� <׳<	��;"�;�{�;���;�=�;X��;�5�;8ӆ;3m;��L;s�,;��;6��:�:>`;:F�~9S�l��c5��g��ʵӺ<���r%���B�O�_��m|�~J����������봻���tzλ��ڻٮ滕C�Q���1��y	�A��ˑ�ve�����!�Q&��[*���.�R�2��t6�9:���=�d[A�<�D�n�G��!K�p-N��#Q�KT���V�+�Y�.p\��0_���a���d�dgg�E"j�t�l�M�o��Er��t���w�Ez�0�|�!�����S��?���]ᄼ'��/m�����������I��9����덼�A��\�������tP��ԫ�����W]��|�������M������ڝ�w��&[�� ����٢�����^������
�>��[���J㫼99��[����篼K?�������볼�?�������㷼4�������һ��!���  �  'O=�]N=��M=�	M=�\L=��K=��J=�MJ=��I=c�H=�7H=��G=��F=�(F=�|E=��D=�*D=t�C==�B=�:B=n�A=��@=L@=��?=<�>=�Q>=j�==~�<=GH<=�;=@�:=6:=�9=I�8=�#8=�s7=W�6=6=�e5=ݵ4==4=QS3=��2=;�1= 01=Us0=��/=��.=?&.=�Y-=�,=k�+=��*=�*=_()=�G(=d'=@|&=ȏ%=͝$=l�#=��"=�!=� =n=�E=A=�=�=6'=��=�K=��=h@=Q�=�	=�_=��=��
=[.	=�c=�=ƹ=!�=j��<�<�4�<�G�<�O�<�M�<�B�<�/�<�<q��<���<l��<���<�q�<SQ�<�2�<��<��<�<wʲ<ñ�<ɗ�<�{�<d]�<�;�<�<�<cđ<f��<�h�<�9�<$
�<��y<�Zq<�i<O�`<�^X<GP<u�G<h�?<�H7<9
/<y�&<��<I<^<��<���;�<�;���;r�;�l�;6�;_o�;4�;��m;�?M;8*-;�P;i�:��:�<:�z�9�i�t�4��3����Ӻg����%���B�� `��|��n��UG��Dا�:���»B�λ��ڻ���sf�>���=���	����Ւ�3c���!�E&�{L*��s.�$y2�]6�:���=�9?A��D��G��K��N��Q�/�S���V�E�Y��g\�o+_���a���d�8lg�q*j�*�l�v�o��Wr�p
u�+�w�K^z��|��������_������!ꄼR.���r��B�������AJ��ߗ���荼=�����푼G���������/P��ţ�����?��=���p͝���Q�������Ң�}���Z��p����識N?��U����竼�?��k�����^J�����P����L��Z����M?��X����ڻ��(���  �  O=�[N=s�M=q	M=�]L=Y�K=iK=8QJ=?�I=��H=�=H=��G=��F=�0F=�E=��D=j2D=e�C=��B=,@B=�A==�@=�N@=��?=��>=nQ>='�==9�<=E<=ɓ;=�:=0:=O~9= �8=J8=Hl7=�6=�6=5_5=@�4=� 4=�O3=Ĝ2=��1=C/1=�s0=�/=��.=X).=�]-=�,=@�+=�*=�*=0)=�O(=l'=�&=�%=H�$=#�#=S�"=�!=�� =�o=�F==��=�=�#=,�='F=L�=9=N�=n=:W=A�=!�
=\&	=h\=��=P�=��=���<��<"2�<�F�<Q�<2Q�<SH�<�7�<� �<C�<"��</��<���<*��<�a�<�B�<�%�<�	�<Z�<ղ<b��<���<���<1`�<�<�<��<��<ž�<���<_�<�-�<���<̘y<N;q<4�h<
�`<�?X<S�O<U�G<�r?<667<��.<��&<L�<G<f<E�<���;bZ�;���;�/�;ݢ�;�!�;Ű�;uT�;6 n;��M;�-;��;�R�:�s�:��=:FŃ9��e� 4�e���?�Ӻ����%��C�9`�w�|�g���y����%U���G»��λ#ۻ��Ɛ�i����J��	�n��Ӕ�[a��
���!�!�%��;*�_.�a2�B6��:�0�=��A��~D���G�	�J���M���P���S��V�C�Y��^\�?&_�}�a�b�d��rg��4j���l���o�nr��#u��w��{z��}�d��.&��4m��Ա����7��dy��������	K��Ŗ���卼 8��6���M䑼x<�������땼JA�������㙼�/���x�� ������E�� ���ˢ�����V��|����識6A��0������G��B���*���pW��K���S��	\��k���l����L������仼�0���  �  ��N=xYN=�M=	M=h^L=�K=)K=UJ=�I=��H=�DH=�G=��F=O9F=~�E==�D=]:D=��C=�B=�EB=��A=��@=$Q@=�?=T�>=�P>=��==��<=AA<=�;=9�:=h):=�v9=�8=�8=�c7=��6=C6=.X5=�4=M�3=gK3=��2=p�1=0.1=�s0=�/=��.=_,.=b-=�,=E�+=�*=U*=!8)=5X(=Nt'=�&=t�%=�$=�#=@�"=��!=y� =�q=G=v=1�=}=�=1�=@=/�=1=��=/�=�M=��=��
=�	=pT=��=F�=��=���<A�<�.�<�E�<6R�<�T�<�M�<�?�<	+�<|�<L��<���<F��<k��<"s�<�S�<�5�<��<��<�߲<<î<O��<S��<�b�<�<�<��<��<H��<���<T�<� �<��<xy<�q<��h<�j`<sX<��O<��G<�Y?<j!7<��.<�&<�}<�C<�<�<��;�x�;i��;�_�;{۸;_a�;��;���;9�n;�`N;@.;V;�E�:�I�:eo?:�9�Eb��y3��Ж��}Ӻ����%�-FC�^y`�:D}��ʌ�鯚�-J�������»| ϻ�]ۻK=绱������\Z��	�������`�����!�4�%��**��I.�LH2��%6�s�9�=���@��\D�c�G���J�&�M���P�n�S��V�w�Y��U\��!_��a�%�d�_zg�Aj��m�+�o�n�r�O?u���w�V�z�'?}����;6��4|��W���� ���@��"�������}L�����㍼G3��[���Mۑ��1��և��uݕ��1��R����ҙ�����h�����t����9��~��.â��	��OS��ퟦ���C��Ț������WP��.����	���e����������l��ྶ�6��[�����𻼲9���  �  ��N=�VN=f�M=vM=�^L=��K=�K=�XJ=��I=e�H=+KH=i�G=z�F=�AF=��E=k�D=,BD=�C=X�B=&KB=�A=�@=bS@=I�?=��>=�O>=��==��<=H=<=�;=L�:=�":=Ho9=�8=�8=m[7=r�6=e�5=�P5=��4=��3=�F3=;�2=�1=�,1=9s0=ܵ/=��.=./.=�e-=�,=&�+=��*=�*=@)=l`(=�|'=Փ&=إ%=��$=Ŷ#=�"=`�!=�� =�r=mG=�=O�=
z=�=��=�9=�=�(=��=��=D=�=��
=�	=HL=U}=�=x�=���<>�<�*�<TD�<�R�<�W�<3S�<CG�<�4�<l�<�<:��<���<w��<+��<[d�<!E�<�&�<{�<Z�<�ˮ<z��<c��<�d�<�<�<H�<��<T��<�}�<�H�<Y�<�ހ<�Vy<��p<��h<�F`<��W<.�O<fxG<	@?<�7<w�.<֧&<�t<�?<�<��<k�;
��;�;���;��;ҟ�;n:�;]�;�Ho;f�N;��.;�;�2�:��:�@:%Q�9w�^���2���� zӺ�����%�VyC��`�{�}�����6蚻���zӵ���»�_ϻ��ۻ;t�������j�d�	�/��a���`�����!�(�%�9*��5.�02�
6���9��^=��@��:D��G�%�J�p�M�Z�P�%�S���V��yY��M\�_���a�طd�W�g��Mj�!m�r�o�e�r��[u��x�a�z�a}�����F������A̓����K��P����Ȉ�
��cN�������/������ґ��&��Y{��Rϕ�"��s������m���X��:���9螼s.���t��˻�����*P��Ԟ����F�����������Y��o������t���ϲ�u(���}���϶�F���i��^���z���IC���  �  /�N=TN=��M=�M=�^L=��K=�K=�[J=��I=y�H=QH=�G=��F=IF=��E=��D=HID=`�C=�B=PB=ħA=�@=@U@=.�?=p�>=�N>=��==��<=h9<=)�;=��:=�:=h9=-�8=�8=]S7=��6=��5=J5=��4=��3=�B3=Ւ2=��1=j+1=�r0=H�/=��.=�1.=`i-=C�,=y�+=��*=�"*=OG)=�g(= �'=�&=��%=��$=��#=%�"=��!=#� =
t=sG=�=S�=w=�=�=�3=�=,!=?�=��=�:=��=��
=h	=�D=hv=��=x�=���<4 �<'�<[B�<S�<�Y�<�W�<�M�<�=�<?(�<��<?��<���<��<���<ts�<HS�<c3�<��<��<�Ү<ư�<���<�e�<�;�<x�<�ݕ<d��<�t�<�=�<g�<Ѐ<j7y<9�p<�xh<�$`<B�W<��O<^\G<a'?<��6<��.<��&<�k<�:<G<��<p'�;��;�2�;���;�D�;�ب;�x�;0'�;�o;�wO;&M/;TP;�
�:֟:mB:F�9$\��q2�����JӺ���\�%��C�la��}��,��������:���û�ϻ?�ۻf�给�7��N{��	���J��b�L��Nz!���%��*�r#.�2���5��9��@=�Y�@�D�bG�=�J�T�M�X�P���S�u�V�,oY��G\��_�;�a�(�d���g�[j�(m��o���r��vu�@.x���z�9�}����V��	����ڃ�X���T��K����Έ�T���P��U���Oߍ��+��Xz��Kˑ�r��p�������d��w���J���;J��Ɠ��9ܞ�$��Sl��_���S ���M��[���}�.J��F������b��Uî��#�������޲�^8��捵��߶�p-��x��'�������L���  �  ��N=yQN=�M=�M=�^L=b�K=`
K=.^J=!�I=�I=VH=��G=��F=�OF=
�E=I�D=JOD=�C=��B=TB=�A=OA=�V@=ê?=1�>=�M>=��==��<=�5<=܀;=w�:=G:=�a9=n�8=��7=[L7=��6=k�5=D5=+�4=��3=�>3=��2=X�1=�)1=r0=y�/=��.={3.=l-=ߠ,=��+=�*=G(*=tM)=En(=X�'=/�&=?�%=ּ$=<�#=��"=�!=Ȗ =�t=OG=�=]�=;t=$=i�=t.=ة=f=߀=(�=�2=	�=��
=	=�==Wp=��=��=S��<���<1#�<c@�<�R�<q[�<:[�<YS�<�D�<91�<M�<��<{��<J��<���<;��<9_�<>�<��<K��<�خ<�<��<if�<�:�<��<6ٕ<���<�l�<�3�<��<_À<�y<?�p<�Zh<�`<��W<�|O<DG<�?<�6<&�.<Վ&<�c<�5<<��<4�;0��;�N�;���;o�;	�;���;O_�;.Bp;v�O;��/;��;Y��:.q�:�C:׋9,�Y�o2����ՋӺ��!&���C��=a�o4~��V��M�����E��X:ûC�ϻvܻO�继G��Z�������	�?������c����yu!���%�_ *�i.��2���5���9��'=�C�@� D��HG��xJ��M�3�P��S���V�gY�C\��_�U�a���d�B�g� gj�67m�Fp���r���u�EHx��z�;�}�����c��Φ��惼�"���]������rԈ�S��S�����Oލ��(���u��!ő�����f���������eW������g��=��i���%Ҟ����_e��0�������L��O���"���|M��*����	���j���̮��.��ˎ��B첼*F��웵�u��:��z���M˺�c���T���  �   �N=rON=u�M=�M=�^L=еK=�K=�_J=��I=�I=�YH=�G=` G=eTF=�E=�D=�SD=�C={ C=WB=L�A=�A=�W@=
�?=��>=�L>=)�==��<=3<=r};=z�:=�:=�\9=<�8=1�7=�F7=j�6=Y�5=l?5=�4=F�3=�;3=E�2=��1=�(1=yq0=y�/=��.=�4.=n-=��,=$�+=�+=�,*=R)=s(=$�'=ͥ&=}�%=��$=u�#=8�"=��!=� =<u=
G=�=��=�q=D=ܣ=A*=�=!=/{=6�=�,=�y=�
=n�=�8=�k=��=|�=���<M��<! �<�>�<rR�<�\�<�]�<`W�<wJ�<8�<Q!�<��<+��<A��<��<ډ�<(h�<7F�<�#�<� �<ݮ<෪<���<�f�<�9�<	�<sՕ<Ӟ�<f�<,�<0�<q��<Ry<۠p<�Ch<��_<��W<�gO<�0G<� ?<��6<�.<��&<�\<�1<�<U�<�<�;���;�c�;C��;��;�-�;�՘;뉈;��p;�?P;50;c;#F�:�:�C:c��9`>X�@�1�bw��p�Ӻ�#�k9&��D�0na��n~�Ax��r��r��n��-dû��ϻd+ܻL���g��v�������	���ڪ��e�L��[r!���%���)�&	.�_�1���5�9��=�~�@�E�C��5G�gJ��M���P���S�]{V�[aY�@\�4_�S�a�Q�d�S�g��pj�?Cm��p�m�r�(�u�d\x�{���}��&��n������&�*���d��P����؈����U�������ݍ� '���r����������_��r�������M�������蚼�4������ʞ�-��5`��s���p����J����������4P��������Jq���Ԯ�U7��^��������P��ߦ��'���E��%���Ժ�"��b[���  �  l�N=NN={�M=YM=�^L=�K=3K=aJ= �I=�I=\H=��G=FG=iWF=��E=E=�VD=��C=�C=�XB=��A=�A=FX@==�?=��>==L>=�==S�<=B1<=B{;=��:=�:=�Y9=�8=��7=qC7=��6=(�5=l<5=E�4=��3=�93=��2=<�1=�'1=q0=t�/= �.=�5.=To-=/�,=.�+=F+=I/*=�T)=v(= �'=��&=2�%=�$=q�#=��"=�!=�� ={u=�F==��=~p=d=��=�'=�=�=�w=d�=�(=v=8�
=��=N5=�h=��=J�=��<o��<(�<�=�<FR�<7]�<Y_�<�Y�<�M�<E<�<N&�<��<6��<|��<D��<��<�m�<*K�<(�<X�<�߮<���<b��<�f�<�8�<Z�<�ҕ<|��<�a�</'�<~�<��<��x<h�p<?5h<2�_<��W<�ZO<�$G<�><W�6<��.<T&<RX</<�<X�<B�;��;Vp�;��;�;�D�;��;Y��;��p;uP;�>0;h0;4��:�,�:�8D:��9|KW�P�1�|u��)�Ӻ�0��L&��D��a�ԓ~���������5�������~ûMлDܻr軎|�Ո������	����ܭ�9g����p!�7�%���)�p.���1��5��s9��=�>�@� �C��)G��[J�#zM��P�܄S�KvV��]Y�P>\�_���a�j�d�.�g��vj��Jm��p���r�
�u�ix��{���}�}-���t���������/��i�������ۈ����|V��[����ݍ��%���p��㽑�+��9[��e���d����G�������⚼�.���z���Ş�:��"]��+�������[J����������R��ǰ��#��ju��gٮ��<��v��������W��ŭ��
����K��F����ٺ����_���  �  ��N=�MN=5�M=-M={^L=$�K=^K=oaJ=��I=]	I=�\H=s�G=>G=gXF=�E=E=�WD=r�C=rC=|YB=2�A=HA=eX@=B�?=��>=L>=ș==��<=�0<=uz;=�:=�:=�X9=��8=��7=PB7=ϓ6=�5=f;5=_�4=�3=�83=�2=��1=�'1=�p0=q�/=�.=�5.=�o-=��,=��+=+=40*=�U)=w(=!�'=��&=�%=��$="�#=N�"=}�!=٘ =�u=�F=�=q�=	p=�=͠=�&=�=�=pv=�=�'=�t=��
=��=;4=�g=�=��=��<���<��<;=�<DR�<g]�<�_�<�Z�<O�<�=�<	(�<��<9��<���<Q��<��<�o�<�L�<q)�<p�<s�<���<y��<pf�<<8�<��<�ѕ<:��<C`�<d%�<��<簀<��x<g�p<�0h<<�_<הW<rVO<� G<��><�6<�.<}&<<W<e.<�<��<FD�;~��;u�;��;���;pL�;O��;$��;��p;��P;�O0;�?;-��:�C�:�]D:�ۍ9�W�Y�1�x��A�ӺA5�ST&��$D���a�h�~�����ᑛ�>��󑶻Їû�л�Lܻ�軪��9�������	�3������g�	��p!�1�%� �)� .�	�1�Ҿ5�p9��=�#~@���C��%G�XJ��vM��P�y�S�}tV��\Y��=\��_���a�Q�d���g�	yj��Mm�5p���r��u�Tmx�k{�^�}��/��w����������1���j��Q����܈�y���V�������ݍ��%��Gp��鼑��
���Y������x����E�����������,���x��QĞ����\��h�������?J��ݞ�������R������N���v��ۮ��>������=���Z�����d���M��V����ۺ����(a���  �  l�N=NN={�M=YM=�^L=�K=3K=aJ= �I=�I=\H=��G=FG=iWF=��E=E=�VD=��C=�C=�XB=��A=�A=FX@==�?=��>==L>=�==S�<=B1<=B{;=��:=�:=�Y9=�8=��7=qC7=��6=(�5=l<5=E�4=��3=�93=��2=<�1=�'1=q0=t�/= �.=�5.=To-=/�,=.�+=F+=I/*=�T)=v(= �'=��&=2�%=�$=r�#=¿"=�!=�� =}u=�F==��=�p=k=��=�'= �=�=�w=x�=)=(v=U�
=�=p5=�h=$�=r�=W��<���<|�<�=�<�R�<�]�<�_�<Z�<N�<s<�<s&�<��<D��<���<<��<ҏ�<�m�<K�<�'�< �<o߮<Z��<��<Jf�<P8�<�<�ҕ<;��<�a�<�&�<S�<���<��x<Q�p<?5h<G�_<ęW<[O<3%G<~�><��6<�.<�&<�X<�/<l<��<�C�;��;@q�;��;���;E�;�;}��;z�p;�tP;�=0;</;4��:)�:q0D:��9�sW���1�{��ҪӺ�3��O&��D���a�^�~�*���Њ��6�������ûл�Dܻ�}�D���I����	�������Qg�#���p!�D�%���)�x.���1��5��s9��=�@�@��C��)G��[J�$zM��P�܄S�KvV��]Y�P>\�_���a�j�d�.�g��vj��Jm��p���r�
�u�ix��{���}�}-���t���������/��i�������ۈ����|V��[����ݍ��%���p��㽑�+��9[��e���d����G�������⚼�.���z���Ş�:��"]��+�������[J����������R��ǰ��#��ju��gٮ��<��v��������W��ŭ��
����K��F����ٺ����_���  �   �N=rON=u�M=�M=�^L=еK=�K=�_J=��I=�I=�YH=�G=` G=eTF=�E=�D=�SD=�C={ C=WB=L�A=�A=�W@=
�?=��>=�L>=)�==��<=3<=r};=z�:=�:=�\9=<�8=1�7=�F7=j�6=Y�5=l?5=�4=F�3=�;3=E�2=��1=�(1=yq0=y�/=��.=�4.=n-=��,=$�+=�+=�,*=R)=s(=$�'=ͥ&=}�%=��$=v�#=9�"=��!=� =@u=G=�=��=	r=Q=�=U*=+�===P{=\�=-="z=:�
=��=�8=�k=�=ɿ=N��<���<� �<U?�<S�<]�<E^�<�W�<�J�<f8�<�!�<1�<H��<H��<���<���<�g�<�E�<v#�<� �<�ܮ<\��<���<	f�<�8�<��<�ԕ<V��<�e�<�+�<��<2��<�y<��p<�Ch<��_<�W<ihO<�1G<|?<x�6<�.<��&<�]<�2<�<r�<�>�;���;ke�;���;X��;r.�;!֘;0��;n�p;�>P;�	0;!�;W@�:ߠ:��C:�Ռ9�X���1����`�Ӻs)��>&�JD�Vsa��s~��z��)t��l���o���eûN�ϻ�,ܻj���h��w�����	�B�����e�q��yr!���%���)�6	.�l�1���5� 9��=���@�I�C��5G�gJ��M���P���S�^{V�\aY�@\�4_�S�a�Q�d�T�g��pj�?Cm��p�m�r�(�u�d\x�{���}��&��n������&�*���d��P����؈����U�������ݍ� '���r����������_��r�������M�������蚼�4������ʞ�-��5`��s���p����J����������4P��������Jq���Ԯ�U7��^��������P��ߦ��'���E��%���Ժ�"��b[���  �  ��N=yQN=�M=�M=�^L=b�K=`
K=.^J=!�I=�I=VH=��G=��F=�OF=
�E=I�D=JOD=�C=��B=TB=�A=OA=�V@=ê?=1�>=�M>=��==��<=�5<=܀;=w�:=G:=�a9=n�8=��7=[L7=��6=j�5=D5=+�4=��3=�>3=��2=X�1=�)1=r0=y�/=��.={3.=l-=ߠ,=��+=�*=G(*=tM)=En(=X�'=/�&=?�%=׼$=>�#=��"=�!=̖ =�t=VG=�=i�=Jt=7=��=�.=��=�=�=^�=83=N�==�
=k	=4>=�p=#�=k�=5��<���<$�<EA�<�S�<@\�<�[�<T�<�E�<�1�<��<`��<���<S��<��<��<�^�<�=�<d�<���</خ<9��<B��<�e�<�9�<�
�<xؕ<G��<�k�<Y3�<���<À<;y<��p<�Zh<�`<�W<t}O<�DG<�?<_�6<��.<U�&<e<m7<�<��<7�;���;.Q�;���;�p�;s
�;z��;�_�;�Ap;7�O;~�/;T�;&��:Qg�: �B:w��9�BZ��62�����L�Ӻ���%&�+�C�Ea�_;~�:Z��P�������G���<ûO�ϻEܻ���I��[��q���	����Ц� d����u!���%�{ *��.�2���5���9��'=�J�@�D��HG��xJ��M�5�P��S��V�gY�C\��_�U�a���d�B�g� gj�67m�Gp���r���u�EHx��z�;�}�����c��Φ��惼�"���]������rԈ�S��S�����Oލ��(���u��!ő�����f���������eW������g��=��i���&Ҟ����_e��0�������L��O���"���|M��*����	���j���̮��.��ˎ��B첼*F��웵�u��:��z���M˺�c���T���  �  /�N=TN=��M=�M=�^L=��K=�K=�[J=��I=y�H=QH=�G=��F=IF=��E=��D=HID=`�C=�B=PB=ħA=�@=@U@=.�?=p�>=�N>=��==��<=h9<=)�;=��:=�:=h9=-�8=�8=]S7=��6=��5=J5=��4=��3=�B3=Ւ2=��1=j+1=�r0=H�/=��.=�1.=`i-=C�,=y�+=��*=�"*=OG)=�g(=�'=�&=��%=��$=��#=(�"=��!=(� =t=|G=�=a�=w=�=�=�3=�=]!=y�="�=1;=E�=�
=�	=E=�v=�=��=���<M�<(�<oC�<T�<�Z�<�X�<�N�<e>�<�(�<�<���<���<'��<���<5s�<�R�<�2�<�<��<Ү<⯪<���<�d�<�:�<��<�ܕ<���<�s�< =�<��<�π<�6y<��p<�xh<E%`<��W<j�O<y]G<�(?<(�6<:�.<��&<�m<�<<@<�<+�;k��;�5�;6��;G�;qڨ;�y�;�'�;��o;dvO;hJ/;iL;� �:�ɟ:��A:&�9��\�'�2�x���;�Ӻo��&�Q�C�V
a���}��0��r!���Ĩ�X���ûc�ϻu�ۻV��G � 9���{�x�	�q�����Xb�����z!���%�*��#.�(2��5�(�9��@=�b�@�D�bG�B�J�X�M�[�P���S�w�V�-oY��G\��_�<�a�)�d���g�[j�(m��o���r��vu�@.x���z�9�}����V��	����ڃ�X���T��K����Έ�T���P��U���Oߍ��+��Xz��Kˑ�r��p�������d��w���J���;J��Ɠ��9ܞ�$��Sl��_���S ���M��[���}�.J��F������b��Uî��#�������޲�^8��捵��߶�p-��x��'�������L���  �  ��N=�VN=f�M=vM=�^L=��K=�K=�XJ=��I=e�H=+KH=i�G=z�F=�AF=��E=k�D=,BD=�C=X�B=&KB=�A=�@=bS@=I�?=��>=�O>=��==��<=H=<=�;=L�:=�":=Ho9=�8=�8=m[7=r�6=e�5=�P5=��4=��3=�F3=;�2=�1=�,1=9s0=ܵ/=��.=./.=�e-=�,=&�+=��*=�*=@)=l`(=�|'=֓&=٥%=��$=Ƕ#=��"=d�!=� =s=wG=�=`�=z=�=�=�9=�=!)=��=�=]D=q�=��
=8	=�L=�}=��=�=���<w�<6,�<�E�<T�<�X�<8T�</H�<�5�<�<��<���<���<���<��<d�<�D�<&�<��<��<�ʮ<|��<W��<{c�<y;�<9�<��<b��<�|�<�G�<��<ހ<&Vy<K�p<��h<NG`<�W< �O<�yG<�A?<R7<`�.<�&<w<�A<(	<�<��;ט�;r�;��;�;���;�;�;��;GHo;��N;��.;��;�'�:o�:�@:�9Z�_�3�Ⱦ��@�Ӻ���r�%���C��`���}�7��]욻芨��ֵ���»ybϻ�ۻdv绳��H���k���	����ʜ�/a���!�X�%�_*��5.�&02�
6� �9��^=��@��:D��G�*�J�t�M�^�P�'�S���V��yY��M\�_���a�طd�X�g��Mj�!m�r�o�e�r��[u��x�a�z�a}�����F������A̓����K��P����Ȉ�
��cN�������/������ґ��&��Y{��Rϕ�"��s������m���X��:���9螼s.���t��˻�����*P��Ԟ����F�����������Y��o������t���ϲ�u(���}���϶�F���i��^���z���IC���  �  ��N=xYN=�M=	M=h^L=�K=)K=UJ=�I=��H=�DH=�G=��F=O9F=~�E==�D=]:D=��C=�B=�EB=��A=��@=$Q@=�?=T�>=�P>=��==��<=AA<=�;=9�:=h):=�v9=�8=�8=�c7=��6=C6=.X5=�4=M�3=gK3=��2=p�1=0.1=�s0=�/=��.=_,.=b-=�,=E�+=�*=U*=!8)=6X(=Ot'=�&=u�%=�$=
�#=C�"=¤!=� =�q=%G=�=B�=#}= =R�==@=_�=V1=͙=|�=N=�=P�
=	=�T=�=ۮ=G�=��<��<0�<G�<jS�<�U�<O�<�@�<�+�<.�<���<<��<��<y��<s�<�S�<%5�<��<W��<߲<I®<H��<>��<�a�<�;�<��<w�<N��<��<NS�<! �<G�<lwy<|q<��h<.k`<X<��O<��G</[?<2#7<��.<�&<�<�E<�<H�<��;x|�;���;c�;�ݸ;Cc�;Z��;��;�n;'_N;�<.;�Q;:�:�;�:DO?:�҅9��b���3��喺��Ӻ����%��PC���`�	N}�Wό�6���"N��G���]�»`#ϻA`ۻ�?绡��o���[���	�6������`��ڈ!�e�%��**��I.�fH2��%6���9�"=���@��\D�i�G���J�*�M���P�p�S��V�x�Y��U\��!_��a�&�d�_zg�Aj��m�+�o�n�r�P?u���w�V�z�'?}����;6��4|��W���� ���@��"�������}L�����㍼G3��[���Mۑ��1��և��uݕ��1��R����ҙ�����h�����t����9��~��.â��	��OS��ퟦ���C��Ț������WP��.����	���e����������l��ྶ�6��[�����𻼲9���  �  O=�[N=s�M=q	M=�]L=Y�K=iK=8QJ=?�I=��H=�=H=��G=��F=�0F=�E=��D=j2D=e�C=��B=,@B=�A==�@=�N@=��?=��>=nQ>='�==9�<=E<=ɓ;=�:=0:=O~9= �8=J8=Hl7=�6=�6=5_5=@�4=� 4=�O3=Ĝ2=��1=C/1=�s0=�/=��.=W).=�]-=�,=@�+=�*=�*=0)=�O(=l'=�&=�%=J�$=%�#=V�"=�!=č =�o=�F==��=�=�#=L�=MF={�=U9=��=�=�W=��=��
=�&	=�\=*�=�=B�=���<�<Z3�<-H�<BR�<LR�<XI�<�8�<�!�<��<���<���<ã�<7��<�a�<�B�<D%�<j	�<��<9Բ<x��<���<��<_�<�;�<��<��<ӽ�<֎�<X^�<1-�<'��<$�y<�:q<1�h<[�`<(@X<E�O<��G<,t?<�77<i�.<�&<s�<6I<�<k�<���;/^�;3��;�2�;H��;S#�;���;�T�;�n;��M;��-;x�;�G�:Df�:��=:&��9�|f��C4���^�Ӻ2��l�%�(!C��B`���|�ݞ��4}��Q���X���J»��λ%ۻ
绦�����tK��	���;���a��
�ב!�Q�%��;*�-_.�6a2�*B6��:�=�=��A��~D���G��J���M���P���S��V�E�Y��^\�@&_�}�a�b�d��rg��4j���l���o�nr��#u��w��{z��}�d��.&��4m��Ա����7��dy��������	K��Ŗ���卼 8��6���M䑼x<�������땼JA�������㙼�/���x�� ������E�� ���ˢ�����V��|����識6A��0������G��B���*���pW��K���S��	\��k���l����L������仼�0���  �  'O=�]N=��M=�	M=�\L=��K=��J=�MJ=��I=c�H=�7H=��G=��F=�(F=�|E=��D=�*D=t�C==�B=�:B=n�A=��@=L@=��?=<�>=�Q>=j�==~�<=GH<=�;=@�:=6:=�9=I�8=�#8=�s7=W�6=6=�e5=ݵ4==4=QS3=��2=;�1= 01=Us0=��/=��.=?&.=�Y-=�,=k�+=��*=�*=_()=�G(=d'=@|&=ɏ%=Ν$=n�#=��"=�!=� =%n=�E=M=*�=*�=M'=��=�K=��=�@=��=2
=K`=T�=��
=�.	=d=��=F�=��=��<��<�5�<�H�<�P�<�N�<�C�<�0�<��<��<4��<ö�<ۓ�<�q�<9Q�<�2�<B�<���<d�<�ɲ<�<喪<�z�<n\�<�:�<�<�<�Ñ<���<Rh�<9�<�	�<��y<�Zq<�i<��`</_X<P<��G<��?<lJ7<�/<Q�&<��<K<W<�<1��;^@�;���;�;�n�;��;pp�;��;��m;R>M;z'-;M;_�:���:-�<:�<�9�j��4�	F����Ӻ���,�%��B��	`���|��r��K���ۧ�X���»ìλ��ڻ���!h򻰝���=��	���2���c�O�"�!�p&��L*��s.�;y2�.]6�$:���=�B?A��D��G��K��N��Q�1�S���V�F�Y��g\�p+_���a���d�9lg�q*j�*�l�w�o��Wr�p
u�+�w�K^z��|��������_������!ꄼR.���r��B�������AJ��ߗ���荼=�����푼G���������/P��ţ�����?��=���p͝���Q�������Ң�}���Z��p����識N?��U����竼�?��k�����^J�����P����L��Z����M?��X����ڻ��(���  �  �O=�_N=9�M=h	M=�[L=��K=�J=JJ=`�I=q�H=�1H=K�G=1�F=�!F=�uE=�D=K$D=[~C=��B= 6B=m�A={�@=�I@=]�?=u�>=�Q>=T�==E�<=�J<=��;=��:=3;:=Ȋ9=u�8=R*8=oz7=��6=�6=�j5=��4=	4=[V3=��2=��1=x01=�r0=��/=��.=f#.=ZV-=��,=E�+=��*=2�)=�!)=A(==]'=�u&=|�%=�$=f�#=Q�"=��!=Z� =ll=�D=R=�=��=*=]�=NP=I�=�F=K�=c=�g=��=#�
=w5	=8j=ߗ=ž=:�=���<%�<�7�<�H�<�N�<�J�<#>�<�)�<��<���<]��<���<��<�c�<�B�<�$�<	�<��<�׶<{��<2��<ϐ�<�v�<�Y�<�9�<��<��<ȑ<��<�p�<C�<9�<C�y<�uq<Yi<�`<jyX<�,P<C�G<B�?<�Y7<�/<d�&<�<�K<r<j�<	��;�$�;>~�;���;�?�;���;�6�;�ӆ;�m;��L;5�,;��;��:9�:�I;:f~9Im���5��v��A�Ӻ���z%�
�B���_��t|��M��� ��O���yM���|λ��ڻm���D�~���e2�Wz	�������e���ޣ!�t&��[*�Ӆ.�e�2��t6�9:��=�k[A�B�D�s�G��!K�s-N��#Q�MT���V�-�Y�/p\��0_���a���d�egg�E"j�t�l�N�o��Er��t���w�Ez�0�|�!�����S��?���]ᄼ'��/m�����������I��9����덼�A��\�������tP��ԫ�����W]��|�������M������ڝ�w��&[�� ����٢�����^������
�>��[���J㫼99��[����篼K?�������볼�?�������㷼4�������һ��!���  �  X
O=�`N=��M=3	M=[L=F�K=��J=^GJ=�I=��H=~-H=p{G=�F=�F=wpE=��D=/D=�yC=v�B=62B=B�A=��@=�G@=
�?=��>=�Q>=�==��<=�L<=+�;=��:=	?:=�9=�8=8/8=T7=v�6=e6=o5=�4=4=�X3=5�2=k�1=�01=�r0=��/=��.=(!.=vS-=�,==�+=B�*=F�)=�)=�;(=�W'=tp&=��%=��$=t�#=�"=�!=I� =�j=+D=<=��=:�=�+=�=�S=T�=jK=Y�=�=Dm=S�=��
=x:	=�n=כ=�=��=���<��<�8�<KH�<M�<�G�<�9�<�#�<��<c��<��<���<_{�<tX�<�7�<�<���<5�<2϶<6��<��<��<s�<~W�<9�<I�<��<^ˑ<롍<�v�<�J�<��<E�y<�q<*3i<��`<*�X<�>P<��G<6�?<e7<�/<��&<��<�K<��<��<̹�;��;�b�;��;5�;?��;b
�;%��;X�l;�fL;V,;��;X��:�W�:_V::H6{9k�o�4�5�����Y�Ӻ����m%��B���_�dF|��1��� ��<���Aɴ�����Wλ��ڻl��=*�oj��*��t	�������g�����!��&��g*�6�.���2�Q�6�8M:�*�=�1qA��D��H��5K��?N�n4Q��T���V���Y�.w\�e5_���a�"�d�Edg�nj���l��o�8r��t��w�2z���|��l����`K��s����ڄ��!��2i��㱈������I��u���`qE��Y���(����W��S���6���g��������X������㝼a$��c��ߠ��7ߢ����a��a�����m=��P����߫�r4��D����௼�6��録��᳼�5��ˈ���ڷ��+��|��b̻����  �  lO=HaN=�M=	M=xZL=F�K=��J=�EJ=�I=�H=�*H=]xG=��F=/F=mE=N�D=�D=�vC=��B=�/B=8�A=C�@=[F@=!�?=@�>=�Q>=8�==H�<=�M<=��;=��:=fA:=Ǒ9=�8=>28=b�7=q�6=6"6=�q5=/�4=�4=�Y3=(�2=��1=�01=?r0=��/=��.=�.=�Q-=�,=��+=]�*=+�)=,)=_8(=�T'= m&=��%=ΐ$=��#=˛"=+�!=� =�i=�C==��=��=--=��=�U=��=DN=��=2=�p=Ž=�=�=	=�q=G�=�=j�=���<��<9�<�G�<�K�<�E�<�6�<8 �<e�<"��<!��< ��<tt�<pQ�<�0�<5�<o��<5�<�ɶ<���<O��<툪<�p�<V�<k8�<��<��<t͑<פ�<�z�<>O�<P#�<Y�y<��q<)@i<��`<��X<DJP<��G<��?<�k7<%/<U�&<$�<�K<��<�<���;� �;Q�;F��;2�;�m�;�;G��;|l;`*L;�,;$R;��:y��:P�9:�3y9|q�aI6�����&�Ӻ���te%���B��_�X)|� ��5왻�s�����y����@λ�ڻ/~���>]��)%�Yq	�������qi���ȯ!�+ &�ho*�^�.�f�2�*�6��Y:���=�)A��D�NH�mBK��KN��>Q��T���V�ǺY��{\�m8_�_�a��d�jbg��j���l�"�o��/r�/�t�؂w�6&z�i�|�e`������E�������ք�}���f��G�������J��j������H������#����\������;���m�������h_������ꝼ*��h��6����⢼�!���c��������<������ݫ��1������,ܯ��1��-����۳��/��ǂ���Է�t&���w���Ȼ����  �  :O=�UN=��M=	�L=SML=Q�K=!�J=:J=Y�I=��H="H=mpG=�F=�F=�cE=;�D=gD= fC=��B=B=�qA=��@=##@=�z?=��>=%>=Lx==�<=�<=|j;=g�:=�:=�U9=\�8=��7=�=7=��6=��5=L"5=�l4=R�3=�2=�C2=W�1=��0=^0=l?/=�u.=h�-=H�,=|,==*+=�N*=�o)=k�(=��'=m�&=�%=��$=Q�#=w�"=T�!=� =��=c�=}u=O?=��=$�=�V=��=�=%=O~=��=�Q=��=��=�G
=C�=��=��=_!=�F=���<j��<�%�<B�<HT�<�\�<b]�<@V�<%I�<q7�<p"�<��<���<n��<��<
��<���<.��<�y�<�h�<wW�<�D�<�0�<��<��<��<�ȕ<7��<}��<]d�<?@�<��<��y<ڤq< ]i<�a<��X<+�P<�QH<@<�7<(�/<rf'<�,<(�<��<v<.l�;���;ql�;n��;���;�"�;ԙ;��;��r;6�R;v33;ϩ;̹�:[��:l�Y:ɂ�9��ӸyX�]���@A���O���g��V8�<�T��q�Ym�����q�������\����ǻ=Ի�߻���h���v� ��'�cO�cQ��/�n��Ճ���"�5S'�+�+�4�/���3�0j7�[;��>��(B�A�E�b�H��K�d�N���Q�)�T��W���Z�@}]�oN`��c���e�7�h��qk��2n���p�8�s�^v��y�V�{�@b~�C����Ӂ��"���p����������[����������R������z��\�� �������p��˕�$���y���̙����g����������l:��j~��~¢����O�������䧼�3���9ث�7-��J����ٯ��0��s����ݳ�'3��#����ܷ�k0��
����׻��+���  �  � O=�UN=��M=�L=vML=��K=r�J=r:J=�I=7�H=�"H=4qG=��F=�F=�dE=�D=5D=�fC=b�B=�B=rA=�@=q#@=�z?=��>=(%>=;x==��<=v<=j;=�:=.:=
U9=��8=��7=�<7=ŉ6=�5=�!5=\l4=۵3=��2=�C2=:�1=��0=y0=�?/=v.=��-=��,=,=�*+=NO*=lp)=<�(=��'=W�&=��%=��$=�#=�"=��!=}� =�=��=�u=Z?=��=�=}V=@�=��=z=�}=!�=�P=��=��=G
=g�=4�=��=� =6F=��<���<\%�<�A�<YT�<Q]�<�]�<W�<DJ�<�8�<�#�<�<���<P��<���<ǲ�<-��<ƌ�<V{�<j�<oX�<�E�<~1�<�<)�<��<�ȕ<¨�<Ά�<|c�<'?�<M�<��y<��q<dYi<ka<��X<!�P<POH<�@<��7<}�/<je'<�+<�<��<�v</n�;Y��;�p�;i��;z��; )�; ۙ;ݣ�;@s;�	S;:B3;W�;���:���:��Y:�ž9s�Ҹ�A�B���w:���L��Lh��Y8���T�� q��p�����v�������b��g�ǻ�Ի��߻v�뻷����� ��(��O�KQ� /�������T�"�lQ'���+�~�/���3��f7�;�'�>��$B��}E�1�H�n�K���N�2�Q�V�T���W�v�Z��|]��M`��c�M�e�'�h�sk�t4n�(�p���s��`v�}y�Խ{��e~������ԁ��#���q������]���[��竉������Q��>���� ��][��"���Y��Po���ɕ��"��.x���ʙ����qe�����r���"9��C}������7���N��X����䧼�3��3����ث��-��<���ۯ� 2��눲�/߳��4��ĉ��	޷��1��,����ػ��,���  �   O=#UN==�M=2�L=�ML=?�K=|�J=�;J=z�I=�H=�$H=zsG=+�F=TF=gE=��D=�D=iC=a�B=mB=�sA=T�@=l$@=Z{?=��>=(%>=�w==J�<=�<=�h;=S�:=^:=S9=z�8=��7=�:7=��6=��5=�5=�j4=u�3=��2=�B2=��1=��0=�0=@/=�v.=ש-=�,=�,=�,+=lQ*=�r)=��(=�'=��&=A�%=��$=#�#=��"=�!=�� =�=V�=�u=c?=6�=D�=~U=��=�~==U{=��=%N=	�=��=}D
=�=��=��==�D= ��<o��<�$�<�A�<�T�<�^�<�_�<�Y�<vM�<f<�<.(�<��<���<Z��<��<׷�<��<A��<W�<�m�<n[�<OH�<]3�<<�<��<��<ȕ<@��<���<�`�<�;�<I�<��y<@�q<�Oi<�	a<6�X<^�P<XGH<�@<c�7<�/<Db'<�)<��<��<�x<�u�;?��;.}�;0�;���;R<�;��;I��;�7s;�5S;;m3;Y�;��:��:�kZ:o��9}и� ����e/��_M���m��c8�p�T��5q��}��#������⡮��s����ǻ1*Ի�
���������� �G+�>Q��Q��-�o�����"��K'�؀+�ɕ/��3��]7�#;�)�>��B�tE�ĲH���K�
�N�c�Q���T�,�W���Z�pz]�M`�c��e��h�'wk��9n���p�A�s�Niv�>y���{��n~�	���ف��'��u���D��H]����������@Q����� ����X��0������`k���ŕ����Gs���ř�����`������C�v5��z�������M��~���䧼/4��I���yګ�C0��+����ޯ�
6��*����㳼h9��4���Mⷼ�5�������ۻ�/���  �  ��N=9TN=بM=A�L=jNL=C�K=��J=�=J=�I=��H=!(H=wG=��F=NF=%kE=��D=_D=lC=��B=2B=�uA==�@=�%@=D|?=j�>=%>=`w==D�<=�<=�f;=ִ:=x:=�O9=�8=�7=77=�6=��5=�5=h4=3�3=��2=�A2=�1=��0=�0=�@/=�w.={�-=:�,=A,=�/+=�T*=Sv)=}�(=�'=��&=�%=��$=h�#=��"=��!=�� =��=D�=ov=Z?=��=:�=�S=��=,|=b�=�w=��=�I=Ǥ=��=L@
=�=m�=��=a=�B=���<G��<k#�<�A�<�U�<�`�<�b�<�]�<tR�<cB�<�.�<1�<w�<���<8��<ؿ�<���<M��<���<s�<`�<�K�<�5�<��<U�<>�<�ƕ<���<�<�[�<6�<��<��y<ňq<9@i<�`<+�X<�wP<�:H<� @<;�7<�/<\]'<H'<��<�<c|<���;�;���;��;���;]Z�;u�;�ۉ;s;�{S;Q�3;6!;��:!^�:U%[:��9�J̸ǣ�<s��� ��N���v��u8��U��Wq�����*:������4����3ȻTCԻ�!��뻮���#� ��/��S�R��,�(��z���"��B'�_v+�l�/�<|3��N7�Y;���>��
B�@dE��H��K���N���Q���T�9�W�3�Z�[w]��K`��c���e��h�~k��Bn�Eq�I�s��vv��(y�v�{�C}~�6����߁�k-��)z��Mƅ�}��s_��ǭ��
���~P��N���k���CU������m
��e������B��bk����������X��Z����鞼�/�� u�������J��C���E䧼�4������1ݫ�4������䯼C<������과�@������:鷼<��O���y໼�2���  �  ��N=�RN=/�M=?�L=OL=��K=��J=B@J=��I=��H=R,H=�{G=��F=cF=HpE=��D=>D=qC=��B=� B=�xA=��@=�'@=q}?=��>=�$>=�v==��<=�<=d;=��:=��9=�K9=Y�8=?�7=B27=;6=$�5=�5=sd4=;�3=��2=�?2=�1=�0=0=�A/=uy.=��-=��,=�
,=�3+=
Y*=�z)=c�(=�'=��&=��%=(�$=��#=��"=�!=V� =k�=��=w=<?=��=��=�Q=��=�x=D�=s=��=�D=8�=(�=�:
=�|=��=��=�=�?=H��<,��<�!�<yA�<W�<c�<�f�<�b�<�X�<J�<�7�<�"�<��<��<���<��<T��<X��<���<z�<�e�<sP�<X9�<��<��<|�<aĕ</��<|�<�U�<�.�<6�<��y<�tq<�+i<��`<��X<�dP<*H<�?<?�7<��/<�V'<B#<��<��<�< ��;��;ש�;8=�;(ٺ;���;�:�;��;J�s;g�S;�4;t;�/�:��:�\:�Y�9t\Ǹ�,�N��u���T�������8�c=U���q�����}Y�������஻
���i5Ȼ�dԻ�@ໄ�������� ��5�nW�FS�7+����s���"�v7'��h+��y/��j3��;7�B�:�C�>��A�,PE���H�l�K���N�|�Q���T��W�חZ��s]��J`�Jc���e���h�/�k�LNn�/q�}�s��v�i;y���{�u�~�i���>聼N5��ۀ���˅�����b������|����O����� ����P��©��}�� ]���������Ya��S�������N�����)ូ&(���n��ĵ�����:H��͔��#䧼	6�������ૼ9�����z민�D������l���bJ�����E�zD��ҕ���滼8���  �  N�N=LQN=P�M=*�L=�OL=�K=��J=CJ=��I=��H=1H=�G=��F=N#F=:vE=q�D=�D=/vC=E�B=�$B=?|A=<�@=�)@=�~?=]�>=�$>=�u==	�<=_<=�`;=��:=�9=fF9=�8=��7=�,7=�y6=��5=�5=4`4=��3=��2=�=2=��1=x�0=40=hB/=
{.=ݯ-=��,=D,=�7+=�]*=X�)=�(=�'=��&=��%=v�$=k�#=��"=��!=)� =|�=ڤ=zw=�>=��=ݪ=O=��=rt=Y�=�m=��=5>=��=��=�4
=�v==�=��=�=`<=���<p��<��<�@�<�W�<�e�<�j�<�h�<9`�<�R�<�A�<�-�<K�<�<���<���<���<���<ؖ�<��<cl�<�U�<�<�<�!�<��<]�<���<͜�<!v�<N�<�%�<��<��y<P]q<ki<��`<5�X<2OP<{H<7�?<��7<R~/<nN'<A<�<�<]�<'��;2�;���;�_�;�;}��;uk�;R;�;�At;�=T;�m4;��;��: ��:�]:E�9~������'������`��8����8��hU���q�4Ά��~���须5�� ޻�A_Ȼ��Ի�d�u�����?� ��=�\��T��)�a���l��"��*'�EY+�h/��V3��%7���:�Ph>��A��8E��zH�Z�K�6�N���Q� �T�ثW���Z��o]��I`�O c���e���h�1�k�i\n��!q�Y�s�!�v�{Qy���{�'�~�\�����~>�������҅���6f��̱��%����N�����=����K��(��������S��p������U��q��������C��e����מ�����g���������kE������$䧼�7�������嫼?������2���sN�����������U��I������kN������u>>���  �  ��N=nON=2�M=��L=/PL=-�K=�J=�EJ=4�I=�H=!6H=x�G=��F=�)F=�|E=��D=�%D=�{C=1�B=�(B=�A=��@=n+@=�?=��>=5$>=?t==��<=u<=,];=3�:=�9=�@9=�8=o�7=T&7=�s6=�5=�5=�[4=��3=r�2=N;2=�1=��0=-0=-C/=�|.=2�-=��,=,=i<+=c*=�)=	�(=�'=��&=��%=�$=��#=1�"=W�!=� =��=�=�w=�>=��=��=L=��=�o=��=�g=�=I7=��=��=�-
=jp=F�=U�==�8=��<*��<�<@�<�X�<Wh�< o�<�n�<�g�<�[�<"L�<@9�<�$�<��<���<Y��<K̾<}��<s��<D��<s�<�Z�<M@�<�#�<��<��<}��<���<qo�<�E�<��<��<�y<�Cq<�h<��`<�rX<�7P<H<X�?<�7<sq/<-E'<4<��<�<͉<$��;�H�;���;!��;�+�;�ݪ;���;|q�;S�t;׫T; �4;�6;Փ�:�!�:R3^:���9�M��L7�6�������r�����i�8�^�U���q�򆻏���Z��`9������ȻR�ԻI�໕
�l3��I��F��a��W�R)�����e��"��'�VI+�1U/�'A3��7�w�:�O>���A�C E��cH��K�[�N��Q��T��W�Q�Z�sl]�yI`�n#c��e�!�h�؞k��kn�B4q���s��v��iy�Q|�ѿ~�V��������H��ّ���م�"���j������Y ��XN�����]F��]���K�9J����������OI��ߚ��>ꚼ�7��0���H͞����`��&���T����B��C����䧼�9������꫼�E��ա������+Y��m������Eb���������@Y��Y�������'E���  �  ��N=^MN=�M=\�L=�PL=V�K=��J=�HJ=��I=V�H=;H=�G=j�F=�/F=��E=��D=�+D=��C=��B=-B=�A=��@=)-@=��?=��>=�#>=�r==��<=x<=hY;=��:=��9=;;9=��8=1�7= 7=zm6=J�5=(	5=�V4=��3=�2=�82=�1=��0=�0=�C/=�}.=a�-= �,=�,=�@+=h*=~�)=�(= �'=��&=l�%=��$=w $=��"=��!=�� =��=.�=3x=�==�=u�=�H=��=k=w�=ma=��=J0=_�=Y�=�&
=�i=�=��=[=�4=���<���<�<�>�<vY�<�j�<;s�<�t�<Ao�<�d�<eV�<�D�<�0�<z�<L�<���<�׾< ��<˩�< ��<�y�<o_�<sC�<F%�<a�<���<ۺ�<s��<sh�<1=�<��<��<�yy<�)q<n�h<��`<SYX<sP<��G<�?<7<Zd/<9;'<�<6�<q�<��<½�;_�;r�;���;/U�;��;�њ;ئ�;�u;AU;V@5;И;4F�:��:9?_:`��9�4��Y���儺����\�������8���U��9r����є�C��Uh��t<����ȻJ�Իi���.�#R����P�h�[��)�[���_���"�I'�:+��B/��,3���6�4�:�#6>�ثA� E��LH�E|K�
�N���Q�}�T���W�b�Z�ri]��I`�'c�� f�	�h��k��{n�)Gq�mt���v��y�n1|���~�i���	��S�������ᅼ+(��.o���������:N�����GZA��Е��M뒼�@��
���Oꖼ.=��x����ݚ��+��,x��hÞ�,���X��g���L�-@��]���\姼<�����L��L��S������+d��*���*���n���¶����Vd��k�������[L���  �  �N=HKN=��M=��L=�PL=?�K=��J=KJ=֜I=5�H=t?H=�G=��F=E5F=s�E=H�D=�0D=܅C=F�B=�0B=�A=��@=�.@=n�?=��>=�">=]q==��<=�
<=�U;=x�:=�9=�59=9�8=D�7=7=�g6=õ5=5=8R4=��3=��2=<62=B~1=��0=�0=*D/=.=?�-=��,=%,=�D+=�l*=��)=W�(=��'=X�&=��%=��$=�$=o#=�!=M� =/�=�=@x====��=(�=�E=��=�f=N�=�[==�=�)=��=��= 
=�c=a�=��=�=�0=���<��<E�<}=�<�Y�<il�<�v�<�y�<v�<m�<�_�<AO�<<�<!'�<��<���<��<�ʺ<Q��<9��<*�<�c�<F�<:&�<��<�ޙ<��<F��<�a�<�4�<!�<�ۀ<4by<�q<D�h<�`<AX<�P<D�G<��?<�~7<�W/<Q1'<=<��<�<̐<W��;�r�;`�;��;�z�;�7�;| �;�׊;��u;�{U;ߠ5;L�;���:�N�:t.`:��9�²�Zf��Є��������v��h9���U��ur��:�������m������i��8�Ȼ]ջ��8Q��o���MY��n�Q^�>*�I���Z���"�C'�,+�62/��3���6��:�4>�ޔA���D��7H�kiK�X�N���Q���T���W�`Z��g]��J`��*c��f���h���k�f�n��Xq�� t���v�W�y�/I|���~��ǀ�����\������%酼'.���s������X��uN��͛��{뎼=�����䒼N8��m����ߖ�2������Қ�� ��n��b���F��yR��f�����.>������T槼\>����������S��q�������n��^ʲ��#���z���ζ�����n��ջ�����jS���  �  ��N=kIN=h�M=4�L=�PL=�K=��J=MJ=q�I=e�H==CH=-�G=^�F=:F=D�E= �D=R5D=�C=��B=�3B=~�A=��@=�/@=��?=��>=">=�o==��<=�<=�R;=��:=��9=519=E|8=&�7=�7=�b6=�5=��4=6N4=-�3=��2=�32=�|1={�0=.0=gD/=�.=ɷ-=��,=�,=5H+=�p*=�)=�(=l�'=�&=M�%=�%=�$=�#=��!=L� =��=��=:x=�<=8�=�=-C=��=�b=��=�V=��=�#=�}=��=h
=&^=Y�=6�=�=}-=I��<���<�<'<�<�Y�<�m�<�y�<�}�<�{�<�s�<�g�<X�<uE�<�0�<��<z�<��<�Һ<T��<��<̓�<�f�<H�<�&�<,�<�ܙ<���<���<�[�<�-�<���<rҀ<�My<��p<��h<%j`<�+X<��O<�G<��?<q7<`L/<�('<<��<��<#�<���;���;1�;���;C��;\�;�'�;��;��u;�U;��5;�>;.r�:�Ů:v�`:�N�9��!�:�������V������
A9�,V��r�BZ�����!���ɻ������eɻ-3ջ�໶o�����'��a��t�
b�O+����TV���"�'�&�x +�f$/��	3�8�6�c|:��>�w�A�&�D�/&H�7YK�yzN��Q���T� �W�M{Z�2f]�9L`��.c�6f���h���k��n��hq�2t��v�P�y��]|���р�M��xe��>�����3���w������	���N��ؚ��,鎼r9��I���ޒ�#1��-����֖��(��by��ɚ����te���������� M��M����꣼�<������h秼�@������p����Y������3���w��#Բ�.������ض��)��x��)ĺ�	���Y���  �  ��N=�GN=i�M=��L=�PL=^�K=��J=�NJ=k�I=��H=FH=U�G=��F=�=F=�E=��D=�8D= �C=��B=*6B=\�A=��@=�0@=J�?=��>=t!>=�n==�<=�<=
P;=��:={�9=�-9=hx8='�7=�7=�^6=2�5=.�4=K4=}�3=��2=22=M{1=��0=�0=�D/=��.=�-=d�,=,=�J+=�s*=�)=m�(=	�'=��&=��%=�%=�$=#	#=��!=�� =~�=!�=x=�;=�=��=A=��=�_=/�=�R=��=�=3y=0�=�
=�Y=z�=��=��=�*=!��<���<R�<;�<�Y�<�n�<�{�<��<��<y�<�m�<�^�<�L�<d8�<I"�<�
�<3�<�غ<���<���<3��<Ci�<aI�<?'�<�<ۙ<��<���<�V�<(�<��<-ˀ<�=y<��p<V�h<AY`<�X<��O<�G<�?<pf7<gC/<�!'<J <��<��<��<D��;n��;�A�;���;n��;]w�;F�;�!�;�v;�V;�/6;�w;��:��:�a:�5�9�x������������������]9�	OV���r��r��j6��X���2گ������,ɻ�OջZử��n���y0��h�qy��d�R,�����S�2�"�L�&��+��/���2���6��m:���=��rA���D��H�0MK�pN�T�Q���T�c�W��xZ��e]�hM`��1c�
f���h���k�e�n�uq��?t��w�	�y��m|���ـ��$��)l��?������7��*{��ӿ��k��/O��V����玼�6������sْ��+��~��Ж�[!��
r���������_��򬞼����I��J��� 飼�;������U觼�B��f���R���|^��.�������~���۲��5��!����඼f1�����ʺ����Z^���  �  E�N=�FN=��M=L�L=�PL=��K=��J=jOJ=��I=X�H=�GH=S�G=��F=�?F=.�E=��D=�:D=�C=d�B=�7B=z�A=��@=51@=��?=w�>=!>=n==޹<=�<=kN;=�:=`�9=O+9=�u8=��7=m7=:\6=ժ5=��4=I4=��3=1�2=�02=_z1=
�0=�0=�D/=�.=��-=X�,=N,=UL+=Tu*=$�)=��(=8�'=��&=��%=	%=x$=�
#= "=�� =�=h�=x=|;=Z�=e�=�?=6�=�]=��=;P=�=�=hv=e�=7
=ZW=
�=��=��=8)=g��<���<��<L:�<�Y�<�o�<
}�<���<���<j|�<�q�<�b�<HQ�<�<�<�&�<>�<i��<�ܺ<���<9��<9��<�j�<9J�<Y'�<��<�ٙ< ��<<��<�S�<X$�<��<�ƀ<�3y<��p<ϓh<�N`<[X<��O<�G<G�?<�_7<�=/<f'<�<��<��<��<��;ڕ�;�K�;��;�»;���;�X�;T5�;q@v;�8V;�U6;}�;h�:W�:w�a:��9�⪸��������������'��o9�nfV�'�r������G���¢�!��¼�r?ɻ	bջN)Ử������6�m��|�g�<-�t���Q�B�"�D�&�R+�V/��2���6�e:���=��iA���D��H��EK�fiN��}Q���T�{�W��vZ�
e]�eN`��3c��f�,�h�s�k�;�n��|q�xHt�7w���y��w|����ހ�4)��lp�� �������:��_}��w���_���O��񙍼�掼Q5��~����֒�[(��4z���˖�����m��M���i��[��V��������F��w����磼;������
駼�C��e���� ���a���®��#��#����಼�:������嶼86�������κ�X��va���  �  ��N=�FN=��M=+�L=�PL=��K=��J=�OJ=�I=��H=jHH= �G=��F=�@F=�E=��D=�;D=��C=��B=8B=܋A=�@=U1@=��?=_�>=� >=�m==��<=<=�M;=A�:=��9=�*9=$u8=��7=7=_[6=�5=3�4=nH4=�3=��2=�02=z1=��0=i0=�D/=	�.=Ź-=��,=�,=�L+=�u*=Ԛ)=F�(=�'=��&=��%=�	%=$=5#=q "=� =C�=u�=x=P;=�=�=:?=��=�\=:�=`O=	�=�=du=c�=O
=}V=8�=��=:�=�(=���<%��<��<:�<�Y�<�o�<�}�<���<s��<�}�<�r�<|d�<�R�<�>�<�(�<��<���<�ݺ<�¶<��<߉�<k�<RJ�<5'�<��<_ٙ<s��<q��<�R�<�"�<e�<�Ā<�0y<��p<�h<�J`<�X<��O<�G<��?<Z]7<8</<'<J�<��<R�<��<���;���;XO�;��;�ǻ;���;>_�;�<�;�Ov;�FV;�b6;S�;�-�:Ph�:Lb:M��9Ǉ��C��~���7�������� v9��oV�o�r�]���N���ɢ�p���ʼ�<Fɻdhջr/���ʰ���7�]n�~��g��-�w��wQ�[�"���&��+�1/���2�Ӹ6�b:���=�)fA���D��H�/CK�8gN�|Q�0�T���W��vZ�
e]��N`��4c��f���h�Q�k���n�nq��Kt�gw�-�y�}{|��"�)����*���q��R���6���`;��~�������O��虍�p掼�4�������Ւ�@'���x��dʖ�l���k�������
���Y��2��������E��ӕ��f磼�:��֐��H駼^D���������b��Į�%������Ⲽ�<�������綼�7��(���-к�����b���  �  E�N=�FN=��M=L�L=�PL=��K=��J=jOJ=��I=X�H=�GH=S�G=��F=�?F=.�E=��D=�:D=�C=d�B=�7B=z�A=��@=51@=��?=w�>=!>=n==޹<=�<=kN;=�:=`�9=O+9=�u8=��7=m7=:\6=ժ5=��4=I4=��3=1�2=�02=_z1=
�0=�0=�D/=�.=��-=X�,=N,=UL+=Tu*=$�)=��(=8�'=��&=��%=	%=x$=�
#= "=�� =�=j�=x=;=]�=j�=�?==�=�]=�=FP=��=�=yv=y�=M
=rW=$�=��= �=V)=���<��<,�<�:�<�Y�<�o�<?}�</��<���<�|�<�q�<c�<SQ�<�<�<�&�<0�<S��<�ܺ<���<��<
��<�j�<J�<"'�<��<�ٙ<쮕<��<�S�<2$�<��<gƀ<�3y<��p<ϓh<�N`<|X<	�O<U�G<��?<�_7<)>/<�'<��<n�<��<$�<���;���;TL�;3�;Eû;��;Y�;n5�;^@v;�8V;U6;��;$�:ST�:1�a:��9C�����ϸ�����@���L�r9�vhV��r�w����H���â���Gü�@ɻ�bջ�)������)6�+m��|�,g�O-�����Q�M�"�L�&�Y+�\/�"�2���6�
e:���=��iA���D��H��EK�giN��}Q���T�|�W��vZ�
e]�fN`��3c��f�,�h�s�k�;�n��|q�xHt�7w���y��w|����ހ�4)��lp�� �������:��_}��w���_���O��񙍼�掼Q5��~����֒�[(��4z���˖�����m��M���i��[��V��������F��w����磼;������
駼�C��e���� ���a���®��#��#����಼�:������嶼86�������κ�X��va���  �  ��N=�GN=i�M=��L=�PL=^�K=��J=�NJ=k�I=��H=FH=U�G=��F=�=F=�E=��D=�8D= �C=��B=*6B=\�A=��@=�0@=J�?=��>=t!>=�n==�<=�<=
P;=��:={�9=�-9=hx8='�7=�7=�^6=2�5=.�4=K4=}�3=��2=22=M{1=��0=�0=�D/=��.=�-=d�,=,=�J+=�s*=�)=m�(=	�'=��&=��%=�%=�$=%	#=��!=�� =��=%�="x=�;=!�=��=A=��=�_=B�=�R=��=�=Uy=W�=$
=+Z=��=��= =+=���<^��<��<�;�<Z�<Oo�<|�<g��<)��<by�<n�<�^�<�L�<j8�<>"�<�
�<�<�غ<^��<<��<ن�<�h�<�H�<�&�<�<�ڙ<���<\��<|V�<�'�<���<�ʀ<�=y<��p<U�h<`Y`<�X<��O<m�G<��?<g7<%D/<�"'<<��<Ѻ<e�<���;��;�B�;���;\��;x�;�F�;�!�;�v;�V;Q.6;/v;���:_�:�a:��9��Q��3�����������a9��RV���r��t��8��߱���ۯ�Ѱ���-ɻ�Pջ;�r������0��h��y�'e�v,����S�F�"�]�&��+�/���2��6��m:���=��rA���D��H�2MK�
pN�U�Q���T�d�W��xZ��e]�hM`��1c�
f���h���k�e�n�uq��?t��w�
�y��m|���ـ��$��)l��?������7��*{��ӿ��k��/O��V����玼�6������sْ��+��~��Ж�[!��
r���������_��򬞼����I��J��� 飼�;������U觼�B��f���R���|^��.�������~���۲��5��!����඼f1�����ʺ����Z^���  �  ��N=kIN=h�M=4�L=�PL=�K=��J=MJ=q�I=e�H==CH=-�G=^�F=:F=D�E= �D=R5D=�C=��B=�3B=~�A=��@=�/@=��?=��>=">=�o==��<=�<=�R;=��:=��9=519=E|8=&�7=�7=�b6=�5=��4=6N4=-�3=��2=�32=�|1={�0=-0=gD/=�.=ɷ-=��,=�,=5H+=�p*=�)=�(=l�'=�&=N�%=�%=�$=�#=��!=O� =��=��=@x=�<=B�=�==C=��=�b=��=�V=��=%$=�}=��=�
=h^=��=��=*=�-=���<���<,�<�<�<cZ�<�n�<6z�<Q~�<|�<Rt�<$h�<IX�<�E�<�0�<��<T�<H�<vҺ<�<���<M��<[f�<�G�<Q&�<��<*ܙ<)��<��<[�<O-�<V��</Ҁ<qMy<l�p<��h<Qj`<X,X<S�O<��G<x�?<r7<kM/<�)'<9<��<��<P�<��;���;�2�;���;���;]�;�(�;��;��u;�U;,�5;z<;�k�:��:S�`:c(�9����2��̄����#���|���F9��1V�Z�r��\�����I���½��]����ɻ�4ջF���p�����:(�b�u�Hb��+����wV��"�?�&�� +�u$/��	3�C�6�k|:��>�|�A�*�D�2&H�:YK�{zN��Q���T�!�W�M{Z�2f]�:L`��.c�7f���h���k��n��hq�2t��v�P�y��]|���р�M��xe��>�����3���w������	���N��ؚ��,鎼r9��I���ޒ�#1��-����֖��(��by��ɚ����te���������� M��M����꣼�<������h秼�@������p����Y������3���w��#Բ�.������ض��)��x��)ĺ�	���Y���  �  �N=HKN=��M=��L=�PL=?�K=��J=KJ=֜I=5�H=t?H=�G=��F=E5F=s�E=H�D=�0D=܅C=F�B=�0B=�A=��@=�.@=n�?=��>=�">=]q==��<=�
<=�U;=x�:=�9=�59=9�8=D�7=7=�g6=õ5=5=8R4=��3=��2=<62=B~1=��0=�0=)D/=.=?�-=��,=%,=�D+=�l*=��)=W�(=��'=X�&=��%=��$=�$=q#=!�!=Q� =3�=�=Gx=F==��=8�=�E= �=�f=o�=�[=j�=�)=Ճ=��=` 
=�c=��=�=*=81=w��<���<�<M>�<xZ�<'m�<tw�<6z�<�v�<�m�<#`�<�O�<(<�<*'�<��<���<;�<6ʺ<ر�<���<�~�<�b�<YE�<�%�<(�<*ޙ<n��<���<a�<w4�<��<�ۀ<�ay<�q<B�h<�`<�AX<R	P<�G<��?<�7<�X/<�2'<�<_�<��<<�<��;u�;��;��;�|�;�8�;G�;P؊;~�u;�zU;̞5;W�;B��:�E�:v`:���9����E���ބ�J��^������o%9�wV�||r��=�������p��z����k��-�Ȼջ��ໍR�#q�����Y�o��^�~*�~���Z���"�`'�,+�I2/��3���6��:�<>��A���D��7H�niK�Z�N���Q���T���W�aZ��g]��J`��*c��f���h���k�f�n��Xq�� t���v�W�y�/I|���~��ǀ�����\������%酼'.���s������X��uN��͛��{뎼=�����䒼N8��m����ߖ�2������Қ�� ��n��b���F��yR��f�����.>������T槼\>����������S��q�������n��^ʲ��#���z���ζ�����n��ջ�����jS���  �  ��N=^MN=�M=\�L=�PL=V�K=��J=�HJ=��I=V�H=;H=�G=j�F=�/F=��E=��D=�+D=��C=��B=-B=�A=��@=)-@=��?=��>=�#>=�r==��<=x<=hY;=��:=��9=;;9=��8=1�7= 7=zm6=J�5=(	5=�V4=��3=�2=�82=�1=��0=�0=�C/=�}.=a�-=��,=�,=�@+=h*=~�)=�(= �'=��&=m�%=��$=x $=��"=��!=�� =��=4�=<x=>=�=��= I=��=<k=��=�a=��=�0=��=��='
=-j=��=C�=�=5=���<���<��<�?�<VZ�<ek�< t�<3u�<�o�<ne�<�V�<E�<1�<��<7�<}��<�׾<���<D��<���<�x�<�^�<�B�<y$�<��<��<��<���<�g�<�<�</�<B�<yy<a)q<l�h<8�`<�YX<( P<��G<$�?<�7<�e/<�<'<D<��<�<Y�<���;�a�;��;ϩ�;�V�;��;�Қ;:��;gu;�U;>5;��;�=�:�:�'_:7X�9���_��f������z�����f 9�>�U��@r���EԔ�F��k���>���Ȼ:�Ի��w0�kS��]��P�}h�V[��)�����_���"�j'�:+��B/��,3���6�?�:�,6>�߫A�E��LH�I|K��N���Q��T���W�c�Z�si]��I`�'c�� f�	�h��k��{n�*Gq�mt���v��y�n1|���~�i���	��S�������ᅼ+(��.o���������:N�����GZA��Е��M뒼�@��
���Oꖼ.=��x����ݚ��+��,x��hÞ�,���X��g���L�-@��]���\姼<�����L��L��S������+d��*���*���n���¶����Vd��k�������[L���  �  ��N=nON=2�M=��L=/PL=-�K=�J=�EJ=4�I=�H=!6H=x�G=��F=�)F=�|E=��D=�%D=�{C=1�B=�(B=�A=��@=n+@=�?=��>=5$>=?t==��<=u<=,];=3�:=�9=�@9=�8=o�7=T&7=�s6=�5=�5=�[4=��3=r�2=N;2=�1=��0=-0=-C/=�|.=2�-=��,=,=i<+=c*=�)=	�(=�'=��&=��%=�$=��#=3�"=Z�!=� =��="�=�w=�>=��=Ө=!L=��=�o= �=�g=P�=�7=ё=��=�-
=�p=��=��=�=�8=���<��<��<A�<�Y�<3i�<�o�<no�<zh�<\�<�L�<�9�<�$�<��<���<#��<�˾<��<矶<���<Qr�<�Y�<~?�<�"�<��<��<���<���<�n�<3E�<R�<��<��y<gCq<�h<ĳ`<FsX<I8P<H<��?<t�7<�r/<�F'<�<5�<��<w�<O��;�K�;_��;h��;�-�;`ߪ;��;�q�;�t;�T;��4;�3;��:,�:^:ڞ�9H8��aV�d�� ��|��������8�8�U�|r�����ݪ��g��+<��m��Y�ȻS�Ի����4����+G�b�X��)�����e�7�"�'�rI+�GU/�9A3��7���:�O>���A�I E��cH��K�^�N�
�Q��T�	�W�R�Z�tl]�zI`�o#c��e�"�h�؞k��kn�B4q���s��v��iy�Q|�ѿ~�V��������H��ّ���م�"���j������Y ��XN�����]F��]���K�9J����������OI��ߚ��>ꚼ�7��0���H͞����`��&���T����B��C����䧼�9������꫼�E��ա������+Y��m������Eb���������@Y��Y�������'E���  �  N�N=LQN=P�M=*�L=�OL=�K=��J=CJ=��I=��H=1H=�G=��F=N#F=:vE=q�D=�D=/vC=E�B=�$B=?|A=<�@=�)@=�~?=]�>=�$>=�u==	�<=_<=�`;=��:=�9=fF9=�8=��7=�,7=�y6=��5=�5=4`4=��3=��2=�=2=��1=x�0=40=hB/=
{.=ݯ-=��,=D,=�7+=�]*=X�)=�(=�'=��&=��%=v�$=l�#=��"=��!=-� =��=�=�w=
?=��=�=#O=��=�t=~�=�m=��=o>=�=��=�4
=Kw=��=�==�<=��<^��<� �<�A�<�X�<�f�<�k�<ci�<�`�<<S�<�A�<.�<u�<#�<���<���<3��<%��<Q��<w��<�k�<�T�<<�<!�<��<��<���<��<}u�<�M�<"%�<���<�y<]q<ii<��`<��X<�OP<gH<U�?<=�7<�/<�O'<�<��<��<��<6��;�4�;z��;�a�;��;ٯ�;Wl�;�;�;wAt;�<T;4k4;8�;���:�u�:�]:��9ڹ¸��k7��~���p��8����8�rpU���q��ц�����졻����໻paȻ��Իlf�������� �*>��\�RU�:*�����l�-�"��*'�_Y+�h/��V3��%7� �:�Xh>��A��8E��zH�^�K�8�N���Q��T�٫W���Z� p]��I`�O c���e���h�2�k�j\n��!q�Z�s�!�v�{Qy���{�'�~�\�����~>�������҅���6f��̱��%����N�����=����K��(��������S��p������U��q��������C��e����מ�����g���������kE������$䧼�7�������嫼?������2���sN�����������U��I������kN������u>>���  �  ��N=�RN=/�M=?�L=OL=��K=��J=B@J=��I=��H=R,H=�{G=��F=cF=HpE=��D=>D=qC=��B=� B=�xA=��@=�'@=q}?=��>=�$>=�v==��<=�<=d;=��:=��9=�K9=Y�8=?�7=B27=;6=$�5=�5=sd4=;�3=��2=�?2=�1=�0=0=�A/=uy.=��-=��,=�
,=�3+=
Y*=�z)=c�(=�'=��&=��%=)�$=��#=��"=�!=Y� =p�=��=w=F?=��=ì=�Q=�=�x=e�=;s=��=�D=s�=k�=7;
=O}=�=��=>=6@=��<��<�"�<JB�<�W�<�c�<^g�<tc�<gY�<�J�<�7�<#�<��<��<���<���<��<���<E��<�y�<Pe�<�O�<�8�<>�<>�<��<�Õ<���<|{�<,U�<.�<��<q�y<�tq<�+i<��`<��X<�eP<�*H<�?<f�7<��/<�W'<�$<-�<+�<T�<���;m�;!��;1?�;�ں;΂�;�;�;:�;�s;=�S;�4;q;(�:|ܫ:��[:�*�9j'ȸ�G� \�����Xc��)����8�0DU�t�q�����Z\��/ġ�K㮻:���^7Ȼ`fԻ1B��������E� �j6��W��S�v+�R���s��"��7'��h+��y/��j3��;7�K�:�J�>��A�1PE�ĐH�o�K���N�~�Q���T���W�ؗZ��s]��J`�Kc���e���h�0�k�MNn�/q�~�s��v�i;y���{�u�~�i���>聼N5��ۀ���˅�����b������|����O����� ����P��©��}�� ]���������Ya��S�������N�����)ូ&(���n��ĵ�����:H��͔��#䧼	6�������ૼ9�����z민�D������l���bJ�����E�zD��ҕ���滼8���  �  ��N=9TN=بM=A�L=jNL=C�K=��J=�=J=�I=��H=!(H=wG=��F=NF=%kE=��D=_D=lC=��B=2B=�uA==�@=�%@=D|?=j�>=%>=`w==D�<=�<=�f;=ִ:=x:=�O9=�8=�7=77=�6=��5=�5=h4=3�3=��2=�A2=�1=��0=�0=�@/=�w.={�-=:�,=A,=�/+=�T*=Sv)=}�(=�'=��&=�%=��$=i�#=��"=��!=�� =��=I�=uv=b?=��=G�=�S=��=C|=}�=�w=��=J=��=��=�@
=Z�=��=�=�=C=e��<���<$�<lB�<�V�<!a�<kc�<1^�<�R�<�B�<+/�<f�<��<���<)��<���<P��<���<L��<�r�<�_�<XK�<j5�<Y�<��<��<ƕ<5��<|��<y[�<�5�<��<E�y<��q<7@i<B�`<��X<xP<z;H<�@<,�7<(�/<|^'<u(< �<C�<�}<���;$
�;���;� �;O��;[[�;�;	܉;�~s;�zS;��3;�;Ӑ�:�V�:/[:ݨ�9��̸¹��~��H,���Y���|�^{8�yU�]q�}����<��顡�-��������Ȼ�DԻ�"���뻟����� �0��S�]R��,�S��;z���"��B'�sv+�|�/�I|3��N7�a;��>��
B�DdE���H��K���N���Q���T�:�W�4�Z�\w]��K`��c���e��h�~k��Bn�Eq�I�s��vv��(y�v�{�C}~�6����߁�k-��)z��Mƅ�}��s_��ǭ��
���~P��N���k���CU������m
��e������B��bk����������X��Z����鞼�/�� u�������J��C���E䧼�4������1ݫ�4������䯼C<������과�@������:鷼<��O���y໼�2���  �   O=#UN==�M=2�L=�ML=?�K=|�J=�;J=z�I=�H=�$H=zsG=+�F=TF=gE=��D=�D=iC=a�B=mB=�sA=T�@=l$@=Z{?=��>=(%>=�w==J�<=�<=�h;=S�:=^:=S9=z�8=��7=�:7=��6=��5=�5=�j4=u�3=��2=�B2=��1=��0=�0=@/=�v.=ש-=�,=�,=�,+=lQ*=�r)=��(=�'=��&=B�%=��$=$�#=��"=��!=�� =
�=Y�=�u=i?==�=M�=�U=�=�~=�=k{=��=CN=+�=%�=�D
="�=+�=�=K=E=y��<���<%�<cB�<qU�<_�<.`�<�Y�<�M�<�<�<b(�<��<���<`��<���<���<ۣ�<��<�<Ym�<[�<�G�<�2�<��<E�<&�<�Ǖ<⦑<O��<L`�<f;�<�<��y<�q<�Oi<�	a<u�X<��P<�GH<e@<�7<ښ/<c'<�*<��<��<�y<cw�;���;�~�;T�;���;=�;�;|��;�7s;�4S;l3;��;��:��:�_Z:nw�9��и������7���U���q��g8�\U��9q�N���$��8���G����t����ǻ2+Ի�໽�뻠����� ��+�rQ��Q�.�������"��K'��+�ԕ/��3��]7�(;�.�>��B�tE�ƲH���K��N�d�Q���T�-�W���Z�qz]�M`�c��e��h�'wk��9n���p�A�s�Niv�>y���{��n~�
���ف��'��u���D��H]����������@Q����� ����X��0������`k���ŕ����Gs���ř�����`������C�v5��z�������M��~���䧼/4��I���yګ�D0��+����ޯ�
6��*����㳼h9��4���Mⷼ�5�������ۻ�/���  �  � O=�UN=��M=�L=vML=��K=r�J=r:J=�I=7�H=�"H=4qG=��F=�F=�dE=�D=5D=�fC=b�B=�B=rA=�@=q#@=�z?=��>=(%>=;x==��<=v<=j;=�:=.:=
U9=��8=��7=�<7=ŉ6=�5=�!5=\l4=۵3=��2=�C2=:�1=��0=y0=�?/=v.=��-=��,=,=�*+=NO*=lp)=<�(=��'=W�&=��%=��$=�#=�"=��!=~� =	�=��=�u=\?=��=��=�V=G�=��=�=�}=.�=�P=��=��=$G
=�=N�=��=� =UF=W��<*��<�%�<.B�<�T�<�]�<^�<=W�<mJ�<�8�<$�<1�<���<S��<���<���<��<���<2{�<�i�<@X�<�E�<H1�<��<��<��<�ȕ<���<���<Vc�<?�<5�<��y<{�q<dYi<|a<��X<R�P<�OH<@<U�7<ޞ/<�e'<b,<��<�<�v<o�;��;Rq�; ��;���;~)�;<ۙ;���;.s;�	S;�A3;u�;w��:���:��Y:Ϸ�9	Ӹ�I�r����>���P��qj��[8���T��"q��q��h���v��M����c����ǻ	Ի%�߻ی������ ��(��O�bQ�/�������_�"�uQ'���+���/���3�g7�;�)�>��$B��}E�2�H�o�K���N�2�Q�W�T���W�v�Z��|]��M`��c�M�e�'�h�sk�t4n�(�p���s��`v�}y�Խ{��e~������ԁ��#���q������]���[��竉������Q��>���� ��][��"���Y��Po���ɕ��"��.x���ʙ����qe�����r���"9��C}������7���N��X����䧼�3��3����ث��-��<���ۯ� 2��눲�/߳��4��ĉ��	޷��1��,����ػ��,���  �  ��N=dKN=P�M=A�L=<AL=*�K=<�J=�.J=�|I=R�H=JH=�fG=,�F=�F=XE=��D=��C=�SC=��B=��A=�UA=��@=� @=�T?=�>=��==�J==�<=��;=6;=��:=��9=F9=>e8=֯7=��6=XC6=0�5=�4=�4=u`3=A�2=	�1=[%1=b0=��/=�.=�.=I4-=�_,=�+=y�*=X�)=��(=A(=�'=�+&=�8%=�@$=:C#=>?"=4!=%! =~=u�=��=Rx=S4=^�=��=�&=�=�<=y�=,*=L�=s�=�G=��	=e�=g=jS=ڄ=�� =��<���<g�<�E�<;e�<�{�<"��<^��<���<���<���<�}�<r�<Re�<�X�<NL�< @�<=4�<x(�<`�<��<��<+�<��<^͝<̷�<��<���<�k�<?O�<2�<��<��y<��q<�yi<CAa<Y<4�P<c�H<�u@<�G8<�0<��'<K�<��<�l<v@<�(�;���;+��;/5�;e��;���;���;��;�<y;}�Y;�:;s�;v_�:���:��x:|��9���7����<h�R��E��|���R.�W�J�{sf��Co����������E]��������ͻF�ٻC��z�e��)��,��2�B�[���w�7���V$��(�S�,���0��4��^8��<���?���B�UF���I�P�L���O���R���U�b�X�<�[��^�Q�a�ld�!Dg�?j�(�l���o�Izr�B<u���w�$�z��f}�����a�������m^������a���Y���������|_��˹����[q���͒��)������ޖ�,5������ۚ�b+���x��Ğ�W��X��㡢��주�8��r���G֧�	(���{���Ы��'��'��9ׯ�p/������d߳��6������䷼:�����滼�<���  �  ��N=CKN=>�M=B�L=OAL=T�K=|�J=�.J=�|I=��H=�H=hgG=��F=AF=�XE=��D=��C=�TC=�B= B=VA=ѫ@=� @=U?=�>=��==�J==�<=H�;=�5;=T�:=P�9=�9=�d8=1�7=>�6=�B6=��5=��4=�4=`3=�2=��1=C%1=b0=��/=,�.= .=�4-=I`,=p�+=�*=��)=0�(=�(=�'=P,&=^9%=^A$=�C#=�?"=�4!=n! =�=��=��=Lx=?4=:�=A�=P&=��=e<=�=�)=��=��=G=G�	=��=�=�R=a�=�� ={��<Q��<+�<�E�<?e�<�{�<��<��<d��<ۏ�<���<�~�<Ds�<�f�<9Z�<�M�<_A�<n5�<�)�<Z�<j�<V�<��<0�<�͝<̷�<<C��<�j�<�N�<I1�<��<��y<|�q<�vi<�>a<�Y<��P<a�H<�s@<EF8< 0<��'<��<d�<�l<�@<O*�;���;9��;�8�;���;�Ƭ;`��;癌;�Iy;:�Y;g:;�;,s�:�Ĺ:f
y:��9)��7v��0h�D�����=���U.��J��wf����r������)���.b��������ͻ��ٻ�E�L}�g����
-��2������v�.���U$��(�v�,�R�0���4�e\8��<���?�	�B��RF�c�I�t�L���O���R��U���X���[��^�^�a�ald��Dg�yj���l�#�o�$|r��>u��w��z�3i}����c������_��E������Z���������B_��Q�������p���̒��(�������ܖ��3�������ښ�<*��{w��Þ�k��?W��O���*주c8��J���@֧�)(��|��yѫ�F(�����د�i0�������೼�7��ӎ��!巼;��ܐ���滼>=���  �  ��N=�JN=��M=F�L=�AL=ёK=;�J=�/J=~I=�H=XH=iG=��F=	F=�ZE=p�D=OD=,VC=��B=gB=8WA=��@=�@=uU?=H�>=��==9J==o�<=��;=�4;="�:=��9=19=c8=��7=��6=,A6=�5=1�4=C4=_3= �2=/�1=�$1=�a0=Л/=z�.=�.=Q5-=Ga,=��+=L�*=t�)=��(=�(=j'=.&=;%=C$=ME#=A"=�5!=\" =i= �=ޱ=Ex=�3=��=t�=K%=[�=�:=5�=�'=��=��=E=^�	=��==aQ=�=�� =ԧ�<��<}�<sE�<�e�<�|�<��<Γ�<���<���<��<3��<�v�<{j�<�]�<=Q�<�D�<�8�<x,�<��<��<&�<��<��<�͝<���<=��<
��<Pi�<WL�<�.�<��<��y<��q<�oi<�7a<�Y<6�P<F�H<�n@<B8<�0<G�'<�<�<im<B<�/�;���;���;�C�;`�;լ;´�;]��;;iy; �Y;�1:;��;��:c��:Ocy:�i�9��7��dh����Y��{���].���J��f������}�� ���=���tn��~���r�ͻj�ٻvO�+��m���V.�_3�l����Wt����YQ$��(�ï,��0���4�5U8�^�;�l�?���B��KF��I�øL���O�n�R���U��X���[�c�^��a��md�]Gg��j���l�7�o��r��Du�dx���z��o}����+f������>��a��ȳ������Z��˯��R��r^���������{n��Rʒ��%��O���aٖ�S0�������֚��&��t��򿞼�
���T��f����꣼Y7������(֧��(���|���ҫ�*��!����گ�h3�������㳼V;�����U跼>������黼?���  �  ��N=JN=��M=L�L=�AL=��K=R�J=`1J=�I=C�H=�H=�kG=f�F=�F=�]E=b�D= D=�XC=�B=uB=�XA=$�@=�@=!V?=��>=��==�I==��<=S�;=,3;=B:=��9=�9=g`8=Ȫ7=��6=j>6=��5=��4=>4=S]3=��2=.�1=B$1=�a0=�/=��.=�.=�6-=�b,=��+=��*=��)=��(=v	(=['=�0&=�=%=�E$=�G#=6C"=~7!=�# =�=��=8�=4x=}3=��=/�=�#=T�=�8=��=�$=��=|�=�A=3�	=��=f= O=�=Ϭ =>��<e��<��<CE�<Cf�<2~�<*��<ɖ�<h��<
��<���<���<�|�<�p�<�c�<>W�<�J�<�=�<61�<$�<�<��<���<*�<FΝ<?��<��<��<vf�<�H�<Z*�<��<�y<�q<�ci<�+a<K�X<��P<֓H<of@<;8<'0<]�'<��<I�<Kn<�D<�7�;���;��;jU�;`�;��;^͜;Ì;�y;��Y;�d:;a;X�:|F�:f�y:�+ :���7r��u�g������� ��l.��J�[�f����F����Л��ͨ��������Tλ��ٻy^��w����T0��3������p�����J$�I�(�v�,��0���4�hI8�G�;�Qy?��B��@F��I�y�L��O���R�}�U�~�X�9�[���^���a�pd�,Kg�"j�Z�l�.�o��r��Nu�]x���z��z}�P��k��1�����Bd��J�������[���������)]�������k��Nƒ�:!��K{���Ӗ�r*���~��	њ�� ���n��!���R��;Q��L���W裼�5��鄦�֧�+)��F~���ԫ��,�������ޯ�$8�����Y鳼�@���������B��̗���컼B���  �  ,�N=IN=�M=8�L=`BL=��K=��J=<3J=/�I= �H=�H=oG=��F=�F=taE=�D=�D=\C=��B=B=)[A=�@=�@=�V?=�>=��==%I==q�<=��;=1;=�|:=��9=�9=�\8=;�7=;�6=�:6=8�5=��4=�4=[3=�2=��1=^#1=<a0=�/=��.=�.=8-=�d,=�+=d�*=�)= �(=
(=#'=�4&=�A%=I$=�J#=�E"=�9!=�% =�=��=��=x=�2=��=v�=b!=��=\5=�=� =��=V�=�==-�	=�=�=�K=T~=�� =���<���<"�<�D�<g�< ��<���<���<3��<Ɯ�<.��<���<��<Px�<�k�<�^�<�Q�<�D�<77�<+)�<c�<+
�<e��<��<�Ν<���<I��<>��<�b�<�C�<�$�< �<$�y<;�q<�Ti<�a<��X<εP<-�H<k[@<�18<�	0<�'<��<�<_o<`H<pB�;v��;���;l�;�3�;	�;R�;��;`�y;{)Z;�:;�T;�u�:���:C�z:�� :���7���հg����2�麻���.�l�J��f��"�������電�稻����M» %λ��ٻ�r�̢�[�����V3��4���4���k���@B$�=~(���,�̘0�{x4��:8��;�j?�X�B�w2F��tI���L���O�x�R��U���X�}�[��^��a�Xsd�oPg�7)j�S�l���o�H�r��[u�Dx���z��}�-���q��'ł�9���h�������
��]��r���L���[����������f�����0���t���̖�#��Lw���ɚ�����g��ƴ��� ���L��z���w壼�3��惦�֧�.*��F����׫��0��u����䯼o>������c�H������M���6I�������F���  �  Y�N=�GN=^�M=�L=�BL=�K=J�J=O5J=ބI=�H=e#H=
sG=5�F=F=�eE=n�D=�D=�_C=e�B=	B=�]A=ر@=S@=�W?=5�>=`�==HH==�<=��;=�.;=�y:=d�9=�9=�X8=��7=��6=�66=>�5=2�4=Q4=BX3=��2=*�1=F"1=�`0=�/='�.=�.=�9-=g,=��+=��*=��)=��(=?(=Z''=�8&=�E%=M$=^N#=I"=�<!=�' =l
=��=�=�w=�1=(�=k�=�=`�=�1=ѫ=\=ƃ=f�=�8=l�	=��=�=H={=� =���<���<d�<nD�<�g�<��<��<��<���<&��<���<��<͌�<0��<�t�<�g�<Z�<7L�<�=�<//�<3�<��<���<��<�Ν<���<)��<�|�<^�<7>�<��<���<_�y<�}q<hBi<�
a<H�X<��P<pxH<EN@<�&8<<0<��'<��<��<Ap<�K<kN�;��;���;Յ�;�Q�;�)�;��;�	�;].z;�vZ;D�:;��;���:��:�g{:pb:@�8�)�oxg���2�����l�.���J��f�;��`�������޽��o'»Cλ�ڻ׊�u��}���~�7��6���v���f�����8$��r(���,�ԉ0�h4�d)8�^�;�fX?��B�"F��eI���L�L�O��R���U���X���[�y�^�ԓa�|wd��Vg��1j�%m�r�o�f�r��ku��+x���z�(�}�U$��?y��̂�]���m����������^��������Z��°������a��$���{��m��kĖ�f���n������0���_����������G��3���3⣼�1������0֧��+������p۫�u5��2���민�E��ş�������P�����[����P��&���l����J���  �  =�N=RFN=��M=��L=/CL=u�K=��J=t7J=��I=]�H=-'H=,wG=��F=�F=|jE=�D=1D=�cC=�B=FB=Q`A=�@=�@=�X?={�>= �==PG==|�<=��;=�+;=jv:=��9=�
9=�T8=m�7=Z�6=G26=�{5=H�4=�4=HU3=;�2=E�1=
!1=�_0=�/=��.=�	.=�;-=li,=��+=��*=��)=�(=�(=�+'=�=&=J%=!Q$=+R#=aL"=C?!=�) ==��=5�=�w=�0=��=�=�=�=�-=Q�=p=�~= �=�3=B�	=��=8
=D=�w=�� =��<���<`�<�C�<Bh�<���<M��<���<n��<��<w��<d��<���<���<*~�<�p�<�b�<\T�<*E�<P5�<*$�<��<���<^�<ϝ<C��<���<�x�<�X�<�7�<��<?��<2�y<�jq<�.i<(�`<]�X<�P<RhH<@@<�8<a�/<��'<��<<q<�N<�Z�;�;���;'��;tq�;�L�;�6�;�1�;��z;��Z;�>;;S�;��:���:#8|:�:�8�p߹C@g�m뮺������R�.�8K�#g��U�������(���)��^ൻiI»�cλk,ڻ<�廮�𻤧��\�_;��8�Y����{a���/$��f(�~,��y0�W4�8���;��E?���B�F��UI�}�L�X�O�[�R�\�U���X�Y�[��^�6�a�|d��]g�F;j��m�E�o�ܴr��|u��=x�J�z�a�}�9-�������ӂ�$��Is��A�1�� a�����X���X����������\��򴒼:���d��ֻ��<��;e������E���W��������wA��ʏ���ޣ��/�����|֧� -��f����߫��:��e���I��M��z�������Y��'������X��s�������P���  �   �N=�DN=��M=��L=sCL=X�K=a�J=�9J==�I=��H=�*H=A{G=�F=BF=oE=��D=�D=�gC=��B=WB=�bA=�@="@=hY?=��>=��===F==Œ<=H�;=);=
s:=̼9=j9=P8=Ǚ7=��6=�-6=�w5=B�4=5
4=6R3=��2=P�1=�1=@_0=�/=/�.=�
.=<=-=�k,=i�+=N�*=O�)=D�(=(=e0'=�A&=xN%=<U$=�U#=�O"=�A!=, =�=n�=k�=w=�/=��=��=�=T�=m)=��=�=`y=��=-.=
}	=��=�=�?=t=� =G��<;��<+�<�B�<�h�<���<t��<��<���<ǰ�< ��<��<
��<���<���<�y�<rk�<?\�<1L�<?;�<)�<x�<���<�<�Ν<ܲ�<ޔ�<�t�<�S�<�1�<��<��<�y<*Wq<i<h�`<i�X<��P<�WH<�1@<�8<��/<�'<+�<[�<aq<R<f�;4)�;���;��;���;�o�;�\�;�Y�;��z;�[;�;;�/;��:�:6}:��:�8��޹�g�6鮺��d���.�o@K��Kg��q��[����I��wL������k»߃λ�Jڻg�廲��Y����!�4@�	;���:���\�����%$��Z(��q,�ej0��E4�8�!�;�$3?���B���E�rFI��zL�ÞO�ܴR�<�U�$�X��[���^���a�4�d��eg�Ej��m�k�o���r���u��Ox��
{��}�?6�����fۂ��*��y���Ɔ����Ic�����H��W��q������W��񮒼-��]��7���7��	\��g���q���mO������M퟼<��f����ۣ��-��_���ק��.��k����㫼�?��Ĝ�������U��.����� c��f�������`��󲺼>��hU���  �  �N=3CN=��M=�L=�CL=�K=��J=s;J=��I=��H=0.H=�~G=�F=y!F=asE=��D=�D=�kC=�B=/B="eA=��@=K	@=Z?=��>=�==(E==�<=�;=<&;=�o:=3�9=n9=�K8=g�7=P�6=_)6=�s5=u�4=�4=?O3=C�2=q�1=I1=�^0=��/=��.=�.=�>-=�m,=��+=\�*=��)=)=(=�4'=,F&=vR%=Y$=3Y#=�R"=dD!=�- =�='�=��=xv=�.=�=r~=�=�=�%=^�=�=qt=��=))=x	=�=R=<=�p=3� =���<���<�<�A�<i�<1��<+��<˫�<&��<���<'��<ԯ�<`��<���<3��<W��<^s�<nc�<�R�<�@�<l-�<��<�<W�<uΝ<o��<��<q�<�N�<Y+�<��<��<��y<�Dq<�i<��`<S�X<�pP<}HH<�#@<�8<#�/<��'<v�<��<Vq<�T<�o�;48�;��;���;��;돭;��;~~�;�{;1d[;��;;�r;��:�}�:ʺ}:K:��8t&޹��f��论@�麥���.��fK�&xg�ً������i��_m���$��Ԍ»<�λ�gڻ��������^(�'E�b=��I���X�����$�,P(�e,�P\0�G64���7���;��!?� �B�%�E�V8I�	nL��O�e�R��U��X�D�[�?�^�{�a�m�d��lg��Nj�r+m��p���r��u�ax�q{���}��>������₼K1���~��Tˆ�)���e��4���c���U��8�������LS��]��������U��>�������vS��讀�X����G��Ǘ��M矼7������٣�,����ק��0��e����竼E��آ��� ���]����������k��!¶�R���h��񹺼c
���Z���  �  ?�N=�AN=��M=��L=�CL=��K=��J=�<J=��I=��H=1H=*�G=n�F=%F=�vE=<�D=�D=�nC=��B=�B=gA=�@=D
@=�Z?=��>=|�==D==��<=,�;=�#;=m:=�9=��8=*H8=��7=��6=�%6=�o5=&�4=�4=�L3=�2=��1=1=�]0=f�/=��.=�.=�?-=ho,=!�+=��*=��)=H)={!(=8'=�I&=�U%=.\$=\#=U"=qF!=�/ =�=��=��= v=�-=��=m|=t=�=+"=��=�	=Ap=k�=�$=�s	=�=��=�8=�m=�� =Ë�<���<�<�@�<<i�<j��<p��<!��<u��<,��<7��<g��<i��<���<|��<e��<z�<�i�<	X�<7E�<1�<H�<��<��<Ν<گ�<���<�m�<J�<�%�<��<�݀<�vy<=5q<_�h<��`<�X<JbP<�:H<�@<|�7<��/<W�'<֥<��<?q<�V<Qx�;�D�;|�;m��;�Ž;W��;!��;���;�\{;�[;<;d�;4��:ټ:�U~:}�:� 8�ݹ�f�쮺���&�/�@�K�B�g�6���P6����������tA��è»9�λπڻQ�廁������.��I�@������@U�]���$�8G(�nZ,�P0�)4���7�{�;�|?�(�B���E�,I�pcL��O�<�R�ӳU�ָX��[��^�G�a�&�d�6sg��Vj��5m�Rp���r�#�u��ox��+{���}�
F�����&邼 7������Qφ�0���g��d������$U��e��������O������@����O����������NL��֞����rA��𑞼L⟼�2��\����֣��*������xا�V2�����(뫼}I��-������qd������&���s���ɶ�}���o��2������B_���  �  ��N=�@N=��M=[�L=�CL=�K=��J=$>J=1�I=��H=13H=��G=�F=�'F=�yE=��D=pD=qC=��B=NB=�hA=�@=�
@=�Z?=��>=
�==RC=={�<=��;=";=�j:=��9=W�8=CE8=��7=�6=�"6=9m5=��4=�4=�J3=k�2=e�1=1=]0=(�/=��.=".=�@-=�p,=��+=��*=��)=�)=&$(=�:'=XL&=}X%=�^$=G^#=�V"=�G!=�0 =�=	�=��=�u=�,=X�=�z=y=��=}=��=�=�l=�=q!=�p	=��=��=6=qk=�� =���<u��<x�<4@�<5i�<;��<��<���<���<��<ƿ�<q��<��<���<$��<��<)�<4n�<\�<�H�<�3�<+�<��<A�<�͝<���<���<�j�<�F�<�!�<���<�؀<�jy<�(q<��h<O�`<��X<.WP<{0H<�@<��7<	�/<h�'<_�<��<�p<�W<\~�;)N�;3!�;���;�׽;��;��;���;��{;*�[;�@<;��;�6�:�:��~:�!:��$8S`ݹ��f�]����k4�/��K�D�g������I��s���D���SX��0�»W�λؓڻ)滋�t����3��L�-B�#�#��S�����$��@(�~R,� G0�!4���7�e~;�f?�#{B���E��"I�z[L�i�O���R��U���X�_�[���^���a���d�vxg��]j�F=m��p���r��u�|{x��7{���}��K��V����;��G����҆����qi��b�������T��$��������L��I���0���K������h��F��T���8뛼�<�������ޟ��/������.գ��)������٧��3������L��T���v���i��YƲ�!���y��|϶�3#���t���ĺ����b���  �  ��N=@N=��M=�L=�CL=O�K=��J=�>J=�I=��H=�4H=�G=��F=i)F=b{E=��D=	 D=�rC=�B=jB=[iA=ĺ@=[@=�Z?=w�>=��==�B==��<=��;=� ;=�i:=
�9=��8=zC8=�7=��6=� 6=pk5=�4= 4=gI3=Z�2=��1=t1=�\0=��/=��.=x.=TA-=kq,=��+=
�*=H�)==
)=�%(=g<'=�M&=
Z%=`$=�_#=X"=�H!=k1 ==G�=��=Iu=^,=��=�y=<=)�=�=�=�=�j=��=m=�n	=�=��=x4=�i=�� =���<���<��<�?�<Ni�<͉�<-��<#��<���<���<���<���<1��<���<���<<��<^��<q�<�^�<�J�<I5�<I�<m�<n�<;͝<ĭ�<>��<�h�<ND�<��<���<Հ<Dcy<O!q<�h<��`<{X<�OP<�)H<�@<��7<��/<"�'<1�<��<�p<�X<"��;T�;�(�;��;��;Fͭ;;č;C�{;.�[;b]<;��;Yh�:�G�::*Y:�5'8�,ݹ�f�����}>�e'/��K�D�g������V�����ƭ���e����»�λj�ڻ6�C'�����6�eO��C�������Q�/��V$�{<(�wM,�<A0��4� �7��w;��?��tB���E�0I�nVL�M�O�ƜR���U�:�X�ִ[�4�^��a�9�d��{g��aj�QBm�Lp�@�r�$�u���x��>{���}�kO��ӡ��'�I>�������Ԇ�9���j���������OT��V�������K�������H��\���1�rC�����蛼�9��׊��8ܟ�.������3ԣ�g)��{����٧��4��}����﫼:O������s���l���ɲ��$��}��Ӷ��&��x���Ǻ����e���  �  ��N=�?N=[�M=�L=�CL=b�K=�J="?J=m�I=S�H=�4H=��G=8�F=*F=|E=3�D=� D=sC=��B=�B=�iA=�@=y@=[?=t�>=��==�B==t�<=W�;=h ;=i:=}�9=�8=�B8=.�7=��6=V 6=�j5=s�4=��3=�H3=��2=D�1=71=�\0=�/=��.=�.=�A-=�q,=	�+=i�*=��)=�
)=D&(=='=�N&=�Z%=�`$=`#=vX"=6I!=�1 =C=O�=y�=3u=;,=B�=}y=�=��=O=H�==8j=*�=�=�m	=Z�=M�=�3=�i=0� =��<���<T�<�?�<Xi�<���<���<���<m��<k��<���<���<^��<]��<ѡ�<]��<q��<r�<Q_�<MK�<�5�<��<��<j�<͝<t��<���<Vh�<}C�<�<}��<�Ӏ<�`y<�q<��h<�`<�xX<|MP<�'H<�@<��7<��/<�'<��<V�<�p<IY<r��;�V�;�+�;-�;q�;�ѭ;�Ɲ;�ɍ;<�{;��[;g<;��;fw�:�T�:�%:�l:��'8-!ݹ�f�����)	�5B��+/���K��g��ā��[������{���l����»��λ�ڻ��*�C����7�LP��C������>Q�c��$�;(��K,�X?0��4���7��t;���>�prB�b�E�PI��TL��~O���R��U���X�ϴ[�Y�^�i�a��d��|g�cj�Dm�.p�~�r�{�u��x��A{���}��P�����C�1?������Ն�����j��"������;T��#���*���qJ��f�����"G��A���	B�����曼{8��󉞼u۟�S-������ӣ�A)��{����٧��4������h��O��ݯ��z��n��˲��%���~��fԶ��'��Cy��ɺ�����e���  �  ��N=@N=��M=�L=�CL=O�K=��J=�>J=�I=��H=�4H=�G=��F=i)F=b{E=��D=	 D=�rC=�B=jB=[iA=ĺ@=[@=�Z?=w�>=��==�B==��<=��;=� ;=�i:=
�9=��8=zC8=�7=��6=� 6=pk5=�4= 4=gI3=Z�2=��1=t1=�\0=��/=��.=x.=TA-=kq,=��+=
�*=H�)==
)=�%(=h<'=�M&=
Z%=`$=�_#=X"=�H!=l1 ==I�=��=Ku=a,=��=�y=B=0�=�=�=�=�j=�=|=�n	=�=��=�4=j=�� =ц�<%��<��<�?�<{i�<���<U��<G��<ս�<���<���<���<9��<���<���<1��<N��<q�<n^�<}J�<&5�<#�<E�<E�<͝<���<��<�h�<-D�<��<~��<�Ԁ<+cy<B!q<�h<Ƭ`<{X<
PP< *H<	@<��7<:�/<q�'<��<�<q<8Y<���;�T�;c)�;@�;��;�ͭ;4;.č;4�{;��[;�\<;N�;�f�:sE�:Y	:�S:&�&8(9ݹ]�f�(���$�@��(/���K���g�8����W������U���yf��]�»t�λƠڻ�滉'�����6�{O��C�������Q�8��^$��<(�|M,�@A0��4�#�7��w;��?��tB���E�1I�nVL�M�O�ƜR���U�:�X�״[�4�^��a�9�d��{g��aj�QBm�Mp�@�r�$�u���x��>{���}�kO��ӡ��'�I>�������Ԇ�9���j���������OT��V�������K�������H��\���1�rC�����蛼�9��׊��8ܟ�.������3ԣ�g)��{����٧��4��}����﫼:O������s���l���ɲ��$��}��Ӷ��&��x���Ǻ����e���  �  ��N=�@N=��M=[�L=�CL=�K=��J=$>J=1�I=��H=13H=��G=�F=�'F=�yE=��D=pD=qC=��B=NB=�hA=�@=�
@=�Z?=��>=
�==RC=={�<=��;=";=�j:=��9=W�8=CE8=��7=�6=�"6=9m5=��4=�4=�J3=k�2=e�1=1=]0='�/=��.=".=�@-=�p,=��+=��*=��)=�)=&$(=�:'=XL&=}X%=�^$=H^#=�V"=�G!=�0 =�=�=��=�u=�,=_�=�z=�=��=�=ї=�=m=�=�!=�p	= �=��=>6=�k=� =���<���<��<�@�<�i�<���<g��<��<��<C��<��<���<��<���<��<Ԏ�<
�<
n�<�[�<_H�<l3�<��<k�<��<D͝<M��<W��<zj�<ZF�<z!�<���<^؀<�jy<�(q<��h<g�`<��X<tWP<�0H<@<�7<��/< �'<��<d�<�q<�X<��;AO�;/"�;���;xؽ;���;Y��;ӵ�;��{;��[;�?<;n�;l3�:#�:��~:�:�	$8�wݹ�f�����2�麑7�+/��K�"�g�W���?K������Y���NY���» �λ��ڻ��������3�M�QB�A�<��(S�����$��@(��R,�G0�'4���7�i~;�j?�&{B���E��"I�|[L�j�O���R��U���X�_�[���^���a���d�vxg��]j�G=m��p���r��u�|{x��7{���}��K��V����;��G����҆����qi��b�������T��$��������L��I���0���K������h��F��T���8뛼�<�������ޟ��/������.գ��)������٧��3������L��T���v���i��YƲ�!���y��|϶�3#���t���ĺ����b���  �  ?�N=�AN=��M=��L=�CL=��K=��J=�<J=��I=��H=1H=*�G=n�F=%F=�vE=<�D=�D=�nC=��B=�B=gA=�@=D
@=�Z?=��>=|�==D==��<=,�;=�#;=m:=�9=��8=*H8=��7=��6=�%6=�o5=&�4=�4=�L3=�2=��1=1=�]0=f�/=��.=�.=�?-=ho,=!�+=��*=��)=H)={!(=8'=�I&=�U%=/\$=\#=U"=rF!=�/ =�=��=��=v=�-=��=z|=�=��=@"=��=�	=bp=��=%=t	=C�=��=�8=�m=�� =E��<G��<��<}A�<�i�<���<ݟ�<���<˸�<t��<o��<���<���<���<q��<I��<�y�<ci�<�W�<�D�<�0�<��<F�<��<�͝<k��<(��<;m�<�I�<�%�<L�<�݀<\vy<5q<^�h<�`<-�X<�bP<W;H<�@<0�7<��/<.�'<��<��<%r<�W<�y�;;F�;��;���;�ƽ;��;���;���;�\{;U�[;�<;��;���:~Ӽ:�H~:�:��8B�ݹ[�f��������y*�b	/�|�K�Q�g�"���8��<���C����B���»U�λˁڻ-��@�e����.��I�5@�����]U�u���$�IG(�{Z,�&P0� )4���7���;��?�,�B���E�,I�rcL��O�>�R�ԳU�׸X��[��^�G�a�&�d�6sg��Vj��5m�Rp���r�#�u��ox��+{���}�
F�����&邼 7������Qφ�0���g��d������$U��e��������O������@����O����������NL��֞����rA��𑞼L⟼�2��\����֣��*������xا�V2�����(뫼}I��-������qd������&���s���ɶ�}���o��2������B_���  �  �N=3CN=��M=�L=�CL=�K=��J=s;J=��I=��H=0.H=�~G=�F=y!F=asE=��D=�D=�kC=�B=/B="eA=��@=K	@=Z?=��>=�==(E==�<=�;=<&;=�o:=3�9=n9=�K8=g�7=P�6=_)6=�s5=u�4=�4=?O3=C�2=q�1=I1=�^0=��/=��.=�.=�>-=�m,=��+=\�*=��)=)=(=�4'=-F&=vR%=Y$=4Y#=�R"=gD!=�- =�=,�=��=�v=�.=�=�~==��=�%=|�=�=�t=��=\)=Xx	=U�=�=f<=�p=�� =[��<y��<��<zB�<�i�<���<���<C��<���<L��<l��<��<|��<���<%��<4��<'s�<$c�<MR�<D@�<�,�<"�<��<��<�͝<簙<���<�p�<(N�<�*�<��<��<7�y<�Dq<�i<��`<��X<xqP<IH<�$@<�8<�/<��'<��<�<pr<�U<�q�;:�;[�;*��;?��;Ӑ�;Z��;�~�;S{;Nc[;�;;�p;*{�:�v�:�}:j9:�8&O޹�g�v�6�����.��kK�}g�3�������k��>o��B&��[�»��λ�hڻ������i����(�pE��=�6�t���X����$�@P(�e,�]\0�Q64���7��;��!?�$�B�(�E�Y8I�nL��O�f�R��U��X�E�[�?�^�|�a�m�d��lg��Nj�r+m��p���r��u�ax�q{���}��>������₼K1���~��Tˆ�)���e��4���c���U��8�������LS��]��������U��>�������vS��讀�X����G��Ǘ��M矼7������٣�,����ק��0��e����竼E��آ��� ���]����������k��!¶�R���h��񹺼c
���Z���  �   �N=�DN=��M=��L=sCL=X�K=a�J=�9J==�I=��H=�*H=A{G=�F=BF=oE=��D=�D=�gC=��B=WB=�bA=�@="@=hY?=��>=��===F==Œ<=H�;=);=
s:=̼9=j9=P8=Ǚ7=��6=�-6=�w5=B�4=5
4=6R3=��2=P�1=�1=@_0=�/=/�.=�
.=<=-=�k,=i�+=N�*=O�)=D�(=(=e0'=�A&=xN%==U$=�U#=�O"=�A!=, =�=s�=s�=w=�/=��=Ȁ=�=m�=�)=ע=�=�y=��=g.=I}	=�=�=?@=et=]� =���<���<��<�C�<ni�<T��<	��<i��<p��<)��<m��<$��<*��<��<r��<�y�<5k�<�[�<�K�<�:�<�(�<��<^��<��</Ν<E��<M��<pt�<DS�<1�<��<��<��y<�Vq<i<��`<İX<��P<�XH<t2@<�8<��/<<�'<_�<��<�r<8S<Yh�;R+�;���;���;�;�p�;w]�;�Y�;��z;�[;[�;;%-;���:Y�:��|:��:�8�޹C+g�S���K��x���.�8FK�;Qg�ft�����L���N��f���m»d�λ2Lڻ��廷��:����!��@�N;���j���\����%$��Z(��q,�tj0�F4�8�)�;�*3?���B���E�uFI��zL�ŞO�ݴR�>�U�%�X��[���^��a�4�d��eg�Ej��m�k�o���r���u��Ox��
{��}�?6�����fۂ��*��y���Ɔ����Ic�����H��W��q������W��񮒼-��]��7���7��	\��g���q���mO������M퟼<��f����ۣ��-��_���ק��.��k����㫼�?��Ĝ�������U��.����� c��f�������`��󲺼>��hU���  �  =�N=RFN=��M=��L=/CL=u�K=��J=t7J=��I=]�H=-'H=,wG=��F=�F=|jE=�D=1D=�cC=�B=FB=Q`A=�@=�@=�X?={�>= �==PG==|�<=��;=�+;=jv:=��9=�
9=�T8=m�7=Z�6=G26=�{5=H�4=�4=HU3=;�2=E�1=
!1=�_0=�/=��.=�	.=�;-=li,=��+=��*=��)=�(=�(=�+'=�=&=J%="Q$=,R#=cL"=E?!=* ==��=<�=�w=�0=��=/�=�=��=�-=u�=�=�~=U�=�3=��	=��=�
=aD=�w=U� =͙�<l��<�<�D�<�h�<���<��<��<��<t��<Ǧ�<���<��<���<~�<�p�<�b�<T�<�D�<�4�<�#�<H�<���<��<dΝ<���<��<fx�<}X�<�7�<.�<��<Ѩy<[jq<�.i<W�`<��X<q�P<	iH<�@@<�8<{�/<��'<>�<�<Tr<7P<]�;A�;���;ڢ�;�r�;�M�;|7�;C2�;M�z;��Z;�<;;��;y�:���:�%|:s�:Ơ
8ğ߹�Xg�����X��I����.�5 K��!g��X��9㎻�*���+��U⵻-K»eλ�-ڻs�廼�𻌨�����;��8�������a�9��9/$��f(��,��y0�W4�!8���;��E?���B�
F��UI���L�Z�O�]�R�]�U���X�Z�[��^�7�a�|d��]g�F;j��m�E�o�ܴr��|u��=x�J�z�a�}�9-�������ӂ�$��Is��A�1�� a�����X���X����������\��򴒼:���d��ֻ��<��;e������E���W��������wA��ʏ���ޣ��/�����|֧� -��f����߫��:��e���I��M��z�������Y��'������X��s�������P���  �  Y�N=�GN=^�M=�L=�BL=�K=J�J=O5J=ބI=�H=e#H=
sG=5�F=F=�eE=n�D=�D=�_C=e�B=	B=�]A=ر@=S@=�W?=5�>=`�==HH==�<=��;=�.;=�y:=d�9=�9=�X8=��7=��6=�66=>�5=2�4=Q4=BX3=��2=*�1=F"1=�`0=�/='�.=�.=�9-=g,=��+=��*=��)=��(=?(=Z''=�8&=�E%=M$=`N#=I"=�<!=�' =p
=��=�=�w=�1=6�=|�=�=y�=�1=�=�=�=��=9=��	=��==lH=m{=D� =\��<���<�<E�<Uh�<���<���<���<)��<���<��<��<��<8��<�t�<`g�<�Y�<�K�<�=�<�.�<��<g�<f��<`�<LΝ<�<���<X|�<�]�<�=�<��<G��<�y<k}q<gBi<�
a<��X< �P<!yH<O@<�'8<M0<��'<й<�<|q<�L<�P�;	�;���;y��;�R�;�*�;N�;�	�;&.z;�uZ;��:;-�;���:J�:9V{:�N:I<8W��g�����k����d�.�y�J���f��=���Ď�
���	��ÿ��$)»�Dλ;ڻ��z��^�����j7��6�!�����f�����8$��r(���,��0�#h4�m)8�e�;�lX?��B�"F��eI���L�M�O��R���U���X���[�y�^�ԓa�}wd��Vg��1j�%m�r�o�f�r��ku��+x���z�(�}�U$��?y��̂�]���m����������^��������Z��°������a��$���{��m��kĖ�f���n������0���_����������G��3���3⣼�1������0֧��+������p۫�u5��2���민�E��ş�������P�����[����P��&���l����J���  �  ,�N=IN=�M=8�L=`BL=��K=��J=<3J=/�I= �H=�H=oG=��F=�F=taE=�D=�D=\C=��B=B=)[A=�@=�@=�V?=�>=��==%I==q�<=��;=1;=�|:=��9=�9=�\8=;�7=;�6=�:6=8�5=��4=�4=[3=�2=��1=^#1=<a0=�/=��.=�.=8-=�d,=�+=d�*=�)= �(=
(=#'=�4&=�A%=I$=�J#=�E"=�9!=�% =�=��=��=x=�2=��=��=u!=��=v5=�=!=��=��=�==f�	=W�== L=�~=� =a��<���<��<�E�<�g�<���<|��<��<���<��<t��<��<5��<Wx�<�k�<�^�<�Q�<VD�<�6�<�(�<��<�	�<���<�<Ν<��<Ǜ�<��<2b�<�C�<T$�<��<��y<�q<�Ti<�a<�X<G�P<̇H<+\@<�28<�
0<�'<ý<1�<yp<tI<}D�;\��;k��;�m�;5�;��;��;��;/�y;�(Z;n�:;�R;p�:��:i�z:ެ :b6�7��	�g����(��.��݄.���J��f�+%��ި���뛻�騻j����	»|&λ#�ٻ�s延��$������3�,5���_���k�*��YB$�Q~(�ǚ,�٘0��x4��:8��;�j?�\�B�{2F��tI���L���O�y�R��U���X�}�[��^��a�Xsd�pPg�7)j�S�l���o�H�r��[u�Dx���z��}�-���q��'ł�9���h�������
��]��r���L���[����������f�����0���t���̖�#��Lw���ɚ�����g��ƴ��� ���L��z���w壼�3��惦�֧�.*��F����׫��0��u����䯼o>������c�H������M���6I�������F���  �  ��N=JN=��M=L�L=�AL=��K=R�J=`1J=�I=C�H=�H=�kG=f�F=�F=�]E=b�D= D=�XC=�B=uB=�XA=$�@=�@=!V?=��>=��==�I==��<=S�;=,3;=B:=��9=�9=g`8=Ȫ7=��6=j>6=��5=��4=>4=S]3=��2=.�1=B$1=�a0=�/=��.=�.=�6-=�b,=��+=��*=��)=��(=v	(=['=�0&=�=%=�E$=�G#=7C"=�7!=�# =�=��=>�=;x=�3=��=<�=�#=f�=�8=��=�$=��=��=B=a�	="�=�=:O=I�=� =���<���<�<�E�<�f�<�~�<���<+��<���<R��<���<ه�<�|�<�p�<�c�<"W�<VJ�<�=�<�0�<�#�<��<j�<w��<��<�͝<ж�<���<���<f�<~H�<*�<n�<��y<�q<�ci<�+a<��X<�P<W�H<g@<�;8<�0<4�'<��</�<1o<�E<�9�;J��;h��;�V�;\�;��;�͜;HÌ;�y;��Y;Qc:;�;���:�@�:u�y:A :��7�����g����z�麓��jp.�'�J�i�f�������dқ�Ϩ�_���Z���pλ��ٻU_廁��_x�����0�4���=���p�����J$�Y�(���,���0���4�nI8�L�;�Vy?��B��@F�	�I�{�L��O���R�~�U��X�9�[���^���a�pd�,Kg�"j�Z�l�.�o��r��Nu�]x���z��z}�P��k��1�����Bd��J�������[���������)]�������k��Nƒ�:!��K{���Ӗ�r*���~��	њ�� ���n��!���R��;Q��L���W裼�5��鄦�֧�+)��F~���ԫ��,�������ޯ�$8�����Y鳼�@���������B��̗���컼B���  �  ��N=�JN=��M=F�L=�AL=ёK=;�J=�/J=~I=�H=XH=iG=��F=	F=�ZE=p�D=OD=,VC=��B=gB=8WA=��@=�@=uU?=H�>=��==9J==o�<=��;=�4;="�:=��9=19=c8=��7=��6=,A6=�5=1�4=C4=_3= �2=/�1=�$1=�a0=Л/=z�.=�.=Q5-=Ga,=��+=L�*=t�)=��(=�(=j'=.&=;%=C$=ME#=A"=�5!=^" =k=#�=�=Ix=�3=��=}�=V%=h�=�:=G�=�'=Տ=��=4E=�	=��=<=�Q=E�=�� =0��<y��<��<�E�<�e�<5}�<4��<��<���<ʒ�<��<O��<�v�<j�<�]�<)Q�<�D�<�8�<D,�<��<U�<��<��<��<�͝<>��<�<Ą�<i�< L�<e.�<]�<��y<��q<�oi<�7a<�Y<|�P<��H<o@<�B8<:0<��'<��<��<n<C<�0�;���;���;�D�;�;�լ;��;���;iy;��Y;�0:;��;���:i�:(Zy:rU�9�<�7z2⹢h������麡���`.���J�ˊf�������M���Q���oo��`���;�ͻ�ٻP廲��n��O��.��3������kt����gQ$��(�̯,��0���4�:U8�a�;�o�?���B��KF��I�ĸL���O�o�R���U��X���[�c�^��a��md�]Gg��j���l�7�o��r��Du�dx���z��o}����+f������>��a��ȳ������Z��˯��R��r^���������{n��Rʒ��%��O���aٖ�S0�������֚��&��t��򿞼�
���T��f����꣼Y7������(֧��(���|���ҫ�*��!����گ�h3�������㳼V;�����U跼>������黼?���  �  ��N=CKN=>�M=B�L=OAL=T�K=|�J=�.J=�|I=��H=�H=hgG=��F=AF=�XE=��D=��C=�TC=�B= B=VA=ѫ@=� @=U?=�>=��==�J==�<=H�;=�5;=T�:=P�9=�9=�d8=1�7=>�6=�B6=��5=��4=�4=`3=�2=��1=C%1=b0=��/=,�.= .=�4-=I`,=p�+=�*=��)=0�(=�(=�'=P,&=^9%=^A$=�C#=�?"=�4!=o! =�=��=��=Nx=B4=>�=F�=U&=��=m<=�=�)=��=��=G=X�	=��=�=�R=w�=�� =���<���<[�<�E�<le�<|�<���<��<���<���<̈�<�~�<Ls�<�f�<5Z�<zM�<OA�<X5�<i)�<;�<G�<0�<��<�<^͝<���<ǟ�<��<�j�<rN�<11�<��<l�y<o�q<�vi<�>a<�Y<�P<��H<,t@<�F8<i0<�'<�<��<2m<4A<�*�;8��;���;89�;��;�Ƭ;���;���;�Iy;��Y;�:;p�;vq�:�¹:�y:���9��77��7h������޸�EW.���J�wyf������s��"��������b������ͻ��ٻ F廒}��g��	�-�3�����v�6���U$��(�{�,�U�0���4�g\8��<���?��B��RF�d�I�t�L���O���R��U���X���[��^�^�a�ald��Dg�yj���l�#�o�$|r��>u��w��z�3i}����c������_��D������Z���������B_��Q�������p���̒��(�������ܖ��3�������ښ�<*��{w��Þ�k��?W��O���*주c8��J���@֧�)(��|��yѫ�F(�����د�i0�������೼�7��ӎ��!巼;��ܐ���滼>=���  �  9�N=�AN=�M=8�L=�5L=r�K=o�J=�"J=�pI=�H=�H=B[G=(�F=��E=JE=^�D=a�C=�?C=�B=I�A=`9A=<�@=s�?=�/?=U�>=��====Jk<=��;=�;=QM:=��9=�8=|(8=?p7=f�6=��5=VC5=��4=��3=�3=�L2=��1=�0=��/=�4/=�g.=��-=��,=6�+=�+=1*=QN)=�g(=^}'=��&=��%=�$=Ѧ#=�"=��!=a� =qr=QR=Z)= �="�=<u=%=��=>f=��==��=Cq=��=U?=ę
=V�=a7=5{=P�=��=a =œ�<���<��<"R�<~�<��<S��<���<���<���<���<���<4��<���<���<���<�߽<�ڹ<<յ<�α<Dǭ<���<O��<J��<m��<���<&y�<*f�<�Q�<+<�<�%�<3�<?�y<-�q<^�i<�ma<mEY<�Q<	�H<��@<ض8<��0<y(<�\ <
@<@$<Y	<$��;���;��;Fe�;�N�;�F�;�N�;rj�;?7;��_;��@;o�!;3�;RC�:�}�:�X:`[9ix���F�3z��-Z׺�P���$�ѕ@�Z(\��Qw�����!��h ��^������ǻ��ӻ�@߻�r��[��r���R+�V5
��������*�g{!���%���)���-���1��5��w9��=�#�@�eD�7[G���J���M�p�P��
T��W��Z��]��`���b��e�P�h�y�k��xn��Lq�Rt�d�v���y�k|�S'���J��f���4����U��������>`����������q���Ώ�,��=���擼�A��v���_���yL��d���Z����E�������䟼n3�����cѣ��!��,s��1Ƨ�����p���ǫ�E ��Gy���ү��,��'����߳��8�������鷼:B��n����򻼆K���  �  �N=�AN=�M=5�L=�5L=��K=��J=&#J=BqI=9�H=DH=�[G=��F=;�E=�JE=ۛD=��C=`@C=^�B=��A=�9A=|�@=��?= 0?=c�>=��====-k<=S�;=�;=M:=��9=��8=(8=�o7=��6=X�5=�B5=i�4=��3=w3=rL2=h�1=��0=��/=�4/=�g.= �-= �,=��+=H+=W1*=�N)=3h(=�}'=:�&=3�%=W�$=0�#=M�"=��!=�� =�r=�R=|)=(�=�=&u=�$=��=�e=B�=�~=^�=�p=�=�>=B�
=��=�6=�z=�=��= =S��<c��<��<R�<~�<F��<���<��<[��<���<���<���<#��<���<���<s��<��<�۹<�յ<vϱ<�ǭ<��<���<���<���<���<y�<�e�<1Q�<�;�<=%�<��<z�y<i�q<��i<la<�CY<Q<��H<F�@<��8<��0<�x(<\ <�?<H$<�	<���;���;���;�g�;�Q�;�I�;aR�;�n�;�@;��_;ۗ@;�!;!�;P�:1��:�n:��9#_��6F��w���X׺�P�b�$���@�,\��Uw�=���$��<��n���'���ȻC�ӻ�B߻�t껚]������z+�p5
������<��/�$z!�U�%�^�)�b�-�E�1�M�5��u9��=�Q�@��D��YG�J�J���M�9�P��	T��W��Z��]��`���b���e�L�h���k��yn�Nq�t��v�5�y��l|�)������K���������V��S������H`����������q��OΏ�|+������c哼%A������m���cK��[������D��𔞼䟼�2�������У�X!��s��4Ƨ�����p��Sȫ�� ���y���ӯ�H-������೼�9��m����근�B�����D�
L���  �  y�N=mAN=��M=9�L=�5L=�K=)�J=�#J=rI=9�H=lH=�\G=�F=��E=�KE=4�D=�C=�AC=~�B=��A=�:A=�@=�?=M0?=��>=��==�==�j<=��;=�;=L:=��9=��8=�&8=�n7=��6=�5=�A5=S�4=��3=�3=�K2=�1=��0=��/=�4/=�g.=��-=��,==�+=0+=`2*=�O)=wi(='=��&=��%=��$=p�#=u�"=��!=�� =hs=S=�)=L�=�=�t=�$=��=%e=D�=w}=�=Uo=��=Q==ė
=Z�=u5=~y=��=��=6 =��<p��<4�<�Q�<>~�<��<���<j��<��<���<��<��<���<���<h��<9��<}�<0޹<'ص<jѱ<}ɭ<\��<���<"��<ƚ�<{��<�x�<�d�<�O�<�9�<0#�<9�<[�y<2�q<�i<�fa</>Y<	Q<�H<)�@<^�8<��0<w(<�Z <p?<�$<�
<M��;���;n��;�o�;w[�;�T�;�]�;�z�;BX;��_;ï@;�!;Y�;�u�:���:c�:_X9y����E��r��RZ׺T���$���@��8\��cw�f���-��W��ާ��:���$ȻL�ӻ@J߻�z�%b���  �w,��5
��q��s����w!���%��)���-��1��5�:p9� =��@���C��TG���J���M�$�P��T�W��Z�]�$`��b���e���h�ʣk��}n�KRq��!t��v�N�y��q|��-�"󀼘M��馃�>���>W��!���|��r`��;������p��͏��)������*㓼�>������񗼺H��������`B������
⟼ 1��4����ϣ�� ���r��Ƨ�/���q��\ɫ�"���{���կ��/��{���㳼:<��锶�C�5E��������cM���  �  ��N=�@N=Y�M=2�L=66L=u�K=��J=�$J=rsI=��H=.H=�^G=��F=��E=&NE=W�D=(�C=CC==�B=�A=�;A=&�@=��?=�0?=��>=��==\==j<=ϵ;=� ;=�J:=��9=��8=�$8=�l7=��6=�5=�?5=��4=%�3=L
3=�J2=!�1=#�0=��/=�4/==h.='�-=��,=d�+=�+=
4*=�Q)=pk(=2�'=��&=��%=��$=e�#=0�"=��!=�� ={t=�S=S*=��=�=�t=�#=��=�c=��=�{=�=%m=O�=�:=Y�
=�=E3=tw=�=��=� = ��<���<e�<�Q�<�~�<��<E��<���<���<���<���<(��<��<��<���<���<��<��<�۵<gԱ<̭<Y©<	��<�<���<��<xw�<Bc�<�M�< 7�<��<��<e�y<��q<;�i<�]a<�5Y<+Q<��H<��@<�8<��0<�s(<�X <�><D%<�<p��;e��;.��;'}�;?j�;�d�;�o�;Z��;;`;Z�@;��!;.�;.��:�ߋ:��:�m9:���|�E��k��^׺�Z���$���@�&L\�{w�f���;�����9���9��ȻR�ӻ�U߻����i��_ �R.�d6
�����������7r!�ȹ%�-�)�7�-���1�J�5�eg9�I=�Y�@�s�C�wMG�&�J� �M�S�P��T�rW��Z��]��`��b���e���h��k�уn�4Yq�Q)t��v���y�
z|��5������P��٩�����1Y������]���`��񹋼��;o��ˏ�\'�������ߓ��:��󔖼v헼UD��T����웼x>������ޟ�J.���}��.Σ�w��r�� Ƨ�����r��˫�`$��`~���د�3��L���糼`@�������H��N��������O���  �  m�N=�?N=�M=�L=�6L=#�K=��J=R&J=%uI=��H=�H=daG=��F=~ F=QE=�D=��C=�EC=��B=�A=q=A=z�@=��?=d1?=�>=y�==�==4i<=��;=�:=�H:=Ñ9=F�8=G"8=�i7=��6=r�5=M=5=@�4=�3=�3=RI2=�1=s�0=9�/=�4/=�h.=�-=��,=��+=Y+=$6*= T)=n(=ك'=m�&=d�%=W�$=�#=��"=��!=�� =�u=�T=�*=��=պ=�s=�"=��=%b=��=Hy=]�=@j==�=�7=?�
=��=]0=�t=��=��=3 =P��<��<U�<[Q�<5�<*��<]��<l��<W��<��<n��<b��<���<���<���</��<��<��<�<5ر<Hϭ<�ĩ<θ�<瑱<,��<���<v�<"a�<�J�<�3�<��<��<��y<e�q<�|i<�Ra<�*Y<�Q<S�H<��@<ڥ8<,�0<�o(<rV <�=<�%<�<��;���;��;��;�}�;�z�;��;o��;h�;�B`;�A;��!;�!;(��:1!�:k:-�96���E�=d���b׺�c�^�$�n�@�$f\�H�w��,���N��2/���ʯ� ���+Ȼ��ӻ�d߻���Ot�� ��0�+7
�����@����k!�]�%�u�)��-�J�1�Z�5�\9���<�i}@���C��CG�m�J���M��P���S�!W�Z�]��	`���b���e�`�h�֯k�͋n�dbq�;3t���v�3�y���|�K@�����rU������
���[��q���n	��a���������qm���ȏ�$$�����=ۓ�6������ 藼�>��ʓ��C盼S9��a����ڟ��*��{��̣���`q��5Ƨ�~��St��Oͫ�['�������ܯ��7��\���k쳼�E��U���7����M�����������R���  �  ��N=�>N=[�M= �L=�6L=��K=*�J=�'J=#wI=)�H=$H=JdG=ʳF=�F=ATE=M�D=��C=�HC=�B=M�A=W?A=��@=��?=2?=(�>=<�==4==h<=�;="�:=sF:=1�9=o�8=>8=�f7=ĭ6=]�5=^:5=�4=��3=�3=�G2=Ɇ1=��0=��/=5/=i.=͙-=��,=��+=n+=�8*=�V)=�p(=��'=��&=��%=q�$=ѯ#=(�"=�!=�� =tw=�U=�+=�=��=Is=�!=�=`=4�=wv=A�=�f=��=4=��
=d�=�,=�q=��=w�=, =��<���<��<�P�<��<���<���<���<n��<���<���<f�<��<t �<.��<���<!�<��<3�<�ܱ<�ҭ<�ǩ<���< ��<Y��<Ĉ�<ct�<{^�<JG�<0/�<��<���<b�y<F�q<joi<Ea<�Y<��P<8�H<��@<��8<n�0<�j(<LS <�<<�&<�<��;��;L��;?��;��;t��;���;���;��;�|`;=A;.";�Q;S�:m�:��:wQ9թ��ϋE�=^���j׺/o���$��@���\���w��A��:e���F���⯻%7���AȻ�Ի�v߻͠껭���� ��3��8
������\����d!���%���)�E�-�?�1�{�5��N9���<��p@���C��8G��J��M���P���S�W
W�Z�]�j`���b���e���h�Էk�Q�n��lq��>t��
w���y�e�|�wL�j���Z��V�������^�������
���a��=������[k���ŏ�p ��o{��1֓�[0�������ᗼ#8��L�������y3������՟��&���w���ɣ�v���p��UƧ����;v��Ы��*��B����᯼M=��R�����L������8���"S����������eV���  �  l�N=�=N=��M=��L=7L=��K=c�J=�)J=7yI=��H=�H=[gG=�F=.F=�WE=��D="�C=�KC=ʝB=��A=OAA=}�@=�?=�2?=S�>=��==s==�f<=a�;=�:=�C:=]�9=L�8=�8=Oc7=Z�6=�5=%75=�|4=�3==3=�E2=[�1=��0=>�/=�4/=|i.=��-=R�,=T�+=�+=;*=�Y)=t(=G�'=��&=�%=��$=ݲ#=��"=h�!=�� =y=(W=`,=2�=\�={r=� =E�=�]=��=fs=��=(c=��=-0=��
=��=F)==n=��=��=� =���<K��<S�<qP�<��<%��<#��<��<���<��<��<��<��<x�<D�<���<���<��<��<N�<�֭<�ʩ<���<���<V��<ɇ�<�r�<�[�<iC�<q*�<
�<���<ٽy<2�q<�`i<�6a<�Y<,�P<�H<�@<��8<|0<ue(<�O <;<'<<6 <��;a��;ȵ�;ϫ�;���;y��;�ߏ;��;�`;�wA;�e";�;��:Ի�:ki :L� 9���kcE�~Z���u׺
|���$���@��\�2�w�]X��_}���_��R���*P��ZȻ&Ի��߻���t���� ��6�!:
�H����b{����d]!���%��)�l�-���1�ۊ5��@9���<��b@��C��,G�uJ��M���P���S�wW�6Z��]�K`�Wc� �e�(�h���k���n��xq��Kt�#w���y��|��Y����]`��\���#��Ob��?���r��Xb���������7i��������v���Г�Z*�� ����ڗ�71��c���Xڛ�N-��W���П��"��zt��ǣ����
p���Ƨ����Lx��ӫ��.��􊮼K篼_C��͞��T����R��P������EY��������aZ���  �  ��N=�<N=��M=��L=S7L=I�K=��J=+J=;{I=�H=�H=pjG=X�F=�
F="[E=�D=^�C=�NC=|�B=�A=>CA=��@=�?==3?=s�>=��==�==�e<=��;=��:=xA:=��9=4�8=�8=�_7=�6=��5=�35=�y4=_�3=�3=�C2=�1=��0=��/=�4/=�i.=~�-=��,=�+=�+=�=*=k\)=#w(=��'=P�&=A�%=�$=�#=��"=֦!=�� =�z=HX=�,=_�=�=�q=)=u�=�[=��=Np=d�={_=��=0,=��
=��=�%=�j=��=�=� =���<���<��<�O�<}��<s��<���<b��<���<�<�	�< �<��<e�<-�<Z�<  �<���<��<��<_ڭ<Jͩ<���<ୡ<<��<���<^p�<�X�<o?�<�%�<g�<j�<>�y<�q<3Ri<�'a<�Y<��P<׿H<$�@<7�8<�t0<�_(<+L <m9<�'<i<� <���;���;��;Sÿ;.ȯ;�ڟ;=��;$2�;��`;��A;<�";��;��:,	�:�� :j"9ᖝ��>E�-W����׺��� �$��A��\�6x��n������y��R���i��>rȻ�.ԻӞ߻��t���L ��:��;
�B�����w�e��V!���%���)���-���1��}5�E39��<��U@�2�C�� G��jJ��M�t�P�~�S��W�bZ�%]�,`�Fc���e���h���k�=�n���q�^Xt��%w�f�y�Ĭ|�g����%f��r�������e��빇�3��c��ݸ�����Kg��¿�����-r��~˓�c$���|��ԗ�b*������ӛ�'���y��̟�d��&q���ģ�m��so��ǧ� ���z��:֫��2�����쯼rI��P���7 ���Y��4���J	��b_�������	��~^���  �  G�N=�;N=H�M=@�L=y7L=�K=��J=�,J=}I==�H=<H=<mG=[�F=�F=Q^E=/�D=W D=�QC=�B=!�A=�DA=Y�@=��?=�3?=|�>=3�==�==bd<=�;=��:=?:=Ά9=D�8={8=�\7=��6=h�5=�05=�v4=ݻ3=��2=B2=v�1=��0="�/=�4/=-j.=5�-=��,=��+=�+=�?*=�^)=�y(=��'=o�&=]�%=�$=��#=D�"=�!=�� =|=LY=�-=}�=��=�p=�=��=zY==�=hm=&�=\=@�=s(=��
=��=("=�g=��=��=� =��<��<�<O�<ǀ�<���<���<b��<���<��<��<��<��<��<��<��<�<��<���<��<�ݭ<�ϩ<��<���<���<���<In�<�U�<�;�<� �<�<{�<[�y<!rq<sDi<+a<6�X<U�P<Y�H<�@<Y�8<�m0<>Z(<�H <�7<�'<{<w
 <���;��;���;�ؿ;9�;���;��;KN�;5-a;d�A;��";	�;�Z�:"O�:\!:�#9���"E��V����׺���%��3A�x�\�I7x�����z�������.��#���0�ȻDԻ��߻������{ �)>��=
�������t�k���O!���%�'�)��-��1�1q5�b&9�:�<�8I@���C�TG�"aJ�%�M���P���S���V��Z��]�<`� 
c�%�e���h���k��n���q�cdt��2w�f�y�ù|��s�����k��C������)i��w�������c��帋�����e�� ���p��n���Ɠ�����v���͗�$��Ry���͛�j!���t���ǟ����-n���£�%��
o���ǧ�h!���|��;٫��6��L�����+O��{������N`���������'e��깺�,��ob���  �  ��N=�:N=��M=��L=�7L=Q�K=\�J=�-J=�~I=�H=dH=�oG=�F=YF=�`E=رD=�D=�SC=
�B=��A=sFA=q�@=��?=4?=��>=��====Mc<=��;=�:==:=s�9=��8=�8=�Y7=ˠ6=��5=B.5=St4=��3=��2=r@2=3�1=��0=��/=�4/=[j.=��-=��,=��+=H+=�A*=5a)=`|(=�'=�&=�%=v�$=�#=q�"=�!=� =M}=Z=�-=��=H�=p=�=7�=�W=
�=�j=V�=�X=!�=4%=�
=��=!=�d=*�=[�=� =�|�<���<��<uN�<ހ�<���<_��<���<��<�	�<\�<��<�<=�< �<��<�<��<���<W�<i�<�ѩ<X��<��<���<���<~l�<�R�<H8�<��<l�<E�<5�y<�fq<R8i<ia<��X<Z�P<G�H<�@<�z8<7g0<�U(<VE <6<�'< <� <C�;���;+��;9�;���;�;"0�;�e�;�\a;$B; �";];��:6��:�!:��$9FŜ��
E� X��:�׺P��Q'%��KA��	]�~Yx�����~���ۦ��DD��ǖ��F�Ȼ�VԻz�߻�������  �LA�w?
������r�[��J!�ۈ%�/�)��-�	�1��f5��9���<��>@���C�$G�,YJ�Y�M���P���S�\�V��Z��]�7`�zc��f���h���k�ּn�p�q��nt�^=w��z���|��~���`p��|Ń�H��0l������w���d������$d���������j����T���q���ȗ�����s���ț����=p���ß�����k������0���n���ǧ��"���~���۫��9��8�������2T��Ѱ��'��	f��.������:j������+���e���  �  ��N=�9N=�M=��L=�7L=��K=�J=�.J=�I=�H=!H=oqG=��F=gF=cE=�D=�D=�UC=��B=G�A=�GA=H�@=L�?=^4?=��>=��==}==ob<=p�;=��:=_;:=��9=��8=�8=�W7=��6=��5=5,5=zr4=�3=S�2=4?2=4�1=��0=!�/=g4/=zj.=3�-=d�,=��+=�+=:C*=�b)=/~(=�'=�&=��%=i�$=�#=�"=S�!=?� =1~=�Z=M.=��=�={o=�=�=V=U�=�h=:�=�V=��=�"=,}
=m�=�=�b=0�=��=8 =Ez�< ��<��<�M�<���<_��<���<���<���<��<��<��<�<r�<W�<�<��<!�<���< �<|�<^ө<H¥<[��<x��<���<k�<�P�<�5�<��<���<V�<x�y<�]q< /i<>a<��X<�P<��H<�@<�t8<Mb0<�Q(<�B <�4<�'<7<N <��;���;+��;$��;p�;��;$B�;0x�;3�a;�8B;�#;�*;|��:F��:�":��%9������D�Z���׺د�Y6%��^A��!]�Qsx�4���hі�<����T�������Ȼ�dԻ��߻��I����# ��C�A
��-���o�C��F!���%�!�)���-���1��^5�K9�)�<��6@��C�7G�"SJ��M�p�P���S�_�V�@Z�U]��`�/c��f���h���k���n���q�wt��Ew��z���|� �����s���ȃ����n���������re���������c��i���d���g��p������n���ė�����o���ě�����l���������i������n���n��_ȧ��#��C���ޫ�<��T�������W������q��pj��{¶���n��
º�V��lh���  �  '�N==9N=M=��L=�7L=�K=_�J=//J=x�I=i�H=
"H=�rG=�F=�F=TdE=�D=�D=�VC=��B=$�A=;HA=˗@=��?=�4?=q�>=O�====�a<=��;=��:=Y::=��9=p�8=V8=NV7=C�6=2�5=�*5=@q4=Ҷ3=]�2=e>2=�1=��0=��/=D4/=�j.=x�-=��,=q�+=L +=-D*=�c)=V(=8�'=K�&=5�%=��$=�#=�"=@�!=�� =�~=[=.=��=Ǹ=o=G=K�=0U=;�=�g=��=+U=,�=.!=�{
=��=[=Ra=��=��=V =�x�<��<��<�M�<��<Ϋ�<���<��<$��<��<��<�<�!�<!�<��<��<I�<M�<���<��<��<6ԩ<�¥<��<2��<��<j�<�O�<�3�<��<w��<�߀<�y<�Wq<c)i<�`<�X<��P<��H<ȅ@<9q8<p_0<�O(<9A <�3<w'<<� <8�;��;���;��;N�;�&�;M�;���;c�a;�NB;�/#;�=;h��:Hэ:`,":�;&9�V����D��\���׺~���?%�nkA��0]�܄x�ɯ���ۖ�����_��S����Ȼ%nԻ�߻a��]���& ��E��A
�t�����n�z���C!�m�%�4�)���-�Ӌ1��Y5�19�
�<��1@�Q�C��G�/OJ��M���P���S�3�V��
Z��]��`��c�-f���h�z�k���n���q�C|t�?Kw��z��|�W�����Sv���ʃ�����o����������e��*���F��fb��j�����(f��m�������k������bm��:�����j���������h��þ������n���ȧ�G$��<���N߫�->��I���E���yZ������#��m��.Ŷ�����p��Wĺ�S��!j���  �  ��N=9N=��M=��L=�7L=�K=w�J=i/J=��I=��H=Y"H=�rG=��F=F=�dE=��D=mD=2WC=�B=o�A=zHA=��@=��?=�4?=q�>=@�==�==�a<=u�;=��:=	::=�9=�8=�8=�U7=��6=��5=�*5=�p4={�3=�2=>2=[1=V�0=��/=:4/=�j.=��-=��,=��+=� +=yD*==d)=�(=��'=��&=��%=�$=w�#=i�"=��!=9� =�~=8[=�.=��=��=�n==�=�T=��=?g=e�=�T=��=� ={
=n�=�=�`=��=9�= =Wx�<���<��<�M�<#��<��<���<���<���<!�<��<��<w"�<�!�<��<k�<�<��<b��<
�<1�<lԩ<�¥<���<��<Ƃ�<�i�<
O�<E3�<!�<���<�ހ<G�y<�Uq<'i<]�`<^�X< �P<�H<w�@<�o8<X^0<�N(<�@ <�3<�'<d<> <<�;�;��;��;��;z*�;�P�;r��;�a;uVB;�5#;1C; �:dڍ:~;":U&9NL��:�D�V^���׺��&D%��pA�d5]��x�粉��ޖ��ţ�_c�� �����Ȼ@qԻ��߻��������& �8F�BB
�������n����}B!�U%���)�\�-��1��W5��9�[�<��/@���C�� G��MJ�ыM���P�$�S� �V��
Z��]�'`��c�#	f��h���k�S�n�(�q��}t�Mw��z�#�|���p ��w���˃�����p������f��/���,��Eb���������e��Ҽ������j��6������l��_������>j��q��� ��Jh����������n���ȧ�|$�������߫��>��睮�����B[��h�����/n��1ƶ����\q��ź�����j���  �  '�N==9N=M=��L=�7L=�K=_�J=//J=x�I=i�H=
"H=�rG=�F=�F=TdE=�D=�D=�VC=��B=$�A=;HA=˗@=��?=�4?=q�>=O�====�a<=��;=��:=Y::=��9=p�8=V8=NV7=C�6=2�5=�*5=@q4=Ҷ3=]�2=e>2=�1=��0=��/=D4/=�j.=x�-=��,=q�+=L +=-D*=�c)=V(=8�'=K�&=5�%=��$=�#=�"=@�!=�� =�~=[=�.=��=ɸ=o=J=O�=5U=@�=�g=��=4U=5�=9!=�{
=��=i=aa=�=��=h = y�<0��<��<�M�<2��<��<���<��<<��<��<�<$�<�!�<!�<��<��<=�<=�<���<l�<��<ԩ<�¥<a��<��<備<�i�<|O�<�3�<��<e��<�߀<܉y<�Wq<c)i<��`<�X<ùP<˝H<�@<jq8<�_0<�O(<vA <4<�'<Q< <��;�;H �;A�;��;�&�;!M�;���;0�a;qNB;n/#;�<;���:ύ:d(":�*&9�_����D�p_��a�׺����@%��lA��1]���x�J����ۖ�����_������A�ȻnnԻC�߻��껍���"& ��E�B
�������n�����C!�r�%�8�)���-�Ջ1��Y5�39��<��1@�R�C��G�/OJ��M���P���S�3�V��
Z��]��`��c�-f���h�z�k���n���q�C|t�?Kw��z��|�W�����Sv���ʃ�����o����������e��*���F��fb��j�����(f��m�������k������bm��:�����j���������h��þ������n���ȧ�G$��<���N߫�->��I���E���yZ������#��m��.Ŷ�����p��Wĺ�S��!j���  �  ��N=�9N=�M=��L=�7L=��K=�J=�.J=�I=�H=!H=oqG=��F=gF=cE=�D=�D=�UC=��B=G�A=�GA=H�@=L�?=^4?=��>=��==}==ob<=p�;=��:=_;:=��9=��8=�8=�W7=��6=��5=5,5=zr4=�3=S�2=4?2=4�1=��0=!�/=g4/=zj.=3�-=d�,=��+=�+=:C*=�b)=/~(=�'=�&=��%=i�$=�#=�"=T�!=@� =3~=�Z=O.=��=�=�o=�=�=(V=_�=�h=I�=�V=��=�"=C}
=��=�=�b=O�=��=Z =�z�<f��<��<;N�<:��<���<���<��<���<��<��<��<(�<v�<Q�<��<��<�<���<��<J�<'ө<¥<��<=��<]��<�j�<�P�<�5�<��<���<<�<T�y<x]q< /i<Oa<��X<D�P<�H<o�@<Uu8<�b0<SR(<=C <E5<
(<�<� <|�;� �;���;���;��;9�;>B�;$x�;πa;�7B;�#;�);{��:ѳ�:��!:&�%9t���@E��^��ޮ׺<���8%�aA��#]�gux�.���PҖ�����U�������ȻCeԻ�߻|�껦����# �D�"A
�+�A��	p�Q��F!���%�)�)��-���1��^5�N9�+�<��6@��C�8G�#SJ��M�q�P���S�_�V�@Z�U]��`�/c��f���h���k���n���q�wt��Ew��z���|� �����s���ȃ����n���������re���������c��i���d���g��p������n���ė�����o���ě�����l���������i������n���n��_ȧ��#��C���ޫ�<��T�������W������q��pj��{¶���n��
º�V��lh���  �  ��N=�:N=��M=��L=�7L=Q�K=\�J=�-J=�~I=�H=dH=�oG=�F=YF=�`E=رD=�D=�SC=
�B=��A=sFA=q�@=��?=4?=��>=��====Mc<=��;=�:==:=s�9=��8=�8=�Y7=ˠ6=��5=B.5=Rt4=��3=��2=r@2=3�1=��0=��/=�4/=[j.=��-=��,=��+=H+=�A*=5a)=`|(=�'=�&=�%=w�$=�#=r�"=�!=� =O}=Z=�-=��=N�=p=�=A�=�W=�=�j=j�=Y=;�=Q%=�
=�=H=�d=V�=��=� =�|�<C��<
�<�N�<<��<��<���<6��<O��<�	�<��<
�<�<B�<�<��<�
�<y�<��<�<"�<�ѩ<��<���<e��<2��</l�<�R�<8�<��<<�<�<�y<xfq<R8i<�a<��X<��P<��H<��@<X{8<�g0<8V(<�E <�6<P(<�<Z <l�;���;��;��;s��;u�;H0�;�e�;M\a;*B;��";�;���:T��:,�!:X�$9gޜ��E��^���׺����*%�OA�]�p\x� �����
���XE������%�Ȼ}WԻ'�߻o�����V  �|A��?
�����r�n��.J!��%�:�)��-��1��f5��9���<��>@���C�&G�-YJ�[�M���P���S�]�V��Z��]�7`�zc��f���h���k�ּn�p�q��nt�^=w��z���|��~���`p��|Ń�H��0l������w���d������$d���������j����T���q���ȗ�����s���ț����=p���ß�����k������0���n���ǧ��"���~���۫��9��8�������2T��Ѱ��'��	f��.������:j������+���e���  �  G�N=�;N=H�M=@�L=y7L=�K=��J=�,J=}I==�H=<H=<mG=[�F=�F=Q^E=/�D=W D=�QC=�B=!�A=�DA=Y�@=��?=�3?=|�>=3�==�==bd<=�;=��:=?:=Ά9=D�8={8=�\7=��6=h�5=�05=�v4=ݻ3=��2=B2=v�1=��0="�/=�4/=-j.=5�-=��,=��+=�+=�?*=�^)=�y(=��'=o�&=^�%=�$=��#=E�"=�!=�� =|=OY=�-=��=��=�p=�=��=�Y=O�=}m=?�=\=`�=�(=�
=(�=X"=�g=�=��=� =��<���<��<�O�<:��<��<��<���<��<��<�<�<��<��<��<��<��<���<h��<��<\ݭ<fϩ<���<-��<���<2��<�m�<?U�<F;�<� �<��<M�<�y<rq<sDi<Ja<t�X<��P<ϴH<x�@<��8<Dn0<[(<]I <l8<u(<H<: <��;J��;���;�ٿ;��;G��;��;7N�;�,a;2�A;��";��;�U�:&I�:�N!:��#9�=��2E�_��٘׺Μ�+%��7A�E�\��:x�7������u���0��T���A�Ȼ�DԻ��߻d�껰���� �d>��=
������t�����O!���%�4�)��-�
�1�8q5�h&9�?�<�<I@���C�WG�$aJ�&�M���P���S���V��Z��]�<`�!
c�&�e���h���k��n���q�cdt��2w�f�y�ù|��s�����k��C������)i��w�������c��帋�����e�� ���p��n���Ɠ�����v���͗�$��Ry���͛�j!���t���ǟ����-n���£�%��
o���ǧ�h!���|��;٫��6��L�����+O��{������N`���������'e��깺�,��ob���  �  ��N=�<N=��M=��L=S7L=I�K=��J=+J=;{I=�H=�H=pjG=X�F=�
F="[E=�D=^�C=�NC=|�B=�A=>CA=��@=�?==3?=s�>=��==�==�e<=��;=��:=xA:=��9=4�8=�8=�_7=�6=��5=�35=�y4=_�3=�3=�C2=�1=��0=��/=�4/=�i.=~�-=��,=�+=�+=�=*=k\)=#w(=��'=P�&=A�%=�$=�#=±"=צ!=�� =�z=KX=-=e�=�=�q=5=��=�[=��=ep=�=�_=�=X,=ˆ
=��=�%=	k=Щ=Z�=� =���<,��<@�<RP�<���<��<���<���<P��<[�<�	�<J�<��<l�<"�<=�<���<]��<��<y�<�٭<�̩<��<m��<Ț�<H��<�o�<$X�<?�<E%�<$�<7�<��y<�q<2Ri<(a<�Y<B�P<\�H<Ĥ@<�8<wu0<�`(<M <X:<p(<N<\ <���;i��;A��;SĿ;�ȯ;2۟;p��;2�;��`;/�A;Y�";C�;��:�:�� :~)"96���qPE�\`���׺2���%�<A�?�\�<x��p��ɗ��J{�����:k��osȻ�/Ի��߻���'���� ��:�<
�q�����w����/V!���%�»)���-���1��}5�K39��<��U@�5�C�� G��jJ��M�v�P��S��W�cZ�%]�,`�Gc���e���h���k�=�n���q�^Xt��%w�f�y�Ĭ|�g����%f��r�������e��빇�3��c��ݸ�����Kg��¿�����-r��~˓�c$���|��ԗ�b*������ӛ�'���y��̟�d��&q���ģ�m��so��ǧ� ���z��:֫��2�����쯼rI��P���7 ���Y��4���J	��b_�������	��~^���  �  l�N=�=N=��M=��L=7L=��K=c�J=�)J=7yI=��H=�H=[gG=�F=.F=�WE=��D="�C=�KC=ʝB=��A=OAA=}�@=�?=�2?=S�>=��==s==�f<=a�;=�:=�C:=]�9=L�8=�8=Oc7=Z�6=�5=%75=�|4=�3==3=�E2=[�1=��0=>�/=�4/=|i.=��-=R�,=T�+=�+=;*=�Y)=t(=G�'=��&=�%=��$=޲#=��"=j�!=�� =y=,W=d,=8�=d�=�r=� =S�=�]=��=~s=��=Hc=��=W0=̊
=��=})=yn=�=�=3 =(��<���<��<�P�<���<���<���<v��<��<N��<��<��<��<~�<8�<u��<i��<g�<B�<��<B֭<"ʩ<@��<~��<ߚ�<T��<r�<#[�<
C�<*�<��<��<��y<�q<�`i<�6a<Y<��P<��H<��@<E�8<�|0<Xf(<�P <<<(<�< <���;���;��;٬�;���;���;��;��;�`;�vA;�c";��;��:봌:Z :g� 9|A���uE��c��׺Ӏ���$���@�M�\�\�w�QZ��0���a�������Q��U[Ȼ=Ի��߻���-���@ �7�[:
�x�����{����{]!���%��)�y�-���1��5��@9���<��b@��C��,G�uJ���M���P���S�xW�7Z��]�K`�Xc� �e�(�h���k���n��xq��Kt�#w���y��|��Y����]`��\���#��Ob��?���r��Xb���������7i��������v���Г�Z*�� ����ڗ�71��c���Xڛ�N-��W���П��"��zt��ǣ����
p���Ƨ����Lx��ӫ��.��􊮼K篼_C��͞��T����R��P������EY��������aZ���  �  ��N=�>N=[�M= �L=�6L=��K=*�J=�'J=#wI=)�H=$H=JdG=ʳF=�F=ATE=M�D=��C=�HC=�B=M�A=W?A=��@=��?=2?=(�>=<�==4==h<=�;="�:=sF:=1�9=o�8=>8=�f7=ĭ6=]�5=^:5=�4=��3=�3=�G2=Ɇ1=��0=��/=5/=i.=̙-=��,=��+=n+=�8*=�V)=�p(=��'=��&=��%=r�$=ү#=*�"=��!=�� =vw=�U=�+=�=��=Rs=�!=�=0`=H�=�v=]�=�f=��=F4=��
=��=1-=�q=�=��=n =���<W��<v�<�Q�<2��<��<&��<��<���<-��<(��<��<�<z �<#��<���<��<d�<��<Rܱ<�ҭ<4ǩ<N��<���<嚝<S��<�s�<^�<�F�<�.�<V�<���<�y<"�q<ioi<2Ea<Y<��P<��H<T�@<Q�8<:�0<�k(<2T <�=<�'<k<���;���;���;y��;��;5��;s��;���;}�;�{`;�;A;%,";TO;@M�:Yf�:�:�9)̞���E�kg��#t׺�s�L�$���@���\���w�dC���f��_H��:䯻y8��CȻ�Ի�w߻���`��� ��3��8
������|����d!���%���)�Q�-�I�1���5��N9���<��p@���C��8G��J��M� �P���S�W
W�Z�]�k`���b���e���h�շk�Q�n��lq��>t��
w���y�e�|�wL�j���Z��V�������^�������
���a��=������[k���ŏ�p ��o{��1֓�[0�������ᗼ#8��L�������y3������՟��&���w���ɣ�v���p��UƧ����;v��Ы��*��B����᯼M=��R�����L������8���"S����������eV���  �  m�N=�?N=�M=�L=�6L=#�K=��J=R&J=%uI=��H=�H=daG=��F=~ F=QE=�D=��C=�EC=��B=�A=q=A=z�@=��?=d1?=�>=y�==�==4i<=��;=�:=�H:=Ñ9=F�8=G"8=�i7=��6=r�5=M=5=@�4=�3=�3=RI2=�1=s�0=9�/=�4/=�h.=�-=��,=��+=Y+=$6*= T)=n(=ڃ'=m�&=e�%=X�$=�#=��"=��!=�� =�u=�T=�*=��=ۺ=t=�"=��=4b=��=]y=u�=]j=]�=�7=g�
=�=�0=�t=��=�=n =ɍ�<���<��<�Q�<��<���<���<���<���<\��<���<���<���<���<|��<��<��<��<�ߵ<�ױ<�έ<pĩ<j��<���<Ś�<2��<�u�<�`�<qJ�<;3�<n�<}�<��y<E�q<�|i<�Ra<+Y<Q<��H<�@<�8<�0<{p(<@W <�><�&<�<���;��;H��;��;�~�;\{�;r��;���;@�;QB`;UA;��!;r;���:5�:�]:>�9�T��'�E�yl���j׺�g�q�$�c�@��i\��w��.��~P���0��E̯�>!���,Ȼ��ӻ�e߻E���t��] ��0�]7
�H����^��0��k!�m�%���)���-�S�1�a�5�\9���<�m}@���C��CG�o�J���M��P���S�"W�Z�]��	`���b���e�`�h�֯k�΋n�dbq�;3t���v�3�y���|�K@�����rU������
���[��q���n	��a���������qm���ȏ�$$�����=ۓ�6������ 藼�>��ʓ��C盼S9��a����ڟ��*��{��̣���`q��5Ƨ�~��St��Oͫ�['�������ܯ��7��\���k쳼�E��U���7����M�����������R���  �  ��N=�@N=Y�M=2�L=66L=u�K=��J=�$J=rsI=��H=.H=�^G=��F=��E=&NE=W�D=(�C=CC==�B=�A=�;A=&�@=��?=�0?=��>=��==\==j<=ϵ;=� ;=�J:=��9=��8=�$8=�l7=��6=�5=�?5=��4=%�3=L
3=�J2=!�1=#�0=��/=�4/==h.='�-=��,=d�+=�+=
4*=�Q)=pk(=2�'=��&=��%=��$=e�#=1�"=��!=� =}t=�S=W*=��=�=�t=�#=��=�c=��=�{="�=<m=i�=;=z�
='�=l3=�w=�=#�= =c��<T��<��<R�<�<C��<���<���<��<��<���<F��<*��<��<���<���<v�<��<v۵<'Ա<�˭<©<���<���<���<Ɖ�<)w�<�b�<oM�<�6�<��<i�<1�y<��q<:�i<^a<6Y<uQ<5�H<?�@<r�8<M�0<mt(<�Y <v?<�%<L<���;���;8��;~�;�j�;�e�;@p�;���;�~;}`;`�@;+�!;i�;��:�ڋ:�:�>9]Ο���E��r���d׺'^��$�Ǵ@�@O\� ~w����;=�����M���2���Ȼ�ӻSV߻@��sj��� ��.��6
������ǆ��Gr!�ֹ%�8�)�@�-���1�P�5�jg9�M=�\�@�v�C�yMG�(�J�!�M�T�P��T�sW��Z��]��`��b���e���h��k�уn�4Yq�Q)t��v���y�
z|��5������P��٩�����1Y������]���`��񹋼��;o��ˏ�\'�������ߓ��:��󔖼v헼UD��T����웼x>������ޟ�J.���}��.Σ�w��r�� Ƨ�����r��˫�`$��`~���د�3��L���糼`@�������H��N��������O���  �  y�N=mAN=��M=9�L=�5L=�K=)�J=�#J=rI=9�H=lH=�\G=�F=��E=�KE=4�D=�C=�AC=~�B=��A=�:A=�@=�?=M0?=��>=��==�==�j<=��;=�;=L:=��9=��8=�&8=�n7=��6=�5=�A5=S�4=��3=�3=�K2=�1=��0=��/=�4/=�g.=��-=��,=<�+=0+=`2*=�O)=wi(='=��&=��%=��$=p�#=v�"=��!=�� =is=S=�)=O�=!�=�t=�$=��=.e=O�=�}=&�=eo=��=f==ۗ
=s�=�5=�y=ض=��=Y =[��<���<z�<:R�<�~�<#��<۽�<���<G��<���<-��<0��<���<���<b��<*��<e�<޹< ص<<ѱ<Jɭ<%��<a��<模<���<A��<Rx�<�d�<�O�<�9�<#�<�<7�y< �q<�i<�fa<S>Y<=Q<F�H<|�@<��8<d�0<xw(<6[ <�?<7%<=<0��;���;*��;�p�;�[�;�T�;^�;�z�;+X;t�_;�@;�!;�;�r�:7��:��:�69>/���F�]w��_׺iV���$�Σ@��:\��ew�`���.��-�����������Ȼ��ӻ�J߻>{껂b���  ��,��5
�'���������w!���%��)���-��1��5�>p9�#=��@���C��TG���J���M�$�P��T�W��Z�]�$`��b���e���h�ʣk��}n�KRq��!t��v�N�y��q|��-�"󀼘M��馃�>���>W��!���|��r`��;������p��͏��)������*㓼�>������񗼺H��������`B������
⟼ 1��4����ϣ�� ���r��Ƨ�/���q��\ɫ�"���{���կ��/��{���㳼:<��锶�C�5E��������cM���  �  �N=�AN=�M=5�L=�5L=��K=��J=&#J=BqI=9�H=DH=�[G=��F=;�E=�JE=ۛD=��C=`@C=^�B=��A=�9A=|�@=��?= 0?=c�>=��====-k<=S�;=�;=M:=��9=��8=(8=�o7=��6=X�5=�B5=i�4=��3=w3=rL2=h�1=��0=��/=�4/=�g.= �-= �,=��+=H+=W1*=�N)=3h(=�}'=:�&=3�%=W�$=1�#=M�"=��!=�� =�r=�R=})=)�= �=(u= %=��=�e=G�=�~=e�=�p="�=�>=N�
=��=�6=�z=��=��= =w��<���<��<1R�<(~�<g��<˼�<��<r��<���<���<���<)��<���<���<l��<��<�۹<�յ<_ϱ<�ǭ<���<���<d��<d��<���<�x�<�e�<Q�<�;�<+%�<v�<h�y<`�q<��i<la<�CY<"Q<��H<q�@<ĵ8<Ԗ0<%y(<I\ <@<�$<�	<��;��;��;h�;R�;J�;�R�;�n�;�@;��_;��@;c�!;{�;�N�:g��:�j:Q�9Vh��F��y��6[׺*R���$��@�@-\��Vw����U%�����Ӟ������jȻ��ӻC߻�t��]�������+�5
������E��6�*z!�Z�%�b�)�f�-�H�1�O�5��u9��=�R�@��D��YG�J�J���M�9�P��	T��W��Z��]��`���b���e�L�h���k��yn�Nq�t��v�5�y��l|�)������K���������V��S������H`����������q��OΏ�|+������c哼%A������m���cK��[������D��𔞼䟼�2�������У�X!��s��4Ƨ�����p��Sȫ�� ���y���ӯ�H-������೼�9��m����근�B�����D�
L���  �  `�N=9N=@�M=��L=�*L=zK=��J=�J=�dI=��H=P H=@NG={�F=#�E=d:E=�D=5�C=�*C=p{B=;�A=�A=�l@=��?=~?=vY>=��==��<=�=<=��;=��:=:=e`9=�8=��7=27=Nv6=��5=�4==4=�|3=�2=Z�1=�11=Ni0=��/=��.=��-=�+-=`T,=Uy+=��*=>�)=��(=��'=S�&=�&=Q%=�$=I#=�	"=�� =�=��=�=�z=qE=1=��=�n=�=��=�A=��=J=r�=�/=ԕ=��	=�J=��=�=�#=)_=1)�<}��<���<�&�<-g�<h��<��<+��<7�<Z.�<C�<hS�<4`�<�i�<�q�<w�<D{�<O~�<��<��<���<�~�<�{�<Cw�<�p�<�h�<?_�<�S�<LG�<U9�<�*�<�<4�<��y<Y�q<	�i<�a<��Y<�fQ<^OI<�9A<�%9<�1<D)<B� <��<D�<��<-� <A��;
�;���;��;峱;��;$�;�z�;��e;`�F;t(;7�	;oP�:��:�e<:�?�9��@� %�Kb����ź�m���>�!�6��:R��!m�̃� ͐�������@V���S»�λٻK��g�ﻁ5���I�vW��D���-�� N����m#� G'�i`+�0]/�N?3��7��:��K>���A��7E� �H���K��O��<R��\U��rX�!�[�d�^��a�|d��mg�*Zj�`@m�}!p���r���u��x�lp{�:8~�9~���ށ��=����������V��	���,���m���ˌ�b*�����萼�F��Ӥ��:��f^��j�������j����������i���������b������	���^��㴧���Ud��x������8r��Dͯ��(�������޳��9��s����8I���������$Y���  �  2�N=�8N=2�M=��L=�*L=zK=��J=,J=eI=زH=� H=�NG=ϜF=x�E=�:E=Y�D=��C=+C=�{B=r�A=�A=.m@=��?=�?=�Y>=�==|�<=y=<=y�;=��:=�:=+`9=Ȧ8=��7=�17=v6=^�5=��4=�<4=�|3=ֺ2=,�1=c11=<i0=n�/=��.= .=�+-=�T,=�y+=�*={�)=:�(=�'=��&=�&=�%=A$=�#=�	"=� =L�=%�=�=�z=|E=.=��=cn=�=[�=�A=p�=3J=�=f/={�=��	=J=a�=��=x#=�^=�(�<��<���<�&�< g�<s��<<��<o��<��<�.�<�C�<�S�<�`�<�j�<r�<�w�<�{�<�~�<���<���<��<p�<=|�<�w�<q�<�h�<-_�<�S�<�F�<9�<*�<��<�
�<x�y<$�q<Ƿi<��a<6Y<�eQ<:NI<�8A<�$9<1<�)<�� <a�<G�<��<�� <̄�;��;o��;]��;b��;��;�&�;A}�;��e;�F;N(;��	;tY�:n�:`v<:�\�9��@���$��a��еź#o���@���6�>R�?$m��̓�Gϐ�풝����WX���U»nλ�ٻ��仡�ﻏ6��2J��W��D�A����EM�����#�F'�%_+�\/��=3�t7�̳:�SJ>���A�@6E��H�#�K�O��;R�N\U��rX��[�Ʌ^�h�a��|d��ng��Zj�Am�p"p���r�&�u�)�x��q{��9~��~�� ߁�>�����]���IV��2���O���m���ˌ�*�������琼)F��I�������]���������i��D���S��Zi������|��cb��Ƶ���	���^��촧�)��{d��ҽ������r���ͯ�)��a���}߳�\:�����|﷼�I���������~Y���  �  ��N=�8N=�M=��L=�*L=[zK==�J=�J=�eI=��H=wH=wOG=ɝF=��E=�;E=h�D=w�C=�+C=�|B=%�A=�A=�m@=�?=�?=�Y>=v�==Q�<=*=<=�;=�:=:=f_9=�8=��7=�07=u6=k�5=��4=<4=�{3==�2=��1=11=i0=P�/=��.=- .=D,-=�T,=z+=��*==�)=!�(=��'=��&=�&=�%=F$=n#=�
"=�� =��=��=p�=�z=�E=*=S�=n=-=��=�@=��=?I=�=G.=L�=n�	=�H=Q�=��=�"=0^=d'�<��<���<O&�<g�<���<���<��<��<�/�<E�<�U�<�b�<�l�<!t�<�y�<
~�<܀�<���<"��<���<���<&}�<+x�<q�<(i�<_�<fS�<8F�<8�<�(�<�<��<��y<"�q<s�i<��a<{Y<�aQ<�JI<�5A<�"9<�1<O)<�� <�<��<��<� <i��;��;Z��;���;-��;��;/0�;@��;��e;y�F;Q)(;v�	;�t�:�)�:��<:3��9O3@���$��]��s�ź^t��
F�d�6��GR��.m�ԃ�֐������R_���\»_λ��ٻ��#��=9���J�X�(D���n���K�����#��B'�k[+�[X/��93�97���:�F>���A��2E��H�s�K��O�E:R�[U��qX��[�,�^�*�a�~d��pg�@]j�{Dm��%p��s���u�3�x�zu{�_=~����������?��)���K����V������j���m��Pˌ�m)��݇��_搼�D�����������[���������g��F���}���g�����2��ka�����P	���^��ߴ��q���d����������s��Mϯ��*��?���e᳼g<������_�wK�����������Z���  �  �N=58N=ĉM=��L=+L=�zK=��J=wJ=�fI=´H=�H=�PG=K�F=�E=N=E=�D=��C=V-C=�}B=L�A=�A=dn@=��?=!?=�Y>=`�==��<=�<<=M�;=�:=�:= ^9=��8=C�7=?/7=}s6=��5=d�4=�:4=�z3=6�2=��1=e01=�h0="�/=��.=h .=�,-=�U,=�z+=��*=r�)=t�(=h�'=(�&=�	&=)%=�$=�#=$"=�� =��=q�=
�=J{=�E=
=�=~m=f=��=�?=5�=�G=_�=�,=��=��	=EG=��=5�=5!=�\=d%�<���<���<�%�<�f�<؞�<���<N��<>�<2�<uG�<mX�<�e�<�o�<jw�<}�<*��<���<u��<���<τ�<u��<�~�<Dy�<r�<Ai�<�^�<�R�<E�<R6�<�&�<��<0�<��y<��q<�i<�a<�tY<\Q<ZEI<�0A<[9<�1<��(<\� <{�<��<3�<|� <��;!��;;��;���;�ʱ;���;�=�;���;Of; 
G;VC(;��	;x��:�P�:e�<:��97�?���$�Y���źr~��QN��7��UR��@m��݃�^���&���F)��j��g»-λ�ٻ���<�ﻉ=��WL��X��C�b�@���H�ӷ�Y	#��='��U+�>R/��33���6� �:��?>���A�-E���H��K�F
O�i7R��XU��pX��[���^�҆a�`�d��sg�Iaj��Hm��*p�+s���u�J�x��{{�C~�X���Cぼ�A���������X��G������lm���ʌ�D(��X���{䐼�B��$��������X����������d��C�������d������#���_������j��1^��񴧼����e��񿫼���v���ѯ�q-�����]䳼o?������/���+N�������U\���  �  :�N=�7N=q�M=��L=F+L=B{K=��J=�J=�gI=F�H=uH=�RG=V�F=*�E=l?E=�D=�C=2/C=|B=��A=�A=bo@=T�?=�?=�Y>=>�==��<=�;<=^�;=��:=�:=v\9=��8=M�7=>-7=�q6=�5=��4=�84=7y3=�2=��1=�/1=h0=�/=��.=� .=N--=tV,=|+=�*=�)=*�(=V�'=(�&=�&=7%=�$=�#=�"=~� =2�={�=˨=�{=�E=�=��=�l=d=p�=>=f�=�E=/�==*=/�=K�	=�D=v�=-�=k=Y[=�"�<y��<:��<�$�<~f�<0��<Z��<���<X�<�4�<�J�<�[�<�i�<�s�<�{�<a��<e��<���<��<��<���<ㄭ<x��<�z�<�r�<]i�<B^�<Q�<iC�<4�<�#�<V�<��<��y<Z�q<��i<v�a<�lY<)TQ<.>I<�*A<�9<�	1<��(<�� <��<W�<��<B� <B��;y��;ע�;ݷ�;�ڱ;��;�O�;O��;$'f;�.G;�e(;��	;��:끚:�1=:͇�9��>���$�*T��#�ź����TY��7�9iR��Wm�냻�볝��7��3y��7u»H+λ��ٻv��	��+C��:N�&Y��C���ʸ�E����#�j7'��N+�EJ/�V+3�G�6���:��7>���A��%E�u�H�z�K��O��3R��VU�WoX�k[���^��a�l�d��wg��fj��Nm��1p��s���u�<�x���{��J~�����恼�D����������rY��(������7m���Ɍ� '��m���␼�?��՜��S����T��o�������`��-�������a�������	���]��(���j���]�������g����������x���ԯ�1��ጲ�j購dC����������Q��B�������^���  �  �N=�6N= �M=��L=�+L=�{K={�J=�J=siI=�H=xH=�TG=��F=��E=�AE=c�D=A�C=N1C=q�B=s�A=0!A=p@=�?=?=
Z>=�==�<=;<=1�;=i�:=�:=�Z9=��8=
�7=�*7=$o6=��5=U�4=�64=]w3=U�2=}�1=�.1=^g0=��/=��.=.=�--=lW,=Q}+=n�*=׽)=3�(=x�'=w '=�&=�%=$=�#=�"=C!=��=��=��=7|=F=�=�=�k=#=�=3<=:�=OC=��=�'=s�=��	=FB=��=��=@=�Y=��<��<��<�#�<5f�<���<c��<���<��<�7�<@N�<
`�<�m�<�x�<���<H��<2��<{��<b��<挵<䊱<���<���<�{�<�s�<si�<�]�<P�<UA�<q1�<� �<}�<E��<��y<��q<��i<|}a< cY<#KQ<�5I<#A<�9<c1<��(< � <��<��<��<�� <���;q��;w��;���;�;| �;�d�;v��;�Qf;�WG;��(;��	;H�:��:�=:+�9r>�F�$��O��A�ź�����g�h%7�3�R�Ysm�'���9���,ŝ��I��p���n�»W:λX�ٻ���j��vJ��}P�-Z�5C�"����@����t�"��/'�kF+�tA/��!3���6���:�6.>��A��E��xH�%�K�R O��/R��SU��mX�*[���^�K�a�O�d��|g��lj�MVm��9p�=s���u���x��{�T~�<����ꁼ/H������ ��D[��8���d���l���Ȍ��%��C���Sߐ�V<������ ���iP����������[������h��u]��
������![��W���?��]��)���T���h���ë����|���د�5��M����H�����������U�������ga���  �  ��N=�5N=��M=k�L=�+L=^|K=g�J=�J=kI=عH=�H=BWG=�F=�E=_DE=�D=��C=�3C=x�B=8�A=�"A=�q@=��?=�?=$Z>=ϥ==��<=/:<=�;=��:=�:=nX9=E�8=��7=\(7=�l6=&�5=��4=�44=gu3=��2=�1=�-1=�f0=&�/=��.=W.=�.-=jX,=�~+=�*=��)=X�(=��'=�'=i&=%=q$=2#=�"=!=5�=��=��=�|=/F=|=t�=�j=�=1�=+:=��=�@=�=�$=t�=��	=d?=,�=J�=�=~W=Q�<R~�<���<{"�<�e�<���<���<o��<K�<�:�<R�<dd�<�r�<�}�<���<���<N��<Y��<���<ݐ�<d��<j��<ń�<p}�<Kt�<li�<�\�<�N�<&?�<�.�<�<a�<���<a�y<�q<��i<�ra<�XY<3AQ<�,I<
A<�9<��0<��(<z� <��<9�<��<"� <~��;O��;���;���;� �;�5�;@{�;!ӂ;Of;��G;z�(;�
;�_�:���: �=:B��9�0=�#y$��L��S�ź����w�d:7��R��m���:��؝��\������w�»�Jλ�ٻ���ѹ�R���R�h[�C��
����<�6����"�('��=+��7/��3�E�6���:�$>�K�A��E�&qH�J�K���N��+R��PU�llX�6[�&�^��a�e�d�t�g�Rsj�^m�uBp�� s���u���x�)�{��]~�������K��ɧ�����&]��r�������l��Ȍ��#�����oܐ��8�������𔼕K�����������V���������7Y��Z���b���X��p���	���\��i���@��3j��ƫ��"������ܯ��9��'����MM������]��tZ��������md���  �  ��N=5N=��M=A�L=�+L=�|K=>�J=J=�lI=��H=�
H=�YG=��F=��E=�FE=o�D=�C=�5C=x�B=��A="$A=�r@=��?=�?=?Z>=��==��<=89<=��;=5�:=:=LV9=�8=�7=�%7=�i6=��5=��4=�24=os3=ݲ2=��1=l,1=�e0=��/=��.=�.==/-=\Y,=�+=��*=��)=p�(=�'=S'=�&=�%=�$=|#=�"=�!=��=�=Y�==}=PF=@=ؼ=�i=u=~�=8=��=->=�=�!=}�=��	=|<=h�=��=�=pU=��<�{�<���<M!�<Ee�<*��<���<-��<� �<>�<�U�<�h�<xw�<���<���<���<]��<4��<G��<Ԕ�<͑�<(��<φ�<�~�<�t�<ci�<\�<M�<�<�<�+�<��<-�<��<5�y<H�q<��i<�ga<�MY<17Q<�#I<�A<�9<Y�0<��(<�� <c�<��<��<a� <��;��;���;��;��;�J�;`��;�;�f;��G;��(;�?
;���:F0�:�P>:�G�9}c<�S\$��I��N�ź����߆�&P7���R���m���t#��띻�o�������»�[λ��ٻ���V��Z���U��\��B�)	���{8�â���"�U '��4+�>./��3���6�8�:�">���A�E�riH���K�b�N�y'R�/NU�kX�4[���^��a���d���g�+zj��em�PKp�Y*s��v�1�x�a�{��g~�����󁼶O�����O��#_��ɸ������l��Bǌ�d"���}���ِ�]5�����2씼�F�����������Q���������U������B ��*V���������;\������9���k��eȫ��%��(����௼,>�����*���lR��Ȭ��B��_��H���T���g���  �  ��N=64N=n�M=�L=,L=X}K=�J=<J=�mI=Y�H=�H=�[G=��F=��E=TIE=��D=M�C=�7C=V�B=��A=t%A=�s@=y�?=[?=JZ>=F�==F�<=J8<=p�;=��:=M:=AT9=ș8=��7=h#7=�g6==�5=N�4=o04=�q3=9�2=I�1=Z+1=e0=L�/=��.=�.=�/-=EZ,=�+=#�*=U�)=`�(=3�'=�'=5&=�%=!$=�#=�"=�!=�=%�=%�=�}=eF=�=4�=�h=&=ޥ=66=m�=�;=��=	=��=��	=�9=ۉ=F�=w=�S=��< y�<���< �<�d�<f��<x��<���<#�<�@�<IY�<�l�<�{�<D��<���<���<��<���<\��<���<���<���<ƈ�<��<�u�<*i�<-[�<�K�<�:�<�(�<�<!�<|��<Ƽy<@�q<�zi<�]a< DY<�-Q<�I<LA<a�8<�0<�(<	� <�<��<�<�� <5��;]��; ��;V��;j&�;O^�;ҥ�;���;��f;~�G;s);�b
;*��:ke�:{�>:mЎ9�;�RE$��I��f�ź�������Zd7�
�R���m��+���4������⁪�����A�»xkλ9�ٻ���o���a��dX�^�#C�������4������"��'��,+��%/�x3�i�6��x:��>��A��E�bH���K�f�N��#R��KU��iX��[�'�^�ԓa���d�D�g���j�Rmm��Sp� 3s�ev���x���{�Dq~�����:���aS��&������a�����,���l���ƌ�!���{�� א�<2��V���(蔼iB����������L��8�������4Q��7���q����S����������[�����?���m���ʫ�u(�������䯼gB����������3W�������
��Oc��I������gj���  �  ��N=�3N=��M=��L=,L=�}K=��J=J=oI=��H='H=n]G=��F=��E=NKE=ǚD=6�C=�9C=�B=��A=�&A=�t@=�?=�?=RZ>=�==��<=�7<=W;=h�:=�:=�R9=ؗ8=��7=R!7=|e6=/�5=L�4=�.4=�o3=ί2=�1=g*1=yd0=�/=��.=	.=80-=�Z,=�+=e�*=��)=
�(=�'=�	'='&=�%=�"$=S #=}"=�!=N�=
�=¬=�}=lF=�=��=h= =r�=�4=��=�9=D�=�=K�=l�	=e7=��=9�=�=�Q=��<�v�<��<��<Jd�<z��<>��<* �< %�<uC�<B\�<p�<��<T��<Ɠ�<���<��<_��<ٝ�<���<���<Ǒ�<P��<���<�u�<�h�<hZ�<CJ�<�8�<2&�<
�<���<��<C�y<��q<�qi<�Ta<];Y<�%Q<�I<�A<��8<J�0< �(<�� <��<��<P�<� <l��;=��;���;@
�;�5�;-o�;z��;��;��f;#�G;8&);��
;o�:c��:��>:[?�93;��2$�4J��+�ź�������v7���R���m�:���C�����ؑ��dѶ�s�»7yλ��ٻ���U���h���Z�h_�?C������t1����y�"��'��%+�!/�l�2�[�6��p:��>���A��D�\H�I�K�M�N�� R��IU�iX��[���^�3�a�`�d��g��j��sm��Zp�;s��v�2�x�V�{�my~�圀������V��а��
���b��$�������l��ƌ����7z���Ԑ��/��8����䔼�>���������H��O���N����M��f��� ���R������0���[��`��� ���n���̫��*������	诼%F������ ��p[���������g����������l���  �  ��N=�2N=��M=��L=,,L=�}K=1�J=�J=pI=̿H=bH=�^G=�F={�E=�LE=A�D=��C=�:C=�B=��A=r'A=Iu@=��?=�?=XZ>=ͤ==M�<=�6<=}~;=]�:=�:=7Q9=_�8==�7=�7=�c6=��5=��4=;-4=�n3=��2=&�1=�)1=�c0=��/=o�.=".=�0-=�[,=т+=]�*=��)=P�(=a�'=�
'=�&=>!%=`$$=�!#=�"=�!=9�=��=;�=G~=lF=�=2�=gg=
=X�=>3=�=8=��=�=r�=��	=�5=م=��==�P=��<u�<���<$�<�c�<���<���<,�<�&�<aE�<x^�<�r�<I��<D��<ٖ�<���<��<<��<���<ѝ�<���<S��<|��<���<7v�<�h�<�Y�<I�<7�<9$�<��<��<��<�y<
�q<�ji<Na<�4Y<�Q<�I<v�@<L�8<��0<B�(<�� <�<��<b�<� <���;���;���;��;�A�;�{�;�Ē;�;vg;�H;�>);Җ
;�>�:$��:�'?:9�:��$$��J��]�ź������g�7�B�R���m��D��O��t������ܶ���»��λ�ٻ�S��Sn���\�w`�QC�c���/�i��i�"��'�� +�w/���2�/�6��j:�>��A���D��WH�?�K��N�@R�,HU��hX��[���^�a�a�@�d���g���j��xm�B`p�*As��v���x���{�r~�㟀�]����X��񲄼���d�����<���l���Ō����x��!Ӑ��-��臓��ᔼ�;������혼�E��w�������bK��C�������P����������[���������#p��AΫ��,��ً���꯼�H������%���^��ϸ������i��=���-���n���  �  E�N=�2N=S�M=��L=-,L="~K=y�J== J=�pI=z�H='H=�_G=�F=t�E=�ME=4�D=��C=�;C=ފB=��A=�'A=�u@=��?=�?=OZ>=��==
�<=s6<=�};=��:=�
:=PP9=s�8=;�7=�7=�b6=��5=��4=O,4=�m3=��2=��1=<)1=�c0=f�/=V�.=1.=�0-=�[,=G�+=�*=��)=�(=@�'=�'=�&=9"%=M%$=�"#=|"=�	!=��=)�=��=d~=mF=[=�=�f=�	=��=r2=%�=7=t�=�=E=f�	=z4=ʄ=��=9=�O=j�<�s�<���<��<�c�<���<*��<��<i'�<�F�<�_�<>t�<��<,��<��<���<���<
��<��<M��<���<P��<(��<(��<Rv�<�h�<UY�<^H�<;6�<�"�<5�<K��<��<�y<��q<Zfi<�Ia<�0Y<�Q<-
I<W�@<��8<��0<��(<�� <g�<��<��</� <���;Z��;���;t�;+I�;���;;͒;'�;r%g;i$H;N);��
;�V�:ɛ:�I?:Ï9�r:��$��K����ź��������7�
 S�Qn��K���V��x ��ᥪ�	嶻0�»��λF�ٻT廯��iq���]�a��C�����-�t��#�"��'�r+��/���2�)�6��f:�'�=�N�A���D��TH���K�,�N��R�kGU�4hX�3�[�e�^���a��d�ԗg�:�j��{m��cp��Ds��v���x��{���~�����/����Z��?�������d����������l��oŌ����4x��$Ґ�H,��f���Z����9��"����똼�C���������I��ܠ������O�����6��u[��ض��L���p��!ϫ�.��@���J쯼�J������D���`�������k���º����)p���  �  �N=W2N=A�M=��L=3,L=0~K=��J=l J=�pI=��H=dH=�_G=a�F=��E="NE=~�D=��C=<C= �B=��A=(A=�u@=��?=?=SZ>=��==��<=H6<=�};=z�:=�
:=P9=+�8=��7=^7=�b6=@�5=��4= ,4=�m3=ǭ2=X�1=)1=oc0=P�/=K�.=E.=�0-=�[,=u�+=�*=��)=N�(=��'=+'=�&=~"%=�%$=�"#=�"=�	!=��=Q�=��=s~=F=L=Ժ=�f=`	=i�=22=ڸ=�6=#�=X=�~=�	=4={�=D�=�=�O=��<�s�<���<��<�c�<Ϡ�<L��<&�<�'�<�F�<z`�<�t�<���<Đ�<��<G��<���<���<���<џ�<��<���<]��<H��<av�<�h�<(Y�<H�<�5�<t"�<��<���<�<��y<�q<1ei<*Ha<\/Y<TQ< 	I<m�@<��8<��0<��(<l� <I�<��<E�<�� <Q��;���;���;��;�K�;���;�ϒ;�)�;�*g;*H;�R);��
;_�:�ϛ:�V?:1Ϗ9�Z:��$��L��@�ź���ع�G�7��S��
n�N��[Y���"�������綻r�»,�λ[�ٻ��n���r��[^�]a��C���Ǩ� -����g�"�o
'��+��/�m�2��6�be:���=�#�A���D��SH�4�K�x�N�JR�GU��gX�P�[���^��a���d���g��j��|m�.ep��Es�B v���x��{��~�C��������Z������K��9e��Ἀ�����l��@Ō�o���w���ѐ��+��م���ߔ�\9������,똼SC��蚛�B�bI��Y�������UO��ʧ����a[����s��-q���ϫ��.�������쯼nK��*������Da���������gl���ú�	���p���  �  E�N=�2N=S�M=��L=-,L="~K=y�J== J=�pI=z�H='H=�_G=�F=t�E=�ME=4�D=��C=�;C=ފB=��A=�'A=�u@=��?=�?=OZ>=��==
�<=s6<=�};=��:=�
:=PP9=s�8=;�7=�7=�b6=��5=��4=O,4=�m3=��2=��1=<)1=�c0=f�/=V�.=1.=�0-=�[,=G�+=�*=��)=�(=@�'=�'=�&=9"%=M%$=�"#=|"=�	!=��=*�=��=e~=oF=]=�=g=�	=��=v2=*�=7=z�=�=N=o�	=�4=Մ=��=E=�O=��<t�<��<��<�c�<���<B��<��<}'�<�F�<�_�<Jt�<(��<1��<��<���<��<��<��<>��<���<=��<��<��<;v�<�h�<>Y�<HH�<&6�<�"�<%�<>��<��<کy<��q<Zfi<�Ia<�0Y<�Q<G
I<w�@<��8<��0<��(<�� <��<�<)�<Z� <���;���;���;��;QI�;ڃ�;E͒;'�;K%g;#$H;�M);}�
;�U�:�Ǜ:�F?:���9r�:��#$��M��m�źk	��w��r�7�� S�%n�3L��W��� ��/���P嶻p�»�λx�ٻ����ﻊq���]�a��C��%���-�y��'�"��'�u+��/���2�*�6��f:�'�=�O�A���D��TH���K�,�N��R�kGU�4hX�3�[�e�^���a��d�ԗg�:�j��{m��cp��Ds��v���x��{���~�����/����Z��?�������d����������l��oŌ����4x��$Ґ�H,��f���Z����9��"����똼�C���������I��ܠ������O�����6��u[��ض��L���p��!ϫ�.��@���J쯼�J������D���`�������k���º����)p���  �  ��N=�2N=��M=��L=,,L=�}K=1�J=�J=pI=̿H=bH=�^G=�F={�E=�LE=A�D=��C=�:C=�B=��A=r'A=Iu@=��?=�?=XZ>=ͤ==M�<=�6<=}~;=]�:=�:=7Q9=_�8==�7=�7=�c6=��5=��4=;-4=�n3=��2=&�1=�)1=�c0=��/=o�.=".=�0-=�[,=т+=]�*=��)=P�(=a�'=�
'=�&=?!%=`$$=�!#=�"=�!=:�=��==�=I~=nF=�=6�=kg= 
=_�=G3=�=8=��=�=��=��	=�5=�=��=6=�P=��<9u�<���<Y�<.d�< �<��<X�<�&�<�E�<�^�<�r�<Y��<M��<ܖ�<���<���<+��<h��<���<o��<-��<S��<���<v�<�h�<�Y�<�H�<�6�<$�<��<���<��<ѭy<��q<�ji<&Na<�4Y<�Q<I<��@<��8<��0<��(<� <^�<D�<��<[� <���;���;W��;7�;�A�;�{�;�Ē;��;)g;H;>);��
;J<�:���:�!?:I��9��:��+$�`N���ź������%�7���R���m��E���O��������wݶ�x�»�λu�ٻo廝�ﻒn���\��`�eC�t����#/�r��q�"��'�� +�|/���2�1�6��j:�>��A���D��WH�@�K��N�AR�,HU��hX��[���^�a�a�@�d���g���j��xm�B`p�*As��v���x���{�r~�㟀�]����X��񲄼���d�����<���l���Ō����x��!Ӑ��-��臓��ᔼ�;������혼�E��w�������bK��C�������P����������[���������#p��AΫ��,��ً���꯼�H������%���^��ϸ������i��=���-���n���  �  ��N=�3N=��M=��L=,L=�}K=��J=J=oI=��H='H=n]G=��F=��E=NKE=ǚD=6�C=�9C=�B=��A=�&A=�t@=�?=�?=RZ>=�==��<=�7<=W;=h�:=�:=�R9=ؗ8=��7=R!7=|e6=/�5=L�4=�.4=�o3=ί2=�1=g*1=yd0=�/=��.=	.=80-=�Z,=�+=e�*=��)=
�(=�'=�	'=(&=�%=�"$=T #=}"=�!=O�=�=Ĭ= ~=pF=�=��=$h=	=|�=�4=��=�9=V�=�=b�=��	=�7=��=Y�=�=R=*�<w�<S��<<�<�d�<���<���<h �<8%�<�C�<k\�</p�<��<a��<ɓ�<���<��<F��<���<`��<W��<���<��<���<�u�<�h�<+Z�<J�<w8�< &�<��<���<�<�y<��q<�qi<�Ta<�;Y<�%Q<�I< A<!�8<��0<��(<9� <]�<R�<��<�� <J��;��;���;�
�;`6�;po�;���;��;y�f;f�G;,%);.
;:�:���:��>:z-�9:E;�r<$�MO��S�ź
���A��}x7�[�R���m�;���D��q������&Ҷ�!�»�yλ/�ٻ 廽��(i���Z��_�[C������1������"�'��%+�'/�q�2�_�6��p:��>���A��D�\H�J�K�N�N�� R��IU�iX��[���^�3�a�`�d��g��j��sm��Zp�;s��v�2�x�V�{�my~�圀������V��а��
���b��$�������l��ƌ����7z���Ԑ��/��8����䔼�>���������H��O���N����M��f��� ���R������0���[��`��� ���n���̫��*������	诼%F������ ��p[���������g����������l���  �  ��N=64N=n�M=�L=,L=X}K=�J=<J=�mI=Y�H=�H=�[G=��F=��E=TIE=��D=M�C=�7C=V�B=��A=t%A=�s@=y�?=[?=JZ>=F�==F�<=J8<=p�;=��:=M:=AT9=ș8=��7=h#7=�g6==�5=N�4=o04=�q3=9�2=I�1=Z+1=e0=L�/=��.=�.=�/-=EZ,=�+=#�*=U�)=`�(=3�'=�'=6&=�%=!$=�#=�"=�!=�=(�=(�=�}=jF=�=;�=�h=0=�=D6=~�=�;=��="=Մ=��	=�9= �=m�=�=�S=�<\y�< ��<g �<e�<���<���<)��<Z#�<9A�<{Y�<�l�<�{�<T��<ď�<x��<��<v��<3��<R��<���<z��<��<��<;u�<�h�<�Z�<@K�<f:�<p(�<��<��<Z��<��y<(�q<�zi<�]a<NDY<6.Q<AI<�A<��8<��0<�(<�� <��<\�<��<� <E��;P��;���;��;�&�;�^�;���;���;#�f;��G;+);a
;<��:�`�:g�>:���9��;�zQ$��O����ź,������`g7���R���m�-���5��
���肪��¶��»6lλ��ٻ������Lb���X�B^�EC��í��4�Ɲ���"�	'��,+��%/�~3�n�6��x:��>��A��E�bH���K�g�N��#R��KU��iX��[�'�^�ԓa���d�D�g���j�Rmm��Sp� 3s�ev���x���{�Dq~�����:���aS��&������a�����,���l���ƌ�!���{�� א�<2��V���(蔼iB����������L��8�������4Q��7���q����S����������[�����?���m���ʫ�u(�������䯼gB����������3W�������
��Oc��I������gj���  �  ��N=5N=��M=A�L=�+L=�|K=>�J=J=�lI=��H=�
H=�YG=��F=��E=�FE=o�D=�C=�5C=x�B=��A="$A=�r@=��?=�?=?Z>=��==��<=89<=��;=5�:=:=LV9=�8=�7=�%7=�i6=��5=��4=�24=os3=ݲ2=��1=l,1=�e0=��/=��.=�.==/-=\Y,=�+=��*=��)=p�(=�'=T'=�&=�%=�$=|#=�"=�!=��=�=\�=A}=UF=F=�=�i=�=��=.8=��=B>=5�=�!=��=��	=�<=��=��=�=�U=T�<|�<���<�!�<�e�<���<���<���<!�<\>�<�U�<�h�<�w�<���<���<���<H��<��<��<���<���<ߌ�<���<~�<�t�<i�<�[�<�L�<�<�<=+�<E�<��<��<�y<.�q<��i<�ga<(NY<}7Q<$I<vA<i9<��0<,�(<d� <�<E�</�<� <>��;���;���;���;�;9K�;���;��;��f;��G;t�(;�=
;���:;+�:�E>:/�9o�<��i$��P��Y�ź����U���S7��R���m�����$��T읻#q�������»�\λy�ٻa����ﻋZ��V��\�C�I	�1���8�֢���"�b '��4+�F./��3���6�=�:�&>���A�E�tiH���K�c�N�z'R�0NU�kX�5[���^��a���d���g�+zj��em�PKp�Y*s��v�1�x�a�{��g~�����󁼶O�����O��#_��ɸ������l��Bǌ�d"���}���ِ�]5�����2씼�F�����������Q���������U������B ��*V���������;\������9���k��eȫ��%��(����௼,>�����*���lR��Ȭ��B��_��H���T���g���  �  ��N=�5N=��M=k�L=�+L=^|K=g�J=�J=kI=عH=�H=BWG=�F=�E=_DE=�D=��C=�3C=x�B=8�A=�"A=�q@=��?=�?=$Z>=ϥ==��<=/:<=�;=��:=�:=nX9=E�8=��7=\(7=�l6=&�5=��4=�44=gu3=��2=�1=�-1=�f0=&�/=��.=W.=�.-=jX,=�~+=�*=��)=X�(=��'=�'=i&=%=q$=3#=�"=!=7�=��=��=�|=4F=�=|�=�j=�=?�=<:=�=�@=��=�$=��=��	=�?=V�=w�=&=�W=��<�~�<���<�"�<"f�<D��<���<���<��<+;�<=R�<�d�<�r�<�}�<���<|��<8��<6��<���<���<!��<��<s��<}�<�s�<i�<�\�<[N�<�>�<:.�<��<-�<s��<+�y<�q<��i<�ra<�XY<�AQ<9-I<�A<l9<��0<��(<,� <E�<��<b�<�� <���;h��;���;t��;j�;6�;g{�;ӂ;�~f;��G;��(;�
;C[�:p�:\�=:���9�f=�,�$��S����źʸ���z��=7�>�R�K�m�������[ٝ�^�����m�»�Kλķٻk��d�ﻞR��0S��[�=C��
�����<�I����"�('��=+��7/��3�K�6���:�$>�N�A��E�(qH�L�K���N��+R��PU�llX�7[�&�^��a�e�d�t�g�Rsj�^m�vBp�� s���u���x�)�{��]~�������K��ɧ�����&]��r�������l��Ȍ��#�����oܐ��8�������𔼕K�����������V���������7Y��Z���b���X��p���	���\��i���@��3j��ƫ��"������ܯ��9��'����MM������]��tZ��������md���  �  �N=�6N= �M=��L=�+L=�{K={�J=�J=siI=�H=xH=�TG=��F=��E=�AE=c�D=A�C=N1C=q�B=s�A=0!A=p@=�?=?=
Z>=�==�<=;<=1�;=i�:=�:=�Z9=��8=
�7=�*7=$o6=��5=U�4=�64=]w3=U�2=}�1=�.1=^g0=��/=��.=.=�--=lW,=Q}+=n�*=׽)=3�(=x�'=w '=�&=�%=$=�#=�"=D!=��=��=��=;|=F=�=�=�k=.=�=C<=M�=dC=ù=�'=��=��	=kB=�=��=n=�Y= �<Y��<���<$�<�f�<���<���<���<�<�7�<xN�<6`�<n�<�x�<���<@��<��<Y��<4��<���<���<Q��<D��<�{�<Fs�<i�<F]�<�O�<	A�<,1�<y �<L�<��<O�y<w�q<��i<�}a<3cY<oKQ<,6I<�#A<F9<�1<��(<�� <t�<��<g�<:� <��;���;a��;���;��;� �;e�;d��;0Qf;�VG;'�(;��	;��:��:Є=:��9g9>�գ$��V��L�ź����)k��(7�q�R�nvm������ ��lƝ��J��x���\�»*;λ�ٻ�������J���P�ZZ�[C�B����@�ҭ���"��/'�uF+�|A/��!3���6���:�:.>��A��E��xH�&�K�S O��/R��SU��mX�*[���^�K�a�O�d��|g��lj�MVm��9p�=s���u���x��{�T~�<����ꁼ/H������ ��D[��8���d���l���Ȍ��%��C���Sߐ�V<������ ���iP����������[������h��u]��
������![��W���?��]��)���T���h���ë����|���د�5��M����H�����������U�������ga���  �  :�N=�7N=q�M=��L=F+L=B{K=��J=�J=�gI=F�H=uH=�RG=V�F=*�E=l?E=�D=�C=2/C=|B=��A=�A=bo@=T�?=�?=�Y>=>�==��<=�;<=^�;=��:=�:=v\9=��8=M�7=>-7=�q6=�5=��4=�84=7y3=�2=��1=�/1=h0=�/=��.=� .=N--=tV,=|+=�*=�)=+�(=W�'=(�&=�&=7%=�$=�#=�"=� =3�=}�=Ψ=�{=�E=�=��=�l=n=|�=>=w�=�E=E�=V*=K�=j�	=E=��=U�=�=�[=&#�<Ճ�<���<&%�<�f�<���<���<)��<��<�4�<�J�<!\�<�i�<�s�<�{�<Y��<R��<ڇ�<눹<܈�<i��<���<1��<8z�<~r�<i�<�]�<7Q�<%C�<�3�<�#�<*�<^�<��y<B�q<��i<��a<�lY<mTQ<�>I<�*A<u9<
1<Q�(<� <Q�<��<l�<�� <Q��;m��;���;���;>۱;��;P�;?��;�&f;�-G;Vd(;B�	;+��:e}�:�'=:�q�9�
?���$�hZ��s�źB���n\��7�!lR��Zm�Y샻�
���9�� z��v»,λ2�ٻ	�仉�ﻚC��iN�OY��C�����E�'���#�u7'��N+�LJ/�\+3�L�6���:��7>���A��%E�v�H�{�K��O��3R��VU�XoX�l[���^��a�l�d��wg��fj��Nm��1p��s���u�<�x���{��J~�����恼�D����������rY��(������7m���Ɍ� '��m���␼�?��՜��S����T��o�������`��-�������a�������	���]��(���j���]�������g����������x���ԯ�1��ጲ�j購dC����������Q��B�������^���  �  �N=58N=ĉM=��L=+L=�zK=��J=wJ=�fI=´H=�H=�PG=K�F=�E=N=E=�D=��C=V-C=�}B=L�A=�A=dn@=��?=!?=�Y>=`�==��<=�<<=M�;=�:=�:= ^9=��8=C�7=?/7=}s6=��5=d�4=�:4=�z3=6�2=��1=e01=�h0="�/=��.=h .=�,-=�U,=�z+=��*=r�)=t�(=h�'=(�&=�	&=)%=�$=�#=%"=�� =��=s�=�=M{=�E==�=�m=n=ŭ=�?=C�=�G=q�=�,=��=��	=`G=Ö=U�=W!=]=�%�<υ�<���<�%�<g�<��<���<���<v�<62�<�G�<�X�<�e�<�o�<nw�<}�<��<׃�<T��<���<���<@��<s~�<y�<�q�<i�<k^�<TR�<�D�< 6�<�&�<t�<�<��y<��q< �i<+�a<%uY<?\Q<�EI<!1A<�9<-1<R�(<�� <��<b�<��<�� <�;��;��;*��;�ʱ;@��;�=�;���;�f;B	G;JB(;3�	;B��:M�:*�<:���9@�?�m�$�+^��>�ź�����P�+7�LXR��Bm�
߃�[ᐻ���*���j���g»�λ��ٻ�令���=��~L��X�	D�y�S���H���d	#��='��U+�DR/��33���6�$�:� @>���A�-E���H��K�F
O�i7R��XU��pX��[���^�҆a�`�d��sg�Iaj��Hm��*p�+s���u�J�x��{{�C~�X���Cぼ�A���������X��G������lm���ʌ�D(��X���{䐼�B��$��������X����������d��C�������d������#���_������j��1^��񴧼����e��񿫼���v���ѯ�q-�����]䳼o?������/���+N�������U\���  �  ��N=�8N=�M=��L=�*L=[zK==�J=�J=�eI=��H=wH=wOG=ɝF=��E=�;E=h�D=w�C=�+C=�|B=%�A=�A=�m@=�?=�?=�Y>=v�==Q�<=*=<=�;=�:=:=f_9=�8=��7=�07=u6=k�5=��4=<4=�{3==�2=��1=11=i0=P�/=��.=- .=D,-=�T,=z+=��*==�)=!�(=��'=��&=�&=�%=F$=o#=�
"=�� =��=��=q�=�z=�E=-=W�=n=3=Ů=�@=��=JI=�=U.=\�=��	=I=f�=��=�"=I^=�'�<N��<��<�&�<@g�<���<���<?��<��<0�<6E�<�U�<�b�<�l�<$t�<�y�<�}�<ʀ�<���<��<j��<j��<�|�<�w�<Sq�<�h�<�^�<<S�<F�<�7�<�(�<��<��<|�y<�q<s�i<��a<9{Y<bQ<�JI<�5A<�"9<<1<�)<D� <u�<��<�<k� <��;���;ӌ�;��;w��;#�;B0�;6��;Q�e;��F;�((;��	;�r�:_'�:�<:���94N@���$�1a���źx���G�"�6�6IR�\0m��ԃ��֐���������_��?]»�λ��ٻk��m��}9���J�-X�;D���|���K�����#��B'�p[+�_X/��93�<7���:�F>���A��2E��H�t�K��O�F:R�[U��qX��[�,�^�*�a�~d��pg�@]j�{Dm��%p��s���u�3�x�zu{�_=~����������?��)���K����V������j���m��Pˌ�m)��݇��_搼�D�����������[���������g��F���}���g�����2��ka�����P	���^��ߴ��q���d����������s��Mϯ��*��?���e᳼g<������_�wK�����������Z���  �  2�N=�8N=2�M=��L=�*L=zK=��J=,J=eI=زH=� H=�NG=ϜF=x�E=�:E=Y�D=��C=+C=�{B=r�A=�A=.m@=��?=�?=�Y>=�==|�<=y=<=y�;=��:=�:=+`9=Ȧ8=��7=�17=v6=^�5=��4=�<4=�|3=ֺ2=,�1=c11=<i0=n�/=��.= .=�+-=�T,=�y+=�*={�)=:�(=�'=��&=�&=�%=A$=�#=�	"=� =M�=&�=�=�z=}E=0=��=fn=�=^�=�A=t�=9J=�=n/=��=��	=$J=l�=��=�#=�^=�(�<1��<���<�&�<;g�<���<U��<���<��<�.�<�C�<T�<�`�<�j�<r�<�w�<�{�<�~�<���<x��<��<]�<(|�<nw�< q�<�h�<_�<�S�<�F�<�8�<
*�<��<�
�<j�y<�q<Ƿi<��a<DY<�eQ<TNI<�8A<%9<51<�)<
� <��<v�<,�<�� <��;5��;���;���;���;��;'�;<}�;��e;��F;�(; �	;GX�:�:\s<:V�9��@���$�fc����źq���A���6��>R�%m�Z΃��ϐ�C�������X��9V»�λE�ٻ��ǔﻰ6��AJ��W��D�J����KM�����#�!F'�(_+�\/��=3�u7�ͳ:�TJ>���A�A6E��H�#�K�O��;R�N\U��rX��[�Ʌ^�h�a��|d��ng��Zj�Am�p"p���r�&�u�)�x��q{��9~��~�� ߁�>�����]���IV��2���O���m���ˌ�*�������琼)F��I�������]���������i��D���S��Zi������|��cb��Ƶ���	���^��촧�)��{d��ҽ������r���ͯ�)��a���}߳�\:�����|﷼�I���������~Y���  �  �N=�0N=$�M=��L=$ L=�nK=�J=�
J=aXI=��H=��G=3@G=��F=Q�E=_)E=swD=��C=�C=/cB=��A=��@=�M@=�?=��>=N3>=+~==��<=�<=�X;=��:=��9=�*9=7o8=��7=�6=�66=�v5=H�4=6�3=�03=]k2=0�1=��0=0=�@/=po.=+�-=��,=��+=]
+=>(*=iB)=�X(=�j'=�x&=�%=��$=4�#=p�"=�t!=�b =J=Z*=�=��=�=�[=�=��= f=	=�=o= �=3=2�=P�
=�U	=��==�O=��=c� =��<���<���<:�<���<R��<���<�1�<�\�<���<��<��<���<3��<'��<K�<~�<�<%�<�,�<p2�<�6�<�9�<;�<�:�<�8�<%5�<0�<�)�<_"�<"�<\�<$�<��y<��q<��i<{�a<�Y<[�Q<��I<��A<}�9<��1<A�)<�!<��<�<%�	<��<�L�;k�;6��;���;��;�^�;�Ô;�=�;!�k;�L;{].;n;D��:��:8xY:�Z�9 �����s�w�B������E0�I�-�۩H�tRc�ۏ}�4����Y���Ǥ����e弻G�ȻF�ӻ�$߻�	����D��p���	�`\�d����i��{ �»$���(��,��0�A�4��n8�<�#�?��'C��F���I��;M��zP���S���V�n�Y�(
]�o`�5c�>f��i�l���n�1�q�K�t� �w��wz�K}����r��ׂ�H:��Y�������	_��￉�!������ ㍼D���������e���Ĕ�#��]����ۘ��6��L����蜼$@��������D��㚣�"�J��ˢ��_����V���������.j���Ư��#������`ݳ��9��������SO������{���e���  �  ��N=�0N=�M=��L=0 L=�nK=/�J=J=�XI=�H=%�G=q@G=�F=��E=})E=�wD=4�C=�C=icB=�A=$ A=�M@=*�?=��>=X3>=~==��<=�<=�X;=��:=��9=�*9=o8=`�7=��6=Z66=�v5=�4=�3=u03=3k2=�1=��0=�0=�@/=uo.=8�-=��,=��+=}
+=k(*=�B)=�X(=k'=�x&=>�%=�$={�#=��"=�t!=�b =EJ=y*==��=�=�[=�=��=�e=�=�='=Ġ=�=�=�
=�U	=��=�=MO=O�=5� =��<\��<���<�9�<���<Y��<���<�1�<�\�<��<���<b��<T��<���<j��<��<�<��<�%�<�,�<�2�<E7�<:�<G;�<�:�<�8�<5�<�/�<�)�<("�<��<��<��<�y<��q<��i<��a<)�Y<k�Q<��I<��A<�9<ݎ1<ɋ)<v�!<J�<�<Z�	<>�<rM�;il�;���;���;��;a�;�Ŕ;�>�;��k;��L;#b.;�;���:��:��Y:hp�9�Ј������w� ������[1�]�-���H��Tc���}����� [��Qɤ�n����漻��Ȼ�ӻ�%߻�
�ӭ���������	�!\� �����{ ��$�|�(��,���0���4�2n8��<�9�?��&C��F���I�>;M�RzP�I�S���V�M�Y�{
]��`��c��f��i��l�_�n���q��t�ޠw��xz��K}����Cs���ׂ��:���������3_������ ��ہ���⍼�C������D��2e��mĔ��"������ۘ�]6������蜼�?������@��C���������I��Т�������V��?������j��9ǯ�$�������ݳ�q:������^󷼼O��,�������e���  �  ��N=�0N=�M=��L=B L=oK={�J=iJ=
YI=n�H=��G=AG=��F=X�E=G*E=�xD=��C=pC=dB=n�A=� A=MN@=p�?=��>=h3>=~==��<=�<=JX;=0�:=�9=,*9=Xn8=��7=�6=�56=v5=a�4=h�3=�/3=�j2=��1=g�0=�0=�@/=}o.=L�-=��,=/�+=�
+=�(*=&C)=yY(=�k'=�y&=�%=��$=A�#=E�"=�u!=~c =�J=�*=Y=��=�=�[=�=��=ve=`=\�={=�=#=�=(�
=�T	=׮==�N=��=�� =t�<���<��<s9�<h��<^��<4 �<^2�<�]�<ւ�<���<���<���<]��<��<^�<��<��<�&�<%.�<�3�<%8�<�:�<�;�<;�<�8�<�4�<�/�<�(�<d!�<��<��<r�<�y<��q<j�i<��a<!�Y<��Q<�I<Z�A<��9<-�1<��)<ɉ!<��<4�<ۓ	<T�<KP�;Vp�;��;��;{�;Eg�;�̔;�E�;R�k;S�L;yn.;Q;|��:�.�:��Y:ƣ�9�Q�������w�头���캶5�f�-���H��\c�ԛ}�����b`���Τ������뼻�ȻԻ�(߻i������������	��[��¤�#��x ���$���(�z�,���0�W�4��j8��<���?�9$C�ՐF���I��9M�yP�_�S�2�V�(�Y��
]�<`�� c�V!f�Ii�6l���n���q���t��w��{z��N}����qt���؂�Z;��_�������j_��2���� ������a⍼5C��֣��<��d��Ô�F!��/~��ژ��4��@����朼c>������@젼C��������I��Т������ZW��������k��Xȯ�S%��W���4߳��;��g�������Q��O����	���f���  �  �N=-0N=M=��L=c L=ioK=�J=J=�YI=N�H=��G=6BG=��F=~�E=w+E=�yD=�C=�C=�dB=I�A=QA=�N@=ۛ?=�>=�3>=~==��<=!<=�W;=x�:=D�9=6)9=Lm8=��7= �6={46=�t5=N�4=b�3=/3=�i2=	�1=��0=0=h@/=~o.=|�-=P�,=��+=�+=�)*=D)=|Z(=�l'=�z&=,�%=Ј$=P�#=\�"=�v!=Zd =�K=p+=�=3�=;�=�[=i=)�=�d=� =n�=s=ٞ=�=ш=��
=VS	=��=� =bM=��=�� =��<_��<7��<�8�<<��<���<� �<=3�<�^�<d��<e��<���<���<���<i��<�	�<��<Y �<)�<0�<�5�<�9�<�;�<�<�<�;�<�8�<�4�</�<(�< �<C�<��<Q�<��y<*�q<��i<��a<r�Y<�Q<�I<ϔA<ˎ9<��1<҈)<��!<��<}�<ݔ	<�<U�;`v�;a��;a��;��;�p�;�֔;ZP�;��k;�M;�.;�.;��:bK�:G�Y:���9Ym��[��]�w�G�������;���-�L�H�>jc���}�j����h���֤�����󼻭�Ȼ�Ի�.߻��<������I��m�	��Z�v����l��u ���$���(���,�D�0���4�4f8�J<��?� C�#�F�]�I��6M��vP�ЪS�T�V��Y�:]��`��"c��#f�Vi��l�� o��q�L�t�M�w��z�
S}����fv��Aڂ��<������n����_��W���� ��&����፼B��u������!b���������{���ט�o2��	����䜼d<�������꠼�A��!����𤼌I��ע�����X��峫�@��m��*ʯ�d'��~���q᳼/>����������S��+���p��h���  �  o�N=�/N=z�M=��L=� L=�oK=|�J=�J=�ZI=u�H=��G=�CG=@�F=
�E=-E=/{D=��C=�C=3fB=e�A=7A=�O@=^�?=j�>=�3>=�}==7�<=�<=W;=��:=1�9=�'9=�k8=!�7=u�6=�26=ws5=�4=�3=�-3=�h2=5�1=W�0=0=3@/=xo.=��-=��,=J�+=U+=�**=9E)=�[(=,n'=5|&=��%=V�$=̉#=Ń"=�w!=}e =sL=*,=S=��=]�=�[==��=d=��=8�==V�=E=�=�
=�Q	=ѫ=+�=�K=>�=|� =��<Ѓ�<��<@8�<���<���<h�<a4�<o`�<_��<���<B��<���<���<���<��<�<L#�<�+�<�2�<�7�<J;�<2=�<|=�<<�<�8�<F4�<'.�<�&�<S�<0�<��<��<��y<��q<=�i<*�a<>�Y<F�Q<��I<�A<��9<��1<X�)<!�!<�<َ<&�	<!�<([�;~�;���;���;�(�;	~�;v�;1^�;!�k;#M;`�.;�E;�H�:�o�:qZ:�P�9;H����@�w�>���U��oD��-���H��{c�ɽ}�ǋ��s��P⤻	�����=�Ȼ�Ի6߻�껂���������J�	��Y������	�pq ��$�h�(���,��0�C�4��_8�<�"�?��C�?�F�8�I��3M�ItP��S�A�V���Y��]�(`��$c��&f�R"i�!l��o�v�q�R�t�w�w�E�z��X}�����x��r܂��>������� ���`������� �����������@������\ ���_��R������x���Ԙ�T/�������᜼�9��b����蠼:@������2�+I����������Y��3�����$o���̯�*��R���|䳼:A�����������U����������i���  �  ��N=/N=#�M=��L=� L=.pK=&�J=�J=�[I=��H=~�G=0EG=�F=��E=�.E=�|D=.�C=rC=�gB=��A=CA=pP@=��?=��>=�3>=�}==��<=�<=#V;=u�:=��9=}&9=]j8=o�7=��6=816=�q5=F�4=��3=~,3=�g2=;�1=��0=�0=�?/=so.=��-=.�,=�+=J+=�+*=�F)=?](=�o'=�}&=p�%=�$=�#=T�"=;y!=�f =�M=-=�=��=z�=r[=�=�='c=n�=ِ=y=��=X=�=�
=�O	=Ω=A�=J=��=� =��<��<���<f7�<���<��</�<�5�<=b�<���<k��<M��<��<3��<.�<��<��<�&�<�.�<h5�<(:�<T=�<�>�<�>�<�<�<�8�<�3�<.-�<@%�<X�<��<��<b��<��y<��q<��i<߳a<�Y<o�Q<5�I<w�A<�9<��1<��)<S�!<�</�<��	<��<@b�;��;˵�;���;�6�;���;��;n�;0�k;bAM;��.;8a;y�:왨:eVZ:ۿ�9V��0����w�˯�����4O���-���H�q�c���}�tӋ�[���碌���v
����ȻRԻ�>߻�����7������	�fX��	�Ü����l �n�$�&�(�c�,���0��4��X8�� <���?��C���F�~�I�}/M�$qP��S�&�V���Y��]��`��'c��*f��&i��l��o��q�+�t�W�w��z��_}�����{��߂��@��Ρ�����~a�����f �����yߍ�?�����������\��,������Su��ј��+�������ޜ��6�������格f>������W祿�H�����8���Z��ж�����q��aϯ� -�������糼�D�����#����X��v������k���  �  ��N=t.N=�M=��L=� L=�pK=տJ=�J=]I=�H=�G=�FG=ǔF=��E=�0E=�~D=��C=(C=,iB=��A=fA=OQ@=��?=�>=�3>=�}==b�<=B<=4U;=H�:=y�9=�$9=�h8=��7=��6=J/6=�o5=|�4=��3=+3=�f2=/�1=��0=0=�?/=oo.=-�-=��,=��+=I+=-*=�G)=�^(=�q'=�&=L�%=�$=M�#=�"=�z!=$h =�N=�-=�=F�=��=I[=-=)�=$b=+�=R�=�=��=E=�=��
=JM	=��=1�=/H=ߎ=�� =�<��<6��<�6�<_��<L��<	�<7�</d�<���<<��<���<���<���<�<v�<i �<S*�<B2�<Y8�<�<�<v?�<m@�<�?�<#=�<�8�<-3�<	,�<�#�<)�<��<��<���<'�y<��q<��i<׫a<�Y<�Q<|�I<\�A<�9<�1<m�)<F�!<V�<z�<��	<S�<�i�;��;��;���;yE�;���;��;�~�;l;ZbM;B�.;�};F��:uǨ:��Z:6�9�у���w�C���u	�Z�1�-�-�H�G�c�s�}�����a���{����+�������Ȼf&Ի9H߻�&����������ވ	�BW�:������yg ���$�r�(�&�,�q�0�Y�4��P8�u�;�\�?��C��|F�V�I�H+M��mP�ΤS��V���Y��]� `��*c��.f��+i�r"l�bo� �q���t��w���z�$g}�Y�����ႼVC������Q��ub��e���B ��?��?ލ�`=��m���R����Y��Ʒ�����q��A͘��'��せ�ۜ��3�����!䠼|<��+���rrH��@�������\[������7��It��hү�s0��J����볼�H��ޤ��� ��=\���������)n���  �  ��N=�-N=ZM=p�L=� L=�pK=~�J=�J='^I={�H=��G=�HG=��F=��E=�2E=��D=��C=�C=�jB=I�A=|A=*R@=5�?=s�>=�3>=_}==��<=�<=;T;=�:=�9=T#9=�f8=��7=��6=b-6=n5=��4=@�3=�)3=5e2=�1=��0=g0=O?/=_o.=`�-=,�,=��+=>+=I.*=aI)=h`(=7s'=��&=*�%=ɏ$=�#=��"=T|!=�i =�O=�.=B=��=��=[=�=`�=a=��=ƍ==��=.=��=��
=K	=y�=�=<F='�=� =w�<�}�<���<�5�<���<���<��<h8�<f�<b��<��<���<��<���<�	�<U�<4$�<�-�<�5�<Z;�<[?�<�A�<B�<�@�<�=�<�8�<�2�<�*�<�!�<��<N�<[�<b��<��y<��q<��i<��a<;�Y<��Q<��I<f~A<�{9<K{1<9})<@�!<g�<��<d�	<�<q�;W��;���;�	�;T�;���;P�;��;�<l;?�M;��.;I�;���:3�:L�Z:;��9 ���}w���w�b���'�f���-�DI�8�c�(~�q�������9��]%��q�Ȼm1Ի�Q߻�.�����N!�����؈	�0V��\���
�nb ���$��(��,��0���4�6I8��;�?�?�sC��vF�N�I�?'M��jP���S��V���Y�]�]"`�$.c�3f�1i�B(l�o�Mr���t���w�X�z��n}����H����䂼�E���������vc������8 ���~��ݍ��;��P��������V����������m��eɘ�($��8~���ל��0��5����ᠼ�:��̓����)H��x��������\��R�������v��wկ��3��푲�fﳼ]L������s���_������v���p���  �  ��N="-N=�~M=K�L=!L=XqK=�J=YJ=-_I=��H=
�G=3JG=I�F=O�E=c4E=l�D=x�C=\C=lB=��A=zA=�R@=��?=��>=�3>=+}==z�<=�<=MS;=�:=��9=�!9=Fe8=	�7=)�6=�+6=@l5=�4=��3=(3= d2=�1=�0=�0=�>/=No.=��-=��,=/�+=(+=[/*=�J)=�a(=�t'=4�&=Ԍ%=s�$=��#=N�"=�}!=�j =�P=�/=�=��=��=�Z=<=��=`=��=Y�=X=��=F=�~=��
=�H	=q�=1�=kD=��=�� =�<�{�<F��<�4�<���<���<z�<�9�<�g�<���<���<���<f��<��<q�<��<�'�<61�<�8�<>�<�A�<uC�<pC�<�A�<>�<�8�<�1�<�)�<. �<��<�
�<V��<�<��y<5�q<��i<�a<��Y<��Q<!}I<�xA<�v9<Kw1<*z)<S!<~�<ޏ<��	<,�<�w�;آ�;j��;A�;�a�;'��;K$�;z��;![l;��M;|/;��;��:5�:u,[:L
�9�w��8d��w�lĴ�3)�`r���-��I���c�c~����ĩ������F���1��=�Ȼ#<Ի�Z߻b6껱���4%�����و	�)U�.�i�����] �:�$��(�v�,��0���4�HB8�#�;��?�dC�|qF���I�k#M��gP��S�)�V��Y�']�q$`�L1c�7f��5i��-l�Po��	r��t���w�w�z��u}� !��V���y炼 H������J��cd��I�) ��~��܍�0:��[���Y���T��q���4��sj���Ř�� ���z��qԜ��-�������ߠ��8�������줼�G������b ���]��������ty��hد�7��F������O��?�������b���������r���  �  )�N=�,N=�~M=&�L=.!L=�qK=��J=J=`I=ͮH=B�G=�KG=��F=��E=�5E=�D=��C=�C=DmB=��A=YA=�S@=3�?=��>=�3>=�|==�<==<=�R;=�:=��9=� 9=�c8=��7=��6=	*6=�j5=��4=_�3=�&3=�b2=1�1=k�0=_0=�>/=<o.=��-=��,=��+=�+=Q0*=�K)=c(=!v'=��&=W�%=��$=.�#=��"=�~!=�k =�Q=_0=P=;�=Ü=�Z=�=�=C_=��=�=�=]�=�=�|=��
=.G	=��=��=�B=�=f� =��<6z�<��<�3�<T��<���<�<�:�<<i�<o��<��<?��<!��<��<��<��<�*�< 4�<8;�<f@�<�C�<	E�<�D�<gB�<h>�<�8�<\1�<�(�<��<��<u�<���<H�<A�y<��q<X�i<~�a<v�Y<�~Q<�wI<�sA<�r9<�s1<�w)<�}!<��<�<��	<0�<}}�;z��;Q��;� �;m�;�Ǥ;�1�;���;Mvl;$�M;�+/;�;~6�:>�:�c[:*b�9�����S�^�w�˴�c6�c|��.�|(I���c�3~�]��d����$��}R���<���ȻWEԻ�b߻�<�����}(������	�^T�}������Y ���$�ȴ(���,��0�l}4�<8��;�+z?�F�B��lF���I�L M��eP�F�S�w�V��Y�@]�/&`��3c�l:f��9i��2l�v$o��r�3�t��w���z��{}�$�������邼J��>������3e���� ���}��8ۍ��8������R����Q��ٮ��o��mg��������w���ќ�1+��}����ݠ�x7������1줼�G������^������t���{���گ��9��I������S��T����
���e�����O���t���  �  ��N=&,N=R~M=�L=6!L=�qK=��J=�J=�`I=��H=2�G=�LG=ΚF=��E=7E=�D=��C=� C=+nB=M�A=A=T@=��?=(�>=�3>=�|==��<=�<=�Q;=-�:=��9=�9=�b8=h�7=q�6=�(6=�i5=i�4=M�3=�%3=b2=��1=��0=�
0=r>/=,o.=ʜ-=9�,=#�+=t+=1*=�L)=d(=)w'=��&=l�%=�$=7�#=��"=�!=�l =sR=�0=�=s�=Ü=�Z=v=��=�^=��=�=�=$�=B=�{=U�
=�E	=c�=/�=�A=�=o� =Y�<�x�<��<43�<��<���<��<j;�<_j�<ݒ�<���<=��<?��<O�<��<A!�<�,�<+6�<;=�<B�<6E�<5F�<�E�<�B�<�>�<�8�<�0�<�'�<��<x�<��<���<�<��y<��q<N�i<��a<��Y<�yQ<rsI<�oA<Bo9<)q1<�u)<*|!<��<�<v�	<��<���;f��;��;�(�;v�;$Ѥ;�;�;Զ�;Z�l;��M;�>/;�;�T�:eX�:5�[:)��9����I���w�\Ѵ��A���o.�5I�~�c��C~��������-���Z���E��$�ȻqLԻ<i߻�A껹���\+��Q����	��S�; �C��F��V �T�$���(���,���0��x4��78���;��u?�7�B��iF���I��M��cP��S��V�B�Y� ]��'`�6c�=f�:=i�p6l��(o�@r���t���w�c�z��}�G&��쉁��낼�K����������e��É� ��X}���ڍ�8��f������O��ά��K	��7e������o���u���Ϝ�H)��炟�dܠ�g6�������뤼�G��#�������_���������i}���ܯ��;������Q���uU���������g��º���v���  �  4�N=�+N=+~M=��L=>!L=�qK=1�J=�J=4aI=�H=��G=6MG=��F=��E=�7E=ƅD=��C=P!C=�nB=ƻA=hA=hT@=��?=B�>=�3>=�|==��<=t<=~Q;=��:=&�9=�9=b8=��7=��6=(6=�h5=��4=��3=Z%3=�a2=�1=��0=�
0=X>/=o.=ٜ-=T�,=f�+=�+=v1*= M)=�d(=�w'=g�&=$�%=��$=�#=J�"={�!=m =�R=?1=�=��=Ɯ=qZ=K=6�=.^=@�=�=)=`�=�
=�z=l�
=�D	=��=o�=�@=\�=�� =X�<x�<{��<�2�<���<���<��<�;�<k�<���<���<n��<���<��<Q�<�"�<_.�<�7�<p>�<4C�<F�<G�<F�<:C�<�>�<r8�<�0�<M'�<��<�<��<���<��<��y<��q<��i<$�a<��Y<wQ<�pI<�mA<"m9<�o1<Et)<q{!<��<�<�	<��<���;ٳ�;X��;�-�;�{�;=פ;�A�;���;8�l;Y�M;�I/;~�;�f�:5h�:��[:���9V�$E���w�մ�KI�����.��<I���c�cM~�-��3Ę��3�� a��~J��5�Ȼ�PԻ'm߻9E�:���1-������	��S���� �����U ��$�V�(��,�Р0��u4��48���;�s?���B�TgF��I�KM��bP���S���V�j�Y�]��(`�`7c��>f�O?i��8l�S+o��r���t���w���z��}��'��9����삼�L��X���"	��Qf��EÉ�) ��'}��5ڍ�f7���������N����������c��"������_t��_Μ� (��ف���۠��5��<����뤼uG��D������X`��[������v~��ޯ�D=��雲�����W��@�����*i��Dú����v���  �  �N=�+N=~M=��L=F!L=	rK=G�J=J=RaI=L�H=��G=kMG=��F=��E=8E=��D=��C=�!C=�nB=��A=�A=�T@=ϟ?=V�>=�3>=�|==z�<=X<=bQ;=�:=��9=�9=�a8=^�7=q�6=�'6=�h5=��4=b�3="%3=`a2=�1=k�0=�
0=H>/=o.=�-=i�,=��+=�+=�1*=]M)=�d(=x'=��&=Z�%=��$=�#=y�"=��!=Zm =�R=\1==��=ל=bZ=6=�=	^=�=J�=�=�=@
=gz=@�
=�D	=/�=/�=�@="�=�� =�<�w�<G��<�2�<ҁ�<��<��</<�<Tk�<��<"��<���<��<&�<��<$#�<�.�<�7�<�>�<�C�<TF�<@G�<9F�<aC�<�>�<X8�<}0�<'�<��<#�<5�<��<�<��y<x�q<t�i<2�a<�Y<vQ<�oI<�lA<nl9<o1<�s)<+{!<r�<B�<?�	<�<���;��;&��;�/�;�}�;+٤;�C�;���;Úl;8�M;�M/;��;$m�:�l�:��[:��9��~�;D�ދw�s״�rL�j��H.��?I�� d� Q~�w���Ř��4��8c��YL��7�Ȼ�RԻ�n߻sF�&���.��ݟ�>�	�BS�a����� ���T ��$���(��,��0�u4��38��;�Mr?��B�ZfF�|�I��M�MbP�;�S�i�V���Y��]�)`��7c�c?f�
@i��9l�Z,o��r���t���w�L�z�B�}�(������)킼M������[	��}f��^É�1 ���|��ڍ�)7��\�����eN��.���y��bc����������s���͜��'��k���V۠�j5�����Y뤼ZG��Z��� ���`������+���~��xޯ��=��l���s���BW���������i���ú���Sw���  �  4�N=�+N=+~M=��L=>!L=�qK=1�J=�J=4aI=�H=��G=6MG=��F=��E=�7E=ƅD=��C=P!C=�nB=ƻA=hA=hT@=��?=B�>=�3>=�|==��<=t<=~Q;=��:=&�9=�9=b8=��7=��6=(6=�h5=��4=��3=Z%3=�a2=�1=��0=�
0=X>/=o.=ٜ-=T�,=f�+=�+=v1*= M)=�d(=�w'=g�&=$�%=��$=�#=J�"={�!= m =�R=@1=�=��=Ȝ=rZ=M=8�=0^=C�=��=-=d�=�
=�z=r�
=�D	=��=w�=�@=f�=�� =l�<,x�<���<�2�<��<��<��<<�<'k�<œ�<���<w��<���<��<R�<�"�<Z.�<�7�<g>�<(C�<F�<�F�<�E�<)C�<�>�<a8�<�0�<='�<��<q�<��<���<��<��y<|�q<��i<)�a<��Y<wQ<�pI<�mA<>m9<�o1<ft)<�{!<<;�<�	<��<���;��;���;�-�;�{�;Oפ;�A�;���;�l;$�M;�I/;�;�e�:/g�::�[:���9{H��G�^�w�~ִ��J�v��:.�d=I���c��M~�u��uĘ��3��7a���J��a�Ȼ�PԻJm߻WE�T���H-�����#�	��S����$�����U ��$�X�(��,�Ҡ0��u4��48���;�s?���B�TgF��I�LM��bP���S���V�j�Y�]��(`�`7c��>f�P?i��8l�S+o��r���t���w���z��}��'��9����삼�L��X���"	��Qf��EÉ�) ��'}��5ڍ�f7���������N����������c��"������_t��_Μ� (��ف���۠��5��<����뤼uG��D������X`��[������v~��ޯ�D=��雲�����W��@�����*i��Dú����v���  �  ��N=&,N=R~M=�L=6!L=�qK=��J=�J=�`I=��H=2�G=�LG=ΚF=��E=7E=�D=��C=� C=+nB=M�A=A=T@=��?=(�>=�3>=�|==��<=�<=�Q;=-�:=��9=�9=�b8=h�7=q�6=�(6=�i5=i�4=M�3=�%3=b2=��1=��0=�
0=r>/=,o.=ʜ-=9�,=#�+=t+=1*=�L)=d(=)w'=��&=l�%=�$=7�#=��"=�!=�l =tR=�0=�=u�=Ŝ=�Z=y=��=�^=��=$�=�=-�=L=�{=a�
=�E	=r�=@�=�A=�=�� =��<y�<6��<\3�<9��<	��<��<�;�<}j�<���<���<N��<K��<V�<��<>!�<�,�<6�<)=�<B�<E�<F�<nE�<�B�<t>�<j8�<�0�<�'�<v�<]�<��<���<��<{�y<�q<N�i<��a<��Y<zQ<�sI<	pA<wo9<dq1<�u)<l|!<A�<J�<��	<��<5��;ϰ�;_��;)�;Jv�;GѤ;�;�;̶�;�l;D�M;>/;N�;�R�:lV�:χ[:���9���+O�-�w�!Դ�hD�����.�V6I���c��D~�������.��6[���E��z�Ȼ�LԻi߻B������+��c���	��S�F �L��N��V �Y�$�İ(���,���0��x4��78���;��u?�8�B��iF���I��M��cP��S��V�B�Y� ]��'`�6c�=f�:=i�q6l��(o�@r���t���w�c�z��}�G&��쉁��낼�K����������e��É� ��X}���ڍ�8��f������O��ά��K	��7e������o���u���Ϝ�H)��炟�dܠ�g6�������뤼�G��#�������_���������i}���ܯ��;������Q���uU���������g��º���v���  �  )�N=�,N=�~M=&�L=.!L=�qK=��J=J=`I=ͮH=B�G=�KG=��F=��E=�5E=�D=��C=�C=DmB=��A=YA=�S@=3�?=��>=�3>=�|==�<==<=�R;=�:=��9=� 9=�c8=��7=��6=	*6=�j5=��4=_�3=�&3=�b2=1�1=k�0=_0=�>/=<o.=��-=��,=��+=�+=Q0*=�K)=c(=!v'=��&=X�%=��$=.�#=��"=�~!=�k =�Q=a0=R=>�=Ɯ=�Z=�=�=I_=��=#�=�=i�=�=�|=��
=AG	=��=��=C=-�=�� =/�<oz�<H��<4�<���<	��<K�<�:�<fi�<���<��<W��<3��<"��<��<��<�*�<�3�<;�<H@�<�C�<�D�<wD�<9B�<9>�<�8�<.1�<~(�<��<��<U�<���<3�<$�y<��q<X�i<��a<��Y<�~Q<�wI<�sA<�r9<)t1<�w)<�}!<�<e�<�	<��<"~�;��;���;!�;am�;�Ǥ;�1�;�;�ul;��M;�*/;�;4�:J;�:_][:�T�9�ˀ�E[��w��δ�M:�Q~��.�L*I���c��4~�!�����]%��S��s=����Ȼ�EԻ@c߻ =�����(�������	�qT��������Y ���$�δ(��,��0�p}4�
<8��;�-z?�G�B��lF���I�M M��eP�G�S�w�V��Y�@]�/&`��3c�l:f��9i��2l�w$o��r�3�t��w���z��{}�$�������邼J��>������3e���� ���}��8ۍ��8������R����Q��ٮ��o��mg��������w���ќ�1+��}����ݠ�x7������1줼�G������^������t���{���گ��9��I������S��T����
���e�����O���t���  �  ��N="-N=�~M=K�L=!L=XqK=�J=YJ=-_I=��H=
�G=3JG=I�F=O�E=c4E=l�D=x�C=\C=lB=��A=zA=�R@=��?=��>=�3>=+}==z�<=�<=MS;=�:=��9=�!9=Fe8=	�7=)�6=�+6=@l5=�4=��3=(3= d2=�1=�0=�0=�>/=No.=��-=��,=/�+=(+=[/*=�J)=�a(=�t'=4�&=Ԍ%=s�$=��#=O�"=�}!=�j =�P=�/=�=��=��=�Z=A=��=$`=��=e�=e=�=W=�~=��
=I	=��=M�=�D=��=�� =I�<!|�<���<�4�<���<���<��<�9�<�g�<���<۱�<���<{��<��<t�<��<�'�<1�<|8�<�=�<uA�<DC�<;C�<gA�<�=�<�8�<�1�<t)�<��<��<�
�<5��<��<h�y<#�q<��i<%�a<�Y<ׄQ<c}I<yA<w9<�w1<�z)<�!<�<T�<�	<��<�x�;���;��;��;b�;c��;c$�;m��;�Zl;�M;�/;��;��:��:�$[:���9J���mm�_�w�8ɴ��-�t���-��I�	�c�d ~� �����������G��[2����Ȼ�<ԻL[߻�6�	����%�������	�@U�B�y�����] �C�$���(�}�,��0���4�LB8�&�;��?�fC�}qF���I�l#M��gP��S�*�V��Y�(]�q$`�L1c�7f��5i��-l�Po��	r��t���w�w�z��u}� !��V���y炼 H������J��cd��I�) ��~��܍�0:��[���Y���T��q���4��sj���Ř�� ���z��qԜ��-�������ߠ��8�������줼�G������b ���]��������ty��hد�7��F������O��?�������b���������r���  �  ��N=�-N=ZM=p�L=� L=�pK=~�J=�J='^I={�H=��G=�HG=��F=��E=�2E=��D=��C=�C=�jB=I�A=|A=*R@=5�?=s�>=�3>=_}==��<=�<=;T;=�:=�9=T#9=�f8=��7=��6=b-6=n5=��4=@�3=�)3=5e2=�1=��0=g0=O?/=_o.=`�-=,�,=��+=>+=I.*=aI)=h`(=8s'=��&=+�%=ɏ$=�#=��"=U|!=�i =�O=�.=E=��=��=[=�=h�=&a=��=ҍ==ė=A=Ҁ=��
=+K	=��=8�=^F=K�=1� =��<&~�<���<�5�<B��<���<�<�8�<Af�<���<9��<���<7��<���<�	�<O�<$$�<�-�<c5�<1;�<*?�<OA�<�A�<v@�<Y=�<�8�<S2�<�*�<�!�<��<!�<6�<E��<g�y<��q<��i<ˣa<a�Y<ËQ<�I<�~A<�{9<�{1<�})<��!<�<%�<�	<[�<�q�;!��;d��;{
�;~T�;Ѭ�;l�;�;<l;{�M;��.;�;n��:c�:��Z:���9����Á�;�w��´��Pi�N�-��I���c�d	~�|w������[:��&���Ȼ 2ԻbR߻A/�(����!�������	�JV��n���
�zb ���$��(��,�
�0���4�9I8��;�A�?�uC��vF�O�I�@'M��jP���S��V���Y�]�]"`�$.c�3f�1i�B(l�o�Mr���t���w�X�z��n}����H����䂼�E���������vc������8 ���~��ݍ��;��P��������V����������m��eɘ�($��8~���ל��0��5����ᠼ�:��̓����)H��x��������\��R�������v��wկ��3��푲�fﳼ]L������s���_������v���p���  �  ��N=t.N=�M=��L=� L=�pK=տJ=�J=]I=�H=�G=�FG=ǔF=��E=�0E=�~D=��C=(C=,iB=��A=fA=OQ@=��?=�>=�3>=�}==b�<=B<=4U;=H�:=y�9=�$9=�h8=��7=��6=J/6=�o5=|�4=��3=+3=�f2=/�1=��0=0=�?/=oo.=,�-=��,=��+=I+=-*=�G)=�^(=�q'=�&=M�%=�$=N�#=�"=�z!=&h =�N=�-=�=J�=��=N[=4=1�=-b=6�=_�=�=��=Y= �=��
=eM	=ħ=R�=RH=�=�� =[�<6��<���<�6�<���<���<Q�<T7�<jd�<1��<g��<���<���<��<�<o�<Y �<9*�<2�<.8�<�<�<>?�<0@�<b?�<�<�<�8�<�2�<�+�<W#�<��<��<Z�<���<��y<��q<��i<�a<F�Y<N�Q<ȊI<��A<K�9<�1<�)<˃!<ވ<�<y�	<ѥ<�j�;���;���;v��;�E�;;��;�~�;�l;�aM;"�.;m|;ר�:�è:ΗZ:�"�9#��d���w�ͻ����T]���-���H���c���}��ዻa���e���U,�����j�Ȼ�&Ի�H߻5'�3���p�������	�]W�Q�������g ���$�{�(�.�,�w�0�]�4��P8�x�;�^�?��C��|F�W�I�I+M��mP�ϤS��V���Y��]� `��*c��.f��+i�r"l�bo�!�q���t��w���z�$g}�Y�����ႼVC������Q��ub��e���B ��?��?ލ�`=��m���R����Y��Ʒ�����q��A͘��'��せ�ۜ��3�����!䠼|<��+���rrH��@�������\[������7��It��hү�s0��J����볼�H��ޤ��� ��=\���������)n���  �  ��N=/N=#�M=��L=� L=.pK=&�J=�J=�[I=��H=~�G=0EG=�F=��E=�.E=�|D=.�C=rC=�gB=��A=CA=pP@=��?=��>=�3>=�}==��<=�<=#V;=u�:=��9=}&9=]j8=o�7=��6=816=�q5=F�4=��3=~,3=�g2=;�1=��0=�0=�?/=so.=��-=.�,=�+=J+=�+*=�F)=?](=�o'=�}&=p�%=�$=��#=T�"=<y!=�f =�M=-=�=��=~�=w[=�=�=0c=y�=�=�=��=k=#�= �
=�O	=�=`�=4J==D� =��<:��<��<�7�<���<^��<t�<�5�<vb�<ʈ�<���<n��<��<A��<1�<��<��<�&�<�.�<>5�<�9�<=�<�>�<L>�<[<�<�8�<�3�<�,�<%�<%�<��<t�<F��<��y<��q<��i<�a<'�Y<��Q<�I<ЊA<i�9< �1<�)<Ӆ!<��<��<	�	<)�<"c�;߇�;y��;��;�6�;���;8��;n�;��k;�@M;��.;�_;�u�:��:�MZ:`��9�a��v��E�w�$�������Q�O�-�6�H�ϒc���}�ԋ�S���𤻏��0��E�Ȼ�Ի%?߻��[������ٚ�8�	�X��	�՜�	��l �x�$�.�(�j�,� �0��4��X8�<���?��C���F��I�~/M�%qP��S�'�V���Y��]��`��'c��*f��&i��l��o��q�+�t�W�w��z��_}�����{��߂��@��Ρ�����~a�����f �����yߍ�?�����������\��,������Su��ј��+�������ޜ��6�������格f>������W祿�H�����8���Z��ж�����q��aϯ� -�������糼�D�����#����X��v������k���  �  o�N=�/N=z�M=��L=� L=�oK=|�J=�J=�ZI=u�H=��G=�CG=@�F=
�E=-E=/{D=��C=�C=3fB=e�A=7A=�O@=^�?=j�>=�3>=�}==7�<=�<=W;=��:=1�9=�'9=�k8=!�7=u�6=�26=ws5=�4=�3=�-3=�h2=5�1=W�0=0=3@/=xo.=��-=��,=J�+=U+=�**=9E)=�[(=,n'=5|&=��%=V�$=̉#=Ń"=�w!=e =uL=,,=V=��=`�=�[==��=#d=��=D�=&=e�=V="�="�
=�Q	=�=H�=�K=^�=�� =;�<��<M��<�8�<B��<��<��<�4�<�`�<���<ئ�<`��<���<���<���<��<�<5#�<�+�<p2�<�7�<;�<�<�<E=�<�;�<�8�<4�<�-�<�&�<%�<�<c�<��<��y<��q<=�i<<�a<a�Y<y�Q<їI<h�A<�9<�1<Ɔ)<��!<b�<N�<��	<��<�[�;�~�;���;]��;;)�;E~�;��;$^�;��k;R"M;g�.;�D;�E�:@l�:�Z::@�9����K����w�	��� ���F�g�-��H��}c�ʿ}�
ȋ��t��㤻�������ҩȻ�Ի�6߻b�ڷ��=�� ��e�	��Y������|q ��$�o�(���,��0�G�4��_8�<�$�?��C�@�F�9�I��3M�JtP��S�A�V���Y��]�(`��$c��&f�R"i�!l��o�v�q�R�t�w�w�E�z��X}�����x��r܂��>������� ���`������� �����������@������\ ���_��R������x���Ԙ�T/�������᜼�9��b����蠼:@������2�+I����������Y��3�����$o���̯�*��R���|䳼:A�����������U����������i���  �  �N=-0N=M=��L=c L=ioK=�J=J=�YI=N�H=��G=6BG=��F=~�E=w+E=�yD=�C=�C=�dB=I�A=QA=�N@=ۛ?=�>=�3>=~==��<=!<=�W;=x�:=D�9=6)9=Lm8=��7= �6={46=�t5=N�4=b�3=/3=�i2=	�1=��0=0=h@/=~o.=|�-=P�,=��+=�+=�)*=D)=|Z(=�l'=�z&=,�%=Ј$=P�#=\�"=�v!=[d =�K=q+=�=6�=>�=�[=n=.�=�d=� =x�=}=�=�=�=��
=jS	=��=� ={M=��=�� =&�<���<p��<09�<t��<���<� �<l3�<_�<���<���<ѿ�<���<���<l��<�	�<��<F �<�(�<�/�<y5�<`9�<�;�<[<�<Q;�<�8�<{4�<�.�<�'�<��<"�<��<<�<��y<�q<��i<��a<��Y<6�Q<�I<�A<�9<�1<,�)<�!<��<ݎ<;�	<[�<�U�;�v�;��;���;F�;q�;ה;OP�;<�k;9M;��.;�-;F�:�H�:�Y:'��9������w�1�������=���-��H��kc�J�}�.���9i���פ�k��o���&�Ȼ�Ի�.߻J껃���5��d����	��Z������w��u ��$���(���,�H�0���4�7f8�L<��?� C�$�F�^�I��6M��vP�ЪS�T�V��Y�:]��`��"c��#f�Vi��l�� o��q�L�t�M�w��z�
S}����fv��Aڂ��<������n����_��W���� ��&����፼B��u������!b���������{���ט�o2��	����䜼d<�������꠼�A��!����𤼌I��ע�����X��峫�@��m��*ʯ�d'��~���q᳼/>����������S��+���p��h���  �  ��N=�0N=�M=��L=B L=oK={�J=iJ=
YI=n�H=��G=AG=��F=X�E=G*E=�xD=��C=pC=dB=n�A=� A=MN@=p�?=��>=h3>=~==��<=�<=JX;=0�:=�9=,*9=Xn8=��7=�6=�56=v5=a�4=h�3=�/3=�j2=��1=g�0=�0=�@/=}o.=L�-=��,=/�+=�
+=�(*=&C)=yY(=�k'=�y&=�%=��$=A�#=F�"=�u!=c =�J=�*=Z=��=!�=�[=�=��={e=e=c�=�=�=-=#�=5�
=�T	=�==�N=��=�� =��<���<G��<�9�<���<���<X �<2�<�]�<���<���<���<���<d��<��<Z�<��<��<�&�<.�<�3�<	8�<�:�<�;�<�:�<�8�<�4�<�/�<�(�<I!�<��<��<c�<�y<��q<j�i<��a<4�Y<��Q</�I<��A<3�9<h�1<��)<�!<A�<x�<�	<��<�P�;�p�;x��;]��;��;hg�;�̔;�E�;�k;��L;�m.;�;���:�,�:��Y:4��9Cz����r�w��������7���-��H�^c���}�C����`��VϤ�!���X켻m�ȻfԻ8)߻��5����������	��[��ˤ�+��x ���$���(�}�,���0�Y�4��j8��<���?�:$C�֐F���I��9M�yP�_�S�2�V�(�Y��
]�<`�� c�V!f�Ii�6l���n���q���t��w��{z��N}����qt���؂�Z;��_�������j_��2���� ������a⍼5C��֣��<��d��Ô�F!��/~��ژ��4��@����朼c>������@젼C��������I��Т������ZW��������k��Xȯ�S%��W���4߳��;��g�������Q��O����	���f���  �  ��N=�0N=�M=��L=0 L=�nK=/�J=J=�XI=�H=%�G=q@G=�F=��E=})E=�wD=4�C=�C=icB=�A=$ A=�M@=*�?=��>=X3>=~==��<=�<=�X;=��:=��9=�*9=o8=`�7=��6=Z66=�v5=�4=�3=u03=3k2=�1=��0=�0=�@/=uo.=8�-=��,=��+=}
+=k(*=�B)=�X(=k'=�x&=>�%=�$={�#=��"=�t!=�b =FJ=y*==��=�=�[=�=��=�e=�=�=*=ɠ=�=��=�
=�U	=��=�=VO=X�=?� =��<q��<���<�9�<���<m��<���<�1�<]�<���<���<k��<[��<���<k��<��<�<��<�%�<�,�<�2�<67�<�9�<6;�<�:�<�8�<�4�<�/�<�)�<"�<��<��<��<��y<��q<��i<��a<3�Y<z�Q<��I<��A<��9<��1<�)<��!<m�<?�<|�	<_�<�M�;�l�;��;���;��;)a�;�Ŕ;�>�;��k;��L;�a.;};���:��:i�Y:uk�9戸n����w�����J��2��-�P�H��Uc�&�}�����b[���ɤ������漻ӓȻ)�ӻ�%߻�
�����������	�(\��#����{ ��$�~�(��,���0���4�3n8��<�:�?��&C��F���I�>;M�RzP�I�S���V�N�Y�{
]��`��c��f��i��l�_�n���q��t�ޠw��xz��K}����Cs���ׂ��:���������3_������ ��ہ���⍼�C������D��2e��mĔ��"������ۘ�]6������蜼�?������@��C���������I��Т�������V��?������j��9ǯ�$�������ݳ�q:������^󷼼O��,�������e���  �  6�N=)N=uxM=e�L=�L=�cK=��J=��I=�KI=d�H=��G=v1G=~F=��E=YE=dD=��C=��B=�JB=�A=6�@=�.@=�y?=P�>=�>=�V==J�<=�;=�*;=�o:=��9=��8=}88=oy7=W�6=/�5=�55=r4=�3=>�2=�2="S1=e�0=A�/=v�.=�.=09-=X^,=�+=l�*=�)=��(=��'=1�&=��%=J%=;$=�"=m�!=�� =��=^�=s�=$f=H4=��=��=on=�=��=�\=��=f|=��=�z=g�=VZ
=�=d=&s=Y�=Z=SQ =;�<��<L��<�U�<��<���<9�<�t�<(��<	��<��<'�<{G�<
d�<�}�<��<=��<;��<<ʸ<uش<��<��<���<���<~�<�	�<@�<q�<f�<n�<�
�<e�<��<z<� r<��i<A�a<��Y<7�Q<��I<��A< :<�	2<�*<�"<.<�><S
<Ej<H�;�J�;Δ�;~��;WP�;UŦ;�K�;&�;�)q;b�R;To4;�\;.��:�:��u:�� :�kN8�˹��W�'&����ۺt	���$��t?�I�Y�!�s��Æ��X�������ѫ������Sû!�λF�ٻռ�aﻕ���>�����M��i~��������K"��{&�l�*�K�.��r2��@6���9���=��+A��D��H��tK�g�N��	R�uBU�TqX���[���^���a�1�d���g��j�+�m�b�p�/�s��v��y�M`|�:���Tq��Rك� @�����8���o��vԊ��8��d�������6c��Ƒ�'(������ꕼ�I��駘�S���a��4������%r��̠��%�����ڤ��4��,���쨼�H��ץ��s��ia������7���|��B۳��9�����Z����T��I�����Mq���  �  &�N=�(N=fxM=i�L=�L=�cK=��J=��I=�KI=��H=#�G=�1G=8~F=��E=~E=NdD=-�C=��B=�JB=-�A=L�@=�.@=z?=Y�>=�>=�V===�<=�;=�*;=�o:=|�9=`�8=N88=Fy7=*�6=��5=�55=�q4=Ƭ3=�2=�2=S1=U�0=4�/=p�.=�.=89-=k^,=0�+=z�*=�)=��(=��'=b�&=��%=q%=`$=:�"=��!=0� =��=��=��=1f=X4=��=��=gn=�=��=�\=��=2|=t�=�z=7�=Z
=��=2=�r="�=$=1Q =�<���<��<�U�<���<���<9�<u�<F��<P��<��<r'�<�G�<sd�<�}�<s��<���<���<�ʸ<�ش<#�<��<���< �<��<�	�</�<_�<P�<R�<p
�<�<U�<Zz<( r<��i<��a<��Y<l�Q<-�I<��A<�:<G	2<A*<["< .<?<%S
<}j<|�;fK�;��;���;�Q�;Ǧ;uM�;z�;o-q;�R;�r4;�_;h �:��:��u:�� :�N8��˹�W�x&����ۺ]t	���$�zv?�x�Y���s��Ć��Y��d����ҫ����UûS�λ�ٻ8��ua�����K����� ��~�h�>��p�OK"��z&���*�m�.�Hr2��?6���9�Κ=��*A���D�H�dtK�#�N�8	R�XBU�qX���[���^���a�t�d�)�g�-�j���m�.�p�Ƿs�۟v�˂y��`|��:�c���q���ك�>@�����R���o��UԊ�r8��C�������
c���ő��'��9����镼%I���������Ka��м������q���ˠ��%������٤��4�����'쨼�H����������a��	������}���۳��9��k�������,U������\��pq���  �  ��N=�(N=MxM=`�L=�L=dK=ڱJ='�I=1LI=�H=��G= 2G=�~F=a�E=E=�dD=��C=r�B=KB=��A=��@=8/@==z?=s�>=�>=zV==#�<=��;=�*;=Mo:=�9=��8=�78=�x7=��6=m�5=55=kq4=\�3=��2=02=�R1=�0=�/=X�.=�.=G9-=�^,=o�+=ɞ*=z�)=K�(=)�'=��&=;�%=%=�$=��"=�!=�� =�=�=Ȑ=if=y4=��=��=An=�=@�={\=C�=�{=��=&z=��=qY
=�=�=Qr=��=�=�P =5�<+��<���<bU�<��<���<Z9�<vu�<ߪ�<��<��<[(�<�H�<�e�<�~�<���<���<���<�˸<�ٴ<��<y�<Q��<h �<��<�	�<�<"�<��<��<�	�<C�<p�<4z<��q<z�i<9�a<�Y<r�Q<e�I<�A< :<�2<s*<�"<�-<)?<�S
<dk<��;xN�;]��;���;�U�;l˦;�R�;��;�7q;��R;�{4;�g;�:���:l�u:I� :ۇO8��˹�W��&����ۺ�w	��$��{?���Y�<�s�pȆ��]��o���s֫�˶��Xû"�λ��ٻ���cﻼ������������Y}�T�������I"�y&���*�A�.��o2��=6�{�9��=��(A��D�sH�sK��N��R�BU�qX�
�[�9�^���a���d���g���j�z�m�8�p�޹s��v� �y��b|��<�.	��nr��5ڃ��@��������!p��AԊ�C8��؛��V���Xb���đ�'��E����蕼H��r������E`��⻜����q��
ˠ�%��.���٤��4��)���Z쨼I��z���?��vb������p��~���ܳ�;��|�������V��j���"��r���  �  ��N=�(N=$xM=V�L=L=SdK=&�J=��I=�LI=��H=R�G=�2G=�F==�E=�E=�eD=��C=I�B=�KB=0�A=*�@=�/@=z?=��>=�>=gV==�<=�;=#*;=�n:=v�9=<�8=78=�w7=Ƿ6=��5=545=�p4=��3=��2=�2=MR1=��0=̶/=9�.=�.=o9-=�^,=ɀ+=>�*=�)=��(=��'=��&=�%=�%=�$=��"=��!=f� =��=e�=4�=�f=�4=��=��=n=,=˿=�[=��=�z=�=5y=��=vX
=�=�=^q=��=�=
P =�<0��<���<�T�<���<���<�9�<v�<���<��<��<�)�<J�<Cg�<���<f��<���<n��<7͸<۴<*�<�<��<� �<)�<�	�<��<��<(�<�
�<}�<��<��<��y<R�q<�i<��a<��Y<�Q<(�I<W�A<��9<E2<�*<�"<S-<\?<@T
<~l<e�;�R�;���;���;:]�;�Ҧ;Z�;d�;Gq;��R;b�4;�u;-(�:bѵ:y�u:�� :c�P8I�˹�W�)����ۺ�{	���$� �?��Y�C t��Ά�d��a����ܫ������]ûO�λ��ٻ��仌eﻘ������`��	��\|������y���F"��u&�3�*�ć.�kl2�:6��9�g�=��%A��D�)H�+qK���N��R�[AU��pX�}�[�B�^��a�e�d���g�u�j���m�c�p�X�s�b�v�W�y�hf|��?��
���s��Iۃ��A��1������Pp��/Ԋ��7��Y�������Ya���Ñ��%�������敼QF���������^��)���.���o���ɠ�,$���~��@٤�n4��6����쨼�I��/���4���c��F¯�!�����Z޳��<��0���j����W��⵺�X��s���  �  �N=(N=�wM=J�L=,L=�dK=��J=1 J=kMI=u�H=A�G=�3G=��F=c�E=E=�fD=��C=B C=�LB=�A=��@=50@=�z?=��>=>=XV==��<=�;=�);=n:=��9=N�8=68=�v7=��6=v�5=35=�o4=��3=!�2=�2=�Q1=E�0=u�/=�.=�.=�9-=_,=H�+=ݟ*=ź)=��(=��'=��&=,�%=�%=�$=� #=��!=L� =��=�=ő=(g=�4=��=k�=�m=�=0�=)[=��=�y=��=x=I�=W
=��=E=/p=��=�
=O =��<��<��<}T�<���<���<*:�<w�<߬�<���<��<�+�<�L�<�i�<��<���<ԭ�<���<4ϸ<�ܴ<��<��<��<��<��<�	�<��<��<1�<h	�<��<��<� �<��y<��q<"�i<��a<k�Y<��Q<,�I<��A<��9<�2<�*<�"<�,<�?<5U
<+n<!�;�X�;��;���;�e�;uܦ;-d�;���;�[q;��R;��4;G�;�H�:��:xv::�R8��˹!�W��+��p�ۺ^�	��$��?��Z�
t�7ֆ�Jl���Ɵ��䫻ķ��dû��λ��ٻ\���h�����7��A��A���z���W��Q��(C"��q&��*�3�.��g2�m56�p�9��=��!A�p�D� H��nK�t�N�?R��@U��pX���[�v�^���a���d���g���j�X�m�\�p���s���v��y��j|��C����du���܃��B��������pp��Ԋ�n7������h���`��!��#�������䕼D��a�������R\�����N���m���Ƞ��"���}���ؤ�.4��I����쨼fJ��1������9e��	į��"�������೼
?��p���}����Y���������~t���  �  [�N=�'N=�wM=4�L=HL=�dK=�J=� J=BNI=f�H=]�G=75G=��F=��E=rE=1hD=ߴC=|C=�MB=�A=��@=�0@=^{?="�>=>=6V==g�<=��;=�(;=Am:=��9=5�8=�48=�u7=]�6=%�5=�15=Pn4=v�3=�2=�2=�P1=��0=�/=��.=�.=�9-=x_,=Ё+=��*=��)=��(= �'=��&=m�%=G%=3$=�#=�!=l� =r�=�=j�=�g=*5=��=K�=ym=<=|�=>Z=��=�x=��=�v=��=�U
=)�=�=�n=<�=�	=N =��<���<��<�S�<H��<��<�:�<�w�<:��<C��<��<&.�<O�<'l�<Ʌ�<|��<w��<%¼<�Ѹ<
ߴ<��<U��<L��<p�<��<�	�<1�<6�< 
�<��<�<��<\��<�y<K�q<��i<T�a<��Y<{�Q<}�I<��A<�9<� 2<*<p"<@,<�?<;V
<p<H�;n_�;׭�;P�;up�;��;�o�;�
�;Ssq;q�R;9�4;w�;�l�:�:�:v:�F:�YT8^i˹S�W�'/����ۺ��	�A�$�̛?�UZ��t��߆��u���П�>�ͷ��mû+�λ�ٻ����l�?��������d��Iy�V�Y�����?"�.m&��*��}.�Sb2�06�6�9� �=��A�h�D�dH��kK�8�N��R��?U��pX���[�ҷ^��a���d�I�g���j���m�~�p���s�.�v��y��o|��H����Ow��`ރ�5D��������p�� Ԋ��6������<���w^��M����!��B���J╼hA����������Y������
��l���Ơ��!���|��ؤ��3��e���w�&K��m�����g��!Ư�R%��V���㳼�A��������� \��͹�����	v���  �  ��N=:'N=^wM=&�L=mL=3eK=��J=�J=)OI=m�H=��G=~6G=P�F=#�E=�E=�iD=6�C=�C=�NB=�A=��@=o1@=�{?=e�>=;>=V==	�<=�;=)(;=bl:=��9=
�8=�38=1t7=�6=��5=w05=�l4=G�3=��2=2=#P1=�0=��/=��.=�.=�9-=�_,=Z�+=M�*=��)=��(=2�'=4�&=� &=�%=�$=D#=Y�!=�� =r�=̶=�=h=n5=��=3�=m=�=��=KY=y�=Sw=*�=�t=1�=�S
=~�=&=+m=ѽ=E=�L =��<��<���< S�<��<;��<];�<�x�<���<��<�
�<�0�<�Q�<�n�<���<a��<I��<�ļ<Ը<A�<��<���<{��<;�<_�<�	�<�
�<Q
�<��<J�<
�<t��<���<~�y<k�q<W�i<U�a<�Y< �Q<^�I<�A<X�9<��1<�
*<�"<�+<!@<LW
<r<� �;�f�;o��;A�;n{�;N�;N|�;�;ǌq;�S;��4;�;p��:�/�:5pv:q:BV8�@˹	�W��4��� ܺ��	���$�Ϫ?��"Z��1t�v醻���F۟������׷�Uvû��λ�ٻp�仝q�J���������w���w���4������:"�4h&��|*�Vx.��\2�Q*6���9�Ԇ=��A��D��H�vhK��N�	R�?U��pX�|�[�}�^���a���d��g�k�j���m���p�=�s��v���y�Du|��M����y��*����E��$������q���ӊ�6��՘������\��R���g������ߕ��>��眘�H���W���������i���Ġ�< ���{��bפ��3��s���L��ͪ���	��i��tȯ��'������峼�D��â��� ��s^��!�������w���  �  �N=�&N=wM=�L=L=�eK=�J=7J=�OI=z�H=��G=�7G=��F=��E=ME= kD=��C=�C=#PB=�A=N�@=2@=I|?=��>=?>=�U==��<=��;=t';=uk:=��9=��8=D28=�r7=��6=J�5=/5=�k4=�3=��2=2=NO1=t�0==�/=d�.=�.=:-=5`,=�+=	�*=t�)=��(=Y�'=v�&= &=%=�$=�#=��!=�� =��=��==�h=�5=��=��=�l==�=NX=N�=v=��=os=��=@R
=ն=�=�k=\�=�=�K =��<���<���<eR�<���<k��<�;�<�y�<��<���<��<�2�<HT�<�q�<���<B��<��<rǼ<�ָ<��<{�<���<���<�<��<�	�<:
�<v	�<p�<��< �<��<8��<��y<r�q<_�i<E�a<.�Y<��Q<C�I<��A<U�9<��1<M*<K"<�*<5@<}X
<t<j&�;�m�;L��;0�;��;��;���;�#�;Υq;M-S;�4;��;��:P�:g�v:��:�:X8�$˹
�W�W9���ܺf�	���$��?��3Z��Dt�}�y����埻���᷻�û�λb�ٻ����u�(���Q���������u�������*6"�gc&�[w*��r.��V2��$6���9���=�>A�w�D��H�meK�|�N�aR�?>U��pX�O�[��^���a�
�d���g���j���m��p���s���v�c�y��z|�)S�����{��	⃼+G��9������gq���ӊ��5�������9[��c�����_}���ܕ��;�����v���ST������T���g��Cà����~z���֤�g3�������M�����p��k���ʯ�G*�������購gG������{���`��t������xy���  �  ^�N=?&N=�vM=��L=�L=�eK=��J=�J=�PI=f�H=��G=�8G=��F=��E=�E=BlD=ظC=#C=.QB=֜A=�@=�2@=�|?=��>=I>=�U==`�<=	�;=�&;=�j:=��9=��8=18=�q7=2�6=��5=�-5=kj4=Х3=��2=2=�N1=߂0=ʴ/=,�.=�.=>:-=�`,=d�+=��*=C�)=��(=r�'=��&=\&=N	%=9
$=�#=��!=�� =o�=g�=g�=�h=�5=��=ٷ=hl=�=4�=bW=9�=�t=O�=�q=	�=�P
=F�==)j=��=�=�J =�<��<���<�Q�<x��<���<r<�<�z�<^��<w��<��<!5�<�V�<@t�<8��<ܤ�<���<ʼ<�ظ<��<1�<���<���<��<�<�	�<�	�<��<;�<��<��<���<���<��y<��q<��i<��a<��Y<@�Q<t�I<[�A<��9<��1<�*<�"<D*<h@<nY
<�u<�+�;Dt�;��;Q%�;���;T
�;ғ�;�/�;��q;�DS;��4;��;���:�n�:��v:��:v�Y8_˹D�W�^>��8ܺɤ	�K�$�4�?��CZ��Vt�����_��������귻Ɉû��λ"ڻ-��z�K���������˾�t�r������/2"��^&�5r*��m.��Q2�B6���9�h|=��A�x�D�h H�ybK�e�N� R�x=U��pX��[���^��a��d�x�g���j�X�m���p��s��v���y��|�X�����}���ー�H��K���R���q���ӊ��5��8��������Y������	��{��`ڕ�J9��`��������Q�����'
���e������l���y��֤�+3��ڐ��屮�M��K������l���̯��,��:���`볼J��@�����vc���������${���  �  ��N=�%N=�vM=��L=�L=fK=�J=fJ=zQI=3�H=��G=�9G=�F=��E=� E=_mD=ݹC=C=RB=��A=��@=63@=}?=�>=P>=�U==�<=��;=)&;=�i:=��9=��8=08=np7=
�6=��5=�,5=Yi4=ۤ3=��2=O2=�M1=S�0=l�/=��.=�.=N:-=�`,=Ӄ+=Q�*=��)=��(=`�'=��&=j&=j
%=U$=�#=��!=�� =7�=�=�=\i=%6=��=��=l==��=�V=F�=�s=0�=�p=��=ZO
=�=�=�h=ڹ=�=�I =w�<���<���<%Q�<>��<���<�<�<�{�<���<���<��<�6�<�X�<sv�<���<+��<��<̼<�ڸ<J�<��<0��<� �<Y�<B�<�	�<Y	�<��<�<��<d��<���<��<�y<�q<��i<��a<�Y<��Q<b�I<��A<t�9<��1<�*<�"<�)<z@<3Z
<6w<0�;z�;���;-�;��;t�;���;�9�;��q;uWS;�	5;�;'��: ��:�w:I�:8[8��ʹj�W�}C��"ܺ��	�K�$���?�QQZ�ret���󜓻N���^�����û��λ'ڻ
��	~�����������_��Hs����������."��Z&�7n*�@i.��L2��6���9�jx=��
A��D�f�G�`K���N���Q�=U�	qX�ܛ[��^�+�a���d���g�s�j�%�m�8�p���s���v�[�y�k�|�D\����e��O僼�I��J������r���ӊ�F5����������nX�����S��y��\ؕ�7������򙼢O��'���P��Rd��@���W���x���դ�3�� ����屮�N��p���n���n���ί��.��e�����eL������4��te���º�z���|���  �  W�N=�%N=RvM=��L=�L=,fK=;�J=�J=�QI=ϟH=i�G=�:G=ևF=��E=�!E=;nD=��C=�C=�RB=4�A=2�@=�3@=R}?=6�>=V>=�U==ۛ<=>�;=�%;=Si:=�9= �8=$/8=�o7=.�6=��5=�+5=wh4=�3=+�2=�2=aM1=�0=-�/=��.=�.=g:-=a,=*�+=��*=��)=`�(=�'=o�&=B&=9%=!$=�#=��!=c� =��=��=L�=�i=S6=�=��=�k=�=
�=�U=��=�r=?�=�o=��=XN
=�=�=�g=�=�=I =K�<ͅ�<"��<�P�<��<���<V=�<B|�<O��<���<��<�8�<iZ�<-x�<1��<��<���<�ͼ<[ܸ<��<��<��<e�<��<u�<�	�<��<C�<A�<� �<��<t��<��<c�y<p�q<�i<�a<G�Y<C�Q<�I<��A<'�9<��1<�*<�"<>)<�@<�Z
<~x<3�;Y~�;��;g3�;Ο�;��;8��;(A�;��q;9fS;15;y�;��:��:h%w:��:I<\8��ʹ��W�G��6)ܺh�	�k�$��?�M\Z�*rt�m��\��������������%�û�λ�ڻ�����ﻊ���Q�������>r�
���M��,"��W&�k*��e.��I2�M6��9�8u=��A�Y�D�&�G�U^K�,�N���Q��<U�qX���[��^���a���d���g�H�j�a�m���p��s��v�ͪy�܇|��_�M������e惼�J������`��Tr���ӊ�5�����������W�������w���֕�]5��q������M���������c��7������#x��Dդ��2�� ����WO��J���r���o��;Я�c0��'���`ﳼN��C����	��'g��ĺ�� ���}���  �  
�N=K%N=2vM=��L=�L=EfK=c�J=	J=RRI=3�H=��G=';G=\�F=Q�E=&"E=�nD=1�C=OC=*SB=��A=��@=�3@=v}?=O�>=[>=zU==��<=��;=d%;=�h:=��9=��8=�.8=o7=��6=U�5=1+5=�g4=��3=��2=P2=
M1=��0=��/=��.=�.=z:-=a,=[�+=�*=޿)=��(=~�'=��&=�&=�%=�$=2#=�!=�� =4�=�=��=�i=g6=�=��=�k=v=��=�U=�=pr=��=/o=�=�M
=A�==`g=d�=j=�H =��<*��<���<fP�<���<���<�=�<�|�<��<���<��<R9�<m[�<:y�<Q��< ��<���<�μ<1ݸ<q�<��<���<��<�<��<p	�<��<��<��<���<L��<���<��<U�y<�q<��i<��a<%�Y<:�Q<C�I<�A<��9<��1<�*< "<�(<�@<5[
<&y<^5�;B��;g��;�6�;ȣ�;M�;�;!F�;t�q;�oS;* 5;��;l �:��:`:w::��\8�ʹ
�W��I��n/ܺ��	� �$���?��bZ��xt�N��ǧ��T��
 �����Ùû�λ�ڻC�����������������q�=	�������|*"�LV&��h*��c.�[G2�6���9�+s=�*A�̇D���G�]K�P�N�V�Q�Q<U�/qX�ߜ[���^���a���d���g���j�I�m���p�7�s�^�v�%�y���|��a�;������4烼`K��z������qr���ӊ��4������j����V��,��� ���v���Օ�P4��T�����L������
��Jb���������w��դ��2��:���>��O��⯫�.���p��ѯ�U1�� �����NO��n����
��h���ĺ��!��S~���  �  �N=9%N=&vM=��L=�L=TfK=r�J=J=dRI=[�H=��G=U;G=��F=}�E=Y"E=�nD=a�C=|C=VSB=��A=��@=�3@=�}?=Z�>=Q>=mU==��<=��;=X%;=�h:=�9=Y�8={.8=�n7=n�6=1�5=�*5=�g4=Z�3=��2='2=�L1=��0=�/=��.=�.={:-=)a,=g�+=�*=��)=��(=��'=�&=�&=�%=�$=U#=1�!=�� =]�=�=��=�i=p6=
�=w�=�k=^=��=�U=��=Cr=w�=�n=��=�M
=�=�=)g=,�=>=rH =b�<���<���<MP�<ާ�<���<�=�<�|�<��<���<��<�9�<�[�<�y�<���<\��<��<ϼ<�ݸ<��<��<���<��< �<��<M	�<��<��<��<���<���<8��<y�<��y<2�q<��i<��a<N�Y<j�Q<��I<]�A<�9<��1<J*<�"<�(<�@<x[
<iy<�5�;���;���;Z8�;Z��;� �;{��;�G�;L�q;�rS;J#5;�;`%�:���:�>w::_]8o�ʹ��W�qK��j1ܺD�	���$�:�?�fZ�|t������o���!������b�ûH�λ�ڻ���d�ﻁ������8��u���q�		�f��r���)"��U&�6h*�c.��F2�K6�S�9�ar=�sA��D�C�G��\K��N�$�Q�H<U�iqX���[��^��a��d�*�g�u�j��m�]�p��s���v�ʭy�׊|�_b����ց��y烼{K����������r���ӊ��4������K����V�������^v��YՕ�4��푘���L��H�������a��^�������w���Ԥ��2��[���R��O������\���p��gѯ��1�������𳼙O��ϭ��U��{h��7ź��!���~���  �  
�N=K%N=2vM=��L=�L=EfK=c�J=	J=RRI=3�H=��G=';G=\�F=Q�E=&"E=�nD=1�C=OC=*SB=��A=��@=�3@=v}?=O�>=[>=zU==��<=��;=d%;=�h:=��9=��8=�.8=o7=��6=U�5=1+5=�g4=��3=��2=P2=
M1=��0=��/=��.=�.=z:-=a,=[�+=�*=޿)=��(=~�'=��&=�&=�%=�$=2#=�!=�� =4�=�=��=�i=h6=�=��=�k=w=��=�U=�=sr=��=3o=�=�M
=F�==fg=k�=q=�H =��<:��<���<vP�<	��<���<�=�<�|�<��<���<��<Y9�<r[�<=y�<R��<���<���<�μ<*ݸ<i�<��<���<��<��<��<c	�<��<��<��<���<C��<���<��<M�y<�q<��i<��a<,�Y<F�Q<R�I<�A<��9<��1<�*<"<)<�@<N[
<>y<�5�;k��;���;�6�;ݣ�;Z�;���;F�;\�q;doS;�5;��;��:K��:�8w:?	:�\8J�ʹ/�W��J���0ܺ.�	���$�?�?�kcZ�syt�����������4 ��3����û#�λ�ڻ[����������������q�A	�������~*"�MV&��h*��c.�\G2�6���9�,s=�*A�̇D���G�]K�P�N�V�Q�Q<U�/qX�ߜ[���^���a���d���g���j�I�m���p�7�s�^�v�%�y���|��a�;������4烼`K��z������qr���ӊ��4������j����V��,��� ���v���Օ�P4��T�����L������
��Jb���������w��դ��2��:���>��O��⯫�.���p��ѯ�U1�� �����NO��n����
��h���ĺ��!��S~���  �  W�N=�%N=RvM=��L=�L=,fK=;�J=�J=�QI=ϟH=i�G=�:G=ևF=��E=�!E=;nD=��C=�C=�RB=4�A=2�@=�3@=R}?=6�>=V>=�U==ۛ<=>�;=�%;=Si:=�9= �8=$/8=�o7=.�6=��5=�+5=wh4=�3=+�2=�2=aM1=�0=-�/=��.=�.=g:-=a,=*�+=��*=��)=`�(=�'=o�&=B&=9%="$=�#=��!=c� =��=��=M�=�i=U6=�=��=�k=�=�=V=��=�r=F�=�o=��=bN
=��=�=�g=��=�="I =i�<��<A��<�P�</��<���<q=�<[|�<e��<��<��<�8�<rZ�<2x�<2��<��<���<�ͼ<Mܸ<��<��<���<N�<��<\�<l	�<��<,�<+�<o �<��<f��<��<T�y<h�q<�i<�a<V�Y<Y�Q<;�I<��A<O�9<+�1<�*<�"<q)<�@<[
<�x<i3�;�~�;U��;�3�;���;��;B��;"A�;��q;�eS;�5;��;��:���:"w:$�:��[8��ʹۖW�(I��Q+ܺs�	�o�$��?�=]Z�st��������1���$������h�ûA�λ�ڻ���'�ﻭ���`�������Hr�
���R��,"��W&�k*��e.��I2�O6��9�:u=��A�Y�D�&�G�V^K�,�N���Q��<U�qX���[��^���a���d���g�H�j�a�m���p��s��v�ͪy�܇|��_�M������e惼�J������`��Tr���ӊ�5�����������W�������w���֕�]5��q������M���������c��7������#x��Dդ��2�� ����WO��J���r���o��;Я�c0��'���`ﳼN��C����	��'g��ĺ�� ���}���  �  ��N=�%N=�vM=��L=�L=fK=�J=fJ=zQI=3�H=��G=�9G=�F=��E=� E=_mD=ݹC=C=RB=��A=��@=63@=}?=�>=P>=�U==�<=��;=)&;=�i:=��9=��8=08=np7=
�6=��5=�,5=Yi4=ۤ3=��2=O2=�M1=S�0=l�/=��.=�.=N:-=�`,=Ӄ+=Q�*=��)=��(=`�'=��&=j&=j
%=U$=�#=��!=�� =8�=�=�=^i='6=��=��=l==��=�V=M�=�s=9�=�p=��=hO
=��=�= i=�=�=�I =��<��<���<PQ�<h��<���<=�<�{�<���<���<��<7�<�X�<{v�<���<(��<��<̼<�ڸ<3�<��<��<� �<7�<�<u	�<7	�<��<��<m�<K��<���<��<��y<�q<��i<��a<�Y<
�Q<��I<��A<��9<=�1<>*<�"<�)<�@<yZ
<yw<�0�;�z�;?��;h-�;E��;��;ɝ�;�9�;O�q;WS;.	5;>�;P��:��:8w:*�:��Z8`�ʹG�W�wF��%ܺ�	���$�5�?��RZ��ft��������������F�L�û��λrڻK��B~����������n��Ts����������."��Z&�;n*�Di.��L2��6���9�kx=��
A��D�g�G�`K���N���Q�=U�	qX�ܛ[��^�+�a���d���g�s�j�%�m�8�p���s���v�[�y�k�|�D\����e��O僼�I��J������r���ӊ�F5����������nX�����S��y��\ؕ�7������򙼢O��'���P��Rd��@���W���x���դ�3�� ����屮�N��p���n���n���ί��.��e�����eL������4��te���º�z���|���  �  ^�N=?&N=�vM=��L=�L=�eK=��J=�J=�PI=f�H=��G=�8G=��F=��E=�E=BlD=ظC=#C=.QB=֜A=�@=�2@=�|?=��>=I>=�U==`�<=	�;=�&;=�j:=��9=��8=18=�q7=2�6=��5=�-5=kj4=Х3=��2=2=�N1=߂0=ʴ/=,�.=�.=>:-=�`,=d�+=��*=C�)=��(=r�'=��&=]&=N	%=:
$=�#=��!=�� =p�=h�=i�= i=�5=�=ݷ=ml=�=;�=jW=B�=�t=[�=
r=�=�P
=X�==>j=�=�=�J =C�<B��<���<�Q�<���<���<�<�<{�<���<���<�<75�<�V�<It�<:��<ؤ�<���<�ɼ<�ظ<s�<�<���<���<��<��<�	�<�	�<d�<�<��<���<���<���<��y<��q<��i<��a<��Y<f�Q<��I<��A<��9<��1<J*<3"<�*<�@<�Y
<�u<T,�;�t�;���;�%�;쐶;�
�;㓗;�/�;=�q;GDS;7�4;��;���: l�:��v:��:��Y8U˹s�W�B���ܺ��	��$���?��EZ�Xt�����
���=�c��Q뷻>�û$�λ~ڻ~��Qzﻇ����� ��޾��t�������72"��^&�;r*��m.��Q2�E6���9�j|=��A�y�D�i H�zbK�f�N� R�x=U��pX��[���^��a��d�x�g���j�X�m���p��s��v���y��|�X�����}���ー�H��L���R���q���ӊ��5��8��������Y������	��{��`ڕ�J9��`��������Q�����'
���e������l���y��֤�+3��ڐ��屮�M��K������l���̯��,��:���`볼J��@�����vc���������${���  �  �N=�&N=wM=�L=L=�eK=�J=7J=�OI=z�H=��G=�7G=��F=��E=ME= kD=��C=�C=#PB=�A=N�@=2@=I|?=��>=?>=�U==��<=��;=t';=uk:=��9=��8=D28=�r7=��6=J�5=/5=�k4=�3=��2=2=NO1=t�0==�/=d�.=�.=:-=5`,=�+=
�*=t�)=��(=Y�'=v�&= &=%=�$=�#=��!=�� =��=��=ē=�h=�5=��=�=�l==��=WX=X�=v=��=~s=��=RR
=�=�=�k=v�==�K =�<���<��<�R�<���<���</<�<)z�<:��<���<�<�2�<YT�<�q�<���<=��<��<_Ǽ<yָ<n�<W�<X��<���<��<��<�	�<

�<I	�<F�<e�<� �< ��<#��<��y<c�q<^�i<S�a<K�Y<��Q<{�I<��A<��9<��1<�*<�"<N+<�@<�X
<ft<'�;en�;ο�;��;f��;K��;���;�#�;w�q;�,S;2�4;��;���:6M�:��v:��:�W8$4˹�W�g=���ܺh�	���$��?�~5Z�\Ft�K�8���j査���ⷻ.�ûw�λ��ٻ���1v�k���n��������u�������36"�nc&�aw*��r.��V2��$6��9���=�@A�x�D��H�neK�}�N�aR�?>U��pX�O�[��^���a�
�d���g���j���m��p���s���v�c�y��z|�)S�����{��	⃼+G��9������gq���ӊ��5�������9[��c�����_}���ܕ��;�����v���ST������T���g��Cà����~z���֤�h3�������M�����p��k���ʯ�G*�������購gG������{���`��t������xy���  �  ��N=:'N=^wM=&�L=mL=3eK=��J=�J=)OI=m�H=��G=~6G=P�F=#�E=�E=�iD=6�C=�C=�NB=�A=��@=o1@=�{?=e�>=;>=V==	�<=�;=)(;=bl:=��9=
�8=�38=1t7=�6=��5=w05=�l4=G�3=��2=2=#P1=�0=��/=��.=�.=�9-=�_,=Z�+=M�*=��)=��(=2�'=5�&=� &=�%=�$=E#=Y�!=�� =s�=Ͷ=�=h=q5=��=8�="m=�=��=TY=��=_w=8�=u=B�=�S
=��=>=Dm=�=a=M =�<C��<,��<]S�<Y��<t��<�;�<y�<��<:��<�
�<�0�<�Q�<o�<���<\��<=��<�ļ<Ը< �<w�<���<M��<�<-�<�	�<
�<"
�<�<"�<��<X��<���<`�y<[�q<W�i<d�a<"�Y<L�Q<��I<R�A<��9<��1<�
*<1"<#,<�@<�W
<cr<X!�;}g�;���;��;�{�;��;b|�;�;m�q;KS;��4;ݯ;א�:�,�:�iv:�i:��U8�P˹U�W��8���ܺՕ	���$�Ŭ?��$Z��3t�Kꆻ΀���۟�/���5ط��vû4�λ�ٻ����qﻐ�������������w��A������:"�;h&��|*�[x.��\2�T*6���9�ֆ=� A��D��H�whK��N�
R�?U��pX�}�[�}�^���a���d��g�k�j���m���p�=�s��v���y�Du|��M����y��*����E��$������q���ӊ�6��՘������\��R���g������ߕ��>��眘�H���W���������i���Ġ�< ���{��bפ��3��s���L��ͪ���	��i��tȯ��'������峼�D��â��� ��s^��!�������w���  �  [�N=�'N=�wM=4�L=HL=�dK=�J=� J=BNI=f�H=]�G=75G=��F=��E=rE=1hD=ߴC=|C=�MB=�A=��@=�0@=^{?="�>=>=6V==g�<=��;=�(;=Am:=��9=5�8=�48=�u7=]�6=%�5=�15=Pn4=v�3=�2=�2=�P1=��0=�/=��.=�.=�9-=x_,=Ё+=��*=��)=��(= �'=��&=m�%=G%=3$=�#=�!=m� =s�=�=l�=�g=,5=��=O�=~m=B=��=GZ=��=�x=��=�v=��=�U
=>�=�=�n=U�=�	=/N =��<ӌ�<W��<	T�<���<H��< ;�<!x�<e��<i��<��<?.�<O�<2l�<̅�<x��<k��<¼<�Ѹ<�޴<z�<,��< ��<A�<��<�	�<�<	�<�	�<��<��<��<G��<��y<<�q<��i<c�a<��Y<��Q<��I<��A<f�9<(2<d*<�"<�,<)@<�V
<up<��;`�;Y��;��;�p�;��;�o�;�
�;�rq;��R;f�4;l�;j�:+
�: 4v:�?:��S8�x˹V�W�83����ۺ��	�8�$���?�%Z��!t�\���ev��<џ��Tη�nû��λm�ٻ(��Cmﻂ������3��y��Zy�e�f�����&?"�5m&��*�~.�Wb2�06�9�9�"�=��A�i�D�eH��kK�9�N��R��?U��pX���[�ҷ^��a���d�I�g���j���m�~�p���s�.�v��y��o|��H����Ow��`ރ�5D��������p�� Ԋ��6������<���w^��M����!��B���J╼hA����������Y������
��l���Ơ��!���|��ؤ��3��e���w�&K��m�����g��!Ư�R%��V���㳼�A��������� \��͹�����	v���  �  �N=(N=�wM=J�L=,L=�dK=��J=1 J=kMI=u�H=A�G=�3G=��F=c�E=E=�fD=��C=B C=�LB=�A=��@=50@=�z?=��>=>=XV==��<=�;=�);=n:=��9=N�8=68=�v7=��6=v�5=35=�o4=��3=!�2=�2=�Q1=E�0=u�/=�.=�.=�9-=_,=H�+=ݟ*=ź)=��(=��'=��&=,�%=�%=�$=� #=��!=L� =��=�=Ƒ=+g=�4=��=o�=�m=�=6�=1[=��=�y=��=x=X�=0W
=��=Y=Ep=��=�
=5O =��<(��<T��<�T�<���<��<X:�<-w�<��<���<��<�+�<�L�<�i�<��<���<ɭ�<���<ϸ<�ܴ<��<��<���<~�<]�<�	�<g�<��<�<F	�<��<��<� �<h�y<��q<"�i<��a<��Y<��Q<^�I< �A<��9<2<J*<!"<9-<�?<�U
<|n<��;
Y�;g��;E��;&f�;�ܦ;>d�;���;P[q;�R;М4;W�;FF�:2�:� v:�:@$R8��˹P�W�]/���ۺ+�	�Ϲ$���?��Z��t��ֆ��l��wǟ�~嫻�ķ�aeû�λ��ٻ���4i����Q��X��T��{���c��Z��0C"��q&���*�7�.��g2�p56�s�9� �=��!A�q�D�H��nK�t�N�@R��@U��pX��[�w�^���a���d���g���j�X�m�\�p���s���v��y��j|��C����du���܃��B��������pp��Ԋ�n7������h���`��!��#�������䕼D��a�������R\�����N���m���Ƞ��"���}���ؤ�.4��I����쨼fJ��1������9e��	į��"�������೼
?��p���}����Y���������~t���  �  ��N=�(N=$xM=V�L=L=SdK=&�J=��I=�LI=��H=R�G=�2G=�F==�E=�E=�eD=��C=I�B=�KB=0�A=*�@=�/@=z?=��>=�>=gV==�<=�;=#*;=�n:=v�9=<�8=78=�w7=Ƿ6=��5=545=�p4=��3=��2=�2=MR1=��0=̶/=9�.=�.=o9-=�^,=ɀ+=>�*=�)=��(=��'=��&=�%=�%=�$=��"=��!=g� =��=f�=5�=�f=�4=��=��=n=0=п=�[=��=�z=�=@y=��=�X
=�=�=pq=��=�=P =I�<[��<)��<U�<��<���<�9�<?v�<٫�<8��<�<*�<�J�<Kg�<À�<c��<���<a��<$͸< ۴<�<a�<���<� �<�<�	�<��<w�<	�<�
�<e�<��<��<��y<G�q<�i<��a< �Y<%�Q<P�I<��A<��9<�2</*<-"<�-<�?<�T
<�l<��;S�;
��;E��;s]�;Ӧ;%Z�;[�;�Fq;_�R;Ȋ4;u;W&�:Eϵ:��u:�� :2�P8��˹��W�,����ۺb}	��$�c�?�d�Y��t�'φ��d��⾟�Gݫ����/^û��λI�ٻ����e��������s����i|���������F"��u&�7�*�Ǉ.�nl2�!:6��9�h�=��%A��D�)H�+qK���N��R�[AU��pX�}�[�B�^��a�e�d���g�u�j���m�c�p�X�s�b�v�W�y�hf|��?��
���s��Iۃ��A��1������Pp��/Ԋ��7��Y�������Ya���Ñ��%�������敼QF���������^��)���.���o���ɠ�,$���~��@٤�n4��6����쨼�I��/���4���c��F¯�!�����Z޳��<��0���j����W��⵺�X��s���  �  ��N=�(N=MxM=`�L=�L=dK=ڱJ='�I=1LI=�H=��G= 2G=�~F=a�E=E=�dD=��C=r�B=KB=��A=��@=8/@==z?=s�>=�>=zV==#�<=��;=�*;=Mo:=�9=��8=�78=�x7=��6=m�5=55=kq4=\�3=��2=02=�R1=�0=�/=X�.=�.=G9-=�^,=o�+=ɞ*=z�)=K�(=)�'=��&=<�%=%=�$=��"=�!=�� =�=�=ɐ=jf=z4=��=��=Dn=�=D�=�\=I�=�{=��=.z=��={Y
=�=�=]r=��=�=�P =S�<J��<���<�U�<��<���<u9�<�u�<���<��<��<h(�<�H�<�e�<�<���<���<���<�˸<�ٴ<��<d�<:��<P �<��<�	�<��<
�<��<��<�	�<5�<e�<$z<��q<z�i<@�a<��Y<��Q<��I<6�A<7 :<+2<�*<�"<�-<\?<�S
<�k<0�;�N�;���;���;V�;�˦;�R�;��;�7q;��R;x{4;=g;��:8��:�u:�� :0JO8��˹4�W��(����ۺ�x	��$��|?���Y��s��Ȇ�H^��ʸ���֫����UXû]�λ�ٻ���Gc��������������b}�\��������I"�y&���*�C�.��o2��=6�}�9��=��(A��D�tH�sK��N��R�BU�qX�
�[�9�^���a���d���g���j�z�m�8�p�޹s��v� �y��b|��<�.	��nr��5ڃ��@��������!p��AԊ�C8��؛��V���Xb���đ�'��E����蕼H��r������E`��⻜����q��
ˠ�%��.���٤��4��)���Z쨼I��z���?��vb������p��~���ܳ�;��|�������V��j���"��r���  �  &�N=�(N=fxM=i�L=�L=�cK=��J=��I=�KI=��H=#�G=�1G=8~F=��E=~E=NdD=-�C=��B=�JB=-�A=L�@=�.@=z?=Y�>=�>=�V===�<=�;=�*;=�o:=|�9=`�8=N88=Fy7=*�6=��5=�55=�q4=Ƭ3=�2=�2=S1=U�0=4�/=p�.=�.=89-=k^,=0�+=z�*=�)=��(=��'=b�&=��%=q%=`$=:�"=��!=1� =��=��=��=1f=Y4=��=��=hn=�=��=�\=��=5|=w�=�z=;�=Z
=��=8=�r=)�=+=8Q =�<ϐ�<-��<�U�<��<���< 9�<u�<R��<Z��<��<y'�<�G�<vd�<�}�<r��<���<���<�ʸ<�ش<�<��<���< �<��<�	�<#�<R�<E�<H�<g
�<�<O�<Rz<$ r<��i<��a<��Y<x�Q<<�I<��A<�:<^	2<Z*<t"<.</?<?S
<�j<��;�K�;3��;��;R�;Ǧ;zM�;w�;X-q;ƸR;�r4;�_;���:G��:�u:�� :�N8�˹�W��'����ۺ�t	�*�$��v?���Y�
�s��Ć�0Z�������ҫ�7���?Uûr�λ0�ٻP�今a�����R�����%��~�l�B��s�RK"��z&���*�o�.�Ir2��?6���9�Κ=��*A���D�H�dtK�#�N�8	R�YBU�qX���[���^���a�t�d�)�g�-�j���m�.�p�Ƿs�۟v�˂y��`|��:�c���q���ك�>@�����R���o��UԊ�r8��C�������
c���ő��'��9����镼%I���������Ka��м������q���ˠ��%������٤��4�����'쨼�H����������a��	������}���۳��9��k�������,U������\��pq���  �  ��N=�!N=pM=4�L=�L=;YK=�J=��I=�>I=׊H=��G=@"G=�mF=X�E=�E=9PD=��C=��B=�1B=F|A=��@=4@=:Y?=��>=�==�/==su<=4�;=��:=�@:={�9=<�8=�8=qA7=�~6=�5=��4=�/4=ig3=��2=��1=61=D40=�a/=̌.=�-=�,=��+=z+=�5*=�L)=g`(=�o'=3{&=*�%=�$= �#=iz"=`m!=�Z =�A=�"=��= �=�=o`==��=�~=J#=�=�T=7�=f=M�=�X=l�	=�.=h�=��=9==ފ=m��<*�<	��<��<z�<]��<,�<�x�<$��<���<�4�<�g�<a��<���<���<��<-$�<�?�<DY�<Qp�<A��<+��<5��<Q��<�Ť<�Ѡ<�ۜ<u�<��<"�<d��<���< �<��<�z<#r<�j<�'b<]2Z<n>R<ZLJ<\B<n:<V�2<��*<�"<��<��<<�4<ž�;A�;��;k��;"��;!�;���;?w�;3�v;�SX;K:;�t;4��:S��:_�:��:i�'9��V�8�5;���w˺�������6��P���j�k������Ԛ��㦻ն���N���ɻ��Ի?�߻O껡���:����k�5H	�;�U���4�ۢ�c���0$��Q(��Z,��L0��(4�3�7�ʡ;�sA?�X�B�DMF���I��M��pP�9�S� �V�C+Z�V]��x`�Q�c�c�f�K�i�|�l�:�o�\�r�5�u��x��x{��\~�W������Cy���䄼�N��㷇�| ��M����vV������~"��ˇ��2쒼�O��ײ������u���ՙ��4��e����WN��H������d������W��!}��Lۨ��9���������<X��"���@��gx���س��8��;���Z����Y��<�����O|���  �  ��N=�!N=pM=<�L=�L=9YK=%�J=��I=�>I=�H=��G=l"G=�mF=��E=�E=cPD=��C=��B=�1B=b|A=��@=:@=FY?=��>=�==�/==eu<=%�;=��:=�@:=`�9=�8=�8=NA7=�~6=�5=��4=P/4=;g3=~�2=��1=11=840=�a/=ʌ.=��-=�,=��+=�+=�5*=�L)=y`(=p'=^{&=P�%=��$=*�#=�z"=�m!=�Z =�A=�"=�='�=�=f`==��=�~=9#=޿=oT=�=�e=�=�X=<�	=�.=>�=F�===��=>��<�)�<ݣ�<��<z�<]��<�+�<�x�<"��<���< 5�<�g�<���<��<3��<��<�$�<Q@�<�Y�<�p�<q��<T��<K��<u��<�Ť<�Ѡ<�ۜ<n�<��<�<_��<���<���<n�<4z<�r<�j<'b<�1Z<�=R<�KJ<�[B<�m:<�2<��*<ر"<��<��<<"5<��;��;���;y��;���;x�;��;�x�;&�v;�VX;XN:;�v;���:���:�`�:�:ȼ'9Pꏹ��8��;��`x˺�������6��P�#�j�S������֚��䦻G���	P���ɻ�ԻK�߻SO����<����k�:H	�����4�����0$�*Q(�VZ,�KL0�	(4���7��;��@?��B��LF���I��M��pP�P�S��V�D+Z�NV]��x`�d�c���f�Ųi�/�l��o�دr�բu���x�.y{�]]~��������_y���䄼�N�����s ��>����[V������k"�������뒼�O�����g��hu��uՙ��4�������.N��&������d������T��}��[ۨ�:���������jX��f�������x��ٳ�19��{�������Z������K��Y|���  �  }�N=s!N=pM=5�L=�L=QYK=T�J=��I=<?I=>�H=�G=�"G=XnF=�E=`E=�PD=�C=<�B=2B=�|A=��@=q@=tY?=��>=�==�/==Ou<= �;=��:=b@:=�9=��8=`8=�@7=P~6=��5=x�4=�.4=�f3=5�2=��1=�1=40=�a/=��.=�-=�,=�+=�+=�5*=@M)=�`(=\p'=�{&=��%=�$=��#=�z"=�m!=![ =HB= #=6�=R�=-�=l`=	=��=b~=�"=��=T=��=�e=��=[X=��	=&.=Ў=��=�<=[�=~��<:)�<f��<k�<�y�<F��<,�<y�<y��<4��<�5�<�h�<b��<���<���<��<T%�<A�<dZ�<Tq�<��<���<ҩ�<渨<!Ƥ<�Ѡ<�ۜ<T�<��<��<���<7��<7��<��<�z<r<)j<e%b<0Z<8<R<jJJ<NZB<�l:<��2<�*<n�"<��<��<O<�5<���; �;+��;=�;���;��;�;X|�;	�v;_]X;'U:;�|;��:���:j�:@�:��'9_ޏ���8�s<���z˺����c�6���P�̱j����ǐ��ٚ�E离Ӻ��=R����ɻJ�Ի<�߻�P껮��������k��G	�x�G���3�1������.$��O(��X,��J0�_&4��7���;�e??���B��KF���I��M�pP��S�	�V�|+Z��V]��y`�o�c�ܧf��i�b�l�r�o�7�r�t�u�#�x��z{��^~�A���d���y�� 儼O��5���� ��5���zV��E����!������`뒼�N��Ʊ������t���ԙ��3��S���-𝼎M����������d������B��}���ۨ�B:����������X������=��|y���ٳ�:��;���i����Z���������|���  �  9�N=;!N=�oM=&�L=L=�YK=��J=?�I=�?I=��H=��G=e#G=oF=��E=	E=oQD=��C=��B=�2B='}A=8�@=�@=�Y?=ԡ>='�==�/==2u<=Ĺ;=f�:=@:=��9=4�8=�8=I@7=�}6=�5=��4=[.4=Tf3=��2=)�1=�1=�30=�a/=��.=�-=:�,=A�+=�+=*6*=�M)=Na(=�p'=W|&=V�%=��$=3�#=�{"=�n!=�[ =�B=}#=��=��=D�=�`=�=��=&~=�"=!�=�S=�=�d=��=�W=�	=c-=�=!�=�;=��=���<m(�<���<��<�y�<��<9,�<9y�<���<���<y6�<�i�<{��<���<G��<�<�&�<wB�<�[�<�r�<7��<ԙ�<���<n��<�Ƥ<Ҡ<�ۜ<1�<@�<%�<$��<b��<��<��<
z<Jr<�j<�"b<T-Z<�9R<�GJ<\XB<�j:<�2<��*<ΰ"<I�< �<�<�6<`��;##�;E��;��;㋸;y!�;Sș;3��;�v;�iX;`:;W�;���:%��:�w�:��:)0(94̏���8��<��]˺�F���6��P�<�j����t����ݚ�P즻>����V��Ѱɻ+�Ի��߻zR�ӹ������k�AG	�����+2�������L,$�M(�V,��G0��#4�U�7�
�;�=?���B��IF��I��M�loP�_�S��V��+Z�NW]��z`���c�k�f���i���l�Һo��r���u���x�F}{� a~�p���\���z���儼�O��t���� ��/����U������*!�����F꒼�M��s���N��Ds��Uә��2������L��ʩ�����d��`�����3}���ۨ��:����������Y�����o���z��۳�E;�����������[��6�������}���  �  ��N=� N=�oM= �L=L=�YK=٦J=��I=$@I=a�H=U�G=$G=�oF=h�E=�E=GRD=��C=��B=Z3B=�}A=��@=2@=�Y?=��>=/�==�/== u<=j�;=��:=t?:=�9=��8=8=�?7=�|6=�5=��4=�-4=�e3=�2=��1=1=d30=Ba/=��.=�-=S�,={�+=Y+=�6*=2N)=�a(=�q'=}&="�%=��$=�#=\|"=9o!=R\ =iC=$=��=��=p�=�`=�=^�=�}=+"=��=�R=T�=�c=�=�V=�	=k,=�=<�=;=��=��<@'�<���<E�<1y�<���<P,�<�y�<���<���<�7�<�j�<ۘ�<u��<���<�	�<i(�< D�<9]�<�s�<���<��<���<3��<Ǥ<@Ҡ<�ۜ<�<��<m�<��<)��<���<
 �<�z<�r<�j<	b<�)Z<k6R<�DJ<�UB<~h:<�}2<n�*<�"<�<�<�<�7<��;'�;���;��; ��;n(�;�ϙ;���;N�v;xX;lm:;��;8��:'��:)��:9:|(9�m�8�?����˺}�j�Ƭ6���P���j�1��^����㚻]��Ĳ��[����ɻs�Ի!�߻U�ʻ��q����k��F	������0�2�����p)$�	J(��R,��D0�< 4��7���;�J:?���B��GF��I��M�inP��S��V�,Z�]X]�|`���c���f���i���l�ܽo�4�r�?�u��x�r�{�d~�١������{���愼MP��⸇�� ��&����)U��κ��$ ��ل���蒼[L��㮕�����q���љ��0�������흼<K���������bc���������<}���ۨ�F;��Ӛ������
[��j������E|���ܳ��<��2���:���`]����������~���  �  [�N=� N=�oM=�L=2L=�YK=;�J=*�I=�@I=�H=*�G=%G=�pF=e�E=�E=@SD=s�C=y�B=#4B=y~A=T�@=�@=IZ?=.�>=@�==t/==�t<=�;=v�:=�>:=J�9=��8= 8=�>7=�{6=�5=�4=�,4=�d3=D�2=��1=�1= 30=�`/=Z�.=�-=p�,=��+=�+= 7*=�N)=�b(={r'= ~&=�%=��$= �#=I}"=p!=2] =D=�$=h�=.�=��=�`=�=�=b}=�!=ܽ=R=l�=�b=��=�U=��	=?+=�=�=:=�=t��<�%�<���<m�<�x�<���<k,�<z�<F��<���<�8�<Dl�<���<J��<���<��<n*�<F�<1_�<�u�<��<l��<���<��<�Ǥ<�Ҡ<�ۜ<��<(�<��<��<���<$��<7��<�z<�	r<�j<�b<�%Z<�2R<~AJ<wRB<�e:<�{2<��*<Ѯ"<�<N�<t<D9<���;�,�;���;��;B��;�0�;vؙ;���;��v;7�X;�~:;z�;T��:�:���:H<:��(9���Ի8��B��c�˺��r�~�6���P���j�
!��|���+뚻 ���
̲�4b��9�ɻm�Ի'�߻�W껢�������|k�F	�U���.�^������%$�2F(��N,�t@0�/4��7�-�;��6?���B��DF��I�mM�mP�^�S��V��,Z�qY]�|}`�c�\�f���i���l���o��r�W�u��x�1�{��g~�t�����}���焼�P��l���!�����xmT��������s���^璼zJ���������o���ϙ�/�������라�I��g�������b��t������Y}��dܨ��;������ ���n\���������3~���޳��>�����(���,_��!���^������  �  ��N=@ N=IoM= �L=IL=#ZK=��J=��I=sAI=׍H=�G=&G=�qF=v�E=�E=TTD=s�C=f�B=�4B=8A=��@=@=�Z?=[�>=R�==[/==t<=��;=��:=5>:=v9=ӿ8=*�7=�=7=�z6=��5=�4=�+4=�c3=b�2=3�1=�1=20=�`/=(�.=�-=��,=�+='+=�7*=�O)=qc(=[s'=�~&=�%=��$= �#=O~"=q!=^ =�D=L%=��=��=�=�`=�=��=�|=!="�==Q=c�=�a=��=JT=��	=*=��=��=9=
�=О�<f$�<���<��<x�<���<~,�<�z�<��<� �<5:�<�m�<n��<:��<��<��<�,�<>H�<*a�<�w�<ȋ�<ꝰ<ڭ�<��<EȤ<�Ҡ<�ۜ<C�<��<��<��<=��<S��<S��<��y<�r<$j<�b<p!Z<|.R<�=J<OB<	c:<2y2<5�*<��"<�<~�<.<�:<���;N2�;���;Q�;d��;�9�;��;��;7�v;~�X;
�:;t�;v�:%,�:���:�]:�*)9�}���8�F��̔˺k �c���6�"Q�b�j�r(�����󚻶 ��pӲ��h����ɻ��Իe�߻u[껾�������Ek�}E	�"�����+�w�����"$�NB(��J,�6<0��4���7�D�;��2?���B��AF���I��M��kP�ӶS���V�o-Z��Z]�g`��c��f��i�~�l���o���r���u��x�N�{��k~�:������f~���脼�Q��򹇼J!��퇊�'�S�������������咼�H��
������{m���͙��,��׋��3ꝼFH���������a��������f}���ܨ��<��˜��/����]������x��6����೼A��*���-��a������� ������  �  P�N=�N=oM=�L=XL=`ZK= �J=7�I=BI=��H=��G=�&G=�rF=��E= 
E=[UD=t�C=N�B=�5B=�A=��@=�@=�Z?=��>=V�==@/==@t<=F�;=]�:=�=:=�~9=�8=8�7=|<7=�y6=�5=��4=�*4=�b3=��2=x�1=U1=20=X`/= �.=ִ-=��,=O�+=�+=B8*=0P)=Hd(=9t'=�&=�%=��$=�#=M"=�q!=�^ =�E=�%=q�=��=�=�`=�=��=�|=s =`�=]P=k�=�`=��=	S=_�	=�(=}�=��=�7=�=��<�"�<S��<��<�w�<U��<�,�<�z�<���<��<~;�<|o�<)��<1��<��<�<�.�<VJ�< c�<�y�<���<@��<��<켨<�Ȥ<Ӡ<�ۜ<��<��<��<x�<��<���<d��<k�y<� r<�j<�b<Z<e*R<�9J<�KB<`:<�v2<`�*<��"<��<��<	<E<<@��;R7�;���;�!�;g��;pB�;�;���;��v;֭X;��:;)�;1�:@D�:�ǈ:c}:3�)9�g��W�8�1I���˺�&�w'�f�6�{Q���j�0��豎���������ڲ��o����ɻ��Ի��߻�^���������Uk��D	�����8)�Ȕ���w$�[>(�cF,��70��4���7�L�;�\/?�)�B�:?F�G�I��M��jP�(�S�	�V��-Z��[]�D�`���c��f�:�i��l���o�H�r���u�P�x���{��o~����S������鄼�R��v����!�������틼"S�������������㒼�F��
���{
��Xk��q˙��*������k蝼�F��̤����� a������T���}��0ݨ�F=��Ɲ�����n_��o���U!��:����⳼/C��O���7���b���º�o"��o����  �  ��N=|N=�nM=ֽL=nL=�ZK=M�J=��I=�BI=V�H=��G=�'G=�sF=u�E=E=JVD=l�C=-�B=�6B=��A=%�@=@=B[?=Ȣ>=a�==%/==�s<=�;=��:=�<:=�}9=�8=F�7=�;7=�x6=��5=��4=�)4=b3=И2=��1=� 1=�10=�_/=֋.=ʴ-=��,=��+=�+=�8*=�P)= e(=u'=π&=�%=��$=�#=0�"=�r!=�_ =UF=~&=��=8�=C�=�`=j=H�=|=�=��=�O=��=�_=~�=�Q=3�	=�'=\�=��=�6=/�=b��<�!�<H��<��<w�<!��<�,�<P{�<���<��<�<�<�p�<ϟ�<��<���<�<�0�<ML�<e�</{�<
��<���<0��<���<wɤ<jӠ<�ۜ<��<�<��<C��<N�<���<o��<{�y<��q<�j<�b<�Z<L&R<46J<�HB<?]:<�t2<��*<~�"<
�<��<�<r=<D��;`<�;���;�(�;=��;�J�;s�;���;��v;i�X;!�:;��;�K�:�[�:pڈ:T�:��)9�O��;�8��M��-�˺�,�R0��6��Q���j�	7��A���������᲻�v��i�ɻ�Ի�߻�a�~�������\k�D	�� ����'�����)$�~:(��B,��30��4���7�p�;�,?�&�B��<F� �I�=M��iP�~�S� �V��.Z�(]]�ɂ`���c���f�0�i���l�H�o�$�r���u�R�x�Y�{�Gs~�˨�����&����ꄼqS������!��懊�\틼�R��8���q��4��kⒼ$E��������Oi���ə�	)������杼7E���������b`�� ������}���ݨ�>�����������`��¯�9#������䳼'E��G������d��Gĺ��#�������  �  j�N=.N=�nM=ǽL=uL=�ZK=��J=�I=2CI=�H=c�G=�(G=�tF=G�E=�E=WD=1�C=��B=M7B=>�A=��@=p@=�[?=�>=e�==/==�s<=��;=j�:=O<:=R}9=`�8=��7=�:7=�w6=�5=#�4=�(4=La3=�2=(�1=D 1=410=�_/=��.=ƴ-=��,=��+=D+=69*=`Q)=�e(=�u'=��&=Ɉ%=M�$=̈#=��"=�s!=T` =�F='=P =��=q�=�`=S=�=�{=m=�=�N=��=�^=��=�P=2�	=�&=g�=��=
6=b�=���<h �<K��<1�<�v�<���<�,�<�{�<��<��<�=�<+r�<6��<���<���<��<^2�<�M�<�f�<�|�<Y��<ġ�<��<f��<�ɤ<�Ӡ<�ۜ<S�<��<��<6�<�<��<���<&�y<H�q<� j<
b<�Z<*#R<*3J<�EB<�Z:<�r2<0�*<��"<��<��<|<�><���;�@�;ȱ�;z.�;���;�Q�;���;���;�w;��X;��:;e�;*c�:�o�:[�:��:�#*9?���8��P����˺�2��7�0�6��%Q�5k��<������u��)���粻�{����ɻ��Ի��߻�d�N�������Hk��C	������&%�Ə����?$�u7(�\?,��00�J4���7�c�;�)?���B�F:F�?�I��M��hP�<�S��V�/Z�*^]�e�`���c��f���i���l�W�o�o�r�#�u���x���{�Iv~�0�����D����넼.T�������!��ᇊ�,틼�Q��z���t��~��ᒼ�C����������g���Ǚ�y'������t坼�C��w���� ���_���������}���ݨ��>������� ��b��jï��$������z泼�F���������:f���ź�%�������  �  �N=�N=}nM=��L=�L=�ZK=ڨJ=^�I=�CI=b�H=��G=+)G=0uF=��E=yE=�WD=ϢC=��B=�7B=��A=��@=�@=�[?=��>=o�==�.==�s<=P�;=�:=�;:=�|9=Ѽ8=��7=	:7=Cw6=n�5=u�4=F(4=�`3=��2=��1=��0=�00=�_/=��.=Ŵ-=��,=��+=�+=9*=�Q)=f(=Jv'=�&=s�%=�$=h�#=��"=-t!=�` =dG=Z'=� =��=��=�`=E=��=~{==��=NN=�=;^=��='P=n�	=�%=��=�=_5=��=��<~�<���<��<9v�<���<�,�<�{�<���<@�<�>�<.s�<^��<���<���<�<�3�<AO�<�g�<�}�<O��<���<���<쾨<.ʤ<�Ӡ<�ۜ<��<7�<3�<u�<�<_�<���<Y�y<w�q<�i<Jb<�Z<� R<�0J<�CB<5Y:<?q2<=�*<��"<H�<��<�<�?<���;�C�;��;S3�;���;7W�;{ �;���;�w;��X;��:;��;Ls�:�}�:���:��:!R*9<.���8��S���˺7��<��6��-Q�Pk��A��pĎ�d��A��{첻?�����ɻ��Ի}�߻�f�T�������5k�dC	������#�0�����$�5(��<,�.0��	4���7� �;��&?���B��8F���I��M�	hP��S��V��/Z��^]���`��c���f��i���l���o�*�r���u�^�x�[�{��x~�N���'������센�T��׻��8"��ч���싼�Q���������7}������B��]������ef���ƙ�*&��t���L䝼C������o ��<_��i�������}��Oި��>��*���|�� c���į��%��
����糼8H��L�����ng���ƺ�&��z����  �  ��N=�N=hnM=��L=�L=�ZK=��J=��I=�CI=��H=?�G=�)G=�uF=P�E=�E=%XD=+�C=��B=!8B=�A=F�@=�@=�[?=�>=u�==�.==zs<=�;=��:=�;:=}|9=z�8=��7=�97=�v6=�5=�4=�'4=^`3=C�2=i�1=��0=�00=d_/=p�.=��-=��,=�+=�+=�9*=
R)=af(=�v'=t�&=ɉ%=P�$=̉#=�"=�t!=+a =�G=�'=� =��=��=�`=:=��=J{=�=X�=�M=��=�]=j�=�O=��	=]%=.�=��=�4=`�=E��<��<��<Y�<	v�<���<�,�<|�<���<��<?�<�s�<���<~��<���<��<{4�<�O�<�h�<u~�<鑴<.��<7��<:��<\ʤ<�Ӡ<�ۜ<��<��<��<��<i��<��<��<��y<��q<J�i<�b<Z<�R<[/J<BBB<�W:<Cp2<p�*<G�"<&�<�<1<0@<���;WF�;���;�5�;���;lZ�;��;9��;w;S�X;��:;�;c~�:���:���:s�:�p*9@%����8�4V���˺F:��@���6��2Q��k��D��uǎ�z����3ﲻ���� �ɻ3�Իf�߻}h껒���?���8k�,C	����`���"����Q���$��3(�2;,�b,0�4��7���;��%?�e�B��7F��I�M��gP���S��V��/Z�^_]�`�`�
�c���f�N�i�V�l�^�o���r�j�u���x�ɗ{�?z~� ����������턼U�����R"��Ǉ���싼nQ������>���|��zߒ��A����������e���ř�r%��Ǆ���㝼�B��$��������^��A�������}��wި�U?������
���c��&ů��&�������購	I��������)h��jǺ��&������  �  ��N=�N=knM=��L=�L=�ZK=
�J=��I=�CI=ŐH=c�G=�)G=�uF=q�E=E=DXD=Z�C=��B=C8B=	�A=K�@=�@=�[?=�>=l�==�.==vs<=�;=��:=�;:=i|9=W�8=a�7=�97=�v6=ܲ5=��4=�'4=3`3=+�2=N�1=��0=�00=U_/=v�.=��-=��,=�+=�+=�9*=R)=}f(=�v'=��&=�%=u�$=�#=�"=�t!=Va =�G=�'=� =��=��=�`=0=��=9{=�=L�=�M=��=�]=9�=�O=Ž	=.%=�=u�=�4=I�=��<��<���<C�<	v�<���<�,�<<|�<���<��<E?�<�s�<T��<���<���<1�<�4�<IP�<�h�<�~�<��<A��<J��<X��<uʤ<�Ӡ<�ۜ<��<��<��<��<0��<s�<��<!�y<&�q<��i<�b<kZ<AR<�.J<�AB<�W:<(p2<6�*<U�"<�<��<]<n@<��;�F�;ٸ�;7�;(¸;�[�;��;���;Cw;�X;��:;Z�;���:��:C �:��:�z*9�(��W�8��V��j�˺�:��A��6��4Q�Jk��E���Ȏ����Q����D�����ɻ�Ի��߻�h��������Rk�7C	�h��)���"��������$��2(��:,��+0�{4��7�;��$?��B�=7F�٩I��M�ZgP���S�.�V��/Z��_]���`�-�c�i�f���i���l��o�B�r��u���x�f�{��z~�K������Ӄ��턼0U��'���M"��؇���싼NQ��w���6��x|��9ߒ��A��D������Be���ř�(%��j���k㝼MB����������^��&�������}��jި�o?������$���c��dů��&������購_I��g���	���h���Ǻ��&��,����  �  ��N=�N=hnM=��L=�L=�ZK=��J=��I=�CI=��H=?�G=�)G=�uF=P�E=�E=%XD=+�C=��B=!8B=�A=F�@=�@=�[?=�>=u�==�.==zs<=�;=��:=�;:=}|9=z�8=��7=�97=�v6=�5=�4=�'4=^`3=C�2=i�1=��0=�00=d_/=p�.=��-=��,=�+=�+=�9*=
R)=af(=�v'=t�&=ɉ%=P�$=̉#=�"=�t!=+a =�G=�'=� =��=��=�`=;=��=K{=�=Z�=�M=��=�]=n�=�O=��	=b%=3�=��=�4=e�=Q��<��<%��<e�<v�<���<�,�<)|�<���<��<'?�<�s�<���<���<���<��<z4�<�O�<~h�<p~�<㑴<'��<.��<1��<Rʤ<�Ӡ<�ۜ<��<��<��<��<b��<��<��<��y<��q<J�i<�b<Z<R<f/J<OBB<X:<Tp2<��*<Z�"<9�<'�<D<B@<���;uF�;��;�5�;���;vZ�;��;6��;w;4�X;Y�:;��;�}�:��:���:�:�j*9k(��S�8�W����˺�:�QA�Y�6�3Q��k��D���ǎ����/��Rﲻ����ɻI�Իy�߻�h껠���L���=k�0C	����c���"����S���$��3(�3;,�c,0�4���7���;��%?�e�B��7F��I�M��gP���S��V��/Z�^_]�`�`�
�c���f�O�i�V�l�^�o���r�j�u���x�ɗ{�?z~� ����������턼U�����R"��Ǉ���싼nQ������>���|��zߒ��A����������e���ř�r%��Ǆ���㝼�B��$��������^��A�������}��wި�U?������
���c��&ů��&�������購	I��������)h��jǺ��&������  �  �N=�N=}nM=��L=�L=�ZK=ڨJ=^�I=�CI=b�H=��G=+)G=0uF=��E=yE=�WD=ϢC=��B=�7B=��A=��@=�@=�[?=��>=o�==�.==�s<=P�;=�:=�;:=�|9=Ѽ8=��7=	:7=Cw6=n�5=u�4=F(4=�`3=��2=��1=��0=�00=�_/=��.=Ŵ-=��,=��+=�+=9*=�Q)=f(=Jv'=�&=s�%=�$=h�#=��"=-t!=�` =eG=['=� =��=��=�`=G=��=�{==��=RN=�=A^=��=-P=u�	=�%=��=�=i5=Ƀ=��<��<���<��<Pv�<���<�,�<|�<���<Q�<�>�<:s�<h��<���<���<�<�3�<=O�<�g�<�}�<C��<���<���<ھ�<ʤ<�Ӡ<�ۜ<��<&�<#�<g�<�<T�<���<M�y<q�q<�i<Ob<�Z<� R<�0J<�CB<SY:<`q2<a�*<ҩ"<n�< �<<�?<���;!D�;���;|3�;ؽ�;JW�;� �;���;`w;��X;O�:;*�;Pr�:�|�:z�:7�:sF*9Y4��@�8��U����˺�7�`=�?�6�h.Q��k�NB���Ď��������첻t�����ɻ��Ի��߻g�p�������?k�mC	�&�����#�4������$�5(��<,�.0��	4���7��;��&?���B��8F���I��M�	hP��S��V��/Z��^]���`��c���f��i���l���o�*�r���u�^�x�[�{��x~�N���'������센�T��׻��8"��ч���싼�Q���������7}������B��]������ef���ƙ�*&��t���L䝼C������o ��<_��i�������}��Oި��>��*���|�� c���į��%��
����糼8H��L�����ng���ƺ�&��z����  �  j�N=.N=�nM=ǽL=uL=�ZK=��J=�I=2CI=�H=c�G=�(G=�tF=G�E=�E=WD=1�C=��B=M7B=>�A=��@=p@=�[?=�>=e�==/==�s<=��;=j�:=O<:=R}9=`�8=��7=�:7=�w6=�5=#�4=�(4=La3=�2=(�1=D 1=410=�_/=��.=ƴ-=��,=��+=D+=69*=`Q)=�e(=�u'=��&=ʈ%=M�$=̈#=��"=�s!=U` =�F='=Q =��=r�=�`=V=�=�{=r=�=�N=��=�^=��=�P==�	=�&=s�=��=6=q�=��<� �<l��<R�<�v�<��<�,�<�{�<6��<��<�=�<=r�<D��<���<���<��<\2�<�M�<�f�<�|�<H��<���<��<N��<�ɤ<oӠ<�ۜ<9�<y�<��<!�<��<r�<���<�y<?�q<� j<%
b<�Z<A#R<H3J<�EB<[:<�r2<b�*<ɪ"<��<�<�<�><���;*A�;��;�.�;���;�Q�;���;�;Zw;6�X;"�:;��;�a�:?n�:��:��:*9�G����8�)S��8�˺�3��8�@�6��&Q�,k�b=��򿎻�������粻A|����ɻ��Ի �߻�d�v�������Vk��C	����#��.%�̏����C$�y7(�^?,��00�K4���7�d�;�)?���B�G:F�?�I��M��hP�<�S��V�/Z�+^]�e�`���c��f���i���l�W�o�o�r�#�u���x���{�Iv~�0�����D����넼.T�������!��ᇊ�,틼�Q��z���t��~��ᒼ�C����������g���Ǚ�y'������t坼�C��w���� ���_���������}���ݨ��>������� ��b��jï��$������z泼�F���������:f���ź�%�������  �  ��N=|N=�nM=ֽL=nL=�ZK=M�J=��I=�BI=V�H=��G=�'G=�sF=u�E=E=JVD=l�C=-�B=�6B=��A=%�@=@=B[?=Ȣ>=a�==%/==�s<=�;=��:=�<:=�}9=�8=F�7=�;7=�x6=��5=��4=�)4=b3=И2=��1=� 1=�10=�_/=֋.=ʴ-=��,=��+=�+=�8*=�P)= e(=u'=π&=�%=��$=�#=0�"=�r!=�_ =VF=&=��=:�=E�=�`=m=L�=|=�=��=�O=��=�_=��=�Q=@�	=�'=l�=��=�6=A�=���<�!�<p��<	�<;w�<H��<�,�<s{�<���<��<�<�<q�<���<#��<���<�<�0�<EL�<�d�<{�<���<~��<��<���<Xɤ<JӠ<�ۜ<�<��<��<*��<8�<���<a��<g�y<��q<�j<�b<
Z<i&R<Y6J<�HB<s]:<u2<؎*<��"<L�<�<+<�=<���;�<�;��;�(�;r��;�J�;��;���;g�v;�X;��:;�;4J�:�Y�:A؈:��:��)9�Z����8�}P���˺�-��1�i�6�Q���j��7��ƹ��}��g�� ⲻ�v����ɻc�ԻM�߻�a껮�������nk� D	�� ����'�!����/$��:(��B,��30��4���7�r�;�,?�'�B��<F�!�I�>M��iP�~�S� �V��.Z�(]]�ɂ`���c���f�0�i���l�H�o�$�r���u�R�x�Y�{�Gs~�˨�����&����ꄼqS������!��懊�\틼�R��8���q��4��kⒼ$E��������Oi���ə�	)������杼7E���������b`�� ������}���ݨ�>�����������`��¯�9#������䳼'E��G������d��Gĺ��#�������  �  P�N=�N=oM=�L=XL=`ZK= �J=7�I=BI=��H=��G=�&G=�rF=��E= 
E=[UD=t�C=N�B=�5B=�A=��@=�@=�Z?=��>=V�==@/==@t<=F�;=]�:=�=:=�~9=�8=8�7=|<7=�y6=�5=��4=�*4=�b3=��2=x�1=U1=20=X`/= �.=ִ-=��,=O�+=�+=B8*=0P)=Hd(=9t'=�&=�%=��$=�#=M"=�q!=�^ =�E=�%=r�=��=�=�`=�=��=�|=y =f�=eP=t�=�`=��=S=m�	=�(=��=��=8='�==��<#�<���<��<�w�<���<�,�<{�<��<��<�;�<�o�<<��<?��<��<�<�.�<MJ�<c�<qy�<j��<%��<���<˼�<�Ȥ<�Ҡ<�ۜ<��<��<o�<[�<��<��<T��<V�y<� r<�j<�b<!Z<�*R<�9J<�KB<@`:<w2<��*<ެ"<��<��<P<�<<���;�7�;��;6"�;���;�B�;�;{��;|�v;d�X;V�:;_�;+/�:B�:ň:x:�r)9�s��l�8�HL���˺w(��(���6��Q�0�j��0��|���2���9	��.۲�p��+�ɻ8�ԻF�߻_�$�������ik��D	���#��B)�Д�$��}$�`>(�gF,��70��4���7�N�;�]/?�*�B�:?F�G�I��M��jP�)�S�
�V��-Z��[]�D�`���c��f�:�i��l���o�H�r���u�P�x���{��o~����S������鄼�R��v����!�������틼"S�������������㒼�F��
���{
��Xk��q˙��*������k蝼�F��̤����� a������T���}��0ݨ�F=��Ɲ�����n_��o���U!��:����⳼/C��O���7���b���º�o"��o����  �  ��N=@ N=IoM= �L=IL=#ZK=��J=��I=sAI=׍H=�G=&G=�qF=v�E=�E=TTD=s�C=f�B=�4B=8A=��@=@=�Z?=[�>=R�==[/==t<=��;=��:=5>:=v9=ӿ8=*�7=�=7=�z6=��5=�4=�+4=�c3=b�2=3�1=�1=20=�`/=(�.=�-=��,=�+='+=�7*=�O)=qc(=\s'=�~&=�%=��$= �#=P~"=q!=^ =�D=M%=��=��=�=�`=�=��=�|=!=)�=EQ=l�=�a=��=WT=��	=*=͊=�=9=�=���<�$�<���<��<Dx�<���<�,�<�z�<-��<� �<R:�<�m�<���<H��<��<��<�,�<5H�<a�<�w�<���<Ν�<���<仨<!Ȥ<�Ҡ<�ۜ<�<b�<c�<��<$��<>��<B��<��y<ur<$j<�b<�!Z<�.R<�=J<:OB<Ec:<ty2<|�*<�"<c�<��<x<;<\��;�2�;X��;��;���;�9�;��;���;��v;	�X;e�:;��;�:�)�:��:0X:�)9���_�8�8I�� �˺"���O�6��Q���j�)��������7���Ӳ�>i��)�ɻ��Ի��߻�[����� ���Yk��E	�1����+�������"$�SB(��J,�9<0��4���7�F�;��2?���B��AF���I��M��kP�ӶS���V�o-Z��Z]�g`��c��f��i�~�l���o���r���u��x�N�{��k~�:������f~���脼�Q��򹇼J!��퇊�'�S�������������咼�H��
������{m���͙��,��׋��3ꝼFH���������a��������f}���ܨ��<��˜��/����]������x��6����೼A��*���-��a������� ������  �  [�N=� N=�oM=�L=2L=�YK=;�J=*�I=�@I=�H=*�G=%G=�pF=e�E=�E=@SD=s�C=y�B=#4B=y~A=T�@=�@=IZ?=.�>=@�==t/==�t<=�;=v�:=�>:=J�9=��8= 8=�>7=�{6=�5=�4=�,4=�d3=D�2=��1=�1= 30=�`/=Z�.=�-=p�,=��+=�+= 7*=�N)=�b(={r'= ~&=�%=��$= �#=I}"=p!=2] =D=�$=j�=0�=��=�`=�=�=g}=�!=�=R=u�=�b=��=�U=��	=O+=�=/�=+:='�=���<&�<��<��<�x�<���<�,�<?z�<j��<���<�8�<\l�<���<W��<���<��<k*�<F�<#_�<�u�<��<Q��<���<���<�Ǥ<hҠ<�ۜ<}�<�<l�<��<���<��<'��<�z<�	r<�j< b<�%Z<�2R<�AJ<�RB<�e:<�{2<:�*<�"<��<��<�<�9<7��;&-�;��;7�;|��;�0�;�ؙ;���;��v;ňX;*~:;��;n��:��:D��:�6:�(9����8��E��{�˺+����6��P�&�j��!������뚻����{̲��b����ɻ��Իn�߻X�ؽ�������k�-F	�c����.�f������%$�7F(��N,�w@0�14� �7�/�;��6?���B��DF��I�nM�mP�_�S��V��,Z�qY]�|}`�c�\�f���i���l���o��r�W�u��x�1�{��g~�t�����}���焼�P��l���!�����xmT��������s���^璼zJ���������o���ϙ�/�������라�I��g�������b��t������Y}��dܨ��;������ ���n\���������3~���޳��>�����(���,_��!���^������  �  ��N=� N=�oM= �L=L=�YK=٦J=��I=$@I=a�H=U�G=$G=�oF=h�E=�E=GRD=��C=��B=Z3B=�}A=��@=2@=�Y?=��>=/�==�/== u<=j�;=��:=t?:=�9=��8=8=�?7=�|6=�5=��4=�-4=�e3=�2=��1=1=d30=Ba/=��.=�-=S�,={�+=Y+=�6*=2N)=�a(=�q'=}&="�%=��$=�#=\|"=9o!=R\ =jC=$=��=��=s�=�`=�=b�=�}=0"=��=�R=\�=�c=�=�V=�	=y,= �=M�=%;=�=;��<g'�<ܡ�<m�<Yy�<��<v,�<�y�<ƿ�<���<�7�<�j�<��<���<���<�	�<f(�<D�<,]�<�s�<���<隰<���<��<�Ƥ< Ҡ<�ۜ<��<��<Q�<��<��<���<���<�z<�r<�j<b<*Z<�6R<EJ<�UB<�h:< ~2<��*<C�"<F�<]�<�<8<���;�'�;��;�;U��;�(�;�ϙ;퉊;�v;�wX;�l:;ϓ;���:2��:���:y:�g(9������8��A��~�˺�����6���P���j����㛎�#䚻��EŲ�S\���ɻ��Ի`�߻UU����������k��F	������&0�:�����v)$�J(��R,��D0�? 4��7���;�K:?���B��GF��I��M�jnP��S��V�,Z�]X]�|`���c���f���i���l�ܽo�4�r�?�u��x�r�{�d~�١������{���愼MP��⸇�� ��&����)U��κ��$ ��ل���蒼[L��㮕�����q���љ��0�������흼<K���������bc���������<}���ۨ�F;��Ӛ������
[��j������E|���ܳ��<��2���:���`]����������~���  �  9�N=;!N=�oM=&�L=L=�YK=��J=?�I=�?I=��H=��G=e#G=oF=��E=	E=oQD=��C=��B=�2B='}A=8�@=�@=�Y?=ԡ>='�==�/==2u<=Ĺ;=f�:=@:=��9=4�8=�8=I@7=�}6=�5=��4=[.4=Tf3=��2=)�1=�1=�30=�a/=��.=�-=:�,=A�+=�+=*6*=�M)=Na(=�p'=W|&=V�%=��$=3�#=�{"=�n!=�[ =�B=~#=��=��=E�=�`=�=��=)~=�"=&�=�S=!�=�d=��=�W=�	=o-=�=/�=�;=ω=���<�(�<Ӣ�<�<�y�<<��<X,�<Vy�<��<���<�6�<�i�<���<���<M��<�<�&�<qB�<�[�<ur�<&��<���<���<V��<{Ƥ<�Ѡ<�ۜ<�<(�<�<��<O��<
��<�<
z<Ar<�j<�"b<d-Z<�9R<HJ<�XB<k:<�2<'�*<�"<�<6�<1<�6<���;v#�;���;%�;��;�!�;]ș;,��;�v;6iX;�_:;;z��:���:v�:��:�(9�ԏ���8�-?����˺��_���6��P�3�j�	��ᕎ��ݚ��즻�����V���ɻf�Իή߻�R�����-����k�MG	���'��22�������P,$�!M(�V,��G0��#4�V�7��;� =?���B��IF��I��M�moP�`�S��V��+Z�NW]��z`���c�k�f���i���l�Һo��r���u���x�F}{� a~�p���\���z���儼�O��t���� ��/����U������*!�����F꒼�M��s���N��Ds��Uә��2������L��ʩ�����d��`�����3}���ۨ��:����������Y�����o���z��۳�E;�����������[��6�������}���  �  }�N=s!N=pM=5�L=�L=QYK=T�J=��I=<?I=>�H=�G=�"G=XnF=�E=`E=�PD=�C=<�B=2B=�|A=��@=q@=tY?=��>=�==�/==Ou<= �;=��:=b@:=�9=��8=`8=�@7=P~6=��5=x�4=�.4=�f3=5�2=��1=�1=40=�a/=��.=�-=�,=�+=�+=�5*=@M)=�`(=\p'=�{&=��%=�$=��#=�z"=�m!=![ =HB=!#=7�=S�=.�=n`==��=e~=#=��=T=��=�e=��=bX=��	=/.=َ=��=�<=f�=���<Q)�<}��<��<�y�<]��<,�<#y�<���<E��<�5�<�h�<l��<���<���<��<R%�<A�<]Z�<Jq�<��<<©�<ո�<Ƥ<�Ѡ<�ۜ<B�<��<��<���<*��<,��<��<�z<r<)j<j%b<0Z<H<R<JJ<hZB<�l:<�2</�*<��"<��<��<t<�5<���;M �;]��;f�;Ά�;��;�;S|�;�v;$]X;�T:;~|;���:���:�h�:��:�'9|䏹�8�>���|˺j�m�#�6���P�{�j�#�����Oٚ��离���rR��'�ɻt�Իa�߻�P�ʸ�������k��G	��M���3�6������.$��O(��X,��J0�a&4��7���;�f??���B��KF���I��M�pP��S�	�V�|+Z��V]��y`�o�c�ܧf��i�b�l�r�o�7�r�t�u�#�x��z{��^~�A���d���y�� 儼O��5���� ��5���zV��E����!������`뒼�N��Ʊ������t���ԙ��3��S���-𝼎M����������d������B��}���ۨ�B:����������X������=��|y���ٳ�:��;���i����Z���������|���  �  ��N=�!N=pM=<�L=�L=9YK=%�J=��I=�>I=�H=��G=l"G=�mF=��E=�E=cPD=��C=��B=�1B=b|A=��@=:@=FY?=��>=�==�/==eu<=%�;=��:=�@:=`�9=�8=�8=NA7=�~6=�5=��4=P/4=;g3=~�2=��1=11=840=�a/=ʌ.=��-=�,=��+=�+=�5*=�L)=y`(=p'=^{&=P�%=��$=+�#=�z"=�m!=�Z =�A=�"=�='�=�=g`==��=�~=:#=�=qT=�=�e=�=�X=@�	=�.=C�=K�===��=J��<�)�<��<��<"z�<h��<
,�<�x�<,��<���<'5�<�g�<���<��<5��<��<�$�<N@�<�Y�<�p�<j��<M��<C��<l��<�Ť<�Ѡ<�ۜ<e�<��<�<X��<���<���<j�<.z<�r<�j<'b<�1Z<�=R<�KJ<�[B<�m:<.�2<*<�"<��<��<<45<��;��;���;���;���;��;��;�x�;�v;�VX;.N:;�v;��:H��:%`�:��:��'9z폹Y�8��<��4y˺	�S���6�w�P�}�j�~��"���<֚��䦻e���$P�� �ɻ1�Ի^�߻dO� ���H����k�>H	��!���4������0$�+Q(�WZ,�LL0�	(4���7��;��@?��B��LF���I��M��pP�P�S��V�D+Z�NV]��x`�d�c���f�Ųi�/�l��o�دr�բu���x�.y{�]]~��������_y���䄼�N�����s ��>����[V������k"�������뒼�O�����g��hu��uՙ��4�������.N��&������d������T��}��[ۨ�:���������jX��f�������x��ٳ�19��{�������Z������K��Y|���  �  ��N=�N=hM=M�L=-L=�NK=��J=��I=�1I=+}H=�G=�G=W]F=��E=��D=<D=�C={�B=�B=�aA=�@=��?=�8?=f>=��==�	==sM<=5�;=��:=�:=cR9=��8=d�7=�
7=�E6=X5=��4=f�3={#3=�V2=,�1=m�0=f�/=�/=�6.=�[-=�},=x�+=�*=��)=�(=r�'=� '=�&=�%=�$=5#=p�!=Q� =��=�=�=�o=�@=�
=a�=��=�<=��=y�=f*=��=qM=��=�R=m�
==;	=?�=�=�e=ϼ=�=���<�>�<���<t8�<ئ�<v�<�i�<���<�<lT�<���<���<.�<�8�<2f�<׏�<��<Nٿ<���<��<=3�<�L�<�c�<:y�<֌�<���<�<ν�<U˔<�א<!�<��<+��<�<�z<�+r< @j<RUb<*lZ<=�R<A�J<+�B</�:<��2<�+<�A#<�j<ߖ<��<��<g�;���;�j�;$��;A��;�U�;e�;.�;˼{;��];��?;ZV";��;�q�:�{�:��7:��9�;,�����℺ ������ ��l.�� H�
�a��{����+��!,��h�ہ����Ļ'�ϻ��ڻ/u廃����~�U��Ӭ�TW�J��b]�����!�*&��>*�=.��%2� �5�ߺ9�.i=�A� �D��H���K���N��:R���U���X�� \�/0_�;Wb�ive��h���k���n�4�q�˩t��w���z���}�D6��)���a������K���he���ш��<������t���z���⏼�J���������$}���ᖼE��ͧ���	���j��h˝�w+��O����꡼oJ������	���i��1ʨ��*��拫�2��N��K���"���s��ֳ��7��������_^�������#��Æ���  �  ��N=tN=hM=M�L=,L=�NK=њJ=��I=2I=6}H='�G=�G=t]F=ۧE=�D='<D=��C=��B=�B=�aA=�@=��?=9?=g>=��==�	==fM<=*�;=��:=�:=LR9=ܐ8=A�7=�
7=�E6=;5=��4=D�3=d#3=�V2=�1=k�0=[�/=�/=�6.=�[-=�},=�+=�*=��)=�(=}�'=� '=	&=�%=$=T#=��!=n� =��=��= �=�o=�@=�
=Z�=��=�<=��=j�=_*=��=WM=��=�R=I�
=;	=�=�=�e=��=�=���<�>�<i��<K8�<Ʀ�<i�<�i�<��<,�<T�<���<
��<b�<9�<of�<��<[��<�ٿ<���<��<Y3�<�L�<d�<ey�<猤<���<���<���<@˔<�א<#�<��< ��<��<Qz<!+r<�?j<�Tb<�kZ<��R<؝J<йB< �:<��2<�+<�A#<�j<ϖ<��<��<fg�;C��;�j�;���;9��;�V�;x�;,�;��{;��];�?;�W";�;ft�:"~�:��7:�904,�D���ㄺ����������~.�%"H���a��{�;����,���,��_���������Ļz�ϻ��ڻuu����K��e�]�����W���]�Ź���!��)&�O>*��<.�]%2���5�g�9��h=��A���D��H���K�|�N��:R���U���X�� \�X0_�DWb��ve�R�h��k��n���q�A�t�T�w�4�z�N�}�q6��S���k�����_����e���ш��<������J��qz���⏼�J����������|��Tᖼ�D������t	���j��=˝�`+��+����꡼KJ�������	���i��Gʨ��*������3��N��w���Y��:t��0ֳ�"8��6���U����^�������#��Æ���  �  `�N=`N=�gM=M�L=6L=�NK=�J=��I=A2I=s}H=j�G=,G=�]F='�E=`�D=s<D=E�C=��B=B=�aA=J�@=�?=$9?=r>=��==�	==TM<=�;=��:=w:=R9=��8=�7=A
7=@E6=�~5=;�4=��3=&#3=~V2=�1=9�0=7�/=�/=�6.=�[-=�},=��+=�*=�)=U�(=��'=$'=S	&=%=I$=�#=��!=�� =��=5�=Y�=�o=�@=�
=^�=��=�<=��==�= *=[�=
M=J�=0R=��
=�:	=Ť=>=[e=f�=�=��<:>�<��<	8�<���<\�<�i�<;��<^�<�T�<��<���<��<�9�<g�<���<���<ڿ<���<b�<�3�<1M�<Xd�<�y�<��<Ӟ�<��<���<˔<Wא<��<N�<���<U�<2z<�)r<?>j<�Sb<njZ<��R<J<��B<5�:<��2<@+<@A#<uj<�<�<j�<{h�;��;�l�;��;���;�X�;�;���;b�{;��];7�?;p\";��;�|�:��:N8:���9\,����䄺1�����񺙱��.�0%H�.�a�+{�8����.���.��L���<���W�Ļ,�ϻ2�ڻnv�x��u��C�!��F���V�\��\�Ǹ���!�z(&�*=*�e;.�4$2���5�K�9��g=��A�ÑD��H��K��N��:R���U���X�4\��0_�Xb�wwe�Q�h��k��n���q�z�t�x�w�>�z�L�}��6��ѩ�����e��������e���ш��<��p�����-z��|⏼J�������b|������HD���������j���ʝ��*������v꡼J��Щ���	���i��aʨ�+��I�����DO����������t���ֳ��8����������_��x���6$��*����  �  )�N=6N=�gM=A�L=CL=�NK=�J=��I=�2I=�}H=��G=�G=9^F=��E=��D=�<D=C=I�B=�B=IbA=��@=D�?=G9?=�>=�==�	==9M<=�;=��:=):=�Q9=3�8=��7=�	7=�D6=p~5=��4=��3=�"3= V2=��1=�0=�/=�/=�6.=�[-=�},=��+=B�*=G�)=��(=�'=�'=�	&=�%=�$=#=M�!=$� =M�=��=��=*p=�@=�
=p�=��=c<=��=��=�)=��=�L=��=�Q=`�
=(:	=.�=�=�d=޻==D��<�=�<���<�7�<]��<;�<�i�<^��<��<JU�<���<K��<��<z:�<�g�<���<���<$ۿ<|��<=�<�4�<�M�<�d�<z�<p��<��<���<���<�ʔ<�֐<.�<��<���<l �<Hz<�'r<<<j<�Qb<lhZ<��R<��J<X�B<��:<��2<q+<�@#<#j< �<��<�<�j�;Q��;�o�;e�;[��;<]�;h"�;_��;2�{;��];@;Pd";h�;���:���:s8:I�9,�[��儺o���]��f���.�+H�9�a��{�����^2��m2������������ĻC�ϻ-�ڻ�w�[�����W��������U�B���Z�����!��&&�#;*�Z9.�("2�}�5�`�9�f=�;A���D��H�K���N�:R���U���X��\��1_� Yb��xe���h�ˡk�߫n���q�i�t�r�w�+�z��}��7��x���s��䊄������e���ш��<��&�������y���ᏼwI��9���F��i{���ߖ�GC���������0i���ɝ�#*��&����顼�I�������	���i���ʨ�q+������-�O����������u���׳��9��Û�������_��Fº��$��Ç���  �  ��N=�N=�gM=<�L=KL=OK=Q�J=V�I=�2I=J~H=X�G=1G=�^F=A�E=��D=�=D=`�C=��B=B=�bA=�@=��?={9?=�>=�==�	==M<=��;=8�:=�:=HQ9=��8=�7=)	7= D6=�}5=�4=��3=)"3=�U2=&�1=��0=��/=i/=�6.=�[-=�},=ݜ+=��*=��)=�(=��'='=]
&=-%=_$=�#=��!=�� =��=�=��=}p=5A=�
=x�=��=?<=:�=��=Z)=r�=L=�=�P=��
=p9	=q�=�=%d=6�=�=1��<�<�<о�<7�<��<�<�i�<���<@�<�U�<r��<@��<�	�<�;�<.i�<���<9��<hܿ<���<]�<�5�<�N�<�e�<�z�<ȍ�<.��< ��<e��<aʔ<g֐<h�<��<���<H��<�z<=%r<�9j<�Nb<�eZ<M~R<��J<Q�B<�:<m�2<=+<'@#<�i<�<��<��<dm�;���;�s�;�	�;U��;�b�;�'�; �;�{;�];�@;En";X;���:���:))8: 0�9��+�2���愺˺����񺡺��$.�t2H��a��"{�W����6���6������}�����Ļ��ϻ��ڻ�y����7��H�<������T����1Y�����!�"$&��8*��6.��2��5��9��c=�:A�ߎD�OH��}K���N��9R���U�9�X��\��2_�~Zb�dze���h��k�#�n�4�q�үt��w���z�H�}��8��d���L������x���:f���ш��<��馋�p��y��3ᏼ�H��2���(��0z���ޖ�B���������h���ȝ�-)��\���5顼?I��B����	���i���ʨ��+��C�����P����������v���س��:���������a��Mú��%�������  �  ��N=�N=�gM=1�L=bL=2OK=��J=��I=c3I=�~H=��G=�G=�_F= �E=F�D=I>D=�C=��B=�B=DcA=`�@=��?=�9?=�>=�==x	==�L<=a�;=��:=J:=�P9=�8=W�7=v7=eC6=}5=h�4=E�3=�!3=U2=��1=)�0=q�/=2/=^6.=�[-=�},=�+=˸*=�)=��(= �'=�'=&=�%=$=k#=��!=]� =q�=��=w�=�p=qA==|�=��=<=��=>�=�(=ֽ=UK=d�=&P=��
=�8	=��==Rc={�=�=���<�;�<��<{6�<���<�<�i�<���<��<�V�<f��<N��<�<=�<�j�<z��<���<�ݿ<��<��<�6�<�O�<}f�<D{�<B��<p��<��< ��<�ɔ<�Ր<���<��<{�<���<�z<>"r<j6j<�Kb<�bZ<x{R<�J<�B<�:<��2<+<C?#<�i<A�<��<��<p�;j��;qx�;%�;&��;�h�;Z.�;��;��{;��];4@;wy";�;e��:[��:B8:Q�9�+����c鄺����$��y��},.��:H���a��,{����a<��<�����������Ļ,�ϻ��ڻ�{�\�����������US�#��W����!�[!&��5*��3.��2��5�/�9�'a=��@���D��H��|K���N�E9R���U���X�a\��3_�\b�`|e��h�V�k��n���q��t��w�q�z��}�
:������>��K�������f��҈��<���������ux��]����G���������x��ݖ��@��?���F���f���ǝ�(��a����衼�H��ۨ��P	��j��˨�b,����לּ�Q��鳯���Bx��hڳ�{<��t���a ��ab��yĺ��&��k����  �   �N=yN=ugM=#�L=pL=ZOK=�J=�I=�3I=eH=��G=�G=K`F=ΪE=�D=?D=ˈC=8�B=?B=�cA=ݫ@=I�?=:?=�>=#�==a	==�L<=�;=n�:=�:=P9=i�8=��7=�7=�B6=I|5=��4=��3=� 3=hT2=!�1=��0=�/=�/=66.=�[-=~,=K�+=#�*=n�)=�(=��'=]'=�&=�%=�$=.	#=X�!=� =�=�=��=5q=�A===��=q�=�;=��=ɋ=G(=8�=�J=��=@O=��
=�7	=��=0=lb=��==ĭ�<�:�<$��<�5�<B��<��<�i�<Z��<P�<wW�<k��<~��<c�<k>�<Cl�<
��<_��<o߿<���<�<8�<�P�<eg�<|�<���<���<���<ۼ�<�ɔ<Ր<�ߌ<��<$�<y��<�z<r<3j<�Hb<�_Z<OxR<:�J<b�B<��:<��2<�+<m>#<9i<Y�<+�<6�<As�;���;A}�;��;)��;Mo�;q5�;��;�{;*�];&@;��";�; ��:���:0]8:Tq�9�+����.넺�Ż�V��X���4.��CH�I�a��7{�3
��B���A�����.�����Ļ��ϻ�ڻi~建�������P������Q�O���T�g��C�!��&��2*��0.�d2���5�\�9�e^=���@���D��	H�Y{K���N��8R���U�:�X�#\�:5_��]b�[~e��h��k��n���q���t���w�v�z�	�}�c;��í��.��&��������f��Q҈��<��s���]���w��mߏ�fF��ά��j��aw��tۖ��>���������Ee��EƝ��&��P����硼H������1	��j��a˨��,���������R��8�������y���۳�
>����������c���ź��'��V����  �  ��N=(N=NgM=�L=�L=�OK=-�J=w�I=`4I=�H=F�G=KG=aF=��E=��D=�?D=��C=��B=�B=`dA=Q�@=��?=E:?="�>=+�==O	==�L<=��;=�:=J:=�O9=��8=��7=�7=�A6=�{5=ڳ4=��3=' 3=�S2=��1=>�0=��/=�/=6.=�[-=,~,=w�+=u�*=��)=��(=R�'='=r&=c%=�$=�	#=�!=�� =��=��=d�=�q=B=Z=��=X�=�;=L�=R�=�'=��=�I=��=iN=��
=�6	=��=C=�a=ڸ=O
=j��<m9�<2��<B5�<ޤ�<��<j�<���<��<AX�<_��<���<��<�?�<�m�<���<��<�<�<{�<W9�<�Q�<Oh�<�|�<��<ܟ�<���<���<�Ȕ<?Ԑ<�ތ<x�<��<
��<�z<�r<�/j<)Eb<D\Z<HuR<f�J<ۭB<��:<,�2<i+<�=#<�h<|�<��<8 <�v�;���;��;W�;v��;�u�;*<�;��;�|;=^;R3@;�";W";���:�ʕ:�s8:#��9Kg+����i턺"ͻ�p	�_��l<.�MH�*�a��B{����G���G�����M���A�Ļлv�ڻ�廍�ﻐ�������/��pP�����R�ڭ�}�!�p&�w/*�x-.�E2���5�G�9��[=��@���D�*H��yK�9�N�M8R���U���X�\��6_��_b���e���h�۫k�Ѷn�/�q��t�$�w���z�ѐ}��<��󮁼C�����W���]g��|҈��<��$�������v���ޏ�YE���������u���ٖ�d=�����7���c���ĝ��%��c����桼qG��,���	��3j���˨�t-��z�����T��������G{���ݳ��?������l��8e��Ǻ�)��_����  �  i�N=�N="gM= �L=�L=�OK=j�J=��I=�4I=��H=��G=�G=�aF=H�E=��D=�@D=D�C=��B=yB=�dA=��@=��?=}:?=J�>=.�==8	==RL<=u�;=��:=�:= O9=�8=8�7=97=A6=�z5=�4=�3=y3=9S2=
�1=մ0=f�/=u/=�5.=�[-=@~,=��+=��*=:�)=��(=��'=�'=&=%=V$=�
#=��!=k� =K�=;�=֚=�q=<B=}=��=8�=o;=��=�=7'=�=)I=��=�M=�
=�5	=՟=h=�`=�=�	=#��<v8�<f��<�4�<~��<w�<1j�<���<h�<�X�<K��<���<��<OA�<'o�<-��<h��<q�<~�<��<�:�<�R�<i�<=}�<���<��<߮�<_��<qȔ<�Ӑ<�݌<d�<���<���<�z<�r<�,j<�Ab<HYZ<[rR<��J<�B<��:<��2<+<�<#<gh<��<o�<-<my�;:��;���;_�;%ƺ;|�;�B�;��;�|;^;"?@;�";w,;���:�ؕ:�8:(��9�G+��������ӻ�������C.�&VH��b�=M{����^M�� M����Y���_�Ļ�лt�ڻ/��^��/���G��M��BO�����P�}���!��&��,*�q*.�12��5�r�9�/Y=���@���D��H��xK�f�N��7R�ĆU��X�\��7_�Eab���e�!�h���k���n�#�q��t�"�w�z�z���}�>�����J �����������g���҈��<��ݥ�����Zv���ݏ�VD��\������nt���ؖ��;������� ��tb���Ý��$��|���&桼�F��˧�����Yj���˨� .�������U������C���|��߳�A���������f��MȺ�"*��K����  �  �N=�N=gM=��L=�L=�OK=��J=�I=55I=��H=a�G=�G=]bF=�E=2�D=-AD=ڊC=�B=�B=WeA= �@=F�?=�:?=_�>=2�==*	==-L<=7�;=M�:=d:=�N9=��8=��7=�7=w@6=z5=��4=~�3=�3=�R2=��1=t�0=�/=E/=�5.=�[-=M~,=֝+=��*=��)=h�(=V�'=!'=�&=�%=�$=>#=S "=�� =��=��=<�=9r=rB=�=��=&�=C;=��=��=�&=c�=�H=N�=�L=h�
=5	=�=�=`=l�=	=��<�7�<���<4�<0��<U�<3j�<<��<��<�Y�<��<���<��<sB�<dp�<_��<���<��<��<� �<�;�<�S�<�i�<�}�<ߏ�<*��<ᮜ<)��<Ȕ<�Ґ<�܌<s�<��<u��<z<�r<�)j<a?b<�VZ<�oR<l�J<i�B<��:<�2<+<)<#<3h<��<��<3<�{�;���;���;�#�;�ʺ;b��;H�;� �;�|;�^;ZI@;�";5;3��:	�:|�8:�͌9B-+������6ػ���4��WJ.��]H�Zb�!V{���R���Q�����~���+�Ļ:
л5�ڻn�廣���������z��N����O������!�O&�**��'.��2���5�(�9�W=���@�ЄD�2H��wK���N��7R�ÆU�g�X��\� 9_��bb�a�e�"�h���k���n���q���t���w��z��}�?�� ���!��y���j���"h���҈��<���������u���܏�rC��[������Es��Oז��:��h�������Va�����#�������塼mF���������aj��1̨�i.��ǐ��`�V������e���}��:೼]B��H������g��Zɺ�+������  �  ��N=�N=�fM=�L=�L=�OK=לJ=V�I=�5I=F�H=��G=�G=�bF=k�E=��D=�AD=N�C=��B=]B=�eA=j�@=z�?=�:?=v�>=>�==	==
L<=
�;=	�:=:= N9=+�8=.�7=7=�?6=�y5=�4=�3=�3=KR2=I�1=1�0=��/=%/=�5.=�[-=\~,=�+=(�*=��)=��(=��'=�'=&=$%=j$=�#=� "=_� =6�=��=~�=sr=�B=�=��=�=;=��=D�=m&=�=H=��=VL=��
=}4	=��==�_=�=�=e��<�6�<.��<�3�<ޣ�<N�<Aj�<n��<(�<"Z�<���<r��<��<TC�<cq�<T��<���<��<��<�!�<*<�<cT�<Kj�<4~�<��<O��<خ�<㻘<�ǔ<wҐ<r܌<��<��<���<z<�r<�'j<H=b<~TZ<�mR<��J<ۧB<��:<��2<[+<|;#<�g<Ɨ<5�<�<�}�; �;8��;Z'�;�κ;x��;�L�;%�;�"|;$^;zQ@;��";�:;���:��:��8:�9�+����&���ܻ��!�����O.�dcH��b�}]{�����U��DU��3������I�Ļ�л!�ڻ��x�������������[M�s���M�7���!��&�"(*��%.��2���5�d�9�=U=�c�@���D�$H� wK��N�b7R���U���X�D\��9_��cb���e�˟h�W�k��n���q���t���w��z�ŗ}��?��ͱ���!���������dh���҈��<���������ku��`܏��B���������`r��N֖��9��h�������w`������#�����塼F��Q������pj��}̨��.��G����󬼴V������?���~��4᳼cC��D���	���h��+ʺ��+�������  �  ��N=eN=�fM=�L=�L=�OK=�J=��I=�5I=��H=�G=0G=cF=��E= �D=�AD=��C=��B=�B=�eA=��@=��?=�:?=��>=;�==	==�K<=�;=��:=�:=�M9=�8=��7=�7=�?6=Sy5=��4=��3=<3=	R2=
�1=��0=��/=	/=�5.=�[-=`~,=�+=D�*=��)=��(=��'=�'=V&=e%=�$= #="=�� =p�=8�=��=�r=�B=�=��=�=�:=a�=�=0&=��=�G=��=L=~�
=&4	=.�=�=1_=��=I=ը�<n6�<׹�<t3�<���<5�<Hj�<���<g�<~Z�<��<���<O�<�C�<�q�<���<E��<6�<�<3"�<�<�<�T�<�j�<g~�<E��<W��<ʮ�<ʻ�<�ǔ<3Ґ<܌<A�<#�<���<��y<�r<~&j<<b<SSZ<�lR<��J<ҦB<��:<\�2<�+<2;#<�g<Ɨ<w�<7<�;��;R��;s)�;�к;ˇ�;�N�;�'�;�'|;)^;�U@;H�";�?;O�:��:P�8:(�9^	+���������޻�a%�)��/S.�(gH�b��a{����X��vW��?������9�Ļ]л��ڻ��9�������������L�����L�2���!��&�'*��$.��2�o�5�[�9�BT=�a�@���D�WH�|vK���N�H7R���U��X��\�h:_��db���e�ˠh�m�k���n���q���t�ùw��z���}�o@��F���$"��V�������h��ӈ��<��{������!u���ۏ�cB�� ���Q���q���Ֆ�9��ٛ������_��d����"�������䡼�E��.�������j���̨��.������U���0W��������j���᳼�C��ܥ�����"i���ʺ�D,������  �  ��N=ON=�fM=�L=�L=PK=��J=��I=�5I=��H=�G=OG=:cF=ǭE=�D=BD=��C=��B=�B=�eA=��@=��?=;?=��>=8�==	==�K<=ۍ;=��:=�:=�M9=ҋ8=��7=�7=�?6=3y5=��4=��3=!3=�Q2=��1=�0=��/=�/=�5.=�[-=d~,=�+=M�*=��)=��(=��'=�'=z&=�%=�$=#=+"=�� =��=J�=��=�r=�B=�=��=�= ;=Q�=	�=!&=��=�G=d�=�K=]�
=4	=	�=�=_=��=;=���<R6�<���<b3�<���<*�<Vj�<���<z�<Z�<4��<��<��<"D�< r�<5��<u��<{�<S�<e"�<�<�<�T�<�j�<}~�<`��<V��<Ȯ�<ǻ�<_ǔ<Ґ<�ی<$�<�<���<n�y< r<&j<;b<�RZ<SlR<9�J<��B<n�:<$�2<�+<$;#<�g<ė<��<l<^�;��; ��;>*�;�Ѻ;�;�O�;�(�;h)|;g+^;�W@;ݳ";�@;��:{��:x�8:@�9
+���� ����໺�&�A���S.��hH��b�_c{�� �� Y��lX����n�����Ļ�л�ڻj���������}��e���L�����L�����!��&��&*�V$.�2���5�Σ9��S=��@���D�KH�VvK��N�47R���U��X��\��:_��db�Ȇe���h�سk�k�n�%�q�M�t�G�w�y�z�V�}��@��^���I"��l���(����h��ӈ��<��j���{��u���ۏ�FB���������q���Ֆ��8�����������_��2���t"�������䡼�E���������j���̨�/������t���KW��0��������⳼2D��������]i���ʺ�],��/����  �  ��N=eN=�fM=�L=�L=�OK=�J=��I=�5I=��H=�G=0G=cF=��E= �D=�AD=��C=��B=�B=�eA=��@=��?=�:?=��>=;�==	==�K<=�;=��:=�:=�M9=�8=��7=�7=�?6=Sy5=��4=��3=<3=	R2=
�1=��0=��/=	/=�5.=�[-=`~,=�+=D�*=��)=��(=��'=�'=V&=e%=�$= #="=�� =p�=8�=��=�r=�B=�=��=�= ;=b�=�=2&=��=�G=��=L=��
=)4	=1�=�=5_=��=M=ި�<w6�<��<}3�<���<>�<Pj�<���<o�<�Z�<��<���<S�<�C�<�q�<���<D��<5�<�</"�<�<�<�T�<�j�<`~�<>��<P��<î�<û�<�ǔ<-Ґ<�ی<<�<�<���<��y<�r<~&j<<b<WSZ<�lR<��J<ܦB<��:<h�2<�+<@;#<�g<ԗ<��<D<4�;��;f��;�)�;�к;҇�;�N�;�'�;�'|;�(^;�U@;�";_?;��:s�:=�8:��9*+���4���m߻�&�x��{S.�qgH�Kb��a{� ��X���W��W������L�Ļnл��ڻ ��E��%�����������L�����L�3���!��&�'*��$.��2�o�5�\�9�CT=�a�@���D�WH�}vK���N�H7R���U��X��\�h:_��db���e�ˠh�m�k���n���q���t�ùw��z���}�o@��F���$"��V�������h��ӈ��<��{������!u���ۏ�cB�� ���Q���q���Ֆ�9��ٛ������_��d����"�������䡼�E��.�������j���̨��.������U���0W��������j���᳼�C��ܥ�����"i���ʺ�D,������  �  ��N=�N=�fM=�L=�L=�OK=לJ=V�I=�5I=F�H=��G=�G=�bF=k�E=��D=�AD=N�C=��B=]B=�eA=j�@=z�?=�:?=v�>=>�==	==
L<=
�;=	�:=:= N9=+�8=.�7=7=�?6=�y5=�4=�3=�3=KR2=I�1=1�0=��/=%/=�5.=�[-=\~,=�+=(�*=��)=��(=��'=�'=&=$%=j$=�#=� "=_� =7�=��=�=tr=�B=�=��= �=;=��=G�=o&=�=H=��=ZL=��
=�4	=��=#=�_=��=�=v��<�6�<@��<�3�<��<_�<Rj�<~��<6�</Z�<���<{��<��<ZC�<fq�<U��<���<��<��<�!�<!<�<XT�<?j�<'~�<��<A��<ˮ�<ջ�<�ǔ<kҐ<g܌<��<��<���<z<�r<�'j<L=b<�TZ<nR<��J<�B<��:<�2<u+<�;#<h<�<Q�<�<�}�;K �;]��;x'�;�κ;���;�L�;%�;�"|;�#^;;Q@;h�";�:;���:��:�8:�݌95+����]���=ݻ��"�}��eP.��cH�wb��]{����V��vU��a������n�Ļ�л>�ڻ3�廎�������������`M�x���M�:���!��&�#(*��%.��2���5�e�9�=U=�c�@���D�%H� wK��N�b7R���U���X�D\��9_��cb���e�˟h�W�k��n���q���t���w��z�ŗ}��?��ͱ���!���������dh���҈��<���������ku��`܏��B���������`r��N֖��9��h�������w`������#�����塼F��Q������pj��}̨��.��G����󬼴V������?���~��4᳼cC��D���	���h��+ʺ��+�������  �  �N=�N=gM=��L=�L=�OK=��J=�I=55I=��H=a�G=�G=]bF=�E=2�D=-AD=ڊC=�B=�B=WeA= �@=F�?=�:?=_�>=2�==*	==-L<=7�;=M�:=d:=�N9=��8=��7=�7=w@6=z5=��4=~�3=�3=�R2=��1=t�0=�/=E/=�5.=�[-=M~,=֝+=��*=��)=h�(=V�'=!'=�&=�%=�$=>#=T "=�� =��=��==�=:r=tB=�=��=(�=E;=��=��=�&=h�=�H=T�=�L=o�
=5	=#�=�=`=w�=	=5��<�7�<˺�<04�<I��<m�<Jj�<R��<��<�Y�<-��<���<�<zB�<hp�<`��<���<��<��<� �<s;�<�S�<�i�<�}�<̏�<��<ͮ�<��<�ǔ<�Ґ<�܌<e�<z�<l��<z<�r<�)j<g?b<�VZ<�oR<��J<��B<��:<<�2<7+<P<#<[h<×<��<X<|�;���;Ί�;�#�;˺;v��;H�;� �;�|;�^;I@;�";�4;���:��:��8:zǌ9_:+����k��ٻ�����'K.�o^H�b��V{�e��`R���Q���������_�Ļh
л^�ڻ��������������&N����O������!�R&� **��'.��2���5�)�9�W=���@�ЄD�2H��wK���N��7R�ÆU�g�X��\� 9_��bb�a�e�"�h���k���n���q���t���w��z��}�?�� ���!��y���j���"h���҈��<���������u���܏�rC��[������Es��Oז��:��h�������Va�����#�������塼mF���������aj��1̨�i.��ǐ��`�V������e���}��:೼]B��H������g��Zɺ�+������  �  i�N=�N="gM= �L=�L=�OK=j�J=��I=�4I=��H=��G=�G=�aF=H�E=��D=�@D=D�C=��B=yB=�dA=��@=��?=}:?=J�>=.�==8	==RL<=u�;=��:=�:= O9=�8=8�7=97=A6=�z5=�4=�3=y3=9S2=
�1=մ0=f�/=u/=�5.=�[-=@~,=��+=��*=:�)=��(=��'=�'=&=%=W$=�
#=��!=k� =L�=<�=ך=�q==B=~=��=:�=r;=��=�=;'=�=0I=��=�M='�
=�5	=��=t=�`=�=�	=A��<�8�<���<�4�<���<��<Nj�<���<��<Y�<_��<���<��<YA�<-o�</��<f��<k�<u�<��<x:�<�R�<	i�<'}�<t��<���<Ǯ�<H��<ZȔ<�Ӑ<�݌<T�<���<���<�z<zr<�,j<Bb<VYZ<prR<ՍJ<��B<��:<��2<H+<�<#<�h<ʗ<��<Z<�y�;���; ��;��;Lƺ;/|�;�B�;��;Y|;�^;�>@;\�";�+;W��:Bו:[�8:|��9�W+������"ջ������D.�WH��b�N{�����M��wM��P��������Ļ,л��ڻ[�廄��P��%�S��W��KO�����P�����!��&��,*�t*.�32��5�t�9�0Y=���@���D��H��xK�f�N��7R�ĆU��X�\��7_�Eab���e�!�h���k���n�#�q��t�"�w�z�z���}�>�����J �����������g���҈��<��ݥ�����Zv���ݏ�VD��\������nt���ؖ��;������� ��tb���Ý��$��|���&桼�F��˧�����Yj���˨� .�������U������C���|��߳�A���������f��MȺ�"*��K����  �  ��N=(N=NgM=�L=�L=�OK=-�J=w�I=`4I=�H=F�G=KG=aF=��E=��D=�?D=��C=��B=�B=`dA=Q�@=��?=E:?="�>=+�==O	==�L<=��;=�:=J:=�O9=��8=��7=�7=�A6=�{5=ڳ4=��3=' 3=�S2=��1=>�0=��/=�/=6.=�[-=,~,=w�+=u�*=��)=��(=R�'='=r&=c%=�$=�	#=�!=�� =��=��=e�=�q=B=\=��=[�=�;=P�=V�=�'=��=�I=��=sN=�
=�6	= =P=�a=�=_
=���<�9�<T��<d5�< ��<��<6j�<���<�<ZX�<u��<���<��<�?�<�m�<���<��<��<�<m�<F9�<�Q�<9h�<�|�<���<���<ޮ�<���<�Ȕ<'Ԑ<�ތ<f�<��<���<�z<�r<�/j<1Eb<T\Z<`uR<��J<�B<��:<[�2<�+<�=#<i<��<��<k <�v�;���;c��;��;���;v�;4<�;��;�|;�^;�2@;J�";�!;���:�ȕ:�o8:���95y+�4���}ϻ������=.�&NH�-�a��C{����<H���G��M��������ĻKл��ڻ9�廷�ﻵ������:��zP�����R�����!�t&�z/*�{-.�G2���5�I�9��[=��@���D�+H��yK�9�N�N8R���U���X�\��6_��_b���e���h�۫k�Ѷn�/�q��t�$�w���z�ѐ}��<��󮁼C�����W���]g��|҈��<��$�������v���ޏ�YE���������u���ٖ�d=�����7���c���ĝ��%��c����桼qG��,���	��3j���˨�t-��z�����T��������G{���ݳ��?������l��8e��Ǻ�)��_����  �   �N=yN=ugM=#�L=pL=ZOK=�J=�I=�3I=eH=��G=�G=K`F=ΪE=�D=?D=ˈC=8�B=?B=�cA=ݫ@=I�?=:?=�>=#�==a	==�L<=�;=n�:=�:=P9=i�8=��7=�7=�B6=I|5=��4=��3=� 3=hT2=!�1=��0=�/=�/=66.=�[-=~,=K�+=#�*=n�)=�(=��'=]'=�&=�%=�$=.	#=Y�!=� =�=�=��=6q=�A=?=��=t�=�;=��=͋=L(=?�=�J=��=IO=��
=�7	=��=>={b=��==��<�:�<H��<6�<e��<��<j�<y��<m�<�W�<���<���<r�<v>�<Jl�<��<]��<i߿<���<�<8�<�P�<Mg�<�{�<���<���<㮜<���<oɔ<�Ԑ<�ߌ<��<�<m��<�z<r<3j<�Hb<�_Z<hxR<Z�J<��B<*�:<-�2<+<�>#<ri<��<b�<k�<�s�;��;�}�;��;V��;io�;{5�;��;��{;��];�%@;�";�;j��:���:Y8:yh�9n�+�����턺Ȼ������5.��DH�V�a��8{��
���B��B��
	��������Ļ5�ϻV�ڻ�~�������^�����Q�X���T�m��H�!��&��2*��0.�f2���5�^�9�f^=���@���D��	H�Z{K���N��8R���U�:�X�#\�:5_��]b�[~e��h��k��n���q���t���w�v�z�	�}�c;��í��.��&��������f��Q҈��<��s���]���w��mߏ�fF��ά��j��aw��tۖ��>���������Ee��EƝ��&��P����硼H������1	��j��a˨��,���������R��8�������y���۳�
>����������c���ź��'��V����  �  ��N=�N=�gM=1�L=bL=2OK=��J=��I=d3I=�~H=��G=�G=�_F= �E=F�D=I>D=�C=��B=�B=DcA=`�@=��?=�9?=�>=�==x	==�L<=a�;=��:=J:=�P9=�8=W�7=v7=eC6=}5=h�4=E�3=�!3=U2=��1=)�0=q�/=2/=^6.=�[-=�},=�+=˸*=�)=��(= �'=�'=&=�%=$=k#=��!=]� =q�=��=x�=�p=rA==�=��=<=��=B�=�(=ܽ=\K=l�=0P=��
=�8	=��=$=`c=��=�=��<�;�<+��<�6�<ץ�<"�<j�<��<��<�V�<|��<a��<�<=�<�j�<|��<���<�ݿ<��<��<�6�<�O�<ff�<+{�<(��<U��<鮜<��<�ɔ<�Ր<z��<��<k�<���<�z<6"r<i6j<�Kb<�bZ<�{R<=�J<�B<>�:< �2<G+<x?#<�i<x�<��<(�<_p�;���;�x�;`�;Q��;�h�;d.�;��;Y�{;^�];�@;�x";�;���:���:>8:�H�9��+�8���넺����z�����-.��;H���a��-{����<��z<��S��H����Ļk�ϻ	�ڻ�{廆��$��+�������_S�,��W���
�!�_!&��5*��3.��2��5�1�9�(a=��@���D��H��|K���N�E9R���U���X�a\��3_�\b�`|e��h�V�k��n���q��t��w�q�z��}�
:������>��K�������f��҈��<���������ux��]����G���������x��ݖ��@��?���F���f���ǝ�(��a����衼�H��ۨ��P	��j��˨�b,����לּ�Q��鳯���Bx��hڳ�{<��t���a ��ab��yĺ��&��k����  �  ��N=�N=�gM=<�L=KL=OK=Q�J=V�I=�2I=J~H=X�G=1G=�^F=A�E=��D=�=D=`�C=��B=B=�bA=�@=��?={9?=�>=�==�	==M<=��;=8�:=�:=HQ9=��8=�7=)	7= D6=�}5=�4=��3=)"3=�U2=&�1=��0=��/=i/=�6.=�[-=�},=ݜ+=��*=��)=�(=��'='=^
&=-%=`$=�#=��!=�� =��=�=��=~p=6A=�
=z�=��=B<=>�=��=_)=x�=L=&�=Q=��
=z9	=|�=�=2d=D�=�=N��<�<�<��<:7�<2��<.�<�i�<���<Y�<V�<���<P��<�	�<�;�<3i�<���<7��<bܿ<���<P�<�5�<�N�<�e�<�z�<���<��<箜<M��<Kʔ<R֐<U�<��<���<>��<�z<5%r<�9j<�Nb<�eZ<b~R<ИJ<s�B</�:<��2<k+<W@#<j<5�<&�<�<�m�;���;5t�;
�;|��;�b�;�'�;���;��{;��];1@;�m";�;��:��:�%8:U(�9��+�V���脺缻���񺨻��%.�i3H��a��#{�����7��M7�����ċ����Ļ��ϻ��ڻ�y���X��V�H�����T����7Y�����!�&$&��8*��6.��2��5��9��c=�;A���D�OH��}K���N��9R���U�9�X��\��2_�~Zb�dze���h��k�#�n�4�q�үt��w���z�H�}��8��d���L������x���:f���ш��<��馋�p��y��3ᏼ�H��2���(��0z���ޖ�B���������h���ȝ�-)��\���5顼?I��B����	���i���ʨ��+��C�����P����������v���س��:���������a��Mú��%�������  �  )�N=6N=�gM=A�L=CL=�NK=�J=��I=�2I=�}H=��G=�G=9^F=��E=��D=�<D=C=I�B=�B=IbA=��@=D�?=G9?=�>=�==�	==9M<=�;=��:=):=�Q9=3�8=��7=�	7=�D6=p~5=��4=��3=�"3= V2=��1=�0=�/=�/=�6.=�[-=�},=��+=B�*=G�)=��(=�'=�'=�	&=�%=�$=#=M�!=$� =M�=��=��=+p=�@=�
=r�=��=f<=��= �=�)=�=�L=��=�Q=g�
=1:	=7�=�=�d=�=!=\��<�=�<���<�7�<v��<S�<�i�<t��<��<\U�<���<X��<��<�:�<h�<���<���<ۿ<u��<3�<�4�<�M�<�d�<z�<]��<�<宜<s��<�ʔ<�֐<�<��<���<d �<<z<�'r<<<j<�Qb<whZ<ʀR<�J<s�B<��:<��2<�+<�@#<Kj<(�<��<&�<�j�;���;+p�;��;{��;P]�;p"�;Y��;�{;��];�@;�c";��;Ɇ�:E��:�8:�99,�����愺(�����=���.��+H���a��{�"����2���2����������3�Ļq�ϻV�ڻ�w�{�����c��������U�H���Z�!����!��&&�%;*�\9.�)"2�~�5�a�9�f=�;A���D��H�K���N�:R���U���X��\��1_� Yb��xe���h�ˡk�߫n���q�i�t�r�w�+�z��}��7��x���s��䊄������e���ш��<��&�������y���ᏼwI��9���F��i{���ߖ�GC���������0i���ɝ�#*��&����顼�I�������	���i���ʨ�q+������-�O����������u���׳��9��Û�������_��Fº��$��Ç���  �  `�N=`N=�gM=M�L=6L=�NK=�J=��I=A2I=s}H=j�G=,G=�]F='�E=`�D=s<D=E�C=��B=B=�aA=J�@=�?=$9?=r>=��==�	==TM<=�;=��:=w:=R9=��8=�7=A
7=@E6=�~5=;�4=��3=&#3=~V2=�1=9�0=7�/=�/=�6.=�[-=�},=��+=�*=�)=U�(=��'=$'=S	&=%=I$=�#=��!=�� =��=6�=Y�=�o=�@=�
=_�=��=�<=��=@�=#*=^�=M=O�=5R=��
=�:	=ˤ=E=ce=n�=�=��<L>�<&��<8�<���<m�<�i�<J��<l�<�T�<��<���<��<�9�<g�<���<���<ڿ<���<[�<�3�<&M�<Md�<�y�<��<Ş�<���<���<˔<Jא<��<E�<y��<O�<*z<�)r<?>j<�Sb<vjZ<��R<ҜJ<˸B<K�:<��2<[+<\A#<�j<��<�<��<�h�;<��;m�;�;���;�X�;�;���;G�{;��];��?;!\";q�;�{�:��::8:w�9�',�	��G儺i���"��0��R.��%H���a��{�s��� /���.��z���e���|�ĻM�ϻO�ڻ�v廎�ﻈ��L�(��L���V�`��\�ʸ���!�|(&�+=*�f;.�5$2���5�L�9��g=��A�ÑD��H��K��N��:R���U���X�4\��0_�Xb�wwe�Q�h��k��n���q�z�t�x�w�>�z�L�}��6��ѩ�����e��������e���ш��<��p�����-z��|⏼J�������b|������HD���������j���ʝ��*������v꡼J��Щ���	���i��aʨ�+��I�����DO����������t���ֳ��8����������_��x���6$��*����  �  ��N=tN=hM=M�L=,L=�NK=њJ=��I=2I=6}H='�G=�G=t]F=ۧE=�D='<D=��C=��B=�B=�aA=�@=��?=9?=g>=��==�	==fM<=*�;=��:=�:=LR9=ܐ8=A�7=�
7=�E6=;5=��4=D�3=d#3=�V2=�1=k�0=[�/=�/=�6.=�[-=�},=�+=�*=��)=�(=}�'=� '=	&=�%=$=T#=��!=n� =��=��= �=�o=�@=�
=[�=��=�<=��=l�=a*=��=YM=��=�R=L�
=;	=!�=�=�e=��=�=���<�>�<r��<T8�<Ϧ�<r�<�i�< ��<3�<�T�<���<��<f�<9�<qf�<��<[��<�ٿ<���<��<T3�<�L�<�c�<^y�<���<���<ﮜ<���<9˔<�א<�<��<���<��<Mz<+r<�?j<�Tb<�kZ<R<��J<ڹB<+�:<��2<�+<�A#<�j<ݖ<��<�<g�;Y��;	k�;���;E��;�V�;{�;*�;�{;��];��?;jW";��;�s�:�}�:��7:��9�8,����-䄺\���{��D���.�n"H�+�a��{�Y����,���,��w���������Ļ��ϻ��ڻ�u���U��i�a�����W���]�ƹ���!��)&�P>*��<.�^%2���5�h�9��h=��A���D��H���K�|�N��:R���U���X�� \�X0_�DWb��ve�R�h��k��n���q�A�t�T�w�4�z�N�}�q6��S���k�����_����e���ш��<������J��qz���⏼�J����������|��Tᖼ�D������t	���j��=˝�`+��+����꡼KJ�������	���i��Gʨ��*������3��N��w���Y��:t��0ֳ�"8��6���U����^�������#��Æ���  �  ��N=�N=R`M=��L=��K=DDK=��J=��I=%I=noH=i�G=4G=�LF=�E=��D=�'D=0pC=G�B=��A=4GA=Ѝ@=��?=1?=�]>=��==f�<=>&<=g;=��:=��9=W#9=�_8=�7=�6=�6=�D5=�z4=�3=B�2=�2=f@1=�l0=͖/=P�.=2�-=+-='$,=�?+=]X*=Km)=�~(=��'=J�&=��%=B�$=r�#=Ԏ"=$�!=:n =�U=v7=)=��=��=�=A=M�=p�=>Z=��=�=�1=��=1H=��=�B
=t�=�!=�=��=�A=Q� =*��<O]�<5��<�e�<���<I�<J��<��<b�<|��<���<n>�<�|�<M��<d��<��<9J�<�t�<���<���<��<Q�<��<g;�<U�< m�<N��<*��<���<!��<�ό<e��<���<� �<� z<�@r<aj<C�b<�Z<��R<j�J<bC<N@;<�l3<�+<n�#<�<�<<�y<c�<�;s��;�?�;���;��;-��;�b�;�W�;"`�;��b;RhE;Q(;��
;y��:E#�:NR:��9�s������9l�Ȁ���D�|��"�%���?�5GY��cr����浑������d���괻8���M˻�+ֻz���?�gv���v�����jk	�������0���� ��$��8(��B,�p70�s4�4�7�;�;��L?���B��sF���I�lbM���P�S T��nW���Z���]�x"a�DMd�pg���j�h�m�k�p�`�s�u�v��y���|���<G��޼���0�������΃����p`��g͌�S9���������nx��ᓼ�H��ܯ�����/{���ߚ�tC��Ʀ��y	���k��Ρ�70��;���P����V����������~���ᬼ�D��K������To��ӳ��6�����������b��Ǻ��+�������  �  ��N=�N=H`M=��L=��K=QDK=��J=��I=$%I=xoH=y�G=@G=�LF=�E=	�D=�'D=;pC=T�B= B==GA=��@=��?=H?=�]>=��==\�<=;&<=g;=�:=��9=D#9=�_8=��7=��6=�6=�D5=�z4=Ԯ3=C�2=�2=Z@1=�l0=/=O�.='�-=(-=*$,=�?+=hX*=Vm)=�~(=��'=^�&=��%=V�$=��#=�"=9�!=An =�U=�7=4=��=��=�=A=M�=c�=;Z=��=��=�1=��=.H=��=fB
=^�=�!=�=��=�A=:� =��<"]�<��<ze�<���<I�<Z��<��<b�<���<���<}>�<�|�<^��<���<��<aJ�<�t�<��<���<��<{�< �<�;�<2U�<m�<D��<��<���<���<�ό<J��<���<| �<� z<[@r<�`j<��b<y�Z<��R<N�J<C<@;<�l3<��+<=�#<�<�<<*z<��<O�;���;@�;K��;���;���;tc�;�W�;�`�;��b;\iE;9(;��
;��:%�: &R:���9��r�7����9l�	����F⺯���%���?��GY��dr�s���^���	���We���괻L8��:N˻�+ֻ��໿?뻷v���v�����2k	������D0�|������$�c8(�=B,�*70�4��7��;��L?���B��sF�[�I�3bM���P�M T�oW���Z���]��"a�pMd�Xpg���j���m�®p���s���v�T�y��|���aG�����0�������ト���Y`��>͌�A9��������[x�������H���������{���ߚ�_C������_	���k���͡�0�����L����V���������~���ᬼ�D��X�������o��0ӳ��6��Ú�������b��Ǻ��+��͐���  �  z�N=�N=<`M=��L=��K=VDK=��J=��I=O%I=�oH=��G=vG=�LF=I�E=@�D=(D=rpC=��B=6 B=fGA=	�@=�?=V?=�]>=��==Z�<=.&<=g;=Ʀ:=��9=#9=�_8=7=��6=k6=�D5=qz4=��3=�2=�2=3@1=�l0=��/=B�.=�-=/-=,$,=@+=|X*=sm)=�~(='�'=��&=��%=��$=��#=�"=y�!=tn =�U=�7=W=��=��=�=A=N�=S�=$Z=��=ϛ=�1=Z�=�G=q�= B
=�=�!=��=��=�A=�� =���<�\�<���<Je�<���<I�<N��<��<0b�<ڱ�<7��<�>�<H}�<Ŷ�<��<0�<�J�<7u�<���<��<�<��<C �<�;�<JU�<m�<X��<��<���<̽�<Oό<�߈<%��< �<�z<{?r<�_j<�b<f�Z<��R<m�J<:C<�?;<l3<��+<��#<�<�<<4z<�<��;R��;pA�; ��;V��;���;�e�;�Y�;Cc�;�c;�mE;-(;��
;y��:�(�:c,R:���9��r�����&:l�Ձ��6I�ܳ���%��?��JY�zhr������������$g��촻�9��PO˻�,ֻi��
@��v���v��}���j	�Q����/�˔����$�[7(�PA,�C60�4�;�7��;�L?��B��rF��I��aM���P�, T�;oW�6�Z��]�&#a��Md�8qg�Ìj���m���p���s���v�K�y�֭|�����G��(���1��<���*��냈���S`��#͌�9��1�������w������]H��*���X���z��ߚ��B��1���	��k���͡��/�����B����V��%�������~���ᬼSE��¨��J���o���ӳ�m7��/���3���5c���Ǻ�&,������  �  R�N=fN=#`M=��L=��K=oDK=яJ=��I=�%I=�oH=��G=�G=RMF=��E=��D=c(D=�pC=ݸB=� B=�GA=?�@=9�?=y?=�]>=��==S�<=&<=�f;=��:=F�9=�"9=<_8=p�7=g�6=6=MD5=z4=C�3=��2=[2=�?1=dl0=��/=�.=�-=+-=7$,=@+=�X*=�m)=�~(=n�'=ݕ&=�%=�$=�#=y�"=ǁ!=�n =AV=�7=�=��=��=�=A=@�=<�=�Y=l�=��=h1=�=�G=�=�A
=��=!=9�=4�=LA=�� =��<I\�<x��<�d�<T��<�H�<Z��<�<�b�<3��<���<e?�<�}�<u��<���<��<�K�<�u�<2��<���<��<P�<� �<<�<�U�<4m�<X��<䗘<F��<���<�Ό<s߈<��<h��<7z<�=r<7^j<�b<�Z<6�R<&�J<'C<�>;<Vk3<��+<�#<�<=<�z<�<��;��;�C�;���;��;���;�h�;l]�;Mf�;�c;esE;�(;��
;>��:R1�:C9R:\�9�Or�9��.>l�����GM� ����%�?�?�MOY��lr������������si��\�;��Q˻S.ֻs��
A�7w���v��A��mj	���+���.��������$�6(��?,��40��4���7�۟;��J?��B�*rF�Q�I�yaM���P�8 T�foW�ǴZ���]��#a��Nd�-rg���j��m���p��s��v���y�$�|���GH������d1������n��������.`���̌��8��ǣ����aw���ߓ��G����������y��gޚ�JB���������k��a͡��/��ܑ��2����V��P�����,��g⬼�E��P�������p��PԳ�8��盶������c��Ⱥ��,������  �  �N==N=`M=��L=��K=�DK=��J=�I=�%I=CpH=^�G=<G=�MF=�E=$�D=�(D=HqC=J�B=� B= HA=��@=u�?=�?=^>=��==I�<=�%<=�f;=a�:=��9={"9=�^8=�7=��6=�6=�C5=�y4=ԭ3=Q�2=�2=�?1= l0=V�/=��.=�-=%-=K$,=?@+=�X*=�m)=F(=Ќ'=B�&=��%=U�$=��#=�"=4�!==o =�V=K8=�=%�=�=�=A=.�=!�=�Y=/�=8�= 1=��=G=��=(A
=�=� =��=��=�@=6� =H��<�[�<���<�d�<��<�H�<q��<<�<�b�<���<H��<@�<�~�<i��<���<��<�L�<�v�<&��<�·<��<��<O!�<�<�<�U�<Ym�<Q��<ϗ�<���<!��<EΌ<�ވ<��<���<_z<�;r<[\j<{}b<�Z<T�R<`�J<�C<'=;<^j3<6�+<�#<S<=<�z<"�<��;w��;�F�;���;���;Ɗ�;�l�;�a�;Tj�;�c;[{E;#(;��
;���:W;�:HHR:(�9��q�Uz���>l������Q���J�%���?�)UY��sr�����ؽ�������l���񴻎>��wS˻40ֻ����A�ow���v��ٟ��i	�����X-������$�44(��=,��20��4���7�/�;�SI?���B�qF��I��`M�0�P�F T��oW�>�Z�W�]��$a�KPd��sg���j���m��p�̺s��v�w�y�Ұ|�����H��L����1��ۣ�����������_���̌�H8��9���P���v��ߓ��F����������x��uݚ�^A��֤�����yj���̡�D/����������V��m���k������⬼uF���������q��Hճ��8��ܜ��� ���d���Ⱥ�I-������  �  ��N=	N=�_M=��L=��K=�DK=0�J=\�I=*&I=�pH=ӺG=�G=TNF=��E=��D=e)D=�qC=ƹB=SB=cHA=ߎ@=��?=�?=%^>=��===�<=�%<=zf;=�:=��9="9=_^8=��7=i�6=6=LC5=y4=O�3=��2=�2=D?1=�k0=�/=ν.=��-=&-=[$,=c@+=Y*=8n)=�(=5�'=��&=�%=�$=�#=t�"=��!=�o =W=�8=,=l�=�=�=A="�=��=�Y=��=Ӛ=�0=�=}F=��=�@
=x�=�=�=�=9@=�� =j��<�Z�<I��<d�<���<�H�<u��<s�<Cc�<A��<���<�@�<��<a��<���< �<�M�<�w�<(��<�÷<Y�<��<�!�<�<�<$V�<�m�<S��<���<���<���<�͌<�݈<��<���<7z<�9r<�Yj<3{b<ٝZ<7�R<g�J<�C<�;;<i3<?�+<��#<<5=<\{<�<�
�;d��;J�;���;,��;f��;�q�;�f�;no�;;c;d�E;�(;j�
;���:{F�:�YR:"?�9�mq�Nu���Al�����HY����%��?�\Y�{r�ʙ����������kp�������A��V˻m2ֻ���C��w��dv�����1i	�������+�Y��#���$��1(��;,��00��4���7�D�;��G?�?�B��oF�z�I�U`M���P�2 T��oW�ڵZ�q�]�:&a��Qd�yug���j���m��p���s��v���y�ʲ|�i���I������u2��[������/������_��>̌��7����������u��ޓ��E��~�������w��bܚ�g@��裝�����i��N̡��.��]����󥼳V���������%����㬼=G���������r��Zֳ� :��흶�����e���ɺ�.�������  �  ��N=�N=�_M=��L=��K=�DK=j�J=��I=�&I=qH=V�G=@G=�NF==�E=@�D=�)D=TrC=O�B=�B=�HA=7�@=��?=?=@^>=��==&�<=�%<=Cf;=å:=@�9=�!9=�]8=��7=��6=v6=�B5=�x4=��3=X�2=2=�>1=xk0=̕/=��.=��-= -=j$,=�@+=LY*=}n)=�(=��'==�&=��%=n�$=��#=�"=L�!=4p =�W=9=�=��=K�=/�="A=�=ʭ=NY=��=f�=0=��=�E=A�=�?
=��=3=Z�=i�=�?="� =i��< Z�<���<�c�<m��<�H�<���<��<�c�<г�<���<�A�<���<l��<���<3!�<�N�<y�<C��<�ķ<C�<��<�"�<�=�<xV�<�m�<I��<f��<J��<��<�̌<݈<��<o��<�z<D7r<VWj<�xb<_�Z<�R<_�J<�C<:;<�g3<P�+<��#<�<L=<�{<Ҿ<��;v��;�M�;.�;�¼;;��;�v�;�k�;�t�;$%c;j�E;�&(;��
;���:�Q�:�mR:�X�9��p��u���El������`���� &���?�	dY�%�r����eƑ������t������E��Y˻�4ֻs�� D뻻x��_v��*��qh	������(*�}������$��/(�=9,�5.0�Q4���7��;��E?���B��nF���I��_M���P�7 T�_pW�|�Z�j�]��'a�LSd�9wg���j��m�K�p�o�s�k�v�սy��|�R���J������3��Τ��0��e���u򉼞_���ˌ�E7��塏�����t��ݓ��D��O���[���v��Eۚ�V?��ܢ�����h���ˡ�`.��������V��깨�-������T䬼H��髯�����s���׳�Z;���������f���ʺ��.��w����  �  C�N=�N=�_M=v�L=��K=�DK=��J=��I=�&I=�qH=ͻG=�G=sOF=јE=��D=�*D=�rC=ԺB=DB=:IA=��@==�?=3?=c^>=��==�<=�%<=	f;=}�:=��9=/!9=_]8=m�7=I�6=�
6=B5=�w4=4�3=��2=�2=n>1=%k0=��/=n�.=��-=-=�$,=�@+=�Y*=�n)=k�(=�'=��&=�%=��$=?�#=��"=Ճ!=�p =X=}9=�=��=|�=I�=/A=��=��=Y=/�=�=�/=��=CE=��=)?
=�=~=��=��=�>=�� =e��<AY�< ��< c�<"��<�H�<���<��<d�<l��<}��<�B�<���<���<��<k"�<P�<Fz�<k��<�ŷ</�<a�<3#�<�=�<�V�<�m�<D��<7��<ᩔ<���<8̌<I܈<��<P��<�z<�4r<�Tj<-vb<�Z<��R<'�J<C<h8;<sf3<A�+<4�#<<y=<X|<��<i�;���;LQ�;)�;|Ǽ;?��;|�;3q�;�y�;�/c;�E;�/(;��
;^��:�]�: R:v�9Jmp�7q��Il�L����f�1���&���?��kY�0�r�y����ʑ������x�������H��'\˻;7ֻ,�໌E�Hy��Uv������g	���&��}(�������6$�T-(��6,��+0�4�t�7�!�;�D?���B�9mF���I��^M�)�P�8 T��pW�C�Z�[�]��(a��Td�yg���j��m���p���s���v��y�5�|�v���K�������3��A����������g�\_��~ˌ��6��2����
���s��
ܓ�yC��/���$��mu��#ښ�:>��록�=��9h��'ˡ��-��ʐ�����V��!������8���嬼�H��謯�����t���س�|<��F������g���˺��/��1����  �   �N=kN=�_M=h�L=��K=EK=ҐJ=9�I=:'I=�qH=@�G=HG=�OF=Y�E=n�D=+D=ksC=O�B=�B=�IA=�@=��?=d?=}^>=��==�<=n%<=�e;=5�:=��9=� 9=�\8=�7=��6=P
6=�A5=\w4=��3=R�2=+2=>1=�j0=J�/=C�.=��-=-=�$,=�@+=�Y*=o)=��(=�'=(�&=��%=~�$=Ě#=!�"=X�!=9q ={X=�9=6=9�=��=a�=4A=��=��=�X=��=��=/=t�=�D=�=>
=m�=�=�=.�=m>=� =~��<yX�<X��<�b�<���<[H�<���</�<�d�<���<%��<~C�<|��<���<��<�#�<(Q�<Y{�<o��<�Ʒ<�<�<�#�<}>�<W�<n�<1��<��<���<��<�ˌ<}ۈ<��<O��<`z<e2r<�Rj<�sb<��Z<t�R<*�J<SC<�6;<@e3<S�+<��#<+<�=<�|<m�<��;?��;�T�;	�;�˼;͝�;ˀ�;Lv�;�~�;#9c;	�E;8(;_;��:�i�:�R:��9Zp��n��LLl�%����m����&�y�?�lrY��r�v����Α�3���3|��- ���K���^˻�9ֻ�໮F뻪y��jv��L��g	���٪�'�����/$�)+(��4,��)0��
4�h�7�>�;�EB?���B��kF�z�I�V^M���P�J T��pW��Z�]�]�*a�oVd��zg���j��m��p���s���v�O�y�$�|�S��jL��G���@4�������������i�._��#ˌ�.6������'
�� s��ۓ�qB�������^t��ٚ�>=�����d���g���ʡ��-���������V��S�����������嬼�I��̭������u���ٳ��=��f������h���̺��0��唽��  �  ��N=AN=y_M=a�L=��K=EK=��J=n�I=�'I=CrH=��G=�G=lPF=ԙE=��D=�+D=�sC=��B=B=�IA=*�@=��?=�?=�^>=��==��<=L%<=�e;=�:=4�9=g 9=�\8={�7=F�6=�	6=A5=�v4=9�3=��2=�2=�=1=�j0=�/= �.=��-=-=�$,=�@+=�Y*=Wo)=�(=ڎ'=��&=��%=�$=6�#=��"=̈́!=�q =�X==:=�=n�=ָ=s�=4A=��=Y�=�X=��=C�=�.=��=3D=y�=�=
=ڰ=I=y�=��=�==�� =���<�W�<���<Jb�<���<GH�<���<^�<�d�<l��<���<;D�<N��<h��<��<r$�<R�<K|�<O��<kǷ<��<��<S$�<�>�<QW�<$n�<5��<ז�<9��<���<�ʌ<�ڈ<.�<j��<Zz<�0r<�Pj<�qb<��Z<��R<|�J<�	C<�5;<#d3<��+<�#<�<�=<}<�<��;ǯ�;�W�;|�;pϼ;���;��;;z�;)��;5Ac;��E;�?(;�;V	�: r�:�R:��9a�o�Km��sPl�񝬺Rt⺵��P&��?�yY��r�䩅�.ґ�tĝ����M���N��ua˻�;ֻ��໛G�Wz��+v�����f	������%�j��Z��x
$�>)(��2,��'0��4���7���;��@?�;�B��jF���I��]M���P�; T�WqW�g�Z�2�]�*+a��Wd�M|g�>�j��m���p���s���v�'�y��|���1M�������4�����
��˄��^�_���ʌ��5��
���~	��7r��=ړ��A��$��� ��js��+ؚ�g<��4�������f�� ʡ�.-��c������V������L��6���I欼jJ����������v���ڳ��>��K������i��fͺ�P1��w����  �  ��N=N=a_M=\�L=��K=9EK="�J=��I=�'I=rH=�G=G=�PF=0�E=6�D=�+D=.tC=�B=bB=.JA=f�@=��?=�?=�^>=¡==��<=2%<=xe;=��:=��9=! 9=9\8=&�7=��6={	6=�@5=�v4=ߪ3=��2=~2=v=1=Tj0=ߔ/=��.=p�-=-=�$,=A+=Z*=�o)=N�(=�'=ߘ&=L�%=D�$=��#=�"=�!=�q =+Y=u:=�=��=��=��=5A=��=>�=qX=X�=�=g.=��=�C=�=�=
=g�=�=�=9�=�==D� =#��<>W�<b��<�a�<f��<;H�<���<��<e�<ӵ�<0 �<�D�<��<
��<���<&%�<�R�<�|�<���<ȷ<O�<E�<�$�<.?�<�W�<6n�<1��<���<�<��<�ʌ<=ڈ<��<���<�z</r<�Nj<epb<?�Z<&�R<6�J<�C<�4;<3c3<�+<��#<�<�=<h}<��<��;ڱ�;�Y�;�;4Ҽ;���;5��;Q}�;Y��;Gc;ԮE;�D(;{;��:�x�:ثR:ɮ�98^o��k��Tl������y⺖��&��?��}Y���r�����Ց��Ɲ�w���u���P��Ec˻/=ֻ�໎H��z��v��ޝ�f	�J����$�t����#	$��'(�B1,�;&0��4�^�7�H�;��??�9�B�&jF�1�I�O]M�z�P�2 T��qW��Z���]��+a��Xd�r}g�c�j�V�m��p�b�s�^�v�n�y�_�|����M��Z�65��q���D������T��^���ʌ��5������	���q���ٓ��@��t���m���r���ך��;������<��uf���ɡ��,��(���~�W��������������欼�J��&���Q��vw��^۳�Y?���������Oj���ͺ��1��啽��  �  w�N=
N=]_M=U�L=��K=EEK=.�J=��I=�'I=�rH=$�G==G=�PF=f�E=u�D=$,D=ltC=B�B=�B=ZJA=��@=��?=�?=�^>=��==��<=(%<=ee;=��:=��9=�9=\8=�7=��6=>	6=z@5=Tv4=��3=`�2=M2=O=1=.j0=Δ/=�.=m�-=	-=�$,=A+=&Z*=�o)=k�(=K�'=�&=��%=�$=ƛ#=!�"=V�!=*r =[Y=�:=�=��=�=��=6A=��=5�=[X=>�=֘=7.=l�=�C=��=J=
=%�=�=͂=��=U==� =���<�V�<(��<�a�<S��< H�<���<��<3e�<��<| �<!E�<P��<���<(��<�%�<JS�<t}�<n��<rȷ<��<��<�$�<P?�<�W�<9n�<$��<���<֨�<���<1ʌ<�و<#�<L��<�z<�-r<�Mj<Job<F�Z<;�R<G�J<�C<�3;<�b3<��+<��#<�<�=<�}<��<��;ò�;Q[�;��;Լ;���;��;�;>��;yKc;��E;�H(;�;�:�|�:��R:��9�Zo��i���Tl�/���|⺵��P&�>�?��Y�(�r�W����֑��ȝ����;��2R��gd˻D>ֻw���H��z��Pv����e	������9$����G��,$��&(�^0,�Q%0��4�f�7�y�;��>?���B��iF���I�]M�[�P�S T��qW� �Z�9�]��,a�VYd�,~g�N�j�-�m���p�C�s�J�v�n�y�9�|����N����m5������^��儈�b��^��zʌ�T5��]������Eq��3ٓ�q@��������Dr��	ך�Q;��6������>f���ɡ��,�����}�W���������Ă��笼@K����������w���۳��?��~���$���j��kκ�)2��:����  �  n�N=�N=P_M=S�L=�K=NEK=4�J=��I=�'I=�rH=)�G=FG=QF=v�E=��D=4,D=�tC=F�B=�B=gJA=��@=
�?=�?=�^>=��==��<=%<=Te;=��:=��9=�9=�[8=�7=��6=+	6=m@5=>v4=��3=O�2=C2=F=1=j0=Ɣ/=ݼ.=b�-=-=�$,=A+=,Z*=�o)=t�(=\�'=�&=��%=��$=֛#=1�"=l�!=7r =XY=�:=�=��=
�=��=>A=��=,�=JX=2�=Ƙ=*.=^�=�C=��=1=
=�=�=��=��=?==� =���<�V�<��<�a�<K��<$H�<֮�<��<Le�<��<� �<4E�<R��<���<K��<�%�<hS�<�}�<���<yȷ<��<��<%�<[?�<�W�<Jn�<��<���<���<㹐<ʌ<�و<	�<0��<�z<�-r<�Mj<�nb<�Z<�R<�J<�C<�3;<�b3<G�+<Y�#<�<�=<�}< �<��;��;�[�;��;iԼ;���;���;3��;ӈ�;�Lc;�E;.I(;�;��:L�:�R:���9�Ao�tj�� Xl�7���v}����.&�h�?���Y�<�r�뮅�ב��ɝ�I������|R���d˻�>ֻ���xI�{��`v������e	���L��$�F��H���$��&(�0,�%0�S4�.�7���;��>?���B�riF���I�]M�5�P�] T��qW�]�Z�^�]��,a��Yd�Y~g���j�M�m�Y�p���s���v���y�Z�|�E��2N�����5������x��너�]��^��uʌ�:5��F������3q��1ٓ�M@��⦖����&r���֚�=;��0������.f��dɡ��,�����k�W��ں�����؂��)笼PK����������w��ܳ��?������B���j���κ�:2��[����  �  w�N=
N=]_M=U�L=��K=EEK=.�J=��I=�'I=�rH=$�G==G=�PF=f�E=u�D=$,D=ltC=B�B=�B=ZJA=��@=��?=�?=�^>=��==��<=(%<=ee;=��:=��9=�9=\8=�7=��6=>	6=z@5=Tv4=��3=`�2=M2=O=1=.j0=Δ/=�.=m�-=	-=�$,=A+=&Z*=�o)=k�(=K�'=�&=��%=�$=ƛ#=!�"=V�!=*r =[Y=�:=�=��=�=��=7A=��=6�=\X=?�=ט=9.=n�=�C=��=L=
='�=�=Ђ=��=X==� =���<�V�</��<�a�<Z��<'H�<Ʈ�<��<9e�<	��<� �<%E�<S��<���<)��<�%�<JS�<s}�<l��<pȷ<��<|�<�$�<K?�<�W�<4n�<��<���<Ѩ�<���<-ʌ<�و< �<J��<�z<�-r<�Mj<Lob<I�Z<@�R<M�J<�C<�3;<�b3<��+<��#<�<�=<�}<��<��;Ӳ�;_[�;��;Լ;���;��;}�;9��;gKc;��E;}H(;�;��:�|�:ٯR:$��9`io��k���Ul������|�����&�v�?�9�Y�Z�r�o����֑��ȝ����L��AR��td˻P>ֻ����H��z��Wv��ŝ��e	������:$����H��-$��&(�^0,�R%0��4�f�7�z�;��>?���B��iF���I�]M�[�P�S T��qW� �Z�9�]��,a�VYd�,~g�N�j�-�m���p�C�s�J�v�n�y�9�|����N����m5������^��儈�b��^��zʌ�T5��]������Eq��3ٓ�q@��������Dr��	ך�Q;��6������>f���ɡ��,�����}�W���������Ă��笼@K����������w���۳��?��~���$���j��kκ�)2��:����  �  ��N=N=a_M=\�L=��K=9EK="�J=��I=�'I=rH=�G=G=�PF=0�E=6�D=�+D=.tC=�B=bB=.JA=f�@=��?=�?=�^>=¡==��<=2%<=xe;=��:=��9=! 9=9\8=&�7=��6={	6=�@5=�v4=ߪ3=��2=~2=v=1=Tj0=ߔ/=��.=p�-=-=�$,=A+=Z*=�o)=N�(=�'=ߘ&=L�%=D�$=��#=�"=�!=�q =+Y=u:=�=��=��=��=6A=��=@�=rX=Z�=�=i.=��=�C=�=�=
=k�=�=�=?�=�==J� =0��<KW�<p��<b�<s��<HH�<Į�<��<e�<ܵ�<8 �<�D�<��<��<���<'%�<�R�<�|�<���<ȷ<H�<=�<�$�<$?�<�W�<,n�<&��<���<ꨔ<��<~ʌ<6ڈ<��<���<�z</r<�Nj<hpb<F�Z</�R<B�J<�C<�4;<Fc3<��+<��#<�<�=<}}<��<�;���;�Y�;�;DҼ;���;8��;N}�;N��;�Fc;��E;~D(;3;��:�w�:E�R:n��9dzo�"o���Ul������z�
���&�x�?�I~Y���r�����>Ց�ǝ���������P��^c˻F=ֻ�໠H��z��!v����f	�N����$�v����%	$��'(�C1,�<&0��4�_�7�I�;��??�:�B�&jF�1�I�O]M�z�P�2 T��qW��Z���]��+a��Xd�r}g�c�j�V�m��p�b�s�^�v�n�y�_�|����M��Z�65��q���D������T��^���ʌ��5������	���q���ٓ��@��t���m���r���ך��;������<��uf���ɡ��,��(���~�W��������������欼�J��&���Q��vw��^۳�Y?���������Oj���ͺ��1��啽��  �  ��N=AN=y_M=a�L=��K=EK=��J=n�I=�'I=CrH=��G=�G=lPF=ԙE=��D=�+D=�sC=��B=B=�IA=*�@=��?=�?=�^>=��==��<=L%<=�e;=�:=4�9=g 9=�\8={�7=F�6=�	6=A5=�v4=9�3=��2=�2=�=1=�j0=�/= �.=��-=-=�$,=�@+=�Y*=Wo)=�(=ڎ'=��&=��%=�$=6�#=��"=̈́!=�q =�X=>:=�=o�=׸=t�=5A=��=[�=�X=��=F�=�.= �=7D=~�=�=
=�=P=��=��=�==�� =���<�W�<���<]b�<���<ZH�<���<n�<�d�<y��<���<ED�<V��<n��<��<s$�<R�<H|�<J��<cǷ<��<��<G$�<�>�<CW�<n�<&��<Ȗ�<+��<|��<�ʌ<�ڈ<&�<d��<Qz<�0r<�Pj<�qb<��Z<��R<��J<�	C<�5;<=d3<��+<1�#<<�=<!}</�<��;���;�W�;��;�ϼ;Ρ�;��;6z�;��;Ac;��E;4?(;\;k�:�p�:ӜR:W��91�o�nr��Sl�A����u�Y���&���?��yY�m�r�%���iґ��ĝ����z���N���a˻�;ֻ��໴G�lz��=v�����f	������%�m��]��{
$�@)(��2,��'0��4���7���;��@?�;�B��jF���I��]M���P�; T�WqW�g�Z�2�]�*+a��Wd�M|g�>�j��m���p���s���v�'�y��|���1M�������4�����
��˄��^�_���ʌ��5��
���~	��7r��=ړ��A��$��� ��js��+ؚ�g<��4�������f�� ʡ�.-��c������V������L��6���I欼jJ����������v���ڳ��>��K������i��fͺ�P1��w����  �   �N=kN=�_M=h�L=��K=EK=ҐJ=9�I=:'I=�qH=@�G=HG=�OF=Y�E=n�D=+D=ksC=O�B=�B=�IA=�@=��?=d?=}^>=��==�<=n%<=�e;=5�:=��9=� 9=�\8=�7=��6=P
6=�A5=\w4=��3=R�2=+2=>1=�j0=J�/=C�.=��-=-=�$,=�@+=�Y*=o)=��(=�'=(�&=��%=~�$=Ś#=!�"=X�!=9q =|X=�9=6=:�=��=b�=6A=��=��=�X=��=��=/=y�=�D=�=�>
=u�=�=�=8�=w>= � =���<�X�<o��<�b�<���<qH�<®�<C�<�d�<��<4��<�C�<���<���<��<�#�<&Q�<U{�<h��<�Ʒ<
�<�<�#�<m>�<W�<�m�<��<���<u��<�<vˌ<qۈ<��<H��<Vz<`2r<�Rj<�sb<ʖZ<��R<?�J<lC<�6;<`e3<u�+<��#<P<�=<�|<��<�;w��;�T�;(	�;�˼;ޝ�;р�;Fv�;�~�;�8c;��E;�7(;� ;���:Xh�:0�R:D��9>p�u��Ol�����Fo⺕���&�5�?�sY���r�Ŧ���Α�w���q|��e ���K��_˻�9ֻ(���F��y���v��U��'g	���ߪ�'�����2$�,+(��4,��)0��
4�i�7�?�;�FB?���B��kF�z�I�V^M���P�K T��pW��Z�^�]�*a�oVd��zg���j��m��p���s���v�O�y�$�|�S��jL��G���@4�������������i�._��#ˌ�.6������'
�� s��ۓ�qB�������^t��ٚ�>=�����d���g���ʡ��-���������V��S�����������嬼�I��̭������u���ٳ��=��f������h���̺��0��唽��  �  C�N=�N=�_M=v�L=��K=�DK=��J=��I=�&I=�qH=ͻG=�G=sOF=јE=��D=�*D=�rC=ԺB=DB=:IA=��@==�?=3?=c^>=��==�<=�%<=	f;=}�:=��9=/!9=_]8=m�7=I�6=�
6=B5=�w4=4�3=��2=�2=n>1=%k0=��/=n�.=��-=-=�$,=�@+=�Y*=�n)=k�(=�'=��&=�%=��$=?�#=��"=փ!=�p =X=}9=�=��=}�=K�=0A= �=��=Y=3�=�=�/=��=IE=��=1?
=�=�=��=��=	?=�� =~��<[Y�<��<:c�<;��<�H�<���<�<!d�<~��<���<�B�<���<���<��<m"�<P�<Az�<c��<�ŷ<"�<R�<"#�<�=�<�V�<�m�<0��<#��<Ω�<r��<(̌<;܈<��<G��<~z<�4r<�Tj<3vb<�Z<��R<?�J<1C<�8;<�f3<h�+<\�#<�<�=<�|<��<��;٪�;�Q�;U�;�Ǽ;S��;|�;-q�;�y�;n/c;��E;/(;W�
;��:\�:|R:�o�9��p�;x���Ll�����h����&���?�alY��r�Ѣ���ʑ�K����x�������H��Y\˻g7ֻS�໮E�fy��nv������g	���-���(�������9$�W-(��6,��+0�4�u�7�"�;�D?���B�:mF���I��^M�)�P�9 T��pW�C�Z�[�]��(a��Td�yg���j��m���p���s���v��y�5�|�v���K�������3��A����������g�\_��~ˌ��6��2����
���s��
ܓ�yC��/���$��mu��#ښ�:>��록�=��9h��'ˡ��-��ʐ�����V��!������8���嬼�H��謯�����t���س�|<��F������g���˺��/��1����  �  ��N=�N=�_M=��L=��K=�DK=j�J=��I=�&I=qH=V�G=@G=�NF==�E=@�D=�)D=TrC=O�B=�B=�HA=7�@=��?=?=@^>=��==&�<=�%<=Cf;=å:=@�9=�!9=�]8=��7=��6=v6=�B5=�x4=��3=X�2=2=�>1=xk0=̕/=��.=��-= -=j$,=�@+=LY*=}n)=�(=��'==�&=��%=n�$=��#=�"=M�!=4p =�W=9=�=��=M�=1�=$A=�=ͭ=RY=��=j�=0=��=�E=I�=�?
=Ȳ===e�=t�=�?=/� =���<Z�<���<�c�<���<�H�<���<��<�c�<��<���<�A�<���<t��<���<4!�<�N�<y�<;��<�ķ<5�<}�<u"�<o=�<dV�<�m�<4��<Q��<7��<�<�̌<݈<��<e��<�z<>7r<VWj<�xb<l�Z<�R<w�J<C<,:;<�g3<x�+<��#<�<v=<�{<��<=�;���;�M�;[�;�¼;P��;�v�;�k�;�t�;�$c;�E;i&(;��
;t��:8P�:{jR:�Q�9)q��|��IIl������b�����&�n�?��dY��r�q����Ƒ�򸝻�t������PE��IY˻5ֻ���CD��x��yv��5��zh	������.*��������$��/(�@9,�7.0�S4���7��;��E?���B��nF���I��_M���P�8 T�_pW�|�Z�j�]��'a�LSd�:wg���j��m�K�p�o�s�k�v�սy��|�R���J������3��Τ��0��e���u򉼞_���ˌ�E7��塏�����t��ݓ��D��O���[���v��Eۚ�V?��ܢ�����h���ˡ�`.��������V��깨�-������T䬼H��髯�����s���׳�Z;���������f���ʺ��.��w����  �  ��N=	N=�_M=��L=��K=�DK=0�J=\�I=*&I=�pH=ӺG=�G=TNF=��E=��D=e)D=�qC=ƹB=SB=cHA=ߎ@=��?=�?=%^>=��===�<=�%<=zf;=�:=��9="9=_^8=��7=i�6=6=LC5=y4=O�3=��2=�2=D?1=�k0=�/=ν.=��-=&-=[$,=c@+=Y*=8n)=�(=5�'=��&=�%=�$=�#=t�"=��!=�o =W=�8=-=m�=�=�=!A=%�=��=�Y=��=ؚ=�0=�=�F=��=�@
=��=�=�="�=E@=�� =���<�Z�<d��<9d�<���<�H�<���<��<Xc�<S��<��<�@�<��<i��<���< �<�M�<�w�< ��<}÷<L�<��<�!�<�<�<V�<qm�<?��<���<���<~��<�͌<�݈<��<}��<+z<�9r<�Yj<9{b<�Z<I�R<~�J<�C<�;;<(i3<e�+<��#<B<^=<�{<�<�;���;HJ�;���;M��;z��;�q�;�f�;Zo�;�c;�E;(;��
;o��:E�:�VR:�8�92�q�Q|��El�V���[�����%���?��\Y��{r�"���B�״���p��;���B��:V˻�2ֻ���3C�x��~v�����;i	�������+�]��'���$��1(��;,��00��4���7�E�;��G?�@�B��oF�{�I�U`M���P�2 T��oW�ڵZ�q�]�:&a��Qd�yug���j���m��p���s��v���y�ʲ|�i���I������u2��[������/������_��>̌��7����������u��ޓ��E��~�������w��bܚ�g@��裝�����i��N̡��.��]����󥼳V���������%����㬼=G���������r��Zֳ� :��흶�����e���ɺ�.�������  �  �N==N=`M=��L=��K=�DK=��J=�I=�%I=CpH=^�G=<G=�MF=�E=$�D=�(D=HqC=J�B=� B= HA=��@=u�?=�?=^>=��==I�<=�%<=�f;=a�:=��9={"9=�^8=�7=��6=�6=�C5=�y4=ԭ3=Q�2=�2=�?1= l0=V�/=��.=�-=%-=K$,=?@+=�X*=�m)=F(=Ќ'=C�&=��%=V�$=��#=�"=4�!==o =�V=K8=�=&�=�=�=A=0�=$�=�Y=2�=<�=1=��=G=��=/A
=&�=� =��=��=�@=A� =^��<�[�<��<�d�</��<�H�<���<P�<�b�<���<W��<)@�<�~�<p��<���<��<�L�<�v�< ��<�·<u�<��<@!�<o<�<�U�<Gm�<?��<���<<��<7Ό<�ވ<��<}��<Uz<�;r<[\j<�}b<!�Z<d�R<t�J<�C<D=;<~j3<Y�+<>�#<x<4=<{<D�<��;���;�F�;��;��;؊�;�l�;�a�;Bj�;�c;{E;�(;L�
;���::�:�ER:8"�9�.r�����Bl�4����S�λ��%���?��UY�1tr�F���!���ܰ���l�����>���S˻[0ֻ���B뻊w���v�����i	���	��]-������$�64(��=,��20��4���7�0�;�TI?���B�qF��I��`M�0�P�F T��oW�>�Z�W�]��$a�KPd��sg���j���m��p�̺s��v�w�y�Ұ|�����H��L����1��ۣ�����������_���̌�H8��9���P���v��ߓ��F����������x��uݚ�^A��֤�����yj���̡�D/����������V��m���k������⬼uF���������q��Hճ��8��ܜ��� ���d���Ⱥ�I-������  �  R�N=fN=#`M=��L=��K=oDK=яJ=��I=�%I=�oH=��G=�G=RMF=��E=��D=c(D=�pC=ݸB=� B=�GA=?�@=9�?=y?=�]>=��==S�<=&<=�f;=��:=F�9=�"9=<_8=p�7=g�6=6=MD5=z4=C�3=��2=[2=�?1=dl0=��/=�.=�-=+-=7$,=@+=�X*=�m)=�~(=n�'=ݕ&=�%=�$=�#=z�"=ǁ!=�n =AV=�7=�=��=��=�=A=B�=>�=�Y=o�=��=l1=�=�G=�=�A
=��="!=A�=<�=TA=�� =)��<\\�<���<�d�<g��<I�<l��<�<�b�<A��<���<o?�<�}�<{��<���<��<�K�<�u�<,��<���<��<D�<� �<	<�<zU�<%m�<I��<՗�<9��<t��<�Ό<h߈<��<a��<.z<�=r<7^j<�b<�Z<C�R<7�J<;C<�>;<qk3<�+<��#<�<!=<�z<��<��;D��;�C�;���;5��;���;�h�;g]�;?f�;�c;"sE;s(;��
;S��:L0�:	7R:�
�9�wr�\����@l�����N�ķ�\�%���?��OY�qmr�Ӓ��ẑ�D����i����;��4Q˻s.ֻ���#A�Mw���v��I��sj	���0���.��������$�6(��?,��40��4���7�ܟ;��J?��B�+rF�R�I�zaM���P�8 T�goW�ǴZ���]��#a��Nd�-rg���j��m���p��s��v���y�$�|���GH������d1������n��������.`���̌��8��ǣ����aw���ߓ��G����������y��gޚ�JB���������k��a͡��/��ܑ��2����V��P�����,��g⬼�E��P�������p��PԳ�8��盶������c��Ⱥ��,������  �  z�N=�N=<`M=��L=��K=VDK=��J=��I=O%I=�oH=��G=vG=�LF=I�E=@�D=(D=rpC=��B=6 B=fGA=	�@=�?=V?=�]>=��==Z�<=.&<=g;=Ʀ:=��9=#9=�_8=7=��6=k6=�D5=qz4=��3=�2=�2=3@1=�l0=��/=B�.=�-=/-=,$,=@+=|X*=sm)=�~(='�'=��&=��%=��$=��#=�"=y�!=tn =�U=�7=W=��=��=�=A=O�=T�=&Z=��=ћ=�1=]�=�G=u�=$B
=�=�!=��=��=�A=�� =���<�\�<���<We�<���<I�<Z��<��<;b�<��<@��<�>�<N}�<ɶ�<��<1�<�J�<4u�<~��<��<�<��<: �<�;�<@U�<m�<N��<���<���<ý�<Gό<�߈<��<	 �<�z<x?r<�_j<�b<m�Z<��R<y�J<IC<�?;<+l3<Û+<�#<�<=<Iz<��<�;r��;�A�;6��;g��;ƃ�;�e�;�Y�;9c�;vc;dmE;�(;��
;ӱ�:�'�:�*R:p��9��r�2����;l�Â��!J�P��8�%���?�BKY��hr�'���B���Ī��Gg��;촻:��jO˻�,ֻ}��@��v���v������j	�U����/�͔����
$�\7(�QA,�D60�4�;�7��;�L?��B��rF��I��aM���P�, T�;oW�6�Z��]�&#a��Md�8qg�Ìj���m���p���s���v�K�y�֭|�����G��(���1��<���*��냈���S`��#͌�9��1�������w������]H��*���X���z��ߚ��B��1���	��k���͡��/�����B����V��%�������~���ᬼSE��¨��J���o���ӳ�m7��/���3���5c���Ǻ�&,������  �  ��N=�N=H`M=��L=��K=QDK=��J=��I=$%I=xoH=y�G=@G=�LF=�E=	�D=�'D=;pC=T�B= B==GA=��@=��?=H?=�]>=��==\�<=;&<=g;=�:=��9=D#9=�_8=��7=��6=�6=�D5=�z4=Ԯ3=C�2=�2=Z@1=�l0=/=O�.='�-=(-=*$,=�?+=hX*=Vm)=�~(=��'=^�&=��%=V�$=��#=�"=9�!=An =�U=�7=4=��=��=�=A=M�=d�=<Z=��=��=�1=��=0H=��=hB
=`�=�!=�=��=�A==� =��<)]�<&��<�e�<���<I�<a��<��<"b�<���<���<�>�<�|�<`��<���<��<aJ�<�t�<��<���<��<w�< �<�;�<-U�<m�<?��<��<���<���<~ό<F��<���<z �<� z<Y@r<�`j<��b<|�Z<��R<T�J<C<#@;<�l3< �+<G�#<�<�<<5z<��<b�;��;'@�;V��;���;Á�;vc�;�W�;�`�;�b;CiE;(;��
;���:�$�:O%R:��9*�r�����:l�����!G���@�%���?��GY�,er�����t������je���괻Z8��GN˻ ,ֻ����?뻿v�� w�����5k	������F0�}������$�c8(�=B,�*70�4��7��;��L?���B��sF�[�I�3bM���P�M T�oW���Z���]��"a�pMd�Xpg���j���m�®p���s���v�T�y��|���aG�����0�������ト���X`��>͌�A9��������[x�������H���������{���ߚ�_C������_	���k���͡�0�����L����V���������~���ᬼ�D��X�������o��0ӳ��6��Ú�������b��Ǻ��+��͐���  �  ��N=�N=�XM=7�L=L�K=:K=|�J=��I=FI=�aH=��G=��F= <F=!�E=��D=fD=�ZC=,�B=S�A=-A=r@=r�?=�>=�<>=�~==�<=��;=�>;=�|:=��9=X�8=�/8=�h7=��6=�5=5=Y?4=q3=נ2=��1=��0=G$0=�K/= p.=6�-=Q�,=n�+=W�*=��)=)=c(=�&'=y-&=�/%=�-$=='#=�"=!=�=��=\�=ݓ=Gg=s4=�=+�=st=�&=Q�=�v=q=�=�:=P�=hE=��	=�5=�==�o=w�=�# =w��<4��<��<��<��<(��<���<�^�<��<�<e�<C��<4��<J7�<�s�<=��<���<�<5@�<=k�<ȓ�<���<�ݫ<	��<��<�<�<�X�<xs�<Ќ�<Y��<���<Pӈ<g�<6��<�)z<NUr<k�j<�b<.�Z<�S<�<K<epC< �;<��3<6,<�W$<f�<��<�(<�v<U��;LG�;��;���;���;.��;N��;���;˂;h;��J;I|-;��;r�:2V�:�Wk:: �9=q:8�;Ź��O�'睺6JӺc� ���7�cQ�tj��W��$q���W��v	��܆��4λ��ƻ��ѻ�aܻ �滄�@��Ls��B����Q��d�������"��G&�p\*��\.��I2�j#6� �9���=��KA�o�D�*oH��K�H^O�*�R��V�;pY�.�\�l�_�n+c�Yf�vi�A�l���o��r���u��x���{���~� 瀼�`���؃�O���Æ�.7��u���j��w���J���dg��`Ԑ��@���������}���痼�O��ڶ�� ��	���C螼=M��ȱ��H���z���ޥ�MC��̧��|��q���լ��:��#���[���j��г�s5������ ���f���̺�j3��T����  �  ��N=�N=�XM=/�L=P�K=:K=��J=��I=VI=�aH=ЪG=��F=<F=0�E=�D=yD=�ZC=6�B=c�A=-A=r@=u�?=�>=�<>=�~==ܿ<=��;=�>;=�|:=��9=H�8=�/8=�h7=��6=�5=�5=P?4=�p3=٠2=��1=��0=,$0=tK/=+p.=,�-=M�,=v�+=c�*=��)=)=p(= ''=�-&=�/%=�-$=G'#=�"=�!=��=�=i�=�=Tg=y4= �=0�=nt=�&=Y�=�v=Q=ߪ=�:=O�=]E=��	=�5=r�=�=�o=u�=�# =U��<��<��<��<b�<$��<���<�^�<��<�<%e�<^��<K��<H7�<�s�<L��<���<�<5@�<^k�<ޓ�<ֹ�<�ݫ<��<��<�<�<�X�<ps�<ߌ�<*��<~��<3ӈ<^�<5��<�)z<'Ur<!�j<��b<�Z<�S<�<K< pC<��;<�3<@,<}W$<>�<��<�(<w<l��;�G�;��;G��;Ϯ�;[��;ԗ�;���;'̂;Nh;��J;�}-;t�;dt�:�V�:�Zk:t�9D�:8K@Ź��O�@睺�MӺ���u�7�)Q��j�X���q���W���	������tλ�o�ƻ��ѻEbܻ�����[��*s��B����$��/�f�����"��G&�C\*��\.�TI2��#6���9���=�UKA�6�D�oH���K�*^O�7�R�/V�pY�j�\���_��+c�QYf�ni�_�l���o�Q�r��u�"�x���{���~�B瀼a���؃�'O���Æ�I7��s���\��b���B���Bg��GԐ�i@���������X���痼�O��˶��"��ꂝ�/螼 M������9���z���ޥ�\C��֧��o��2q��#֬�;��-���[���j��г��5��,���� ���f��ͺ��3��x����  �  ��N=�N=�XM=.�L=S�K=":K=��J=��I=tI=�aH=��G=��F=7<F=d�E=&�D=�D=�ZC=f�B=��A=%-A=/r@=��?=�>=�<>=�~==ֿ<=��;=�>;=�|:=��9=!�8=�/8=�h7=y�6=��5=�5=*?4=�p3=��2=��1=�0= $0=`K/=#p.=�-=S�,=v�+=l�*=�)=!)=�(=''=�-&=0%=.$=r'#="=�!=%�=7�=��=�=hg=�4='�=+�=ot=�&=K�=�v=;=Ȫ=N:=�=E=��	=�5=;�=�=ao=A�=�# =0��<���<��<��<?�<"��<���< _�<���<L�<Re�<���<���<�7�<Kt�<���<Z��<��<�@�<�k�<��<��<�ݫ<C��<��<�<�<�X�<^s�<ӌ�< ��<m��<�҈<�<���<�(z<�Tr<W�j<V�b</�Z<�
S<<K<�oC<�;<��3<
,<HW$</�<��<�(<Lw<��;�H�;��;���;O��;��;���;<��;΂;�h;��J;m�-;��;y�:�Y�:�`k:�	�9��:8�>Ź��O��睺KOӺ'�����7�"Q�Cj�5Y���r���X��;������ϻ���ƻμѻ�bܻ������s�vB����ƕ��������o"��F&��[*��[.�kH2��"6��9��=��JA���D��nH���K�+^O��R�aV�0pY���\��_��+c�Zf��i�7�l�A�o��r���u���x���{���~��瀼"a��"ك�DO���Æ�[7��f���^��D���(���g��Ԑ� @��<�������~���痼PO��`�����������瞼�L���������z���ޥ�WC������_q��6֬�N;���������k��eг��5��x���K��-g��Yͺ��3�������  �  ��N=�N=�XM=0�L=W�K=4:K=��J=��I=�I=bH=1�G=��F=u<F=��E=p�D=�D=�ZC=��B=��A=[-A=Zr@=��?=>�>=�<>=�~==ٿ<=��;=�>;=�|:=]�9=��8=X/8=oh7=@�6=��5=�5=�>4=�p3=v�2=d�1=H�0=�#0=?K/=p.=�-=V�,=z�+=��*=(�)=J)=�(=N''=�-&=I0%=G.$=�'#=T"=�!=e�=f�=��=2�=�g=�4=<�=)�=kt=�&=$�=�v==��=:=��=�D=L�	=85=�=�=o=�=P# =���<R��<:�<���<.�<��<���</_�<:��<��<�e�< ��<��<8�<�t�<*��<���<�<A�<.l�<���<}��<ޫ<���<�<�<�<�X�<Ls�<���<���<��<�҈<��<`��<�'z<fSr<0j<-�b<6�Z<�	S<;;K<�nC<��;<�3<o,<�V$<'�<��< )<�w<0��;.J�;q	�;{��;\��;1��;���;Ϋ�;%Ђ;.h;�J;Y�-;��;��:H`�:lk:��9��:8k7Ź0�O�^ꝺ)RӺ�-�C�7�7%Q�Vj�![���t���Z���������
ѻ���ƻ�ѻ�cܻ���#����s�B�������������]"��E&�Z*��Z.��G2��!6�J�9�7�=�JA�.�D�KnH�6�K�^O�
�R�aV��pY�.�\���_��,c��Zf��i�&�l�1�o�&�r���u���x���{�]�~��瀼�a��kك��O��)Ć�U7��c���L����������f���Ӑ��?��Ҫ����w~��痼�N��굚�M��$����瞼�L��F������Zz���ޥ�SC���������q���֬��;��䠯�*���k���г��6���������g���ͺ�+4��򚽼�  �  ��N=�N=�XM="�L=c�K=O:K=ʄJ=��I=�I=ZbH={�G=S�F=�<F=��E=��D=@D=S[C=�B=�A=�-A=�r@=ʶ?=R�>==>=�~==ʿ<=��;=�>;=p|:= �9=��8=/8=h7=�6=B�5=+5=�>4=9p3="�2=!�1=�0=�#0=K/=�o.=
�-=J�,=��+=��*=A�)=r)=�(=�''=2.&=�0%=�.$=(#=�"=L!=��=��=��=d�=�g=�4=I�=6�=Wt=�&=�=gv=�=9�=�9=u�=pD=ڿ	=�4=z�==�n=��=�" =��<؃�<��<^��<��<���<���<B_�<a��<��<)f�<���<���<�8�<cu�<���<���<��<�A�<�l�<,��<<jޫ<���<D�<�<�<�X�<5s�<j��<��<���<҈<�<���<�&z<�Qr<�}j<��b<��Z<^S<�9K<�mC<��;<\�3<�,<�V$<ۘ<��<c)<x<R��;�K�;��;���;.��;L��;Ϟ�;V��;;ӂ;�h;��J;�-;��;���:2f�:uk:,�9�?;867Ź7�O��읺�UӺ�U���7��)Q�j#j��]��jw���]��K�������һ�7�ƻ��ѻ�dܻ&��~����r��A����f����օ�����"��D&��X*�4Y.�*F2�T 6��9���=�#IA���D��mH���K��]O�-�R��V��pY���\���_��-c��[f�@�i�v�l���o���r�B�u�,�x���{���~�q耼b���ك��O��PĆ�p7��d�����ۉ������]f��#Ӑ�?��4���_���}��C旼N��6�����������枼 L���������%z���ޥ�nC��!�������q��׬�/<��w������7l���ѳ�27��Ɯ��l��Ih��Sκ��4��g����  �  F�N=�N=yXM=�L=m�K=_:K=��J=<�I=I=�bH=ѫG=��F=7=F=d�E=6�D=�D=�[C=G�B=`�A=�-A=�r@=�?=y�>=#=>=�~==��<=��;=q>;=5|:=�9=`�8=�.8=�g7=}�6=��5=�
5=%>4=�o3=Ɵ2=��1=��0=�#0=�J/=�o.=��-=J�,=��+=��*=s�)=�)=5(=�''=�.&=�0%=/$=p(#="=�!=�=��=I�=��=�g=�4=V�=<�=Mt=�&=��=!v=~=�=X9=�=D=a�	=R4=�=�=An=-�=�" =k��<@��<S�<��<��<��<��<n_�<���<W�<�f�<0��<L��<�9�<=v�<���<e��<��<�B�<m�<͕�<���<�ޫ<. �<r�<�<�<�X�<s�<"��<��<+��<�ш<X�<���<�$z<2Pr<|j<�b<�Z<�S<k8K<DlC<��;<Q�3<.,<.V$<��<�<�)<�x<c��;N�;>�;���;:��;ͤ�;v��;���;ׂ;� h;��J;z�-;W�;��:	p�:b�k:Q=�9��;8>5Ź�O�W�A[Ӻ����j�7��.Q�.)j��`��?z��P`����������ջ��ƻ�ѻfܻ������Or�:A����N�������K��~"��B&�`W*��W.�hD2��6���9���=�HA�t�D�mH�|�K�p]O� �R��V�iqY���\�h�_��.c�%]f���i��l�J�o�&�r���u���x�Y�{��~�逼�b��6ڃ�%P���Ć��7��W����������+����e���Ґ�t>����������|���嗼MM��b������䀝�`枼�K��w���K��z���ޥ�vC��M���>��Zr��y׬��<��(�������l��tҳ��7������7��i��Ϻ�B5��ԛ���  �  �N=cN=`XM=�L=v�K=x:K='�J=m�I=`I=�bH=8�G=�F=�=F=ׅE=��D=D=\C=��B=��A=1.A=s@=7�?=��>=6=>=�~==��<=��;=M>;=�{:=��9=�8=X.8=Vg7=�6=n�5=Q
5=�=4=lo3=i�2=s�1=o�0=C#0=�J/=�o.=�-=K�,=��+=��*=��)=�)=�(=;('=�.&=_1%=o/$=�(#=}"=!=v�=e�=��=�=h=5=t�=;�=Et=j&=��=�u=,=~�=�8=��=C=�	=�3=z�==�m=��=-" =���<���<��<���<�<Ҍ�<��<�_�<��<��<)g�<ڲ�<��<W:�<w�<���<O��<s�<]C�<Zn�<w��<#��<j߫<� �<��<=�<�X�<�r�<勔<���<���<�Ј<��<)��<#z<eNr<zj<�b<.�Z<S<�6K<�jC<G�;<Z�3<�,<�U$<��<&�<�)<�y<���;dP�;��;A��;׻�;h��;m��;���;ۂ;q(h;y�J;��-;?�;S��:wx�:��k:P�9�<8r0Źy�O���f`Ӻ��$���7��4Q�6/j��c���}��^c��$��3����׻���ƻ��ѻcgܻ���N���r��@����d����0������"�!A&��U*��U.��B2�66���9�R�=��FA���D�:lH���K�A]O��R� V��qY�7�\�i�_�0c�q^f��i���l���o���r���u�{�x��{�q�~��逼(c���ڃ�rP���Ć��7��J������>�������Re��Ґ��=���������|���䗼gL������������垼K���������y���ޥ�{C��y������r��ج�t=��Ϣ��M���m��Nӳ��8��f������i���Ϻ��5��g����  �  �N=4N=IXM=�L={�K=�:K=K�J=��I=�I=HcH=��G={�F=>F=F�E=�D=�D=�\C=�B=�A=�.A=Vs@=i�?=��>=I=>=�~==��<=b�;=>;=�{:=N�9=��8=�-8=�f7=��6=��5=�	5=I=4= o3=��2=�1="�0=#0=�J/=�o.=ב-=D�,=��+=��*=��)=$)=�(=�('=F/&=�1%=�/$=L)#=�"=�!=��=��=�=4�=Qh=$5=��=:�=2t=P&=o�=�u=�=�=�8=�=�B=]�	=F3=�=�
=@m=A�=�! =���<��<U�<>��<J�<���<��<�_�<T��<8�<�g�<u��<���<1;�<�w�<��<4��<R�<2D�<o�<,��<ɼ�<�߫<� �<��<$=�<�X�<�r�<���<K��<��<6Ј<��<I��<d!z<�Lr<Dxj<%�b<h�Z<IS<=5K<jiC<�;<v�3<�,<;U$<P�<+�<Q*<z<���;�R�;��;��;;��;%��;G��;���;�ނ;_0h;��J;��-;ܞ;c��:��:�k:c�9T[<8�,ŹD�O�����dӺh�B(���7�g:Q�"5j��f�������f��=��_���tڻ���ƻ��ѻ�hܻ��滔�����q�@�%��a��B�ځ�,��"�n?&��S*�
T.��@2�{6���9��=�{EA���D��kH�W�K�]O� �R�P V��rY���\�X�_�B1c��_f�Ɇi�K�l���o���r�_�u�%�x���{��~�fꀼ�c��ۃ��P��ņ��7��L����������j����d��Tѐ�=��꧓����4{���㗼�K������L��h��垼fJ����������y���ޥ��C���������!s���ج�>������&	���n��4Գ��9��L�������j��wк��6����  �  ��N=N=9XM=�L=��K=�:K=u�J=��I=�I=�cH=�G=��F=s>F=��E=�D=�D=�\C=o�B=l�A=�.A=�s@=��?=��>=_=>=�~==��<=P�;=�=;=�{:=	�9=n�8=�-8=�f7=<�6=��5=�	5=�<4=�n3=��2=��1=��0=�"0=MJ/=`o.=Ñ-=>�,=��+=	�*=��)=[)=(=�('=�/&=!2%=;0$=�)#=K"=�!=3�=�=2�=h�=h=P5=��=C�="t=1&=G�=_u=�=˨=#8=��=�B=ڽ	=�2=x�=
=�l=��=b! =,��<c��<��<���<�<���<��<`�<���<��<Gh�<��<���<�;�<�x�<H��<���<%�<�D�<�o�<ؗ�<B��<e�<R�<0 �<C=�<�X�<�r�<>��<Ѣ�<���<�ψ<1�<���<�z<�Jr<�vj<^�b<��Z<�S<�3K<,hC<֞;<V�3<�,<�T$<�<>�<�*<�z<���;�T�;S�;��;f¾;���;���;=��;l�;g7h;?�J;��-;v�;J��:o��:��k:sv�9��<8z*Ź�O�i���wkӺ��>,�s�7�A?Q�,;j��i��~����i�����򖰻�ܻ���ƻ��ѻMjܻ��������q��?�P��t��S�w������"��=&�.R*�rR.�]?2�6�"�9���=��DA���D��jH���K��\O�.�R�� V��rY�ѻ\�h�_�I2c�af�1�i���l�l�o�:�r���u���x��{�{�~�뀼Id���ۃ�<Q��.ņ��7��J��������������_d���А�b<��2���4��qz���◼�J��籚�����~��s䞼�I��+���G��ay��uޥ��C������.���s��٬��>��?����	��po��ճ��:��!������Qk��#Ѻ�7������  �  |�N=�N=XM=��L=��K=�:K=��J=�I=I=�cH=2�G=,�F=�>F=	�E=��D=ND=C]C=ģB=��A=/A=�s@=ķ?=�>=o=>= ==��<=6�;=�=;=`{:=շ9="�8=N-8=;f7=�6=9�5=	5=�<4=Fn3=S�2=w�1=��0=�"0=/J/=Ko.=��-=@�,=��+=�*=�)=�)=F(=)'=�/&=q2%=�0$=*#=�"=B!=��=\�=n�=��=�h=i5=��=H�=t=&=%�=5u=R=��=�7=P�=%B=s�	=[2=
�=�	=hl=z�=! =���<���<}�<���<��<���<(��<`�<��<��<�h�<���<$��<�<�<xy�<���<���<��<�E�<op�<[��<ý�<��<��<\ �<h=�<�X�<}r�<��<���<*��<ψ<��<���<Cz<IIr<�tj<�b<+�Z<] S<z2K<�fC<��;<��3<x,<eT$<�<o�<�*<#{<͠�;�V�;d�;���;?ž;���;��;Y��;��;�=h;]�J;ީ-;;�;��:g��:�k:+��9�=8�+ŹD�O������nӺx�`0�i�7�8DQ�@@j�l��_���Gl�����6���#߻���ƻ��ѻkܻ\�滹���>q�7?�������V�j�`��J"�B<&��P*��P.��=2��6���9���=��CA���D�4jH���K��\O��R�� V�JsY�F�\��_�53c�Qbf�_�i�#�l���o���r�l�u�:�x�|�{���~��뀼�d���ۃ�nQ��\ņ��7��1���g�����������c��PА��;����������y��>◼J��2������~���㞼~I��ڮ����=y��Vޥ��C������W���s��x٬�%?��٤��|
��+p���ճ�P;��Ѡ��e���k���Ѻ��7��᝽��  �  U�N=�N=XM=��L=��K=�:K=��J=%�I=SI=dH=d�G=g�F=?F=N�E=�D=�D=|]C=��B=��A=C/A=�s@=�?=#�>=x=>=�~==��<=!�;=�=;=6{:=��9=��8=-8=�e7=��6=��5=�5=L<4=n3=�2=B�1=i�0=h"0=J/=,o.=��-=>�,=��+=4�*=9�)=�)=(=K)'=!0&=�2%=�0$=H*#=�"=y!=��=��=��=ҕ=�h=�5=��=@�=t=�%=��=u==A�=�7=�=�A=0�	=2=��=c	=l=:�=�  =$��<���<$�<g��<��<���<$��<M`�<��<F�<i�<���<���<=�<�y�<���<H��<S�<F�<�p�<���<8��<�<��<� �<e=�<�X�<ar�<ي�<?��<Ѹ�<�Έ<)�<o��<3z<QHr<�sj<�b<�Z<\�R<�1K< fC<2�;<�3<�,<T$<ȗ<`�<&+<�{<��;TX�;�;a��;?Ǿ;���;m��;�Ñ;>�;�Ah;r�J;n�-;�;���:㕮:��k:Ď�9c1=8k)ŹG�O������rӺ!�c3�D�7��GQ�yCj�Wn��{����m����������໻�ƻ�ѻ/lܻ9������?q��>�=����e��~����T"�Y;&��O*��O.��<2��6���9���=��BA�>�D��iH�"�K��\O��R�!V��sY�׼\���_�4c�cf�-�i�2�l���o���r�u�u��x���{�p�~�쀼e��B܃��Q���ņ�8��9���\��O���u����c���ϐ�};�������+y���ᗼxI������r���}���㞼I���������y��]ޥ��C��������.t���٬��?��>����
���p��/ֳ��;��J������nl��#Һ�8��:����  �  D�N=�N=XM=��L=��K=�:K=��J=;�I=[I='dH=��G=��F=5?F=u�E=M�D=�D=�]C=*�B=�A=\/A= t@=��?=+�>=�=>=�~==��<=�;=�=;="{:=��9=��8=�,8=�e7=q�6=��5=�5=<4=�m3=�2=�1=N�0=N"0=�I/=o.=��-=6�,=��+=<�*=H�)=�)=�(=u)'=J0&=�2%=�0$=t*#="=�!=��=��=��=ܕ=�h=�5=��=G�=t=�%=��=�t= =�=`7=ٿ=�A=�	=�1=��=#	=�k=�=�  =���<R��<��<K��<��<j��<3��<S`�<<��<V�<Ai�<L��<���<i=�<Dz�<��<���<��<�F�</q�<��<K��<4�<��<� �<p=�<�X�<ar�<���<!��<���<tΈ<��<��<rz<oGr<'sj<�b<K�Z<��R<�0K<�eC<��;<��3<�,<T$<��<c�<I+<�{<���;�X�;'�;���;�Ⱦ;H��;Ǵ�;oő;��;NEh;��J;��-;�;���:h��:h�k:��9�;=8�'Źg�O�� ���tӺ�"��4���7�GJQ��Fj��o�������o��� ��%����ỻ��ƻ��ѻ�lܻ��������q��>����ʎ�8�~����z"��:&��N*�%O.�H<2��6�N�9�+�=�wBA���D�qiH��K�T\O�8�R�!V��sY��\��_�|4c��cf��i�תl���o���r�.�u���x�-�{�2�~�A쀼Se��m܃��Q���ņ�8��E���E��@���K���~c���ϐ�";��¥������x��Sᗼ'I��b�����]}��M㞼�H��m������y��Tޥ��C��������Lt��ڬ��?������I��q���ֳ�*<������F���l��wҺ�H8��w����  �  A�N=�N=XM=�L=��K=�:K=��J=X�I=lI=7dH=��G=��F=>?F=}�E=^�D=�D=�]C=)�B=�A=k/A=t@=�?=$�>=�=>= ==��<=�;=�=;={:=y�9=��8=�,8=�e7=h�6=��5=�5=<4=�m3=��2=�1=A�0=="0=�I/=o.=��-=6�,=��+=5�*=S�)=�)=�(=�)'=H0&=�2%=�0$=~*#="=�!=��=��=ϼ=�=�h=�5=��=S�=t=�%=��=�t=�=�=P7=ȿ=�A=ݼ	=�1=x�=	=�k=��=�  =���<>��<��<2��<��<s��<F��<@`�<c��<��<[i�<]��<���<~=�<Xz�<
��<���<��<�F�<.q�</��<i��<q�<��<� �<�=�<�X�<Pr�<���<��<t��<^Έ<��<���<gz<"Gr<sj<��b<:�Z<�R<�0K<meC<n�;<��3<|,<�S$<��<��<K+<�{<���;2Y�;��;���;�Ⱦ;���;��;Ƒ;��;Fh;��J;�-;�;���:u��:��k:ߛ�9�Y=8m*Ź��O����tuӺi#�T5���7�JQ�7Gj�6p��Ӊ��p��� ������⻻E�ƻ`�ѻ�lܻ���������p��>����J����}����q"��:&��N*��N.�(<2��6�V�9��=�CBA���D�:iH�'�K�\O�2�R�%!V�$tY�"�\�U�_��4c��cf�-�i�êl���o���r�\�u�(�x��{�r�~�X쀼me��܃��Q���ņ�8��;���1��S���#���Mc���ϐ�;��ƥ������x��2ᗼI��R�����^}��+㞼�H��0������y��<ޥ��C��%������Qt��)ڬ��?������\��q���ֳ�:<��ӡ��M���l���Һ�[8�������  �  D�N=�N=XM=��L=��K=�:K=��J=;�I=[I='dH=��G=��F=5?F=u�E=M�D=�D=�]C=*�B=�A=\/A= t@=��?=+�>=�=>=�~==��<=�;=�=;="{:=��9=��8=�,8=�e7=q�6=��5=�5=<4=�m3=�2=�1=N�0=N"0=�I/=o.=��-=6�,=��+=<�*=H�)=�)=�(=u)'=J0&=�2%=�0$=t*#="=�!=��=��=��=ܕ=�h=�5=��=H�=t=�%=��=�t== �=b7=ڿ=�A=�	=�1=��=%	=�k=�=�  =���<X��<�<P��<��<o��<8��<X`�<@��<Z�<Di�<O��<���<j=�<Ez�<��<���<��<�F�<-q�<��<H��<1�<��<� �<l=�<�X�<]r�<���<��<���<qΈ<��<��<oz<nGr<'sj<�b<M�Z<��R<�0K<�eC<��;<��3<�,<T$<��<k�<Q+<�{<���;�X�;2�;���;�Ⱦ;L��;ȴ�;nő;��;@Eh;��J;�-;��;s��:��:��k:���9�0=8)Ź!�O�T��)uӺ�"��4��7�pJQ��Fj��o�������o��� ��2����ỻ��ƻ��ѻ�lܻ��������q��>����̎�9�~����{"��:&��N*�%O.�H<2��6�O�9�+�=�wBA���D�riH��K�T\O�8�R�!V��sY��\��_�|4c��cf��i�תl���o���r�.�u���x�-�{�2�~�A쀼Se��m܃��Q���ņ�8��E���E��@���K���~c���ϐ�";��¥������x��Sᗼ'I��b�����]}��M㞼�H��m������y��Tޥ��C��������Lt��ڬ��?������I��q���ֳ�*<������F���l��wҺ�H8��w����  �  U�N=�N=XM=��L=��K=�:K=��J=%�I=SI=dH=d�G=g�F=?F=N�E=�D=�D=|]C=��B=��A=C/A=�s@=�?=#�>=x=>=�~==��<=!�;=�=;=6{:=��9=��8=-8=�e7=��6=��5=�5=L<4=n3=�2=B�1=i�0=h"0=J/=,o.=��-=>�,=��+=4�*=9�)=�)=�(=K)'=!0&=�2%=�0$=H*#=�"=y!=��=��=��=ӕ=�h=�5=��=@�=t= &= �=u= =C�=�7=�=�A=3�	=2=��=g	=l=?�=�  =.��<���</�<r��<��<���<.��<U`�<!��<M�<!i�<���<���<=�<�y�<���<H��<Q�<F�<�p�<���<2��<�<��< �<^=�<�X�<Zr�<Ҋ�<8��<˸�<�Έ<$�<l��<.z<NHr<�sj<�b<!�Z<b�R<�1K<fC<>�;<�3<�,<'T$<ؗ<p�<6+<�{<���;lX�;�;r��;KǾ;���;p��;�Ñ;7�;�Ah;N�J;@�-;ެ;'��:V��:��k:7��9=8-,Ź��O�V ���sӺg!��3���7�HQ��Cj�{n�������m�����К���໻/�ƻ-�ѻ?lܻG������Cq��>�@����g��~����U"�[;&��O*��O.��<2��6���9���=��BA�>�D��iH�"�K��\O��R�!V��sY�׼\���_�4c�cf�-�i�2�l���o���r�u�u��x���{�p�~�쀼e��B܃��Q���ņ�8��9���\��O���u����c���ϐ�};�������+y���ᗼxI������r���}���㞼I���������y��]ޥ��C��������.t���٬��?��>����
���p��/ֳ��;��J������nl��#Һ�8��:����  �  |�N=�N=XM=��L=��K=�:K=��J=�I=I=�cH=2�G=,�F=�>F=	�E=��D=ND=C]C=ģB=��A=/A=�s@=ķ?=�>=o=>= ==��<=6�;=�=;=`{:=շ9="�8=N-8=;f7=�6=9�5=	5=�<4=Fn3=S�2=w�1=��0=�"0=/J/=Ko.=��-=@�,=��+=�*=�)=�)=F(=)'=�/&=q2%=�0$=*#=�"=B!=��=]�=o�=��=�h=j5=��=I�=t=&='�=7u=U=��=�7=T�=)B=w�	=`2=�=�	=nl=��=! =���<��<��<���<��<���<6��<&`�<��<��<�h�<���<*��<�<�<{y�<���<���<��<�E�<ip�<T��<���<��<��<Q �<]=�<�X�<rr�<��<���<!��<ψ<��<���<<z<FIr<�tj<�b<2�Z<g S<�2K<�fC<	�;<��3<�,<{T$<��<��<�*<8{<��;�V�;��;���;Qž;���;��;V��;��;b=h;*�J;��-;�;e��:���:g�k:���9��<8�/ŹA�O������oӺ���0���7��DQ��@j��l������ql�����Y���C߻���ƻ�ѻ,kܻp������Eq�=?�������Z�m�b��L"�C<&��P*� Q.��=2��6���9���=��CA���D�5jH���K��\O��R�� V�JsY�F�\��_�53c�Qbf�_�i�#�l���o���r�l�u�:�x�|�{���~��뀼�d���ۃ�nQ��\ņ��7��1���g�����������c��PА��;����������y��>◼J��2������~���㞼~I��ڮ����=y��Vޥ��C������W���s��x٬�%?��٤��|
��+p���ճ�P;��Ѡ��e���k���Ѻ��7��᝽��  �  ��N=N=9XM=�L=��K=�:K=u�J=��I=�I=�cH=�G=��F=s>F=��E=�D=�D=�\C=o�B=l�A=�.A=�s@=��?=��>=_=>=�~==��<=P�;=�=;=�{:=	�9=n�8=�-8=�f7=<�6=��5=�	5=�<4=�n3=��2=��1=��0=�"0=MJ/=`o.=Ñ-=>�,=��+=	�*=��)=[)=(=�('=�/&=!2%=<0$=�)#=L"=�!=3�=�=3�=h�=�h=Q5=��=E�=$t=3&=I�=bu=�=Ϩ='8=��=�B=�	=�2=�=
=�l=��=k! =>��<t��<��<��<!�<���<.��<`�<���<��<Sh�<'��<���<�;�<�x�<I��<���<"�<�D�<�o�<ϗ�<8��<Z�<E�<# �<5=�<�X�<�r�<2��<Ţ�<}��<�ψ<*�<���<�z<�Jr<�vj<b�b<��Z<�S<�3K<?hC<�;<n�3<�,<U$<4�<Y�<�*<�z<ǟ�;�T�;v�;2��;{¾;���;���;9��;^�;:7h;�J;3�-;�;p��:|��:��k:
r�9��<8B/Ź��O������lӺ���,��7��?Q��;j�+j������j�������ݻ���ƻ��ѻhjܻ��������q��?�V��y��W�z������"��=&�0R*�sR.�^?2�6�#�9���=��DA���D��jH���K��\O�.�R�� V��rY�һ\�h�_�I2c�af�1�i���l�l�o�:�r���u���x��{�{�~�뀼Id���ۃ�<Q��.ņ��7��J��������������_d���А�b<��2���4��qz���◼�J��籚�����~��s䞼�I��+���G��ay��uޥ��C������.���s��٬��>��?����	��po��ճ��:��!������Qk��#Ѻ�7������  �  �N=4N=IXM=�L={�K=�:K=K�J=��I=�I=HcH=��G={�F=>F=F�E=�D=�D=�\C=�B=�A=�.A=Vs@=i�?=��>=I=>=�~==��<=b�;=>;=�{:=N�9=��8=�-8=�f7=��6=��5=�	5=I=4= o3=��2=�1="�0=#0=�J/=�o.=ב-=D�,=��+=��*=��)=$)=�(=�('=F/&=�1%=�/$=L)#=�"=�!=��=��=�=5�=Rh=%5=��=<�=4t=R&=r�=�u=�="�=�8=�=C=c�	=M3=��=�
=Hm=J�=�! =���<��<i�<R��<^�<Č�<��<�_�<c��<F�<�g�<��<���<7;�<�w�<���<2��<O�<,D�<o�<"��<���<�߫<� �<��<=�<�X�<�r�<��<>��<��<+Ј<��<B��<[!z<|Lr<Dxj<*�b<q�Z<WS<N5K<iC<.�;<��3<�,<YU$<n�<I�<o*<-z<��; S�;��;?��;S��;4��;L��;���;�ނ;-0h;=�J;��-;s�;p��:��:˝k:'^�92<8�1Ź��O�`���HfӺ��(�V�7� ;Q��5j�Ag��򀍻�f��s�������ڻ���ƻ��ѻ�hܻ�滬�����q�@�,��g��G�݁�/��"�p?&��S*�T.� A2�|6���9��=�|EA���D��kH�W�K�]O� �R�P V��rY���\�X�_�B1c��_f�Ɇi�K�l���o���r�_�u�%�x���{��~�fꀼ�c��ۃ��P��ņ��7��L����������j����d��Tѐ�=��꧓����4{���㗼�K������L��h��垼fJ����������y���ޥ��C���������!s���ج�>������&	���n��4Գ��9��L�������j��wк��6����  �  �N=cN=`XM=�L=v�K=x:K='�J=m�I=`I=�bH=8�G=�F=�=F=ׅE=��D=D=\C=��B=��A=1.A=s@=7�?=��>=6=>=�~==��<=��;=M>;=�{:=��9=�8=X.8=Vg7=�6=n�5=Q
5=�=4=lo3=i�2=s�1=o�0=C#0=�J/=�o.=�-=K�,=��+=��*=��)=�)=�(=;('=�.&=_1%=o/$=�(#=}"=!=w�=f�=��=�=h=5=v�=<�=Gt=m&=��=�u=0=��=�8=��=�C=�	=�3=��==�m=��=6" =���<���<��<���<��<��<��<�_�<��<��<6g�<��<&��<]:�<#w�<���<M��<o�<WC�<Rn�<m��<��<]߫<� �<��<�<�<�X�<�r�<׋�<���<���<�Ј<��<"��<#z<`Nr<zj<�b<7�Z<)S<7K<�jC<`�;<u�3<�,<�U$<��<E�<*<�y<,��;�P�;��;b��;�;x��;r��;���;ۂ;=(h;0�J;?�-;ї;W��:_w�:�k:�J�9
�;8�5ŹI�O�?����aӺ^��$���7�05Q��/j�d���}���c��\��e���ػ���ƻ�ѻ�gܻ���f����r��@����j����4������"�#A&��U*��U.��B2�76���9�S�=��FA���D�:lH���K�B]O��R� V��qY�7�\�i�_�0c�q^f��i���l���o���r���u�{�x��{�q�~��逼(c���ڃ�rP���Ć��7��J������>�������Re��Ґ��=���������|���䗼gL������������垼K���������y���ޥ�{C��y������r��ج�t=��Ϣ��M���m��Nӳ��8��f������i���Ϻ��5��g����  �  F�N=�N=yXM=�L=m�K=_:K=��J=<�I=I=�bH=ѫG=��F=7=F=d�E=6�D=�D=�[C=G�B=`�A=�-A=�r@=�?=y�>=#=>=�~==��<=��;=q>;=5|:=�9=`�8=�.8=�g7=}�6=��5=�
5=%>4=�o3=Ɵ2=��1=��0=�#0=�J/=�o.=��-=J�,=��+=��*=s�)=�)=5(=�''=�.&=�0%=/$=p(#="=�!=�=��=I�=��=�g=�4=X�==�=Ot=�&=��=$v=�=�=]9=�=D=g�	=Y4=	�=�=In=6�=�" =~��<S��<g�<��<��<���<��<_�<Ͻ�<e�<�f�<:��<T��<�9�<@v�<���<d��<��<|B�<wm�<Õ�<{��<�ޫ<  �<d�<�<�<�X�<s�<��< ��< ��<yш<P�<���<�$z<-Pr<|j<�b<�Z<�S<}8K<YlC<��;<l�3<K,<LV$<˘<2�<�)<�x<���;NN�;f�;���;R��;ܤ�;{��;���;�ւ;� h;V�J;"�-;�;��:�n�:�k:f8�9nz;8�:Ź��O��񝺝\ӺQ�N �
�7�k/Q��)j��`��~z���`��#�������ջ�D�ƻ2�ѻ>fܻ�����Xr�BA����S�������N���"��B&�bW*��W.�iD2��6���9���=�HA�u�D�mH�|�K�p]O� �R��V�iqY���\�h�_��.c�%]f���i��l�J�o�&�r���u���x�Y�{��~�逼�b��6ڃ�%P���Ć��7��W����������+����e���Ґ�t>����������|���嗼MM��b������䀝�`枼�K��w���K��z���ޥ�vC��M���>��Zr��y׬��<��(�������l��tҳ��7������7��i��Ϻ�B5��ԛ���  �  ��N=�N=�XM="�L=c�K=O:K=ʄJ=��I=�I=ZbH={�G=S�F=�<F=��E=��D=@D=S[C=�B=�A=�-A=�r@=ʶ?=R�>==>=�~==ʿ<=��;=�>;=p|:= �9=��8=/8=h7=�6=B�5=+5=�>4=9p3="�2=!�1=�0=�#0=K/=�o.=
�-=J�,=��+=��*=A�)=r)=�(=�''=2.&=�0%=�.$=(#=�"=L!=��=��=��=e�=�g=�4=J�=8�=Yt=�&=�=iv=�=<�=�9=z�=uD=�	=�4=��==�n=��=# =��<��<��<p��<	�<��<��<Q_�<p��<��<5f�<���<���<�8�<fu�<���<���<��<�A�<�l�<$��<㺯<^ޫ<���<7�<�<�<�X�<(s�<]��<s��<���<҈<�<���<&z<�Qr<�}j<��b<��Z<jS< :K<�mC<��;<t�3<,<�V$<��<�<~)<1x<���;�K�; �;��;C��;Z��;Ӟ�;R��;.ӂ;�h;��J;̉-;��;��:?e�:sk:�'�9�;8�;Ź��O��흺�VӺ�����7�H*Q��#j�^���w���]��{�����ӻ�Z�ƻ��ѻ�dܻ>�滓�,���r��A����k����څ�����"��D&��X*�5Y.�+F2�U 6��9���=�#IA���D��mH���K��]O�-�R��V��pY���\���_��-c��[f�@�i�v�l���o���r�B�u�,�x���{���~�q耼b���ك��O��PĆ�p7��d�����ۉ������]f��#Ӑ�?��4���_���}��C旼N��6�����������枼 L���������%z���ޥ�nC��!�������q��׬�/<��w������7l���ѳ�27��Ɯ��l��Ih��Sκ��4��g����  �  ��N=�N=�XM=0�L=W�K=4:K=��J=��I=�I=bH=1�G=��F=u<F=��E=p�D=�D=�ZC=��B=��A=[-A=Zr@=��?=>�>=�<>=�~==ٿ<=��;=�>;=�|:=]�9=��8=X/8=oh7=@�6=��5=�5=�>4=�p3=v�2=d�1=H�0=�#0=?K/=p.=�-=V�,=z�+=��*=(�)=J)=�(=N''=�-&=I0%=G.$=�'#=U"=�!=f�=f�=��=2�=�g=�4==�=*�=lt=�&=&�=�v==��=:=��=�D=Q�	==5=�=�=o=�=W# =���<a��<H�<���<=�<��<���<;_�<E��<��<�e�<��<��<8�<�t�<+��<���<�<A�<(l�<���<t��<ޫ<���<��<�<�<�X�<Bs�<���<���<���<�҈<��<[��<�'z<cSr<0j<0�b<=�Z<�	S<H;K<�nC<��;<�3<�,<W$<>�<��<)<�w<V��;PJ�;�	�;���;n��;<��;ě�;ʫ�;Ђ;	h;�J;�-;O�;L�:�_�:Tjk:-�9��:8Q;Ź-�O�^띺(SӺ������7��%Q��j�S[��
u���Z��
������*ѻ���ƻ1�ѻ�cܻ���4����s�B� �����������_"��E&��Z*��Z.��G2��!6�K�9�7�=�JA�/�D�LnH�6�K�^O�
�R�aV��pY�.�\���_��,c��Zf��i�&�l�1�o�&�r���u���x���{�]�~��瀼�a��kك��O��)Ć�U7��c���L����������f���Ӑ��?��Ҫ����w~��痼�N��굚�M��$����瞼�L��F������Zz���ޥ�SC���������q���֬��;��䠯�*���k���г��6���������g���ͺ�+4��򚽼�  �  ��N=�N=�XM=.�L=S�K=":K=��J=��I=tI=�aH=��G=��F=7<F=d�E=&�D=�D=�ZC=f�B=��A=%-A=/r@=��?=�>=�<>=�~==ֿ<=��;=�>;=�|:=��9=!�8=�/8=�h7=y�6=��5=�5=*?4=�p3=��2=��1=�0= $0=`K/=#p.=�-=S�,=v�+=l�*=�)=!)=�(=''=�-&=0%=.$=r'#="=�!=%�=7�=��=�=hg=�4=(�=,�=pt=�&=M�=�v===ʪ=Q:=�=!E=��	=�5=?�=�=eo=F�=�# =:��<���<��<���<I�<,��<���<	_�<��<S�<Xe�<���<���<�7�<Mt�<���<Z��<��<�@�<�k�<��<��<�ݫ<<��<��<�<�<�X�<Ws�<̌�<���<g��<�҈<�<���<�(z<�Tr<W�j<Y�b<3�Z<�
S<"<K<�oC<��;<��3<,<XW$<?�<��<�(<[w<��;�H�;��;���;\��;��;���;9��;΂;jh;ٯJ;?�-;L�;�x�:;Y�:�_k:l�9��:8�AŹC�O��蝺�OӺ��2��7�S"Q��j�XY��s��Y��W��&����ϻ��ƻ�ѻ�bܻ���,� ��#s�yB����ɕ���������p"��F&��[*��[.�lH2��"6��9��=��JA���D��nH���K�+^O��R�aV�0pY���\��_��+c�Zf��i�7�l�A�o��r���u���x���{���~��瀼"a��"ك�DO���Æ�[7��f���^��D���(���g��Ԑ� @��<�������~���痼PO��`�����������瞼�L���������z���ޥ�WC������_q��6֬�N;���������k��eг��5��x���K��-g��Yͺ��3�������  �  ��N=�N=�XM=/�L=P�K=:K=��J=��I=VI=�aH=ЪG=��F=<F=0�E=�D=yD=�ZC=6�B=c�A=-A=r@=u�?=�>=�<>=�~==ܿ<=��;=�>;=�|:=��9=H�8=�/8=�h7=��6=�5=�5=P?4=�p3=٠2=��1=��0=,$0=tK/=+p.=,�-=M�,=v�+=c�*=��)=)=p(= ''=�-&=�/%=�-$=G'#=�"=�!=��=�=i�=�=Tg=y4= �=1�=nt=�&=Z�=�v=Q=�=�:=Q�=^E=��	=�5=t�=�=�o=w�=�# =Z��<��<��<��<g�<)��<���<�^�<��<#�<)e�<a��<M��<J7�<�s�<L��<���<�<3@�<\k�<ܓ�<ӹ�<�ݫ<��<��<�<�<�X�<ls�<܌�<'��<{��<0ӈ<[�<3��<�)z<&Ur<!�j<��b<�Z<�S<�<K<&pC<��;<�3<H,<�W$<F�<��<�(<w<z��;�G�;��;P��;ծ�;_��;֗�;���;#̂;Ah;��J;k}-;X�;#t�:�V�:;Zk:"�92x:8�AŹw�O��睺NӺA����7�RQ��j� X���q���W���	��ˆ���λ�z�ƻ��ѻMbܻ�����a��,s��B����&��1�g�����"��G&�C\*��\.�TI2��#6���9���=�UKA�6�D�oH���K�*^O�7�R�/V�pY�j�\���_��+c�QYf�ni�_�l���o�Q�r��u�"�x���{���~�B瀼a���؃�'O���Æ�I7��s���\��b���B���Bg��GԐ�i@���������X���痼�O��˶��"��ꂝ�/螼 M������9���z���ޥ�\C��֧��o��2q��#֬�;��-���[���j��г��5��,���� ���f��ͺ��3��x����  �  Z�N=vN=bQM=�L=(�K=0K=�yJ=��I=�I=TH=/�G=��F=c+F=arE=��D=:�C=
EC=K�B=�A=0A=�V@=u�?=p�>=�>=�\==0�<=p�;=�;=�S:=��9=p�8=� 8=�77=�m6=�5=��4=�4=�43=1b2=��1=�0=��/=x/=i$.=�C-='`,=�y+=Ï*=��)=�(=��'=��&=U�%=�$=c�#=6�"=O�!={� =��=Ke=�B==��=9�=�|=y;=��=¥=�P=p�=;�=T*=к=�D=,�
=7E	=�=�,=��=��=.\=�l�<G�<��<	L�<���<�\�<���<_L�<u��<��<�{�<I��<�&�<�s�<��<r��<�>�<1z�<��<��<�<�F�<�r�<���<"ħ<��<I�<I/�<�O�<�n�<��<5��<�ƈ<y�<���<�2z<�ir<��j<��b<5[<�LS<x�K<1�C<	<<�L4<,�,<E�$<�*<>|<`�<-<�;���;��;<��;1��;"��;_��;��;!�;Y�l;ƾO;+�2;��;���:j�:�ρ::��9x��,|4��⏺��ĺ'Y��&��R0��OI��'b���z�F\��J7��qߠ�
U��Ö��̤»�~ͻ%ػ,�⻠�� ���M^ �Q2���	�R��)�֑�H��k8 ��k$�P�(��,�ތ0�,r4�}F8��	<�ٽ?��bC���F���J�� N��rQ���T��5X���[���^�Fb�]Ie��yh�u�k�h�n�x�q���t��x�b{�$~���������������:u���뇼�a���Պ��H������a+������	���w��Q䔼TP��b����%���������,`���Ǟ�,/���������Nc���ɥ�>0������C����c��`ʬ�1��엯������e���̳�4��l�������j���Һ��:�������  �  L�N=~N=bQM=�L=-�K=0K=�yJ=��I=�I=%TH=>�G=�F=c+F=qrE=�D=J�C=	EC=T�B=�A=:A=�V@=z�?=r�>=�>=�\==.�<=t�;=�;=�S:=��9=c�8=� 8=�77=�m6=ء5=��4=�4=�43=-b2=��1=ֶ0=��/=j/=r$.=�C-=)`,=�y+=ď*=��)=��(=��'=��&=b�%=�$=k�#=B�"=Z�!=�� =��=Ve=�B==��=?�=�|=u;=��=��=�P=b�=$�=I*=ĺ=�D=�
=.E	=�=�,=��=��=&\=sl�<+�<׵�<�K�<���<�\�<���<KL�<t��<��<|�<]��<�&�<�s�<���<���<�>�<Pz�<��<��<%�<�F�<�r�<���<(ħ<��<R�<N/�<�O�<�n�<��<��<�ƈ<j�<���<�2z<lir<��j<��b<[<�LS<U�K<��C<�<<�L4<H�,<?�$<�*<M|<O�<-<��;���;O��;���;\��;)��;踢;�;�!�;a�l;t�O;�2;_�;#��:\�:OЁ:X:$�99��`z4��ᏺ��ĺ8Z��Ώ��0�>PI�(b�D�z��\��r7���ߠ�!U������»�ͻz%ػ֗⻺�����I^ �H2���	� ���������r8 ��k$��(��,���0�3r4�NF8��	<���?��bC���F���J�� N��rQ��T�^5X�Ӈ[�!�^�kb��Ie��yh���k���n���q���t��x��{�:~�������ւ������-u��쇼�a���Պ��H��~���D+�������	��{w��T䔼6P��E���}%��
�������`���Ǟ�/���������Sc���ɥ�;0������.����c��~ʬ�'1�����������e���̳�/4��}�������j���Һ��:�������  �  >�N=sN=PQM=�L=5�K=0K=�yJ=��I=�I=5TH=Z�G="�F=�+F=�rE=)�D=o�C=(EC=u�B=(�A=JA=�V@=��?=��>=�>=�\==$�<=e�;=�;=�S:=��9=H�8=� 8=�77=m6=��5=^�4=j4=�43=b2=u�1=Ƕ0=��/=]/=i$.=�C-=.`,=�y+=Ώ*=��)=	�(=��'=��&=��%=1�$=��#=`�"=u�!=�� =��=we=�B=*=��=E�=�|=u;=��=��=�P=O�=�=9*=��=�D=��
=
E	=ۻ=�,=t�=��=\=.l�<�<���<�K�<���<�\�<���<NL�<���<��<)|�<y��<�&�<"t�<7��<���<?�<�z�<`��<��<f�<G�<#s�<ɜ�<Nħ<��<c�<N/�<�O�<�n�<錐<��<eƈ<.�<���<2z<�hr<�j<M�b<�[<HLS<ՈK<��C<�<<EL4<�,<��$<�*<i|<n�<Y-<��;!��;ѿ�;���;n��;O��;��;�;�"�;��l;��O;��2;��;���:o�:�Ӂ:�:��9����|4��⏺K�ĺBZ��.��0�5RI��)b��z��]��58���࠻�U��՗��u�»�ͻ�%ػ��4������2^ �2���	�����n������7 ��j$���(�r�,��0��q4��E8��	<�]�?��bC���F�[�J�� N�wrQ�M�T��5X��[�8�^��b��Ie�0zh�8�k���n�G�q�B�t�\x�#{��~�Q�����肃�����Eu��쇼xa���Պ��H��k���(+��Ԛ���	��9w��䔼�O�����:%��Î�������_���Ǟ��.��액�����@c���ɥ�?0��ʖ��C����c���ʬ�S1��7������'f��2ͳ�w4������C���j���Һ�.;��ɣ���  �  (�N=]N=OQM=�L=3�K='0K=�yJ=��I=�I=bTH=��G=L�F=�+F=�rE=c�D=��C=\EC=��B=R�A=wA=�V@=��?=��>=�>=�\==$�<=_�;=�;=�S:=u�9= �8=� 8=�77=Om6=��5=0�4=44=z43=�a2=L�1=��0=��/=G/=V$.=�C-=-`,=�y+=ݏ*=Ƣ)=)�(=�'=��&=��%=_�$=��#=��"=��!=֚ =�=�e=�B=N=��=Z�=�|=r;=��=��=�P=2�=�=�)=n�=YD=��
=�D	=��=a,=8�=J�=�[=�k�<��<n��<�K�<���<�\�<}��<ML�<���<��<d|�<���<A'�<pt�<���<4 �<�?�<�z�<Ų�<F�<��<eG�<ps�<��<~ħ<��<f�<R/�<�O�<�n�<���<ũ�<ƈ<��<X��<N1z<hr<T�j<j�b<�[<�KS<+�K<��C<�<<�K4<��,<��$<�*<U|<��<�-<��;E��;L��;��;��;��;ǻ�;	�;�$�;k�l;��O;�2; ;d��::�:�ց:�:��9��|4��䏺n�ĺ_��1���0�kTI�g,b�ޥz�_���9���ᠻW������Ѧ»�ͻ_&ػ���������$^ ��1��	�c����������27 �?j$���(���,�Y�0��p4�E8��<���?��aC�#�F� �J�� N�|rQ�N�T��5X�[�[���^�Ub��Je��zh��k���n��q��t�!x��{�C~�����a��������Xu��쇼�a���Պ�rH��5����*��~���8	���v���㔼�O�������$��a���=����_��AǞ��.������{���(c���ɥ�@0��ʖ��m���d���ʬ��1������u����f���ͳ��4��&������Lk��7Ӻ��;������  �  �N=CN=AQM=�L=;�K=;0K=�yJ=$�I=I=�TH=��G=��F=�+F=sE=��D=��C=�EC=ߊB=��A=�A=
W@=ř?=��>=�>=�\==�<=N�;=l;=vS:=I�9=��8=R 8=^77=m6=@�5=��4=�4=<43=�a2=�1=n�0=�/=*/=@$.=�C-=%`,=�y+=��*=�)=M�(=	�'=��&=��%=��$=��#=ӻ"=�!=� ='�=�e= C=n=��=r�=�|={;=��=��=�P=�==�)=7�=D=p�
=zD	=S�=,=�=��=�[=Zk�<)�<��<IK�<T��<�\�<n��<`L�<���<�<�|�<��<�'�<�t�<(��<� �<@�<z{�<O��<��<2�<�G�<�s�<b��<�ħ<�<��<G/�<�O�<�n�<���<q��<�ň<t�<���<M0z<�fr<I�j<E�b<�[<jJS<4�K<�C<8<<RK4<,�,<��$<m*<k|<��<�-<�;d��;���;��;$��;a��;���;��;�&�;c�l;��O;r�2;z;g��:G"�:cځ:�:D9!���}4��揺��ĺPc��0��V#0��WI�0b���z��`���;���㠻Y��D�����»��ͻ%'ػ��U�������] �x1���	�Ə�i�؏����6 �4i$���(�}�,�V�0��o4�/D8��<�"�?�daC���F�΂J�{ N��rQ�v�T�6X�̈[�C�^��b�IKe��{h�ߤk���n��q��t�1x��{�G~�􉀼���`���J���~u��0쇼{a��rՊ�PH����*��.������kv�� 㔼O�����W$��ڍ������_���ƞ�W.��a���N��� c���ɥ�Q0��疨�����Kd��(ˬ��1��혯������f��&γ�M5���������k���Ӻ��;��t����  �  ߺN=(N=.QM=�L=B�K=G0K=�yJ=K�I=7I=�TH=��G=��F=G,F=SsE=��D=- D=�EC= �B=��A=�A=?W@=�?=��>=�>=�\==�<=:�;=O;=JS:=�9=��8= 8=77=�l6=�5=��4=�4=�33=ca2=ی1=5�0=T�/=/=+$.=�C-=)`,=�y+= �*=��)=|�(=C�'=7�&=#�%=��$=I�#=�"=4�!=`� =c�=f=:C=�=&�=��=�|=|;=��=u�=�P=��=��=�)=�=�C=�
=D	=�=�+=��=��=2[=�j�<��<���<�J�<��<c\�<b��<ZL�<Ը�<E�<�|�<q��<$(�<`u�<���<Q�<�@�<|�<볾<]�<��<KH�<4t�<���<�ħ</�<��<P/�<�O�<hn�<4��<��<@ň<���<G��</z<�er<�j<��b<g[<MIS<�K< �C<x<<�J4<��,<3�$<V*<||<��<o.<[�;'��;���;$��;a��;�;���; �;�)�;��l;~�O;8�2;�;���:�(�:�߁:S#:�!9���.4��菺��ĺ�g������&0�l[I�*4b��z�c���=���堻�Z��)�����»��ͻ4(ػ��⻭�컬����] �*1��	����s�َ����5 ��g$���(�H�,��0��n4�$C8��<�5�?��`C��F�}�J�T N�xrQ���T�g6X�]�[���^��b�XLe��|h���k��n�G�q�J�t�Zx��{�K~�x��������������u��E쇼oa��cՊ�H������0*������D���u���┼mN��{����#��B���0����^��hƞ��-���������b���ɥ�N0����������d��{ˬ�u2��r���} ���g���γ��5��H������Ql��-Ժ�Q<��Ǥ���  �  ��N=N=QM=ޛL=J�K=\0K=zJ=k�I=oI=UH=G�G=�F=�,F=�sE=J�D=� D=4FC=m�B=�A=A=rW@=�?=��>=�>=�\==�<=%�;=1;=S:=�9=s�8=��7=�67=nl6=��5=H�4=S4=�33=a2=��1=��0=#�/=�/=$.=�C-=(`,=�y+=�*="�)=��(=w�'=o�&=m�%=-�$=��#=s�"=��!=�� =��=Wf=pC=�=J�=��=�|={;=��=Z�=^P=��=L�==)=��=cC=��
=�C	=��=Q+=(�=F�=�Z=j�<�<��<�J�<���<9\�<P��<\L�<��<p�<N}�<���<�(�<�u�<;��<��<SA�<�|�<���<��<Z�<�H�<�t�<	��<Hŧ<g�<��<P/�<_O�<>n�<܋�<���<�Ĉ<c��<���<�-z<adr<u�j<��b<�[<�GS<�K<��C<�<<�I4<8�,<��$<7*<�|<K�<�.<g�;���;���;���;���;���;�â;#�;�,�;��l;�O;d�2;W;���:-.�:��:�*:�49M���4��ꏺ��ĺ�l����^*0��_I��8b�q�z��e��@��N蠻�\�����C�»!�ͻI)ػ?��$�컈���v] ��0�|�	�Q����������3 ��f$��(��,�Ǉ0��m4��A8��<�^�?��_C���F��J�/ N�qrQ���T��6X��[���^��b�`Me�	~h�S�k�M�n���q���t��x�#{�^~����������������u��U쇼ia��JՊ��G��j����)��L������Nu��┼�M��и��#�����������]���Ş�z-��ʔ�������b���ɥ�T0��2��������d���ˬ��2��������=h��\ϳ��6��坶�\���l���Ժ��<��/����  �  ��N=�N=QM=֛L=O�K=q0K=3zJ=��I=�I=EUH=��G=m�F=�,F=�sE=��D=� D=�FC=��B=T�A=PA=�W@=4�?=��>=�>=�\==�<=�;=;=�R:=��9=:�8=��7=~67=l6=L�5=��4=4=T33=�`2=X�1=µ0=��/=�/=�#.=yC-=%`,=�y+=/�*=A�)=в(=��'=��&=��%=��$=��#=��"=ٮ!=�� =��=�f=�C==q�=��=�|=�;=��=E�=5P=|�=�=�(=H�=C=\�
=\C	=&�=�*=Ǖ=��=�Z={i�<��<���<.J�<z��<\�<:��<nL�< ��<��<�}�<C��<)�<�v�<��<��<B�<j}�<7��<��<��<OI�<u�<t��<�ŧ<��<��<I/�<CO�<�m�<���<N��<LĈ<�߄<
��<m,z<�br<�j<8�b<�[<�FS<��K<��C<�<<"I4<��,<l�$<*<�|<��<[/<� �;���;���;İ�;���;��;~Ƣ;*�;�/�;m;��O;Z�2;�;��:t5�:��:+3:E9�
��(�4��폺Z�ĺKr����f.0�dI�1=b�S�z�h��mB��W꠻$_������լ»q�ͻ*ػ��_�����@] �L0���	������Ќ����q2 �Ze$�Ƀ(���,�z�0�8l4��@8��<�y�?�/_C�	�F���J���M�wrQ��T�97X�q�[�b�^��b�UNe�<h�t�k���n���q���t��	x�S{��~�s������c������v��f쇼ha��#Պ��G�����l)��Ԙ��;���t��Wᔼ)M��"���m"����������q]��sŞ�-��h��������b��ɥ�`0��T���E���9e��J̬�f3����������h��	г�P7����������m��?պ�C=�������  �  k�N=�N=�PM=ϛL=S�K=�0K=NzJ=��I=�I=�UH=̝G=��F=4-F=EtE=��D=D=�FC=��B=��A=�A=�W@=^�?=�>=�>=�\==��<= �;=�;=�R:=v�9=��8=>�7==67=�k6=��5=��4=�4=33=�`2=�1=��0=��/=�/=�#.=pC-=`,=�y+=C�*=a�)=��(=޾'=��&=��%=��$=/�#=�"=%�!=B� =;�=�f=�C=4=��=ݷ=�|=�;=��=2�=P=O�=ӑ=�(=��=�B=�
=�B	=˹=�*=j�=��=.Z=�h�<��<:��<�I�<D��<�[�<��<{L�<8��<��<�}�<���<�)�<�v�<r��<*�<�B�<~�<ѵ�<)�<p�<�I�<}u�<ў�<�ŧ<��<��<A/�<5O�<�m�<W��<㧌<�È<O߄<���<?+z<�ar<טj<��b<m
[<�ES<��K<��C<�<<tH4<�,<1�$<�)<�|<��<�/<N"�;��;���;��;��;��;)ɢ;��;92�;�m;S�O;E�2;o;���:U<�:�:�::XO9���E�4�����ź#x����20��gI�}Ab�лz�%j���D��G젻�`������y�»�ͻ+ػ��⻀�컔���] ��/�c�	�Ό���������_1 �+d$���(�L�,�I�0�"k4��?8��<���?�y^C�y�F�Z�J���M��rQ�4�T��7X���[�,�^��b�UOe�@�h�{�k���n�'�q�%�t�x�Z{��~�틀�h	����K���$v��z쇼na��Պ�G��ȸ��)��b������=t�������L��}����!��h���t����\���Ğ��,�����X���fb��qɥ�n0��e��������e���̬��3�����/��di���г��7��4������	n���պ��=��	����  �  F�N=�N=�PM=țL=\�K=�0K=hzJ=��I=�I=�UH=�G=��F=s-F=�tE=2�D=bD=GC=;�B=��A=�A=�W@=z�?=-�>=>=�\==�<=��;=�;=�R:=S�9=��8=�7=�57=�k6=��5=`�4=p4=�23=O`2=ދ1=a�0=��/=v/=�#.=^C-=`,=�y+=V�*=|�)=�(=�'=�&=0�%=��$=q�#=L�"=c�!=�� =v�=g=D=Y=��=�=�|=�;=��=�=�O=%�=��=�(=��=pB=��
=�B	=z�==*=�=E�=�Y=bh�<��<ز�<�I�<��<�[�<��<�L�<V��<�<0~�<���<�)�<w�<��<��<#C�<�~�<V��<��<��<0J�<�u�<��<Ƨ<��<��<7/�<O�<�m�<��<���<�È<�ބ<���<*z<�`r<��j<��b<G	[<tDS<��K<�C<<<�G4<��,<��$<�)<�|<�<20<?#�;|��;O��;���;��;?��;�ˢ;H��;�4�;�m;4�O;"�2;�;]�:5A�:��:�@:b9�	���4���ź\{�����:50��kI�BEb�t�z�/l���F��c�b��_�����»��ͻ,ػ4����컁����\ ��/���	�;��%���s��[0 �c$�~�(�E�,�7�0�$j4��>8�3<��?��]C��F��J���M�rQ�v�T��7X�v�[���^�b�3Pe�.�h���k���n�7�q�(�t�%x�v{��~�V����	���������Nv���쇼_a���Ԋ�RG�������(�����W���s��H���L�����J!��抚���q\���Ğ�^,��Փ��#���Gb��]ɥ�|0�����������e���̬�-4��y�������i��'ѳ�p8���������n��;ֺ�>��N����  �  '�N=�N=�PM=˛L=\�K=�0K=zJ=��I=%I=�UH=,�G=�F=�-F=�tE=_�D=�D=>GC=h�B=��A=�A=X@=��?=B�>=>=�\==�<=��;=�;=�R:=/�9=��8=��7=�57=_k6=��5='�4=C4=�23=%`2=��1=7�0=w�/=[/=�#.=WC-= `,=�y+=a�*=��)=8�(=8�'=B�&=W�%='�$=��#={�"=��!=�� =��=:g=6D=�=��=�=�|=�;=��=�=�O=�=y�=O(=��=>B={�
=zB	=8�=�)=�=�=�Y=�g�<B�<���<II�<���<�[�<��<uL�<u��<?�<m~�<L��<9*�<�w�<@��<�<�C�<�~�<���<�<>�<�J�<:v�<H��<7Ƨ<��<��<C/�<O�<~m�<Ԋ�<U��<$È<}ބ<���<A)z<�_r<��j<�b<j[<�CS<�K<Z�C<r<<GG4<S�,<��$<�)<�|<�<�0<$�;���;���;B��;���;ڴ�;[͢;���;�6�;'m;}�O;�2;;�:E�:4��:�B:&j9�����4���7
ź$��%��;70�nI��Gb�W�z��m���G����c������Ȱ»��ͻ�,ػ�����U����\ �a/���	�ǋ�]�h������/ �Ib$���(���,�e�0�ti4�>8��<�,�?�r]C���F�ŀJ���M�vrQ���T�8X�ދ[�J�^��b��Pe�сh�i�k���n��q���t��x�1{�~������	��L�������kv���쇼_a���Ԋ�*G��e����(��������Ys���ߔ��K������� ��������&\��NĞ�,����������<b��]ɥ�r0����������f��Aͬ��4��͛����Xj���ѳ��8�����z���n���ֺ�l>�������  �  �N=�N=�PM=L=b�K=�0K=�zJ=�I=*I=�UH=H�G=<�F=�-F=�tE=��D=�D=aGC=��B=�A=�A= X@=��?=K�>=>=�\==�<=��;=�;=yR:=�9=��8=��7=�57=:k6=i�5=�4=4=u23=`2=��1=%�0=j�/=R/=�#.=QC-=`,=�y+=k�*=��)=?�(=?�'=]�&=p�%=M�$=��#=��"=��!=М ==Qg=QD=�=��=�=�|=�;=��=�=�O=��=h�=8(=j�=B=W�
=LB	=�=�)=��=��=�Y=�g�<�<d��<'I�<���<�[�<��<�L�<���<U�<o~�<i��<r*�<x�<���<R�<�C�<;�<���<N�<x�<�J�<Gv�<a��<OƧ<�<�<0/�<�N�<Wm�<���<1��<È<Kބ<_��<�(z<;_r<?�j<q�b<�[<2CS<q�K<�C<<<G4<�,<��$<�)<�|<d�<�0<p$�;"��;���;6��;���;��;u΢;"��;�7�;�m;��O;2�2;�;	�:>G�:���:QH:o9J���4�<���`źq���	��90��oI�Jb�4�z��n��I�����d��<���E�»T�ͻ-ػ��?�컟����\ �2/�V�	����<����c��/ ��a$�,�(��,��0��h4��=8�<��?�V]C�}�F���J�[�M��rQ���T�O8X��[�|�^�b�2Qe�\�h��k�#�n���q�y�t�zx��{��~�ӌ��#
��e�������v���쇼ca���Ԋ�G��J���}(���������&s���ߔ�dK��^���� ��E���W��[��Ğ��+����������b��Mɥ��0����������f��cͬ��4������G���j���ѳ�9��W������"o���ֺ��>�������  �  �N=�N=�PM=��L=d�K=�0K=�zJ=�I=6I=�UH=O�G=C�F=�-F=�tE=��D=�D=lGC=��B=�A=A=1X@=��?=A�>=>=�\==�<=��;=�;=rR:=�9=��8=��7=�57=6k6=[�5= �4=4=w23=�_2=��1=�0=\�/=M/=�#.=XC-=`,=�y+=d�*=��)=T�(=I�'=h�&=t�%=W�$=��#=��"=¯!=՜ =̈́=Tg=ZD=�=��=�=�|=�;=��=�=�O=��=X�=+(=a�=	B=X�
=?B	=	�=�)=��=��=�Y=�g�<��<N��<I�<���<�[�<���<�L�<j��<r�<�~�<���<�*�<x�<���<a�<�C�<T�<��<_�<��<�J�<]v�<���<DƧ<�<�<"/�<�N�<Tm�<���<��<�<0ބ<O��<�(z<�^r<��j<.�b<�[<CS<5�K<�C<�<<G4<��,<��$<~)<�|<a�<�0<�$�;���;���;w��;���;E��;�΢;���;�7�;Ym;��O;��2;�;@�:%I�:���:�H:n9���k�4�d���ź#���d���90��oI�XJb��z��n��uI����9e��������»ͻ1-ػ!���컾����\ �P/�E�	�O���ɉ�N���. ��a$��(���,�Ղ0��h4��=8��<��?� ]C�U�F�ĀJ�F�M��rQ���T�V8X��[���^�2b�NQe���h�٫k�T�n���q���t��x��{��~�ߌ��=
��y��������v���쇼ga���Ԋ�.G��,���V(��x������s���ߔ�VK��9���� ��7���F��[�� Ğ��+��i�������"b��Hɥ��0����������%f���ͬ��4�����U���j���ѳ�:9��x������.o���ֺ��>��ݦ���  �  �N=�N=�PM=L=b�K=�0K=�zJ=�I=*I=�UH=H�G=<�F=�-F=�tE=��D=�D=aGC=��B=�A=�A= X@=��?=K�>=>=�\==�<=��;=�;=yR:=�9=��8=��7=�57=:k6=i�5=�4=4=u23=`2=��1=%�0=j�/=R/=�#.=QC-=`,=�y+=k�*=��)=?�(=?�'=]�&=p�%=M�$=��#=��"=��!=М ==Qg=QD=�=��=�=�|=�;=��=�=�O=��=i�=9(=j�=B=X�
=NB	=�=�)=��=��=�Y=�g�<�<h��<+I�<���<�[�<��<�L�<���<X�<r~�<l��<t*�<x�<���<S�<�C�<;�<���<M�<w�<�J�<Ev�<_��<LƧ<�<�<-/�<�N�<Tm�<���</��<È<Jބ<^��<�(z<:_r<?�j<r�b<�[<5CS<t�K<�C<$<<G4<�,<��$<�)<�|<j�<�0<z$�;+��;���;=��;���;��;u΢;!��;�7�;�m;~�O; �2;�;��:G�:���:�G:�l9a��y�4������ź����+��=90�pI�3Jb�P�z��n��I�����d��E���M�»[�ͻ-ػ��D�컣����\ �4/�W�	����=����d��/ ��a$�,�(��,��0��h4��=8�<��?�V]C�}�F���J�[�M��rQ���T�O8X��[�|�^�b�2Qe�\�h��k�#�n���q�y�t�zx��{��~�ӌ��#
��e�������v���쇼ca���Ԋ�G��J���}(���������&s���ߔ�dK��^���� ��E���W��[��Ğ��+����������b��Mɥ��0����������f��cͬ��4������G���j���ѳ�9��W������"o���ֺ��>�������  �  '�N=�N=�PM=˛L=\�K=�0K=zJ=��I=%I=�UH=,�G=�F=�-F=�tE=_�D=�D=>GC=h�B=��A=�A=X@=��?=B�>=>=�\==�<=��;=�;=�R:=/�9=��8=��7=�57=_k6=��5='�4=C4=�23=%`2=��1=7�0=w�/=[/=�#.=WC-= `,=�y+=a�*=��)=8�(=8�'=B�&=W�%='�$=��#={�"=��!=�� =��=:g=6D=�=��=�=�|=�;=��=�=�O=�={�=Q(=��=@B=}�
=|B	=;�=*=�=�=�Y=�g�<J�<���<QI�<���<�[�<��<|L�<{��<E�<r~�<Q��<=*�<�w�<B��<�<�C�<�~�<���<�<;�<�J�<5v�<C��<1Ƨ<��<��<=/�<�N�<ym�<ϊ�<Q��< È<zބ<���<>)z<�_r<��j<	�b<m[<�CS<�K<b�C<{<<RG4<^�,<��$<�)<�|<*�<�0<$�;���;���;O��;���;ߴ�;\͢;���;�6�;m;b�O;��2;�;��:�D�:���:�A:f9�����4�P��
ź���g��{70�XnI�/Hb���z��m���G����c������ذ»�ͻ�,ػ���%��]����\ �d/���	�ɋ�^�j������/ �Jb$���(���,�f�0�ui4�>8��<�,�?�r]C���F�ŀJ���M�vrQ���T�8X�ދ[�J�^��b��Pe�сh�i�k���n��q���t��x�1{�~������	��L�������kv���쇼_a���Ԋ�*G��e����(��������Ys���ߔ��K������� ��������&\��NĞ�,����������<b��]ɥ�r0����������f��Aͬ��4��͛����Xj���ѳ��8�����z���n���ֺ�l>�������  �  F�N=�N=�PM=țL=\�K=�0K=hzJ=��I=�I=�UH=�G=��F=s-F=�tE=2�D=bD=GC=;�B=��A=�A=�W@=z�?=-�>=>=�\==�<=��;=�;=�R:=S�9=��8=�7=�57=�k6=��5=`�4=p4=�23=O`2=ދ1=a�0=��/=v/=�#.=^C-=`,=�y+=V�*=|�)=�(=�'=�&=0�%=��$=q�#=L�"=c�!=�� =v�=g=D=Z=��=�=�|=�;=��=�=�O='�=��=�(=��=sB=��
=�B	=~�=A*=�=I�=�Y=lh�<��<��<�I�<��<�[�<%��<�L�<`��<'�<8~�<���<�)�<�w�<��<��<$C�<�~�<T��<��<��<+J�<�u�<��<�ŧ<��<��<//�<O�<�m�<��<���<zÈ<�ބ<���<*z<�`r<��j<��b<L	[<|DS<��K<(�C<<<�G4<��,<��$<�)<�|<(�<A0<\#�;���;e��;��;"��;F��;�ˢ;E��;�4�;�m;�O;��2;�;��:�@�:��:s?:S\9�����4����ź|�����50��kI��Eb���z�Sl���F����b��x�����»�ͻ,ػD���컍����\ ��/���	�>��(���u��]0 �c$��(�F�,�8�0�$j4��>8�4<��?��]C�	�F��J���M�rQ�w�T��7X�v�[���^�b�3Pe�.�h���k���n�7�q�(�t�%x�v{��~�V����	���������Nv���쇼_a���Ԋ�RG�������(�����W���s��H���L�����J!��抚���q\���Ğ�^,��Փ��#���Gb��]ɥ�|0�����������e���̬�-4��y�������i��'ѳ�p8���������n��;ֺ�>��N����  �  k�N=�N=�PM=ϛL=S�K=�0K=NzJ=��I=�I=�UH=̝G=��F=4-F=EtE=��D=D=�FC=��B=��A=�A=�W@=^�?=�>=�>=�\==��<= �;=�;=�R:=v�9=��8=>�7==67=�k6=��5=��4=�4=33=�`2=�1=��0=��/=�/=�#.=pC-=`,=�y+=C�*=a�)=��(=޾'=��&=��%=��$=/�#=�"=%�!=B� =;�=�f=�C=4=��=޷=�|=�;=��=3�=P=Q�=֑=�(=��=�B=�
= C	=й=�*=o�=��=4Z=�h�<�<G��<�I�<Q��<�[�<+��<�L�<D��<��<�}�<���<�)�<�v�<v��<,�<�B�<~�<ϵ�<%�<k�<�I�<vu�<ɞ�<�ŧ<��<��<7/�<+O�<�m�<N��<ۧ�<�È<J߄<~��<9+z<�ar<טj<��b<s
[<�ES<��K<��C<�<<�H4<�,<E�$<�)<�|<��<�/<q"�;3��;��;��;��;��;,ɢ;��;/2�;em;#�O;	�2;';��:�;�:N�:9:PH9m���4�����qźy������20�hI��Ab�.�z�Qj���D��l젻a��ݡ����»�ͻ++ػԛ⻑�컢���] ��/�h�	�Ҍ���������a1 �-d$���(�M�,�J�0�#k4��?8��<���?�y^C�z�F�Z�J���M��rQ�4�T��7X���[�,�^��b�UOe�@�h�{�k���n�'�q�%�t�x�Z{��~�틀�h	����K���$v��z쇼na��Պ�G��ȸ��)��b������=t�������L��}����!��h���t����\���Ğ��,�����X���fb��qɥ�n0��e��������e���̬��3�����/��di���г��7��4������	n���պ��=��	����  �  ��N=�N=QM=֛L=O�K=q0K=3zJ=��I=�I=EUH=��G=m�F=�,F=�sE=��D=� D=�FC=��B=T�A=PA=�W@=4�?=��>=�>=�\==�<=�;=;=�R:=��9=:�8=��7=~67=l6=L�5=��4=4=T33=�`2=X�1=µ0=��/=�/=�#.=yC-=%`,=�y+=/�*=A�)=в(=��'=��&=��%=��$=��#=��"=ٮ!=�� =��=�f=�C==r�=·=�|=�;=��=G�=7P=�=�=�(=L�=
C=a�
=aC	=+�=�*=͕=��=�Z=�i�<��<ó�<=J�<���<\�<H��<|L�<-��<��<�}�<L��<")�<�v�<��<��<B�<i}�<5��<��<��<HI�<u�<j��<ŧ<��<��<>/�<8O�<�m�<���<F��<DĈ<�߄<��<g,z<�br<�j<;�b<�[<�FS<K<��C<�<<5I4<��,<��$<*<�|<��<p/<
!�;���;���;ܰ�;���;���;�Ƣ;&�;u/�;�m;Z�O;�2;�;M��:�4�:��:M1:+=9���:�4��c źPs��r���.0��dI��=b���z�6h���B���꠻J_������»��ͻ5*ػ0��r�컏���G] �S0���	������ӌ����s2 �\e$�˃(���,�{�0�8l4��@8��<�z�?�/_C�	�F���J���M�wrQ��T�97X�q�[�b�^��b�UNe�<h�t�k���n���q���t��	x�S{��~�s������c������v��f쇼ia��#Պ��G�����l)��Ԙ��;���t��Wᔼ)M��"���m"����������q]��sŞ�-��h��������b��ɥ�`0��T���E���9e��J̬�f3����������h��	г�P7����������m��?պ�C=�������  �  ��N=N=QM=ޛL=J�K=\0K=zJ=k�I=oI=UH=G�G=�F=�,F=�sE=J�D=� D=4FC=m�B=�A=A=rW@=�?=��>=�>=�\==�<=%�;=1;=S:=�9=s�8=��7=�67=nl6=��5=H�4=S4=�33=a2=��1=��0=#�/=�/=$.=�C-=(`,=�y+=�*="�)=��(=w�'=o�&=m�%=-�$=��#=s�"=��!=�� =��=Xf=pC=�=J�=��=�|=|;=��=[�=`P=��=O�=@)=��=gC=��
=�C	=��=W+=/�=M�=�Z=j�<+�<-��<�J�<���<H\�<_��<kL�<��<|�<Y}�<���<�(�<�u�<?��<��<TA�<�|�<���<��<T�<�H�<�t�< ��<=ŧ<\�<��<D/�<TO�<3n�<ҋ�<���<�Ĉ<\��<���<�-z<]dr<u�j<��b<�[<HS<��K<��C<�<<�I4<N�,<��$<N*<�|<b�</<��;��;���;���;��;���;�â;�;�,�;��l;��O;�2;;!��:X-�:��:�(:�,9��2�4��돺��ĺn������*0�a`I�B9b�ݲz��e��K@��y蠻]��&���c�»=�ͻc)ػU��7�컙���}] ��0���	�V����������3 ��f$��(��,�ȇ0��m4��A8� <�^�?��_C���F��J�0 N�qrQ���T��6X��[���^��b�`Me�	~h�S�k�M�n���q���t��x�#{�^~����������������u��U쇼ia��JՊ��G��j����)��L������Nu��┼�M��и��#�����������]���Ş�z-��ʔ�������b���ɥ�T0��2��������d���ˬ��2��������=h��\ϳ��6��坶�\���l���Ժ��<��/����  �  ߺN=(N=.QM=�L=B�K=G0K=�yJ=K�I=7I=�TH=��G=��F=G,F=SsE=��D=- D=�EC= �B=��A=�A=?W@=�?=��>=�>=�\==�<=:�;=O;=JS:=�9=��8= 8=77=�l6=�5=��4=�4=�33=ca2=ی1=5�0=T�/=/=+$.=�C-=)`,=�y+= �*=��)=|�(=C�'=7�&=#�%=��$=I�#=�"=4�!=`� =d�=f=:C=�='�=��=�|=};=��=w�=�P=��=��=�)=�=�C= �
=$D	=��=�+=��=��=9[=�j�<��<���<�J�<!��<r\�<p��<hL�<��<Q�<}�<{��<,(�<fu�<���<T�<�@�<|�<鳾<X�<��<DH�<,t�<���<�ħ<$�<��<E/�<wO�<^n�<*��<��<8ň<���<B��<
/z<�er<�j<�b<n[<WIS<�K<�C<�<<�J4<Ñ,<J�$<m*<�|<�<�.<��;J��;���;<��;r��;���;���;�;�)�;f�l;H�O;��2;o;���:�'�:�ށ:u!:�9���?�4��鏺��ĺ�h��#��X'0��[I��4b�k�z�Pc���=���堻�Z��K�����»ۂͻL(ػ��⻿�컼����] �01��	����w�܎����5 ��g$���(�J�,��0��n4�%C8��<�6�?��`C��F�}�J�T N�xrQ���T�g6X�]�[���^��b�XLe��|h���k��n�G�q�K�t�Zx��{�K~�x��������������u��E쇼oa��cՊ�H������0*������D���u���┼mN��{����#��B���0����^��hƞ��-���������b���ɥ�N0����������d��{ˬ�u2��r���} ���g���γ��5��H������Ql��-Ժ�Q<��Ǥ���  �  �N=CN=AQM=�L=;�K=;0K=�yJ=$�I=I=�TH=��G=��F=�+F=sE=��D=��C=�EC=ߊB=��A=�A=
W@=ř?=��>=�>=�\==�<=N�;=l;=vS:=I�9=��8=R 8=^77=m6=@�5=��4=�4=<43=�a2=�1=n�0=�/=*/=@$.=�C-=%`,=�y+=��*=�)=M�(=	�'=��&=��%=��$=��#=ӻ"=�!=� ='�=�e= C=o=��=s�=�|=|;=��=��=�P=�=Ē=�)=:�=D=t�
=~D	=X�=,=�=�=�[=gk�<6�<��<VK�<b��<�\�<{��<lL�<���<�<�|�<��<�'�<�t�<,��<� �<@�<y{�<M��<��<,�<�G�<�s�<Z��<�ħ<�<x�<=/�<�O�<�n�<���<i��<�ň<n�<���<G0z<�fr<I�j<H�b<�[<sJS<?�K< �C<H<<dK4<?�,<��$<�*<|<��<.<>�;���;��;���;3��;k��;���;��;�&�;@�l;u�O;6�2;2;���:�!�:�ف:9:<9���[4�}珺��ĺ;d������#0�]XI�v0b��z��`���;���㠻/Y��b����»��ͻ;'ػ1��f�������] �~1���	�ʏ�m�ۏ����6 �6i$���(�~�,�W�0��o4�/D8��<�#�?�eaC���F�ςJ�| N��rQ�v�T�6X�̈[�C�^��b�JKe��{h�ߤk���n��q��t�1x��{�G~�􉀼���`���J���~u��0쇼{a��rՊ�PH����*��.������kv�� 㔼O�����W$��ڍ������_���ƞ�W.��a���N��� c���ɥ�Q0��疨�����Kd��(ˬ��1��혯������f��&γ�M5���������k���Ӻ��;��t����  �  (�N=]N=OQM=�L=3�K='0K=�yJ=��I=�I=bTH=��G=L�F=�+F=�rE=c�D=��C=\EC=��B=R�A=wA=�V@=��?=��>=�>=�\==$�<=_�;=�;=�S:=u�9= �8=� 8=�77=Om6=��5=0�4=44=z43=�a2=L�1=��0=��/=G/=V$.=�C-=-`,=�y+=ݏ*=Ƣ)=)�(=�'=��&=��%=_�$=��#=��"=��!=֚ =�=�e=�B=O=��=Z�=�|=s;=��=��=�P=4�=��=*=q�=\D=��
=�D	=��=e,=<�=O�=�[=�k�<��<y��<�K�<���<�\�<���<WL�<���<��<l|�<���<G'�<ut�<���<6 �<�?�<�z�<ò�<C�<��<`G�<js�<��<vħ<��<^�<J/�<�O�<�n�<���<���<ƈ<��<T��<I1z<hr<T�j<l�b<�[<�KS<5�K<��C<<<�K4<��,<��$<�*<f|<��<�-<�;_��;a��;���;��;��;ʻ�;�;�$�;O�l;��O;��2;��;���:��: ց:q:�9���}4�R叺0�ĺ�_�����R 0��TI��,b�+�z�3_���9��⠻'W������»��ͻp&ػ���(������)^ ��1��	�g�� �������47 �Aj$�(���,�Z�0��p4�E8��<���?��aC�#�F� �J�� N�|rQ�N�T��5X�[�[���^�Ub��Je��zh��k���n��q��t�!x��{�C~�����a��������Xu��쇼�a���Պ�rH��5����*��~���8	���v���㔼�O�������$��a���=����_��AǞ��.������{���(c���ɥ�@0��ʖ��m���d���ʬ��1������u����f���ͳ��4��&������Lk��7Ӻ��;������  �  >�N=sN=PQM=�L=5�K=0K=�yJ=��I=�I=5TH=Z�G="�F=�+F=�rE=)�D=o�C=(EC=u�B=(�A=JA=�V@=��?=��>=�>=�\==$�<=e�;=�;=�S:=��9=H�8=� 8=�77=m6=��5=^�4=j4=�43=b2=u�1=Ƕ0=��/=]/=i$.=�C-=.`,=�y+=Ώ*=��)=	�(=��'=��&=��%=1�$=��#=`�"=u�!=�� =��=we=�B=*=��=E�=�|=v;=��=��=�P=P�=�=:*=��=�D=��
=E	=޻=�,=w�=��=\=5l�<�<���<�K�<���<�\�<���<UL�<���<��</|�<~��<�&�<%t�<:��<���<?�<�z�<_��<��<c�<G�<s�<Ĝ�<Iħ<��<]�<H/�<�O�<�n�<䌐<��<aƈ<+�<���<2z<�hr<�j<O�b<�[<MLS<܈K<��C<�<<PL4<�,<��$<�*<u|<z�<d-<
�;3��;��;���;w��;T��;��;�;�"�;��l;��O;��2;��;���:�:Ӂ:�:��9����}4�-㏺��ĺ�Z��p��G0�rRI�*b�A�z��]��M8���࠻�U��旷���»�ͻ�%ػ��=������6^ �2���	�����o������7 ��j$���(�r�,��0��q4��E8��	<�^�?��bC���F�[�J�� N�wrQ�M�T��5X��[�8�^��b��Ie�0zh�8�k���n�G�q�B�t�\x�#{��~�Q�����肃�����Eu��쇼xa���Պ��H��k���(+��Ԛ���	��9w��䔼�O�����:%��Î�������_���Ǟ��.��액�����@c���ɥ�?0��ʖ��C����c���ʬ�S1��7������'f��2ͳ�w4������C���j���Һ�.;��ɣ���  �  L�N=~N=bQM=�L=-�K=0K=�yJ=��I=�I=%TH=>�G=�F=c+F=qrE=�D=J�C=	EC=T�B=�A=:A=�V@=z�?=r�>=�>=�\==.�<=t�;=�;=�S:=��9=c�8=� 8=�77=�m6=ء5=��4=�4=�43=-b2=��1=ֶ0=��/=j/=r$.=�C-=)`,=�y+=ď*=��)=��(=��'=��&=b�%=�$=k�#=B�"=Z�!=�� =��=Ve=�B==��=?�=�|=u;=��=��=�P=b�=%�=I*=ź=�D=�
=0E	=�=�,=��=��=(\=wl�</�<۵�<L�<���<�\�<���<OL�<x��<��<|�<_��<�&�<�s�<���<���<�>�<Pz�<��<��<#�<�F�<�r�<���<%ħ<��<O�<K/�<�O�<�n�< ��<��<�ƈ<h�<���<�2z<kir<��j<��b<[<�LS<X�K<��C<�<<�L4<N�,<E�$<�*<S|<U�<-<��;���;W��;���;a��;,��;鸢;�;�!�;W�l;f�O; �2;I�;���:%�:Ё:�:
�9O���z4�5⏺��ĺ~Z������0�^PI�#(b�`�z��\��7���ߠ�+U�����"�»�ͻ�%ػܗ⻿�����K^ �I2���	�!���������s8 ��k$��(��,���0�4r4�OF8��	<���?��bC���F���J�� N��rQ��T�^5X�Ӈ[�!�^�kb��Ie��yh���k���n���q���t��x��{�:~�������ւ������-u��쇼�a���Պ��H��~���D+�������	��{w��T䔼6P��E���}%��
�������`���Ǟ�/���������Sc���ɥ�;0������.����c��~ʬ�'1�����������e���̳�/4��}�������j���Һ��:�������  �  �N=1 N=0JM=ۓL=@�K=L&K=�nJ=4�I=�H=�FH=ƍG=��F=�F=�`E=A�D=G�C=�/C=�sB=�A=��@=�;@=}?=|�>=�==�;==Iy<=�;=Y�:=�+:=�d9=��8=(�7=M7=�;6=n5=��4=Y�3=W�2=^%2=XN1=*u0=��/=��.=&�-=��,=�,=�(+=%<*=dL)=*Y(=@b'=�g&=�h%=f$=�^#=_S"=C!=	. =�=��=��=��=�u=�?=�=��=My=�*=��=z=-=ܯ= A=�=�P
=c�=�G=��=�'=��=�� =��<SJ�<���<���<��<��<"+�<���<T�<1��<g��<H�<ˡ�<���<�D�<���<���<p�<�T�<p��<Ƕ<���<�-�<{]�<Ŋ�<��<jߟ<��<%-�<�Q�<�u�<Y��<P��<�ۄ<���<u;z<5}r<��j<�c<�F[<w�S<��K<cD<ii<<'�4<�	-<_%<��<H<w<��<���;�w�;i�;7h�;�v�;���;=Ƥ;�	�;a�;��q;ءT;��7;�?;y��:Fa�:�|�:�%,:�#y9m:��B�o��l%��1@��\�B�(���A���Z���r�v��F��=圻wS��	�������sɻEԻЍ޻[���������49����Ϣ�%5�Ͱ���zg�p�"�r�&��*���.��2��6��:��>>� �A�M�E�Y&I���L��+P�9�S�4W�aZ���]��`�Ad�{g�`�j���m���p��t��2w��Dz��Q}�-������m.��*���(��Z�����F���[��}������c��`ԑ��D������Z"��㏗�����_h���ӛ�$>���������z���㢼\L��䴥�h������bV��Ͼ��B'��Ǐ��M����`���ɳ��2���������Vn�� غ�4B�������  �  �N=7 N=3JM=�L=<�K=<&K=�nJ=:�I=#�H=�FH=ύG=��F=�F=�`E=R�D=S�C=�/C=�sB=�A=��@=�;@=}?=|�>=�==�;==Oy<=�;=`�:=�+:=�d9=��8=!�7=<7=�;6=n5=��4=V�3=G�2=Q%2=NN1="u0=��/=��.=,�-=��,=�,=�(+=<*=iL)=2Y(=Ob'=�g&=�h%=#f$=_#=pS"=-C!=. =�=��=��=��=�u=�?=�=��=Ty=�*=��=z=*=ѯ=A=
�=�P
=\�=�G=��=�'=��=�� =��<>J�<���<���<��<��<%+�<f��<M�<:��<|��<�H�<ԡ�<���<�D�<Ύ�<���<��<�T�<���<&Ƕ<���<�-�<�]�<Ί�<���<`ߟ<	�<--�<�Q�<�u�<P��<D��<�ۄ<���<?;z< }r<O�j<jc<�F[<8�S<��K<@D<Li<<�4<�	-<_%<�<5<�v<��<͓�;x�;<i�;~h�;$w�;�;�Ƥ;
�;�a�;�q;��T;j�7;�@;z��:fb�:�|�:�!,:�'y9�:�UA��m���%���@�]���(���A��Z�z�r�v��*F���圻�S��T�������$sɻKԻ��޻+�軔��4���R9��������4������Sg�I�"�,�&���*���.���2�Ͱ6�~:��>>���A�;�E�r&I���L��+P�"�S�%W�aZ���]�/�`�BAd�<{g���j���m�%�p�
t��2w�3Ez�R}�-��ͮ��u.�����(��N�����k���_��}�������b��Uԑ��D������E"������d���Sh��yӛ�>���������z���㢼vL��𴥼V������lV��ؾ��O'��Տ��i���a���ɳ��2���������tn��.غ�CB�������  �  ۵N=) N=#JM=��L=D�K=G&K=�nJ=>�I=/�H=�FH=�G=��F=�F=�`E=_�D=g�C=�/C=�sB=+�A=��@=�;@=}?=��>=�==�;==Iy<=ӵ;=Q�:=�+:=�d9=��8=�7=)7=�;6=�m5=r�4=A�3=/�2=C%2=?N1=u0=��/=��.=�-=��,=�,=�(+=.<*=xL)=7Y(=^b'=�g&=i%=:f$=_#=~S"=;C!=&. ==��=��=��=�u=�?=�=��=Uy=�*=��=z==��=�@=��=�P
=C�=�G=��=s'=ǎ=�� =՚�<J�<���<���<��<���<,+�<r��<o�<G��<���<�H�<��<���<�D�<���<���<��<�T�<���<SǶ<��<.�<�]�<���<��<rߟ<	�<-�<�Q�<|u�<7��< ��<�ۄ<���<�:z<�|r<��j<c<9F[<�S<t�K<�D<i<<��4<�	-<�^%<�<Q<w<��<��;ix�;�i�;+i�; x�;���;vǤ;�
�;?b�;��q;��T;��7;�A;M��:�c�:��:�%,:�4y9�:�*D�o��:'��B��]�(�(���A�?�Z�j�r��v���F��]朻1T������<���xsɻ�Ի��޻���y������9�a������4����T��f���"���&���*�h�.�~�2�n�6�A:�G>>���A��E�$&I�ۮL��+P�S�S�VW�TaZ�ٴ]�w�`��Ad�u{g���j��m�l�p�Pt�+3w��Ez�FR}�5-����.��?���-(��_�����X���6���|�������b��6ԑ�hD��Ƴ��"������?���(h��Gӛ��=����������z���㢼ZL��ᴥ�Y��х��(�V��񾬼r'����������Aa���ɳ��2��蛶�&���n��Hغ�gB��Ь���  �  εN= N=)JM=ۓL=C�K=M&K=�nJ=S�I=G�H=�FH=�G=��F=%F=aE=��D=��C=	0C=�sB=O�A=�@=�;@=,}?=��>=�==�;==Ey<=ص;=B�:=�+:=�d9=m�8=��7=7=�;6=�m5=L�4=�3=�2=%2=N1=�t0=|�/=��.=�-=��,=�,=�(+=/<*=�L)=NY(=wb'=�g&="i%=Yf$=A_#=�S"=iC!=M. =$=��=�=��=�u=�?=�=��=Hy=�*=�=�y=�=��=�@=��=�P
=�=�G=M�=<'=��=�� =���<�I�<L��<[��<�<��<+�<y��<^�<Z��<���<�H�<7��< ��<E�<H��<.��<�<9U�<���<�Ƕ<U��<F.�<�]�<��<*��<zߟ<�<-�<�Q�<cu�<��<幈<Gۄ<K��<L:z<�{r<d�j<Jc<�E[<U�S<��K<nD<�h<<�4<r	-<�^%<�<F<w<��<���;,y�;�j�;?j�;�x�;��;�Ȥ;N�;�c�;w�q;��T;y�7;xD;M��:�f�:���:x),:"5y9:�A�0p��n(���D�|_�M�(�Q�A���Z���r�x��;H��,眻QU���������1tɻ#Ի�޻n�軡������8�9��.��:4�ݯ���mf�P�"�4�&���*���.���2��6��~:��=>�Y�A�ԐE�%&I���L��+P�X�S�_W��aZ�;�]���`�Bd�|g�l�j���m��p��t��3w��Ez��R}�s-��%����.��a���'(��f�����E���<���|��M����b���ӑ�0D��z����!��@��������g��ӛ��=������U���z���㢼QL��ݴ��c��ą��9�V��(����'��6��������a��^ʳ�+3��G���q���n���غ��B������  �  ��N= N=JM=דL=K�K=`&K=oJ=z�I=b�H=�FH=-�G=��F=TF=AaE=æD=��C=80C=#tB=w�A=�@=<@=S}?=��>=)�==�;==@y<=Ƶ;=(�:=w+:=~d9=R�8=��7=�7=;6=�m5= �4=��3=��2=�$2=�M1=�t0=c�/=~�.=��-=��,=�,=�(+=@<*=�L)=pY(=�b'=�g&=Li%=�f$=l_#=�S"=�C!=u. =S=��=5�=ԥ=�u=�?=�=��=By=�*=_�=�y=�=p�=�@=��=LP
=��=iG=�='=j�=S� =:��<wI�<��<��<H�<Ũ�<+�<���<{�<���<���<I�<���<q��<`E�<���<���<g�<�U�<_��<�Ƕ<���<~.�<^�<8��<T��<�ߟ<��<-�<�Q�<8u�<Ǘ�<���<�ڄ<���<�9z<0{r<��j< c<�D[<v�S<�K<�D<h<<�4<�-<�^%<ӷ<[<\w<G�<Е�;z�;�k�;�k�;�z�;���;`ʤ;�;4e�;�q;�T;x�7;�F;���:�l�:d��:�/,:�Cy9�:�vC�Yr��.*���G뺵`���(���A���Z���r�By���I��G蜻�V������֜���tɻ�ԻЎ޻��軒��P����8��������3�L��)��e���"�n�&� �*��.�0�2�S�6�~:�|=>���A�b�E��%I���L��+P�m�S��W��aZ���]�` a�|Bd��|g��j���m���p��t��4w��Fz��S}��-��e����.������M(��p�����(������|�����lb���ӑ��C�����x!��ߎ������wg���қ�P=��h���!��Mz��a㢼,L��д��k��߅��q�V��b����'������=����a���ʳ��3���������Bo���غ��B��E����  �  ��N=��M=JM=ٓL=K�K=i&K=+oJ=��I=��H=+GH=`�G=-�F=�F=�aE=��D=��C=t0C=YtB=��A=O�@=7<@=`}?=��>=,�==�;===y<=��;=�:=V+:=Td9=�8=��7=�7=F;6=Zm5=ݝ4=��3=��2=�$2=�M1=�t0=A�/=f�.=��-=��,=�,=�(+=T<*=�L)=�Y(=�b'=h&=�i%=�f$=�_#=T"=�C!=�. =�=%�=[�=�=�u=�?=�=��=@y=z*=J�=�y=�=5�=u@=V�=P
=��=G=ǹ=�&='�= � =���<I�<���<��<�<���<+�<x��<��<���<��<kI�<Ԣ�<���<�E�<��< ��<��<V�<ː�<Zȶ<���<�.�<A^�<i��<u��<�ߟ<
�<�,�<�Q�<u�<���<B��<�ڄ<���<�8z<9zr<��j<��b<�C[<��S<P�K<D<^g<<��4<�-<\^%<η<V<|w<��<D��;r{�;tm�;Vm�;`|�;���;�̤;�;zg�;,�q;�T;�7;XJ;���:�o�:Ԉ�:&3,:�Ry9�:��D�s��-��	L�gc���(���A��Z��r�'{�� K��ꜻ�W��퓳�L����uɻgԻ�޻���P��M���N8�r��9��3����N��d���"�|�&��*��.�C�2�x�6�[}:��<>�o�A� �E�z%I���L��+P���S��W�DbZ��]�"a�?Cd��}g��j�b�m���p��t�q5w��Gz�QT}�.������&/������j(��w��� ��(������v|���b��?ӑ�oC������� ��n������g��Cқ��<��������*z��6㢼L��д��d�������W������N(��㐯�����Ob��1˳�4�����<���o��Bٺ�@C�������  �  o�N=��M=�IM=ГL=O�K=v&K=GoJ=��I=��H=XGH=��G=d�F=�F=�aE=;�D=:�C=�0C=�tB=طA={�@=d<@=x}?=ֽ>=7�==�;==0y<=��;= �:=,+:=7d9=�8=^�7=g7=;6="m5=��4=n�3=l�2=�$2=�M1=�t0=�/=@�.=��-=��,=�,=�(+=e<*=�L)=�Y(=�b'=Ih&=�i%=�f$=�_#=MT"=
D!=�. =�=Y�=��=+�=v=�?=�=��=6y=]*=4�=�y=~=�=3@=�=�O
=F�=�F=��=v&=ڍ=�� =;��<�H�<I��<���<��<v��<�*�<}��<��<ʄ�<g��<�I�<.��<B��<?F�<���<���<i�<�V�<=��<�ȶ<W��<B/�<�^�<���<���<�ߟ<�<�,�<jQ�<�t�<@��<���<%ڄ<��<�7z<Vyr<��j<��b<�B[<��S<b�K<TD<�f<<ӵ4<^-<^%<��<\<�w<�<5��;�|�;�n�;o�;D~�;���;�Τ;I�;�i�;/�q;�T;��7;�M;���:)t�:���:�8,:<_y9K:��E��t��-1���N��e���(�0�A���Z��r��|���L���뜻�Y������.����vɻtԻX�޻N��O������7������G2�٭�h��c���"���&��*��.�m�2���6��|:��;>���A���E�+%I�u�L��+P�֝S�'W��bZ���]��a�Dd�^~g��j�H�m�� q��t�m6w��Hz�$U}�x.������x/��묄��(���������������D|��}�a���ґ��B��4���z ��퍗������f���ћ��<������i���y��㢼�K��ƴ��p������bW��鿬��(��P�������b���˳��4���������p���ٺ��C��̭���  �  S�N=��M=�IM=͓L=Y�K=�&K=[oJ=зI=��H=�GH=ɎG=��F=	F=�aE=x�D=o�C=�0C=�tB=�A=��@=�<@=�}?=�>=J�==�;==+y<=��;=��:=+:=
d9=��8=(�7=17=�:6=�l5=`�4=.�3=6�2=M$2=dM1=Ut0=�/='�.=��-=��,=�,=�(+=s<*=�L)=�Y(=c'=}h&=�i%=0g$=`#=�T"=CD!="/ =�=��=��=C�=#v=@=�=��=/y=L*=�=cy=M=ծ=�?=��=wO
=��=�F=5�=,&=��=�� =Ƙ�<DH�<���<K��<��<V��<�*�<���<��<
��<���<�I�<���<���<�F�<���<���<��<W�<���<8ɶ<���<�/�<�^�<؋�<���<�ߟ<�<�,�<6Q�<|t�<斌<���<�ل<���<�6z<Kxr<u�j<��b<�A[<��S<��K<�D<	f<<Q�4<�-<�]%<��<{<�w<^�<���;�}�;]p�;�p�;]��;;�Ф;q�;�k�;ذq;K�T;��7;�P;B��:�z�:Đ�:L@,:oy9w:�rG��v���3��(S�=h���(�!�A���Z���r��~��~N��^휻%[��䖳�j����wɻ Ի�޻���B��]����7��������1�������b���"���&�#�*�0�.�j�2���6��{:�;>�9�A�-�E��$I�%�L��+P���S�xW�7cZ�R�]�La��Dd�@g�ٱj�F�m��q��t�a7w�\Iz�V}��.��P����/������(���������ꑊ�����{��6la��oґ��B������ ��s���&���f��Vћ�<��W���/���y���⢼�K������u��4�����W��C����(������x���@c��̳�5�����.���p��ں��C��(����  �  F�N=��M=�IM=̓L=X�K=�&K=foJ=�I=��H=�GH=��G=��F=CF=3bE=��D=��C=(1C=�tB=?�A=��@=�<@=�}?=�>=U�==�;==+y<=��;=��:=�*:=�c9=��8=��7=�7=�:6=�l5='�4=��3=��2=$2=7M1="t0=Ә/=�.=��-=��,=�,=�(+=�<*=�L)=�Y(=2c'=�h&=j%=fg$=Q`#=�T"=�D!=V/ =/=��=��=m�=@v=!@=�=��="y=F*=��=Jy='=��=�?=��=0O
=��=@F=�=�%=V�=Z� =[��<�G�<���<��<p�<H��<�*�<���<��<1��<���<RJ�<��<���<3G�<o��<���<T�<�W�<#��<�ɶ<(��<�/�<"_�<���<޶�<�ߟ<��<�,�<Q�<dt�<���<8��<Zل<&��<�5z<<wr<��j<s�b<�@[<ІS<��K<�D<Pe<<�4<s-<�]%<y�<q<x<��<���;.�;r�;ar�;���;롳;�Ҥ;��;�m�;�q;r�T;��7;�T;���:U�:D��:�E,:uy9q�9�I�ux��=5��
X뺅j�v�(���A�8�Z�+s�E���OP��$�\��,���桾��xɻ}Ի��޻f��\��'���u7�/��i��1�-�����a�͝"���&��*�Q�.�{�2��6��z:��:>���A�َE��$I��L��+P��S��W�wcZ���]�a��Ed��g�ʲj�>�m��q�� t�M8w�4Jz��V}�)/�������/��C����(������ ��ؑ������{���a��ґ�=B��9������쌗������e���Л��;������Zy���⢼�K������|��;���塚�W������S)����������c���̳�w5����������p��wں�JD��{����  �  �N=��M=�IM=œL=\�K=�&K=�oJ=�I= I=�GH="�G=�F=oF=cbE=�D=��C=P1C=*uB=e�A=��@=�<@=�}?=�>=a�==�;==$y<=v�;=��:=�*:=�c9=s�8=��7=�7=a:6=wl5=��4=��3=��2=�#2=M1=
t0=��/=��.=��-=��,=�,=�(+=�<*=M)=Z(=Pc'=�h&=Aj%=�g$=|`#=�T"=�D!=�/ =X=��= �=��=Rv=1@==��=y=4*=��=%y==w�=�?=[�=�N
=~�=F=��=�%=�=%� =��<�G�<U��<ɉ�<>�<)��<�*�<���<�<V��<��<�J�<2��<`��<G�<ɑ�<���<��<�W�<���<�ɶ<a��<0�<S_�<3��<��<�ߟ<��<�,�<�P�<t�<_��<��<ل<���<�4z<�vr<��j<��b<@[<	�S<��K<CD<�d<<b�4<-<L]%<W�<~<Yx<��<E��;6��;s�;�s�;���;q��;sԤ;b�;ko�;�q;5�T;W�7;�V;h��:&��:×�:�J,:a�y9��9��K��z��)9��oZ�9l���(���A�̥Z��s�����mQ�����]��I��������yɻqԻ5�޻���[�����7�������0�����?a��"���&�\�*���.���2�K�6�{z:�F:>�R�A���E�a$I���L��+P��S�'W��cZ�:�]�wa�Fd�Àg���j���m�Zq�G!t�9w��Jz��W}�o/��㰁�.0��y����(���������ő��G���{����`���ё��A��바�=������L���Be���Л�c;���������-y���⢼�K���������^���6塚�W�������)��d���=���d���̳��5��ޞ����Kq���ں��D�������  �  
�N=��M=�IM=ǓL=a�K=�&K=�oJ=�I=: I=�GH=G�G=%�F=�F=�bE=�D=�C=r1C=QuB=��A=�@=�<@=�}?=�>=\�==�;==!y<=s�;=��:=�*:=�c9=K�8=��7=�7=8:6=Ll5=Ɯ4=��3=��2=�#2=�L1=�s0=��/=�.=��-=��,=�,=�(+=�<*=M)=Z(=kc'=�h&=ij%=�g$=�`#=U"=�D!=�/ =q=�=�=��=fv=?@==��=y=%*=��=y=�=U�=c?=9�=�N
=N�=�E=��=}%=�= � =���<HG�<��<���<.�<��<�*�<���<�<k��<7��<�J�<m��<���<�G�<2��<#��<�</X�<̒�<Bʶ<���<W0�<t_�<S��<���<�ߟ<�<�,�<�P�<�s�<.��<���<�؄<���<H4z<�ur<۷j<�b<`?[<��S<e�K<�D<jd<<�4<-<(]%<Y�<�<Ax<0�<���; ��;�s�;!u�;ӄ�;¤�;֤;��;2q�;��q;��T;��7;
Y;���:���:y��:�J,:��y9y�9��J��z��;���\�hn�k�(�U�A�+�Z�.s�����R���񜻬^��q���j���lzɻ�Ի�޻�����ο��7�������0�9��s��`�U�"�"�&���*���.�Y�2���6��y:��9>���A�<�E�[$I��L��+P�?�S� W�dZ���]��a��Fd�.�g��j���m�q��!t��9w�wKz��W}��/�����\0�������(���������ˑ��<��z{����`���ё��A���������J��������d��RЛ�;��}���f��y��d⢼�K������}��m���4塚 X�������)������t���dd��Aͳ�@6��.���T���q��ۺ��D��⮽��  �  �N=��M=�IM=��L=e�K=�&K=�oJ=#�I=H I=HH=T�G=6�F=�F=�bE= �D= �C=�1C=`uB=��A=�@=�<@=�}?=!�>=l�==�;==y<=d�;=��:=�*:=�c9==�8=��7=�7=":6=:l5=��4=��3=��2=�#2=�L1=�s0=��/=ݺ.=��-=��,=�,=�(+=�<*=)M)=&Z(=|c'=�h&=vj%=�g$=�`#=)U"=�D!=�/ =�=�=,�=��=pv=L@==��=y=*=��=y=�=B�=P?=�=�N
=5�=�E=l�=d%=،=�� =~��<"G�<	��<���<�<���<�*�<���<�<���<L��<�J�<���<���<�G�<[��<H��<6�<ZX�<�<]ʶ<���<u0�<�_�<q��<��<�ߟ<��<t,�<�P�<�s�<��<���<�؄<Y��<�3z<�ur<��j<��b<�>[<�S<�K<`D<8d<<�4<�-<�\%<9�<�<�x<m�<A��;���;�t�;�u�;q��;���;�֤;\�;�q�;=�q;!�T;��7;YZ;���:H��:���:�O,:T�y9��9�N��|��P;��2^�!o���(���A�\�Z�&s�y���7S��C�k_��ޚ��ޣ���zɻԻ��޻?��A��y����6�C�����/���;�}`���"���&�u�*�|�.��2�k�6��y:��9>���A���E�'$I�íL��+P�`�S�oW�PdZ���]�$a� Gd���g�s�j���m�Vq�8"t��9w��Kz�QX}��/��3���e0������)��ˢ���������"��Y{��ql`��jё�gA��|������%��������d��-Л��:��Y���J���x��H⢼�K�������������^塚+X������)��ђ�������d��iͳ�Z6��V�������q��5ۺ��D�������  �   �N=��M=�IM=��L=]�K=�&K=�oJ=)�I=N I=	HH=\�G=F�F=�F=�bE=/�D=$�C=�1C=muB=��A=$�@=�<@=�}?=�>=h�==�;=="y<=o�;=��:=�*:=�c9=:�8=��7=�7=:6=)l5=��4=~�3=��2=�#2=�L1=�s0=��/=غ.=��-=��,=�,=�(+=�<*=%M)=*Z(=�c'=�h&=j%=�g$=�`#=6U"=�D!=�/ =�=�=4�=��=rv=J@==��=y=)*=��=�x=�=3�=K?=�=�N
=)�=�E=Y�=Z%=͌=�� =w��<G�<���<|��<�<��<�*�<���<�<���<S��<�J�<���<���<	H�<b��<f��<J�<mX�<��<mʶ<���<�0�<�_�<b��<��<�ߟ<��<�,�<�P�<�s�<���<���<�؄<B��<�3z<Qur<^�j<~�b<�>[<�S<��K<HD<�c<<׳4<�-<A]%<A�<|<vx<V�<v��;΁�;�t�;�u�;��;女;	פ;��;r�;1�q;
�T;s�7;�Z;0��:��:��:�N,:2�y96�9�K��|��5<��$`�Mo�I�(�k�A�ͩZ�As�	����S��m��_�����8����zɻBԻ��޻���f�򻤿���6�R��o���/�Ԫ��6`��"���&�=�*�i�.���2�B�6��y:�g9>���A��E�4$I�حL��+P� �S�\W�adZ��]�\a�Gd���g���j��m��q��"t�:w��Kz�zX}��/��R���u0������)������������.��R{��j]`��Wё�MA��]��������������d��Л��:��M���=���x��V⢼�K���������^���^塚8X��,����)��ݒ�������d���ͳ�z6��t�������q��Dۺ��D������  �  �N=��M=�IM=��L=e�K=�&K=�oJ=#�I=H I=HH=T�G=6�F=�F=�bE= �D= �C=�1C=`uB=��A=�@=�<@=�}?=!�>=l�==�;==y<=d�;=��:=�*:=�c9==�8=��7=�7=":6=:l5=��4=��3=��2=�#2=�L1=�s0=��/=ݺ.=��-=��,=�,=�(+=�<*=)M)=&Z(=|c'=�h&=vj%=�g$=�`#=)U"=�D!=�/ =�=�=,�=��=pv=M@==��=y=*=��=y=�=B�=P?=�=�N
=6�=�E=m�=f%=ٌ=�� =���<%G�<��<���<�<��<�*�<���<�<���<N��<�J�<���<���<�G�<[��<H��<5�<ZX�<�<\ʶ<���<s0�<�_�<n��<��<�ߟ<��<r,�<�P�<�s�<��<���<�؄<X��<�3z<�ur<��j<��b<�>[<�S<�K<cD<;d<<��4<�-< ]%<=�<�<�x<q�<I��;���;�t�;�u�;u��;���;�֤;[�;�q�;5�q;�T;��7;IZ;i��:��:}��:OO,:��y9g�9�~N��|���;��g^�<o���(���A�s�Z�<s�����AS��L�s_��嚳�䣾��zɻ Ի��޻C��D��|����6�D������/���<�}`���"���&�u�*�|�.��2�k�6��y:��9>���A���E�'$I�íL��+P�`�S�oW�PdZ���]�$a� Gd���g�s�j���m�Vq�8"t��9w��Kz�QX}��/��3���e0������)��ˢ���������"��Y{��ql`��jё�gA��|������%��������d��-Л��:��Y���J���x��H⢼�K�������������^塚+X������)��ђ�������d��iͳ�Z6��V�������q��5ۺ��D�������  �  
�N=��M=�IM=ǓL=a�K=�&K=�oJ=�I=: I=�GH=G�G=%�F=�F=�bE=�D=�C=r1C=QuB=��A=�@=�<@=�}?=�>=\�==�;==!y<=s�;=��:=�*:=�c9=K�8=��7=�7=7:6=Ll5=Ɯ4=��3=��2=�#2=�L1=�s0=��/=�.=��-=��,=�,=�(+=�<*=M)=Z(=kc'=�h&=ij%=�g$=�`#=U"=�D!=�/ =r=�=�=��=fv=?@==��=y=&*=��=y=�=W�=d?=;�=�N
=P�=�E=��=%=��=� =���<NG�< ��<���<4�<��<�*�<���<
�<o��<;��<�J�<q��<���<�G�<3��<$��<�<.X�<ʒ�<@ʶ<���<T0�<q_�<O��<���<�ߟ<��<�,�<�P�<�s�<*��<���<�؄<���<F4z<�ur<۷j<�b<b?[<��S<j�K<�D<qd<<�4<-<1]%<b�<�<Ix<9�<ǚ�;.��;t�;*u�;ڄ�;Ƥ�;	֤;��;.q�;|�q;�T;��7;�X;M��:N��:!��:J,:��y9��9��K��z���;��]뺚n���(���A�X�Z�Xs�'����R���񜻻^�����v���wzɻ�Ի�޻����Կ��!7������� 0�:��t��`�U�"�#�&���*���.�Z�2���6��y:��9>���A�<�E�[$I��L��+P�?�S� W�dZ���]��a��Fd�.�g��j���m�q��!t��9w�wKz��W}��/�����\0�������(���������ˑ��<��z{����`���ё��A���������J��������d��RЛ�;��}���f��y��d⢼�K������}��m���4塚 X�������)������t���dd��Aͳ�@6��.���T���q��ۺ��D��⮽��  �  �N=��M=�IM=œL=\�K=�&K=�oJ=�I= I=�GH="�G=�F=oF=cbE=�D=��C=P1C=*uB=e�A=��@=�<@=�}?=�>=a�==�;==$y<=v�;=��:=�*:=�c9=s�8=��7=�7=a:6=wl5=��4=��3=��2=�#2=M1=
t0=��/=��.=��-=��,=�,=�(+=�<*=M)=Z(=Pc'=�h&=Aj%=�g$=|`#=�T"=�D!=�/ =Y=��= �=��=Sv=1@==��=y=5*=��='y==y�=�?=]�=�N
=��=	F=��=�%=�=)� =
��<�G�<]��<҉�<F�<1��<�*�<���<	�<]��<��<�J�<6��<d��<�G�<ˑ�<���<��<�W�<���<�ɶ<]��<0�<N_�<-��<���<�ߟ<��<�,�<�P�<t�<Z��<���<ل<���<�4z<�vr<��j<��b<@[<�S<��K<LD<�d<<m�4<-<X]%<c�<�<ex<	�<Z��;I��;s�;�s�;���;v��;tԤ;_�;eo�;��q;�T;2�7;�V;��:���:F��:�I,:|y95 :��L�i{���9��[뺀l��(���A��Z��s������Q�����]��\��������yɻԻA�޻���d������"7�������0�����@a��"���&�]�*���.���2�K�6�{z:�F:>�S�A���E�b$I���L��+P��S�'W��cZ�:�]�wa�Fd�Àg���j���m�Zq�G!t�9w��Jz��W}�o/��㰁�.0��y����(���������ő��G���{����`���ё��A��바�=������L���Be���Л�c;���������-y���⢼�K���������^���6塚�W�������)��d���=���d���̳��5��ޞ����Kq���ں��D�������  �  F�N=��M=�IM=̓L=X�K=�&K=foJ=�I=��H=�GH=��G=��F=CF=3bE=��D=��C=(1C=�tB=?�A=��@=�<@=�}?=�>=U�==�;==+y<=��;=��:=�*:=�c9=��8=��7=�7=�:6=�l5='�4=��3=��2=$2=7M1="t0=Ә/=�.=��-=��,=�,=�(+=�<*=�L)=�Y(=2c'=�h&=j%=fg$=Q`#=�T"=�D!=V/ =0=��=��=n�=Av="@=�=��=#y=G*=��=Ly=)=��=�?=��=3O
=��=DF=�=�%=Z�=_� =e��<�G�<���<��<{�<R��<�*�<���<��<9��<���<XJ�<���<���<6G�<q��<���<S�<�W�< ��<�ɶ<#��<�/�<_�<�<׶�<�ߟ<��<�,�< Q�<]t�<���<3��<Vل<"��<�5z<9wr<��j<u�b<�@[<׆S<��K<�D<]e<<�4<�-<�]%<��<�<*x<��<���;E�;0r�;qr�;���;�;�Ҥ;��;�m�;��q;M�T;W�7;WT;i��:�~�:���:?D,:�oy9�:�uJ�+y���5���X��j���(�K�A���Z�ts�g���nP��A�\��C��������xɻ�Ի��޻s��g��1���y7�3��m��1�/�����a�Ν"���&��*�R�.�|�2��6��z:��:>���A�َE��$I��L��+P��S��W�wcZ���]�a��Ed��g�ʲj�>�m��q�� t�M8w�4Jz��V}�)/�������/��C����(������ ��ؑ������{���a��ґ�=B��9������쌗������e���Л��;������Zy���⢼�K������|��;���塚�W������S)����������c���̳�w5����������p��wں�JD��{����  �  S�N=��M=�IM=͓L=Y�K=�&K=[oJ=зI=��H=�GH=ɎG=��F=	F=�aE=x�D=o�C=�0C=�tB=�A=��@=�<@=�}?=�>=J�==�;==+y<=��;=��:=+:=
d9=��8=(�7=17=�:6=�l5=`�4=.�3=6�2=M$2=dM1=Ut0=�/='�.=��-=��,=�,=�(+=s<*=�L)=�Y(=c'=}h&=�i%=0g$=`#=�T"=CD!=#/ =�=��=��=C�=#v=@=�=��=0y=M*=�=ey=O=׮=�?=��={O
=��=�F=:�=1&=��=�� =ј�<OH�<���<W��<��<a��<�*�<���<��<��<���<�I�<���<���<�F�<���<���<��<
W�<���<4ɶ<���<{/�<�^�<Ћ�<���<�ߟ<��<�,�<.Q�<ut�<ߖ�<���<�ل<���<�6z<Ixr<u�j<��b<�A[<��S<��K<�D<f<<`�4<�-<�]%<��<�<�w<m�<���;~�;sp�;�p�;j��;���;�Ф;n�;�k�;��q;"�T;��7;eP;���:�y�:��:�>,:(iy9�:�I��w���4���S뺟h�
�(�{�A�O�Z���r��~���N��~휻B[����������xɻ3Ի�޻���N��i����7��������1�������b���"���&�$�*�1�.�k�2���6��{:�;>�:�A�.�E��$I�%�L��+P���S�yW�7cZ�R�]�La��Dd�@g�ٱj�F�m��q��t�a7w�\Iz�V}��.��P����/������(���������ꑊ�����{��6la��oґ��B������ ��s���&���f��Vћ�<��W���/���y���⢼�K������u��4�����W��C����(������x���@c��̳�5�����.���p��ں��C��(����  �  o�N=��M=�IM=ГL=O�K=v&K=GoJ=��I=��H=XGH=��G=d�F=�F=�aE=;�D=:�C=�0C=�tB=طA={�@=d<@=x}?=ֽ>=7�==�;==0y<=��;= �:=,+:=7d9=�8=^�7=g7=;6="m5=��4=n�3=l�2=�$2=�M1=�t0=�/=@�.=��-=��,=�,=�(+=e<*=�L)=�Y(=�b'=Ih&=�i%=�f$=�_#=MT"=D!=�. =�=Z�=��=,�=v=�?=�=��=7y=^*=5�=�y=�=�=6@=�=�O
=J�=�F=��={&=ߍ=�� =F��<�H�<T��<���<��<���<�*�<���<��<ӄ�<p��<�I�<4��<G��<CF�<���<���<h�<�V�<9��<�ȶ<Q��<</�<|^�<���<���<�ߟ<��<�,�<bQ�<�t�<9��<�< ڄ<	��<�7z<Tyr<��j<��b<�B[<��S<l�K<`D<�f<<�4<o-<^%<��<n<�w<�<S��;}�;o�;%o�;R~�;���;�Τ;F�;�i�;�q;�T;��7;�M;;��:�s�:ь�:*7,:Yy9�:��G��u���1��ZO�[f�3�(���A���Z�i�r��|���L���뜻�Y������F����vɻ�Իi�޻^��\�����8������J2�ۭ�j��c���"���&��*� �.�n�2���6��|:��;>���A���E�+%I�v�L��+P�֝S�(W��bZ���]��a�Dd�^~g��j�H�m�� q��t�m6w��Hz�$U}�x.������x/��묄��(���������������D|��}�a���ґ��B��4���z ��퍗������f���ћ��<������i���y��㢼�K��ƴ��p������bW��鿬��(��P�������b���˳��4���������p���ٺ��C��̭���  �  ��N=��M=JM=ٓL=K�K=i&K=+oJ=��I=��H=+GH=`�G=-�F=�F=�aE=��D=��C=t0C=YtB=��A=O�@=7<@=`}?=��>=,�==�;===y<=��;=�:=V+:=Td9=�8=��7=�7=F;6=Zm5=ݝ4=��3=��2=�$2=�M1=�t0=A�/=f�.=��-=��,=�,=�(+=T<*=�L)=�Y(=�b'=h&=�i%=�f$=�_#=T"=�C!=�. =�=%�=\�=�=�u=�?=�=��=Ay={*=K�=�y=�=8�=x@=Y�=P
=��=G=˹=�&=,�=%� =ə�<I�<���<��<!�<���<+�<���<��<���<%��<rI�<ڢ�<���<�E�<��<��<��<V�<Ȑ�<Uȶ<���<�.�<:^�<a��<m��<�ߟ<�<�,�<�Q�<�t�<z��<<��<�ڄ<���<�8z<7zr<��j<��b<�C[<��S<Z�K<D<kg<<��4<�-<m^%<߷<g<�w<��<a��;�{�;�m�;hm�;m|�;ě�;�̤;�;qg�;�q;��T;��7;J;V��:o�:*��:�1,:�Ly9�:�#F��s���-���L��c�V�(��A�j�Z�X�r�M{��CK��%ꜻX�����d����uɻzԻ�޻���]��Y���S8�v��=��3����P��d���"�~�&��*��.�D�2�y�6�[}:��<>�o�A� �E�z%I���L��+P���S��W�DbZ��]�"a�?Cd��}g��j�b�m���p��t�q5w��Gz�QT}�.������&/������j(��w��� ��(������v|���b��?ӑ�oC������� ��n������g��Cқ��<��������*z��6㢼L��д��d�������W������N(��㐯�����Ob��1˳�4�����<���o��Bٺ�@C�������  �  ��N= N=JM=דL=K�K=`&K=oJ=z�I=b�H=�FH=-�G=��F=TF=AaE=æD=��C=80C=#tB=w�A=�@=<@=S}?=��>=)�==�;==@y<=Ƶ;=(�:=w+:=~d9=R�8=��7=�7=;6=�m5= �4=��3=��2=�$2=�M1=�t0=c�/=~�.=��-=��,=�,=�(+=@<*=�L)=pY(=�b'=�g&=Li%=�f$=l_#=�S"=�C!=u. =S=��=5�=ԥ=�u=�?=�=��=Cy=�*=`�=�y=�=r�=�@=��=OP
=��=lG=�=
'=n�=X� =D��<�I�<��<&��<R�<Ϩ�<+�<���<��<���<���<I�<���<v��<cE�<���<���<g�<�U�<\��<�Ƕ<���<x.�<^�<1��<M��<�ߟ<��< -�<�Q�<2u�<���<���<�ڄ<���<�9z<.{r<��j<� c<�D[<|�S<"�K<�D<h<<&�4<	-<�^%<�<j<kw<V�<��;#z�;�k�;�k�;�z�;ř�;bʤ;�;,e�;ʣq;��T;J�7;YF;q��:/l�:˃�:�.,:�>y9!:��D�s���*���H�a�<�(�M�A�B�Z���r�dy���I��d蜻�V������윾��tɻ�Իߎ޻��軝��Z����8��������3�N��+��e���"�o�&��*��.�0�2�S�6�	~:�|=>���A�b�E��%I���L��+P�m�S��W��aZ���]�` a�|Bd��|g��j���m���p��t��4w��Fz��S}��-��e����.������M(��p�����(������|�����lb���ӑ��C�����x!��ߎ������wg���қ�P=��h���!��Mz��a㢼,L��д��k��߅��q�V��b����'������=����a���ʳ��3���������Bo���غ��B��E����  �  εN= N=)JM=ۓL=C�K=M&K=�nJ=S�I=G�H=�FH=�G=��F=%F=aE=��D=��C=	0C=�sB=O�A=�@=�;@=,}?=��>=�==�;==Ey<=ص;=B�:=�+:=�d9=m�8=��7=7=�;6=�m5=L�4=�3=�2=%2=N1=�t0=|�/=��.=�-=��,=�,=�(+=/<*=�L)=NY(=wb'=�g&="i%=Yf$=A_#=�S"=iC!=M. =$=��=�=��=�u=�?=�=��=Hy=�*=��=�y=�=��=�@=��=�P
=
�=�G=P�=?'=��=�� =���<�I�<U��<d��<��<��<+�<���<e�<a��<���<�H�<;��<#��<E�<I��<.��<�<8U�<���<�Ƕ<Q��<A.�<�]�<���<$��<tߟ<��<-�<�Q�<^u�<���<Ṉ<Dۄ<H��<H:z<�{r<d�j<Kc<�E[<[�S<��K<wD<�h<<��4<~	-<�^%<��<R<"w<��<���;?y�;k�;Mj�;	y�; ��;�Ȥ;K�;�c�;b�q;��T;T�7;KD;��:Kf�:)��:n(,:�0y9�:�CB��p��)��eE��_���(���A���Z�&�r�&x��UH��D眻gU������#���Atɻ1Ի�޻y�軫������8�<��1��<4�߯���of�Q�"�5�&���*���.���2��6��~:��=>�Y�A�ԐE�%&I���L��+P�X�S�_W��aZ�;�]���`�Bd�|g�l�j���m��p��t��3w��Ez��R}�s-��%����.��a���'(��f�����E���<���|��M����b���ӑ�0D��z����!��@��������g��ӛ��=������U���z���㢼QL��ݴ��c��ą��9�V��(����'��6��������a��^ʳ�+3��G���q���n���غ��B������  �  ۵N=) N=#JM=��L=D�K=G&K=�nJ=>�I=/�H=�FH=�G=��F=�F=�`E=_�D=g�C=�/C=�sB=+�A=��@=�;@=}?=��>=�==�;==Iy<=ӵ;=Q�:=�+:=�d9=��8=�7=)7=�;6=�m5=r�4=A�3=/�2=C%2=?N1=u0=��/=��.=�-=��,=�,=�(+=.<*=xL)=7Y(=^b'=�g&=i%=:f$=_#=S"=;C!=&. ==��=��=��=�u=�?=�=��=Vy=�*=��=	z==��=A=��=�P
=E�=�G=��=v'=ʎ=�� =ښ�<J�<���<���<��<���<2+�<w��<t�<L��<���<�H�<��<���<�D�<���<���<��<�T�<���<QǶ< ��<.�<�]�<�<��<nߟ<�<
-�<�Q�<xu�<4��<��<�ۄ<���<�:z<�|r<��j<c<;F[<�S<y�K<�D<i<<ɷ4<�	-<�^%<�<Y<w<��<���;vx�;�i�;5i�;x�;���;wǤ;�
�;:b�;��q;r�T;��7;�A;��:{c�:��:�$,:�1y9�:��D��o���'���B�%^�X�(���A�k�Z���r�w���F��n朻@T��ɐ��I����sɻ�Ի �޻���������9�c������4����U��f���"���&���*�i�.��2�o�6�A:�G>>���A��E�$&I�ܮL��+P�S�S�VW�TaZ�ٴ]�w�`��Ad�u{g���j��m�l�p�Pt�+3w��Ez�FR}�5-����.��?���-(��_�����X���6���|�������b��6ԑ�hD��Ƴ��"������?���(h��Gӛ��=����������z���㢼ZL��ᴥ�Y��х��(�V��񾬼r'����������Aa���ɳ��2��蛶�&���n��Hغ�gB��Ь���  �  �N=7 N=3JM=�L=<�K=<&K=�nJ=:�I=#�H=�FH=ύG=��F=�F=�`E=R�D=S�C=�/C=�sB=�A=��@=�;@=}?=|�>=�==�;==Oy<=�;=`�:=�+:=�d9=��8=!�7=<7=�;6=n5=��4=V�3=G�2=Q%2=NN1="u0=��/=��.=,�-=��,=�,=�(+=<*=iL)=2Y(=Ob'=�g&=�h%=#f$=_#=pS"=-C!=. =�=��=��=��=�u=�?=�=��=Ty=�*=��=z=*=ү=A=�=�P
=]�=�G=��=�'=�=�� =��<AJ�<���<���<��<��<(+�<i��<O�<=��<~��<�H�<ա�<���<�D�<Ύ�<���<��<�T�<���<%Ƕ<���<�-�<�]�<̊�<���<^ߟ<�<+-�<�Q�<�u�<N��<B��<�ۄ<���<>;z<}r<O�j<kc<�F[<:�S<��K<CD<Pi<<�4<�	-<#_%< �<9<�v<��<Փ�;x�;Bi�;�h�;'w�;�;�Ƥ;
�;�a�;ݛq;��T;\�7;�@;U��:<b�:�|�:g!,:G&y9T:��A�n�� &��A�7]���(���A�6�Z���r��v��4F���圻�S��[���Ú��*sɻPԻ��޻/�軗��7���T9��������4�°���Sg�J�"�,�&���*���.���2�Ͱ6�~:��>>���A�;�E�r&I���L��+P�"�S�%W�aZ���]�/�`�BAd�<{g���j���m�%�p�
t��2w�3Ez�R}�-��ͮ��u.�����(��N�����k���_��}�������b��Uԑ��D������E"������d���Sh��yӛ�>���������z���㢼vL��𴥼V������lV��ؾ��O'��Տ��i���a���ɳ��2���������tn��.غ�CB�������  �  ��N=�M=2CM=�L=��K=�K=ddJ=ΫI=��H=f9H=�G=O�F=�
F=nOE=ƓD=��C=�C=�]B=��A=��@=y!@=Ha?=1�>=B�==H==HW<=<�;=�:=�:=�;9=r8=��7=��6=�6=�;5=)j4=��3=��2=[�1=
1=�50=�W/=Fw.=S�-=��,=��+=\�*=��)=L�(=�(=E
'=5&=&%=�$=��"=��!=A� =�=�=��=4b=@6=�=��=��=�M=�=p�=.`=�=
�=>;=@�=4Y=�	=_=Q�=�M=��=-&=d� =���<I��< 2�<���<Zl�<���<Є�<[�<n~�<���<V\�<���<�!�<�{�<��<�!�<�m�<ɵ�<��<�:�<~x�<��<��<( �<S�<�<в�<�ߛ<��<�5�<�^�<���<b��<7Մ<���<�Cz<;�r<U�j<�*c<�y[<��S<L<+pD<��<<C 5<�|-<�%<A<z�<�<y�<B  <���;��;��;�A�;�x�;��;`�;���;W v;VY;E�<;�Q ;�;�=�:Q��:�EC:�5�9�Q�����k�����ݺ]y���!�O�:�yNS�(�k�|���ς�����․�h���������Ż�<л��ڻ�����>����V���9�
��b�����Q�c���� �@%��<)�XH-�TB1�Y+5�C9���<���@��5D�R�G�XhK���N��kR���U��CY��\��_��@c�ۃf�S�i���l�^ p��Fs�Kgv���y���|�����X��$܂�c]���܅�IZ��)ֈ�uP��uɋ��@��G���\,��:�����Ԅ������e��}Ԙ��B��!������%�������6`��9ˢ��5��]����
���t��(ߩ�FI��e������������6\���Ƴ�1��盶�����q��fݺ�=I��x����  �  ��N=�M=4CM=�L=}�K=�K=edJ=̫I=��H=f9H=�G=W�F=�
F={OE=ғD=��C=�C=�]B=��A=��@=!@=Ea?=0�>=3�==F==MW<=<�;=�:=�:=�;9=r8=��7=��6=�6=�;5=j4=��3=��2=R�1=1=50=�W/=Kw.=U�-=��,=�+=O�*=v�)=G�(=�(=R
'=6&=,%=$=��"=��!=R� =�=�=��=4b=K6=�=��=��=�M=�=s�=,`=�=�=7;=8�=*Y=�	=_=<�=�M=��=&=[� =���<@��<2�<���<Tl�<���<Є�<=�<g~�<���<[\�<���<�!�<�{�< ��<�!�<�m�<��<*��<�:�<�x�<��<��<' �<S�<݃�<���<�ߛ<��<�5�<�^�<��<Z��<'Մ<���<�Cz<(�r<�j<�*c<�y[<��S<�L<pD<��<<D 5<�|-<�%<+A<\�<O<x�<;  <!��;��;��;7B�;�x�;���;��;��;� v;�VY;x�<;[R ;R;�=�:b��:qBC:�5�9�D��2�'k�c���ݺ�y�N�!��:��NS�k����҂�����"�����������K�Ż�<л��ڻn�什ﻥ����V���>�
�[b�����Q�?��h� ��%��<)�=H-�7B1�9+5�@9���<���@��5D�m�G��hK���N��kR���U��CY��\�/�_��@c���f���i���l�� p�$Gs�Xgv�ցy���|�����X��܂�W]���܅�AZ��&ֈ��P��yɋ�A��?���L,��7������Ȅ������be��^Ԙ��B��������%�������9`��:ˢ��5��o����
���t��ߩ�BI��_������������H\���Ƴ�C1��󛶼���r��tݺ�FI��u����  �  ��N=�M=*CM=�L=��K=�K={dJ=ӫI=��H=p9H=�G=g�F=�
F=�OE=ܓD=��C=�C=�]B=��A=��@=�!@=Na?=E�>=<�==H==IW<=2�;= �:=�:=�;9=�q8=��7=��6=�6=�;5=j4=��3=r�2=C�1=�1=p50=�W/=<w.=I�-=��,=��+=S�*=��)=X�(=�(=_
'=?&=;%=$=��"=��!=]� =$�=�=ǈ=<b=X6=�=��=��=�M=�=h�=`=�=��=#;=+�=Y=��	=_=*�=�M=��=
&=I� =���<��<�1�<��<:l�<���<ʄ�<E�<�~�<���<j\�<���<�!�<	|�<>��<�!�<�m�<��<D��<;�<�x�<)��<�<5 �<=S�<���<ʲ�<�ߛ<v�<�5�<�^�<ꆌ<<��<Մ<o��<\Cz<��r<��j<�*c<Hy[<�S<�L<�oD<��<< 5<�|-<��%<A<g�<<Έ<U  <���;&�;B�;�B�;uy�;¦;)�;���;�!v;�WY;x�<;ES ;5;0?�:���:�EC:n8�9�F����k����ݺ^z���!�߳:�\OS�S�k�m������Q������丯������Ż=л�ڻ��仂�u����V���"�
�"b�����Q����6� ��%��<)�H-��A1��*5�9���<���@�|5D��G�|hK���N��kR���U��CY�'�\�o�_��@c�1�f�ʿi���l�� p�SGs��gv��y��|�ɦ��X��7܂�n]���܅�MZ��&ֈ��P��Pɋ��@��,���3,��!����������n���Pe��CԘ��B��𯛼����������-`��ˢ��5��g����
��	u��.ߩ�_I��w������͇���h\���Ƴ�]1��������)r���ݺ�bI�������  �  ��N=�M=.CM=��L=��K=�K=wdJ=�I=��H=�9H=�G=��F=�
F=�OE= �D=��C=C=�]B=��A=
�@=�!@=^a?=@�>=F�==H==GW<=6�;=��:=�:=�;9=�q8=�7=��6=c6={;5=�i4=��3=_�2=$�1=�1=_50=�W/=2w.=J�-=��,=��+=^�*=��)=\�(=�(=m
'=\&=P%=1$=��"=��!=z� =H�=!�=ڈ=Xb=c6=�=��=��=�M=�=g�=`=�=�=;=�=�X=��	=�^=�=~M=f�=�%=!� =���<��<�1�<_��<8l�<���<���<P�<x~�<���<�\�<��<�!�</|�<|��<
"�<*n�<@��<���<P;�<�x�<f��<'�<d �<>S�< ��<۲�<�ߛ<�<�5�<�^�<Ɔ�<��<�Ԅ<;��<�Bz<R�r<P�j<�)c<�x[<�S<,L<|oD<H�<<�5<�|-<��%<�@<r�<�<��<�  <	��;
�;�;�C�;�z�;æ;b�;���;5$v;�YY;|�<;�T ;�;�A�:���:qIC:8;�9�>��v��k�a����ݺG{���!��:�EQS�g�k�4���B������l������������ŻE=лɲڻ��仲�����V�����
��a�#��<Q�y���� �N%�<)�uG-�lA1��*5��9�S�<�D�@�^5D�4�G�LhK���N��kR���U��CY�d�\���_�8Ac���f��i�V�l�[!p��Gs�'hv�a�y�p�|���Y��N܂��]���܅�LZ��+ֈ�oP��[ɋ��@�����,��蟑����i���+���e��Ԙ�7B���������׈������`��ˢ��5��X����
��u��8ߩ�pI������������I򰼔\��ǳ��1��W���.��Wr���ݺ��I�������  �  ��N=��M=!CM=��L=��K=�K=�dJ=��I= �H=�9H=�G=��F=�
F=�OE='�D=��C=7C=�]B=۟A=$�@=�!@=ta?=L�>=P�==H==@W<=%�;=��:=w:=�;9=�q8=_�7=��6=F6=Y;5=�i4=h�3=B�2=��1=�1=D50=pW/="w.=4�-=��,=��+=g�*=��)=l�(=�(=�
'={&=n%=O$=��"=�!=�� =d�=?�=��=wb=x6=�=��=��=�M==X�=`==΢=�:=��=�X=��	=�^=��=UM=@�=�%=�� =U��<���<�1�<%��<l�<g��<���<[�<�~�<���<�\�<B��<"�<l|�<���<G"�<zn�<���<���<�;�<y�<���<S�<� �<[S�<��<벟<�ߛ<j�<�5�<�^�<���<魈<�Ԅ<���<|Bz<��r<��j<O)c<Px[<x�S<�L<oD<��<<�5<>|-<��%<�@<~�<�<�< <���;��;+�;�D�;�{�;=Ħ;��;ӎ�;�&v;
\Y;��<;�V ;V!;�E�:���:�MC:�>�9�>��3��k�������ݺ;|�W�!���:��RS�A�k����G������~���C���Q�����Ż�=лj�ڻ��们ﻻ���oV�B�X�
��a�����P����"� ��%�u;)��F-��@1�'*5�9���<�ۇ@�5D��G�#hK���N��kR��U�FDY���\�!�_��Ac�H�f���i���l��!p�dHs��hv��y���|�o��IY��v܂��]���܅�ZZ��+ֈ�YP��Aɋ��@��ܶ���+������r��%��������d���Ә��A��z���X������}����_���ʢ��5��M����
��u��gߩ��I��г�����>������\��]ǳ��1������l���r��޺��I��鵽��  �  m�N=��M=CM=��L=��K=�K=�dJ=�I=!�H=�9H= �G=��F=F=�OE=O�D= �C=`C=^B=��A=G�@=�!@=}a?=e�>=Q�==K==AW<=�;=��:=a:=�;9=�q8=B�7=g�6=6=-;5=�i4=A�3=�2=��1=�1=50=VW/=w.=)�-=��,=��+=`�*=��)=~�(=�(=�
'=�&=�%=w$=�"=;�!=�� =��=e�=�=�b=�6==��=��=�M==J�=�_=i=��=�:=��=�X=�	=z^=��=M=�=�%=҉ =���<N��<K1�<���<�k�<S��<���<J�<�~�<���<�\�<���<P"�<�|�<��<�"�<�n�<��<,��<�;�<hy�<ೲ<��<� �<�S�<;��<鲟<�ߛ<X�<u5�<h^�<\��<���<[Ԅ<���<�Az<�r< �j<�(c<}w[<��S<%L<onD<I�<<'5<|-<|�%<�@<u�<�<F�<. <���;��;i�;.F�;F}�;�Ŧ;4!�;y��;�)v;(_Y;}�<;�Y ;�#;�G�:
��:PC:rD�9d.�����k�������ݺU~���!�]�:�RUS���k�p���Z���/��S���9���bº�r�Ż%>л��ڻ��l�����V���#�
��`�4��P�L��i� ��%��:)�GF-�D@1�z)5��9�c�<���@��4D���G�9hK���N��kR�J�U��DY��\���_�4Bc���f�^�i�~�l��"p�Is�Hiv���y�h�|����Y���܂��]���܅�_Z��!ֈ�^P��ɋ��@�������+��j�����҃������id��hӘ��A��$�����e���9����_���ʢ��5��R����
��.u��xߩ��I�����I��|�����8]���ǳ�52�������r��@޺�J��#����  �  Q�N=��M=CM=��L=��K=�K=�dJ=$�I=E�H=�9H='�G=��F=KF=(PE=|�D=R�C=�C=,^B=�A=c�@=�!@=�a?=w�>=V�==T==8W<=�;=��:=F:=�;9=yq8=�7=?�6=�
6=�:5=ii4=�3=��2=��1=s1=50=AW/=�v.="�-=v�,=�+=e�*=��)=��(=�(=�
'=�&=�%=�$=B�"=f�!=�� =��=��=E�=�b=�6= =��=��=�M=�=8�=�_=H=��=�:=��=qX=J�	=G^=j�=�L=ػ=W%=�� =���< ��<1�<���<�k�<.��<���<G�<�~�<��<]�<���<�"�<}�<[��<#�<&o�<@��<���<=<�<�y�<!��<��<� �<�S�<M��<���<�ߛ<?�<`5�<0^�<9��<U��<�ӄ<R��<�@z<^�r<�j<�'c<�v[<(�S<bL<�mD<��<<�5<�{-<<�%<�@<��<�<��<� <���;��;� �;�G�;�~�;�Ǧ;�"�;B��;�,v;>bY;.�<;�[ ;Y&;�K�:n��:}SC:%M�9�/��t�k�D���n�ݺ�����!���:��WS�=�k�����y���w��d�������ú� �Ż�>л˳ڻJ��'ﻝ����U�����
�U`����bO������ �J%�:)�xE-��?1��(5�*9���<��@�|4D�s�G�hK�}�N�lR�d�U��DY�|�\���_��Bc�Q�f��i�!�l�]#p��Is��iv�Z�y��|�����Y���܂��]��݅�uZ��ֈ�SP���ȋ�b@��e���V+��$����������,���d��
Ә�CA��ծ�����'����󟼁_���ʢ��5��E����
��Iu���ߩ��I��(������و��)󰼗]��ȳ��2��F���+��;s���޺�MJ��B����  �  7�N=��M=CM=�L=��K=�K=�dJ=@�I=T�H=
:H=S�G=�F=xF=TPE=��D=}�C=�C=S^B=N�A=��@="@=�a?=��>=c�==R==2W<=�;=��:=&:=m;9=Zq8=�7=�6=�
6=�:5=<i4=�3=��2=��1=Q1=�40=W/=�v.=�-=q�,=��+=p�*=��)=��(=(=�
'=�&=�%=�$=j�"=��!="� =��=��=g�=�b=�6=5=��=��=�M=r=+�=�_=+=e�=x:=`�=?X=�	=
^=4�=�L=��=&%=n� =4��<���<�0�<���<�k�<��<���<R�<�~�<K��<3]�<���<�"�<T}�<���<U#�<�o�<���<���<�<�<z�<w��<	�<+!�<�S�<g��<��<�ߛ<7�<;5�<�]�<<��<�ӄ<���<8@z<��r<c�j<'c< v[<r�S<�L<KmD<c�<<25<t{-<�%<�@<��<<҉< <r �;?
�;0"�;�H�;R��;ɦ;�$�;͓�;0v;eY;��<;[^ ; (;�P�:�:�XC:DP�9�+��~�� k�`���`�ݺ ���!���:�-ZS�˝k�Á�����������������ú���Ż�?л4�ڻ`��[�1����U�?�$�
�`�����N����� ��%�>9)��D-��>1�8(5�k9���<���@�4D�W�G��gK���N�lR���U�:EY� �\���_�yCc���f���i���l�$p��Js��jv��y���|�@���Y��݂�^��݅�Z��ֈ�<P���ȋ�*@��=���$+��Ğ��}��&����󕼩c���Ҙ��@������g��Շ����K_���ʢ�}5��6����
��Su���ߩ�&J��q������ ���|��]��fȳ��2����������s���޺��J�������  �  -�N=��M=�BM=�L=��K=�K=�dJ=U�I=q�H=2:H=o�G=D�F=�F=}PE=ߔD=��C=�C=t^B=n�A=��@="@=�a?=��>=n�==M==6W<=��;=��:=:=K;9=>q8=ɥ7=��6=�
6=�:5=i4=��3=��2=e�1=51=�40=W/=�v.=��-=t�,=��+=s�*=��)=��(=.(=�
'=&=�%=�$=��"=��!=N� =�=�=��=�b=�6=H=��=��=�M=f=+�=�_==L�=M:=>�=X=��	=�]=��=vL=g�=�$=<� =���<i��<�0�<T��<ak�<��<~��<\�<�~�<e��<^]�<*��<(#�<�}�<��<�#�<�o�<��<@��<�<�<Nz�<˴�<J�<Z!�<�S�<���<��<�ߛ<5�<5�<�]�<���<Ӭ�<kӄ<���<�?z<Ƌr<��j<M&c<Mu[<��S<L<�lD<��<<�5<{-<��%<�@<��<G<��<i <i�;��;-#�;PJ�;���;�ʦ;;&�;1��;�3v;�gY;�<;Xa ;%*;�S�:�Ę:O]C:PQ�9���!��#k�������ݺ{��3�!��:��\S�{�k�Nā�5���� ��ˇ��V����ĺ���Ż�?л�ڻ2��w�����U����
��_�M��PN�%��I� ��%��8)�.D-�>1��'5�� 9� �<�R�@��3D�)�G��gK���N�lR���U�pEY�F�\��_��Cc���f�O�i���l��$p�GKs�ikv���y�P�|����6Z��/݂�<^��H݅�tZ��%ֈ�&P���ȋ�@��
����*������?��������Lc��YҘ��@��*���.�������� _��pʢ�h5��9����
��Xu���ߩ�9J������	��f�����9^���ȳ�J3���������s��.ߺ��J��ɶ���  �  �N=��M=�BM=�L=��K=�K=�dJ=f�I=��H=F:H=��G=i�F=�F=�PE= �D=��C=
C=�^B=��A=��@=5"@=�a?=��>=x�==P==/W<=�;=��:=:=6;9=!q8=��7=��6=s
6=�:5=�h4=��3=k�2=E�1=1=�40=�V/=�v.=�-=h�,=��+=z�*=��)=��(=B(='=&=!%=$=��"=��!=m� =*�=�=��=c=�6=Z=��=̐=�M=b=�=�_=�=-�=.:=�=�W=��	=�]=��=ML=A�=�$=� =���<0��<J0�<)��<@k�<���<x��<g�<�~�<���<�]�<X��<X#�<�}�<V��<�#�<,p�<8��<{��<6=�<�z�<���<��<�!�<$T�<���<��<�ߛ<�<�4�<�]�<���<���<(ӄ<_��<�>z<C�r<�j<�%c<�t[<,�S<�L<FlD<y�<<�5<�z-<��%<�@<��<~<Q�<� <_�;A�;8$�;�K�;��;�˦;k'�;v��;	6v;mjY;#�<; c ;,;�V�:xȘ:�aC:�U�9��*#��%k� ����ݺ�����!���:�l^S�E�k�qŁ�����!������U����ź�>�Żd@л<�ڻ~��iﻼ���)U���p�
�	_�����M������ �G%��7)��C-��=1�2'5�g 9���<���@��3D���G��gK���N�/lR�(�U��EY���\�u�_�gDc�!�f���i��l�[%p��Ks��kv��y�˚|�%��bZ��`݂�[^��^݅��Z��"ֈ�P���ȋ��?��ڵ���*��M���������D�c��Ҙ�T@��䭛����]���Y��^��Dʢ�H5��-����
��ou���ߩ�hJ��Ѵ��<����������^��ɳ��3��F���	��&t��mߺ��J��񶽼�  �  �N=��M=�BM=�L=��K=�K=�dJ=o�I=��H=Z:H=��G=�F=�F=�PE=�D=��C=C=�^B=��A=��@=G"@=�a?=��>=u�==W==&W<=�;=��:=�:=';9=q8=��7=��6=N
6=c:5=�h4=w�3=J�2=0�1=�1=�40=�V/=�v.=�-=^�,=��+=y�*=��)=��(=N(=%'=.&=A%=)$=��"=��!=�� =R�=�==!c=7=e=�=Đ=�M=d=�=�_=�=�=:=��=�W=��	=�]=��=)L=�=�$=�� =\��<��<0�<��<<k�<���<���<X�<�~�<���<�]�<x��<�#�<~�<{��<8$�<dp�<���<���<a=�<�z�<��<��<�!�<7T�<���<"��<�ߛ<�<�4�<�]�<j��<o��<�҄<0��<j>z<Êr<y�j<B%c<$t[<��S<%L<�kD<4�<<D5<�z-<��%<}@<��<m<o�<� <��;��;E%�;QL�;��;ͦ;o(�;ٗ�;�7v;dlY;�<;�d ;�-;�X�:�ɘ:�aC:�[�9W��"�%k���I�ݺ����!�<�:��`S���k�fƁ�����"��H���-���ƺ�țŻ�@л��ڻ���@﻽���6U�}�:�
��^����9M�X��)� ��%�}7)� C-�X=1��&5� 9�F�<���@�k3D���G��gK���N�]lR��U��EY���\���_��Dc�t�f�Y�i���l��%p�CLs�xlv���y�&�|����Z���݂�a^��X݅��Z��ֈ�P���ȋ��?�������*��������Y������b���ј�@���������6���8��^��4ʢ�P5��'����
��u���ߩ��J������j��܉��@����^��>ɳ��3������]	��Ut���ߺ�0K������  �  ��N=��M=�BM=�L=��K=�K=�dJ=~�I=��H=h:H=��G=��F=�F=�PE=*�D=��C=/C=�^B=��A=��@=S"@=�a?=��>=��==Y=="W<=ޑ;=z�:=�:=;9=�p8=��7=��6=A
6=V:5=�h4=i�3=:�2=�1=�1=�40=�V/=�v.=ݓ-=X�,=��+=�*=��)=��(=[(=4'=9&=N%=9$=��"=�!=�� =]�="�=ω=)c=7=q=�=͐=�M=c=�=�_=�=	�=
:=��=�W=��	=w]=��=L=�=�$=� =C��<��< 0�<���<k�<���<~��<i�<�<���<�]�<���<�#�<-~�<���<N$�<p�<���<���<�=�<�z�<=��<��<�!�<MT�<���<+��<�ߛ<�
�<�4�<�]�<R��<X��<�҄<��<->z<��r<K�j<%c<�s[<}�S<�L<�kD<��<<#5<�z-<x�%<p@<��<�<��< <[�;f�;�%�;�L�;���;}ͦ;�(�;E��;�8v;hmY;�<;�e ;z.;�Z�:�ʘ:OeC:�]�90#��:%�R)k������ݺ����!�"�:�;aS���k��Ɓ�u���#��É��u���|ƺ��ŻAл��ڻ���5ﻄ���U�M��
��^�m��M����� ��%�G7)��B-�=1�s&5���8��<���@�63D���G��gK���N�llR�`�U�FY��\���_�Ec���f���i���l�&p�wLs��lv�نy�^�|�����Z���݂��^��{݅��Z��ֈ�P���ȋ��?������a*��������7����򕼵b���ј��?��������������^��ʢ�;5������
���u��੼�J������������b����^��]ɳ��3������y	��vt���ߺ�FK��)����  �  ��N=��M=�BM=�L=��K=�K=�dJ=}�I=��H=m:H=��G=��F=�F=�PE=>�D=��C=8C=�^B=��A=��@=O"@=�a?=��>=}�==Q==-W<=�;=|�:=�:=;9=�p8=��7=��6=;
6=F:5=�h4=_�3=4�2=�1=�1=�40=�V/=�v.=ߓ-=e�,=��+={�*=��)=��(=U(=7'=?&=V%=F$=��"=�!=�� =^�=.�=։=/c=7=j=�=ΐ=�M=[=�=�_=�=�=�9=��=�W=}�	=n]=��=L= �=�$=� =>��<˄�<0�<���<*k�<���<l��<a�<�~�<���<�]�<���<�#�<B~�<���<R$�<�p�<���<���<�=�<�z�<I��<��<�!�<BT�<���<!��<�ߛ<�<�4�<�]�<C��<Q��<�҄<���<>z<M�r<�j<�$c<�s[<\�S<�L<�kD<��<<*5<�z-<��%<�@<��<�<��< <V�;��;�%�;GM�;Ą�;�ͦ;�)�;j��;g9v;BnY;��<;f ;E.;sZ�:sʘ:�dC:cZ�9��"��(k����*�ݺ��&�!���:��aS���k�"ǁ���N#����������ƺ��Ż�@л��ڻ���Uﻥ���	U�b��
�z^�V���L����� �L%��6)��B-��<1�R&5���8���<���@�M3D���G��gK���N�7lR�L�U�FY��\��_�Ec�ӈf���i���l�H&p��Ls��lv���y�w�|�ƪ��Z���݂�~^��d݅��Z�� ֈ�P���ȋ��?������Z*���������%����򕼍b���ј��?��������������^��*ʢ�<5��)����
��uu��੼�J������������r����^��vɳ�
4�������	���t���ߺ�HK��<����  �  ��N=��M=�BM=�L=��K=�K=�dJ=~�I=��H=h:H=��G=��F=�F=�PE=*�D=��C=/C=�^B=��A=��@=S"@=�a?=��>=��==Y=="W<=ޑ;=z�:=�:=;9=�p8=��7=��6=A
6=V:5=�h4=i�3=:�2=�1=�1=�40=�V/=�v.=ݓ-=X�,=��+=�*=��)=��(=[(=4'=9&=N%=9$=��"=�!=�� =]�="�=ω=)c=7=q=�=͐=�M=c=�=�_=�=	�=
:=��=�W=��	=w]=��=L=�=�$=� =E��<��<0�<���<k�<���<���<k�<�<���<�]�<���<�#�<.~�<���<O$�<�p�<���<���<=�<�z�<<��<��<�!�<KT�<���<)��<�ߛ<�
�<�4�<�]�<Q��<W��<�҄<��<,>z<��r<K�j<%c<�s[<�S<�L<�kD< �<<&5<�z-<{�%<s@<��<�<��< <`�;k�;�%�;�L�;���;}ͦ;�(�;D��;�8v;`mY;��<;�e ;k.;�Z�:�ʘ:eC:O]�9�%���%��)k�����ݺ(����!�5�:�MaS�ɤk��Ɓ�|���&#��ɉ��{����ƺ�
�ŻAл��ڻ���8ﻆ���U�N��
��^�n��M����� ��%�G7)��B-�=1�s&5���8��<���@�63D���G��gK���N�llR�`�U�FY��\���_�Ec���f���i���l�&p�wLs��lv�نy�^�|�����Z���݂��^��{݅��Z��ֈ�P���ȋ��?������a*��������7����򕼵b���ј��?��������������^��ʢ�;5������
���u��੼�J������������b����^��]ɳ��3������y	��vt���ߺ�FK��)����  �  �N=��M=�BM=�L=��K=�K=�dJ=o�I=��H=Z:H=��G=�F=�F=�PE=�D=��C=C=�^B=��A=��@=G"@=�a?=��>=u�==W==&W<=�;=��:=�:=';9=q8=��7=��6=N
6=c:5=�h4=w�3=J�2=0�1=�1=�40=�V/=�v.=�-=^�,=��+=y�*=��)=��(=N(=%'=.&=A%=)$=��"= �!=�� =R�=�==!c=7=f=�=Đ=�M=d=�=�_=�=�=:=��=�W=��	=�]=��=+L=�=�$=�� =`��<��<0�<��<Ak�<���<���<\�<�~�<���<�]�<{��<�#�<~�<|��<9$�<dp�<���<���<`=�<�z�<��<��<�!�<4T�<���<��<�ߛ<�<�4�<�]�<g��<m��<�҄</��<h>z<r<y�j<C%c<&t[<��S<)L<�kD<9�<<J5<�z-<��%<�@<��<s<u�<� <�;��;K%�;VL�;��;ͦ;m(�;՗�;�7v;TlY;�<;�d ;o-;QX�:=ɘ:`aC:hZ�92$���"��%k������ݺ���C�!�_�:��`S��k�uƁ�#����"��S���8���(ƺ�ЛŻ�@л�ڻ���F�����8U��;�
��^����:M�Y��*� ��%�}7)� C-�X=1��&5� 9�F�<���@�k3D���G��gK���N�]lR��U��EY���\���_��Dc�t�f�Y�i���l��%p�CLs�xlv���y�&�|����Z���݂�a^��X݅��Z��ֈ�P���ȋ��?�������*��������Y������b���ј�@���������6���8��^��4ʢ�P5��'����
��u���ߩ��J������j��܉��@����^��>ɳ��3������]	��Ut���ߺ�0K������  �  �N=��M=�BM=�L=��K=�K=�dJ=f�I=��H=F:H=��G=i�F=�F=�PE= �D=��C=
C=�^B=��A=��@=5"@=�a?=��>=x�==P==/W<=�;=��:=:=6;9=!q8=��7=��6=s
6=�:5=�h4=��3=k�2=E�1=1=�40=�V/=�v.=�-=h�,=��+=z�*=��)=��(=B(='=&=!%=$=��"=��!=m� =+�=�=��=c=�6=Z=��=̐=�M=c=�=�_=�=.�=0:=�=�W=��	=�]=��=OL=D�=�$=� =���<6��<Q0�</��<Fk�<���<~��<m�<�~�<���<�]�<\��<\#�<�}�<X��<�#�<-p�<7��<z��<4=�<�z�<�<��<~!�< T�<���<��<�ߛ<�<�4�<�]�<���<���<%ӄ<]��<�>z<A�r<�j<�%c<�t[<0�S<�L<LlD<��<<�5<�z-<��%<�@<��<�<Y�<� <m�;M�;A$�;�K�;��;�˦;i'�;p��;�5v;VjY;�<;�b ;�+;�V�:Ș:�`C:)T�9���
$��&k�� ��9�ݺ0��	�!���:��^S�s�k��Ł�(����!��ǈ��e����ź�J�Żo@лF�ڻ���q�����,U���r�
�_�����M������ �H%��7)��C-��=1�2'5�g 9���<���@��3D���G��gK���N�/lR�(�U��EY���\�u�_�gDc�!�f���i��l�[%p��Ks��kv��y�˚|�%��bZ��`݂�[^��^݅��Z��"ֈ�P���ȋ��?��ڵ���*��M���������D�c��Ҙ�T@��䭛����]���Y��^��Dʢ�H5��-����
��ou���ߩ�hJ��Ѵ��<����������^��ɳ��3��F���	��&t��mߺ��J��񶽼�  �  -�N=��M=�BM=�L=��K=�K=�dJ=U�I=q�H=2:H=o�G=D�F=�F=}PE=ߔD=��C=�C=t^B=n�A=��@="@=�a?=��>=n�==M==6W<=��;=��:=:=K;9=>q8=ɥ7=��6=�
6=�:5=i4=��3=��2=e�1=51=�40=W/=�v.=��-=t�,=��+=s�*=��)=��(=.(=�
'=&=�%=�$=��"=��!=N� =�=�=��=�b=�6=H=��=��=�M=g=,�=�_==N�=O:=@�=X=��	=�]=�=yL=k�=�$=?� =���<q��<�0�<\��<ik�<��<���<c�<�~�<k��<c]�</��<,#�<�}�< ��<�#�<�o�<��<>��<�<�<Lz�<Ǵ�<F�<V!�<�S�<{��<��<�ߛ<0�<5�<�]�<���<Ь�<hӄ<���<�?z<ŋr<��j<O&c<Qu[<��S<%L<�lD<��<<5<{-<�%<�@<��<R< �<r <z�;��;9#�;XJ�;���;�ʦ;9&�;*��;�3v;�gY;��<;.a ;�);kS�:JĘ:X\C:IO�9l���"� %k�5���_�ݺ���t�!�1�:��\S���k�hā�M���� ��߇��i���ź���Ż�?л�ڻ<�什�����U�	���
��_�O��RN�&��K� ��%��8)�/D-�>1��'5�� 9� �<�S�@��3D�)�G��gK���N�lR���U�pEY�F�\��_��Cc���f�O�i���l��$p�GKs�ikv���y�P�|����6Z��/݂�<^��H݅�tZ��%ֈ�&P���ȋ�@��
����*������?��������Lc��YҘ��@��*���.�������� _��pʢ�h5��9����
��Xu���ߩ�9J������	��f�����9^���ȳ�J3���������s��.ߺ��J��ɶ���  �  7�N=��M=CM=�L=��K=�K=�dJ=@�I=T�H=
:H=S�G=�F=xF=TPE=��D=}�C=�C=S^B=N�A=��@="@=�a?=��>=c�==R==2W<=�;=��:=&:=m;9=Zq8=�7=�6=�
6=�:5=<i4=�3=��2=��1=Q1=�40=W/=�v.=�-=q�,=��+=p�*=��)=��(=(=�
'=�&=�%=�$=j�"=��!="� =��=��=h�=�b=�6=6=��=��=�M=s=-�=�_=-=g�=z:=b�=AX=�	=^=7�=�L=��=*%=r� =<��<Ʌ�<�0�<���<�k�<��<���<Z�<�~�<R��<9]�<���<�"�<X}�<���<W#�<�o�<���<���<�<�<z�<s��<�<&!�<�S�<a��<��<�ߛ<1�<55�<�]�<ꅌ<��<�ӄ<���<4@z<��r<c�j<'c<v[<x�S<�L<SmD<m�<<>5<�{-<+�%<�@<��<)<މ< <� �;O
�;="�;�H�;W��;ɦ;�$�;Ɠ�; 0v;�dY;u�<;-^ ;�';P�:+:�WC: N�965��� ��!k�������ݺk��_�!�۽:�oZS�	�k�8Á����������������ú��Ż�?лA�ڻk��e�:����U�B�'�
�`�����N����� ��%�?9)��D-��>1�9(5�l9���<���@�4D�W�G��gK���N�lR���U�:EY� �\���_�yCc���f���i���l�$p��Js��jv��y���|�@���Y��݂�^��݅�Z��ֈ�<P���ȋ�*@��=���$+��Ğ��}��&����󕼩c���Ҙ��@������g��Շ����K_���ʢ�}5��6����
��Su���ߩ�&J��q������ ���|��]��fȳ��2����������s���޺��J�������  �  Q�N=��M=CM=��L=��K=�K=�dJ=$�I=E�H=�9H='�G=��F=KF=(PE=|�D=R�C=�C=,^B=�A=c�@=�!@=�a?=w�>=V�==T==8W<=�;=��:=F:=�;9=yq8=�7=?�6=�
6=�:5=ii4=�3=��2=��1=s1=50=AW/=�v.="�-=v�,=�+=e�*=��)=��(=�(=�
'=�&=�%=�$=B�"=f�!=�� =��=��=F�=�b=�6= =��=��=�M=�=9�=�_=J=��=�:=��=tX=M�	=J^=m�=�L=ܻ=Z%=�� =���<)��<1�<���<�k�<7��<���<P�<�~�<$��<]�<���<�"�<}�<^��<#�<&o�<?��<���<;<�<�y�<��<��<� �<�S�<G��<�<�ߛ<9�<Z5�<*^�<4��<P��<�ӄ<O��<�@z<\�r<�j<�'c<�v[<.�S<jL<�mD<�<<�5<�{-<I�%<�@<��<�<��<� < �;	�;� �;�G�;�~�;�Ǧ;�"�;:��;�,v;bY;�<;�[ ;"&;�K�:还:_RC:�J�9�9��� �Mk������ݺ׀�1�!�ɻ:��WS�}�k������������|�������ú��Ż�>лٳڻV��2ﻦ����U�����
�X`����cO������ �K%�:)�xE-��?1��(5�*9���<��@�|4D�s�G�hK�}�N�lR�d�U��DY�|�\���_��Bc�Q�f��i�!�l�]#p��Is��iv�Z�y��|�����Y���܂��]��݅�uZ��ֈ�SP���ȋ�b@��e���V+��$����������,���d��
Ә�CA��ծ�����'����󟼁_���ʢ��5��E����
��Iu���ߩ��I��(������و��)󰼗]��ȳ��2��F���+��;s���޺�MJ��B����  �  m�N=��M=CM=��L=��K=�K=�dJ=�I=!�H=�9H= �G=��F=F=�OE=O�D= �C=`C=^B=��A=G�@=�!@=}a?=e�>=Q�==K==AW<=�;=��:=a:=�;9=�q8=B�7=g�6=6=-;5=�i4=A�3=�2=��1=�1=50=VW/=w.=)�-=��,=��+=`�*=��)=~�(=�(=�
'=�&=�%=x$=�"=<�!=�� =��=e�=�=�b=�6==��=��=�M=�=K�=�_=j=��=�:=��=�X=��	=}^=��=!M=�=�%=։ =���<V��<T1�<��<�k�<\��<���<R�<�~�<���<�\�<���<T"�<�|�<��<�"�<�n�<��<+��<�;�<ey�<ܳ�<��<� �<�S�<5��<㲟<�ߛ<R�<o5�<c^�<W��<���<XԄ<���<�Az<�r< �j<�(c<�w[<��S<,L<xnD<S�<<25<|-<��%<�@<��<�<R�<9 <���;�;v�;8F�;K}�;�Ŧ;2!�;r��;�)v;	_Y;V�<;~Y ;V#;IG�:���:OC:/B�9�7����k�m���O�ݺ�~��!���:��US���k�����u���H��j���N���uº���Ż4>л��ڻ��w�����V���&�
��`�6��P�M��j� � %��:)�HF-�D@1�{)5��9�d�<���@��4D���G�9hK���N��kR�J�U��DY��\���_�4Bc���f�^�i�~�l��"p�Is�Hiv���y�h�|����Y���܂��]���܅�_Z��!ֈ�^P��ɋ��@�������+��j�����҃������id��hӘ��A��$�����e���9����_���ʢ��5��R����
��.u��xߩ��I�����I��|�����8]���ǳ�52�������r��@޺�J��#����  �  ��N=��M=!CM=��L=��K=�K=�dJ=��I= �H=�9H=�G=��F=�
F=�OE='�D=��C=7C=�]B=۟A=$�@=�!@=ta?=L�>=P�==H==@W<=%�;=��:=w:=�;9=�q8=_�7=��6=F6=Y;5=�i4=h�3=B�2=��1=�1=D50=pW/="w.=4�-=��,=��+=g�*=��)=l�(=�(=�
'={&=n%=O$=��"=�!=�� =e�=?�=��=xb=x6=�=��=��=�M=�=Y�=`=�=Т=�:=��=�X=��	=�^=��=XM=C�=�%=�� =\��<���<�1�<-��<
l�<n��<���<b�<�~�<���<�\�<G��<"�<o|�<���<H"�<{n�<���<���<�;�<y�<���<O�<� �<VS�<��<岟<�ߛ<e�<~5�<�^�<���<孈<�Ԅ<���<yBz<��r<��j<Q)c<Tx[<}�S<�L<'oD<��<<�5<I|-<��%<�@<��<�<��< <���;��;7�;�D�;�{�;?Ħ;��;͎�;�&v;�[Y;��<;�V ;&!;0E�:���:�LC:�<�9EG��F��k�z���>�ݺ~|���!���:�	SS�y�k�9���`����������V���b���ϗŻ�=лv�ڻ��仵�����rV�E�[�
��a�����P����#� ��%�u;)��F-��@1�(*5�9���<�܇@�5D��G�#hK���N��kR��U�FDY���\�!�_��Ac�H�f���i���l��!p�dHs��hv��y���|�o��IY��v܂��]���܅�ZZ��+ֈ�YP��Aɋ��@��ܶ���+������r��%��������d���Ә��A��z���X������}����_���ʢ��5��M����
��u��gߩ��I��г�����>������\��]ǳ��1������l���r��޺��I��鵽��  �  ��N=�M=.CM=��L=��K=�K=wdJ=�I=��H=�9H=�G=��F=�
F=�OE= �D=��C=C=�]B=��A=
�@=�!@=^a?=@�>=F�==H==GW<=6�;=��:=�:=�;9=�q8=�7=��6=c6={;5=�i4=��3=_�2=$�1=�1=_50=�W/=2w.=J�-=��,=��+=^�*=��)=\�(=�(=m
'=\&=P%=1$=��"=��!=z� =I�="�=ۈ=Yb=c6=�=��=��=�M=�=h�=`=�=�=;=�=�X=��	=�^=�=�M=i�=�%=$� =���<���<�1�<f��<?l�<���<���<V�<}~�<���<�\�<��<�!�<2|�<~��<"�<+n�<@��<���<N;�<�x�<d��<#�<` �<:S�<���<ײ�<�ߛ<z�<�5�<�^�<Æ�<��<�Ԅ<9��<�Bz<P�r<Q�j<�)c<�x[<�S<2L<�oD<O�<<�5<�|-<��%<A<{�<�<Ȉ<�  <��;�;)�;�C�;�z�;æ;`�;���;%$v;�YY;`�<;�T ;�;�A�:2��:�HC:�9�9�E��W��k�������ݺ~{���!��:�uQS���k�I���V������}�����������*�ŻP=лӲڻ��仺�����V�����
��a�%��=Q�z���� �N%�<)�uG-�lA1��*5��9�S�<�D�@�^5D�5�G�LhK���N��kR���U��CY�d�\���_�8Ac���f��i�V�l�[!p��Gs�'hv�a�y�p�|���Y��N܂��]���܅�LZ��+ֈ�oP��[ɋ��@�����,��蟑����i���+���e��Ԙ�7B���������׈������`��ˢ��5��X����
��u��8ߩ�pI������������I򰼔\��ǳ��1��W���.��Wr���ݺ��I�������  �  ��N=�M=*CM=�L=��K=�K={dJ=ӫI=��H=p9H=�G=g�F=�
F=�OE=ܓD=��C=�C=�]B=��A=��@=�!@=Na?=E�>=<�==H==IW<=2�;= �:=�:=�;9=�q8=��7=��6=�6=�;5=j4=��3=r�2=C�1=�1=p50=�W/=<w.=I�-=��,=��+=S�*=��)=X�(=�(=_
'=?&=;%=$=��"=��!=]� =$�=�=ǈ==b=X6=�=��=��=�M=�=h�=`=�= �=$;=,�=Y=��	=_=,�=�M=��=&=K� =���<��<�1�<���<?l�<���<τ�<I�<�~�<���<m\�<���<�!�<|�<?��<�!�<�m�<��<D��<;�<�x�<'��<�<2 �<:S�<���<ǲ�<�ߛ<r�<�5�<�^�<熌<:��<Մ<n��<ZCz<��r<��j<�*c<Jy[<��S<�L<�oD<��<<	 5<�|-<��%<A<m�<�<Ԉ<[  <���;/�;I�;�B�;xy�;¦;(�;���;�!v;�WY;d�<;-S ;;�>�:A��:EC:B7�9qK��n��k�.���]�ݺ�z��!��:�OS�t�k�}���)���^������︯�&�����Ż=л�ڻ��仇�y����V���$�
�#b�����Q����7� ��%��<)�H-��A1��*5�9���<���@�|5D��G�|hK���N��kR���U��CY�'�\�o�_��@c�1�f�ʿi���l�� p�SGs��gv��y��|�ɦ��X��7܂�n]���܅�MZ��&ֈ��P��Pɋ��@��,���3,��!����������n���Pe��CԘ��B��𯛼����������-`��ˢ��5��g����
��	u��.ߩ�_I��w������͇���h\���Ƴ�]1��������)r���ݺ�bI�������  �  ��N=�M=4CM=�L=}�K=�K=edJ=̫I=��H=f9H=�G=W�F=�
F={OE=ғD=��C=�C=�]B=��A=��@=!@=Ea?=0�>=3�==F==MW<=<�;=�:=�:=�;9=r8=��7=��6=�6=�;5=j4=��3=��2=R�1=1=50=�W/=Kw.=U�-=��,=�+=O�*=v�)=G�(=�(=R
'=6&=-%=$=��"=��!=R� =�=�=��=4b=K6=�=��=��=�M=�=s�=,`=�=�=7;=9�=+Y=�	=_==�=�M=��=&=\� =���<B��<2�<���<Vl�<���<ӄ�<?�<i~�<���<]\�<���<�!�<�{�<!��<�!�<�m�<��<*��<�:�<�x�<��<��<& �<S�<ۃ�<���<�ߛ<��<�5�<�^�< ��<Y��<&Մ<���<�Cz<'�r<�j<�*c<�y[<��S<�L<pD<��<<G 5<�|-<�%</A<`�<R<{�<>  <&��;��;��;:B�;�x�;���;��;��;� v;�VY;n�<;NR ;D;~=�:@��:'BC:�4�9DG����yk�����ݺ�y�a�!�#�:��NS�ґk����ق�����(�����������P�Ż�<л��ڻq�仃ﻧ����V���?�
�[b�����Q�@��h� ��%��<)�=H-�7B1�:+5�@9���<���@��5D�m�G��hK���N��kR���U��CY��\�/�_��@c���f���i���l�� p�$Gs�Xgv�ցy���|�����X��܂�W]���܅�AZ��&ֈ��P��yɋ�A��?���L,��7������Ȅ������be��^Ԙ��B��������%�������9`��:ˢ��5��o����
���t��ߩ�BI��_������������H\���Ƴ�C1��󛶼���r��tݺ�FI��u����  �  ��N=�M=f<M=V�L=��K=:K=ZJ=��I=��H=^,H=�qG=T�F=��E=^>E=��D=E�C=`C=�GB=��A=��@=�@=+F?=��>=+�==��<=06<=�o;=��:=��9=M9=�H8=w{7=ܬ6=��5=�
5=K74=�a3=��2=*�1=��0=��/=�/=65.=�O-=�g,=�|+=��*=̝)=K�(=Q�'=��&=W�%=�$=��#=�"=-�!=�{ =�b=�D=�!=o�=��=.�=�`=�"=��=Z�=�E=i�= �=�3=B�=�^=��
=�r	=$�=�o=��=�V=:�=�( =��<���<�|�<�#�<���<�W�<S��<�k�<���<c�<���<:@�<��<f�<�a�<8��<f
�<SX�<~��<	�<I,�<�l�<۩�<��<�<MS�<���<��<��<w�<�H�<2v�<Ӣ�<�΄<i��<�Kz<��r<�j<�Qc<�[<hT<�aL<_�D<N!=<=�5<T�-<W&<��<�8<��<�-<�� <�r�;��;^��;`��;J�;"��;m�;��;yz;z�];�mA;�0%;�'	;3��:sv�:BrY:���9�K�6QҹvdR�fP����кJ�����3�aL�}�d��]|��뉻�z���۠�a��`��������̻,׻�MỲh�hU������S��	�Ť�1-���� �tL�5�#�r�'�ѿ+���/�q�3��7�Yk;�0?���B���F��-J���M�;DQ��T��/X�;�[���^�Hb�]�e�k�h�(l�kJo�2yr���u���x�~�{���~����������1���������N�����Y��`��	���om���Ⓖ�V��ʕ�0<������������������j���؟�(F��2������L���y���zd��kЩ�E<������������밼~W���ó��/��������xu���⺼
P�������  �  ��N=�M=_<M=X�L=��K=<K=ZJ=��I=��H=_,H=�qG=Y�F=��E=f>E=��D=N�C=bC=�GB=��A=��@=�@=!F?=��>=/�==��<=16<=�o;=��:=��9=Q9=�H8=w{7=ڬ6=��5=�
5=974=�a3=��2=.�1=��0=��/=�/=55.=�O-=�g,=�|+=��*=͝)=F�(=M�'=��&=U�%=�$=��#=$�"=.�!=�{ =�b=�D=�!=l�=�=+�=�`=�"=��=a�=�E=i�=��=�3=@�=�^=��
=�r	=$�=�o=��=�V=5�=�( =��<���<�|�<�#�<���<�W�<b��<�k�<���<�b�<���<B@�<��<n�<�a�<K��<d
�<]X�<���<�<U,�<�l�<�<��<�<PS�<���<��<��<y�<�H�<3v�<Ƣ�<�΄<n��<�Kz<��r<��j<�Qc<�[<jT<�aL<=�D<Q!=<2�5<R�-<�V&<��<�8<��<�-<e� <�r�;���;���;���;BJ�;b��;h�;p��;Kyz;��];�mA;�0%;�'	;��:�v�:�sY:)��9��6\ҹfdR�ZP��:�к������3��`L��d��^|��뉻�z���۠����v������ƍ̻#׻N�wh�RU������S�	����7-����z �[L�.�#�h�'���+���/�Z�3��7�Ck;�0?��B���F��-J���M�JDQ��T��/X�:�[���^�/Hb�Q�e�t�h�#l��Jo�Zyr���u���x�y�{���~�	��⋂����5������񒈼F�����m��Y������om���Ⓖ�V��ʕ�1<��y���������������j���؟�7F��8������E���q����d��kЩ�J<������������밼|W���ó��/��������vu���⺼P�������  �  ��N=�M=Z<M=W�L=��K=>K=$ZJ=��I=��H=h,H=�qG=d�F=��E=x>E=��D=`�C=hC=�GB=��A=��@=�@=%F?=��>=.�==��<=-6<=�o;=��:=��9=J9=�H8=o{7=Ȭ6=��5=�
5=+74=�a3=u�2=#�1=��0=��/=�/=+5.=�O-=�g,=�|+=��*=ԝ)=O�(=U�'=ĵ&=`�%=�$=��#=.�"=>�!=�{ =�b=�D=�!=v�=�=3�=�`=�"=��=`�=�E=e�=�=�3=2�=�^=��
=�r	=�=�o=��=�V=�=�( =��<���<�|�<u#�<���<rW�<\��<�k�<���<�b�<���<V@�<'��<��<�a�<m��<�
�<�X�<���<'�<y,�<�l�<��<��<"�<ZS�<���<��<��<u�<�H�<$v�<���<�΄<R��<wKz<b�r<��j<�Qc<��[<'T<�aL<�D<0!=<��5<E�-<�V&<��<�8<��<�-<t� <;s�;B��;��;���;�J�;��;��;��;�yz;��];�nA;�1%;�(	;��:0x�: tY:��9�{�6�ҹ�dR��Q����кn��]���3��aL�T�d�\_|��뉻G{��"ܠ������������̻)׻:N�fh�_U��j���S��	�n��-����a �1L��#�%�'��+���/��3�ė7�
k;��/?���B�p�F��-J���M�_DQ��T��/X�g�[���^�`Hb�z�e���h�Ll��Jo�}yr�ơu��x���{���~����������;������򒈼I������a��C������Tm���Ⓖ�V���ɕ�<��T����������t����j���؟�0F��&������F���p����d��oЩ�_<��&���������밼�W���ó��/��/�������u���⺼3P������  �  }�N=�M=W<M=V�L=��K=@K=*ZJ=��I=��H=u,H=�qG=y�F=��E=�>E=āD=p�C=�C=�GB=��A=��@=�@=8F?=��>=1�==��<=-6<=~o;=��:=��9=:9=H8=Z{7=��6=��5=�
5=74=�a3=e�2=�1=��0=��/=�/=$5.=�O-=�g,=�|+=��*=՝)=X�(=b�'=ǵ&=o�%=,�$=ԫ#=D�"=S�!=�{ =�b=�D=�!=��=�==�=�`=�"=��=[�=�E=U�=�=�3=�=�^=��
=�r	=��=�o=��=�V=
�=f( =��<���<�|�<^#�<���<kW�<Y��<�k�<���<c�<���<e@�<E��<��<b�<���<�
�<�X�<̢�<V�<�,�<�l�<��<��<4�<`S�<���<��<��<\�<�H�<v�<���<�΄<-��<%Kz<��r<G�j<-Qc<A�[<�T<HaL<˿D<� =<ۄ5<�-<�V&<��<�8<��<�-<ð <qs�;���;���;���;aK�;���;��;���;�{z;@�];pA;�2%;�)	;٭�: y�:�uY:f��9��6�ҹ�eR�,R��T�к���k���3��bL���d�`|��쉻�{���ܠ�G��,������2�̻�׻#NỂh�1U��T��kS��	�^���,�x������K���#�Ԫ'�0�+�E�/�۴3���7��j;��/?���B�k�F��-J���M�ZDQ�C�T��/X�|�[��^��Hb�Дe��h��l�Ko��yr�'�u�[�x���{�/�~�<��������N�������@������A��2������4m��vⒼ�V���ɕ��;��/������V���W����j���؟�
F��������?���v����d���Щ�m<��=���������밼�W���ó��/��`�������u���⺼MP��$����  �  s�N=�M=V<M=S�L=��K=IK=3ZJ=��I=��H=�,H=�qG=��F=��E=�>E=�D=��C=�C=HB=��A=��@=�@=FF?=��>=<�==��<=,6<=zo;=��:=��9=#9=kH8=@{7=��6=h�5=�
5= 74=�a3=N�2=��1=~�0=��/=�/=5.=�O-=�g,=�|+=�*=ݝ)=d�(=t�'=ܵ&=��%=>�$=�#=\�"=m�!=�{ =�b=�D=�!=��='�=L�=�`=�"= �=S�=�E=I�=֔=k3=�=�^=��
=�r	=��=�o=��=iV=��=G( =c�<}��<e|�<<#�<l��<]W�<K��<�k�<���<$c�<���<�@�<r��<��<@b�<���<�
�<�X�<��<��<�,�<�l�<=��<�<I�<tS�<���<��<��<L�<�H�<�u�<h��<`΄<���<�Jz<w�r<��j<�Pc<�[<pT<�`L<o�D<� =<��5<��-<�V&<��<�8<Ѱ<�-< � <�s�;���;S��;|��;\L�;���;��;���;�}z;��];�qA;�4%;+	;P��:�z�:�yY:���9=}�6@ҹEgR��R����к�������3�OdL�F�d��a|��퉻P|��qݠ�������������̻�׻NỐh��T����6S�[	���K,�&�����jK�!�#�Y�'�ƾ+���/���3��7��j;�v/?��B�M�F�h-J���M�^DQ�b�T��/X�ǖ[�g�^��Hb�6�e�]�h�,l��Ko�Hzr���u���x�Y�{��~�k��"������Z��� ��򒈼,���$��������m��IⒼXV���ɕ��;������j��"���/����j���؟��E��������6���}����d���Щ��<��i���H��$���
찼�W��ĳ�90������	���u��㺼vP��Q����  �  ^�N=��M=M<M=Q�L=��K=PK=FZJ=ΠI=��H=�,H=�qG=��F=��E=�>E=�D=��C=�C="HB=؈A=��@=�@=SF?=ƃ>=?�==��<=&6<=uo;=��:=v�9=9=RH8=){7=z�6=I�5=q
5=�64=|a3=(�2=ذ1=h�0=��/=�/=5.=�O-=�g,=�|+= �*=�)=t�(=��'=�&=��%=`�$=�#=z�"=��!=| =�b=�D=�!=��=:�=X�=�`=�"=��=P�=�E=@�=��=Q3=��=�^=i�
=dr	=��=^o=��=DV=��=)( =!�<R��<.|�<#�<Z��<EW�<A��<�k�<���<8c�<��<�@�<���<�<ib�<��<,�<#Y�<<��<��<-�<"m�<p��<�<s�<�S�<���<��<��<:�<qH�<�u�<B��<3΄<���<-Jz<�r<5�j<:Pc<F�[<�T<l`L<�D<E =<M�5<��-<�V&<��<�8<�<K.<5� <�t�;J��;P��;���;HM�;Ĭ�;��;֤�;�z;G�];�sA;16%;�,	;���:�}�:&|Y:���9���6�ҹYiR��T����кA�����3�	fL�ϐd��c|�Am}��9ޠ����@�������̻�׻]N�uh��T������R� 	�����+�������J���#�Щ'�D�+�o�/���3���7�Cj;�6/?�A�B� �F�t-J���M��DQ�o�T�90X��[���^�QIb���e���h��l�Lo��zr�	�u�R�x���{���~����L������`�����򒈼+��΋��
���~������l��Ⓖ.V��Gɕ�i;������1��錛�����hj��T؟��E��޲�����;���~����d���Щ��<������m��O���J찼DX��Kĳ�0��ќ��c	��0v��3㺼�P��q����  �  J�N=��M=@<M=Q�L=�K=SK=OZJ=ܠI=�H=�,H=rG=ӶF= �E=�>E=�D=��C=�C=FHB=�A=��@=@=_F?=σ>=@�==��<= 6<=eo;=��:=a�9=�9=.H8={7=^�6=*�5=K
5=�64=[a3=�2=��1=F�0=��/=�/=�4.=�O-=�g,=�|+=�*=�)=}�(=��'=�&=��%=��$='�#=��"=��!=/| =c=�D=�!=��=Q�=i�=�`=�"=��=V�=�E=,�=��=83=��=q^=H�
==r	=��=,o=U�=V=��=( =��<��<�{�<�"�<.��<*W�<P��<�k�<���<Gc�<4��<�@�<Φ�<Y�<�b�<S��<^�<hY�<���<�<I-�<Km�<���<@�<��<�S�<���<��<��<!�<MH�<�u�<���<�̈́<���<�Iz<��r<~�j<�Oc<��[<iT<�_L<~�D<�=<�5<m�-<^V&<��<�8<��<m.<p� <�u�;���;U��;� �;�N�;��;��;@��;�z;��];�uA;8%;�.	;
��:}�: ~Y:��9���6�ҹfkR��V����к&��O���3��gL��d�f|�#X~���ޠ���������w�̻.׻�N�%h뻳T��i���R��	�3���+�
�����GJ��#�[�'���+���/�k�3�d�7��i;��.?��B���F�d-J�z�M��DQ���T�}0X�a�[��^��Ib��e�{�h�l��Lo�]{r���u���x��{�y�~����w�����������ْ��&����������~��N����l���ᒼ�U���ȕ�6;��p��������������Bj�� ؟��E��˲�����*���w����d���Щ��<�������������{찼�X���ĳ��0������	��bv��n㺼�P�������  �  <�N=��M=><M=F�L=�K=`K=[ZJ=�I= �H=�,H=%rG=�F=@�E=?E=J�D=��C=�C=^HB=�A=�@=)@=rF?=݃>=M�==��<=6<=ao;={�:=Q�9=�9=H8=�z7==�6=�5=*
5=�64=2a3=�2=��1=,�0=|�/=u/=�4.=�O-=�g,=�|+=�*=��)=��(=��'="�&=Զ%=��$=D�#=��"=ѐ!=W| =(c=E="=��=f�=z�= a=�"=��=E�=�E=�=��=3=��=U^=�
=r	=\�=	o=-�=�U=s�=�' =��<���<�{�<�"�<��<W�<7��<�k�<��<ac�<P��<A�<��<��<�b�<���<��<�Y�<ɣ�<D�<�-�<�m�<Ԫ�<m�<��<�S�<���<���<��<�<5H�<hu�<ѡ�<�̈́<5��<Iz<ޟr<�j<Oc<!�[<�T<i_L< �D<v=<��5<B�-<MV&<Q�<�8<&�<�.<ñ <>v�;!��;M��;��;�O�;A��;[!�;f��;o�z;��];LxA;t:%;G0	;+��:��:�Y:���9�x�6�ҹQlR�8X��s�к����V�3��iL���d�fg|�Q���B���ߠ�6�����'�����̻s׻�N�zh�dT�����~R�w	�Ԣ�+�������I�w�#���'�!�+�o�/��3�ҕ7�ti;��.?���B���F�<-J���M��DQ�ҿT��0X���[�p�^�5Jb���e���h��l�%Mo��{r�!�u�H�x���{���~��������������'��撈�����������~�����Zl���ᒼ�U���ȕ��:��&������o���w����i���ן��E���������!��������d���Щ��<��⨬����ɀ���찼�X���ĳ�1��`����	���v���㺼Q��;���  �  /�N=��M=8<M=G�L=�K=iK=hZJ=�I=/�H=�,H=<rG=�F=c�E=)?E=l�D=�C=!C=}HB=*�A=�@=:@=�F?=�>=X�==��<=6<=Yo;=h�:=D�9=�9=H8=�z7=!�6=��5=
5=x64=a3=щ2=y�1=�0=h�/=a/=�4.=�O-=�g,=�|+=�*=��)=��(=��'=0�&=�%=��$=k�#=٠"=�!=u| =Bc=@E=-"=��=r�=��=a=�"=�=@�=�E=�=��=3=��=8^=��
=�q	=5�=�n=�=�U=Q�=�' =a�<���<�{�<�"�<���<W�<*��<�k�<	��<�c�<p��<0A�<4��<��<1c�<���<��<�Y�<��<��<�-�<�m�<���<��<��<�S�<Ǉ�<���<��<��<H�<:u�<���<�̈́<���<�Hz<G�r<��j<mNc<��[<OT<�^L<ͽD<=<w�5<��-<.V&<P�<�8<G�<�.<� <�v�;ٖ�;��;��;�P�;0��;�"�;Q��;�z;�];�yA;�;%;�1	;T��:ă�:&�Y:x��9!w�68ҹ�oR�(Y����к�������3�wkL���d�@i|�B�����࠻���M�������̻�׻�N�mh�!T�����<R�!	�����*�=��{��UI���#�2�'���+�Ϳ/���3�q�7�9i;�A.?���B���F�-J���M��DQ��T��0X���[���^��Jb� �e�X�h�5l��Mo�f|r���u���x�/�{��~�������3������!��ꒈ�����������l~������0l��Tᒼ^U���ȕ��:��齃�d��#���I����i���ן�]E������z����������d�� ѩ�=����� ��������X��"ų�E1������
���v���㺼2Q�������  �  !�N=��M=.<M=G�L=	�K=jK=rZJ=�I=F�H=-H=WrG=)�F=y�E=G?E=��D=/�C=7C=�HB=D�A=,�@=P@=�F?=�>=W�==��<=6<=Po;=^�:=4�9=�9=�G8=�z7=�6=��5=�	5=W64=�`3=��2=d�1=��0=Q�/=N/=�4.=�O-=�g,=�|+=�*=�)=��(=ɱ'=G�&= �%=ɳ$=�#=��"=�!=�| =^c=SE=D"=�=��=��=a=�"=��=@�=�E= �=s�=�2=u�=^=��
=�q	=�=�n=��=�U=0�=�' =�<e��<q{�<v"�<���<�V�<)��<�k�<��<�c�<���<ZA�<a��<��<\c�<��<2�<(Z�<=��<��<�-�<�m�<%��<��<��<�S�<͇�<���<��<��<�G�<u�<s��<P̈́<���</Hz<۞r<�j<�Mc<5�[<�T<�^L<P�D<�=<4�5<��-<V&<J�<�8<J�<�.<F� <�w�;���;��;��;�Q�;@��;�#�;z��;Ĉz;�];�{A;�=%;h3	;2��:s��:G�Y:���93K�6>ҹ�pR��Z����к�����B�3��lL�&�d�(k|�򉻿����ᠻ������=���{�̻�׻�N�Kh�T�����
R��	�5��U*�ם�$���H��#���'�8�+�w�/�8�3��7��h;��-?�b�B���F�-J���M��DQ��T�1X�C�[��^��Jb�q�e���h��l�)No��|r��u� �x�}�{���~�A��֌��J������2��㒈�����������C~�������k��ᒼ1U��Bȕ�a:������5����������i���ן�HE������t����������d��ѩ�=��/���8��+���0�7Y��Uų��1��ܝ��X
��w��亼lQ������  �  �N=��M=,<M=D�L=
�K=nK=~ZJ=�I=U�H=-H=jrG=9�F=��E=_?E=��D=F�C=IC=�HB=U�A=:�@=Z@=�F?=��>=W�==��<=6<=No;=V�:=!�9=�9=�G8=�z7=�6=��5=�	5=D64=�`3=��2=T�1=��0=H�/=E/=�4.=�O-=�g,=�|+=�*=�)=��(=α'=V�&=�%=߳$=��#=�"=�!=�| =uc=bE=Y"=�=��=��=a=�"=��=>�=�E=��=d�=�2=k�=^=��
=�q	=��=�n=��=�U=�=�' =��<U��<J{�<]"�<���<�V�<-��<�k�<)��<�c�<���<sA�<���<�<|c�<0��<M�<WZ�<k��<��<.�<n�<G��<��<��<�S�<·�<���<��<��<�G�<	u�<[��<1̈́<���<�Gz<��r<��j<�Mc<Ȧ[<�T<M^L<�D<�=<�5<��-<�U&<;�<�8<Z�<+/<i� <x�;���;���;7�;_R�;��;$�;L��;�z;W�];&}A;�>%;@4	;���:���:�Y:���9�L�6�ҹGrR��\����кH������3�GnL�=�d�:l|�u򉻃����ᠻ��5��z����̻׻O�Sh�T��,���Q��	���*�z�����~H�0�#�t�'�ӻ+�4�/�ݱ3��7��h;��-?�I�B�d�F�-J���M��DQ�#�T�G1X�m�[�8�^�?Kb���e�8�h��l�wNo�#}r�b�u���x���{���~�H������\������;��ْ�����g������5~�������k������U��ȕ�F:��������Ջ�������i���ן�6E��l���f����������d��ѩ�E=��?���O��I���W�kY��tų��1�������
��?w��,亼�Q��'����  �  	�N=��M=+<M=D�L=�K=tK=�ZJ=$�I=\�H= -H=rrG=J�F=��E=h?E=��D=O�C=_C=�HB=^�A=E�@=b@=�F?=��>=\�==��<=6<=Io;=M�:=�9=�9=�G8=�z7=�6=��5=�	5=464=�`3=��2=D�1=��0=<�/=:/=�4.=�O-=�g,=�|+=�*=�)=��(=۱'=`�&=�%=�$=��#=�"=&�!=�| =c=vE=b"=%�=��=��= a=�"= �=;�=�E=��=Z�=�2=[�=�]=��
=�q	=��=�n=��=�U=
�=t' =��<5��<9{�<G"�<���<�V�<'��<�k�<*��<�c�<���<�A�<���<)�<�c�<D��<j�<iZ�<���<�<!.�<(n�<T��<��<��<�S�<Շ�<���<��<��<�G�<�t�<G��<̈́<���<�Gz<K�r<k�j<lMc<��[<[T<^L<�D<n=<ς5<��-<�U&<:�<�8<q�<5/<�� <<x�;e��;���;��;S�;i��;�$�;���;��z;I�];�}A;?%;�4	;"��:!��:�Y:1��91��6�ҹtR��\��m�к������3��nL�L�d�m|��򉻭���m⠻n����������̻E׻�N�Ih��S�����Q��	�ȡ��)�S�����OH�	�#�E�'���+��/���3���7�mh;��-?�&�B�\�F��,J���M��DQ�E�T�f1X���[�m�^�mKb��e�P�h�l��No�j}r���u���x���{���~�d�����n������7��ܒ�����d���r�� ~�������k�������T���Ǖ�):��q��������������oi��}ן�E��g���]����������d��%ѩ�N=��Z���b��g���p�vY���ų��1��!����
��Uw��L亼�Q��E����  �  �N=��M=(<M=>�L=
�K=yK=�ZJ=&�I=Z�H=(-H=srG=J�F=��E=m?E=��D=R�C=^C=�HB=c�A=K�@=b@=�F?=��>=c�==��<=6<=Ho;=P�:=$�9=�9=�G8=�z7=�6=��5=�	5=564=�`3=��2=?�1=��0=7�/=8/=�4.=�O-=�g,=�|+=�*=�)=��(=۱'=^�&= �%=�$=��#=�"=1�!=�| =~c=xE=^"=*�=��=��="a=�"=�=2�=�E=��=a�=�2=V�=�]=��
=�q	=��=�n=��={U=�=n' =��<$��<B{�<M"�<���<�V�<��<�k�<&��<�c�<���<�A�<���<$�<�c�<F��<��<uZ�<���<�<".�<9n�<N��<��<��<�S�<҇�<칛<��<��<�G�<�t�<A��<
̈́<v��<�Gz<%�r<p�j<IMc<��[<DT<�]L<�D<R=<��5<��-<�U&<$�<�8<��<5/<�� <1x�;���;���;��;S�;���;>%�;���;��z;$�];+~A;�?%;�4	;r��:��:��Y:���9 P�6�ҹ>sR�\����к�����S�3�oL���d�m|�:󉻼����⠻e���������̻̐K׻Oốh��S�����Q��	�Ρ��)�Z�����OH�܀#��'���+�ؾ/���3���7�mh;��-?��B�Z�F��,J���M��DQ�L�T�F1X���[���^�eKb��e�X�h�Bl��No�p}r���u���x��{���~�s������f����;��蒈����f���q��~�������k�������T���Ǖ�:��e��������������]i���ן�E��g���V����������d��%ѩ�9=��f���h��n���{�|Y���ų��1��1����
��`w��V亼�Q��R����  �  	�N=��M=+<M=D�L=�K=tK=�ZJ=$�I=\�H= -H=rrG=J�F=��E=h?E=��D=O�C=_C=�HB=^�A=E�@=b@=�F?=��>=\�==��<=6<=Io;=M�:=�9=�9=�G8=�z7=�6=��5=�	5=464=�`3=��2=D�1=��0=<�/=:/=�4.=�O-=�g,=�|+=�*=�)=��(=۱'=`�&=�%=�$=��#=�"=&�!=�| =c=vE=b"=%�=��=��= a=�"= �=<�=�E=��=Z�=�2=[�=�]=��
=�q	=��=�n=��=�U=�=u' =��<6��<;{�<I"�<���<�V�<(��<�k�<+��<�c�<���<�A�<���<*�<�c�<D��<j�<iZ�<���<�<!.�<'n�<S��<��<��<�S�<ԇ�<���<��<��<�G�<�t�<F��<̈́<���<�Gz<K�r<k�j<lMc<��[<\T<	^L<�D<p=<҂5<��-<�U&<=�<�8<s�<8/<�� <@x�;h��;���;��;S�;i��;�$�;���;��z;B�];�}A;u?%;�4	;
��:��:��Y:���9r��6zҹGtR�]����к������3��nL�Y�d�%m|��򉻲���r⠻r����������̻H׻�N�Lh��S�����Q��	�ɡ��)�S�����OH�	�#�F�'���+��/���3���7�mh;��-?�'�B�\�F��,J���M��DQ�E�T�f1X���[�m�^�mKb��e�P�h�l��No�j}r���u���x���{���~�d�����n������7��ܒ�����d���r�� ~�������k�������T���Ǖ�):��q��������������oi��}ן�E��g���]����������d��%ѩ�N=��Z���b��g���p�vY���ų��1��!����
��Uw��L亼�Q��E����  �  �N=��M=,<M=D�L=
�K=nK=~ZJ=�I=U�H=-H=jrG=9�F=��E=_?E=��D=F�C=IC=�HB=U�A=:�@=Z@=�F?=��>=W�==��<=6<=No;=V�:=!�9=�9=�G8=�z7=�6=��5=�	5=D64=�`3=��2=T�1=��0=H�/=E/=�4.=�O-=�g,=�|+=�*=�)=��(=α'=V�&=�%=߳$=��#=�"=�!=�| =uc=bE=Y"=�=��=��=a=�"=��=>�=�E=��=d�=�2=k�=^=��
=�q	= �=�n=��=�U=�=�' =��<Y��<M{�<a"�<���<�V�<0��<�k�<,��<�c�<���<uA�<���<�<}c�<1��<M�<WZ�<k��<��<.�<n�<E��<��<��<�S�<̇�<���<��<��<�G�<u�<Y��</̈́<���<�Gz<��r<��j<�Mc<ʦ[<�T<P^L<�D<�=<�5<��-<�U&<@�<�8<^�<0/<m� <
x�;���;���;;�;aR�;��;$�;J��;�z;K�];}A;�>%;+4	;g��:j��:��Y:���9w�6�ҹ�rR��\��,�кf������3�anL�V�d�Ql|��򉻍��� ⠻��<�������̻	׻	O�Wh�T��/���Q��	���� *�z�����H�0�#�u�'�Ի+�4�/�ݱ3��7��h;��-?�I�B�d�F�-J���M��DQ�#�T�G1X�m�[�8�^�?Kb���e�8�h��l�wNo�#}r�b�u���x���{���~�H������\������;��ْ�����g������5~�������k������U��ȕ�F:��������Ջ�������i���ן�6E��l���f����������d��ѩ�E=��?���O��I���W�kY��tų��1�������
��?w��,亼�Q��'����  �  !�N=��M=.<M=G�L=	�K=jK=rZJ=�I=F�H=-H=WrG=)�F=y�E=G?E=��D=/�C=7C=�HB=D�A=,�@=P@=�F?=�>=W�==��<=6<=Po;=^�:=4�9=�9=�G8=�z7=�6=��5=�	5=W64=�`3=��2=d�1=��0=Q�/=N/=�4.=�O-=�g,=�|+=�*=�)=��(=ɱ'=G�&=�%=ɳ$=�#=��"=�!=�| =^c=SE=D"=�=��=��=a=�"= �=@�=�E= �=t�=�2=v�=^=��
=�q	=�=�n=��=�U=2�=�' = �<i��<v{�<{"�<���<�V�<-��<�k�<��<�c�<���<]A�<c��<��<^c�<��<2�<(Z�<<��<��<�-�<�m�<#��<��<��<�S�<ʇ�<���<��<��<�G�<u�<q��<N̈́<���<,Hz<ڞr<�j<�Mc<7�[<�T<�^L<U�D<�=<:�5<��-<	V&<Q�<�8<Q�</<L� <�w�;���;��;��;�Q�;@��;�#�;v��;��z;��];�{A;�=%;J3	;��:+��:��Y:[��9���6�ҹ�qR��Z���к����i�3�mL�I�d�Ik|��̀���ᠻ�����G�����̻׻�N�Qh�T�����R��	�6��V*�؝�$���H��#���'�8�+�w�/�9�3��7��h;��-?�b�B���F�-J���M��DQ��T�1X�C�[��^��Jb�q�e���h��l�)No��|r��u� �x�}�{���~�A��֌��J������2��㒈�����������C~�������k��ᒼ1U��Bȕ�a:������5����������i���ן�HE������t����������d��ѩ�=��/���8��+���0�7Y��Uų��1��ܝ��X
��w��亼lQ������  �  /�N=��M=8<M=G�L=�K=iK=hZJ=�I=/�H=�,H=<rG=�F=c�E=)?E=l�D=�C=!C=}HB=*�A=�@=:@=�F?=�>=X�==��<=6<=Yo;=h�:=D�9=�9=H8=�z7=!�6=��5=
5=x64=a3=щ2=y�1=�0=h�/=a/=�4.=�O-=�g,=�|+=�*=��)=��(=��'=0�&=�%=��$=k�#=ڠ"=�!=u| =Bc=@E=-"=��=r�=��=a=�"=�=A�=�E=�=��=3=��=:^=��
=�q	=7�=�n=�=�U=T�=�' =g�<���<�{�<�"�<���<W�<0��<�k�<��<�c�<u��<4A�<7��<��<3c�<¹�<��<�Y�<��<��<�-�<�m�<�<��<��<�S�<Ç�<���<��<��<H�<6u�<���<̈́<���<�Hz<F�r<��j<oNc<��[<RT<�^L<ӽD<=<�5<��-<7V&<X�<�8<O�<�.<%� <�v�;��;"��;��;�P�;1��;�"�;L��;�z;��];�yA;�;%;�1	;��:l��:k�Y:���9��6�ҹ�pR��Y��c�к-��� �3��kL��d�hi|�U�����࠻���Z������"�̻�׻�N�th�'T�����>R�#	�����*�>��|��UI���#�2�'���+�Ϳ/���3�q�7�:i;�A.?���B���F�-J���M��DQ��T��0X���[���^��Jb� �e�X�h�5l��Mo�f|r���u���x�/�{��~�������3������!��ꒈ�����������l~������0l��Tᒼ^U���ȕ��:��齃�d��#���I����i���ן�]E������z����������d�� ѩ�=����� ��������X��"ų�E1������
���v���㺼2Q�������  �  <�N=��M=><M=F�L=�K=`K=[ZJ=�I= �H=�,H=%rG=�F=@�E=?E=J�D=��C=�C=^HB=�A=�@=)@=rF?=݃>=M�==��<=6<=ao;={�:=Q�9=�9=H8=�z7==�6=�5=*
5=�64=2a3=�2=��1=,�0=|�/=u/=�4.=�O-=�g,=�|+=�*=��)=��(=��'="�&=Զ%=��$=D�#=��"=ѐ!=W| =(c=E="=��=g�=z�=a=�"=��=F�=�E=�=��=3=��=V^= �
=r	=^�=o=0�=�U=v�=�' =��<���<�{�<�"�<��<W�<=��<�k�<��<gc�<T��<A�<��<��<�b�<���<��<�Y�<ȣ�<B�<-�<�m�<Ъ�<i�<��<�S�<���<���<��<�<1H�<du�<Ρ�<�̈́<2��<Iz<ݟr<�j<
Oc<$�[<�T<o_L<'�D<~=<��5<K�-<VV&<[�<�8</�<�.<˱ <Lv�;-��;W��;��;�O�;B��;X!�;a��;^�z;��];.xA;P:%;0	;ѷ�:���:�Y:?��9��6�ҹ=mR��X����к6��U���3�jL��d��g|�g���U���ߠ�F�����4���ʏ̻}׻�NỂh�kT������R�z	�֢�+���� ���I�x�#���'�"�+�p�/��3�ӕ7�ti;��.?���B���F�=-J���M��DQ�ҿT��0X���[�p�^�5Jb���e���h��l�%Mo��{r�!�u�H�x���{���~��������������'��撈�����������~�����Zl���ᒼ�U���ȕ��:��&������o���w����i���ן��E���������!��������d���Щ��<��⨬����ɀ���찼�X���ĳ�1��`����	���v���㺼Q��;���  �  J�N=��M=@<M=Q�L=�K=SK=OZJ=ܠI=�H=�,H=rG=ӶF= �E=�>E=�D=��C=�C=FHB=�A=��@=@=_F?=σ>=@�==��<= 6<=eo;=��:=a�9=�9=.H8={7=^�6=*�5=K
5=�64=[a3=�2=��1=F�0=��/=�/=�4.=�O-=�g,=�|+=�*=�)=}�(=��'=�&=��%=��$='�#=��"=��!=0| =c=�D=�!=��=Q�=j�=�`=�"=��=V�=�E=-�=��=93=��=s^=J�
=?r	=��=.o=W�=!V=��=
( =��<��<�{�<�"�<5��<0W�<V��<�k�<���<Lc�<9��<�@�<Ҧ�<[�<�b�<T��<_�<hY�<���<
�<F-�<Hm�<���<<�<��<�S�<���<	��<��<�<HH�<�u�<���<�̈́<~��<�Iz<��r<~�j<�Oc<��[<mT<�_L<��D<�=<��5<v�-<hV&<��<�8<��<v.<x� <�u�;��;_��;� �;�N�;��;��;;��;�z;��];�uA;�7%;�.	;���:�:G}Y:J��9��6yҹZlR�MW��E�кa������3��gL��d�4f|�9l~���ޠ������������̻9׻�N�.h뻺T��o���R��	�5���+������HJ��#�\�'���+���/�k�3�d�7��i;��.?��B���F�d-J�z�M��DQ���T�}0X�a�[��^��Ib��e�{�h�l��Lo�]{r���u���x��{�y�~����w�����������ْ��&����������~��N����l���ᒼ�U���ȕ�6;��p��������������Bj�� ؟��E��˲�����*���w����d���Щ��<�������������{찼�X���ĳ��0������	��bv��n㺼�P�������  �  ^�N=��M=M<M=Q�L=��K=PK=FZJ=ΠI=��H=�,H=�qG=��F=��E=�>E=�D=��C=�C="HB=؈A=��@=�@=SF?=ƃ>=?�==��<=&6<=uo;=��:=v�9=9=RH8=){7=z�6=I�5=q
5=�64=|a3=(�2=ذ1=h�0=��/=�/=5.=�O-=�g,=�|+= �*=�)=t�(=��'=�&=��%=`�$=�#=z�"=��!=| =�b=�D=�!=��=:�=Y�=�`=�"=��=Q�=�E=A�==R3=��=�^=k�
=fr	=��=`o=��=GV=��=,( ='�<Y��<5|�<#�<a��<LW�<H��<�k�<���<>c�<��<�@�<���<�<kb�<��<,�<#Y�<;��<��<-�<m�<l��<�<n�<�S�<���< ��<��<5�<mH�<�u�<>��<0΄<���<*Jz<�r<5�j<;Pc<I�[<�T<r`L<�D<L =<U�5<��-<�V&<��<�8<��<T.<=� <�t�;V��;Z��;���;LM�;Ŭ�;��;Ѥ�;�z;0�];�sA;6%;�,	;[��:*}�:U{Y:���9M&�6�ҹEjR�]U��f�кz��+�E�3�<fL���d��c|�V�}��Kޠ����O�����
�̻�׻fN�}h��T������R�"	�����+�������J���#�Щ'�D�+�p�/���3���7�Cj;�6/?�A�B�!�F�t-J���M��DQ�o�T�90X��[���^�QIb���e���h��l�Lo��zr�	�u�R�x���{���~����L������`�����򒈼+��΋��
���~������l��Ⓖ.V��Gɕ�i;������1��錛�����hj��T؟��E��޲�����;���~����d���Щ��<������m��O���J찼DX��Kĳ�0��ќ��c	��0v��3㺼�P��q����  �  s�N=�M=V<M=S�L=��K=IK=3ZJ=��I=��H=�,H=�qG=��F=��E=�>E=�D=��C=�C=HB=��A=��@=�@=FF?=��>=<�==��<=,6<=zo;=��:=��9=#9=kH8=@{7=��6=h�5=�
5= 74=�a3=N�2=��1=~�0=��/=�/=5.=�O-=�g,=�|+=�*=ݝ)=d�(=t�'=ܵ&=��%=>�$=�#=]�"=m�!=�{ =�b=�D=�!=��='�=L�=�`=�"= �=T�=�E=J�=ؔ=l3=�=�^=��
=�r	=��=�o=��=kV=��=J( =h�<���<k|�<B#�<r��<bW�<Q��<�k�<���<)c�<���<�@�<u��<��<Bb�<���<�
�<�X�<��<��<�,�<�l�<:��<��<F�<pS�<���< ��<��<H�<�H�<�u�<e��<]΄<���<�Jz<v�r<��j<�Pc<�[<tT<�`L<u�D<� =<��5<��-<�V&<��<�8<ٰ<.<� < t�;���;[��;���;`L�;���;��;���;�}z;��];�qA;�4%;�*	;���:-z�:1yY:
��9��6�ҹhR�PS���к,����3�}dL�q�d��a|��퉻a|���ݠ�������������̻�׻Nỗh��T����9S�]	���M,�'�����kK�"�#�Z�'�ƾ+���/���3��7��j;�v/?��B�M�F�h-J���M�^DQ�b�T��/X�ǖ[�g�^��Hb�6�e�]�h�,l��Ko�Hzr���u���x�Y�{��~�k��"������Z��� ��򒈼,���$��������m��IⒼXV���ɕ��;������j��"���/����j���؟��E��������6���}����d���Щ��<��i���H��$���
찼�W��ĳ�90������	���u��㺼vP��Q����  �  }�N=�M=W<M=V�L=��K=@K=*ZJ=��I=��H=u,H=�qG=y�F=��E=�>E=āD=p�C=�C=�GB=��A=��@=�@=8F?=��>=1�==��<=-6<=~o;=��:=��9=:9=H8=Z{7=��6=��5=�
5=74=�a3=e�2=�1=��0=��/=�/=$5.=�O-=�g,=�|+=��*=՝)=X�(=b�'=ǵ&=o�%=,�$=ԫ#=D�"=S�!=�{ =�b=�D=�!=��=�==�=�`=�"=��=\�=�E=V�=�=�3=�=�^=��
=�r	=��=�o=��=�V=�=i( =��<���<�|�<c#�<���<pW�<^��<�k�<���<c�<���<h@�<G��<��<b�<���<�
�<�X�<ˢ�<U�<�,�<�l�<��<��<1�<]S�<���<��<��<Y�<�H�<v�<���<�΄<,��<#Kz<��r<G�j<.Qc<C�[<�T<LaL<пD<� =<�5<�-<�V&<��<�8<��<�-<ɰ <{s�;���;���;���;dK�;���;��;���;�{z;/�];�oA;�2%;�)	;���:�x�:auY:$��9��6Gҹ�fR��R����к(������3�#cL���d�5`|��쉻�{���ܠ�S��7�� ���:�̻�׻*NỈh�6U��X��mS��	�_���,�y������K���#�Ԫ'�0�+�F�/�۴3���7��j;��/?���B�k�F��-J���M�ZDQ�C�T��/X�|�[��^��Hb�Дe��h��l�Ko��yr�'�u�[�x���{�/�~�<��������N�������@������A��2������4m��vⒼ�V���ɕ��;��/������V���W����j���؟�
F��������?���v����d���Щ�m<��=���������밼�W���ó��/��`�������u���⺼MP��$����  �  ��N=�M=Z<M=W�L=��K=>K=$ZJ=��I=��H=h,H=�qG=d�F=��E=x>E=��D=`�C=hC=�GB=��A=��@=�@=%F?=��>=.�==��<=-6<=�o;=��:=��9=J9=�H8=o{7=Ǭ6=��5=�
5=+74=�a3=u�2=#�1=��0=��/=�/=+5.=�O-=�g,=�|+=��*=ԝ)=O�(=U�'=ĵ&=`�%=�$=��#=.�"=>�!=�{ =�b=�D=�!=v�=�=4�=�`=�"=��=`�=�E=e�=�=�3=3�=�^=��
=�r	=�=�o=��=�V=!�=�( =��<���<�|�<x#�<���<uW�<_��<�k�<���<�b�<���<X@�<)��<��<�a�<n��<�
�<�X�<���<&�<w,�<�l�<	��<��< �<WS�<���<
��<��<s�<�H�<#v�<���<�΄<Q��<uKz<a�r<��j<�Qc<��[<)T<�aL<	�D<4!=<�5<I�-<�V&<��<�8<��<�-<x� <Cs�;H��;��;���;�J�;��;��;��;�yz;��];�nA;�1%;�(	;֪�:�w�:�sY:��9�@�6�ҹ	eR��Q����к���z��3��aL�m�d�s_|�
쉻Q{��+ܠ������������̻.׻?N�kh�cU��m���S��	�o��	-����b �2L��#�&�'��+���/��3�ŗ7�
k;��/?���B�q�F��-J���M�_DQ��T��/X�g�[���^�`Hb�z�e���h�Ll��Jo�}yr�ơu��x���{���~����������;������򒈼I������a��C������Tm���Ⓖ�V���ɕ�<��T����������t����j���؟�0F��&������F���p����d��oЩ�_<��&���������밼�W���ó��/��/�������u���⺼3P������  �  ��N=�M=_<M=X�L=��K=<K=ZJ=��I=��H=_,H=�qG=Y�F=��E=f>E=��D=N�C=bC=�GB=��A=��@=�@=!F?=��>=/�==��<=16<=�o;=��:=��9=Q9=�H8=w{7=ڬ6=��5=�
5=974=�a3=��2=.�1=��0=��/=�/=55.=�O-=�g,=�|+=��*=͝)=F�(=M�'=��&=U�%=�$=��#=$�"=.�!=�{ =�b=�D=�!=l�=�=+�=�`=�"=��=a�=�E=i�=��=�3=@�=�^=��
=�r	=%�=�o=��=�V=6�=�( =��<���<�|�<�#�<���<�W�<d��<�k�<���<�b�<���<C@�<��<o�<�a�<L��<e
�<]X�<���<�<T,�<�l�<쩮<��<�<OS�<���<	��<��<w�<�H�<2v�<Ţ�<�΄<m��<�Kz<��r<��j<�Qc<�[<kT<�aL<?�D<S!=<5�5<T�-<�V&<��<�8<��<�-<h� <�r�;���;���;���;CJ�;b��;g�;o��;Fyz;��];�mA;�0%;�'	;���:�v�:[sY:���9nw�6�ҹ�dR�zP��Z�к�����3��`L��d��^|��뉻�z���۠����z������ɍ̻%׻N�yh�TU������S�	����8-����z �[L�.�#�i�'���+���/�Z�3��7�Dk;�0?��B���F��-J���M�JDQ��T��/X�:�[���^�/Hb�Q�e�t�h�#l��Jo�Zyr���u���x�y�{���~�	��⋂����5������񒈼F�����m��Y������om���Ⓖ�V��ʕ�1<��y���������������j���؟�7F��8������E���q����d��kЩ�J<������������밼|W���ó��/��������vu���⺼P�������  �  ��N=P�M=�5M=�|L=��K=
K=PJ=��I=��H=�H=�cG=��F=��E=�-E=�oD=[�C=M�B=�2B=rA=Ű@=��?=�+?=�g>=�==��<=<=�M;=v�:=Թ9=��8=u 8=�Q7=,�6=,�5=t�4=�4=�.3=YU2=�y1=k�0=��/=I�.=��-=-=�#,=�6+=sF*=S)=^\(=8b'=sd&=�b%=�]$=+T#=�F"=�4!=a =R=��=�=r�=�f=�2=!�=-�=�u=�+=��=�=�*=��=�b="�=��
=�	=^�=s=&�=��=�b=���<�]�<!�<���<]{�<��<���<�L�<���<]�<��<eR�<���<W/�<c��<���<�R�<���<&��<�M�<���<��<a(�<k�<,��<��<8$�<�]�<Y��<o˗< �<�3�<�e�<���<�Ȅ<:��<�Sz<1�r<�k<Wwc<��[<�>T<C�L<�E<�x=<��5<�W.<��&<�E<�<SE<��<eZ<���;��;�S�;Y��;�	�;y~�;��;á�;c�~;�2b;��E;�);��;1��:�ŭ:{�n:��:K/�8�����:�<���ĺ)2��ޣ�Q]-��E�I�]���u����,���b��`���Ǒ��e��ɻ�ӻ?�ݻB��u�񻨦�����qX�W��\�����i�����!�+&�H*�|S.��N2�H:6��:���=� �A�.XE�u�H�ƘL�i'P���S��$W�v�Z���]��Wa���d���g��=k�2{n�űq���t��x��/{��M~������=���Ń��K��|φ��Q���щ�^P��X͌��H��Ï��;������3*�������������@���l��)ݜ��M�������,��Л��\
���x���榼PT��©��/�����q
���w��e尼�R������:.��D���^
���x���纼�V��Jƽ��  �  ��N=L�M=�5M=�|L=��K=
K=PJ=��I=��H=�H=�cG=��F=��E=�-E=�oD=`�C=P�B=�2B=rA=��@=��?=�+?=�g>=��==�<=�<=�M;=m�:=˹9=��8=j 8=�Q7=.�6=*�5=w�4= 4=�.3=WU2=�y1=b�0=��/=E�.=v�-=-=�#,=�6+=|F*=S)=e\(=;b'=qd&=�b%=�]$=/T#=�F"=�4!=Q =]=��=
�=k�=�f=�2=%�=7�=�u=�+=��=�=�*=��=�b=�=Ń
=�	=_�=t=)�=��=�b=���<�]�<,�<���<I{�<|�<���<�L�<���<1]�<��<qR�<���<N/�<n��<���<�R�<���<��<�M�<���<��<R(�<k�<0��<��<Q$�<�]�<V��<S˗<���<r3�<�e�<���<�Ȅ<J��<�Sz<D�r<�k<hwc<��[<�>T<?�L<�E<�x=<��5<�W.<��&<�E<5�<�E<�<fZ<���;��;�S�;w��;�	�;�~�;E�;硍;��~;3b;��E;��);��;V��:�ƭ:��n:�:}%�8�����:�{=��_�ĺv3����� ]-��E��]�i�u����9���b����������e��_ɻ�ӻ��ݻ9��*��C���{��gX�\��������i����&�!�Q+&��G*�pS.��N2�f:6��:���=��A�XE�R�H���L��'P���S�%W���Z���]��Wa�~�d���g��=k�({n���q���t��x��/{��M~������=���Ń��K���φ�|Q���щ�KP��U͌��H��$Ï�<������0*������!������.���l��$ݜ��M��z����,������D
���x���榼lT��
©��/�����y
���w��U尼�R������<.��;���^
���x���纼�V��Dƽ��  �  ��N=V�M=�5M=�|L=��K=
K=PJ=��I=��H=�H=�cG=��F=��E=�-E=�oD=u�C=U�B=�2B=rA=ɰ@=��?=�+?=�g>=�==�<=�<=�M;=s�:=¹9=��8=\ 8=�Q7=�6=�5=m�4=�4=�.3=BU2=�y1=T�0=��/==�.=s�-=-=�#,=�6+=sF*=S)=c\(=Ab'=�d&=�b%=�]$=1T#=�F"=�4!=a =q=��=�=t�=�f=�2=#�=3�=�u=�+=��= �=�*=��=�b=�=��
=�	=S�=`=�=��=�b=���<x]�<&�<���<J{�<��<���<�L�<���<.]�<��<�R�<���<c/�<���<���<�R�<���<E��<�M�<	��<��<`(�<,k�<7��<��<F$�<�]�<_��<\˗< �<d3�<�e�<~��<�Ȅ<2��<1Sz<$�r<Gk<Dwc<8�[<�>T<�L<�E<�x=<��5<X.<��&<�E<�<`E<
�<jZ<Q��;��;;T�;���;
�;0�;��;���;�~;4b;�E;��);��;���:Cǭ:ǲn:��:p)�8����:�b>��4�ĺ�4�����^-���E���]�f�u��������b���������Ye��qɻ��ӻ��ݻ��g��e���~��KX� ��]��>��i�x����!�+&��G*�kS.��N2�;:6��:���=��A�XE�u�H���L��'P�O�S�%W���Z���]�Xa���d�3�g��=k�n{n��q���t��x��/{�8N~������=���Ń��K���φ�Q���щ�KP��S͌��H��Ï��;������+*������ ��y�������k��ݜ��M��]����,������Q
���x���榼dT�������/������
���w��m尼�R������a.��K����
���x���纼�V��Jƽ��  �  ��N=E�M=�5M=�|L=��K=
K=PJ=��I=��H=�H=�cG=ŧF=�E=�-E=�oD={�C=f�B=�2B=rA=հ@=��?=�+?=�g>=�==�<=�<=�M;=i�:=��9=��8=W 8=|Q7=�6=�5=_�4=�4=�.3=6U2=�y1=M�0=u�/=5�.=n�-=�-=�#,=�6+=vF*="S)=m\(=Gb'=�d&=	c%=�]$=AT#=�F"=�4!=o =s=��=$�=�=�f=�2=+�=>�=�u=�+=��=�=�*=��=�b=��=��
=�	=E�=O=�=��=�b=i��<f]�<�<{��<1{�<]�<}��<�L�<���<A]�<��<�R�<���<w/�<���<���<�R�<Ī�<Y��<N�<,��<��<|(�<5k�<I��<��<[$�<�]�<]��<O˗<���<Z3�<�e�<m��<zȄ<��<�Rz<�r<k<wc<�[<~>T<�L<gE<~x=<k�5<�W.<��&<�E<&�<�E<6�<�Z<k��;)�;�T�;D��;�
�;~�;b�;ࢍ;<�~;�4b;J�E;~�);�;h��:ɭ:��n:5�:0�8�����:�?����ĺR5��u���^-�@�E�^�]�(�u�/���(��c��6�������e���ɻU�ӻ��ݻ��E������U��/X� ��)���]i�e����!��*&�G*�&S.�eN2�	:6��:���=��A��WE�h�H���L��'P���S�"%W�ɔZ���]�'Xa�Ĭd�g�g�>k��{n�%�q��t��x��/{�MN~�ɳ��>���Ń��K���φ�{Q���щ�4P��=͌��H�����;��~���*��|������e�������k���ܜ�qM��U����,������<
���x���榼rT��©��/��$����
��x���尼S������z.��f����
��y���纼�V��cƽ��  �  ��N==�M=�5M=�|L=��K=
K=PJ=ŕI=��H=�H=dG=ڧF=&�E=�-E=pD=��C=��B=�2B=.rA=�@=��?=�+?=�g>=��==�<=�<=�M;=a�:=��9=��8=D 8=dQ7=�6=��5=C�4=�4=p.3=&U2=�y1=;�0=d�/='�.=h�-=�-=�#,=�6+=}F*=#S)=q\(=Qb'=�d&=c%=�]$=_T#=�F"=�4!=� =�=��=,�=��=�f=�2=/�=<�=�u=�+=��=��=�*=t�=�b=��=��
=�	=#�=3=�=b�=�b=.��<9]�<��<a��<{�<U�<y��<�L�<���<7]�<#��<�R�<��<�/�<���<���<S�<��<���<FN�<_��<�<�(�<Qk�<_��<��<e$�<�]�<W��<U˗<���<S3�<�e�<G��<MȄ<���<�Rz<r�r<�k<�vc<��[<@>T<��L<E<3x=<U�5<�W.<��&<�E<.�<�E<2�<�Z<���;��;�T�;���;v�;-��;=�;���;2�~;6b;~�E;&�); ;	��:oɭ:��n:��:99�8r�����:�`?��"�ĺ17�����v_-���E���]�W�u��������c�����������e���ɻr�ӻ��ݻ2�������?��X����Ո����h���L�!�q*&�"G*��R.�>N2��96�W:�~�=�ϤA��WE�K�H���L��'P���S�>%W���Z�4�]�lXa��d���g��>k� |n���q��t�6x�30{��N~�賀�>���Ń��K���φ��Q���щ�7P��.͌��H�����;��g����)��U������<��������k���ܜ�AM��;����,������5
���x���榼mT��)©��/��D����
��3x���尼9S�������.�������
��$y���纼W���ƽ��  �  p�N=8�M=�5M=�|L=��K=
K=)PJ=ՕI=�H=�H= dG=�F=5�E=�-E="pD=��C=��B=�2B=GrA=��@=��?=�+?=�g>=�==�<=�<=�M;=V�:=��9=��8=4 8=QQ7=�6=�5=1�4=�4=].3=U2=�y1=#�0=\�/=�.=W�-=�-=�#,=�6+=�F*=&S)=�\(=ab'=�d&=0c%=�]$=kT#=�F"=�4!=� =�=��=D�=��=�f=�2=;�=?�=�u=+=��=��=�*=`�=}b=��=w�
=�	=
�==ς=G�=�b=���<	]�<��<2��<�z�<H�<\��<�L�<���<F]�<<��<�R�<��<�/�<��<���<IS�<!��<���<iN�<~��<4�<�(�<uk�<���<�<p$�<�]�<O��<G˗<���<.3�<�e�<2��<Ȅ<���<NRz<!�r<Nk<?vc<E�[<�=T<-�L<�E<x=<�5<zW.<��&<�E<4�<�E<f�<�Z<a��;d�;�U�;���;�;)��;	�;���;I�~;�7b;H�E;�);|;���:b˭:c�n:��:�/�8����z�:�6A��v�ĺ�8������`-���E���]���u�����1	��Nd��f�������Hf��/ɻf�ӻ��ݻ/�������������W����������h������!�*&��F*�nR.��M2�l96�:�<�=���A��WE�&�H���L��'P���S�%W�5�Z�R�]��Xa�u�d���g��>k�W|n�ݲq���t��x�~0{��N~�����9>��ƃ��K���φ��Q���щ�"P��͌��H�����;��5����)����������������k���ܜ�$M������,������,
��~x���榼}T��/©��/��[����
��`x���尼jS������.��Ŝ���
��Vy��躼W���ƽ��  �  d�N=/�M=�5M=�|L=��K=
K=6PJ=ܕI=�H=�H=8dG=�F=R�E=.E=3pD=ɱC=��B=�2B=YrA=	�@=��?=�+?=�g>= �==
�<=�<=�M;=N�:=��9=��8= 8=@Q7=π6=ˮ5=�4=�4=F.3=�T2=�y1=�0=A�/=
�.=L�-=�-=�#,=�6+=�F*=0S)=�\(=jb'=�d&=<c%=�]$=�T#=�F"=5!=� =�=��=^�=��=�f=�2=B�=F�=�u=�+=��=�=~*=M�=^b=��=_�
=g	=�=�
=��=(�=�b=Е�<�\�<��<��<�z�<)�<S��<�L�<���<U]�<D��<�R�<7��<�/�<��<.��<�S�<B��<���<�N�<���<i�<�(�<�k�<���<-�<}$�<�]�<Y��<=˗<���<3�<ue�<���<�Ǆ<���<�Qz<��r<�k<�uc<��[<t=T<�L<rE<�w=<��5<QW.<`�&<�E<;�<�E<��<[<��;��;�V�;���;��;+��;�	�;���;>�~;�9b;��E;��);�;���:�ͭ:g�n:��:!=�8n���H�:�_B��щĺF;�����$b-�&�E�S�]�k�u�+����	���d��咨������f��vɻ��ӻ��ݻ������i���˟��W�-��O���Jh�+����!��)&�AF*�R.�eM2�496��:��=�i�A��WE�3�H���L��'P��S��%W�n�Z���]�Ya���d�h�g�.?k��|n�L�q�7�t� x��0{�=O~�%���T>��&ƃ��K���φ�vQ���щ�P��͌�vH����f;������~)��ߞ��_��͆��u���Uk��vܜ�M��򼟼t,��p���!
��{x���榼�T��C©��/��|������x��氼�S��;���/������ ���y��5躼KW���ƽ��  �  \�N="�M=�5M=�|L=��K=&
K=?PJ=�I=1�H=�H=IdG=�F=j�E=*.E=SpD=�C=��B=�2B=jrA=#�@=��?=�+?=�g>=�==�<=�<=�M;=C�:=��9=|�8= 8=%Q7=��6=��5=��4=�4=(.3=�T2=�y1=�0=.�/=��.=D�-=�-=�#,=�6+=�F*=:S)=�\(=vb'=�d&=Qc%=�]$=�T#=G"=)5!=� =�=�=n�=��=�f=�2=G�=N�=�u=w+=��=݅=q*=<�=Eb=��=>�
=I	=ɍ=�
=��=�=cb=���<�\�<S�<���<�z�<�<K��<�L�<���<d]�<U��<�R�<h��<�/�<?��<c��<�S�<���<&��<�N�<暹<��<)�<�k�<���<?�<�$�<�]�<O��<>˗<���<3�<Qe�<ږ�<�Ǆ<\��<tQz<>�r<{k<Zuc<g�[<�<T<{�L<%E<ew=<��5<W.<O�&<�E<-�<�E<��<Q[<���;��;0W�;P��;��;��;�
�;z��;"�~;i;b;�E;r�);;!��:|ϭ:۾n:��:D�8|�����:��B����ĺd<�����xc-���E���]�T�u�����
���e��I������g���ɻ�ӻ��ݻ�绷��������YW���������g�ʺ��!�?)&��E*��Q.�M2��86�c:���=�G�A�eWE�'�H�L��'P��S��%W���Z��]�MYa�0�d���g��?k�!}n���q���t�`x�51{�mO~�M���e>��;ƃ��K���φ��Q���щ��O���̌�VH��^�C;��ղ��G)������������D���#k��Sܜ��L��Ǽ��Y,��a���
���x���榼�T��^©� 0������)���x��:氼�S��z���9/��0���W���y��c躼mW���ƽ��  �  M�N=�M=�5M=�|L=��K=+
K=FPJ=��I=9�H= H=]dG=7�F=��E==.E=lpD=�C=��B=3B=�rA=+�@=�?=�+?=�g>=�==	�<=�<=�M;=3�:=|�9=l�8=  8=Q7=��6=��5=��4=j4=.3=�T2=fy1=�0="�/=��.=4�-=�-=�#,=�6+=�F*=;S)=�\(=�b'=�d&=dc%=^$=�T#=!G"=<5!=� =�=)�=��=ӕ=�f=�2=T�=K�=�u=s+=��=҅=]*='�=3b=��=�
=6	=��=�
=o�=��=Qb=M��<}\�<)�<���<�z�<��<7��<�L�<���<_]�<t��<�R�<s��<)0�<o��<���<�S�<���<J��<O�<��<��<<)�<�k�<֫�<T�<�$�<�]�<O��<2˗<���<�2�<.e�<Ö�<�Ǆ<,��<6Qz<Ǳr<k<�tc<#�[<�<T<�L<�E<w=<b�5<�V.<7�&<}E<H�<�E<��<�[<���;,�;�W�;#��;��;���;��;-��;կ~;M=b;��E;?�););��:BЭ:�n:��:	C�8������:�>D��X�ĺ�=��\��#d-���E�\�]���u�܃����\f������\����g��ɻ8�ӻ��ݻ��X������m��W�������p�{g�r����!��(&��E*�GQ.��L2��86�F:���=��A�eWE���H���L��'P�*�S�&W��Z�>�]��Ya���d���g�@k�}n��q� �t��x��1{��O~�m����>��\ƃ��K���φ�|Q���щ��O���̌�=H��O�;������)���������u�������j��,ܜ��L������3,��M���

��nx���榼�T��s©�0������?���x��i氼�S������f/��j���v���y���躼�W��ǽ��  �  D�N=�M=�5M=�|L=��K=*
K=MPJ= �I=J�H= H=tdG=D�F=��E=Z.E=�pD=�C=��B= 3B=�rA=>�@=�?=,?=h>=�==�<=�<=�M;=1�:=r�9=^�8=�8=Q7=��6=��5=��4=T4=�-3=�T2=\y1=ٛ0=�/=��.=-�-=�-=�#,=�6+=�F*=;S)=�\(=�b'=�d&=vc%=%^$=�T#=;G"=U5!=� = =7�=��=�=g=�2=Y�=K�=�u=v+=y�=υ=S*=�=b=n�=�
=	=��=�
=T�=��=/b=1��<J\�<�<���<�z�<��<#��<�L�<���<d]�<y��<S�<���<L0�<���<���<T�<۫�<���<6O�<3��<��<c)�<�k�<㫪<e�<�$�<�]�<S��<$˗<���<�2�<e�<���<�Ǆ<��<�Pz<w�r<�k<�tc<��[<S<T<آL<�E<�v=<6�5<�V.<�&<sE<M�<�E<��<�[<z��;��;�X�;���;e�;���;m�;3��;�~;q>b;P�E;��);d;���:�ѭ:_�n:��:]@�8I�����:�E����ĺc@�����e-�;�E���]��u�h�������f��o���ꔳ��g��Eɻ"�ӻ2�ݻ���k�����O���V�e��V���=g���T�!��(&�E*�Q.�eL2�B86�:�f�=��A�\WE��H���L�(P�*�S�&W�
�Z���]��Ya���d�|�g�i@k��}n�p�q�e�t�	x��1{�
P~������>��dƃ� L���φ�pQ���щ��O���̌�!H��+��:�������(��P������=��������j���ۜ��L������),��=���	
��nx���榼�T��p©�10��ٝ��m���x���氼%T�������/���������z���躼�W��ǽ��  �  9�N=�M=�5M=�|L=��K=6
K=\PJ=�I=V�H=! H=dG=T�F=��E=g.E=�pD=�C=��B=.3B=�rA=H�@=�?=,?=h>=�==�<=�<=�M;=(�:=j�9=Y�8=�8=�P7=}�6=y�5=��4=C4=�-3=�T2=Py1=Λ0=�/=��.="�-=�-=�#,=�6+=�F*=PS)=�\(=�b'=�d&=zc%=3^$=�T#=CG"=b5!= =	=D�=��=�=g=�2=^�=`�=�u=s+=s�=��=F*=�=b=_�=�
=�
	=��=�
=E�=��=b=��<*\�<��<���<lz�<��<��<�L�<���<�]�<���<$S�<���<Z0�<���<���<*T�<���<���<JO�<Q��<�<n)�<l�<�<~�<�$�<�]�<N��<˗<���<�2�<e�<y��<nǄ<���<�Pz<Y�r<ck<ntc<q�[<<T<��L<PE<�v=<�5<�V.<��&<dE<Q�<F<6�<�[<���;	�;Y�;)��;��;)��;��;���;��~;x?b;��E;l�);8;���:~ԭ:E�n:��:�>�8c���b�:��E���ĺ�A��P���f-���E� �]��u�x���i���f������C����g���ɻ}�ӻU�ݻ���a��@���*���V�*��?��� �g�޹��!�P(&��D*��P.�,L2�+86��:�G�=�УA� WE�	�H���L�(P�]�S�E&W��Z���]�Za��d���g�t@k�~n���q�z�t�Mx��1{�?P~������>��wƃ�L���φ�nQ���щ��O���̌�H����:��e����(��7������!��������j���ۜ��L��~���,��%����	��nx���榼�T���©�H0��۝�����
y���氼FT�������/���������'z���躼�W��ǽ��  �  8�N=�M=�5M=�|L=��K=0
K=SPJ=�I=Y�H=- H=�dG=b�F=��E=p.E=�pD=%�C=�B=93B=�rA=N�@=$�?=,?=h>=�==�<=�<=�M;=(�:=f�9=K�8=�8=�P7=y�6=n�5=��4=24=�-3=�T2=@y1=0=��/=��.=!�-=�-=�#,=�6+=�F*=ES)=�\(=�b'=�d&=�c%=6^$=�T#=OG"=p5!= ==U�=��=��=g=�2=^�=R�=�u=n+={�=��=E*=�=b=R�=��
=�
	=r�={
=0�=��=b=��<\�<��<���<kz�<��<%��<�L�<���<s]�<���<2S�<���<t0�<���<���<9T�<��<���<eO�<q��<�<�)�<l�<��<p�<�$�<�]�<W��<'˗<���<�2�<�d�<j��<SǄ<���<kPz<�r<+k<tc<T�[<�;T<s�L<7E<�v=<�5<�V.<�&<wE<E�<�E<�<�[<���;l�;KY�;���;P�;u��;��;���;b�~;E@b;��E;��);�;���:Eӭ:��n:?�:7O�8������:�F����ĺ�B��E���f-�G�E�M�]��u�%���s��pg���������:h���ɻu�ӻ�ݻ���O�񻏤��-���V�$�� ��� ��f������!�(&��D*��P.�L2��76��:� �=�ʣA�3WE��H���L��'P�U�S�C&W�B�Z���]�FZa�-�d���g��@k�^~n��q���t�Wx�02{�`P~������>��tƃ�L���φ�yQ���щ��O���̌� H����:��U����(��'��������������j���ۜ�pL��|���,��5����	��ox���榼�T���©�G0��󝬼���%y���氼PT��³��/��ȝ�����7z���躼�W��9ǽ��  �  7�N= �M=�5M=�|L=��K=:
K=YPJ=�I=V�H=5 H=�dG=]�F=��E=l.E=�pD=�C=�B=03B=�rA=P�@=$�?=,?=h>=�==�<=�<=�M;=�:=d�9=G�8=�8=�P7=u�6=c�5=��4=E4=�-3=�T2=;y1=ț0=��/=��.=�-=�-=�#,=�6+=�F*=FS)=�\(=�b'=�d&=�c%=1^$=�T#=OG"=m5!= ==V�=��=�=g=�2=h�=Q�=�u=k+=q�=��=A*=�=b=X�=�
=�
	=g�=�
=;�=��=b=��<)\�<��<���<[z�<��<��<�L�<���<v]�<���<7S�<���<�0�<���<���</T�<��<���<gO�<j��<�<�)�<l�<��<�<�$�<�]�<D��<˗<q��<�2�<�d�<t��<TǄ<���<YPz<�r<vk<tc<;�[<�;T<l�L<PE<�v=< �5<~V.<��&<WE<T�<&F<)�<\<���;��;IY�;x��;X�;X��;��;Ϩ�;a�~;�?b;#�E;�);�;5��:�ӭ:��n:��:�>�8����S�:�MF���ĺkA��m��g-���E���]���u�\���z���g��씨�f���lh���ɻ��ӻQ�ݻ���񻄤�����V�@��ӆ�� ��f������!�(&��D*��P.�4L2��76��:��=���A�5WE���H�ŘL�(P�~�S�R&W�S�Z���]�,Za�D�d���g��@k�~n���q���t�gx�=2{�7P~������>���ƃ�&L���φ�yQ��cщ��O���̌��G����:��c����(��1��������������j���ۜ�ZL�������+��%����	��fx���榼�T���©�I0��������#y���氼YT��³��/��̝�����?z���躼�W��Fǽ��  �  8�N=�M=�5M=�|L=��K=0
K=SPJ=�I=Y�H=- H=�dG=b�F=��E=p.E=�pD=%�C=�B=93B=�rA=N�@=$�?=,?=h>=�==�<=�<=�M;=(�:=f�9=K�8=�8=�P7=y�6=n�5=��4=24=�-3=�T2=@y1=0=��/=��.=!�-=�-=�#,=�6+=�F*=ES)=�\(=�b'=�d&=�c%=6^$=�T#=OG"=p5!= ==U�=��=��=g=�2=^�=R�=�u=o+={�=��=E*=�=b=S�=�
=�
	=r�=|
=1�=��=b=��<\�<��<���<mz�<��<&��<�L�<���<t]�<���<3S�<���<u0�<���<���<:T�<��<���<eO�<q��<�<�)�<l�<��<o�<�$�<�]�<V��<&˗<���<�2�<�d�<j��<SǄ<���<jPz<�r<+k<tc<T�[<�;T<t�L<8E<�v=<�5<�V.<�&<yE<G�<�E<�<�[<���;o�;MY�;���;Q�;v��;��;���;^�~;@@b;��E;��);�;��:1ӭ:��n:�:�M�8����*�:�&F����ĺ�B��P���f-�R�E�W�]��u�)���w��sg���������=h���ɻx�ӻ�ݻ���P�񻑤��.���V�%�� ��� ��f������!�(&��D*��P.�L2��76��:� �=�ʣA�3WE��H���L��'P�U�S�C&W�B�Z���]�FZa�-�d���g��@k�^~n��q���t�Wx�02{�`P~������>��tƃ�L���φ�yQ���щ��O���̌� H����:��U����(��'��������������j���ۜ�pL��|���,��5����	��ox���榼�T���©�G0��󝬼���%y���氼PT��³��/��ȝ�����7z���躼�W��9ǽ��  �  9�N=�M=�5M=�|L=��K=6
K=\PJ=�I=V�H=! H=dG=T�F=��E=g.E=�pD=�C=��B=.3B=�rA=H�@=�?=,?=h>=�==�<=�<=�M;=(�:=j�9=Y�8=�8=�P7=}�6=y�5=��4=C4=�-3=�T2=Py1=Λ0=�/=��.="�-=�-=�#,=�6+=�F*=PS)=�\(=�b'=�d&=zc%=3^$=�T#=CG"=b5!= =	=D�=��=�=g=�2=^�=`�=�u=t+=s�=��=G*=�=b=`�=�
=�
	=��=�
=F�=��=b=��<,\�<��<���<oz�<��<��<�L�<���<�]�<���<&S�<���<[0�<���<���<*T�<���<���<JO�<Q��< �<m)�<l�<�<|�<�$�<�]�<L��<˗<���<�2�<e�<x��<mǄ<���<�Pz<X�r<ck<otc<r�[<<T<��L<SE<�v=<	�5<�V.<��&<hE<T�<F<:�<�[<���;�;
Y�;,��;��;)��;��;���;��~;o?b;��E;^�);(;ַ�:Xԭ:��n:��:�;�8�����:��E���ĺ�A��f���f-���E�4�]��u�����p���f��ǔ��I����g���ɻ��ӻY�ݻ���d��B���+���V�+��@��� �g�߹��!�P(&��D*��P.�,L2�,86��:�G�=�УA� WE�	�H���L�(P�]�S�E&W��Z���]�Za��d���g�t@k�~n���q�z�t�Mx��1{�?P~������>��wƃ�L���φ�nQ���щ��O���̌�H����:��e����(��7������!��������j���ۜ��L��~���,��%����	��nx���榼�T���©�H0��۝�����
y���氼FT�������/���������'z���躼�W��ǽ��  �  D�N=�M=�5M=�|L=��K=*
K=MPJ= �I=J�H= H=tdG=D�F=��E=Z.E=�pD=�C=��B= 3B=�rA=>�@=�?=,?=h>=�==�<=�<=�M;=1�:=r�9=^�8=�8=Q7=��6=��5=��4=T4=�-3=�T2=\y1=ٛ0=�/=��.=-�-=�-=�#,=�6+=�F*=;S)=�\(=�b'=�d&=vc%=&^$=�T#=;G"=U5!=� = =7�=��=�=g=�2=Y�=K�=�u=w+=y�=υ=T*=�= b=o�=�
=	=��=�
=V�=��=1b=4��<M\�<�<���<�z�<��<'��<�L�<���<g]�<|��<S�<���<N0�<���<���<T�<۫�<���<6O�<2��<��<b)�<�k�<᫪<c�<�$�<�]�<Q��<"˗<���<�2�<e�<���<�Ǆ<	��<�Pz<w�r<�k<�tc<��[<V<T<ۢL<�E<�v=<:�5<�V.<�&<xE<S�<�E<��<�[<���;��;�X�;���;g�;���;l�;0��;��~;d>b;@�E;��);N;˶�:Pѭ:��n:m�:e<�8N����:�VE����ĺ�@������e-�W�E���]��u�t�������f��x���򔳻�g��Lɻ(�ӻ7�ݻ���o�����P���V�g��W���>g���U�!��(&�E*�Q.�eL2�B86�:�f�=��A�\WE��H���L�(P�*�S�&W�
�Z���]��Ya���d�|�g�i@k��}n�p�q�e�t�	x��1{�
P~������>��dƃ� L���φ�pQ���щ��O���̌�!H��+��:�������(��P������=��������j���ۜ��L������),��=���	
��nx���榼�T��p©�10��ٝ��m���x���氼%T�������/���������z���躼�W��ǽ��  �  M�N=�M=�5M=�|L=��K=+
K=FPJ=��I=9�H= H=]dG=7�F=��E==.E=lpD=�C=��B=3B=�rA=+�@=�?=�+?=�g>=�==	�<=�<=�M;=3�:=|�9=l�8=  8=Q7=��6=��5=��4=j4=.3=�T2=fy1=�0="�/=��.=4�-=�-=�#,=�6+=�F*=;S)=�\(=�b'=�d&=dc%=^$=�T#=!G"=<5!=� =�=)�=��=ԕ=�f=�2=U�=K�=�u=t+=��=Ӆ=^*=(�=4b=��=!�
=8	=��=�
=q�=��=Sb=R��<�\�<-�<���<�z�<�<;��<�L�<���<b]�<w��< S�<u��<+0�<q��<���<�S�<���<J��<O�<��<��<:)�<�k�<ԫ�<R�<�$�<�]�<L��</˗<���<�2�<,e�<���<�Ǆ<+��<4Qz<Ʊr<k<�tc<%�[<�<T<�L<�E<w=<h�5<�V.<>�&<�E<N�<�E<��<�[<���;4�;�W�;'��;��;���;��;*��;ɯ~;<=b;��E;'�);;ʵ�:�ϭ:�n:'�:*>�8������:��D����ĺ$>�����Hd-���E�~�]�şu�ꃆ���if�����f����g��!ɻ@�ӻ�ݻ��]������o��W�������q�|g�s����!��(&��E*�GQ.��L2��86�F:���=��A�eWE���H���L��'P�*�S�&W��Z�>�]��Ya���d���g�@k�}n��q� �t��x��1{��O~�m����>��\ƃ��K���φ�|Q���щ��O���̌�=H��O�;������)���������u�������j��,ܜ��L������3,��M���

��ox���榼�T��s©�0������?���x��i氼�S������f/��j���v���y���躼�W��ǽ��  �  \�N="�M=�5M=�|L=��K=&
K=?PJ=�I=1�H=�H=IdG=�F=j�E=*.E=SpD=�C=��B=�2B=jrA=#�@=��?=�+?=�g>=�==�<=�<=�M;=C�:=��9=|�8= 8=%Q7=��6=��5=��4=�4=(.3=�T2=�y1=�0=.�/=��.=D�-=�-=�#,=�6+=�F*=:S)=�\(=vb'=�d&=Qc%=�]$=�T#=G"=)5!=� =�=�=n�=��=�f=�2=H�=O�=�u=x+=��=ޅ=q*==�=Fb=��=?�
=K	=ˍ=�
=��=�=eb=���<�\�<X�<���<�z�<�<P��<�L�<���<h]�<Y��<�R�<k��<�/�<A��<d��<�S�<���<&��<�N�<嚹<��<)�<�k�<���<<�<�$�<�]�<L��<:˗<���<3�<Oe�<ؖ�<�Ǆ<[��<rQz<=�r<{k<[uc<i�[<=T<�L<*E<jw=<��5<W.<U�&<�E<4�<�E<��<W[<���;��;7W�;U��;��;��;�
�;v��;�~;W;b;��E;X�);�;ܲ�:2ϭ:;�n:�:�>�8������:�C���ĺ�<��$���c-���E���]�w�u�����
���e��U������)g���ɻ��ӻ��ݻ%�绽��������[W���������g�˺��!�@)&��E*��Q.�M2��86�d:���=�G�A�eWE�'�H�L��'P��S��%W���Z��]�MYa�0�d���g��?k�!}n���q���t�`x�51{�mO~�M���e>��;ƃ��K���φ��Q���щ��O���̌�VH��^�C;��ղ��G)������������D���#k��Sܜ��L��Ǽ��Y,��a���
���x���榼�T��^©� 0������)���x��:氼�S��z���9/��0���W���y��c躼mW���ƽ��  �  d�N=/�M=�5M=�|L=��K=
K=6PJ=ܕI=�H=�H=8dG=�F=R�E=.E=3pD=ɱC=��B=�2B=YrA=	�@=��?=�+?=�g>= �==
�<=�<=�M;=N�:=��9=��8= 8=@Q7=π6=ˮ5=�4=�4=F.3=�T2=�y1=�0=A�/=
�.=L�-=�-=�#,=�6+=�F*=0S)=�\(=jb'=�d&=<c%=�]$=�T#=�F"=5!=� =�=��=^�=��=�f=�2=B�=F�=�u=�+=��=�=*=N�=_b=��=a�
=i	=�=�
=��=+�=�b=Օ�<�\�<��<��<�z�</�<X��<�L�<���<Z]�<H��<�R�<:��<�/�<��<0��<�S�<B��<���<�N�<���<h�<�(�<�k�<���<*�<z$�<�]�<U��<:˗<���<3�<re�<���<�Ǆ<���<�Qz<��r<�k<�uc<��[<x=T<�L<wE<�w=<��5<WW.<g�&<�E<C�<�E<��<"[<��;��;�V�;���; �;,��;�	�;���;0�~;�9b;��E;t�);�;���:Kͭ:»n:��:7�8�����:��B��-�ĺ�;�����Nb-�N�E�y�]���u�<���
���d��򒨻�����f���ɻ��ӻ��ݻ������n���͟��W�/��P���Kh�,����!��)&�AF*�R.�eM2�496��:��=�i�A��WE�3�H���L��'P��S��%W�n�Z���]�Ya���d�h�g�.?k��|n�L�q�7�t� x��0{�=O~�%���T>��&ƃ��K���φ�vQ���щ�P��͌�vH����f;������~)��ߞ��_��̆��u���Uk��vܜ�M��򼟼t,��p���!
��{x���榼�T��C©��/��|������x��氼�S��;���/������ ���y��5躼KW���ƽ��  �  p�N=8�M=�5M=�|L=��K=
K=)PJ=ՕI=�H=�H= dG=�F=5�E=�-E="pD=��C=��B=�2B=GrA=��@=��?=�+?=�g>=�==�<=�<=�M;=V�:=��9=��8=4 8=QQ7=�6=�5=1�4=�4=].3=U2=�y1=#�0=\�/=�.=W�-=�-=�#,=�6+=�F*=&S)=�\(=ab'=�d&=0c%=�]$=kT#=�F"=�4!=� =�=��=D�=��=�f=�2=<�=?�=�u=+=��=��=�*=a�=~b=��=y�
=�	=�==т=I�=�b=��<]�<��<7��<�z�<M�<a��<�L�<���<J]�<@��<�R�<��<�/�<��<���<JS�<!��<���<iN�<}��<2�<�(�<rk�<~��<�<l$�<�]�<K��<C˗<���<+3�<�e�<0��<Ȅ<���<LRz< �r<Nk<@vc<G�[<�=T<1�L<�E<x=<	�5<�W.<��&<�E<;�<�E<l�<[<k��;m�;�U�;���;	�;*��;	�;���;<�~;�7b;1�E;��);];B��:˭:ĺn:2�:6*�8����.�:��A��χĺ9��ݦ��`-���E��]���u�����@	��\d��s���͒��Rf��8ɻn�ӻ��ݻ6�����ť������W����������h������!�*&��F*�oR.��M2�l96�:�<�=���A��WE�&�H���L��'P���S�%W�5�Z�R�]��Xa�u�d���g��>k�W|n�ݲq���t��x�~0{��N~�����9>��ƃ��K���φ��Q���щ�"P��͌��H�����;��5����)����������������k���ܜ�$M������,������,
��~x���榼}T��/©��/��[����
��`x���尼jS������.��Ŝ���
��Vy��躼W���ƽ��  �  ��N==�M=�5M=�|L=��K=
K=PJ=ŕI=��H=�H=dG=ڧF=&�E=�-E=pD=��C=��B=�2B=.rA=�@=��?=�+?=�g>=��==�<=�<=�M;=a�:=��9=��8=D 8=dQ7=�6=��5=C�4=�4=p.3=&U2=�y1=;�0=d�/='�.=h�-=�-=�#,=�6+=}F*=#S)=q\(=Qb'=�d&=c%=�]$=_T#=�F"=�4!=� =�=��=,�=��=�f=�2=/�==�=�u=�+=��= �=�*=u�=�b=��=��
=�	=%�=5=�=d�=�b=2��<=]�<��<e��<{�<Y�<~��<�L�<���<;]�<&��<�R�<��<�/�<���<���<S�<��<���<EN�<^��<��<�(�<Ok�<\��<��<b$�<�]�<T��<R˗<���<Q3�<�e�<E��<KȄ<���<�Rz<q�r<�k<�vc<��[<C>T<��L<E<8x=<[�5<�W.<��&<�E<4�<�E<8�<�Z<���;��;�T�;���;x�;-��;<�;���;&�~;6b;i�E;�);  ;ˬ�:,ɭ:�n:�:\4�8����^�:��?��r�ĺ7�����_-���E��]�v�u��������c��ő�������e���ɻy�ӻ��ݻ8�������A��X����ֈ����h���M�!�q*&�#G*��R.�>N2��96�W:�~�=�ФA��WE�K�H���L��'P���S�>%W���Z�4�]�lXa��d���g��>k� |n���q��t�6x�30{��N~�賀�>���Ń��K���φ��Q���щ�7P��.͌��H�����;��g����)��U������<��������k���ܜ�AM��;����,������5
���x���榼mT��)©��/��D����
��3x���尼9S�������.�������
��$y���纼W���ƽ��  �  ��N=E�M=�5M=�|L=��K=
K=PJ=��I=��H=�H=�cG=ŧF=�E=�-E=�oD={�C=f�B=�2B=rA=հ@=��?=�+?=�g>=�==�<=�<=�M;=i�:=��9=��8=W 8=|Q7=�6=�5=_�4=�4=�.3=6U2=�y1=M�0=u�/=5�.=n�-=�-=�#,=�6+=vF*="S)=m\(=Gb'=�d&=	c%=�]$=AT#=�F"=�4!=o =s=��=$�=�=�f=�2=,�=>�=�u=�+=��=�=�*=��=�b=��=��
=�	=F�=P=�=��=�b=m��<j]�<�<~��<5{�<a�<���<�L�<���<D]�<��<�R�<���<y/�<���<���<�R�<Ū�<Y��<N�<+��<��<z(�<3k�<G��<��<Y$�<�]�<Z��<M˗<���<W3�<�e�<k��<xȄ<��<�Rz<�r<k<wc<�[<�>T<�L<kE<�x=<o�5<�W.<��&<�E<+�<�E<;�<�Z<s��;0�;�T�;H��;�
�;�;`�;ݢ�;2�~;�4b;9�E;j�);	�;6��:�ȭ:�n:��:,�8���i�:�P?���ĺ�5������^-�\�E�z�]�B�u�;���3��c��?��� ����e���ɻ[�ӻ��ݻ
��I������W��1X���*���^i�f����!��*&�G*�&S.�fN2�	:6��:���=��A��WE�h�H���L��'P���S�"%W�ɔZ���]�'Xa�Ĭd�g�g�>k��{n�%�q��t��x��/{�MN~�ɳ��>���Ń��K���φ�{Q���щ�4P��=͌��H�����;��~���*��|������e�������k���ܜ�qM��U����,������<
���x���榼rT��©��/��$����
��x���尼S������z.��f����
��y���纼�V��cƽ��  �  ��N=V�M=�5M=�|L=��K=
K=PJ=��I=��H=�H=�cG=��F=��E=�-E=�oD=u�C=U�B=�2B=rA=ɰ@=��?=�+?=�g>=�==�<=�<=�M;=s�:=¹9=��8=\ 8=�Q7=�6=�5=m�4=�4=�.3=BU2=�y1=T�0=��/==�.=s�-=-=�#,=�6+=sF*=S)=c\(=Ab'=�d&=�b%=�]$=1T#=�F"=�4!=a =q=��=�=t�=�f=�2=#�=3�=�u=�+=��=!�=�*=��=�b=�=��
=�	=T�=a=�=��=�b=���<{]�<)�<���<M{�<��<���<�L�<���<0]�<	��<�R�<���<e/�<���<���<�R�<���<D��<�M�<	��<��<_(�<*k�<5��<��<D$�<�]�<]��<Z˗< �<c3�<�e�<}��<�Ȅ<1��<0Sz<#�r<Gk<Ewc<9�[<�>T<�L<�E<�x=<��5<X.<��&<�E<�<cE<�<mZ<V��;��;>T�;���;
�;0�;��;���;�~;�3b;t�E;u�);��;���:ǭ:u�n:{�:�&�8>�B�:��>��b�ĺ5��ң�^-���E���]�x�u��������b�������^e��vɻ��ӻ��ݻ��j��g������LX�!��^��?��i�x����!�+&��G*�kS.��N2�;:6��:���=��A�XE�u�H���L��'P�O�S�%W���Z���]�Xa���d�3�g��=k�n{n��q���t��x��/{�8N~������=���Ń��K���φ�Q���щ�KP��S͌��H��Ï��;������+*������ ��y�������k��ݜ��M��]����,������Q
���x���榼dT�������/������
���w��m尼�R������a.��K����
���x���纼�V��Jƽ��  �  ��N=L�M=�5M=�|L=��K=
K=PJ=��I=��H=�H=�cG=��F=��E=�-E=�oD=`�C=P�B=�2B=rA=��@=��?=�+?=�g>=��==�<=�<=�M;=m�:=˹9=��8=j 8=�Q7=.�6=*�5=w�4= 4=�.3=WU2=�y1=b�0=��/=E�.=v�-=-=�#,=�6+=|F*=S)=e\(=;b'=qd&=�b%=�]$=/T#=�F"=�4!=Q =]=��=
�=k�=�f=�2=%�=7�=�u=�+=��=�=�*=��=�b=�=Ń
=�	=`�=u=)�=��=�b=���<�]�<-�<���<J{�<}�<���<�L�<���<2]�<	��<rR�<���<N/�<n��<���<�R�<���<��<�M�<���<��<Q(�<k�</��<��<P$�<�]�<U��<R˗<���<q3�<�e�<���<�Ȅ<I��<�Sz<D�r<�k<hwc<��[<�>T<@�L<�E<�x=<��5<�W.<��&<�E<6�<�E<
�<hZ<���;��;�S�;y��;�	�;�~�;D�;桍;��~;3b;��E;��);��;C��:�ƭ:~�n:��:$�8����N�:��=��w�ĺ�3�����+]-��E��]�r�u����=���b���������� e��aɻ�ӻ��ݻ;��,��D���|��gX�]��������i����&�!�Q+&��G*�pS.��N2�f:6��:���=��A�XE�R�H���L��'P���S�%W���Z���]��Wa�~�d���g��=k�({n���q���t��x��/{��M~������=���Ń��K���φ�|Q���щ�KP��U͌��H��$Ï�<������0*������!������.���l��$ݜ��M��z����,������D
���x���榼lT��
©��/�����y
���w��U尼�R������<.��;���^
���x���纼�V��Dƽ��  �  ˡN=��M=S/M=�uL=��K=K=7FJ=��I=L�H=-H=|VG=V�F=��E=TE=^D=�C=��B=�B=\A=��@=A�?=�?=�L>=��==6�<=��;=*-;=Db:=�9=w�8=��7=�(7=�V6=,�5=��4=]�3='�2=�!2=�D1=#e0=5�/=�.=$�-=��,=Z�+=�*=� *=O)=�(=Z'=�&=%=�$=g #=��!=9� =!�=o�=1�=a=6==��=n�=�V=�=��=�v=!=��=�d=^�=s�=� 
=��=�-=�=%=2�=I=���<��<�q�<�*�<���<Ƃ�<�"�<��<�K�<���<�X�<���<WL�<T��<�(�<k��<��<]N�<B��<J��<�M�<���<��<h.�<�s�<K��<���<J5�<�q�<���<}�<��<%V�<���<�<��<�Zz<A�r<0k<��c<x\<^vT<b�L<vXE<�=<�D6<��.<�>'<;�<�H<��<Mf	<��<_7�;ـ�;B��;�?�;���;!A�;�ݝ;���;#S�;[\f;�AJ;YW.;y�;>:�:z��:̓�:h�:"}59��o�u;$���������2�:��E('��x?��wW��#o�u=�����j=��<�������Ż�-лQ{ڻ8��L���a��������e
�	��y�R��3?�e� ��$�o�(���,���0�X�4�t�8�(�<�&p@��+D���G��}K�BO���R��#V���Y��
]��o`���c�� g��mj���m���p�
(t��Xw��z�:�}��d��'�N}��3������������P���	������ ����������v��햼�b���י�mK�������0��٢��������S���Ye��զ��D��鳩�#��8���7��%p��E߰�=N�������,��]������|��e캼#]��]ν��  �  ¡N=��M=F/M=�uL=��K=K=FFJ=�I=N�H=%H=~VG=V�F=��E=UE=p^D=�C=��B=�B=\A=��@=C�?=?=�L>=��==8�<=��;= -;=:b:=�9=��8=��7=�(7=�V6=%�5=��4=h�3='�2=�!2=�D1=e0=;�/=��.=�-=��,=I�+=�*=� *=Z)=�(=]'=�&=%=�$=c #=��!=1� =�=u�=-�=a=6=	=��=y�=�V=�=��=�v=!=��=�d=e�=e�=� 
=�=�-=��="%=-�=D=���<��<�q�<�*�<���<���<�"�<��<�K�<���<�X�<���<ML�<S��<�(�<k��<��<?N�<B��<W��<�M�<���<��<g.�<�s�<g��<���<O5�<�q�<ᬗ<p�<��<6V�<���<�<��<�Zz<H�r<E0k<��c<C\<YvT<T�L<nXE<*�=<�D6<��.<[>'<)�<�H<��<�f	<��<l7�;���;Q��;�?�;���;2A�;�ݝ;ύ�;1S�;�\f;�AJ;�V.;��;;�:$��:I��:�:;t59t�o��=$�N���ؾ��3���c('��x?�wW��"o�n=��B�������=���;�������Ż�-л�{ڻB��6��~a�������e
����x�`��?��� ��$�W�(���,�s�0�a�4�z�8��<��o@��+D���G�~K��O��R�$V���Y��
]��o`���c�� g��mj���m���p�(t�Yw��z�e�}��d��1�c}��E��������𔉼6��ᕌ������� ��	��������v��3햼�b���י�oK������1��ۢ����ᄢ�D���Ue��զ��D������ #��&���6��2p��C߰�VN�������,��W�����|��k캼&]��Hν��  �  ��N=��M=I/M=�uL=��K=K=BFJ= �I=X�H=)H=�VG=Z�F=��E=eE=z^D=��C=��B=�B=#\A=��@=K�?=�?=�L>=��==:�<=��;='-;=Ab:=�9=��8=r�7=�(7=�V6=�5=��4=R�3=!�2=�!2=�D1=
e0=:�/=�.=�-=��,=I�+=�*=� *=R)=�(=^'=�&=%=�$=a #=��!=@� =!�=��=*�=a=6==��=q�=�V=�=��=�v=!=��=�d=d�=U�=� 
=�=�-=�=%=#�=8=���<ʯ�<�q�<{*�<���<Â�<�"�<��<�K�<���<�X�<���<WL�<Z��<�(�<h��<2��<RN�<_��<i��<�M�<ț�<��<}.�<�s�<_��<���<I5�<�q�<欗<��<��<-V�<���<�<��<�Zz<*�r<�/k<��c<$\<MvT<0�L<CXE<�=<�D6<ʿ.<h>'<9�<�H<��<yf	<��<�7�;���;���;�?�;귺;�A�;�ݝ;c��;BS�;5]f;BJ;jW.;;�;�:�:ޥ�:b��:*�:rx59��o��;$��������5�E���('�[y?�RxW�)$o��=���������/>���;������Żv-л�{ڻ��o�a�������e
����x�f���>�D� �߻$��(���,�L�0�\�4�_�8��<�p@��+D���G��}K��O��R�!$V��Y��
]�p`���c�!g��mj��m���p�8(t�5Yw��z���}��d��A�W}��2�������� ���?��알�������������������lv�� 햼�b��vי�jK��}����0��Ƣ����ꄢ�W���\e��զ��D��ݳ��,#��0���D��Hp��D߰�fN�������,��i���'�� |��|캼:]��Nν��  �  ��N=��M=A/M=�uL=��K=K=LFJ=	�I=\�H=7H=�VG=h�F=��E=jE=�^D=��C=��B=�B=+\A=��@=P�?=?=�L>=��==9�<=��;=-;=9b:=�9=u�8=r�7=�(7=�V6=�5=��4=G�3=�2=�!2=�D1=e0=1�/=�.=�-=��,=E�+=�*=� *=c)=�(=f'=�&=%=�$=r #=��!=G� =,�=��=;�=&a=6==��=z�=�V=�=��=�v=� =��=�d=W�=Q�=� 
=ө=�-=٫=%=�='=���<Ư�<�q�<i*�<���<���<�"�<��<�K�<���<�X�<���<lL�<i��<)�<���<8��<pN�<i��<w��<�M�<؛�<��<�.�<�s�<v��<���<S5�<�q�<ڬ�<n�<��<V�<���<}<���<�Zz<�r<�/k<f�c<\<vT<�L<5XE<��=<�D6<��.<C>'<&�<�H<��<�f	<�<�7�;.��;���;U@�;?��;�A�;jޝ;���;�S�;^f;�BJ;dX.;��;a<�:���:n��:��:�y59�o� =$�G��������4����)'�yy?��xW��$o��=��þ��_��@>��+<��L���Ż�-л�{ڻ��/��-a����ǽ�be
�����x����>�$� ���$��(���,� �0�4�4�9�8��<��o@��+D���G��}K��O�#�R�$$V�D�Y��
]�p`���c�L!g��mj��m��p�G(t�mYw�R�z���}��d��M�d}��O��������蔉�#��ؕ��������������������ev��햼�b��gי�KK��o����0��������Ԅ��7���Re��զ��D������,#��I���M��Xp��i߰�qN������-��w���/��D|���캼?]��gν��  �  ��N=��M=G/M=�uL=��K=K=IFJ=�I=c�H=EH=�VG=x�F=��E=yE=�^D=�C=��B=�B=7\A=��@=W�?=?=�L>=��==2�<=��;=-;=4b:=��9=d�8=f�7=�(7=�V6=�5=��4=?�3=�2=�!2=~D1=�d0=#�/=ڞ.=�-=��,=N�+=�*=� *=[)=�(=p'=�&=-%=�$=� #=�!=X� ==�=��=Q�=,a=-6= =��=}�=�V=�=��=�v=� =��=�d=E�=C�=� 
=ĩ=j-=˫=�$=�==���<���<iq�<W*�<���<���<�"�<Һ�<�K�<���<�X�<���<�L�<���<)�<���<S��<�N�<���<���<N�<曵<��<�.�<�s�<u��<���<P5�<�q�<鬗<[�<��<�U�<���<f<���<>Zz<��r<�/k<�c<�\<�uT<��L<XE<��=<�D6<r�.<V>'<(�<yH<��<�f	<I�<$8�;���;4��;�@�;︺;mB�;ߝ;��;�T�;_f;�CJ;QY.;S�;?>�:8��:���:��:U�59 �o��=$����������5뺘��
*'��z?��yW�$%o�^>��(������>���<����� �Ż.л�{ڻ:��3��_a�������?e
����~x�����>�څ �f�$���(�I�,��0���4��8�Ʀ<��o@��+D���G�~K�jO�3�R�+$V�a�Y��
]�@p`��c�z!g�nj�3�m�F�p��(t��Yw���z�̩}��d��X�m}��Q��������ꔉ�2��Õ�����������΅������Jv���얼�b��@י�'K��a����0���������ք��>���We��զ��D�����0#��a���c��op��߰��N��ͽ��-������Y��X|���캼U]���ν��  �  ��N=��M=</M=�uL=��K=!K=PFJ= �I=o�H=NH=�VG=��F=��E=�E=�^D=#�C=��B=�B=K\A=Ù@=c�?=?=�L>=��==;�<=��;=-;=,b:=�9=\�8=V�7=�(7=�V6=�5=w�4=,�3=��2=�!2=rD1=�d0=�/=О.=�-=��,=A�+=�*=� *=`)=�(=z'=�&=;%=�$=� #=�!=h� =K�=��=Y�==a=<6='=��=��=�V=�=��=�v=� =��=�d=8�=*�=� 
=��=S-=��=�$=�==}��<|��<Rq�<5*�<���<~��<�"�<ۺ�<�K�<���<�X�<���<�L�<���<?)�<Ə�<}��<�N�<���<���<!N�<��<��<�.�<�s�<���<���<f5�<�q�<Ӭ�<U�<��<�U�<n��<=<���<�Yz<i�r<J/k<Śc<j\<�uT<|�L<�WE<~�=<>D6<Z�.<(>'<�<�H<��<�f	<r�<�8�;��;���;nA�;m��;C�;�ߝ;Ώ�;�T�;W`f;EJ;Z.;C�;�?�:P��:+��:��:q}59��o��>$�ḅ�¸��7뺆���*'��{?��zW�/&o��>��������?���<�����t�Ż5.л�{ڻ.��Ĕ�3a��n�p��e
�h��+x����@>��� �+�$��(�!�,���0���4���8���<��o@��+D���G��}K��O�P�R�e$V���Y�
]��p`�>�c��!g�jnj�z�m���p��(t��Yw�΄z��}��d��r򁼀}��d��"������֔��)���������k����������s���v���얼fb��"י�	K��6����0���������Ǆ��7���Be��!զ��D�����O#��u���|���p���߰��N���:-����|��q|���캼r]���ν��  �  ��N=��M=7/M=�uL=��K=#K=_FJ=%�I=~�H=]H=�VG=��F=��E=�E=�^D=9�C=��B=B=W\A=ԙ@=p�?=%?=�L>=��==:�<=��;=-;=(b:=�9=Q�8=F�7=�(7=�V6=��5=e�4=�3=��2=�!2=`D1=�d0=
�/=Ȟ.=��-=��,==�+=�*=� *=g)=�(=�'=�&=F%=�$=� #=2�!=|� =_�=��=f�=Pa=F6=6= �=��=�V=�=��=�v=� =��=�d=%�=�=� 
=��=@-=��=�$=ט=�=X��<W��</q�<*�<z��<s��<~"�<Ӻ�<�K�<���<	Y�<���<�L�<���<c)�<��<���<�N�<ܧ�<���<AN�<6��<��<�.�<�s�<���<��<b5�<�q�<ˬ�<P�<��<�U�<L��< <���<�Yz<%�r<�.k<�c<\<>uT<<�L<}WE<O�=<D6<I�.<>'<�<�H<�<�f	<��<9�;v��;m��;�A�;��;�C�;+��;���;�U�;�af;FJ;`[.;S�;>A�:���:l��:B�:��59��o��>$�t���ø�39�7��,'��|?��{W��'o�J?��E������w?��;=��	����ŻK.л
|ڻ��ߔ��`��7�M���d
�6���w�Z���=�?� �պ$�&�(���,�c�0���4���8�x�<�yo@�s+D���G��}K��O�Y�R�w$V���Y�E]��p`���c�"g��nj�ֳm���p�.)t�+Zw��z�N�}�e���򁼇}��h��!������ޔ�����������I����������V����u���얼8b���֙��J������0��t����������-���He�� զ��D�����^#����������p���߰��N�����p-��✶�����|���캼�]���ν��  �  ��N=��M=6/M=�uL=��K=)K=cFJ=.�I=��H=mH=�VG=��F=��E=�E=�^D=I�C=�B="B=d\A=�@=y�?=,?=�L>=��==9�<=��;=	-;=b:=�9=?�8=9�7=�(7=�V6=̂5=N�4= �3=��2=�!2=LD1=�d0=��/=��.=��-=u�,=A�+=�*=� *=i)=�(=�'=�&=S%=$=� #=A�!=�� =t�=ɨ=}�=^a=P6=C=�=��=�V=�=��=�v=� =��=�d=�=�={ 
=��=%-=��=�$=��=�=)��<6��<q�<*�<V��<^��<"�<ʺ�<�K�<���<Y�<���<�L�<н�<�)�<��<���<O�< ��<��<nN�<T��<�<�.�<t�<���<��<c5�<�q�<Ϭ�<1�<��<�U�<*��<<u��<YYz<��r<�.k<�c<�\<�tT<��L<:WE<�=<�C6<�.<>'<�<�H<�<�f	<��<[9�;���;���;�B�;���;�D�;�;,��;QV�;cf;GJ;�\.;�;�B�:���:j��:�:}�59��o��A$�㹅� Ÿ��:�/���,'��}?��|W��(o��?������$���?���=��S��ҴŻ�.л�{ڻ��ה��`��'�(���d
�����w�����=�� �z�$���(���,�#�0�R�4�k�8�U�<�io@�k+D���G��}K��O���R��$V�ҜY��]��p`���c�R"g��nj�)�m�1�p�)t�gZw�R�z��}�9e���򁼣}��v��������Ք�����������*���v��`���)����u��i얼b���֙��J������u0��^����������$���He��զ��D��8���k#����������p���߰�O��<����-���������|����]���ν��  �  ��N=�M=0/M=�uL=��K=3K=hFJ==�I=��H=|H=�VG=��F=
�E=�E=�^D=Z�C=#�B=/B=y\A=�@=��?=<?=�L>=��==;�<=��;=-;=b:=ٕ9=4�8=.�7=�(7=�V6=��5=<�4=��3=��2=�!2=;D1=�d0=�/=��.=�-=r�,=6�+=�*=� *=r)=�(=�'=�&=e%=$=� #=Q�!=�� =��=ڨ=��=ja=c6=J=�=��=�V=�=��=�v=� =x�=�d=�=��=f 
=t�=-=n�=�$=��=�=���<��<�p�<�)�<<��<N��<`"�<Ǻ�<�K�<���<-Y�<���<�L�<���<�)�<-��<���<-O�<!��<*��<�N�<y��<<�<�.�<&t�<���<��<s5�<�q�<���<'�<t�<�U�<��<���<P��<'Yz<m�r<[.k<ƙc<�\<�tT<��L<WE<��=<�C6<�.<�='<��<�H<=�<g	<��<�9�;~��;���;*C�;Q��;E�;��;ʑ�;�V�;df;�HJ;�].;��;	E�:q��:D��:r�:,�59��o��B$������Ÿ�v;�b���-'��~?��}W�W)o��@���������K@���=������Ż�.л+|ڻ<��p�`��� ����rd
����_w����a=��� �4�$���(�G�,���0���4�F�8�'�<�2o@�J+D�~�G�~K��O���R��$V���Y��]�5q`��c�x"g�Noj�_�m�u�p��)t��Zw���z���}�Le���򁼶}����2�������������r���������J��H�������u��C얼�a���֙��J��ӽ��U0��N�������������9e��.զ��D��C���~#����������p��఼O��e����-��:�������|��1��]���ν��  �  ��N=��M=2/M=�uL=��K=.K=pFJ=@�I=��H=�H=�VG=ęF= �E=�E=�^D=q�C=6�B=;B=�\A=��@=��?==?=�L>=��===�<=��;=
-;=b:=Ε9=.�8=�7=�(7=pV6=��5=+�4=��3=��2=y!2=2D1=�d0=�/=��.=�-=y�,=7�+=�*=� *=s)=�(=�'=�&=p%= $=� #=i�!=�� =��=�=��=xa=l6=X=�=��=�V=�=��=�v=� =n�={d=��=�=[ 
=Z�=�,=X�=�$=��=�=���<��<�p�<�)�<4��<U��<]"�<ʺ�<�K�<���<+Y�<��<�L�<	��<�)�<L��<��<:O�<G��<Y��<�N�<���<T�< /�</t�<̶�<��<k5�<�q�<ì�<3�<Z�<�U�<���<���<5��<�Xz<1�r<
.k<��c<8\<qtT<~�L<�VE<��=<�C6<��.<�='<��<�H<*�<1g	<��<(:�;ރ�;���;�C�;��;�E�;��;���;�W�;�df;nIJ;r^.;إ;�E�:���:���:��:�59�o�DB$�л��|Ƹ�!=뺦���.'��?��~W�t*o��@����������@��L>�����_�Żu.л|ڻ��仩��t`��� �ۼ�1d
����"w�����<�j� ��$�7�(��,���0���4�	�8��<�(o@�<+D���G��}K��O�r�R��$V�(�Y��]�rq`�9�c��"g��oj���m���p�*t��Zw���z��}�[e���򁼸}��s��0������Δ�����q���v������8��-��������u��5얼�a���֙��J������>0��-�������������Be��"զ��D��7����#��Ȓ�����	q��఼HO�������-��W���
���|��B��]���ν��  �  y�N=y�M=#/M=�uL=��K=8K={FJ=B�I=��H=�H=�VG=֙F=$�E=�E=�^D=w�C=<�B=MB=�\A=�@=��?=<?= M>=��==A�<=��;=�,;=b:=Õ9='�8=�7=�(7=`V6=��5=&�4=��3=��2=i!2=&D1=�d0=؂/=��.=ַ-=j�,=,�+=�*=� *=�)=�(=�'=�&=o%=.$=� #=m�!=�� =��=��=��=�a=k6=a=�=��=�V=�=��=�v=� =a�=rd=��=ؑ=M 
=F�=�,=I�=w$=��=�=���<Ԯ�<�p�<�)�<��</��<L"�<κ�<�K�<���<&Y�<(��<M�<��<�)�<\��< ��<RO�<T��<`��<�N�<���<V�<8/�<7t�<߶�<4��<o5�<�q�<���<�<F�<�U�<㋈<���<��<�Xz< �r<�-k<r�c<
\<9tT<[�L<�VE<��=<rC6<ʾ.<�='<��<�H<P�<^g	<�<�:�;��;U��;D�;7��;F�;p�;Ӓ�;�W�;7ff;�IJ;�^.;ʦ;�E�:��:���:�:�59��o��D$�޼��Ǹ�g>�����/'��?��~W�Q+o��@���4���@���>������Ż�.лm|ڻڝ仞���_��� ����d
�����v�\���<�L� �ݹ$�(�(���,�j�0���4���8��<�o@��*D���G��}K��O���R�%V�C�Y� ]��q`�g�c�#g��oj�ߴm���p�*t�1[w�݅z��}�ke�����}�����=������Ŕ�����s���[��쏏�/���������xu��얼�a���֙�oJ������=0��������t�������>e��"զ��D��M����#��В����q��8఼aO�������-��`��� ��}��R��]���ν��  �  }�N=|�M=,/M=�uL=��K=3K=pFJ=J�I=��H=�H=�VG=ٙF=+�E=�E=_D=}�C=D�B=MB=�\A=�@=��?=B?=�L>=��==;�<=��;=-;=b:=ĕ9=�8=�7=~(7=^V6=��5=�4=��3=��2=k!2=D1=�d0=҂/=��.=ܷ-=o�,=4�+=�*=� *=x)=�(=�'=�&=~%=/$=� #=s�!=�� =��=��=��=�a=z6=`=$�=��=�V=�=��=�v=� =g�=nd=��=Ց=C 
=G�=�,=<�=g$=~�=�=���<̮�<�p�<�)�<!��<=��<X"�<���<�K�<���<-Y�<1��<M�<,��<�)�<l��<,��<}O�<o��<o��<�N�<���<q�<9/�<Gt�<϶�<(��<j5�<�q�<���<%�<M�<yU�<׋�<���<��<�Xz<��r<�-k</�c<�\<$tT<2�L<�VE<�=<~C6<׾.<�='<��<�H<=�<5g	<$�<�:�;T��;���;:D�;w��;jF�;*�;��;$X�;Cff;�JJ;]_.;/�;�F�:���:���:�:׆59	�o�'C$�����Iȸ��>뺮���/'�n�?��W��+o�xA������r��A���>��0��w�Ż�.л(|ڻ�仦��D`��� ����d
�D���v�3���<�� ���$��(���,�q�0���4���8�ǥ<�"o@�++D���G��}K��O���R��$V�O�Y�]��q`���c�#g��oj��m��p�M*t�.[w��z�%�}�~e�����}�����/������ǔ�����j���P��珏���	�������ku���떼�a��r֙�bJ������"0���������������De��$զ��D��F����#��㒬���'q��F఼eO������.������(�� }��e�^��Ͻ��  �  x�N=n�M=&/M=�uL=��K=@K=yFJ=S�I=��H=�H=�VG=ۙF=8�E=�E=_D=|�C=P�B=KB=�\A=�@=��?=L?=�L>=��==>�<=��;=�,;=�a:=9=�8=�7=y(7=`V6=��5=�4=��3=��2=k!2=D1=�d0=ւ/=��.=շ-=b�,=1�+=
�*=� *=�)=�(=�'=�&=�%=-$=� #=v�!=�� =��=��=��=�a=�6=W=%�=��=�V=�=��=�v=� =]�=jd=��=֑=; 
=I�=�,=H�=k$=w�=�=���<ծ�<�p�<�)�<��<)��<R"�<���<�K�<���<EY�<%��<�L�<A��<�)�<���<+��<hO�<f��<���<�N�<���<�<&/�<Ut�<ⶦ<?��<z5�<�q�<���<	�<B�<tU�<勈<���<��<�Xz<��r<�-k<$�c<�\<tT<.�L<�VE<t�=<lC6<��.<�='<��<�H<t�<Yg	<F�<O:�;n��;���;JD�;Ἲ;PF�;��;��;�X�;*ff;WKJ;8_.;��;�G�:e��:���:��:�59C�o�uF$�׼��+ȸ��=���r/'��?��W��*o��A���������A���>��B����Ż!/лB|ڻ��6��`��� ����%d
����v����<�+� ���$��(���,�{�0�`�4� �8�å<��n@�+D�Y�G��}K��O�͢R�%V�\�Y�]��q`���c�#g��oj�شm��p�k*t�[w�&�z��}�|e�����}�����5�������������R���]��򏏼�
���������mu��얼�a��_֙�_J������0��'���u��r�������4e��(զ��D��a����#��璬� ��'q��L఼hO�������-������/��#}��g��]��Ͻ��  �  }�N=|�M=,/M=�uL=��K=3K=pFJ=J�I=��H=�H=�VG=ٙF=+�E=�E=_D=}�C=D�B=MB=�\A=�@=��?=B?=�L>=��==;�<=��;=-;=b:=ĕ9=�8=�7=~(7=^V6=��5=�4=��3=��2=k!2=D1=�d0=҂/=��.=ܷ-=o�,=4�+=�*=� *=x)=�(=�'=�&=~%=/$=� #=s�!=�� =��=��=��=�a=z6=`=$�=��=�V=�=��=�v=� =g�=nd=��=֑=C 
=G�=�,=<�=g$=�=�=���<ͮ�<�p�<�)�<"��<>��<Y"�<���<�K�<���<.Y�<2��<M�<,��<�)�<l��<,��<~O�<o��<o��<�N�<���<q�<9/�<Ft�<ζ�<(��<i5�<�q�<���<$�<M�<xU�<׋�<���<��<�Xz<��r<�-k</�c<�\<$tT<3�L<�VE<��=<C6<ؾ.<�='<��<�H<?�<6g	<%�<�:�;V��;���;;D�;x��;jF�;*�;��;"X�;?ff;�JJ;W_.;)�;�F�:���:���:�:K�59��o�LC$�����[ȸ��>뺷���/'�v�?��W��+o�{A�� �u��A���>��2��y�Ż�.л*|ڻ�仨��E`��� ����d
�E���v�3���<�� ���$��(���,�q�0���4���8�ǥ<�#o@�++D���G��}K��O���R��$V�O�Y�]��q`���c�#g��oj��m��p�M*t�.[w��z�%�}�~e�����}�����/������ǔ�����j���P��珏���	�������ku���떼�a��r֙�bJ������"0���������������De��$զ��D��F����#��㒬���'q��F఼eO������.������(�� }��e�^��Ͻ��  �  y�N=y�M=#/M=�uL=��K=8K={FJ=B�I=��H=�H=�VG=֙F=$�E=�E=�^D=w�C=<�B=MB=�\A=�@=��?=<?= M>=��==A�<=��;=�,;=b:=Õ9='�8=�7=�(7=`V6=��5=&�4=��3=��2=i!2=&D1=�d0=؂/=��.=ַ-=j�,=,�+=�*=� *=�)=�(=�'=�&=o%=.$=� #=m�!=�� =��=��=��=�a=k6=a=�=��=�V=�=��=�v=� =b�=rd=��=ّ=N 
=F�=�,=I�=x$=��=�=���<֮�<�p�<�)�<��<1��<N"�<Ϻ�<�K�<���<(Y�<)��<M�<��<�)�<\��<!��<RO�<T��<_��<�N�<���<U�<7/�<5t�<޶�<3��<n5�<�q�<���<�<E�<�U�<⋈<���<��<�Xz< �r<�-k<r�c<\<:tT<]�L<�VE<��=<tC6<̾.<�='<��<�H<S�<`g	<�<�:�;���;X��;D�;8��;F�;o�;ђ�;�W�;0ff;�IJ;�^.;��;�E�:���:���:پ:�59��o��D$����AǸ��>����/'��?�W�_+o��@���:���@���>������Ż�.лp|ڻݝ仠���_��� ����d
�����v�\���<�L� �ݹ$�(�(���,�j�0���4���8��<�o@��*D���G��}K��O���R�%V�C�Y� ]��q`�g�c�#g��oj�ߴm���p�*t�1[w�݅z��}�ke�����}�����=������Ŕ�����s���[��쏏�/���������xu��얼�a���֙�oJ������=0��������t�������>e��"զ��D��M����#��В����q��8఼aO�������-��`��� ��}��R��]���ν��  �  ��N=��M=2/M=�uL=��K=.K=pFJ=@�I=��H=�H=�VG=ęF= �E=�E=�^D=q�C=6�B=;B=�\A=��@=��?==?=�L>=��===�<=��;=
-;=b:=Ε9=.�8=�7=�(7=pV6=��5=+�4=��3=��2=y!2=2D1=�d0=�/=��.=�-=y�,=7�+=�*=� *=s)=�(=�'=�&=p%= $=� #=i�!=�� =��=�=��=ya=l6=X=�=��=�V=�=��=�v=� =o�=|d=��=�=\ 
=[�=�,=Y�=�$=��=�=���<��<�p�<�)�<7��<X��<`"�<̺�<�K�<���<-Y�<��<�L�<��<�)�<M��<��<:O�<G��<X��<�N�<���<S�</�<-t�<˶�<��<i5�<�q�<���<1�<X�<�U�<���<���<4��<�Xz<0�r<
.k<��c<9\<stT<��L<�VE<��=<�C6<��.<�='<��<�H<.�<4g	<��<.:�;��;���;�C�;��;�E�;��;���;�W�;�df;bIJ;c^.;ǥ;`E�:ͭ�:���:$�:i�59��o��B$�����Ƹ�R=뺾���.'��?��~W��*o��@����������@��R>�����e�Żz.л"|ڻ��们��w`��� �ܼ�1d
����"w�����<�k� ��$�7�(��,���0���4�	�8��<�(o@�<+D���G��}K��O�r�R��$V�(�Y��]�rq`�9�c��"g��oj���m���p�*t��Zw���z��}�[e���򁼸}��s��0������Δ�����q���v������8��-��������u��5얼�a���֙��J������>0��-�������������Be��"զ��D��7����#��Ȓ�����	q��఼HO�������-��W���
���|��B��]���ν��  �  ��N=�M=0/M=�uL=��K=3K=hFJ==�I=��H=|H=�VG=��F=
�E=�E=�^D=Z�C=#�B=/B=y\A=�@=��?=<?=�L>=��==;�<=��;=-;=b:=ٕ9=4�8=.�7=�(7=�V6=��5=<�4=��3=��2=�!2=;D1=�d0=�/=��.=�-=r�,=6�+=�*=� *=r)=�(=�'=�&=e%=$=� #=Q�!=�� =��=ڨ=��=ka=c6=J=�=��=�V=�=��=�v=� =x�=�d=�=��=g 
=u�=-=p�=�$=��=�=���<��<�p�<�)�<?��<Q��<d"�<ʺ�<�K�<���<0Y�<���<�L�<���<�)�<.��<���<-O�<!��<)��<�N�<x��<;�<�.�<$t�<���<��<q5�<�q�<���<$�<r�<�U�<��<���<O��<&Yz<m�r<[.k<Ǚc<�\<�tT<��L<WE<��=<�C6<�.<�='<��<�H<B�<g	<��<�9�;���;���;-C�;S��;E�;��;Ǒ�;�V�;�cf;�HJ;�].;ߤ;�D�:>��:��: �:Q~59h�o�mC$�����7Ƹ��;����-'��~?��}W�p)o��@���������T@��>�����#�Ż�.л1|ڻA��t�`��� ����td
����`w����b=��� �5�$���(�G�,���0���4�F�8�'�<�2o@�J+D�~�G�~K��O���R��$V���Y��]�5q`��c�x"g�Noj�_�m�u�p��)t��Zw���z���}�Le���򁼶}����2�������������r���������J��H�������u��C얼�a���֙��J��ӽ��U0��N�������������9e��.զ��D��C���~#����������p��఼O��e����-��:�������|��1��]���ν��  �  ��N=��M=6/M=�uL=��K=)K=cFJ=.�I=��H=mH=�VG=��F=��E=�E=�^D=I�C=�B="B=d\A=�@=y�?=,?=�L>=��==9�<=��;=	-;=b:=�9=?�8=9�7=�(7=�V6=̂5=N�4= �3=��2=�!2=LD1=�d0=��/=��.=��-=u�,=A�+=�*=� *=i)=�(=�'=�&=S%=$=� #=A�!=�� =t�=ʨ=}�=_a=P6=C=�=��=�V=�=��=�v=� =��=�d=�=�=} 
=��='-=��=�$=��=�=,��<9��<q�<
*�<Z��<b��<�"�<κ�<�K�<���<Y�<���<�L�<ҽ�<�)�<��<���<O�< ��<��<mN�<R��<�<�.�<t�<���<	��<`5�<�q�<̬�</�<��<�U�<(��<<t��<WYz<��r<�.k<�c<�\<�tT<�L<>WE<�=<D6<�.<>'<�<�H<�<g	<��<c9�;��;���;�B�;���;�D�;�;(��;LV�;�bf;GJ;�\.;�;nB�:V��:.��:h�:k�59�o�GB$�(���EŸ��:�P���,'��}?��|W��(o��?������/���?���=��[��ٴŻ�.л�{ڻ��۔��`��)�*���d
� ���w�����=�� �{�$���(���,�#�0�R�4�l�8�U�<�io@�k+D���G��}K��O���R��$V�ҜY��]��p`���c�R"g��nj�)�m�1�p�)t�gZw�R�z��}�9e���򁼣}��v��������Ք�����������*���v��`���)����u��i얼b���֙��J������u0��^����������$���He��զ��D��8���k#����������p���߰�O��<����-���������|����]���ν��  �  ��N=��M=7/M=�uL=��K=#K=_FJ=%�I=~�H=]H=�VG=��F=��E=�E=�^D=9�C=��B=B=W\A=ԙ@=p�?=%?=�L>=��==:�<=��;=-;=(b:=�9=Q�8=F�7=�(7=�V6=��5=e�4=�3=��2=�!2=`D1=�d0=
�/=Ȟ.=��-=��,==�+=�*=� *=g)=�(=�'=�&=F%=�$=� #=2�!=|� =_�=��=f�=Pa=F6=6= �=��=�V=�=��=�v=� =��=�d=&�=�=� 
=��=A-=��=�$=ؘ=�=\��<Z��<3q�<!*�<~��<w��<�"�<׺�<�K�<���<Y�<���<�L�<���<d)�<��<���<�N�<ܧ�<���<@N�<5��<��<�.�<�s�<���<���<_5�<�q�<ɬ�<M�<��<�U�<J��<<���<�Yz<$�r<�.k<��c<\<AuT<@�L<�WE<T�=<D6<N�.<>'<�<�H<�<�f	<��<
9�;}��;s��;�A�;	��;�C�;*��;���;U�;�af;�EJ;K[.;;�;A�:{��:-��:��:\59��o�g?$�����fø�y9�Y��#,'��|?��{W��'o�W?��Q�������?��D=������ŻQ.л|ڻ$�����`��8�N���d
�8���w�[���=�?� �պ$�&�(���,�d�0���4���8�y�<�zo@�s+D���G��}K��O�Y�R�w$V���Y�E]��p`���c�"g��nj�ֳm���p�.)t�+Zw��z�N�}�e���򁼇}��h��!������ޔ�����������I����������V����u���얼8b���֙��J������0��t����������-���He�� զ��D�����^#����������p���߰��N�����p-��✶�����|���캼�]���ν��  �  ��N=��M=</M=�uL=��K=!K=PFJ= �I=o�H=NH=�VG=��F=��E=�E=�^D=#�C=��B=�B=K\A=Ù@=c�?=?=�L>=��==;�<=��;=-;=,b:=�9=\�8=V�7=�(7=�V6=�5=w�4=,�3=��2=�!2=rD1=�d0=�/=О.=�-=��,=A�+=�*=� *=`)=�(=z'=�&=;%=�$=� #=�!=h� =K�=��=Y�==a=<6='=��=��=�V=�=��=�v=� =��=�d=9�=,�=� 
=��=T-=��=�$=�=	=���<���<Vq�<9*�<���<���<�"�<޺�<�K�<���<Y�<���<�L�<���<@)�<Ǐ�<~��<�N�<���<���< N�<��<��<�.�<�s�<���<���<c5�<�q�<Ѭ�<S�<��<�U�<l��<;<���<�Yz<i�r<J/k<ƚc<l\<�uT<�L<�WE<��=<CD6<_�.<->'<�<�H<��<�f	<v�<�8�;���;���;rA�;o��;C�;�ߝ;ˏ�;�T�;J`f;EJ;Z.;,�;�?�:��::�:`{59��o�5?$�%���^¸��7뺧���*'��{?��zW�J&o��>��������(?���<�����{�Ż<.л�{ڻ3��Ȕ�6a��p�r��e
�i��,x����A>��� �,�$���(�"�,���0���4���8���<��o@��+D���G��}K��O�P�R�e$V���Y�
]��p`�>�c��!g�jnj�z�m���p��(t��Yw�΄z��}��d��r򁼀}��d��"������֔��)���������k����������s���v���얼fb��"י�	K��6����0���������Ǆ��7���Be��!զ��D�����O#��u���|���p���߰��N���:-����|��q|���캼r]���ν��  �  ��N=��M=G/M=�uL=��K=K=IFJ=�I=c�H=EH=�VG=x�F=��E=yE=�^D=�C=��B=�B=7\A=��@=W�?=?=�L>=��==2�<=��;=-;=4b:=��9=d�8=f�7=�(7=�V6=�5=��4=?�3=�2=�!2=~D1=�d0=#�/=ڞ.=�-=��,=N�+=�*=� *=[)=�(=p'=�&=-%=�$=� #=�!=Y� =>�=��=Q�=,a=-6= =��=~�=�V=�=��=�v=� =��=�d=F�=D�=� 
=ũ=k-=̫=�$=�==���<���<mq�<[*�<���<���<�"�<պ�<�K�<���<�X�<���<�L�<���<)�<���<S��<�N�<���<���<N�<囵<��<�.�<�s�<s��<���<M5�<�q�<笗<Y�<��<�U�<���<e<���<<Zz<��r<�/k<�c<�\<�uT<��L<XE<��=<�D6<v�.<[>'<-�<~H<��<�f	<M�<+8�;���;9��;�@�;�;mB�;ߝ;	��;�T�;�^f;�CJ;?Y.;>�;>�:��:p��:2�:{�59�o�&>$���������36뺵��&*'��z?��yW�<%o�i>��3�������>���<������Ż.л�{ڻ?��7��ca�������@e
����x�����>�څ �g�$���(�I�,��0���4��8�Ʀ<��o@��+D���G�~K�jO�3�R�+$V�a�Y��
]�@p`��c�z!g�nj�3�m�F�p��(t��Yw���z�̩}��d��X�m}��Q��������ꔉ�2��Õ�����������΅������Jv���얼�b��@י�'K��a����0���������ք��>���We��զ��D�����0#��a���c��op��߰��N��ͽ��-������Y��X|���캼U]���ν��  �  ��N=��M=A/M=�uL=��K=K=LFJ=	�I=\�H=7H=�VG=h�F=��E=jE=�^D=��C=��B=�B=+\A=��@=P�?=?=�L>=��==9�<=��;=-;=9b:=�9=u�8=r�7=�(7=�V6=�5=��4=G�3=�2=�!2=�D1=e0=1�/=�.=�-=��,=E�+=�*=� *=c)=�(=f'=�&=%=�$=r #=��!=G� =,�=��=;�=&a=6==��=z�=�V=�=��=�v=� =��=�d=X�=R�=� 
=ԩ=�-=۫=%=�=(=���<ȯ�<�q�<l*�<���<���<�"�<��<�K�<���<�X�<���<nL�<j��<)�<���<9��<pN�<i��<w��<�M�<כ�<��<�.�<�s�<t��<���<Q5�<�q�<ج�<l�<��<V�<���<|<���<�Zz<�r<�/k<f�c<\<vT<�L<8XE<��=<�D6<��.<F>'<*�<�H<��<�f	<�<�7�;3��;���;W@�;A��;�A�;iޝ;���;�S�;^f;�BJ;UX.;��;;<�:���:B��::�:%x59��o�d=$�y�����5�����)'��y?��xW��$o��=��˾��g��G>��1<��R���Ż�-л�{ڻ��3��0a����Ƚ�ce
�����x����>�$� ���$��(���,� �0�4�4�9�8��<��o@��+D���G��}K��O�#�R�$$V�D�Y��
]�p`���c�L!g��mj��m��p�G(t�mYw�R�z���}��d��M�d}��O��������蔉�#��ؕ��������������������ev��햼�b��gי�KK��o����0��������Ԅ��7���Re��զ��D������,#��I���M��Xp��i߰�qN������-��w���/��D|���캼?]��gν��  �  ��N=��M=I/M=�uL=��K=K=BFJ= �I=X�H=)H=�VG=Z�F=��E=eE=z^D=��C=��B=�B=#\A=��@=K�?=�?=�L>=��==:�<=��;='-;=Ab:=�9=��8=r�7=�(7=�V6=�5=��4=R�3=!�2=�!2=�D1=
e0=:�/=�.=�-=��,=I�+=�*=� *=R)=�(=^'=�&=%=�$=a #=��!=@� ="�=��=*�=a=6==��=q�=�V=�=��=�v=!=��=�d=d�=U�=� 
=�=�-=�=%=$�=9=���<̯�<�q�<}*�<���<ł�<�"�<��<�K�<���<�X�<���<XL�<[��<�(�<i��<3��<RN�<_��<h��<�M�<ț�<��<|.�<�s�<^��<���<H5�<�q�<嬗<��<��<,V�<���<�<��<�Zz<)�r<�/k<��c<$\<NvT<2�L<EXE<�=<�D6<Ϳ.<j>'<<�<�H<��<|f	<��<�7�;���;���;�?�;췺;�A�;�ݝ;b��;@S�;.]f;BJ;_W.;/�;�:�:���:C��:�:`w59��o��;$�0���ʾ��95�V���('�jy?�`xW�7$o��=���������4>���;������Żz-л�{ڻ��r�a�������e
����x�g���>�D� �߻$��(���,�L�0�\�4�_�8��<�p@��+D���G��}K��O��R�!$V��Y��
]�p`���c�!g��mj��m���p�8(t�6Yw��z���}��d��A�W}��2�������� ���?��알�������������������lv�� 햼�b��vי�jK��}����0��Ƣ����ꄢ�W���\e��զ��D��ݳ��,#��0���D��Hp��D߰�fN�������,��i���'�� |��|캼:]��Nν��  �  ¡N=��M=F/M=�uL=��K=K=FFJ=�I=N�H=%H=~VG=V�F=��E=UE=p^D=�C=��B=�B=\A=��@=C�?=?=�L>=��==8�<=��;= -;=:b:=�9=��8=��7=�(7=�V6=%�5=��4=h�3='�2=�!2=�D1=e0=;�/=��.=�-=��,=I�+=�*=� *=Z)=�(=]'=�&=%=�$=c #=��!=1� =�=u�=-�=a=6=	=��=y�=�V=�=��=�v=!=��=�d=e�=f�=� 
=�=�-=��=#%=-�=D=���<��<�q�<�*�<���<���<�"�<��<�K�<���<�X�<���<ML�<T��<�(�<l��<��<?N�<B��<W��<�M�<���<��<g.�<�s�<g��<���<N5�<�q�<ଗ<o�<��<6V�<���<�<��<�Zz<H�r<E0k<��c<D\<ZvT<U�L<oXE<+�=<�D6<��.<]>'<*�<�H<��<�f	<��<n7�;���;S��;�?�;���;2A�;�ݝ;ύ�;/S�;�\f;�AJ;�V.;��;�:�:��:9��:�:�s59�o��=$�`���꾸��3�!��l('��x?��wW��"o�q=��E�������=���;�������Ż�-л�{ڻD��8��a�������e
����x�`��?��� ��$�W�(���,�s�0�a�4�z�8��<��o@��+D���G�~K��O��R�$V���Y��
]��o`���c�� g��mj���m���p�(t�Yw��z�e�}��d��1�c}��E��������𔉼6��ᕌ������� ��	��������v��3햼�b���י�oK������1��ۢ����ᄢ�D���Ue��զ��D������ #��&���6��2p��C߰�VN�������,��W�����|��k캼&]��Hν��  �  �N=1�M=)M=|nL=��K=`�J=�<J=��I=�H=H=oIG=\�F=��E=jE=�MD=��C=��B=�	B=�FA=�@=��?=�>=�2>=k==X�<=��;=�;='A:=�s9=f�8=��7=�7=.6=�X5=x�4=n�3=v�2=|�1=>1=�/0=L/=�e.=#}-=��,=e�+=-�*=��)=��(=��'=��&=��%=��$=a�#=M�"=�!=�� =�o=�Q=/=�=B�=�=�s=�8=�=c�=Lg=�=�=�e=2=(�=�3=��	=�L=��=8Q=��=PA=� =�;�<�
�<>��<E��<�A�<4��<���<�/�<g��<T�<K��<(^�<���<P�<���<|,�<J��<���<�S�<뭼<b�<LW�<$��< ��<,>�<���<ˢ<\�<�O�<���<�͓<�
�<�F�<6��<ռ�<���<
bz<��r<�Ik<}�c<�4\<ëT<�$M<T�E<:><Y�6<�#/<ɫ'<�7 <��<�^<��	<4�<X��;��;7M�;^��;T�;+�;J��;�d�;�=�;mXj;�cN;^�2;�;�`�:��:H:�:��+:���9o�����6pu�ȇ����ߺ.��/?!��y9�UeQ���h��#�������f������෻%�»<ͻvQ׻�w�s�VE��;���7�O���{��s����� �m]#���'��+�:�/���3���7��v;��G?��C��F�onJ�N���Q��,U�ެX�0#\�>�_���b�~Pf���i� �l�T6p��ts�t�v�\�y�+
}�Y��騁�7�����L��Tԇ�Z���݊�+`�������_���ݐ��Y���ԓ��N��rǖ�3?��뵙��+������M����������n���ࣼ�R��Ħ�65��0����������0����h��Iٰ��I������q+��t������<���dc��'ֽ��  �  �N=0�M=)M=}nL=��K=_�J=�<J=��I=�H=H=zIG=^�F=��E=rE=�MD=��C=��B=�	B=�FA=#�@=��?=�>=�2>=�j==Y�<=��;=|;=(A:=�s9=o�8=��7=�7=.6=�X5=z�4=t�3=r�2=h�1=?1=�/0=L/=�e.= }-=��,=b�+=2�*=��)=��(=��'=��&=��%=��$=o�#=I�"=�!=�� =�o=�Q=�.=�=K�=�=�s=�8=$�=`�=Pg=�=�=�e=5=(�=�3=��	=�L=��=<Q=��=IA=�� =�;�<�
�<J��<D��<�A�<(��<���<�/�<]��<6T�<P��< ^�<���<!P�<���<{,�<Z��<���<�S�<譼<_�<eW�<0��<��<!>�<ʅ�<ˢ<W�<�O�<���<�͓<�
�<G�<5��<˼�<���<�az<��r<�Ik<�c<T4\<��T<�$M<N�E<[><J�6<�#/<��'<�7 <��<�^<
�	<�<R��; ��;�M�;p��;T�;m�;c��;;e�;�=�;�Xj;]dN;��2;�;�`�:/�:�9�:��+:��9���T���ou�������ߺ2���?!�:z9�'eQ�(�h��#��W����������p෻;�»>ͻ�Q׻aw�%s�E������)7�8���{�� � s���� �W]#�؈'��+��/�ת3��7��v;��G?��C��F�]nJ�N�ĢQ��,U�ϬX�-#\�X�_���b��Pf���i��l�K6p��ts���v�W�y�5
}�K��騁�7�����L��Qԇ�Z���݊�%`�������_��oݐ��Y���ԓ��N��iǖ�?����+��⠜�B����������n���ࣼ�R��Ħ�?5��1����������1����h��Rٰ��I������b+��s������J��$�gc��ֽ��  �  �N=4�M=�(M=�nL=��K=[�J=�<J=��I=�H=H=}IG=b�F=��E=yE=�MD=�C=��B=�	B=�FA=(�@=��?=�>=�2>=�j==`�<=��;=|;=)A:=xs9=i�8=��7=�7=.6=�X5=t�4=h�3=p�2=f�1=H1=�/0=L/=�e.=}-=��,=a�+=8�*=�)=��(=��'=��&=�%=��$=s�#=K�"=�!=�� =�o=�Q=/=�=H�=$�=�s=�8= �=Z�=Vg=�=�=�e=/= �=�3=��	=�L=��=/Q=��=IA=�� =�;�<�
�<=��</��<�A�<(��<���<�/�<P��<0T�<M��<,^�<��<P�<���<z,�<i��<���<�S�<�<e�<nW�<1��<��<!>�<Ʌ�<ˢ<]�<�O�<|��<�͓<�
�<�F�<%��<Ǽ�<��<�az<��r<�Ik<l�c<L4\<ëT<�$M<(�E<B><'�6<�#/<��'<8 <��<�^<�	< �<���;0��;�M�;���;%T�;��;p��;�e�;�=�;1Yj;udN;�2;-;�`�:�:�9�:�+:�9������"ru�6�����ߺ	���?!�+z9��eQ���h��#��g���f���&���෻i�»!ͻ�Q׻,w�9s�/E������"7����{�� �s����� �I]#���'��+���/��3���7��v;��G?��C�,�F�BnJ�N���Q��,U��X�F#\�w�_���b��Pf���i�;�l�q6p��ts���v�H�y�Y
}�W������7�����L��@ԇ�Z���݊�(`�������_��qݐ��Y���ԓ��N��hǖ�?��浙��+��ؠ��A��戟�����n���ࣼ�R��	Ħ�E5��,���������@����h��@ٰ��I������{+��|������;��%�xc��!ֽ��  �  �N=+�M=�(M={nL=��K=e�J=�<J=��I=�H=H=�IG=o�F=��E=~E=�MD=�C=��B=�	B=�FA=-�@=��?=�>=�2>=k==[�<=��;=u;="A:=ws9=a�8=��7=�7= .6=�X5=m�4=b�3=f�2=^�1=21=�/0=L/=�e.=}-=��,=]�+=/�*=��)=��(=��'=��&=�%=��$=y�#=Z�"=$�!=�� =�o=�Q=/=�=Q�=$�=�s=�8=#�=d�=Kg=�=�=�e=&=�=�3=��	=�L=��=&Q=��=:A=� =�;�<v
�<,��<'��<�A�<��<���<�/�<f��<.T�<U��<2^�<��<.P�<���<�,�<s��<���<�S�<��<��<zW�<A��<��<2>�<̅�<#ˢ<f�<�O�<x��<�͓<�
�<�F�<!��<���<���<�az<b�r<zIk<K�c<#4\<y�T<�$M<�E<><*�6<|#/<��'<�7 <��<�^<�	<A�<���;k��;�M�;��;�T�;��;ʡ�;�e�;T>�;Zj;	eN;}�2;q;�a�:E�:K;�:�+:��98��,���qu�ᇭ��ߺѷ�X@!��z9��eQ�/ i�#$���������0���෻c�»eͻ�Q׻mw��r��D������7����{�� ��r����� �+]#���'���+�Ԯ/���3���7��v;��G?��C���F�gnJ�-N��Q��,U���X�V#\���_���b��Pf��i�U�l��6p��ts�Ҭv���y�f
}�c������)7��Ä��L��Oԇ� Z���݊�`�������_��_ݐ��Y���ԓ��N��Tǖ�?��˵���+��͠��2��鈟�����n���ࣼ�R��Ħ�J5��=���������D����h��hٰ�J�������+���������_��;�}c��2ֽ��  �  �N="�M=)M=~nL=��K=e�J=�<J=��I=�H=H=�IG=r�F=��E=�E=�MD=�C=��B=�	B=�FA=7�@=��?="�>=�2>=	k==S�<=��;=y;=A:=vs9=V�8=��7=�7=�-6=�X5=_�4=X�3=U�2=X�1=)1=�/0=L/=�e.=}-=��,=i�+=-�*=��)=��(=��'=��&=�%=��$=~�#=^�"=+�!=ʉ =p=�Q=/=�=_�='�=�s=�8= �=b�=Fg=�= �=�e==�=�3=��	=�L=~�=Q=��=(A=� =�;�<h
�<��<��<�A�<��<���<�/�<f��<+T�<j��<9^�<��<EP�<���<�,�<���<���<�S�<��<��<�W�<a��<��<K>�<ׅ�<$ˢ<Y�<�O�<���<�͓<�
�<�F�<��<���<���<caz<�r<WIk<�c<�3\<T�T<�$M<�E<�><#�6<V#/<��'<�7 <��<�^<�	<t�<���;���;+N�;#��;�T�;N�;l��;f�;�>�;fZj;�eN;9�2;�;�c�:��:�;�:��+:]��9���ۻ��qu����d�ߺA���@!��{9��fQ�� i��$������I��t���෻k�»�ͻFQ׻xw��r�E�������6� ��>{�� ��r����n ��\#�}�'���+�Ʈ/�z�3���7�pv;��G?��C���F�vnJ� N��Q��,U��X��#\���_��b��Pf�.�i���l��6p�(us��v���y�w
}�{�����/7��Ä��L��]ԇ��Y���݊�`�������_��Gݐ��Y���ԓ�|N��-ǖ��>�������+��������㈟������n���ࣼ�R��Ħ�35��O�����Ƈ��T����h��zٰ�J��к���+���������o��L񺼉c��Gֽ��  �  �N=!�M=�(M=}nL=��K=l�J=�<J=��I=&�H=!H=�IG=��F=��E=�E=�MD=!�C=��B=�	B=�FA=@�@=��?=$�>=�2>=k==]�<=��;=o;=A:=ks9=O�8=��7=�7=�-6=�X5=P�4=G�3=L�2=G�1=$1=�/0=�K/=�e.=}-=��,=`�+=0�*=��)=��(=��'=��&=�%=��$=��#=o�"=;�!=҉ =p=�Q=$/=�=c�=0�=�s=�8=$�=c�=Jg=�=��=�e==�=�3=��	=�L=r�=Q=��=A=ұ =�;�<F
�<���<��<�A�<���<���<�/�<i��<1T�<k��<F^�<(��<PP�<��<�,�<���<���<T�<8��<��<�W�<l��<:��<P>�<Ⅶ<3ˢ<j�<�O�<z��<�͓<�
�<�F�<���<���<���<2az<��r<�Hk<ӽc<�3\<,�T<N$M<џE<�><��6<L#/<��'<�7 <��<�^<1�	<z�<#��;��;�N�;���;\U�;��;���;�f�;/?�;�[j;�fN;�2;�;nd�:��:�<�:�+:_��9��ܻ��su�������ߺ��TA!�	|9�ygQ��i��$��:���m������0᷻��»�ͻ�Q׻Uw��r��D������6����0{�= �~r�[��K ��\#�1�'�I�+�}�/�g�3�}�7�^v;�~G?��C���F�]nJ�N��Q�-U�4�X��#\�֐_�3�b�BQf�R�i���l��6p�Ous� �v���y��
}�������77��Ä��L��Kԇ��Y���݊��_�������_��:ݐ�zY���ԓ�YN��"ǖ��>�������+������	��Ɉ�������n���ࣼ�R��Ħ�J5��S�����҇��i����h���ٰ�-J��庳��+��Ĝ��������h񺼞c��Qֽ��  �  ��N=!�M=�(M=znL=��K=i�J=�<J=��I=4�H=.H=�IG=��F=��E=�E=�MD=3�C=��B=�	B=�FA=M�@=��?=(�>=�2>=
k==Z�<=�;=n;=A:=^s9=M�8=��7=�7=�-6=sX5=E�4=9�3=D�2=3�1=1=�/0=�K/=�e.=}-=��,=Y�+=/�*=��)=��(=��'=��&=&�%=��$=��#=w�"=K�!=�� =%p=�Q=*/=�=l�=?�=�s=�8=*�=_�=Fg=�=��=�e==��=�3=��	=�L=g�=�P=y�=A=�� =t;�<%
�<���<��<�A�<���<���<�/�<`��<BT�<r��<V^�<B��<dP�<9��<�,�<ɓ�<��<9T�<U��<��<�W�<���<Y��<Y>�<���<3ˢ<e�<�O�<m��<�͓<�
�<�F�<ꁈ<o��<���<�`z<��r<�Hk<��c<s3\<�T<$M<��E<�><��6<J#/<q�'<�7 <��<�^<U�	<��<���;���;�N�;��;�U�;i�;8��;Pg�;�?�;�\j;jgN;��2;|;^e�:g�:�<�:հ+:���9i��3��`vu�������ߺT��GB!��|9��gQ�hi�%��ʟ���������p᷻�»�ͻ�Q׻Vw��r뻟D��G����6����{�	 �[r��� �}\#��'�,�+�D�/�;�3�<�7�Bv;�eG?�qC���F�`nJ�;N���Q�8-U�c�X��#\��_�`�b��Qf�r�i���l�/7p�us�h�v��y��
}����3���E7��Ä��L��Pԇ��Y���݊��_������|_��$ݐ�[Y��sԓ�3N�� ǖ��>������p+������������������n���ࣼ�R��Ħ�W5��O���/��އ��z���i���ٰ�TJ�������+��Ӝ��$�����}񺼲c��\ֽ��  �  �N=�M=�(M=|nL=��K=m�J=�<J=ÀI=9�H=8H=�IG=��F=��E=�E=�MD=;�C=��B=�	B=GA=U�@=��?=3�>=�2>=k==\�<=��;=n;=A:=Ys9==�8=��7=�7=�-6=dX5=5�4='�3=1�2=,�1=1=�/0=�K/=�e.= }-=��,=[�+=1�*=�)=��(=��'=��&=)�%=��$=��#=��"=U�!=� =2p= R=</=�=x�=C�=	t=�8=&�=d�=Eg=�=��=�e=�=�=s3=��	=�L=R�=�P=f�=�@=�� =U;�<
�<���<Ҍ�<pA�<���<���<�/�<j��<6T�<���<c^�<M��<|P�<R��<�,�<ٓ�<0��<LT�<v��<��<�W�<���<a��<u>�<���<7ˢ<p�<�O�<u��<�͓<�
�<�F�<Ё�<Z��<{��<�`z<��r<}Hk<g�c<A3\<��T<�#M<m�E<�><��6<$#/<z�'<�7 <��<�^<U�	<Û<Ć�;���;SO�;���;hV�;��;���;�g�;C@�;�]j;ZhN;��2;
;g�:|�:�=�:�+:���9l������vu�>����ߺ߹��B!��}9��hQ�ci��%������6�)��N���᷻�»�ͻ�Q׻=wộr뻜D�����|6�|���z����r������G\#�ɇ'�ޢ+��/��3�'�7�v;�DG?�xC���F�\nJ�3N��Q�P-U���X��#\�5�_���b��Qf���i�;�l�m7p��us���v�2�y�}����<���T7��Ä��L��Nԇ��Y���݊��_��p���o_��
ݐ�@Y��Kԓ�"N���Ɩ��>��a���N+��x���������������n���ࣼ�R��Ħ�P5��a���7����������,i���ٰ�iJ������+������;��������c��wֽ��  �  �N=�M=�(M=snL=��K=y�J=�<J=̀I=>�H=CH=�IG=��F=�E=�E=�MD=D�C=��B=�	B=GA=_�@=��?==�>=�2>=k==[�<={�;=f;=	A:=Ws9=0�8=��7=~7=�-6=TX5=*�4="�3=�2=�1=�1=�/0=�K/=�e.=�|-=��,=W�+=(�*=�)=��(=��'=��&=/�%=��$=��#=��"=]�!=�� =Ap=	R=L/=�=��=H�=t=�8=)�=i�=<g=�=��=�e=�=ڞ=l3=��	=�L=<�=�P=Z�=�@=�� =.;�<�	�<���<ǌ�<cA�<���<{��<�/�<x��<8T�<���<q^�<^��<�P�<[��<-�<��<T��<iT�<���<��<�W�<���<n��<�>�< ��<Nˢ<y�<�O�<j��<�͓<�
�<�F�<���<D��<W��<y`z<<�r<aHk<$�c<3\<h�T<�#M<L�E<S><��6<#/<^�'<�7 <��<_<]�	<�<��;9��;�O�;��;�V�;.��;p��;�g�;�@�;A^j;aiN;n�2;�;�h�:�:�?�:y�+:S��9������vu�����B�ߺ����C!��~9�uiQ��i�&��u�����N������᷻�»�ͻ�Q׻|w�fr�eD������R6�_���z�����q������\#���'���+���/�ȩ3��7��u;�(G?�eC���F�wnJ�=N�1�Q�]-U���X�$\�H�_���b��Qf��i�U�l��7p�vs�ԭv�t�y�}����B���[7��*Ä��L��Sԇ��Y���݊��_��`���\_���ܐ�6Y��,ԓ�N���Ɩ��>��N���3+��^��������������|n���ࣼ�R��*Ħ�[5��n���:��
�������Ai���ٰ��J��;���,�����X��������c���ֽ��  �  �N=�M=�(M=|nL=��K=p�J=�<J=΀I=H�H=IH=�IG=��F=�E=�E=�MD=U�C=�B=�	B=GA=h�@=ʾ?=>�>=�2>=k==Z�<=��;=f;=A:=Ks9=-�8=��7=w7=�-6=NX5=�4=�3=�2=�1=�1=�/0=�K/=�e.=�|-=��,=U�+=/�*=��)=��(=��'=��&=;�%=��$=��#=��"=m�!=	� =Lp=R=O/=�=��=R�=t=�8=*�=\�=?g=�=��=�e=�=Ӟ=[3=��	=}L=2�=�P=G�=�@=�� =;�<�	�<���<���<RA�<���<��<�/�<]��<FT�<���<}^�<o��<�P�<k��<$-�<	��<f��<�T�<���<
�< X�<���<���<�>�<��<Dˢ<k�<�O�<h��<�͓<�
�<�F�<���</��<P��<T`z<�r<Hk<�c<�2\<W�T<�#M<�E<E><m�6<�"/<Z�'<�7 <��<�^<~�	<�<I��;k��;P�;O��;-W�;���;���;�h�;A�;�^j;�iN;�2;Z;i�:u�:Y>�:ݲ+:s9�����Fyu�͌��*�ߺ���C!��~9�OjQ��i�B&�������𖻮����� ⷻl�»�ͻ�Q׻CwỶr�ZD������F6�.��|z�����q����_��[#�_�'���+�խ/���3�ߖ7��u;�G?�ZC���F�dnJ�AN�+�Q��-U���X�0$\���_���b�
Rf��i���l��7p�vs�߭v���y�b}����Y���h7��&Ä��L��Qԇ��Y���݊��_��Q���I_���ܐ�$Y��ԓ��M���Ɩ�d>��6���'+��L��������������pn���ࣼ�R��Ħ�]5��r���T���������Vi���ٰ��J��P���/,��.���h��������c���ֽ��  �  ۜN=�M=�(M=|nL=��K=t�J=�<J=̀I=P�H=KH=�IG=ËF=�E=�E=�MD=^�C=�B=
B=$GA=j�@=Ҿ?==�>=�2>=k==c�<=|�;=`;=A:=Ds9=.�8=��7=q7=�-6=AX5=�4=�3=�2=�1=�1=�/0=�K/=�e.=�|-=��,=H�+=7�*= �)=��(=��'=��&=@�%=��$=Ƚ#=��"=y�!=� =Qp=$R=X/=�=��=V�=t=�8=3�=_�=Gg=�=��=�e=�=ў=O3=��	=mL=(�=�P=?�=�@=�� =;�<�	�<���<���<IA�<���<l��<�/�<`��<VT�<���<�^�<q��<�P�<���<2-�<��<t��<�T�<���<(�<X�<ŧ�<���<�>�<��<Pˢ<x�<�O�<Q��<�͓<�
�<�F�<���< ��<6��<`z<��r<�Gk<ڼc<�2\<#�T<y#M<��E<@><H�6<�"/<.�'<�7 <��<�^<��	<�<���;~��;|P�;���;�W�;���; ��;�h�;cA�;Y`j;�jN;R�2;�;i�:��:�>�:��+:���9�������zu�i�����ߺZ���D!��9��jQ�Ri�k&������������$ⷻ��»�ͻR׻�vỎr�D������76���lz�D���q�R��H��[#�0�'�b�+�}�/���3�˖7��u;�G?�3C���F�>nJ�rN�;�Q��-U�ŭX�5$\���_��b�CRf�=�i���l��7p�Nvs��v���y��}����e���m7��2Ä��L��>ԇ��Y���݊��_��B���F_���ܐ��X��ԓ��M���Ɩ�V>�����	+��1������s�������`n���ࣼ�R��Ħ�u5��q���c���������ci��ڰ��J��X���B,��7����������� d���ֽ��  �  ܜN=�M=�(M=vnL=��K=w�J=�<J=րI=V�H=TH=�IG=��F=�E=�E=�MD=a�C=�B=
B='GA=q�@=ؾ?=F�>=�2>=k==^�<={�;=c;=A:=Ds9=$�8=��7=l7=�-6=<X5=�4=�3=�2=�1=�1=�/0=�K/=�e.=�|-=��,=N�+=/�*=��)=��(=��'=��&=E�%=��$=Ľ#=��"=x�!=� =]p=#R=Z/=�=��=[�=t=�8=0�=^�=?g=�=��=�e=�=ƞ=P3=��	=jL=!�=�P=9�=�@=�� =;�<�	�<���<���<HA�<���<m��<�/�<c��<OT�<���<�^�<��<�P�<���<8-�<"��<���<�T�<���<!�<X�<ק�<���<�>�<��<Qˢ<q�<�O�<X��<�͓<�
�<rF�<���<��<-��<`z<��r<�Gk<��c<�2\<�T<m#M<�E<><I�6<�"/<?�'<�7 <��<	_<��	<�<�;���;�P�;���;�W�;$��;h��; i�;zA�;�_j;�jN;ҥ2;g;Uj�:��:W?�:I�+:\��9������zu�������ߺ����D!��9��jQ�Ui��&�����1������Sⷻ��»�ͻ�Q׻>wỗr�D������6� ��Iz�W���q�U����[#�1�'�Y�+���/���3���7��u;�G?�:C���F�[nJ�ZN�-�Q��-U�٭X�Z$\���_�#�b�HRf�X�i���l� 8p�avs�&�v���y�~}����f���m7��+Ä��L��Kԇ��Y���݊��_��6���7_���ܐ�Y��	ԓ��M���Ɩ�K>�����+��4������g�������dn���ࣼ�R�� Ħ�m5��o���b��%�������fi��ڰ��J��i���E,��E�����������d���ֽ��  �  �N=�M=�(M=xnL=��K=|�J=�<J=؀I=M�H=UH=�IG=ËF=(�E=�E=�MD=d�C=%�B=
B=-GA=r�@=о?=I�>=�2>=k==Y�<=}�;=_;=�@:=Is9=!�8=��7=`7=�-6=>X5=�4=��3=�2=�1=�1=}/0=�K/=�e.=�|-=~�,=R�+=,�*=�)=��(= �'=��&=A�%=��$=��#=��"=|�!=� =Xp='R=h/=�=��=Y�=t=�8=3�=b�=;g=�=��=�e=�=��=F3=v�	=jL=�=�P=0�=�@=�� =�:�<�	�<|��<���<5A�<���<q��<~/�<h��<OT�<���<�^�<���<�P�<���<`-�<)��<��<�T�<Ю�<3�<X�<ڧ�<���<�>�<��<Zˢ<t�<�O�<`��<�͓<�
�<yF�<���<��<!��<`z<��r<�Gk<��c<�2\< �T<D#M<�E<><[�6<�"/<D�'<�7 <��<_<��	<�<y��;���;�P�;���;X�;��;/��;i�;B�;`j;8kN;�2;�;�j�:��:�?�:L�+:���9��9��)yu�������ߺg���D!��9��kQ��i��&������2��4��/ⷻ��»=ͻ�Q׻Ow�nr��C��t���6���<z�_��Zq�A��(��[#�"�'��+���/�s�3���7��u;��F?�,C���F�lnJ�MN�\�Q��-U�ȭX�t$\�Ǒ_�T�b�FRf�g�i���l� 8p�Vvs��v���y��}����^���7��8Ä��L��Uԇ��Y���݊��_��F���4_���ܐ�
Y���ӓ��M���Ɩ�P>������*��0������z�������en���ࣼ�R��Ħ�f5������^���������{i��ڰ��J��y���J,��U�����������d���ֽ��  �  ܜN=�M=�(M=vnL=��K=w�J=�<J=րI=V�H=TH=�IG=��F=�E=�E=�MD=a�C=�B=
B='GA=q�@=ؾ?=F�>=�2>=k==^�<={�;=c;=A:=Ds9=$�8=��7=l7=�-6=<X5=�4=�3=�2=�1=�1=�/0=�K/=�e.=�|-=��,=N�+=/�*=��)=��(=��'=��&=E�%=��$=Ľ#=��"=x�!=� =]p=#R=Z/=�=��=[�=t=�8=0�=^�=?g=�=��=�e=�=ƞ=P3=��	=kL=!�=�P=9�=�@=�� =;�<�	�<���<���<IA�<���<m��<�/�<c��<OT�<���<�^�<���<�P�<���<8-�<"��<���<�T�<���<!�<X�<ק�<���<�>�<��<Qˢ<p�<�O�<X��<�͓<�
�<qF�<���<��<-��<`z<��r<�Gk<��c<�2\<�T<n#M<�E<><J�6<�"/<@�'<�7 <��<
_<��	<�<ć�;���;�P�;���;�W�;$��;h��;�h�;yA�;�_j;�jN;ͥ2;b;Kj�:|�:J?�:/�+:%��9}��Ӿ��zu�������ߺ����D!��9��jQ�[i��&�����3����	��Uⷻ��»�ͻ�Q׻?wỘr�D������6� ��Iz�W���q�U����[#�1�'�Y�+���/���3���7��u;�G?�:C���F�[nJ�ZN�-�Q��-U�٭X�Z$\���_�#�b�HRf�X�i���l� 8p�avs�&�v���y�~}����f���m7��+Ä��L��Kԇ��Y���݊��_��6���7_���ܐ�Y��	ԓ��M���Ɩ�K>�����+��4������g�������dn���ࣼ�R�� Ħ�m5��o���b��%�������fi��ڰ��J��i���E,��E�����������d���ֽ��  �  ۜN=�M=�(M=|nL=��K=t�J=�<J=̀I=P�H=KH=�IG=ËF=�E=�E=�MD=^�C=�B=
B=$GA=j�@=Ҿ?==�>=�2>=k==d�<=|�;=`;=A:=Ds9=.�8=��7=q7=�-6=AX5=�4=�3=�2=�1=�1=�/0=�K/=�e.=�|-=��,=H�+=7�*= �)=��(=��'=��&=@�%=��$=Ƚ#=��"=y�!=� =Rp=$R=X/=�=��=V�=t=�8=3�=_�=Gg=�=��=�e=�=ў=O3=��	=mL=)�=�P=@�=�@=�� =;�<�	�<���<���<JA�<���<m��<�/�<a��<WT�<���<�^�<r��<�P�<���<3-�<��<t��<�T�<���<(�<X�<ħ�<���<�>�<��<Oˢ<w�<�O�<P��<�͓<�
�<�F�<���< ��<6��<`z<��r<�Gk<ۼc<�2\<$�T<z#M<��E<B><I�6<�"/<0�'<�7 <��< _<��	<�<���;���;~P�;���;�W�;���;���;�h�;aA�;T`j;�jN;J�2;�;�h�:��:�>�:^�+:]��9���/���zu������ߺg���D!��9��jQ�]i�p&�����"�������(ⷻ��»�ͻR׻ wỐr�D������86���lz�E���q�R��H��[#�0�'�b�+�}�/���3�˖7��u;�G?�3C���F�>nJ�sN�;�Q��-U�ŭX�5$\���_��b�CRf�=�i���l��7p�Nvs��v���y��}����e���m7��2Ä��L��>ԇ��Y���݊��_��B���F_���ܐ��X��ԓ��M���Ɩ�V>�����	+��1������s�������`n���ࣼ�R��Ħ�u5��q���c���������ci��ڰ��J��X���B,��7����������� d���ֽ��  �  �N=�M=�(M=|nL=��K=p�J=�<J=΀I=H�H=IH=�IG=��F=�E=�E=�MD=U�C=�B=�	B=GA=h�@=ʾ?=>�>=�2>=k==Z�<=��;=f;=A:=Ks9=-�8=��7=w7=�-6=NX5=�4=�3=�2=�1=�1=�/0=�K/=�e.=�|-=��,=U�+=/�*=��)=��(=��'=��&=;�%=��$=��#=��"=m�!=	� =Lp=R=O/=�=��=R�=t=�8=*�=]�=@g=�=��=�e=�=Ԟ=[3=��	=~L=3�=�P=H�=�@=�� =;�<�	�<���<���<TA�<���<���<�/�<^��<HT�<���<^�<p��<�P�<l��<%-�<
��<f��<�T�<���<	�<�W�<���<���<�>�<��<Cˢ<j�<�O�<g��<�͓<�
�<�F�<���<.��<O��<S`z<�r<Hk<�c<�2\<Y�T<�#M<�E<H><p�6<�"/<]�'<�7 <��<�^<��	<��<M��;o��;P�;Q��;.W�;���;���;�h�;A�;�^j;�iN;�2;M;�h�:V�:7>�:��+:���9���T���yu�󌭺P�ߺ"���C!��~9�_jQ��i�I&�������𖻴�����ⷻp�»�ͻ�Q׻Fwỹr�\D������G6�/��}z�����q����_��[#�`�'���+�խ/���3�ߖ7��u;�G?�ZC���F�dnJ�AN�+�Q��-U���X�0$\���_���b�
Rf��i���l��7p�vs�߭v���y�b}����Y���h7��&Ä��L��Qԇ��Y���݊��_��Q���I_���ܐ�$Y��ԓ��M���Ɩ�d>��6���'+��L��������������pn���ࣼ�R��Ħ�]5��r���T���������Vi���ٰ��J��P���/,��.���h��������c���ֽ��  �  �N=�M=�(M=snL=��K=y�J=�<J=̀I=>�H=CH=�IG=��F=�E=�E=�MD=D�C=��B=�	B=GA=_�@=��?==�>=�2>=k==[�<={�;=f;=	A:=Ws9=0�8=��7=~7=�-6=TX5=*�4="�3=�2=�1=�1=�/0=�K/=�e.=�|-=��,=W�+=(�*=�)=��(=��'=��&=/�%=��$=��#=��"=]�!=�� =Ap=	R=L/=�=��=H�=t=�8=)�=j�==g=�=��=�e=�=۞=l3=��	=�L==�=�P=[�=�@=�� =0;�<�	�<���<Ɍ�<fA�<���<}��<�/�<{��<:T�<���<r^�<`��<�P�<\��<-�<��<T��<iT�<���<��<�W�<���<l��<�>�<���<Lˢ<w�<�O�<i��<�͓<�
�<�F�<���<C��<V��<x`z<;�r<aHk<$�c<3\<i�T<�#M<O�E<V><��6<#/<a�'<�7 <��<_<`�	<�<���;>��;�O�;��;�V�;.��;o��;�g�;�@�;7^j;ViN;`�2;�;�h�:��:u?�:"�+:���97��i��.wu�����p�ߺѺ��C!��~9��iQ��i�&��}�����T������᷻�»�ͻ�Q׻�w�jr�gD������S6�`���z�����q������\#���'���+���/�ȩ3��7��u;�(G?�eC���F�wnJ�=N�1�Q�]-U���X�$\�H�_���b��Qf��i�U�l��7p�vs�ԭv�t�y�}����B���[7��*Ä��L��Sԇ��Y���݊��_��`���\_���ܐ�6Y��,ԓ�N���Ɩ��>��N���3+��^��������������|n���ࣼ�R��*Ħ�[5��n���:��
�������Ai���ٰ��J��;���,�����X��������c���ֽ��  �  �N=�M=�(M=|nL=��K=m�J=�<J=ÀI=9�H=8H=�IG=��F=��E=�E=�MD=;�C=��B=�	B=GA=U�@=��?=3�>=�2>=k==\�<=��;=n;=A:=Ys9==�8=��7=�7=�-6=dX5=5�4='�3=1�2=,�1=1=�/0=�K/=�e.= }-=��,=[�+=1�*=�)=��(=��'=��&=)�%=��$=��#=��"=U�!=� =2p= R=</=�=x�=C�=	t=�8=&�=e�=Fg=�=��=�e=�=�=t3=��	=�L=S�=�P=g�=�@=�� =X;�<
�<���<Ռ�<sA�<���<���<�/�<m��<9T�<���<e^�<O��<}P�<S��<�,�<ٓ�<1��<LT�<u��<��<�W�<���<_��<s>�<���<5ˢ<n�<�O�<s��<�͓<�
�<�F�<ρ�<Y��<z��<�`z<��r<}Hk<h�c<B3\<��T<�#M<p�E<�><��6<(#/<~�'<�7 <��<�^<X�	<Ǜ<ʆ�;���;WO�;���;jV�;��;���;�g�;?@�;�]j;MhN;��2;�;�f�:Q�:�=�:��+:���9	�����Hwu�r���A�ߺ����B!��}9��hQ�xi��%�����?�0��U���᷻�»�ͻ�Q׻Awờr뻟D�����}6�}���z����r������G\#�ʇ'�ߢ+��/��3�'�7�v;�DG?�xC���F�\nJ�3N��Q�P-U���X��#\�5�_���b��Qf���i�;�l�m7p��us���v�2�y�}����<���T7��Ä��L��Nԇ��Y���݊��_��p���o_��
ݐ�@Y��Kԓ�"N���Ɩ��>��a���N+��x���������������n���ࣼ�R��Ħ�P5��a���7����������,i���ٰ�iJ������+������;��������c��wֽ��  �  ��N=!�M=�(M=znL=��K=i�J=�<J=��I=4�H=.H=�IG=��F=��E=�E=�MD=3�C=��B=�	B=�FA=M�@=��?=(�>=�2>=
k==Z�<=�;=n;=A:=^s9=M�8=��7=�7=�-6=sX5=E�4=9�3=D�2=3�1=1=�/0=�K/=�e.=}-=��,=Y�+=/�*=��)=��(=��'=��&=&�%=��$=��#=w�"=K�!=�� =%p=�Q=*/=�=l�=?�=�s=�8=*�=_�=Gg=�=��=�e==��=�3=��	=�L=h�=�P=z�=A=�� =w;�<(
�<���<��<�A�<���<���<�/�<c��<DT�<t��<X^�<D��<eP�<:��<�,�<ʓ�<��<9T�<T��<��<�W�<���<X��<X>�<�<1ˢ<c�<�O�<k��<�͓<�
�<�F�<遈<n��<���<�`z<��r<�Hk<��c<u3\<�T<"$M<��E<�><��6<N#/<u�'<�7 <��<�^<X�	<��<���;���;�N�;��;�U�;i�;7��;Mg�;�?�;�\j;]gN;�2;i;5e�::�:�<�:q�+:뼃9������vu�Չ���ߺn��`B!��|9�hQ�}i�%��ԟ���������w᷻�»�ͻ�Q׻Zw��r뻢D��J����6����{�
 �\r��� �}\#��'�,�+�D�/�;�3�<�7�Bv;�eG?�qC���F�`nJ�;N���Q�8-U�c�X��#\��_�`�b��Qf�r�i���l�/7p�us�h�v��y��
}����3���E7��Ä��L��Pԇ��Y���݊��_������|_��$ݐ�[Y��sԓ�3N�� ǖ��>������p+������������������n���ࣼ�R��Ħ�W5��O���/��އ��z���i���ٰ�TJ�������+��Ӝ��$�����}񺼲c��\ֽ��  �  �N=!�M=�(M=}nL=��K=l�J=�<J=��I=&�H=!H=�IG=��F=��E=�E=�MD=!�C=��B=�	B=�FA=@�@=��?=$�>=�2>=k==]�<=��;=o;=A:=ks9=O�8=��7=�7=�-6=�X5=P�4=G�3=L�2=G�1=$1=�/0=�K/=�e.=}-=��,=`�+=0�*=��)=��(=��'=��&=�%=��$=��#=o�"=;�!=҉ =p=�Q=$/=�=c�=1�=�s=�8=%�=d�=Jg=�=��=�e==�=�3=��	=�L=s�=Q=��=A=ӱ =�;�<I
�<���<��<�A�<���<���<�/�<l��<4T�<n��<H^�<*��<RP�<��<�,�<���<���<T�<8��<��<�W�<k��<8��<N>�<ᅦ<1ˢ<h�<�O�<x��<�͓<�
�<�F�<���<���<���<1az<��r<�Hk<Խc<�3\<.�T<P$M<ԟE<�><��6<O#/<��'<�7 <��<�^<5�	<}�<)��;��;�N�;���;^U�;��;���;�f�;+?�;�[j;�fN;�2;�;Fd�:��:�<�:��+:���9���D��.tu�щ����ߺ��lA!�!|9��gQ��i��$��C���u������6᷻��»�ͻ�Q׻Yw��r��D�������6����1{�> �r�\��K ��\#�2�'�I�+�~�/�g�3�~�7�^v;�G?��C���F�]nJ�N��Q�-U�4�X��#\�֐_�3�b�BQf�R�i���l��6p�Ous� �v���y��
}�������77��Ä��L��Kԇ��Y���݊��_�������_��:ݐ�zY���ԓ�YN��"ǖ��>�������+������	��Ɉ�������n���ࣼ�R��Ħ�J5��S�����҇��i����h���ٰ�-J��庳��+��Ĝ��������h񺼞c��Qֽ��  �  �N="�M=)M=~nL=��K=e�J=�<J=��I=�H=H=�IG=r�F=��E=�E=�MD=�C=��B=�	B=�FA=7�@=��?="�>=�2>=	k==S�<=��;=y;=A:=vs9=V�8=��7=�7=�-6=�X5=_�4=X�3=U�2=X�1=)1=�/0=L/=�e.=}-=��,=i�+=-�*=��)=��(=��'=��&=�%=��$=~�#=^�"=+�!=ʉ =p=�Q=/=�=`�='�=�s=�8= �=c�=Fg=�=�=�e==�=�3=��	=�L=�=Q=��=)A=� =�;�<k
�<��<!��<�A�<��<���<�/�<h��<-T�<l��<;^�<��<FP�<���<�,�<���<���<�S�<��<��<�W�<`��<��<J>�<օ�<"ˢ<W�<�O�<���<�͓<�
�<�F�<��<���<���<baz<�r<WIk<�c<�3\<V�T<�$M<�E<�><'�6<Y#/<��'<�7 <��<�^<�	<w�<ǅ�;���;/N�;&��;�T�;O�;k��;f�;�>�;]Zj;�eN;+�2;�;�c�:��:�;�:N�+:���9���9���qu�D�����ߺW���@!��{9��fQ�� i��$��ɞ��Q��{���෻p�»�ͻJQ׻|w��r�E�������6���?{�� ��r����n ��\#�}�'���+�Ʈ/�z�3���7�pv;��G?��C���F�vnJ�N��Q��,U��X��#\���_��b��Pf�.�i���l��6p�(us��v���y�w
}�{�����/7��Ä��L��]ԇ��Y���݊�`�������_��Gݐ��Y���ԓ�|N��-ǖ��>�������+��������∟������n���ࣼ�R��Ħ�35��O�����Ƈ��T����h��zٰ�J��к���+���������o��L񺼉c��Gֽ��  �  �N=+�M=�(M={nL=��K=e�J=�<J=��I=�H=H=�IG=o�F=��E=~E=�MD=�C=��B=�	B=�FA=-�@=��?=�>=�2>=k==[�<=��;=u;="A:=ws9=a�8=��7=�7= .6=�X5=m�4=b�3=f�2=^�1=21=�/0=L/=�e.=}-=��,=]�+=/�*=��)=��(=��'=��&=�%=��$=y�#=Z�"=%�!=�� =�o=�Q=/=�=Q�=$�=�s=�8=#�=d�=Lg=�=�=�e='=�=�3=��	=�L=��='Q=��=;A=� =�;�<x
�<.��<)��<�A�<��<���<�/�<h��<0T�<W��<3^�<��</P�<���<�,�<t��<���<�S�<��<��<zW�<@��<��<1>�<˅�<!ˢ<e�<�O�<w��<�͓<�
�<�F�< ��<���<���<�az<b�r<zIk<L�c<#4\<z�T<�$M<�E<><,�6<#/<��'<�7 <��<�^<
�	<D�<���;n��;�M�;��;�T�;��;ɡ�;�e�;Q>�;Zj; eN;r�2;d;�a�:&�:);�:��+:���9f��x��)ru����7�ߺ��j@!��z9��eQ�> i�*$���������5���෻g�»iͻ�Q׻pw��r� E������7����{�� ��r����� �,]#���'���+�Ԯ/���3���7��v;��G?��C���F�gnJ�-N��Q��,U���X�V#\���_���b��Pf��i�U�l��6p��ts�Ҭv���y�f
}�c������)7��Ä��L��Oԇ� Z���݊�`�������_��_ݐ��Y���ԓ��N��Tǖ�?��˵���+��͠��2��鈟�����n���ࣼ�R��Ħ�J5��=���������D����h��hٰ�J�������+���������_��;�}c��2ֽ��  �  �N=4�M=�(M=�nL=��K=[�J=�<J=��I=�H=H=}IG=b�F=��E=yE=�MD=�C=��B=�	B=�FA=(�@=��?=�>=�2>=�j==`�<=��;=|;=)A:=xs9=i�8=��7=�7=.6=�X5=t�4=h�3=p�2=f�1=H1=�/0=L/=�e.=}-=��,=a�+=8�*=�)=��(=��'=��&=�%=��$=s�#=K�"=�!=�� =�o=�Q=/=�=H�=$�=�s=�8= �=Z�=Vg=�=�=�e=/=!�=�3=��	=�L=��=0Q=��=IA=�� =�;�<�
�<>��<1��<�A�<*��<���<�/�<Q��<1T�<N��<-^�<��<P�<���<{,�<j��<���<�S�<�<e�<nW�<0��<��< >�<ȅ�<ˢ<\�<�O�<{��<�͓<�
�<�F�<%��<Ƽ�< ��<�az<��r<�Ik<m�c<M4\<īT<�$M<)�E<D><(�6<�#/<��'<8 <��<�^<�	<"�<���;3��;�M�;���;%T�;��;o��;�e�;�=�;+Yj;odN;	�2;$;�`�:	�:x9�:��+:���9�����Xru�P����ߺ���?!�7z9��eQ���h��#��l���k���*���෻l�»$ͻ�Q׻.w�:s�1E������"7����{�� �s����� �I]#���'��+���/��3���7��v;��G?��C�,�F�BnJ�N���Q��,U��X�F#\�w�_���b��Pf���i�;�l�q6p��ts���v�H�y�Y
}�W������7�����L��@ԇ�Z���݊�(`�������_��qݐ��Y���ԓ��N��hǖ�?��浙��+��ؠ��A��戟�����n���ࣼ�R��	Ħ�E5��,���������@����h��@ٰ��I������{+��|������;��%�xc��!ֽ��  �  �N=0�M=)M=}nL=��K=_�J=�<J=��I=�H=H=zIG=^�F=��E=rE=�MD=��C=��B=�	B=�FA=#�@=��?=�>=�2>=�j==Y�<=��;=|;=(A:=�s9=o�8=��7=�7=.6=�X5=z�4=t�3=r�2=h�1=?1=�/0=L/=�e.= }-=��,=b�+=2�*=��)=��(=��'=��&=��%=��$=o�#=I�"=�!=�� =�o=�Q=�.=�=K�=�=�s=�8=$�=`�=Pg=�=�=�e=5=(�=�3=��	=�L=��=<Q=��=JA=�� =�;�<�
�<K��<E��<�A�<)��<���<�/�<^��<6T�<Q��< ^�<���<"P�<���<|,�<[��<���<�S�<譼<_�<dW�<0��<��<!>�<ʅ�<ˢ<V�<�O�<���<�͓<�
�<G�<5��<ʼ�<���<�az<��r<�Ik<�c<T4\<��T<�$M<N�E<\><K�6<�#/<��'<�7 <��<�^<�	< �<T��;!��;�M�;p��;T�;m�;c��;;e�;�=�;�Xj;ZdN;��2;�;�`�:#�:�9�:��+:ۺ�9Y��p��pu�������ߺ8���?!�@z9�-eQ�.�h��#��Y����������r෻=�»?ͻ�Q׻bw�&s�E������)7�9���{�� � s���� �W]#�؈'��+��/�ת3��7��v;��G?��C��F�]nJ�N�ĢQ��,U�ϬX�-#\�X�_���b��Pf���i��l�K6p��ts���v�W�y�5
}�K��騁�7�����L��Qԇ�Z���݊�%`�������_��oݐ��Y���ԓ��N��iǖ�?����+��⠜�B����������n���ࣼ�R��Ħ�?5��1����������1����h��Rٰ��I������b+��s������J��$�gc��ֽ��  �  ��N=��M=�"M=�gL=��K=��J=k3J=�vI=!�H=6�G=�<G=�}F=6�E=��D==D=�{C=3�B=�A='2A=Wm@=��?=��>=+>=gP==t�<=M�;=��:=2!:= R9=��8=��7=��6=�6=�/5=�V4=;|3=��2=��1=��0=��/=*/=/.=�D-=2W,=g+=
t*=�})=��(='�'=;�&=��%=�}$=�r#=�c"=Q!=: =�=-�=�=X�=�=�R=�={�=K�=X=�=�=f=�
=s�=�D=��
=�i	=��=`z=�=�v=��=` =I��<lm�<�6�<���<��<�`�<�	�<��<5E�<���<se�<��<�l�<���<7]�<���<|9�<���<��<�b�<齸<��<Oj�<໭<�
�<�V�<���<��<�.�<=s�<��<���<O8�<x�<0��<���<�hz<%�r<Sbk<��c<�^\<�T<aM<l�E<Bl><8�6<{�/<�(<� <D<�<i�
<2<���;�4�;Ʋ�;@�;�޽;���;qQ�;�'�;�;�'n;oWR;ȶ6;�H;� ;��:J~�:�>:�Ϫ9�d��,|��	�`��٢���Ժ].�C����3���K�9)c��cz�⥈���������ܴ�|���c�ɻ�OԻ�x޻�x�7P�S���M���s�������-x�C��$"�;A&�Ec*��u.��x2�(m6�US:�3,>���A��E�jI�xM�ԭP��?T��W��D[�p�^�%b��e�S�h��6l���o���r�v�P>y��p|���+b��E�����h������!������,������0��s����.��%���(��𢖼���^���=��:���h����o���䠼5Y��
ͣ�m@������O&��ߘ��*��]}��aﭼpa��qӰ��E��÷���)������B��A�������ki���ݽ��  �  ��N=��M=�"M=�gL=��K=��J=q3J=vI=�H=;�G=�<G=�}F=4�E=��D==D=�{C=2�B=�A=/2A=[m@=��?=��>=3>=bP==r�<=O�;=��:=9!:="R9=��8=��7=��6=�6=�/5=�V4=4|3=��2=��1=��0=��/='/=/.=�D-=7W,=g+=t*=�})=��(=$�'=,�&=��%=�}$=�r#=�c"=Q!=: =�=/�=�=`�=�=�R=�=u�=P�=X=�=�=f=�
=u�=�D=��
=�i	=��=_z=�=�v=��=` =?��<hm�<�6�<���<&��<�`�<�	�<��<&E�<���<ae�<���<�l�<���<F]�<���<�9�<���<��<�b�<�<��<Uj�<໭<�
�<W�<���<��<�.�<Bs�<%��<���<W8�<x�<)��<���<ihz<0�r<7bk<��c<�^\<��T<aM<_�E<Kl><:�6<��/<�(<� <�C<��<��
<�1<n��;�4�;��;�@�;�޽;���;�Q�;�'�;�;0(n;�WR;�6;hH;  ;��:�}�:��>:�Ъ9�`���x��k�`�0٢���Ժ�.�2���3���K��)c�xcz�N������������۴�\���>�ɻ�OԻ�x޻�x� P�d�������s��������)x����"�2A&�9c*�iu.��x2�$m6��S:�H,>���A��E��iI�qM�ĭP�z?T��W��D[�n�^�%b�R�e�R�h��6l���o���r�Pv�b>y��p|���%b��8�����d������!��|���0,��)����0��i����.��&���(��⢖����c���3��%���b����o���䠼.Y��	ͣ�z@������J&��Ϙ��%��V}��hﭼwa���Ӱ��E������*������L��U�������pi���ݽ��  �  ��N=��M=�"M=�gL=��K=��J=|3J=�vI=)�H=7�G=�<G=�}F=4�E=�D==D=�{C=4�B=�A=&2A=]m@=��?=��>=;>=`P==t�<=M�;=��:=6!:=R9=��8=��7=��6=�6=�/5=�V4=-|3=��2=��1=��0=��/=!/=/.=�D-=4W,=g+=t*=�})=��(=.�'=4�&=��%=�}$=�r#=�c"=Q!=: =�=0�=�=^�=�=�R=�=~�=T�=X=�=�=f=�
=q�=�D=��
=�i	=��=cz=�=�v=��=` =B��<^m�<�6�<���<��<�`�<}	�<��<E�<���<qe�<��<�l�<���<H]�<���<�9�<���<��<�b�<���<��<Ij�<���<�
�<W�< ��<��<�.�<7s�<"��<���<R8�<x�<'��<���<ehz<7�r<bk<��c<�^\<��T<�`M<K�E<@l><�6<��/<�(<� <�C<��<��
<�1<���;�4�;��;�@�;�޽;��;�Q�;(�;�;F(n;nWR;J�6;"I;� ;�:�}�:U�>:�Ъ9jg���y���`��٢�%�Ժ�.�����3�ٟK�*c�cz�O�����������ܴ�����S�ɻ�OԻ�x޻�x�P����h��s���Ț�w�"x����"�.A&�,c*�qu.��x2��l6�uS:�#,>���A��E��iI��M�ЭP��?T�$�W��D[�u�^�%b�T�e�?�h��6l�˂o���r�Nv�X>y��p|�-��1b��>�����h������!��m���,�����0��y����.��"���(��碖����b���.��0���n����o���䠼Y��ͣ�{@������U&��Ҙ��3��Z}��tﭼza���Ӱ��E������*������M��T�������yi���ݽ��  �  ��N=��M=�"M=�gL=��K=��J=s3J=�vI=%�H=@�G=�<G=�}F=B�E=�D=$=D=�{C=A�B=&�A=12A=`m@=��?=��>=0>=gP==s�<=K�;=��:=3!:=R9=��8=��7=��6=�6=�/5=�V4=-|3=z�2=��1=��0=��/= /=/.=D-=5W,=g+=t*=�})=��(=*�'=7�&=��%=�}$=�r#=�c"=Q!=: =�=;�=�=d�=��=�R=�=|�=I�=X=�=�=f=�
=o�=�D=��
=�i	=��=Mz=
�=�v=��=�_ ="��<Rm�<�6�<���<��<�`�<z	�<��</E�<���<te�<��<�l�<���<W]�<���<�9�<ʠ�<��<�b�<��<��<_j�<�<�
�<W�<���<��<�.�<As�<��<���<N8�<	x�<��<���<<hz<��r<bk<��c<q^\<��T<�`M<B�E<5l><&�6<��/<�(<�� <	D<�<��
<2<���;5�;3��;A�;b߽;P��;�Q�;j(�;��;�(n;7XR;��6;I;� ;��:�~�:^�>:\Ъ9M[��z���`��٢�v�Ժ=/�H����3�@�K��)c�Edz�r����*�����ܴ�����B�ɻ�OԻ�x޻�x�;P�4���X���s������M��w����"��@&��b*�Uu.�x2�m6�gS:�(,>���A��E�jI�qM�ɭP��?T�#�W��D[���^�G%b�`�e���h��6l��o��r�]v��>y��p|�1��/b��D��i������!������,�����~0��`����.������'��Ԣ�����H����� ���Y����o���䠼'Y��
ͣ�m@������L&��ט��/��_}��wﭼ�a���Ӱ��E��ط��*������g��e�������}i���ݽ��  �  ��N=��M=�"M=�gL=��K=��J=w3J=�vI=(�H=N�G=�<G=�}F=E�E=�D=0=D=�{C=D�B=%�A=<2A=mm@=��?=��>=6>=nP==o�<=L�;=��:=(!:=R9=��8=��7=��6=�6=�/5=�V4=$|3=r�2=��1=��0=��/=/=/.=zD-=*W,=g+=t*=�})=��(=1�'==�&=��%=�}$=�r#=�c"=Q!=: =�=?�= �=f�=�=�R=�=��=N�=X=�=�=�e=�
=e�=�D=��
=�i	=��=Ez=�=�v=��=�_ =��<Fm�<�6�<w��<���<�`�<y	�<٪�<:E�<���<�e�<��<�l�<���<T]�<���<�9�<��<��<�b�<��<��<}j�<���<�
�<W�<
��<��<�.�<?s�<��<���<68�<�w�<
��<���<Dhz<��r<�ak<��c<s^\<��T<�`M<$�E<�k><�6<O�/<�(<� <D<�<��
<)2<���;�5�;u��;A�;�߽;���;OR�;�(�;��;	)n; YR;v�6;fI; ;��:��: �>:�Ѫ9�a���~����`��ڢ���Ժ�/�_����3���K�p*c��dz�_���2�T��3��Kܴ�������ɻ�OԻ�x޻dx�P�����=��|s�Q����F��w�����"��@&��b*�Ku.�Kx2��l6�RS:�,>���A�ͶE�jI�oM��P��?T�D�W�'E[���^�e%b�a�e���h��6l��o��r�dv��>y��p|�]��<b��X�����f������� ��x���
,�����g0��G����.������'������}��?��������<����o���䠼Y���̣�n@������O&��𘩼7��v}���ﭼ�a���Ӱ��E��鷳�-*������e��l��������i���ݽ��  �  ~�N=��M=�"M=�gL=��K=��J=|3J=�vI=8�H=L�G=�<G=�}F=Q�E=�D=2=D=�{C=Q�B=8�A=<2A=rm@=��?=��>==>=gP==r�<=K�;=��:=,!:=R9=��8=~�7=��6=�6=�/5=�V4=|3=q�2=��1=��0=��/=/=/.=yD-=*W,=g+=
t*=�})=��(=3�'=B�&=Є%=�}$=�r#=�c"=!Q!=%: =�=I�=/�=u�=��=�R=�=��=U�=X=�=�=�e=�
=`�=�D=��
=�i	=��=Az=��=�v=��=�_ =���<+m�<�6�<h��< ��<�`�<o	�<ݪ�<&E�<���<|e�<!��<�l�<���<x]�<��<�9�<��<��<�b�<4��<��<sj�<��<�
�<W�<��<��<�.�<2s�<��<���<28�<�w�<���<���<�gz<��r<�ak<t�c<8^\<t�T<�`M<��E<�k><�6<]�/<�(<�� <D<�<��
<%2<J��;�5�;���;�A�;�߽;���;oR�;)�;'�;S*n;!YR;�6;=J;} ;��:%�:/�>:YҪ94g���{����`�3ۢ���Ժ�/�b��D�3�J�K�]+c��dz����~򓻬��Q��^ܴ�������ɻ�OԻ�x޻�x��O�����(��9s�l�a����w�����"��@&��b*�u.�ex2��l6�6S:�,>���A���E�jI��M���P��?T�R�W�9E[�Ϲ^��%b���e���h�.7l�2�o�)�r��v��>y��p|�o��Fb��Q����l������!��i���,������T0��M����.��㫓��'������e��%���������F����o���䠼Y���̣�r@������\&��阩�=��{}���ﭼ�a���Ӱ��E��񷳼Q*��Ü��������������i���ݽ��  �  o�N=��M=�"M=�gL=��K=��J=�3J=�vI=>�H=T�G=�<G=�}F=U�E=*�D=@=D=�{C=Q�B=A�A=H2A=zm@=��?=��>=G>=gP==w�<=H�;=��:=)!:=R9=��8=n�7=��6=�6=�/5=�V4=
|3=e�2=��1=��0=��/=/=/.=mD-=-W,=
g+=t*=�})=��(=7�'=C�&=ل%=�}$=�r#=�c"=+Q!=2: =�=U�=-�=��=�=�R=�=��=[�=X=�=ڻ=�e=�
=R�=�D=��
=�i	=p�=1z=��=�v=��=�_ =��<m�<�6�<J��<��<�`�<c	�<��<!E�<���<~e�<'��<�l�<���<�]�<���<�9�<��<
�<�b�<:��<�<�j�<)��<�
�<.W�<��<��<�.�<)s�<��<���<(8�<�w�<䶄<���<�gz<��r<zak<U�c<�]\<\�T<v`M<��E<�k><��6<[�/<}(<�� <D<"�<ч
<,2<���;�5�; ��;�A�;�;���;�R�;�)�;6�;+n;�YR;��6;�J;� ;b�:x�:�>:�Ѫ9�c���|��چ`��ڢ���Ժ0����:�3���K��+c�Rez�z���|���_���ܴ����m�ɻ�OԻ�x޻�x軔O����!��s�@�*����w����d"��@&��b*��t.�?x2��l6�.S:��+>���A���E��iI��M��P��?T�~�W�;E[�
�^��%b���e���h�W7l�S�o�g�r��v��>y�%q|�i��`b��]����u������!��V���,������E0��7����.��竓��'������I��������ボ�4����o���䠼Y���̣�q@������f&��嘩�[���}���ﭼ�a���Ӱ��E�����e*��ќ��������������i���ݽ��  �  m�N=��M=�"M=�gL=��K=��J=�3J=�vI=?�H=a�G=�<G=�}F=g�E=1�D=J=D=�{C=b�B=C�A=Q2A=�m@=��?=
�>=D>=mP==t�<=H�;=��:=!!:=R9=�8=d�7=��6=�6=�/5=�V4=�{3=W�2=��1=��0=��/=/=/.=kD-=$W,=g+=t*=�})=��(==�'=O�&=ք%=�}$=�r#=d"=9Q!=9: =�=b�=:�=��=�=�R=�=��=V�=X=�=ٻ=�e=�
=M�=�D=��
=�i	=o�=!z=��=�v=��=�_ =Қ�<�l�<q6�<C��<��<`�<a	�<ڪ�<)E�<���<�e�<7��<�l�<���<�]�<��<�9�<��<�<c�<N��<�<�j�<)��<�
�<3W�<��<��<�.�<'s�<���<���<8�<�w�<ʶ�<~��<�gz<`�r<@ak<�c<�]\<<�T<8`M<��E<�k><��6<2�/<s(<� <D<-�<ԇ
<j2<���;66�;Z��;)B�;��;�;FS�;�)�;��;D+n;�ZR;�6;BK;� ;R�:]��:߻>:Ӫ9�f��S����`��ۢ���Ժ�0������3�`�K��,c�fz�^�����L������ܴ������ɻ�OԻ�x޻px軞O�~������s� �$����Dw�]��<"�S@&�}b*��t.�x2��l6�S:��+>���A�߶E�jI��M��P��?T���W�ZE[�/�^��%b��e��h��7l���o���r��v�
?y�Nq|����bb��g�
���s������� ��]����+��⮍�=0�� ����.��ǫ���'������=���������ك������o���䠼 Y���̣�l@������h&������_���}���ﭼ�a���Ӱ��E������*��������������i���ݽ��  �  n�N=��M=�"M=�gL=��K=��J=�3J=�vI=B�H=k�G=�<G=~F=s�E=8�D=\=D=�{C=v�B=Q�A=\2A=�m@=ç?=�>=A>=tP==o�<=L�;=��:=!:=R9=o�8=j�7=��6=w6=v/5=�V4=�{3=L�2=��1=��0=��/=�/=�..=kD-=W,=g+=t*=�})=��(=:�'=T�&=ۄ%=�}$=�r#=d"=<Q!=E: =	=c�=P�=��=�=�R=�=��=W�=X=�=�=�e=�
=D�=�D=��
=�i	=]�=z=��=�v=��=�_ =���<�l�<L6�<8��<ٯ�<o`�<h	�<ʪ�<5E�<���<�e�<;��<�l�<���<�]�<F��<�9�<7��<*�<)c�<p��<"�<�j�<1��<�<,W�<'��<��<�.�<3s�<�<���<8�<�w�<Ƕ�<X��<xgz<-�r<3ak<��c<�]\<��T<'`M<��E<�k><��6<�/<|(<� <D<F�<ć
<|2<���;�6�;���;�B�;�;��;�S�;*�;w�;;,n;�[R;��6;�K; ;A�:���:�>:�ժ9Vj�����h�`�]ݢ���Ժc1���J�3�
�K��,c��fz�ԧ��T�)������ܴ������ɻ�OԻ�x޻Lx軇O�������s�����w�7w�*��"�J@&�#b*��t.��w2��l6��R:��+>���A�ȶE�jI�tM�'�P��?T���W��E[��^��%b�-�e�E�h��7l���o���r�*v�>?y�2q|�͝�hb��k����g����� ��_����+��ܮ��30��
����.�������'��e���)��甙����σ������o���䠼Y���̣�l@������\&�����Z���}���ﭼ�a���Ӱ�F��7����*��������Ƃ������i��޽��  �  g�N=��M=�"M=�gL=��K=��J=�3J=�vI=O�H=q�G==G=~F=r�E=A�D=e=D=�{C=s�B=U�A=b2A=�m@=ͧ?=�>=N>=uP==r�<=K�;=��:=!:=�Q9=l�8=\�7=��6=u6=r/5=�V4=�{3=F�2=��1=��0=x�/=�/=�..=cD-=W,=g+=t*=�})=Ȅ(=C�'=Z�&=�%=�}$=�r#=d"=?Q!=M: ==h�=O�=��= �=�R=�=��=_�=	X=�=ڻ=�e=�
=>�=�D=��
=�i	=Y�=z=��=�v=��=�_ =���<�l�<C6�<%��<Ư�<^`�<a	�<Ϊ�<2E�<���<�e�<L��<m�<	��<�]�<A��< :�<I��<;�<)c�<w��<4�<�j�<I��<�<DW�<.��<��<�.�<$s�<浓<���<�7�<�w�<���<W��<kgz<�r<ak<��c<�]\<��T<`M<k�E<zk><��6<�/<](<� <D<N�<�
<�2<��;�6�;ٴ�;�B�;�;Y��;0T�;[*�;n�;�,n;�[R;A�6;VL;w ; �:Ӂ�:-�>:>֪9	t��_���
�`��ݢ�4�Ժ�1����~�3�}�K��-c�	gz�ᧈ�D󓻉��3��ݴ�C����ɻ�OԻ�x޻Sx�BO�G�������r�����q�(w�	���"�5@&�!b*��t.��w2�Ql6��R:��+>��A�̶E�jI��M�?�P� @T���W��E[�K�^��%b�7�e�X�h��7l�փo���r�0v�R?y�dq|�֝�wb��z�$���k������� ��H����+��ɮ��0������{.�������'��T�����攙�������������o���䠼�X���̣�n@������k&�����j���}���ﭼ�a���Ӱ�F��C����*��������ǂ��%����i��޽��  �  b�N=��M=�"M=�gL= �K=��J=�3J=�vI=R�H=s�G==G=~F=��E=L�D=c=D=�{C=|�B=`�A=j2A=�m@=ϧ?=�>=O>=pP==w�<=C�;=��:=!:=�Q9=q�8=P�7=��6=k6=e/5=�V4=�{3=;�2=}�1=��0=k�/=�/=�..=bD-="W,=g+=t*=�})=ń(=F�'=Y�&=�%=�}$=�r#=d"=RQ!=Q: ==|�=Q�=��=$�=�R=�=��=\�=X=�=λ=�e=�
=9�=�D=��
=�i	=K�= z=��=�v=r�=�_ =���<�l�<H6�<��<ί�<h`�<K	�<ت�<&E�<���<�e�<L��<m�<��<�]�<N��<':�<G��<L�<Lc�<���<L�<�j�<M��<�<JW�<&��<��<�.�<s�<���<x��<8�<�w�<���<B��<4gz<��r<�`k<��c<d]\<��T<�_M<N�E<�k><��6<-�/<Q(<� <D<>�<�
<�2<+��;�6�;-��;C�;��;���;*T�;�*�;��;\-n;�\R;m�6;�L;s ;\�:b��:ܽ>:�Ҫ9�k��A~��߈`��ܢ���Ժ%2����A�3�ȣK�.c��gz�E���~����+��ݴ�H�����ɻPԻzx޻Vx�ZO�*�������r������e��v�����"��?&�b*�`t.��w2�Nl6��R:��+>���A�׶E��iI��M��P��?T���W��E[���^�&b�h�e���h��7l��o��r�Vv�n?y��q|�ǝ�b��o����������� ��I����+��Ǯ��0��﯐�c.������m'��U�����Ô��������������o���䠼�X���̣�h@������v&������r���}���ﭼ b��	԰�,F��U����*��#������݂��8����i�� ޽��  �  Z�N=��M=�"M=�gL=�K= �J=�3J=�vI=U�H=w�G==G=~F=��E=M�D=l=D=�{C=}�B=`�A=j2A=�m@=ѧ?=�>=Q>=uP==x�<=C�;=��:=!:=�Q9=c�8=W�7=��6=h6=d/5=�V4=�{3=:�2=z�1=��0=s�/=�/=�..=YD-=W,=g+=
t*=�})=Ǆ(=I�'=^�&=�%=�}$=�r#=d"=NQ!=U: ==w�=Q�=��='�=�R=�=��=^�=X=�=л=�e=�
=0�=�D=��
=�i	=G�=�y=��=v=p�=�_ =���<�l�<-6�<	��<���<b`�<K	�<ת�<1E�<���<�e�<Q��<m�<��<�]�<O��<:�<V��<Q�<Ic�<��<J�<�j�<W��<�<NW�</��<��<�.�<s�<鵓<f��<�7�<�w�<���<@��<.gz<��r<�`k<��c<b]\<��T<�_M<T�E<Zk><e�6<�/<T(<� <D<T�<�
<�2<F��;�6�;3��;C�;��;đ�;xT�;�*�;��;Z-n;�\R;ۻ6;�L;� ;��:-��:
�>:#Ӫ92n��<�����`��ޢ���Ժ�1����F�3�ۣK��-c��gz�V����󓻫��S��]ݴ�������ɻ�OԻ�x޻@x�CO��������r������c��v�����"��?&�b*�gt.��w2�9l6��R:��+>�{�A�ʶE��iI��M�(�P�#@T���W��E[�e�^�&b�s�e���h��7l��o�	�r�gv�]?y�q|�����b�������~������� ��D����+��®��0��﯐�c.������y'��E�����ǔ��������������o��{䠼�X���̣�e@������s&���������}���ﭼ�a��
԰�.F��\����*��*������߂��*����i��޽��  �  g�N=��M=�"M=�gL=��K=��J=�3J=�vI=S�H=z�G==G=~F=��E=M�D=s=D=�{C=��B=g�A=m2A=�m@=Χ?=�>=J>=tP==u�<=K�;=��:=!:=�Q9=c�8=U�7=��6=b6=f/5=�V4=�{3=7�2={�1=��0=o�/=�/=�..=`D-=W,=g+=	t*=�})=Ą(=C�'=[�&=�%=�}$=�r#=-d"=PQ!=[: ==x�=a�=��=&�=�R=�=��=Z�=X=�=ֻ=�e=�
=@�=�D=��
=�i	=E�=�y=��=uv=p�=�_ =���<�l�<*6�<'��<���<]`�<Z	�<Ъ�<.E�<���<�e�<J��<m�<��<�]�<g��<:�<f��<U�<Pc�<���<U�<�j�<S��<�<AW�<-��<��<�.�<&s�<۵�<~��<�7�<�w�<���<2��<3gz<��r<�`k<y�c<h]\<��T<�_M<?�E<kk><��6<�/<^(<�� <D<G�<�
<�2<7��;7�;^��;_C�;��;���;�T�;�*�;�;�-n;�\R;!�6;�L;� ;��:��:a�>:2ת9n��-�����`�}ޢ���Ժw2�
��!�3�]�K�U.c��gz�S��������g���ܴ�T���#�ɻ�OԻ�x޻Rx�^O�B�������r������ ��v�����"��?&��a*�Tt.��w2�6l6��R:��+>���A�ҶE� jI��M�B�P�@T���W��E[�l�^�7&b�z�e���h�8l��o��r��v��?y��q|����pb���� ���n������� ��O����+��Ȯ��	0����W.��y���'��6����������������������o��~䠼�X���̣�i@������i&�����l���}���ﭼ�a��԰�,F��f����*��9������ꂹ�=����i��޽��  �  Z�N=��M=�"M=�gL=�K= �J=�3J=�vI=U�H=w�G==G=~F=��E=M�D=l=D=�{C=}�B=`�A=j2A=�m@=ѧ?=�>=Q>=uP==x�<=C�;=��:=!:=�Q9=c�8=W�7=��6=h6=d/5=�V4=�{3=:�2=z�1=��0=s�/=�/=�..=YD-=W,=g+=
t*=�})=Ǆ(=I�'=^�&=�%=�}$=�r#=d"=NQ!=U: ==w�=Q�=��='�=�R=�=��=^�=X=�=л=�e=�
=0�=�D=��
=�i	=G�=�y=��=v=p�=�_ =���<�l�<-6�<
��<���<b`�<L	�<ت�<1E�<���<�e�<Q��<m�<��<�]�<O��<:�<V��<Q�<Hc�<��<I�<�j�<V��<�<NW�</��<��<�.�<s�<鵓<f��<�7�<�w�<���<@��<.gz<��r<�`k<��c<b]\<��T<�_M<U�E<Zk><e�6<�/<U(<� <D<U�<�
<�2<G��;�6�;4��;C�;��;đ�;xT�;�*�;��;W-n;�\R;ػ6;�L;� ;��:$��:��>:�Ҫ9�n��f�����`��ޢ���Ժ�1����K�3��K��-c��gz�X����󓻬��U��_ݴ�������ɻ�OԻ�x޻Ax�DO��������r������c��v�����"��?&�b*�gt.��w2�9l6��R:��+>�{�A�ʶE��iI��M�(�P�#@T���W��E[�e�^�&b�s�e���h��7l��o�	�r�gv�]?y�q|�����b�������~������� ��D����+��®��0��﯐�c.������y'��E�����ǔ��������������o��{䠼�X���̣�e@������s&���������}���ﭼ�a��
԰�.F��\����*��*������߂��*����i��޽��  �  b�N=��M=�"M=�gL= �K=��J=�3J=�vI=R�H=s�G==G=~F=��E=L�D=c=D=�{C=|�B=`�A=j2A=�m@=ϧ?=�>=O>=pP==w�<=C�;=��:=!:=�Q9=q�8=P�7=��6=k6=e/5=�V4=�{3=;�2=}�1=��0=k�/=�/=�..=bD-="W,=g+=t*=�})=ń(=F�'=Y�&=�%=�}$=�r#=d"=RQ!=R: ==|�=Q�=��=$�=�R=�=��=\�=X=�=λ=�e=�
=:�=�D=��
=�i	=K�= z=��=�v=r�=�_ =���<�l�<I6�<��<ϯ�<i`�<L	�<٪�<'E�<���<�e�<M��<m�<��<�]�<N��<':�<G��<L�<Lc�<���<K�<�j�<L��<�<IW�<%��<��<�.�<s�<���<w��<8�<�w�<���<B��<3gz<��r<�`k<��c<e]\<��T<�_M<O�E<�k><��6</�/<R(<� <D<@�<�
<�2<.��;�6�;.��;C�;��;���;)T�;�*�;��;X-n;�\R;g�6;zL;k ;K�:P��:��>:JҪ9�l���~��	�`��ܢ���Ժ/2����K�3�ѣK�
.c��gz�I��������.��ݴ�J�����ɻPԻ{x޻Wx�[O�+�������r������f��v�����"��?&�b*�`t.��w2�Nl6��R:��+>���A�׶E��iI��M��P��?T���W��E[���^�&b�h�e���h��7l��o��r�Vv�n?y��q|�ǝ�b��o����������� ��I����+��Ǯ��0��﯐�c.������m'��U�����Ô��������������o���䠼�X���̣�h@������v&������r���}���ﭼ b��	԰�,F��U����*��#������݂��8����i�� ޽��  �  g�N=��M=�"M=�gL=��K=��J=�3J=�vI=O�H=q�G==G=~F=r�E=A�D=e=D=�{C=s�B=U�A=b2A=�m@=ͧ?=�>=N>=uP==r�<=K�;=��:=!:=�Q9=l�8=\�7=��6=u6=r/5=�V4=�{3=F�2=��1=��0=x�/=�/=�..=cD-=W,=g+=t*=�})=Ȅ(=C�'=Z�&=�%=�}$=�r#=d"=?Q!=M: ==h�=O�=��= �=�R=�=��=_�=	X=�=ڻ=�e=�
=>�=�D=��
=�i	=Y�=z=��=�v=��=�_ =���<�l�<E6�<'��<ȯ�<``�<c	�<Ъ�<3E�<���<�e�<M��<m�<
��<�]�<B��< :�<I��<;�<)c�<v��<4�<�j�<I��<�<CW�<-��<��<�.�<#s�<嵓<��<�7�<�w�<���<V��<jgz<�r<ak<��c<�]\<��T<`M<l�E<|k><��6<�/<_(<� <D<P�<��
<�2<��;�6�;ܴ�;�B�;�;Y��;/T�;Y*�;l�;�,n;�[R;9�6;LL;l ;��:���:��>:�ժ9�u��Ԃ��E�`��ݢ�Q�Ժ�1�����3���K��-c�gz�槈�I󓻍��7��ݴ�F����ɻ�OԻ�x޻Vx�DO�H�������r�����r�(w�	���"�6@&�!b*��t.��w2�Ql6��R:��+>��A�̶E�jI��M�?�P� @T���W��E[�K�^��%b�7�e�X�h��7l�փo���r�0v�R?y�dq|�֝�wb��z�$���k������� ��H����+��ɮ��0������{.�������'��T�����攙�������������o���䠼�X���̣�n@������k&�����j���}���ﭼ�a���Ӱ�F��C����*��������ǂ��%����i��޽��  �  n�N=��M=�"M=�gL=��K=��J=�3J=�vI=B�H=k�G=�<G=~F=s�E=8�D=\=D=�{C=v�B=Q�A=\2A=�m@=ç?=�>=A>=tP==o�<=L�;=��:=!:=R9=o�8=j�7=��6=w6=v/5=�V4=�{3=L�2=��1=��0=��/=�/=�..=kD-=W,=g+=t*=�})=��(=:�'=T�&=ۄ%=�}$=�r#=d"=<Q!=E: =	=d�=P�=��=�=�R=�=��=W�=X=�=�=�e=�
=D�=�D=��
=�i	=^�=z=��=�v=��=�_ =���<�l�<N6�<:��<ۯ�<q`�<j	�<̪�<7E�<���<�e�<<��<�l�<���<�]�<F��<�9�<7��<*�<(c�<p��<"�<�j�<0��<�<+W�<%��<��<�.�<2s�<ﵓ<���<8�<�w�<ƶ�<W��<wgz<-�r<3ak<��c<�]\<��T<)`M<��E<�k><��6<�/<~(<� <D<H�<Ǉ
<2<���;�6�;���;�B�;�;��;�S�;*�;u�;4,n;w[R;��6;�K; ;#�:e��:��>:'ժ9�l��������`��ݢ���Ժu1���Z�3��K��,c��fz�ۧ��Y�/�����ݴ������ɻ�OԻ�x޻Ox軉O�������s�����x�7w�+��"�J@&�#b*��t.��w2��l6��R:��+>���A�ȶE�jI�tM�'�P��?T���W��E[��^��%b�-�e�E�h��7l���o���r�*v�>?y�3q|�͝�hb��k����g����� ��_����+��ܮ��30��
����.�������'��e���)��甙����σ������o���䠼Y���̣�l@������\&�����Z���}���ﭼ�a���Ӱ�F��7����*��������Ƃ������i��޽��  �  m�N=��M=�"M=�gL=��K=��J=�3J=�vI=?�H=a�G=�<G=�}F=g�E=1�D=J=D=�{C=b�B=C�A=Q2A=�m@=��?=
�>=D>=mP==t�<=H�;=��:=!!:=R9=�8=d�7=��6=�6=�/5=�V4=�{3=W�2=��1=��0=��/=/=/.=kD-=$W,=g+=t*=�})=��(==�'=O�&=ք%=�}$=�r#=d"=9Q!=:: =�=b�=:�=��=�=�R=�=��=W�=X=�=ٻ=�e=�
=N�=�D=��
=�i	=p�="z=��=�v=��=�_ =Ԛ�<�l�<s6�<E��<��<�`�<c	�<ܪ�<+E�<���<�e�<9��<�l�<���<�]�<��<�9�<��<�<c�<M��<�<�j�<(��<�
�<2W�<��<��<�.�<&s�<���<���<8�<�w�<ʶ�<}��<�gz<`�r<@ak<�c<�]\<=�T<:`M<��E<�k><��6<5�/<v(<� <D</�<ׇ
<m2<���;:6�;]��;+B�;��;�;ES�;�)�;��;<+n;�ZR;�6;4K;� ;1�::��:��>:uҪ9i�������`��ۢ���Ժ�0�����3�q�K��,c�*fz�e�����R������ܴ������ɻ�OԻ�x޻sx軡O�������s��$����Ew�]��<"�T@&�~b*��t.�x2��l6�S:��+>���A�߶E�jI��M��P��?T���W�ZE[�/�^��%b��e��h��7l���o���r��v�
?y�Nq|����bb��g�
���s������� ��]����+��⮍�=0�� ����.��ǫ���'������=���������ك������o���䠼 Y���̣�l@������h&������_���}���ﭼ�a���Ӱ��E������*��������������i���ݽ��  �  o�N=��M=�"M=�gL=��K=��J=�3J=�vI=>�H=T�G=�<G=�}F=U�E=*�D=@=D=�{C=Q�B=A�A=H2A=zm@=��?=��>=G>=gP==w�<=H�;=��:=)!:=R9=��8=n�7=��6=�6=�/5=�V4=
|3=e�2=��1=��0=��/=/=/.=mD-=-W,=
g+=t*=�})=��(=7�'=C�&=ل%=�}$=�r#=�c"=+Q!=2: =�=U�=-�=��=�=�R=�=��=[�=X=�=ڻ=�e=�
=S�=�D=��
=�i	=q�=2z=��=�v=��=�_ =���<	m�<�6�<L��<��<�`�<e	�<��<#E�<���<�e�<)��<�l�<���<�]�<���<�9�<��<
�<�b�<9��<�<�j�<'��<�
�<,W�<��<��<�.�<'s�<��<���<'8�<�w�<㶄<���<�gz<��r<zak<U�c<�]\<^�T<x`M<��E<�k><��6<^�/<�(<�� <D<%�<ԇ
</2<���;�5�;#��;�A�;�;���;�R�;�)�;3�;�*n;�YR;�6;�J;� ;@�:S�:��>:KѪ9#f��7}��-�`�ۢ���Ժ!0���L�3���K��+c�bez���������d���ܴ�
���q�ɻ�OԻ�x޻�x軖O����"��s�A�+����w����e"��@&��b*��t.�?x2��l6�.S:��+>���A���E��iI��M��P��?T�~�W�;E[�
�^��%b���e���h�W7l�S�o�g�r��v��>y�%q|�i��`b��]����u������!��V���,������E0��7����.��竓��'������I��������ボ�4����o���䠼Y���̣�q@������f&��嘩�[���}���ﭼ�a���Ӱ��E�����e*��ќ��������������i���ݽ��  �  ~�N=��M=�"M=�gL=��K=��J=|3J=�vI=8�H=L�G=�<G=�}F=Q�E=�D=2=D=�{C=Q�B=8�A=<2A=rm@=��?=��>==>=gP==r�<=K�;=��:=,!:=R9=��8=~�7=��6=�6=�/5=�V4=|3=q�2=��1=��0=��/=/=/.=yD-=*W,=g+=
t*=�})=��(=3�'=B�&=Є%=�}$=�r#=�c"=!Q!=%: =�=I�=/�=u�=��=�R=�=��=U�=X=�=�=�e=�
=`�=�D=��
=�i	=��=Bz=��=�v=��=�_ =���<-m�<�6�<j��<��<�`�<q	�<ߪ�<(E�<���<~e�<"��<�l�<���<y]�<��<�9�<��<��<�b�<3��<��<rj�<��<�
�<W�<��<��<�.�<0s�<��<���<18�<�w�<���<���<�gz<��r<�ak<t�c<9^\<u�T<�`M<��E<�k><�6<`�/<�(<�� <D<�<��
<(2<N��;�5�;���;�A�;�߽;���;oR�;)�;$�;K*n;YR;�6;/J;n ;��:�:�>:�Ѫ9�i���|���`�Zۢ��Ժ�/�u��V�3�[�K�m+c��dz�����򓻲��W��cܴ�������ɻ�OԻ�x޻�x��O�����)��:s�l�a����w�����"��@&��b*�u.�ex2��l6�6S:�,>���A���E�jI��M���P��?T�R�W�9E[�Ϲ^��%b���e���h�.7l�2�o�)�r��v��>y��p|�o��Fb��Q����l������!��i���,������T0��M����.��㫓��'������e��%���������F����o���䠼Y���̣�r@������\&��阩�=��{}���ﭼ�a���Ӱ��E��񷳼Q*��Ü��������������i���ݽ��  �  ��N=��M=�"M=�gL=��K=��J=w3J=�vI=(�H=N�G=�<G=�}F=E�E=�D=0=D=�{C=D�B=%�A=<2A=mm@=��?=��>=6>=nP==o�<=L�;=��:=(!:=R9=��8=��7=��6=�6=�/5=�V4=$|3=r�2=��1=��0=��/=/=/.=zD-=*W,=g+=t*=�})=��(=1�'=>�&=��%=�}$=�r#=�c"=Q!=: =�=?�= �=f�=�=�R=�=��=N�=X=�=�=�e=�
=f�=�D=��
=�i	=��=Fz=�=�v=��=�_ =��<Hm�<�6�<y��<���<�`�<{	�<۪�<<E�<���<�e�<��<�l�<���<U]�<���<�9�<��<��<�b�<��<��<|j�<���<�
�<W�<	��<��<�.�<>s�<��<���<58�<�w�<	��<���<Chz<��r<�ak<��c<t^\<��T<�`M<&�E<�k><�6<R�/<�(<�� <D< �<��
<,2<���;�5�;x��;A�;�߽;���;NR�;�(�;��;)n;�XR;k�6;ZI;q ;��:��:��>:?Ѫ9�c��s��(�`�ۢ���Ժ�/�p��	�3�ŠK�*c��dz�f���8�Y��8��Pܴ�������ɻ�OԻ�x޻fx�P�����=��}s�Q����F��w�����"��@&��b*�Lu.�Lx2��l6�RS:�,>���A�ͶE�jI�oM��P��?T�D�W�'E[���^�e%b�a�e���h��6l��o��r�dv��>y��p|�]��<b��X�����f������� ��x���
,�����g0��G����.������'������}��?��������<����o���䠼Y���̣�n@������O&��𘩼7��v}���ﭼ�a���Ӱ��E��鷳�-*������e��l��������i���ݽ��  �  ��N=��M=�"M=�gL=��K=��J=s3J=�vI=%�H=@�G=�<G=�}F=B�E=�D=$=D=�{C=A�B=&�A=12A=`m@=��?=��>=0>=gP==s�<=K�;=��:=3!:=R9=��8=��7=��6=�6=�/5=�V4=-|3=z�2=��1=��0=��/= /=/.=D-=5W,=g+=t*=�})=��(=*�'=7�&=��%=�}$=�r#=�c"=Q!=: =�=;�=�=d�=��=�R=�=|�=J�=X=�=�=f=�
=p�=�D=��
=�i	=��=Nz=�=�v=��=�_ =$��<Tm�<�6�<���<��<�`�<|	�<��<0E�<���<ue�<��<�l�<���<W]�<���<�9�<ʠ�<��<�b�<��<��<_j�<�<�
�<W�<���<��<�.�<@s�<��<���<M8�<x�<��<���<<hz<��r<bk<��c<r^\<��T<�`M<D�E<7l><(�6<��/<�(<�� <D<�<��
<2<���;5�;5��;A�;c߽;P��;�Q�;i(�;��;�(n;0XR;��6;I;� ;��:~�:'�>:�Ϫ9]��yz��'�`��٢���ԺK/�U���3�L�K�*c�Pdz�w����.�����ܴ�����E�ɻ�OԻ�x޻�x�=P�6���Y���s������N��w����"��@&��b*�Uu.�x2�	m6�gS:�(,>���A��E�jI�rM�ɭP��?T�#�W��D[���^�G%b�`�e���h��6l��o��r�]v��>y��p|�1��/b��D��i������!������,�����~0��`����.������'��Ԣ�����H����� ���Y����o���䠼'Y��
ͣ�n@������L&��ט��/��_}��wﭼ�a���Ӱ��E��ط��*������g��e�������}i���ݽ��  �  ��N=��M=�"M=�gL=��K=��J=|3J=�vI=)�H=7�G=�<G=�}F=4�E=�D==D=�{C=4�B=�A=&2A=]m@=��?=��>=;>=`P==t�<=M�;=��:=6!:=R9=��8=��7=��6=�6=�/5=�V4=-|3=��2=��1=��0=��/=!/=/.=�D-=4W,=g+=t*=�})=��(=.�'=4�&=��%=�}$=�r#=�c"=Q!=: =�=0�=�=^�=�=�R=�=~�=T�=X=�=�=f=�
=q�=�D=��
=�i	=��=cz=�=�v=��=` =C��<_m�<�6�<���<��<�`�<	�<��< E�<���<re�<��<�l�<���<I]�<���<�9�<���<��<�b�<���<��<Ij�<���<�
�<W�<���<��<�.�<6s�<"��<���<R8�<x�<&��<���<ehz<7�r<bk<��c<�^\<��T< aM<L�E<Al><�6<��/<�(<� <�C<��<��
<�1<���;�4�;��;�@�;�޽;��;�Q�;(�;�;B(n;iWR;D�6;I;� ;��:y}�:.�>:RЪ9�h���y��8�`��٢�:�Ժ�.�����3��K�	*c�cz�S����������ܴ�����U�ɻ�OԻ�x޻�x�P����h��s���Ț�w�"x����"�.A&�,c*�qu.��x2� m6�uS:�#,>���A��E��iI��M�ѭP��?T�$�W��D[�u�^�%b�T�e�?�h��6l�˂o���r�Nv�X>y��p|�-��1b��>�����h������!��m���,�����0��y����.��"���(��碖����b���.��0���n����o���䠼Y��ͣ�{@������U&��Ҙ��3��Z}��tﭼza���Ӱ��E������*������M��T�������yi���ݽ��  �  ��N=��M=�"M=�gL=��K=��J=q3J=vI=�H=;�G=�<G=�}F=4�E=��D==D=�{C=2�B=�A=/2A=[m@=��?=��>=3>=bP==r�<=O�;=��:=9!:="R9=��8=��7=��6=�6=�/5=�V4=4|3=��2=��1=��0=��/='/=/.=�D-=7W,=g+=t*=�})=��(=$�'=,�&=��%=�}$=�r#=�c"=Q!=: =�=/�=�=`�=�=�R=�=u�=Q�=X=�=�=f=�
=u�=�D=��
=�i	=��=`z=�=�v=��=` =@��<im�<�6�<���<'��<�`�<�	�<��<&E�<���<be�<���<�l�<���<F]�<���<�9�<���<��<�b�<�<��<Uj�<߻�<�
�<W�<���<��<�.�<Bs�<%��<���<V8�<x�<)��<���<ihz<0�r<7bk<��c<�^\<��T<aM<`�E<Kl><;�6<��/<�(<� <�C<��<��
<�1<o��;�4�;��;�@�;�޽;���;�Q�;�'�;�;.(n;�WR;�6;eH;� ;��:�}�:r�>:�Ъ9-a���x����`�;٢���Ժ�.�7��!�3���K��)c�|cz�P������������۴�]���?�ɻ�OԻ�x޻�x�!P�e�������s��������)x����"�2A&�9c*�iu.��x2�$m6��S:�H,>���A��E��iI�qM�ĭP�z?T��W��D[�n�^�%b�R�e�R�h��6l���o���r�Pv�b>y��p|���%b��8�����d������!��|���0,��)����0��i����.��&���(��⢖����c���3��%���b����o���䠼.Y��	ͣ�z@������J&��Ϙ��%��V}��hﭼwa���Ӱ��E������*������L��U�������pi���ݽ��  �  '�N=��M=M=�`L=��K=��J=z*J=�lI=��H=��G=�0G=�pF=+�E=�D=6-D=�jC=T�B=(�A=2A=NX@=w�?=��>=� >=�6==�k<= �;=r�:=j:=�19=`8=��7=��6=��5=Q5=�-4=�Q3=ms2=�1=��0=��/=c�.=��-=N-==,=h-+=�8*=�@)=�E(=�G'=�E&=�@%=�7$=c+#="=�!=;�=��=��=J�=da=�2=��=��=�=&I=f=��=�e=�=��=�T=6�=Ԅ
=r	=�=�'=v�=k&=��=P =��<0��<���<di�<�%�<%��<��<�,�<��<�b�<2��<3�<Z�<��<��<Hs�<���<zO�<��<��<sz�<�ִ< 0�<��<�٩<0*�<�x�<�Ğ<P�<X�<O��<Z�<C*�<Vn�<���<��<�nz<�r<�yk<��c<5�\<U<��M<�'F<�><�I7<r�/<Jy(<B!<��<�a<<x�<���;y�;��;��;gX�;��;��;<֔;ӆ;�q;mV;�:;�P;[8;��:Q�:�P:�9��44�͹�L����ٍʺ����7J��].�<%F�Y�]���t�Յ�����:��&1������F���!ǻuѻR�ۻ���a��\6��@b�����
��F�@��>.����� �-	%��1)��J-��T1�
P5�S=9�F=�9�@���D��pH��L�?�O�\S���V��oZ�C�]��]a���d��)h�g�k���n��!r�
fu�n�x���{������ձ��?C��R҅�C_��ꈼ�r������8������������؄��������V����u���xh��i����W��7Π�QD��ι���.���������틩�����^s���歼rZ���Ͱ�cA�������(���������;������Ko���佼�  �  '�N=��M=M= aL=��K=��J=w*J=�lI=��H=��G=�0G=�pF=,�E=�D=3-D=�jC=T�B=0�A=3A=OX@=s�?=��>=� >=�6==�k<=$�;=u�:=o:=�19=`8=��7=��6=��5=S5=�-4=�Q3=rs2=�1=��0=��/=c�.=��-=P-=D,=g-+=�8*=�@)=�E(=�G'=�E&=�@%=�7$=h+#=	"=�!=;�=��=��=L�=ja=�2=��=��=�="I=_=��=�e=�=��=T=6�=ׄ
=p	=�=�'=m�=g&=��=H =��<*��<���<di�<�%�</��<��<�,�<��<�b�<��<'�<]�<��<��<Es�<���<vO�<��<��<�z�<�ִ<�/�<��<_٩<%*�<�x�<�Ğ<Z�<X�<\��<Z�<>*�<Sn�<���<��<�nz<�r<�yk<��c<<�\<U<��M<�'F<��><�I7<��/<Ly(<S!<��<�a<<9�<���;y�;��;G��;lX�;�;l�;Q֔;ӆ;{�q;�V;��:;�P;]7;ϧ�:�P�:��P:��9@5t�͹��L�Q���6�ʺ�����J��].�B%F��]�N�t�%Յ�����:��$1��
���0���� ǻ uѻ.�ۻ*��w�ﻤ6��xb�|���
��F�3��0.����� �	%��1)��J-��T1��O5�~=9�p=�E�@���D��pH��L�&�O�\S���V��oZ�7�]��]a���d�)h���k�	�n�u!r�-fu�n�x���{������˱��5C��L҅�>_��ꈼ�r������D������������ۄ��������S����u���lh��n����W��XΠ�\D��Թ���.���������ߋ������cs���歼hZ���Ͱ�bA�������(���������C������No���佼�  �   �N=��M=M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=,�E=�D=4-D=�jC=S�B=4�A=2A=SX@=|�?=��>=� >=�6==�k<= �;=l�:=g:=�19=`8=��7=��6=��5=T5=�-4=�Q3=ts2=�1=z�0=��/=`�.=��-=I-==,=_-+=�8*=�@)=�E(=�G'=�E&=�@%=�7$=l+#="=�!=>�=��=��=J�=oa=�2=��=��=�=+I=a=��=�e=�=��={T=2�=҄
=k	=��=�'=g�=e&=��=C =��<!��<��<Yi�<�%�<��<���<�,�<��<�b�<��<:�<i�<��<(��<Ds�<���<yO�<��<��<�z�<�ִ<�/�<&��<e٩<8*�<�x�<�Ğ<[�<X�<O��<L�<>*�<Ln�<���<��<�nz<&�r<ryk<��c<2�\<�U<��M<s'F<��><yI7<n�/<'y(<P!<��<�a<%<B�<0��;y�;��;_��;nX�;:�;w�;|֔;ӆ;��q;{V;A�:;eQ;�7;��:�P�:A�P:]�9j��4K�͹͛L�)���|�ʺm����J��].�@%F���]�$�t�/Յ����:��<1�����f���!ǻauѻ�ۻ��:��Q6��ab�T���
�xF�9��-.����� �	%��1)�J-��T1��O5�`=9�J=�#�@���D��pH��L�F�O�/\S���V��oZ�I�]��]a���d�v)h���k��n�k!r�;fu�m�x���{������ޱ��IC��[҅�:_��ꈼ�r������0������������܄��������H����u���jh��p����W��RΠ�ID��ι���.���������싩�����cs���歼kZ���Ͱ�hA��𴳼�(���������M������Uo���佼�  �  "�N=��M=M=�`L=��K=��J=z*J=�lI=��H=��G=�0G=�pF=0�E=�D==-D=�jC=Y�B=7�A=<A=VX@=y�?=��>=� >=�6==�k<="�;=v�:=j:=�19=`8=��7=��6=��5=H5=�-4=�Q3=bs2=	�1=v�0=��/=[�.=��-=I-=A,=h-+=�8*=�@)=�E(=�G'=�E&=�@%=�7$=q+#="=�!=G�=��=��=P�=qa=�2=��=��=�= I=d=��=�e=�=��={T=,�=΄
=e	=��=�'=g�=^&=��=D =��<��<��<Zi�<�%�<)��<��<�,�<��<�b�<#��<4�<h�<���<,��<Qs�<���<�O�<��<��<�z�<�ִ<0�<��<o٩<0*�<�x�<�Ğ<X�<X�<T��<M�<:*�<En�<���<��<�nz<��r<�yk<��c<�\<�U<}�M<f'F<�><}I7<v�/<Ty(<I!<�<�a<<W�<��;Ty�;	�;���;�X�;X�;��;�֔;7ӆ;�q;,V;��:;7Q;8;3��:�P�:��P:��915b�͹�L�������ʺo����J�e^.��%F�.�]�5�t�7Յ�4��;��]1�����d���� ǻuѻ2�ۻ���{��Z6��Ub�i���
�bF�$��.������ �		%��1)�rJ-�dT1��O5�`=9�G=�J�@���D��pH��L�-�O�*\S���V��oZ�U�]��]a���d��)h���k�%�n��!r�5fu���x���{�����ױ��6C��S҅�=_��ꈼ�r������5�����䄐����΄��������=����u���\h��Z����W��HΠ�QD��׹���.���������狩�����hs���歼xZ���Ͱ�sA������(���������M���'���[o��彼�  �  �N=��M=
M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=9�E=�D=D-D=�jC=a�B=:�A=?A=[X@=z�?=��>=� >=�6==�k<=�;=o�:=b:=�19=`8=��7=��6=��5=D5=�-4=�Q3=\s2=�1=n�0=��/=U�.=��-=E-=:,=d-+=�8*=�@)=�E(=�G'=�E&=�@%=�7$=q+#="=�!=H�=��=��=Z�=qa=�2=��=��=�=#I=h=��=�e=�=��=sT=#�=̈́
=Y	=��=�'=`�=U&=��=< =��<��<Ѥ�<Mi�<�%�<��<���<�,�<"��<�b�<1��<6�<o�<��<-��<cs�<���<�O�<!��<��<�z�<�ִ<0�<��<٩<<*�<�x�<�Ğ<O�<X�<F��<H�<&*�<An�<���<��<�nz<��r<uyk<��c<�\<�U<g�M<d'F<ɶ><qI7<V�/<<y(<7!<�<�a<#<{�<��;�y�;+	�;���;�X�;x�;�;�֔;�ӆ;E�q;oV;�:;dQ;�8;Ȩ�:�Q�:\�P:��9�g�4˅͹"�L�Ǵ��_�ʺ(���K��^.�&F�\�]���t�JՅ�p���:���1��P������'!ǻ*uѻM�ۻϤ�N��'6��Ab�^�{�
�aF����.������ ��%�W1)�oJ-�KT1��O5�Q=9�-=�9�@�u�D��pH��L�K�O�<\S���V��oZ�R�]�^a���d��)h���k�A�n��!r�Kfu���x���{�7���求�FC��W҅�<_���鈼�r������2�����ڄ���������������:����u���\h��P����W��9Π�ED��ʹ���.�����������������zs���歼Z���Ͱ�tA�� ����(��ǜ�����[���1���[o��彼�  �  �N=��M=M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=?�E=�D=I-D=�jC=g�B=G�A=?A=_X@=��?=��>=� >=�6==�k<= �;=n�:=e:=�19=`8=��7=��6=��5=?5=�-4=�Q3=^s2=��1=i�0=��/=R�.=��-=E-=<,=_-+=�8*=�@)=�E(=�G'=�E&=�@%=�7$={+#="=�!=S�=��=��=]�=}a=�2=��=��=��=&I=^=��=�e=�=��=pT=�=Ä
=V	=�=�'=O�=J&=��=+ =��< ��<ˤ�<Gi�<�%�<��<���<�,�<��<�b�<+��<I�<z�<���<H��<ls�<���<�O�<:��<��<�z�< ״<0�<=��<~٩<A*�<�x�<�Ğ<]�<X�<K��<B�<&*�<5n�<���<~�<hnz<��r<?yk<��c<چ\<�U<X�M<C'F<Ƕ><aI7<^�/<-y(<J!<��<�a<0<y�<���;�y�;S	�;��;Y�;��;6�;)ה;�ӆ;8�q;�V;<�:;NR;�8;���:�P�:��P:N�9 5u�͹��L�������ʺ����K��^.�n&F�G�]�\�t��Յ����-;���1��R���x���!ǻMuѻ��ۻ��I��,6��;b�#���
�2F�����-����]� ��%�G1)�<J-�VT1��O5�@=9�5=�)�@���D��pH��L�F�O�8\S���V��oZ�q�]�^a��d��)h��k�g�n��!r��fu���x���{�=���᱂�HC��Z҅�7_��ꈼ�r�����������݄��k���������u��!����u��tNh��Q����W��;Π�BD��չ���.���������񋩼����{s��筼�Z��ΰ��A������(��ʜ�����u���8���jo��彼�  �  �N=��M=M= aL=��K=��J=�*J=�lI=��H=��G=�0G=�pF=A�E=)�D=N-D=�jC=h�B=S�A=MA=bX@=��?=��>=� >=�6==�k<=�;=k�:=c:=�19=`8=��7=��6=��5=25=�-4=�Q3=Ts2=�1=m�0=��/=L�.=��-=:-=<,=Z-+=�8*=�@)=�E(=�G'=�E&=�@%=�7$=�+#="=�!=Z�=��=ð=^�=�a=�2=��=��=�=-I=]=��=�e=�=��=dT=�=��
=X	=ڠ=�'=H�=D&=��=! =��<���<Ĥ�<*i�<�%�<��<��<�,�<��<�b�<&��<L�<�<��<c��<ls�<���<�O�<P��<��<�z�<$״<0�<G��<~٩<N*�<�x�<�Ğ<c�<X�<O��<+�<*�< n�<���<��<4nz<��r<yk<z�c<��\<�U<J�M<'F<��><.I7<`�/<y(<M!<�<�a<L<s�<���;�y�;�	�;N��;4Y�;F�;d�;�ה;�ӆ;�q;xV;��:;�R;�8;���:�Q�:��P:��9���4��͹�L�{����ʺ����*L��_.��&F���]���t�օ�k���;���1������Ǥ��!ǻsuѻʠۻ����6��/b��m�
��E�����-�j��E� ��%�@1)��I-�8T1��O5�3=9�,=�
�@���D��pH��L�C�O�]\S��V�pZ���]��]a�J�d��)h���k�x�n��!r��fu���x��{�D���豂�JC��a҅�'_��ꈼ�r�����������Ƅ��O���������l������u��k*h��L����W��;Π�6D��ȹ���.��������������s��筼�Z��ΰ��A��-����(��֜����s���=����o��彼�  �  �N=��M=�M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=N�E=/�D=V-D=�jC=t�B=O�A=TA=lX@=��?=��>=� >=�6==�k<=�;=d�:=]:=�19=`8=��7=q�6=��5=-5=�-4=�Q3=Js2=�1=^�0=|�/=H�.=��-=;-=5,=Z-+=�8*=�@)=�E(=�G'=�E&=�@%=8$=�+#=%"=�!=^�=��=ΰ=h�=�a=
3=��=��=��=*I=`=��=�e=�=��=_T=�=��
=E	=נ={'=A�=9&=x�= =u�<���<���<!i�<�%�<���<��<�,�<��<�b�<9��<V�<��<&��<Z��<�s�<���<�O�<Z��<��<�z�<"״<70�<I��<�٩<P*�<�x�<�Ğ<W�<�W�<?��<0�<*�<n�<n��<o�<.nz<t�r<yk<H�c<��\<zU<�M<'F<��><5I7<C�/<	y(<:!<�<�a<J<��<���;z�;�	�;V��;�Y�;|�;��;�ה;?Ԇ;��q;V;E�:;�R;j9;���:OR�:K�P:B�9���4��͹��L�Ĵ���ʺ����LL��_.�;'F�ء]���t�
օ�����;���1����������@!ǻnuѻ�ۻ�����5���a��6�
��E�����-�X��2� �%�1)�J-�T1��O5�=9�=��@���D��pH��L�a�O�a\S�(�V�pZ���]�B^a�O�d� *h��k���n�"r��fu��x��{�M�$��󱂼YC��e҅�1_��ꈼ�r���������������W���������\������u��c,h��5����W�� Π�3D�������.������������������s��$筼�Z��ΰ��A��E���)��휶�������^����o��$彼�  �  �N=��M=M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=X�E=1�D=d-D=�jC=��B=Y�A=YA=qX@=��?=��>=� >=�6==�k<=#�;=h�:=\:=�19=�_8=��7=i�6=��5=(5=�-4=�Q3=?s2=�1=P�0=�/=A�.=��-==-=/,=c-+=�8*=�@)=�E(=�G'=�E&=�@%=8$=�+#=4"=�!=i�=��=Ͱ=v�=�a=3=��=��=��=)I=c=��=�e=�=��=XT=	�=��
=6	=Ѡ=p'=5�=+&=p�= =\�<���<���<i�<~%�<���<���<y,�<��<�b�<7��<V�<��<3��<g��<�s�<���<�O�<d��<��<�z�<%״<M0�<G��<�٩<J*�<�x�<�Ğ<[�<X�<4��<2�<�)�<n�<l��<T�<nz<C�r<�xk<�c<��\<JU<��M<'F<i�><6I7<1�/<)y(<H!<��<�a<?<��<���;Oz�;
�;̩�;�Y�;��;)�;�ה;�Ԇ;��q;vV;��:;S;�9;Ϊ�:S�:��P:Y�9�;�4~�͹>�L�����ϐʺ�����L�`.��'F�L�]��t�'օ�F���;��2����������m!ǻ#uѻ'�ۻ̤�����5���a���
��E�y���-�*���� ��%��0)�J-��S1��O5�=9�=��@�v�D��pH��L�u�O�W\S�=�V�7pZ���]�x^a�^�d�C*h�;�k���n�)"r��fu��x��{���$��򱂼WC��S҅�C_���鈼�r������
���������I��}������=�������u��F*h������W��Π�:D�������.�����������������s��(筼�Z��8ΰ��A��\���)�����#������d����o��C彼�  �  
�N=��M=�M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=Z�E=:�D=i-D=�jC=��B=`�A=\A=sX@=��?=��>=� >=�6==�k<=�;=b�:=V:=�19=�_8=~�7=i�6=��5= 5=�-4=�Q3=;s2=ܒ1=O�0=y�/==�.=��-=6-=+,=]-+=�8*=�@)=�E(=�G'=�E&=�@%=8$=�+#=9"=�!=o�=��=Ѱ=z�=�a=3=��=��=��=0I=e=��=�e=�=��=TT=�=��
=4	=Ơ=i'=1�=(&=g�=	 =Z�<���<���<i�<p%�<���<��<�,�<!��<�b�<>��<h�<��<3��<w��<�s�<���<�O�<t��<�<�z�<1״<L0�<]��<�٩<Z*�<�x�<�Ğ<V�<�W�<,��<#�<�)�<n�<h��<N�<�mz<2�r<�xk<�c<^�\<6U<�M<�&F<f�><I7<�/<y(<8!<	�<b<^<��<��;Kz�;9
�;
��;Z�;��;W�;'ؔ;�Ԇ;�q;�V;�:;�S;�9;��:�S�:1�P:O�9���4��͹��L�����G�ʺ����9M�v`.��'F���]�V�t�qօ�G���;��-2������ؤ���!ǻQuѻ�ۻ��廵�ﻯ5���a����
��E�c��z-����� �l%��0)��I-��S1�mO5��<9��=���@�h�D��pH��L���O�r\S�I�V�GpZ���]�z^a���d�W*h�H�k���n�D"r��fu��x�,�{���/������bC��]҅�:_���鈼�r�������~���������9��x���z��6�������u��9h��!���oW��Π�*D�������.�����������������s��3筼�Z��>ΰ��A��e���)�����4������g����o��C彼�  �  �N=��M= M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=b�E=E�D=b-D=�jC=��B=b�A=bA=xX@=��?=��>=� >=�6==�k<=�;=g�:=Y:=�19=�_8=s�7=b�6=��5=5=�-4=|Q3=8s2=֒1=M�0=p�/=>�.=��-=2-=5,=[-+=�8*=�@)=�E(=�G'=�E&=�@%=8$=�+#=7"=�!=s�=��=�=y�=�a=3=��=��=��=(I=\=��=�e=�=��=ST=�=��
=0	=��=d'=%�=&=b�= =L�<���<���<i�<r%�<���<���<�,�<��<�b�<<��<i�<��<;��<|��<�s�<��<�O�<���<�<�z�<D״<P0�<f��<�٩<V*�<�x�<�Ğ<U�< X�<<��<�<*�<�m�<T��<F�<�mz<&�r<�xk<��c<H�\<$U<ΙM<�&F<|�><�H7<5�/<y(<4!<�<�a<U<��<*��;fz�;�
�;��;UZ�;B�;)�;�ؔ;�Ԇ;I�q; V;?�:;�S;�9;���:�R�:�P:R�9� 5��͹��L�ǵ����ʺ@���eM��`.�R(F��]�x�t��օ�R��(<��2����������5!ǻYuѻ�ۻ������5���a����
��E�i��8-������ �#%��0)��I-��S1�[O5��<9�=��@���D��pH��L�\�O�z\S�F�V�6pZ���]��^a���d�g*h�p�k���n�U"r�gu�-�x�X�{�}�6������SC��d҅�4_��ꈼ�r�������~���������3��s���X��A������~u��<h�����fW��Π�/D��Ĺ���.�����������������s��=筼�Z��Eΰ��A��j���,)�����?������w����o��8彼�  �  �N=��M=�M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=d�E=D�D=k-D=�jC=��B=h�A=cA={X@=��?=��>=� >=�6==�k<=�;=c�:=P:=�19=�_8=t�7=a�6=��5=5=�-4=yQ3=4s2=֒1=G�0=q�/=6�.={�-=,-=+,=Y-+=�8*=�@)=�E(=�G'=�E&=�@%=8$=�+#=;"=�!=t�=��=�={�=�a=3=��=��= �=0I=d=��=�e=�=��=KT=��=��
=*	=��=b'=#�=&=`�= =E�<���<���<�h�<\%�<���<݆�<,�<��<�b�<J��<i�<��<@��<���<�s�<��<�O�<���<�<�z�<D״<V0�<e��<�٩<g*�<�x�< Ş<R�< X�<*��<�<�)�<�m�<V��<>�<�mz<�r<�xk<��c<I�\<U<ЙM<�&F<S�><�H7<�/<	y(</!<�<�a<u<��<&��;�z�;�
�;.��;gZ�;>�;r�;�ؔ;Ն;��q;> V;z�:;�S;y:;���:�S�:��P:Q�9�6�4I�͹M�L����n�ʺ_���dM��`.��(F�6�]���t��օ���<��Y2�� ��%����!ǻkuѻ�ۻ��廪��u5���a�����
��E�Z��B-������ �.%��0)��I-��S1�PO5��<9��=���@�g�D��pH��L���O��\S�f�V�ZpZ���]��^a���d�n*h�y�k� �n�Y"r��fu�8�x�U�{���?�����`C��f҅�9_���鈼�r�������~���������'��n���]��1������~u��4h�����gW��Π�D�������.�����������������s��B筼�Z��Lΰ��A��u���-)�����>������v����o��L彼�  �  �N=��M=M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=b�E=B�D=y-D=�jC=��B=j�A=_A=|X@=��?=��>=� >=�6==�k<=�;=f�:=V:=�19=�_8=w�7=[�6=��5=5=�-4=zQ3=1s2=ג1=A�0=q�/=4�.=��-=;-=-,=_-+=�8*=�@)=�E(=�G'=�E&=�@%=8$=�+#=B"=�!=y�=��=۰=��=�a=3=��=��=��=*I=d=��=�e=�=��=TT=��=��
=%	=��=^'=#�=&=]�=� =:�<���<���<i�<m%�<���<��<v,�<��<�b�<H��<n�<��<7��<���<�s�<��< P�<���<�<�z�<?״<Z0�<j��<�٩<Z*�<�x�<�Ğ<O�<X�<+��<0�<�)�<�m�<Q��<0�<�mz<�r<�xk<��c<H�\<�U<��M<�&F<X�></I7<�/<y(<.!< �<�a<\<��<:��;�z�;o
�;^��;XZ�;,�;��;uؔ;Ն;��q;�V;��:;!T;s:;���:�S�:��P:��9���4�͹D�L�����ʺ%����M��`.��(F��]���t��օ����<��k2����������m!ǻ:uѻ6�ۻ���؀ﻜ5���a����
��E�:��U-����� �B%��0)��I-��S1�QO5��<9��=��@�g�D��pH��L�t�O�l\S�@�V�fpZ���]��^a���d�{*h�v�k� �n�f"r�gu�N�x�I�{���������[C��\҅�B_���鈼�r�������~���������#��j���g���������u��%h�����bW��Π�*D�������.�����������������s��D筼�Z��[ΰ��A��{���')��%���>����������o��J彼�  �  �N=��M=�M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=d�E=D�D=k-D=�jC=��B=h�A=cA={X@=��?=��>=� >=�6==�k<=�;=c�:=P:=�19=�_8=t�7=a�6=��5=5=�-4=yQ3=4s2=֒1=G�0=q�/=6�.={�-=,-=+,=Y-+=�8*=�@)=�E(=�G'=�E&=�@%=8$=�+#=;"=�!=t�=��=�={�=�a=3=��=��= �=0I=d=��=�e=�=��=KT=��=��
=*	=��=b'=#�=&=a�= =E�<���<���<�h�<]%�<���<݆�<,�<��<�b�<K��<j�<��<A��<���<�s�<��<�O�<���<�<�z�<D״<V0�<e��<�٩<f*�<�x�< Ş<Q�< X�<*��<�<�)�<�m�<V��<>�<�mz<�r<�xk<��c<I�\<U<љM<�&F<S�><�H7<�/<	y(</!<�<�a<v<��<'��;�z�;�
�;/��;hZ�;>�;r�;�ؔ;Ն;��q;; V;w�:;�S;v:;���:�S�:��P:1�9?��4j�͹^�L����v�ʺg���hM��`.��(F�:�]���t��օ���� <��Z2�� ��&����!ǻkuѻ�ۻ��廫��u5���a�����
��E�Z��B-������ �.%��0)��I-��S1�PO5��<9��=���@�g�D��pH��L���O��\S�f�V�ZpZ���]��^a���d�n*h�y�k� �n�Y"r��fu�8�x�U�{���?�����`C��f҅�9_���鈼�r�������~���������'��n���]��1������~u��4h�����gW��Π�D�������.�����������������s��B筼�Z��Lΰ��A��u���-)�����>������v����o��L彼�  �  �N=��M= M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=b�E=E�D=b-D=�jC=��B=b�A=bA=xX@=��?=��>=� >=�6==�k<=�;=g�:=Y:=�19=�_8=s�7=b�6=��5=5=�-4=|Q3=8s2=֒1=M�0=p�/=>�.=��-=2-=5,=[-+=�8*=�@)=�E(=�G'=�E&=�@%=8$=�+#=7"=�!=s�=��=�=y�=�a=3=��=��=��=(I=\=��=�e=�=��=TT=�=��
=0	=��=e'=&�=&=b�= =M�<���<���<i�<s%�<���<��<�,�<��<�b�<=��<j�<��<;��<|��<�s�<��<�O�<���<�<�z�<D״<O0�<f��<�٩<V*�<�x�<�Ğ<U�<�W�<;��<�<*�<�m�<T��<F�<�mz<%�r<�xk<��c<H�\<$U<ϙM<�&F<}�><�H7<6�/<y(<6!<�<�a<V<��<+��;gz�;�
�;��;VZ�;B�;(�;�ؔ;�Ԇ;F�q; V;;�:;�S;�9;���:�R�:��P:�9T 5�͹��L�׵����ʺO���lM��`.�Y(F��]�~�t��օ�T��+<��2����������7!ǻ[uѻ�ۻ������5���a���	�
��E�i��8-������ �#%��0)��I-��S1�[O5��<9�=��@���D��pH��L�\�O�z\S�F�V�6pZ���]��^a���d�g*h�p�k���n�U"r�gu�-�x�X�{�}�6������SC��d҅�4_��ꈼ�r�������~���������3��s���X��A������~u��<h�����fW��Π�/D��Ĺ���.�����������������s��=筼�Z��Eΰ��A��j���,)�����?������w����o��8彼�  �  
�N=��M=�M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=Z�E=:�D=i-D=�jC=��B=`�A=\A=sX@=��?=��>=� >=�6==�k<=�;=b�:=V:=�19=�_8=~�7=i�6=��5= 5=�-4=�Q3=;s2=ܒ1=O�0=y�/==�.=��-=6-=+,=]-+=�8*=�@)=�E(=�G'=�E&=�@%=8$=�+#=9"=�!=o�=��=Ѱ=z�=�a=3=��=��=��=0I=e=��=�e=�=��=TT=�=��
=4	=Ơ=j'=1�=)&=h�=
 =[�<���<���<i�<r%�<���<��<�,�<"��<�b�<?��<i�<��<4��<w��<�s�<���<�O�<t��<�<�z�<1״<K0�<\��<�٩<Z*�<�x�<�Ğ<U�<�W�<+��<"�<�)�<n�<g��<M�<�mz<1�r<�xk<�c<^�\<7U<�M<�&F<h�><I7<�/<
y(<:!<
�<b<`<��<��;Mz�;:
�;��;Z�;��;V�;&ؔ;�Ԇ;�q;�V;�:;�S;�9;ϫ�:�S�:�P:��9�"�4�͹ݟL�����]�ʺ����CM��`.�(F���]�_�t�uօ�K���;��02������ڤ���!ǻSuѻ�ۻ��廷�ﻰ5���a����
��E�c��z-����� �l%��0)��I-��S1�nO5��<9��=���@�h�D��pH��L���O�r\S�I�V�GpZ���]�z^a���d�W*h�H�k���n�D"r��fu��x�,�{���/������bC��]҅�:_���鈼�r�������~���������9��x���z��6�������u��9h��!���oW��Π�*D�������.�����������������s��3筼�Z��>ΰ��A��e���)�����4������g����o��C彼�  �  �N=��M=M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=X�E=1�D=d-D=�jC=��B=Y�A=YA=qX@=��?=��>=� >=�6==�k<=#�;=h�:=\:=�19=�_8=��7=i�6=��5=(5=�-4=�Q3=?s2=�1=P�0=�/=A�.=��-==-=/,=c-+=�8*=�@)=�E(=�G'=�E&=�@%=8$=�+#=4"=�!=i�=��=Ͱ=v�=�a=3=��=��=��=)I=c=��=�e=�=��=YT=
�=��
=6	=Ҡ=q'=6�=,&=p�= =^�<���<���<i�<%�<���<���<{,�<��<�b�<9��<W�<��<4��<h��<�s�<���<�O�<d��<��<�z�<$״<L0�<G��<�٩<I*�<�x�<�Ğ<Z�<X�<3��<1�<�)�<n�<l��<T�<nz<C�r<�xk<�c<��\<KU<��M<'F<k�><7I7<3�/<+y(<J!<��<�a<@<��<���;Rz�;

�;ͩ�;�Y�;��;(�;�ה;�Ԇ;��q;oV;��:;S;�9;���:�R�:��P:��92��4�͹u�L�϶���ʺ�����L�`.��'F�W�]�"�t�,օ�J���;��2����������p!ǻ%uѻ)�ۻΤ�����5���a���
��E�y���-�+���� ��%��0)�J-��S1��O5�=9�=��@�v�D��pH��L�u�O�X\S�=�V�7pZ���]�x^a�^�d�C*h�;�k���n�)"r��fu��x��{���$��򱂼WC��S҅�C_���鈼�r������
���������I��}������=�������u��F*h������W��Π�:D�������.�����������������s��(筼�Z��8ΰ��A��\���)�����#������d����o��C彼�  �  �N=��M=�M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=N�E=/�D=V-D=�jC=t�B=O�A=TA=lX@=��?=��>=� >=�6==�k<=�;=d�:=]:=�19=`8=��7=q�6=��5=-5=�-4=�Q3=Js2=�1=^�0=|�/=H�.=��-=;-=5,=Z-+=�8*=�@)=�E(=�G'=�E&=�@%=8$=�+#=%"=�!=^�=��=ΰ=i�=�a=
3=��=��=��=*I=`=��=�e=�=��=_T=�=��
=F	=ؠ={'=B�=:&=y�= =w�<���<���<#i�<�%�<���<��<�,�<��<�b�<:��<W�<��<'��<[��<�s�<���<�O�<Z��<��<�z�<"״<60�<H��<�٩<O*�<�x�<�Ğ<V�<�W�<>��</�<*�<n�<n��<n�<-nz<t�r<yk<H�c<��\<{U<	�M<'F<��><7I7<E�/<y(<<!<�<�a<L<��<���;	z�;�	�;W��;�Y�;|�;��;�ה;=Ԇ;��q;�V;<�:;�R;_9;۪�:4R�:�P:��9��4�͹��L�ⴘ�+�ʺ����ZL��_.�H'F��]���t�օ�����;���1����������C!ǻquѻ�ۻ�����5���a��7�
��E�����-�X��2� �%�1)�J-�T1��O5�=9�=��@���D��pH��L�a�O�a\S�(�V�pZ���]�B^a�O�d� *h��k���n�"r��fu��x��{�M�$��󱂼YC��e҅�1_��ꈼ�r���������������W���������\������u��c,h��5����W�� Π�3D�������.������������������s��$筼�Z��ΰ��A��E���)��휶�������^����o��$彼�  �  �N=��M=M= aL=��K=��J=�*J=�lI=��H=��G=�0G=�pF=A�E=)�D=N-D=�jC=h�B=S�A=MA=bX@=��?=��>=� >=�6==�k<=�;=k�:=c:=�19=`8=��7=��6=��5=25=�-4=�Q3=Ts2=�1=m�0=��/=L�.=��-=:-=<,=Z-+=�8*=�@)=�E(=�G'=�E&=�@%=�7$=�+#="=�!=Z�=��=ð=^�=�a=�2=��=��=�=-I=]=��=�e=�=��=eT=�=��
=Y	=۠=�'=I�=D&=��=" =��<���<Ť�<+i�<�%�<��<��<�,�<��<�b�<'��<M�<��<��<d��<ms�<���<�O�<P��<��<�z�<#״<0�<F��<}٩<M*�<�x�<�Ğ<b�<X�<N��<*�<*�<n�<���<��<4nz<��r<yk<z�c<��\<�U<L�M<'F<��><0I7<b�/< y(<O!<�<�a<N<u�<���;�y�;�	�;P��;5Y�;F�;d�;�ה;�ӆ;�q;pV;��:;�R;�8;ڪ�:pQ�:��P:C�9u��4�͹/�L������ʺ����9L��_.��&F���]���t�օ�p���;���1������ʤ��!ǻvuѻ͠ۻ
��	��6��/b��m�
��E�����-�j��E� ��%�@1)��I-�8T1��O5�3=9�,=�
�@���D��pH��L�C�O�]\S��V�pZ���]��]a�J�d��)h���k�x�n��!r��fu���x��{�D���豂�JC��a҅�'_��ꈼ�r�����������Ƅ��O���������l������u��k*h��L����W��;Π�6D��ȹ���.��������������s��筼�Z��ΰ��A��-����(��֜����s���=����o��彼�  �  �N=��M=M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=?�E=�D=I-D=�jC=g�B=G�A=?A=_X@=��?=��>=� >=�6==�k<= �;=n�:=e:=�19=`8=��7=��6=��5=?5=�-4=�Q3=^s2=��1=i�0=��/=R�.=��-=E-=<,=_-+=�8*=�@)=�E(=�G'=�E&=�@%=�7$={+#="=�!=S�=��=��=]�=}a=�2=��=��=��=&I=^=��=�e=�=��=pT= �=Ą
=W	=�=�'=P�=K&=��=, =��<��<ͤ�<Ii�<�%�<��<���<�,�<��<�b�<-��<J�<{�<���<I��<ls�<���<�O�<:��<��<�z�<�ִ<0�<=��<}٩<@*�<�x�<�Ğ<\�<
X�<J��<A�<%*�<4n�<���<~�<gnz<��r<?yk<��c<ۆ\<�U<Y�M<D'F<ȶ><cI7<`�/</y(<M!<��<�a<2<{�<���;�y�;U	�;��;Y�;��;5�;(ה;�ӆ;2�q;zV;3�:;DR;�8;���:�P�:t�P:��9$6�4�͹;�L�������ʺ*����K��^.�{&F�S�]�h�t��Յ����1;���1��V���|���!ǻPuѻ�ۻ��K��.6��<b�#���
�3F�����-����]� ��%�G1)�<J-�VT1��O5�A=9�5=�)�@���D��pH��L�F�O�8\S���V��oZ�q�]�^a��d��)h��k�g�n��!r��fu���x���{�=���᱂�HC��Z҅�7_��ꈼ�r�����������݄��k���������u��!����u��tNh��Q����W��;Π�BD��չ���.���������񋩼����{s��筼�Z��ΰ��A������(��ʜ�����u���8���jo��彼�  �  �N=��M=
M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=9�E=�D=D-D=�jC=a�B=:�A=?A=[X@=z�?=��>=� >=�6==�k<=�;=o�:=b:=�19=`8=��7=��6=��5=D5=�-4=�Q3=\s2=�1=n�0=��/=U�.=��-=E-=:,=d-+=�8*=�@)=�E(=�G'=�E&=�@%=�7$=q+#="=�!=H�=��=��=Z�=qa=�2=��=��=�=#I=h=��=�e=�=��=sT=$�=̈́
=Z	=��=�'=a�=V&=��== =��<��<Ӥ�<Ni�<�%�<��<���<�,�<#��<�b�<2��<7�<p�<��<.��<cs�<���<�O�<!��<��<�z�<�ִ<0�<��<~٩<<*�<�x�<�Ğ<N�<X�<E��<G�<&*�<An�<���<��<�nz<��r<uyk<��c<�\<�U<h�M<f'F<˶><sI7<X�/<>y(<9!<�<�a<%<}�<��;�y�;,	�;���;�X�;x�;�;�֔;�ӆ;?�q;hV;�:;[Q;�8;���:�Q�:*�P:J�9z��48�͹Y�L�㴘�z�ʺB���K��^.� &F�g�]���t�OՅ�u�� ;���1��S�������*!ǻ-uѻO�ۻѤ�O��(6��Bb�_�|�
�aF����.������ ��%�W1)�oJ-�LT1��O5�Q=9�-=�9�@�u�D��pH��L�K�O�<\S���V��oZ�R�]�^a���d��)h���k�A�n��!r�Kfu���x���{�7���求�FC��W҅�<_���鈼�r������2�����ڄ���������������:����u���\h��P����W��9Π�ED��ʹ���.�����������������zs���歼Z���Ͱ�tA�� ����(��ǜ�����[���1���[o��彼�  �  "�N=��M=M=�`L=��K=��J=z*J=�lI=��H=��G=�0G=�pF=0�E=�D==-D=�jC=Y�B=7�A=<A=VX@=y�?=��>=� >=�6==�k<="�;=v�:=j:=�19=`8=��7=��6=��5=H5=�-4=�Q3=bs2=	�1=v�0=��/=[�.=��-=I-=A,=h-+=�8*=�@)=�E(=�G'=�E&=�@%=�7$=q+#="=�!=G�=��=��=P�=qa=�2=��=��=�= I=d=��=�e=�=��={T=-�=΄
=e	=��=�'=h�=_&=��=D =��<��<��<[i�<�%�<+��<��<�,�<��<�b�<$��<5�<i�<���<,��<Qs�<���<�O�<��<��<�z�<�ִ<0�<��<n٩<0*�<�x�<�Ğ<W�<X�<T��<L�<9*�<Dn�<���<��<�nz<��r<�yk<��c<�\<�U<~�M<g'F<�><~I7<w�/<Uy(<K!<�<�a<<X�<��;Vy�;	�;���;�X�;X�;��;�֔;5ӆ;�q;&V;��:;0Q;8;!��:�P�:h�P:N�9O�5��͹H�L�������ʺ�����J�o^.��%F�7�]�=�t�;Յ�8��;��`1�����f���� ǻuѻ4�ۻ���}��[6��Vb�i���
�cF�$��.������ �
	%��1)�rJ-�eT1��O5�`=9�G=�J�@���D��pH��L�-�O�*\S���V��oZ�U�]��]a���d��)h���k�%�n��!r�5fu���x���{�����ױ��6C��S҅�<_��ꈼ�r������5�����䄐����΄��������=����u���\h��Z����W��HΠ�QD��׹���.���������狩�����hs���歼xZ���Ͱ�sA������(���������M���'���[o��彼�  �   �N=��M=M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=,�E=�D=4-D=�jC=S�B=4�A=2A=SX@=|�?=��>=� >=�6==�k<= �;=l�:=g:=�19=`8=��7=��6=��5=T5=�-4=�Q3=ts2=�1=z�0=��/=`�.=��-=I-==,=_-+=�8*=�@)=�E(=�G'=�E&=�@%=�7$=l+#="=�!=>�=��=��=J�=oa=�2=��=��=�=+I=a=��=�e=�=��={T=2�=҄
=k	=��=�'=h�=f&=��=D =��<!��<���<Zi�<�%�<��<���<�,�<��<�b�<��<;�<i�<��<)��<Ds�<���<yO�<��<��<�z�<�ִ<�/�<&��<e٩<7*�<�x�<�Ğ<[�<X�<O��<K�<>*�<Ln�<���<��<�nz<%�r<ryk<��c<2�\<�U<��M<t'F<��><zI7<o�/<(y(<Q!<��<�a<&<C�<1��;y�;��;`��;oX�;:�;w�;{֔;ӆ;��q;wV;<�:;`Q;�7;	��:�P�:#�P:!�9N��4��͹�L�9�����ʺ|����J��].�F%F���]�*�t�2Յ����:��>1�����h���!ǻbuѻ�ۻ��;��R6��bb�T���
�xF�:��-.����� �	%��1)�J-��T1��O5�`=9�J=�#�@���D��pH��L�F�O�/\S���V��oZ�I�]��]a���d�v)h���k��n�k!r�;fu�m�x���{������ޱ��IC��[҅�:_��ꈼ�r������0������������܄��������H����u���jh��p����W��RΠ�ID��ι���.���������싩�����cs���歼kZ���Ͱ�hA��𴳼�(���������M������Uo���佼�  �  '�N=��M=M= aL=��K=��J=w*J=�lI=��H=��G=�0G=�pF=,�E=�D=3-D=�jC=T�B=0�A=3A=OX@=s�?=��>=� >=�6==�k<=$�;=u�:=o:=�19=`8=��7=��6=��5=S5=�-4=�Q3=rs2=�1=��0=��/=c�.=��-=P-=D,=g-+=�8*=�@)=�E(=�G'=�E&=�@%=�7$=h+#=	"=�!=;�=��=��=L�=ja=�2=��=��=�=#I=_=��=�e=�=��=T=6�=ׄ
=p	=�=�'=m�=g&=��=H =��<*��<���<di�<�%�</��<��<�,�<��<�b�<��<(�<]�<��<��<Fs�<���<vO�<��<��<�z�<�ִ<�/�<��<_٩<%*�<�x�<�Ğ<Z�<X�<\��<Z�<=*�<Rn�<���<��<�nz<�r<�yk<��c<<�\<U<��M<�'F<��><�I7<��/<My(<T!<��<�a<<9�<���;y�;��;H��;lX�;�;k�;P֔;ӆ;y�q;�V;��:;�P;Z7;ȧ�:�P�:��P:��9��5��͹
�L�Y���>�ʺ�����J��].�E%F��]�Q�t�&Յ�����:��%1�����1���� ǻ uѻ/�ۻ+��x�ﻥ6��xb�|���
��F�3��1.����� � 	%��1)��J-��T1��O5�~=9�p=�E�@���D��pH��L�&�O�\S���V��oZ�7�]��]a���d�)h���k�	�n�u!r�-fu�n�x���{������˱��5C��L҅�>_��ꈼ�r������D������������ۄ��������S����u���lh��n����W��XΠ�\D��Թ���.���������ߋ������cs���歼hZ���Ͱ�bA�������(���������C������No���佼�  �  �N=��M=aM=�ZL=j�K=��J=�!J=QcI=F�H=��G=�$G=�cF=��E=��D=�D=QZC=�B=��A=�
A=D@=|?=.�>="�====�Q<=
�;=�:=��9=9=�?8=k7=��6=~�5=��4=�4=�(3=-I2=Cg1=�0=��/=ӳ.=v�-=��,=��+=S�*=��)=n)=�	(=�	'=�&=��$=��#=��"=��!=�� =:�=M�=f=�?=�=3�=�=Rx=�:=�=S�=,e='=�="c=*=9�=Y4
=��=�Q=a�=&\=7�=�S=D��<Br�<�J�<��<���<S��<eZ�<�<���<W�<���<U��<��<��<�$�<m��<�<���<��<�m�<�ջ<:�<���<8��<�R�<7��<>��<�Q�<���<�<>�<r��<�ӏ<��<�d�<w��<��<�tz<<s<�k<od<��\<�>U<��M<�fF<~�><C�7<O70<��(<�!<�*<��<��<3L<;�;���;%O�;m��;g��;Œ�;'x�;Ip�;�}�;�@u;N�Y;�T>;�&#;,-;B��: ��:Kb:�W�9���8���� �9���F������T;��<)�Z�@��`X�Ȁo��)���l��#���8|���H����~kĻ�λ��ػ3��+�컯���� �[��`p	���Ԅ����S�,����#��(�&.,�U>0�x@4��48�<���?���C��G��8K��N���R�V���Y��%]���`�Pd�|wg���j�a0n��q�{�t��x�`N{�n�~�b܀��r����������'�����Y@���ɋ�/Q���֎�[���ݑ��^��ߔ��]��7ۗ��W��Ӛ��M��_ǝ�g@������<0��H����������	��s�������i���ޭ��S��tȰ�S=��Q���g'������C�����^����t��
콼�  �  �N=��M=bM=�ZL=k�K=��J=�!J=ScI=Q�H=��G=�$G=�cF=��E=��D=�D=VZC=�B=��A=�
A=D@=|?=.�>="�==�==�Q<=�;=�:=��9=9=�?8=k7=��6=��5=��4=�4=�(3=0I2=Cg1="�0=��/=ӳ.=q�-=�,=��+=R�*=��)=j)=�	(=�	'=�&=��$=��#=��"=��!=� =5�=G�=f=�?=�=-�=�=Zx=�:=z�=L�=0e='="�=$c=&=9�=X4
=��=�Q=e�=#\=8�=�S=J��<Xr�<�J�<��<���<_��<yZ�<!�<���<W�<���<U��<��<��<�$�<o��<��<���<��<�m�<�ջ<
:�<���</��<�R�<=��<=��<�Q�<���<$�<>�<���<�ӏ<��<�d�<���<��<�tz<Gs<��k<}d<�\<�>U<��M<�fF<s�><=�7<w70<��(<�!<�*<��<��<9L<��;j��;O�;f��;]��;���;�w�;rp�;�}�;�@u;�Y;�T>;h'#;'-;-��:z��:b:�W�9/��8�����9�?�����+��;��<)��@��`X���o��)���l�����>|���H����%kĻ
�λ��ػT��I�컷���� �9��rp	���������S�C��{�#��(�#.,�l>0�b@4�f48�<���?���C��G��8K���N���R�&V���Y��%]�֞`�Hd�mwg���j�^0n�ہq�m�t��x�qN{�q�~�h܀��r����������'�� ���\@���ɋ�Q���֎�[���ݑ�_���ޔ��]��<ۗ��W��#Ӛ��M��hǝ�R@������=0��R����������	��_�������i���ޭ��S��lȰ�X=��L���r'������G�����O����t��콼�  �  �N=��M=ZM=�ZL=m�K=��J=�!J=OcI=T�H=��G=�$G=�cF=��E=��D=�D=bZC=�B=��A=�
A=D@= |?=)�>=)�==�==�Q<=�;=�:=��9=9=�?8=k7=��6=w�5=��4=�4=�(3=-I2=8g1=�0=��/=ҳ.=t�-=|�,=��+=K�*=��)=i)=�	(=�	'=�&=��$=��#=��"=��!=
� =8�=I�=#f=�?=�=.�=�=Vx=�:=��=L�=6e= = �= c='=;�=P4
=��=�Q=`�=\=4�=�S=2��<Sr�<�J�<��<~��<T��<qZ�<�<���<W�<���<K��<��<��<�$�<��<��<���<��<�m�<�ջ<
:�<Κ�<-��<�R�<7��<H��<�Q�<���<*�<	>�<���<�ӏ<��<�d�<{��<��<�tz<Fs<�k<d<˭\<�>U<��M<�fF<��><6�7<p70<h�(<�!<�*<��<��<(L<��;]��;MO�;���;w��;��;�w�;�p�;�}�;Au;m�Y;�T>;�'#;�,;?��:���:Ab:�V�9W��8ق���9�^������O��;�0=)��@��`X�Ào�>*���l��L���>|���H����$kĻ@�λ��ػX���컪���� �3��qp	�m�������S�;��T�#��(��-,�g>0�_@4�s48�<���?���C��G��8K���N���R� V���Y��%]���`�td�|wg���j�h0n��q���t��x��N{�X�~�i܀��r����������'�����L@���ɋ�Q���֎�[���ݑ�
_���ޔ��]��/ۗ��W��#Ӛ��M��jǝ�M@������20��I����������	��_�������i���ޭ��S��vȰ�k=��L���w'������Z��&���S����t��콼�  �  �N=��M=_M=�ZL=h�K=��J=�!J=UcI=T�H=��G=�$G=�cF=��E=��D=�D=]ZC=�B=��A=�
A=D@=|?=/�>=(�==�==�Q<=�;=�:=��9=9=�?8=k7=��6=z�5=��4=�4=�(3=)I2=>g1=�0=��/=̳.=s�-=}�,=��+=O�*=��)=e)=�	(=�	'=�&=��$=��#=��"=��!=� ==�=N�=f=�?=�=/�=�=Xx=�:=��=H�=/e=#=�= c=%=2�=P4
=��=�Q=\�=\=-�=�S=8��<Cr�<�J�<��<z��<S��<nZ�<�<���<W�<���<T��<��<��<�$�<w��<��<���<��<�m�<�ջ<:�<͚�<8��<�R�<B��<E��<�Q�<x��<"�<>�<{��<�ӏ<��<�d�<s��<��<�tz<+s<�k<]d<ۭ\<�>U<��M<�fF<h�><2�7<`70<{�(<�!<�*<��<��<CL<��;���;HO�;���;���;��;*x�;�p�;�}�;�@u;��Y;�T>;�'#;N-;4��:���:Qb:�W�9~��8V����9��������2��;��<)���@��`X���o�
*���l��G���m|���H����NkĻ�λ��ػr��"�컬���� �1��hp	�w��������S�%��g�#��(�.,�`>0�T@4�h48�<���?���C�	�G��8K��N���R�#V���Y��%]��`�_d��wg���j��0n��q���t��x��N{���~�k܀��r����������'��%���M@���ɋ�Q���֎�[���ݑ� _���ޔ��]��+ۗ��W��Ӛ��M��^ǝ�N@������60��K����������	��j�������i���ޭ��S��tȰ�`=��Y���s'��Ĝ��Q��#���]����t��콼�  �  �N=��M=^M=�ZL=l�K=��J=�!J=[cI=R�H=��G=�$G=�cF=��E=��D=�D=_ZC=%�B=��A=�
A=D@=|?=4�>=&�====�Q<=�;=�:=��9=9=�?8=k7=��6=s�5=��4=�4=�(3=I2=8g1=�0=��/=ʳ.=o�-={�,=��+=N�*=��)=m)=�	(=�	'=�&=��$=��#=��"=��!=� =?�=Q�="f=�?=�=7�=�=]x=�:=��=O�=,e="=�=c=!=.�=P4
=x�=�Q=Q�=\='�=�S=)��</r�<�J�<��<w��<K��<fZ�<�<���<W�<���<\��<��<��<�$�<���<�<���<�<�m�<�ջ<':�<̚�<E��<�R�<O��<F��<�Q�<���<�<>�<v��<�ӏ<��<�d�<k��<s�<�tz<�s<�k<0d<ĭ\<�>U<��M<�fF<N�><6�7<S70<s�(<�!<�*<��<��<[L<��;���;XO�;���;���;��;rx�;�p�;[~�;|Au;�Y;JU>;�'#;�-;��:���:�b:�V�9���8����Q�9�-���������;�c=)��@��`X���o�6*��m��M���x|���H����gkĻ�λ��ػ/���컈���z �&��Gp	�z��������S���T�#��(��-,�?>0�I@4�Q48��<���?���C��G��8K��N���R�/V�ϣY��%]�#�`�sd��wg���j��0n��q���t��x�|N{���~�k܀��r����������'�����Q@���ɋ�Q���֎�[���ݑ��^���ޔ��]��&ۗ��W��Ӛ��M��Rǝ�P@������50��D����������	��o�������i���ޭ��S���Ȱ�l=��p���v'��ڜ��\��9���h����t�� 콼�  �  ��N=��M=\M=�ZL=l�K=��J=�!J=WcI=Y�H=��G=�$G=�cF=��E=��D=�D=iZC=�B=��A=A=D@=&|?=2�>=-�====�Q<=�;=�:=��9=9=�?8=k7=��6=o�5=~�4=�4=�(3=I2=5g1=�0=��/=ų.=n�-=s�,=��+=L�*=��)=j)=�	(=�	'=�&=��$=��#=��"=��!=� =F�=Y�=+f=�?=�==�="�=]x=�:=��=K�=/e==�=c==)�=E4
=u�=�Q=N�=\="�=�S=��<(r�<�J�<��<m��<:��<hZ�<�<���<W�<���<W��<��<"��<%�<���<�<Α�<�<�m�<�ջ< :�<ܚ�<W��<�R�<G��<U��<�Q�<���<#�<>�<s��<�ӏ<��<�d�<a��<s�<�tz<�s<��k<-d<��\<�>U<|�M<�fF<U�><�7<F70<i�(<�!<�*<��<��<LL<��;��;�O�;���;���;l��;�x�;q�;+~�;�Au;n�Y;�U>;"(#;�-;��:���:;b:LX�9ڼ�8����d�9����w���6��<�x=)��@��aX���o�E*��m�������|��I��PkĻ*�λ��ػF�����g���� ���$p	�c��������S����.�#��(��-,�!>0�7@4�O48��<���?���C��G��8K��N�ՂR�7V�ۣY�&]�'�`��d��wg���j��0n��q���t��x��N{���~�s܀�s����������'�����E@���ɋ�Q���֎��Z���ݑ��^���ޔ��]��ۗ��W��Ӛ��M��@ǝ�C@������&0��B����������	��r�������i���ޭ��S���Ȱ�o=��q����'��ۜ��_��<���p���u��콼�  �  ؏N=��M=YM=�ZL=k�K=��J=�!J=XcI=b�H=��G=�$G=dF=��E=��D=�D=sZC=&�B=�A=A=D@=.|?=2�>=0�==�==�Q<=�;=�:=��9=9=�?8=�j7=��6=h�5=y�4=�4=�(3=I2=*g1=�0=��/=��.=m�-=p�,=��+=F�*=��)=h)=�	(=�	'=�&= %=��#=��"=��!=� =J�=Z�=4f=�?=�=9�=&�=cx=�:=��=G�=,e==�=c==#�==4
=r�=�Q=L�=\=�=�S=��< r�<�J�<��<]��<<��<eZ�<�<���<W�<���<V��<��<#��<%�<���<�<��<
�<n�<ֻ<4:�<뚴<L��<�R�<J��<Y��<R�<���< �<>�<y��<�ӏ<��<�d�<X��<e�<dtz<�s<��k<d<��\<�>U<l�M<mfF<N�><��7<S70<]�(<�!<�*<��<��<NL< �;��;�O�; �;+��;���;�x�;vq�;u~�;JBu;��Y;�U>;�(#;�-;���:j��:�b:�V�9*��8���9�9����<���Y��u<��=)�a�@�
bX���o��*��'m�������|��I��+;kĻX�λ��ػR�����Y���m ����<p	�;����z���S����#��(��-,�1>0�%@4�548��<���?���C��G��8K� �N�ۂR�>V��Y�&]�0�`��d��wg��j��0n�'�q���t��x��N{���~��܀��r����������'�����=@���ɋ��P���֎��Z���ݑ��^���ޔ��]��ۗ�zW���Қ��M��Kǝ�3@������#0��>����������	��m�������i���ޭ��S���Ȱ��=��w����'��㜶�p��J���w���u��콼�  �  ؏N=��M=XM=�ZL=o�K=��J=�!J=`cI=d�H=��G=�$G=dF=��E=��D=�D=vZC=1�B=�A=
A=D@=/|?=9�>=.�====�Q<=�;=�:=��9=	9=�?8=k7=��6=^�5=o�4=�4=�(3=I2="g1=�0=��/=��.=e�-=n�,=��+=J�*=��)=n)=�	(=�	'=�&=	 %=��#=��"=��!=� =R�=b�=5f=�?=�=?�=)�=ex=�:=��=M�=,e==�=c==�=>4
=f�=�Q=?�=\=�=�S=���<	r�<�J�<��<S��<7��<\Z�<�<���<W�<���<_��<��<,��<%�<���<0�<��<�<n�<ֻ<B:�<<[��<�R�<\��<R��<R�<���< �<>�<r��<�ӏ<��<�d�<S��<O�<Btz<�s<��k<�d<w�\<e>U<Z�M<zfF<&�><��7<A70<X�(<�!<�*< �<��<pL<0�;��;�O�;^ �;p��;⓲;�x�;�q�;�~�;�Bu;��Y;/V>;�(#;=.;���:2��:Nb:UX�9p��8*���h�9����P���9���<�M>)���@��aX�Q�o��*��wm�������|��CI��2\kĻ4�λ��ػ�����c���X ����p	�0�v��o��hS�͡���#�s(��-,�>0�@4�*48��<���?���C��G��8K��N��R�[V���Y�&]�V�`��d��wg��j��0n�Q�q���t�x��N{���~��܀��r����������'�����A@���ɋ��P���֎��Z���ݑ��^���ޔ�s]���ڗ�nW���Қ��M��>ǝ�,@��u���*0��;����������	��t�������i���ޭ��S���Ȱ��=�������'���������]�������u��2콼�  �  ۏN=��M=XM=�ZL=l�K=��J=�!J=gcI=a�H=��G=�$G=dF=��E=��D=�D=vZC=2�B=�A=A=D@=/|?=A�>=/�====�Q<=�;=�:=��9=9=�?8=�j7=��6=b�5=m�4=�4=�(3=I2=+g1=��0=��/=��.=`�-=p�,=��+=K�*=��)=m)=�	(=�	'=�&= %=��#=��"=��!= � =W�=j�=7f=�?=�=I�=*�=fx=�:=��=M�=(e==�=c==�=64
=a�=�Q=4�=�[=	�=�S=���<�q�<xJ�<v�<V��<)��<XZ�<�<|��<W�<���<n��<��<8��<%�<���<4�<��<2�<n�<ֻ<I:�<���<w��<�R�<h��<^��<R�<���<�<	>�<d��<�ӏ<��<�d�<B��<Q�<Vtz<�s<��k<�d<~�\<j>U<3�M<XfF<	�><�7<%70<Y�(<�!<�*<�<��<�L<!�;���;P�;u �;���;;Wy�;�q�;�~�;�Bu;^�Y;�V>;�(#;�.;���:���:�b:�Y�9>��8A���=�9�n��]�����<�[>)�;�@�<bX��o��*���m��ш���|��fI��$�kĻ'�λ��ػ�����%���K �����o	�)�f��d��QS������#�`(��-,��=0�@4�!48��<���?���C��G��8K� �N���R�bV��Y�0&]�f�`��d�xg�:�j��0n�c�q���t�x��N{�φ~��܀�
s����������'�����D@��wɋ��P���֎��Z���ݑ��^���ޔ�^]���ڗ�jW���Қ�yM��!ǝ�2@��i���0��:����������	����������i���ޭ��S���Ȱ��=�������'�����|��Z�������&u��@콼�  �  ֏N=��M=TM=�ZL=o�K=��J=�!J=ecI=g�H=��G=�$G=dF=��E=��D= D=�ZC=8�B=�A=A=D@=4|?=@�>=2�====�Q<=��;=�:=��9=9=�?8=�j7=��6=U�5=d�4=�4=�(3=I2=g1=��0=��/=��.=]�-=k�,=��+=C�*=��)=o)=�	(=�	'=�&= %=��#=��"=��!=)� =Z�=l�=?f=�?=�=G�=.�=hx=�:=��=M�=)e==�=c=	=�=-4
=]�=�Q=/�=�[=�=|S=ߐ�<�q�<fJ�<o�<G��<!��<NZ�<�
�<���<W�<���<m��<��<8��< %�<���<@�<���<7�<+n�<"ֻ<Z:�<��<n��<�R�<e��<c��<R�<���<�<�=�<i��<�ӏ<��<�d�<9��<A�<tz<�s<\�k<�d<M�\<C>U<'�M<DfF<�><�7<*70<H�(<�!<�*<�<Đ<�L<P�;j��;AP�;� �;���;E��;ky�; r�;�;�Cu;��Y;�V>;P)#;�.;G��:׵�:�b:�V�9j��8Y�����9�R��������s=��>)�\�@��bX��o�+���m����� }��vI��D{kĻ`�λ��ػ��������D �����o	���N��A��DS������#�M(�-,��=0��?4�48��<���?���C�	�G��8K�$�N��R�uV��Y�O&]�r�`��d�xg�M�j��0n�~�q��t�x��N{�؆~��܀�s���������'�����=@��wɋ��P���֎��Z��wݑ��^���ޔ�Y]���ڗ�]W���Қ�mM��*ǝ�'@��m���0��6����������	��}�������i���ޭ��S���Ȱ��=�������'��
������m�������0u��:콼�  �  ϏN=��M=UM=�ZL=p�K=��J=�!J=fcI=p�H=��G=�$G=dF=��E=��D=�D=�ZC=2�B=�A=A=$D@=8|?=?�>=7�====�Q<=�;=�:=��9=9=�?8=�j7=��6=R�5=e�4=�4=�(3=
I2=g1=��0=��/=��.=\�-=f�,=��+=F�*=��)=l)=�	(=�	'=�&= %=��#=��"=��!=)� =_�=n�=Af=�?=�=F�=6�=hx=�:=��=I�=.e==�=c==�=*4
=`�=�Q=3�=�[= �=}S=Ր�<�q�<_J�<o�<=��<"��<QZ�<�<���<W�<���<k��<��<D��<"%�<���<3�<��<7�<=n�<ֻ<T:�<��<o��<�R�<g��<g��<R�<���<&�<>�<j��<xӏ<��<�d�<8��<E�<tz<�s<A�k<�d<C�\<F>U<+�M<*fF<�><Θ7<.70<K�(<�!<�*<��<Ԑ<�L<��;��;vP�;� �;���;���;dy�;4r�;�~�;�Cu;ܵY;.W>;�)#;�.;��:R��:b:�Y�9˹�8T�����9�+���������=��>)���@� cX���o�%+���m����� }��|I��gnkĻH�λ��ػ#�⻿�����@ �����o	���_��@��/S������#�`(�o-,��=0��?4�48��<���?���C��G��8K��N���R�}V�&�Y�W&]�a�`��d�xg�e�j�1n�v�q�-�t�x� O{�ֆ~��܀�s����������'�����2@��xɋ��P���֎��Z��uݑ��^���ޔ�Y]���ڗ�dW���Қ�^M��)ǝ�@��j���0��;����������	��{�������i���ޭ��S���Ȱ��=�������'��������k�������<u��:콼�  �  ӏN=��M=RM=�ZL=p�K=��J=�!J=gcI=j�H=��G=�$G=dF=ĢE=��D=D=�ZC=<�B=�A=A=&D@=3|?=B�>=7�==	==�Q<=�;=�:=��9=9=�?8=�j7={�6=S�5=_�4=�4=�(3=�H2=g1=�0=��/=��.=]�-=j�,=��+=F�*=��)=q)=�	(=
'=�&= %=��#=��"=��!=-� =b�=q�=Ef=�?=�=L�=3�=gx=�:=��=O�=(e==�=c=	=�=(4
=U�=�Q=(�=�[=��=uS=א�<�q�<_J�<j�<B��<��<DZ�< �<~��<W�<���<p��<��<F��<.%�<ģ�<G�<��<<�<<n�<,ֻ<g:�<��<|��<�R�<j��<p��<R�<���<�<�=�<\��<�ӏ<��<�d�<,��<8�<tz<us<>�k<�d<9�\<1>U<�M</fF<�><ޘ7<70<@�(<�!<�*<�<ܐ<�L<i�;���;�P�;� �;���;���;{y�;=r�;D�;�Cu;,�Y;^W>;W)#;	/;	��:K��:Qb:�Y�9E��87�����9�e��~������=�?)���@�cX�V�o�+���m��+���}��vI��F�kĻI�λ��ػ��⻨�����? �����o	���/��,��#S������#�2(�g-,��=0��?4�48��<�}�?���C�
�G��8K�>�N���R�sV�(�Y�]&]���`��d�0xg�l�j�"1n���q�%�t�=x��N{�܆~��܀�s��
�������'��	���2@��rɋ��P���֎��Z��oݑ��^���ޔ�T]���ڗ�SW���Қ�ZM��ǝ�@��h���0��1����������	����������i���ޭ��S���Ȱ��=�������'��������u�������9u��A콼�  �  ӏN=��M=XM=�ZL=n�K=��J=�!J=icI=m�H=��G=�$G=dF=ŢE=��D=D=�ZC=>�B=�A=A=)D@=7|?=E�>=,�==
==�Q<=�;=�:=��9=9=�?8=�j7=|�6=X�5=]�4=�4=�(3=�H2=g1=�0=��/=��.=S�-=k�,=��+=L�*=��)=p)=�	(=�	'=�&= %=��#=��"=��!=*� =c�=t�=Bf=�?=�=M�=2�=kx=�:=|�=N�=#e==	�=c=�=�=.4
=T�=�Q=!�=�[= �=pS=��<�q�<hJ�<W�<8��<��<LZ�<�<u��<W�<���<t��<��<H��<)%�<���<H�<��<A�<2n�<,ֻ<`:�< ��<���<�R�<o��<_��<R�<���<�<>�<\��<�ӏ<r�<�d�<3��<7�<tz<ds<]�k<�d<C�\<3>U<�M<FfF<��><ܘ7<70<W�(<�!<�*<�<��<�L<��;ү�;<P�;� �;���;h��;�y�;*r�;V�;�Cu;�Y;�W>;�)#;1/;���:o��:�b:bY�9:��8���û9�����������==�>?)���@��bX�ǃo��*���m������#}���I��@�kĻ�λ��ػ�������3 �����o	�	�<��;��S�}����#�<(��-,��=0��?4�48��<���?���C��G��8K�.�N��R��V�:�Y�E&]���`��d�Mxg�R�j�1n���q��t�=x��N{��~��܀�s���������'�����H@��oɋ��P���֎��Z��|ݑ��^���ޔ�O]���ڗ�SW���Қ�qM��ǝ�@��b���0��<����������	���������
j���ޭ��S���Ȱ��=�������'��������t�������.u��V콼�  �  ӏN=��M=RM=�ZL=p�K=��J=�!J=gcI=j�H=��G=�$G=dF=ĢE=��D=D=�ZC=<�B=�A=A=&D@=3|?=B�>=7�==	==�Q<=�;=�:=��9=9=�?8=�j7={�6=S�5=_�4=�4=�(3=�H2=g1=�0=��/=��.=]�-=j�,=��+=F�*=��)=q)=�	(=
'=�&= %=��#=��"=��!=-� =b�=q�=Ef=�?=�=L�=3�=gx=�:=��=O�=(e==�=c=	=�=(4
=U�=�Q=)�=�[=��=uS=ؐ�<�q�<_J�<k�<C��<��<DZ�<�<��<W�<���<p��<��<F��<.%�<ģ�<G�<��<<�<<n�<,ֻ<g:�<��<|��<�R�<j��<o��<R�<���<�<�=�<[��<�ӏ<��<�d�<,��<8�<tz<ts<>�k<�d<9�\<1>U<�M<0fF<�><ߘ7<70<@�(<�!<�*<�<ݐ<�L<j�;���;�P�;� �;���;���;{y�;=r�;D�;�Cu;*�Y;\W>;T)#;/;��:F��:Eb:{Y�9䰑8Q�����9�k���������=� ?)���@�cX�X�o�+���m��,���}��wI��F�kĻJ�λ��ػ��⻨�����? �����o	���0��,��#S������#�2(�g-,��=0��?4�48��<�}�?���C�
�G��8K�>�N���R�sV�(�Y�]&]���`��d�0xg�l�j�"1n���q�%�t�=x��N{�܆~��܀�s��
�������'��	���2@��rɋ��P���֎��Z��oݑ��^���ޔ�T]���ڗ�SW���Қ�ZM��ǝ�@��h���0��1����������	����������i���ޭ��S���Ȱ��=�������'��������u�������9u��A콼�  �  ϏN=��M=UM=�ZL=p�K=��J=�!J=fcI=p�H=��G=�$G=dF=��E=��D=�D=�ZC=2�B=�A=A=$D@=8|?=?�>=7�====�Q<=�;=�:=��9=9=�?8=�j7=��6=R�5=e�4=�4=�(3=
I2=g1=��0=��/=��.=\�-=f�,=��+=F�*=��)=l)=�	(=�	'=�&= %=��#=��"=��!=)� =_�=n�=Af=�?=�=F�=6�=hx=�:=��=I�=.e==�=c==�=*4
=a�=�Q=4�=�[= �=}S=Ր�<�q�<`J�<o�<>��<"��<RZ�<�<���<	W�<���<l��<��<D��<"%�<���<3�<��<7�<=n�<ֻ<T:�<��<o��<�R�<g��<g��<R�<���<%�<>�<j��<xӏ<��<�d�<8��<E�<tz<�s<A�k<�d<C�\<F>U<+�M<+fF<�><Θ7</70<L�(<�!<�*<��<Ԑ<�L<��;���;wP�;� �;���;���;dy�;3r�;�~�;�Cu;ٵY;+W>;�)#;�.;���:H��:�b:aY�9��8����Ż9�7���������=��>)���@�cX���o�'+���m�����!}��~I��hpkĻI�λ��ػ$��������@ �����o	���_��@��/S������#�`(�o-,��=0��?4�48��<���?���C��G��8K��N���R�}V�&�Y�W&]�a�`��d�xg�e�j�1n�v�q�-�t�x� O{�ֆ~��܀�s����������'�����2@��xɋ��P���֎��Z��uݑ��^���ޔ�Y]���ڗ�dW���Қ�^M��)ǝ�@��j���0��;����������	��{�������i���ޭ��S���Ȱ��=�������'��������k�������<u��:콼�  �  ֏N=��M=TM=�ZL=o�K=��J=�!J=ecI=g�H=��G=�$G=dF=��E=��D= D=�ZC=8�B=�A=A=D@=4|?=@�>=2�====�Q<=��;=�:=��9=9=�?8=�j7=��6=U�5=d�4=�4=�(3=I2=g1=��0=��/=��.=]�-=k�,=��+=C�*=��)=o)=�	(=�	'=�&= %=��#=��"=��!=)� =Z�=l�=?f=�?=�=G�=.�=hx=�:=��=M�=)e==�=c=	=�=-4
=]�=�Q=/�=�[=�=|S=���<�q�<gJ�<p�<H��<"��<OZ�<�
�<���<W�<���<m��<��<9��<!%�<���<@�<���<7�<+n�<"ֻ<Y:�<��<n��<�R�<e��<b��<
R�<���<�<�=�<h��<�ӏ<��<�d�<9��<A�<tz<�s<\�k<�d<N�\<D>U<(�M<EfF<�><�7<+70<I�(<�!<�*<�<Ő<�L<R�;k��;BP�;� �;���;E��;jy�;�q�;�;�Cu;��Y;�V>;J)#;�.;9��:ȵ�:�b:iV�9]��8������9�d��*������|=��>)�d�@��bX��o�+���m��
���}��yI��F|kĻa�λ��ػ��������E �����o	���O��A��DS������#�M(�-,��=0��?4�48��<���?���C�	�G��8K�$�N��R�uV��Y�O&]�r�`��d�xg�M�j��0n�~�q��t�x��N{�؆~��܀�s���������'�����=@��wɋ��P���֎��Z��wݑ��^���ޔ�Y]���ڗ�]W���Қ�mM��*ǝ�'@��m���0��6����������	��}�������i���ޭ��S���Ȱ��=�������'��
������m�������0u��:콼�  �  ۏN=��M=XM=�ZL=l�K=��J=�!J=gcI=a�H=��G=�$G=dF=��E=��D=�D=vZC=2�B=�A=A=D@=/|?=A�>=/�====�Q<=�;=�:=��9=9=�?8=�j7=��6=b�5=m�4=�4=�(3=I2=+g1=��0=��/=��.=`�-=p�,=��+=K�*=��)=m)=�	(=�	'=�&= %=��#=��"=��!= � =W�=j�=7f=�?=�=I�=*�=fx=�:=��=M�=(e==�=c==�=64
=b�=�Q=4�=�[=
�=�S=���<�q�<zJ�<w�<W��<+��<YZ�<�<}��<W�<���<o��<��<9��<%�<���<4�<��<2�<n�<ֻ<I:�<���<v��<�R�<h��<^��<R�<���<�<	>�<c��<�ӏ<��<�d�<A��<Q�<Vtz<�s<��k<�d<~�\<j>U<4�M<YfF<�><�7<&70<[�(<�!<�*<�<��<�L<$�;���;P�;v �;���;;Vy�;�q�;�~�;�Bu;Y�Y;�V>;�(#;�.;���:���:�b:vY�9���8����g�9����q�����<�e>)�D�@�EbX���o��*���m��Ո���|��iI��&�kĻ)�λ��ػ �����&���K �����o	�)�f��d��RS������#�`(��-,��=0�@4�!48��<���?���C��G��8K� �N���R�bV��Y�0&]�f�`��d�xg�:�j��0n�c�q���t�x��N{�φ~��܀�
s����������'�����D@��wɋ��P���֎��Z���ݑ��^���ޔ�^]���ڗ�jW���Қ�yM��!ǝ�2@��i���0��:����������	����������i���ޭ��S���Ȱ��=�������'�����|��Z�������&u��@콼�  �  ؏N=��M=XM=�ZL=o�K=��J=�!J=`cI=d�H=��G=�$G=dF=��E=��D=�D=vZC=1�B=�A=
A=D@=/|?=9�>=.�====�Q<=�;=�:=��9=	9=�?8=k7=��6=^�5=o�4=�4=�(3=I2="g1=�0=��/=��.=e�-=n�,=��+=J�*=��)=n)=�	(=�	'=�&=	 %=��#=��"=��!=� =R�=b�=5f=�?=�=?�=*�=ex=�:=��=M�=,e==�=c==�=>4
=g�=�Q=@�=\=�=�S=���<r�<�J�<��<T��<8��<]Z�<�<���<W�<���<`��<��<-��<%�<���<1�<��<�<n�<ֻ<B:�<<Z��<�R�<\��<Q��<R�<���< �<>�<q��<�ӏ<��<�d�<R��<O�<Btz<�s<��k<�d<x�\<e>U<[�M<{fF<'�><��7<C70<Z�(<�!<�*<�<��<rL<3�;��;�O�;_ �;p��;⓲;�x�;�q�;�~�;�Bu;�Y;(V>;�(#;5.;|��:��:#b:�W�9��8������9����g���P��	=�W>)���@��aX�Z�o��*��{m�������|��FI��4^kĻ7�λ��ػ!�����e���X ����p	�0�v��o��iS�͡���#�s(��-,�>0�@4�*48��<���?���C��G��8K��N��R�[V���Y�&]�V�`��d��wg��j��0n�Q�q���t�x��N{���~��܀��r����������'�����A@���ɋ��P���֎��Z���ݑ��^���ޔ�s]���ڗ�nW���Қ��M��>ǝ�,@��u���*0��;����������	��t�������i���ޭ��S���Ȱ��=�������'���������]�������u��2콼�  �  ؏N=��M=YM=�ZL=k�K=��J=�!J=XcI=b�H=��G=�$G=dF=��E=��D=�D=sZC=&�B=�A=A=D@=.|?=2�>=0�==�==�Q<=�;=�:=��9=9=�?8=�j7=��6=h�5=y�4=�4=�(3=I2=*g1=�0=��/=��.=m�-=p�,=��+=F�*=��)=h)=�	(=�	'=�&= %=��#=��"=��!=� =J�=Z�=5f=�?=�=9�=&�=cx=�:=��=G�=,e==�=c==#�==4
=r�=�Q=L�=\=�=�S=��<!r�<�J�<��<_��<>��<fZ�<�<���<W�<���<W��<��<#��<%�<���<�<��<
�<n�<ֻ<3:�<ꚴ<L��<�R�<I��<X��<R�<���<�<>�<x��<�ӏ<��<�d�<W��<e�<dtz<�s<��k<d<��\<�>U<m�M<nfF<O�><��7<T70<_�(<�!<�*<��<��<OL<#�;��;�O�;  �;,��;���;�x�;uq�;s~�;EBu;��Y;�U>;�(#;�-;���:U��:{b:�V�9���8���j�9���T���p��<��=)�k�@�bX���o��*��+m�������|��I��.>kĻZ�λ��ػT�����[���n ����<p	�<����z���S����#��(��-,�1>0�%@4�548��<���?���C��G��8K� �N�ۂR�>V��Y�&]�0�`��d��wg��j��0n�'�q���t��x��N{���~��܀��r����������'�����=@���ɋ��P���֎��Z���ݑ��^���ޔ��]��ۗ�zW���Қ��M��Kǝ�3@������#0��>����������	��m�������i���ޭ��S���Ȱ��=��w����'��㜶�p��J���w���u��콼�  �  ��N=��M=\M=�ZL=l�K=��J=�!J=WcI=Y�H=��G=�$G=�cF=��E=��D=�D=iZC=�B=��A=A=D@=&|?=2�>=-�====�Q<=�;=�:=��9=9=�?8=k7=��6=o�5=~�4=�4=�(3=I2=5g1=�0=��/=ų.=n�-=s�,=��+=L�*=��)=j)=�	(=�	'=�&=��$=��#=��"=��!=� =F�=Y�=+f=�?=�=>�="�=]x=�:=��=L�=/e==�=c==)�=E4
=v�=�Q=N�=\=#�=�S=��<)r�<�J�<��<n��<;��<iZ�<�<���<W�<���<X��<��<"��<	%�<���<�<Α�<�<�m�<�ջ< :�<ܚ�<W��<�R�<G��<T��<�Q�<���<"�<>�<r��<�ӏ<��<�d�<`��<r�<�tz<�s<��k<-d<��\<�>U<}�M<�fF<V�><�7<G70<k�(<�!<�*<��<��<ML<��;��;�O�;���;���;l��;�x�;q�;*~�;{Au;h�Y;�U>;(#;�-;��:���:b:�W�9k��8ކ����9��������M��!<��=)��@��aX���o�I*��m�������|��
I��RkĻ,�λ��ػH�����i���� ���$p	�d��������S����.�#��(��-,�!>0�8@4�P48��<���?���C��G��8K��N�ՂR�7V�ۣY�&]�'�`��d��wg���j��0n��q���t��x��N{���~�s܀�s����������'�����E@���ɋ�Q���֎��Z���ݑ��^���ޔ��]��ۗ��W��Ӛ��M��@ǝ�C@������&0��B����������	��r�������i���ޭ��S���Ȱ�o=��q����'��ۜ��_��<���p���u��콼�  �  �N=��M=^M=�ZL=l�K=��J=�!J=[cI=R�H=��G=�$G=�cF=��E=��D=�D=_ZC=%�B=��A=�
A=D@=|?=4�>=&�====�Q<=�;=�:=��9=9=�?8=k7=��6=s�5=��4=�4=�(3=I2=8g1=�0=��/=ʳ.=o�-={�,=��+=N�*=��)=m)=�	(=�	'=�&=��$=��#=��"=��!=� =?�=Q�="f=�?=�=7�=�=]x=�:=��=O�=,e="=�=c=!=.�=P4
=x�=�Q=R�=\=(�=�S=*��<0r�<�J�<��<x��<L��<gZ�<�<���<W�<���<]��<��<��<�$�<���<�<���<�<�m�<�ջ<':�<̚�<E��<�R�<N��<E��<�Q�<���<�<>�<u��<�ӏ<��<�d�<k��<s�<�tz<�s<�k<0d<ŭ\<�>U<��M<�fF<O�><7�7<T70<t�(<�!<�*<��<��<\L<��;���;YO�;���;���;��;qx�;�p�;Y~�;xAu;۳Y;CU>;�'#;�-;��:z��:�b:zV�9W��8部�{�9�B����������;�m=)�
�@��`X���o�:*��"m��Q���{|��I����ikĻ�λ��ػ1���컉���{ �&��Gp	�{��������S���T�#��(��-,�?>0�J@4�Q48��<���?���C��G��8K��N���R�/V�ϣY��%]�#�`�sd��wg���j��0n��q���t��x�|N{���~�k܀��r����������'�����Q@���ɋ�Q���֎�[���ݑ��^���ޔ��]��&ۗ��W��Ӛ��M��Rǝ�P@������50��D����������	��o�������i���ޭ��S���Ȱ�l=��p���v'��ڜ��\��9���h����t�� 콼�  �  �N=��M=_M=�ZL=h�K=��J=�!J=UcI=T�H=��G=�$G=�cF=��E=��D=�D=]ZC=�B=��A=�
A=D@=|?=/�>=(�==�==�Q<=�;=�:=��9=9=�?8=k7=��6=z�5=��4=�4=�(3=)I2=>g1=�0=��/=̳.=s�-=}�,=��+=O�*=��)=e)=�	(=�	'=�&=��$=��#=��"=��!=� ==�=N�=f=�?=�=/�=�=Xx=�:=��=H�=/e=$=�= c=%=2�=Q4
=��=�Q=\�=\=.�=�S=9��<Dr�<�J�<��<{��<T��<oZ�<�<���<W�<���<T��<��<��<�$�<x��<��<���<��<�m�<�ջ<:�<̚�<8��<�R�<A��<D��<�Q�<x��<"�<>�<z��<�ӏ<��<�d�<r��<��<�tz<*s<�k<]d<ܭ\<�>U<��M<�fF<i�><3�7<b70<|�(<�!<�*<��<��<DL<��;���;IO�;���;���;��;*x�;�p�;�}�;�@u;��Y;�T>;�'#;H-;&��:|��:2b:^W�9r��8����*�9��������C��;�=)���@��`X��o�*���l��J���p|���H����PkĻ�λ��ػs��#�컭���� �1��hp	�w��������S�%��g�#��(�.,�`>0�U@4�h48�<���?���C�	�G��8K��N���R�#V���Y��%]��`�_d��wg���j��0n��q���t��x��N{���~�k܀��r����������'��%���M@���ɋ�Q���֎�[���ݑ� _���ޔ��]��+ۗ��W��Ӛ��M��^ǝ�N@������60��K����������	��j�������i���ޭ��S��tȰ�`=��Y���s'��Ĝ��Q��#���]����t��콼�  �  �N=��M=ZM=�ZL=m�K=��J=�!J=OcI=T�H=��G=�$G=�cF=��E=��D=�D=bZC=�B=��A=�
A=D@= |?=)�>=)�==�==�Q<=�;=�:=��9=9=�?8=k7=��6=w�5=��4=�4=�(3=-I2=8g1=�0=��/=ҳ.=t�-=|�,=��+=K�*=��)=i)=�	(=�	'=�&=��$=��#=��"=��!=
� =8�=I�=#f=�?=�=.�=�=Vx=�:=��=L�=6e=!=!�=!c='=;�=Q4
=��=�Q=`�= \=5�=�S=2��<Tr�<�J�<��<~��<U��<rZ�<�<���<W�<���<K��<��<��<�$�<��<��<���<��<�m�<�ջ<
:�<Κ�<-��<�R�<6��<H��<�Q�<���<*�<	>�<���<�ӏ<��<�d�<z��<��<�tz<Es<�k<d<̭\<�>U<��M<�fF<��><7�7<q70<i�(<�!<�*<��<��<)L<��;^��;NO�;���;w��;��;�w�;�p�;�}�;Au;j�Y;�T>;�'#;�,;5��:���:+b:�V�9���8
�����9�j������[���;�6=)��@��`X�Ȁo�A*���l��N���@|���H����%kĻA�λ��ػY���컫���� �3��qp	�m�������S�<��T�#��(��-,�g>0�_@4�s48�<���?���C��G��8K���N���R� V���Y��%]���`�td�|wg���j�h0n��q���t��x��N{�X�~�i܀��r����������'�����L@���ɋ�Q���֎�[���ݑ�
_���ޔ��]��/ۗ��W��#Ӛ��M��jǝ�M@������20��I����������	��_�������i���ޭ��S��vȰ�k=��L���w'������Z��&���S����t��콼�  �  �N=��M=bM=�ZL=k�K=��J=�!J=ScI=Q�H=��G=�$G=�cF=��E=��D=�D=VZC=�B=��A=�
A=D@=|?=.�>="�==�==�Q<=�;=�:=��9=9=�?8=k7=��6=��5=��4=�4=�(3=0I2=Cg1="�0=��/=ӳ.=q�-=�,=��+=R�*=��)=j)=�	(=�	'=�&=��$=��#=��"=��!=� =5�=G�=f=�?=�=-�=�=Zx=�:={�=L�=0e='="�=$c=&=9�=X4
=��=�Q=e�=#\=8�=�S=K��<Yr�<�J�<��<���<_��<yZ�<!�<���<W�<���<U��<��<��<�$�<p��<��<���<��<�m�<�ջ<
:�<���<.��<�R�<=��<=��<�Q�<���<$�<>�<���<�ӏ<��<�d�<���<��<�tz<Gs<��k<}d<�\<�>U<��M<�fF<s�><=�7<w70<��(<�!<�*<��<��<:L<��;k��;O�;f��;^��;���;�w�;rp�;�}�;�@u;�Y;�T>;f'#;%-;(��:u��:b:�W�9̽�8#���Ʒ9�E������1��;��<)��@��`X���o��)���l�����?|���H����%kĻ�λ��ػU��I�컷���� �9��rp	���������S�C��{�#��(�#.,�l>0�b@4�f48�<���?���C��G��8K���N���R�&V���Y��%]�֞`�Hd�mwg���j�^0n�ہq�m�t��x�qN{�q�~�h܀��r����������'�� ���\@���ɋ�Q���֎�[���ݑ�_���ޔ��]��<ۗ��W��#Ӛ��M��hǝ�R@������=0��R����������	��_�������i���ޭ��S��lȰ�X=��L���r'������G�����O����t��콼�  �  ߋN=�M=�M=jTL=��K=?�J=vJ=3ZI=n�H=*�G=>G=�WF=��E=��D=D=�JC=�B=j�A=r�@=�0@=�g?=��>=��==I==�8<=j;=�:=s�9=��8= !8=�J7=)s6=��5=e�4=3�3=3=� 2=i=1=�W0=�o/={�.=��-= �,=ض+=��*=��)=��(=��'=V�&=��%=f�$=��#==�"=�!=�| =�a=�B=r=��=��=��=�f=/-=�=?�=�d=C=�=�p=!=Z�=�Q=T�	=
z==i�==3�=�=��<���<���<ݗ�<�b�<�%�<v��<���<�B�<��<���<�!�<(��<�B�<���<:M�<���<�C�<��<$(�<@��<���<la�<ð<p!�< }�<H֥<-�<���<CԚ<=%�<�t�<�<��<\�<u��<j�<izz<�s<X�k<�;d<��\<�kU<=N<;�F<�B?<p�7<6�0<D5)<m�!<_�<sN<�<��<3�;k��;��;UF�;�;O��;r�;s��;��;�x;"];��A;\�&;��;���:Y��:bir:�l
:�s9Gt����'���uv��t��q�eb$��
<��iS��~j�룀��⋻�����[����\��U���_2̻�cֻ~n໥S�&��Э�����c:����%W�����/�F����"���&��+�6/�A>3��87�d%;�e?���B�z�F�A\J�=N�"�Q��NU���X�$i\���_�_c�>�f�]3j��m��p�g9t��w��z��~�y����6��̓�a����C������?����$�������2�������:�������<��]����:�������3��C����)���������o������,���`���ds���骼{`���֭�M��Bð�n9��ï��*&��Ӝ�����犹�o��Wz�����  �  ыN=�M=�M=fTL=��K=7�J=zJ=@ZI=}�H=%�G=:G=�WF=��E=��D=D=�JC=u�B=e�A=l�@=�0@=�g?=��>=��==B==�8<=j;=�:=t�9=}�8= !8=�J7=1s6=��5=f�4=3�3=3=� 2=l=1=�W0=�o/=y�.=��-=�,=ܶ+=��*=��)=��(=��'=\�&=��%=o�$=��#=;�"=	�!=�| =�a=�B=v=��=��=��=�f=@-=�=?�=�d=F=�=q==R�=�Q=J�	=z==l�==3�=�=��<���<���<ڗ�<�b�<�%�<x��<���<�B�<���<���<"�<N��<�B�<���<5M�<���<�C�<��<)(�<=��<���<ga�<�°<�!�<<}�<Q֥<�,�<���<=Ԛ<3%�<�t�<�<��<�[�<p��<|�<nzz<�s<O�k<�;d<��\<�kU<=N< �F<�B?<8�7<I�0<95)<^�!<Z�<VN<<��<�3�;=��;���;
F�;��;l��;Q�;���;C�;ˊx;�];��A;��&;g�;Ȍ�:|��:�ir:�j
:t9�s��k�'��󅺵w��s�8q�Nb$��
<��iS��~j�ͣ���⋻#��������]��.����2̻�cֻ�n໸S����L�������:����ZW�����/�L����"���&��+�56/�->3�U87�D%;�e?���B�p�F�a\J�.N�B�Q�OU���X�Hi\�z�_��^c�0�f�a3j��m��p�F9t��w�G�z��~������6��̓�a����P������'����$�������2�������:������=��X����:��Ʒ���3��O����)���������|������1���k���Ys��ꪼ�`���֭�M��0ð�k9������/&��͜�����֊��n��ez�����  �  ͋N=�M=�M=gTL=��K=9�J=|J=3ZI=u�H="�G=GG=�WF=��E=��D=	D=�JC=v�B=o�A=w�@=0@=�g?=��>=��==?==�8<=j;=�:=w�9={�8=!8=�J7=0s6=��5=^�4=1�3=3=� 2=]=1=�W0=�o/=�.=��-=�,=�+=��*=��)=��(=��'=W�&=��%=i�$=��#=I�"=�!=} =�a=�B=�=��=��=��=�f=5-=�=E�=�d=J=
�=q==U�=�Q=D�	=z==h�==1�=�=��<���<���<��<�b�<�%�<~��<���<�B�<���<���<�!�<:��<�B�<���<LM�<���<�C�<��<1(�<M��<���<�a�<�°<}!�<"}�<P֥<-�<���<DԚ<-%�<�t�<�<��<�[�<e��<u�<@zz<�s<B�k<�;d<��\<�kU<,N<�F<�B?<)�7<b�0<15)<c�!<\�<ZN<<�<O3�;%��;0��;9F�;�;���;%�;���;N�;q�x;z];s�A;�&;��;e��:<��:�jr:Ij
:dv9�q����'�`�Qx��$s��q��b$��
<�jS��~j�F����⋻S����졻T���-]�������2̻�cֻ�n໌S�����������:�u��SW�����/�P����"��&��+�06/�C>3��87�a%;�L?���B�]�F�x\J�N�F�Q�OU���X�bi\�~�_�2_c�>�f�a3j��m�2�p�}9t���w�b�z�k~������6��̓�"a����V������@����$�������2��r����:��p���=��O����:�������3��V����)���������w������+���q���Js��ꪼo`���֭�M��7ð��9������5&��Μ���������v��iz�����  �  ΋N=�M=�M=kTL=��K=>�J=}J=:ZI=}�H=)�G=BG=�WF=��E=��D=D=�JC={�B=g�A=s�@=�0@=�g?=��>=��==A==�8<=	j;=�:=q�9={�8= !8=�J7=.s6=��5=h�4=+�3=�3=� 2=c=1=�W0=�o/=v�.=��-=�,=ܶ+=��*=��)=��(=��'=Y�&=��%=u�$=��#=@�"=�!=�| =�a=�B=|=��=��=��=�f=>-=�=H�=�d=J=�=�p==N�=�Q=G�	=z==k�==*�=�=��<���<���<ؗ�<�b�<�%�<q��<���<�B�<���<���<�!�<K��<�B�<���<:M�<���<�C�<��<.(�<I��<���<ua�< ð<�!�<3}�<Q֥<-�<���<JԚ</%�<�t�<�<��<�[�<k��<q�<bzz<�s< �k<~;d<��\<�kU<2N<�F<�B?<,�7<;�0<-5)<q�!<P�<pN<<��<�3�;a��;��;.F�;'�;���;t�;���;}�;�x;8];�A;��&;�;ލ�:���:�jr:�k
:�r9	u����'����w��=s躶q�b$�B<�sjS�~j�����⋻-���"�����/]��1����2̻�cֻ�n�dS���\������z:����EW�����/�>����"���&��+�%6/�>3�[87�U%;�<?���B�\�F�`\J�5N�J�Q�!OU���X�Qi\���_�_c�.�f�~3j� �m��p�l9t���w�R�z��~������6��̓�a����T������5����$�������2�������:��x����<��S����:�������3��K����)���������i������%���o���_s��ꪼ�`���֭�M��;ð�q9��į��F&��؜�����䊹�s��hz�����  �  ԋN=�M=�M=hTL=��K=?�J=tJ=@ZI=|�H=*�G=DG=�WF=��E=��D=D=�JC=��B=p�A=w�@=�0@=�g?=��>=��==F==�8<=j;=�:=r�9=��8=� 8=�J7='s6=��5=^�4='�3=�3=� 2=b=1=�W0=�o/=u�.=��-=�,=ڶ+=��*=��)=��(=��'=T�&=��%=n�$=��#=C�"=�!=�| =�a=�B={=��=��=��=�f=?-=�=A�=�d=E=�=�p==P�=�Q=G�	=z==^�==&�=�=��<���<���<͗�<�b�<�%�<p��<���<�B�<��<���<�!�<K��<�B�<���<FM�<���<�C�<*��<2(�<T��<���<za�<	ð<�!�<@}�<A֥<-�<���<BԚ<5%�<�t�<�<��<�[�<f��<Y�<Lzz<�s<=�k<b;d<��\<mkU<#N<�F<�B?<B�7<:�0<55)<f�!<V�<rN<�<��<�3�;p��;��;�F�;m�;���;��;���;��;��x;�];�A;��&;c�;ӌ�:8��:/jr:�k
:tt9�s���'�V􅺙w��t�r��b$�s<�7jS�-j����㋻,���)������\��;����2̻�cֻ�n່S�3��C������a:����W�����/�����"���&��+�6/�0>3�U87�_%;�U?���B�l�F�]\J�9N�7�Q�OU���X�Oi\���_�_c�_�f�|3j��m�=�p�~9t� �w�J�z��~������6��̓�a����H������/����$�������2��w����:��~����<��N���|:�������3��C����)���������l������.���j���bs���骼�`���֭�M��Sð�|9��կ��6&��朶��������z��fz�����  �  ʋN=�M=�M=iTL=��K=?�J=}J=@ZI=z�H=/�G=LG=�WF=��E=��D=D=�JC=��B=o�A=��@=�0@=�g?=��>=��==G==�8<=j;=�:=k�9=v�8=� 8=�J7='s6=��5=T�4=&�3=�3=� 2=_=1=�W0=�o/=p�.=��-=�,=۶+=��*=��)=��(=��'=[�&=��%=k�$=��#=I�"=�!=} =�a=�B=�=��=��=��=�f=@-=�=C�=�d=E=�=�p==J�=�Q=@�	=z==T�==%�=�=��<���<���<̗�<�b�<�%�<t��<���<�B�<��<���<�!�<G��<�B�<���<FM�<���<�C�<'��<<(�<\��<���<�a�<ð<�!�<A}�<S֥<-�<���<DԚ<3%�<�t�<�<��<�[�<b��<c�<6zz<qs<6�k<O;d<��\<�kU<"N<�F<�B?<�7<3�0<35)<i�!<]�<tN<<��<{3�;���;^��;hF�;�;���;��;��;��;��x;M];H�A;��&;{�;���:s��:�jr:�k
:�v9�v����'��zx���s��q�Lc$�v<�4jS��j�+����⋻N���K�����[]��0����2̻�cֻwnເS����5������>:�s��"W�����/�����"���&��+��5/�2>3�O87�H%;�L?���B�h�F�d\J�1N�f�Q�)OU��X�ei\���_�'_c���f�x3j��m�f�p�|9t��w�h�z��~������6��̓�a����G������-����$�������2��v����:��j����<��D���s:�������3��7����)���������n������+���k���as��ꪼ�`���֭�M��Hð��9��௳�:&�������z��yz�����  �  ɋN=�M=�M=hTL=��K=<�J=�J=BZI=��H=.�G=LG=�WF=��E=��D=D=�JC=��B=t�A=~�@=�0@=�g?=��>=��==C==�8<=j;=�:=o�9=y�8=� 8=�J7=!s6=��5=W�4=�3=�3=� 2=X=1=�W0=�o/=l�.=��-=�,=۶+=��*=��)=��(=��'=]�&=��%=x�$=��#=L�"=�!=} =�a=�B=�=��=�=��=�f=E-=�=E�=�d=G=�=�p==N�=�Q=;�	=�y==X�=�=�=�=��<��<���<Ǘ�<�b�<�%�<g��<���<�B�<���<���<"�<X��<�B�<���<QM�<���<�C�<)��<F(�<g��<���<�a�<ð<�!�<E}�<]֥<-�<���<DԚ<(%�<�t�<�<��<�[�<U��<N�<(zz<ws<��k<J;d<��\<UkU<N<ݢF<�B?<�7<<�0<5)<c�!<W�<hN<#<��<�3�;���;^��;�F�;��;��;��;K��;�;�x;];��A;W�&;��;m��:��:Nkr:�k
:Wr9�t����'���y���t�Ur�c$��<�kS�Jj�X���!㋻n���f�|���U]��(����2̻�cֻ�n�pS�������p��K:�d��W�����/�����"���&��+��5/�>3�987�A%;�??���B�_�F�s\J�6N�c�Q�OU��X�vi\���_�C_c�n�f��3j�0�m�T�p��9t�8�w�z�z��~������6��̓�a����P������(����$�������2��k����:��Y����<��:���i:�������3��<����)���������p������,���v���]s��ꪼ�`���֭�"M��^ð��9��ݯ��V&��𜶼����������z�����  �  ȋN= �M=�M=iTL=��K=B�J=J=AZI=��H=3�G=SG=�WF=��E=��D=*D=�JC=��B=�A=��@=�0@=�g?=��>=��==H==�8<=j;=�:=k�9=v�8=� 8=�J7=s6=��5=Q�4=�3=�3=� 2=S=1=�W0=�o/=f�.=��-=�,=ֶ+=��*=��)=��(=��'=\�&=��%=z�$=��#=R�"=#�!=} =b=�B=�=��=�=��=�f=?-=�=G�=�d=C=�=�p=
=G�=�Q=>�	=�y=�=N�=�=�=�=��<x��<���<���<�b�<�%�<b��<���<�B�<��<���<"�<N��<�B�<���<cM�<��<�C�<E��<R(�<c��<���<�a�<ð<�!�<A}�<V֥<-�<���<DԚ<0%�<�t�<�<��<�[�<\��<C�<zz<Vs<��k<,;d<��\<<kU<
N<�F<dB?<�7<)�0<*5)<g�!<\�<~N<<��<�3�;���;���;�F�;��;��;H�;:��;/�;��x;�];��A;*�&;��;U��:�:Xkr:~l
:ms9v����'�_����x���t躹r�^c$� <�kS��j�}���N㋻L���������b]��M����2̻�cֻtn�GS����7���h��9:�J���V����[/�߂���"���&��+��5/��=3�N87�E%;�5?���B�h�F�d\J�GN�j�Q�.OU�8�X�gi\���_�Z_c���f��3j�;�m�o�p��9t�B�w�m�z��~������6��̓�a����E������)����$�������2��X����:��b����<��.���m:�������3��0����)���������e������,���o���fs��ꪼ�`���֭�M��hð��9����T&����������������z�����  �  ɋN=��M=�M=gTL=��K=B�J=�J=LZI=��H=<�G=RG=�WF=��E=��D=,D=�JC=��B=y�A=��@=�0@=�g?=��>=��==I==�8<=j;=�:=b�9=v�8=� 8=�J7=s6=��5=L�4=�3=�3=� 2=X=1=�W0=�o/=d�.=��-=	�,=Ӷ+=��*=��)=��(=��'=e�&=��%=z�$=¶#=Q�"=#�!=} =b=�B=�=��=�=��=�f=E-=$�=D�=�d=B=
�=�p==E�=�Q=2�	=�y==E�=�=�=�=��<k��<���<���<�b�<�%�<a��<���<�B�<��<���<"�<Q��<�B�<���<ZM�<��<�C�<F��<V(�<v��<���<�a�<,ð<�!�<V}�<b֥<-�<���<AԚ<.%�<�t�<�<��<�[�<F��<G�<zz<0s<��k<;d<��\<LkU<�N<͢F<iB?<�7<�0<&5)<_�!<Z�<}N<%<��<�3�;	��;���;�F�;��;?��;[�;u��;[�;b�x;�];q�A;0�&;q�;T��:��:Xkr:Bl
:�t99z����'���Yy��qu�Zr��c$�R<��jS�]�j�Q���X㋻����������n]��g����2̻�cֻjn�_S껛������e��:�M���V����_/�����"���&��+��5/��=3�487�%;�>?���B�m�F�d\J�QN�|�Q�1OU�9�X��i\���_�F_c���f��3j�E�m���p��9t�Y�w���z��~������6��̓�a����B����������$�������2��a���z:��R����<��*���Z:�������3�� ����)���������g������/���q���us��ꪼ�`���֭�0M��cð��9������V&���������������z�����  �  N= �M=�M=fTL=��K=?�J=�J=FZI=��H=<�G=VG=�WF=��E=��D=%D=�JC=��B=��A=��@=�0@=�g?=��>=��==G==�8<=j;=�:=j�9=p�8=� 8=�J7=s6=��5=H�4=�3=�3=� 2=J=1=�W0=�o/=h�.=��-=�,=ڶ+=��*=��)=��(=��'=b�&=��%=~�$=��#=Z�"=&�!=} =b=�B=�=��=�=��=�f=A-=�=D�=�d=E=�=�p==C�=�Q=,�	=�y=�=F�=�=�=�=��<b��<���<���<�b�<�%�<g��<���<�B�<���<���<
"�<O��<�B�<���<pM�<��<�C�<=��<^(�<���<���<�a�<*ð<�!�<K}�<`֥<-�<���<CԚ<'%�<�t�<�<��<�[�<>��<4�<�yz<?s<Ҥk<;d<b�\< kU<�N<ɢF<lB?<��7<*�0<5)<Z�!<b�<uN<!<��<�3�;��;���;"G�;8�;r��;&�;���;��;*�x;�];u�A;_�&;%�;���::�lr:�k
:�x9�u���'�&��y���u�s��c$��<�kS�+�j�����z㋻���������y]��(����2̻�cֻ\n�`S껵�����T��$:�(���V�M��W/����T�"���&�v+��5/��=3�B87�)%;�<?���B�^�F�\J�6N�w�Q�7OU� �X��i\���_�_c���f��3j�a�m���p��9t�f�w���z��~������6��̓�'a����F����������$�������2��J���v:��<����<��!���G:�������3��#����)���������i������-���x���bs��#ꪼ�`���֭�8M��vð��9������j&���������������z�����  �  ��N=��M=�M=iTL=��K=A�J=�J=EZI=��H=:�G=VG=�WF=��E=��D=,D=�JC=��B=��A=��@=�0@=�g?=��>=��==E==�8<=j;=�:=i�9=g�8=� 8=�J7=s6=��5=K�4=�3=�3=� 2=D=1=�W0=�o/=]�.=��-=�,=ֶ+=��*=��)=��(=��'=f�&=��%=��$=��#=\�"=!�!=} =
b=�B=�=��=�=��=�f=E-=!�=J�=�d=E=�=�p==9�=�Q=*�	=�y=�=I�=�=	�=�=��<r��<���<���<�b�<�%�<[��<���<�B�<���<���<
"�<b��<�B�<���<vM�<��<�C�<J��<i(�<t��<���<�a�<%ð<�!�<J}�<n֥<-�<���<GԚ<!%�<�t�<�<��<�[�<H��<@�<�yz<Js<��k<;d<X�\<,kU<�N<��F<LB?<��7<&�0<5)<f�!<S�<~N<F<��<>4�;���;���;/G�;��;���;i�;���;E�;\�x;�];��A;�&;(�;��:���:3lr:%l
:fr9v��M�'�e���vz���t�.s��c$�t<��kS��j��/㋻�����������]��F����2̻�cֻ�n�)S껏������*��4:� ���V�n��9/��i�"���&�k+��5/��=3�.87� %;�!?���B�[�F�|\J�DN���Q�\OU�O�X��i\���_��_c���f��3j�d�m�~�p��9t�C�w���z��~������6��!̓�#a����O����������$��s����2��D����:��=����<�����\:�������3��(����)���������c������)���~���gs��0ꪼ�`��׭�-M��jð��9��񯳼}&���������������z����  �  ɋN=��M=�M=hTL=��K=B�J=�J=IZI=��H==�G=YG=�WF=��E=��D=0D=�JC=��B=��A=��@=�0@=�g?=��>=��==I==�8<=j;=�:=j�9=t�8=� 8=�J7=s6=��5=B�4=�3=�3=� 2=D=1=�W0=�o/=c�.=��-=�,=Ѷ+=��*=��)=��(=��'=e�&=��%=~�$=ö#=]�"=0�!=} =
b=�B=�=�=�=��=�f=C-=!�=E�=�d=?=�=�p=
=C�=�Q='�	=�y=�=?�=�=�=�=��<T��<���<���<�b�<�%�<Q��<���<�B�<���<���<"�<V��<�B�<���<yM�<��<�C�<O��<m(�<���<���<�a�<.ð<�!�<P}�<g֥<-�<���<@Ԛ<%%�<�t�<�<��<�[�<1��<.�<�yz<)s<��k< ;d<J�\<kU<�N<��F<iB?<�7<�0<
5)<`�!<P�<�N</<��<�3�;��;ц�;dG�;;�;���;��;���;��;��x;];��A;��&;Z�;��:J��:Ykr:�l
:no9�t����'����y��sv�ks�5d$��<��kS�~�j�餀��㋻����������C]��m����2̻�cֻon�ES껚������S��:����V�T��9/�ł�X�"�X�&�e+��5/��=3�887�%;�4?���B�o�F�n\J�\N�b�Q�1OU�7�X��i\��_��_c���f��3j�i�m���p��9t�~�w���z��~������6��*̓�a����D����������$��|����2��@���g:��;����<�����J:��t����3������)���������d������0���z���os��ꪼ�`���֭�EM��|ð��9�����q&��������#�������z�����  �  ��N=��M=�M=hTL=��K=D�J=�J=VZI=��H=E�G=WG=�WF=��E=��D=2D=�JC=��B=��A=��@=�0@=�g?=��>=��==O==�8<=	j;=�:=f�9=e�8=� 8=�J7=s6=��5=B�4=�3=�3=� 2=P=1=�W0=�o/=c�.=y�-=�,=϶+=��*=��)=��(=��'=h�&=��%=��$=ζ#=R�"=)�!=} =
b=�B=�=�=�=��=�f=L-=(�=B�=�d===
�=�p= =1�=�Q=/�	=�y=�=:�=�=�=�=��<X��<���<���<�b�<�%�<Y��<���<�B�<��<���<#"�<^��<�B�<���<dM�<��<�C�<R��<l(�<���<���<�a�<Bð<�!�<h}�<a֥<-�<���<>Ԛ<3%�<�t�<�<��<�[�<<��<:�<�yz<s<դk<�:d<b�\<1kU<�N<ʢF<(B?<��7<	�0<*5)<b�!<c�<�N<<�<�3�;S��;�;!G�;6�;���;��;���;��;�x;P];��A;��&;�;k��:#��:�kr:wm
:}u9,w����'����0y��6v躬r�3d$��<�ukS�ŀj������㋻������?����]������2̻�cֻ&n�TS껀������K���9�E���V�]��9/��d�"�r�&��+��5/��=3�87�%;�@?���B�y�F�]\J�aN���Q�xOU�C�X��i\��_�\_c���f��3j�k�m���p��9t�u�w���z��~������6��"̓�a����4����������$��w����2��V���n:��C����<�����L:�������3������)��z������d���{��2���k���ts��-ꪼ�`���֭�9M��pð��9��
���h&���������������z����  �  ɋN=��M=�M=hTL=��K=B�J=�J=IZI=��H==�G=YG=�WF=��E=��D=0D=�JC=��B=��A=��@=�0@=�g?=��>=��==I==�8<=j;=�:=j�9=t�8=� 8=�J7=s6=��5=B�4=�3=�3=� 2=D=1=�W0=�o/=c�.=��-=�,=Ѷ+=��*=��)=��(=��'=e�&=��%=~�$=ö#=]�"=0�!=} =
b=�B=�=�=�=��=�f=C-=!�=E�=�d=@=�=�p=
=C�=�Q='�	=�y=�=?�=�=�=�=��<U��<���<���<�b�<�%�<Q��<���<�B�<���<���<"�<V��<�B�<���<yM�<��<�C�<O��<m(�<���<���<�a�<-ð<�!�<O}�<g֥<-�<���<@Ԛ<$%�<�t�<�<��<�[�<1��<.�<�yz<)s<��k< ;d<J�\<kU<�N<��F<iB?<�7<�0<
5)<`�!<P�<�N</<��<�3�;��;ц�;dG�;;�;���;��;���;��;��x;];��A;��&;X�;��:F��:Pkr:�l
:Ho9u���'����y��xv�ms�8d$��<��kS���j�꤀��㋻����������C]��n����2̻�cֻpn�FS껛������S��:����V�T��9/�ł�X�"�X�&�e+��5/��=3�887�%;�4?���B�o�F�n\J�\N�b�Q�1OU�7�X��i\��_��_c���f��3j�i�m���p��9t�~�w���z��~������6��*̓�a����D����������$��|����2��@���g:��;����<�����J:��t����3������)���������d������0���z���os��ꪼ�`���֭�EM��|ð��9�����q&��������#�������z�����  �  ��N=��M=�M=iTL=��K=A�J=�J=EZI=��H=:�G=VG=�WF=��E=��D=,D=�JC=��B=��A=��@=�0@=�g?=��>=��==E==�8<=j;=�:=i�9=g�8=� 8=�J7=s6=��5=K�4=�3=�3=� 2=D=1=�W0=�o/=]�.=��-=�,=ֶ+=��*=��)=��(=��'=f�&=��%=��$=��#=\�"=!�!=} =
b=�B=�=��=�=��=�f=F-=!�=J�=�d=E=�=�p==9�=�Q=*�	=�y=�=J�=�=
�=�=��<s��<���<���<�b�<�%�<[��<���<�B�<���<���<"�<c��<�B�<���<vM�<��<�C�<J��<i(�<t��<���<�a�<%ð<�!�<J}�<n֥<-�<���<GԚ< %�<�t�<�<��<�[�<H��<@�<�yz<Js<��k<;d<X�\<-kU<�N<��F<MB?<��7<'�0<5)<g�!<S�<~N<F<��<?4�;���;���;/G�;��;���;i�;���;E�;Z�x;�];��A;�&;%�;���:���:"lr:l
:r9+v��_�'�n���z���t�3s��c$�x<��kS��j�𤀻1㋻�����������]��G����2̻�cֻ�n�)S껐������+��4:� ���V�n��9/��i�"���&�k+��5/��=3�.87� %;�!?���B�[�F�|\J�DN���Q�\OU�O�X��i\���_��_c���f��3j�d�m�~�p��9t�C�w���z��~������6��!̓�#a����O����������$��s����2��D����:��=����<�����\:�������3��(����)���������c������)���~���gs��0ꪼ�`��׭�-M��jð��9��񯳼}&���������������z����  �  N= �M=�M=fTL=��K=?�J=�J=FZI=��H=<�G=VG=�WF=��E=��D=%D=�JC=��B=��A=��@=�0@=�g?=��>=��==G==�8<=j;=�:=j�9=p�8=� 8=�J7=s6=��5=H�4=�3=�3=� 2=J=1=�W0=�o/=h�.=��-=�,=ڶ+=��*=��)=��(=��'=b�&=��%=~�$=��#=Z�"=&�!=} =b=�B=�=��=�=��=�f=A-=�=D�=�d=E=�=�p==C�=�Q=,�	=�y=�=F�=�=�=�=��<c��<���<���<�b�<�%�<h��<���<�B�<���<���<"�<P��<�B�<���<pM�<��<�C�<=��<^(�<���<���<�a�<)ð<�!�<J}�<_֥<-�<���<CԚ<&%�<�t�<�<��<�[�<>��<4�<�yz<?s<Ҥk<;d<b�\< kU<�N<ɢF<mB?<��7<+�0<5)<[�!<c�<vN<"<��<�3�;��;���;"G�;8�;r��;&�;���;��;'�x;�];q�A;[�&; �;���:㩭:�lr:�k
:6x9�u��9�'�3��y���u�s��c$��<��kS�0�j�����|㋻����������{]��)����2̻�cֻ]n�aS껶�����T��$:�)���V�M��W/����T�"���&�v+��5/��=3�B87�)%;�<?���B�^�F�\J�6N�w�Q�7OU� �X��i\���_�_c���f��3j�a�m���p��9t�f�w���z��~������6��̓�'a����F����������$�������2��J���v:��<����<��!���G:�������3��#����)���������i������-���x���bs��#ꪼ�`���֭�8M��vð��9������j&���������������z�����  �  ɋN=��M=�M=gTL=��K=B�J=�J=LZI=��H=<�G=RG=�WF=��E=��D=,D=�JC=��B=y�A=��@=�0@=�g?=��>=��==I==�8<=j;=�:=b�9=v�8=� 8=�J7=s6=��5=L�4=�3=�3=� 2=X=1=�W0=�o/=d�.=��-=	�,=Ӷ+=��*=��)=��(=��'=e�&=��%=z�$=¶#=Q�"=#�!=} =b=�B=�=��=�=��=�f=E-=$�=D�=�d=B=
�=�p==E�=�Q=2�	=�y==E�=�=�=�=��<k��<���<���<�b�<�%�<a��<���<�B�<��<���<"�<Q��<�B�<���<ZM�<��<�C�<F��<V(�<u��<���<�a�<,ð<�!�<V}�<a֥<-�<���<@Ԛ<-%�<�t�<�<��<�[�<F��<G�<zz<0s<��k<;d<��\<MkU<�N<͢F<jB?<�7<�0<'5)<`�!<[�<~N<&<��<�3�;
��;���;�F�;��;?��;[�;u��;Z�;_�x;�];m�A;+�&;k�;G��:��:;kr:$l
:>t9yz���'���iy���u�br��c$�Y<��jS�d�j�T���[㋻����������p]��i����2̻�cֻln�`S껜������f��:�N���V����`/�����"���&��+��5/��=3�487�%;�>?���B�m�F�d\J�QN�|�Q�1OU�9�X��i\���_�F_c���f��3j�E�m���p��9t�Y�w���z��~������6��̓�a����B����������$�������2��a���z:��R����<��*���Z:�������3�� ����)���������g������/���q���us��ꪼ�`���֭�0M��cð��9������V&���������������z�����  �  ȋN= �M=�M=iTL=��K=B�J=J=AZI=��H=3�G=SG=�WF=��E=��D=*D=�JC=��B=�A=��@=�0@=�g?=��>=��==H==�8<=j;=�:=k�9=v�8=� 8=�J7=s6=��5=Q�4=�3=�3=� 2=S=1=�W0=�o/=f�.=��-=�,=ֶ+=��*=��)=��(=��'=\�&=��%=z�$=��#=R�"=#�!=} =b=�B=�=��=�=��=�f=?-=�=G�=�d=D=�=�p==G�=�Q=>�	=�y=�=O�=�=�=�=��<y��<���<���<�b�<�%�<c��<���<�B�<��<���<"�<O��<�B�<���<dM�<��<�C�<E��<R(�<c��<���<�a�<ð<�!�<A}�<U֥<-�<���<CԚ</%�<�t�<�<��<�[�<\��<C�<zz<Vs<��k<,;d<��\<=kU<N<�F<eB?<�7<*�0<+5)<h�!<]�<N<<��<�3�;���;���;�F�;��;��;H�;9��;-�;��x;|];��A;$�&;��;F��:੭:8kr:\l
:�r9^v���'�q����x���t��r�fc$�(<�kS��j�����Q㋻O���������d]��O����2̻�cֻvn�HS����8���h��::�J���V����[/�߂���"���&��+��5/��=3�N87�E%;�5?���B�h�F�d\J�GN�j�Q�.OU�8�X�gi\���_�Z_c���f��3j�;�m�o�p��9t�B�w�m�z��~������6��̓�a����E������)����$�������2��X����:��b����<��.���m:�������3��0����)���������e������,���o���fs��ꪼ�`���֭�M��hð��9����T&����������������z�����  �  ɋN=�M=�M=hTL=��K=<�J=�J=BZI=��H=.�G=LG=�WF=��E=��D=D=�JC=��B=t�A=~�@=�0@=�g?=��>=��==C==�8<=j;=�:=o�9=y�8=� 8=�J7=!s6=��5=W�4=�3=�3=� 2=X=1=�W0=�o/=l�.=��-=�,=۶+=��*=��)=��(=��'=]�&=��%=x�$=��#=L�"=�!=} =�a=�B=�=��=�=��=�f=E-=�=E�=�d=G=	�=�p==N�=�Q=;�	=�y==X�= =�=�=��<���<���<ȗ�<�b�<�%�<h��<���<�B�<���<���<"�<Y��<�B�<���<RM�<���<�C�<)��<F(�<g��<���<�a�<ð<�!�<E}�<\֥<-�<���<CԚ<(%�<�t�<�<��<�[�<U��<M�<(zz<ws<��k<J;d<��\<VkU<N<ޢF<�B?<�7<=�0<5)<d�!<X�<iN<$<��<�3�;���;`��;�F�;��;��;��;J��;�;�x;];��A;P�&;��;^��:��:,kr:�k
:�q9�t����'���"y���t�]r�c$��<�kS�Qj�\���$㋻q���h�~���W]��*����2̻�cֻ�n�qS�������q��L:�e��W�����/�����"���&��+��5/�>3�987�A%;�??���B�_�F�s\J�7N�d�Q�OU��X�vi\���_�C_c�n�f��3j�0�m�T�p��9t�8�w�z�z��~������6��̓�a����P������(����$�������2��k����:��Y����<��:���i:�������3��<����)���������p������,���v���]s��ꪼ�`���֭�"M��^ð��9��ݯ��V&��𜶼����������z�����  �  ʋN=�M=�M=iTL=��K=?�J=}J=@ZI=z�H=/�G=LG=�WF=��E=��D=D=�JC=��B=o�A=��@=�0@=�g?=��>=��==G==�8<=j;=�:=k�9=v�8=� 8=�J7='s6=��5=T�4=&�3=�3=� 2=_=1=�W0=�o/=p�.=��-=�,=۶+=��*=��)=��(=��'=[�&=��%=k�$=��#=I�"=�!=} =�a=�B=�=��=��=��=�f=@-=�=C�=�d=F=�=�p==J�=�Q=@�	=z==T�==&�=�=��<���<���<͗�<�b�<�%�<u��<���<�B�<��<���< "�<H��<�B�<���<GM�<���<�C�<'��<<(�<\��<���<�a�<ð<�!�<@}�<S֥<-�<���<CԚ<3%�<�t�<�<��<�[�<a��<c�<6zz<qs<6�k<O;d<��\<�kU<"N<��F<�B?<�7<4�0<45)<j�!<_�<uN<<��<}3�;���;_��;iF�;��;���;��;��;��;��x;I];C�A;��&;t�;���:d��:�jr:�k
:Hv9�v����'�􅺌x���s��q�Tc$�~<�;jS��j�.����⋻Q���N�����]]��2����2̻�cֻxnແS����6������?:�s��"W�����/�����"���&��+��5/�2>3�O87�H%;�L?���B�h�F�d\J�1N�f�Q�)OU��X�ei\���_�'_c���f�x3j��m�f�p�|9t��w�h�z��~������6��̓�a����G������-����$�������2��v����:��j����<��D���s:�������3��7����)���������n������+���k���as��ꪼ�`���֭�M��Hð��9��௳�:&�������z��yz�����  �  ԋN=�M=�M=hTL=��K=?�J=tJ=@ZI=|�H=*�G=DG=�WF=��E=��D=D=�JC=��B=p�A=w�@=�0@=�g?=��>=��==F==�8<=j;=�:=r�9=��8=� 8=�J7='s6=��5=^�4='�3=�3=� 2=b=1=�W0=�o/=u�.=��-=�,=ڶ+=��*=��)=��(=��'=T�&=��%=n�$=��#=C�"=�!=�| =�a=�B={=��=��=��=�f=?-=�=B�=�d=E=�=�p==P�=�Q=G�	=z==^�==&�=�=��<���<���<Η�<�b�<�%�<q��<���<�B�<��<���<�!�<L��<�B�<���<FM�<���<�C�<*��<2(�<T��<���<za�<ð<�!�<@}�<@֥<-�<���<AԚ<4%�<�t�<�<��<�[�<f��<Y�<Lzz<�s<>�k<b;d<��\<nkU<$N<�F<�B?<C�7<;�0<65)<g�!<W�<sN<�<��<�3�;q��;��;�F�;m�;���;��;���;��;��x;�];
�A;��&;]�;ƌ�:*��:jr:�k
:�s9�s��5�'�f􅺨w��,t�r��b$�z<�>jS�3j����㋻/���+������\��=����2̻�cֻ�n້S�4��D������a:����W�����/�����"���&��+�6/�0>3�U87�_%;�U?���B�l�F�]\J�9N�7�Q�OU���X�Oi\���_�_c�_�f�|3j��m�=�p�~9t� �w�J�z��~������6��̓�a����H������/����$�������2��w����:��~����<��N���|:�������3��C����)���������l������.���j���bs���骼�`���֭�M��Sð�|9��կ��6&��朶��������z��fz�����  �  ΋N=�M=�M=kTL=��K=>�J=}J=:ZI=}�H=)�G=BG=�WF=��E=��D=D=�JC={�B=g�A=s�@=�0@=�g?=��>=��==A==�8<=	j;=�:=q�9={�8= !8=�J7=.s6=��5=h�4=+�3=�3=� 2=c=1=�W0=�o/=v�.=��-=�,=ܶ+=��*=��)=��(=��'=Y�&=��%=u�$=��#=@�"=�!=�| =�a=�B=|=��=��=��=�f=>-=�=H�=�d=J=�=�p==N�=�Q=G�	=z==l�==*�=�=��<���<���<ٗ�<�b�<�%�<r��<���<�B�<���<���<�!�<K��<�B�<���<;M�<���<�C�<��<.(�<H��<���<ua�< ð<�!�<3}�<Q֥<-�<���<JԚ<.%�<�t�<�<��<�[�<j��<q�<bzz<�s< �k<;d<��\<�kU<3N<�F<�B?<-�7<<�0<.5)<r�!<Q�<qN<<��<�3�;b��;��;/F�;(�;���;s�;���;|�; �x;5];�A;��&;�;Ӎ�:���:ojr:�k
:Jr9=u����'����w��Is躼q�#b$�G<�yjS��~j�����⋻/���$�����0]��2����2̻�cֻ�n�eS���]������z:����FW�����/�>����"���&��+�%6/�>3�[87�U%;�<?���B�\�F�`\J�5N�J�Q�!OU���X�Qi\���_�_c�.�f�~3j� �m��p�l9t���w�R�z��~������6��̓�a����T������5����$�������2�������:��x����<��S����:�������3��K����)���������i������%���o���_s��ꪼ�`���֭�M��;ð�q9��į��F&��؜�����䊹�s��hz�����  �  ͋N=�M=�M=gTL=��K=9�J=|J=3ZI=u�H="�G=GG=�WF=��E=��D=	D=�JC=v�B=o�A=w�@=0@=�g?=��>=��==?==�8<=j;=�:=w�9={�8=!8=�J7=0s6=��5=^�4=1�3=3=� 2=]=1=�W0=�o/=�.=��-=�,=�+=��*=��)=��(=��'=W�&=��%=j�$=��#=I�"=�!=} =�a=�B=�=��=��=��=�f=5-=�=E�=�d=J=
�=q==U�=�Q=D�	=z==h�==2�=�=��<���<���<��<�b�<�%�<~��<���<�B�<���<���<�!�<;��<�B�<���<LM�<���<�C�<��<1(�<M��<���<�a�<�°<}!�<!}�<P֥<-�<���<DԚ<-%�<�t�<�<��<�[�<d��<u�<?zz<�s<B�k<�;d<��\<�kU<-N<�F<�B?<*�7<c�0<25)<d�!<]�<[N<<�<P3�;&��;0��;9F�;�;���;%�;���;N�;o�x;w];p�A;�&;��;]��:4��:�jr:8j
:v9r����'�i�[x��-s��q��b$��
<�jS��~j�H����⋻U����졻U���/]�������2̻�cֻ�nໍS�����������:�u��SW�����/�Q����"��&��+�06/�C>3��87�a%;�L?���B�]�F�x\J�N�F�Q�OU���X�bi\�~�_�2_c�>�f�a3j��m�2�p�}9t���w�b�z�k~������6��̓�"a����V������@����$�������2��r����:��p���=��O����:�������3��V����)���������w������+���q���Js��ꪼo`���֭�M��7ð��9������5&��Μ���������v��iz�����  �  ыN=�M=�M=fTL=��K=7�J=zJ=@ZI=}�H=%�G=:G=�WF=��E=��D=D=�JC=u�B=e�A=l�@=�0@=�g?=��>=��==B==�8<=j;=�:=t�9=}�8= !8=�J7=1s6=��5=f�4=3�3=3=� 2=l=1=�W0=�o/=y�.=��-=�,=ܶ+=��*=��)=��(=��'=\�&=��%=o�$=��#=;�"=	�!=�| =�a=�B=v=��=��=��=�f=@-=�=?�=�d=F=�=q==R�=�Q=K�	=z==l�==3�=�=��<���<���<ڗ�<�b�<�%�<y��<���<�B�< ��<���<"�<O��<�B�<���<5M�<���<�C�<��<)(�<=��<���<ga�<�°<�!�<<}�<Q֥<�,�<���<=Ԛ<3%�<�t�<�<��<�[�<o��<|�<nzz<�s<O�k<�;d<��\<�kU<=N< �F<�B?<8�7<I�0<95)<^�!<[�<VN<<��<�3�;=��;���;F�;��;l��;Q�;���;C�;ʊx;�];��A;��&;e�;Č�:x��:�ir:�j
:�s9�s��t�'��󅺺w��s�;q�Pb$��
<��iS��~j�Σ���⋻$��������]��.����2̻�cֻ�n໸S����L�������:����ZW�����/�L����"���&��+�56/�->3�V87�D%;�e?���B�p�F�a\J�.N�B�Q�OU���X�Hi\�z�_��^c�0�f�a3j��m��p�F9t��w�G�z��~������6��̓�a����P������'����$�������2�������:������=��X����:��Ʒ���3��O����)���������|������1���k���Ys��ꪼ�`���֭�M��0ð�k9������/&��͜�����֊��n��ez�����  �  ��N=o�M=�M=|NL=�K=��J=uJ={QI=��H=��G=FG=�KF=�E=I�D=� D=�;C=�uB=��A=��@=�@=�S?=�>=ּ==��<=� <=-Q;=�:=P�9=@�8=�8=C,7==S6={x5=��4=`�3=��2=@�1=�1=z.0=.E/=\Y.=k-=!z,=l�+=��*=��)=�(=��'=��&=��%=�$= {#=Aj"=�U!=�= =G!=	=��=&�=E�=V=n =H�=��=Sd=b=��=j~=K(=�=�m=�	=��	=�2=��=�I=9�=CN=�� =w��<�h�<�F�<C�<@��<]��< o�<�&�<��<ـ�<$�<��<�W�<;��<�t�<o��<�|�<���<�q�<��<�U�<8·<�*�<^��<��<HR�<F��<�	�<Fb�<���<��<�`�<���<l�<gS�<���<T�<�z<ns<��k<6Wd<��\<�U<H8N<��F<p�?<�-8<�0<��)<5B"<��<8�<^�<|L<<�;e��;��;�|�;n\�;�M�;vQ�;�h�;I��;©{;�W`;�3E;H?*;~;���:81�:<�:`E:uZN94�H�#���z����K�ߺ���j���g7�ֹN���e���|�c}�����������L����o����ɻJ�ӻ�	޻������V��gi���n���9���m��s�G�!�s�%��*��;.�mI2�|I6�<:�">���A�'�E���I��AM���P���T�r'X���[��:_��b��*f�|�i���l�VWp��s���v��Cz��}�]a�����������+������Q��;ቼ�n��w���:���S��ܒ�����}������Ӟ�����m���P��4���[������K
��W��������v��m識�g���ߪ��W��+ϭ��F��>����5��O����$��蜶�������T�����i����  �  �N=n�M=�M=|NL=��K=��J=wJ=�QI=�H=��G=DG=�KF=��E=R�D=� D=�;C=�uB=��A=��@=�@=�S?=��>=׼==��<=!<=(Q;=�:=L�9=2�8=�8=:,7=<S6=�x5=�4=\�3=��2=D�1=�1=�.0=$E/=YY.=k-=z,=l�+=�*=��)=�(=��'=&=��%=�$=�z#=Dj"=�U!=�= =L!==��=�=G�=V=v =T�=��=Sd=b=��=c~=J(=t�=�m=�	=��	=�2=��=�I=/�==N=�� =���<�h�<�F�<J�<)��<P��<o�<�&�<��<Հ�<$�<��<X�<A��<�t�<j��<�|�<���<�q�<��<�U�<(·<�*�<W��<��<YR�<L��<�	�<Qb�<���<��<�`�<���<s�<bS�<���<g�<�z<ws<y�k<3Wd<�\<?�U<;8N<��F<��?<�-8<�0<��)<2B"<��<1�<g�<�L<|<�;T��;��;i|�;R\�;�M�;�Q�;�h�;��;��{;JW`;�3E;,@*;\~;���:�0�:���:GD:�TN94�H�{����z����i�ߺm���� h7���N�R�e�:�|�"}��В��ł���L��d��o����ɻ�ӻ�	޻������V��Ai���d��:���V��s�D�!���%��*��;.�LI2�LI6�<:�">�}�A�
�E���I��AM���P���T�u'X���[��:_��b��*f���i���l�DWp�̬s���v�$Dz�p�}�ta����������,�������Q��9ቼ�n��[���4���\���������r�����������~���P��<���D������F
��Z��������v��z識�g���ߪ��W��/ϭ��F��+����5��K���%��Ꜷ���|���[�����a����  �  �N=y�M=�M=|NL=�K=��J=yJ=wQI=�H=��G=NG=�KF=�E=S�D=� D=�;C=�uB=��A=��@=�@=�S?=�>=ݼ==��<=!<=&Q;=�:=W�9=0�8=�8=6,7==S6=yx5=�4=a�3=��2=H�1=|1=�.0= E/=_Y.=k-=z,=v�+=�*=��)=�(=��'=��&=��%=�$=�z#=Oj"=�U!=�= =J!=	=��=�=R�=V=r =K�=��=Td=]=��=]~=S(=x�=�m=�	=��	=�2=��=�I=1�=AN=�� =o��<�h�<zF�<\�<)��<b��<o�<�&�<"��<̀�<$�<���<X�<<��<�t�<|��<�|�<���<�q�<��<�U�<2·<�*�<V��<��<AR�<L��<�	�<Ob�<¸�<{�<�`�<���<��<cS�<���<c�<�z<�s<��k<EWd<��\<0�U<58N<��F<��?<�-8<5�0<~�)<3B"<��<%�<o�<jL<Z<�;J��;Q��;�|�;h\�;�M�;ZQ�;�h�;%��;(�{;�W`;3E;�?*;�};���:30�:�:�C:=XN9f�H����G�z�����1�ߺ���D���g7�p�N��e��|�}��뒔������L��Y񴻤o����ɻ��ӻ
޻�����W��Qi���4��:���^��s�5�!���%��*��;.�XI2�qI6�-<:��!>���A���E��I��AM���P���T�U'X���[��:_��b��*f���i���l�OWp��s���v�8Dz�K�}�sa����������,����Q��1ቼ�n��h���9���R��Β�����n�������������t���:��=���K������F
��\��������v���識�g���ߪ��W��/ϭ��F��/����5��A��� %������������]�����N����  �  �N=q�M=�M=�NL=�K=��J=|J=�QI=�H=��G=HG=�KF=�E=S�D=� D=�;C=�uB=��A=��@=�@=�S?=�>=߼==��<=!<=+Q;=�:=O�9=1�8=�8=7,7=@S6=wx5=�4=\�3=��2=C�1=}1=.0=#E/=WY.=k-=z,=n�+=�*=��)=�(=��'=Ɨ&=��%=�$={#=Dj"=�U!=�= =N!==��=!�=H�=V=w =S�=��=Wd=\=��=a~=K(=s�=�m=�	=��	=�2=��=�I=*�=;N=�� =k��<�h�<|F�<D�<"��<Q��<o�<�&�<��<΀�<$�<��<X�<F��<�t�<n��<�|�<���<�q�<��<�U�<.·<�*�<c��<��<SR�<U��<�	�<Fb�<˸�<}�<�`�<���<l�<[S�<���<Z�<�z<us<l�k<2Wd<��\<!�U<C8N<|�F<t�?<�-8<�0<z�)<GB"<��<2�<x�<�L<�<�;w��;"��;||�;�\�;�M�;�Q�;�h�;N��;ǩ{;�W`;�3E;;@*;)~;���:�0�:i��:/E:�TN9��H�����z�u���Ĉߺ ��B���g7�̺N�W�e�҄|�8}��ϒ��Ђ��M��f��o����ɻ��ӻ
޻���۶�V��:i�|�`��	:�ܲ�M��s�2�!���%��*��;.�CI2�NI6�<:��!>���A���E��I��AM���P���T�|'X���[��:_��b��*f���i���l�OWp���s���v�1Dz�x�}�ya����������,�������Q��-ቼ�n��Y���.���N��ܒ�����m�������������x���L��0���@������=
��U��������v���識�g���ߪ��W��7ϭ��F��8����5��K���%��霶�������V�����g����  �  �N=o�M=�M=|NL=�K=��J=tJ=�QI=�H=��G=LG= LF=�E=O�D=� D=�;C=�uB=��A=��@=�@=�S?=��>=׼==��<= !<=)Q;=�:=N�9=7�8=�8=7,7=3S6=tx5=ߛ4=X�3=��2==�1=�1=u.0=!E/=XY.=
k-=z,=j�+=�*=��)=�(=��'=��&=��%=�$={#=Gj"=�U!=�= =Q!==��=)�=I�=V=o =S�=��=Sd=a=��=a~=G(=x�=�m=�	=��	=�2=��=�I=*�=8N=�� =g��<�h�<zF�<A�<0��<T��<o�<�&�<��<ۀ�<$�<��<X�<:��<u�<r��<�|�<���<r�<��<�U�<;·<�*�<g��<��<ZR�<H��<�	�<Hb�<���<��<�`�<���<n�<[S�<���<K�<�z<_s<v�k<Wd<��\<�U<8N<��F<w�?<�-8<	�0<~�)<2B"<��<L�<[�<�L<^<�;|��;F��;�|�;�\�;�M�;	R�;�h�;o��;��{;X`;�3E;%@*;d~;���:�1�:F��:�D:TTN9ĜH�����z�h���U�ߺ%��Y��#h7���N���e���|��}��ᒔ�Ȃ���L��3�p����ɻ)�ӻ�	޻�����V��\i�q�S���9���A��s�D�!�b�%��*��;.�cI2�MI6�<:�">�~�A��E��I��AM���P���T�y'X���[��:_��b��*f���i���l�\Wp���s���v�2Dz�z�}�ja����������	,�������Q��<ቼ�n��]���9���G��ؒ�����|�������������k���B��,���O������J
��M��������v��~識�g���ߪ��W��6ϭ��F��G����5��V���%������������h�����e����  �  ߇N=r�M=�M=zNL=�K=��J={J=�QI=�H=��G=QG= LF=�E=W�D=� D=�;C=�uB=��A=��@=�@=�S?=��>=ݼ==��<=!<=&Q;=�:=R�9=*�8=�8=4,7=8S6=wx5=֛4=U�3=��2=6�1=y1=z.0=E/=TY.=k-=z,=n�+=�*=��)=�(=��'=ŗ&=��%=�$={#=Lj"=�U!=�= =U!==��=(�=L�=V=t =X�=��=Wd=^=��=]~=J(=r�=�m=�	=��	=�2=��=�I=*�=5N=�� =h��<�h�<rF�<7�<��<T��<o�<�&�<��<Ѐ�<$�<��<X�<A��<u�<y��<}�<���<�q�<��<V�<9·<�*�<i��<��<aR�<Q��<�	�<Kb�<���<~�<�`�<���<h�<SS�<���<R�<�z<?s<v�k< Wd<��\<�U<&8N<o�F<p�?<n-8<�0<{�)<-B"<��<=�<t�<�L<t<�;���;u��;�|�;�\�;N�;�Q�;�h�;���;/�{;SX`;�3E;Y@*;�~;���:*1�:���:.D:�WN9��H�����z�������ߺ������Qh7���N�!�e� �|�Z}��璔�₟�M��q��o����ɻ�ӻ�	޻�����tV��Ii�i�A���9�ʲ�0��s�#�!�e�%��*��;.�NI2�8I6�<:��!>���A��E��I��AM���P���T��'X���[��:_�"�b�+f���i���l�~Wp���s���v�>Dz���}��a����������,�������Q��0ቼ�n��W���1���@��В�����h�������������m���8��*���G������B
��P��������v���識�g���ߪ��W��>ϭ��F��?����5��f���%�����%������d�����h����  �  އN=q�M=�M=�NL=�K=��J=}J=�QI=�H=��G=SG=LF=�E=]�D=� D=�;C=�uB=��A=��@=�@=�S?=��>=�==��<=!<=(Q;=�:=O�9=,�8=�8=/,7=3S6=nx5=؛4=S�3=��2=:�1=v1=t.0=E/=RY.=k-=z,=n�+=�*=��)=�(=��'=ŗ&=��%=�$={#=Oj"=�U!=�= =V!==��=)�=Q�=V=y =V�=��=Vd=\=��=Z~=H(=n�=�m=�	=��	=�2=��=�I=!�=0N=�� =V��<�h�<iF�<;�<��<L��<o�<�&�<"��<ɀ�<$�<��<X�<K��<u�<���< }�<���< r�<�<V�<A·<+�<k��<��<[R�<W��<�	�<Ob�<θ�<p�<�`�<���<o�<MS�<���<F�<�z<Ks<Q�k<	Wd<��\<��U<8N<]�F<{�?<i-8<�0<[�)<EB"<��<,�<�<�L<�<�;���;���;�|�;�\�;AN�;R�;8i�;���;��{;TX`;D4E;�@*;�~;-��:�0�:x�:�D:eQN9W�H�u����z�/���)�ߺ{�����`h7��N���e�,�|��}���������M��z��o����ɻ��ӻ
޻�����V��)i�l�2���9����*�{s��!�]�%��*��;.�5I2�>I6�<:��!>���A���E��I��AM� �P���T��'X�ֵ[��:_�4�b��*f�Жi���l�tWp��s���v�NDz���}�~a����������,��鿆��Q��,ቼ�n��P���'���D��ǒ�����Z�������������f���4��(���4������;
��W��������v���識�g���ߪ��W��Dϭ��F��K����5��_���%������"������k�����b����  �  �N=o�M=�M={NL=�K=��J=~J=�QI=�H=��G=WG=
LF=�E=[�D=� D=�;C=�uB=��A=��@=�@=�S?=��>=�==��<= !<='Q;=�:=M�9=/�8=z8=/,7=1S6=jx5=֛4=P�3=��2=4�1=v1=o.0=E/=MY.=k-=z,=k�+=�*=��)=�(=��'=ȗ&=��%=�$=
{#=Tj"=�U!=�= =Z!==��=.�=V�= V=y =T�=��=Wd=]=��=[~=G(=o�=�m=�	=��	=�2=��=�I=�=-N=�� =N��<�h�<iF�<(�<��<H��<o�<�&�<��<Ԁ�<$�<��<X�<O��<u�<���<}�<���<r�<�<V�<R·<
+�<v��<��<ZR�<[��<�	�<Hb�<���<x�<�`�<���<b�<DS�<���<<�<�z</s<I�k<�Vd<��\<�U<8N<P�F<Y�?<z-8<�0<n�)<-B"<��<L�<��<�L<�<�;���;���;
}�;�\�;5N�;RR�;i�;���;�{;�X`;z4E;�@*;�~;Z��:�1�:���:E:�UN9N�H�����z�#���W�ߺ�������h7�;�N�)�e�#�|��}���������M��d��o����ɻ�ӻ
޻���¶�V��0i�\����9�����^s��!�I�%��*�s;.�6I2�AI6��;:��!>���A��E��I��AM���P���T��'X�˵[��:_�9�b�+f�ٖi���l��Wp�"�s���v�JDz���}�wa����������,�������Q��+ቼ�n��T���"���:���������d�������������T���,�����:������8
��H��������v���識�g���ߪ��W��Mϭ��F��U����5��m���%��
���%������n�����s����  �  ��N=h�M=�M=zNL=�K=��J={J=�QI=�H= �G=TG=LF=�E=b�D=� D=�;C=�uB=��A=��@=�@=�S?=�>=ܼ==��<= !<=&Q;=�:=I�9=+�8=u8=.,7=,S6=lx5=Λ4=I�3=��2=*�1=s1=k.0=E/=HY.=�j-=z,=f�+=�*=��)=�(=��'=ɗ&=��%=!�$={#=Oj"=�U!=�= =\!==��=1�=Q�=!V=| =]�=��=Sd=`=��=]~=A(=i�=�m=�	=��	=�2=��=�I=�='N=�� =R��<vh�<cF�<�<��<=��<o�<�&�<
��<׀�<$�<#��<X�<U��<u�<���<}�<���<r�<�<V�<M·<+�<{��<��<uR�<S��<�	�<Nb�<���<��<�`�<���<]�<@S�<���<8�<jz<s<U�k<�Vd<��\<�U<�7N<I�F<M�?<o-8<��0<{�)<*B"<��<J�<u�<�L<�<�;���;���;�|�;-]�;lN�;TR�;bi�;��;��{;�X`;�4E;�@*;k;���:2�:���:�D:�VN9��H�j���z�5����ߺ���Q���h7��N���e�G�|��}�����8���+M����p����ɻ�ӻ�	޻��绸��<V��i�P�.���9�����^s���!�<�%��*�k;.�'I2�I6��;:��!>�x�A��E��I��AM��P�ȏT��'X�ֵ[�;_�:�b�=+f�ܖi���l��Wp��s��v�RDz���}��a����������,�������Q��3ቼ�n��J������9��Ò�����T����������}��Y���4�����5������@
��L��������v��識�g���ߪ��W��Qϭ��F��Y����5��}���%�����1������y�����x����  �  ۇN=p�M=�M={NL=�K=��J=}J=�QI=�H=��G=^G=LF=�E=g�D=� D=�;C=�uB=��A=��@=�@=�S?=��>=�==��<=!<=$Q;=�:=O�9='�8=}8=+,7='S6=ex5=Λ4=I�3=��2=1�1=n1=i.0=E/=OY.=k-=z,=m�+=�*=��)=�(=��'=Ɨ&=��%=!�$={#=\j"=�U!=�= =^!==��=0�=]�=#V={ =V�=��=Vd=`=��=W~=E(=k�=�m=�	=��	=�2=z�=�I=�=$N=�� =?��<lh�<]F�<.�<��<J��<o�<�&�<��<Ӏ�<$�<��<X�<S��<u�<���<}�<���<r�<�<V�<T·<+�<{��<��<gR�<V��<�	�<Sb�<¸�<r�<�`�<���<`�<ES�<z��<1�<[z<&s<1�k<�Vd<��\<͕U<�7N<L�F<[�?<^-8<�0<a�)<.B"<��<H�<��<�L<�<�;���;��;-}�; ]�;�N�;AR�;�i�;���;D�{;Y`;�4E;�@*;;n��:�1�:}�:�D:OTN9ØH�D����z�t���x�ߺ���A���h7�t�N�P�e���|��}��+������M�����o����ɻ�ӻ�	޻���Ѷ�yV��i�L�����9�����^s��!�?�%�~*�d;.�(I2�5I6�<:��!>�v�A��E��I��AM��P�ďT��'X��[�;_�V�b�'+f��i���l��Wp�:�s��v�\Dz���}��a����������,��񿆼�Q��+ቼ�n��P������2���������I����������{��R��������4������=
��K��������v���識�g���ߪ��W��Lϭ��F��`����5��q���'%�����7������������q����  �  ӇN=n�M=�M=�NL=�K=��J=�J=�QI=�H=�G=[G=LF=�E=k�D=� D=�;C=�uB=��A=��@=�@=T?=��>=�==��<=!<=)Q;=�:=J�9=�8=x8=$,7=1S6=ex5=͛4=H�3=��2=1�1=i1=q.0=E/=JY.=�j-=z,=j�+=�*=��)=�(=��'=͗&=��%=,�$={#=\j"=�U!=�= =c!=#=��=/�=_�= V=� =^�=��=]d=Z=��=V~=B(=c�=�m=�	=��	=�2=u�=�I=�=!N=�� =;��<�h�<MF�<!�<���<;��<�n�<�&�<��<̀�<)$�<��<(X�<`��<u�<���<	}�<���<r�<!�<V�<Y·<+�<}��<��<fR�<g��<�	�<Jb�<͸�<l�<�`�<}��<V�<9S�<}��<<�<Iz<%s<��k<�Vd<��\<ݕU<�7N<4�F<F�?<;-8<�0<S�)<CB"<��<N�<��<�L<=�;���;ɭ�;D}�;]�;�N�;tR�;�i�;Д�;��{;�X`;!5E;�A*;�~;t��:�1�: �:�E:3QN9U�H�'����z�J���(�ߺ���U��i7��N�I�e��|��}��>���*���WM�����o����ɻ��ӻ
޻��绔��VV���h�T�����9������Fs��!�A�%�u*�n;.��H2�I6��;:��!>���A���E��I��AM�"�P��T��'X���[��:_�g�b�)+f��i�
�l��Wp�@�s���v�zDz���}��a������Ǖ��,�������Q��ቼ�n��<������8���������?����������{��M���"�����������,
��E��������v���識�g���ߪ��W��Xϭ��F��T����5��q���@%�����?������x�����{����  �  ߇N=k�M=�M=NL=�K=��J=zJ=�QI=�H=�G=[G=LF=�E=f�D=� D=�;C=�uB=��A=��@=�@=�S?=��>=ܼ==��<=!<=+Q;=�:=J�9=*�8={8=$,7=&S6=ax5=ɛ4=G�3=��2=.�1=h1=g.0=E/=LY.= k-=z,=g�+=�*=��)=�(=��'=ŗ&=��%=#�$={#=Yj"=�U!=�= =`!=!=��=9�=\�=#V=| =Y�=��=Td=_=��=[~=?(=j�=�m=�	=}�	=�2=t�=�I=�=!N=�� =4��<jh�<KF�<(�<��<?��<�n�<�&�<��<׀�<$�<��<X�<W��<u�<���<}�<���<r�<�<#V�<g·<+�<���<��<kR�<Q��<�	�<Mb�<ȸ�<u�<�`�<���<a�<=S�<l��<,�<Az<s<&�k<�Vd<��\<ĕU<�7N<<�F<Z�?<j-8<��0<a�)<=B"<��<R�<r�<�L<�<�;
��;Э�;k}�;Q]�;�N�;bR�;�i�;/��;��{;
Y`;5E;A*;#;$��:Y2�:���:^F:nQN9��H�5��6�z�B�����ߺ �����i7���N�v�e���|��}��`������!M��{�p����ɻ��ӻ�	޻���׶�aV��i�B����9������Ns��!��%��*�`;.�"I2�)I6�<:��!>�w�A��E�	�I��AM��P�ƏT��'X��[�;_�l�b�8+f���i��l��Wp�M�s��v�}Dz���}��a������ɕ��,�������Q��/ቼ�n��J������2���������H����������r��?���$�����/������B
��I��������v���識�g���ߪ��W��Sϭ��F��d����5��u���,%�����B������������q����  �  ؇N=i�M=�M=wNL=�K=��J={J=�QI=
�H=	�G=^G=LF=�E=h�D= D=�;C=�uB=��A=��@=�@=�S?=�>=ݼ==��<=� <=&Q;=�:=H�9="�8=p8=),7=%S6=jx5=͛4=@�3=��2=*�1=p1=h.0=E/=HY.=�j-=z,=f�+=�*=��)=#�(=��'=̗&=��%= �$={#=Uj"=�U!=�= =f!=*=��=3�=V�=.V=| =`�=��=Vd=g=��=[~=?(=h�=�m=�	=��	=�2=|�=�I=�=N=�� =F��<fh�<UF�<�<���<;��<�n�<�&�<��<��<$�<0��<X�<\��<'u�<���<}�<���<-r�<�<V�<X·<+�<���<��<�R�<W��<�	�<Tb�<���<|�<�`�<���<E�<>S�<t��<3�<Xz<�s<�k<�Vd<��\<֕U<�7N<C�F<"�?<Q-8<��0<l�)<B"<��<m�<y�<�L<�<�;/��;��;)}�;(]�;�N�;�R�;�i�;
��;�{;jY`;"5E;�@*;�;%��:;3�:���::E:SN96�H�j����z�������ߺ���G��ui7���N���e�y�|��}��;���8����M����p����ɻH�ӻ�	޻��绠��V��i�����9������+s��!�0�%��*�4;.�#I2�I6��;:��!>�V�A�'�E�	�I��AM��P���T��'X��[�;_�I�b�?+f��i��l��Wp�'�s��v�hDz���}��a������ƕ��,������Q��0ቼ�n��I������ ���������O���w������~��N��� �����8��n���<
��<��������v���識�g���ߪ��W��Rϭ��F��]����5������7%��%���:�����������������  �  ߇N=k�M=�M=NL=�K=��J=zJ=�QI=�H=�G=[G=LF=�E=f�D=� D=�;C=�uB=��A=��@=�@=�S?=��>=ܼ==��<=!<=+Q;=�:=J�9=*�8={8=$,7=&S6=ax5=ɛ4=G�3=��2=.�1=h1=g.0=E/=LY.= k-=z,=g�+=�*=��)=�(=��'=ŗ&=��%=#�$={#=Yj"=�U!=�= =`!=!=��=9�=\�=#V=| =Y�=��=Td=_=��=[~=?(=j�=�m=�	=}�	=�2=t�=�I=�="N=�� =4��<kh�<KF�<(�<��<?��<�n�<�&�<��<׀�<$�<��<X�<W��<u�<���<}�<���<r�<�<#V�<g·<+�<���<��<kR�<Q��<�	�<Mb�<Ǹ�<u�<�`�<���<a�<=S�<l��<,�<Az<s<&�k<�Vd<��\<ĕU<�7N<=�F<[�?<j-8<��0<b�)<>B"<��<S�<r�<�L<�<�;
��;Э�;k}�;Q]�;�N�;bR�;�i�;/��;��{;	Y`;5E;A*;!;!��:U2�:���:WF:QQN9��H�<��=�z�E�����ߺ"�����i7���N�w�e���|��}��a������!M��|�p����ɻ��ӻ�	޻���׶�bV��i�B����9������Ns��!��%��*�`;.�"I2�)I6�<:��!>�w�A��E�	�I��AM��P�ƏT��'X��[�;_�l�b�8+f���i��l��Wp�M�s��v�}Dz���}��a������ɕ��,�������Q��/ቼ�n��J������2���������H����������r��?���$�����/������B
��I��������v���識�g���ߪ��W��Sϭ��F��d����5��u���,%�����B������������q����  �  ӇN=n�M=�M=�NL=�K=��J=�J=�QI=�H=�G=[G=LF=�E=k�D=� D=�;C=�uB=��A=��@=�@=T?=��>=�==��<=!<=)Q;=�:=J�9=�8=x8=$,7=1S6=ex5=͛4=H�3=��2=1�1=i1=q.0=E/=JY.=�j-=z,=j�+=�*=��)=�(=��'=͗&=��%=,�$={#=\j"=�U!=�= =c!=#=��=/�=_�= V=� =^�=��=]d=Z=��=V~=B(=c�=�m=�	=��	=�2=u�=�I=�=!N=�� =;��<�h�<MF�<!�<���<<��<�n�<�&�<��<̀�<)$�<��<(X�<`��<u�<���<	}�<���<r�<!�<V�<Y·<+�<}��<��<eR�<g��<�	�<Jb�<͸�<l�<�`�<}��<V�<8S�<}��<<�<Iz<%s<��k<�Vd<��\<ݕU<�7N<4�F<G�?<;-8<�0<S�)<CB"<��<O�<��<�L<=�;���;ʭ�;D}�;]�;�N�;tR�;�i�;Д�;��{;�X`;5E;�A*;�~;n��:�1�:�:�E:�PN9��H�5���z�Q���/�ߺ���X��i7��N�L�e��|��}��?���+���XM�����o����ɻ��ӻ
޻��绕��VV���h�T�����9������Fs��!�A�%�u*�n;.��H2�I6��;:��!>���A���E��I��AM�"�P��T��'X���[��:_�g�b�)+f��i�
�l��Wp�@�s���v�zDz���}��a������Ǖ��,�������Q��ቼ�n��<������8���������?����������{��M���"�����������,
��E��������v���識�g���ߪ��W��Xϭ��F��T����5��q���@%�����?������x�����{����  �  ۇN=p�M=�M={NL=�K=��J=}J=�QI=�H=��G=^G=LF=�E=g�D=� D=�;C=�uB=��A=��@=�@=�S?=��>=�==��<=!<=$Q;=�:=O�9='�8=}8=+,7='S6=ex5=Λ4=I�3=��2=1�1=n1=i.0=E/=OY.=k-=z,=m�+=�*=��)=�(=��'=Ɨ&=��%=!�$={#=\j"=�U!=�= =^!==��=0�=]�=#V={ =V�=��=Vd=`=��=W~=E(=k�=�m=�	=��	=�2=z�=�I=�=%N=�� =?��<mh�<]F�<.�<	��<K��<o�<�&�<��<Ԁ�<$�<��<X�<T��<u�<���<}�<���<r�<�<V�<T·<+�<{��<��<gR�<V��<�	�<Sb�<¸�<q�<�`�<���<`�<ES�<z��<1�<Zz<&s<1�k<�Vd<��\<͕U<�7N<M�F<\�?<^-8<�0<b�)</B"<��<I�<��<�L<�<�;���;��;-}�; ]�;�N�;AR�;�i�;ߔ�;B�{;Y`;�4E;�@*;;f��:�1�:t�:~D:TN9�H�X����z�~�����ߺ���E���h7�x�N�T�e���|��}��,������M�����o����ɻ�ӻ�	޻���Ҷ�zV��i�M�����9�����^s��!�?�%�~*�d;.�(I2�5I6�<:��!>�v�A��E��I��AM��P�ďT��'X��[�;_�V�b�'+f��i���l��Wp�:�s��v�\Dz���}��a����������,��񿆼�Q��+ቼ�n��P������2���������I����������{��R��������4������=
��K��������v���識�g���ߪ��W��Lϭ��F��`����5��q���'%�����7������������q����  �  ��N=h�M=�M=zNL=�K=��J={J=�QI=�H= �G=TG=LF=�E=b�D=� D=�;C=�uB=��A=��@=�@=�S?=�>=ܼ==��<= !<=&Q;=�:=I�9=+�8=u8=.,7=,S6=lx5=Λ4=I�3=��2=*�1=s1=k.0=E/=HY.=�j-=z,=f�+=�*=��)=�(=��'=ɗ&=��%=!�$={#=Oj"=�U!=�= =\!==��=1�=Q�=!V=| =]�=��=Sd=`=��=]~=A(=j�=�m=�	=��	=�2=��=�I=�=(N=�� =S��<wh�<dF�<�<��<>��<o�<�&�<��<׀�<$�<#��<X�<U��<u�<���<}�<���<r�<�<V�<M·<+�<{��<��<tR�<S��<�	�<Mb�<���<��<�`�<���<\�<@S�<���<8�<jz<s<U�k<�Vd<��\<�U<�7N<J�F<M�?<o-8<��0<|�)<+B"<��<J�<u�<�L<�<�;���;���;�|�;-]�;lN�;TR�;ai�;��;��{;�X`;�4E;�@*;f;���:	2�:���:�D:hVN9�H������z�A����ߺ���V���h7�$�N���e�L�|��}�����:���,M����p����ɻ�ӻ�	޻��绹��=V��i�Q�.���9�����^s���!�<�%��*�k;.�'I2�I6��;:��!>�x�A��E��I��AM��P�ȏT��'X�ֵ[�;_�:�b�=+f�ܖi���l��Wp��s��v�RDz���}��a����������,�������Q��3ቼ�n��J������9��Ò�����T����������}��Y���4�����5������@
��L��������v��識�g���ߪ��W��Qϭ��F��Y����5��}���%�����1������y�����x����  �  �N=o�M=�M={NL=�K=��J=~J=�QI=�H=��G=WG=
LF=�E=[�D=� D=�;C=�uB=��A=��@=�@=�S?=��>=�==��<= !<='Q;=�:=M�9=/�8=z8=/,7=1S6=jx5=֛4=P�3=��2=4�1=v1=o.0=E/=MY.=k-=z,=k�+=�*=��)=�(=��'=ȗ&=��%=�$=
{#=Tj"=�U!=�= =Z!==��=.�=V�= V=y =T�=��=Xd=]=��=[~=G(=p�=�m=�	=��	=�2=��=�I=�=-N=�� =O��<�h�<iF�<)�<��<I��<o�<�&�<��<Հ�<$�<��<X�<P��<u�<���<}�<���<r�<�<V�<R·<
+�<u��<��<YR�<Z��<�	�<Hb�<���<w�<�`�<���<a�<CS�<���<<�<z</s<I�k<�Vd<��\<�U<8N<Q�F<Z�?<z-8<�0<o�)<.B"<��<M�<��<�L<�<�;���;���;}�;�\�;5N�;QR�;i�;���;�{;�X`;v4E;�@*;�~;O��:�1�:|��:�D:AUN9��H�����z�0���d�ߺ�������h7�A�N�/�e�(�|��}���������M��f��o����ɻ�ӻ
޻���¶�V��0i�\����9�����^s��!�J�%��*�s;.�6I2�AI6��;:��!>���A��E��I��AM���P���T��'X�˵[��:_�9�b�+f�ٖi���l��Wp�"�s���v�JDz���}�wa����������,�������Q��+ቼ�n��T���"���:���������d�������������T���,�����9������8
��H��������v���識�g���ߪ��W��Mϭ��F��U����5��m���%��
���%������n�����s����  �  އN=q�M=�M=�NL=�K=��J=}J=�QI=�H=��G=SG=LF=�E=]�D=� D=�;C=�uB=��A=��@=�@=�S?=��>=�==��<=!<=(Q;=�:=O�9=,�8=�8=/,7=3S6=nx5=؛4=S�3=��2=:�1=v1=t.0=E/=RY.=k-=z,=n�+=�*=��)=�(=��'=ŗ&=��%=�$={#=Oj"=�U!=�= =V!==��=*�=Q�=V=y =V�=��=Vd=\=��=Z~=H(=n�=�m=�	=��	=�2=��=�I=!�=0N=�� =V��<�h�<jF�<<�<��<M��<o�<�&�<#��<ɀ�<$�<��<X�<K��<u�<���< }�<���< r�<�<V�<A·<+�<k��<��<[R�<W��<�	�<Ob�<͸�<o�<�`�<���<n�<MS�<���<E�<�z<Ks<Q�k<	Wd<��\<��U<8N<]�F<|�?<j-8<�0<\�)<FB"<��<-�<��<�L<�<�;���;���;�|�;�\�;AN�;R�;7i�;���;��{;QX`;@4E;�@*;|~;!��:�0�:k�:�D:�PN9ǚH����éz�=���6�ߺ������fh7�$�N���e�1�|��}�����򂟻M��|��o����ɻ��ӻ

޻�����V��)i�l�2���9����*�{s��!�]�%��*��;.�6I2�>I6�<:��!>���A���E��I��AM� �P���T��'X�ֵ[��:_�4�b��*f�Жi���l�tWp��s���v�NDz���}�~a����������,��鿆��Q��,ቼ�n��P���'���D��ǒ�����Z�������������f���4��(���4������;
��W��������v���識�g���ߪ��W��Dϭ��F��K����5��_���%������"������k�����b����  �  ߇N=r�M=�M=zNL=�K=��J={J=�QI=�H=��G=QG= LF=�E=W�D=� D=�;C=�uB=��A=��@=�@=�S?=��>=ݼ==��<=!<=&Q;=�:=R�9=*�8=�8=4,7=8S6=wx5=֛4=U�3=��2=6�1=y1=z.0=E/=TY.=k-=z,=n�+=�*=��)=�(=��'=ŗ&=��%=�$={#=Lj"=�U!=�= =U!==��=(�=L�=V=t =X�=��=Wd=^=��=]~=J(=r�=�m=�	=��	=�2=��=�I=*�=5N=�� =i��<�h�<sF�<7�<��<U��<o�<�&�<��<р�<$�<��<X�<B��<u�<y��<}�<���<�q�<��<V�<9·<�*�<i��<��<aR�<P��<�	�<Jb�<���<~�<�`�<���<h�<SS�<���<R�<�z<?s<v�k< Wd<��\<�U<&8N<o�F<q�?<o-8<�0<|�)<.B"<��<>�<u�<�L<v<�;���;v��;�|�;�\�;N�;�Q�;�h�;���;-�{;PX`;�3E;U@*;�~;���:1�:���:D:iWN9�H� ��˪z�������ߺ������Wh7���N�'�e��|�]}��钔�䂟�M��r��o����ɻ�ӻ�	޻�����uV��Ji�i�A���9�ʲ�1��s�#�!�f�%��*��;.�NI2�8I6�<:��!>���A��E��I��AM���P���T��'X���[��:_�"�b�+f���i���l�~Wp���s���v�>Dz���}��a����������,�������Q��0ቼ�n��W���1���@��В�����h�������������m���8��*���G������B
��P��������v���識�g���ߪ��W��>ϭ��F��?����5��f���%�����%������d�����h����  �  �N=o�M=�M=|NL=�K=��J=tJ=�QI=�H=��G=LG= LF=�E=O�D=� D=�;C=�uB=��A=��@=�@=�S?=��>=׼==��<= !<=)Q;=�:=N�9=7�8=�8=7,7=3S6=tx5=ߛ4=X�3=��2==�1=�1=u.0=!E/=XY.=
k-=z,=j�+=�*=��)=�(=��'=��&=��%=�$={#=Gj"=�U!=�= =Q!==��=)�=I�=V=o =S�=��=Sd=a=��=a~=G(=x�=�m=�	=��	=�2=��=�I=*�=8N=�� =h��<�h�<{F�<B�<0��<U��<o�<�&�<��<ۀ�<$�<��<X�<:��<u�<r��<�|�<���<r�<��<�U�<;·<�*�<g��<��<YR�<G��<�	�<Gb�<���<��<�`�<���<m�<[S�<���<K�<�z<_s<v�k<Wd<��\<�U<8N<��F<x�?<�-8<
�0<�)<3B"<��<M�<\�<�L<`<�;}��;F��;�|�;�\�;�M�;	R�;�h�;n��;��{;X`;�3E;!@*;`~;���:�1�:;��:�D:�SN9&�H���7�z�u���a�ߺ+��^��(h7���N���e���|��}��㒔�ɂ���L��5�p����ɻ*�ӻ�	޻�����V��\i�q�S���9���A��s�D�!�c�%��*��;.�dI2�MI6�<:�">�~�A��E��I��AM���P���T�y'X���[��:_��b��*f���i���l�\Wp���s���v�2Dz�z�}�ja����������	,�������Q��<ቼ�n��]���9���G��ؒ�����|�������������k���B��,���O������J
��M��������v��~識�g���ߪ��W��6ϭ��F��G����5��V���%������������h�����e����  �  �N=q�M=�M=�NL=�K=��J=|J=�QI=�H=��G=HG=�KF=�E=S�D=� D=�;C=�uB=��A=��@=�@=�S?=�>=߼==��<=!<=+Q;=�:=O�9=1�8=�8=7,7=@S6=wx5=�4=\�3=��2=C�1=}1=.0=#E/=WY.=k-=z,=n�+=�*=��)=�(=��'=Ɨ&=��%=�$={#=Dj"=�U!=�= =N!==��=!�=H�=V=w =S�=��=Wd=]=��=a~=K(=s�=�m=�	=��	=�2=��=�I=*�=<N=�� =l��<�h�<|F�<D�<"��<R��<o�<�&�<��<΀�<$�<��<X�<F��<�t�<n��<�|�<���<�q�<��<�U�<.·<�*�<c��<��<RR�<U��<�	�<Fb�<˸�<}�<�`�<���<l�<ZS�<���<Z�<�z<us<l�k<2Wd<��\<"�U<C8N<|�F<t�?<�-8<�0<{�)<HB"<��<3�<y�<�L<�<�;x��;"��;}|�;�\�;�M�;�Q�;�h�;M��;ũ{;�W`;�3E;7@*;&~;���:�0�:`��:E:|TN9��H����!�z����Έߺ��F���g7�кN�[�e�ք|�9}��ђ��т��M��h��o����ɻ��ӻ
޻���۶�V��:i�}�`��	:�ܲ�M��s�2�!���%��*��;.�CI2�NI6�<:��!>���A���E��I��AM���P���T�|'X���[��:_��b��*f���i���l�NWp���s���v�1Dz�x�}�ya����������,�������Q��-ቼ�n��Y���.���N��ܒ�����m�������������x���L��0���@������=
��U��������v���識�g���ߪ��W��7ϭ��F��8����5��K���%��霶�������V�����g����  �  �N=y�M=�M=|NL=�K=��J=yJ=wQI=�H=��G=NG=�KF=�E=S�D=� D=�;C=�uB=��A=��@=�@=�S?=�>=ݼ==��<=!<=&Q;=�:=W�9=0�8=�8=6,7==S6=yx5=�4=a�3=��2=H�1=|1=�.0= E/=_Y.=k-=z,=v�+=�*=��)=�(=��'=��&=��%=�$=�z#=Oj"=�U!=�= =J!=	=��=�=R�=V=r =K�=��=Ud=]=��=]~=S(=x�=�m=�	=��	=�2=��=�I=1�=AN=�� =o��<�h�<zF�<\�<)��<c��<o�<�&�<"��<̀�<$�<���<X�<<��<�t�<|��<�|�<���<�q�<��<�U�<2·<�*�<U��<��<AR�<L��<�	�<Ob�<¸�<{�<�`�<���<��<cS�<���<c�<�z<�s<��k<EWd<��\<0�U<68N<��F<��?<�-8<5�0<�)<4B"<��<&�<o�<jL<[<�;J��;R��;�|�;h\�;�M�;ZQ�;�h�;%��;'�{;�W`;}3E;�?*;�};|��:-0�:���:�C:XN9��H����U�z�����8�ߺ���H���g7�s�N��e��|�}��쒔������L��Z񴻤o����ɻ��ӻ
޻�����W��Qi���4��:���^��s�5�!���%��*��;.�XI2�qI6�-<:��!>���A���E��I��AM���P���T�U'X���[��:_��b��*f���i���l�OWp��s���v�8Dz�K�}�sa����������,����Q��1ቼ�n��h���9���R��Β�����n�������������t���:��=���K������F
��\��������v���識�g���ߪ��W��/ϭ��F��/����5��A��� %������������]�����N����  �  �N=n�M=�M=|NL=��K=��J=wJ=�QI=�H=��G=DG=�KF=��E=R�D=� D=�;C=�uB=��A=��@=�@=�S?=��>=׼==��<=!<=(Q;=�:=L�9=2�8=�8=:,7=<S6=�x5=�4=\�3=��2=D�1=�1=�.0=$E/=YY.=k-=z,=l�+=�*=��)=�(=��'=&=��%=�$=�z#=Dj"=�U!=�= =L!==��=�=G�=V=v =T�=��=Sd=b=��=c~=J(=t�=�m=�	=��	=�2=��=�I=/�==N=�� =���<�h�<�F�<J�<)��<P��<o�<�&�<��<ր�<$�<��<X�<A��<�t�<j��<�|�<���<�q�<��<�U�<(·<�*�<W��<��<YR�<L��<�	�<Qb�<���<��<�`�<���<s�<bS�<���<g�<�z<ws<y�k<3Wd<�\<@�U<;8N<��F<��?<�-8<�0<��)<3B"<��<1�<g�<�L<|<�;T��;��;j|�;R\�;�M�;�Q�;�h�;��;��{;IW`;�3E;+@*;Z~;���:�0�:���:@D:�TN9R�H������z����l�ߺo����h7���N�S�e�<�|�#}��В��Ƃ���L��d��o����ɻ�ӻ�	޻������V��Bi���d��:���W��s�E�!���%��*��;.�LI2�LI6�<:�">�}�A�
�E���I��AM���P���T�u'X���[��:_��b��*f���i���l�DWp�̬s���v�$Dz�p�}�ta����������,�������Q��9ቼ�n��[���4���\���������r�����������~���P��<���D������F
��Z��������v��z識�g���ߪ��W��/ϭ��F��+����5��K���%��Ꜷ���|���[�����a����  �  .�N=
�M=�M=�HL=��K=��J=�	J=*II=�H=0�G=�G=�@F=}E=��D=I�C=9-C=TfB=��A=��@=�@=$A?=Bu>=%�==��<=L
<=l9;=/g:=s�9=B�8=e�7=�7=�46=�X5={4=O�3=��2=��1=��0=E0=�/={/.=�?-=�M,=X+=�`*=�e)=$h(==g'='c&=�[%=�P$=�B#=�0"=!=� =F�=�=��=5t=�F=�==�=��=Vd=� =V�=p�=�9=��=&�=�)=��
=)]	=��=@~= =`�=P=� =��< ��<|��<ŧ�<~x�<~A�<8�<���<nq�<��<��<�e�<���<���<�#�<��<%3�<���<r/�<!��<��<Ċ�<6��<^`�<^Ƭ<�)�<>��<y�<�D�<���<��<�M�<]��<���<<K�<��<P��<��z<�(s<��k<wqd<I]<��U<�gN<G<��?<Qr8<�&1<h�)<�"<�]<j$<��<�<a7�;���;���;V��;���;ꏶ;���;�ƚ;8 �;�~;fc;�\H;ނ-;��;���:aN�:<�:�8):ȅ9�
�5��Tjj��l���"׺����{�5	3��OJ�yPa��x��;��EN��\<��{��n����(��łǻf�ѻ��ۻp�廮}�x"��R�B���
��,�˩�{�9s�t� ���$��-)��N-��a1�g5�:_9��J=��)A��D�}�H��L��2P���S�QwW��
[���^�1b���e�_i��jl���o�'s��zv��y�S}�(���Ł��`��t�������9#��ڴ��JD���ь��]���珼�o�������{�������������c�������������o|�������s���;i��㧼�\���ժ�O���ǭ��@��f���2��쪳��#������Y�����
�����������  �  (�N=�M=�M=�HL=��K=��J=�	J=#II=�H=,�G=�G=�@F=}E=��D=Q�C=@-C=TfB=��A=��@=�@='A?=:u>=&�==��<=V
<=p9;=-g:=r�9=<�8=n�7=�7=�46=�X5={4=H�3=��2=��1=��0=E0=�/=z/.=�?-=�M,=�X+=�`*=�e)=$h(=>g'=$c&=�[%=�P$=�B#=�0"=!=� =M�=�=��=7t=�F=�=D�=��=Qd=� =U�=y�=�9=��=!�=�)=��
=']	=��=<~==R�=G=� =��<��<z��<ԧ�<qx�<yA�<5�<ʽ�<�q�<{�<��<te�<���<���<�#�<��<&3�<���<�/�<0��<��<Ɋ�<8��<S`�<jƬ<�)�<<��<y�<�D�<���<��<�M�<Q��<���<9K�<���<Q��<��z<�(s<��k<kqd<L]<��U<�gN<G<�?<6r8<�&1<`�)<$�"<�]<d$<��<��<�7�;���;���;n��;���;#��;��;ǚ;6 �;B�~;�ec;�\H;�-;��;���:�M�:a=�:�9):Vǅ9x
����!hj��l���"׺����{��	3��PJ�lPa�x��;��TN��`<����������(����ǻ$�ѻ��ۻd���}�x"���Q�Y��
��,�Ʃ�]�s�h� ���$��-)��N-��a1�g5�N_9��J=��)A���D�w�H��L��2P���S�HwW�[���^�Cb�y�e��i��jl�}�o�'s��zv��y�4}�'(���Ł��`��k���s���B#��ٴ��ZD���ь��]���珼�o�������{������{������^������$�������w|�������s���-i��㧼�\���ժ�	O���ǭ��@��e���2��𪳼�#�� ���W�����"
�����������  �  &�N=�M=�M=�HL=��K=��J=�	J="II=��H=*�G=�G=�@F=�|E=��D=I�C=>-C=RfB=��A=��@=�@=+A?=:u>=/�==��<=U
<=k9;=+g:=z�9=9�8=p�7=�7=�46=�X5={4=P�3=��2=��1=��0=H0=�/=x/.=�?-=�M,=�X+=�`*=�e)=!h(=Ag'=(c&=�[%=�P$=�B#=�0"=!=� =I�=�=��=7t=�F=�=E�=��=Sd=� =Q�=z�=�9=��="�=�)=��
=#]	=��=7~==V�=M=� =��<"��<p��<ק�<nx�<�A�<5�<���<�q�<r�<��<we�<���<���<�#�<��<$3�<���<r/�<(��<��<͊�<9��<M`�<sƬ<�)�<I��<x�<�D�<���<���<�M�<L��<���<.K�< ��<P��<��z<�(s<��k<�qd<6]<��U<�gN<�G<"�?</r8<�&1<J�)<�"<�]<\$<��<��<�7�;���;���;���;m��;��;š�;�ƚ;( �;K�~;�ec;�\H;Z�-;��;���:cM�:Q=�:�8):Rƅ9�
�S���gj�{m��F"׺���{�	3��PJ��Oa�Xx�z;��ZN��q<��m�������(���ǻ,�ѻ�ۻP�廪}ﻄ"���Q�i�z�
��,�Ω�l�3s�n� ���$��-)��N-��a1�g5�E_9��J=��)A���D���H�݀L��2P���S�KwW�[���^�Vb�e�e��i��jl�{�o�('s��zv�2�y�-}�*(���Ł��`��u���t���J#��Ǵ��XD���ь��]���珼�o�������{������������Z������*�������z|��|����s���3i��#㧼�\�� ֪�O���ǭ��@��f���)2��᪳��#���c�����
�����������  �  '�N=�M=�M=�HL=��K=��J=�	J=(II=��H=.�G=�G=�@F=}E=��D=P�C=A-C=ZfB=��A=��@=�@=*A?=?u>=(�==��<=P
<=n9;=-g:=t�9=:�8=h�7=�7=�46=�X5={4=I�3=��2=��1=��0=G0=�/=v/.=�?-=�M,=�X+=�`*=�e)=#h(=:g'=)c&=�[%=�P$=�B#=�0"=!=� =O�=�=��=;t=�F=�=@�=��=Vd=� =T�=v�=�9=��= �=�)=��
=$]	=��=7~=�=T�=H=� =��<"��<n��<ǧ�<mx�<{A�<4�<Ž�<tq�<y�<��<~e�<���<���<�#�<	��<23�<���</�<0��<��<ϊ�<5��<[`�<iƬ<�)�<E��<p�<�D�<���<���<�M�<N��<���<,K�<��<P��<��z<(s<��k<gqd<!]<��U<�gN<�G<�?<3r8<�&1<S�)<#�"<�]<V$<��<�<�7�;���;���;���;���;&��;���;ǚ;j �;8�~;fc;�\H;O�-;W�;��:�M�:�<�:�9):qǅ9�
���jij�vm��"׺Ȩ�Z|�	3��PJ��Pa�:x�{;��RN���<����������(��ڂǻ2�ѻ��ۻ��廝}�i"���Q�H���
��,����W�s�Y� �t�$��-)��N-��a1�g5�8_9��J=��)A���D���H��L��2P���S�]wW�[���^�Rb���e��i��jl���o�%'s��zv�3�y�L}�*(���Ł��`��o�������B#��մ��OD���ь��]���珼�o�������{������{������X�������������q|������s���/i�� 㧼�\���ժ�O���ǭ��@��e���-2�������#�����m�����
�����������  �  (�N=�M=�M=�HL=��K=��J=�	J=)II=�H=4�G=�G=�@F=	}E=��D=T�C=>-C=]fB=��A=��@=�@='A?=>u>=%�==��<=P
<=q9;=-g:=m�9==�8=l�7=�7=�46=�X5={4=G�3=��2=��1=��0=?0=�/=w/.=�?-=�M,=|X+=�`*=�e)=(h(=?g'=%c&=�[%=�P$=�B#=�0"=!=� =K�=�=��=@t=�F=�=@�=��=Sd=� =Z�=t�= :=��=�=�)=��
=#]	=��=;~=�=T�=F=� =��<��<t��<̧�<qx�<mA�</�<ͽ�<sq�<��<��<{e�<���<���<$�<��<73�<���<�/�<'��<��<֊�<=��<e`�<bƬ<�)�<>��<~�<�D�<���<��<�M�<P��<���<2K�<���<G��<��z<t(s<��k<Wqd<F]<y�U<�gN<G<�?<8r8<�&1<[�)<"�"<�]<w$<��<�<r7�;��;��;���;ǐ�;��;%��;�ƚ;� �;[�~;�fc;�\H;(�-;U�;���:�N�:�<�:o:):zǅ9'
�2��ohj��l��V#׺����{��	3��PJ��Pa��x��;��dN��y<��|�������(����ǻ:�ѻ��ۻ_�廹}�V"���Q�.���
��,����e�"s�d� �`�$��-)��N-��a1�
g5�D_9��J=��)A���D�j�H���L��2P���S�VwW�[���^�Cb���e��i��jl���o�#'s�	{v�%�y�?}�%(���Ł��`��f�������3#��ش��QD���ь��]��x珼�o�������{�������������R�������������m|�������s���/i��㧼�\���ժ�
O���ǭ��@��o���2�������#��	���Z�����)
�����������  �  #�N=�M=�M=�HL=��K=��J=�	J=(II=��H=3�G=�G=�@F=
}E=��D=T�C=D-C=\fB=��A=��@= @=.A?==u>=.�==��<=Q
<=l9;=+g:=v�9=7�8=i�7=�7=�46=�X5=	{4=B�3=|�2=��1=��0=A0=�/=s/.=�?-=�M,=�X+=�`*=�e)= h(=Fg'=%c&=�[%=�P$=�B#=�0"=
!=� =P�=
�=��=?t=�F=�=J�=��=Rd=� =P�=u�=�9=��=�=�)=��
=]	=��=2~=�=L�=?=� =��<��<i��<ǧ�<fx�<zA�</�<���<uq�<v�<��<ye�<���<���<�#�<��<43�<���<�/�<4��<��<Պ�<B��<_`�<zƬ<�)�<E��<��<�D�<���<���<�M�<I��<���<'K�<���<C��<��z<w(s<��k<Uqd<-]<m�U<�gN<�G<	�?<!r8<�&1<P�)<�"<�]<n$<��<
�<�7�;��;
��;���;ѐ�;?��;%��;1ǚ;� �;w�~;Ufc;<]H;��-;O�;���:N�: =�:a9):ǅ9!
�����hj��m���"׺ ���{��	3�QJ��Pa�lx��;��yN���<����������(��̂ǻ:�ѻ�ۻ �建}�T"���Q�@�t�
��,����N�s�J� �d�$��-)��N-��a1�g5�F_9��J=��)A���D�}�H��L��2P���S�`wW�[���^�cb���e��i��jl���o�9's��zv�9�y�G}�/(���Ł��`��r���}���D#��ƴ��SD���ь��]���珼�o�������{������w������R�������������o|�������s���3i�� 㧼�\��֪�O���ǭ��@��r���-2�������#��	���f�����(
�����������  �  �N=�M=�M=�HL=��K=��J=�	J=#II=��H=0�G=�G=�@F=
}E=��D=R�C=K-C=ZfB=��A=��@=�@=/A?=9u>=0�==��<=X
<=m9;=)g:=r�9=/�8=l�7=�7=�46=�X5={4=C�3=x�2=��1=��0=C0=�/=v/.=�?-=|M,=�X+=�`*=�e)=h(=Dg'='c&=�[%=�P$=�B#=�0"=!=� =Q�=
�=��=;t=�F=�=J�=��=Rd=� =M�=|�=�9=��=�=�)=��
=]	=��=+~=�=H�=>=� =��<��<W��<˧�<Vx�<qA�<.�<���<�q�<n�<��<qe�<���<���<�#�<��<03�<���<�/�<>��<��<׊�<K��<Z`�<|Ƭ<�)�<K��<z�<�D�<���<���<�M�<:��<���<#K�<�<A��<��z<u(s<v�k<Uqd<]<b�U<�gN<�G<�?<r8<�&1<9�)<3�"<�]<_$<��<��<�7�;���;-��;���;ِ�;n��;��;gǚ;y �;�~;�fc;%]H;��-;�;/��:�M�:�=�:�9):9ƅ9
�_���gj�rn���"׺J��!|��	3�GQJ��Pa��x��;���N��}<�����٩���(���ǻ�ѻ�ۻ-�廧}�m"���Q�F�[�
��,����I�s�7� �q�$��-)��N-��a1�g5�E_9��J=��)A���D���H��L��2P�	�S�TwW�9[���^�}b���e��i��jl���o�O's��zv�Z�y�<}�=(���Ł��`��x���n���J#��ƴ��ZD���ь��]���珼�o�������{������n������P�������������z|��z����s���#i��.㧼�\��֪�O���ǭ��@��u���52�������#��	���o�����(
�����������  �  !�N=�M=�M=�HL=��K=��J=�	J=)II=��H=5�G=�G=�@F=}E=��D=W�C=L-C=_fB=��A=��@=�@=0A?=Au>=/�==��<=O
<=l9;=-g:=p�9=5�8=l�7=�7=�46=�X5={4=?�3=z�2=��1=��0=<0=�/=v/.=�?-=M,=�X+=�`*=�e)="h(=Cg'=+c&=�[%=�P$=�B#=�0"=!=� =Q�=�=��=At=�F=�=G�=��=Wd=� =T�=t�=�9=��=�=�)=��
=]	=��=-~=�=H�=;=�� =��<��<Y��<ʧ�<]x�<jA�<2�<���<pq�<�<��<e�<���<���<$�<��<;3�<���<�/�<<��<��<���<H��<h`�<uƬ<�)�<P��<��<�D�<���<���<�M�<B��<���<'K�<을<4��<��z<\(s<�k<=qd<]<N�U<gN<�G<�?<r8<�&1<H�)<�"<�]<t$<��<�<�7�;��;*��;΢�; ��;p��;F��;pǚ;� �;��~;�fc;:]H;у-;��;��:�N�:�<�:�9):�ȅ9R
�����gj�n��^#׺E��E|�
3�"QJ��Pa��x��;���N��w<����������(����ǻ+�ѻ��ۻ2�廄}�;"���Q�%�^�
��,����G�s�/� �W�$��-)��N-��a1��f5�0_9��J=��)A���D���H��L��2P��S�VwW�8[���^�pb���e��i��jl���o�I's�{v�R�y�=}�5(���Ł��`��v�������9#��Ǵ��KD���ь��]��w珼�o�������{������o������G�������������k|��u����s���1i��&㧼�\��	֪�O���ǭ��@������22������#�����n��'���/
�����������  �  "�N=�M=�M=�HL=��K=��J=�	J=/II=��H=;�G=�G=�@F=}E=��D=\�C=J-C=gfB=��A=��@=@=2A?=Du>='�==��<=Q
<=r9;=)g:=m�9=6�8=`�7=�7=�46=�X5= {4=8�3=y�2=��1=��0=90=�/=n/.=�?-=M,=yX+=�`*=�e)=(h(=Bg'=%c&=�[%=�P$=�B#=�0"=!=� =Y�=�=��=It=�F=�=I�=��=Rd=� =Y�=r�=�9=��=�=�)=��
=]	=��=.~=�=D�=5=ۊ =��<���<a��<���<]x�<hA�<#�<Ƚ�<pq�<��<��<�e�<���<���<
$�<��<K3�<���<�/�<B��<��<銷<F��<t`�<zƬ<�)�<>��<��<�D�<���<��<�M�<E��<���<!K�<�<2��<��z<@(s<��k<"qd<]<M�U<�gN<�G<��?<r8<�&1<U�)<!�"<�]<{$<��<)�<�7�;L��;%��;��;(��;|��;p��;iǚ;� �;�~;�fc;�]H;�-;��;(��:;O�:3=�:;):�ƅ9�
�l���jj��m���#׺1��h|�n
3�8QJ�QQa�}x��;��vN���<����������(����ǻ8�ѻ��ۻ=�廴}�"���Q��l�
��,����(��r�,� �8�$��-)��N-��a1��f5�A_9��J=��)A���D�m�H��L��2P��S�{wW� [�ϕ^�kb���e��i�kl���o�D's�{v�B�y�k}�4(���Ł��`��g������1#��մ��ID���ь��]��s珼�o��u����{������h������>�������������^|�������s���0i��㧼�\��֪� O���ǭ��@������32������#��"���p��(���.
�����������  �  #�N=�M=�M=�HL=��K=��J=�	J=-II=��H=7�G=�G=�@F=
}E=��D=]�C=L-C=afB=��A=��@=@=/A?=Cu>=-�==��<=Q
<=n9;="g:=q�9=4�8=b�7=�7=�46=�X5={4==�3=w�2=��1=��0=60=�/=k/.=�?-=�M,={X+=�`*=�e)=#h(=Eg'=+c&=�[%=�P$=�B#=�0"=!=� =Y�=�=��=Et=�F=�=F�=��=Ud=� =R�=s�=�9=��=�=�)=��
=]	=��=)~=�=D�=9=݊ =��<���<T��<���<Xx�<oA�<�<���<qq�<{�<��<�e�<���<���<$�<(��<@3�<���<�/�<H��<��<銷<Z��<k`�<sƬ<�)�<L��<��<�D�<���<���<�M�<E��<���<K�<䝄</��<z�z<M(s<o�k<1qd<]<H�U<igN<�G<��?<r8<�&1<4�)<�"<�]<w$<��<"�<�7�;,��;r��;���;ܐ�;���;|��;|ǚ;� �;l�~;1gc;o]H;׃-;��;��:�N�:C=�:K:):�Å9%
����jj�&n��$׺h��M|�
3�QQJ�%Qa��x��;���N���<����������(���ǻ2�ѻ��ۻ$�廃}�&"���Q��D�
��,����&��r�:� �F�$��-)��N-��a1��f5�1_9��J=��)A���D���H�	�L��2P��S��wW�=[�ە^�}b���e��i��jl���o�W's�({v�X�y�e}�9(���Ł�a��p���}���<#��ɴ��HD���ь��]��l珼�o�������{������c������?�������������d|��y����s���2i��,㧼�\��֪�O��ȭ��@������82������#�����s��*���:
�����������  �  �N=�M=�M=�HL=��K=��J=�	J=,II=�H=7�G=�G=�@F=}E=��D=\�C=W-C=afB=��A=��@=@=4A?=Bu>=2�==��<=P
<=o9;='g:=r�9=0�8=i�7=�7=�46=�X5=�z4=9�3=p�2=��1=��0=90=�/=o/.=�?-=}M,=�X+=�`*=�e)= h(=Fg'=/c&=�[%=�P$=�B#=�0"=!=� =\�=�=ĝ=Dt=�F=�=L�=��=Xd=� =O�=w�=�9=��=�=�)=��
=]	=��=$~=�==�=3=Պ =y�<���<D��<���<Px�<lA�<#�<���<pq�<v�< ��<�e�<  �<���<$�<(��<>3�<���<�/�<W��<��<抷<W��<l`�<�Ƭ<�)�<W��<��<�D�<���<���<�M�<:��<���<K�<ܝ�<1��<Y�z<B(s<Q�k<$qd<�]<J�U<cgN<�G<��?<r8<�&1<4�)<'�"<�]<n$<��<�<�7�;/��;\��;���;��;搶;s��;�ǚ;� �;t�~;gc;�]H;.�-;��;���:�N�:4=�:�:):Zƅ9�
����vhj��n���#׺����|�`
3��QJ�[Qa�	x��;���N���<�����ȩ���(���ǻ�ѻ��ۻ��_}�!"���Q��F�
��,�t����r�� �H�$��-)��N-��a1��f5�%_9��J=��)A���D���H���L��2P��S�owW�_[�˕^��b���e��i�
kl���o�d's�{v�x�y�K}�@(���Ł��`��s���}���@#������ID���ь��]��m珼�o�������{������S������B�������������f|��o����s���)i��/㧼�\��֪�O��ȭ��@������H2�����$�� ������)���<
�����������  �  �N=�M=�M=�HL=��K=��J=�	J=.II=��H==�G=�G=�@F=}E=��D=X�C=O-C=gfB=��A=��@=@=1A?=Du>=,�==��<=S
<=q9;='g:=m�9=1�8=d�7=�7=�46=�X5=�z4==�3=w�2=��1=��0=80=�/=n/.=�?-={M,=yX+=�`*=�e)=%h(=Eg'=)c&=�[%=�P$=�B#=�0"=!=� =W�=�=��=It=�F=�=K�=��=Td=� =T�=v�=�9=��=�=�)=��
=]	=��=#~=�=D�=6=׊ =w�<���<J��<���<Rx�<eA�< �<���<tq�<��<��<�e�<���<�<$�<#��<I3�<���<�/�<G��<�<튷<Q��<w`�<~Ƭ<�)�<G��<��<�D�<���<���<�M�<:��<���<K�<❄</��<c�z<K(s<q�k<0qd<�]<@�U<igN<�G<��?<r8<�&1<?�)<.�"<�]<�$<��<%�<�7�;a��;K��;��;?��;���;R��;�ǚ;� �;g�~;gc;�]H;��-;��;���:}O�:�=�:);):Zƅ9�
�����ij��n���#׺����|�
3�AQJ�5Qa� 	x��;���N���<�����֩���(���ǻ�ѻ��ۻ#�廏}�"���Q��Q�
��,�{��-��r� � �5�$��-)��N-��a1��f5�4_9��J=��)A���D���H��L��2P��S�rwW�I[�˕^��b���e��i��jl���o�h's�{v�j�y�Z}�=(���Ł��`��l���z���2#��˴��HD���ь�{]��l珼�o��w����{������d������;������ �������b|��~����s���(i��'㧼�\��֪�O��ȭ��@������D2������#��������.���9
�����������  �  $�N=	�M=�M=�HL=��K=��J=�	J=4II=��H=>�G=�G=�@F=}E=��D=k�C=P-C=ifB=��A=��@=	@=-A?=Ju>=(�==��<=K
<=l9;='g:=n�9=3�8=^�7=�7=�46=�X5=�z4=6�3=p�2=��1=��0=50=�/=j/.=�?-=�M,=yX+=�`*=�e)=!h(=Eg'=,c&=�[%=�P$=�B#=�0"=!=� =a�=�=��=Lt=�F=�=H�=��=Yd=� =R�=m�=�9=��=�=�)=��
=]	=��="~=�==�=/=׊ =s�<���<V��<���<Sx�<iA�<�<���<cq�<��<��<�e�<���<Ĕ�<$�<#��<R3�<���<�/�<R��<��<���<S��<x`�<nƬ<�)�<H��<��<�D�<���<���<�M�<L��<���<K�<杄<)��<f�z<.(s<Q�k<qd<�]<4�U<ngN<�G<��?<$r8<�&1<G�)<�"<�]<�$<��<>�<�7�;f��;S��;��;0��;���;�;�ǚ;� �;c�~;Kgc;�]H;��-;M�;z��:oO�:�<�::):sƅ9�
����	kj��m���#׺����|��
3��QJ��Qa�	x��;���N���<����������(��ǻS�ѻ��ۻ#��z}��!���Q��H�
��,������r�*� �'�$��-)�xN-��a1��f5�#_9��J=��)A��D�}�H��L��2P��S��wW�5[�ڕ^��b�̐e��i�kl���o�n's�%{v�Q�y�x}�<(���Ł��`��q�������4#��Ѵ��;D���ь�y]��h珼�o��n����{������Y������8������ �������U|��~����s���9i�� 㧼�\�� ֪�&O��ȭ��@������B2�����$��)���|��4���7
�����������  �  �N=�M=�M=�HL=��K=��J=�	J=.II=��H==�G=�G=�@F=}E=��D=X�C=O-C=gfB=��A=��@=@=1A?=Du>=,�==��<=S
<=q9;='g:=m�9=1�8=d�7=�7=�46=�X5=�z4==�3=w�2=��1=��0=80=�/=n/.=�?-={M,=yX+=�`*=�e)=%h(=Eg'=)c&=�[%=�P$=�B#=�0"=!=� =W�=�=��=It=�F=�=K�=��=Td=� =T�=v�=�9=��=�=�)=��
=]	=��=#~=�=D�=6=׊ =w�<���<J��<���<Sx�<eA�< �<���<tq�<��<��<�e�<���<�<$�<#��<I3�<���<�/�<G��<�<튷<Q��<w`�<~Ƭ<�)�<G��<��<�D�<���<���<�M�<:��<���<K�<❄</��<c�z<K(s<q�k<0qd<�]<@�U<jgN<�G<��?<r8<�&1<@�)<.�"<�]<�$<��<%�<�7�;b��;L��;��;?��;���;R��;�ǚ;� �;f�~;gc;�]H;��-;��;���:zO�:�=�:#;):Oƅ9�
�����ij��n���#׺����|�
3�CQJ�7Qa�	x��;���N���<�����֩���(���ǻ�ѻ��ۻ#�廏}�"���Q��Q�
��,�{��-��r� � �5�$��-)��N-��a1��f5�4_9��J=��)A���D���H��L��2P��S�rwW�I[�˕^��b���e��i��jl���o�h's�{v�j�y�Z}�=(���Ł��`��l���z���2#��˴��HD���ь�{]��l珼�o��w����{������d������;������ �������b|��~����s���(i��'㧼�\��֪�O��ȭ��@������D2������#��������.���9
�����������  �  �N=�M=�M=�HL=��K=��J=�	J=,II=�H=7�G=�G=�@F=}E=��D=\�C=W-C=afB=��A=��@=@=4A?=Bu>=2�==��<=P
<=o9;='g:=r�9=0�8=i�7=�7=�46=�X5=�z4=9�3=p�2=��1=��0=90=�/=o/.=�?-=}M,=�X+=�`*=�e)= h(=Fg'=/c&=�[%=�P$=�B#=�0"=!=� =\�=�=ĝ=Dt=�F=�=L�=��=Xd=� =O�=w�=�9=��=�=�)=��
=]	=��=$~=�==�=3=Պ =y�<���<D��<���<Px�<mA�<#�<���<qq�<v�< ��<�e�<  �<���<$�<(��<>3�<���<�/�<W��<��<抷<W��<l`�<�Ƭ<�)�<W��<��<�D�<���<���<�M�<:��<���<K�<ܝ�<1��<Y�z<B(s<Q�k<$qd<�]<J�U<cgN<�G<��?<r8<�&1<4�)<'�"<�]<n$<��<�<�7�;0��;]��;���;��;搶;s��;�ǚ;� �;s�~;gc;�]H;,�-;��;���:�N�:/=�:�:):Eƅ9�
�����hj�o���#׺����|�c
3��QJ�]Qa�	x��;���N���<�����ɩ���(���ǻ�ѻ��ۻ��_}�""���Q��F�
��,�t����r�� �H�$��-)��N-��a1��f5�%_9��J=��)A���D���H���L��2P��S�owW�_[�˕^��b�e��i�
kl���o�d's�{v�x�y�K}�@(���Ł��`��s���}���@#������ID���ь��]��m珼�o�������{������S������B�������������f|��o����s���)i��/㧼�\��֪�O��ȭ��@������H2�����$�� ������)���<
�����������  �  #�N=�M=�M=�HL=��K=��J=�	J=-II=��H=7�G=�G=�@F=
}E=��D=]�C=L-C=afB=��A=��@=@=/A?=Cu>=-�==��<=Q
<=n9;="g:=q�9=4�8=b�7=�7=�46=�X5={4==�3=w�2=��1=��0=60=�/=k/.=�?-=�M,={X+=�`*=�e)=#h(=Eg'=+c&=�[%=�P$=�B#=�0"=!=� =Y�=�=��=Et=�F=�=F�=��=Vd=� =R�=s�=�9=��=�=�)=��
=]	=��=)~=�=D�=9=݊ =��<���<U��<���<Xx�<oA�<�<���<qq�<{�<��<�e�<���<���<$�<(��<@3�<���<�/�<H��<��<銷<Z��<k`�<sƬ<�)�<K��<��<�D�<���<���<�M�<E��<���<K�<䝄</��<z�z<M(s<o�k<1qd<]<H�U<igN<�G<��?<r8<�&1<4�)<�"<�]<w$<��<"�<�7�;,��;r��;���;ܐ�;���;{��;|ǚ;� �;k�~;/gc;l]H;Ճ-;��;��:�N�:<=�:<:):tÅ9a
� �� jj�.n��!$׺l��P|�
3�TQJ�(Qa��x��;���N���<����������(���ǻ2�ѻ��ۻ$�廄}�'"���Q��E�
��,����&��r�:� �F�$��-)��N-��a1��f5�1_9��J=��)A���D���H�	�L��2P��S��wW�>[�ە^�}b���e��i��jl���o�W's�({v�X�y�e}�9(���Ł�a��p���}���<#��ɴ��HD���ь��]��l珼�o�������{������c������?�������������d|��y����s���2i��,㧼�\��֪�O��ȭ��@������82������#�����s��*���:
�����������  �  "�N=�M=�M=�HL=��K=��J=�	J=/II=��H=;�G=�G=�@F=}E=��D=\�C=J-C=gfB=��A=��@=@=2A?=Du>='�==��<=Q
<=r9;=)g:=m�9=6�8=`�7=�7=�46=�X5= {4=8�3=y�2=��1=��0=90=�/=n/.=�?-=M,=yX+=�`*=�e)=(h(=Bg'=%c&=�[%=�P$=�B#=�0"=!=� =Y�=�=��=It=�F=�=I�=��=Rd=� =Y�=r�=�9=��=�=�)=��
=]	=��=.~=�=D�=5=ۊ =��<���<a��<���<^x�<hA�<#�<ɽ�<qq�<��<��<�e�<���<���<
$�<��<L3�<���<�/�<B��<��<銷<F��<t`�<zƬ<�)�<>��<��<�D�<���< ��<�M�<E��<���<!K�<�<2��<��z<@(s<��k<"qd<]<M�U<�gN<�G<��?<r8<�&1<V�)<!�"<�]<|$<��<)�<�7�;L��;&��;��;(��;|��;p��;hǚ;� �;�~;�fc;�]H;�-;��;!��:3O�:*=�:;):�ƅ9+
����jj��m���#׺6��l|�r
3�<QJ�UQa��x��;��xN���<����������(����ǻ9�ѻ��ۻ=�廵}�"���Q��l�
��,����(��r�,� �8�$��-)��N-��a1��f5�A_9��J=��)A���D�m�H��L��2P��S�{wW� [�ϕ^�kb���e��i�kl���o�D's�{v�B�y�k}�4(���Ł��`��g������1#��մ��ID���ь��]��s珼�o��u����{������h������>�������������^|�������s���0i��㧼�\��֪� O���ǭ��@������32������#��"���p��(���.
�����������  �  !�N=�M=�M=�HL=��K=��J=�	J=)II=��H=5�G=�G=�@F=}E=��D=W�C=L-C=_fB=��A=��@=�@=0A?=Au>=/�==��<=O
<=l9;=-g:=p�9=5�8=l�7=�7=�46=�X5={4=?�3=z�2=��1=��0=<0=�/=v/.=�?-=M,=�X+=�`*=�e)="h(=Cg'=+c&=�[%=�P$=�B#=�0"=!=� =Q�=�=��=At=�F=�=G�=��=Wd=� =T�=t�=�9=��=�=�)=��
=]	=��=.~=�=H�=<=� =��<��<Z��<ʧ�<^x�<kA�<3�<���<pq�<�<��<�e�<���<���<$�<��<;3�<���<�/�<<��<��<���<H��<g`�<uƬ<�)�<P��<��<�D�<���<���<�M�<B��<���<'K�<을<4��<��z<\(s<�k<=qd<]<N�U<gN<�G<�?<r8<�&1<H�)<�"<�]<u$<��<�<�7�;��;+��;΢�; ��;p��;F��;pǚ;� �;��~;�fc;7]H;΃-;��;��:�N�:�<�:�9):[ȅ9�
����	hj�n��h#׺J��J|�
3�&QJ��Pa��x��;���N��x<����������(����ǻ,�ѻ��ۻ3�廅}�;"���Q�&�_�
��,����G�s�/� �W�$��-)��N-��a1��f5�0_9��J=��)A���D���H��L��2P��S�VwW�8[���^�pb���e��i��jl���o�I's�{v�R�y�=}�5(���Ł��`��v�������9#��Ǵ��KD���ь��]��w珼�o�������{������o������G�������������k|��u����s���1i��&㧼�\��	֪�O���ǭ��@������22������#�����n��'���/
�����������  �  �N=�M=�M=�HL=��K=��J=�	J=#II=��H=0�G=�G=�@F=
}E=��D=R�C=K-C=ZfB=��A=��@=�@=/A?=9u>=0�==��<=X
<=m9;=)g:=r�9=/�8=l�7=�7=�46=�X5={4=C�3=x�2=��1=��0=C0=�/=v/.=�?-=|M,=�X+=�`*=�e)=h(=Dg'='c&=�[%=�P$=�B#=�0"=!=� =Q�=
�=��=;t=�F=�=J�=��=Rd=� =N�=|�=�9=��=�=�)=��
=]	=��=+~=�=H�=?=� =��<��<X��<̧�<Wx�<qA�</�<���<�q�<o�<��<qe�<���<���<�#�< ��<03�<���<�/�<>��<��<׊�<J��<Y`�<{Ƭ<�)�<K��<z�<�D�<���<���<�M�<:��<���<#K�<�<@��<��z<u(s<v�k<Uqd<]<b�U<�gN<�G<�?<	r8<�&1<9�)<4�"<�]<`$<��<��<�7�;���;.��;���;ِ�;n��;��;gǚ;y �;�~;�fc;"]H;��-;�;&��:�M�:�=�:�9):ƅ9s
�u��	hj�}n���"׺O��&|��	3�KQJ��Pa��x��;���N��~<�����ک���(���ǻ�ѻ�ۻ.�廨}�n"���Q�F�[�
��,����I�s�7� �r�$��-)��N-��a1�g5�E_9��J=��)A���D���H��L��2P�	�S�TwW�9[���^�}b���e��i��jl���o�O's��zv�Z�y�<}�=(���Ł��`��x���n���J#��ƴ��ZD���ь��]���珼�o�������{������n������P�������������z|��z����s���#i��.㧼�\��֪�O���ǭ��@��u���52�������#��	���o�����(
�����������  �  #�N=�M=�M=�HL=��K=��J=�	J=(II=��H=3�G=�G=�@F=
}E=��D=T�C=D-C=\fB=��A=��@= @=.A?==u>=.�==��<=Q
<=l9;=+g:=v�9=7�8=i�7=�7=�46=�X5=	{4=B�3=|�2=��1=��0=A0=�/=s/.=�?-=�M,=�X+=�`*=�e)= h(=Fg'=%c&=�[%=�P$=�B#=�0"=
!=� =P�=
�=��=?t=�F=�=J�=��=Rd=� =P�=u�=�9=��=�=�)=��
=]	=��=2~=�=L�=?=� =��<��<i��<ǧ�<fx�<zA�</�<���<vq�<w�<��<ye�<���<���<�#�<��<53�<���<�/�<4��<��<Պ�<B��<_`�<zƬ<�)�<D��<��<�D�<���<���<�M�<H��<���<&K�<���<C��<��z<w(s<��k<Vqd<.]<m�U<�gN<�G<	�?<!r8<�&1<Q�)<�"<�]<o$<��<
�<�7�;��;��;���;ѐ�;?��;%��;0ǚ;� �;u�~;Rfc;9]H;��-;L�;���:N�:�<�:M9):�ƅ9u
�����hj��m��	#׺���{��	3�QJ��Pa�px��;��{N���<����������(��͂ǻ;�ѻ�ۻ �建}�U"���Q�@�t�
��,����N�s�J� �d�$��-)��N-��a1�g5�F_9��J=��)A���D�}�H��L��2P���S�`wW�[���^�cb���e��i��jl���o�9's��zv�9�y�G}�/(���Ł��`��r���}���D#��ƴ��SD���ь��]���珼�o�������{������w������R�������������o|�������s���3i�� 㧼�\��֪�O���ǭ��@��r���-2�������#��	���f�����(
�����������  �  (�N=�M=�M=�HL=��K=��J=�	J=)II=�H=4�G=�G=�@F=	}E=��D=T�C=>-C=]fB=��A=��@=�@='A?=>u>=%�==��<=P
<=q9;=-g:=m�9==�8=l�7=�7=�46=�X5={4=G�3=��2=��1=��0=?0=�/=w/.=�?-=�M,=|X+=�`*=�e)=(h(=?g'=%c&=�[%=�P$=�B#=�0"=!=� =K�=�=��=@t=�F=�=@�=��=Sd=� =Z�=t�= :=��=�=�)=��
=#]	=��=;~=�=T�=F=� =��<��<u��<ͧ�<rx�<mA�<0�<ͽ�<sq�<��<��<|e�<���<���<$�<��<73�<���<�/�<'��<��<֊�<=��<d`�<aƬ<�)�<=��<~�<�D�<���<��<�M�<P��<���<1K�<���<F��<��z<t(s<��k<Wqd<F]<y�U<�gN<G<�?<9r8<�&1<[�)<#�"<�]<x$<��<�<s7�;��;��;���;ǐ�;��;$��;�ƚ;� �;Y�~;�fc;�\H;%�-;R�;���:�N�:�<�:]:):Vǅ9p
�E���hj��l��`#׺����{��	3��PJ��Pa��x��;��eN��z<��~�������(����ǻ;�ѻ��ۻ`�建}�W"���Q�/���
��,����e�"s�d� �`�$��-)��N-��a1�
g5�D_9��J=��)A���D�j�H���L��2P���S�VwW�[���^�Cb���e��i��jl���o�#'s�	{v�%�y�?}�%(���Ł��`��f�������3#��ش��QD���ь��]��x珼�o�������{�������������R�������������m|�������s���/i��㧼�\���ժ�
O���ǭ��@��o���2�������#��	���Z�����)
�����������  �  '�N=�M=�M=�HL=��K=��J=�	J=(II=��H=.�G=�G=�@F=}E=��D=P�C=A-C=ZfB=��A=��@=�@=*A?=?u>=(�==��<=P
<=n9;=-g:=t�9=:�8=h�7=�7=�46=�X5={4=I�3=��2=��1=��0=G0=�/=v/.=�?-=�M,=�X+=�`*=�e)=#h(=:g'=)c&=�[%=�P$=�B#=�0"=!=� =O�=�=��=;t=�F=�=@�=��=Vd=� =T�=v�=�9=��= �=�)=��
=$]	=��=8~=�=T�=H=� =��<#��<o��<ǧ�<nx�<{A�<4�<Ž�<tq�<z�<��<e�<���<���<�#�<	��<23�<���</�<0��<��<ϊ�<4��<Z`�<hƬ<�)�<E��<o�<�D�<���<���<�M�<N��<���<,K�<��<P��<��z<(s<��k<gqd<!]<��U<�gN<�G<�?<4r8<�&1<S�)<$�"<�]<V$<��<�<�7�;���;���;���;���;&��;���;ǚ;i �;7�~;fc;�\H;L�-;T�;��:�M�:�<�:w9):Sǅ9�
���zij�~m��"׺˨�^|��	3��PJ��Pa�=x�|;��SN���<����������(��ۂǻ2�ѻ��ۻ��廝}�j"���Q�H���
��,����W�s�Y� �u�$��-)��N-��a1�g5�8_9��J=��)A���D���H��L��2P���S�]wW�[���^�Rb���e��i��jl���o�%'s��zv�3�y�L}�*(���Ł��`��o�������B#��մ��OD���ь��]���珼�o�������{������{������X�������������q|������s���/i�� 㧼�\���ժ�O���ǭ��@��e���-2�������#�����m�����
�����������  �  &�N=�M=�M=�HL=��K=��J=�	J="II=��H=*�G=�G=�@F=�|E=��D=I�C=>-C=RfB=��A=��@=�@=+A?=:u>=/�==��<=U
<=k9;=+g:=z�9=9�8=p�7=�7=�46=�X5={4=P�3=��2=��1=��0=H0=�/=x/.=�?-=�M,=�X+=�`*=�e)=!h(=Ag'=(c&=�[%=�P$=�B#=�0"=!=� =I�=�=��=7t=�F=�=E�=��=Sd=� =Q�=z�=�9=��=#�=�)=��
=$]	=��=7~==V�=M=� =��<"��<p��<ا�<nx�<�A�<5�<���<�q�<r�<��<we�<���<���<�#�<��<$3�<���<r/�<(��<��<͊�<9��<M`�<sƬ<�)�<H��<x�<�D�<���<���<�M�<L��<���<.K�< ��<P��<��z<�(s<��k<�qd<6]<��U<�gN<�G<#�?</r8<�&1<K�)<�"<�]<\$<��<��<�7�;���;���;���;n��;��;š�;�ƚ;' �;J�~;�ec;�\H;X�-;��;���:_M�:L=�:�8):=ƅ9�
�^���gj��m��L"׺���{� 	3��PJ��Oa�Zx�{;��[N��r<��n�������(����ǻ,�ѻ�ۻQ�廪}ﻄ"���Q�i�z�
��,�Ω�l�3s�n� ���$��-)��N-��a1�g5�E_9��J=��)A���D���H�݀L��2P���S�KwW�[���^�Vb�e�e��i��jl�{�o�('s��zv�2�y�-}�*(���Ł��`��u���t���J#��Ǵ��XD���ь��]���珼�o�������{������������Z������*�������z|��|����s���3i��#㧼�\�� ֪�O���ǭ��@��f���)2��᪳��#���c�����
�����������  �  (�N=�M=�M=�HL=��K=��J=�	J=#II=�H=,�G=�G=�@F=}E=��D=Q�C=@-C=TfB=��A=��@=�@='A?=:u>=&�==��<=V
<=p9;=-g:=r�9=<�8=n�7=�7=�46=�X5={4=H�3=��2=��1=��0=E0=�/=z/.=�?-=�M,=�X+=�`*=�e)=$h(=>g'=$c&=�[%=�P$=�B#=�0"=!=� =M�=�=��=7t=�F=�=D�=��=Qd=� =U�=y�=�9=��=!�=�)=��
=']	=��=<~==S�=G=� =��<��<z��<ԧ�<rx�<yA�<6�<ʽ�<�q�<{�<��<ue�<���<���<�#�<��<&3�<���<�/�<0��<��<Ɋ�<8��<S`�<jƬ<�)�<<��<y�<�D�<���<��<�M�<Q��<���<9K�<���<Q��<��z<�(s<��k<kqd<L]<��U<�gN<G<�?<6r8<�&1<`�)<$�"<�]<d$<��<��<�7�;���;���;n��;���;#��;��;ǚ;6 �;B�~;�ec;�\H;�-;��;���:�M�:^=�:�9):Kǅ9�
����'hj��l���"׺����{��	3��PJ�mPa�x��;��TN��`<����������(����ǻ$�ѻ��ۻd���}�x"���Q�Y��
��,�Ʃ�]�s�h� ���$��-)��N-��a1�g5�N_9��J=��)A���D�w�H��L��2P���S�HwW�[���^�Cb�y�e��i��jl�}�o�'s��zv��y�4}�'(���Ł��`��k���s���B#��ٴ��ZD���ь��]���珼�o�������{������{������^������$�������w|�������s���-i��㧼�\���ժ�	O���ǭ��@��e���2��𪳼�#������W�����"
�����������  �  ��N=��M=�M=eCL=��K=H�J=yJ=6AI=PH=޼G=��F= 6F=�qE=X�D=_�C=�C=�WB=*�A=��@=��?=J/?=�b>=v�==G�<=��;=�";=�O:=�z9=��8=��7=7�6=�6=�:5=�[4=�z3=
�2=�1=��0=$�/=0�.=�.=�-=^#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=i#=S�!=�� =(�=٪=��=hb=8=�	=�=�=�d=%=��=v�=^K=��=��=�H=��=�
=�	=�=�?=]�=wP=>�=�O =d��<�|�<�_�<W:�<��<3��<���<$[�<��<���<�k�<;�<��<�D�<���<�d�<���<Vq�<���<�k�<�<dV�<LƳ<�2�<l��<1�<3g�<�ȡ<e(�<څ�<��<�;�<͔�<��<zC�<���<V�<e�z<�3s<��k<2�d<�6]<��U<q�N<�FG<H�?<1�8<kn1<�-*<#�"<��<��<�Y<3<�$�;���;��;׷�;���;��;Tߩ;]�;�W�;���;�Gf;NWK;u�0;�;�Q�:��:W�:�M7:���9�k������[�m����<Ϻ�M���l�k�.��*F��!]���s����S-��j���᥻<������`ŻX�ϻp�ٻa�㻀f���MK �p���	��/�9��� ����+���$��I(�Ro,�?�0�x�4�ǎ8�o<��c@� <D��H���K�q�O��-S���V��iZ�&�]��a�.�d�th�7�k��Ho��r�� v�rRy���|�p�������.��UɄ�`a������������Q����8���ď��N���֒��]��a㕼�g���꘼~l��G훼m��잼j���硼Od��r़&\��Uק�'R���̪��F�������:��Ŵ���.�������"��������k������Z�������  �  ��N=��M=�M=jCL=��K=A�J=yJ=)AI=NH=ܼG=��F=6F=�qE=[�D=^�C=�C=�WB=4�A=��@=��?=D/?=sb>=y�==>�<=��;=�";=�O:=�z9=��8=��7=9�6=�6=�:5=�[4=�z3=�2=�1=��0=!�/=8�.=�.=�-=b#,=-+=�3*=�7)=�8(=�6'=}1&=�(%=�$=d#=X�!=�� =-�=ݪ=��=lb= 8=�	=��=�=�d=%= �=l�=_K=��=��=I=��=�
=�	=�=�?=`�=rP=;�=�O =R��<�|�<�_�<^:�<��<=��<���</[�<��<���<�k�<%�<٬�<�D�<���<e�<���<\q�<���<�k�<�<tV�<TƳ<�2�<l��<�<.g�<�ȡ<U(�<ㅚ<��<�;�<Д�<��<wC�<���<K�<K�z<�3s<��k<<�d<�6]<��U<��N<�FG<T�?<1�8<~n1<�-*<8�"<p�<ۆ<�Y<�2<�$�;���;!��;��;���;3��;Jߩ;l�;�W�;粀;�Gf;\WK;�0;�; R�:� �:��:O7:��9a�����[�7���U<ϺsN��m�t�.�+F�\!]�N�s����-��N��j᥻������`ŻF�ϻ��ٻZ�㻫f�
��JK ����ߞ	��/�%��� �������$��I(�_o,�:�0���4���8�g<��c@��;D��H�r�K�_�O��-S�~�V�oiZ�)�]��a�"�d�'th�?�k��Ho�7�r�� v�fRy��|�r�������.��JɄ�ca�� ���������a����8���ď��N���֒��]��a㕼�g���꘼nl��?훼m��잼8j���硼Zd���़\��Nק�R���̪��F�������:��д���.�������"��������w������\�������  �  ��N=��M=�M=iCL=��K=D�J=�J=)AI=WH=ܼG=��F=6F=�qE=]�D=^�C=�C=�WB=4�A=��@=��?=L/?=tb>=��==?�<=��;=�";=�O:=�z9=��8=��7=3�6=�6=�:5=�[4=�z3=�2=��1=��0=!�/=6�.=�.=�-=[#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=b#=Y�!=�� =)�=ڪ=��=jb=8=�	=��=�=�d=%=�=k�=aK=��=��=�H=��=�
=�	=�=�?=f�=qP==�=�O =U��<�|�<�_�<X:�<z�<4��<���<'[�<��<���<�k�<,�<��<�D�<���<e�<���<\q�<���<�k�<�<pV�<TƳ<�2�<~��<�<<g�<�ȡ<V(�<ᅚ<��<�;�<Ô�<��<nC�<���<L�<Y�z<4s<��k<T�d<�6]<��U<��N<�FG<P�?<�8<nn1<�-*<5�"<t�<�<Z<�2<%�;���;��;��;m��;I��;Pߩ;{�;�W�;벀;�Gf;�WK;��0;;/S�:� �:<�:aN7:]��9ci����L[�٦��K<Ϻ4N���l�F�.�4+F�� ]�8�s����&-��w���᥻P������#`Ż<�ϻ��ٻ"�㻁f����%K ����ܞ	��/�4��� ����"���$��I(�do,��0���4�Ɏ8�I<��c@��;D��H���K�y�O�.S���V�|iZ�'�]��a��d�)th�7�k��Ho�/�r�� v�xRy���|���������.��QɄ�_a��!����������T����8���ď��N���֒��]��b㕼�g���꘼sl��?훼m���랼5j���硼Pd���़ \��Wק�(R���̪��F�������:��ϴ���.�������"��������u������f�������  �  ��N=��M=�M=fCL=��K=F�J=wJ=-AI=OH=߼G=��F=6F=�qE=_�D=a�C=�C=�WB=2�A=��@=��?=G/?=xb>=s�==E�<=��;=�";=�O:=�z9=��8=��7=7�6=�6=�:5=�[4=�z3=�2=�1=��0=�/=3�.=�.=�-=`#,=-+=�3*=�7)=�8(=�6'=1&=�(%=�$=i#=[�!=�� =+�=ߪ=��=kb=8=�	=�=�=�d=%=��=t�=\K=��=��=I=��=�
=�	=�=�?=X�=rP=9�=�O =\��<�|�<�_�<Z:�<��<;��<���<([�<��<���<�k�</�<��<�D�<���<e�<���<]q�<���<�k�<�<qV�<ZƳ<�2�<l��<"�<.g�<�ȡ<d(�<م�<��<�;�<˔�<��<vC�<���<I�<[�z<�3s<��k<*�d<�6]<��U<g�N<�FG<T�?<*�8<un1<�-*<&�"<��<�<�Y<�2<�$�;���;:��;��;���;Y��;dߩ;}�;�W�;ݲ�;'Hf;eWK;M�0;b;yQ�:��:��:kN7:Z��9fd�����[�b���G=Ϻ�M��m���.��*F��!]��s����=-��^��d᥻+������`Żg�ϻt�ٻh�㻞f����HK �m��Ҟ	��/�-��� �������$��I(�Fo,�3�0���4�ӎ8�v<��c@�<D��H�v�K�c�O��-S���V��iZ�7�]��a�=�d�&th�H�k��Ho� �r�� v�nRy���|�h�������.��OɄ�_a������������Z����8��{ď��N���֒��]��[㕼�g���꘼ql��9훼m��잼-j���硼Sd��r़(\��Mק�!R���̪��F�������:��Ҵ���.�������"��������u������]�������  �  ��N=��M=�M=fCL=��K=F�J=xJ=6AI=NH=�G=��F=6F=�qE=\�D=b�C=�C=�WB=1�A=��@=��?=H/?=�b>=v�==F�<=��;=�";=�O:=�z9=��8=��7=:�6=�6=�:5=�[4=�z3=�2=�1=��0=�/=8�.=�.=�-=\#,=-+= 4*=�7)=�8(=�6'=�1&=�(%=�$=l#=W�!=�� =+�=ߪ=��=jb=!8=�	=�=�=�d=%=��=u�=WK=��=��=�H=��=�
=�	=�=�?=V�=sP=8�=�O =Z��<�|�<�_�<G:�<|�</��<���<,[�<��<���<�k�<=�<��<�D�<���<�d�<���<[q�<���<�k�<�<qV�<SƳ<�2�<n��<2�<0g�<�ȡ<a(�<م�<��<�;�<Ɣ�<��<tC�<���<B�<U�z<�3s<��k<�d<�6]<��U<i�N<�FG<0�?<#�8<[n1<�-*<)�"<{�<��<�Y<3<�$�;���;%��;��;���;@��;nߩ;l�;�W�;Բ�;Hf;�WK;[�0;�;�Q�:��:��:�N7:���9cp��7�﹜ [�󥞺P=ϺN��m���.��*F��!]��s����-��y���᥻F�������_Ży�ϻp�ٻ`��vf���FK �a���	��/�,��� �������$��I(�Do,�2�0�{�4���8�t<��c@�<D��H���K�t�O�.S���V�qiZ�D�]��a�E�d� th�J�k��Ho�"�r�� v�`Ry��|��������.��KɄ�la������������U����8��|ď��N���֒��]��Y㕼�g���꘼ql��A훼m��잼j���硼Sd��v़(\��Jק�/R���̪��F�������:��ٴ���.�������"��������|������\�������  �  ��N=��M=�M=hCL=��K=E�J=}J=.AI=VH=޼G=��F=6F=�qE=b�D=f�C=�C=�WB=9�A=��@=��?=K/?=wb>=}�==@�<=��;=�";=�O:=�z9=��8=��7=2�6=�6=�:5=�[4=�z3=��2=�1=��0=�/=4�.=�.=�-=_#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=d#=^�!=�� =-�=�=��=nb=!8=�	=��=�=�d=%=�=m�=^K=��=��=�H=��=�
=�	=�=�?=\�=kP=5�=�O =A��<�|�<�_�<M:�<��<5��<���<*[�<��<���<�k�<+�<��<�D�<���<e�<���<eq�<���<�k�<�<|V�<YƳ<�2�<}��<!�<6g�<�ȡ<U(�<���<��<�;�<˔�<��<hC�<���<<�<@�z<�3s<��k<2�d<�6]<��U<z�N<�FG<B�?<)�8<in1<�-*<1�"<r�<�<�Y<�2<%�;���;'��;F��;���;u��;�ߩ;��;�W�;��;�Gf;�WK;��0;U;�R�:� �:G�:O7:�9�g��r��s[�٦���<ϺUO��0m���.�W+F�f!]���s����/-�����x᥻)������`ŻD�ϻ��ٻ=�㻌f����-K ����ƞ	��/� ��� �}�����$��I(�do,� �0���4�ю8�Y<��c@��;D��H���K�g�O��-S���V��iZ�:�]��a�+�d�<th�R�k��Ho�Q�r�� v�Ry��|�q�������.��LɄ�ba������������V����8���ď�yN���֒��]��S㕼�g���꘼gl��;훼m���랼.j���硼Qd���़!\��Uק�(R���̪��F������:��޴���.�������"���������������j�������  �  ��N=��M=�M=iCL=��K=C�J=�J=,AI=ZH=ݼG=��F=6F=�qE=g�D=_�C=�C=�WB=?�A=��@=��?=O/?=wb>=��==>�<=��;=�";=�O:=�z9=��8=��7=+�6=�6=�:5=�[4=�z3=��2=�1=��0=%�/=.�.=�.=�-=X#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=d#=g�!=�� =/�=�=��=rb=8=�	=��=�=�d=%=�=k�=cK=��=��=�H=��=�
=�	=�=�?=Z�=iP=5�=�O =>��<�|�<u_�<V:�<s�<5��<���<![�<��<���<�k�<,�<��<�D�<���<e�<���<qq�<���<�k�<�<|V�<nƳ<�2�<���<"�<>g�<�ȡ<Z(�<煚<��<�;�<���<��<`C�<���<H�<)�z<�3s<��k<.�d<�6]<��U<w�N<jFG<P�?<�8<vn1<�-*<3�"<x�<�<Z<�2<2%�;���;s��;U��;���;���;]ߩ;��;�W�;H��;IHf;�WK;֖0;Y;WS�:� �:�:kN7:r��9�a������[������;ϺO��[m���.�w+F�!]���s����]-��~���᥻g������;`Ż�ϻ��ٻ0��rf����K ������	��/���� �|�� ���$�dI(�Yo,��0���4�Ď8�P<��c@��;D��H�x�K�z�O�.S���V��iZ��]��a�2�d�Ath�Q�k��Ho�U�r�� v��Ry���|���������.��TɄ�Ta��!����������N����8��}ď�iN���֒��]��]㕼�g���꘼fl��&훼m���랼-j���硼Rd��}़\��]ק�R���̪��F��	����:��Ӵ���.�������"��������������u�������  �  ��N=��M=�M=gCL=��K=D�J=~J=6AI=UH=�G=��F=6F=�qE=h�D=c�C=�C=�WB=8�A=��@=��?=N/?=�b>=|�==B�<=��;=�";=�O:=�z9=��8=��7=+�6=�6=�:5=�[4=�z3=��2=�1=��0=�/=)�.=�.=�-=W#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=l#=_�!=�� =1�=�=��=sb="8=�	=�=�=�d=%=��=p�=]K=��=��=�H=��=
�
=�	=�=�?=U�=jP=1�=�O =B��<�|�<s_�<N:�<m�<-��<���<[�<��<���<�k�<=�<��<�D�<���<e�<���<tq�<���<�k�<�<wV�<eƳ<�2�<y��<5�<:g�<�ȡ<_(�<ޅ�<��<�;�<���<��<cC�<���<?�<3�z<�3s<��k<�d<�6]<��U<V�N<pFG<@�?<�8<gn1<�-*<)�"<{�<�<�Y<3<%�;���;k��;=��;���;���;�ߩ;��;�W�;��;�Hf;�WK;֖0;�;�R�:p�:��:�M7:a��9�h���﹠[�����+=Ϻ�N��bm���.�7+F��!]���s�����-������᥻j������'`ŻI�ϻ��ٻI��if���0K �`����	��/���� �x������$��I(�>o,� �0�p�4���8�e<��c@��;D��H���K���O�.S���V��iZ�:�]��a�C�d�<th�^�k��Ho�J�r�� v��Ry��|���������.��XɄ�`a������������L����8��rď�zN���֒��]��W㕼�g���꘼kl��/훼	m��잼j���硼Ud��x़#\��Yק�&R���̪��F����� ;��ܴ���.�������"��!�������������r�������  �  ��N=��M=�M=hCL=��K=J�J=zJ=4AI=QH=�G=��F=6F=�qE=d�D=n�C=�C=�WB=:�A=��@=�?=I/?=|b>=y�==H�<=��;=�";=�O:=�z9=��8=��7=2�6=�6=�:5=�[4=�z3=��2=�1=��0=�/=0�.=�.=�-=_#,=-+= 4*=�7)=�8(=�6'=�1&=�(%=�$=s#=[�!=�� =/�=�=��=nb=+8=�	=�=�=�d=%=�=r�=VK=��=��=�H=��=�
=�	=�=�?=P�=hP=-�=�O =<��<�|�<�_�<@:�<{�</��<���<-[�<��<���<�k�<5�<��<�D�<���<e�<���<dq�<���<�k�<�<�V�<[Ƴ<3�<p��</�<1g�<�ȡ<](�<څ�<��<�;�<̔�<~�<dC�<���</�<<�z<�3s<��k<��d<�6]<z�U<Y�N<{FG<$�?<)�8<Rn1<�-*<-�"<u�< �<�Y<3<�$�;��;F��;p��;��;���;�ߩ;��; X�;%��;�Hf;4XK;�0;�;aR�:'�:�:�O7:���98l�����u [�Ǧ���=ϺbO��km�#�.�Y+F�"]���s�7��K-������᥻)������_Żx�ϻ~�ٻ+�㻅f���:K �A��͞	�n/���� �c����u$��I(�#o,�"�0�~�4�Ŏ8�[<��c@�<D��H���K�l�O�	.S���V��iZ�_�]��a�T�d�Dth�k�k�Io�V�r�� v�Ry�!�|�z�������.��GɄ�ja������������W����8��mď�zN���֒��]��B㕼�g���꘼Yl��9훼�l��잼 j���硼Id��z़'\��Nק�4R���̪��F������:��봰��.��ͨ���"��/�������������l�������  �  ��N=��M=�M=jCL=��K=I�J=�J=6AI=[H=�G=��F=6F=�qE=f�D=j�C=�C=�WB==�A=��@=�?=Q/?=�b>=��==F�<=��;=�";=�O:=�z9=��8=��7=.�6=�6=�:5=�[4=�z3=��2=�1=��0=�/=0�.=�.=�-=X#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=p#=]�!=�� =0�=�=��=ob=+8=�	=�=�=�d=!%=�=o�=ZK=��=��=�H=��=�
=�	=�=�?=Q�=fP=-�=�O =:��<�|�<{_�<=:�<n�<'��<���<-[�<��<���<�k�<;�<��< E�<���<e�<���<iq�<���<�k�<�<�V�<[Ƴ<3�<���<6�<>g�<�ȡ<Z(�<䅚<��<�;�<���<�<]C�<���<1�<.�z<�3s<��k<	�d<�6]<z�U<`�N<kFG<$�?<�8<Jn1<�-*<8�"<r�<��<Z<3<7%�;��;F��;���;��;���;�ߩ;��;*X�;D��;^Hf;OXK;�0;�;US�:��:5�:<P7:-��91n��_�﹚ [�2���=ϺdO���m��.�g+F�	"]���s���H-������᥻c������_ŻD�ϻ��ٻ"��Xf�}��K �N��ƞ	�m/���� �f����v$��I(�3o,�
�0�_�4���8�L<��c@�<D��H���K���O�.S���V��iZ�O�]��a�P�d�Ith�k�k�Io�X�r�� v��Ry�$�|���������.��FɄ�ga������������F����8��vď�tN���֒��]��J㕼�g���꘼Sl��8훼 m���랼j���硼Jd��}़\��Qק�9R���̪��F������:��鴰��.��Ǩ���"��(�������������s�������  �  ��N=��M=�M=gCL=��K=D�J=J=1AI=ZH=�G=��F=6F=�qE=p�D=d�C=�C=�WB=?�A=��@=�?=P/?=|b>=|�==A�<=��;=�";=�O:=�z9=��8=��7=)�6=�6=�:5=�[4=�z3=��2=�1=��0=�/=*�.=�.=�-=W#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=o#=c�!=�� =:�=�=��=|b=(8=�	=�=�=�d=%=��=l�=^K=��=��=�H=��=�
=�	=�=�?=O�=aP=(�=�O =4��<�|�<l_�<O:�<h�<.��<���<[�<��<���<�k�<3�<��<�D�<���<e�<���<�q�<���<l�<&�<�V�<lƳ<�2�<���<*�<:g�<�ȡ<^(�<߅�<��<�;�<���<��<`C�<���<4�<�z<�3s<��k<�d<z6]<}�U<R�N<gFG<A�?<��8<wn1<�-*<,�"<}�<�<�Y<3<0%�;���;���;���;���;���;�ߩ;.�;#X�;W��;�Hf;XK;��0;�;�R�:[�:��:;N7:���9b��3��I[�ۧ��l=Ϻ�O���m�5�.��+F�"]���s���x-������᥻f������;`Ż=�ϻ��ٻI�㻂f���!K �T����	�|/���| �b������$�uI(�1o,��0�}�4�Ȏ8�a<��c@��;D��H�q�K�~�O�.S���V��iZ�O�]�%�a�V�d�]th�}�k�Io�d�r�� v��Ry���|���������.��WɄ�]a������������K����8��pď�oN���֒��]��S㕼vg��x꘼Xl��(훼m���랼&j���硼Td��z़"\��[ק�R���̪��F��	���;��洰��.��Ȩ���"��*�������������v�������  �  ��N=��M=�M=fCL=��K=J�J=�J=7AI=ZH=�G=��F=6F=�qE=j�D=i�C=�C=�WB=?�A=��@=�?=Q/?=�b>=��==E�<=��;=�";=�O:=�z9=��8=��7=*�6=�6=�:5=�[4=�z3=��2=�1=��0=�/=+�.=�.=�-=S#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=s#=b�!=�� =4�=�=��=ub=&8=�	=�=�=�d=!%=�=p�=\K=��=��=�H=��=�
=�	=�=�?=P�=cP=*�=�O =:��<�|�<p_�<=:�<b�<$��<���<[�<��<���<�k�<?�<��<E�<���<e�<���<vq�<���<�k�<�<�V�<kƳ<3�<���<4�<Bg�<�ȡ<b(�<ۅ�<��<�;�<���<y�<[C�<���<4�<-�z<�3s<��k<��d<�6]<~�U<T�N<bFG<"�?<��8<Vn1<�-*<'�"<��<��<Z<3<6%�;��;���;~��;۳�;���;�ߩ;��;X�;U��;�Hf;dXK;
�0;-;jS�:��:��:.N7:듢9+o�����k [�����p=Ϻ-O��Xm�5�.��+F�"]���s���l-������᥻�������5`ŻL�ϻ~�ٻ��Uf���K �C����	��/� ��� �d������$�yI(�"o,� �0�j�4���8�D<��c@��;D��H���K���O�+.S���V��iZ�W�]��a�R�d�Tth�u�k��Ho�U�r�� v��Ry�#�|���������.��XɄ�^a������������G����8��mď�nN���֒��]��K㕼}g���꘼\l��)훼�l���랼j���硼Gd��u़%\��]ק�.R���̪��F������:��洰��.��̨���"��0�������������x�������  �  ��N=��M=�M=kCL=��K=E�J=~J=7AI=WH=�G=��F=6F=�qE=i�D=r�C=�C=�WB=C�A=��@=�?=M/?=�b>=|�==B�<=��;=�";=�O:=�z9=��8=��7=.�6=�6=�:5=�[4=�z3=��2=�1=��0=�/=+�.=�.=�-=\#,=-+=4*=�7)=�8(=�6'=�1&=�(%=�$=o#=a�!=�� =5�=�=��=tb=08=�	=�=�=�d=%=�=m�=[K=��=��=�H=��=�
=�	=�=�?=L�=aP=%�=�O =.��<�|�<z_�<;:�<z�<.��<���<,[�<��<���<�k�<9�<��<�D�<���< e�<���<oq�<���<�k�<%�<�V�<bƳ<3�<��<4�<9g�<�ȡ<W(�<ㅚ<��<�;�<͔�<��<[C�<���<!�<)�z<�3s<��k<�d<�6]<^�U<H�N<gFG<.�?<'�8<Pn1<�-*<;�"<m�<�<�Y<3<%�;��;_��;���;���;���;�ߩ;��;KX�;y��;WHf;pXK;Ԗ0;;�R�:��:]�:UP7:��9�g�����~ [�,���>ϺP���m���.��+F�B"]���s�[��o-������᥻;�������_ŻE�ϻ��ٻ,��wf���"K �R����	�]/����x �V�����a$�xI(�:o,��0�o�4���8�U<��c@��;D��H���K�w�O�.S���V��iZ�s�]��a�a�d�[th���k�Io�n�r�� v��Ry�&�|�y�������.��FɄ�ca������������O����8��{ď�hN���֒��]��=㕼}g��y꘼Ml��2훼�l���랼j���硼Pd���़\��Mק�4R���̪��F�����;�������.��Ϩ���"��5�������������u�������  �  ��N=��M=�M=fCL=��K=J�J=�J=7AI=ZH=�G=��F=6F=�qE=j�D=i�C=�C=�WB=?�A=��@=�?=Q/?=�b>=��==E�<=��;=�";=�O:=�z9=��8=��7=*�6=�6=�:5=�[4=�z3=��2=�1=��0=�/=+�.=�.=�-=S#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=s#=b�!=�� =4�=�=��=ub=&8=�	=�=�=�d=!%=�=p�=\K=��=��=�H=��=�
=�	=�=�?=P�=cP=*�=�O =:��<�|�<q_�<=:�<b�<$��<���<[�<��<���<�k�<?�<��<E�<���<e�<���<vq�<���<�k�<�<�V�<kƳ<3�<���<4�<Bg�<�ȡ<b(�<ۅ�<��<�;�<���<y�<[C�<���<4�<,�z<�3s<��k<��d<�6]<~�U<T�N<bFG<"�?<��8<Wn1<�-*<'�"<��<��<Z<3<6%�;��;���;~��;ܳ�;���;�ߩ;��;X�;U��;�Hf;cXK;
�0;,;hS�:��:��:*N7:ⓢ9Mo�� ��o [�����r=Ϻ/O��Ym�6�.��+F�"]���s���l-������᥻�������5`ŻL�ϻ~�ٻ��Uf���K �C����	��/� ��� �d������$�yI(�"o,� �0�j�4���8�D<��c@��;D��H���K���O�+.S���V��iZ�W�]��a�R�d�Tth�u�k��Ho�U�r�� v��Ry�#�|���������.��XɄ�^a������������G����8��mď�nN���֒��]��K㕼}g���꘼\l��)훼�l���랼j���硼Gd��u़%\��]ק�.R���̪��F������:��洰��.��̨���"��0�������������x�������  �  ��N=��M=�M=gCL=��K=D�J=J=1AI=ZH=�G=��F=6F=�qE=p�D=d�C=�C=�WB=?�A=��@=�?=P/?=|b>=|�==A�<=��;=�";=�O:=�z9=��8=��7=)�6=�6=�:5=�[4=�z3=��2=�1=��0=�/=*�.=�.=�-=W#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=o#=c�!=�� =:�=�=��=|b=(8=�	=�=�=�d=%=��=l�=^K=��=��=�H=��=�
=�	=�=�?=O�=aP=(�=�O =4��<�|�<l_�<P:�<h�</��<���<[�<��<���<�k�<3�<��<�D�<���<e�<���<�q�<���<l�<&�<�V�<lƳ<�2�<���<*�<:g�<�ȡ<](�<߅�<��<�;�<���<��<_C�<���<4�<�z<�3s<��k<�d<z6]<}�U<R�N<gFG<A�?<��8<wn1<�-*<,�"<}�<�<�Y<3<1%�;���;���;���;���;���;�ߩ;-�;#X�;V��;�Hf;XK;��0;�;�R�:X�:��:3N7:q��9Gb��D��Q[�ߧ��p=Ϻ�O���m�7�.��+F�"]���s���y-������᥻f������<`Ż=�ϻ��ٻJ�㻂f���!K �T����	�|/���| �b������$�uI(�1o,��0�}�4�Ȏ8�a<��c@��;D��H�q�K�~�O�.S���V��iZ�O�]�%�a�V�d�]th�}�k�Io�d�r�� v��Ry���|���������.��WɄ�]a������������K����8��pď�oN���֒��]��S㕼vg��x꘼Xl��(훼m���랼&j���硼Td��z़"\��[ק�R���̪��F��	���;��洰��.��Ȩ���"��*�������������v�������  �  ��N=��M=�M=jCL=��K=I�J=�J=6AI=[H=�G=��F=6F=�qE=f�D=j�C=�C=�WB==�A=��@=�?=Q/?=�b>=��==F�<=��;=�";=�O:=�z9=��8=��7=.�6=�6=�:5=�[4=�z3=��2=�1=��0=�/=0�.=�.=�-=X#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=p#=]�!=�� =0�=�=��=ob=+8=�	=�=�=�d=!%=�=o�=ZK=��=��=�H=��=�
=�	=�=�?=Q�=fP=-�=�O =:��<�|�<{_�<=:�<n�<'��<���<-[�<��<���<�k�<;�<��< E�<���<e�<���<jq�<���<�k�<�<�V�<[Ƴ<3�<���<6�<>g�<�ȡ<Z(�<䅚<��<�;�<���<�<]C�<���<1�<-�z<�3s<��k<	�d<�6]<{�U<`�N<lFG<$�?<�8<Kn1<�-*<8�"<r�<��<Z<3<7%�;��;F��;���;��;���;�ߩ;��;*X�;D��;\Hf;NXK;�0;�;PS�:��:0�:1P7:��9�n��w�﹥ [�8���=ϺjO���m�
�.�i+F�"]���s���I-������᥻d������_ŻD�ϻ��ٻ"��Xf�}��K �N��ƞ	�m/���� �f����v$��I(�3o,�
�0�_�4���8�L<��c@�<D��H���K���O�.S���V��iZ�O�]��a�P�d�Ith�k�k�Io�X�r�� v��Ry�$�|���������.��FɄ�ga������������F����8��vď�tN���֒��]��J㕼�g���꘼Sl��8훼 m���랼j���硼Jd��}़\��Qק�9R���̪��F������:��鴰��.��Ǩ���"��(�������������s�������  �  ��N=��M=�M=hCL=��K=J�J=zJ=4AI=QH=�G=��F=6F=�qE=d�D=n�C=�C=�WB=:�A=��@=�?=I/?=|b>=y�==H�<=��;=�";=�O:=�z9=��8=��7=2�6=�6=�:5=�[4=�z3=��2=�1=��0=�/=0�.=�.=�-=_#,=-+= 4*=�7)=�8(=�6'=�1&=�(%=�$=s#=[�!=�� =/�=�=��=nb=+8=�	=�=�=�d=%=�=r�=VK=��=��=�H=��=�
=�	=�=�?=P�=hP=-�=�O =<��<�|�<�_�<@:�<|�<0��<���<-[�<��<���<�k�<5�<��<�D�<���<e�<���<dq�<���<�k�<�<�V�<ZƳ<3�<p��</�<1g�<�ȡ<](�<څ�<��<�;�<̔�<~�<dC�<���</�<<�z<�3s<��k<��d<�6]<{�U<Y�N<{FG<$�?<)�8<Sn1<�-*<-�"<u�< �<�Y<3<�$�;��;F��;q��;��;���;�ߩ;��; X�;%��;�Hf;2XK;}�0;�;[R�:!�:�:�O7:k��9�l����﹃ [�Φ���=ϺiO��nm�&�.�\+F�"]���s�8��L-������᥻*������_Żx�ϻ�ٻ,�㻅f���;K �A��͞	�n/���� �c����u$��I(�#o,�"�0�~�4�Ŏ8�[<��c@�<D��H���K�l�O�	.S���V��iZ�_�]��a�T�d�Dth�k�k�Io�V�r�� v�Ry�!�|�z�������.��GɄ�ja������������W����8��mď�zN���֒��]��B㕼�g���꘼Yl��9훼�l��잼 j���硼Id��z़'\��Nק�4R���̪��F������:��봰��.��ͨ���"��/�������������l�������  �  ��N=��M=�M=gCL=��K=D�J=~J=6AI=UH=�G=��F=6F=�qE=h�D=c�C=�C=�WB=8�A=��@=��?=N/?=�b>=|�==B�<=��;=�";=�O:=�z9=��8=��7=+�6=�6=�:5=�[4=�z3=��2=�1=��0=�/=)�.=�.=�-=W#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=l#=_�!=�� =1�=�=��=sb="8=�	=�=�=�d=%=��=p�=]K=��=��=�H=��=
�
=�	=�=�?=U�=jP=1�=�O =C��<�|�<t_�<O:�<n�<.��<���<[�<��<���<�k�<=�<��<�D�<���<e�<���<tq�<���<�k�<�<wV�<eƳ<�2�<y��<5�<9g�<�ȡ<_(�<݅�<��<�;�<���<��<cC�<���<?�<3�z<�3s<��k<�d<�6]<��U<V�N<pFG<@�?<�8<hn1<�-*<*�"<{�<�<�Y<3<%�;���;k��;=��;���;���;�ߩ;��;�W�;��;�Hf;�WK;Ӗ0;�;�R�:i�:��:�M7:A��9Ki��$�ﹰ[�����3=Ϻ�N��fm���.�:+F��!]���s�����-������᥻k������(`ŻJ�ϻ��ٻI��if���0K �`����	��/���� �x������$��I(�>o,� �0�p�4���8�e<��c@��;D��H���K���O�.S���V��iZ�:�]��a�C�d�<th�^�k��Ho�J�r�� v��Ry��|���������.��XɄ�`a������������L����8��rď�zN���֒��]��W㕼�g���꘼kl��/훼	m��잼j���硼Ud��x़#\��Yק�&R���̪��F����� ;��ܴ���.�������"��!�������������r�������  �  ��N=��M=�M=iCL=��K=C�J=�J=,AI=ZH=ݼG=��F=6F=�qE=g�D=_�C=�C=�WB=?�A=��@=��?=O/?=wb>=��==>�<=��;=�";=�O:=�z9=��8=��7=+�6=�6=�:5=�[4=�z3=��2=�1=��0=%�/=.�.=�.=�-=X#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=d#=g�!=�� =/�=�=��=rb=8=�	=��=�=�d=%=�=k�=dK=��=��=�H=��=�
=�	=�=�?=Z�=jP=5�=�O =?��<�|�<u_�<W:�<t�<5��<���<"[�<��<���<�k�<,�<��<�D�<���<e�<���<qq�<���<�k�<�<|V�<mƳ<�2�<���<"�<>g�<�ȡ<Z(�<煚<��<�;�<���<��<`C�<���<G�<)�z<�3s<��k<.�d<�6]<��U<x�N<kFG<P�?<�8<vn1<�-*<3�"<y�<�<Z<�2<3%�;���;t��;V��;���;���;]ߩ;��;�W�;H��;GHf;�WK;Ӗ0;V;PS�:� �:�:[N7:R��9b������[�Ƨ���;ϺO��_m���.�{+F��!]���s����^-�����᥻h������<`Ż�ϻ��ٻ1��rf����K ������	��/���� �|�� ���$�dI(�Yo,��0���4�Ď8�P<��c@��;D��H�y�K�z�O�.S���V��iZ��]��a�2�d�Ath�Q�k��Ho�U�r�� v��Ry���|���������.��TɄ�Ta��!����������N����8��}ď�iN���֒��]��]㕼�g���꘼fl��&훼m���랼-j���硼Rd��}़\��]ק�R���̪��F��	����:��Ӵ���.�������"��������������u�������  �  ��N=��M=�M=hCL=��K=E�J=}J=.AI=VH=޼G=��F=6F=�qE=b�D=f�C=�C=�WB=9�A=��@=��?=K/?=wb>=}�==@�<=��;=�";=�O:=�z9=��8=��7=2�6=�6=�:5=�[4=�z3=��2=�1=��0=�/=4�.=�.=�-=_#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=d#=^�!=�� =-�=�=��=nb=!8=�	=��=�=�d=%=�=m�=^K=��=��=�H=��=�
=�	=�=�?=\�=kP=5�=�O =B��<�|�<�_�<N:�<��<6��<���<+[�<��<���<�k�<,�<��<�D�<���<e�<���<eq�<���<�k�<�<{V�<XƳ<�2�<}��<!�<6g�<�ȡ<U(�<���<��<�;�<˔�<��<gC�<���<<�<@�z<�3s<��k<2�d<�6]<��U<z�N<�FG<B�?<*�8<jn1<�-*<2�"<r�<�<�Y<�2<%�;���;'��;G��;���;u��;�ߩ;��;�W�;��;�Gf;�WK;��0;R;�R�:� �:@�:O7:ԓ�9h����﹃[�ᦞ��<Ϻ]O��4m���.�Z+F�i!]���s����1-�����y᥻*������`ŻE�ϻ��ٻ=�㻌f����-K ����ƞ	��/�!��� �}�����$��I(�do,� �0���4�ю8�Y<��c@��;D��H���K�g�O��-S���V��iZ�:�]��a�+�d�<th�R�k��Ho�Q�r�� v�Ry��|�q�������.��LɄ�ba������������V����8���ď�yN���֒��]��S㕼�g���꘼gl��;훼m���랼.j���硼Qd���़!\��Uק�(R���̪��F������:��޴���.�������"���������������j�������  �  ��N=��M=�M=fCL=��K=F�J=xJ=6AI=NH=�G=��F=6F=�qE=\�D=b�C=�C=�WB=1�A=��@=��?=H/?=�b>=v�==F�<=��;=�";=�O:=�z9=��8=��7=:�6=�6=�:5=�[4=�z3=�2=�1=��0=�/=8�.=�.=�-=\#,=-+= 4*=�7)=�8(=�6'=�1&=�(%=�$=l#=W�!=�� =+�=ߪ=��=jb=!8=�	=�=�=�d=%=��=u�=WK=��=��=�H=��=�
=�	=�=�?=V�=sP=8�=�O =Z��<�|�<�_�<G:�<}�<0��<���<,[�<��<���<�k�<=�<��<�D�<���<�d�<���<[q�<���<�k�<�<qV�<SƳ<�2�<m��<2�<0g�<�ȡ<a(�<م�<��<�;�<Ɣ�<��<tC�<���<B�<U�z<�3s<��k<�d<�6]<��U<i�N<�FG<0�?<#�8<[n1<�-*<)�"<|�<�<�Y<3<�$�;���;%��;��;���;@��;nߩ;l�;�W�;Ӳ�;Hf;�WK;X�0;�;�Q�:��:��:�N7:���9�p��T�﹪ [�����W=Ϻ
N��m���.��*F��!]��s����-��{���᥻G�������_Ży�ϻp�ٻa��vf���FK �b���	��/�,��� �������$��I(�Eo,�2�0�{�4���8�t<��c@�<D��H���K�t�O�.S���V�qiZ�D�]��a�E�d� th�J�k��Ho�"�r�� v�`Ry��|��������.��KɄ�la������������U����8��|ď��N���֒��]��Y㕼�g���꘼ql��A훼m��잼j���硼Sd��v़(\��Jק�/R���̪��F�������:��ٴ���.�������"��������|������\�������  �  ��N=��M=�M=fCL=��K=F�J=wJ=-AI=OH=߼G=��F=6F=�qE=_�D=a�C=�C=�WB=2�A=��@=��?=G/?=xb>=s�==E�<=��;=�";=�O:=�z9=��8=��7=7�6=�6=�:5=�[4=�z3=�2=�1=��0=�/=3�.=�.=�-=`#,=-+=�3*=�7)=�8(=�6'=1&=�(%=�$=i#=[�!=�� =+�=ߪ=��=kb=8=�	=�=�=�d=%=��=t�=\K=��=��=I=��=�
=�	=�=�?=Y�=rP=9�=�O =\��<�|�<�_�<Z:�<��<<��<���<([�<��<���<�k�</�<��<�D�<���<e�<���<^q�<���<�k�<�<qV�<ZƳ<�2�<l��<"�<-g�<�ȡ<d(�<م�<��<�;�<˔�<��<vC�<���<I�<[�z<�3s<��k<*�d<�6]<��U<g�N<�FG<U�?<*�8<vn1<�-*<'�"<��<�<�Y<�2<�$�;���;:��;��;���;Y��;dߩ;|�;�W�;ݲ�;%Hf;dWK;K�0;`;uQ�:|�:��:`N7:D��9�d�����![�g���M=Ϻ�M��m���.��*F��!]��s����>-��_��e᥻,������	`Żg�ϻu�ٻh�㻞f����HK �m��Ҟ	��/�-��� �������$��I(�Fo,�3�0���4�ӎ8�v<��c@�<D��H�v�K�c�O��-S���V��iZ�7�]��a�=�d�&th�H�k��Ho� �r�� v�nRy���|�h�������.��OɄ�_a������������Z����8��{ď��N���֒��]��[㕼�g���꘼ql��9훼m��잼-j���硼Sd��r़(\��Mק�!R���̪��F�������:��Ҵ���.�������"��������u������]�������  �  ��N=��M=�M=iCL=��K=D�J=�J=)AI=WH=ܼG=��F=6F=�qE=]�D=^�C=�C=�WB=4�A=��@=��?=L/?=tb>=��==?�<=��;=�";=�O:=�z9=��8=��7=3�6=�6=�:5=�[4=�z3=�2=��1=��0=!�/=6�.=�.=�-=[#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=b#=Y�!=�� =)�=ڪ=��=jb=8=�	=��=�=�d=%=�=k�=aK=��=��=�H=��=�
=�	=�=�?=f�=qP==�=�O =U��<�|�<�_�<X:�<z�<4��<���<'[�<��<���<�k�<,�<��<�D�<���<e�<���<]q�<���<�k�<�<pV�<TƳ<�2�<}��<�<<g�<�ȡ<V(�<ᅚ<��<�;�<�<��<nC�<���<L�<Y�z<4s<��k<T�d<�6]<��U<��N<�FG<P�?<�8<nn1<�-*<5�"<t�<�<Z<�2<%�;���;��;��;m��;I��;Pߩ;{�;�W�;검;�Gf;�WK;��0;;,S�:� �:8�:ZN7:M��9�i����T[�ަ��O<Ϻ8N���l�H�.�6+F�� ]�:�s����'-��x���᥻P������$`Ż=�ϻ��ٻ"�㻂f����%K ����ܞ	��/�4��� ����#���$��I(�do,��0���4�Ɏ8�I<��c@��;D��H���K�y�O�.S���V�|iZ�'�]��a��d�)th�7�k��Ho�/�r�� v�xRy���|���������.��QɄ�_a��!����������T����8���ď��N���֒��]��b㕼�g���꘼sl��?훼m���랼5j���硼Pd���़ \��Wק�(R���̪��F�������:��ϴ���.�������"��������u������f�������  �  ��N=��M=�M=jCL=��K=A�J=yJ=)AI=OH=ܼG=��F=6F=�qE=[�D=^�C=�C=�WB=4�A=��@=��?=D/?=sb>=y�==>�<=��;=�";=�O:=�z9=��8=��7=9�6=�6=�:5=�[4=�z3=�2=�1=��0=!�/=8�.=�.=�-=b#,=-+=�3*=�7)=�8(=�6'=}1&=�(%=�$=d#=X�!=�� =-�=ݪ=��=lb= 8=�	=��=�=�d=%= �=l�=_K=��=��=I=��=�
=�	=�=�?=`�=rP=;�=�O =R��<�|�<�_�<^:�<��<=��<���</[�<��<���<�k�<%�<٬�<�D�<���<e�<���<\q�<���<�k�<�<tV�<TƳ<�2�<l��<�<.g�<�ȡ<U(�<ㅚ<��<�;�<Д�<��<wC�<���<K�<K�z<�3s<��k<<�d<�6]<��U<��N<�FG<T�?<1�8<~n1<�-*<8�"<q�<ۆ<�Y<�2<�$�;���;!��;��;���;3��;Jߩ;l�;�W�;粀;�Gf;\WK;�0;�;R�:� �:��:
O7:��94a�����[�9���W<ϺvN��m�u�.�+F�\!]�O�s����-��N��j᥻������`ŻF�ϻ��ٻZ�㻫f�
��JK ����ߞ	��/�%��� �������$��I(�_o,�:�0���4���8�g<��c@��;D��H�r�K�_�O��-S�~�V�oiZ�)�]��a�"�d�'th�?�k��Ho�7�r�� v�fRy��|�r�������.��JɄ�ca�� ���������a����8���ď��N���֒��]��a㕼�g���꘼nl��?훼m��잼8j���硼Zd���़\��Nק�R���̪��F�������:��д���.�������"��������w������\�������  �  )}N=�M=H�L=E>L=�}K=�J=��I=�9I=wH=�G=F�F=�+F=�fE=ʠD=!�C=�C=JB=��A=J�@=��?=X?=�P>=́==��<=P�;=�;=L9:=�c9=Y�8=��7=��6=��5=�5=u>4=k\3=\x2=*�1=ǩ0=�/=��.=u�-=W�,=��+=)+=�	*=�)=�(=?	'=�&=�$=��#=n�"=M�!=�� =)�=�t=�Q=�*=��=��=O�=�e=*=��=o�=�\=[=��=�g=�=�=wJ
=��=Jv=�=��=p=��=e =r%�<��<���<���<;��<gw�<{>�<���<��<�j�<��<(��<�^�<���<ŏ�<K �<��<3�<���<4�<r��<%�<=��<�<�t�<�ި<F�<��<��<�n�<�͖<�*�<��<�<!<�<h��<X�<ɍz<�>s<��k<��d<xT]<�V<��N<6wG<+2@<E�8<�1<w*<]A#<<��<��<��<�;���;���;c��;`��;y޸;=
�;-H�;ɚ�;��;��h;6$N;z3;{ ;/q�:�K�:��:��D:Ԛ�9���N�ӹ&�L�\����Ǻ����2��+�gHB�<6Y�T�o�n ���.�����>ࣻ̓������_ûؘͻ>�׻&��q�9��ީ���	�5��B���:����[���:#�Rs'�?�+���/���3���7��;���?�H�C��WG��K�|�N���R�93V��Y�we]���`��sd���g�Mak�Q�n�0r��u��x��2|�~|�,`��G��������5��=͇��b������Ȇ�����E����.��ܸ��dA��Oȕ�N��Ҙ��U���כ�Y��dٞ��X���ס�~U���Ҥ��O��̧�!H���ê�/?��X����5��l���q+�������!��+����������*��㍼�?���  �  0}N=�M=H�L=E>L=�}K=�J=��I=�9I=wH=�G=I�F=�+F=�fE=ɠD=�C=�C=JB=��A=H�@=��?=T?=�P>=Ձ==��<=J�;=�;=Q9:=�c9=_�8=��7=��6=��5={5=o>4=t\3=dx2=0�1=��0=�/=��.=u�-=]�,=��+=/+=�	*=�)=�(=A	'=�&=�$=��#=l�"=T�!=�� =-�=�t=�Q=�*=��=��=L�=�e=�)=��=s�=�\=Y=��=�g=�=�=xJ
=��=Mv=�=��=v=�=` =_%�<�<���<���<J��<�w�<�>�<���<��<�j�<��<��<�^�<���<���<V �<��<3�<���<4�<y��<%�<D��<�<�t�<�ި<&F�<	��<��<�n�<~͖<�*�<��<	�<<�<v��<Q�<��z<�>s<��k<��d<NT]<�V<;N<)wG<72@<d�8<�1<�w*<`A#<�<��<�<f�<t�;���;���;r��;n��;l޸;�	�;*H�;���;��;f�h;$N;�y3; ;Gr�:�J�:@��:x�D:��9lſ�J�ӹ �L��\����Ǻ������~+��GB��5Y���o�` ��p.�����ࣻm���c���_û٘ͻ��׻��q뻓�������	���B����":�ɞ�O���:#�5s'�I�+�¹/���3���7���;��?�N�C��WG��K�G�N�R�43V���Y�ke]��`��sd�z�g�2ak�c�n�+0r��u��x��2|�a|�`��;��������5��H͇��b������҆�����K����.��渒�dA��gȕ�N��yҘ��U���כ�Y��gٞ��X��}ס��U���Ҥ��O�� ̧�H���ê�*?��^���r5��t����+�������!��������Ŕ����ꍼ�:���  �  *}N=�M=E�L=J>L=�}K=�J=��I=�9I=%wH=�G=F�F=�+F=�fE=РD=�C=�C=JB=��A=D�@=��?=\?=�P>=ف==��<=O�;=�;=N9:=�c9=Y�8=~�7=��6=��5=|5=r>4=p\3=Xx2=/�1=��0=�/=��.=q�-=X�,=��+=*+=�	*=�)=�(=C	'=�&=�$=��#=i�"=U�!=�� =1�=�t=�Q=�*=��=��=F�=�e=�)=��=u�=�\=a=��=�g=�=�=tJ
=��=Pv=�=��=k=��=c =a%�<�<���<���<<��<ow�<>�<���<��<�j�<��<��<�^�<���<���<Z �<��< 3�<���<4�<y��<%�<B��<�<�t�<�ި<-F�<
��<��<�n�<|͖<�*�<��<�<<�<y��<T�<��z<�>s<��k<��d<QT]<�V<־N<wG<22@<I�8<�1<sw*<tA#<�<��<)�<k�<��;���;���;]��;i��;�޸;�	�;zH�;���;��;+�h;$N;`z3;4 ;�r�:�J�::?�D:���9���e�ӹy�L��\��W�Ǻ����f���+��HB��5Y���o�J ���.����8ࣻ��������_û��ͻ��׻���p�j�������	���'B����:����5��;#�,s'�_�+���/���3���7��;�$�?�/�C��WG��K�h�N�ۋR�B3V��Y�^e]�
�`��sd���g�Gak�W�n�'0r�،u�!�x��2|�{|�#`��B��������5��K͇��b�����������V����.���PA��bȕ�N��yҘ��U���כ�#Y��Tٞ��X��wס��U���Ҥ��O��"̧� H���ê�/?��c���n5��p����+�������!�� ����������������<���  �  0}N=�M=J�L=B>L=�}K=�J=��I=�9I=wH=�G=J�F=�+F=�fE=͠D=�C=�C=JB=��A=J�@=��?=S?=�P>=ρ==��<=M�;=�;=Q9:=�c9=`�8=��7=��6=��5=|5=r>4=n\3=ax2=,�1=ũ0=�/=��.=w�-=]�,=��+=,+=�	*=�)=�(=@	'=�&=�$=��#=i�"=W�!=�� =.�=�t=�Q=�*=��=��=H�=�e=�)=��=o�=�\=Z=��=�g=�=�=zJ
=��=Fv=�=��=s=��=a =b%�<��<���<���<G��<rw�<�>�<���<��<�j�<��<!��<�^�<���<���<\ �<��<3�<���<4�<u��<"%�<I��<�<�t�<�ި<F�<��<��<}n�<�͖<�*�<��<
�<!<�<e��<K�<��z<�>s<��k<��d<cT]<�V<��N<7wG<92@<d�8<��1<�w*<PA#<�<��<�<p�<~�;���;��;���;d��;�޸;�	�;ZH�;���;��;��h;($N;�y3;I ;�q�:�K�:���:)�D:h��9�뿷�ӹ��L��[����Ǻ����a���+�HB�6Y�t�o�� ���.�����ࣻ����x���_û�ͻk�׻%��q뻄������	���B����:�Þ�D���:#�(s'�W�+���/���3���7��;��?�L�C��WG��K�]�N�ȋR�+3V�
�Y��e]���`��sd���g�Aak�]�n�$0r��u�
�x��2|�d|�`��<��������5��?͇��b������Ն�����L����.��丒�ZA��aȕ�N��|Ҙ��U���כ�"Y��eٞ��X���ס�U���Ҥ��O��̧�H���ê�*?��X����5��z���z+�������!��*������Ɣ��-��㍼�9���  �  2}N=�M=J�L=A>L=�}K=�J=��I=�9I=wH=
�G=F�F=�+F=�fE=ΠD=�C=�C=JB=��A=G�@=��?=S?=�P>=с==��<=H�;=�;=Q9:=�c9=_�8=s�7=��6=��5=�5=m>4=j\3=bx2=$�1=ǩ0=�/=��.=p�-=U�,=��+='+=�	*=�)=�(=?	'=�&=�$=��#=p�"=P�!=�� =0�=�t=�Q=�*=��=��=N�=�e=�)=��=n�=�\=T=��=�g=�=�=qJ
=��=Ev=�=��=r=��=[ =k%�<��<���<���<@��<qw�<>�<���<���<�j�<��<7��<�^�<��<���<R �<��<3�<���<4�<|��<"%�<?��<)�<�t�<�ި<(F�<��<��<yn�<�͖<�*�<��<��<<�<q��<O�<��z<�>s<��k<t�d<YT]<�V<��N<1wG<2@<g�8<�1<�w*<NA#<�<��<�<��<v�;��;���;|��;��;�޸;
�;SH�;ٚ�;��;b�h;�$N;�y3;� ;�q�:�K�:&��:�D:Z��9����E�ӹ!�L��[��y�ǺJ������+�HB��6Y�T�o�� ��m.����Mࣻ��������_û��ͻ[�׻)���p�Y��ة���	�*��B����:����B���:#�Bs'�>�+���/���3���7��;���?�`�C��WG��K�X�N��R�N3V���Y��e]���`�td���g�Kak�r�n�0r��u��x��2|�r|� `��A��������5��:͇��b������҆�����J����.��۸��]A��Yȕ�N��uҘ��U���כ�Y��fٞ��X��{ס�U���Ҥ��O��̧�#H���ê�@?��^���v5��v���{+�������!��5����������"��捼�R���  �  0}N=�M=G�L=I>L=�}K=�J=��I=�9I=wH=	�G=H�F=�+F=�fE=РD=�C=�C=JB=��A=H�@=��?=V?=�P>=Ӂ==��<=O�;=�;=M9:=�c9=_�8=|�7=��6=��5={5=p>4=n\3=Wx2=,�1=é0=�/=��.=q�-=Z�,=��+=&+=�	*=�)=�(=>	'=�&=�$=��#=m�"=W�!=�� =2�=�t=�Q=�*=��=��=K�=�e=�)=��=n�=�\=\=��=�g=�=�=tJ
=��=Cv=�=��=k=��=` =^%�<��<���<���<A��<lw�<x>�<���<��<�j�<��<#��<�^�<��<���<g �<��<3�<���<4�<{��<*%�<F��<$�<�t�<�ި<)F�<��<��<�n�<͖<�*�<��<�<<�<l��<C�<��z<�>s<��k<��d<YT]<�V<��N< wG<*2@<b�8<�1<{w*<mA#<�<��<�<j�<��;
��;���;���;r��;�޸;
�;rH�;���;�;r�h;�$N;z3;W ;r�:hK�:��:a�D:蛽9���%�ӹ��L��\��x�Ǻ���n���+��HB�6Y���o�� ���.����(ࣻ��������_û��ͻ`�׻*���p뻁�������	���B����:����1���:#� s'�I�+���/���3���7��;�
�?�A�C��WG��K�^�N�֋R�?3V��Y��e]��`��sd���g�Fak�^�n�*0r��u��x��2|�n|�$`��G��������5��A͇��b������φ�����K����.��⸒�TA��\ȕ�	N��wҘ��U���כ�Y��bٞ��X��{ס��U���Ҥ��O��̧�%H���ê�0?��c���{5������}+�������!��'������̔��$���@���  �  '}N=�M=H�L=C>L=�}K=�J=��I=�9I=%wH=�G=K�F=�+F=�fE=נD=�C=�C=JB=��A=I�@=��?=\?=�P>=؁==��<=L�;=�;=P9:=�c9=V�8=��7=��6=��5=w5=m>4=m\3=Ux2=.�1=��0=�/=��.=r�-=Y�,=��+=.+=�	*=�)=�(=C	'=�&=�$= �#=j�"=[�!=�� =4�=�t=�Q=�*=��=��=H�=�e=�)=��=t�=�\=Y=��=�g=�=�=uJ
=��=Gv=�=��=h=��=] =S%�<��<���<���<4��<qw�<�>�<���<��<�j�<��<"��<�^�<��<���<f �<	��<*3�<���<4�<{��<&%�<L��<�<�t�<�ި<-F�<��<��<�n�<|͖<�*�<��<
�<<�<i��<I�<��z<�>s<��k<��d<?T]<�V<��N<wG<92@<;�8< �1<}w*<WA#<�<��<(�<i�<��;���;��;���;m��;�޸;�	�;�H�;���;�;��h;�$N;lz3;Q ;�r�:9K�:ď�:�D:���9ῷ6�ӹ��L�]��+�Ǻb�������+��HB��5Y��o�x ���.����(ࣻ����b���_ûӘͻ{�׻���p�y�������	����B����:���� ���:#�s'�U�+���/���3���7��;��?�L�C�XG��K�f�N�ߋR�93V�!�Y�ze]�&�`��sd���g�Oak�g�n�>0r��u�1�x��2|��|�`��?��������5��G͇��b������ņ�����L����.��긒�EA��bȕ��M��wҘ��U���כ�Y��Sٞ��X��wס�yU���Ҥ��O��#̧�H���ê�)?��g���~5��{����+�������!��$������ɔ��'��􍼼8���  �  '}N=�M=F�L=F>L=�}K=�J=��I=�9I=!wH=
�G=K�F=�+F=�fE=נD=�C=�C=JB=��A=K�@=��?=Y?=�P>=Ё==��<=Q�;=�;=M9:=�c9=V�8=y�7=��6=��5=y5=l>4=h\3=Wx2='�1=��0=�/=��.=p�-=U�,=��+='+=�	*=�)=�(=>	'=�&=�$=��#=o�"=V�!=�� =5�=�t=�Q=�*=��=��=M�=�e=�)=��=m�=�\=[=��=�g=�=�=rJ
=��=Ev=�=��=g=��=[ =V%�<��<���<���<1��<ow�<w>�<���<��<�j�<��<+��<�^�<��<���<\ �<��<%3�<���<4�<���<+%�<J��<%�<�t�<�ި<!F�<��<��<�n�<}͖<�*�<��<��<<�<e��<L�<��z<�>s<��k<t�d<CT]<�V<��N<wG<2@<=�8<�1<vw*<bA#<
<��<�<��<��;��;��;���;���;�޸;�	�;�H�;�;��;��h;�$N;Ez3;� ;�q�:�K�:i��:�D:�9鿷W�ӹd�L��\����Ǻ������!+��HB�_6Y���o�w ���.����Hࣻ��������_û��ͻT�׻*���p�N�������	����A�����9����"���:#�)s'�B�+���/���3���7��;��?�A�C��WG��K�e�N��R�C3V��Y��e]��`��sd���g�`ak�n�n�50r��u�$�x��2|��|� `��G��������5��?͇��b������ǆ�����H����.��ظ��JA��^ȕ��M��oҘ��U���כ�Y��[ٞ��X���ס�~U���Ҥ��O��!̧� H���ê�5?��e����5��x����+�������!��4������Ŕ��,������E���  �  3}N=�M=G�L=A>L=�}K=�J=��I=�9I=wH=�G=L�F=�+F=�fE=РD=&�C=�C=JB=��A=N�@=��?=R?=�P>=ҁ==��<=H�;=�;=M9:=�c9=_�8=w�7=��6=��5=v5=m>4=h\3=Xx2="�1=��0=�/=��.=o�-=U�,=��+=&+=�	*=�)=�(=A	'=�&=�$=��#=u�"=V�!=�� =0�=�t=�Q=�*=��=��=S�=�e=�)=��=o�=�\=S=��=�g=�=�=pJ
=��=;v=�=��=h=��=Z =S%�<��<���<���<=��<qw�<w>�<���<���<�j�<��</��<�^�<��<ɏ�<f �<"��<3�<Ƶ�<4�<}��<7%�<K��<3�<�t�<�ި<&F�<��<��<yn�<�͖<�*�<��<��<<�<c��<8�<��z<|>s<��k<k�d<NT]<�V<��N< wG<2@<k�8<�1<zw*<LA#<�<��<�<��<T�;>��;��;н�;���;�޸;q
�;hH�;��;"�;��h;�$N;�y3;� ;r�:L�:D��:�D:O��9�濷ɺӹ��L�(\���Ǻ~������+��HB��6Y���o�� ���.�� ��Jࣻb�������_û��ͻc�׻���p�[������	����A�����9����:���:#�#s'�(�+���/���3���7���;��?�a�C��WG��K�J�N��R�M3V��Y��e]��`�td���g�[ak�r�n�:0r�"�u��x��2|�r|�`��F��������5��9͇��b������ц�����@����.��и��ZA��Eȕ�N��tҘ��U���כ�Y��oٞ��X��~ס�wU���Ҥ��O��̧�"H���ê�:?��c����5�������+�������!��8������Ք��0��퍼�J���  �  (}N=�M=H�L=E>L=�}K=�J=��I=�9I=$wH=�G=G�F=�+F=�fE=ՠD=#�C=�C=JB=��A=H�@=��?=\?=�P>=ց==��<=J�;=�;=M9:=�c9=W�8=w�7=��6=��5=v5=i>4=e\3=Tx2=#�1=��0=�/=��.=j�-=S�,=��+=&+=�	*=�)=�(=D	'=�&=�$= �#=s�"=U�!=�� =6�=�t=�Q=�*=��=��=N�=�e=*=��=r�=�\=Y=��=�g=�=�=jJ
=��=Av=�=��=d=�=W =R%�<��<���<���<1��<`w�<x>�<���<��<�j�<��<-��<�^�<��<���<d �<��<$3�<õ�<4�<���<.%�<B��<3�<�t�<�ި<,F�<��<��<�n�<�͖<�*�<��<��<	<�<j��<?�<��z<~>s<��k<i�d<@T]<�V<��N<wG<2@<A�8<ڱ1<{w*<\A#<�<��<#�<��<��;B��;���;���;���;�޸;[
�;�H�;��;�;��h;�$N;z3;� ;�r�:�K�:���:��D:d��9��2�ӹ��L�5]��Q�Ǻf���Ο�L+��HB��6Y���o�� ���.��G��Zࣻ��������_ûȘͻ\�׻����p�4�������	����A�����9���� ���:#�"s'�:�+���/���3���7��;��?�I�C��WG��K�w�N��R�`3V�!�Y��e]��`�td���g�iak�z�n�;0r��u�3�x��2|��|�.`��E��������5��;͇��b�������������J����.��Ը��JA��Iȕ� N��kҘ��U���כ�Y��Sٞ��X��xס�xU���Ҥ��O��̧�(H���ê�:?��o���}5�������+�������!��9������є��'������H���  �  '}N=�M=C�L=D>L=�}K=�J=��I=�9I=#wH=	�G=S�F=�+F=�fE=٠D=�C=�C=JB=��A=Q�@=��?=Y?=�P>=Ӂ==��<=V�;=�;=M9:=�c9=X�8=�7=��6=��5=o5=k>4=g\3=Ux2=)�1=��0=
�/=��.=m�-=[�,=��+=-+=�	*=�)=�(=A	'=�&=�$=��#=n�"=b�!=�� =7�=�t=�Q=�*=��=��=L�=�e=�)=��=p�=�\=^=��=�g=�=�=oJ
=��=@v=�=��=f=�=Y =A%�<��<���<���<5��<kw�<{>�<���<��<�j�<��<"��<�^�<��<ɏ�<r �<��<-3�<���<#4�<���</%�<\��<"�<�t�<�ި<'F�<��<��<�n�<v͖<�*�< ��<
�<<�<_��<:�<��z<�>s<��k<w�d<>T]<zV<��N<�vG<92@<<�8<�1<kw*<\A#<<��<�<w�<��;��;W��;ƽ�;���;�޸;	
�;�H�;ך�;D�;�h;�$N;Kz3;~ ;Rr�:|K�:��:9�D:���9�ۿ��ӹ��L�W]����ǺR������-+��HB�86Y�>�o�� ���.��2��ࣻÃ��e���_û��ͻ^�׻���p�]�������	�ޭ��A�����9�������:#��r'�B�+���/���3���7���;�
�?�1�C�XG��K�u�N�ԋR�L3V�*�Y��e]�5�`��sd���g�bak�r�n�]0r��u�8�x��2|��|�#`��A���Û���5��C͇��b������Ɇ�����@����.��ݸ��BA��\ȕ��M��nҘ��U���כ�Y��Xٞ��X��}ס�U���Ҥ��O��)̧�H���ê�)?��r����5�������+�������!��2������ٔ��/������8���  �  &}N=�M=D�L=@>L=�}K=�J=��I=�9I=$wH=�G=Q�F=�+F=�fE=ݠD=%�C=�C=JB=��A=P�@=��?=\?=�P>=ف==��<=M�;=�;=M9:=�c9=V�8=v�7=��6=��5=t5=k>4=b\3=Rx2=�1=��0=�/=��.=h�-=T�,=��+=,+=�	*=�)=�(=E	'=�&=�$=��#=r�"=^�!=�� =5�=u=�Q=�*=��=��=P�=�e=*=��=t�=�\=W=��=�g=�=�=hJ
=��==v=�=��=b=�=V =M%�<��<���<���<,��<dw�<x>�<���<��<�j�<��<1��<�^�<��<ˏ�<m �<��<.3�<ȵ�<*4�<~��<-%�<W��<)�<�t�<�ި<5F�<��<��<{n�<y͖<�*�<���<��<<�<f��<;�<��z<g>s<��k<V�d<DT]<�V<��N<wG<2@<6�8<��1<nw*<GA#<�<��<1�<��<��;"��;A��;���;���;߸;p
�;�H�;Қ�;7�;
�h;�$N;}z3;� ;"s�:�K�:��:	�D:R��9����ӹ��L��\����Ǻ�������x+��HB��6Y���o�� ���.��U��RࣻɃ��t���_û֘ͻi�׻�Ữp�*�������	����A�����9�������:#�s'�3�+���/���3�}�7��;��?�N�C�
XG��K�y�N��R�g3V��Y��e]��`�td���g�qak�~�n�C0r��u�)�x��2|��|�(`��D���Û���5��B͇��b�������������>����.��߸��AA��Cȕ��M��sҘ��U���כ�Y��Uٞ��X��oס�yU���Ҥ��O��&̧�H���ê�9?��s����5�������+�������!��B������֔��*������J���  �  ,}N=�M=J�L=G>L=�}K=�J=��I=�9I="wH=�G=I�F=�+F=�fE=ԠD=�C=�C=JB=��A=I�@=��?=X?=�P>=Ӂ==��<=M�;=�;=M9:=�c9=_�8=w�7=��6=��5=u5=g>4=e\3=]x2=�1=��0=�/=��.=l�-=Z�,=��+=$+=�	*=�)=�(=>	'=�&=�$=��#=r�"=X�!=�� =8�=�t=�Q=�*=��=��=N�=�e=�)=��=m�=�\=Y=��=�g=�=�=mJ
=��=7v=�=��=j=�=R =Q%�<��<���<���<C��<bw�<v>�<���<��<�j�<��<��<�^�<��<�<l �<"��< 3�<���<4�<���<=%�<I��</�<�t�<�ި<!F�<
��<��<�n�<�͖<�*�<	��< �<<�<g��<4�<��z<i>s<��k<Z�d<@T]<wV<��N<wG<2@<P�8<ձ1<�w*<fA#<�<��<�<v�<��;A��;��;��;���;�޸;(
�;�H�; ��;I�;��h;�$N;Dz3;h ;Tr�:�K�:���:3�D:y��92��O�ӹ��L��\��9�Ǻ������@+�EHB��6Y���o�� ��}.��9��ࣻ��������_û��ͻV�׻&��q�j�������	����A�����9�������:#�s'�:�+���/���3���7��;��?�E�C��WG��K�h�N�ʋR�V3V��Y��e]��`�"td���g�aak���n�<0r�)�u�'�x��2|�e|�+`��F��������5��=͇��b������ˆ�����G����.��ϸ��NA��Rȕ�N��dҘ��U���כ�
Y��Wٞ��X���ס��U���Ҥ��O��̧�.H���ê�3?��m����5�������+�������!��A������ڔ��-������E���  �  &}N=�M=D�L=@>L=�}K=�J=��I=�9I=$wH=�G=Q�F=�+F=�fE=ݠD=%�C=�C=JB=��A=P�@=��?=\?=�P>=ف==��<=M�;=�;=M9:=�c9=V�8=v�7=��6=��5=t5=k>4=b\3=Rx2=�1=��0=�/=��.=h�-=T�,=��+=,+=�	*=�)=�(=E	'=�&=�$=��#=r�"=^�!=�� =5�=u=�Q=�*=��=��=P�=�e=*=��=t�=�\=W=��=�g=�=�=hJ
=��==v=�=��=b=�=V =M%�<��<���<���<,��<dw�<x>�<���<��<�j�<��<1��<�^�<��<ˏ�<m �<��<.3�<ȵ�<*4�<~��<-%�<W��<(�<�t�<�ި<5F�<��<��<{n�<y͖<�*�<���<��<<�<f��<;�<��z<g>s<��k<V�d<DT]<�V<��N<wG<2@<6�8<��1<nw*<GA#<�<��<1�<��<��;"��;A��;���;���;߸;p
�;�H�;Қ�;7�;	�h;�$N;}z3;� ;!s�:�K�:��:�D:K��9O��ӹ��L��\����Ǻ�������x+��HB��6Y���o�� ���.��U��RࣻɃ��t���_ûטͻi�׻�ữp�+�������	����A�����9�������:#�s'�3�+���/���3�~�7��;��?�N�C�
XG��K�y�N��R�g3V��Y��e]��`�td���g�qak�}�n�C0r��u�)�x��2|��|�(`��D���Û���5��B͇��b�������������>����.��߸��AA��Cȕ��M��sҘ��U���כ�Y��Uٞ��X��oס�yU���Ҥ��O��&̧�H���ê�9?��s����5�������+�������!��B������֔��*������J���  �  '}N=�M=C�L=D>L=�}K=�J=��I=�9I=#wH=	�G=S�F=�+F=�fE=٠D=�C=�C=JB=��A=Q�@=��?=Y?=�P>=Ӂ==��<=V�;=�;=M9:=�c9=X�8=�7=��6=��5=o5=k>4=g\3=Ux2=)�1=��0=
�/=��.=m�-=[�,=��+=-+=�	*=�)=�(=A	'=�&=�$=��#=n�"=b�!=�� =7�=�t=�Q=�*=��=��=L�=�e=�)=��=p�=�\=^=��=�g=�=�=oJ
=��=@v=�=��=f=�=Y =A%�<��<���<���<5��<kw�<|>�<���<��<�j�<��<"��<�^�<��<ɏ�<r �<��<-3�<���<#4�<���</%�<\��<"�<�t�<�ި<'F�<��<��<�n�<u͖<�*�< ��<
�<<�<_��<:�<��z<�>s<��k<w�d<>T]<zV<��N<�vG<92@<=�8<�1<kw*<\A#<<��<�<w�<��;��;X��;ƽ�;���;�޸;	
�;�H�;ך�;D�;�h;�$N;Jz3;} ;Or�:zK�:
��:3�D:~��9�ܿ��ӹ��L�[]����ǺU������.+��HB�96Y�?�o�� ���.��2��ࣻă��e���_û��ͻ^�׻���p�]�������	�ޭ��A�����9�������:#��r'�B�+���/���3���7���;�
�?�1�C�XG��K�u�N�ԋR�L3V�*�Y��e]�6�`��sd���g�bak�r�n�]0r��u�8�x��2|��|�#`��A���Û���5��C͇��b������Ɇ�����@����.��ݸ��BA��\ȕ��M��nҘ��U���כ�Y��Xٞ��X��}ס�U���Ҥ��O��)̧�H���ê�)?��r����5�������+�������!��2������ٔ��/������8���  �  (}N=�M=H�L=E>L=�}K=�J=��I=�9I=$wH=�G=G�F=�+F=�fE=ՠD=#�C=�C=JB=��A=H�@=��?=\?=�P>=ց==��<=J�;=�;=M9:=�c9=W�8=w�7=��6=��5=v5=i>4=e\3=Tx2=#�1=��0=�/=��.=j�-=S�,=��+=&+=�	*=�)=�(=D	'=�&=�$= �#=s�"=U�!=�� =6�=�t=�Q=�*=��=��=N�=�e=*=��=s�=�\=Y=��=�g=�=�=kJ
=��=Av=�=��=e=�=X =R%�<��<���<���<1��<`w�<x>�<���<��<�j�<��<-��<�^�<��<���<d �<��<$3�<õ�<4�<���<.%�<B��<3�<�t�<�ި<,F�<��<��<�n�<�͖<�*�<��<��<	<�<j��<?�<��z<~>s<��k<i�d<@T]<�V<��N<wG<2@<A�8<۱1<{w*<\A#<�<��<$�<��<��;C��;���;���;���;�޸;[
�;�H�;��;�;��h;�$N;~z3;� ;�r�:�K�:���:��D:R��96��D�ӹ��L�9]��U�Ǻj���П�N+��HB��6Y���o�� ���.��G��[ࣻ��������_ûɘͻ\�׻����p�4�������	����A�����9���� ���:#�"s'�:�+���/���3���7��;��?�I�C��WG��K�w�N��R�`3V�!�Y��e]��`�td���g�iak�z�n�;0r��u�3�x��2|��|�.`��E��������5��;͇��b�������������J����.��Ը��JA��Iȕ� N��kҘ��U���כ�Y��Sٞ��X��xס�xU���Ҥ��O��̧�(H���ê�:?��o���}5�������+�������!��9������є��'������H���  �  3}N=�M=G�L=A>L=�}K=�J=��I=�9I=wH=�G=L�F=�+F=�fE=РD=&�C=�C=JB=��A=N�@=��?=R?=�P>=ҁ==��<=H�;=�;=M9:=�c9=_�8=w�7=��6=��5=v5=m>4=h\3=Xx2="�1=��0=�/=��.=o�-=U�,=��+=&+=�	*=�)=�(=A	'=�&=�$=��#=u�"=V�!=�� =0�=�t=�Q=�*=��=��=S�=�e=�)=��=o�=�\=S=��=�g=�=�=pJ
=��=<v=�=��=h=��=Z =T%�<��<���<���<=��<qw�<x>�<���<���<�j�<��<0��<�^�<��<ɏ�<f �<"��<3�<Ƶ�<4�<}��<6%�<K��<3�<�t�<�ި<&F�<��<��<yn�<�͖<�*�<��<��<<�<b��<8�<��z<|>s<��k<k�d<NT]<�V<��N<!wG<2@<k�8<�1<zw*<MA#<�<��<�<��<T�;>��;��;ѽ�;���;�޸;q
�;hH�;��;!�;��h;�$N;�y3;� ;r�:�K�:?��:؅D::��9�翷ߺӹ��L�-\��"�Ǻ�������+��HB��6Y���o�� ���.��!��Jࣻc�������_û��ͻc�׻���p�[������	����A�����9����:���:#�#s'�(�+���/���3���7���;��?�a�C��WG��K�J�N��R�M3V��Y��e]��`�td���g�[ak�r�n�:0r�"�u��x��2|�r|�`��F��������5��9͇��b������ц�����@����.��и��ZA��Eȕ�N��tҘ��U���כ�Y��oٞ��X��~ס�wU���Ҥ��O��̧�"H���ê�:?��c����5�������+�������!��8������Ք��0��퍼�J���  �  '}N=�M=F�L=F>L=�}K=�J=��I=�9I=!wH=
�G=K�F=�+F=�fE=נD=�C=�C=JB=��A=K�@=��?=Y?=�P>=Ё==��<=Q�;=�;=M9:=�c9=V�8=y�7=��6=��5=y5=l>4=h\3=Wx2='�1=��0=�/=��.=p�-=U�,=��+='+=�	*=�)=�(=>	'=�&=�$=��#=o�"=V�!=�� =5�=�t=�Q=�*=��=��=M�=�e=�)=��=m�=�\=[=��=�g=�=�=sJ
=��=Ev=�=��=g=��=[ =W%�<��<���<���<2��<ow�<w>�<���<��<�j�<��<+��<�^�<��<���<\ �<��<%3�<���<4�<���<+%�<J��<%�<�t�<�ި<!F�<��<��<�n�<}͖<�*�<��<��<<�<e��<L�<��z<�>s<��k<t�d<CT]<�V<��N<wG<2@<=�8<�1<vw*<cA#<
<��<�<��<��;��;��;���;���;�޸;�	�;�H�;�;��;��h;�$N;Cz3;� ;�q�:�K�:d��:��D:ٛ�9�꿷p�ӹp�L��\����Ǻ"������$+��HB�a6Y���o�x ���.����Iࣻ��������_û��ͻT�׻*���p�O�������	����A�����9����"���:#�)s'�B�+���/���3���7��;��?�B�C��WG��K�e�N��R�C3V��Y��e]��`��sd���g�`ak�n�n�50r��u�$�x��2|��|� `��G��������5��?͇��b������ǆ�����H����.��ظ��JA��^ȕ��M��oҘ��U���כ�Y��[ٞ��X���ס�~U���Ҥ��O��!̧� H���ê�5?��e����5��x����+�������!��4������Ŕ��,������E���  �  '}N=�M=H�L=C>L=�}K=�J=��I=�9I=%wH=�G=K�F=�+F=�fE=נD=�C=�C=JB=��A=I�@=��?=\?=�P>=؁==��<=L�;=�;=P9:=�c9=V�8=��7=��6=��5=w5=m>4=m\3=Ux2=.�1=��0=�/=��.=r�-=Y�,=��+=.+=�	*=�)=�(=C	'=�&=�$= �#=j�"=[�!=�� =4�=�t=�Q=�*=��=��=H�=�e=�)=��=t�=�\=Y=��=�g=�=�=uJ
=��=Hv=�=��=h=��=] =S%�<��<���<���<4��<qw�<�>�<���<��<�j�<��<"��<�^�<��<���<f �<	��<*3�<���<4�<{��<&%�<L��<�<�t�<�ި<-F�<��<��<�n�<{͖<�*�<��<
�<<�<h��<I�<��z<�>s<��k<��d<?T]<�V<��N<wG<92@<;�8<�1<~w*<WA#<�<��<)�<i�<��;���;��;���;m��;�޸;�	�;�H�;���;�;��h;�$N;iz3;O ;�r�:4K�:���:�D:g��9�⿷O�ӹ��L�]��1�Ǻh�������+��HB��5Y��o�y ���.����)ࣻ����b���_ûԘͻ|�׻���p�y�������	����B����:���� ���:#�s'�U�+���/���3���7��;��?�L�C�XG��K�f�N�ߋR�93V�!�Y�ze]�&�`��sd���g�Oak�g�n�>0r��u�1�x��2|��|�`��?��������5��G͇��b������ņ�����L����.��긒�EA��bȕ��M��wҘ��U���כ�Y��Sٞ��X��wס�yU���Ҥ��O��#̧�H���ê�)?��g���~5��{����+�������!��$������ɔ��'��􍼼8���  �  0}N=�M=G�L=I>L=�}K=�J=��I=�9I=wH=	�G=H�F=�+F=�fE=РD=�C=�C=JB=��A=H�@=��?=V?=�P>=Ӂ==��<=O�;=�;=M9:=�c9=_�8=|�7=��6=��5={5=p>4=n\3=Wx2=,�1=é0=�/=��.=q�-=Z�,=��+=&+=�	*=�)=�(=>	'=�&=�$=��#=m�"=W�!=�� =2�=�t=�Q=�*=��=��=K�=�e=�)=��=n�=�\=\=��=�g=�=�=tJ
=��=Cv=�=��=k=��=` =^%�<��<���<���<B��<lw�<y>�<���<��<�j�<��<#��<�^�<��<���<g �<��<3�<���<4�<{��<*%�<E��<$�<�t�<�ި<)F�<��<��<�n�<͖<�*�<��<�<<�<l��<C�<��z<�>s<��k<��d<YT]<�V<��N< wG<*2@<b�8<�1<|w*<mA#<�<��<�<j�<��;��;���;���;r��;�޸;
�;rH�;���;�;q�h;�$N;z3;U ;r�:bK�:
��:U�D:ћ�9u��>�ӹ��L��\��~�Ǻ	���q���+��HB�6Y���o�� ���.����)ࣻ��������_û��ͻ`�׻+���p뻁�������	���B����:����1���:#� s'�I�+���/���3���7��;�
�?�A�C��WG��K�^�N�֋R�?3V��Y��e]��`��sd���g�Fak�^�n�*0r��u��x��2|�n|�$`��G��������5��A͇��b������φ�����K����.��⸒�TA��\ȕ�	N��wҘ��U���כ�Y��cٞ��X��{ס��U���Ҥ��O��̧�%H���ê�0?��c���{5������}+�������!��'������̔��$���@���  �  2}N=�M=J�L=A>L=�}K=�J=��I=�9I=wH=
�G=F�F=�+F=�fE=ΠD=�C=�C=JB=��A=G�@=��?=S?=�P>=с==��<=H�;=�;=Q9:=�c9=_�8=s�7=��6=��5=�5=m>4=j\3=bx2=$�1=ǩ0=�/=��.=p�-=U�,=��+='+=�	*=�)=�(=?	'=�&=�$=��#=p�"=P�!=�� =0�=�t=�Q=�*=��=��=N�=�e=�)=��=o�=�\=T=��=�g=�=�=qJ
=��=Ev=�=��=s=��=\ =k%�<��<���<���<@��<qw�<�>�<���< ��<�j�<��<7��<�^�<��<���<R �<��<3�<���<4�<|��<"%�<?��<)�<�t�<�ި<(F�<��<��<yn�<�͖<�*�<��<��<<�<q��<O�<��z<�>s<��k<t�d<ZT]<�V<��N<1wG<2@<h�8<�1<�w*<NA#<�<��<�<��<w�;��;���;}��;��;�޸;
�;SH�;ٚ�;��;`�h;�$N;�y3;� ;�q�:�K�:!��:��D:D��9Y���[�ӹ,�L��[��~�ǺO������+�HB��6Y�V�o�� ��n.����Nࣻ��������_û��ͻ[�׻*���p�Z��ة���	�*��B����:����B���:#�Bs'�>�+���/���3���7��;���?�`�C��WG��K�X�N��R�N3V���Y��e]���`�td���g�Kak�r�n�0r��u��x��2|�r|� `��A��������5��:͇��b������҆�����J����.��۸��]A��Yȕ�N��uҘ��U���כ�Y��fٞ��X��{ס�U���Ҥ��O��̧�#H���ê�@?��^���v5��v���{+�������!��5����������"��捼�R���  �  0}N=�M=J�L=B>L=�}K=�J=��I=�9I=wH=�G=J�F=�+F=�fE=͠D=�C=�C=JB=��A=J�@=��?=S?=�P>=ρ==��<=M�;=�;=Q9:=�c9=`�8=��7=��6=��5=|5=r>4=n\3=ax2=,�1=ũ0=�/=��.=w�-=]�,=��+=,+=�	*=�)=�(=@	'=�&=�$=��#=i�"=W�!=�� =.�=�t=�Q=�*=��=��=H�=�e=�)=��=o�=�\=Z=��=�g=�=�=zJ
=��=Fv=�=��=s=��=a =b%�<��<���<���<H��<sw�<�>�<���<��<�j�<��<!��<�^�<���<���<\ �<��<3�<���<4�<u��<"%�<I��<�<�t�<�ި<F�<��<��<}n�<�͖<�*�<��<
�<!<�<e��<K�<��z<�>s<��k<��d<cT]<�V<��N<7wG<92@<d�8<��1<�w*<QA#<�<��<�<p�<�;���;��;���;d��;�޸;�	�;ZH�;���;��;��h;'$N;�y3;G ;�q�:�K�:���: �D:W��9��ӹ��L��[�� �Ǻ����c���+�HB�!6Y�u�o�� ���.�����ࣻ����y���_û�ͻk�׻%��q뻅������	���B����:�Þ�D���:#�(s'�W�+���/���3���7��;��?�L�C��WG��K�]�N�ȋR�+3V�
�Y��e]���`��sd���g�Aak�]�n�$0r��u�
�x��2|�d|�`��<��������5��?͇��b������Ն�����L����.��丒�ZA��aȕ�N��|Ҙ��U���כ�"Y��eٞ��X���ס�U���Ҥ��O��̧�H���ê�*?��X����5��z���z+�������!��*������Ɣ��-��㍼�9���  �  *}N=�M=E�L=J>L=�}K=�J=��I=�9I=%wH=�G=F�F=�+F=�fE=РD=�C=�C=JB=��A=D�@=��?=\?=�P>=ف==��<=O�;=�;=N9:=�c9=Y�8=~�7=��6=��5=|5=r>4=p\3=Xx2=/�1=��0=�/=��.=q�-=X�,=��+=*+=�	*=�)=�(=C	'=�&=�$=��#=i�"=U�!=�� =1�=�t=�Q=�*=��=��=F�=�e=�)=��=u�=�\=a=��=�g=�=�=tJ
=��=Pv=�=��=k=��=c =b%�<�<���<���<=��<ow�<>�<���<��<�j�<��<��<�^�<���<���<Z �<��< 3�<���<4�<y��<%�<B��<�<�t�<�ި<-F�<	��<��<�n�<|͖<�*�<��<�<<�<y��<T�<��z<�>s<��k<��d<QT]<�V<׾N<wG<32@<I�8<�1<tw*<tA#<�<��<*�<k�<��;���;���;]��;i��;�޸;�	�;zH�;���;��;*�h;$N;^z3;3 ;�r�:�J�:돕:9�D:���9����q�ӹ�L��\��Z�Ǻ����h���+��HB��5Y���o�J ���.����9ࣻ��������_û��ͻ��׻���p�j�������	���'B����:����5��;#�,s'�_�+���/���3���7��;�$�?�/�C��WG��K�h�N�ۋR�B3V��Y�^e]�
�`��sd���g�Gak�W�n�'0r�،u�!�x��2|�{|�#`��B��������5��K͇��b�����������V����.���PA��bȕ�N��yҘ��U���כ�#Y��Tٞ��X��wס��U���Ҥ��O��"̧� H���ê�/?��c���n5��p����+�������!�� ����������������<���  �  0}N=�M=H�L=E>L=�}K=�J=��I=�9I=wH=�G=I�F=�+F=�fE=ɠD=�C=�C=JB=��A=H�@=��?=T?=�P>=Ձ==��<=J�;=�;=Q9:=�c9=_�8=��7=��6=��5={5=o>4=t\3=dx2=0�1=��0=�/=��.=u�-=]�,=��+=/+=�	*=�)=�(=A	'=�&=�$=��#=m�"=T�!=�� =-�=�t=�Q=�*=��=��=L�=�e=�)=��=s�=�\=Y=��=�g=�=�=xJ
=��=Mv=�=��=v=�=` =`%�<�<���<���<J��<�w�<�>�<���<��<�j�<��<��<�^�<���<���<V �<��<3�<���<4�<y��<%�<D��<�<�t�<�ި<&F�<	��<��<�n�<~͖<�*�<��<	�<<�<v��<Q�<��z<�>s<��k<��d<NT]<�V<;N<)wG<72@<d�8<�1<�w*<`A#<�<��<�<g�<t�;���;���;r��;n��;k޸;�	�;*H�;���;��;f�h;$N;�y3; ;Er�:�J�:?��:u�D:��9�ſ�P�ӹ#�L��\����Ǻ������+��GB��5Y���o�` ��p.�����ࣻm���c���_ûژͻ��׻��q뻔�������	���B����":�ɞ�O���:#�5s'�I�+�¹/���3���7���;��?�N�C��WG��K�G�N�R�43V���Y�ke]��`��sd�z�g�2ak�c�n�+0r��u��x��2|�a|�`��;��������5��H͇��b������҆�����K����.��渒�dA��gȕ�N��yҘ��U���כ�Y��gٞ��X��}ס��U���Ҥ��O�� ̧�H���ê�*?��^���r5��t����+�������!��������Ŕ����ꍼ�:���  �  �yN=#�M=�L=i9L=fxK=�J=��I=u2I=\oH=��G=F�F=;"F=q\E=ܕD=��C=2C==B=�rA=ϧ@=��?=T?=�?>=1p==F�<=�;=c�:=J$:=�M9=u8=��7=5�6=��5=�5=�"4=�?3=�Z2=Vs1=�0=�/=��.=S�-=!�,=O�+=��*=n�)=�(=��'=��&=��%=C�$=$�#=��"=��!=�~ =�b=�B=�=��=�=;�=ag=R/=�=��=�m=�$=Y�=��=t/=��=v=�
=O�=d?=C�=�Z=6�=ze=`��<���<��<ٔ�<�s�<�K�<�<���</��<d�<��<���<Ir�<��<ɳ�<wL�<���<�n�<���<]~�<���<}�<���<�l�<�߯<�O�<���<'�<��<���<�X�<���<��<!z�<؋<65�<���<Z�<ߑz<�Hs<��k<c�d<Mp]<q*V<u�N<�G<�e@<�)9<U�1<��*<��#<(a<�:<<}�<d��;���;;��;���;7��;��;/"�;sk�;�ɐ;w;�;�k;U�P;f.6;��;1�;�-�:U��:��P:��9Q��7ul���c?�������������s~'�ߧ>�L�U�v.l��E��~Q���:��� �����Y$��=����˻��ջW�߻��點M����&�&���c����?b�^���#�n"���&���*�)�.�W3��7��;��>���B�бF�}J�o=N�n�Q�Z�U��AY���\�sj`���c��pg���j�Wn� �q� u��yx���{�O�p1��j҂��p��}��ʥ���<���ъ�Ld�����탏���w���~&��ɮ���5������G@���Û�<F���Ǟ�dH��Xȡ�zG��Ƥ�D��q����>��`����7�����D0��[���_(������� ��F������𖹼[��)�������  �  �yN=(�M=��L=c9L=hxK=�J=��I=o2I=YoH=��G=L�F=8"F=p\E=ەD=y�C=6C==B=�rA=ҧ@=��?=S?=�?>=9p==I�<=�;=Z�:=D$:=�M9=�u8=��7=-�6=��5=�5=�"4=�?3=�Z2=[s1=މ0=�/=�.=P�-=$�,=R�+=��*=b�)=�(=��'=��&=�%=?�$= �#=��"=��!=�~ =�b=�B=�=��=�=E�=bg=O/=�=��=�m=�$=[�=��=t/=��=v=�
=F�=g?=<�=�Z=C�=�e=]��<���<��<ǔ�<�s�<�K�<�<���<��<d�<��<���<Dr�<��<Ƴ�<zL�<���<�n�<���<B~�<���<}�<���<	m�<�߯<�O�<���<'�<��<���<�X�<���<�<)z�<$؋<+5�<���<[�<őz<�Hs<��k<��d<7p]<l*V<v�N<ƤG<�e@<�)9<l�1<Ӽ*<��#<2a<�:<5<g�<J��;���;n��;���;,��;��;�!�;�k�;Uɐ;�;�;,�k;N�P;[.6;s�;��;2.�:˘�::�P:���9��7�j��b?�����.���R�����}'�%�>���U��.l��E���Q���:��� ��룬�=$�������˻��ջ�߻_���M����&�����c����jb�����#�.n"�]�&���*�5�.�h3��7�i;���>���B��F�}J�d=N�f�Q�^�U��AY���\��j`���c��pg���j�Wn��q��u� zx���{�A�k1��s҂��p��v��å���<���ъ�Pd�����ꃏ�������v&��䮕��5������R@���Û�<F���Ǟ�pH��Dȡ�nG��Ƥ�
D�������>��W����7��%���I0��Z���l(��~���� ��/������򖹼[��7�������  �  �yN=+�M=��L=i9L=jxK=�J=��I=n2I=aoH=��G=L�F=7"F=p\E=�D=y�C=AC==B=�rA=ͧ@=��?=[?=�?>=6p==A�<=	�;=\�:=G$:=�M9=}u8=��7=)�6=��5=�5=�"4=�?3=�Z2=Xs1=ډ0=!�/=�.=R�-=!�,=M�+=��*=`�)=&�(=��'=��&=�%=D�$='�#=��"=��!=�~ =�b=�B=�=��=�=H�=[g=V/=�=��=�m=�$=a�=��=y/=��=v=�
=C�=o?=9�=�Z=6�=~e=]��<���<)��<���<�s�<�K�<�<���<��<&d�<��<���<?r�<��<˳�<oL�<��<�n�<���<G~�<���<'}�<���<m�<�߯<�O�<���<'�<���<���<�X�<���<�<z�<"؋<)5�<���<f�<��z<�Hs<��k<��d<4p]<|*V<��N<��G<�e@<�)9<u�1<Ӽ*<��#<:a<�:<-<c�<���;i��;j��;y��;3��;(�;�!�;�k�;1ɐ;�;�;�k;Q�P;�.6;O�;��;$-�:h��:��P:���9��78m���a?�(���<������"~'��>�"�U�/l��E���Q���:��� �����$������Ի˻��ջG�߻j�黚M�g��� &�����c����Kb�w���#�Kn"�R�&���*��.�I3��7�z;��>���B��F�}J�t=N�v�Q�S�U��AY�u�\��j`���c��pg���j�Wn��q��u�4zx���{�V�o1��h҂��p��k��ӥ���<���ъ�@d���������������^&��߮���5������W@���Û�FF���Ǟ�nH��Hȡ�G�� Ƥ��C�������>��d����7��'���G0��O���o(������� ��7������ꖹ�U��>�������  �  �yN=$�M=��L=f9L=gxK=�J=��I=p2I=]oH=��G=L�F=@"F=o\E=ܕD=x�C=7C==B=�rA=Χ@=��?=T?=�?>=9p==F�<=�;=]�:=G$:=�M9=u8=��7=.�6=��5=�5=�"4=�?3=�Z2=\s1=ى0=�/=�.=S�-= �,=N�+=��*=c�)=�(=��'=��&=�%=@�$='�#=��"=��!=�~ =�b=�B=�=��=�=G�=]g=V/=�=��=�m=�$=Y�=��=s/=��=v=�
=F�=f?=8�=�Z=>�=�e=b��<���<��<ǔ�<�s�<�K�<�<���<��<d�<��<���<Gr�<��<г�<rL�<	��<�n�<���<A~�<���<}�<���<	m�<�߯<�O�<���<'�<
��<���<�X�<���<��<z�<؋<15�<���<Z�<őz<�Hs<��k<��d<;p]<b*V<q�N<ͤG<�e@<�)9<Z�1<޼*<��#</a<�:</<h�<k��;y��;m��;���;'��;��;�!�;�k�;Dɐ;�;�;��k;z�P;l.6;��;Ö;�-�:���:��P:���9���7ul���b?�~���8���������}'�Z�>��U�'/l��E���Q���:��� �����M$�������˻��ջ�߻f�黹M�m���&�����c����]b�����#�+n"�S�&���*��.�b3��7�i;��>���B���F�}J�t=N�r�Q�V�U��AY���\��j`���c��pg���j�Wn�$�q��u�zx���{�P�v1��l҂��p��{��˥���<���ъ�Pd�����򃏼������s&��宕��5������D@���Û�CF���Ǟ�oH��Iȡ�sG��Ƥ�D�������>��a����7�����L0��[���l(������� ��4����������]��3�������  �  �yN=!�M=��L=f9L=hxK=�J=��I=s2I=XoH=��G=F�F=;"F=s\E=�D=��C=:C==B=�rA=ͧ@=��?=P?=�?>=3p==I�<=�;=_�:=G$:=�M9=�u8=��7=0�6=��5=�5=�"4=�?3=�Z2=Qs1=މ0=�/=�.=M�-=�,=T�+=��*=k�)=�(=��'=��&=�%=?�$=&�#=��"=��!=�~ =�b=�B=�=��=�=A�=cg=V/=�=��=�m=�$=X�=��=p/=��=v=�
=I�=f?==�=�Z=;�=|e=P��<���<��<̔�<�s�<�K�<�<���<&��<d�<��<���<Nr�<��<׳�<tL�<���<�n�<���<V~�<���<#}�<���<�l�<�߯<�O�<���<'�<
��<���<�X�<���<��<.z�<؋</5�<���<^�<z<�Hs<��k<^�d<1p]<r*V<u�N<ФG<�e@<�)9<N�1<�*<��#<0a<�:<%<v�<B��;»�;@��;���;G��;�;"�;�k�;uɐ;�;�;�k;��P;7.6;��;e�;:.�:���:��P:���9��7)i���c?�,���a������<�W~'�|�>���U��.l��E���Q���:��� ��֣��b$��V����˻��ջA�߻^�黾M�r����%����c����Cb�g���#�n"�n�&���*��.�n3��7��;���>���B�ݱF�#}J�_=N�o�Q�p�U��AY���\��j`���c��pg���j�0Wn��q��u�zx���{�;�q1��p҂��p��{��¥���<���ъ�Wd�����������~���m&��Ю���5������I@���Û�0F���Ǟ�hH��Jȡ�tG�� Ƥ�D��y����>��S����7��!���G0��V���n(������� ��H�������[��1�������  �  �yN=#�M=��L=g9L=lxK=�J=��I=u2I=[oH=��G=J�F=?"F=q\E=��D=y�C=<C==B=�rA=Ч@=��?=U?=�?>=2p==I�<=�;=^�:=G$:=�M9=~u8=��7=-�6=��5=�5=�"4=�?3=�Z2=Us1=߉0=�/=�.=S�-=�,=M�+=��*=g�)=�(=��'=��&=�%=B�$=&�#=��"=��!=�~ =�b=�B=�=��=�=G�=`g=U/=�=��=�m=�$=[�=��=r/=��=v=�
=E�=e?==�=�Z=8�=~e=T��<���<��<Ɣ�<�s�<�K�<�<���<"��<d�<��<���<Mr�<��<ѳ�<vL�<��<�n�<���<G~�<���<#}�<���<m�<�߯<�O�<¼�<'�<���<���<�X�<���<��<z�<؋<15�<z��<Y�<Ƒz<�Hs<��k<x�d<5p]<h*V<]�N<ɤG<�e@<�)9<V�1<ܼ*<��#<@a<�:<#<��<[��;���;d��;���;:��;	�;�!�;�k�;Vɐ;�;�;�k;��P;�.6;��;U�;..�:S��:k�P:��9��7�l���a?�������������~'���>�M�U��.l��E���Q���:��� �����O$��t����˻��ջ_�߻Z�黥M�t���&�����c����Mb�v���#�(n"�R�&���*��.�]3��7��;���>���B��F�}J�u=N�u�Q�S�U��AY���\��j`���c��pg���j�&Wn��q�	 u�zx���{�S�s1��n҂��p��r�������<���ъ�Kd��
����	������h&��߮���5������C@���Û�2F���Ǟ�aH��Kȡ�G���Ť� D�������>��c����7�����R0��\���k(������� ��;������󖹼g��5�������  �  �yN=+�M=��L=c9L=cxK=�J=��I=q2I=^oH=��G=K�F=?"F=o\E=�D=|�C=DC==B=�rA=ϧ@=��?=V?=�?>==p==G�<=��;=Z�:=G$:=�M9={u8=��7=*�6=��5=�5=�"4=�?3=�Z2=Xs1=։0=�/=�.=O�-=�,=L�+=��*=d�)=�(=��'=��&=�%==�$=)�#=��"=��!=�~ =�b=�B=�=��=�=J�=]g=W/=�=��=�m=�$=T�=��=v/=��=v=�
=A�=f?=4�=�Z=7�=|e=Q��<���<��<���<�s�<�K�<�<���<��<
d�<��< ��<Fr�<��<ҳ�<tL�<	��<�n�<���<J~�<���<!}�<���<m�<�߯<�O�<���<'�<��<���<�X�<���<�<z�<؋<(5�<|��<Y�<��z<�Hs<��k<��d<p]<d*V<f�N<��G<�e@<�)9<u�1<ּ*<��#<a<�:<D<o�<y��;���;g��;���;.��;G�;�!�;l�;Aɐ;�;�;�k;��P;�.6;��;�;.�:/��:��P:��9\�7$n��Xb?�󌐺����~��T�"~'�§>��U�Z/l��E���Q���:��� �����$������7�˻��ջ�߻G���M�Z���&�����c����Db�r���#�5n"�G�&���*��.�j3��7�h;��>���B���F�	}J�v=N���Q�d�U��AY���\��j`���c��pg���j�*Wn�)�q��u�0zx���{�e�n1��j҂��p�����ǥ���<���ъ�Md���������������\&��ܮ���5������F@���Û�:F���Ǟ�mH��?ȡ�sG��
Ƥ�
D�������>��g����7��(���P0��[���{(������� ��6����������b��<�������  �  �yN="�M=��L=k9L=gxK=�J=��I=t2I=_oH=��G=H�F=A"F=u\E=�D=|�C=?C==B=�rA=ϧ@=��?=V?=�?>=5p==I�<=�;=c�:=A$:=�M9=�u8=��7=-�6=��5=�5=�"4=�?3=�Z2=Ss1=ى0=�/=�.=M�-=�,=O�+=��*=h�)="�(=��'=��&=�%=B�$=,�#=��"=��!=�~ =�b=�B=�=��=�=G�=bg=[/=�=��=�m=�$=[�=��=k/=��=v=�
=C�=c?=7�=�Z=6�=ye=O��<���<��<�<�s�<�K�<�<v��<)��<d�<��<���<Gr�<��<۳�<wL�<��<�n�<���<L~�<���<*}�<���<m�<�߯<�O�<���<'�<��<���<�X�<���<��<!z�<؋<)5�<}��<Y�<��z<�Hs<��k<b�d<p]<b*V<e�N<ĤG<�e@<�)9<Q�1<ϼ*<��#<,a<�:<'<y�<���;���;T��;Ѳ�;a��;;�;�!�;�k�;�ɐ;�;�;�k;��P;�.6;��;��;W.�:�:��P:���9���7�j��Oc?�m�������*��C�m~'�ѧ>�n�U�(/l��E���Q���:��� ������z$��h����˻��ջ0�߻T�黧M�?����%�����c����Bb�q���#�n"�P�&���*��.�[3��7�x;���>���B��F�3}J�q=N�v�Q�m�U��AY���\��j`���c��pg���j�-Wn��q� u�#zx���{�M�t1��z҂��p��x��¥���<���ъ�Ld����샏���z���c&��ٮ���5������>@���Û�3F���Ǟ�gH��Jȡ�rG��Ƥ��C�������>��`����7��'���P0��\���w(������� ��F����������b��7�������  �  �yN=#�M=��L=h9L=gxK=�J=��I={2I=ZoH=��G=N�F=C"F=t\E=ߕD=��C=9C==B=�rA=ԧ@=��?=T?=�?>=2p==M�<=�;=_�:=F$:=�M9=~u8=��7=/�6=��5=�5=�"4=�?3=�Z2=Ps1=݉0=�/=�.=P�-=�,=O�+=��*=g�)=�(=��'=��&=�%=F�$=$�#=��"=��!=�~ =�b=�B=�=��=�=I�=eg=T/=�=��=�m=�$=W�=��=n/=��=v=�
=E�=[?=;�=�Z=;�={e=H��<���<��<Ɣ�<�s�<�K�<�<��<!��<d�<��<���<Vr�<��<ҳ�<}L�<��<�n�<���<U~�<���<'}�<���<m�<�߯<�O�<˼�<'�<��<���<�X�<���<��< z�<؋<05�<w��<M�<��z<�Hs<��k<h�d<*p]<N*V<W�N<ͤG<�e@<�)9<T�1<޼*<��#<-a<�:<!<��<U��;ͻ�;���;��;Y��;�;"�;�k�;ɐ;�;�;`�k;��P;�.6;@�;g�;�.�:���:��P:���9���7sl���c?�C���?���f��W�A~'�g�>���U��.l� F���Q���:��������_$��r����˻��ջ<�߻B�黀M�}����%�����c����Db�j���#�n"�K�&�x�*��.�Q3��7�};���>���B��F�%}J�r=N���Q�f�U��AY���\��j`���c��pg���j�;Wn��q� u�zx���{�Y�u1��q҂��p��~�������<���ъ�Ld�����惏���|���m&��Ѯ���5������<@���Û�-F���Ǟ�WH��Jȡ�pG�� Ƥ�D�������>��`����7�� ���U0��h���o(������� ��B������ ���j��2�������  �  �yN=&�M=��L=h9L=fxK=�J=��I=t2I=^oH=��G=N�F=>"F=w\E=�D=��C=DC==B=�rA=ѧ@=��?=W?=�?>=5p==H�<=�;=]�:=G$:=�M9={u8=��7=%�6=��5=�5=�"4=�?3=�Z2=Ms1=؉0=�/=�.=M�-=�,=L�+=��*=b�)=�(=��'=��&=�%=B�$=*�#=��"=��!=�~ =�b=�B=�=��=�=I�=bg=Z/=�=��=�m=�$=X�=��=u/=��=v=�
=?�=c?=6�=�Z=2�=ue=F��<���<��<���<�s�<�K�<�<���<��<d�<��<���<Ir�<��<ٳ�<yL�<
��<�n�<���<X~�<���<2}�<���<m�<�߯<�O�<���<'�<��<���<�X�<���<�<z�<؋<"5�<|��<Y�<��z<�Hs<��k<S�d<p]<d*V<h�N<��G<�e@<�)9<`�1<׼*<��#<)a<�:<+<}�<w��;���;~��;���;s��;V�;("�;l�;~ɐ;�;�;@�k;��P;�.6;��;��;8.�:ޘ�:i�P:A��9E��7�m���b?�s���g���4��k��~'���>���U�4/l��E���Q���:��� �����&$�������˻��ջ'�߻^�黣M�O����%�����c����/b�[��}#�,n"�J�&���*��.�Y3��7�t;��>���B���F�}J�|=N�{�Q�j�U��AY���\��j`���c��pg���j�>Wn� �q� u�@zx���{�[�v1��k҂��p��y��ȥ���<���ъ�Id�� ���ꃏ�������V&��ͮ���5������G@���Û�1F���Ǟ�eH��Hȡ�rG��Ƥ�D�������>��h����7��-���P0��\���z(������� ��M����������a��D�������  �  �yN=%�M=��L=k9L=hxK=�J=��I=r2I=coH=��G=S�F=D"F=v\E=�D=v�C=BC==B=�rA=ӧ@=��?=Z?=�?>=>p==E�<=�;=^�:=A$:=�M9=|u8=��7=$�6=��5=�5=�"4=�?3=�Z2=Xs1=Ӊ0=�/=�.=K�-=%�,=H�+=��*=^�)=&�(=��'=��&=�%=A�$=-�#=��"=��!=�~ =�b=�B=�=��=�=Q�=^g=[/=�=��=�m=�$=`�=��=p/=��=v=�
==�=b?=/�=�Z=5�=ze=T��<���<��<���<�s�<�K�<�<z��<��<"d�<��<��<Gr�<��<׳�<xL�<��<�n�<���<@~�<���<-}�<���<m�<�߯<�O�<���<!'�<
��<���<�X�<���<�<z�<#؋<5�<z��<M�<��z<�Hs<��k<q�d<p]<E*V<e�N<��G<�e@<�)9<]�1<��*<��#<0a<�:<E<t�<���;���;���;��;e��;H�;�!�;�k�;vɐ;<�;T�k;��P;�.6;��;&�;�-�:p��:��P:��9���7im��0b?�����2���h���/~'�ԧ>��U��/l��E���Q���:��� ��3���I$������ϻ˻��ջ�߻K�黭M�5���&�����c����Fb�z���#�$n"�(�&���*���.�^3��7�^;��>���B��F�}J��=N�`�Q�m�U��AY���\��j`���c��pg���j�!Wn�F�q��u�Czx���{�P�v1��v҂��p��l��Υ���<���ъ�Gd�����냏��������]&��宕��5������=@���Û�<F���Ǟ�iH��>ȡ�sG��Ƥ��C�������>��o����7��2���S0��g���}(������� ��>���������b��H�������  �  �yN='�M=��L=h9L=cxK=�J=��I=y2I=boH=��G=N�F=A"F=w\E=�D=��C=FC==B=�rA=ӧ@=��?=[?=�?>=:p==E�<= �;=^�:=I$:=�M9=zu8=��7=*�6=��5=�5=�"4=�?3=�Z2=Ks1=ى0=�/=�.=G�-=�,=J�+=��*=f�)= �(=��'=��&=
�%=F�$=+�#=��"=��!=�~ =�b=�B=�=��=�=I�=ag=Y/=�=��=�m=�$=Y�=��=t/=��=v=�
=D�=_?=5�=�Z=0�=qe=D��<���<��<���<�s�<�K�<�<���<��<d�<��<���<Qr�<��<ӳ�<wL�<	��<�n�<���<^~�<���</}�<���<m�<�߯<�O�<Ƽ�< '�<��<���<�X�<���<�<z�<؋< 5�<���<I�<��z<~Hs<��k<O�d<p]<F*V<m�N<��G<�e@<�)9<e�1<߼*<��#<a<�:<<<��<���;���;���;Ҳ�;m��;l�;@"�;l�;�ɐ;�;�;U�k;��P;/6;!�;�;�-�:n��:��P:��9��7	n��*d?�ӌ��[������v��~'�	�>�ٍU�/l�	F���Q���:��� ��"���,$��w�����˻��ջ7�߻5�黃M�E����%�����c����b�I���#�n"�I�&���*��.�K3��7�s;��>���B��F�}J��=N���Q���U��AY���\��j`���c��pg���j�AWn�1�q� u�+zx���{�`�s1��h҂��p��~��˥���<���ъ�Ad�����냏���|���V&��Ǯ���5������B@���Û�4F���Ǟ�]H��?ȡ�wG��
Ƥ� D�������>��j����7��/���K0��k���u(������� ��O���������_��A�������  �  �yN=�M=��L=e9L=jxK=��J=��I=u2I=]oH=��G=M�F=C"F=|\E=��D=z�C=>C==B=�rA=֧@=��?=X?=�?>=3p==Q�<=�;=\�:=C$:=�M9=�u8=��7=)�6=��5=�5=�"4=�?3=�Z2=Hs1=��0=�/=�.=I�-=�,=L�+=��*=b�)=�(=��'=��&=�%=B�$=(�#=��"=��!=�~ =�b=�B=�=��=�=F�=kg=X/=�=��=�m=�$=W�=��=k/=��=v=�
=C�=V?=<�=�Z==�={e=C��<���<���<���<�s�<�K�< �<y��<��<d�<��<���<Jr�<��<ڳ�<�L�<��<�n�<���<G~�<���<8}�<���<
m�<�<�O�<���<'�<��<���<�X�<���<��<z�<؋< 5�<z��<G�<��z<tHs<��k<L�d<%p]<K*V<V�N<��G<�e@<�)9<?�1<Ҽ*<��#<9a< ;<'<��<l��;��;~��;��;���;�;�!�;�k�;�ɐ;�;�;��k;�P;�.6;��;y�;o/�:���:S�P:S��9���7Pk��,c?�����g���<��u�R~'�&�>��U��.l�@F���Q���:��� �����r$�������˻��ջ�߻I�黠M�`����%�����c����Pb�|���#�n"�S�&�_�*��.�T3��7�p;���>���B���F�2}J��=N�p�Q�|�U��AY���\��j`��c��pg���j�AWn��q�, u�/zx���{�K��1��w҂��p��|�������<���ъ�Fd����݃����n���b&��ޮ���5������;@���Û�$F���Ǟ�dH��Hȡ�jG���Ť�D�������>��a����7��/���R0��n���m(������� ��P���������j��A�������  �  �yN='�M=��L=h9L=cxK=�J=��I=y2I=boH=��G=N�F=A"F=w\E=�D=��C=FC==B=�rA=ӧ@=��?=[?=�?>=:p==E�<= �;=^�:=I$:=�M9=zu8=��7=*�6=��5=�5=�"4=�?3=�Z2=Ks1=ى0=�/=�.=G�-=�,=J�+=��*=f�)= �(=��'=��&=
�%=F�$=+�#=��"=��!=�~ =�b=�B=�=��=�=I�=ag=Y/=�=��=�m=�$=Y�=��=t/=��=v=�
=D�=_?=6�=�Z=0�=qe=D��<���<��<���<�s�<�K�<�<���<��<d�<��<���<Qr�<��<ӳ�<wL�<	��<�n�<���<^~�<���</}�<���<m�<�߯<�O�<Ƽ�< '�<��<���<�X�<���<�<z�<؋< 5�<���<I�<��z<~Hs<��k<O�d<p]<F*V<m�N<��G<�e@<�)9<e�1<߼*<��#<a<�:<<<��<���;���;���;Ҳ�;m��;l�;@"�;l�;�ɐ;�;�;T�k;��P;/6; �;�;�-�:m��:��P:{��9��7n��-d?�Ԍ��\������w��~'�
�>�ٍU�/l�	F���Q���:��� ��#���,$��w�����˻��ջ7�߻5�黃M�E����%�����c����b�I���#�n"�I�&���*��.�K3��7�s;��>���B��F�}J��=N���Q���U��AY���\��j`���c��pg���j�AWn�1�q� u�+zx���{�`�s1��h҂��p��~��˥���<���ъ�Ad�����냏���|���V&��Ǯ���5������B@���Û�4F���Ǟ�]H��?ȡ�wG��
Ƥ� D�������>��j����7��/���K0��k���u(������� ��O���������_��A�������  �  �yN=%�M=��L=k9L=hxK=�J=��I=r2I=coH=��G=S�F=D"F=v\E=�D=v�C=BC==B=�rA=ӧ@=��?=Z?=�?>=>p==E�<=�;=^�:=A$:=�M9=|u8=��7=$�6=��5=�5=�"4=�?3=�Z2=Xs1=Ӊ0=�/=�.=K�-=%�,=H�+=��*=^�)=&�(=��'=��&=�%=A�$=-�#=��"=��!=�~ =�b=�B=�=��=�=Q�=^g=[/=�=��=�m=�$=`�=��=p/=��=v=�
==�=b?=/�=�Z=5�=ze=T��<���<��<���<�s�<�K�<�<z��<��<"d�<��<��<Gr�<��<׳�<xL�<��<�n�<���<@~�<���<-}�<���<m�<�߯<�O�<���<!'�<
��<���<�X�<���<�<z�<#؋<5�<z��<M�<��z<�Hs<��k<r�d<p]<E*V<e�N<��G<�e@<�)9<]�1<��*<��#<0a<�:<E<t�<���;���;���;��;e��;H�;�!�;�k�;vɐ;<�;T�k;��P;�.6;��;%�;�-�:n��:��P:u��9���7sm��4b?�����4���j���0~'�է>��U��/l��E���Q���:��� ��4���J$������ϻ˻��ջ�߻K�黭M�5���&�����c����Fb�z���#�$n"�(�&���*���.�^3��7�^;��>���B��F�}J��=N�`�Q�m�U��AY���\��j`���c��pg���j�!Wn�F�q��u�Dzx���{�P�v1��v҂��p��l��Υ���<���ъ�Gd�����냏��������]&��宕��5������=@���Û�<F���Ǟ�iH��>ȡ�sG��Ƥ��C�������>��o����7��2���S0��g���}(������� ��>���������b��H�������  �  �yN=&�M=��L=h9L=fxK=�J=��I=t2I=^oH=��G=N�F=>"F=w\E=�D=��C=DC==B=�rA=ѧ@=��?=W?=�?>=5p==H�<=�;=]�:=G$:=�M9={u8=��7=%�6=��5=�5=�"4=�?3=�Z2=Ms1=؉0=�/=�.=M�-=�,=L�+=��*=b�)=�(=��'=��&=�%=B�$=*�#=��"=��!=�~ =�b=�B=�=��=�=I�=bg=Z/=�=��=�m=�$=X�=��=u/=��=v=�
=?�=c?=6�=�Z=2�=ue=F��<���<��<���<�s�<�K�<�<���<��<d�<��<���<Ir�<��<ڳ�<yL�<
��<�n�<���<X~�<���<2}�<���<m�<�߯<�O�<���<'�<��<���<�X�<���<�<z�<؋<"5�<|��<Y�<��z<�Hs<��k<S�d<p]<d*V<h�N<��G<�e@<�)9<`�1<׼*<��#<*a<�:<+<}�<w��;���;~��;���;s��;V�;'"�;l�;~ɐ;�;�;?�k;��P;�.6;��;��;5.�:ۘ�:b�P:4��9n��7�m���b?�v���j���8��l��~'��>���U�6/l��E���Q���:��� �����&$�������˻��ջ'�߻^�黣M�O����%�����c����/b�[��}#�,n"�J�&���*��.�Y3��7�t;��>���B���F�}J�|=N�{�Q�j�U��AY���\��j`���c��pg���j�>Wn� �q� u�@zx���{�[�v1��k҂��p��y��ȥ���<���ъ�Id�� ���ꃏ�������V&��ͮ���5������G@���Û�1F���Ǟ�eH��Hȡ�rG��Ƥ�D�������>��h����7��-���P0��\���z(������� ��M����������a��D�������  �  �yN=#�M=��L=h9L=gxK=�J=��I={2I=ZoH=��G=N�F=C"F=t\E=ߕD=��C=9C==B=�rA=ԧ@=��?=T?=�?>=2p==M�<=�;=_�:=F$:=�M9=~u8=��7=/�6=��5=�5=�"4=�?3=�Z2=Ps1=݉0=�/=�.=P�-=�,=O�+=��*=g�)=�(=��'=��&=�%=F�$=$�#=��"=��!=�~ =�b=�B=�=��=�=I�=eg=T/=�=��=�m=�$=W�=��=n/=��=v=�
=E�=\?=;�=�Z=;�={e=H��<���<��<Ɣ�<�s�<�K�<�<��<!��<d�<��<���<Vr�<��<ҳ�<}L�<��<�n�<���<U~�<���<'}�<���<m�<�߯<�O�<˼�<'�<��<���<�X�<���<��< z�<؋<05�<w��<M�<��z<�Hs<��k<h�d<*p]<N*V<W�N<ͤG<�e@<�)9<T�1<޼*<��#<-a<�:<!<��<U��;ͻ�;���;��;Y��;�;"�;�k�;~ɐ;�;�;_�k;��P;�.6;>�;f�;�.�:���:��P:~��9���7�l���c?�G���C���j��Y�B~'�i�>���U��.l�!F���Q���:��������`$��s����˻��ջ=�߻B�黁M�~����%�����c����Db�j���#�n"�K�&�x�*��.�Q3��7�};���>���B��F�%}J�r=N���Q�f�U��AY���\��j`���c��pg���j�;Wn��q� u�zx���{�Y�u1��q҂��p��~�������<���ъ�Ld�����惏���|���m&��Ѯ���5������<@���Û�-F���Ǟ�WH��Jȡ�pG�� Ƥ�D�������>��`����7�� ���U0��h���o(������� ��B������ ���j��2�������  �  �yN="�M=��L=k9L=gxK=�J=��I=t2I=_oH=��G=H�F=A"F=u\E=�D=|�C=?C==B=�rA=ϧ@=��?=V?=�?>=5p==I�<=�;=c�:=A$:=�M9=�u8=��7=-�6=��5=�5=�"4=�?3=�Z2=Ss1=ى0=�/=�.=M�-=�,=O�+=��*=h�)="�(=��'=��&=�%=B�$=,�#=��"=��!=�~ =�b=�B=�=��=�=G�=bg=[/=�=��=�m=�$=[�=��=k/=��=v=�
=C�=c?=7�=�Z=6�=ye=P��<���<��<Ô�<�s�<�K�<�<w��<)��<d�<��<���<Gr�<��<۳�<wL�<��<�n�<���<L~�<���<*}�<���<m�<�߯<�O�<���<'�<��<���<�X�<���<��<!z�<؋<)5�<}��<Y�<��z<�Hs<��k<b�d<p]<b*V<e�N<ĤG<�e@<�)9<R�1<ϼ*<��#<,a<�:<'<z�<���;���;U��;Ѳ�;a��;;�;�!�;�k�;�ɐ;�;�;�k;��P;�.6;��;��;S.�::��P:���9���7�j��Xc?�r�������.��E�o~'�ӧ>�p�U�*/l��E���Q���:��� ������{$��i����˻��ջ0�߻T�黧M�@����%�����c����Bb�q���#�n"�P�&���*��.�[3��7�x;���>���B��F�3}J�q=N�v�Q�m�U��AY���\��j`���c��pg���j�-Wn��q� u�#zx���{�M�t1��z҂��p��x��¥���<���ъ�Ld����샏���z���c&��ٮ���5������>@���Û�3F���Ǟ�gH��Jȡ�rG��Ƥ��C�������>��`����7��'���P0��\���w(������� ��F����������b��7�������  �  �yN=+�M=��L=c9L=cxK=�J=��I=q2I=^oH=��G=K�F=?"F=o\E=�D=|�C=DC==B=�rA=ϧ@=��?=V?=�?>==p==G�<=��;=Z�:=G$:=�M9={u8=��7=*�6=��5=�5=�"4=�?3=�Z2=Xs1=։0=�/=�.=O�-=�,=L�+=��*=d�)=�(=��'=��&=�%==�$=)�#=��"=��!=�~ =�b=�B=�=��=�=J�=]g=W/=�=��=�m=�$=T�=��=v/=��=v=�
=A�=f?=4�=�Z=7�=}e=R��<���<��<���<�s�<�K�<�<���<��<d�<��< ��<Fr�<��<ҳ�<tL�<	��<�n�<���<J~�<���<!}�<���<m�<�߯<�O�<���<'�<
��<���<�X�<���<�<z�<؋<(5�<|��<Y�<��z<�Hs<��k<��d<p]<d*V<f�N<��G<�e@<�)9<u�1<ּ*<��#<a<�:<D<o�<z��;���;g��;���;.��;G�;�!�;l�;@ɐ;�;�;�k;��P;�.6;��;�;�-�:+��:{�P:��9(�77n��bb?������������V�$~'�ħ>��U�\/l��E���Q���:��� �����$������7�˻��ջ�߻G���M�Z���&�����c����Db�s���#�5n"�G�&���*��.�j3��7�h;��>���B���F�	}J�v=N���Q�d�U��AY���\��j`���c��pg���j�*Wn�)�q��u�0zx���{�e�n1��j҂��p�����ǥ���<���ъ�Md���������������\&��ܮ���5������F@���Û�:F���Ǟ�mH��?ȡ�sG��
Ƥ�
D�������>��g����7��(���P0��[���{(������� ��6����������b��<�������  �  �yN=#�M=��L=g9L=lxK=�J=��I=u2I=[oH=��G=J�F=?"F=q\E=��D=y�C=<C==B=�rA=Ч@=��?=U?=�?>=2p==I�<=�;=^�:=G$:=�M9=~u8=��7=-�6=��5=�5=�"4=�?3=�Z2=Us1=߉0=�/=�.=S�-=�,=M�+=��*=g�)=�(=��'=��&=�%=B�$=&�#=��"=��!=�~ =�b=�B=�=��=�=G�=`g=U/=�=��=�m=�$=[�=��=r/=��=v=�
=F�=e?==�=�Z=8�=~e=T��<���<��<Ɣ�<�s�<�K�<�<���<#��<d�<��<���<Mr�<��<ѳ�<vL�<��<�n�<���<G~�<���<#}�<���<m�<�߯<�O�<���<'�<���<���<�X�<���<��<z�<؋<15�<z��<Y�<Ƒz<�Hs<��k<x�d<5p]<h*V<]�N<ɤG<�e@<�)9<V�1<ܼ*<��#<@a<�:<$<��<[��;���;d��;���;:��;	�;�!�;�k�;Uɐ;�;�;�k;��P;�.6;��;S�;*.�:O��:b�P:���9���7�l��b?�������������~'���>�O�U��.l��E���Q���:��� �����P$��u����˻��ջ_�߻[�黥M�t���&�����c����Mb�v���#�(n"�R�&���*��.�]3��7��;���>���B��F�}J�u=N�u�Q�S�U��AY���\��j`���c��pg���j�&Wn��q�	 u�zx���{�S�s1��n҂��p��r�������<���ъ�Kd��
����	������h&��߮���5������C@���Û�2F���Ǟ�aH��Kȡ�G���Ť� D�������>��c����7�����R0��\���k(������� ��;������󖹼g��5�������  �  �yN=!�M=��L=f9L=hxK=�J=��I=s2I=XoH=��G=F�F=;"F=s\E=�D=��C=:C==B=�rA=ͧ@=��?=P?=�?>=3p==I�<=�;=_�:=G$:=�M9=�u8=��7=0�6=��5=�5=�"4=�?3=�Z2=Qs1=މ0=�/=�.=M�-=�,=T�+=��*=k�)=�(=��'=��&=�%=?�$=&�#=��"=��!=�~ =�b=�B=�=��=�=A�=cg=V/=�=��=�m=�$=X�=��=p/=��=v=�
=I�=f?==�=�Z=;�=|e=P��<���<��<͔�<�s�<�K�<�<���<&��<d�<��<���<Nr�<��<׳�<tL�<���<�n�<���<V~�<���<#}�<���<�l�<�߯<�O�<���<'�<	��<���<�X�<���<��<.z�<؋</5�<���<^�<z<�Hs<��k<^�d<2p]<r*V<u�N<ФG<�e@<�)9<N�1<�*<��#<1a<�:<&<v�<C��;û�;@��;���;G��;�;"�;�k�;tɐ;�;�;�k;��P;6.6;��;c�;6.�:���:��P:���9
��7:i���c?�0���e������>�Y~'�~�>���U��.l��E���Q���:��� ��֣��b$��V����˻��ջB�߻_�黾M�r����%����c����Cb�g���#�n"�n�&���*��.�n3��7��;���>���B�ݱF�#}J�_=N�o�Q�p�U��AY���\��j`���c��pg���j�0Wn��q��u�zx���{�;�q1��p҂��p��{��¥���<���ъ�Wd�����������~���m&��Ю���5������I@���Û�0F���Ǟ�hH��Jȡ�tG�� Ƥ�D��y����>��S����7��!���G0��V���n(������� ��H�������[��1�������  �  �yN=$�M=��L=f9L=gxK=�J=��I=p2I=]oH=��G=L�F=@"F=o\E=ܕD=x�C=7C==B=�rA=Χ@=��?=T?=�?>=9p==F�<=�;=]�:=G$:=�M9=u8=��7=.�6=��5=�5=�"4=�?3=�Z2=\s1=ى0=�/=�.=S�-= �,=N�+=��*=c�)=�(=��'=��&=�%=@�$='�#=��"=��!=�~ =�b=�B=�=��=�=G�=]g=V/=�=��=�m=�$=Y�=��=s/=��=v=�
=F�=f?=8�=�Z=>�=�e=b��<���<��<ǔ�<�s�<�K�<�<���<��<d�<��<���<Gr�<��<г�<rL�<	��<�n�<���<A~�<���<}�<���<	m�<�߯<�O�<���<'�<
��<���<�X�<���<��<z�<؋<15�<���<Z�<őz<�Hs<��k<��d<;p]<b*V<q�N<ͤG<�e@<�)9<[�1<޼*<��#</a<�:</<i�<k��;y��;m��;���;'��;��;�!�;�k�;Dɐ;�;�;��k;y�P;k.6;��;;�-�:���:��P:��9���7�l���b?�����<���������}'�[�>��U�(/l��E���Q���:��� �����M$�������˻��ջ�߻g�黹M�m���&�����c����]b�����#�+n"�S�&���*��.�b3��7�i;��>���B���F�}J�t=N�r�Q�V�U��AY���\��j`���c��pg���j�Wn�$�q��u�zx���{�P�v1��l҂��p��{��˥���<���ъ�Pd�����򃏼������s&��宕��5������D@���Û�CF���Ǟ�oH��Iȡ�sG��Ƥ�D�������>��a����7�����L0��[���l(������� ��4����������]��3�������  �  �yN=+�M=��L=i9L=jxK=�J=��I=n2I=aoH=��G=L�F=7"F=p\E=�D=y�C=AC==B=�rA=ͧ@=��?=[?=�?>=6p==A�<=	�;=\�:=G$:=�M9=}u8=��7=)�6=��5=�5=�"4=�?3=�Z2=Xs1=ډ0=!�/=�.=R�-=!�,=M�+=��*=`�)=&�(=��'=��&=�%=D�$='�#=��"=��!=�~ =�b=�B=�=��=�=H�=[g=V/=�=��=�m=�$=a�=��=y/=��=v=�
=D�=o?=9�=�Z=6�=~e=]��<���<)��<���<�s�<�K�<�<���<��<&d�<��<���<?r�<��<˳�<oL�<��<�n�<���<G~�<���<'}�<���<m�<�߯<�O�<���<'�<���<���<�X�<���<�<z�<"؋<)5�<���<f�<��z<�Hs<��k<��d<4p]<|*V<��N<��G<�e@<�)9<u�1<Լ*<��#<:a<�:<-<c�<���;i��;j��;z��;3��;(�;�!�;�k�;1ɐ;�;�;�k;P�P;�.6;N�;��;"-�:f��:��P:���9�7Am���a?�+���?������#~'��>�#�U� /l��E���Q���:��� �����$������ջ˻��ջG�߻j�黚M�h��� &���� d����Kb�w���#�Kn"�R�&���*��.�J3��7�z;��>���B��F�}J�t=N�v�Q�S�U��AY�u�\��j`���c��pg���j�Wn��q��u�4zx���{�V�o1��h҂��p��k��ӥ���<���ъ�@d���������������^&��߮���5������W@���Û�FF���Ǟ�nH��Hȡ�G�� Ƥ��C�������>��d����7��'���G0��O���o(������� ��7������ꖹ�U��>�������  �  �yN=(�M=��L=c9L=hxK=�J=��I=o2I=YoH=��G=L�F=8"F=p\E=ەD=y�C=6C==B=�rA=ҧ@=��?=S?=�?>=9p==I�<=�;=Z�:=D$:=�M9=�u8=��7=-�6=��5=�5=�"4=�?3=�Z2=[s1=މ0=�/=�.=P�-=$�,=R�+=��*=b�)=�(=��'=��&=�%=?�$= �#=��"=��!=�~ =�b=�B=�=��=�=E�=bg=O/=�=��=�m=�$=[�=��=t/=��=v=�
=F�=g?=<�=�Z=C�=�e=]��<���<��<ǔ�<�s�<�K�<�<���<��<d�<��<���<Dr�<��<Ƴ�<{L�<���<�n�<���<B~�<���<}�<���<	m�<�߯<�O�<���<'�<��<���<�X�<���<�<)z�<$؋<+5�<���<[�<őz<�Hs<��k<��d<7p]<l*V<v�N<ƤG<�e@<�)9<l�1<Ӽ*<��#<2a<�:<5<g�<J��;���;n��;���;,��;��;�!�;�k�;Uɐ;�;�;+�k;M�P;[.6;s�;��;1.�:ʘ�:8�P:���9��7�j��b?�����/���S�����}'�%�>���U��.l��E���Q���:��� ��룬�=$�������˻��ջ�߻_���M����&�����c����jb�����#�.n"�]�&���*�5�.�h3��7�i;���>���B��F�}J�d=N�f�Q�^�U��AY���\��j`���c��pg���j�Wn��q��u� zx���{�A�k1��s҂��p��v��å���<���ъ�Pd�����ꃏ�������v&��䮕��5������R@���Û�<F���Ǟ�pH��Dȡ�nG��Ƥ�
D�������>��W����7��%���I0��Z���l(��~���� ��/������򖹼[��7�������  �  �vN=��M=��L=�4L=GsK=E�J=��I=�+I=hH=ţG=��F=,F=�RE=��D=��C=��B=�0B=�eA=.�@=L�?=J�>=0>=�_==�<=ߺ;=v�:=�:=99=`8=R�7=��6=��5=��4=�4=�$3=�>2=mV1=l0=7/=�.=k�-=>�,=s�+=ֹ*=��)=1�(=�'=��&=#�%=q�$=f�#=��"=�j!=�Q =f4=�=��=j�=
�=�i=35=��=�=/=:=��=E�={Q=P�=�=,B="�	=�w=^=��=�(=Ű=�4=)i�<a�<-Q�<�9�<��<|��<
��<���<�W�<��<���<��<�+�<���<Ur�<��<��<l5�<��<�J�<�ν<O�<�˶<�D�<V��<-�<ܜ�<�	�<�t�<]ݝ<D�<䨖<�<n�<�΋<�.�<䍄<p�<��z<�Qs<�l<��d<J�]<�IV<�O<��G<ؕ@<�_9<�,2<��*<�#<�<I�<q<\<<M <���;7��;���;/��;z�;g'�;k{�;��;7`�;��m;q5S;L�8;�b;B;ĩ�:t7�:Rf\:�p�9�b�8�堹��2�84���y���@�����&$�MG;�)&R���h���ϕ���}��C���媻�f��IĿ�� ʻRԻL޻^�����0���Q���������=����Aa�"�!�.�%�� *�eE.��\2��f6��d:�yV>�f<B��F��I���M��dQ�U�F�X��X\�~�_�xc��f�vj�=�m��Tq���t�|x�o{���~����O���IH���兼����Q�������C��֍�yf�����ˁ��*��і��C��C���,��ఛ�u4��'����8�����J:��빤��8��w����5��_���1��C���X+�����%���������W���������\��:�������  �  �vN=��M=��L=�4L=OsK=L�J=��I=�+I=
hH=ţG=��F=+F=�RE=��D=��C=��B=�0B=fA=6�@=L�?=F�>=0>=�_==��<=�;=n�:=�:=99=`8=\�7=��6=��5=��4=�4=�$3=�>2=sV1=l0=8/=�.=o�-==�,=e�+=Թ*=w�)=3�(=��'=��&=)�%=n�$=e�#=��"=k!=�Q =h4=�=��=n�=�=�i=65=��=�=2=(:=��=J�=pQ=L�=ݠ=(B=(�	=�w=_=��=�(=̰=�4=,i�<a�<*Q�<�9�<��<j��<���<���<�W�<��<���<��<�+�<���<Vr�<��<��<b5�<'��<�J�<�ν<O�<�˶<�D�<U��<�,�<Ӝ�<
�<�t�<kݝ<�C�<Ѩ�<�<n�<�΋<�.�<ԍ�<s�<��z< Rs<�l<��d<?�]<�IV<�O<v�G<��@<�_9<�,2<��*<��#</�<e�<7q<�[<3M <���;���;���;��;��;"'�;�{�;��;_`�;4�m;|5S;�8;�b;�B;d��:�8�:Zd\:�l�9�T�8S령N�2�)5��Tz���@����P&$��F;��%R���h���*����}��C��
檻�f���Ŀ�u ʻԻ�޻4��$���0���Q�f������Y����2a�4�!�
�%�� *�gE.��\2��f6��d:�fV>�R<B��F�&�I���M��dQ��U�q�X��X\���_��wc���f��uj�6�m�Uq�ǹt��x��n{��~����^���\H���兼����=�������C��֍�jf�����ԁ����㖕�E��F���,��̰��w4��,����8��󹡼=:��ݹ���8�������5��{����0��C���h+��|����%���������M����������h��?�������  �  �vN=��M=��L=�4L=MsK=A�J=��I=�+I=hH=��G=��F=)F=�RE=��D=��C=��B=�0B=fA=3�@=J�?=J�>=0>=�_==�<=�;=m�:=�:=99=`8=e�7=�6=��5=��4=�4=�$3=�>2=wV1=�k0=A/=�.=u�-=@�,=f�+=�*=v�)=7�(=�'=��&=!�%=k�$=g�#=��"=k!=�Q =m4=�=��=u�= �=�i=/5=��=�=+= :=��=O�=oQ=[�=�=)B=0�	=�w=i=��=�(=°=�4=-i�<a�<6Q�<�9�<��<e��<
��<���<�W�<��<���<��<�+�<���<Sr�<��<���<S5�<8��<�J�<�ν<O�<�˶<�D�<J��<-�<͜�<
�<�t�<fݝ<�C�<Ө�<-�<�m�<�΋<�.�<э�<~�<��z<Rs<�l<��d<;�]<JV<�O<q�G<�@<}_9<�,2<��*<�#<(�<8�<.q<�[<MM <���;���;���;��;��;%'�;�{�;��;p`�; �m;[5S;O�8;Hb;eB;���:�8�:d\:q�9�k�8>�7�2��5���y���@�����&$��G;��%R�(�h�V�F����}���B�� 檻f���Ŀ�Z ʻ]ԻF޻p��7���0��R�X������A����a�N�!� �%�!*�dE.��\2�g6��d:��V>�?<B��F���I���M��dQ��U���X�mX\���_��wc��f�vj�5�m�Uq���t��x��n{�'�~����H���^H���兼����F�������C��!֍�uf������䁒���▕�3��E���&,��Ȱ���4�� ����8������S:��㹤��8�������5�������0��@���k+��q����%���������L��� ������f��B�������  �  �vN=��M=��L=�4L=KsK=J�J=��I=�+I=hH=ģG=��F=.F=�RE=��D=��C=��B=�0B=	fA=0�@=M�?=J�>=0>=�_==�<=�;=p�:=�:=99=`8=\�7=�6=��5=��4=�4=�$3=�>2=zV1=�k0=</=�.=o�-=<�,=h�+=׹*=v�)=6�(=�'=��&=(�%=m�$=i�#=�"=
k!=�Q =e4=�=��=m�=�=�i=35=��=�=1=(:=��=L�=pQ=O�=�=(B=)�	=�w=d=��=�(=Ű=�4=3i�<a�<3Q�<�9�<��<j��<��<���<�W�<��<���<��<�+�<���<Yr�<��<���<\5�<'��<�J�<�ν<O�<�˶<�D�<S��<-�<Ҝ�<
�<�t�<gݝ<�C�<Ϩ�<�<n�<�΋<�.�<؍�<p�<��z<Rs<�l<�d<<�]<�IV<�O<p�G<��@<�_9<�,2<��*<
�#< �<\�<Gq<�[<NM <���;u��;���;��;��;5'�;�{�;��;�`�;��m;�5S;W�8;�b;�B;$��:�8�:�d\:Wm�9M`�8�꠹.�2�h5���y��TA����J&$�zG;�P%R�H�h���.����}��C���媻uf���Ŀ�c ʻ8Ի�޻5��%���0���Q�\������K����6a�4�!���%�� *�\E.��\2��f6��d:�qV>�I<B��F��I���M��dQ��U�t�X�X\���_��wc� �f��uj�(�m�Uq���t��x��n{��~����[���\H���兼����9�������C��֍�wf������ځ��������=��M���,��Ͱ��y4������8��칡�=:��⹤��8�������5��x����0��C���e+��~����%���������E��� �����`��C�������  �  �vN=��M=��L=�4L=HsK=J�J=��I=�+I=
hH=ɣG=��F=,F=�RE=��D=��C=��B=�0B=fA=2�@=P�?=F�>=0>=�_==�<=�;=t�:=�:=99=`8=Y�7=��6=��5=��4=�4=�$3=�>2=rV1=�k0=:/=�.=n�-=>�,=m�+=Թ*=�)=/�(=�'=��&=%�%=m�$=c�#=��"=k!=�Q =f4=�=��=m�=�=�i=55=��=�=/=!:=��=E�=xQ=M�=�=*B=&�	=�w=a=��=�(=ð=�4=)i�<a�<+Q�<�9�<��<s��<��<���<�W�<��<���<��<�+�<���<[r�<��<��<e5�<*��<�J�<�ν<	O�<�˶<�D�<^��<�,�<Ҝ�<
�<�t�<^ݝ<�C�<ᨖ<�<n�<�΋<�.�<ҍ�<q�<��z<�Qs<�l<��d<@�]<�IV<�O<o�G<�@<�_9<�,2<��*<�#<�<^�<!q<�[<3M <͊�;`��;���;��;��;i'�;�{�;��;_`�;��m;�5S;�8;�b;3B;)��:�7�:�e\:�n�9b]�8*蠹��2�.5��1z���@�����&$��G;��%R��h���*����}��C���媻�f��_Ŀ�� ʻBԻ"޻N��$���0���Q�x������8����5a�*�!��%�� *�gE.��\2��f6��d:�rV>�e<B��F� �I���M��dQ�U�r�X��X\���_�xc��f��uj�:�m�Uq�ùt��x�o{�
�~����Y���MH���兼����L�������C��֍�rf�����ҁ����Җ��8��I���,��ְ��n4��-����8������@:��깤��8��z����5��j����0��F���j+��}����%���������S���������i��C�������  �  �vN=��M=��L=�4L=OsK=I�J=��I=�+I=hH=ãG=��F=/F=�RE=��D=��C=��B=�0B=fA=3�@=K�?=J�>=0>=�_==�<=�;=k�:=�:=99=`8=[�7=��6=��5=��4=�4=�$3=�>2=rV1=�k0=:/=�.=r�-=<�,=h�+=׹*=v�)=0�(=��'=��&='�%=v�$=d�#=�"=
k!=�Q =i4=�=��=o�=�=�i=25=��=�=3= :=��=F�=oQ=N�=�=%B=*�	=�w=`=��=�(=ǰ=�4=%i�<a�<)Q�<�9�<��<b��<��<���<�W�<��<���<��<�+�<���<Sr�<��<���<a5�<.��<�J�<�ν<O�<�˶<�D�<Q��<�,�<木<
�<�t�<mݝ<�C�<Ѩ�<�<n�<�΋<�.�<̍�<w�<��z<�Qs<�l<��d<0�]<JV<�O<z�G<��@<�_9<�,2<��*<��#<0�<W�<!q<$\<?M <���;|��;���;,��;��;"'�;�{�;��;�`�;�m;v5S;\�8;c;5B;1��:�8�:�c\:�m�9@e�8�젹a�2�)5��<z���@�,��o&$�DG;��%R�;�h���G����}��C���媻tf���Ŀ�� ʻԻ1޻=������0���Q�[������D����,a�1�!���%� !*�hE.��\2��f6��d:�`V>�_<B��F��I���M��dQ��U���X��X\���_��wc���f��uj�A�m�Uq�ƹt��x��n{�*�~����[���`H���兼����K�������C�� ֍�rf������Ձ����▕�6��B���,��Ͱ��{4��*����8������E:��۹��9�������5��|����0��@���p+��x����%���������P���������m��>�������  �  �vN=��M=��L=�4L=OsK=H�J=��I=�+I=hH=ţG=��F=1F=�RE=��D=��C=��B=�0B=fA=5�@=N�?=I�>=0>=�_==�<=�;=s�:=�:=99=	`8=Z�7=�6=��5=��4=�4=�$3=�>2=tV1=�k0=@/=�.=n�-=;�,=h�+=ٹ*=x�)=7�(=�'=��&=(�%=o�$=h�#=�"=k!=�Q =j4=�=��=r�=�=�i=25=��=�=2=$:=��=M�=qQ=P�=�=&B=(�	=�w=f=��=�(=ð=�4=%i�<a�<5Q�<�9�<��<e��<��<���<�W�<��<���<��<�+�<���<Yr�<��<��<Y5�<4��<�J�<�ν<O�<�˶<�D�<U��<-�<Ӝ�<
�<�t�<jݝ<D�<Ψ�<�<n�<�΋<�.�<ԍ�<z�<q�z<Rs<�l<��d<"�]<JV<�O<g�G<�@<�_9<�,2<��*<�#<-�<V�<6q<�[<AM <���;���;ȗ�;��;��;>'�;�{�;��;�`�;+�m;�5S;F�8;�b;�B;���:�8�:�e\:�m�9�g�8�령��2��5��xy��A�"��i&$��G;��%R�t�h�n�B����}��C���媻df���Ŀ�Q ʻ5Ի޻4�����0���Q�F������8����a�=�!���%�� *�WE.��\2��f6��d:�tV>�D<B��F��I���M��dQ��U��X�uX\���_��wc��f��uj�@�m�Uq���t��x��n{�%�~����Z���VH���兼����B�������C��֍�rf������݁����ܖ��/��I���,��°��w4��&����8��򹡼B:��߹���8�������5��|����0��H���h+��t����%���������L���������b��G�������  �  �vN=��M=��L=�4L=EsK=K�J=��I=�+I=hH=ʣG=��F=0F=�RE=��D=��C=��B=�0B=
fA=2�@=R�?=J�>=0>=�_==�<=�;=u�:=�:=99=`8=X�7=�6=��5=��4=�4=�$3=�>2=pV1=�k0=;/=�.=k�-=?�,=m�+=չ*={�)=1�(=�'=��&='�%=m�$=i�#=��"=k!=�Q =j4=�=��=q�=�=�i=25=��=�=0=":=��=F�=vQ=L�=�=+B=$�	=�w=`=��=�(=��=�4=&i�<	a�<*Q�<�9�<��<t��<���<���<�W�<��<���<��<�+�<���<ar�<��<���<a5�<1��<�J�<�ν<	O�<�˶<�D�<^��<-�<М�<
�<�t�<Yݝ<D�<Ө�<�<n�<�΋<�.�<ύ�<q�<��z<�Qs<�l<��d<9�]<�IV<�O<\�G<�@<�_9<�,2<��*<�#<�<_�<4q<�[<EM <Պ�;u��;Ɨ�;��;��;g'�;�{�;��;�`�;��m;�5S;Y�8;�b;|B;��:�7�:7f\:�l�9i^�8`砹<�2��5��(z��A�����&$��G;��%R�7�h���?����}���B���媻�f��|Ŀ�� ʻUԻ޻@��'��0���Q�`��ݔ���-����"a�,�!��%�� *�RE.��\2��f6��d:��V>�^<B��F�!�I���M��dQ�U���X��X\���_�	xc��f�vj�>�m�Uq�ùt��x�o{��~����_���OH���兼����F�������C��֍�tf������Ձ����Ӗ��2��H���,��ΰ��o4��#����8��󹡼@:��﹤��8�������5��k����0��M���m+��~����%���������R��� �����k��L�������  �  �vN=��M=��L=�4L=KsK=O�J=��I=�+I=hH=ȣG=��F=/F=�RE=��D=��C=��B=�0B=fA=5�@=N�?=I�>=0>=�_==��<=�;=m�:=�:=99=`8=V�7=��6=��5=��4=�4=�$3=�>2=nV1=�k0=4/=�.=n�-=9�,=f�+=Թ*=x�)=/�(=��'=��&='�%=t�$=d�#=��"=	k!=�Q =j4=�=��=q�=
�=�i=55=��=�=2=!:=��=D�=rQ=K�=ߠ=$B=%�	=�w=Y=��=�(=Ű=�4=i�<
a�<Q�<�9�<��<b��<���<���<�W�<��<���<��<�+�<���<Xr�<��<���<f5�<0��<�J�<�ν<O�<�˶<�D�<\��<-�<䜨<
�<�t�<iݝ<�C�<Ө�<�<n�<�΋<�.�<̍�<i�<��z<�Qs<�l<��d<3�]<�IV<�O<t�G<�@<�_9<�,2<��*<��#<�<o�<$q<!\<?M <Ŋ�;���;���;8��;��;V'�;�{�;��;�`�;4�m;�5S;L�8;.c;EB;%��:
8�:wd\:�m�9�]�85젹��2�5���z��A�3���&$�8G;�&R��h��9����}��)C���媻�f���Ŀ�� ʻԻ޻;�����0���Q�\��ؔ���7����%a� �!���%�� *�eE.��\2��f6��d:�XV>�e<B��F�#�I���M��dQ�	U�w�X��X\���_�xc���f��uj�M�m�Uq�ܹt��x�o{�(�~����[���[H���兼����L�������C��֍�lf������Ё����ږ��5��@���,��̰��p4��'����8������<:��߹���8�������5��z���1��C���p+�������%���������W�����
���p��@�������  �  �vN=��M=��L=�4L=KsK=I�J=��I=�+I=hH=ǣG=��F=,F=�RE=��D=��C=��B=�0B=fA=7�@=P�?=J�>=0>=�_==�<=�;=q�:=�:=99=`8=]�7=�6=��5=��4=�4=�$3=�>2=mV1=�k0=;/=�.=n�-=<�,=f�+=ݹ*=x�)=6�(=�'=��&='�%=p�$=i�#=��"=k!=�Q =o4=�=��=x�=�=�i=55=��=�=1=":=��=K�=qQ=S�=�=%B=&�	=�w=`=��=�(=��=�4=i�<a�<(Q�<�9�<��<a��<��<���<�W�<��<���<��<�+�<���<[r�<��<���<`5�<A��<�J�<�ν<O�<�˶<�D�<Y��<-�<؜�<
�<�t�<cݝ<�C�<Ө�<%�<n�<�΋<�.�<ʍ�<t�<x�z<�Qs<�l<��d<'�]<�IV<�O<_�G<��@<�_9<�,2<��*<
�#<�<W�<)q<\<IM <Ê�;���;���;9��;��;V'�;|�;��;�`�;[�m;�5S;a�8;�b;tB;��:�8�:e\:�o�9m�8>젹��2��5��(z��A�O���&$��G;�&R�X�h���M����}��C���媻@f���Ŀ�[ ʻJԻ޻<��
��0���Q�M������0����	a�5�!���%�� *�WE.��\2��f6��d:�{V>�H<B��F��I���M��dQ�U��X��X\���_�xc��f�vj�Q�m�Uq�Ĺt��x��n{�*�~����R���WH���兼����F�������C��֍�lf������ց����ٖ��*��<���,��ð��s4��!����8������C:��湤��8�������5��|����0��L���r+��z����%���������[���
�����m��K�������  �  �vN=��M=��L=�4L=IsK=N�J=��I=�+I=hH=ƣG=��F=3F=�RE=��D=��C=��B=�0B=fA=4�@=R�?=P�>=0>=�_==�<=�;=p�:=|:=99=`8=\�7=�6=��5=��4=�4=�$3=�>2=uV1=�k0=8/=�.=k�-=;�,=b�+=׹*=p�)=9�(=�'=��&=)�%=n�$=q�#=�"=k!=�Q =l4=�=��=u�=�=�i=25=��=�=1=-:=��=N�=iQ=L�=۠=#B=$�	=�w=_=��=�(=��=�4=*i�<�`�<+Q�<�9�<��<\��<���<���<�W�<��<���<��<�+�<���<er�<��<��<d5�<:��<�J�<�ν<O�<�˶<�D�<T��<-�<Μ�<
�<�t�<_ݝ<D�<���<�<�m�<�΋<�.�<ύ�<l�<q�z<Rs<�l<��d<)�]<�IV<�O<U�G<��@<z_9<�,2<��*<�#<�<k�<Nq<�[<gM <���;���;ޗ�;/��;��;;'�;�{�;��;�`�;#�m;�5S;��8;�b;1C;2��:�8�:e\:j�9�_�8���2�06���y���A�����&$��G;��%R���h���O����}��C��檻qf���Ŀ�? ʻOԻ�޻)����~0���Q�C��ݔ���A����a�*�!���%�� *�;E.��\2��f6��d:�}V>�<<B��F��I���M��dQ�U���X��X\���_��wc��f� vj�4�m�-Uq���t��x��n{�3�~����g���^H���兼����.�������C��֍�rf������ҁ����ߖ��3��B���,��Ű��x4������8��빡�5:��깤��8�������5�������0��P���m+�������%���������M��������i��P�������  �  �vN=��M=��L=�4L=IsK=I�J=��I=�+I=hH=ɣG=��F=0F=�RE=��D=��C=��B=�0B=fA=6�@=P�?=J�>=0>=�_==�<=�;=t�:=�:=99=`8=W�7=�6=��5=��4=�4=�$3=�>2=mV1=�k0=6/=�.=l�-=:�,=g�+=ܹ*={�)=4�(=�'=��&=!�%=o�$=h�#=��"=k!=�Q =k4=�=��=r�=�=�i=55=��=�=+=:=��=I�=tQ=R�=�=$B=$�	=�w=\=��=�(=��=�4=!i�<a�<%Q�<�9�<��<b��<��<���<�W�<��<���<��<�+�<���<Zr�<��<���<i5�<1��<�J�<�ν<O�<�˶<�D�<]��<-�<ל�<�	�<�t�<`ݝ<D�<ר�<�<n�<�΋<�.�<ԍ�<i�<��z<�Qs<�l<��d<3�]<�IV<�O<f�G<�@<�_9<�,2<��*<�#<�<Y�<q<\<HM <ӊ�;���;ȗ�;5��;��;�'�;�{�;��;�`�;I�m;�5S;e�8;�b;6B;,��:e8�:f\:wo�9Oh�8�령)�2��5��#z��MA���'$��G;�&R�)�h��� ����}��"C���媻Lf��xĿ�k ʻGԻ,޻m�����0���Q�`��Ք�����z�a��!��%�� *�ZE.��\2� g6��d:�{V>�P<B��F��I���M��dQ�U�r�X��X\���_�xc��f�vj�E�m�Uq�ɹt��x�o{�(�~����S���QH���兼����N�������C��֍�kf������́����ǖ��-��A���,��Ͱ��o4��!����8�����D:��鹤��8�������5��|���1��K���h+�������%���������_�����
���g��G�������  �  �vN=��M=��L=�4L=NsK=Q�J=��I=�+I=hH=ΣG=��F=0F=�RE=��D=��C=��B=�0B=fA=?�@=N�?=F�>=$0>=�_==��<=�;=m�:=�:=99=`8=Z�7=�6=��5=��4=�4=�$3=�>2=gV1=l0=./=�.=k�-=>�,=g�+=ѹ*=x�)=,�(=��'=��&=,�%=w�$=`�#=�"=	k!=�Q =i4=�=��=n�=�=�i=?5=��=�=8=$:=��=C�=pQ=H�=ߠ='B=#�	=�w=T=��=�(=Ű=�4=i�<
a�<Q�<�9�<��<h��<���<���<�W�<��<���<��<�+�<���<Sr�<��<��<r5�<%��<�J�<�ν<O�<�˶<�D�<k��<�,�<휨<
�<�t�<nݝ<�C�<̨�<�<n�<�΋<�.�<�<c�<��z<�Qs<�l<��d<?�]<�IV<mO<a�G<�@<�_9<�,2<��*<��#<(�<y�<&q<6\<$M <���;���;�;E��;��;�'�;�{�;�;�`�;��m;�5S;#�8;�c;CB;w��:�8�:|d\:#l�9�[�8�頹��2�]5��c{���@�	���&$�'G;�m&R���h�z�Q����}��C���媻�f���Ŀ�� ʻ�Ի�޻��М�1���Q�_��Ŕ���=����.a��!�	�%�� *�tE.��\2��f6��d:�QV>�i<B��F�/�I���M��dQ�U���X��X\���_�"xc���f�vj�I�m�Uq��t��x�o{��~����e���^H���兼����K�������C��֍�Uf������ā����Ж��9��?���,��İ��a4��5����8������3:��۹��9�������5��s����0��L���z+�������%���������d���������z��I�������  �  �vN=��M=��L=�4L=IsK=I�J=��I=�+I=hH=ɣG=��F=0F=�RE=��D=��C=��B=�0B=fA=6�@=P�?=J�>=0>=�_==�<=�;=t�:=�:=99=`8=W�7=�6=��5=��4=�4=�$3=�>2=mV1=�k0=6/=�.=l�-=:�,=g�+=ܹ*={�)=4�(=�'=��&=!�%=o�$=h�#=��"=k!=�Q =k4=�=��=r�=�=�i=55=��=�=+=:=��=I�=tQ=R�=�=$B=$�	=�w=\=��=�(=��=�4=!i�<a�<%Q�<�9�<��<b��<��<���<�W�<��<���<��<�+�<���<Zr�<��<���<i5�<1��<�J�<�ν<O�<�˶<�D�<]��<-�<ל�<�	�<�t�<`ݝ<D�<ר�<�<n�<�΋<�.�<ԍ�<i�<��z<�Qs<�l<��d<3�]<�IV<�O<f�G<�@<�_9<�,2<��*<�#<�<Y�<q<\<HM <ӊ�;���;ȗ�;5��;��;�'�;�{�;��;�`�;I�m;�5S;d�8;�b;6B;+��:d8�:f\:so�9?h�8�령+�2��5��$z��NA���'$��G;�&R�*�h��� ����}��"C���媻Mf��xĿ�k ʻGԻ-޻m�����0���Q�`��Ք�����z�a��!��%�� *�ZE.��\2� g6��d:�{V>�P<B��F��I���M��dQ�U�r�X��X\���_�xc��f�vj�E�m�Uq�ɹt��x�o{�(�~����S���QH���兼����N�������C��֍�kf������́����ǖ��-��A���,��Ͱ��o4��!����8�����D:��鹤��8�������5��|���1��K���h+�������%���������_�����
���g��G�������  �  �vN=��M=��L=�4L=IsK=N�J=��I=�+I=hH=ƣG=��F=3F=�RE=��D=��C=��B=�0B=fA=4�@=R�?=P�>=0>=�_==�<=�;=p�:=|:=99=`8=\�7=�6=��5=��4=�4=�$3=�>2=uV1=�k0=8/=�.=k�-=;�,=b�+=׹*=p�)=9�(=�'=��&=)�%=n�$=q�#=�"=k!=�Q =l4=�=��=u�=�=�i=25=��=�=1=-:=��=N�=iQ=L�=۠=#B=$�	=�w=_=��=�(=��=�4=*i�<�`�<+Q�<�9�<��<\��<���<���<�W�<��<���<��<�+�<���<er�<��<��<d5�<:��<�J�<�ν<O�<�˶<�D�<T��<-�<Μ�<
�<�t�<_ݝ<D�<���<�<�m�<�΋<�.�<ύ�<l�<q�z<Rs<�l<��d<)�]<�IV<�O<U�G<��@<z_9<�,2<��*<�#<�<k�<Nq<�[<gM <���;���;ޗ�;/��;��;;'�;�{�;��;�`�;#�m;�5S;��8;b;0C;1��:�8�:e\:j�9�_�8���2�26���y���A�����&$��G;��%R���h���O����}��C��檻qf���Ŀ�? ʻOԻ�޻)����~0���Q�C��ݔ���A����a�*�!���%�� *�;E.��\2��f6��d:�}V>�<<B��F��I���M��dQ�U���X��X\���_��wc��f� vj�4�m�-Uq���t��x��n{�3�~����g���^H���兼����.�������C��֍�rf������ҁ����ߖ��3��B���,��Ű��x4������8��빡�5:��깤��8�������5�������0��P���m+�������%���������M��������i��P�������  �  �vN=��M=��L=�4L=KsK=I�J=��I=�+I=hH=ǣG=��F=,F=�RE=��D=��C=��B=�0B=fA=7�@=P�?=J�>=0>=�_==�<=�;=q�:=�:=99=`8=]�7=�6=��5=��4=�4=�$3=�>2=mV1=�k0=;/=�.=n�-=<�,=f�+=ݹ*=x�)=6�(=�'=��&='�%=p�$=i�#=��"=k!=�Q =o4=�=��=x�=�=�i=55=��=�=1=":=��=K�=qQ=S�=�=%B=&�	=�w=`=��=�(=��=�4=i�<a�<(Q�<�9�<��<a��<��<���<�W�<��<���<��<�+�<���<[r�<��<���<`5�<A��<�J�<�ν<O�<�˶<�D�<Y��<-�<؜�<
�<�t�<cݝ<�C�<Ө�<%�<n�<�΋<�.�<ʍ�<t�<x�z<�Qs<�l<��d<'�]<�IV<�O<_�G<��@<�_9<�,2<��*<
�#<�<W�<)q<\<IM <Ê�;���;���;9��;��;V'�;|�;��;�`�;Z�m;�5S;`�8;�b;sB;��:�8�:ze\:�o�9�l�8H젹��2��5��+z��A�P���&$��G;�&R�Y�h���M����}��C���媻@f���Ŀ�\ ʻKԻ޻<����0���Q�M������1����	a�5�!���%�� *�WE.��\2��f6��d:�{V>�H<B��F��I���M��dQ�U��X��X\���_�xc��f�vj�Q�m�Uq�Ĺt��x��n{�*�~����R���WH���兼����F�������C��֍�lf������ց����ٖ��*��<���,��ð��s4��!����8������C:��湤��8�������5��|����0��L���r+��z����%���������[���
�����m��K�������  �  �vN=��M=��L=�4L=KsK=O�J=��I=�+I=hH=ȣG=��F=/F=�RE=��D=��C=��B=�0B=fA=5�@=N�?=I�>=0>=�_==��<=�;=m�:=�:=99=`8=V�7=��6=��5=��4=�4=�$3=�>2=nV1=�k0=4/=�.=n�-=9�,=f�+=Թ*=x�)=/�(=��'=��&='�%=t�$=d�#=��"=	k!=�Q =j4=�=��=q�=
�=�i=55=��=	�=2=!:=��=D�=rQ=K�=ߠ=$B=%�	=�w=Y=��=�(=Ű=�4=i�<
a�<Q�<�9�<��<b��<���<���<�W�<��<���<��<�+�<���<Xr�<��<���<f5�<0��<�J�<�ν<O�<�˶<�D�<\��<-�<䜨<
�<�t�<iݝ<�C�<Ө�<�<n�<�΋<�.�<̍�<i�<��z<�Qs<�l<��d<3�]<�IV<�O<t�G<�@<�_9<�,2<��*<��#< �<p�<$q<!\<?M <Ŋ�;���;���;8��;��;V'�;�{�;��;�`�;3�m;�5S;K�8;,c;CB;"��:8�:qd\:�m�9�]�8B젹��2�5���z��A�4���&$�9G;�	&R��h��9����}��*C���媻�f���Ŀ�� ʻ	Ի޻;�����0���Q�\��ؔ���7����%a� �!���%�� *�eE.��\2��f6��d:�XV>�e<B��F�#�I���M��dQ�	U�w�X��X\���_�xc���f��uj�M�m�Uq�ܹt��x�o{�(�~����[���[H���兼����L�������C��֍�lf������Ё����ږ��5��@���,��̰��p4��'����8������<:��߹���8�������5��z���1��C���p+�������%���������W�����
���p��@�������  �  �vN=��M=��L=�4L=EsK=K�J=��I=�+I=hH=ʣG=��F=0F=�RE=��D=��C=��B=�0B=
fA=2�@=R�?=J�>=0>=�_==�<=�;=u�:=�:=99=`8=X�7=�6=��5=��4=�4=�$3=�>2=pV1=�k0=;/=�.=k�-=?�,=m�+=չ*={�)=1�(=�'=��&='�%=m�$=i�#=��"=k!=�Q =j4=�=��=q�=�=�i=25=��=�=0=":=��=F�=vQ=L�=�=+B=$�	=�w=a=��=�(=��=�4=&i�<	a�<*Q�<�9�<��<t��<���<���<�W�<��<���<��<�+�<���<ar�<��<���<a5�<1��<�J�<�ν<	O�<�˶<�D�<^��<-�<М�<
�<�t�<Yݝ<D�<Ҩ�<�<n�<�΋<�.�<ύ�<p�<��z<�Qs<�l<��d<9�]<�IV<�O<\�G<�@<�_9<�,2<��*<�#<�<_�<4q<�[<EM <Պ�;u��;Ɨ�;��;��;g'�;�{�;��;�`�;��m;�5S;X�8;�b;zB;��:�7�:0f\:�l�90^�8n砹C�2��5��+z��A�����&$��G;��%R�9�h���@����}���B���媻�f��}Ŀ�� ʻVԻ޻@��(��0���Q�`��ݔ���-����"a�,�!��%�� *�RE.��\2��f6��d:��V>�^<B��F�!�I���M��dQ�U���X��X\���_�	xc��f�vj�>�m�Uq�ùt��x�o{��~����_���OH���兼����F�������C��֍�tf������Ձ����Ӗ��2��H���,��ΰ��o4��#����8��󹡼@:��﹤��8�������5��k����0��M���m+��~����%���������R��� �����k��L�������  �  �vN=��M=��L=�4L=OsK=H�J=��I=�+I=hH=ţG=��F=1F=�RE=��D=��C=��B=�0B=fA=5�@=N�?=I�>=0>=�_==�<=�;=s�:=�:=99=	`8=Z�7=�6=��5=��4=�4=�$3=�>2=tV1=�k0=@/=�.=n�-=;�,=h�+=ٹ*=x�)=7�(=�'=��&=(�%=o�$=h�#=�"=k!=�Q =j4=�=��=r�=�=�i=25=��=�=2=$:=��=M�=qQ=P�=�=&B=(�	=�w=f=��=�(=ð=�4=%i�<a�<5Q�<�9�<��<e��<��<���<�W�<��<���<��<�+�<���<Yr�<��<��<Y5�<4��<�J�<�ν<O�<�˶<�D�<U��<-�<Ӝ�<
�<�t�<jݝ<D�<Ψ�<�<n�<�΋<�.�<ԍ�<z�<q�z<Rs<�l<��d<"�]<JV<�O<g�G<�@<�_9<�,2<��*<�#<-�<V�<7q<�[<AM <���;���;ȗ�;��;��;>'�;�{�;��;�`�;*�m;�5S;E�8;�b;�B;��:�8�:�e\:�m�9�g�8�령��2��5��|y�� A�$��k&$��G;��%R�u�h�o�C����}��C���媻ef���Ŀ�R ʻ6Ի޻4�����0���Q�F������8����a�=�!���%�� *�WE.��\2��f6��d:�tV>�D<B��F��I���M��dQ��U��X�uX\���_��wc��f��uj�@�m�Uq���t��x��n{�%�~����Z���VH���兼����B�������C��֍�rf������݁����ܖ��/��I���,��°��w4��&����8��򹡼B:��߹���8�������5��|����0��H���h+��t����%���������L���������b��G�������  �  �vN=��M=��L=�4L=OsK=I�J=��I=�+I=hH=ãG=��F=/F=�RE=��D=��C=��B=�0B=fA=3�@=K�?=J�>=0>=�_==�<=�;=k�:=�:=99=`8=[�7=��6=��5=��4=�4=�$3=�>2=rV1=�k0=:/=�.=r�-=<�,=h�+=׹*=v�)=0�(=��'=��&='�%=v�$=d�#=�"=
k!=�Q =i4=�=��=o�=�=�i=25=��=�=3= :=��=F�=oQ=N�=�=&B=*�	=�w=`=��=�(=ǰ=�4=&i�<a�<)Q�<�9�<��<c��<��<���<�W�<��<���<��<�+�<���<Sr�<��<���<b5�<.��<�J�<�ν<O�<�˶<�D�<Q��<�,�<在<
�<�t�<mݝ<�C�<Ѩ�<�<n�<�΋<�.�<̍�<w�<��z<�Qs<�l<��d<0�]<JV<�O<z�G<��@<�_9<�,2<��*<��#<0�<W�<!q<$\<?M <���;|��;���;,��;��;"'�;�{�;��;�`�;�m;u5S;[�8;c;4B;-��:�8�:�c\:�m�9e�8�젹h�2�-5��?z���@�-��p&$�FG;��%R�<�h���H����}��C���媻uf���Ŀ�� ʻԻ1޻=�����0���Q�[������D����,a�1�!���%� !*�hE.��\2��f6��d:�`V>�_<B��F��I���M��dQ��U���X��X\���_��wc���f��uj�A�m�Uq�ƹt��x��n{�*�~����[���`H���兼����K�������C�� ֍�rf������Ձ����▕�6��B���,��Ͱ��{4��*����8������E:��۹��9�������5��|����0��@���p+��x����%���������P���������m��>�������  �  �vN=��M=��L=�4L=HsK=J�J=��I=�+I=
hH=ɣG=��F=,F=�RE=��D=��C=��B=�0B=fA=2�@=P�?=F�>=0>=�_==�<=�;=t�:=�:=99=`8=Y�7=��6=��5=��4=�4=�$3=�>2=rV1=�k0=:/=�.=n�-=>�,=m�+=Թ*=�)=/�(=�'=��&=%�%=m�$=c�#=��"=k!=�Q =f4=�=��=m�=�=�i=55=��=�=/=!:=��=E�=yQ=M�=�=*B=&�	=�w=a=��=�(=ð=�4=*i�<a�<+Q�<�9�<��<s��<��<���<�W�<��<���<��<�+�<���<[r�<��<��<e5�<*��<�J�<�ν<	O�<�˶<�D�<^��<�,�<Ҝ�<
�<�t�<^ݝ<�C�<ᨖ<�<n�<�΋<�.�<ҍ�<q�<��z<�Qs<�l<��d<@�]<�IV<�O<o�G<�@<�_9<�,2<��*<�#<�<^�<!q<�[<3M <͊�;a��;���;��;��;h'�;�{�;��;_`�;��m;�5S;�8;�b;2B;&��:�7�:�e\:xn�9/]�87蠹��2�15��4z���@�����&$��G;��%R��h���*����}��C���媻�f��_Ŀ�� ʻCԻ#޻O��$���0���Q�x������8����5a�*�!��%�� *�hE.��\2��f6��d:�rV>�e<B��F� �I���M��dQ�U�r�X��X\���_�xc��f��uj�:�m�Uq�ùt��x�o{�
�~����Y���MH���兼����L�������C��֍�rf�����ҁ����Җ��8��I���,��ְ��n4��-����8������@:��깤��8��z����5��j����0��F���j+��}����%���������S���������i��C�������  �  �vN=��M=��L=�4L=KsK=J�J=��I=�+I=hH=ģG=��F=.F=�RE=��D=��C=��B=�0B=	fA=0�@=M�?=J�>=0>=�_==�<=�;=p�:=�:=99=`8=\�7=�6=��5=��4=�4=�$3=�>2=zV1=�k0=</=�.=o�-=<�,=h�+=׹*=v�)=6�(=�'=��&=(�%=m�$=i�#=�"=
k!=�Q =e4=�=��=m�=�=�i=35=��=�=1=(:=��=L�=pQ=O�=�=(B=)�	=�w=d=��=�(=Ű=�4=3i�<a�<3Q�<�9�<��<k��<��<���<�W�<��<���<��<�+�<���<Yr�<��<���<\5�<'��<�J�<�ν<O�<�˶<�D�<S��<-�<Ҝ�<
�<�t�<fݝ<�C�<Ϩ�<�<n�<�΋<�.�<؍�<p�<��z<Rs<�l<�d<<�]<�IV<�O<p�G<��@<�_9<�,2<��*<
�#< �<\�<Gq<�[<NM <���;u��;���;��;��;5'�;�{�;��;�`�;��m;�5S;V�8;�b;�B;"��:�8�:�d\:Mm�9#`�8�꠹3�2�j5���y��WA����K&$�{G;�Q%R�I�h���.����}��C���媻uf���Ŀ�c ʻ9Ի�޻5��%���0���Q�]������K����6a�4�!���%�� *�\E.��\2��f6��d:�qV>�I<B��F��I���M��dQ��U�t�X��X\���_��wc� �f��uj�(�m�Uq���t��x��n{��~����[���\H���兼����9�������C��֍�wf������ځ��������=��M���,��Ͱ��y4������8��칡�=:��⹤��8�������5��x����0��C���e+��~����%���������E��� �����`��C�������  �  �vN=��M=��L=�4L=MsK=A�J=��I=�+I=hH=��G=��F=)F=�RE=��D=��C=��B=�0B=fA=3�@=J�?=J�>=0>=�_==�<=�;=m�:=�:=99=`8=e�7=�6=��5=��4=�4=�$3=�>2=wV1=�k0=A/=�.=u�-=@�,=f�+=�*=v�)=7�(=�'=��&=!�%=k�$=g�#=��"=k!=�Q =m4=�=��=u�= �=�i=/5=��=�=+= :=��=O�=pQ=[�=�=)B=0�	=�w=i=��=�(=°=�4=-i�<a�<6Q�<�9�<��<e��<
��<���<�W�<��<���<��<�+�<���<Sr�<��<���<S5�<8��<�J�<�ν<O�<�˶<�D�<J��<-�<͜�<
�<�t�<eݝ<�C�<Ө�<-�<�m�<�΋<�.�<э�<~�<��z<Rs<�l<��d<;�]<JV<�O<q�G<�@<}_9<�,2<��*<�#<(�<8�<.q<�[<MM <���;���;���;��;��;%'�;�{�;��;o`�; �m;[5S;O�8;Gb;dB;���:�8�:d\:�p�9�k�8E�;�2��5���y���@�����&$��G;��%R�(�h�V�G����}���B�� 檻f���Ŀ�[ ʻ]ԻF޻p��7���0��R�X������A����a�N�!� �%�!*�dE.��\2�g6��d:��V>�?<B��F���I���M��dQ��U���X�mX\���_��wc��f�vj�5�m�Uq���t��x��n{�'�~����H���^H���兼����F�������C��!֍�uf������䁒���▕�3��E���&,��Ȱ���4�� ����8������S:��㹤��8�������5�������0��@���k+��q����%���������L��� ������f��B�������  �  �vN=��M=��L=�4L=OsK=L�J=��I=�+I=
hH=ţG=��F=+F=�RE=��D=��C=��B=�0B=fA=6�@=L�?=F�>=0>=�_==��<=�;=n�:=�:=99=`8=\�7=��6=��5=��4=�4=�$3=�>2=sV1=l0=8/=�.=o�-==�,=e�+=Թ*=w�)=3�(=��'=��&=)�%=n�$=e�#=��"=k!=�Q =h4=�=��=n�=�=�i=65=��=�=2=(:=��=J�=pQ=L�=ݠ=)B=(�	=�w=_=��=�(=̰=�4=,i�<a�<*Q�<�9�<��<j��<���<���<�W�<��<���<��<�+�<���<Vr�<��<��<b5�<'��<�J�<�ν<O�<�˶<�D�<U��<�,�<Ӝ�<
�<�t�<kݝ<�C�<Ѩ�<�<n�<�΋<�.�<ԍ�<s�<��z< Rs<�l<��d<?�]<�IV<�O<w�G<��@<�_9<�,2<��*<��#</�<e�<7q<�[<3M <���;���;���;��;��;"'�;�{�;��;_`�;4�m;|5S;�8;�b;�B;c��:�8�:Yd\:�l�9�T�8W령P�2�*5��Uz���@����Q&$��F;��%R���h���*����}��C��
檻�f���Ŀ�u ʻԻ�޻4��$���0���Q�f������Y����2a�4�!�
�%�� *�gE.��\2��f6��d:�fV>�R<B��F�&�I���M��dQ��U�q�X��X\���_��wc���f��uj�6�m�Uq�ǹt��x��n{��~����^���\H���兼����=�������C��֍�jf�����ԁ����㖕�E��F���,��̰��w4��,����8��󹡼=:��ݹ���8�������5��{����0��C���h+��|����%���������M����������h��?�������  �  'tN=H�M=!�L=�0L=�nK=��J=��I=c%I=0aH=g�G=��F=�F=�IE=�D=]�C=��B=`%B=�YA=w�@=�?=5�>=P!>=)P==�}<=��;=��:=�9=�%9=L8=xp7=K�6=9�5=U�4={�3=�3=�$2=�;1=2P0=rb/=ir.=�-=��,=��+=o�*=$�)=�(=Ɨ'=��&=*�%=�{$=�k#=mX"=�A!=k' =�	=��=��=��=�l=�;=�=��=��=�O=<
=��=s=2!=�=�p="=J�	=[H=$�=�m=q�=�=�=�<|	�<��<S��<���<���<1x�<�E�<��<V��<���<�;�<���<{��<�5�<e��<'l�<& �<s��<��<F��<-$�<O��<��<d��<��<!�<��<`\�<�ǝ<�0�<R��<4��<�b�<Ƌ<�(�<d��<��<6�z<�Zs<�l<��d<��]<ZgV<'.O<5�G<��@<�9<�c2< :+<�$<��<*�<�<�<]� <hK�;+T�;ll�;��;~λ;Z�;$x�;-�;Tp�;�p;�zU;�;;�� ;e�;1��:Qo�:jg:�!:���8�,��K\'�;T��8���J4���	��!�|&8���N���e�s�{�@����ᓻ"���pH��}ɳ�U(���eȻ�һu{ܻFT�E�ѣ��^��9��
��a����M�Ŭ��� � A%�yv)���-�J�1�U�5���9�J�=�#�A�H�E��YI��!M��P�9�T�J>X�n�[�w_�ec��f��j���m��p�fZt���w��{��j~��܀�����"�������]��'���菊��%��1����J���ڐ��h��v���[���
��:���?������#�������*�������-�������.��)���M-��𫪼�*�������&��ᤰ��"��砳����g������𚹼@�����o���  �  tN=C�M=�L=�0L=�nK=�J=��I=c%I=5aH=c�G=��F=�F=�IE=�D=V�C=��B=_%B=�YA=w�@=�?=5�>=S!>=4P==�}<=��;=��:=�9=�%9=L8=�p7=I�6=:�5=W�4=z�3=�3=�$2=�;1=,P0=wb/=fr.=�-=��,=�+=k�*=!�)=�(=Ǘ'=��&=/�%=�{$=�k#=jX"=�A!=k' =�	=��=��=��=�l=�;=�=��=��=�O=E
=��=s=/!=�=�p= =R�	=WH=(�=�m=p�=��== �<{	�<��<M��<��<���<"x�<�E�<��<`��<���<�;�<���<{��<�5�<e��<-l�<% �<}��<~�<J��<0$�<T��< �<]��<��<"�<��<h\�<�ǝ<�0�<P��<)��<�b�<*Ƌ<�(�<`��<��<�z<�Zs<�l<��d<��]<dgV< .O<8�G<��@<��9<�c2<:+<�$<��<0�<*�<�<q� <IK�;BT�;l�;
��;�λ;#�;Cx�;$�;ap�;�p;�zU;�;;�� ;�;���:�o�:�g:�!:ly�8w3��Z'�vT�����4���	� !��&8���N��e��{�\����ᓻ����H���ɳ�h(���eȻ�һ2{ܻT�7𻘣��l��	9��
�}a����
M������ �A%��v)�i�-�A�1�?�5���9�S�=��A�T�E��YI�"M��P��T�]>X�]�[�-w_�lc��f��j���m��p�ZZt���w�~{��j~��܀�����"������^�����⏊��%��-����J���ڐ��h��l���f��� 
��7���;������#�������*�������-�������.��,���X-������*�������&��٤���"��砳���j������뚹�C�����_���  �  tN=R�M=�L=�0L=�nK=��J=��I=^%I=9aH=_�G=��F=�F=�IE=�D=P�C=��B=\%B=�YA=u�@=�?=8�>=P!>=5P==�}<=��;=��:=�9=�%9=�K8=�p7=C�6==�5=U�4=y�3=�3=�$2=�;1=&P0=}b/=`r.=�-=��,=�+=v�*=�)=�(=��'=��&=,�%=�{$=�k#=eX"=�A!=g' =�	=��=��=��=�l=�;=�=��=��=�O=D
=��=s=,!=�=�p==R�	=PH=-�=�m=t�=��=�=!�<v	�<$��<@��<��<���<7x�<�E�<��<c��<���<�;�<���<|��<�5�<^��<+l�< �<���<r�<N��<+$�<O��< �<R��<��<�<��<[\�<�ǝ<�0�<N��<D��<�b�<1Ƌ<�(�<]��<��<�z<�Zs<�l<�d<p�]<mgV<!.O<"�G<��@<��9<d2<:+<�$<��<�<+�< �<�� <(K�;>T�;ql�;���;�λ;��;\x�;
�;Sp�;�p;�zU;�;;�� ;�;���:�o�: g:�":*��8�5��Y'�8U������Q4��	��!��&8�v�N�C�e���{������ᓻ����H��Bɳ�|(���eȻJ�һJ{ܻ/T�P𻂣��}��9��
��a����M����� �A%��v)�d�-�L�1�M�5���9�u�=��A�a�E�jYI��!M��P��T�y>X�G�[�?w_�Yc��f��j���m��p�JZt���w�p{��j~��܀������"������^�����鏊��%��-����J���ڐ��h��f���r����	��<���@������#�������*�������-�������.��-���=-�����|*��Ǩ���&��Ѥ���"��٠����]�����皹�C�����V���  �  tN=H�M=�L=�0L=�nK= �J=��I=a%I=5aH=b�G=��F=�F=�IE=�D=V�C=��B=b%B=�YA=v�@=�?=8�>=Q!>=1P==�}<=��;=��:=�9=�%9=L8=�p7=G�6=>�5=R�4=w�3=�3=�$2=�;1=&P0=xb/=dr.=�-=��,=�+=k�*=�)=�(=Ɨ'=��&=/�%=�{$=�k#=kX"=�A!=m' =�	=��=��=��=�l=�;=�=��=��=�O=D
=��=s=+!=	�=�p==O�	=SH=)�=�m=r�=��=�=�<r	�< ��<H��<��<���<,x�<�E�<��<c��<���<�;�<���<���<�5�<c��<.l�<) �<���<|�<N��<2$�<X��<��<Z��<��< �<��<b\�<�ǝ<�0�<A��<0��<�b�<%Ƌ<�(�<f��<��<�z<�Zs<|l<��d<n�]<_gV<0.O<&�G<��@<��9<�c2<�9+<�$<��<*�<)�<�<s� <>K�;4T�;�l�; ��;�λ;!�;Xx�;=�;bp�;�p;�zU;�;;�� ;�;���:p�:?g:�:3��8�3��,Z'��T�������4�0�	��!�'8���N�<�e��{�j����ᓻ)����H���ɳ��(���eȻ�һ@{ܻT�/𻪣��h��9���
�|a����M������ �A%�v)�u�-�9�1�C�5���9�P�=��A�g�E��YI�"M��P�#�T�h>X�Y�[�@w_�`c��f��j���m��p�SZt���w��{��j~��܀�����"������ ^�����揊��%��0����J���ڐ��h��f���h����	��6���7������#�������*�������-�������.��;���Q-������*��Ũ���&��٤���"��ߠ����`������;�����b���  �  tN=E�M="�L=�0L=~nK= �J=��I=d%I=2aH=h�G=��F=�F=�IE=�D=W�C=��B=a%B=�YA={�@=�?=5�>=S!>=-P==�}<=�;=��:=�9=�%9=L8=~p7=I�6=9�5=W�4=z�3=�3=�$2=�;1=.P0=xb/=fr.=�-=��,=�+=l�*=*�)=�(=ė'=��&=*�%=�{$=�k#=qX"=�A!=o' =�	=��=��=��=�l=�;=�=��=��=�O=@
=��=s=8!=�=�p==R�	=WH='�=�m=q�=��==�<{	�<��<O��<��<���<*x�<�E�<��<R��<���<�;�<���<|��<�5�<l��<'l�<( �<x��<~�<F��<1$�<[��<��<g��<��<'�<��<b\�<�ǝ<�0�<Z��<)��<�b�< Ƌ<�(�<a��<��<"�z<�Zs<�l<��d<��]<dgV<".O<0�G<��@<��9<�c2<":+<�$<��<-�<�<�<i� <mK�;JT�;�l�;��;uλ;/�;-x�;5�;Qp�;�p;�zU;�;;�� ;��;7��:�n�:�g:F":���8�2���Z'��T��#���4��	��!��&8���N���e��{�W����ᓻ0����H���ɳ�"(���eȻ �һV{ܻFT�+𻻣��O��9���
�ya����M������ �(A%�hv)�z�-�:�1�P�5���9�V�=��A�0�E��YI�"M��P��T�X>X�_�[�"w_�gc��f��j���m��p�aZt���w��{��j~��܀�����"�������]�����䏊��%��0����J���ڐ��h��q���f���
��6���3������#������|*�������-�������.��"���X-��	����*�������&��٤���"��⠳���d������뚹�B��	���g���  �  tN=L�M=�L=�0L=�nK=�J=��I=d%I=5aH=d�G=��F=�F=�IE=��D=V�C=��B=b%B=�YA=x�@=�?=6�>=S!>=3P==�}<=��;=��:=�9=�%9= L8=�p7=E�6=9�5=T�4=y�3=�3=�$2=�;1=&P0=xb/=_r.=�-=��,=�+=q�*= �)=�(=ŗ'=��&=+�%=�{$=�k#=mX"=�A!=k' =�	=��=��=��=�l=�;=�=��=��=�O=F
=��=s=-!=�=�p==Q�	=PH=(�=�m=r�=��=}=�<t	�<��<C��<��<���<1x�<�E�<��<W��<���<�;�<���<y��<�5�<f��<)l�<' �<���<|�<P��<1$�<R��< �<^��<��<%�<��<o\�<�ǝ<�0�<M��<7��<�b�<'Ƌ<�(�<Y��<��<	�z<�Zs<�l<��d<q�]<bgV<.O<,�G<��@<��9<�c2<:+<|$<��<=�<!�<�<r� <MK�;DT�;zl�;��;�λ;&�;lx�;<�;Xp�;�p;�zU;�;;�� ;�;?��:�o�:g:Z!:���8u4���Y'��T��5���h4��	�!��&8���N�3�e��{������ᓻ;����H��oɳ�r(���eȻ�һ{ܻ<T�8𻚣��_��9��
�pa����M������ �A%�wv)�k�-�E�1�P�5���9�T�=��A�Z�E��YI��!M��P��T�t>X�]�[�;w_�bc�$�f��j���m��p�_Zt���w�w{��j~��܀�����"�������]�����䏊��%��+����J���ڐ��h��b���i����	��6���=������#������~*�������-�������.��.���J-������*�������&��ؤ���"��⠳���d��� ��욹�H��
���_���  �  tN=J�M=�L=�0L=�nK=��J=��I=`%I=9aH=d�G=��F=�F=�IE=��D=Q�C=��B=^%B=�YA=v�@=�?=8�>=O!>=2P==�}<=��;=��:=�9=�%9=�K8=�p7=B�6=<�5=O�4=z�3=�3=�$2=�;1=$P0=zb/=_r.=�-=��,=�+=m�*=�)=��(=��'=��&=,�%=�{$=�k#=iX"=�A!=i' =�	=��=��=��=�l=�;=�=��=��=�O=B
=��= s=*!=�=�p==T�	=OH=+�=�m=u�=��=}=!�<i	�<!��<=��<��<���<*x�<�E�<��<n��<���<�;�<���<~��<�5�<`��<3l�<  �<���<u�<Q��<3$�<S��<�<\��<��<�<��<^\�<�ǝ<�0�<E��<4��<�b�<+Ƌ<�(�<Z��<��<�z<�Zs<ml<��d<k�]<WgV<.O<$�G<��@<��9<�c2<�9+<�$<��<�<#�<�<�� <OK�;CT�;�l�;��;�λ;��;vx�;#�;yp�;�p;{U;�;;�� ;��;[��:�p�:�g:� :���8�5���X'�EU������5���	��!�O'8�c�N�Y�e���{������ᓻ/����H���ɳ��(��GeȻ3�һF{ܻ4T�H�q���m���8�	�
�ia����M������ �A%��v)�Y�-�I�1�N�5���9�g�=��A�g�E��YI�"M��P��T�z>X�P�[�Kw_�Tc�1�f��j���m�'�p�OZt�»w�j{�k~��܀�
����"��}���^�����돊��%��#����J���ڐ��h��^���p����	��4���;������#�������*�������-�������.��6���M-������*��¨���&��ڤ���"��ݠ����`�����򚹼E�����Z���  �  tN=I�M=!�L=�0L=~nK= �J=��I=e%I=7aH=g�G=��F=�F=�IE=�D=X�C=��B=`%B=�YA=u�@=�?=7�>=U!>=3P==�}<=��;=��:=�9=�%9=L8=�p7=D�6=:�5=N�4=x�3=�3=�$2=�;1='P0=ub/=br.=�-=��,=�+=q�*="�)=�(='=��&=/�%=�{$=�k#=mX"=�A!=n' =�	=��=��=��=�l=�;=�=��=��=�O=E
=��=s=/!=�=�p==P�	=RH=&�=�m=s�=��=|=�<k	�<��<C��<��<���<'x�<�E�<��<U��<���<�;�<���<z��<�5�<_��<0l�<% �<���<��<N��<3$�<]��<��<a��<��<$�< �<d\�<�ǝ<�0�<S��<5��<�b�<$Ƌ<�(�<]��<��<�z<�Zs<�l<��d<s�]<PgV<.O<"�G<��@<��9<�c2<:+<�$<��<,�<.�<�<{� <dK�;5T�;�l�;��;�λ;6�;bx�;0�;{p�;�p;{U;�;;�� ;�;���:Xo�:�g:�":���854���Y'�U������5��	��!�'8���N�$�e�1�{�t����ᓻ>����H��mɳ�^(���eȻ0�һ1{ܻT�;𻉣��`��9���
�ua����	M������ �A%�{v)�e�-�E�1�<�5���9�]�=��A�S�E�YI�"M� �P��T�l>X�`�[�=w_�\c�*�f��j���m�$�p�\Zt���w�{��j~��܀������"������^����������%��(����J���ڐ��h��e���d����	��5���1������#������*�������-�������.��)���K-������*��ƨ���&��ᤰ��"��ߠ��
��c����������C�����c���  �  tN=E�M=�L=�0L=�nK=�J=��I=h%I=2aH=h�G=��F=�F=�IE=��D=X�C=��B=g%B=�YA=z�@=�?=5�>=V!>=-P==�}<=��;=��:=�9=�%9=L8=}p7=I�6=8�5=T�4=x�3=�3=�$2=�;1=(P0=sb/=er.=�-=��,=�+=j�*=#�)=�(=͗'=��&=,�%=�{$=�k#=rX"=�A!=r' =�	=��=��=��=�l=�;=�=��=��=�O=C
=��=s=/!=	�=�p==L�	=UH="�=�m=n�=��={=�<t	�<��<K��<��<���<$x�<�E�<��<Y��<���<�;�<���<z��<�5�<l��</l�<3 �<���<��<R��<6$�<a��<��<g��<��<,�<��<m\�<�ǝ<�0�<R��<*��<�b�< Ƌ<�(�<c��<��<
�z<�Zs<�l<��d<p�]<VgV<$.O<,�G<��@<��9<�c2<:+<{$<��<=�<�<&�<h� <mK�;JT�;�l�;:��;�λ;7�;cx�;h�;yp�;�p;{U;�;;� ;��;���:�o�:�g:-!:��8f3���Z'�eT��5���_4��	�+!�'8���N��e�X�{�\����ᓻ/����H���ɳ�Z(���eȻ׀һ0{ܻ3T�𻗣��I��9���
�wa����M������ �A%�bv)�e�-�5�1�G�5���9�2�=�!�A�R�E��YI�
"M��P�,�T�^>X�p�[�5w_�pc�&�f��j���m��p�mZt���w��{��j~��܀�����"�������]����������%��$����J���ڐ��h��f���b����	��2���-������#������x*�������-��~����.��)���W-������*��Ĩ���&��ᤰ��"��𠳼��s��� ��򚹼A��
���g���  �  tN=K�M=�L=�0L=�nK=��J=��I=f%I=5aH=e�G=��F=�F=�IE=��D=T�C=��B=_%B=�YA={�@=�?=7�>=V!>=/P==�}<=��;=��:=�9=�%9=�K8=p7=B�6=8�5=R�4=x�3=�3=�$2=�;1=(P0=wb/=`r.=�-=��,=�+=n�*="�)=�(=��'=��&=,�%=�{$=�k#=nX"=�A!=m' =�	= �=��=��=�l=�;=�=��=��=�O=>
=��=s=0!=�=�p==L�	=PH=&�=�m=p�=��=|=�<o	�<��<?��<��<���<0x�<�E�<��<`��<���<�;�<���<~��<�5�<i��<0l�<$ �<���<|�<V��<.$�<Y��<�<c��<��<(�<��<Y\�<�ǝ<�0�<O��<3��<�b�<(Ƌ<�(�<Z��<��<�z<�Zs<l<��d<u�]<UgV<.O<�G<��@<��9<�c2<:+<�$<��<�<!�<!�<t� <]K�;hT�;�l�;��;�λ;�;lx�;-�;zp�;p;�zU;�;;� ;ؼ;;��:�o�:�g:)!:��8�4��FZ'�8U��.����4��	��!�'8���N��e��{������ᓻ����H���ɳ�[(��{eȻ<�һg{ܻ/T�.𻜣��Z��9���
�ta�����L������ �A%�rv)�o�-�?�1�H�5���9�h�=��A�M�E��YI�"M��P�)�T�t>X�`�[�:w_�fc�*�f��j���m��p�bZt���w��{��j~��܀�����"������^�����Ꮚ��%��+����J���ڐ��h��e���h����	��9���5������#������|*�������-�������.��,���N-������*��ɨ���&��ߤ���"��䠳���h������򚹼G�����`���  �  tN=L�M=�L=�0L=�nK=�J=�I=a%I=;aH=d�G=��F=�F=�IE=��D=Z�C=��B=_%B=�YA=w�@=�?=<�>=Q!>=:P==�}<=��;=��:=�9=�%9=�K8=�p7=>�6=;�5=M�4=u�3=�3=�$2=�;1="P0=vb/=]r.=�-=��,=�+=p�*=�)=�(=��'=��&=1�%=�{$=�k#=jX"=�A!=n' =�	= �=��=��=�l=�;=�=��=��=�O=J
=��=s=&!=�=�p==P�	=KH=&�=�m=p�=��={=�<d	�<��<3��<��<���<+x�<�E�<��<\��<���<�;�<���<���<�5�<a��<9l�<# �<���<��<W��<2$�<_��<�<]��<��<�<	�<n\�<�ǝ<�0�<=��<:��<�b�<)Ƌ<�(�<Y��<��<��z<�Zs<gl<��d<b�]<KgV<.O<�G<��@<��9<�c2<�9+<�$<��<5�<D�<�<�� <PK�;KT�;�l�;��;�λ;I�;�x�;+�;�p�;�p;�zU;;;�� ;��;���:�o�:�g:� :l��8�6���X'��U��ڂ��B5�D�	�!�X'8���N�x�e�'�{������ᓻ7����H��oɳ��(��zeȻ4�һ{ܻT�.�~���i���8���
�la�����L������ ��@%��v)�a�-�6�1�>�5���9�b�=��A�v�E��YI�"M�#�P��T��>X�^�[�Uw_�fc�3�f��j���m�0�p�WZt�Իw�q{�k~��܀�����"������^�����珊��%��*����J���ڐ��h��^���_����	��6���/��
����#�������*�������-�������.��?���G-������*��ʨ���&��⤰��"��⠳���e���������E�����[���  �  tN=K�M=�L=�0L=�nK=�J=��I=e%I=6aH=j�G=��F=�F=�IE=�D=Z�C=��B=e%B=�YA=z�@=�?=9�>=Q!>=-P==�}<=��;=��:=�9=�%9= L8=�p7=C�6=;�5=O�4=x�3=�3=�$2=�;1=&P0=wb/=ar.=�-=��,=�+=o�*=!�)=�(=ŗ'=��&='�%=�{$=�k#=pX"=�A!=q' =�	=��=��=��=�l=�;=�=��=��=�O=A
=��=s=/!=�=�p==P�	=OH='�=�m=n�=��={=�<k	�<��<<��<��<���</x�<�E�<��<[��<���<�;�<���<���<�5�<k��<.l�</ �<}��<��<N��<7$�<a��<��<h��<��<(�<��<f\�<�ǝ<�0�<N��<8��<�b�<"Ƌ<�(�<]��<��<�z<�Zs<�l<��d<h�]<RgV<.O<�G<��@<��9<�c2<:+<�$<��<1�<�<�<x� <~K�;FT�;�l�;9��;�λ;H�;Ox�;[�;xp�;�p;8{U;�;;�� ;��;��:�o�:�g:�!:��8�4���Y'�"U��ゴ��4��	�!�'8���N�0�e��{�z����ᓻ2����H��vɳ�e(���eȻ�һG{ܻTT�𻕣��P��	9���
�ta�����L������ �A%�hv)�f�-�.�1�[�5���9�U�=��A�R�E��YI��!M��P��T�t>X�]�[�Bw_�mc�$�f��j���m�!�p�ZZt�»w�}{��j~��܀�����"������ ^�����쏊��%��#����J���ڐ��h��k���^����	��1���-������#������{*�������-�������.��-���H-������*��ɨ���&��ޤ���"��頳���k�����󚹼D�����c���  �  tN=C�M=�L=�0L=�nK=�J=��I=u%I=-aH=j�G=��F=�F=�IE=�D=_�C=��B=l%B=�YA={�@=�?=4�>=c!>=3P==�}<=�;=��:=�9=�%9=�K8=yp7=G�6=8�5=N�4=u�3=�3=�$2=|;1='P0=tb/=ar.=�-=��,=�+=e�*=%�)=�(=Ɨ'=��&=0�%=�{$=�k#=tX"=�A!=s' =�	=�=��=��=�l=�;=�=��=��=�O=D
=��=s=2!=�=�p==J�	=PH=$�=�m=i�=��=z=�<j	�<��<D��<���<���<$x�<�E�<��<N��<���<�;�<��<|��<�5�<p��<#l�<< �<}��<��<P��<:$�<^��<��<l��<��<F�<��<l\�<�ǝ<�0�<S��<$��<�b�<"Ƌ<�(�<Z��<��<�z<�Zs<�l<��d<m�]<LgV<.O<,�G<��@<��9<�c2<:+<�$<��<?�< �<Z�<V� <}K�;MT�;�l�;\��;�λ;p�;Nx�;��;Up�;p;�zU;�;;�� ;�;?��:o�:�g:� :�8�4���['��T��I���"5�?�	�<!��&8�(�N�(�e�F�{�v����ᓻ8����H���ɳ�D(���eȻ�һ4{ܻT���ԣ��@��9���
�sa�����L������ �#A%�Tv)���-�!�1�.�5���9�K�=�!�A�F�E��YI�"M�$�P�2�T�p>X�i�[�@w_��c��f��j���m�$�p�fZt���w��{��j~��܀�����"�������]�����ɏ���%��/����J���ڐ��h��k���T����	��-���0������#������^*�������-�������.��)���]-������*��Ĩ���&��ᤰ��"��𠳼���p���������I��
���j���  �  tN=K�M=�L=�0L=�nK=�J=��I=e%I=6aH=j�G=��F=�F=�IE=�D=Z�C=��B=e%B=�YA=z�@=�?=9�>=Q!>=-P==�}<=��;=��:=�9=�%9= L8=�p7=C�6=;�5=O�4=x�3=�3=�$2=�;1=&P0=wb/=ar.=�-=��,=�+=o�*=!�)=�(=ŗ'=��&='�%=�{$=�k#=pX"=�A!=q' =�	=��=��=��=�l=�;=�=��=��=�O=A
=��=s=/!=�=�p==P�	=OH='�=�m=n�=��={=�<k	�<��<<��<��<���</x�<�E�<��<[��<���<�;�<���<���<�5�<k��<.l�</ �<}��<��<N��<7$�<a��<��<h��<��<(�<��<f\�<�ǝ<�0�<N��<8��<�b�<"Ƌ<�(�<]��<��<�z<�Zs<�l<��d<h�]<RgV<.O<�G<��@<��9<�c2<:+<�$<��<1�<�<�<x� <~K�;FT�;�l�;9��;�λ;H�;Ox�;[�;xp�;�p;8{U;�;;�� ;��;��:�o�:�g:�!:t��8�4���Y'�#U��ゴ��4��	�!�'8���N�0�e��{�z����ᓻ2����H��vɳ�e(���eȻ�һG{ܻTT�𻕣��P��	9���
�ta�����L������ �A%�hv)�f�-�.�1�[�5���9�U�=��A�R�E��YI��!M��P��T�t>X�]�[�Bw_�mc�$�f��j���m�!�p�ZZt�»w�}{��j~��܀�����"������ ^�����쏊��%��#����J���ڐ��h��k���^����	��1���-������#������{*�������-�������.��-���H-������*��ɨ���&��ޤ���"��頳���k�����󚹼D�����c���  �  tN=L�M=�L=�0L=�nK=�J=�I=a%I=;aH=d�G=��F=�F=�IE=��D=Z�C=��B=_%B=�YA=w�@=�?=<�>=Q!>=:P==�}<=��;=��:=�9=�%9=�K8=�p7=>�6=;�5=M�4=u�3=�3=�$2=�;1="P0=vb/=]r.=�-=��,=�+=p�*=�)=�(=��'=��&=1�%=�{$=�k#=jX"=�A!=n' =�	= �=��=��=�l=�;=�=��=��=�O=J
=��=s=&!=�=�p==P�	=KH=&�=�m=p�=��=|=�<d	�<��<3��<��<���<+x�<�E�<��<]��<���<�;�<���<���<�5�<a��<9l�<# �<���<��<W��<2$�<_��<�<]��<��<�<	�<n\�<�ǝ<�0�<=��<:��<�b�<)Ƌ<�(�<Y��<��<��z<�Zs<gl<��d<b�]<KgV<.O<�G<��@<��9<�c2<�9+<�$<��<5�<D�<�<�� <PK�;KT�;�l�;��;�λ;I�;�x�;+�;�p�;�p;�zU;;;�� ;��;���:�o�:�g:� :U��8�6���X'��U��ۂ��C5�E�	�!�Y'8���N�x�e�'�{������ᓻ7����H��oɳ��(��zeȻ4�һ{ܻT�/�~���i���8���
�la�����L������ ��@%��v)�a�-�6�1�>�5���9�b�=��A�v�E��YI�"M�#�P��T��>X�_�[�Uw_�fc�3�f��j���m�0�p�WZt�Իw�q{�k~��܀�����"������^�����珊��%��*����J���ڐ��h��^���_����	��6���/��
����#�������*�������-�������.��?���G-������*��ʨ���&��⤰��"��⠳���e���������E�����[���  �  tN=K�M=�L=�0L=�nK=��J=��I=f%I=5aH=e�G=��F=�F=�IE=��D=T�C=��B=_%B=�YA={�@=�?=7�>=V!>=/P==�}<=��;=��:=�9=�%9=�K8=p7=B�6=8�5=R�4=x�3=�3=�$2=�;1=(P0=wb/=`r.=�-=��,=�+=n�*="�)=�(=��'=��&=,�%=�{$=�k#=nX"=�A!=m' =�	= �=��=��=�l=�;=�=��=��=�O=>
=��=s=0!=�=�p==L�	=PH=&�=�m=p�=��=|=�<o	�<��<?��<��<���<0x�<�E�<��<`��<���<�;�<���<~��<�5�<i��<0l�<$ �<���<|�<V��<.$�<Y��<�<c��<��<'�<��<Y\�<�ǝ<�0�<O��<3��<�b�<(Ƌ<�(�<Z��<��<�z<�Zs<l<��d<u�]<UgV<.O<�G<��@<��9<�c2<:+<�$<��<�<!�<!�<t� <]K�;hT�;�l�;��;�λ;�;lx�;,�;zp�;p;�zU;�;;� ;׼;:��:�o�:�g:%!:Ɗ�8�4��JZ'�:U��0����4��	��!�'8���N��e��{������ᓻ����H���ɳ�[(��{eȻ<�һg{ܻ/T�/𻜣��Z��9���
�ta�����L������ �A%�rv)�o�-�?�1�H�5���9�h�=��A�M�E��YI�"M��P�)�T�t>X�`�[�:w_�fc�*�f��j���m��p�bZt���w��{��j~��܀�����"������^�����Ꮚ��%��+����J���ڐ��h��e���h����	��9���5������#������|*�������-�������.��,���N-������*��ɨ���&��ߤ���"��䠳���h������򚹼G�����`���  �  tN=E�M=�L=�0L=�nK=�J=��I=h%I=2aH=h�G=��F=�F=�IE=��D=X�C=��B=g%B=�YA=z�@=�?=5�>=V!>=-P==�}<=��;=��:=�9=�%9=L8=}p7=I�6=8�5=T�4=x�3=�3=�$2=�;1=(P0=sb/=er.=�-=��,=�+=j�*=#�)=�(=͗'=��&=,�%=�{$=�k#=rX"=�A!=r' =�	=��=��=��=�l=�;=�=��=��=�O=C
=��=s=/!=	�=�p==L�	=UH="�=�m=n�=��={=�<t	�<��<K��<��<���<$x�<�E�<��<Y��<���<�;�<���<z��<�5�<l��</l�<3 �<���<��<R��<6$�<a��<��<g��<��<,�<��<m\�<�ǝ<�0�<R��<*��<�b�< Ƌ<�(�<c��<��<
�z<�Zs<�l<��d<p�]<VgV<$.O<,�G<��@<��9<�c2<:+<{$<��<=�<�<'�<h� <mK�;JT�;�l�;:��;�λ;7�;cx�;h�;xp�;�p;{U;�;;� ;��;���:�o�:�g:(!:��8p3���Z'�hT��7���b4��	�,!�	'8���N��e�Y�{�\����ᓻ0����H���ɳ�Z(���eȻ׀һ0{ܻ3T�𻘣��I��9���
�wa����M������ �A%�bv)�e�-�5�1�G�5���9�2�=�!�A�R�E��YI�
"M��P�,�T�^>X�p�[�5w_�pc�&�f��j���m��p�mZt���w��{��j~��܀�����"�������]����������%��$����J���ڐ��h��f���b����	��2���-������#������x*�������-��~����.��)���W-������*��Ĩ���&��ᤰ��"��𠳼��s��� ��򚹼A��
���g���  �  tN=I�M=!�L=�0L=~nK= �J=��I=e%I=7aH=g�G=��F=�F=�IE=�D=X�C=��B=`%B=�YA=u�@=�?=7�>=U!>=3P==�}<=��;=��:=�9=�%9=L8=�p7=D�6=:�5=N�4=x�3=�3=�$2=�;1='P0=ub/=br.=�-=��,=�+=q�*="�)=�(='=��&=/�%=�{$=�k#=mX"=�A!=n' =�	=��=��=��=�l=�;=�=��=��=�O=E
=��=s=/!=�=�p==P�	=RH='�=�m=s�=��=|=�<k	�<��<C��<��<���<'x�<�E�<��<U��<���<�;�<���<z��<�5�<_��<0l�<% �<���<��<N��<3$�<]��<��<a��<��<$�<��<d\�<�ǝ<�0�<S��<5��<�b�<$Ƌ<�(�<]��<��<�z<�Zs<�l<��d<s�]<PgV<.O<"�G<��@<��9<�c2<:+<�$<��<,�<.�<�<{� <dK�;5T�;�l�;��;�λ;6�;bx�;0�;zp�;�p;{U;�;;�� ;�;���:Vo�:�g:�":���8@4���Y'�U������5��	��!�'8���N�%�e�2�{�t����ᓻ>����H��mɳ�_(���eȻ0�һ1{ܻT�;𻉣��`��9���
�ua����	M������ �A%�{v)�e�-�E�1�=�5���9�]�=��A�S�E�YI�"M� �P��T�l>X�`�[�=w_�\c�*�f��j���m�$�p�\Zt���w�{��j~��܀������"������^����������%��(����J���ڐ��h��e���d����	��5���1������#������*�������-�������.��)���K-������*��ƨ���&��ᤰ��"��ߠ��
��c����������C�����c���  �  tN=J�M=�L=�0L=�nK=��J=��I=`%I=9aH=d�G=��F=�F=�IE=��D=Q�C=��B=^%B=�YA=v�@=�?=8�>=O!>=2P==�}<=��;=��:=�9=�%9=�K8=�p7=B�6=<�5=O�4=z�3=�3=�$2=�;1=$P0=zb/=_r.=�-=��,=�+=m�*=�)=��(=��'=��&=,�%=�{$=�k#=iX"=�A!=i' =�	=��=��=��=�l=�;=�=��=��=�O=B
=��= s=*!=�=�p==T�	=OH=+�=�m=u�=��=}=!�<j	�<!��<=��<��<���<*x�<�E�<��<n��<���<�;�<���<~��<�5�<`��<3l�<  �<���<u�<Q��<3$�<S��<�<\��<��<�<��<^\�<�ǝ<�0�<E��<4��<�b�<+Ƌ<�(�<Z��<��<�z<�Zs<ml<��d<k�]<WgV<.O<$�G<��@<��9<�c2<�9+<�$<��<�<#�<�<�� <PK�;CT�;�l�;��;�λ;��;vx�;"�;yp�;�p;{U;�;;�� ;��;Y��:�p�:�g:� :{��86���X'�HU������5���	��!�Q'8�e�N�Z�e���{������ᓻ/����H���ɳ��(��GeȻ3�һG{ܻ4T�I�q���m���8�	�
�ia����M������ �A%��v)�Y�-�I�1�N�5���9�g�=��A�g�E��YI�"M��P��T�z>X�P�[�Kw_�Tc�1�f��j���m�'�p�OZt�»w�j{�k~��܀�
����"��}���^�����돊��%��#����J���ڐ��h��^���p����	��4���;������#�������*�������-�������.��6���M-������*��¨���&��ڤ���"��ݠ����`�����򚹼E�����Z���  �  tN=L�M=�L=�0L=�nK=�J=��I=d%I=5aH=d�G=��F=�F=�IE=��D=V�C=��B=b%B=�YA=x�@=�?=6�>=S!>=3P==�}<=��;=��:=�9=�%9= L8=�p7=E�6=9�5=T�4=y�3=�3=�$2=�;1=&P0=xb/=_r.=�-=��,=�+=q�*= �)=�(=ŗ'=��&=+�%=�{$=�k#=mX"=�A!=k' =�	=��=��=��=�l=�;=�=��=��=�O=F
=��=s=-!=�=�p==Q�	=PH=(�=�m=r�=��=}=�<t	�<��<D��<��<���<1x�<�E�<��<X��<���<�;�<���<y��<�5�<f��<*l�<' �<���<|�<P��<1$�<R��< �<^��<��<%�<��<o\�<�ǝ<�0�<M��<7��<�b�<'Ƌ<�(�<Y��<��<	�z<�Zs<�l<��d<q�]<bgV<.O<,�G<��@<��9<�c2<:+<}$<��<=�<"�<�<r� <MK�;ET�;zl�;��;�λ;&�;lx�;<�;Wp�;�p;�zU;�;;�� ;�;=��:~o�:g:T!:]��8�4���Y'��T��7���k4��	�!��&8���N�4�e��{������ᓻ<����H��oɳ�r(���eȻ�һ{ܻ=T�8𻚣��_��9��
�pa����M������ �A%�wv)�k�-�E�1�P�5���9�T�=��A�Z�E��YI��!M��P��T�t>X�]�[�;w_�bc�$�f��j���m��p�_Zt���w�w{��j~��܀�����"�������]�����䏊��%��+����J���ڐ��h��b���i����	��6���=������#������~*�������-�������.��.���J-������*�������&��ؤ���"��⠳���d��� ��욹�H��
���_���  �  tN=E�M="�L=�0L=~nK= �J=��I=d%I=2aH=h�G=��F=�F=�IE=�D=W�C=��B=a%B=�YA={�@=�?=5�>=S!>=-P==�}<=�;=��:=�9=�%9=L8=~p7=I�6=9�5=W�4=z�3=�3=�$2=�;1=.P0=xb/=fr.=�-=��,=�+=l�*=*�)=�(=ė'=��&=*�%=�{$=�k#=qX"=�A!=o' =�	=��=��=��=�l=�;=�=��=��=�O=@
=��=s=8!=�=�p==R�	=WH='�=�m=q�=��==�<{	�<��<O��<��<���<*x�<�E�<��<R��<���<�;�<���<|��<�5�<l��<'l�<( �<x��<~�<F��<1$�<[��<��<g��<��<'�<��<b\�<�ǝ<�0�<Z��<)��<�b�< Ƌ<�(�<a��<��<"�z<�Zs<�l<��d<��]<dgV<#.O<0�G<��@<��9<�c2<":+<�$<��<-�<�<�<i� <mK�;JT�;�l�;��;uλ;/�;-x�;5�;Qp�;�p;�zU;�;;�� ;��;5��:�n�:�g:A":���8�2���Z'��T��&���4��	��!��&8���N���e��{�W����ᓻ1����H���ɳ�"(���eȻ �һV{ܻFT�+𻻣��O��9���
�ya����M������ �(A%�hv)�z�-�:�1�P�5���9�V�=��A�0�E��YI�"M��P��T�X>X�_�[�"w_�gc��f��j���m��p�aZt���w��{��j~��܀�����"�������]�����䏊��%��0����J���ڐ��h��q���f���
��6���3������#������|*�������-�������.��!���X-��	����*�������&��٤���"��⠳���d������뚹�B��	���g���  �  tN=H�M=�L=�0L=�nK= �J=��I=a%I=5aH=b�G=��F=�F=�IE=�D=V�C=��B=b%B=�YA=v�@=�?=8�>=Q!>=1P==�}<=��;=��:=�9=�%9=L8=�p7=G�6=>�5=R�4=w�3=�3=�$2=�;1=&P0=xb/=dr.=�-=��,=�+=k�*=�)=�(=Ɨ'=��&=/�%=�{$=�k#=kX"=�A!=m' =�	=��=��=��=�l=�;=�=��=��=�O=D
=��=s=+!=	�=�p==O�	=SH=)�=�m=r�=��=�=�<r	�< ��<H��<��<���<,x�<�E�<��<c��<���<�;�<���<���<�5�<c��<.l�<) �<���<|�<N��<2$�<X��<��<Z��<��< �<��<b\�<�ǝ<�0�<A��<0��<�b�<%Ƌ<�(�<f��<��<�z<�Zs<|l<��d<n�]<_gV<0.O<&�G<��@<��9<�c2<�9+<�$<��<*�<)�<�<s� <>K�;4T�;�l�; ��;�λ;!�;Xx�;=�;bp�;�p;�zU;�;;�� ;�;���:p�:;g:�:��8�3��0Z'��T�������4�1�	��!�'8���N�=�e��{�k����ᓻ)����H���ɳ��(���eȻ�һ@{ܻT�/𻪣��h��9���
�|a����M������ �A%�v)�u�-�9�1�C�5���9�P�=��A�g�E��YI�"M��P�#�T�h>X�Y�[�@w_�`c��f��j���m��p�SZt���w��{��j~��܀�����"������ ^�����揊��%��0����J���ڐ��h��f���h����	��6���7������#�������*�������-�������.��;���Q-������*��Ũ���&��٤���"��ߠ����`������;�����b���  �  tN=R�M=�L=�0L=�nK=��J=��I=^%I=9aH=_�G=��F=�F=�IE=�D=P�C=��B=\%B=�YA=u�@=�?=8�>=P!>=5P==�}<=��;=��:=�9=�%9=�K8=�p7=C�6==�5=U�4=y�3=�3=�$2=�;1=&P0=}b/=`r.=�-=��,=�+=v�*=�)=�(=��'=��&=,�%=�{$=�k#=eX"=�A!=g' =�	=��=��=��=�l=�;=�=��=��=�O=D
=��=s=,!=�=�p==R�	=PH=-�=�m=t�=��=�=!�<v	�<$��<@��<��<���<7x�<�E�<��<c��<���<�;�<���<|��<�5�<^��<+l�< �<���<s�<N��<+$�<O��< �<R��<��<�<��<[\�<�ǝ<�0�<N��<D��<�b�<1Ƌ<�(�<]��<��<�z<�Zs<�l<�d<p�]<mgV<!.O<"�G<��@<��9<d2<:+<�$<��<�<+�< �<�� <(K�;>T�;ql�;���;�λ;��;[x�;
�;Sp�;�p;�zU;�;;�� ;�;���:�o�:�g:�":��8�5��Y'�9U������S4��	��!��&8�w�N�D�e���{������ᓻ����H��Bɳ�|(���eȻJ�һJ{ܻ/T�Q𻂣��}��9��
��a����M����� �A%��v)�d�-�L�1�M�5���9�u�=��A�a�E�jYI��!M��P��T�y>X�G�[�?w_�Yc��f��j���m��p�JZt���w�p{��j~��܀������"������^�����鏊��%��-����J���ڐ��h��f���r����	��<���@������#�������*�������-�������.��-���=-�����|*��Ǩ���&��Ѥ���"��٠����]�����皹�C�����V���  �  tN=C�M=�L=�0L=�nK=�J=��I=c%I=5aH=c�G=��F=�F=�IE=�D=V�C=��B=_%B=�YA=w�@=�?=5�>=S!>=4P==�}<=��;=��:=�9=�%9=L8=�p7=I�6=:�5=W�4=z�3=�3=�$2=�;1=,P0=wb/=fr.=�-=��,=�+=k�*=!�)=�(=Ǘ'=��&=/�%=�{$=�k#=jX"=�A!=k' =�	=��=��=��=�l=�;=�=��=��=�O=E
=��=s=/!=�=�p= =R�	=WH=(�=�m=p�=��== �<{	�<��<M��<��<���<"x�<�E�<��<`��<���<�;�<���<{��<�5�<e��<-l�<% �<}��<~�<J��<0$�<T��< �<]��<��<"�<��<h\�<�ǝ<�0�<P��<)��<�b�<*Ƌ<�(�<`��<��<�z<�Zs<�l<��d<��]<dgV< .O<8�G<��@<��9<�c2<:+<�$<��<0�<*�<�<q� <IK�;BT�;l�;
��;�λ;#�;Cx�;$�;ap�;�p;�zU;�;;�� ;�;���:�o�:�g:�!:_y�8y3��Z'�vT�����4���	�!��&8���N��e��{�\����ᓻ����H���ɳ�h(���eȻ�һ2{ܻT�7𻘣��l��	9��
�}a����
M������ �A%��v)�i�-�A�1�?�5���9�S�=��A�T�E��YI�"M��P��T�]>X�]�[�-w_�lc��f��j���m��p�ZZt���w�~{��j~��܀�����"������^�����⏊��%��-����J���ڐ��h��l���f��� 
��7���;������#�������*�������-�������.��,���X-������*�������&��٤���"��砳���j������뚹�C�����_���  �  rqN=1�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=LAE=�xD=ͯC=��B=�B=�NA=��@=s�?=�>=�>=�A==�n<=<�;=O�:=��9=�9=f98= ]7=+6=Q�5=��4=��3=O�2=�2=�"1=b60=�G/=�V.=vc-=ym,=�t+=�y*=\{)=Lz(=Uv'=@o&=e%=�W$= G#= 3"=�!=�  =��=ÿ=ؙ=)p=�B=6=��=�=#e=�#=%�=��=�F=��=��=OD=��
=@�	=�=��=�B=��=�X=�� =��<���<ʫ�<���<�{�<)Y�<x/�<��<���<r��<�F�<���<b��<X�<k��<���<�8�<���<�`�<��<5w�<���<~�<8��<w�<��<�c�<�դ<�E�<x��<�<��<R�<IX�<��<#�<(��<��<S�z<�bs<y)l<��d<�]<��V<NO<�H<N�@<�9<��2<�q+<Q$<65<[<�<�<�� <���;��;O1�;1c�;ǥ�;t��;�a�;�ܓ;}k�;�r;��W;�4=;�#;l	;�s�:�?�:��p:"4:(Z!9��j�G����}����J�޺u��I3��D5��L���b���x�����f���)��$̧�M�������ƻ�ѻRۻ��仏��y5��
� �Ѕ��#
�ٲ��2�����>Z �v�$���(�8-�J"1��35��89��1=��A�� E�r�H���L�.eP��T���W� o[�X
_��b�('f�C�i��#m�>�p��t�Jfw�`�z��~�����z\������򟅼�=��Bو�\r��a	��I���/1��W��Q��hߓ��k��F�������������T��3��������^"������%��s����%��+����$�������"��}���K ��7���.��t���������������������  �  rqN=0�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=MAE=�xD=үC=��B=�B=�NA=��@=p�?=!�>=�>=�A==�n<==�;=R�:=��9=�9=i98=(]7=*6=W�5=��4=��3=I�2=2=�"1=]60=�G/=�V.=zc-=�m,=�t+=�y*=]{)=Sz(=Nv'=>o&=e%=�W$=G#=�2"=�!=�  =��=ȿ=ݙ=-p=�B=7=��=��="e=�#=%�=~�=�F=��=��=OD=��
=D�	=�=��=�B=��=�X=�� =��<���<ի�<���<�{�<0Y�<z/�<	��<���<x��<�F�<���<X��<X�<l��<���<�8�<���<�`�<��<Cw�<���<~�</��<�v�<��<�c�<�դ<�E�<o��<�<��<P�<JX�<$��<#�<0��<��<E�z<�bs<G)l<��d<�]<��V<(NO<�H<n�@<�9<�2<�q+</Q$<,5<F<<�<�� <J��;��;g1�;;c�;���;���;�a�;�ܓ;�k�;Cr;l�W;35=;�#;�	;�r�:@�:��p:}3:�[!9Ӏj�b����}����b�޺����3��E5��L��b���x������e���)��!̧�M��������ƻ ѻ]ۻ��仡��G5��*� �҅��#
�ʲ��2�����:Z �s�$��(�&-�K"1��35��89��1=��A�� E�t�H���L�eP��T���W�
o[�g
_��b�Q'f�]�i��#m�J�p��t�Nfw�G�z��~�����~\������쟅��=��>و�er��[	��I���A1��S��Q��]ߓ��k��8�������������d��"��������d"�������$��v����%��*���~$�������"��v���R ��:���G��x���������������������  �  oqN=5�M=��L=�,L=jK=�J=��I={I=�ZH=��G=��F=�F=HAE=�xD=ͯC=��B=�B=�NA=��@=t�?="�>=�>=�A==�n<=>�;=S�:=��9=�9=f98=']7=$6=X�5=��4=��3=Q�2=�2=�"1=Z60=�G/=�V.=tc-=}m,=�t+=�y*=Y{)=Tz(=Lv'=Eo&=e%=�W$=	G#=�2"=�!=�  =��=Ŀ=ٙ=)p=�B=<=��=��= e=�#=-�=|�=�F=��=��=PD=��
=A�	=�=��=�B=��=�X=�� =��<���<ګ�<{��<�{�<+Y�<}/�<��<���<{��<�F�<��<P��<X�<u��<���<�8�<���<�`�<��<>w�<���<~�<=��<�v�<��<�c�<�դ<�E�<i��<�<���<X�<HX�<!��<�"�<-��<��<?�z<�bs<Z)l<��d<ݸ]<��V<%NO<�H<h�@<�9<�2<�q+<2Q$<&5<Q<<�<�� <f��;��;j1�;c�;�;x��;�a�;|ܓ;�k�;�r;��W;65=;@#;�	;�r�:C@�:��p:�2:�^!9��j������}������޺v��&3�UE5�RL��b�X�x�����(f���)��̧��L��������ƻ2ѻ%ۻ������05��#� �����#
�ݲ��2�����BZ �]�$��(�-�U"1��35��89��1=��A�� E�n�H���L�%eP��T���W��n[�r
_��b�6'f�=�i�#m�T�p��t�efw�O�z��~������\������韅��=��0و�nr��\	��@���81��K��Q��cߓ��k��<�������������^����������["������$��}���|%��,����$�������"��s���U ��*���>��g���������������������  �  qqN=4�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=NAE=�xD=ԯC=��B=�B=�NA=��@=p�?= �>=�>=�A==�n<=<�;=S�:=��9=�9=h98=&]7=(6=S�5=��4=��3=K�2=�2=�"1=^60=�G/=�V.=yc-=}m,=�t+=�y*=Z{)=Pz(=Qv'=?o&=e%=�W$= G#=�2"=�!=�  =��=ɿ=ޙ=+p=�B=5=��=�=$e=�#=%�=��=�F=��=��=SD=��
=C�	=�=��=�B=��=�X=�� =��<���<ϫ�<���<�{�<.Y�<~/�<��<���<s��<�F�<���<Y��<X�<i��<���<�8�<���<�`�<��<Bw�<���<~�<3��<w�<��<�c�<�դ<�E�<s��<�<���<V�<MX�<��<#�<*��<��<J�z<�bs<V)l<��d<�]<��V<NO<�H<f�@<�9<�2<�q+<'Q$<05<R<�<�<�� <s��;��;E1�;Dc�;���;���;�a�;�ܓ;xk�;�r;s�W;5=;�#;f	;Ts�:�?�:��p:�2:�^!9n�j�ذ�_�}�8���޺����3�xE5��L�ۦb���x�퀇�f���)�� ̧�M��������ƻѻ[ۻ��仔��u5��� �҅��#
�ϲ��2�����9Z �z�$���(�5-�F"1��35��89��1=��A�� E�s�H�w�L�eP��T���W�o[�a
_��b�E'f�S�i��#m�=�p��t�Tfw�O�z��~������\������🅼�=��Bو�dr��^	��K���21��Y��Q��^ߓ��k��8�������������X��-��������a"������%��z���~%��(����$�������"��x���O ��=���@��w���������������������  �  rqN=.�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=OAE=�xD=կC=��B=�B=�NA=��@=p�?=!�>=�>=�A==�n<=7�;=V�:=��9=�9=h98=#]7=,6=P�5=��4=��3=L�2=�2=�"1=a60=�G/=�V.=xc-=}m,=�t+=y*=_{)=Mz(=Sv'=>o&=e%=�W$= G#=3"=�!=�  =��=ſ=ܙ=%p=�B=4=��=~�=(e=�#=$�=��=�F=��=��=QD=��
=@�	=�=��=�B=��=�X=�� =��<ĸ�<ƫ�<���<�{�</Y�<y/�<��<���<l��<�F�<���<c��< X�<h��<���<�8�<���<�`�<��<7w�<���<~�<,��<w�<��<�c�<�դ<�E�<r��<�<��<I�<MX�<��<#�<&��<��<R�z<�bs<t)l<��d<�]<��V<NO<H<Y�@<��9<�2<�q+<2Q$<(5<U<�<�<�� <t��;��;^1�;Hc�;ƥ�;���;�a�;�ܓ;�k�;�r;j�W;15=;#;?	;�s�:e?�:��p:�2:�Z!9u�j�����}������޺���q3�E5�L���b���x�����	f���)��̧�)M��}���	�ƻ�ѻ\ۻ���d��t5��� �څ��#
����2�����.Z ��$���(�;-�5"1��35��89��1=��A�� E���H���L� eP��T���W�(o[�W
_��b�*'f�F�i��#m�6�p��t�Ifw�]�z��~������\�����������=��Hو�Zr��X	��M���/1��Z��Q��lߓ�k��D�������������V��-���������`"�������$��r����%��(����$�������"�����L ��A���1��z���������������������  �  sqN=2�M=��L=�,L=	jK=�J=��I=|I=�ZH=��G=��F=�F=KAE=�xD=ׯC=��B=�B=�NA=��@=s�?= �>=�>=�A==�n<=:�;=U�:=��9=�9=h98=$]7=&6=W�5=��4=��3=K�2=�2=�"1=Y60=�G/=�V.=uc-=|m,=�t+=�y*=[{)=Qz(=Lv'=Go&=e%=�W$=G#=�2"=�!=�  =��=˿=�=)p=�B=8=��=��=!e=�#=-�=|�=�F=��=��=QD=��
=>�	=�=��=�B=��=�X=�� =��<���<ի�<��<�{�<,Y�<~/�<��<���<t��<�F�<���<T��<X�<p��<���<�8�<���<�`�<��<Cw�<���<~�<8��<w�<��<�c�<�դ<�E�<g��<�<���<U�<OX�<��<�"�</��<��<:�z<�bs<\)l<��d<ظ]<��V<$NO<�H<Z�@<��9<��2<�q+<7Q$<5<_<<�<�� <}��;��;d1�;/c�;���;���;�a�;�ܓ;�k�;�r;��W;%5=;h#;�	;*s�:�?�:��p:�2:�^!9�j�-����}����{�޺����3�TE5��L�$�b�b�x�����&f���)��̧�M��������ƻ2ѻۻ��仮��S5��� �Ņ��#
�ڲ��2�����:Z �n�$���(�(-�O"1��35��89��1=��A�� E�y�H�~�L�$eP��T���W��n[�r
_��b�;'f�P�i��#m�M�p��t�]fw�Z�z��~������\������🅼�=��5و�ir��^	��E���81��S��Q��`ߓ�zk��7�������������Z��'��������V"������$��z���%��%����$�������"��w���W ��;���=��x���������������������  �  mqN=6�M=��L=�,L=jK=�J=��I=~I=�ZH=��G=��F=�F=NAE=�xD=ͯC=��B=�B=�NA=��@=s�?=%�>=�>=�A==�n<=?�;=O�:=��9=�9=c98=+]7= 6=X�5=��4=��3=M�2=�2=�"1=X60=�G/=�V.=zc-=m,=�t+=�y*=S{)=Wz(=Iv'=Bo&=e%=�W$=	G#=�2"=�!=�  = �=ȿ=ܙ=.p=�B=<=��=��=%e=�#=*�=w�=�F=��=��=PD=��
=E�	=�=��=�B=��=�X=�� =��<���<ث�<q��<�{�<%Y�<~/�<��<���<��<�F�<���<V��<#X�<r��<���<�8�<���<�`�<��<Ew�<���<~�<;��<�v�<��<�c�<�դ<�E�<k��<!�<�<[�<CX�<%��<�"�<)��<��<@�z<�bs<B)l<��d<�]<��V<NO<�H<u�@<�9<	�2<�q+<1Q$<+5<@<<�<�� <_��;��;n1�;Hc�;
��;v��;�a�;�ܓ;�k�;�r;��W;l5=;{#;�	;Cr�:s@�:�p:�2:3`!9*�j�d��k�}������޺v��n3��E5��L�;�b�d�x�����e���)��%̧��L��۬����ƻJѻ<ۻ��仟��05��.� ����$
�²��2������DZ �^�$��(�-�A"1��35��89��1=��A�� E�o�H���L�eP��T���W��n[�|
_��b�J'f�O�i��#m�V�p��t�xfw�>�z��~������\������䟅��=��3و�gr��U	��B���;1��J��Q��Uߓ��k��6�������������b����������d"������$������y%��1���}$�������"��w���T ��3���I��r���������������������  �  kqN=5�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=LAE=�xD=ӯC=��B=�B=�NA=��@=q�?=�>=�>=�A==�n<=<�;=N�:=��9=�9=b98=%]7=%6=W�5=��4=��3=L�2=�2=�"1=[60=�G/=�V.=wc-={m,=�t+=�y*=Z{)=Qz(=Pv'=Ao&=e%=�W$=G#=�2"=�!=�  =��=ɿ=ޙ=+p=�B=<=��=��=#e=�#='�=�=�F=��=��=ND=��
=A�	=�=��=�B=��=�X=�� =��<���<ӫ�<{��<�{�<"Y�<{/�<��<���<t��<�F�<���<^��<X�<j��<���<�8�<���<�`�<��<Aw�<���<~�<9��<w�<��<�c�<�դ<�E�<v��<�<��<X�<AX�<��<#�<*��<��<B�z<�bs<h)l<��d<׸]<��V<NO<�H<_�@<ٿ9<�2<�q+< Q$<75<M<<�<�� <p��;��;r1�;5c�;���;���;�a�;�ܓ;�k�;�r;��W;5=;�#;�	;*s�:@�:��p:@4:�^!9��j���J�}����h�޺���l3�E5��L��b���x����f���)��1̧��L��������ƻѻHۻ��仌��h5��� �����#
�Ѳ��2����	�8Z �_�$���(�3-�E"1��35��89��1=��A�� E�b�H���L�.eP��T���W�o[�q
_��b�0'f�J�i��#m�N�p��t�dfw�Q�z��~�����v\��������=��9و�_r��]	��J���11��J��Q��_ߓ��k��9�������������X��)��������a"������%��x���|%��3����$�������"��|���S ��A���6��z���������������������  �  xqN=-�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=MAE=�xD=ٯC=��B=�B=�NA=��@=x�?= �>=�>=�A==�n<=:�;=U�:=��9=�9=n98="]7='6=P�5=��4=��3=G�2=�2=�"1=^60=�G/=�V.=sc-=m,=�t+=}y*=`{)=Lz(=Sv'=?o&=e%=�W$=G#=3"=!=�  =��=˿=�=(p=�B=2=��=��=%e=�#=%�=��=�F=��=��=QD=��
=<�	=�=��=�B=��=�X=�� =
��<���<ǫ�<���<�{�<7Y�<v/�<���<���<m��<�F�<���<\��<X�<t��<���<�8�< ��<�`�<��<Bw�<���<$~�<,��<w�<��<�c�<�դ<�E�<v��<�<��<G�<XX�<��<�"�<+��<��<N�z<�bs<g)l<w�d<�]<��V<NO<�H<Y�@<�9<�2<�q+<$Q$<35<Z<�<�<�� <���;��;p1�;Cc�;���;���;�a�;�ܓ;�k�;�r;��W;5=;�#;a	;�s�:�?�:��p:�2:�Z!9}{j�Ʊ���}����\�޺����3�UE5�EL�զb���x� �4f���)���˧�4M��z����ƻ�ѻRۻ�����l5��� �����#
�ֲ��2�����Z ���$���(�/-�?"1��35��89��1=��A�� E���H�}�L�eP��T���W�!o[�f
_�*�b�A'f�a�i��#m�E�p��t�Rfw�b�z��~������\�����������=��Dو�`r��\	��@���51��Y��Q��dߓ�vk��8�������������L��,��������^"������%��s����%������$�������"������M ��M���7������������������������  �  qqN=/�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=MAE=�xD=үC=��B=�B=�NA=��@=v�?=!�>=�>=�A==�n<=:�;=U�:=��9=�9=g98="]7=&6=S�5=��4=��3=L�2=�2=�"1=[60=�G/=�V.=tc-=|m,=�t+=y*=]{)=Pz(=Ov'=Bo&=e%=�W$=G#= 3"=�!=�  =��=ǿ=ܙ=)p=�B=7=��=��=$e=�#=)�=}�=�F=��=��=ND=��
=>�	=�=��=�B=��=�X=�� =��<���<̫�<}��<�{�<*Y�<w/�<���<���<q��<�F�<���<`��<X�<t��<���<�8�<���<�`�<��<Bw�<���<&~�<2��<	w�<��<�c�<�դ<�E�<o��<�<��<K�<JX�<��<�"�<,��<��<J�z<�bs<_)l<��d<�]<y�V<NO<�H<X�@<�9<�2<�q+<1Q$<(5<O<<�<�� <���;��;�1�;?c�;���;���;�a�;�ܓ;�k�;�r;ۓW;<5=;�#;�	;%s�:�?�:��p:�2:\!9q�j�Ʊ���}�2��¡޺���t3�JE5��L��b���x�򀇻,f���)�� ̧�#M��������ƻѻ:ۻ��仇��M5��� �΅��#
�ղ��2�����)Z �r�$���(�!-�A"1��35��89��1=��A�� E���H���L�$eP��T���W�o[�q
_��b�;'f�N�i��#m�R�p��t�^fw�b�z��~������\������񟅼�=��:و�]r��Z	��@���11��Q��Q��`ߓ��k��8�������������S��%��������b"�������$��w����%��*����$�������"������O ��<���;��w������Ĝ�������������  �  jqN=6�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=NAE=yD=ӯC=��B=�B=�NA=��@=p�?=#�>=�>=�A==�n<==�;=O�:=��9=�9=_98=+]7="6=Y�5=��4=��3=I�2=2=�"1=X60=�G/=�V.=zc-={m,=�t+=�y*=X{)=Tz(=Mv'=Bo&=e%=�W$=G#=�2"=�!=�  =�=̿=��=2p=�B===��=��=#e=�#=*�={�=�F=��=��=MD=��
=E�	=�=��=�B=��=�X=�� =
��<���<ث�<u��<�{�<Y�<|/�<
��<���<y��<�F�<���<Z��<X�<h��<���<�8�<���<�`�<��<Ow�<���<~�<<��<�v�<��<�c�<�դ<�E�<q��<�<���<\�<>X�<!��< #�<-��<��<3�z<�bs<C)l<��d<ȸ]<��V<'NO<�H<p�@<ҿ9<�2<�q+<,Q$<05<K<<�<�� <a��;��;x1�;Dc�;:��;���;#b�;�ܓ;�k�;�r;s�W;R5=;�#;�	;s�:/@�:5�p:�3:�`!9̉j������}�x��q�޺����3��E5��L�9�b�e�x�����e���)��>̧��L��������ƻ#ѻ;ۻ��仕��Q5��� �����#
�����2������9Z �Z�$���(�)-�H"1��35��89��1=��A�� E�c�H���L�/eP��T���W��n[�{
_��b�T'f�]�i��#m�R�p��t�nfw�?�z��~�����{\������韅��=��6و�cr��Y	��L���41��G��Q��Lߓ��k��,�������������\��$���
�����b"�������$�����x%��7����$�������"��x���[ ��?���I��z���������������������  �  pqN=1�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=NAE=�xD=ͯC=��B=�B=�NA=��@=w�?=$�>=�>=�A==�n<==�;=R�:=��9=�9=e98=(]7= 6=R�5=��4=��3=L�2=�2=�"1=[60=�G/=�V.=vc-=|m,=�t+=�y*=Y{)=Sz(=Ov'=Co&=e%=�W$=G#=3"=�!=�  =��=ſ=ٙ=,p=�B=9=��=��=&e=�#=)�=�=�F=��=��=ND=��
=@�	==��=�B=��=�X=�� =��<���<˫�<r��<�{�<&Y�<v/�<���<���<v��<�F�<���<Y��<%X�<u��<���<�8�<���<�`�<��<>w�<���<!~�<9��<w�<��<�c�<�դ<�E�<p��<�<���<Q�<HX�<��<�"�<!��<��<C�z<�bs<X)l<��d<ܸ]<��V<NO<�H<h�@<�9<��2<�q+<.Q$<-5<X<<�<�� <���;��;x1�;Hc�;���;}��;�a�;�ܓ;�k�;�r;�W;p5=;�#;�	;{s�:.@�:��p:�2:&\!9΃j�E��W�}�F��x�޺���r3�cE5��L��b���x�/���f���)�� ̧�M��������ƻѻ5ۻ���|��>5��� �Å��#
�Ȳ��2�����0Z �h�$���(�-�9"1��35��89��1=��A�� E���H���L�)eP��T���W�o[�q
_��b�A'f�P�i��#m�N�p��t�tfw�I�z��~������\������쟅��=��<و�dr��R	��>���11��L��Q��]ߓ��k��<�������������O��!��������["�������$�������%��,����$�������"��|���S ��:���?��v���������������������  �  rqN=/�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=PAE=�xD=گC=��B=�B=�NA=��@=u�?=�>=�>=�A==�n<=7�;=X�:=��9=�9=i98=]7=(6=V�5=��4=��3=E�2=�2=�"1=Z60=�G/=�V.=tc-=ym,=�t+=y*=`{)=Nz(=Mv'=Eo&=e%=�W$=G#=3"=�!=�  =��=̿=�=,p=�B=3=��=��=!e=�#=*�=~�=�F=��=��=SD=��
==�	=�=��=�B=��=�X=�� =��<���<Ϋ�<���<�{�<+Y�<{/�< ��<���<j��<�F�<���<X��<X�<o��<���<�8�<��<�`�<��<Hw�<���<!~�<.��<w�<��<�c�<�դ<�E�<h��<�<��<L�<NX�<��<#�<-��<��<<�z<�bs<B)l<z�d<׸]<�V< NO<�H<O�@<�9<�2<�q+<6Q$<5<c<�<�<�� <���;��;j1�;Uc�;	��;���;�a�;�ܓ;�k�;�r;̓W;�4=;�#;�	;�s�:u?�:A�p:3:R]!9)�j�O��V�}����ԡ޺����3��E5�L��b���x�倇�%f���)���˧�"M��t��� �ƻ#ѻ"ۻ��代��k5��� �؅��#
�Ʋ��2�����$Z ��$���(�1-�O"1��35��89��1=��A�� E���H�w�L�,eP��T���W�o[�v
_��b�T'f�j�i��#m�W�p��t�Sfw�e�z��~������\�����������=��:و�er��c	��D���51��V��Q��Zߓ�tk��2�������������O��1��������U"������$��s����%��'����$�������"������V ��H���I������������������������  �  pqN=1�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=NAE=�xD=ͯC=��B=�B=�NA=��@=w�?=$�>=�>=�A==�n<==�;=R�:=��9=�9=e98=(]7= 6=R�5=��4=��3=L�2=�2=�"1=[60=�G/=�V.=vc-=|m,=�t+=�y*=Y{)=Sz(=Ov'=Co&=e%=�W$=G#=3"=�!=�  =��=ſ=ٙ=,p=�B=9=��=��=&e=�#=)�=�=�F=��=��=ND=��
=@�	==��=�B=��=�X=�� =��<���<˫�<r��<�{�<&Y�<v/�<���<���<v��<�F�<���<Y��<%X�<u��<���<�8�<���<�`�<��<>w�<���<!~�<9��<w�<��<�c�<�դ<�E�<p��<�<���<Q�<HX�<��<�"�<!��<��<C�z<�bs<X)l<��d<ܸ]<��V<NO<�H<h�@<�9<��2<�q+<.Q$<-5<X<<�<�� <���;��;x1�;Hc�;���;}��;�a�;�ܓ;�k�;�r;�W;p5=;�#;�	;{s�:.@�:��p:�2:"\!9Ӄj�F��X�}�G��y�޺���r3�dE5��L��b���x�/���f���)��!̧�M��������ƻѻ5ۻ���|��>5��� �Å��#
�Ȳ��2�����0Z �h�$���(�-�9"1��35��89��1=��A�� E���H���L�)eP��T���W�o[�q
_��b�A'f�P�i��#m�N�p��t�tfw�I�z��~������\������쟅��=��<و�dr��R	��>���11��L��Q��]ߓ��k��<�������������O��!��������["�������$�������%��,����$�������"��|���S ��:���?��v���������������������  �  jqN=6�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=NAE=yD=ӯC=��B=�B=�NA=��@=p�?=#�>=�>=�A==�n<==�;=O�:=��9=�9=_98=+]7="6=Y�5=��4=��3=I�2=2=�"1=X60=�G/=�V.=zc-={m,=�t+=�y*=X{)=Tz(=Mv'=Bo&=e%=�W$=G#=�2"=�!=�  =�=̿=��=2p=�B===��=��=#e=�#=*�=|�=�F=��=��=MD=��
=E�	=�=��=�B=��=�X=�� =
��<���<ث�<u��<�{�<Y�<|/�<
��<���<y��<�F�<���<Z��<X�<h��<���<�8�<���<�`�<��<Ow�<���<~�<<��<�v�<��<�c�<�դ<�E�<q��<�<���<\�<>X�<!��< #�<-��<��<3�z<�bs<C)l<��d<ȸ]<��V<'NO<�H<p�@<ҿ9<�2<�q+<,Q$<05<K<<�<�� <b��;��;x1�;Dc�;:��;���;#b�;�ܓ;�k�;�r;r�W;Q5=;�#;�	;s�:.@�:3�p:�3:�`!9։j������}�y��r�޺����3��E5��L�:�b�f�x�����e���)��>̧��L��������ƻ$ѻ;ۻ��仕��Q5��� �����#
�����2������9Z �Z�$���(�)-�H"1��35��89��1=��A�� E�c�H���L�/eP��T���W��n[�{
_��b�T'f�]�i��#m�R�p��t�nfw�?�z��~�����{\������韅��=��6و�cr��Y	��L���41��G��Q��Lߓ��k��,�������������\��$���
�����b"�������$�����x%��7����$�������"��x���[ ��?���I��z���������������������  �  qqN=/�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=MAE=�xD=үC=��B=�B=�NA=��@=v�?=!�>=�>=�A==�n<=:�;=U�:=��9=�9=g98="]7=&6=S�5=��4=��3=L�2=�2=�"1=[60=�G/=�V.=tc-=|m,=�t+=y*=]{)=Pz(=Ov'=Bo&=e%=�W$=G#= 3"=�!=�  =��=ǿ=ܙ=)p=�B=7=��=��=$e=�#=)�=}�=�F=��=��=ND=��
=>�	=�=��=�B=��=�X=�� =��<���<̫�<}��<�{�<*Y�<w/�<���<���<q��<�F�<���<`��<X�<t��<���<�8�<���<�`�<��<Bw�<���<&~�<2��<	w�<��<�c�<�դ<�E�<o��<�<��<K�<JX�<��<�"�<,��<��<J�z<�bs<_)l<��d<�]<y�V<NO<�H<X�@<�9<�2<�q+<1Q$<(5<O<<�<�� <���;��;�1�;?c�;���;���;�a�;�ܓ;�k�;�r;ۓW;<5=;�#;�	;$s�:�?�:��p:�2:\!9}�j�ɱ���}�3��ġ޺���u3�KE5��L��b���x�󀇻,f���)�� ̧�$M��������ƻѻ;ۻ��仇��M5��� �΅��#
�ղ��2�����)Z �r�$���(�!-�A"1��35��89��1=��A�� E���H���L�$eP��T���W�o[�q
_��b�;'f�N�i��#m�R�p��t�^fw�b�z��~������\������񟅼�=��:و�]r��Z	��@���11��Q��Q��`ߓ��k��8�������������S��%��������b"�������$��w����%��*����$�������"������O ��<���;��w������Ĝ�������������  �  xqN=-�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=MAE=�xD=ٯC=��B=�B=�NA=��@=x�?= �>=�>=�A==�n<=:�;=U�:=��9=�9=n98="]7='6=P�5=��4=��3=G�2=�2=�"1=^60=�G/=�V.=sc-=m,=�t+=}y*=`{)=Lz(=Sv'=?o&=e%=�W$=G#=3"=!=�  =��=˿=�=(p=�B=2=��=��=%e=�#=%�=��=�F=��=��=QD=��
=<�	=�=��=�B=��=�X=�� =
��<���<ȫ�<���<�{�<7Y�<v/�<���<���<n��<�F�<���<\��<X�<t��<���<�8�< ��<�`�<��<Bw�<���<$~�<,��<w�<��<�c�<�դ<�E�<v��<�<��<G�<XX�<��<�"�<+��<��<N�z<�bs<g)l<w�d<�]<��V<NO<�H<Y�@<�9<�2<�q+<$Q$<35<[<�<�<�� <���;��;p1�;Cc�;���;���;�a�;�ܓ;�k�;�r;��W;5=;�#;a	;�s�:�?�:��p:�2:qZ!9�{j�ʱ���}����^�޺����3�UE5�FL�֦b���x� �4f���)���˧�4M��z����ƻ�ѻRۻ�����l5��� �����#
�ֲ��2�����Z ���$���(�/-�?"1��35��89��1=��A�� E���H�}�L�eP��T���W�!o[�f
_�*�b�A'f�a�i��#m�E�p��t�Rfw�b�z��~������\�����������=��Dو�`r��\	��@���51��Y��Q��dߓ�vk��8�������������L��,��������^"������%��s����%������$�������"������M ��M���7������������������������  �  kqN=5�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=LAE=�xD=ӯC=��B=�B=�NA=��@=q�?=�>=�>=�A==�n<=<�;=N�:=��9=�9=b98=%]7=%6=W�5=��4=��3=L�2=�2=�"1=[60=�G/=�V.=wc-={m,=�t+=�y*=Z{)=Qz(=Pv'=Ao&=e%=�W$=G#=�2"=�!=�  =��=ɿ=ޙ=+p=�B=<=��=��=#e=�#='�=�=�F=��=��=ND=��
=A�	=�=��=�B=��=�X=�� =��<���<ӫ�<{��<�{�<"Y�<{/�<��<���<t��<�F�<���<^��<X�<j��<���<�8�<���<�`�<��<Aw�<���<~�<9��<w�<��<�c�<�դ<�E�<v��<�<��<X�<AX�<��<#�<*��<��<B�z<�bs<h)l<��d<׸]<��V<NO<�H<_�@<ٿ9<�2<�q+< Q$<75<M<<�<�� <q��;��;r1�;5c�;���;���;�a�;�ܓ;�k�;�r;��W;5=;�#;�	;)s�:@�:��p:<4:�^!9�j���N�}����j�޺���m3�E5��L��b���x����f���)��1̧��L��������ƻѻIۻ��仌��i5��� �����#
�Ѳ��2����	�8Z �_�$���(�3-�E"1��35��89��1=��A�� E�b�H���L�.eP��T���W�o[�q
_��b�0'f�J�i��#m�N�p��t�dfw�Q�z��~�����v\��������=��9و�_r��]	��J���11��J��Q��_ߓ��k��9�������������X��)��������a"������%��x���|%��3����$�������"��|���S ��A���6��z���������������������  �  mqN=6�M=��L=�,L=jK=�J=��I=~I=�ZH=��G=��F=�F=NAE=�xD=ͯC=��B=�B=�NA=��@=s�?=%�>=�>=�A==�n<=?�;=O�:=��9=�9=c98=+]7= 6=X�5=��4=��3=M�2=�2=�"1=X60=�G/=�V.=zc-=m,=�t+=�y*=S{)=Wz(=Iv'=Bo&=e%=�W$=	G#=�2"=�!=�  = �=ȿ=ܙ=.p=�B=<=��=��=%e=�#=*�=w�=�F=��=��=PD=��
=E�	=�=��=�B=��=�X=�� =��<���<ث�<q��<�{�<&Y�<~/�<��<���<���<�F�<���<V��<#X�<r��<���<�8�<���<�`�<��<Ew�<���<~�<;��<�v�<��<�c�<�դ<�E�<k��<!�<�<[�<CX�<%��<�"�<)��<��<@�z<�bs<B)l<��d<�]<��V<NO<�H<u�@<�9<	�2<�q+<1Q$<+5<@<<�<�� <_��;��;n1�;Hc�;
��;v��;�a�;�ܓ;�k�;�r;��W;l5=;{#;�	;Br�:q@�:�p:�2:"`!9;�j�h��p�}������޺w��o3��E5��L�<�b�e�x�����e���)��%̧��L��۬����ƻJѻ<ۻ��仟��05��.� ����$
�²��2������DZ �^�$��(�-�A"1��35��89��1=��A�� E�o�H���L�eP��T���W��n[�|
_��b�J'f�O�i��#m�V�p��t�xfw�>�z��~������\������䟅��=��3و�gr��U	��B���;1��J��Q��Uߓ��k��6�������������b����������d"������$������y%��1���}$�������"��w���T ��3���I��r���������������������  �  sqN=2�M=��L=�,L=	jK=�J=��I=|I=�ZH=��G=��F=�F=KAE=�xD=ׯC=��B=�B=�NA=��@=s�?= �>=�>=�A==�n<=:�;=U�:=��9=�9=h98=$]7=&6=W�5=��4=��3=K�2=�2=�"1=Y60=�G/=�V.=uc-=|m,=�t+=�y*=[{)=Qz(=Lv'=Go&=e%=�W$=G#=�2"=�!=�  =��=˿=�=)p=�B=8=��=��=!e=�#=-�=|�=�F=��=��=QD=��
=>�	=�=��=�B=��=�X=�� =��<���<ի�<��<�{�<,Y�<~/�<��<���<t��<�F�<���<T��<X�<p��<���<�8�<���<�`�<��<Cw�<���<~�<8��<w�<��<�c�<�դ<�E�<g��<�<���<U�<OX�<��<�"�</��<��<:�z<�bs<\)l<��d<ظ]<��V<$NO<�H<Z�@<��9<��2<�q+<7Q$<5<_<<�<�� <}��;��;d1�;/c�;���;���;�a�;�ܓ;�k�;�r;��W;$5=;g#;�	;(s�:�?�:��p:�2:�^!9 �j�1����}����}�޺����3�UE5��L�%�b�b�x�����'f���)��̧�M��������ƻ2ѻۻ��仮��S5��� �Ņ��#
�ڲ��2�����:Z �n�$���(�(-�O"1��35��89��1=��A�� E�y�H�~�L�$eP��T���W��n[�r
_��b�;'f�P�i��#m�M�p��t�]fw�Y�z��~������\������🅼�=��5و�ir��^	��E���81��S��Q��`ߓ�zk��7�������������Z��'��������V"������$��z���%��%����$�������"��w���W ��;���=��x���������������������  �  rqN=.�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=OAE=�xD=կC=��B=�B=�NA=��@=p�?=!�>=�>=�A==�n<=7�;=V�:=��9=�9=h98=#]7=,6=P�5=��4=��3=M�2=�2=�"1=a60=�G/=�V.=xc-=}m,=�t+=y*=_{)=Mz(=Sv'=>o&=e%=�W$= G#=3"=�!=�  =��=ſ=ܙ=%p=�B=4=��=~�=(e=�#=$�=��=�F=��=��=QD=��
=@�	=�=��=�B=��=�X=�� =��<ĸ�<ƫ�<���<�{�</Y�<y/�<��<���<l��<�F�<���<c��< X�<h��<���<�8�<���<�`�<��<7w�<���<~�<,��<w�<��<�c�<�դ<�E�<r��<�<��<I�<MX�<��<#�<&��<��<R�z<�bs<t)l<��d<�]<��V<NO<H<Z�@<��9<�2<�q+<2Q$<(5<V<�<�<�� <t��;��;_1�;Hc�;ƥ�;���;�a�;�ܓ;�k�;�r;i�W;15=;#;?	;�s�:d?�:��p:�2:�Z!9��j������}������޺���r3�E5�L���b���x�����	f���)��̧�)M��}���	�ƻ�ѻ\ۻ���d��t5��� �څ��#
����2�����.Z ��$���(�;-�5"1��35��89��1=��A�� E���H���L� eP��T���W�(o[�W
_��b�*'f�F�i��#m�6�p��t�Ifw�]�z��~������\�����������=��Hو�Zr��X	��M���/1��Z��Q��lߓ�k��D�������������V��-���������`"�������$��r����%��(����$�������"�����L ��A���1��z���������������������  �  qqN=4�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=NAE=�xD=ԯC=��B=�B=�NA=��@=p�?= �>=�>=�A==�n<=<�;=S�:=��9=�9=h98=&]7=(6=S�5=��4=��3=K�2=�2=�"1=^60=�G/=�V.=yc-=}m,=�t+=�y*=Z{)=Pz(=Qv'=?o&=e%=�W$= G#=�2"=�!=�  =��=ɿ=ޙ=+p=�B=5=��=�=$e=�#=%�=��=�F=��=��=SD=��
=C�	=�=��=�B=��=�X=�� =��<���<ϫ�<���<�{�</Y�<~/�<��<���<s��<�F�<���<Y��<X�<i��<���<�8�<���<�`�<��<Bw�<���<~�<3��<w�<��<�c�<�դ<�E�<s��<�<���<V�<MX�<��<#�<*��<��<J�z<�bs<V)l<��d<�]<��V<NO<�H<f�@<�9<�2<�q+<(Q$<05<S<�<�<�� <s��;��;F1�;Dc�;���;���;�a�;�ܓ;xk�;�r;s�W;5=;�#;f	;Rs�:�?�:��p:�2:�^!9z�j�۰�b�}�:���޺����3�yE5��L�ܦb���x��f���)��̧�M��������ƻѻ[ۻ��仔��u5��� �҅��#
�ϲ��2�����9Z �z�$���(�5-�F"1��35��89��1=��A�� E�s�H�w�L�eP��T���W�o[�a
_��b�E'f�S�i��#m�=�p��t�Tfw�O�z��~������\������🅼�=��Bو�dr��^	��K���21��Y��Q��^ߓ��k��8�������������X��-��������a"������%��z���~%��(����$�������"��x���O ��=���@��w���������������������  �  oqN=5�M=��L=�,L=jK=�J=��I={I=�ZH=��G=��F=�F=HAE=�xD=ͯC=��B=�B=�NA=��@=t�?="�>=�>=�A==�n<=>�;=S�:=��9=�9=f98=']7=$6=X�5=��4=��3=Q�2=�2=�"1=Z60=�G/=�V.=tc-=}m,=�t+=�y*=Y{)=Tz(=Lv'=Eo&=e%=�W$=	G#=�2"=�!=�  =��=Ŀ=ٙ=)p=�B=<=��=��= e=�#=-�=|�=�F=��=��=PD=��
=A�	=�=��=�B=��=�X=�� =��<���<ګ�<{��<�{�<+Y�<}/�<��<���<{��<�F�<��<P��<X�<u��<���<�8�<���<�`�<��<>w�<���<~�<=��<�v�<��<�c�<�դ<�E�<i��<�<���<X�<HX�<!��<�"�<-��<��<?�z<�bs<Z)l<��d<ݸ]<��V<%NO<�H<h�@<�9<�2<�q+<2Q$<&5<Q<<�<�� <f��;��;j1�;c�;�;x��;�a�;|ܓ;�k�;�r;��W;65=;@#;�	;�r�:B@�:��p:�2:�^!9��j������}������޺v��'3�UE5�RL��b�Y�x�����(f���)��̧��L��������ƻ2ѻ%ۻ������05��#� �����#
�ݲ��2�����BZ �]�$��(�-�U"1��35��89��1=��A�� E�n�H���L�%eP��T���W��n[�r
_��b�6'f�=�i�#m�T�p��t�efw�O�z��~������\������韅��=��0و�nr��\	��@���81��K��Q��cߓ��k��<�������������^����������["������$��}���|%��,����$�������"��s���U ��*���>��g���������������������  �  rqN=0�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=MAE=�xD=үC=��B=�B=�NA=��@=p�?=!�>=�>=�A==�n<==�;=R�:=��9=�9=i98=(]7=*6=W�5=��4=��3=I�2=2=�"1=]60=�G/=�V.=zc-=�m,=�t+=�y*=]{)=Sz(=Nv'=>o&=e%=�W$=G#=�2"=�!=�  =��=ȿ=ݙ=-p=�B=7=��=��="e=�#=%�=~�=�F=��=��=OD=��
=D�	=�=��=�B=��=�X=�� =��<���<ի�<���<�{�<0Y�<z/�<	��<���<x��<�F�<���<X��<X�<l��<���<�8�<���<�`�<��<Cw�<���<~�</��<�v�<��<�c�<�դ<�E�<o��<�<��<P�<JX�<$��<#�<0��<��<E�z<�bs<G)l<��d<�]<��V<(NO<�H<n�@<�9<�2<�q+</Q$<,5<G<<�<�� <J��;��;g1�;;c�;���;���;�a�;�ܓ;�k�;Br;l�W;35=;�#;�	;�r�:@�:��p:|3:�[!9׀j�c����}����b�޺����3��E5��L��b���x������e���)��!̧�M��������ƻ ѻ]ۻ��仡��G5��*� �҅��#
�ʲ��2�����:Z �s�$��(�&-�K"1��35��89��1=��A�� E�t�H���L�eP��T���W�
o[�g
_��b�Q'f�]�i��#m�J�p��t�Nfw�G�z��~�����~\������쟅��=��>و�er��[	��I���A1��S��Q��]ߓ��k��8�������������d��"��������d"�������$��v����%��*���~$�������"��v���R ��:���G��x���������������������  �  �nN=T�M=N�L=�(L=�eK=��J=��I=I=�TH=0�G=��F={F=�9E=�pD=�C=k�B=�B=KDA=�v@=��?=�>=�>=�4==�`<=��;=(�:=�9={9=9(8=NK7=�l6=�5=��4=>�3=��2=T�1=�1=�0=P//=�=.=eI-=�R,=3Y+=]*=(^)=S\(=�W'=�O&=�D%=�6$=V%#=�"=|� =��=��=�=mt=7J=8=X�=��=�z=6==��=ɵ=�k==�=�u=�=Y�
=�Z	=o�=��=K=��=82=ȷ =�r�<�n�<1c�<?P�< 6�<��<���<��<Ɉ�<M�<G�<r��<�u�<�"�<���<1l�<N	�<ʡ�<�5�<-��<�P�<ع<�[�<?ܲ<PY�<4ӫ<hJ�<꾤<1�<頝<��<�z�<r�<�N�<���<��<3��<�<+�z<js<C5l<� e<k�]<��V<|kO<�=H<�A<p�9<��2<Q�+<��$<Xq<�^<�Q<�J<CJ<[��;=��;3��;� �;�k�;�ȯ;+8�;0��;R�;�s;d�Y;�0?;�%; ;,��:��:4�y:�n:	G9�!D�e����s�!����ٺ�K���E�2��mI��_�PCv�b&��?
��p͛��o���𰻴P��0�Ż��ϻ��ٻ;���G�����1 �}����	���Ȕ�5�2m����$�:H(�~v,���0��4�1�8�P�<�٠@�ԅD��_H�+/L��O�ӮS��_W��[�8�^�<b�D�e�|Ni���l��Ap�.�s��w�xz��}������:��3߃�逅� ������W��^h���v��˫��6<��˓�BX���㖼Sn��h���A�����Ӌ������������/�����h���R��Ӟ�����㞭����N���������r���������X���e��֠���"���  �  oN=[�M=K�L=�(L=�eK=�J=��I=I=�TH=&�G=��F=|F=�9E=�pD=�C=p�B=�B=MDA=�v@=�?=�>=�>=�4==�`<=��;=)�:=�9=�9=B(8=OK7=�l6=�5=��4=A�3=��2=H�1=�1=�0=Q//=�=.=cI-=�R,=<Y+=]*=%^)=X\(=�W'=�O&=�D%=�6$=X%#=�"=z� =��=��=�=rt=:J=5=W�=��=�z=6==��=��=�k==	�=�u=�=_�
=�Z	=l�=�=I=��=-2=· =�r�<�n�<9c�<8P�<!6�<��<���<��<Ɉ�<M�<8�<d��<�u�<�"�<���<l�<Q	�<ơ�<�5�<9��<�P�<ع<�[�</ܲ<9Y�<@ӫ<]J�<ݾ�<�0�<ޠ�<��<�z�<�<�N�<���<��<6��<�<1�z<js<5l<� e<u�]<��V<�kO<�=H<�A<��9<
�2<G�+<�$<Lq<�^<�Q<�J<cJ<��;���;:��;� �;�k�;�ȯ;Q8�;&��;*R�;S�s;�Y;,1?;1%;�;/��:��:�y:�n:�G9D�:���s�������ٺ�K�C��	�2�WmI��_�ACv�s&��L
��?͛�=o��u��P���ŻϮϻ׬ٻ|���G���� 2 ������	������#�%m���$�rH(��v,���0�,�4�T�8�s�<�Ơ@�مD��_H�
/L���O�ڮS� `W��[�@�^�<b�o�e��Ni���l��Ap��s��w�~xz���}������:��3߃�倅� ��ɼ��-W��Qp������ɫ��:<���ʓ�6X���㖼Tn��j���P����ǋ������������:�����o���E���������鞭����R������������}������\���]��ݠ���"���  �  �nN=S�M=G�L=�(L=�eK=��J=��I=I=�TH=(�G=��F=F=9E=�pD=�C=l�B=�B=SDA=�v@=�?=�>=�>=�4==�`<=��;=*�:=�9=z9=<(8=NK7=�l6=�5=��4=B�3=��2=J�1=�1=�0=M//=�=.=cI-=�R,=2Y+=]*=!^)=\\(=�W'=�O&=�D%=�6$=\%#=�"=�� =��=��=�=mt=9J=3=`�=��=�z=5==��=̵=�k==�=�u=�=[�
=�Z	=l�=�=A=��=02=Ʒ =�r�<�n�<<c�<8P�<6�<��<���<��<ƈ�<!M�<>�<x��<�u�<�"�<���<l�<a	�<���<�5�<0��<�P�<ع<�[�<?ܲ<:Y�<Eӫ<XJ�<�<1�<ߠ�<��<�z�<r�<�N�<���<��<;��<�<%�z<0js<
5l<� e<i�]<��V<�kO<�=H<�A<}�9<��2<4�+<��$<Kq<�^<�Q<�J<iJ<��;.��;Q��;y �;�k�;�ȯ;38�;��;^R�;��s;/�Y;71?;	%;P ;���:��:��y:im:�G9GD����"�s�R���m�ٺ�K� ���2�mI�W�_�vCv�p&��K
��a͛��o�����P���Ż��ϻ�ٻP���G�����1 �f����	���˔�7�*m����$�iH(�vv,���0��4�%�8�j�<���@��D��_H�3/L��O�ܮS�`W��[�]�^��;b�c�e��Ni���l��Ap��s��w��xz���}������:��6߃� � ������.W��Pl����������A<��˓�?X���㖼Xn��f���@����Ë������������9�����x���R��Ϟ�����螭����]������������w������h���X��ݠ���"���  �  �nN=X�M=R�L=�(L=�eK=��J=��I=I=�TH=,�G=��F=yF=�9E=�pD=�C=m�B=�B=IDA=�v@=�?=�>=�>=�4==�`<=��;=,�:=%�9=9=>(8=NK7=�l6=�5=��4=B�3=��2=K�1=�1=�0=O//=�=.=fI-=�R,=5Y+=]*=,^)=T\(=�W'=�O&=�D%=�6$=V%#=�"=z� =��=��=�=qt=;J=6=V�=��=�z=5==��=õ=�k=
=�=�u=�=]�
=�Z	=p�=��=N=��=.2=�� =�r�<�n�<2c�<CP�< 6�<��<���<*��<Ј�<M�<=�<h��<�u�<�"�<���<!l�<I	�<ɡ�<�5�<8��<�P�<#ع<�[�<9ܲ<FY�<6ӫ<eJ�<ݾ�<�0�<ޠ�<��<�z�<}�<�N�<���<��<4��<�<@�z<	js<#5l<� e<�]<��V<�kO<�=H<�A<��9<��2<c�+<�$<Eq<�^<�Q<�J<NJ<7��;!��;��;� �;�k�;�ȯ;:8�;.��;	R�;��s;,�Y;�0?;�%;�;���:~��:�y:gp:"G9OD�M����s����*�ٺ�K����ڡ2��mI���_�`Cv�V&��:
��\͛�so��d𰻏P��%�Ż��ϻ��ٻs���G�����1 ������	������#� m���$�[H(��v,���0�"�4�G�8�k�<�Ӡ@�ÅD��_H�$/L��O�֮S��_W��[�+�^�<b�m�e��Ni���l��Ap�+�s��w�~xz���}������:��+߃�퀅� ��ļ��#W��[p������Ы��8<��˓�7X���㖼On��n���G����ы������������:�����_���G��͞������������S��������������������Y���c��Ԡ���"���  �  oN=T�M=K�L=�(L=�eK=��J=��I=I=�TH=,�G=��F=~F=�9E=�pD=
�C=h�B=�B=LDA=�v@=�?=
�>=�>=�4==�`<=��;=%�:=�9=|9=A(8=IK7=�l6=�5=��4=B�3=��2=Q�1=�1=�0=G//=�=.=`I-=�R,=8Y+=]*=&^)=R\(=�W'=�O&=�D%=�6$=T%#=�"=y� =��=��=�=pt=5J=>=V�=��=�z=:==��=µ=�k=	=�=�u=�=^�
=�Z	=o�=׉=O=��=42=÷ =�r�<�n�<$c�<FP�<6�<��<���<��<���<M�<N�<_��<�u�<�"�<���<%l�<N	�<ڡ�<�5�<<��<�P�<%ع<�[�<3ܲ<HY�<4ӫ<nJ�<۾�<1�<ꠝ<��<�z�<s�<�N�<���<��</��<�<I�z< js<>5l<� e<��]<��V<ukO<�=H<�A<��9<��2<D�+<҈$<Zq<�^<�Q<K<MJ<8��;��;I��;� �;�k�;�ȯ;8�;n��;"R�;��s;P�Y;�0?;�%;�;���:���:e�y:�m:�
G9�D����>�s�����n�ٺ�K�b��q�2��mI���_��Cv�j&��h
��O͛�Zo�����P��7�Ż{�ϻ��ٻ]���G������1 ������	���Ŕ�*�8m����$�NH(��v,���0��4�K�8�F�<�֠@���D��_H� /L��O��S��_W��[�&�^�<b�R�e��Ni���l��Ap�G�s��w��xz���}������:��;߃�逅�  ��̼��W��Tm������˫��&<��˓�3X��䖼Mn��c���L����Ӌ������������.���%��n���Q�������枭����\����������u���������b���i��ՠ���"���  �  �nN=T�M=L�L=�(L=�eK=��J=��I=I=�TH=+�G=��F=F=�9E=�pD=	�C=i�B=�B=PDA=�v@=�?=�>=�>=�4==�`<=��;=.�:=�9=|9=>(8=IK7=�l6=�5=��4=A�3=��2=K�1=�1=�0=M//=�=.=`I-=�R,=4Y+=]*=(^)=[\(=�W'=�O&=�D%=�6$=Z%#=�"=~� =��=��=�=rt=6J=9=[�=��=�z=5==��=ĵ=�k==�=�u=�=^�
=�Z	=s�=߉=G=��=/2=�� =�r�<�n�<:c�<CP�<6�<��<���<��<Ј�<M�<:�<m��<�u�<�"�<���< l�<Y	�<ʡ�<�5�<<��<�P�<ع<�[�<;ܲ<BY�<Aӫ<YJ�<侤<�0�<ܠ�<��<�z�<s�<�N�<���<��<B��<�<2�z<js<5l<� e<s�]<��V<�kO<�=H<�A<��9<��2<J�+<�$<Fq<�^<�Q<�J<bJ</��;%��;O��;� �;�k�;�ȯ;8�;*��;AR�;��s;I�Y;1?;%;�;���:���:��y:_n:?
G9�D�����s�:���+�ٺ�K�R��ҡ2�umI���_�}Cv�7&��a
��H͛�o���𰻳P���ŻǮϻ��ٻi���G�����1 �v����	������!�4m�����$�]H(�|v,���0�(�4�B�8�p�<���@�ЅD��_H�./L��O��S��_W��[�H�^�<b�f�e��Ni���l��Ap��s��w��xz���}������:��,߃�倅� ������.W��Tl����������6<��˓�3X���㖼Vn��c���D����Ƌ������������<�����m���P��̞�����랭����Z�������������������g���S��ܠ���"���  �  �nN=[�M=H�L=�(L=�eK=��J=��I=I=�TH=%�G=��F=}F=�9E=�pD=�C=s�B=�B=PDA=�v@=�?=�>=�>=�4==�`<=��;=*�:=�9=�9=<(8=RK7=�l6=�5=��4=B�3=��2=F�1=�1=�0=N//=�=.=`I-=�R,=2Y+=]*= ^)=\\(=�W'=�O&=�D%=�6$=^%#=�"=�� =��=��=�=mt=>J=5=^�=��=�z=8==��=ɵ=�k==�=�u=�=^�
=�Z	=i�=�=F=��=+2=�� =�r�<�n�<9c�<2P�<&6�<��<���<��<Ĉ�<%M�<5�<w��<�u�<�"�<���<l�<Y	�<á�<�5�<-��<�P�<"ع<�[�<@ܲ<4Y�<Kӫ<]J�<뾤<�0�<⠝<��<�z�<��<�N�<Ķ�<��<5��<�<,�z<$js<5l<� e<s�]<��V<�kO<�=H<�A<x�9<	�2<:�+<��$<Tq<�^<�Q<�J<yJ<���;/��;>��;� �;�k�;�ȯ;k8�;��;BR�;��s;�Y;r1?;(%;M ;7��:��:��y:tn:�G9�D�T����s�����A�ٺ�K�T���2�AmI��_�gCv��&��e
��;͛��o��U��P���Żîϻ��ٻi���G�x���2 �f����	���Ȕ�6�m�	���$�pH(�sv,���0�*�4�,�8�p�<���@��D��_H�3/L� �O�ޮS�`W��[�K�^��;b�w�e��Ni���l��Ap��s��w�qxz���}������:��7߃�݀�� ������.W��Kr����������=<���ʓ�BX���㖼Pn��l���?������������������6�����w���@��Ҟ�����𞭼���Z������������������e���^��堼��"���  �  �nN=W�M=J�L=�(L=�eK=��J=��I=I=�TH=*�G=��F=|F=�9E=�pD=�C=o�B=�B=ODA=�v@=�?=�>=�>=�4==�`<=��;='�:=�9=}9=:(8=NK7=�l6=�5=��4=?�3=��2=N�1=�1=�0=N//=�=.=bI-=�R,=2Y+=]*="^)=X\(=�W'=�O&=�D%=�6$=W%#=�"=�� =��=��=�=pt=:J=5=]�=��=�z=8==��=Ƶ=�k==�=�u=�=[�
=�Z	=n�=މ=J=��=12=· =�r�<�n�<0c�<<P�<6�<��<���<��<�<&M�<C�<f��<�u�<�"�<���<-l�<V	�<ǡ�<�5�<6��<�P�< ع<�[�<Gܲ<CY�<9ӫ<bJ�<ᾤ<�0�<頝<��<�z�<z�<�N�<���<��<5��<�<1�z< js<,5l<� e<p�]<��V<�kO<�=H<�A<s�9<��2<@�+<�$<`q<�^<�Q<�J<UJ<+��;T��;9��;� �;�k�;�ȯ;O8�;(��;AR�;�s;+�Y;1?;T%;�;���:���:�y:�m:G9� D�i��K�s�������ٺ�K�\����2��mI���_�mCv�h&��V
��U͛��o�����P���Ż��ϻ��ٻq���G�����1 �h����	������(�#m����$�KH(��v,���0�(�4�;�8�V�<���@��D��_H�//L��O��S��_W��[�9�^� <b�^�e��Ni���l��Ap�+�s��w��xz���}������:��9߃�܀�� ��ż��*W��Qo���z��«��9<���ʓ�9X���㖼Rn��l���8��
��΋������������/�����q���J��Ԟ�����螭����Z���������~���������b���`��۠���"���  �  oN=P�M=O�L=�(L=�eK=��J=��I=I=�TH=.�G=��F=F=�9E=�pD=�C=i�B=�B=MDA=�v@=�?=�>=�>=�4==�`<=��;=/�:=�9=z9=C(8=GK7=�l6=�5=��4=B�3=��2=M�1=�1=�0=H//=�=.=`I-=�R,=:Y+=]*=,^)=U\(=�W'=�O&=�D%=�6$=U%#=�"=w� =��=��=�=ut=8J===T�=��=�z=8==��=��=�k=	=�=�u=�=^�
=�Z	=q�=ى=P=��=/2=�� =�r�<�n�<'c�<DP�<6�<��<���<��<Ԉ�<M�<@�<b��<�u�<�"�<���<l�<L	�<֡�<�5�<C��<�P�<$ع<�[�</ܲ<JY�<8ӫ<iJ�<ᾤ<�0�<֠�<��<�z�<j�<�N�<���<��<5��<	�<S�z<�is<.5l<� e<��]<��V<�kO<�=H<�A<��9<��2<W�+<��$<4q<�^<�Q<�J<TJ<H��;���;V��;� �;�k�;�ȯ; 8�;[��;-R�;��s;H�Y;1?;�%;�;���:��:��y:�n:�G9TD���Z�s�}���x�ٺ�K������2��mI�`�_��Cv�O&��^
��M͛�No���𰻋P���ŻŮϻѬٻe���G������1 ������	�������/m����$�TH(��v,���0��4�P�8�i�<�Ԡ@���D��_H�/L���O��S��_W��[� �^�%<b�f�e��Ni���l��Ap�?�s��w��xz���}������:��'߃�򀅼 ��ɼ��W��To������̫��*<��˓�,X���㖼Nn��a���P����ϋ������������B�����c���Z���������枭����`����������|���������e���c��ؠ���"���  �   oN=S�M=J�L=�(L=�eK=��J=��I=I=�TH=-�G=��F=�F=�9E=�pD=�C=l�B=�B=RDA=�v@=��?=�>=�>=�4==�`<=��;=)�:=�9=z9=?(8=IK7=�l6=�5=��4=C�3=��2=L�1=�1=�0=E//=�=.=_I-=�R,=6Y+=]*=$^)=T\(=�W'=�O&=�D%=�6$=\%#=�"=~� =��=��=�=ot=8J=<=\�=��=�z=8==��=˵=�k=
=�=�u=�=Y�
=�Z	=n�=؉=G=��=02=· =�r�<�n�<*c�<@P�<6�<��<���<��<Ĉ�<M�<L�<r��<�u�<�"�<���<$l�<Z	�<ѡ�<�5�<7��<�P�<#ع<�[�<8ܲ<FY�<Cӫ<aJ�<群<1�<㠝<��<�z�<s�<�N�<���<��<6��<�<7�z<js<!5l<� e<z�]<x�V<�kO<�=H<�A<��9<��2<B�+<�$<Iq<�^<�Q<�J<gJ<C��;��;u��;� �;�k�;�ȯ;78�;H��;XR�;��s;��Y;1?;Z%; ;���:ǩ�:w�y:$n:b	G9SD������s����@�ٺ�K�_����2��mI���_��Cv�f&��i
��n͛�ho�����P��$�Ż��ϻs�ٻU���G�����1 �u����	���Ĕ�.�-m�����$�SH(�rv,���0��4�&�8�M�<�Ѡ@��D��_H�&/L��O��S��_W��[�F�^�<b�b�e��Ni���l��Ap�9�s��w��xz���}������:��6߃�쀅�  ������'W��Ud����������/<��˓�8X���㖼Pn��[���H����ċ������������5�����p���Q��ƞ�����Ɬ����g��������������������n���`��٠���"���  �  �nN=\�M=M�L=�(L=�eK=��J=��I=I=�TH=(�G=��F={F=�9E=�pD=�C=v�B=�B=ODA=�v@=�?=�>=�>=�4==�`<=��;=(�:= �9=�9=9(8=PK7=�l6=�5=��4=>�3=��2=H�1=�1=�0=R//=�=.=cI-=�R,=3Y+=]*=$^)=Z\(=�W'=�O&=�D%=�6$=[%#=�"=�� =��=��=�=rt=@J=0=^�=��=�z=5==�=��=�k==�=�u=�=[�
=�Z	=j�=�=D=��=+2=�� =�r�<�n�<7c�<6P�<!6�<��<���<%��<È�<%M�<6�<d��<�u�<�"�<���< l�<W	�<���<�5�<2��<�P�<ع<�[�<Eܲ<;Y�<@ӫ<]J�<ݾ�<�0�<㠝<��<�z�<��<�N�<���<��<5��<�< �z<js<5l<� e<e�]<��V<�kO<�=H<�A<o�9<�2<O�+<�$<Yq<�^<�Q<�J<cJ<��;I��;1��;� �;l�;�ȯ;�8�;��;>R�;��s;P�Y;1?;F%;�;5��:���:L�y:Qo:�G9� D����-�s�����օٺ�K�s�� �2��mI�5�_�#Cv�w&��N
��K͛��o��P��P����Ż��ϻɬٻ}���G�����1 �d����	������ �m����$�fH(�wv,���0�-�4�L�8�o�<���@��D��_H�&/L��O�ܮS�`W��[�R�^�<b�u�e��Ni���l��Ap��s��w�{xz���}������:��7߃�݀�� ��Ǽ��,W��Vj������«��C<���ʓ�=X���㖼Sn��o���:����ǋ������������5�����k���?��֞�����잭����S���
����������������_���^��ߠ���"���  �  �nN=S�M=G�L=�(L=�eK=��J=��I=I=�TH=)�G=��F=�F=�9E=�pD=�C=r�B=�B=SDA=�v@=�?=�>=�>=�4==�`<=��;='�:=�9=z9=<(8=MK7=�l6=�5=��4=@�3=��2=L�1=�1=�0=I//=�=.=`I-=�R,=2Y+=]*=!^)=X\(=�W'=�O&=�D%=�6$=\%#=�"=�� =��=��=�=nt=<J=7=_�=��=�z=:==��=Ƶ=�k==�=�u=�=[�
=�Z	=g�=ډ=F=��=02=÷ =�r�<�n�<'c�<3P�<6�<��<���<��<���<M�<>�<o��<�u�<�"�<���<l�<^	�<ġ�<�5�<.��<�P�<ع<�[�<@ܲ<=Y�<Cӫ<kJ�<<�0�<᠝<��<�z�<p�<�N�<���<��<+��<�<2�z<js<#5l<� e<t�]<��V<qkO<�=H<�A<~�9<��2<4�+<�$<Pq<�^<�Q<K<jJ<!��;2��;`��;� �;�k�;�ȯ;c8�;#��;eR�;��s;I�Y;E1?;�%;% ;���:+��:*�y:m:�G9�D�p��_�s������ٺ�K�;����2�pmI��_��Cv��&��`
��N͛��o�����P���Ż��ϻ��ٻ/���G�����1 �f����	������/�m�����$�eH(�uv,���0��4�8�8�`�<�Š@��D��_H�2/L�
�O��S�`W��[�I�^�<b�b�e��Ni���l��Ap�>�s��w��xz���}������:��:߃�倅� ������W��Nk����������<<���ʓ�AX���㖼Rn��b���?����ċ������������7�����w���T��Ϟ�����힭����^�������������������f���k��⠼��"���  �  oN=X�M=N�L=�(L=�eK=��J=��I=I=�TH=,�G=��F=�F=9E=�pD=�C=n�B=�B=UDA=�v@=��?=�>=�>=�4==�`<=��;=.�:=�9=�9=@(8=GK7=�l6=�5=��4=@�3=��2=F�1=�1=�0=I//=�=.=dI-=�R,=;Y+=]*=)^)=U\(=�W'=�O&=�D%=�6$=\%#=�"=~� =��=��=�=xt=7J=:=\�=��=�z=3==��=µ=�k==�=�u=�=Z�
=�Z	=v�=ډ=H=��=+2=�� =�r�<�n�<.c�<LP�<6�<��<���<!��<ш�<M�<E�<d��<�u�<�"�<���<"l�<^	�<á�<�5�<I��<�P�<ع<�[�<8ܲ<EY�<Aӫ<XJ�<޾�< 1�<ܠ�<��<�z�<{�<�N�<���<��<A��<�<6�z<js<
5l<� e<u�]<��V<�kO<�=H<yA<��9<��2<R�+<��$<>q<�^<�Q<�J<aJ<>��;��;~��; �;�k�;ɯ;F8�;��;oR�;��s;x�Y;1?;2%;�;8��:���:��y:0o:�G9�D����y�s�����хٺ�K�����2��mI���_��Cv�!&��D
��r͛�Co��r𰻥P��!�Ż��ϻ��ٻo��H�����1 �v����	������	�/m�����$�[H(�pv,���0�%�4�H�8�]�<�ؠ@�ɅD��_H�/L��O�߮S��_W��[�?�^�<b�u�e��Ni���l��Ap�.�s��w��xz���}������:��)߃�퀅� ��Ǽ��,W��Yf����������=<��˓�'X���㖼Yn��Y���G����ǋ������������<�����h���I��������➭����b��������������������j���X��Р���"���  �  �nN=S�M=G�L=�(L=�eK=��J=��I=I=�TH=)�G=��F=�F=�9E=�pD=�C=r�B=�B=SDA=�v@=�?=�>=�>=�4==�`<=��;='�:=�9=z9=<(8=MK7=�l6=�5=��4=@�3=��2=L�1=�1=�0=I//=�=.=`I-=�R,=2Y+=]*=!^)=X\(=�W'=�O&=�D%=�6$=\%#=�"=�� =��=��=�=nt=<J=7=_�=��=�z=:==��=Ƶ=�k==�=�u=�=[�
=�Z	=g�=ډ=F=��=02=÷ =�r�<�n�<'c�<3P�<6�<��<���<��<���<M�<>�<o��<�u�<�"�<���<l�<^	�<ġ�<�5�<.��<�P�<ع<�[�<@ܲ<=Y�<Cӫ<kJ�<<�0�<᠝<��<�z�<p�<�N�<���<��<+��<�<2�z<js<#5l<� e<t�]<��V<qkO<�=H<�A<~�9<��2<4�+<�$<Qq<�^<�Q<K<jJ<!��;2��;`��;� �;�k�;�ȯ;c8�;#��;eR�;��s;I�Y;D1?;�%;% ;���:*��:)�y:m:�G9�D�q��`�s������ٺ�K�;����2�pmI��_��Cv��&��`
��N͛��o�����P���Ż��ϻ��ٻ/���G�����1 �f����	������/�m�����$�eH(�uv,���0��4�8�8�`�<�Š@��D��_H�2/L�
�O��S�`W��[�I�^�<b�b�e��Ni���l��Ap�>�s��w��xz���}������:��:߃�倅� ������W��Nk����������<<���ʓ�AX���㖼Rn��b���?����ċ������������7�����w���T��Ϟ�����힭����^�������������������f���k��⠼��"���  �  �nN=\�M=M�L=�(L=�eK=��J=��I=I=�TH=(�G=��F={F=�9E=�pD=�C=v�B=�B=ODA=�v@=�?=�>=�>=�4==�`<=��;=(�:= �9=�9=9(8=PK7=�l6=�5=��4=>�3=��2=H�1=�1=�0=R//=�=.=cI-=�R,=3Y+=]*=$^)=Z\(=�W'=�O&=�D%=�6$=[%#=�"=�� =��=��=�=rt=@J=0=^�=��=�z=5==�=��=�k==�=�u=�=[�
=�Z	=k�=�=D=��=+2=�� =�r�<�n�<7c�<6P�<!6�<��<���<%��<È�<%M�<6�<d��<�u�<�"�<���< l�<W	�<���<�5�<2��<�P�<ع<�[�<Eܲ<;Y�<@ӫ<]J�<ݾ�<�0�<㠝<��<�z�<��<�N�<���<��<5��<�< �z<js<5l<� e<e�]<��V<�kO<�=H<�A<o�9<�2<O�+<�$<Yq<�^<�Q<�J<cJ<��;I��;1��;� �;l�;�ȯ;�8�;��;>R�;��s;P�Y;1?;F%;�;5��:���:J�y:Oo:�G9� D����/�s�����ׅٺ�K�s���2��mI�5�_�#Cv�w&��N
��K͛��o��P��P����Ż��ϻɬٻ}���G�����1 �d����	������ �m����$�fH(�wv,���0�-�4�L�8�o�<���@��D��_H�&/L��O�ܮS�`W��[�R�^�<b�u�e��Ni���l��Ap��s��w�{xz���}������:��7߃�݀�� ��Ǽ��,W��Vj������«��C<���ʓ�=X���㖼Sn��o���:����ǋ������������5�����k���?��֞�����잭����S���
����������������_���^��ߠ���"���  �   oN=S�M=J�L=�(L=�eK=��J=��I=I=�TH=-�G=��F=�F=�9E=�pD=�C=l�B=�B=RDA=�v@=��?=�>=�>=�4==�`<=��;=)�:=�9=z9=?(8=IK7=�l6=�5=��4=C�3=��2=L�1=�1=�0=E//=�=.=_I-=�R,=6Y+=]*=$^)=T\(=�W'=�O&=�D%=�6$=\%#=�"=~� =��=��=�=ot=8J=<=\�=��=�z=8==��=˵=�k=
=�=�u=�=Y�
=�Z	=n�=؉=G=��=02=· =�r�<�n�<*c�<@P�<6�<��<���<��<Ĉ�<M�<M�<r��<�u�<�"�<���<$l�<Z	�<ѡ�<�5�<7��<�P�<#ع<�[�<8ܲ<FY�<Cӫ<aJ�<群<1�<㠝<��<�z�<s�<�N�<���<��<6��<�<7�z<js<!5l<� e<{�]<x�V<�kO<�=H<�A<��9<��2<B�+<�$<Jq<�^<�Q<�J<gJ<C��;��;u��;� �;�k�;�ȯ;78�;H��;XR�;��s;��Y;1?;Z%; ;���:Ʃ�:u�y:"n:Y	G9]D������s����B�ٺ�K�`����2��mI���_��Cv�f&��i
��n͛�ho�����P��%�Ż��ϻs�ٻU���G�����1 �u����	���Ĕ�.�-m�����$�SH(�rv,���0��4�&�8�M�<�Ѡ@��D��_H�&/L��O��S��_W��[�F�^�
<b�b�e��Ni���l��Ap�9�s��w��xz���}������:��6߃�쀅�  ������'W��Ud����������/<��˓�8X���㖼Pn��[���H����ċ������������5�����p���Q��ƞ�����Ɬ����g��������������������n���`��٠���"���  �  oN=P�M=O�L=�(L=�eK=��J=��I=I=�TH=.�G=��F=F=�9E=�pD=�C=i�B=�B=MDA=�v@=�?=�>=�>=�4==�`<=��;=/�:=�9=z9=C(8=GK7=�l6=�5=��4=B�3=��2=M�1=�1=�0=H//=�=.=`I-=�R,=:Y+=]*=,^)=U\(=�W'=�O&=�D%=�6$=U%#=�"=w� =��=��=�=ut=8J===T�=��=�z=8==��=��=�k=	=�=�u=�=^�
=�Z	=q�=ى=P=��=/2=�� =�r�<�n�<'c�<DP�<6�<��<���<��<Ԉ�<M�<@�<b��<�u�<�"�<���<l�<L	�<֡�<�5�<C��<�P�<$ع<�[�</ܲ<JY�<8ӫ<iJ�<ᾤ<�0�<֠�<��<�z�<i�<�N�<���<��<5��<	�<S�z<�is<.5l<� e<��]<��V<�kO<�=H<�A<��9<��2<W�+<��$<4q<�^<�Q<�J<TJ<I��;���;V��;� �;�k�;�ȯ; 8�;[��;-R�;�s;H�Y;1?;�%;�;���:��:��y:�n:�G9_D���]�s�~���y�ٺ�K������2��mI�a�_��Cv�O&��_
��M͛�Oo���𰻌P���ŻŮϻѬٻe���G������1 ������	�������/m����$�TH(��v,���0��4�P�8�i�<�Ԡ@���D��_H�/L���O��S��_W��[� �^�%<b�f�e��Ni���l��Ap�?�s��w��xz���}������:��'߃�򀅼 ��ɼ��W��To������̫��*<��˓�,X���㖼Nn��a���P����ϋ������������B�����c���Z���������枭����`����������|���������e���c��ؠ���"���  �  �nN=W�M=J�L=�(L=�eK=��J=��I=I=�TH=*�G=��F=|F=�9E=�pD=�C=o�B=�B=ODA=�v@=�?=�>=�>=�4==�`<=��;='�:=�9=}9=:(8=NK7=�l6=�5=��4=?�3=��2=N�1=�1=�0=N//=�=.=bI-=�R,=2Y+=]*="^)=X\(=�W'=�O&=�D%=�6$=W%#=�"=�� =��=��=�=pt=:J=5=]�=��=�z=8==��=Ƶ=�k==�=�u=�=[�
=�Z	=n�=މ=J=��=12=· =�r�<�n�<0c�<<P�<6�<��<���<��<�<&M�<C�<g��<�u�<�"�<���<-l�<V	�<ǡ�<�5�<6��<�P�< ع<�[�<Gܲ<CY�<9ӫ<bJ�<ᾤ<�0�<頝<��<�z�<z�<�N�<���<��<5��<�<1�z< js<,5l<� e<p�]<��V<�kO<�=H<�A<s�9<��2<A�+<�$<`q<�^<�Q<�J<UJ<+��;T��;9��;� �;�k�;�ȯ;O8�;(��;AR�;�s;*�Y;1?;T%;�;���:���:�y:�m:G9� D�l��N�s�������ٺ�K�]����2��mI���_�mCv�h&��W
��U͛��o�����P���Ż��ϻ��ٻq���G�����1 �h����	������(�#m����$�KH(��v,���0�(�4�;�8�V�<���@��D��_H�//L��O��S��_W��[�9�^� <b�^�e��Ni���l��Ap�+�s��w��xz���}������:��9߃�܀�� ��ż��*W��Qo���z��«��9<���ʓ�9X���㖼Rn��l���8��
��΋������������/�����q���J��Ԟ�����螭����Z���������~���������b���`��۠���"���  �  �nN=[�M=H�L=�(L=�eK=��J=��I=I=�TH=%�G=��F=}F=�9E=�pD=�C=s�B=�B=PDA=�v@=�?=�>=�>=�4==�`<=��;=)�:=�9=�9=<(8=RK7=�l6=�5=��4=B�3=��2=F�1=�1=�0=N//=�=.=`I-=�R,=2Y+=]*= ^)=\\(=�W'=�O&=�D%=�6$=^%#=�"=�� =��=��=�=mt=>J=5=^�=��=�z=8==��=ɵ=�k==�=�u=�=^�
=�Z	=i�=�=F=��=+2=�� =�r�<�n�<9c�<2P�<&6�<��<���<��<ň�<%M�<5�<w��<�u�<�"�<���<l�<Y	�<á�<�5�<-��<�P�<"ع<�[�<@ܲ<4Y�<Kӫ<]J�<뾤<�0�<⠝<��<�z�<��<�N�<Ķ�<��<5��<�<,�z<$js<5l<� e<s�]<��V<�kO<�=H<�A<x�9<	�2<;�+<��$<Tq<�^<�Q<�J<yJ<���;/��;>��;� �;�k�;�ȯ;k8�;��;BR�;��s;�Y;q1?;'%;L ;6��:~��:��y:qn:�G9�D�X����s�����B�ٺ�K�U���2�BmI��_�hCv��&��f
��;͛��o��U��P���Żîϻ��ٻi���G�x���2 �f����	���Ȕ�6�m�	���$�pH(�sv,���0�*�4�,�8�p�<���@��D��_H�3/L� �O�ޮS�`W��[�K�^��;b�w�e��Ni���l��Ap��s��w�qxz���}������:��7߃�݀�� ������.W��Kr����������=<���ʓ�BX���㖼Pn��l���?������������������6�����w���@��Ҟ�����𞭼���Z������������������e���^��堼��"���  �  �nN=T�M=L�L=�(L=�eK=��J=��I=I=�TH=+�G=��F=F=�9E=�pD=	�C=i�B=�B=PDA=�v@=�?=�>=�>=�4==�`<=��;=.�:=�9=|9=>(8=IK7=�l6=�5=��4=A�3=��2=K�1=�1=�0=M//=�=.=`I-=�R,=4Y+=]*=(^)=[\(=�W'=�O&=�D%=�6$=Z%#=�"=~� =��=��=�=rt=6J=9=[�=��=�z=5==��=ĵ=�k==�=�u=�=^�
=�Z	=s�=��=G=��=/2=�� =�r�<�n�<:c�<CP�<6�<��<���<��<Ј�<M�<:�<m��<�u�<�"�<���< l�<Y	�<ʡ�<�5�<<��<�P�<ع<�[�<;ܲ<BY�<Aӫ<YJ�<侤<�0�<ܠ�<��<�z�<s�<�N�<���<��<B��<�<2�z<js<5l<� e<s�]<��V<�kO<�=H<�A<��9<��2<J�+<�$<Fq<�^<�Q<�J<bJ</��;%��;O��;� �;�k�;�ȯ;8�;*��;AR�;��s;I�Y;1?;%;�;���:���:��y:\n:2
G9�D�����s�<���,�ٺ�K�S��ӡ2�vmI���_�}Cv�8&��a
��H͛�o���𰻳P���ŻȮϻ��ٻi���G�����1 �v����	������!�4m�����$�]H(�|v,���0�(�4�B�8�p�<���@�ЅD��_H�./L��O��S��_W��[�H�^�<b�f�e��Ni���l��Ap��s��w��xz���}������:��,߃�倅� ������.W��Tl����������6<��˓�3X���㖼Vn��c���D����Ƌ������������<�����m���P��̞�����랭����Z�������������������g���S��ܠ���"���  �  oN=T�M=K�L=�(L=�eK=��J=��I=I=�TH=,�G=��F=~F=�9E=�pD=
�C=h�B=�B=LDA=�v@=�?=
�>=�>=�4==�`<=��;=%�:=�9=|9=A(8=IK7=�l6=�5=��4=B�3=��2=Q�1=�1=�0=G//=�=.=`I-=�R,=8Y+=]*=&^)=R\(=�W'=�O&=�D%=�6$=T%#=�"=y� =��=��=�=pt=5J=>=V�=��=�z=:==��=µ=�k=	=�=�u=�=^�
=�Z	=o�=׉=O=��=42=÷ =�r�<�n�<$c�<FP�<6�<��<���<��<���<M�<N�<`��<�u�<�"�<���<%l�<N	�<ڡ�<�5�<<��<�P�<%ع<�[�<3ܲ<HY�<4ӫ<nJ�<۾�<1�<ꠝ<��<�z�<s�<�N�<���<��</��<�<I�z< js<>5l<� e<��]<��V<ukO<�=H<�A<��9<��2<D�+<҈$<Zq<�^<�Q<K<MJ<8��;��;I��;� �;�k�;�ȯ;8�;n��;!R�;��s;O�Y;�0?;�%;�;���:���:b�y:�m:�
G9�D����A�s�����o�ٺ�K�b��r�2��mI���_��Cv�j&��h
��P͛�Zo�����P��7�Ż{�ϻ��ٻ]���G������1 ������	���Ɣ�*�8m����$�NH(��v,���0��4�K�8�F�<�֠@���D��_H� /L��O��S��_W��[�&�^�<b�R�e��Ni���l��Ap�G�s��w��xz���}������:��;߃�逅�  ��̼��W��Tm������˫��&<��˓�3X��䖼Mn��c���L����Ӌ������������.���%��n���Q�������枭����\����������u���������b���i��ՠ���"���  �  �nN=X�M=R�L=�(L=�eK=��J=��I=I=�TH=,�G=��F=yF=�9E=�pD=�C=m�B=�B=IDA=�v@=�?=�>=�>=�4==�`<=��;=,�:=%�9=9=>(8=NK7=�l6=�5=��4=B�3=��2=K�1=�1=�0=O//=�=.=fI-=�R,=5Y+=]*=,^)=T\(=�W'=�O&=�D%=�6$=V%#=�"=z� =��=��=�=qt=<J=6=V�=��=�z=5==��=õ=�k=
=�=�u=�=]�
=�Z	=p�=��=N=��=.2=�� =�r�<�n�<2c�<CP�< 6�<��<���<*��<Ј�<M�<=�<h��<�u�<�"�<���<!l�<I	�<ɡ�<�5�<8��<�P�<#ع<�[�<9ܲ<FY�<6ӫ<eJ�<ݾ�<�0�<ޠ�<��<�z�<}�<�N�<���<��<4��<�<@�z<	js<#5l<� e<�]<��V<�kO<�=H<�A<��9<��2<c�+<�$<Eq<�^<�Q<�J<NJ<7��;!��;��;� �;�k�;�ȯ;:8�;.��;	R�;��s;+�Y;�0?;�%;�;���:}��:�y:ep:G9YD�P����s����+�ٺ�K����ڡ2��mI���_�aCv�W&��:
��\͛�so��d𰻐P��%�Ż��ϻ��ٻs���G�����1 ������	������#� m���$�[H(��v,���0�"�4�G�8�k�<�Ӡ@�ÅD��_H�$/L��O�֮S��_W��[�+�^�<b�m�e��Ni���l��Ap�+�s��w�~xz���}������:��+߃�퀅� ��ļ��#W��[p������Ы��8<��˓�7X���㖼On��n���G����ы������������:�����_���G��͞������������S��������������������Y���c��Ԡ���"���  �  �nN=S�M=G�L=�(L=�eK=��J=��I=I=�TH=(�G=��F=F=9E=�pD=�C=l�B=�B=SDA=�v@=�?=�>=�>=�4==�`<=��;=*�:=�9=z9=<(8=NK7=�l6=�5=��4=B�3=��2=J�1=�1=�0=M//=�=.=cI-=�R,=2Y+=]*=!^)=\\(=�W'=�O&=�D%=�6$=\%#=�"=�� =��=��=�=mt=9J=3=`�=��=�z=5==��=̵=�k==�=�u=�=[�
=�Z	=l�=�=A=��=02=Ʒ =�r�<�n�<<c�<8P�<6�<��<���<��<ƈ�<!M�<>�<x��<�u�<�"�<���<l�<a	�<���<�5�<0��<�P�<ع<�[�<?ܲ<:Y�<Eӫ<XJ�<�<1�<ߠ�<��<�z�<r�<�N�<���<��<;��<�<%�z<0js<
5l<� e<i�]<��V<�kO<�=H<�A<}�9<��2<4�+<��$<Kq<�^<�Q<�J<iJ<��;.��;Q��;y �;�k�;�ȯ;38�;��;^R�;��s;/�Y;71?;	%;O ;���:��:��y:gm:�G9ND����#�s�S���n�ٺ�K� ���2�mI�X�_�vCv�p&��K
��a͛��o�����P���Ż��ϻ�ٻP���G�����1 �f����	���˔�7�*m����$�iH(�vv,���0��4�%�8�j�<���@��D��_H�3/L��O�ܮS�`W��[�]�^��;b�c�e��Ni���l��Ap��s��w��xz���}������:��6߃� � ������.W��Pl����������A<��˓�?X���㖼Xn��f���@����Ë������������9�����x���R��Ϟ�����螭����]������������w������h���X��ݠ���"���  �  oN=[�M=K�L=�(L=�eK=�J=��I=I=�TH=&�G=��F=|F=�9E=�pD=�C=p�B=�B=MDA=�v@=�?=�>=�>=�4==�`<=��;=)�:=�9=�9=B(8=OK7=�l6=�5=��4=A�3=��2=H�1=�1=�0=Q//=�=.=cI-=�R,=<Y+=]*=%^)=X\(=�W'=�O&=�D%=�6$=X%#=�"=z� =��=��=�=rt=:J=5=W�=��=�z=6==��=��=�k==	�=�u=�=_�
=�Z	=l�=�=I=��=-2=· =�r�<�n�<9c�<8P�<!6�<��<���<��<Ɉ�<M�<8�<d��<�u�<�"�<���<l�<Q	�<ơ�<�5�<9��<�P�<ع<�[�</ܲ<8Y�<@ӫ<]J�<ݾ�<�0�<ޠ�<��<�z�<�<�N�<���<��<6��<�<1�z<js<5l<� e<u�]<��V<�kO<�=H<�A<��9<
�2<G�+<�$<Lq<�^<�Q<�J<cJ<��;���;:��;� �;�k�;�ȯ;Q8�;&��;*R�;S�s;�Y;,1?;1%;�;.��:��:~�y:�n:�G9D�;���s�������ٺ�K�C��	�2�XmI��_�ACv�s&��L
��?͛�=o��u��P���ŻϮϻ׬ٻ|���G���� 2 ������	������#�%m���$�rH(��v,���0�,�4�T�8�s�<�Ơ@�مD��_H�
/L���O�ڮS� `W��[�@�^�<b�o�e��Ni���l��Ap��s��w�~xz���}������:��3߃�倅� ��ɼ��-W��Qp������ɫ��:<���ʓ�6X���㖼Tn��j���P����ǋ������������:�����o���E���������鞭����R������������}������\���]��ݠ���"���  �  �lN=��M=K�L=r%L=#bK=[�J=�I=I=�OH=Z�G=o�F=��E=^2E=iD=��C=��B=�B=�:A=�l@=g�?=��>=S�==a(==T<=h~;=J�:=��9=d�8=�8=�:7=�[6=mz5=_�4=H�3=3�2=��1=��0=�0=�/=x&.=�1-=:,=�?+=C*=�C)=�@(=�;'=3&=t'%=�$=�#=X�!=�� =k�=��=Xy=`R=�'=I�=��=�=�V=�=��=�=G=�=�=�P=��=��
=M6	=��=�e=j�=/�==� =�.�<�+�<!�<|�<���<���<=��<���<SO�<?�<(��<��<.C�<���<���<?�<6��<�x�<l�<��<d-�<䶹<�<�<��<%>�<��<P3�<ީ�<�<<���<n�<�ڒ<�E�<���<$�<y��<c�<ءz<�ps<�?l<�e<4�]<p�V<N�O<�\H<�5A<c:<��2<*�+<ʻ$<$�<��<��<��<��<�6�;8Y�;@��;C��; �;̄�;���;��;[$�;o�u;A[;"�@;��&;,	;t��:E��:��:��:�Qi9�,!�R
�>�j�$d���Ժ2���5�B;0�9G��]�!�s�S넻�͏�����a2������9���TĻqtλ!tػ�S���i���K5���K��������z����;���#���'�u�+�K0��04�i;8�a:<��-@��D���G���K�ȌO�wJS���V�B�Z��J^�{�a��se���h��{l�C�o��es���v� 3z�4�}��s��	�������d���������0>���׋��n���������(��d����F��<Ӗ��^��~虼Oq���������/���������B������������񘪼���������y������S�������������⟹��!��ʣ���&���  �  �lN=��M=L�L=s%L=$bK=U�J=��I=I=�OH=Y�G=o�F=��E=Z2E=iD=��C=��B=�B=�:A=�l@=g�?=��>=O�==\(==T<=k~;=K�:=��9=o�8=�8=�:7=�[6=sz5=`�4=Q�3=5�2=��1=��0=�0=�/=w&.=�1-=:,=�?+=(C*=�C)=�@(=�;'=	3&=r'%=�$=�#=S�!=�� =c�=��=Yy=aR=�'=A�=��=��=�V=�=��=�=G=�=�=�P=��=��
=H6	=��=�e=n�=8�==� =�.�<�+�<,!�<r�<���<���<T��<��<SO�<G�<��<���<(C�<���<���<?�<7��<�x�<s�<���<c-�<߶�<�<�<	��<!>�<$��<M3�<ש�<��<폝<���<n�<�ڒ<�E�<ꯋ<�<z��<h�<�z<�ps<�?l<�e<O�]<t�V<U�O<�\H<g5A<l:<��2</�+<һ$<(�<��<��<��< �<�6�;9Y�;1��;#��; �;���;���;慕;U$�;�u;�@[;��@;`�&;�;���:���:��:��:�]i9�-!��
��j��c����Ժ����5��;0��G�ˈ]���s�[넻$Ώ�����;2������O���TĻ�tλTtػ T⻿�:���s5���K��������z����+;���#���'�c�+�20��04��;8�v:<��-@��D���G���K�ԌO��JS���V��Z��J^�V�a��se���h��{l�<�o�xes���v�33z�<�}�us���������}d���������6>��w׋��n���������(��]����F��=Ӗ��^���虼Kq���������1���������D������������옪����������t������C������������������!��ڣ���&���  �  �lN=��M=D�L=s%L=%bK=X�J=�I=I=�OH=S�G=r�F=��E=]2E=iD=�C=��B=�B=�:A=�l@=c�?=��>=M�==f(==T<=m~;=E�:=��9=i�8=�8=�:7=�[6=wz5=W�4=N�3=7�2=��1=��0=�0=�/=v&.=�1-=:,=�?+=$C*=yC)=A(=�;'=3&=w'%=�$=�#=O�!=�� =a�=��=Wy=^R=�'=>�=�=ߐ=�V=�=��=�=G=�=�=�P=��=��
=M6	=��=�e=c�=8�==� =�.�<�+�</!�<p�<���<���<E��<��<CO�<M�<��<��<'C�<���<���<?�<F��<�x�<�<���<g-�<趹<�<�<��<>�<'��<J3�<橤<�<���<���<�m�<�ڒ<�E�<���<�<��<a�<Сz<�ps<�?l<�e<8�]<\�V<c�O<�\H<5A<_:<��2<�+<ϻ$<-�<��<ʐ<��<%�<c6�;JY�;G��;;��;- �;���;���;煕;�$�;2�u;�@[;��@;E�&;x	;��:��:��:$�:�Vi9�.!��
���j��b���Ժ����5��;0��G�|�]���s�d넻�͏�~���n2����������TĻ�tλtػ�S���.����5���K����р�	��z����6;���#���'�^�+�60�}04�c;8�r:<��-@��D���G���K���O�xJS���V�#�Z��J^�X�a��se���h��{l�_�o�pes���v�3z�=�}��s���������vd���������7>��x׋��n���������(��Q����F��9Ӗ��^���虼Bq���������5������A�������������������������|������B�������������쟹��!��գ���&���  �  �lN=��M=P�L=u%L=#bK=S�J=��I=I=�OH=X�G=p�F=��E=^2E=iD=��C=��B=�B=�:A=�l@=i�?=��>=P�==_(==T<=k~;=J�:=��9=g�8=�8=�:7=�[6=tz5=^�4=N�3=3�2= �1=��0=�0=�/=x&.=�1-=:,=�?+=$C*=�C)=�@(=�;'=
3&=r'%=�$=�#=S�!=�� =a�=��=Wy=_R=�'=?�=��=�=�V=�=��=
�=G=�=�=�P=��=��
=H6	=��=�e=l�=3�==� =�.�<�+�<*!�<r�<���<���<C��<��<PO�<F�<��<��<)C�<���<��<?�<6��<�x�<v�<���<d-�<綹<�<�<	��<>�<!��<P3�<ש�<��<菝<���<n�<�ڒ<�E�<���<�<��<i�<ߡz<�ps<�?l<�e<B�]<r�V<^�O<�\H<u5A<i:<��2<?�+<׻$<%�<��<��<��<�<�6�;9Y�;'��;@��; �;���;���;���;X$�;=�u;-A[;��@;j�&;	;:��:���:��:�:SUi9/-!�7
���j�\c��6�Ժ����5�%;0�G��]���s�S넻*Ώ�|���i2������?���TĻ�tλJtػ�S���+���t5���K����݀�	��z����0;���#���'�X�+�?0��04�};8��:<��-@��D���G���K���O��JS���V�'�Z��J^�k�a��se���h��{l�@�o�{es���v�13z�7�}��s���������|d���������5>��~׋��n���������(��Z����F��<Ӗ��^���虼Kq���������/���������H����������������������s������O�������������៹��!��ۣ���&���  �  �lN=��M=K�L=n%L=*bK=\�J=��I=I=�OH=[�G=q�F=��E=`2E=iD=��C=��B=�B=�:A=�l@=i�?=��>=T�==](==T<=o~;=E�:=��9=g�8=�8=�:7=�[6=nz5=]�4=O�3=1�2= �1=��0=�0=�/=~&.=�1-=:,=�?+=!C*=�C)=�@(=�;'=3&=v'%=�$=�#=W�!=�� =h�=��=Xy=aR=�'=G�=��=�=�V=�=��=�=G=�=
�=�P=��=��
=F6	=�=�e=o�=/�==� =�.�<�+�<!�<~�<���<���<E��<��<HO�<J�<)��< ��<0C�<���<��<?�<1��<�x�<m�<��<^-�<趹<�<�<	��<&>�<��<S3�<۩�<�<���<���<n�<�ڒ<�E�<<�<���<\�<�z<�ps<�?l<}e<P�]<^�V<X�O<�\H<e5A<|:<��2<+�+<��$<@�<��<��<��<�<�6�;BY�;9��;O��;��;Ą�;���;!��;M$�;I�u;/A[;\�@;��&;�;���:A��:��:��:�Ui9F(!�%	
���j�d��\�Ժ����5�&;0�PG���]�@�s�$넻9Ώ�����F2������g���TĻZtλ+tػ�S���Q���O5���K���������z����;���#���'�i�+�?0�y04�u;8�Z:<��-@��D���G���K���O��JS���V�F�Z��J^�y�a��se���h��{l�?�o��es���v�<3z�(�}��s���������yd���������/>���׋��n�����!����(��b����F��BӖ��^���虼Jq���������+���������8������
������昪�����������������U�������������럹��!��ף���&���  �  �lN=��M=N�L=s%L="bK=T�J=�I=I=�OH=X�G=q�F=��E=]2E=iD=��C=��B=�B=�:A=�l@=g�?=��>=P�==c(==T<=i~;=I�:=��9=g�8=�8=�:7=�[6=tz5=[�4=P�3=3�2=��1=��0=�0=�/=}&.=�1-=:,=�?+=&C*=�C)= A(=�;'=
3&=w'%=�$=�#=V�!=�� =a�=��=Yy=bR=�'=?�=��=�=�V=�=��=�=G=�=�=�P=��=��
=H6	=��=�e=k�=4�==� =�.�<�+�<(!�<u�<���<���<B��<��<MO�<D�<��<��<)C�<���<��<?�<5��<�x�<u�<��<d-�<涹<�<�<	��<!>�<$��<L3�<㩤<��<ꏝ<���<n�<�ڒ<�E�<���<�<���<Z�<�z<�ps<�?l<�e<I�]<W�V<g�O<�\H<|5A<`:<��2<7�+<ѻ$<�<��<<��<�<�6�;FY�;.��;:��; �;���;���;���;^$�;f�u;A[;��@;p�&;H	;���:r��:g�:5�:TUi9�+!��
���j�Gc����Ժ����5��;0�G���]�7�s�*넻%Ώ�y���u2������^���TĻ�tλKtػ�S���.���V5���K����؀���z����/;���#���'�_�+�>0�|04�z;8�~:<��-@��D���G���K���O��JS���V�<�Z��J^�g�a��se���h��{l�L�o�}es���v�03z�1�}��s���������d���������5>��|׋��n���������(��[����F��=Ӗ��^���虼Jq���������2��򉡼���G��������������������������������M���������������!��֣���&���  �  �lN=��M=H�L=q%L=#bK=U�J=�I=I=�OH=Q�G=r�F=��E=^2E=iD=�C=��B=�B=�:A=�l@=c�?=��>=K�==f(==T<=j~;=F�:=��9=i�8=�8=�:7=�[6=tz5=Y�4=P�3=4�2=��1=��0=�0=�/=x&.=�1-=:,=�?+=)C*=|C)= A(=�;'=3&=t'%=�$=�#=N�!=�� =`�=��=Xy=`R=�'=?�=�=ސ=�V=�=��=�=G=�=�=�P=��=��
=G6	=��=�e=h�=9�==� =�.�<�+�<+!�<i�<���<���<D��<��<FO�<G�<��<��<C�<���<���<?�<;��<�x�<��<���<i-�<궹<�<�<��<>�<.��<G3�<੤<��<ꏝ<���<n�<�ڒ<�E�< ��<�<}��<a�<ڡz<�ps<�?l<�e<@�]<a�V<\�O<{\H<�5A<O:<��2<"�+<ɻ$<%�<��<Đ<��<3�<Y6�;KY�;3��;B��;: �;���;���;���;j$�;:�u;�@[; A;�&;�	;q��:���:�:?�:+Wi9
0!��
���j�Pc����Ժ����5��;0��G�&�]���s�Q넻5Ώ�l����2��u�������TĻ�tλtػ�S���'����5���K����Ȁ���z����1;���#���'�`�+�;0��04�c;8��:<��-@��D���G���K���O��JS���V�/�Z��J^�S�a��se���h��{l�V�o�xes���v�%3z�?�}��s���������|d���������?>��t׋��n���������(��N����F��7Ӗ��^���虼Dq������{��8���������G�������������������������{������D�������������ꟹ��!��䣼��&���  �  �lN=��M=G�L=p%L=%bK=Z�J=��I=I=�OH=Y�G=t�F=��E=`2E=iD=��C=��B=�B=�:A=�l@=h�?=��>=N�==a(==T<=m~;=F�:=��9=k�8=�8=�:7=�[6=pz5=Z�4=M�3=2�2=��1=��0=�0=�/=|&.=�1-=:,=�?+=$C*=~C)=�@(=�;'=3&=t'%=�$=�#=T�!=�� =c�=��=Xy=`R=�'=A�=��=�=�V=�=��=�=G=�=�=�P=��=��
=G6	=��=�e=h�=2�==� =�.�<�+�<!!�<y�<���<���<I��< ��<HO�<I�<��<	��<&C�<���<��<?�<3��<�x�<w�<���<e-�<붹<�<�<��<>�<%��<P3�<۩�<�<<���<n�<�ڒ<�E�<���<�<���<^�<ۡz<�ps<�?l<�e<?�]<]�V<]�O<�\H<v5A<^:<��2<�+<û$<,�<��<��<��<!�<�6�;aY�;(��;P��;( �;���;���;��;J$�;�u;"A[;��@;W�&;3	;(��: ��:#�:D�:*Yi9�-!��
� �j��c����Ժ����5�F;0�G�0�]�0�s�/넻'Ώ�����j2������z���TĻ�tλtػ�S���3���f5���K����Ѐ���z����';���#���'�_�+�30��04�e;8�r:<��-@��D���G���K�ČO��JS���V�D�Z��J^�m�a��se���h��{l�Q�o��es���v�-3z�<�}��s���������yd���������8>��x׋��n���������(��Y����F��;Ӗ��^���虼Aq���������/���������B������������󘪼���������~������N�������������쟹��!��٣���&���  �  �lN=��M=O�L=x%L= bK=W�J=��I=I=�OH=Y�G=p�F=��E=a2E=iD=��C=��B=�B=�:A=�l@=g�?=��>=V�==](==T<=f~;=N�:=��9=h�8=�8=�:7=�[6=oz5=^�4=M�3=0�2=��1=��0=�0=�/=z&.=�1-=:,=�?+="C*=�C)= A(=�;'=3&=u'%=�$=�#=Y�!=�� =g�=��=Xy=bR=�'=F�=��=�=�V=�=��=
�=G=�=�=�P=��=��
=E6	=��=�e=p�=/�==� =�.�<�+�<!�<{�<���<���<F��<��<WO�<=�<��<���<3C�<���<���<?�<2��<�x�<m�<��<`-�<붹<�<�<��<#>�<��<Y3�<ک�<��<珝<���<n�<�ڒ<�E�<鯋<�<��<[�<�z<�ps<�?l<{e<K�]<^�V<Y�O<�\H<]5A<n:<��2<=�+<�$<�<��<��<̍<	�<�6�;;Y�;7��;\��; �;΄�;���;(��;Q$�;u�u;A[;��@;��&;�;���:&��:�:�:QVi9�*!��	
���j��c��-�Ժ����5�0;0�KG���]�P�s�>넻*Ώ�����U2������0���TĻ�tλAtػ�S⻸�F���B5���K����߀���z����;���#���'�g�+�50�x04�};8�|:<��-@��D���G���K�ȌO��JS���V�J�Z��J^�x�a��se���h��{l�:�o��es���v�A3z�4�}��s����������d���������*>��~׋��n���������(��c����F��@Ӗ��^���虼Mq���������&���������I������ ������옪�����������������X�������������럹��!��ң���&���  �  �lN=��M=F�L=r%L='bK=\�J=��I=I=�OH=W�G=r�F=��E=^2E=iD=��C=��B=�B=�:A=�l@=f�?=��>=Q�==_(==T<=l~;=E�:=��9=e�8=�8=�:7=�[6=pz5=Y�4=N�3=2�2=��1=��0=�0=�/=y&.=�1-=:,=�?+=!C*={C)=�@(=�;'=3&=t'%=�$=�#=R�!=�� =f�=��=[y=cR=�'=C�=�=��=�V=�=��=�=G=�=�=�P=��=��
=I6	=��=�e=h�=2�==� =�.�<�+�<#!�<q�<���<���<>��<��<DO�<G�<&��<��<*C�<���< ��<?�<B��<�x�<s�<��<d-�<涹<�<�<��<>�<$��<O3�<۩�<�<�<���< n�<�ڒ<�E�<�<�<}��<\�<ܡz<�ps<�?l<�e<A�]<Z�V<U�O<�\H<n5A<d:<��2<�+<ʻ$<3�<��<��<��<�<�6�;OY�;W��;B��; �;ӄ�;���;��;�$�;K�u;A[;��@;��&;	;���:ݮ�:��:T�:�Si9,!�B
���j��c����Ժ����5�z;0�G��]��s�I넻Ώ�����k2����������TĻytλ#tػ�S���5���y5���K����܀����z����;���#���'�`�+�90��04�n;8�g:<��-@��D���G���K�ǌO��JS���V�=�Z��J^�m�a��se���h��{l�T�o��es���v�.3z�6�}��s���������|d���������4>��y׋��n���������(��\����F��;Ӗ��^��~虼Dq���������0���������?������������򘪼���������������O�������������ퟹ��!��أ���&���  �  �lN=��M=K�L=s%L=$bK=Q�J= �I=I=�OH=Y�G=t�F=��E=\2E=iD=�C=��B=�B=�:A=�l@=l�?=��>=O�==b(==T<=n~;=I�:=��9=l�8=�8=�:7=�[6=uz5=[�4=O�3=3�2=��1=��0=�0=�/=w&.=�1-=:,=�?+=(C*=�C)=A(=�;'=
3&=u'%=�$=�#=Q�!=�� =]�=��=Zy=`R=�'=:�=�=ߐ=�V=�=��=
�=G=�=�=�P=��=��
=G6	=��=�e=f�=6�==� =�.�<�+�</!�<i�<���<���<H��<��<MO�<N�<��<��<(C�<���<��<?�<@��<�x�<��<���<n-�<涹<�<�<��<>�<,��<K3�<ީ�<��<ꏝ<���<n�<�ڒ<�E�<���<�<|��<i�<֡z<�ps<�?l<�e<=�]<l�V<Z�O<�\H<�5A<T:<��2<.�+<ѻ$<)�<��<��<��<(�<�6�;`Y�;+��;3��;K �;���;���;ޅ�;p$�;<�u;YA[;��@;h�&;:	;���:+��:��:��:�Zi97.!��
���j�c����Ժ����5��;0��G�N�]���s�T넻3Ώ�w���n2��|���h���TĻ�tλKtػ�S���	����5���K����̀����z����E;���#���'�I�+�<0��04�{;8��:<��-@��D���G���K���O��JS���V��Z��J^�\�a��se���h��{l�P�o�oes���v�.3z�7�}�s���������ud���������6>��z׋��n���������(��P����F��2Ӗ��^���虼>q������~��3��������G������
�������������������s������F�������������䟹��!��᣼��&���  �  �lN=��M=H�L=r%L=&bK=X�J=�I=I=�OH=W�G=p�F=��E=a2E=iD=�C=��B=�B=�:A=�l@=h�?=��>=T�==f(==T<=k~;=H�:=��9=f�8=�8=�:7=�[6=pz5=[�4=J�3=3�2=��1=��0=�0=�/=w&.=�1-=:,=�?+=C*=C)=�@(=�;'=3&=|'%=�$=�#=R�!=�� =g�=��=Wy=^R=�'=D�=�=�=�V=�=�=�=G=�=
�=�P=��=��
=F6	=��=�e=i�=0�==� =�.�<�+�<!!�<s�<���<���<=��<���<JO�<F�<!��<��<3C�<���<��<?�<E��<�x�<��<���<k-�<�<�<�<��<>�<��<O3�<멤<�<�<���<n�<�ڒ<�E�<���<�<z��<]�<ӡz<�ps<�?l<�e<3�]<\�V<S�O<�\H<{5A<^:<��2<!�+<˻$<0�<��<ϐ<��<�<�6�;;Y�;_��;\��;> �;���;���;&��;�$�;$�u;A[;b�@;��&;�	;.��:ɮ�:`�:��:wTi9�,!�
�'�j��c����Ժ���5�r;0�G�4�]��s�Z넻0Ώ�u���u2��ĳ��j���TĻltλtػ�S���5���v5���K����ʀ���z����;���#���'�^�+�K0�d04�h;8�e:<��-@��D���G���K���O��JS���V�=�Z��J^�s�a��se���h��{l�K�o��es���v�23z�0�}��s���������|d���������*>���׋��n���������(��N����F��4Ӗ�^��z虼Hq���������0��ꉡ����>��������������������������������R�������������쟹��!��ף���&���  �  �lN=��M=O�L=q%L=%bK=U�J=��I=I=�OH=_�G=m�F=��E=Y2E=iD=��C=��B=�B=�:A=�l@=n�?=��>=Q�==W(==T<=f~;=I�:=��9=i�8=�8=�:7=�[6=nz5=`�4=K�3=3�2=��1=��0=�0=�/=|&.=�1-=:,=�?+=%C*=�C)=�@(=�;'=3&=r'%=�$=�#=V�!=�� =e�=��=[y=dR=�'=B�=��=�=�V=�=��=�=G=�=�=�P=��=��
=B6	= �=�e=q�=-�==� =�.�<�+�<!�<|�<���<���<B��<��<QO�<>�<%��<���<+C�<���<��<?�<8��<�x�<q�<��<c-�<۶�<�<�<��<+>�<*��<N3�<ө�<��<���<���<n�<�ڒ<�E�<ᯋ<�<���<^�<�z<�ps<�?l<�e<G�]<d�V<Y�O<�\H<P5A<r:<��2<;�+<ǻ$<*�<��<��<��<(�<�6�;*Y�;]��;��; �;���;���;���;n$�;#�u;~A[;��@;~�&;�;\��:1��:��:�:[Wi9�,!�_

���j�d����Ժ����5�R;0�ZG���]�!�s�-넻<Ώ�����Y2������6���TĻhtλ�tػ�S������Y5���K���������z����%;���#���'�J�+�@0��04��;8�]:<��-@��D���G���K�֌O��JS���V�B�Z��J^���a��se���h��{l�1�o��es���v�N3z�6�}��s����������d���������2>��z׋��n���������(��_����F��<Ӗ��^��{虼Qq���������0�������@������������옪����������~������V�������������蟹��!��գ���&���  �  �lN=��M=H�L=r%L=&bK=X�J=�I=I=�OH=W�G=p�F=��E=a2E=iD=�C=��B=�B=�:A=�l@=h�?=��>=T�==f(==T<=k~;=H�:=��9=f�8=�8=�:7=�[6=pz5=[�4=J�3=3�2=��1=��0=�0=�/=w&.=�1-=:,=�?+=C*=C)=�@(=�;'=3&=|'%=�$=�#=R�!=�� =g�=��=Wy=^R=�'=D�=�=�=�V=�=�=�=G=�=
�=�P=��=��
=F6	=��=�e=i�=0�==� =�.�<�+�<!!�<s�<���<���<=��<���<JO�<F�<!��<��<3C�<���<��<?�<E��<�x�<��<���<k-�<�<�<�<��<>�<��<O3�<멤<�<�<���<n�<�ڒ<�E�<���<�<z��<]�<ӡz<�ps<�?l<�e<3�]<\�V<S�O<�\H<{5A<^:<��2<!�+<˻$<0�<��<ϐ<��<�<�6�;;Y�;_��;\��;> �;���;���;&��;�$�;$�u;A[;a�@;��&;�	;.��:Ȯ�:`�:��:uTi9�,!�
�(�j��c����Ժ���5�r;0�G�4�]��s�Z넻0Ώ�u���u2��ĳ��j���TĻltλtػ�S���5���v5���K����ʀ���z����;���#���'�^�+�K0�d04�h;8�e:<��-@��D���G���K���O��JS���V�=�Z��J^�s�a��se���h��{l�K�o��es���v�23z�0�}��s���������|d���������*>���׋��n���������(��N����F��4Ӗ�^��z虼Hq���������0��ꉡ����>��������������������������������R�������������쟹��!��ף���&���  �  �lN=��M=K�L=s%L=$bK=Q�J= �I=I=�OH=Y�G=t�F=��E=\2E=iD=�C=��B=�B=�:A=�l@=l�?=��>=O�==b(==T<=n~;=I�:=��9=l�8=�8=�:7=�[6=uz5=[�4=O�3=3�2=��1=��0=�0=�/=w&.=�1-=:,=�?+=(C*=�C)=A(=�;'=
3&=u'%=�$=�#=Q�!=�� =]�=��=Zy=`R=�'=:�=�=ߐ=�V=�=��=
�=G=�=�=�P=��=��
=G6	=��=�e=f�=6�==� =�.�<�+�</!�<i�<���<���<I��<��<MO�<N�<��<��<(C�<���<��<?�<@��<�x�<��<���<n-�<涹<�<�<��<>�<,��<K3�<ީ�<��<ꏝ<���<n�<�ڒ<�E�<���<�<|��<i�<֡z<�ps<�?l<�e<=�]<l�V<Z�O<�\H<�5A<T:<��2<.�+<ѻ$<*�<��<��<��<(�<�6�;`Y�;+��;3��;K �;���;���;ޅ�;p$�;<�u;YA[;��@;h�&;:	;���:*��:�:��:�Zi9<.!��
���j�c����Ժ����5��;0��G�N�]���s�T넻3Ώ�w���n2��|���h���TĻ�tλKtػ�S���	����5���K����̀����z����E;���#���'�I�+�<0��04�{;8��:<��-@��D���G���K���O��JS���V��Z��J^�\�a��se���h��{l�P�o�oes���v�.3z�7�}�s���������ud���������6>��z׋��n���������(��P����F��2Ӗ��^���虼>q������~��3��������G������
�������������������s������F�������������䟹��!��᣼��&���  �  �lN=��M=F�L=r%L='bK=\�J=��I=I=�OH=W�G=r�F=��E=^2E=iD=��C=��B=�B=�:A=�l@=f�?=��>=Q�==_(==T<=l~;=E�:=��9=e�8=�8=�:7=�[6=pz5=Y�4=N�3=2�2=��1=��0=�0=�/=y&.=�1-=:,=�?+=!C*={C)=�@(=�;'=3&=t'%=�$=�#=R�!=�� =f�=��=[y=cR=�'=C�=�=��=�V=�=��=�=G=�=�=�P=��=��
=I6	=��=�e=h�=2�==� =�.�<�+�<#!�<q�<���<���<>��<��<DO�<G�<&��<��<*C�<���< ��<?�<B��<�x�<s�<��<d-�<涹<�<�<��<>�<#��<O3�<۩�<�<�<���< n�<�ڒ<�E�<�<�<}��<\�<ܡz<�ps<�?l<�e<A�]<Z�V<U�O<�\H<n5A<d:<��2<�+<ʻ$<3�<��<��<��<�<�6�;OY�;W��;B��; �;҄�;���;��;�$�;J�u;A[;��@;��&;	;���:ܮ�:��:R�:�Si9
,!�C
���j��c����Ժ����5�{;0�G��]��s�I넻Ώ�����k2����������TĻztλ#tػ�S���5���y5���K����܀����z����;���#���'�`�+�90��04�n;8�g:<��-@��D���G���K�ǌO��JS���V�=�Z��J^�m�a��se���h��{l�T�o��es���v�.3z�6�}��s���������|d���������4>��y׋��n���������(��\����F��;Ӗ��^��~虼Dq���������0���������?������������򘪼���������������O�������������ퟹ��!��أ���&���  �  �lN=��M=O�L=x%L= bK=W�J=��I=I=�OH=Y�G=p�F=��E=a2E=iD=��C=��B=�B=�:A=�l@=g�?=��>=V�==](==T<=f~;=N�:=��9=h�8=�8=�:7=�[6=oz5=^�4=M�3=0�2=��1=��0=�0=�/=z&.=�1-=:,=�?+="C*=�C)= A(=�;'=3&=u'%=�$=�#=Y�!=�� =g�=��=Xy=bR=�'=F�=��=�=�V=�=��=
�=G=�=�=�P=��=��
=E6	=��=�e=p�=/�==� =�.�<�+�<!�<{�<���<���<F��<��<XO�<=�<��<���<3C�<���<���<?�<3��<�x�<m�<��<`-�<붹<�<�<��<#>�<��<Y3�<ک�<��<珝<���<n�<�ڒ<�E�<鯋<�<��<[�<�z<�ps<�?l<{e<K�]<^�V<Y�O<�\H<]5A<n:<��2<>�+<�$<�<��<��<̍<	�<�6�;;Y�;8��;\��; �;΄�;���;(��;Q$�;u�u;A[;��@;��&;�;���:%��:�:�:IVi9�*!��	
���j��c��.�Ժ����5�0;0�LG���]�Q�s�>넻*Ώ�����V2������0���TĻ�tλAtػ�S⻸�F���B5���K����߀���z����;���#���'�g�+�50�x04�};8�|:<��-@��D���G���K�ȌO��JS���V�J�Z��J^�y�a��se���h��{l�:�o��es���v�A3z�4�}��s����������d���������*>��~׋��n���������(��c����F��@Ӗ��^���虼Mq���������&���������I������ ������옪�����������������X�������������럹��!��ң���&���  �  �lN=��M=G�L=p%L=%bK=Z�J=��I=I=�OH=Y�G=t�F=��E=`2E=iD=��C=��B=�B=�:A=�l@=h�?=��>=N�==a(==T<=m~;=F�:=��9=k�8=�8=�:7=�[6=pz5=Z�4=M�3=2�2=��1=��0=�0=�/=|&.=�1-=:,=�?+=$C*=~C)=�@(=�;'=3&=t'%=�$=�#=T�!=�� =c�=��=Xy=`R=�'=A�=��=�=�V=�=��=�=G=�=�=�P=��=��
=G6	=��=�e=h�=2�==� =�.�<�+�<!!�<y�<���<���<I��< ��<HO�<I�<��<	��<&C�<���<��<?�<3��<�x�<w�<���<e-�<붹<�<�<��<>�<%��<P3�<۩�<�<<���<n�<�ڒ<�E�<���<�<���<^�<ۡz<�ps<�?l<�e<?�]<]�V<]�O<�\H<v5A<^:<��2<�+<û$<-�<��<��<��<!�<�6�;aY�;(��;P��;( �;���;���;��;J$�;�u;!A[;��@;V�&;2	;'��:���:!�:B�: Yi9�-!�
�"�j��c����Ժ����5�G;0�G�1�]�1�s�0넻'Ώ�����j2������z���TĻ�tλtػ�S���4���f5���K����Ѐ���z����';���#���'�_�+�30��04�e;8�r:<��-@��D���G���K�ČO��JS���V�D�Z��J^�m�a��se���h��{l�Q�o��es���v�-3z�<�}��s���������yd���������8>��x׋��n���������(��Y����F��;Ӗ��^���虼Aq���������/���������B������������󘪼���������~������N�������������쟹��!��٣���&���  �  �lN=��M=H�L=q%L=#bK=U�J=�I=I=�OH=Q�G=r�F=��E=^2E=iD=�C=��B=�B=�:A=�l@=c�?=��>=K�==f(==T<=j~;=F�:=��9=i�8=�8=�:7=�[6=tz5=Y�4=P�3=4�2=��1=��0=�0=�/=x&.=�1-=:,=�?+=)C*=|C)= A(=�;'=3&=t'%=�$=�#=N�!=�� =`�=��=Xy=`R=�'=?�=�=ސ=�V=�=��=�=G=�=�=�P=��=��
=G6	=��=�e=h�=9�==� =�.�<�+�<+!�<i�<���<���<D��<��<FO�<G�<��<��<C�<���<���<?�<;��<�x�<��<���<i-�<궹<�<�<��<>�<.��<G3�<੤<��<ꏝ<���<n�<�ڒ<�E�< ��<�<}��<a�<ڡz<�ps<�?l<�e<@�]<a�V<\�O<{\H<�5A<O:<��2<"�+<ɻ$<%�<��<Đ<��<4�<Y6�;KY�;3��;B��;: �;���;���;���;j$�;:�u;�@[; A;�&;�	;p��:���:�:<�:"Wi90!��
���j�Qc����Ժ����5��;0��G�'�]���s�R넻5Ώ�l����2��u�������TĻ�tλtػ�S���'����5���K����Ȁ���z����1;���#���'�`�+�;0��04�c;8��:<��-@��D���G���K���O��JS���V�/�Z��J^�S�a��se���h��{l�V�o�xes���v�%3z�?�}��s���������|d���������?>��t׋��n���������(��N����F��7Ӗ��^���虼Dq������{��8���������G�������������������������{������D�������������ꟹ��!��䣼��&���  �  �lN=��M=N�L=s%L="bK=T�J=�I=I=�OH=X�G=q�F=��E=]2E=iD=��C=��B=�B=�:A=�l@=g�?=��>=P�==c(==T<=i~;=I�:=��9=g�8=�8=�:7=�[6=tz5=[�4=P�3=3�2=��1=��0=�0=�/=}&.=�1-=:,=�?+=&C*=�C)= A(=�;'=
3&=w'%=�$=�#=V�!=�� =a�=��=Yy=bR=�'=?�=��=�=�V=�=��=�=G=�=�=�P=��=��
=H6	=��=�e=k�=4�==� =�.�<�+�<(!�<u�<���<���<B��<��<NO�<D�<��<��<)C�<���<��<?�<5��<�x�<u�<��<d-�<涹<�<�<	��<!>�<$��<L3�<㩤<��<ꏝ<���<n�<�ڒ<�E�<���<�<���<Y�<�z<�ps<�?l<�e<J�]<W�V<g�O<�\H<|5A<`:<��2<7�+<ѻ$<�<��<<��<�<�6�;FY�;.��;:��; �;���;���;���;^$�;f�u;A[;��@;p�&;H	;���:q��:f�:3�:JUi9�+!��
���j�Hc����Ժ����5��;0�G���]�8�s�+넻%Ώ�y���u2������^���TĻ�tλKtػ�S���/���W5���K����؀���z����/;���#���'�_�+�>0�|04�z;8�:<��-@��D���G���K���O��JS���V�<�Z��J^�g�a��se���h��{l�L�o�}es���v�03z�1�}��s���������d���������5>��|׋��n���������(��[����F��=Ӗ��^���虼Jq���������2��򉡼���F��������������������������������M���������������!��֣���&���  �  �lN=��M=K�L=n%L=*bK=\�J=��I=I=�OH=[�G=q�F=��E=`2E=iD=��C=��B=�B=�:A=�l@=i�?=��>=T�==](==T<=o~;=E�:=��9=g�8=�8=�:7=�[6=nz5=]�4=O�3=1�2= �1=��0=�0=�/=~&.=�1-=:,=�?+=!C*=�C)=�@(=�;'=3&=v'%=�$=�#=W�!=�� =h�=��=Xy=aR=�'=G�=��=�=�V=�=��=�=G=�=
�=�P=��=��
=F6	=�=�e=o�=/�==� =�.�<�+�<!�<~�<���<���<E��<��<HO�<J�<)��< ��<0C�<���<��<?�<1��<�x�<m�<��<^-�<趹<�<�<	��<&>�<��<S3�<۩�<�<���<���<n�<�ڒ<�E�<<�<���<\�<�z<�ps<�?l<}e<Q�]<^�V<X�O<�\H<e5A<|:<��2<+�+<��$<@�<��<��<��<�<�6�;BY�;9��;O��;��;Ą�;���;!��;M$�;H�u;.A[;\�@;��&;�;���:@��:��:��:�Ui9O(!�(	
���j�d��]�Ժ����5�';0�QG���]�A�s�$넻9Ώ�����G2������h���TĻZtλ+tػ�S���Q���O5���K���������z����;���#���'�i�+�?0�y04�u;8�Z:<��-@��D���G���K���O��JS���V�F�Z��J^�y�a��se���h��{l�?�o��es���v�<3z�(�}��s���������yd���������/>���׋��n�����!����(��b����F��BӖ��^���虼Jq���������+���������8������
������昪�����������������U�������������럹��!��ף���&���  �  �lN=��M=P�L=u%L=#bK=S�J=��I=I=�OH=X�G=p�F=��E=^2E=iD=��C=��B=�B=�:A=�l@=i�?=��>=P�==_(==T<=k~;=J�:=��9=g�8=�8=�:7=�[6=tz5=^�4=N�3=3�2= �1=��0=�0=�/=x&.=�1-=:,=�?+=$C*=�C)=�@(=�;'=
3&=r'%=�$=�#=S�!=�� =a�=��=Wy=_R=�'=?�=��=�=�V=�=��=
�=G=�=�=�P=��=��
=H6	=��=�e=l�=3�==� =�.�<�+�<*!�<r�<���<���<C��<��<QO�<F�<��<��<)C�<���<��<?�<6��<�x�<v�<���<d-�<綹<�<�<	��<>�<!��<P3�<ש�<��<菝<���<n�<�ڒ<�E�<���<�<��<i�<ߡz<�ps<�?l<�e<B�]<r�V<^�O<�\H<u5A<i:<��2<?�+<׻$<%�<��<��<��<�<�6�;9Y�;'��;@��; �;���;���;���;X$�;=�u;-A[;��@;j�&;	;9��:���:��:�:LUi97-!�9
���j�]c��7�Ժ����5�%;0�G��]���s�S넻*Ώ�|���i2������?���TĻ�tλKtػ�S���+���t5���K����݀�	��z����0;���#���'�X�+�?0��04�};8��:<��-@��D���G���K���O��JS���V�'�Z��J^�k�a��se���h��{l�@�o�{es���v�13z�7�}��s���������|d���������5>��~׋��n���������(��Z����F��<Ӗ��^���虼Kq���������/���������H����������������������s������O�������������៹��!��ۣ���&���  �  �lN=��M=D�L=s%L=%bK=X�J=�I=I=�OH=S�G=r�F=��E=]2E=iD=�C=��B=�B=�:A=�l@=c�?=��>=M�==f(==T<=m~;=E�:=��9=i�8=�8=�:7=�[6=wz5=W�4=N�3=7�2=��1=��0=�0=�/=v&.=�1-=:,=�?+=$C*=yC)=A(=�;'=3&=w'%=�$=�#=O�!=�� =a�=��=Wy=^R=�'=>�=�=ߐ=�V=�=��=�=G=�=�=�P=��=��
=M6	=��=�e=c�=8�==� =�.�<�+�</!�<p�<���<���<E��<��<CO�<M�<��<��<'C�<���<���<?�<F��<�x�<�<���<g-�<趹<�<�<��<>�<'��<J3�<橤<�<���<���<�m�<�ڒ<�E�<���<�<��<a�<Сz<�ps<�?l<�e<8�]<\�V<c�O<�\H<5A<_:<��2<�+<ϻ$<-�<��<ʐ<��<%�<c6�;JY�;G��;;��;- �;���;���;慕;�$�;2�u;�@[;��@;E�&;x	;��:��:��:"�:�Vi9�.!��
���j��b���Ժ����5��;0��G�}�]���s�d넻�͏�~���o2����������TĻ�tλtػ�S���.����5���K����р�	��z����6;���#���'�^�+�60�}04�c;8�r:<��-@��D���G���K���O�xJS���V�#�Z��J^�X�a��se���h��{l�_�o�pes���v�3z�=�}��s���������vd���������7>��x׋��n���������(��Q����F��9Ӗ��^���虼Bq���������5������A�������������������������|������B�������������쟹��!��գ���&���  �  �lN=��M=L�L=s%L=$bK=U�J=��I=I=�OH=Y�G=o�F=��E=Z2E=iD=��C=��B=�B=�:A=�l@=g�?=��>=O�==\(==T<=k~;=K�:=��9=o�8=�8=�:7=�[6=sz5=`�4=Q�3=5�2=��1=��0=�0=�/=w&.=�1-=:,=�?+=(C*=�C)=�@(=�;'=	3&=r'%=�$=�#=S�!=�� =c�=��=Yy=aR=�'=A�=��=��=�V=�=��=�=G=�=�=�P=��=��
=H6	=��=�e=n�=8�==� =�.�<�+�<,!�<r�<���<���<T��<��<SO�<G�<��<���<(C�<���<���<?�<7��<�x�<s�<���<c-�<߶�<�<�<	��<!>�<$��<M3�<ש�<��<폝<���<n�<�ڒ<�E�<ꯋ<�<z��<h�<�z<�ps<�?l<�e<O�]<t�V<U�O<�\H<g5A<l:<��2</�+<һ$<(�<��<��<��< �<�6�;9Y�;1��;#��; �;���;���;慕;U$�;�u;�@[;��@;`�&;�;���:���:��:��:�]i9�-!��
��j��c����Ժ����5��;0��G�̈]���s�[넻$Ώ�����<2������O���TĻ�tλTtػ T⻿�:���s5���K��������z����+;���#���'�c�+�20��04��;8�v:<��-@��D���G���K�ԌO��JS���V��Z��J^�V�a��se���h��{l�<�o�xes���v�33z�<�}�us���������}d���������6>��w׋��n���������(��]����F��=Ӗ��^���虼Kq���������1���������D������������옪����������t������C������������������!��ڣ���&���  �  �jN=K�M=��L=^"L=�^K=��J=��I=�I=�JH=�G=��F=��E=�+E=/bD=��C=�B=��A=%2A=�c@=Փ?=��>=��==S==�H<=Tr;=��:=|�9=��8=Y
8=',7=FL6=uj5=̆4=!�3=n�2=��1=��0=C�/=�/=�.=-=�#,=0)+=�+*=o+)=@((=6"'=&=�%=��#=��"=�!=�� =�=�~=[=�3=�=��=�=�p=]6=.�=�=�o=�%=��=��=�/=��=hw
=E	=+�=E=�=2e=v�=�u =��<��<���<��<g��<���<�y�<�M�<�<���<R��<�_�<��<���<�p�<e�<D��<}S�<��<g~�<��<㘹<� �<���<�%�<a��<}�<ϖ�<��<���<_�<mb�<�В<>�<թ�<��<�<��<H�z<�vs<�Il<�e<A�]<��V<��O<�xH<�TA<�4:<x3<��+<��$<��<��<p�<-�<��<{��;��;p �;li�;�¾;�.�;��;t=�;'�;a7w;9�\;��B;��(;f�;�8�:N�:�̈́:7h%:!�9�����o�b�B���к�����d.���D��V[�֚q�σ�����r��G��e������{8û2YͻnZ׻�;��������$��*��{h�N��H�����@d�~��m#��M'�р+��/���3�N�7���;���?�A�C��G��dK�6/O���R�i�V��SZ���]�.�a��%e�w�h�,3l�%�o��!s�a�v�^�y��S}�gV�� �������J��솼����'������Z��+���]������s���o6��Ė�)P���ڙ��d��휼st������d�����������M����������<���������꘰�������2������M��R����#������*���  �  �jN=T�M=��L=_"L=�^K=��J=��I=�I=�JH=�G=üF=��E=�+E=1bD=��C=!�B=��A=$2A=�c@=ړ?=��>=��==T==�H<=Xr;=��:=��9=��8=H
8=#,7=AL6=yj5=І4=&�3=o�2=��1=��0=C�/=�/=�.=-=�#,=%)+=�+*=n+)=E((=4"'=&=�%=��#=��"=�!=ǻ =�=�~=[=�3=�=��=�=�p=e6=2�=�=�o=�%=��=��=�/=��=Yw
=A	=(�=E=�=8e=u�=�u =$��<��<���<��<b��<מ�<�y�<�M�<|�<���<F��<�_�<��<���<�p�<u�<F��<iS�<��<V~�<��<ژ�<� �<���<�%�<p��<y�<Җ�<��<���<b�<nb�<�В<�=�<©�<��<�<��<M�z<�vs<�Il<�e<H�]<�V<��O<�xH<�TA<�4:<�3<��+<��$<��<��<t�<%�<�<���;X��;G �;1i�;�¾;\.�;(��;$=�;�;�7w;{�\;J�B;s�(;w�;�7�:�N�:~̈́:Dj%:�"�9-����÷b��A����к�����.�a�D��V[�J�q�%σ�"���@s������������T8ûAYͻ�Z׻�;���껭����$�����h�T��R�����?d����W#��M'���+���/���3�T�7���;���?�H�C��G��dK�u/O���R�r�V��SZ���]��a��%e�u�h�3l��o��!s�r�v�j�y��S}�hV�����������J��솼����'�������Y�����Z������m���6��Ė�2P���ڙ��d���으ct������a�����������L����������O���������ܘ��������:������J��F����#������*���  �  �jN=Y�M=��L=["L=�^K=��J=��I=�I=�JH=�G=ļF=��E=�+E=:bD=��C=,�B=��A='2A=�c@=ғ?=��>=��==[==�H<=_r;=��:=��9=��8=M
8=2,7=<L6=zj5=ˆ4="�3=l�2=��1=��0==�/=�/=�.=-=�#,=&)+=�+*=c+)=I((=3"'=&=�%=��#=��"=�!=ͻ =�=�~=[=�3=�=��=!�=�p=`6=(�=
�=�o=�%=��=��=�/=��=cw
=J	=$�=E=�=8e=q�=�u =��<���<���<��<~��<��<�y�<�M�<l�<���<B��<�_�<x�<���<�p�<i�<L��<eS�<��<P~�<��<☹<~ �<���<�%�<l��<f�<ܖ�<��<���<`�<[b�<�В<�=�<ߩ�<��<�<��<8�z<�vs<�Il<�e<8�]<�V<��O<�xH<UA<�4:<�3<��+<��$<��<��<��<�<�<V��;b��;H �;?i�;Aþ;;.�;���;=�;1�;�7w;��\;�B;�(;��;�7�:mO�:�̄:i%:e$�9�����̸b�uA��6�кQ���5��.�T�D��V[��q�Fσ�ﰎ��r�����ҕ��b���58ûIYͻpZ׻�;�$��̠���$������h�3��L�����d����C#��M'�Ȁ+�#�/���3�C�7���;���?�p�C�ޏG��dK�M/O���R���V��SZ���]��a��%e���h�!3l�6�o��!s���v�1�y��S}�dV�����������J��솼�����'������Z��&���U������W����6�� Ė�*P�� ۙ��d��휼gt������W�����������`����������1���������٘��������C������R��F����#�������)���  �  �jN=R�M=��L=^"L=�^K=��J=��I=�I=�JH=�G=��F=��E=�+E=3bD=��C="�B=��A=)2A=�c@=ٓ?=��>=��==Z==�H<=\r;=��:=��9=��8=O
8=',7=:L6=|j5=͆4=%�3=n�2=��1=��0=C�/=�/=�.= -=�#,=')+=�+*=k+)=I((=1"'=&=�%=��#=��"=�!=˻ =�=�~=[=�3=�=��= �=�p=f6=0�=�=�o=�%=��=��=�/=��=aw
=?	=%�=E=�=7e=u�=�u =��<��<���<��<e��<��<�y�<�M�<w�<���<>��<�_�<|�<���<�p�<i�<P��<fS�<��<Y~�<��<ؘ�<� �<���<�%�<z��<q�<ٖ�<��<���<g�<hb�<�В<�=�<ҩ�<��<	�<��<K�z<�vs<�Il<�e<E�]<
�V<��O<nxH<�TA<�4:<�3<��+<��$<��<��<��<�<�<���;K��;[ �;"i�;þ;e.�;2��;=�;B�;�7w;m�\;v�B;,�(;��;�7�:O�:<̈́:Oi%:s"�9 ����`�b�;A���к����z.�^�D��V[�I�q�>σ�E����r��������#���.8û\YͻvZ׻�;���껚����$������h�R��L�����>d����H#��M'���+��/���3�H�7���;���?�Q�C��G��dK�S/O���R��V��SZ���]��a��%e�w�h�3l�"�o��!s���v�c�y��S}�iV��  �������J��"솼����'�������Y��&���Q������m���}6��	Ė�5P���ڙ��d��휼Zt������Z�����#���~��R����������?���������ޘ��������<������K��J����#������*���  �  �jN=O�M=��L=\"L=�^K=��J=��I=�I=�JH=�G=��F=��E=�+E=2bD=��C= �B=��A='2A=�c@=ԓ?=��>=��==W==�H<=Yr;=��:=��9=��8=P
8=&,7=FL6=zj5=ˆ4=$�3=i�2=��1=��0=E�/=�/=�.=-=�#,=))+=�+*=l+)=D((=6"'=&=�%=��#=��"=�!=Ȼ =�=�~=[=�3=�=��=�=�p=^6=.�=�=�o=�%=��=��=�/=��=`w
=B	=/�=E=�=3e=v�=�u =��<��<���<��<f��<��<�y�<�M�<w�<���<G��<�_�<��<���<�p�<l�<L��<rS�<��<a~�<��<ޘ�<� �<���<�%�<g��<t�<Ԗ�<��<���<_�<kb�<�В<�=�<ʩ�<��<�<��<T�z<�vs<�Il<�e<J�]<��V<��O<�xH<�TA<�4:<�3<��+<��$<��<��<~�<�<��<���;;��;\ �;Ei�;þ;�.�; ��;D=�;6�;�7w;%�\;�B;i�(;��;8�:�N�:̈́:�i%:!�9�����x�b��A��)�к���`�g.���D�wV[�Úq��΃����s�����������U8û3Yͻ~Z׻�;��������$��	���h�S��H�����Bd����Q#��M'�΀+��/���3�M�7���;���?�K�C���G��dK�W/O���R�W�V��SZ���]�*�a��%e���h�$3l�%�o��!s�]�v�a�y��S}�lV�����������J��솼����'������Z��#���U������q���t6��
Ė�.P���ڙ��d��휼mt������_�����������P����������G���������혰�������9������I��S����#������	*���  �  �jN=U�M=��L=\"L=�^K=��J=��I=�I=�JH=�G=üF=��E=�+E=4bD=��C='�B=��A=$2A=�c@=֓?=��>=��==V==�H<=]r;=��:=��9=��8=N
8=*,7=<L6=xj5=Ά4="�3=l�2=��1=��0=E�/=�/=�.=-=�#,=%)+=�+*=g+)=G((=4"'=&=�%=��#=��"=�!=Ȼ =�=�~=[=�3=�=��=�=�p=a6=0�=�=�o=�%=��=��=�/=~�=bw
=@	=$�=E=�=2e=w�=�u =��<��<���<��<k��<��<�y�<�M�<n�<���<C��<�_�<��<���<�p�<t�<F��<mS�<��<U~�<��<䘹< �<���<�%�<l��<t�<ږ�<��<���<_�<cb�<�В<�=�<ҩ�<��<�<��<R�z<�vs<�Il<�e<G�]<�V<��O<vxH<�TA<�4:<�3<��+<��$<��<��<��< �<�<���;X��;? �;Vi�;þ;Z.�;T��;5=�;�;�7w;A�\;Y�B;l�(;��;�7�:'O�:�̄:�i%:�!�9ɧ���ڸb��A���к[���:�B.���D�vV[�i�q�Hσ�3����r�����핮�?���D8û?Yͻ~Z׻�;����à���$�����h�D��V�����1d����U#��M'���+��/���3�J�7���;���?�`�C��G��dK�Q/O���R���V��SZ���]�,�a��%e�{�h�(3l�"�o��!s���v�U�y��S}�nV�����������J��솼����'������Z�����[������d����6��	Ė�(P�� ۙ��d��휼ht������Y�����������W����������?�������������������3������K��H����#������*���  �  �jN=V�M=��L=a"L=�^K=��J=��I=�I=�JH=	�G=ƼF=��E=�+E=3bD=��C=$�B=��A=,2A=�c@=ԓ?=��>=��==Z==�H<=`r;=��:=��9=��8=J
8=+,7=;L6=�j5=͆4="�3=m�2=��1=��0=@�/=�/=�.=-=�#,=#)+=�+*=f+)=M((=1"'=&=�%=��#=��"=�!=л =�=�~=[=�3=�=��=$�=�p=c6=0�=�=�o=�%=��=��=�/=�=cw
=B	='�=E=�=3e=s�=�u =��<��<���<��<m��<���<�y�<�M�<q�<���<>��<�_�<v�<���<�p�<p�<W��<iS�<
��<Y~�<��<ܘ�<� �<���<�%�<q��<i�<ږ�<��<���<l�<ab�<�В<�=�<֩�<��<�<��<<�z<�vs<�Il<�e<5�]<�V<��O<mxH<UA<{4:<�3<��+<��$<��<��<��<�<�<m��;s��;l �;3i�;
þ;e.�;<��; =�;Z�;�7w;"�\;f�B;��(;��;�7�:�O�:3̈́:�i%:C#�9\����4�b��@���кd���$��.���D��V[���q�-σ�0����r�����핮�G���8ûYYͻkZ׻�;���껸����$������h�M��L�����;d����4#��M'���+��/���3�D�7���;���?�f�C��G��dK�K/O���R�x�V��SZ���]�)�a��%e�{�h�'3l�+�o��!s���v�R�y��S}�hV�����������J��!솼 ����'������Z�� ���J������k���}6��Ė�0P���ڙ��d��	휼ct������Y��������y��Z����������:���������ؘ��������A������S��C����#�������)���  �  �jN=T�M=��L=_"L=�^K=��J=��I=�I=�JH=�G=��F=��E=�+E=2bD=��C=!�B=��A=&2A=�c@=Փ?=��>=��==Z==�H<=Yr;=��:=�9=��8=O
8=(,7=>L6=zj5=ˆ4=%�3=k�2=��1=��0=B�/=�/=�.=-=�#,=))+=�+*=i+)=I((=0"'=&=�%=��#=��"=�!=ɻ =�=�~=[=�3=�=��=�=�p=a6=/�=	�=�o=�%=��=��=�/=��=cw
=@	=*�=E=�=6e=r�=�u =��< ��<���<��<i��<��<�y�<�M�<v�<���<@��<�_�<}�<���<�p�<h�<J��<tS�<��<e~�<��<ߘ�<� �<���<�%�<o��<t�<֖�<��<���<f�<bb�<�В<�=�<թ�<��<�<��<H�z<�vs<�Il<�e<F�]<��V<��O<{xH<�TA<�4:<�3<��+<��$<��<��<��<�<�<z��;;��;^ �;Mi�;þ;�.�;%��;O=�;0�;�7w;7�\;C�B;M�(;��;�7�:�N�:3̈́:i%:�#�91��n�A�b�nA��=�к����<��.�k�D��V[���q�σ�2����r��������3���08û_YͻxZ׻�;���������$�����h�N��F�����=d����O#��M'�À+��/���3�J�7���;���?�X�C��G��dK�M/O���R�i�V��SZ���]��a��%e���h�3l�0�o��!s�w�v�Z�y��S}�fV�� �������J�� 솼�����'������Z��'���W������q���q6��
Ė�-P���ڙ��d��휼dt������]�����"�����X����������<���������昰�������D������K��O����#������ *���  �  �jN=S�M=��L=\"L=�^K=��J=��I=�I=�JH=�G=ļF=��E=�+E=0bD=��C=!�B=��A= 2A=�c@=ړ?=��>=��==T==�H<=Zr;=��:=��9=��8=O
8=&,7=>L6=xj5=І4=!�3=l�2=��1=��0=E�/=�/=�.=-=�#,=')+=�+*=k+)=D((=5"'=&=�%=��#=��"=�!=ƻ =�=�~=[=�3=�=��=�=�p=a6=.�=�=�o=�%=��=��=�/=��=`w
=>	='�=E=�=0e=w�=�u =��<
��<���<��<b��<��<�y�<�M�<x�<���<J��<�_�<��<���<�p�<}�<=��<tS�<��<`~�<��<㘹< �<���<�%�<f��<x�<Ж�<��<���<_�<fb�<�В<�=�<̩�<��<�<��<M�z<�vs<�Il<�e<B�]<�V<��O<xxH<�TA<�4:<�3<��+<��$<��<��<p�<*�<��<���;_��;7 �;Xi�;�¾;�.�;*��;T=�;��;/8w;��\;�B;y�(;p�;Y8�:�N�:B̈́:�i%:�!�9G����k�b��A����к`���4�Q.���D�tV[�^�q�2σ�=���s��������"���W8û8YͻpZ׻�;����Ϡ��p$�����h�K��N�����;d����c#�yM'���+�
�/���3�M�7���;���?�O�C��G��dK�W/O���R�v�V��SZ���]�1�a��%e�{�h�+3l��o��!s�}�v�g�y��S}�lV��  �������J��솼����'�������Y�����c������n���u6��Ė�)P�� ۙ��d���으mt������c����� ������T����������E���������ߘ��������7������M��I����#������*���  �  �jN=V�M=��L=]"L=�^K=��J=��I=�I=�JH=	�G=üF=��E=�+E=6bD=��C=&�B=��A=(2A=�c@=ѓ?=��>=��==V==�H<=]r;=��:=��9=��8=M
8=0,7==L6={j5=ˆ4=�3=l�2=��1=��0=?�/=�/=�.=-=�#,=%)+=�+*=f+)=H((=5"'=&=�%=��#=��"=�!=̻ =�=�~=[=�3=�=��= �=�p=_6=/�=�=�o=�%=��=��=�/=��=cw
=F	=%�=E=�=2e=t�=�u =��< ��<���<��<t��<��<�y�<�M�<o�<���<F��<�_�<�<���<�p�<k�<N��<nS�<��<]~�<��<䘹<� �<���<�%�<h��<u�<֖�<��<���<d�<]b�<�В<�=�<ک�<��<�<��<7�z<�vs<�Il<�e</�]<�V<��O<~xH<UA<�4:<�3<��+<��$<��<��<~�< �<�<p��;Y��;T �;Ui�; þ;|.�;P��;==�;A�;�7w;��\;I�B;Q�(;��;(8�:>O�:�̄:xi%:�"�9ۨ�����b�]A��"�к����,��.���D��V[�9�q�@σ�����r�����󕮻I���58û9YͻxZ׻�;����נ���$������h�B��F�����,d����F#��M'�ɀ+��/���3�K�7���;���?�e�C��G��dK�L/O���R�~�V��SZ���]�-�a��%e�}�h�.3l�1�o��!s���v�C�y��S}�iV�����������J��솼����'������
Z��$���R������c���x6��Ė�(P���ڙ��d��휼kt������]�����������]����������7���������ܘ�����	���@������V��G����#�������)���  �  �jN=W�M=��L=a"L=�^K=��J=��I=�I=�JH=�G=��F=��E=�+E=5bD=��C=&�B=��A=+2A=�c@=ړ?=��>=��==^==�H<=Zr;=��:=��9=��8=G
8=),7=8L6=}j5=ʆ4=%�3=p�2=��1=��0==�/=�/=�.=-=�#,=#)+=�+*=i+)=K((=/"'=&=�%=��#=��"=�!=̻ =�=�~=[=�3=�=��="�=�p=k6=/�=�=�o=�%=��=��=�/=~�=[w
=>	="�=E=�=;e=p�=�u =$��<���<���<���<h��<מ�<�y�<�M�<s�<���<6��<�_�<|�<���<�p�<h�<T��<bS�<��<T~�<��<ޘ�<� �<���<�%�<~��<p�<���<��<���<k�<ab�<�В<�=�<Ω�<��<�<��<=�z<�vs<vIl<e<:�]<�V<��O<cxH<�TA<~4:<�3<��+<��$<��<��<��<�<(�<���;H��;^ �;:i�;þ;[.�;O��;=�;X�;�7w;��\;��B;$�(;�;D7�:�N�:4̈́:�i%:�#�9f��3�˹b�A��W�к������.��D��V[�O�q�Iσ�@���s�����䕮�.���!8ûkYͻjZ׻�;����u����$������h�D��Q�����)d����=#��M'���+��/���3�<�7���;���?�W�C��G��dK�k/O���R���V��SZ���]��a��%e�x�h�3l�7�o��!s���v�\�y��S}�hV�����������J��)솼�����'�������Y��'���L������b����6��	Ė�.P���ڙ��d��휼Ut������S�����%���z��Y����������C���������ᘰ��������L������Q��L����#������*���  �  �jN=P�M=��L=\"L=�^K=��J=��I=�I=�JH=�G=��F=��E=�+E=5bD=��C=%�B=��A=)2A=�c@=ؓ?=��>=��==X==�H<=[r;=��:=�9=��8=Q
8=+,7=BL6=yj5=ˆ4= �3=k�2=��1=��0=?�/=�/=�.=-=�#,=))+=�+*=k+)=B((=7"'=&=�%=��#=��"=�!=ɻ =�=�~=[=�3=�=��=�=�p=`6=&�=�=�o=�%=��=��=�/=��=dw
=E	=+�=E=�=2e=r�=�u =��<���<���<��<n��<��<�y�<�M�<u�<���<L��<�_�<{�<���<�p�<q�<N��<oS�<��<\~�<��<䘹<� �<���<�%�<`��<h�<ז�<��<���<]�<eb�<�В<�=�<ԩ�<��<�<��<>�z<�vs<�Il<�e<7�]<�V<��O<�xH<�TA<�4:<�3<��+<��$<��<��<��<�<��<���;M��;i �;Xi�;þ;.�;J��;A=�;D�;�7w;d�\;��B;%�(;��;�8�:�N�:/̈́:i%:�!�9�����^�b��A��!�к����E��.���D��V[���q�σ�����r��}�����%���d8û*Yͻ^Z׻�;�(��ޠ���$�����h�9��E�����&d����J#��M'�Ā+�*�/���3�B�7���;���?�S�C���G��dK�F/O���R�f�V��SZ���]�,�a��%e���h�.3l�1�o��!s�i�v�O�y��S}�jV�� �������J��솼����'�������Y�����R������d���y6��Ė�(P���ڙ��d���으st������\�����������U����������=���������嘰�������C������R��N����#�������)���  �  �jN=O�M=��L=Y"L=�^K=��J=��I=�I=�JH=�G=��F=��E=�+E=4bD=��C= �B=��A="2A=�c@=ړ?=��>=��==K==�H<=Xr;=��:=��9=��8=S
8=#,7==L6=oj5=ӆ4=#�3=k�2=��1=��0=J�/=�/=�.=-=�#,=))+=�+*=p+)=>((=9"'=&=�%=��#=��"=�!=û =�=�~=[=�3=�=��=�=�p=d6=6�=�=�o=�%=��=��=�/=��=_w
==	=&�=E= �=1e=w�=�u =��<��<���<
��<]��<��<�y�<�M�<w�<���<O��<�_�<��<���<�p�<r�<>��<mS�<��<b~�<��<ܘ�<� �<���<�%�<h��<��<ϖ�<��<���<U�<rb�<�В<�=�<ɩ�<��<�~�<��<e�z<�vs<�Il<�e<W�]<�V<}�O<uxH<�TA<�4:<�3<��+<��$<��<��<e�<O�<�<���;C��;< �;Ci�;þ;�.�;"��;:=�;�;�7w;��\;h�B;�(;��;�8�:�N�:5̈́:j%:� �9j������b��B��3�к)���A�9.���D�&V[���q�Iσ�8���s��~����������8ûYͻ�Z׻�;ụ�� ��z$�����h�S��F�����Ad����i#��M'���+��/���3�s�7���;���?�D�C���G��dK�Y/O���R�y�V��SZ���]�0�a��%e�}�h�&3l��o�"s�{�v�p�y��S}�mV�����������J��솼���y'�������Y�����c������q���s6��Ė�1P���ڙ��d���으lt������d���!��������H����������H�������������������.������B��F����#������*���  �  �jN=P�M=��L=\"L=�^K=��J=��I=�I=�JH=�G=��F=��E=�+E=5bD=��C=%�B=��A=)2A=�c@=ؓ?=��>=��==X==�H<=[r;=��:=�9=��8=Q
8=+,7=BL6=yj5=ˆ4= �3=k�2=��1=��0=?�/=�/=�.=-=�#,=))+=�+*=k+)=B((=7"'=&=�%=��#=��"=�!=ɻ =�=�~=[=�3=�=��=�=�p=`6=&�=�=�o=�%=��=��=�/=��=dw
=E	=+�=E=�=2e=r�=�u =��<���<���<��<n��<��<�y�<�M�<u�<���<L��<�_�<{�<���<�p�<q�<N��<oS�<��<\~�<��<䘹<� �<���<�%�<`��<h�<ז�<��<���<]�<eb�<�В<�=�<ԩ�<��<�<��<>�z<�vs<�Il<�e<7�]<�V<��O<�xH<�TA<�4:<�3<��+<��$<��<��<��<�<��<���;M��;i �;Xi�;þ;.�;J��;A=�;D�;�7w;d�\;��B;%�(;��;�8�:�N�:/̈́:i%:�!�9�����^�b��A��!�к����E��.���D��V[���q�σ�����r��}�����%���d8û*Yͻ^Z׻�;�(��ޠ���$�����h�9��E�����&d����J#��M'�Ā+�*�/���3�B�7���;���?�S�C���G��dK�F/O���R�f�V��SZ���]�,�a��%e���h�.3l�1�o��!s�i�v�O�y��S}�jV�� �������J��솼����'�������Y�����R������d���y6��Ė�(P���ڙ��d���으st������\�����������U����������=���������嘰�������C������R��N����#�������)���  �  �jN=W�M=��L=a"L=�^K=��J=��I=�I=�JH=�G=��F=��E=�+E=5bD=��C=&�B=��A=+2A=�c@=ړ?=��>=��==^==�H<=Zr;=��:=��9=��8=G
8=),7=8L6=}j5=ʆ4=%�3=p�2=��1=��0==�/=�/=�.=-=�#,=#)+=�+*=i+)=K((=/"'=&=�%=��#=��"=�!=̻ =�=�~=[=�3=�=��="�=�p=k6=/�=�=�o=�%=��=��=�/=~�=[w
=>	="�=E=�=;e=p�=�u =$��<���<���<���<h��<מ�<�y�<�M�<s�<���<6��<�_�<|�<���<�p�<h�<T��<bS�<��<T~�<��<ޘ�<� �<���<�%�<~��<p�<���<��<���<k�<ab�<�В<�=�<Ω�<��<�<��<=�z<�vs<vIl<e<:�]<�V<��O<cxH<�TA<~4:<�3<��+<��$<��<��<��<�<(�<���;H��;^ �;:i�;þ;[.�;O��;=�;W�;�7w;��\;��B;$�(;�;D7�:�N�:3̈́:�i%:�#�9j��4�̹b�A��X�к������.��D��V[�O�q�Iσ�@���s�����䕮�.���!8ûkYͻjZ׻�;����u����$������h�D��Q�����)d����=#��M'���+��/���3�<�7���;���?�W�C��G��dK�k/O���R���V��SZ���]��a��%e�x�h�3l�7�o��!s���v�\�y��S}�hV�����������J��)솼�����'�������Y��'���L������b����6��	Ė�.P���ڙ��d��휼Ut������S�����%���z��Y����������C���������ᘰ��������L������Q��L����#������*���  �  �jN=V�M=��L=]"L=�^K=��J=��I=�I=�JH=	�G=üF=��E=�+E=6bD=��C=&�B=��A=(2A=�c@=ѓ?=��>=��==V==�H<=]r;=��:=��9=��8=M
8=0,7==L6={j5=ˆ4=�3=l�2=��1=��0=?�/=�/=�.=-=�#,=%)+=�+*=f+)=H((=5"'=&=�%=��#=��"=�!=̻ =�=�~=[=�3=�=��= �=�p=_6=/�=�=�o=�%=��=��=�/=��=cw
=F	=%�=E=�=2e=t�=�u =��< ��<���<��<u��<��<�y�<�M�<o�<���<F��<�_�<��<���<�p�<k�<N��<nS�<��<]~�<��<䘹<� �<���<�%�<h��<u�<֖�<��<���<d�<]b�<�В<�=�<ک�<��<�<��<7�z<�vs<�Il<�e</�]<�V<��O<~xH<UA<�4:<�3<��+<��$<��<��<~�< �<�<p��;Y��;T �;Ui�; þ;|.�;P��;==�;A�;�7w;��\;I�B;P�(;��;'8�:=O�:�̄:wi%:�"�9������b�^A��#�к����,��.���D��V[�9�q�Aσ�����r�����󕮻I���58û9YͻxZ׻�;����ؠ���$������h�B��G�����,d����F#��M'�ɀ+��/���3�K�7���;���?�e�C��G��dK�L/O���R�~�V��SZ���]�-�a��%e�}�h�.3l�1�o��!s���v�C�y��S}�iV�����������J��솼����'������
Z��$���R������c���x6��Ė�(P���ڙ��d��휼kt������]�����������]����������7���������ܘ�����	���@������V��G����#�������)���  �  �jN=S�M=��L=\"L=�^K=��J=��I=�I=�JH=�G=ļF=��E=�+E=0bD=��C=!�B=��A= 2A=�c@=ړ?=��>=��==T==�H<=Zr;=��:=��9=��8=O
8=&,7=>L6=xj5=І4=!�3=l�2=��1=��0=E�/=�/=�.=-=�#,=')+=�+*=k+)=D((=5"'=&=�%=��#=��"=�!=ƻ =�=�~=[=�3=�=��=�=�p=a6=.�=�=�o=�%=��=��=�/=��=`w
=>	='�=E=�=0e=w�=�u =��<
��<���<	��<c��<��<�y�<�M�<x�<���<J��<�_�<��<���<�p�<}�<=��<tS�<��<`~�<��<㘹< �<���<�%�<f��<x�<Ж�<��<���<_�<fb�<�В<�=�<̩�<��<�<��<M�z<�vs<�Il<�e<B�]<�V<��O<xxH<�TA<�4:<�3<��+<��$<��<��<p�<*�<��<���;_��;7 �;Xi�;�¾;�.�;*��;T=�;��;/8w;��\;
�B;x�(;p�;X8�:�N�:Ä́:�i%:�!�9N����l�b��A����кa���4�R.���D�tV[�_�q�2σ�=���s��������"���W8û8YͻpZ׻�;����Ϡ��p$�����h�K��N�����;d����c#�yM'���+�
�/���3�M�7���;���?�O�C��G��dK�W/O���R�v�V��SZ���]�1�a��%e�{�h�+3l��o��!s�}�v�g�y��S}�lV��  �������J��솼����'�������Y�����c������n���u6��Ė�)P�� ۙ��d���으mt������c����� ������T����������E���������ߘ��������7������M��I����#������*���  �  �jN=T�M=��L=_"L=�^K=��J=��I=�I=�JH=�G=��F=��E=�+E=2bD=��C=!�B=��A=&2A=�c@=Փ?=��>=��==Z==�H<=Yr;=��:=�9=��8=O
8=(,7=>L6=zj5=ˆ4=%�3=k�2=��1=��0=B�/=�/=�.=-=�#,=))+=�+*=i+)=I((=0"'=&=�%=��#=��"=�!=ɻ =�=�~=[=�3=�=��=�=�p=a6=/�=	�=�o=�%=��=��=�/=��=cw
=@	=*�=E=�=6e=r�=�u =��< ��<���<��<i��<��<�y�<�M�<v�<���<@��<�_�<}�<���<�p�<h�<J��<tS�<��<e~�<��<ߘ�<� �<���<�%�<o��<t�<֖�<��<���<f�<bb�<�В<�=�<թ�<��<�<��<H�z<�vs<�Il<�e<F�]<��V<��O<{xH<�TA<�4:<�3<��+<��$<��<��<��<�<�<z��;;��;^ �;Mi�;þ;�.�;%��;O=�;0�;�7w;7�\;C�B;M�(;��;�7�:�N�:3̈́:	i%:�#�99��o�C�b�oA��>�к ���<��.�l�D��V[���q�σ�2����r��������3���08û_YͻxZ׻�;���������$�����h�N��F�����=d����O#��M'�À+��/���3�J�7���;���?�X�C��G��dK�M/O���R�i�V��SZ���]��a��%e���h�3l�0�o��!s�w�v�Z�y��S}�fV�� �������J�� 솼�����'������Z��'���W������q���q6��
Ė�-P���ڙ��d��휼dt������]�����"�����X����������<���������昰�������D������K��O����#������ *���  �  �jN=V�M=��L=a"L=�^K=��J=��I=�I=�JH=	�G=ƼF=��E=�+E=3bD=��C=$�B=��A=,2A=�c@=ԓ?=��>=��==Z==�H<=`r;=��:=��9=��8=J
8=+,7=;L6=�j5=͆4="�3=m�2=��1=��0=@�/=�/=�.=-=�#,=#)+=�+*=f+)=M((=1"'=&=�%=��#=��"=�!=л =�=�~=[=�3=�=��=$�=�p=c6=0�=�=�o=�%=��=��=�/=�=cw
=B	='�=E=�=3e=s�=�u =��<��<���<��<m��<���<�y�<�M�<q�<���<>��<�_�<v�<���<�p�<p�<W��<iS�<
��<Y~�<��<ܘ�<� �<���<�%�<q��<i�<ږ�<��<���<l�<ab�<�В<�=�<֩�<��<�<��<<�z<�vs<�Il<�e<5�]<�V<��O<nxH<UA<{4:<�3<��+<��$<��<��<��<�<�<m��;s��;m �;3i�;
þ;e.�;<��; =�;Z�;�7w;!�\;f�B;��(;��;�7�:�O�:2̈́:�i%:?#�9d����6�b��@���кd���%��.���D��V[� �q�-σ�0����r�����핮�G���8ûYYͻkZ׻�;���껸����$������h�M��L�����<d����4#��M'���+��/���3�D�7���;���?�f�C��G��dK�K/O���R�x�V��SZ���]�)�a��%e�{�h�'3l�+�o��!s���v�R�y��S}�hV�����������J��!솼 ����'������Z�� ���J������k���}6��Ė�0P���ڙ��d��	휼ct������Y��������y��Z����������:���������ؘ��������A������S��C����#�������)���  �  �jN=U�M=��L=\"L=�^K=��J=��I=�I=�JH=�G=üF=��E=�+E=4bD=��C='�B=��A=$2A=�c@=֓?=��>=��==V==�H<=]r;=��:=��9=��8=N
8=*,7=<L6=xj5=Ά4="�3=l�2=��1=��0=E�/=�/=�.=-=�#,=%)+=�+*=g+)=G((=4"'=&=�%=��#=��"=�!=Ȼ =�=�~=[=�3=�=��=�=�p=a6=0�=�=�o=�%=��=��=�/=~�=bw
=@	=$�=E=�=2e=w�=�u =��<��<���<��<l��<��<�y�<�M�<n�<���<C��<�_�<��<���<�p�<t�<F��<mS�<��<U~�<��<䘹< �<���<�%�<l��<t�<ږ�<��<���<_�<cb�<�В<�=�<ҩ�<��<�<��<R�z<�vs<�Il<�e<G�]<�V<��O<vxH<�TA<�4:<�3<��+<��$<��<��<��< �<�<���;X��;? �;Vi�;þ;Z.�;T��;5=�;�;�7w;A�\;X�B;l�(;��;�7�:&O�:�̄:�i%:�!�9Ч���ܸb��A���к[���;�B.���D�vV[�j�q�Hσ�3����r�����핮�?���D8û?Yͻ~Z׻�;����à���$�����h�D��V�����1d����U#��M'���+��/���3�J�7���;���?�`�C��G��dK�Q/O���R���V��SZ���]�,�a��%e�{�h�(3l�"�o��!s���v�U�y��S}�nV�����������J��솼����'������Z�����[������d����6��	Ė�(P�� ۙ��d��휼ht������Y�����������W����������?�������������������3������K��H����#������*���  �  �jN=O�M=��L=\"L=�^K=��J=��I=�I=�JH=�G=��F=��E=�+E=2bD=��C= �B=��A='2A=�c@=ԓ?=��>=��==W==�H<=Yr;=��:=��9=��8=P
8=&,7=FL6=zj5=ˆ4=$�3=i�2=��1=��0=E�/=�/=�.=-=�#,=))+=�+*=l+)=D((=6"'=&=�%=��#=��"=�!=Ȼ =�=�~=[=�3=�=��=�=�p=^6=.�=�=�o=�%=��=��=�/=��=`w
=B	=/�=E=�=3e=v�=�u =��<��<���<��<f��<��<�y�<�M�<w�<���<G��<�_�<��<���<�p�<l�<L��<rS�<��<a~�<��<ޘ�<� �<���<�%�<g��<t�<Ԗ�<��<���<_�<kb�<�В<�=�<ʩ�<��<�<��<T�z<�vs<�Il<�e<J�]<��V<��O<�xH<�TA<�4:<�3<��+<��$<��<��<~�<�<��<���;;��;\ �;Ei�;þ;�.�;��;D=�;6�;�7w;$�\;�B;h�(;��;8�:�N�:̈́:�i%:!�9����z�b��A��*�к���`�g.���D�wV[�Úq��΃����s�����������U8û3Yͻ~Z׻�;��������$��	���h�S��H�����Bd����Q#��M'�΀+��/���3�M�7���;���?�K�C���G��dK�W/O���R�W�V��SZ���]�*�a��%e���h�$3l�%�o��!s�]�v�a�y��S}�lV�����������J��솼����'������Z��#���U������q���t6��
Ė�.P���ڙ��d��휼mt������_�����������P����������G���������혰�������9������I��S����#������	*���  �  �jN=R�M=��L=^"L=�^K=��J=��I=�I=�JH=�G=��F=��E=�+E=3bD=��C="�B=��A=)2A=�c@=ٓ?=��>=��==Z==�H<=\r;=��:=��9=��8=O
8=',7=:L6=|j5=͆4=%�3=n�2=��1=��0=C�/=�/=�.= -=�#,=')+=�+*=k+)=I((=1"'=&=�%=��#=��"=�!=˻ =�=�~=[=�3=�=��= �=�p=f6=0�=�=�o=�%=��=��=�/=��=aw
=?	=%�=E=�=7e=u�=�u =��<��<���<��<e��<��<�y�<�M�<w�<���<>��<�_�<|�<���<�p�<i�<P��<fS�<��<Y~�<��<ؘ�<� �<���<�%�<z��<q�<ٖ�<��<���<g�<hb�<�В<�=�<ҩ�<��<	�<��<K�z<�vs<�Il<�e<F�]<
�V<��O<nxH<�TA<�4:<�3<��+<��$<��<��<��<�<�<���;K��;[ �;"i�;þ;e.�;2��;=�;B�;�7w;m�\;v�B;+�(;��;7�:O�:;̈́:Ni%:p"�9&����a�b�;A���к����{.�_�D��V[�I�q�?σ�E����r��������#���/8û\YͻvZ׻�;���껚����$������h�R��L�����>d����H#��M'���+��/���3�H�7���;���?�Q�C��G��dK�S/O���R��V��SZ���]��a��%e�w�h�3l�"�o��!s���v�c�y��S}�iV��  �������J��"솼����'�������Y��&���Q������m���}6��	Ė�5P���ڙ��d��휼Zt������Z�����#���~��R����������?���������ޘ��������<������K��J����#������*���  �  �jN=Y�M=��L=["L=�^K=��J=��I=�I=�JH=�G=ļF=��E=�+E=:bD=��C=,�B=��A='2A=�c@=ғ?=��>=��==[==�H<=_r;=��:=��9=��8=M
8=2,7=<L6=zj5=ˆ4="�3=l�2=��1=��0==�/=�/=�.=-=�#,=&)+=�+*=c+)=I((=3"'=&=�%=��#=��"=�!=ͻ =�=�~=[=�3=�=��=!�=�p=`6=(�=
�=�o=�%=��=��=�/=��=cw
=J	=$�=E=�=8e=q�=�u =��<���<���<��<~��<��<�y�<�M�<l�<���<C��<�_�<x�<���<�p�<i�<L��<eS�<��<P~�<��<☹<~ �<���<�%�<l��<f�<ܖ�<��<���<`�<[b�<�В<�=�<ߩ�<��<�<��<8�z<�vs<�Il<�e<8�]<�V<��O<�xH<UA<�4:<�3<��+<��$<��<��<��<�<�<V��;b��;H �;?i�;Aþ;;.�;���;=�;1�;�7w;��\;�B;�(;��;�7�:mO�:�̄:i%:c$�9�����͸b�uA��6�кR���5��.�T�D� W[��q�Fσ�ﰎ��r�����ҕ��b���58ûIYͻpZ׻�;�$��͠���$������h�3��L�����d����C#��M'�Ȁ+�#�/���3�C�7���;���?�p�C�ޏG��dK�M/O���R���V��SZ���]��a��%e���h�!3l�6�o��!s���v�1�y��S}�dV�����������J��솼�����'������Z��&���U������W����6�� Ė�*P�� ۙ��d��휼gt������W�����������`����������1���������٘��������C������R��F����#�������)���  �  �jN=T�M=��L=_"L=�^K=��J=��I=�I=�JH=�G=üF=��E=�+E=1bD=��C=!�B=��A=$2A=�c@=ړ?=��>=��==T==�H<=Xr;=��:=��9=��8=H
8=#,7=AL6=yj5=І4=&�3=o�2=��1=��0=C�/=�/=�.=-=�#,=%)+=�+*=n+)=E((=4"'=&=�%=��#=��"=�!=ǻ =�=�~=[=�3=�=��=�=�p=e6=2�=�=�o=�%=��=��=�/=��=Yw
=A	=(�=E=�=8e=u�=�u =$��<��<���<��<b��<מ�<�y�<�M�<|�<���<F��<�_�<��<���<�p�<u�<F��<iS�<��<V~�<��<ژ�<� �<���<�%�<p��<y�<Җ�<��<���<b�<nb�<�В<�=�<©�<��<�<��<M�z<�vs<�Il<�e<H�]<�V<��O<�xH<�TA<�4:<�3<��+<��$<��<��<t�<%�<�<���;X��;G �;1i�;�¾;\.�;(��;$=�;�;�7w;{�\;J�B;s�(;w�;�7�:�N�:~̈́:Cj%:�"�9/����÷b��A����к�����.�a�D��V[�J�q�%σ�"���@s������������T8ûAYͻ�Z׻�;���껭����$�����h�T��R�����?d����W#��M'���+���/���3�T�7���;���?�H�C��G��dK�u/O���R�r�V��SZ���]��a��%e�u�h�3l��o��!s�r�v�j�y��S}�hV�����������J��솼����'�������Y�����Z������m���6��Ė�2P���ڙ��d���으ct������a�����������L����������O���������ܘ��������:������J��F����#������*���  �  �hN=+�M=�L=�L=�[K='�J=�I=zI=2FH=PG=��F=C�E=&E=�[D=�C=(�B=R�A=d*A=^[@=A�?=�>=W�==i===><=�g;=k�:=��9=x�8=��7=�7=y>6=*\5=�w4=Ñ3=��2=�1=��0=��/=y�.=��-=�-=,=�+=�*=�)=)(=�'=�&=-�$=M�#=/�"=һ!=� =�=;d=@=:=��=��=��=�S=d=��=��=kR=I=�=h=�=�=�Y
=��=�=	(=R�=�H=A�=Z =5��<
��<���<���<Y��<m�<�H�<3�<9��<��<�x�<v5�<���<]��<�J�<��<��<=2�<]��<V`�<�<~�<Q�<��<��<��<��<ȅ�<|��<�r�<H�<X�<Ȓ<�6�<P��<��<�|�<,�<��z<4|s<ARl<�(e<� ^<w�V<[�O<n�H<qA<HT:<9:3<�$,<�%<"<��<1�< 	<
<T6�;#f�;���;���;tT�;PƱ;�I�;�;���;�x;%@^;�D;*;RL;�a�:#��:��:#-,:8�9@�ʸ����Fs[�ё��'�̺����'��#,���B��`Y���o��т�#���4t��P��m��������:»�\̻<_ֻLB�$�6��B1���L����߇���ň����0Q� �"�O�&��+�A/��\3��l7�mp;��h?��UC��7G��K���N���R�|WV�,Z���]�MKa�W�d�5mh�!�k�Coo�B�r��Sv��y�<}�L<���恼�����3���Ն��u��=��~���}G���ގ��s�����?���(��p���HC���Ι�2Y��H✼vj�����w�����Ё�����G���V������������������!��陳����������������%�����-���  �  �hN=,�M=�L=�L=�[K="�J=�I=}I=7FH=OG=��F=?�E=&E=\D=�C=-�B=L�A=e*A=h[@=D�?=�>=Z�==q==6><=�g;=g�:=��9=s�8=��7=�7=w>6=,\5=�w4=��3=��2= �1=��0=��/=w�.=��-=�-=
,=�+=�*=�)=-(=�'=�&=5�$=Q�#=8�"=ջ!=� =�=9d=@=8=��=��=��=�S=l=��=��=oR=E=�=h=�=շ=�Y
=��=�=(=H�=�H=D�=Z =5��<��<���<���<\��<�l�<�H�<4�<.��<��<�x�<�5�<���<e��<�J�<$��<���</2�<c��<L`�<�<~�<E�<��<��<��<��<օ�<t��<�r�<P�<�W�<Ȓ<�6�<Q��<��<�|�<1�<k�z<=|s<IRl<�(e<p ^<�V<X�O<s�H<&qA<�S:<<:3<�$,<�%<"<t�<N�<$ 	<.
<L6�;_f�;t��;���;�T�;)Ʊ;�I�;���;���;��x;c@^;D;E*;�L;a�:@��:~�:d-,:�9�˸�����s[�����N�̺f����'�o#,���B�;aY��o��т����jt�����Q��������:»�\̻0_ֻB����/1���L��������͈���QQ��"�<�&�+�A/��\3��l7�p;��h?��UC��7G��K���N���R��WV�1Z���]�HKa�M�d�)mh� �k�Qoo�:�r� Tv��y��}�\<���恼�����3���Ն��u��6��u���pG��nގ��s�����9���(��d���PC���Ι�&Y��J✼ij��~񟼹w��$���Ё�����J���Q��ގ��������������3��噳����������������%�����-���  �  �hN=4�M=�L=�L=�[K=�J=�I=uI=8FH=FG=��F=?�E=&E=\D=�C=4�B=L�A=e*A=b[@==�?=�>=S�==s==/><=�g;=f�:=��9={�8=��7=�7=r>6=-\5=�w4=��3=��2=�1=��0=��/=|�.=��-=�-=,=�+=�*=�)=1(=�'=�&=3�$=J�#=8�"=˻!=� =�=?d=@=5=��=��=��=�S=j=��=��=oR=?=!�=�g=�=ط=�Y
=��=ޑ=(=F�=�H=A�=Z =7��<���<���<��<r��<�l�<�H�<9�<*��<���<�x�<�5�<���<b��<�J�<��<���</2�<s��<<`�<$�<
~�<F�<��<��< ��<��<؅�<k��<�r�<U�<�W�<Ȓ<�6�<g��<��<�|�<8�<\�z<N|s<9Rl<�(e<e ^<��V<N�O<k�H<UqA<�S:<_:3<s$,<�%<5<a�<U�< 	<3
<6�;Pf�;x��;���;�T�;�ű;(J�;���;���;<�x;�?^;
D;�*;�L;0`�:��:L�:[-,:��9T˸ϵ���t[�k���g�̺i����'��#,�Q�B�eaY�ġo��т�ݲ��$t�������������:»�\̻8_ֻ B�@���~1���L����͇���ۈ����OQ��"�a�&��+�A/��\3��l7��p;��h?��UC��7G��K���N�o�R��WV�Z���]�:Ka�Z�d�*mh��k�Yoo�-�r�Tv��y�v}�P<���恼�����3���Ն��u��B��w���|G��~ގ��s�����)���!(��^���JC���Ι�'Y��^✼gj���񟼷w��,���́�����V���>��㎪�������������;��ݙ�����������������%������,���  �  �hN=0�M=�L=�L=�[K=#�J=�I=vI==FH=NG=��F=D�E=&E=\D=�C=.�B=K�A=g*A=b[@=C�?=�>=S�==u==5><=�g;=i�:=��9=x�8=��7=�7=s>6=.\5=�w4=đ3=��2=�1=��0=��/=y�.=��-=�-=,=�+=�*=�)=.(=�'=�&=5�$=Q�#=<�"=һ!=� =�=:d=@=8=��=��=��=�S=o=�=��=sR=B=�= h=�=ٷ=�Y
=��=�=
(=J�=�H=?�=Z ==��< ��<���<��<[��<�l�<�H�<3�<0��<��<�x�<�5�<���<q��<�J�<��<���</2�<f��<K`�<�<~�<O�<��<��<)��<��<ۅ�<x��<�r�<Q�<�W�<Ȓ<�6�<R��<��<�|�<0�<r�z<O|s<-Rl<�(e<w ^<|�V<\�O<`�H<"qA<�S:<L:3<v$,<�%<,<{�<Y�< 	<G
<E6�;Cf�;���;���;�T�;Ʊ;�I�;���;ȋ�;8�x;W@^;vD;�*;M;�`�:���:��:-,:q�9˸Ļ���t[�K�����̺�����'��#,�i�B�aY��o��т�#���ft�����C��������:»�\̻_ֻB��˪�E1���L���������ψ����LQ��"�J�&�t+��@/��\3��l7��p;��h?��UC��7G��K���N���R��WV�'Z���]�<Ka�a�d�)mh��k�Woo�/�r�Tv��y�|}�T<���恼�����3���Ն��u��A��i���rG��zގ�}s�����6���(��f���PC���Ι�)Y��O✼_j���񟼴w�����Ё�����Q���H��܎��������������0��ܙ�����������������%�����-���  �  �hN=+�M= �L=�L=�[K=#�J=�I=zI=4FH=KG=��F=D�E=&E= \D=�C=,�B=P�A=g*A=e[@=@�?=�>=T�==o==8><=�g;=k�:=��9=v�8=��7=�7=}>6=)\5=�w4=đ3=��2=�1=��0=��/=r�.=��-=�-=,=�+=�*=�)=*(=�'=�&=.�$=P�#=2�"=ӻ!=� =�=:d=@=:=��=��=��=�S=e=��=��=nR=D=�=h=�=۷=�Y
=��=�=(=K�=�H=A�=Z =;��<���<���<��<^��<�l�<�H�<8�<7��<��<�x�<�5�<���<c��<�J�<��<���<82�<a��<R`�<�<~�<O�<��<��<��<��<̅�<u��<�r�<O�<X�<Ȓ<�6�<S��< �<�|�<(�<y�z<5|s<@Rl<�(e<~ ^<r�V<Y�O<��H<%qA<T:<::3<�$,<�%<<|�<>�< 	<#
<26�;?f�;���;���;�T�;AƱ;�I�;���;Ƌ�;f�x;@^;�D;�*;�L;Qa�:���:��:�-,:��99˸~���r[�䑝���̺�����'��#,���B��`Y�e�o��т�沍�Lt�����W��������:»�\̻3_ֻHB����:1���L������~�ƈ���=Q���"�A�&��+� A/��\3��l7��p;��h?��UC��7G��K���N���R�yWV�DZ���]�FKa�W�d�3mh��k�Woo�H�r��Sv��y�k}�T<���恼�����3���Ն��u��C��v���|G��tގ��s�����;���(��f���LC���Ι�-Y��P✼qj�����w��#���ҁ�����D���R��ӎ��������������,��陳����������������%������-���  �  �hN=0�M=�L=�L=�[K=#�J=�I=|I=9FH=LG=��F==�E=&E=\D=
�C=1�B=P�A=_*A=d[@=B�?=�>=X�==o==6><=�g;=f�:=��9=y�8=��7=�7=s>6='\5=�w4=Ñ3=�2="�1=��0=��/=z�.=��-=�-=,=�+=�*=�)=-(=�'=�&=/�$=R�#=7�"=ѻ!=� =�=@d=@=6=��=��=��=�S=i= �=��=pR=C=�= h=�=ٷ=�Y
=��=ߑ=(=L�=�H=C�=Z =9��<��<���<��<a��<�l�<�H�<5�<,��<��<�x�<�5�<���<i��<�J�<��<w��<82�<n��<A`�<�<~�<D�<��<��<"��<��<υ�<u��<�r�<L�<�W�<Ȓ<�6�<V��<��<�|�<9�<u�z<0|s<VRl<�(e<y ^<��V<=�O<j�H<,qA<T:<M:3<t$,<�%<2<z�<@�<! 	<7
<66�;Jf�;f��;���;�T�;�ű;J�;���;���;Y�x;8@^;)D;$*;�L;a�:�:W�:�,,:��9�˸ʺ���t[�����̺����'�P#,���B��`Y��o�҂����Kt�����<��������:»�\̻%_ֻ=B�����I1���L����ʇ���ֈ����>Q��"�I�&��+��@/��\3��l7��p;��h?��UC��7G��K���N���R��WV�-Z���]�HKa�O�d�4mh��k�Ioo�C�r�Tv��y�q}�R<���恼�����3���Ն��u��=��p���wG��vގ��s�����.���(��c���EC���Ι�+Y��O✼ej��~��w��"���ʁ�����R���J��׎��������������.��왳����������������%�����-���  �  �hN=3�M=�L=�L=�[K= �J=�I=wI=:FH=MG=��F=@�E=&E=\D=�C=/�B=I�A=f*A=e[@=C�?=�>=S�==u==2><=�g;=f�:=��9=z�8=��7=�7=u>6=.\5=�w4=��3=��2=�1=��0=��/=z�.=��-=�-=,=�+=�*=�)=1(=�'=�&=1�$=M�#=:�"=ѻ!=� =�=;d=@=9=��=��=��=�S=m=��=��=uR=?= �=�g=�=׷=�Y
=��=�=
(=D�=�H=A�=Z =7��<���<���<��<h��<�l�<�H�<9�<)��<���<�x�<�5�<���<g��<�J�<��<���<*2�<g��<M`�<�<~�<F�<��<��<%��<��<م�<r��<�r�<U�<�W�<Ȓ<�6�<V��<��<�|�<1�<Z�z<E|s<BRl<�(e<d ^<u�V<\�O<u�H<2qA<�S:<X:3<r$,<�%<#<n�<Z�< 	<<
<;6�;^f�;{��;���;�T�;*Ʊ;�I�;���;���;e�x;I@^;+D;�*;M;�`�:̋�:h�:-,:��9�˸¸��!t[�<�����̺z����'��#,���B�zaY��o��т�벍�Zt����� ��������:»�\̻_ֻ-B�%�ߪ�N1���L����އ�|�Ɉ����UQ��"�L�&�}+�
A/��\3��l7��p;��h?��UC��7G��K���N�}�R��WV�'Z���]�DKa�W�d�,mh��k�doo�-�r�Tv���y��}�Q<���恼�����3���Ն��u��D��r���tG��uގ�~s�����4���(��b���RC���Ι�$Y��Q✼cj���񟼵w��&���Ӂ�����S���D��ߎ��������������<��ᙳ����������������%�����-���  �  �hN=,�M=�L=�L=�[K= �J=�I={I=8FH=JG=��F=F�E=&E=�[D=�C=*�B=Q�A=i*A=_[@=?�?=�>=W�==r==3><=�g;=k�:=��9=v�8=��7=�7=v>6=*\5=�w4=Ƒ3=��2=�1=��0=��/=r�.=��-=�-=,=�+=�*=�)=/(=�'=�&=1�$=Q�#=6�"=ϻ!=� =�=;d=@=:=��=��=��=�S=j= �=��=rR=B=�=h=�=ط=�Y
=��=�=(=K�=�H=>�=Z =A��<���<���<��<c��<�l�<�H�<5�<3��<��<�x�<�5�<���<j��<�J�<��<���<<2�<b��<W`�<�<~�<T�<��<��<��<��<Յ�<p��<�r�<V�<�W�<Ȓ<�6�<U��<��<�|�<$�<t�z<L|s<&Rl<�(e<~ ^<f�V<U�O<q�H</qA<T:<>:3<�$,<%<<n�<O�< 	<3
<)6�;f�;���;���;�T�;SƱ;�I�;���;ڋ�;�x;@^;1D;*;�L;�`�:6��:��:;-,:U�9˸Z����s[�ב����̺�����'��#,�A�B�aY�Z�o��т�����Lt�����J��������:»�\̻"_ֻ-B�����[1���L����އ���ǈ����7Q���"�U�&��+��@/��\3��l7��p;��h?��UC��7G��K���N���R��WV�@Z���]�1Ka�e�d�4mh��k�\oo�C�r�Tv���y�n}�V<���恼�����3���Ն��u��?��o���zG���ގ�|s�����:���(��h���HC���Ι�3Y��U✼jj���񟼺w��(���ց�����K���Q��Վ��������������/��ޙ�����������������%�����-���  �  �hN=,�M=�L=�L=�[K='�J=�I=~I=6FH=SG=��F=@�E=&E= \D=�C=+�B=R�A=`*A=h[@=E�?=�>=Y�==n==:><=�g;=h�:=��9=t�8=��7=�7=v>6=)\5=�w4=3=��2= �1=��0=��/=w�.=��-=�-=,=�+=�*=�)=((=�'=�&=1�$=S�#=5�"=ڻ!=� =�=<d=@=9=��=��=��=�S=j=�=��=oR=H=�=h=�=ַ=�Y
=��=�=(=K�=�H=C�=Z =7��<��<���<���<X��<�l�<�H�<2�</��<��<�x�<5�<���<i��<�J�<(��<v��<;2�<a��<L`�<�<~�<J�<��<��<��<��<υ�<|��<�r�<G�<X�<Ȓ<�6�<M��<��<�|�<4�<q�z<8|s<ORl<�(e<u ^<��V<P�O<m�H<qA< T:<>:3<�$,<�%<)<��<<�<' 	<+
<k6�;Qf�;���;���;�T�;&Ʊ;�I�;�;���;��x;v@^;D;;*;�L;�a�:G��:��:-,:��9�˸�����s[�呝�M�̺-����'�u#,���B�aY��o��т����_t�����Q��������:»�\̻!_ֻ.B�����1���L����ڇ���ʈ����>Q��"�+�&��+��@/��\3��l7�rp;��h?��UC��7G��K���N���R��WV�4Z���]�QKa�Q�d�0mh��k�Poo�?�r� Tv��y�v}�Y<���恼�����3���Ն��u��9��q���qG��jގ��s�����:���(��h���FC���Ι�+Y��A✼lj��|��w�����́�����H���O��܎��������������0��虳����������������%�����-���  �  �hN=2�M=�L=�L=�[K=!�J=�I=yI=5FH=HG=��F=B�E=&E=\D=�C=1�B=P�A=e*A=g[@==�?=�>=T�==s==4><=�g;=h�:=��9=|�8=��7=�7=v>6=+\5=�w4=��3=��2=�1=��0=��/=y�.=��-=�-=,=�+=�*=�)=-(=�'=�&=0�$=O�#=3�"=ѻ!=� =�==d=@=8=��=��=��=�S=e=��=��=nR=B=�= h=�=۷=�Y
=��=�=	(=G�=�H=@�=Z =6��<���<���<��<m��<�l�<�H�<;�</��<��<�x�<�5�<���<d��<�J�<!��<���<72�<k��<D`�<$�<~�<K�<��<��<��<��<ԅ�<t��<�r�<S�<�W�<Ȓ<�6�<_��<��<�|�<4�<_�z<@|s<9Rl<�(e<e ^<��V<O�O<y�H<@qA<�S:<W:3<�$,<�%<&<s�<L�< 	<*
<6�;^f�;���;���;�T�;�ű;J�;���;���;��x;�?^;D;�*;�L;�`�:���:��:�-,:R�9�˸����s[�����b�̺g����'��#,���B�NaY��o��т�಍�3t�����)��������:»�\̻2_ֻ5B����L1���L����ԇ�}�Ј����BQ��"�H�&��+�A/��\3��l7��p;��h?��UC��7G��K���N�u�R��WV�+Z���]�CKa�\�d�6mh��k�Zoo�7�r�Tv��y�y}�K<���恼�����3���Ն��u��A��u����G��rގ��s�����1���(��^���HC���Ι�$Y��V✼mj���񟼻w��#���ρ�����L���E��������
����������9��䙳����������������%�� ���-���  �  �hN=2�M=�L=�L=�[K=!�J=�I=vI=BFH=JG=��F=E�E=
&E=\D=�C=2�B=K�A=i*A=a[@=B�?=�>=Q�==x==0><=�g;=i�:=��9=z�8=��7=�7=n>6=,\5=�w4=đ3=��2=�1=��0=��/=y�.=��-=�-=
,=�+=�*=�)=2(=�'=�&=2�$=Q�#=>�"=ͻ!=� =�=;d=@=8=��=��=��=�S=p=�=��=tR=?= �=�g=�=ٷ=�Y
=��=ݑ=
(=F�=�H=<�=Z =>��<���<���<��<d��<�l�<�H�</�<,��<���<�x�<�5�<���<v��<�J�<��<���<-2�<n��<J`�<!�<~�<O�<��<��<3��<��<ۅ�<v��<�r�<Z�<�W�<Ȓ<�6�<S��<��<�|�<-�<b�z<Z|s<Rl<�(e<l ^<q�V<U�O<Y�H<)qA<�S:<T:3<e$,<%<"<r�<_�< 	<]
<#6�;Ef�;���;���;�T�;Ʊ;J�;���;ڋ�;/�x;;@^;�D;�*;JM;_`�:ы�:��:G,,:��9�˸ֹ���u[�r�����̺�����'�$,�"�B�LaY��o�҂����pt�����@��������:»�\̻_ֻ(B�껼��k1���L����܇�}�̈����PQ��"�[�&�n+��@/��\3��l7��p;��h?��UC��7G��K���N���R��WV�'Z���]�,Ka�l�d�2mh��k�boo�2�r�!Tv���y��}�O<���恼�����3���Ն��u��F��c���rG��|ގ�ys�����.���(��`���PC���Ι�'Y��V✼Uj���񟼴w��"���Ձ�����Y���F������������������8��֙�����������������%�����-���  �  �hN=0�M=�L=�L=�[K=$�J=�I=xI=6FH=MG=��F=C�E=&E=\D=�C=.�B=N�A=e*A=e[@=@�?=�>=S�==o==6><=�g;=i�:=��9=z�8=��7=�7=y>6=-\5=�w4=��3=��2=�1=��0=��/=y�.=��-=�-=,=�+=�*=�)=,(=�'=�&=,�$=M�#=4�"=һ!=� =�=:d=	@=;=��=��=��=�S=g=��=��=oR=D=�=h=�=ݷ=�Y
=��=�=	(=F�=�H=@�=Z =3��<���<���<���<b��<�l�<�H�<3�<2��<��<�x�<�5�<���<b��<�J�<��<���<32�<e��<Q`�<�<~�<O�<��<��<��<��<ʅ�<w��<�r�<N�<�W�<Ȓ<�6�<Q��<��<�|�<.�<a�z<>|s<DRl<�(e<k ^<r�V<a�O<|�H<'qA<T:<L:3<{$,<�%<#<��<=�< 	<-
<A6�;Vf�;���;���;�T�;9Ʊ;�I�;���;���;g�x;%@^;D;�*;�L;a�:\��:��:-,:F�9�˸����6s[�n�����̺t����'��#,���B�PaY��o��т�߲��[t�����O��������:»�\̻,_ֻTB�'���A1���L������w�������FQ���"�G�&��+�A/�]3��l7��p;��h?��UC��7G��K���N�|�R��WV�(Z���]�KKa�[�d�1mh�$�k�boo�2�r��Sv���y�q}�L<���恼�����3���Ն��u��E��w���{G��uގ��s�����6���(��f���OC���Ι�(Y��M✼mj�����w�� ���Ӂ�����L���L��Ҏ����	����������8��䙳����������������%������-���  �  �hN=(�M="�L=�L=�[K=$�J=�I=�I=2FH=LG=��F=A�E=&E= \D=�C=+�B=X�A=d*A=g[@=>�?=�>=g�==l==9><=�g;=j�:=��9=s�8=��7=�7=y>6='\5=�w4=Ñ3=}�2="�1=��0=��/=u�.=��-=�-=,=�+=�*=�)=+(=�'=�&=6�$=]�#=2�"=׻!=� =�=9d=@=8=��=��=��=�S=e=�=��=lR=I=�=h=�=ط=�Y
=��=��=(=N�=�H=C�=Z =8��<
��<���<���<R��<�l�<�H�<3�<5��<��<�x�<z5�<���<l��<�J�<&��<���<G2�<a��<N`�<�<~�<Q�<��<��<��<��<х�<v��<�r�<M�<X�<�ǒ<�6�<K��<��<�|�<0�<{�z<%|s<VRl<�(e<~ ^<}�V<>�O<|�H<qA<T:<,:3<�$,<�%<"<|�<<�<\ 	<
<96�;Rf�;���;���;�T�;,Ʊ;�I�;.�;���;��x; @^;#D;*;�L;{a�:���:��:�-,:��9�˸ӽ���r[������̺	��� (�V#,���B��`Y�0�o�҂�����t�����{��������:»{\̻8_ֻB໧���1���L��������͈���&Q���"�.�&��+��@/��\3��l7�kp;��h?��UC��7G��K���N���R��WV�<Z���]�IKa�O�d�6mh��k�Aoo�G�r��Sv��y�|}�[<���恼�����3���Ն��u��"��m����G��lގ��s�����;���(��g���FC���Ι�*Y��L✼tj��_񟼾w��"���́�����>���[��؎��"������������+��񙳼���������������%������-���  �  �hN=0�M=�L=�L=�[K=$�J=�I=xI=6FH=MG=��F=C�E=&E=\D=�C=.�B=N�A=e*A=e[@=@�?=�>=S�==o==6><=�g;=i�:=��9=z�8=��7=�7=y>6=-\5=�w4=��3=��2=�1=��0=��/=y�.=��-=�-=,=�+=�*=�)=,(=�'=�&=,�$=M�#=4�"=һ!=� =�=:d=	@=;=��=��=��=�S=g=��=��=oR=D=�=h=�=ݷ=�Y
=��=�=	(=F�=�H=@�=Z =3��<���<���<���<b��<�l�<�H�<3�<2��<��<�x�<�5�<���<b��<�J�<��<���<32�<e��<Q`�<�<~�<O�<��<��<��<��<ʅ�<w��<�r�<N�<�W�<Ȓ<�6�<Q��<��<�|�<.�<a�z<>|s<DRl<�(e<k ^<r�V<a�O<|�H<'qA<T:<L:3<{$,<�%<#<��<=�< 	<-
<A6�;Vf�;���;���;�T�;9Ʊ;�I�;���;���;g�x;%@^;D;�*;�L;a�:\��:��:-,:E�9�˸����6s[�n�����̺t����'��#,���B�PaY��o��т�߲��[t�����O��������:»�\̻,_ֻTB�'���B1���L������w�������FQ���"�G�&��+�A/�]3��l7��p;��h?��UC��7G��K���N�|�R��WV�(Z���]�KKa�[�d�1mh�$�k�boo�2�r��Sv���y�q}�L<���恼�����3���Ն��u��E��w���{G��uގ��s�����6���(��f���OC���Ι�(Y��M✼mj�����w�� ���ҁ�����L���L��Ҏ����	����������8��䙳����������������%������-���  �  �hN=2�M=�L=�L=�[K=!�J=�I=vI=BFH=JG=��F=E�E=
&E=\D=�C=2�B=K�A=i*A=a[@=B�?=�>=Q�==x==0><=�g;=i�:=��9=z�8=��7=�7=n>6=,\5=�w4=đ3=��2=�1=��0=��/=y�.=��-=�-=
,=�+=�*=�)=2(=�'=�&=2�$=Q�#=>�"=ͻ!=� =�=;d=@=8=��=��=��=�S=p=�=��=tR=?= �=�g=�=ٷ=�Y
=��=ݑ=
(=F�=�H=<�=Z =>��<���<���<��<d��<�l�<�H�</�<,��<���<�x�<�5�<���<v��<�J�<��<���<-2�<n��<J`�<!�<~�<O�<��<��<3��<��<ۅ�<v��<�r�<Z�<�W�<Ȓ<�6�<S��<��<�|�<-�<b�z<Z|s<Rl<�(e<l ^<q�V<U�O<Y�H<)qA<�S:<T:3<e$,<%<"<r�<_�< 	<]
<#6�;Ef�;���;���;�T�;Ʊ;J�;���;ڋ�;/�x;;@^;�D;�*;JM;_`�:Ћ�:��:G,,:��9�˸ع���u[�s�����̺�����'�$,�"�B�MaY��o�҂����pt�����@��������:»�\̻_ֻ(B�껼��k1���L����܇�}�̈����PQ��"�[�&�n+��@/��\3��l7��p;��h?��UC��7G��K���N���R��WV�'Z���]�,Ka�l�d�2mh��k�boo�2�r�!Tv���y��}�O<���恼�����3���Ն��u��F��c���rG��|ގ�ys�����.���(��`���PC���Ι�'Y��V✼Uj���񟼴w��"���Ձ�����Y���F������������������8��֙�����������������%�����-���  �  �hN=2�M=�L=�L=�[K=!�J=�I=yI=5FH=HG=��F=B�E=&E=\D=�C=1�B=P�A=e*A=g[@==�?=�>=T�==s==4><=�g;=h�:=��9=|�8=��7=�7=v>6=+\5=�w4=��3=��2=�1=��0=��/=y�.=��-=�-=,=�+=�*=�)=-(=�'=�&=0�$=O�#=3�"=ѻ!=� =�==d=@=8=��=��=��=�S=e=��=��=nR=B=�= h=�=۷=�Y
=��=�=	(=G�=�H=@�=Z =6��<���<���<��<m��<�l�<�H�<;�</��<��<�x�<�5�<���<d��<�J�<!��<���<72�<k��<D`�<$�<~�<K�<��<��<��<��<ԅ�<t��<�r�<S�<�W�<Ȓ<�6�<_��<��<�|�<4�<_�z<@|s<9Rl<�(e<e ^<��V<O�O<y�H<@qA<�S:<W:3<�$,<�%<&<s�<L�< 	<*
<6�;^f�;���;���;�T�;�ű;J�;���;���;��x;�?^;D;�*;�L;�`�:���:��:�-,:P�9�˸����s[�����c�̺g����'��#,���B�NaY��o��т�಍�3t�����)��������:»�\̻2_ֻ5B����L1���L����ԇ�}�Ј����BQ��"�H�&��+�A/��\3��l7��p;��h?��UC��7G��K���N�u�R��WV�+Z���]�CKa�\�d�6mh��k�Zoo�7�r�Tv��y�y}�K<���恼�����3���Ն��u��A��u����G��rގ��s�����1���(��^���HC���Ι�$Y��V✼mj���񟼻w��#���ρ�����L���E��������
����������9��䙳����������������%�� ���-���  �  �hN=,�M=�L=�L=�[K='�J=�I=~I=6FH=SG=��F=@�E=&E= \D=�C=+�B=R�A=`*A=h[@=E�?=�>=Y�==n==:><=�g;=h�:=��9=t�8=��7=�7=v>6=)\5=�w4=3=��2= �1=��0=��/=w�.=��-=�-=,=�+=�*=�)=((=�'=�&=1�$=S�#=5�"=ڻ!=� =�=<d=@=9=��=��=��=�S=j=�=��=oR=H=�=h=�=ַ=�Y
=��=�=(=K�=�H=C�=Z =7��<��<���<���<X��<�l�<�H�<2�<0��<��<�x�<5�<���<i��<�J�<(��<v��<;2�<a��<L`�<�<~�<J�<��<��<��<��<υ�<|��<�r�<G�<X�<Ȓ<�6�<M��<��<�|�<4�<q�z<8|s<ORl<�(e<u ^<��V<P�O<m�H<qA< T:<>:3<�$,<�%<)<��<<�<' 	<+
<k6�;Qf�;���;���;�T�;&Ʊ;�I�;�;���;��x;v@^;D;;*;�L;�a�:G��:��:-,:��9�˸�����s[�呝�M�̺-����'�v#,���B�aY��o��т����_t�����Q��������:»�\̻!_ֻ.B�����1���L����ڇ���ʈ����>Q��"�+�&��+��@/��\3��l7�rp;��h?��UC��7G��K���N���R��WV�4Z���]�QKa�Q�d�0mh��k�Poo�?�r� Tv��y�v}�Y<���恼�����3���Ն��u��9��q���qG��jގ��s�����:���(��h���FC���Ι�+Y��A✼lj��|��w�����́�����H���O��܎��������������0��虳����������������%�����-���  �  �hN=,�M=�L=�L=�[K= �J=�I={I=8FH=JG=��F=F�E=&E=�[D=�C=*�B=Q�A=i*A=_[@=?�?=�>=W�==r==3><=�g;=k�:=��9=v�8=��7=�7=v>6=*\5=�w4=Ƒ3=��2=�1=��0=��/=r�.=��-=�-=,=�+=�*=�)=/(=�'=�&=1�$=Q�#=6�"=ϻ!=� =�=;d=@=:=��=��=��=�S=j= �=��=rR=B=�=h=�=ط=�Y
=��=�=(=K�=�H=>�=Z =A��<���<���<��<c��<�l�<�H�<5�<3��<��<�x�<�5�<���<j��<�J�<��<���<<2�<b��<W`�<�<~�<T�<��<��<��<��<Յ�<p��<�r�<V�<�W�<Ȓ<�6�<U��<��<�|�<$�<t�z<L|s<&Rl<�(e<~ ^<f�V<U�O<q�H</qA<T:<>:3<�$,<%<<n�<O�< 	<3
<)6�;f�;���;���;�T�;SƱ;�I�;���;ڋ�;�x;@^;1D;*;�L;�`�:6��:��::-,:R�9˸^����s[�ؑ����̺�����'��#,�A�B�aY�Z�o��т�����Lt�����J��������:»�\̻"_ֻ-B�����[1���L����އ���ǈ����7Q���"�U�&��+��@/��\3��l7��p;��h?��UC��7G��K���N���R��WV�@Z���]�1Ka�e�d�4mh��k�\oo�C�r�Tv���y�n}�V<���恼�����3���Ն��u��?��o���zG���ގ�|s�����:���(��h���HC���Ι�3Y��U✼jj���񟼺w��(���ց�����K���Q��Վ��������������/��ޙ�����������������%�����-���  �  �hN=3�M=�L=�L=�[K= �J=�I=wI=:FH=MG=��F=@�E=&E=\D=�C=/�B=I�A=f*A=e[@=C�?=�>=S�==u==2><=�g;=f�:=��9=z�8=��7=�7=u>6=.\5=�w4=��3=��2=�1=��0=��/=z�.=��-=�-=,=�+=�*=�)=1(=�'=�&=1�$=M�#=:�"=ѻ!=� =�=;d=@=9=��=��=��=�S=m=��=��=uR=?= �=�g=�=׷=�Y
=��=�=
(=D�=�H=A�=Z =7��<���<���<��<h��<�l�<�H�<9�<)��<���<�x�<�5�<���<g��<�J�<��<���<*2�<g��<M`�<�<~�<F�<��<��<%��<��<م�<r��<�r�<U�<�W�<Ȓ<�6�<V��<��<�|�<1�<Z�z<E|s<BRl<�(e<d ^<u�V<\�O<u�H<2qA<�S:<X:3<r$,<�%<#<n�<Z�< 	<<
<;6�;^f�;{��;���;�T�;*Ʊ;�I�;���;���;d�x;I@^;+D;�*;M;�`�:ˋ�:h�:
-,:��9�˸Ÿ��"t[�=�����̺{����'��#,���B�{aY��o��т�벍�Zt����� ��������:»�\̻_ֻ-B�%�ߪ�N1���L����އ�|�Ɉ����UQ��"�L�&�}+�
A/��\3��l7��p;��h?��UC��7G��K���N�}�R��WV�'Z���]�DKa�W�d�,mh��k�doo�-�r�Tv���y��}�Q<���恼�����3���Ն��u��D��r���tG��uގ�~s�����4���(��b���RC���Ι�$Y��Q✼cj���񟼵w��&���Ӂ�����S���D��ߎ��������������<��ᙳ����������������%�����-���  �  �hN=0�M=�L=�L=�[K=#�J=�I=|I=9FH=LG=��F==�E=&E=\D=
�C=1�B=P�A=_*A=d[@=B�?=�>=X�==o==6><=�g;=f�:=��9=y�8=��7=�7=s>6='\5=�w4=Ñ3=�2="�1=��0=��/=z�.=��-=�-=,=�+=�*=�)=-(=�'=�&=/�$=R�#=7�"=ѻ!=� =�=@d=@=6=��=��=��=�S=i= �=��=pR=C=�= h=�=ٷ=�Y
=��=ߑ=(=L�=�H=C�=Z =9��<��<���<��<a��<�l�<�H�<5�<,��<��<�x�<�5�<���<i��<�J�<��<w��<82�<n��<A`�<�<~�<D�<��<��<"��<��<υ�<u��<�r�<L�<�W�<Ȓ<�6�<V��<��<�|�<9�<u�z<0|s<VRl<�(e<y ^<��V<=�O<j�H<,qA<T:<N:3<t$,<�%<2<z�<@�<! 	<7
<66�;Jf�;f��;���;�T�;�ű;J�;���;���;Y�x;8@^;)D;$*;�L;a�:���:W�:�,,:��9�˸ͺ���t[�����̺����'�P#,���B��`Y��o�҂����Kt�����<��������:»�\̻%_ֻ=B�����I1���L����ʇ���ֈ����>Q��"�I�&��+��@/��\3��l7��p;��h?��UC��7G��K���N���R��WV�-Z���]�HKa�O�d�4mh��k�Ioo�C�r�Tv��y�q}�R<���恼�����3���Ն��u��=��p���wG��vގ��s�����.���(��c���EC���Ι�+Y��O✼ej��~��w��"���ʁ�����R���J��׎��������������.��왳����������������%�����-���  �  �hN=+�M= �L=�L=�[K=#�J=�I=zI=4FH=KG=��F=D�E=&E= \D=�C=,�B=P�A=g*A=e[@=@�?=�>=T�==o==8><=�g;=k�:=��9=v�8=��7=�7=}>6=)\5=�w4=đ3=��2=�1=��0=��/=r�.=��-=�-=,=�+=�*=�)=*(=�'=�&=.�$=P�#=2�"=ӻ!=� =�=:d=@=:=��=��=��=�S=e=��=��=nR=D=�=h=�=۷=�Y
=��=�=(=K�=�H=A�=Z =;��<���<���<��<^��<�l�<�H�<8�<7��<��<�x�<�5�<���<c��<�J�<��<���<82�<a��<R`�<�<~�<O�<��<��<��<��<̅�<u��<�r�<O�<X�<Ȓ<�6�<S��< �<�|�<(�<y�z<5|s<@Rl<�(e<~ ^<r�V<Y�O<��H<%qA<T:<::3<�$,<�%<<|�<>�< 	<#
<26�;?f�;���;���;�T�;AƱ;�I�;���;Ƌ�;f�x;@^;�D;�*;�L;Qa�:���:��:�-,:��9C˸����r[�䑝���̺�����'��#,���B��`Y�f�o��т�沍�Mt�����X��������:»�\̻3_ֻHB����:1���L������~�ƈ���=Q���"�A�&��+� A/��\3��l7��p;��h?��UC��7G��K���N���R�yWV�DZ���]�FKa�W�d�3mh��k�Woo�H�r��Sv��y�k}�T<���恼�����3���Ն��u��C��v���|G��tގ��s�����;���(��f���LC���Ι�-Y��P✼qj�����w��#���ҁ�����E���R��ӎ��������������,��陳����������������%������-���  �  �hN=0�M=�L=�L=�[K=#�J=�I=vI==FH=NG=��F=D�E=&E=\D=�C=.�B=K�A=g*A=b[@=C�?=�>=S�==u==5><=�g;=i�:=��9=x�8=��7=�7=s>6=.\5=�w4=đ3=��2=�1=��0=��/=y�.=��-=�-=,=�+=�*=�)=.(=�'=�&=5�$=Q�#=<�"=һ!=� =�=:d=@=8=��=��=��=�S=o=�=��=sR=B=�= h=�=ٷ=�Y
=��=�=
(=J�=�H=?�=Z ==��< ��<���<��<[��<�l�<�H�<3�<0��<��<�x�<�5�<���<q��<�J�<��<���</2�<f��<K`�<�<~�<O�<��<��<)��<��<ۅ�<x��<�r�<Q�<�W�<Ȓ<�6�<R��<��<�|�<0�<r�z<O|s<-Rl<�(e<w ^<|�V<\�O<`�H<"qA<�S:<L:3<v$,<�%<,<{�<Y�< 	<G
<E6�;Cf�;���;���;�T�;Ʊ;�I�;���;ȋ�;7�x;W@^;vD;�*;M;�`�:���:��:-,:o�9˸ƻ���t[�L�����̺�����'��#,�i�B�aY��o��т�#���ft�����C��������:»�\̻_ֻB��˪�E1���L���������ψ����LQ��"�J�&�t+��@/��\3��l7��p;��h?��UC��7G��K���N���R��WV�'Z���]�<Ka�a�d�)mh��k�Woo�/�r�Tv��y�|}�T<���恼�����3���Ն��u��A��i���rG��zގ�}s�����5���(��f���PC���Ι�)Y��O✼_j���񟼴w�����Ё�����Q���H��܎��������������0��ܙ�����������������%�����-���  �  �hN=4�M=�L=�L=�[K=�J=�I=uI=8FH=FG=��F=?�E=&E=\D=�C=4�B=L�A=e*A=b[@==�?=�>=S�==s==/><=�g;=f�:=��9={�8=��7=�7=r>6=-\5=�w4=��3=��2=�1=��0=��/=|�.=��-=�-=,=�+=�*=�)=1(=�'=�&=3�$=J�#=8�"=˻!=� =�=?d=@=5=��=��=��=�S=j=��=��=oR=?=!�=�g=�=ط=�Y
=��=ޑ=(=F�=�H=A�=Z =7��<���<���<��<s��<�l�<�H�<9�<*��<���<�x�<�5�<���<b��<�J�<��<���</2�<s��<<`�<$�<
~�<F�<��<��< ��<��<؅�<k��<�r�<U�<�W�<Ȓ<�6�<g��<��<�|�<8�<\�z<N|s<9Rl<�(e<e ^<��V<N�O<k�H<UqA<�S:<_:3<s$,<�%<5<a�<U�< 	<3
<6�;Pf�;x��;���;�T�;�ű;(J�;���;���;;�x;�?^;
D;�*;�L;0`�: ��:L�:[-,:��9[˸ѵ���t[�l���g�̺i����'��#,�Q�B�eaY�ġo��т�ݲ��$t�������������:»�\̻8_ֻ B�@���~1���L����͇���ۈ����OQ��"�a�&��+�A/��\3��l7��p;��h?��UC��7G��K���N�o�R��WV�Z���]�:Ka�Z�d�*mh��k�Yoo�-�r�Tv��y�v}�P<���恼�����3���Ն��u��B��w���|G��~ގ��s�����)���!(��^���JC���Ι�'Y��^✼gj���񟼷w��,���́�����V���>��㎪�������������;��ݙ�����������������%������,���  �  �hN=,�M=�L=�L=�[K="�J=�I=}I=7FH=OG=��F=?�E=&E=\D=�C=-�B=L�A=e*A=h[@=D�?=�>=Z�==q==6><=�g;=g�:=��9=s�8=��7=�7=w>6=,\5=�w4=��3=��2= �1=��0=��/=w�.=��-=�-=
,=�+=�*=�)=-(=�'=�&=5�$=Q�#=8�"=ջ!=� =�=9d=@=8=��=��=��=�S=l=��=��=oR=E=�=h=�=շ=�Y
=��=�=(=H�=�H=D�=Z =5��<��<���<���<\��<�l�<�H�<4�<.��<��<�x�<�5�<���<e��<�J�<$��<���</2�<c��<L`�<�<~�<E�<��<��<��<��<օ�<t��<�r�<P�<�W�<Ȓ<�6�<Q��<��<�|�<1�<k�z<=|s<IRl<�(e<p ^<�V<X�O<s�H<&qA<�S:<<:3<�$,<�%<"<t�<N�<$ 	<.
<L6�;_f�;t��;���;�T�;)Ʊ;�I�;���;���;��x;c@^;D;E*;�L;a�:@��:~�:d-,:�9�˸»���s[�����N�̺f����'�o#,���B�;aY��o��т����jt�����Q��������:»�\̻0_ֻB����/1���L��������͈���QQ��"�<�&�+�A/��\3��l7�p;��h?��UC��7G��K���N���R��WV�1Z���]�HKa�M�d�)mh� �k�Qoo�:�r� Tv��y��}�\<���恼�����3���Ն��u��6��u���pG��nގ��s�����9���(��d���PC���Ι�&Y��J✼ij��~񟼹w��$���Ё�����J���Q��ގ��������������3��噳����������������%�����-���  �  @gN=H�M=��L=%L=�XK=�J=��I=�I=NBH={G=�F=l�E=� E=�VD=>�C=�B=��A=�#A=)T@=��?=�>=��==�
==5<=�];=n�:=Y�9=��8=D�7=&7=L26=�O5=�j4=2�3=p�2=��1=}�0=,�/=o�.=X�-=��,=��+=�+=1*=�)=��'=��&=u�%=G�$=��#=i�"=��!=f� =�m=�L=6(= =K�=֤=�q=�:=��=R�=�~=v8=8�=��=�M=��=ĝ=�?
=��=)x=t=��=�/=t�=�A =���<���<́�<(s�<o]�<A�<��<f��<z��<X��<HR�<P�<���<�{�<�)�<��<�u�<��<��<�E�<�׼<gf�<�<Cx�<M��<1}�<U��<�v�<��<�f�<�ۙ<�N�<L��<x0�<s��<��<�z�<��<i�z<��s<�Yl<Q3e<�^<��V<{�O<��H<��A<�o:<�X3<�E,<=7%<O-<k(<�(<�/	<�<<���; ��;��;�o�;�Կ;�K�;�Ԥ;&q�;!�;�y;_;�^E;l+;��;�(�:�d�:��:�"2:/�9�����&��U�mS����ɺ�����y��p*��+A���W���m���iӌ�d����5�� �������[��P~˻ �ջ|f߻�+黪��[�������v ����k$�!�����A"���&���*��.��3��7�x;��?��C���F��J��N��VR��V���Y�l]��a��d��1h���k��7o���r�I v�N�y���|�H%���Ё�Ry��1��[�c��E��G���7���Ύ��d������Ɗ��T��`����7��ę�O���؜��a��F韼"p�����V{��������������u��叭�?���������蘳�5��Ɲ��{ ������-'��)����/���  �  >gN=J�M=��L=$L=�XK=�J=��I=�I=QBH={G=#�F=m�E=� E=�VD=B�C=�B=��A=�#A=)T@=��?=�>=��==�
==5<=�];=k�:=V�9=��8=D�7=-7=I26=�O5=�j4=.�3=q�2=��1=~�0=%�/=r�.=U�-=��,=��+=�+=1*=�)=��'=��&={�%=M�$=��#=j�"=��!=l� =�m=�L==(= =K�=Ӥ=�q=�:=��=P�=�~=~8=7�= �=�M=��==�?
=��=&x=y=�=�/=t�=�A =��<x��<ҁ�<!s�<|]�<
A�<��<`��<o��<_��<JR�<b�<���<�{�<)�<��<�u�<��<���<�E�<ؼ<`f�<�<Lx�<B��<7}�<U��<�v�<��<�f�<�ۙ<�N�<P��<w0�<���<��<�z�<��<J�z<�s<�Yl<c3e<�^<��V<{�O<w�H<�A<�o:<�X3<�E,<87%<F-<p(<()<�/	<�<<���;;��;�;�o�;տ;�K�;�Ԥ;q�;!�;�y;�~_;�^E;�k+;F�; )�:e�:q�:�!2:��9�����"鹆U�4S��)�ɺW���iy��p*�o+A��W�[�m��Yӌ�6����5����� ���[��\~˻�ջOf߻�+黡��&[�������{ ����P$�����uA"���&���*��.��3��7�|;��?��C���F��J��N��VR��V���Y�(l]��a��d��1h���k��7o���r�V v�5�y���|�E%���Ё�\y��+��X�c��G��H���7���Ύ��d����������K��O����7��ę�O���؜��a��G韼p�����Z{�����������������d��鏭�@��|������☳�3������� ������-'��.����/���  �  <gN=P�M=��L=(L=�XK=�J=��I=�I=XBH={G=$�F=o�E=� E=�VD=8�C=�B=��A=�#A=(T@=��?=��>=��==�
==5<=�];=m�:=V�9=��8=A�7=/7=C26=�O5=�j4=/�3=u�2=��1=��0=%�/=z�.=R�-=��,=��+=�+=7*=�)=��'=��&=v�%=I�$=��#=n�"=��!=n� =�m=�L=9(= =L�=Ӥ=�q=�:=��=P�=�~=z8=2�=�=�M=��=ŝ=�?
=��="x=�=�=�/=r�=�A =���<{��<݁�<s�<]�<A�<��<f��<s��<i��<=R�<^�<���<�{�<�)�<��<�u�<��<���<�E�<
ؼ<^f�<�<Qx�<?��<E}�<M��<�v�<��<�f�<�ۙ<�N�<[��<t0�<���<��<�z�<��<G�z<�s<�Yl<y3e<�^<��V<�O<`�H< �A<�o:<�X3<�E,<K7%<I-<U(<)<�/	<�<<���;D��;�;�o�;տ;�K�;դ;q�;7!�;�y;�~_;�^E;�k+;%�;I(�:�e�:��:�!2:��9ך���!�+U��R��ǩɺ���3y�,q*�+A���W���m��iӌ�,����5��񶬻)��N[��w~˻�ջmf߻�+黀��?[�������x ����a$�����kA"���&���*��.��3��7��;��?��C���F��J��N��VR�V���Y�'l]��a��d��1h���k��7o���r�p v�.�y���|�;%���Ё�Yy��!��e�c��N��A���7���Ύ��d����������\��R����7��ę�
O���؜��a��N韼p�� ���Y{���������w������`��􏭼A��r������֘��?������� ������*'��:����/���  �  ?gN=K�M=��L=$L=�XK=�J=��I=�I=PBH={G=�F=l�E=� E=�VD=A�C=�B=��A=�#A=*T@=��?=�>=��==�
==5<=�];=l�:=R�9=��8=B�7=,7=I26=�O5=�j4=+�3=s�2=��1=��0=$�/=s�.=W�-=��,=��+=�+=2*=�)=��'=��&=x�%=I�$=��#=g�"=��!=i� =�m=�L=:(= =N�=֤=�q=�:=��=N�=�~={8=8�= �=�M=��=ĝ=�?
=��='x=z=�=�/=t�=�A =���<x��<ԁ�< s�<{]�<A�<��<[��<r��<]��<JR�<[�<���<�{�<|)�< ��<�u�<��<���<�E�<ؼ<ef�<�<Dx�<I��<4}�<S��<�v�<��<�f�<�ۙ<�N�<R��<z0�<}��<��<�z�<��<D�z<�s<�Yl<j3e<�^<��V<��O<w�H<�A<�o:<�X3<�E,<:7%<G-<m(<)<�/	<�<<���;��;��;�o�;տ;�K�;դ;q�;!�;!�y;�~_;�^E;�k+;	�;+)�:�d�:��:� 2:�9���E#鹬U��R����ɺ����Ny�
q*�W+A��W�K�m���fӌ�O����5��������[��T~˻�ջnf߻�+黺��[�������p ����X$������A"���&���*��.��3��7�x;��?��C���F��J��N��VR��V���Y�*l]��a��d��1h���k��7o���r�W v�7�y���|�C%���Ё�Zy��,��X�c��I��I���7���Ύ��d����������N��T����7��ę�O���؜��a��H韼p�����X{����������������j��쏭�;��{������ޘ��>������� ������''��.����/���  �  EgN=F�M=��L=%L=�XK=�J=��I=�I=LBH={G=#�F=l�E=� E=�VD=D�C= �B=��A=�#A=-T@=��?=�>=��==�
==5<=�];=q�:=U�9=��8=H�7=)7=J26=�O5=�j4=,�3=r�2=��1=}�0=(�/=q�.=U�-=��,=��+=�+=-*=�)=��'=��&=x�%=J�$=��#=c�"=��!=g� =�m=�L=:(= =G�=֤=�q=�:=��=R�=�~=y8=:�=��=�M=��=Ɲ=�?
=��=&x=w=��=�/=w�=�A =��<��<́�<$s�<t]�<A�<��<[��<}��<V��<RR�<S�<���<�{�<})�<%��<�u�<��<y��<�E�<ؼ<]f�<�<Ix�<R��<*}�<]��<�v�<��<�f�<�ۙ<�N�<F��<�0�<|��<��<�z�<��<R�z<�s<�Yl<`3e<�^<��V<n�O<x�H<�A<�o:<�X3<�E,<@7%<:-<u(<)<�/	<�<<���;<��;��;�o�;�Կ; L�;�Ԥ;q�;� �;U�y;�~_;p^E;5l+;§;�)�:|d�:=�:r!2:c�9�����$�aU��S����ɺ����^y��p*�~+A�ϧW�m�m���xӌ�G���b5��@�������[��L~˻�ջff߻�+�����Z�������� ����S$�0�����A"���&�Ƽ*��.��3��7�n;��?��C���F���J��N��VR��V���Y�l]��a�ۢd��1h���k��7o���r�Q v�C�y�y�|�D%���Ё�Oy��3��P�c��D��I���7���Ύ��d������͊��H��Z����7��ę�O���؜��a��>韼p�����\{�����������������k��폭�F��{������㘳�,������� ������3'��-����/���  �  ?gN=H�M=��L='L=�XK=�J=��I=�I=QBH={G=#�F=n�E=� E=�VD=<�C=�B=��A=�#A=*T@=��?=�>=��==�
==5<=�];=q�:=T�9=��8=C�7=+7=I26=�O5=�j4=0�3=o�2=��1=��0=%�/=w�.=T�-=��,=��+=�+=/*=�)=��'=��&=z�%=J�$=��#=i�"=��!=j� =�m=�L=9(= =K�=ؤ=�q=�:=��=T�=�~={8=6�=�=�M=��=ĝ=�?
=��=%x=}=�=�/=q�=�A =���<���<ׁ�<s�<v]�<A�<��<]��<z��<^��<HR�<Z�<���<�{�<})�<��<�u�<��<���<�E�<	ؼ<cf�<�<Lx�<B��<7}�<V��<�v�<��<�f�<�ۙ<�N�<J��<y0�<~��<��<�z�<��<N�z<�s<�Yl<X3e<�^<��V<y�O<x�H<�A<�o:<�X3<�E,<G7%<I-<r(<)<�/	<�<<���;@��;�;�o�;տ;�K�;�Ԥ;2q�;%!�;�y;�~_;�^E;)l+;��;)�:�d�:4�:U!2:h�9͖��$鹙U��R����ɺ����y�:q*�W+A���W��m��dӌ�L����5��/�����i[��]~˻��ջbf߻�+黬��[�����߈�z ����_$� ����|A"���&���*��.��3��7�};��?��C���F��J���N��VR��V���Y�"l]��a���d��1h���k��7o���r�\ v�?�y���|�C%���Ё�Ry��+��Z�	c��D��E���7���Ύ��d��������U��S����7��ę�O���؜��a��E韼p�����W{�����������������i��ꏭ�D��s������☳�>����� ������.'��-����/���  �  <gN=O�M=��L=$L=�XK=�J=��I=�I=SBH={G=%�F=k�E=� E=�VD=<�C=�B=��A=�#A=+T@=��?=�>=��==�
==
5<=�];=j�:=V�9=��8=>�7=.7=F26=�O5=�j4=.�3=t�2=��1=��0= �/=v�.=T�-=��,=��+=�+=7*=�)=��'=��&={�%=J�$=��#=k�"=��!=l� =�m=�L=;(= =O�=Ф=�q=�:=��=M�=�~=8=0�=�=�M=��=ĝ=�?
=��=$x=}=�=�/=s�=�A =���<r��<؁�<s�<]�<�@�<��<b��<l��<]��<@R�<g�<���<�{�<�)�<��<�u�<��<���<�E�<ؼ<af�<�<Ox�<C��<<}�<I��<�v�<��<�f�<�ۙ<�N�<Z��<u0�<}��<��<�z�<��<B�z<�s<�Yl<x3e<�^<��V<��O<q�H<�A<�o:<�X3<�E,<87%<@-<l(<()<�/	<�<<���;M��;��;�o�;'տ;�K�;*դ;�p�;!�;7�y;_;�^E;�k+;g�;�(�:�d�:j�:�!2:��95���G"�nU��R��D�ɺF���9y�%q*��*A�M�W��m��Pӌ�^����5��񶬻0��r[���~˻�ջ`f߻,默��[��������q ����Y$���)��qA"���&���*�!�.��3��7��;��?��C���F��J��N��VR��V���Y�:l]��a��d��1h���k��7o���r�e v�/�y���|�@%���Ё�_y��,��b��b��M��K���7���Ύ��d����������V��M����7��!ę�O���؜��a��R韼p�����]{����������y������j��鏭�A��y������՘��>������� ������*'��1����/���  �  CgN=G�M=��L=&L=�XK=�J=��I=�I=QBH={G=#�F=p�E=� E=�VD=<�C=�B=��A=�#A=*T@=��?=�>=��==�
==5<=�];=o�:=V�9=��8=E�7=,7=F26=�O5=�j4=.�3=r�2=��1=��0=(�/=u�.=T�-=��,=��+=�+=0*=�)=��'=��&=x�%=J�$=��#=g�"=��!=l� =�m=�L=8(= =M�=֤=�q=�:=��=Q�=�~=z8=6�=�=�M=��=Ɲ=�?
=��=%x=z=��=�/=r�=�A =��<��<ԁ�<s�<y]�<A�<��<a��<w��<b��<KR�<W�<���<�{�<�)�<��<�u�<��<���<�E�<ؼ<df�<�<Mx�<I��<5}�<R��<�v�<��<�f�<�ۙ<�N�<K��<�0�<}��<��<�z�<��<Y�z<�s<�Yl<b3e<�^<��V<z�O<i�H<�A<�o:<�X3<�E,<@7%<P-<n(<)<�/	<�<<���;>��;�;�o�;�Կ;�K�;�Ԥ;q�;/!�;"�y;�~_;�^E;�k+;�;V)�:Ee�:��:�!2:��99����#�cU��R����ɺ@���ay�q*�V+A�ȧW�,�m��hӌ�<���m5��"�����v[��X~˻�ջgf߻�+黷��[�����ވ�q ����b$�����rA"���&���*��.��3��7�;��?��C���F���J��N��VR��V���Y�l]��a��d��1h���k��7o���r�` v�:�y��|�C%���Ё�Uy��'��W�c��K��F���7���Ύ��d��������X��Z����7��ę�O���؜��a��I韼p�����S{�����������������j������D��v������☳�>������� ������-'��5����/���  �  FgN=G�M=��L="L=�XK= �J=��I=�I=OBH={G= �F=m�E=� E=�VD=E�C=�B=��A=�#A=*T@=��?=�>=��==�
==5<=�];=m�:=U�9=��8=I�7=%7=N26=�O5=�j4=+�3=o�2=��1=z�0=&�/=p�.=Y�-=��,=��+=�+=-*=�)=��'=��&=v�%=J�$=��#=f�"=��!=g� =�m=�L=<(= =I�=ؤ=�q=�:=��=S�=�~=x8=:�=��=�M=��=Ɲ=�?
=��=*x=v=�=�/=v�=�A =��<{��<ρ�<)s�<m]�<A�<��<^��<x��<V��<QR�<S�<���<�{�<z)�<��<�u�<��<��<�E�<	ؼ<^f�<�<Cx�<J��<1}�<]��<�v�<��<�f�<�ۙ<�N�<F��<�0�<v��<��<�z�<��<J�z<�s<�Yl<O3e<�^<��V<~�O<��H<��A<�o:<�X3<�E,<07%<K-<x(<	)<�/	<�<<���;"��; �;�o�; տ;L�;�Ԥ;'q�;!�;#�y;�~_;�^E;8l+;ͧ;�)�:�d�:��:�!2:��9Ћ��'�fU�;S���ɺ�����y��p*��+A��W�y�m���vӌ�O���m5��<�������[��C~˻�ջcf߻�+�����Z�����܈�� ����N$�(��	���A"���&���*�
�.��3��7�n;��?��C���F���J���N��VR��V���Y�!l]��a�ߢd��1h���k��7o���r�E v�R�y�{�|�C%���Ё�Sy��3��Q�c��A��F���7���Ύ��d������Ɗ��F��S����7��ę�O���؜��a��>韼p�����S{������򃧼�������q��菭�>��~������옳�-��Ɲ��� ������+'��)����/���  �  @gN=K�M=��L=%L=�XK=�J=��I=�I=QBH={G=&�F=l�E=� E=�VD==�C=�B=��A=�#A=/T@=��?=�>=��==�
==
5<=�];=n�:=T�9=��8=C�7=*7=I26=�O5=�j4=0�3=q�2=��1=��0=&�/=s�.=U�-=��,=��+=�+=1*=�)=��'=��&=x�%=J�$=��#=i�"=��!=j� =�m=�L=;(= =K�=Ԥ=�q=�:=��=O�=�~={8=4�= �=�M=��=Ý=�?
=��=&x=y=�=�/=t�=�A =���<z��<Ё�<s�<v]�<A�<��<]��<x��<[��<BR�<]�<���<�{�<~)�<$��<�u�<��<���<�E�<ؼ<Zf�<�<Nx�<H��<8}�<Q��<�v�<��<�f�<�ۙ<�N�<O��<{0�<}��<��<�z�<��<P�z<�s<�Yl<f3e<�^<��V<n�O<u�H<�A<�o:<�X3<�E,<?7%<B-<`(<)<�/	<�<<���;Q��;��;�o�;տ;�K�;դ;	q�;!�;n�y;�~_;�^E;�k+;#�;�(�:�d�:��:O!2:��9�����$鹛U�bS���ɺ	���ky��p*�:+A��W�P�m���nӌ�U���5�������z[��l~˻
�ջdf߻�+黪�� [�������| ����Y$�����~A"���&���*��.��3��7��;��?��C���F��J��N��VR��V���Y�#l]��a��d��1h���k��7o���r�\ v�?�y���|�D%���Ё�Ty��.��`�c��J��G���7���Ύ��d����������S��P����7��ę�O���؜��a��J韼p�����[{�����������������j��폭�F��{������ޘ��5������� ������3'��/����/���  �  <gN=L�M=��L='L=�XK=�J=��I=�I=VBH={G=%�F=o�E=� E=�VD=<�C=�B=��A=�#A=+T@=��?=��>=��==�
==	5<= ^;=m�:=P�9=��8=A�7=27=C26=�O5=�j4=-�3=r�2=��1=��0=#�/=x�.=Q�-=��,=��+=�+=2*=�)=��'=��&=}�%=M�$=��#=k�"=��!=o� =�m=�L=:(= =P�=դ=�q=�:=��=R�=�~=�8=3�=�=�M=��=Ý=�?
=��= x==�=�/=p�=�A =��<z��<܁�<s�<�]�<A�<��<W��<q��<h��<AR�<h�<���<�{�<|)�<��<�u�<��<���<�E�<ؼ<cf�<�<Qx�<<��<?}�<M��<�v�<��<�f�<�ۙ<�N�<S��<t0�<���<��<�z�<��<F�z<�s<�Yl<g3e<�^<��V<z�O<h�H<&�A<�o:<�X3<�E,<E7%<O-<e(<-)<�/	<�<<q��;L��;�;�o�;0տ;�K�; դ;q�;7!�;1�y;�~_;�^E;�k+;u�;�(�:�e�:��:b 2:��9>���* ��U��R����ɺt���\y�Lq*�H+A�#�W���m�!�Uӌ�=����5�����:��N[��m~˻܁ջMf߻�+黗��/[�������k ����\$�����fA"���&���*��.��3��7��;��?��C���F��J���N��VR�V���Y�0l]��a���d��1h���k��7o���r�u v�!�y���|�C%���Ё�Zy�� ��a��b��O��>���7���Ύ��d����������V��K����7��ę�O���؜��a��N韼p�����W{����������������`������F��r������ݘ��F������� ������-'��5����/���  �  AgN=N�M=��L=&L=�XK=�J=��I=�I=TBH={G=#�F=k�E=� E=�VD=A�C=�B=��A=�#A=,T@=��?=�>=��==�
==5<=�];=m�:=V�9=��8=D�7=,7=E26=�O5=�j4=-�3=t�2=��1=��0=#�/=u�.=R�-=��,=��+=�+=4*=�)=��'=��&=y�%=H�$=��#=j�"=��!=i� =�m=�L=;(= =K�=Ԥ=�q=�:=��=S�=�~={8=3�= �=�M=��=Ɲ=�?
=��=!x=|=�=�/=v�=�A =��<w��<ց�<s�<{]�<A�<��<a��<w��<[��<DR�<]�<���<�{�<�)�<��<�u�<��<���<�E�<ؼ<af�<�<Ix�<I��<;}�<Q��<�v�<��<�f�<�ۙ<�N�<V��<}0�<|��<��<�z�<��<F�z<
�s<�Yl<f3e<�^<��V<x�O<l�H<�A<�o:<�X3<�E,<@7%<?-<l(<)<�/	<�<<���;>��;��;�o�;տ;�K�;�Ԥ;q�;	!�;>�y;_;�^E;�k+;�;�(�:�d�:��:�!2:R�9<����#鹀U��R����ɺc���<y��p*�P+A��W�$�m��`ӌ�R���r5�������x[��z~˻��ջsf߻�+黠���Z�������{ ����W$�!�����A"���&���*��.��3��7��;��?��C���F���J���N��VR�V���Y�.l]��a�ߢd��1h���k��7o���r�i v�5�y���|�=%���Ё�Uy��.��^�c��N��A���7���Ύ��d������Ċ��N��T����7�� ę�O���؜��a��J韼p�����^{����������}������k��폭�E��w������ߘ��2������� ������.'��3����/���  �  BgN=D�M=��L='L=�XK=!�J=��I=�I=LBH={G="�F=l�E=� E=�VD=A�C=�B=��A=�#A=-T@=��?=�>=��==�
==5<=�];=o�:=S�9=��8=E�7=)7=K26=�O5=�j4=1�3=l�2=��1=~�0='�/=s�.=T�-=��,=��+=�+=,*=�)=��'=��&=|�%=G�$=��#=d�"=��!=e� =�m=�L=;(= =L�=ۤ=�q=�:=��=O�=�~=}8=8�=��=�M=��=ĝ=�?
=��=$x=x=��=�/=p�=�A =���<{��<́�<!s�<x]�<A�<��<W��<z��<W��<PR�<Z�<���<�{�<�)�<%��<�u�<��<~��<�E�<ؼ<kf�<�<Fx�<O��<,}�<T��<�v�<��<�f�<�ۙ<�N�<C��<�0�<y��<��<�z�<��<X�z<�s<�Yl<J3e<�^<��V<l�O<|�H<�A<�o:<�X3<�E,<E7%<F-<~(<)<�/	<�<<���;6��;��;�o�;�Կ;�K�;�Ԥ;Rq�;� �;Y�y;!_;G^E;�k+; �;�)�:�d�:��:!2:�9s����$�U��S��ݩɺ�����y�"q*�p+A�קW�L�m��Rӌ�I���r5��G������[��N~˻�ջwf߻�+�����Z�����Ԉ�o ����X$�������A"���&�ü*��.��3��7�u;��?��C���F��J���N��VR��V���Y�l]��a���d��1h���k��7o���r�U v�<�y���|�J%���Ё�Qy��1��Q�	c��J��O���7���Ύ��d������Ǌ��N��Y����7��ę�O���؜��a��G韼 p�����X{�����������������n��班�G��z������똳�:��ɝ�� ������4'��+����/���  �  AgN=N�M=��L=&L=�XK=�J=��I=�I=TBH={G=#�F=k�E=� E=�VD=A�C=�B=��A=�#A=,T@=��?=�>=��==�
==5<=�];=m�:=V�9=��8=D�7=,7=E26=�O5=�j4=-�3=t�2=��1=��0=#�/=u�.=R�-=��,=��+=�+=4*=�)=��'=��&=y�%=H�$=��#=j�"=��!=i� =�m=�L=;(= =K�=Ԥ=�q=�:=��=S�=�~={8=3�= �=�M=��=Ɲ=�?
=��=!x=|=�=�/=v�=�A =��<w��<ց�<s�<{]�<A�<��<a��<w��<[��<DR�<]�<���<�{�<�)�<��<�u�<��<���<�E�<ؼ<af�<�<Ix�<I��<;}�<Q��<�v�<��<�f�<�ۙ<�N�<V��<}0�<|��<��<�z�<��<F�z<
�s<�Yl<f3e<�^<��V<x�O<l�H<�A<�o:<�X3<�E,<@7%<?-<l(<)<�/	<�<<���;>��;��;�o�;տ;�K�;�Ԥ;q�;	!�;>�y;_;�^E;�k+;�;�(�:�d�:��:�!2:Q�9?����#鹁U��R����ɺc���<y��p*�P+A��W�$�m��`ӌ�R���r5�������x[��z~˻��ջsf߻�+黠���Z�������{ ����W$�!�����A"���&���*��.��3��7��;��?��C���F���J���N��VR�V���Y�.l]��a�ߢd��1h���k��7o���r�h v�5�y���|�=%���Ё�Uy��.��^�c��N��A���7���Ύ��d������Ċ��N��T����7�� ę�O���؜��a��J韼p�����^{����������}������k��폭�E��w������ߘ��2������� ������.'��3����/���  �  <gN=L�M=��L='L=�XK=�J=��I=�I=VBH={G=%�F=o�E=� E=�VD=<�C=�B=��A=�#A=+T@=��?=��>=��==�
==	5<= ^;=m�:=P�9=��8=A�7=27=C26=�O5=�j4=-�3=r�2=��1=��0=#�/=x�.=Q�-=��,=��+=�+=2*=�)=��'=��&=}�%=M�$=��#=k�"=��!=o� =�m=�L=:(= =P�=դ=�q=�:=��=R�=�~=�8=3�=�=�M=��=Ý=�?
=��= x==�=�/=p�=�A =��<z��<܁�<s�<�]�<A�<��<W��<q��<h��<AR�<h�<���<�{�<|)�<��<�u�<��<���<�E�<ؼ<cf�<�<Qx�<<��<?}�<M��<�v�<��<�f�<�ۙ<�N�<S��<t0�<���<��<�z�<��<F�z<�s<�Yl<g3e<�^<��V<z�O<h�H<&�A<�o:<�X3<�E,<E7%<O-<e(<-)<�/	<�<<q��;L��;�;�o�;0տ;�K�; դ;q�;7!�;1�y;�~_;�^E;�k+;u�;�(�:�e�:��:a 2:��9B���+ ��U��R����ɺt���\y�Mq*�H+A�#�W���m�!�Uӌ�=����5�����:��N[��m~˻݁ջMf߻�+黗��/[�������k ����\$�����fA"���&���*��.��3��7��;��?��C���F��J���N��VR�V���Y�0l]��a���d��1h���k��7o���r�u v�!�y���|�C%���Ё�Zy�� ��a��b��O��>���7���Ύ��d����������V��K����7��ę�O���؜��a��N韼p�����W{����������������`������F��r������ݘ��F������� ������-'��5����/���  �  @gN=K�M=��L=%L=�XK=�J=��I=�I=QBH={G=&�F=l�E=� E=�VD==�C=�B=��A=�#A=/T@=��?=�>=��==�
==
5<=�];=n�:=T�9=��8=C�7=*7=I26=�O5=�j4=0�3=q�2=��1=��0=&�/=s�.=U�-=��,=��+=�+=1*=�)=��'=��&=x�%=J�$=��#=i�"=��!=j� =�m=�L=;(= =K�=Ԥ=�q=�:=��=O�=�~={8=4�= �=�M=��=Ý=�?
=��=&x=y=�=�/=t�=�A =���<z��<Ё�<s�<v]�<A�<��<]��<x��<[��<CR�<]�<���<�{�<~)�<$��<�u�<��<���<�E�<ؼ<Zf�<�<Nx�<H��<8}�<Q��<�v�<��<�f�<�ۙ<�N�<O��<{0�<}��<��<�z�<��<P�z<�s<�Yl<f3e<�^<��V<n�O<u�H<�A<�o:<�X3<�E,<?7%<B-<`(<)<�/	<�<<���;Q��;��;�o�;տ;�K�;դ;	q�;!�;m�y;�~_;�^E;�k+;#�;�(�:�d�:��:N!2:��9�����$鹜U�cS���ɺ
���ky��p*�:+A��W�P�m���nӌ�V���5�������z[��l~˻
�ջdf߻�+黪�� [�������| ����Y$�����~A"���&���*��.��3��7��;��?��C���F��J��N��VR��V���Y�#l]��a��d��1h���k��7o���r�\ v�?�y���|�D%���Ё�Ty��.��`�c��J��G���7���Ύ��d����������S��P����7��ę�O���؜��a��J韼p�����[{�����������������j��폭�F��{������ޘ��5������� ������3'��/����/���  �  FgN=G�M=��L="L=�XK= �J=��I=�I=OBH={G= �F=m�E=� E=�VD=E�C=�B=��A=�#A=*T@=��?=�>=��==�
==5<=�];=m�:=U�9=��8=I�7=%7=N26=�O5=�j4=+�3=o�2=��1=z�0=&�/=p�.=Y�-=��,=��+=�+=-*=�)=��'=��&=v�%=J�$=��#=f�"=��!=g� =�m=�L=<(= =I�=ؤ=�q=�:=��=S�=�~=x8=:�=��=�M=��=Ɲ=�?
=��=*x=v=�=�/=v�=�A =��<{��<ρ�<)s�<m]�<A�<��<^��<x��<V��<QR�<S�<���<�{�<z)�<��<�u�<��<��<�E�<	ؼ<^f�<�<Cx�<J��<1}�<]��<�v�<��<�f�<�ۙ<�N�<F��<�0�<v��<��<�z�<��<J�z<�s<�Yl<O3e<�^<��V<~�O<��H<��A<�o:<�X3<�E,<07%<K-<x(<	)<�/	<�<<���;"��; �;�o�; տ;L�;�Ԥ;'q�;!�;#�y;�~_;�^E;8l+;ͧ;�)�:�d�:��:�!2:��9ً��'�gU�<S���ɺ�����y��p*��+A��W�y�m���vӌ�O���m5��<�������[��C~˻�ջcf߻�+�����Z�����܈�� ����N$�(��	���A"���&���*�
�.��3��7�n;��?��C���F���J���N��VR��V���Y�!l]��a�ߢd��1h���k��7o���r�E v�R�y�{�|�C%���Ё�Sy��3��Q�c��A��F���7���Ύ��d������Ɗ��F��S����7��ę�O���؜��a��>韼p�����S{������򃧼�������q��菭�>��~������옳�-��Ɲ��� ������+'��)����/���  �  CgN=G�M=��L=&L=�XK=�J=��I=�I=QBH={G=#�F=p�E=� E=�VD=<�C=�B=��A=�#A=*T@=��?=�>=��==�
==5<=�];=o�:=V�9=��8=E�7=,7=F26=�O5=�j4=.�3=r�2=��1=��0=(�/=u�.=T�-=��,=��+=�+=0*=�)=��'=��&=x�%=J�$=��#=g�"=��!=l� =�m=�L=8(= =M�=֤=�q=�:=��=Q�=�~=z8=6�=�=�M=��=Ɲ=�?
=��=%x=z=��=�/=r�=�A =��<��<ԁ�<s�<y]�<A�<��<a��<w��<b��<KR�<X�<���<�{�<�)�<��<�u�<��<���<�E�<ؼ<df�<�<Mx�<I��<5}�<R��<�v�<��<�f�<�ۙ<�N�<K��<�0�<}��<��<�z�<��<Y�z<�s<�Yl<b3e<�^<��V<z�O<i�H<�A<�o:<�X3<�E,<@7%<P-<n(<)<�/	<�<<���;>��;�;�o�;�Կ;�K�;�Ԥ;q�;/!�;"�y;�~_;�^E;�k+;�;V)�:Ee�:��:�!2:��9A����#�dU��R����ɺA���by�q*�V+A�ȧW�,�m��hӌ�<���n5��"�����v[��X~˻�ջgf߻�+黸��[�����ވ�q ����b$�����rA"���&���*��.��3��7�;��?��C���F���J��N��VR��V���Y�l]��a��d��1h���k��7o���r�` v�:�y��|�C%���Ё�Uy��'��W�c��K��F���7���Ύ��d��������X��Z����7��ę�O���؜��a��I韼p�����S{�����������������j������D��v������☳�>������� ������-'��5����/���  �  <gN=O�M=��L=$L=�XK=�J=��I=�I=SBH={G=%�F=k�E=� E=�VD=<�C=�B=��A=�#A=+T@=��?=�>=��==�
==
5<=�];=j�:=V�9=��8=>�7=.7=F26=�O5=�j4=.�3=t�2=��1=��0= �/=v�.=T�-=��,=��+=�+=7*=�)=��'=��&={�%=J�$=��#=k�"=��!=l� =�m=�L=;(= =O�=Ф=�q=�:=��=M�=�~=8=0�=�=�M=��=ĝ=�?
=��=$x=}=�=�/=s�=�A =���<r��<؁�<s�<]�<�@�<��<b��<l��<]��<@R�<g�<���<�{�<�)�<��<�u�<��<���<�E�<ؼ<af�<�<Ox�<C��<<}�<I��<�v�<��<�f�<�ۙ<�N�<Z��<u0�<}��<��<�z�<��<B�z<�s<�Yl<x3e<�^<��V<��O<q�H<�A<�o:<�X3<�E,<87%<@-<l(<()<�/	<�<<���;M��;��;�o�;'տ;�K�;*դ;�p�;!�;7�y;_;�^E;�k+;g�;�(�:�d�:i�:�!2:��9>���J"�oU��R��E�ɺF���9y�%q*��*A�M�W��m��Pӌ�^����5��񶬻0��r[���~˻�ջ`f߻,默��[��������q ����Y$���)��qA"���&���*�!�.��3��7��;��?��C���F��J��N��VR��V���Y�:l]��a��d��1h���k��7o���r�e v�/�y���|�@%���Ё�_y��,��b��b��M��K���7���Ύ��d����������V��M����7��!ę�O���؜��a��R韼p�����]{����������y������j��鏭�A��y������՘��>������� ������*'��1����/���  �  ?gN=H�M=��L='L=�XK=�J=��I=�I=QBH={G=#�F=n�E=� E=�VD=<�C=�B=��A=�#A=*T@=��?=�>=��==�
==5<=�];=q�:=T�9=��8=C�7=+7=I26=�O5=�j4=0�3=o�2=��1=��0=%�/=w�.=T�-=��,=��+=�+=/*=�)=��'=��&=z�%=J�$=��#=i�"=��!=j� =�m=�L=9(= =K�=ؤ=�q=�:=��=T�=�~={8=6�=�=�M=��=ĝ=�?
=��=%x=}=�=�/=q�=�A =���<���<ׁ�<s�<v]�<A�<��<]��<z��<^��<HR�<Z�<���<�{�<})�<��<�u�<��<���<�E�<	ؼ<cf�<�<Lx�<B��<7}�<V��<�v�<��<�f�<�ۙ<�N�<J��<y0�<~��<��<�z�<��<N�z<�s<�Yl<X3e<�^<��V<y�O<x�H<�A<�o:<�X3<�E,<G7%<I-<r(<)<�/	<�<<���;@��;�;�o�;տ;�K�;�Ԥ;2q�;%!�;�y;�~_;�^E;(l+;��;)�:�d�:3�:T!2:e�9ז�� $鹛U��R����ɺ����y�:q*�W+A���W��m��dӌ�L����5��/�����i[��]~˻��ջbf߻�+黬��[�����߈�z ����_$� ����|A"���&���*��.��3��7�};��?��C���F��J���N��VR��V���Y�"l]��a���d��1h���k��7o���r�\ v�?�y���|�C%���Ё�Ry��+��Z�	c��D��E���7���Ύ��d��������U��S����7��ę�O���؜��a��E韼p�����W{�����������������i��ꏭ�D��s������☳�>����� ������.'��-����/���  �  EgN=F�M=��L=%L=�XK=�J=��I=�I=LBH={G=#�F=l�E=� E=�VD=D�C= �B=��A=�#A=-T@=��?=�>=��==�
==5<=�];=q�:=U�9=��8=H�7=)7=J26=�O5=�j4=,�3=r�2=��1=}�0=(�/=q�.=U�-=��,=��+=�+=-*=�)=��'=��&=x�%=J�$=��#=c�"=��!=g� =�m=�L=:(= =G�=֤=�q=�:=��=R�=�~=y8=:�=��=�M=��=Ɲ=�?
=��=&x=w=��=�/=w�=�A =��<��<́�<$s�<t]�<A�<��<[��<}��<V��<SR�<S�<���<�{�<})�<%��<�u�<��<y��<�E�<ؼ<]f�<�<Ix�<R��<*}�<]��<�v�<��<�f�<�ۙ<�N�<F��<�0�<|��<��<�z�<��<R�z<�s<�Yl<`3e<�^<��V<n�O<x�H<�A<�o:<�X3<�E,<@7%<:-<u(<)<�/	<�<<���;<��;��;�o�;�Կ; L�;�Ԥ;q�;� �;U�y;�~_;o^E;5l+;§;�)�:|d�:<�:p!2:b�9�����$�bU��S����ɺ����_y��p*�~+A�ϧW�m�m���xӌ�G���b5��@�������[��L~˻�ջff߻�+�����Z�������� ����S$�0�����A"���&�Ƽ*��.��3��7�n;��?��C���F���J��N��VR��V���Y�l]��a�ۢd��1h���k��7o���r�Q v�C�y�y�|�D%���Ё�Oy��3��P�c��D��I���7���Ύ��d������͊��H��Z����7��ę�O���؜��a��>韼p�����\{�����������������k��폭�F��{������㘳�,������� ������3'��-����/���  �  ?gN=K�M=��L=$L=�XK=�J=��I=�I=PBH={G=�F=l�E=� E=�VD=A�C=�B=��A=�#A=*T@=��?=�>=��==�
==5<=�];=l�:=R�9=��8=B�7=,7=I26=�O5=�j4=+�3=s�2=��1=��0=$�/=s�.=W�-=��,=��+=�+=2*=�)=��'=��&=x�%=I�$=��#=g�"=��!=i� =�m=�L=:(= =N�=֤=�q=�:=��=N�=�~={8=8�= �=�M=��=ĝ=�?
=��='x=z=�=�/=t�=�A =���<x��<ԁ�< s�<{]�<A�<��<[��<r��<]��<JR�<[�<���<�{�<|)�< ��<�u�<��<���<�E�<ؼ<ef�<�<Dx�<I��<4}�<S��<�v�<��<�f�<�ۙ<�N�<R��<z0�<}��<��<�z�<��<D�z<�s<�Yl<j3e<�^<��V<��O<w�H<�A<�o:<�X3<�E,<:7%<G-<m(<)<�/	<�<<���;��;��;�o�;տ;�K�;դ;q�;!�;!�y;�~_;�^E;�k+;	�;*)�:�d�:��:� 2:
�9����G#鹬U��R����ɺ����Ny�
q*�X+A��W�K�m���fӌ�O����5��������[��T~˻�ջnf߻�+黺��[�������p ����X$������A"���&���*��.��3��7�x;��?��C���F��J��N��VR��V���Y�*l]��a��d��1h���k��7o���r�W v�7�y���|�C%���Ё�Zy��,��X�c��I��I���7���Ύ��d����������N��T����7��ę�O���؜��a��H韼p�����X{����������������j��쏭�;��{������ޘ��>������� ������''��.����/���  �  <gN=P�M=��L=(L=�XK=�J=��I=�I=XBH={G=$�F=o�E=� E=�VD=8�C=�B=��A=�#A=(T@=��?=��>=��==�
==5<=�];=m�:=V�9=��8=A�7=/7=C26=�O5=�j4=/�3=u�2=��1=��0=%�/=z�.=R�-=��,=��+=�+=7*=�)=��'=��&=v�%=I�$=��#=n�"=��!=n� =�m=�L=9(= =L�=Ӥ=�q=�:=��=P�=�~=z8=2�=�=�M=��=ŝ=�?
=��="x=�=�=�/=r�=�A =���<{��<݁�<s�<]�<A�<��<f��<s��<i��<=R�<^�<���<�{�<�)�<��<�u�<��<���<�E�<
ؼ<^f�<�<Qx�<?��<E}�<M��<�v�<��<�f�<�ۙ<�N�<[��<t0�<���<��<�z�<��<G�z<�s<�Yl<y3e<�^<��V<�O<`�H< �A<�o:<�X3<�E,<K7%<I-<U(<)<�/	<�<<���;D��;�;�o�;տ;�K�;դ;q�;7!�;�y;�~_;�^E;�k+;%�;I(�:�e�:��:�!2:��9ܚ���!�+U��R��ǩɺ���3y�,q*�+A���W���m��jӌ�,����5��񶬻)��N[��w~˻�ջmf߻�+黀��?[�������x ����a$�����kA"���&���*��.��3��7��;��?��C���F��J��N��VR�V���Y�'l]��a��d��1h���k��7o���r�p v�.�y���|�;%���Ё�Yy��!��e�c��N��A���7���Ύ��d����������\��R����7��ę�
O���؜��a��N韼p�� ���Y{���������w������`��􏭼A��r������֘��?������� ������*'��:����/���  �  >gN=J�M=��L=$L=�XK=�J=��I=�I=QBH={G=#�F=m�E=� E=�VD=B�C=�B=��A=�#A=)T@=��?=�>=��==�
==5<=�];=k�:=V�9=��8=D�7=-7=I26=�O5=�j4=.�3=q�2=��1=~�0=%�/=r�.=U�-=��,=��+=�+=1*=�)=��'=��&={�%=M�$=��#=j�"=��!=l� =�m=�L==(= =K�=Ӥ=�q=�:=��=P�=�~=~8=7�= �=�M=��==�?
=��=&x=y=�=�/=t�=�A =��<x��<ҁ�<!s�<|]�<
A�<��<`��<o��<_��<JR�<b�<���<�{�<)�<��<�u�<��<���<�E�<ؼ<`f�<�<Lx�<B��<7}�<U��<�v�<��<�f�<�ۙ<�N�<P��<w0�<���<��<�z�<��<J�z<�s<�Yl<c3e<�^<��V<{�O<w�H<�A<�o:<�X3<�E,<87%<F-<p(<()<�/	<�<<���;;��;�;�o�;տ;�K�;�Ԥ;q�;!�;�y;�~_;�^E;�k+;F�; )�:e�:q�:�!2:��9�����"鹆U�4S��)�ɺW���iy��p*�p+A��W�[�m��Yӌ�6����5����� ���[��\~˻�ջOf߻�+黡��&[�������{ ����P$�����uA"���&���*��.��3��7�|;��?��C���F��J��N��VR��V���Y�(l]��a��d��1h���k��7o���r�V v�5�y���|�E%���Ё�\y��+��X�c��G��H���7���Ύ��d����������K��O����7��ę�O���؜��a��G韼p�����Z{�����������������d��鏭�@��|������☳�3������� ������-'��.����/���  �  �eN=��M=�L=L=�VK=w�J=��I=�I=�>H=swG=8�F=7�E=nE=�QD=.�C=��B=)�A=�A=�M@=}?=�>=��====-<=�U;=�|:=P�9=:�8=w�7=�7=�'6=�D5=_4=hx3=>�2=��1=t�0=��/=��.=�-=��,=[�+=�*=*�)=o�(=��'=N�&=��%=1�$=|�#=��"=]�!=�w =�Y=�8=�=/�=$�=k�=�[=�$=��=$�=�h="=��=q�=J7=7�=8�=S)
=��=�a=_�=�=�=�=g, =;`�<p`�<mY�<�K�<�6�<�<���<6��<?��<$l�<1�<1��<é�<�]�<��<|��<T[�<���<[��<�.�<L¼<�Q�<�ݵ<Hf�<��<�m�<"�<�i�<�<Q\�<tҙ<�F�<���<+�<H��<�
�<0y�<>�<��z<�s<�`l<n<e<�^<��V<	�O<��H<��A<��:<fs3<�b,<�V%<4O<�L<�O<	Y	<Mh<���;=7�;���;"��;D�;t��;<M�;�;I��;��z;�`;�zF;��,;K�;���:Aܿ:K��:�H7:w��9͛]�B޹҆O�*�����ƺ����U���(���?�J*V�gl�[2��%���Җ��s��W����W������3�ʻ��Իa�޻o軗򻔡����S.���aQ�~���;������!�m4&�-m*�!�.���2�:�6���:���>�i�B�2�F�X�J�RN��R���U�(�Y�H3]���`��md�5�g�ˆk��o�@�r���u�_y���|�C��}����f��m��_����R����W����(��2����W��@쑼��F��ܟ���-��ʺ��JF���М��Y��⟼{i��𢼴u������U��\������9
��2���������K��	������ѝ��� �������(����� 2���  �  �eN=��M=�L=L=�VK=��J=��I=�I=�>H=iwG=5�F=9�E=kE=�QD=3�C=��B=%�A=�A=�M@=}?=�>=��====-<=�U;=�|:=J�9=<�8=��7=	7=�'6=�D5=y_4=fx3=?�2=��1=w�0=��/=��.=�-=��,=c�+=#�*=,�)=h�(=��'=K�&=��%=/�$=p�#=��"=S�!=�w =�Y=�8=�=4�='�=l�=\=�$=��=�=�h="=��=r�=E7=6�==�=\)
=��=�a=f�=�=�=�=f, =8`�<c`�<yY�<�K�<�6�<�<���<.��<8��<'l�<1�<@��<���<�]�<��<h��<X[�<���<d��<�.�<U¼<�Q�<�ݵ<Gf�<x�<�m�<�<�i�<.�<I\�<nҙ<�F�<���<+�<V��<�
�<7y�<@�<�z<�s<�`l<y<e<v^<��V<�O<�H<��A<Ӈ:<os3<�b,<�V%<,O<�L<�O<�X	<Ah<���;!7�;���;
��;.D�;���;ZM�;��;R��;L�z;��`;�zF;�,;��;0��:;ܿ:���:2G7:җ�9�z]��>޹K�O�����v�ƺ����N�<�(���?��*V��fl�I2����xҖ��s��M����W������E�ʻ��Իp�޻xo���������P.����PQ�l���;������!��4&�Jm*�L�.�ϸ2��6���:���>�~�B�5�F�E�J��QN��R���U��Y�^3]���`��md�:�g�҆k��o�)�r���u��^y���|�<�������f��j��X����R����d����(��G����W��C쑼��:��ԟ���-��ź��KF���М��Y��*⟼si����u������b��X���+
��6����������U��������˝��!�������(�����2���  �  �eN=��M=	�L=	L=�VK=~�J=��I=�I=�>H=mwG=9�F=;�E=fE=�QD=0�C=��B= �A=�A=�M@=}?=�>=��====-<=�U;=�|:=K�9=;�8=w�7=�7=�'6=�D5=y_4=kx3=@�2=�1=|�0=��/=��.=�-=��,=Z�+=�*=-�)=j�(=��'=H�&=��%=0�$=w�#=��"=U�!=�w =�Y=�8=�=0�="�=g�=\=�$=��="�=�h="=��=t�=F7=6�=7�=R)
=��=�a=h�=	�=�=�=f, =D`�<b`�<}Y�<tK�<�6�<�<���</��<<��<'l�<1�<?��<���<�]�<��<n��<`[�<���<]��<�.�<P¼<�Q�<�ݵ<Of�<�<�m�<	�<�i�<,�<C\�<zҙ<�F�<���<�*�<I��<�
�<5y�<A�<�z<8�s<k`l<�<e<~^<��V<�O<n�H<��A<��:<os3<�b,<�V%<#O<�L<�O<�X	<gh<���;F7�;���;���;D�;���;@M�;��;t��;��z;�`;Q{F;�,;��;���:%ܿ:���:�G7:0��9֞]��A޹��O�v���w�ƺU���4���(�E�?��*V��fl�l2��N���Җ��s��C����W��i���]�ʻ��Իc�޻@o�h�С����c.���\Q�z���;�����!��4&� m*�(�.�Ǹ2��6���:���>�{�B�3�F�^�J�RN��R���U��Y�h3]���`��md�8�g���k��o�!�r���u�_y��|�C�������f��j��b����R����Q����(��?����W��M쑼��A��ٟ��	.��Ǻ��CF���М��Y��(⟼ti����u������\��W������8
��>����������R�������������!�������(�����!2���  �  �eN=��M=�L=L=�VK=�J=��I=�I=�>H=lwG=6�F=8�E=qE=�QD=1�C=��B=*�A=�A=�M@=}?=��>=��====-<=�U;=�|:=M�9=<�8={�7=	7=�'6=�D5=}_4=fx3==�2=��1=v�0=��/=��.=�-=�,=`�+=�*=*�)=l�(=��'=O�&=��%=0�$=x�#=��"=W�!=�w =�Y=�8=�=2�=&�=n�=�[=�$=��=�=�h="=��=o�=G7=5�=;�=X)
=��=�a=a�=�=�=�=d, =8`�<j`�<qY�<�K�<�6�<�<���<2��<=��<#l�<1�<5��<���<�]�<��<r��<T[�<���<`��<�.�<Q¼<�Q�<�ݵ<Ef�<��<�m�<�<�i�<+�<O\�<qҙ<�F�<���<+�<Q��<�
�<1y�<>�<�z<�s<�`l<u<e<w^<��V<
�O<��H<��A<��:<fs3<�b,<�V%<1O<�L<�O<�X	<(h<���;,7�;���;7��;D�;���;GM�;�;H��;��z;��`;zzF;��,;c�;K��:ܿ:I��:�G7:���9��]��>޹I�O� �����ƺ���j�W�(���?��*V��fl�U2������Җ��s��]����W������)�ʻ��Իe�޻8o���ȡ����N.����WQ�t���;�����!��4&�Km*�5�.���2�-�6���:���>�u�B�8�F�M�J�RN��R���U��Y�^3]���`��md�>�g�Іk��o�8�r���u��^y���|�=�������f��n��V����R����f����(��=����W��;쑼��?��؟���-��ɺ��NF���М��Y��⟼{i����u������X��]������0
��&��� ������S��������͝��!�������(�����2���  �  �eN=��M=�L=L=�VK=��J=��I=�I=�>H=vwG=4�F=7�E=nE=�QD=6�C=��B=+�A=�A=�M@=}?=�>=��====-<=�U;=�|:=M�9=:�8=}�7=�7=�'6=�D5=�_4=ex3=@�2=��1=s�0=��/=��.=�-=��,=[�+="�*=(�)=q�(=��'=O�&=��%=0�$={�#=��"=]�!=�w =�Y=�8=�=5�=!�=p�=�[=�$=��=!�=�h="=��=k�=M7=4�=<�=U)
=��=�a=d�=�=�=	�=h, =3`�<t`�<pY�<|K�<�6�<�<���<0��<A��<l�<1�<+��<ȩ�<�]�<��<s��<M[�<���<T��<�.�<J¼<�Q�<�ݵ<Af�<��<�m�< �<�i�<*�<K\�<jҙ<�F�<���<+�<B��<�
�<-y�<G�<��z<�s<�`l<y<e<^<��V<�O<~�H<��A<ԇ:<]s3<�b,<�V%<(O<�L<�O<Y	<3h<���;7�;���;&��;�C�;���; M�;�;,��;��z;�`;�zF;��,;�;���:�ۿ:R��:�G7:Ɩ�9�]�HC޹��O�L���k�ƺ���2���(�ְ?�:*V��fl�i2��7���Җ��s��n���wW������'�ʻ��Իg�޻!o軲򻒡����F.���UQ�h���;�����!�s4&�:m*�*�.���2�:�6���:���>�_�B�>�F�I�J�RN��R���U��Y�C3]���`��md�/�g�ۆk��o�;�r���u�_y���|�?�������f��x��Q����R����^����(��;����W��9쑼��5��ߟ���-��Ǻ��QF���М��Y��⟼}i����u������S��a��솪�@
��5���������N��������˝��!�������(�����)2���  �  �eN=��M=	�L=L=�VK=}�J=��I=�I=�>H=lwG=4�F=?�E=iE=�QD=6�C=��B=%�A=�A=�M@=}?=�>=��====-<=�U;=�|:=J�9=:�8={�7=	7=�'6=�D5=w_4=fx3=B�2=�1=z�0=��/=��.=�-=��,=_�+=!�*=(�)=k�(=��'=L�&=��%=.�$=u�#=��"=S�!=�w =�Y=�8=�=4�= �=n�=\=�$=��=�=�h=
"=��=r�=H7=4�=:�=X)
=��=�a=e�=�=�=�=g, =9`�<^`�<xY�<�K�<�6�<�<���<,��<@��<#l�<1�<2��<���<�]�<��<h��<e[�<���<V��<�.�<O¼<�Q�<�ݵ<Ff�<|�<�m�<�<�i�<&�<H\�<uҙ<�F�<���<	+�<K��<�
�<8y�<<�<�z<5�s<l`l<�<e<q^<��V<�O<��H<��A<ʇ:<`s3<�b,<�V%<'O<�L<�O<�X	<Oh<���;7�;��;���;D�;���;.M�;��;���;O�z;��`;�zF;&�,;M�;P��:ܿ:���:$G7:���9��]��?޹چO�������ƺ��� ���(�h�?��*V��fl�V2�����Җ��s��j����W������<�ʻ��Իu�޻Qo軥�������@.���RQ�k���;�����!��4&�<m*�:�.�˸2�2�6���:���>�s�B�?�F�N�J�RN��R���U��Y�m3]���`��md�5�g�Άk��o�+�r���u��^y���|�@�������f��n��V����R����]����(��F����W��C쑼��7��ٟ��.������MF���М��Y��#⟼wi����u������[��_��򆪼6
��-����������X�������������
!�������(�����2���  �  �eN=��M=�L=L=�VK=z�J=��I=�I=�>H=iwG=7�F=8�E=iE=�QD=+�C=��B=�A=�A=�M@=}?=�>=��====-<=�U;=�|:=L�9=?�8=x�7=	7=�'6=�D5=x_4=fx3=C�2=�1=~�0=��/=��.=��-=��,=_�+=�*=-�)=h�(=��'=K�&=��%=2�$=u�#=��"=R�!=�w =�Y=�8=�=/�=)�=f�=\=�$=��=�=�h="=��=u�=D7=8�=9�=V)
=��=�a=h�=�=�= �=h, =<`�<``�<|Y�<tK�<�6�<
�<���<1��<:��<,l�<1�<>��<���<�]�<��<f��<`[�<���<o��<�.�<Z¼<�Q�<�ݵ<Mf�<w�<�m�<�<�i�<#�<L\�<vҙ<�F�<���<�*�<Q��<�
�</y�<A�<֩z<A�s<k`l<�<e<d^<��V<�O<q�H<��A<��:<zs3<�b,<�V%<2O<�L<�O<�X	<\h<���;57�;���;���;HD�;b��;�M�;��;j��;[�z;��`;{F;#�,;��;���:�ܿ:C��:�G7:�9ؘ]��=޹ňO�������ƺ��� ���(��?��*V�vfl��2�� ���Җ��s��@����W��f���C�ʻ��ԻV�޻Oo軁������b.����VQ�{��~;�����!��4&�-m*�7�.�¸2�"�6���:���>���B�,�F�S�J�RN��R���U� �Y�r3]���`��md�1�g�Ȇk��o�#�r���u��^y���|�:�������f��e��_����R����Z����(��H����W��O쑼��H��ϟ�� .��̺��FF���М��Y��&⟼ki����u������_��R������1
��7���������`��󗳼�������!�������(�����2���  �  �eN=��M=�L=L=�VK=z�J=��I=�I=�>H=pwG=:�F=6�E=kE=�QD=+�C=��B=#�A=�A=�M@=}?=�>=��====-<=�U;=�|:=L�9=9�8=y�7= 	7=�'6=�D5=�_4=cx3=?�2=��1=r�0=��/=��.= �-=��,=^�+=�*=(�)=m�(=��'=O�&=��%=0�$=w�#=��"=X�!=�w =�Y=�8=�=0�=&�=g�=\=�$=��= �=�h=
"=��=q�=H7=3�=8�=U)
=��=�a=g�=�=�=�=g, =2`�<q`�<vY�<wK�<�6�<
�<���</��<:��<&l�<1�<2��<���<�]�<��<q��<Y[�<���<f��<�.�<U¼<�Q�<�ݵ<Of�<��<�m�<�<�i�<!�<Q\�<oҙ<�F�<���<+�<N��<�
�<,y�<L�<�z<�s<�`l<w<e<n^<��V<�O<{�H<��A<��:<_s3<�b,<�V%<:O<�L<�O<�X	<Jh<���;I7�;���;��;5D�;c��;gM�;��;T��;��z;�`;�zF;n�,;U�;���:Uܿ:��:�G7:��9��]�i@޹:�O�������ƺS���A�1�(��?��*V�]fl�{2��/���Җ��s��j����W������)�ʻ��Իf�޻>o軏򻻡�����c.���WQ�z���;�����!��4&�.m*�/�.���2�3�6���:���>�t�B�>�F�Y�J�RN��R���U��Y�U3]���`��md�4�g�݆k��o�/�r���u�_y���|�D�������f��k��Z����R����\����(��=����W��J쑼��G��ӟ���-��Ϻ��CF���М��Y��⟼vi����u������U��a������4
��5���������V��������̝��!�������(�����2���  �  �eN=��M=�L=L=�VK=~�J=��I=�I=�>H=mwG=2�F=>�E=mE=�QD=9�C=��B=)�A=�A=�M@=}?=�>=��====-<=�U;=�|:=M�9=6�8=��7=�7=�'6=�D5=|_4=fx3==�2=��1=r�0=��/=��.=�-=��,=_�+=%�*=$�)=o�(=��'=P�&=��%=1�$=w�#=��"=U�!=�w =�Y=�8=�=6�= �=r�= \=�$=��=�=�h=
"=��=k�=J7=1�==�=Y)
=��=�a=^�=�=�=�=e, =6`�<k`�<hY�<�K�<�6�<�<���<.��<?��<l�<1�<1��<©�<�]�<��<k��<^[�<���<W��<�.�<Q¼<�Q�<�ݵ<Bf�<��<�m�<�<�i�<(�<K\�<jҙ<�F�<���<+�<E��<�
�<3y�<4�<��z<�s<�`l<k<e<�^<��V<�O<��H<��A<߇:<Ks3<�b,<�V%<(O<�L<�O<�X	<2h<���;7�;؀�;��;D�;п�;*M�;�;w��;Z�z;��`;�zF;��,;E�;���:�ۿ:T��:
H7:���9�r]��B޹-�O�u���"�ƺ���g��(��?�@*V�gl�C2�����Җ��s�������W�������ʻ��Ի_�޻Ao���ѡ����9.���KQ�b���;�����!��4&�Fm*�8�.���2�2�6���:���>�i�B�I�F�B�J�RN��R���U�+�Y�I3]���`��md�:�g�Ԇk��o�I�r�n�u�_y���|�C�������f��v��O����R����d����(��C����W��9쑼��0��ן���-������QF���М��Y��⟼ui����u������O��j��熪�=
��'����������K��������ҝ��!�������(�����(2���  �  �eN=��M=�L=L=�VK=}�J=��I=�I=�>H=twG=5�F=;�E=lE=�QD=1�C=��B=&�A=�A=�M@=}?=�>=��====-<=�U;=�|:=O�9=8�8=}�7=�7=�'6=�D5=z_4=kx3=@�2=��1=x�0=��/=��.=�-=��,=[�+=!�*=)�)=m�(=��'=M�&=��%=1�$=w�#=��"=Y�!=�w =�Y=�8=�=2�=#�=l�=�[=�$=��= �=�h="=��=o�=I7=5�=;�=U)
=��=�a=b�=�=�=�=f, =@`�<g`�<qY�<}K�<�6�<�<���<1��<@��<"l�<1�<6��<���<�]�<��<p��<T[�<���<]��<�.�<J¼<�Q�<�ݵ<Ef�<��<�m�<�<�i�<'�<L\�<qҙ<�F�<���<+�<>��<�
�<5y�<;�<��z<%�s<�`l<}<e<�^<��V<�O<y�H<~�A<҇:<Zs3<�b,<�V%</O<�L<�O<�X	<Vh<���;#7�;���;��;D�;���;>M�;��;Q��;{�z;+�`;{F;H�,;s�;'��:#ܿ:���:[H7:���9�]�	D޹u�O�6���L�ƺR���:�a�(���?�X*V��fl�U2��H���Җ��s��_����W������6�ʻ��Ի\�޻Ao�r򻲡����O.�	��ZQ�s���;������!��4&�m*�0�.���2�+�6���:���>�n�B�:�F�K�J�RN��R���U��Y�R3]���`��md�7�g�k��o�9�r���u�_y���|�A�������f��n��Y����R����X����(��>����W��C쑼��>��ޟ���-��º��MF���М��Y�� ⟼qi����u������U��_���D
��9����������K��������ɝ��� �������(�����-2���  �  �eN=��M=�L=L=�VK={�J=��I=�I=�>H=iwG=9�F=8�E=nE=�QD=+�C=��B=&�A=�A=�M@=
}?=�>=��====-<=�U;=�|:=P�9=:�8=w�7=	7=�'6=�D5=z_4=ax3=?�2=��1=v�0=��/=��.=�-=��,=c�+=�*=.�)=g�(=��'=L�&=��%=.�$=q�#=��"=R�!=�w =�Y=�8=�=0�=)�=h�=\=�$=��=�=�h="=��=t�=C7=9�=8�=[)
=��=�a=h�=�=�=�=e, =1`�<``�<}Y�<{K�<�6�<�<���<6��<3��<,l�<1�<<��<���<�]�<��<m��<_[�<���<i��<�.�<S¼<�Q�<�ݵ<Of�<w�<�m�<
�<�i�<#�<Q\�<qҙ<�F�<���<�*�<Z��<�
�<5y�<E�<֩z<!�s<�`l<|<e<_^<��V<�O<��H<��A<��:<ns3<�b,<�V%<@O<�L<�O<�X	<Ah<���;E7�;���;&��;2D�;c��;oM�;��;k��;��z;h�`;�zF;�,;��;ܐ�:�ܿ:���:�H7:䖨9��]�=޹؇O�s���]�ƺ����E�u�(���?��*V�yfl�b2����sҖ��s��8����W��z���A�ʻ��Իt�޻ko軴������].����YQ�y��};�����!��4&�Fm*�G�.�͸2�+�6���:���>���B�*�F�Y�J��QN��R���U���Y�q3]���`��md�<�g�ކk��o�!�r���u��^y���|�?��|����f��e��]����R����c����(��A����W��G쑼	��G��֟���-��ɺ��DF���М��Y��'⟼pi����u������^��T�����'
��0����������`��������ɝ��!�������(�����2���  �  �eN=��M=�L=L=�VK=y�J=��I=�I=�>H=mwG=9�F=8�E=lE=�QD=3�C=��B=%�A=�A=�M@=}?=�>=��====-<=�U;=�|:=Q�9=;�8=u�7=�7=�'6=�D5=|_4=fx3=A�2=��1=z�0=��/=��.= �-=��,=Z�+=�*=.�)=l�(=��'=K�&=��%=2�$=|�#=��"=X�!=�w =�Y=�8=�=2�=#�=k�=\=�$=��=$�=�h="=��=r�=G7=9�=6�=Q)
=��=�a=d�=�=�=�=g, =;`�<h`�<tY�<wK�<�6�< �<���<8��<8��<"l�<
1�<:��<é�<�]�<��<s��<][�<���<]��<�.�<N¼<�Q�<�ݵ<Of�<��<�m�<�<�i�<!�<H\�<sҙ<�F�<���<�*�<H��<�
�<.y�<=�<�z<-�s<�`l<�<e<q^<��V<�O<p�H<��A<��:<os3<�b,<�V%<(O<�L<�O<�X	<Xh<���;G7�;���;��;D�;���;:M�;��;i��;��z;��`;>{F;��,;��;���:ܿ:��:�H7:��9ӣ]�B޹��O���ƺ����?�(�c�?��*V��fl�}2��J���Җ��s��8����W��}���I�ʻ��ԻR�޻o軈򻽡�����Z.�
��YQ�q���;������!��4&�/m*��.���2�+�6���:���>�v�B�)�F�_�J�#RN��R���U��Y�\3]���`��md�2�g�ʆk��o�2�r���u�_y��|�A��y����f��n��`����R����S����(��;����W��D쑼��9��ڟ���-��ɺ��DF���М��Y��⟼oi����u������V��T�����9
��:���������U���������ĝ��
!�������(�����!2���  �  �eN=��M=�L=L=�VK=��J=��I=�I=�>H=pwG=5�F=;�E=oE=�QD=;�C=��B=*�A=�A=�M@=}?=�>=��====-<=�U;=�|:=G�9=7�8=��7=	7=�'6=�D5=z_4=gx3==�2=�1=u�0=��/=��.=�-=��,=b�+=#�*='�)=i�(=��'=N�&=��%=.�$=s�#=��"=X�!=�w =�Y=�8=�=5�=#�=q�=�[=�$=��=�=�h="=��=p�=F7=1�=<�=[)
=��=�a=a�=�=�= �=c, =;`�<f`�<pY�<�K�<�6�<�<���<)��<>��<&l�<1�<6��<���<�]�<��<n��<R[�<���<Y��<�.�<K¼<�Q�<�ݵ<Ff�<��<�m�<
�<�i�<.�<K\�<sҙ<�F�<���<+�<M��<�
�<<y�<9�<��z< �s<w`l<{<e<�^<��V<�O<��H<��A<�:<Vs3<�b,<�V%</O<�L<�O<�X	<Ch<���;$7�;���;/��;�C�;޿�;*M�;�;P��;o�z;ƒ`;�zF;)�,;w�;]��:Kܿ:���:zF7:V��9�m]��?޹�O����c�ƺ����k���(���?��*V��fl�'2����Җ��s��u����W������+�ʻ��Իt�޻`o軻򻼡����?.���RQ�e���;�����!��4&�=m*�A�.�ɸ2�#�6���:���>�z�B�H�F�F�J��QN��R���U��Y�_3]���`��md�C�g�ˆk��o�;�r�s�u�_y���|�A�������f��k��R����R����d����(��@����W��:쑼��.��ݟ���-������MF���М��Y��&⟼ui����u������a��a��ꆪ�4
��-����������M��������ʝ��!�������(�����2���  �  �eN=��M=�L=L=�VK=y�J=��I=�I=�>H=mwG=9�F=8�E=lE=�QD=3�C=��B=%�A=�A=�M@=}?=�>=��====-<=�U;=�|:=Q�9=;�8=u�7=�7=�'6=�D5=|_4=fx3=A�2=��1=z�0=��/=��.= �-=��,=Z�+=�*=.�)=l�(=��'=K�&=��%=2�$=|�#=��"=X�!=�w =�Y=�8=�=2�=#�=k�=\=�$=��=$�=�h="=��=r�=G7=9�=6�=Q)
=��=�a=d�=�=�=�=g, =;`�<h`�<tY�<wK�<�6�< �<���<8��<8��<"l�<
1�<:��<é�<�]�<��<s��<][�<���<]��<�.�<N¼<�Q�<�ݵ<Of�<��<�m�<�<�i�<!�<H\�<sҙ<�F�<���<�*�<H��<�
�<.y�<=�<�z<-�s<�`l<�<e<q^<��V<�O<p�H<��A<��:<os3<�b,<�V%<(O<�L<�O<�X	<Xh<���;G7�;���;��;D�;���;:M�;��;i��;��z;��`;>{F;��,;��;���:ܿ:��:�H7:��9֣]�B޹��O���ƺ����?�(�c�?��*V��fl�}2��J���Җ��s��8����W��}���J�ʻ��ԻR�޻o軈򻽡�����Z.�
��YQ�q���;������!��4&�/m*��.���2�+�6���:���>�v�B�)�F�_�J�#RN��R���U��Y�\3]���`��md�2�g�ʆk��o�2�r���u�_y��|�A��y����f��n��`����R����S����(��;����W��D쑼��9��ڟ���-��ɺ��DF���М��Y��⟼oi����u������V��T�����9
��:���������U���������ĝ��
!�������(�����!2���  �  �eN=��M=�L=L=�VK={�J=��I=�I=�>H=iwG=9�F=8�E=nE=�QD=+�C=��B=&�A=�A=�M@=
}?=�>=��====-<=�U;=�|:=P�9=:�8=w�7=	7=�'6=�D5=z_4=ax3=?�2=��1=v�0=��/=��.=�-=��,=c�+=�*=.�)=g�(=��'=L�&=��%=.�$=q�#=��"=R�!=�w =�Y=�8=�=0�=)�=h�=\=�$=��=�=�h="=��=t�=C7=9�=8�=[)
=��=�a=h�=�=�=�=e, =1`�<``�<}Y�<{K�<�6�<�<���<6��<3��<,l�<1�<<��<���<�]�<��<m��<_[�<���<i��<�.�<S¼<�Q�<�ݵ<Of�<w�<�m�<
�<�i�<#�<Q\�<qҙ<�F�<���<�*�<Z��<�
�<5y�<E�<֩z<!�s<�`l<|<e<_^<��V<�O<��H<��A<��:<ns3<�b,<�V%<@O<�L<�O<�X	<Ah<���;E7�;���;&��;2D�;c��;oM�;��;k��;��z;h�`;�zF;�,;��;ܐ�:�ܿ:���:�H7:㖨9��]�=޹؇O�s���]�ƺ����E�u�(���?��*V�yfl�c2����sҖ��s��8����W��z���A�ʻ��Իt�޻ko軴������].����YQ�y��};�����!��4&�Fm*�G�.�͸2�+�6���:���>���B�*�F�Y�J��QN��R���U���Y�q3]���`��md�<�g�ކk��o�!�r���u��^y���|�?��|����f��e��]����R����c����(��A����W��G쑼	��G��֟���-��ɺ��DF���М��Y��'⟼pi����u������^��T�����'
��0����������`��������ɝ��!�������(�����2���  �  �eN=��M=�L=L=�VK=}�J=��I=�I=�>H=twG=5�F=;�E=lE=�QD=1�C=��B=&�A=�A=�M@=}?=�>=��====-<=�U;=�|:=O�9=8�8=}�7=�7=�'6=�D5=z_4=kx3=@�2=��1=x�0=��/=��.=�-=��,=[�+=!�*=)�)=m�(=��'=M�&=��%=1�$=w�#=��"=Y�!=�w =�Y=�8=�=2�=#�=l�=�[=�$=��= �=�h="=��=o�=I7=5�=;�=U)
=��=�a=b�=�=�=�=f, =@`�<g`�<qY�<}K�<�6�<�<���<1��<@��<"l�<1�<6��<���<�]�<��<p��<T[�<���<]��<�.�<J¼<�Q�<�ݵ<Ef�<��<�m�<�<�i�<'�<L\�<qҙ<�F�<���<+�<>��<�
�<5y�<;�<��z<%�s<�`l<}<e<�^<��V<�O<y�H<~�A<҇:<Zs3<�b,<�V%</O<�L<�O<�X	<Vh<���;#7�;���;��;D�;���;>M�;��;Q��;{�z;+�`;{F;H�,;s�;'��:"ܿ:���:ZH7:���9�]�D޹v�O�6���L�ƺS���;�a�(���?�X*V��fl�U2��H���Җ��s��_����W������6�ʻ��Ի\�޻Ao�r򻲡����O.�	��ZQ�s���;������!��4&�m*�0�.���2�+�6���:���>�n�B�:�F�K�J�RN��R���U��Y�R3]���`��md�7�g�k��o�9�r���u�_y���|�A�������f��n��Y����R����X����(��>����W��C쑼��>��ޟ���-��º��MF���М��Y�� ⟼qi����u������U��_���D
��9����������K��������ɝ��� �������(�����-2���  �  �eN=��M=�L=L=�VK=~�J=��I=�I=�>H=mwG=2�F=>�E=mE=�QD=9�C=��B=)�A=�A=�M@=}?=�>=��====-<=�U;=�|:=M�9=6�8=��7=�7=�'6=�D5=|_4=fx3==�2=��1=r�0=��/=��.=�-=��,=_�+=%�*=$�)=o�(=��'=P�&=��%=1�$=w�#=��"=U�!=�w =�Y=�8=�=6�= �=r�= \=�$=��=�=�h=
"=��=k�=J7=1�==�=Y)
=��=�a=^�=�=�=�=e, =6`�<k`�<hY�<�K�<�6�<�<���<.��<?��<l�<1�<1��<©�<�]�<��<k��<^[�<���<W��<�.�<Q¼<�Q�<�ݵ<Bf�<��<�m�<�<�i�<(�<K\�<jҙ<�F�<���<+�<E��<�
�<3y�<4�<��z<�s<�`l<k<e<�^<��V<�O<��H<��A<߇:<Ks3<�b,<�V%<(O<�L<�O<�X	<2h<���;7�;؀�;��;D�;п�;*M�;�;w��;Y�z;��`;�zF;��,;E�;���:�ۿ:T��:	H7:���9�r]��B޹.�O�v���"�ƺ���g��(��?�@*V�gl�C2�����Җ��s�������W�������ʻ��Ի_�޻Bo���ѡ����9.���KQ�b���;�����!��4&�Fm*�8�.���2�2�6���:���>�i�B�I�F�B�J�RN��R���U�+�Y�I3]���`��md�:�g�Ԇk��o�I�r�n�u�_y���|�C�������f��v��O����R����d����(��C����W��9쑼��0��ן���-������QF���М��Y��⟼ui����u������O��j��熪�=
��'����������K��������ҝ��!�������(�����(2���  �  �eN=��M=�L=L=�VK=z�J=��I=�I=�>H=pwG=:�F=6�E=kE=�QD=+�C=��B=#�A=�A=�M@=}?=�>=��====-<=�U;=�|:=L�9=9�8=y�7= 	7=�'6=�D5=�_4=cx3=?�2=��1=r�0=��/=��.= �-=��,=^�+=�*=(�)=m�(=��'=O�&=��%=0�$=w�#=��"=X�!=�w =�Y=�8=�=0�=&�=g�=\=�$=��= �=�h=
"=��=q�=H7=3�=8�=U)
=��=�a=g�=�=�=�=g, =2`�<q`�<vY�<wK�<�6�<
�<���</��<:��<&l�<1�<2��<���<�]�<��<q��<Y[�<���<f��<�.�<U¼<�Q�<�ݵ<Of�<��<�m�<�<�i�<!�<Q\�<oҙ<�F�<���<+�<N��<�
�<,y�<L�<�z<�s<�`l<w<e<n^<��V<�O<{�H<��A<��:<_s3<�b,<�V%<:O<�L<�O<�X	<Jh<���;I7�;���;��;4D�;c��;gM�;��;T��;��z;�`;�zF;n�,;T�;���:Uܿ:��:�G7:��9œ]�k@޹;�O�������ƺS���B�1�(��?��*V�]fl�{2��/���Җ��s��j����W������)�ʻ��Իf�޻>o軏򻻡�����c.���WQ�z���;�����!��4&�.m*�/�.���2�3�6���:���>�t�B�>�F�Y�J�RN��R���U��Y�U3]���`��md�4�g�݆k��o�/�r���u�_y���|�D�������f��k��Z����R����\����(��=����W��J쑼��G��ӟ���-��Ϻ��CF���М��Y��⟼vi����u������U��a������4
��5���������V��������̝��!�������(�����2���  �  �eN=��M=�L=L=�VK=z�J=��I=�I=�>H=iwG=7�F=8�E=iE=�QD=+�C=��B=�A=�A=�M@=}?=�>=��====-<=�U;=�|:=L�9=?�8=x�7=	7=�'6=�D5=x_4=fx3=C�2=�1=~�0=��/=��.=��-=��,=_�+=�*=-�)=h�(=��'=K�&=��%=2�$=u�#=��"=R�!=�w =�Y=�8=�=/�=)�=f�=\=�$=��=�=�h="=��=u�=D7=8�=9�=V)
=��=�a=h�=�=�= �=h, =<`�<``�<|Y�<tK�<�6�<
�<���<1��<:��<,l�<1�<>��<���<�]�<��<f��<`[�<���<o��<�.�<Z¼<�Q�<�ݵ<Mf�<w�<�m�<�<�i�<#�<L\�<vҙ<�F�<���<�*�<Q��<�
�</y�<A�<֩z<A�s<k`l<�<e<d^<��V<�O<q�H<��A<��:<zs3<�b,<�V%<2O<�L<�O<�X	<\h<���;57�;���;���;HD�;b��;�M�;��;j��;[�z;��`;{F;#�,;��;���:�ܿ:C��:�G7:9�]��=޹ƈO�������ƺ��� ���(��?��*V�vfl��2�� ���Җ��s��@����W��f���C�ʻ��ԻV�޻Oo軁������b.����VQ�{��~;�����!��4&�-m*�7�.�¸2�"�6���:���>���B�,�F�S�J�RN��R���U� �Y�r3]���`��md�1�g�Ȇk��o�#�r���u��^y���|�:�������f��e��_����R����Z����(��H����W��O쑼��H��ϟ�� .��̺��FF���М��Y��&⟼ki����u������_��R������1
��7���������`��󗳼�������!�������(�����2���  �  �eN=��M=	�L=L=�VK=}�J=��I=�I=�>H=lwG=4�F=?�E=iE=�QD=6�C=��B=%�A=�A=�M@=}?=�>=��====-<=�U;=�|:=J�9=:�8={�7=	7=�'6=�D5=w_4=fx3=B�2=�1=z�0=��/=��.=�-=��,=_�+=!�*=(�)=k�(=��'=L�&=��%=.�$=u�#=��"=S�!=�w =�Y=�8=�=4�= �=n�=\=�$=��=�=�h=
"=��=r�=H7=4�=:�=X)
=��=�a=e�=�=�=�=g, =9`�<^`�<xY�<�K�<�6�<�<���<,��<A��<#l�<1�<2��<���<�]�<��<h��<e[�<���<V��<�.�<O¼<�Q�<�ݵ<Ff�<|�<�m�<�<�i�<&�<H\�<uҙ<�F�<���<	+�<K��<�
�<8y�<<�<�z<5�s<l`l<�<e<q^<��V<�O<��H<��A<ʇ:<`s3<�b,<�V%<'O<�L<�O<�X	<Oh<���;7�;��;���;D�;���;.M�;��;���;O�z;��`;�zF;%�,;M�;P��:ܿ:���:#G7:���9Ɍ]��?޹ۆO�������ƺ��� ���(�h�?��*V��fl�V2�����Җ��s��j����W������<�ʻ��Իu�޻Qo軦�������@.���RQ�k���;�����!��4&�<m*�:�.�˸2�2�6���:���>�s�B�?�F�N�J�RN��R���U��Y�m3]���`��md�5�g�Άk��o�+�r���u��^y���|�@�������f��n��V����R����]����(��F����W��C쑼��7��ٟ��.������MF���М��Y��#⟼wi����u������[��_��򆪼6
��-����������X�������������
!�������(�����2���  �  �eN=��M=�L=L=�VK=��J=��I=�I=�>H=vwG=4�F=7�E=nE=�QD=6�C=��B=+�A=�A=�M@=}?=�>=��====-<=�U;=�|:=M�9=:�8=}�7=�7=�'6=�D5=�_4=ex3=@�2=��1=s�0=��/=��.=�-=��,=[�+="�*=(�)=q�(=��'=O�&=��%=0�$={�#=��"=]�!=�w =�Y=�8=�=5�=!�=p�=�[=�$=��=!�=�h="=��=k�=M7=4�=<�=U)
=��=�a=d�=�=�=	�=h, =3`�<t`�<pY�<|K�<�6�<�<���<0��<A��<l�<1�<+��<ȩ�<�]�<��<s��<M[�<���<T��<�.�<J¼<�Q�<�ݵ<Af�<��<�m�< �<�i�<*�<K\�<jҙ<�F�<���<+�<B��<�
�<-y�<G�<��z<�s<�`l<y<e<^<��V<�O<~�H<��A<ԇ:<]s3<�b,<�V%<(O<�L<�O<Y	<3h<���;7�;���;&��;�C�;���; M�;�;,��;��z;�`;�zF;��,;�;���:�ۿ:R��:�G7:Ė�9�]�IC޹��O�L���k�ƺ���3���(�ְ?�:*V��fl�i2��8���Җ��s��n���wW������'�ʻ��Իg�޻!o軲򻒡����F.���UQ�h���;�����!�s4&�:m*�*�.���2�:�6���:���>�_�B�>�F�I�J�RN��R���U��Y�C3]���`��md�/�g�ۆk��o�;�r���u�_y���|�?�������f��x��Q����R����^����(��;����W��9쑼��5��ߟ���-��Ǻ��QF���М��Y��⟼}i����u������S��a��솪�@
��5���������N��������˝��!�������(�����)2���  �  �eN=��M=�L=L=�VK=�J=��I=�I=�>H=lwG=6�F=8�E=qE=�QD=1�C=��B=*�A=�A=�M@=}?=��>=��====-<=�U;=�|:=M�9=<�8={�7=	7=�'6=�D5=}_4=fx3==�2=��1=v�0=��/=��.=�-=�,=`�+=�*=*�)=l�(=��'=O�&=��%=0�$=x�#=��"=W�!=�w =�Y=�8=�=2�=&�=n�=�[=�$=��=�=�h="=��=o�=G7=5�=;�=X)
=��=�a=a�=�=�=�=d, =8`�<j`�<qY�<�K�<�6�<�<���<2��<=��<#l�<1�<5��<���<�]�<��<r��<T[�<���<`��<�.�<Q¼<�Q�<�ݵ<Ef�<��<�m�<�<�i�<+�<O\�<qҙ<�F�<���<+�<Q��<�
�<1y�<>�<�z<�s<�`l<u<e<w^<��V<
�O<��H<��A<��:<fs3<�b,<�V%<1O<�L<�O<�X	<(h<���;,7�;���;7��;D�;���;GM�;�;H��;��z;��`;zzF;��,;c�;K��:ܿ:I��:�G7:���9��]��>޹J�O� �����ƺ���k�W�(���?��*V��fl�U2������Җ��s��]����W������)�ʻ��Իe�޻8o���ȡ����N.����WQ�t���;�����!��4&�Km*�5�.���2�-�6���:���>�u�B�8�F�M�J�RN��R���U��Y�^3]���`��md�>�g�Іk��o�8�r���u��^y���|�=�������f��n��V����R����f����(��=����W��;쑼��?��؟���-��ɺ��NF���М��Y��⟼{i����u������X��]������0
��&��� ������S��������͝��!�������(�����2���  �  �eN=��M=	�L=	L=�VK=~�J=��I=�I=�>H=mwG=9�F=;�E=fE=�QD=0�C=��B= �A=�A=�M@=}?=�>=��====-<=�U;=�|:=K�9=;�8=w�7=�7=�'6=�D5=y_4=kx3=@�2=�1=|�0=��/=��.=�-=��,=Z�+=�*=-�)=j�(=��'=H�&=��%=0�$=w�#=��"=U�!=�w =�Y=�8=�=0�="�=g�=\=�$=��="�=�h="=��=t�=F7=6�=7�=R)
=��=�a=h�=	�=�=�=f, =D`�<b`�<}Y�<tK�<�6�<�<���</��<<��<'l�<1�<?��<���<�]�<��<n��<`[�<���<]��<�.�<P¼<�Q�<�ݵ<Of�<�<�m�<�<�i�<,�<C\�<zҙ<�F�<���<�*�<I��<�
�<5y�<A�<�z<8�s<k`l<�<e<~^<��V<�O<n�H<��A<��:<os3<�b,<�V%<#O<�L<�O<�X	<gh<���;F7�;���;���;D�;���;@M�;��;t��;��z;�`;P{F;�,;��;���:$ܿ:���:�G7:/��9۞]��A޹��O�v���x�ƺU���5���(�E�?��*V��fl�l2��N���Җ��s��C����W��i���]�ʻ��Իc�޻@o�i�С����c.���\Q�z���;�����!��4&� m*�(�.�Ǹ2��6���:���>�{�B�3�F�^�J�RN��R���U��Y�h3]���`��md�8�g���k��o�!�r���u�_y��|�C�������f��j��b����R����Q����(��?����W��M쑼��A��ٟ��	.��Ǻ��CF���М��Y��(⟼ti����u������\��W������8
��>����������R�������������!�������(�����!2���  �  �eN=��M=�L=L=�VK=��J=��I=�I=�>H=iwG=5�F=9�E=kE=�QD=3�C=��B=%�A=�A=�M@=}?=�>=��====-<=�U;=�|:=J�9=<�8=��7=	7=�'6=�D5=y_4=fx3=?�2=��1=w�0=��/=��.=�-=��,=c�+=#�*=,�)=h�(=��'=K�&=��%=/�$=p�#=��"=S�!=�w =�Y=�8=�=4�='�=l�=\=�$=��=�=�h="=��=r�=E7=6�==�=\)
=��=�a=f�=�=�=�=f, =8`�<c`�<yY�<�K�<�6�<�<���<.��<8��<'l�<1�<@��<���<�]�<��<h��<X[�<���<d��<�.�<U¼<�Q�<�ݵ<Gf�<x�<�m�<�<�i�<.�<I\�<nҙ<�F�<���<+�<V��<�
�<7y�<@�<�z<�s<�`l<y<e<v^<��V<�O<�H<��A<Ӈ:<os3<�b,<�V%<,O<�L<�O<�X	<Ah<���;!7�;���;
��;/D�;���;ZM�;��;R��;L�z;��`;�zF;�,;��;0��:;ܿ:���:2G7:ї�9�z]��>޹K�O�����v�ƺ����N�<�(���?��*V��fl�I2����xҖ��s��M����W������E�ʻ��Իp�޻xo���������P.����PQ�l���;������!��4&�Jm*�L�.�ϸ2��6���:���>�~�B�5�F�E�J��QN��R���U��Y�^3]���`��md�:�g�҆k��o�)�r���u��^y���|�<�������f��j��X����R����d����(��G����W��C쑼��:��ԟ���-��ź��KF���М��Y��*⟼si����u������b��X���+
��6����������U��������˝��!�������(�����2���  �  �dN==�M=u�L=4L=�TK=C�J=w�I=I=	<H=YtG=�F=��E=�E=�MD=�C=�B=[�A=~A=�H@=xw?=)�>=��==��<=_&<=�N;=ku:=��9=B�8=,�7=] 7=�6=B;5=�U4=mn3=�2=K�1=i�0=T�/=��.=��-=z�,=��+=��*=��)=��(=��'=��&=��%=�$=�#=��"=�!=<g =	I=\'=C=��=>�=W}=�I=i=D�=j�=�U==��=dv=7$=%�=1t=[
=��=!O=��=�x=�=�=� =�<�<�=�<X7�<
*�<��<���<���<���<y��<;O�<	�<��<���<�D�<G��<��<�D�<.��<��<��<���<�@�<�͵<W�<cݮ<�`�<�<�^�<5ڠ<mS�<�ʙ<@�<鳒<b&�<���<�<�w�<��<k�z<��s<7fl<#De<a#^<�W<�O<��H<ȱA<�:<ʉ3<r{,<Aq%<�k<�k<�p<�{	<&�<�J�;M��;���;�3�;��;�!�;ղ�;sW�;f�;ظ{;�{a;6kG;Ї-;��;͙�:R��:9��: �;:!v�9�O�jչ^�J�'��Xkĺ�;�%����'�+q>��T��"k�����&o��</��Р��Q��7��������ʻi!Ի�޻����y����9�����{������j���T��!���%�**�=W.�Hx2�8�6�'�:���>�ۅB�$mF��IJ�N�;�Q���U��WY�-]�C�`�~@d���g��\k���n��Yr���u��:y���|�N ��2���4W��c���뢆��D��n䉼������������L���ᑼ6u�����񖖼�%��㲙��>���ɜ�cS���۟��c���ꢼ�p��~���d{������߃�����銭���*���#��N���g��ڝ��h!��m����)������$4���  �  �dN==�M=o�L=7L=~TK=E�J=y�I=I=	<H=RtG=�F=��E=�E=�MD=�C="�B=`�A=�A=�H@=rw?=&�>=��==��<=_&<=�N;=mu:=��9=B�8=4�7=e 7=�6=J;5=�U4=ln3=�2=I�1=l�0=L�/=��.=��-=��,=��+=��*=��)=��(=��'=��&=��%=߾$=ӭ#=��"=�!=>g =I=e'===��=F�=\}=�I=a=A�=_�=�U==��=fv=5$=&�=5t=f
=��="O=��=�x=�=�=� =�<�<�=�<e7�<
*�<��<��<���<���<}��<=O�<�<��<s��<~D�<=��<
��<�D�<8��<���<u�<�<�@�<�͵<
W�<Rݮ<�`�<��<�^�<<ڠ<iS�<�ʙ<@�<곒<j&�<Ɨ�<�<�w�<��<R�z<��s<$fl<-De<K#^<�W<,�O<��H<�A<�:<̉3<^{,<Mq%<�k<�k<�p<�{	<&�<�J�;��;���;/4�;��;N!�;���;�W�;��;g�{;{{a;kG;�-;C�;���:=��:{��:1�;:"v�9@2�aչ�J�
&���kĺ-<����'��p>���T��"k������n���.���Ϡ��Q��W�������ʻE!Ի޻���y�S���9����s{�����G���T��!��%�**�hW.�ex2�%�6�4�:���>��B�"mF��IJ��N��Q���U�zWY�K]�9�`��@d���g��\k���n��Yr���u�c:y���|�J ��4���1W��b�����D���䉼������������L���ᑼ+u����������%��ײ���>���ɜ�cS��ܟ��c���ꢼ�p��w���n{������փ��w��㊭���,���/��G���q��՝��r!��o����)������4���  �  �dN=?�M=p�L=9L=xTK=C�J=|�I=I=<H=TtG=�F=��E=�E=�MD=�C=&�B=X�A=�A=�H@=yw?=0�>=��==��<=[&<=�N;=nu:=��9=A�8=-�7=` 7=�6=L;5=�U4=on3=�2=H�1=s�0=H�/=��.=��-=}�,=��+=��*=��)=��(=��'=��&=��%=�$=ح#=��"=�!=@g =I=e'=A=��=G�=R}=�I=b=K�=f�=�U==��=gv=6$=)�=1t=]
=��=O=��=�x=�=�=� ==�<�=�<i7�<*�<��<���<���<���<~��<9O�<��<��<u��<�D�<M��<
��<�D�<$��<���<~�<���<�@�<�͵<W�<Uݮ<�`�<�<�^�<9ڠ<^S�<�ʙ<@�<ﳒ<_&�<���<�<�w�<��<K�z<��s<fl<EDe<K#^<�W<'�O<��H<ԱA<�:<Ӊ3<a{,<Vq%<�k<�k<�p<�{	<W�<�J�;*��;���; 4�;&��;w!�;��;XW�;��;g�{;�{a;�kG;2�-;�;?��:���:���:��;:�u�9�O��չ��J��%��Tlĺ�;����,�'��p>���T��"k�����o��)/��'Р��Q��R�������*ʻ<!Ի�޻���xy�P���9����v{��� ��C���T��!� �%��)*�LW.�\x2��6�H�:���>�߅B�mF��IJ� N�-�Q���U�tWY�X]�!�`��@d���g��\k��n��Yr���u�v:y���|�O ��1���0W��e��������D���䉼������������L���ᑼ'u�������%��ⲙ��>���ɜ�IS��ܟ��c���ꢼq��q���l{������ც����銭���,���3��;���s��ɝ��s!��r����)������4���  �  �dN=>�M=q�L=4L=TK=E�J=u�I=I=<H=RtG=�F=��E=�E=�MD=�C=!�B=^�A=�A=�H@=tw?=#�>=��==��<=a&<=�N;=ku:=��9=C�8=2�7=e 7=�6=C;5=�U4=nn3=�2=K�1=m�0=O�/=��.=��-=��,=��+=��*=��)=��(=��'=��&=��%=�$=խ#=��"=�!=Bg =I=c'=?=��=D�=X}=�I=a=@�=`�=�U==��=ev=6$=%�=7t=c
=��="O=��=�x=�=�=� = =�<�=�<Z7�<*�<��< ��<���<���<z��<>O�<�<
��<{��<zD�<@��<��<�D�<2��<��<{�<�<�@�<�͵<W�<Qݮ<�`�<
�<�^�<:ڠ<jS�<�ʙ<@�<곒<k&�<×�<(�<�w�<��<X�z<��s<7fl<-De<R#^<�W<	�O<��H<�A<�:<Љ3<f{,<Cq%<�k<�k<�p<�{	<�<�J�;F��;���;4�;��;f!�;鲥;�W�;��;��{;�{a;�jG;{�-;��;���:g��:G��:��;:�v�9�:�lչ��J��&��lĺ�;�	����'��p>�V�T��"k������n���.���Ϡ��Q��S��������ʻR!Ի޻����y�P���9����|{�����P���T��!��%�"**�fW.�^x2�/�6�'�:���>��B�%mF��IJ��N��Q���U��WY�>]�4�`��@d���g��\k���n��Yr���u�^:y���|�G ��5���3W��a���袆��D��z䉼������������L���ᑼ0u����������%��۲���>���ɜ�hS��ܟ��c���ꢼ�p��|���k{������Ճ��z��ڊ����)���,��H���g��՝��o!��l����)������4���  �  �dN=;�M=u�L=4L=TK=G�J=s�I=I=<H=[tG=ޫF=��E=�E=�MD=�C= �B=c�A=�A=�H@=}w?=$�>=��==��<=b&<=�N;=nu:=��9=@�8=0�7=\ 7=�6=E;5=�U4=kn3=�2=K�1=g�0=R�/=��.=��-=~�,=��+=��*=��)=��(=��'=��&=��%=�$=׭#=��"=�!=9g =I=c'===��=C�=[}=�I=g=I�=c�=�U==��=av=;$=#�=4t=[
=��=!O=��=�x=�=�=� =�<�<�=�<[7�<*�<��<���<���<���<���<2O�<�<��<���<|D�<S��<��<�D�<;��<��<��<�<�@�<�͵<W�<cݮ<�`�<�<�^�<=ڠ<mS�<�ʙ<@�<峒<k&�<���<"�<�w�<��<[�z<��s</fl<De<N#^<�W<�O<��H<��A<�:<ŉ3<t{,<Aq%<�k<�k<�p<�{	<#�<�J�;��;���;74�;���;|!�;㲥;�W�;s�;k�{;/|a;�jG;��-;��;.��:���:���:�;:{u�9�@�չ~�J��&��kĺ4<�*����'�Cq>�/�T��"k�����o��E/��Р��Q����������ʻT!Ի�޻��绥y����9����}{�����T���T�(�!���%��)*�[W.�Ox2�4�6�#�:���>�˅B�,mF��IJ�N�6�Q���U��WY�0]�I�`��@d���g��\k���n��Yr���u��:y���|�M ��3���,W��l���梆��D��r䉼������������L���ᑼ0u����������%��ݲ���>���ɜ�bS��ܟ��c���ꢼ�p��~���a{������Ճ�����������#���+��T���k��ߝ��q!��e����)������*4���  �  �dN=>�M=p�L=6L=|TK=E�J=}�I=I=<H=VtG=�F=��E=�E=�MD=�C="�B=W�A=�A=�H@=zw?='�>=��==��<=a&<=�N;=lu:=��9=C�8=0�7=c 7=�6=H;5=�U4=mn3=��2=G�1=s�0=I�/=��.=��-=��,=��+=��*=��)=��(=��'=��&=��%=�$=ѭ#=��"=�!=?g =	I=a'=A=��=C�=V}=�I=`=H�=^�=�U==��=bv=6$='�=4t=_
=��="O=��=�x=�=�=� ==�<�=�<^7�<*�<��<���<���<���<{��<3O�<�<��<v��<}D�<M��<��<�D�<&��<��<��<���<�@�<�͵<
W�<Xݮ<�`�<��<�^�<;ڠ<hS�<�ʙ<@�<볒<k&�<���<#�<�w�<��<M�z<��s<fl<MDe<J#^<�W< �O<��H<ڱA<�:<щ3<`{,<Kq%<�k<�k<�p<�{	<5�<�J�;��;���;�3�;��;�!�;�;SW�;��;L�{;�{a;kG;#�-;g�;��:���:a��:B�;:�v�9/@��չ��J�^&��7lĺ�;����9�'��p>���T��"k������n�� /��Р��Q��P��������ʻA!Ի�޻�统y�N���9�����{������R���T�	�!��%�**�mW.�Yx2�#�6�-�:���>���B�mF��IJ��N��Q���U��WY�X]�"�`��@d���g��\k��n��Yr���u�g:y���|�J ��4���2W��k���袆��D���䉼������������L���ᑼ.u�����򖖼�%��ڲ���>���ɜ�XS��ܟ��c���ꢼ�p��y���n{������Ճ�����ߊ����.���1��8���y��ŝ��s!��t����)������4���  �  �dN=C�M=m�L=7L=�TK=?�J=~�I=I=<H=PtG=�F=��E=�E=�MD=��C=*�B=X�A=�A=�H@=uw?=+�>=��==��<=Y&<=�N;=mu:=��9=F�8=,�7=e 7=�6=L;5=�U4=nn3=�2=A�1=v�0=H�/=��.=��-=��,=��+=��*=��)=~�(=��'=��&=��%=�$=ԭ#=��"=�!=Eg =I=h'=>=��=K�=T}=�I=\=I�=a�=�U==��=gv=4$=*�=3t=a
=��=O=��=�x=�=�=� ==�<�=�<j7�<�)�<��<���<���<���<z��<@O�<��<��<w��<�D�<I��<��<�D�<&��<��<l�<���<�@�<�͵<W�<Jݮ<�`�<��<�^�<1ڠ<lS�<�ʙ<@�<�<`&�<ȗ�<�<�w�<��<B�z<��s<�el<LDe<@#^<�W<�O<��H<�A<�:<�3<T{,<Pq%<�k<sk<�p<�{	<G�<�J�;>��;���;4�;7��;)!�;1��;ZW�;��;K�{;�{a;ZkG;,�-;u�;��:���:i��:�;:Tx�9�P�չ@�J��%���kĺ�;������'�Vp>���T�t"k�ҏ���n��/��Р��Q��f�������ʻM!Ի�޻�绐y�z��}9����i{�����3���T��!��%��)*�`W.�Ux2�"�6�:�:���>��B�mF��IJ��N��Q���U�fWY�U]��`��@d���g��\k���n��Yr���u�c:y���|�F ��4���4W��^��������D��~䉼�������µ���L���ᑼu�������%��ڲ���>���ɜ�QS��ܟ��c���ꢼ�p��t���t{����������v��ꊭ������7��7������Ɲ��x!��e����)������4���  �  �dN=B�M=s�L=2L=TK=B�J=z�I=I=<H=UtG=�F=��E=�E=�MD=�C=)�B=[�A=�A=�H@=zw?=&�>=��==��<=\&<=�N;=ku:=��9=D�8=,�7=b 7=�6=E;5=�U4=jn3=�2=L�1=m�0=I�/=��.=��-=��,=��+=��*=��)=��(=��'=��&=��%=�$=ԭ#=��"=�!=?g =I=f'=@=��=I�=S}=�I=c=I�=a�=�U==��=bv=8$=)�=2t=\
=��=O=��=�x=�=�=� =�<�<�=�<]7�<
*�<��<���<���<���<z��<7O�<�<��<��<~D�<O��<��<�D�<)��< ��<y�<���<�@�<�͵<W�<Uݮ<�`�<�<�^�<5ڠ<lS�<�ʙ<@�<�<`&�<���<"�<�w�<��<?�z<��s<0fl<4De<<#^<�W<�O<��H<ٱA<�:<މ3<l{,<;q%<�k<k<�p<�{	<7�<�J�;6��;���;4�;;��;Z!�;'��;rW�;��;z�{; |a;kG;��-;;�;m��:2��:9��:�;:Nw�9sQ��չ��J��&���kĺn<�����'��p>���T��"k������n��-/��Р��Q��3��������ʻU!Ի�޻��绕y�>���9����p{�����>���T��!���%��)*�bW.�Rx2�-�6�2�:���>�ׅB�mF��IJ�N��Q���U�}WY�P]�7�`�|@d���g��\k���n��Yr���u�l:y���|�J ��/���3W��g���𢆼�D��w䉼������������L���ᑼ!u�����떖��%��岙��>���ɜ�XS��ܟ��c���ꢼ�p������e{������ც����������#���9��F���j��ҝ��z!��f����)������4���  �  �dN=8�M=v�L=5L=}TK=G�J=w�I=I=<H=VtG=�F=��E=�E=�MD=�C=�B=_�A=�A=�H@=yw?= �>=��==��<=c&<=�N;=nu:=��9=>�8=5�7=^ 7=�6=A;5=�U4=on3=�2=J�1=l�0=S�/=��.=��-=��,=��+=��*=��)=��(=��'=��&=��%=�$=ӭ#=��"=�!=>g =I=a'=?=��=@�=]}=�I=b=B�=^�=�U==��=`v=:$=$�=6t=`
=��=%O=��=�x=�=�=� = =�<�=�<Q7�<*�<��< ��<���<���<��<4O�<�<��<~��<tD�<G��<��<�D�<7��<��<��<쯼<�@�<�͵<
W�<Yݮ<�`�<�<�^�<<ڠ<lS�<�ʙ<@�<೒<s&�<���<+�<�w�<��<k�z<��s<%fl<(De<a#^<�W<�O<��H<ȱA</�:<��3<w{,<Eq%<�k<�k<�p<�{	<�<�J�;��;���;4�;ܡ�;�!�;���;�W�;��;P�{;�{a;�jG;}�-;�;K��:���:���:�;:Yt�9�/��չ4�J�E'���kĺ�;�$���'��p>��T�Q#k������n��#/���Ϡ��Q��(��������ʻX!Ի�޻	���y�@���9�����{������_���T��!���%�**�nW.�Sx2�7�6��:���>�υB�)mF��IJ��N��Q�z�U��WY�5]�9�`��@d���g��\k���n��Yr�x�u�s:y���|�N ��2���.W��k���⢆��D��w䉼Ł����������L���ᑼ;u����������%��Ӳ���>���ɜ�fS��ܟ��c���ꢼ�p�����b{������΃�����׊����1���#��J���p��؝��g!��r����)������%4���  �  �dN=9�M=t�L=6L=}TK=C�J=y�I=I=<H=XtG=ޫF=��E=�E=�MD=�C=!�B=^�A=�A=�H@=}w?=*�>=��==��<=^&<=�N;=lu:=��9=?�8=4�7=Z 7=�6=J;5=�U4=mn3=�2=G�1=m�0=N�/=��.=��-=z�,=��+=��*=��)=��(=��'=��&=��%=�$=ح#=��"=�!=>g =	I=d'=?=��=E�=X}=�I=c=K�=d�=�U==��=ev=9$=&�=2t=]
=��= O=��=�x=�=�=� =�<�<�=�<c7�<*�<��<���<~��<���<|��<8O�<�<��<���<�D�<R��<��<�D�<3��<��<��<�<�@�<�͵<W�<^ݮ<�`�<�<�^�<8ڠ<iS�<�ʙ<@�<䳒<n&�<���<�<�w�<��<X�z<��s<fl<.De<O#^<�W<&�O<��H<��A<(�:<��3<n{,<Hq%<�k<�k<�p<�{	<@�<�J�;	��;���; 4�; ��;�!�;첥;�W�;��;?�{;)|a;EkG;��-;3�;���:��:b��:�;:�t�9"3��չ;�J�&���kĺ<���/�'��p>�h�T��"k�����%o��0/��Р��Q��0��������ʻW!Ի�޻��练y�9���9����y{��� ��L���T��!���%��)*�TW.�Jx2�2�6�2�:���>�ӅB�"mF��IJ��N�=�Q���U�~WY�B]�6�`��@d���g��\k���n��Yr���u��:y���|�Q ��2���1W��f�����D��t䉼������������L���ᑼ.u����������%��ಙ��>���ɜ�TS��ܟ��c���ꢼ�p��x���e{������Ӄ�����銭���*���-��H���t��՝��q!��m����)������(4���  �  �dN=A�M=p�L=0L=�TK=B�J=y�I=I=<H=PtG=�F=��E=�E=�MD=�C=(�B=Z�A=�A=�H@=uw?=%�>=��==��<=]&<=�N;=eu:=��9=C�8=2�7=i 7=�6=H;5=�U4=ln3=�2=I�1=q�0=G�/=��.=��-=��,=��+=��*=��)=|�(=��'=��&=��%=�$=ҭ#=��"=�!=Dg =I=g'=@=��=I�=R}=�I=_=D�=^�=�U==��=fv=1$=*�=1t=e
=��=!O=��=�x=�=�=� = =�<�=�<`7�<	*�<��<���<���<���<o��<CO�<�<��<t��<}D�<D��<
��<�D�<'��<���<{�<���<�@�<͵<W�<Mݮ<�`�<��<�^�<7ڠ<oS�<�ʙ<	@�<�<b&�<З�<�<�w�<��<A�z<��s<%fl<BDe<A#^<�W<�O<��H<��A<�:<ۉ3<`{,<1q%<�k<�k<�p<�{	<1�<�J�;H��;���;4�;*��;j!�;!��;iW�;��;��{;�{a;�jG;�-;W�;���:���:���:ޡ;:�v�9�:�չ�J�f&��*lĺ0<�����'��p>���T��"k������n���.��!Р��Q��v��������ʻE!Ի�޻�绸y�k���9����k{�����;���T���!��%�**�lW.�_x2�$�6�/�:���>���B�mF��IJ��N��Q���U�{WY�]]�'�`��@d���g��\k��n��Yr���u�U:y���|�M ��/���>W��\���𢆼�D���䉼������������L���ᑼ"u�������%��岙��>���ɜ�\S��ܟ��c���ꢼ�p������p{������ރ��m��㊭���)���7��>���p��˝��x!��o����)������4���  �  �dN=>�M=s�L=5L=�TK=A�J=x�I=I=<H=TtG=�F=��E=�E=�MD=�C=!�B=\�A=�A=�H@=xw?=,�>=��==��<=]&<=�N;=ku:=��9=@�8=,�7=] 7=�6=E;5=�U4=on3=�2=E�1=o�0=Q�/=��.=��-=z�,=��+=��*=��)=��(=��'=��&=��%=�$=ۭ#=��"=�!=Bg =	I=b'=@=��=C�=V}=�I=b=I�=g�=�U==��=fv=6$=(�=0t=]
=��=!O=��=�x=�=�=� ==�<�=�<[7�<*�<��<���<}��<���<y��<>O�<�<
��<~��<�D�<K��<��<�D�<.��<��<~�<�<�@�<�͵<W�<Tݮ<�`�<�<�^�<4ڠ<mS�<�ʙ<@�<쳒<^&�<���<�<�w�<��<b�z<��s<fl<1De<[#^<�W<�O<��H<ͱA<�:<Ή3<m{,<Dq%<�k<{k<�p<�{	<D�<�J�;L��;���;4�;��;u!�;;}W�;��;��{;�{a;`kG;r�-;,�;���:y��:O��:9�;:�u�9�O�Uչ2�J��&��Pkĺ�;���Z�'��p>�6�T��"k�����*o��$/��*Р��Q��L��������ʻU!Ի�޻��绑y�H���9����{������R���T��!���%��)*�HW.�Ox2�/�6�2�:���>��B�mF��IJ��N�<�Q���U��WY�6]�-�`��@d���g��\k���n��Yr���u��:y���|�R ��/���4W��`���񢆼�D��w䉼������������L���ᑼ/u����������%��޲���>���ɜ�RS��ܟ��c���ꢼ�p��{���h{������⃪�������'���'��E���{��ӝ��k!��j����)������"4���  �  �dN=<�M=q�L=6L=}TK=F�J=x�I=I=	<H=RtG=߫F=��E=�E=�MD=�C=�B=c�A=�A=�H@=tw?=#�>=��==��<=b&<=�N;=nu:=��9=B�8=:�7=] 7=�6=G;5=�U4=gn3=�2=N�1=h�0=M�/=��.=��-=~�,=��+=��*=��)=��(=��'=��&=��%=�$=ѭ#=��"=�!=<g =I=a'=?=��=A�=^}=�I=b=A�=\�=�U==��=dv=9$=$�=8t=g
=��=(O=��=�x=�=�=� =�<�<�=�<Z7�<*�<��<��<���<���<~��<8O�<�<��<w��<xD�<@��<��<�D�<=��<��<��<ﯼ<�@�<�͵<W�<Pݮ<�`�<��<�^�<<ڠ<hS�<�ʙ<@�<䳒<v&�<���<!�<�w�<��<L�z<��s<2fl<,De<A#^<�W<.�O<��H<ϱA<;�:<Ɖ3<f{,<Jq%<�k<�k<�p<�{	<%�<�J�;��;���;64�;��;�!�;ϲ�;�W�;��;\�{;�{a;�jG;6�-;)�;��:��:���:3�;:zv�9X�Sչ�J�m&��lĺ�<����ƻ'�-q>��T�H#k�{���	o���.���Ϡ��Q��9��������ʻT!Ի�޻���y�C���9�����{������[���T��!���%�**�sW.�ax2�1�6�.�:���>�ԅB�*mF��IJ��N�.�Q�p�U��WY�G]�N�`�r@d���g��\k���n��Yr�v�u�}:y���|�J ��8���/W��f���袆��D��~䉼������������L���ᑼ7u����������%��ٲ���>���ɜ�cS��ܟ��c���ꢼ�p��y���i{������ʃ��~��ክ���4���3��L���j��֝��w!��u����)������!4���  �  �dN=>�M=s�L=5L=�TK=A�J=x�I=I=<H=TtG=�F=��E=�E=�MD=�C=!�B=\�A=�A=�H@=xw?=,�>=��==��<=]&<=�N;=ku:=��9=@�8=,�7=] 7=�6=E;5=�U4=on3=�2=E�1=o�0=Q�/=��.=��-=z�,=��+=��*=��)=��(=��'=��&=��%=�$=ۭ#=��"=�!=Bg =	I=b'=@=��=C�=V}=�I=b=I�=g�=�U==��=fv=6$=(�=0t=]
=��=!O=��=�x=�=�=� ==�<�=�<[7�<*�<��<���<}��<���<y��<>O�<�<
��<~��<�D�<K��<��<�D�<.��<��<~�<�<�@�<�͵<W�<Tݮ<�`�<�<�^�<4ڠ<mS�<�ʙ<@�<쳒<^&�<���<�<�w�<��<b�z<��s<fl<1De<[#^<�W<�O<��H<ͱA<�:<Ή3<m{,<Dq%<�k<{k<�p<�{	<D�<�J�;L��;���;4�;��;u!�;;}W�;��;��{;�{a;`kG;r�-;,�;���:y��:O��:9�;:�u�9�O�Uչ3�J��&��Pkĺ�;���Z�'��p>�6�T��"k�����*o��$/��*Р��Q��L��������ʻU!Ի�޻��绑y�H���9����{������R���T��!���%��)*�HW.�Ox2�/�6�2�:���>��B�mF��IJ��N�<�Q���U��WY�6]�-�`��@d���g��\k���n��Yr���u��:y���|�R ��/���4W��`���񢆼�D��w䉼������������L���ᑼ/u����������%��޲���>���ɜ�RS��ܟ��c���ꢼ�p��{���h{������⃪�������'���'��E���{��ӝ��k!��j����)������"4���  �  �dN=A�M=p�L=0L=�TK=B�J=y�I=I=<H=PtG=�F=��E=�E=�MD=�C=(�B=Z�A=�A=�H@=uw?=%�>=��==��<=]&<=�N;=eu:=��9=C�8=2�7=i 7=�6=H;5=�U4=ln3=�2=I�1=q�0=G�/=��.=��-=��,=��+=��*=��)=|�(=��'=��&=��%=�$=ҭ#=��"=�!=Dg =I=g'=@=��=I�=R}=�I=_=D�=^�=�U==��=fv=1$=*�=1t=e
=��=!O=��=�x=�=�=� = =�<�=�<`7�<	*�<��<���<���<���<o��<CO�<�<��<t��<}D�<D��<
��<�D�<'��<���<{�<���<�@�<͵<W�<Mݮ<�`�<��<�^�<7ڠ<oS�<�ʙ<	@�<�<b&�<З�<�<�w�<��<A�z<��s<%fl<BDe<A#^<�W<�O<��H<��A<�:<ۉ3<a{,<1q%<�k<�k<�p<�{	<1�<�J�;H��;���;4�;*��;j!�;!��;iW�;��;��{;�{a;�jG;�-;W�;���:���:���:ޡ;:�v�9;�չ�J�f&��*lĺ1<�����'��p>���T��"k������n���.��!Р��Q��v��������ʻE!Ի�޻�绸y�k���9����k{�����;���T���!��%�**�lW.�_x2�$�6�/�:���>���B�mF��IJ��N��Q���U�{WY�]]�'�`��@d���g��\k��n��Yr���u�U:y���|�M ��/���>W��\���𢆼�D���䉼������������L���ᑼ"u�������%��岙��>���ɜ�\S��ܟ��c���ꢼ�p������p{������ރ��m��㊭���)���7��>���p��˝��x!��o����)������4���  �  �dN=9�M=t�L=6L=}TK=C�J=y�I=I=<H=XtG=ޫF=��E=�E=�MD=�C=!�B=^�A=�A=�H@=}w?=*�>=��==��<=^&<=�N;=lu:=��9=?�8=4�7=Z 7=�6=J;5=�U4=mn3=�2=G�1=m�0=N�/=��.=��-=z�,=��+=��*=��)=��(=��'=��&=��%=�$=ح#=��"=�!=>g =	I=d'=?=��=E�=X}=�I=c=K�=d�=�U==��=ev=9$=&�=2t=]
=��= O=��=�x=�=�=� =�<�<�=�<d7�<*�<��<���<~��<���<|��<8O�<�<��<���<�D�<R��<��<�D�<3��<��<��<�<�@�<�͵<W�<^ݮ<�`�<�<�^�<8ڠ<iS�<�ʙ<@�<䳒<n&�<���<�<�w�<��<X�z<��s<fl<.De<O#^<�W<&�O<��H<��A<(�:<��3<n{,<Hq%<�k<�k<�p<�{	<@�<�J�;	��;���; 4�; ��;�!�;첥;�W�;��;?�{;)|a;EkG;��-;3�;���:��:b��:�;:�t�9,3��չ<�J�&���kĺ<���/�'��p>�h�T��"k�����%o��0/��Р��Q��0��������ʻW!Ի�޻��练y�9���9����y{��� ��L���T��!���%��)*�TW.�Jx2�2�6�2�:���>�ӅB�"mF��IJ��N�=�Q���U�~WY�B]�6�`��@d���g��\k���n��Yr���u��:y���|�Q ��2���1W��f�����D��t䉼������������L���ᑼ.u����������%��ಙ��>���ɜ�TS��ܟ��c���ꢼ�p��x���e{������Ӄ�����銭���*���-��H���t��՝��q!��m����)������(4���  �  �dN=8�M=v�L=5L=}TK=G�J=w�I=I=<H=VtG=�F=��E=�E=�MD=�C=�B=_�A=�A=�H@=yw?= �>=��==��<=c&<=�N;=nu:=��9=>�8=5�7=^ 7=�6=A;5=�U4=on3=�2=J�1=l�0=S�/=��.=��-=��,=��+=��*=��)=��(=��'=��&=��%=�$=ӭ#=��"=�!=>g =I=a'=?=��=@�=]}=�I=b=B�=^�=�U==��=`v=:$=$�=6t=`
=��=%O=��=�x=�=�=� = =�<�=�<Q7�<*�<��< ��<���<���<��<4O�<�<��<��<tD�<G��<��<�D�<7��<��<��<쯼<�@�<�͵<
W�<Yݮ<�`�<�<�^�<<ڠ<lS�<�ʙ<@�<೒<s&�<���<+�<�w�<��<k�z<��s<%fl<(De<a#^<�W<�O<��H<ȱA</�:<��3<w{,<Eq%<�k<�k<�p<�{	<�<�J�;��;���;4�;ܡ�;�!�;���;�W�;��;P�{;�{a;�jG;}�-;�;J��:���:���:�;:Wt�9�/��չ5�J�E'���kĺ�;�$���'��p>��T�Q#k������n��#/���Ϡ��Q��(��������ʻX!Ի�޻	���y�@���9�����{������_���T��!���%�**�nW.�Sx2�8�6��:���>�υB�*mF��IJ��N��Q�z�U��WY�5]�9�`��@d���g��\k���n��Yr�x�u�s:y���|�N ��2���.W��k���⢆��D��w䉼Ł����������L���ᑼ;u����������%��Ӳ���>���ɜ�fS��ܟ��c���ꢼ�p�����b{������΃�����׊����1���#��J���p��؝��g!��r����)������%4���  �  �dN=B�M=s�L=2L=TK=B�J=z�I=I=<H=UtG=�F=��E=�E=�MD=�C=)�B=[�A=�A=�H@=zw?=&�>=��==��<=\&<=�N;=ku:=��9=D�8=,�7=b 7=�6=E;5=�U4=jn3=�2=L�1=m�0=I�/=��.=��-=��,=��+=��*=��)=��(=��'=��&=��%=�$=ԭ#=��"=�!=?g =I=f'=@=��=I�=S}=�I=c=I�=a�=�U==��=bv=8$=)�=2t=\
=��=O=��=�x=�=�=� =�<�<�=�<]7�<
*�<��<���<���<���<z��<7O�<�<��<��<~D�<O��<��<�D�<)��< ��<y�<���<�@�<�͵<W�<Uݮ<�`�<�<�^�<5ڠ<lS�<�ʙ<@�<�<`&�<���<"�<�w�<��<?�z<��s<0fl<4De<<#^<�W<�O<��H<ٱA<�:<މ3<l{,<;q%<�k<k<�p<�{	<7�<�J�;6��;���;4�;;��;Z!�;'��;qW�;��;y�{; |a;kG;��-;:�;l��:1��:9��:�;:Mw�9Q��չ��J��&���kĺn<�����'��p>���T��"k������n��-/��Р��Q��3��������ʻU!Ի�޻��绕y�>���9����p{�����>���T��!���%��)*�bW.�Rx2�-�6�2�:���>�ׅB�mF��IJ�N��Q���U�}WY�P]�7�`�|@d���g��\k���n��Yr���u�l:y���|�J ��/���3W��g���𢆼�D��w䉼������������L���ᑼ!u�����떖��%��岙��>���ɜ�XS��ܟ��c���ꢼ�p������e{������ც����������#���9��F���j��ҝ��z!��f����)������4���  �  �dN=C�M=m�L=7L=�TK=?�J=~�I=I=<H=PtG=�F=��E=�E=�MD=��C=*�B=X�A=�A=�H@=uw?=+�>=��==��<=Y&<=�N;=mu:=��9=F�8=,�7=e 7=�6=L;5=�U4=nn3=�2=A�1=v�0=H�/=��.=��-=��,=��+=��*=��)=~�(=��'=��&=��%=�$=ԭ#=��"=�!=Eg =I=h'=>=��=K�=T}=�I=\=I�=a�=�U==��=gv=4$=*�=3t=a
=��=O=��=�x=�=�=� ==�<�=�<j7�<�)�<��<���<���<���<z��<@O�<��<��<w��<�D�<I��<��<�D�<&��<��<l�<���<�@�<�͵<W�<Jݮ<�`�<��<�^�<1ڠ<lS�<�ʙ<@�<�<`&�<ȗ�<�<�w�<��<B�z<��s<�el<LDe<@#^<�W<�O<��H<�A<�:<�3<T{,<Pq%<�k<sk<�p<�{	<G�<�J�;>��;���;4�;7��;)!�;1��;ZW�;��;K�{;�{a;YkG;,�-;u�;��:���:i��:�;:Sx�9�P�չ@�J��%���kĺ�;������'�Vp>���T�t"k�ҏ���n��/��Р��Q��f�������ʻM!Ի�޻�绐y�z��}9����i{�����3���T��!��%��)*�`W.�Ux2�"�6�:�:���>��B�mF��IJ��N��Q���U�fWY�U]��`��@d���g��\k���n��Yr���u�c:y���|�F ��4���4W��^��������D��~䉼�������µ���L���ᑼu�������%��ڲ���>���ɜ�QS��ܟ��c���ꢼ�p��t���t{����������v��ꊭ������7��7������Ɲ��x!��e����)������4���  �  �dN=>�M=p�L=6L=|TK=E�J=}�I=I=<H=VtG=�F=��E=�E=�MD=�C="�B=W�A=�A=�H@=zw?='�>=��==��<=a&<=�N;=lu:=��9=C�8=0�7=c 7=�6=H;5=�U4=mn3=��2=G�1=s�0=I�/=��.=��-=��,=��+=��*=��)=��(=��'=��&=��%=�$=ѭ#=��"=�!=?g =	I=a'=B=��=C�=V}=�I=`=H�=^�=�U==��=bv=6$='�=4t=_
=��="O=��=�x=�=�=� ==�<�=�<^7�<*�<��<���<���<���<{��<3O�<�<��<v��<}D�<M��<��<�D�<&��<��<��<���<�@�<�͵<
W�<Xݮ<�`�<��<�^�<;ڠ<hS�<�ʙ<@�<볒<k&�<���<#�<�w�<��<M�z<��s<fl<MDe<J#^<�W< �O<��H<ڱA<�:<щ3<`{,<Kq%<�k<�k<�p<�{	<5�<�J�;��;���;�3�;��;�!�;�;SW�;��;L�{;�{a;kG;#�-;g�;��:���:a��:B�;:�v�9:@��չ��J�_&��7lĺ�;����9�'��p>���T��"k������n�� /��Р��Q��P��������ʻA!Ի�޻�统y�N���9�����{������R���T�	�!��%�**�mW.�Yx2�#�6�-�:���>���B�mF��IJ��N��Q���U��WY�X]�"�`��@d���g��\k��n��Yr���u�g:y���|�J ��4���2W��k���袆��D���䉼������������L���ᑼ.u�����򖖼�%��ڲ���>���ɜ�XS��ܟ��c���ꢼ�p��y���n{������Ճ�����ߊ����.���1��8���y��ŝ��s!��t����)������4���  �  �dN=;�M=u�L=4L=TK=G�J=s�I=I=<H=[tG=ޫF=��E=�E=�MD=�C= �B=c�A=�A=�H@=}w?=$�>=��==��<=b&<=�N;=nu:=��9=@�8=0�7=\ 7=�6=E;5=�U4=kn3=�2=K�1=g�0=R�/=��.=��-=~�,=��+=��*=��)=��(=��'=��&=��%=�$=׭#=��"=�!=9g =I=c'===��=C�=[}=�I=g=I�=c�=�U==��=av=;$=#�=4t=[
=��=!O=��=�x=�=�=� =�<�<�=�<[7�<*�<��<���<���<���<���<2O�<�<��<���<|D�<S��<��<�D�<;��<��<��<�<�@�<�͵<W�<cݮ<�`�<�<�^�<=ڠ<mS�<�ʙ<@�<峒<k&�<���<"�<�w�<��<[�z<��s</fl<De<N#^<�W<�O<��H<��A<�:<ŉ3<t{,<Aq%<�k<�k<�p<�{	<#�<�J�;��;���;74�;���;|!�;㲥;�W�;s�;k�{;/|a;�jG;��-;��;-��:���:���:�;:zu�9A�չ�J��&��kĺ5<�*����'�Cq>�/�T��"k�����o��E/��Р��Q����������ʻT!Ի�޻��绥y����9����}{�����T���T�(�!���%��)*�[W.�Ox2�4�6�#�:���>�˅B�,mF��IJ�N�6�Q���U��WY�0]�I�`��@d���g��\k���n��Yr���u��:y���|�M ��3���,W��l���梆��D��r䉼������������L���ᑼ0u����������%��ݲ���>���ɜ�bS��ܟ��c���ꢼ�p��~���a{������Ճ�����������#���+��T���k��ߝ��q!��e����)������*4���  �  �dN=>�M=q�L=4L=TK=E�J=u�I=I=<H=RtG=�F=��E=�E=�MD=�C=!�B=^�A=�A=�H@=tw?=#�>=��==��<=a&<=�N;=ku:=��9=C�8=2�7=e 7=�6=C;5=�U4=nn3=�2=K�1=m�0=O�/=��.=��-=��,=��+=��*=��)=��(=��'=��&=��%=�$=խ#=��"=�!=Bg =I=c'=?=��=D�=X}=�I=a=@�=`�=�U==��=ev=6$=%�=7t=c
=��="O=��=�x=�=�=� = =�<�=�<Z7�<*�<��< ��<���<���<z��<>O�<�<
��<{��<zD�<@��<��<�D�<2��<��<{�<�<�@�<�͵<W�<Qݮ<�`�<
�<�^�<:ڠ<jS�<�ʙ<@�<곒<k&�<×�<(�<�w�<��<X�z<��s<7fl<-De<R#^<�W<	�O<��H<�A<�:<Љ3<f{,<Cq%<�k<�k<�p<�{	<�<�J�;F��;���;4�;��;f!�;鲥;�W�;��;��{;�{a;�jG;{�-;��;���:g��:G��:��;:�v�9�:�mչ��J��&��lĺ�;�	����'��p>�V�T��"k������n���.���Ϡ��Q��S��������ʻR!Ի޻����y�P���9����|{�����P���T��!��%�"**�fW.�^x2�/�6�'�:���>��B�%mF��IJ��N��Q���U��WY�>]�4�`��@d���g��\k���n��Yr���u�^:y���|�G ��5���3W��a���袆��D��z䉼������������L���ᑼ0u����������%��۲���>���ɜ�hS��ܟ��c���ꢼ�p��|���k{������Ճ��z��ڊ����)���,��H���g��՝��o!��l����)������4���  �  �dN=?�M=p�L=9L=xTK=C�J=|�I=I=<H=TtG=�F=��E=�E=�MD=�C=&�B=X�A=�A=�H@=yw?=0�>=��==��<=[&<=�N;=nu:=��9=A�8=-�7=` 7=�6=L;5=�U4=on3=�2=H�1=s�0=H�/=��.=��-=}�,=��+=��*=��)=��(=��'=��&=��%=�$=ح#=��"=�!=@g =I=e'=A=��=G�=R}=�I=b=K�=f�=�U==��=gv=6$=)�=1t=]
=��=O=��=�x=�=�=� ==�<�=�<i7�<*�<��<���<���<���<~��<9O�<��<��<u��<�D�<M��<
��<�D�<$��<���<~�<���<�@�<�͵<W�<Uݮ<�`�<�<�^�<9ڠ<^S�<�ʙ<@�<ﳒ<_&�<���<�<�w�<��<K�z<��s<fl<EDe<K#^<�W<'�O<��H<ԱA<�:<Ӊ3<a{,<Vq%<�k<�k<�p<�{	<W�<�J�;*��;���; 4�;&��;w!�;��;XW�;��;g�{;�{a;�kG;2�-;�;?��:���:���:��;:�u�9�O��չ��J��%��Tlĺ�;����,�'��p>���T��"k�����o��)/��'Р��Q��R�������*ʻ<!Ի�޻���xy�P���9����v{��� ��C���T��!� �%��)*�LW.�\x2��6�H�:���>�߅B�mF��IJ� N�-�Q���U�tWY�X]�!�`��@d���g��\k��n��Yr���u�v:y���|�O ��1���0W��e��������D���䉼������������L���ᑼ'u�������%��ⲙ��>���ɜ�IS��ܟ��c���ꢼq��q���l{������ც����銭���,���3��;���s��ɝ��s!��r����)������4���  �  �dN==�M=o�L=7L=~TK=E�J=y�I=I=	<H=RtG=�F=��E=�E=�MD=�C="�B=`�A=�A=�H@=rw?=&�>=��==��<=_&<=�N;=mu:=��9=B�8=4�7=e 7=�6=J;5=�U4=ln3=�2=I�1=l�0=L�/=��.=��-=��,=��+=��*=��)=��(=��'=��&=��%=߾$=ӭ#=��"=�!=>g =I=e'===��=F�=\}=�I=a=A�=_�=�U==��=fv=5$=&�=5t=f
=��="O=��=�x=�=�=� =�<�<�=�<e7�<
*�<��<��<���<���<}��<=O�<�<��<s��<~D�<=��<
��<�D�<8��<���<u�<�<�@�<�͵<
W�<Rݮ<�`�<��<�^�<<ڠ<iS�<�ʙ<@�<곒<j&�<Ɨ�<�<�w�<��<R�z<��s<$fl<-De<K#^<�W<,�O<��H<�A<�:<̉3<^{,<Mq%<�k<�k<�p<�{	<&�<�J�;��;���;/4�;��;N!�;���;�W�;��;g�{;{{a;kG;�-;C�;���:=��:{��:1�;:"v�9F2�bչ�J�
&���kĺ-<����'��p>���T��"k������n���.���Ϡ��Q��W�������ʻE!Ի޻���y�S���9����s{�����G���T��!��%�**�hW.�ex2�%�6�4�:���>��B�"mF��IJ��N��Q���U�zWY�K]�9�`��@d���g��\k���n��Yr���u�c:y���|�J ��4���1W��b�����D���䉼������������L���ᑼ+u����������%��ײ���>���ɜ�cS��ܟ��c���ꢼ�p��w���n{������փ��w��㊭���,���/��G���q��՝��r!��o����)������4���  �  �cN=�M=&�L=�L=�RK=u�J=s�I=� I=�9H=�qG="�F=��E=E=gJD=y~C=f�B=o�A=YA=8D@=�r?=W�>=��==\�<=� <=�H;=go:=d�9=��8=f�7=N�6=w6=�35=�M4=Ef3=w|2=��1=c�0=��/=-�.=�-=I�,=�+="�*=��)=#�(=��'=��&=��%=]�$=�#=��"=�t!=�Y =F;=]=�=1�=��=�n=�:=S=�=�=BF=��=,�=�f=�=��=�d=�
=>�=�?=��=i=��=&�=� == �<n!�<�<��<��<���<��<���<-k�<�7�<#��<Ѿ�<z�<�/�<^��<��<�2�<���<9r�<��<�<]2�<7��<�J�<�Ѯ<�U�<1ק<�U�<Ҡ<%L�<1ę<�:�<F��<�"�<Δ�<�<�v�<��<��z<`�s<�jl<mJe<e+^<}W<��O<��H<��A<��:<'�3<��,<�%<B�<��<r�<f�	<Q�<o��;��;��;�}�;���;r�;��;���;�h�;q|;n:b;N/H;�Q.;@�;�C�:#��:�j�:�/?:]��9�^���͹�	G�r7���uº�?�z���&��k=�7�S��j��
���銻����\J��̪��.���r��d�ɻl�ӻ��ݻ�M����I���u��>���=�����G�X����p!��%�*�)�!.��C2��Y6��c:��b>��UB�\>F�9J���M�-�Q��xU�/Y���\��`��d�ڮg�:k���n��9r�`�u��y�؃|����ӟ��^J�������9���ى�]w�����J����C��Bّ�m������������a����8���Ü�N��ן�?_��{梼m����'x������G���N������x������8������!��䝶��!������*�������5���  �  �cN=�M=!�L=�L=�RK=p�J=v�I=� I=�9H=�qG=&�F=��E=�E=cJD=`~C=g�B=t�A=bA=;D@=�r?=V�>=��==a�<=� <=�H;=ko:=b�9=��8=g�7=V�6=o6=�35=�M4=Df3=z|2=��1=g�0=��/=-�.=��-=L�,=�+=�*=��)=�(=��'=��&=��%=_�$=�#=��"=�t!=�Y =J;=e=�=�=��=�n=�:=R=�=�=BF=��=*�=�f=�=��=�d=�
=D�=�?=��=zi=��='�=� =? �<i!�<��<��<��<���<��<���</k�<�7�<��<ܾ�<z�<�/�<]��<���<�2�<���<?r�<��<㠼<p2�<A��<�J�<�Ѯ<�U�<&ק<�U�<Ҡ<,L�<Bę<�:�<C��<�"�<ݔ�<�<�v�<��<z�z<{�s<�jl<�Je<\+^<|W<��O<��H<��A<��:<#�3<o�,<�%<R�<��<~�<R�	<_�<n��;)��;�;�}�;���;Aq�;��;筘;�h�;?q|;Z:b;G/H;IQ.;��;
C�:��:k�:Z/?:`��9TY��I�͹eG�l7���uº�?�M���&��k=�z�S��j��
���銻q���}J��/̪��.���r��f�ɻ`�ӻ�ݻ�M绱��\���]��.���=���H�@����p!��%��)��!.��C2��Y6��c:��b>��UB�k>F�HJ���M��Q��xU�/Y���\��`��d�Үg�
:k���n��9r��u�py�΃|����ڟ��]J�������9���ى�`w�����G����C��=ّ�m��2����������W����8���Ü�N��ן�<_���梼	m����3x������M���>�������������=������!��ٝ���!������*�������5���  �  �cN=�M=�L=�L=�RK=n�J=}�I=� I=�9H=�qG=&�F=��E=�E=lJD=e~C=q�B=k�A=_A=7D@=�r?=Z�>=��==f�<=� <=�H;=ho:=e�9=��8=d�7=U�6=j6=�35=�M4=Bf3=w|2=��1=g�0=��/=6�.=��-=J�,=�+=�*=��)=�(=��'=��&=��%=a�$=�#=��"=�t!=�Y =?;=g=�='�=��=�n=�:=M=�=�=CF=��=%�=�f=�=��=�d=�
=B�=�?=��=xi=��=!�=� == �<i!�<��<��<��<���<��<���<*k�<�7�<��<��<z�<�/�<\��<��<�2�<���<Sr�<��<���<j2�<0��<�J�<�Ѯ<�U�<ק<�U�<Ҡ<)L�<Dę<�:�<S��<�"�<ٔ�<�<�v�<��<g�z<x�s<�jl<�Je<N+^<�W<��O<��H<��A<��:<>�3<j�,<�%<N�<��<��<B�	<n�<N��;&��;��;�}�;���;iq�;Q�;���;�h�;�p|;C:b;�/H;Q.;ڡ;�B�:	��:�j�:50?:��9'u��f�͹�G�s6���uº)@�w��U�&��k=���S�j��
���銻�����J���˪��.��{r����ɻd�ӻބݻ�M绅�𻇅��V��Y���=�����G�)�����o!��%��)��!.��C2��Y6��c:�tb>��UB�P>F�IJ���M��Q��xU��.Y���\��`��d��g�:k���n��9r���u�qy���|����П��aJ���(����9���ى�[w�����Q����C��Rّ� m��$����������h����8���Ü��M��ן�2_���梼m����9x������S���B�����z��㏰�F������2��ڝ���!������*������5���  �  �cN=�M=�L=�L=�RK=r�J=x�I=� I=�9H=�qG=)�F=��E=~E=gJD=h~C=i�B=k�A=eA=8D@=�r?=Y�>=��==`�<=� <=�H;=eo:=_�9=��8=i�7=Q�6=n6=�35=�M4=Df3=z|2=��1=f�0=��/=1�.=��-=H�,=�+=!�*=��)=�(=��'=��&=��%=_�$=�#=��"=�t!=�Y =E;=`=	�=&�=��=�n=�:=N=�=�=BF=��=+�=�f=�=��=�d=�
=@�=�?=��=yi=��=(�=� => �<f!�<��<��<��<���<��<���<&k�<�7�<��<ھ�<z�<�/�<\��<��<�2�<���<Ar�<��<<^2�<<��<�J�<�Ѯ<�U�< ק<�U�<Ҡ<+L�<<ę<�:�<E��<�"�<Ք�<�<�v�<��<t�z<w�s<�jl<�Je<Y+^<�W<��O<��H<��A<��:<(�3<g�,<�%<Q�<��<��<E�	<`�<U��;@��;�;}�;���;~q�;�;���;
i�;q|;V:b;j/H;(Q.;z�;0C�:��:cj�:�.?:$��9�L���͹�G�.7���uº@�H��׸&��k=���S�xj��
���銻����^J��(̪��.���r��e�ɻl�ӻ�ݻ�M绪�𻀅��E��C���=�����G�F�����o!���%� �)��!.��C2��Y6��c:��b>��UB�k>F�<J���M�(�Q��xU��.Y���\��`��d�Ѯg�:k���n��9r���u�y�Ѓ|����ݟ��eJ�������9���ى�\w�����L����C��Mّ�m��#����������\����8���Ü�N��ן�9_��梼
m����8x������F���F��������鏰�@������"��ٝ���!������*������5���  �  �cN=�M=%�L=�L=�RK=p�J=u�I=� I=�9H=�qG=#�F=��E=�E=hJD=g~C=i�B=r�A=`A=7D@=�r?=V�>=��==^�<=� <=�H;=mo:=b�9=��8=j�7=O�6=t6=�35=�M4=Bf3=u|2=��1=b�0=��/=.�.=�-=K�,=�+="�*=~�)=%�(=��'=��&=��%=b�$=�#=��"=�t!=�Y =G;=f=
�=&�=��=�n=�:=Q=�=�=GF=��=+�=�f=�=��=�d=�
=A�=�?=��=}i=��='�=� =7 �<p!�<��<��<��<���<��<���<8k�<�7�<��<Ӿ�<z�<�/�<_��<��<�2�<���<Ar�<��<<m2�<<��<�J�<�Ѯ<�U�<.ק<�U�<Ҡ<(L�<>ę<�:�<8��<�"�<є�<�<�v�<��<|�z<h�s<�jl<mJe<\+^<�W<��O<��H<��A<Ƭ:<�3<��,<�%<G�<��<{�<d�	<[�<o��;��;�;�}�;���;|q�;�;ӭ�;�h�;q|;h:b;;/H;�Q.;X�;�B�:���:ek�:x/?:��9=����͹
G�B7���uºC@���ٸ&��k=�N�S��j��
���銻����WJ��X̪��.���r��g�ɻ��ӻфݻ�M绯��h���h��9���=�����G�:����
p!���%��)��!.��C2��Y6��c:��b>��UB�{>F�9J���M�#�Q��xU�/Y���\�#�`��d��g�:k���n��9r�k�u��y�ƃ|����ܟ��SJ�������9���ى�aw�����L����C��@ّ�m��%����������\����8���Ü�N��	ן�;_���梼m����'x�����E���J������}��쏰�<��������䝶��!������*�������5���  �  �cN=�M=#�L=�L=�RK=p�J=z�I=� I=�9H=�qG=(�F=��E=�E=kJD=e~C=n�B=l�A=`A=9D@=�r?=V�>=��==c�<=� <=�H;=jo:=d�9=��8=g�7=T�6=o6=�35=�M4=Bf3=z|2=��1=g�0=��/=1�.=��-=K�,=�+=!�*=��)=!�(=��'=��&=��%=c�$=�#=��"=�t!=�Y =B;=d=
�=&�=��=�n=�:=P=�=�=GF=��=+�=�f=�=��=�d=�
=B�=�?=��=zi=��=(�=� =; �<i!�<��<��<��<���<��<���</k�<�7�<��<ܾ�<z�<�/�<^��<��<�2�<���<Kr�<��<���<f2�<5��<�J�<�Ѯ<�U�<%ק<�U�<Ҡ<(L�<;ę<�:�<G��<�"�<Ԕ�<�<�v�<��<j�z<|�s<�jl<�Je<Q+^<�W<��O<��H<��A<��:<'�3<z�,<�%<J�<��<��<S�	<[�<f��;9��;��;�}�;���;kq�;7�;���;�h�; q|;]:b;</H;]Q.;��; C�:���:�j�:�/?:���9dY��,�͹pG�{7���uº(@�R��߸&��k=���S�uj��
���銻����bJ��#̪��.���r��f�ɻx�ӻɄݻ�M绣��k���N��P���=�����G�6�����o!���%��)��!.��C2��Y6��c:��b>��UB�g>F�:J���M��Q��xU��.Y���\��`��d�Ԯg�:k���n��9r�~�u�wy�҃|����֟��\J�������9���ى�bw�����L����C��Lّ�	m��%����������c����8���Ü�N��ן�2_���梼m����-x������K���G���������쏰�E������"��ٝ���!������*�������5���  �  �cN=�M=�L=�L=�RK=m�J=y�I=� I=�9H=�qG=)�F=��E=�E=kJD=^~C=n�B=l�A=fA=7D@=�r?=[�>=��==b�<=� <=�H;=jo:=_�9=��8=c�7=U�6=j6=�35=�M4=Bf3=y|2=��1=h�0=��/=8�.=��-=J�,=	�+=�*=��)=�(=��'=��&=��%=`�$=�#=��"=�t!=�Y =C;=e=�="�=��=�n=�:=J=�=�=CF=��='�=�f=�=��=�d=�
=B�=�?=��=vi=��=!�=� =< �<g!�<��<��<��<���<��<���<,k�<�7�<��<۾�<z�<�/�<]��<��<�2�<���<Jr�<��<�<f2�<:��<�J�<�Ѯ<�U�<ק<�U�<Ҡ<+L�<Eę<�:�<G��<�"�<ܔ�<�<�v�<��<g�z<��s<�jl<�Je<K+^<�W<��O<��H<��A<��:<(�3<f�,<�%<V�<��<��<>�	<t�<C��;<��;�;�}�;���;5q�;6�;���;i�;q|;H:b;�/H;Q.;��;�B�:D��:�j�:�.?:��9�{��<�͹�G��6���uº8@�`��j�&��k=���S�j��
���銻����{J��.̪�/��ur��x�ɻ��ӻ�ݻ�M绊�𻝅��?��L���=����H�5�����o!��%��)��!.��C2��Y6��c:�nb>��UB�q>F�FJ���M��Q��xU��.Y���\��`��d�ݮg�:k���n��9r���u�oy�݃|����ޟ��_J���&����9���ى�[w�����R����C��Nّ�
m��2����������^����8���Ü��M��ן�6_���梼
m����8x������T���?��������ߏ��F������7��՝���!������*������5���  �  �cN=�M=!�L=�L=�RK=r�J=y�I=� I=�9H=�qG=%�F=��E=�E=iJD=i~C=l�B=m�A=_A=7D@=�r?=W�>=��==c�<=� <=�H;=io:=b�9=��8=g�7=Q�6=p6=�35=�M4=Bf3={|2=��1=h�0=��/=2�.=��-=J�,=�+="�*=��)= �(=��'=��&=��%=b�$=�#=��"=�t!=�Y =D;=d=�=(�=��=�n=�:=P=�=�=EF=��=*�=�f=�=��=�d=�
=A�=�?=��=wi=��=&�=� =: �<d!�<��<��<��<���<��<���<0k�<�7�<��<ݾ�<	z�<�/�<`��<��<�2�<���<Hr�<��<�<h2�<8��<�J�<�Ѯ<�U�<%ק<�U�<Ҡ<)L�<<ę<�:�<H��<�"�<Д�<�<�v�<��<d�z<��s<�jl<�Je<G+^<�W<��O<��H<��A<��:<+�3<o�,<�%<H�<��<��<P�	<h�<Y��;��;��;�}�;���;�q�;$�;���;�h�;q|;n:b;W/H;MQ.;��;HC�:���:�j�:g/?:B��9*Z����͹G��6��vºG@�=���&��k=���S�fj��
���銻����UJ��,̪��.���r��i�ɻk�ӻτݻ�M绚��q���[��F���=�����G�8�����o!���%��)��!.��C2��Y6��c:��b>��UB�m>F�4J���M�!�Q��xU��.Y���\��`��d�Үg�:k���n��9r�y�u�}y�Ӄ|����ڟ��[J�������9���ى�`w�����M����C��Iّ�m������������`����8���Ü� N��ן�4_��~梼m����2x������I���K������~��돰�H������*��֝���!������*�������5���  �  �cN=�M=!�L=�L=�RK=s�J=s�I=� I=�9H=�qG=(�F=��E=�E=dJD=k~C=g�B=r�A=_A=:D@=�r?=V�>=��==[�<=� <=�H;=io:=a�9=��8=k�7=P�6=q6=�35=�M4=Df3=x|2=��1=d�0=��/=/�.=��-=J�,=�+=%�*=�)= �(=��'=��&=��%=`�$=�#=��"=�t!=�Y =H;=b=�=&�=��=�n=�:=T=�=�=EF=��=/�=�f=�=��=�d=�
=A�=�?=��=}i=��=%�=� => �<o!�<~�<��<��<���<��<���<0k�<�7�<%��<Ͼ�<z�<�/�<`��<���<�2�<���<=r�<��<蠼<h2�<=��<�J�<�Ѯ<�U�<-ק<�U�<Ҡ<0L�<<ę<�:�<=��<�"�<Д�<�<�v�<��<{�z<r�s<�jl<|Je<]+^<�W<��O<��H<��A<ά:<�3<p�,<�%<S�<��<r�<_�	<Y�<��;7��;�;�}�;���;�q�;��;׭�;�h�;6q|;�:b;H/H;wQ.;2�;�C�:¤�:�j�:9/?:r��9S9��؍͹�
G��7���uº�?�j���&��k=�O�S��j��
���銻����BJ��N̪��.���r��D�ɻ��ӻ�ݻ�M绷��M���a��6���=�����G�I����p!��%��)��!.��C2��Y6��c:��b>��UB�z>F�1J���M�$�Q��xU�/Y���\��`��d�خg�:k���n��9r�w�u��y�ƃ|����ݟ��\J�������9���ى�^w�����G����C��@ّ�m������������[����8���Ü�
N��
ן�@_���梼m����2x������?���K���������鏰�<������$��ݝ���!������*�������5���  �  �cN=�M=#�L=�L=�RK=m�J=y�I=� I=�9H=�qG=(�F=��E=�E=jJD=i~C=j�B=p�A=aA=8D@=�r?=X�>=��==a�<=� <=�H;=jo:=c�9=��8=e�7=P�6=n6=�35=�M4==f3=x|2=��1=c�0=��/=6�.=��-=I�,=�+=�*=��)=!�(=��'=��&=��%=a�$=�#=��"=�t!=�Y =B;=f=�=(�=��=�n=�:=N=�=�=EF=��='�=�f=�=��=�d=�
=@�=�?=��=yi=��=&�=� =2 �<k!�<��<��<��<���<��<���<1k�<�7�<��<۾�<z�<�/�<Y��<��<�2�<���<Er�<��<���<j2�<6��<�J�<�Ѯ<�U�<*ק<�U�<Ҡ<"L�<Bę<�:�<A��<�"�<֔�<�<�v�<��<_�z<q�s<�jl<|Je<A+^<�W<��O<��H<��A<��:< �3<z�,<�%<D�<��<��<Y�	<d�<O��;6��;��;�}�;���;�q�;�;ĭ�;�h�;q|;1:b;b/H;rQ.;��;�B�:���:k�:�/?:o��9=h����͹�G��6���uº�@�i����&��k=���S�j��
���銻����xJ��/̪��.���r����ɻ��ӻلݻ�M绩��y���[��L���=�����G�9���� p!���%��)��!.��C2��Y6��c:��b>��UB�k>F�GJ���M�'�Q��xU��.Y���\��`��d�خg�$:k���n��9r���u��y�׃|����ן��[J���&����9���ى�^w�����L����C��Fّ�m������������b����8���Ü�N��ן�6_���梼m����.x������O���F��������Ᏸ�J������$��ݝ���!������*�� ����5���  �  �cN=�M=�L=�L=�RK=o�J=�I=� I=�9H=�qG=,�F=��E=�E=hJD=a~C=k�B=m�A=dA=:D@=�r?=Z�>=��==i�<=� <=�H;=io:=a�9=��8=e�7=U�6=m6=�35=�M4=Df3=||2=��1=m�0=��/=1�.=��-=J�,=	�+=�*=��)=�(=��'=��&=��%=a�$=�#=��"=�t!=�Y =C;=f=�=!�=��=�n=�:=M=�=�=BF=��='�=�f=�=��=�d=�
=C�=�?=��=ti=��=&�=� =? �<_!�<��<��<��<���<��<���<(k�<�7�<��<��<�y�<�/�<\��<��<�2�<���<Hr�<��<<g2�<<��<�J�<�Ѯ<�U�<ק<�U�<Ҡ<(L�<Bę<�:�<M��<�"�<ٔ�<�<�v�<��<c�z<��s<�jl<�Je<L+^<{W<��O<��H<��A<��:<5�3<g�,<
�%<P�<��<��<=�	<q�<;��;Y��;�;�}�;���;Hq�;�;���;i�;;q|;7:b;z/H;Q.;�;B�:K��:�j�:(/?:ܶ�9i��Y�͹
G�C7��lvº�?�%����&�?k=���S�xj��
���銻����}J��̪�/���r����ɻN�ӻ؄ݻ�M绌�𻋅��<��H���=����H�3�����o!��%��)��!.��C2��Y6��c:�ub>�VB�[>F�FJ���M��Q��xU��.Y��\��`��d�ˮg�	:k���n��9r���u�my�Ӄ|����ן��cJ���%����9���ى�]w�����K����C��Jّ�m��/����������]����8���Ü��M��ן�-_��~梼m����7x������Q���B��������폰�I������+��ҝ���!������*������5���  �  �cN=�M=!�L=�L=�RK=p�J=x�I=� I=�9H=�qG='�F=��E=�E=iJD=i~C=l�B=q�A=\A=8D@=�r?=\�>=��==a�<=� <=�H;=ko:=c�9=��8=h�7=P�6=q6=�35=�M4=Ff3=r|2=��1=c�0=��/=1�.=�-=J�,=�+=�*=��)= �(=��'=��&=��%=_�$=�#=��"=�t!=�Y =D;=f=�='�=��=�n=�:=O=�=�=BF=��=)�=�f=�=��=�d=�
=@�=�?=��=i=��=�=� => �<t!�<��<��<��<���<��<���<0k�<�7�<��<ھ�<z�<�/�<b��<��<�2�<���<Hr�<��<�<k2�<7��<�J�<�Ѯ<�U�<%ק<�U�<Ҡ<,L�<Aę<�:�<C��<�"�<Ҕ�<�<�v�<��<��z<g�s<�jl<kJe<g+^<�W<��O<��H<��A<��:<�3<s�,<�%<S�<��<��<M�	<s�<a��;-��;��;�}�;���;�q�;#�;ϭ�;�h�;q|;n:b;�/H;7Q.;��;�B�:���:k�:�/?:���9(T����͹�
G�p7��>uº�?����y�&��k=�4�S�vj��
���銻����pJ��&̪��.���r��r�ɻy�ӻ�ݻ�M绊��u���c��E���=�����G�3����p!���%��)��!.��C2��Y6��c:��b>��UB�d>F�GJ���M�%�Q��xU��.Y���\��`��d��g�:k�z�n��9r�u�u��y�΃|����՟��[J���"����9���ى�Vw�����M����C��Eّ�m�� ����������b����8���Ü��M��ן�8_���梼	m����0x������J���I������}��台�7������3��坶��!������*�������5���  �  �cN=�M=&�L=�L=�RK=t�J=z�I=� I=�9H=�qG=(�F=��E=�E=eJD=i~C=e�B=t�A=]A==D@=�r?=T�>=��==b�<=� <=�H;=ho:=d�9=��8=m�7=L�6=s6=�35=�M4=<f3={|2=��1=_�0=��/=*�.= �-=J�,=	�+=!�*=�)=$�(=��'=��&=��%=b�$=�#=��"=�t!=�Y =G;=d=	�=%�=��=�n=�:=V=�=�=FF=��=,�=�f=�=��=�d=�
=>�=�?=�=~i=��=3�=� =+ �<k!�<y�<��<
��<���<��<���</k�<�7�<"��<��<z�<�/�<\��<���<�2�<���<>r�<��<�<n2�<8��<�J�<�Ѯ<�U�<&ק<�U�<Ҡ<$L�<5ę<�:�<:��<�"�<є�<�<�v�<��<l�z<g�s<kl<wJe<G+^<yW<��O<��H<��A<ͬ:<�3<��,<��%<<�<��<��<V�	<S�<���;7��;��;�}�;���;�q�;��;歘;�h�;mq|;e:b;#/H;iQ.;��;�C�:��:�j�:0?:��9],��׏͹p
G��7���uº�@�3���&�l=�K�S��j��
���銻����aJ��O̪��.���r��j�ɻ\�ӻфݻ�M����9���h��9���=����H�C����p!�޷%�(�)��!.��C2��Y6��c:��b>��UB�v>F�GJ���M�.�Q��xU�/Y���\�1�`�dd���g�1:k���n��9r�j�u��y���|����֟��\J��"�����9���ى�fw�����?����C��>ّ�m������������`����8���Ü�N��ן�5_��}梼m����(x������B���K�������������D������ ��ߝ���!������*�������5���  �  �cN=�M=!�L=�L=�RK=p�J=x�I=� I=�9H=�qG='�F=��E=�E=iJD=i~C=k�B=q�A=\A=8D@=�r?=\�>=��==a�<=� <=�H;=ko:=c�9=��8=h�7=P�6=q6=�35=�M4=Ff3=r|2=��1=c�0=��/=1�.=�-=J�,=�+=�*=��)= �(=��'=��&=��%=_�$=�#=��"=�t!=�Y =D;=f=�='�=��=�n=�:=O=�=�=BF=��=)�=�f=�=��=�d=�
=@�=�?=��=i=��=�=� => �<t!�<��<��<��<���<��<���<0k�<�7�<��<ھ�<z�<�/�<b��<��<�2�<���<Hr�<��<�<k2�<7��<�J�<�Ѯ<�U�<%ק<�U�<Ҡ<,L�<Aę<�:�<C��<�"�<Ҕ�<�<�v�<��<��z<g�s<�jl<kJe<g+^<�W<��O<��H<��A<��:<�3<s�,<�%<S�<��<��<M�	<s�<a��;-��;��;�}�;���;�q�;#�;ϭ�;�h�;q|;n:b;�/H;7Q.;��;�B�:���:k�:�/?:���9-T����͹�
G�q7��>uº�?����y�&��k=�4�S�vj��
���銻����pJ��&̪��.���r��r�ɻy�ӻ�ݻ�M绊��u���c��E���=�����G�3����p!���%��)��!.��C2��Y6��c:��b>��UB�d>F�GJ���M�%�Q��xU��.Y���\��`��d��g�:k�z�n��9r�u�u��y�΃|����՟��[J���"����9���ى�Vw�����M����C��Eّ�m�� ����������b����8���Ü��M��ן�8_���梼	m����0x������J���I������}��台�7������3��坶��!������*�������5���  �  �cN=�M=�L=�L=�RK=o�J=�I=� I=�9H=�qG=,�F=��E=�E=hJD=a~C=k�B=m�A=dA=:D@=�r?=Z�>=��==i�<=� <=�H;=io:=a�9=��8=e�7=U�6=m6=�35=�M4=Df3=||2=��1=m�0=��/=1�.=��-=J�,=	�+=�*=��)=�(=��'=��&=��%=a�$=�#=��"=�t!=�Y =C;=f=�=!�=��=�n=�:=M=�=�=BF=��='�=�f=�=��=�d=�
=C�=�?=��=ti=��=&�=� =? �<_!�<��<��<��<���<��<���<(k�<�7�<��<��<�y�<�/�<\��<��<�2�<���<Hr�<��<<g2�<<��<�J�<�Ѯ<�U�<ק<�U�<Ҡ<(L�<Bę<�:�<M��<�"�<ٔ�<�<�v�<��<c�z<��s<�jl<�Je<L+^<{W<��O<��H<��A<��:<5�3<g�,<
�%<P�<��<��<=�	<q�<;��;Y��;�;�}�;���;Hq�;�;���;i�;;q|;7:b;z/H;Q.;�;B�:K��:�j�:(/?:ܶ�9i��Z�͹
G�C7��lvº�?�%����&�?k=���S�xj��
���銻����}J��̪�/���r����ɻN�ӻ؄ݻ�M绌�𻋅��<��H���=����H�3�����o!��%��)��!.��C2��Y6��c:�ub>�VB�[>F�FJ���M��Q��xU��.Y��\��`��d�ˮg�	:k���n��9r���u�my�Ӄ|����ן��cJ���%����9���ى�]w�����K����C��Jّ�m��/����������]����8���Ü��M��ן�-_��~梼m����7x������Q���B��������폰�I������+��ҝ���!������*������5���  �  �cN=�M=#�L=�L=�RK=m�J=y�I=� I=�9H=�qG=(�F=��E=�E=jJD=i~C=j�B=p�A=aA=8D@=�r?=X�>=��==a�<=� <=�H;=jo:=c�9=��8=e�7=P�6=n6=�35=�M4==f3=x|2=��1=c�0=��/=6�.=��-=I�,=�+=�*=��)=!�(=��'=��&=��%=a�$=�#=��"=�t!=�Y =B;=f=�=(�=��=�n=�:=N=�=�=EF=��='�=�f=�=��=�d=�
=@�=�?=��=yi=��=&�=� =2 �<k!�<��<��<��<���<��<���<1k�<�7�<��<۾�<z�<�/�<Y��<��<�2�<���<Er�<��<���<j2�<6��<�J�<�Ѯ<�U�<*ק<�U�<Ҡ<"L�<Bę<�:�<A��<�"�<֔�<�<�v�<��<_�z<q�s<�jl<|Je<A+^<�W<��O<��H<��A<��:< �3<z�,<�%<D�<��<��<Y�	<d�<O��;6��;��;�}�;���;�q�;�;ĭ�;�h�;q|;1:b;b/H;rQ.;��;�B�:���:k�:�/?:o��9Eh����͹�G��6���uº�@�i����&��k=���S�j��
���銻����xJ��/̪��.���r����ɻ��ӻلݻ�M绩��y���[��L���=�����G�9���� p!���%��)��!.��C2��Y6��c:��b>��UB�k>F�GJ���M�'�Q��xU��.Y���\��`��d�خg�$:k���n��9r���u��y�׃|����ן��[J���&����9���ى�^w�����L����C��Fّ�m������������b����8���Ü�N��ן�6_���梼m����.x������O���F��������Ᏸ�J������$��ݝ���!������*�� ����5���  �  �cN=�M=!�L=�L=�RK=s�J=s�I=� I=�9H=�qG=(�F=��E=�E=dJD=k~C=g�B=r�A=_A=:D@=�r?=V�>=��==[�<=� <=�H;=io:=a�9=��8=k�7=P�6=q6=�35=�M4=Df3=x|2=��1=d�0=��/=/�.=��-=J�,=�+=%�*=�)= �(=��'=��&=��%=`�$=�#=��"=�t!=�Y =H;=b=�=&�=��=�n=�:=T=�=�=EF=��=/�=�f=�=��=�d=�
=A�=�?=��=}i=��=%�=� => �<o!�<~�<��<��<���<��<���<0k�<�7�<%��<Ͼ�<z�<�/�<`��<���<�2�<���<=r�<��<蠼<h2�<=��<�J�<�Ѯ<�U�<-ק<�U�<Ҡ<0L�<<ę<�:�<=��<�"�<Д�<�<�v�<��<{�z<r�s<�jl<|Je<]+^<�W<��O<��H<��A<ά:<�3<p�,<�%<S�<��<r�<_�	<Y�<��;7��;�;�}�;���;�q�;��;׭�;�h�;6q|;�:b;H/H;wQ.;2�;�C�:¤�:�j�:9/?:q��9d9��ٍ͹�
G��7���uº�?�j���&��k=�O�S��j��
���銻����BJ��N̪��.���r��D�ɻ��ӻ�ݻ�M绷��M���a��6���=�����G�I����p!��%��)��!.��C2��Y6��c:��b>��UB�z>F�1J���M�$�Q��xU�/Y���\��`��d�خg�:k���n��9r�w�u��y�ƃ|����ݟ��\J�������9���ى�^w�����G����C��@ّ�m������������[����8���Ü�
N��
ן�@_���梼m����2x������?���K���������鏰�<������$��ݝ���!������*�������5���  �  �cN=�M=!�L=�L=�RK=r�J=y�I=� I=�9H=�qG=%�F=��E=�E=iJD=i~C=l�B=m�A=_A=7D@=�r?=W�>=��==c�<=� <=�H;=io:=b�9=��8=g�7=Q�6=p6=�35=�M4=Bf3={|2=��1=h�0=��/=2�.=��-=J�,=�+="�*=��)= �(=��'=��&=��%=b�$=�#=��"=�t!=�Y =D;=d=�=(�=��=�n=�:=P=�=�=EF=��=*�=�f=�=��=�d=�
=A�=�?=��=wi=��=&�=� =: �<d!�<��<��<��<���<��<���<0k�<�7�<��<ݾ�<	z�<�/�<`��<��<�2�<���<Hr�<��<�<h2�<8��<�J�<�Ѯ<�U�<%ק<�U�<Ҡ<)L�<<ę<�:�<H��<�"�<Д�<�<�v�<��<d�z<��s<�jl<�Je<G+^<�W<��O<��H<��A<��:<+�3<o�,<�%<H�<��<��<P�	<h�<Y��;��;��;�}�;���;�q�;$�;���;�h�;q|;n:b;W/H;MQ.;��;HC�:���:�j�:g/?:@��99Z����͹G��6��vºG@�>���&��k=���S�fj��
���銻����UJ��,̪��.���r��i�ɻl�ӻτݻ�M绚��q���[��F���=�����G�8�����o!���%��)��!.��C2��Y6��c:��b>��UB�m>F�4J���M�!�Q��xU��.Y���\��`��d�Үg�:k���n��9r�y�u�}y�Ӄ|����ڟ��[J�������9���ى�`w�����M����C��Iّ�m������������`����8���Ü� N��ן�4_��~梼m����2x������I���K������~��돰�H������*��֝���!������*�������5���  �  �cN=�M=�L=�L=�RK=m�J=y�I=� I=�9H=�qG=)�F=��E=�E=kJD=^~C=n�B=l�A=fA=7D@=�r?=[�>=��==b�<=� <=�H;=jo:=_�9=��8=c�7=U�6=j6=�35=�M4=Bf3=y|2=��1=h�0=��/=8�.=��-=J�,=	�+=�*=��)=�(=��'=��&=��%=`�$=�#=��"=�t!=�Y =C;=e=�="�=��=�n=�:=J=�=�=CF=��='�=�f=�=��=�d=�
=B�=�?=��=vi=��=!�=� =< �<g!�<��<��<��<���<��<���<,k�<�7�<��<۾�<z�<�/�<]��<��<�2�<���<Jr�<��<�<f2�<:��<�J�<�Ѯ<�U�<ק<�U�<Ҡ<+L�<Eę<�:�<G��<�"�<ܔ�<�<�v�<��<g�z<��s<�jl<�Je<K+^<�W<��O<��H<��A<��:<(�3<f�,<�%<V�<��<��<>�	<t�<C��;<��;�;�}�;���;5q�;6�;���;i�;q|;H:b;�/H;Q.;��;�B�:D��:�j�:�.?:��9�{��=�͹�G��6���uº8@�`��j�&��k=���S�j��
���銻����{J��.̪�/��ur��x�ɻ��ӻ�ݻ�M绊�𻝅��?��L���=����H�5�����o!��%��)��!.��C2��Y6��c:�nb>��UB�q>F�FJ���M��Q��xU��.Y���\��`��d�ݮg�:k���n��9r���u�oy�݃|����ޟ��_J���&����9���ى�[w�����R����C��Nّ�
m��2����������^����8���Ü��M��ן�6_���梼
m����8x������T���?��������ߏ��F������7��՝���!������*������5���  �  �cN=�M=#�L=�L=�RK=p�J=z�I=� I=�9H=�qG=(�F=��E=�E=kJD=e~C=n�B=l�A=`A=9D@=�r?=V�>=��==c�<=� <=�H;=jo:=d�9=��8=g�7=T�6=o6=�35=�M4=Bf3=z|2=��1=g�0=��/=1�.=��-=K�,=�+=!�*=��)=!�(=��'=��&=��%=c�$=�#=��"=�t!=�Y =B;=d=
�=&�=��=�n=�:=P=�=�=GF=��=+�=�f=�=��=�d=�
=B�=�?=��=zi=��=(�=� =; �<i!�<��<��<��<���<��<���</k�<�7�<��<ܾ�<z�<�/�<^��<��<�2�<���<Kr�<��<���<f2�<5��<�J�<�Ѯ<�U�<%ק<�U�<Ҡ<(L�<;ę<�:�<G��<�"�<Ԕ�<�<�v�<��<j�z<|�s<�jl<�Je<Q+^<�W<��O<��H<��A<��:<'�3<z�,<�%<J�<��<��<S�	<[�<f��;9��;��;�}�;���;kq�;7�;���;�h�; q|;]:b;</H;]Q.;��; C�:���:�j�:�/?:���9{Y��-�͹pG�|7���uº(@�S��߸&��k=���S�uj��
���銻����bJ��#̪��.���r��f�ɻx�ӻɄݻ�M绣��k���N��P���=�����G�6�����o!���%��)��!.��C2��Y6��c:��b>��UB�g>F�:J���M��Q��xU��.Y���\��`��d�Ԯg�:k���n��9r�~�u�wy�҃|����֟��\J�������9���ى�bw�����L����C��Lّ�	m��%����������c����8���Ü�N��ן�2_���梼m����-x������K���G���������쏰�E������"��ٝ���!������*�������5���  �  �cN=�M=%�L=�L=�RK=p�J=u�I=� I=�9H=�qG=#�F=��E=�E=hJD=g~C=i�B=r�A=`A=7D@=�r?=V�>=��==^�<=� <=�H;=mo:=b�9=��8=j�7=O�6=t6=�35=�M4=Bf3=u|2=��1=b�0=��/=.�.=�-=K�,=�+="�*=~�)=%�(=��'=��&=��%=b�$=�#=��"=�t!=�Y =G;=f=
�=&�=��=�n=�:=Q=�=�=GF=��=+�=�f=�=��=�d=�
=A�=�?=��=}i=��='�=� =7 �<p!�<��<��<��<���<��<���<8k�<�7�<��<Ӿ�<z�<�/�<_��<��<�2�<���<Ar�<��<<m2�<<��<�J�<�Ѯ<�U�<.ק<�U�<Ҡ<(L�<>ę<�:�<8��<�"�<є�<�<�v�<��<|�z<h�s<�jl<mJe<\+^<�W<��O<��H<��A<Ƭ:<�3<��,<�%<G�<��<{�<d�	<[�<o��;��;�;�}�;���;|q�;�;ӭ�;�h�;q|;h:b;;/H;�Q.;X�;�B�:���:ek�:x/?:
��9=����͹
G�C7���uºC@���ڸ&��k=�N�S��j��
���銻����WJ��X̪��.���r��g�ɻ��ӻфݻ�M绯��h���h��9���=�����G�:����
p!���%��)��!.��C2��Y6��c:��b>��UB�{>F�9J���M�#�Q��xU�/Y���\�#�`��d��g�:k���n��9r�k�u��y�ƃ|����ܟ��SJ�������9���ى�aw�����L����C��@ّ�m��%����������\����8���Ü�N��	ן�;_���梼m����'x�����E���J������}��쏰�<��������䝶��!������*�������5���  �  �cN=�M=�L=�L=�RK=r�J=x�I=� I=�9H=�qG=)�F=��E=~E=gJD=h~C=i�B=k�A=eA=8D@=�r?=Y�>=��==`�<=� <=�H;=eo:=_�9=��8=i�7=Q�6=n6=�35=�M4=Df3=z|2=��1=f�0=��/=1�.=��-=H�,=�+=!�*=��)=�(=��'=��&=��%=_�$=�#=��"=�t!=�Y =E;=`=	�=&�=��=�n=�:=N=�=�=BF=��=+�=�f=�=��=�d=�
=@�=�?=��=yi=��=(�=� => �<f!�<��<��<��<���<��<���<&k�<�7�<��<ھ�<z�<�/�<\��<��<�2�<���<Ar�<��<<^2�<<��<�J�<�Ѯ<�U�< ק<�U�<Ҡ<+L�<<ę<�:�<E��<�"�<Ք�<�<�v�<��<t�z<w�s<�jl<�Je<Y+^<�W<��O<��H<��A<��:<(�3<g�,<�%<Q�<��<��<E�	<`�<V��;@��;�;}�;���;~q�;�;���;
i�;q|;V:b;i/H;(Q.;z�;0C�:��:cj�:�.?:#��9�L����͹�G�.7���uº@�H��׸&��k=���S�xj��
���銻����^J��(̪��.���r��e�ɻl�ӻ�ݻ�M绪�𻀅��E��C���=�����G�F�����o!���%� �)��!.��C2��Y6��c:��b>��UB�k>F�<J���M�(�Q��xU��.Y���\��`��d�Ѯg�:k���n��9r���u�y�Ѓ|����ݟ��eJ�������9���ى�\w�����L����C��Mّ�m��#����������\����8���Ü�N��ן�9_��梼
m����8x������F���F��������鏰�@������"��ٝ���!������*������5���  �  �cN=�M=�L=�L=�RK=n�J=}�I=� I=�9H=�qG=&�F=��E=�E=lJD=e~C=q�B=k�A=_A=7D@=�r?=Z�>=��==f�<=� <=�H;=ho:=e�9=��8=d�7=U�6=j6=�35=�M4=Bf3=w|2=��1=g�0=��/=6�.=��-=J�,=�+=�*=��)=�(=��'=��&=��%=a�$=�#=��"=�t!=�Y =?;=g=�='�=��=�n=�:=M=�=�=CF=��=%�=�f=�=��=�d=�
=B�=�?=��=xi=��=!�=� == �<i!�<��<��<��<���<��<���<*k�<�7�<��<��<z�<�/�<\��<��<�2�<���<Sr�<��<���<j2�<0��<�J�<�Ѯ<�U�<ק<�U�<Ҡ<)L�<Dę<�:�<S��<�"�<ٔ�<�<�v�<��<g�z<x�s<�jl<�Je<N+^<�W<��O<��H<��A<��:<>�3<j�,<�%<N�<��<��<B�	<n�<N��;&��;��;�}�;���;iq�;Q�;���;�h�;�p|;C:b;�/H;Q.;ڡ;�B�:	��:�j�:50?:��96u��f�͹�G�s6���uº*@�w��U�&��k=���S�j��
���銻�����J���˪��.��{r����ɻd�ӻބݻ�M绅�𻇅��V��Y���=�����G�)�����o!��%��)��!.��C2��Y6��c:�tb>��UB�P>F�IJ���M��Q��xU��.Y���\��`��d��g�:k���n��9r���u�qy���|����П��aJ���(����9���ى�[w�����Q����C��Rّ� m��$����������h����8���Ü��M��ן�2_���梼m����9x������S���B�����z��㏰�F������2��ڝ���!������*������5���  �  �cN=�M=!�L=�L=�RK=p�J=v�I=� I=�9H=�qG=&�F=��E=�E=cJD=`~C=g�B=t�A=bA=;D@=�r?=V�>=��==a�<=� <=�H;=ko:=b�9=��8=g�7=V�6=o6=�35=�M4=Df3=z|2=��1=g�0=��/=-�.=��-=L�,=�+=�*=��)=�(=��'=��&=��%=_�$=�#=��"=�t!=�Y =J;=e=�=�=��=�n=�:=R=�=�=BF=��=*�=�f=�=��=�d=�
=D�=�?=��=zi=��='�=� =? �<i!�<��<��<��<���<��<���</k�<�7�<��<ܾ�<z�<�/�<]��<���<�2�<���<?r�<��<㠼<p2�<A��<�J�<�Ѯ<�U�<&ק<�U�<Ҡ<,L�<Bę<�:�<C��<�"�<ݔ�<�<�v�<��<z�z<{�s<�jl<�Je<\+^<|W<��O<��H<��A<��:<#�3<o�,<�%<R�<��<~�<R�	<_�<n��;)��;�;�}�;���;Aq�;��;筘;�h�;?q|;Z:b;G/H;IQ.;��;
C�:��:k�:Z/?:_��9QY��I�͹eG�l7���uº�?�M���&��k=�z�S��j��
���銻q���}J��/̪��.���r��f�ɻ`�ӻ�ݻ�M绱��\���]��.���=���H�@����p!��%��)��!.��C2��Y6��c:��b>��UB�k>F�HJ���M��Q��xU�/Y���\��`��d�Ѯg�
:k���n��9r��u�py�σ|����ڟ��]J�������9���ى�`w�����G����C��=ّ�m��2����������W����8���Ü�N��ן�<_���梼	m����3x������M���>�������������=������!��ٝ���!������*�������5���  �  �bN=1�M=�L=�L=�QK=�J=��I=6�H=�7H=�oG=�F=y�E=E=�GD=�{C=�B=f�A=&A=�@@=Ro?=��>=��==B�<=�<=^D;=�j:=��9=��8=&�7=��6=�6=�-5=�G4=�_3=�u2=��1=Z�0=��/=��.=T�-=X�,=��+=��*=��)=L�(=��'=n�&=�%=��$= �#=d�"=vj!=*O =�0=�=�=��=Q�=c=,/=��=B�=/}=L:=��=�=�Z=�=��=�X=��	=E�=�3=��=�]=�=�x=�  =�	�<q�<��<���<;��<|��<��<M��<[X�<3%�<Y��<���<\i�<��<���<}�<Z$�<��<Ae�<g��<D��<h'�<䵵<�@�<�Ȯ<xM�<zϧ<�N�<�ˠ<}F�<F��<G6�<���<��<���<��<�u�<S�<T�z<��s<Pnl<GOe<�1^<!W<��O<)�H<=�A<ƹ:<\�3<�,<��%<q�<T�<P�<�	<��<���; �;�S�;��;p*�;���;�F�;��;O��;% };s�b;��H;'�.;�B;i��:D��:�Œ:��A:2X�9)�0���ǹ�D�޵���������u���%�0�<�S� Mi��F�M����A��o⟻rd��Ǵ�Z���0ɻ�6ӻ1ݻ��滆��"��N���r������K�_������C!�m�%�x�)���-��2��16��<:�a<>��0B�F���I�A�M���Q�XU�aY�H�\�~b`���c��g�=k���n� r�$�u�Fy�?m|�&��p���R@���脼�����0��8щ�Uo��3�������<���ґ��f��������W��M���4��w����I��1ӟ��[��%㢼j��#𥼦u������>���������6������@������𝶼"�������+������7���  �  �bN=2�M=�L=�L=�QK=�J=��I=9�H=�7H=�oG=�F=x�E=E=�GD=�{C=��B=`�A=(A=�@@=Vo?=��>=��==E�<=�<=gD;=�j:=|�9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=É1=a�0=��/=��.=D�-=V�,=��+=��*=��)=D�(=��'=n�&=�%=��$="�#=i�"=xj!=2O =�0=�=��=�=T�=c=3/=��=G�=2}=Q:=��=�=�Z=�=~�=�X=��	=E�=�3=��=�]=�=�x=�  =�	�<j�<��<z��<G��<p��<��<>��<MX�<E%�<L��<���<di�<��<���<}�<a$�<��<Ie�<K��<@��<e'�<޵�<�@�<�Ȯ<�M�<�ϧ<�N�<�ˠ<�F�<J��<96�<���<��<���<v�<�u�<Q�<Y�z<��s<]nl<oOe<�1^<W<i�O<	�H<]�A<��:<`�3<��,<��%<��<4�<d�<��	<��<	��;j �;�S�;ض�;x*�;���;�F�;��;Z��;� };��b;��H;i�.;�B;g��:m��:�Ē:��A:\V�9�51�4�ǹ�D����:����������%���<�,S�)Mi��G�]����A���⟻{d��^Ǵ�'���0ɻ7ӻݻ���^��"��,���r������m�V������C!�`�%�b�)���-��2��16��<:�?<>��0B�'F���I�I�M���Q�PXU�rY�R�\�cb`���c���g�-k���n�� r�X�u�.y�Xm|�>�����`@��y脼퍆��0��0щ�Mo��(��癩��<���ґ��f��,������Y��S����3��s����I��*ӟ��[��1㢼j�� 𥼵u������R���������R��򎰼���,������ݝ��"�������+�����7���  �  �bN=<�M=�L=�L=�QK=��J=��I=1�H=�7H=�oG=	�F=t�E=E=�GD=�{C=��B=[�A=&A=�@@=Po?=��>=��==J�<=�<=kD;=�j:=��9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=��1=`�0=��/=��.=H�-=]�,=��+=��*=��)=@�(=��'=j�&=�%=��$=�#=h�"=oj!=4O =�0=�=�=��=Y�=c=5/=��=E�=+}=O:=��=�=�Z=�=��=�X=��	=M�=�3=��=�]=�=�x=�  =�	�<k�<��<|��<Z��<g��<��<O��<EX�<N%�<@��<���<Xi�<��<���<}�<`$�<��<^e�<J��<Q��<e'�<ֵ�<�@�<�Ȯ<M�<oϧ<�N�<�ˠ<�F�<F��<76�<���<��<���<}�<�u�<]�<D�z<��s<2nl<jOe<�1^<-W<��O<�H<{�A<��:<��3<��,<�%<��<#�<y�<k�	<��<Ż�;^ �;�S�;ȶ�;�*�;���;�F�;��;P��;r };V�b;��H;��.;�B;���:���:tĒ:S�A:~Y�9�1�c�ǹWD�ᵑ���������%�Ġ<�gS��Li�sG�$����A���⟻"d���Ǵ�%���0ɻ7ӻݻ���j��N"��%���r������^�?������C!���%�k�)���-��2��16��<:�7<>��0B��F���I�D�M���Q�FXU�IY�]�\�gb`���c��g�4k���n�t r�T�u�	y�jm|�(��n���i@��q脼�����0��<щ�To��2�������<���ґ��f��,���󉖼Y��[����3�������I��<ӟ��[��8㢼j��#𥼷u������`��}������E��掰����,������ߝ��"�������+������6���  �  �bN=4�M=�L=�L=�QK=�J=��I=0�H=�7H=�oG=�F=}�E=E=�GD=�{C=��B=^�A=-A=�@@=Vo?=��>=��==K�<=�<=dD;=�j:=��9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=��1=b�0=��/=��.=I�-=X�,=��+=��*=��)=F�(=��'=o�&=�%=��$= �#=p�"=tj!=2O =�0=�=��=�=R�=c=5/=��=M�=2}=Q:=��=�=�Z=�=��=�X=��	=F�=�3=��=�]=�=�x=�  =�	�<f�<��<}��<H��<k��<��<M��<LX�<?%�<L��<���<Yi�<��<���<	}�<i$�<��<Ne�<L��<F��<b'�<浵<�@�<�Ȯ<�M�<qϧ<�N�<�ˠ<�F�<I��<A6�<���<��<���<x�<�u�<J�<K�z<��s<Bnl<wOe<�1^<
W<��O<
�H<Y�A<��:<j�3<�,<��%<��<9�<v�<g�	<��<���;@ �;�S�;˶�;�*�;���;�F�;��;���;c };��b;&�H;��.;
C;~��:"��: Œ:��A:)W�9�D1���ǹgD�c���a����������%���<�pS�8Mi�eG�Q����A���⟻Wd��OǴ�@��y0ɻ�6ӻ�ݻ���$��$"��,���r������k�Z������C!�s�%�I�)���-��2��16��<:�N<>��0B�F���I�K�M���Q�AXU�kY�_�\�^b`���c��g�&k���n�� r�R�u�,y�am|�9��o���a@��脼썆��0��;щ�Go��%�������<���ґ��f��+�������\��K���4��x����I��;ӟ��[��.㢼j��!𥼮u������U���������C���������'������ٝ��"�������+�����7���  �  �bN=.�M=�L=�L=�QK=�J=��I=6�H=�7H=�oG=�F=y�E=E=�GD=�{C=��B=`�A='A=�@@=Ro?=��>=��==C�<=�<=bD;=�j:=��9=��8=$�7=��6=�6=�-5=�G4=�_3=�u2=��1=]�0=��/=��.=N�-=Z�,=��+=��*=��)=K�(=��'=p�&=�%=��$=�#=f�"=uj!=,O =�0=�= �=��=T�=c=-/=��=D�=.}=O:=��=�=�Z=�=�=�X=��	=G�=�3=��=�]=�=�x=�  =�	�<o�<��<���<D��<{��<��<H��<UX�<;%�<R��<���<_i�<��<���<	}�<[$�<��<Le�<V��<G��<e'�<⵵<�@�<�Ȯ<}M�<{ϧ<�N�<�ˠ<�F�<D��<F6�<���<��<���<�<�u�<M�<g�z<��s<Fnl<_Oe<�1^<W<��O<!�H<P�A<��:<R�3<�,<��%<��<8�<a�<��	<��<��;1 �;�S�;ٶ�;�*�;���;�F�;��;P��;` };m�b;��H;;�.;�B;���:���:8Œ:,�A:�U�9`�0���ǹ�D��������_��7���%���<��S�5Mi�G�@����A���⟻�d��#Ǵ�c��u0ɻ"7ӻݻ���u��"��D���r������X�S������C!�r�%�o�)���-��2��16��<:�`<>��0B�$F���I�:�M���Q�,XU�qY�>�\�pb`���c��g�-k���n�� r�9�u�5y�Cm|�;��u���X@���脼獆��0��5щ�So��2�������<���ґ��f��!�������Y��O���4��x����I��0ӟ��[��3㢼j��&𥼨u������C���������B������|��5������坶�"�������+������7���  �  �bN=6�M=�L=�L=�QK=�J=��I=8�H=�7H=�oG=�F=v�E=E=�GD=�{C=��B=`�A=&A=�@@=So?=��>=��==C�<=�<=gD;=�j:=��9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=1=\�0=��/=��.=H�-=Y�,=��+=��*=��)=E�(=��'=r�&=�%=��$= �#=g�"=uj!=3O =�0=�=��=�=V�=c=4/=��=E�=/}=P:=��= �=�Z=�=��=�X=��	=G�=�3=��=�]=�=�x=�  =�	�<n�<��<���<F��<i��<��<L��<DX�<A%�<Q��<���<`i�<��<���<}�<_$�<��<Se�<L��<G��<e'�<ܵ�<�@�<�Ȯ<zM�<ϧ<�N�<�ˠ<�F�<;��<?6�<���<��<���<|�<�u�<X�<O�z<��s<\nl<XOe<�1^<(W<|�O<�H<N�A<��:<r�3<
�,<ؗ%<��<<�<Y�<��	<��<��;j �;�S�;۶�;�*�;���;�F�;��;L��;� };��b;��H;K�.;�B;���:y��:2Ē:s�A:vX�9�U1���ǹ}D���������������%��<�%S� Mi�zG�D����A���⟻Od��RǴ�e��c0ɻ	7ӻݻ���m��"��'���r������h�K������C!�j�%�i�)���-��2��16��<:�Z<>��0B�F���I�U�M���Q�DXU�gY�K�\�ub`���c��g�3k���n�� r�I�u�0y�fm|�-��q���i@��}脼荆��0��4щ�Po��.��癩��<���ґ��f��+�������Y��U����3��z����I��,ӟ��[��0㢼�i��/𥼯u������N���������I��뎰����9������蝶�"�������+�����7���  �  �bN=4�M=�L=�L=�QK=�J=��I=4�H=�7H=�oG=�F=w�E=E=�GD=�{C=��B=]�A=(A=�@@=So?=��>=��==G�<=�<=hD;=�j:=��9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=��1=a�0=��/=��.=E�-=^�,=��+=��*=��)=D�(=��'=n�&=�%=��$=�#=o�"=pj!=1O =�0=�= �=��=V�=c=3/=��=L�=0}=O:=��=�=�Z=�=��=�X=��	=N�=�3=��=�]=�=�x=�  =�	�<g�<��<y��<W��<l��<
��<K��<KX�<G%�<I��<���<Xi�<��<���<}�<`$�<��<Qe�<S��<K��<c'�<ݵ�<�@�<�Ȯ<�M�<xϧ<�N�<�ˠ<�F�<J��<=6�<���<��<���<��<�u�<T�<F�z<��s<Gnl<tOe<�1^<W<x�O<�H<l�A<��:<i�3<�,<�%<��<6�<f�<y�	<��<��;D �;�S�;ζ�;�*�;���;�F�;��;Z��;b };��b;�H;�.;�B;K��:���:�Ē:B�A:�W�9+71�i�ǹ�D�m���?����������%���<�vS��Li��G�����A���⟻Wd��ZǴ�0���0ɻ�6ӻݻ���/��C"��/���r������[�N������C!���%�P�)���-��2��16��<:�C<>��0B�F���I�H�M���Q�QXU�`Y�b�\�cb`���c��g�,k���n�� r�Z�u�y�_m|�4��q���b@��w脼�����0��;щ�Ho��*�������<���ґ��f��$�������[��U���4������I��3ӟ��[��1㢼j�� 𥼱u������R���������L������+������ڝ��"�������+������6���  �  �bN=0�M=�L=�L=�QK=�J=��I=4�H=�7H=�oG=�F={�E=E=�GD=�{C=��B=`�A=)A=�@@=Po?=��>=��==H�<=�<=`D;=�j:=��9=��8= �7=��6=�6=�-5=�G4=�_3=�u2=��1=b�0=��/=��.=K�-=[�,=��+=��*=��)=I�(=��'=k�&=�%=��$=�#=g�"=tj!=/O =�0=�= �=��=Q�=c=1/=��=E�=.}=P:=��=�=�Z=�=��=�X=��	=H�=�3=��=�]=�=�x=�  =�	�<i�<��<���<F��<p��<��<I��<TX�<8%�<K��<���<]i�<��<���<}�<`$�<��<Ge�<Y��<C��<d'�<㵵<�@�<�Ȯ<|M�<uϧ<�N�<�ˠ<vF�<L��<C6�<���<��<���<�<�u�<P�<O�z<��s<5nl<sOe<�1^<W<��O<�H<K�A<��:<\�3<�,< �%<o�<:�<q�<w�	<��<��;E �;�S�;ն�;p*�;ʯ�;�F�;��;f��;� };Y�b;��H;*�.;�B;k��:���:fŒ:/�A:�V�9�
1��ǹ�D�����4������� �%���<�DS��Li�GG�3����A���⟻rd��2Ǵ�K���0ɻ�6ӻݻ���o��#"��8���r������T�^������C!�r�%�k�)���-��2��16��<:�X<>��0B�F���I�O�M���Q�:XU�^Y�W�\�_b`���c��g�,k���n�~ r�I�u�1y�Xm|�2��t���Y@���脼��0��7щ�Ro��3�������<���ґ��f��������Z��N���4��x����I��6ӟ��[��0㢼j��𥼫u������J���������A��򎰼���)������۝��"�������+�����7���  �  �bN=2�M=�L=�L=�QK=�J=��I=;�H=�7H=�oG=�F=u�E=E=�GD=�{C=��B=f�A=$A=�@@=Ro?=��>=��==@�<=�<=cD;=�j:=�9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=��1=_�0=��/=��.=G�-=Y�,=��+=��*=��)=I�(=��'=t�&=�%=��$=&�#=f�"=zj!=-O =�0=�=��=�=S�=c=//=��=D�=5}=N:=��=!�=�Z=�=~�=�X=��	=G�=�3=��=�]=�=�x=�  =�	�<n�<��<���<E��<m��<��<B��<NX�<:%�<U��<���<bi�<��<���<}�<W$�<��<Ie�<P��<@��<m'�<ݵ�<�@�<�Ȯ<yM�<�ϧ<�N�<�ˠ<�F�<B��<C6�<���<��<���<�<�u�<T�<N�z<��s<Nnl<fOe<�1^<#W<r�O<�H<P�A<��:<a�3<
�,<�%<��<>�<Q�<��	<��< ��;N �;�S�;��;v*�;���;�F�;��;>��;� };s�b;��H;v�.;^B;���:���:�Ē:��A:�V�9)'1�~�ǹ�D���������������%�ڠ<�8S�/Mi��G�F����A���⟻zd��2Ǵ�b��W0ɻ7ӻݻ���t���!��>���r������e�X������C!�Z�%�l�)���-��2��16��<:�_<>��0B�%F���I�S�M���Q�EXU�uY�P�\�ib`���c��g�.k���n�� r�H�u�3y�]m|�7��z���_@���脼㍆��0��1щ�Io��0��뤎��<���ґ��f��'������R��U���4��r����I��'ӟ��[��/㢼�i��(𥼬u������L���������M������1������᝶�"�������+�����7���  �  �bN=8�M=�L=�L=�QK=�J=��I=3�H=�7H=�oG=	�F=t�E=E=�GD=�{C=��B=^�A="A=�@@=Oo?=��>=��==G�<=�<=fD;=�j:=��9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=��1=_�0=��/=��.=G�-=`�,=��+=��*=��)=F�(=��'=n�&=�%=��$=�#=g�"=sj!=0O =�0=�=�=��=W�=c=1/=��=D�=0}=L:=��=�=�Z=�=��=�X=��	=P�=�3=��=�]=�=�x=�  =�	�<o�<��<���<Y��<l��<��<M��<OX�<D%�<L��<���<Ui�<��<���<}�<V$�<��<Te�<R��<J��<g'�<ص�<�@�<�Ȯ<�M�<uϧ<�N�<�ˠ<�F�<D��<?6�<���<��<���<��<�u�<_�<G�z<��s<9nl<kOe<�1^<4W<w�O<"�H<s�A<��:<y�3<�,<�%<��<8�<g�<s�	<��<л�;` �;�S�;޶�;�*�;���;�F�;��;0��;� };@�b;��H;��.;�B;���:f��:�Ē:��A:Y�9�c1���ǹ�D�y�����������%�Ӡ<�OS��Li��G�
����A���⟻Hd��LǴ�L���0ɻ�6ӻݻ���l��-"��4���r������U�I������C!�r�%�n�)���-��2��16��<:�P<>��0B�F���I�@�M���Q�EXU�UY�W�\�nb`���c��g�6k���n�� r�K�u�
y�`m|�*��o���_@��{脼퍆��0��?щ�No��5��󤎼�<���ґ��f��$�������W��Y����3������I��6ӟ��[��.㢼 j��&𥼯u������V�����}���M��㎰����.������ߝ��"�������+�������6���  �  �bN=8�M=�L=�L=�QK=�J=��I=,�H=�7H=�oG=
�F={�E=E=�GD=�{C=��B=]�A=-A=�@@=Ro?=��>=��==O�<=�<=fD;=�j:=~�9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=��1=g�0=��/=��.=D�-=Z�,=��+=��*=��)=@�(=��'=j�&=�%=��$=�#=p�"=rj!=6O =�0=�=��=�=T�=c=9/=��=K�=0}=O:=��=�=�Z=�=��=�X=��	=G�=�3=��=�]=�=�x=�  =�	�<a�<��<u��<H��<c��<��<F��<FX�<G%�<@��<���<Ri�<��<���<}�<k$�<��<Pe�<H��<D��<a'�<⵵<�@�<�Ȯ<�M�<iϧ<�N�<�ˠ<}F�<P��<36�<���<��<���<z�<�u�<Q�<<�z<ҍs<5nl<�Oe<�1^<W<��O<	�H<S�A<��:<z�3<�,< �%<��<,�<��<W�	< �<ۻ�;f �;�S�;ƶ�;�*�;z��;�F�;��;���;� };}�b;N�H;��.;MC;��:`��:�Ē:��A:�Y�9m�1���ǹ;D����������������%�V�<��S��Li��G�?����A���⟻Od��yǴ����0ɻ�6ӻ�ݻ���)��5"�����r������l�S������C!�w�%�R�)���-��2��16��<:�5<>��0B�F���I�\�M���Q�UXU�XY�j�\�Pb`���c���g�%k���n�{ r�a�u�,y�rm|�*��w���h@��v脼�����0��Aщ�Eo��+�������<���ґ��f��/������]��O����3��~����I��Bӟ��[��2㢼j��𥼻u������T���������I��򎰼���������Н��"�������+�����
7���  �  �bN=3�M=�L=�L=�QK= �J=��I=3�H=�7H=�oG=�F=v�E=E=�GD=�{C=��B=b�A=&A=�@@=Mo?=��>=��==D�<=�<=gD;=�j:=��9=��8=!�7=��6=�6=�-5=�G4=�_3=�u2=��1=]�0=��/=��.=L�-=]�,=��+=��*=��)=F�(=��'=n�&=�%=��$=!�#=g�"=qj!=,O =�0=�=�=��=V�=c=./=��=C�=0}=L:=��=�=�Z=�=��=�X=��	=J�=�3=��=�]=�=�x=�  =�	�<k�<��<���<K��<t��<��<I��<KX�<H%�<G��<���<Xi�<��<���<}�<[$�<��<Qe�<[��<J��<h'�<ܵ�<�@�<�Ȯ<M�<wϧ<�N�<�ˠ<�F�<H��<>6�<���<��<���<��<�u�<T�<N�z<��s<9nl<_Oe<�1^<W<��O<*�H<Y�A<��:<f�3<�,<�%<��<)�<^�<u�	<��<˻�; �;�S�;��;�*�;ϯ�;�F�;��;K��;8 };+�b;�H;�.;�B; ��:x��:�Ē:>�A:�W�9�0�0�ǹ�D����������A��%��<�>S��Li�;G�#����A���⟻dd��JǴ�2���0ɻ.7ӻ'ݻ���o��<"��C���r������Q�M������C!�~�%�s�)���-��2��16��<:�A<>��0B�F���I�F�M���Q�1XU�^Y�T�\�lb`���c��g�/k���n�� r�;�u�'y�Qm|�-��s���b@��v脼򍆼�0��<щ�Ko��9�������<���ґ��f���������V��V���4�������I��4ӟ��[��;㢼j��!𥼰u������F�����{���C������5������䝶�"�������+������7���  �  �bN=.�M="�L=�L=�QK=�J=��I=>�H=�7H=�oG=�F=y�E=E=�GD=�{C=~�B=a�A='A=�@@=Ro?=��>=��==C�<=�<=eD;=�j:=��9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=ɉ1=Z�0=��/=��.=F�-=X�,=��+=��*=��)=L�(=��'=v�&=�%=��$=&�#=b�"=j!=2O =�0=�=��=�=P�=c=3/=��=A�=4}=S:=��=#�=�Z=�=��=�X=��	=E�=�3=��=�]=�=�x=�  =�	�<t�<��<���<A��<o��<��<M��<JX�<>%�<W��<���<ii�<��<���<!}�<_$�<��<Ae�<S��<7��<b'�<䵵<�@�<�Ȯ<qM�<�ϧ<�N�<�ˠ<�F�<7��<N6�<���<��<���<��<�u�<T�<c�z<��s<tnl<WOe<�1^<"W<d�O<�H<F�A<��:<R�3<$�,<֗%<��<@�<\�<��	<��<��;� �;�S�;ڶ�;I*�;���;~F�;��;U��;};s�b;��H;��.;�B;��:=��:�Ē:y�A:�T�9�1���ǹ[D�6�����������2�%�.�<��S�5Mi��G�P����A���⟻|d��Ǵ�{��B0ɻ�6ӻ�ݻ��滕���!��*���r������g�f������C!�B�%�y�)���-��2��16��<:�c<>��0B�F���I�Q�M���Q�AXU�{Y�D�\�xb`���c��g�0k���n�� r�B�u�;y�Zm|�F��o���b@���脼⍆��0��*щ�Oo��3��ऎ��<���ґ��f��$������]��M����3��k����I��"ӟ��[��.㢼�i��2𥼠u������N���������U���~��;������蝶�"�������+�� ���7���  �  �bN=3�M=�L=�L=�QK= �J=��I=3�H=�7H=�oG=�F=v�E=E=�GD=�{C=��B=b�A=&A=�@@=Mo?=��>=��==D�<=�<=gD;=�j:=��9=��8=!�7=��6=�6=�-5=�G4=�_3=�u2=��1=]�0=��/=��.=L�-=]�,=��+=��*=��)=F�(=��'=n�&=�%=��$=!�#=g�"=qj!=,O =�0=�=�=��=V�=c=./=��=C�=0}=L:=��=�=�Z=�=��=�X=��	=J�=�3=��=�]=�=�x=�  =�	�<k�<��<���<K��<t��<��<I��<KX�<H%�<G��<���<Xi�<��<���<}�<[$�<��<Qe�<[��<J��<h'�<ܵ�<�@�<�Ȯ<M�<wϧ<�N�<�ˠ<�F�<H��<>6�<���<��<���<��<�u�<T�<N�z<��s<9nl<_Oe<�1^<W<��O<*�H<Y�A<��:<f�3<�,<�%<��<)�<^�<u�	<��<˻�; �;�S�;��;�*�;ϯ�;�F�;��;K��;8 };+�b;�H;�.;�B; ��:x��:�Ē:=�A:�W�9�0�0�ǹ�D����������A��%��<�>S��Li�;G�#����A���⟻dd��JǴ�2���0ɻ.7ӻ'ݻ���o��<"��C���r������Q�M������C!�~�%�s�)���-��2��16��<:�A<>��0B�F���I�F�M���Q�1XU�^Y�T�\�lb`���c��g�/k���n�� r�;�u�'y�Qm|�-��s���b@��v脼򍆼�0��<щ�Ko��9�������<���ґ��f���������V��V���4�������I��4ӟ��[��;㢼j��!𥼰u������F�����{���C������5������䝶�"�������+������7���  �  �bN=8�M=�L=�L=�QK=�J=��I=,�H=�7H=�oG=
�F={�E=E=�GD=�{C=��B=]�A=-A=�@@=Ro?=��>=��==O�<=�<=fD;=�j:=~�9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=��1=g�0=��/=��.=D�-=Z�,=��+=��*=��)=@�(=��'=j�&=�%=��$=�#=p�"=rj!=6O =�0=�=��=�=T�=c=9/=��=K�=0}=O:=��=�=�Z=�=��=�X=��	=G�=�3=��=�]=�=�x=�  =�	�<a�<��<u��<H��<c��<��<F��<FX�<G%�<@��<���<Ri�<��<���<}�<k$�<��<Pe�<H��<D��<a'�<⵵<�@�<�Ȯ<�M�<iϧ<�N�<�ˠ<}F�<P��<36�<���<��<���<z�<�u�<Q�<<�z<ҍs<5nl<�Oe<�1^<W<��O<	�H<S�A<��:<z�3<�,< �%<��<,�<��<W�	< �<ۻ�;f �;�S�;ƶ�;�*�;z��;�F�;��;���;� };}�b;N�H;��.;MC;��:`��:�Ē:��A:�Y�9x�1���ǹ;D����������������%�V�<��S��Li��G�?����A���⟻Od��yǴ����0ɻ�6ӻ�ݻ���)��5"�����r������l�S������C!�w�%�R�)���-��2��16��<:�5<>��0B�F���I�\�M���Q�UXU�XY�j�\�Pb`���c���g�%k���n�{ r�a�u�,y�rm|�*��w���h@��v脼�����0��Aщ�Eo��+�������<���ґ��f��/������]��O����3��~����I��Bӟ��[��2㢼j��𥼻u������T���������I��򎰼���������Н��"�������+�����
7���  �  �bN=8�M=�L=�L=�QK=�J=��I=3�H=�7H=�oG=	�F=t�E=E=�GD=�{C=��B=^�A="A=�@@=Oo?=��>=��==G�<=�<=fD;=�j:=��9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=��1=_�0=��/=��.=G�-=`�,=��+=��*=��)=F�(=��'=n�&=�%=��$=�#=g�"=sj!=0O =�0=�=�=��=W�=c=1/=��=D�=0}=L:=��=�=�Z=�=��=�X=��	=P�=�3=��=�]=�=�x=�  =�	�<o�<��<���<Y��<l��<��<M��<OX�<D%�<L��<���<Ui�<��<���<}�<V$�<��<Te�<R��<J��<g'�<ص�<�@�<�Ȯ<�M�<uϧ<�N�<�ˠ<�F�<D��<?6�<���<��<���<��<�u�<_�<G�z<��s<9nl<kOe<�1^<4W<w�O<"�H<s�A<��:<y�3<�,<�%<��<8�<g�<s�	<��<л�;` �;�S�;޶�;�*�;���;�F�;��;0��;� };@�b;��H;��.;�B;���:f��:�Ē:��A:Y�9�c1���ǹ�D�y�����������%�Ӡ<�OS��Li��G�
����A���⟻Hd��LǴ�L���0ɻ�6ӻݻ���l��-"��4���r������U�I������C!�r�%�n�)���-��2��16��<:�P<>��0B�F���I�@�M���Q�EXU�UY�W�\�nb`���c��g�6k���n�� r�K�u�
y�`m|�*��o���_@��{脼퍆��0��?щ�No��5��󤎼�<���ґ��f��$�������W��Y����3������I��6ӟ��[��.㢼 j��&𥼯u������V�����}���M��㎰����.������ߝ��"�������+�������6���  �  �bN=2�M=�L=�L=�QK=�J=��I=;�H=�7H=�oG=�F=u�E=E=�GD=�{C=��B=f�A=$A=�@@=Ro?=��>=��==@�<=�<=cD;=�j:=�9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=��1=_�0=��/=��.=G�-=Y�,=��+=��*=��)=I�(=��'=t�&=�%=��$=&�#=f�"=zj!=-O =�0=�=��=�=S�=c=//=��=D�=5}=N:=��=!�=�Z=�=~�=�X=��	=G�=�3=��=�]=�=�x=�  =�	�<n�<��<���<E��<m��<��<B��<NX�<:%�<U��<���<bi�<��<���<}�<W$�<��<Ie�<P��<@��<m'�<ݵ�<�@�<�Ȯ<yM�<�ϧ<�N�<�ˠ<�F�<B��<B6�<���<��<���<�<�u�<T�<N�z<��s<Nnl<fOe<�1^<#W<r�O<�H<P�A<��:<a�3<
�,<�%<��<>�<Q�<��	<��< ��;N �;�S�;��;v*�;���;�F�;��;>��;� };s�b;��H;v�.;^B;���:���:�Ē:��A:�V�9O'1��ǹ�D���������������%�ڠ<�8S�/Mi��G�F����A���⟻zd��2Ǵ�b��W0ɻ7ӻݻ���t���!��>���r������e�X������C!�Z�%�l�)���-��2��16��<:�_<>��0B�%F���I�S�M���Q�EXU�uY�P�\�ib`���c��g�.k���n�� r�H�u�3y�]m|�7��z���_@���脼㍆��0��1щ�Io��0��뤎��<���ґ��f��'������R��U���4��r����I��'ӟ��[��/㢼�i��(𥼬u������L���������M������1������᝶�"�������+�����7���  �  �bN=0�M=�L=�L=�QK=�J=��I=4�H=�7H=�oG=�F={�E=E=�GD=�{C=��B=`�A=)A=�@@=Po?=��>=��==H�<=�<=`D;=�j:=��9=��8= �7=��6=�6=�-5=�G4=�_3=�u2=��1=b�0=��/=��.=K�-=[�,=��+=��*=��)=I�(=��'=k�&=�%=��$=�#=g�"=tj!=/O =�0=�= �=��=Q�=c=1/=��=E�=.}=P:=��=�=�Z=�=��=�X=��	=H�=�3=��=�]=�=�x=�  =�	�<i�<��<���<F��<p��<��<I��<TX�<8%�<K��<���<]i�<��<���<}�<`$�<��<Ge�<Y��<C��<d'�<㵵<�@�<�Ȯ<|M�<uϧ<�N�<�ˠ<vF�<L��<C6�<���<��<���<�<�u�<P�<O�z<��s<5nl<sOe<�1^<W<��O<�H<L�A<��:<\�3<�,< �%<o�<:�<q�<w�	<��<��;E �;�S�;ն�;p*�;ʯ�;�F�;��;e��;� };Y�b;��H;*�.;�B;k��:���:eŒ:/�A:�V�9�
1��ǹ�D�����4������� �%���<�DS��Li�GG�3����A���⟻rd��2Ǵ�K���0ɻ�6ӻݻ���o��#"��8���r������U�^������C!�r�%�k�)���-��2��16��<:�X<>��0B�F���I�O�M���Q�:XU�^Y�W�\�_b`���c��g�,k���n�~ r�I�u�1y�Xm|�2��t���Y@���脼��0��7щ�Ro��3�������<���ґ��f��������Z��N���4��x����I��6ӟ��[��0㢼j��𥼫u������J���������A��򎰼���)������۝��"�������+�����7���  �  �bN=4�M=�L=�L=�QK=�J=��I=4�H=�7H=�oG=�F=w�E=E=�GD=�{C=��B=]�A=(A=�@@=So?=��>=��==G�<=�<=hD;=�j:=��9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=��1=a�0=��/=��.=E�-=^�,=��+=��*=��)=D�(=��'=n�&=�%=��$=�#=o�"=pj!=1O =�0=�= �=��=V�=c=3/=��=L�=0}=O:=��=�=�Z=�=��=�X=��	=N�=�3=��=�]=�=�x=�  =�	�<g�<��<y��<W��<l��<
��<K��<KX�<G%�<I��<���<Xi�<��<���<}�<`$�<��<Qe�<S��<K��<c'�<ݵ�<�@�<�Ȯ<�M�<xϧ<�N�<�ˠ<�F�<J��<=6�<���<��<���<��<�u�<T�<F�z<��s<Gnl<tOe<�1^<W<x�O<�H<l�A<��:<i�3<�,<�%<��<6�<f�<y�	<��<��;D �;�S�;ζ�;�*�;���;�F�;��;Z��;b };��b;�H;�.;�B;K��:���:�Ē:B�A:�W�9K71�k�ǹ�D�m���?����������%���<�vS��Li��G�����A���⟻Wd��ZǴ�0���0ɻ�6ӻݻ���/��C"��/���r������[�N������C!���%�P�)���-��2��16��<:�C<>��0B�F���I�H�M���Q�QXU�`Y�b�\�cb`���c��g�,k���n�� r�Z�u�y�_m|�4��q���b@��w脼�����0��;щ�Ho��*�������<���ґ��f��$�������[��U���4������I��3ӟ��[��1㢼j�� 𥼱u������R���������L������+������ڝ��"�������+������6���  �  �bN=6�M=�L=�L=�QK=�J=��I=8�H=�7H=�oG=�F=v�E=E=�GD=�{C=��B=`�A=&A=�@@=So?=��>=��==C�<=�<=gD;=�j:=��9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=1=\�0=��/=��.=H�-=Y�,=��+=��*=��)=E�(=��'=r�&=�%=��$= �#=g�"=uj!=3O =�0=�=��=�=V�=c=4/=��=E�=/}=P:=��= �=�Z=�=��=�X=��	=G�=�3=��=�]=�=�x=�  =�	�<n�<��<���<F��<i��<��<L��<DX�<A%�<Q��<���<`i�<��<���<}�<_$�<��<Se�<L��<G��<e'�<ܵ�<�@�<�Ȯ<zM�<ϧ<�N�<�ˠ<�F�<;��<?6�<���<��<���<|�<�u�<X�<O�z<��s<\nl<XOe<�1^<(W<|�O<�H<N�A<��:<r�3<
�,<ؗ%<��<<�<Y�<��	<��<��;j �;�S�;۶�;�*�;���;�F�;��;L��;� };��b;��H;K�.;�B;���:y��:2Ē:s�A:uX�9�U1���ǹ}D���������������%��<�%S� Mi�zG�D����A���⟻Od��RǴ�e��c0ɻ	7ӻݻ���m��"��'���r������h�K������C!�j�%�i�)���-��2��16��<:�Z<>��0B�F���I�U�M���Q�DXU�gY�K�\�ub`���c��g�3k���n�� r�I�u�0y�fm|�-��q���i@��}脼荆��0��4щ�Po��.��癩��<���ґ��f��+�������Y��U����3��z����I��,ӟ��[��0㢼�i��/𥼯u������N���������I��뎰����9������蝶�"�������+�����7���  �  �bN=.�M=�L=�L=�QK=�J=��I=6�H=�7H=�oG=�F=y�E=E=�GD=�{C=��B=`�A='A=�@@=Ro?=��>=��==C�<=�<=bD;=�j:=��9=��8=$�7=��6=�6=�-5=�G4=�_3=�u2=��1=]�0=��/=��.=N�-=Z�,=��+=��*=��)=K�(=��'=p�&=�%=��$=�#=f�"=uj!=,O =�0=�= �=��=T�=c=-/=��=D�=.}=O:=��=�=�Z=�=�=�X=��	=G�=�3=��=�]=�=�x=�  =�	�<o�<��<���<D��<{��<��<H��<UX�<;%�<R��<���<_i�<��<���<	}�<[$�<��<Le�<V��<G��<e'�<⵵<�@�<�Ȯ<}M�<{ϧ<�N�<�ˠ<�F�<D��<F6�<���<��<���<�<�u�<M�<g�z<��s<Fnl<_Oe<�1^<W<��O<!�H<P�A<��:<R�3<�,<��%<��<8�<a�<��	<��<��;1 �;�S�;ٶ�;�*�;���;�F�;��;P��;` };m�b;��H;;�.;�B;���:���:8Œ:+�A:�U�9u�0���ǹ�D��������`��7���%���<��S�5Mi�G�@����A���⟻�d��$Ǵ�c��u0ɻ"7ӻݻ���u��"��D���r������X�S������C!�r�%�o�)���-��2��16��<:�`<>��0B�%F���I�:�M���Q�,XU�qY�>�\�pb`���c��g�-k���n�� r�9�u�5y�Cm|�;��u���X@���脼獆��0��5щ�So��2�������<���ґ��f��!�������Y��O���4��x����I��0ӟ��[��3㢼j��&𥼨u������C���������B������|��5������坶�"�������+������7���  �  �bN=4�M=�L=�L=�QK=�J=��I=0�H=�7H=�oG=�F=}�E=E=�GD=�{C=��B=^�A=-A=�@@=Vo?=��>=��==K�<=�<=dD;=�j:=��9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=��1=b�0=��/=��.=I�-=X�,=��+=��*=��)=F�(=��'=o�&=�%=��$= �#=p�"=tj!=2O =�0=�=��=�=R�=c=5/=��=M�=2}=Q:=��=�=�Z=�=��=�X=��	=F�=�3=��=�]=�=�x=�  =�	�<f�<��<}��<H��<k��<��<M��<LX�<?%�<L��<���<Yi�<��<���<	}�<i$�<��<Ne�<L��<F��<b'�<浵<�@�<�Ȯ<�M�<qϧ<�N�<�ˠ<�F�<I��<A6�<���<��<���<x�<�u�<J�<K�z<��s<Bnl<wOe<�1^<
W<��O<
�H<Y�A<��:<j�3<�,<��%<��<9�<v�<g�	<��<���;@ �;�S�;˶�;�*�;���;�F�;��;���;c };��b;&�H;��.;
C;~��:"��: Œ:��A:(W�9�D1���ǹgD�c���a����������%���<�pS�8Mi�eG�Q����A���⟻Wd��OǴ�@��y0ɻ�6ӻ�ݻ���$��$"��,���r������k�Z������C!�s�%�I�)���-��2��16��<:�N<>��0B�F���I�K�M���Q�AXU�kY�_�\�^b`���c��g�&k���n�� r�R�u�,y�am|�9��o���a@��脼썆��0��;щ�Go��%�������<���ґ��f��+�������\��K���4��x����I��;ӟ��[��.㢼j��!𥼮u������U���������C���������'������ٝ��"�������+�����7���  �  �bN=<�M=�L=�L=�QK=��J=��I=1�H=�7H=�oG=	�F=t�E=E=�GD=�{C=��B=[�A=&A=�@@=Po?=��>=��==J�<=�<=kD;=�j:=��9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=��1=`�0=��/=��.=H�-=]�,=��+=��*=��)=@�(=��'=j�&=�%=��$=�#=h�"=oj!=4O =�0=�=�=��=Y�=c=5/=��=E�=+}=O:=��=�=�Z=�=��=�X=��	=M�=�3=��=�]=�=�x=�  =�	�<k�<��<|��<Z��<g��<��<O��<EX�<N%�<@��<���<Xi�<��<���<}�<`$�<��<^e�<J��<Q��<e'�<ֵ�<�@�<�Ȯ<M�<oϧ<�N�<�ˠ<�F�<F��<76�<���<��<���<}�<�u�<]�<D�z<��s<2nl<jOe<�1^<-W<��O<�H<{�A<��:<��3<��,<�%<��<#�<y�<k�	<��<Ż�;^ �;�S�;ȶ�;�*�;���;�F�;��;P��;r };V�b;��H;��.;�B;���:���:tĒ:S�A:}Y�9
�1�d�ǹWD�ᵑ���������%�Ġ<�gS��Li�sG�$����A���⟻"d���Ǵ�%���0ɻ7ӻݻ���j��O"��%���r������^�?������C!���%�k�)���-��2��16��<:�7<>��0B��F���I�D�M���Q�FXU�IY�]�\�gb`���c��g�4k���n�t r�T�u�
y�jm|�(��n���i@��q脼�����0��<щ�To��2�������<���ґ��f��,���󉖼Y��[����3�������I��<ӟ��[��8㢼j��#𥼷u������`��}������E��掰����,������ߝ��"�������+������6���  �  �bN=2�M=�L=�L=�QK=�J=��I=9�H=�7H=�oG=�F=x�E=E=�GD=�{C=��B=`�A=(A=�@@=Vo?=��>=��==E�<=�<=gD;=�j:=|�9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=É1=a�0=��/=��.=D�-=V�,=��+=��*=��)=D�(=��'=n�&=�%=��$="�#=i�"=xj!=2O =�0=�=��=�=T�=c=3/=��=G�=2}=Q:=��=�=�Z=�=~�=�X=��	=E�=�3=��=�]=�=�x=�  =�	�<j�<��<z��<G��<p��<��<>��<MX�<E%�<L��<���<di�<��<���<}�<a$�<��<Ie�<K��<@��<e'�<޵�<�@�<�Ȯ<�M�<�ϧ<�N�<�ˠ<�F�<J��<96�<���<��<���<v�<�u�<Q�<Y�z<��s<]nl<oOe<�1^<W<i�O<	�H<]�A<��:<`�3<��,<��%<��<4�<d�<��	<��<	��;j �;�S�;ض�;x*�;���;�F�;��;Z��;� };��b;��H;h�.;�B;g��:m��:�Ē:��A:\V�9�51�4�ǹ�D����:����������%���<�,S�)Mi��G�]����A���⟻{d��^Ǵ�'���0ɻ7ӻݻ���^��"��,���r������m�V������C!�`�%�b�)���-��2��16��<:�?<>��0B�'F���I�I�M���Q�PXU�rY�R�\�cb`���c���g�-k���n�� r�X�u�.y�Xm|�>�����`@��y脼퍆��0��0щ�Mo��(��癩��<���ґ��f��,������Y��S����3��s����I��*ӟ��[��1㢼j�� 𥼵u������R���������R��򎰼���,������ݝ��"�������+�����7���  �  `bN=��M=c�L=�L=�PK=�J=��I=��H=�6H=enG=}�F=��E=`E=�ED=�yC=q�B=4�A=�A=c>@=�l?=�>=��==Q�<=�<='A;=ig:=�9= �8=]�7=��6=�6=�)5=uC4=^[3=/q2=�1=V�0=��/=\�.=̼-=��,=	�+=��*=��)=��(=Q�'=ͻ&=I�%=��$=�#=){"=c!=�G =�(=�=�=�=<�=�Z=�&=>�=ֳ=�t=�1=�=��=R=��=ߩ=P=L�	=��=l+=D�=hU=��=}p=��<���<���<{��<g��<m��<��<֝�<rw�<�J�<�<���<F��<x]�<9�<���<lr�<4�<a��<\�<}��<猼<��<���<�9�<J®<�G�<�ɧ<�I�<JǠ<rB�<���<43�<��<��<됋<g�<u�<#�<��z<9�s<�pl<�Re<6^<�W<� P<��H<��A<��:<�3<5�,<�%<v�<H�<<�<N�	<��<P��;^%�;�z�;���;U�;�۳;�t�;� �;�ߋ;�f};"8c;z4I;/^/;j�;Cz�:���:���:�C:�Y�9Vs7�|�ù_�A�ۣ���ٿ�>��u�9`%�a<�R�R���h��~�P8������t������=}�������Ȼ��һ{�ܻ����L�S���/���O���
��x�#���i�\��$!�`m%���)���-��1�6�� :�!!>��B�9 F���I���M��Q��@U���X�n�\�GM`�X�c�8g��k���n��r��u���x�;]|�ȿ����19���ᄼM����*��0ˉ��i����������7���͑�;b����������{�������0��J����F��pП�Y���ࢼ�g��#�s��%����}��V��j���^
��B������ޕ�����띶�@"������,�������7���  �  XbN=��M=_�L=�L=�PK=�J=��I=�H=�6H=dnG=��F=��E=WE= FD=�yC=x�B=+�A=�A=e>@=�l?=�>=��==S�<=}<=/A;=cg:=�9=�8=V�7=��6=�6=�)5=sC4=`[3=5q2=�1=[�0=��/=]�.=ļ-=��,=�+=��*=��)=��(=W�'=̻&=H�%=��$=�#=1{"=c!=�G =�(=�= �=��==�=�Z=�&=@�=޳=�t=�1=�=��=%R=��=�=�O=F�	=��=e+=E�=fU=��=~p=��<���<���<y��<W��<p��<��<ܝ�<rw�<�J�<&�<���<J��<]�<G�<���<qr�<6�<P��<\�<���<���<��<s��<:�<I®<�G�<ʧ<�I�<BǠ<yB�<���<.3�<��<��<�<Z�<u�<&�<�z<F�s<�pl<�Re<6^<�W<� P<h�H<��A<��:<��3<(�,<�%<��<1�<J�<\�	<��<I��;�%�;�z�;���;FU�;ܳ;u�;z �;�ߋ;�f};E8c;�4I;j^/;��;}y�:���:���:��C:!]�9u9��ù1�A�����ٿ��t�-`%�<���R���h�b�~�s8����������[��^}������Ȼ��һZ�ܻ}�滷L�F�����P���
��x����i�~���#!�Ym%�۩)���-�p�1�6�� :�!>�B�' F���I���M��Q�AU���X�v�\�4M`�Q�c�$g��k��n��r��u���x�U]|�������<9���ᄼY����*��(ˉ��i����������7���͑�/b������酖���������0��K����F��hП�Y���ࢼ�g��#�s������}��Q��v���m
��?�����ؕ�����᝶�A"������$,�������7���  �  RbN=��M=]�L=�L=�PK=��J=��I=��H=�6H=]nG=��F=��E=WE=FD=�yC={�B=+�A=�A=d>@=�l?=�>=��==W�<=w<=6A;=_g:=�9=�8=Q�7=��6=�6=�)5=sC4=\[3=4q2=��1=^�0=��/=c�.=Ƽ-=��,=�+=��*=��)=��(=Z�'=ʻ&=G�%=��$=�#=.{"=c!=�G =�(=�=�=��=A�=�Z=�&=9�=ڳ=�t=�1=�=�=)R=��=�= P=J�	=Đ=e+=K�=aU=��=zp=��<���<���<���<V��<���<��<��<xw�<�J�<4�<���<Q��<t]�<=�<���<ir�<>�<N��<\�<x��<���<��<x��<	:�<:®<�G�<�ɧ<�I�<;Ǡ<}B�<���<&3�<!��<��<��<]�<
u�<0�<٭z<Q�s<�pl<�Re<�5^<�W<� P<k�H<��A<��:<��3<�,<�%<��< �<R�<D�	<��<��;�%�;�z�;���;\U�;�۳;u�;z �;	��;�f};�7c;�4I;^/;ε;�x�:v��:y��:��C:�_�9�/:��ù,�A�B����ٿ�g�t�t`%��<�ڃR�$�h�?�~�A8����������0���}��h����Ȼ��һm�ܻ ��L����
��P�|�
��x���}i�����#!�vm%��)���-�~�1�6�� :�� >�)B� F���I���M��Q�AU���X���\�1M`�c�c�+g��k��n��r��u�b�x�\]|�������E9���ᄼc���|*��3ˉ��i����������7���͑�+b������煖���������0��Z����F��uП�Y���ࢼ�g��%�s��
����}��@��s���e
��4�����ҕ�����ޝ��K"������,�������7���  �  VbN=��M=`�L=�L=�PK=��J=��I=��H=�6H=dnG=�F=��E=ZE=�ED=�yC=u�B=/�A=�A=b>@=�l?=�>=��==X�<={<=.A;=dg:=�9=�8=U�7=��6=�6=�)5=rC4=^[3=4q2=�1=^�0=��/=^�.=Ƽ-=��,=�+=��*=��)=��(=W�'=˻&=I�%=��$=�#=1{"=c!=�G =�(=�=�=��=?�=�Z=�&=>�=޳=�t=�1=�=��=%R=��=�=�O=H�	=��=f+=F�=dU=��=|p=��<���<���<��<W��<r��<��<ם�<sw�<�J�<&�<���<R��<v]�<C�<���<lr�<7�<X��<\�<{��<���<��<���<�9�<H®<�G�<�ɧ<�I�<?Ǡ<xB�<���<.3�<��<��<���<U�<
u�<$�<�z<Q�s<�pl<�Re<6^<�W<� P<]�H<��A<��:<��3<*�,<
�%<��<)�<T�<H�	<��<J��;l%�;�z�;���;1U�;�۳;�t�;� �;�ߋ;�f};N8c;�4I;^/;ݵ;9y�:���: ��:��C:�[�9�B9���ù]�A�ƣ��ڿ�5�t�H`%��<���R�x�h�E�~�y8����������]��]}�������Ȼ��һ_�ܻ��滵L�P���%��P���
��x� ���i�j���#!�am%�ک)���-�x�1��6�� :�!>�B�% F���I���M��Q�AU���X�}�\�.M`�Z�c�,g��k��n��r��u���x�Q]|�ǿ����;9���ᄼ[���{*��1ˉ��i����������7���͑�4b������񅖼��������0��L����F��qП�Y���ࢼ�g��%�s������}��M��{���e
��@�����ҕ���������F"������,��Ʊ���7���  �  _bN=��M=a�L=�L=�PK=�J=��I=��H=�6H=fnG=��F=��E=XE=�ED=�yC=s�B=/�A=�A=e>@=�l?=�>=��==S�<=�<=-A;=eg:=�9=�8=^�7=��6=�6=�)5=sC4=_[3=2q2=�1=W�0=��/=[�.=ʼ-=��,=�+=��*=��)=��(=S�'=ϻ&=G�%=��$=�#=){"=c!=�G =�(=�=!�=��=:�=�Z=�&=C�=׳=�t=�1=�=��=!R=��=�=P=K�	=��=k+=C�=hU=��=|p=��<���<���<w��<d��<n��<���<ٝ�<qw�<�J�<!�<���<G��<y]�<=�<���<rr�<.�<X��<	\�<���<�<��<z��<�9�<O®<�G�<�ɧ<�I�<BǠ<{B�<���<33�<
��<��<�<\�<	u�<!�<��z<3�s<�pl<�Re<6^<~W<� P<t�H<��A<��:<��3</�,<�%<��<5�<I�<S�	<��<Y��;o%�;�z�;���;)U�;:ܳ;�t�;� �;�ߋ;�f};,8c;�4I;;^/;��;�y�:c��:2��:��C:J[�9%7���ù��A�1����ٿ����t�F`%�P<�M�R���h��~�z8������x���y��;}��������Ȼ��һf�ܻ����L�(���,��P���
��x����i�i���#!�Pm%���)���-�w�1�6�� :�!>� B�5 F���I���M��Q��@U���X�k�\�BM`�Y�c�0g��k��n��r��u���x�6]|�Ŀ����79���ᄼQ����*��.ˉ��i����������7���͑�9b���������������0��E����F��mП�Y���ࢼ�g��)�s��!����}��P��u���e
��C������╳����띶�="�����,�������7���  �  UbN=��M=a�L=�L=�PK=��J=��I=�H=�6H=enG=��F=��E=\E=�ED=�yC=r�B=1�A=�A=h>@=�l?=�>=��==T�<=|<=2A;=`g:=�9=�8=S�7=��6=�6=�)5=uC4=[[3=1q2=�1=X�0=��/=^�.=ȼ-=��,=�+=��*=��)=��(=U�'=λ&=H�%=��$=
�#=,{"=c!=�G =�(=�=�=�=<�=�Z=�&=@�=ٳ=�t=�1=�=��=#R=��=�=�O=F�	=��=h+=F�=fU=��=}p=��<���<���<���<_��<o��<��<ܝ�<vw�<�J�<*�<���<L��<|]�<A�<���<tr�<8�<Z��<	\�<{��<팼<��<|��<:�<L®<�G�<ʧ<�I�<@Ǡ<�B�<���<03�<��<��<<_�<	u�<*�<�z<;�s<�pl<�Re<6^<�W<� P<t�H<��A<��:<��3<.�,<��%<��<,�<D�<\�	<��<P��;�%�;�z�;���;U�;�۳;�t�;� �;�ߋ;%g};8c;�4I;Y^/;��;\y�:���:���:@�C:�\�9��9�>�ùa�A������ٿ�����t�1`%�A<���R�x�h�!�~�e8����������_��c}��������Ȼ��һb�ܻ����L�A�����P���
��x�$���i�k���#!�Xm%��)���-�s�1�6�� :�
!>�B�) F���I���M��Q�AU���X�w�\�CM`�X�c�1g�k��n��r���u���x�\]|�������A9���ᄼY����*��+ˉ��i����������7���͑�9b������􅖼��������0��H����F��iП�Y���ࢼ�g��)�s������}��S��r���f
��;�����ݕ�����靶�E"������,�������7���  �  VbN=��M=^�L=�L=�PK=��J=��I=��H=�6H=bnG=��F=��E=[E=�ED=�yC=w�B=/�A=�A=c>@=�l?=�>=��==Y�<=y<=2A;=ag:=�9=�8=T�7=��6=�6=�)5=sC4=_[3=4q2=�1=_�0=��/=`�.=ļ-=��,=�+=��*=��)=��(=Y�'=ɻ&=J�%=��$=�#=2{"=c!=�G =�(=�=�=��=A�=�Z=�&=<�=޳=�t=�1=�=��='R=��=�=�O=G�	==d+=H�=cU=��=|p=��<���<���<~��<T��<~��<��<ܝ�<ww�<�J�<.�<���<W��<s]�<C�<���<kr�<5�<V��<\�<���<�<��<z��<�9�<C®<�G�<�ɧ<�I�<CǠ<xB�<���<)3�<��<��<���<[�<u�<'�<�z<O�s<�pl<�Re<6^<�W<� P<f�H<��A<��:<��3<$�,<�%<��<,�<U�<E�	<��<7��;s%�;�z�;���;;U�;�۳;�t�;� �;�ߋ;�f};,8c;�4I;^/;�;�x�:��:���:�C:�\�9�u9�h�ù��A�꣐��ٿ�	���t�S`%��<���R�_�h�j�~�R8����������@��x}��q���#�Ȼ��һg�ܻ��滰L�d�����P��
��x���~i�t���#!�hm%�ة)���-�~�1��6�� :�� >�B� F���I���M��Q�AU���X��\�&M`�[�c�.g��k��n��r��u�i�x�V]|�������B9���ᄼa���v*��4ˉ��i����������7���͑�.b������텖���������0��Q����F��rП�
Y���ࢼ�g��$�s������}��J��u���m
��=�����ӕ���������D"������#,��±���7���  �  \bN=��M=_�L=�L=�PK=�J=��I=��H=�6H=fnG=��F=��E=YE=�ED=�yC=q�B=1�A=�A=f>@=�l?=�>=��==V�<=|<=0A;=eg:=�9=�8=X�7=��6=�6=�)5=tC4=_[3=1q2=ބ1=Z�0=��/=`�.=ȼ-=��,=�+=��*=��)=��(=V�'=ʻ&=I�%=��$=�#=+{"=c!=�G =�(=�=�=��=:�=�Z=�&=A�=س=�t=�1=�=��=#R=��=�=P=I�	=��=h+=H�=eU=��=yp=��<���<���<���<\��<q��<��<ܝ�<sw�<�J�<'�<���<O��<s]�<>�<���<tr�<4�<[��<\�<���<팼<��<���<:�<K®<�G�<�ɧ<�I�<EǠ<wB�<���<.3�<��<��<�<Z�<u�<+�<�z<@�s<�pl<�Re<6^<�W<� P<n�H<��A<��:<��3<(�,<�%<��<4�<Q�<C�	<��<X��;�%�;�z�;���;U�; ܳ;�t�;� �;�ߋ;g};88c;�4I;�]/;õ;ky�:���:A��:��C:0\�9r8�͎ùa�A������ٿ����t��`%�)<���R�W�h�%�~�g8���������h��X}�������Ȼ��һh�ܻ����L�;�����P���
��x����i�j���#!�Um%��)���-�z�1�6�� :�
!>�B�, F���I���M��Q�AU���X�x�\�;M`�h�c�6g��k��n��r� �u���x�H]|�������89���ᄼZ���~*��4ˉ��i����������7���͑�;b������󅖼��������0��I����F��tП�Y���ࢼ�g��#�s������}��Q��v���c
��9�����ە�����睶�@"������,�������7���  �  YbN=��M=b�L=�L=�PK=�J=��I=�H=�6H=fnG=��F=��E=]E=�ED=�yC=o�B=4�A=�A=g>@=�l?=�>=��==R�<=<=/A;=cg:=�9=�8=W�7=��6=�6=�)5=sC4=Z[3=4q2=�1=Y�0=��/=[�.=ȼ-=��,=�+=��*=��)=��(=R�'=л&=F�%=��$=�#=*{"=c!=�G =�(=�=�=��=;�=�Z=�&=D�=ֳ=�t=�1=�=��=!R=��=ߩ= P=F�	=��=i+=D�=fU=��=�p=��<���<���<w��<c��<k��<��<ܝ�<rw�<�J�<#�<���<G��<]�<D�<���<vr�<-�<a��<\�<���<<��<z��<�9�<P®<�G�<ʧ<�I�<BǠ<B�<���<53�<��<��<쐋<^�<u�<#�<�z<C�s<�pl<�Re<�5^<�W<� P<s�H<��A<��:<��3<3�,<��%<��<2�<?�<j�	<��<]��;{%�;�z�;���;U�;ܳ;�t�;� �;�ߋ;g};8c;�4I;w^/;��;�y�:���:��:��C:�\�9�8���ù��A�:����ٿ���t��_%�+<���R���h�%�~�k8����������|��8}��������Ȼ��һm�ܻu���L�'���.��P���
��x����i�a��$!�Jm%���)���-�u�1�6�� :�!>� B�5 F���I���M��Q� AU���X�v�\�BM`�G�c�$g�k��n��r��u���x�O]|�������89���ᄼR����*��(ˉ��i����������7���͑�?b������򅖼��������0��D����F��_П�Y���ࢼ�g��-�s������}��U��s���j
��B�����ڕ�����坶�I"�� ���",�������7���  �  VbN=��M=_�L=�L=�PK= �J=��I=��H=�6H=`nG=��F=��E=YE=�ED=�yC=w�B=/�A=�A=g>@=�l?=�>=��==V�<={<=1A;=ag:=�9=�8=U�7=��6=�6=�)5=vC4=^[3=2q2=ބ1=\�0=��/=`�.=ļ-=��,=�+=��*=��)=��(=U�'=̻&=H�%=��$=�#=,{"=c!=�G =�(=�=�=��=?�=�Z=�&=>�=س=�t=�1=�=��=$R=��=�=�O=G�	==e+=G�=eU=��=yp=��<���<���<z��<Y��<}��<��<ޝ�<tw�<�J�<*�<���<O��<r]�<C�<���<pr�<3�<X��<\�<���<�<��<y��<:�<B®<�G�<�ɧ<�I�<BǠ<B�<���<,3�<��<��<���<`�< u�<,�<�z<K�s<�pl<�Re<6^<�W<� P<p�H<��A<��:<��3<%�,<��%<��</�<M�<I�	<��<*��;�%�;�z�;���;<U�;ܳ;�t�;� �;�ߋ;g};�7c;�4I;	^/;��;Py�:���:���:��C:�]�9�S9��ù��A�����ٿ�4���t��`%��<���R�`�h�a�~�F8����������S��a}�������Ȼ��һz�ܻ����L�Y�����P���
��x����i�q���#!�am%��)���-���1�6�� :�!>�B�# F���I���M��Q�AU���X�w�\�/M`�f�c�4g��k���n��r��u�k�x�T]|�������?9���ᄼZ���}*��5ˉ��i����������7���͑�0b������텖���������0��Q����F��pП�Y���ࢼ�g��,�s������}��H��q���n
��8�����Օ�����❶�E"������$,�������7���  �  VbN=��M=\�L=�L=�PK=��J=��I=��H=�6H=cnG=��F=��E=WE= FD=�yC=w�B=+�A=�A=f>@=�l?=�>=��==]�<=w<=2A;=bg:=�9=�8=R�7=��6=�6=�)5=qC4=][3=6q2=݄1=`�0=��/=d�.=¼-=��,=�+=��*=��)=��(=\�'=ǻ&=K�%=��$=�#=3{"=c!=�G =�(=�=�=��=>�=�Z=�&=>�=�=�t=�1=�=}�=*R=��=�=�O=D�	=��=a+=L�=_U=��=yp=��<���<���<���<L��<v��<߽�<۝�<qw�<�J�<0�<���<Z��<q]�<K�<���<qr�<>�<O��<\�<��<���<��<{��<	:�<F®<�G�<�ɧ<�I�<?Ǡ<vB�<Ļ�<&3�<��<��<�<S�<u�</�<ڭz<c�s<�pl<Se<�5^<�W<� P<T�H<��A<��:<��3<�,<�%<��<%�<k�<6�	<��<A��;�%�;�z�;���;CU�;�۳;�t�;z �;��;g};C8c;/5I;�]/;*�;�x�:��:뻓:3�C:�\�9d�9���ù��A�@���&ڿ�F�t��`%��<��R��h���~�l8����������X���}��]���3�Ȼ��һI�ܻ��滢L�[�����P���
��x����i�|���#!�cm%�ѩ)���-�r�1��6�� :�� >�#B�& F���I�ŴM��Q�"AU���X���\�&M`�f�c�&g��k��n��r�"�u�w�x�`]|�������@9���ᄼf���r*��6ˉ��i����������7���͑�0b������셖���������0��N����F��yП��X���ࢼ�g���s������}��N��~���h
��5�����ɕ�����ם��K"������,��˱���7���  �  \bN=��M=a�L=�L=�PK= �J=��I=��H=�6H=cnG=�F=��E=\E=�ED=�yC=t�B=0�A=�A=c>@=�l?=�>=��==W�<=|<=2A;=ag:=�9=�8=Z�7=��6=�6=�)5=oC4=[[3=6q2=�1=]�0=��/=`�.=Ǽ-=��,=
�+=��*=��)=��(=U�'=̻&=H�%=��$=�#=+{"=c!=�G =�(=�= �=��=>�=�Z=�&==�=س=�t=�1=�=��=$R=��=�=P=L�	==g+=H�=aU=��=~p=��<���<���<���<[��<{��<��<ޝ�<uw�<�J�<,�<���<P��<v]�<>�<���<lr�<1�<Z��<\�<���<���<��<z��<�9�<F®<�G�<�ɧ<�I�<@Ǡ<}B�<���<13�<��<��<���<_�<u�<'�<حz<U�s<�pl<�Re<�5^<�W<� P<n�H<��A<��:<��3<.�,< �%<��<.�<Q�<O�	<��<?��;m%�;�z�;���;;U�;ܳ;�t�;� �;�ߋ;�f};8c;�4I;^/;ʵ;^y�:��:���:��C:�\�9�"8���ù��A�����|ڿ���t�&`%��<�׃R�]�h�/�~�K8������t���n��^}������
�Ȼ��һi�ܻ����L�Z���(��P���
��x����i�k���#!�em%��)���-�|�1�6�� :�!>�B�, F���I���M��Q�AU���X���\�4M`�Q�c�#g��k��n��r��u�o�x�>]|�������=9���ᄼZ���}*��1ˉ��i����������7���͑�7b������ꅖ��������0��N����F��nП�
Y���ࢼ�g��)�s������}��K��r���g
��=�����Е�����ݝ��K"�����,�������7���  �  XbN=��M=g�L=�L=�PK=�J=��I=�H=�6H=jnG=��F=��E=\E=�ED=�yC=q�B=3�A=�A=k>@=�l?=�>=��==P�<=<=0A;=_g:=�9=�8=U�7=��6=�6=�)5=wC4=a[3=.q2=߄1=Y�0=��/=]�.=ż-=��,=�+=��*=��)=��(=M�'=һ&=F�%=��$=�#=*{"=c!=�G =�(=�=�=��=9�=�Z=�&=E�=ٳ=�t=�1=�=��=R=��=�=�O=E�	=��=e+=C�=iU=��=yp=
��<���<���<u��<X��<k��<��<՝�<ww�<�J�<"�<���<C��<]�<C�<���<{r�<-�<a��<\�<���<錼<��<~��<:�<S®<�G�<ʧ<�I�<FǠ<�B�<���<>3�<	��<��<ꐋ<]�< u�<-�<��z<:�s<�pl<�Re<6^<�W<� P<p�H<��A<��:<��3<E�,<�%<��<7�<4�<p�	<��<u��;�%�;�z�;���;U�;ܳ;�t�;� �;�ߋ;Tg};�8c;�4I;�^/;b�;�y�:���:���:��C:�Z�9|39�Y�ù��A�z���kٿ����u��`%�8<�P�R���h�X�~�w8����������x��-}��������Ȼ��һt�ܻu���L����&���O���
��x����i�c���#!�Dm%��)���-�v�1�6�� :�$!>�B�. F���I�´M��Q�AU���X�g�\�>M`�f�c�=g��k���n��r��u���x�R]|�ʿ����>9���ᄼR����*��(ˉ��i����������7���͑�?b������������������0��A����F��`П�Y���ࢼ�g��8�s��#����}��X��t���n
��8������ޕ�����읶�:"������&,�������7���  �  \bN=��M=a�L=�L=�PK= �J=��I=��H=�6H=cnG=�F=��E=\E=�ED=�yC=t�B=0�A=�A=c>@=�l?=�>=��==W�<=|<=2A;=ag:=�9=�8=Z�7=��6=�6=�)5=oC4=[[3=6q2=�1=]�0=��/=`�.=Ǽ-=��,=
�+=��*=��)=��(=U�'=̻&=H�%=��$=�#=+{"=c!=�G =�(=�= �=��=>�=�Z=�&==�=س=�t=�1=�=��=$R=��=�=P=L�	==g+=H�=aU=��=~p=��<���<���<���<[��<{��<��<ޝ�<uw�<�J�<,�<���<P��<v]�<>�<���<lr�<1�<Z��<\�<���<���<��<z��<�9�<F®<�G�<�ɧ<�I�<@Ǡ<}B�<���<13�<��<��<���<_�<u�<'�<حz<U�s<�pl<�Re<�5^<�W<� P<n�H<��A<��:<��3<.�,< �%<��<.�<Q�<O�	<��<?��;m%�;�z�;���;;U�;ܳ;�t�;� �;�ߋ;�f};8c;�4I;^/;ʵ;^y�:��:���:��C:�\�9�"8���ù��A�����|ڿ���t�&`%��<�׃R�]�h�/�~�K8������t���n��^}������
�Ȼ��һi�ܻ����L�Z���(��P���
��x����i�k���#!�em%��)���-�|�1�6�� :�!>�B�, F���I���M��Q�AU���X���\�4M`�Q�c�#g��k��n��r��u�o�x�>]|�������=9���ᄼZ���}*��1ˉ��i����������7���͑�7b������ꅖ��������0��N����F��nП�
Y���ࢼ�g��)�s������}��K��r���g
��=�����Е�����ݝ��K"�����,�������7���  �  VbN=��M=\�L=�L=�PK=��J=��I=��H=�6H=cnG=��F=��E=WE= FD=�yC=w�B=+�A=�A=f>@=�l?=�>=��==]�<=w<=2A;=bg:=�9=�8=R�7=��6=�6=�)5=qC4=][3=6q2=݄1=`�0=��/=d�.=¼-=��,=�+=��*=��)=��(=\�'=ǻ&=K�%=��$=�#=3{"=c!=�G =�(=�=�=��=>�=�Z=�&=>�=�=�t=�1=�=}�=*R=��=�=�O=D�	=��=a+=L�=_U=��=yp=��<���<���<���<L��<v��<߽�<۝�<qw�<�J�<0�<���<Z��<q]�<K�<���<qr�<>�<O��<\�<��<���<��<{��<	:�<F®<�G�<�ɧ<�I�<?Ǡ<vB�<Ļ�<&3�<��<��<�<S�<u�</�<ڭz<c�s<�pl<Se<�5^<�W<� P<T�H<��A<��:<��3<�,<�%<��<%�<k�<6�	<��<A��;�%�;�z�;���;CU�;�۳;�t�;z �;��;g};C8c;/5I;�]/;*�;�x�:��:뻓:3�C:�\�9��9���ù��A�@���&ڿ�F�t��`%��<��R��h���~�l8����������X���}��]���3�Ȼ��һI�ܻ��滢L�[�����P���
��x����i�|���#!�cm%�ѩ)���-�r�1��6�� :�� >�#B�& F���I�ŴM��Q�"AU���X���\�&M`�f�c�&g��k��n��r�"�u�w�x�`]|�������@9���ᄼf���r*��6ˉ��i����������7���͑�0b������셖���������0��N����F��yП��X���ࢼ�g���s������}��N��~���h
��5�����ɕ�����ם��K"������,��˱���7���  �  VbN=��M=_�L=�L=�PK= �J=��I=��H=�6H=`nG=��F=��E=YE=�ED=�yC=w�B=/�A=�A=g>@=�l?=�>=��==V�<={<=1A;=ag:=�9=�8=U�7=��6=�6=�)5=vC4=^[3=2q2=ބ1=\�0=��/=`�.=ļ-=��,=�+=��*=��)=��(=U�'=̻&=H�%=��$=�#=,{"=c!=�G =�(=�=�=��=?�=�Z=�&=>�=س=�t=�1=�=��=$R=��=�=�O=G�	==e+=G�=eU=��=yp=��<���<���<z��<Y��<}��<��<ޝ�<tw�<�J�<*�<���<O��<r]�<C�<���<pr�<3�<X��<\�<���<�<��<y��<:�<B®<�G�<�ɧ<�I�<BǠ<B�<���<,3�<��<��<���<`�< u�<,�<�z<K�s<�pl<�Re<6^<�W<� P<p�H<��A<��:<��3<%�,<��%<��</�<M�<I�	<��<*��;�%�;�z�;���;<U�;ܳ;�t�;� �;�ߋ;g};�7c;�4I;	^/;��;Py�:���:���:��C:�]�9.T9��ù��A�����ٿ�4���t��`%��<���R�`�h�a�~�F8����������S��a}�������Ȼ��һz�ܻ����L�Y�����P���
��x����i�q���#!�am%��)���-���1�6�� :�!>�B�# F���I���M��Q�AU���X�w�\�/M`�f�c�4g��k���n��r��u�k�x�T]|�������?9���ᄼZ���}*��5ˉ��i����������7���͑�0b������텖���������0��Q����F��pП�Y���ࢼ�g��,�s������}��H��q���n
��8�����Օ�����❶�E"������$,�������7���  �  YbN=��M=b�L=�L=�PK=�J=��I=�H=�6H=fnG=��F=��E=]E=�ED=�yC=o�B=4�A=�A=g>@=�l?=�>=��==R�<=<=/A;=cg:=�9=�8=W�7=��6=�6=�)5=sC4=Z[3=4q2=�1=Y�0=��/=[�.=ȼ-=��,=�+=��*=��)=��(=R�'=л&=F�%=��$=�#=*{"=c!=�G =�(=�=�=��=;�=�Z=�&=D�=ֳ=�t=�1=�=��=!R=��=ߩ= P=F�	=��=i+=D�=fU=��=�p=��<���<���<w��<c��<k��<��<ܝ�<rw�<�J�<#�<���<G��<]�<D�<���<vr�<-�<a��<\�<���<<��<z��<�9�<P®<�G�<ʧ<�I�<BǠ<B�<���<53�<��<��<쐋<^�<u�<#�<�z<C�s<�pl<�Re<�5^<�W<� P<s�H<��A<��:<��3<3�,<��%<��<2�<?�<j�	<��<]��;{%�;�z�;���;U�;ܳ;�t�;� �;�ߋ;g};8c;�4I;w^/;��;�y�:���:��:��C:�\�9`�8���ù��A�:����ٿ���t��_%�+<���R���h�%�~�k8����������|��8}��������Ȼ��һm�ܻu���L�'���.��P���
��x����i�a��$!�Jm%���)���-�u�1�6�� :�!>� B�5 F���I���M��Q� AU���X�v�\�BM`�G�c�$g�k��n��r��u���x�O]|�������89���ᄼR����*��(ˉ��i����������7���͑�?b������򅖼��������0��D����F��_П�Y���ࢼ�g��-�s������}��U��s���j
��B�����ڕ�����坶�I"�� ���",�������7���  �  \bN=��M=_�L=�L=�PK=�J=��I=��H=�6H=fnG=��F=��E=YE=�ED=�yC=q�B=1�A=�A=f>@=�l?=�>=��==V�<=|<=0A;=eg:=�9=�8=X�7=��6=�6=�)5=tC4=_[3=1q2=ބ1=Z�0=��/=`�.=ȼ-=��,=�+=��*=��)=��(=V�'=ʻ&=I�%=��$=�#=+{"=c!=�G =�(=�=�=��=:�=�Z=�&=A�=س=�t=�1=�=��=#R=��=�=P=I�	=��=h+=H�=eU=��=yp=��<���<���<���<\��<q��<��<ܝ�<sw�<�J�<'�<���<O��<s]�<>�<���<tr�<4�<[��<\�<���<팼<��<���<:�<K®<�G�<�ɧ<�I�<EǠ<wB�<���<.3�<��<��<�<Z�<u�<+�<�z<@�s<�pl<�Re<6^<�W<� P<n�H<��A<��:<��3<(�,<�%<��<4�<Q�<C�	<��<X��;�%�;�z�;���;U�; ܳ;�t�;� �;�ߋ;g};88c;�4I;�]/;µ;ky�:���:A��:��C:/\�9pr8�Ύùb�A������ٿ����t��`%�)<���R�W�h�%�~�g8���������h��X}�������Ȼ��һh�ܻ����L�;�����P���
��x����i�j���#!�Um%��)���-�z�1�6�� :�
!>�B�, F���I���M��Q�AU���X�x�\�;M`�h�c�6g��k��n��r� �u���x�H]|�������89���ᄼZ���}*��4ˉ��i����������7���͑�;b������󅖼��������0��I����F��tП�Y���ࢼ�g��#�s������}��Q��v���c
��9�����ە�����睶�@"������,�������7���  �  VbN=��M=^�L=�L=�PK=��J=��I=��H=�6H=bnG=��F=��E=[E=�ED=�yC=w�B=/�A=�A=c>@=�l?=�>=��==Y�<=y<=2A;=ag:=�9=�8=T�7=��6=�6=�)5=sC4=_[3=4q2=�1=_�0=��/=`�.=ļ-=��,=�+=��*=��)=��(=Y�'=ɻ&=J�%=��$=�#=2{"=c!=�G =�(=�=�=��=A�=�Z=�&=<�=޳=�t=�1=�=��='R=��=�=�O=G�	==d+=H�=cU=��=|p=��<���<���<~��<T��<~��<��<ܝ�<ww�<�J�<.�<���<W��<s]�<C�<���<kr�<5�<V��<\�<���<�<��<z��<�9�<C®<�G�<�ɧ<�I�<CǠ<xB�<���<)3�<��<��<���<[�<u�<'�<�z<O�s<�pl<�Re<6^<�W<� P<f�H<��A<��:<��3<$�,<�%<��<,�<U�<E�	<��<7��;s%�;�z�;���;;U�;�۳;�t�;� �;�ߋ;�f};,8c;�4I;^/;�;�x�:��:���:�C:�\�9�v9�i�ù��A�꣐��ٿ�	���t�T`%��<���R�`�h�j�~�R8����������@��x}��q���#�Ȼ��һg�ܻ��滰L�d�����P��
��x���~i�t���#!�hm%�ة)���-�~�1��6�� :�� >�B� F���I���M��Q�AU���X��\�&M`�[�c�.g��k��n��r��u�i�x�V]|�������B9���ᄼa���v*��4ˉ��i����������7���͑�.b������텖���������0��Q����F��rП�
Y���ࢼ�g��$�s������}��J��u���m
��=�����ӕ���������D"������#,��±���7���  �  UbN=��M=a�L=�L=�PK=��J=��I=�H=�6H=enG=��F=��E=\E=�ED=�yC=r�B=1�A=�A=h>@=�l?=�>=��==T�<=|<=2A;=`g:=�9=�8=S�7=��6=�6=�)5=uC4=[[3=1q2=�1=X�0=��/=^�.=ȼ-=��,=�+=��*=��)=��(=U�'=λ&=H�%=��$=
�#=,{"=c!=�G =�(=�=�=�=<�=�Z=�&=@�=ٳ=�t=�1=�=��=#R=��=�=�O=F�	=��=h+=F�=fU=��=}p=��<���<���<���<_��<o��<��<ܝ�<vw�<�J�<*�<���<L��<|]�<A�<���<tr�<8�<Z��<	\�<{��<팼<��<|��<:�<L®<�G�<ʧ<�I�<@Ǡ<�B�<���<03�<��<��<<_�<	u�<*�<�z<;�s<�pl<�Re<6^<�W<� P<t�H<��A<��:<��3<.�,<��%<��<,�<D�<\�	<��<P��;�%�;�z�;���;U�;�۳;�t�;� �;�ߋ;%g};8c;�4I;Y^/;��;\y�:���:���:?�C:�\�9�9�?�ùa�A������ٿ�����t�1`%�A<���R�x�h�!�~�e8����������_��c}��������Ȼ��һb�ܻ����L�A�����P���
��x�$���i�k���#!�Xm%��)���-�s�1�6�� :�
!>�B�) F���I���M��Q�AU���X�w�\�CM`�X�c�1g�k��n��r���u���x�\]|�������A9���ᄼY����*��+ˉ��i����������7���͑�9b������􅖼��������0��H����F��iП�Y���ࢼ�g��)�s������}��S��r���f
��;�����ݕ�����靶�E"������,�������7���  �  _bN=��M=a�L=�L=�PK=�J=��I=��H=�6H=fnG=��F=��E=XE=�ED=�yC=s�B=/�A=�A=e>@=�l?=�>=��==S�<=�<=-A;=eg:=�9=�8=^�7=��6=�6=�)5=sC4=_[3=2q2=�1=W�0=��/=[�.=ʼ-=��,=�+=��*=��)=��(=S�'=ϻ&=G�%=��$=�#=){"=c!=�G =�(=�=!�=��=:�=�Z=�&=C�=׳=�t=�1=�=��=!R=��=�=P=K�	=��=k+=C�=hU=��=|p=��<���<���<w��<d��<n��<���<ٝ�<qw�<�J�<!�<���<G��<y]�<=�<���<rr�<.�<X��<	\�<���<�<��<z��<�9�<O®<�G�<�ɧ<�I�<BǠ<{B�<���<33�<
��<��<�<\�<	u�<!�<��z<3�s<�pl<�Re<6^<~W<� P<t�H<��A<��:<��3</�,<�%<��<5�<I�<S�	<��<Y��;o%�;�z�;���;)U�;:ܳ;�t�;� �;�ߋ;�f};,8c;�4I;;^/;��;�y�:c��:2��:��C:I[�9o%7���ù��A�1����ٿ����t�F`%�P<�M�R���h��~�z8������x���y��;}��������Ȼ��һf�ܻ����L�(���,��P���
��x����i�i���#!�Pm%���)���-�w�1�6�� :�!>� B�5 F���I���M��Q��@U���X�k�\�BM`�Y�c�0g��k��n��r��u���x�6]|�Ŀ����79���ᄼQ����*��.ˉ��i����������7���͑�9b���������������0��E����F��mП�Y���ࢼ�g��)�s��!����}��P��u���e
��C������╳����띶�="�����,�������7���  �  VbN=��M=`�L=�L=�PK=��J=��I=��H=�6H=dnG=�F=��E=ZE=�ED=�yC=u�B=/�A=�A=b>@=�l?=�>=��==X�<={<=.A;=dg:=�9=�8=U�7=��6=�6=�)5=rC4=^[3=4q2=�1=^�0=��/=^�.=Ƽ-=��,=�+=��*=��)=��(=W�'=˻&=I�%=��$=�#=1{"=c!=�G =�(=�=�=��=?�=�Z=�&=>�=޳=�t=�1=�=��=%R=��=�=�O=H�	=��=f+=F�=dU=��=|p=��<���<���<��<W��<r��<��<ם�<sw�<�J�<&�<���<R��<v]�<C�<���<lr�<7�<X��<\�<{��<���<��<���<�9�<H®<�G�<�ɧ<�I�<?Ǡ<xB�<���<.3�<��<��<���<U�<
u�<$�<�z<Q�s<�pl<�Re<6^<�W<� P<]�H<��A<��:<��3<*�,<
�%<��<)�<T�<H�	<��<J��;l%�;�z�;���;1U�;�۳;�t�;� �;�ߋ;�f};N8c;�4I;^/;ݵ;9y�:���: ��:��C:�[�9�B9���ù]�A�ƣ��ڿ�5�t�H`%��<���R�y�h�E�~�y8����������]��]}�������Ȼ��һ_�ܻ��滵L�Q���%��P���
��x� ���i�j���#!�am%�ک)���-�x�1��6�� :�!>�B�% F���I���M��Q�AU���X�}�\�.M`�Z�c�,g��k��n��r��u���x�Q]|�ǿ����;9���ᄼ[���{*��1ˉ��i����������7���͑�4b������񅖼��������0��L����F��qП�Y���ࢼ�g��%�s������}��M��{���e
��@�����ҕ���������F"������,��Ʊ���7���  �  RbN=��M=]�L=�L=�PK=��J=��I=��H=�6H=]nG=��F=��E=WE=FD=�yC={�B=+�A=�A=d>@=�l?=�>=��==W�<=w<=6A;=_g:=�9=�8=Q�7=��6=�6=�)5=sC4=\[3=4q2=��1=^�0=��/=c�.=Ƽ-=��,=�+=��*=��)=��(=Z�'=ʻ&=G�%=��$=�#=.{"=c!=�G =�(=�=�=��=A�=�Z=�&=9�=ڳ=�t=�1=�=�=)R=��=�= P=J�	=Đ=e+=K�=aU=��=zp=��<���<���<���<V��<���<��<��<xw�<�J�<4�<���<Q��<t]�<=�<���<ir�<>�<N��<\�<x��<���<��<x��<	:�<:®<�G�<�ɧ<�I�<;Ǡ<}B�<���<&3�<!��<��<��<]�<
u�<0�<٭z<Q�s<�pl<�Re<�5^<�W<� P<k�H<��A<��:<��3<�,<�%<��< �<R�<D�	<��<��;�%�;�z�;���;\U�;�۳;u�;z �;	��;�f};�7c;�4I;^/;ε;�x�:v��:x��:��C:�_�9�/:��ù,�A�C����ٿ�g�t�t`%��<�ڃR�$�h�?�~�A8����������0���}��h����Ȼ��һm�ܻ ��L����
��P�|�
��x���}i�����#!�vm%��)���-�~�1�6�� :�� >�)B� F���I���M��Q�AU���X���\�1M`�c�c�+g��k��n��r��u�c�x�\]|�������E9���ᄼc���|*��3ˉ��i����������7���͑�+b������煖���������0��Z����F��uП�Y���ࢼ�g��%�s��
����}��@��s���e
��4�����ҕ�����ޝ��K"������,�������7���  �  XbN=��M=_�L=�L=�PK=�J=��I=�H=�6H=dnG=��F=��E=WE= FD=�yC=x�B=+�A=�A=e>@=�l?=�>=��==S�<=}<=/A;=cg:=�9=�8=V�7=��6=�6=�)5=sC4=`[3=5q2=�1=[�0=��/=]�.=ļ-=��,=�+=��*=��)=��(=W�'=̻&=H�%=��$=�#=1{"=c!=�G =�(=�= �=��==�=�Z=�&=@�=޳=�t=�1=�=��=%R=��=�=�O=F�	=��=e+=E�=fU=��=~p=��<���<���<y��<W��<p��<��<ܝ�<rw�<�J�<&�<���<J��<]�<G�<���<qr�<6�<P��<\�<���<���<��<s��<:�<I®<�G�<ʧ<�I�<BǠ<yB�<���<.3�<��<��<�<Z�<u�<&�<�z<F�s<�pl<�Re<6^<�W<� P<h�H<��A<��:<��3<(�,<�%<��<1�<J�<\�	<��<I��;�%�;�z�;���;FU�;ܳ;u�;z �;�ߋ;�f};E8c;�4I;j^/;��;}y�:���:���:��C:!]�9�9��ù1�A�����ٿ��t�-`%�<���R���h�b�~�s8����������[��^}������Ȼ��һZ�ܻ}�滷L�F�����P���
��x����i�~���#!�Ym%�۩)���-�p�1�6�� :�!>�B�' F���I���M��Q�AU���X�v�\�4M`�Q�c�$g��k��n��r��u���x�U]|�������<9���ᄼY����*��(ˉ��i����������7���͑�/b������酖���������0��K����F��hП�Y���ࢼ�g��#�s������}��Q��v���m
��?�����ؕ�����᝶�A"������$,�������7���  �  bN=(�M=��L==L=PK=e�J=�I=I�H=�5H=�mG=��F=��E=PE=�DD=�xC=6�B=��A=vA=�<@=@k?=K�>="�==��<=�<=A?;=ae:=�9=Ӭ8=�7=��6=76=�&5=�@4=�X3=bn2= �1=W�0=s�/=$�.=v�-=J�,=��+=$�*=�)=-�(=m�'=׷&=3�%=��$=Ƌ#=�v"=�^!=,C =]$==a�=(�=a�=V=�!=B�=ˮ=�o=�,=��=b�=�L=��=��=�J=%�	=��=N&=2�=eP=��=�k=e��<g��<Q��</��<J��<���<8��<U��<o�<�B�<H�<��<��<`V�<W�<>��<l�<�<���<V�<3�<퇼<��<��<�5�<y��<�C�<�Ƨ<�F�<�Ġ<@�<���<X1�<{��<[�<���<��<�t�<�<Y�z<=�s<orl<Ue<�8^<�W<�P<��H<��A<w�:<��3<Ӱ,<8�%<_�<��</�<��	<��<���;�;�;1��;-��;�n�;��;���;X=�;���;��};�wc;�uI;��/;Y�;��:Hy�:P�:E:(��9��6����@�. ��=3��l��s��	%�W�;��+R��bh�(\~���|˔�l��%�P������ӺȻ0�һ˪ܻtu�"𻣰����-;��
��d�.���U����!��Z%���)� �-���1��6��:��>�B���E�t�I��M�fqQ�"3U�m�X�K�\��@`���c�:sg�r k��n��r��zu�r�x��S|���������4���݄�Z����&���ǉ�f��\�������4���ʑ�_��T򔼄���7�������.��U���E���Ο��W��eߢ��f���쥼�r��-��� }�����΅���	��׍������������䝶�]"��9����,��+���}8���  �  bN=0�M=��L=?L=PK=d�J= �I=D�H=�5H=�mG=��F=��E=LE=�DD=�xC=:�B=��A=xA=�<@=>k?=O�>=�==��<=�<=A?;=ae:=�9=۬8=�7=��6=66='5=�@4=�X3=^n2=��1=X�0=o�/=,�.=|�-=I�,=��+=$�*=�)=-�(=p�'=ҷ&=4�%=��$=ǋ#=�v"=�^!=-C =V$==g�=.�=c�=�U=�!=;�=Ϯ=�o=�,=��=\�=�L=��=��=�J=�	=��=R&=;�=cP=��=�k=Z��<g��<S��<E��<K��<���<-��<`��<-o�<�B�<I�<���<��<UV�<^�<<��<l�<�<}��<�V�<B�<���<��<��<�5�<m��<�C�<�Ƨ<�F�<�Ġ<@�<���<[1�<���<T�<���<��<�t�<�<J�z<:�s<Crl<Ue<�8^<�W<�P<��H<��A<g�:<��3<ܰ,<>�%<X�<��<6�<��	<��<���;�;�;$��;��;�n�;���;���;.=�;���;.�};�wc;�uI;Y�/;��;�:Dy�:P�:�E:���9�m 6����@�����3������o
%�F�;�(,R�jbh��[~����˔�l�����P��q�����Ȼ'�һ�ܻlu��!�ٰ����G;��
��d����U�"���!��Z%���)���-���1��6��:��>�B���E�o�I��M�fqQ�3U�G�X�V�\�~@`��c�Psg�r k��n��r��zu�u�x��S|�k�������4���݄�c����&���ǉ�f��^�������4��
ˑ�x_��F�x���=�������.��a���E���Ο��W��eߢ��f���쥼�r�����}�����Ѕ���	��͍������������睶�c"��2���m,��-����8���  �  bN=.�M=��L=BL=PK=e�J=#�I=@�H=�5H=�mG=��F=��E=ME=�DD=�xC=8�B=��A=~A=�<@=>k?=R�>=�==��<=�<=E?;=`e:=�9=ڬ8=�7=��6=.6=�&5=�@4=�X3=cn2=��1=^�0=j�/=+�.=u�-=H�,=��+=!�*=
�)='�(=v�'=ѷ&=9�%=��$=ǋ#=�v"=�^!=3C =W$==`�=&�=d�=�U=�!=:�=Ү=�o=�,=��=Z�=�L=��=��=�J="�	=��=K&=:�=]P=��=�k=d��<l��<I��<C��<<��<���</��<\��<!o�<�B�<R�<���<���<QV�<a�<=��<l�<+�<}��<�V�<1�<�<��<��<�5�<h��<D�<�Ƨ<�F�<�Ġ<@�<���<N1�<���<R�<���<��<�t�<�<@�z<O�s<Frl<Ue<�8^<�W<�P<��H<��A<d�:<��3<Ű,<K�%<b�<��<D�<��	<��<{��;�;�;F��;��;�n�;j��;���;1=�;���;P�};�wc;'vI;!�/;��;��:�y�:	P�:3E:x��9� 6���ݴ@�����3��b��a�]
%��;��,R�|bh�;\~����˔�0l����$Q��@����Ȼ��һتܻhu��!������E;��
��d�9���U�%���!��Z%���)���-���1��6�:��>�&B���E�}�I���M�dqQ�-3U�L�X�n�\�k@`��c�<sg�h k���n��r��zu�k�x��S|�s�������4���݄�g����&���ǉ�f��\�������4��
ˑ�x_��V򔼀���9�������.��f���E���Ο��W��`ߢ��f���쥼�r��"���	}�����م���	��э������������ܝ��e"��8���s,��8���x8���  �  bN=-�M=��L=AL=PK=d�J=�I=F�H=�5H=�mG=��F=��E=OE=�DD=�xC=8�B=��A=tA=�<@==k?=N�>=�==��<=�<=B?;=be:=�9=ج8=�7=��6=46=�&5=�@4=�X3=_n2=��1=V�0=p�/=.�.=x�-=H�,=��+=$�*=
�)=+�(=r�'=Ϸ&=3�%=��$=ɋ#=�v"=�^!=+C =V$==e�=,�=d�=�U=�!=>�=̮=�o=�,=��=Y�=�L=��=��=�J=#�	=��=P&=<�=cP=��=�k=]��<f��<W��<B��<G��<���<3��<\��<#o�<�B�<L�<���<��<\V�<]�<:��<l�<�<���<�V�<@�<���<��<	��<�5�<n��<�C�<�Ƨ<�F�<�Ġ<@�<���<V1�<���<W�<���<��<�t�<�<Q�z</�s<Url<�Te<�8^<�W<�P<��H<��A<l�:<��3<հ,<H�%<]�<��<3�<��	<��<���;�;�;��;(��;�n�;���;���;H=�;���;v�};�wc;�uI;��/;y�;��:sy�:4P�:�E:���9^6J��v�@�����2��}���M
%�e�;�,R�Obh��[~����˔�l����Q��Z����Ȼ,�һ֪ܻVu��!𻿰��%��F;��
��d����U���!��Z%���)���-���1��6�
:��>�B���E�s�I���M�jqQ�3U�F�X�T�\��@`��c�Isg�t k�څn��r��zu�~�x��S|�t�������4���݄�h����&���ǉ�f��`�������4��ˑ�z_��G�|���7�������.��_���E���Ο��W��fߢ��f���쥼�r��$���}�����Ӆ���	��ɍ������������띶�_"��-���r,��0���8���  �  bN=,�M=��L=>L=PK=h�J=�I=I�H=�5H=�mG=��F=��E=QE=�DD=�xC=1�B=��A=vA=�<@=>k?=N�>="�==��<=�<=@?;=ae:=�9=׬8=�7=��6=:6=�&5=�@4=�X3=bn2=��1=U�0=q�/=%�.={�-=I�,=��+=&�*=�)=,�(=o�'=շ&=4�%=��$=̋#=�v"=�^!=+C =^$==d�=,�=^�=V=�!=B�=ʮ=�o=�,=��=_�=�L=��=��=�J=#�	=��=S&=3�=dP=��=�k=e��<d��<U��<4��<O��<���<6��<[��<%o�<�B�<F�<��<��<_V�<^�<9��<l�<�<���<uV�<E�<<��<��<�5�<u��<�C�<�Ƨ<�F�<�Ġ<@�<���<[1�<���<Z�<���<��<�t�<	�<R�z<-�s<trl<�Te<�8^<�W<�P<��H<��A<v�:<��3<۰,<;�%<[�<��<+�<��	<��<���;�;�;)��;7��;�n�;���;k��;s=�;���;��};�wc;�uI;��/;\�;��:;y�:P�:�E:��9��6	���@������2�����|��	%�t�;�,R��bh��[~����˔�	l���P��z����Ȼ"�һ٪ܻ>u�"𻢰��$��);��
��d����U����!��Z%���)���-���1��6��:��>�B���E�i�I���M�lqQ�3U�g�X�Q�\��@`���c�9sg�x k�܅n��r��zu���x��S|�u�������4���݄�[����&���ǉ�f��a�������4���ʑ��_��B򔼃���8�������.��X��� E���Ο��W��`ߢ��f���쥼�r��&���}�����̅���	��֍������������띶�_"��7���w,��)����8���  �  bN=,�M=��L=DL=PK=a�J="�I=D�H=�5H=�mG=��F=��E=QE=�DD=�xC=5�B=��A=wA=�<@==k?=Q�>=�==��<=�<=C?;=de:=�9=֬8=�7=��6=46=�&5=�@4=�X3=bn2=��1=Z�0=o�/=*�.=z�-=H�,=��+=#�*=�)=,�(=v�'=η&=4�%=��$=ɋ#=�v"=�^!=+C =X$==e�=,�=b�=�U=�!=;�=ή=�o=�,=��=W�=�L=��=��=�J=&�	=��=P&=9�=bP=��=�k=a��<f��<Q��<?��<D��<���<8��<Z��<&o�<�B�<P�<���<��<UV�<b�<9��<l�<�<���<V�<A�<�<��<��<�5�<m��<�C�<�Ƨ<�F�<�Ġ<	@�<���<Y1�<���<S�<��<��<�t�<�<J�z<A�s<Mrl<Ue<�8^<�W<�P<��H<��A<m�:<��3<ְ,<S�%<S�<��<?�<��	<��<���;�;�;"��;3��;�n�;���;���;W=�;���;A�};�wc;!vI;P�/;��;z�:�y�:�P�:�E:���9P�6�����@�@���&3�����w�D
%�/�;�2,R��bh��[~���g˔�"l��
�P��>����Ȼ%�һ�ܻVu��!�ϰ��"��>;� �
��d����U����!��Z%���)���-���1��6�:��>�B���E�t�I��M�iqQ�3U�P�X�Z�\�z@`��c�Bsg�s k��n��r��zu�t�x��S|�x�������4���݄�n����&���ǉ�f��a�������4��ˑ�_��G����4�������.��a���E���Ο��W��hߢ��f���쥼�r��%���}�����ԅ���	��ԍ������������❶�a"��7���r,��3���v8���  �   bN=3�M=��L=AL=PK=`�J=&�I=?�H=�5H=�mG=��F=��E=NE=�DD=�xC=:�B=��A=yA=�<@=:k?=R�>=�==��<=�<=F?;=]e:=�9=ڬ8=�7=��6=16='5=�@4=�X3=cn2=��1=]�0=j�/=.�.=w�-=G�,=��+= �*=�)=%�(=x�'=η&=6�%=��$=Ƌ#=�v"=�^!=2C =S$==c�=)�=f�=�U=�!=:�=ή=�o=�,=��=V�=�L=��=��=�J="�	=��=L&==�=\P=��=�k=a��<i��<J��<G��<?��<���<.��<\��<'o�<�B�<W�<���<���<OV�<b�<6��<l�<#�<|��<�V�<6�<���<��<��<�5�<d��<�C�<�Ƨ<�F�<�Ġ<@�<���<O1�<���<J�<���<��<�t�<�<:�z<J�s<Arl<Ue<�8^<�W<�P<��H<��A<W�:<Ⱥ3<ɰ,<H�%<]�<��<P�<��	<��<`��;�;�;��;��;�n�;}��;���;0=�;���;r�};bwc;1vI;	�/;	�;.�:�y�:�O�:�E:���9P= 6M��6�@�����y3��{��i�g
%� �;��,R�Nbh�\~�'��˔�8l����6Q��.����Ȼ�һ֪ܻtu��!������R;���
��d�)���U�.���!��Z%���)���-���1��6�:��>�,B���E�}�I���M�nqQ�(3U�@�X�o�\�o@`��c�Asg�m k��n��r��zu�s�x��S|�s�������4��}݄�s����&���ǉ�f��d�������4��ˑ�u_��Q�{���9�������.��j���E���Ο�zW��hߢ��f���쥼�r�����}�����؅���	��ύ������������ߝ��g"��5���m,��6���v8���  �  bN=.�M=��L=>L=PK=c�J= �I=E�H=�5H=�mG=��F=��E=PE=�DD=�xC=8�B=��A=uA=�<@==k?=T�>=�==��<=�<=G?;=\e:=�9=׬8=�7=��6=66=�&5=�@4=�X3=bn2=��1=X�0=o�/=)�.=v�-=H�,=��+=#�*=
�)='�(=t�'=շ&=4�%=��$=ʋ#=�v"=�^!=.C =X$==d�=*�=c�=�U=�!==�=ή=�o=�,=��=^�=�L=��=��=�J=%�	=��=M&=7�=aP=��=�k=c��<i��<R��<9��<G��<���<6��<W��<$o�<�B�<T�<���<��<UV�<g�<:��<l�<�<���<�V�<;�<�<��<��<�5�<i��<�C�<�Ƨ<�F�<�Ġ<@�<���<S1�<���<T�<���<��<�t�<�<M�z<6�s<`rl< Ue<�8^<�W<�P<��H<��A<k�:<��3<ΰ,<;�%<n�<��<7�<��	<��<q��;�;�;��;1��;�n�;���;���;R=�;���;z�};�wc;CvI;P�/;��;��:z�:�O�:�E:"��9�h6���	�@�����3��J��z�!
%�P�;�2,R��bh� \~���v˔�$l����%Q��J����Ȼ"�һ֪ܻMu��!�Ѱ����@;��
��d�%���U����!��Z%���)���-���1��6��:��>�'B���E�w�I��M�mqQ�$3U�Y�X�[�\�@`��c�=sg�n k��n��r��zu�w�x��S|�|�������4��݄�e����&���ǉ�f��`�������4��ˑ�{_��L�}���7�������.��e���E���Ο��W��fߢ�}f���쥼�r�� ���}�����҅���	��э������������蝶�`"��4���w,��.���x8���  �  
bN=(�M=��L=?L=PK=d�J= �I=F�H=�5H=�mG=��F=��E=QE=�DD=�xC=3�B=��A=tA=�<@=?k?=N�>= �==��<=�<=@?;=be:=�9=լ8=�7=��6=:6=�&5=�@4=�X3=`n2=��1=S�0=t�/=)�.=}�-=G�,=��+='�*=�)=0�(=o�'=ӷ&=4�%=��$=ɋ#=�v"=�^!=(C =Z$==g�=0�=`�=V=�!=A�=ͮ=�o=�,=��=]�=�L=��=��=�J=%�	=��=T&=6�=gP=��=�k=a��<`��<\��<9��<Q��<���<=��<X��<'o�<�B�<G�<���<��<]V�<\�<=��<l�<�<���<yV�<L�<�<��<��<�5�<t��<�C�<�Ƨ<�F�<�Ġ<@�<���<c1�<z��<_�<�<��<�t�<�<X�z<(�s<lrl<�Te<�8^<�W<�P<��H<��A<��:<��3<�,<>�%<Y�<��<7�<��	<��<���;�;�; ��;3��;�n�;���;x��;d=�;���;h�};�wc;�uI;��/;��;�:1y�:9P�:E:W��9�6F����@�n����2������
%���;��+R��bh��[~�&��~˔�l��!�P��x����Ȼ&�һ˪ܻWu��!𻩰��/��8;�	�
��d����U���!��Z%���)���-���1��6��:��>�B���E�i�I��M�wqQ�3U�[�X�D�\��@`� �c�Bsg�� k�υn��r��zu���x��S|�|�������4���݄�c����&���ǉ�f��]�������4���ʑ��_��<򔼀���8�������.��Z���E���Ο��W��fߢ��f���쥼�r��.����|�����υ���	��ҍ������������흶�]"��4���q,��)����8���  �  bN=+�M=��L=@L=PK=b�J=!�I=C�H=�5H=�mG=��F=��E=QE=�DD=�xC=3�B=��A={A=�<@==k?=O�>=�==��<=�<=D?;=_e:=�9=֬8=�7=��6=66=�&5=�@4=�X3=cn2=��1=Z�0=n�/='�.=z�-=H�,=��+=&�*=�)=*�(=r�'=ӷ&=4�%=��$=ȋ#=�v"=�^!=0C =Z$==b�=)�=a�= V=�!==�=ͮ=�o=�,=��=\�=�L=��=��=�J=#�	=��=P&=6�=aP=��=�k=d��<f��<N��<9��<J��<���<6��<Y��<#o�<�B�<N�<���<��<XV�<]�<;��<l�<%�<���<{V�<<�<퇼<��<��<�5�<i��<�C�<�Ƨ<�F�<�Ġ<@�<���<Y1�<~��<Z�<���<��<�t�<�<G�z<B�s<Yrl<Ue<�8^<�W<�P<��H<��A<v�:<��3<۰,<B�%<b�<��<=�<��	<��<}��;�;�;<��;3��;�n�;���;~��;c=�;���;e�};�wc;�uI;n�/;��;��:�y�:�O�:�E:���9�6���@�r���U3�����e� 
%�)�;�A,R��bh��[~����˔�l��Q��^����Ȼ'�һӪܻbu��!�ʰ����7;��
��d�)���U����!��Z%���)���-���1��6��:��>�B���E�n�I���M�qqQ�3U�]�X�^�\�x@`��c�<sg�s k��n��r��zu���x��S|�y�������4���݄�f����&���ǉ�f��_�������4���ʑ��_��L򔼅���7�������.��e���E���Ο�W��iߢ��f���쥼�r��)���}�����х���	��׍������������᝶�c"��:���r,��.����8���  �  bN=0�M=��L=AL=PK=_�J="�I=A�H=�5H=�mG=��F=��E=NE=�DD=�xC=<�B=��A=wA=�<@=:k?=R�>=�==��<=�<=F?;=be:=�9=ج8=�7=��6=36= '5=�@4=�X3=`n2=�1=[�0=k�/=1�.=v�-=J�,=��+=!�*=�)=*�(=u�'=Ϸ&=2�%=��$=Ƌ#=�v"=�^!=0C =S$==e�=+�=g�=�U=�!=9�=Ю=�o=�,=��=X�=�L=��=��=�J=$�	=��=L&=?�=^P=��=�k=[��<g��<Q��<H��<A��<���<0��<Z��<.o�<�B�<S�<���<��<SV�<`�<8��<l�<�<|��<�V�<8�<���<��<��<�5�<^��< D�<�Ƨ<�F�<�Ġ<@�<���<Z1�<���<M�<���<��<�t�<�<:�z<A�s<9rl<Ue<�8^<�W<�P<��H<��A<\�:<��3<ް,<I�%<d�<}�<A�<��	<��<X��;�;�;��;!��;�n�;���;���;7=�;���;A�};Zwc;#vI;M�/;��;>�:�y�:8P�:�E:���9� 6���˳@������2�������
%��;�o,R�bh�(\~�	��~˔�3l����Q��B����Ȼ2�һتܻpu��!������R;���
��d�#���U�,���!��Z%���)���-���1��6�:��>�B���E�y�I���M�]qQ�(3U�7�X�g�\�w@`��c�Nsg�r k��n��r��zu�h�x��S|�w�������4���݄�o����&���ǉ�f��b�������4��ˑ�s_��P�z���7�������.��o���E���Ο�}W��nߢ��f���쥼�r�����}�����х���	��č������������䝶�h"��*���q,��/���w8���  �  bN=,�M=��L=>L=PK=e�J=$�I=B�H=�5H=�mG=��F=��E=OE=�DD=�xC=6�B=��A=yA=�<@=>k?=M�>=�==��<=�<=B?;=ae:=�9=֬8=�7=��6=56=�&5=�@4=�X3=en2=��1=[�0=k�/=*�.=v�-=I�,=��+="�*=�)=,�(=q�'=ӷ&=8�%=��$=ŋ#=�v"=�^!=1C =Y$==`�='�=c�= V=�!=@�=Ϯ=�o=�,=��=^�=�L=��=��=�J="�	=��=M&=8�=_P=��=�k=g��<d��<O��<=��<D��<���<1��<W��<$o�<�B�<H�<���<���<WV�<X�<<��<l�< �<���<�V�<6�<쇼<��<��<�5�<n��<�C�<�Ƨ<�F�<�Ġ<@�<���<\1�<���<T�<���<��<�t�<�<8�z<J�s<\rl<Ue<�8^<�W<�P<��H<��A<j�:<��3<ܰ,<;�%<Y�<��<G�<��	<��<���;�;�;*��;&��;�n�;��;���;T=�;���;��};�wc;�uI;]�/;��;�:hy�:P�:E:���9g-62��6�@�u���3�����L�
%��;�i,R��bh�+\~����˔�(l��	�P��h����Ȼ �һ��ܻ{u��!𻹰����=;��
��d�1���U����!��Z%���)��-���1��6��:��>�B���E�y�I���M�fqQ�'3U�S�X�d�\�{@`���c�4sg�x k��n��r��zu�v�x��S|�|�������4���݄�b����&���ǉ�f��^�������4�� ˑ�~_��Q򔼅���8�������.��`���E���Ο�{W��bߢ��f���쥼�r��&���}�����Ѕ���	��Ѝ������������ޝ��j"��3���z,��-���}8���  �  bN=)�M=��L=?L=PK=a�J=�I=F�H=�5H=�mG=��F=��E=QE=�DD=�xC=6�B=��A=sA=�<@=?k?=P�>=�==��<=�<=??;=ce:=�9=׬8=�7=��6=;6=�&5=�@4=�X3=_n2=�1=X�0=s�/=)�.=}�-=I�,=��+='�*=�)=1�(=p�'=ӷ&=0�%=��$=ʋ#=�v"=�^!=&C =Y$==f�=/�=a�=V=�!=<�=Ϯ=�o=�,=��=^�=�L=��=��=�J= �	=��=T&=7�=hP=��=�k=\��<e��<[��<<��<Q��<���<2��<\��<#o�<�B�<C�<���<��<YV�<`�<>��<l�<�<���<~V�<M�<�<��<	��<�5�<o��<�C�<�Ƨ<�F�<�Ġ<@�<���<a1�<z��<`�<<��<�t�<�<K�z<;�s<Erl<Ue<�8^<�W<�P<��H<��A<��:<��3<�,<A�%<V�<��<+�<��	<��<���;�;�;��;8��;�n�;���;���;v=�;���;�};�wc;	vI;��/;]�;��:	y�:`P�:E:Y��9��6�����@�j���{2��x����
%�N�;��+R��bh��[~����˔�l���P��n����ȻD�һ�ܻNu��!�ǰ��6��=;��
��d����U���!��Z%���)���-���1��6��:��>��B���E�k�I��M�pqQ�
3U�W�X�B�\��@`��c�Lsg�u k�хn��r��zu���x��S|�s�������4���݄�c����&���ǉ�f��\�������4���ʑ�_��;�~���5�������.��^���E���Ο��W��mߢ��f���쥼�r��-����|�����ʅ���	��ҍ������������杶�a"��2���r,��$����8���  �  bN=,�M=��L=>L=PK=e�J=$�I=B�H=�5H=�mG=��F=��E=OE=�DD=�xC=6�B=��A=yA=�<@=>k?=M�>=�==��<=�<=B?;=ae:=�9=֬8=�7=��6=56=�&5=�@4=�X3=en2=��1=[�0=k�/=*�.=v�-=I�,=��+="�*=�)=,�(=q�'=ӷ&=8�%=��$=ŋ#=�v"=�^!=1C =Y$==`�='�=c�= V=�!=@�=Ϯ=�o=�,=��=^�=�L=��=��=�J="�	=��=L&=8�=_P=��=�k=g��<d��<O��<=��<D��<���<1��<W��<$o�<�B�<H�<���<���<WV�<X�<<��<l�< �<���<�V�<6�<쇼<��<��<�5�<n��<�C�<�Ƨ<�F�<�Ġ<@�<���<\1�<���<T�<���<��<�t�<�<8�z<J�s<\rl<Ue<�8^<�W<�P<��H<��A<j�:<��3<ܰ,<;�%<Y�<��<G�<��	<��<���;�;�;*��;&��;�n�;��;���;T=�;���;��};�wc;�uI;]�/;��;�:hy�:P�:E:���9+-62��6�@�u���3�����L�
%��;�i,R��bh�+\~����˔�(l��	�P��h����Ȼ �һ��ܻ{u��!𻹰����=;��
��d�1���U����!��Z%���)��-���1��6��:��>�B���E�y�I���M�fqQ�'3U�S�X�d�\�{@`���c�4sg�x k��n��r��zu�v�x��S|�|�������4���݄�b����&���ǉ�f��^�������4�� ˑ�~_��Q򔼅���8�������.��`���E���Ο�{W��bߢ��f���쥼�r��&���}�����Ѕ���	��Ѝ������������ޝ��j"��3���z,��-���}8���  �  bN=0�M=��L=AL=PK=_�J="�I=A�H=�5H=�mG=��F=��E=NE=�DD=�xC=<�B=��A=wA=�<@=:k?=R�>=�==��<=�<=F?;=be:=�9=ج8=�7=��6=36= '5=�@4=�X3=`n2=�1=[�0=k�/=1�.=v�-=J�,=��+=!�*=�)=*�(=u�'=Ϸ&=2�%=��$=Ƌ#=�v"=�^!=0C =S$==e�=+�=g�=�U=�!=9�=Ю=�o=�,=��=X�=�L=��=��=�J=$�	=��=L&=?�=^P=��=�k=[��<g��<Q��<H��<A��<���<0��<Z��<.o�<�B�<S�<���<��<SV�<`�<8��<l�<�<|��<�V�<8�<���<��<��<�5�<^��< D�<�Ƨ<�F�<�Ġ<@�<���<Z1�<���<M�<���<��<�t�<�<:�z<A�s<9rl<Ue<�8^<�W<�P<��H<��A<\�:<��3<ް,<I�%<d�<}�<A�<��	<��<X��;�;�;��;!��;�n�;���;���;7=�;���;A�};Zwc;#vI;M�/;��;>�:�y�:8P�:�E:���9� 6���˳@������2�������
%��;�o,R�bh�(\~�	��~˔�3l����Q��B����Ȼ2�һتܻpu��!������R;���
��d�#���U�,���!��Z%���)���-���1��6�:��>�B���E�y�I���M�]qQ�(3U�7�X�g�\�w@`��c�Nsg�r k��n��r��zu�h�x��S|�w�������4���݄�o����&���ǉ�f��b�������4��ˑ�s_��P�z���7�������.��o���E���Ο�}W��nߢ��f���쥼�r�����}�����х���	��č������������䝶�h"��*���q,��/���w8���  �  bN=+�M=��L=@L=PK=b�J=!�I=C�H=�5H=�mG=��F=��E=QE=�DD=�xC=3�B=��A={A=�<@==k?=O�>=�==��<=�<=D?;=_e:=�9=֬8=�7=��6=66=�&5=�@4=�X3=cn2=��1=Z�0=n�/='�.=z�-=H�,=��+=&�*=�)=*�(=r�'=ӷ&=4�%=��$=ȋ#=�v"=�^!=0C =Z$==b�=)�=a�= V=�!==�=ͮ=�o=�,=��=\�=�L=��=��=�J=#�	=��=P&=6�=aP=��=�k=d��<f��<N��<9��<J��<���<6��<Y��<#o�<�B�<N�<���<��<XV�<]�<;��<l�<%�<���<{V�<<�<퇼<��<��<�5�<i��<�C�<�Ƨ<�F�<�Ġ<@�<���<Y1�<~��<Z�<���<��<�t�<�<G�z<B�s<Yrl<Ue<�8^<�W<�P<��H<��A<v�:<��3<۰,<B�%<b�<��<=�<��	<��<}��;�;�;<��;3��;�n�;���;~��;c=�;���;e�};�wc;�uI;n�/;��;��:�y�:�O�:�E:���9��6���@�r���U3�����e� 
%�)�;�A,R��bh��[~����˔�l��Q��^����Ȼ'�һӪܻbu��!�ʰ����7;��
��d�)���U����!��Z%���)���-���1��6��:��>�B���E�n�I���M�qqQ�3U�]�X�^�\�x@`��c�<sg�s k��n��r��zu���x��S|�y�������4���݄�f����&���ǉ�f��_�������4���ʑ��_��L򔼅���7�������.��e���E���Ο�W��iߢ��f���쥼�r��)���}�����х���	��׍������������᝶�c"��:���r,��.����8���  �  
bN=(�M=��L=?L=PK=d�J= �I=F�H=�5H=�mG=��F=��E=QE=�DD=�xC=3�B=��A=tA=�<@=?k?=N�>= �==��<=�<=@?;=be:=�9=լ8=�7=��6=:6=�&5=�@4=�X3=`n2=��1=S�0=t�/=)�.=}�-=G�,=��+='�*=�)=0�(=o�'=ӷ&=4�%=��$=ɋ#=�v"=�^!=(C =Z$==g�=0�=`�=V=�!=A�=ͮ=�o=�,=��=]�=�L=��=��=�J=%�	=��=T&=6�=gP=��=�k=a��<`��<\��<9��<Q��<���<=��<X��<'o�<�B�<G�<���<��<]V�<\�<=��<l�<�<���<yV�<L�<�<��<��<�5�<t��<�C�<�Ƨ<�F�<�Ġ<@�<���<c1�<z��<_�<�<��<�t�<�<X�z<(�s<lrl<�Te<�8^<�W<�P<��H<��A<��:<��3<�,<>�%<Y�<��<7�<��	<��<���;�;�; ��;3��;�n�;���;x��;d=�;���;h�};�wc;�uI;��/;��;�:1y�:8P�:E:V��9��6F����@�n����2������
%���;��+R��bh��[~�&��~˔�l��!�P��x����Ȼ&�һ˪ܻWu��!𻩰��/��8;�	�
��d����U���!��Z%���)���-���1��6��:��>�B���E�i�I��M�wqQ�3U�[�X�D�\��@`� �c�Bsg�� k�υn��r��zu���x��S|�|�������4���݄�c����&���ǉ�f��]�������4���ʑ��_��<򔼀���8�������.��Z���E���Ο��W��fߢ��f���쥼�r��.����|�����υ���	��ҍ������������흶�]"��4���q,��)����8���  �  bN=.�M=��L=>L=PK=c�J= �I=E�H=�5H=�mG=��F=��E=PE=�DD=�xC=8�B=��A=uA=�<@==k?=T�>=�==��<=�<=G?;=\e:=�9=׬8=�7=��6=66=�&5=�@4=�X3=bn2=��1=X�0=o�/=)�.=v�-=H�,=��+=#�*=
�)='�(=t�'=շ&=4�%=��$=ʋ#=�v"=�^!=.C =X$==d�=*�=c�=�U=�!==�=ή=�o=�,=��=^�=�L=��=��=�J=%�	=��=M&=7�=aP=��=�k=c��<i��<R��<9��<G��<���<6��<X��<$o�<�B�<T�<���<��<UV�<g�<:��<l�<�<���<�V�<;�<�<��<��<�5�<i��<�C�<�Ƨ<�F�<�Ġ<@�<���<S1�<���<T�<���<��<�t�<�<M�z<6�s<`rl< Ue<�8^<�W<�P<��H<��A<k�:<��3<ΰ,<;�%<n�<��<7�<��	<��<q��;�;�;��;1��;�n�;���;���;R=�;���;y�};�wc;CvI;P�/;��;��:z�:�O�:�E:!��9�h6���
�@�����3��J��z�!
%�P�;�2,R��bh� \~���v˔�$l����%Q��K����Ȼ"�һ֪ܻMu��!�Ѱ����@;��
��d�%���U����!��Z%���)���-���1��6��:��>�'B���E�w�I��M�mqQ�$3U�Y�X�[�\�@`��c�=sg�n k��n��r��zu�w�x��S|�|�������4��݄�e����&���ǉ�f��`�������4��ˑ�{_��L�}���7�������.��e���E���Ο��W��fߢ�}f���쥼�r�� ���}�����҅���	��э������������蝶�`"��4���w,��.���x8���  �   bN=3�M=��L=AL=PK=`�J=&�I=?�H=�5H=�mG=��F=��E=NE=�DD=�xC=:�B=��A=yA=�<@=:k?=R�>=�==��<=�<=F?;=]e:=�9=ڬ8=�7=��6=16='5=�@4=�X3=cn2=��1=]�0=j�/=.�.=w�-=G�,=��+= �*=�)=%�(=x�'=η&=6�%=��$=Ƌ#=�v"=�^!=2C =S$==c�=)�=f�=�U=�!=:�=ή=�o=�,=��=V�=�L=��=��=�J="�	=��=L&==�=\P=��=�k=a��<i��<J��<G��<?��<���<.��<\��<'o�<�B�<W�<���<���<OV�<b�<6��<l�<#�<|��<�V�<6�<���<��<��<�5�<d��<�C�<�Ƨ<�F�<�Ġ<@�<���<O1�<���<J�<���<��<�t�<�<:�z<J�s<Arl<Ue<�8^<�W<�P<��H<��A<W�:<Ⱥ3<ɰ,<H�%<]�<��<P�<��	<��<`��;�;�;��;��;�n�;}��;���;0=�;���;r�};bwc;1vI;	�/;	�;.�:�y�:�O�:�E:���9�< 6M��6�@�����z3��{��j�g
%� �;��,R�Nbh�\~�'��˔�8l����6Q��.����Ȼ�һ֪ܻtu��!������R;���
��d�)���U�.���!��Z%���)���-���1��6�:��>�,B���E�}�I���M�nqQ�(3U�@�X�o�\�o@`��c�Asg�m k��n��r��zu�s�x��S|�s�������4��}݄�s����&���ǉ�f��d�������4��ˑ�u_��Q�{���9�������.��j���E���Ο�zW��hߢ��f���쥼�r�����}�����؅���	��ύ������������ߝ��g"��5���m,��6���v8���  �  bN=,�M=��L=DL=PK=a�J="�I=D�H=�5H=�mG=��F=��E=QE=�DD=�xC=5�B=��A=wA=�<@==k?=Q�>=�==��<=�<=C?;=de:=�9=֬8=�7=��6=46=�&5=�@4=�X3=bn2=��1=Z�0=o�/=*�.=z�-=H�,=��+=#�*=�)=,�(=v�'=η&=4�%=��$=ɋ#=�v"=�^!=+C =X$==e�=,�=b�=�U=�!=;�=ή=�o=�,=��=W�=�L=��=��=�J=&�	=��=P&=9�=bP=��=�k=a��<f��<Q��<?��<D��<���<8��<Z��<&o�<�B�<P�<���<��<UV�<c�<9��<l�<�<���<V�<A�<�<��<��<�5�<m��<�C�<�Ƨ<�F�<�Ġ<	@�<���<Y1�<���<S�<��<��<�t�<�<J�z<A�s<Mrl<Ue<�8^<�W<�P<��H<��A<m�:<��3<ְ,<S�%<S�<��<?�<��	<��<���;�;�;"��;3��;�n�;���;���;W=�;���;A�};�wc;!vI;P�/;��;z�:�y�:�P�:�E:���9�6�����@�@���'3�����w�D
%�/�;�2,R��bh��[~���g˔�#l��
�P��>����Ȼ%�һ�ܻVu��!�ϰ��"��>;� �
��d����U����!��Z%���)���-���1��6�:��>�B���E�t�I��M�iqQ�3U�P�X�Z�\�z@`��c�Bsg�s k��n��r��zu�t�x��S|�x�������4���݄�n����&���ǉ�f��a�������4��ˑ�_��G����4�������.��a���E���Ο��W��hߢ��f���쥼�r��%���}�����ԅ���	��ԍ������������❶�a"��7���r,��3���v8���  �  bN=,�M=��L=>L=PK=h�J=�I=I�H=�5H=�mG=��F=��E=QE=�DD=�xC=1�B=��A=vA=�<@=>k?=N�>="�==��<=�<=@?;=ae:=�9=׬8=�7=��6=:6=�&5=�@4=�X3=bn2=��1=U�0=q�/=%�.={�-=I�,=��+=&�*=�)=,�(=o�'=շ&=4�%=��$=̋#=�v"=�^!=+C =^$==d�=,�=^�=V=�!=B�=ʮ=�o=�,=��=_�=�L=��=��=�J=#�	=��=S&=3�=dP=��=�k=e��<d��<U��<4��<O��<���<6��<[��<%o�<�B�<F�<��<��<_V�<^�<9��<l�<�<���<uV�<E�<<��<��<�5�<u��<�C�<�Ƨ<�F�<�Ġ<@�<���<[1�<���<Z�<���<��<�t�<	�<R�z<-�s<trl<�Te<�8^<�W<�P<��H<��A<v�:<��3<۰,<;�%<[�<��<+�<��	<��<���;�;�;)��;7��;�n�;���;k��;s=�;���;��};�wc;�uI;��/;\�;��:;y�:P�:�E:��9b�6	���@������2�����|��	%�t�;�,R��bh��[~����˔�	l���P��z����Ȼ"�һ٪ܻ>u�"𻢰��$��);��
��d����U����!��Z%���)���-���1��6��:��>�B���E�i�I���M�lqQ�3U�g�X�Q�\��@`���c�9sg�x k�܅n��r��zu���x��S|�u�������4���݄�[����&���ǉ�f��a�������4���ʑ��_��B򔼃���8�������.��X��� E���Ο��W��`ߢ��f���쥼�r��&���}�����̅���	��֍������������띶�_"��7���w,��)����8���  �  bN=-�M=��L=AL=PK=d�J=�I=F�H=�5H=�mG=��F=��E=OE=�DD=�xC=8�B=��A=tA=�<@==k?=N�>=�==��<=�<=B?;=be:=�9=ج8=�7=��6=46=�&5=�@4=�X3=_n2=��1=V�0=p�/=.�.=x�-=H�,=��+=$�*=
�)=+�(=r�'=Ϸ&=3�%=��$=ɋ#=�v"=�^!=+C =V$==e�=,�=d�=�U=�!=>�=̮=�o=�,=��=Y�=�L=��=��=�J=#�	=��=P&=<�=cP=��=�k=]��<f��<W��<B��<G��<���<3��<\��<#o�<�B�<L�<���<��<\V�<]�<:��<l�<�<���<�V�<@�<���<��<	��<�5�<n��<�C�<�Ƨ<�F�<�Ġ<@�<���<V1�<���<W�<���<��<�t�<�<Q�z</�s<Url<�Te<�8^<�W<�P<��H<��A<l�:<��3<հ,<H�%<]�<��<3�<��	<��<���;�;�;��;(��;�n�;���;���;H=�;���;v�};�wc;�uI;��/;y�;��:sy�:4P�:�E:���96K��w�@�����2��}���M
%�e�;�,R�Obh��[~����˔�l����Q��Z����Ȼ,�һ֪ܻVu��!𻿰��%��F;��
��d����U���!��Z%���)���-���1��6�
:��>�B���E�s�I���M�jqQ�3U�F�X�T�\��@`��c�Isg�t k�څn��r��zu�~�x��S|�t�������4���݄�h����&���ǉ�f��`�������4��ˑ�z_��G�|���7�������.��_���E���Ο��W��fߢ��f���쥼�r��$���}�����Ӆ���	��ɍ������������띶�_"��-���r,��0���8���  �  bN=.�M=��L=BL=PK=e�J=#�I=@�H=�5H=�mG=��F=��E=ME=�DD=�xC=8�B=��A=~A=�<@=>k?=R�>=�==��<=�<=E?;=`e:=�9=ڬ8=�7=��6=.6=�&5=�@4=�X3=cn2=��1=^�0=j�/=+�.=u�-=H�,=��+=!�*=
�)='�(=v�'=ѷ&=9�%=��$=ǋ#=�v"=�^!=3C =W$==`�=&�=d�=�U=�!=:�=Ү=�o=�,=��=Z�=�L=��=��=�J="�	=��=K&=:�=]P=��=�k=d��<l��<I��<C��<<��<���</��<\��<!o�<�B�<R�<���<���<QV�<a�<=��<l�<+�<}��<�V�<1�<�<��<��<�5�<h��<D�<�Ƨ<�F�<�Ġ<@�<���<N1�<���<R�<���<��<�t�<�<@�z<O�s<Frl<Ue<�8^<�W<�P<��H<��A<d�:<��3<Ű,<K�%<b�<��<D�<��	<��<{��;�;�;F��;��;�n�;j��;���;1=�;���;P�};�wc;'vI;!�/;��;��:�y�:	P�:3E:x��9֔ 6���ݴ@�����3��c��a�]
%��;��,R�|bh�;\~����˔�0l����$Q��@����Ȼ��һتܻhu��!������E;��
��d�9���U�%���!��Z%���)���-���1��6�:��>�&B���E�}�I���M�dqQ�-3U�L�X�n�\�k@`��c�<sg�h k���n��r��zu�k�x��S|�s�������4���݄�g����&���ǉ�f��\�������4��
ˑ�x_��V򔼀���9�������.��f���E���Ο��W��`ߢ��f���쥼�r��"���	}�����م���	��э������������ܝ��e"��8���s,��8���x8���  �  bN=0�M=��L=?L=PK=d�J= �I=D�H=�5H=�mG=��F=��E=LE=�DD=�xC=:�B=��A=xA=�<@=>k?=O�>=�==��<=�<=A?;=ae:=�9=۬8=�7=��6=66='5=�@4=�X3=^n2=��1=X�0=o�/=,�.=|�-=I�,=��+=$�*=�)=-�(=p�'=ҷ&=4�%=��$=ǋ#=�v"=�^!=-C =V$==g�=.�=c�=�U=�!=;�=Ϯ=�o=�,=��=\�=�L=��=��=�J=�	=��=R&=;�=cP=��=�k=Z��<g��<S��<E��<K��<���<-��<`��<-o�<�B�<I�<���<��<UV�<^�<<��<l�<�<}��<�V�<B�<���<��<��<�5�<m��<�C�<�Ƨ<�F�<�Ġ<@�<���<[1�<���<T�<���<��<�t�<�<J�z<:�s<Crl<Ue<�8^<�W<�P<��H<��A<g�:<��3<ܰ,<>�%<X�<��<6�<��	<��<���;�;�;$��;��;�n�;���;���;.=�;���;.�};�wc;�uI;Y�/;��;�:Dy�:P�:�E:���9�m 6����@�����3������o
%�F�;�(,R�jbh��[~����˔�l�����P��q�����Ȼ'�һ�ܻlu��!�ٰ����G;��
��d����U�"���!��Z%���)���-���1��6��:��>�B���E�o�I��M�fqQ�3U�G�X�V�\�~@`��c�Psg�r k��n��r��zu�u�x��S|�k�������4���݄�c����&���ǉ�f��^�������4��
ˑ�x_��F�x���=�������.��a���E���Ο��W��eߢ��f���쥼�r�����}�����Ѕ���	��͍������������睶�c"��2���m,��-����8���  �  �aN=
�M=��L=L=�OK=.�J=��I=�H=s5H=HmG=K�F=��E=�E=�DD= xC=ʪB=q�A=A=v<@=�j?=>=��==��<=	<=�>;=�d:=4�9=!�8=T�7=��6=b
6=&5=�?4=�W3=tm2=�1=R�0=f�/=�.=X�-=#�,=]�+=��*=��)=��(='�'=��&=Ԫ%=4�$=a�#=du"=8]!=�A =�"=� =��=��=��=_T=K =��= �=�m=+=.�=��=@K=�=��= I=m�	=�=�$=��=�N='�=�i=1��<8��<2��<��<8��<���<Q��<���<Sl�<@�<��<t��<m��<T�<�<��<�i�<�<���<�T�<x�<N��<6�<���<u4�<1��<�B�<�ŧ<�E�<�à<T?�<߸�<�0�<���<��<���<o�<ot�<�<e�z<{�s<�rl<�Ue<�9^<�W<�P<C�H<G�A<G�:<��3<�,<��%<�<T�<1�< �	<��<���;JC�;���;9 �;Vw�;d��;���;�F�;��;
�};��c;y�I;p�/;W;E6�:l��:���:�|E:���9�j60:���G@�dɏ�]���������$���;�R��Eh�?~�t�������L]��yߩ�/B�������Ȼ��һ��ܻ�f滨�Q���$��G4�:�
��]����kO�����
!�]T%���)���-���1�=�5�Q
:�8>�� B���E�c�I��M��lQ��.U���X��\�P<`���c�3og���j�(�n�\ r�=wu�/�x�mP|�X��"����3��#܄����~%��EƉ��d��?��x����3��ʑ��^��r񔼩���{��͠���-�������D��(Ο��V���ޢ�f���쥼or�������|��L�������	����������������靶�n"��F����,��X����8���  �  �aN=�M=��L=L=�OK=-�J=��I=�H=y5H=BmG=D�F=��E=�E=�DD=$xC=̪B=n�A=A=l<@=�j?=ė>=��==��<=<=�>;=�d:=;�9="�8=N�7=��6=f
6=,&5=�?4=�W3=lm2=��1=U�0=e�/=�.=d�-=(�,=[�+=��*=��)=��(=$�'=}�&=Ԫ%=*�$=Z�#=cu"=+]!=�A =�"=� =��=��=Ą=[T=K =��=�=�m=�*=/�=��==K=�= �=$I=k�	=�=�$=��=�N=)�=�i=��<5��<2��<9��<D��<���<G��<���<gl�<@�<��<k��<s��<�S�<�<��<�i�<�<���<�T�<|�<O��<8�<���<l4�<!��<�B�<�ŧ<�E�<�à<??�<޸�<�0�<��<��<���<y�<�t�<�<`�z<��s<�rl<�Ue<�9^<�W<P<V�H<;�A<?�:<ż3<"�,<��%<��<R�<5�<��	<��<���;C�;��;= �;_w�;���;ϙ�;�F�;��;k�};��c;��I;��/;�;�5�:k��:���:P~E:��9�i67:���F@�mǏ�5���\��^���$��;�#R��Dh�7>~�J���ü��@]��0ߩ�,B������X�Ȼ��һP�ܻg滲𻿢��*��P4�+�
��]�m��[O�����
!��T%���)��-��1�7�5�r
:�E>�� B�e�E�T�I��M��lQ�e.U���X���\�K<`���c�[og���j�'�n�% r�'wu�(�x��P|�N�����3��.܄����x%��^Ɖ��d��F�������3��ʑ��^��n񔼨���y��̠���-�������D��9Ο��V���ޢ�f���쥼jr�������|��T�������	����������������ꝶ�q"��>����,��O����8���  �  �aN=
�M=��L=L=�OK=0�J=��I=�H=5H=DmG=G�F=��E=�E=�DD=xC=ͪB=m�A=A=p<@=�j?=ʗ>=��==�<=<=�>;=�d:=4�9=�8=P�7=��6=_
6=$&5=�?4=�W3=xm2=�1=_�0=`�/=�.=X�-=&�,=^�+=��*=��)=��(=)�'=|�&=ު%=+�$=\�#=hu"=-]!=�A =�"=� =��=��=Ǆ=\T=U =��="�=�m=�*=8�=��=CK=
�=��= I=n�	=�=�$=��=�N=2�=�i=1��<@��<!��<'��<2��<���<L��<���<Wl�<@�<��<m��<���<�S�<�<��<�i�<"�<���<�T�<q�<D��<>�<���<w4�<&��<�B�<�ŧ<�E�<�à<8?�<縙<�0�<���<��<���<r�<{t�<��<`�z<��s<�rl<�Ue<�9^<�W<�P<>�H<K�A<I�:<��3<�,<��%<�<Z�<I�<��	<�<���;*C�;��;K �;Cw�;`��;ә�;�F�;��;��};��c;�I;��/;�;�5�:t��:恔:�|E:���99�i6�6��nH@��ȏ�v���ĺ��h�$�ۛ;�kR�`Eh�?~�V�������X]��Wߩ�NB������b�Ȼ]�һJ�ܻ�f滉𻭢����P4�%�
��]����QO�����
!��T%�y�)���-��1��5�t
:�,>�� B�}�E�e�I��M��lQ��.U���X��\�%<`���c�3og���j�K�n�I r�Jwu��x�vP|�h������3��*܄����i%��bƉ��d��;�������3��ʑ��^��y񔼳���s��ʠ���-������vD��8Ο��V���ޢ�f���쥼vr�������|��M�������	����������������֝��m"��U����,��Z����8���  �  �aN=�M=��L=L=�OK=.�J=��I=�H=v5H=CmG=I�F=��E=�E=�DD=)xC=ΪB=o�A=�A=t<@=�j?=×>=��==��<=<=�>;=�d:=;�9="�8=Q�7=��6=i
6=%&5=�?4=�W3=mm2=��1=R�0=g�/=�.=^�-=+�,=[�+=��*=��)=��(=(�'=}�&=ת%=(�$=^�#=_u"=2]!=�A =�"=� =��=��=ń=YT=I =��=�=�m=�*=0�=��=AK=�= �="I=m�	=�=�$=��=�N='�=�i= ��<5��<4��<,��<G��<���<M��<���<gl�<@�<��<o��<m��<�S�<�<��<�i�<�<���<�T�<��<O��<?�<���<s4�<(��<�B�<�ŧ<�E�<�à<=?�<帙<�0�<��<��<���<��<t�<�<p�z<t�s<�rl<�Ue<�9^<�W<�P<c�H<>�A<G�:<ü3<�,<��%<�<U�<'�<�	<��<���;9C�;���;Q �;\w�;���;���;�F�;T�;�};��c;��I;�/;S;6�:���:䁔:^~E:X��9g�i6�8���E@�Iȏ�F���K��M���$���;��R�Eh��>~�3���ż��E]��*ߩ�%B������Z�Ȼ��һ]�ܻ�f��𻃢��'��`4�(�
��]�j��XO�����
!�xT%���)���-��1�6�5�q
:�5>�� B�c�E�Z�I��M��lQ�t.U���X��\�R<`���c�Uog���j�#�n�? r�!wu��x�uP|�L�����{3��*܄����~%��VƉ��d��I�������3��ʑ��^��e񔼨���r��ܠ���-�������D��-Ο�W���ޢ�f���쥼jr�������|��R�������	����������������񝶼i"��D����,��H����8���  �  �aN=�M=��L=L=�OK=6�J=��I=�H=x5H=EmG=J�F=��E=�E={DD= xC=ªB=x�A=A=v<@=�j?=ė>=��==��<=<=�>;=�d:=:�9=�8=L�7=��6=i
6=&5=�?4=�W3=nm2=�1=T�0=h�/=�.=^�-='�,=U�+=��*=��)=��(="�'=��&=۪%='�$=a�#=_u"=4]!=�A =�"=� =��=��=��=dT=J =��=�=�m=�*=4�=��=;K=
�=��=I=f�	=�=�$=��=�N='�=�i=&��<2��<4��<��<J��<���<C��<���<bl�<@�<��<���<n��<�S�<�<��<�i�<�<���<�T�<u�<:��<A�<���<u4�<*��<�B�<�ŧ<�E�<�à<H?�<ظ�<�0�<���<��<���<z�<|t�<�<p�z<�s<�rl<�Ue<�9^<�W<�P<Z�H<%�A<=�:<��3<�,<��%<��<r�<�<�	<��<���;@C�;��;y �;w�;f��;{��;(G�;��;	�};��c;��I;�/;E;7�:\��:%��:~E:���9��h6�<���E@�*ɏ�[���y��:�2�$���;��R��Eh��>~�N���򼔻Y]��?ߩ�@B��Ɇ���Ȼs�һl�ܻ�f���t���'��04�:�
��]����pO�����
!�kT%���)���-��1�%�5�L
:�L>�� B�p�E�j�I�'�M��lQ�r.U���X��\�Q<`���c�Hog���j�"�n�^ r�wu�4�x��P|�]������3��2܄����|%��VƉ��d��H��z����3���ɑ��^��u񔼽���p��Ơ���-�������D��(Ο�W���ޢ�f���쥼or�������|��]�������	�����������������l"��K����,��L����8���  �  �aN=�M=��L=L=�OK=1�J=��I= �H=~5H=AmG=E�F=��E=�E=�DD=*xC=̪B=o�A=�A=o<@=�j?=ʗ>=��==��<=<=�>;=�d:=6�9=�8=T�7=��6=a
6=%&5=�?4=�W3=rm2=��1=Y�0=g�/=�.=\�-=#�,=_�+=��*=��)=��(=)�'=z�&=ު%=(�$=\�#=gu"=/]!=�A =�"=� =��=��=Ƅ=\T=K =��="�=�m=�*=7�=��=BK=�=��=I=o�	=�=�$=��=�N=-�=�i=&��<<��<1��<*��<:��<���<R��<���<]l�<@�<��<l��<}��<�S�<�<��<�i�<�<���<�T�<��<H��<<�<���<o4�< ��<�B�<�ŧ<�E�<�à<=?�<鸙<�0�<���<��<���<g�<�t�<�<n�z<��s<�rl<�Ue<�9^<�W<�P<4�H<Q�A<L�:<��3<�,<��%<�<`�<<�<��	<�<���;C�;��;P �;Hw�;���;ϙ�;�F�;q�;��};��c;�I;_�/;�;�5�:���:Ձ�:}E:S��9��j6X8���G@�_ȏ�{���ں�	���$�C�;��R�0Eh��>~�q�������\]��>ߩ�8B������m�Ȼa�һd�ܻg滐𻝢��(��T4�,�
��]�r��RO�����
!��T%�|�)���-�%�1��5�x
:�0>�� B�p�E�l�I��M��lQ��.U���X���\�;<`���c�Jog���j�*�n�D r�:wu��x�jP|�f������3��)܄����n%��gƉ��d��?�������3��ʑ��^��c񔼯���u��Ѡ���-������yD��<Ο��V���ޢ�f���쥼wr�������|��H�������	����������������❶�i"��J����,��_����8���  �  �aN=�M=��L=L=�OK=-�J=��I=��H=5H=>mG=S�F=��E=�E=�DD=xC=ѪB=i�A=A=x<@=�j?=ʗ>=��==�<=<=�>;=�d:=;�9=#�8=K�7=��6=b
6=.&5=�?4=�W3=sm2=��1=[�0=^�/=�.=`�-=&�,=]�+=��*=��)=��(=)�'=z�&=ު%=,�$=Z�#=eu"=,]!=�A =�"=� =��=��=Ƅ=UT=W =��= �=�m=�*=:�=��=CK=�=�=I=m�	=�=�$=��=�N=.�=�i=(��<9��<%��<;��<<��<���<D��<���<kl�<	@�<��<d��<���<�S�<�<��<�i�< �<���<�T�<q�<N��<9�<���<�4�<��<�B�<�ŧ<�E�<�à<??�<鸙<�0�<��<��<���<m�<�t�<�<U�z<��s<�rl<�Ue<�9^<�W<P<;�H<K�A<$�:<ؼ3<�,<��%<��<P�<T�<��	<�<y��;�C�;��;6 �;lw�;T��;���;�F�;��;+�};��c;�I;R�/;(;i5�:T��:;��:W~E:ҕ�9��h6e9���G@�(Ǐ�����}������$�(�;��R��Dh�~>~�Y�������~]���ީ�rB������r�Ȼ[�һB�ܻg滜𻰢�����h4�%�
��]����RO�ĳ�
!��T%���)���-��1��5��
:�+>�� B�O�E�m�I��M��lQ�w.U���X��\�7<`���c�Eog���j�B�n�" r�5wu�"�x��P|�S������3��!܄�!���d%��fƉ��d��H��|����3��ʑ��^��y񔼩���x��Ԡ���-��Ĺ��{D��AΟ��V���ޢ�f���쥼{r�������|��J�������	����������������۝��u"��H���,��\����8���  �  �aN=�M=��L=L=�OK=,�J=��I=�H=�5H==mG=L�F=��E=�E=�DD=xC=ΪB=p�A=A=t<@=�j?=˗>=��==��<=<=�>;=�d:==�9=�8=N�7=��6=d
6=&5=�?4=�W3=qm2=�1=Y�0=f�/=�.=\�-=*�,=]�+=��*=��)=��(='�'=��&=ת%=(�$=`�#=fu"=+]!=�A =�"=� =��=��=Ƅ=]T=O =��=�=�m=�*=2�=��=AK=�=�=I=l�	=�=�$=��=�N=-�=�i='��<7��<.��<��<A��<���<I��<���<kl�<@�<��<p��<u��<�S�<�<���<�i�<�<���<�T�<l�<K��<E�<���<x4�<��<�B�<�ŧ<�E�<�à<I?�<ݸ�<�0�<��<��<���<y�<vt�< �<i�z<��s<�rl<�Ue<�9^<�W<�P<J�H<I�A<-�:<ü3<�,<��%<
�<N�<1�<�	<�<q��;QC�;��;g �;Vw�;<��;ߙ�;�F�;��;�};Q�c;�I;ַ/;�;�5�:6��:��:�~E:���9�*i6�8��GG@� ɏ�����Z���;�$�8�;�R�|Eh��>~�;��������]��ߩ�OB������?�Ȼ��һ^�ܻ�f滗𻻢����M4�#�
��]����TO�����
!��T%���)���-��1�/�5�f
:�2>�� B�[�E�z�I��M��lQ�z.U���X���\�8<`���c�Fog���j�0�n�X r�,wu��x�|P|�f������3��#܄����v%��[Ɖ��d��M�������3��ʑ��^��}񔼭���l��Ѡ���-��Ź��wD��.Ο� W���ޢ�f���쥼sr�������|��K�������	����������������杶�m"��M����,��T����8���  �  �aN=�M=��L=L=�OK=1�J=��I=�H=v5H=FmG=G�F=��E=�E=DD=,xC=ɪB=q�A=�A=r<@=�j?=��>=��==��<=<=�>;=�d:=>�9=�8=W�7=��6=h
6="&5=�?4=�W3=jm2=��1=N�0=n�/=�.=b�-=$�,=Z�+=��*=��)=��(="�'=|�&=ت%=*�$=W�#=au"=3]!=�A =�"=� =��=��=��=_T=H =��=�=�m=�*=2�=��=;K=�=��=I=m�	=�=�$=��=�N=$�=�i=��<2��<@��<!��<K��<���<W��<|��<hl�<@�<��<p��<t��<�S�<�<	��<�i�<�<���<�T�<��<B��<<�<���<m4�<-��<�B�<�ŧ<�E�<�à<=?�<ܸ�<�0�<�<��<���<v�<�t�<�<��z<b�s<�rl<�Ue<�9^<�W<�P<V�H<1�A<_�:<��3</�,<��%<�<`�<:�<��	<��<���;'C�;��;Q �;'w�;���;���;�F�;s�;ȸ};݌c;t�I;��/;�;(6�:1��:联:�~E:���9^k6<��F@��ȏ�����7��|���$��;��R�mEh�Z>~�i���Ǽ��K]��Lߩ��A��ʆ��^�Ȼ��һO�ܻ#g滼�{���0��E4�8�
��]�p��iO�����
!�xT%���)��-��1�,�5�q
:�L>�� B�n�E�i�I��M��lQ�d.U���X�ؕ\�\<`���c�\og���j��n�T r�wu�9�x�bP|�p�����z3��2܄����w%��[Ɖ��d��A�������3��ʑ��^��b񔼵���u��Ϡ���-�������D��<Ο��V���ޢ�f���쥼ar�������|��X�������	��������������������a"��D����,��O����8���  �  �aN=�M=��L=L=�OK=1�J=��I=�H=}5H=HmG=J�F=��E=�E=~DD=#xC=ƪB=p�A=A=r<@=�j?=Ɨ>=��==��<=<=�>;=�d:=8�9=�8=T�7=��6=h
6="&5=�?4=�W3=um2=�1=Y�0=c�/=�.=_�-=$�,=Y�+=��*=��)=��(=%�'=��&=ܪ%=.�$=]�#=fu"=1]!=�A =�"=� =��=��=��=^T=R =��=!�=�m=�*=6�=��=@K=	�=��=I=l�	=�=�$=��=�N=+�=�i=1��<9��<'��<!��<H��<���<Q��<���<^l�<@�<��<v��<y��<�S�<�<��<�i�<�<���<�T�<x�<A��<?�<���<z4�<.��<�B�<�ŧ<�E�<�à<I?�<޸�<�0�<���<��<���<r�<�t�<��<k�z<��s<�rl<�Ue<�9^<�W<�P<M�H<&�A<]�:<��3<�,<��%<��<b�<A�<��	<�<���;BC�;���;c �; w�;y��;���;�F�;��;Ը};�c;I;Ƿ/;�;�6�:���:/��:�}E:���9f�j6�<��-F@��ȏ�0���)����C�$�A�;�8R��Eh��>~�k���ϼ��K]��Zߩ�GB������(�Ȼq�һ-�ܻ�f滚𻋢����G4�3�
��]����iO�����
!�{T%�~�)���-��1��5�[
:�6>�� B�|�E�h�I��M��lQ�p.U���X��\�?<`���c�3og���j�>�n�U r�wu�;�x�mP|�f������3��&܄����q%��XƉ��d��;�������3��ʑ��^��r񔼶���r��͠���-������yD��6Ο��V���ޢ�f���쥼rr�������|��\�������	����������������❶�m"��V����,��S����8���  �  �aN=�M=��L=L=�OK=+�J=��I=�H=�5H=>mG=H�F=��E=�E=�DD=$xC=ժB=l�A=�A=p<@=�j?=ɗ>=��==��<=<=�>;=�d:=<�9=!�8=O�7=��6=e
6=%&5=�?4=�W3=nm2=��1=Y�0=d�/= �.=\�-=+�,=^�+=��*=��)=��(=&�'=�&=Ԫ%=(�$=^�#=gu"=']!=�A =�"=� =��=��=ʄ=UT=M =��= �=�m=�*=/�=��=BK=�=�=I=m�	=�=�$=��=�N=.�=�i= ��<:��<1��<.��<?��<���<J��<���<kl�<
@�<��<l��<o��<�S�<�<��<�i�<�<���<�T�<~�<W��<E�<���<v4�<��<�B�<�ŧ<�E�<�à<J?�<ڸ�<�0�<
��<��<���<|�<yt�<�<c�z<��s<�rl<�Ue<�9^<�W<�P<W�H<L�A<7�:<μ3<�,<��%<
�<K�<,�<�	<�<t��;5C�;���;] �;�w�;���;��;�F�;c�;��};��c;�I;��/;w;�5�:��:Ԁ�:�~E:Ԕ�9މi6"8���F@�Qȏ�;���/��D���$�:�;�0R��Dh��>~�0�������r]��	ߩ�NB������J�Ȼ��һ]�ܻ�f滌�ܢ����p4��
��]�l��BO�ó��
!��T%���)���-��1�:�5�n
:�0>�� B�W�E�o�I��M��lQ�.U���X���\�7<`���c�Uog���j�*�n�; r�0wu��x�{P|�W������3��"܄����|%��\Ɖ��d��E�������3��ʑ��^��l񔼠���l��ߠ���-��ɹ��qD��7Ο�W���ޢ�f���쥼tr�������|��J�������	����������������杶�o"��?����,��N����8���  �  �aN=�M=��L=L=�OK=2�J=��I=�H={5H=DmG=Q�F=��E=�E=�DD= xC=˪B=m�A=A={<@=�j?=Ɨ>=��==��<=<=�>;=�d:=6�9=�8=O�7=��6=c
6=&5=�?4=�W3=tm2=�1=V�0=d�/=�.=X�-=%�,=Y�+=��*=��)=��(=$�'=��&=۪%=.�$=Z�#=du"=1]!=�A =�"=� =��=��==\T=T =��=�=�m=�*=5�=��==K=�=��=I=i�	=�=�$=��=�N=+�=�i=+��<6��<1��<��<:��<���<G��<���<Yl�<@�<��<u��<w��<�S�<�<	��<j�< �<���<�T�<s�<@��<=�<���<�4�<&��<�B�<�ŧ<�E�<�à<H?�<ݸ�<�0�<���<��<���<v�<rt�<�<g�z<��s<�rl<�Ue<�9^<�W<�P<L�H<2�A<>�:<��3<�,<��%<��<f�<C�<��	<�<���;~C�;��;D �;2w�;b��;ƙ�;�F�;��;W�};ތc;ŋI;��/;�;�6�:���:H��:}E:͒�9�oi6q;��hG@�ɏ�D��������q�$�m�;�5R�NEh��>~�_���Ҽ��]]��Gߩ�RB������;�Ȼr�һ.�ܻg滣𻌢�����N4�2�
��]����dO�����
!�pT%���)� �-��1�!�5�`
:�E>�� B�w�E�g�I��M��lQ��.U���X��\�B<`���c�>og���j�)�n�[ r�:wu�-�x��P|�^������3��-܄����s%��WƉ��d��A��t����3��ʑ��^��w񔼷���t��ʠ���-������D��;Ο��V���ޢ�f���쥼ur�������|��W�������	����������������᝶�q"��B����,��S����8���  �  �aN=
�M=��L=L=�OK=.�J=��I=�H=~5H=AmG=?�F=��E=�E=�DD=+xC=ƪB=o�A= A=k<@=�j?=ʗ>=��==��<=	<=�>;=�d:=6�9= �8=W�7=��6=l
6=!&5=�?4=�W3=sm2=��1=T�0=i�/=�.=d�-=(�,=Z�+=��*=��)=��(=(�'=~�&=Ѫ%=+�$=^�#=cu"=*]!=�A =�"=� =��=��=��=^T=I =��=�=�m=�*=*�=��=@K=�=��=+I=m�	=�=�$=��=�N='�=�i=$��<0��<3��<!��<T��<���<V��<���<Yl�<"@�<��<t��<g��<�S�<�<���<�i�<�<���<�T�<��<L��<@�<���<g4�<��<�B�<�ŧ<�E�<�à<C?�<<�0�<���< �<���<~�<�t�<�<l�z<��s<�rl<�Ue<�9^<�W<�P<^�H<�A<l�:<��3<�,<̭%<��<U�<4�< �	<�<���;�B�;���;S �;Hw�;���;���;�F�;��;W�};��c;��I;ѷ/;P;O6�:���:���:}E:v��9+]k6m<���D@��ȏ�T���һ�����$���;��R�`Eh�5>~�E���˼���\��]ߩ�,B������K�ȻųһJ�ܻ�f滲�����.��K4�/�
��]�Z��fO�����
!��T%���)���-��1�L�5�f
:�8>�� B��E�7�I�	�M��lQ�U.U���X��\�Q<`���c�Log���j�&�n�U r�wu�*�x�dP|�?�����r3��'܄�����%��XƉ��d��L�������3��ʑ��^��]񔼫���p��Ϡ���-��¹��|D��0Ο��V���ޢ�f���쥼pr�������|��^�������	����������������坶�q"��F����,��J����8���  �  �aN=�M=��L=L=�OK=2�J=��I=�H={5H=DmG=Q�F=��E=�E=�DD= xC=˪B=m�A=A={<@=�j?=Ɨ>=��==��<=<=�>;=�d:=6�9=�8=O�7=��6=c
6=&5=�?4=�W3=tm2=�1=V�0=d�/=�.=X�-=%�,=Y�+=��*=��)=��(=$�'=��&=۪%=.�$=Z�#=du"=1]!=�A =�"=� =��=��==\T=T =��=�=�m=�*=5�=��==K=�=��=I=i�	=�=�$=��=�N=+�=�i=+��<6��<1��<��<:��<���<G��<���<Yl�<@�<��<u��<w��<�S�<�<	��<j�< �<���<�T�<s�<@��<=�<���<�4�<&��<�B�<�ŧ<�E�<�à<H?�<ݸ�<�0�<���<��<���<v�<rt�<�<g�z<��s<�rl<�Ue<�9^<�W<�P<L�H<2�A<>�:<��3<�,<��%<��<f�<C�<��	<�<���;~C�;��;D �;2w�;b��;ƙ�;�F�;��;W�};ތc;ŋI;��/;�;�6�:���:H��:}E:͒�9�oi6q;��iG@�ɏ�D��������q�$�m�;�5R�NEh��>~�_���Ҽ��]]��Gߩ�RB������;�Ȼr�һ.�ܻg滣𻌢�����N4�2�
��]����dO�����
!�pT%���)� �-��1�!�5�`
:�E>�� B�w�E�g�I��M��lQ��.U���X��\�B<`���c�>og���j�)�n�[ r�:wu�-�x��P|�^������3��-܄����s%��WƉ��d��A��t����3��ʑ��^��w񔼷���t��ʠ���-������D��;Ο��V���ޢ�f���쥼ur�������|��W�������	����������������᝶�q"��B����,��S����8���  �  �aN=�M=��L=L=�OK=+�J=��I=�H=�5H=>mG=H�F=��E=�E=�DD=$xC=ժB=l�A=�A=p<@=�j?=ɗ>=��==��<=<=�>;=�d:=<�9=!�8=O�7=��6=e
6=%&5=�?4=�W3=nm2=��1=Y�0=d�/= �.=\�-=+�,=^�+=��*=��)=��(=&�'=�&=Ԫ%=(�$=^�#=gu"=']!=�A =�"=� =��=��=ʄ=UT=M =��= �=�m=�*=/�=��=BK=�=�=I=m�	=�=�$=��=�N=.�=�i= ��<:��<1��<.��<?��<���<J��<���<kl�<
@�<��<l��<o��<�S�<�<��<�i�<�<���<�T�<~�<W��<E�<���<v4�<��<�B�<�ŧ<�E�<�à<J?�<ڸ�<�0�<
��<��<���<|�<yt�<�<c�z<��s<�rl<�Ue<�9^<�W<�P<W�H<L�A<7�:<μ3<�,<��%<
�<K�<,�<�	<�<t��;5C�;���;] �;�w�;���;��;�F�;c�;��};��c;�I;��/;w;�5�:��:Ԁ�:�~E:Ӕ�9ԉi6#8���F@�Qȏ�<���/��E���$�:�;�0R��Dh��>~�0�������r]��	ߩ�NB������J�Ȼ��һ]�ܻ�f滌�ܢ����p4��
��]�l��BO�ó��
!��T%���)���-��1�:�5�n
:�0>�� B�W�E�o�I��M��lQ�.U���X���\�7<`���c�Uog���j�*�n�; r�0wu��x�{P|�W������3��"܄����|%��\Ɖ��d��E�������3��ʑ��^��l񔼠���l��ߠ���-��ɹ��qD��7Ο�W���ޢ�f���쥼tr�������|��J�������	����������������杶�o"��?����,��N����8���  �  �aN=�M=��L=L=�OK=1�J=��I=�H=}5H=HmG=J�F=��E=�E=~DD=#xC=ƪB=p�A=A=r<@=�j?=Ɨ>=��==��<=<=�>;=�d:=8�9=�8=T�7=��6=h
6="&5=�?4=�W3=um2=�1=Y�0=c�/=�.=_�-=$�,=Y�+=��*=��)=��(=%�'=��&=ܪ%=.�$=]�#=fu"=1]!=�A =�"=� =��=��=��=^T=R =��=!�=�m=�*=6�=��=@K=	�=��=I=l�	=�=�$=��=�N=+�=�i=1��<9��<'��<!��<H��<���<Q��<���<^l�<@�<��<w��<y��<�S�<�<��<�i�<�<���<�T�<x�<A��<?�<���<z4�<.��<�B�<�ŧ<�E�<�à<I?�<޸�<�0�<���<��<���<r�<�t�<��<k�z<��s<�rl<�Ue<�9^<�W<�P<M�H<&�A<]�:<��3<�,<��%<��<b�<A�<��	<�<���;BC�;���;c �; w�;y��;���;�F�;��;Ը};�c;I;Ƿ/;�;�6�:���:/��:�}E:���9F�j6�<��-F@��ȏ�0���)����C�$�A�;�8R��Eh��>~�k���ϼ��K]��Zߩ�GB������(�Ȼq�һ-�ܻ�f滚𻋢����G4�3�
��]����iO�����
!�{T%�~�)���-��1��5�[
:�6>�� B�|�E�h�I��M��lQ�p.U���X��\�?<`���c�3og���j�>�n�U r�wu�;�x�mP|�f������3��&܄����q%��XƉ��d��;�������3��ʑ��^��r񔼶���r��͠���-������yD��6Ο��V���ޢ�f���쥼rr�������|��\�������	����������������❶�m"��V����,��S����8���  �  �aN=�M=��L=L=�OK=1�J=��I=�H=v5H=FmG=G�F=��E=�E=DD=,xC=ɪB=q�A=�A=r<@=�j?=��>=��==��<=<=�>;=�d:=>�9=�8=W�7=��6=h
6="&5=�?4=�W3=jm2=��1=N�0=n�/=�.=b�-=$�,=Z�+=��*=��)=��(="�'=|�&=ت%=*�$=W�#=au"=3]!=�A =�"=� =��=��=��=_T=H =��=�=�m=�*=2�=��=;K=�=��=I=m�	=�=�$=��=�N=$�=�i=��<2��<@��<!��<K��<���<W��<|��<hl�<@�<��<p��<t��<�S�<�<	��<�i�<�<���<�T�<��<B��<<�<���<m4�<-��<�B�<�ŧ<�E�<�à<=?�<ܸ�<�0�<�<��<���<v�<�t�<�<��z<b�s<�rl<�Ue<�9^<�W<�P<V�H<0�A<_�:<��3</�,<��%<�<`�<:�<��	<��<���;'C�;��;Q �;'w�;���;���;�F�;s�;ȸ};܌c;t�I;��/;�;(6�:1��:联:�~E:���9�]k6<��F@��ȏ�����7��|���$��;��R�mEh�Z>~�i���Ǽ��K]��Lߩ��A��ʆ��^�Ȼ��һO�ܻ#g滼�{���0��E4�8�
��]�p��iO�����
!�xT%���)��-��1�,�5�q
:�L>�� B�n�E�i�I��M��lQ�d.U���X�ؕ\�\<`���c�\og���j��n�T r�wu�9�x�bP|�p�����z3��2܄����w%��[Ɖ��d��A�������3��ʑ��^��b񔼵���u��Ϡ���-�������D��<Ο��V���ޢ�f���쥼ar�������|��X�������	��������������������a"��D����,��O����8���  �  �aN=�M=��L=L=�OK=,�J=��I=�H=�5H==mG=L�F=��E=�E=�DD=xC=ΪB=p�A=A=t<@=�j?=˗>=��==��<=<=�>;=�d:==�9=�8=N�7=��6=d
6=&5=�?4=�W3=qm2=�1=Y�0=f�/=�.=\�-=*�,=]�+=��*=��)=��(='�'=��&=ת%=(�$=`�#=fu"=+]!=�A =�"=� =��=��=Ƅ=]T=O =��=�=�m=�*=2�=��=AK=�=�=I=l�	=�=�$=��=�N=-�=�i='��<7��<.��< ��<A��<���<I��<���<kl�<@�<��<p��<u��<�S�<�<���<�i�<�<���<�T�<l�<K��<E�<���<x4�<��<�B�<�ŧ<�E�<�à<I?�<ݸ�<�0�<��<��<���<y�<vt�< �<i�z<��s<�rl<�Ue<�9^<�W<�P<J�H<I�A<-�:<ü3<�,<��%<
�<N�<1�<�	<�<q��;QC�;��;g �;Vw�;<��;ߙ�;�F�;��;�};Q�c;�I;շ/;�;�5�:6��:��:�~E:���9�)i6�8��GG@� ɏ�����Z���;�$�8�;�R�|Eh��>~�;��������]��ߩ�OB������?�Ȼ��һ^�ܻ�f滗𻻢����M4�#�
��]����TO�����
!��T%���)���-��1�/�5�f
:�2>�� B�[�E�z�I��M��lQ�z.U���X���\�8<`���c�Fog���j�0�n�X r�,wu��x�|P|�f������3��#܄����v%��[Ɖ��d��M�������3��ʑ��^��}񔼭���l��Ѡ���-��Ź��wD��.Ο� W���ޢ�f���쥼sr�������|��K�������	����������������杶�m"��M����,��T����8���  �  �aN=�M=��L=L=�OK=-�J=��I=��H=5H=>mG=S�F=��E=�E=�DD=xC=ѪB=i�A=A=x<@=�j?=ʗ>=��==�<=<=�>;=�d:=;�9=#�8=K�7=��6=b
6=.&5=�?4=�W3=sm2=��1=[�0=^�/=�.=`�-=&�,=]�+=��*=��)=��(=)�'=z�&=ު%=,�$=Z�#=eu"=,]!=�A =�"=� =��=��=Ƅ=UT=W =��= �=�m=�*=:�=��=CK=�=�=I=m�	=�=�$=��=�N=.�=�i=(��<9��<%��<;��<<��<���<D��<���<kl�<	@�<��<d��<���<�S�<�<��<�i�< �<���<�T�<q�<N��<9�<���<�4�<��<�B�<�ŧ<�E�<�à<??�<鸙<�0�<��<��<���<m�<�t�<�<U�z<��s<�rl<�Ue<�9^<�W<P<;�H<K�A<$�:<ؼ3<�,<��%<��<Q�<T�<��	<�<y��;�C�;��;6 �;lw�;T��;���;�F�;��;+�};��c;�I;R�/;(;i5�:S��:;��:V~E:ҕ�9\�h6e9���G@�(Ǐ�����}������$�(�;��R��Dh�~>~�Y�������~]���ީ�rB������r�Ȼ[�һB�ܻg滝𻰢�����h4�%�
��]����RO�ĳ�
!��T%���)���-��1��5��
:�+>�� B�O�E�m�I��M��lQ�w.U���X��\�7<`���c�Eog���j�B�n�" r�5wu�"�x��P|�S������3��!܄�!���d%��fƉ��d��H��|����3��ʑ��^��y񔼩���x��Ԡ���-��Ĺ��{D��AΟ��V���ޢ�f���쥼{r�������|��J�������	����������������۝��u"��H���,��\����8���  �  �aN=�M=��L=L=�OK=1�J=��I= �H=~5H=AmG=E�F=��E=�E=�DD=*xC=̪B=o�A=�A=o<@=�j?=ʗ>=��==��<=<=�>;=�d:=6�9=�8=T�7=��6=a
6=%&5=�?4=�W3=rm2=��1=Y�0=g�/=�.=\�-=#�,=_�+=��*=��)=��(=)�'=z�&=ު%=(�$=\�#=gu"=/]!=�A =�"=� =��=��=Ƅ=\T=K =��="�=�m=�*=7�=��=BK=�=��=I=o�	=�=�$=��=�N=-�=�i=&��<<��<1��<*��<:��<���<R��<���<]l�<@�<��<l��<}��<�S�<�<��<�i�<�<���<�T�<��<H��<<�<���<o4�< ��<�B�<�ŧ<�E�<�à<=?�<鸙<�0�<���<��<���<g�<�t�<�<n�z<��s<�rl<�Ue<�9^<�W<�P<4�H<Q�A<L�:<��3<�,<��%<�<`�<<�<��	<�<���;C�;��;P �;Hw�;���;ϙ�;�F�;q�;��};��c;�I;_�/;�;�5�:���:Ձ�:}E:R��9��j6Y8���G@�_ȏ�{���ں�	���$�C�;��R�0Eh��>~�q�������\]��>ߩ�9B������m�Ȼa�һd�ܻg滐𻝢��(��T4�,�
��]�r��RO�����
!��T%�|�)���-�%�1��5�x
:�0>�� B�p�E�l�I��M��lQ��.U���X���\�;<`���c�Jog���j�*�n�D r�:wu��x�jP|�f������3��)܄����n%��gƉ��d��?�������3��ʑ��^��c񔼯���u��Ѡ���-������yD��<Ο��V���ޢ�f���쥼wr�������|��H�������	����������������❶�i"��J����,��_����8���  �  �aN=�M=��L=L=�OK=6�J=��I=�H=x5H=EmG=J�F=��E=�E={DD= xC=ªB=x�A=A=v<@=�j?=ė>=��==��<=<=�>;=�d:=:�9=�8=L�7=��6=i
6=&5=�?4=�W3=nm2=�1=T�0=h�/=�.=^�-='�,=U�+=��*=��)=��(="�'=��&=۪%='�$=a�#=_u"=4]!=�A =�"=� =��=��=��=dT=J =��=�=�m=�*=4�=��=;K=
�=��=I=f�	=�=�$=��=�N='�=�i=&��<2��<4��<��<K��<���<C��<���<bl�<@�<��<���<n��<�S�<�<��<�i�<�<���<�T�<u�<:��<A�<���<u4�<*��<�B�<�ŧ<�E�<�à<H?�<ظ�<�0�<���<��<���<z�<|t�<�<p�z<�s<�rl<�Ue<�9^<�W<�P<Z�H<%�A<=�:<��3<�,<��%<��<r�<�<�	<��<���;@C�;��;y �;w�;f��;{��;(G�;��;	�};��c;��I;�/;E;7�:\��:%��:~E:���9��h6�<���E@�*ɏ�[���y��:�2�$���;��R��Eh��>~�N���򼔻Y]��?ߩ�@B��Ɇ���Ȼs�һl�ܻ�f���t���'��04�:�
��]����pO�����
!�kT%���)���-��1�%�5�L
:�L>�� B�p�E�j�I�'�M��lQ�r.U���X��\�Q<`���c�Hog���j�"�n�^ r�wu�4�x��P|�]������3��2܄����|%��VƉ��d��H��z����3���ɑ��^��u񔼽���p��Ơ���-�������D��(Ο�W���ޢ�f���쥼or�������|��]�������	�����������������l"��K����,��L����8���  �  �aN=�M=��L=L=�OK=.�J=��I=�H=v5H=CmG=I�F=��E=�E=�DD=)xC=ΪB=o�A=�A=t<@=�j?=×>=��==��<=<=�>;=�d:=<�9="�8=Q�7=��6=i
6=%&5=�?4=�W3=mm2=��1=R�0=g�/=�.=^�-=+�,=[�+=��*=��)=��(=(�'=}�&=ת%=(�$=^�#=_u"=2]!=�A =�"=� =��=��=ń=YT=I =��=�=�m=�*=0�=��=AK=�= �="I=m�	=�=�$=��=�N='�=�i= ��<5��<4��<,��<G��<���<M��<���<gl�<@�<��<o��<m��<�S�<�<��<�i�<�<���<�T�<��<O��<?�<���<s4�<(��<�B�<�ŧ<�E�<�à<=?�<帙<�0�<��<��<���<��<t�<�<p�z<t�s<�rl<�Ue<�9^<�W<�P<c�H<>�A<G�:<ü3<�,<��%<�<U�<'�<�	<��<���;9C�;���;Q �;\w�;���;���;�F�;T�;�};��c;��I;�/;S;6�:���:ご:^~E:W��9*�i6�8���E@�Iȏ�F���K��M���$���;��R�Eh��>~�3���ż��E]��*ߩ�%B������Z�Ȼ��һ]�ܻ�f��𻃢��'��`4�(�
��]�j��XO�����
!�xT%���)���-��1�6�5�q
:�5>�� B�c�E�Z�I��M��lQ�t.U���X��\�R<`���c�Uog���j�#�n�? r�!wu��x�uP|�L�����{3��*܄����~%��VƉ��d��I�������3��ʑ��^��e񔼨���r��ܠ���-�������D��-Ο�W���ޢ�f���쥼jr�������|��R�������	����������������񝶼i"��D����,��H����8���  �  �aN=
�M=��L=L=�OK=0�J=��I=�H=5H=DmG=G�F=��E=�E=�DD=xC=ͪB=m�A=A=p<@=�j?=ʗ>=��==�<=<=�>;=�d:=4�9=�8=P�7=��6=_
6=$&5=�?4=�W3=xm2=�1=_�0=`�/=�.=X�-=&�,=^�+=��*=��)=��(=)�'=|�&=ު%=+�$=\�#=hu"=-]!=�A =�"=� =��=��=Ǆ=\T=U =��="�=�m=�*=8�=��=CK=
�=��= I=n�	=�=�$=��=�N=2�=�i=1��<@��<!��<'��<2��<���<L��<���<Wl�<@�<��<m��<���<�S�<�<��<�i�<"�<���<�T�<q�<D��<>�<���<w4�<&��<�B�<�ŧ<�E�<�à<8?�<縙<�0�<���<��<���<r�<{t�<��<`�z<��s<�rl<�Ue<�9^<�W<�P<>�H<K�A<I�:<��3<�,<��%<�<Z�<I�<��	<�<���;*C�;��;K �;Cw�;`��;ә�;�F�;��;��};��c;�I;��/;�;�5�:t��:恔:�|E:���9�i6�6��nH@��ȏ�v���ĺ��h�$�ۛ;�kR�`Eh�?~�V�������X]��Wߩ�NB������b�Ȼ]�һJ�ܻ�f滉𻭢����P4�%�
��]����QO�����
!��T%�y�)���-��1��5�t
:�,>�� B�}�E�e�I��M��lQ��.U���X��\�%<`���c�3og���j�K�n�I r�Jwu��x�vP|�h������3��*܄����i%��bƉ��d��;�������3��ʑ��^��y񔼳���s��ʠ���-������vD��8Ο��V���ޢ�f���쥼vr�������|��M�������	����������������֝��m"��U����,��Z����8���  �  �aN=�M=��L=L=�OK=-�J=��I=�H=y5H=BmG=D�F=��E=�E=�DD=$xC=̪B=n�A=A=l<@=�j?=ė>=��==��<=<=�>;=�d:=;�9="�8=N�7=��6=f
6=,&5=�?4=�W3=lm2=��1=U�0=e�/=�.=d�-=(�,=[�+=��*=��)=��(=$�'=}�&=Ԫ%=*�$=Z�#=cu"=+]!=�A =�"=� =��=��=Ą=[T=K =��=�=�m=�*=/�=��==K=�= �=$I=k�	=�=�$=��=�N=)�=�i=��<5��<2��<9��<D��<���<F��<���<gl�<@�<��<k��<s��<�S�<�<��<�i�<�<���<�T�<|�<O��<8�<���<l4�<!��<�B�<�ŧ<�E�<�à<??�<޸�<�0�<��<��<���<y�<�t�<�<`�z<��s<�rl<�Ue<�9^<�W<P<V�H<;�A<?�:<ż3<"�,<��%<��<R�<5�<��	<��<���;C�;��;= �;_w�;���;ϙ�;�F�;��;k�};��c;��I;��/;�;�5�:k��:���:P~E:��9�i67:���F@�mǏ�5���\��^���$��;�#R��Dh�7>~�J���ü��@]��0ߩ�,B������X�Ȼ��һP�ܻg滲𻿢��*��P4�+�
��]�m��[O�����
!��T%���)��-��1�7�5�r
:�E>�� B�e�E�T�I��M��lQ�e.U���X���\�K<`���c�[og���j�'�n�% r�'wu�(�x��P|�N�����3��.܄����x%��^Ɖ��d��F�������3��ʑ��^��n񔼨���y��̠���-�������D��9Ο��V���ޢ�f���쥼jr�������|��S�������	����������������ꝶ�q"��>����,��O����8���  �  bN=(�M=��L==L=PK=e�J=�I=I�H=�5H=�mG=��F=��E=PE=�DD=�xC=6�B=��A=vA=�<@=@k?=K�>="�==��<=�<=A?;=ae:=�9=Ӭ8=�7=��6=76=�&5=�@4=�X3=bn2= �1=W�0=s�/=$�.=v�-=J�,=��+=$�*=�)=-�(=m�'=׷&=3�%=��$=Ƌ#=�v"=�^!=,C =]$==a�=(�=a�=V=�!=B�=ˮ=�o=�,=��=b�=�L=��=��=�J=%�	=��=N&=2�=eP=��=�k=e��<g��<Q��</��<J��<���<8��<U��<o�<�B�<H�<��<��<`V�<W�<>��<l�<�<���<V�<3�<퇼<��<��<�5�<y��<�C�<�Ƨ<�F�<�Ġ<@�<���<X1�<{��<[�<���<��<�t�<�<Y�z<=�s<orl<Ue<�8^<�W<�P<��H<��A<w�:<��3<Ӱ,<8�%<_�<��</�<��	<��<���;�;�;1��;-��;�n�;��;���;X=�;���;��};�wc;�uI;��/;Y�;��:Hy�:P�:E:(��9��6����@�. ��=3��l��s��	%�W�;��+R��bh�(\~���|˔�l��%�P������ӺȻ0�һ˪ܻtu�"𻣰����-;��
��d�.���U����!��Z%���)� �-���1��6��:��>�B���E�t�I��M�fqQ�"3U�m�X�K�\��@`���c�:sg�r k��n��r��zu�r�x��S|���������4���݄�Z����&���ǉ�f��\�������4���ʑ�_��T򔼄���7�������.��U���E���Ο��W��eߢ��f���쥼�r��-��� }�����΅���	��׍������������䝶�]"��9����,��+���}8���  �  bN=0�M=��L=?L=PK=d�J= �I=D�H=�5H=�mG=��F=��E=LE=�DD=�xC=:�B=��A=xA=�<@=>k?=O�>=�==��<=�<=A?;=ae:=�9=۬8=�7=��6=66='5=�@4=�X3=^n2=��1=X�0=o�/=,�.=|�-=I�,=��+=$�*=�)=-�(=p�'=ҷ&=4�%=��$=ǋ#=�v"=�^!=-C =V$==g�=.�=c�=�U=�!=;�=Ϯ=�o=�,=��=\�=�L=��=��=�J=�	=��=R&=;�=cP=��=�k=Z��<g��<S��<E��<K��<���<-��<`��<-o�<�B�<I�<���<��<UV�<^�<<��<l�<�<}��<�V�<B�<���<��<��<�5�<m��<�C�<�Ƨ<�F�<�Ġ<@�<���<[1�<���<T�<���<��<�t�<�<J�z<:�s<Crl<Ue<�8^<�W<�P<��H<��A<g�:<��3<ܰ,<>�%<X�<��<6�<��	<��<���;�;�;$��;��;�n�;���;���;.=�;���;.�};�wc;�uI;Y�/;��;�:Dy�:P�:�E:���9�m 6����@�����3������o
%�F�;�(,R�jbh��[~����˔�l�����P��q�����Ȼ'�һ�ܻlu��!�ٰ����G;��
��d����U�"���!��Z%���)���-���1��6��:��>�B���E�o�I��M�fqQ�3U�G�X�V�\�~@`��c�Psg�r k��n��r��zu�u�x��S|�k�������4���݄�c����&���ǉ�f��^�������4��
ˑ�x_��F�x���=�������.��a���E���Ο��W��eߢ��f���쥼�r�����}�����Ѕ���	��͍������������睶�c"��2���m,��-����8���  �  bN=.�M=��L=BL=PK=e�J=#�I=@�H=�5H=�mG=��F=��E=ME=�DD=�xC=8�B=��A=~A=�<@=>k?=R�>=�==��<=�<=E?;=`e:=�9=ڬ8=�7=��6=.6=�&5=�@4=�X3=cn2=��1=^�0=j�/=+�.=u�-=H�,=��+=!�*=
�)='�(=v�'=ѷ&=9�%=��$=ǋ#=�v"=�^!=3C =W$==`�=&�=d�=�U=�!=:�=Ү=�o=�,=��=Z�=�L=��=��=�J="�	=��=K&=:�=]P=��=�k=d��<l��<I��<C��<<��<���</��<\��<!o�<�B�<R�<���<���<QV�<a�<=��<l�<+�<}��<�V�<1�<�<��<��<�5�<h��<D�<�Ƨ<�F�<�Ġ<@�<���<N1�<���<R�<���<��<�t�<�<@�z<O�s<Frl<Ue<�8^<�W<�P<��H<��A<d�:<��3<Ű,<K�%<b�<��<D�<��	<��<{��;�;�;F��;��;�n�;j��;���;1=�;���;P�};�wc;'vI;!�/;��;��:�y�:	P�:3E:x��9� 6���ݴ@�����3��b��a�]
%��;��,R�|bh�;\~����˔�0l����$Q��@����Ȼ��һتܻhu��!������E;��
��d�9���U�%���!��Z%���)���-���1��6�:��>�&B���E�}�I���M�dqQ�-3U�L�X�n�\�k@`��c�<sg�h k���n��r��zu�k�x��S|�s�������4���݄�g����&���ǉ�f��\�������4��
ˑ�x_��V򔼀���9�������.��f���E���Ο��W��`ߢ��f���쥼�r��"���	}�����م���	��э������������ܝ��e"��8���s,��8���x8���  �  bN=-�M=��L=AL=PK=d�J=�I=F�H=�5H=�mG=��F=��E=OE=�DD=�xC=8�B=��A=tA=�<@==k?=N�>=�==��<=�<=B?;=be:=�9=ج8=�7=��6=46=�&5=�@4=�X3=_n2=��1=V�0=p�/=.�.=x�-=H�,=��+=$�*=
�)=+�(=r�'=Ϸ&=3�%=��$=ɋ#=�v"=�^!=+C =V$==e�=,�=d�=�U=�!=>�=̮=�o=�,=��=Y�=�L=��=��=�J=#�	=��=P&=<�=cP=��=�k=]��<f��<W��<B��<G��<���<3��<\��<#o�<�B�<L�<���<��<\V�<]�<:��<l�<�<���<�V�<@�<���<��<	��<�5�<n��<�C�<�Ƨ<�F�<�Ġ<@�<���<V1�<���<W�<���<��<�t�<�<Q�z</�s<Url<�Te<�8^<�W<�P<��H<��A<l�:<��3<հ,<H�%<]�<��<3�<��	<��<���;�;�;��;(��;�n�;���;���;H=�;���;v�};�wc;�uI;��/;y�;��:sy�:4P�:�E:���9^6J��v�@�����2��}���M
%�e�;�,R�Obh��[~����˔�l����Q��Z����Ȼ,�һ֪ܻVu��!𻿰��%��F;��
��d����U���!��Z%���)���-���1��6�
:��>�B���E�s�I���M�jqQ�3U�F�X�T�\��@`��c�Isg�t k�څn��r��zu�~�x��S|�t�������4���݄�h����&���ǉ�f��`�������4��ˑ�z_��G�|���7�������.��_���E���Ο��W��fߢ��f���쥼�r��$���}�����Ӆ���	��ɍ������������띶�_"��-���r,��0���8���  �  bN=,�M=��L=>L=PK=h�J=�I=I�H=�5H=�mG=��F=��E=QE=�DD=�xC=1�B=��A=vA=�<@=>k?=N�>="�==��<=�<=@?;=ae:=�9=׬8=�7=��6=:6=�&5=�@4=�X3=bn2=��1=U�0=q�/=%�.={�-=I�,=��+=&�*=�)=,�(=o�'=շ&=4�%=��$=̋#=�v"=�^!=+C =^$==d�=,�=^�=V=�!=B�=ʮ=�o=�,=��=_�=�L=��=��=�J=#�	=��=S&=3�=dP=��=�k=e��<d��<U��<4��<O��<���<6��<[��<%o�<�B�<F�<��<��<_V�<^�<9��<l�<�<���<uV�<E�<<��<��<�5�<u��<�C�<�Ƨ<�F�<�Ġ<@�<���<[1�<���<Z�<���<��<�t�<	�<R�z<-�s<trl<�Te<�8^<�W<�P<��H<��A<v�:<��3<۰,<;�%<[�<��<+�<��	<��<���;�;�;)��;7��;�n�;���;k��;s=�;���;��};�wc;�uI;��/;\�;��:;y�:P�:�E:��9��6	���@������2�����|��	%�t�;�,R��bh��[~����˔�	l���P��z����Ȼ"�һ٪ܻ>u�"𻢰��$��);��
��d����U����!��Z%���)���-���1��6��:��>�B���E�i�I���M�lqQ�3U�g�X�Q�\��@`���c�9sg�x k�܅n��r��zu���x��S|�u�������4���݄�[����&���ǉ�f��a�������4���ʑ��_��B򔼃���8�������.��X��� E���Ο��W��`ߢ��f���쥼�r��&���}�����̅���	��֍������������띶�_"��7���w,��)����8���  �  bN=,�M=��L=DL=PK=a�J="�I=D�H=�5H=�mG=��F=��E=QE=�DD=�xC=5�B=��A=wA=�<@==k?=Q�>=�==��<=�<=C?;=de:=�9=֬8=�7=��6=46=�&5=�@4=�X3=bn2=��1=Z�0=o�/=*�.=z�-=H�,=��+=#�*=�)=,�(=v�'=η&=4�%=��$=ɋ#=�v"=�^!=+C =X$==e�=,�=b�=�U=�!=;�=ή=�o=�,=��=W�=�L=��=��=�J=&�	=��=P&=9�=bP=��=�k=a��<f��<Q��<?��<D��<���<8��<Z��<&o�<�B�<P�<���<��<UV�<b�<9��<l�<�<���<V�<A�<�<��<��<�5�<m��<�C�<�Ƨ<�F�<�Ġ<	@�<���<Y1�<���<S�<��<��<�t�<�<J�z<A�s<Mrl<Ue<�8^<�W<�P<��H<��A<m�:<��3<ְ,<S�%<S�<��<?�<��	<��<���;�;�;"��;3��;�n�;���;���;W=�;���;A�};�wc;!vI;P�/;��;z�:�y�:�P�:�E:���9P�6�����@�@���&3�����w�D
%�/�;�2,R��bh��[~���g˔�"l��
�P��>����Ȼ%�һ�ܻVu��!�ϰ��"��>;� �
��d����U����!��Z%���)���-���1��6�:��>�B���E�t�I��M�iqQ�3U�P�X�Z�\�z@`��c�Bsg�s k��n��r��zu�t�x��S|�x�������4���݄�n����&���ǉ�f��a�������4��ˑ�_��G����4�������.��a���E���Ο��W��hߢ��f���쥼�r��%���}�����ԅ���	��ԍ������������❶�a"��7���r,��3���v8���  �   bN=3�M=��L=AL=PK=`�J=&�I=?�H=�5H=�mG=��F=��E=NE=�DD=�xC=:�B=��A=yA=�<@=:k?=R�>=�==��<=�<=F?;=]e:=�9=ڬ8=�7=��6=16='5=�@4=�X3=cn2=��1=]�0=j�/=.�.=w�-=G�,=��+= �*=�)=%�(=x�'=η&=6�%=��$=Ƌ#=�v"=�^!=2C =S$==c�=)�=f�=�U=�!=:�=ή=�o=�,=��=V�=�L=��=��=�J="�	=��=L&==�=\P=��=�k=a��<i��<J��<G��<?��<���<.��<\��<'o�<�B�<W�<���<���<OV�<b�<6��<l�<#�<|��<�V�<6�<���<��<��<�5�<d��<�C�<�Ƨ<�F�<�Ġ<@�<���<O1�<���<J�<���<��<�t�<�<:�z<J�s<Arl<Ue<�8^<�W<�P<��H<��A<W�:<Ⱥ3<ɰ,<H�%<]�<��<P�<��	<��<`��;�;�;��;��;�n�;}��;���;0=�;���;r�};bwc;1vI;	�/;	�;.�:�y�:�O�:�E:���9P= 6M��6�@�����y3��{��i�g
%� �;��,R�Nbh�\~�'��˔�8l����6Q��.����Ȼ�һ֪ܻtu��!������R;���
��d�)���U�.���!��Z%���)���-���1��6�:��>�,B���E�}�I���M�nqQ�(3U�@�X�o�\�o@`��c�Asg�m k��n��r��zu�s�x��S|�s�������4��}݄�s����&���ǉ�f��d�������4��ˑ�u_��Q�{���9�������.��j���E���Ο�zW��hߢ��f���쥼�r�����}�����؅���	��ύ������������ߝ��g"��5���m,��6���v8���  �  bN=.�M=��L=>L=PK=c�J= �I=E�H=�5H=�mG=��F=��E=PE=�DD=�xC=8�B=��A=uA=�<@==k?=T�>=�==��<=�<=G?;=\e:=�9=׬8=�7=��6=66=�&5=�@4=�X3=bn2=��1=X�0=o�/=)�.=v�-=H�,=��+=#�*=
�)='�(=t�'=շ&=4�%=��$=ʋ#=�v"=�^!=.C =X$==d�=*�=c�=�U=�!==�=ή=�o=�,=��=^�=�L=��=��=�J=%�	=��=M&=7�=aP=��=�k=c��<i��<R��<9��<G��<���<6��<W��<$o�<�B�<T�<���<��<UV�<g�<:��<l�<�<���<�V�<;�<�<��<��<�5�<i��<�C�<�Ƨ<�F�<�Ġ<@�<���<S1�<���<T�<���<��<�t�<�<M�z<6�s<`rl< Ue<�8^<�W<�P<��H<��A<k�:<��3<ΰ,<;�%<n�<��<7�<��	<��<q��;�;�;��;1��;�n�;���;���;R=�;���;z�};�wc;CvI;P�/;��;��:z�:�O�:�E:"��9�h6���	�@�����3��J��z�!
%�P�;�2,R��bh� \~���v˔�$l����%Q��J����Ȼ"�һ֪ܻMu��!�Ѱ����@;��
��d�%���U����!��Z%���)���-���1��6��:��>�'B���E�w�I��M�mqQ�$3U�Y�X�[�\�@`��c�=sg�n k��n��r��zu�w�x��S|�|�������4��݄�e����&���ǉ�f��`�������4��ˑ�{_��L�}���7�������.��e���E���Ο��W��fߢ�}f���쥼�r�� ���}�����҅���	��э������������蝶�`"��4���w,��.���x8���  �  
bN=(�M=��L=?L=PK=d�J= �I=F�H=�5H=�mG=��F=��E=QE=�DD=�xC=3�B=��A=tA=�<@=?k?=N�>= �==��<=�<=@?;=be:=�9=լ8=�7=��6=:6=�&5=�@4=�X3=`n2=��1=S�0=t�/=)�.=}�-=G�,=��+='�*=�)=0�(=o�'=ӷ&=4�%=��$=ɋ#=�v"=�^!=(C =Z$==g�=0�=`�=V=�!=A�=ͮ=�o=�,=��=]�=�L=��=��=�J=%�	=��=T&=6�=gP=��=�k=a��<`��<\��<9��<Q��<���<=��<X��<'o�<�B�<G�<���<��<]V�<\�<=��<l�<�<���<yV�<L�<�<��<��<�5�<t��<�C�<�Ƨ<�F�<�Ġ<@�<���<c1�<z��<_�<�<��<�t�<�<X�z<(�s<lrl<�Te<�8^<�W<�P<��H<��A<��:<��3<�,<>�%<Y�<��<7�<��	<��<���;�;�; ��;3��;�n�;���;x��;d=�;���;h�};�wc;�uI;��/;��;�:1y�:9P�:E:W��9�6F����@�n����2������
%���;��+R��bh��[~�&��~˔�l��!�P��x����Ȼ&�һ˪ܻWu��!𻩰��/��8;�	�
��d����U���!��Z%���)���-���1��6��:��>�B���E�i�I��M�wqQ�3U�[�X�D�\��@`� �c�Bsg�� k�υn��r��zu���x��S|�|�������4���݄�c����&���ǉ�f��]�������4���ʑ��_��<򔼀���8�������.��Z���E���Ο��W��fߢ��f���쥼�r��.����|�����υ���	��ҍ������������흶�]"��4���q,��)����8���  �  bN=+�M=��L=@L=PK=b�J=!�I=C�H=�5H=�mG=��F=��E=QE=�DD=�xC=3�B=��A={A=�<@==k?=O�>=�==��<=�<=D?;=_e:=�9=֬8=�7=��6=66=�&5=�@4=�X3=cn2=��1=Z�0=n�/='�.=z�-=H�,=��+=&�*=�)=*�(=r�'=ӷ&=4�%=��$=ȋ#=�v"=�^!=0C =Z$==b�=)�=a�= V=�!==�=ͮ=�o=�,=��=\�=�L=��=��=�J=#�	=��=P&=6�=aP=��=�k=d��<f��<N��<9��<J��<���<6��<Y��<#o�<�B�<N�<���<��<XV�<]�<;��<l�<%�<���<{V�<<�<퇼<��<��<�5�<i��<�C�<�Ƨ<�F�<�Ġ<@�<���<Y1�<~��<Z�<���<��<�t�<�<G�z<B�s<Yrl<Ue<�8^<�W<�P<��H<��A<v�:<��3<۰,<B�%<b�<��<=�<��	<��<}��;�;�;<��;3��;�n�;���;~��;c=�;���;e�};�wc;�uI;n�/;��;��:�y�:�O�:�E:���9�6���@�r���U3�����e� 
%�)�;�A,R��bh��[~����˔�l��Q��^����Ȼ'�һӪܻbu��!�ʰ����7;��
��d�)���U����!��Z%���)���-���1��6��:��>�B���E�n�I���M�qqQ�3U�]�X�^�\�x@`��c�<sg�s k��n��r��zu���x��S|�y�������4���݄�f����&���ǉ�f��_�������4���ʑ��_��L򔼅���7�������.��e���E���Ο�W��iߢ��f���쥼�r��)���}�����х���	��׍������������᝶�c"��:���r,��.����8���  �  bN=0�M=��L=AL=PK=_�J="�I=A�H=�5H=�mG=��F=��E=NE=�DD=�xC=<�B=��A=wA=�<@=:k?=R�>=�==��<=�<=F?;=be:=�9=ج8=�7=��6=36= '5=�@4=�X3=`n2=�1=[�0=k�/=1�.=v�-=J�,=��+=!�*=�)=*�(=u�'=Ϸ&=2�%=��$=Ƌ#=�v"=�^!=0C =S$==e�=+�=g�=�U=�!=9�=Ю=�o=�,=��=X�=�L=��=��=�J=$�	=��=L&=?�=^P=��=�k=[��<g��<Q��<H��<A��<���<0��<Z��<.o�<�B�<S�<���<��<SV�<`�<8��<l�<�<|��<�V�<8�<���<��<��<�5�<^��< D�<�Ƨ<�F�<�Ġ<@�<���<Z1�<���<M�<���<��<�t�<�<:�z<A�s<9rl<Ue<�8^<�W<�P<��H<��A<\�:<��3<ް,<I�%<d�<}�<A�<��	<��<X��;�;�;��;!��;�n�;���;���;7=�;���;A�};Zwc;#vI;M�/;��;>�:�y�:8P�:�E:���9� 6���˳@������2�������
%��;�o,R�bh�(\~�	��~˔�3l����Q��B����Ȼ2�һتܻpu��!������R;���
��d�#���U�,���!��Z%���)���-���1��6�:��>�B���E�y�I���M�]qQ�(3U�7�X�g�\�w@`��c�Nsg�r k��n��r��zu�h�x��S|�w�������4���݄�o����&���ǉ�f��b�������4��ˑ�s_��P�z���7�������.��o���E���Ο�}W��nߢ��f���쥼�r�����}�����х���	��č������������䝶�h"��*���q,��/���w8���  �  bN=,�M=��L=>L=PK=e�J=$�I=B�H=�5H=�mG=��F=��E=OE=�DD=�xC=6�B=��A=yA=�<@=>k?=M�>=�==��<=�<=B?;=ae:=�9=֬8=�7=��6=56=�&5=�@4=�X3=en2=��1=[�0=k�/=*�.=v�-=I�,=��+="�*=�)=,�(=q�'=ӷ&=8�%=��$=ŋ#=�v"=�^!=1C =Y$==`�='�=c�= V=�!=@�=Ϯ=�o=�,=��=^�=�L=��=��=�J="�	=��=M&=8�=_P=��=�k=g��<d��<O��<=��<D��<���<1��<W��<$o�<�B�<H�<���<���<WV�<X�<<��<l�< �<���<�V�<6�<쇼<��<��<�5�<n��<�C�<�Ƨ<�F�<�Ġ<@�<���<\1�<���<T�<���<��<�t�<�<8�z<J�s<\rl<Ue<�8^<�W<�P<��H<��A<j�:<��3<ܰ,<;�%<Y�<��<G�<��	<��<���;�;�;*��;&��;�n�;��;���;T=�;���;��};�wc;�uI;]�/;��;�:hy�:P�:E:���9g-62��6�@�u���3�����L�
%��;�i,R��bh�+\~����˔�(l��	�P��h����Ȼ �һ��ܻ{u��!𻹰����=;��
��d�1���U����!��Z%���)��-���1��6��:��>�B���E�y�I���M�fqQ�'3U�S�X�d�\�{@`���c�4sg�x k��n��r��zu�v�x��S|�|�������4���݄�b����&���ǉ�f��^�������4�� ˑ�~_��Q򔼅���8�������.��`���E���Ο�{W��bߢ��f���쥼�r��&���}�����Ѕ���	��Ѝ������������ޝ��j"��3���z,��-���}8���  �  bN=)�M=��L=?L=PK=a�J=�I=F�H=�5H=�mG=��F=��E=QE=�DD=�xC=6�B=��A=sA=�<@=?k?=P�>=�==��<=�<=??;=ce:=�9=׬8=�7=��6=;6=�&5=�@4=�X3=_n2=�1=X�0=s�/=)�.=}�-=I�,=��+='�*=�)=1�(=p�'=ӷ&=0�%=��$=ʋ#=�v"=�^!=&C =Y$==f�=/�=a�=V=�!=<�=Ϯ=�o=�,=��=^�=�L=��=��=�J= �	=��=T&=7�=hP=��=�k=\��<e��<[��<<��<Q��<���<2��<\��<#o�<�B�<C�<���<��<YV�<`�<>��<l�<�<���<~V�<M�<�<��<	��<�5�<o��<�C�<�Ƨ<�F�<�Ġ<@�<���<a1�<z��<`�<<��<�t�<�<K�z<;�s<Erl<Ue<�8^<�W<�P<��H<��A<��:<��3<�,<A�%<V�<��<+�<��	<��<���;�;�;��;8��;�n�;���;���;v=�;���;�};�wc;	vI;��/;]�;��:	y�:`P�:E:Y��9��6�����@�j���{2��x����
%�N�;��+R��bh��[~����˔�l���P��n����ȻD�һ�ܻNu��!�ǰ��6��=;��
��d����U���!��Z%���)���-���1��6��:��>��B���E�k�I��M�pqQ�
3U�W�X�B�\��@`��c�Lsg�u k�хn��r��zu���x��S|�s�������4���݄�c����&���ǉ�f��\�������4���ʑ�_��;�~���5�������.��^���E���Ο��W��mߢ��f���쥼�r��-����|�����ʅ���	��ҍ������������杶�a"��2���r,��$����8���  �  bN=,�M=��L=>L=PK=e�J=$�I=B�H=�5H=�mG=��F=��E=OE=�DD=�xC=6�B=��A=yA=�<@=>k?=M�>=�==��<=�<=B?;=ae:=�9=֬8=�7=��6=56=�&5=�@4=�X3=en2=��1=[�0=k�/=*�.=v�-=I�,=��+="�*=�)=,�(=q�'=ӷ&=8�%=��$=ŋ#=�v"=�^!=1C =Y$==`�='�=c�= V=�!=@�=Ϯ=�o=�,=��=^�=�L=��=��=�J="�	=��=L&=8�=_P=��=�k=g��<d��<O��<=��<D��<���<1��<W��<$o�<�B�<H�<���<���<WV�<X�<<��<l�< �<���<�V�<6�<쇼<��<��<�5�<n��<�C�<�Ƨ<�F�<�Ġ<@�<���<\1�<���<T�<���<��<�t�<�<8�z<J�s<\rl<Ue<�8^<�W<�P<��H<��A<j�:<��3<ܰ,<;�%<Y�<��<G�<��	<��<���;�;�;*��;&��;�n�;��;���;T=�;���;��};�wc;�uI;]�/;��;�:hy�:P�:E:���9+-62��6�@�u���3�����L�
%��;�i,R��bh�+\~����˔�(l��	�P��h����Ȼ �һ��ܻ{u��!𻹰����=;��
��d�1���U����!��Z%���)��-���1��6��:��>�B���E�y�I���M�fqQ�'3U�S�X�d�\�{@`���c�4sg�x k��n��r��zu�v�x��S|�|�������4���݄�b����&���ǉ�f��^�������4�� ˑ�~_��Q򔼅���8�������.��`���E���Ο�{W��bߢ��f���쥼�r��&���}�����Ѕ���	��Ѝ������������ޝ��j"��3���z,��-���}8���  �  bN=0�M=��L=AL=PK=_�J="�I=A�H=�5H=�mG=��F=��E=NE=�DD=�xC=<�B=��A=wA=�<@=:k?=R�>=�==��<=�<=F?;=be:=�9=ج8=�7=��6=36= '5=�@4=�X3=`n2=�1=[�0=k�/=1�.=v�-=J�,=��+=!�*=�)=*�(=u�'=Ϸ&=2�%=��$=Ƌ#=�v"=�^!=0C =S$==e�=+�=g�=�U=�!=9�=Ю=�o=�,=��=X�=�L=��=��=�J=$�	=��=L&=?�=^P=��=�k=[��<g��<Q��<H��<A��<���<0��<Z��<.o�<�B�<S�<���<��<SV�<`�<8��<l�<�<|��<�V�<8�<���<��<��<�5�<^��< D�<�Ƨ<�F�<�Ġ<@�<���<Z1�<���<M�<���<��<�t�<�<:�z<A�s<9rl<Ue<�8^<�W<�P<��H<��A<\�:<��3<ް,<I�%<d�<}�<A�<��	<��<X��;�;�;��;!��;�n�;���;���;7=�;���;A�};Zwc;#vI;M�/;��;>�:�y�:8P�:�E:���9� 6���˳@������2�������
%��;�o,R�bh�(\~�	��~˔�3l����Q��B����Ȼ2�һتܻpu��!������R;���
��d�#���U�,���!��Z%���)���-���1��6�:��>�B���E�y�I���M�]qQ�(3U�7�X�g�\�w@`��c�Nsg�r k��n��r��zu�h�x��S|�w�������4���݄�o����&���ǉ�f��b�������4��ˑ�s_��P�z���7�������.��o���E���Ο�}W��nߢ��f���쥼�r�����}�����х���	��č������������䝶�h"��*���q,��/���w8���  �  bN=+�M=��L=@L=PK=b�J=!�I=C�H=�5H=�mG=��F=��E=QE=�DD=�xC=3�B=��A={A=�<@==k?=O�>=�==��<=�<=D?;=_e:=�9=֬8=�7=��6=66=�&5=�@4=�X3=cn2=��1=Z�0=n�/='�.=z�-=H�,=��+=&�*=�)=*�(=r�'=ӷ&=4�%=��$=ȋ#=�v"=�^!=0C =Z$==b�=)�=a�= V=�!==�=ͮ=�o=�,=��=\�=�L=��=��=�J=#�	=��=P&=6�=aP=��=�k=d��<f��<N��<9��<J��<���<6��<Y��<#o�<�B�<N�<���<��<XV�<]�<;��<l�<%�<���<{V�<<�<퇼<��<��<�5�<i��<�C�<�Ƨ<�F�<�Ġ<@�<���<Y1�<~��<Z�<���<��<�t�<�<G�z<B�s<Yrl<Ue<�8^<�W<�P<��H<��A<v�:<��3<۰,<B�%<b�<��<=�<��	<��<}��;�;�;<��;3��;�n�;���;~��;c=�;���;e�};�wc;�uI;n�/;��;��:�y�:�O�:�E:���9��6���@�r���U3�����e� 
%�)�;�A,R��bh��[~����˔�l��Q��^����Ȼ'�һӪܻbu��!�ʰ����7;��
��d�)���U����!��Z%���)���-���1��6��:��>�B���E�n�I���M�qqQ�3U�]�X�^�\�x@`��c�<sg�s k��n��r��zu���x��S|�y�������4���݄�f����&���ǉ�f��_�������4���ʑ��_��L򔼅���7�������.��e���E���Ο�W��iߢ��f���쥼�r��)���}�����х���	��׍������������᝶�c"��:���r,��.����8���  �  
bN=(�M=��L=?L=PK=d�J= �I=F�H=�5H=�mG=��F=��E=QE=�DD=�xC=3�B=��A=tA=�<@=?k?=N�>= �==��<=�<=@?;=be:=�9=լ8=�7=��6=:6=�&5=�@4=�X3=`n2=��1=S�0=t�/=)�.=}�-=G�,=��+='�*=�)=0�(=o�'=ӷ&=4�%=��$=ɋ#=�v"=�^!=(C =Z$==g�=0�=`�=V=�!=A�=ͮ=�o=�,=��=]�=�L=��=��=�J=%�	=��=T&=6�=gP=��=�k=a��<`��<\��<9��<Q��<���<=��<X��<'o�<�B�<G�<���<��<]V�<\�<=��<l�<�<���<yV�<L�<�<��<��<�5�<t��<�C�<�Ƨ<�F�<�Ġ<@�<���<c1�<z��<_�<�<��<�t�<�<X�z<(�s<lrl<�Te<�8^<�W<�P<��H<��A<��:<��3<�,<>�%<Y�<��<7�<��	<��<���;�;�; ��;3��;�n�;���;x��;d=�;���;h�};�wc;�uI;��/;��;�:1y�:8P�:E:V��9��6F����@�n����2������
%���;��+R��bh��[~�&��~˔�l��!�P��x����Ȼ&�һ˪ܻWu��!𻩰��/��8;�	�
��d����U���!��Z%���)���-���1��6��:��>�B���E�i�I��M�wqQ�3U�[�X�D�\��@`� �c�Bsg�� k�υn��r��zu���x��S|�|�������4���݄�c����&���ǉ�f��]�������4���ʑ��_��<򔼀���8�������.��Z���E���Ο��W��fߢ��f���쥼�r��.����|�����υ���	��ҍ������������흶�]"��4���q,��)����8���  �  bN=.�M=��L=>L=PK=c�J= �I=E�H=�5H=�mG=��F=��E=PE=�DD=�xC=8�B=��A=uA=�<@==k?=T�>=�==��<=�<=G?;=\e:=�9=׬8=�7=��6=66=�&5=�@4=�X3=bn2=��1=X�0=o�/=)�.=v�-=H�,=��+=#�*=
�)='�(=t�'=շ&=4�%=��$=ʋ#=�v"=�^!=.C =X$==d�=*�=c�=�U=�!==�=ή=�o=�,=��=^�=�L=��=��=�J=%�	=��=M&=7�=aP=��=�k=c��<i��<R��<9��<G��<���<6��<X��<$o�<�B�<T�<���<��<UV�<g�<:��<l�<�<���<�V�<;�<�<��<��<�5�<i��<�C�<�Ƨ<�F�<�Ġ<@�<���<S1�<���<T�<���<��<�t�<�<M�z<6�s<`rl< Ue<�8^<�W<�P<��H<��A<k�:<��3<ΰ,<;�%<n�<��<7�<��	<��<q��;�;�;��;1��;�n�;���;���;R=�;���;y�};�wc;CvI;P�/;��;��:z�:�O�:�E:!��9�h6���
�@�����3��J��z�!
%�P�;�2,R��bh� \~���v˔�$l����%Q��K����Ȼ"�һ֪ܻMu��!�Ѱ����@;��
��d�%���U����!��Z%���)���-���1��6��:��>�'B���E�w�I��M�mqQ�$3U�Y�X�[�\�@`��c�=sg�n k��n��r��zu�w�x��S|�|�������4��݄�e����&���ǉ�f��`�������4��ˑ�{_��L�}���7�������.��e���E���Ο��W��fߢ�}f���쥼�r�� ���}�����҅���	��э������������蝶�`"��4���w,��.���x8���  �   bN=3�M=��L=AL=PK=`�J=&�I=?�H=�5H=�mG=��F=��E=NE=�DD=�xC=:�B=��A=yA=�<@=:k?=R�>=�==��<=�<=F?;=]e:=�9=ڬ8=�7=��6=16='5=�@4=�X3=cn2=��1=]�0=j�/=.�.=w�-=G�,=��+= �*=�)=%�(=x�'=η&=6�%=��$=Ƌ#=�v"=�^!=2C =S$==c�=)�=f�=�U=�!=:�=ή=�o=�,=��=V�=�L=��=��=�J="�	=��=L&==�=\P=��=�k=a��<i��<J��<G��<?��<���<.��<\��<'o�<�B�<W�<���<���<OV�<b�<6��<l�<#�<|��<�V�<6�<���<��<��<�5�<d��<�C�<�Ƨ<�F�<�Ġ<@�<���<O1�<���<J�<���<��<�t�<�<:�z<J�s<Arl<Ue<�8^<�W<�P<��H<��A<W�:<Ⱥ3<ɰ,<H�%<]�<��<P�<��	<��<`��;�;�;��;��;�n�;}��;���;0=�;���;r�};bwc;1vI;	�/;	�;.�:�y�:�O�:�E:���9�< 6M��6�@�����z3��{��j�g
%� �;��,R�Nbh�\~�'��˔�8l����6Q��.����Ȼ�һ֪ܻtu��!������R;���
��d�)���U�.���!��Z%���)���-���1��6�:��>�,B���E�}�I���M�nqQ�(3U�@�X�o�\�o@`��c�Asg�m k��n��r��zu�s�x��S|�s�������4��}݄�s����&���ǉ�f��d�������4��ˑ�u_��Q�{���9�������.��j���E���Ο�zW��hߢ��f���쥼�r�����}�����؅���	��ύ������������ߝ��g"��5���m,��6���v8���  �  bN=,�M=��L=DL=PK=a�J="�I=D�H=�5H=�mG=��F=��E=QE=�DD=�xC=5�B=��A=wA=�<@==k?=Q�>=�==��<=�<=C?;=de:=�9=֬8=�7=��6=46=�&5=�@4=�X3=bn2=��1=Z�0=o�/=*�.=z�-=H�,=��+=#�*=�)=,�(=v�'=η&=4�%=��$=ɋ#=�v"=�^!=+C =X$==e�=,�=b�=�U=�!=;�=ή=�o=�,=��=W�=�L=��=��=�J=&�	=��=P&=9�=bP=��=�k=a��<f��<Q��<?��<D��<���<8��<Z��<&o�<�B�<P�<���<��<UV�<c�<9��<l�<�<���<V�<A�<�<��<��<�5�<m��<�C�<�Ƨ<�F�<�Ġ<	@�<���<Y1�<���<S�<��<��<�t�<�<J�z<A�s<Mrl<Ue<�8^<�W<�P<��H<��A<m�:<��3<ְ,<S�%<S�<��<?�<��	<��<���;�;�;"��;3��;�n�;���;���;W=�;���;A�};�wc;!vI;P�/;��;z�:�y�:�P�:�E:���9�6�����@�@���'3�����w�D
%�/�;�2,R��bh��[~���g˔�#l��
�P��>����Ȼ%�һ�ܻVu��!�ϰ��"��>;� �
��d����U����!��Z%���)���-���1��6�:��>�B���E�t�I��M�iqQ�3U�P�X�Z�\�z@`��c�Bsg�s k��n��r��zu�t�x��S|�x�������4���݄�n����&���ǉ�f��a�������4��ˑ�_��G����4�������.��a���E���Ο��W��hߢ��f���쥼�r��%���}�����ԅ���	��ԍ������������❶�a"��7���r,��3���v8���  �  bN=,�M=��L=>L=PK=h�J=�I=I�H=�5H=�mG=��F=��E=QE=�DD=�xC=1�B=��A=vA=�<@=>k?=N�>="�==��<=�<=@?;=ae:=�9=׬8=�7=��6=:6=�&5=�@4=�X3=bn2=��1=U�0=q�/=%�.={�-=I�,=��+=&�*=�)=,�(=o�'=շ&=4�%=��$=̋#=�v"=�^!=+C =^$==d�=,�=^�=V=�!=B�=ʮ=�o=�,=��=_�=�L=��=��=�J=#�	=��=S&=3�=dP=��=�k=e��<d��<U��<4��<O��<���<6��<[��<%o�<�B�<F�<��<��<_V�<^�<9��<l�<�<���<uV�<E�<<��<��<�5�<u��<�C�<�Ƨ<�F�<�Ġ<@�<���<[1�<���<Z�<���<��<�t�<	�<R�z<-�s<trl<�Te<�8^<�W<�P<��H<��A<v�:<��3<۰,<;�%<[�<��<+�<��	<��<���;�;�;)��;7��;�n�;���;k��;s=�;���;��};�wc;�uI;��/;\�;��:;y�:P�:�E:��9a�6	���@������2�����|��	%�t�;�,R��bh��[~����˔�	l���P��z����Ȼ"�һ٪ܻ>u�"𻢰��$��);��
��d����U����!��Z%���)���-���1��6��:��>�B���E�i�I���M�lqQ�3U�g�X�Q�\��@`���c�9sg�x k�܅n��r��zu���x��S|�u�������4���݄�[����&���ǉ�f��a�������4���ʑ��_��B򔼃���8�������.��X��� E���Ο��W��`ߢ��f���쥼�r��&���}�����̅���	��֍������������띶�_"��7���w,��)����8���  �  bN=-�M=��L=AL=PK=d�J=�I=F�H=�5H=�mG=��F=��E=OE=�DD=�xC=8�B=��A=tA=�<@==k?=N�>=�==��<=�<=B?;=be:=�9=ج8=�7=��6=46=�&5=�@4=�X3=_n2=��1=V�0=p�/=.�.=x�-=H�,=��+=$�*=
�)=+�(=r�'=Ϸ&=3�%=��$=ɋ#=�v"=�^!=+C =V$==e�=,�=d�=�U=�!=>�=̮=�o=�,=��=Y�=�L=��=��=�J=#�	=��=P&=<�=cP=��=�k=]��<f��<W��<B��<G��<���<3��<\��<#o�<�B�<L�<���<��<\V�<]�<:��<l�<�<���<�V�<@�<���<��<	��<�5�<n��<�C�<�Ƨ<�F�<�Ġ<@�<���<V1�<���<W�<���<��<�t�<�<Q�z</�s<Url<�Te<�8^<�W<�P<��H<��A<l�:<��3<հ,<H�%<]�<��<3�<��	<��<���;�;�;��;(��;�n�;���;���;H=�;���;v�};�wc;�uI;��/;y�;��:sy�:4P�:�E:���9
6K��w�@�����2��}���M
%�e�;�,R�Obh��[~����˔�l����Q��Z����Ȼ,�һ֪ܻVu��!𻿰��%��F;��
��d����U���!��Z%���)���-���1��6�
:��>�B���E�s�I���M�jqQ�3U�F�X�T�\��@`��c�Isg�t k�څn��r��zu�~�x��S|�t�������4���݄�h����&���ǉ�f��`�������4��ˑ�z_��G�|���7�������.��`���E���Ο��W��fߢ��f���쥼�r��$���}�����Ӆ���	��ɍ������������띶�_"��-���r,��0���8���  �  bN=.�M=��L=BL=PK=e�J=#�I=@�H=�5H=�mG=��F=��E=ME=�DD=�xC=8�B=��A=~A=�<@=>k?=R�>=�==��<=�<=E?;=`e:=�9=ڬ8=�7=��6=.6=�&5=�@4=�X3=cn2=��1=^�0=j�/=+�.=u�-=H�,=��+=!�*=
�)='�(=v�'=ѷ&=9�%=��$=ǋ#=�v"=�^!=3C =W$==`�=&�=d�=�U=�!=:�=Ү=�o=�,=��=Z�=�L=��=��=�J="�	=��=K&=:�=]P=��=�k=d��<l��<I��<C��<<��<���</��<\��<!o�<�B�<R�<���<���<QV�<a�<=��<l�<+�<}��<�V�<1�<�<��<��<�5�<h��<D�<�Ƨ<�F�<�Ġ<@�<���<N1�<���<R�<���<��<�t�<�<@�z<O�s<Frl<Ue<�8^<�W<�P<��H<��A<d�:<��3<Ű,<K�%<b�<��<D�<��	<��<{��;�;�;F��;��;�n�;j��;���;1=�;���;P�};�wc;'vI;!�/;��;��:�y�:	P�:3E:x��9֔ 6���ݴ@�����3��c��a�]
%��;��,R�|bh�;\~����˔�0l����$Q��@����Ȼ��һتܻhu��!������E;��
��d�9���U�%���!��Z%���)���-���1��6�:��>�&B���E�}�I���M�dqQ�-3U�L�X�n�\�k@`��c�<sg�h k���n��r��zu�k�x��S|�s�������4���݄�g����&���ǉ�f��\�������4��
ˑ�x_��V򔼀���9�������.��f���E���Ο��W��`ߢ��f���쥼�r��"���	}�����م���	��э������������ܝ��e"��8���s,��8���x8���  �  bN=0�M=��L=?L=PK=d�J= �I=D�H=�5H=�mG=��F=��E=LE=�DD=�xC=:�B=��A=xA=�<@=>k?=O�>=�==��<=�<=A?;=ae:=�9=۬8=�7=��6=66='5=�@4=�X3=^n2=��1=X�0=o�/=,�.=|�-=I�,=��+=$�*=�)=-�(=p�'=ҷ&=4�%=��$=ǋ#=�v"=�^!=-C =V$==g�=.�=c�=�U=�!=;�=Ϯ=�o=�,=��=\�=�L=��=��=�J=�	=��=R&=;�=cP=��=�k=Z��<g��<S��<E��<K��<���<-��<`��<-o�<�B�<I�<���<��<UV�<^�<<��<l�<�<}��<�V�<B�<���<��<��<�5�<m��<�C�<�Ƨ<�F�<�Ġ<@�<���<[1�<���<T�<���<��<�t�<�<J�z<:�s<Crl<Ue<�8^<�W<�P<��H<��A<g�:<��3<ܰ,<>�%<X�<��<6�<��	<��<���;�;�;$��;��;�n�;���;���;.=�;���;.�};�wc;�uI;Y�/;��;�:Dy�:P�:�E:���9�m 6����@�����3������o
%�F�;�(,R�jbh��[~����˔�l�����P��q�����Ȼ'�һ�ܻlu��!�ٰ����G;��
��d����U�"���!��Z%���)���-���1��6��:��>�B���E�o�I��M�fqQ�3U�G�X�V�\�~@`��c�Psg�r k��n��r��zu�u�x��S|�k�������4���݄�c����&���ǉ�f��^�������4��
ˑ�x_��F�x���=�������.��a���E���Ο��W��eߢ��f���쥼�r�����}�����Ѕ���	��͍������������睶�c"��2���m,��-����8���  �  `bN=��M=c�L=�L=�PK=�J=��I=��H=�6H=enG=}�F=��E=`E=�ED=�yC=q�B=4�A=�A=c>@=�l?=�>=��==Q�<=�<='A;=ig:=�9= �8=]�7=��6=�6=�)5=uC4=^[3=/q2=�1=V�0=��/=\�.=̼-=��,=	�+=��*=��)=��(=Q�'=ͻ&=I�%=��$=�#=){"=c!=�G =�(=�=�=�=<�=�Z=�&=>�=ֳ=�t=�1=�=��=R=��=ߩ=P=L�	=��=l+=D�=hU=��=}p=��<���<���<{��<g��<m��<��<֝�<rw�<�J�<�<���<F��<x]�<9�<���<lr�<4�<a��<\�<}��<猼<��<���<�9�<J®<�G�<�ɧ<�I�<JǠ<rB�<���<43�<��<��<됋<g�<u�<#�<��z<9�s<�pl<�Re<6^<�W<� P<��H<��A<��:<�3<5�,<�%<v�<H�<<�<N�	<��<P��;^%�;�z�;���;U�;�۳;�t�;� �;�ߋ;�f};"8c;z4I;/^/;j�;Cz�:���:���:�C:�Y�9Ws7�|�ù_�A�ۣ���ٿ�>��u�9`%�a<�R�R���h��~�P8������t������=}�������Ȼ��һ{�ܻ����L�S���/���O���
��x�#���i�\��$!�`m%���)���-��1�6�� :�!!>��B�9 F���I���M��Q��@U���X�n�\�GM`�X�c�8g��k���n��r��u���x�;]|�ȿ����19���ᄼM����*��0ˉ��i����������7���͑�;b����������{�������0��J����F��pП�Y���ࢼ�g��#�s��%����}��V��j���^
��B������ޕ�����띶�@"������,�������7���  �  XbN=��M=_�L=�L=�PK=�J=��I=�H=�6H=dnG=��F=��E=WE= FD=�yC=x�B=+�A=�A=e>@=�l?=�>=��==S�<=}<=/A;=cg:=�9=�8=V�7=��6=�6=�)5=sC4=`[3=5q2=�1=[�0=��/=]�.=ļ-=��,=�+=��*=��)=��(=W�'=̻&=H�%=��$=�#=1{"=c!=�G =�(=�= �=��==�=�Z=�&=@�=޳=�t=�1=�=��=%R=��=�=�O=F�	=��=e+=E�=fU=��=~p=��<���<���<y��<W��<p��<��<ܝ�<rw�<�J�<&�<���<J��<]�<G�<���<qr�<6�<P��<\�<���<���<��<s��<:�<I®<�G�<ʧ<�I�<BǠ<yB�<���<.3�<��<��<�<Z�<u�<&�<�z<F�s<�pl<�Re<6^<�W<� P<h�H<��A<��:<��3<(�,<�%<��<1�<J�<\�	<��<I��;�%�;�z�;���;FU�;ܳ;u�;z �;�ߋ;�f};E8c;�4I;j^/;��;}y�:���:���:��C:!]�9v9��ù1�A�����ٿ��t�-`%�<���R���h�b�~�s8����������[��^}������Ȼ��һZ�ܻ}�滷L�F�����P���
��x����i�~���#!�Ym%�۩)���-�p�1�6�� :�!>�B�' F���I���M��Q�AU���X�v�\�4M`�Q�c�$g��k��n��r��u���x�U]|�������<9���ᄼY����*��(ˉ��i����������7���͑�/b������酖���������0��K����F��hП�Y���ࢼ�g��#�s������}��Q��v���m
��?�����ؕ�����᝶�A"������$,�������7���  �  RbN=��M=]�L=�L=�PK=��J=��I=��H=�6H=]nG=��F=��E=WE=FD=�yC={�B=+�A=�A=d>@=�l?=�>=��==W�<=w<=6A;=_g:=�9=�8=Q�7=��6=�6=�)5=sC4=\[3=4q2=��1=^�0=��/=c�.=Ƽ-=��,=�+=��*=��)=��(=Z�'=ʻ&=G�%=��$=�#=.{"=c!=�G =�(=�=�=��=A�=�Z=�&=9�=ڳ=�t=�1=�=�=)R=��=�= P=J�	=Đ=e+=K�=aU=��=zp=��<���<���<���<V��<���<��<��<xw�<�J�<4�<���<Q��<t]�<=�<���<ir�<>�<N��<\�<x��<���<��<x��<	:�<:®<�G�<�ɧ<�I�<;Ǡ<}B�<���<&3�<!��<��<��<]�<
u�<0�<٭z<Q�s<�pl<�Re<�5^<�W<� P<k�H<��A<��:<��3<�,<�%<��< �<R�<D�	<��<��;�%�;�z�;���;\U�;�۳;u�;z �;	��;�f};�7c;�4I;^/;ε;�x�:v��:y��:��C:�_�9�/:��ù,�A�B����ٿ�g�t�t`%��<�ڃR�$�h�?�~�A8����������0���}��h����Ȼ��һm�ܻ ��L����
��P�|�
��x���}i�����#!�vm%��)���-�~�1�6�� :�� >�)B� F���I���M��Q�AU���X���\�1M`�c�c�+g��k��n��r��u�b�x�\]|�������E9���ᄼc���|*��3ˉ��i����������7���͑�+b������煖���������0��Z����F��uП�Y���ࢼ�g��%�s��
����}��@��s���e
��4�����ҕ�����ޝ��K"������,�������7���  �  VbN=��M=`�L=�L=�PK=��J=��I=��H=�6H=dnG=�F=��E=ZE=�ED=�yC=u�B=/�A=�A=b>@=�l?=�>=��==X�<={<=.A;=dg:=�9=�8=U�7=��6=�6=�)5=rC4=^[3=4q2=�1=^�0=��/=^�.=Ƽ-=��,=�+=��*=��)=��(=W�'=˻&=I�%=��$=�#=1{"=c!=�G =�(=�=�=��=?�=�Z=�&=>�=޳=�t=�1=�=��=%R=��=�=�O=H�	=��=f+=F�=dU=��=|p=��<���<���<��<W��<r��<��<ם�<sw�<�J�<&�<���<R��<v]�<C�<���<lr�<7�<X��<\�<{��<���<��<���<�9�<H®<�G�<�ɧ<�I�<?Ǡ<xB�<���<.3�<��<��<���<U�<
u�<$�<�z<Q�s<�pl<�Re<6^<�W<� P<]�H<��A<��:<��3<*�,<
�%<��<)�<T�<H�	<��<J��;l%�;�z�;���;1U�;�۳;�t�;� �;�ߋ;�f};N8c;�4I;^/;ݵ;9y�:���: ��:��C:�[�9�B9���ù]�A�ƣ��ڿ�5�t�H`%��<���R�x�h�E�~�y8����������]��]}�������Ȼ��һ_�ܻ��滵L�P���%��P���
��x� ���i�j���#!�am%�ک)���-�x�1��6�� :�!>�B�% F���I���M��Q�AU���X�}�\�.M`�Z�c�,g��k��n��r��u���x�Q]|�ǿ����;9���ᄼ[���{*��1ˉ��i����������7���͑�4b������񅖼��������0��L����F��qП�Y���ࢼ�g��%�s������}��M��{���e
��@�����ҕ���������F"������,��Ʊ���7���  �  _bN=��M=a�L=�L=�PK=�J=��I=��H=�6H=fnG=��F=��E=XE=�ED=�yC=s�B=/�A=�A=e>@=�l?=�>=��==S�<=�<=-A;=eg:=�9=�8=^�7=��6=�6=�)5=sC4=_[3=2q2=�1=W�0=��/=[�.=ʼ-=��,=�+=��*=��)=��(=S�'=ϻ&=G�%=��$=�#=){"=c!=�G =�(=�=!�=��=:�=�Z=�&=C�=׳=�t=�1=�=��=!R=��=�=P=K�	=��=k+=C�=hU=��=|p=��<���<���<w��<d��<n��<���<ٝ�<qw�<�J�<!�<���<G��<y]�<=�<���<rr�<.�<X��<	\�<���<�<��<z��<�9�<O®<�G�<�ɧ<�I�<BǠ<{B�<���<33�<
��<��<�<\�<	u�<!�<��z<3�s<�pl<�Re<6^<~W<� P<t�H<��A<��:<��3</�,<�%<��<5�<I�<S�	<��<Y��;o%�;�z�;���;)U�;:ܳ;�t�;� �;�ߋ;�f};,8c;�4I;;^/;��;�y�:c��:2��:��C:J[�9%7���ù��A�1����ٿ����t�F`%�P<�M�R���h��~�z8������x���y��;}��������Ȼ��һf�ܻ����L�(���,��P���
��x����i�i���#!�Pm%���)���-�w�1�6�� :�!>� B�5 F���I���M��Q��@U���X�k�\�BM`�Y�c�0g��k��n��r��u���x�6]|�Ŀ����79���ᄼQ����*��.ˉ��i����������7���͑�9b���������������0��E����F��mП�Y���ࢼ�g��)�s��!����}��P��u���e
��C������╳����띶�="�����,�������7���  �  UbN=��M=a�L=�L=�PK=��J=��I=�H=�6H=enG=��F=��E=\E=�ED=�yC=r�B=1�A=�A=h>@=�l?=�>=��==T�<=|<=2A;=`g:=�9=�8=S�7=��6=�6=�)5=uC4=[[3=1q2=�1=X�0=��/=^�.=ȼ-=��,=�+=��*=��)=��(=U�'=λ&=H�%=��$=
�#=,{"=c!=�G =�(=�=�=�=<�=�Z=�&=@�=ٳ=�t=�1=�=��=#R=��=�=�O=F�	=��=h+=F�=fU=��=}p=��<���<���<���<_��<o��<��<ܝ�<vw�<�J�<*�<���<L��<|]�<A�<���<tr�<8�<Z��<	\�<{��<팼<��<|��<:�<L®<�G�<ʧ<�I�<@Ǡ<�B�<���<03�<��<��<<_�<	u�<*�<�z<;�s<�pl<�Re<6^<�W<� P<t�H<��A<��:<��3<.�,<��%<��<,�<D�<\�	<��<P��;�%�;�z�;���;U�;�۳;�t�;� �;�ߋ;%g};8c;�4I;Y^/;��;\y�:���:���:@�C:�\�9��9�>�ùa�A������ٿ�����t�1`%�A<���R�x�h�!�~�e8����������_��c}��������Ȼ��һb�ܻ����L�A�����P���
��x�$���i�k���#!�Xm%��)���-�s�1�6�� :�
!>�B�) F���I���M��Q�AU���X�w�\�CM`�X�c�1g�k��n��r���u���x�\]|�������A9���ᄼY����*��+ˉ��i����������7���͑�9b������􅖼��������0��H����F��iП�Y���ࢼ�g��)�s������}��S��r���f
��;�����ݕ�����靶�E"������,�������7���  �  VbN=��M=^�L=�L=�PK=��J=��I=��H=�6H=bnG=��F=��E=[E=�ED=�yC=w�B=/�A=�A=c>@=�l?=�>=��==Y�<=y<=2A;=ag:=�9=�8=T�7=��6=�6=�)5=sC4=_[3=4q2=�1=_�0=��/=`�.=ļ-=��,=�+=��*=��)=��(=Y�'=ɻ&=J�%=��$=�#=2{"=c!=�G =�(=�=�=��=A�=�Z=�&=<�=޳=�t=�1=�=��='R=��=�=�O=G�	==d+=H�=cU=��=|p=��<���<���<~��<T��<~��<��<ܝ�<ww�<�J�<.�<���<W��<s]�<C�<���<kr�<5�<V��<\�<���<�<��<z��<�9�<C®<�G�<�ɧ<�I�<CǠ<xB�<���<)3�<��<��<���<[�<u�<'�<�z<O�s<�pl<�Re<6^<�W<� P<f�H<��A<��:<��3<$�,<�%<��<,�<U�<E�	<��<7��;s%�;�z�;���;;U�;�۳;�t�;� �;�ߋ;�f};,8c;�4I;^/;�;�x�:��:���:�C:�\�9�u9�h�ù��A�꣐��ٿ�	���t�S`%��<���R�_�h�j�~�R8����������@��x}��q���#�Ȼ��һg�ܻ��滰L�d�����P��
��x���~i�t���#!�hm%�ة)���-�~�1��6�� :�� >�B� F���I���M��Q�AU���X��\�&M`�[�c�.g��k��n��r��u�i�x�V]|�������B9���ᄼa���v*��4ˉ��i����������7���͑�.b������텖���������0��Q����F��rП�
Y���ࢼ�g��$�s������}��J��u���m
��=�����ӕ���������D"������#,��±���7���  �  \bN=��M=_�L=�L=�PK=�J=��I=��H=�6H=fnG=��F=��E=YE=�ED=�yC=q�B=1�A=�A=f>@=�l?=�>=��==V�<=|<=0A;=eg:=�9=�8=X�7=��6=�6=�)5=tC4=_[3=1q2=ބ1=Z�0=��/=`�.=ȼ-=��,=�+=��*=��)=��(=V�'=ʻ&=I�%=��$=�#=+{"=c!=�G =�(=�=�=��=:�=�Z=�&=A�=س=�t=�1=�=��=#R=��=�=P=I�	=��=h+=H�=eU=��=yp=��<���<���<���<\��<q��<��<ܝ�<sw�<�J�<'�<���<O��<s]�<>�<���<tr�<4�<[��<\�<���<팼<��<���<:�<K®<�G�<�ɧ<�I�<EǠ<wB�<���<.3�<��<��<�<Z�<u�<+�<�z<@�s<�pl<�Re<6^<�W<� P<n�H<��A<��:<��3<(�,<�%<��<4�<Q�<C�	<��<X��;�%�;�z�;���;U�; ܳ;�t�;� �;�ߋ;g};88c;�4I;�]/;õ;ky�:���:A��:��C:0\�9r8�͎ùa�A������ٿ����t��`%�)<���R�W�h�%�~�g8���������h��X}�������Ȼ��һh�ܻ����L�;�����P���
��x����i�j���#!�Um%��)���-�z�1�6�� :�
!>�B�, F���I���M��Q�AU���X�x�\�;M`�h�c�6g��k��n��r� �u���x�H]|�������89���ᄼZ���~*��4ˉ��i����������7���͑�;b������󅖼��������0��I����F��tП�Y���ࢼ�g��#�s������}��Q��v���c
��9�����ە�����睶�@"������,�������7���  �  YbN=��M=b�L=�L=�PK=�J=��I=�H=�6H=fnG=��F=��E=]E=�ED=�yC=o�B=4�A=�A=g>@=�l?=�>=��==R�<=<=/A;=cg:=�9=�8=W�7=��6=�6=�)5=sC4=Z[3=4q2=�1=Y�0=��/=[�.=ȼ-=��,=�+=��*=��)=��(=R�'=л&=F�%=��$=�#=*{"=c!=�G =�(=�=�=��=;�=�Z=�&=D�=ֳ=�t=�1=�=��=!R=��=ߩ= P=F�	=��=i+=D�=fU=��=�p=��<���<���<w��<c��<k��<��<ܝ�<rw�<�J�<#�<���<G��<]�<D�<���<vr�<-�<a��<\�<���<<��<z��<�9�<P®<�G�<ʧ<�I�<BǠ<B�<���<53�<��<��<쐋<^�<u�<#�<�z<C�s<�pl<�Re<�5^<�W<� P<s�H<��A<��:<��3<3�,<��%<��<2�<?�<j�	<��<]��;{%�;�z�;���;U�;ܳ;�t�;� �;�ߋ;g};8c;�4I;w^/;��;�y�:���:��:��C:�\�9�8���ù��A�:����ٿ���t��_%�+<���R���h�%�~�k8����������|��8}��������Ȼ��һm�ܻu���L�'���.��P���
��x����i�a��$!�Jm%���)���-�u�1�6�� :�!>� B�5 F���I���M��Q� AU���X�v�\�BM`�G�c�$g�k��n��r��u���x�O]|�������89���ᄼR����*��(ˉ��i����������7���͑�?b������򅖼��������0��D����F��_П�Y���ࢼ�g��-�s������}��U��s���j
��B�����ڕ�����坶�I"�� ���",�������7���  �  VbN=��M=_�L=�L=�PK= �J=��I=��H=�6H=`nG=��F=��E=YE=�ED=�yC=w�B=/�A=�A=g>@=�l?=�>=��==V�<={<=1A;=ag:=�9=�8=U�7=��6=�6=�)5=vC4=^[3=2q2=ބ1=\�0=��/=`�.=ļ-=��,=�+=��*=��)=��(=U�'=̻&=H�%=��$=�#=,{"=c!=�G =�(=�=�=��=?�=�Z=�&=>�=س=�t=�1=�=��=$R=��=�=�O=G�	==e+=G�=eU=��=yp=��<���<���<z��<Y��<}��<��<ޝ�<tw�<�J�<*�<���<O��<r]�<C�<���<pr�<3�<X��<\�<���<�<��<y��<:�<B®<�G�<�ɧ<�I�<BǠ<B�<���<,3�<��<��<���<`�< u�<,�<�z<K�s<�pl<�Re<6^<�W<� P<p�H<��A<��:<��3<%�,<��%<��</�<M�<I�	<��<*��;�%�;�z�;���;<U�;ܳ;�t�;� �;�ߋ;g};�7c;�4I;	^/;��;Py�:���:���:��C:�]�9�S9��ù��A�����ٿ�4���t��`%��<���R�`�h�a�~�F8����������S��a}�������Ȼ��һz�ܻ����L�Y�����P���
��x����i�q���#!�am%��)���-���1�6�� :�!>�B�# F���I���M��Q�AU���X�w�\�/M`�f�c�4g��k���n��r��u�k�x�T]|�������?9���ᄼZ���}*��5ˉ��i����������7���͑�0b������텖���������0��Q����F��pП�Y���ࢼ�g��,�s������}��H��q���n
��8�����Օ�����❶�E"������$,�������7���  �  VbN=��M=\�L=�L=�PK=��J=��I=��H=�6H=cnG=��F=��E=WE= FD=�yC=w�B=+�A=�A=f>@=�l?=�>=��==]�<=w<=2A;=bg:=�9=�8=R�7=��6=�6=�)5=qC4=][3=6q2=݄1=`�0=��/=d�.=¼-=��,=�+=��*=��)=��(=\�'=ǻ&=K�%=��$=�#=3{"=c!=�G =�(=�=�=��=>�=�Z=�&=>�=�=�t=�1=�=}�=*R=��=�=�O=D�	=��=a+=L�=_U=��=yp=��<���<���<���<L��<v��<߽�<۝�<qw�<�J�<0�<���<Z��<q]�<K�<���<qr�<>�<O��<\�<��<���<��<{��<	:�<F®<�G�<�ɧ<�I�<?Ǡ<vB�<Ļ�<&3�<��<��<�<S�<u�</�<ڭz<c�s<�pl<Se<�5^<�W<� P<T�H<��A<��:<��3<�,<�%<��<%�<k�<6�	<��<A��;�%�;�z�;���;CU�;�۳;�t�;z �;��;g};C8c;/5I;�]/;*�;�x�:��:뻓:3�C:�\�9e�9���ù��A�@���&ڿ�F�t��`%��<��R��h���~�l8����������X���}��]���3�Ȼ��һI�ܻ��滢L�[�����P���
��x����i�|���#!�cm%�ѩ)���-�r�1��6�� :�� >�#B�& F���I�ŴM��Q�"AU���X���\�&M`�f�c�&g��k��n��r�"�u�w�x�`]|�������@9���ᄼf���r*��6ˉ��i����������7���͑�0b������셖���������0��N����F��yП��X���ࢼ�g���s������}��N��~���h
��5�����ɕ�����ם��K"������,��˱���7���  �  \bN=��M=a�L=�L=�PK= �J=��I=��H=�6H=cnG=�F=��E=\E=�ED=�yC=t�B=0�A=�A=c>@=�l?=�>=��==W�<=|<=2A;=ag:=�9=�8=Z�7=��6=�6=�)5=oC4=[[3=6q2=�1=]�0=��/=`�.=Ǽ-=��,=
�+=��*=��)=��(=U�'=̻&=H�%=��$=�#=+{"=c!=�G =�(=�= �=��=>�=�Z=�&==�=س=�t=�1=�=��=$R=��=�=P=L�	==g+=H�=aU=��=~p=��<���<���<���<[��<{��<��<ޝ�<uw�<�J�<,�<���<P��<v]�<>�<���<lr�<1�<Z��<\�<���<���<��<z��<�9�<F®<�G�<�ɧ<�I�<@Ǡ<}B�<���<13�<��<��<���<_�<u�<'�<حz<U�s<�pl<�Re<�5^<�W<� P<n�H<��A<��:<��3<.�,< �%<��<.�<Q�<O�	<��<?��;m%�;�z�;���;;U�;ܳ;�t�;� �;�ߋ;�f};8c;�4I;^/;ʵ;^y�:��:���:��C:�\�9�"8���ù��A�����|ڿ���t�&`%��<�׃R�]�h�/�~�K8������t���n��^}������
�Ȼ��һi�ܻ����L�Z���(��P���
��x����i�k���#!�em%��)���-�|�1�6�� :�!>�B�, F���I���M��Q�AU���X���\�4M`�Q�c�#g��k��n��r��u�o�x�>]|�������=9���ᄼZ���}*��1ˉ��i����������7���͑�7b������ꅖ��������0��N����F��nП�
Y���ࢼ�g��)�s������}��K��r���g
��=�����Е�����ݝ��K"�����,�������7���  �  XbN=��M=g�L=�L=�PK=�J=��I=�H=�6H=jnG=��F=��E=\E=�ED=�yC=q�B=3�A=�A=k>@=�l?=�>=��==P�<=<=0A;=_g:=�9=�8=U�7=��6=�6=�)5=wC4=a[3=.q2=߄1=Y�0=��/=]�.=ż-=��,=�+=��*=��)=��(=M�'=һ&=F�%=��$=�#=*{"=c!=�G =�(=�=�=��=9�=�Z=�&=E�=ٳ=�t=�1=�=��=R=��=�=�O=E�	=��=e+=C�=iU=��=yp=
��<���<���<u��<X��<k��<��<՝�<ww�<�J�<"�<���<C��<]�<C�<���<{r�<-�<a��<\�<���<錼<��<~��<:�<S®<�G�<ʧ<�I�<FǠ<�B�<���<>3�<	��<��<ꐋ<]�< u�<-�<��z<:�s<�pl<�Re<6^<�W<� P<p�H<��A<��:<��3<E�,<�%<��<7�<4�<p�	<��<u��;�%�;�z�;���;U�;ܳ;�t�;� �;�ߋ;Tg};�8c;�4I;�^/;b�;�y�:���:���:��C:�Z�9}39�Y�ù��A�z���kٿ����u��`%�8<�P�R���h�X�~�w8����������x��-}��������Ȼ��һt�ܻu���L����&���O���
��x����i�c���#!�Dm%��)���-�v�1�6�� :�$!>�B�. F���I�´M��Q�AU���X�g�\�>M`�f�c�=g��k���n��r��u���x�R]|�ʿ����>9���ᄼR����*��(ˉ��i����������7���͑�?b������������������0��A����F��`П�Y���ࢼ�g��8�s��#����}��X��t���n
��8������ޕ�����읶�:"������&,�������7���  �  \bN=��M=a�L=�L=�PK= �J=��I=��H=�6H=cnG=�F=��E=\E=�ED=�yC=t�B=0�A=�A=c>@=�l?=�>=��==W�<=|<=2A;=ag:=�9=�8=Z�7=��6=�6=�)5=oC4=[[3=6q2=�1=]�0=��/=`�.=Ǽ-=��,=
�+=��*=��)=��(=U�'=̻&=H�%=��$=�#=+{"=c!=�G =�(=�= �=��=>�=�Z=�&==�=س=�t=�1=�=��=$R=��=�=P=L�	==g+=H�=aU=��=~p=��<���<���<���<[��<{��<��<ޝ�<uw�<�J�<,�<���<P��<v]�<>�<���<lr�<1�<Z��<\�<���<���<��<z��<�9�<F®<�G�<�ɧ<�I�<@Ǡ<}B�<���<13�<��<��<���<_�<u�<'�<حz<U�s<�pl<�Re<�5^<�W<� P<n�H<��A<��:<��3<.�,< �%<��<.�<Q�<O�	<��<?��;m%�;�z�;���;;U�;ܳ;�t�;� �;�ߋ;�f};8c;�4I;^/;ʵ;^y�:��:���:��C:�\�9�"8���ù��A�����|ڿ���t�&`%��<�׃R�]�h�/�~�K8������t���n��^}������
�Ȼ��һi�ܻ����L�Z���(��P���
��x����i�k���#!�em%��)���-�|�1�6�� :�!>�B�, F���I���M��Q�AU���X���\�4M`�Q�c�#g��k��n��r��u�o�x�>]|�������=9���ᄼZ���}*��1ˉ��i����������7���͑�7b������ꅖ��������0��N����F��nП�
Y���ࢼ�g��)�s������}��K��r���g
��=�����Е�����ݝ��K"�����,�������7���  �  VbN=��M=\�L=�L=�PK=��J=��I=��H=�6H=cnG=��F=��E=WE= FD=�yC=w�B=+�A=�A=f>@=�l?=�>=��==]�<=w<=2A;=bg:=�9=�8=R�7=��6=�6=�)5=qC4=][3=6q2=݄1=`�0=��/=d�.=¼-=��,=�+=��*=��)=��(=\�'=ǻ&=K�%=��$=�#=3{"=c!=�G =�(=�=�=��=>�=�Z=�&=>�=�=�t=�1=�=}�=*R=��=�=�O=D�	=��=a+=L�=_U=��=yp=��<���<���<���<L��<v��<߽�<۝�<qw�<�J�<0�<���<Z��<q]�<K�<���<qr�<>�<O��<\�<��<���<��<{��<	:�<F®<�G�<�ɧ<�I�<?Ǡ<vB�<Ļ�<&3�<��<��<�<S�<u�</�<ڭz<c�s<�pl<Se<�5^<�W<� P<T�H<��A<��:<��3<�,<�%<��<%�<k�<6�	<��<A��;�%�;�z�;���;CU�;�۳;�t�;z �;��;g};C8c;/5I;�]/;*�;�x�:��:뻓:3�C:�\�9��9���ù��A�@���&ڿ�F�t��`%��<��R��h���~�l8����������X���}��]���3�Ȼ��һI�ܻ��滢L�[�����P���
��x����i�|���#!�cm%�ѩ)���-�r�1��6�� :�� >�#B�& F���I�ŴM��Q�"AU���X���\�&M`�f�c�&g��k��n��r�"�u�w�x�`]|�������@9���ᄼf���r*��6ˉ��i����������7���͑�0b������셖���������0��N����F��yП��X���ࢼ�g���s������}��N��~���h
��5�����ɕ�����ם��K"������,��˱���7���  �  VbN=��M=_�L=�L=�PK= �J=��I=��H=�6H=`nG=��F=��E=YE=�ED=�yC=w�B=/�A=�A=g>@=�l?=�>=��==V�<={<=1A;=ag:=�9=�8=U�7=��6=�6=�)5=vC4=^[3=2q2=ބ1=\�0=��/=`�.=ļ-=��,=�+=��*=��)=��(=U�'=̻&=H�%=��$=�#=,{"=c!=�G =�(=�=�=��=?�=�Z=�&=>�=س=�t=�1=�=��=$R=��=�=�O=G�	==e+=G�=eU=��=yp=��<���<���<z��<Y��<}��<��<ޝ�<tw�<�J�<*�<���<O��<r]�<C�<���<pr�<3�<X��<\�<���<�<��<y��<:�<B®<�G�<�ɧ<�I�<BǠ<B�<���<,3�<��<��<���<`�< u�<,�<�z<K�s<�pl<�Re<6^<�W<� P<p�H<��A<��:<��3<%�,<��%<��</�<M�<I�	<��<*��;�%�;�z�;���;<U�;ܳ;�t�;� �;�ߋ;g};�7c;�4I;	^/;��;Py�:���:���:��C:�]�9.T9��ù��A�����ٿ�4���t��`%��<���R�`�h�a�~�F8����������S��a}�������Ȼ��һz�ܻ����L�Y�����P���
��x����i�q���#!�am%��)���-���1�6�� :�!>�B�# F���I���M��Q�AU���X�w�\�/M`�f�c�4g��k���n��r��u�k�x�T]|�������?9���ᄼZ���}*��5ˉ��i����������7���͑�0b������텖���������0��Q����F��pП�Y���ࢼ�g��,�s������}��H��q���n
��8�����Օ�����❶�E"������$,�������7���  �  YbN=��M=b�L=�L=�PK=�J=��I=�H=�6H=fnG=��F=��E=]E=�ED=�yC=o�B=4�A=�A=g>@=�l?=�>=��==R�<=<=/A;=cg:=�9=�8=W�7=��6=�6=�)5=sC4=Z[3=4q2=�1=Y�0=��/=[�.=ȼ-=��,=�+=��*=��)=��(=R�'=л&=F�%=��$=�#=*{"=c!=�G =�(=�=�=��=;�=�Z=�&=D�=ֳ=�t=�1=�=��=!R=��=ߩ= P=F�	=��=i+=D�=fU=��=�p=��<���<���<w��<c��<k��<��<ܝ�<rw�<�J�<#�<���<G��<]�<D�<���<vr�<-�<a��<\�<���<<��<z��<�9�<P®<�G�<ʧ<�I�<BǠ<B�<���<53�<��<��<쐋<^�<u�<#�<�z<C�s<�pl<�Re<�5^<�W<� P<s�H<��A<��:<��3<3�,<��%<��<2�<?�<j�	<��<]��;{%�;�z�;���;U�;ܳ;�t�;� �;�ߋ;g};8c;�4I;w^/;��;�y�:���:��:��C:�\�9`�8���ù��A�:����ٿ���t��_%�+<���R���h�%�~�k8����������|��8}��������Ȼ��һm�ܻu���L�'���.��P���
��x����i�a��$!�Jm%���)���-�u�1�6�� :�!>� B�5 F���I���M��Q� AU���X�v�\�BM`�G�c�$g�k��n��r��u���x�O]|�������89���ᄼR����*��(ˉ��i����������7���͑�?b������򅖼��������0��D����F��_П�Y���ࢼ�g��-�s������}��U��s���j
��B�����ڕ�����坶�I"�� ���",�������7���  �  \bN=��M=_�L=�L=�PK=�J=��I=��H=�6H=fnG=��F=��E=YE=�ED=�yC=q�B=1�A=�A=f>@=�l?=�>=��==V�<=|<=0A;=eg:=�9=�8=X�7=��6=�6=�)5=tC4=_[3=1q2=ބ1=Z�0=��/=`�.=ȼ-=��,=�+=��*=��)=��(=V�'=ʻ&=I�%=��$=�#=+{"=c!=�G =�(=�=�=��=:�=�Z=�&=A�=س=�t=�1=�=��=#R=��=�=P=I�	=��=h+=H�=eU=��=yp=��<���<���<���<\��<q��<��<ܝ�<sw�<�J�<'�<���<O��<s]�<>�<���<tr�<4�<[��<\�<���<팼<��<���<:�<K®<�G�<�ɧ<�I�<EǠ<wB�<���<.3�<��<��<�<Z�<u�<+�<�z<@�s<�pl<�Re<6^<�W<� P<n�H<��A<��:<��3<(�,<�%<��<4�<Q�<C�	<��<X��;�%�;�z�;���;U�; ܳ;�t�;� �;�ߋ;g};88c;�4I;�]/;µ;ky�:���:A��:��C:/\�9pr8�Ύùb�A������ٿ����t��`%�)<���R�W�h�%�~�g8���������h��X}�������Ȼ��һh�ܻ����L�;�����P���
��x����i�j���#!�Um%��)���-�z�1�6�� :�
!>�B�, F���I���M��Q�AU���X�x�\�;M`�h�c�6g��k��n��r� �u���x�H]|�������89���ᄼZ���}*��4ˉ��i����������7���͑�;b������󅖼��������0��I����F��tП�Y���ࢼ�g��#�s������}��Q��v���c
��9�����ە�����睶�@"������,�������7���  �  VbN=��M=^�L=�L=�PK=��J=��I=��H=�6H=bnG=��F=��E=[E=�ED=�yC=w�B=/�A=�A=c>@=�l?=�>=��==Y�<=y<=2A;=ag:=�9=�8=T�7=��6=�6=�)5=sC4=_[3=4q2=�1=_�0=��/=`�.=ļ-=��,=�+=��*=��)=��(=Y�'=ɻ&=J�%=��$=�#=2{"=c!=�G =�(=�=�=��=A�=�Z=�&=<�=޳=�t=�1=�=��='R=��=�=�O=G�	==d+=H�=cU=��=|p=��<���<���<~��<T��<~��<��<ܝ�<ww�<�J�<.�<���<W��<s]�<C�<���<kr�<5�<V��<\�<���<�<��<z��<�9�<C®<�G�<�ɧ<�I�<CǠ<xB�<���<)3�<��<��<���<[�<u�<'�<�z<O�s<�pl<�Re<6^<�W<� P<f�H<��A<��:<��3<$�,<�%<��<,�<U�<E�	<��<7��;s%�;�z�;���;;U�;�۳;�t�;� �;�ߋ;�f};,8c;�4I;^/;�;�x�:��:���:�C:�\�9�v9�i�ù��A�꣐��ٿ�	���t�T`%��<���R�`�h�j�~�R8����������@��x}��q���#�Ȼ��һg�ܻ��滰L�d�����P��
��x���~i�t���#!�hm%�ة)���-�~�1��6�� :�� >�B� F���I���M��Q�AU���X��\�&M`�[�c�.g��k��n��r��u�i�x�V]|�������B9���ᄼa���v*��4ˉ��i����������7���͑�.b������텖���������0��Q����F��rП�
Y���ࢼ�g��$�s������}��J��u���m
��=�����ӕ���������D"������#,��±���7���  �  UbN=��M=a�L=�L=�PK=��J=��I=�H=�6H=enG=��F=��E=\E=�ED=�yC=r�B=1�A=�A=h>@=�l?=�>=��==T�<=|<=2A;=`g:=�9=�8=S�7=��6=�6=�)5=uC4=[[3=1q2=�1=X�0=��/=^�.=ȼ-=��,=�+=��*=��)=��(=U�'=λ&=H�%=��$=
�#=,{"=c!=�G =�(=�=�=�=<�=�Z=�&=@�=ٳ=�t=�1=�=��=#R=��=�=�O=F�	=��=h+=F�=fU=��=}p=��<���<���<���<_��<o��<��<ܝ�<vw�<�J�<*�<���<L��<|]�<A�<���<tr�<8�<Z��<	\�<{��<팼<��<|��<:�<L®<�G�<ʧ<�I�<@Ǡ<�B�<���<03�<��<��<<_�<	u�<*�<�z<;�s<�pl<�Re<6^<�W<� P<t�H<��A<��:<��3<.�,<��%<��<,�<D�<\�	<��<P��;�%�;�z�;���;U�;�۳;�t�;� �;�ߋ;%g};8c;�4I;Y^/;��;\y�:���:���:?�C:�\�9�9�?�ùa�A������ٿ�����t�1`%�A<���R�x�h�!�~�e8����������_��c}��������Ȼ��һb�ܻ����L�A�����P���
��x�$���i�k���#!�Xm%��)���-�s�1�6�� :�
!>�B�) F���I���M��Q�AU���X�w�\�CM`�X�c�1g�k��n��r���u���x�\]|�������A9���ᄼY����*��+ˉ��i����������7���͑�9b������􅖼��������0��H����F��iП�Y���ࢼ�g��)�s������}��S��r���f
��;�����ݕ�����靶�E"������,�������7���  �  _bN=��M=a�L=�L=�PK=�J=��I=��H=�6H=fnG=��F=��E=XE=�ED=�yC=s�B=/�A=�A=e>@=�l?=�>=��==S�<=�<=-A;=eg:=�9=�8=^�7=��6=�6=�)5=sC4=_[3=2q2=�1=W�0=��/=[�.=ʼ-=��,=�+=��*=��)=��(=S�'=ϻ&=G�%=��$=�#=){"=c!=�G =�(=�=!�=��=:�=�Z=�&=C�=׳=�t=�1=�=��=!R=��=�=P=K�	=��=k+=C�=hU=��=|p=��<���<���<w��<d��<n��<���<ٝ�<qw�<�J�<!�<���<G��<y]�<=�<���<rr�<.�<X��<	\�<���<�<��<z��<�9�<O®<�G�<�ɧ<�I�<BǠ<{B�<���<33�<
��<��<�<\�<	u�<!�<��z<3�s<�pl<�Re<6^<~W<� P<t�H<��A<��:<��3</�,<�%<��<5�<I�<S�	<��<Y��;o%�;�z�;���;)U�;:ܳ;�t�;� �;�ߋ;�f};,8c;�4I;;^/;��;�y�:c��:2��:��C:I[�9p%7���ù��A�1����ٿ����t�F`%�P<�M�R���h��~�z8������x���y��;}��������Ȼ��һf�ܻ����L�(���,��P���
��x����i�i���#!�Pm%���)���-�w�1�6�� :�!>� B�5 F���I���M��Q��@U���X�k�\�BM`�Y�c�0g��k��n��r��u���x�6]|�Ŀ����79���ᄼQ����*��.ˉ��i����������7���͑�9b���������������0��E����F��mП�Y���ࢼ�g��)�s��!����}��P��u���e
��C������╳����띶�="�����,�������7���  �  VbN=��M=`�L=�L=�PK=��J=��I=��H=�6H=dnG=�F=��E=ZE=�ED=�yC=u�B=/�A=�A=b>@=�l?=�>=��==X�<={<=.A;=dg:=�9=�8=U�7=��6=�6=�)5=rC4=^[3=4q2=�1=^�0=��/=^�.=Ƽ-=��,=�+=��*=��)=��(=W�'=˻&=I�%=��$=�#=1{"=c!=�G =�(=�=�=��=?�=�Z=�&=>�=޳=�t=�1=�=��=%R=��=�=�O=H�	=��=f+=F�=dU=��=|p=��<���<���<��<W��<r��<��<ם�<sw�<�J�<&�<���<R��<v]�<C�<���<lr�<7�<X��<\�<{��<���<��<���<�9�<H®<�G�<�ɧ<�I�<?Ǡ<xB�<���<.3�<��<��<���<U�<
u�<$�<�z<Q�s<�pl<�Re<6^<�W<� P<]�H<��A<��:<��3<*�,<
�%<��<)�<T�<H�	<��<J��;l%�;�z�;���;1U�;�۳;�t�;� �;�ߋ;�f};N8c;�4I;^/;ݵ;9y�:���: ��:��C:�[�9�B9���ù]�A�ƣ��ڿ�5�t�H`%��<���R�y�h�E�~�y8����������]��]}�������Ȼ��һ_�ܻ��滵L�Q���%��P���
��x� ���i�j���#!�am%�ک)���-�x�1��6�� :�!>�B�% F���I���M��Q�AU���X�}�\�.M`�Z�c�,g��k��n��r��u���x�Q]|�ǿ����;9���ᄼ[���{*��1ˉ��i����������7���͑�4b������񅖼��������0��L����F��qП�Y���ࢼ�g��%�s������}��M��{���e
��@�����ҕ���������F"������,��Ʊ���7���  �  RbN=��M=]�L=�L=�PK=��J=��I=��H=�6H=]nG=��F=��E=WE=FD=�yC={�B=+�A=�A=d>@=�l?=�>=��==W�<=w<=6A;=_g:=�9=�8=Q�7=��6=�6=�)5=sC4=\[3=4q2=��1=^�0=��/=c�.=Ƽ-=��,=�+=��*=��)=��(=Z�'=ʻ&=G�%=��$=�#=.{"=c!=�G =�(=�=�=��=A�=�Z=�&=9�=ڳ=�t=�1=�=�=)R=��=�= P=J�	=Đ=e+=K�=aU=��=zp=��<���<���<���<V��<���<��<��<xw�<�J�<4�<���<Q��<t]�<=�<���<ir�<>�<N��<\�<x��<���<��<x��<	:�<:®<�G�<�ɧ<�I�<;Ǡ<}B�<���<&3�<!��<��<��<]�<
u�<0�<٭z<Q�s<�pl<�Re<�5^<�W<� P<k�H<��A<��:<��3<�,<�%<��< �<R�<D�	<��<��;�%�;�z�;���;\U�;�۳;u�;z �;	��;�f};�7c;�4I;^/;ε;�x�:v��:x��:��C:�_�9�/:��ù,�A�C����ٿ�g�t�t`%��<�ڃR�$�h�?�~�A8����������0���}��h����Ȼ��һm�ܻ ��L����
��P�|�
��x���}i�����#!�vm%��)���-�~�1�6�� :�� >�)B� F���I���M��Q�AU���X���\�1M`�c�c�+g��k��n��r��u�c�x�\]|�������E9���ᄼc���|*��3ˉ��i����������7���͑�+b������煖���������0��Z����F��uП�Y���ࢼ�g��%�s��
����}��@��s���e
��4�����ҕ�����ޝ��K"������,�������7���  �  XbN=��M=_�L=�L=�PK=�J=��I=�H=�6H=dnG=��F=��E=WE= FD=�yC=x�B=+�A=�A=e>@=�l?=�>=��==S�<=}<=/A;=cg:=�9=�8=V�7=��6=�6=�)5=sC4=`[3=5q2=�1=[�0=��/=]�.=ļ-=��,=�+=��*=��)=��(=W�'=̻&=H�%=��$=�#=1{"=c!=�G =�(=�= �=��==�=�Z=�&=@�=޳=�t=�1=�=��=%R=��=�=�O=F�	=��=e+=E�=fU=��=~p=��<���<���<y��<W��<p��<��<ܝ�<rw�<�J�<&�<���<J��<]�<G�<���<qr�<6�<P��<\�<���<���<��<s��<:�<I®<�G�<ʧ<�I�<BǠ<yB�<���<.3�<��<��<�<Z�<u�<&�<�z<F�s<�pl<�Re<6^<�W<� P<h�H<��A<��:<��3<(�,<�%<��<1�<J�<\�	<��<I��;�%�;�z�;���;FU�;ܳ;u�;z �;�ߋ;�f};E8c;�4I;j^/;��;}y�:���:���:��C:!]�9�9��ù1�A�����ٿ��t�-`%�<���R���h�b�~�s8����������[��^}������Ȼ��һZ�ܻ}�滷L�F�����P���
��x����i�~���#!�Ym%�۩)���-�p�1�6�� :�!>�B�' F���I���M��Q�AU���X�v�\�4M`�Q�c�$g��k��n��r��u���x�U]|�������<9���ᄼY����*��(ˉ��i����������7���͑�/b������酖���������0��K����F��hП�Y���ࢼ�g��#�s������}��Q��v���m
��?�����ؕ�����᝶�A"������$,�������7���  �  �bN=1�M=�L=�L=�QK=�J=��I=6�H=�7H=�oG=�F=y�E=E=�GD=�{C=�B=f�A=&A=�@@=Ro?=��>=��==B�<=�<=^D;=�j:=��9=��8=&�7=��6=�6=�-5=�G4=�_3=�u2=��1=Z�0=��/=��.=T�-=X�,=��+=��*=��)=L�(=��'=n�&=�%=��$= �#=d�"=vj!=*O =�0=�=�=��=Q�=c=,/=��=B�=/}=L:=��=�=�Z=�=��=�X=��	=E�=�3=��=�]=�=�x=�  =�	�<q�<��<���<;��<|��<��<M��<[X�<3%�<Y��<���<\i�<��<���<}�<Z$�<��<Ae�<g��<D��<h'�<䵵<�@�<�Ȯ<xM�<zϧ<�N�<�ˠ<}F�<F��<G6�<���<��<���<��<�u�<S�<T�z<��s<Pnl<GOe<�1^<!W<��O<)�H<=�A<ƹ:<\�3<�,<��%<q�<T�<P�<�	<��<���; �;�S�;��;p*�;���;�F�;��;O��;% };s�b;��H;'�.;�B;i��:D��:�Œ:��A:2X�9)�0���ǹ�D�޵���������u���%�0�<�S� Mi��F�M����A��o⟻rd��Ǵ�Z���0ɻ�6ӻ1ݻ��滆��"��N���r������K�_������C!�m�%�x�)���-��2��16��<:�a<>��0B�F���I�A�M���Q�XU�aY�H�\�~b`���c��g�=k���n� r�$�u�Fy�?m|�&��p���R@���脼�����0��8щ�Uo��3�������<���ґ��f��������W��M���4��w����I��1ӟ��[��%㢼j��#𥼦u������>���������6������@������𝶼"�������+������7���  �  �bN=2�M=�L=�L=�QK=�J=��I=9�H=�7H=�oG=�F=x�E=E=�GD=�{C=��B=`�A=(A=�@@=Vo?=��>=��==E�<=�<=gD;=�j:=|�9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=É1=a�0=��/=��.=D�-=V�,=��+=��*=��)=D�(=��'=n�&=�%=��$="�#=i�"=xj!=2O =�0=�=��=�=T�=c=3/=��=G�=2}=Q:=��=�=�Z=�=~�=�X=��	=E�=�3=��=�]=�=�x=�  =�	�<j�<��<z��<G��<p��<��<>��<MX�<E%�<L��<���<di�<��<���<}�<a$�<��<Ie�<K��<@��<e'�<޵�<�@�<�Ȯ<�M�<�ϧ<�N�<�ˠ<�F�<J��<96�<���<��<���<v�<�u�<Q�<Y�z<��s<]nl<oOe<�1^<W<i�O<	�H<]�A<��:<`�3<��,<��%<��<4�<d�<��	<��<	��;j �;�S�;ض�;x*�;���;�F�;��;Z��;� };��b;��H;i�.;�B;g��:m��:�Ē:��A:\V�9�51�4�ǹ�D����:����������%���<�,S�)Mi��G�]����A���⟻{d��^Ǵ�'���0ɻ7ӻݻ���^��"��,���r������m�V������C!�`�%�b�)���-��2��16��<:�?<>��0B�'F���I�I�M���Q�PXU�rY�R�\�cb`���c���g�-k���n�� r�X�u�.y�Xm|�>�����`@��y脼퍆��0��0щ�Mo��(��癩��<���ґ��f��,������Y��S����3��s����I��*ӟ��[��1㢼j�� 𥼵u������R���������R��򎰼���,������ݝ��"�������+�����7���  �  �bN=<�M=�L=�L=�QK=��J=��I=1�H=�7H=�oG=	�F=t�E=E=�GD=�{C=��B=[�A=&A=�@@=Po?=��>=��==J�<=�<=kD;=�j:=��9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=��1=`�0=��/=��.=H�-=]�,=��+=��*=��)=@�(=��'=j�&=�%=��$=�#=h�"=oj!=4O =�0=�=�=��=Y�=c=5/=��=E�=+}=O:=��=�=�Z=�=��=�X=��	=M�=�3=��=�]=�=�x=�  =�	�<k�<��<|��<Z��<g��<��<O��<EX�<N%�<@��<���<Xi�<��<���<}�<`$�<��<^e�<J��<Q��<e'�<ֵ�<�@�<�Ȯ<M�<oϧ<�N�<�ˠ<�F�<F��<76�<���<��<���<}�<�u�<]�<D�z<��s<2nl<jOe<�1^<-W<��O<�H<{�A<��:<��3<��,<�%<��<#�<y�<k�	<��<Ż�;^ �;�S�;ȶ�;�*�;���;�F�;��;P��;r };V�b;��H;��.;�B;���:���:tĒ:S�A:~Y�9�1�c�ǹWD�ᵑ���������%�Ġ<�gS��Li�sG�$����A���⟻"d���Ǵ�%���0ɻ7ӻݻ���j��N"��%���r������^�?������C!���%�k�)���-��2��16��<:�7<>��0B��F���I�D�M���Q�FXU�IY�]�\�gb`���c��g�4k���n�t r�T�u�	y�jm|�(��n���i@��q脼�����0��<щ�To��2�������<���ґ��f��,���󉖼Y��[����3�������I��<ӟ��[��8㢼j��#𥼷u������`��}������E��掰����,������ߝ��"�������+������6���  �  �bN=4�M=�L=�L=�QK=�J=��I=0�H=�7H=�oG=�F=}�E=E=�GD=�{C=��B=^�A=-A=�@@=Vo?=��>=��==K�<=�<=dD;=�j:=��9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=��1=b�0=��/=��.=I�-=X�,=��+=��*=��)=F�(=��'=o�&=�%=��$= �#=p�"=tj!=2O =�0=�=��=�=R�=c=5/=��=M�=2}=Q:=��=�=�Z=�=��=�X=��	=F�=�3=��=�]=�=�x=�  =�	�<f�<��<}��<H��<k��<��<M��<LX�<?%�<L��<���<Yi�<��<���<	}�<i$�<��<Ne�<L��<F��<b'�<浵<�@�<�Ȯ<�M�<qϧ<�N�<�ˠ<�F�<I��<A6�<���<��<���<x�<�u�<J�<K�z<��s<Bnl<wOe<�1^<
W<��O<
�H<Y�A<��:<j�3<�,<��%<��<9�<v�<g�	<��<���;@ �;�S�;˶�;�*�;���;�F�;��;���;c };��b;&�H;��.;
C;~��:"��: Œ:��A:)W�9�D1���ǹgD�c���a����������%���<�pS�8Mi�eG�Q����A���⟻Wd��OǴ�@��y0ɻ�6ӻ�ݻ���$��$"��,���r������k�Z������C!�s�%�I�)���-��2��16��<:�N<>��0B�F���I�K�M���Q�AXU�kY�_�\�^b`���c��g�&k���n�� r�R�u�,y�am|�9��o���a@��脼썆��0��;щ�Go��%�������<���ґ��f��+�������\��K���4��x����I��;ӟ��[��.㢼j��!𥼮u������U���������C���������'������ٝ��"�������+�����7���  �  �bN=.�M=�L=�L=�QK=�J=��I=6�H=�7H=�oG=�F=y�E=E=�GD=�{C=��B=`�A='A=�@@=Ro?=��>=��==C�<=�<=bD;=�j:=��9=��8=$�7=��6=�6=�-5=�G4=�_3=�u2=��1=]�0=��/=��.=N�-=Z�,=��+=��*=��)=K�(=��'=p�&=�%=��$=�#=f�"=uj!=,O =�0=�= �=��=T�=c=-/=��=D�=.}=O:=��=�=�Z=�=�=�X=��	=G�=�3=��=�]=�=�x=�  =�	�<o�<��<���<D��<{��<��<H��<UX�<;%�<R��<���<_i�<��<���<	}�<[$�<��<Le�<V��<G��<e'�<⵵<�@�<�Ȯ<}M�<{ϧ<�N�<�ˠ<�F�<D��<F6�<���<��<���<�<�u�<M�<g�z<��s<Fnl<_Oe<�1^<W<��O<!�H<P�A<��:<R�3<�,<��%<��<8�<a�<��	<��<��;1 �;�S�;ٶ�;�*�;���;�F�;��;P��;` };m�b;��H;;�.;�B;���:���:8Œ:,�A:�U�9`�0���ǹ�D��������_��7���%���<��S�5Mi�G�@����A���⟻�d��#Ǵ�c��u0ɻ"7ӻݻ���u��"��D���r������X�S������C!�r�%�o�)���-��2��16��<:�`<>��0B�$F���I�:�M���Q�,XU�qY�>�\�pb`���c��g�-k���n�� r�9�u�5y�Cm|�;��u���X@���脼獆��0��5щ�So��2�������<���ґ��f��!�������Y��O���4��x����I��0ӟ��[��3㢼j��&𥼨u������C���������B������|��5������坶�"�������+������7���  �  �bN=6�M=�L=�L=�QK=�J=��I=8�H=�7H=�oG=�F=v�E=E=�GD=�{C=��B=`�A=&A=�@@=So?=��>=��==C�<=�<=gD;=�j:=��9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=1=\�0=��/=��.=H�-=Y�,=��+=��*=��)=E�(=��'=r�&=�%=��$= �#=g�"=uj!=3O =�0=�=��=�=V�=c=4/=��=E�=/}=P:=��= �=�Z=�=��=�X=��	=G�=�3=��=�]=�=�x=�  =�	�<n�<��<���<F��<i��<��<L��<DX�<A%�<Q��<���<`i�<��<���<}�<_$�<��<Se�<L��<G��<e'�<ܵ�<�@�<�Ȯ<zM�<ϧ<�N�<�ˠ<�F�<;��<?6�<���<��<���<|�<�u�<X�<O�z<��s<\nl<XOe<�1^<(W<|�O<�H<N�A<��:<r�3<
�,<ؗ%<��<<�<Y�<��	<��<��;j �;�S�;۶�;�*�;���;�F�;��;L��;� };��b;��H;K�.;�B;���:y��:2Ē:s�A:vX�9�U1���ǹ}D���������������%��<�%S� Mi�zG�D����A���⟻Od��RǴ�e��c0ɻ	7ӻݻ���m��"��'���r������h�K������C!�j�%�i�)���-��2��16��<:�Z<>��0B�F���I�U�M���Q�DXU�gY�K�\�ub`���c��g�3k���n�� r�I�u�0y�fm|�-��q���i@��}脼荆��0��4щ�Po��.��癩��<���ґ��f��+�������Y��U����3��z����I��,ӟ��[��0㢼�i��/𥼯u������N���������I��뎰����9������蝶�"�������+�����7���  �  �bN=4�M=�L=�L=�QK=�J=��I=4�H=�7H=�oG=�F=w�E=E=�GD=�{C=��B=]�A=(A=�@@=So?=��>=��==G�<=�<=hD;=�j:=��9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=��1=a�0=��/=��.=E�-=^�,=��+=��*=��)=D�(=��'=n�&=�%=��$=�#=o�"=pj!=1O =�0=�= �=��=V�=c=3/=��=L�=0}=O:=��=�=�Z=�=��=�X=��	=N�=�3=��=�]=�=�x=�  =�	�<g�<��<y��<W��<l��<
��<K��<KX�<G%�<I��<���<Xi�<��<���<}�<`$�<��<Qe�<S��<K��<c'�<ݵ�<�@�<�Ȯ<�M�<xϧ<�N�<�ˠ<�F�<J��<=6�<���<��<���<��<�u�<T�<F�z<��s<Gnl<tOe<�1^<W<x�O<�H<l�A<��:<i�3<�,<�%<��<6�<f�<y�	<��<��;D �;�S�;ζ�;�*�;���;�F�;��;Z��;b };��b;�H;�.;�B;K��:���:�Ē:B�A:�W�9+71�i�ǹ�D�m���?����������%���<�vS��Li��G�����A���⟻Wd��ZǴ�0���0ɻ�6ӻݻ���/��C"��/���r������[�N������C!���%�P�)���-��2��16��<:�C<>��0B�F���I�H�M���Q�QXU�`Y�b�\�cb`���c��g�,k���n�� r�Z�u�y�_m|�4��q���b@��w脼�����0��;щ�Ho��*�������<���ґ��f��$�������[��U���4������I��3ӟ��[��1㢼j�� 𥼱u������R���������L������+������ڝ��"�������+������6���  �  �bN=0�M=�L=�L=�QK=�J=��I=4�H=�7H=�oG=�F={�E=E=�GD=�{C=��B=`�A=)A=�@@=Po?=��>=��==H�<=�<=`D;=�j:=��9=��8= �7=��6=�6=�-5=�G4=�_3=�u2=��1=b�0=��/=��.=K�-=[�,=��+=��*=��)=I�(=��'=k�&=�%=��$=�#=g�"=tj!=/O =�0=�= �=��=Q�=c=1/=��=E�=.}=P:=��=�=�Z=�=��=�X=��	=H�=�3=��=�]=�=�x=�  =�	�<i�<��<���<F��<p��<��<I��<TX�<8%�<K��<���<]i�<��<���<}�<`$�<��<Ge�<Y��<C��<d'�<㵵<�@�<�Ȯ<|M�<uϧ<�N�<�ˠ<vF�<L��<C6�<���<��<���<�<�u�<P�<O�z<��s<5nl<sOe<�1^<W<��O<�H<K�A<��:<\�3<�,< �%<o�<:�<q�<w�	<��<��;E �;�S�;ն�;p*�;ʯ�;�F�;��;f��;� };Y�b;��H;*�.;�B;k��:���:fŒ:/�A:�V�9�
1��ǹ�D�����4������� �%���<�DS��Li�GG�3����A���⟻rd��2Ǵ�K���0ɻ�6ӻݻ���o��#"��8���r������T�^������C!�r�%�k�)���-��2��16��<:�X<>��0B�F���I�O�M���Q�:XU�^Y�W�\�_b`���c��g�,k���n�~ r�I�u�1y�Xm|�2��t���Y@���脼��0��7щ�Ro��3�������<���ґ��f��������Z��N���4��x����I��6ӟ��[��0㢼j��𥼫u������J���������A��򎰼���)������۝��"�������+�����7���  �  �bN=2�M=�L=�L=�QK=�J=��I=;�H=�7H=�oG=�F=u�E=E=�GD=�{C=��B=f�A=$A=�@@=Ro?=��>=��==@�<=�<=cD;=�j:=�9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=��1=_�0=��/=��.=G�-=Y�,=��+=��*=��)=I�(=��'=t�&=�%=��$=&�#=f�"=zj!=-O =�0=�=��=�=S�=c=//=��=D�=5}=N:=��=!�=�Z=�=~�=�X=��	=G�=�3=��=�]=�=�x=�  =�	�<n�<��<���<E��<m��<��<B��<NX�<:%�<U��<���<bi�<��<���<}�<W$�<��<Ie�<P��<@��<m'�<ݵ�<�@�<�Ȯ<yM�<�ϧ<�N�<�ˠ<�F�<B��<C6�<���<��<���<�<�u�<T�<N�z<��s<Nnl<fOe<�1^<#W<r�O<�H<P�A<��:<a�3<
�,<�%<��<>�<Q�<��	<��< ��;N �;�S�;��;v*�;���;�F�;��;>��;� };s�b;��H;v�.;^B;���:���:�Ē:��A:�V�9*'1�~�ǹ�D���������������%�ڠ<�8S�/Mi��G�F����A���⟻zd��2Ǵ�b��W0ɻ7ӻݻ���t���!��>���r������e�X������C!�Z�%�l�)���-��2��16��<:�_<>��0B�%F���I�S�M���Q�EXU�uY�P�\�ib`���c��g�.k���n�� r�H�u�3y�]m|�7��z���_@���脼㍆��0��1щ�Io��0��뤎��<���ґ��f��'������R��U���4��r����I��'ӟ��[��/㢼�i��(𥼬u������L���������M������1������᝶�"�������+�����7���  �  �bN=8�M=�L=�L=�QK=�J=��I=3�H=�7H=�oG=	�F=t�E=E=�GD=�{C=��B=^�A="A=�@@=Oo?=��>=��==G�<=�<=fD;=�j:=��9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=��1=_�0=��/=��.=G�-=`�,=��+=��*=��)=F�(=��'=n�&=�%=��$=�#=g�"=sj!=0O =�0=�=�=��=W�=c=1/=��=D�=0}=L:=��=�=�Z=�=��=�X=��	=P�=�3=��=�]=�=�x=�  =�	�<o�<��<���<Y��<l��<��<M��<OX�<D%�<L��<���<Ui�<��<���<}�<V$�<��<Te�<R��<J��<g'�<ص�<�@�<�Ȯ<�M�<uϧ<�N�<�ˠ<�F�<D��<?6�<���<��<���<��<�u�<_�<G�z<��s<9nl<kOe<�1^<4W<w�O<"�H<s�A<��:<y�3<�,<�%<��<8�<g�<s�	<��<л�;` �;�S�;޶�;�*�;���;�F�;��;0��;� };@�b;��H;��.;�B;���:f��:�Ē:��A:Y�9�c1���ǹ�D�y�����������%�Ӡ<�OS��Li��G�
����A���⟻Hd��LǴ�L���0ɻ�6ӻݻ���l��-"��4���r������U�I������C!�r�%�n�)���-��2��16��<:�P<>��0B�F���I�@�M���Q�EXU�UY�W�\�nb`���c��g�6k���n�� r�K�u�
y�`m|�*��o���_@��{脼퍆��0��?щ�No��5��󤎼�<���ґ��f��$�������W��Y����3������I��6ӟ��[��.㢼 j��&𥼯u������V�����}���M��㎰����.������ߝ��"�������+�������6���  �  �bN=8�M=�L=�L=�QK=�J=��I=,�H=�7H=�oG=
�F={�E=E=�GD=�{C=��B=]�A=-A=�@@=Ro?=��>=��==O�<=�<=fD;=�j:=~�9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=��1=g�0=��/=��.=D�-=Z�,=��+=��*=��)=@�(=��'=j�&=�%=��$=�#=p�"=rj!=6O =�0=�=��=�=T�=c=9/=��=K�=0}=O:=��=�=�Z=�=��=�X=��	=G�=�3=��=�]=�=�x=�  =�	�<a�<��<u��<H��<c��<��<F��<FX�<G%�<@��<���<Ri�<��<���<}�<k$�<��<Pe�<H��<D��<a'�<⵵<�@�<�Ȯ<�M�<iϧ<�N�<�ˠ<}F�<P��<36�<���<��<���<z�<�u�<Q�<<�z<ҍs<5nl<�Oe<�1^<W<��O<	�H<S�A<��:<z�3<�,< �%<��<,�<��<W�	< �<ۻ�;f �;�S�;ƶ�;�*�;z��;�F�;��;���;� };}�b;N�H;��.;MC;��:`��:�Ē:��A:�Y�9m�1���ǹ;D����������������%�V�<��S��Li��G�?����A���⟻Od��yǴ����0ɻ�6ӻ�ݻ���)��5"�����r������l�S������C!�w�%�R�)���-��2��16��<:�5<>��0B�F���I�\�M���Q�UXU�XY�j�\�Pb`���c���g�%k���n�{ r�a�u�,y�rm|�*��w���h@��v脼�����0��Aщ�Eo��+�������<���ґ��f��/������]��O����3��~����I��Bӟ��[��2㢼j��𥼻u������T���������I��򎰼���������Н��"�������+�����
7���  �  �bN=3�M=�L=�L=�QK= �J=��I=3�H=�7H=�oG=�F=v�E=E=�GD=�{C=��B=b�A=&A=�@@=Mo?=��>=��==D�<=�<=gD;=�j:=��9=��8=!�7=��6=�6=�-5=�G4=�_3=�u2=��1=]�0=��/=��.=L�-=]�,=��+=��*=��)=F�(=��'=n�&=�%=��$=!�#=g�"=qj!=,O =�0=�=�=��=V�=c=./=��=C�=0}=L:=��=�=�Z=�=��=�X=��	=J�=�3=��=�]=�=�x=�  =�	�<k�<��<���<K��<t��<��<I��<KX�<H%�<G��<���<Xi�<��<���<}�<[$�<��<Qe�<[��<J��<h'�<ܵ�<�@�<�Ȯ<M�<wϧ<�N�<�ˠ<�F�<H��<>6�<���<��<���<��<�u�<T�<N�z<��s<9nl<_Oe<�1^<W<��O<*�H<Y�A<��:<f�3<�,<�%<��<)�<^�<u�	<��<˻�; �;�S�;��;�*�;ϯ�;�F�;��;K��;8 };+�b;�H;�.;�B; ��:x��:�Ē:>�A:�W�9�0�0�ǹ�D����������A��%��<�>S��Li�;G�#����A���⟻dd��JǴ�2���0ɻ.7ӻ'ݻ���o��<"��C���r������Q�M������C!�~�%�s�)���-��2��16��<:�A<>��0B�F���I�F�M���Q�1XU�^Y�T�\�lb`���c��g�/k���n�� r�;�u�'y�Qm|�-��s���b@��v脼򍆼�0��<щ�Ko��9�������<���ґ��f���������V��V���4�������I��4ӟ��[��;㢼j��!𥼰u������F�����{���C������5������䝶�"�������+������7���  �  �bN=.�M="�L=�L=�QK=�J=��I=>�H=�7H=�oG=�F=y�E=E=�GD=�{C=~�B=a�A='A=�@@=Ro?=��>=��==C�<=�<=eD;=�j:=��9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=ɉ1=Z�0=��/=��.=F�-=X�,=��+=��*=��)=L�(=��'=v�&=�%=��$=&�#=b�"=j!=2O =�0=�=��=�=P�=c=3/=��=A�=4}=S:=��=#�=�Z=�=��=�X=��	=E�=�3=��=�]=�=�x=�  =�	�<t�<��<���<A��<o��<��<M��<JX�<>%�<W��<���<ii�<��<���<!}�<_$�<��<Ae�<S��<7��<b'�<䵵<�@�<�Ȯ<qM�<�ϧ<�N�<�ˠ<�F�<7��<N6�<���<��<���<��<�u�<T�<c�z<��s<tnl<WOe<�1^<"W<d�O<�H<F�A<��:<R�3<$�,<֗%<��<@�<\�<��	<��<��;� �;�S�;ڶ�;I*�;���;~F�;��;U��;};s�b;��H;��.;�B;��:=��:�Ē:y�A:�T�9�1���ǹ[D�6�����������2�%�.�<��S�5Mi��G�P����A���⟻|d��Ǵ�{��B0ɻ�6ӻ�ݻ��滕���!��*���r������g�f������C!�B�%�y�)���-��2��16��<:�c<>��0B�F���I�Q�M���Q�AXU�{Y�D�\�xb`���c��g�0k���n�� r�B�u�;y�Zm|�F��o���b@���脼⍆��0��*щ�Oo��3��ऎ��<���ґ��f��$������]��M����3��k����I��"ӟ��[��.㢼�i��2𥼠u������N���������U���~��;������蝶�"�������+�� ���7���  �  �bN=3�M=�L=�L=�QK= �J=��I=3�H=�7H=�oG=�F=v�E=E=�GD=�{C=��B=b�A=&A=�@@=Mo?=��>=��==D�<=�<=gD;=�j:=��9=��8=!�7=��6=�6=�-5=�G4=�_3=�u2=��1=]�0=��/=��.=L�-=]�,=��+=��*=��)=F�(=��'=n�&=�%=��$=!�#=g�"=qj!=,O =�0=�=�=��=V�=c=./=��=C�=0}=L:=��=�=�Z=�=��=�X=��	=J�=�3=��=�]=�=�x=�  =�	�<k�<��<���<K��<t��<��<I��<KX�<H%�<G��<���<Xi�<��<���<}�<[$�<��<Qe�<[��<J��<h'�<ܵ�<�@�<�Ȯ<M�<wϧ<�N�<�ˠ<�F�<H��<>6�<���<��<���<��<�u�<T�<N�z<��s<9nl<_Oe<�1^<W<��O<*�H<Y�A<��:<f�3<�,<�%<��<)�<^�<u�	<��<˻�; �;�S�;��;�*�;ϯ�;�F�;��;K��;8 };+�b;�H;�.;�B; ��:x��:�Ē:=�A:�W�9�0�0�ǹ�D����������A��%��<�>S��Li�;G�#����A���⟻dd��JǴ�2���0ɻ.7ӻ'ݻ���o��<"��C���r������Q�M������C!�~�%�s�)���-��2��16��<:�A<>��0B�F���I�F�M���Q�1XU�^Y�T�\�lb`���c��g�/k���n�� r�;�u�'y�Qm|�-��s���b@��v脼򍆼�0��<щ�Ko��9�������<���ґ��f���������V��V���4�������I��4ӟ��[��;㢼j��!𥼰u������F�����{���C������5������䝶�"�������+������7���  �  �bN=8�M=�L=�L=�QK=�J=��I=,�H=�7H=�oG=
�F={�E=E=�GD=�{C=��B=]�A=-A=�@@=Ro?=��>=��==O�<=�<=fD;=�j:=~�9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=��1=g�0=��/=��.=D�-=Z�,=��+=��*=��)=@�(=��'=j�&=�%=��$=�#=p�"=rj!=6O =�0=�=��=�=T�=c=9/=��=K�=0}=O:=��=�=�Z=�=��=�X=��	=G�=�3=��=�]=�=�x=�  =�	�<a�<��<u��<H��<c��<��<F��<FX�<G%�<@��<���<Ri�<��<���<}�<k$�<��<Pe�<H��<D��<a'�<⵵<�@�<�Ȯ<�M�<iϧ<�N�<�ˠ<}F�<P��<36�<���<��<���<z�<�u�<Q�<<�z<ҍs<5nl<�Oe<�1^<W<��O<	�H<S�A<��:<z�3<�,< �%<��<,�<��<W�	< �<ۻ�;f �;�S�;ƶ�;�*�;z��;�F�;��;���;� };}�b;N�H;��.;MC;��:`��:�Ē:��A:�Y�9x�1���ǹ;D����������������%�V�<��S��Li��G�?����A���⟻Od��yǴ����0ɻ�6ӻ�ݻ���)��5"�����r������l�S������C!�w�%�R�)���-��2��16��<:�5<>��0B�F���I�\�M���Q�UXU�XY�j�\�Pb`���c���g�%k���n�{ r�a�u�,y�rm|�*��w���h@��v脼�����0��Aщ�Eo��+�������<���ґ��f��/������]��O����3��~����I��Bӟ��[��2㢼j��𥼻u������T���������I��򎰼���������Н��"�������+�����
7���  �  �bN=8�M=�L=�L=�QK=�J=��I=3�H=�7H=�oG=	�F=t�E=E=�GD=�{C=��B=^�A="A=�@@=Oo?=��>=��==G�<=�<=fD;=�j:=��9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=��1=_�0=��/=��.=G�-=`�,=��+=��*=��)=F�(=��'=n�&=�%=��$=�#=g�"=sj!=0O =�0=�=�=��=W�=c=1/=��=D�=0}=L:=��=�=�Z=�=��=�X=��	=P�=�3=��=�]=�=�x=�  =�	�<o�<��<���<Y��<l��<��<M��<OX�<D%�<L��<���<Ui�<��<���<}�<V$�<��<Te�<R��<J��<g'�<ص�<�@�<�Ȯ<�M�<uϧ<�N�<�ˠ<�F�<D��<?6�<���<��<���<��<�u�<_�<G�z<��s<9nl<kOe<�1^<4W<w�O<"�H<s�A<��:<y�3<�,<�%<��<8�<g�<s�	<��<л�;` �;�S�;޶�;�*�;���;�F�;��;0��;� };@�b;��H;��.;�B;���:f��:�Ē:��A:Y�9�c1���ǹ�D�y�����������%�Ӡ<�OS��Li��G�
����A���⟻Hd��LǴ�L���0ɻ�6ӻݻ���l��-"��4���r������U�I������C!�r�%�n�)���-��2��16��<:�P<>��0B�F���I�@�M���Q�EXU�UY�W�\�nb`���c��g�6k���n�� r�K�u�
y�`m|�*��o���_@��{脼퍆��0��?щ�No��5��󤎼�<���ґ��f��$�������W��Y����3������I��6ӟ��[��.㢼 j��&𥼯u������V�����}���M��㎰����.������ߝ��"�������+�������6���  �  �bN=2�M=�L=�L=�QK=�J=��I=;�H=�7H=�oG=�F=u�E=E=�GD=�{C=��B=f�A=$A=�@@=Ro?=��>=��==@�<=�<=cD;=�j:=�9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=��1=_�0=��/=��.=G�-=Y�,=��+=��*=��)=I�(=��'=t�&=�%=��$=&�#=f�"=zj!=-O =�0=�=��=�=S�=c=//=��=D�=5}=N:=��=!�=�Z=�=~�=�X=��	=G�=�3=��=�]=�=�x=�  =�	�<n�<��<���<E��<m��<��<B��<NX�<:%�<U��<���<bi�<��<���<}�<W$�<��<Ie�<P��<@��<m'�<ݵ�<�@�<�Ȯ<yM�<�ϧ<�N�<�ˠ<�F�<B��<B6�<���<��<���<�<�u�<T�<N�z<��s<Nnl<fOe<�1^<#W<r�O<�H<P�A<��:<a�3<
�,<�%<��<>�<Q�<��	<��< ��;N �;�S�;��;v*�;���;�F�;��;>��;� };s�b;��H;v�.;^B;���:���:�Ē:��A:�V�9O'1��ǹ�D���������������%�ڠ<�8S�/Mi��G�F����A���⟻zd��2Ǵ�b��W0ɻ7ӻݻ���t���!��>���r������e�X������C!�Z�%�l�)���-��2��16��<:�_<>��0B�%F���I�S�M���Q�EXU�uY�P�\�ib`���c��g�.k���n�� r�H�u�3y�]m|�7��z���_@���脼㍆��0��1щ�Io��0��뤎��<���ґ��f��'������R��U���4��r����I��'ӟ��[��/㢼�i��(𥼬u������L���������M������1������᝶�"�������+�����7���  �  �bN=0�M=�L=�L=�QK=�J=��I=4�H=�7H=�oG=�F={�E=E=�GD=�{C=��B=`�A=)A=�@@=Po?=��>=��==H�<=�<=`D;=�j:=��9=��8= �7=��6=�6=�-5=�G4=�_3=�u2=��1=b�0=��/=��.=K�-=[�,=��+=��*=��)=I�(=��'=k�&=�%=��$=�#=g�"=tj!=/O =�0=�= �=��=Q�=c=1/=��=E�=.}=P:=��=�=�Z=�=��=�X=��	=H�=�3=��=�]=�=�x=�  =�	�<i�<��<���<F��<p��<��<I��<TX�<8%�<K��<���<]i�<��<���<}�<`$�<��<Ge�<Y��<C��<d'�<㵵<�@�<�Ȯ<|M�<uϧ<�N�<�ˠ<vF�<L��<C6�<���<��<���<�<�u�<P�<O�z<��s<5nl<sOe<�1^<W<��O<�H<L�A<��:<\�3<�,< �%<o�<:�<q�<w�	<��<��;E �;�S�;ն�;p*�;ʯ�;�F�;��;e��;� };Y�b;��H;*�.;�B;k��:���:eŒ:/�A:�V�9�
1��ǹ�D�����4������� �%���<�DS��Li�GG�3����A���⟻rd��2Ǵ�K���0ɻ�6ӻݻ���o��#"��8���r������U�^������C!�r�%�k�)���-��2��16��<:�X<>��0B�F���I�O�M���Q�:XU�^Y�W�\�_b`���c��g�,k���n�~ r�I�u�1y�Xm|�2��t���Y@���脼��0��7щ�Ro��3�������<���ґ��f��������Z��N���4��x����I��6ӟ��[��0㢼j��𥼫u������J���������A��򎰼���)������۝��"�������+�����7���  �  �bN=4�M=�L=�L=�QK=�J=��I=4�H=�7H=�oG=�F=w�E=E=�GD=�{C=��B=]�A=(A=�@@=So?=��>=��==G�<=�<=hD;=�j:=��9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=��1=a�0=��/=��.=E�-=^�,=��+=��*=��)=D�(=��'=n�&=�%=��$=�#=o�"=pj!=1O =�0=�= �=��=V�=c=3/=��=L�=0}=O:=��=�=�Z=�=��=�X=��	=N�=�3=��=�]=�=�x=�  =�	�<g�<��<y��<W��<l��<
��<K��<KX�<G%�<I��<���<Xi�<��<���<}�<`$�<��<Qe�<S��<K��<c'�<ݵ�<�@�<�Ȯ<�M�<xϧ<�N�<�ˠ<�F�<J��<=6�<���<��<���<��<�u�<T�<F�z<��s<Gnl<tOe<�1^<W<x�O<�H<l�A<��:<i�3<�,<�%<��<6�<f�<y�	<��<��;D �;�S�;ζ�;�*�;���;�F�;��;Z��;b };��b;�H;�.;�B;K��:���:�Ē:B�A:�W�9K71�k�ǹ�D�m���?����������%���<�vS��Li��G�����A���⟻Wd��ZǴ�0���0ɻ�6ӻݻ���/��C"��/���r������[�N������C!���%�P�)���-��2��16��<:�C<>��0B�F���I�H�M���Q�QXU�`Y�b�\�cb`���c��g�,k���n�� r�Z�u�y�_m|�4��q���b@��w脼�����0��;щ�Ho��*�������<���ґ��f��$�������[��U���4������I��3ӟ��[��1㢼j�� 𥼱u������R���������L������+������ڝ��"�������+������6���  �  �bN=6�M=�L=�L=�QK=�J=��I=8�H=�7H=�oG=�F=v�E=E=�GD=�{C=��B=`�A=&A=�@@=So?=��>=��==C�<=�<=gD;=�j:=��9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=1=\�0=��/=��.=H�-=Y�,=��+=��*=��)=E�(=��'=r�&=�%=��$= �#=g�"=uj!=3O =�0=�=��=�=V�=c=4/=��=E�=/}=P:=��= �=�Z=�=��=�X=��	=G�=�3=��=�]=�=�x=�  =�	�<n�<��<���<F��<i��<��<L��<DX�<A%�<Q��<���<`i�<��<���<}�<_$�<��<Se�<L��<G��<e'�<ܵ�<�@�<�Ȯ<zM�<ϧ<�N�<�ˠ<�F�<;��<?6�<���<��<���<|�<�u�<X�<O�z<��s<\nl<XOe<�1^<(W<|�O<�H<N�A<��:<r�3<
�,<ؗ%<��<<�<Y�<��	<��<��;j �;�S�;۶�;�*�;���;�F�;��;L��;� };��b;��H;K�.;�B;���:y��:2Ē:s�A:uX�9�U1���ǹ}D���������������%��<�%S� Mi�zG�D����A���⟻Od��RǴ�e��c0ɻ	7ӻݻ���m��"��'���r������h�K������C!�j�%�i�)���-��2��16��<:�Z<>��0B�F���I�U�M���Q�DXU�gY�K�\�ub`���c��g�3k���n�� r�I�u�0y�fm|�-��q���i@��}脼荆��0��4щ�Po��.��癩��<���ґ��f��+�������Y��U����3��z����I��,ӟ��[��0㢼�i��/𥼯u������N���������I��뎰����9������蝶�"�������+�����7���  �  �bN=.�M=�L=�L=�QK=�J=��I=6�H=�7H=�oG=�F=y�E=E=�GD=�{C=��B=`�A='A=�@@=Ro?=��>=��==C�<=�<=bD;=�j:=��9=��8=$�7=��6=�6=�-5=�G4=�_3=�u2=��1=]�0=��/=��.=N�-=Z�,=��+=��*=��)=K�(=��'=p�&=�%=��$=�#=f�"=uj!=,O =�0=�= �=��=T�=c=-/=��=D�=.}=O:=��=�=�Z=�=�=�X=��	=G�=�3=��=�]=�=�x=�  =�	�<o�<��<���<D��<{��<��<H��<UX�<;%�<R��<���<_i�<��<���<	}�<[$�<��<Le�<V��<G��<e'�<⵵<�@�<�Ȯ<}M�<{ϧ<�N�<�ˠ<�F�<D��<F6�<���<��<���<�<�u�<M�<g�z<��s<Fnl<_Oe<�1^<W<��O<!�H<P�A<��:<R�3<�,<��%<��<8�<a�<��	<��<��;1 �;�S�;ٶ�;�*�;���;�F�;��;P��;` };m�b;��H;;�.;�B;���:���:8Œ:+�A:�U�9u�0���ǹ�D��������`��7���%���<��S�5Mi�G�@����A���⟻�d��$Ǵ�c��u0ɻ"7ӻݻ���u��"��D���r������X�S������C!�r�%�o�)���-��2��16��<:�`<>��0B�%F���I�:�M���Q�,XU�qY�>�\�pb`���c��g�-k���n�� r�9�u�5y�Cm|�;��u���X@���脼獆��0��5щ�So��2�������<���ґ��f��!�������Y��O���4��x����I��0ӟ��[��3㢼j��&𥼨u������C���������B������|��5������坶�"�������+������7���  �  �bN=4�M=�L=�L=�QK=�J=��I=0�H=�7H=�oG=�F=}�E=E=�GD=�{C=��B=^�A=-A=�@@=Vo?=��>=��==K�<=�<=dD;=�j:=��9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=��1=b�0=��/=��.=I�-=X�,=��+=��*=��)=F�(=��'=o�&=�%=��$= �#=p�"=tj!=2O =�0=�=��=�=R�=c=5/=��=M�=2}=Q:=��=�=�Z=�=��=�X=��	=F�=�3=��=�]=�=�x=�  =�	�<f�<��<}��<H��<k��<��<M��<LX�<?%�<L��<���<Yi�<��<���<	}�<i$�<��<Ne�<L��<F��<b'�<浵<�@�<�Ȯ<�M�<qϧ<�N�<�ˠ<�F�<I��<A6�<���<��<���<x�<�u�<J�<K�z<��s<Bnl<wOe<�1^<
W<��O<
�H<Y�A<��:<j�3<�,<��%<��<9�<v�<g�	<��<���;@ �;�S�;˶�;�*�;���;�F�;��;���;c };��b;&�H;��.;
C;~��:"��: Œ:��A:(W�9�D1���ǹgD�c���a����������%���<�pS�8Mi�eG�Q����A���⟻Wd��OǴ�@��y0ɻ�6ӻ�ݻ���$��$"��,���r������k�Z������C!�s�%�I�)���-��2��16��<:�N<>��0B�F���I�K�M���Q�AXU�kY�_�\�^b`���c��g�&k���n�� r�R�u�,y�am|�9��o���a@��脼썆��0��;щ�Go��%�������<���ґ��f��+�������\��K���4��x����I��;ӟ��[��.㢼j��!𥼮u������U���������C���������'������ٝ��"�������+�����7���  �  �bN=<�M=�L=�L=�QK=��J=��I=1�H=�7H=�oG=	�F=t�E=E=�GD=�{C=��B=[�A=&A=�@@=Po?=��>=��==J�<=�<=kD;=�j:=��9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=��1=`�0=��/=��.=H�-=]�,=��+=��*=��)=@�(=��'=j�&=�%=��$=�#=h�"=oj!=4O =�0=�=�=��=Y�=c=5/=��=E�=+}=O:=��=�=�Z=�=��=�X=��	=M�=�3=��=�]=�=�x=�  =�	�<k�<��<|��<Z��<g��<��<O��<EX�<N%�<@��<���<Xi�<��<���<}�<`$�<��<^e�<J��<Q��<e'�<ֵ�<�@�<�Ȯ<M�<oϧ<�N�<�ˠ<�F�<F��<76�<���<��<���<}�<�u�<]�<D�z<��s<2nl<jOe<�1^<-W<��O<�H<{�A<��:<��3<��,<�%<��<#�<y�<k�	<��<Ż�;^ �;�S�;ȶ�;�*�;���;�F�;��;P��;r };V�b;��H;��.;�B;���:���:tĒ:S�A:}Y�9
�1�d�ǹWD�ᵑ���������%�Ġ<�gS��Li�sG�$����A���⟻"d���Ǵ�%���0ɻ7ӻݻ���j��O"��%���r������^�?������C!���%�k�)���-��2��16��<:�7<>��0B��F���I�D�M���Q�FXU�IY�]�\�gb`���c��g�4k���n�t r�T�u�
y�jm|�(��n���i@��q脼�����0��<щ�To��2�������<���ґ��f��,���󉖼Y��[����3�������I��<ӟ��[��8㢼j��#𥼷u������`��}������E��掰����,������ߝ��"�������+������6���  �  �bN=2�M=�L=�L=�QK=�J=��I=9�H=�7H=�oG=�F=x�E=E=�GD=�{C=��B=`�A=(A=�@@=Vo?=��>=��==E�<=�<=gD;=�j:=|�9=��8=�7=��6=�6=�-5=�G4=�_3=�u2=É1=a�0=��/=��.=D�-=V�,=��+=��*=��)=D�(=��'=n�&=�%=��$="�#=i�"=xj!=2O =�0=�=��=�=T�=c=3/=��=G�=2}=Q:=��=�=�Z=�=~�=�X=��	=E�=�3=��=�]=�=�x=�  =�	�<j�<��<z��<G��<p��<��<>��<MX�<E%�<L��<���<di�<��<���<}�<a$�<��<Ie�<K��<@��<e'�<޵�<�@�<�Ȯ<�M�<�ϧ<�N�<�ˠ<�F�<J��<96�<���<��<���<v�<�u�<Q�<Y�z<��s<]nl<oOe<�1^<W<i�O<	�H<]�A<��:<`�3<��,<��%<��<4�<d�<��	<��<	��;j �;�S�;ض�;x*�;���;�F�;��;Z��;� };��b;��H;h�.;�B;g��:m��:�Ē:��A:\V�9�51�4�ǹ�D����:����������%���<�,S�)Mi��G�]����A���⟻{d��^Ǵ�'���0ɻ7ӻݻ���^��"��,���r������m�V������C!�`�%�b�)���-��2��16��<:�?<>��0B�'F���I�I�M���Q�PXU�rY�R�\�cb`���c���g�-k���n�� r�X�u�.y�Xm|�>�����`@��y脼퍆��0��0щ�Mo��(��癩��<���ґ��f��,������Y��S����3��s����I��*ӟ��[��1㢼j�� 𥼵u������R���������R��򎰼���,������ݝ��"�������+�����7���  �  �cN=�M=&�L=�L=�RK=u�J=s�I=� I=�9H=�qG="�F=��E=E=gJD=y~C=f�B=o�A=YA=8D@=�r?=W�>=��==\�<=� <=�H;=go:=d�9=��8=f�7=N�6=w6=�35=�M4=Ef3=w|2=��1=c�0=��/=-�.=�-=I�,=�+="�*=��)=#�(=��'=��&=��%=]�$=�#=��"=�t!=�Y =F;=]=�=1�=��=�n=�:=S=�=�=BF=��=,�=�f=�=��=�d=�
=>�=�?=��=i=��=&�=� == �<n!�<�<��<��<���<��<���<-k�<�7�<#��<Ѿ�<z�<�/�<^��<��<�2�<���<9r�<��<�<]2�<7��<�J�<�Ѯ<�U�<1ק<�U�<Ҡ<%L�<1ę<�:�<F��<�"�<Δ�<�<�v�<��<��z<`�s<�jl<mJe<e+^<}W<��O<��H<��A<��:<'�3<��,<�%<B�<��<r�<f�	<Q�<o��;��;��;�}�;���;r�;��;���;�h�;q|;n:b;N/H;�Q.;@�;�C�:#��:�j�:�/?:]��9�^���͹�	G�r7���uº�?�z���&��k=�7�S��j��
���銻����\J��̪��.���r��d�ɻl�ӻ��ݻ�M����I���u��>���=�����G�X����p!��%�*�)�!.��C2��Y6��c:��b>��UB�\>F�9J���M�-�Q��xU�/Y���\��`��d�ڮg�:k���n��9r�`�u��y�؃|����ӟ��^J�������9���ى�]w�����J����C��Bّ�m������������a����8���Ü�N��ן�?_��{梼m����'x������G���N������x������8������!��䝶��!������*�������5���  �  �cN=�M=!�L=�L=�RK=p�J=v�I=� I=�9H=�qG=&�F=��E=�E=cJD=`~C=g�B=t�A=bA=;D@=�r?=V�>=��==a�<=� <=�H;=ko:=b�9=��8=g�7=V�6=o6=�35=�M4=Df3=z|2=��1=g�0=��/=-�.=��-=L�,=�+=�*=��)=�(=��'=��&=��%=_�$=�#=��"=�t!=�Y =J;=e=�=�=��=�n=�:=R=�=�=BF=��=*�=�f=�=��=�d=�
=D�=�?=��=zi=��='�=� =? �<i!�<��<��<��<���<��<���</k�<�7�<��<ܾ�<z�<�/�<]��<���<�2�<���<?r�<��<㠼<p2�<A��<�J�<�Ѯ<�U�<&ק<�U�<Ҡ<,L�<Bę<�:�<C��<�"�<ݔ�<�<�v�<��<z�z<{�s<�jl<�Je<\+^<|W<��O<��H<��A<��:<#�3<o�,<�%<R�<��<~�<R�	<_�<n��;)��;�;�}�;���;Aq�;��;筘;�h�;?q|;Z:b;G/H;IQ.;��;
C�:��:k�:Z/?:`��9TY��I�͹eG�l7���uº�?�M���&��k=�z�S��j��
���銻q���}J��/̪��.���r��f�ɻ`�ӻ�ݻ�M绱��\���]��.���=���H�@����p!��%��)��!.��C2��Y6��c:��b>��UB�k>F�HJ���M��Q��xU�/Y���\��`��d�Үg�
:k���n��9r��u�py�΃|����ڟ��]J�������9���ى�`w�����G����C��=ّ�m��2����������W����8���Ü�N��ן�<_���梼	m����3x������M���>�������������=������!��ٝ���!������*�������5���  �  �cN=�M=�L=�L=�RK=n�J=}�I=� I=�9H=�qG=&�F=��E=�E=lJD=e~C=q�B=k�A=_A=7D@=�r?=Z�>=��==f�<=� <=�H;=ho:=e�9=��8=d�7=U�6=j6=�35=�M4=Bf3=w|2=��1=g�0=��/=6�.=��-=J�,=�+=�*=��)=�(=��'=��&=��%=a�$=�#=��"=�t!=�Y =?;=g=�='�=��=�n=�:=M=�=�=CF=��=%�=�f=�=��=�d=�
=B�=�?=��=xi=��=!�=� == �<i!�<��<��<��<���<��<���<*k�<�7�<��<��<z�<�/�<\��<��<�2�<���<Sr�<��<���<j2�<0��<�J�<�Ѯ<�U�<ק<�U�<Ҡ<)L�<Dę<�:�<S��<�"�<ٔ�<�<�v�<��<g�z<x�s<�jl<�Je<N+^<�W<��O<��H<��A<��:<>�3<j�,<�%<N�<��<��<B�	<n�<N��;&��;��;�}�;���;iq�;Q�;���;�h�;�p|;C:b;�/H;Q.;ڡ;�B�:	��:�j�:50?:��9'u��f�͹�G�s6���uº)@�w��U�&��k=���S�j��
���銻�����J���˪��.��{r����ɻd�ӻބݻ�M绅�𻇅��V��Y���=�����G�)�����o!��%��)��!.��C2��Y6��c:�tb>��UB�P>F�IJ���M��Q��xU��.Y���\��`��d��g�:k���n��9r���u�qy���|����П��aJ���(����9���ى�[w�����Q����C��Rّ� m��$����������h����8���Ü��M��ן�2_���梼m����9x������S���B�����z��㏰�F������2��ڝ���!������*������5���  �  �cN=�M=�L=�L=�RK=r�J=x�I=� I=�9H=�qG=)�F=��E=~E=gJD=h~C=i�B=k�A=eA=8D@=�r?=Y�>=��==`�<=� <=�H;=eo:=_�9=��8=i�7=Q�6=n6=�35=�M4=Df3=z|2=��1=f�0=��/=1�.=��-=H�,=�+=!�*=��)=�(=��'=��&=��%=_�$=�#=��"=�t!=�Y =E;=`=	�=&�=��=�n=�:=N=�=�=BF=��=+�=�f=�=��=�d=�
=@�=�?=��=yi=��=(�=� => �<f!�<��<��<��<���<��<���<&k�<�7�<��<ھ�<z�<�/�<\��<��<�2�<���<Ar�<��<<^2�<<��<�J�<�Ѯ<�U�< ק<�U�<Ҡ<+L�<<ę<�:�<E��<�"�<Ք�<�<�v�<��<t�z<w�s<�jl<�Je<Y+^<�W<��O<��H<��A<��:<(�3<g�,<�%<Q�<��<��<E�	<`�<U��;@��;�;}�;���;~q�;�;���;
i�;q|;V:b;j/H;(Q.;z�;0C�:��:cj�:�.?:$��9�L���͹�G�.7���uº@�H��׸&��k=���S�xj��
���銻����^J��(̪��.���r��e�ɻl�ӻ�ݻ�M绪�𻀅��E��C���=�����G�F�����o!���%� �)��!.��C2��Y6��c:��b>��UB�k>F�<J���M�(�Q��xU��.Y���\��`��d�Ѯg�:k���n��9r���u�y�Ѓ|����ݟ��eJ�������9���ى�\w�����L����C��Mّ�m��#����������\����8���Ü�N��ן�9_��梼
m����8x������F���F��������鏰�@������"��ٝ���!������*������5���  �  �cN=�M=%�L=�L=�RK=p�J=u�I=� I=�9H=�qG=#�F=��E=�E=hJD=g~C=i�B=r�A=`A=7D@=�r?=V�>=��==^�<=� <=�H;=mo:=b�9=��8=j�7=O�6=t6=�35=�M4=Bf3=u|2=��1=b�0=��/=.�.=�-=K�,=�+="�*=~�)=%�(=��'=��&=��%=b�$=�#=��"=�t!=�Y =G;=f=
�=&�=��=�n=�:=Q=�=�=GF=��=+�=�f=�=��=�d=�
=A�=�?=��=}i=��='�=� =7 �<p!�<��<��<��<���<��<���<8k�<�7�<��<Ӿ�<z�<�/�<_��<��<�2�<���<Ar�<��<<m2�<<��<�J�<�Ѯ<�U�<.ק<�U�<Ҡ<(L�<>ę<�:�<8��<�"�<є�<�<�v�<��<|�z<h�s<�jl<mJe<\+^<�W<��O<��H<��A<Ƭ:<�3<��,<�%<G�<��<{�<d�	<[�<o��;��;�;�}�;���;|q�;�;ӭ�;�h�;q|;h:b;;/H;�Q.;X�;�B�:���:ek�:x/?:��9=����͹
G�B7���uºC@���ٸ&��k=�N�S��j��
���銻����WJ��X̪��.���r��g�ɻ��ӻфݻ�M绯��h���h��9���=�����G�:����
p!���%��)��!.��C2��Y6��c:��b>��UB�{>F�9J���M�#�Q��xU�/Y���\�#�`��d��g�:k���n��9r�k�u��y�ƃ|����ܟ��SJ�������9���ى�aw�����L����C��@ّ�m��%����������\����8���Ü�N��	ן�;_���梼m����'x�����E���J������}��쏰�<��������䝶��!������*�������5���  �  �cN=�M=#�L=�L=�RK=p�J=z�I=� I=�9H=�qG=(�F=��E=�E=kJD=e~C=n�B=l�A=`A=9D@=�r?=V�>=��==c�<=� <=�H;=jo:=d�9=��8=g�7=T�6=o6=�35=�M4=Bf3=z|2=��1=g�0=��/=1�.=��-=K�,=�+=!�*=��)=!�(=��'=��&=��%=c�$=�#=��"=�t!=�Y =B;=d=
�=&�=��=�n=�:=P=�=�=GF=��=+�=�f=�=��=�d=�
=B�=�?=��=zi=��=(�=� =; �<i!�<��<��<��<���<��<���</k�<�7�<��<ܾ�<z�<�/�<^��<��<�2�<���<Kr�<��<���<f2�<5��<�J�<�Ѯ<�U�<%ק<�U�<Ҡ<(L�<;ę<�:�<G��<�"�<Ԕ�<�<�v�<��<j�z<|�s<�jl<�Je<Q+^<�W<��O<��H<��A<��:<'�3<z�,<�%<J�<��<��<S�	<[�<f��;9��;��;�}�;���;kq�;7�;���;�h�; q|;]:b;</H;]Q.;��; C�:���:�j�:�/?:���9dY��,�͹pG�{7���uº(@�R��߸&��k=���S�uj��
���銻����bJ��#̪��.���r��f�ɻx�ӻɄݻ�M绣��k���N��P���=�����G�6�����o!���%��)��!.��C2��Y6��c:��b>��UB�g>F�:J���M��Q��xU��.Y���\��`��d�Ԯg�:k���n��9r�~�u�wy�҃|����֟��\J�������9���ى�bw�����L����C��Lّ�	m��%����������c����8���Ü�N��ן�2_���梼m����-x������K���G���������쏰�E������"��ٝ���!������*�������5���  �  �cN=�M=�L=�L=�RK=m�J=y�I=� I=�9H=�qG=)�F=��E=�E=kJD=^~C=n�B=l�A=fA=7D@=�r?=[�>=��==b�<=� <=�H;=jo:=_�9=��8=c�7=U�6=j6=�35=�M4=Bf3=y|2=��1=h�0=��/=8�.=��-=J�,=	�+=�*=��)=�(=��'=��&=��%=`�$=�#=��"=�t!=�Y =C;=e=�="�=��=�n=�:=J=�=�=CF=��='�=�f=�=��=�d=�
=B�=�?=��=vi=��=!�=� =< �<g!�<��<��<��<���<��<���<,k�<�7�<��<۾�<z�<�/�<]��<��<�2�<���<Jr�<��<�<f2�<:��<�J�<�Ѯ<�U�<ק<�U�<Ҡ<+L�<Eę<�:�<G��<�"�<ܔ�<�<�v�<��<g�z<��s<�jl<�Je<K+^<�W<��O<��H<��A<��:<(�3<f�,<�%<V�<��<��<>�	<t�<C��;<��;�;�}�;���;5q�;6�;���;i�;q|;H:b;�/H;Q.;��;�B�:D��:�j�:�.?:��9�{��<�͹�G��6���uº8@�`��j�&��k=���S�j��
���銻����{J��.̪�/��ur��x�ɻ��ӻ�ݻ�M绊�𻝅��?��L���=����H�5�����o!��%��)��!.��C2��Y6��c:�nb>��UB�q>F�FJ���M��Q��xU��.Y���\��`��d�ݮg�:k���n��9r���u�oy�݃|����ޟ��_J���&����9���ى�[w�����R����C��Nّ�
m��2����������^����8���Ü��M��ן�6_���梼
m����8x������T���?��������ߏ��F������7��՝���!������*������5���  �  �cN=�M=!�L=�L=�RK=r�J=y�I=� I=�9H=�qG=%�F=��E=�E=iJD=i~C=l�B=m�A=_A=7D@=�r?=W�>=��==c�<=� <=�H;=io:=b�9=��8=g�7=Q�6=p6=�35=�M4=Bf3={|2=��1=h�0=��/=2�.=��-=J�,=�+="�*=��)= �(=��'=��&=��%=b�$=�#=��"=�t!=�Y =D;=d=�=(�=��=�n=�:=P=�=�=EF=��=*�=�f=�=��=�d=�
=A�=�?=��=wi=��=&�=� =: �<d!�<��<��<��<���<��<���<0k�<�7�<��<ݾ�<	z�<�/�<`��<��<�2�<���<Hr�<��<�<h2�<8��<�J�<�Ѯ<�U�<%ק<�U�<Ҡ<)L�<<ę<�:�<H��<�"�<Д�<�<�v�<��<d�z<��s<�jl<�Je<G+^<�W<��O<��H<��A<��:<+�3<o�,<�%<H�<��<��<P�	<h�<Y��;��;��;�}�;���;�q�;$�;���;�h�;q|;n:b;W/H;MQ.;��;HC�:���:�j�:g/?:B��9*Z����͹G��6��vºG@�=���&��k=���S�fj��
���銻����UJ��,̪��.���r��i�ɻk�ӻτݻ�M绚��q���[��F���=�����G�8�����o!���%��)��!.��C2��Y6��c:��b>��UB�m>F�4J���M�!�Q��xU��.Y���\��`��d�Үg�:k���n��9r�y�u�}y�Ӄ|����ڟ��[J�������9���ى�`w�����M����C��Iّ�m������������`����8���Ü� N��ן�4_��~梼m����2x������I���K������~��돰�H������*��֝���!������*�������5���  �  �cN=�M=!�L=�L=�RK=s�J=s�I=� I=�9H=�qG=(�F=��E=�E=dJD=k~C=g�B=r�A=_A=:D@=�r?=V�>=��==[�<=� <=�H;=io:=a�9=��8=k�7=P�6=q6=�35=�M4=Df3=x|2=��1=d�0=��/=/�.=��-=J�,=�+=%�*=�)= �(=��'=��&=��%=`�$=�#=��"=�t!=�Y =H;=b=�=&�=��=�n=�:=T=�=�=EF=��=/�=�f=�=��=�d=�
=A�=�?=��=}i=��=%�=� => �<o!�<~�<��<��<���<��<���<0k�<�7�<%��<Ͼ�<z�<�/�<`��<���<�2�<���<=r�<��<蠼<h2�<=��<�J�<�Ѯ<�U�<-ק<�U�<Ҡ<0L�<<ę<�:�<=��<�"�<Д�<�<�v�<��<{�z<r�s<�jl<|Je<]+^<�W<��O<��H<��A<ά:<�3<p�,<�%<S�<��<r�<_�	<Y�<��;7��;�;�}�;���;�q�;��;׭�;�h�;6q|;�:b;H/H;wQ.;2�;�C�:¤�:�j�:9/?:r��9S9��؍͹�
G��7���uº�?�j���&��k=�O�S��j��
���銻����BJ��N̪��.���r��D�ɻ��ӻ�ݻ�M绷��M���a��6���=�����G�I����p!��%��)��!.��C2��Y6��c:��b>��UB�z>F�1J���M�$�Q��xU�/Y���\��`��d�خg�:k���n��9r�w�u��y�ƃ|����ݟ��\J�������9���ى�^w�����G����C��@ّ�m������������[����8���Ü�
N��
ן�@_���梼m����2x������?���K���������鏰�<������$��ݝ���!������*�������5���  �  �cN=�M=#�L=�L=�RK=m�J=y�I=� I=�9H=�qG=(�F=��E=�E=jJD=i~C=j�B=p�A=aA=8D@=�r?=X�>=��==a�<=� <=�H;=jo:=c�9=��8=e�7=P�6=n6=�35=�M4==f3=x|2=��1=c�0=��/=6�.=��-=I�,=�+=�*=��)=!�(=��'=��&=��%=a�$=�#=��"=�t!=�Y =B;=f=�=(�=��=�n=�:=N=�=�=EF=��='�=�f=�=��=�d=�
=@�=�?=��=yi=��=&�=� =2 �<k!�<��<��<��<���<��<���<1k�<�7�<��<۾�<z�<�/�<Y��<��<�2�<���<Er�<��<���<j2�<6��<�J�<�Ѯ<�U�<*ק<�U�<Ҡ<"L�<Bę<�:�<A��<�"�<֔�<�<�v�<��<_�z<q�s<�jl<|Je<A+^<�W<��O<��H<��A<��:< �3<z�,<�%<D�<��<��<Y�	<d�<O��;6��;��;�}�;���;�q�;�;ĭ�;�h�;q|;1:b;b/H;rQ.;��;�B�:���:k�:�/?:o��9=h����͹�G��6���uº�@�i����&��k=���S�j��
���銻����xJ��/̪��.���r����ɻ��ӻلݻ�M绩��y���[��L���=�����G�9���� p!���%��)��!.��C2��Y6��c:��b>��UB�k>F�GJ���M�'�Q��xU��.Y���\��`��d�خg�$:k���n��9r���u��y�׃|����ן��[J���&����9���ى�^w�����L����C��Fّ�m������������b����8���Ü�N��ן�6_���梼m����.x������O���F��������Ᏸ�J������$��ݝ���!������*�� ����5���  �  �cN=�M=�L=�L=�RK=o�J=�I=� I=�9H=�qG=,�F=��E=�E=hJD=a~C=k�B=m�A=dA=:D@=�r?=Z�>=��==i�<=� <=�H;=io:=a�9=��8=e�7=U�6=m6=�35=�M4=Df3=||2=��1=m�0=��/=1�.=��-=J�,=	�+=�*=��)=�(=��'=��&=��%=a�$=�#=��"=�t!=�Y =C;=f=�=!�=��=�n=�:=M=�=�=BF=��='�=�f=�=��=�d=�
=C�=�?=��=ti=��=&�=� =? �<_!�<��<��<��<���<��<���<(k�<�7�<��<��<�y�<�/�<\��<��<�2�<���<Hr�<��<<g2�<<��<�J�<�Ѯ<�U�<ק<�U�<Ҡ<(L�<Bę<�:�<M��<�"�<ٔ�<�<�v�<��<c�z<��s<�jl<�Je<L+^<{W<��O<��H<��A<��:<5�3<g�,<
�%<P�<��<��<=�	<q�<;��;Y��;�;�}�;���;Hq�;�;���;i�;;q|;7:b;z/H;Q.;�;B�:K��:�j�:(/?:ܶ�9i��Y�͹
G�C7��lvº�?�%����&�?k=���S�xj��
���銻����}J��̪�/���r����ɻN�ӻ؄ݻ�M绌�𻋅��<��H���=����H�3�����o!��%��)��!.��C2��Y6��c:�ub>�VB�[>F�FJ���M��Q��xU��.Y��\��`��d�ˮg�	:k���n��9r���u�my�Ӄ|����ן��cJ���%����9���ى�]w�����K����C��Jّ�m��/����������]����8���Ü��M��ן�-_��~梼m����7x������Q���B��������폰�I������+��ҝ���!������*������5���  �  �cN=�M=!�L=�L=�RK=p�J=x�I=� I=�9H=�qG='�F=��E=�E=iJD=i~C=l�B=q�A=\A=8D@=�r?=\�>=��==a�<=� <=�H;=ko:=c�9=��8=h�7=P�6=q6=�35=�M4=Ff3=r|2=��1=c�0=��/=1�.=�-=J�,=�+=�*=��)= �(=��'=��&=��%=_�$=�#=��"=�t!=�Y =D;=f=�='�=��=�n=�:=O=�=�=BF=��=)�=�f=�=��=�d=�
=@�=�?=��=i=��=�=� => �<t!�<��<��<��<���<��<���<0k�<�7�<��<ھ�<z�<�/�<b��<��<�2�<���<Hr�<��<�<k2�<7��<�J�<�Ѯ<�U�<%ק<�U�<Ҡ<,L�<Aę<�:�<C��<�"�<Ҕ�<�<�v�<��<��z<g�s<�jl<kJe<g+^<�W<��O<��H<��A<��:<�3<s�,<�%<S�<��<��<M�	<s�<a��;-��;��;�}�;���;�q�;#�;ϭ�;�h�;q|;n:b;�/H;7Q.;��;�B�:���:k�:�/?:���9(T����͹�
G�p7��>uº�?����y�&��k=�4�S�vj��
���銻����pJ��&̪��.���r��r�ɻy�ӻ�ݻ�M绊��u���c��E���=�����G�3����p!���%��)��!.��C2��Y6��c:��b>��UB�d>F�GJ���M�%�Q��xU��.Y���\��`��d��g�:k�z�n��9r�u�u��y�΃|����՟��[J���"����9���ى�Vw�����M����C��Eّ�m�� ����������b����8���Ü��M��ן�8_���梼	m����0x������J���I������}��台�7������3��坶��!������*�������5���  �  �cN=�M=&�L=�L=�RK=t�J=z�I=� I=�9H=�qG=(�F=��E=�E=eJD=i~C=e�B=t�A=]A==D@=�r?=T�>=��==b�<=� <=�H;=ho:=d�9=��8=m�7=L�6=s6=�35=�M4=<f3={|2=��1=_�0=��/=*�.= �-=J�,=	�+=!�*=�)=$�(=��'=��&=��%=b�$=�#=��"=�t!=�Y =G;=d=	�=%�=��=�n=�:=V=�=�=FF=��=,�=�f=�=��=�d=�
=>�=�?=�=~i=��=3�=� =+ �<k!�<y�<��<
��<���<��<���</k�<�7�<"��<��<z�<�/�<\��<���<�2�<���<>r�<��<�<n2�<8��<�J�<�Ѯ<�U�<&ק<�U�<Ҡ<$L�<5ę<�:�<:��<�"�<є�<�<�v�<��<l�z<g�s<kl<wJe<G+^<yW<��O<��H<��A<ͬ:<�3<��,<��%<<�<��<��<V�	<S�<���;7��;��;�}�;���;�q�;��;歘;�h�;mq|;e:b;#/H;iQ.;��;�C�:��:�j�:0?:��9],��׏͹p
G��7���uº�@�3���&�l=�K�S��j��
���銻����aJ��O̪��.���r��j�ɻ\�ӻфݻ�M����9���h��9���=����H�C����p!�޷%�(�)��!.��C2��Y6��c:��b>��UB�v>F�GJ���M�.�Q��xU�/Y���\�1�`�dd���g�1:k���n��9r�j�u��y���|����֟��\J��"�����9���ى�fw�����?����C��>ّ�m������������`����8���Ü�N��ן�5_��}梼m����(x������B���K�������������D������ ��ߝ���!������*�������5���  �  �cN=�M=!�L=�L=�RK=p�J=x�I=� I=�9H=�qG='�F=��E=�E=iJD=i~C=k�B=q�A=\A=8D@=�r?=\�>=��==a�<=� <=�H;=ko:=c�9=��8=h�7=P�6=q6=�35=�M4=Ff3=r|2=��1=c�0=��/=1�.=�-=J�,=�+=�*=��)= �(=��'=��&=��%=_�$=�#=��"=�t!=�Y =D;=f=�='�=��=�n=�:=O=�=�=BF=��=)�=�f=�=��=�d=�
=@�=�?=��=i=��=�=� => �<t!�<��<��<��<���<��<���<0k�<�7�<��<ھ�<z�<�/�<b��<��<�2�<���<Hr�<��<�<k2�<7��<�J�<�Ѯ<�U�<%ק<�U�<Ҡ<,L�<Aę<�:�<C��<�"�<Ҕ�<�<�v�<��<��z<g�s<�jl<kJe<g+^<�W<��O<��H<��A<��:<�3<s�,<�%<S�<��<��<M�	<s�<a��;-��;��;�}�;���;�q�;#�;ϭ�;�h�;q|;n:b;�/H;7Q.;��;�B�:���:k�:�/?:���9-T����͹�
G�q7��>uº�?����y�&��k=�4�S�vj��
���銻����pJ��&̪��.���r��r�ɻy�ӻ�ݻ�M绊��u���c��E���=�����G�3����p!���%��)��!.��C2��Y6��c:��b>��UB�d>F�GJ���M�%�Q��xU��.Y���\��`��d��g�:k�z�n��9r�u�u��y�΃|����՟��[J���"����9���ى�Vw�����M����C��Eّ�m�� ����������b����8���Ü��M��ן�8_���梼	m����0x������J���I������}��台�7������3��坶��!������*�������5���  �  �cN=�M=�L=�L=�RK=o�J=�I=� I=�9H=�qG=,�F=��E=�E=hJD=a~C=k�B=m�A=dA=:D@=�r?=Z�>=��==i�<=� <=�H;=io:=a�9=��8=e�7=U�6=m6=�35=�M4=Df3=||2=��1=m�0=��/=1�.=��-=J�,=	�+=�*=��)=�(=��'=��&=��%=a�$=�#=��"=�t!=�Y =C;=f=�=!�=��=�n=�:=M=�=�=BF=��='�=�f=�=��=�d=�
=C�=�?=��=ti=��=&�=� =? �<_!�<��<��<��<���<��<���<(k�<�7�<��<��<�y�<�/�<\��<��<�2�<���<Hr�<��<<g2�<<��<�J�<�Ѯ<�U�<ק<�U�<Ҡ<(L�<Bę<�:�<M��<�"�<ٔ�<�<�v�<��<c�z<��s<�jl<�Je<L+^<{W<��O<��H<��A<��:<5�3<g�,<
�%<P�<��<��<=�	<q�<;��;Y��;�;�}�;���;Hq�;�;���;i�;;q|;7:b;z/H;Q.;�;B�:K��:�j�:(/?:ܶ�9i��Z�͹
G�C7��lvº�?�%����&�?k=���S�xj��
���銻����}J��̪�/���r����ɻN�ӻ؄ݻ�M绌�𻋅��<��H���=����H�3�����o!��%��)��!.��C2��Y6��c:�ub>�VB�[>F�FJ���M��Q��xU��.Y��\��`��d�ˮg�	:k���n��9r���u�my�Ӄ|����ן��cJ���%����9���ى�]w�����K����C��Jّ�m��/����������]����8���Ü��M��ן�-_��~梼m����7x������Q���B��������폰�I������+��ҝ���!������*������5���  �  �cN=�M=#�L=�L=�RK=m�J=y�I=� I=�9H=�qG=(�F=��E=�E=jJD=i~C=j�B=p�A=aA=8D@=�r?=X�>=��==a�<=� <=�H;=jo:=c�9=��8=e�7=P�6=n6=�35=�M4==f3=x|2=��1=c�0=��/=6�.=��-=I�,=�+=�*=��)=!�(=��'=��&=��%=a�$=�#=��"=�t!=�Y =B;=f=�=(�=��=�n=�:=N=�=�=EF=��='�=�f=�=��=�d=�
=@�=�?=��=yi=��=&�=� =2 �<k!�<��<��<��<���<��<���<1k�<�7�<��<۾�<z�<�/�<Y��<��<�2�<���<Er�<��<���<j2�<6��<�J�<�Ѯ<�U�<*ק<�U�<Ҡ<"L�<Bę<�:�<A��<�"�<֔�<�<�v�<��<_�z<q�s<�jl<|Je<A+^<�W<��O<��H<��A<��:< �3<z�,<�%<D�<��<��<Y�	<d�<O��;6��;��;�}�;���;�q�;�;ĭ�;�h�;q|;1:b;b/H;rQ.;��;�B�:���:k�:�/?:o��9Eh����͹�G��6���uº�@�i����&��k=���S�j��
���銻����xJ��/̪��.���r����ɻ��ӻلݻ�M绩��y���[��L���=�����G�9���� p!���%��)��!.��C2��Y6��c:��b>��UB�k>F�GJ���M�'�Q��xU��.Y���\��`��d�خg�$:k���n��9r���u��y�׃|����ן��[J���&����9���ى�^w�����L����C��Fّ�m������������b����8���Ü�N��ן�6_���梼m����.x������O���F��������Ᏸ�J������$��ݝ���!������*�� ����5���  �  �cN=�M=!�L=�L=�RK=s�J=s�I=� I=�9H=�qG=(�F=��E=�E=dJD=k~C=g�B=r�A=_A=:D@=�r?=V�>=��==[�<=� <=�H;=io:=a�9=��8=k�7=P�6=q6=�35=�M4=Df3=x|2=��1=d�0=��/=/�.=��-=J�,=�+=%�*=�)= �(=��'=��&=��%=`�$=�#=��"=�t!=�Y =H;=b=�=&�=��=�n=�:=T=�=�=EF=��=/�=�f=�=��=�d=�
=A�=�?=��=}i=��=%�=� => �<o!�<~�<��<��<���<��<���<0k�<�7�<%��<Ͼ�<z�<�/�<`��<���<�2�<���<=r�<��<蠼<h2�<=��<�J�<�Ѯ<�U�<-ק<�U�<Ҡ<0L�<<ę<�:�<=��<�"�<Д�<�<�v�<��<{�z<r�s<�jl<|Je<]+^<�W<��O<��H<��A<ά:<�3<p�,<�%<S�<��<r�<_�	<Y�<��;7��;�;�}�;���;�q�;��;׭�;�h�;6q|;�:b;H/H;wQ.;2�;�C�:¤�:�j�:9/?:q��9d9��ٍ͹�
G��7���uº�?�j���&��k=�O�S��j��
���銻����BJ��N̪��.���r��D�ɻ��ӻ�ݻ�M绷��M���a��6���=�����G�I����p!��%��)��!.��C2��Y6��c:��b>��UB�z>F�1J���M�$�Q��xU�/Y���\��`��d�خg�:k���n��9r�w�u��y�ƃ|����ݟ��\J�������9���ى�^w�����G����C��@ّ�m������������[����8���Ü�
N��
ן�@_���梼m����2x������?���K���������鏰�<������$��ݝ���!������*�������5���  �  �cN=�M=!�L=�L=�RK=r�J=y�I=� I=�9H=�qG=%�F=��E=�E=iJD=i~C=l�B=m�A=_A=7D@=�r?=W�>=��==c�<=� <=�H;=io:=b�9=��8=g�7=Q�6=p6=�35=�M4=Bf3={|2=��1=h�0=��/=2�.=��-=J�,=�+="�*=��)= �(=��'=��&=��%=b�$=�#=��"=�t!=�Y =D;=d=�=(�=��=�n=�:=P=�=�=EF=��=*�=�f=�=��=�d=�
=A�=�?=��=wi=��=&�=� =: �<d!�<��<��<��<���<��<���<0k�<�7�<��<ݾ�<	z�<�/�<`��<��<�2�<���<Hr�<��<�<h2�<8��<�J�<�Ѯ<�U�<%ק<�U�<Ҡ<)L�<<ę<�:�<H��<�"�<Д�<�<�v�<��<d�z<��s<�jl<�Je<G+^<�W<��O<��H<��A<��:<+�3<o�,<�%<H�<��<��<P�	<h�<Y��;��;��;�}�;���;�q�;$�;���;�h�;q|;n:b;W/H;MQ.;��;HC�:���:�j�:g/?:@��99Z����͹G��6��vºG@�>���&��k=���S�fj��
���銻����UJ��,̪��.���r��i�ɻl�ӻτݻ�M绚��q���[��F���=�����G�8�����o!���%��)��!.��C2��Y6��c:��b>��UB�m>F�4J���M�!�Q��xU��.Y���\��`��d�Үg�:k���n��9r�y�u�}y�Ӄ|����ڟ��[J�������9���ى�`w�����M����C��Iّ�m������������`����8���Ü� N��ן�4_��~梼m����2x������I���K������~��돰�H������*��֝���!������*�������5���  �  �cN=�M=�L=�L=�RK=m�J=y�I=� I=�9H=�qG=)�F=��E=�E=kJD=^~C=n�B=l�A=fA=7D@=�r?=[�>=��==b�<=� <=�H;=jo:=_�9=��8=c�7=U�6=j6=�35=�M4=Bf3=y|2=��1=h�0=��/=8�.=��-=J�,=	�+=�*=��)=�(=��'=��&=��%=`�$=�#=��"=�t!=�Y =C;=e=�="�=��=�n=�:=J=�=�=CF=��='�=�f=�=��=�d=�
=B�=�?=��=vi=��=!�=� =< �<g!�<��<��<��<���<��<���<,k�<�7�<��<۾�<z�<�/�<]��<��<�2�<���<Jr�<��<�<f2�<:��<�J�<�Ѯ<�U�<ק<�U�<Ҡ<+L�<Eę<�:�<G��<�"�<ܔ�<�<�v�<��<g�z<��s<�jl<�Je<K+^<�W<��O<��H<��A<��:<(�3<f�,<�%<V�<��<��<>�	<t�<C��;<��;�;�}�;���;5q�;6�;���;i�;q|;H:b;�/H;Q.;��;�B�:D��:�j�:�.?:��9�{��=�͹�G��6���uº8@�`��j�&��k=���S�j��
���銻����{J��.̪�/��ur��x�ɻ��ӻ�ݻ�M绊�𻝅��?��L���=����H�5�����o!��%��)��!.��C2��Y6��c:�nb>��UB�q>F�FJ���M��Q��xU��.Y���\��`��d�ݮg�:k���n��9r���u�oy�݃|����ޟ��_J���&����9���ى�[w�����R����C��Nّ�
m��2����������^����8���Ü��M��ן�6_���梼
m����8x������T���?��������ߏ��F������7��՝���!������*������5���  �  �cN=�M=#�L=�L=�RK=p�J=z�I=� I=�9H=�qG=(�F=��E=�E=kJD=e~C=n�B=l�A=`A=9D@=�r?=V�>=��==c�<=� <=�H;=jo:=d�9=��8=g�7=T�6=o6=�35=�M4=Bf3=z|2=��1=g�0=��/=1�.=��-=K�,=�+=!�*=��)=!�(=��'=��&=��%=c�$=�#=��"=�t!=�Y =B;=d=
�=&�=��=�n=�:=P=�=�=GF=��=+�=�f=�=��=�d=�
=B�=�?=��=zi=��=(�=� =; �<i!�<��<��<��<���<��<���</k�<�7�<��<ܾ�<z�<�/�<^��<��<�2�<���<Kr�<��<���<f2�<5��<�J�<�Ѯ<�U�<%ק<�U�<Ҡ<(L�<;ę<�:�<G��<�"�<Ԕ�<�<�v�<��<j�z<|�s<�jl<�Je<Q+^<�W<��O<��H<��A<��:<'�3<z�,<�%<J�<��<��<S�	<[�<f��;9��;��;�}�;���;kq�;7�;���;�h�; q|;]:b;</H;]Q.;��; C�:���:�j�:�/?:���9{Y��-�͹pG�|7���uº(@�S��߸&��k=���S�uj��
���銻����bJ��#̪��.���r��f�ɻx�ӻɄݻ�M绣��k���N��P���=�����G�6�����o!���%��)��!.��C2��Y6��c:��b>��UB�g>F�:J���M��Q��xU��.Y���\��`��d�Ԯg�:k���n��9r�~�u�wy�҃|����֟��\J�������9���ى�bw�����L����C��Lّ�	m��%����������c����8���Ü�N��ן�2_���梼m����-x������K���G���������쏰�E������"��ٝ���!������*�������5���  �  �cN=�M=%�L=�L=�RK=p�J=u�I=� I=�9H=�qG=#�F=��E=�E=hJD=g~C=i�B=r�A=`A=7D@=�r?=V�>=��==^�<=� <=�H;=mo:=b�9=��8=j�7=O�6=t6=�35=�M4=Bf3=u|2=��1=b�0=��/=.�.=�-=K�,=�+="�*=~�)=%�(=��'=��&=��%=b�$=�#=��"=�t!=�Y =G;=f=
�=&�=��=�n=�:=Q=�=�=GF=��=+�=�f=�=��=�d=�
=A�=�?=��=}i=��='�=� =7 �<p!�<��<��<��<���<��<���<8k�<�7�<��<Ӿ�<z�<�/�<_��<��<�2�<���<Ar�<��<<m2�<<��<�J�<�Ѯ<�U�<.ק<�U�<Ҡ<(L�<>ę<�:�<8��<�"�<є�<�<�v�<��<|�z<h�s<�jl<mJe<\+^<�W<��O<��H<��A<Ƭ:<�3<��,<�%<G�<��<{�<d�	<[�<o��;��;�;�}�;���;|q�;�;ӭ�;�h�;q|;h:b;;/H;�Q.;X�;�B�:���:ek�:x/?:
��9=����͹
G�C7���uºC@���ڸ&��k=�N�S��j��
���銻����WJ��X̪��.���r��g�ɻ��ӻфݻ�M绯��h���h��9���=�����G�:����
p!���%��)��!.��C2��Y6��c:��b>��UB�{>F�9J���M�#�Q��xU�/Y���\�#�`��d��g�:k���n��9r�k�u��y�ƃ|����ܟ��SJ�������9���ى�aw�����L����C��@ّ�m��%����������\����8���Ü�N��	ן�;_���梼m����'x�����E���J������}��쏰�<��������䝶��!������*�������5���  �  �cN=�M=�L=�L=�RK=r�J=x�I=� I=�9H=�qG=)�F=��E=~E=gJD=h~C=i�B=k�A=eA=8D@=�r?=Y�>=��==`�<=� <=�H;=eo:=_�9=��8=i�7=Q�6=n6=�35=�M4=Df3=z|2=��1=f�0=��/=1�.=��-=H�,=�+=!�*=��)=�(=��'=��&=��%=_�$=�#=��"=�t!=�Y =E;=`=	�=&�=��=�n=�:=N=�=�=BF=��=+�=�f=�=��=�d=�
=@�=�?=��=yi=��=(�=� => �<f!�<��<��<��<���<��<���<&k�<�7�<��<ھ�<z�<�/�<\��<��<�2�<���<Ar�<��<<^2�<<��<�J�<�Ѯ<�U�< ק<�U�<Ҡ<+L�<<ę<�:�<E��<�"�<Ք�<�<�v�<��<t�z<w�s<�jl<�Je<Y+^<�W<��O<��H<��A<��:<(�3<g�,<�%<Q�<��<��<E�	<`�<V��;@��;�;}�;���;~q�;�;���;
i�;q|;V:b;i/H;(Q.;z�;0C�:��:cj�:�.?:#��9�L����͹�G�.7���uº@�H��׸&��k=���S�xj��
���銻����^J��(̪��.���r��e�ɻl�ӻ�ݻ�M绪�𻀅��E��C���=�����G�F�����o!���%� �)��!.��C2��Y6��c:��b>��UB�k>F�<J���M�(�Q��xU��.Y���\��`��d�Ѯg�:k���n��9r���u�y�Ѓ|����ݟ��eJ�������9���ى�\w�����L����C��Mّ�m��#����������\����8���Ü�N��ן�9_��梼
m����8x������F���F��������鏰�@������"��ٝ���!������*������5���  �  �cN=�M=�L=�L=�RK=n�J=}�I=� I=�9H=�qG=&�F=��E=�E=lJD=e~C=q�B=k�A=_A=7D@=�r?=Z�>=��==f�<=� <=�H;=ho:=e�9=��8=d�7=U�6=j6=�35=�M4=Bf3=w|2=��1=g�0=��/=6�.=��-=J�,=�+=�*=��)=�(=��'=��&=��%=a�$=�#=��"=�t!=�Y =?;=g=�='�=��=�n=�:=M=�=�=CF=��=%�=�f=�=��=�d=�
=B�=�?=��=xi=��=!�=� == �<i!�<��<��<��<���<��<���<*k�<�7�<��<��<z�<�/�<\��<��<�2�<���<Sr�<��<���<j2�<0��<�J�<�Ѯ<�U�<ק<�U�<Ҡ<)L�<Dę<�:�<S��<�"�<ٔ�<�<�v�<��<g�z<x�s<�jl<�Je<N+^<�W<��O<��H<��A<��:<>�3<j�,<�%<N�<��<��<B�	<n�<N��;&��;��;�}�;���;iq�;Q�;���;�h�;�p|;C:b;�/H;Q.;ڡ;�B�:	��:�j�:50?:��96u��f�͹�G�s6���uº*@�w��U�&��k=���S�j��
���銻�����J���˪��.��{r����ɻd�ӻބݻ�M绅�𻇅��V��Y���=�����G�)�����o!��%��)��!.��C2��Y6��c:�tb>��UB�P>F�IJ���M��Q��xU��.Y���\��`��d��g�:k���n��9r���u�qy���|����П��aJ���(����9���ى�[w�����Q����C��Rّ� m��$����������h����8���Ü��M��ן�2_���梼m����9x������S���B�����z��㏰�F������2��ڝ���!������*������5���  �  �cN=�M=!�L=�L=�RK=p�J=v�I=� I=�9H=�qG=&�F=��E=�E=cJD=`~C=g�B=t�A=bA=;D@=�r?=V�>=��==a�<=� <=�H;=ko:=b�9=��8=g�7=V�6=o6=�35=�M4=Df3=z|2=��1=g�0=��/=-�.=��-=L�,=�+=�*=��)=�(=��'=��&=��%=_�$=�#=��"=�t!=�Y =J;=e=�=�=��=�n=�:=R=�=�=BF=��=*�=�f=�=��=�d=�
=D�=�?=��=zi=��='�=� =? �<i!�<��<��<��<���<��<���</k�<�7�<��<ܾ�<z�<�/�<]��<���<�2�<���<?r�<��<㠼<p2�<A��<�J�<�Ѯ<�U�<&ק<�U�<Ҡ<,L�<Bę<�:�<C��<�"�<ݔ�<�<�v�<��<z�z<{�s<�jl<�Je<\+^<|W<��O<��H<��A<��:<#�3<o�,<�%<R�<��<~�<R�	<_�<n��;)��;�;�}�;���;Aq�;��;筘;�h�;?q|;Z:b;G/H;IQ.;��;
C�:��:k�:Z/?:_��9QY��I�͹eG�l7���uº�?�M���&��k=�z�S��j��
���銻q���}J��/̪��.���r��f�ɻ`�ӻ�ݻ�M绱��\���]��.���=���H�@����p!��%��)��!.��C2��Y6��c:��b>��UB�k>F�HJ���M��Q��xU�/Y���\��`��d�Ѯg�
:k���n��9r��u�py�σ|����ڟ��]J�������9���ى�`w�����G����C��=ّ�m��2����������W����8���Ü�N��ן�<_���梼	m����3x������M���>�������������=������!��ٝ���!������*�������5���  �  �dN==�M=u�L=4L=�TK=C�J=w�I=I=	<H=YtG=�F=��E=�E=�MD=�C=�B=[�A=~A=�H@=xw?=)�>=��==��<=_&<=�N;=ku:=��9=B�8=,�7=] 7=�6=B;5=�U4=mn3=�2=K�1=i�0=T�/=��.=��-=z�,=��+=��*=��)=��(=��'=��&=��%=�$=�#=��"=�!=<g =	I=\'=C=��=>�=W}=�I=i=D�=j�=�U==��=dv=7$=%�=1t=[
=��=!O=��=�x=�=�=� =�<�<�=�<X7�<
*�<��<���<���<���<y��<;O�<	�<��<���<�D�<G��<��<�D�<.��<��<��<���<�@�<�͵<W�<cݮ<�`�<�<�^�<5ڠ<mS�<�ʙ<@�<鳒<b&�<���<�<�w�<��<k�z<��s<7fl<#De<a#^<�W<�O<��H<ȱA<�:<ʉ3<r{,<Aq%<�k<�k<�p<�{	<&�<�J�;M��;���;�3�;��;�!�;ղ�;sW�;f�;ظ{;�{a;6kG;Ї-;��;͙�:Q��:9��: �;:!v�9�O�jչ^�J�'��Xkĺ�;�%����'�+q>��T��"k�����&o��</��Р��Q��7��������ʻi!Ի�޻����y����9�����{������j���T��!���%�**�=W.�Hx2�8�6�'�:���>�ۅB�$mF��IJ�N�;�Q���U��WY�-]�C�`�~@d���g��\k���n��Yr���u��:y���|�N ��2���4W��c���뢆��D��n䉼������������L���ᑼ6u�����񖖼�%��㲙��>���ɜ�cS���۟��c���ꢼ�p��~���d{������߃�����銭���*���#��N���g��ڝ��h!��m����)������$4���  �  �dN==�M=o�L=7L=~TK=E�J=y�I=I=	<H=RtG=�F=��E=�E=�MD=�C="�B=`�A=�A=�H@=rw?=&�>=��==��<=_&<=�N;=mu:=��9=B�8=4�7=e 7=�6=J;5=�U4=ln3=�2=I�1=l�0=L�/=��.=��-=��,=��+=��*=��)=��(=��'=��&=��%=߾$=ӭ#=��"=�!=>g =I=e'===��=F�=\}=�I=a=A�=_�=�U==��=fv=5$=&�=5t=f
=��="O=��=�x=�=�=� =�<�<�=�<e7�<
*�<��<��<���<���<}��<=O�<�<��<s��<~D�<=��<
��<�D�<8��<���<u�<�<�@�<�͵<
W�<Rݮ<�`�<��<�^�<<ڠ<iS�<�ʙ<@�<곒<j&�<Ɨ�<�<�w�<��<R�z<��s<$fl<-De<K#^<�W<,�O<��H<�A<�:<̉3<^{,<Mq%<�k<�k<�p<�{	<&�<�J�;��;���;/4�;��;N!�;���;�W�;��;g�{;{{a;kG;�-;C�;���:=��:{��:1�;:"v�9@2�aչ�J�
&���kĺ-<����'��p>���T��"k������n���.���Ϡ��Q��W�������ʻE!Ի޻���y�S���9����s{�����G���T��!��%�**�hW.�ex2�%�6�4�:���>��B�"mF��IJ��N��Q���U�zWY�K]�9�`��@d���g��\k���n��Yr���u�c:y���|�J ��4���1W��b�����D���䉼������������L���ᑼ+u����������%��ײ���>���ɜ�cS��ܟ��c���ꢼ�p��w���n{������փ��w��㊭���,���/��G���q��՝��r!��o����)������4���  �  �dN=?�M=p�L=9L=xTK=C�J=|�I=I=<H=TtG=�F=��E=�E=�MD=�C=&�B=X�A=�A=�H@=yw?=0�>=��==��<=[&<=�N;=nu:=��9=A�8=-�7=` 7=�6=L;5=�U4=on3=�2=H�1=s�0=H�/=��.=��-=}�,=��+=��*=��)=��(=��'=��&=��%=�$=ح#=��"=�!=@g =I=e'=A=��=G�=R}=�I=b=K�=f�=�U==��=gv=6$=)�=1t=]
=��=O=��=�x=�=�=� ==�<�=�<i7�<*�<��<���<���<���<~��<9O�<��<��<u��<�D�<M��<
��<�D�<$��<���<~�<���<�@�<�͵<W�<Uݮ<�`�<�<�^�<9ڠ<^S�<�ʙ<@�<ﳒ<_&�<���<�<�w�<��<K�z<��s<fl<EDe<K#^<�W<'�O<��H<ԱA<�:<Ӊ3<a{,<Vq%<�k<�k<�p<�{	<W�<�J�;*��;���; 4�;&��;w!�;��;XW�;��;g�{;�{a;�kG;2�-;�;?��:���:���:��;:�u�9�O��չ��J��%��Tlĺ�;����,�'��p>���T��"k�����o��)/��'Р��Q��R�������*ʻ<!Ի�޻���xy�P���9����v{��� ��C���T��!� �%��)*�LW.�\x2��6�H�:���>�߅B�mF��IJ� N�-�Q���U�tWY�X]�!�`��@d���g��\k��n��Yr���u�v:y���|�O ��1���0W��e��������D���䉼������������L���ᑼ'u�������%��ⲙ��>���ɜ�IS��ܟ��c���ꢼq��q���l{������ც����銭���,���3��;���s��ɝ��s!��r����)������4���  �  �dN=>�M=q�L=4L=TK=E�J=u�I=I=<H=RtG=�F=��E=�E=�MD=�C=!�B=^�A=�A=�H@=tw?=#�>=��==��<=a&<=�N;=ku:=��9=C�8=2�7=e 7=�6=C;5=�U4=nn3=�2=K�1=m�0=O�/=��.=��-=��,=��+=��*=��)=��(=��'=��&=��%=�$=խ#=��"=�!=Bg =I=c'=?=��=D�=X}=�I=a=@�=`�=�U==��=ev=6$=%�=7t=c
=��="O=��=�x=�=�=� = =�<�=�<Z7�<*�<��< ��<���<���<z��<>O�<�<
��<{��<zD�<@��<��<�D�<2��<��<{�<�<�@�<�͵<W�<Qݮ<�`�<
�<�^�<:ڠ<jS�<�ʙ<@�<곒<k&�<×�<(�<�w�<��<X�z<��s<7fl<-De<R#^<�W<	�O<��H<�A<�:<Љ3<f{,<Cq%<�k<�k<�p<�{	<�<�J�;F��;���;4�;��;f!�;鲥;�W�;��;��{;�{a;�jG;{�-;��;���:g��:G��:��;:�v�9�:�lչ��J��&��lĺ�;�	����'��p>�V�T��"k������n���.���Ϡ��Q��S��������ʻR!Ի޻����y�P���9����|{�����P���T��!��%�"**�fW.�^x2�/�6�'�:���>��B�%mF��IJ��N��Q���U��WY�>]�4�`��@d���g��\k���n��Yr���u�^:y���|�G ��5���3W��a���袆��D��z䉼������������L���ᑼ0u����������%��۲���>���ɜ�hS��ܟ��c���ꢼ�p��|���k{������Ճ��z��ڊ����)���,��H���g��՝��o!��l����)������4���  �  �dN=;�M=u�L=4L=TK=G�J=s�I=I=<H=[tG=ޫF=��E=�E=�MD=�C= �B=c�A=�A=�H@=}w?=$�>=��==��<=b&<=�N;=nu:=��9=@�8=0�7=\ 7=�6=E;5=�U4=kn3=�2=K�1=g�0=R�/=��.=��-=~�,=��+=��*=��)=��(=��'=��&=��%=�$=׭#=��"=�!=9g =I=c'===��=C�=[}=�I=g=I�=c�=�U==��=av=;$=#�=4t=[
=��=!O=��=�x=�=�=� =�<�<�=�<[7�<*�<��<���<���<���<���<2O�<�<��<���<|D�<S��<��<�D�<;��<��<��<�<�@�<�͵<W�<cݮ<�`�<�<�^�<=ڠ<mS�<�ʙ<@�<峒<k&�<���<"�<�w�<��<[�z<��s</fl<De<N#^<�W<�O<��H<��A<�:<ŉ3<t{,<Aq%<�k<�k<�p<�{	<#�<�J�;��;���;74�;���;|!�;㲥;�W�;s�;k�{;/|a;�jG;��-;��;.��:���:���:�;:{u�9�@�չ~�J��&��kĺ4<�*����'�Cq>�/�T��"k�����o��E/��Р��Q����������ʻT!Ի�޻��绥y����9����}{�����T���T�(�!���%��)*�[W.�Ox2�4�6�#�:���>�˅B�,mF��IJ�N�6�Q���U��WY�0]�I�`��@d���g��\k���n��Yr���u��:y���|�M ��3���,W��l���梆��D��r䉼������������L���ᑼ0u����������%��ݲ���>���ɜ�bS��ܟ��c���ꢼ�p��~���a{������Ճ�����������#���+��T���k��ߝ��q!��e����)������*4���  �  �dN=>�M=p�L=6L=|TK=E�J=}�I=I=<H=VtG=�F=��E=�E=�MD=�C="�B=W�A=�A=�H@=zw?='�>=��==��<=a&<=�N;=lu:=��9=C�8=0�7=c 7=�6=H;5=�U4=mn3=��2=G�1=s�0=I�/=��.=��-=��,=��+=��*=��)=��(=��'=��&=��%=�$=ѭ#=��"=�!=?g =	I=a'=A=��=C�=V}=�I=`=H�=^�=�U==��=bv=6$='�=4t=_
=��="O=��=�x=�=�=� ==�<�=�<^7�<*�<��<���<���<���<{��<3O�<�<��<v��<}D�<M��<��<�D�<&��<��<��<���<�@�<�͵<
W�<Xݮ<�`�<��<�^�<;ڠ<hS�<�ʙ<@�<볒<k&�<���<#�<�w�<��<M�z<��s<fl<MDe<J#^<�W< �O<��H<ڱA<�:<щ3<`{,<Kq%<�k<�k<�p<�{	<5�<�J�;��;���;�3�;��;�!�;�;SW�;��;L�{;�{a;kG;#�-;g�;��:���:a��:B�;:�v�9/@��չ��J�^&��7lĺ�;����9�'��p>���T��"k������n�� /��Р��Q��P��������ʻA!Ի�޻�统y�N���9�����{������R���T�	�!��%�**�mW.�Yx2�#�6�-�:���>���B�mF��IJ��N��Q���U��WY�X]�"�`��@d���g��\k��n��Yr���u�g:y���|�J ��4���2W��k���袆��D���䉼������������L���ᑼ.u�����򖖼�%��ڲ���>���ɜ�XS��ܟ��c���ꢼ�p��y���n{������Ճ�����ߊ����.���1��8���y��ŝ��s!��t����)������4���  �  �dN=C�M=m�L=7L=�TK=?�J=~�I=I=<H=PtG=�F=��E=�E=�MD=��C=*�B=X�A=�A=�H@=uw?=+�>=��==��<=Y&<=�N;=mu:=��9=F�8=,�7=e 7=�6=L;5=�U4=nn3=�2=A�1=v�0=H�/=��.=��-=��,=��+=��*=��)=~�(=��'=��&=��%=�$=ԭ#=��"=�!=Eg =I=h'=>=��=K�=T}=�I=\=I�=a�=�U==��=gv=4$=*�=3t=a
=��=O=��=�x=�=�=� ==�<�=�<j7�<�)�<��<���<���<���<z��<@O�<��<��<w��<�D�<I��<��<�D�<&��<��<l�<���<�@�<�͵<W�<Jݮ<�`�<��<�^�<1ڠ<lS�<�ʙ<@�<�<`&�<ȗ�<�<�w�<��<B�z<��s<�el<LDe<@#^<�W<�O<��H<�A<�:<�3<T{,<Pq%<�k<sk<�p<�{	<G�<�J�;>��;���;4�;7��;)!�;1��;ZW�;��;K�{;�{a;ZkG;,�-;u�;��:���:i��:�;:Tx�9�P�չ@�J��%���kĺ�;������'�Vp>���T�t"k�ҏ���n��/��Р��Q��f�������ʻM!Ի�޻�绐y�z��}9����i{�����3���T��!��%��)*�`W.�Ux2�"�6�:�:���>��B�mF��IJ��N��Q���U�fWY�U]��`��@d���g��\k���n��Yr���u�c:y���|�F ��4���4W��^��������D��~䉼�������µ���L���ᑼu�������%��ڲ���>���ɜ�QS��ܟ��c���ꢼ�p��t���t{����������v��ꊭ������7��7������Ɲ��x!��e����)������4���  �  �dN=B�M=s�L=2L=TK=B�J=z�I=I=<H=UtG=�F=��E=�E=�MD=�C=)�B=[�A=�A=�H@=zw?=&�>=��==��<=\&<=�N;=ku:=��9=D�8=,�7=b 7=�6=E;5=�U4=jn3=�2=L�1=m�0=I�/=��.=��-=��,=��+=��*=��)=��(=��'=��&=��%=�$=ԭ#=��"=�!=?g =I=f'=@=��=I�=S}=�I=c=I�=a�=�U==��=bv=8$=)�=2t=\
=��=O=��=�x=�=�=� =�<�<�=�<]7�<
*�<��<���<���<���<z��<7O�<�<��<��<~D�<O��<��<�D�<)��< ��<y�<���<�@�<�͵<W�<Uݮ<�`�<�<�^�<5ڠ<lS�<�ʙ<@�<�<`&�<���<"�<�w�<��<?�z<��s<0fl<4De<<#^<�W<�O<��H<ٱA<�:<މ3<l{,<;q%<�k<k<�p<�{	<7�<�J�;6��;���;4�;;��;Z!�;'��;rW�;��;z�{; |a;kG;��-;;�;m��:2��:9��:�;:Nw�9tQ��չ��J��&���kĺn<�����'��p>���T��"k������n��-/��Р��Q��3��������ʻU!Ի�޻��绕y�>���9����p{�����>���T��!���%��)*�bW.�Rx2�-�6�2�:���>�ׅB�mF��IJ�N��Q���U�}WY�P]�7�`�|@d���g��\k���n��Yr���u�l:y���|�J ��/���3W��g���𢆼�D��w䉼������������L���ᑼ!u�����떖��%��岙��>���ɜ�XS��ܟ��c���ꢼ�p������e{������ც����������#���9��F���j��ҝ��z!��f����)������4���  �  �dN=8�M=v�L=5L=}TK=G�J=w�I=I=<H=VtG=�F=��E=�E=�MD=�C=�B=_�A=�A=�H@=yw?= �>=��==��<=c&<=�N;=nu:=��9=>�8=5�7=^ 7=�6=A;5=�U4=on3=�2=J�1=l�0=S�/=��.=��-=��,=��+=��*=��)=��(=��'=��&=��%=�$=ӭ#=��"=�!=>g =I=a'=?=��=@�=]}=�I=b=B�=^�=�U==��=`v=:$=$�=6t=`
=��=%O=��=�x=�=�=� = =�<�=�<Q7�<*�<��< ��<���<���<��<4O�<�<��<~��<tD�<G��<��<�D�<7��<��<��<쯼<�@�<�͵<
W�<Yݮ<�`�<�<�^�<<ڠ<lS�<�ʙ<@�<೒<s&�<���<+�<�w�<��<k�z<��s<%fl<(De<a#^<�W<�O<��H<ȱA</�:<��3<w{,<Eq%<�k<�k<�p<�{	<�<�J�;��;���;4�;ܡ�;�!�;���;�W�;��;P�{;�{a;�jG;}�-;�;K��:���:���:�;:Yt�9�/��չ4�J�E'���kĺ�;�$���'��p>��T�Q#k������n��#/���Ϡ��Q��(��������ʻX!Ի�޻	���y�@���9�����{������_���T��!���%�**�nW.�Sx2�7�6��:���>�υB�)mF��IJ��N��Q�z�U��WY�5]�9�`��@d���g��\k���n��Yr�x�u�s:y���|�N ��2���.W��k���⢆��D��w䉼Ł����������L���ᑼ;u����������%��Ӳ���>���ɜ�fS��ܟ��c���ꢼ�p�����b{������΃�����׊����1���#��J���p��؝��g!��r����)������%4���  �  �dN=9�M=t�L=6L=}TK=C�J=y�I=I=<H=XtG=ޫF=��E=�E=�MD=�C=!�B=^�A=�A=�H@=}w?=*�>=��==��<=^&<=�N;=lu:=��9=?�8=4�7=Z 7=�6=J;5=�U4=mn3=�2=G�1=m�0=N�/=��.=��-=z�,=��+=��*=��)=��(=��'=��&=��%=�$=ح#=��"=�!=>g =	I=d'=?=��=E�=X}=�I=c=K�=d�=�U==��=ev=9$=&�=2t=]
=��= O=��=�x=�=�=� =�<�<�=�<c7�<*�<��<���<~��<���<|��<8O�<�<��<���<�D�<R��<��<�D�<3��<��<��<�<�@�<�͵<W�<^ݮ<�`�<�<�^�<8ڠ<iS�<�ʙ<@�<䳒<n&�<���<�<�w�<��<X�z<��s<fl<.De<O#^<�W<&�O<��H<��A<(�:<��3<n{,<Hq%<�k<�k<�p<�{	<@�<�J�;	��;���; 4�; ��;�!�;첥;�W�;��;?�{;)|a;EkG;��-;3�;���:��:b��:�;:�t�9"3��չ;�J�&���kĺ<���/�'��p>�h�T��"k�����%o��0/��Р��Q��0��������ʻW!Ի�޻��练y�9���9����y{��� ��L���T��!���%��)*�TW.�Jx2�2�6�2�:���>�ӅB�"mF��IJ��N�=�Q���U�~WY�B]�6�`��@d���g��\k���n��Yr���u��:y���|�Q ��2���1W��f�����D��t䉼������������L���ᑼ.u����������%��ಙ��>���ɜ�TS��ܟ��c���ꢼ�p��x���e{������Ӄ�����銭���*���-��H���t��՝��q!��m����)������(4���  �  �dN=A�M=p�L=0L=�TK=B�J=y�I=I=<H=PtG=�F=��E=�E=�MD=�C=(�B=Z�A=�A=�H@=uw?=%�>=��==��<=]&<=�N;=eu:=��9=C�8=2�7=i 7=�6=H;5=�U4=ln3=�2=I�1=q�0=G�/=��.=��-=��,=��+=��*=��)=|�(=��'=��&=��%=�$=ҭ#=��"=�!=Dg =I=g'=@=��=I�=R}=�I=_=D�=^�=�U==��=fv=1$=*�=1t=e
=��=!O=��=�x=�=�=� = =�<�=�<`7�<	*�<��<���<���<���<o��<CO�<�<��<t��<}D�<D��<
��<�D�<'��<���<{�<���<�@�<͵<W�<Mݮ<�`�<��<�^�<7ڠ<oS�<�ʙ<	@�<�<b&�<З�<�<�w�<��<A�z<��s<%fl<BDe<A#^<�W<�O<��H<��A<�:<ۉ3<`{,<1q%<�k<�k<�p<�{	<1�<�J�;H��;���;4�;*��;j!�;!��;iW�;��;��{;�{a;�jG;�-;W�;���:���:���:ޡ;:�v�9�:�չ�J�f&��*lĺ0<�����'��p>���T��"k������n���.��!Р��Q��v��������ʻE!Ի�޻�绸y�k���9����k{�����;���T���!��%�**�lW.�_x2�$�6�/�:���>���B�mF��IJ��N��Q���U�{WY�]]�'�`��@d���g��\k��n��Yr���u�U:y���|�M ��/���>W��\���𢆼�D���䉼������������L���ᑼ"u�������%��岙��>���ɜ�\S��ܟ��c���ꢼ�p������p{������ރ��m��㊭���)���7��>���p��˝��x!��o����)������4���  �  �dN=>�M=s�L=5L=�TK=A�J=x�I=I=<H=TtG=�F=��E=�E=�MD=�C=!�B=\�A=�A=�H@=xw?=,�>=��==��<=]&<=�N;=ku:=��9=@�8=,�7=] 7=�6=E;5=�U4=on3=�2=E�1=o�0=Q�/=��.=��-=z�,=��+=��*=��)=��(=��'=��&=��%=�$=ۭ#=��"=�!=Bg =	I=b'=@=��=C�=V}=�I=b=I�=g�=�U==��=fv=6$=(�=0t=]
=��=!O=��=�x=�=�=� ==�<�=�<[7�<*�<��<���<}��<���<y��<>O�<�<
��<~��<�D�<K��<��<�D�<.��<��<~�<�<�@�<�͵<W�<Tݮ<�`�<�<�^�<4ڠ<mS�<�ʙ<@�<쳒<^&�<���<�<�w�<��<b�z<��s<fl<1De<[#^<�W<�O<��H<ͱA<�:<Ή3<m{,<Dq%<�k<{k<�p<�{	<D�<�J�;L��;���;4�;��;u!�;;}W�;��;��{;�{a;`kG;r�-;,�;���:y��:O��:9�;:�u�9�O�Uչ2�J��&��Pkĺ�;���Z�'��p>�6�T��"k�����*o��$/��*Р��Q��L��������ʻU!Ի�޻��绑y�H���9����{������R���T��!���%��)*�HW.�Ox2�/�6�2�:���>��B�mF��IJ��N�<�Q���U��WY�6]�-�`��@d���g��\k���n��Yr���u��:y���|�R ��/���4W��`���񢆼�D��w䉼������������L���ᑼ/u����������%��޲���>���ɜ�RS��ܟ��c���ꢼ�p��{���h{������⃪�������'���'��E���{��ӝ��k!��j����)������"4���  �  �dN=<�M=q�L=6L=}TK=F�J=x�I=I=	<H=RtG=߫F=��E=�E=�MD=�C=�B=c�A=�A=�H@=tw?=#�>=��==��<=b&<=�N;=nu:=��9=B�8=:�7=] 7=�6=G;5=�U4=gn3=�2=N�1=h�0=M�/=��.=��-=~�,=��+=��*=��)=��(=��'=��&=��%=�$=ѭ#=��"=�!=<g =I=a'=?=��=A�=^}=�I=b=A�=\�=�U==��=dv=9$=$�=8t=g
=��=(O=��=�x=�=�=� =�<�<�=�<Z7�<*�<��<��<���<���<~��<8O�<�<��<w��<xD�<@��<��<�D�<=��<��<��<ﯼ<�@�<�͵<W�<Pݮ<�`�<��<�^�<<ڠ<hS�<�ʙ<@�<䳒<v&�<���<!�<�w�<��<L�z<��s<2fl<,De<A#^<�W<.�O<��H<ϱA<;�:<Ɖ3<f{,<Jq%<�k<�k<�p<�{	<%�<�J�;��;���;64�;��;�!�;ϲ�;�W�;��;\�{;�{a;�jG;6�-;)�;��:��:���:3�;:zv�9X�Sչ�J�m&��lĺ�<����ƻ'�-q>��T�H#k�{���	o���.���Ϡ��Q��9��������ʻT!Ի�޻���y�C���9�����{������[���T��!���%�**�sW.�ax2�1�6�.�:���>�ԅB�*mF��IJ��N�.�Q�p�U��WY�G]�N�`�r@d���g��\k���n��Yr�v�u�}:y���|�J ��8���/W��f���袆��D��~䉼������������L���ᑼ7u����������%��ٲ���>���ɜ�cS��ܟ��c���ꢼ�p��y���i{������ʃ��~��ክ���4���3��L���j��֝��w!��u����)������!4���  �  �dN=>�M=s�L=5L=�TK=A�J=x�I=I=<H=TtG=�F=��E=�E=�MD=�C=!�B=\�A=�A=�H@=xw?=,�>=��==��<=]&<=�N;=ku:=��9=@�8=,�7=] 7=�6=E;5=�U4=on3=�2=E�1=o�0=Q�/=��.=��-=z�,=��+=��*=��)=��(=��'=��&=��%=�$=ۭ#=��"=�!=Bg =	I=b'=@=��=C�=V}=�I=b=I�=g�=�U==��=fv=6$=(�=0t=]
=��=!O=��=�x=�=�=� ==�<�=�<[7�<*�<��<���<}��<���<y��<>O�<�<
��<~��<�D�<K��<��<�D�<.��<��<~�<�<�@�<�͵<W�<Tݮ<�`�<�<�^�<4ڠ<mS�<�ʙ<@�<쳒<^&�<���<�<�w�<��<b�z<��s<fl<1De<[#^<�W<�O<��H<ͱA<�:<Ή3<m{,<Dq%<�k<{k<�p<�{	<D�<�J�;L��;���;4�;��;u!�;;}W�;��;��{;�{a;`kG;r�-;,�;���:y��:O��:9�;:�u�9�O�Uչ3�J��&��Pkĺ�;���Z�'��p>�6�T��"k�����*o��$/��*Р��Q��L��������ʻU!Ի�޻��绑y�H���9����{������R���T��!���%��)*�HW.�Ox2�/�6�2�:���>��B�mF��IJ��N�<�Q���U��WY�6]�-�`��@d���g��\k���n��Yr���u��:y���|�R ��/���4W��`���񢆼�D��w䉼������������L���ᑼ/u����������%��޲���>���ɜ�RS��ܟ��c���ꢼ�p��{���h{������⃪�������'���'��E���{��ӝ��k!��j����)������"4���  �  �dN=A�M=p�L=0L=�TK=B�J=y�I=I=<H=PtG=�F=��E=�E=�MD=�C=(�B=Z�A=�A=�H@=uw?=%�>=��==��<=]&<=�N;=eu:=��9=C�8=2�7=i 7=�6=H;5=�U4=ln3=�2=I�1=q�0=G�/=��.=��-=��,=��+=��*=��)=|�(=��'=��&=��%=�$=ҭ#=��"=�!=Dg =I=g'=@=��=I�=R}=�I=_=D�=^�=�U==��=fv=1$=*�=1t=e
=��=!O=��=�x=�=�=� = =�<�=�<`7�<	*�<��<���<���<���<o��<CO�<�<��<t��<}D�<D��<
��<�D�<'��<���<{�<���<�@�<͵<W�<Mݮ<�`�<��<�^�<7ڠ<oS�<�ʙ<	@�<�<b&�<З�<�<�w�<��<A�z<��s<%fl<BDe<A#^<�W<�O<��H<��A<�:<ۉ3<a{,<1q%<�k<�k<�p<�{	<1�<�J�;H��;���;4�;*��;j!�;!��;iW�;��;��{;�{a;�jG;�-;W�;���:���:���:ޡ;:�v�9;�չ�J�f&��*lĺ1<�����'��p>���T��"k������n���.��!Р��Q��v��������ʻE!Ի�޻�绸y�k���9����k{�����;���T���!��%�**�lW.�_x2�$�6�/�:���>���B�mF��IJ��N��Q���U�{WY�]]�'�`��@d���g��\k��n��Yr���u�U:y���|�M ��/���>W��\���𢆼�D���䉼������������L���ᑼ"u�������%��岙��>���ɜ�\S��ܟ��c���ꢼ�p������p{������ރ��m��㊭���)���7��>���p��˝��x!��o����)������4���  �  �dN=9�M=t�L=6L=}TK=C�J=y�I=I=<H=XtG=ޫF=��E=�E=�MD=�C=!�B=^�A=�A=�H@=}w?=*�>=��==��<=^&<=�N;=lu:=��9=?�8=4�7=Z 7=�6=J;5=�U4=mn3=�2=G�1=m�0=N�/=��.=��-=z�,=��+=��*=��)=��(=��'=��&=��%=�$=ح#=��"=�!=>g =	I=d'=?=��=E�=X}=�I=c=K�=d�=�U==��=ev=9$=&�=2t=]
=��= O=��=�x=�=�=� =�<�<�=�<c7�<*�<��<���<~��<���<|��<8O�<�<��<���<�D�<R��<��<�D�<3��<��<��<�<�@�<�͵<W�<^ݮ<�`�<�<�^�<8ڠ<iS�<�ʙ<@�<䳒<n&�<���<�<�w�<��<X�z<��s<fl<.De<O#^<�W<&�O<��H<��A<(�:<��3<n{,<Hq%<�k<�k<�p<�{	<@�<�J�;	��;���; 4�; ��;�!�;첥;�W�;��;?�{;)|a;EkG;��-;3�;���:��:b��:�;:�t�9,3��չ<�J�&���kĺ<���/�'��p>�h�T��"k�����%o��0/��Р��Q��0��������ʻW!Ի�޻��练y�9���9����y{��� ��L���T��!���%��)*�TW.�Jx2�2�6�2�:���>�ӅB�"mF��IJ��N�=�Q���U�~WY�B]�6�`��@d���g��\k���n��Yr���u��:y���|�Q ��2���1W��f�����D��t䉼������������L���ᑼ.u����������%��ಙ��>���ɜ�TS��ܟ��c���ꢼ�p��x���e{������Ӄ�����銭���*���-��H���t��՝��q!��m����)������(4���  �  �dN=8�M=v�L=5L=}TK=G�J=w�I=I=<H=VtG=�F=��E=�E=�MD=�C=�B=_�A=�A=�H@=yw?= �>=��==��<=c&<=�N;=nu:=��9=>�8=5�7=^ 7=�6=A;5=�U4=on3=�2=J�1=l�0=S�/=��.=��-=��,=��+=��*=��)=��(=��'=��&=��%=�$=ӭ#=��"=�!=>g =I=a'=?=��=@�=]}=�I=b=B�=^�=�U==��=`v=:$=$�=6t=`
=��=%O=��=�x=�=�=� = =�<�=�<Q7�<*�<��< ��<���<���<��<4O�<�<��<��<tD�<G��<��<�D�<7��<��<��<쯼<�@�<�͵<
W�<Yݮ<�`�<�<�^�<<ڠ<lS�<�ʙ<@�<೒<s&�<���<+�<�w�<��<k�z<��s<%fl<(De<a#^<�W<�O<��H<ȱA</�:<��3<w{,<Eq%<�k<�k<�p<�{	<�<�J�;��;���;4�;ܡ�;�!�;���;�W�;��;P�{;�{a;�jG;}�-;�;J��:���:���:�;:Wt�9�/��չ5�J�E'���kĺ�;�$���'��p>��T�Q#k������n��#/���Ϡ��Q��(��������ʻX!Ի�޻	���y�@���9�����{������_���T��!���%�**�nW.�Sx2�8�6��:���>�υB�*mF��IJ��N��Q�z�U��WY�5]�9�`��@d���g��\k���n��Yr�x�u�s:y���|�N ��2���.W��k���⢆��D��w䉼Ł����������L���ᑼ;u����������%��Ӳ���>���ɜ�fS��ܟ��c���ꢼ�p�����b{������΃�����׊����1���#��J���p��؝��g!��r����)������%4���  �  �dN=B�M=s�L=2L=TK=B�J=z�I=I=<H=UtG=�F=��E=�E=�MD=�C=)�B=[�A=�A=�H@=zw?=&�>=��==��<=\&<=�N;=ku:=��9=D�8=,�7=b 7=�6=E;5=�U4=jn3=�2=L�1=m�0=I�/=��.=��-=��,=��+=��*=��)=��(=��'=��&=��%=�$=ԭ#=��"=�!=?g =I=f'=@=��=I�=S}=�I=c=I�=a�=�U==��=bv=8$=)�=2t=\
=��=O=��=�x=�=�=� =�<�<�=�<]7�<
*�<��<���<���<���<z��<7O�<�<��<��<~D�<O��<��<�D�<)��< ��<y�<���<�@�<�͵<W�<Uݮ<�`�<�<�^�<5ڠ<lS�<�ʙ<@�<�<`&�<���<"�<�w�<��<?�z<��s<0fl<4De<<#^<�W<�O<��H<ٱA<�:<މ3<l{,<;q%<�k<k<�p<�{	<7�<�J�;6��;���;4�;;��;Z!�;'��;qW�;��;y�{; |a;kG;��-;:�;l��:1��:9��:�;:Mw�9Q��չ��J��&���kĺn<�����'��p>���T��"k������n��-/��Р��Q��3��������ʻU!Ի�޻��绕y�>���9����p{�����>���T��!���%��)*�bW.�Rx2�-�6�2�:���>�ׅB�mF��IJ�N��Q���U�}WY�P]�7�`�|@d���g��\k���n��Yr���u�l:y���|�J ��/���3W��g���𢆼�D��w䉼������������L���ᑼ!u�����떖��%��岙��>���ɜ�XS��ܟ��c���ꢼ�p������e{������ც����������#���9��F���j��ҝ��z!��f����)������4���  �  �dN=C�M=m�L=7L=�TK=?�J=~�I=I=<H=PtG=�F=��E=�E=�MD=��C=*�B=X�A=�A=�H@=uw?=+�>=��==��<=Y&<=�N;=mu:=��9=F�8=,�7=e 7=�6=L;5=�U4=nn3=�2=A�1=v�0=H�/=��.=��-=��,=��+=��*=��)=~�(=��'=��&=��%=�$=ԭ#=��"=�!=Eg =I=h'=>=��=K�=T}=�I=\=I�=a�=�U==��=gv=4$=*�=3t=a
=��=O=��=�x=�=�=� ==�<�=�<j7�<�)�<��<���<���<���<z��<@O�<��<��<w��<�D�<I��<��<�D�<&��<��<l�<���<�@�<�͵<W�<Jݮ<�`�<��<�^�<1ڠ<lS�<�ʙ<@�<�<`&�<ȗ�<�<�w�<��<B�z<��s<�el<LDe<@#^<�W<�O<��H<�A<�:<�3<T{,<Pq%<�k<sk<�p<�{	<G�<�J�;>��;���;4�;7��;)!�;1��;ZW�;��;K�{;�{a;YkG;,�-;u�;��:���:i��:�;:Sx�9�P�չ@�J��%���kĺ�;������'�Vp>���T�t"k�ҏ���n��/��Р��Q��f�������ʻM!Ի�޻�绐y�z��}9����i{�����3���T��!��%��)*�`W.�Ux2�"�6�:�:���>��B�mF��IJ��N��Q���U�fWY�U]��`��@d���g��\k���n��Yr���u�c:y���|�F ��4���4W��^��������D��~䉼�������µ���L���ᑼu�������%��ڲ���>���ɜ�QS��ܟ��c���ꢼ�p��t���t{����������v��ꊭ������7��7������Ɲ��x!��e����)������4���  �  �dN=>�M=p�L=6L=|TK=E�J=}�I=I=<H=VtG=�F=��E=�E=�MD=�C="�B=W�A=�A=�H@=zw?='�>=��==��<=a&<=�N;=lu:=��9=C�8=0�7=c 7=�6=H;5=�U4=mn3=��2=G�1=s�0=I�/=��.=��-=��,=��+=��*=��)=��(=��'=��&=��%=�$=ѭ#=��"=�!=?g =	I=a'=B=��=C�=V}=�I=`=H�=^�=�U==��=bv=6$='�=4t=_
=��="O=��=�x=�=�=� ==�<�=�<^7�<*�<��<���<���<���<{��<3O�<�<��<v��<}D�<M��<��<�D�<&��<��<��<���<�@�<�͵<
W�<Xݮ<�`�<��<�^�<;ڠ<hS�<�ʙ<@�<볒<k&�<���<#�<�w�<��<M�z<��s<fl<MDe<J#^<�W< �O<��H<ڱA<�:<щ3<`{,<Kq%<�k<�k<�p<�{	<5�<�J�;��;���;�3�;��;�!�;�;SW�;��;L�{;�{a;kG;#�-;g�;��:���:a��:B�;:�v�9:@��չ��J�_&��7lĺ�;����9�'��p>���T��"k������n�� /��Р��Q��P��������ʻA!Ի�޻�统y�N���9�����{������R���T�	�!��%�**�mW.�Yx2�#�6�-�:���>���B�mF��IJ��N��Q���U��WY�X]�"�`��@d���g��\k��n��Yr���u�g:y���|�J ��4���2W��k���袆��D���䉼������������L���ᑼ.u�����򖖼�%��ڲ���>���ɜ�XS��ܟ��c���ꢼ�p��y���n{������Ճ�����ߊ����.���1��8���y��ŝ��s!��t����)������4���  �  �dN=;�M=u�L=4L=TK=G�J=s�I=I=<H=[tG=ޫF=��E=�E=�MD=�C= �B=c�A=�A=�H@=}w?=$�>=��==��<=b&<=�N;=nu:=��9=@�8=0�7=\ 7=�6=E;5=�U4=kn3=�2=K�1=g�0=R�/=��.=��-=~�,=��+=��*=��)=��(=��'=��&=��%=�$=׭#=��"=�!=9g =I=c'===��=C�=[}=�I=g=I�=c�=�U==��=av=;$=#�=4t=[
=��=!O=��=�x=�=�=� =�<�<�=�<[7�<*�<��<���<���<���<���<2O�<�<��<���<|D�<S��<��<�D�<;��<��<��<�<�@�<�͵<W�<cݮ<�`�<�<�^�<=ڠ<mS�<�ʙ<@�<峒<k&�<���<"�<�w�<��<[�z<��s</fl<De<N#^<�W<�O<��H<��A<�:<ŉ3<t{,<Aq%<�k<�k<�p<�{	<#�<�J�;��;���;74�;���;|!�;㲥;�W�;s�;k�{;/|a;�jG;��-;��;-��:���:���:�;:zu�9A�չ�J��&��kĺ5<�*����'�Cq>�/�T��"k�����o��E/��Р��Q����������ʻT!Ի�޻��绥y����9����}{�����T���T�(�!���%��)*�[W.�Ox2�4�6�#�:���>�˅B�,mF��IJ�N�6�Q���U��WY�0]�I�`��@d���g��\k���n��Yr���u��:y���|�M ��3���,W��l���梆��D��r䉼������������L���ᑼ0u����������%��ݲ���>���ɜ�bS��ܟ��c���ꢼ�p��~���a{������Ճ�����������#���+��T���k��ߝ��q!��e����)������*4���  �  �dN=>�M=q�L=4L=TK=E�J=u�I=I=<H=RtG=�F=��E=�E=�MD=�C=!�B=^�A=�A=�H@=tw?=#�>=��==��<=a&<=�N;=ku:=��9=C�8=2�7=e 7=�6=C;5=�U4=nn3=�2=K�1=m�0=O�/=��.=��-=��,=��+=��*=��)=��(=��'=��&=��%=�$=խ#=��"=�!=Bg =I=c'=?=��=D�=X}=�I=a=@�=`�=�U==��=ev=6$=%�=7t=c
=��="O=��=�x=�=�=� = =�<�=�<Z7�<*�<��< ��<���<���<z��<>O�<�<
��<{��<zD�<@��<��<�D�<2��<��<{�<�<�@�<�͵<W�<Qݮ<�`�<
�<�^�<:ڠ<jS�<�ʙ<@�<곒<k&�<×�<(�<�w�<��<X�z<��s<7fl<-De<R#^<�W<	�O<��H<�A<�:<Љ3<f{,<Cq%<�k<�k<�p<�{	<�<�J�;F��;���;4�;��;f!�;鲥;�W�;��;��{;�{a;�jG;{�-;��;���:g��:G��:��;:�v�9�:�mչ��J��&��lĺ�;�	����'��p>�V�T��"k������n���.���Ϡ��Q��S��������ʻR!Ի޻����y�P���9����|{�����P���T��!��%�"**�fW.�^x2�/�6�'�:���>��B�%mF��IJ��N��Q���U��WY�>]�4�`��@d���g��\k���n��Yr���u�^:y���|�G ��5���3W��a���袆��D��z䉼������������L���ᑼ0u����������%��۲���>���ɜ�hS��ܟ��c���ꢼ�p��|���k{������Ճ��z��ڊ����)���,��H���g��՝��o!��l����)������4���  �  �dN=?�M=p�L=9L=xTK=C�J=|�I=I=<H=TtG=�F=��E=�E=�MD=�C=&�B=X�A=�A=�H@=yw?=0�>=��==��<=[&<=�N;=nu:=��9=A�8=-�7=` 7=�6=L;5=�U4=on3=�2=H�1=s�0=H�/=��.=��-=}�,=��+=��*=��)=��(=��'=��&=��%=�$=ح#=��"=�!=@g =I=e'=A=��=G�=R}=�I=b=K�=f�=�U==��=gv=6$=)�=1t=]
=��=O=��=�x=�=�=� ==�<�=�<i7�<*�<��<���<���<���<~��<9O�<��<��<u��<�D�<M��<
��<�D�<$��<���<~�<���<�@�<�͵<W�<Uݮ<�`�<�<�^�<9ڠ<^S�<�ʙ<@�<ﳒ<_&�<���<�<�w�<��<K�z<��s<fl<EDe<K#^<�W<'�O<��H<ԱA<�:<Ӊ3<a{,<Vq%<�k<�k<�p<�{	<W�<�J�;*��;���; 4�;&��;w!�;��;XW�;��;g�{;�{a;�kG;2�-;�;?��:���:���:��;:�u�9�O��չ��J��%��Tlĺ�;����,�'��p>���T��"k�����o��)/��'Р��Q��R�������*ʻ<!Ի�޻���xy�P���9����v{��� ��C���T��!� �%��)*�LW.�\x2��6�H�:���>�߅B�mF��IJ� N�-�Q���U�tWY�X]�!�`��@d���g��\k��n��Yr���u�v:y���|�O ��1���0W��e��������D���䉼������������L���ᑼ'u�������%��ⲙ��>���ɜ�IS��ܟ��c���ꢼq��q���l{������ც����銭���,���3��;���s��ɝ��s!��r����)������4���  �  �dN==�M=o�L=7L=~TK=E�J=y�I=I=	<H=RtG=�F=��E=�E=�MD=�C="�B=`�A=�A=�H@=rw?=&�>=��==��<=_&<=�N;=mu:=��9=B�8=4�7=e 7=�6=J;5=�U4=ln3=�2=I�1=l�0=L�/=��.=��-=��,=��+=��*=��)=��(=��'=��&=��%=߾$=ӭ#=��"=�!=>g =I=e'===��=F�=\}=�I=a=A�=_�=�U==��=fv=5$=&�=5t=f
=��="O=��=�x=�=�=� =�<�<�=�<e7�<
*�<��<��<���<���<}��<=O�<�<��<s��<~D�<=��<
��<�D�<8��<���<u�<�<�@�<�͵<
W�<Rݮ<�`�<��<�^�<<ڠ<iS�<�ʙ<@�<곒<j&�<Ɨ�<�<�w�<��<R�z<��s<$fl<-De<K#^<�W<,�O<��H<�A<�:<̉3<^{,<Mq%<�k<�k<�p<�{	<&�<�J�;��;���;/4�;��;N!�;���;�W�;��;g�{;{{a;kG;�-;C�;���:=��:{��:1�;:"v�9F2�bչ�J�
&���kĺ-<����'��p>���T��"k������n���.���Ϡ��Q��W�������ʻE!Ի޻���y�S���9����s{�����G���T��!��%�**�hW.�ex2�%�6�4�:���>��B�"mF��IJ��N��Q���U�zWY�K]�9�`��@d���g��\k���n��Yr���u�c:y���|�J ��4���1W��b�����D���䉼������������L���ᑼ+u����������%��ײ���>���ɜ�cS��ܟ��c���ꢼ�p��w���n{������փ��w��㊭���,���/��G���q��՝��r!��o����)������4���  �  �eN=��M=�L=L=�VK=w�J=��I=�I=�>H=swG=8�F=7�E=nE=�QD=.�C=��B=)�A=�A=�M@=}?=�>=��====-<=�U;=�|:=P�9=:�8=w�7=�7=�'6=�D5=_4=hx3=>�2=��1=t�0=��/=��.=�-=��,=[�+=�*=*�)=o�(=��'=N�&=��%=1�$=|�#=��"=]�!=�w =�Y=�8=�=/�=$�=k�=�[=�$=��=$�=�h="=��=q�=J7=7�=8�=S)
=��=�a=_�=�=�=�=g, =;`�<p`�<mY�<�K�<�6�<�<���<6��<?��<$l�<1�<1��<é�<�]�<��<|��<T[�<���<[��<�.�<L¼<�Q�<�ݵ<Hf�<��<�m�<"�<�i�<�<Q\�<tҙ<�F�<���<+�<H��<�
�<0y�<>�<��z<�s<�`l<n<e<�^<��V<	�O<��H<��A<��:<fs3<�b,<�V%<4O<�L<�O<	Y	<Mh<���;=7�;���;"��;D�;t��;<M�;�;I��;��z;�`;�zF;��,;K�;���:Aܿ:K��:�H7:w��9͛]�B޹҆O�*�����ƺ����U���(���?�J*V�gl�[2��%���Җ��s��W����W������3�ʻ��Իa�޻o軗򻔡����S.���aQ�~���;������!�m4&�-m*�!�.���2�:�6���:���>�i�B�2�F�X�J�RN��R���U�(�Y�H3]���`��md�5�g�ˆk��o�@�r���u�_y���|�C��}����f��m��_����R����W����(��2����W��@쑼��F��ܟ���-��ʺ��JF���М��Y��⟼{i��𢼴u������U��\������9
��2���������K��	������ѝ��� �������(����� 2���  �  �eN=��M=�L=L=�VK=��J=��I=�I=�>H=iwG=5�F=9�E=kE=�QD=3�C=��B=%�A=�A=�M@=}?=�>=��====-<=�U;=�|:=J�9=<�8=��7=	7=�'6=�D5=y_4=fx3=?�2=��1=w�0=��/=��.=�-=��,=c�+=#�*=,�)=h�(=��'=K�&=��%=/�$=p�#=��"=S�!=�w =�Y=�8=�=4�='�=l�=\=�$=��=�=�h="=��=r�=E7=6�==�=\)
=��=�a=f�=�=�=�=f, =8`�<c`�<yY�<�K�<�6�<�<���<.��<8��<'l�<1�<@��<���<�]�<��<h��<X[�<���<d��<�.�<U¼<�Q�<�ݵ<Gf�<x�<�m�<�<�i�<.�<I\�<nҙ<�F�<���<+�<V��<�
�<7y�<@�<�z<�s<�`l<y<e<v^<��V<�O<�H<��A<Ӈ:<os3<�b,<�V%<,O<�L<�O<�X	<Ah<���;!7�;���;
��;.D�;���;ZM�;��;R��;L�z;��`;�zF;�,;��;0��:;ܿ:���:2G7:җ�9�z]��>޹K�O�����v�ƺ����N�<�(���?��*V��fl�I2����xҖ��s��M����W������E�ʻ��Իp�޻xo���������P.����PQ�l���;������!��4&�Jm*�L�.�ϸ2��6���:���>�~�B�5�F�E�J��QN��R���U��Y�^3]���`��md�:�g�҆k��o�)�r���u��^y���|�<�������f��j��X����R����d����(��G����W��C쑼��:��ԟ���-��ź��KF���М��Y��*⟼si����u������b��X���+
��6����������U��������˝��!�������(�����2���  �  �eN=��M=	�L=	L=�VK=~�J=��I=�I=�>H=mwG=9�F=;�E=fE=�QD=0�C=��B= �A=�A=�M@=}?=�>=��====-<=�U;=�|:=K�9=;�8=w�7=�7=�'6=�D5=y_4=kx3=@�2=�1=|�0=��/=��.=�-=��,=Z�+=�*=-�)=j�(=��'=H�&=��%=0�$=w�#=��"=U�!=�w =�Y=�8=�=0�="�=g�=\=�$=��="�=�h="=��=t�=F7=6�=7�=R)
=��=�a=h�=	�=�=�=f, =D`�<b`�<}Y�<tK�<�6�<�<���</��<<��<'l�<1�<?��<���<�]�<��<n��<`[�<���<]��<�.�<P¼<�Q�<�ݵ<Of�<�<�m�<	�<�i�<,�<C\�<zҙ<�F�<���<�*�<I��<�
�<5y�<A�<�z<8�s<k`l<�<e<~^<��V<�O<n�H<��A<��:<os3<�b,<�V%<#O<�L<�O<�X	<gh<���;F7�;���;���;D�;���;@M�;��;t��;��z;�`;Q{F;�,;��;���:%ܿ:���:�G7:0��9֞]��A޹��O�v���w�ƺU���4���(�E�?��*V��fl�l2��N���Җ��s��C����W��i���]�ʻ��Իc�޻@o�i�С����c.���\Q�z���;�����!��4&� m*�(�.�Ǹ2��6���:���>�{�B�3�F�^�J�RN��R���U��Y�h3]���`��md�8�g���k��o�!�r���u�_y��|�C�������f��j��b����R����Q����(��?����W��M쑼��A��ٟ��	.��Ǻ��CF���М��Y��(⟼ti����u������\��W������8
��>����������R�������������!�������(�����!2���  �  �eN=��M=�L=L=�VK=�J=��I=�I=�>H=lwG=6�F=8�E=qE=�QD=1�C=��B=*�A=�A=�M@=}?=��>=��====-<=�U;=�|:=M�9=<�8={�7=	7=�'6=�D5=}_4=fx3==�2=��1=v�0=��/=��.=�-=�,=`�+=�*=*�)=l�(=��'=O�&=��%=0�$=x�#=��"=W�!=�w =�Y=�8=�=2�=&�=n�=�[=�$=��=�=�h="=��=o�=G7=5�=;�=X)
=��=�a=a�=�=�=�=d, =8`�<j`�<qY�<�K�<�6�<�<���<2��<=��<#l�<1�<5��<���<�]�<��<r��<T[�<���<`��<�.�<Q¼<�Q�<�ݵ<Ef�<��<�m�<�<�i�<+�<O\�<qҙ<�F�<���<+�<Q��<�
�<1y�<>�<�z<�s<�`l<u<e<w^<��V<
�O<��H<��A<��:<fs3<�b,<�V%<1O<�L<�O<�X	<(h<���;,7�;���;7��;D�;���;GM�;�;H��;��z;��`;zzF;��,;c�;K��:ܿ:I��:�G7:���9��]��>޹I�O� �����ƺ���j�W�(���?��*V��fl�U2������Җ��s��]����W������)�ʻ��Իe�޻8o���ȡ����N.����WQ�t���;�����!��4&�Km*�5�.���2�-�6���:���>�u�B�8�F�M�J�RN��R���U��Y�^3]���`��md�>�g�Іk��o�8�r���u��^y���|�=�������f��n��V����R����f����(��=����W��;쑼��?��؟���-��ɺ��NF���М��Y��⟼{i����u������X��]������0
��&��� ������S��������͝��!�������(�����2���  �  �eN=��M=�L=L=�VK=��J=��I=�I=�>H=vwG=4�F=7�E=nE=�QD=6�C=��B=+�A=�A=�M@=}?=�>=��====-<=�U;=�|:=M�9=:�8=}�7=�7=�'6=�D5=�_4=ex3=@�2=��1=s�0=��/=��.=�-=��,=[�+="�*=(�)=q�(=��'=O�&=��%=0�$={�#=��"=]�!=�w =�Y=�8=�=5�=!�=p�=�[=�$=��=!�=�h="=��=k�=M7=4�=<�=U)
=��=�a=d�=�=�=	�=h, =3`�<t`�<pY�<|K�<�6�<�<���<0��<A��<l�<1�<+��<ȩ�<�]�<��<s��<M[�<���<T��<�.�<J¼<�Q�<�ݵ<Af�<��<�m�< �<�i�<*�<K\�<jҙ<�F�<���<+�<B��<�
�<-y�<G�<��z<�s<�`l<y<e<^<��V<�O<~�H<��A<ԇ:<]s3<�b,<�V%<(O<�L<�O<Y	<3h<���;7�;���;&��;�C�;���; M�;�;,��;��z;�`;�zF;��,;�;���:�ۿ:R��:�G7:Ɩ�9�]�HC޹��O�L���k�ƺ���2���(�ְ?�:*V��fl�i2��7���Җ��s��n���wW������'�ʻ��Իg�޻!o軲򻒡����F.���UQ�h���;�����!�s4&�:m*�*�.���2�:�6���:���>�_�B�>�F�I�J�RN��R���U��Y�C3]���`��md�/�g�ۆk��o�;�r���u�_y���|�?�������f��x��Q����R����^����(��;����W��9쑼��5��ߟ���-��Ǻ��QF���М��Y��⟼}i����u������S��a��솪�@
��5���������N��������˝��!�������(�����)2���  �  �eN=��M=	�L=L=�VK=}�J=��I=�I=�>H=lwG=4�F=?�E=iE=�QD=6�C=��B=%�A=�A=�M@=}?=�>=��====-<=�U;=�|:=J�9=:�8={�7=	7=�'6=�D5=w_4=fx3=B�2=�1=z�0=��/=��.=�-=��,=_�+=!�*=(�)=k�(=��'=L�&=��%=.�$=u�#=��"=S�!=�w =�Y=�8=�=4�= �=n�=\=�$=��=�=�h=
"=��=r�=H7=4�=:�=X)
=��=�a=e�=�=�=�=g, =9`�<^`�<xY�<�K�<�6�<�<���<,��<@��<#l�<1�<2��<���<�]�<��<h��<e[�<���<V��<�.�<O¼<�Q�<�ݵ<Ff�<|�<�m�<�<�i�<&�<H\�<uҙ<�F�<���<	+�<K��<�
�<8y�<<�<�z<5�s<l`l<�<e<q^<��V<�O<��H<��A<ʇ:<`s3<�b,<�V%<'O<�L<�O<�X	<Oh<���;7�;��;���;D�;���;.M�;��;���;O�z;��`;�zF;&�,;M�;P��:ܿ:���:$G7:���9��]��?޹چO�������ƺ��� ���(�h�?��*V��fl�V2�����Җ��s��j����W������<�ʻ��Իu�޻Qo軥�������@.���RQ�k���;�����!��4&�<m*�:�.�˸2�2�6���:���>�s�B�?�F�N�J�RN��R���U��Y�m3]���`��md�5�g�Άk��o�+�r���u��^y���|�@�������f��n��V����R����]����(��F����W��C쑼��7��ٟ��.������MF���М��Y��#⟼wi����u������[��_��򆪼6
��-����������X�������������
!�������(�����2���  �  �eN=��M=�L=L=�VK=z�J=��I=�I=�>H=iwG=7�F=8�E=iE=�QD=+�C=��B=�A=�A=�M@=}?=�>=��====-<=�U;=�|:=L�9=?�8=x�7=	7=�'6=�D5=x_4=fx3=C�2=�1=~�0=��/=��.=��-=��,=_�+=�*=-�)=h�(=��'=K�&=��%=2�$=u�#=��"=R�!=�w =�Y=�8=�=/�=)�=f�=\=�$=��=�=�h="=��=u�=D7=8�=9�=V)
=��=�a=h�=�=�= �=h, =<`�<``�<|Y�<tK�<�6�<
�<���<1��<:��<,l�<1�<>��<���<�]�<��<f��<`[�<���<o��<�.�<Z¼<�Q�<�ݵ<Mf�<w�<�m�<�<�i�<#�<L\�<vҙ<�F�<���<�*�<Q��<�
�</y�<A�<֩z<A�s<k`l<�<e<d^<��V<�O<q�H<��A<��:<zs3<�b,<�V%<2O<�L<�O<�X	<\h<���;57�;���;���;HD�;b��;�M�;��;j��;[�z;��`;{F;#�,;��;���:�ܿ:C��:�G7:�9ؘ]��=޹ňO�������ƺ��� ���(��?��*V�vfl��2�� ���Җ��s��@����W��f���C�ʻ��ԻV�޻Oo軁������b.����VQ�{��~;�����!��4&�-m*�7�.�¸2�"�6���:���>���B�,�F�S�J�RN��R���U� �Y�r3]���`��md�1�g�Ȇk��o�#�r���u��^y���|�:�������f��e��_����R����Z����(��H����W��O쑼��H��ϟ�� .��̺��FF���М��Y��&⟼ki����u������_��R������1
��7���������`��󗳼�������!�������(�����2���  �  �eN=��M=�L=L=�VK=z�J=��I=�I=�>H=pwG=:�F=6�E=kE=�QD=+�C=��B=#�A=�A=�M@=}?=�>=��====-<=�U;=�|:=L�9=9�8=y�7= 	7=�'6=�D5=�_4=cx3=?�2=��1=r�0=��/=��.= �-=��,=^�+=�*=(�)=m�(=��'=O�&=��%=0�$=w�#=��"=X�!=�w =�Y=�8=�=0�=&�=g�=\=�$=��= �=�h=
"=��=q�=H7=3�=8�=U)
=��=�a=g�=�=�=�=g, =2`�<q`�<vY�<wK�<�6�<
�<���</��<:��<&l�<1�<2��<���<�]�<��<q��<Y[�<���<f��<�.�<U¼<�Q�<�ݵ<Of�<��<�m�<�<�i�<!�<Q\�<oҙ<�F�<���<+�<N��<�
�<,y�<L�<�z<�s<�`l<w<e<n^<��V<�O<{�H<��A<��:<_s3<�b,<�V%<:O<�L<�O<�X	<Jh<���;I7�;���;��;5D�;c��;gM�;��;T��;��z;�`;�zF;n�,;U�;���:Uܿ:��:�G7:��9��]�i@޹:�O�������ƺS���A�1�(��?��*V�]fl�{2��/���Җ��s��j����W������)�ʻ��Իf�޻>o軏򻻡�����c.���WQ�z���;�����!��4&�.m*�/�.���2�3�6���:���>�t�B�>�F�Y�J�RN��R���U��Y�U3]���`��md�4�g�݆k��o�/�r���u�_y���|�D�������f��k��Z����R����\����(��=����W��J쑼��G��ӟ���-��Ϻ��CF���М��Y��⟼vi����u������U��a������4
��5���������V��������̝��!�������(�����2���  �  �eN=��M=�L=L=�VK=~�J=��I=�I=�>H=mwG=2�F=>�E=mE=�QD=9�C=��B=)�A=�A=�M@=}?=�>=��====-<=�U;=�|:=M�9=6�8=��7=�7=�'6=�D5=|_4=fx3==�2=��1=r�0=��/=��.=�-=��,=_�+=%�*=$�)=o�(=��'=P�&=��%=1�$=w�#=��"=U�!=�w =�Y=�8=�=6�= �=r�= \=�$=��=�=�h=
"=��=k�=J7=1�==�=Y)
=��=�a=^�=�=�=�=e, =6`�<k`�<hY�<�K�<�6�<�<���<.��<?��<l�<1�<1��<©�<�]�<��<k��<^[�<���<W��<�.�<Q¼<�Q�<�ݵ<Bf�<��<�m�<�<�i�<(�<K\�<jҙ<�F�<���<+�<E��<�
�<3y�<4�<��z<�s<�`l<k<e<�^<��V<�O<��H<��A<߇:<Ks3<�b,<�V%<(O<�L<�O<�X	<2h<���;7�;؀�;��;D�;п�;*M�;�;w��;Z�z;��`;�zF;��,;E�;���:�ۿ:T��:
H7:���9�r]��B޹-�O�u���"�ƺ���g��(��?�@*V�gl�C2�����Җ��s�������W�������ʻ��Ի_�޻Ao���ѡ����9.���KQ�b���;�����!��4&�Fm*�8�.���2�2�6���:���>�i�B�I�F�B�J�RN��R���U�+�Y�I3]���`��md�:�g�Ԇk��o�I�r�n�u�_y���|�C�������f��v��O����R����d����(��C����W��9쑼��0��ן���-������QF���М��Y��⟼ui����u������O��j��熪�=
��'����������K��������ҝ��!�������(�����(2���  �  �eN=��M=�L=L=�VK=}�J=��I=�I=�>H=twG=5�F=;�E=lE=�QD=1�C=��B=&�A=�A=�M@=}?=�>=��====-<=�U;=�|:=O�9=8�8=}�7=�7=�'6=�D5=z_4=kx3=@�2=��1=x�0=��/=��.=�-=��,=[�+=!�*=)�)=m�(=��'=M�&=��%=1�$=w�#=��"=Y�!=�w =�Y=�8=�=2�=#�=l�=�[=�$=��= �=�h="=��=o�=I7=5�=;�=U)
=��=�a=b�=�=�=�=f, =@`�<g`�<qY�<}K�<�6�<�<���<1��<@��<"l�<1�<6��<���<�]�<��<p��<T[�<���<]��<�.�<J¼<�Q�<�ݵ<Ef�<��<�m�<�<�i�<'�<L\�<qҙ<�F�<���<+�<>��<�
�<5y�<;�<��z<%�s<�`l<}<e<�^<��V<�O<y�H<~�A<҇:<Zs3<�b,<�V%</O<�L<�O<�X	<Vh<���;#7�;���;��;D�;���;>M�;��;Q��;{�z;+�`;{F;H�,;s�;'��:#ܿ:���:[H7:���9�]�	D޹u�O�6���L�ƺR���:�a�(���?�X*V��fl�U2��H���Җ��s��_����W������6�ʻ��Ի\�޻Ao�r򻲡����O.�	��ZQ�s���;������!��4&�m*�0�.���2�+�6���:���>�n�B�:�F�K�J�RN��R���U��Y�R3]���`��md�7�g�k��o�9�r���u�_y���|�A�������f��n��Y����R����X����(��>����W��C쑼��>��ޟ���-��º��MF���М��Y�� ⟼qi����u������U��_���D
��9����������K��������ɝ��� �������(�����-2���  �  �eN=��M=�L=L=�VK={�J=��I=�I=�>H=iwG=9�F=8�E=nE=�QD=+�C=��B=&�A=�A=�M@=
}?=�>=��====-<=�U;=�|:=P�9=:�8=w�7=	7=�'6=�D5=z_4=ax3=?�2=��1=v�0=��/=��.=�-=��,=c�+=�*=.�)=g�(=��'=L�&=��%=.�$=q�#=��"=R�!=�w =�Y=�8=�=0�=)�=h�=\=�$=��=�=�h="=��=t�=C7=9�=8�=[)
=��=�a=h�=�=�=�=e, =1`�<``�<}Y�<{K�<�6�<�<���<6��<3��<,l�<1�<<��<���<�]�<��<m��<_[�<���<i��<�.�<S¼<�Q�<�ݵ<Of�<w�<�m�<
�<�i�<#�<Q\�<qҙ<�F�<���<�*�<Z��<�
�<5y�<E�<֩z<!�s<�`l<|<e<_^<��V<�O<��H<��A<��:<ns3<�b,<�V%<@O<�L<�O<�X	<Ah<���;E7�;���;&��;2D�;c��;oM�;��;k��;��z;h�`;�zF;�,;��;ܐ�:�ܿ:���:�H7:䖨9��]�=޹؇O�s���]�ƺ����E�u�(���?��*V�yfl�b2����sҖ��s��8����W��z���A�ʻ��Իt�޻ko軴������].����YQ�y��};�����!��4&�Fm*�G�.�͸2�+�6���:���>���B�*�F�Y�J��QN��R���U���Y�q3]���`��md�<�g�ކk��o�!�r���u��^y���|�?��|����f��e��]����R����c����(��A����W��G쑼	��G��֟���-��ɺ��DF���М��Y��'⟼pi����u������^��T�����'
��0����������`��������ɝ��!�������(�����2���  �  �eN=��M=�L=L=�VK=y�J=��I=�I=�>H=mwG=9�F=8�E=lE=�QD=3�C=��B=%�A=�A=�M@=}?=�>=��====-<=�U;=�|:=Q�9=;�8=u�7=�7=�'6=�D5=|_4=fx3=A�2=��1=z�0=��/=��.= �-=��,=Z�+=�*=.�)=l�(=��'=K�&=��%=2�$=|�#=��"=X�!=�w =�Y=�8=�=2�=#�=k�=\=�$=��=$�=�h="=��=r�=G7=9�=6�=Q)
=��=�a=d�=�=�=�=g, =;`�<h`�<tY�<wK�<�6�< �<���<8��<8��<"l�<
1�<:��<é�<�]�<��<s��<][�<���<]��<�.�<N¼<�Q�<�ݵ<Of�<��<�m�<�<�i�<!�<H\�<sҙ<�F�<���<�*�<H��<�
�<.y�<=�<�z<-�s<�`l<�<e<q^<��V<�O<p�H<��A<��:<os3<�b,<�V%<(O<�L<�O<�X	<Xh<���;G7�;���;��;D�;���;:M�;��;i��;��z;��`;>{F;��,;��;���:ܿ:��:�H7:��9ӣ]�B޹��O���ƺ����?�(�c�?��*V��fl�}2��J���Җ��s��8����W��}���I�ʻ��ԻR�޻o軈򻽡�����Z.�
��YQ�q���;������!��4&�/m*��.���2�+�6���:���>�v�B�)�F�_�J�#RN��R���U��Y�\3]���`��md�2�g�ʆk��o�2�r���u�_y��|�A��y����f��n��`����R����S����(��;����W��D쑼��9��ڟ���-��ɺ��DF���М��Y��⟼oi����u������V��T�����9
��:���������U���������ĝ��
!�������(�����!2���  �  �eN=��M=�L=L=�VK=��J=��I=�I=�>H=pwG=5�F=;�E=oE=�QD=;�C=��B=*�A=�A=�M@=}?=�>=��====-<=�U;=�|:=G�9=7�8=��7=	7=�'6=�D5=z_4=gx3==�2=�1=u�0=��/=��.=�-=��,=b�+=#�*='�)=i�(=��'=N�&=��%=.�$=s�#=��"=X�!=�w =�Y=�8=�=5�=#�=q�=�[=�$=��=�=�h="=��=p�=F7=1�=<�=[)
=��=�a=a�=�=�= �=c, =;`�<f`�<pY�<�K�<�6�<�<���<)��<>��<&l�<1�<6��<���<�]�<��<n��<R[�<���<Y��<�.�<K¼<�Q�<�ݵ<Ff�<��<�m�<
�<�i�<.�<K\�<sҙ<�F�<���<+�<M��<�
�<<y�<9�<��z< �s<w`l<{<e<�^<��V<�O<��H<��A<�:<Vs3<�b,<�V%</O<�L<�O<�X	<Ch<���;$7�;���;/��;�C�;޿�;*M�;�;P��;o�z;ƒ`;�zF;)�,;w�;]��:Kܿ:���:zF7:V��9�m]��?޹�O����c�ƺ����k���(���?��*V��fl�'2����Җ��s��u����W������+�ʻ��Իt�޻`o軻򻼡����?.���RQ�e���;�����!��4&�=m*�A�.�ɸ2�#�6���:���>�z�B�H�F�F�J��QN��R���U��Y�_3]���`��md�C�g�ˆk��o�;�r�s�u�_y���|�A�������f��k��R����R����d����(��@����W��:쑼��.��ݟ���-������MF���М��Y��&⟼ui����u������a��a��ꆪ�4
��-����������M��������ʝ��!�������(�����2���  �  �eN=��M=�L=L=�VK=y�J=��I=�I=�>H=mwG=9�F=8�E=lE=�QD=3�C=��B=%�A=�A=�M@=}?=�>=��====-<=�U;=�|:=Q�9=;�8=u�7=�7=�'6=�D5=|_4=fx3=A�2=��1=z�0=��/=��.= �-=��,=Z�+=�*=.�)=l�(=��'=K�&=��%=2�$=|�#=��"=X�!=�w =�Y=�8=�=2�=#�=k�=\=�$=��=$�=�h="=��=r�=G7=9�=6�=Q)
=��=�a=d�=�=�=�=g, =;`�<h`�<tY�<wK�<�6�< �<���<8��<8��<"l�<
1�<:��<é�<�]�<��<s��<][�<���<]��<�.�<N¼<�Q�<�ݵ<Of�<��<�m�<�<�i�<!�<H\�<sҙ<�F�<���<�*�<H��<�
�<.y�<=�<�z<-�s<�`l<�<e<q^<��V<�O<p�H<��A<��:<os3<�b,<�V%<(O<�L<�O<�X	<Xh<���;G7�;���;��;D�;���;:M�;��;i��;��z;��`;>{F;��,;��;���:ܿ:��:�H7:��9֣]�B޹��O���ƺ����?�(�c�?��*V��fl�}2��J���Җ��s��8����W��}���J�ʻ��ԻR�޻o軈򻽡�����Z.�
��YQ�q���;������!��4&�/m*��.���2�+�6���:���>�v�B�)�F�_�J�#RN��R���U��Y�\3]���`��md�2�g�ʆk��o�2�r���u�_y��|�A��y����f��n��`����R����S����(��;����W��D쑼��9��ڟ���-��ɺ��DF���М��Y��⟼oi����u������V��T�����9
��:���������U���������ĝ��
!�������(�����!2���  �  �eN=��M=�L=L=�VK={�J=��I=�I=�>H=iwG=9�F=8�E=nE=�QD=+�C=��B=&�A=�A=�M@=
}?=�>=��====-<=�U;=�|:=P�9=:�8=w�7=	7=�'6=�D5=z_4=ax3=?�2=��1=v�0=��/=��.=�-=��,=c�+=�*=.�)=g�(=��'=L�&=��%=.�$=q�#=��"=R�!=�w =�Y=�8=�=0�=)�=h�=\=�$=��=�=�h="=��=t�=C7=9�=8�=[)
=��=�a=h�=�=�=�=e, =1`�<``�<}Y�<{K�<�6�<�<���<6��<3��<,l�<1�<<��<���<�]�<��<m��<_[�<���<i��<�.�<S¼<�Q�<�ݵ<Of�<w�<�m�<
�<�i�<#�<Q\�<qҙ<�F�<���<�*�<Z��<�
�<5y�<E�<֩z<!�s<�`l<|<e<_^<��V<�O<��H<��A<��:<ns3<�b,<�V%<@O<�L<�O<�X	<Ah<���;E7�;���;&��;2D�;c��;oM�;��;k��;��z;h�`;�zF;�,;��;ܐ�:�ܿ:���:�H7:㖨9��]�=޹؇O�s���]�ƺ����E�u�(���?��*V�yfl�c2����sҖ��s��8����W��z���A�ʻ��Իt�޻ko軴������].����YQ�y��};�����!��4&�Fm*�G�.�͸2�+�6���:���>���B�*�F�Y�J��QN��R���U���Y�q3]���`��md�<�g�ކk��o�!�r���u��^y���|�?��|����f��e��]����R����c����(��A����W��G쑼	��G��֟���-��ɺ��DF���М��Y��'⟼pi����u������^��T�����'
��0����������`��������ɝ��!�������(�����2���  �  �eN=��M=�L=L=�VK=}�J=��I=�I=�>H=twG=5�F=;�E=lE=�QD=1�C=��B=&�A=�A=�M@=}?=�>=��====-<=�U;=�|:=O�9=8�8=}�7=�7=�'6=�D5=z_4=kx3=@�2=��1=x�0=��/=��.=�-=��,=[�+=!�*=)�)=m�(=��'=M�&=��%=1�$=w�#=��"=Y�!=�w =�Y=�8=�=2�=#�=l�=�[=�$=��= �=�h="=��=o�=I7=5�=;�=U)
=��=�a=b�=�=�=�=f, =@`�<g`�<qY�<}K�<�6�<�<���<1��<@��<"l�<1�<6��<���<�]�<��<p��<T[�<���<]��<�.�<J¼<�Q�<�ݵ<Ef�<��<�m�<�<�i�<'�<L\�<qҙ<�F�<���<+�<>��<�
�<5y�<;�<��z<%�s<�`l<}<e<�^<��V<�O<y�H<~�A<҇:<Zs3<�b,<�V%</O<�L<�O<�X	<Vh<���;#7�;���;��;D�;���;>M�;��;Q��;{�z;+�`;{F;H�,;s�;'��:"ܿ:���:ZH7:���9�]�D޹v�O�6���L�ƺS���;�a�(���?�X*V��fl�U2��H���Җ��s��_����W������6�ʻ��Ի\�޻Ao�r򻲡����O.�	��ZQ�s���;������!��4&�m*�0�.���2�+�6���:���>�n�B�:�F�K�J�RN��R���U��Y�R3]���`��md�7�g�k��o�9�r���u�_y���|�A�������f��n��Y����R����X����(��>����W��C쑼��>��ޟ���-��º��MF���М��Y�� ⟼qi����u������U��_���D
��9����������K��������ɝ��� �������(�����-2���  �  �eN=��M=�L=L=�VK=~�J=��I=�I=�>H=mwG=2�F=>�E=mE=�QD=9�C=��B=)�A=�A=�M@=}?=�>=��====-<=�U;=�|:=M�9=6�8=��7=�7=�'6=�D5=|_4=fx3==�2=��1=r�0=��/=��.=�-=��,=_�+=%�*=$�)=o�(=��'=P�&=��%=1�$=w�#=��"=U�!=�w =�Y=�8=�=6�= �=r�= \=�$=��=�=�h=
"=��=k�=J7=1�==�=Y)
=��=�a=^�=�=�=�=e, =6`�<k`�<hY�<�K�<�6�<�<���<.��<?��<l�<1�<1��<©�<�]�<��<k��<^[�<���<W��<�.�<Q¼<�Q�<�ݵ<Bf�<��<�m�<�<�i�<(�<K\�<jҙ<�F�<���<+�<E��<�
�<3y�<4�<��z<�s<�`l<k<e<�^<��V<�O<��H<��A<߇:<Ks3<�b,<�V%<(O<�L<�O<�X	<2h<���;7�;؀�;��;D�;п�;*M�;�;w��;Y�z;��`;�zF;��,;E�;���:�ۿ:T��:	H7:���9�r]��B޹.�O�v���"�ƺ���g��(��?�@*V�gl�C2�����Җ��s�������W�������ʻ��Ի_�޻Bo���ѡ����9.���KQ�b���;�����!��4&�Fm*�8�.���2�2�6���:���>�i�B�I�F�B�J�RN��R���U�+�Y�I3]���`��md�:�g�Ԇk��o�I�r�n�u�_y���|�C�������f��v��O����R����d����(��C����W��9쑼��0��ן���-������QF���М��Y��⟼ui����u������O��j��熪�=
��'����������K��������ҝ��!�������(�����(2���  �  �eN=��M=�L=L=�VK=z�J=��I=�I=�>H=pwG=:�F=6�E=kE=�QD=+�C=��B=#�A=�A=�M@=}?=�>=��====-<=�U;=�|:=L�9=9�8=y�7= 	7=�'6=�D5=�_4=cx3=?�2=��1=r�0=��/=��.= �-=��,=^�+=�*=(�)=m�(=��'=O�&=��%=0�$=w�#=��"=X�!=�w =�Y=�8=�=0�=&�=g�=\=�$=��= �=�h=
"=��=q�=H7=3�=8�=U)
=��=�a=g�=�=�=�=g, =2`�<q`�<vY�<wK�<�6�<
�<���</��<:��<&l�<1�<2��<���<�]�<��<q��<Y[�<���<f��<�.�<U¼<�Q�<�ݵ<Of�<��<�m�<�<�i�<!�<Q\�<oҙ<�F�<���<+�<N��<�
�<,y�<L�<�z<�s<�`l<w<e<n^<��V<�O<{�H<��A<��:<_s3<�b,<�V%<:O<�L<�O<�X	<Jh<���;I7�;���;��;4D�;c��;gM�;��;T��;��z;�`;�zF;n�,;T�;���:Uܿ:��:�G7:��9Ɠ]�k@޹;�O�������ƺS���B�1�(��?��*V�]fl�{2��/���Җ��s��j����W������)�ʻ��Իf�޻>o軏򻻡�����c.���WQ�z���;�����!��4&�.m*�/�.���2�3�6���:���>�t�B�>�F�Y�J�RN��R���U��Y�U3]���`��md�4�g�݆k��o�/�r���u�_y���|�D�������f��k��Z����R����\����(��=����W��J쑼��G��ӟ���-��Ϻ��CF���М��Y��⟼vi����u������U��a������4
��5���������V��������̝��!�������(�����2���  �  �eN=��M=�L=L=�VK=z�J=��I=�I=�>H=iwG=7�F=8�E=iE=�QD=+�C=��B=�A=�A=�M@=}?=�>=��====-<=�U;=�|:=L�9=?�8=x�7=	7=�'6=�D5=x_4=fx3=C�2=�1=~�0=��/=��.=��-=��,=_�+=�*=-�)=h�(=��'=K�&=��%=2�$=u�#=��"=R�!=�w =�Y=�8=�=/�=)�=f�=\=�$=��=�=�h="=��=u�=D7=8�=9�=V)
=��=�a=h�=�=�= �=h, =<`�<``�<|Y�<tK�<�6�<
�<���<1��<:��<,l�<1�<>��<���<�]�<��<f��<`[�<���<o��<�.�<Z¼<�Q�<�ݵ<Mf�<w�<�m�<�<�i�<#�<L\�<vҙ<�F�<���<�*�<Q��<�
�</y�<A�<֩z<A�s<k`l<�<e<d^<��V<�O<q�H<��A<��:<zs3<�b,<�V%<2O<�L<�O<�X	<\h<���;57�;���;���;HD�;b��;�M�;��;j��;[�z;��`;{F;#�,;��;���:�ܿ:C��:�G7:9�]��=޹ƈO�������ƺ��� ���(��?��*V�vfl��2�� ���Җ��s��@����W��f���C�ʻ��ԻV�޻Oo軁������b.����VQ�{��~;�����!��4&�-m*�7�.�¸2�"�6���:���>���B�,�F�S�J�RN��R���U� �Y�r3]���`��md�1�g�Ȇk��o�#�r���u��^y���|�:�������f��e��_����R����Z����(��H����W��O쑼��H��ϟ�� .��̺��FF���М��Y��&⟼ki����u������_��R������1
��7���������`��󗳼�������!�������(�����2���  �  �eN=��M=	�L=L=�VK=}�J=��I=�I=�>H=lwG=4�F=?�E=iE=�QD=6�C=��B=%�A=�A=�M@=}?=�>=��====-<=�U;=�|:=J�9=:�8={�7=	7=�'6=�D5=w_4=fx3=B�2=�1=z�0=��/=��.=�-=��,=_�+=!�*=(�)=k�(=��'=L�&=��%=.�$=u�#=��"=S�!=�w =�Y=�8=�=4�= �=n�=\=�$=��=�=�h=
"=��=r�=H7=4�=:�=X)
=��=�a=e�=�=�=�=g, =9`�<^`�<xY�<�K�<�6�<�<���<,��<A��<#l�<1�<2��<���<�]�<��<h��<e[�<���<V��<�.�<O¼<�Q�<�ݵ<Ff�<|�<�m�<�<�i�<&�<H\�<uҙ<�F�<���<	+�<K��<�
�<8y�<<�<�z<5�s<l`l<�<e<q^<��V<�O<��H<��A<ʇ:<`s3<�b,<�V%<'O<�L<�O<�X	<Oh<���;7�;��;���;D�;���;.M�;��;���;O�z;��`;�zF;%�,;M�;P��:ܿ:���:#G7:���9Ɍ]��?޹ۆO�������ƺ��� ���(�h�?��*V��fl�V2�����Җ��s��j����W������<�ʻ��Իu�޻Qo軦�������@.���RQ�k���;�����!��4&�<m*�:�.�˸2�2�6���:���>�s�B�?�F�N�J�RN��R���U��Y�m3]���`��md�5�g�Άk��o�+�r���u��^y���|�@�������f��n��V����R����]����(��F����W��C쑼��7��ٟ��.������MF���М��Y��#⟼wi����u������[��_��򆪼6
��-����������X�������������
!�������(�����2���  �  �eN=��M=�L=L=�VK=��J=��I=�I=�>H=vwG=4�F=7�E=nE=�QD=6�C=��B=+�A=�A=�M@=}?=�>=��====-<=�U;=�|:=M�9=:�8=}�7=�7=�'6=�D5=�_4=ex3=@�2=��1=s�0=��/=��.=�-=��,=[�+="�*=(�)=q�(=��'=O�&=��%=0�$={�#=��"=]�!=�w =�Y=�8=�=5�=!�=p�=�[=�$=��=!�=�h="=��=k�=M7=4�=<�=U)
=��=�a=d�=�=�=	�=h, =3`�<t`�<pY�<|K�<�6�<�<���<0��<A��<l�<1�<+��<ȩ�<�]�<��<s��<M[�<���<T��<�.�<J¼<�Q�<�ݵ<Af�<��<�m�< �<�i�<*�<K\�<jҙ<�F�<���<+�<B��<�
�<-y�<G�<��z<�s<�`l<y<e<^<��V<�O<~�H<��A<ԇ:<]s3<�b,<�V%<(O<�L<�O<Y	<3h<���;7�;���;&��;�C�;���; M�;�;,��;��z;�`;�zF;��,;�;���:�ۿ:R��:�G7:Ė�9�]�IC޹��O�L���k�ƺ���3���(�ְ?�:*V��fl�i2��8���Җ��s��n���wW������'�ʻ��Իg�޻!o軲򻒡����F.���UQ�h���;�����!�s4&�:m*�*�.���2�:�6���:���>�_�B�>�F�I�J�RN��R���U��Y�C3]���`��md�/�g�ۆk��o�;�r���u�_y���|�?�������f��x��Q����R����^����(��;����W��9쑼��5��ߟ���-��Ǻ��QF���М��Y��⟼}i����u������S��a��솪�@
��5���������N��������˝��!�������(�����)2���  �  �eN=��M=�L=L=�VK=�J=��I=�I=�>H=lwG=6�F=8�E=qE=�QD=1�C=��B=*�A=�A=�M@=}?=��>=��====-<=�U;=�|:=M�9=<�8={�7=	7=�'6=�D5=}_4=fx3==�2=��1=v�0=��/=��.=�-=�,=`�+=�*=*�)=l�(=��'=O�&=��%=0�$=x�#=��"=W�!=�w =�Y=�8=�=2�=&�=n�=�[=�$=��=�=�h="=��=o�=G7=5�=;�=X)
=��=�a=a�=�=�=�=d, =8`�<j`�<qY�<�K�<�6�<�<���<2��<=��<#l�<1�<5��<���<�]�<��<r��<T[�<���<`��<�.�<Q¼<�Q�<�ݵ<Ef�<��<�m�<�<�i�<+�<O\�<qҙ<�F�<���<+�<Q��<�
�<1y�<>�<�z<�s<�`l<u<e<w^<��V<
�O<��H<��A<��:<fs3<�b,<�V%<1O<�L<�O<�X	<(h<���;,7�;���;7��;D�;���;GM�;�;H��;��z;��`;zzF;��,;c�;K��:ܿ:I��:�G7:���9��]��>޹J�O� �����ƺ���k�W�(���?��*V��fl�U2������Җ��s��]����W������)�ʻ��Իe�޻8o���ȡ����N.����WQ�t���;�����!��4&�Km*�5�.���2�-�6���:���>�u�B�8�F�M�J�RN��R���U��Y�^3]���`��md�>�g�Іk��o�8�r���u��^y���|�=�������f��n��V����R����f����(��=����W��;쑼��?��؟���-��ɺ��NF���М��Y��⟼{i����u������X��]������0
��&��� ������S��������͝��!�������(�����2���  �  �eN=��M=	�L=	L=�VK=~�J=��I=�I=�>H=mwG=9�F=;�E=fE=�QD=0�C=��B= �A=�A=�M@=}?=�>=��====-<=�U;=�|:=K�9=;�8=w�7=�7=�'6=�D5=y_4=kx3=@�2=�1=|�0=��/=��.=�-=��,=Z�+=�*=-�)=j�(=��'=H�&=��%=0�$=w�#=��"=U�!=�w =�Y=�8=�=0�="�=g�=\=�$=��="�=�h="=��=t�=F7=6�=7�=R)
=��=�a=h�=	�=�=�=f, =D`�<b`�<}Y�<tK�<�6�<�<���</��<<��<'l�<1�<?��<���<�]�<��<n��<`[�<���<]��<�.�<P¼<�Q�<�ݵ<Of�<�<�m�<�<�i�<,�<C\�<zҙ<�F�<���<�*�<I��<�
�<5y�<A�<�z<8�s<k`l<�<e<~^<��V<�O<n�H<��A<��:<os3<�b,<�V%<#O<�L<�O<�X	<gh<���;F7�;���;���;D�;���;@M�;��;t��;��z;�`;P{F;�,;��;���:$ܿ:���:�G7:/��9۞]��A޹��O�v���x�ƺU���5���(�E�?��*V��fl�l2��N���Җ��s��C����W��i���]�ʻ��Իc�޻@o�i�С����c.���\Q�z���;�����!��4&� m*�(�.�Ǹ2��6���:���>�{�B�3�F�^�J�RN��R���U��Y�h3]���`��md�8�g���k��o�!�r���u�_y��|�C�������f��j��b����R����Q����(��?����W��M쑼��A��ٟ��	.��Ǻ��CF���М��Y��(⟼ti����u������\��W������8
��>����������R�������������!�������(�����!2���  �  �eN=��M=�L=L=�VK=��J=��I=�I=�>H=iwG=5�F=9�E=kE=�QD=3�C=��B=%�A=�A=�M@=}?=�>=��====-<=�U;=�|:=J�9=<�8=��7=	7=�'6=�D5=y_4=fx3=?�2=��1=w�0=��/=��.=�-=��,=c�+=#�*=,�)=h�(=��'=K�&=��%=/�$=p�#=��"=S�!=�w =�Y=�8=�=4�='�=l�=\=�$=��=�=�h="=��=r�=E7=6�==�=\)
=��=�a=f�=�=�=�=f, =8`�<c`�<yY�<�K�<�6�<�<���<.��<8��<'l�<1�<@��<���<�]�<��<h��<X[�<���<d��<�.�<U¼<�Q�<�ݵ<Gf�<x�<�m�<�<�i�<.�<I\�<nҙ<�F�<���<+�<V��<�
�<7y�<@�<�z<�s<�`l<y<e<v^<��V<�O<�H<��A<Ӈ:<os3<�b,<�V%<,O<�L<�O<�X	<Ah<���;!7�;���;
��;/D�;���;ZM�;��;R��;L�z;��`;�zF;�,;��;0��:;ܿ:���:2G7:ї�9�z]��>޹K�O�����v�ƺ����N�<�(���?��*V��fl�I2����xҖ��s��M����W������E�ʻ��Իp�޻xo���������P.����PQ�l���;������!��4&�Jm*�L�.�ϸ2��6���:���>�~�B�5�F�E�J��QN��R���U��Y�^3]���`��md�:�g�҆k��o�)�r���u��^y���|�<�������f��j��X����R����d����(��G����W��C쑼��:��ԟ���-��ź��KF���М��Y��*⟼si����u������b��X���+
��6����������U��������˝��!�������(�����2���  �  @gN=H�M=��L=%L=�XK=�J=��I=�I=NBH={G=�F=l�E=� E=�VD=>�C=�B=��A=�#A=)T@=��?=�>=��==�
==5<=�];=n�:=Y�9=��8=D�7=&7=L26=�O5=�j4=2�3=p�2=��1=}�0=,�/=o�.=X�-=��,=��+=�+=1*=�)=��'=��&=u�%=G�$=��#=i�"=��!=f� =�m=�L=6(= =K�=֤=�q=�:=��=R�=�~=v8=8�=��=�M=��=ĝ=�?
=��=)x=t=��=�/=t�=�A =���<���<́�<(s�<o]�<A�<��<f��<z��<X��<HR�<P�<���<�{�<�)�<��<�u�<��<��<�E�<�׼<gf�<�<Cx�<M��<1}�<U��<�v�<��<�f�<�ۙ<�N�<L��<x0�<s��<��<�z�<��<i�z<��s<�Yl<Q3e<�^<��V<{�O<��H<��A<�o:<�X3<�E,<=7%<O-<k(<�(<�/	<�<<���; ��;��;�o�;�Կ;�K�;�Ԥ;&q�;!�;�y;_;�^E;l+;��;�(�:�d�:��:�"2:/�9�����&��U�nS����ɺ�����y��p*��+A���W���m���iӌ�d����5�� �������[��P~˻ �ջ|f߻�+黪��[�������v ����k$�!�����A"���&���*��.��3��7�x;��?��C���F��J��N��VR��V���Y�l]��a��d��1h���k��7o���r�I v�N�y���|�H%���Ё�Ry��1��[�c��E��G���7���Ύ��d������Ɗ��T��`����7��ę�O���؜��a��F韼"p�����V{��������������u��叭�?���������蘳�5��Ɲ��{ ������-'��)����/���  �  >gN=J�M=��L=$L=�XK=�J=��I=�I=QBH={G=#�F=m�E=� E=�VD=B�C=�B=��A=�#A=)T@=��?=�>=��==�
==5<=�];=k�:=V�9=��8=D�7=-7=I26=�O5=�j4=.�3=q�2=��1=~�0=%�/=r�.=U�-=��,=��+=�+=1*=�)=��'=��&={�%=M�$=��#=j�"=��!=l� =�m=�L==(= =K�=Ӥ=�q=�:=��=P�=�~=~8=7�= �=�M=��==�?
=��=&x=y=�=�/=t�=�A =��<x��<ҁ�<!s�<|]�<
A�<��<`��<o��<_��<JR�<b�<���<�{�<)�<��<�u�<��<���<�E�<ؼ<`f�<�<Lx�<B��<7}�<U��<�v�<��<�f�<�ۙ<�N�<P��<w0�<���<��<�z�<��<J�z<�s<�Yl<c3e<�^<��V<{�O<w�H<�A<�o:<�X3<�E,<87%<F-<p(<()<�/	<�<<���;;��;�;�o�;տ;�K�;�Ԥ;q�;!�;�y;�~_;�^E;�k+;F�; )�:e�:q�:�!2:��9�����"鹆U�4S��)�ɺW���iy��p*�o+A��W�[�m��Yӌ�6����5����� ���[��\~˻�ջOf߻�+黡��&[�������{ ����P$�����uA"���&���*��.��3��7�|;��?��C���F��J��N��VR��V���Y�(l]��a��d��1h���k��7o���r�V v�5�y���|�E%���Ё�\y��+��X�c��G��H���7���Ύ��d����������K��O����7��ę�O���؜��a��G韼p�����Z{�����������������d��鏭�@��|������☳�3������� ������-'��.����/���  �  <gN=P�M=��L=(L=�XK=�J=��I=�I=XBH={G=$�F=o�E=� E=�VD=8�C=�B=��A=�#A=(T@=��?=��>=��==�
==5<=�];=m�:=V�9=��8=A�7=/7=C26=�O5=�j4=/�3=u�2=��1=��0=%�/=z�.=R�-=��,=��+=�+=7*=�)=��'=��&=v�%=I�$=��#=n�"=��!=n� =�m=�L=9(= =L�=Ӥ=�q=�:=��=P�=�~=z8=2�=�=�M=��=ŝ=�?
=��="x=�=�=�/=r�=�A =���<{��<݁�<s�<]�<A�<��<f��<s��<i��<=R�<^�<���<�{�<�)�<��<�u�<��<���<�E�<
ؼ<^f�<�<Qx�<?��<E}�<M��<�v�<��<�f�<�ۙ<�N�<[��<t0�<���<��<�z�<��<G�z<�s<�Yl<y3e<�^<��V<�O<`�H< �A<�o:<�X3<�E,<K7%<I-<U(<)<�/	<�<<���;D��;�;�o�;տ;�K�;դ;q�;7!�;�y;�~_;�^E;�k+;%�;I(�:�e�:��:�!2:��9ך���!�+U��R��ǩɺ���3y�,q*�+A���W���m��iӌ�,����5��񶬻)��N[��w~˻�ջmf߻�+黀��?[�������x ����a$�����kA"���&���*��.��3��7��;��?��C���F��J��N��VR�V���Y�'l]��a��d��1h���k��7o���r�p v�.�y���|�;%���Ё�Yy��!��e�c��N��A���7���Ύ��d����������\��R����7��ę�
O���؜��a��N韼p�� ���Y{���������w������`��􏭼A��r������֘��?������� ������*'��:����/���  �  ?gN=K�M=��L=$L=�XK=�J=��I=�I=PBH={G=�F=l�E=� E=�VD=A�C=�B=��A=�#A=*T@=��?=�>=��==�
==5<=�];=l�:=R�9=��8=B�7=,7=I26=�O5=�j4=+�3=s�2=��1=��0=$�/=s�.=W�-=��,=��+=�+=2*=�)=��'=��&=x�%=I�$=��#=g�"=��!=i� =�m=�L=:(= =N�=֤=�q=�:=��=N�=�~={8=8�= �=�M=��=ĝ=�?
=��='x=z=�=�/=t�=�A =���<x��<ԁ�< s�<{]�<A�<��<[��<r��<]��<JR�<[�<���<�{�<|)�< ��<�u�<��<���<�E�<ؼ<ef�<�<Dx�<I��<4}�<S��<�v�<��<�f�<�ۙ<�N�<R��<z0�<}��<��<�z�<��<D�z<�s<�Yl<j3e<�^<��V<��O<w�H<�A<�o:<�X3<�E,<:7%<G-<m(<)<�/	<�<<���;��;��;�o�;տ;�K�;դ;q�;!�;!�y;�~_;�^E;�k+;	�;+)�:�d�:��:� 2:�9���E#鹬U��R����ɺ����Ny�
q*�W+A��W�K�m���fӌ�O����5��������[��T~˻�ջnf߻�+黺��[�������p ����X$������A"���&���*��.��3��7�x;��?��C���F��J��N��VR��V���Y�*l]��a��d��1h���k��7o���r�W v�7�y���|�C%���Ё�Zy��,��X�c��I��I���7���Ύ��d����������N��T����7��ę�O���؜��a��H韼p�����X{����������������j��쏭�;��{������ޘ��>������� ������''��.����/���  �  EgN=F�M=��L=%L=�XK=�J=��I=�I=LBH={G=#�F=l�E=� E=�VD=D�C= �B=��A=�#A=-T@=��?=�>=��==�
==5<=�];=q�:=U�9=��8=H�7=)7=J26=�O5=�j4=,�3=r�2=��1=}�0=(�/=q�.=U�-=��,=��+=�+=-*=�)=��'=��&=x�%=J�$=��#=c�"=��!=g� =�m=�L=:(= =G�=֤=�q=�:=��=R�=�~=y8=:�=��=�M=��=Ɲ=�?
=��=&x=w=��=�/=w�=�A =��<��<́�<$s�<t]�<A�<��<[��<}��<V��<RR�<S�<���<�{�<})�<%��<�u�<��<y��<�E�<ؼ<]f�<�<Ix�<R��<*}�<]��<�v�<��<�f�<�ۙ<�N�<F��<�0�<|��<��<�z�<��<R�z<�s<�Yl<`3e<�^<��V<n�O<x�H<�A<�o:<�X3<�E,<@7%<:-<u(<)<�/	<�<<���;<��;��;�o�;�Կ; L�;�Ԥ;q�;� �;U�y;�~_;p^E;5l+;§;�)�:|d�:=�:q!2:c�9�����$�aU��S����ɺ����^y��p*�~+A�ϧW�m�m���xӌ�G���b5��@�������[��L~˻�ջff߻�+�����Z�������� ����S$�0�����A"���&�Ƽ*��.��3��7�n;��?��C���F���J��N��VR��V���Y�l]��a�ۢd��1h���k��7o���r�Q v�C�y�y�|�D%���Ё�Oy��3��P�c��D��I���7���Ύ��d������͊��H��Z����7��ę�O���؜��a��>韼p�����\{�����������������k��폭�F��{������㘳�,������� ������3'��-����/���  �  ?gN=H�M=��L='L=�XK=�J=��I=�I=QBH={G=#�F=n�E=� E=�VD=<�C=�B=��A=�#A=*T@=��?=�>=��==�
==5<=�];=q�:=T�9=��8=C�7=+7=I26=�O5=�j4=0�3=o�2=��1=��0=%�/=w�.=T�-=��,=��+=�+=/*=�)=��'=��&=z�%=J�$=��#=i�"=��!=j� =�m=�L=9(= =K�=ؤ=�q=�:=��=T�=�~={8=6�=�=�M=��=ĝ=�?
=��=%x=}=�=�/=q�=�A =���<���<ׁ�<s�<v]�<A�<��<]��<z��<^��<HR�<Z�<���<�{�<})�<��<�u�<��<���<�E�<	ؼ<cf�<�<Lx�<B��<7}�<V��<�v�<��<�f�<�ۙ<�N�<J��<y0�<~��<��<�z�<��<N�z<�s<�Yl<X3e<�^<��V<y�O<x�H<�A<�o:<�X3<�E,<G7%<I-<r(<)<�/	<�<<���;@��;�;�o�;տ;�K�;�Ԥ;2q�;%!�;�y;�~_;�^E;)l+;��;)�:�d�:4�:U!2:h�9͖��$鹙U��R����ɺ����y�:q*�W+A���W��m��dӌ�L����5��/�����i[��]~˻��ջbf߻�+黬��[�����߈�z ����_$� ����|A"���&���*��.��3��7�};��?��C���F��J���N��VR��V���Y�"l]��a���d��1h���k��7o���r�\ v�?�y���|�C%���Ё�Ry��+��Z�	c��D��E���7���Ύ��d��������U��S����7��ę�O���؜��a��E韼p�����W{�����������������i��ꏭ�D��s������☳�>����� ������.'��-����/���  �  <gN=O�M=��L=$L=�XK=�J=��I=�I=SBH={G=%�F=k�E=� E=�VD=<�C=�B=��A=�#A=+T@=��?=�>=��==�
==
5<=�];=j�:=V�9=��8=>�7=.7=F26=�O5=�j4=.�3=t�2=��1=��0= �/=v�.=T�-=��,=��+=�+=7*=�)=��'=��&={�%=J�$=��#=k�"=��!=l� =�m=�L=;(= =O�=Ф=�q=�:=��=M�=�~=8=0�=�=�M=��=ĝ=�?
=��=$x=}=�=�/=s�=�A =���<r��<؁�<s�<]�<�@�<��<b��<l��<]��<@R�<g�<���<�{�<�)�<��<�u�<��<���<�E�<ؼ<af�<�<Ox�<C��<<}�<I��<�v�<��<�f�<�ۙ<�N�<Z��<u0�<}��<��<�z�<��<B�z<�s<�Yl<x3e<�^<��V<��O<q�H<�A<�o:<�X3<�E,<87%<@-<l(<()<�/	<�<<���;M��;��;�o�;'տ;�K�;*դ;�p�;!�;7�y;_;�^E;�k+;g�;�(�:�d�:j�:�!2:��95���G"�nU��R��D�ɺF���9y�%q*��*A�M�W��m��Pӌ�^����5��񶬻0��r[���~˻�ջ`f߻,默��[��������q ����Y$���)��qA"���&���*�!�.��3��7��;��?��C���F��J��N��VR��V���Y�:l]��a��d��1h���k��7o���r�e v�/�y���|�@%���Ё�_y��,��b��b��M��K���7���Ύ��d����������V��M����7��!ę�O���؜��a��R韼p�����]{����������y������j��鏭�A��y������՘��>������� ������*'��1����/���  �  CgN=G�M=��L=&L=�XK=�J=��I=�I=QBH={G=#�F=p�E=� E=�VD=<�C=�B=��A=�#A=*T@=��?=�>=��==�
==5<=�];=o�:=V�9=��8=E�7=,7=F26=�O5=�j4=.�3=r�2=��1=��0=(�/=u�.=T�-=��,=��+=�+=0*=�)=��'=��&=x�%=J�$=��#=g�"=��!=l� =�m=�L=8(= =M�=֤=�q=�:=��=Q�=�~=z8=6�=�=�M=��=Ɲ=�?
=��=%x=z=��=�/=r�=�A =��<��<ԁ�<s�<y]�<A�<��<a��<w��<b��<KR�<W�<���<�{�<�)�<��<�u�<��<���<�E�<ؼ<df�<�<Mx�<I��<5}�<R��<�v�<��<�f�<�ۙ<�N�<K��<�0�<}��<��<�z�<��<Y�z<�s<�Yl<b3e<�^<��V<z�O<i�H<�A<�o:<�X3<�E,<@7%<P-<n(<)<�/	<�<<���;>��;�;�o�;�Կ;�K�;�Ԥ;q�;/!�;"�y;�~_;�^E;�k+;�;V)�:Ee�:��:�!2:��99����#�cU��R����ɺ@���ay�q*�V+A�ȧW�,�m��hӌ�<���m5��"�����v[��X~˻�ջgf߻�+黷��[�����ވ�q ����b$�����rA"���&���*��.��3��7�;��?��C���F���J��N��VR��V���Y�l]��a��d��1h���k��7o���r�` v�:�y��|�C%���Ё�Uy��'��W�c��K��F���7���Ύ��d��������X��Z����7��ę�O���؜��a��I韼p�����S{�����������������j������D��v������☳�>������� ������-'��5����/���  �  FgN=G�M=��L="L=�XK= �J=��I=�I=OBH={G= �F=m�E=� E=�VD=E�C=�B=��A=�#A=*T@=��?=�>=��==�
==5<=�];=m�:=U�9=��8=I�7=%7=N26=�O5=�j4=+�3=o�2=��1=z�0=&�/=p�.=Y�-=��,=��+=�+=-*=�)=��'=��&=v�%=J�$=��#=f�"=��!=g� =�m=�L=<(= =I�=ؤ=�q=�:=��=S�=�~=x8=:�=��=�M=��=Ɲ=�?
=��=*x=v=�=�/=v�=�A =��<{��<ρ�<)s�<m]�<A�<��<^��<x��<V��<QR�<S�<���<�{�<z)�<��<�u�<��<��<�E�<	ؼ<^f�<�<Cx�<J��<1}�<]��<�v�<��<�f�<�ۙ<�N�<F��<�0�<v��<��<�z�<��<J�z<�s<�Yl<O3e<�^<��V<~�O<��H<��A<�o:<�X3<�E,<07%<K-<x(<	)<�/	<�<<���;"��; �;�o�; տ;L�;�Ԥ;'q�;!�;#�y;�~_;�^E;8l+;ͧ;�)�:�d�:��:�!2:��9Ћ��'�fU�;S���ɺ�����y��p*��+A��W�y�m���vӌ�O���m5��<�������[��C~˻�ջcf߻�+�����Z�����܈�� ����N$�(��	���A"���&���*�
�.��3��7�n;��?��C���F���J���N��VR��V���Y�!l]��a�ߢd��1h���k��7o���r�E v�R�y�{�|�C%���Ё�Sy��3��Q�c��A��F���7���Ύ��d������Ɗ��F��S����7��ę�O���؜��a��>韼p�����S{������򃧼�������q��菭�>��~������옳�-��Ɲ��� ������+'��)����/���  �  @gN=K�M=��L=%L=�XK=�J=��I=�I=QBH={G=&�F=l�E=� E=�VD==�C=�B=��A=�#A=/T@=��?=�>=��==�
==
5<=�];=n�:=T�9=��8=C�7=*7=I26=�O5=�j4=0�3=q�2=��1=��0=&�/=s�.=U�-=��,=��+=�+=1*=�)=��'=��&=x�%=J�$=��#=i�"=��!=j� =�m=�L=;(= =K�=Ԥ=�q=�:=��=O�=�~={8=4�= �=�M=��=Ý=�?
=��=&x=y=�=�/=t�=�A =���<z��<Ё�<s�<v]�<A�<��<]��<x��<[��<BR�<]�<���<�{�<~)�<$��<�u�<��<���<�E�<ؼ<Zf�<�<Nx�<H��<8}�<Q��<�v�<��<�f�<�ۙ<�N�<O��<{0�<}��<��<�z�<��<P�z<�s<�Yl<f3e<�^<��V<n�O<u�H<�A<�o:<�X3<�E,<?7%<B-<`(<)<�/	<�<<���;Q��;��;�o�;տ;�K�;դ;	q�;!�;n�y;�~_;�^E;�k+;#�;�(�:�d�:��:O!2:��9�����$鹛U�bS���ɺ	���ky��p*�:+A��W�P�m���nӌ�U���5�������z[��l~˻
�ջdf߻�+黪�� [�������| ����Y$�����~A"���&���*��.��3��7��;��?��C���F��J��N��VR��V���Y�#l]��a��d��1h���k��7o���r�\ v�?�y���|�D%���Ё�Ty��.��`�c��J��G���7���Ύ��d����������S��P����7��ę�O���؜��a��J韼p�����[{�����������������j��폭�F��{������ޘ��5������� ������3'��/����/���  �  <gN=L�M=��L='L=�XK=�J=��I=�I=VBH={G=%�F=o�E=� E=�VD=<�C=�B=��A=�#A=+T@=��?=��>=��==�
==	5<= ^;=m�:=P�9=��8=A�7=27=C26=�O5=�j4=-�3=r�2=��1=��0=#�/=x�.=Q�-=��,=��+=�+=2*=�)=��'=��&=}�%=M�$=��#=k�"=��!=o� =�m=�L=:(= =P�=դ=�q=�:=��=R�=�~=�8=3�=�=�M=��=Ý=�?
=��= x==�=�/=p�=�A =��<z��<܁�<s�<�]�<A�<��<W��<q��<h��<AR�<h�<���<�{�<|)�<��<�u�<��<���<�E�<ؼ<cf�<�<Qx�<<��<?}�<M��<�v�<��<�f�<�ۙ<�N�<S��<t0�<���<��<�z�<��<F�z<�s<�Yl<g3e<�^<��V<z�O<h�H<&�A<�o:<�X3<�E,<E7%<O-<e(<-)<�/	<�<<q��;L��;�;�o�;0տ;�K�; դ;q�;7!�;1�y;�~_;�^E;�k+;u�;�(�:�e�:��:b 2:��9>���* ��U��R����ɺt���\y�Lq*�H+A�#�W���m�!�Uӌ�=����5�����:��N[��m~˻܁ջMf߻�+黗��/[�������k ����\$�����fA"���&���*��.��3��7��;��?��C���F��J���N��VR�V���Y�0l]��a���d��1h���k��7o���r�u v�!�y���|�C%���Ё�Zy�� ��a��b��O��>���7���Ύ��d����������V��K����7��ę�O���؜��a��N韼p�����W{����������������`������F��r������ݘ��F������� ������-'��5����/���  �  AgN=N�M=��L=&L=�XK=�J=��I=�I=TBH={G=#�F=k�E=� E=�VD=A�C=�B=��A=�#A=,T@=��?=�>=��==�
==5<=�];=m�:=V�9=��8=D�7=,7=E26=�O5=�j4=-�3=t�2=��1=��0=#�/=u�.=R�-=��,=��+=�+=4*=�)=��'=��&=y�%=H�$=��#=j�"=��!=i� =�m=�L=;(= =K�=Ԥ=�q=�:=��=S�=�~={8=3�= �=�M=��=Ɲ=�?
=��=!x=|=�=�/=v�=�A =��<w��<ց�<s�<{]�<A�<��<a��<w��<[��<DR�<]�<���<�{�<�)�<��<�u�<��<���<�E�<ؼ<af�<�<Ix�<I��<;}�<Q��<�v�<��<�f�<�ۙ<�N�<V��<}0�<|��<��<�z�<��<F�z<
�s<�Yl<f3e<�^<��V<x�O<l�H<�A<�o:<�X3<�E,<@7%<?-<l(<)<�/	<�<<���;>��;��;�o�;տ;�K�;�Ԥ;q�;	!�;>�y;_;�^E;�k+;�;�(�:�d�:��:�!2:R�9<����#鹀U��R����ɺc���<y��p*�P+A��W�$�m��`ӌ�R���r5�������x[��z~˻��ջsf߻�+黠���Z�������{ ����W$�!�����A"���&���*��.��3��7��;��?��C���F���J���N��VR�V���Y�.l]��a�ߢd��1h���k��7o���r�i v�5�y���|�=%���Ё�Uy��.��^�c��N��A���7���Ύ��d������Ċ��N��T����7�� ę�O���؜��a��J韼p�����^{����������}������k��폭�E��w������ߘ��2������� ������.'��3����/���  �  BgN=D�M=��L='L=�XK=!�J=��I=�I=LBH={G="�F=l�E=� E=�VD=A�C=�B=��A=�#A=-T@=��?=�>=��==�
==5<=�];=o�:=S�9=��8=E�7=)7=K26=�O5=�j4=1�3=l�2=��1=~�0='�/=s�.=T�-=��,=��+=�+=,*=�)=��'=��&=|�%=G�$=��#=d�"=��!=e� =�m=�L=;(= =L�=ۤ=�q=�:=��=O�=�~=}8=8�=��=�M=��=ĝ=�?
=��=$x=x=��=�/=p�=�A =���<{��<́�<!s�<x]�<A�<��<W��<z��<W��<PR�<Z�<���<�{�<�)�<%��<�u�<��<~��<�E�<ؼ<kf�<�<Fx�<O��<,}�<T��<�v�<��<�f�<�ۙ<�N�<C��<�0�<y��<��<�z�<��<X�z<�s<�Yl<J3e<�^<��V<l�O<|�H<�A<�o:<�X3<�E,<E7%<F-<~(<)<�/	<�<<���;6��;��;�o�;�Կ;�K�;�Ԥ;Rq�;� �;Y�y;!_;G^E;�k+; �;�)�:�d�:��:!2:�9s����$�U��S��ݩɺ�����y�"q*�p+A�קW�L�m��Rӌ�I���r5��G������[��N~˻�ջwf߻�+�����Z�����Ԉ�o ����X$�������A"���&�ü*��.��3��7�u;��?��C���F��J���N��VR��V���Y�l]��a���d��1h���k��7o���r�U v�<�y���|�J%���Ё�Qy��1��Q�	c��J��O���7���Ύ��d������Ǌ��N��Y����7��ę�O���؜��a��G韼 p�����X{�����������������n��班�G��z������똳�:��ɝ�� ������4'��+����/���  �  AgN=N�M=��L=&L=�XK=�J=��I=�I=TBH={G=#�F=k�E=� E=�VD=A�C=�B=��A=�#A=,T@=��?=�>=��==�
==5<=�];=m�:=V�9=��8=D�7=,7=E26=�O5=�j4=-�3=t�2=��1=��0=#�/=u�.=R�-=��,=��+=�+=4*=�)=��'=��&=y�%=H�$=��#=j�"=��!=i� =�m=�L=;(= =K�=Ԥ=�q=�:=��=S�=�~={8=3�= �=�M=��=Ɲ=�?
=��=!x=|=�=�/=v�=�A =��<w��<ց�<s�<{]�<A�<��<a��<w��<[��<DR�<]�<���<�{�<�)�<��<�u�<��<���<�E�<ؼ<af�<�<Ix�<I��<;}�<Q��<�v�<��<�f�<�ۙ<�N�<V��<}0�<|��<��<�z�<��<F�z<
�s<�Yl<f3e<�^<��V<x�O<l�H<�A<�o:<�X3<�E,<@7%<?-<l(<)<�/	<�<<���;>��;��;�o�;տ;�K�;�Ԥ;q�;	!�;>�y;_;�^E;�k+;�;�(�:�d�:��:�!2:Q�9?����#鹁U��R����ɺc���<y��p*�P+A��W�$�m��`ӌ�R���r5�������x[��z~˻��ջsf߻�+黠���Z�������{ ����W$�!�����A"���&���*��.��3��7��;��?��C���F���J���N��VR�V���Y�.l]��a�ߢd��1h���k��7o���r�h v�5�y���|�=%���Ё�Uy��.��^�c��N��A���7���Ύ��d������Ċ��N��T����7�� ę�O���؜��a��J韼p�����^{����������}������k��폭�E��w������ߘ��2������� ������.'��3����/���  �  <gN=L�M=��L='L=�XK=�J=��I=�I=VBH={G=%�F=o�E=� E=�VD=<�C=�B=��A=�#A=+T@=��?=��>=��==�
==	5<= ^;=m�:=P�9=��8=A�7=27=C26=�O5=�j4=-�3=r�2=��1=��0=#�/=x�.=Q�-=��,=��+=�+=2*=�)=��'=��&=}�%=M�$=��#=k�"=��!=o� =�m=�L=:(= =P�=դ=�q=�:=��=R�=�~=�8=3�=�=�M=��=Ý=�?
=��= x==�=�/=p�=�A =��<z��<܁�<s�<�]�<A�<��<W��<q��<h��<AR�<h�<���<�{�<|)�<��<�u�<��<���<�E�<ؼ<cf�<�<Qx�<<��<?}�<M��<�v�<��<�f�<�ۙ<�N�<S��<t0�<���<��<�z�<��<F�z<�s<�Yl<g3e<�^<��V<z�O<h�H<&�A<�o:<�X3<�E,<E7%<O-<e(<-)<�/	<�<<q��;L��;�;�o�;0տ;�K�; դ;q�;7!�;1�y;�~_;�^E;�k+;u�;�(�:�e�:��:a 2:��9B���+ ��U��R����ɺt���\y�Mq*�H+A�#�W���m�!�Uӌ�=����5�����:��N[��m~˻݁ջMf߻�+黗��/[�������k ����\$�����fA"���&���*��.��3��7��;��?��C���F��J���N��VR�V���Y�0l]��a���d��1h���k��7o���r�u v�!�y���|�C%���Ё�Zy�� ��a��b��O��>���7���Ύ��d����������V��K����7��ę�O���؜��a��N韼p�����W{����������������`������F��r������ݘ��F������� ������-'��5����/���  �  @gN=K�M=��L=%L=�XK=�J=��I=�I=QBH={G=&�F=l�E=� E=�VD==�C=�B=��A=�#A=/T@=��?=�>=��==�
==
5<=�];=n�:=T�9=��8=C�7=*7=I26=�O5=�j4=0�3=q�2=��1=��0=&�/=s�.=U�-=��,=��+=�+=1*=�)=��'=��&=x�%=J�$=��#=i�"=��!=j� =�m=�L=;(= =K�=Ԥ=�q=�:=��=O�=�~={8=4�= �=�M=��=Ý=�?
=��=&x=y=�=�/=t�=�A =���<z��<Ё�<s�<v]�<A�<��<]��<x��<[��<CR�<]�<���<�{�<~)�<$��<�u�<��<���<�E�<ؼ<Zf�<�<Nx�<H��<8}�<Q��<�v�<��<�f�<�ۙ<�N�<O��<{0�<}��<��<�z�<��<P�z<�s<�Yl<f3e<�^<��V<n�O<u�H<�A<�o:<�X3<�E,<?7%<B-<`(<)<�/	<�<<���;Q��;��;�o�;տ;�K�;դ;	q�;!�;m�y;�~_;�^E;�k+;#�;�(�:�d�:��:N!2:��9�����$鹜U�cS���ɺ
���ky��p*�:+A��W�P�m���nӌ�V���5�������z[��l~˻
�ջdf߻�+黪�� [�������| ����Y$�����~A"���&���*��.��3��7��;��?��C���F��J��N��VR��V���Y�#l]��a��d��1h���k��7o���r�\ v�?�y���|�D%���Ё�Ty��.��`�c��J��G���7���Ύ��d����������S��P����7��ę�O���؜��a��J韼p�����[{�����������������j��폭�F��{������ޘ��5������� ������3'��/����/���  �  FgN=G�M=��L="L=�XK= �J=��I=�I=OBH={G= �F=m�E=� E=�VD=E�C=�B=��A=�#A=*T@=��?=�>=��==�
==5<=�];=m�:=U�9=��8=I�7=%7=N26=�O5=�j4=+�3=o�2=��1=z�0=&�/=p�.=Y�-=��,=��+=�+=-*=�)=��'=��&=v�%=J�$=��#=f�"=��!=g� =�m=�L=<(= =I�=ؤ=�q=�:=��=S�=�~=x8=:�=��=�M=��=Ɲ=�?
=��=*x=v=�=�/=v�=�A =��<{��<ρ�<)s�<m]�<A�<��<^��<x��<V��<QR�<S�<���<�{�<z)�<��<�u�<��<��<�E�<	ؼ<^f�<�<Cx�<J��<1}�<]��<�v�<��<�f�<�ۙ<�N�<F��<�0�<v��<��<�z�<��<J�z<�s<�Yl<O3e<�^<��V<~�O<��H<��A<�o:<�X3<�E,<07%<K-<x(<	)<�/	<�<<���;"��; �;�o�; տ;L�;�Ԥ;'q�;!�;#�y;�~_;�^E;8l+;ͧ;�)�:�d�:��:�!2:��9ً��'�gU�<S���ɺ�����y��p*��+A��W�y�m���vӌ�O���m5��<�������[��C~˻�ջcf߻�+�����Z�����܈�� ����N$�(��	���A"���&���*�
�.��3��7�n;��?��C���F���J���N��VR��V���Y�!l]��a�ߢd��1h���k��7o���r�E v�R�y�{�|�C%���Ё�Sy��3��Q�c��A��F���7���Ύ��d������Ɗ��F��S����7��ę�O���؜��a��>韼p�����S{������򃧼�������q��菭�>��~������옳�-��Ɲ��� ������+'��)����/���  �  CgN=G�M=��L=&L=�XK=�J=��I=�I=QBH={G=#�F=p�E=� E=�VD=<�C=�B=��A=�#A=*T@=��?=�>=��==�
==5<=�];=o�:=V�9=��8=E�7=,7=F26=�O5=�j4=.�3=r�2=��1=��0=(�/=u�.=T�-=��,=��+=�+=0*=�)=��'=��&=x�%=J�$=��#=g�"=��!=l� =�m=�L=8(= =M�=֤=�q=�:=��=Q�=�~=z8=6�=�=�M=��=Ɲ=�?
=��=%x=z=��=�/=r�=�A =��<��<ԁ�<s�<y]�<A�<��<a��<w��<b��<KR�<X�<���<�{�<�)�<��<�u�<��<���<�E�<ؼ<df�<�<Mx�<I��<5}�<R��<�v�<��<�f�<�ۙ<�N�<K��<�0�<}��<��<�z�<��<Y�z<�s<�Yl<b3e<�^<��V<z�O<i�H<�A<�o:<�X3<�E,<@7%<P-<n(<)<�/	<�<<���;>��;�;�o�;�Կ;�K�;�Ԥ;q�;/!�;"�y;�~_;�^E;�k+;�;V)�:Ee�:��:�!2:��9A����#�dU��R����ɺA���by�q*�V+A�ȧW�,�m��hӌ�<���n5��"�����v[��X~˻�ջgf߻�+黸��[�����ވ�q ����b$�����rA"���&���*��.��3��7�;��?��C���F���J��N��VR��V���Y�l]��a��d��1h���k��7o���r�` v�:�y��|�C%���Ё�Uy��'��W�c��K��F���7���Ύ��d��������X��Z����7��ę�O���؜��a��I韼p�����S{�����������������j������D��v������☳�>������� ������-'��5����/���  �  <gN=O�M=��L=$L=�XK=�J=��I=�I=SBH={G=%�F=k�E=� E=�VD=<�C=�B=��A=�#A=+T@=��?=�>=��==�
==
5<=�];=j�:=V�9=��8=>�7=.7=F26=�O5=�j4=.�3=t�2=��1=��0= �/=v�.=T�-=��,=��+=�+=7*=�)=��'=��&={�%=J�$=��#=k�"=��!=l� =�m=�L=;(= =O�=Ф=�q=�:=��=M�=�~=8=0�=�=�M=��=ĝ=�?
=��=$x=}=�=�/=s�=�A =���<r��<؁�<s�<]�<�@�<��<b��<l��<]��<@R�<g�<���<�{�<�)�<��<�u�<��<���<�E�<ؼ<af�<�<Ox�<C��<<}�<I��<�v�<��<�f�<�ۙ<�N�<Z��<u0�<}��<��<�z�<��<B�z<�s<�Yl<x3e<�^<��V<��O<q�H<�A<�o:<�X3<�E,<87%<@-<l(<()<�/	<�<<���;M��;��;�o�;'տ;�K�;*դ;�p�;!�;7�y;_;�^E;�k+;g�;�(�:�d�:i�:�!2:��9>���J"�oU��R��E�ɺF���9y�%q*��*A�M�W��m��Pӌ�^����5��񶬻0��r[���~˻�ջ`f߻,默��[��������q ����Y$���)��qA"���&���*�!�.��3��7��;��?��C���F��J��N��VR��V���Y�:l]��a��d��1h���k��7o���r�e v�/�y���|�@%���Ё�_y��,��b��b��M��K���7���Ύ��d����������V��M����7��!ę�O���؜��a��R韼p�����]{����������y������j��鏭�A��y������՘��>������� ������*'��1����/���  �  ?gN=H�M=��L='L=�XK=�J=��I=�I=QBH={G=#�F=n�E=� E=�VD=<�C=�B=��A=�#A=*T@=��?=�>=��==�
==5<=�];=q�:=T�9=��8=C�7=+7=I26=�O5=�j4=0�3=o�2=��1=��0=%�/=w�.=T�-=��,=��+=�+=/*=�)=��'=��&=z�%=J�$=��#=i�"=��!=j� =�m=�L=9(= =K�=ؤ=�q=�:=��=T�=�~={8=6�=�=�M=��=ĝ=�?
=��=%x=}=�=�/=q�=�A =���<���<ׁ�<s�<v]�<A�<��<]��<z��<^��<HR�<Z�<���<�{�<})�<��<�u�<��<���<�E�<	ؼ<cf�<�<Lx�<B��<7}�<V��<�v�<��<�f�<�ۙ<�N�<J��<y0�<~��<��<�z�<��<N�z<�s<�Yl<X3e<�^<��V<y�O<x�H<�A<�o:<�X3<�E,<G7%<I-<r(<)<�/	<�<<���;@��;�;�o�;տ;�K�;�Ԥ;2q�;%!�;�y;�~_;�^E;(l+;��;)�:�d�:3�:T!2:e�9ז�� $鹛U��R����ɺ����y�:q*�W+A���W��m��dӌ�L����5��/�����i[��]~˻��ջbf߻�+黬��[�����߈�z ����_$� ����|A"���&���*��.��3��7�};��?��C���F��J���N��VR��V���Y�"l]��a���d��1h���k��7o���r�\ v�?�y���|�C%���Ё�Ry��+��Z�	c��D��E���7���Ύ��d��������U��S����7��ę�O���؜��a��E韼p�����W{�����������������i��ꏭ�D��s������☳�>����� ������.'��-����/���  �  EgN=F�M=��L=%L=�XK=�J=��I=�I=LBH={G=#�F=l�E=� E=�VD=D�C= �B=��A=�#A=-T@=��?=�>=��==�
==5<=�];=q�:=U�9=��8=H�7=)7=J26=�O5=�j4=,�3=r�2=��1=}�0=(�/=q�.=U�-=��,=��+=�+=-*=�)=��'=��&=x�%=J�$=��#=c�"=��!=g� =�m=�L=:(= =G�=֤=�q=�:=��=R�=�~=y8=:�=��=�M=��=Ɲ=�?
=��=&x=w=��=�/=w�=�A =��<��<́�<$s�<t]�<A�<��<[��<}��<V��<SR�<S�<���<�{�<})�<%��<�u�<��<y��<�E�<ؼ<]f�<�<Ix�<R��<*}�<]��<�v�<��<�f�<�ۙ<�N�<F��<�0�<|��<��<�z�<��<R�z<�s<�Yl<`3e<�^<��V<n�O<x�H<�A<�o:<�X3<�E,<@7%<:-<u(<)<�/	<�<<���;<��;��;�o�;�Կ; L�;�Ԥ;q�;� �;U�y;�~_;o^E;5l+;§;�)�:|d�:<�:p!2:b�9�����$�bU��S����ɺ����_y��p*�~+A�ϧW�m�m���xӌ�G���b5��@�������[��L~˻�ջff߻�+�����Z�������� ����S$�0�����A"���&�Ƽ*��.��3��7�n;��?��C���F���J��N��VR��V���Y�l]��a�ۢd��1h���k��7o���r�Q v�C�y�y�|�D%���Ё�Oy��3��P�c��D��I���7���Ύ��d������͊��H��Z����7��ę�O���؜��a��>韼p�����\{�����������������k��폭�F��{������㘳�,������� ������3'��-����/���  �  ?gN=K�M=��L=$L=�XK=�J=��I=�I=PBH={G=�F=l�E=� E=�VD=A�C=�B=��A=�#A=*T@=��?=�>=��==�
==5<=�];=l�:=R�9=��8=B�7=,7=I26=�O5=�j4=+�3=s�2=��1=��0=$�/=s�.=W�-=��,=��+=�+=2*=�)=��'=��&=x�%=I�$=��#=g�"=��!=i� =�m=�L=:(= =N�=֤=�q=�:=��=N�=�~={8=8�= �=�M=��=ĝ=�?
=��='x=z=�=�/=t�=�A =���<x��<ԁ�< s�<{]�<A�<��<[��<r��<]��<JR�<[�<���<�{�<|)�< ��<�u�<��<���<�E�<ؼ<ef�<�<Dx�<I��<4}�<S��<�v�<��<�f�<�ۙ<�N�<R��<z0�<}��<��<�z�<��<D�z<�s<�Yl<j3e<�^<��V<��O<w�H<�A<�o:<�X3<�E,<:7%<G-<m(<)<�/	<�<<���;��;��;�o�;տ;�K�;դ;q�;!�;!�y;�~_;�^E;�k+;	�;*)�:�d�:��:� 2:
�9����G#鹬U��R����ɺ����Ny�
q*�X+A��W�K�m���fӌ�O����5��������[��T~˻�ջnf߻�+黺��[�������p ����X$������A"���&���*��.��3��7�x;��?��C���F��J��N��VR��V���Y�*l]��a��d��1h���k��7o���r�W v�7�y���|�C%���Ё�Zy��,��X�c��I��I���7���Ύ��d����������N��T����7��ę�O���؜��a��H韼p�����X{����������������j��쏭�;��{������ޘ��>������� ������''��.����/���  �  <gN=P�M=��L=(L=�XK=�J=��I=�I=XBH={G=$�F=o�E=� E=�VD=8�C=�B=��A=�#A=(T@=��?=��>=��==�
==5<=�];=m�:=V�9=��8=A�7=/7=C26=�O5=�j4=/�3=u�2=��1=��0=%�/=z�.=R�-=��,=��+=�+=7*=�)=��'=��&=v�%=I�$=��#=n�"=��!=n� =�m=�L=9(= =L�=Ӥ=�q=�:=��=P�=�~=z8=2�=�=�M=��=ŝ=�?
=��="x=�=�=�/=r�=�A =���<{��<݁�<s�<]�<A�<��<f��<s��<i��<=R�<^�<���<�{�<�)�<��<�u�<��<���<�E�<
ؼ<^f�<�<Qx�<?��<E}�<M��<�v�<��<�f�<�ۙ<�N�<[��<t0�<���<��<�z�<��<G�z<�s<�Yl<y3e<�^<��V<�O<`�H< �A<�o:<�X3<�E,<K7%<I-<U(<)<�/	<�<<���;D��;�;�o�;տ;�K�;դ;q�;7!�;�y;�~_;�^E;�k+;%�;I(�:�e�:��:�!2:��9ܚ���!�+U��R��ǩɺ���3y�,q*�+A���W���m��jӌ�,����5��񶬻)��N[��w~˻�ջmf߻�+黀��?[�������x ����a$�����kA"���&���*��.��3��7��;��?��C���F��J��N��VR�V���Y�'l]��a��d��1h���k��7o���r�p v�.�y���|�;%���Ё�Yy��!��e�c��N��A���7���Ύ��d����������\��R����7��ę�
O���؜��a��N韼p�� ���Y{���������w������`��􏭼A��r������֘��?������� ������*'��:����/���  �  >gN=J�M=��L=$L=�XK=�J=��I=�I=QBH={G=#�F=m�E=� E=�VD=B�C=�B=��A=�#A=)T@=��?=�>=��==�
==5<=�];=k�:=V�9=��8=D�7=-7=I26=�O5=�j4=.�3=q�2=��1=~�0=%�/=r�.=U�-=��,=��+=�+=1*=�)=��'=��&={�%=M�$=��#=j�"=��!=l� =�m=�L==(= =K�=Ӥ=�q=�:=��=P�=�~=~8=7�= �=�M=��==�?
=��=&x=y=�=�/=t�=�A =��<x��<ҁ�<!s�<|]�<
A�<��<`��<o��<_��<JR�<b�<���<�{�<)�<��<�u�<��<���<�E�<ؼ<`f�<�<Lx�<B��<7}�<U��<�v�<��<�f�<�ۙ<�N�<P��<w0�<���<��<�z�<��<J�z<�s<�Yl<c3e<�^<��V<{�O<w�H<�A<�o:<�X3<�E,<87%<F-<p(<()<�/	<�<<���;;��;�;�o�;տ;�K�;�Ԥ;q�;!�;�y;�~_;�^E;�k+;F�; )�:e�:q�:�!2:��9�����"鹆U�4S��)�ɺW���iy��p*�p+A��W�[�m��Yӌ�6����5����� ���[��\~˻�ջOf߻�+黡��&[�������{ ����P$�����uA"���&���*��.��3��7�|;��?��C���F��J��N��VR��V���Y�(l]��a��d��1h���k��7o���r�V v�5�y���|�E%���Ё�\y��+��X�c��G��H���7���Ύ��d����������K��O����7��ę�O���؜��a��G韼p�����Z{�����������������d��鏭�@��|������☳�3������� ������-'��.����/���  �  �hN=+�M=�L=�L=�[K='�J=�I=zI=2FH=PG=��F=C�E=&E=�[D=�C=(�B=R�A=d*A=^[@=A�?=�>=W�==i===><=�g;=k�:=��9=x�8=��7=�7=y>6=*\5=�w4=Ñ3=��2=�1=��0=��/=y�.=��-=�-=,=�+=�*=�)=)(=�'=�&=-�$=M�#=/�"=һ!=� =�=;d=@=:=��=��=��=�S=d=��=��=kR=I=�=h=�=�=�Y
=��=�=	(=R�=�H=A�=Z =5��<
��<���<���<Y��<m�<�H�<3�<9��<��<�x�<v5�<���<]��<�J�<��<��<=2�<]��<V`�<�<~�<Q�<��<��<��<��<ȅ�<|��<�r�<H�<X�<Ȓ<�6�<P��<��<�|�<,�<��z<4|s<ARl<�(e<� ^<w�V<[�O<n�H<qA<HT:<9:3<�$,<�%<"<��<1�< 	<
<T6�;#f�;���;���;tT�;PƱ;�I�;�;���;�x;%@^;�D;*;RL;�a�:#��:��:#-,:8�9@�ʸ����Fs[�ё��'�̺����'��#,���B��`Y���o��т�#���4t��P��m��������:»�\̻<_ֻLB�$�6��B1���L����߇���ň����0Q� �"�O�&��+�A/��\3��l7�mp;��h?��UC��7G��K���N���R�|WV�,Z���]�MKa�W�d�5mh�!�k�Coo�B�r��Sv��y�<}�L<���恼�����3���Ն��u��=��~���}G���ގ��s�����?���(��p���HC���Ι�2Y��H✼vj�����w�����Ё�����G���V������������������!��陳����������������%�����-���  �  �hN=,�M=�L=�L=�[K="�J=�I=}I=7FH=OG=��F=?�E=&E=\D=�C=-�B=L�A=e*A=h[@=D�?=�>=Z�==q==6><=�g;=g�:=��9=s�8=��7=�7=w>6=,\5=�w4=��3=��2= �1=��0=��/=w�.=��-=�-=
,=�+=�*=�)=-(=�'=�&=5�$=Q�#=8�"=ջ!=� =�=9d=@=8=��=��=��=�S=l=��=��=oR=E=�=h=�=շ=�Y
=��=�=(=H�=�H=D�=Z =5��<��<���<���<\��<�l�<�H�<4�<.��<��<�x�<�5�<���<e��<�J�<$��<���</2�<c��<L`�<�<~�<E�<��<��<��<��<օ�<t��<�r�<P�<�W�<Ȓ<�6�<Q��<��<�|�<1�<k�z<=|s<IRl<�(e<p ^<�V<X�O<s�H<&qA<�S:<<:3<�$,<�%<"<t�<N�<$ 	<.
<L6�;_f�;t��;���;�T�;)Ʊ;�I�;���;���;��x;c@^;D;E*;�L;a�:@��:~�:d-,:�9�˸�����s[�����N�̺f����'�o#,���B�;aY��o��т����jt�����Q��������:»�\̻0_ֻB����/1���L��������͈���QQ��"�<�&�+�A/��\3��l7�p;��h?��UC��7G��K���N���R��WV�1Z���]�HKa�M�d�)mh� �k�Qoo�:�r� Tv��y��}�\<���恼�����3���Ն��u��6��u���pG��nގ��s�����9���(��d���PC���Ι�&Y��J✼ij��~񟼹w��$���Ё�����J���Q��ގ��������������3��噳����������������%�����-���  �  �hN=4�M=�L=�L=�[K=�J=�I=uI=8FH=FG=��F=?�E=&E=\D=�C=4�B=L�A=e*A=b[@==�?=�>=S�==s==/><=�g;=f�:=��9={�8=��7=�7=r>6=-\5=�w4=��3=��2=�1=��0=��/=|�.=��-=�-=,=�+=�*=�)=1(=�'=�&=3�$=J�#=8�"=˻!=� =�=?d=@=5=��=��=��=�S=j=��=��=oR=?=!�=�g=�=ط=�Y
=��=ޑ=(=F�=�H=A�=Z =7��<���<���<��<r��<�l�<�H�<9�<*��<���<�x�<�5�<���<b��<�J�<��<���</2�<s��<<`�<$�<
~�<F�<��<��< ��<��<؅�<k��<�r�<U�<�W�<Ȓ<�6�<g��<��<�|�<8�<\�z<N|s<9Rl<�(e<e ^<��V<N�O<k�H<UqA<�S:<_:3<s$,<�%<5<a�<U�< 	<3
<6�;Pf�;x��;���;�T�;�ű;(J�;���;���;<�x;�?^;
D;�*;�L;0`�:��:L�:[-,:��9T˸ϵ���t[�k���g�̺i����'��#,�Q�B�eaY�ġo��т�ݲ��$t�������������:»�\̻8_ֻ B�@���~1���L����͇���ۈ����OQ��"�a�&��+�A/��\3��l7��p;��h?��UC��7G��K���N�o�R��WV�Z���]�:Ka�Z�d�*mh��k�Yoo�-�r�Tv��y�v}�P<���恼�����3���Ն��u��B��w���|G��~ގ��s�����)���!(��^���JC���Ι�'Y��^✼gj���񟼷w��,���́�����V���>��㎪�������������;��ݙ�����������������%������,���  �  �hN=0�M=�L=�L=�[K=#�J=�I=vI==FH=NG=��F=D�E=&E=\D=�C=.�B=K�A=g*A=b[@=C�?=�>=S�==u==5><=�g;=i�:=��9=x�8=��7=�7=s>6=.\5=�w4=đ3=��2=�1=��0=��/=y�.=��-=�-=,=�+=�*=�)=.(=�'=�&=5�$=Q�#=<�"=һ!=� =�=:d=@=8=��=��=��=�S=o=�=��=sR=B=�= h=�=ٷ=�Y
=��=�=
(=J�=�H=?�=Z ==��< ��<���<��<[��<�l�<�H�<3�<0��<��<�x�<�5�<���<q��<�J�<��<���</2�<f��<K`�<�<~�<O�<��<��<)��<��<ۅ�<x��<�r�<Q�<�W�<Ȓ<�6�<R��<��<�|�<0�<r�z<O|s<-Rl<�(e<w ^<|�V<\�O<`�H<"qA<�S:<L:3<v$,<�%<,<{�<Y�< 	<G
<E6�;Cf�;���;���;�T�;Ʊ;�I�;���;ȋ�;8�x;W@^;vD;�*;M;�`�:���:��:-,:q�9˸Ļ���t[�K�����̺�����'��#,�i�B�aY��o��т�#���ft�����C��������:»�\̻_ֻB��˪�E1���L���������ψ����LQ��"�J�&�t+��@/��\3��l7��p;��h?��UC��7G��K���N���R��WV�'Z���]�<Ka�a�d�)mh��k�Woo�/�r�Tv��y�|}�T<���恼�����3���Ն��u��A��i���rG��zގ�}s�����6���(��f���PC���Ι�)Y��O✼_j���񟼴w�����Ё�����Q���H��܎��������������0��ܙ�����������������%�����-���  �  �hN=+�M= �L=�L=�[K=#�J=�I=zI=4FH=KG=��F=D�E=&E= \D=�C=,�B=P�A=g*A=e[@=@�?=�>=T�==o==8><=�g;=k�:=��9=v�8=��7=�7=}>6=)\5=�w4=đ3=��2=�1=��0=��/=r�.=��-=�-=,=�+=�*=�)=*(=�'=�&=.�$=P�#=2�"=ӻ!=� =�=:d=@=:=��=��=��=�S=e=��=��=nR=D=�=h=�=۷=�Y
=��=�=(=K�=�H=A�=Z =;��<���<���<��<^��<�l�<�H�<8�<7��<��<�x�<�5�<���<c��<�J�<��<���<82�<a��<R`�<�<~�<O�<��<��<��<��<̅�<u��<�r�<O�<X�<Ȓ<�6�<S��< �<�|�<(�<y�z<5|s<@Rl<�(e<~ ^<r�V<Y�O<��H<%qA<T:<::3<�$,<�%<<|�<>�< 	<#
<26�;?f�;���;���;�T�;AƱ;�I�;���;Ƌ�;f�x;@^;�D;�*;�L;Qa�:���:��:�-,:��99˸~���r[�䑝���̺�����'��#,���B��`Y�e�o��т�沍�Lt�����W��������:»�\̻3_ֻHB����:1���L������~�ƈ���=Q���"�A�&��+� A/��\3��l7��p;��h?��UC��7G��K���N���R�yWV�DZ���]�FKa�W�d�3mh��k�Woo�H�r��Sv��y�k}�T<���恼�����3���Ն��u��C��v���|G��tގ��s�����;���(��f���LC���Ι�-Y��P✼qj�����w��#���ҁ�����D���R��ӎ��������������,��陳����������������%������-���  �  �hN=0�M=�L=�L=�[K=#�J=�I=|I=9FH=LG=��F==�E=&E=\D=
�C=1�B=P�A=_*A=d[@=B�?=�>=X�==o==6><=�g;=f�:=��9=y�8=��7=�7=s>6='\5=�w4=Ñ3=�2="�1=��0=��/=z�.=��-=�-=,=�+=�*=�)=-(=�'=�&=/�$=R�#=7�"=ѻ!=� =�=@d=@=6=��=��=��=�S=i= �=��=pR=C=�= h=�=ٷ=�Y
=��=ߑ=(=L�=�H=C�=Z =9��<��<���<��<a��<�l�<�H�<5�<,��<��<�x�<�5�<���<i��<�J�<��<w��<82�<n��<A`�<�<~�<D�<��<��<"��<��<υ�<u��<�r�<L�<�W�<Ȓ<�6�<V��<��<�|�<9�<u�z<0|s<VRl<�(e<y ^<��V<=�O<j�H<,qA<T:<M:3<t$,<�%<2<z�<@�<! 	<7
<66�;Jf�;f��;���;�T�;�ű;J�;���;���;Y�x;8@^;)D;$*;�L;a�:�:W�:�,,:��9�˸ʺ���t[�����̺����'�P#,���B��`Y��o�҂����Kt�����<��������:»�\̻%_ֻ=B�����I1���L����ʇ���ֈ����>Q��"�I�&��+��@/��\3��l7��p;��h?��UC��7G��K���N���R��WV�-Z���]�HKa�O�d�4mh��k�Ioo�C�r�Tv��y�q}�R<���恼�����3���Ն��u��=��p���wG��vގ��s�����.���(��c���EC���Ι�+Y��O✼ej��~��w��"���ʁ�����R���J��׎��������������.��왳����������������%�����-���  �  �hN=3�M=�L=�L=�[K= �J=�I=wI=:FH=MG=��F=@�E=&E=\D=�C=/�B=I�A=f*A=e[@=C�?=�>=S�==u==2><=�g;=f�:=��9=z�8=��7=�7=u>6=.\5=�w4=��3=��2=�1=��0=��/=z�.=��-=�-=,=�+=�*=�)=1(=�'=�&=1�$=M�#=:�"=ѻ!=� =�=;d=@=9=��=��=��=�S=m=��=��=uR=?= �=�g=�=׷=�Y
=��=�=
(=D�=�H=A�=Z =7��<���<���<��<h��<�l�<�H�<9�<)��<���<�x�<�5�<���<g��<�J�<��<���<*2�<g��<M`�<�<~�<F�<��<��<%��<��<م�<r��<�r�<U�<�W�<Ȓ<�6�<V��<��<�|�<1�<Z�z<E|s<BRl<�(e<d ^<u�V<\�O<u�H<2qA<�S:<X:3<r$,<�%<#<n�<Z�< 	<<
<;6�;^f�;{��;���;�T�;*Ʊ;�I�;���;���;e�x;I@^;+D;�*;M;�`�:̋�:h�:-,:��9�˸¸��!t[�<�����̺z����'��#,���B�zaY��o��т�벍�Zt����� ��������:»�\̻_ֻ-B�%�ߪ�N1���L����އ�|�Ɉ����UQ��"�L�&�}+�
A/��\3��l7��p;��h?��UC��7G��K���N�}�R��WV�'Z���]�DKa�W�d�,mh��k�eoo�-�r�Tv���y��}�Q<���恼�����3���Ն��u��D��r���tG��uގ�~s�����4���(��b���RC���Ι�$Y��Q✼cj���񟼵w��&���Ӂ�����S���D��ߎ��������������<��ᙳ����������������%�����-���  �  �hN=,�M=�L=�L=�[K= �J=�I={I=8FH=JG=��F=F�E=&E=�[D=�C=*�B=Q�A=i*A=_[@=?�?=�>=W�==r==3><=�g;=k�:=��9=v�8=��7=�7=v>6=*\5=�w4=Ƒ3=��2=�1=��0=��/=r�.=��-=�-=,=�+=�*=�)=/(=�'=�&=1�$=Q�#=6�"=ϻ!=� =�=;d=@=:=��=��=��=�S=j= �=��=rR=B=�=h=�=ط=�Y
=��=�=(=K�=�H=>�=Z =A��<���<���<��<c��<�l�<�H�<5�<3��<��<�x�<�5�<���<j��<�J�<��<���<<2�<b��<W`�<�<~�<T�<��<��<��<��<Յ�<p��<�r�<V�<�W�<Ȓ<�6�<U��<��<�|�<$�<t�z<L|s<&Rl<�(e<~ ^<f�V<U�O<q�H</qA<T:<>:3<�$,<%<<n�<O�< 	<3
<)6�;f�;���;���;�T�;SƱ;�I�;���;ڋ�;�x;@^;1D;*;�L;�`�:6��:��:;-,:U�9˸Z����s[�ב����̺�����'��#,�A�B�aY�Z�o��т�����Lt�����J��������:»�\̻"_ֻ-B�����[1���L����އ���ǈ����7Q���"�U�&��+��@/��\3��l7��p;��h?��UC��7G��K���N���R��WV�@Z���]�1Ka�e�d�4mh��k�\oo�C�r�Tv���y�n}�V<���恼�����3���Ն��u��?��o���zG���ގ�|s�����:���(��h���HC���Ι�3Y��U✼jj���񟼺w��(���ց�����K���Q��Վ��������������/��ޙ�����������������%�����-���  �  �hN=,�M=�L=�L=�[K='�J=�I=~I=6FH=SG=��F=@�E=&E= \D=�C=+�B=R�A=`*A=h[@=E�?=�>=Y�==n==:><=�g;=h�:=��9=t�8=��7=�7=v>6=)\5=�w4=3=��2= �1=��0=��/=w�.=��-=�-=,=�+=�*=�)=((=�'=�&=1�$=S�#=5�"=ڻ!=� =�=<d=@=9=��=��=��=�S=j=�=��=oR=H=�=h=�=ַ=�Y
=��=�=(=K�=�H=C�=Z =7��<��<���<���<X��<�l�<�H�<2�</��<��<�x�<5�<���<i��<�J�<(��<v��<;2�<a��<L`�<�<~�<J�<��<��<��<��<υ�<|��<�r�<G�<X�<Ȓ<�6�<M��<��<�|�<4�<q�z<8|s<ORl<�(e<u ^<��V<P�O<m�H<qA< T:<>:3<�$,<�%<)<��<<�<' 	<+
<k6�;Qf�;���;���;�T�;&Ʊ;�I�;�;���;��x;v@^;D;;*;�L;�a�:G��:��:-,:��9�˸�����s[�呝�M�̺-����'�u#,���B�aY��o��т����_t�����Q��������:»�\̻!_ֻ.B�����1���L����ڇ���ʈ����>Q��"�+�&��+��@/��\3��l7�rp;��h?��UC��7G��K���N���R��WV�4Z���]�QKa�Q�d�0mh��k�Poo�?�r� Tv��y�v}�Y<���恼�����3���Ն��u��9��q���qG��jގ��s�����:���(��h���FC���Ι�+Y��A✼lj��|��w�����́�����H���O��܎��������������0��虳����������������%�����-���  �  �hN=2�M=�L=�L=�[K=!�J=�I=yI=5FH=HG=��F=B�E=&E=\D=�C=1�B=P�A=e*A=g[@==�?=�>=T�==s==4><=�g;=h�:=��9=|�8=��7=�7=v>6=+\5=�w4=��3=��2=�1=��0=��/=y�.=��-=�-=,=�+=�*=�)=-(=�'=�&=0�$=O�#=3�"=ѻ!=� =�==d=@=8=��=��=��=�S=e=��=��=nR=B=�= h=�=۷=�Y
=��=�=	(=G�=�H=@�=Z =6��<���<���<��<m��<�l�<�H�<;�</��<��<�x�<�5�<���<d��<�J�<!��<���<72�<k��<D`�<$�<~�<K�<��<��<��<��<ԅ�<t��<�r�<S�<�W�<Ȓ<�6�<_��<��<�|�<4�<_�z<@|s<9Rl<�(e<e ^<��V<O�O<y�H<@qA<�S:<W:3<�$,<�%<&<s�<L�< 	<*
<6�;^f�;���;���;�T�;�ű;J�;���;���;��x;�?^;D;�*;�L;�`�:���:��:�-,:R�9�˸����s[�����c�̺g����'��#,���B�NaY��o��т�಍�3t�����)��������:»�\̻2_ֻ5B����L1���L����ԇ�}�Ј����BQ��"�H�&��+�A/��\3��l7��p;��h?��UC��7G��K���N�u�R��WV�+Z���]�CKa�\�d�6mh��k�Zoo�7�r�Tv��y�y}�K<���恼�����3���Ն��u��A��u����G��rގ��s�����1���(��^���HC���Ι�$Y��V✼mj���񟼻w��#���ρ�����L���E��������
����������9��䙳����������������%�� ���-���  �  �hN=2�M=�L=�L=�[K=!�J=�I=vI=BFH=JG=��F=E�E=
&E=\D=�C=2�B=K�A=i*A=a[@=B�?=�>=Q�==x==0><=�g;=i�:=��9=z�8=��7=�7=n>6=,\5=�w4=đ3=��2=�1=��0=��/=y�.=��-=�-=
,=�+=�*=�)=2(=�'=�&=2�$=Q�#=>�"=ͻ!=� =�=;d=@=8=��=��=��=�S=p=�=��=tR=?= �=�g=�=ٷ=�Y
=��=ݑ=
(=F�=�H=<�=Z =>��<���<���<��<d��<�l�<�H�</�<,��<���<�x�<�5�<���<v��<�J�<��<���<-2�<n��<J`�<!�<~�<O�<��<��<3��<��<ۅ�<v��<�r�<Z�<�W�<Ȓ<�6�<S��<��<�|�<-�<b�z<Z|s<Rl<�(e<l ^<q�V<U�O<Y�H<)qA<�S:<T:3<e$,<%<"<r�<_�< 	<]
<#6�;Ef�;���;���;�T�;Ʊ;J�;���;ڋ�;/�x;;@^;�D;�*;JM;_`�:ы�:��:G,,:��9�˸ֹ���u[�r�����̺�����'�$,�"�B�LaY��o�҂����pt�����@��������:»�\̻_ֻ(B�껼��k1���L����܇�}�̈����PQ��"�[�&�n+��@/��\3��l7��p;��h?��UC��7G��K���N���R��WV�'Z���]�,Ka�l�d�2mh��k�boo�2�r�!Tv���y��}�O<���恼�����3���Ն��u��F��c���rG��|ގ�ys�����.���(��`���PC���Ι�'Y��V✼Uj���񟼴w��"���Ձ�����Y���F������������������8��֙�����������������%�����-���  �  �hN=0�M=�L=�L=�[K=$�J=�I=xI=6FH=MG=��F=C�E=&E=\D=�C=.�B=N�A=e*A=e[@=@�?=�>=S�==o==6><=�g;=i�:=��9=z�8=��7=�7=y>6=-\5=�w4=��3=��2=�1=��0=��/=y�.=��-=�-=,=�+=�*=�)=,(=�'=�&=,�$=M�#=4�"=һ!=� =�=:d=	@=;=��=��=��=�S=g=��=��=oR=D=�=h=�=ݷ=�Y
=��=�=	(=F�=�H=@�=Z =3��<���<���<���<b��<�l�<�H�<3�<2��<��<�x�<�5�<���<b��<�J�<��<���<32�<e��<Q`�<�<~�<O�<��<��<��<��<ʅ�<w��<�r�<N�<�W�<Ȓ<�6�<Q��<��<�|�<.�<a�z<>|s<DRl<�(e<k ^<r�V<a�O<|�H<'qA<T:<L:3<{$,<�%<#<��<=�< 	<-
<A6�;Vf�;���;���;�T�;9Ʊ;�I�;���;���;g�x;%@^;D;�*;�L;a�:\��:��:-,:E�9�˸����6s[�n�����̺t����'��#,���B�PaY��o��т�߲��[t�����O��������:»�\̻,_ֻTB�'���A1���L������w�������FQ���"�G�&��+�A/�]3��l7��p;��h?��UC��7G��K���N�|�R��WV�(Z���]�KKa�[�d�1mh�$�k�boo�2�r��Sv���y�q}�L<���恼�����3���Ն��u��E��w���{G��uގ��s�����6���(��f���OC���Ι�(Y��M✼mj�����w�� ���Ӂ�����L���L��Ҏ����	����������8��䙳����������������%������-���  �  �hN=(�M="�L=�L=�[K=$�J=�I=�I=2FH=LG=��F=A�E=&E= \D=�C=+�B=X�A=d*A=g[@=>�?=�>=g�==l==9><=�g;=j�:=��9=s�8=��7=�7=y>6='\5=�w4=Ñ3=}�2="�1=��0=��/=u�.=��-=�-=,=�+=�*=�)=+(=�'=�&=6�$=]�#=2�"=׻!=� =�=9d=@=8=��=��=��=�S=e=�=��=lR=I=�=h=�=ط=�Y
=��=��=(=N�=�H=C�=Z =8��<
��<���<���<R��<�l�<�H�<3�<5��<��<�x�<z5�<���<l��<�J�<&��<���<G2�<a��<N`�<�<~�<Q�<��<��<��<��<х�<v��<�r�<M�<X�<�ǒ<�6�<K��<��<�|�<0�<{�z<%|s<VRl<�(e<~ ^<}�V<>�O<|�H<qA<T:<,:3<�$,<�%<"<|�<<�<\ 	<
<96�;Rf�;���;���;�T�;,Ʊ;�I�;.�;���;��x; @^;#D;*;�L;{a�:���:��:�-,:��9�˸ӽ���r[������̺	��� (�V#,���B��`Y�0�o�҂�����t�����{��������:»{\̻8_ֻB໧���1���L��������͈���&Q���"�.�&��+��@/��\3��l7�kp;��h?��UC��7G��K���N���R��WV�<Z���]�IKa�O�d�6mh��k�Aoo�G�r��Sv��y�|}�[<���恼�����3���Ն��u��"��m����G��lގ��s�����;���(��g���FC���Ι�*Y��L✼tj��_񟼾w��"���́�����>���[��؎��"������������+��񙳼���������������%������-���  �  �hN=0�M=�L=�L=�[K=$�J=�I=xI=6FH=MG=��F=C�E=&E=\D=�C=.�B=N�A=e*A=e[@=@�?=�>=S�==o==6><=�g;=i�:=��9=z�8=��7=�7=y>6=-\5=�w4=��3=��2=�1=��0=��/=y�.=��-=�-=,=�+=�*=�)=,(=�'=�&=,�$=M�#=4�"=һ!=� =�=:d=	@=;=��=��=��=�S=g=��=��=oR=D=�=h=�=ݷ=�Y
=��=�=	(=F�=�H=@�=Z =3��<���<���<���<b��<�l�<�H�<3�<2��<��<�x�<�5�<���<b��<�J�<��<���<32�<e��<Q`�<�<~�<O�<��<��<��<��<ʅ�<w��<�r�<N�<�W�<Ȓ<�6�<Q��<��<�|�<.�<a�z<>|s<DRl<�(e<k ^<r�V<a�O<|�H<'qA<T:<L:3<{$,<�%<#<��<=�< 	<-
<A6�;Vf�;���;���;�T�;9Ʊ;�I�;���;���;g�x;%@^;D;�*;�L;a�:\��:��:-,:E�9�˸����6s[�n�����̺t����'��#,���B�PaY��o��т�߲��[t�����O��������:»�\̻,_ֻTB�'���B1���L������w�������FQ���"�G�&��+�A/�]3��l7��p;��h?��UC��7G��K���N�|�R��WV�(Z���]�KKa�[�d�1mh�$�k�boo�2�r��Sv���y�q}�L<���恼�����3���Ն��u��E��w���{G��uގ��s�����6���(��f���OC���Ι�(Y��M✼mj�����w�� ���ҁ�����L���L��Ҏ����	����������8��䙳����������������%������-���  �  �hN=2�M=�L=�L=�[K=!�J=�I=vI=BFH=JG=��F=E�E=
&E=\D=�C=2�B=K�A=i*A=a[@=B�?=�>=Q�==x==0><=�g;=i�:=��9=z�8=��7=�7=n>6=,\5=�w4=đ3=��2=�1=��0=��/=y�.=��-=�-=
,=�+=�*=�)=2(=�'=�&=2�$=Q�#=>�"=ͻ!=� =�=;d=@=8=��=��=��=�S=p=�=��=tR=?= �=�g=�=ٷ=�Y
=��=ݑ=
(=F�=�H=<�=Z =>��<���<���<��<d��<�l�<�H�</�<,��<���<�x�<�5�<���<v��<�J�<��<���<-2�<n��<J`�<!�<~�<O�<��<��<3��<��<ۅ�<v��<�r�<Z�<�W�<Ȓ<�6�<S��<��<�|�<-�<b�z<Z|s<Rl<�(e<l ^<q�V<U�O<Y�H<)qA<�S:<T:3<e$,<%<"<r�<_�< 	<]
<#6�;Ef�;���;���;�T�;Ʊ;J�;���;ڋ�;/�x;;@^;�D;�*;JM;_`�:Ћ�:��:G,,:��9�˸ع���u[�s�����̺�����'�$,�"�B�MaY��o�҂����pt�����@��������:»�\̻_ֻ(B�껼��k1���L����܇�}�̈����PQ��"�[�&�n+��@/��\3��l7��p;��h?��UC��7G��K���N���R��WV�'Z���]�,Ka�l�d�2mh��k�boo�2�r�!Tv���y��}�O<���恼�����3���Ն��u��F��c���rG��|ގ�ys�����.���(��`���PC���Ι�'Y��V✼Uj���񟼴w��"���Ձ�����Y���F������������������8��֙�����������������%�����-���  �  �hN=2�M=�L=�L=�[K=!�J=�I=yI=5FH=HG=��F=B�E=&E=\D=�C=1�B=P�A=e*A=g[@==�?=�>=T�==s==4><=�g;=h�:=��9=|�8=��7=�7=v>6=+\5=�w4=��3=��2=�1=��0=��/=y�.=��-=�-=,=�+=�*=�)=-(=�'=�&=0�$=O�#=3�"=ѻ!=� =�==d=@=8=��=��=��=�S=e=��=��=nR=B=�= h=�=۷=�Y
=��=�=	(=G�=�H=@�=Z =6��<���<���<��<m��<�l�<�H�<;�</��<��<�x�<�5�<���<d��<�J�<!��<���<72�<k��<D`�<$�<~�<K�<��<��<��<��<ԅ�<t��<�r�<S�<�W�<Ȓ<�6�<_��<��<�|�<4�<_�z<@|s<9Rl<�(e<e ^<��V<O�O<y�H<@qA<�S:<W:3<�$,<�%<&<s�<L�< 	<*
<6�;^f�;���;���;�T�;�ű;J�;���;���;��x;�?^;D;�*;�L;�`�:���:��:�-,:P�9�˸����s[�����c�̺g����'��#,���B�NaY��o��т�಍�3t�����)��������:»�\̻2_ֻ5B����L1���L����ԇ�}�Ј����BQ��"�H�&��+�A/��\3��l7��p;��h?��UC��7G��K���N�u�R��WV�+Z���]�CKa�\�d�6mh��k�Zoo�7�r�Tv��y�y}�K<���恼�����3���Ն��u��A��u����G��rގ��s�����1���(��^���HC���Ι�$Y��V✼mj���񟼻w��#���ρ�����L���E��������
����������9��䙳����������������%�� ���-���  �  �hN=,�M=�L=�L=�[K='�J=�I=~I=6FH=SG=��F=@�E=&E= \D=�C=+�B=R�A=`*A=h[@=E�?=�>=Y�==n==:><=�g;=h�:=��9=t�8=��7=�7=v>6=)\5=�w4=3=��2= �1=��0=��/=w�.=��-=�-=,=�+=�*=�)=((=�'=�&=1�$=S�#=5�"=ڻ!=� =�=<d=@=9=��=��=��=�S=j=�=��=oR=H=�=h=�=ַ=�Y
=��=�=(=K�=�H=C�=Z =7��<��<���<���<X��<�l�<�H�<2�<0��<��<�x�<5�<���<i��<�J�<(��<v��<;2�<a��<L`�<�<~�<J�<��<��<��<��<υ�<|��<�r�<G�<X�<Ȓ<�6�<M��<��<�|�<4�<q�z<8|s<ORl<�(e<u ^<��V<P�O<m�H<qA< T:<>:3<�$,<�%<)<��<<�<' 	<+
<k6�;Qf�;���;���;�T�;&Ʊ;�I�;�;���;��x;v@^;D;;*;�L;�a�:G��:��:-,:��9�˸�����s[�呝�M�̺-����'�v#,���B�aY��o��т����_t�����Q��������:»�\̻!_ֻ.B�����1���L����ڇ���ʈ����>Q��"�+�&��+��@/��\3��l7�rp;��h?��UC��7G��K���N���R��WV�4Z���]�QKa�Q�d�0mh��k�Poo�?�r� Tv��y�v}�Y<���恼�����3���Ն��u��9��q���qG��jގ��s�����:���(��h���FC���Ι�+Y��A✼lj��|��w�����́�����H���O��܎��������������0��虳����������������%�����-���  �  �hN=,�M=�L=�L=�[K= �J=�I={I=8FH=JG=��F=F�E=&E=�[D=�C=*�B=Q�A=i*A=_[@=?�?=�>=W�==r==3><=�g;=k�:=��9=v�8=��7=�7=v>6=*\5=�w4=Ƒ3=��2=�1=��0=��/=r�.=��-=�-=,=�+=�*=�)=/(=�'=�&=1�$=Q�#=6�"=ϻ!=� =�=;d=@=:=��=��=��=�S=j= �=��=rR=B=�=h=�=ط=�Y
=��=�=(=K�=�H=>�=Z =A��<���<���<��<c��<�l�<�H�<5�<3��<��<�x�<�5�<���<j��<�J�<��<���<<2�<b��<W`�<�<~�<T�<��<��<��<��<Յ�<p��<�r�<V�<�W�<Ȓ<�6�<U��<��<�|�<$�<t�z<L|s<&Rl<�(e<~ ^<f�V<U�O<q�H</qA<T:<>:3<�$,<%<<n�<O�< 	<3
<)6�;f�;���;���;�T�;SƱ;�I�;���;ڋ�;�x;@^;1D;*;�L;�`�:6��:��::-,:R�9˸^����s[�ؑ����̺�����'��#,�A�B�aY�Z�o��т�����Lt�����J��������:»�\̻"_ֻ-B�����[1���L����އ���ǈ����7Q���"�U�&��+��@/��\3��l7��p;��h?��UC��7G��K���N���R��WV�@Z���]�1Ka�e�d�4mh��k�\oo�C�r�Tv���y�n}�V<���恼�����3���Ն��u��?��o���zG���ގ�|s�����:���(��h���HC���Ι�3Y��U✼jj���񟼺w��(���ց�����K���Q��Վ��������������/��ޙ�����������������%�����-���  �  �hN=3�M=�L=�L=�[K= �J=�I=wI=:FH=MG=��F=@�E=&E=\D=�C=/�B=I�A=f*A=e[@=C�?=�>=S�==u==2><=�g;=f�:=��9=z�8=��7=�7=u>6=.\5=�w4=��3=��2=�1=��0=��/=z�.=��-=�-=,=�+=�*=�)=1(=�'=�&=1�$=M�#=:�"=ѻ!=� =�=;d=@=9=��=��=��=�S=m=��=��=uR=?= �=�g=�=׷=�Y
=��=�=
(=D�=�H=A�=Z =7��<���<���<��<h��<�l�<�H�<9�<)��<���<�x�<�5�<���<g��<�J�<��<���<*2�<g��<M`�<�<~�<F�<��<��<%��<��<م�<r��<�r�<U�<�W�<Ȓ<�6�<V��<��<�|�<1�<Z�z<E|s<BRl<�(e<d ^<u�V<\�O<u�H<2qA<�S:<X:3<r$,<�%<#<n�<Z�< 	<<
<;6�;^f�;{��;���;�T�;*Ʊ;�I�;���;���;d�x;I@^;+D;�*;M;�`�:ˋ�:h�:
-,:��9�˸Ÿ��"t[�=�����̺{����'��#,���B�{aY��o��т�벍�Zt����� ��������:»�\̻_ֻ-B�%�ߪ�N1���L����އ�|�Ɉ����UQ��"�L�&�}+�
A/��\3��l7��p;��h?��UC��7G��K���N�}�R��WV�'Z���]�DKa�W�d�,mh��k�doo�-�r�Tv���y��}�Q<���恼�����3���Ն��u��D��r���tG��uގ�~s�����4���(��b���RC���Ι�$Y��Q✼cj���񟼵w��&���Ӂ�����S���D��ߎ��������������<��ᙳ����������������%�����-���  �  �hN=0�M=�L=�L=�[K=#�J=�I=|I=9FH=LG=��F==�E=&E=\D=
�C=1�B=P�A=_*A=d[@=B�?=�>=X�==o==6><=�g;=f�:=��9=y�8=��7=�7=s>6='\5=�w4=Ñ3=�2="�1=��0=��/=z�.=��-=�-=,=�+=�*=�)=-(=�'=�&=/�$=R�#=7�"=ѻ!=� =�=@d=@=6=��=��=��=�S=i= �=��=pR=C=�= h=�=ٷ=�Y
=��=ߑ=(=L�=�H=C�=Z =9��<��<���<��<a��<�l�<�H�<5�<,��<��<�x�<�5�<���<i��<�J�<��<w��<82�<n��<A`�<�<~�<D�<��<��<"��<��<υ�<u��<�r�<L�<�W�<Ȓ<�6�<V��<��<�|�<9�<u�z<0|s<VRl<�(e<y ^<��V<=�O<j�H<,qA<T:<N:3<t$,<�%<2<z�<@�<! 	<7
<66�;Jf�;f��;���;�T�;�ű;J�;���;���;Y�x;8@^;)D;$*;�L;a�:���:W�:�,,:��9�˸ͺ���t[�����̺����'�P#,���B��`Y��o�҂����Kt�����<��������:»�\̻%_ֻ=B�����I1���L����ʇ���ֈ����>Q��"�I�&��+��@/��\3��l7��p;��h?��UC��7G��K���N���R��WV�-Z���]�HKa�O�d�4mh��k�Ioo�C�r�Tv��y�q}�R<���恼�����3���Ն��u��=��p���wG��vގ��s�����.���(��c���EC���Ι�+Y��O✼ej��~��w��"���ʁ�����R���J��׎��������������.��왳����������������%�����-���  �  �hN=+�M= �L=�L=�[K=#�J=�I=zI=4FH=KG=��F=D�E=&E= \D=�C=,�B=P�A=g*A=e[@=@�?=�>=T�==o==8><=�g;=k�:=��9=v�8=��7=�7=}>6=)\5=�w4=đ3=��2=�1=��0=��/=r�.=��-=�-=,=�+=�*=�)=*(=�'=�&=.�$=P�#=2�"=ӻ!=� =�=:d=@=:=��=��=��=�S=e=��=��=nR=D=�=h=�=۷=�Y
=��=�=(=K�=�H=A�=Z =;��<���<���<��<^��<�l�<�H�<8�<7��<��<�x�<�5�<���<c��<�J�<��<���<82�<a��<R`�<�<~�<O�<��<��<��<��<̅�<u��<�r�<O�<X�<Ȓ<�6�<S��< �<�|�<(�<y�z<5|s<@Rl<�(e<~ ^<r�V<Y�O<��H<%qA<T:<::3<�$,<�%<<|�<>�< 	<#
<26�;?f�;���;���;�T�;AƱ;�I�;���;Ƌ�;f�x;@^;�D;�*;�L;Qa�:���:��:�-,:��9C˸����r[�䑝���̺�����'��#,���B��`Y�f�o��т�沍�Mt�����X��������:»�\̻3_ֻHB����:1���L������~�ƈ���=Q���"�A�&��+� A/��\3��l7��p;��h?��UC��7G��K���N���R�yWV�DZ���]�FKa�W�d�3mh��k�Woo�H�r��Sv��y�k}�T<���恼�����3���Ն��u��C��v���|G��tގ��s�����;���(��f���LC���Ι�-Y��P✼qj�����w��#���ҁ�����E���R��ӎ��������������,��陳����������������%������-���  �  �hN=0�M=�L=�L=�[K=#�J=�I=vI==FH=NG=��F=D�E=&E=\D=�C=.�B=K�A=g*A=b[@=C�?=�>=S�==u==5><=�g;=i�:=��9=x�8=��7=�7=s>6=.\5=�w4=đ3=��2=�1=��0=��/=y�.=��-=�-=,=�+=�*=�)=.(=�'=�&=5�$=Q�#=<�"=һ!=� =�=:d=@=8=��=��=��=�S=o=�=��=sR=B=�= h=�=ٷ=�Y
=��=�=
(=J�=�H=?�=Z ==��< ��<���<��<[��<�l�<�H�<3�<0��<��<�x�<�5�<���<q��<�J�<��<���</2�<f��<K`�<�<~�<O�<��<��<)��<��<ۅ�<x��<�r�<Q�<�W�<Ȓ<�6�<R��<��<�|�<0�<r�z<O|s<-Rl<�(e<w ^<|�V<\�O<`�H<"qA<�S:<L:3<v$,<�%<,<{�<Y�< 	<G
<E6�;Cf�;���;���;�T�;Ʊ;�I�;���;ȋ�;7�x;W@^;vD;�*;M;�`�:���:��:-,:o�9˸ƻ���t[�L�����̺�����'��#,�i�B�aY��o��т�#���ft�����C��������:»�\̻_ֻB��˪�E1���L���������ψ����LQ��"�J�&�t+��@/��\3��l7��p;��h?��UC��7G��K���N���R��WV�'Z���]�<Ka�a�d�)mh��k�Woo�/�r�Tv��y�|}�T<���恼�����3���Ն��u��A��i���rG��zގ�}s�����5���(��f���PC���Ι�)Y��O✼_j���񟼴w�����Ё�����Q���H��܎��������������0��ܙ�����������������%�����-���  �  �hN=4�M=�L=�L=�[K=�J=�I=uI=8FH=FG=��F=?�E=&E=\D=�C=4�B=L�A=e*A=b[@==�?=�>=S�==s==/><=�g;=f�:=��9={�8=��7=�7=r>6=-\5=�w4=��3=��2=�1=��0=��/=|�.=��-=�-=,=�+=�*=�)=1(=�'=�&=3�$=J�#=8�"=˻!=� =�=?d=@=5=��=��=��=�S=j=��=��=oR=?=!�=�g=�=ط=�Y
=��=ޑ=(=F�=�H=A�=Z =7��<���<���<��<s��<�l�<�H�<9�<*��<���<�x�<�5�<���<b��<�J�<��<���</2�<s��<<`�<$�<
~�<F�<��<��< ��<��<؅�<k��<�r�<U�<�W�<Ȓ<�6�<g��<��<�|�<8�<\�z<N|s<9Rl<�(e<e ^<��V<N�O<k�H<UqA<�S:<_:3<s$,<�%<5<a�<U�< 	<3
<6�;Pf�;x��;���;�T�;�ű;(J�;���;���;;�x;�?^;
D;�*;�L;0`�: ��:L�:[-,:��9[˸ѵ���t[�l���g�̺i����'��#,�Q�B�eaY�ġo��т�ݲ��$t�������������:»�\̻8_ֻ B�@���~1���L����͇���ۈ����OQ��"�a�&��+�A/��\3��l7��p;��h?��UC��7G��K���N�o�R��WV�Z���]�:Ka�Z�d�*mh��k�Yoo�-�r�Tv��y�v}�P<���恼�����3���Ն��u��B��w���|G��~ގ��s�����)���!(��^���JC���Ι�'Y��^✼gj���񟼷w��,���́�����V���>��㎪�������������;��ݙ�����������������%������,���  �  �hN=,�M=�L=�L=�[K="�J=�I=}I=7FH=OG=��F=?�E=&E=\D=�C=-�B=L�A=e*A=h[@=D�?=�>=Z�==q==6><=�g;=g�:=��9=s�8=��7=�7=w>6=,\5=�w4=��3=��2= �1=��0=��/=w�.=��-=�-=
,=�+=�*=�)=-(=�'=�&=5�$=Q�#=8�"=ջ!=� =�=9d=@=8=��=��=��=�S=l=��=��=oR=E=�=h=�=շ=�Y
=��=�=(=H�=�H=D�=Z =5��<��<���<���<\��<�l�<�H�<4�<.��<��<�x�<�5�<���<e��<�J�<$��<���</2�<c��<L`�<�<~�<E�<��<��<��<��<օ�<t��<�r�<P�<�W�<Ȓ<�6�<Q��<��<�|�<1�<k�z<=|s<IRl<�(e<p ^<�V<X�O<s�H<&qA<�S:<<:3<�$,<�%<"<t�<N�<$ 	<.
<L6�;_f�;t��;���;�T�;)Ʊ;�I�;���;���;��x;c@^;D;E*;�L;a�:@��:~�:d-,:�9�˸»���s[�����N�̺f����'�o#,���B�;aY��o��т����jt�����Q��������:»�\̻0_ֻB����/1���L��������͈���QQ��"�<�&�+�A/��\3��l7�p;��h?��UC��7G��K���N���R��WV�1Z���]�HKa�M�d�)mh� �k�Qoo�:�r� Tv��y��}�\<���恼�����3���Ն��u��6��u���pG��nގ��s�����9���(��d���PC���Ι�&Y��J✼ij��~񟼹w��$���Ё�����J���Q��ގ��������������3��噳����������������%�����-���  �  �jN=K�M=��L=^"L=�^K=��J=��I=�I=�JH=�G=��F=��E=�+E=/bD=��C=�B=��A=%2A=�c@=Փ?=��>=��==S==�H<=Tr;=��:=|�9=��8=Y
8=',7=FL6=uj5=̆4=!�3=n�2=��1=��0=C�/=�/=�.=-=�#,=0)+=�+*=o+)=@((=6"'=&=�%=��#=��"=�!=�� =�=�~=[=�3=�=��=�=�p=]6=.�=�=�o=�%=��=��=�/=��=hw
=E	=+�=E=�=2e=v�=�u =��<��<���<��<g��<���<�y�<�M�<�<���<R��<�_�<��<���<�p�<e�<D��<}S�<��<g~�<��<㘹<� �<���<�%�<a��<}�<ϖ�<��<���<_�<mb�<�В<>�<թ�<��<�<��<H�z<�vs<�Il<�e<A�]<��V<��O<�xH<�TA<�4:<x3<��+<��$<��<��<p�<-�<��<{��;��;p �;li�;�¾;�.�;��;t=�;'�;a7w;9�\;��B;��(;f�;�8�:N�:�̈́:7h%:!�9�����o�b�B���к�����d.���D��V[�֚q�σ�����r��G��e������{8û2YͻnZ׻�;��������$��*��{h�N��H�����@d�~��m#��M'�р+��/���3�N�7���;���?�A�C��G��dK�6/O���R�i�V��SZ���]�.�a��%e�w�h�,3l�%�o��!s�a�v�^�y��S}�gV�� �������J��솼����'������Z��+���]������s���o6��Ė�)P���ڙ��d��휼st������d�����������M����������<���������꘰�������2������M��R����#������*���  �  �jN=T�M=��L=_"L=�^K=��J=��I=�I=�JH=�G=üF=��E=�+E=1bD=��C=!�B=��A=$2A=�c@=ړ?=��>=��==T==�H<=Xr;=��:=��9=��8=H
8=#,7=AL6=yj5=І4=&�3=o�2=��1=��0=C�/=�/=�.=-=�#,=%)+=�+*=n+)=E((=4"'=&=�%=��#=��"=�!=ǻ =�=�~=[=�3=�=��=�=�p=e6=2�=�=�o=�%=��=��=�/=��=Yw
=A	=(�=E=�=8e=u�=�u =$��<��<���<��<b��<מ�<�y�<�M�<|�<���<F��<�_�<��<���<�p�<u�<F��<iS�<��<V~�<��<ژ�<� �<���<�%�<p��<y�<Җ�<��<���<b�<nb�<�В<�=�<©�<��<�<��<M�z<�vs<�Il<�e<H�]<�V<��O<�xH<�TA<�4:<�3<��+<��$<��<��<t�<%�<�<���;X��;G �;1i�;�¾;\.�;(��;$=�;�;�7w;{�\;J�B;s�(;w�;�7�:�N�:~̈́:Dj%:�"�9-����÷b��A����к�����.�a�D��V[�J�q�%σ�"���@s������������T8ûAYͻ�Z׻�;���껭����$�����h�T��R�����?d����W#��M'���+���/���3�T�7���;���?�H�C��G��dK�u/O���R�r�V��SZ���]��a��%e�u�h�3l��o��!s�r�v�j�y��S}�hV�����������J��솼����'�������Y�����Z������m���6��Ė�2P���ڙ��d���으ct������a�����������L����������O���������ܘ��������:������J��F����#������*���  �  �jN=Y�M=��L=["L=�^K=��J=��I=�I=�JH=�G=ļF=��E=�+E=:bD=��C=,�B=��A='2A=�c@=ғ?=��>=��==[==�H<=_r;=��:=��9=��8=M
8=2,7=<L6=zj5=ˆ4="�3=l�2=��1=��0==�/=�/=�.=-=�#,=&)+=�+*=c+)=I((=3"'=&=�%=��#=��"=�!=ͻ =�=�~=[=�3=�=��=!�=�p=`6=(�=
�=�o=�%=��=��=�/=��=cw
=J	=$�=E=�=8e=q�=�u =��<���<���<��<~��<��<�y�<�M�<l�<���<B��<�_�<x�<���<�p�<i�<L��<eS�<��<P~�<��<☹<~ �<���<�%�<l��<f�<ܖ�<��<���<`�<[b�<�В<�=�<ߩ�<��<�<��<8�z<�vs<�Il<�e<8�]<�V<��O<�xH<UA<�4:<�3<��+<��$<��<��<��<�<�<V��;b��;H �;?i�;Aþ;;.�;���;=�;1�;�7w;��\;�B;�(;��;�7�:mO�:�̄:i%:e$�9�����̸b�uA��6�кQ���5��.�T�D��V[��q�Fσ�ﰎ��r�����ҕ��b���58ûIYͻpZ׻�;�$��̠���$������h�3��L�����d����C#��M'�Ȁ+�#�/���3�C�7���;���?�p�C�ޏG��dK�M/O���R���V��SZ���]��a��%e���h�!3l�6�o��!s���v�1�y��S}�dV�����������J��솼�����'������Z��&���U������W����6�� Ė�*P�� ۙ��d��휼gt������W�����������`����������1���������٘��������C������R��F����#�������)���  �  �jN=R�M=��L=^"L=�^K=��J=��I=�I=�JH=�G=��F=��E=�+E=3bD=��C="�B=��A=)2A=�c@=ٓ?=��>=��==Z==�H<=\r;=��:=��9=��8=O
8=',7=:L6=|j5=͆4=%�3=n�2=��1=��0=C�/=�/=�.= -=�#,=')+=�+*=k+)=I((=1"'=&=�%=��#=��"=�!=˻ =�=�~=[=�3=�=��= �=�p=f6=0�=�=�o=�%=��=��=�/=��=aw
=?	=%�=E=�=7e=u�=�u =��<��<���<��<e��<��<�y�<�M�<w�<���<>��<�_�<|�<���<�p�<i�<P��<fS�<��<Y~�<��<ؘ�<� �<���<�%�<z��<q�<ٖ�<��<���<g�<hb�<�В<�=�<ҩ�<��<	�<��<K�z<�vs<�Il<�e<E�]<
�V<��O<nxH<�TA<�4:<�3<��+<��$<��<��<��<�<�<���;K��;[ �;"i�;þ;e.�;2��;=�;B�;�7w;m�\;v�B;,�(;��;�7�:O�:<̈́:Oi%:s"�9 ����`�b�;A���к����z.�^�D��V[�I�q�>σ�E����r��������#���/8û\YͻvZ׻�;���껚����$������h�R��L�����>d����H#��M'���+��/���3�H�7���;���?�Q�C��G��dK�S/O���R��V��SZ���]��a��%e�w�h�3l�"�o��!s���v�c�y��S}�iV��  �������J��"솼����'�������Y��&���Q������m���}6��	Ė�5P���ڙ��d��휼Zt������Z�����#���~��R����������?���������ޘ��������<������K��J����#������*���  �  �jN=O�M=��L=\"L=�^K=��J=��I=�I=�JH=�G=��F=��E=�+E=2bD=��C= �B=��A='2A=�c@=ԓ?=��>=��==W==�H<=Yr;=��:=��9=��8=P
8=&,7=FL6=zj5=ˆ4=$�3=i�2=��1=��0=E�/=�/=�.=-=�#,=))+=�+*=l+)=D((=6"'=&=�%=��#=��"=�!=Ȼ =�=�~=[=�3=�=��=�=�p=^6=.�=�=�o=�%=��=��=�/=��=`w
=B	=/�=E=�=3e=v�=�u =��<��<���<��<f��<��<�y�<�M�<w�<���<G��<�_�<��<���<�p�<l�<L��<rS�<��<a~�<��<ޘ�<� �<���<�%�<g��<t�<Ԗ�<��<���<_�<kb�<�В<�=�<ʩ�<��<�<��<T�z<�vs<�Il<�e<J�]<��V<��O<�xH<�TA<�4:<�3<��+<��$<��<��<~�<�<��<���;;��;\ �;Ei�;þ;�.�; ��;D=�;6�;�7w;%�\;�B;i�(;��;8�:�N�:̈́:�i%:!�9�����x�b��A��)�к���`�g.���D�wV[�Úq��΃����s�����������U8û3Yͻ~Z׻�;��������$��	���h�S��H�����Bd����Q#��M'�΀+��/���3�M�7���;���?�K�C���G��dK�W/O���R�W�V��SZ���]�*�a��%e���h�$3l�%�o��!s�]�v�a�y��S}�lV�����������J��솼����'������Z��#���U������q���t6��
Ė�.P���ڙ��d��휼mt������_�����������P����������G���������혰�������9������I��S����#������	*���  �  �jN=U�M=��L=\"L=�^K=��J=��I=�I=�JH=�G=üF=��E=�+E=4bD=��C='�B=��A=$2A=�c@=֓?=��>=��==V==�H<=]r;=��:=��9=��8=N
8=*,7=<L6=xj5=Ά4="�3=l�2=��1=��0=E�/=�/=�.=-=�#,=%)+=�+*=g+)=G((=4"'=&=�%=��#=��"=�!=Ȼ =�=�~=[=�3=�=��=�=�p=a6=0�=�=�o=�%=��=��=�/=~�=bw
=@	=$�=E=�=2e=w�=�u =��<��<���<��<k��<��<�y�<�M�<n�<���<C��<�_�<��<���<�p�<t�<F��<mS�<��<U~�<��<䘹< �<���<�%�<l��<t�<ږ�<��<���<_�<cb�<�В<�=�<ҩ�<��<�<��<R�z<�vs<�Il<�e<G�]<�V<��O<vxH<�TA<�4:<�3<��+<��$<��<��<��< �<�<���;X��;? �;Vi�;þ;Z.�;T��;5=�;�;�7w;A�\;Y�B;l�(;��;�7�:'O�:�̄:�i%:�!�9ɧ���ڸb��A���к[���:�B.���D�vV[�i�q�Hσ�3����r�����핮�?���D8û?Yͻ~Z׻�;����à���$�����h�D��V�����1d����U#��M'���+��/���3�J�7���;���?�`�C��G��dK�Q/O���R���V��SZ���]�,�a��%e�{�h�(3l�"�o��!s���v�U�y��S}�nV�����������J��솼����'������Z�����[������d����6��	Ė�(P�� ۙ��d��휼ht������Y�����������W����������?�������������������3������K��H����#������*���  �  �jN=V�M=��L=a"L=�^K=��J=��I=�I=�JH=	�G=ƼF=��E=�+E=3bD=��C=$�B=��A=,2A=�c@=ԓ?=��>=��==Z==�H<=`r;=��:=��9=��8=J
8=+,7=;L6=�j5=͆4="�3=m�2=��1=��0=@�/=�/=�.=-=�#,=#)+=�+*=f+)=M((=1"'=&=�%=��#=��"=�!=л =�=�~=[=�3=�=��=$�=�p=c6=0�=�=�o=�%=��=��=�/=�=cw
=B	='�=E=�=3e=s�=�u =��<��<���<��<m��<���<�y�<�M�<q�<���<>��<�_�<v�<���<�p�<p�<W��<iS�<
��<Y~�<��<ܘ�<� �<���<�%�<q��<i�<ږ�<��<���<l�<ab�<�В<�=�<֩�<��<�<��<<�z<�vs<�Il<�e<5�]<�V<��O<mxH<UA<{4:<�3<��+<��$<��<��<��<�<�<m��;s��;l �;3i�;
þ;e.�;<��; =�;Z�;�7w;"�\;f�B;��(;��;�7�:�O�:3̈́:�i%:C#�9\����4�b��@���кd���$��.���D��V[���q�-σ�0����r�����핮�G���8ûYYͻkZ׻�;���껸����$������h�M��L�����;d����4#��M'���+��/���3�D�7���;���?�f�C��G��dK�K/O���R�x�V��SZ���]�)�a��%e�{�h�'3l�+�o��!s���v�R�y��S}�hV�����������J��!솼 ����'������Z�� ���J������k���}6��Ė�0P���ڙ��d��	휼ct������Y��������y��Z����������:���������ؘ��������A������S��C����#�������)���  �  �jN=T�M=��L=_"L=�^K=��J=��I=�I=�JH=�G=��F=��E=�+E=2bD=��C=!�B=��A=&2A=�c@=Փ?=��>=��==Z==�H<=Yr;=��:=�9=��8=O
8=(,7=>L6=zj5=ˆ4=%�3=k�2=��1=��0=B�/=�/=�.=-=�#,=))+=�+*=i+)=I((=0"'=&=�%=��#=��"=�!=ɻ =�=�~=[=�3=�=��=�=�p=a6=/�=	�=�o=�%=��=��=�/=��=cw
=@	=*�=E=�=6e=r�=�u =��< ��<���<��<i��<��<�y�<�M�<v�<���<@��<�_�<}�<���<�p�<h�<J��<tS�<��<e~�<��<ߘ�<� �<���<�%�<o��<t�<֖�<��<���<f�<bb�<�В<�=�<թ�<��<�<��<H�z<�vs<�Il<�e<F�]<��V<��O<{xH<�TA<�4:<�3<��+<��$<��<��<��<�<�<z��;;��;^ �;Mi�;þ;�.�;%��;O=�;0�;�7w;7�\;C�B;M�(;��;�7�:�N�:3̈́:i%:�#�91��n�A�b�nA��=�к����<��.�k�D��V[���q�σ�2����r��������3���08û_YͻxZ׻�;���������$�����h�N��F�����=d����O#��M'�À+��/���3�J�7���;���?�X�C��G��dK�M/O���R�i�V��SZ���]��a��%e���h�3l�0�o��!s�w�v�Z�y��S}�fV�� �������J�� 솼�����'������Z��'���W������q���q6��
Ė�-P���ڙ��d��휼dt������]�����"�����X����������<���������昰�������D������K��O����#������ *���  �  �jN=S�M=��L=\"L=�^K=��J=��I=�I=�JH=�G=ļF=��E=�+E=0bD=��C=!�B=��A= 2A=�c@=ړ?=��>=��==T==�H<=Zr;=��:=��9=��8=O
8=&,7=>L6=xj5=І4=!�3=l�2=��1=��0=E�/=�/=�.=-=�#,=')+=�+*=k+)=D((=5"'=&=�%=��#=��"=�!=ƻ =�=�~=[=�3=�=��=�=�p=a6=.�=�=�o=�%=��=��=�/=��=`w
=>	='�=E=�=0e=w�=�u =��<
��<���<��<b��<��<�y�<�M�<x�<���<J��<�_�<��<���<�p�<}�<=��<tS�<��<`~�<��<㘹< �<���<�%�<f��<x�<Ж�<��<���<_�<fb�<�В<�=�<̩�<��<�<��<M�z<�vs<�Il<�e<B�]<�V<��O<xxH<�TA<�4:<�3<��+<��$<��<��<p�<*�<��<���;_��;7 �;Xi�;�¾;�.�;*��;T=�;��;/8w;��\;�B;y�(;p�;Y8�:�N�:B̈́:�i%:�!�9G����k�b��A����к`���4�Q.���D�tV[�^�q�2σ�=���s��������"���W8û8YͻpZ׻�;����Ϡ��p$�����h�K��N�����;d����c#�yM'���+�
�/���3�M�7���;���?�O�C��G��dK�W/O���R�v�V��SZ���]�1�a��%e�{�h�+3l��o��!s�}�v�g�y��S}�lV��  �������J��솼����'�������Y�����c������n���u6��Ė�)P�� ۙ��d���으mt������c����� ������T����������E���������ߘ��������7������M��I����#������*���  �  �jN=V�M=��L=]"L=�^K=��J=��I=�I=�JH=	�G=üF=��E=�+E=6bD=��C=&�B=��A=(2A=�c@=ѓ?=��>=��==V==�H<=]r;=��:=��9=��8=M
8=0,7==L6={j5=ˆ4=�3=l�2=��1=��0=?�/=�/=�.=-=�#,=%)+=�+*=f+)=H((=5"'=&=�%=��#=��"=�!=̻ =�=�~=[=�3=�=��= �=�p=_6=/�=�=�o=�%=��=��=�/=��=cw
=F	=%�=E=�=2e=t�=�u =��< ��<���<��<t��<��<�y�<�M�<o�<���<F��<�_�<�<���<�p�<k�<N��<nS�<��<]~�<��<䘹<� �<���<�%�<h��<u�<֖�<��<���<d�<]b�<�В<�=�<ک�<��<�<��<7�z<�vs<�Il<�e</�]<�V<��O<~xH<UA<�4:<�3<��+<��$<��<��<~�< �<�<p��;Y��;T �;Ui�; þ;|.�;P��;==�;A�;�7w;��\;I�B;Q�(;��;(8�:>O�:�̄:xi%:�"�9ۨ�����b�]A��"�к����,��.���D��V[�9�q�@σ�����r�����󕮻I���58û9YͻxZ׻�;����נ���$������h�B��G�����,d����F#��M'�ɀ+��/���3�K�7���;���?�e�C��G��dK�L/O���R�~�V��SZ���]�-�a��%e�}�h�.3l�1�o��!s���v�C�y��S}�iV�����������J��솼����'������
Z��$���R������c���x6��Ė�(P���ڙ��d��휼kt������]�����������]����������7���������ܘ�����	���@������V��G����#�������)���  �  �jN=W�M=��L=a"L=�^K=��J=��I=�I=�JH=�G=��F=��E=�+E=5bD=��C=&�B=��A=+2A=�c@=ړ?=��>=��==^==�H<=Zr;=��:=��9=��8=G
8=),7=8L6=}j5=ʆ4=%�3=p�2=��1=��0==�/=�/=�.=-=�#,=#)+=�+*=i+)=K((=/"'=&=�%=��#=��"=�!=̻ =�=�~=[=�3=�=��="�=�p=k6=/�=�=�o=�%=��=��=�/=~�=[w
=>	="�=E=�=;e=p�=�u =$��<���<���<���<h��<מ�<�y�<�M�<s�<���<6��<�_�<|�<���<�p�<h�<T��<bS�<��<T~�<��<ޘ�<� �<���<�%�<~��<p�<���<��<���<k�<ab�<�В<�=�<Ω�<��<�<��<=�z<�vs<vIl<e<:�]<�V<��O<cxH<�TA<~4:<�3<��+<��$<��<��<��<�<(�<���;H��;^ �;:i�;þ;[.�;O��;=�;X�;�7w;��\;��B;$�(;�;D7�:�N�:4̈́:�i%:�#�9f��3�˹b�A��W�к������.��D��V[�O�q�Iσ�@���s�����䕮�.���!8ûkYͻjZ׻�;����u����$������h�D��Q�����)d����=#��M'���+��/���3�<�7���;���?�W�C��G��dK�k/O���R���V��SZ���]��a��%e�x�h�3l�7�o��!s���v�\�y��S}�hV�����������J��)솼�����'�������Y��'���L������b����6��	Ė�.P���ڙ��d��휼Ut������S�����%���z��Y����������C���������ᘰ��������L������Q��L����#������*���  �  �jN=P�M=��L=\"L=�^K=��J=��I=�I=�JH=�G=��F=��E=�+E=5bD=��C=%�B=��A=)2A=�c@=ؓ?=��>=��==X==�H<=[r;=��:=�9=��8=Q
8=+,7=BL6=yj5=ˆ4= �3=k�2=��1=��0=?�/=�/=�.=-=�#,=))+=�+*=k+)=B((=7"'=&=�%=��#=��"=�!=ɻ =�=�~=[=�3=�=��=�=�p=`6=&�=�=�o=�%=��=��=�/=��=dw
=E	=+�=E=�=2e=r�=�u =��<���<���<��<n��<��<�y�<�M�<u�<���<L��<�_�<{�<���<�p�<q�<N��<oS�<��<\~�<��<䘹<� �<���<�%�<`��<h�<ז�<��<���<]�<eb�<�В<�=�<ԩ�<��<�<��<>�z<�vs<�Il<�e<7�]<�V<��O<�xH<�TA<�4:<�3<��+<��$<��<��<��<�<��<���;M��;i �;Xi�;þ;.�;J��;A=�;D�;�7w;d�\;��B;%�(;��;�8�:�N�:/̈́:i%:�!�9�����^�b��A��!�к����E��.���D��V[���q�σ�����r��}�����%���d8û*Yͻ^Z׻�;�(��ޠ���$�����h�9��E�����&d����J#��M'�Ā+�*�/���3�B�7���;���?�S�C���G��dK�F/O���R�f�V��SZ���]�,�a��%e���h�.3l�1�o��!s�i�v�O�y��S}�jV�� �������J��솼����'�������Y�����R������d���y6��Ė�(P���ڙ��d���으st������\�����������U����������=���������嘰�������C������R��N����#�������)���  �  �jN=O�M=��L=Y"L=�^K=��J=��I=�I=�JH=�G=��F=��E=�+E=4bD=��C= �B=��A="2A=�c@=ړ?=��>=��==K==�H<=Xr;=��:=��9=��8=S
8=#,7==L6=oj5=ӆ4=#�3=k�2=��1=��0=J�/=�/=�.=-=�#,=))+=�+*=p+)=>((=9"'=&=�%=��#=��"=�!=û =�=�~=[=�3=�=��=�=�p=d6=6�=�=�o=�%=��=��=�/=��=_w
==	=&�=E= �=1e=w�=�u =��<��<���<
��<]��<��<�y�<�M�<w�<���<O��<�_�<��<���<�p�<r�<>��<mS�<��<b~�<��<ܘ�<� �<���<�%�<h��<��<ϖ�<��<���<U�<rb�<�В<�=�<ɩ�<��<�~�<��<e�z<�vs<�Il<�e<W�]<�V<}�O<uxH<�TA<�4:<�3<��+<��$<��<��<e�<O�<�<���;C��;< �;Ci�;þ;�.�;"��;:=�;�;�7w;��\;h�B;�(;��;�8�:�N�:5̈́:j%:� �9j������b��B��3�к)���A�9.���D�&V[���q�Iσ�8���s��~����������8ûYͻ�Z׻�;ụ�� ��z$�����h�S��F�����Ad����i#��M'���+��/���3�s�7���;���?�D�C���G��dK�Y/O���R�y�V��SZ���]�0�a��%e�}�h�&3l��o�"s�{�v�p�y��S}�mV�����������J��솼���y'�������Y�����c������q���s6��Ė�1P���ڙ��d���으lt������d���!��������H����������H�������������������.������B��F����#������*���  �  �jN=P�M=��L=\"L=�^K=��J=��I=�I=�JH=�G=��F=��E=�+E=5bD=��C=%�B=��A=)2A=�c@=ؓ?=��>=��==X==�H<=[r;=��:=�9=��8=Q
8=+,7=BL6=yj5=ˆ4= �3=k�2=��1=��0=?�/=�/=�.=-=�#,=))+=�+*=k+)=B((=7"'=&=�%=��#=��"=�!=ɻ =�=�~=[=�3=�=��=�=�p=`6=&�=�=�o=�%=��=��=�/=��=dw
=E	=+�=E=�=2e=r�=�u =��<���<���<��<n��<��<�y�<�M�<u�<���<L��<�_�<{�<���<�p�<q�<N��<oS�<��<\~�<��<䘹<� �<���<�%�<`��<h�<ז�<��<���<]�<eb�<�В<�=�<ԩ�<��<�<��<>�z<�vs<�Il<�e<7�]<�V<��O<�xH<�TA<�4:<�3<��+<��$<��<��<��<�<��<���;M��;i �;Xi�;þ;.�;J��;A=�;D�;�7w;d�\;��B;%�(;��;�8�:�N�:/̈́:i%:�!�9�����^�b��A��!�к����E��.���D��V[���q�σ�����r��}�����%���d8û*Yͻ^Z׻�;�(��ޠ���$�����h�9��E�����&d����J#��M'�Ā+�*�/���3�B�7���;���?�S�C���G��dK�F/O���R�f�V��SZ���]�,�a��%e���h�.3l�1�o��!s�i�v�O�y��S}�jV�� �������J��솼����'�������Y�����R������d���y6��Ė�(P���ڙ��d���으st������\�����������U����������=���������嘰�������C������R��N����#�������)���  �  �jN=W�M=��L=a"L=�^K=��J=��I=�I=�JH=�G=��F=��E=�+E=5bD=��C=&�B=��A=+2A=�c@=ړ?=��>=��==^==�H<=Zr;=��:=��9=��8=G
8=),7=8L6=}j5=ʆ4=%�3=p�2=��1=��0==�/=�/=�.=-=�#,=#)+=�+*=i+)=K((=/"'=&=�%=��#=��"=�!=̻ =�=�~=[=�3=�=��="�=�p=k6=/�=�=�o=�%=��=��=�/=~�=[w
=>	="�=E=�=;e=p�=�u =$��<���<���<���<h��<מ�<�y�<�M�<s�<���<6��<�_�<|�<���<�p�<h�<T��<bS�<��<T~�<��<ޘ�<� �<���<�%�<~��<p�<���<��<���<k�<ab�<�В<�=�<Ω�<��<�<��<=�z<�vs<vIl<e<:�]<�V<��O<cxH<�TA<~4:<�3<��+<��$<��<��<��<�<(�<���;H��;^ �;:i�;þ;[.�;O��;=�;W�;�7w;��\;��B;$�(;�;D7�:�N�:3̈́:�i%:�#�9j��4�̹b�A��X�к������.��D��V[�O�q�Iσ�@���s�����䕮�.���!8ûkYͻjZ׻�;����u����$������h�D��Q�����)d����=#��M'���+��/���3�<�7���;���?�W�C��G��dK�k/O���R���V��SZ���]��a��%e�x�h�3l�7�o��!s���v�\�y��S}�hV�����������J��)솼�����'�������Y��'���L������b����6��	Ė�.P���ڙ��d��휼Ut������S�����%���z��Y����������C���������ᘰ��������L������Q��L����#������*���  �  �jN=V�M=��L=]"L=�^K=��J=��I=�I=�JH=	�G=üF=��E=�+E=6bD=��C=&�B=��A=(2A=�c@=ѓ?=��>=��==V==�H<=]r;=��:=��9=��8=M
8=0,7==L6={j5=ˆ4=�3=l�2=��1=��0=?�/=�/=�.=-=�#,=%)+=�+*=f+)=H((=5"'=&=�%=��#=��"=�!=̻ =�=�~=[=�3=�=��= �=�p=_6=/�=�=�o=�%=��=��=�/=��=cw
=F	=%�=E=�=2e=t�=�u =��< ��<���<��<u��<��<�y�<�M�<o�<���<F��<�_�<��<���<�p�<k�<N��<nS�<��<]~�<��<䘹<� �<���<�%�<h��<u�<֖�<��<���<d�<]b�<�В<�=�<ک�<��<�<��<7�z<�vs<�Il<�e</�]<�V<��O<~xH<UA<�4:<�3<��+<��$<��<��<~�< �<�<p��;Y��;T �;Ui�; þ;|.�;P��;==�;A�;�7w;��\;I�B;P�(;��;'8�:=O�:�̄:wi%:�"�9������b�^A��#�к����,��.���D��V[�9�q�Aσ�����r�����󕮻I���58û9YͻxZ׻�;����ؠ���$������h�B��G�����,d����F#��M'�ɀ+��/���3�K�7���;���?�e�C��G��dK�L/O���R�~�V��SZ���]�-�a��%e�}�h�.3l�1�o��!s���v�C�y��S}�iV�����������J��솼����'������
Z��$���R������c���x6��Ė�(P���ڙ��d��휼kt������]�����������]����������7���������ܘ�����	���@������V��G����#�������)���  �  �jN=S�M=��L=\"L=�^K=��J=��I=�I=�JH=�G=ļF=��E=�+E=0bD=��C=!�B=��A= 2A=�c@=ړ?=��>=��==T==�H<=Zr;=��:=��9=��8=O
8=&,7=>L6=xj5=І4=!�3=l�2=��1=��0=E�/=�/=�.=-=�#,=')+=�+*=k+)=D((=5"'=&=�%=��#=��"=�!=ƻ =�=�~=[=�3=�=��=�=�p=a6=.�=�=�o=�%=��=��=�/=��=`w
=>	='�=E=�=0e=w�=�u =��<
��<���<	��<c��<��<�y�<�M�<x�<���<J��<�_�<��<���<�p�<}�<=��<tS�<��<`~�<��<㘹< �<���<�%�<f��<x�<Ж�<��<���<_�<fb�<�В<�=�<̩�<��<�<��<M�z<�vs<�Il<�e<B�]<�V<��O<xxH<�TA<�4:<�3<��+<��$<��<��<p�<*�<��<���;_��;7 �;Xi�;�¾;�.�;*��;T=�;��;/8w;��\;
�B;x�(;p�;X8�:�N�:Ä́:�i%:�!�9N����l�b��A����кa���4�R.���D�tV[�_�q�2σ�=���s��������"���W8û8YͻpZ׻�;����Ϡ��p$�����h�K��N�����;d����c#�yM'���+�
�/���3�M�7���;���?�O�C��G��dK�W/O���R�v�V��SZ���]�1�a��%e�{�h�+3l��o��!s�}�v�g�y��S}�lV��  �������J��솼����'�������Y�����c������n���u6��Ė�)P�� ۙ��d���으mt������c����� ������T����������E���������ߘ��������7������M��I����#������*���  �  �jN=T�M=��L=_"L=�^K=��J=��I=�I=�JH=�G=��F=��E=�+E=2bD=��C=!�B=��A=&2A=�c@=Փ?=��>=��==Z==�H<=Yr;=��:=�9=��8=O
8=(,7=>L6=zj5=ˆ4=%�3=k�2=��1=��0=B�/=�/=�.=-=�#,=))+=�+*=i+)=I((=0"'=&=�%=��#=��"=�!=ɻ =�=�~=[=�3=�=��=�=�p=a6=/�=	�=�o=�%=��=��=�/=��=cw
=@	=*�=E=�=6e=r�=�u =��< ��<���<��<i��<��<�y�<�M�<v�<���<@��<�_�<}�<���<�p�<h�<J��<tS�<��<e~�<��<ߘ�<� �<���<�%�<o��<t�<֖�<��<���<f�<bb�<�В<�=�<թ�<��<�<��<H�z<�vs<�Il<�e<F�]<��V<��O<{xH<�TA<�4:<�3<��+<��$<��<��<��<�<�<z��;;��;^ �;Mi�;þ;�.�;%��;O=�;0�;�7w;7�\;C�B;M�(;��;�7�:�N�:3̈́:	i%:�#�99��o�C�b�oA��>�к ���<��.�l�D��V[���q�σ�2����r��������3���08û_YͻxZ׻�;���������$�����h�N��F�����=d����O#��M'�À+��/���3�J�7���;���?�X�C��G��dK�M/O���R�i�V��SZ���]��a��%e���h�3l�0�o��!s�w�v�Z�y��S}�fV�� �������J�� 솼�����'������Z��'���W������q���q6��
Ė�-P���ڙ��d��휼dt������]�����"�����X����������<���������昰�������D������K��O����#������ *���  �  �jN=V�M=��L=a"L=�^K=��J=��I=�I=�JH=	�G=ƼF=��E=�+E=3bD=��C=$�B=��A=,2A=�c@=ԓ?=��>=��==Z==�H<=`r;=��:=��9=��8=J
8=+,7=;L6=�j5=͆4="�3=m�2=��1=��0=@�/=�/=�.=-=�#,=#)+=�+*=f+)=M((=1"'=&=�%=��#=��"=�!=л =�=�~=[=�3=�=��=$�=�p=c6=0�=�=�o=�%=��=��=�/=�=cw
=B	='�=E=�=3e=s�=�u =��<��<���<��<m��<���<�y�<�M�<q�<���<>��<�_�<v�<���<�p�<p�<W��<iS�<
��<Y~�<��<ܘ�<� �<���<�%�<q��<i�<ږ�<��<���<l�<ab�<�В<�=�<֩�<��<�<��<<�z<�vs<�Il<�e<5�]<�V<��O<nxH<UA<{4:<�3<��+<��$<��<��<��<�<�<m��;s��;m �;3i�;
þ;e.�;<��; =�;Z�;�7w;!�\;f�B;��(;��;�7�:�O�:2̈́:�i%:?#�9d����6�b��@���кd���%��.���D��V[� �q�-σ�0����r�����핮�G���8ûYYͻkZ׻�;���껸����$������h�M��L�����<d����4#��M'���+��/���3�D�7���;���?�f�C��G��dK�K/O���R�x�V��SZ���]�)�a��%e�{�h�'3l�+�o��!s���v�R�y��S}�hV�����������J��!솼 ����'������Z�� ���J������k���}6��Ė�0P���ڙ��d��	휼ct������Y��������y��Z����������:���������ؘ��������A������S��C����#�������)���  �  �jN=U�M=��L=\"L=�^K=��J=��I=�I=�JH=�G=üF=��E=�+E=4bD=��C='�B=��A=$2A=�c@=֓?=��>=��==V==�H<=]r;=��:=��9=��8=N
8=*,7=<L6=xj5=Ά4="�3=l�2=��1=��0=E�/=�/=�.=-=�#,=%)+=�+*=g+)=G((=4"'=&=�%=��#=��"=�!=Ȼ =�=�~=[=�3=�=��=�=�p=a6=0�=�=�o=�%=��=��=�/=~�=bw
=@	=$�=E=�=2e=w�=�u =��<��<���<��<l��<��<�y�<�M�<n�<���<C��<�_�<��<���<�p�<t�<F��<mS�<��<U~�<��<䘹< �<���<�%�<l��<t�<ږ�<��<���<_�<cb�<�В<�=�<ҩ�<��<�<��<R�z<�vs<�Il<�e<G�]<�V<��O<vxH<�TA<�4:<�3<��+<��$<��<��<��< �<�<���;X��;? �;Vi�;þ;Z.�;T��;5=�;�;�7w;A�\;X�B;l�(;��;�7�:&O�:�̄:�i%:�!�9Ч���ܸb��A���к[���;�B.���D�vV[�j�q�Hσ�3����r�����핮�?���D8û?Yͻ~Z׻�;����à���$�����h�D��V�����1d����U#��M'���+��/���3�J�7���;���?�`�C��G��dK�Q/O���R���V��SZ���]�,�a��%e�{�h�(3l�"�o��!s���v�U�y��S}�nV�����������J��솼����'������Z�����[������d����6��	Ė�(P�� ۙ��d��휼ht������Y�����������W����������?�������������������3������K��H����#������*���  �  �jN=O�M=��L=\"L=�^K=��J=��I=�I=�JH=�G=��F=��E=�+E=2bD=��C= �B=��A='2A=�c@=ԓ?=��>=��==W==�H<=Yr;=��:=��9=��8=P
8=&,7=FL6=zj5=ˆ4=$�3=i�2=��1=��0=E�/=�/=�.=-=�#,=))+=�+*=l+)=D((=6"'=&=�%=��#=��"=�!=Ȼ =�=�~=[=�3=�=��=�=�p=^6=.�=�=�o=�%=��=��=�/=��=`w
=B	=/�=E=�=3e=v�=�u =��<��<���<��<f��<��<�y�<�M�<w�<���<G��<�_�<��<���<�p�<l�<L��<rS�<��<a~�<��<ޘ�<� �<���<�%�<g��<t�<Ԗ�<��<���<_�<kb�<�В<�=�<ʩ�<��<�<��<T�z<�vs<�Il<�e<J�]<��V<��O<�xH<�TA<�4:<�3<��+<��$<��<��<~�<�<��<���;;��;\ �;Ei�;þ;�.�;��;D=�;6�;�7w;$�\;�B;h�(;��;8�:�N�:̈́:�i%:!�9����z�b��A��*�к���`�g.���D�wV[�Úq��΃����s�����������U8û3Yͻ~Z׻�;��������$��	���h�S��H�����Bd����Q#��M'�΀+��/���3�M�7���;���?�K�C���G��dK�W/O���R�W�V��SZ���]�*�a��%e���h�$3l�%�o��!s�]�v�a�y��S}�lV�����������J��솼����'������Z��#���U������q���t6��
Ė�.P���ڙ��d��휼mt������_�����������P����������G���������혰�������9������I��S����#������	*���  �  �jN=R�M=��L=^"L=�^K=��J=��I=�I=�JH=�G=��F=��E=�+E=3bD=��C="�B=��A=)2A=�c@=ٓ?=��>=��==Z==�H<=\r;=��:=��9=��8=O
8=',7=:L6=|j5=͆4=%�3=n�2=��1=��0=C�/=�/=�.= -=�#,=')+=�+*=k+)=I((=1"'=&=�%=��#=��"=�!=˻ =�=�~=[=�3=�=��= �=�p=f6=0�=�=�o=�%=��=��=�/=��=aw
=?	=%�=E=�=7e=u�=�u =��<��<���<��<e��<��<�y�<�M�<w�<���<>��<�_�<|�<���<�p�<i�<P��<fS�<��<Y~�<��<ؘ�<� �<���<�%�<z��<q�<ٖ�<��<���<g�<hb�<�В<�=�<ҩ�<��<	�<��<K�z<�vs<�Il<�e<F�]<
�V<��O<nxH<�TA<�4:<�3<��+<��$<��<��<��<�<�<���;K��;[ �;"i�;þ;e.�;2��;=�;B�;�7w;m�\;v�B;+�(;��;7�:O�:;̈́:Ni%:p"�9&����a�b�;A���к����{.�_�D��V[�I�q�?σ�E����r��������#���/8û\YͻvZ׻�;���껚����$������h�R��L�����>d����H#��M'���+��/���3�H�7���;���?�Q�C��G��dK�S/O���R��V��SZ���]��a��%e�w�h�3l�"�o��!s���v�c�y��S}�iV��  �������J��"솼����'�������Y��&���Q������m���}6��	Ė�5P���ڙ��d��휼Zt������Z�����#���~��R����������?���������ޘ��������<������K��J����#������*���  �  �jN=Y�M=��L=["L=�^K=��J=��I=�I=�JH=�G=ļF=��E=�+E=:bD=��C=,�B=��A='2A=�c@=ғ?=��>=��==[==�H<=_r;=��:=��9=��8=M
8=2,7=<L6=zj5=ˆ4="�3=l�2=��1=��0==�/=�/=�.=-=�#,=&)+=�+*=c+)=I((=3"'=&=�%=��#=��"=�!=ͻ =�=�~=[=�3=�=��=!�=�p=`6=(�=
�=�o=�%=��=��=�/=��=cw
=J	=$�=E=�=8e=q�=�u =��<���<���<��<~��<��<�y�<�M�<l�<���<C��<�_�<x�<���<�p�<i�<L��<eS�<��<P~�<��<☹<~ �<���<�%�<l��<f�<ܖ�<��<���<`�<[b�<�В<�=�<ߩ�<��<�<��<8�z<�vs<�Il<�e<8�]<�V<��O<�xH<UA<�4:<�3<��+<��$<��<��<��<�<�<V��;b��;H �;?i�;Aþ;;.�;���;=�;1�;�7w;��\;�B;�(;��;�7�:mO�:�̄:i%:c$�9�����͸b�uA��6�кR���5��.�T�D� W[��q�Fσ�ﰎ��r�����ҕ��b���58ûIYͻpZ׻�;�$��͠���$������h�3��L�����d����C#��M'�Ȁ+�#�/���3�C�7���;���?�p�C�ޏG��dK�M/O���R���V��SZ���]��a��%e���h�!3l�6�o��!s���v�1�y��S}�dV�����������J��솼�����'������Z��&���U������W����6�� Ė�*P�� ۙ��d��휼gt������W�����������`����������1���������٘��������C������R��F����#�������)���  �  �jN=T�M=��L=_"L=�^K=��J=��I=�I=�JH=�G=üF=��E=�+E=1bD=��C=!�B=��A=$2A=�c@=ړ?=��>=��==T==�H<=Xr;=��:=��9=��8=H
8=#,7=AL6=yj5=І4=&�3=o�2=��1=��0=C�/=�/=�.=-=�#,=%)+=�+*=n+)=E((=4"'=&=�%=��#=��"=�!=ǻ =�=�~=[=�3=�=��=�=�p=e6=2�=�=�o=�%=��=��=�/=��=Yw
=A	=(�=E=�=8e=u�=�u =$��<��<���<��<b��<מ�<�y�<�M�<|�<���<F��<�_�<��<���<�p�<u�<F��<iS�<��<V~�<��<ژ�<� �<���<�%�<p��<y�<Җ�<��<���<b�<nb�<�В<�=�<©�<��<�<��<M�z<�vs<�Il<�e<H�]<�V<��O<�xH<�TA<�4:<�3<��+<��$<��<��<t�<%�<�<���;X��;G �;1i�;�¾;\.�;(��;$=�;�;�7w;{�\;J�B;s�(;w�;�7�:�N�:~̈́:Cj%:�"�9/����÷b��A����к�����.�a�D��V[�J�q�%σ�"���@s������������T8ûAYͻ�Z׻�;���껭����$�����h�T��R�����?d����W#��M'���+���/���3�T�7���;���?�H�C��G��dK�u/O���R�r�V��SZ���]��a��%e�u�h�3l��o��!s�r�v�j�y��S}�hV�����������J��솼����'�������Y�����Z������m���6��Ė�2P���ڙ��d���으ct������a�����������L����������O���������ܘ��������:������J��F����#������*���  �  �lN=��M=K�L=r%L=#bK=[�J=�I=I=�OH=Z�G=o�F=��E=^2E=iD=��C=��B=�B=�:A=�l@=g�?=��>=S�==a(==T<=h~;=J�:=��9=d�8=�8=�:7=�[6=mz5=_�4=H�3=3�2=��1=��0=�0=�/=x&.=�1-=:,=�?+=C*=�C)=�@(=�;'=3&=t'%=�$=�#=X�!=�� =k�=��=Xy=`R=�'=I�=��=�=�V=�=��=�=G=�=�=�P=��=��
=M6	=��=�e=j�=/�==� =�.�<�+�<!�<|�<���<���<=��<���<SO�<?�<(��<��<.C�<���<���<?�<6��<�x�<l�<��<d-�<䶹<�<�<��<%>�<��<P3�<ީ�<�<<���<n�<�ڒ<�E�<���<$�<y��<c�<ءz<�ps<�?l<�e<4�]<p�V<N�O<�\H<�5A<c:<��2<*�+<ʻ$<$�<��<��<��<��<�6�;8Y�;@��;C��; �;̄�;���;��;[$�;o�u;A[;"�@;��&;,	;t��:E��:��:��:�Qi9�,!�R
�>�j�$d���Ժ2���5�B;0�9G��]�!�s�S넻�͏�����a2������9���TĻqtλ!tػ�S���i���K5���K��������z����;���#���'�u�+�K0��04�i;8�a:<��-@��D���G���K�ȌO�wJS���V�B�Z��J^�{�a��se���h��{l�C�o��es���v� 3z�4�}��s��	�������d���������0>���׋��n���������(��d����F��<Ӗ��^��~虼Oq���������/���������B������������񘪼���������y������S�������������⟹��!��ʣ���&���  �  �lN=��M=L�L=s%L=$bK=U�J=��I=I=�OH=Y�G=o�F=��E=Z2E=iD=��C=��B=�B=�:A=�l@=g�?=��>=O�==\(==T<=k~;=K�:=��9=o�8=�8=�:7=�[6=sz5=`�4=Q�3=5�2=��1=��0=�0=�/=w&.=�1-=:,=�?+=(C*=�C)=�@(=�;'=	3&=r'%=�$=�#=S�!=�� =c�=��=Yy=aR=�'=A�=��=��=�V=�=��=�=G=�=�=�P=��=��
=H6	=��=�e=n�=8�==� =�.�<�+�<,!�<r�<���<���<T��<��<SO�<G�<��<���<(C�<���<���<?�<7��<�x�<s�<���<c-�<߶�<�<�<	��<!>�<$��<M3�<ש�<��<폝<���<n�<�ڒ<�E�<ꯋ<�<z��<h�<�z<�ps<�?l<�e<O�]<t�V<U�O<�\H<g5A<l:<��2</�+<һ$<(�<��<��<��< �<�6�;9Y�;1��;#��; �;���;���;慕;U$�;�u;�@[;��@;`�&;�;���:���:��:��:�]i9�-!��
��j��c����Ժ����5��;0��G�ˈ]���s�[넻$Ώ�����;2������O���TĻ�tλTtػ T⻿�:���s5���K��������z����+;���#���'�c�+�20��04��;8�v:<��-@��D���G���K�ԌO��JS���V��Z��J^�V�a��se���h��{l�<�o�xes���v�33z�<�}�us���������}d���������6>��w׋��n���������(��]����F��=Ӗ��^���虼Kq���������1���������D������������옪����������t������C������������������!��ڣ���&���  �  �lN=��M=D�L=s%L=%bK=X�J=�I=I=�OH=S�G=r�F=��E=]2E=iD=�C=��B=�B=�:A=�l@=c�?=��>=M�==f(==T<=m~;=E�:=��9=i�8=�8=�:7=�[6=wz5=W�4=N�3=7�2=��1=��0=�0=�/=v&.=�1-=:,=�?+=$C*=yC)=A(=�;'=3&=w'%=�$=�#=O�!=�� =a�=��=Wy=^R=�'=>�=�=ߐ=�V=�=��=�=G=�=�=�P=��=��
=M6	=��=�e=c�=8�==� =�.�<�+�</!�<p�<���<���<E��<��<CO�<M�<��<��<'C�<���<���<?�<F��<�x�<�<���<g-�<趹<�<�<��<>�<'��<J3�<橤<�<���<���<�m�<�ڒ<�E�<���<�<��<a�<Сz<�ps<�?l<�e<8�]<\�V<c�O<�\H<5A<_:<��2<�+<ϻ$<-�<��<ʐ<��<%�<c6�;JY�;G��;;��;- �;���;���;煕;�$�;2�u;�@[;��@;E�&;x	;��:��:��:$�:�Vi9�.!��
���j��b���Ժ����5��;0��G�|�]���s�d넻�͏�~���n2����������TĻ�tλtػ�S���.����5���K����р�	��z����6;���#���'�^�+�60�}04�c;8�r:<��-@��D���G���K���O�xJS���V�#�Z��J^�X�a��se���h��{l�_�o�pes���v�3z�=�}��s���������vd���������7>��x׋��n���������(��Q����F��9Ӗ��^���虼Bq���������5������A�������������������������|������B�������������쟹��!��գ���&���  �  �lN=��M=P�L=u%L=#bK=S�J=��I=I=�OH=X�G=p�F=��E=^2E=iD=��C=��B=�B=�:A=�l@=i�?=��>=P�==_(==T<=k~;=J�:=��9=g�8=�8=�:7=�[6=tz5=^�4=N�3=3�2= �1=��0=�0=�/=x&.=�1-=:,=�?+=$C*=�C)=�@(=�;'=
3&=r'%=�$=�#=S�!=�� =a�=��=Wy=_R=�'=?�=��=�=�V=�=��=
�=G=�=�=�P=��=��
=H6	=��=�e=l�=3�==� =�.�<�+�<*!�<r�<���<���<C��<��<PO�<F�<��<��<)C�<���<��<?�<6��<�x�<v�<���<d-�<綹<�<�<	��<>�<!��<P3�<ש�<��<菝<���<n�<�ڒ<�E�<���<�<��<i�<ߡz<�ps<�?l<�e<B�]<r�V<^�O<�\H<u5A<i:<��2<?�+<׻$<%�<��<��<��<�<�6�;9Y�;'��;@��; �;���;���;���;X$�;=�u;-A[;��@;j�&;	;9��:���:��:�:SUi9/-!�7
���j�\c��6�Ժ����5�%;0�G��]���s�S넻*Ώ�|���i2������?���TĻ�tλJtػ�S���+���t5���K����݀�	��z����0;���#���'�X�+�?0��04�};8��:<��-@��D���G���K���O��JS���V�'�Z��J^�k�a��se���h��{l�@�o�{es���v�13z�7�}��s���������|d���������5>��~׋��n���������(��Z����F��<Ӗ��^���虼Kq���������/���������H����������������������s������O�������������៹��!��ۣ���&���  �  �lN=��M=K�L=n%L=*bK=\�J=��I=I=�OH=[�G=q�F=��E=`2E=iD=��C=��B=�B=�:A=�l@=i�?=��>=T�==](==T<=o~;=E�:=��9=g�8=�8=�:7=�[6=nz5=]�4=O�3=1�2= �1=��0=�0=�/=~&.=�1-=:,=�?+=!C*=�C)=�@(=�;'=3&=v'%=�$=�#=W�!=�� =h�=��=Xy=aR=�'=G�=��=�=�V=�=��=�=G=�=
�=�P=��=��
=F6	=�=�e=o�=/�==� =�.�<�+�<!�<~�<���<���<E��<��<HO�<J�<)��< ��<0C�<���<��<?�<1��<�x�<m�<��<^-�<趹<�<�<	��<&>�<��<S3�<۩�<�<���<���<n�<�ڒ<�E�<<�<���<\�<�z<�ps<�?l<}e<P�]<^�V<X�O<�\H<e5A<|:<��2<+�+<��$<@�<��<��<��<�<�6�;BY�;9��;O��;��;Ą�;���;!��;M$�;I�u;/A[;\�@;��&;�;���:A��:��:��:�Ui9F(!�%	
���j�d��\�Ժ����5�&;0�PG���]�@�s�$넻9Ώ�����F2������g���TĻZtλ+tػ�S���Q���O5���K���������z����;���#���'�i�+�?0�y04�u;8�Z:<��-@��D���G���K���O��JS���V�F�Z��J^�y�a��se���h��{l�@�o��es���v�<3z�(�}��s���������yd���������/>���׋��n�����!����(��b����F��BӖ��^���虼Jq���������+���������8������
������昪�����������������U�������������럹��!��ף���&���  �  �lN=��M=N�L=s%L="bK=T�J=�I=I=�OH=X�G=q�F=��E=]2E=iD=��C=��B=�B=�:A=�l@=g�?=��>=P�==c(==T<=i~;=I�:=��9=g�8=�8=�:7=�[6=tz5=[�4=P�3=3�2=��1=��0=�0=�/=}&.=�1-=:,=�?+=&C*=�C)= A(=�;'=
3&=w'%=�$=�#=V�!=�� =a�=��=Yy=bR=�'=?�=��=�=�V=�=��=�=G=�=�=�P=��=��
=H6	=��=�e=k�=4�==� =�.�<�+�<(!�<u�<���<���<B��<��<MO�<D�<��<��<)C�<���<��<?�<5��<�x�<u�<��<d-�<涹<�<�<	��<!>�<$��<L3�<㩤<��<ꏝ<���<n�<�ڒ<�E�<���<�<���<Z�<�z<�ps<�?l<�e<I�]<W�V<g�O<�\H<|5A<`:<��2<7�+<ѻ$<�<��<<��<�<�6�;FY�;.��;:��; �;���;���;���;^$�;f�u;A[;��@;p�&;H	;���:r��:g�:5�:TUi9�+!��
���j�Gc����Ժ����5��;0�G���]�7�s�*넻%Ώ�y���u2������^���TĻ�tλKtػ�S���.���V5���K����؀���z����/;���#���'�_�+�>0�|04�z;8�~:<��-@��D���G���K���O��JS���V�<�Z��J^�g�a��se���h��{l�L�o�}es���v�03z�1�}��s���������d���������5>��|׋��n���������(��[����F��=Ӗ��^���虼Jq���������2��򉡼���G��������������������������������M���������������!��֣���&���  �  �lN=��M=H�L=q%L=#bK=U�J=�I=I=�OH=Q�G=r�F=��E=^2E=iD=�C=��B=�B=�:A=�l@=c�?=��>=K�==f(==T<=j~;=F�:=��9=i�8=�8=�:7=�[6=tz5=Y�4=P�3=4�2=��1=��0=�0=�/=x&.=�1-=:,=�?+=)C*=|C)= A(=�;'=3&=t'%=�$=�#=N�!=�� =`�=��=Xy=`R=�'=?�=�=ސ=�V=�=��=�=G=�=�=�P=��=��
=G6	=��=�e=h�=9�==� =�.�<�+�<+!�<i�<���<���<D��<��<FO�<G�<��<��<C�<���<���<?�<;��<�x�<��<���<i-�<궹<�<�<��<>�<.��<G3�<੤<��<ꏝ<���<n�<�ڒ<�E�< ��<�<}��<a�<ڡz<�ps<�?l<�e<@�]<a�V<\�O<{\H<�5A<O:<��2<"�+<ɻ$<%�<��<Đ<��<3�<Y6�;KY�;3��;B��;: �;���;���;���;j$�;:�u;�@[; A;�&;�	;q��:���:�:?�:+Wi9
0!��
���j�Pc����Ժ����5��;0��G�&�]���s�Q넻5Ώ�l����2��u�������TĻ�tλtػ�S���'����5���K����Ȁ���z����1;���#���'�`�+�;0��04�c;8��:<��-@��D���G���K���O��JS���V�/�Z��J^�S�a��se���h��{l�V�o�xes���v�%3z�?�}��s���������|d���������?>��t׋��n���������(��N����F��7Ӗ��^���虼Dq������{��8���������G�������������������������{������D�������������ꟹ��!��䣼��&���  �  �lN=��M=G�L=p%L=%bK=Z�J=��I=I=�OH=Y�G=t�F=��E=`2E=iD=��C=��B=�B=�:A=�l@=h�?=��>=N�==a(==T<=m~;=F�:=��9=k�8=�8=�:7=�[6=pz5=Z�4=M�3=2�2=��1=��0=�0=�/=|&.=�1-=:,=�?+=$C*=~C)=�@(=�;'=3&=t'%=�$=�#=T�!=�� =c�=��=Xy=`R=�'=A�=��=�=�V=�=��=�=G=�=�=�P=��=��
=G6	=��=�e=h�=2�==� =�.�<�+�<!!�<y�<���<���<I��< ��<HO�<I�<��<	��<&C�<���<��<?�<3��<�x�<w�<���<e-�<붹<�<�<��<>�<%��<P3�<۩�<�<<���<n�<�ڒ<�E�<���<�<���<^�<ۡz<�ps<�?l<�e<?�]<]�V<]�O<�\H<v5A<^:<��2<�+<û$<,�<��<��<��<!�<�6�;aY�;(��;P��;( �;���;���;��;J$�;�u;!A[;��@;W�&;3	;(��: ��:#�:D�:*Yi9�-!��
� �j��c����Ժ����5�F;0�G�0�]�0�s�0넻'Ώ�����j2������z���TĻ�tλtػ�S���3���f5���K����Ѐ���z����';���#���'�_�+�30��04�e;8�r:<��-@��D���G���K�ČO��JS���V�D�Z��J^�m�a��se���h��{l�Q�o��es���v�-3z�<�}��s���������yd���������8>��x׋��n���������(��Y����F��;Ӗ��^���虼Aq���������/���������B������������󘪼���������~������N�������������쟹��!��٣���&���  �  �lN=��M=O�L=x%L= bK=W�J=��I=I=�OH=Y�G=p�F=��E=a2E=iD=��C=��B=�B=�:A=�l@=g�?=��>=V�==](==T<=f~;=N�:=��9=h�8=�8=�:7=�[6=oz5=^�4=M�3=0�2=��1=��0=�0=�/=z&.=�1-=:,=�?+="C*=�C)= A(=�;'=3&=u'%=�$=�#=Y�!=�� =g�=��=Xy=bR=�'=F�=��=�=�V=�=��=
�=G=�=�=�P=��=��
=E6	=��=�e=p�=/�==� =�.�<�+�<!�<{�<���<���<F��<��<WO�<=�<��<���<3C�<���<���<?�<2��<�x�<m�<��<`-�<붹<�<�<��<#>�<��<Y3�<ک�<��<珝<���<n�<�ڒ<�E�<鯋<�<��<[�<�z<�ps<�?l<{e<K�]<^�V<Y�O<�\H<]5A<n:<��2<=�+<�$<�<��<��<̍<	�<�6�;;Y�;7��;\��; �;΄�;���;(��;Q$�;u�u;A[;��@;��&;�;���:&��:�:�:QVi9�*!��	
���j��c��-�Ժ����5�0;0�KG���]�P�s�>넻*Ώ�����U2������0���TĻ�tλAtػ�S⻸�F���B5���K����߀���z����;���#���'�g�+�50�x04�};8�|:<��-@��D���G���K�ȌO��JS���V�J�Z��J^�x�a��se���h��{l�:�o��es���v�A3z�4�}��s����������d���������*>��~׋��n���������(��c����F��@Ӗ��^���虼Mq���������&���������I������ ������옪�����������������X�������������럹��!��ң���&���  �  �lN=��M=F�L=r%L='bK=\�J=��I=I=�OH=W�G=r�F=��E=^2E=iD=��C=��B=�B=�:A=�l@=f�?=��>=Q�==_(==T<=l~;=E�:=��9=e�8=�8=�:7=�[6=pz5=Y�4=N�3=2�2=��1=��0=�0=�/=y&.=�1-=:,=�?+=!C*={C)=�@(=�;'=3&=t'%=�$=�#=R�!=�� =f�=��=[y=cR=�'=C�=�=��=�V=�=��=�=G=�=�=�P=��=��
=I6	=��=�e=h�=2�==� =�.�<�+�<#!�<q�<���<���<>��<��<DO�<G�<&��<��<*C�<���< ��<?�<B��<�x�<s�<��<d-�<涹<�<�<��<>�<$��<O3�<۩�<�<�<���< n�<�ڒ<�E�<�<�<}��<\�<ܡz<�ps<�?l<�e<A�]<Z�V<U�O<�\H<n5A<d:<��2<�+<ʻ$<3�<��<��<��<�<�6�;OY�;W��;B��; �;ӄ�;���;��;�$�;K�u;A[;��@;��&;	;���:ݮ�:��:T�:�Si9,!�B
���j��c����Ժ����5�z;0�G��]��s�I넻Ώ�����k2����������TĻytλ#tػ�S���5���y5���K����܀����z����;���#���'�`�+�90��04�n;8�g:<��-@��D���G���K�ǌO��JS���V�=�Z��J^�m�a��se���h��{l�T�o��es���v�.3z�6�}��s���������|d���������4>��y׋��n���������(��\����F��;Ӗ��^��~虼Dq���������0���������?������������򘪼���������������O�������������ퟹ��!��أ���&���  �  �lN=��M=K�L=s%L=$bK=Q�J= �I=I=�OH=Y�G=t�F=��E=\2E=iD=�C=��B=�B=�:A=�l@=l�?=��>=O�==b(==T<=n~;=I�:=��9=l�8=�8=�:7=�[6=uz5=[�4=O�3=3�2=��1=��0=�0=�/=w&.=�1-=:,=�?+=(C*=�C)=A(=�;'=
3&=u'%=�$=�#=Q�!=�� =]�=��=Zy=`R=�'=:�=�=ߐ=�V=�=��=
�=G=�=�=�P=��=��
=G6	=��=�e=f�=6�==� =�.�<�+�</!�<i�<���<���<H��<��<MO�<N�<��<��<(C�<���<��<?�<@��<�x�<��<���<n-�<涹<�<�<��<>�<,��<K3�<ީ�<��<ꏝ<���<n�<�ڒ<�E�<���<�<|��<i�<֡z<�ps<�?l<�e<=�]<l�V<Z�O<�\H<�5A<T:<��2<.�+<ѻ$<)�<��<��<��<(�<�6�;`Y�;+��;3��;K �;���;���;ޅ�;p$�;<�u;YA[;��@;h�&;:	;���:+��:��:��:�Zi97.!��
���j�c����Ժ����5��;0��G�N�]���s�T넻3Ώ�w���n2��|���h���TĻ�tλKtػ�S���	����5���K����̀����z����E;���#���'�I�+�<0��04�{;8��:<��-@��D���G���K���O��JS���V��Z��J^�\�a��se���h��{l�P�o�oes���v�.3z�7�}�s���������ud���������6>��z׋��n���������(��P����F��2Ӗ��^���虼>q������~��3��������G������
�������������������s������F�������������䟹��!��᣼��&���  �  �lN=��M=H�L=r%L=&bK=X�J=�I=I=�OH=W�G=p�F=��E=a2E=iD=�C=��B=�B=�:A=�l@=h�?=��>=T�==f(==T<=k~;=H�:=��9=f�8=�8=�:7=�[6=pz5=[�4=J�3=3�2=��1=��0=�0=�/=w&.=�1-=:,=�?+=C*=C)=�@(=�;'=3&=|'%=�$=�#=R�!=�� =g�=��=Wy=^R=�'=D�=�=�=�V=�=�=�=G=�=
�=�P=��=��
=F6	=��=�e=i�=0�==� =�.�<�+�<!!�<s�<���<���<=��<���<JO�<F�<!��<��<3C�<���<��<?�<E��<�x�<��<���<k-�<�<�<�<��<>�<��<O3�<멤<�<�<���<n�<�ڒ<�E�<���<�<z��<]�<ӡz<�ps<�?l<�e<3�]<\�V<S�O<�\H<{5A<^:<��2<!�+<˻$<0�<��<ϐ<��<�<�6�;;Y�;_��;\��;> �;���;���;&��;�$�;$�u;A[;b�@;��&;�	;.��:ɮ�:`�:��:wTi9�,!�
�'�j��c����Ժ���5�r;0�G�4�]��s�Z넻0Ώ�u���u2��ĳ��j���TĻltλtػ�S���5���v5���K����ʀ���z����;���#���'�^�+�K0�d04�h;8�e:<��-@��D���G���K���O��JS���V�=�Z��J^�s�a��se���h��{l�K�o��es���v�23z�0�}��s���������|d���������*>���׋��n���������(��N����F��4Ӗ�^��z虼Hq���������0��ꉡ����>��������������������������������R�������������쟹��!��ף���&���  �  �lN=��M=O�L=q%L=%bK=U�J=��I=I=�OH=_�G=m�F=��E=Y2E=iD=��C=��B=�B=�:A=�l@=n�?=��>=Q�==W(==T<=f~;=I�:=��9=i�8=�8=�:7=�[6=nz5=`�4=K�3=3�2=��1=��0=�0=�/=|&.=�1-=:,=�?+=%C*=�C)=�@(=�;'=3&=r'%=�$=�#=V�!=�� =e�=��=[y=dR=�'=B�=��=�=�V=�=��=�=G=�=�=�P=��=��
=B6	= �=�e=q�=-�==� =�.�<�+�<!�<|�<���<���<B��<��<QO�<>�<%��<���<+C�<���<��<?�<8��<�x�<q�<��<c-�<۶�<�<�<��<+>�<*��<N3�<ө�<��<���<���<n�<�ڒ<�E�<ᯋ<�<���<^�<�z<�ps<�?l<�e<G�]<d�V<Y�O<�\H<P5A<r:<��2<;�+<ǻ$<*�<��<��<��<(�<�6�;*Y�;]��;��; �;���;���;���;n$�;#�u;~A[;��@;~�&;�;\��:1��:��:�:[Wi9�,!�_

���j�d����Ժ����5�R;0�ZG���]�!�s�-넻<Ώ�����Y2������6���TĻhtλ�tػ�S������Y5���K���������z����%;���#���'�J�+�@0��04��;8�]:<��-@��D���G���K�֌O��JS���V�B�Z��J^���a��se���h��{l�1�o��es���v�N3z�6�}��s����������d���������2>��z׋��n���������(��_����F��<Ӗ��^��{虼Qq���������0�������@������������옪����������~������V�������������蟹��!��գ���&���  �  �lN=��M=H�L=r%L=&bK=X�J=�I=I=�OH=W�G=p�F=��E=a2E=iD=�C=��B=�B=�:A=�l@=h�?=��>=T�==f(==T<=k~;=H�:=��9=f�8=�8=�:7=�[6=pz5=[�4=J�3=3�2=��1=��0=�0=�/=w&.=�1-=:,=�?+=C*=C)=�@(=�;'=3&=|'%=�$=�#=R�!=�� =g�=��=Wy=^R=�'=D�=�=�=�V=�=�=�=G=�=
�=�P=��=��
=F6	=��=�e=i�=0�==� =�.�<�+�<!!�<s�<���<���<=��<���<JO�<F�<!��<��<3C�<���<��<?�<E��<�x�<��<���<k-�<�<�<�<��<>�<��<O3�<멤<�<�<���<n�<�ڒ<�E�<���<�<z��<]�<ӡz<�ps<�?l<�e<3�]<\�V<S�O<�\H<{5A<^:<��2<!�+<˻$<0�<��<ϐ<��<�<�6�;;Y�;_��;\��;> �;���;���;&��;�$�;$�u;A[;a�@;��&;�	;.��:Ȯ�:`�:��:uTi9�,!�
�(�j��c����Ժ���5�r;0�G�4�]��s�Z넻0Ώ�u���u2��ĳ��j���TĻltλtػ�S���5���v5���K����ʀ���z����;���#���'�^�+�K0�d04�h;8�e:<��-@��D���G���K���O��JS���V�=�Z��J^�s�a��se���h��{l�K�o��es���v�23z�0�}��s���������|d���������*>���׋��n���������(��N����F��4Ӗ�^��z虼Hq���������0��ꉡ����>��������������������������������R�������������쟹��!��ף���&���  �  �lN=��M=K�L=s%L=$bK=Q�J= �I=I=�OH=Y�G=t�F=��E=\2E=iD=�C=��B=�B=�:A=�l@=l�?=��>=O�==b(==T<=n~;=I�:=��9=l�8=�8=�:7=�[6=uz5=[�4=O�3=3�2=��1=��0=�0=�/=w&.=�1-=:,=�?+=(C*=�C)=A(=�;'=
3&=u'%=�$=�#=Q�!=�� =]�=��=Zy=`R=�'=:�=�=ߐ=�V=�=��=
�=G=�=�=�P=��=��
=G6	=��=�e=f�=6�==� =�.�<�+�</!�<i�<���<���<I��<��<MO�<N�<��<��<(C�<���<��<?�<@��<�x�<��<���<n-�<涹<�<�<��<>�<,��<K3�<ީ�<��<ꏝ<���<n�<�ڒ<�E�<���<�<|��<i�<֡z<�ps<�?l<�e<=�]<l�V<Z�O<�\H<�5A<T:<��2<.�+<ѻ$<*�<��<��<��<(�<�6�;`Y�;+��;3��;K �;���;���;ޅ�;p$�;<�u;YA[;��@;h�&;:	;���:*��:�:��:�Zi9<.!��
���j�c����Ժ����5��;0��G�O�]���s�T넻3Ώ�w���n2��|���h���TĻ�tλKtػ�S���	����5���K����̀����z����E;���#���'�I�+�<0��04�{;8��:<��-@��D���G���K���O��JS���V��Z��J^�\�a��se���h��{l�P�o�oes���v�.3z�7�}�s���������ud���������6>��z׋��n���������(��P����F��2Ӗ��^���虼>q������~��3��������G������
�������������������s������F�������������䟹��!��᣼��&���  �  �lN=��M=F�L=r%L='bK=\�J=��I=I=�OH=W�G=r�F=��E=^2E=iD=��C=��B=�B=�:A=�l@=f�?=��>=Q�==_(==T<=l~;=E�:=��9=e�8=�8=�:7=�[6=pz5=Y�4=N�3=2�2=��1=��0=�0=�/=y&.=�1-=:,=�?+=!C*={C)=�@(=�;'=3&=t'%=�$=�#=R�!=�� =f�=��=[y=cR=�'=C�=�=��=�V=�=��=�=G=�=�=�P=��=��
=I6	=��=�e=h�=2�==� =�.�<�+�<#!�<q�<���<���<>��<��<DO�<G�<&��<��<*C�<���< ��<?�<B��<�x�<s�<��<d-�<涹<�<�<��<>�<#��<O3�<۩�<�<�<���< n�<�ڒ<�E�<�<�<}��<\�<ܡz<�ps<�?l<�e<A�]<Z�V<U�O<�\H<n5A<d:<��2<�+<ʻ$<3�<��<��<��<�<�6�;OY�;W��;B��; �;҄�;���;��;�$�;J�u;A[;��@;��&;	;���:ܮ�:��:R�:�Si9
,!�C
���j��c����Ժ����5�{;0�G��]��s�I넻Ώ�����k2����������TĻztλ#tػ�S���5���y5���K����܀����z����;���#���'�`�+�90��04�n;8�g:<��-@��D���G���K�ǌO��JS���V�=�Z��J^�m�a��se���h��{l�T�o��es���v�.3z�6�}��s���������|d���������4>��y׋��n���������(��\����F��;Ӗ��^��~虼Dq���������0���������?������������򘪼���������������O�������������ퟹ��!��أ���&���  �  �lN=��M=O�L=x%L= bK=W�J=��I=I=�OH=Y�G=p�F=��E=a2E=iD=��C=��B=�B=�:A=�l@=g�?=��>=V�==](==T<=f~;=N�:=��9=h�8=�8=�:7=�[6=oz5=^�4=M�3=0�2=��1=��0=�0=�/=z&.=�1-=:,=�?+="C*=�C)= A(=�;'=3&=u'%=�$=�#=Y�!=�� =g�=��=Xy=bR=�'=F�=��=�=�V=�=��=
�=G=�=�=�P=��=��
=E6	=��=�e=p�=/�==� =�.�<�+�<!�<{�<���<���<F��<��<XO�<=�<��<���<3C�<���<���<?�<3��<�x�<m�<��<`-�<붹<�<�<��<#>�<��<Y3�<ک�<��<珝<���<n�<�ڒ<�E�<鯋<�<��<[�<�z<�ps<�?l<{e<K�]<^�V<Y�O<�\H<]5A<n:<��2<>�+<�$<�<��<��<̍<	�<�6�;;Y�;8��;\��; �;΄�;���;(��;Q$�;u�u;A[;��@;��&;�;���:%��:�:�:IVi9�*!��	
���j��c��.�Ժ����5�0;0�LG���]�Q�s�>넻*Ώ�����V2������0���TĻ�tλAtػ�S⻸�F���B5���K����߀���z����;���#���'�g�+�50�x04�};8�|:<��-@��D���G���K�ȌO��JS���V�J�Z��J^�y�a��se���h��{l�:�o��es���v�A3z�4�}��s����������d���������*>��~׋��n���������(��c����F��@Ӗ��^���虼Mq���������&���������I������ ������옪�����������������X�������������럹��!��ң���&���  �  �lN=��M=G�L=p%L=%bK=Z�J=��I=I=�OH=Y�G=t�F=��E=`2E=iD=��C=��B=�B=�:A=�l@=h�?=��>=N�==a(==T<=m~;=F�:=��9=k�8=�8=�:7=�[6=pz5=Z�4=M�3=2�2=��1=��0=�0=�/=|&.=�1-=:,=�?+=$C*=~C)=�@(=�;'=3&=t'%=�$=�#=T�!=�� =c�=��=Xy=`R=�'=A�=��=�=�V=�=��=�=G=�=�=�P=��=��
=G6	=��=�e=h�=2�==� =�.�<�+�<!!�<y�<���<���<I��< ��<HO�<I�<��<	��<&C�<���<��<?�<3��<�x�<w�<���<e-�<붹<�<�<��<>�<%��<P3�<۩�<�<<���<n�<�ڒ<�E�<���<�<���<^�<ۡz<�ps<�?l<�e<?�]<]�V<]�O<�\H<v5A<^:<��2<�+<û$<-�<��<��<��<!�<�6�;aY�;(��;P��;( �;���;���;��;J$�;�u;!A[;��@;V�&;2	;'��:���:!�:B�: Yi9�-!�
�#�j��c����Ժ����5�G;0�G�1�]�1�s�0넻'Ώ�����j2������z���TĻ�tλtػ�S���4���f5���K����Ѐ���z����';���#���'�_�+�30��04�e;8�r:<��-@��D���G���K�ČO��JS���V�D�Z��J^�m�a��se���h��{l�Q�o��es���v�-3z�<�}��s���������yd���������8>��x׋��n���������(��Y����F��;Ӗ��^���虼Aq���������/���������B������������󘪼���������~������N�������������쟹��!��٣���&���  �  �lN=��M=H�L=q%L=#bK=U�J=�I=I=�OH=Q�G=r�F=��E=^2E=iD=�C=��B=�B=�:A=�l@=c�?=��>=K�==f(==T<=j~;=F�:=��9=i�8=�8=�:7=�[6=tz5=Y�4=P�3=4�2=��1=��0=�0=�/=x&.=�1-=:,=�?+=)C*=|C)= A(=�;'=3&=t'%=�$=�#=N�!=�� =`�=��=Xy=`R=�'=?�=�=ސ=�V=�=��=�=G=�=�=�P=��=��
=G6	=��=�e=h�=9�==� =�.�<�+�<+!�<i�<���<���<D��<��<FO�<G�<��<��<C�<���<���<?�<;��<�x�<��<���<i-�<궹<�<�<��<>�<.��<G3�<੤<��<ꏝ<���<n�<�ڒ<�E�< ��<�<}��<a�<ڡz<�ps<�?l<�e<@�]<a�V<\�O<{\H<�5A<O:<��2<"�+<ɻ$<%�<��<Đ<��<4�<Y6�;KY�;3��;B��;: �;���;���;���;j$�;:�u;�@[; A;�&;�	;p��:���:�:<�:"Wi90!��
���j�Qc����Ժ����5��;0��G�'�]���s�R넻5Ώ�l����2��u�������TĻ�tλtػ�S���'����5���K����Ȁ���z����1;���#���'�`�+�;0��04�c;8��:<��-@��D���G���K���O��JS���V�/�Z��J^�S�a��se���h��{l�V�o�xes���v�%3z�?�}��s���������|d���������?>��t׋��n���������(��N����F��7Ӗ��^���虼Dq������{��8���������G�������������������������{������D�������������ꟹ��!��䣼��&���  �  �lN=��M=N�L=s%L="bK=T�J=�I=I=�OH=X�G=q�F=��E=]2E=iD=��C=��B=�B=�:A=�l@=g�?=��>=P�==c(==T<=i~;=I�:=��9=g�8=�8=�:7=�[6=tz5=[�4=P�3=3�2=��1=��0=�0=�/=}&.=�1-=:,=�?+=&C*=�C)= A(=�;'=
3&=w'%=�$=�#=V�!=�� =a�=��=Yy=bR=�'=?�=��=�=�V=�=��=�=G=�=�=�P=��=��
=H6	=��=�e=k�=4�==� =�.�<�+�<(!�<u�<���<���<B��<��<NO�<D�<��<��<)C�<���<��<?�<5��<�x�<u�<��<d-�<涹<�<�<	��<!>�<$��<L3�<㩤<��<ꏝ<���<n�<�ڒ<�E�<���<�<���<Y�<�z<�ps<�?l<�e<J�]<W�V<g�O<�\H<|5A<`:<��2<7�+<ѻ$<�<��<<��<�<�6�;FY�;.��;:��; �;���;���;���;^$�;f�u;A[;��@;p�&;H	;���:q��:f�:3�:JUi9�+!��
���j�Hc����Ժ����5��;0�G���]�8�s�+넻%Ώ�y���u2������^���TĻ�tλKtػ�S���/���W5���K����؀���z����/;���#���'�_�+�>0�|04�z;8�:<��-@��D���G���K���O��JS���V�<�Z��J^�g�a��se���h��{l�L�o�}es���v�03z�1�}��s���������d���������5>��|׋��n���������(��[����F��=Ӗ��^���虼Jq���������2��򉡼���F��������������������������������M���������������!��֣���&���  �  �lN=��M=K�L=n%L=*bK=\�J=��I=I=�OH=[�G=q�F=��E=`2E=iD=��C=��B=�B=�:A=�l@=i�?=��>=T�==](==T<=o~;=E�:=��9=g�8=�8=�:7=�[6=nz5=]�4=O�3=1�2= �1=��0=�0=�/=~&.=�1-=:,=�?+=!C*=�C)=�@(=�;'=3&=v'%=�$=�#=W�!=�� =h�=��=Xy=aR=�'=G�=��=�=�V=�=��=�=G=�=
�=�P=��=��
=F6	=�=�e=o�=/�==� =�.�<�+�<!�<~�<���<���<E��<��<HO�<J�<)��< ��<0C�<���<��<?�<1��<�x�<m�<��<^-�<趹<�<�<	��<&>�<��<S3�<۩�<�<���<���<n�<�ڒ<�E�<<�<���<\�<�z<�ps<�?l<}e<Q�]<^�V<X�O<�\H<e5A<|:<��2<+�+<��$<@�<��<��<��<�<�6�;BY�;9��;O��;��;Ą�;���;!��;M$�;H�u;.A[;\�@;��&;�;���:@��:��:��:�Ui9O(!�(	
���j�d��]�Ժ����5�';0�QG���]�A�s�$넻9Ώ�����G2������h���TĻZtλ+tػ�S���Q���O5���K���������z����;���#���'�i�+�?0�y04�u;8�Z:<��-@��D���G���K���O��JS���V�F�Z��J^�y�a��se���h��{l�?�o��es���v�<3z�(�}��s���������yd���������/>���׋��n�����!����(��b����F��BӖ��^���虼Jq���������+���������8������
������昪�����������������U�������������럹��!��ף���&���  �  �lN=��M=P�L=u%L=#bK=S�J=��I=I=�OH=X�G=p�F=��E=^2E=iD=��C=��B=�B=�:A=�l@=i�?=��>=P�==_(==T<=k~;=J�:=��9=g�8=�8=�:7=�[6=tz5=^�4=N�3=3�2= �1=��0=�0=�/=x&.=�1-=:,=�?+=$C*=�C)=�@(=�;'=
3&=r'%=�$=�#=S�!=�� =a�=��=Wy=_R=�'=?�=��=�=�V=�=��=
�=G=�=�=�P=��=��
=H6	=��=�e=l�=3�==� =�.�<�+�<*!�<r�<���<���<C��<��<QO�<F�<��<��<)C�<���<��<?�<6��<�x�<v�<���<d-�<綹<�<�<	��<>�<!��<P3�<ש�<��<菝<���<n�<�ڒ<�E�<���<�<��<i�<ߡz<�ps<�?l<�e<B�]<r�V<^�O<�\H<u5A<i:<��2<?�+<׻$<%�<��<��<��<�<�6�;9Y�;'��;@��; �;���;���;���;X$�;=�u;-A[;��@;j�&;	;9��:���:��:�:LUi97-!�9
���j�]c��7�Ժ����5�%;0�G��]���s�S넻*Ώ�|���i2������?���TĻ�tλKtػ�S���+���t5���K����݀�	��z����0;���#���'�X�+�?0��04�};8��:<��-@��D���G���K���O��JS���V�'�Z��J^�k�a��se���h��{l�@�o�{es���v�13z�7�}��s���������|d���������5>��~׋��n���������(��Z����F��<Ӗ��^���虼Kq���������/���������H����������������������s������O�������������៹��!��ۣ���&���  �  �lN=��M=D�L=s%L=%bK=X�J=�I=I=�OH=S�G=r�F=��E=]2E=iD=�C=��B=�B=�:A=�l@=c�?=��>=M�==f(==T<=m~;=E�:=��9=i�8=�8=�:7=�[6=wz5=W�4=N�3=7�2=��1=��0=�0=�/=v&.=�1-=:,=�?+=$C*=yC)=A(=�;'=3&=w'%=�$=�#=O�!=�� =a�=��=Wy=^R=�'=>�=�=ߐ=�V=�=��=�=G=�=�=�P=��=��
=M6	=��=�e=c�=8�==� =�.�<�+�</!�<p�<���<���<E��<��<CO�<M�<��<��<'C�<���<���<?�<F��<�x�<�<���<g-�<趹<�<�<��<>�<'��<J3�<橤<�<���<���<�m�<�ڒ<�E�<���<�<��<a�<Сz<�ps<�?l<�e<8�]<\�V<c�O<�\H<5A<_:<��2<�+<ϻ$<-�<��<ʐ<��<%�<c6�;JY�;G��;;��;- �;���;���;慕;�$�;2�u;�@[;��@;E�&;x	;��:��:��:"�:�Vi9�.!��
���j��b���Ժ����5��;0��G�}�]���s�d넻�͏�~���o2����������TĻ�tλtػ�S���.����5���K����р�	��z����6;���#���'�^�+�60�}04�c;8�r:<��-@��D���G���K���O�xJS���V�#�Z��J^�X�a��se���h��{l�_�o�pes���v�3z�=�}��s���������vd���������7>��x׋��n���������(��Q����F��9Ӗ��^���虼Bq���������5������A�������������������������|������B�������������쟹��!��գ���&���  �  �lN=��M=L�L=s%L=$bK=U�J=��I=I=�OH=Y�G=o�F=��E=Z2E=iD=��C=��B=�B=�:A=�l@=g�?=��>=O�==\(==T<=k~;=K�:=��9=o�8=�8=�:7=�[6=sz5=`�4=Q�3=5�2=��1=��0=�0=�/=w&.=�1-=:,=�?+=(C*=�C)=�@(=�;'=	3&=r'%=�$=�#=S�!=�� =c�=��=Yy=aR=�'=A�=��=��=�V=�=��=�=G=�=�=�P=��=��
=H6	=��=�e=n�=8�==� =�.�<�+�<,!�<r�<���<���<T��<��<SO�<G�<��<���<(C�<���<���<?�<7��<�x�<s�<���<c-�<߶�<�<�<	��<!>�<$��<M3�<ש�<��<폝<���<n�<�ڒ<�E�<ꯋ<�<z��<h�<�z<�ps<�?l<�e<O�]<t�V<U�O<�\H<g5A<l:<��2</�+<һ$<(�<��<��<��< �<�6�;9Y�;1��;#��; �;���;���;慕;U$�;�u;�@[;��@;`�&;�;���:���:��:��:�]i9�-!��
��j��c����Ժ����5��;0��G�̈]���s�[넻$Ώ�����<2������O���TĻ�tλTtػ T⻿�:���s5���K��������z����+;���#���'�c�+�20��04��;8�v:<��-@��D���G���K�ԌO��JS���V��Z��J^�V�a��se���h��{l�<�o�xes���v�33z�<�}�us���������}d���������6>��w׋��n���������(��]����F��=Ӗ��^���虼Kq���������1���������D������������옪����������t������C������������������!��ڣ���&���  �  �nN=T�M=N�L=�(L=�eK=��J=��I=I=�TH=0�G=��F={F=�9E=�pD=�C=k�B=�B=KDA=�v@=��?=�>=�>=�4==�`<=��;=(�:=�9={9=9(8=NK7=�l6=�5=��4=>�3=��2=T�1=�1=�0=P//=�=.=eI-=�R,=3Y+=]*=(^)=S\(=�W'=�O&=�D%=�6$=V%#=�"=|� =��=��=�=mt=7J=8=X�=��=�z=6==��=ɵ=�k==�=�u=�=Y�
=�Z	=o�=��=K=��=82=ȷ =�r�<�n�<1c�<?P�< 6�<��<���<��<Ɉ�<M�<G�<r��<�u�<�"�<���<1l�<N	�<ʡ�<�5�<-��<�P�<ع<�[�<?ܲ<PY�<4ӫ<hJ�<꾤<1�<頝<��<�z�<r�<�N�<���<��<3��<�<+�z<js<C5l<� e<k�]<��V<|kO<�=H<�A<p�9<��2<Q�+<��$<Xq<�^<�Q<�J<CJ<[��;=��;3��;� �;�k�;�ȯ;+8�;0��;R�;�s;d�Y;�0?;�%; ;,��:��:4�y:�n:	G9�!D�e����s�!����ٺ�K���E�2��mI��_�PCv�b&��?
��p͛��o���𰻴P��0�Ż��ϻ��ٻ;���G�����1 �}����	���Ȕ�5�2m����$�:H(�~v,���0��4�1�8�P�<�٠@�ԅD��_H�+/L��O�ӮS��_W��[�8�^�<b�D�e�|Ni���l��Ap�.�s��w�xz��}������:��3߃�逅� ������W��^h���v��˫��6<��˓�BX���㖼Sn��h���A�����Ӌ������������/�����h���R��Ӟ�����㞭����N���������r���������X���e��֠���"���  �  oN=[�M=K�L=�(L=�eK=�J=��I=I=�TH=&�G=��F=|F=�9E=�pD=�C=p�B=�B=MDA=�v@=�?=�>=�>=�4==�`<=��;=)�:=�9=�9=B(8=OK7=�l6=�5=��4=A�3=��2=H�1=�1=�0=Q//=�=.=cI-=�R,=<Y+=]*=%^)=X\(=�W'=�O&=�D%=�6$=X%#=�"=z� =��=��=�=rt=:J=5=W�=��=�z=6==��=��=�k==	�=�u=�=_�
=�Z	=l�=�=I=��=-2=· =�r�<�n�<9c�<8P�<!6�<��<���<��<Ɉ�<M�<8�<d��<�u�<�"�<���<l�<Q	�<ơ�<�5�<9��<�P�<ع<�[�</ܲ<9Y�<@ӫ<]J�<ݾ�<�0�<ޠ�<��<�z�<�<�N�<���<��<6��<�<1�z<js<5l<� e<u�]<��V<�kO<�=H<�A<��9<
�2<G�+<�$<Lq<�^<�Q<�J<cJ<��;���;:��;� �;�k�;�ȯ;Q8�;&��;*R�;S�s;�Y;,1?;1%;�;/��:��:�y:�n:�G9D�:���s�������ٺ�K�C��	�2�WmI��_�ACv�s&��L
��?͛�=o��u��P���ŻϮϻ׬ٻ|���G���� 2 ������	������#�%m���$�rH(��v,���0�,�4�T�8�s�<�Ơ@�مD��_H�
/L���O�ڮS� `W��[�@�^�<b�o�e��Ni���l��Ap��s��w�~xz���}������:��3߃�倅� ��ɼ��-W��Qp������ɫ��:<���ʓ�6X���㖼Tn��j���P����ǋ������������:�����o���E���������鞭����R������������}������\���]��ݠ���"���  �  �nN=S�M=G�L=�(L=�eK=��J=��I=I=�TH=(�G=��F=F=9E=�pD=�C=l�B=�B=SDA=�v@=�?=�>=�>=�4==�`<=��;=*�:=�9=z9=<(8=NK7=�l6=�5=��4=B�3=��2=J�1=�1=�0=M//=�=.=cI-=�R,=2Y+=]*=!^)=\\(=�W'=�O&=�D%=�6$=\%#=�"=�� =��=��=�=mt=9J=3=`�=��=�z=5==��=̵=�k==�=�u=�=[�
=�Z	=l�=�=A=��=02=Ʒ =�r�<�n�<<c�<7P�<6�<��<���<��<ƈ�<!M�<>�<x��<�u�<�"�<���<l�<a	�<���<�5�<0��<�P�<ع<�[�<?ܲ<:Y�<Eӫ<XJ�<�<1�<ߠ�<��<�z�<r�<�N�<���<��<;��<�<%�z<0js<
5l<� e<i�]<��V<�kO<�=H<�A<}�9<��2<4�+<��$<Kq<�^<�Q<�J<iJ<��;.��;Q��;y �;�k�;�ȯ;38�;��;^R�;��s;/�Y;71?;	%;P ;���:��:��y:im:�G9GD����"�s�R���m�ٺ�K� ���2�mI�W�_�vCv�p&��K
��a͛��o�����P���Ż��ϻ�ٻP���G�����1 �f����	���˔�7�*m����$�iH(�vv,���0��4�%�8�j�<���@��D��_H�3/L��O�ܮS�`W��[�]�^��;b�c�e��Ni���l��Ap��s��w��xz���}������:��6߃� � ������.W��Pl����������A<��˓�?X���㖼Xn��f���@����Ë������������9�����x���R��Ϟ�����螭����]������������w������h���X��ݠ���"���  �  �nN=X�M=R�L=�(L=�eK=��J=��I=I=�TH=,�G=��F=yF=�9E=�pD=�C=m�B=�B=IDA=�v@=�?=�>=�>=�4==�`<=��;=,�:=%�9=9=>(8=NK7=�l6=�5=��4=B�3=��2=K�1=�1=�0=O//=�=.=fI-=�R,=5Y+=]*=,^)=T\(=�W'=�O&=�D%=�6$=V%#=�"=z� =��=��=�=qt=;J=6=V�=��=�z=5==��=õ=�k=
=�=�u=�=]�
=�Z	=p�=��=N=��=.2=�� =�r�<�n�<2c�<CP�< 6�<��<���<*��<Ј�<M�<=�<h��<�u�<�"�<���<!l�<I	�<ɡ�<�5�<8��<�P�<#ع<�[�<9ܲ<FY�<6ӫ<eJ�<ݾ�<�0�<ޠ�<��<�z�<}�<�N�<���<��<4��<�<@�z<	js<#5l<� e<�]<��V<�kO<�=H<�A<��9<��2<c�+<�$<Eq<�^<�Q<�J<NJ<7��;!��;��;� �;�k�;�ȯ;:8�;.��;	R�;��s;,�Y;�0?;�%;�;���:~��:�y:gp:"G9OD�M����s����*�ٺ�K����ڡ2��mI���_�`Cv�V&��:
��\͛�so��d𰻏P��%�Ż��ϻ��ٻs���G�����1 ������	������#� m���$�[H(��v,���0�"�4�G�8�k�<�Ӡ@�ÅD��_H�$/L��O�֮S��_W��[�+�^�<b�m�e��Ni���l��Ap�+�s��w�~xz���}������:��+߃�퀅� ��ļ��#W��[p������Ы��8<��˓�7X���㖼On��n���G����ы������������:�����_���G��͞������������S��������������������Y���c��Ԡ���"���  �  oN=T�M=K�L=�(L=�eK=��J=��I=I=�TH=,�G=��F=~F=�9E=�pD=
�C=h�B=�B=LDA=�v@=�?=
�>=�>=�4==�`<=��;=%�:=�9=|9=A(8=IK7=�l6=�5=��4=B�3=��2=Q�1=�1=�0=G//=�=.=`I-=�R,=8Y+=]*=&^)=R\(=�W'=�O&=�D%=�6$=T%#=�"=y� =��=��=�=pt=5J=>=V�=��=�z=:==��=µ=�k=	=�=�u=�=^�
=�Z	=o�=׉=O=��=42=÷ =�r�<�n�<$c�<FP�<6�<��<���<��<���<M�<N�<_��<�u�<�"�<���<%l�<N	�<ڡ�<�5�<<��<�P�<%ع<�[�<3ܲ<HY�<4ӫ<nJ�<۾�<1�<ꠝ<��<�z�<s�<�N�<���<��</��<�<I�z< js<>5l<� e<��]<��V<ukO<�=H<�A<��9<��2<D�+<҈$<Zq<�^<�Q<K<MJ<8��;��;I��;� �;�k�;�ȯ;8�;n��;"R�;��s;P�Y;�0?;�%;�;���:���:e�y:�m:�
G9�D����>�s�����n�ٺ�K�b��q�2��mI���_��Cv�j&��h
��O͛�Zo�����P��7�Ż{�ϻ��ٻ]���G������1 ������	���Ɣ�*�8m����$�NH(��v,���0��4�K�8�F�<�֠@���D��_H� /L��O��S��_W��[�&�^�<b�R�e��Ni���l��Ap�G�s��w��xz���}������:��;߃�逅�  ��̼��W��Tm������˫��&<��˓�3X��䖼Mn��c���L����Ӌ������������.���%��n���Q�������枭����\����������u���������b���i��ՠ���"���  �  �nN=T�M=L�L=�(L=�eK=��J=��I=I=�TH=+�G=��F=F=�9E=�pD=	�C=i�B=�B=PDA=�v@=�?=�>=�>=�4==�`<=��;=.�:=�9=|9=>(8=IK7=�l6=�5=��4=A�3=��2=K�1=�1=�0=M//=�=.=`I-=�R,=4Y+=]*=(^)=[\(=�W'=�O&=�D%=�6$=Z%#=�"=~� =��=��=�=rt=6J=9=[�=��=�z=5==��=ĵ=�k==�=�u=�=^�
=�Z	=s�=߉=G=��=/2=�� =�r�<�n�<:c�<CP�<6�<��<���<��<Ј�<M�<:�<m��<�u�<�"�<���< l�<Y	�<ʡ�<�5�<<��<�P�<ع<�[�<;ܲ<BY�<Aӫ<YJ�<侤<�0�<ܠ�<��<�z�<s�<�N�<���<��<B��<�<2�z<js<5l<� e<s�]<��V<�kO<�=H<�A<��9<��2<J�+<�$<Fq<�^<�Q<�J<bJ</��;%��;O��;� �;�k�;�ȯ;8�;*��;AR�;��s;I�Y;1?;%;�;���:���:��y:_n:?
G9�D�����s�:���+�ٺ�K�R��ҡ2�umI���_�}Cv�7&��a
��H͛�o���𰻳P���ŻǮϻ��ٻi���G�����1 �v����	������!�4m�����$�]H(�|v,���0�(�4�B�8�p�<���@�ЅD��_H�./L��O��S��_W��[�H�^�<b�f�e��Ni���l��Ap��s��w��xz���}������:��,߃�倅� ������.W��Tl����������6<��˓�3X���㖼Vn��c���D����Ƌ������������<�����m���P��̞�����랭����Z�������������������g���S��ܠ���"���  �  �nN=[�M=H�L=�(L=�eK=��J=��I=I=�TH=%�G=��F=}F=�9E=�pD=�C=s�B=�B=PDA=�v@=�?=�>=�>=�4==�`<=��;=)�:=�9=�9=<(8=RK7=�l6=�5=��4=B�3=��2=F�1=�1=�0=N//=�=.=`I-=�R,=2Y+=]*= ^)=\\(=�W'=�O&=�D%=�6$=^%#=�"=�� =��=��=�=mt=>J=5=^�=��=�z=8==��=ɵ=�k==�=�u=�=^�
=�Z	=i�=�=F=��=+2=�� =�r�<�n�<9c�<2P�<&6�<��<���<��<Ĉ�<%M�<5�<w��<�u�<�"�<���<l�<Y	�<á�<�5�<-��<�P�<"ع<�[�<@ܲ<4Y�<Kӫ<]J�<뾤<�0�<⠝<��<�z�<��<�N�<Ķ�<��<5��<�<,�z<$js<5l<� e<s�]<��V<�kO<�=H<�A<x�9<	�2<:�+<��$<Tq<�^<�Q<�J<yJ<���;/��;>��;� �;�k�;�ȯ;k8�;��;BR�;��s;�Y;r1?;(%;M ;7��:��:��y:tn:�G9�D�T����s�����A�ٺ�K�T���2�AmI��_�gCv��&��e
��;͛��o��U��P���Żîϻ��ٻi���G�x���2 �f����	���Ȕ�6�m�	���$�pH(�sv,���0�*�4�,�8�p�<���@��D��_H�3/L� �O�ޮS�`W��[�K�^��;b�w�e��Ni���l��Ap��s��w�qxz���}������:��7߃�݀�� ������.W��Kr����������=<���ʓ�BX���㖼Pn��l���?������������������6�����w���@��Ҟ�����𞭼���Z������������������e���^��堼��"���  �  �nN=W�M=J�L=�(L=�eK=��J=��I=I=�TH=*�G=��F=|F=�9E=�pD=�C=o�B=�B=ODA=�v@=�?=�>=�>=�4==�`<=��;='�:=�9=}9=:(8=NK7=�l6=�5=��4=?�3=��2=N�1=�1=�0=N//=�=.=bI-=�R,=2Y+=]*="^)=X\(=�W'=�O&=�D%=�6$=W%#=�"=�� =��=��=�=pt=:J=5=]�=��=�z=8==��=Ƶ=�k==�=�u=�=[�
=�Z	=n�=މ=J=��=12=· =�r�<�n�<0c�<<P�<6�<��<���<��<�<&M�<C�<f��<�u�<�"�<���<-l�<V	�<ǡ�<�5�<6��<�P�< ع<�[�<Gܲ<CY�<9ӫ<bJ�<ᾤ<�0�<頝<��<�z�<z�<�N�<���<��<5��<�<1�z< js<,5l<� e<p�]<��V<�kO<�=H<�A<s�9<��2<@�+<�$<`q<�^<�Q<�J<UJ<+��;T��;9��;� �;�k�;�ȯ;O8�;(��;AR�;�s;+�Y;1?;T%;�;���:���:�y:�m:G9� D�i��K�s�������ٺ�K�\����2��mI���_�mCv�h&��V
��U͛��o�����P���Ż��ϻ��ٻq���G�����1 �h����	������(�#m����$�KH(��v,���0�(�4�;�8�V�<���@��D��_H�//L��O��S��_W��[�9�^� <b�^�e��Ni���l��Ap�+�s��w��xz���}������:��9߃�܀�� ��ż��*W��Qo���z��«��9<���ʓ�9X���㖼Rn��l���8��
��΋������������/�����q���J��Ԟ�����螭����Z���������~���������b���`��۠���"���  �  oN=P�M=O�L=�(L=�eK=��J=��I=I=�TH=.�G=��F=F=�9E=�pD=�C=i�B=�B=MDA=�v@=�?=�>=�>=�4==�`<=��;=/�:=�9=z9=C(8=GK7=�l6=�5=��4=B�3=��2=M�1=�1=�0=H//=�=.=`I-=�R,=:Y+=]*=,^)=U\(=�W'=�O&=�D%=�6$=U%#=�"=w� =��=��=�=ut=8J===T�=��=�z=8==��=��=�k=	=�=�u=�=^�
=�Z	=q�=ى=P=��=/2=�� =�r�<�n�<'c�<DP�<6�<��<���<��<Ԉ�<M�<@�<b��<�u�<�"�<���<l�<L	�<֡�<�5�<C��<�P�<$ع<�[�</ܲ<JY�<8ӫ<iJ�<ᾤ<�0�<֠�<��<�z�<j�<�N�<���<��<5��<	�<S�z<�is<.5l<� e<��]<��V<�kO<�=H<�A<��9<��2<W�+<��$<4q<�^<�Q<�J<TJ<H��;���;V��;� �;�k�;�ȯ; 8�;[��;-R�;��s;H�Y;1?;�%;�;���:��:��y:�n:�G9TD���Z�s�}���x�ٺ�K������2��mI�`�_��Cv�O&��^
��M͛�No���𰻋P���ŻŮϻѬٻe���G������1 ������	�������/m����$�TH(��v,���0��4�P�8�i�<�Ԡ@���D��_H�/L���O��S��_W��[� �^�%<b�f�e��Ni���l��Ap�?�s��w��xz���}������:��'߃�򀅼 ��ɼ��W��To������̫��*<��˓�,X���㖼Nn��a���P����ϋ������������B�����c���Z���������枭����`����������|���������e���c��ؠ���"���  �   oN=S�M=J�L=�(L=�eK=��J=��I=I=�TH=-�G=��F=�F=�9E=�pD=�C=l�B=�B=RDA=�v@=��?=�>=�>=�4==�`<=��;=)�:=�9=z9=?(8=IK7=�l6=�5=��4=C�3=��2=L�1=�1=�0=E//=�=.=_I-=�R,=6Y+=]*=$^)=T\(=�W'=�O&=�D%=�6$=\%#=�"=~� =��=��=�=ot=8J=<=\�=��=�z=8==��=˵=�k=
=�=�u=�=Y�
=�Z	=n�=؉=G=��=02=· =�r�<�n�<*c�<@P�<6�<��<���<��<Ĉ�<M�<L�<r��<�u�<�"�<���<$l�<Z	�<ѡ�<�5�<7��<�P�<#ع<�[�<8ܲ<FY�<Cӫ<aJ�<群<1�<㠝<��<�z�<s�<�N�<���<��<6��<�<7�z<js<!5l<� e<z�]<x�V<�kO<�=H<�A<��9<��2<B�+<�$<Iq<�^<�Q<�J<gJ<C��;��;u��;� �;�k�;�ȯ;78�;H��;XR�;��s;��Y;1?;Z%; ;���:ǩ�:w�y:$n:b	G9SD������s����@�ٺ�K�_����2��mI���_��Cv�f&��i
��n͛�ho�����P��$�Ż��ϻs�ٻU���G�����1 �u����	���Ĕ�.�-m�����$�SH(�rv,���0��4�&�8�M�<�Ѡ@��D��_H�&/L��O��S��_W��[�F�^�<b�b�e��Ni���l��Ap�9�s��w��xz���}������:��6߃�쀅�  ������'W��Ud����������/<��˓�8X���㖼Pn��[���H����ċ������������5�����p���Q��ƞ�����Ɬ����g��������������������n���`��٠���"���  �  �nN=\�M=M�L=�(L=�eK=��J=��I=I=�TH=(�G=��F={F=�9E=�pD=�C=v�B=�B=ODA=�v@=�?=�>=�>=�4==�`<=��;=(�:= �9=�9=9(8=PK7=�l6=�5=��4=>�3=��2=H�1=�1=�0=R//=�=.=cI-=�R,=3Y+=]*=$^)=Z\(=�W'=�O&=�D%=�6$=[%#=�"=�� =��=��=�=rt=@J=0=^�=��=�z=5==�=��=�k==�=�u=�=[�
=�Z	=j�=�=D=��=+2=�� =�r�<�n�<7c�<6P�<!6�<��<���<%��<È�<%M�<6�<d��<�u�<�"�<���< l�<W	�<���<�5�<2��<�P�<ع<�[�<Eܲ<;Y�<@ӫ<]J�<ݾ�<�0�<㠝<��<�z�<��<�N�<���<��<5��<�< �z<js<5l<� e<e�]<��V<�kO<�=H<�A<o�9<�2<O�+<�$<Yq<�^<�Q<�J<cJ<��;I��;1��;� �;l�;�ȯ;�8�;��;>R�;��s;P�Y;1?;F%;�;5��:���:L�y:Qo:�G9� D����-�s�����օٺ�K�s�� �2��mI�5�_�#Cv�w&��N
��K͛��o��P��P����Ż��ϻɬٻ}���G�����1 �d����	������ �m����$�fH(�wv,���0�-�4�L�8�o�<���@��D��_H�&/L��O�ܮS�`W��[�R�^�<b�u�e��Ni���l��Ap��s��w�{xz���}������:��7߃�݀�� ��Ǽ��,W��Vj������«��C<���ʓ�=X���㖼Sn��o���:����ǋ������������5�����k���?��֞�����잭����S���
����������������_���^��ߠ���"���  �  �nN=S�M=G�L=�(L=�eK=��J=��I=I=�TH=)�G=��F=�F=�9E=�pD=�C=r�B=�B=SDA=�v@=�?=�>=�>=�4==�`<=��;='�:=�9=z9=<(8=MK7=�l6=�5=��4=@�3=��2=L�1=�1=�0=I//=�=.=`I-=�R,=2Y+=]*=!^)=X\(=�W'=�O&=�D%=�6$=\%#=�"=�� =��=��=�=nt=<J=7=_�=��=�z=:==��=Ƶ=�k==�=�u=�=[�
=�Z	=g�=ډ=F=��=02=÷ =�r�<�n�<'c�<3P�<6�<��<���<��<���<M�<>�<o��<�u�<�"�<���<l�<^	�<ġ�<�5�<.��<�P�<ع<�[�<@ܲ<=Y�<Cӫ<kJ�<<�0�<᠝<��<�z�<p�<�N�<���<��<+��<�<2�z<js<#5l<� e<t�]<��V<qkO<�=H<�A<~�9<��2<4�+<�$<Pq<�^<�Q<K<jJ< ��;2��;`��;� �;�k�;�ȯ;c8�;#��;eR�;��s;I�Y;E1?;�%;% ;���:+��:*�y:m:�G9�D�p��_�s������ٺ�K�;����2�pmI��_��Cv��&��`
��N͛��o�����P���Ż��ϻ��ٻ/���G�����1 �f����	������/�m�����$�eH(�uv,���0��4�8�8�`�<�Š@��D��_H�2/L�
�O��S�`W��[�I�^�<b�b�e��Ni���l��Ap�>�s��w��xz���}������:��:߃�倅� ������W��Nk����������<<���ʓ�AX���㖼Rn��b���?����ċ������������7�����w���T��Ϟ�����힭����^�������������������f���k��⠼��"���  �  oN=X�M=N�L=�(L=�eK=��J=��I=I=�TH=,�G=��F=�F=9E=�pD=�C=n�B=�B=UDA=�v@=��?=�>=�>=�4==�`<=��;=.�:=�9=�9=@(8=GK7=�l6=�5=��4=@�3=��2=F�1=�1=�0=I//=�=.=dI-=�R,=;Y+=]*=)^)=U\(=�W'=�O&=�D%=�6$=\%#=�"=~� =��=��=�=xt=7J=:=\�=��=�z=3==��=µ=�k==�=�u=�=Z�
=�Z	=v�=ډ=H=��=+2=�� =�r�<�n�<.c�<LP�<6�<��<���<!��<ш�<M�<E�<d��<�u�<�"�<���<"l�<^	�<á�<�5�<I��<�P�<ع<�[�<8ܲ<EY�<Aӫ<XJ�<޾�< 1�<ܠ�<��<�z�<{�<�N�<���<��<A��<�<6�z<js<
5l<� e<u�]<��V<�kO<�=H<yA<��9<��2<R�+<��$<>q<�^<�Q<�J<aJ<>��;��;~��; �;�k�;ɯ;F8�;��;oR�;��s;x�Y;1?;2%;�;8��:���:��y:0o:�G9�D����y�s�����хٺ�K�����2��mI���_��Cv�!&��D
��r͛�Co��r𰻥P��!�Ż��ϻ��ٻo��H�����1 �v����	������	�/m�����$�[H(�pv,���0�%�4�H�8�]�<�ؠ@�ɅD��_H�/L��O�߮S��_W��[�?�^�<b�u�e��Ni���l��Ap�.�s��w��xz���}������:��)߃�퀅� ��Ǽ��,W��Yf����������=<��˓�'X���㖼Yn��Y���G����ǋ������������<�����h���I��������➭����b��������������������j���X��Р���"���  �  �nN=S�M=G�L=�(L=�eK=��J=��I=I=�TH=)�G=��F=�F=�9E=�pD=�C=r�B=�B=SDA=�v@=�?=�>=�>=�4==�`<=��;='�:=�9=z9=<(8=MK7=�l6=�5=��4=@�3=��2=L�1=�1=�0=I//=�=.=`I-=�R,=2Y+=]*=!^)=X\(=�W'=�O&=�D%=�6$=\%#=�"=�� =��=��=�=nt=<J=7=_�=��=�z=:==��=Ƶ=�k==�=�u=�=[�
=�Z	=g�=ډ=F=��=02=÷ =�r�<�n�<'c�<3P�<6�<��<���<��<���<M�<>�<o��<�u�<�"�<���<l�<^	�<ġ�<�5�<.��<�P�<ع<�[�<@ܲ<=Y�<Cӫ<kJ�<<�0�<᠝<��<�z�<p�<�N�<���<��<+��<�<2�z<js<#5l<� e<t�]<��V<qkO<�=H<�A<~�9<��2<4�+<�$<Qq<�^<�Q<K<jJ<!��;2��;`��;� �;�k�;�ȯ;c8�;#��;eR�;��s;I�Y;D1?;�%;% ;���:*��:)�y:m:�G9�D�q��`�s������ٺ�K�;����2�pmI��_��Cv��&��`
��N͛��o�����P���Ż��ϻ��ٻ/���G�����1 �f����	������/�m�����$�eH(�uv,���0��4�8�8�`�<�Š@��D��_H�2/L�
�O��S�`W��[�I�^�<b�b�e��Ni���l��Ap�>�s��w��xz���}������:��:߃�倅� ������W��Nk����������<<���ʓ�AX���㖼Rn��b���?����ċ������������7�����w���T��Ϟ�����힭����^�������������������f���k��⠼��"���  �  �nN=\�M=M�L=�(L=�eK=��J=��I=I=�TH=(�G=��F={F=�9E=�pD=�C=v�B=�B=ODA=�v@=�?=�>=�>=�4==�`<=��;=(�:= �9=�9=9(8=PK7=�l6=�5=��4=>�3=��2=H�1=�1=�0=R//=�=.=cI-=�R,=3Y+=]*=$^)=Z\(=�W'=�O&=�D%=�6$=[%#=�"=�� =��=��=�=rt=@J=0=^�=��=�z=5==�=��=�k==�=�u=�=[�
=�Z	=k�=�=D=��=+2=�� =�r�<�n�<7c�<6P�<!6�<��<���<%��<È�<%M�<6�<d��<�u�<�"�<���< l�<W	�<���<�5�<2��<�P�<ع<�[�<Eܲ<;Y�<@ӫ<]J�<ݾ�<�0�<㠝<��<�z�<��<�N�<���<��<5��<�< �z<js<5l<� e<e�]<��V<�kO<�=H<�A<o�9<�2<O�+<�$<Yq<�^<�Q<�J<cJ<��;I��;1��;� �;l�;�ȯ;�8�;��;>R�;��s;P�Y;1?;F%;�;5��:���:J�y:Oo:�G9� D����/�s�����ׅٺ�K�s���2��mI�5�_�#Cv�w&��N
��K͛��o��P��P����Ż��ϻɬٻ}���G�����1 �d����	������ �m����$�fH(�wv,���0�-�4�L�8�o�<���@��D��_H�&/L��O�ܮS�`W��[�R�^�<b�u�e��Ni���l��Ap��s��w�{xz���}������:��7߃�݀�� ��Ǽ��,W��Vj������«��C<���ʓ�=X���㖼Sn��o���:����ǋ������������5�����k���?��֞�����잭����S���
����������������_���^��ߠ���"���  �   oN=S�M=J�L=�(L=�eK=��J=��I=I=�TH=-�G=��F=�F=�9E=�pD=�C=l�B=�B=RDA=�v@=��?=�>=�>=�4==�`<=��;=)�:=�9=z9=?(8=IK7=�l6=�5=��4=C�3=��2=L�1=�1=�0=E//=�=.=_I-=�R,=6Y+=]*=$^)=T\(=�W'=�O&=�D%=�6$=\%#=�"=~� =��=��=�=ot=8J=<=\�=��=�z=8==��=˵=�k=
=�=�u=�=Y�
=�Z	=n�=؉=G=��=02=· =�r�<�n�<*c�<@P�<6�<��<���<��<Ĉ�<M�<M�<r��<�u�<�"�<���<$l�<Z	�<ѡ�<�5�<7��<�P�<#ع<�[�<8ܲ<FY�<Cӫ<aJ�<群<1�<㠝<��<�z�<s�<�N�<���<��<6��<�<7�z<js<!5l<� e<{�]<x�V<�kO<�=H<�A<��9<��2<B�+<�$<Jq<�^<�Q<�J<gJ<C��;��;u��;� �;�k�;�ȯ;78�;H��;XR�;��s;��Y;1?;Z%; ;���:Ʃ�:u�y:"n:Y	G9]D������s����B�ٺ�K�`����2��mI���_��Cv�f&��i
��n͛�ho�����P��%�Ż��ϻs�ٻU���G�����1 �u����	���Ĕ�.�-m�����$�SH(�rv,���0��4�&�8�M�<�Ѡ@��D��_H�&/L��O��S��_W��[�F�^�
<b�b�e��Ni���l��Ap�9�s��w��xz���}������:��6߃�쀅�  ������'W��Ud����������/<��˓�8X���㖼Pn��[���H����ċ������������5�����p���Q��ƞ�����Ɬ����g��������������������n���`��٠���"���  �  oN=P�M=O�L=�(L=�eK=��J=��I=I=�TH=.�G=��F=F=�9E=�pD=�C=i�B=�B=MDA=�v@=�?=�>=�>=�4==�`<=��;=/�:=�9=z9=C(8=GK7=�l6=�5=��4=B�3=��2=M�1=�1=�0=H//=�=.=`I-=�R,=:Y+=]*=,^)=U\(=�W'=�O&=�D%=�6$=U%#=�"=w� =��=��=�=ut=8J===T�=��=�z=8==��=��=�k=	=�=�u=�=^�
=�Z	=q�=ى=P=��=/2=�� =�r�<�n�<'c�<DP�<6�<��<���<��<Ԉ�<M�<@�<b��<�u�<�"�<���<l�<L	�<֡�<�5�<C��<�P�<$ع<�[�</ܲ<JY�<8ӫ<iJ�<ᾤ<�0�<֠�<��<�z�<i�<�N�<���<��<5��<	�<S�z<�is<.5l<� e<��]<��V<�kO<�=H<�A<��9<��2<W�+<��$<4q<�^<�Q<�J<TJ<I��;���;V��;� �;�k�;�ȯ; 8�;[��;-R�;�s;H�Y;1?;�%;�;���:��:��y:�n:�G9_D���]�s�~���y�ٺ�K������2��mI�a�_��Cv�O&��_
��M͛�Oo���𰻌P���ŻŮϻѬٻe���G������1 ������	�������/m����$�TH(��v,���0��4�P�8�i�<�Ԡ@���D��_H�/L���O��S��_W��[� �^�%<b�f�e��Ni���l��Ap�?�s��w��xz���}������:��'߃�򀅼 ��ɼ��W��To������̫��*<��˓�,X���㖼Nn��a���P����ϋ������������B�����c���Z���������枭����`����������|���������e���c��ؠ���"���  �  �nN=W�M=J�L=�(L=�eK=��J=��I=I=�TH=*�G=��F=|F=�9E=�pD=�C=o�B=�B=ODA=�v@=�?=�>=�>=�4==�`<=��;='�:=�9=}9=:(8=NK7=�l6=�5=��4=?�3=��2=N�1=�1=�0=N//=�=.=bI-=�R,=2Y+=]*="^)=X\(=�W'=�O&=�D%=�6$=W%#=�"=�� =��=��=�=pt=:J=5=]�=��=�z=8==��=Ƶ=�k==�=�u=�=[�
=�Z	=n�=މ=J=��=12=· =�r�<�n�<0c�<<P�<6�<��<���<��<�<&M�<C�<g��<�u�<�"�<���<-l�<V	�<ǡ�<�5�<6��<�P�< ع<�[�<Gܲ<CY�<9ӫ<bJ�<ᾤ<�0�<頝<��<�z�<z�<�N�<���<��<5��<�<1�z< js<,5l<� e<p�]<��V<�kO<�=H<�A<s�9<��2<A�+<�$<`q<�^<�Q<�J<UJ<+��;T��;9��;� �;�k�;�ȯ;O8�;(��;AR�;�s;*�Y;1?;T%;�;���:���:�y:�m:G9� D�l��N�s�������ٺ�K�]����2��mI���_�mCv�h&��W
��U͛��o�����P���Ż��ϻ��ٻq���G�����1 �h����	������(�#m����$�KH(��v,���0�(�4�;�8�V�<���@��D��_H�//L��O��S��_W��[�9�^� <b�^�e��Ni���l��Ap�+�s��w��xz���}������:��9߃�܀�� ��ż��*W��Qo���z��«��9<���ʓ�9X���㖼Rn��l���8��
��΋������������/�����q���J��Ԟ�����螭����Z���������~���������b���`��۠���"���  �  �nN=[�M=H�L=�(L=�eK=��J=��I=I=�TH=%�G=��F=}F=�9E=�pD=�C=s�B=�B=PDA=�v@=�?=�>=�>=�4==�`<=��;=)�:=�9=�9=<(8=RK7=�l6=�5=��4=B�3=��2=F�1=�1=�0=N//=�=.=`I-=�R,=2Y+=]*= ^)=\\(=�W'=�O&=�D%=�6$=^%#=�"=�� =��=��=�=mt=>J=5=^�=��=�z=8==��=ɵ=�k==�=�u=�=^�
=�Z	=i�=�=F=��=+2=�� =�r�<�n�<9c�<2P�<&6�<��<���<��<ň�<%M�<5�<w��<�u�<�"�<���<l�<Y	�<á�<�5�<-��<�P�<"ع<�[�<@ܲ<4Y�<Kӫ<]J�<뾤<�0�<⠝<��<�z�<��<�N�<Ķ�<��<5��<�<,�z<$js<5l<� e<s�]<��V<�kO<�=H<�A<x�9<	�2<;�+<��$<Tq<�^<�Q<�J<yJ<���;/��;>��;� �;�k�;�ȯ;k8�;��;BR�;��s;�Y;q1?;'%;L ;6��:~��:��y:qn:�G9�D�X����s�����B�ٺ�K�U���2�BmI��_�hCv��&��f
��;͛��o��U��P���Żîϻ��ٻi���G�x���2 �f����	���Ȕ�6�m�	���$�pH(�sv,���0�*�4�,�8�p�<���@��D��_H�3/L� �O�ޮS�`W��[�K�^��;b�w�e��Ni���l��Ap��s��w�qxz���}������:��7߃�݀�� ������.W��Kr����������=<���ʓ�BX���㖼Pn��l���?������������������6�����w���@��Ҟ�����𞭼���Z������������������e���^��堼��"���  �  �nN=T�M=L�L=�(L=�eK=��J=��I=I=�TH=+�G=��F=F=�9E=�pD=	�C=i�B=�B=PDA=�v@=�?=�>=�>=�4==�`<=��;=.�:=�9=|9=>(8=IK7=�l6=�5=��4=A�3=��2=K�1=�1=�0=M//=�=.=`I-=�R,=4Y+=]*=(^)=[\(=�W'=�O&=�D%=�6$=Z%#=�"=~� =��=��=�=rt=6J=9=[�=��=�z=5==��=ĵ=�k==�=�u=�=^�
=�Z	=s�=��=G=��=/2=�� =�r�<�n�<:c�<CP�<6�<��<���<��<Ј�<M�<:�<m��<�u�<�"�<���< l�<Y	�<ʡ�<�5�<<��<�P�<ع<�[�<;ܲ<BY�<Aӫ<YJ�<侤<�0�<ܠ�<��<�z�<s�<�N�<���<��<B��<�<2�z<js<5l<� e<s�]<��V<�kO<�=H<�A<��9<��2<J�+<�$<Fq<�^<�Q<�J<bJ</��;%��;O��;� �;�k�;�ȯ;8�;*��;AR�;��s;I�Y;1?;%;�;���:���:��y:\n:2
G9�D�����s�<���,�ٺ�K�S��ӡ2�vmI���_�}Cv�8&��a
��H͛�o���𰻳P���ŻȮϻ��ٻi���G�����1 �v����	������!�4m�����$�]H(�|v,���0�(�4�B�8�p�<���@�ЅD��_H�./L��O��S��_W��[�H�^�<b�f�e��Ni���l��Ap��s��w��xz���}������:��,߃�倅� ������.W��Tl����������6<��˓�3X���㖼Vn��c���D����Ƌ������������<�����m���P��̞�����랭����Z�������������������g���S��ܠ���"���  �  oN=T�M=K�L=�(L=�eK=��J=��I=I=�TH=,�G=��F=~F=�9E=�pD=
�C=h�B=�B=LDA=�v@=�?=
�>=�>=�4==�`<=��;=%�:=�9=|9=A(8=IK7=�l6=�5=��4=B�3=��2=Q�1=�1=�0=G//=�=.=`I-=�R,=8Y+=]*=&^)=R\(=�W'=�O&=�D%=�6$=T%#=�"=y� =��=��=�=pt=5J=>=V�=��=�z=:==��=µ=�k=	=�=�u=�=^�
=�Z	=o�=׉=O=��=42=÷ =�r�<�n�<$c�<FP�<6�<��<���<��<���<M�<N�<`��<�u�<�"�<���<%l�<N	�<ڡ�<�5�<<��<�P�<%ع<�[�<3ܲ<HY�<4ӫ<nJ�<۾�<1�<ꠝ<��<�z�<s�<�N�<���<��</��<�<I�z< js<>5l<� e<��]<��V<ukO<�=H<�A<��9<��2<D�+<҈$<Zq<�^<�Q<K<MJ<8��;��;I��;� �;�k�;�ȯ;8�;n��;!R�;��s;O�Y;�0?;�%;�;���:���:b�y:�m:�
G9�D����A�s�����o�ٺ�K�b��r�2��mI���_��Cv�j&��h
��P͛�Zo�����P��7�Ż{�ϻ��ٻ]���G������1 ������	���Ɣ�*�8m����$�NH(��v,���0��4�K�8�F�<�֠@���D��_H� /L��O��S��_W��[�&�^�<b�R�e��Ni���l��Ap�G�s��w��xz���}������:��;߃�逅�  ��̼��W��Tm������˫��&<��˓�3X��䖼Mn��c���L����Ӌ������������.���%��n���Q�������枭����\����������u���������b���i��ՠ���"���  �  �nN=X�M=R�L=�(L=�eK=��J=��I=I=�TH=,�G=��F=yF=�9E=�pD=�C=m�B=�B=IDA=�v@=�?=�>=�>=�4==�`<=��;=,�:=%�9=9=>(8=NK7=�l6=�5=��4=B�3=��2=K�1=�1=�0=O//=�=.=fI-=�R,=5Y+=]*=,^)=T\(=�W'=�O&=�D%=�6$=V%#=�"=z� =��=��=�=qt=<J=6=V�=��=�z=5==��=õ=�k=
=�=�u=�=]�
=�Z	=p�=��=N=��=.2=�� =�r�<�n�<2c�<CP�< 6�<��<���<*��<Ј�<M�<=�<h��<�u�<�"�<���<!l�<I	�<ɡ�<�5�<8��<�P�<#ع<�[�<9ܲ<FY�<6ӫ<eJ�<ݾ�<�0�<ޠ�<��<�z�<}�<�N�<���<��<4��<�<@�z<	js<#5l<� e<�]<��V<�kO<�=H<�A<��9<��2<c�+<�$<Eq<�^<�Q<�J<NJ<7��;!��;��;� �;�k�;�ȯ;:8�;.��;	R�;��s;+�Y;�0?;�%;�;���:}��:�y:ep:G9YD�P����s����+�ٺ�K����ڡ2��mI���_�aCv�W&��:
��\͛�so��d𰻐P��%�Ż��ϻ��ٻs���G�����1 ������	������#� m���$�[H(��v,���0�"�4�G�8�k�<�Ӡ@�ÅD��_H�$/L��O�֮S��_W��[�+�^�<b�m�e��Ni���l��Ap�+�s��w�~xz���}������:��+߃�퀅� ��ļ��#W��[p������Ы��8<��˓�7X���㖼On��n���G����ы������������:�����_���G��͞������������S��������������������Y���c��Ԡ���"���  �  �nN=S�M=G�L=�(L=�eK=��J=��I=I=�TH=(�G=��F=F=9E=�pD=�C=l�B=�B=SDA=�v@=�?=�>=�>=�4==�`<=��;=*�:=�9=z9=<(8=NK7=�l6=�5=��4=B�3=��2=J�1=�1=�0=M//=�=.=cI-=�R,=2Y+=]*=!^)=\\(=�W'=�O&=�D%=�6$=\%#=�"=�� =��=��=�=mt=9J=3=`�=��=�z=5==��=̵=�k==�=�u=�=[�
=�Z	=l�=�=A=��=02=Ʒ =�r�<�n�<<c�<8P�<6�<��<���<��<ƈ�<!M�<>�<x��<�u�<�"�<���<l�<a	�<���<�5�<0��<�P�<ع<�[�<?ܲ<:Y�<Eӫ<XJ�<�<1�<ߠ�<��<�z�<r�<�N�<���<��<;��<�<%�z<0js<
5l<� e<i�]<��V<�kO<�=H<�A<}�9<��2<4�+<��$<Kq<�^<�Q<�J<iJ<��;.��;Q��;y �;�k�;�ȯ;38�;��;^R�;��s;/�Y;71?;	%;O ;���:��:��y:gm:�G9ND����#�s�S���n�ٺ�K� ���2�mI�X�_�vCv�p&��K
��a͛��o�����P���Ż��ϻ�ٻP���G�����1 �f����	���˔�7�*m����$�iH(�vv,���0��4�%�8�j�<���@��D��_H�3/L��O�ܮS�`W��[�]�^��;b�c�e��Ni���l��Ap��s��w��xz���}������:��6߃� � ������.W��Pl����������A<��˓�?X���㖼Xn��f���@����Ë������������9�����x���R��Ϟ�����螭����]������������w������h���X��ݠ���"���  �  oN=[�M=K�L=�(L=�eK=�J=��I=I=�TH=&�G=��F=|F=�9E=�pD=�C=p�B=�B=MDA=�v@=�?=�>=�>=�4==�`<=��;=)�:=�9=�9=B(8=OK7=�l6=�5=��4=A�3=��2=H�1=�1=�0=Q//=�=.=cI-=�R,=<Y+=]*=%^)=X\(=�W'=�O&=�D%=�6$=X%#=�"=z� =��=��=�=rt=:J=5=W�=��=�z=6==��=��=�k==	�=�u=�=_�
=�Z	=l�=�=I=��=-2=· =�r�<�n�<9c�<8P�<!6�<��<���<��<Ɉ�<M�<8�<d��<�u�<�"�<���<l�<Q	�<ơ�<�5�<9��<�P�<ع<�[�</ܲ<8Y�<@ӫ<]J�<ݾ�<�0�<ޠ�<��<�z�<�<�N�<���<��<6��<�<1�z<js<5l<� e<u�]<��V<�kO<�=H<�A<��9<
�2<G�+<�$<Lq<�^<�Q<�J<cJ<��;���;:��;� �;�k�;�ȯ;Q8�;&��;*R�;S�s;�Y;,1?;1%;�;.��:��:~�y:�n:�G9D�;���s�������ٺ�K�C��	�2�XmI��_�ACv�s&��L
��?͛�=o��u��P���ŻϮϻ׬ٻ|���G���� 2 ������	������#�%m���$�rH(��v,���0�,�4�T�8�s�<�Ơ@�مD��_H�
/L���O�ڮS� `W��[�@�^�<b�o�e��Ni���l��Ap��s��w�~xz���}������:��3߃�倅� ��ɼ��-W��Qp������ɫ��:<���ʓ�6X���㖼Tn��j���P����ǋ������������:�����o���E���������鞭����R������������}������\���]��ݠ���"���  �  rqN=1�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=LAE=�xD=ͯC=��B=�B=�NA=��@=s�?=�>=�>=�A==�n<=<�;=O�:=��9=�9=f98= ]7=+6=Q�5=��4=��3=O�2=�2=�"1=b60=�G/=�V.=vc-=ym,=�t+=�y*=\{)=Lz(=Uv'=@o&=e%=�W$= G#= 3"=�!=�  =��=ÿ=ؙ=)p=�B=6=��=�=#e=�#=%�=��=�F=��=��=OD=��
=@�	=�=��=�B=��=�X=�� =��<���<ʫ�<���<�{�<)Y�<x/�<��<���<r��<�F�<���<b��<X�<k��<���<�8�<���<�`�<��<5w�<���<~�<8��<w�<��<�c�<�դ<�E�<x��<�<��<R�<IX�<��<#�<(��<��<S�z<�bs<y)l<��d<�]<��V<NO<�H<N�@<�9<��2<�q+<Q$<65<[<�<�<�� <���;��;O1�;1c�;ǥ�;t��;�a�;�ܓ;}k�;�r;��W;�4=;�#;l	;�s�:�?�:��p:"4:(Z!9��j�G����}����J�޺u��I3��D5��L���b���x�����f���)��$̧�M�������ƻ�ѻRۻ��仏��y5��
� �Ѕ��#
�ٲ��2�����>Z �v�$���(�8-�J"1��35��89��1=��A�� E�r�H���L�.eP��T���W� o[�X
_��b�('f�C�i��#m�>�p��t�Jfw�`�z��~�����z\������򟅼�=��Bو�\r��a	��I���/1��W��Q��hߓ��k��F�������������T��3��������^"������%��s����%��+����$�������"��}���K ��7���.��t���������������������  �  rqN=0�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=MAE=�xD=үC=��B=�B=�NA=��@=p�?=!�>=�>=�A==�n<==�;=R�:=��9=�9=i98=(]7=*6=W�5=��4=��3=I�2=2=�"1=]60=�G/=�V.=zc-=�m,=�t+=�y*=]{)=Sz(=Nv'=>o&=e%=�W$=G#=�2"=�!=�  =��=ȿ=ݙ=-p=�B=7=��=��="e=�#=%�=~�=�F=��=��=OD=��
=D�	=�=��=�B=��=�X=�� =��<���<ի�<���<�{�<0Y�<z/�<	��<���<x��<�F�<���<X��<X�<l��<���<�8�<���<�`�<��<Cw�<���<~�</��<�v�<��<�c�<�դ<�E�<o��<�<��<P�<JX�<$��<#�<0��<��<E�z<�bs<G)l<��d<�]<��V<(NO<�H<n�@<�9<�2<�q+</Q$<,5<F<<�<�� <J��;��;g1�;;c�;���;���;�a�;�ܓ;�k�;Cr;l�W;35=;�#;�	;�r�:@�:��p:}3:�[!9Ӏj�b����}����b�޺����3��E5��L��b���x������e���)��!̧�M��������ƻ ѻ]ۻ��仡��G5��*� �҅��#
�ʲ��2�����:Z �s�$��(�&-�K"1��35��89��1=��A�� E�t�H���L�eP��T���W�
o[�g
_��b�Q'f�]�i��#m�J�p��t�Nfw�G�z��~�����~\������쟅��=��>و�er��[	��I���A1��S��Q��]ߓ��k��8�������������d��"��������d"�������$��v����%��*���~$�������"��v���R ��:���G��x���������������������  �  oqN=5�M=��L=�,L=jK=�J=��I={I=�ZH=��G=��F=�F=HAE=�xD=ͯC=��B=�B=�NA=��@=t�?="�>=�>=�A==�n<=>�;=S�:=��9=�9=f98=']7=$6=X�5=��4=��3=Q�2=�2=�"1=Z60=�G/=�V.=tc-=}m,=�t+=�y*=Y{)=Tz(=Lv'=Eo&=e%=�W$=	G#=�2"=�!=�  =��=Ŀ=ٙ=)p=�B=<=��=��= e=�#=-�=|�=�F=��=��=PD=��
=A�	=�=��=�B=��=�X=�� =��<���<ګ�<{��<�{�<+Y�<}/�<��<���<{��<�F�<��<P��<X�<u��<���<�8�<���<�`�<��<>w�<���<~�<=��<�v�<��<�c�<�դ<�E�<i��<�<���<X�<HX�<!��<�"�<-��<��<?�z<�bs<Z)l<��d<ݸ]<��V<%NO<�H<h�@<�9<�2<�q+<2Q$<&5<Q<<�<�� <f��;��;j1�;c�;�;x��;�a�;|ܓ;�k�;�r;��W;65=;@#;�	;�r�:C@�:��p:�2:�^!9��j������}������޺v��&3�UE5�RL��b�X�x�����(f���)��̧��L��������ƻ2ѻ%ۻ������05��#� �����#
�ݲ��2�����BZ �]�$��(�-�U"1��35��89��1=��A�� E�n�H���L�%eP��T���W��n[�r
_��b�6'f�=�i�#m�T�p��t�efw�O�z��~������\������韅��=��0و�nr��\	��@���81��K��Q��cߓ��k��<�������������^����������["������$��}���|%��,����$�������"��s���U ��*���>��g���������������������  �  qqN=4�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=NAE=�xD=ԯC=��B=�B=�NA=��@=p�?= �>=�>=�A==�n<=<�;=S�:=��9=�9=h98=&]7=(6=S�5=��4=��3=K�2=�2=�"1=^60=�G/=�V.=yc-=}m,=�t+=�y*=Z{)=Pz(=Qv'=?o&=e%=�W$= G#=�2"=�!=�  =��=ɿ=ޙ=+p=�B=5=��=�=$e=�#=%�=��=�F=��=��=SD=��
=C�	=�=��=�B=��=�X=�� =��<���<ϫ�<���<�{�<.Y�<~/�<��<���<s��<�F�<���<Y��<X�<i��<���<�8�<���<�`�<��<Bw�<���<~�<3��<w�<��<�c�<�դ<�E�<s��<�<���<V�<MX�<��<#�<*��<��<J�z<�bs<V)l<��d<�]<��V<NO<�H<f�@<�9<�2<�q+<'Q$<05<R<�<�<�� <s��;��;E1�;Dc�;���;���;�a�;�ܓ;xk�;�r;s�W;5=;�#;f	;Ts�:�?�:��p:�2:�^!9n�j�ذ�_�}�8���޺����3�xE5��L�ۦb���x�퀇�f���)�� ̧�M��������ƻѻ[ۻ��仔��u5��� �҅��#
�ϲ��2�����9Z �z�$���(�5-�F"1��35��89��1=��A�� E�s�H�w�L�eP��T���W�o[�a
_��b�E'f�S�i��#m�=�p��t�Tfw�O�z��~������\������🅼�=��Bو�dr��^	��K���21��Y��Q��^ߓ��k��8�������������X��-��������a"������%��z���~%��(����$�������"��x���O ��=���@��w���������������������  �  rqN=.�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=OAE=�xD=կC=��B=�B=�NA=��@=p�?=!�>=�>=�A==�n<=7�;=V�:=��9=�9=h98=#]7=,6=P�5=��4=��3=L�2=�2=�"1=a60=�G/=�V.=xc-=}m,=�t+=y*=_{)=Mz(=Sv'=>o&=e%=�W$= G#=3"=�!=�  =��=ſ=ܙ=%p=�B=4=��=~�=(e=�#=$�=��=�F=��=��=QD=��
=@�	=�=��=�B=��=�X=�� =��<ĸ�<ƫ�<���<�{�</Y�<y/�<��<���<l��<�F�<���<c��< X�<h��<���<�8�<���<�`�<��<7w�<���<~�<,��<w�<��<�c�<�դ<�E�<r��<�<��<I�<MX�<��<#�<&��<��<R�z<�bs<t)l<��d<�]<��V<NO<H<Y�@<��9<�2<�q+<2Q$<(5<U<�<�<�� <t��;��;^1�;Hc�;ƥ�;���;�a�;�ܓ;�k�;�r;j�W;15=;#;?	;�s�:e?�:��p:�2:�Z!9u�j�����}������޺���q3�E5�L���b���x�����	f���)��̧�)M��}���	�ƻ�ѻ\ۻ���d��t5��� �څ��#
����2�����.Z ��$���(�;-�5"1��35��89��1=��A�� E���H���L� eP��T���W�(o[�W
_��b�*'f�F�i��#m�6�p��t�Ifw�]�z��~������\�����������=��Hو�Zr��X	��M���/1��Z��Q��lߓ�k��D�������������V��-���������`"�������$��r����%��(����$�������"�����L ��A���1��z���������������������  �  sqN=2�M=��L=�,L=	jK=�J=��I=|I=�ZH=��G=��F=�F=KAE=�xD=ׯC=��B=�B=�NA=��@=s�?= �>=�>=�A==�n<=:�;=U�:=��9=�9=h98=$]7=&6=W�5=��4=��3=K�2=�2=�"1=Y60=�G/=�V.=uc-=|m,=�t+=�y*=[{)=Qz(=Lv'=Go&=e%=�W$=G#=�2"=�!=�  =��=˿=�=)p=�B=8=��=��=!e=�#=-�=|�=�F=��=��=QD=��
=>�	=�=��=�B=��=�X=�� =��<���<ի�<��<�{�<,Y�<~/�<��<���<t��<�F�<���<T��<X�<p��<���<�8�<���<�`�<��<Cw�<���<~�<8��<w�<��<�c�<�դ<�E�<g��<�<���<U�<OX�<��<�"�</��<��<:�z<�bs<\)l<��d<ظ]<��V<$NO<�H<Z�@<��9<��2<�q+<7Q$<5<_<<�<�� <}��;��;d1�;/c�;���;���;�a�;�ܓ;�k�;�r;��W;%5=;h#;�	;*s�:�?�:��p:�2:�^!9�j�-����}����{�޺����3�TE5��L�$�b�b�x�����&f���)��̧�M��������ƻ2ѻۻ��仮��S5��� �Ņ��#
�ڲ��2�����:Z �n�$���(�(-�O"1��35��89��1=��A�� E�y�H�~�L�$eP��T���W��n[�r
_��b�;'f�P�i��#m�M�p��t�]fw�Z�z��~������\������🅼�=��5و�ir��^	��E���81��S��Q��`ߓ�zk��7�������������Z��'��������V"������$��z���%��%����$�������"��w���W ��;���=��x���������������������  �  mqN=6�M=��L=�,L=jK=�J=��I=~I=�ZH=��G=��F=�F=NAE=�xD=ͯC=��B=�B=�NA=��@=s�?=%�>=�>=�A==�n<=?�;=O�:=��9=�9=c98=+]7= 6=X�5=��4=��3=M�2=�2=�"1=X60=�G/=�V.=zc-=m,=�t+=�y*=S{)=Wz(=Iv'=Bo&=e%=�W$=	G#=�2"=�!=�  = �=ȿ=ܙ=.p=�B=<=��=��=%e=�#=*�=w�=�F=��=��=PD=��
=E�	=�=��=�B=��=�X=�� =��<���<ث�<q��<�{�<%Y�<~/�<��<���<��<�F�<���<V��<#X�<r��<���<�8�<���<�`�<��<Ew�<���<~�<;��<�v�<��<�c�<�դ<�E�<k��<!�<�<[�<CX�<%��<�"�<)��<��<@�z<�bs<B)l<��d<�]<��V<NO<�H<u�@<�9<	�2<�q+<1Q$<+5<@<<�<�� <_��;��;n1�;Hc�;
��;v��;�a�;�ܓ;�k�;�r;��W;l5=;{#;�	;Cr�:s@�:�p:�2:3`!9*�j�d��k�}������޺v��n3��E5��L�;�b�d�x�����e���)��%̧��L��۬����ƻJѻ<ۻ��仟��05��.� ����$
�²��2������DZ �^�$��(�-�A"1��35��89��1=��A�� E�o�H���L�eP��T���W��n[�|
_��b�J'f�O�i��#m�V�p��t�xfw�>�z��~������\������䟅��=��3و�gr��U	��B���;1��J��Q��Uߓ��k��6�������������b����������d"������$������y%��1���}$�������"��w���T ��3���I��r���������������������  �  kqN=5�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=LAE=�xD=ӯC=��B=�B=�NA=��@=q�?=�>=�>=�A==�n<=<�;=N�:=��9=�9=b98=%]7=%6=W�5=��4=��3=L�2=�2=�"1=[60=�G/=�V.=wc-={m,=�t+=�y*=Z{)=Qz(=Pv'=Ao&=e%=�W$=G#=�2"=�!=�  =��=ɿ=ޙ=+p=�B=<=��=��=#e=�#='�=�=�F=��=��=ND=��
=A�	=�=��=�B=��=�X=�� =��<���<ӫ�<{��<�{�<"Y�<{/�<��<���<t��<�F�<���<^��<X�<j��<���<�8�<���<�`�<��<Aw�<���<~�<9��<w�<��<�c�<�դ<�E�<v��<�<��<X�<AX�<��<#�<*��<��<B�z<�bs<h)l<��d<׸]<��V<NO<�H<_�@<ٿ9<�2<�q+< Q$<75<M<<�<�� <p��;��;r1�;5c�;���;���;�a�;�ܓ;�k�;�r;��W;5=;�#;�	;*s�:@�:��p:@4:�^!9��j���J�}����h�޺���l3�E5��L��b���x����f���)��1̧��L��������ƻѻHۻ��仌��h5��� �����#
�Ѳ��2����	�8Z �_�$���(�3-�E"1��35��89��1=��A�� E�b�H���L�.eP��T���W�o[�q
_��b�0'f�J�i��#m�N�p��t�dfw�Q�z��~�����v\��������=��9و�_r��]	��J���11��J��Q��_ߓ��k��9�������������X��)��������a"������%��x���|%��3����$�������"��|���S ��A���6��z���������������������  �  xqN=-�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=MAE=�xD=ٯC=��B=�B=�NA=��@=x�?= �>=�>=�A==�n<=:�;=U�:=��9=�9=n98="]7='6=P�5=��4=��3=G�2=�2=�"1=^60=�G/=�V.=sc-=m,=�t+=}y*=`{)=Lz(=Sv'=?o&=e%=�W$=G#=3"=!=�  =��=˿=�=(p=�B=2=��=��=%e=�#=%�=��=�F=��=��=QD=��
=<�	=�=��=�B=��=�X=�� =
��<���<ǫ�<���<�{�<7Y�<v/�<���<���<m��<�F�<���<\��<X�<t��<���<�8�< ��<�`�<��<Bw�<���<$~�<,��<w�<��<�c�<�դ<�E�<v��<�<��<G�<XX�<��<�"�<+��<��<N�z<�bs<g)l<w�d<�]<��V<NO<�H<Y�@<�9<�2<�q+<$Q$<35<Z<�<�<�� <���;��;p1�;Cc�;���;���;�a�;�ܓ;�k�;�r;��W;5=;�#;a	;�s�:�?�:��p:�2:�Z!9}{j�Ʊ���}����\�޺����3�UE5�EL�զb���x� �4f���)���˧�4M��z����ƻ�ѻRۻ�����l5��� �����#
�ֲ��2�����Z ���$���(�/-�?"1��35��89��1=��A�� E���H�}�L�eP��T���W�!o[�f
_�*�b�A'f�a�i��#m�E�p��t�Rfw�b�z��~������\�����������=��Dو�`r��\	��@���51��Y��Q��dߓ�vk��8�������������L��,��������^"������%��s����%������$�������"������M ��M���7������������������������  �  qqN=/�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=MAE=�xD=үC=��B=�B=�NA=��@=v�?=!�>=�>=�A==�n<=:�;=U�:=��9=�9=g98="]7=&6=S�5=��4=��3=L�2=�2=�"1=[60=�G/=�V.=tc-=|m,=�t+=y*=]{)=Pz(=Ov'=Bo&=e%=�W$=G#= 3"=�!=�  =��=ǿ=ܙ=)p=�B=7=��=��=$e=�#=)�=}�=�F=��=��=ND=��
=>�	=�=��=�B=��=�X=�� =��<���<̫�<}��<�{�<*Y�<w/�<���<���<q��<�F�<���<`��<X�<t��<���<�8�<���<�`�<��<Bw�<���<&~�<2��<	w�<��<�c�<�դ<�E�<o��<�<��<K�<JX�<��<�"�<,��<��<J�z<�bs<_)l<��d<�]<y�V<NO<�H<X�@<�9<�2<�q+<1Q$<(5<O<<�<�� <���;��;�1�;?c�;���;���;�a�;�ܓ;�k�;�r;ۓW;<5=;�#;�	;%s�:�?�:��p:�2:\!9q�j�Ʊ���}�2��¡޺���t3�JE5��L��b���x�򀇻,f���)�� ̧�#M��������ƻѻ:ۻ��仇��M5��� �΅��#
�ղ��2�����)Z �r�$���(�!-�A"1��35��89��1=��A�� E���H���L�$eP��T���W�o[�q
_��b�;'f�N�i��#m�R�p��t�^fw�b�z��~������\������񟅼�=��:و�]r��Z	��@���11��Q��Q��`ߓ��k��8�������������S��%��������b"�������$��w����%��*����$�������"������O ��<���;��w������Ĝ�������������  �  jqN=6�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=NAE=yD=ӯC=��B=�B=�NA=��@=p�?=#�>=�>=�A==�n<==�;=O�:=��9=�9=_98=+]7="6=Y�5=��4=��3=I�2=2=�"1=X60=�G/=�V.=zc-={m,=�t+=�y*=X{)=Tz(=Mv'=Bo&=e%=�W$=G#=�2"=�!=�  =�=̿=��=2p=�B===��=��=#e=�#=*�={�=�F=��=��=MD=��
=E�	=�=��=�B=��=�X=�� =
��<���<ث�<u��<�{�<Y�<|/�<
��<���<y��<�F�<���<Z��<X�<h��<���<�8�<���<�`�<��<Ow�<���<~�<<��<�v�<��<�c�<�դ<�E�<q��<�<���<\�<>X�<!��< #�<-��<��<3�z<�bs<C)l<��d<ȸ]<��V<'NO<�H<p�@<ҿ9<�2<�q+<,Q$<05<K<<�<�� <a��;��;x1�;Dc�;:��;���;#b�;�ܓ;�k�;�r;s�W;R5=;�#;�	;s�:/@�:5�p:�3:�`!9͉j������}�x��q�޺����3��E5��L�9�b�e�x�����e���)��>̧��L��������ƻ#ѻ;ۻ��仕��Q5��� �����#
�����2������9Z �Z�$���(�)-�H"1��35��89��1=��A�� E�c�H���L�/eP��T���W��n[�{
_��b�T'f�]�i��#m�R�p��t�nfw�?�z��~�����{\������韅��=��6و�cr��Y	��L���41��G��Q��Lߓ��k��,�������������\��$���
�����b"�������$�����x%��7����$�������"��x���[ ��?���I��z���������������������  �  pqN=1�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=NAE=�xD=ͯC=��B=�B=�NA=��@=w�?=$�>=�>=�A==�n<==�;=R�:=��9=�9=e98=(]7= 6=R�5=��4=��3=L�2=�2=�"1=[60=�G/=�V.=vc-=|m,=�t+=�y*=Y{)=Sz(=Ov'=Co&=e%=�W$=G#=3"=�!=�  =��=ſ=ٙ=,p=�B=9=��=��=&e=�#=)�=�=�F=��=��=ND=��
=@�	==��=�B=��=�X=�� =��<���<˫�<r��<�{�<&Y�<v/�<���<���<v��<�F�<���<Y��<%X�<u��<���<�8�<���<�`�<��<>w�<���<!~�<9��<w�<��<�c�<�դ<�E�<p��<�<���<Q�<HX�<��<�"�<!��<��<C�z<�bs<X)l<��d<ܸ]<��V<NO<�H<h�@<�9<��2<�q+<.Q$<-5<X<<�<�� <���;��;x1�;Hc�;���;}��;�a�;�ܓ;�k�;�r;�W;p5=;�#;�	;{s�:.@�:��p:�2:&\!9΃j�E��W�}�F��x�޺���r3�cE5��L��b���x�/���f���)�� ̧�M��������ƻѻ5ۻ���|��>5��� �Å��#
�Ȳ��2�����0Z �h�$���(�-�9"1��35��89��1=��A�� E���H���L�)eP��T���W�o[�q
_��b�A'f�P�i��#m�N�p��t�tfw�I�z��~������\������쟅��=��<و�dr��R	��>���11��L��Q��]ߓ��k��<�������������O��!��������["�������$�������%��,����$�������"��|���S ��:���?��v���������������������  �  rqN=/�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=PAE=�xD=گC=��B=�B=�NA=��@=u�?=�>=�>=�A==�n<=7�;=X�:=��9=�9=i98=]7=(6=V�5=��4=��3=E�2=�2=�"1=Z60=�G/=�V.=tc-=ym,=�t+=y*=`{)=Nz(=Mv'=Eo&=e%=�W$=G#=3"=�!=�  =��=̿=�=,p=�B=3=��=��=!e=�#=*�=~�=�F=��=��=SD=��
==�	=�=��=�B=��=�X=�� =��<���<Ϋ�<���<�{�<+Y�<{/�< ��<���<j��<�F�<���<X��<X�<o��<���<�8�<��<�`�<��<Hw�<���<!~�<.��<w�<��<�c�<�դ<�E�<h��<�<��<L�<NX�<��<#�<-��<��<<�z<�bs<B)l<z�d<׸]<�V< NO<�H<O�@<�9<�2<�q+<6Q$<5<c<�<�<�� <���;��;j1�;Uc�;	��;���;�a�;�ܓ;�k�;�r;̓W;�4=;�#;�	;�s�:u?�:A�p:3:R]!9)�j�O��V�}����ԡ޺����3��E5�L��b���x�倇�%f���)���˧�"M��t��� �ƻ#ѻ"ۻ��代��k5��� �؅��#
�Ʋ��2�����$Z ��$���(�1-�O"1��35��89��1=��A�� E���H�w�L�,eP��T���W�o[�v
_��b�T'f�j�i��#m�W�p��t�Sfw�e�z��~������\�����������=��:و�er��c	��D���51��V��Q��Zߓ�tk��2�������������O��1��������U"������$��s����%��'����$�������"������V ��H���I������������������������  �  pqN=1�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=NAE=�xD=ͯC=��B=�B=�NA=��@=w�?=$�>=�>=�A==�n<==�;=R�:=��9=�9=e98=(]7= 6=R�5=��4=��3=L�2=�2=�"1=[60=�G/=�V.=vc-=|m,=�t+=�y*=Y{)=Sz(=Ov'=Co&=e%=�W$=G#=3"=�!=�  =��=ſ=ٙ=,p=�B=9=��=��=&e=�#=)�=�=�F=��=��=ND=��
=@�	==��=�B=��=�X=�� =��<���<˫�<r��<�{�<&Y�<v/�<���<���<v��<�F�<���<Y��<%X�<u��<���<�8�<���<�`�<��<>w�<���<!~�<9��<w�<��<�c�<�դ<�E�<p��<�<���<Q�<HX�<��<�"�<!��<��<C�z<�bs<X)l<��d<ܸ]<��V<NO<�H<h�@<�9<��2<�q+<.Q$<-5<X<<�<�� <���;��;x1�;Hc�;���;}��;�a�;�ܓ;�k�;�r;�W;p5=;�#;�	;{s�:.@�:��p:�2:"\!9Ӄj�F��X�}�G��y�޺���r3�dE5��L��b���x�/���f���)��!̧�M��������ƻѻ5ۻ���|��>5��� �Å��#
�Ȳ��2�����0Z �h�$���(�-�9"1��35��89��1=��A�� E���H���L�)eP��T���W�o[�q
_��b�A'f�P�i��#m�N�p��t�tfw�I�z��~������\������쟅��=��<و�dr��R	��>���11��L��Q��]ߓ��k��<�������������O��!��������["�������$�������%��,����$�������"��|���S ��:���?��v���������������������  �  jqN=6�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=NAE=yD=ӯC=��B=�B=�NA=��@=p�?=#�>=�>=�A==�n<==�;=O�:=��9=�9=_98=+]7="6=Y�5=��4=��3=I�2=2=�"1=X60=�G/=�V.=zc-={m,=�t+=�y*=X{)=Tz(=Mv'=Bo&=e%=�W$=G#=�2"=�!=�  =�=̿=��=2p=�B===��=��=#e=�#=*�=|�=�F=��=��=MD=��
=E�	=�=��=�B=��=�X=�� =
��<���<ث�<u��<�{�<Y�<|/�<
��<���<y��<�F�<���<Z��<X�<h��<���<�8�<���<�`�<��<Ow�<���<~�<<��<�v�<��<�c�<�դ<�E�<q��<�<���<\�<>X�<!��< #�<-��<��<3�z<�bs<C)l<��d<ȸ]<��V<'NO<�H<p�@<ҿ9<�2<�q+<,Q$<05<K<<�<�� <b��;��;x1�;Dc�;:��;���;#b�;�ܓ;�k�;�r;r�W;Q5=;�#;�	;s�:.@�:3�p:�3:�`!9։j������}�y��r�޺����3��E5��L�:�b�f�x�����e���)��>̧��L��������ƻ$ѻ;ۻ��仕��Q5��� �����#
�����2������9Z �Z�$���(�)-�H"1��35��89��1=��A�� E�c�H���L�/eP��T���W��n[�{
_��b�T'f�]�i��#m�R�p��t�nfw�?�z��~�����{\������韅��=��6و�cr��Y	��L���41��G��Q��Lߓ��k��,�������������\��$���
�����b"�������$�����x%��7����$�������"��x���[ ��?���I��z���������������������  �  qqN=/�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=MAE=�xD=үC=��B=�B=�NA=��@=v�?=!�>=�>=�A==�n<=:�;=U�:=��9=�9=g98="]7=&6=S�5=��4=��3=L�2=�2=�"1=[60=�G/=�V.=tc-=|m,=�t+=y*=]{)=Pz(=Ov'=Bo&=e%=�W$=G#= 3"=�!=�  =��=ǿ=ܙ=)p=�B=7=��=��=$e=�#=)�=}�=�F=��=��=ND=��
=>�	=�=��=�B=��=�X=�� =��<���<̫�<}��<�{�<*Y�<w/�<���<���<q��<�F�<���<`��<X�<t��<���<�8�<���<�`�<��<Bw�<���<&~�<2��<	w�<��<�c�<�դ<�E�<o��<�<��<K�<JX�<��<�"�<,��<��<J�z<�bs<_)l<��d<�]<y�V<NO<�H<X�@<�9<�2<�q+<1Q$<(5<O<<�<�� <���;��;�1�;?c�;���;���;�a�;�ܓ;�k�;�r;ۓW;<5=;�#;�	;$s�:�?�:��p:�2:\!9}�j�ɱ���}�3��ġ޺���u3�KE5��L��b���x�󀇻,f���)�� ̧�$M��������ƻѻ;ۻ��仇��M5��� �΅��#
�ղ��2�����)Z �r�$���(�!-�A"1��35��89��1=��A�� E���H���L�$eP��T���W�o[�q
_��b�;'f�N�i��#m�R�p��t�^fw�b�z��~������\������񟅼�=��:و�]r��Z	��@���11��Q��Q��`ߓ��k��8�������������S��%��������b"�������$��w����%��*����$�������"������O ��<���;��w������Ĝ�������������  �  xqN=-�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=MAE=�xD=ٯC=��B=�B=�NA=��@=x�?= �>=�>=�A==�n<=:�;=U�:=��9=�9=n98="]7='6=P�5=��4=��3=G�2=�2=�"1=^60=�G/=�V.=sc-=m,=�t+=}y*=`{)=Lz(=Sv'=?o&=e%=�W$=G#=3"=!=�  =��=˿=�=(p=�B=2=��=��=%e=�#=%�=��=�F=��=��=QD=��
=<�	=�=��=�B=��=�X=�� =
��<���<ȫ�<���<�{�<7Y�<v/�<���<���<n��<�F�<���<\��<X�<t��<���<�8�< ��<�`�<��<Bw�<���<$~�<,��<w�<��<�c�<�դ<�E�<v��<�<��<G�<XX�<��<�"�<+��<��<N�z<�bs<g)l<w�d<�]<��V<NO<�H<Y�@<�9<�2<�q+<$Q$<35<[<�<�<�� <���;��;p1�;Cc�;���;���;�a�;�ܓ;�k�;�r;��W;5=;�#;a	;�s�:�?�:��p:�2:qZ!9�{j�ʱ���}����^�޺����3�UE5�FL�֦b���x� �4f���)���˧�4M��z����ƻ�ѻRۻ�����l5��� �����#
�ֲ��2�����Z ���$���(�/-�?"1��35��89��1=��A�� E���H�}�L�eP��T���W�!o[�f
_�*�b�A'f�a�i��#m�E�p��t�Rfw�b�z��~������\�����������=��Dو�`r��\	��@���51��Y��Q��dߓ�vk��8�������������L��,��������^"������%��s����%������$�������"������M ��M���7������������������������  �  kqN=5�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=LAE=�xD=ӯC=��B=�B=�NA=��@=q�?=�>=�>=�A==�n<=<�;=N�:=��9=�9=b98=%]7=%6=W�5=��4=��3=L�2=�2=�"1=[60=�G/=�V.=wc-={m,=�t+=�y*=Z{)=Qz(=Pv'=Ao&=e%=�W$=G#=�2"=�!=�  =��=ɿ=ޙ=+p=�B=<=��=��=#e=�#='�=�=�F=��=��=ND=��
=A�	=�=��=�B=��=�X=�� =��<���<ӫ�<{��<�{�<"Y�<{/�<��<���<t��<�F�<���<^��<X�<j��<���<�8�<���<�`�<��<Aw�<���<~�<9��<w�<��<�c�<�դ<�E�<v��<�<��<X�<AX�<��<#�<*��<��<B�z<�bs<h)l<��d<׸]<��V<NO<�H<_�@<ٿ9<�2<�q+< Q$<75<M<<�<�� <q��;��;r1�;5c�;���;���;�a�;�ܓ;�k�;�r;��W;5=;�#;�	;)s�:@�:��p:<4:�^!9�j���N�}����j�޺���m3�E5��L��b���x����f���)��1̧��L��������ƻѻIۻ��仌��i5��� �����#
�Ѳ��2����	�8Z �_�$���(�3-�E"1��35��89��1=��A�� E�b�H���L�.eP��T���W�o[�q
_��b�0'f�J�i��#m�N�p��t�dfw�Q�z��~�����v\��������=��9و�_r��]	��J���11��J��Q��_ߓ��k��9�������������X��)��������a"������%��x���|%��3����$�������"��|���S ��A���6��z���������������������  �  mqN=6�M=��L=�,L=jK=�J=��I=~I=�ZH=��G=��F=�F=NAE=�xD=ͯC=��B=�B=�NA=��@=s�?=%�>=�>=�A==�n<=?�;=O�:=��9=�9=c98=+]7= 6=X�5=��4=��3=M�2=�2=�"1=X60=�G/=�V.=zc-=m,=�t+=�y*=S{)=Wz(=Iv'=Bo&=e%=�W$=	G#=�2"=�!=�  = �=ȿ=ܙ=.p=�B=<=��=��=%e=�#=*�=w�=�F=��=��=PD=��
=E�	=�=��=�B=��=�X=�� =��<���<ث�<q��<�{�<&Y�<~/�<��<���<���<�F�<���<V��<#X�<r��<���<�8�<���<�`�<��<Ew�<���<~�<;��<�v�<��<�c�<�դ<�E�<k��<!�<�<[�<CX�<%��<�"�<)��<��<@�z<�bs<B)l<��d<�]<��V<NO<�H<u�@<�9<	�2<�q+<1Q$<+5<@<<�<�� <_��;��;n1�;Hc�;
��;v��;�a�;�ܓ;�k�;�r;��W;l5=;{#;�	;Br�:q@�:�p:�2:!`!9;�j�h��p�}������޺w��o3��E5��L�<�b�e�x�����e���)��%̧��L��۬����ƻJѻ<ۻ��仟��05��.� ����$
�²��2������DZ �^�$��(�-�A"1��35��89��1=��A�� E�o�H���L�eP��T���W��n[�|
_��b�J'f�O�i��#m�V�p��t�xfw�>�z��~������\������䟅��=��3و�gr��U	��B���;1��J��Q��Uߓ��k��6�������������b����������d"������$������y%��1���}$�������"��w���T ��3���I��r���������������������  �  sqN=2�M=��L=�,L=	jK=�J=��I=|I=�ZH=��G=��F=�F=KAE=�xD=ׯC=��B=�B=�NA=��@=s�?= �>=�>=�A==�n<=:�;=U�:=��9=�9=h98=$]7=&6=W�5=��4=��3=K�2=�2=�"1=Y60=�G/=�V.=uc-=|m,=�t+=�y*=[{)=Qz(=Lv'=Go&=e%=�W$=G#=�2"=�!=�  =��=˿=�=)p=�B=8=��=��=!e=�#=-�=|�=�F=��=��=QD=��
=>�	=�=��=�B=��=�X=�� =��<���<ի�<��<�{�<,Y�<~/�<��<���<t��<�F�<���<T��<X�<p��<���<�8�<���<�`�<��<Cw�<���<~�<8��<w�<��<�c�<�դ<�E�<g��<�<���<U�<OX�<��<�"�</��<��<:�z<�bs<\)l<��d<ظ]<��V<$NO<�H<Z�@<��9<��2<�q+<7Q$<5<_<<�<�� <}��;��;d1�;/c�;���;���;�a�;�ܓ;�k�;�r;��W;$5=;g#;�	;(s�:�?�:��p:�2:�^!9 �j�1����}����}�޺����3�UE5��L�%�b�b�x�����'f���)��̧�M��������ƻ2ѻۻ��仮��S5��� �Ņ��#
�ڲ��2�����:Z �n�$���(�(-�O"1��35��89��1=��A�� E�y�H�~�L�$eP��T���W��n[�r
_��b�;'f�P�i��#m�M�p��t�]fw�Y�z��~������\������🅼�=��5و�ir��^	��E���81��S��Q��`ߓ�zk��7�������������Z��'��������V"������$��z���%��%����$�������"��w���W ��;���=��x���������������������  �  rqN=.�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=OAE=�xD=կC=��B=�B=�NA=��@=p�?=!�>=�>=�A==�n<=7�;=V�:=��9=�9=h98=#]7=,6=P�5=��4=��3=L�2=�2=�"1=a60=�G/=�V.=xc-=}m,=�t+=y*=_{)=Mz(=Sv'=>o&=e%=�W$= G#=3"=�!=�  =��=ſ=ܙ=%p=�B=4=��=~�=(e=�#=$�=��=�F=��=��=QD=��
=@�	=�=��=�B=��=�X=�� =��<ĸ�<ƫ�<���<�{�</Y�<y/�<��<���<l��<�F�<���<c��< X�<h��<���<�8�<���<�`�<��<7w�<���<~�<,��<w�<��<�c�<�դ<�E�<r��<�<��<I�<MX�<��<#�<&��<��<R�z<�bs<t)l<��d<�]<��V<NO<H<Z�@<��9<�2<�q+<2Q$<(5<V<�<�<�� <t��;��;_1�;Hc�;ƥ�;���;�a�;�ܓ;�k�;�r;i�W;15=;#;?	;�s�:d?�:��p:�2:�Z!9��j������}������޺���r3�E5�L���b���x�����	f���)��̧�)M��}���	�ƻ�ѻ\ۻ���d��t5��� �څ��#
����2�����.Z ��$���(�;-�5"1��35��89��1=��A�� E���H���L� eP��T���W�(o[�W
_��b�*'f�F�i��#m�6�p��t�Ifw�]�z��~������\�����������=��Hو�Zr��X	��M���/1��Z��Q��lߓ�k��D�������������V��-���������`"�������$��r����%��(����$�������"�����L ��A���1��z���������������������  �  qqN=4�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=NAE=�xD=ԯC=��B=�B=�NA=��@=p�?= �>=�>=�A==�n<=<�;=S�:=��9=�9=h98=&]7=(6=S�5=��4=��3=K�2=�2=�"1=^60=�G/=�V.=yc-=}m,=�t+=�y*=Z{)=Pz(=Qv'=?o&=e%=�W$= G#=�2"=�!=�  =��=ɿ=ޙ=+p=�B=5=��=�=$e=�#=%�=��=�F=��=��=SD=��
=C�	=�=��=�B=��=�X=�� =��<���<ϫ�<���<�{�</Y�<~/�<��<���<s��<�F�<���<Y��<X�<i��<���<�8�<���<�`�<��<Bw�<���<~�<3��<w�<��<�c�<�դ<�E�<s��<�<���<V�<MX�<��<#�<*��<��<J�z<�bs<V)l<��d<�]<��V<NO<�H<f�@<�9<�2<�q+<(Q$<05<S<�<�<�� <s��;��;F1�;Dc�;���;���;�a�;�ܓ;xk�;�r;s�W;5=;�#;f	;Rs�:�?�:��p:�2:�^!9z�j�۰�b�}�:���޺����3�yE5��L�ܦb���x��f���)��̧�M��������ƻѻ[ۻ��仔��u5��� �҅��#
�ϲ��2�����9Z �z�$���(�5-�F"1��35��89��1=��A�� E�s�H�w�L�eP��T���W�o[�a
_��b�E'f�S�i��#m�=�p��t�Tfw�O�z��~������\������🅼�=��Bو�dr��^	��K���21��Y��Q��^ߓ��k��8�������������X��-��������a"������%��z���~%��(����$�������"��x���O ��=���@��w���������������������  �  oqN=5�M=��L=�,L=jK=�J=��I={I=�ZH=��G=��F=�F=HAE=�xD=ͯC=��B=�B=�NA=��@=t�?="�>=�>=�A==�n<=>�;=S�:=��9=�9=f98=']7=$6=X�5=��4=��3=Q�2=�2=�"1=Z60=�G/=�V.=tc-=}m,=�t+=�y*=Y{)=Tz(=Lv'=Eo&=e%=�W$=	G#=�2"=�!=�  =��=Ŀ=ٙ=)p=�B=<=��=��= e=�#=-�=|�=�F=��=��=PD=��
=A�	=�=��=�B=��=�X=�� =��<���<ګ�<{��<�{�<+Y�<}/�<��<���<{��<�F�<��<P��<X�<u��<���<�8�<���<�`�<��<>w�<���<~�<=��<�v�<��<�c�<�դ<�E�<i��<�<���<X�<HX�<!��<�"�<-��<��<?�z<�bs<Z)l<��d<ݸ]<��V<%NO<�H<h�@<�9<�2<�q+<2Q$<&5<Q<<�<�� <f��;��;j1�;c�;�;x��;�a�;|ܓ;�k�;�r;��W;65=;@#;�	;�r�:B@�:��p:�2:�^!9��j������}������޺v��'3�UE5�RL��b�Y�x�����(f���)��̧��L��������ƻ2ѻ%ۻ������05��#� �����#
�ݲ��2�����BZ �]�$��(�-�U"1��35��89��1=��A�� E�n�H���L�%eP��T���W��n[�r
_��b�6'f�=�i�#m�T�p��t�efw�O�z��~������\������韅��=��0و�nr��\	��@���81��K��Q��cߓ��k��<�������������^����������["������$��}���|%��,����$�������"��s���U ��*���>��g���������������������  �  rqN=0�M=��L=�,L=jK=�J=��I=�I=�ZH=��G=��F=�F=MAE=�xD=үC=��B=�B=�NA=��@=p�?=!�>=�>=�A==�n<==�;=R�:=��9=�9=i98=(]7=*6=W�5=��4=��3=I�2=2=�"1=]60=�G/=�V.=zc-=�m,=�t+=�y*=]{)=Sz(=Nv'=>o&=e%=�W$=G#=�2"=�!=�  =��=ȿ=ݙ=-p=�B=7=��=��="e=�#=%�=~�=�F=��=��=OD=��
=D�	=�=��=�B=��=�X=�� =��<���<ի�<���<�{�<0Y�<z/�<	��<���<x��<�F�<���<X��<X�<l��<���<�8�<���<�`�<��<Cw�<���<~�</��<�v�<��<�c�<�դ<�E�<o��<�<��<P�<JX�<$��<#�<0��<��<E�z<�bs<G)l<��d<�]<��V<(NO<�H<n�@<�9<�2<�q+</Q$<,5<G<<�<�� <J��;��;g1�;;c�;���;���;�a�;�ܓ;�k�;Br;l�W;35=;�#;�	;�r�:@�:��p:|3:�[!9׀j�c����}����b�޺����3��E5��L��b���x������e���)��!̧�M��������ƻ ѻ]ۻ��仡��G5��*� �҅��#
�ʲ��2�����:Z �s�$��(�&-�K"1��35��89��1=��A�� E�t�H���L�eP��T���W�
o[�g
_��b�Q'f�]�i��#m�J�p��t�Nfw�G�z��~�����~\������쟅��=��>و�er��[	��I���A1��S��Q��]ߓ��k��8�������������d��"��������d"�������$��v����%��*���~$�������"��v���R ��:���G��x���������������������  �  'tN=H�M=!�L=�0L=�nK=��J=��I=c%I=0aH=g�G=��F=�F=�IE=�D=]�C=��B=`%B=�YA=w�@=�?=5�>=P!>=)P==�}<=��;=��:=�9=�%9=L8=xp7=K�6=9�5=U�4={�3=�3=�$2=�;1=2P0=rb/=ir.=�-=��,=��+=o�*=$�)=�(=Ɨ'=��&=*�%=�{$=�k#=mX"=�A!=k' =�	=��=��=��=�l=�;=�=��=��=�O=<
=��=s=2!=�=�p="=J�	=[H=$�=�m=q�=�=�=�<|	�<��<S��<���<���<1x�<�E�<��<V��<���<�;�<���<{��<�5�<e��<'l�<& �<s��<��<F��<-$�<O��<��<d��<��<!�<��<`\�<�ǝ<�0�<R��<4��<�b�<Ƌ<�(�<d��<��<6�z<�Zs<�l<��d<��]<ZgV<'.O<5�G<��@<�9<�c2< :+<�$<��<*�<�<�<]� <hK�;+T�;ll�;��;~λ;Z�;$x�;-�;Tp�;�p;�zU;�;;�� ;e�;1��:Qo�:jg:�!:���8�,��K\'�;T��8���J4���	��!�|&8���N���e�s�{�@����ᓻ"���pH��}ɳ�U(���eȻ�һu{ܻFT�E�ѣ��^��9��
��a����M�Ŭ��� � A%�yv)���-�J�1�U�5���9�J�=�#�A�H�E��YI��!M��P�9�T�J>X�n�[�w_�ec��f��j���m��p�fZt���w��{��j~��܀�����"�������]��'���菊��%��1����J���ڐ��h��v���[���
��:���?������#�������*�������-�������.��)���M-��𫪼�*�������&��ᤰ��"��砳����g������𚹼@�����o���  �  tN=C�M=�L=�0L=�nK=�J=��I=c%I=5aH=c�G=��F=�F=�IE=�D=V�C=��B=_%B=�YA=w�@=�?=5�>=S!>=4P==�}<=��;=��:=�9=�%9=L8=�p7=I�6=:�5=W�4=z�3=�3=�$2=�;1=,P0=wb/=fr.=�-=��,=�+=k�*=!�)=�(=Ǘ'=��&=/�%=�{$=�k#=jX"=�A!=k' =�	=��=��=��=�l=�;=�=��=��=�O=E
=��=s=/!=�=�p= =R�	=WH=(�=�m=p�=��== �<{	�<��<M��<��<���<"x�<�E�<��<`��<���<�;�<���<{��<�5�<e��<-l�<% �<}��<~�<J��<0$�<T��< �<]��<��<"�<��<h\�<�ǝ<�0�<P��<)��<�b�<*Ƌ<�(�<`��<��<�z<�Zs<�l<��d<��]<dgV< .O<8�G<��@<��9<�c2<:+<�$<��<0�<*�<�<q� <IK�;BT�;l�;
��;�λ;#�;Cx�;$�;ap�;�p;�zU;�;;�� ;�;���:�o�:�g:�!:ly�8w3��Z'�vT�����4���	� !��&8���N��e��{�\����ᓻ����H���ɳ�h(���eȻ�һ2{ܻT�7𻘣��l��	9��
�}a����
M������ �A%��v)�i�-�A�1�?�5���9�S�=��A�T�E��YI�"M��P��T�]>X�]�[�-w_�lc��f��j���m��p�ZZt���w�~{��j~��܀�����"������^�����⏊��%��-����J���ڐ��h��l���f��� 
��7���;������#�������*�������-�������.��,���X-������*�������&��٤���"��砳���j������뚹�C�����_���  �  tN=R�M=�L=�0L=�nK=��J=��I=^%I=9aH=_�G=��F=�F=�IE=�D=P�C=��B=\%B=�YA=u�@=�?=8�>=P!>=5P==�}<=��;=��:=�9=�%9=�K8=�p7=C�6==�5=U�4=y�3=�3=�$2=�;1=&P0=}b/=`r.=�-=��,=�+=v�*=�)=�(=��'=��&=,�%=�{$=�k#=eX"=�A!=g' =�	=��=��=��=�l=�;=�=��=��=�O=D
=��=s=,!=�=�p==R�	=PH=-�=�m=t�=��=�=!�<v	�<$��<@��<��<���<7x�<�E�<��<c��<���<�;�<���<|��<�5�<^��<+l�< �<���<r�<N��<+$�<O��< �<R��<��<�<��<[\�<�ǝ<�0�<N��<D��<�b�<1Ƌ<�(�<]��<��<�z<�Zs<�l<�d<p�]<mgV<!.O<"�G<��@<��9<d2<:+<�$<��<�<+�< �<�� <(K�;>T�;ql�;���;�λ;��;\x�;
�;Sp�;�p;�zU;�;;�� ;�;���:�o�: g:�":*��8�5��Y'�8U������Q4��	��!��&8�v�N�C�e���{������ᓻ����H��Bɳ�|(���eȻJ�һJ{ܻ/T�P𻂣��}��9��
��a����M����� �A%��v)�d�-�L�1�M�5���9�u�=��A�a�E�jYI��!M��P��T�y>X�G�[�?w_�Yc��f��j���m��p�JZt���w�p{��j~��܀������"������^�����鏊��%��-����J���ڐ��h��f���r����	��<���@������#�������*�������-�������.��-���=-�����|*��Ǩ���&��Ѥ���"��٠����]�����皹�C�����V���  �  tN=H�M=�L=�0L=�nK= �J=��I=a%I=5aH=b�G=��F=�F=�IE=�D=V�C=��B=b%B=�YA=v�@=�?=8�>=Q!>=1P==�}<=��;=��:=�9=�%9=L8=�p7=G�6=>�5=R�4=w�3=�3=�$2=�;1=&P0=xb/=dr.=�-=��,=�+=k�*=�)=�(=Ɨ'=��&=/�%=�{$=�k#=kX"=�A!=m' =�	=��=��=��=�l=�;=�=��=��=�O=D
=��=s=+!=	�=�p==O�	=SH=)�=�m=r�=��=�=�<r	�< ��<H��<��<���<,x�<�E�<��<c��<���<�;�<���<���<�5�<c��<.l�<) �<���<|�<N��<2$�<X��<��<Z��<��< �<��<b\�<�ǝ<�0�<A��<0��<�b�<%Ƌ<�(�<f��<��<�z<�Zs<|l<��d<n�]<_gV<0.O<&�G<��@<��9<�c2<�9+<�$<��<*�<)�<�<s� <>K�;4T�;�l�; ��;�λ;!�;Xx�;=�;bp�;�p;�zU;�;;�� ;�;���:p�:?g:�:3��8�3��,Z'��T�������4�0�	��!�'8���N�<�e��{�j����ᓻ)����H���ɳ��(���eȻ�һ@{ܻT�/𻪣��h��9���
�|a����M������ �A%�v)�u�-�9�1�C�5���9�P�=��A�g�E��YI�"M��P�#�T�h>X�Y�[�@w_�`c��f��j���m��p�SZt���w��{��j~��܀�����"������ ^�����揊��%��0����J���ڐ��h��f���h����	��6���7������#�������*�������-�������.��;���Q-������*��Ũ���&��٤���"��ߠ����`������;�����b���  �  tN=E�M="�L=�0L=~nK= �J=��I=d%I=2aH=h�G=��F=�F=�IE=�D=W�C=��B=a%B=�YA={�@=�?=5�>=S!>=-P==�}<=�;=��:=�9=�%9=L8=~p7=I�6=9�5=W�4=z�3=�3=�$2=�;1=.P0=xb/=fr.=�-=��,=�+=l�*=*�)=�(=ė'=��&=*�%=�{$=�k#=qX"=�A!=o' =�	=��=��=��=�l=�;=�=��=��=�O=@
=��=s=8!=�=�p==R�	=WH='�=�m=q�=��==�<{	�<��<O��<��<���<*x�<�E�<��<R��<���<�;�<���<|��<�5�<l��<'l�<( �<x��<~�<F��<1$�<[��<��<g��<��<'�<��<b\�<�ǝ<�0�<Z��<)��<�b�< Ƌ<�(�<a��<��<"�z<�Zs<�l<��d<��]<dgV<".O<0�G<��@<��9<�c2<":+<�$<��<-�<�<�<i� <mK�;JT�;�l�;��;uλ;/�;-x�;5�;Qp�;�p;�zU;�;;�� ;��;7��:�n�:�g:F":���8�2���Z'��T��#���4��	��!��&8���N���e��{�W����ᓻ0����H���ɳ�"(���eȻ �һV{ܻFT�+𻻣��O��9���
�ya����M������ �(A%�hv)�z�-�:�1�P�5���9�V�=��A�0�E��YI�"M��P��T�X>X�_�[�"w_�gc��f��j���m��p�aZt���w��{��j~��܀�����"�������]�����䏊��%��0����J���ڐ��h��q���f���
��6���3������#������|*�������-�������.��"���X-��	����*�������&��٤���"��⠳���d������뚹�B��	���g���  �  tN=L�M=�L=�0L=�nK=�J=��I=d%I=5aH=d�G=��F=�F=�IE=��D=V�C=��B=b%B=�YA=x�@=�?=6�>=S!>=3P==�}<=��;=��:=�9=�%9= L8=�p7=E�6=9�5=T�4=y�3=�3=�$2=�;1=&P0=xb/=_r.=�-=��,=�+=q�*= �)=�(=ŗ'=��&=+�%=�{$=�k#=mX"=�A!=k' =�	=��=��=��=�l=�;=�=��=��=�O=F
=��=s=-!=�=�p==Q�	=PH=(�=�m=r�=��=}=�<t	�<��<C��<��<���<1x�<�E�<��<W��<���<�;�<���<y��<�5�<f��<)l�<' �<���<|�<P��<1$�<R��< �<^��<��<%�<��<o\�<�ǝ<�0�<M��<7��<�b�<'Ƌ<�(�<Y��<��<	�z<�Zs<�l<��d<q�]<bgV<.O<,�G<��@<��9<�c2<:+<|$<��<=�<!�<�<r� <MK�;DT�;zl�;��;�λ;&�;lx�;<�;Xp�;�p;�zU;�;;�� ;�;?��:�o�:g:Z!:���8u4���Y'��T��5���h4��	�!��&8���N�3�e��{������ᓻ;����H��oɳ�r(���eȻ�һ{ܻ=T�8𻚣��_��9��
�pa����M������ �A%�wv)�k�-�E�1�P�5���9�T�=��A�Z�E��YI��!M��P��T�t>X�]�[�;w_�bc�$�f��j���m��p�_Zt���w�w{��j~��܀�����"�������]�����䏊��%��+����J���ڐ��h��b���i����	��6���=������#������~*�������-�������.��.���J-������*�������&��ؤ���"��⠳���d��� ��욹�H��
���_���  �  tN=J�M=�L=�0L=�nK=��J=��I=`%I=9aH=d�G=��F=�F=�IE=��D=Q�C=��B=^%B=�YA=v�@=�?=8�>=O!>=2P==�}<=��;=��:=�9=�%9=�K8=�p7=B�6=<�5=O�4=z�3=�3=�$2=�;1=$P0=zb/=_r.=�-=��,=�+=m�*=�)=��(=��'=��&=,�%=�{$=�k#=iX"=�A!=i' =�	=��=��=��=�l=�;=�=��=��=�O=B
=��= s=*!=�=�p==T�	=OH=+�=�m=u�=��=}=!�<i	�<!��<=��<��<���<*x�<�E�<��<n��<���<�;�<���<~��<�5�<`��<3l�<  �<���<u�<Q��<3$�<S��<�<\��<��<�<��<^\�<�ǝ<�0�<E��<4��<�b�<+Ƌ<�(�<Z��<��<�z<�Zs<ml<��d<k�]<WgV<.O<$�G<��@<��9<�c2<�9+<�$<��<�<#�<�<�� <OK�;CT�;�l�;��;�λ;��;vx�;#�;yp�;�p;{U;�;;�� ;��;[��:�p�:�g:� :���8�5���X'�EU������5���	��!�O'8�c�N�Y�e���{������ᓻ/����H���ɳ��(��GeȻ3�һF{ܻ4T�H�q���m���8�	�
�ia����M������ �A%��v)�Y�-�I�1�N�5���9�g�=��A�g�E��YI�"M��P��T�z>X�P�[�Kw_�Tc�1�f��j���m�'�p�OZt�»w�j{�k~��܀�
����"��}���^�����돊��%��#����J���ڐ��h��^���p����	��4���;������#�������*�������-�������.��6���M-������*��¨���&��ڤ���"��ݠ����`�����򚹼E�����Z���  �  tN=I�M=!�L=�0L=~nK= �J=��I=e%I=7aH=g�G=��F=�F=�IE=�D=X�C=��B=`%B=�YA=u�@=�?=7�>=U!>=3P==�}<=��;=��:=�9=�%9=L8=�p7=D�6=:�5=N�4=x�3=�3=�$2=�;1='P0=ub/=br.=�-=��,=�+=q�*="�)=�(='=��&=/�%=�{$=�k#=mX"=�A!=n' =�	=��=��=��=�l=�;=�=��=��=�O=E
=��=s=/!=�=�p==P�	=RH=&�=�m=s�=��=|=�<k	�<��<C��<��<���<'x�<�E�<��<U��<���<�;�<���<z��<�5�<_��<0l�<% �<���<��<N��<3$�<]��<��<a��<��<$�< �<d\�<�ǝ<�0�<S��<5��<�b�<$Ƌ<�(�<]��<��<�z<�Zs<�l<��d<s�]<PgV<.O<"�G<��@<��9<�c2<:+<�$<��<,�<.�<�<{� <dK�;5T�;�l�;��;�λ;6�;bx�;0�;{p�;�p;{U;�;;�� ;�;���:Xo�:�g:�":���854���Y'�U������5��	��!�'8���N�$�e�1�{�t����ᓻ>����H��mɳ�^(���eȻ0�һ1{ܻT�;𻉣��`��9���
�ua����	M������ �A%�{v)�e�-�E�1�<�5���9�]�=��A�S�E�YI�"M� �P��T�l>X�`�[�=w_�\c�*�f��j���m�$�p�\Zt���w�{��j~��܀������"������^����������%��(����J���ڐ��h��e���d����	��5���1������#������*�������-�������.��)���K-������*��ƨ���&��ᤰ��"��ߠ��
��c����������C�����c���  �  tN=E�M=�L=�0L=�nK=�J=��I=h%I=2aH=h�G=��F=�F=�IE=��D=X�C=��B=g%B=�YA=z�@=�?=5�>=V!>=-P==�}<=��;=��:=�9=�%9=L8=}p7=I�6=8�5=T�4=x�3=�3=�$2=�;1=(P0=sb/=er.=�-=��,=�+=j�*=#�)=�(=͗'=��&=,�%=�{$=�k#=rX"=�A!=r' =�	=��=��=��=�l=�;=�=��=��=�O=C
=��=s=/!=	�=�p==L�	=UH="�=�m=n�=��={=�<t	�<��<K��<��<���<$x�<�E�<��<Y��<���<�;�<���<z��<�5�<l��</l�<3 �<���<��<R��<6$�<a��<��<g��<��<,�<��<m\�<�ǝ<�0�<R��<*��<�b�< Ƌ<�(�<c��<��<
�z<�Zs<�l<��d<p�]<VgV<$.O<,�G<��@<��9<�c2<:+<{$<��<=�<�<&�<h� <mK�;JT�;�l�;:��;�λ;7�;cx�;h�;yp�;�p;{U;�;;� ;��;���:�o�:�g:-!:��8f3���Z'�eT��5���_4��	�+!�'8���N��e�X�{�\����ᓻ/����H���ɳ�Z(���eȻ׀һ0{ܻ3T�𻗣��I��9���
�wa����M������ �A%�bv)�e�-�5�1�G�5���9�2�=�!�A�R�E��YI�
"M��P�,�T�^>X�p�[�5w_�pc�&�f��j���m��p�mZt���w��{��j~��܀�����"�������]����������%��$����J���ڐ��h��f���b����	��2���-������#������x*�������-��~����.��)���W-������*��Ĩ���&��ᤰ��"��𠳼��s��� ��򚹼A��
���g���  �  tN=K�M=�L=�0L=�nK=��J=��I=f%I=5aH=e�G=��F=�F=�IE=��D=T�C=��B=_%B=�YA={�@=�?=7�>=V!>=/P==�}<=��;=��:=�9=�%9=�K8=p7=B�6=8�5=R�4=x�3=�3=�$2=�;1=(P0=wb/=`r.=�-=��,=�+=n�*="�)=�(=��'=��&=,�%=�{$=�k#=nX"=�A!=m' =�	= �=��=��=�l=�;=�=��=��=�O=>
=��=s=0!=�=�p==L�	=PH=&�=�m=p�=��=|=�<o	�<��<?��<��<���<0x�<�E�<��<`��<���<�;�<���<~��<�5�<i��<0l�<$ �<���<|�<V��<.$�<Y��<�<c��<��<(�<��<Y\�<�ǝ<�0�<O��<3��<�b�<(Ƌ<�(�<Z��<��<�z<�Zs<l<��d<u�]<UgV<.O<�G<��@<��9<�c2<:+<�$<��<�<!�<!�<t� <]K�;hT�;�l�;��;�λ;�;lx�;-�;zp�;p;�zU;�;;� ;ؼ;;��:�o�:�g:)!:��8�4��FZ'�8U��.����4��	��!�'8���N��e��{������ᓻ����H���ɳ�[(��{eȻ<�һg{ܻ/T�.𻜣��Z��9���
�ta�����L������ �A%�rv)�o�-�?�1�H�5���9�h�=��A�M�E��YI�"M��P�)�T�t>X�`�[�:w_�fc�*�f��j���m��p�bZt���w��{��j~��܀�����"������^�����Ꮚ��%��+����J���ڐ��h��e���h����	��9���5������#������|*�������-�������.��,���N-������*��ɨ���&��ߤ���"��䠳���h������򚹼G�����`���  �  tN=L�M=�L=�0L=�nK=�J=�I=a%I=;aH=d�G=��F=�F=�IE=��D=Z�C=��B=_%B=�YA=w�@=�?=<�>=Q!>=:P==�}<=��;=��:=�9=�%9=�K8=�p7=>�6=;�5=M�4=u�3=�3=�$2=�;1="P0=vb/=]r.=�-=��,=�+=p�*=�)=�(=��'=��&=1�%=�{$=�k#=jX"=�A!=n' =�	= �=��=��=�l=�;=�=��=��=�O=J
=��=s=&!=�=�p==P�	=KH=&�=�m=p�=��={=�<d	�<��<3��<��<���<+x�<�E�<��<\��<���<�;�<���<���<�5�<a��<9l�<# �<���<��<W��<2$�<_��<�<]��<��<�<	�<n\�<�ǝ<�0�<=��<:��<�b�<)Ƌ<�(�<Y��<��<��z<�Zs<gl<��d<b�]<KgV<.O<�G<��@<��9<�c2<�9+<�$<��<5�<D�<�<�� <PK�;KT�;�l�;��;�λ;I�;�x�;+�;�p�;�p;�zU;;;�� ;��;���:�o�:�g:� :l��8�6���X'��U��ڂ��B5�D�	�!�X'8���N�x�e�'�{������ᓻ7����H��oɳ��(��zeȻ4�һ{ܻT�.�~���i���8���
�la�����L������ ��@%��v)�a�-�6�1�>�5���9�b�=��A�v�E��YI�"M�#�P��T��>X�^�[�Uw_�fc�3�f��j���m�0�p�WZt�Իw�q{�k~��܀�����"������^�����珊��%��*����J���ڐ��h��^���_����	��6���/��
����#�������*�������-�������.��?���G-������*��ʨ���&��⤰��"��⠳���e���������E�����[���  �  tN=K�M=�L=�0L=�nK=�J=��I=e%I=6aH=j�G=��F=�F=�IE=�D=Z�C=��B=e%B=�YA=z�@=�?=9�>=Q!>=-P==�}<=��;=��:=�9=�%9= L8=�p7=C�6=;�5=O�4=x�3=�3=�$2=�;1=&P0=wb/=ar.=�-=��,=�+=o�*=!�)=�(=ŗ'=��&='�%=�{$=�k#=pX"=�A!=q' =�	=��=��=��=�l=�;=�=��=��=�O=A
=��=s=/!=�=�p==P�	=OH='�=�m=n�=��={=�<k	�<��<<��<��<���</x�<�E�<��<[��<���<�;�<���<���<�5�<k��<.l�</ �<}��<��<N��<7$�<a��<��<h��<��<(�<��<f\�<�ǝ<�0�<N��<8��<�b�<"Ƌ<�(�<]��<��<�z<�Zs<�l<��d<h�]<RgV<.O<�G<��@<��9<�c2<:+<�$<��<1�<�<�<x� <~K�;FT�;�l�;9��;�λ;H�;Ox�;[�;xp�;�p;8{U;�;;�� ;��;��:�o�:�g:�!:��8�4���Y'�"U��ゴ��4��	�!�'8���N�0�e��{�z����ᓻ2����H��vɳ�e(���eȻ�һG{ܻTT�𻕣��P��	9���
�ta�����L������ �A%�hv)�f�-�.�1�[�5���9�U�=��A�R�E��YI��!M��P��T�t>X�]�[�Bw_�mc�$�f��j���m�!�p�ZZt�»w�}{��j~��܀�����"������ ^�����쏊��%��#����J���ڐ��h��k���^����	��1���-������#������{*�������-�������.��-���H-������*��ɨ���&��ޤ���"��頳���k�����󚹼D�����c���  �  tN=C�M=�L=�0L=�nK=�J=��I=u%I=-aH=j�G=��F=�F=�IE=�D=_�C=��B=l%B=�YA={�@=�?=4�>=c!>=3P==�}<=�;=��:=�9=�%9=�K8=yp7=G�6=8�5=N�4=u�3=�3=�$2=|;1='P0=tb/=ar.=�-=��,=�+=e�*=%�)=�(=Ɨ'=��&=0�%=�{$=�k#=tX"=�A!=s' =�	=�=��=��=�l=�;=�=��=��=�O=D
=��=s=2!=�=�p==J�	=PH=$�=�m=i�=��=z=�<j	�<��<D��<���<���<$x�<�E�<��<N��<���<�;�<��<|��<�5�<p��<#l�<< �<}��<��<P��<:$�<^��<��<l��<��<F�<��<l\�<�ǝ<�0�<S��<$��<�b�<"Ƌ<�(�<Z��<��<�z<�Zs<�l<��d<m�]<LgV<.O<,�G<��@<��9<�c2<:+<�$<��<?�< �<Z�<V� <}K�;MT�;�l�;\��;�λ;p�;Nx�;��;Up�;p;�zU;�;;�� ;�;?��:o�:�g:� :�8�4���['��T��I���"5�?�	�<!��&8�(�N�(�e�F�{�v����ᓻ8����H���ɳ�D(���eȻ�һ4{ܻT���ԣ��@��9���
�sa�����L������ �#A%�Tv)���-�!�1�.�5���9�K�=�!�A�F�E��YI�"M�$�P�2�T�p>X�i�[�@w_��c��f��j���m�$�p�fZt���w��{��j~��܀�����"�������]�����ɏ���%��/����J���ڐ��h��k���T����	��-���0������#������^*�������-�������.��)���]-������*��Ĩ���&��ᤰ��"��𠳼���p���������I��
���j���  �  tN=K�M=�L=�0L=�nK=�J=��I=e%I=6aH=j�G=��F=�F=�IE=�D=Z�C=��B=e%B=�YA=z�@=�?=9�>=Q!>=-P==�}<=��;=��:=�9=�%9= L8=�p7=C�6=;�5=O�4=x�3=�3=�$2=�;1=&P0=wb/=ar.=�-=��,=�+=o�*=!�)=�(=ŗ'=��&='�%=�{$=�k#=pX"=�A!=q' =�	=��=��=��=�l=�;=�=��=��=�O=A
=��=s=/!=�=�p==P�	=OH='�=�m=n�=��={=�<k	�<��<<��<��<���</x�<�E�<��<[��<���<�;�<���<���<�5�<k��<.l�</ �<}��<��<N��<7$�<a��<��<h��<��<(�<��<f\�<�ǝ<�0�<N��<8��<�b�<"Ƌ<�(�<]��<��<�z<�Zs<�l<��d<h�]<RgV<.O<�G<��@<��9<�c2<:+<�$<��<1�<�<�<x� <~K�;FT�;�l�;9��;�λ;H�;Ox�;[�;xp�;�p;8{U;�;;�� ;��;��:�o�:�g:�!:t��8�4���Y'�#U��ゴ��4��	�!�'8���N�0�e��{�z����ᓻ2����H��vɳ�e(���eȻ�һG{ܻTT�𻕣��P��	9���
�ta�����L������ �A%�hv)�f�-�.�1�[�5���9�U�=��A�R�E��YI��!M��P��T�t>X�]�[�Bw_�mc�$�f��j���m�!�p�ZZt�»w�}{��j~��܀�����"������ ^�����쏊��%��#����J���ڐ��h��k���^����	��1���-������#������{*�������-�������.��-���H-������*��ɨ���&��ޤ���"��頳���k�����󚹼D�����c���  �  tN=L�M=�L=�0L=�nK=�J=�I=a%I=;aH=d�G=��F=�F=�IE=��D=Z�C=��B=_%B=�YA=w�@=�?=<�>=Q!>=:P==�}<=��;=��:=�9=�%9=�K8=�p7=>�6=;�5=M�4=u�3=�3=�$2=�;1="P0=vb/=]r.=�-=��,=�+=p�*=�)=�(=��'=��&=1�%=�{$=�k#=jX"=�A!=n' =�	= �=��=��=�l=�;=�=��=��=�O=J
=��=s=&!=�=�p==P�	=KH=&�=�m=p�=��=|=�<d	�<��<3��<��<���<+x�<�E�<��<]��<���<�;�<���<���<�5�<a��<9l�<# �<���<��<W��<2$�<_��<�<]��<��<�<	�<n\�<�ǝ<�0�<=��<:��<�b�<)Ƌ<�(�<Y��<��<��z<�Zs<gl<��d<b�]<KgV<.O<�G<��@<��9<�c2<�9+<�$<��<5�<D�<�<�� <PK�;KT�;�l�;��;�λ;I�;�x�;+�;�p�;�p;�zU;;;�� ;��;���:�o�:�g:� :U��8�6���X'��U��ۂ��C5�E�	�!�Y'8���N�x�e�'�{������ᓻ7����H��oɳ��(��zeȻ4�һ{ܻT�/�~���i���8���
�la�����L������ ��@%��v)�a�-�6�1�>�5���9�b�=��A�v�E��YI�"M�#�P��T��>X�_�[�Uw_�fc�3�f��j���m�0�p�WZt�Իw�q{�k~��܀�����"������^�����珊��%��*����J���ڐ��h��^���_����	��6���/��
����#�������*�������-�������.��?���G-������*��ʨ���&��⤰��"��⠳���e���������E�����[���  �  tN=K�M=�L=�0L=�nK=��J=��I=f%I=5aH=e�G=��F=�F=�IE=��D=T�C=��B=_%B=�YA={�@=�?=7�>=V!>=/P==�}<=��;=��:=�9=�%9=�K8=p7=B�6=8�5=R�4=x�3=�3=�$2=�;1=(P0=wb/=`r.=�-=��,=�+=n�*="�)=�(=��'=��&=,�%=�{$=�k#=nX"=�A!=m' =�	= �=��=��=�l=�;=�=��=��=�O=>
=��=s=0!=�=�p==L�	=PH=&�=�m=p�=��=|=�<o	�<��<?��<��<���<0x�<�E�<��<`��<���<�;�<���<~��<�5�<i��<0l�<$ �<���<|�<V��<.$�<Y��<�<c��<��<'�<��<Y\�<�ǝ<�0�<O��<3��<�b�<(Ƌ<�(�<Z��<��<�z<�Zs<l<��d<u�]<UgV<.O<�G<��@<��9<�c2<:+<�$<��<�<!�<!�<t� <]K�;hT�;�l�;��;�λ;�;lx�;,�;zp�;p;�zU;�;;� ;׼;9��:�o�:�g:%!:Ɗ�8�4��JZ'�:U��0����4��	��!�'8���N��e��{������ᓻ����H���ɳ�[(��{eȻ<�һg{ܻ/T�/𻜣��Z��9���
�ta�����L������ �A%�rv)�o�-�?�1�H�5���9�h�=��A�M�E��YI�"M��P�)�T�t>X�`�[�:w_�fc�*�f��j���m��p�bZt���w��{��j~��܀�����"������^�����Ꮚ��%��+����J���ڐ��h��e���h����	��9���5������#������|*�������-�������.��,���N-������*��ɨ���&��ߤ���"��䠳���h������򚹼G�����`���  �  tN=E�M=�L=�0L=�nK=�J=��I=h%I=2aH=h�G=��F=�F=�IE=��D=X�C=��B=g%B=�YA=z�@=�?=5�>=V!>=-P==�}<=��;=��:=�9=�%9=L8=}p7=I�6=8�5=T�4=x�3=�3=�$2=�;1=(P0=sb/=er.=�-=��,=�+=j�*=#�)=�(=͗'=��&=,�%=�{$=�k#=rX"=�A!=r' =�	=��=��=��=�l=�;=�=��=��=�O=C
=��=s=/!=	�=�p==L�	=UH="�=�m=n�=��={=�<t	�<��<K��<��<���<$x�<�E�<��<Y��<���<�;�<���<z��<�5�<l��</l�<3 �<���<��<R��<6$�<a��<��<g��<��<,�<��<m\�<�ǝ<�0�<R��<*��<�b�< Ƌ<�(�<c��<��<
�z<�Zs<�l<��d<p�]<VgV<$.O<,�G<��@<��9<�c2<:+<{$<��<=�<�<'�<h� <mK�;JT�;�l�;:��;�λ;7�;cx�;h�;xp�;�p;{U;�;;� ;��;���:�o�:�g:(!:��8p3���Z'�hT��7���b4��	�,!�	'8���N��e�Y�{�\����ᓻ0����H���ɳ�Z(���eȻ׀һ0{ܻ3T�𻘣��I��9���
�wa����M������ �A%�bv)�e�-�5�1�G�5���9�2�=�!�A�R�E��YI�
"M��P�,�T�^>X�p�[�5w_�pc�&�f��j���m��p�mZt���w��{��j~��܀�����"�������]����������%��$����J���ڐ��h��f���b����	��2���-������#������x*�������-��~����.��)���W-������*��Ĩ���&��ᤰ��"��𠳼��s��� ��򚹼A��
���g���  �  tN=I�M=!�L=�0L=~nK= �J=��I=e%I=7aH=g�G=��F=�F=�IE=�D=X�C=��B=`%B=�YA=u�@=�?=7�>=U!>=3P==�}<=��;=��:=�9=�%9=L8=�p7=D�6=:�5=N�4=x�3=�3=�$2=�;1='P0=ub/=br.=�-=��,=�+=q�*="�)=�(='=��&=/�%=�{$=�k#=mX"=�A!=n' =�	=��=��=��=�l=�;=�=��=��=�O=E
=��=s=/!=�=�p==P�	=RH='�=�m=s�=��=|=�<k	�<��<C��<��<���<'x�<�E�<��<U��<���<�;�<���<z��<�5�<_��<0l�<% �<���<��<N��<3$�<]��<��<a��<��<$�<��<d\�<�ǝ<�0�<S��<5��<�b�<$Ƌ<�(�<]��<��<�z<�Zs<�l<��d<s�]<PgV<.O<"�G<��@<��9<�c2<:+<�$<��<,�<.�<�<{� <dK�;5T�;�l�;��;�λ;6�;bx�;0�;zp�;�p;{U;�;;�� ;�;���:Vo�:�g:�":���8@4���Y'�U������5��	��!�'8���N�%�e�2�{�t����ᓻ>����H��mɳ�_(���eȻ0�һ1{ܻT�;𻉣��`��9���
�ua����	M������ �A%�{v)�e�-�E�1�=�5���9�]�=��A�S�E�YI�"M� �P��T�l>X�`�[�=w_�\c�*�f��j���m�$�p�\Zt���w�{��j~��܀������"������^����������%��(����J���ڐ��h��e���d����	��5���1������#������*�������-�������.��)���K-������*��ƨ���&��ᤰ��"��ߠ��
��c����������C�����c���  �  tN=J�M=�L=�0L=�nK=��J=��I=`%I=9aH=d�G=��F=�F=�IE=��D=Q�C=��B=^%B=�YA=v�@=�?=8�>=O!>=2P==�}<=��;=��:=�9=�%9=�K8=�p7=B�6=<�5=O�4=z�3=�3=�$2=�;1=$P0=zb/=_r.=�-=��,=�+=m�*=�)=��(=��'=��&=,�%=�{$=�k#=iX"=�A!=i' =�	=��=��=��=�l=�;=�=��=��=�O=B
=��= s=*!=�=�p==T�	=OH=+�=�m=u�=��=}=!�<j	�<!��<=��<��<���<*x�<�E�<��<n��<���<�;�<���<~��<�5�<`��<3l�<  �<���<u�<Q��<3$�<S��<�<\��<��<�<��<^\�<�ǝ<�0�<E��<4��<�b�<+Ƌ<�(�<Z��<��<�z<�Zs<ml<��d<k�]<WgV<.O<$�G<��@<��9<�c2<�9+<�$<��<�<#�<�<�� <PK�;CT�;�l�;��;�λ;��;vx�;"�;yp�;�p;{U;�;;�� ;��;Y��:�p�:�g:� :{��86���X'�HU������5���	��!�Q'8�e�N�Z�e���{������ᓻ/����H���ɳ��(��GeȻ3�һG{ܻ4T�I�q���m���8�	�
�ia����M������ �A%��v)�Y�-�I�1�N�5���9�g�=��A�g�E��YI�"M��P��T�z>X�P�[�Kw_�Tc�1�f��j���m�'�p�OZt�»w�j{�k~��܀�
����"��}���^�����돊��%��#����J���ڐ��h��^���p����	��4���;������#�������*�������-�������.��6���M-������*��¨���&��ڤ���"��ݠ����`�����򚹼E�����Z���  �  tN=L�M=�L=�0L=�nK=�J=��I=d%I=5aH=d�G=��F=�F=�IE=��D=V�C=��B=b%B=�YA=x�@=�?=6�>=S!>=3P==�}<=��;=��:=�9=�%9= L8=�p7=E�6=9�5=T�4=y�3=�3=�$2=�;1=&P0=xb/=_r.=�-=��,=�+=q�*= �)=�(=ŗ'=��&=+�%=�{$=�k#=mX"=�A!=k' =�	=��=��=��=�l=�;=�=��=��=�O=F
=��=s=-!=�=�p==Q�	=PH=(�=�m=r�=��=}=�<t	�<��<D��<��<���<1x�<�E�<��<X��<���<�;�<���<y��<�5�<f��<*l�<' �<���<|�<P��<1$�<R��< �<^��<��<%�<��<o\�<�ǝ<�0�<M��<7��<�b�<'Ƌ<�(�<Y��<��<	�z<�Zs<�l<��d<q�]<bgV<.O<,�G<��@<��9<�c2<:+<}$<��<=�<"�<�<r� <MK�;ET�;zl�;��;�λ;&�;lx�;<�;Wp�;�p;�zU;�;;�� ;�;=��:~o�:g:T!:]��8�4���Y'��T��7���k4��	�!��&8���N�4�e��{������ᓻ<����H��oɳ�r(���eȻ�һ{ܻ=T�8𻚣��_��9��
�pa����M������ �A%�wv)�k�-�E�1�P�5���9�T�=��A�Z�E��YI��!M��P��T�t>X�]�[�;w_�bc�$�f��j���m��p�_Zt���w�w{��j~��܀�����"�������]�����䏊��%��+����J���ڐ��h��b���i����	��6���=������#������~*�������-�������.��.���J-������*�������&��ؤ���"��⠳���d��� ��욹�H��
���_���  �  tN=E�M="�L=�0L=~nK= �J=��I=d%I=2aH=h�G=��F=�F=�IE=�D=W�C=��B=a%B=�YA={�@=�?=5�>=S!>=-P==�}<=�;=��:=�9=�%9=L8=~p7=I�6=9�5=W�4=z�3=�3=�$2=�;1=.P0=xb/=fr.=�-=��,=�+=l�*=*�)=�(=ė'=��&=*�%=�{$=�k#=qX"=�A!=o' =�	=��=��=��=�l=�;=�=��=��=�O=@
=��=s=8!=�=�p==R�	=WH='�=�m=q�=��==�<{	�<��<O��<��<���<*x�<�E�<��<R��<���<�;�<���<|��<�5�<l��<'l�<( �<x��<~�<F��<1$�<[��<��<g��<��<'�<��<b\�<�ǝ<�0�<Z��<)��<�b�< Ƌ<�(�<a��<��<"�z<�Zs<�l<��d<��]<dgV<#.O<0�G<��@<��9<�c2<":+<�$<��<-�<�<�<i� <mK�;JT�;�l�;��;uλ;/�;-x�;5�;Qp�;�p;�zU;�;;�� ;��;5��:�n�:�g:A":���8�2���Z'��T��&���4��	��!��&8���N���e��{�W����ᓻ1����H���ɳ�"(���eȻ �һV{ܻFT�+𻻣��O��9���
�ya����M������ �(A%�hv)�z�-�:�1�P�5���9�V�=��A�0�E��YI�"M��P��T�X>X�_�[�"w_�gc��f��j���m��p�aZt���w��{��j~��܀�����"�������]�����䏊��%��0����J���ڐ��h��q���f���
��6���3������#������|*�������-�������.��!���X-��	����*�������&��٤���"��⠳���d������뚹�B��	���g���  �  tN=H�M=�L=�0L=�nK= �J=��I=a%I=5aH=b�G=��F=�F=�IE=�D=V�C=��B=b%B=�YA=v�@=�?=8�>=Q!>=1P==�}<=��;=��:=�9=�%9=L8=�p7=G�6=>�5=R�4=w�3=�3=�$2=�;1=&P0=xb/=dr.=�-=��,=�+=k�*=�)=�(=Ɨ'=��&=/�%=�{$=�k#=kX"=�A!=m' =�	=��=��=��=�l=�;=�=��=��=�O=D
=��=s=+!=	�=�p==O�	=SH=)�=�m=r�=��=�=�<r	�< ��<H��<��<���<,x�<�E�<��<c��<���<�;�<���<���<�5�<c��<.l�<) �<���<|�<N��<2$�<X��<��<Z��<��< �<��<b\�<�ǝ<�0�<A��<0��<�b�<%Ƌ<�(�<f��<��<�z<�Zs<|l<��d<n�]<_gV<0.O<&�G<��@<��9<�c2<�9+<�$<��<*�<)�<�<s� <>K�;4T�;�l�; ��;�λ;!�;Xx�;=�;bp�;�p;�zU;�;;�� ;�;���:p�:;g:�:��8�3��0Z'��T�������4�1�	��!�'8���N�=�e��{�k����ᓻ)����H���ɳ��(���eȻ�һ@{ܻT�/𻪣��h��9���
�|a����M������ �A%�v)�u�-�9�1�C�5���9�P�=��A�g�E��YI�"M��P�#�T�h>X�Y�[�@w_�`c��f��j���m��p�SZt���w��{��j~��܀�����"������ ^�����揊��%��0����J���ڐ��h��f���h����	��6���7������#�������*�������-�������.��;���Q-������*��Ũ���&��٤���"��ߠ����`������;�����b���  �  tN=R�M=�L=�0L=�nK=��J=��I=^%I=9aH=_�G=��F=�F=�IE=�D=P�C=��B=\%B=�YA=u�@=�?=8�>=P!>=5P==�}<=��;=��:=�9=�%9=�K8=�p7=C�6==�5=U�4=y�3=�3=�$2=�;1=&P0=}b/=`r.=�-=��,=�+=v�*=�)=�(=��'=��&=,�%=�{$=�k#=eX"=�A!=g' =�	=��=��=��=�l=�;=�=��=��=�O=D
=��=s=,!=�=�p==R�	=PH=-�=�m=t�=��=�=!�<v	�<$��<@��<��<���<7x�<�E�<��<c��<���<�;�<���<|��<�5�<^��<+l�< �<���<s�<N��<+$�<O��< �<R��<��<�<��<[\�<�ǝ<�0�<N��<D��<�b�<1Ƌ<�(�<]��<��<�z<�Zs<�l<�d<p�]<mgV<!.O<"�G<��@<��9<d2<:+<�$<��<�<+�< �<�� <(K�;>T�;ql�;���;�λ;��;[x�;
�;Sp�;�p;�zU;�;;�� ;�;���:�o�:�g:�":��8�5��Y'�9U������S4��	��!��&8�w�N�D�e���{������ᓻ����H��Bɳ�|(���eȻJ�һJ{ܻ/T�Q𻂣��}��9��
��a����M����� �A%��v)�d�-�L�1�M�5���9�u�=��A�a�E�jYI��!M��P��T�y>X�G�[�?w_�Yc��f��j���m��p�JZt���w�p{��j~��܀������"������^�����鏊��%��-����J���ڐ��h��f���r����	��<���@������#�������*�������-�������.��-���=-�����|*��Ǩ���&��Ѥ���"��٠����]�����皹�C�����V���  �  tN=C�M=�L=�0L=�nK=�J=��I=c%I=5aH=c�G=��F=�F=�IE=�D=V�C=��B=_%B=�YA=w�@=�?=5�>=S!>=4P==�}<=��;=��:=�9=�%9=L8=�p7=I�6=:�5=W�4=z�3=�3=�$2=�;1=,P0=wb/=fr.=�-=��,=�+=k�*=!�)=�(=Ǘ'=��&=/�%=�{$=�k#=jX"=�A!=k' =�	=��=��=��=�l=�;=�=��=��=�O=E
=��=s=/!=�=�p= =R�	=WH=(�=�m=p�=��== �<{	�<��<M��<��<���<"x�<�E�<��<`��<���<�;�<���<{��<�5�<e��<-l�<% �<}��<~�<J��<0$�<T��< �<]��<��<"�<��<h\�<�ǝ<�0�<P��<)��<�b�<*Ƌ<�(�<`��<��<�z<�Zs<�l<��d<��]<dgV< .O<8�G<��@<��9<�c2<:+<�$<��<0�<*�<�<q� <IK�;BT�;l�;
��;�λ;#�;Cx�;$�;ap�;�p;�zU;�;;�� ;�;���:�o�:�g:�!:^y�8y3��Z'�vT�����4���	�!��&8���N��e��{�\����ᓻ����H���ɳ�h(���eȻ�һ2{ܻT�7𻘣��l��	9��
�}a����
M������ �A%��v)�i�-�A�1�?�5���9�S�=��A�T�E��YI�"M��P��T�]>X�]�[�-w_�lc��f��j���m��p�ZZt���w�~{��j~��܀�����"������^�����⏊��%��-����J���ڐ��h��l���f��� 
��7���;������#�������*�������-�������.��,���X-������*�������&��٤���"��砳���j������뚹�C�����_���  �  �vN=��M=��L=�4L=GsK=E�J=��I=�+I=hH=ţG=��F=,F=�RE=��D=��C=��B=�0B=�eA=.�@=L�?=J�>=0>=�_==�<=ߺ;=v�:=�:=99=`8=R�7=��6=��5=��4=�4=�$3=�>2=mV1=l0=7/=�.=k�-=>�,=s�+=ֹ*=��)=1�(=�'=��&=#�%=q�$=f�#=��"=�j!=�Q =f4=�=��=j�=
�=�i=35=��=�=/=:=��=E�={Q=P�=�=,B="�	=�w=^=��=�(=Ű=�4=)i�<a�<-Q�<�9�<��<|��<
��<���<�W�<��<���<��<�+�<���<Ur�<��<��<l5�<��<�J�<�ν<O�<�˶<�D�<V��<-�<ܜ�<�	�<�t�<]ݝ<D�<䨖<�<n�<�΋<�.�<䍄<p�<��z<�Qs<�l<��d<J�]<�IV<�O<��G<ؕ@<�_9<�,2<��*<�#<�<I�<q<\<<M <���;7��;���;/��;z�;g'�;k{�;��;7`�;��m;q5S;L�8;�b;B;ĩ�:t7�:Rf\:�p�9�b�8�堹��2�84���y���@�����&$�MG;�)&R���h���ϕ���}��C���媻�f��IĿ�� ʻRԻL޻^�����0���Q���������=����Aa�"�!�.�%�� *�eE.��\2��f6��d:�yV>�f<B��F��I���M��dQ�U�F�X��X\�~�_�xc��f�vj�=�m��Tq���t�|x�o{���~����O���IH���兼����Q�������C��֍�yf�����ˁ��*��і��C��C���,��ఛ�u4��'����8�����J:��빤��8��w����5��_���1��C���X+�����%���������W���������\��:�������  �  �vN=��M=��L=�4L=OsK=L�J=��I=�+I=
hH=ţG=��F=+F=�RE=��D=��C=��B=�0B=fA=6�@=L�?=F�>=0>=�_==��<=�;=n�:=�:=99=`8=\�7=��6=��5=��4=�4=�$3=�>2=sV1=l0=8/=�.=o�-==�,=e�+=Թ*=w�)=3�(=��'=��&=)�%=n�$=e�#=��"=k!=�Q =h4=�=��=n�=�=�i=65=��=�=2=(:=��=J�=pQ=L�=ݠ=(B=(�	=�w=_=��=�(=̰=�4=,i�<a�<*Q�<�9�<��<j��<���<���<�W�<��<���<��<�+�<���<Vr�<��<��<b5�<'��<�J�<�ν<O�<�˶<�D�<U��<�,�<Ӝ�<
�<�t�<kݝ<�C�<Ѩ�<�<n�<�΋<�.�<ԍ�<s�<��z< Rs<�l<��d<?�]<�IV<�O<v�G<��@<�_9<�,2<��*<��#</�<e�<7q<�[<3M <���;���;���;��;��;"'�;�{�;��;_`�;4�m;|5S;�8;�b;�B;d��:�8�:Zd\:�l�9�T�8S령N�2�)5��Tz���@����P&$��F;��%R���h���*����}��C��
檻�f���Ŀ�u ʻԻ�޻4��$���0���Q�f������Y����2a�4�!�
�%�� *�gE.��\2��f6��d:�fV>�R<B��F�&�I���M��dQ��U�q�X��X\���_��wc���f��uj�6�m�Uq�ǹt��x��n{��~����^���\H���兼����=�������C��֍�jf�����ԁ����㖕�E��F���,��̰��w4��,����8��󹡼=:��ݹ���8�������5��{����0��C���h+��|����%���������M����������h��?�������  �  �vN=��M=��L=�4L=MsK=A�J=��I=�+I=hH=��G=��F=)F=�RE=��D=��C=��B=�0B=fA=3�@=J�?=J�>=0>=�_==�<=�;=m�:=�:=99=`8=e�7=�6=��5=��4=�4=�$3=�>2=wV1=�k0=A/=�.=u�-=@�,=f�+=�*=v�)=7�(=�'=��&=!�%=k�$=g�#=��"=k!=�Q =m4=�=��=u�= �=�i=/5=��=�=+= :=��=O�=oQ=[�=�=)B=0�	=�w=i=��=�(=°=�4=-i�<a�<6Q�<�9�<��<e��<
��<���<�W�<��<���<��<�+�<���<Sr�<��<���<S5�<8��<�J�<�ν<O�<�˶<�D�<J��<-�<͜�<
�<�t�<fݝ<�C�<Ө�<-�<�m�<�΋<�.�<э�<~�<��z<Rs<�l<��d<;�]<JV<�O<q�G<�@<}_9<�,2<��*<�#<(�<8�<.q<�[<MM <���;���;���;��;��;%'�;�{�;��;p`�; �m;[5S;O�8;Hb;eB;���:�8�:d\:q�9�k�8>�7�2��5���y���@�����&$��G;��%R�(�h�V�F����}���B�� 檻f���Ŀ�Z ʻ]ԻF޻p��7���0��R�X������A����a�N�!� �%�!*�dE.��\2�g6��d:��V>�?<B��F���I���M��dQ��U���X�mX\���_��wc��f�vj�5�m�Uq���t��x��n{�'�~����H���^H���兼����F�������C��!֍�uf������䁒���▕�3��E���&,��Ȱ���4�� ����8������S:��㹤��8�������5�������0��@���k+��q����%���������L��� ������f��B�������  �  �vN=��M=��L=�4L=KsK=J�J=��I=�+I=hH=ģG=��F=.F=�RE=��D=��C=��B=�0B=	fA=0�@=M�?=J�>=0>=�_==�<=�;=p�:=�:=99=`8=\�7=�6=��5=��4=�4=�$3=�>2=zV1=�k0=</=�.=o�-=<�,=h�+=׹*=v�)=6�(=�'=��&=(�%=m�$=i�#=�"=
k!=�Q =e4=�=��=m�=�=�i=35=��=�=1=(:=��=L�=pQ=O�=�=(B=)�	=�w=d=��=�(=Ű=�4=3i�<a�<3Q�<�9�<��<j��<��<���<�W�<��<���<��<�+�<���<Yr�<��<���<\5�<'��<�J�<�ν<O�<�˶<�D�<S��<-�<Ҝ�<
�<�t�<gݝ<�C�<Ϩ�<�<n�<�΋<�.�<؍�<p�<��z<Rs<�l<�d<<�]<�IV<�O<p�G<��@<�_9<�,2<��*<
�#< �<\�<Gq<�[<NM <���;u��;���;��;��;5'�;�{�;��;�`�;��m;�5S;W�8;�b;�B;$��:�8�:�d\:Wm�9M`�8�꠹.�2�h5���y��TA����J&$�zG;�P%R�H�h���.����}��C���媻uf���Ŀ�c ʻ8Ի�޻5��%���0���Q�\������K����6a�4�!���%�� *�\E.��\2��f6��d:�qV>�I<B��F��I���M��dQ��U�t�X�X\���_��wc� �f��uj�(�m�Uq���t��x��n{��~����[���\H���兼����9�������C��֍�wf������ځ��������=��M���,��Ͱ��y4������8��칡�=:��⹤��8�������5��x����0��C���e+��~����%���������E��� �����`��C�������  �  �vN=��M=��L=�4L=HsK=J�J=��I=�+I=
hH=ɣG=��F=,F=�RE=��D=��C=��B=�0B=fA=2�@=P�?=F�>=0>=�_==�<=�;=t�:=�:=99=`8=Y�7=��6=��5=��4=�4=�$3=�>2=rV1=�k0=:/=�.=n�-=>�,=m�+=Թ*=�)=/�(=�'=��&=%�%=m�$=c�#=��"=k!=�Q =f4=�=��=m�=�=�i=55=��=�=/=!:=��=E�=xQ=M�=�=*B=&�	=�w=a=��=�(=ð=�4=)i�<a�<+Q�<�9�<��<s��<��<���<�W�<��<���<��<�+�<���<[r�<��<��<e5�<*��<�J�<�ν<	O�<�˶<�D�<^��<�,�<Ҝ�<
�<�t�<^ݝ<�C�<ᨖ<�<n�<�΋<�.�<ҍ�<q�<��z<�Qs<�l<��d<@�]<�IV<�O<o�G<�@<�_9<�,2<��*<�#<�<^�<!q<�[<3M <͊�;`��;���;��;��;i'�;�{�;��;_`�;��m;�5S;�8;�b;3B;)��:�7�:�e\:�n�9b]�8*蠹��2�.5��1z���@�����&$��G;��%R��h���*����}��C���媻�f��_Ŀ�� ʻBԻ"޻N��$���0���Q�x������8����5a�*�!��%�� *�gE.��\2��f6��d:�rV>�e<B��F� �I���M��dQ�U�r�X��X\���_�xc��f��uj�:�m�Uq�ùt��x�o{�
�~����Y���MH���兼����L�������C��֍�rf�����ҁ����Җ��8��I���,��ְ��n4��-����8������@:��깤��8��z����5��j����0��F���j+��}����%���������S���������i��C�������  �  �vN=��M=��L=�4L=OsK=I�J=��I=�+I=hH=ãG=��F=/F=�RE=��D=��C=��B=�0B=fA=3�@=K�?=J�>=0>=�_==�<=�;=k�:=�:=99=`8=[�7=��6=��5=��4=�4=�$3=�>2=rV1=�k0=:/=�.=r�-=<�,=h�+=׹*=v�)=0�(=��'=��&='�%=v�$=d�#=�"=
k!=�Q =i4=�=��=o�=�=�i=25=��=�=3= :=��=F�=oQ=N�=�=%B=*�	=�w=`=��=�(=ǰ=�4=%i�<a�<)Q�<�9�<��<b��<��<���<�W�<��<���<��<�+�<���<Sr�<��<���<a5�<.��<�J�<�ν<O�<�˶<�D�<Q��<�,�<木<
�<�t�<mݝ<�C�<Ѩ�<�<n�<�΋<�.�<̍�<w�<��z<�Qs<�l<��d<0�]<JV<�O<z�G<��@<�_9<�,2<��*<��#<0�<W�<!q<$\<?M <���;|��;���;,��;��;"'�;�{�;��;�`�;�m;v5S;\�8;c;5B;1��:�8�:�c\:�m�9@e�8�젹a�2�)5��<z���@�,��o&$�DG;��%R�;�h���G����}��C���媻tf���Ŀ�� ʻԻ1޻=������0���Q�[������D����,a�1�!���%� !*�hE.��\2��f6��d:�`V>�_<B��F��I���M��dQ��U���X��X\���_��wc���f��uj�A�m�Uq�ƹt��x��n{�*�~����[���`H���兼����K�������C�� ֍�rf������Ձ����▕�6��B���,��Ͱ��{4��*����8������E:��۹��9�������5��|����0��@���p+��x����%���������P���������m��>�������  �  �vN=��M=��L=�4L=OsK=H�J=��I=�+I=hH=ţG=��F=1F=�RE=��D=��C=��B=�0B=fA=5�@=N�?=I�>=0>=�_==�<=�;=s�:=�:=99=	`8=Z�7=�6=��5=��4=�4=�$3=�>2=tV1=�k0=@/=�.=n�-=;�,=h�+=ٹ*=x�)=7�(=�'=��&=(�%=o�$=h�#=�"=k!=�Q =j4=�=��=r�=�=�i=25=��=�=2=$:=��=M�=qQ=P�=�=&B=(�	=�w=f=��=�(=ð=�4=%i�<a�<5Q�<�9�<��<e��<��<���<�W�<��<���<��<�+�<���<Yr�<��<��<Y5�<4��<�J�<�ν<O�<�˶<�D�<U��<-�<Ӝ�<
�<�t�<jݝ<D�<Ψ�<�<n�<�΋<�.�<ԍ�<z�<q�z<Rs<�l<��d<"�]<JV<�O<g�G<�@<�_9<�,2<��*<�#<-�<V�<6q<�[<AM <���;���;ȗ�;��;��;>'�;�{�;��;�`�;+�m;�5S;F�8;�b;�B;���:�8�:�e\:�m�9�g�8�령��2��5��xy��A�"��i&$��G;��%R�t�h�n�B����}��C���媻df���Ŀ�Q ʻ5Ի޻4�����0���Q�F������8����a�=�!���%�� *�WE.��\2��f6��d:�tV>�D<B��F��I���M��dQ��U��X�uX\���_��wc��f��uj�@�m�Uq���t��x��n{�%�~����Z���VH���兼����B�������C��֍�rf������݁����ܖ��/��I���,��°��w4��&����8��򹡼B:��߹���8�������5��|����0��H���h+��t����%���������L���������b��G�������  �  �vN=��M=��L=�4L=EsK=K�J=��I=�+I=hH=ʣG=��F=0F=�RE=��D=��C=��B=�0B=
fA=2�@=R�?=J�>=0>=�_==�<=�;=u�:=�:=99=`8=X�7=�6=��5=��4=�4=�$3=�>2=pV1=�k0=;/=�.=k�-=?�,=m�+=չ*={�)=1�(=�'=��&='�%=m�$=i�#=��"=k!=�Q =j4=�=��=q�=�=�i=25=��=�=0=":=��=F�=vQ=L�=�=+B=$�	=�w=`=��=�(=��=�4=&i�<	a�<*Q�<�9�<��<t��<���<���<�W�<��<���<��<�+�<���<ar�<��<���<a5�<1��<�J�<�ν<	O�<�˶<�D�<^��<-�<М�<
�<�t�<Yݝ<D�<Ө�<�<n�<�΋<�.�<ύ�<q�<��z<�Qs<�l<��d<9�]<�IV<�O<\�G<�@<�_9<�,2<��*<�#<�<_�<4q<�[<EM <Պ�;u��;Ɨ�;��;��;g'�;�{�;��;�`�;��m;�5S;Y�8;�b;|B;��:�7�:7f\:�l�9i^�8`砹<�2��5��(z��A�����&$��G;��%R�7�h���?����}���B���媻�f��|Ŀ�� ʻUԻ޻@��'��0���Q�`��ݔ���-����"a�,�!��%�� *�RE.��\2��f6��d:��V>�^<B��F�!�I���M��dQ�U���X��X\���_�	xc��f�vj�>�m�Uq�ùt��x�o{��~����_���OH���兼����F�������C��֍�tf������Ձ����Ӗ��2��H���,��ΰ��o4��#����8��󹡼@:��﹤��8�������5��k����0��M���m+��~����%���������R��� �����k��L�������  �  �vN=��M=��L=�4L=KsK=O�J=��I=�+I=hH=ȣG=��F=/F=�RE=��D=��C=��B=�0B=fA=5�@=N�?=I�>=0>=�_==��<=�;=m�:=�:=99=`8=V�7=��6=��5=��4=�4=�$3=�>2=nV1=�k0=4/=�.=n�-=9�,=f�+=Թ*=x�)=/�(=��'=��&='�%=t�$=d�#=��"=	k!=�Q =j4=�=��=q�=
�=�i=55=��=�=2=!:=��=D�=rQ=K�=ߠ=$B=%�	=�w=Y=��=�(=Ű=�4=i�<
a�<Q�<�9�<��<b��<���<���<�W�<��<���<��<�+�<���<Xr�<��<���<f5�<0��<�J�<�ν<O�<�˶<�D�<\��<-�<䜨<
�<�t�<iݝ<�C�<Ө�<�<n�<�΋<�.�<̍�<i�<��z<�Qs<�l<��d<3�]<�IV<�O<t�G<�@<�_9<�,2<��*<��#<�<o�<$q<!\<?M <Ŋ�;���;���;8��;��;V'�;�{�;��;�`�;4�m;�5S;L�8;.c;EB;%��:
8�:wd\:�m�9�]�85젹��2�5���z��A�3���&$�8G;�&R��h��9����}��)C���媻�f���Ŀ�� ʻԻ޻;�����0���Q�\��ؔ���7����%a� �!���%�� *�eE.��\2��f6��d:�XV>�e<B��F�#�I���M��dQ�	U�w�X��X\���_�xc���f��uj�M�m�Uq�ܹt��x�o{�(�~����[���[H���兼����L�������C��֍�lf������Ё����ږ��5��@���,��̰��p4��'����8������<:��߹���8�������5��z���1��C���p+�������%���������W�����
���p��@�������  �  �vN=��M=��L=�4L=KsK=I�J=��I=�+I=hH=ǣG=��F=,F=�RE=��D=��C=��B=�0B=fA=7�@=P�?=J�>=0>=�_==�<=�;=q�:=�:=99=`8=]�7=�6=��5=��4=�4=�$3=�>2=mV1=�k0=;/=�.=n�-=<�,=f�+=ݹ*=x�)=6�(=�'=��&='�%=p�$=i�#=��"=k!=�Q =o4=�=��=x�=�=�i=55=��=�=1=":=��=K�=qQ=S�=�=%B=&�	=�w=`=��=�(=��=�4=i�<a�<(Q�<�9�<��<a��<��<���<�W�<��<���<��<�+�<���<[r�<��<���<`5�<A��<�J�<�ν<O�<�˶<�D�<Y��<-�<؜�<
�<�t�<cݝ<�C�<Ө�<%�<n�<�΋<�.�<ʍ�<t�<x�z<�Qs<�l<��d<'�]<�IV<�O<_�G<��@<�_9<�,2<��*<
�#<�<W�<)q<\<IM <Ê�;���;���;9��;��;V'�;|�;��;�`�;[�m;�5S;a�8;�b;tB;��:�8�:e\:�o�9m�8>젹��2��5��(z��A�O���&$��G;�&R�X�h���M����}��C���媻@f���Ŀ�[ ʻJԻ޻<����0���Q�M������0����	a�5�!���%�� *�WE.��\2��f6��d:�{V>�H<B��F��I���M��dQ�U��X��X\���_�xc��f�vj�Q�m�Uq�Ĺt��x��n{�*�~����R���WH���兼����F�������C��֍�lf������ց����ٖ��*��<���,��ð��s4��!����8������C:��湤��8�������5��|����0��L���r+��z����%���������[���
�����m��K�������  �  �vN=��M=��L=�4L=IsK=N�J=��I=�+I=hH=ƣG=��F=3F=�RE=��D=��C=��B=�0B=fA=4�@=R�?=P�>=0>=�_==�<=�;=p�:=|:=99=`8=\�7=�6=��5=��4=�4=�$3=�>2=uV1=�k0=8/=�.=k�-=;�,=b�+=׹*=p�)=9�(=�'=��&=)�%=n�$=q�#=�"=k!=�Q =l4=�=��=u�=�=�i=25=��=�=1=-:=��=N�=iQ=L�=۠=#B=$�	=�w=_=��=�(=��=�4=*i�<�`�<+Q�<�9�<��<\��<���<���<�W�<��<���<��<�+�<���<er�<��<��<d5�<:��<�J�<�ν<O�<�˶<�D�<T��<-�<Μ�<
�<�t�<_ݝ<D�<���<�<�m�<�΋<�.�<ύ�<l�<q�z<Rs<�l<��d<)�]<�IV<�O<U�G<��@<z_9<�,2<��*<�#<�<k�<Nq<�[<gM <���;���;ޗ�;/��;��;;'�;�{�;��;�`�;#�m;�5S;��8;�b;1C;2��:�8�:e\:j�9�_�8���2�06���y���A�����&$��G;��%R���h���O����}��C��檻qf���Ŀ�? ʻOԻ�޻)����~0���Q�C��ݔ���A����a�*�!���%�� *�;E.��\2��f6��d:�}V>�<<B��F��I���M��dQ�U���X��X\���_��wc��f� vj�4�m�-Uq���t��x��n{�3�~����g���^H���兼����.�������C��֍�rf������ҁ����ߖ��3��B���,��Ű��x4������8��빡�5:��깤��8�������5�������0��P���m+�������%���������M��������i��P�������  �  �vN=��M=��L=�4L=IsK=I�J=��I=�+I=hH=ɣG=��F=0F=�RE=��D=��C=��B=�0B=fA=6�@=P�?=J�>=0>=�_==�<=�;=t�:=�:=99=`8=W�7=�6=��5=��4=�4=�$3=�>2=mV1=�k0=6/=�.=l�-=:�,=g�+=ܹ*={�)=4�(=�'=��&=!�%=o�$=h�#=��"=k!=�Q =k4=�=��=r�=�=�i=55=��=�=+=:=��=I�=tQ=R�=�=$B=$�	=�w=\=��=�(=��=�4=!i�<a�<%Q�<�9�<��<b��<��<���<�W�<��<���<��<�+�<���<Zr�<��<���<i5�<1��<�J�<�ν<O�<�˶<�D�<]��<-�<ל�<�	�<�t�<`ݝ<D�<ר�<�<n�<�΋<�.�<ԍ�<i�<��z<�Qs<�l<��d<3�]<�IV<�O<f�G<�@<�_9<�,2<��*<�#<�<Y�<q<\<HM <ӊ�;���;ȗ�;5��;��;�'�;�{�;��;�`�;I�m;�5S;e�8;�b;6B;,��:e8�:f\:wo�9Nh�8�령)�2��5��#z��MA���'$��G;�&R�)�h��� ����}��"C���媻Lf��xĿ�k ʻGԻ,޻m�����0���Q�`��Ք�����z�a��!��%�� *�ZE.��\2� g6��d:�{V>�P<B��F��I���M��dQ�U�r�X��X\���_�xc��f�vj�E�m�Uq�ɹt��x�o{�(�~����S���QH���兼����N�������C��֍�kf������́����ǖ��-��A���,��Ͱ��o4��!����8�����D:��鹤��8�������5��|���1��K���h+�������%���������_�����
���g��G�������  �  �vN=��M=��L=�4L=NsK=Q�J=��I=�+I=hH=ΣG=��F=0F=�RE=��D=��C=��B=�0B=fA=?�@=N�?=F�>=$0>=�_==��<=�;=m�:=�:=99=`8=Z�7=�6=��5=��4=�4=�$3=�>2=gV1=l0=./=�.=k�-=>�,=g�+=ѹ*=x�)=,�(=��'=��&=,�%=w�$=`�#=�"=	k!=�Q =i4=�=��=n�=�=�i=?5=��=�=8=$:=��=C�=pQ=H�=ߠ='B=#�	=�w=T=��=�(=Ű=�4=i�<
a�<Q�<�9�<��<h��<���<���<�W�<��<���<��<�+�<���<Sr�<��<��<r5�<%��<�J�<�ν<O�<�˶<�D�<k��<�,�<휨<
�<�t�<nݝ<�C�<̨�<�<n�<�΋<�.�<�<c�<��z<�Qs<�l<��d<?�]<�IV<mO<a�G<�@<�_9<�,2<��*<��#<(�<y�<&q<6\<$M <���;���;�;E��;��;�'�;�{�;�;�`�;��m;�5S;#�8;�c;CB;w��:�8�:|d\:#l�9�[�8�頹��2�]5��c{���@�	���&$�'G;�m&R���h�z�Q����}��C���媻�f���Ŀ�� ʻ�Ի�޻��М�1���Q�_��Ŕ���=����.a��!�	�%�� *�tE.��\2��f6��d:�QV>�i<B��F�/�I���M��dQ�U���X��X\���_�"xc���f�vj�I�m�Uq��t��x�o{��~����e���^H���兼����K�������C��֍�Uf������ā����Ж��9��?���,��İ��a4��5����8������3:��۹��9�������5��s����0��L���z+�������%���������d���������z��I�������  �  �vN=��M=��L=�4L=IsK=I�J=��I=�+I=hH=ɣG=��F=0F=�RE=��D=��C=��B=�0B=fA=6�@=P�?=J�>=0>=�_==�<=�;=t�:=�:=99=`8=W�7=�6=��5=��4=�4=�$3=�>2=mV1=�k0=6/=�.=l�-=:�,=g�+=ܹ*={�)=4�(=�'=��&=!�%=o�$=h�#=��"=k!=�Q =k4=�=��=r�=�=�i=55=��=�=+=:=��=I�=tQ=R�=�=$B=$�	=�w=\=��=�(=��=�4=!i�<a�<%Q�<�9�<��<b��<��<���<�W�<��<���<��<�+�<���<Zr�<��<���<i5�<1��<�J�<�ν<O�<�˶<�D�<]��<-�<ל�<�	�<�t�<`ݝ<D�<ר�<�<n�<�΋<�.�<ԍ�<i�<��z<�Qs<�l<��d<3�]<�IV<�O<f�G<�@<�_9<�,2<��*<�#<�<Y�<q<\<HM <ӊ�;���;ȗ�;5��;��;�'�;�{�;��;�`�;I�m;�5S;d�8;�b;6B;+��:d8�:f\:so�9>h�8�령+�2��5��$z��NA���'$��G;�&R�*�h��� ����}��"C���媻Mf��xĿ�k ʻGԻ-޻m�����0���Q�`��Ք�����z�a��!��%�� *�ZE.��\2� g6��d:�{V>�P<B��F��I���M��dQ�U�r�X��X\���_�xc��f�vj�E�m�Uq�ɹt��x�o{�(�~����S���QH���兼����N�������C��֍�kf������́����ǖ��-��A���,��Ͱ��o4��!����8�����D:��鹤��8�������5��|���1��K���h+�������%���������_�����
���g��G�������  �  �vN=��M=��L=�4L=IsK=N�J=��I=�+I=hH=ƣG=��F=3F=�RE=��D=��C=��B=�0B=fA=4�@=R�?=P�>=0>=�_==�<=�;=p�:=|:=99=`8=\�7=�6=��5=��4=�4=�$3=�>2=uV1=�k0=8/=�.=k�-=;�,=b�+=׹*=p�)=9�(=�'=��&=)�%=n�$=q�#=�"=k!=�Q =l4=�=��=u�=�=�i=25=��=�=1=-:=��=N�=iQ=L�=۠=#B=$�	=�w=_=��=�(=��=�4=*i�<�`�<+Q�<�9�<��<\��<���<���<�W�<��<���<��<�+�<���<er�<��<��<d5�<:��<�J�<�ν<O�<�˶<�D�<T��<-�<Μ�<
�<�t�<_ݝ<D�<���<�<�m�<�΋<�.�<ύ�<l�<q�z<Rs<�l<��d<)�]<�IV<�O<U�G<��@<z_9<�,2<��*<�#<�<k�<Nq<�[<gM <���;���;ޗ�;/��;��;;'�;�{�;��;�`�;#�m;�5S;��8;b;0C;1��:�8�:e\:j�9�_�8���2�26���y���A�����&$��G;��%R���h���O����}��C��檻qf���Ŀ�? ʻOԻ�޻)����~0���Q�C��ݔ���A����a�*�!���%�� *�;E.��\2��f6��d:�}V>�<<B��F��I���M��dQ�U���X��X\���_��wc��f� vj�4�m�-Uq���t��x��n{�3�~����g���^H���兼����.�������C��֍�rf������ҁ����ߖ��3��B���,��Ű��x4������8��빡�5:��깤��8�������5�������0��P���m+�������%���������M��������i��P�������  �  �vN=��M=��L=�4L=KsK=I�J=��I=�+I=hH=ǣG=��F=,F=�RE=��D=��C=��B=�0B=fA=7�@=P�?=J�>=0>=�_==�<=�;=q�:=�:=99=`8=]�7=�6=��5=��4=�4=�$3=�>2=mV1=�k0=;/=�.=n�-=<�,=f�+=ݹ*=x�)=6�(=�'=��&='�%=p�$=i�#=��"=k!=�Q =o4=�=��=x�=�=�i=55=��=�=1=":=��=K�=qQ=S�=�=%B=&�	=�w=`=��=�(=��=�4=i�<a�<(Q�<�9�<��<a��<��<���<�W�<��<���<��<�+�<���<[r�<��<���<`5�<A��<�J�<�ν<O�<�˶<�D�<Y��<-�<؜�<
�<�t�<cݝ<�C�<Ө�<%�<n�<�΋<�.�<ʍ�<t�<x�z<�Qs<�l<��d<'�]<�IV<�O<_�G<��@<�_9<�,2<��*<
�#<�<W�<)q<\<IM <Ê�;���;���;9��;��;V'�;|�;��;�`�;Z�m;�5S;`�8;�b;sB;��:�8�:ze\:�o�9�l�8H젹��2��5��+z��A�P���&$��G;�&R�Y�h���M����}��C���媻@f���Ŀ�\ ʻKԻ޻<����0���Q�M������1����	a�5�!���%�� *�WE.��\2��f6��d:�{V>�H<B��F��I���M��dQ�U��X��X\���_�xc��f�vj�Q�m�Uq�Ĺt��x��n{�*�~����R���WH���兼����F�������C��֍�lf������ց����ٖ��*��<���,��ð��s4��!����8������C:��湤��8�������5��|����0��L���r+��z����%���������[���
�����m��K�������  �  �vN=��M=��L=�4L=KsK=O�J=��I=�+I=hH=ȣG=��F=/F=�RE=��D=��C=��B=�0B=fA=5�@=N�?=I�>=0>=�_==��<=�;=m�:=�:=99=`8=V�7=��6=��5=��4=�4=�$3=�>2=nV1=�k0=4/=�.=n�-=9�,=f�+=Թ*=x�)=/�(=��'=��&='�%=t�$=d�#=��"=	k!=�Q =j4=�=��=q�=
�=�i=55=��=	�=2=!:=��=D�=rQ=K�=ߠ=$B=%�	=�w=Y=��=�(=Ű=�4=i�<
a�<Q�<�9�<��<b��<���<���<�W�<��<���<��<�+�<���<Xr�<��<���<f5�<0��<�J�<�ν<O�<�˶<�D�<\��<-�<䜨<
�<�t�<iݝ<�C�<Ө�<�<n�<�΋<�.�<̍�<i�<��z<�Qs<�l<��d<3�]<�IV<�O<t�G<�@<�_9<�,2<��*<��#< �<p�<$q<!\<?M <Ŋ�;���;���;8��;��;V'�;�{�;��;�`�;3�m;�5S;K�8;,c;CB;"��:8�:qd\:�m�9�]�8B젹��2�5���z��A�4���&$�9G;�	&R��h��9����}��*C���媻�f���Ŀ�� ʻ	Ի޻;�����0���Q�\��ؔ���7����%a� �!���%�� *�eE.��\2��f6��d:�XV>�e<B��F�#�I���M��dQ�	U�w�X��X\���_�xc���f��uj�M�m�Uq�ܹt��x�o{�(�~����[���[H���兼����L�������C��֍�lf������Ё����ږ��5��@���,��̰��p4��'����8������<:��߹���8�������5��z���1��C���p+�������%���������W�����
���p��@�������  �  �vN=��M=��L=�4L=EsK=K�J=��I=�+I=hH=ʣG=��F=0F=�RE=��D=��C=��B=�0B=
fA=2�@=R�?=J�>=0>=�_==�<=�;=u�:=�:=99=`8=X�7=�6=��5=��4=�4=�$3=�>2=pV1=�k0=;/=�.=k�-=?�,=m�+=չ*={�)=1�(=�'=��&='�%=m�$=i�#=��"=k!=�Q =j4=�=��=q�=�=�i=25=��=�=0=":=��=F�=vQ=L�=�=+B=$�	=�w=a=��=�(=��=�4=&i�<	a�<*Q�<�9�<��<t��<���<���<�W�<��<���<��<�+�<���<ar�<��<���<a5�<1��<�J�<�ν<	O�<�˶<�D�<^��<-�<М�<
�<�t�<Yݝ<D�<Ҩ�<�<n�<�΋<�.�<ύ�<p�<��z<�Qs<�l<��d<9�]<�IV<�O<\�G<�@<�_9<�,2<��*<�#<�<_�<4q<�[<EM <Պ�;u��;Ɨ�;��;��;g'�;�{�;��;�`�;��m;�5S;X�8;�b;zB;��:�7�:0f\:�l�90^�8n砹C�2��5��+z��A�����&$��G;��%R�9�h���@����}���B���媻�f��}Ŀ�� ʻVԻ޻@��(��0���Q�`��ݔ���-����"a�,�!��%�� *�RE.��\2��f6��d:��V>�^<B��F�!�I���M��dQ�U���X��X\���_�	xc��f�vj�>�m�Uq�ùt��x�o{��~����_���OH���兼����F�������C��֍�tf������Ձ����Ӗ��2��H���,��ΰ��o4��#����8��󹡼@:��﹤��8�������5��k����0��M���m+��~����%���������R��� �����k��L�������  �  �vN=��M=��L=�4L=OsK=H�J=��I=�+I=hH=ţG=��F=1F=�RE=��D=��C=��B=�0B=fA=5�@=N�?=I�>=0>=�_==�<=�;=s�:=�:=99=	`8=Z�7=�6=��5=��4=�4=�$3=�>2=tV1=�k0=@/=�.=n�-=;�,=h�+=ٹ*=x�)=7�(=�'=��&=(�%=o�$=h�#=�"=k!=�Q =j4=�=��=r�=�=�i=25=��=�=2=$:=��=M�=qQ=P�=�=&B=(�	=�w=f=��=�(=ð=�4=%i�<a�<5Q�<�9�<��<e��<��<���<�W�<��<���<��<�+�<���<Yr�<��<��<Y5�<4��<�J�<�ν<O�<�˶<�D�<U��<-�<Ӝ�<
�<�t�<jݝ<D�<Ψ�<�<n�<�΋<�.�<ԍ�<z�<q�z<Rs<�l<��d<"�]<JV<�O<g�G<�@<�_9<�,2<��*<�#<-�<V�<7q<�[<AM <���;���;ȗ�;��;��;>'�;�{�;��;�`�;*�m;�5S;E�8;�b;�B;��:�8�:�e\:�m�9�g�8�령��2��5��|y�� A�$��k&$��G;��%R�u�h�o�C����}��C���媻ef���Ŀ�R ʻ6Ի޻4�����0���Q�F������8����a�=�!���%�� *�WE.��\2��f6��d:�tV>�D<B��F��I���M��dQ��U��X�uX\���_��wc��f��uj�@�m�Uq���t��x��n{�%�~����Z���VH���兼����B�������C��֍�rf������݁����ܖ��/��I���,��°��w4��&����8��򹡼B:��߹���8�������5��|����0��H���h+��t����%���������L���������b��G�������  �  �vN=��M=��L=�4L=OsK=I�J=��I=�+I=hH=ãG=��F=/F=�RE=��D=��C=��B=�0B=fA=3�@=K�?=J�>=0>=�_==�<=�;=k�:=�:=99=`8=[�7=��6=��5=��4=�4=�$3=�>2=rV1=�k0=:/=�.=r�-=<�,=h�+=׹*=v�)=0�(=��'=��&='�%=v�$=d�#=�"=
k!=�Q =i4=�=��=o�=�=�i=25=��=�=3= :=��=F�=oQ=N�=�=&B=*�	=�w=`=��=�(=ǰ=�4=&i�<a�<)Q�<�9�<��<c��<��<���<�W�<��<���<��<�+�<���<Sr�<��<���<b5�<.��<�J�<�ν<O�<�˶<�D�<Q��<�,�<在<
�<�t�<mݝ<�C�<Ѩ�<�<n�<�΋<�.�<̍�<w�<��z<�Qs<�l<��d<0�]<JV<�O<z�G<��@<�_9<�,2<��*<��#<0�<W�<!q<$\<?M <���;|��;���;,��;��;"'�;�{�;��;�`�;�m;u5S;[�8;c;4B;-��:�8�:�c\:�m�9e�8�젹h�2�-5��?z���@�-��p&$�FG;��%R�<�h���H����}��C���媻uf���Ŀ�� ʻԻ1޻=�����0���Q�[������D����,a�1�!���%� !*�hE.��\2��f6��d:�`V>�_<B��F��I���M��dQ��U���X��X\���_��wc���f��uj�A�m�Uq�ƹt��x��n{�*�~����[���`H���兼����K�������C�� ֍�rf������Ձ����▕�6��B���,��Ͱ��{4��*����8������E:��۹��9�������5��|����0��@���p+��x����%���������P���������m��>�������  �  �vN=��M=��L=�4L=HsK=J�J=��I=�+I=
hH=ɣG=��F=,F=�RE=��D=��C=��B=�0B=fA=2�@=P�?=F�>=0>=�_==�<=�;=t�:=�:=99=`8=Y�7=��6=��5=��4=�4=�$3=�>2=rV1=�k0=:/=�.=n�-=>�,=m�+=Թ*=�)=/�(=�'=��&=%�%=m�$=c�#=��"=k!=�Q =f4=�=��=m�=�=�i=55=��=�=/=!:=��=E�=yQ=M�=�=*B=&�	=�w=a=��=�(=ð=�4=*i�<a�<+Q�<�9�<��<s��<��<���<�W�<��<���<��<�+�<���<[r�<��<��<e5�<*��<�J�<�ν<	O�<�˶<�D�<^��<�,�<Ҝ�<
�<�t�<^ݝ<�C�<ᨖ<�<n�<�΋<�.�<ҍ�<q�<��z<�Qs<�l<��d<@�]<�IV<�O<o�G<�@<�_9<�,2<��*<�#<�<^�<!q<�[<3M <͊�;a��;���;��;��;h'�;�{�;��;_`�;��m;�5S;�8;�b;2B;&��:�7�:�e\:xn�9.]�87蠹��2�15��4z���@�����&$��G;��%R��h���*����}��C���媻�f��_Ŀ�� ʻCԻ#޻O��$���0���Q�x������8����5a�*�!��%�� *�hE.��\2��f6��d:�rV>�e<B��F� �I���M��dQ�U�r�X��X\���_�xc��f��uj�:�m�Uq�ùt��x�o{�
�~����Y���MH���兼����L�������C��֍�rf�����ҁ����Җ��8��I���,��ְ��n4��-����8������@:��깤��8��z����5��j����0��F���j+��}����%���������S���������i��C�������  �  �vN=��M=��L=�4L=KsK=J�J=��I=�+I=hH=ģG=��F=.F=�RE=��D=��C=��B=�0B=	fA=0�@=M�?=J�>=0>=�_==�<=�;=p�:=�:=99=`8=\�7=�6=��5=��4=�4=�$3=�>2=zV1=�k0=</=�.=o�-=<�,=h�+=׹*=v�)=6�(=�'=��&=(�%=m�$=i�#=�"=
k!=�Q =e4=�=��=m�=�=�i=35=��=�=1=(:=��=L�=pQ=O�=�=(B=)�	=�w=d=��=�(=Ű=�4=3i�<a�<3Q�<�9�<��<k��<��<���<�W�<��<���<��<�+�<���<Yr�<��<���<\5�<'��<�J�<�ν<O�<�˶<�D�<S��<-�<Ҝ�<
�<�t�<fݝ<�C�<Ϩ�<�<n�<�΋<�.�<؍�<p�<��z<Rs<�l<�d<<�]<�IV<�O<p�G<��@<�_9<�,2<��*<
�#< �<\�<Gq<�[<NM <���;u��;���;��;��;5'�;�{�;��;�`�;��m;�5S;V�8;�b;�B;"��:�8�:�d\:Mm�9#`�8�꠹3�2�j5���y��WA����K&$�{G;�Q%R�I�h���.����}��C���媻uf���Ŀ�c ʻ9Ի�޻5��%���0���Q�]������K����6a�4�!���%�� *�\E.��\2��f6��d:�qV>�I<B��F��I���M��dQ��U�t�X��X\���_��wc� �f��uj�(�m�Uq���t��x��n{��~����[���\H���兼����9�������C��֍�wf������ځ��������=��M���,��Ͱ��y4������8��칡�=:��⹤��8�������5��x����0��C���e+��~����%���������E��� �����`��C�������  �  �vN=��M=��L=�4L=MsK=A�J=��I=�+I=hH=��G=��F=)F=�RE=��D=��C=��B=�0B=fA=3�@=J�?=J�>=0>=�_==�<=�;=m�:=�:=99=`8=e�7=�6=��5=��4=�4=�$3=�>2=wV1=�k0=A/=�.=u�-=@�,=f�+=�*=v�)=7�(=�'=��&=!�%=k�$=g�#=��"=k!=�Q =m4=�=��=u�= �=�i=/5=��=�=+= :=��=O�=pQ=[�=�=)B=0�	=�w=i=��=�(=°=�4=-i�<a�<6Q�<�9�<��<e��<
��<���<�W�<��<���<��<�+�<���<Sr�<��<���<S5�<8��<�J�<�ν<O�<�˶<�D�<J��<-�<͜�<
�<�t�<eݝ<�C�<Ө�<-�<�m�<�΋<�.�<э�<~�<��z<Rs<�l<��d<;�]<JV<�O<q�G<�@<}_9<�,2<��*<�#<(�<8�<.q<�[<MM <���;���;���;��;��;%'�;�{�;��;o`�; �m;[5S;O�8;Gb;dB;���:�8�:d\:�p�9�k�8E�;�2��5���y���@�����&$��G;��%R�(�h�V�G����}���B�� 檻f���Ŀ�[ ʻ]ԻF޻p��7���0��R�X������A����a�N�!� �%�!*�dE.��\2�g6��d:��V>�?<B��F���I���M��dQ��U���X�mX\���_��wc��f�vj�5�m�Uq���t��x��n{�'�~����H���^H���兼����F�������C��!֍�uf������䁒���▕�3��E���&,��Ȱ���4�� ����8������S:��㹤��8�������5�������0��@���k+��q����%���������L��� ������f��B�������  �  �vN=��M=��L=�4L=OsK=L�J=��I=�+I=
hH=ţG=��F=+F=�RE=��D=��C=��B=�0B=fA=6�@=L�?=F�>=0>=�_==��<=�;=n�:=�:=99=`8=\�7=��6=��5=��4=�4=�$3=�>2=sV1=l0=8/=�.=o�-==�,=e�+=Թ*=w�)=3�(=��'=��&=)�%=n�$=e�#=��"=k!=�Q =h4=�=��=n�=�=�i=65=��=�=2=(:=��=J�=pQ=L�=ݠ=)B=(�	=�w=_=��=�(=̰=�4=,i�<a�<*Q�<�9�<��<j��<���<���<�W�<��<���<��<�+�<���<Vr�<��<��<b5�<'��<�J�<�ν<O�<�˶<�D�<U��<�,�<Ӝ�<
�<�t�<kݝ<�C�<Ѩ�<�<n�<�΋<�.�<ԍ�<s�<��z< Rs<�l<��d<?�]<�IV<�O<w�G<��@<�_9<�,2<��*<��#</�<e�<7q<�[<3M <���;���;���;��;��;"'�;�{�;��;_`�;4�m;|5S;�8;�b;�B;c��:�8�:Yd\:�l�9�T�8W령P�2�*5��Uz���@����Q&$��F;��%R���h���*����}��C��
檻�f���Ŀ�u ʻԻ�޻4��$���0���Q�f������Y����2a�4�!�
�%�� *�gE.��\2��f6��d:�fV>�R<B��F�&�I���M��dQ��U�q�X��X\���_��wc���f��uj�6�m�Uq�ǹt��x��n{��~����^���\H���兼����=�������C��֍�jf�����ԁ����㖕�E��F���,��̰��w4��,����8��󹡼=:��ݹ���8�������5��{����0��C���h+��|����%���������M����������h��?�������  �  �yN=#�M=�L=i9L=fxK=�J=��I=u2I=\oH=��G=F�F=;"F=q\E=ܕD=��C=2C==B=�rA=ϧ@=��?=T?=�?>=1p==F�<=�;=c�:=J$:=�M9=u8=��7=5�6=��5=�5=�"4=�?3=�Z2=Vs1=�0=�/=��.=S�-=!�,=O�+=��*=n�)=�(=��'=��&=��%=C�$=$�#=��"=��!=�~ =�b=�B=�=��=�=;�=ag=R/=�=��=�m=�$=Y�=��=t/=��=v=�
=O�=d?=C�=�Z=6�=ze=`��<���<��<ٔ�<�s�<�K�<�<���</��<d�<��<���<Ir�<��<ɳ�<wL�<���<�n�<���<]~�<���<}�<���<�l�<�߯<�O�<���<'�<��<���<�X�<���<��<!z�<؋<65�<���<Z�<ߑz<�Hs<��k<c�d<Mp]<q*V<u�N<�G<�e@<�)9<U�1<��*<��#<(a<�:<<}�<d��;���;;��;���;7��;��;/"�;sk�;�ɐ;w;�;�k;U�P;f.6;��;1�;�-�:U��:��P:��9Q��7ul���c?�������������s~'�ߧ>�L�U�v.l��E��~Q���:��� �����Y$��=����˻��ջW�߻��點M����&�&���c����?b�^���#�n"���&���*�)�.�W3��7��;��>���B�бF�}J�o=N�n�Q�Z�U��AY���\�sj`���c��pg���j�Wn� �q� u��yx���{�O�p1��j҂��p��}��ʥ���<���ъ�Ld�����탏���w���~&��ɮ���5������G@���Û�<F���Ǟ�dH��Xȡ�zG��Ƥ�D��q����>��`����7�����D0��[���_(������� ��F������𖹼[��)�������  �  �yN=(�M=��L=c9L=hxK=�J=��I=o2I=YoH=��G=L�F=8"F=p\E=ەD=y�C=6C==B=�rA=ҧ@=��?=S?=�?>=9p==I�<=�;=Z�:=D$:=�M9=�u8=��7=-�6=��5=�5=�"4=�?3=�Z2=[s1=މ0=�/=�.=P�-=$�,=R�+=��*=b�)=�(=��'=��&=�%=?�$= �#=��"=��!=�~ =�b=�B=�=��=�=E�=bg=O/=�=��=�m=�$=[�=��=t/=��=v=�
=F�=g?=<�=�Z=C�=�e=]��<���<��<ǔ�<�s�<�K�<�<���<��<d�<��<���<Dr�<��<Ƴ�<zL�<���<�n�<���<B~�<���<}�<���<	m�<�߯<�O�<���<'�<��<���<�X�<���<�<)z�<$؋<+5�<���<[�<őz<�Hs<��k<��d<7p]<l*V<v�N<ƤG<�e@<�)9<l�1<Ӽ*<��#<2a<�:<5<g�<J��;���;n��;���;,��;��;�!�;�k�;Uɐ;�;�;,�k;N�P;[.6;s�;��;2.�:˘�::�P:���9��7�j��b?�����.���R�����}'�%�>���U��.l��E���Q���:��� ��룬�=$�������˻��ջ�߻_���M����&�����c����jb�����#�.n"�]�&���*�5�.�h3��7�i;���>���B��F�}J�d=N�f�Q�^�U��AY���\��j`���c��pg���j�Wn��q��u� zx���{�A�k1��s҂��p��v��å���<���ъ�Pd�����ꃏ�������v&��䮕��5������R@���Û�<F���Ǟ�pH��Dȡ�nG��Ƥ�
D�������>��W����7��%���I0��Z���l(��~���� ��/������򖹼[��7�������  �  �yN=+�M=��L=i9L=jxK=�J=��I=n2I=aoH=��G=L�F=7"F=p\E=�D=y�C=AC==B=�rA=ͧ@=��?=[?=�?>=6p==A�<=	�;=\�:=G$:=�M9=}u8=��7=)�6=��5=�5=�"4=�?3=�Z2=Xs1=ډ0=!�/=�.=R�-=!�,=M�+=��*=`�)=&�(=��'=��&=�%=D�$='�#=��"=��!=�~ =�b=�B=�=��=�=H�=[g=V/=�=��=�m=�$=a�=��=y/=��=v=�
=C�=o?=9�=�Z=6�=~e=]��<���<)��<���<�s�<�K�<�<���<��<&d�<��<���<?r�<��<˳�<oL�<��<�n�<���<G~�<���<'}�<���<m�<�߯<�O�<���<'�<���<���<�X�<���<�<z�<"؋<)5�<���<f�<��z<�Hs<��k<��d<4p]<|*V<��N<��G<�e@<�)9<u�1<Ӽ*<��#<:a<�:<-<c�<���;i��;j��;y��;3��;(�;�!�;�k�;1ɐ;�;�;�k;Q�P;�.6;O�;��;$-�:h��:��P:���9��78m���a?�(���<������"~'��>�"�U�/l��E���Q���:��� �����$������Ի˻��ջG�߻j�黚M�g��� &�����c����Kb�w���#�Kn"�R�&���*��.�I3��7�z;��>���B��F�}J�t=N�v�Q�S�U��AY�u�\��j`���c��pg���j�Wn��q��u�4zx���{�V�o1��h҂��p��k��ӥ���<���ъ�@d���������������^&��߮���5������W@���Û�FF���Ǟ�nH��Hȡ�G�� Ƥ��C�������>��d����7��'���G0��O���o(������� ��7������ꖹ�U��>�������  �  �yN=$�M=��L=f9L=gxK=�J=��I=p2I=]oH=��G=L�F=@"F=o\E=ܕD=x�C=7C==B=�rA=Χ@=��?=T?=�?>=9p==F�<=�;=]�:=G$:=�M9=u8=��7=.�6=��5=�5=�"4=�?3=�Z2=\s1=ى0=�/=�.=S�-= �,=N�+=��*=c�)=�(=��'=��&=�%=@�$='�#=��"=��!=�~ =�b=�B=�=��=�=G�=]g=V/=�=��=�m=�$=Y�=��=s/=��=v=�
=F�=f?=8�=�Z=>�=�e=b��<���<��<ǔ�<�s�<�K�<�<���<��<d�<��<���<Gr�<��<г�<rL�<	��<�n�<���<A~�<���<}�<���<	m�<�߯<�O�<���<'�<
��<���<�X�<���<��<z�<؋<15�<���<Z�<őz<�Hs<��k<��d<;p]<b*V<q�N<ͤG<�e@<�)9<Z�1<޼*<��#</a<�:</<h�<k��;y��;m��;���;'��;��;�!�;�k�;Dɐ;�;�;��k;z�P;l.6;��;Ö;�-�:���:��P:���9���7ul���b?�~���8���������}'�Z�>��U�'/l��E���Q���:��� �����M$�������˻��ջ�߻f�黹M�m���&�����c����]b�����#�+n"�S�&���*��.�b3��7�i;��>���B���F�}J�t=N�r�Q�V�U��AY���\��j`���c��pg���j�Wn�$�q��u�zx���{�P�v1��l҂��p��{��˥���<���ъ�Pd�����򃏼������s&��宕��5������D@���Û�CF���Ǟ�oH��Iȡ�sG��Ƥ�D�������>��a����7�����L0��[���l(������� ��4����������]��3�������  �  �yN=!�M=��L=f9L=hxK=�J=��I=s2I=XoH=��G=F�F=;"F=s\E=�D=��C=:C==B=�rA=ͧ@=��?=P?=�?>=3p==I�<=�;=_�:=G$:=�M9=�u8=��7=0�6=��5=�5=�"4=�?3=�Z2=Qs1=މ0=�/=�.=M�-=�,=T�+=��*=k�)=�(=��'=��&=�%=?�$=&�#=��"=��!=�~ =�b=�B=�=��=�=A�=cg=V/=�=��=�m=�$=X�=��=p/=��=v=�
=I�=f?==�=�Z=;�=|e=P��<���<��<̔�<�s�<�K�<�<���<&��<d�<��<���<Nr�<��<׳�<tL�<���<�n�<���<V~�<���<#}�<���<�l�<�߯<�O�<���<'�<
��<���<�X�<���<��<.z�<؋</5�<���<^�<z<�Hs<��k<^�d<1p]<r*V<u�N<ФG<�e@<�)9<N�1<�*<��#<0a<�:<%<v�<B��;»�;@��;���;G��;�;"�;�k�;uɐ;�;�;�k;��P;7.6;��;e�;:.�:���:��P:���9��7)i���c?�,���a������<�W~'�|�>���U��.l��E���Q���:��� ��֣��b$��V����˻��ջA�߻^�黾M�r����%����c����Cb�g���#�n"�n�&���*��.�n3��7��;���>���B�ݱF�#}J�_=N�o�Q�p�U��AY���\��j`���c��pg���j�0Wn��q��u�zx���{�;�q1��p҂��p��{��¥���<���ъ�Wd�����������~���m&��Ю���5������I@���Û�0F���Ǟ�hH��Jȡ�tG�� Ƥ�D��y����>��S����7��!���G0��V���n(������� ��H�������[��1�������  �  �yN=#�M=��L=g9L=lxK=�J=��I=u2I=[oH=��G=J�F=?"F=q\E=��D=y�C=<C==B=�rA=Ч@=��?=U?=�?>=2p==I�<=�;=^�:=G$:=�M9=~u8=��7=-�6=��5=�5=�"4=�?3=�Z2=Us1=߉0=�/=�.=S�-=�,=M�+=��*=g�)=�(=��'=��&=�%=B�$=&�#=��"=��!=�~ =�b=�B=�=��=�=G�=`g=U/=�=��=�m=�$=[�=��=r/=��=v=�
=E�=e?==�=�Z=8�=~e=T��<���<��<Ɣ�<�s�<�K�<�<���<"��<d�<��<���<Mr�<��<ѳ�<vL�<��<�n�<���<G~�<���<#}�<���<m�<�߯<�O�<¼�<'�<���<���<�X�<���<��<z�<؋<15�<z��<Y�<Ƒz<�Hs<��k<x�d<5p]<h*V<]�N<ɤG<�e@<�)9<V�1<ܼ*<��#<@a<�:<#<��<[��;���;d��;���;:��;	�;�!�;�k�;Vɐ;�;�;�k;��P;�.6;��;U�;..�:S��:k�P:��9��7�l���a?�������������~'���>�M�U��.l��E���Q���:��� �����O$��t����˻��ջ_�߻Z�黥M�t���&�����c����Mb�v���#�(n"�R�&���*��.�]3��7��;���>���B��F�}J�u=N�u�Q�S�U��AY���\��j`���c��pg���j�&Wn��q�	 u�zx���{�S�s1��n҂��p��r�������<���ъ�Kd��
����	������h&��߮���5������C@���Û�2F���Ǟ�aH��Kȡ�G���Ť� D�������>��c����7�����R0��\���k(������� ��;������󖹼g��5�������  �  �yN=+�M=��L=c9L=cxK=�J=��I=q2I=^oH=��G=K�F=?"F=o\E=�D=|�C=DC==B=�rA=ϧ@=��?=V?=�?>==p==G�<=��;=Z�:=G$:=�M9={u8=��7=*�6=��5=�5=�"4=�?3=�Z2=Xs1=։0=�/=�.=O�-=�,=L�+=��*=d�)=�(=��'=��&=�%==�$=)�#=��"=��!=�~ =�b=�B=�=��=�=J�=]g=W/=�=��=�m=�$=T�=��=v/=��=v=�
=A�=f?=4�=�Z=7�=|e=Q��<���<��<���<�s�<�K�<�<���<��<
d�<��< ��<Fr�<��<ҳ�<tL�<	��<�n�<���<J~�<���<!}�<���<m�<�߯<�O�<���<'�<��<���<�X�<���<�<z�<؋<(5�<|��<Y�<��z<�Hs<��k<��d<p]<d*V<f�N<��G<�e@<�)9<u�1<ּ*<��#<a<�:<D<o�<y��;���;g��;���;.��;G�;�!�;l�;Aɐ;�;�;�k;��P;�.6;��;�;.�:/��:��P:��9[�7$n��Yb?�󌐺����~��T�"~'�§>��U�Z/l��E���Q���:��� �����$������7�˻��ջ�߻G���M�Z���&�����c����Db�s���#�5n"�G�&���*��.�j3��7�h;��>���B���F�	}J�v=N���Q�d�U��AY���\��j`���c��pg���j�*Wn�)�q��u�0zx���{�e�n1��j҂��p�����ǥ���<���ъ�Md���������������\&��ܮ���5������F@���Û�:F���Ǟ�mH��?ȡ�sG��
Ƥ�
D�������>��g����7��(���P0��[���{(������� ��6����������b��<�������  �  �yN="�M=��L=k9L=gxK=�J=��I=t2I=_oH=��G=H�F=A"F=u\E=�D=|�C=?C==B=�rA=ϧ@=��?=V?=�?>=5p==I�<=�;=c�:=A$:=�M9=�u8=��7=-�6=��5=�5=�"4=�?3=�Z2=Ss1=ى0=�/=�.=M�-=�,=O�+=��*=h�)="�(=��'=��&=�%=B�$=,�#=��"=��!=�~ =�b=�B=�=��=�=G�=bg=[/=�=��=�m=�$=[�=��=k/=��=v=�
=C�=c?=7�=�Z=6�=ye=O��<���<��<�<�s�<�K�<�<v��<)��<d�<��<���<Gr�<��<۳�<wL�<��<�n�<���<L~�<���<*}�<���<m�<�߯<�O�<���<'�<��<���<�X�<���<��<!z�<؋<)5�<}��<Y�<��z<�Hs<��k<b�d<p]<b*V<e�N<ĤG<�e@<�)9<Q�1<ϼ*<��#<,a<�:<'<y�<���;���;T��;Ѳ�;a��;;�;�!�;�k�;�ɐ;�;�;�k;��P;�.6;��;��;W.�:�:��P:���9���7�j��Oc?�m�������*��C�m~'�ѧ>�n�U�(/l��E���Q���:��� ������z$��h����˻��ջ0�߻T�黧M�?����%�����c����Bb�q���#�n"�P�&���*��.�[3��7�x;���>���B��F�3}J�q=N�v�Q�m�U��AY���\��j`���c��pg���j�-Wn��q� u�#zx���{�M�t1��z҂��p��x��¥���<���ъ�Ld����샏���z���c&��ٮ���5������>@���Û�3F���Ǟ�gH��Jȡ�rG��Ƥ��C�������>��`����7��'���P0��\���w(������� ��F����������b��7�������  �  �yN=#�M=��L=h9L=gxK=�J=��I={2I=ZoH=��G=N�F=C"F=t\E=ߕD=��C=9C==B=�rA=ԧ@=��?=T?=�?>=2p==M�<=�;=_�:=F$:=�M9=~u8=��7=/�6=��5=�5=�"4=�?3=�Z2=Ps1=݉0=�/=�.=P�-=�,=O�+=��*=g�)=�(=��'=��&=�%=F�$=$�#=��"=��!=�~ =�b=�B=�=��=�=I�=eg=T/=�=��=�m=�$=W�=��=n/=��=v=�
=E�=[?=;�=�Z=;�={e=H��<���<��<Ɣ�<�s�<�K�<�<��<!��<d�<��<���<Vr�<��<ҳ�<}L�<��<�n�<���<U~�<���<'}�<���<m�<�߯<�O�<˼�<'�<��<���<�X�<���<��< z�<؋<05�<w��<M�<��z<�Hs<��k<h�d<*p]<N*V<W�N<ͤG<�e@<�)9<T�1<޼*<��#<-a<�:<!<��<U��;ͻ�;���;��;Y��;�;"�;�k�;ɐ;�;�;`�k;��P;�.6;@�;g�;�.�:���:��P:���9���7sl���c?�C���?���f��W�A~'�g�>���U��.l� F���Q���:��������_$��r����˻��ջ<�߻B�黀M�}����%�����c����Db�j���#�n"�K�&�x�*��.�Q3��7�};���>���B��F�%}J�r=N���Q�f�U��AY���\��j`���c��pg���j�;Wn��q� u�zx���{�Y�u1��q҂��p��~�������<���ъ�Ld�����惏���|���m&��Ѯ���5������<@���Û�-F���Ǟ�WH��Jȡ�pG�� Ƥ�D�������>��`����7�� ���U0��h���o(������� ��B������ ���j��2�������  �  �yN=&�M=��L=h9L=fxK=�J=��I=t2I=^oH=��G=N�F=>"F=w\E=�D=��C=DC==B=�rA=ѧ@=��?=W?=�?>=5p==H�<=�;=]�:=G$:=�M9={u8=��7=%�6=��5=�5=�"4=�?3=�Z2=Ms1=؉0=�/=�.=M�-=�,=L�+=��*=b�)=�(=��'=��&=�%=B�$=*�#=��"=��!=�~ =�b=�B=�=��=�=I�=bg=Z/=�=��=�m=�$=X�=��=u/=��=v=�
=?�=c?=6�=�Z=2�=ue=F��<���<��<���<�s�<�K�<�<���<��<d�<��<���<Ir�<��<ٳ�<yL�<
��<�n�<���<X~�<���<2}�<���<m�<�߯<�O�<���<'�<��<���<�X�<���<�<z�<؋<"5�<|��<Y�<��z<�Hs<��k<S�d<p]<d*V<h�N<��G<�e@<�)9<`�1<׼*<��#<)a<�:<+<}�<w��;���;~��;���;s��;V�;("�;l�;~ɐ;�;�;@�k;��P;�.6;��;��;8.�:ޘ�:i�P:A��9E��7�m���b?�s���g���4��k��~'���>���U�4/l��E���Q���:��� �����&$�������˻��ջ'�߻^�黣M�O����%�����c����/b�[��}#�,n"�J�&���*��.�Y3��7�t;��>���B���F�}J�|=N�{�Q�j�U��AY���\��j`���c��pg���j�>Wn� �q� u�@zx���{�[�v1��k҂��p��y��ȥ���<���ъ�Id�� ���ꃏ�������V&��ͮ���5������G@���Û�1F���Ǟ�eH��Hȡ�rG��Ƥ�D�������>��h����7��-���P0��\���z(������� ��M����������a��D�������  �  �yN=%�M=��L=k9L=hxK=�J=��I=r2I=coH=��G=S�F=D"F=v\E=�D=v�C=BC==B=�rA=ӧ@=��?=Z?=�?>=>p==E�<=�;=^�:=A$:=�M9=|u8=��7=$�6=��5=�5=�"4=�?3=�Z2=Xs1=Ӊ0=�/=�.=K�-=%�,=H�+=��*=^�)=&�(=��'=��&=�%=A�$=-�#=��"=��!=�~ =�b=�B=�=��=�=Q�=^g=[/=�=��=�m=�$=`�=��=p/=��=v=�
==�=b?=/�=�Z=5�=ze=T��<���<��<���<�s�<�K�<�<z��<��<"d�<��<��<Gr�<��<׳�<xL�<��<�n�<���<@~�<���<-}�<���<m�<�߯<�O�<���<!'�<
��<���<�X�<���<�<z�<#؋<5�<z��<M�<��z<�Hs<��k<q�d<p]<E*V<e�N<��G<�e@<�)9<]�1<��*<��#<0a<�:<E<t�<���;���;���;��;e��;H�;�!�;�k�;vɐ;<�;T�k;��P;�.6;��;&�;�-�:p��:��P:��9���7im��0b?�����2���h���/~'�ԧ>��U��/l��E���Q���:��� ��3���I$������ϻ˻��ջ�߻K�黭M�5���&�����c����Fb�z���#�$n"�(�&���*���.�^3��7�^;��>���B��F�}J��=N�`�Q�m�U��AY���\��j`���c��pg���j�!Wn�F�q��u�Czx���{�P�v1��v҂��p��l��Υ���<���ъ�Gd�����냏��������]&��宕��5������=@���Û�<F���Ǟ�iH��>ȡ�sG��Ƥ��C�������>��o����7��2���S0��g���}(������� ��>���������b��H�������  �  �yN='�M=��L=h9L=cxK=�J=��I=y2I=boH=��G=N�F=A"F=w\E=�D=��C=FC==B=�rA=ӧ@=��?=[?=�?>=:p==E�<= �;=^�:=I$:=�M9=zu8=��7=*�6=��5=�5=�"4=�?3=�Z2=Ks1=ى0=�/=�.=G�-=�,=J�+=��*=f�)= �(=��'=��&=
�%=F�$=+�#=��"=��!=�~ =�b=�B=�=��=�=I�=ag=Y/=�=��=�m=�$=Y�=��=t/=��=v=�
=D�=_?=5�=�Z=0�=qe=D��<���<��<���<�s�<�K�<�<���<��<d�<��<���<Qr�<��<ӳ�<wL�<	��<�n�<���<^~�<���</}�<���<m�<�߯<�O�<Ƽ�< '�<��<���<�X�<���<�<z�<؋< 5�<���<I�<��z<~Hs<��k<O�d<p]<F*V<m�N<��G<�e@<�)9<e�1<߼*<��#<a<�:<<<��<���;���;���;Ҳ�;m��;l�;@"�;l�;�ɐ;�;�;U�k;��P;/6;!�;�;�-�:n��:��P:��9��7	n��*d?�ӌ��[������v��~'�	�>�ٍU�/l�	F���Q���:��� ��"���,$��w�����˻��ջ7�߻5�黃M�E����%�����c����b�I���#�n"�I�&���*��.�K3��7�s;��>���B��F�}J��=N���Q���U��AY���\��j`���c��pg���j�AWn�1�q� u�+zx���{�`�s1��h҂��p��~��˥���<���ъ�Ad�����냏���|���V&��Ǯ���5������B@���Û�4F���Ǟ�]H��?ȡ�wG��
Ƥ� D�������>��j����7��/���K0��k���u(������� ��O���������_��A�������  �  �yN=�M=��L=e9L=jxK=��J=��I=u2I=]oH=��G=M�F=C"F=|\E=��D=z�C=>C==B=�rA=֧@=��?=X?=�?>=3p==Q�<=�;=\�:=C$:=�M9=�u8=��7=)�6=��5=�5=�"4=�?3=�Z2=Hs1=��0=�/=�.=I�-=�,=L�+=��*=b�)=�(=��'=��&=�%=B�$=(�#=��"=��!=�~ =�b=�B=�=��=�=F�=kg=X/=�=��=�m=�$=W�=��=k/=��=v=�
=C�=V?=<�=�Z==�={e=C��<���<���<���<�s�<�K�< �<y��<��<d�<��<���<Jr�<��<ڳ�<�L�<��<�n�<���<G~�<���<8}�<���<
m�<�<�O�<���<'�<��<���<�X�<���<��<z�<؋< 5�<z��<G�<��z<tHs<��k<L�d<%p]<K*V<V�N<��G<�e@<�)9<?�1<Ҽ*<��#<9a< ;<'<��<l��;��;~��;��;���;�;�!�;�k�;�ɐ;�;�;��k;�P;�.6;��;y�;o/�:���:S�P:S��9���7Pk��,c?�����g���<��u�R~'�&�>��U��.l�@F���Q���:��� �����r$�������˻��ջ�߻I�黠M�`����%�����c����Pb�|���#�n"�S�&�_�*��.�T3��7�p;���>���B���F�2}J��=N�p�Q�|�U��AY���\��j`��c��pg���j�AWn��q�, u�/zx���{�K��1��w҂��p��|�������<���ъ�Fd����݃����n���b&��ޮ���5������;@���Û�$F���Ǟ�dH��Hȡ�jG���Ť�D�������>��a����7��/���R0��n���m(������� ��P���������j��A�������  �  �yN='�M=��L=h9L=cxK=�J=��I=y2I=boH=��G=N�F=A"F=w\E=�D=��C=FC==B=�rA=ӧ@=��?=[?=�?>=:p==E�<= �;=^�:=I$:=�M9=zu8=��7=*�6=��5=�5=�"4=�?3=�Z2=Ks1=ى0=�/=�.=G�-=�,=J�+=��*=f�)= �(=��'=��&=
�%=F�$=+�#=��"=��!=�~ =�b=�B=�=��=�=I�=ag=Y/=�=��=�m=�$=Y�=��=t/=��=v=�
=D�=_?=6�=�Z=0�=qe=D��<���<��<���<�s�<�K�<�<���<��<d�<��<���<Qr�<��<ӳ�<wL�<	��<�n�<���<^~�<���</}�<���<m�<�߯<�O�<Ƽ�< '�<��<���<�X�<���<�<z�<؋< 5�<���<I�<��z<~Hs<��k<O�d<p]<F*V<m�N<��G<�e@<�)9<e�1<߼*<��#<a<�:<<<��<���;���;���;Ҳ�;m��;l�;@"�;l�;�ɐ;�;�;T�k;��P;/6; �;�;�-�:m��:��P:{��9��7n��-d?�Ԍ��\������w��~'�
�>�ڍU�/l�	F���Q���:��� ��#���,$��w�����˻��ջ7�߻5�黃M�E����%�����c����b�I���#�n"�I�&���*��.�K3��7�s;��>���B��F�}J��=N���Q���U��AY���\��j`���c��pg���j�AWn�1�q� u�+zx���{�`�s1��h҂��p��~��˥���<���ъ�Ad�����냏���|���V&��Ǯ���5������B@���Û�4F���Ǟ�]H��?ȡ�wG��
Ƥ� D�������>��j����7��/���K0��k���u(������� ��O���������_��A�������  �  �yN=%�M=��L=k9L=hxK=�J=��I=r2I=coH=��G=S�F=D"F=v\E=�D=v�C=BC==B=�rA=ӧ@=��?=Z?=�?>=>p==E�<=�;=^�:=A$:=�M9=|u8=��7=$�6=��5=�5=�"4=�?3=�Z2=Xs1=Ӊ0=�/=�.=K�-=%�,=H�+=��*=^�)=&�(=��'=��&=�%=A�$=-�#=��"=��!=�~ =�b=�B=�=��=�=Q�=^g=[/=�=��=�m=�$=`�=��=p/=��=v=�
==�=b?=/�=�Z=5�=ze=T��<���<��<���<�s�<�K�<�<z��<��<"d�<��<��<Gr�<��<׳�<xL�<��<�n�<���<@~�<���<-}�<���<m�<�߯<�O�<���<!'�<
��<���<�X�<���<�<z�<#؋<5�<z��<M�<��z<�Hs<��k<r�d<p]<E*V<e�N<��G<�e@<�)9<]�1<��*<��#<0a<�:<E<t�<���;���;���;��;e��;H�;�!�;�k�;vɐ;<�;T�k;��P;�.6;��;%�;�-�:n��:��P:u��9���7sm��4b?�����4���j���0~'�է>��U��/l��E���Q���:��� ��4���J$������ϻ˻��ջ�߻K�黭M�5���&�����c����Fb�z���#�$n"�(�&���*���.�^3��7�^;��>���B��F�}J��=N�`�Q�m�U��AY���\��j`���c��pg���j�!Wn�F�q��u�Dzx���{�P�v1��v҂��p��l��Υ���<���ъ�Gd�����냏��������]&��宕��5������=@���Û�<F���Ǟ�iH��>ȡ�sG��Ƥ��C�������>��o����7��2���S0��g���}(������� ��>���������b��H�������  �  �yN=&�M=��L=h9L=fxK=�J=��I=t2I=^oH=��G=N�F=>"F=w\E=�D=��C=DC==B=�rA=ѧ@=��?=W?=�?>=5p==H�<=�;=]�:=G$:=�M9={u8=��7=%�6=��5=�5=�"4=�?3=�Z2=Ms1=؉0=�/=�.=M�-=�,=L�+=��*=b�)=�(=��'=��&=�%=B�$=*�#=��"=��!=�~ =�b=�B=�=��=�=I�=bg=Z/=�=��=�m=�$=X�=��=u/=��=v=�
=?�=c?=6�=�Z=2�=ue=F��<���<��<���<�s�<�K�<�<���<��<d�<��<���<Ir�<��<ڳ�<yL�<
��<�n�<���<X~�<���<2}�<���<m�<�߯<�O�<���<'�<��<���<�X�<���<�<z�<؋<"5�<|��<Y�<��z<�Hs<��k<S�d<p]<d*V<h�N<��G<�e@<�)9<`�1<׼*<��#<*a<�:<+<}�<w��;���;~��;���;s��;V�;'"�;l�;~ɐ;�;�;?�k;��P;�.6;��;��;5.�:ۘ�:b�P:4��9m��7�m���b?�v���j���8��l��~'��>���U�6/l��E���Q���:��� �����&$�������˻��ջ'�߻^�黣M�O����%�����c����/b�[��}#�,n"�J�&���*��.�Y3��7�t;��>���B���F�}J�|=N�{�Q�j�U��AY���\��j`���c��pg���j�>Wn� �q� u�@zx���{�[�v1��k҂��p��y��ȥ���<���ъ�Id�� ���ꃏ�������V&��ͮ���5������G@���Û�1F���Ǟ�eH��Hȡ�rG��Ƥ�D�������>��h����7��-���P0��\���z(������� ��M����������a��D�������  �  �yN=#�M=��L=h9L=gxK=�J=��I={2I=ZoH=��G=N�F=C"F=t\E=ߕD=��C=9C==B=�rA=ԧ@=��?=T?=�?>=2p==M�<=�;=_�:=F$:=�M9=~u8=��7=/�6=��5=�5=�"4=�?3=�Z2=Ps1=݉0=�/=�.=P�-=�,=O�+=��*=g�)=�(=��'=��&=�%=F�$=$�#=��"=��!=�~ =�b=�B=�=��=�=I�=eg=T/=�=��=�m=�$=W�=��=n/=��=v=�
=E�=\?=;�=�Z=;�={e=H��<���<��<Ɣ�<�s�<�K�<�<��<!��<d�<��<���<Vr�<��<ҳ�<}L�<��<�n�<���<U~�<���<'}�<���<m�<�߯<�O�<˼�<'�<��<���<�X�<���<��< z�<؋<05�<w��<M�<��z<�Hs<��k<h�d<*p]<N*V<W�N<ͤG<�e@<�)9<T�1<޼*<��#<-a<�:<!<��<U��;ͻ�;���;��;Y��;�;"�;�k�;~ɐ;�;�;_�k;��P;�.6;>�;f�;�.�:���:��P:~��9���7�l���c?�G���C���j��Y�B~'�i�>���U��.l�!F���Q���:��������`$��s����˻��ջ=�߻B�黁M�~����%�����c����Db�j���#�n"�K�&�x�*��.�Q3��7�};���>���B��F�%}J�r=N���Q�f�U��AY���\��j`���c��pg���j�;Wn��q� u�zx���{�Y�u1��q҂��p��~�������<���ъ�Ld�����惏���|���m&��Ѯ���5������<@���Û�-F���Ǟ�WH��Jȡ�pG�� Ƥ�D�������>��`����7�� ���U0��h���o(������� ��B������ ���j��2�������  �  �yN="�M=��L=k9L=gxK=�J=��I=t2I=_oH=��G=H�F=A"F=u\E=�D=|�C=?C==B=�rA=ϧ@=��?=V?=�?>=5p==I�<=�;=c�:=A$:=�M9=�u8=��7=-�6=��5=�5=�"4=�?3=�Z2=Ss1=ى0=�/=�.=M�-=�,=O�+=��*=h�)="�(=��'=��&=�%=B�$=,�#=��"=��!=�~ =�b=�B=�=��=�=G�=bg=[/=�=��=�m=�$=[�=��=k/=��=v=�
=C�=c?=7�=�Z=6�=ye=P��<���<��<Ô�<�s�<�K�<�<w��<)��<d�<��<���<Gr�<��<۳�<wL�<��<�n�<���<L~�<���<*}�<���<m�<�߯<�O�<���<'�<��<���<�X�<���<��<!z�<؋<)5�<}��<Y�<��z<�Hs<��k<b�d<p]<b*V<e�N<ĤG<�e@<�)9<R�1<ϼ*<��#<,a<�:<'<z�<���;���;U��;Ѳ�;a��;;�;�!�;�k�;�ɐ;�;�;�k;��P;�.6;��;��;S.�::��P:���9���7�j��Xc?�r�������.��E�o~'�ӧ>�p�U�*/l��E���Q���:��� ������{$��i����˻��ջ0�߻T�黨M�@����%�����c����Bb�q���#�n"�P�&���*��.�[3��7�x;���>���B��F�3}J�q=N�v�Q�m�U��AY���\��j`���c��pg���j�-Wn��q� u�#zx���{�M�t1��z҂��p��x��¥���<���ъ�Ld����샏���z���c&��ٮ���5������>@���Û�3F���Ǟ�gH��Jȡ�rG��Ƥ��C�������>��`����7��'���P0��\���w(������� ��F����������b��7�������  �  �yN=+�M=��L=c9L=cxK=�J=��I=q2I=^oH=��G=K�F=?"F=o\E=�D=|�C=DC==B=�rA=ϧ@=��?=V?=�?>==p==G�<=��;=Z�:=G$:=�M9={u8=��7=*�6=��5=�5=�"4=�?3=�Z2=Xs1=։0=�/=�.=O�-=�,=L�+=��*=d�)=�(=��'=��&=�%==�$=)�#=��"=��!=�~ =�b=�B=�=��=�=J�=]g=W/=�=��=�m=�$=T�=��=v/=��=v=�
=A�=f?=4�=�Z=7�=}e=R��<���<��<���<�s�<�K�<�<���<��<d�<��< ��<Fr�<��<ҳ�<tL�<	��<�n�<���<J~�<���<!}�<���<m�<�߯<�O�<���<'�<
��<���<�X�<���<�<z�<؋<(5�<|��<Y�<��z<�Hs<��k<��d<p]<d*V<f�N<��G<�e@<�)9<u�1<ּ*<��#<a<�:<D<o�<z��;���;g��;���;.��;G�;�!�;l�;@ɐ;�;�;�k;��P;�.6;��;�;�-�:+��:{�P:��9(�77n��bb?������������V�$~'�ħ>��U�\/l��E���Q���:��� �����$������7�˻��ջ�߻G���M�Z���&�����c����Db�s���#�5n"�G�&���*��.�j3��7�h;��>���B���F�	}J�v=N���Q�d�U��AY���\��j`���c��pg���j�*Wn�)�q��u�0zx���{�e�n1��j҂��p�����ǥ���<���ъ�Md���������������\&��ܮ���5������F@���Û�:F���Ǟ�mH��?ȡ�sG��
Ƥ�
D�������>��g����7��(���P0��[���{(������� ��6����������b��<�������  �  �yN=#�M=��L=g9L=lxK=�J=��I=u2I=[oH=��G=J�F=?"F=q\E=��D=y�C=<C==B=�rA=Ч@=��?=U?=�?>=2p==I�<=�;=^�:=G$:=�M9=~u8=��7=-�6=��5=�5=�"4=�?3=�Z2=Us1=߉0=�/=�.=S�-=�,=M�+=��*=g�)=�(=��'=��&=�%=B�$=&�#=��"=��!=�~ =�b=�B=�=��=�=G�=`g=U/=�=��=�m=�$=[�=��=r/=��=v=�
=F�=e?==�=�Z=8�=~e=T��<���<��<Ɣ�<�s�<�K�<�<���<#��<d�<��<���<Mr�<��<ѳ�<vL�<��<�n�<���<G~�<���<#}�<���<m�<�߯<�O�<���<'�<���<���<�X�<���<��<z�<؋<15�<z��<Y�<Ƒz<�Hs<��k<x�d<5p]<h*V<]�N<ɤG<�e@<�)9<V�1<ܼ*<��#<@a<�:<$<��<[��;���;d��;���;:��;	�;�!�;�k�;Uɐ;�;�;�k;��P;�.6;��;S�;*.�:O��:b�P:���9���7�l��b?�������������~'���>�O�U��.l��E���Q���:��� �����P$��u����˻��ջ_�߻[�黥M�t���&�����c����Mb�v���#�(n"�R�&���*��.�]3��7��;���>���B��F�}J�u=N�u�Q�S�U��AY���\��j`���c��pg���j�&Wn��q�	 u�zx���{�S�s1��n҂��p��r�������<���ъ�Kd��
����	������h&��߮���5������C@���Û�2F���Ǟ�aH��Kȡ�G���Ť� D�������>��c����7�����R0��\���k(������� ��;������󖹼g��5�������  �  �yN=!�M=��L=f9L=hxK=�J=��I=s2I=XoH=��G=F�F=;"F=s\E=�D=��C=:C==B=�rA=ͧ@=��?=P?=�?>=3p==I�<=�;=_�:=G$:=�M9=�u8=��7=0�6=��5=�5=�"4=�?3=�Z2=Qs1=މ0=�/=�.=M�-=�,=T�+=��*=k�)=�(=��'=��&=�%=?�$=&�#=��"=��!=�~ =�b=�B=�=��=�=A�=cg=V/=�=��=�m=�$=X�=��=p/=��=v=�
=I�=f?==�=�Z=;�=|e=P��<���<��<͔�<�s�<�K�<�<���<&��<d�<��<���<Nr�<��<׳�<tL�<���<�n�<���<V~�<���<#}�<���<�l�<�߯<�O�<���<'�<	��<���<�X�<���<��<.z�<؋</5�<���<^�<z<�Hs<��k<^�d<2p]<r*V<u�N<ФG<�e@<�)9<N�1<�*<��#<1a<�:<&<v�<C��;û�;@��;���;G��;�;"�;�k�;tɐ;�;�;�k;��P;6.6;��;c�;6.�:���:��P:���9
��7:i���c?�0���e������>�Y~'�~�>���U��.l��E���Q���:��� ��֣��b$��V����˻��ջB�߻_�黾M�r����%����c����Cb�g���#�n"�n�&���*��.�n3��7��;���>���B�ݱF�#}J�_=N�o�Q�p�U��AY���\��j`���c��pg���j�0Wn��q��u�zx���{�;�q1��p҂��p��{��¥���<���ъ�Wd�����������~���m&��Ю���5������I@���Û�0F���Ǟ�hH��Jȡ�tG�� Ƥ�D��y����>��S����7��!���G0��V���n(������� ��H�������[��1�������  �  �yN=$�M=��L=f9L=gxK=�J=��I=p2I=]oH=��G=L�F=@"F=o\E=ܕD=x�C=7C==B=�rA=Χ@=��?=T?=�?>=9p==F�<=�;=]�:=G$:=�M9=u8=��7=.�6=��5=�5=�"4=�?3=�Z2=\s1=ى0=�/=�.=S�-= �,=N�+=��*=c�)=�(=��'=��&=�%=@�$='�#=��"=��!=�~ =�b=�B=�=��=�=G�=]g=V/=�=��=�m=�$=Y�=��=s/=��=v=�
=F�=f?=8�=�Z=>�=�e=b��<���<��<ǔ�<�s�<�K�<�<���<��<d�<��<���<Gr�<��<г�<rL�<	��<�n�<���<A~�<���<}�<���<	m�<�߯<�O�<���<'�<
��<���<�X�<���<��<z�<؋<15�<���<Z�<őz<�Hs<��k<��d<;p]<b*V<q�N<ͤG<�e@<�)9<[�1<޼*<��#</a<�:</<i�<k��;y��;m��;���;'��;��;�!�;�k�;Dɐ;�;�;��k;y�P;k.6;��;;�-�:���:��P:��9���7�l���b?�����<���������}'�[�>��U�(/l��E���Q���:��� �����M$�������˻��ջ�߻g�黹M�m���&�����c����]b�����#�+n"�S�&���*��.�b3��7�i;��>���B���F�}J�t=N�r�Q�V�U��AY���\��j`���c��pg���j�Wn�$�q��u�zx���{�P�v1��l҂��p��{��˥���<���ъ�Pd�����򃏼������s&��宕��5������D@���Û�CF���Ǟ�oH��Iȡ�sG��Ƥ�D�������>��a����7�����L0��[���l(������� ��4����������]��3�������  �  �yN=+�M=��L=i9L=jxK=�J=��I=n2I=aoH=��G=L�F=7"F=p\E=�D=y�C=AC==B=�rA=ͧ@=��?=[?=�?>=6p==A�<=	�;=\�:=G$:=�M9=}u8=��7=)�6=��5=�5=�"4=�?3=�Z2=Xs1=ډ0=!�/=�.=R�-=!�,=M�+=��*=`�)=&�(=��'=��&=�%=D�$='�#=��"=��!=�~ =�b=�B=�=��=�=H�=[g=V/=�=��=�m=�$=a�=��=y/=��=v=�
=D�=o?=9�=�Z=6�=~e=]��<���<)��<���<�s�<�K�<�<���<��<&d�<��<���<?r�<��<˳�<oL�<��<�n�<���<G~�<���<'}�<���<m�<�߯<�O�<���<'�<���<���<�X�<���<�<z�<"؋<)5�<���<f�<��z<�Hs<��k<��d<4p]<|*V<��N<��G<�e@<�)9<u�1<Լ*<��#<:a<�:<-<c�<���;i��;j��;z��;3��;(�;�!�;�k�;1ɐ;�;�;�k;P�P;�.6;N�;��;"-�:f��:��P:���9�7Am���a?�+���?������#~'��>�#�U� /l��E���Q���:��� �����$������ջ˻��ջG�߻j�黚M�h��� &���� d����Kb�w���#�Kn"�R�&���*��.�J3��7�z;��>���B��F�}J�t=N�v�Q�S�U��AY�u�\��j`���c��pg���j�Wn��q��u�4zx���{�V�o1��h҂��p��k��ӥ���<���ъ�@d���������������^&��߮���5������W@���Û�FF���Ǟ�nH��Hȡ�G�� Ƥ��C�������>��d����7��'���G0��O���o(������� ��7������ꖹ�U��>�������  �  �yN=(�M=��L=c9L=hxK=�J=��I=o2I=YoH=��G=L�F=8"F=p\E=ەD=y�C=6C==B=�rA=ҧ@=��?=S?=�?>=9p==I�<=�;=Z�:=D$:=�M9=�u8=��7=-�6=��5=�5=�"4=�?3=�Z2=[s1=މ0=�/=�.=P�-=$�,=R�+=��*=b�)=�(=��'=��&=�%=?�$= �#=��"=��!=�~ =�b=�B=�=��=�=E�=bg=O/=�=��=�m=�$=[�=��=t/=��=v=�
=F�=g?=<�=�Z=C�=�e=]��<���<��<ǔ�<�s�<�K�<�<���<��<d�<��<���<Dr�<��<Ƴ�<{L�<���<�n�<���<B~�<���<}�<���<	m�<�߯<�O�<���<'�<��<���<�X�<���<�<)z�<$؋<+5�<���<[�<őz<�Hs<��k<��d<7p]<l*V<v�N<ƤG<�e@<�)9<l�1<Ӽ*<��#<2a<�:<5<g�<J��;���;n��;���;,��;��;�!�;�k�;Uɐ;�;�;+�k;M�P;[.6;s�;��;1.�:ʘ�:8�P:���9��7�j��b?�����/���S�����}'�%�>���U��.l��E���Q���:��� ��룬�=$�������˻��ջ�߻_���M����&�����c����jb�����#�.n"�]�&���*�5�.�h3��7�i;���>���B��F�}J�d=N�f�Q�^�U��AY���\��j`���c��pg���j�Wn��q��u� zx���{�A�k1��s҂��p��v��å���<���ъ�Pd�����ꃏ�������v&��䮕��5������R@���Û�<F���Ǟ�pH��Dȡ�nG��Ƥ�
D�������>��W����7��%���I0��Z���l(��~���� ��/������򖹼[��7�������  �  )}N=�M=H�L=E>L=�}K=�J=��I=�9I=wH=�G=F�F=�+F=�fE=ʠD=!�C=�C=JB=��A=J�@=��?=X?=�P>=́==��<=P�;=�;=L9:=�c9=Y�8=��7=��6=��5=�5=u>4=k\3=\x2=*�1=ǩ0=�/=��.=u�-=W�,=��+=)+=�	*=�)=�(=?	'=�&=�$=��#=n�"=M�!=�� =)�=�t=�Q=�*=��=��=O�=�e=*=��=o�=�\=[=��=�g=�=�=wJ
=��=Jv=�=��=p=��=e =r%�<��<���<���<;��<gw�<{>�<���<��<�j�<��<(��<�^�<���<ŏ�<K �<��<3�<���<4�<r��<%�<=��<�<�t�<�ި<F�<��<��<�n�<�͖<�*�<��<�<!<�<h��<X�<ɍz<�>s<��k<��d<xT]<�V<��N<6wG<+2@<E�8<�1<w*<]A#<<��<��<��<�;���;���;c��;`��;y޸;=
�;-H�;ɚ�;��;��h;6$N;z3;{ ;/q�:�K�:��:��D:Ԛ�9���O�ӹ&�L�\����Ǻ����2��+�gHB�<6Y�T�o�n ���.�����>ࣻ̓������_ûؘͻ>�׻&��q�9��ީ���	�5��B���:����[���:#�Rs'�?�+���/���3���7��;���?�H�C��WG��K�|�N���R�93V��Y�we]���`��sd���g�Mak�Q�n�0r��u��x��2|�~|�,`��G��������5��=͇��b������Ȇ�����E����.��ܸ��dA��Oȕ�N��Ҙ��U���כ�Y��dٞ��X���ס�~U���Ҥ��O��̧�!H���ê�/?��X����5��l���q+�������!��+����������*��㍼�?���  �  0}N=�M=H�L=E>L=�}K=�J=��I=�9I=wH=�G=I�F=�+F=�fE=ɠD=�C=�C=JB=��A=H�@=��?=T?=�P>=Ձ==��<=J�;=�;=Q9:=�c9=_�8=��7=��6=��5={5=o>4=t\3=dx2=0�1=��0=�/=��.=u�-=]�,=��+=/+=�	*=�)=�(=A	'=�&=�$=��#=l�"=T�!=�� =-�=�t=�Q=�*=��=��=L�=�e=�)=��=s�=�\=Y=��=�g=�=�=xJ
=��=Mv=�=��=v=�=` =_%�<�<���<���<J��<�w�<�>�<���<��<�j�<��<��<�^�<���<���<V �<��<3�<���<4�<y��<%�<D��<�<�t�<�ި<&F�<	��<��<�n�<~͖<�*�<��<	�<<�<v��<Q�<��z<�>s<��k<��d<NT]<�V<;N<)wG<72@<d�8<�1<�w*<`A#<�<��<�<f�<t�;���;���;r��;n��;l޸;�	�;*H�;���;��;f�h;$N;�y3; ;Gr�:�J�:@��:x�D:��9lſ�J�ӹ �L��\����Ǻ������~+��GB��5Y���o�` ��p.�����ࣻm���c���_û٘ͻ��׻��q뻓�������	���B����":�ɞ�O���:#�5s'�I�+�¹/���3���7���;��?�N�C��WG��K�G�N�R�43V���Y�ke]��`��sd�z�g�2ak�c�n�+0r��u��x��2|�a|�`��;��������5��H͇��b������҆�����K����.��渒�dA��gȕ�N��yҘ��U���כ�Y��gٞ��X��}ס��U���Ҥ��O�� ̧�H���ê�*?��^���r5��t����+�������!��������Ŕ����ꍼ�:���  �  *}N=�M=E�L=J>L=�}K=�J=��I=�9I=%wH=�G=F�F=�+F=�fE=РD=�C=�C=JB=��A=D�@=��?=\?=�P>=؁==��<=O�;=�;=N9:=�c9=Y�8=~�7=��6=��5=|5=r>4=p\3=Xx2=/�1=��0=�/=��.=q�-=X�,=��+=*+=�	*=�)=�(=C	'=�&=�$=��#=i�"=U�!=�� =1�=�t=�Q=�*=��=��=F�=�e=�)=��=u�=�\=a=��=�g=�=�=tJ
=��=Pv=�=��=k=��=c =a%�<�<���<���<<��<ow�<>�<���<��<�j�<��<��<�^�<���<���<Z �<��< 3�<���<4�<y��<%�<B��<�<�t�<�ި<-F�<
��<��<�n�<|͖<�*�<��<�<<�<y��<T�<��z<�>s<��k<��d<QT]<�V<־N<wG<22@<I�8<�1<sw*<tA#<�<��<)�<k�<��;���;���;]��;i��;�޸;�	�;zH�;���;��;+�h;$N;`z3;4 ;�r�:�J�::?�D:���9���e�ӹy�L��\��W�Ǻ����f���+��HB��5Y���o�J ���.����8ࣻ��������_û��ͻ��׻���p�j�������	���'B����:����5��;#�,s'�_�+���/���3���7��;�$�?�/�C��WG��K�h�N�ۋR�B3V��Y�^e]�
�`��sd���g�Gak�W�n�'0r�،u�!�x��2|�{|�#`��B��������5��K͇��b�����������V����.���PA��bȕ�N��yҘ��U���כ�#Y��Tٞ��X��wס��U���Ҥ��O��"̧� H���ê�/?��c���n5��p����+�������!�� ����������������<���  �  0}N=�M=J�L=B>L=�}K=�J=��I=�9I=wH=�G=J�F=�+F=�fE=͠D=�C=�C=JB=��A=J�@=��?=S?=�P>=ρ==��<=M�;=�;=Q9:=�c9=`�8=��7=��6=��5=|5=r>4=n\3=ax2=,�1=ũ0=�/=��.=w�-=]�,=��+=,+=�	*=�)=�(=@	'=�&=�$=��#=i�"=W�!=�� =.�=�t=�Q=�*=��=��=H�=�e=�)=��=o�=�\=Z=��=�g=�=�=zJ
=��=Fv=�=��=s=��=a =b%�<��<���<���<G��<rw�<�>�<���<��<�j�<��<!��<�^�<���<���<\ �<��<3�<���<4�<u��<"%�<I��<�<�t�<�ި<F�<��<��<}n�<�͖<�*�<��<
�<!<�<e��<K�<��z<�>s<��k<��d<cT]<�V<��N<7wG<92@<d�8<��1<�w*<PA#<�<��<�<p�<~�;���;��;���;d��;�޸;�	�;ZH�;���;��;��h;($N;�y3;I ;�q�:�K�:���:)�D:h��9�뿷�ӹ��L��[����Ǻ����a���+�HB�6Y�t�o�� ���.�����ࣻ����x���_û�ͻk�׻%��q뻄������	���B����:�Þ�D���:#�(s'�W�+���/���3���7��;��?�L�C��WG��K�]�N�ȋR�+3V�
�Y��e]���`��sd���g�Aak�]�n�$0r��u�
�x��2|�d|�`��<��������5��?͇��b������Ն�����L����.��丒�ZA��aȕ�N��|Ҙ��U���כ�"Y��eٞ��X���ס�U���Ҥ��O��̧�H���ê�*?��X����5��z���z+�������!��*������Ɣ��-��㍼�9���  �  2}N=�M=J�L=A>L=�}K=�J=��I=�9I=wH=
�G=F�F=�+F=�fE=ΠD=�C=�C=JB=��A=G�@=��?=S?=�P>=с==��<=H�;=�;=Q9:=�c9=_�8=s�7=��6=��5=�5=m>4=j\3=bx2=$�1=ǩ0=�/=��.=p�-=U�,=��+='+=�	*=�)=�(=?	'=�&=�$=��#=p�"=P�!=�� =0�=�t=�Q=�*=��=��=N�=�e=�)=��=n�=�\=T=��=�g=�=�=qJ
=��=Ev=�=��=r=��=[ =k%�<��<���<���<@��<qw�<>�<���<���<�j�<��<7��<�^�<��<���<R �<��<3�<���<4�<|��<"%�<?��<)�<�t�<�ި<(F�<��<��<yn�<�͖<�*�<��<��<<�<q��<O�<��z<�>s<��k<t�d<YT]<�V<��N<1wG<2@<g�8<�1<�w*<NA#<�<��<�<��<v�;��;���;|��;��;�޸;
�;SH�;ٚ�;��;b�h;�$N;�y3;� ;�q�:�K�:&��:�D:Z��9����E�ӹ!�L��[��y�ǺJ������+�HB��6Y�T�o�� ��m.����Mࣻ��������_û��ͻ[�׻)���p�Y��ة���	�*��B����:����B���:#�Bs'�>�+���/���3���7��;���?�`�C��WG��K�X�N��R�N3V���Y��e]���`�td���g�Kak�r�n�0r��u��x��2|�r|� `��A��������5��:͇��b������҆�����J����.��۸��]A��Yȕ�N��uҘ��U���כ�Y��fٞ��X��{ס�U���Ҥ��O��̧�#H���ê�@?��^���v5��v���{+�������!��5����������"��捼�R���  �  0}N=�M=G�L=I>L=�}K=�J=��I=�9I=wH=	�G=H�F=�+F=�fE=РD=�C=�C=JB=��A=H�@=��?=V?=�P>=Ӂ==��<=O�;=�;=M9:=�c9=_�8=|�7=��6=��5={5=p>4=n\3=Wx2=,�1=é0=�/=��.=q�-=Z�,=��+=&+=�	*=�)=�(=>	'=�&=�$=��#=m�"=W�!=�� =2�=�t=�Q=�*=��=��=K�=�e=�)=��=n�=�\=\=��=�g=�=�=tJ
=��=Cv=�=��=k=��=` =^%�<��<���<���<A��<lw�<x>�<���<��<�j�<��<#��<�^�<��<���<g �<��<3�<���<4�<{��<*%�<F��<$�<�t�<�ި<)F�<��<��<�n�<͖<�*�<��<�<<�<l��<C�<��z<�>s<��k<��d<YT]<�V<��N< wG<*2@<b�8<�1<{w*<mA#<�<��<�<j�<��;
��;���;���;r��;�޸;
�;rH�;���;�;r�h;�$N;z3;W ;r�:hK�:��:a�D:蛽9���%�ӹ��L��\��x�Ǻ���n���+��HB�6Y���o�� ���.����(ࣻ��������_û��ͻ`�׻*���p뻁�������	���B����:����1���:#� s'�I�+���/���3���7��;�
�?�A�C��WG��K�^�N�֋R�?3V��Y��e]��`��sd���g�Fak�^�n�*0r��u��x��2|�n|�$`��G��������5��A͇��b������φ�����K����.��⸒�TA��\ȕ�	N��wҘ��U���כ�Y��bٞ��X��{ס��U���Ҥ��O��̧�%H���ê�0?��c���{5������}+�������!��'������̔��$���@���  �  '}N=�M=H�L=C>L=�}K=�J=��I=�9I=%wH=�G=K�F=�+F=�fE=נD=�C=�C=JB=��A=I�@=��?=\?=�P>=؁==��<=L�;=�;=P9:=�c9=V�8=��7=��6=��5=w5=m>4=m\3=Ux2=.�1=��0=�/=��.=r�-=Y�,=��+=.+=�	*=�)=�(=C	'=�&=�$= �#=j�"=[�!=�� =4�=�t=�Q=�*=��=��=H�=�e=�)=��=t�=�\=Y=��=�g=�=�=uJ
=��=Gv=�=��=h=��=] =S%�<��<���<���<4��<qw�<�>�<���<��<�j�<��<"��<�^�<��<���<f �<	��<*3�<���<4�<{��<&%�<L��<�<�t�<�ި<-F�<��<��<�n�<|͖<�*�<��<
�<<�<i��<I�<��z<�>s<��k<��d<?T]<�V<��N<wG<92@<;�8< �1<}w*<WA#<�<��<(�<i�<��;���;��;���;m��;�޸;�	�;�H�;���;�;��h;�$N;lz3;Q ;�r�:9K�:ď�:�D:���9ῷ6�ӹ��L�]��+�Ǻb�������+��HB��5Y��o�x ���.����(ࣻ����b���_ûӘͻ{�׻���p�y�������	����B����:���� ���:#�s'�U�+���/���3���7��;��?�L�C�XG��K�f�N�ߋR�93V�!�Y�ze]�&�`��sd���g�Oak�g�n�>0r��u�1�x��2|��|�`��?��������5��G͇��b������ņ�����L����.��긒�EA��bȕ��M��wҘ��U���כ�Y��Sٞ��X��wס�yU���Ҥ��O��#̧�H���ê�)?��g���~5��{����+�������!��$������ɔ��'��􍼼8���  �  '}N=�M=F�L=F>L=�}K=�J=��I=�9I=!wH=
�G=K�F=�+F=�fE=נD=�C=�C=JB=��A=K�@=��?=Y?=�P>=Ё==��<=Q�;=�;=M9:=�c9=V�8=y�7=��6=��5=y5=l>4=h\3=Wx2='�1=��0=�/=��.=p�-=U�,=��+='+=�	*=�)=�(=>	'=�&=�$=��#=o�"=V�!=�� =5�=�t=�Q=�*=��=��=M�=�e=�)=��=m�=�\=[=��=�g=�=�=rJ
=��=Ev=�=��=g=��=[ =V%�<��<���<���<1��<ow�<w>�<���<��<�j�<��<+��<�^�<��<���<\ �<��<%3�<���<4�<���<+%�<J��<%�<�t�<�ި<!F�<��<��<�n�<}͖<�*�<��<��<<�<e��<L�<��z<�>s<��k<t�d<CT]<�V<��N<wG<2@<=�8<�1<vw*<bA#<
<��<�<��<��;��;��;���;���;�޸;�	�;�H�;�;��;��h;�$N;Ez3;� ;�q�:�K�:i��:�D:�9鿷W�ӹd�L��\����Ǻ������!+��HB�_6Y���o�w ���.����Hࣻ��������_û��ͻT�׻*���p�N�������	����A�����9����"���:#�)s'�B�+���/���3���7��;��?�B�C��WG��K�e�N��R�C3V��Y��e]��`��sd���g�`ak�n�n�50r��u�$�x��2|��|� `��G��������5��?͇��b������ǆ�����H����.��ظ��JA��^ȕ��M��oҘ��U���כ�Y��[ٞ��X���ס�~U���Ҥ��O��!̧� H���ê�5?��e����5��x����+�������!��4������Ŕ��,������E���  �  3}N=�M=G�L=A>L=�}K=�J=��I=�9I=wH=�G=L�F=�+F=�fE=РD=&�C=�C=JB=��A=N�@=��?=R?=�P>=ҁ==��<=H�;=�;=M9:=�c9=_�8=w�7=��6=��5=v5=m>4=h\3=Xx2="�1=��0=�/=��.=o�-=U�,=��+=&+=�	*=�)=�(=A	'=�&=�$=��#=u�"=V�!=�� =0�=�t=�Q=�*=��=��=S�=�e=�)=��=o�=�\=S=��=�g=�=�=pJ
=��=;v=�=��=h=��=Z =S%�<��<���<���<=��<qw�<w>�<���<���<�j�<��</��<�^�<��<ɏ�<f �<"��<3�<Ƶ�<4�<}��<7%�<K��<3�<�t�<�ި<&F�<��<��<yn�<�͖<�*�<��<��<<�<c��<8�<��z<|>s<��k<k�d<NT]<�V<��N< wG<2@<k�8<�1<zw*<LA#<�<��<�<��<T�;>��;��;н�;���;�޸;q
�;hH�;��;"�;��h;�$N;�y3;� ;r�:L�:D��:�D:O��9�濷ɺӹ��L�(\���Ǻ~������+��HB��6Y���o�� ���.�� ��Jࣻb�������_û��ͻc�׻���p�[������	����A�����9����:���:#�#s'�(�+���/���3���7���;��?�a�C��WG��K�J�N��R�M3V��Y��e]��`�td���g�[ak�r�n�:0r�"�u��x��2|�r|�`��F��������5��9͇��b������ц�����@����.��и��ZA��Eȕ�N��tҘ��U���כ�Y��oٞ��X��~ס�wU���Ҥ��O��̧�"H���ê�:?��c����5�������+�������!��8������Ք��0��퍼�J���  �  (}N=�M=H�L=E>L=�}K=�J=��I=�9I=$wH=�G=G�F=�+F=�fE=ՠD=#�C=�C=JB=��A=H�@=��?=\?=�P>=ց==��<=J�;=�;=M9:=�c9=W�8=w�7=��6=��5=v5=i>4=e\3=Tx2=#�1=��0=�/=��.=j�-=S�,=��+=&+=�	*=�)=�(=D	'=�&=�$= �#=s�"=U�!=�� =6�=�t=�Q=�*=��=��=N�=�e=*=��=r�=�\=Y=��=�g=�=�=jJ
=��=Av=�=��=d=�=W =R%�<��<���<���<1��<`w�<x>�<���<��<�j�<��<-��<�^�<��<���<d �<��<$3�<õ�<4�<���<.%�<B��<3�<�t�<�ި<,F�<��<��<�n�<�͖<�*�<��<��<	<�<j��<?�<��z<~>s<��k<i�d<@T]<�V<��N<wG<2@<A�8<ڱ1<{w*<\A#<�<��<#�<��<��;B��;���;���;���;�޸;[
�;�H�;��;�;��h;�$N;z3;� ;�r�:�K�:���:��D:d��9��2�ӹ��L�5]��Q�Ǻf���Ο�L+��HB��6Y���o�� ���.��G��Zࣻ��������_ûȘͻ\�׻����p�4�������	����A�����9���� ���:#�"s'�:�+���/���3���7��;��?�I�C��WG��K�w�N��R�`3V�!�Y��e]��`�td���g�iak�z�n�;0r��u�3�x��2|��|�.`��E��������5��;͇��b�������������J����.��Ը��JA��Iȕ� N��kҘ��U���כ�Y��Sٞ��X��xס�xU���Ҥ��O��̧�(H���ê�:?��o���}5�������+�������!��9������є��'������H���  �  '}N=�M=C�L=D>L=�}K=�J=��I=�9I=#wH=	�G=S�F=�+F=�fE=٠D=�C=�C=JB=��A=Q�@=��?=Y?=�P>=Ӂ==��<=V�;=�;=M9:=�c9=X�8=�7=��6=��5=o5=k>4=g\3=Ux2=)�1=��0=
�/=��.=m�-=[�,=��+=-+=�	*=�)=�(=A	'=�&=�$=��#=n�"=b�!=�� =7�=�t=�Q=�*=��=��=L�=�e=�)=��=p�=�\=^=��=�g=�=�=oJ
=��=@v=�=��=f=�=Y =A%�<��<���<���<5��<kw�<{>�<���<��<�j�<��<"��<�^�<��<ɏ�<r �<��<-3�<���<#4�<���</%�<\��<"�<�t�<�ި<'F�<��<��<�n�<v͖<�*�< ��<
�<<�<_��<:�<��z<�>s<��k<w�d<>T]<zV<��N<�vG<92@<<�8<�1<kw*<\A#<<��<�<w�<��;��;W��;ƽ�;���;�޸;	
�;�H�;ך�;D�;�h;�$N;Kz3;~ ;Rr�:|K�:��:9�D:���9�ۿ��ӹ��L�W]����ǺR������-+��HB�86Y�>�o�� ���.��2��ࣻÃ��e���_û��ͻ^�׻���p�]�������	�ޭ��A�����9�������:#��r'�B�+���/���3���7���;�
�?�1�C�XG��K�u�N�ԋR�L3V�*�Y��e]�5�`��sd���g�bak�r�n�]0r��u�8�x��2|��|�#`��A���Û���5��C͇��b������Ɇ�����@����.��ݸ��BA��\ȕ��M��nҘ��U���כ�Y��Xٞ��X��}ס�U���Ҥ��O��)̧�H���ê�)?��r����5�������+�������!��2������ٔ��/������8���  �  &}N=�M=D�L=@>L=�}K=�J=��I=�9I=$wH=�G=Q�F=�+F=�fE=ݠD=%�C=�C=JB=��A=P�@=��?=\?=�P>=ف==��<=M�;=�;=M9:=�c9=V�8=v�7=��6=��5=t5=k>4=b\3=Rx2=�1=��0=�/=��.=h�-=T�,=��+=,+=�	*=�)=�(=E	'=�&=�$=��#=r�"=^�!=�� =5�=u=�Q=�*=��=��=P�=�e=*=��=t�=�\=W=��=�g=�=�=hJ
=��==v=�=��=b=�=V =M%�<��<���<���<,��<dw�<x>�<���<��<�j�<��<1��<�^�<��<ˏ�<m �<��<.3�<ȵ�<*4�<~��<-%�<W��<)�<�t�<�ި<5F�<��<��<{n�<y͖<�*�<���<��<<�<f��<;�<��z<g>s<��k<V�d<DT]<�V<��N<wG<2@<6�8<��1<nw*<GA#<�<��<1�<��<��;"��;A��;���;���;߸;p
�;�H�;Қ�;7�;
�h;�$N;}z3;� ;"s�:�K�:��:	�D:R��9����ӹ��L��\����Ǻ�������x+��HB��6Y���o�� ���.��U��RࣻɃ��t���_û֘ͻi�׻�Ữp�*�������	����A�����9�������:#�s'�3�+���/���3�}�7��;��?�N�C�
XG��K�y�N��R�g3V��Y��e]��`�td���g�qak�~�n�C0r��u�)�x��2|��|�(`��D���Û���5��B͇��b�������������>����.��߸��AA��Cȕ��M��sҘ��U���כ�Y��Uٞ��X��oס�yU���Ҥ��O��&̧�H���ê�9?��s����5�������+�������!��B������֔��*������J���  �  ,}N=�M=J�L=G>L=�}K=�J=��I=�9I="wH=�G=I�F=�+F=�fE=ԠD=�C=�C=JB=��A=I�@=��?=X?=�P>=Ӂ==��<=M�;=�;=M9:=�c9=_�8=w�7=��6=��5=u5=g>4=e\3=]x2=�1=��0=�/=��.=l�-=Z�,=��+=$+=�	*=�)=�(=>	'=�&=�$=��#=r�"=X�!=�� =8�=�t=�Q=�*=��=��=N�=�e=�)=��=m�=�\=Y=��=�g=�=�=mJ
=��=7v=�=��=j=�=R =Q%�<��<���<���<C��<bw�<v>�<���<��<�j�<��<��<�^�<��<�<l �<"��< 3�<���<4�<���<=%�<I��</�<�t�<�ި<!F�<
��<��<�n�<�͖<�*�<	��< �<<�<g��<4�<��z<i>s<��k<Z�d<@T]<wV<��N<wG<2@<P�8<ձ1<�w*<fA#<�<��<�<v�<��;A��;��;��;���;�޸;(
�;�H�; ��;I�;��h;�$N;Dz3;h ;Tr�:�K�:���:3�D:y��92��O�ӹ��L��\��9�Ǻ������@+�EHB��6Y���o�� ��}.��9��ࣻ��������_û��ͻV�׻&��q�j�������	����A�����9�������:#�s'�:�+���/���3���7��;��?�E�C��WG��K�h�N�ʋR�V3V��Y��e]��`�"td���g�aak���n�<0r�)�u�'�x��2|�e|�+`��F��������5��=͇��b������ˆ�����G����.��ϸ��NA��Rȕ�N��dҘ��U���כ�
Y��Wٞ��X���ס��U���Ҥ��O��̧�.H���ê�3?��m����5�������+�������!��A������ڔ��-������E���  �  &}N=�M=D�L=@>L=�}K=�J=��I=�9I=$wH=�G=Q�F=�+F=�fE=ݠD=%�C=�C=JB=��A=P�@=��?=\?=�P>=ف==��<=M�;=�;=M9:=�c9=V�8=v�7=��6=��5=t5=k>4=b\3=Rx2=�1=��0=�/=��.=h�-=T�,=��+=,+=�	*=�)=�(=E	'=�&=�$=��#=r�"=^�!=�� =5�=u=�Q=�*=��=��=P�=�e=*=��=t�=�\=W=��=�g=�=�=hJ
=��==v=�=��=b=�=V =M%�<��<���<���<,��<dw�<x>�<���<��<�j�<��<1��<�^�<��<ˏ�<m �<��<.3�<ȵ�<*4�<~��<-%�<W��<(�<�t�<�ި<5F�<��<��<{n�<y͖<�*�<���<��<<�<f��<;�<��z<g>s<��k<V�d<DT]<�V<��N<wG<2@<6�8<��1<nw*<GA#<�<��<1�<��<��;"��;A��;���;���;߸;p
�;�H�;Қ�;7�;	�h;�$N;}z3;� ;!s�:�K�:��:�D:K��9P��ӹ��L��\����Ǻ�������x+��HB��6Y���o�� ���.��U��RࣻɃ��t���_ûטͻi�׻�ữp�+�������	����A�����9�������:#�s'�3�+���/���3�~�7��;��?�N�C�
XG��K�y�N��R�g3V��Y��e]��`�td���g�qak�}�n�C0r��u�)�x��2|��|�(`��D���Û���5��B͇��b�������������>����.��߸��AA��Cȕ��M��sҘ��U���כ�Y��Uٞ��X��oס�yU���Ҥ��O��&̧�H���ê�9?��s����5�������+�������!��B������֔��*������J���  �  '}N=�M=C�L=D>L=�}K=�J=��I=�9I=#wH=	�G=S�F=�+F=�fE=٠D=�C=�C=JB=��A=Q�@=��?=Y?=�P>=Ӂ==��<=V�;=�;=M9:=�c9=X�8=�7=��6=��5=o5=k>4=g\3=Ux2=)�1=��0=
�/=��.=m�-=[�,=��+=-+=�	*=�)=�(=A	'=�&=�$=��#=n�"=b�!=�� =7�=�t=�Q=�*=��=��=L�=�e=�)=��=p�=�\=^=��=�g=�=�=oJ
=��=@v=�=��=f=�=Y =A%�<��<���<���<5��<kw�<|>�<���<��<�j�<��<"��<�^�<��<ɏ�<r �<��<-3�<���<#4�<���</%�<\��<"�<�t�<�ި<'F�<��<��<�n�<u͖<�*�< ��<
�<<�<_��<:�<��z<�>s<��k<w�d<>T]<zV<��N<�vG<92@<=�8<�1<kw*<\A#<<��<�<w�<��;��;X��;ƽ�;���;�޸;	
�;�H�;ך�;D�;�h;�$N;Jz3;} ;Or�:zK�:
��:3�D:~��9�ܿ��ӹ��L�[]����ǺU������.+��HB�96Y�?�o�� ���.��2��ࣻă��e���_û��ͻ^�׻���p�]�������	�ޭ��A�����9�������:#��r'�B�+���/���3���7���;�
�?�1�C�XG��K�u�N�ԋR�L3V�*�Y��e]�6�`��sd���g�bak�r�n�]0r��u�8�x��2|��|�#`��A���Û���5��C͇��b������Ɇ�����@����.��ݸ��BA��\ȕ��M��nҘ��U���כ�Y��Xٞ��X��}ס�U���Ҥ��O��)̧�H���ê�)?��r����5�������+�������!��2������ٔ��/������8���  �  (}N=�M=H�L=E>L=�}K=�J=��I=�9I=$wH=�G=G�F=�+F=�fE=ՠD=#�C=�C=JB=��A=H�@=��?=\?=�P>=ց==��<=J�;=�;=M9:=�c9=W�8=w�7=��6=��5=v5=i>4=e\3=Tx2=#�1=��0=�/=��.=j�-=S�,=��+=&+=�	*=�)=�(=D	'=�&=�$= �#=s�"=U�!=�� =6�=�t=�Q=�*=��=��=N�=�e=*=��=s�=�\=Y=��=�g=�=�=kJ
=��=Av=�=��=e=�=X =R%�<��<���<���<1��<`w�<x>�<���<��<�j�<��<-��<�^�<��<���<d �<��<$3�<õ�<4�<���<.%�<B��<3�<�t�<�ި<,F�<��<��<�n�<�͖<�*�<��<��<	<�<j��<?�<��z<~>s<��k<i�d<@T]<�V<��N<wG<2@<A�8<۱1<{w*<\A#<�<��<$�<��<��;C��;���;���;���;�޸;[
�;�H�;��;�;��h;�$N;~z3;� ;�r�:�K�:���:��D:R��96��D�ӹ��L�9]��U�Ǻj���П�N+��HB��6Y���o�� ���.��G��[ࣻ��������_ûɘͻ\�׻����p�4�������	����A�����9���� ���:#�"s'�:�+���/���3���7��;��?�I�C��WG��K�w�N��R�`3V�!�Y��e]��`�td���g�iak�z�n�;0r��u�3�x��2|��|�.`��E��������5��;͇��b�������������J����.��Ը��JA��Iȕ� N��kҘ��U���כ�Y��Sٞ��X��xס�xU���Ҥ��O��̧�(H���ê�:?��o���}5�������+�������!��9������є��'������H���  �  3}N=�M=G�L=A>L=�}K=�J=��I=�9I=wH=�G=L�F=�+F=�fE=РD=&�C=�C=JB=��A=N�@=��?=R?=�P>=ҁ==��<=H�;=�;=M9:=�c9=_�8=w�7=��6=��5=v5=m>4=h\3=Xx2="�1=��0=�/=��.=o�-=U�,=��+=&+=�	*=�)=�(=A	'=�&=�$=��#=u�"=V�!=�� =0�=�t=�Q=�*=��=��=S�=�e=�)=��=o�=�\=S=��=�g=�=�=pJ
=��=<v=�=��=h=��=Z =T%�<��<���<���<=��<qw�<x>�<���<���<�j�<��<0��<�^�<��<ɏ�<f �<"��<3�<Ƶ�<4�<}��<6%�<K��<3�<�t�<�ި<&F�<��<��<yn�<�͖<�*�<��<��<<�<b��<8�<��z<|>s<��k<k�d<NT]<�V<��N<!wG<2@<k�8<�1<zw*<MA#<�<��<�<��<T�;>��;��;ѽ�;���;�޸;q
�;hH�;��;!�;��h;�$N;�y3;� ;r�:�K�:?��:؅D::��9�翷ߺӹ��L�-\��"�Ǻ�������+��HB��6Y���o�� ���.��!��Jࣻc�������_û��ͻc�׻���p�[������	����A�����9����:���:#�#s'�(�+���/���3���7���;��?�a�C��WG��K�J�N��R�M3V��Y��e]��`�td���g�[ak�r�n�:0r�"�u��x��2|�r|�`��F��������5��9͇��b������ц�����@����.��и��ZA��Eȕ�N��tҘ��U���כ�Y��oٞ��X��~ס�wU���Ҥ��O��̧�"H���ê�:?��c����5�������+�������!��8������Ք��0��퍼�J���  �  '}N=�M=F�L=F>L=�}K=�J=��I=�9I=!wH=
�G=K�F=�+F=�fE=נD=�C=�C=JB=��A=K�@=��?=Y?=�P>=Ё==��<=Q�;=�;=M9:=�c9=V�8=y�7=��6=��5=y5=l>4=h\3=Wx2='�1=��0=�/=��.=p�-=U�,=��+='+=�	*=�)=�(=>	'=�&=�$=��#=o�"=V�!=�� =5�=�t=�Q=�*=��=��=M�=�e=�)=��=m�=�\=[=��=�g=�=�=sJ
=��=Ev=�=��=g=��=[ =W%�<��<���<���<2��<ow�<w>�<���<��<�j�<��<+��<�^�<��<���<\ �<��<%3�<���<4�<���<+%�<J��<%�<�t�<�ި<!F�<��<��<�n�<}͖<�*�<��<��<<�<e��<L�<��z<�>s<��k<t�d<CT]<�V<��N<wG<2@<=�8<�1<vw*<cA#<
<��<�<��<��;��;��;���;���;�޸;�	�;�H�;�;��;��h;�$N;Cz3;� ;�q�:�K�:d��:��D:ٛ�9�꿷p�ӹp�L��\����Ǻ"������$+��HB�a6Y���o�x ���.����Iࣻ��������_û��ͻT�׻*���p�O�������	����A�����9����"���:#�)s'�B�+���/���3���7��;��?�B�C��WG��K�e�N��R�C3V��Y��e]��`��sd���g�`ak�n�n�50r��u�$�x��2|��|� `��G��������5��?͇��b������ǆ�����H����.��ظ��JA��^ȕ��M��oҘ��U���כ�Y��[ٞ��X���ס�~U���Ҥ��O��!̧� H���ê�5?��e����5��x����+�������!��4������Ŕ��,������E���  �  '}N=�M=H�L=C>L=�}K=�J=��I=�9I=%wH=�G=K�F=�+F=�fE=נD=�C=�C=JB=��A=I�@=��?=\?=�P>=؁==��<=L�;=�;=P9:=�c9=V�8=��7=��6=��5=w5=m>4=m\3=Ux2=.�1=��0=�/=��.=r�-=Y�,=��+=.+=�	*=�)=�(=C	'=�&=�$= �#=j�"=[�!=�� =4�=�t=�Q=�*=��=��=H�=�e=�)=��=t�=�\=Y=��=�g=�=�=uJ
=��=Hv=�=��=h=��=] =S%�<��<���<���<4��<qw�<�>�<���<��<�j�<��<"��<�^�<��<���<f �<	��<*3�<���<4�<{��<&%�<L��<�<�t�<�ި<-F�<��<��<�n�<{͖<�*�<��<
�<<�<h��<I�<��z<�>s<��k<��d<?T]<�V<��N<wG<92@<;�8<�1<~w*<WA#<�<��<)�<i�<��;���;��;���;m��;�޸;�	�;�H�;���;�;��h;�$N;iz3;O ;�r�:4K�:���:�D:g��9�⿷O�ӹ��L�]��1�Ǻh�������+��HB��5Y��o�y ���.����)ࣻ����b���_ûԘͻ|�׻���p�y�������	����B����:���� ���:#�s'�U�+���/���3���7��;��?�L�C�XG��K�f�N�ߋR�93V�!�Y�ze]�&�`��sd���g�Oak�g�n�>0r��u�1�x��2|��|�`��?��������5��G͇��b������ņ�����L����.��긒�EA��bȕ��M��wҘ��U���כ�Y��Sٞ��X��wס�yU���Ҥ��O��#̧�H���ê�)?��g���~5��{����+�������!��$������ɔ��'��􍼼8���  �  0}N=�M=G�L=I>L=�}K=�J=��I=�9I=wH=	�G=H�F=�+F=�fE=РD=�C=�C=JB=��A=H�@=��?=V?=�P>=Ӂ==��<=O�;=�;=M9:=�c9=_�8=|�7=��6=��5={5=p>4=n\3=Wx2=,�1=é0=�/=��.=q�-=Z�,=��+=&+=�	*=�)=�(=>	'=�&=�$=��#=m�"=W�!=�� =2�=�t=�Q=�*=��=��=K�=�e=�)=��=n�=�\=\=��=�g=�=�=tJ
=��=Cv=�=��=k=��=` =^%�<��<���<���<B��<lw�<y>�<���<��<�j�<��<#��<�^�<��<���<g �<��<3�<���<4�<{��<*%�<E��<$�<�t�<�ި<)F�<��<��<�n�<͖<�*�<��<�<<�<l��<C�<��z<�>s<��k<��d<YT]<�V<��N< wG<*2@<b�8<�1<|w*<mA#<�<��<�<j�<��;��;���;���;r��;�޸;
�;rH�;���;�;q�h;�$N;z3;U ;r�:bK�:
��:U�D:ћ�9u��>�ӹ��L��\��~�Ǻ	���q���+��HB�6Y���o�� ���.����)ࣻ��������_û��ͻ`�׻+���p뻁�������	���B����:����1���:#� s'�I�+���/���3���7��;�
�?�A�C��WG��K�^�N�֋R�?3V��Y��e]��`��sd���g�Fak�^�n�*0r��u��x��2|�n|�$`��G��������5��A͇��b������φ�����K����.��⸒�TA��\ȕ�	N��wҘ��U���כ�Y��cٞ��X��{ס��U���Ҥ��O��̧�%H���ê�0?��c���{5������}+�������!��'������̔��$���@���  �  2}N=�M=J�L=A>L=�}K=�J=��I=�9I=wH=
�G=F�F=�+F=�fE=ΠD=�C=�C=JB=��A=G�@=��?=S?=�P>=с==��<=H�;=�;=Q9:=�c9=_�8=s�7=��6=��5=�5=m>4=j\3=bx2=$�1=ǩ0=�/=��.=p�-=U�,=��+='+=�	*=�)=�(=?	'=�&=�$=��#=p�"=P�!=�� =0�=�t=�Q=�*=��=��=N�=�e=�)=��=o�=�\=T=��=�g=�=�=qJ
=��=Ev=�=��=s=��=\ =k%�<��<���<���<@��<qw�<�>�<���< ��<�j�<��<7��<�^�<��<���<R �<��<3�<���<4�<|��<"%�<?��<)�<�t�<�ި<(F�<��<��<yn�<�͖<�*�<��<��<<�<q��<O�<��z<�>s<��k<t�d<ZT]<�V<��N<1wG<2@<h�8<�1<�w*<NA#<�<��<�<��<w�;��;���;}��;��;�޸;
�;SH�;ٚ�;��;`�h;�$N;�y3;� ;�q�:�K�:!��:��D:D��9Y���[�ӹ,�L��[��~�ǺP������+�HB��6Y�V�o�� ��n.����Nࣻ��������_û��ͻ[�׻*���p�Z��ة���	�*��B����:����B���:#�Bs'�>�+���/���3���7��;���?�`�C��WG��K�X�N��R�N3V���Y��e]���`�td���g�Kak�r�n�0r��u��x��2|�r|� `��A��������5��:͇��b������҆�����J����.��۸��]A��Yȕ�N��uҘ��U���כ�Y��fٞ��X��{ס�U���Ҥ��O��̧�#H���ê�@?��^���v5��v���{+�������!��5����������"��捼�R���  �  0}N=�M=J�L=B>L=�}K=�J=��I=�9I=wH=�G=J�F=�+F=�fE=͠D=�C=�C=JB=��A=J�@=��?=S?=�P>=ρ==��<=M�;=�;=Q9:=�c9=`�8=��7=��6=��5=|5=r>4=n\3=ax2=,�1=ũ0=�/=��.=w�-=]�,=��+=,+=�	*=�)=�(=@	'=�&=�$=��#=i�"=W�!=�� =.�=�t=�Q=�*=��=��=H�=�e=�)=��=o�=�\=Z=��=�g=�=�=zJ
=��=Fv=�=��=s=��=a =b%�<��<���<���<H��<sw�<�>�<���<��<�j�<��<!��<�^�<���<���<\ �<��<3�<���<4�<u��<"%�<I��<�<�t�<�ި<F�<��<��<}n�<�͖<�*�<��<
�<!<�<e��<K�<��z<�>s<��k<��d<cT]<�V<��N<7wG<92@<d�8<��1<�w*<QA#<�<��<�<p�<�;���;��;���;d��;�޸;�	�;ZH�;���;��;��h;'$N;�y3;G ;�q�:�K�:���: �D:W��9��ӹ��L��[�� �Ǻ����c���+�HB�!6Y�u�o�� ���.�����ࣻ����y���_û�ͻk�׻%��q뻅������	���B����:�Þ�D���:#�(s'�W�+���/���3���7��;��?�L�C��WG��K�]�N�ȋR�+3V�
�Y��e]���`��sd���g�Aak�]�n�$0r��u�
�x��2|�d|�`��<��������5��?͇��b������Ն�����L����.��丒�ZA��aȕ�N��|Ҙ��U���כ�"Y��eٞ��X���ס�U���Ҥ��O��̧�H���ê�*?��X����5��z���z+�������!��*������Ɣ��-��㍼�9���  �  *}N=�M=E�L=J>L=�}K=�J=��I=�9I=%wH=�G=F�F=�+F=�fE=РD=�C=�C=JB=��A=D�@=��?=\?=�P>=ف==��<=O�;=�;=N9:=�c9=Y�8=~�7=��6=��5=|5=r>4=p\3=Xx2=/�1=��0=�/=��.=q�-=X�,=��+=*+=�	*=�)=�(=C	'=�&=�$=��#=i�"=U�!=�� =1�=�t=�Q=�*=��=��=F�=�e=�)=��=u�=�\=a=��=�g=�=�=tJ
=��=Pv=�=��=k=��=c =b%�<�<���<���<=��<ow�<>�<���<��<�j�<��<��<�^�<���<���<Z �<��< 3�<���<4�<y��<%�<B��<�<�t�<�ި<-F�<	��<��<�n�<|͖<�*�<��<�<<�<y��<T�<��z<�>s<��k<��d<QT]<�V<׾N<wG<32@<I�8<�1<tw*<tA#<�<��<*�<k�<��;���;���;]��;i��;�޸;�	�;zH�;���;��;*�h;$N;^z3;3 ;�r�:�J�:돕:9�D:���9����q�ӹ�L��\��Z�Ǻ����h���+��HB��5Y���o�J ���.����9ࣻ��������_û��ͻ��׻���p�j�������	���'B����:����5��;#�,s'�_�+���/���3���7��;�$�?�/�C��WG��K�h�N�ۋR�B3V��Y�^e]�
�`��sd���g�Gak�W�n�'0r�،u�!�x��2|�{|�#`��B��������5��K͇��b�����������V����.���PA��bȕ�N��yҘ��U���כ�#Y��Tٞ��X��wס��U���Ҥ��O��"̧� H���ê�/?��c���n5��p����+�������!�� ����������������<���  �  0}N=�M=H�L=E>L=�}K=�J=��I=�9I=wH=�G=I�F=�+F=�fE=ɠD=�C=�C=JB=��A=H�@=��?=T?=�P>=Ձ==��<=J�;=�;=Q9:=�c9=_�8=��7=��6=��5={5=o>4=t\3=dx2=0�1=��0=�/=��.=u�-=]�,=��+=/+=�	*=�)=�(=A	'=�&=�$=��#=m�"=T�!=�� =-�=�t=�Q=�*=��=��=L�=�e=�)=��=s�=�\=Y=��=�g=�=�=xJ
=��=Mv=�=��=v=�=` =`%�<�<���<���<J��<�w�<�>�<���<��<�j�<��<��<�^�<���<���<V �<��<3�<���<4�<y��<%�<D��<�<�t�<�ި<&F�<	��<��<�n�<~͖<�*�<��<	�<<�<v��<Q�<��z<�>s<��k<��d<NT]<�V<;N<)wG<72@<d�8<�1<�w*<`A#<�<��<�<g�<t�;���;���;r��;n��;k޸;�	�;*H�;���;��;f�h;$N;�y3; ;Er�:�J�:?��:u�D:��9�ſ�P�ӹ#�L��\����Ǻ������+��GB��5Y���o�` ��p.�����ࣻm���c���_ûژͻ��׻��q뻔�������	���B����":�ɞ�O���:#�5s'�I�+�¹/���3���7���;��?�N�C��WG��K�G�N�R�43V���Y�ke]��`��sd�z�g�2ak�c�n�+0r��u��x��2|�a|�`��;��������5��H͇��b������҆�����K����.��渒�dA��gȕ�N��yҘ��U���כ�Y��gٞ��X��}ס��U���Ҥ��O�� ̧�H���ê�*?��^���r5��t����+�������!��������Ŕ����ꍼ�:���  �  ��N=��M=�M=eCL=��K=H�J=yJ=6AI=PH=޼G=��F= 6F=�qE=X�D=_�C=�C=�WB=*�A=��@=��?=J/?=�b>=v�==G�<=��;=�";=�O:=�z9=��8=��7=7�6=�6=�:5=�[4=�z3=
�2=�1=��0=$�/=0�.=�.=�-=^#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=i#=S�!=�� =(�=٪=��=hb=8=�	=�=�=�d=%=��=v�=^K=��=��=�H=��=�
=�	=�=�?=]�=wP=>�=�O =d��<�|�<�_�<W:�<��<3��<���<$[�<��<���<�k�<;�<��<�D�<���<�d�<���<Vq�<���<�k�<�<dV�<LƳ<�2�<l��<1�<3g�<�ȡ<e(�<څ�<��<�;�<͔�<��<zC�<���<V�<e�z<�3s<��k<2�d<�6]<��U<q�N<�FG<H�?<1�8<kn1<�-*<#�"<��<��<�Y<3<�$�;���;��;׷�;���;��;Tߩ;]�;�W�;���;�Gf;NWK;u�0;�;�Q�:��:W�:�M7:���9�k������[�m����<Ϻ�M���l�k�.��*F��!]���s����S-��j���᥻<������`ŻX�ϻp�ٻa�㻀f���MK �p���	��/�9��� ����+���$��I(�Ro,�?�0�x�4�ǎ8�o<��c@� <D��H���K�q�O��-S���V��iZ�&�]��a�.�d�th�7�k��Ho��r�� v�rRy���|�p�������.��UɄ�`a������������Q����8���ď��N���֒��]��a㕼�g���꘼~l��G훼m��잼j���硼Od��r़&\��Uק�'R���̪��F�������:��Ŵ���.�������"��������k������Z�������  �  ��N=��M=�M=jCL=��K=A�J=yJ=)AI=NH=ܼG=��F=6F=�qE=[�D=^�C=�C=�WB=4�A=��@=��?=D/?=sb>=y�==>�<=��;=�";=�O:=�z9=��8=��7=9�6=�6=�:5=�[4=�z3=�2=�1=��0=!�/=8�.=�.=�-=b#,=-+=�3*=�7)=�8(=�6'=}1&=�(%=�$=d#=X�!=�� =-�=ݪ=��=lb= 8=�	=��=�=�d=%= �=l�=_K=��=��=I=��=�
=�	=�=�?=`�=rP=;�=�O =R��<�|�<�_�<^:�<��<=��<���</[�<��<���<�k�<%�<٬�<�D�<���<e�<���<\q�<���<�k�<�<tV�<TƳ<�2�<l��<�<.g�<�ȡ<U(�<ㅚ<��<�;�<Д�<��<wC�<���<K�<K�z<�3s<��k<<�d<�6]<��U<��N<�FG<T�?<1�8<~n1<�-*<8�"<p�<ۆ<�Y<�2<�$�;���;!��;��;���;3��;Jߩ;l�;�W�;粀;�Gf;\WK;�0;�; R�:� �:��:O7:��9a�����[�7���U<ϺsN��m�t�.�+F�\!]�N�s����-��N��j᥻������`ŻF�ϻ��ٻZ�㻫f�
��JK ����ߞ	��/�%��� �������$��I(�_o,�:�0���4���8�g<��c@��;D��H�r�K�_�O��-S�~�V�oiZ�)�]��a�"�d�'th�?�k��Ho�7�r�� v�fRy��|�r�������.��JɄ�ca�� ���������a����8���ď��N���֒��]��a㕼�g���꘼nl��?훼m��잼8j���硼Zd���़\��Nק�R���̪��F�������:��д���.�������"��������w������\�������  �  ��N=��M=�M=iCL=��K=D�J=�J=)AI=WH=ܼG=��F=6F=�qE=]�D=^�C=�C=�WB=4�A=��@=��?=L/?=tb>=��==?�<=��;=�";=�O:=�z9=��8=��7=3�6=�6=�:5=�[4=�z3=�2=��1=��0=!�/=6�.=�.=�-=[#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=b#=Y�!=�� =)�=ڪ=��=jb=8=�	=��=�=�d=%=�=k�=aK=��=��=�H=��=�
=�	=�=�?=f�=qP==�=�O =U��<�|�<�_�<X:�<z�<4��<���<'[�<��<���<�k�<,�<��<�D�<���<e�<���<\q�<���<�k�<�<pV�<TƳ<�2�<~��<�<<g�<�ȡ<V(�<ᅚ<��<�;�<Ô�<��<nC�<���<L�<Y�z<4s<��k<T�d<�6]<��U<��N<�FG<P�?<�8<nn1<�-*<5�"<t�<�<Z<�2<%�;���;��;��;m��;I��;Pߩ;{�;�W�;벀;�Gf;�WK;��0;;/S�:� �:<�:aN7:]��9ci����L[�٦��K<Ϻ4N���l�F�.�4+F�� ]�8�s����&-��w���᥻P������#`Ż<�ϻ��ٻ"�㻁f����%K ����ܞ	��/�4��� ����"���$��I(�do,��0���4�Ɏ8�I<��c@��;D��H���K�y�O�.S���V�|iZ�'�]��a��d�)th�7�k��Ho�/�r�� v�xRy���|���������.��QɄ�_a��!����������T����8���ď��N���֒��]��b㕼�g���꘼sl��?훼m���랼5j���硼Pd���़ \��Wק�(R���̪��F�������:��ϴ���.�������"��������u������f�������  �  ��N=��M=�M=fCL=��K=F�J=wJ=-AI=OH=߼G=��F=6F=�qE=_�D=a�C=�C=�WB=2�A=��@=��?=G/?=xb>=s�==E�<=��;=�";=�O:=�z9=��8=��7=7�6=�6=�:5=�[4=�z3=�2=�1=��0=�/=3�.=�.=�-=`#,=-+=�3*=�7)=�8(=�6'=1&=�(%=�$=i#=[�!=�� =+�=ߪ=��=kb=8=�	=�=�=�d=%=��=t�=\K=��=��=I=��=�
=�	=�=�?=X�=rP=9�=�O =\��<�|�<�_�<Z:�<��<;��<���<([�<��<���<�k�</�<��<�D�<���<e�<���<]q�<���<�k�<�<qV�<ZƳ<�2�<l��<"�<.g�<�ȡ<d(�<م�<��<�;�<˔�<��<vC�<���<I�<[�z<�3s<��k<*�d<�6]<��U<g�N<�FG<T�?<*�8<un1<�-*<&�"<��<�<�Y<�2<�$�;���;:��;��;���;Y��;dߩ;}�;�W�;ݲ�;'Hf;eWK;M�0;b;yQ�:��:��:kN7:Z��9fd�����[�b���G=Ϻ�M��m���.��*F��!]��s����=-��^��d᥻+������`Żg�ϻt�ٻh�㻞f����HK �m��Ҟ	��/�-��� �������$��I(�Fo,�3�0���4�ӎ8�v<��c@�<D��H�v�K�c�O��-S���V��iZ�7�]��a�=�d�&th�H�k��Ho� �r�� v�nRy���|�h�������.��OɄ�_a������������Z����8��{ď��N���֒��]��[㕼�g���꘼ql��9훼m��잼-j���硼Sd��r़(\��Mק�!R���̪��F�������:��Ҵ���.�������"��������u������]�������  �  ��N=��M=�M=fCL=��K=F�J=xJ=6AI=NH=�G=��F=6F=�qE=\�D=b�C=�C=�WB=1�A=��@=��?=H/?=�b>=v�==F�<=��;=�";=�O:=�z9=��8=��7=:�6=�6=�:5=�[4=�z3=�2=�1=��0=�/=8�.=�.=�-=\#,=-+= 4*=�7)=�8(=�6'=�1&=�(%=�$=l#=W�!=�� =+�=ߪ=��=jb=!8=�	=�=�=�d=%=��=u�=WK=��=��=�H=��=�
=�	=�=�?=V�=sP=8�=�O =Z��<�|�<�_�<G:�<|�</��<���<,[�<��<���<�k�<=�<��<�D�<���<�d�<���<[q�<���<�k�<�<qV�<SƳ<�2�<n��<2�<0g�<�ȡ<a(�<م�<��<�;�<Ɣ�<��<tC�<���<B�<U�z<�3s<��k<�d<�6]<��U<i�N<�FG<0�?<#�8<[n1<�-*<)�"<{�<��<�Y<3<�$�;���;%��;��;���;@��;nߩ;l�;�W�;Բ�;Hf;�WK;[�0;�;�Q�:��:��:�N7:���9cp��7�﹜ [�󥞺P=ϺN��m���.��*F��!]��s����-��y���᥻F�������_Ży�ϻp�ٻ`��vf���FK �a���	��/�,��� �������$��I(�Do,�2�0�{�4���8�t<��c@�<D��H���K�t�O�.S���V�qiZ�D�]��a�E�d� th�J�k��Ho�"�r�� v�`Ry��|��������.��KɄ�la������������U����8��|ď��N���֒��]��Y㕼�g���꘼ql��A훼m��잼j���硼Sd��v़(\��Jק�/R���̪��F�������:��ٴ���.�������"��������|������\�������  �  ��N=��M=�M=hCL=��K=E�J=}J=.AI=VH=޼G=��F=6F=�qE=b�D=f�C=�C=�WB=9�A=��@=��?=K/?=wb>=}�==@�<=��;=�";=�O:=�z9=��8=��7=2�6=�6=�:5=�[4=�z3=��2=�1=��0=�/=4�.=�.=�-=_#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=d#=^�!=�� =-�=�=��=nb=!8=�	=��=�=�d=%=�=m�=^K=��=��=�H=��=�
=�	=�=�?=\�=kP=5�=�O =A��<�|�<�_�<M:�<��<5��<���<*[�<��<���<�k�<+�<��<�D�<���<e�<���<eq�<���<�k�<�<|V�<YƳ<�2�<}��<!�<6g�<�ȡ<U(�<���<��<�;�<˔�<��<hC�<���<<�<@�z<�3s<��k<2�d<�6]<��U<z�N<�FG<B�?<)�8<in1<�-*<1�"<r�<�<�Y<�2<%�;���;'��;F��;���;u��;�ߩ;��;�W�;��;�Gf;�WK;��0;U;�R�:� �:G�:O7:�9�g��r��s[�ڦ���<ϺUO��0m���.�W+F�f!]���s����/-�����x᥻)������`ŻD�ϻ��ٻ=�㻌f����-K ����ƞ	��/� ��� �}�����$��I(�do,� �0���4�ю8�Y<��c@��;D��H���K�g�O��-S���V��iZ�:�]��a�+�d�<th�R�k��Ho�Q�r�� v�Ry��|�q�������.��LɄ�ba������������V����8���ď�yN���֒��]��S㕼�g���꘼gl��;훼m���랼.j���硼Qd���़!\��Uק�(R���̪��F������:��޴���.�������"���������������j�������  �  ��N=��M=�M=iCL=��K=C�J=�J=,AI=ZH=ݼG=��F=6F=�qE=g�D=_�C=�C=�WB=?�A=��@=��?=O/?=wb>=��==>�<=��;=�";=�O:=�z9=��8=��7=+�6=�6=�:5=�[4=�z3=��2=�1=��0=%�/=.�.=�.=�-=X#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=d#=g�!=�� =/�=�=��=rb=8=�	=��=�=�d=%=�=k�=cK=��=��=�H=��=�
=�	=�=�?=Z�=iP=5�=�O =>��<�|�<u_�<V:�<s�<5��<���<![�<��<���<�k�<,�<��<�D�<���<e�<���<qq�<���<�k�<�<|V�<nƳ<�2�<���<"�<>g�<�ȡ<Z(�<煚<��<�;�<���<��<`C�<���<H�<)�z<�3s<��k<.�d<�6]<��U<w�N<jFG<P�?<�8<vn1<�-*<3�"<x�<�<Z<�2<2%�;���;s��;U��;���;���;]ߩ;��;�W�;H��;IHf;�WK;֖0;Y;WS�:� �:�:kN7:r��9�a������[������;ϺO��[m���.�w+F�!]���s����]-��~���᥻g������;`Ż�ϻ��ٻ0��rf����K ������	��/���� �|�� ���$�dI(�Yo,��0���4�Ď8�P<��c@��;D��H�x�K�z�O�.S���V��iZ��]��a�2�d�Ath�Q�k��Ho�U�r�� v��Ry���|���������.��TɄ�Ta��!����������N����8��}ď�iN���֒��]��]㕼�g���꘼fl��&훼m���랼-j���硼Rd��}़\��]ק�R���̪��F��	����:��Ӵ���.�������"��������������u�������  �  ��N=��M=�M=gCL=��K=D�J=~J=6AI=UH=�G=��F=6F=�qE=h�D=c�C=�C=�WB=8�A=��@=��?=N/?=�b>=|�==B�<=��;=�";=�O:=�z9=��8=��7=+�6=�6=�:5=�[4=�z3=��2=�1=��0=�/=)�.=�.=�-=W#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=l#=_�!=�� =1�=�=��=sb="8=�	=�=�=�d=%=��=p�=]K=��=��=�H=��=
�
=�	=�=�?=U�=jP=1�=�O =B��<�|�<s_�<N:�<m�<-��<���<[�<��<���<�k�<=�<��<�D�<���<e�<���<tq�<���<�k�<�<wV�<eƳ<�2�<y��<5�<:g�<�ȡ<_(�<ޅ�<��<�;�<���<��<cC�<���<?�<3�z<�3s<��k<�d<�6]<��U<V�N<pFG<@�?<�8<gn1<�-*<)�"<{�<�<�Y<3<%�;���;k��;=��;���;���;�ߩ;��;�W�;��;�Hf;�WK;֖0;�;�R�:p�:��:�M7:a��9�h���﹠[�����+=Ϻ�N��bm���.�7+F��!]���s�����-������᥻j������'`ŻI�ϻ��ٻI��if���0K �`����	��/���� �x������$��I(�>o,� �0�p�4���8�e<��c@��;D��H���K���O�.S���V��iZ�:�]��a�C�d�<th�^�k��Ho�J�r�� v��Ry��|���������.��XɄ�`a������������L����8��rď�zN���֒��]��W㕼�g���꘼kl��/훼	m��잼j���硼Ud��x़#\��Yק�&R���̪��F����� ;��ܴ���.�������"��!�������������r�������  �  ��N=��M=�M=hCL=��K=J�J=zJ=4AI=QH=�G=��F=6F=�qE=d�D=n�C=�C=�WB=:�A=��@=�?=I/?=|b>=y�==H�<=��;=�";=�O:=�z9=��8=��7=2�6=�6=�:5=�[4=�z3=��2=�1=��0=�/=0�.=�.=�-=_#,=-+= 4*=�7)=�8(=�6'=�1&=�(%=�$=s#=[�!=�� =/�=�=��=nb=+8=�	=�=�=�d=%=�=r�=VK=��=��=�H=��=�
=�	=�=�?=P�=hP=-�=�O =<��<�|�<�_�<@:�<{�</��<���<-[�<��<���<�k�<5�<��<�D�<���<e�<���<dq�<���<�k�<�<�V�<[Ƴ<3�<p��</�<1g�<�ȡ<](�<څ�<��<�;�<̔�<~�<dC�<���</�<<�z<�3s<��k<��d<�6]<z�U<Y�N<{FG<$�?<)�8<Rn1<�-*<-�"<u�< �<�Y<3<�$�;��;F��;p��;��;���;�ߩ;��; X�;%��;�Hf;4XK;�0;�;aR�:'�:�:�O7:���98l�����u [�Ǧ���=ϺbO��km�#�.�Y+F�"]���s�7��K-������᥻)������_Żx�ϻ~�ٻ+�㻅f���:K �A��͞	�n/���� �c����u$��I(�#o,�"�0�~�4�Ŏ8�[<��c@�<D��H���K�l�O�	.S���V��iZ�_�]��a�T�d�Dth�k�k�Io�V�r�� v�Ry�!�|�z�������.��GɄ�ja������������W����8��mď�zN���֒��]��B㕼�g���꘼Yl��9훼�l��잼 j���硼Id��z़'\��Nק�4R���̪��F������:��봰��.��ͨ���"��/�������������l�������  �  ��N=��M=�M=jCL=��K=I�J=�J=6AI=[H=�G=��F=6F=�qE=f�D=j�C=�C=�WB==�A=��@=�?=Q/?=�b>=��==F�<=��;=�";=�O:=�z9=��8=��7=.�6=�6=�:5=�[4=�z3=��2=�1=��0=�/=0�.=�.=�-=X#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=p#=]�!=�� =0�=�=��=ob=+8=�	=�=�=�d=!%=�=o�=ZK=��=��=�H=��=�
=�	=�=�?=Q�=fP=-�=�O =:��<�|�<{_�<=:�<n�<'��<���<-[�<��<���<�k�<;�<��< E�<���<e�<���<iq�<���<�k�<�<�V�<[Ƴ<3�<���<6�<>g�<�ȡ<Z(�<䅚<��<�;�<���<�<]C�<���<1�<.�z<�3s<��k<	�d<�6]<z�U<`�N<kFG<$�?<�8<Jn1<�-*<8�"<r�<��<Z<3<7%�;��;F��;���;��;���;�ߩ;��;*X�;D��;^Hf;OXK;�0;�;US�:��:5�:<P7:-��91n��_�﹚ [�2���=ϺdO���m��.�g+F�	"]���s���H-������᥻c������_ŻD�ϻ��ٻ"��Xf�}��K �N��ƞ	�m/���� �f����v$��I(�3o,�
�0�_�4���8�L<��c@�<D��H���K���O�.S���V��iZ�O�]��a�P�d�Ith�k�k�Io�X�r�� v��Ry�$�|���������.��FɄ�ga������������F����8��vď�tN���֒��]��J㕼�g���꘼Sl��8훼 m���랼j���硼Jd��}़\��Qק�9R���̪��F������:��鴰��.��Ǩ���"��(�������������s�������  �  ��N=��M=�M=gCL=��K=D�J=J=1AI=ZH=�G=��F=6F=�qE=p�D=d�C=�C=�WB=?�A=��@=�?=P/?=|b>=|�==A�<=��;=�";=�O:=�z9=��8=��7=)�6=�6=�:5=�[4=�z3=��2=�1=��0=�/=*�.=�.=�-=W#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=o#=c�!=�� =:�=�=��=|b=(8=�	=�=�=�d=%=��=l�=^K=��=��=�H=��=�
=�	=�=�?=O�=aP=(�=�O =4��<�|�<l_�<O:�<h�<.��<���<[�<��<���<�k�<3�<��<�D�<���<e�<���<�q�<���<l�<&�<�V�<lƳ<�2�<���<*�<:g�<�ȡ<^(�<߅�<��<�;�<���<��<`C�<���<4�<�z<�3s<��k<�d<z6]<}�U<R�N<gFG<A�?<��8<wn1<�-*<,�"<}�<�<�Y<3<0%�;���;���;���;���;���;�ߩ;.�;#X�;W��;�Hf;XK;��0;�;�R�:[�:��:;N7:���9b��3��I[�ۧ��l=Ϻ�O���m�5�.��+F�"]���s���x-������᥻f������;`Ż=�ϻ��ٻI�㻂f���!K �T����	�|/���| �b������$�uI(�1o,��0�}�4�Ȏ8�a<��c@��;D��H�q�K�~�O�.S���V��iZ�O�]�%�a�V�d�]th�}�k�Io�d�r�� v��Ry���|���������.��WɄ�]a������������K����8��pď�oN���֒��]��S㕼vg��x꘼Xl��(훼m���랼&j���硼Td��z़"\��[ק�R���̪��F��	���;��洰��.��Ȩ���"��*�������������v�������  �  ��N=��M=�M=fCL=��K=J�J=�J=7AI=ZH=�G=��F=6F=�qE=j�D=i�C=�C=�WB=?�A=��@=�?=Q/?=�b>=��==E�<=��;=�";=�O:=�z9=��8=��7=*�6=�6=�:5=�[4=�z3=��2=�1=��0=�/=+�.=�.=�-=S#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=s#=b�!=�� =4�=�=��=ub=&8=�	=�=�=�d=!%=�=p�=\K=��=��=�H=��=�
=�	=�=�?=P�=cP=*�=�O =:��<�|�<p_�<=:�<b�<$��<���<[�<��<���<�k�<?�<��<E�<���<e�<���<vq�<���<�k�<�<�V�<kƳ<3�<���<4�<Bg�<�ȡ<b(�<ۅ�<��<�;�<���<y�<[C�<���<4�<-�z<�3s<��k<��d<�6]<~�U<T�N<bFG<"�?<��8<Vn1<�-*<'�"<��<��<Z<3<6%�;��;���;~��;۳�;���;�ߩ;��;X�;U��;�Hf;dXK;
�0;-;jS�:��:��:.N7:듢9+o�����k [�����p=Ϻ-O��Xm�5�.��+F�"]���s���l-������᥻�������5`ŻL�ϻ~�ٻ��Uf���K �C����	��/� ��� �d������$�yI(�"o,� �0�j�4���8�D<��c@��;D��H���K���O�+.S���V��iZ�W�]��a�R�d�Tth�u�k��Ho�U�r�� v��Ry�#�|���������.��XɄ�^a������������G����8��mď�nN���֒��]��K㕼}g���꘼\l��)훼�l���랼j���硼Gd��u़%\��]ק�.R���̪��F������:��洰��.��̨���"��0�������������x�������  �  ��N=��M=�M=kCL=��K=E�J=~J=7AI=WH=�G=��F=6F=�qE=i�D=r�C=�C=�WB=C�A=��@=�?=M/?=�b>=|�==B�<=��;=�";=�O:=�z9=��8=��7=.�6=�6=�:5=�[4=�z3=��2=�1=��0=�/=+�.=�.=�-=\#,=-+=4*=�7)=�8(=�6'=�1&=�(%=�$=o#=a�!=�� =5�=�=��=tb=08=�	=�=�=�d=%=�=m�=[K=��=��=�H=��=�
=�	=�=�?=L�=aP=%�=�O =.��<�|�<z_�<;:�<z�<.��<���<,[�<��<���<�k�<9�<��<�D�<���< e�<���<oq�<���<�k�<%�<�V�<bƳ<3�<��<4�<9g�<�ȡ<W(�<ㅚ<��<�;�<͔�<��<[C�<���<!�<)�z<�3s<��k<�d<�6]<^�U<H�N<gFG<.�?<'�8<Pn1<�-*<;�"<m�<�<�Y<3<%�;��;_��;���;���;���;�ߩ;��;KX�;y��;WHf;pXK;Ԗ0;;�R�:��:]�:UP7:��9�g�����~ [�,���>ϺP���m���.��+F�B"]���s�[��o-������᥻;�������_ŻE�ϻ��ٻ,��wf���"K �R����	�]/����x �V�����a$�xI(�:o,��0�o�4���8�U<��c@��;D��H���K�w�O�.S���V��iZ�s�]��a�a�d�[th���k�Io�n�r�� v��Ry�&�|�y�������.��FɄ�ca������������O����8��{ď�hN���֒��]��=㕼}g��y꘼Ml��2훼�l���랼j���硼Pd���़\��Mק�4R���̪��F�����;�������.��Ϩ���"��5�������������u�������  �  ��N=��M=�M=fCL=��K=J�J=�J=7AI=ZH=�G=��F=6F=�qE=j�D=i�C=�C=�WB=?�A=��@=�?=Q/?=�b>=��==E�<=��;=�";=�O:=�z9=��8=��7=*�6=�6=�:5=�[4=�z3=��2=�1=��0=�/=+�.=�.=�-=S#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=s#=b�!=�� =4�=�=��=ub=&8=�	=�=�=�d=!%=�=p�=\K=��=��=�H=��=�
=�	=�=�?=P�=cP=*�=�O =:��<�|�<q_�<=:�<b�<$��<���<[�<��<���<�k�<?�<��<E�<���<e�<���<vq�<���<�k�<�<�V�<kƳ<3�<���<4�<Bg�<�ȡ<b(�<ۅ�<��<�;�<���<y�<[C�<���<4�<,�z<�3s<��k<��d<�6]<~�U<T�N<bFG<"�?<��8<Wn1<�-*<'�"<��<��<Z<3<6%�;��;���;~��;ܳ�;���;�ߩ;��;X�;U��;�Hf;cXK;
�0;,;hS�:��:��:*N7:ⓢ9Mo�� ��o [�����r=Ϻ/O��Ym�6�.��+F�"]���s���l-������᥻�������5`ŻL�ϻ~�ٻ��Uf���K �C����	��/� ��� �d������$�yI(�"o,� �0�j�4���8�D<��c@��;D��H���K���O�+.S���V��iZ�W�]��a�R�d�Tth�u�k��Ho�U�r�� v��Ry�#�|���������.��XɄ�^a������������G����8��mď�nN���֒��]��K㕼}g���꘼\l��)훼�l���랼j���硼Gd��u़%\��]ק�.R���̪��F������:��洰��.��̨���"��0�������������x�������  �  ��N=��M=�M=gCL=��K=D�J=J=1AI=ZH=�G=��F=6F=�qE=p�D=d�C=�C=�WB=?�A=��@=�?=P/?=|b>=|�==A�<=��;=�";=�O:=�z9=��8=��7=)�6=�6=�:5=�[4=�z3=��2=�1=��0=�/=*�.=�.=�-=W#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=o#=c�!=�� =:�=�=��=|b=(8=�	=�=�=�d=%=��=l�=^K=��=��=�H=��=�
=�	=�=�?=O�=aP=(�=�O =4��<�|�<l_�<P:�<h�</��<���<[�<��<���<�k�<3�<��<�D�<���<e�<���<�q�<���<l�<&�<�V�<lƳ<�2�<���<*�<:g�<�ȡ<](�<߅�<��<�;�<���<��<_C�<���<4�<�z<�3s<��k<�d<z6]<}�U<R�N<gFG<A�?<��8<wn1<�-*<,�"<}�<�<�Y<3<1%�;���;���;���;���;���;�ߩ;-�;#X�;V��;�Hf;XK;��0;�;�R�:X�:��:3N7:q��9Gb��D��Q[�ߧ��p=Ϻ�O���m�7�.��+F�"]���s���y-������᥻f������<`Ż=�ϻ��ٻJ�㻂f���!K �T����	�|/���| �b������$�uI(�1o,��0�}�4�Ȏ8�a<��c@��;D��H�q�K�~�O�.S���V��iZ�O�]�%�a�V�d�]th�}�k�Io�d�r�� v��Ry���|���������.��WɄ�]a������������K����8��pď�oN���֒��]��S㕼vg��x꘼Xl��(훼m���랼&j���硼Td��z़"\��[ק�R���̪��F��	���;��洰��.��Ȩ���"��*�������������v�������  �  ��N=��M=�M=jCL=��K=I�J=�J=6AI=[H=�G=��F=6F=�qE=f�D=j�C=�C=�WB==�A=��@=�?=Q/?=�b>=��==F�<=��;=�";=�O:=�z9=��8=��7=.�6=�6=�:5=�[4=�z3=��2=�1=��0=�/=0�.=�.=�-=X#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=p#=]�!=�� =0�=�=��=ob=+8=�	=�=�=�d=!%=�=o�=ZK=��=��=�H=��=�
=�	=�=�?=Q�=fP=-�=�O =:��<�|�<{_�<=:�<n�<'��<���<-[�<��<���<�k�<;�<��< E�<���<e�<���<jq�<���<�k�<�<�V�<[Ƴ<3�<���<6�<>g�<�ȡ<Z(�<䅚<��<�;�<���<�<]C�<���<1�<-�z<�3s<��k<	�d<�6]<{�U<`�N<lFG<$�?<�8<Kn1<�-*<8�"<r�<��<Z<3<7%�;��;F��;���;��;���;�ߩ;��;*X�;D��;\Hf;NXK;�0;�;PS�:��:0�:1P7:��9�n��w�﹥ [�8���=ϺjO���m�
�.�i+F�"]���s���I-������᥻d������_ŻD�ϻ��ٻ"��Xf�}��K �N��ƞ	�m/���� �f����v$��I(�3o,�
�0�_�4���8�L<��c@�<D��H���K���O�.S���V��iZ�O�]��a�P�d�Ith�k�k�Io�X�r�� v��Ry�$�|���������.��FɄ�ga������������F����8��vď�tN���֒��]��J㕼�g���꘼Sl��8훼 m���랼j���硼Jd��}़\��Qק�9R���̪��F������:��鴰��.��Ǩ���"��(�������������s�������  �  ��N=��M=�M=hCL=��K=J�J=zJ=4AI=QH=�G=��F=6F=�qE=d�D=n�C=�C=�WB=:�A=��@=�?=I/?=|b>=y�==H�<=��;=�";=�O:=�z9=��8=��7=2�6=�6=�:5=�[4=�z3=��2=�1=��0=�/=0�.=�.=�-=_#,=-+= 4*=�7)=�8(=�6'=�1&=�(%=�$=s#=[�!=�� =/�=�=��=nb=+8=�	=�=�=�d=%=�=r�=VK=��=��=�H=��=�
=�	=�=�?=P�=hP=-�=�O =<��<�|�<�_�<@:�<|�<0��<���<-[�<��<���<�k�<5�<��<�D�<���<e�<���<dq�<���<�k�<�<�V�<ZƳ<3�<p��</�<1g�<�ȡ<](�<څ�<��<�;�<̔�<~�<dC�<���</�<<�z<�3s<��k<��d<�6]<{�U<Y�N<{FG<$�?<)�8<Sn1<�-*<-�"<u�< �<�Y<3<�$�;��;F��;q��;��;���;�ߩ;��; X�;%��;�Hf;2XK;}�0;�;[R�:!�:�:�O7:k��9�l����﹃ [�Φ���=ϺiO��nm�&�.�\+F�"]���s�8��L-������᥻*������_Żx�ϻ�ٻ,�㻅f���;K �A��͞	�n/���� �c����u$��I(�#o,�"�0�~�4�Ŏ8�[<��c@�<D��H���K�m�O�	.S���V��iZ�_�]��a�T�d�Dth�k�k�Io�V�r�� v�Ry�!�|�z�������.��GɄ�ja������������W����8��mď�zN���֒��]��B㕼�g���꘼Yl��9훼�l��잼 j���硼Id��z़'\��Nק�4R���̪��F������:��봰��.��ͨ���"��/�������������l�������  �  ��N=��M=�M=gCL=��K=D�J=~J=6AI=UH=�G=��F=6F=�qE=h�D=c�C=�C=�WB=8�A=��@=��?=N/?=�b>=|�==B�<=��;=�";=�O:=�z9=��8=��7=+�6=�6=�:5=�[4=�z3=��2=�1=��0=�/=)�.=�.=�-=W#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=l#=_�!=�� =1�=�=��=sb="8=�	=�=�=�d=%=��=p�=]K=��=��=�H=��=
�
=�	=�=�?=U�=jP=1�=�O =C��<�|�<t_�<O:�<n�<.��<���<[�<��<���<�k�<=�<��<�D�<���<e�<���<tq�<���<�k�<�<wV�<eƳ<�2�<y��<5�<9g�<�ȡ<_(�<݅�<��<�;�<���<��<cC�<���<?�<3�z<�3s<��k<�d<�6]<��U<V�N<pFG<@�?<�8<hn1<�-*<*�"<{�<�<�Y<3<%�;���;k��;=��;���;���;�ߩ;��;�W�;��;�Hf;�WK;Ӗ0;�;�R�:i�:��:�M7:A��9Ki��$�ﹰ[�����3=Ϻ�N��fm���.�:+F��!]���s�����-������᥻k������(`ŻJ�ϻ��ٻI��if���0K �`����	��/���� �x������$��I(�>o,� �0�p�4���8�e<��c@��;D��H���K���O�.S���V��iZ�:�]��a�C�d�<th�^�k��Ho�J�r�� v��Ry��|���������.��XɄ�`a������������L����8��rď�zN���֒��]��W㕼�g���꘼kl��/훼	m��잼j���硼Ud��x़#\��Yק�&R���̪��F����� ;��ܴ���.�������"��!�������������r�������  �  ��N=��M=�M=iCL=��K=C�J=�J=,AI=ZH=ݼG=��F=6F=�qE=g�D=_�C=�C=�WB=?�A=��@=��?=O/?=wb>=��==>�<=��;=�";=�O:=�z9=��8=��7=+�6=�6=�:5=�[4=�z3=��2=�1=��0=%�/=.�.=�.=�-=X#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=d#=g�!=�� =/�=�=��=rb=8=�	=��=�=�d=%=�=k�=dK=��=��=�H=��=�
=�	=�=�?=Z�=jP=5�=�O =?��<�|�<u_�<W:�<t�<5��<���<"[�<��<���<�k�<,�<��<�D�<���<e�<���<qq�<���<�k�<�<|V�<mƳ<�2�<���<"�<>g�<�ȡ<Z(�<煚<��<�;�<���<��<`C�<���<G�<)�z<�3s<��k<.�d<�6]<��U<x�N<kFG<P�?<�8<vn1<�-*<3�"<y�<�<Z<�2<3%�;���;t��;V��;���;���;]ߩ;��;�W�;H��;GHf;�WK;Ӗ0;V;PS�:� �:�:[N7:R��9b������[�Ƨ���;ϺO��_m���.�{+F��!]���s����^-�����᥻h������<`Ż�ϻ��ٻ1��rf����K ������	��/���� �|�� ���$�dI(�Yo,��0���4�Ď8�P<��c@��;D��H�y�K�z�O�.S���V��iZ��]��a�2�d�Ath�Q�k��Ho�U�r�� v��Ry���|���������.��TɄ�Ta��!����������N����8��}ď�iN���֒��]��]㕼�g���꘼fl��&훼m���랼-j���硼Rd��}़\��]ק�R���̪��F��	����:��Ӵ���.�������"��������������u�������  �  ��N=��M=�M=hCL=��K=E�J=}J=.AI=VH=޼G=��F=6F=�qE=b�D=f�C=�C=�WB=9�A=��@=��?=K/?=wb>=}�==@�<=��;=�";=�O:=�z9=��8=��7=2�6=�6=�:5=�[4=�z3=��2=�1=��0=�/=4�.=�.=�-=_#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=d#=^�!=�� =-�=�=��=nb=!8=�	=��=�=�d=%=�=m�=^K=��=��=�H=��=�
=�	=�=�?=\�=kP=5�=�O =B��<�|�<�_�<N:�<��<6��<���<+[�<��<���<�k�<,�<��<�D�<���<e�<���<eq�<���<�k�<�<{V�<XƳ<�2�<}��<!�<6g�<�ȡ<U(�<���<��<�;�<˔�<��<gC�<���<<�<@�z<�3s<��k<2�d<�6]<��U<z�N<�FG<B�?<*�8<jn1<�-*<2�"<r�<�<�Y<�2<%�;���;'��;G��;���;u��;�ߩ;��;�W�;��;�Gf;�WK;��0;R;�R�:� �:@�:O7:ԓ�9h����﹃[�ᦞ��<Ϻ]O��4m���.�Z+F�i!]���s����1-�����y᥻*������`ŻE�ϻ��ٻ=�㻌f����-K ����ƞ	��/�!��� �}�����$��I(�do,� �0���4�ю8�Y<��c@��;D��H���K�g�O��-S���V��iZ�:�]��a�+�d�<th�R�k��Ho�Q�r�� v�Ry��|�q�������.��LɄ�ba������������V����8���ď�yN���֒��]��S㕼�g���꘼gl��;훼m���랼.j���硼Qd���़!\��Uק�(R���̪��F������:��޴���.�������"���������������j�������  �  ��N=��M=�M=fCL=��K=F�J=xJ=6AI=NH=�G=��F=6F=�qE=\�D=b�C=�C=�WB=1�A=��@=��?=H/?=�b>=v�==F�<=��;=�";=�O:=�z9=��8=��7=:�6=�6=�:5=�[4=�z3=�2=�1=��0=�/=8�.=�.=�-=\#,=-+= 4*=�7)=�8(=�6'=�1&=�(%=�$=l#=W�!=�� =+�=ߪ=��=jb=!8=�	=�=�=�d=%=��=u�=WK=��=��=�H=��=�
=�	=�=�?=V�=sP=8�=�O =Z��<�|�<�_�<G:�<}�<0��<���<,[�<��<���<�k�<=�<��<�D�<���<�d�<���<[q�<���<�k�<�<qV�<SƳ<�2�<m��<2�<0g�<�ȡ<a(�<م�<��<�;�<Ɣ�<��<tC�<���<B�<U�z<�3s<��k<�d<�6]<��U<i�N<�FG<0�?<#�8<[n1<�-*<)�"<|�<�<�Y<3<�$�;���;%��;��;���;@��;nߩ;l�;�W�;Ӳ�;Hf;�WK;X�0;�;�Q�:��:��:�N7:���9�p��T�﹪ [�����W=Ϻ
N��m���.��*F��!]��s����-��{���᥻G�������_Ży�ϻp�ٻa��vf���FK �b���	��/�,��� �������$��I(�Eo,�2�0�{�4���8�t<��c@�<D��H���K�t�O�.S���V�qiZ�D�]��a�E�d� th�J�k��Ho�"�r�� v�`Ry��|��������.��KɄ�la������������U����8��|ď��N���֒��]��Y㕼�g���꘼ql��A훼m��잼j���硼Sd��v़(\��Jק�/R���̪��F�������:��ٴ���.�������"��������|������\�������  �  ��N=��M=�M=fCL=��K=F�J=wJ=-AI=OH=߼G=��F=6F=�qE=_�D=a�C=�C=�WB=2�A=��@=��?=G/?=xb>=s�==E�<=��;=�";=�O:=�z9=��8=��7=7�6=�6=�:5=�[4=�z3=�2=�1=��0=�/=3�.=�.=�-=`#,=-+=�3*=�7)=�8(=�6'=1&=�(%=�$=i#=[�!=�� =+�=ߪ=��=kb=8=�	=�=�=�d=%=��=t�=\K=��=��=I=��=�
=�	=�=�?=Y�=rP=9�=�O =\��<�|�<�_�<Z:�<��<<��<���<([�<��<���<�k�</�<��<�D�<���<e�<���<^q�<���<�k�<�<qV�<ZƳ<�2�<l��<"�<-g�<�ȡ<d(�<م�<��<�;�<˔�<��<vC�<���<I�<[�z<�3s<��k<*�d<�6]<��U<g�N<�FG<U�?<*�8<vn1<�-*<'�"<��<�<�Y<�2<�$�;���;:��;��;���;Y��;dߩ;|�;�W�;ݲ�;%Hf;dWK;K�0;`;uQ�:|�:��:`N7:D��9�d�����![�g���M=Ϻ�M��m���.��*F��!]��s����>-��_��e᥻,������	`Żg�ϻu�ٻh�㻞f����HK �m��Ҟ	��/�-��� �������$��I(�Fo,�3�0���4�ӎ8�v<��c@�<D��H�v�K�c�O��-S���V��iZ�7�]��a�=�d�&th�H�k��Ho� �r�� v�nRy���|�h�������.��OɄ�_a������������Z����8��{ď��N���֒��]��[㕼�g���꘼ql��9훼m��잼-j���硼Sd��r़(\��Mק�!R���̪��F�������:��Ҵ���.�������"��������u������]�������  �  ��N=��M=�M=iCL=��K=D�J=�J=)AI=WH=ܼG=��F=6F=�qE=]�D=^�C=�C=�WB=4�A=��@=��?=L/?=tb>=��==?�<=��;=�";=�O:=�z9=��8=��7=3�6=�6=�:5=�[4=�z3=�2=��1=��0=!�/=6�.=�.=�-=[#,=-+=�3*=�7)=�8(=�6'=�1&=�(%=�$=b#=Y�!=�� =)�=ڪ=��=jb=8=�	=��=�=�d=%=�=k�=aK=��=��=�H=��=�
=�	=�=�?=f�=qP==�=�O =U��<�|�<�_�<X:�<z�<4��<���<'[�<��<���<�k�<,�<��<�D�<���<e�<���<]q�<���<�k�<�<pV�<TƳ<�2�<}��<�<<g�<�ȡ<V(�<ᅚ<��<�;�<�<��<nC�<���<L�<Y�z<4s<��k<T�d<�6]<��U<��N<�FG<P�?<�8<nn1<�-*<5�"<t�<�<Z<�2<%�;���;��;��;m��;I��;Pߩ;{�;�W�;검;�Gf;�WK;��0;;,S�:� �:8�:ZN7:M��9�i����T[�ަ��O<Ϻ8N���l�H�.�6+F�� ]�:�s����'-��x���᥻P������$`Ż=�ϻ��ٻ"�㻂f����%K ����ܞ	��/�4��� ����#���$��I(�do,��0���4�Ɏ8�I<��c@��;D��H���K�y�O�.S���V�|iZ�'�]��a��d�)th�7�k��Ho�/�r�� v�xRy���|���������.��QɄ�_a��!����������T����8���ď��N���֒��]��b㕼�g���꘼sl��?훼m���랼5j���硼Pd���़ \��Wק�(R���̪��F�������:��ϴ���.�������"��������u������f�������  �  ��N=��M=�M=jCL=��K=A�J=yJ=)AI=OH=ܼG=��F=6F=�qE=[�D=^�C=�C=�WB=4�A=��@=��?=D/?=sb>=y�==>�<=��;=�";=�O:=�z9=��8=��7=9�6=�6=�:5=�[4=�z3=�2=�1=��0=!�/=8�.=�.=�-=b#,=-+=�3*=�7)=�8(=�6'=}1&=�(%=�$=d#=X�!=�� =-�=ݪ=��=lb= 8=�	=��=�=�d=%= �=l�=_K=��=��=I=��=�
=�	=�=�?=`�=rP=;�=�O =R��<�|�<�_�<^:�<��<=��<���</[�<��<���<�k�<%�<٬�<�D�<���<e�<���<\q�<���<�k�<�<tV�<TƳ<�2�<l��<�<.g�<�ȡ<U(�<ㅚ<��<�;�<Д�<��<wC�<���<K�<K�z<�3s<��k<<�d<�6]<��U<��N<�FG<T�?<1�8<~n1<�-*<8�"<q�<ۆ<�Y<�2<�$�;���;!��;��;���;3��;Jߩ;l�;�W�;粀;�Gf;\WK;�0;�;R�:� �:��:
O7:��94a�����[�9���W<ϺvN��m�u�.�+F�]!]�O�s����-��N��j᥻������`ŻF�ϻ��ٻZ�㻫f�
��JK ����ߞ	��/�%��� �������$��I(�_o,�:�0���4���8�g<��c@��;D��H�r�K�_�O��-S�~�V�oiZ�)�]��a�"�d�'th�?�k��Ho�7�r�� v�fRy��|�r�������.��JɄ�ca�� ���������a����8���ď��N���֒��]��a㕼�g���꘼nl��?훼m��잼8j���硼Zd���़\��Nק�R���̪��F�������:��д���.�������"��������w������\�������  �  .�N=
�M=�M=�HL=��K=��J=�	J=*II=�H=0�G=�G=�@F=}E=��D=I�C=9-C=TfB=��A=��@=�@=$A?=Bu>=%�==��<=L
<=l9;=/g:=s�9=B�8=e�7=�7=�46=�X5={4=O�3=��2=��1=��0=E0=�/={/.=�?-=�M,=X+=�`*=�e)=$h(==g'='c&=�[%=�P$=�B#=�0"=!=� =F�=�=��=5t=�F=�==�=��=Vd=� =V�=p�=�9=��=&�=�)=��
=)]	=��=@~= =`�=P=� =��< ��<|��<ŧ�<~x�<~A�<8�<���<nq�<��<��<�e�<���<���<�#�<��<%3�<���<r/�<!��<��<Ċ�<6��<^`�<^Ƭ<�)�<>��<y�<�D�<���<��<�M�<]��<���<<K�<��<P��<��z<�(s<��k<wqd<I]<��U<�gN<G<��?<Qr8<�&1<h�)<�"<�]<j$<��<�<a7�;���;���;V��;���;ꏶ;���;�ƚ;8 �;�~;fc;�\H;ނ-;��;���:aN�:<�:�8):ȅ9�
�5��Tjj��l���"׺����{�5	3��OJ�yPa��x��;��EN��\<��{��n����(��łǻf�ѻ��ۻp�廮}�x"��R�B���
��,�˩�{�9s�t� ���$��-)��N-��a1�g5�:_9��J=��)A��D�}�H��L��2P���S�QwW��
[���^�1b���e�_i��jl���o�'s��zv��y�S}�(���Ł��`��t�������9#��ڴ��JD���ь��]���珼�o�������{�������������c�������������o|�������s���;i��㧼�\���ժ�O���ǭ��@��f���2��쪳��#������Y�����
�����������  �  (�N=�M=�M=�HL=��K=��J=�	J=#II=�H=,�G=�G=�@F=}E=��D=Q�C=@-C=TfB=��A=��@=�@='A?=:u>=&�==��<=V
<=p9;=-g:=r�9=<�8=n�7=�7=�46=�X5={4=H�3=��2=��1=��0=E0=�/=z/.=�?-=�M,=�X+=�`*=�e)=$h(=>g'=$c&=�[%=�P$=�B#=�0"=!=� =M�=�=��=7t=�F=�=D�=��=Qd=� =U�=y�=�9=��=!�=�)=��
=']	=��=<~==R�=G=� =��<��<z��<ԧ�<qx�<yA�<5�<ʽ�<�q�<{�<��<te�<���<���<�#�<��<&3�<���<�/�<0��<��<Ɋ�<8��<S`�<jƬ<�)�<<��<y�<�D�<���<��<�M�<Q��<���<9K�<���<Q��<��z<�(s<��k<kqd<L]<��U<�gN<G<�?<6r8<�&1<`�)<$�"<�]<d$<��<��<�7�;���;���;n��;���;#��;��;ǚ;6 �;B�~;�ec;�\H;�-;��;���:�M�:a=�:�9):Uǅ9x
����!hj��l���"׺����{��	3��PJ�lPa�x��;��TN��`<����������(����ǻ$�ѻ��ۻd���}�x"���Q�Y��
��,�Ʃ�]�s�h� ���$��-)��N-��a1�g5�N_9��J=��)A���D�w�H��L��2P���S�HwW�[���^�Cb�y�e��i��jl�}�o�'s��zv��y�4}�'(���Ł��`��k���s���B#��ٴ��ZD���ь��]���珼�o�������{������{������^������$�������w|�������s���-i��㧼�\���ժ�	O���ǭ��@��e���2��𪳼�#�� ���W�����"
�����������  �  &�N=�M=�M=�HL=��K=��J=�	J="II=��H=*�G=�G=�@F=�|E=��D=I�C=>-C=RfB=��A=��@=�@=+A?=:u>=/�==��<=U
<=k9;=+g:=z�9=9�8=p�7=�7=�46=�X5={4=P�3=��2=��1=��0=H0=�/=x/.=�?-=�M,=�X+=�`*=�e)=!h(=Ag'=(c&=�[%=�P$=�B#=�0"=!=� =I�=�=��=7t=�F=�=E�=��=Sd=� =Q�=z�=�9=��="�=�)=��
=#]	=��=7~==V�=M=� =��<"��<p��<ק�<nx�<�A�<5�<���<�q�<r�<��<we�<���<���<�#�<��<$3�<���<r/�<(��<��<͊�<9��<M`�<sƬ<�)�<I��<x�<�D�<���<���<�M�<L��<���<.K�< ��<P��<��z<�(s<��k<�qd<6]<��U<�gN<�G<"�?</r8<�&1<J�)<�"<�]<\$<��<��<�7�;���;���;���;m��;��;š�;�ƚ;( �;K�~;�ec;�\H;Z�-;��;���:cM�:Q=�:�8):Rƅ9�
�S���gj�{m��F"׺���{�	3��PJ��Oa�Xx�z;��ZN��q<��m�������(���ǻ,�ѻ�ۻP�廪}ﻄ"���Q�i�z�
��,�Ω�l�3s�n� ���$��-)��N-��a1�g5�E_9��J=��)A���D���H�݀L��2P���S�KwW�[���^�Vb�e�e��i��jl�{�o�('s��zv�2�y�-}�*(���Ł��`��u���t���J#��Ǵ��XD���ь��]���珼�o�������{������������Z������*�������z|��|����s���3i��#㧼�\�� ֪�O���ǭ��@��f���)2��᪳��#���c�����
�����������  �  '�N=�M=�M=�HL=��K=��J=�	J=(II=��H=.�G=�G=�@F=}E=��D=P�C=A-C=ZfB=��A=��@=�@=*A?=?u>=(�==��<=P
<=n9;=-g:=t�9=:�8=h�7=�7=�46=�X5={4=I�3=��2=��1=��0=G0=�/=v/.=�?-=�M,=�X+=�`*=�e)=#h(=:g'=)c&=�[%=�P$=�B#=�0"=!=� =O�=�=��=;t=�F=�=@�=��=Vd=� =T�=v�=�9=��= �=�)=��
=$]	=��=7~=�=T�=H=� =��<"��<n��<ǧ�<mx�<{A�<4�<Ž�<tq�<y�<��<~e�<���<���<�#�<	��<23�<���</�<0��<��<ϊ�<5��<[`�<iƬ<�)�<E��<p�<�D�<���<���<�M�<N��<���<,K�<��<P��<��z<(s<��k<gqd<!]<��U<�gN<�G<�?<3r8<�&1<S�)<#�"<�]<V$<��<�<�7�;���;���;���;���;&��;���;ǚ;j �;8�~;fc;�\H;O�-;W�;��:�M�:�<�:�9):qǅ9�
���jij�vm��"׺Ȩ�Z|�	3��PJ��Pa�:x�{;��RN���<����������(��ڂǻ2�ѻ��ۻ��廝}�i"���Q�H���
��,����W�s�Y� �t�$��-)��N-��a1�g5�8_9��J=��)A���D���H��L��2P���S�]wW�[���^�Rb���e��i��jl���o�%'s��zv�3�y�L}�*(���Ł��`��o�������B#��մ��OD���ь��]���珼�o�������{������{������X�������������q|������s���/i�� 㧼�\���ժ�O���ǭ��@��e���-2�������#�����m�����
�����������  �  (�N=�M=�M=�HL=��K=��J=�	J=)II=�H=4�G=�G=�@F=	}E=��D=T�C=>-C=]fB=��A=��@=�@='A?=>u>=%�==��<=P
<=q9;=-g:=m�9==�8=l�7=�7=�46=�X5={4=G�3=��2=��1=��0=?0=�/=w/.=�?-=�M,=|X+=�`*=�e)=(h(=?g'=%c&=�[%=�P$=�B#=�0"=!=� =K�=�=��=@t=�F=�=@�=��=Sd=� =Z�=t�= :=��=�=�)=��
=#]	=��=;~=�=T�=F=� =��<��<t��<̧�<qx�<mA�</�<ͽ�<sq�<��<��<{e�<���<���<$�<��<73�<���<�/�<'��<��<֊�<=��<e`�<bƬ<�)�<>��<~�<�D�<���<��<�M�<P��<���<2K�<���<G��<��z<t(s<��k<Wqd<F]<y�U<�gN<G<�?<8r8<�&1<[�)<"�"<�]<w$<��<�<r7�;��;��;���;ǐ�;��;%��;�ƚ;� �;[�~;�fc;�\H;(�-;U�;���:�N�:�<�:o:):zǅ9'
�2��ohj��l��V#׺����{��	3��PJ��Pa��x��;��dN��y<��|�������(����ǻ:�ѻ��ۻ_�廹}�V"���Q�.���
��,����e�"s�d� �`�$��-)��N-��a1�
g5�D_9��J=��)A���D�j�H���L��2P���S�VwW�[���^�Cb���e��i��jl���o�#'s�	{v�%�y�?}�%(���Ł��`��f�������3#��ش��QD���ь��]��x珼�o�������{�������������R�������������m|�������s���/i��㧼�\���ժ�
O���ǭ��@��o���2�������#��	���Z�����)
�����������  �  #�N=�M=�M=�HL=��K=��J=�	J=(II=��H=3�G=�G=�@F=
}E=��D=T�C=D-C=\fB=��A=��@= @=.A?==u>=.�==��<=Q
<=l9;=+g:=v�9=7�8=i�7=�7=�46=�X5=	{4=B�3=|�2=��1=��0=A0=�/=s/.=�?-=�M,=�X+=�`*=�e)= h(=Fg'=%c&=�[%=�P$=�B#=�0"=
!=� =P�=
�=��=?t=�F=�=J�=��=Rd=� =P�=u�=�9=��=�=�)=��
=]	=��=2~=�=L�=?=� =��<��<i��<ǧ�<fx�<zA�</�<���<uq�<v�<��<ye�<���<���<�#�<��<43�<���<�/�<4��<��<Պ�<B��<_`�<zƬ<�)�<E��<��<�D�<���<���<�M�<I��<���<'K�<���<C��<��z<w(s<��k<Uqd<-]<m�U<�gN<�G<	�?<!r8<�&1<P�)<�"<�]<n$<��<
�<�7�;��;
��;���;ѐ�;?��;%��;1ǚ;� �;w�~;Ufc;<]H;��-;O�;���:N�: =�:a9):ǅ9"
�����hj��m���"׺ ���{��	3�QJ��Pa�lx��;��yN���<����������(��̂ǻ:�ѻ�ۻ �建}�T"���Q�@�t�
��,����N�s�J� �d�$��-)��N-��a1�g5�F_9��J=��)A���D�}�H��L��2P���S�`wW�[���^�cb���e��i��jl���o�9's��zv�9�y�G}�/(���Ł��`��r���}���D#��ƴ��SD���ь��]���珼�o�������{������w������R�������������o|�������s���3i�� 㧼�\��֪�O���ǭ��@��r���-2�������#��	���f�����(
�����������  �  �N=�M=�M=�HL=��K=��J=�	J=#II=��H=0�G=�G=�@F=
}E=��D=R�C=K-C=ZfB=��A=��@=�@=/A?=9u>=0�==��<=X
<=m9;=)g:=r�9=/�8=l�7=�7=�46=�X5={4=C�3=x�2=��1=��0=C0=�/=v/.=�?-=|M,=�X+=�`*=�e)=h(=Dg'='c&=�[%=�P$=�B#=�0"=!=� =Q�=
�=��=;t=�F=�=J�=��=Rd=� =M�=|�=�9=��=�=�)=��
=]	=��=+~=�=H�=>=� =��<��<W��<˧�<Vx�<qA�<.�<���<�q�<n�<��<qe�<���<���<�#�<��<03�<���<�/�<>��<��<׊�<K��<Z`�<|Ƭ<�)�<K��<z�<�D�<���<���<�M�<:��<���<#K�<�<A��<��z<u(s<v�k<Uqd<]<b�U<�gN<�G<�?<r8<�&1<9�)<3�"<�]<_$<��<��<�7�;���;-��;���;ِ�;n��;��;gǚ;y �;�~;�fc;%]H;��-;�;/��:�M�:�=�:�9):9ƅ9
�_���gj�rn���"׺J��!|��	3�GQJ��Pa��x��;���N��}<�����٩���(���ǻ�ѻ�ۻ-�廧}�m"���Q�F�[�
��,����I�s�7� �q�$��-)��N-��a1�g5�E_9��J=��)A���D���H��L��2P�	�S�TwW�9[���^�}b���e��i��jl���o�O's��zv�Z�y�<}�=(���Ł��`��x���n���J#��ƴ��ZD���ь��]���珼�o�������{������n������P�������������z|��z����s���#i��.㧼�\��֪�O���ǭ��@��u���52�������#��	���o�����(
�����������  �  !�N=�M=�M=�HL=��K=��J=�	J=)II=��H=5�G=�G=�@F=}E=��D=W�C=L-C=_fB=��A=��@=�@=0A?=Au>=/�==��<=O
<=l9;=-g:=p�9=5�8=l�7=�7=�46=�X5={4=?�3=z�2=��1=��0=<0=�/=v/.=�?-=M,=�X+=�`*=�e)="h(=Cg'=+c&=�[%=�P$=�B#=�0"=!=� =Q�=�=��=At=�F=�=G�=��=Wd=� =T�=t�=�9=��=�=�)=��
=]	=��=-~=�=H�=;=�� =��<��<Y��<ʧ�<]x�<jA�<2�<���<pq�<�<��<e�<���<���<$�<��<;3�<���<�/�<<��<��<���<H��<h`�<uƬ<�)�<P��<��<�D�<���<���<�M�<B��<���<'K�<을<4��<��z<\(s<�k<=qd<]<N�U<gN<�G<�?<r8<�&1<H�)<�"<�]<t$<��<�<�7�;��;*��;΢�; ��;p��;F��;pǚ;� �;��~;�fc;:]H;у-;��;��:�N�:�<�:�9):�ȅ9R
�����gj�n��^#׺E��E|�
3�"QJ��Pa��x��;���N��w<����������(����ǻ+�ѻ��ۻ2�廄}�;"���Q�%�^�
��,����G�s�/� �W�$��-)��N-��a1��f5�0_9��J=��)A���D���H��L��2P��S�VwW�8[���^�pb���e��i��jl���o�I's�{v�R�y�=}�5(���Ł��`��v�������9#��Ǵ��KD���ь��]��w珼�o�������{������o������G�������������k|��u����s���1i��&㧼�\��	֪�O���ǭ��@������22������#�����n��'���/
�����������  �  "�N=�M=�M=�HL=��K=��J=�	J=/II=��H=;�G=�G=�@F=}E=��D=\�C=J-C=gfB=��A=��@=@=2A?=Du>='�==��<=Q
<=r9;=)g:=m�9=6�8=`�7=�7=�46=�X5= {4=8�3=y�2=��1=��0=90=�/=n/.=�?-=M,=yX+=�`*=�e)=(h(=Bg'=%c&=�[%=�P$=�B#=�0"=!=� =Y�=�=��=It=�F=�=I�=��=Rd=� =Y�=r�=�9=��=�=�)=��
=]	=��=.~=�=D�=5=ۊ =��<���<a��<���<]x�<hA�<#�<Ƚ�<pq�<��<��<�e�<���<���<
$�<��<K3�<���<�/�<B��<��<銷<F��<t`�<zƬ<�)�<>��<��<�D�<���<��<�M�<E��<���<!K�<�<2��<��z<@(s<��k<"qd<]<M�U<�gN<�G<��?<r8<�&1<U�)<!�"<�]<{$<��<)�<�7�;L��;%��;��;(��;|��;p��;iǚ;� �;�~;�fc;�]H;�-;��;(��:;O�:3=�:;):�ƅ9�
�l���jj��m���#׺1��h|�n
3�8QJ�QQa�}x��;��vN���<����������(����ǻ8�ѻ��ۻ=�廴}�"���Q��l�
��,����(��r�,� �8�$��-)��N-��a1��f5�A_9��J=��)A���D�m�H��L��2P��S�{wW� [�ϕ^�kb���e��i�kl���o�D's�{v�B�y�k}�4(���Ł��`��g������1#��մ��ID���ь��]��s珼�o��u����{������h������>�������������^|�������s���0i��㧼�\��֪� O���ǭ��@������32������#��"���p��(���.
�����������  �  #�N=�M=�M=�HL=��K=��J=�	J=-II=��H=7�G=�G=�@F=
}E=��D=]�C=L-C=afB=��A=��@=@=/A?=Cu>=-�==��<=Q
<=n9;="g:=q�9=4�8=b�7=�7=�46=�X5={4==�3=w�2=��1=��0=60=�/=k/.=�?-=�M,={X+=�`*=�e)=#h(=Eg'=+c&=�[%=�P$=�B#=�0"=!=� =Y�=�=��=Et=�F=�=F�=��=Ud=� =R�=s�=�9=��=�=�)=��
=]	=��=)~=�=D�=9=݊ =��<���<T��<���<Xx�<oA�<�<���<qq�<{�<��<�e�<���<���<$�<(��<@3�<���<�/�<H��<��<銷<Z��<k`�<sƬ<�)�<L��<��<�D�<���<���<�M�<E��<���<K�<䝄</��<z�z<M(s<o�k<1qd<]<H�U<igN<�G<��?<r8<�&1<4�)<�"<�]<w$<��<"�<�7�;,��;r��;���;ܐ�;���;|��;|ǚ;� �;l�~;1gc;o]H;׃-;��;��:�N�:C=�:K:):�Å9%
����jj�&n��$׺h��M|�
3�QQJ�%Qa��x��;���N���<����������(���ǻ2�ѻ��ۻ$�廃}�&"���Q��D�
��,����&��r�:� �F�$��-)��N-��a1��f5�1_9��J=��)A���D���H�	�L��2P��S��wW�>[�ە^�}b���e��i��jl���o�W's�({v�X�y�e}�9(���Ł�a��p���}���<#��ɴ��HD���ь��]��l珼�o�������{������c������?�������������d|��y����s���2i��,㧼�\��֪�O��ȭ��@������82������#�����s��*���:
�����������  �  �N=�M=�M=�HL=��K=��J=�	J=,II=�H=7�G=�G=�@F=}E=��D=\�C=W-C=afB=��A=��@=@=4A?=Bu>=2�==��<=P
<=o9;='g:=r�9=0�8=i�7=�7=�46=�X5=�z4=9�3=p�2=��1=��0=90=�/=o/.=�?-=}M,=�X+=�`*=�e)= h(=Fg'=/c&=�[%=�P$=�B#=�0"=!=� =\�=�=ĝ=Dt=�F=�=L�=��=Xd=� =O�=w�=�9=��=�=�)=��
=]	=��=$~=�==�=3=Պ =y�<���<D��<���<Px�<lA�<#�<���<pq�<v�< ��<�e�<  �<���<$�<(��<>3�<���<�/�<W��<��<抷<W��<l`�<�Ƭ<�)�<W��<��<�D�<���<���<�M�<:��<���<K�<ܝ�<1��<Y�z<B(s<Q�k<$qd<�]<J�U<cgN<�G<��?<r8<�&1<4�)<'�"<�]<n$<��<�<�7�;/��;\��;���;��;搶;s��;�ǚ;� �;t�~;gc;�]H;.�-;��;���:�N�:4=�:�:):Zƅ9�
����vhj��n���#׺����|�`
3��QJ�[Qa�	x��;���N���<�����ȩ���(���ǻ�ѻ��ۻ��_}�!"���Q��F�
��,�t����r�� �H�$��-)��N-��a1��f5�%_9��J=��)A���D���H���L��2P��S�owW�_[�˕^��b���e��i�
kl���o�d's�{v�x�y�K}�@(���Ł��`��s���}���@#������ID���ь��]��m珼�o�������{������S������B�������������f|��o����s���)i��/㧼�\��֪�O��ȭ��@������H2�����$�� ������)���<
�����������  �  �N=�M=�M=�HL=��K=��J=�	J=.II=��H==�G=�G=�@F=}E=��D=X�C=O-C=gfB=��A=��@=@=1A?=Du>=,�==��<=S
<=q9;='g:=m�9=1�8=d�7=�7=�46=�X5=�z4==�3=w�2=��1=��0=80=�/=n/.=�?-={M,=yX+=�`*=�e)=%h(=Eg'=)c&=�[%=�P$=�B#=�0"=!=� =W�=�=��=It=�F=�=K�=��=Td=� =T�=v�=�9=��=�=�)=��
=]	=��=#~=�=D�=6=׊ =w�<���<J��<���<Rx�<eA�< �<���<tq�<��<��<�e�<���<�<$�<#��<I3�<���<�/�<G��<�<튷<Q��<w`�<~Ƭ<�)�<G��<��<�D�<���<���<�M�<:��<���<K�<❄</��<c�z<K(s<q�k<0qd<�]<@�U<igN<�G<��?<r8<�&1<?�)<.�"<�]<�$<��<%�<�7�;a��;K��;��;?��;���;R��;�ǚ;� �;g�~;gc;�]H;��-;��;���:}O�:�=�:);):Zƅ9�
�����ij��n���#׺����|�
3�AQJ�5Qa� 	x��;���N���<�����֩���(���ǻ�ѻ��ۻ#�廏}�"���Q��Q�
��,�{��-��r� � �5�$��-)��N-��a1��f5�4_9��J=��)A���D���H��L��2P��S�rwW�I[�˕^��b���e��i��jl���o�h's�{v�j�y�Z}�=(���Ł��`��l���z���2#��˴��HD���ь�{]��l珼�o��w����{������d������;������ �������b|��~����s���(i��'㧼�\��֪�O��ȭ��@������D2������#��������.���9
�����������  �  $�N=	�M=�M=�HL=��K=��J=�	J=4II=��H=>�G=�G=�@F=}E=��D=k�C=P-C=ifB=��A=��@=	@=-A?=Ju>=(�==��<=K
<=l9;='g:=n�9=3�8=^�7=�7=�46=�X5=�z4=6�3=p�2=��1=��0=50=�/=j/.=�?-=�M,=yX+=�`*=�e)=!h(=Eg'=,c&=�[%=�P$=�B#=�0"=!=� =a�=�=��=Lt=�F=�=H�=��=Yd=� =R�=m�=�9=��=�=�)=��
=]	=��="~=�==�=/=׊ =s�<���<V��<���<Sx�<iA�<�<���<cq�<��<��<�e�<���<Ĕ�<$�<#��<R3�<���<�/�<R��<��<���<S��<x`�<nƬ<�)�<H��<��<�D�<���<���<�M�<L��<���<K�<杄<)��<f�z<.(s<Q�k<qd<�]<4�U<ngN<�G<��?<$r8<�&1<G�)<�"<�]<�$<��<>�<�7�;f��;S��;��;0��;���;�;�ǚ;� �;c�~;Kgc;�]H;��-;M�;z��:oO�:�<�::):sƅ9�
����	kj��m���#׺����|��
3��QJ��Qa�	x��;���N���<����������(��ǻS�ѻ��ۻ#��z}��!���Q��H�
��,������r�*� �'�$��-)�xN-��a1��f5�#_9��J=��)A��D�}�H��L��2P��S��wW�5[�ڕ^��b�̐e��i�kl���o�n's�%{v�Q�y�x}�<(���Ł��`��q�������4#��Ѵ��;D���ь�y]��h珼�o��n����{������Y������8������ �������U|��~����s���9i�� 㧼�\�� ֪�&O��ȭ��@������B2�����$��)���|��4���7
�����������  �  �N=�M=�M=�HL=��K=��J=�	J=.II=��H==�G=�G=�@F=}E=��D=X�C=O-C=gfB=��A=��@=@=1A?=Du>=,�==��<=S
<=q9;='g:=m�9=1�8=d�7=�7=�46=�X5=�z4==�3=w�2=��1=��0=80=�/=n/.=�?-={M,=yX+=�`*=�e)=%h(=Eg'=)c&=�[%=�P$=�B#=�0"=!=� =W�=�=��=It=�F=�=K�=��=Td=� =T�=v�=�9=��=�=�)=��
=]	=��=#~=�=D�=6=׊ =w�<���<J��<���<Sx�<eA�< �<���<tq�<��<��<�e�<���<�<$�<#��<I3�<���<�/�<G��<�<튷<Q��<w`�<~Ƭ<�)�<G��<��<�D�<���<���<�M�<:��<���<K�<❄</��<c�z<K(s<q�k<0qd<�]<@�U<jgN<�G<��?<r8<�&1<@�)<.�"<�]<�$<��<%�<�7�;b��;L��;��;?��;���;R��;�ǚ;� �;f�~;gc;�]H;��-;��;���:zO�:�=�:#;):Oƅ9�
�����ij��n���#׺����|�
3�CQJ�7Qa�	x��;���N���<�����֩���(���ǻ�ѻ��ۻ#�廏}�"���Q��Q�
��,�{��-��r� � �5�$��-)��N-��a1��f5�4_9��J=��)A���D���H��L��2P��S�rwW�I[�˕^��b���e��i��jl���o�h's�{v�j�y�Z}�=(���Ł��`��l���z���2#��˴��HD���ь�{]��l珼�o��w����{������d������;������ �������b|��~����s���(i��'㧼�\��֪�O��ȭ��@������D2������#��������.���9
�����������  �  �N=�M=�M=�HL=��K=��J=�	J=,II=�H=7�G=�G=�@F=}E=��D=\�C=W-C=afB=��A=��@=@=4A?=Bu>=2�==��<=P
<=o9;='g:=r�9=0�8=i�7=�7=�46=�X5=�z4=9�3=p�2=��1=��0=90=�/=o/.=�?-=}M,=�X+=�`*=�e)= h(=Fg'=/c&=�[%=�P$=�B#=�0"=!=� =\�=�=ĝ=Dt=�F=�=L�=��=Xd=� =O�=w�=�9=��=�=�)=��
=]	=��=$~=�==�=3=Պ =y�<���<D��<���<Px�<mA�<#�<���<qq�<v�< ��<�e�<  �<���<$�<(��<>3�<���<�/�<W��<��<抷<W��<l`�<�Ƭ<�)�<W��<��<�D�<���<���<�M�<:��<���<K�<ܝ�<1��<Y�z<B(s<Q�k<$qd<�]<J�U<cgN<�G<��?<r8<�&1<4�)<'�"<�]<n$<��<�<�7�;0��;]��;���;��;搶;s��;�ǚ;� �;s�~;gc;�]H;,�-;��;���:�N�:/=�:�:):Eƅ9�
�����hj�o���#׺����|�c
3��QJ�]Qa�	x��;���N���<�����ɩ���(���ǻ�ѻ��ۻ��_}�""���Q��F�
��,�t����r�� �H�$��-)��N-��a1��f5�%_9��J=��)A���D���H���L��2P��S�owW�_[�˕^��b�e��i�
kl���o�d's�{v�x�y�K}�@(���Ł��`��s���}���@#������ID���ь��]��m珼�o�������{������S������B�������������f|��o����s���)i��/㧼�\��֪�O��ȭ��@������H2�����$�� ������)���<
�����������  �  #�N=�M=�M=�HL=��K=��J=�	J=-II=��H=7�G=�G=�@F=
}E=��D=]�C=L-C=afB=��A=��@=@=/A?=Cu>=-�==��<=Q
<=n9;="g:=q�9=4�8=b�7=�7=�46=�X5={4==�3=w�2=��1=��0=60=�/=k/.=�?-=�M,={X+=�`*=�e)=#h(=Eg'=+c&=�[%=�P$=�B#=�0"=!=� =Y�=�=��=Et=�F=�=F�=��=Vd=� =R�=s�=�9=��=�=�)=��
=]	=��=)~=�=D�=9=݊ =��<���<U��<���<Xx�<oA�<�<���<qq�<{�<��<�e�<���<���<$�<(��<@3�<���<�/�<H��<��<銷<Z��<k`�<sƬ<�)�<K��<��<�D�<���<���<�M�<E��<���<K�<䝄</��<z�z<M(s<o�k<1qd<]<H�U<igN<�G<��?<r8<�&1<4�)<�"<�]<w$<��<"�<�7�;,��;r��;���;ܐ�;���;{��;|ǚ;� �;k�~;/gc;l]H;Ճ-;��;��:�N�:<=�:<:):tÅ9a
� �� jj�.n��!$׺l��P|�
3�TQJ�(Qa��x��;���N���<����������(���ǻ2�ѻ��ۻ$�廄}�'"���Q��E�
��,����&��r�:� �F�$��-)��N-��a1��f5�1_9��J=��)A���D���H�	�L��2P��S��wW�>[�ە^�}b���e��i��jl���o�W's�({v�X�y�e}�9(���Ł�a��p���}���<#��ɴ��HD���ь��]��l珼�o�������{������c������?�������������d|��y����s���2i��,㧼�\��֪�O��ȭ��@������82������#�����s��*���:
�����������  �  "�N=�M=�M=�HL=��K=��J=�	J=/II=��H=;�G=�G=�@F=}E=��D=\�C=J-C=gfB=��A=��@=@=2A?=Du>='�==��<=Q
<=r9;=)g:=m�9=6�8=`�7=�7=�46=�X5= {4=8�3=y�2=��1=��0=90=�/=n/.=�?-=M,=yX+=�`*=�e)=(h(=Bg'=%c&=�[%=�P$=�B#=�0"=!=� =Y�=�=��=It=�F=�=I�=��=Rd=� =Y�=r�=�9=��=�=�)=��
=]	=��=.~=�=D�=5=ۊ =��<���<a��<���<^x�<hA�<#�<ɽ�<qq�<��<��<�e�<���<���<
$�<��<L3�<���<�/�<B��<��<銷<F��<t`�<zƬ<�)�<>��<��<�D�<���< ��<�M�<E��<���<!K�<�<2��<��z<@(s<��k<"qd<]<M�U<�gN<�G<��?<r8<�&1<V�)<!�"<�]<|$<��<)�<�7�;L��;&��;��;(��;|��;p��;hǚ;� �;�~;�fc;�]H;�-;��;!��:3O�:*=�:;):�ƅ9+
����jj��m���#׺6��l|�r
3�<QJ�UQa��x��;��xN���<����������(����ǻ9�ѻ��ۻ=�廵}�"���Q��l�
��,����(��r�,� �8�$��-)��N-��a1��f5�A_9��J=��)A���D�m�H��L��2P��S�{wW� [�ϕ^�kb���e��i�kl���o�D's�{v�B�y�k}�4(���Ł��`��g������1#��մ��ID���ь��]��s珼�o��u����{������h������>�������������^|�������s���0i��㧼�\��֪� O���ǭ��@������32������#��"���p��(���.
�����������  �  !�N=�M=�M=�HL=��K=��J=�	J=)II=��H=5�G=�G=�@F=}E=��D=W�C=L-C=_fB=��A=��@=�@=0A?=Au>=/�==��<=O
<=l9;=-g:=p�9=5�8=l�7=�7=�46=�X5={4=?�3=z�2=��1=��0=<0=�/=v/.=�?-=M,=�X+=�`*=�e)="h(=Cg'=+c&=�[%=�P$=�B#=�0"=!=� =Q�=�=��=At=�F=�=G�=��=Wd=� =T�=t�=�9=��=�=�)=��
=]	=��=.~=�=H�=<=� =��<��<Z��<ʧ�<^x�<kA�<3�<���<pq�<�<��<�e�<���<���<$�<��<;3�<���<�/�<<��<��<���<H��<g`�<uƬ<�)�<P��<��<�D�<���<���<�M�<B��<���<'K�<을<4��<��z<\(s<�k<=qd<]<N�U<gN<�G<�?<r8<�&1<H�)<�"<�]<u$<��<�<�7�;��;+��;΢�; ��;p��;F��;pǚ;� �;��~;�fc;7]H;΃-;��;��:�N�:�<�:�9):[ȅ9�
����	hj�n��h#׺J��J|�
3�&QJ��Pa��x��;���N��x<����������(����ǻ,�ѻ��ۻ3�廅}�;"���Q�&�_�
��,����G�s�/� �W�$��-)��N-��a1��f5�0_9��J=��)A���D���H��L��2P��S�VwW�8[���^�pb���e��i��jl���o�I's�{v�R�y�=}�5(���Ł��`��v�������9#��Ǵ��KD���ь��]��w珼�o�������{������o������G�������������k|��u����s���1i��&㧼�\��	֪�O���ǭ��@������22������#�����n��'���/
�����������  �  �N=�M=�M=�HL=��K=��J=�	J=#II=��H=0�G=�G=�@F=
}E=��D=R�C=K-C=ZfB=��A=��@=�@=/A?=9u>=0�==��<=X
<=m9;=)g:=r�9=/�8=l�7=�7=�46=�X5={4=C�3=x�2=��1=��0=C0=�/=v/.=�?-=|M,=�X+=�`*=�e)=h(=Dg'='c&=�[%=�P$=�B#=�0"=!=� =Q�=
�=��=;t=�F=�=J�=��=Rd=� =N�=|�=�9=��=�=�)=��
=]	=��=+~=�=H�=?=� =��<��<X��<̧�<Wx�<qA�</�<���<�q�<o�<��<qe�<���<���<�#�< ��<03�<���<�/�<>��<��<׊�<J��<Y`�<{Ƭ<�)�<K��<z�<�D�<���<���<�M�<:��<���<#K�<�<@��<��z<u(s<v�k<Uqd<]<b�U<�gN<�G<�?<	r8<�&1<9�)<4�"<�]<`$<��<��<�7�;���;.��;���;ِ�;n��;��;gǚ;y �;�~;�fc;"]H;��-;�;&��:�M�:�=�:�9):ƅ9s
�u��	hj�}n���"׺O��&|��	3�KQJ��Pa��x��;���N��~<�����ک���(���ǻ�ѻ�ۻ.�廨}�n"���Q�F�[�
��,����I�s�7� �r�$��-)��N-��a1�g5�E_9��J=��)A���D���H��L��2P�	�S�TwW�9[���^�}b���e��i��jl���o�O's��zv�Z�y�<}�=(���Ł��`��x���n���J#��ƴ��ZD���ь��]���珼�o�������{������n������P�������������z|��z����s���#i��.㧼�\��֪�O���ǭ��@��u���52�������#��	���o�����(
�����������  �  #�N=�M=�M=�HL=��K=��J=�	J=(II=��H=3�G=�G=�@F=
}E=��D=T�C=D-C=\fB=��A=��@= @=.A?==u>=.�==��<=Q
<=l9;=+g:=v�9=7�8=i�7=�7=�46=�X5=	{4=B�3=|�2=��1=��0=A0=�/=s/.=�?-=�M,=�X+=�`*=�e)= h(=Fg'=%c&=�[%=�P$=�B#=�0"=
!=� =P�=
�=��=?t=�F=�=J�=��=Rd=� =P�=u�=�9=��=�=�)=��
=]	=��=2~=�=L�=?=� =��<��<i��<ǧ�<fx�<zA�</�<���<vq�<w�<��<ye�<���<���<�#�<��<53�<���<�/�<4��<��<Պ�<B��<_`�<zƬ<�)�<D��<��<�D�<���<���<�M�<H��<���<&K�<���<C��<��z<w(s<��k<Vqd<.]<m�U<�gN<�G<	�?<!r8<�&1<Q�)<�"<�]<o$<��<
�<�7�;��;��;���;ѐ�;?��;%��;0ǚ;� �;u�~;Rfc;9]H;��-;L�;���:N�:�<�:M9):�ƅ9u
�����hj��m��	#׺���{��	3�QJ��Pa�px��;��{N���<����������(��͂ǻ;�ѻ�ۻ �建}�U"���Q�@�t�
��,����N�s�J� �d�$��-)��N-��a1�g5�F_9��J=��)A���D�}�H��L��2P���S�`wW�[���^�cb���e��i��jl���o�9's��zv�9�y�G}�/(���Ł��`��r���}���D#��ƴ��SD���ь��]���珼�o�������{������w������R�������������o|�������s���3i�� 㧼�\��֪�O���ǭ��@��r���-2�������#��	���f�����(
�����������  �  (�N=�M=�M=�HL=��K=��J=�	J=)II=�H=4�G=�G=�@F=	}E=��D=T�C=>-C=]fB=��A=��@=�@='A?=>u>=%�==��<=P
<=q9;=-g:=m�9==�8=l�7=�7=�46=�X5={4=G�3=��2=��1=��0=?0=�/=w/.=�?-=�M,=|X+=�`*=�e)=(h(=?g'=%c&=�[%=�P$=�B#=�0"=!=� =K�=�=��=@t=�F=�=@�=��=Sd=� =Z�=t�= :=��=�=�)=��
=#]	=��=;~=�=T�=F=� =��<��<u��<ͧ�<rx�<mA�<0�<ͽ�<sq�<��<��<|e�<���<���<$�<��<73�<���<�/�<'��<��<֊�<=��<d`�<aƬ<�)�<=��<~�<�D�<���<��<�M�<P��<���<1K�<���<F��<��z<t(s<��k<Wqd<F]<y�U<�gN<G<�?<9r8<�&1<[�)<#�"<�]<x$<��<�<s7�;��;��;���;ǐ�;��;$��;�ƚ;� �;Y�~;�fc;�\H;%�-;R�;���:�N�:�<�:]:):Vǅ9p
�E���hj��l��`#׺����{��	3��PJ��Pa��x��;��eN��z<��~�������(����ǻ;�ѻ��ۻ`�建}�W"���Q�/���
��,����e�"s�d� �`�$��-)��N-��a1�
g5�D_9��J=��)A���D�j�H���L��2P���S�VwW�[���^�Cb���e��i��jl���o�#'s�	{v�%�y�?}�%(���Ł��`��f�������3#��ش��QD���ь��]��x珼�o�������{�������������R�������������m|�������s���/i��㧼�\���ժ�
O���ǭ��@��o���2�������#��	���Z�����)
�����������  �  '�N=�M=�M=�HL=��K=��J=�	J=(II=��H=.�G=�G=�@F=}E=��D=P�C=A-C=ZfB=��A=��@=�@=*A?=?u>=(�==��<=P
<=n9;=-g:=t�9=:�8=h�7=�7=�46=�X5={4=I�3=��2=��1=��0=G0=�/=v/.=�?-=�M,=�X+=�`*=�e)=#h(=:g'=)c&=�[%=�P$=�B#=�0"=!=� =O�=�=��=;t=�F=�=@�=��=Vd=� =T�=v�=�9=��= �=�)=��
=$]	=��=8~=�=T�=H=� =��<#��<o��<ǧ�<nx�<{A�<4�<Ž�<tq�<z�<��<e�<���<���<�#�<	��<23�<���</�<0��<��<ϊ�<4��<Z`�<hƬ<�)�<E��<o�<�D�<���<���<�M�<N��<���<,K�<��<P��<��z<(s<��k<gqd<!]<��U<�gN<�G<�?<4r8<�&1<S�)<$�"<�]<V$<��<�<�7�;���;���;���;���;&��;���;ǚ;i �;7�~;fc;�\H;L�-;T�;��:�M�:�<�:w9):Sǅ9�
���zij�~m��"׺˨�^|��	3��PJ��Pa�=x�|;��SN���<����������(��ۂǻ2�ѻ��ۻ��廝}�j"���Q�H���
��,����W�s�Y� �u�$��-)��N-��a1�g5�8_9��J=��)A���D���H��L��2P���S�]wW�[���^�Rb���e��i��jl���o�%'s��zv�3�y�L}�*(���Ł��`��o�������B#��մ��OD���ь��]���珼�o�������{������{������X�������������q|������s���/i�� 㧼�\���ժ�O���ǭ��@��e���-2�������#�����m�����
�����������  �  &�N=�M=�M=�HL=��K=��J=�	J="II=��H=*�G=�G=�@F=�|E=��D=I�C=>-C=RfB=��A=��@=�@=+A?=:u>=/�==��<=U
<=k9;=+g:=z�9=9�8=p�7=�7=�46=�X5={4=P�3=��2=��1=��0=H0=�/=x/.=�?-=�M,=�X+=�`*=�e)=!h(=Ag'=(c&=�[%=�P$=�B#=�0"=!=� =I�=�=��=7t=�F=�=E�=��=Sd=� =Q�=z�=�9=��=#�=�)=��
=$]	=��=7~==V�=M=� =��<"��<p��<ا�<nx�<�A�<5�<���<�q�<r�<��<we�<���<���<�#�<��<$3�<���<r/�<(��<��<͊�<9��<M`�<sƬ<�)�<H��<x�<�D�<���<���<�M�<L��<���<.K�< ��<P��<��z<�(s<��k<�qd<6]<��U<�gN<�G<#�?</r8<�&1<K�)<�"<�]<\$<��<��<�7�;���;���;���;n��;��;š�;�ƚ;' �;J�~;�ec;�\H;X�-;��;���:_M�:L=�:�8):=ƅ9�
�^���gj��m��L"׺���{� 	3��PJ��Oa�Zx�{;��[N��r<��n�������(����ǻ,�ѻ�ۻQ�廪}ﻄ"���Q�i�z�
��,�Ω�l�3s�n� ���$��-)��N-��a1�g5�E_9��J=��)A���D���H�݀L��2P���S�KwW�[���^�Vb�e�e��i��jl�{�o�('s��zv�2�y�-}�*(���Ł��`��u���t���J#��Ǵ��XD���ь��]���珼�o�������{������������Z������*�������z|��|����s���3i��#㧼�\�� ֪�O���ǭ��@��f���)2��᪳��#���c�����
�����������  �  (�N=�M=�M=�HL=��K=��J=�	J=#II=�H=,�G=�G=�@F=}E=��D=Q�C=@-C=TfB=��A=��@=�@='A?=:u>=&�==��<=V
<=p9;=-g:=r�9=<�8=n�7=�7=�46=�X5={4=H�3=��2=��1=��0=E0=�/=z/.=�?-=�M,=�X+=�`*=�e)=$h(=>g'=$c&=�[%=�P$=�B#=�0"=!=� =M�=�=��=7t=�F=�=D�=��=Qd=� =U�=y�=�9=��=!�=�)=��
=']	=��=<~==S�=G=� =��<��<z��<ԧ�<rx�<yA�<6�<ʽ�<�q�<{�<��<ue�<���<���<�#�<��<&3�<���<�/�<0��<��<Ɋ�<8��<S`�<jƬ<�)�<<��<y�<�D�<���<��<�M�<Q��<���<9K�<���<Q��<��z<�(s<��k<kqd<L]<��U<�gN<G<�?<6r8<�&1<`�)<$�"<�]<d$<��<��<�7�;���;���;n��;���;#��;��;ǚ;6 �;B�~;�ec;�\H;�-;��;���:�M�:^=�:�9):Kǅ9�
����'hj��l���"׺����{��	3��PJ�mPa�x��;��TN��`<����������(����ǻ$�ѻ��ۻd���}�x"���Q�Y��
��,�Ʃ�]�s�h� ���$��-)��N-��a1�g5�N_9��J=��)A���D�w�H��L��2P���S�HwW�[���^�Cb�y�e��i��jl�}�o�'s��zv��y�4}�'(���Ł��`��k���s���B#��ٴ��ZD���ь��]���珼�o�������{������{������^������$�������w|�������s���-i��㧼�\���ժ�	O���ǭ��@��e���2��𪳼�#������W�����"
�����������  �  ��N=o�M=�M=|NL=�K=��J=uJ={QI=��H=��G=FG=�KF=�E=I�D=� D=�;C=�uB=��A=��@=�@=�S?=�>=ּ==��<=� <=-Q;=�:=P�9=@�8=�8=C,7==S6={x5=��4=`�3=��2=@�1=�1=z.0=.E/=\Y.=k-=!z,=l�+=��*=��)=�(=��'=��&=��%=�$= {#=Aj"=�U!=�= =G!=	=��=&�=E�=V=n =H�=��=Sd=b=��=j~=K(=�=�m=�	=��	=�2=��=�I=9�=CN=�� =w��<�h�<�F�<C�<@��<]��< o�<�&�<��<ـ�<$�<��<�W�<;��<�t�<o��<�|�<���<�q�<��<�U�<8·<�*�<^��<��<HR�<F��<�	�<Fb�<���<��<�`�<���<l�<gS�<���<T�<�z<ns<��k<6Wd<��\<�U<H8N<��F<p�?<�-8<�0<��)<5B"<��<8�<^�<|L<<�;e��;��;�|�;n\�;�M�;vQ�;�h�;I��;©{;�W`;�3E;H?*;~;���:81�:<�:`E:uZN94�H�#���z����K�ߺ���j���g7�ֹN���e���|�c}�����������L����o����ɻJ�ӻ�	޻������V��gi���n���9���m��s�G�!�s�%��*��;.�mI2�|I6�<:�">���A�'�E���I��AM���P���T�r'X���[��:_��b��*f�|�i���l�VWp��s���v��Cz��}�]a�����������+������Q��;ቼ�n��w���:���S��ܒ�����}������Ӟ�����m���P��4���[������K
��W��������v��m識�g���ߪ��W��+ϭ��F��>����5��O����$��蜶�������T�����i����  �  �N=n�M=�M=|NL=��K=��J=wJ=�QI=�H=��G=DG=�KF=��E=R�D=� D=�;C=�uB=��A=��@=�@=�S?=��>=׼==��<=!<=(Q;=�:=L�9=2�8=�8=:,7=<S6=�x5=�4=\�3=��2=D�1=�1=�.0=$E/=YY.=k-=z,=l�+=�*=��)=�(=��'=&=��%=�$=�z#=Dj"=�U!=�= =L!==��=�=G�=V=v =T�=��=Sd=b=��=c~=J(=t�=�m=�	=��	=�2=��=�I=/�==N=�� =���<�h�<�F�<J�<)��<P��<o�<�&�<��<Հ�<$�<��<X�<A��<�t�<j��<�|�<���<�q�<��<�U�<(·<�*�<W��<��<YR�<L��<�	�<Qb�<���<��<�`�<���<s�<bS�<���<g�<�z<ws<y�k<3Wd<�\<?�U<;8N<��F<��?<�-8<�0<��)<2B"<��<1�<g�<�L<|<�;T��;��;i|�;R\�;�M�;�Q�;�h�;��;��{;JW`;�3E;,@*;\~;���:�0�:���:GD:�TN94�H�{����z����i�ߺm���� h7���N�R�e�:�|�"}��В��ł���L��d��o����ɻ�ӻ�	޻������V��Ai���d��:���V��s�D�!���%��*��;.�LI2�LI6�<:�">�}�A�
�E���I��AM���P���T�u'X���[��:_��b��*f���i���l�DWp�̬s���v�$Dz�p�}�ta����������,�������Q��9ቼ�n��[���4���\���������r�����������~���P��<���D������F
��Z��������v��z識�g���ߪ��W��/ϭ��F��+����5��K���%��Ꜷ���|���[�����a����  �  �N=y�M=�M=|NL=�K=��J=yJ=wQI=�H=��G=NG=�KF=�E=S�D=� D=�;C=�uB=��A=��@=�@=�S?=�>=ݼ==��<=!<=&Q;=�:=W�9=0�8=�8=6,7==S6=yx5=�4=a�3=��2=H�1=|1=�.0= E/=_Y.=k-=z,=v�+=�*=��)=�(=��'=��&=��%=�$=�z#=Oj"=�U!=�= =J!=	=��=�=R�=V=r =K�=��=Td=]=��=]~=S(=x�=�m=�	=��	=�2=��=�I=1�=AN=�� =o��<�h�<zF�<\�<)��<b��<o�<�&�<"��<̀�<$�<���<X�<<��<�t�<|��<�|�<���<�q�<��<�U�<2·<�*�<V��<��<AR�<L��<�	�<Ob�<¸�<{�<�`�<���<��<cS�<���<c�<�z<�s<��k<EWd<��\<0�U<58N<��F<��?<�-8<5�0<~�)<3B"<��<%�<o�<jL<Z<�;J��;Q��;�|�;h\�;�M�;ZQ�;�h�;%��;(�{;�W`;3E;�?*;�};���:30�:�:�C:=XN9f�H����G�z�����1�ߺ���D���g7�p�N��e��|�}��뒔������L��Y񴻤o����ɻ��ӻ
޻�����W��Qi���4��:���^��s�5�!���%��*��;.�XI2�qI6�-<:��!>���A���E��I��AM���P���T�U'X���[��:_��b��*f���i���l�OWp��s���v�8Dz�K�}�sa����������,����Q��1ቼ�n��h���9���R��Β�����n�������������t���:��=���K������F
��\��������v���識�g���ߪ��W��/ϭ��F��/����5��A��� %������������]�����N����  �  �N=q�M=�M=�NL=�K=��J=|J=�QI=�H=��G=HG=�KF=�E=S�D=� D=�;C=�uB=��A=��@=�@=�S?=�>=߼==��<=!<=+Q;=�:=O�9=1�8=�8=7,7=@S6=wx5=�4=\�3=��2=C�1=}1=.0=#E/=WY.=k-=z,=n�+=�*=��)=�(=��'=Ɨ&=��%=�$={#=Dj"=�U!=�= =N!==��=!�=H�=V=w =S�=��=Wd=\=��=a~=K(=s�=�m=�	=��	=�2=��=�I=*�=;N=�� =k��<�h�<|F�<D�<"��<Q��<o�<�&�<��<΀�<$�<��<X�<F��<�t�<n��<�|�<���<�q�<��<�U�<.·<�*�<c��<��<SR�<U��<�	�<Fb�<˸�<}�<�`�<���<l�<[S�<���<Z�<�z<us<l�k<2Wd<��\<!�U<C8N<|�F<t�?<�-8<�0<z�)<GB"<��<2�<x�<�L<�<�;w��;"��;||�;�\�;�M�;�Q�;�h�;N��;ǩ{;�W`;�3E;;@*;)~;���:�0�:i��:/E:�TN9��H�����z�u���Ĉߺ ��B���g7�̺N�W�e�҄|�8}��ϒ��Ђ��M��f��o����ɻ��ӻ
޻���۶�V��:i�|�`��	:�ܲ�M��s�2�!���%��*��;.�CI2�NI6�<:��!>���A���E��I��AM���P���T�|'X���[��:_��b��*f���i���l�OWp���s���v�1Dz�x�}�ya����������,�������Q��-ቼ�n��Y���.���N��ܒ�����m�������������x���L��0���@������=
��U��������v���識�g���ߪ��W��7ϭ��F��8����5��K���%��霶�������V�����g����  �  �N=o�M=�M=|NL=�K=��J=tJ=�QI=�H=��G=LG= LF=�E=O�D=� D=�;C=�uB=��A=��@=�@=�S?=��>=׼==��<= !<=)Q;=�:=N�9=7�8=�8=7,7=3S6=tx5=ߛ4=X�3=��2==�1=�1=u.0=!E/=XY.=
k-=z,=j�+=�*=��)=�(=��'=��&=��%=�$={#=Gj"=�U!=�= =Q!==��=)�=I�=V=o =S�=��=Sd=a=��=a~=G(=x�=�m=�	=��	=�2=��=�I=*�=8N=�� =g��<�h�<zF�<A�<0��<T��<o�<�&�<��<ۀ�<$�<��<X�<:��<u�<r��<�|�<���<r�<��<�U�<;·<�*�<g��<��<ZR�<H��<�	�<Hb�<���<��<�`�<���<n�<[S�<���<K�<�z<_s<v�k<Wd<��\<�U<8N<��F<w�?<�-8<	�0<~�)<2B"<��<L�<[�<�L<^<�;|��;F��;�|�;�\�;�M�;	R�;�h�;o��;��{;X`;�3E;%@*;d~;���:�1�:F��:�D:TTN9ĜH�����z�h���U�ߺ%��Y��#h7���N���e���|��}��ᒔ�Ȃ���L��3�p����ɻ)�ӻ�	޻�����V��\i�q�S���9���A��s�D�!�b�%��*��;.�cI2�MI6�<:�">�~�A��E��I��AM���P���T�y'X���[��:_��b��*f���i���l�\Wp���s���v�2Dz�z�}�ja����������	,�������Q��<ቼ�n��]���9���G��ؒ�����|�������������k���B��,���O������J
��M��������v��~識�g���ߪ��W��6ϭ��F��G����5��V���%������������h�����e����  �  ߇N=r�M=�M=zNL=�K=��J={J=�QI=�H=��G=QG= LF=�E=W�D=� D=�;C=�uB=��A=��@=�@=�S?=��>=ݼ==��<=!<=&Q;=�:=R�9=*�8=�8=4,7=8S6=wx5=֛4=U�3=��2=6�1=y1=z.0=E/=TY.=k-=z,=n�+=�*=��)=�(=��'=ė&=��%=�$={#=Lj"=�U!=�= =U!==��=(�=L�=V=t =X�=��=Wd=^=��=]~=J(=r�=�m=�	=��	=�2=��=�I=*�=5N=�� =h��<�h�<rF�<7�<��<T��<o�<�&�<��<Ѐ�<$�<��<X�<A��<u�<y��<}�<���<�q�<��<V�<9·<�*�<i��<��<aR�<Q��<�	�<Kb�<���<~�<�`�<���<h�<SS�<���<R�<�z<?s<v�k< Wd<��\<�U<&8N<o�F<p�?<n-8<�0<{�)<-B"<��<=�<t�<�L<t<�;���;u��;�|�;�\�;N�;�Q�;�h�;���;/�{;SX`;�3E;Y@*;�~;���:*1�:���:.D:�WN9��H�����z�������ߺ������Qh7���N�!�e� �|�Z}��璔�₟�M��q��o����ɻ�ӻ�	޻�����tV��Ii�i�A���9�ʲ�0��s�#�!�e�%��*��;.�NI2�8I6�<:��!>���A��E��I��AM���P���T��'X���[��:_�"�b�+f���i���l�~Wp���s���v�>Dz���}��a����������,�������Q��0ቼ�n��W���1���@��В�����h�������������m���8��*���G������B
��P��������v���識�g���ߪ��W��>ϭ��F��?����5��f���%�����%������d�����h����  �  އN=q�M=�M=�NL=�K=��J=}J=�QI=�H=��G=SG=LF=�E=]�D=� D=�;C=�uB=��A=��@=�@=�S?=��>=�==��<=!<=(Q;=�:=O�9=,�8=�8=/,7=3S6=nx5=؛4=S�3=��2=:�1=v1=t.0=E/=RY.=k-=z,=n�+=�*=��)=�(=��'=ŗ&=��%=�$={#=Oj"=�U!=�= =V!==��=)�=Q�=V=y =V�=��=Vd=\=��=Z~=H(=n�=�m=�	=��	=�2=��=�I=!�=0N=�� =V��<�h�<iF�<;�<��<L��<o�<�&�<"��<ɀ�<$�<��<X�<K��<u�<���< }�<���< r�<�<V�<A·<+�<k��<��<[R�<W��<�	�<Ob�<θ�<p�<�`�<���<o�<MS�<���<F�<�z<Ks<Q�k<	Wd<��\<��U<8N<]�F<{�?<i-8<�0<[�)<EB"<��<,�<�<�L<�<�;���;���;�|�;�\�;AN�;R�;8i�;���;��{;TX`;D4E;�@*;�~;-��:�0�:x�:�D:eQN9W�H�u����z�/���)�ߺ{�����`h7��N���e�,�|��}���������M��z��o����ɻ��ӻ
޻�����V��)i�l�2���9����*�{s��!�]�%��*��;.�5I2�>I6�<:��!>���A���E��I��AM� �P���T��'X�ֵ[��:_�4�b��*f�Жi���l�tWp��s���v�NDz���}�~a����������,��鿆��Q��,ቼ�n��P���'���D��ǒ�����Z�������������f���4��(���4������;
��W��������v���識�g���ߪ��W��Dϭ��F��K����5��_���%������"������k�����b����  �  �N=o�M=�M={NL=�K=��J=~J=�QI=�H=��G=WG=
LF=�E=[�D=� D=�;C=�uB=��A=��@=�@=�S?=��>=�==��<= !<='Q;=�:=M�9=/�8=z8=/,7=1S6=jx5=֛4=P�3=��2=4�1=v1=o.0=E/=MY.=k-=z,=k�+=�*=��)=�(=��'=ȗ&=��%=�$=
{#=Tj"=�U!=�= =Z!==��=.�=V�= V=y =T�=��=Wd=]=��=[~=G(=o�=�m=�	=��	=�2=��=�I=�=-N=�� =N��<�h�<iF�<(�<��<H��<o�<�&�<��<Ԁ�<$�<��<X�<O��<u�<���<}�<���<r�<�<V�<R·<
+�<v��<��<ZR�<[��<�	�<Hb�<���<x�<�`�<���<b�<DS�<���<<�<�z</s<I�k<�Vd<��\<�U<8N<P�F<Y�?<z-8<�0<n�)<-B"<��<L�<��<�L<�<�;���;���;
}�;�\�;5N�;RR�;i�;���;�{;�X`;z4E;�@*;�~;Z��:�1�:���:E:�UN9N�H�����z�#���W�ߺ�������h7�;�N�)�e�#�|��}���������M��d��o����ɻ�ӻ
޻���¶�V��0i�\����9�����^s��!�I�%��*�s;.�6I2�AI6��;:��!>���A��E��I��AM���P���T��'X�˵[��:_�9�b�+f�ٖi���l��Wp�"�s���v�JDz���}�wa����������,�������Q��+ቼ�n��T���"���:���������d�������������T���,�����:������8
��H��������v���識�g���ߪ��W��Mϭ��F��U����5��m���%��
���%������n�����s����  �  ��N=h�M=�M=zNL=�K=��J={J=�QI=�H= �G=TG=LF=�E=b�D=� D=�;C=�uB=��A=��@=�@=�S?=�>=ܼ==��<= !<=&Q;=�:=I�9=+�8=u8=.,7=,S6=lx5=Λ4=I�3=��2=*�1=s1=k.0=E/=HY.=�j-=z,=f�+=�*=��)=�(=��'=ɗ&=��%=!�$={#=Oj"=�U!=�= =\!==��=1�=Q�=!V=| =]�=��=Sd=`=��=]~=A(=i�=�m=�	=��	=�2=��=�I=�='N=�� =R��<vh�<cF�<�<��<=��<o�<�&�<
��<׀�<$�<#��<X�<U��<u�<���<}�<���<r�<�<V�<M·<+�<{��<��<uR�<S��<�	�<Nb�<���<��<�`�<���<]�<@S�<���<8�<jz<s<U�k<�Vd<��\<�U<�7N<I�F<M�?<o-8<��0<{�)<*B"<��<J�<u�<�L<�<�;���;���;�|�;-]�;lN�;TR�;bi�;��;��{;�X`;�4E;�@*;k;���:2�:���:�D:�VN9��H�j���z�5����ߺ���Q���h7��N���e�G�|��}�����8���+M����p����ɻ�ӻ�	޻��绸��<V��i�P�.���9�����^s���!�<�%��*�k;.�'I2�I6��;:��!>�x�A��E��I��AM��P�ȏT��'X�ֵ[�;_�:�b�=+f�ܖi���l��Wp��s��v�RDz���}��a����������,�������Q��3ቼ�n��J������9��Ò�����T����������}��Y���4�����5������@
��L��������v��識�g���ߪ��W��Qϭ��F��Y����5��}���%�����1������y�����x����  �  ۇN=p�M=�M={NL=�K=��J=}J=�QI=�H=��G=^G=LF=�E=g�D=� D=�;C=�uB=��A=��@=�@=�S?=��>=�==��<=!<=$Q;=�:=O�9='�8=}8=+,7='S6=ex5=Λ4=I�3=��2=1�1=n1=i.0=E/=OY.=k-=z,=m�+=�*=��)=�(=��'=Ɨ&=��%=!�$={#=\j"=�U!=�= =^!==��=0�=]�=#V={ =V�=��=Vd=`=��=W~=E(=k�=�m=�	=��	=�2=z�=�I=�=$N=�� =?��<lh�<]F�<.�<��<J��<o�<�&�<��<Ӏ�<$�<��<X�<S��<u�<���<}�<���<r�<�<V�<T·<+�<{��<��<gR�<V��<�	�<Sb�<¸�<r�<�`�<���<`�<ES�<z��<1�<[z<&s<1�k<�Vd<��\<͕U<�7N<L�F<[�?<^-8<�0<a�)<.B"<��<H�<��<�L<�<�;���;��;-}�; ]�;�N�;AR�;�i�;���;D�{;Y`;�4E;�@*;;n��:�1�:}�:�D:OTN9ØH�D����z�t���x�ߺ���A���h7�t�N�P�e���|��}��+������M�����o����ɻ�ӻ�	޻���Ѷ�yV��i�L�����9�����^s��!�?�%�~*�d;.�(I2�5I6�<:��!>�v�A��E��I��AM��P�ďT��'X��[�;_�V�b�'+f��i���l��Wp�:�s��v�\Dz���}��a����������,��񿆼�Q��+ቼ�n��P������2���������I����������{��R��������4������=
��K��������v���識�g���ߪ��W��Lϭ��F��`����5��q���'%�����7������������q����  �  ӇN=n�M=�M=�NL=�K=��J=�J=�QI=�H=�G=[G=LF=�E=k�D=� D=�;C=�uB=��A=��@=�@=T?=��>=�==��<=!<=)Q;=�:=J�9=�8=x8=$,7=1S6=ex5=͛4=H�3=��2=1�1=i1=q.0=E/=JY.=�j-=z,=j�+=�*=��)=�(=��'=͗&=��%=,�$={#=\j"=�U!=�= =c!=#=��=/�=_�= V=� =^�=��=]d=Z=��=V~=B(=c�=�m=�	=��	=�2=u�=�I=�=!N=�� =;��<�h�<MF�<!�<���<;��<�n�<�&�<��<̀�<)$�<��<(X�<`��<u�<���<	}�<���<r�<!�<V�<Y·<+�<}��<��<fR�<g��<�	�<Jb�<͸�<l�<�`�<}��<V�<9S�<}��<<�<Iz<%s<��k<�Vd<��\<ݕU<�7N<4�F<F�?<;-8<�0<S�)<CB"<��<N�<��<�L<=�;���;ɭ�;D}�;]�;�N�;tR�;�i�;Д�;��{;�X`;!5E;�A*;�~;t��:�1�: �:�E:2QN9U�H�'����z�J���(�ߺ���U��i7��N�I�e��|��}��>���*���WM�����o����ɻ��ӻ
޻��绔��VV���h�T�����9������Fs��!�A�%�u*�n;.��H2�I6��;:��!>���A���E��I��AM�"�P��T��'X���[��:_�g�b�)+f��i�
�l��Wp�@�s���v�zDz���}��a������Ǖ��,�������Q��ቼ�n��<������8���������?����������{��M���"�����������,
��E��������v���識�g���ߪ��W��Xϭ��F��T����5��q���@%�����?������x�����{����  �  ߇N=k�M=�M=NL=�K=��J=zJ=�QI=�H=�G=[G=LF=�E=f�D=� D=�;C=�uB=��A=��@=�@=�S?=��>=ܼ==��<=!<=+Q;=�:=J�9=*�8={8=$,7=&S6=ax5=ɛ4=G�3=��2=.�1=h1=g.0=E/=LY.= k-=z,=g�+=�*=��)=�(=��'=ŗ&=��%=#�$={#=Yj"=�U!=�= =`!=!=��=9�=\�=#V=| =Y�=��=Td=_=��=[~=?(=j�=�m=�	=}�	=�2=t�=�I=�=!N=�� =4��<jh�<KF�<(�<��<?��<�n�<�&�<��<׀�<$�<��<X�<W��<u�<���<}�<���<r�<�<#V�<g·<+�<���<��<kR�<Q��<�	�<Mb�<ȸ�<u�<�`�<���<a�<=S�<l��<,�<Az<s<&�k<�Vd<��\<ĕU<�7N<<�F<Z�?<j-8<��0<a�)<=B"<��<R�<r�<�L<�<�;
��;Э�;k}�;Q]�;�N�;bR�;�i�;/��;��{;
Y`;5E;A*;#;$��:Y2�:���:^F:nQN9��H�5��6�z�B�����ߺ �����i7���N�v�e���|��}��`������!M��{�p����ɻ��ӻ�	޻���׶�aV��i�B����9������Ns��!��%��*�`;.�"I2�)I6�<:��!>�w�A��E�	�I��AM��P�ƏT��'X��[�;_�l�b�8+f���i��l��Wp�M�s��v�}Dz���}��a������ɕ��,�������Q��/ቼ�n��J������2���������H����������r��?���$�����/������B
��I��������v���識�g���ߪ��W��Sϭ��F��d����5��u���,%�����B������������q����  �  ؇N=i�M=�M=wNL=�K=��J={J=�QI=
�H=	�G=^G=LF=�E=h�D= D=�;C=�uB=��A=��@=�@=�S?=�>=ݼ==��<=� <=&Q;=�:=H�9="�8=p8=),7=%S6=jx5=͛4=@�3=��2=*�1=p1=h.0=E/=HY.=�j-=z,=f�+=�*=��)=#�(=��'=̗&=��%= �$={#=Uj"=�U!=�= =f!=*=��=3�=V�=.V=| =`�=��=Vd=g=��=[~=?(=h�=�m=�	=��	=�2=|�=�I=�=N=�� =F��<fh�<UF�<�<���<;��<�n�<�&�<��<��<$�<0��<X�<\��<'u�<���<}�<���<-r�<�<V�<X·<+�<���<��<�R�<W��<�	�<Tb�<���<|�<�`�<���<E�<>S�<t��<3�<Xz<�s<�k<�Vd<��\<֕U<�7N<C�F<"�?<Q-8<��0<l�)<B"<��<m�<y�<�L<�<�;/��;��;)}�;(]�;�N�;�R�;�i�;
��;�{;jY`;"5E;�@*;�;%��:;3�:���::E:SN96�H�j����z�������ߺ���G��ui7���N���e�y�|��}��;���8����M����p����ɻH�ӻ�	޻��绠��V��i�����9������+s��!�0�%��*�4;.�#I2�I6��;:��!>�V�A�'�E�	�I��AM��P���T��'X��[�;_�I�b�?+f��i��l��Wp�'�s��v�hDz���}��a������ƕ��,������Q��0ቼ�n��I������ ���������O���w������~��N��� �����8��n���<
��<��������v���識�g���ߪ��W��Rϭ��F��]����5������7%��%���:�����������������  �  ߇N=k�M=�M=NL=�K=��J=zJ=�QI=�H=�G=[G=LF=�E=f�D=� D=�;C=�uB=��A=��@=�@=�S?=��>=ܼ==��<=!<=+Q;=�:=J�9=*�8={8=$,7=&S6=ax5=ɛ4=G�3=��2=.�1=h1=g.0=E/=LY.= k-=z,=g�+=�*=��)=�(=��'=ŗ&=��%=#�$={#=Yj"=�U!=�= =`!=!=��=9�=\�=#V=| =Y�=��=Td=_=��=[~=?(=j�=�m=�	=}�	=�2=t�=�I=�="N=�� =4��<kh�<KF�<(�<��<?��<�n�<�&�<��<׀�<$�<��<X�<W��<u�<���<}�<���<r�<�<#V�<g·<+�<���<��<kR�<Q��<�	�<Mb�<Ǹ�<u�<�`�<���<a�<=S�<l��<,�<Az<s<&�k<�Vd<��\<ĕU<�7N<=�F<[�?<j-8<��0<b�)<>B"<��<S�<r�<�L<�<�;
��;Э�;k}�;Q]�;�N�;bR�;�i�;/��;��{;	Y`;5E;A*;!;!��:U2�:���:WF:QQN9��H�<��=�z�E�����ߺ"�����i7���N�w�e���|��}��a������!M��|�p����ɻ��ӻ�	޻���׶�bV��i�B����9������Ns��!��%��*�`;.�"I2�)I6�<:��!>�w�A��E�	�I��AM��P�ƏT��'X��[�;_�l�b�8+f���i��l��Wp�M�s��v�}Dz���}��a������ɕ��,�������Q��/ቼ�n��J������2���������H����������r��?���$�����/������B
��I��������v���識�g���ߪ��W��Sϭ��F��d����5��u���,%�����B������������q����  �  ӇN=n�M=�M=�NL=�K=��J=�J=�QI=�H=�G=[G=LF=�E=k�D=� D=�;C=�uB=��A=��@=�@=T?=��>=�==��<=!<=)Q;=�:=J�9=�8=x8=$,7=1S6=ex5=͛4=H�3=��2=1�1=i1=q.0=E/=JY.=�j-=z,=j�+=�*=��)=�(=��'=͗&=��%=,�$={#=\j"=�U!=�= =c!=#=��=/�=_�= V=� =^�=��=]d=Z=��=V~=B(=c�=�m=�	=��	=�2=u�=�I=�=!N=�� =;��<�h�<MF�<!�<���<<��<�n�<�&�<��<̀�<)$�<��<(X�<`��<u�<���<	}�<���<r�<!�<V�<Y·<+�<}��<��<eR�<g��<�	�<Jb�<͸�<l�<�`�<}��<V�<8S�<}��<<�<Iz<%s<��k<�Vd<��\<ݕU<�7N<4�F<G�?<;-8<�0<S�)<CB"<��<O�<��<�L<=�;���;ʭ�;D}�;]�;�N�;tR�;�i�;Д�;��{;�X`;5E;�A*;�~;n��:�1�:�:�E:�PN9��H�5���z�Q���/�ߺ���X��i7��N�L�e��|��}��?���+���XM�����o����ɻ��ӻ
޻��绕��VV���h�T�����9������Fs��!�A�%�u*�n;.��H2�I6��;:��!>���A���E��I��AM�"�P��T��'X���[��:_�g�b�)+f��i�
�l��Wp�@�s���v�zDz���}��a������Ǖ��,�������Q��ቼ�n��<������8���������?����������{��M���"�����������,
��E��������v���識�g���ߪ��W��Xϭ��F��T����5��q���@%�����?������x�����{����  �  ۇN=p�M=�M={NL=�K=��J=}J=�QI=�H=��G=^G=LF=�E=g�D=� D=�;C=�uB=��A=��@=�@=�S?=��>=�==��<=!<=$Q;=�:=O�9='�8=}8=+,7='S6=ex5=Λ4=I�3=��2=1�1=n1=i.0=E/=OY.=k-=z,=m�+=�*=��)=�(=��'=Ɨ&=��%=!�$={#=\j"=�U!=�= =^!==��=0�=]�=#V={ =V�=��=Vd=`=��=W~=E(=k�=�m=�	=��	=�2=z�=�I=�=%N=�� =?��<mh�<]F�<.�<	��<K��<o�<�&�<��<Ԁ�<$�<��<X�<T��<u�<���<}�<���<r�<�<V�<T·<+�<{��<��<gR�<V��<�	�<Sb�<¸�<q�<�`�<���<`�<ES�<z��<1�<Zz<&s<1�k<�Vd<��\<͕U<�7N<M�F<\�?<^-8<�0<b�)</B"<��<I�<��<�L<�<�;���;��;-}�; ]�;�N�;AR�;�i�;ߔ�;B�{;Y`;�4E;�@*;;f��:�1�:t�:~D:TN9�H�X����z�~�����ߺ���E���h7�x�N�T�e���|��}��,������M�����o����ɻ�ӻ�	޻���Ҷ�zV��i�M�����9�����^s��!�?�%�~*�d;.�(I2�5I6�<:��!>�v�A��E��I��AM��P�ďT��'X��[�;_�V�b�'+f��i���l��Wp�:�s��v�\Dz���}��a����������,��񿆼�Q��+ቼ�n��P������2���������I����������{��R��������4������=
��K��������v���識�g���ߪ��W��Lϭ��F��`����5��q���'%�����7������������q����  �  ��N=h�M=�M=zNL=�K=��J={J=�QI=�H= �G=TG=LF=�E=b�D=� D=�;C=�uB=��A=��@=�@=�S?=�>=ܼ==��<= !<=&Q;=�:=I�9=+�8=u8=.,7=,S6=lx5=Λ4=I�3=��2=*�1=s1=k.0=E/=HY.=�j-=z,=f�+=�*=��)=�(=��'=ɗ&=��%=!�$={#=Oj"=�U!=�= =\!==��=1�=Q�=!V=| =]�=��=Sd=`=��=]~=A(=j�=�m=�	=��	=�2=��=�I=�=(N=�� =S��<wh�<dF�<�<��<>��<o�<�&�<��<׀�<$�<#��<X�<U��<u�<���<}�<���<r�<�<V�<M·<+�<{��<��<tR�<S��<�	�<Mb�<���<��<�`�<���<\�<@S�<���<8�<jz<s<U�k<�Vd<��\<�U<�7N<J�F<M�?<o-8<��0<|�)<+B"<��<J�<u�<�L<�<�;���;���;�|�;-]�;lN�;TR�;ai�;��;��{;�X`;�4E;�@*;f;���:	2�:���:�D:hVN9�H������z�A����ߺ���V���h7�$�N���e�L�|��}�����:���,M����p����ɻ�ӻ�	޻��绹��=V��i�Q�.���9�����^s���!�<�%��*�k;.�'I2�I6��;:��!>�x�A��E��I��AM��P�ȏT��'X�ֵ[�;_�:�b�=+f�ܖi���l��Wp��s��v�RDz���}��a����������,�������Q��3ቼ�n��J������9��Ò�����T����������}��Y���4�����5������@
��L��������v��識�g���ߪ��W��Qϭ��F��Y����5��}���%�����1������y�����x����  �  �N=o�M=�M={NL=�K=��J=~J=�QI=�H=��G=WG=
LF=�E=[�D=� D=�;C=�uB=��A=��@=�@=�S?=��>=�==��<= !<='Q;=�:=M�9=/�8=z8=/,7=1S6=jx5=֛4=P�3=��2=4�1=v1=o.0=E/=MY.=k-=z,=k�+=�*=��)=�(=��'=ȗ&=��%=�$=
{#=Tj"=�U!=�= =Z!==��=.�=V�= V=y =T�=��=Xd=]=��=[~=G(=p�=�m=�	=��	=�2=��=�I=�=-N=�� =O��<�h�<iF�<)�<��<I��<o�<�&�<��<Հ�<$�<��<X�<P��<u�<���<}�<���<r�<�<V�<R·<
+�<u��<��<YR�<Z��<�	�<Hb�<���<w�<�`�<���<a�<CS�<���<<�<z</s<I�k<�Vd<��\<�U<8N<Q�F<Z�?<z-8<�0<o�)<.B"<��<M�<��<�L<�<�;���;���;}�;�\�;5N�;QR�;i�;���;�{;�X`;v4E;�@*;�~;O��:�1�:|��:�D:AUN9��H�����z�0���d�ߺ�������h7�A�N�/�e�(�|��}���������M��f��o����ɻ�ӻ
޻���¶�V��0i�\����9�����^s��!�J�%��*�s;.�6I2�AI6��;:��!>���A��E��I��AM���P���T��'X�˵[��:_�9�b�+f�ٖi���l��Wp�"�s���v�JDz���}�wa����������,�������Q��+ቼ�n��T���"���:���������d�������������T���,�����:������8
��H��������v���識�g���ߪ��W��Mϭ��F��U����5��m���%��
���%������n�����s����  �  އN=q�M=�M=�NL=�K=��J=}J=�QI=�H=��G=SG=LF=�E=]�D=� D=�;C=�uB=��A=��@=�@=�S?=��>=�==��<=!<=(Q;=�:=O�9=,�8=�8=/,7=3S6=nx5=؛4=S�3=��2=:�1=v1=t.0=E/=RY.=k-=z,=n�+=�*=��)=�(=��'=ŗ&=��%=�$={#=Oj"=�U!=�= =V!==��=*�=Q�=V=y =V�=��=Vd=\=��=Z~=H(=n�=�m=�	=��	=�2=��=�I=!�=0N=�� =V��<�h�<jF�<<�<��<M��<o�<�&�<#��<ɀ�<$�<��<X�<K��<u�<���< }�<���< r�<�<V�<A·<+�<k��<��<[R�<W��<�	�<Ob�<͸�<o�<�`�<���<n�<MS�<���<E�<�z<Ks<Q�k<	Wd<��\<��U<8N<]�F<|�?<j-8<�0<\�)<FB"<��<-�<��<�L<�<�;���;���;�|�;�\�;AN�;R�;7i�;���;��{;QX`;@4E;�@*;|~;!��:�0�:k�:�D:�PN9ǚH����éz�=���6�ߺ������fh7�$�N���e�1�|��}�����򂟻M��|��o����ɻ��ӻ

޻�����V��)i�l�2���9����*�{s��!�]�%��*��;.�6I2�>I6�<:��!>���A���E��I��AM� �P���T��'X�ֵ[��:_�4�b��*f�Жi���l�tWp��s���v�NDz���}�~a����������,��鿆��Q��,ቼ�n��P���'���D��ǒ�����Z�������������f���4��(���4������;
��W��������v���識�g���ߪ��W��Dϭ��F��K����5��_���%������"������k�����b����  �  ߇N=r�M=�M=zNL=�K=��J={J=�QI=�H=��G=QG= LF=�E=W�D=� D=�;C=�uB=��A=��@=�@=�S?=��>=ݼ==��<=!<=&Q;=�:=R�9=*�8=�8=4,7=8S6=wx5=֛4=U�3=��2=6�1=y1=z.0=E/=TY.=k-=z,=n�+=�*=��)=�(=��'=ŗ&=��%=�$={#=Lj"=�U!=�= =U!==��=(�=L�=V=t =X�=��=Wd=^=��=]~=J(=r�=�m=�	=��	=�2=��=�I=*�=5N=�� =i��<�h�<sF�<7�<��<U��<o�<�&�<��<р�<$�<��<X�<B��<u�<y��<}�<���<�q�<��<V�<9·<�*�<i��<��<aR�<P��<�	�<Jb�<���<~�<�`�<���<h�<SS�<���<R�<�z<?s<v�k< Wd<��\<�U<&8N<o�F<q�?<o-8<�0<|�)<.B"<��<>�<u�<�L<v<�;���;v��;�|�;�\�;N�;�Q�;�h�;���;-�{;PX`;�3E;U@*;�~;���:1�:���:D:iWN9�H� ��˪z�������ߺ������Wh7���N�'�e��|�]}��钔�䂟�M��r��o����ɻ�ӻ�	޻�����uV��Ji�i�A���9�ʲ�1��s�#�!�f�%��*��;.�NI2�8I6�<:��!>���A��E��I��AM���P���T��'X���[��:_�"�b�+f���i���l�~Wp���s���v�>Dz���}��a����������,�������Q��0ቼ�n��W���1���@��В�����h�������������m���8��*���G������B
��P��������v���識�g���ߪ��W��>ϭ��F��?����5��f���%�����%������d�����h����  �  �N=o�M=�M=|NL=�K=��J=tJ=�QI=�H=��G=LG= LF=�E=O�D=� D=�;C=�uB=��A=��@=�@=�S?=��>=׼==��<= !<=)Q;=�:=N�9=7�8=�8=7,7=3S6=tx5=ߛ4=X�3=��2==�1=�1=u.0=!E/=XY.=
k-=z,=j�+=�*=��)=�(=��'=��&=��%=�$={#=Gj"=�U!=�= =Q!==��=)�=I�=V=o =S�=��=Sd=a=��=a~=G(=x�=�m=�	=��	=�2=��=�I=*�=8N=�� =h��<�h�<{F�<B�<0��<U��<o�<�&�<��<ۀ�<$�<��<X�<:��<u�<r��<�|�<���<r�<��<�U�<;·<�*�<g��<��<YR�<G��<�	�<Gb�<���<��<�`�<���<m�<[S�<���<K�<�z<_s<v�k<Wd<��\<�U<8N<��F<x�?<�-8<
�0<�)<3B"<��<M�<\�<�L<`<�;}��;F��;�|�;�\�;�M�;	R�;�h�;n��;��{;X`;�3E;!@*;`~;���:�1�:;��:�D:�SN9&�H���7�z�u���a�ߺ+��^��(h7���N���e���|��}��㒔�ɂ���L��5�p����ɻ*�ӻ�	޻�����V��\i�q�S���9���A��s�D�!�c�%��*��;.�dI2�MI6�<:�">�~�A��E��I��AM���P���T�y'X���[��:_��b��*f���i���l�\Wp���s���v�2Dz�z�}�ja����������	,�������Q��<ቼ�n��]���9���G��ؒ�����|�������������k���B��,���O������J
��M��������v��~識�g���ߪ��W��6ϭ��F��G����5��V���%������������h�����e����  �  �N=q�M=�M=�NL=�K=��J=|J=�QI=�H=��G=HG=�KF=�E=S�D=� D=�;C=�uB=��A=��@=�@=�S?=�>=߼==��<=!<=+Q;=�:=O�9=1�8=�8=7,7=@S6=wx5=�4=\�3=��2=C�1=}1=.0=#E/=WY.=k-=z,=n�+=�*=��)=�(=��'=Ɨ&=��%=�$={#=Dj"=�U!=�= =N!==��=!�=H�=V=w =S�=��=Wd=]=��=a~=K(=s�=�m=�	=��	=�2=��=�I=*�=<N=�� =l��<�h�<|F�<D�<"��<R��<o�<�&�<��<΀�<$�<��<X�<F��<�t�<n��<�|�<���<�q�<��<�U�<.·<�*�<c��<��<RR�<U��<�	�<Fb�<˸�<}�<�`�<���<l�<ZS�<���<Z�<�z<us<l�k<2Wd<��\<"�U<C8N<|�F<t�?<�-8<�0<{�)<HB"<��<3�<y�<�L<�<�;x��;"��;}|�;�\�;�M�;�Q�;�h�;M��;ũ{;�W`;�3E;7@*;&~;���:�0�:`��:E:|TN9��H����!�z����Έߺ��F���g7�кN�[�e�ք|�9}��ђ��т��M��h��o����ɻ��ӻ
޻���۶�V��:i�}�`��	:�ܲ�M��s�2�!���%��*��;.�CI2�NI6�<:��!>���A���E��I��AM���P���T�|'X���[��:_��b��*f���i���l�NWp���s���v�1Dz�x�}�ya����������,�������Q��-ቼ�n��Y���.���N��ܒ�����m�������������x���L��0���@������=
��U��������v���識�g���ߪ��W��7ϭ��F��8����5��K���%��霶�������V�����g����  �  �N=y�M=�M=|NL=�K=��J=yJ=wQI=�H=��G=NG=�KF=�E=S�D=� D=�;C=�uB=��A=��@=�@=�S?=�>=ݼ==��<=!<=&Q;=�:=W�9=0�8=�8=6,7==S6=yx5=�4=a�3=��2=H�1=|1=�.0= E/=_Y.=k-=z,=v�+=�*=��)=�(=��'=��&=��%=�$=�z#=Oj"=�U!=�= =J!=	=��=�=R�=V=r =K�=��=Ud=]=��=]~=S(=x�=�m=�	=��	=�2=��=�I=1�=AN=�� =o��<�h�<zF�<\�<)��<c��<o�<�&�<"��<̀�<$�<���<X�<<��<�t�<|��<�|�<���<�q�<��<�U�<2·<�*�<U��<��<AR�<L��<�	�<Ob�<¸�<{�<�`�<���<��<cS�<���<c�<�z<�s<��k<EWd<��\<0�U<68N<��F<��?<�-8<5�0<�)<4B"<��<&�<o�<jL<[<�;J��;R��;�|�;h\�;�M�;ZQ�;�h�;%��;'�{;�W`;}3E;�?*;�};|��:-0�:���:�C:XN9��H����U�z�����8�ߺ���H���g7�s�N��e��|�}��쒔������L��Z񴻤o����ɻ��ӻ
޻�����W��Qi���4��:���^��s�5�!���%��*��;.�XI2�qI6�-<:��!>���A���E��I��AM���P���T�U'X���[��:_��b��*f���i���l�OWp��s���v�8Dz�K�}�sa����������,����Q��1ቼ�n��h���9���R��Β�����n�������������t���:��=���K������F
��\��������v���識�g���ߪ��W��/ϭ��F��/����5��A��� %������������]�����N����  �  �N=n�M=�M=|NL=��K=��J=wJ=�QI=�H=��G=DG=�KF=��E=R�D=� D=�;C=�uB=��A=��@=�@=�S?=��>=׼==��<=!<=(Q;=�:=L�9=2�8=�8=:,7=<S6=�x5=�4=\�3=��2=D�1=�1=�.0=$E/=YY.=k-=z,=l�+=�*=��)=�(=��'=&=��%=�$=�z#=Dj"=�U!=�= =L!==��=�=G�=V=v =T�=��=Sd=b=��=c~=J(=t�=�m=�	=��	=�2=��=�I=/�==N=�� =���<�h�<�F�<J�<)��<P��<o�<�&�<��<ր�<$�<��<X�<A��<�t�<j��<�|�<���<�q�<��<�U�<(·<�*�<W��<��<YR�<L��<�	�<Qb�<���<��<�`�<���<s�<bS�<���<g�<�z<ws<y�k<3Wd<�\<@�U<;8N<��F<��?<�-8<�0<��)<3B"<��<1�<g�<�L<|<�;T��;��;j|�;R\�;�M�;�Q�;�h�;��;��{;IW`;�3E;+@*;Z~;���:�0�:���:@D:�TN9R�H������z����l�ߺo����h7���N�S�e�<�|�#}��В��Ƃ���L��d��o����ɻ�ӻ�	޻������V��Bi���d��:���W��s�E�!���%��*��;.�LI2�LI6�<:�">�}�A�
�E���I��AM���P���T�u'X���[��:_��b��*f���i���l�DWp�̬s���v�$Dz�p�}�ta����������,�������Q��9ቼ�n��[���4���\���������s�����������~���P��<���D������F
��Z��������v��z識�g���ߪ��W��/ϭ��F��+����5��K���%��Ꜷ���|���[�����a����  �  ߋN=�M=�M=jTL=��K=?�J=vJ=3ZI=n�H=*�G=>G=�WF=��E=��D=D=�JC=�B=j�A=r�@=�0@=�g?=��>=��==I==�8<=j;=�:=s�9=��8= !8=�J7=)s6=��5=e�4=3�3=3=� 2=i=1=�W0=�o/={�.=��-= �,=ض+=��*=��)=��(=��'=V�&=��%=f�$=��#==�"=�!=�| =�a=�B=r=��=��=��=�f=/-=�=?�=�d=C=�=�p=!=Z�=�Q=T�	=
z==i�==3�=�=��<���<���<ݗ�<�b�<�%�<v��<���<�B�<��<���<�!�<(��<�B�<���<:M�<���<�C�<��<$(�<@��<���<la�<ð<p!�< }�<H֥<-�<���<CԚ<=%�<�t�<�<��<\�<u��<j�<izz<�s<X�k<�;d<��\<�kU<=N<;�F<�B?<p�7<6�0<D5)<m�!<_�<sN<�<��<3�;k��;��;UF�;�;O��;r�;s��;��;�x;"];��A;\�&;��;���:Y��:bir:�l
:�s9Gt����'���uv��t��q�eb$��
<��iS��~j�룀��⋻�����[����\��U���_2̻�cֻ~n໥S�&��Э�����c:����%W�����/�F����"���&��+�6/�A>3��87�d%;�e?���B�z�F�A\J�=N�"�Q��NU���X�$i\���_�_c�>�f�]3j��m��p�g9t��w��z��~�y����6��̓�a����C������?����$�������2�������:�������<��]����:�������3��C����)���������o������,���`���ds���骼{`���֭�M��Bð�n9��ï��*&��Ӝ�����犹�o��Wz�����  �  ыN=�M=�M=fTL=��K=7�J=zJ=@ZI=}�H=%�G=:G=�WF=��E=��D=D=�JC=u�B=e�A=l�@=�0@=�g?=��>=��==B==�8<=j;=�:=t�9=}�8= !8=�J7=1s6=��5=f�4=3�3=3=� 2=l=1=�W0=�o/=y�.=��-=�,=ܶ+=��*=��)=��(=��'=\�&=��%=o�$=��#=;�"=	�!=�| =�a=�B=v=��=��=��=�f=@-=�=?�=�d=F=�=q==R�=�Q=J�	=z==l�==3�=�=��<���<���<ڗ�<�b�<�%�<x��<���<�B�<���<���<"�<N��<�B�<���<5M�<���<�C�<��<)(�<=��<���<ga�<�°<�!�<<}�<Q֥<�,�<���<=Ԛ<3%�<�t�<�<��<�[�<p��<|�<nzz<�s<O�k<�;d<��\<�kU<=N< �F<�B?<8�7<I�0<95)<^�!<Z�<VN<<��<�3�;=��;���;
F�;��;l��;Q�;���;C�;ˊx;�];��A;��&;g�;Ȍ�:|��:�ir:�j
:t9�s��k�'��󅺵w��s�8q�Nb$��
<��iS��~j�ͣ���⋻#��������]��.����2̻�cֻ�n໸S����L�������:����ZW�����/�L����"���&��+�56/�->3�U87�D%;�e?���B�p�F�a\J�.N�B�Q�OU���X�Hi\�z�_��^c�0�f�a3j��m��p�F9t��w�G�z��~������6��̓�a����P������'����$�������2�������:������=��X����:��Ʒ���3��O����)���������|������1���k���Ys��ꪼ�`���֭�M��0ð�k9������/&��͜�����֊��n��ez�����  �  ͋N=�M=�M=gTL=��K=9�J=|J=3ZI=u�H="�G=GG=�WF=��E=��D=	D=�JC=v�B=o�A=w�@=0@=�g?=��>=��==?==�8<=j;=�:=w�9={�8=!8=�J7=0s6=��5=^�4=1�3=3=� 2=]=1=�W0=�o/=�.=��-=�,=�+=��*=��)=��(=��'=W�&=��%=i�$=��#=I�"=�!=} =�a=�B=�=��=��=��=�f=5-=�=E�=�d=J=
�=q==U�=�Q=D�	=z==h�==1�=�=��<���<���<��<�b�<�%�<~��<���<�B�<���<���<�!�<:��<�B�<���<LM�<���<�C�<��<1(�<M��<���<�a�<�°<}!�<"}�<P֥<-�<���<DԚ<-%�<�t�<�<��<�[�<e��<u�<@zz<�s<B�k<�;d<��\<�kU<,N<�F<�B?<)�7<b�0<15)<c�!<\�<ZN<<�<O3�;%��;0��;9F�;�;���;%�;���;N�;q�x;z];s�A;�&;��;e��:<��:�jr:Ij
:dv9�q����'�`�Qx��$s��q��b$��
<�jS��~j�F����⋻S����졻T���-]�������2̻�cֻ�n໌S�����������:�u��SW�����/�P����"��&��+�06/�C>3��87�a%;�L?���B�]�F�x\J�N�F�Q�OU���X�bi\�~�_�2_c�>�f�a3j��m�2�p�}9t���w�b�z�k~������6��̓�"a����V������@����$�������2��r����:��p���=��O����:�������3��V����)���������w������+���q���Js��ꪼo`���֭�M��7ð��9������5&��Μ���������v��iz�����  �  ΋N=�M=�M=kTL=��K=>�J=}J=:ZI=}�H=)�G=BG=�WF=��E=��D=D=�JC={�B=g�A=s�@=�0@=�g?=��>=��==A==�8<=	j;=�:=q�9={�8= !8=�J7=.s6=��5=h�4=+�3=�3=� 2=c=1=�W0=�o/=v�.=��-=�,=ܶ+=��*=��)=��(=��'=Y�&=��%=u�$=��#=@�"=�!=�| =�a=�B=|=��=��=��=�f=>-=�=H�=�d=J=�=�p==N�=�Q=G�	=z==k�==*�=�=��<���<���<ؗ�<�b�<�%�<q��<���<�B�<���<���<�!�<K��<�B�<���<:M�<���<�C�<��<.(�<I��<���<ua�< ð<�!�<3}�<Q֥<-�<���<JԚ</%�<�t�<�<��<�[�<k��<q�<bzz<�s< �k<~;d<��\<�kU<2N<�F<�B?<,�7<;�0<-5)<q�!<P�<pN<<��<�3�;a��;��;.F�;'�;���;t�;���;}�;�x;8];�A;��&;�;ލ�:���:�jr:�k
:�r9	u����'����w��=s躶q�b$�B<�sjS�~j�����⋻-���"�����/]��1����2̻�cֻ�n�dS���\������z:����EW�����/�>����"���&��+�%6/�>3�[87�U%;�<?���B�\�F�`\J�5N�J�Q�!OU���X�Qi\���_�_c�.�f�~3j� �m��p�l9t���w�R�z��~������6��̓�a����T������5����$�������2�������:��x����<��S����:�������3��K����)���������i������%���o���_s��ꪼ�`���֭�M��;ð�q9��į��F&��؜�����䊹�s��hz�����  �  ԋN=�M=�M=hTL=��K=?�J=tJ=@ZI=|�H=*�G=DG=�WF=��E=��D=D=�JC=��B=p�A=w�@=�0@=�g?=��>=��==F==�8<=j;=�:=r�9=��8=� 8=�J7='s6=��5=^�4='�3=�3=� 2=b=1=�W0=�o/=u�.=��-=�,=ڶ+=��*=��)=��(=��'=T�&=��%=n�$=��#=C�"=�!=�| =�a=�B={=��=��=��=�f=?-=�=A�=�d=E=�=�p==P�=�Q=G�	=z==^�==&�=�=��<���<���<͗�<�b�<�%�<p��<���<�B�<��<���<�!�<K��<�B�<���<FM�<���<�C�<*��<2(�<T��<���<za�<	ð<�!�<@}�<A֥<-�<���<BԚ<5%�<�t�<�<��<�[�<f��<Y�<Lzz<�s<=�k<b;d<��\<mkU<#N<�F<�B?<B�7<:�0<55)<f�!<V�<rN<�<��<�3�;p��;��;�F�;m�;���;��;���;��;��x;�];�A;��&;c�;ӌ�:8��:/jr:�k
:tt9�s���'�V􅺙w��t�r��b$�s<�7jS�-j����㋻,���)������\��;����2̻�cֻ�n່S�3��C������a:����W�����/�����"���&��+�6/�0>3�U87�_%;�U?���B�l�F�]\J�9N�7�Q�OU���X�Oi\���_�_c�_�f�|3j��m�=�p�~9t� �w�J�z��~������6��̓�a����H������/����$�������2��w����:��~����<��N���|:�������3��C����)���������l������.���j���bs���骼�`���֭�M��Sð�|9��կ��6&��朶��������z��fz�����  �  ʋN=�M=�M=iTL=��K=?�J=}J=@ZI=z�H=/�G=LG=�WF=��E=��D=D=�JC=��B=o�A=��@=�0@=�g?=��>=��==G==�8<=j;=�:=k�9=v�8=� 8=�J7='s6=��5=T�4=&�3=�3=� 2=_=1=�W0=�o/=p�.=��-=�,=۶+=��*=��)=��(=��'=[�&=��%=k�$=��#=I�"=�!=} =�a=�B=�=��=��=��=�f=@-=�=C�=�d=E=�=�p==J�=�Q=@�	=z==T�==%�=�=��<���<���<̗�<�b�<�%�<t��<���<�B�<��<���<�!�<G��<�B�<���<FM�<���<�C�<'��<<(�<\��<���<�a�<ð<�!�<A}�<S֥<-�<���<DԚ<3%�<�t�<�<��<�[�<b��<c�<6zz<qs<6�k<O;d<��\<�kU<"N<�F<�B?<�7<3�0<35)<i�!<]�<tN<<��<{3�;���;^��;hF�;�;���;��;��;��;��x;M];H�A;��&;{�;���:s��:�jr:�k
:�v9�v����'��zx���s��q�Lc$�v<�4jS��j�+����⋻N���K�����[]��0����2̻�cֻwnເS����5������>:�s��"W�����/�����"���&��+��5/�2>3�O87�H%;�L?���B�h�F�d\J�1N�f�Q�)OU��X�ei\���_�'_c���f�x3j��m�f�p�|9t��w�h�z��~������6��̓�a����G������-����$�������2��v����:��j����<��D���s:�������3��7����)���������n������+���k���as��ꪼ�`���֭�M��Hð��9��௳�:&�������z��yz�����  �  ɋN=�M=�M=hTL=��K=<�J=�J=BZI=��H=.�G=LG=�WF=��E=��D=D=�JC=��B=t�A=~�@=�0@=�g?=��>=��==C==�8<=j;=�:=o�9=y�8=� 8=�J7=!s6=��5=W�4=�3=�3=� 2=X=1=�W0=�o/=l�.=��-=�,=۶+=��*=��)=��(=��'=]�&=��%=x�$=��#=L�"=�!=} =�a=�B=�=��=�=��=�f=E-=�=E�=�d=G=�=�p==N�=�Q=;�	=�y==X�=�=�=�=��<��<���<Ǘ�<�b�<�%�<g��<���<�B�<���<���<"�<X��<�B�<���<QM�<���<�C�<)��<F(�<g��<���<�a�<ð<�!�<E}�<]֥<-�<���<DԚ<(%�<�t�<�<��<�[�<U��<N�<(zz<ws<��k<J;d<��\<UkU<N<ݢF<�B?<�7<<�0<5)<c�!<W�<hN<#<��<�3�;���;^��;�F�;��;��;��;K��;�;�x;];��A;W�&;��;m��:��:Nkr:�k
:Wr9�t����'���y���t�Ur�c$��<�kS�Jj�X���!㋻n���f�|���U]��(����2̻�cֻ�n�pS�������p��K:�d��W�����/�����"���&��+��5/�>3�987�A%;�??���B�_�F�s\J�6N�c�Q�OU��X�vi\���_�C_c�n�f��3j�0�m�T�p��9t�8�w�z�z��~������6��̓�a����P������(����$�������2��k����:��Y����<��:���i:�������3��<����)���������p������,���v���]s��ꪼ�`���֭�"M��^ð��9��ݯ��V&��𜶼����������z�����  �  ȋN= �M=�M=iTL=��K=B�J=J=AZI=��H=3�G=SG=�WF=��E=��D=*D=�JC=��B=�A=��@=�0@=�g?=��>=��==H==�8<=j;=�:=k�9=v�8=� 8=�J7=s6=��5=Q�4=�3=�3=� 2=S=1=�W0=�o/=f�.=��-=�,=ֶ+=��*=��)=��(=��'=\�&=��%=z�$=��#=R�"=#�!=} =b=�B=�=��=�=��=�f=?-=�=G�=�d=C=�=�p=
=G�=�Q=>�	=�y=�=N�=�=�=�=��<x��<���<���<�b�<�%�<b��<���<�B�<��<���<"�<N��<�B�<���<cM�<��<�C�<E��<R(�<c��<���<�a�<ð<�!�<A}�<V֥<-�<���<DԚ<0%�<�t�<�<��<�[�<\��<C�<zz<Vs<��k<,;d<��\<<kU<
N<�F<dB?<�7<)�0<*5)<g�!<\�<~N<<��<�3�;���;���;�F�;��;��;H�;:��;/�;��x;�];��A;*�&;��;U��:�:Xkr:~l
:ms9v����'�_����x���t躹r�^c$� <�kS��j�}���N㋻L���������b]��M����2̻�cֻtn�GS����7���h��9:�J���V����[/�߂���"���&��+��5/��=3�N87�E%;�5?���B�h�F�d\J�GN�j�Q�.OU�8�X�gi\���_�Z_c���f��3j�;�m�o�p��9t�B�w�m�z��~������6��̓�a����E������)����$�������2��X����:��b����<��.���m:�������3��0����)���������e������,���o���fs��ꪼ�`���֭�M��hð��9����T&����������������z�����  �  ɋN=��M=�M=gTL=��K=B�J=�J=LZI=��H=<�G=RG=�WF=��E=��D=,D=�JC=��B=y�A=��@=�0@=�g?=��>=��==I==�8<=j;=�:=b�9=v�8=� 8=�J7=s6=��5=L�4=�3=�3=� 2=X=1=�W0=�o/=d�.=��-=	�,=Ӷ+=��*=��)=��(=��'=e�&=��%=z�$=¶#=Q�"=#�!=} =b=�B=�=��=�=��=�f=E-=$�=D�=�d=B=
�=�p==E�=�Q=2�	=�y==E�=�=�=�=��<k��<���<���<�b�<�%�<a��<���<�B�<��<���<"�<Q��<�B�<���<ZM�<��<�C�<F��<V(�<v��<���<�a�<,ð<�!�<V}�<b֥<-�<���<AԚ<.%�<�t�<�<��<�[�<F��<G�<zz<0s<��k<;d<��\<LkU<�N<͢F<iB?<�7<�0<&5)<_�!<Z�<}N<%<��<�3�;	��;���;�F�;��;?��;[�;u��;[�;b�x;�];q�A;0�&;q�;T��:��:Xkr:Bl
:�t99z����'���Yy��qu�Zr��c$�R<��jS�]�j�Q���X㋻����������n]��g����2̻�cֻjn�_S껛������e��:�M���V����_/�����"���&��+��5/��=3�487�%;�>?���B�m�F�d\J�QN�|�Q�1OU�9�X��i\���_�F_c���f��3j�E�m���p��9t�Y�w���z��~������6��̓�a����B����������$�������2��a���z:��R����<��*���Z:�������3�� ����)���������g������/���q���us��ꪼ�`���֭�0M��cð��9������V&���������������z�����  �  N= �M=�M=fTL=��K=?�J=�J=FZI=��H=<�G=VG=�WF=��E=��D=%D=�JC=��B=��A=��@=�0@=�g?=��>=��==G==�8<=j;=�:=j�9=p�8=� 8=�J7=s6=��5=H�4=�3=�3=� 2=J=1=�W0=�o/=h�.=��-=�,=ڶ+=��*=��)=��(=��'=b�&=��%=~�$=��#=Z�"=&�!=} =b=�B=�=��=�=��=�f=A-=�=D�=�d=E=�=�p==C�=�Q=,�	=�y=�=F�=�=�=�=��<b��<���<���<�b�<�%�<g��<���<�B�<���<���<
"�<O��<�B�<���<pM�<��<�C�<=��<^(�<���<���<�a�<*ð<�!�<K}�<`֥<-�<���<CԚ<'%�<�t�<�<��<�[�<>��<4�<�yz<?s<Ҥk<;d<b�\< kU<�N<ɢF<lB?<��7<*�0<5)<Z�!<b�<uN<!<��<�3�;��;���;"G�;8�;r��;&�;���;��;*�x;�];u�A;_�&;%�;���::�lr:�k
:�x9�u���'�&��y���u�s��c$��<�kS�+�j�����z㋻���������y]��(����2̻�cֻ\n�`S껵�����T��$:�(���V�M��W/����T�"���&�v+��5/��=3�B87�)%;�<?���B�^�F�\J�6N�w�Q�7OU� �X��i\���_�_c���f��3j�a�m���p��9t�f�w���z��~������6��̓�'a����F����������$�������2��J���v:��<����<��!���G:�������3��#����)���������i������-���x���bs��#ꪼ�`���֭�8M��vð��9������j&���������������z�����  �  ��N=��M=�M=iTL=��K=A�J=�J=EZI=��H=:�G=VG=�WF=��E=��D=,D=�JC=��B=��A=��@=�0@=�g?=��>=��==E==�8<=j;=�:=i�9=g�8=� 8=�J7=s6=��5=K�4=�3=�3=� 2=D=1=�W0=�o/=]�.=��-=�,=ֶ+=��*=��)=��(=��'=f�&=��%=��$=��#=\�"=!�!=} =
b=�B=�=��=�=��=�f=E-=!�=J�=�d=E=�=�p==9�=�Q=*�	=�y=�=I�=�=	�=�=��<r��<���<���<�b�<�%�<[��<���<�B�<���<���<
"�<b��<�B�<���<vM�<��<�C�<J��<i(�<t��<���<�a�<%ð<�!�<J}�<n֥<-�<���<GԚ<!%�<�t�<�<��<�[�<H��<@�<�yz<Js<��k<;d<X�\<,kU<�N<��F<LB?<��7<&�0<5)<f�!<S�<~N<F<��<>4�;���;���;/G�;��;���;i�;���;E�;\�x;�];��A;�&;(�;��:���:3lr:%l
:fr9v��M�'�e���vz���t�.s��c$�t<��kS��j��/㋻�����������]��F����2̻�cֻ�n�)S껏������*��4:� ���V�n��9/��i�"���&�k+��5/��=3�.87� %;�!?���B�[�F�|\J�DN���Q�\OU�O�X��i\���_��_c���f��3j�d�m�~�p��9t�C�w���z��~������6��!̓�#a����O����������$��s����2��D����:��=����<�����\:�������3��(����)���������c������)���~���gs��0ꪼ�`��׭�-M��jð��9��񯳼}&���������������z����  �  ɋN=��M=�M=hTL=��K=B�J=�J=IZI=��H==�G=YG=�WF=��E=��D=0D=�JC=��B=��A=��@=�0@=�g?=��>=��==I==�8<=j;=�:=j�9=t�8=� 8=�J7=s6=��5=B�4=�3=�3=� 2=D=1=�W0=�o/=c�.=��-=�,=Ѷ+=��*=��)=��(=��'=e�&=��%=~�$=ö#=]�"=0�!=} =
b=�B=�=�=�=��=�f=C-=!�=E�=�d=?=�=�p=
=C�=�Q='�	=�y=�=?�=�=�=�=��<T��<���<���<�b�<�%�<Q��<���<�B�<���<���<"�<V��<�B�<���<yM�<��<�C�<O��<m(�<���<���<�a�<.ð<�!�<P}�<g֥<-�<���<@Ԛ<%%�<�t�<�<��<�[�<1��<.�<�yz<)s<��k< ;d<J�\<kU<�N<��F<iB?<�7<�0<
5)<`�!<P�<�N</<��<�3�;��;ц�;dG�;;�;���;��;���;��;��x;];��A;��&;Z�;��:J��:Ykr:�l
:no9�t����'����y��sv�ks�5d$��<��kS�~�j�餀��㋻����������C]��m����2̻�cֻon�ES껚������S��:����V�T��9/�ł�X�"�X�&�e+��5/��=3�887�%;�4?���B�o�F�n\J�\N�b�Q�1OU�7�X��i\��_��_c���f��3j�i�m���p��9t�~�w���z��~������6��*̓�a����D����������$��|����2��@���g:��;����<�����J:��t����3������)���������d������0���z���os��ꪼ�`���֭�EM��|ð��9�����q&��������#�������z�����  �  ��N=��M=�M=hTL=��K=D�J=�J=VZI=��H=E�G=WG=�WF=��E=��D=2D=�JC=��B=��A=��@=�0@=�g?=��>=��==O==�8<=	j;=�:=f�9=e�8=� 8=�J7=s6=��5=B�4=�3=�3=� 2=P=1=�W0=�o/=c�.=y�-=�,=϶+=��*=��)=��(=��'=h�&=��%=��$=ζ#=R�"=)�!=} =
b=�B=�=�=�=��=�f=L-=(�=B�=�d===
�=�p= =1�=�Q=/�	=�y=�=:�=�=�=�=��<X��<���<���<�b�<�%�<Y��<���<�B�<��<���<#"�<^��<�B�<���<dM�<��<�C�<R��<l(�<���<���<�a�<Bð<�!�<h}�<a֥<-�<���<>Ԛ<3%�<�t�<�<��<�[�<<��<:�<�yz<s<դk<�:d<b�\<1kU<�N<ʢF<(B?<��7<	�0<*5)<b�!<c�<�N<<�<�3�;S��;�;!G�;6�;���;��;���;��;�x;P];��A;��&;�;k��:#��:�kr:wm
:}u9,w����'����0y��6v躬r�3d$��<�ukS�ŀj������㋻������?����]������2̻�cֻ&n�TS껀������K���9�E���V�]��9/��d�"�r�&��+��5/��=3�87�%;�@?���B�y�F�]\J�aN���Q�xOU�C�X��i\��_�\_c���f��3j�k�m���p��9t�u�w���z��~������6��"̓�a����4����������$��w����2��V���n:��C����<�����L:�������3������)��z������d���{��2���k���ts��-ꪼ�`���֭�9M��pð��9��
���h&���������������z����  �  ɋN=��M=�M=hTL=��K=B�J=�J=IZI=��H==�G=YG=�WF=��E=��D=0D=�JC=��B=��A=��@=�0@=�g?=��>=��==I==�8<=j;=�:=j�9=t�8=� 8=�J7=s6=��5=B�4=�3=�3=� 2=D=1=�W0=�o/=c�.=��-=�,=Ѷ+=��*=��)=��(=��'=e�&=��%=~�$=ö#=]�"=0�!=} =
b=�B=�=�=�=��=�f=C-=!�=E�=�d=@=�=�p=
=C�=�Q='�	=�y=�=?�=�=�=�=��<U��<���<���<�b�<�%�<Q��<���<�B�<���<���<"�<V��<�B�<���<yM�<��<�C�<O��<m(�<���<���<�a�<-ð<�!�<O}�<g֥<-�<���<@Ԛ<$%�<�t�<�<��<�[�<1��<.�<�yz<)s<��k< ;d<J�\<kU<�N<��F<iB?<�7<�0<
5)<`�!<P�<�N</<��<�3�;��;ц�;dG�;;�;���;��;���;��;��x;];��A;��&;X�;��:F��:Pkr:�l
:Ho9u���'����y��xv�ms�8d$��<��kS���j�꤀��㋻����������C]��n����2̻�cֻpn�FS껛������S��:����V�T��9/�ł�X�"�X�&�e+��5/��=3�887�%;�4?���B�o�F�n\J�\N�b�Q�1OU�7�X��i\��_��_c���f��3j�i�m���p��9t�~�w���z��~������6��*̓�a����D����������$��|����2��@���g:��;����<�����J:��t����3������)���������d������0���z���os��ꪼ�`���֭�EM��|ð��9�����q&��������#�������z�����  �  ��N=��M=�M=iTL=��K=A�J=�J=EZI=��H=:�G=VG=�WF=��E=��D=,D=�JC=��B=��A=��@=�0@=�g?=��>=��==E==�8<=j;=�:=i�9=g�8=� 8=�J7=s6=��5=K�4=�3=�3=� 2=D=1=�W0=�o/=]�.=��-=�,=ֶ+=��*=��)=��(=��'=f�&=��%=��$=��#=\�"=!�!=} =
b=�B=�=��=�=��=�f=F-=!�=J�=�d=E=�=�p==9�=�Q=*�	=�y=�=J�=�=
�=�=��<s��<���<���<�b�<�%�<[��<���<�B�<���<���<"�<c��<�B�<���<vM�<��<�C�<J��<i(�<t��<���<�a�<%ð<�!�<J}�<n֥<-�<���<GԚ< %�<�t�<�<��<�[�<H��<@�<�yz<Js<��k<;d<X�\<-kU<�N<��F<MB?<��7<'�0<5)<g�!<S�<~N<F<��<?4�;���;���;/G�;��;���;i�;���;E�;Z�x;�];��A;�&;%�;���:���:"lr:l
:r9+v��_�'�n���z���t�3s��c$�x<��kS��j�𤀻1㋻�����������]��G����2̻�cֻ�n�)S껐������+��4:� ���V�n��9/��i�"���&�k+��5/��=3�.87� %;�!?���B�[�F�|\J�DN���Q�\OU�O�X��i\���_��_c���f��3j�d�m�~�p��9t�C�w���z��~������6��!̓�#a����O����������$��s����2��D����:��=����<�����\:�������3��(����)���������c������)���~���gs��0ꪼ�`��׭�-M��jð��9��񯳼}&���������������z����  �  N= �M=�M=fTL=��K=?�J=�J=FZI=��H=<�G=VG=�WF=��E=��D=%D=�JC=��B=��A=��@=�0@=�g?=��>=��==G==�8<=j;=�:=j�9=p�8=� 8=�J7=s6=��5=H�4=�3=�3=� 2=J=1=�W0=�o/=h�.=��-=�,=ڶ+=��*=��)=��(=��'=b�&=��%=~�$=��#=Z�"=&�!=} =b=�B=�=��=�=��=�f=A-=�=D�=�d=E=�=�p==C�=�Q=,�	=�y=�=F�=�=�=�=��<c��<���<���<�b�<�%�<h��<���<�B�<���<���<"�<P��<�B�<���<pM�<��<�C�<=��<^(�<���<���<�a�<)ð<�!�<J}�<_֥<-�<���<CԚ<&%�<�t�<�<��<�[�<>��<4�<�yz<?s<Ҥk<;d<b�\< kU<�N<ɢF<mB?<��7<+�0<5)<[�!<c�<vN<"<��<�3�;��;���;"G�;8�;r��;&�;���;��;'�x;�];q�A;[�&; �;���:㩭:�lr:�k
:6x9�u��9�'�3��y���u�s��c$��<��kS�0�j�����|㋻����������{]��)����2̻�cֻ]n�aS껶�����T��$:�)���V�M��W/����T�"���&�v+��5/��=3�B87�)%;�<?���B�^�F�\J�6N�w�Q�7OU� �X��i\���_�_c���f��3j�a�m���p��9t�f�w���z��~������6��̓�'a����F����������$�������2��J���v:��<����<��!���G:�������3��#����)���������i������-���x���bs��#ꪼ�`���֭�8M��vð��9������j&���������������z�����  �  ɋN=��M=�M=gTL=��K=B�J=�J=LZI=��H=<�G=RG=�WF=��E=��D=,D=�JC=��B=y�A=��@=�0@=�g?=��>=��==I==�8<=j;=�:=b�9=v�8=� 8=�J7=s6=��5=L�4=�3=�3=� 2=X=1=�W0=�o/=d�.=��-=	�,=Ӷ+=��*=��)=��(=��'=e�&=��%=z�$=¶#=Q�"=#�!=} =b=�B=�=��=�=��=�f=E-=$�=D�=�d=B=
�=�p==E�=�Q=2�	=�y==E�=�=�=�=��<k��<���<���<�b�<�%�<a��<���<�B�<��<���<"�<Q��<�B�<���<ZM�<��<�C�<F��<V(�<u��<���<�a�<,ð<�!�<V}�<a֥<-�<���<@Ԛ<-%�<�t�<�<��<�[�<F��<G�<zz<0s<��k<;d<��\<MkU<�N<͢F<jB?<�7<�0<'5)<`�!<[�<~N<&<��<�3�;
��;���;�F�;��;?��;[�;u��;Z�;_�x;�];m�A;+�&;k�;G��:��:;kr:$l
:>t9yz���'���iy���u�br��c$�Y<��jS�d�j�T���[㋻����������p]��i����2̻�cֻln�`S껜������f��:�N���V����`/�����"���&��+��5/��=3�487�%;�>?���B�m�F�d\J�QN�|�Q�1OU�9�X��i\���_�F_c���f��3j�E�m���p��9t�Y�w���z��~������6��̓�a����B����������$�������2��a���z:��R����<��*���Z:�������3�� ����)���������g������/���q���us��ꪼ�`���֭�0M��cð��9������V&���������������z�����  �  ȋN= �M=�M=iTL=��K=B�J=J=AZI=��H=3�G=SG=�WF=��E=��D=*D=�JC=��B=�A=��@=�0@=�g?=��>=��==H==�8<=j;=�:=k�9=v�8=� 8=�J7=s6=��5=Q�4=�3=�3=� 2=S=1=�W0=�o/=f�.=��-=�,=ֶ+=��*=��)=��(=��'=\�&=��%=z�$=��#=R�"=#�!=} =b=�B=�=��=�=��=�f=?-=�=G�=�d=D=�=�p==G�=�Q=>�	=�y=�=O�=�=�=�=��<y��<���<���<�b�<�%�<c��<���<�B�<��<���<"�<O��<�B�<���<dM�<��<�C�<E��<R(�<c��<���<�a�<ð<�!�<A}�<U֥<-�<���<CԚ</%�<�t�<�<��<�[�<\��<C�<zz<Vs<��k<,;d<��\<=kU<N<�F<eB?<�7<*�0<+5)<h�!<]�<N<<��<�3�;���;���;�F�;��;��;H�;9��;-�;��x;|];��A;$�&;��;F��:੭:8kr:\l
:�r9^v���'�q����x���t��r�fc$�(<�kS��j�����Q㋻O���������d]��O����2̻�cֻvn�HS����8���h��::�J���V����[/�߂���"���&��+��5/��=3�N87�E%;�5?���B�h�F�d\J�GN�j�Q�.OU�8�X�gi\���_�Z_c���f��3j�;�m�o�p��9t�B�w�m�z��~������6��̓�a����E������)����$�������2��X����:��b����<��.���m:�������3��0����)���������e������,���o���fs��ꪼ�`���֭�M��hð��9����T&����������������z�����  �  ɋN=�M=�M=hTL=��K=<�J=�J=BZI=��H=.�G=LG=�WF=��E=��D=D=�JC=��B=t�A=~�@=�0@=�g?=��>=��==C==�8<=j;=�:=o�9=y�8=� 8=�J7=!s6=��5=W�4=�3=�3=� 2=X=1=�W0=�o/=l�.=��-=�,=۶+=��*=��)=��(=��'=]�&=��%=x�$=��#=L�"=�!=} =�a=�B=�=��=�=��=�f=E-=�=E�=�d=G=	�=�p==N�=�Q=;�	=�y==X�= =�=�=��<���<���<ȗ�<�b�<�%�<h��<���<�B�<���<���<"�<Y��<�B�<���<RM�<���<�C�<)��<F(�<g��<���<�a�<ð<�!�<E}�<\֥<-�<���<CԚ<(%�<�t�<�<��<�[�<U��<M�<(zz<ws<��k<J;d<��\<VkU<N<ޢF<�B?<�7<=�0<5)<d�!<X�<iN<$<��<�3�;���;`��;�F�;��;��;��;J��;�;�x;];��A;P�&;��;^��:��:,kr:�k
:�q9�t����'���"y���t�]r�c$��<�kS�Qj�\���$㋻q���h�~���W]��*����2̻�cֻ�n�qS�������q��L:�e��W�����/�����"���&��+��5/�>3�987�A%;�??���B�_�F�s\J�7N�d�Q�OU��X�vi\���_�C_c�n�f��3j�0�m�T�p��9t�8�w�z�z��~������6��̓�a����P������(����$�������2��k����:��Y����<��:���i:�������3��<����)���������p������,���v���]s��ꪼ�`���֭�"M��^ð��9��ݯ��V&��𜶼����������z�����  �  ʋN=�M=�M=iTL=��K=?�J=}J=@ZI=z�H=/�G=LG=�WF=��E=��D=D=�JC=��B=o�A=��@=�0@=�g?=��>=��==G==�8<=j;=�:=k�9=v�8=� 8=�J7='s6=��5=T�4=&�3=�3=� 2=_=1=�W0=�o/=p�.=��-=�,=۶+=��*=��)=��(=��'=[�&=��%=k�$=��#=I�"=�!=} =�a=�B=�=��=��=��=�f=@-=�=C�=�d=F=�=�p==J�=�Q=@�	=z==T�==&�=�=��<���<���<͗�<�b�<�%�<u��<���<�B�<��<���< "�<H��<�B�<���<GM�<���<�C�<'��<<(�<\��<���<�a�<ð<�!�<@}�<S֥<-�<���<CԚ<3%�<�t�<�<��<�[�<a��<c�<6zz<qs<6�k<O;d<��\<�kU<"N<��F<�B?<�7<4�0<45)<j�!<_�<uN<<��<}3�;���;_��;iF�;��;���;��;��;��;��x;H];C�A;��&;t�;���:d��:�jr:�k
:Hv9�v����'�􅺌x���s��q�Tc$�~<�;jS��j�.����⋻Q���N�����]]��2����2̻�cֻxnແS����6������?:�s��"W�����/�����"���&��+��5/�2>3�O87�H%;�L?���B�h�F�d\J�1N�f�Q�)OU��X�ei\���_�'_c���f�x3j��m�f�p�|9t��w�h�z��~������6��̓�a����G������-����$�������2��v����:��j����<��D���s:�������3��7����)���������n������+���k���as��ꪼ�`���֭�M��Hð��9��௳�:&�������z��yz�����  �  ԋN=�M=�M=hTL=��K=?�J=tJ=@ZI=|�H=*�G=DG=�WF=��E=��D=D=�JC=��B=p�A=w�@=�0@=�g?=��>=��==F==�8<=j;=�:=r�9=��8=� 8=�J7='s6=��5=^�4='�3=�3=� 2=b=1=�W0=�o/=u�.=��-=�,=ڶ+=��*=��)=��(=��'=T�&=��%=n�$=��#=C�"=�!=�| =�a=�B={=��=��=��=�f=?-=�=B�=�d=E=�=�p==P�=�Q=G�	=z==^�==&�=�=��<���<���<Η�<�b�<�%�<q��<���<�B�<��<���<�!�<L��<�B�<���<FM�<���<�C�<*��<2(�<T��<���<za�<ð<�!�<@}�<@֥<-�<���<AԚ<4%�<�t�<�<��<�[�<f��<Y�<Lzz<�s<>�k<b;d<��\<nkU<$N<�F<�B?<C�7<;�0<65)<g�!<W�<sN<�<��<�3�;q��;��;�F�;m�;���;��;���;��;��x;�];
�A;��&;]�;ƌ�:*��:jr:�k
:�s9�s��6�'�f􅺨w��,t�r��b$�z<�>jS�3j����㋻/���+������\��=����2̻�cֻ�n້S�4��D������a:����W�����/�����"���&��+�6/�0>3�U87�_%;�U?���B�l�F�]\J�9N�7�Q�OU���X�Oi\���_�_c�_�f�|3j��m�=�p�~9t� �w�J�z��~������6��̓�a����H������/����$�������2��w����:��~����<��N���|:�������3��C����)���������l������.���j���bs���骼�`���֭�M��Sð�|9��կ��6&��朶��������z��fz�����  �  ΋N=�M=�M=kTL=��K=>�J=}J=:ZI=}�H=)�G=BG=�WF=��E=��D=D=�JC={�B=g�A=s�@=�0@=�g?=��>=��==A==�8<=	j;=�:=q�9={�8= !8=�J7=.s6=��5=h�4=+�3=�3=� 2=c=1=�W0=�o/=v�.=��-=�,=ܶ+=��*=��)=��(=��'=Y�&=��%=u�$=��#=@�"=�!=�| =�a=�B=|=��=��=��=�f=>-=�=H�=�d=J=�=�p==N�=�Q=G�	=z==l�==*�=�=��<���<���<ٗ�<�b�<�%�<r��<���<�B�<���<���<�!�<K��<�B�<���<;M�<���<�C�<��<.(�<H��<���<ua�< ð<�!�<3}�<Q֥<-�<���<JԚ<.%�<�t�<�<��<�[�<j��<q�<bzz<�s< �k<;d<��\<�kU<3N<�F<�B?<-�7<<�0<.5)<r�!<Q�<qN<<��<�3�;b��;��;/F�;(�;���;s�;���;|�; �x;5];�A;��&;�;Ӎ�:���:ojr:�k
:Jr9=u����'����w��Is躼q�#b$�G<�yjS��~j�����⋻/���$�����0]��2����2̻�cֻ�n�eS���]������z:����FW�����/�>����"���&��+�%6/�>3�[87�U%;�=?���B�\�F�`\J�5N�J�Q�!OU���X�Qi\���_�_c�.�f�~3j� �m��p�l9t���w�R�z��~������6��̓�a����T������5����$�������2�������:��x����<��S����:�������3��K����)���������i������%���o���_s��ꪼ�`���֭�M��;ð�q9��į��F&��؜�����䊹�s��hz�����  �  ͋N=�M=�M=gTL=��K=9�J=|J=3ZI=u�H="�G=GG=�WF=��E=��D=	D=�JC=v�B=o�A=w�@=0@=�g?=��>=��==?==�8<=j;=�:=w�9={�8=!8=�J7=0s6=��5=^�4=1�3=3=� 2=]=1=�W0=�o/=�.=��-=�,=�+=��*=��)=��(=��'=W�&=��%=i�$=��#=I�"=�!=} =�a=�B=�=��=��=��=�f=5-=�=E�=�d=J=
�=q==U�=�Q=D�	=z==h�==2�=�=��<���<���<��<�b�<�%�<~��<���<�B�<���<���<�!�<;��<�B�<���<LM�<���<�C�<��<1(�<M��<���<�a�<�°<}!�<!}�<P֥<-�<���<DԚ<-%�<�t�<�<��<�[�<d��<u�<?zz<�s<B�k<�;d<��\<�kU<-N<�F<�B?<*�7<c�0<25)<d�!<]�<[N<<�<P3�;&��;0��;9F�;�;���;%�;���;N�;o�x;w];p�A;�&;��;]��:4��:�jr:8j
:v9r����'�i�[x��-s��q��b$��
<�jS��~j�H����⋻U����졻U���/]�������2̻�cֻ�nໍS�����������:�u��SW�����/�Q����"��&��+�06/�C>3��87�a%;�L?���B�]�F�x\J�N�F�Q�OU���X�bi\�~�_�2_c�>�f�a3j��m�2�p�}9t���w�b�z�k~������6��̓�"a����V������@����$�������2��r����:��p���=��O����:�������3��V����)���������w������+���q���Js��ꪼo`���֭�M��7ð��9������5&��Μ���������v��iz�����  �  ыN=�M=�M=fTL=��K=7�J=zJ=@ZI=}�H=%�G=:G=�WF=��E=��D=D=�JC=u�B=e�A=l�@=�0@=�g?=��>=��==B==�8<=j;=�:=t�9=}�8= !8=�J7=1s6=��5=f�4=3�3=3=� 2=l=1=�W0=�o/=y�.=��-=�,=ܶ+=��*=��)=��(=��'=\�&=��%=o�$=��#=;�"=	�!=�| =�a=�B=v=��=��=��=�f=@-=�=?�=�d=F=�=q==R�=�Q=K�	=z==l�==3�=�=��<���<���<ڗ�<�b�<�%�<y��<���<�B�< ��<���<"�<O��<�B�<���<5M�<���<�C�<��<)(�<=��<���<ga�<�°<�!�<<}�<Q֥<�,�<���<=Ԛ<3%�<�t�<�<��<�[�<o��<|�<nzz<�s<O�k<�;d<��\<�kU<=N< �F<�B?<8�7<I�0<95)<^�!<[�<VN<<��<�3�;=��;���;F�;��;l��;Q�;���;C�;ʊx;�];��A;��&;e�;Č�:x��:�ir:�j
:�s9�s��t�'��󅺺w��s�;q�Pb$��
<��iS��~j�Σ���⋻$��������]��.����2̻�cֻ�n໸S����M�������:����ZW�����/�L����"���&��+�56/�->3�V87�D%;�e?���B�p�F�a\J�.N�B�Q�OU���X�Hi\�z�_��^c�0�f�a3j��m��p�F9t��w�G�z��~������6��̓�a����P������'����$�������2�������:������=��X����:��Ʒ���3��O����)���������|������1���k���Ys��ꪼ�`���֭�M��0ð�k9������/&��͜�����֊��n��ez�����  �  �N=��M=aM=�ZL=j�K=��J=�!J=QcI=F�H=��G=�$G=�cF=��E=��D=�D=QZC=�B=��A=�
A=D@=|?=.�>="�====�Q<=
�;=�:=��9=9=�?8=k7=��6=~�5=��4=�4=�(3=-I2=Cg1=�0=��/=ӳ.=v�-=��,=��+=S�*=��)=n)=�	(=�	'=�&=��$=��#=��"=��!=�� =:�=M�=f=�?=�=3�=�=Rx=�:=�=S�=,e='=�="c=*=9�=Y4
=��=�Q=a�=&\=7�=�S=D��<Br�<�J�<��<���<S��<eZ�<�<���<W�<���<U��<��<��<�$�<m��<�<���<��<�m�<�ջ<:�<���<8��<�R�<7��<>��<�Q�<���<�<>�<r��<�ӏ<��<�d�<w��<��<�tz<<s<�k<od<��\<�>U<��M<�fF<~�><C�7<O70<��(<�!<�*<��<��<3L<;�;���;%O�;m��;g��;Œ�;'x�;Ip�;�}�;�@u;N�Y;�T>;�&#;,-;B��: ��:Kb:�W�9���8���� �9���F������T;��<)�Z�@��`X�Ȁo��)���l��#���8|���H����~kĻ�λ��ػ3��+�컯���� �[��`p	���Ԅ����S�,����#��(�&.,�U>0�x@4��48�<���?���C��G��8K��N���R�V���Y��%]���`�Pd�|wg���j�a0n��q�{�t��x�`N{�n�~�b܀��r����������'�����Y@���ɋ�/Q���֎�[���ݑ��^��ߔ��]��7ۗ��W��Ӛ��M��_ǝ�g@������<0��H����������	��s�������i���ޭ��S��tȰ�S=��Q���g'������C�����^����t��
콼�  �  �N=��M=bM=�ZL=k�K=��J=�!J=ScI=Q�H=��G=�$G=�cF=��E=��D=�D=VZC=�B=��A=�
A=D@=|?=.�>="�==�==�Q<=�;=�:=��9=9=�?8=k7=��6=��5=��4=�4=�(3=0I2=Cg1="�0=��/=ӳ.=q�-=�,=��+=R�*=��)=j)=�	(=�	'=�&=��$=��#=��"=��!=� =5�=G�=f=�?=�=-�=�=Zx=�:=z�=L�=0e='="�=$c=&=9�=X4
=��=�Q=e�=#\=8�=�S=J��<Xr�<�J�<��<���<_��<yZ�<!�<���<W�<���<U��<��<��<�$�<o��<��<���<��<�m�<�ջ<
:�<���</��<�R�<=��<=��<�Q�<���<$�<>�<���<�ӏ<��<�d�<���<��<�tz<Gs<��k<}d<�\<�>U<��M<�fF<s�><=�7<w70<��(<�!<�*<��<��<9L<��;j��;O�;f��;]��;���;�w�;rp�;�}�;�@u;�Y;�T>;h'#;'-;-��:z��:b:�W�9/��8�����9�?�����+��;��<)��@��`X���o��)���l�����>|���H����%kĻ
�λ��ػT��I�컷���� �9��rp	���������S�C��{�#��(�#.,�l>0�b@4�f48�<���?���C��G��8K���N���R�&V���Y��%]�֞`�Hd�mwg���j�^0n�ہq�m�t��x�qN{�q�~�h܀��r����������'�� ���\@���ɋ�Q���֎�[���ݑ�_���ޔ��]��<ۗ��W��#Ӛ��M��hǝ�R@������=0��R����������	��_�������i���ޭ��S��lȰ�X=��L���r'������G�����O����t��콼�  �  �N=��M=ZM=�ZL=m�K=��J=�!J=OcI=T�H=��G=�$G=�cF=��E=��D=�D=bZC=�B=��A=�
A=D@= |?=)�>=)�==�==�Q<=�;=�:=��9=9=�?8=k7=��6=w�5=��4=�4=�(3=-I2=8g1=�0=��/=ҳ.=t�-=|�,=��+=K�*=��)=i)=�	(=�	'=�&=��$=��#=��"=��!=
� =8�=I�=#f=�?=�=.�=�=Vx=�:=��=L�=6e= = �= c='=;�=P4
=��=�Q=`�=\=4�=�S=2��<Sr�<�J�<��<~��<T��<qZ�<�<���<W�<���<K��<��<��<�$�<��<��<���<��<�m�<�ջ<
:�<Κ�<-��<�R�<7��<H��<�Q�<���<*�<	>�<���<�ӏ<��<�d�<{��<��<�tz<Fs<�k<d<˭\<�>U<��M<�fF<��><6�7<p70<h�(<�!<�*<��<��<(L<��;]��;MO�;���;w��;��;�w�;�p�;�}�;Au;m�Y;�T>;�'#;�,;?��:���:Ab:�V�9V��8ق���9�^������O��;�0=)��@��`X�Ào�>*���l��L���>|���H����$kĻ@�λ��ػX���컪���� �3��qp	�m�������S�;��T�#��(��-,�g>0�_@4�s48�<���?���C��G��8K���N���R� V���Y��%]���`�td�|wg���j�h0n��q���t��x��N{�X�~�i܀��r����������'�����L@���ɋ�Q���֎�[���ݑ�
_���ޔ��]��/ۗ��W��#Ӛ��M��jǝ�M@������20��I����������	��_�������i���ޭ��S��vȰ�k=��L���w'������Z��&���S����t��콼�  �  �N=��M=_M=�ZL=h�K=��J=�!J=UcI=T�H=��G=�$G=�cF=��E=��D=�D=]ZC=�B=��A=�
A=D@=|?=/�>=(�==�==�Q<=�;=�:=��9=9=�?8=k7=��6=z�5=��4=�4=�(3=)I2=>g1=�0=��/=̳.=s�-=}�,=��+=O�*=��)=e)=�	(=�	'=�&=��$=��#=��"=��!=� ==�=N�=f=�?=�=/�=�=Xx=�:=��=H�=/e=#=�= c=%=2�=P4
=��=�Q=\�=\=-�=�S=8��<Cr�<�J�<��<z��<S��<nZ�<�<���<W�<���<T��<��<��<�$�<w��<��<���<��<�m�<�ջ<:�<͚�<8��<�R�<B��<E��<�Q�<x��<"�<>�<{��<�ӏ<��<�d�<s��<��<�tz<+s<�k<]d<ۭ\<�>U<��M<�fF<h�><2�7<`70<{�(<�!<�*<��<��<CL<��;���;HO�;���;���;��;*x�;�p�;�}�;�@u;��Y;�T>;�'#;N-;4��:���:Qb:�W�9~��8V����9��������2��;��<)���@��`X���o�
*���l��G���m|���H����NkĻ�λ��ػr��"�컬���� �1��hp	�w��������S�%��g�#��(�.,�`>0�T@4�h48�<���?���C�	�G��8K��N���R�#V���Y��%]��`�_d��wg���j��0n��q���t��x��N{���~�k܀��r����������'��%���M@���ɋ�Q���֎�[���ݑ� _���ޔ��]��+ۗ��W��Ӛ��M��^ǝ�N@������60��K����������	��j�������i���ޭ��S��tȰ�`=��Y���s'��Ĝ��Q��#���]����t��콼�  �  �N=��M=^M=�ZL=l�K=��J=�!J=[cI=R�H=��G=�$G=�cF=��E=��D=�D=_ZC=%�B=��A=�
A=D@=|?=4�>=&�====�Q<=�;=�:=��9=9=�?8=k7=��6=s�5=��4=�4=�(3=I2=8g1=�0=��/=ʳ.=o�-={�,=��+=N�*=��)=m)=�	(=�	'=�&=��$=��#=��"=��!=� =?�=Q�="f=�?=�=7�=�=]x=�:=��=O�=,e="=�=c=!=.�=P4
=x�=�Q=Q�=\='�=�S=)��</r�<�J�<��<w��<K��<fZ�<�<���<W�<���<\��<��<��<�$�<���<�<���<�<�m�<�ջ<':�<̚�<E��<�R�<O��<F��<�Q�<���<�<>�<v��<�ӏ<��<�d�<k��<s�<�tz<�s<�k<0d<ĭ\<�>U<��M<�fF<N�><6�7<S70<s�(<�!<�*<��<��<[L<��;���;XO�;���;���;��;rx�;�p�;[~�;|Au;�Y;JU>;�'#;�-;��:���:�b:�V�9���8����Q�9�-���������;�c=)��@��`X���o�6*��m��M���x|���H����gkĻ�λ��ػ/���컈���z �&��Gp	�z��������S���T�#��(��-,�?>0�I@4�Q48��<���?���C��G��8K��N���R�/V�ϣY��%]�#�`�sd��wg���j��0n��q���t��x�|N{���~�k܀��r����������'�����Q@���ɋ�Q���֎�[���ݑ��^���ޔ��]��&ۗ��W��Ӛ��M��Rǝ�P@������50��D����������	��o�������i���ޭ��S���Ȱ�l=��p���v'��ڜ��\��9���h����t�� 콼�  �  ��N=��M=[M=�ZL=l�K=��J=�!J=WcI=Y�H=��G=�$G=�cF=��E=��D=�D=iZC=�B=��A=A=D@=&|?=2�>=-�====�Q<=�;=�:=��9=9=�?8=k7=��6=o�5=~�4=�4=�(3=I2=5g1=�0=��/=ų.=n�-=s�,=��+=L�*=��)=j)=�	(=�	'=�&=��$=��#=��"=��!=� =F�=Y�=+f=�?=�==�="�=]x=�:=��=K�=/e==�=c==)�=E4
=u�=�Q=N�=\="�=�S=��<(r�<�J�<��<m��<:��<hZ�<�<���<W�<���<W��<��<"��<%�<���<�<Α�<�<�m�<�ջ< :�<ܚ�<W��<�R�<G��<U��<�Q�<���<#�<>�<s��<�ӏ<��<�d�<a��<s�<�tz<�s<��k<-d<��\<�>U<|�M<�fF<U�><�7<F70<i�(<�!<�*<��<��<LL<��;��;�O�;���;���;l��;�x�;q�;+~�;�Au;n�Y;�U>;"(#;�-;��:���:;b:LX�9ڼ�8����d�9����w���6��<�x=)��@��aX���o�E*��m�������|��I��PkĻ*�λ��ػF�����g���� ���$p	�c��������S����.�#��(��-,�!>0�7@4�P48��<���?���C��G��8K��N�ՂR�7V�ۣY�&]�'�`��d��wg���j��0n��q���t��x��N{���~�s܀�s����������'�����E@���ɋ�Q���֎��Z���ݑ��^���ޔ��]��ۗ��W��Ӛ��M��@ǝ�C@������&0��B����������	��r�������i���ޭ��S���Ȱ�o=��q����'��ۜ��_��<���p���u��콼�  �  ؏N=��M=YM=�ZL=k�K=��J=�!J=XcI=b�H=��G=�$G=dF=��E=��D=�D=sZC=&�B=�A=A=D@=.|?=2�>=0�==�==�Q<=�;=�:=��9=9=�?8=�j7=��6=h�5=y�4=�4=�(3=I2=*g1=�0=��/=��.=m�-=p�,=��+=F�*=��)=h)=�	(=�	'=�&= %=��#=��"=��!=� =J�=Z�=4f=�?=�=9�=&�=cx=�:=��=G�=,e==�=c==#�==4
=r�=�Q=L�=\=�=�S=��< r�<�J�<��<]��<<��<eZ�<�<���<W�<���<V��<��<#��<%�<���<�<��<
�<n�<ֻ<4:�<뚴<L��<�R�<J��<Y��<R�<���< �<>�<y��<�ӏ<��<�d�<X��<e�<dtz<�s<��k<d<��\<�>U<l�M<mfF<N�><��7<S70<]�(<�!<�*<��<��<NL< �;��;�O�; �;+��;���;�x�;vq�;u~�;JBu;��Y;�U>;�(#;�-;���:j��:�b:�V�9*��8���9�9����<���Y��u<��=)�a�@�
bX���o��*��'m�������|��I��+;kĻX�λ��ػR�����Y���m ����<p	�;����z���S����#��(��-,�1>0�%@4�548��<���?���C��G��8K� �N�ۂR�>V��Y�&]�0�`��d��wg��j��0n�'�q���t��x��N{���~��܀��r����������'�����=@���ɋ��P���֎��Z���ݑ��^���ޔ��]��ۗ�zW���Қ��M��Kǝ�3@������#0��>����������	��m�������i���ޭ��S���Ȱ��=��w����'��㜶�p��J���w���u��콼�  �  ؏N=��M=XM=�ZL=o�K=��J=�!J=`cI=d�H=��G=�$G=dF=��E=��D=�D=vZC=1�B=�A=
A=D@=/|?=9�>=.�====�Q<=�;=�:=��9=	9=�?8=k7=��6=^�5=o�4=�4=�(3=I2="g1=�0=��/=��.=e�-=n�,=��+=J�*=��)=n)=�	(=�	'=�&=	 %=��#=��"=��!=� =R�=b�=5f=�?=�=?�=)�=ex=�:=��=M�=,e==�=c==�=>4
=f�=�Q=?�=\=�=�S=���<	r�<�J�<��<S��<7��<\Z�<�<���<W�<���<_��<��<,��<%�<���<0�<��<�<n�<ֻ<B:�<<[��<�R�<\��<R��<R�<���< �<>�<r��<�ӏ<��<�d�<S��<O�<Btz<�s<��k<�d<w�\<e>U<Z�M<zfF<&�><��7<A70<X�(<�!<�*< �<��<pL<0�;��;�O�;^ �;p��;⓲;�x�;�q�;�~�;�Bu;��Y;/V>;�(#;=.;���:2��:Nb:UX�9o��8+���h�9����P���9���<�M>)���@��aX�Q�o��*��wm�������|��CI��2\kĻ5�λ��ػ�����c���X ����p	�0�v��o��hS�͡���#�s(��-,�>0�@4�*48��<���?���C��G��8K��N��R�[V���Y�&]�V�`��d��wg��j��0n�Q�q���t�x��N{���~��܀��r����������'�����A@���ɋ��P���֎��Z���ݑ��^���ޔ�s]���ڗ�nW���Қ��M��>ǝ�,@��u���*0��;����������	��t�������i���ޭ��S���Ȱ��=�������'���������]�������u��2콼�  �  ۏN=��M=XM=�ZL=l�K=��J=�!J=gcI=a�H=��G=�$G=dF=��E=��D=�D=vZC=2�B=�A=A=D@=/|?=A�>=/�====�Q<=�;=�:=��9=9=�?8=�j7=��6=b�5=m�4=�4=�(3=I2=+g1=��0=��/=��.=`�-=p�,=��+=K�*=��)=m)=�	(=�	'=�&= %=��#=��"=��!= � =W�=j�=7f=�?=�=I�=*�=fx=�:=��=M�=(e==�=c==�=64
=a�=�Q=4�=�[=	�=�S=���<�q�<xJ�<v�<V��<)��<XZ�<�<|��<W�<���<n��<��<8��<%�<���<4�<��<2�<n�<ֻ<I:�<���<w��<�R�<h��<^��<R�<���<�<	>�<d��<�ӏ<��<�d�<B��<Q�<Vtz<�s<��k<�d<~�\<j>U<3�M<XfF<	�><�7<%70<Y�(<�!<�*<�<��<�L<!�;���;P�;u �;���;;Wy�;�q�;�~�;�Bu;^�Y;�V>;�(#;�.;���:���:�b:�Y�9>��8A���=�9�n��]�����<�[>)�;�@�<bX��o��*���m��ш���|��fI��$�kĻ'�λ��ػ�����%���K �����o	�)�f��d��QS������#�`(��-,��=0�@4�!48��<���?���C��G��8K� �N���R�bV��Y�0&]�f�`��d�xg�:�j��0n�c�q���t�x��N{�φ~��܀�
s����������'�����D@��wɋ��P���֎��Z���ݑ��^���ޔ�^]���ڗ�jW���Қ�yM��!ǝ�2@��i���0��:����������	����������i���ޭ��S���Ȱ��=�������'�����|��Z�������&u��@콼�  �  ֏N=��M=TM=�ZL=o�K=��J=�!J=ecI=g�H=��G=�$G=dF=��E=��D= D=�ZC=8�B=�A=A=D@=4|?=@�>=2�====�Q<=��;=�:=��9=9=�?8=�j7=��6=U�5=d�4=�4=�(3=I2=g1=��0=��/=��.=]�-=k�,=��+=C�*=��)=o)=�	(=�	'=�&= %=��#=��"=��!=)� =Z�=l�=?f=�?=�=G�=.�=hx=�:=��=M�=)e==�=c=	=�=-4
=]�=�Q=/�=�[=�=|S=ߐ�<�q�<fJ�<o�<G��<!��<NZ�<�
�<���<W�<���<m��<��<8��< %�<���<@�<���<7�<+n�<"ֻ<Z:�<��<n��<�R�<e��<c��<R�<���<�<�=�<i��<�ӏ<��<�d�<9��<A�<tz<�s<\�k<�d<M�\<C>U<'�M<DfF<�><�7<*70<H�(<�!<�*<�<Đ<�L<P�;j��;AP�;� �;���;E��;ky�; r�;�;�Cu;��Y;�V>;P)#;�.;G��:׵�:�b:�V�9j��8Y�����9�R��������s=��>)�\�@��bX��o�+���m����� }��vI��D{kĻ`�λ��ػ��������D �����o	���N��A��DS������#�M(�-,��=0��?4�48��<���?���C�	�G��8K�$�N��R�uV��Y�O&]�r�`��d�xg�M�j��0n�~�q��t�x��N{�؆~��܀�s���������'�����=@��wɋ��P���֎��Z��wݑ��^���ޔ�Y]���ڗ�]W���Қ�mM��*ǝ�'@��m���0��6����������	��}�������i���ޭ��S���Ȱ��=�������'��
������m�������0u��:콼�  �  ϏN=��M=UM=�ZL=p�K=��J=�!J=fcI=p�H=��G=�$G=dF=��E=��D=�D=�ZC=2�B=�A=A=$D@=8|?=?�>=7�====�Q<=�;=�:=��9=9=�?8=�j7=��6=R�5=e�4=�4=�(3=
I2=g1=��0=��/=��.=\�-=f�,=��+=F�*=��)=l)=�	(=�	'=�&= %=��#=��"=��!=)� =_�=n�=Af=�?=�=F�=6�=hx=�:=��=I�=.e==�=c==�=*4
=`�=�Q=3�=�[= �=}S=Ր�<�q�<_J�<o�<=��<"��<QZ�<�<���<W�<���<k��<��<D��<"%�<���<3�<��<7�<=n�<ֻ<T:�<��<o��<�R�<g��<g��<R�<���<&�<>�<j��<xӏ<��<�d�<8��<E�<tz<�s<A�k<�d<C�\<F>U<+�M<*fF<�><Θ7<.70<K�(<�!<�*<��<Ԑ<�L<��;��;vP�;� �;���;���;dy�;4r�;�~�;�Cu;ܵY;.W>;�)#;�.;��:R��:b:�Y�9˹�8T�����9�+���������=��>)���@� cX���o�%+���m����� }��|I��gnkĻH�λ��ػ#�⻿�����@ �����o	���_��@��/S������#�`(�o-,��=0��?4�48��<���?���C��G��8K��N���R�}V�&�Y�W&]�a�`��d�xg�e�j�1n�v�q�-�t�x� O{�ֆ~��܀�s����������'�����2@��xɋ��P���֎��Z��uݑ��^���ޔ�Y]���ڗ�dW���Қ�^M��)ǝ�@��j���0��;����������	��{�������i���ޭ��S���Ȱ��=�������'��������k�������<u��:콼�  �  ӏN=��M=RM=�ZL=p�K=��J=�!J=gcI=j�H=��G=�$G=dF=ĢE=��D=D=�ZC=<�B=�A=A=&D@=3|?=B�>=7�==	==�Q<=�;=�:=��9=9=�?8=�j7={�6=S�5=_�4=�4=�(3=�H2=g1=�0=��/=��.=]�-=j�,=��+=F�*=��)=q)=�	(=
'=�&= %=��#=��"=��!=-� =b�=q�=Ef=�?=�=L�=3�=gx=�:=��=O�=(e==�=c=	=�=(4
=U�=�Q=(�=�[=��=uS=א�<�q�<_J�<j�<B��<��<DZ�< �<~��<W�<���<p��<��<F��<.%�<ģ�<G�<��<<�<<n�<,ֻ<g:�<��<|��<�R�<j��<p��<R�<���<�<�=�<\��<�ӏ<��<�d�<,��<8�<tz<us<>�k<�d<9�\<1>U<�M</fF<�><ޘ7<70<@�(<�!<�*<�<ܐ<�L<i�;���;�P�;� �;���;���;{y�;=r�;D�;�Cu;,�Y;^W>;W)#;	/;	��:K��:Qb:�Y�9E��87�����9�e��~������=�?)���@�cX�V�o�+���m��+���}��vI��F�kĻI�λ��ػ��⻨�����? �����o	���/��,��#S������#�2(�g-,��=0��?4�48��<�}�?���C�
�G��8K�>�N���R�sV�(�Y�]&]���`��d�0xg�l�j�"1n���q�%�t�=x��N{�܆~��܀�s��
�������'��	���2@��rɋ��P���֎��Z��oݑ��^���ޔ�T]���ڗ�SW���Қ�ZM��ǝ�@��h���0��1����������	����������i���ޭ��S���Ȱ��=�������'��������u�������9u��A콼�  �  ӏN=��M=XM=�ZL=n�K=��J=�!J=icI=m�H=��G=�$G=dF=ŢE=��D=D=�ZC=>�B=�A=A=)D@=7|?=E�>=,�==
==�Q<=�;=�:=��9=9=�?8=�j7=|�6=X�5=]�4=�4=�(3=�H2=g1=�0=��/=��.=S�-=k�,=��+=L�*=��)=p)=�	(=�	'=�&= %=��#=��"=��!=*� =c�=t�=Bf=�?=�=M�=2�=kx=�:=|�=N�=#e==	�=c=�=�=.4
=T�=�Q=!�=�[= �=pS=��<�q�<hJ�<W�<8��<��<LZ�<�<u��<W�<���<t��<��<H��<)%�<���<H�<��<A�<2n�<,ֻ<`:�< ��<���<�R�<o��<_��<R�<���<�<>�<\��<�ӏ<r�<�d�<3��<7�<tz<ds<]�k<�d<C�\<3>U<�M<FfF<��><ܘ7<70<W�(<�!<�*<�<��<�L<��;ү�;<P�;� �;���;h��;�y�;*r�;V�;�Cu;�Y;�W>;�)#;1/;���:o��:�b:bY�9:��8���û9�����������==�>?)���@��bX�ǃo��*���m������#}���I��@�kĻ�λ��ػ�������3 �����o	�	�<��;��S�}����#�<(��-,��=0��?4�48��<���?���C��G��8K�.�N��R��V�:�Y�E&]���`��d�Mxg�R�j�1n���q��t�=x��N{��~��܀�s���������'�����H@��oɋ��P���֎��Z��|ݑ��^���ޔ�O]���ڗ�SW���Қ�qM��ǝ�@��b���0��<����������	���������
j���ޭ��S���Ȱ��=�������'��������t�������.u��V콼�  �  ӏN=��M=RM=�ZL=p�K=��J=�!J=gcI=j�H=��G=�$G=dF=ĢE=��D=D=�ZC=<�B=�A=A=&D@=3|?=B�>=7�==	==�Q<=�;=�:=��9=9=�?8=�j7={�6=S�5=_�4=�4=�(3=�H2=g1=�0=��/=��.=]�-=j�,=��+=F�*=��)=q)=�	(=
'=�&= %=��#=��"=��!=-� =b�=q�=Ef=�?=�=L�=3�=gx=�:=��=O�=(e==�=c=	=�=(4
=U�=�Q=)�=�[=��=uS=ؐ�<�q�<_J�<k�<C��<��<DZ�<�<��<W�<���<p��<��<F��<.%�<ģ�<G�<��<<�<<n�<,ֻ<g:�<��<|��<�R�<j��<o��<R�<���<�<�=�<[��<�ӏ<��<�d�<,��<8�<tz<ts<>�k<�d<9�\<1>U<�M<0fF<�><ߘ7<70<@�(<�!<�*<�<ݐ<�L<j�;���;�P�;� �;���;���;{y�;=r�;D�;�Cu;*�Y;\W>;T)#;/;��:F��:Eb:{Y�9㰑8Q�����9�k���������=� ?)���@�cX�X�o�+���m��,���}��wI��F�kĻJ�λ��ػ��⻨�����? �����o	���0��,��#S������#�2(�g-,��=0��?4�48��<�}�?���C�
�G��8K�>�N���R�sV�(�Y�]&]���`��d�0xg�l�j�"1n���q�%�t�=x��N{�܆~��܀�s��
�������'��	���2@��rɋ��P���֎��Z��oݑ��^���ޔ�T]���ڗ�SW���Қ�ZM��ǝ�@��h���0��1����������	����������i���ޭ��S���Ȱ��=�������'��������u�������9u��A콼�  �  ϏN=��M=UM=�ZL=p�K=��J=�!J=fcI=p�H=��G=�$G=dF=��E=��D=�D=�ZC=2�B=�A=A=$D@=8|?=?�>=7�====�Q<=�;=�:=��9=9=�?8=�j7=��6=R�5=e�4=�4=�(3=
I2=g1=��0=��/=��.=\�-=f�,=��+=F�*=��)=l)=�	(=�	'=�&= %=��#=��"=��!=)� =_�=n�=Af=�?=�=F�=6�=hx=�:=��=I�=.e==�=c==�=*4
=a�=�Q=4�=�[= �=}S=Ր�<�q�<`J�<o�<>��<"��<RZ�<�<���<	W�<���<l��<��<D��<"%�<���<3�<��<7�<=n�<ֻ<T:�<��<o��<�R�<g��<g��<R�<���<%�<>�<j��<xӏ<��<�d�<8��<E�<tz<�s<A�k<�d<C�\<F>U<+�M<+fF<�><Θ7</70<L�(<�!<�*<��<Ԑ<�L<��;���;wP�;� �;���;���;dy�;3r�;�~�;�Cu;ٵY;+W>;�)#;�.;���:H��:�b:aY�9��8����Ż9�7���������=��>)���@�cX���o�'+���m�����!}��~I��hpkĻI�λ��ػ$��������@ �����o	���_��@��/S������#�`(�o-,��=0��?4�48��<���?���C��G��8K��N���R�}V�&�Y�W&]�a�`��d�xg�e�j�1n�v�q�-�t�x� O{�ֆ~��܀�s����������'�����2@��xɋ��P���֎��Z��uݑ��^���ޔ�Y]���ڗ�dW���Қ�^M��)ǝ�@��j���0��;����������	��{�������i���ޭ��S���Ȱ��=�������'��������k�������<u��:콼�  �  ֏N=��M=TM=�ZL=o�K=��J=�!J=ecI=g�H=��G=�$G=dF=��E=��D= D=�ZC=8�B=�A=A=D@=4|?=@�>=2�====�Q<=��;=�:=��9=9=�?8=�j7=��6=U�5=d�4=�4=�(3=I2=g1=��0=��/=��.=]�-=k�,=��+=C�*=��)=o)=�	(=�	'=�&= %=��#=��"=��!=)� =Z�=l�=?f=�?=�=G�=.�=hx=�:=��=M�=)e==�=c=	=�=-4
=]�=�Q=/�=�[=�=|S=���<�q�<gJ�<p�<H��<"��<OZ�<�
�<���<W�<���<m��<��<9��<!%�<���<@�<���<7�<+n�<"ֻ<Y:�<��<n��<�R�<e��<b��<
R�<���<�<�=�<h��<�ӏ<��<�d�<9��<A�<tz<�s<\�k<�d<N�\<D>U<(�M<EfF<�><�7<+70<I�(<�!<�*<�<Ő<�L<R�;k��;BP�;� �;���;E��;jy�;�q�;�;�Cu;��Y;�V>;J)#;�.;9��:ȵ�:�b:iV�9]��8������9�d��*������|=��>)�d�@��bX��o�+���m��
���}��yI��F|kĻa�λ��ػ��������E �����o	���O��A��DS������#�M(�-,��=0��?4�48��<���?���C�	�G��8K�$�N��R�uV��Y�O&]�r�`��d�xg�M�j��0n�~�q��t�x��N{�؆~��܀�s���������'�����=@��wɋ��P���֎��Z��wݑ��^���ޔ�Y]���ڗ�]W���Қ�mM��*ǝ�'@��m���0��6����������	��}�������i���ޭ��S���Ȱ��=�������'��
������m�������0u��:콼�  �  ۏN=��M=XM=�ZL=l�K=��J=�!J=gcI=a�H=��G=�$G=dF=��E=��D=�D=vZC=2�B=�A=A=D@=/|?=A�>=/�====�Q<=�;=�:=��9=9=�?8=�j7=��6=b�5=m�4=�4=�(3=I2=+g1=��0=��/=��.=`�-=p�,=��+=K�*=��)=m)=�	(=�	'=�&= %=��#=��"=��!= � =W�=j�=7f=�?=�=I�=*�=fx=�:=��=M�=(e==�=c==�=64
=b�=�Q=4�=�[=
�=�S=���<�q�<zJ�<w�<W��<+��<YZ�<�<}��<W�<���<o��<��<9��<%�<���<4�<��<2�<n�<ֻ<I:�<���<v��<�R�<h��<^��<R�<���<�<	>�<c��<�ӏ<��<�d�<A��<Q�<Vtz<�s<��k<�d<~�\<j>U<4�M<YfF<�><�7<&70<[�(<�!<�*<�<��<�L<$�;���;P�;v �;���;;Vy�;�q�;�~�;�Bu;Y�Y;�V>;�(#;�.;���:���:�b:vY�9���8����g�9����q�����<�e>)�D�@�EbX���o��*���m��Ո���|��iI��&�kĻ)�λ��ػ �����&���K �����o	�)�f��d��RS������#�`(��-,��=0�@4�!48��<���?���C��G��8K� �N���R�bV��Y�0&]�f�`��d�xg�:�j��0n�c�q���t�x��N{�φ~��܀�
s����������'�����D@��wɋ��P���֎��Z���ݑ��^���ޔ�^]���ڗ�jW���Қ�yM��!ǝ�2@��i���0��:����������	����������i���ޭ��S���Ȱ��=�������'�����|��Z�������&u��@콼�  �  ؏N=��M=XM=�ZL=o�K=��J=�!J=`cI=d�H=��G=�$G=dF=��E=��D=�D=vZC=1�B=�A=
A=D@=/|?=9�>=.�====�Q<=�;=�:=��9=	9=�?8=k7=��6=^�5=o�4=�4=�(3=I2="g1=�0=��/=��.=e�-=n�,=��+=J�*=��)=n)=�	(=�	'=�&=	 %=��#=��"=��!=� =R�=b�=5f=�?=�=?�=*�=ex=�:=��=M�=,e==�=c==�=>4
=g�=�Q=@�=\=�=�S=���<r�<�J�<��<T��<8��<]Z�<�<���<W�<���<`��<��<-��<%�<���<1�<��<�<n�<ֻ<B:�<<Z��<�R�<\��<Q��<R�<���< �<>�<q��<�ӏ<��<�d�<R��<O�<Btz<�s<��k<�d<x�\<e>U<[�M<{fF<'�><��7<C70<Z�(<�!<�*<�<��<rL<3�;��;�O�;_ �;p��;⓲;�x�;�q�;�~�;�Bu;�Y;(V>;�(#;5.;|��:��:#b:�W�9 ��8������9����g���P��	=�W>)���@��aX�Z�o��*��{m�������|��FI��4^kĻ7�λ��ػ!�����e���X ����p	�0�v��o��iS�͡���#�s(��-,�>0�@4�*48��<���?���C��G��8K��N��R�[V���Y�&]�V�`��d��wg��j��0n�Q�q���t�x��N{���~��܀��r����������'�����A@���ɋ��P���֎��Z���ݑ��^���ޔ�s]���ڗ�nW���Қ��M��>ǝ�,@��u���*0��;����������	��t�������i���ޭ��S���Ȱ��=�������'���������]�������u��2콼�  �  ؏N=��M=YM=�ZL=k�K=��J=�!J=XcI=b�H=��G=�$G=dF=��E=��D=�D=sZC=&�B=�A=A=D@=.|?=2�>=0�==�==�Q<=�;=�:=��9=9=�?8=�j7=��6=h�5=y�4=�4=�(3=I2=*g1=�0=��/=��.=m�-=p�,=��+=F�*=��)=h)=�	(=�	'=�&= %=��#=��"=��!=� =J�=Z�=5f=�?=�=9�=&�=cx=�:=��=G�=,e==�=c==#�==4
=r�=�Q=L�=\=�=�S=��<!r�<�J�<��<_��<>��<fZ�<�<���<W�<���<W��<��<#��<%�<���<�<��<
�<n�<ֻ<3:�<ꚴ<L��<�R�<I��<X��<R�<���<�<>�<x��<�ӏ<��<�d�<W��<e�<dtz<�s<��k<d<��\<�>U<m�M<nfF<O�><��7<T70<_�(<�!<�*<��<��<OL<#�;��;�O�;  �;,��;���;�x�;uq�;s~�;EBu;��Y;�U>;�(#;�-;���:U��:{b:�V�9���8����j�9���T���p��<��=)�k�@�bX���o��*��+m�������|��I��.>kĻZ�λ��ػT�����[���n ����<p	�<����z���S����#��(��-,�1>0�%@4�548��<���?���C��G��8K� �N�ۂR�>V��Y�&]�0�`��d��wg��j��0n�'�q���t��x��N{���~��܀��r����������'�����=@���ɋ��P���֎��Z���ݑ��^���ޔ��]��ۗ�zW���Қ��M��Kǝ�3@������#0��>����������	��m�������i���ޭ��S���Ȱ��=��w����'��㜶�p��J���w���u��콼�  �  ��N=��M=\M=�ZL=l�K=��J=�!J=WcI=Y�H=��G=�$G=�cF=��E=��D=�D=iZC=�B=��A=A=D@=&|?=2�>=-�====�Q<=�;=�:=��9=9=�?8=k7=��6=o�5=~�4=�4=�(3=I2=5g1=�0=��/=ų.=n�-=s�,=��+=L�*=��)=j)=�	(=�	'=�&=��$=��#=��"=��!=� =F�=Y�=+f=�?=�=>�="�=]x=�:=��=L�=/e==�=c==)�=E4
=v�=�Q=N�=\=#�=�S=��<)r�<�J�<��<n��<;��<iZ�<�<���<W�<���<X��<��<"��<	%�<���<�<Α�<�<�m�<�ջ< :�<ܚ�<W��<�R�<G��<T��<�Q�<���<"�<>�<r��<�ӏ<��<�d�<`��<r�<�tz<�s<��k<-d<��\<�>U<}�M<�fF<V�><�7<G70<k�(<�!<�*<��<��<ML<��;��;�O�;���;���;l��;�x�;q�;*~�;{Au;h�Y;�U>;(#;�-;��:���:b:�W�9k��8ކ����9��������M��!<��=)��@��aX���o�I*��m�������|��
I��RkĻ,�λ��ػH�����i���� ���$p	�d��������S����.�#��(��-,�!>0�8@4�P48��<���?���C��G��8K��N�ՂR�7V�ۣY�&]�'�`��d��wg���j��0n��q���t��x��N{���~�s܀�s����������'�����E@���ɋ�Q���֎��Z���ݑ��^���ޔ��]��ۗ��W��Ӛ��M��@ǝ�C@������&0��B����������	��r�������i���ޭ��S���Ȱ�o=��q����'��ۜ��_��<���p���u��콼�  �  �N=��M=^M=�ZL=l�K=��J=�!J=[cI=R�H=��G=�$G=�cF=��E=��D=�D=_ZC=%�B=��A=�
A=D@=|?=4�>=&�====�Q<=�;=�:=��9=9=�?8=k7=��6=s�5=��4=�4=�(3=I2=8g1=�0=��/=ʳ.=o�-={�,=��+=N�*=��)=m)=�	(=�	'=�&=��$=��#=��"=��!=� =?�=Q�="f=�?=�=7�=�=]x=�:=��=O�=,e="=�=c=!=.�=P4
=x�=�Q=R�=\=(�=�S=*��<0r�<�J�<��<x��<L��<gZ�<�<���<W�<���<]��<��<��<�$�<���<�<���<�<�m�<�ջ<':�<̚�<E��<�R�<N��<E��<�Q�<���<�<>�<u��<�ӏ<��<�d�<k��<s�<�tz<�s<�k<0d<ŭ\<�>U<��M<�fF<O�><7�7<T70<t�(<�!<�*<��<��<\L<��;���;YO�;���;���;��;qx�;�p�;Y~�;xAu;۳Y;CU>;�'#;�-;��:z��:�b:zV�9W��8部�{�9�B����������;�m=)��@��`X���o�:*��"m��Q���{|��I����ikĻ�λ��ػ1���컉���{ �&��Gp	�{��������S���T�#��(��-,�?>0�J@4�Q48��<���?���C��G��8K��N���R�/V�ϣY��%]�#�`�sd��wg���j��0n��q���t��x�|N{���~�k܀��r����������'�����Q@���ɋ�Q���֎�[���ݑ��^���ޔ��]��&ۗ��W��Ӛ��M��Rǝ�P@������50��D����������	��o�������i���ޭ��S���Ȱ�l=��p���v'��ڜ��\��9���h����t�� 콼�  �  �N=��M=_M=�ZL=h�K=��J=�!J=UcI=T�H=��G=�$G=�cF=��E=��D=�D=]ZC=�B=��A=�
A=D@=|?=/�>=(�==�==�Q<=�;=�:=��9=9=�?8=k7=��6=z�5=��4=�4=�(3=)I2=>g1=�0=��/=̳.=s�-=}�,=��+=O�*=��)=e)=�	(=�	'=�&=��$=��#=��"=��!=� ==�=N�=f=�?=�=/�=�=Xx=�:=��=H�=/e=$=�= c=%=2�=Q4
=��=�Q=\�=\=.�=�S=9��<Dr�<�J�<��<{��<T��<oZ�<�<���<W�<���<T��<��<��<�$�<x��<��<���<��<�m�<�ջ<:�<̚�<8��<�R�<A��<D��<�Q�<x��<"�<>�<z��<�ӏ<��<�d�<r��<��<�tz<*s<�k<]d<ܭ\<�>U<��M<�fF<i�><3�7<b70<|�(<�!<�*<��<��<DL<��;���;IO�;���;���;��;*x�;�p�;�}�;�@u;��Y;�T>;�'#;H-;&��:|��:2b:]W�9r��8����*�9��������C��;�=)���@��`X��o�*���l��J���p|���H����PkĻ�λ��ػs��#�컭���� �1��hp	�w��������S�%��g�#��(�.,�`>0�U@4�h48�<���?���C�	�G��8K��N���R�#V���Y��%]��`�_d��wg���j��0n��q���t��x��N{���~�k܀��r����������'��%���M@���ɋ�Q���֎�[���ݑ� _���ޔ��]��+ۗ��W��Ӛ��M��^ǝ�N@������60��K����������	��j�������i���ޭ��S��tȰ�`=��Y���s'��Ĝ��Q��#���]����t��콼�  �  �N=��M=ZM=�ZL=m�K=��J=�!J=OcI=T�H=��G=�$G=�cF=��E=��D=�D=bZC=�B=��A=�
A=D@= |?=)�>=)�==�==�Q<=�;=�:=��9=9=�?8=k7=��6=w�5=��4=�4=�(3=-I2=8g1=�0=��/=ҳ.=t�-=|�,=��+=K�*=��)=i)=�	(=�	'=�&=��$=��#=��"=��!=
� =8�=I�=#f=�?=�=.�=�=Vx=�:=��=L�=6e=!=!�=!c='=;�=Q4
=��=�Q=`�= \=5�=�S=2��<Tr�<�J�<��<~��<U��<rZ�<�<���<W�<���<K��<��<��<�$�<��<��<���<��<�m�<�ջ<
:�<Κ�<-��<�R�<6��<H��<�Q�<���<*�<	>�<���<�ӏ<��<�d�<z��<��<�tz<Es<�k<d<̭\<�>U<��M<�fF<��><7�7<q70<i�(<�!<�*<��<��<)L<��;^��;NO�;���;w��;��;�w�;�p�;�}�;Au;j�Y;�T>;�'#;�,;5��:���:+b:�V�9���8
�����9�j������[���;�6=)��@��`X�Ȁo�A*���l��N���@|���H����%kĻA�λ��ػY���컫���� �3��qp	�m�������S�<��T�#��(��-,�g>0�_@4�s48�<���?���C��G��8K���N���R� V���Y��%]���`�td�|wg���j�h0n��q���t��x��N{�X�~�i܀��r����������'�����L@���ɋ�Q���֎�[���ݑ�
_���ޔ��]��/ۗ��W��#Ӛ��M��jǝ�M@������20��I����������	��_�������i���ޭ��S��vȰ�k=��L���w'������Z��&���S����t��콼�  �  �N=��M=bM=�ZL=k�K=��J=�!J=ScI=Q�H=��G=�$G=�cF=��E=��D=�D=VZC=�B=��A=�
A=D@=|?=.�>="�==�==�Q<=�;=�:=��9=9=�?8=k7=��6=��5=��4=�4=�(3=0I2=Cg1="�0=��/=ӳ.=q�-=�,=��+=R�*=��)=j)=�	(=�	'=�&=��$=��#=��"=��!=� =5�=G�=f=�?=�=-�=�=Zx=�:={�=L�=0e='="�=$c=&=9�=X4
=��=�Q=e�=#\=8�=�S=K��<Yr�<�J�<��<���<_��<yZ�<!�<���<W�<���<U��<��<��<�$�<p��<��<���<��<�m�<�ջ<
:�<���<.��<�R�<=��<=��<�Q�<���<$�<>�<���<�ӏ<��<�d�<���<��<�tz<Gs<��k<}d<�\<�>U<��M<�fF<s�><=�7<w70<��(<�!<�*<��<��<:L<��;k��;O�;f��;^��;���;�w�;rp�;�}�;�@u;�Y;�T>;f'#;%-;(��:u��:b:�W�9̽�8#���Ʒ9�E������1��;��<)��@��`X���o��)���l�����?|���H����%kĻ�λ��ػU��I�컷���� �9��rp	���������S�C��{�#��(�#.,�l>0�b@4�f48�<���?���C��G��8K���N���R�&V���Y��%]�֞`�Hd�mwg���j�^0n�ہq�m�t��x�qN{�q�~�h܀��r����������'�� ���\@���ɋ�Q���֎�[���ݑ�_���ޔ��]��<ۗ��W��#Ӛ��M��hǝ�R@������=0��R����������	��_�������i���ޭ��S��lȰ�X=��L���r'������G�����O����t��콼�  �  '�N=��M=M=�`L=��K=��J=z*J=�lI=��H=��G=�0G=�pF=+�E=�D=6-D=�jC=T�B=(�A=2A=NX@=w�?=��>=� >=�6==�k<= �;=r�:=j:=�19=`8=��7=��6=��5=Q5=�-4=�Q3=ms2=�1=��0=��/=c�.=��-=N-==,=h-+=�8*=�@)=�E(=�G'=�E&=�@%=�7$=c+#="=�!=;�=��=��=J�=da=�2=��=��=�=&I=f=��=�e=�=��=�T=6�=Ԅ
=r	=�=�'=v�=k&=��=P =��<0��<���<di�<�%�<%��<��<�,�<��<�b�<2��<3�<Z�<��<��<Hs�<���<zO�<��<��<sz�<�ִ< 0�<��<�٩<0*�<�x�<�Ğ<P�<X�<O��<Z�<C*�<Vn�<���<��<�nz<�r<�yk<��c<5�\<U<��M<�'F<�><�I7<r�/<Jy(<B!<��<�a<<x�<���;y�;��;��;gX�;��;��;<֔;ӆ;�q;mV;�:;�P;[8;��:Q�:�P:�9ߙ�44�͹�L����ٍʺ����7J��].�<%F�Y�]���t�Յ�����:��&1������F���!ǻuѻR�ۻ���a��\6��@b�����
��F�@��>.����� �.	%��1)��J-��T1�
P5�S=9�F=�9�@���D��pH��L�?�O�\S���V��oZ�C�]��]a���d��)h�g�k���n��!r�
fu�n�x���{������ձ��?C��R҅�C_��ꈼ�r������8������������؄��������V����u���xh��i����W��7Π�QD��ι���.���������틩�����^s���歼rZ���Ͱ�cA�������(���������;������Ko���佼�  �  '�N=��M=M= aL=��K=��J=w*J=�lI=��H=��G=�0G=�pF=,�E=�D=3-D=�jC=T�B=0�A=3A=OX@=s�?=��>=� >=�6==�k<=$�;=u�:=o:=�19=`8=��7=��6=��5=S5=�-4=�Q3=rs2=�1=��0=��/=c�.=��-=P-=D,=g-+=�8*=�@)=�E(=�G'=�E&=�@%=�7$=h+#=	"=�!=;�=��=��=L�=ja=�2=��=��=�="I=_=��=�e=�=��=T=6�=ׄ
=p	=�=�'=m�=g&=��=H =��<*��<���<di�<�%�</��<��<�,�<��<�b�<��<'�<]�<��<��<Es�<���<vO�<��<��<�z�<�ִ<�/�<��<_٩<%*�<�x�<�Ğ<Z�<X�<\��<Z�<>*�<Sn�<���<��<�nz<�r<�yk<��c<<�\<U<��M<�'F<��><�I7<��/<Ly(<S!<��<�a<<9�<���;y�;��;G��;lX�;�;l�;Q֔;ӆ;{�q;�V;��:;�P;]7;ϧ�:�P�:��P:��9/5t�͹��L�Q���6�ʺ�����J��].�B%F��]�N�t�%Յ�����:��$1��
���0���� ǻ uѻ.�ۻ*��w�ﻤ6��xb�|���
��F�3��0.����� �	%��1)��J-��T1��O5�~=9�p=�E�@���D��pH��L�&�O�\S���V��oZ�7�]��]a���d�)h���k�	�n�u!r�-fu�n�x���{������˱��5C��L҅�>_��ꈼ�r������D������������ۄ��������S����u���lh��n����W��XΠ�\D��Թ���.���������ߋ������cs���歼hZ���Ͱ�bA�������(���������C������No���佼�  �   �N=��M=M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=,�E=�D=4-D=�jC=S�B=4�A=2A=SX@=|�?=��>=� >=�6==�k<= �;=l�:=g:=�19=`8=��7=��6=��5=T5=�-4=�Q3=ts2=�1=z�0=��/=`�.=��-=I-==,=_-+=�8*=�@)=�E(=�G'=�E&=�@%=�7$=l+#="=�!=>�=��=��=J�=oa=�2=��=��=�=+I=a=��=�e=�=��={T=2�=҄
=k	=��=�'=g�=e&=��=C =��<!��<��<Yi�<�%�<��<���<�,�<��<�b�<��<:�<i�<��<(��<Ds�<���<yO�<��<��<�z�<�ִ<�/�<&��<e٩<8*�<�x�<�Ğ<[�<X�<O��<L�<>*�<Ln�<���<��<�nz<&�r<ryk<��c<2�\<�U<��M<s'F<��><yI7<n�/<'y(<P!<��<�a<%<B�<0��;y�;��;_��;nX�;:�;w�;|֔;ӆ;��q;{V;A�:;eQ;�7;��:�P�:A�P:]�9H��4K�͹͛L�)���|�ʺm����J��].�@%F���]�$�t�/Յ����:��<1�����f���!ǻauѻ�ۻ��:��Q6��ab�T���
�xF�9��-.����� �	%��1)�J-��T1��O5�`=9�J=�#�@���D��pH��L�F�O�/\S���V��oZ�I�]��]a���d�v)h���k��n�k!r�;fu�m�x���{������ޱ��IC��[҅�:_��ꈼ�r������0������������܄��������H����u���jh��p����W��RΠ�ID��ι���.���������싩�����cs���歼kZ���Ͱ�hA��𴳼�(���������M������Uo���佼�  �  "�N=��M=M=�`L=��K=��J=z*J=�lI=��H=��G=�0G=�pF=0�E=�D==-D=�jC=Y�B=7�A=<A=VX@=y�?=��>=� >=�6==�k<="�;=v�:=j:=�19=`8=��7=��6=��5=H5=�-4=�Q3=bs2=	�1=v�0=��/=[�.=��-=I-=A,=h-+=�8*=�@)=�E(=�G'=�E&=�@%=�7$=q+#="=�!=G�=��=��=P�=qa=�2=��=��=�= I=d=��=�e=�=��={T=,�=΄
=e	=��=�'=g�=^&=��=D =��<��<��<Zi�<�%�<)��<��<�,�<��<�b�<#��<4�<h�<���<,��<Qs�<���<�O�<��<��<�z�<�ִ<0�<��<o٩<0*�<�x�<�Ğ<X�<X�<T��<M�<:*�<En�<���<��<�nz<��r<�yk<��c<�\<�U<}�M<f'F<�><}I7<v�/<Ty(<I!<�<�a<<W�<��;Ty�;	�;���;�X�;X�;��;�֔;7ӆ;�q;,V;��:;7Q;8;3��:�P�:��P:��915b�͹�L�������ʺo����J�e^.��%F�.�]�5�t�7Յ�4��;��]1�����d���� ǻuѻ2�ۻ���{��Z6��Ub�i���
�bF�$��.������ �		%��1)�rJ-�dT1��O5�`=9�G=�J�@���D��pH��L�-�O�*\S���V��oZ�U�]��]a���d��)h���k�%�n��!r�5fu���x���{�����ױ��6C��S҅�=_��ꈼ�r������5�����䄐����΄��������=����u���\h��Z����W��HΠ�QD��׹���.���������狩�����hs���歼xZ���Ͱ�sA������(���������M���'���[o��彼�  �  �N=��M=
M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=9�E=�D=D-D=�jC=a�B=:�A=?A=[X@=z�?=��>=� >=�6==�k<=�;=o�:=b:=�19=`8=��7=��6=��5=D5=�-4=�Q3=\s2=�1=n�0=��/=U�.=��-=E-=:,=d-+=�8*=�@)=�E(=�G'=�E&=�@%=�7$=q+#="=�!=H�=��=��=Z�=qa=�2=��=��=�=#I=h=��=�e=�=��=sT=#�=̈́
=Y	=��=�'=`�=U&=��=< =��<��<Ѥ�<Mi�<�%�<��<���<�,�<"��<�b�<1��<6�<o�<��<-��<cs�<���<�O�<!��<��<�z�<�ִ<0�<��<٩<<*�<�x�<�Ğ<O�<X�<F��<H�<&*�<An�<���<��<�nz<��r<uyk<��c<�\<�U<g�M<d'F<ɶ><qI7<V�/<<y(<7!<�<�a<#<{�<��;�y�;+	�;���;�X�;x�;�;�֔;�ӆ;E�q;oV;�:;dQ;�8;Ȩ�:�Q�:\�P:��9~g�4˅͹"�L�Ǵ��_�ʺ(���K��^.�&F�\�]���t�JՅ�p���:���1��P������'!ǻ*uѻM�ۻϤ�N��'6��Ab�^�{�
�aF����.������ ��%�W1)�oJ-�KT1��O5�Q=9�-=�9�@�u�D��pH��L�K�O�<\S���V��oZ�R�]�^a���d��)h���k�A�n��!r�Kfu���x���{�7���求�FC��W҅�<_���鈼�r������2�����ڄ���������������:����u���\h��P����W��9Π�ED��ʹ���.�����������������zs���歼Z���Ͱ�tA�� ����(��ǜ�����[���1���[o��彼�  �  �N=��M=M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=?�E=�D=I-D=�jC=g�B=G�A=?A=_X@=��?=��>=� >=�6==�k<= �;=n�:=e:=�19=`8=��7=��6=��5=?5=�-4=�Q3=^s2=��1=i�0=��/=R�.=��-=E-=<,=_-+=�8*=�@)=�E(=�G'=�E&=�@%=�7$={+#="=�!=S�=��=��=]�=}a=�2=��=��=��=&I=^=��=�e=�=��=pT=�=Ä
=V	=�=�'=O�=J&=��=+ =��< ��<ˤ�<Gi�<�%�<��<���<�,�<��<�b�<+��<I�<z�<���<H��<ls�<���<�O�<:��<��<�z�< ״<0�<=��<~٩<A*�<�x�<�Ğ<]�<X�<K��<B�<&*�<5n�<���<~�<hnz<��r<?yk<��c<چ\<�U<X�M<C'F<Ƕ><aI7<^�/<-y(<J!<��<�a<0<y�<���;�y�;S	�;��;Y�;��;6�;)ה;�ӆ;8�q;�V;<�:;NR;�8;���:�P�:��P:N�9�
 5u�͹��L�������ʺ����K��^.�n&F�G�]�\�t��Յ����-;���1��R���x���!ǻMuѻ��ۻ��I��,6��;b�#���
�2F�����-����]� ��%�G1)�<J-�VT1��O5�@=9�5=�)�@���D��pH��L�F�O�8\S���V��oZ�q�]�^a��d��)h��k�g�n��!r��fu���x���{�=���᱂�HC��Z҅�7_��ꈼ�r�����������݄��k���������u��!����u��tNh��Q����W��;Π�BD��չ���.���������񋩼����{s��筼�Z��ΰ��A������(��ʜ�����u���8���jo��彼�  �  �N=��M=M= aL=��K=��J=�*J=�lI=��H=��G=�0G=�pF=A�E=)�D=N-D=�jC=h�B=S�A=MA=bX@=��?=��>=� >=�6==�k<=�;=k�:=c:=�19=`8=��7=��6=��5=25=�-4=�Q3=Ts2=�1=m�0=��/=L�.=��-=:-=<,=Z-+=�8*=�@)=�E(=�G'=�E&=�@%=�7$=�+#="=�!=Z�=��=ð=^�=�a=�2=��=��=�=-I=]=��=�e=�=��=dT=�=��
=X	=ڠ=�'=H�=D&=��=! =��<���<Ĥ�<*i�<�%�<��<��<�,�<��<�b�<&��<L�<�<��<c��<ls�<���<�O�<P��<��<�z�<$״<0�<G��<~٩<N*�<�x�<�Ğ<c�<X�<O��<+�<*�< n�<���<��<4nz<��r<yk<z�c<��\<�U<J�M<'F<��><.I7<`�/<y(<M!<�<�a<L<s�<���;�y�;�	�;N��;4Y�;F�;d�;�ה;�ӆ;�q;xV;��:;�R;�8;���:�Q�:��P:��9z��4��͹�L�{����ʺ����*L��_.��&F���]���t�օ�k���;���1������Ǥ��!ǻsuѻʠۻ����6��/b��m�
��E�����-�j��E� ��%�@1)��I-�8T1��O5�3=9�,=�
�@���D��pH��L�C�O�]\S��V�pZ���]��]a�J�d��)h���k�x�n��!r��fu���x��{�D���豂�JC��a҅�'_��ꈼ�r�����������Ƅ��O���������l������u��k*h��L����W��;Π�6D��ȹ���.��������������s��筼�Z��ΰ��A��-����(��֜����s���=����o��彼�  �  �N=��M=�M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=N�E=/�D=V-D=�jC=t�B=O�A=TA=lX@=��?=��>=� >=�6==�k<=�;=d�:=]:=�19=`8=��7=q�6=��5=-5=�-4=�Q3=Js2=�1=^�0=|�/=H�.=��-=;-=5,=Z-+=�8*=�@)=�E(=�G'=�E&=�@%=8$=�+#=%"=�!=^�=��=ΰ=h�=�a=
3=��=��=��=*I=`=��=�e=�=��=_T=�=��
=E	=נ={'=A�=9&=x�= =u�<���<���<!i�<�%�<���<��<�,�<��<�b�<9��<V�<��<&��<Z��<�s�<���<�O�<Z��<��<�z�<"״<70�<I��<�٩<P*�<�x�<�Ğ<W�<�W�<?��<0�<*�<n�<n��<o�<.nz<t�r<yk<H�c<��\<zU<�M<'F<��><5I7<C�/<	y(<:!<�<�a<J<��<���;z�;�	�;V��;�Y�;|�;��;�ה;?Ԇ;��q;V;E�:;�R;j9;���:OR�:K�P:B�9���4��͹��L�Ĵ���ʺ����LL��_.�;'F�ء]���t�
օ�����;���1����������@!ǻnuѻ�ۻ�����5���a��6�
��E�����-�X��2� �%�1)�J-�T1��O5�=9�=��@���D��pH��L�a�O�a\S�(�V�pZ���]�B^a�O�d� *h��k���n�"r��fu��x��{�M�$��󱂼YC��e҅�1_��ꈼ�r���������������W���������\������u��c,h��5����W�� Π�3D�������.������������������s��$筼�Z��ΰ��A��E���)��휶�������^����o��$彼�  �  �N=��M=M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=X�E=1�D=d-D=�jC=��B=Y�A=YA=qX@=��?=��>=� >=�6==�k<=#�;=h�:=\:=�19=�_8=��7=i�6=��5=(5=�-4=�Q3=?s2=�1=P�0=�/=A�.=��-==-=/,=c-+=�8*=�@)=�E(=�G'=�E&=�@%=8$=�+#=4"=�!=i�=��=Ͱ=v�=�a=3=��=��=��=)I=c=��=�e=�=��=XT=	�=��
=6	=Ѡ=p'=5�=+&=p�= =\�<���<���<i�<~%�<���<���<y,�<��<�b�<7��<V�<��<3��<g��<�s�<���<�O�<d��<��<�z�<%״<M0�<G��<�٩<J*�<�x�<�Ğ<[�<X�<4��<2�<�)�<n�<l��<T�<nz<C�r<�xk<�c<��\<JU<��M<'F<i�><6I7<1�/<)y(<H!<��<�a<?<��<���;Oz�;
�;̩�;�Y�;��;)�;�ה;�Ԇ;��q;vV;��:;S;�9;Ϊ�:S�:��P:Y�9�;�4~�͹>�L�����ϐʺ�����L�`.��'F�L�]��t�'օ�F���;��2����������m!ǻ#uѻ'�ۻ̤�����5���a���
��E�y���-�*���� ��%��0)�J-��S1��O5�=9�=��@�v�D��pH��L�u�O�W\S�=�V�7pZ���]�x^a�^�d�C*h�;�k���n�)"r��fu��x��{���$��򱂼WC��S҅�C_���鈼�r������
���������I��}������=�������u��F*h������W��Π�:D�������.�����������������s��(筼�Z��8ΰ��A��\���)�����#������d����o��C彼�  �  
�N=��M=�M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=Z�E=:�D=i-D=�jC=��B=`�A=\A=sX@=��?=��>=� >=�6==�k<=�;=b�:=V:=�19=�_8=~�7=i�6=��5= 5=�-4=�Q3=;s2=ܒ1=O�0=y�/==�.=��-=6-=+,=]-+=�8*=�@)=�E(=�G'=�E&=�@%=8$=�+#=9"=�!=o�=��=Ѱ=z�=�a=3=��=��=��=0I=e=��=�e=�=��=TT=�=��
=4	=Ơ=i'=1�=(&=g�=	 =Z�<���<���<i�<p%�<���<��<�,�<!��<�b�<>��<h�<��<3��<w��<�s�<���<�O�<t��<�<�z�<1״<L0�<]��<�٩<Z*�<�x�<�Ğ<V�<�W�<,��<#�<�)�<n�<h��<N�<�mz<2�r<�xk<�c<^�\<6U<�M<�&F<f�><I7<�/<y(<8!<	�<b<^<��<��;Kz�;9
�;
��;Z�;��;W�;'ؔ;�Ԇ;�q;�V;�:;�S;�9;��:�S�:1�P:O�9���4��͹��L�����G�ʺ����9M�v`.��'F���]�V�t�qօ�G���;��-2������ؤ���!ǻQuѻ�ۻ��廵�ﻯ5���a����
��E�c��z-����� �l%��0)��I-��S1�mO5��<9��=���@�h�D��pH��L���O�r\S�I�V�GpZ���]�z^a���d�W*h�H�k���n�D"r��fu��x�,�{���/������bC��]҅�:_���鈼�r�������~���������9��x���z��6�������u��9h��!���oW��Π�*D�������.�����������������s��3筼�Z��>ΰ��A��e���)�����4������g����o��C彼�  �  �N=��M= M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=b�E=E�D=b-D=�jC=��B=b�A=bA=xX@=��?=��>=� >=�6==�k<=�;=g�:=Y:=�19=�_8=s�7=b�6=��5=5=�-4=|Q3=8s2=֒1=M�0=p�/=>�.=��-=2-=5,=[-+=�8*=�@)=�E(=�G'=�E&=�@%=8$=�+#=7"=�!=s�=��=�=y�=�a=3=��=��=��=(I=\=��=�e=�=��=ST=�=��
=0	=��=d'=%�=&=b�= =L�<���<���<i�<r%�<���<���<�,�<��<�b�<<��<i�<��<;��<|��<�s�<��<�O�<���<�<�z�<D״<P0�<f��<�٩<V*�<�x�<�Ğ<U�< X�<<��<�<*�<�m�<T��<F�<�mz<&�r<�xk<��c<H�\<$U<ΙM<�&F<|�><�H7<5�/<y(<4!<�<�a<U<��<*��;fz�;�
�;��;UZ�;B�;)�;�ؔ;�Ԇ;I�q; V;?�:;�S;�9;���:�R�:�P:R�9� 5��͹��L�ǵ����ʺ@���eM��`.�R(F��]�y�t��օ�R��(<��2����������5!ǻYuѻ�ۻ������5���a����
��E�i��8-������ �#%��0)��I-��S1�[O5��<9�=��@���D��pH��L�\�O�z\S�F�V�6pZ���]��^a���d�g*h�p�k���n�U"r�gu�-�x�X�{�}�6������SC��d҅�4_��ꈼ�r�������~���������3��s���X��A������~u��<h�����fW��Π�/D��Ĺ���.�����������������s��=筼�Z��Eΰ��A��j���,)�����?������w����o��8彼�  �  �N=��M=�M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=d�E=D�D=k-D=�jC=��B=h�A=cA={X@=��?=��>=� >=�6==�k<=�;=c�:=P:=�19=�_8=t�7=a�6=��5=5=�-4=yQ3=4s2=֒1=G�0=q�/=6�.={�-=,-=+,=Y-+=�8*=�@)=�E(=�G'=�E&=�@%=8$=�+#=;"=�!=t�=��=�={�=�a=3=��=��= �=0I=d=��=�e=�=��=KT=��=��
=*	=��=b'=#�=&=`�= =E�<���<���<�h�<\%�<���<݆�<,�<��<�b�<J��<i�<��<@��<���<�s�<��<�O�<���<�<�z�<D״<V0�<e��<�٩<g*�<�x�< Ş<R�< X�<*��<�<�)�<�m�<V��<>�<�mz<�r<�xk<��c<I�\<U<ЙM<�&F<S�><�H7<�/<	y(</!<�<�a<u<��<&��;�z�;�
�;.��;gZ�;>�;r�;�ؔ;Ն;��q;> V;z�:;�S;y:;���:�S�:��P:Q�9l6�4I�͹M�L����n�ʺ_���dM��`.��(F�6�]���t��օ���<��Y2�� ��%����!ǻkuѻ�ۻ��廪��u5���a�����
��E�Z��B-������ �.%��0)��I-��S1�PO5��<9��=���@�g�D��pH��L���O��\S�f�V�ZpZ���]��^a���d�n*h�y�k� �n�Y"r��fu�8�x�V�{���?�����`C��f҅�9_���鈼�r�������~���������'��n���]��1������~u��4h�����gW��Π�D�������.�����������������s��B筼�Z��Lΰ��A��u���-)�����>������v����o��L彼�  �  �N=��M=M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=b�E=B�D=y-D=�jC=��B=j�A=_A=|X@=��?=��>=� >=�6==�k<=�;=f�:=V:=�19=�_8=w�7=[�6=��5=5=�-4=zQ3=1s2=ג1=A�0=q�/=4�.=��-=;-=-,=_-+=�8*=�@)=�E(=�G'=�E&=�@%=8$=�+#=B"=�!=y�=��=۰=��=�a=3=��=��=��=*I=d=��=�e=�=��=TT=��=��
=%	=��=^'=#�=&=]�=� =:�<���<���<i�<m%�<���<��<v,�<��<�b�<H��<n�<��<7��<���<�s�<��< P�<���<�<�z�<?״<Z0�<j��<�٩<Z*�<�x�<�Ğ<O�<X�<+��<0�<�)�<�m�<Q��<0�<�mz<�r<�xk<��c<H�\<�U<��M<�&F<X�></I7<�/<y(<.!< �<�a<\<��<:��;�z�;o
�;^��;XZ�;,�;��;uؔ;Ն;��q;�V;��:;!T;s:;���:�S�:��P:��9h��4�͹D�L�����ʺ%����M��`.��(F��]���t��օ����<��k2����������m!ǻ:uѻ6�ۻ���؀ﻜ5���a����
��E�:��U-����� �B%��0)��I-��S1�QO5��<9��=��@�g�D��pH��L�t�O�l\S�@�V�fpZ���]��^a���d�{*h�v�k� �n�f"r�gu�N�x�I�{���������[C��\҅�B_���鈼�r�������~���������#��j���g���������u��%h�����bW��Π�*D�������.�����������������s��D筼�Z��[ΰ��A��{���')��%���>����������o��J彼�  �  �N=��M=�M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=d�E=D�D=k-D=�jC=��B=h�A=cA={X@=��?=��>=� >=�6==�k<=�;=c�:=P:=�19=�_8=t�7=a�6=��5=5=�-4=yQ3=4s2=֒1=G�0=q�/=6�.={�-=,-=+,=Y-+=�8*=�@)=�E(=�G'=�E&=�@%=8$=�+#=;"=�!=t�=��=�={�=�a=3=��=��= �=0I=d=��=�e=�=��=KT=��=��
=*	=��=b'=#�=&=a�= =E�<���<���<�h�<]%�<���<݆�<,�<��<�b�<K��<j�<��<A��<���<�s�<��<�O�<���<�<�z�<D״<V0�<e��<�٩<f*�<�x�< Ş<Q�< X�<*��<�<�)�<�m�<V��<>�<�mz<�r<�xk<��c<I�\<U<љM<�&F<S�><�H7<�/<	y(</!<�<�a<v<��<'��;�z�;�
�;/��;hZ�;>�;r�;�ؔ;Ն;��q;; V;w�:;�S;v:;���:�S�:��P:1�9��4j�͹^�L����v�ʺg���hM��`.��(F�:�]���t��օ���� <��Z2�� ��&����!ǻkuѻ�ۻ��廫��u5���a�����
��E�Z��B-������ �.%��0)��I-��S1�PO5��<9��=���@�g�D��pH��L���O��\S�f�V�ZpZ���]��^a���d�n*h�y�k� �n�Y"r��fu�8�x�U�{���?�����`C��f҅�9_���鈼�r�������~���������'��n���]��1������~u��4h�����gW��Π�D�������.�����������������s��B筼�Z��Lΰ��A��u���-)�����>������v����o��L彼�  �  �N=��M= M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=b�E=E�D=b-D=�jC=��B=b�A=bA=xX@=��?=��>=� >=�6==�k<=�;=g�:=Y:=�19=�_8=s�7=b�6=��5=5=�-4=|Q3=8s2=֒1=M�0=p�/=>�.=��-=2-=5,=[-+=�8*=�@)=�E(=�G'=�E&=�@%=8$=�+#=7"=�!=s�=��=�=y�=�a=3=��=��=��=(I=\=��=�e=�=��=TT=�=��
=0	=��=e'=&�=&=b�= =M�<���<���<i�<s%�<���<��<�,�<��<�b�<=��<j�<��<;��<|��<�s�<��<�O�<���<�<�z�<D״<O0�<f��<�٩<V*�<�x�<�Ğ<U�<�W�<;��<�<*�<�m�<T��<F�<�mz<%�r<�xk<��c<H�\<$U<ϙM<�&F<}�><�H7<6�/<y(<6!<�<�a<V<��<+��;gz�;�
�;��;VZ�;B�;(�;�ؔ;�Ԇ;F�q; V;;�:;�S;�9;���:�R�:��P:�9C 5�͹��L�׵����ʺO���lM��`.�Y(F��]�~�t��օ�T��+<��2����������7!ǻ[uѻ�ۻ������5���a���	�
��E�i��8-������ �#%��0)��I-��S1�[O5��<9�=��@���D��pH��L�\�O�z\S�F�V�6pZ���]��^a���d�g*h�p�k���n�U"r�gu�-�x�X�{�}�6������SC��d҅�4_��ꈼ�r�������~���������3��s���X��A������~u��<h�����fW��Π�/D��Ĺ���.�����������������s��=筼�Z��Eΰ��A��j���,)�����?������w����o��8彼�  �  
�N=��M=�M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=Z�E=:�D=i-D=�jC=��B=`�A=\A=sX@=��?=��>=� >=�6==�k<=�;=b�:=V:=�19=�_8=~�7=i�6=��5= 5=�-4=�Q3=;s2=ܒ1=O�0=y�/==�.=��-=6-=+,=]-+=�8*=�@)=�E(=�G'=�E&=�@%=8$=�+#=9"=�!=o�=��=Ѱ=z�=�a=3=��=��=��=0I=e=��=�e=�=��=TT=�=��
=4	=Ơ=j'=1�=)&=h�=
 =[�<���<���<i�<r%�<���<��<�,�<"��<�b�<?��<i�<��<4��<w��<�s�<���<�O�<t��<�<�z�<1״<K0�<\��<�٩<Z*�<�x�<�Ğ<U�<�W�<+��<"�<�)�<n�<g��<M�<�mz<1�r<�xk<�c<^�\<7U<�M<�&F<h�><I7<�/<
y(<:!<
�<b<`<��<��;Mz�;:
�;��;Z�;��;V�;&ؔ;�Ԇ;�q;�V;�:;�S;�9;ϫ�:�S�:�P:��9"�4�͹ݟL�����]�ʺ����CM��`.�(F���]�_�t�uօ�K���;��02������ڤ���!ǻSuѻ�ۻ��廷�ﻰ5���a����
��E�c��z-����� �l%��0)��I-��S1�nO5��<9��=���@�h�D��pH��L���O�r\S�I�V�GpZ���]�z^a���d�W*h�H�k���n�D"r��fu��x�,�{���/������bC��]҅�:_���鈼�r�������~���������9��x���z��6�������u��9h��!���oW��Π�*D�������.�����������������s��3筼�Z��>ΰ��A��e���)�����4������g����o��C彼�  �  �N=��M=M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=X�E=1�D=d-D=�jC=��B=Y�A=YA=qX@=��?=��>=� >=�6==�k<=#�;=h�:=\:=�19=�_8=��7=i�6=��5=(5=�-4=�Q3=?s2=�1=P�0=�/=A�.=��-==-=/,=c-+=�8*=�@)=�E(=�G'=�E&=�@%=8$=�+#=4"=�!=i�=��=Ͱ=v�=�a=3=��=��=��=)I=c=��=�e=�=��=YT=
�=��
=6	=Ҡ=q'=6�=,&=p�= =^�<���<���<i�<%�<���<���<{,�<��<�b�<9��<W�<��<4��<h��<�s�<���<�O�<d��<��<�z�<$״<L0�<G��<�٩<I*�<�x�<�Ğ<Z�<X�<3��<1�<�)�<n�<l��<T�<nz<C�r<�xk<�c<��\<KU<��M<'F<k�><7I7<3�/<+y(<J!<��<�a<@<��<���;Rz�;

�;ͩ�;�Y�;��;(�;�ה;�Ԇ;��q;oV;��:;S;�9;���:�R�:��P:��9��4�͹v�L�϶���ʺ�����L�`.��'F�W�]�"�t�,օ�J���;��2����������p!ǻ%uѻ)�ۻΤ�����5���a���
��E�y���-�+���� ��%��0)�J-��S1��O5�=9�=��@�v�D��pH��L�u�O�X\S�=�V�7pZ���]�x^a�^�d�C*h�;�k���n�)"r��fu��x��{���$��򱂼WC��S҅�C_���鈼�r������
���������I��}������=�������u��F*h������W��Π�:D�������.�����������������s��(筼�Z��8ΰ��A��\���)�����#������d����o��C彼�  �  �N=��M=�M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=N�E=/�D=V-D=�jC=t�B=O�A=TA=lX@=��?=��>=� >=�6==�k<=�;=d�:=]:=�19=`8=��7=q�6=��5=-5=�-4=�Q3=Js2=�1=^�0=|�/=H�.=��-=;-=5,=Z-+=�8*=�@)=�E(=�G'=�E&=�@%=8$=�+#=%"=�!=^�=��=ΰ=i�=�a=
3=��=��=��=*I=`=��=�e=�=��=_T=�=��
=F	=ؠ={'=B�=:&=y�= =w�<���<���<#i�<�%�<���<��<�,�<��<�b�<:��<W�<��<'��<[��<�s�<���<�O�<Z��<��<�z�<"״<60�<H��<�٩<O*�<�x�<�Ğ<V�<�W�<>��</�<*�<n�<n��<n�<-nz<t�r<yk<H�c<��\<{U<	�M<'F<��><7I7<E�/<y(<<!<�<�a<L<��<���;	z�;�	�;W��;�Y�;|�;��;�ה;=Ԇ;��q;�V;<�:;�R;_9;۪�:4R�:�P:��9��4�͹��L�ⴘ�+�ʺ����ZL��_.�H'F��]���t�օ�����;���1����������C!ǻquѻ�ۻ�����5���a��7�
��E�����-�X��2� �%�1)�J-�T1��O5�=9�=��@���D��pH��L�a�O�a\S�(�V�pZ���]�B^a�O�d� *h��k���n�"r��fu��x��{�M�$��󱂼YC��e҅�1_��ꈼ�r���������������W���������\������u��c,h��5����W�� Π�3D�������.������������������s��$筼�Z��ΰ��A��E���)��휶�������^����o��$彼�  �  �N=��M=M= aL=��K=��J=�*J=�lI=��H=��G=�0G=�pF=A�E=)�D=N-D=�jC=h�B=S�A=MA=bX@=��?=��>=� >=�6==�k<=�;=k�:=c:=�19=`8=��7=��6=��5=25=�-4=�Q3=Ts2=�1=m�0=��/=L�.=��-=:-=<,=Z-+=�8*=�@)=�E(=�G'=�E&=�@%=�7$=�+#="=�!=Z�=��=ð=^�=�a=�2=��=��=�=-I=]=��=�e=�=��=eT=�=��
=Y	=۠=�'=I�=D&=��=" =��<���<Ť�<+i�<�%�<��<��<�,�<��<�b�<'��<M�<��<��<d��<ms�<���<�O�<P��<��<�z�<#״<0�<F��<}٩<M*�<�x�<�Ğ<b�<X�<N��<*�<*�<n�<���<��<4nz<��r<yk<z�c<��\<�U<L�M<'F<��><0I7<b�/< y(<O!<�<�a<N<u�<���;�y�;�	�;P��;5Y�;F�;d�;�ה;�ӆ;�q;pV;��:;�R;�8;ڪ�:pQ�:��P:C�9S��4�͹/�L������ʺ����9L��_.��&F���]���t�օ�p���;���1������ʤ��!ǻvuѻ͠ۻ
��	��6��/b��m�
��E�����-�j��E� ��%�@1)��I-�8T1��O5�3=9�,=�
�@���D��pH��L�C�O�]\S��V�pZ���]��]a�J�d��)h���k�x�n��!r��fu���x��{�D���豂�JC��a҅�'_��ꈼ�r�����������Ƅ��O���������l������u��k*h��L����W��;Π�6D��ȹ���.��������������s��筼�Z��ΰ��A��-����(��֜����s���=����o��彼�  �  �N=��M=M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=?�E=�D=I-D=�jC=g�B=G�A=?A=_X@=��?=��>=� >=�6==�k<= �;=n�:=e:=�19=`8=��7=��6=��5=?5=�-4=�Q3=^s2=��1=i�0=��/=R�.=��-=E-=<,=_-+=�8*=�@)=�E(=�G'=�E&=�@%=�7$={+#="=�!=S�=��=��=]�=}a=�2=��=��=��=&I=^=��=�e=�=��=pT= �=Ą
=W	=�=�'=P�=K&=��=, =��<��<ͤ�<Ii�<�%�<��<���<�,�<��<�b�<-��<J�<{�<���<I��<ls�<���<�O�<:��<��<�z�<�ִ<0�<=��<}٩<@*�<�x�<�Ğ<\�<
X�<J��<A�<%*�<4n�<���<~�<gnz<��r<?yk<��c<ۆ\<�U<Y�M<D'F<ȶ><cI7<`�/</y(<M!<��<�a<2<{�<���;�y�;U	�;��;Y�;��;5�;(ה;�ӆ;2�q;zV;3�:;DR;�8;���:�P�:t�P:��96�4�͹;�L�������ʺ*����K��^.�{&F�S�]�h�t��Յ����1;���1��V���|���!ǻPuѻ�ۻ��K��.6��<b�#���
�3F�����-����^� ��%�G1)�<J-�VT1��O5�A=9�5=�)�@���D��pH��L�F�O�8\S���V��oZ�q�]�^a��d��)h��k�g�n��!r��fu���x���{�=���᱂�HC��Z҅�7_��ꈼ�r�����������݄��k���������u��!����u��tNh��Q����W��;Π�BD��չ���.���������񋩼����{s��筼�Z��ΰ��A������(��ʜ�����u���8���jo��彼�  �  �N=��M=
M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=9�E=�D=D-D=�jC=a�B=:�A=?A=[X@=z�?=��>=� >=�6==�k<=�;=o�:=b:=�19=`8=��7=��6=��5=D5=�-4=�Q3=\s2=�1=n�0=��/=U�.=��-=E-=:,=d-+=�8*=�@)=�E(=�G'=�E&=�@%=�7$=q+#="=�!=H�=��=��=Z�=qa=�2=��=��=�=#I=h=��=�e=�=��=sT=$�=̈́
=Z	=��=�'=a�=V&=��== =��<��<Ӥ�<Ni�<�%�<��<���<�,�<#��<�b�<2��<7�<p�<��<.��<cs�<���<�O�<!��<��<�z�<�ִ<0�<��<~٩<<*�<�x�<�Ğ<N�<X�<E��<G�<&*�<An�<���<��<�nz<��r<uyk<��c<�\<�U<h�M<f'F<˶><sI7<X�/<>y(<9!<�<�a<%<}�<��;�y�;,	�;���;�X�;x�;�;�֔;�ӆ;?�q;hV;�:;[Q;�8;���:�Q�:*�P:J�9X��48�͹Y�L�㴘�z�ʺB���K��^.� &F�g�]���t�OՅ�u�� ;���1��S�������*!ǻ-uѻO�ۻѤ�O��(6��Bb�_�|�
�aF����.������ ��%�W1)�oJ-�LT1��O5�Q=9�-=�9�@�u�D��pH��L�K�O�<\S���V��oZ�R�]�^a���d��)h���k�A�n��!r�Kfu���x���{�7���求�FC��W҅�<_���鈼�r������2�����ڄ���������������:����u���\h��P����W��9Π�ED��ʹ���.�����������������zs���歼Z���Ͱ�tA�� ����(��ǜ�����[���1���[o��彼�  �  "�N=��M=M=�`L=��K=��J=z*J=�lI=��H=��G=�0G=�pF=0�E=�D==-D=�jC=Y�B=7�A=<A=VX@=y�?=��>=� >=�6==�k<="�;=v�:=j:=�19=`8=��7=��6=��5=H5=�-4=�Q3=bs2=	�1=v�0=��/=[�.=��-=I-=A,=h-+=�8*=�@)=�E(=�G'=�E&=�@%=�7$=q+#="=�!=G�=��=��=P�=qa=�2=��=��=�= I=d=��=�e=�=��={T=-�=΄
=e	=��=�'=h�=_&=��=D =��<��<��<[i�<�%�<+��<��<�,�<��<�b�<$��<5�<i�<���<,��<Qs�<���<�O�<��<��<�z�<�ִ<0�<��<n٩<0*�<�x�<�Ğ<W�<X�<T��<L�<9*�<Dn�<���<��<�nz<��r<�yk<��c<�\<�U<~�M<g'F<�><~I7<w�/<Uy(<K!<�<�a<<X�<��;Vy�;	�;���;�X�;X�;��;�֔;5ӆ;�q;&V;��:;0Q;8;!��:�P�:h�P:N�9>�5��͹H�L�������ʺ�����J�o^.��%F�7�]�=�t�;Յ�8��;��`1�����f���� ǻuѻ4�ۻ���}��[6��Vb�i���
�cF�$��.������ �
	%��1)�rJ-�eT1��O5�`=9�G=�J�@���D��pH��L�-�O�*\S���V��oZ�U�]��]a���d��)h���k�%�n��!r�5fu���x���{�����ױ��6C��S҅�<_��ꈼ�r������5�����䄐����΄��������=����u���\h��Z����W��HΠ�QD��׹���.���������狩�����hs���歼xZ���Ͱ�sA������(���������M���'���[o��彼�  �   �N=��M=M=�`L=��K=��J=�*J=�lI=��H=��G=�0G=�pF=,�E=�D=4-D=�jC=S�B=4�A=2A=SX@=|�?=��>=� >=�6==�k<= �;=l�:=g:=�19=`8=��7=��6=��5=T5=�-4=�Q3=ts2=�1=z�0=��/=`�.=��-=I-==,=_-+=�8*=�@)=�E(=�G'=�E&=�@%=�7$=l+#="=�!=>�=��=��=J�=oa=�2=��=��=�=+I=a=��=�e=�=��={T=2�=҄
=k	=��=�'=h�=f&=��=D =��<!��<���<Zi�<�%�<��<���<�,�<��<�b�<��<;�<i�<��<)��<Ds�<���<yO�<��<��<�z�<�ִ<�/�<&��<e٩<7*�<�x�<�Ğ<[�<X�<O��<K�<>*�<Ln�<���<��<�nz<%�r<ryk<��c<2�\<�U<��M<t'F<��><zI7<o�/<(y(<Q!<��<�a<&<C�<1��;y�;��;`��;oX�;:�;w�;{֔;ӆ;��q;wV;<�:;`Q;�7;	��:�P�:#�P:!�9,��4��͹�L�9�����ʺ|����J��].�F%F���]�*�t�2Յ����:��>1�����h���!ǻbuѻ�ۻ��;��R6��bb�T���
�xF�:��-.����� �	%��1)�J-��T1��O5�`=9�J=�#�@���D��pH��L�F�O�/\S���V��oZ�I�]��]a���d�v)h���k��n�k!r�;fu�m�x���{������ޱ��IC��[҅�:_��ꈼ�r������0������������܄��������H����u���jh��p����W��RΠ�ID��ι���.���������싩�����cs���歼kZ���Ͱ�hA��𴳼�(���������M������Uo���佼�  �  '�N=��M=M= aL=��K=��J=w*J=�lI=��H=��G=�0G=�pF=,�E=�D=3-D=�jC=T�B=0�A=3A=OX@=s�?=��>=� >=�6==�k<=$�;=u�:=o:=�19=`8=��7=��6=��5=S5=�-4=�Q3=rs2=�1=��0=��/=c�.=��-=P-=D,=g-+=�8*=�@)=�E(=�G'=�E&=�@%=�7$=h+#=	"=�!=;�=��=��=L�=ja=�2=��=��=�=#I=_=��=�e=�=��=T=6�=ׄ
=p	=�=�'=m�=g&=��=H =��<*��<���<di�<�%�</��<��<�,�<��<�b�<��<(�<]�<��<��<Fs�<���<vO�<��<��<�z�<�ִ<�/�<��<_٩<%*�<�x�<�Ğ<Z�<X�<\��<Z�<=*�<Rn�<���<��<�nz<�r<�yk<��c<<�\<U<��M<�'F<��><�I7<��/<My(<T!<��<�a<<9�<���;y�;��;H��;lX�;�;k�;P֔;ӆ;y�q;�V;��:;�P;Z7;ȧ�:�P�:��P:��9��5��͹
�L�Y���>�ʺ�����J��].�E%F��]�Q�t�&Յ�����:��%1�����1���� ǻ uѻ/�ۻ+��x�ﻥ6��xb�|���
��F�3��1.����� � 	%��1)��J-��T1��O5�~=9�p=�E�@���D��pH��L�&�O�\S���V��oZ�7�]��]a���d�)h���k�	�n�u!r�-fu�n�x���{������˱��5C��L҅�>_��ꈼ�r������D������������ۄ��������S����u���lh��n����W��XΠ�\D��Թ���.���������ߋ������cs���歼hZ���Ͱ�bA�������(���������C������No���佼�  �  ��N=��M=�"M=�gL=��K=��J=k3J=�vI=!�H=6�G=�<G=�}F=6�E=��D==D=�{C=3�B=�A='2A=Wm@=��?=��>=+>=gP==t�<=M�;=��:=2!:= R9=��8=��7=��6=�6=�/5=�V4=;|3=��2=��1=��0=��/=*/=/.=�D-=2W,=g+=
t*=�})=��(='�'=;�&=��%=�}$=�r#=�c"=Q!=: =�=-�=�=X�=�=�R=�={�=K�=X=�=�=f=�
=s�=�D=��
=�i	=��=`z=�=�v=��=` =I��<lm�<�6�<���<��<�`�<�	�<��<5E�<���<se�<��<�l�<���<7]�<���<|9�<���<��<�b�<齸<��<Oj�<໭<�
�<�V�<���<��<�.�<=s�<��<���<O8�<x�<0��<���<�hz<%�r<Sbk<��c<�^\<�T<aM<l�E<Bl><8�6<{�/<�(<� <D<�<i�
<2<���;�4�;Ʋ�;@�;�޽;���;qQ�;�'�;�;�'n;oWR;ȶ6;�H;� ;��:J~�:�>:�Ϫ9�d��,|��	�`��٢���Ժ].�C����3���K�9)c��cz�⥈���������ܴ�|���c�ɻ�OԻ�x޻�x�7P�S���M���s�������-x�C��$"�;A&�Ec*��u.��x2�(m6�US:�3,>���A��E�jI�xM�ԭP��?T��W��D[�p�^�%b��e�S�h��6l���o���r�v�Q>y��p|���+b��E�����h������!������,������0��s����.��%���(��𢖼���^���=��:���h����o���䠼5Y��
ͣ�m@������O&��ߘ��*��]}��aﭼpa��qӰ��E��÷���)������B��A�������ki���ݽ��  �  ��N=��M=�"M=�gL=��K=��J=q3J=vI=�H=;�G=�<G=�}F=4�E=��D==D=�{C=2�B=�A=/2A=[m@=��?=��>=3>=bP==r�<=O�;=��:=9!:="R9=��8=��7=��6=�6=�/5=�V4=4|3=��2=��1=��0=��/='/=/.=�D-=7W,=g+=t*=�})=��(=$�'=,�&=��%=�}$=�r#=�c"=Q!=: =�=/�=�=`�=�=�R=�=u�=P�=X=�=�=f=�
=u�=�D=��
=�i	=��=_z=�=�v=��=` =?��<hm�<�6�<���<&��<�`�<�	�<��<&E�<���<ae�<���<�l�<���<F]�<���<�9�<���<��<�b�<�<��<Uj�<໭<�
�<W�<���<��<�.�<Bs�<%��<���<W8�<x�<)��<���<ihz<0�r<7bk<��c<�^\<��T<aM<_�E<Kl><:�6<��/<�(<� <�C<��<��
<�1<n��;�4�;��;�@�;�޽;���;�Q�;�'�;�;0(n;�WR;�6;hH;  ;��:�}�:��>:�Ъ9�`���x��k�`�0٢���Ժ�.�2���3���K��)c�xcz�N������������۴�\���>�ɻ�OԻ�x޻�x� P�d�������s��������)x����"�2A&�9c*�iu.��x2�$m6��S:�H,>���A��E��iI�qM�ĭP�z?T��W��D[�n�^�%b�R�e�R�h��6l���o���r�Pv�b>y��p|���%b��8�����d������!��|���0,��)����0��i����.��&���(��⢖����c���3��%���b����o���䠼.Y��	ͣ�z@������J&��Ϙ��%��V}��hﭼwa���Ӱ��E������*������L��U�������pi���ݽ��  �  ��N=��M=�"M=�gL=��K=��J=|3J=�vI=)�H=7�G=�<G=�}F=4�E=�D==D=�{C=4�B=�A=&2A=]m@=��?=��>=;>=`P==t�<=M�;=��:=6!:=R9=��8=��7=��6=�6=�/5=�V4=-|3=��2=��1=��0=��/=!/=/.=�D-=4W,=g+=t*=�})=��(=.�'=4�&=��%=�}$=�r#=�c"=Q!=: =�=0�=�=^�=�=�R=�=~�=T�=X=�=�=f=�
=q�=�D=��
=�i	=��=cz=�=�v=��=` =B��<^m�<�6�<���<��<�`�<}	�<��<E�<���<qe�<��<�l�<���<H]�<���<�9�<���<��<�b�<���<��<Ij�<���<�
�<W�< ��<��<�.�<7s�<"��<���<R8�<x�<'��<���<ehz<7�r<bk<��c<�^\<��T<�`M<K�E<@l><�6<��/<�(<� <�C<��<��
<�1<���;�4�;��;�@�;�޽;��;�Q�;(�;�;F(n;nWR;J�6;"I;� ;�:�}�:U�>:�Ъ9jg���y���`��٢�%�Ժ�.�����3�ٟK�*c�cz�O�����������ܴ�����S�ɻ�OԻ�x޻�x�P����h��s���Ț�w�"x����"�.A&�,c*�qu.��x2��l6�uS:�#,>���A��E��iI��M�ѭP��?T�$�W��D[�u�^�%b�T�e�?�h��6l�˂o���r�Nv�X>y��p|�-��1b��>�����h������!��m���,�����0��y����.��"���(��碖����b���.��0���n����o���䠼Y��ͣ�{@������U&��Ҙ��3��Z}��tﭼza���Ӱ��E������*������M��T�������yi���ݽ��  �  ��N=��M=�"M=�gL=��K=��J=s3J=�vI=%�H=@�G=�<G=�}F=B�E=�D=$=D=�{C=A�B=&�A=12A=`m@=��?=��>=0>=gP==s�<=K�;=��:=3!:=R9=��8=��7=��6=�6=�/5=�V4=-|3=z�2=��1=��0=��/= /=/.=D-=5W,=g+=t*=�})=��(=*�'=7�&=��%=�}$=�r#=�c"=Q!=: =�=;�=�=d�=��=�R=�=|�=I�=X=�=�=f=�
=o�=�D=��
=�i	=��=Mz=
�=�v=��=�_ ="��<Rm�<�6�<���<��<�`�<z	�<��</E�<���<te�<��<�l�<���<W]�<���<�9�<ʠ�<��<�b�<��<��<_j�<�<�
�<W�<���<��<�.�<As�<��<���<N8�<	x�<��<���<<hz<��r<bk<��c<q^\<��T<�`M<B�E<5l><&�6<��/<�(<�� <	D<�<��
<2<���;5�;3��;A�;b߽;P��;�Q�;j(�;��;�(n;7XR;��6;I;� ;��:�~�:^�>:\Ъ9M[��z���`��٢�v�Ժ=/�H����3�@�K��)c�Edz�r����*�����ܴ�����B�ɻ�OԻ�x޻�x�;P�4���X���s������M��w����"��@&��b*�Uu.�x2�m6�gS:�(,>���A��E�jI�qM�ɭP��?T�#�W��D[���^�G%b�`�e���h��6l��o��r�]v��>y��p|�1��/b��D��i������!������,�����~0��`����.������'��Ԣ�����H����� ���Y����o���䠼'Y��
ͣ�m@������L&��ט��/��_}��wﭼ�a���Ӱ��E��ط��*������g��e�������}i���ݽ��  �  ��N=��M=�"M=�gL=��K=��J=w3J=�vI=(�H=N�G=�<G=�}F=E�E=�D=0=D=�{C=D�B=%�A=<2A=mm@=��?=��>=6>=nP==o�<=L�;=��:=(!:=R9=��8=��7=��6=�6=�/5=�V4=$|3=r�2=��1=��0=��/=/=/.=zD-=*W,=g+=t*=�})=��(=1�'==�&=��%=�}$=�r#=�c"=Q!=: =�=?�= �=f�=�=�R=�=��=N�=X=�=�=�e=�
=e�=�D=��
=�i	=��=Ez=�=�v=��=�_ =��<Fm�<�6�<w��<���<�`�<y	�<٪�<:E�<���<�e�<��<�l�<���<T]�<���<�9�<��<��<�b�<��<��<}j�<���<�
�<W�<
��<��<�.�<?s�<��<���<68�<�w�<
��<���<Dhz<��r<�ak<��c<s^\<��T<�`M<$�E<�k><�6<O�/<�(<� <D<�<��
<)2<���;�5�;u��;A�;�߽;���;OR�;�(�;��;	)n; YR;v�6;fI; ;��:��: �>:�Ѫ9�a���~����`��ڢ���Ժ�/�_����3���K�p*c��dz�_���2�T��3��Kܴ�������ɻ�OԻ�x޻dx�P�����=��|s�Q����F��w�����"��@&��b*�Ku.�Kx2��l6�RS:�,>���A�ͶE�jI�oM��P��?T�D�W�'E[���^�e%b�a�e���h��6l��o��r�dv��>y��p|�]��<b��X�����f������� ��x���
,�����g0��G����.������'������}��?��������<����o���䠼Y���̣�n@������O&��𘩼7��v}���ﭼ�a���Ӱ��E��鷳�-*������e��l��������i���ݽ��  �  ~�N=��M=�"M=�gL=��K=��J=|3J=�vI=8�H=L�G=�<G=�}F=Q�E=�D=2=D=�{C=Q�B=8�A=<2A=rm@=��?=��>==>=gP==r�<=K�;=��:=,!:=R9=��8=~�7=��6=�6=�/5=�V4=|3=q�2=��1=��0=��/=/=/.=yD-=*W,=g+=
t*=�})=��(=3�'=B�&=Є%=�}$=�r#=�c"=!Q!=%: =�=I�=/�=u�=��=�R=�=��=U�=X=�=�=�e=�
=`�=�D=��
=�i	=��=Az=��=�v=��=�_ =���<+m�<�6�<h��< ��<�`�<o	�<ݪ�<&E�<���<|e�<!��<�l�<���<x]�<��<�9�<��<��<�b�<4��<��<sj�<��<�
�<W�<��<��<�.�<2s�<��<���<28�<�w�<���<���<�gz<��r<�ak<t�c<8^\<t�T<�`M<��E<�k><�6<]�/<�(<�� <D<�<��
<%2<J��;�5�;���;�A�;�߽;���;oR�;)�;'�;S*n;!YR;�6;=J;} ;��:%�:/�>:YҪ94g���{����`�3ۢ���Ժ�/�b��D�3�J�K�]+c��dz����~򓻬��Q��^ܴ�������ɻ�OԻ�x޻�x��O�����(��9s�l�a����w�����"��@&��b*�u.�ex2��l6�6S:�,>���A���E�jI��M���P��?T�R�W�9E[�Ϲ^��%b���e���h�.7l�2�o�)�r��v��>y��p|�o��Fb��Q����l������!��i���,������T0��M����.��㫓��'������e��%���������F����o���䠼Y���̣�r@������\&��阩�=��{}���ﭼ�a���Ӱ��E��񷳼Q*��Ü��������������i���ݽ��  �  o�N=��M=�"M=�gL=��K=��J=�3J=�vI=>�H=T�G=�<G=�}F=U�E=*�D=@=D=�{C=Q�B=A�A=H2A=zm@=��?=��>=G>=gP==w�<=H�;=��:=)!:=R9=��8=n�7=��6=�6=�/5=�V4=
|3=e�2=��1=��0=��/=/=/.=mD-=-W,=
g+=t*=�})=��(=7�'=C�&=ل%=�}$=�r#=�c"=+Q!=2: =�=U�=-�=��=�=�R=�=��=[�=X=�=ڻ=�e=�
=R�=�D=��
=�i	=p�=1z=��=�v=��=�_ =��<m�<�6�<J��<��<�`�<c	�<��<!E�<���<~e�<'��<�l�<���<�]�<���<�9�<��<
�<�b�<:��<�<�j�<)��<�
�<.W�<��<��<�.�<)s�<��<���<(8�<�w�<䶄<���<�gz<��r<zak<U�c<�]\<\�T<v`M<��E<�k><��6<[�/<}(<�� <D<"�<ч
<,2<���;�5�; ��;�A�;�;���;�R�;�)�;6�;+n;�YR;��6;�J;� ;b�:x�:�>:�Ѫ9�c���|��چ`��ڢ���Ժ0����:�3���K��+c�Rez�z���|���_���ܴ����m�ɻ�OԻ�x޻�x軔O����!��s�@�*����w����d"��@&��b*��t.�?x2��l6�.S:��+>���A���E��iI��M��P��?T�~�W�;E[�
�^��%b���e���h�W7l�S�o�g�r��v��>y�%q|�i��`b��]����u������!��V���,������E0��7����.��竓��'������I��������ボ�4����o���䠼Y���̣�q@������f&��嘩�[���}���ﭼ�a���Ӱ��E�����e*��ќ��������������i���ݽ��  �  m�N=��M=�"M=�gL=��K=��J=�3J=�vI=?�H=a�G=�<G=�}F=g�E=1�D=J=D=�{C=b�B=C�A=Q2A=�m@=��?=
�>=D>=mP==t�<=H�;=��:=!!:=R9=�8=d�7=��6=�6=�/5=�V4=�{3=W�2=��1=��0=��/=/=/.=kD-=$W,=g+=t*=�})=��(==�'=O�&=ք%=�}$=�r#=d"=9Q!=9: =�=b�=:�=��=�=�R=�=��=V�=X=�=ٻ=�e=�
=M�=�D=��
=�i	=o�=!z=��=�v=��=�_ =Қ�<�l�<q6�<C��<��<`�<a	�<ڪ�<)E�<���<�e�<7��<�l�<���<�]�<��<�9�<��<�<c�<N��<�<�j�<)��<�
�<3W�<��<��<�.�<'s�<���<���<8�<�w�<ʶ�<~��<�gz<`�r<@ak<�c<�]\<<�T<8`M<��E<�k><��6<2�/<s(<� <D<-�<ԇ
<j2<���;66�;Z��;)B�;��;�;FS�;�)�;��;D+n;�ZR;�6;BK;� ;R�:]��:߻>:Ӫ9�f��S����`��ۢ���Ժ�0������3�`�K��,c�fz�^�����L������ܴ������ɻ�OԻ�x޻px軞O�~������s� �$����Dw�]��<"�S@&�}b*��t.�x2��l6�S:��+>���A�߶E�jI��M��P��?T���W�ZE[�/�^��%b��e��h��7l���o���r��v�
?y�Nq|����bb��g�
���s������� ��]����+��⮍�=0�� ����.��ǫ���'������=���������ك������o���䠼 Y���̣�l@������h&������_���}���ﭼ�a���Ӱ��E������*��������������i���ݽ��  �  n�N=��M=�"M=�gL=��K=��J=�3J=�vI=B�H=k�G=�<G=~F=s�E=8�D=\=D=�{C=v�B=Q�A=\2A=�m@=ç?=�>=A>=tP==o�<=L�;=��:=!:=R9=o�8=j�7=��6=w6=v/5=�V4=�{3=L�2=��1=��0=��/=�/=�..=kD-=W,=g+=t*=�})=��(=:�'=T�&=ۄ%=�}$=�r#=d"=<Q!=E: =	=c�=P�=��=�=�R=�=��=W�=X=�=�=�e=�
=D�=�D=��
=�i	=]�=z=��=�v=��=�_ =���<�l�<L6�<8��<ٯ�<o`�<h	�<ʪ�<5E�<���<�e�<;��<�l�<���<�]�<F��<�9�<7��<*�<)c�<p��<"�<�j�<1��<�<,W�<'��<��<�.�<3s�<�<���<8�<�w�<Ƕ�<X��<xgz<-�r<3ak<��c<�]\<��T<'`M<��E<�k><��6<�/<|(<� <D<F�<ć
<|2<���;�6�;���;�B�;�;��;�S�;*�;w�;;,n;�[R;��6;�K; ;A�:���:�>:�ժ9Vj�����h�`�]ݢ���Ժc1���J�3�
�K��,c��fz�ԧ��T�)������ܴ������ɻ�OԻ�x޻Lx軇O�������s�����w�7w�*��"�J@&�#b*��t.��w2��l6��R:��+>���A�ȶE�jI�tM�'�P��?T���W��E[��^��%b�-�e�E�h��7l���o���r�*v�>?y�3q|�͝�hb��k����g����� ��_����+��ܮ��30��
����.�������'��e���)��甙����σ������o���䠼Y���̣�l@������\&�����Z���}���ﭼ�a���Ӱ�F��7����*��������Ƃ������i��޽��  �  g�N=��M=�"M=�gL=��K=��J=�3J=�vI=O�H=q�G==G=~F=r�E=A�D=e=D=�{C=s�B=U�A=b2A=�m@=ͧ?=�>=N>=uP==r�<=K�;=��:=!:=�Q9=l�8=\�7=��6=u6=r/5=�V4=�{3=F�2=��1=��0=x�/=�/=�..=cD-=W,=g+=t*=�})=Ȅ(=C�'=Z�&=�%=�}$=�r#=d"=?Q!=M: ==h�=O�=��= �=�R=�=��=_�=	X=�=ڻ=�e=�
=>�=�D=��
=�i	=Y�=z=��=�v=��=�_ =���<�l�<C6�<%��<Ư�<^`�<a	�<Ϊ�<2E�<���<�e�<L��<m�<	��<�]�<A��< :�<I��<;�<)c�<w��<4�<�j�<I��<�<DW�<.��<��<�.�<$s�<浓<���<�7�<�w�<���<W��<kgz<�r<ak<��c<�]\<��T<`M<k�E<zk><��6<�/<](<� <D<N�<�
<�2<��;�6�;ٴ�;�B�;�;Y��;0T�;[*�;n�;�,n;�[R;A�6;VL;w ; �:Ӂ�:-�>:>֪9	t��_���
�`��ݢ�4�Ժ�1����~�3�}�K��-c�	gz�ᧈ�D󓻉��3��ݴ�C����ɻ�OԻ�x޻Sx�BO�G�������r�����q�(w�	���"�5@&�!b*��t.��w2�Ql6��R:��+>��A�̶E�jI��M�?�P� @T���W��E[�K�^��%b�7�e�X�h��7l�փo���r�0v�R?y�dq|�֝�wb��z�$���k������� ��H����+��ɮ��0������{.�������'��T�����攙�������������o���䠼�X���̣�n@������k&�����j���}���ﭼ�a���Ӱ�F��C����*��������ǂ��%����i��޽��  �  b�N=��M=�"M=�gL= �K=��J=�3J=�vI=R�H=s�G==G=~F=��E=L�D=c=D=�{C=|�B=`�A=j2A=�m@=ϧ?=�>=O>=pP==w�<=C�;=��:=!:=�Q9=q�8=P�7=��6=k6=e/5=�V4=�{3=;�2=}�1=��0=k�/=�/=�..=bD-="W,=g+=t*=�})=ń(=F�'=Y�&=�%=�}$=�r#=d"=RQ!=Q: ==|�=Q�=��=$�=�R=�=��=\�=X=�=λ=�e=�
=9�=�D=��
=�i	=K�= z=��=�v=r�=�_ =���<�l�<H6�<��<ί�<h`�<K	�<ت�<&E�<���<�e�<L��<m�<��<�]�<N��<':�<G��<L�<Lc�<���<L�<�j�<M��<�<JW�<&��<��<�.�<s�<���<x��<8�<�w�<���<B��<4gz<��r<�`k<��c<d]\<��T<�_M<N�E<�k><��6<-�/<Q(<� <D<>�<�
<�2<+��;�6�;-��;C�;��;���;*T�;�*�;��;\-n;�\R;m�6;�L;s ;\�:b��:ܽ>:�Ҫ9�k��A~��߈`��ܢ���Ժ%2����A�3�ȣK�.c��gz�E���~����+��ݴ�H�����ɻPԻzx޻Vx�ZO�*�������r������e��v�����"��?&�b*�`t.��w2�Nl6��R:��+>���A�׶E��iI��M��P��?T���W��E[���^�&b�h�e���h��7l��o��r�Vv�n?y��q|�ǝ�b��o����������� ��I����+��Ǯ��0��﯐�c.������m'��U�����Ô��������������o���䠼�X���̣�h@������v&������r���}���ﭼ b��	԰�,F��U����*��#������݂��8����i�� ޽��  �  Z�N=��M=�"M=�gL=�K= �J=�3J=�vI=U�H=w�G==G=~F=��E=M�D=l=D=�{C=}�B=`�A=j2A=�m@=ѧ?=�>=Q>=uP==x�<=C�;=��:=!:=�Q9=c�8=W�7=��6=h6=d/5=�V4=�{3=:�2=z�1=��0=s�/=�/=�..=YD-=W,=g+=
t*=�})=Ǆ(=I�'=^�&=�%=�}$=�r#=d"=NQ!=U: ==w�=Q�=��='�=�R=�=��=^�=X=�=л=�e=�
=0�=�D=��
=�i	=G�=�y=��=v=p�=�_ =���<�l�<-6�<	��<���<b`�<K	�<ת�<1E�<���<�e�<Q��<m�<��<�]�<O��<:�<V��<Q�<Ic�<��<J�<�j�<W��<�<NW�</��<��<�.�<s�<鵓<f��<�7�<�w�<���<@��<.gz<��r<�`k<��c<b]\<��T<�_M<T�E<Zk><e�6<�/<T(<� <D<T�<�
<�2<F��;�6�;3��;C�;��;đ�;xT�;�*�;��;Z-n;�\R;ۻ6;�L;� ;��:-��:
�>:#Ӫ92n��<�����`��ޢ���Ժ�1����F�3�ۣK��-c��gz�V����󓻫��S��]ݴ�������ɻ�OԻ�x޻@x�CO��������r������c��v�����"��?&�b*�gt.��w2�9l6��R:��+>�{�A�ʶE��iI��M�(�P�#@T���W��E[�e�^�&b�s�e���h��7l��o�	�r�gv�]?y�q|�����b�������~������� ��D����+��®��0��﯐�c.������y'��E�����ǔ��������������o��{䠼�X���̣�e@������s&���������}���ﭼ�a��
԰�.F��\����*��*������߂��*����i��޽��  �  g�N=��M=�"M=�gL=��K=��J=�3J=�vI=S�H=z�G==G=~F=��E=M�D=s=D=�{C=��B=g�A=m2A=�m@=Χ?=�>=J>=tP==u�<=K�;=��:=!:=�Q9=c�8=U�7=��6=b6=f/5=�V4=�{3=7�2={�1=��0=o�/=�/=�..=`D-=W,=g+=	t*=�})=Ą(=C�'=[�&=�%=�}$=�r#=-d"=PQ!=[: ==x�=a�=��=&�=�R=�=��=Z�=X=�=ֻ=�e=�
=@�=�D=��
=�i	=E�=�y=��=uv=p�=�_ =���<�l�<*6�<'��<���<]`�<Z	�<Ъ�<.E�<���<�e�<J��<m�<��<�]�<g��<:�<f��<U�<Pc�<���<U�<�j�<S��<�<AW�<-��<��<�.�<&s�<۵�<~��<�7�<�w�<���<2��<3gz<��r<�`k<y�c<h]\<��T<�_M<?�E<kk><��6<�/<^(<�� <D<G�<�
<�2<7��;7�;^��;_C�;��;���;�T�;�*�;�;�-n;�\R;!�6;�L;� ;��:��:a�>:2ת9n��-�����`�}ޢ���Ժw2�
��!�3�]�K�U.c��gz�S��������g���ܴ�T���#�ɻ�OԻ�x޻Rx�^O�B�������r������ ��v�����"��?&��a*�Tt.��w2�6l6��R:��+>���A�ҶE� jI��M�B�P�@T���W��E[�l�^�7&b�z�e���h�8l��o��r��v��?y��q|����pb���� ���n������� ��O����+��Ȯ��	0����W.��y���'��6����������������������o��~䠼�X���̣�i@������i&�����l���}���ﭼ�a��԰�,F��f����*��9������ꂹ�=����i��޽��  �  Z�N=��M=�"M=�gL=�K= �J=�3J=�vI=U�H=w�G==G=~F=��E=M�D=l=D=�{C=}�B=`�A=j2A=�m@=ѧ?=�>=Q>=uP==x�<=C�;=��:=!:=�Q9=c�8=W�7=��6=h6=d/5=�V4=�{3=:�2=z�1=��0=s�/=�/=�..=YD-=W,=g+=
t*=�})=Ǆ(=I�'=^�&=�%=�}$=�r#=d"=NQ!=U: ==w�=Q�=��='�=�R=�=��=^�=X=�=л=�e=�
=0�=�D=��
=�i	=G�=�y=��=v=p�=�_ =���<�l�<-6�<
��<���<b`�<L	�<ت�<1E�<���<�e�<Q��<m�<��<�]�<O��<:�<V��<Q�<Hc�<��<I�<�j�<V��<�<NW�</��<��<�.�<s�<鵓<f��<�7�<�w�<���<@��<.gz<��r<�`k<��c<b]\<��T<�_M<U�E<Zk><e�6<�/<U(<� <D<U�<�
<�2<G��;�6�;4��;C�;��;đ�;xT�;�*�;��;W-n;�\R;ػ6;�L;� ;��:$��:��>:�Ҫ9�n��f�����`��ޢ���Ժ�1����K�3��K��-c��gz�X����󓻬��U��_ݴ�������ɻ�OԻ�x޻Ax�DO��������r������c��v�����"��?&�b*�gt.��w2�9l6��R:��+>�{�A�ʶE��iI��M�(�P�#@T���W��E[�e�^�&b�s�e���h��7l��o�	�r�gv�]?y�q|�����b�������~������� ��D����+��®��0��﯐�c.������y'��E�����ǔ��������������o��{䠼�X���̣�e@������s&���������}���ﭼ�a��
԰�.F��\����*��*������߂��*����i��޽��  �  b�N=��M=�"M=�gL= �K=��J=�3J=�vI=R�H=s�G==G=~F=��E=L�D=c=D=�{C=|�B=`�A=j2A=�m@=ϧ?=�>=O>=pP==w�<=C�;=��:=!:=�Q9=q�8=P�7=��6=k6=e/5=�V4=�{3=;�2=}�1=��0=k�/=�/=�..=bD-="W,=g+=t*=�})=ń(=F�'=Y�&=�%=�}$=�r#=d"=RQ!=R: ==|�=Q�=��=$�=�R=�=��=\�=X=�=λ=�e=�
=:�=�D=��
=�i	=K�= z=��=�v=r�=�_ =���<�l�<I6�<��<ϯ�<i`�<L	�<٪�<'E�<���<�e�<M��<m�<��<�]�<N��<':�<G��<L�<Lc�<���<K�<�j�<L��<�<IW�<%��<��<�.�<s�<���<w��<8�<�w�<���<B��<3gz<��r<�`k<��c<e]\<��T<�_M<O�E<�k><��6</�/<R(<� <D<@�<�
<�2<.��;�6�;.��;C�;��;���;)T�;�*�;��;X-n;�\R;g�6;zL;k ;K�:P��:��>:JҪ9�l���~��	�`��ܢ���Ժ/2����K�3�ѣK�
.c��gz�I��������.��ݴ�J�����ɻPԻ{x޻Wx�[O�+�������r������f��v�����"��?&�b*�`t.��w2�Nl6��R:��+>���A�׶E��iI��M��P��?T���W��E[���^�&b�h�e���h��7l��o��r�Vv�n?y��q|�ǝ�b��o����������� ��I����+��Ǯ��0��﯐�c.������m'��U�����Ô��������������o���䠼�X���̣�h@������v&������r���}���ﭼ b��	԰�,F��U����*��#������݂��8����i�� ޽��  �  g�N=��M=�"M=�gL=��K=��J=�3J=�vI=O�H=q�G==G=~F=r�E=A�D=e=D=�{C=s�B=U�A=b2A=�m@=ͧ?=�>=N>=uP==r�<=K�;=��:=!:=�Q9=l�8=\�7=��6=u6=r/5=�V4=�{3=F�2=��1=��0=x�/=�/=�..=cD-=W,=g+=t*=�})=Ȅ(=C�'=Z�&=�%=�}$=�r#=d"=?Q!=M: ==h�=O�=��= �=�R=�=��=_�=	X=�=ڻ=�e=�
=>�=�D=��
=�i	=Y�=z=��=�v=��=�_ =���<�l�<E6�<'��<ȯ�<``�<c	�<Ъ�<3E�<���<�e�<M��<m�<
��<�]�<B��< :�<I��<;�<)c�<v��<4�<�j�<I��<�<CW�<-��<��<�.�<#s�<嵓<��<�7�<�w�<���<V��<jgz<�r<ak<��c<�]\<��T<`M<l�E<|k><��6<�/<_(<� <D<P�<��
<�2<��;�6�;ܴ�;�B�;�;Y��;/T�;Y*�;l�;�,n;�[R;9�6;LL;l ;��:���:��>:�ժ9�u��Ԃ��E�`��ݢ�Q�Ժ�1�����3���K��-c�gz�槈�I󓻍��7��ݴ�F����ɻ�OԻ�x޻Vx�DO�H�������r�����r�(w�	���"�6@&�!b*��t.��w2�Ql6��R:��+>��A�̶E�jI��M�?�P� @T���W��E[�K�^��%b�7�e�X�h��7l�փo���r�0v�R?y�dq|�֝�wb��z�$���k������� ��H����+��ɮ��0������{.�������'��T�����攙�������������o���䠼�X���̣�n@������k&�����j���}���ﭼ�a���Ӱ�F��C����*��������ǂ��%����i��޽��  �  n�N=��M=�"M=�gL=��K=��J=�3J=�vI=B�H=k�G=�<G=~F=s�E=8�D=\=D=�{C=v�B=Q�A=\2A=�m@=ç?=�>=A>=tP==o�<=L�;=��:=!:=R9=o�8=j�7=��6=w6=v/5=�V4=�{3=L�2=��1=��0=��/=�/=�..=kD-=W,=g+=t*=�})=��(=:�'=T�&=ۄ%=�}$=�r#=d"=<Q!=E: =	=d�=P�=��=�=�R=�=��=W�=X=�=�=�e=�
=D�=�D=��
=�i	=^�=z=��=�v=��=�_ =���<�l�<N6�<:��<ۯ�<q`�<j	�<̪�<7E�<���<�e�<<��<�l�<���<�]�<F��<�9�<7��<*�<(c�<p��<"�<�j�<0��<�<+W�<%��<��<�.�<2s�<ﵓ<���<8�<�w�<ƶ�<W��<wgz<-�r<3ak<��c<�]\<��T<)`M<��E<�k><��6<�/<~(<� <D<H�<Ǉ
<2<���;�6�;���;�B�;�;��;�S�;*�;u�;4,n;w[R;��6;�K; ;#�:e��:��>:'ժ9�l��������`��ݢ���Ժu1���Z�3��K��,c��fz�ۧ��Y�/�����ݴ������ɻ�OԻ�x޻Ox軉O�������s�����x�7w�+��"�J@&�#b*��t.��w2��l6��R:��+>���A�ȶE�jI�tM�'�P��?T���W��E[��^��%b�-�e�E�h��7l���o���r�*v�>?y�3q|�͝�hb��k����g����� ��_����+��ܮ��30��
����.�������'��e���)��甙����σ������o���䠼Y���̣�l@������\&�����Z���}���ﭼ�a���Ӱ�F��7����*��������Ƃ������i��޽��  �  m�N=��M=�"M=�gL=��K=��J=�3J=�vI=?�H=a�G=�<G=�}F=g�E=1�D=J=D=�{C=b�B=C�A=Q2A=�m@=��?=
�>=D>=mP==t�<=H�;=��:=!!:=R9=�8=d�7=��6=�6=�/5=�V4=�{3=W�2=��1=��0=��/=/=/.=kD-=$W,=g+=t*=�})=��(==�'=O�&=ք%=�}$=�r#=d"=9Q!=:: =�=b�=:�=��=�=�R=�=��=W�=X=�=ٻ=�e=�
=N�=�D=��
=�i	=p�="z=��=�v=��=�_ =Ԛ�<�l�<s6�<E��<��<�`�<c	�<ܪ�<+E�<���<�e�<9��<�l�<���<�]�<��<�9�<��<�<c�<M��<�<�j�<(��<�
�<2W�<��<��<�.�<&s�<���<���<8�<�w�<ʶ�<}��<�gz<`�r<@ak<�c<�]\<=�T<:`M<��E<�k><��6<5�/<v(<� <D</�<ׇ
<m2<���;:6�;]��;+B�;��;�;ES�;�)�;��;<+n;�ZR;�6;4K;� ;1�::��:��>:uҪ9i�������`��ۢ���Ժ�0�����3�q�K��,c�*fz�e�����R������ܴ������ɻ�OԻ�x޻sx軡O�������s��$����Ew�]��<"�T@&�~b*��t.�x2��l6�S:��+>���A�߶E�jI��M��P��?T���W�ZE[�/�^��%b��e��h��7l���o���r��v�
?y�Nq|����bb��g�
���s������� ��]����+��⮍�=0�� ����.��ǫ���'������=���������ك������o���䠼 Y���̣�l@������h&������_���}���ﭼ�a���Ӱ��E������*��������������i���ݽ��  �  o�N=��M=�"M=�gL=��K=��J=�3J=�vI=>�H=T�G=�<G=�}F=U�E=*�D=@=D=�{C=Q�B=A�A=H2A=zm@=��?=��>=G>=gP==w�<=H�;=��:=)!:=R9=��8=n�7=��6=�6=�/5=�V4=
|3=e�2=��1=��0=��/=/=/.=mD-=-W,=
g+=t*=�})=��(=7�'=C�&=ل%=�}$=�r#=�c"=+Q!=2: =�=U�=-�=��=�=�R=�=��=[�=X=�=ڻ=�e=�
=S�=�D=��
=�i	=q�=2z=��=�v=��=�_ =���<	m�<�6�<L��<��<�`�<e	�<��<#E�<���<�e�<)��<�l�<���<�]�<���<�9�<��<
�<�b�<9��<�<�j�<'��<�
�<,W�<��<��<�.�<'s�<��<���<'8�<�w�<㶄<���<�gz<��r<zak<U�c<�]\<^�T<x`M<��E<�k><��6<^�/<�(<�� <D<%�<ԇ
</2<���;�5�;#��;�A�;�;���;�R�;�)�;3�;�*n;�YR;�6;�J;� ;@�:S�:��>:KѪ9#f��7}��-�`�ۢ���Ժ!0���L�3���K��+c�bez���������d���ܴ�
���q�ɻ�OԻ�x޻�x軖O����"��s�A�+����w����e"��@&��b*��t.�?x2��l6�.S:��+>���A���E��iI��M��P��?T�~�W�;E[�
�^��%b���e���h�W7l�S�o�g�r��v��>y�%q|�i��`b��]����u������!��V���,������E0��7����.��竓��'������I��������ボ�4����o���䠼Y���̣�q@������f&��嘩�[���}���ﭼ�a���Ӱ��E�����e*��ќ��������������i���ݽ��  �  ~�N=��M=�"M=�gL=��K=��J=|3J=�vI=8�H=L�G=�<G=�}F=Q�E=�D=2=D=�{C=Q�B=8�A=<2A=rm@=��?=��>==>=gP==r�<=K�;=��:=,!:=R9=��8=~�7=��6=�6=�/5=�V4=|3=q�2=��1=��0=��/=/=/.=yD-=*W,=g+=
t*=�})=��(=3�'=B�&=Є%=�}$=�r#=�c"=!Q!=%: =�=I�=/�=u�=��=�R=�=��=U�=X=�=�=�e=�
=`�=�D=��
=�i	=��=Bz=��=�v=��=�_ =���<-m�<�6�<j��<��<�`�<q	�<ߪ�<(E�<���<~e�<"��<�l�<���<y]�<��<�9�<��<��<�b�<3��<��<rj�<��<�
�<W�<��<��<�.�<0s�<��<���<18�<�w�<���<���<�gz<��r<�ak<t�c<9^\<u�T<�`M<��E<�k><�6<`�/<�(<�� <D<�<��
<(2<N��;�5�;���;�A�;�߽;���;oR�;)�;$�;K*n;YR;�6;/J;n ;��:�:�>:�Ѫ9�i���|���`�Zۢ��Ժ�/�u��V�3�[�K�m+c��dz�����򓻲��W��cܴ�������ɻ�OԻ�x޻�x��O�����)��:s�l�a����w�����"��@&��b*�u.�ex2��l6�6S:�,>���A���E�jI��M���P��?T�R�W�9E[�Ϲ^��%b���e���h�.7l�2�o�)�r��v��>y��p|�o��Fb��Q����l������!��i���,������T0��M����.��㫓��'������e��%���������F����o���䠼Y���̣�r@������\&��阩�=��{}���ﭼ�a���Ӱ��E��񷳼Q*��Ü��������������i���ݽ��  �  ��N=��M=�"M=�gL=��K=��J=w3J=�vI=(�H=N�G=�<G=�}F=E�E=�D=0=D=�{C=D�B=%�A=<2A=mm@=��?=��>=6>=nP==o�<=L�;=��:=(!:=R9=��8=��7=��6=�6=�/5=�V4=$|3=r�2=��1=��0=��/=/=/.=zD-=*W,=g+=t*=�})=��(=1�'=>�&=��%=�}$=�r#=�c"=Q!=: =�=?�= �=f�=�=�R=�=��=N�=X=�=�=�e=�
=f�=�D=��
=�i	=��=Fz=�=�v=��=�_ =��<Hm�<�6�<y��<���<�`�<{	�<۪�<<E�<���<�e�<��<�l�<���<U]�<���<�9�<��<��<�b�<��<��<|j�<���<�
�<W�<	��<��<�.�<>s�<��<���<58�<�w�<	��<���<Chz<��r<�ak<��c<t^\<��T<�`M<&�E<�k><�6<R�/<�(<�� <D< �<��
<,2<���;�5�;x��;A�;�߽;���;NR�;�(�;��;)n;�XR;k�6;ZI;q ;��:��:��>:?Ѫ9�c��s��(�`�ۢ���Ժ�/�p��	�3�ŠK�*c��dz�f���8�Y��8��Pܴ�������ɻ�OԻ�x޻fx�P�����=��}s�Q����F��w�����"��@&��b*�Lu.�Lx2��l6�RS:�,>���A�ͶE�jI�oM��P��?T�D�W�'E[���^�e%b�a�e���h��6l��o��r�dv��>y��p|�]��<b��X�����f������� ��x���
,�����g0��G����.������'������}��?��������<����o���䠼Y���̣�n@������O&��𘩼7��v}���ﭼ�a���Ӱ��E��鷳�-*������e��l��������i���ݽ��  �  ��N=��M=�"M=�gL=��K=��J=s3J=�vI=%�H=@�G=�<G=�}F=B�E=�D=$=D=�{C=A�B=&�A=12A=`m@=��?=��>=0>=gP==s�<=K�;=��:=3!:=R9=��8=��7=��6=�6=�/5=�V4=-|3=z�2=��1=��0=��/= /=/.=D-=5W,=g+=t*=�})=��(=*�'=7�&=��%=�}$=�r#=�c"=Q!=: =�=;�=�=d�=��=�R=�=|�=J�=X=�=�=f=�
=p�=�D=��
=�i	=��=Nz=�=�v=��=�_ =$��<Tm�<�6�<���<��<�`�<|	�<��<0E�<���<ue�<��<�l�<���<W]�<���<�9�<ʠ�<��<�b�<��<��<_j�<�<�
�<W�<���<��<�.�<@s�<��<���<M8�<x�<��<���<<hz<��r<bk<��c<r^\<��T<�`M<D�E<7l><(�6<��/<�(<�� <D<�<��
<2<���;5�;5��;A�;c߽;P��;�Q�;i(�;��;�(n;0XR;��6;I;� ;��:~�:'�>:�Ϫ9]��yz��'�`��٢���ԺK/�U���3�L�K�*c�Pdz�w����.�����ܴ�����E�ɻ�OԻ�x޻�x�=P�6���Y���s������N��w����"��@&��b*�Uu.�x2�	m6�gS:�(,>���A��E�jI�rM�ɭP��?T�#�W��D[���^�G%b�`�e���h��6l��o��r�]v��>y��p|�1��/b��D��i������!������,�����~0��`����.������'��Ԣ�����H����� ���Y����o���䠼'Y��
ͣ�n@������L&��ט��/��_}��wﭼ�a���Ӱ��E��ط��*������g��e�������}i���ݽ��  �  ��N=��M=�"M=�gL=��K=��J=|3J=�vI=)�H=7�G=�<G=�}F=4�E=�D==D=�{C=4�B=�A=&2A=]m@=��?=��>=;>=`P==t�<=M�;=��:=6!:=R9=��8=��7=��6=�6=�/5=�V4=-|3=��2=��1=��0=��/=!/=/.=�D-=4W,=g+=t*=�})=��(=.�'=4�&=��%=�}$=�r#=�c"=Q!=: =�=0�=�=^�=�=�R=�=~�=T�=X=�=�=f=�
=q�=�D=��
=�i	=��=cz=�=�v=��=` =C��<_m�<�6�<���<��<�`�<	�<��< E�<���<re�<��<�l�<���<I]�<���<�9�<���<��<�b�<���<��<Ij�<���<�
�<W�<���<��<�.�<6s�<"��<���<R8�<x�<&��<���<ehz<7�r<bk<��c<�^\<��T< aM<L�E<Al><�6<��/<�(<� <�C<��<��
<�1<���;�4�;��;�@�;�޽;��;�Q�;(�;�;B(n;iWR;D�6;I;� ;��:y}�:.�>:RЪ9�h���y��8�`��٢�:�Ժ�.�����3��K�	*c�cz�S����������ܴ�����U�ɻ�OԻ�x޻�x�P����h��s���Ț�w�"x����"�.A&�,c*�qu.��x2� m6�uS:�#,>���A��E��iI��M�ѭP��?T�$�W��D[�u�^�%b�T�e�?�h��6l�˂o���r�Nv�X>y��p|�-��1b��>�����h������!��m���,�����0��y����.��"���(��碖����b���.��0���n����o���䠼Y��ͣ�{@������U&��Ҙ��3��Z}��tﭼza���Ӱ��E������*������M��T�������yi���ݽ��  �  ��N=��M=�"M=�gL=��K=��J=q3J=vI=�H=;�G=�<G=�}F=4�E=��D==D=�{C=2�B=�A=/2A=[m@=��?=��>=3>=bP==r�<=O�;=��:=9!:="R9=��8=��7=��6=�6=�/5=�V4=4|3=��2=��1=��0=��/='/=/.=�D-=7W,=g+=t*=�})=��(=$�'=,�&=��%=�}$=�r#=�c"=Q!=: =�=/�=�=`�=�=�R=�=u�=Q�=X=�=�=f=�
=u�=�D=��
=�i	=��=`z=�=�v=��=` =@��<im�<�6�<���<'��<�`�<�	�<��<&E�<���<be�<���<�l�<���<F]�<���<�9�<���<��<�b�<�<��<Uj�<߻�<�
�<W�<���<��<�.�<Bs�<%��<���<V8�<x�<)��<���<ihz<0�r<7bk<��c<�^\<��T<aM<`�E<Kl><;�6<��/<�(<� <�C<��<��
<�1<o��;�4�;��;�@�;�޽;���;�Q�;�'�;�;.(n;�WR;�6;eH;� ;��:�}�:r�>:�Ъ9-a���x����`�;٢���Ժ�.�7��!�3���K��)c�|cz�P������������۴�]���?�ɻ�OԻ�x޻�x�!P�e�������s��������)x����"�2A&�9c*�iu.��x2�$m6��S:�H,>���A��E��iI�qM�ĭP�z?T��W��D[�n�^�%b�R�e�R�h��6l���o���r�Pv�b>y��p|���%b��8�����d������!��|���0,��)����0��i����.��&���(��⢖����c���3��%���b����o���䠼.Y��	ͣ�z@������J&��Ϙ��%��V}��hﭼwa���Ӱ��E������*������L��U�������pi���ݽ��  �  �N=1�M=)M=|nL=��K=`�J=�<J=��I=�H=H=oIG=\�F=��E=jE=�MD=��C=��B=�	B=�FA=�@=��?=�>=�2>=k==X�<=��;=�;='A:=�s9=f�8=��7=�7=.6=�X5=x�4=n�3=v�2=|�1=>1=�/0=L/=�e.=#}-=��,=e�+=-�*=��)=��(=��'=��&=��%=��$=a�#=M�"=�!=�� =�o=�Q=/=�=B�=�=�s=�8=�=c�=Lg=�=�=�e=2=(�=�3=��	=�L=��=8Q=��=PA=� =�;�<�
�<>��<E��<�A�<4��<���<�/�<g��<T�<K��<(^�<���<P�<���<|,�<J��<���<�S�<뭼<b�<LW�<$��< ��<,>�<���<ˢ<\�<�O�<���<�͓<�
�<�F�<6��<ռ�<���<
bz<��r<�Ik<}�c<�4\<ëT<�$M<T�E<:><Y�6<�#/<ɫ'<�7 <��<�^<��	<4�<X��;��;7M�;^��;T�;+�;J��;�d�;�=�;mXj;�cN;^�2;�;�`�:��:H:�:��+:���9o�����6pu�ȇ����ߺ.��/?!��y9�UeQ���h��#�������f������෻%�»<ͻvQ׻�w�s�VE��;���7�O���{��s����� �m]#���'��+�:�/���3���7��v;��G?��C��F�onJ�N���Q��,U�ެX�0#\�>�_���b�~Pf���i� �l�T6p��ts�t�v�\�y�+
}�Y��騁�7�����L��Tԇ�Z���݊�+`�������_���ݐ��Y���ԓ��N��rǖ�3?��뵙��+������M����������n���ࣼ�R��Ħ�65��0����������0����h��Iٰ��I������q+��t������<���dc��'ֽ��  �  �N=0�M=)M=}nL=��K=_�J=�<J=��I=�H=H=zIG=^�F=��E=rE=�MD=��C=��B=�	B=�FA=#�@=��?=�>=�2>=�j==Y�<=��;=|;=(A:=�s9=o�8=��7=�7=.6=�X5=z�4=t�3=r�2=h�1=?1=�/0=L/=�e.= }-=��,=b�+=2�*=��)=��(=��'=��&=��%=��$=o�#=I�"=�!=�� =�o=�Q=�.=�=K�=�=�s=�8=$�=`�=Pg=�=�=�e=5=(�=�3=��	=�L=��=<Q=��=IA=�� =�;�<�
�<J��<D��<�A�<(��<���<�/�<]��<6T�<P��< ^�<���<!P�<���<{,�<Z��<���<�S�<譼<_�<eW�<0��<��<!>�<ʅ�<ˢ<W�<�O�<���<�͓<�
�<G�<5��<˼�<���<�az<��r<�Ik<�c<T4\<��T<�$M<N�E<[><J�6<�#/<��'<�7 <��<�^<
�	<�<R��; ��;�M�;p��;T�;m�;c��;;e�;�=�;�Xj;]dN;��2;�;�`�:/�:�9�:��+:��9���T���ou�������ߺ2���?!�:z9�'eQ�(�h��#��W����������p෻;�»>ͻ�Q׻aw�%s�E������)7�8���{�� � s���� �W]#�؈'��+��/�ת3��7��v;��G?��C��F�]nJ�N�ĢQ��,U�ϬX�-#\�X�_���b��Pf���i��l�K6p��ts���v�W�y�5
}�K��騁�7�����L��Qԇ�Z���݊�%`�������_��oݐ��Y���ԓ��N��iǖ�?����+��⠜�B����������n���ࣼ�R��Ħ�?5��1����������1����h��Rٰ��I������b+��s������J��$�gc��ֽ��  �  �N=4�M=�(M=�nL=��K=[�J=�<J=��I=�H=H=}IG=b�F=��E=yE=�MD=�C=��B=�	B=�FA=(�@=��?=�>=�2>=�j==`�<=��;=|;=)A:=xs9=i�8=��7=�7=.6=�X5=t�4=h�3=p�2=f�1=H1=�/0=L/=�e.=}-=��,=a�+=8�*=�)=��(=��'=��&=�%=��$=s�#=K�"=�!=�� =�o=�Q=/=�=H�=$�=�s=�8= �=Z�=Vg=�=�=�e=/= �=�3=��	=�L=��=/Q=��=IA=�� =�;�<�
�<=��</��<�A�<(��<���<�/�<P��<0T�<M��<,^�<��<P�<���<z,�<i��<���<�S�<�<e�<nW�<1��<��<!>�<Ʌ�<ˢ<]�<�O�<|��<�͓<�
�<�F�<%��<Ǽ�<��<�az<��r<�Ik<l�c<L4\<ëT<�$M<(�E<B><'�6<�#/<��'<8 <��<�^<�	< �<���;0��;�M�;���;%T�;��;p��;�e�;�=�;1Yj;udN;�2;-;�`�:�:�9�:�+:�9������"ru�6�����ߺ	���?!�+z9��eQ���h��#��g���f���&���෻i�»!ͻ�Q׻,w�9s�/E������"7����{�� �s����� �I]#���'��+���/��3���7��v;��G?��C�,�F�BnJ�N���Q��,U��X�F#\�w�_���b��Pf���i�;�l�q6p��ts���v�I�y�Y
}�W������7�����L��@ԇ�Z���݊�(`�������_��qݐ��Y���ԓ��N��hǖ�?��浙��+��ؠ��A��戟�����n���ࣼ�R��	Ħ�E5��,���������@����h��@ٰ��I������{+��|������;��%�xc��!ֽ��  �  �N=+�M=�(M={nL=��K=e�J=�<J=��I=�H=H=�IG=o�F=��E=~E=�MD=�C=��B=�	B=�FA=-�@=��?=�>=�2>=k==[�<=��;=u;="A:=ws9=a�8=��7=�7= .6=�X5=m�4=b�3=f�2=^�1=21=�/0=L/=�e.=}-=��,=]�+=/�*=��)=��(=��'=��&=�%=��$=y�#=Z�"=$�!=�� =�o=�Q=/=�=Q�=$�=�s=�8=#�=d�=Kg=�=�=�e=&=�=�3=��	=�L=��=&Q=��=:A=� =�;�<v
�<,��<'��<�A�<��<���<�/�<f��<.T�<U��<2^�<��<.P�<���<�,�<s��<���<�S�<��<��<zW�<A��<��<2>�<̅�<#ˢ<f�<�O�<x��<�͓<�
�<�F�<!��<���<���<�az<b�r<zIk<K�c<#4\<y�T<�$M<�E<><*�6<|#/<��'<�7 <��<�^<�	<A�<���;k��;�M�;��;�T�;��;ʡ�;�e�;T>�;Zj;	eN;}�2;q;�a�:E�:K;�:�+:��98��,���qu�ᇭ��ߺѷ�Y@!��z9��eQ�/ i�#$���������0���෻c�»eͻ�Q׻mw��r��D������7����{�� ��r����� �+]#���'���+�Ԯ/���3���7��v;��G?��C���F�gnJ�-N��Q��,U���X�V#\���_���b��Pf��i�U�l��6p��ts�Ҭv���y�f
}�c������)7��Ä��L��Oԇ� Z���݊�`�������_��_ݐ��Y���ԓ��N��Tǖ�?��˵���+��͠��2��鈟�����n���ࣼ�R��Ħ�J5��=���������D����h��hٰ�J�������+���������_��;�}c��2ֽ��  �  �N="�M=)M=~nL=��K=e�J=�<J=��I=�H=H=�IG=r�F=��E=�E=�MD=�C=��B=�	B=�FA=7�@=��?="�>=�2>=	k==S�<=��;=y;=A:=vs9=V�8=��7=�7=�-6=�X5=_�4=X�3=U�2=X�1=)1=�/0=L/=�e.=}-=��,=i�+=-�*=��)=��(=��'=��&=�%=��$=~�#=^�"=+�!=ʉ =p=�Q=/=�=_�='�=�s=�8= �=b�=Fg=�= �=�e==�=�3=��	=�L=~�=Q=��=(A=� =�;�<h
�<��<��<�A�<��<���<�/�<f��<+T�<j��<9^�<��<EP�<���<�,�<���<���<�S�<��<��<�W�<a��<��<K>�<ׅ�<$ˢ<Y�<�O�<���<�͓<�
�<�F�<��<���<���<caz<�r<WIk<�c<�3\<T�T<�$M<�E<�><#�6<V#/<��'<�7 <��<�^<�	<t�<���;���;+N�;#��;�T�;N�;l��;f�;�>�;fZj;�eN;9�2;�;�c�:��:�;�:��+:]��9���ۻ��qu����d�ߺA���@!��{9��fQ�� i��$������I��t���෻k�»�ͻFQ׻xw��r�E�������6� ��>{�� ��r����n ��\#�}�'���+�Ʈ/�z�3���7�pv;��G?��C���F�vnJ� N��Q��,U��X��#\���_��b��Pf�.�i���l��6p�(us��v���y�w
}�{�����/7��Ä��L��]ԇ��Y���݊�`�������_��Gݐ��Y���ԓ�|N��-ǖ��>�������+��������㈟������n���ࣼ�R��Ħ�35��O�����Ƈ��T����h��zٰ�J��к���+���������o��L񺼉c��Gֽ��  �  �N=!�M=�(M=}nL=��K=l�J=�<J=��I=&�H=!H=�IG=��F=��E=�E=�MD=!�C=��B=�	B=�FA=@�@=��?=$�>=�2>=k==]�<=��;=o;=A:=ks9=O�8=��7=�7=�-6=�X5=P�4=G�3=L�2=G�1=$1=�/0=�K/=�e.=}-=��,=`�+=0�*=��)=��(=��'=��&=�%=��$=��#=o�"=;�!=҉ =p=�Q=$/=�=c�=0�=�s=�8=$�=c�=Jg=�=��=�e==�=�3=��	=�L=r�=Q=��=A=ұ =�;�<F
�<���<��<�A�<���<���<�/�<i��<1T�<k��<F^�<(��<PP�<��<�,�<���<���<T�<8��<��<�W�<l��<:��<P>�<Ⅶ<3ˢ<j�<�O�<z��<�͓<�
�<�F�<���<���<���<2az<��r<�Hk<ӽc<�3\<,�T<N$M<џE<�><��6<L#/<��'<�7 <��<�^<1�	<z�<#��;��;�N�;���;\U�;��;���;�f�;/?�;�[j;�fN;�2;�;nd�:��:�<�:�+:_��9��ܻ��su�������ߺ��TA!�	|9�ygQ��i��$��:���m������0᷻��»�ͻ�Q׻Uw��r��D������6����0{�= �~r�[��K ��\#�1�'�I�+�}�/�g�3�}�7�^v;�~G?��C���F�]nJ�N��Q�-U�4�X��#\�֐_�3�b�BQf�R�i���l��6p�Ous� �v���y��
}�������77��Ä��L��Kԇ��Y���݊��_�������_��:ݐ�zY���ԓ�YN��"ǖ��>�������+������	��Ɉ�������n���ࣼ�R��Ħ�J5��S�����҇��i����h���ٰ�-J��庳��+��Ĝ��������h񺼞c��Qֽ��  �  ��N=!�M=�(M=znL=��K=i�J=�<J=��I=4�H=.H=�IG=��F=��E=�E=�MD=3�C=��B=�	B=�FA=M�@=��?=(�>=�2>=
k==Z�<=�;=n;=A:=^s9=M�8=��7=�7=�-6=sX5=E�4=9�3=D�2=3�1=1=�/0=�K/=�e.=}-=��,=Y�+=/�*=��)=��(=��'=��&=&�%=��$=��#=w�"=K�!=�� =%p=�Q=*/=�=l�=?�=�s=�8=*�=_�=Fg=�=��=�e==��=�3=��	=�L=g�=�P=y�=A=�� =t;�<%
�<���<��<�A�<���<���<�/�<`��<BT�<r��<V^�<B��<dP�<9��<�,�<ɓ�<��<9T�<U��<��<�W�<���<Y��<Y>�<���<3ˢ<e�<�O�<m��<�͓<�
�<�F�<ꁈ<o��<���<�`z<��r<�Hk<��c<s3\<�T<$M<��E<�><��6<J#/<q�'<�7 <��<�^<U�	<��<���;���;�N�;��;�U�;i�;8��;Pg�;�?�;�\j;jgN;��2;|;^e�:g�:�<�:հ+:���9i��3��`vu�������ߺT��GB!��|9��gQ�hi�%��ʟ���������p᷻�»�ͻ�Q׻Vw��r뻟D��G����6����{�	 �[r��� �}\#��'�,�+�D�/�;�3�<�7�Bv;�eG?�qC���F�`nJ�;N���Q�8-U�c�X��#\��_�`�b��Qf�r�i���l�/7p�us�h�v��y��
}����3���E7��Ä��L��Pԇ��Y���݊��_������|_��$ݐ�[Y��sԓ�3N�� ǖ��>������p+������������������n���ࣼ�R��Ħ�W5��O���/��އ��z���i���ٰ�TJ�������+��Ӝ��$�����}񺼲c��\ֽ��  �  �N=�M=�(M=|nL=��K=m�J=�<J=ÀI=9�H=8H=�IG=��F=��E=�E=�MD=;�C=��B=�	B=GA=U�@=��?=3�>=�2>=k==\�<=��;=n;=A:=Ys9==�8=��7=�7=�-6=dX5=5�4='�3=1�2=,�1=1=�/0=�K/=�e.= }-=��,=[�+=1�*=�)=��(=��'=��&=)�%=��$=��#=��"=U�!=� =2p= R=</=�=x�=C�=	t=�8=&�=d�=Eg=�=��=�e=�=�=s3=��	=�L=R�=�P=f�=�@=�� =U;�<
�<���<Ҍ�<pA�<���<���<�/�<j��<6T�<���<c^�<M��<|P�<R��<�,�<ٓ�<0��<LT�<v��<��<�W�<���<a��<u>�<���<7ˢ<p�<�O�<u��<�͓<�
�<�F�<Ё�<Z��<{��<�`z<��r<}Hk<g�c<A3\<��T<�#M<m�E<�><��6<$#/<z�'<�7 <��<�^<U�	<Û<Ć�;���;SO�;���;hV�;��;���;�g�;C@�;�]j;ZhN;��2;
;g�:|�:�=�:�+:���9l������vu�>����ߺ߹��B!��}9��hQ�ci��%������6�)��N���᷻�»�ͻ�Q׻=wộr뻜D�����|6�|���z����r������G\#�ɇ'�ޢ+��/��3�'�7�v;�DG?�xC���F�\nJ�3N��Q�P-U���X��#\�5�_���b��Qf���i�;�l�m7p��us���v�2�y�}����<���T7��Ä��L��Nԇ��Y���݊��_��p���o_��
ݐ�@Y��Kԓ�"N���Ɩ��>��a���N+��x���������������n���ࣼ�R��Ħ�P5��a���7����������,i���ٰ�iJ������+������;��������c��wֽ��  �  �N=�M=�(M=snL=��K=y�J=�<J=̀I=>�H=CH=�IG=��F=�E=�E=�MD=D�C=��B=�	B=GA=_�@=��?==�>=�2>=k==[�<={�;=f;=	A:=Ws9=0�8=��7=~7=�-6=TX5=*�4="�3=�2=�1=�1=�/0=�K/=�e.=�|-=��,=W�+=(�*=�)=��(=��'=��&=/�%=��$=��#=��"=]�!=�� =Ap=	R=L/=�=��=H�=t=�8=)�=i�=<g=�=��=�e=�=ڞ=l3=��	=�L=<�=�P=Z�=�@=�� =.;�<�	�<���<ǌ�<cA�<���<{��<�/�<x��<8T�<���<q^�<^��<�P�<[��<-�<��<T��<iT�<���<��<�W�<���<n��<�>�< ��<Nˢ<y�<�O�<j��<�͓<�
�<�F�<���<D��<W��<y`z<<�r<aHk<$�c<3\<h�T<�#M<L�E<S><��6<#/<^�'<�7 <��<_<]�	<�<��;9��;�O�;��;�V�;.��;p��;�g�;�@�;A^j;aiN;n�2;�;�h�:�:�?�:y�+:S��9������vu�����B�ߺ����C!��~9�uiQ��i�&��u�����N������᷻�»�ͻ�Q׻|w�fr�eD������R6�_���z�����q������\#���'���+���/�ȩ3��7��u;�(G?�eC���F�wnJ�=N�1�Q�]-U���X�$\�H�_���b��Qf��i�U�l��7p�vs�ԭv�t�y�}����B���[7��*Ä��L��Sԇ��Y���݊��_��`���\_���ܐ�6Y��,ԓ�N���Ɩ��>��N���3+��^��������������|n���ࣼ�R��*Ħ�[5��n���:��
�������Ai���ٰ��J��;���,�����X��������c���ֽ��  �  �N=�M=�(M=|nL=��K=p�J=�<J=΀I=H�H=IH=�IG=��F=�E=�E=�MD=U�C=�B=�	B=GA=h�@=ʾ?=>�>=�2>=k==Z�<=��;=f;=A:=Ks9=-�8=��7=w7=�-6=NX5=�4=�3=�2=�1=�1=�/0=�K/=�e.=�|-=��,=U�+=/�*=��)=��(=��'=��&=;�%=��$=��#=��"=m�!=	� =Lp=R=O/=�=��=R�=t=�8=*�=\�=?g=�=��=�e=�=Ӟ=[3=��	=}L=2�=�P=G�=�@=�� =;�<�	�<���<���<RA�<���<��<�/�<]��<FT�<���<}^�<o��<�P�<k��<$-�<	��<f��<�T�<���<
�< X�<���<���<�>�<��<Dˢ<k�<�O�<h��<�͓<�
�<�F�<���</��<P��<T`z<�r<Hk<�c<�2\<W�T<�#M<�E<E><m�6<�"/<Z�'<�7 <��<�^<~�	<�<I��;k��;P�;O��;-W�;���;���;�h�;A�;�^j;�iN;�2;Z;i�:u�:Y>�:ݲ+:s9�����Fyu�͌��*�ߺ���C!��~9�OjQ��i�B&�������𖻮����� ⷻl�»�ͻ�Q׻CwỶr�ZD������F6�.��|z�����q����_��[#�_�'���+�խ/���3�ߖ7��u;�G?�ZC���F�dnJ�AN�+�Q��-U���X�0$\���_���b�
Rf��i���l��7p�vs�߭v���y�b}����Y���h7��&Ä��L��Qԇ��Y���݊��_��Q���I_���ܐ�$Y��ԓ��M���Ɩ�d>��6���'+��L��������������pn���ࣼ�R��Ħ�]5��r���T���������Vi���ٰ��J��P���/,��.���h��������c���ֽ��  �  ۜN=�M=�(M=|nL=��K=t�J=�<J=̀I=P�H=KH=�IG=ËF=�E=�E=�MD=^�C=�B=
B=$GA=j�@=Ҿ?==�>=�2>=k==c�<=|�;=`;=A:=Ds9=.�8=��7=q7=�-6=AX5=�4=�3=�2=�1=�1=�/0=�K/=�e.=�|-=��,=H�+=7�*= �)=��(=��'=��&=@�%=��$=Ƚ#=��"=y�!=� =Qp=$R=X/=�=��=V�=t=�8=3�=_�=Gg=�=��=�e=�=ў=O3=��	=mL=(�=�P=?�=�@=�� =;�<�	�<���<���<IA�<���<l��<�/�<`��<VT�<���<�^�<q��<�P�<���<2-�<��<t��<�T�<���<(�<X�<ŧ�<���<�>�<��<Pˢ<x�<�O�<Q��<�͓<�
�<�F�<���< ��<6��<`z<��r<�Gk<ڼc<�2\<#�T<y#M<��E<@><H�6<�"/<.�'<�7 <��<�^<��	<�<���;~��;|P�;���;�W�;���; ��;�h�;cA�;Y`j;�jN;R�2;�;i�:��:�>�:��+:���9�������zu�i�����ߺZ���D!��9��jQ�Ri�k&������������$ⷻ��»�ͻR׻�vỎr�D������76���lz�E���q�R��H��[#�0�'�b�+�}�/���3�˖7��u;�G?�3C���F�>nJ�rN�;�Q��-U�ŭX�5$\���_��b�CRf�=�i���l��7p�Nvs��v���y��}����e���m7��2Ä��L��>ԇ��Y���݊��_��B���F_���ܐ��X��ԓ��M���Ɩ�V>�����	+��1������s�������`n���ࣼ�R��Ħ�u5��q���c���������ci��ڰ��J��X���B,��7����������� d���ֽ��  �  ܜN=�M=�(M=vnL=��K=w�J=�<J=րI=V�H=TH=�IG=��F=�E=�E=�MD=a�C=�B=
B='GA=q�@=ؾ?=F�>=�2>=k==^�<={�;=c;=A:=Ds9=$�8=��7=l7=�-6=<X5=�4=�3=�2=�1=�1=�/0=�K/=�e.=�|-=��,=N�+=/�*=��)=��(=��'=��&=E�%=��$=Ľ#=��"=x�!=� =]p=#R=Z/=�=��=[�=t=�8=0�=^�=?g=�=��=�e=�=ƞ=P3=��	=jL=!�=�P=9�=�@=�� =;�<�	�<���<���<HA�<���<m��<�/�<c��<OT�<���<�^�<��<�P�<���<8-�<"��<���<�T�<���<!�<X�<ק�<���<�>�<��<Qˢ<q�<�O�<X��<�͓<�
�<rF�<���<��<-��<`z<��r<�Gk<��c<�2\<�T<m#M<�E<><I�6<�"/<?�'<�7 <��<	_<��	<�<�;���;�P�;���;�W�;$��;h��; i�;zA�;�_j;�jN;ҥ2;g;Uj�:��:W?�:I�+:[��9������zu�������ߺ����D!��9��jQ�Ui��&�����1������Sⷻ��»�ͻ�Q׻>wỗr�D������6� ��Iz�W���q�U����[#�1�'�Y�+���/���3���7��u;�G?�:C���F�[nJ�ZN�-�Q��-U�٭X�Z$\���_�#�b�HRf�X�i���l� 8p�avs�&�v���y�~}����f���m7��+Ä��L��Kԇ��Y���݊��_��6���7_���ܐ�Y��	ԓ��M���Ɩ�K>�����+��4������g�������dn���ࣼ�R�� Ħ�m5��o���b��%�������fi��ڰ��J��i���E,��E�����������d���ֽ��  �  �N=�M=�(M=xnL=��K=|�J=�<J=؀I=M�H=UH=�IG=ËF=(�E=�E=�MD=d�C=%�B=
B=-GA=r�@=о?=I�>=�2>=k==Y�<=}�;=_;=�@:=Is9=!�8=��7=`7=�-6=>X5=�4=��3=�2=�1=�1=}/0=�K/=�e.=�|-=~�,=R�+=,�*=�)=��(= �'=��&=A�%=��$=��#=��"=|�!=� =Xp='R=h/=�=��=Y�=t=�8=3�=b�=;g=�=��=�e=�=��=F3=v�	=jL=�=�P=0�=�@=�� =�:�<�	�<|��<���<5A�<���<q��<~/�<h��<OT�<���<�^�<���<�P�<���<`-�<)��<��<�T�<Ю�<3�<X�<ڧ�<���<�>�<��<Zˢ<t�<�O�<`��<�͓<�
�<yF�<���<��<!��<`z<��r<�Gk<��c<�2\< �T<D#M<�E<><[�6<�"/<D�'<�7 <��<_<��	<�<y��;���;�P�;���;X�;��;/��;i�;B�;`j;8kN;�2;�;�j�:��:�?�:L�+:���9��9��)yu�������ߺg���D!��9��kQ��i��&������2��4��/ⷻ��»=ͻ�Q׻Ow�nr��C��t���6���<z�_��Zq�A��(��[#�"�'��+���/�s�3���7��u;��F?�,C���F�lnJ�MN�\�Q��-U�ȭX�t$\�Ǒ_�T�b�FRf�g�i���l� 8p�Vvs��v���y��}����^���7��8Ä��L��Uԇ��Y���݊��_��F���4_���ܐ�
Y���ӓ��M���Ɩ�P>������*��0������z�������en���ࣼ�R��Ħ�f5������^���������{i��ڰ��J��y���J,��U�����������d���ֽ��  �  ܜN=�M=�(M=vnL=��K=w�J=�<J=րI=V�H=TH=�IG=��F=�E=�E=�MD=a�C=�B=
B='GA=q�@=ؾ?=F�>=�2>=k==^�<={�;=c;=A:=Ds9=$�8=��7=l7=�-6=<X5=�4=�3=�2=�1=�1=�/0=�K/=�e.=�|-=��,=N�+=/�*=��)=��(=��'=��&=E�%=��$=Ľ#=��"=x�!=� =]p=#R=Z/=�=��=[�=t=�8=0�=^�=?g=�=��=�e=�=ƞ=P3=��	=kL=!�=�P=9�=�@=�� =;�<�	�<���<���<IA�<���<m��<�/�<c��<OT�<���<�^�<���<�P�<���<8-�<"��<���<�T�<���<!�<X�<ק�<���<�>�<��<Qˢ<p�<�O�<X��<�͓<�
�<qF�<���<��<-��<`z<��r<�Gk<��c<�2\<�T<n#M<�E<><J�6<�"/<@�'<�7 <��<
_<��	<�<ć�;���;�P�;���;�W�;$��;h��;�h�;yA�;�_j;�jN;ͥ2;b;Kj�:|�:J?�:/�+:%��9}��Ӿ��zu�������ߺ����D!��9��jQ�[i��&�����3����	��Uⷻ��»�ͻ�Q׻?wỘr�D������6� ��Iz�W���q�U����[#�1�'�Y�+���/���3���7��u;�G?�:C���F�[nJ�ZN�-�Q��-U�٭X�Z$\���_�#�b�HRf�X�i���l� 8p�avs�&�v���y�~}����f���m7��+Ä��L��Kԇ��Y���݊��_��6���7_���ܐ�Y��	ԓ��M���Ɩ�K>�����+��4������g�������dn���ࣼ�R�� Ħ�m5��o���b��%�������fi��ڰ��J��i���E,��E�����������d���ֽ��  �  ۜN=�M=�(M=|nL=��K=t�J=�<J=̀I=P�H=KH=�IG=ËF=�E=�E=�MD=^�C=�B=
B=$GA=j�@=Ҿ?==�>=�2>=k==c�<=|�;=`;=A:=Ds9=.�8=��7=q7=�-6=AX5=�4=�3=�2=�1=�1=�/0=�K/=�e.=�|-=��,=H�+=7�*= �)=��(=��'=��&=@�%=��$=Ƚ#=��"=y�!=� =Rp=$R=X/=�=��=V�=t=�8=3�=_�=Gg=�=��=�e=�=ў=O3=��	=mL=)�=�P=@�=�@=�� =;�<�	�<���<���<JA�<���<m��<�/�<a��<WT�<���<�^�<r��<�P�<���<3-�<��<t��<�T�<���<(�<X�<ħ�<���<�>�<��<Oˢ<w�<�O�<P��<�͓<�
�<�F�<���< ��<6��<`z<��r<�Gk<ۼc<�2\<$�T<z#M<��E<B><I�6<�"/<0�'<�7 <��< _<��	<�<���;���;~P�;���;�W�;���;���;�h�;aA�;T`j;�jN;J�2;�;�h�:��:�>�:^�+:\��9���/���zu������ߺg���D!��9��jQ�]i�p&�����"�������(ⷻ��»�ͻR׻ wỐr�D������86���lz�E���q�R��H��[#�0�'�b�+�}�/���3�˖7��u;�G?�3C���F�>nJ�sN�;�Q��-U�ŭX�5$\���_��b�CRf�=�i���l��7p�Nvs��v���y��}����e���m7��2Ä��L��>ԇ��Y���݊��_��B���F_���ܐ��X��ԓ��M���Ɩ�V>�����	+��1������s�������`n���ࣼ�R��Ħ�u5��q���c���������ci��ڰ��J��X���B,��7����������� d���ֽ��  �  �N=�M=�(M=|nL=��K=p�J=�<J=΀I=H�H=IH=�IG=��F=�E=�E=�MD=U�C=�B=�	B=GA=h�@=ʾ?=>�>=�2>=k==Z�<=��;=f;=A:=Ks9=-�8=��7=w7=�-6=NX5=�4=�3=�2=�1=�1=�/0=�K/=�e.=�|-=��,=U�+=/�*=��)=��(=��'=��&=;�%=��$=��#=��"=m�!=	� =Lp=R=O/=�=��=R�=t=�8=*�=]�=@g=�=��=�e=�=Ԟ=[3=��	=~L=3�=�P=H�=�@=�� =;�<�	�<���<���<TA�<���<���<�/�<^��<HT�<���<^�<p��<�P�<l��<%-�<
��<f��<�T�<���<	�<�W�<���<���<�>�<��<Cˢ<j�<�O�<g��<�͓<�
�<�F�<���<.��<O��<S`z<�r<Hk<�c<�2\<Y�T<�#M<�E<H><p�6<�"/<]�'<�7 <��<�^<��	<��<M��;o��;P�;Q��;.W�;���;���;�h�;A�;�^j;�iN;�2;M;�h�:V�:7>�:��+:���9���T���yu�󌭺P�ߺ"���C!��~9�_jQ��i�I&�������𖻴�����ⷻp�»�ͻ�Q׻Fwỹr�\D������G6�/��}z�����q����_��[#�`�'���+�խ/���3�ߖ7��u;�G?�ZC���F�dnJ�AN�+�Q��-U���X�0$\���_���b�
Rf��i���l��7p�vs�߭v���y�b}����Y���h7��&Ä��L��Qԇ��Y���݊��_��Q���I_���ܐ�$Y��ԓ��M���Ɩ�d>��6���'+��L��������������pn���ࣼ�R��Ħ�]5��r���T���������Vi���ٰ��J��P���/,��.���h��������c���ֽ��  �  �N=�M=�(M=snL=��K=y�J=�<J=̀I=>�H=CH=�IG=��F=�E=�E=�MD=D�C=��B=�	B=GA=_�@=��?==�>=�2>=k==[�<={�;=f;=	A:=Ws9=0�8=��7=~7=�-6=TX5=*�4="�3=�2=�1=�1=�/0=�K/=�e.=�|-=��,=W�+=(�*=�)=��(=��'=��&=/�%=��$=��#=��"=]�!=�� =Ap=	R=L/=�=��=H�=t=�8=)�=j�==g=�=��=�e=�=۞=l3=��	=�L==�=�P=[�=�@=�� =0;�<�	�<���<Ɍ�<fA�<���<}��<�/�<{��<:T�<���<r^�<`��<�P�<\��<-�<��<T��<iT�<���<��<�W�<���<l��<�>�<���<Lˢ<w�<�O�<i��<�͓<�
�<�F�<���<C��<V��<x`z<;�r<aHk<$�c<3\<i�T<�#M<O�E<V><��6<#/<a�'<�7 <��<_<`�	<�<���;>��;�O�;��;�V�;.��;o��;�g�;�@�;7^j;ViN;`�2;�;�h�:��:u?�:"�+:���97��i��.wu�����p�ߺѺ��C!��~9��iQ��i�&��}�����T������᷻�»�ͻ�Q׻�w�jr�gD������S6�`���z�����q������\#���'���+���/�ȩ3��7��u;�(G?�eC���F�wnJ�=N�1�Q�]-U���X�$\�H�_���b��Qf��i�U�l��7p�vs�ԭv�t�y�}����B���[7��*Ä��L��Sԇ��Y���݊��_��`���\_���ܐ�6Y��,ԓ�N���Ɩ��>��N���3+��^��������������|n���ࣼ�R��*Ħ�[5��n���:��
�������Ai���ٰ��J��;���,�����X��������c���ֽ��  �  �N=�M=�(M=|nL=��K=m�J=�<J=ÀI=9�H=8H=�IG=��F=��E=�E=�MD=;�C=��B=�	B=GA=U�@=��?=3�>=�2>=k==\�<=��;=n;=A:=Ys9==�8=��7=�7=�-6=dX5=5�4='�3=1�2=,�1=1=�/0=�K/=�e.= }-=��,=[�+=1�*=�)=��(=��'=��&=)�%=��$=��#=��"=U�!=� =2p= R=</=�=x�=C�=	t=�8=&�=e�=Fg=�=��=�e=�=�=t3=��	=�L=S�=�P=g�=�@=�� =X;�<
�<���<Ռ�<sA�<���<���<�/�<m��<9T�<���<e^�<O��<}P�<S��<�,�<ٓ�<1��<LT�<u��<��<�W�<���<_��<s>�<���<5ˢ<n�<�O�<s��<�͓<�
�<�F�<ρ�<Y��<z��<�`z<��r<}Hk<h�c<B3\<��T<�#M<p�E<�><��6<(#/<~�'<�7 <��<�^<X�	<Ǜ<ʆ�;���;WO�;���;jV�;��;���;�g�;?@�;�]j;MhN;��2;�;�f�:Q�:�=�:��+:���9	�����Hwu�r���A�ߺ����B!��}9��hQ�xi��%�����?�0��U���᷻�»�ͻ�Q׻Awờr뻟D�����}6�}���z����r������G\#�ʇ'�ߢ+��/��3�'�7�v;�DG?�xC���F�\nJ�3N��Q�P-U���X��#\�5�_���b��Qf���i�;�l�m7p��us���v�2�y�}����<���T7��Ä��L��Nԇ��Y���݊��_��p���o_��
ݐ�@Y��Kԓ�"N���Ɩ��>��a���N+��x���������������n���ࣼ�R��Ħ�P5��a���7����������,i���ٰ�iJ������+������;��������c��wֽ��  �  ��N=!�M=�(M=znL=��K=i�J=�<J=��I=4�H=.H=�IG=��F=��E=�E=�MD=3�C=��B=�	B=�FA=M�@=��?=(�>=�2>=
k==Z�<=�;=n;=A:=^s9=M�8=��7=�7=�-6=sX5=E�4=9�3=D�2=3�1=1=�/0=�K/=�e.=}-=��,=Y�+=/�*=��)=��(=��'=��&=&�%=��$=��#=w�"=K�!=�� =%p=�Q=*/=�=l�=?�=�s=�8=*�=_�=Gg=�=��=�e==��=�3=��	=�L=h�=�P=z�=A=�� =w;�<(
�<���<��<�A�<���<���<�/�<c��<DT�<t��<X^�<D��<eP�<:��<�,�<ʓ�<��<9T�<T��<��<�W�<���<X��<X>�<�<1ˢ<c�<�O�<k��<�͓<�
�<�F�<遈<n��<���<�`z<��r<�Hk<��c<u3\<�T<"$M<��E<�><��6<N#/<u�'<�7 <��<�^<X�	<��<���;���;�N�;��;�U�;i�;7��;Mg�;�?�;�\j;]gN;�2;i;5e�::�:�<�:q�+:뼃9������vu�Չ���ߺn��`B!��|9�hQ�}i�%��ԟ���������w᷻�»�ͻ�Q׻Zw��r뻢D��J����6����{�
 �\r��� �}\#��'�,�+�D�/�;�3�<�7�Bv;�eG?�qC���F�`nJ�;N���Q�8-U�c�X��#\��_�`�b��Qf�r�i���l�/7p�us�h�v��y��
}����3���E7��Ä��L��Pԇ��Y���݊��_������|_��$ݐ�[Y��sԓ�3N�� ǖ��>������p+������������������n���ࣼ�R��Ħ�W5��O���/��އ��z���i���ٰ�TJ�������+��Ӝ��$�����}񺼲c��\ֽ��  �  �N=!�M=�(M=}nL=��K=l�J=�<J=��I=&�H=!H=�IG=��F=��E=�E=�MD=!�C=��B=�	B=�FA=@�@=��?=$�>=�2>=k==]�<=��;=o;=A:=ks9=O�8=��7=�7=�-6=�X5=P�4=G�3=L�2=G�1=$1=�/0=�K/=�e.=}-=��,=`�+=0�*=��)=��(=��'=��&=�%=��$=��#=o�"=;�!=҉ =p=�Q=$/=�=c�=1�=�s=�8=%�=d�=Jg=�=��=�e==�=�3=��	=�L=s�=Q=��=A=ӱ =�;�<I
�<���<��<�A�<���<���<�/�<l��<4T�<n��<H^�<*��<RP�<��<�,�<���<���<T�<8��<��<�W�<k��<8��<N>�<ᅦ<1ˢ<h�<�O�<x��<�͓<�
�<�F�<���<���<���<1az<��r<�Hk<Խc<�3\<.�T<P$M<ԟE<�><��6<O#/<��'<�7 <��<�^<5�	<}�<)��;��;�N�;���;^U�;��;���;�f�;+?�;�[j;�fN;�2;�;Fd�:��:�<�:��+:���9���D��.tu�щ����ߺ��lA!�!|9��gQ��i��$��C���u������6᷻��»�ͻ�Q׻Yw��r��D�������6����1{�> �r�\��K ��\#�2�'�I�+�~�/�g�3�~�7�^v;�G?��C���F�]nJ�N��Q�-U�4�X��#\�֐_�3�b�BQf�R�i���l��6p�Ous� �v���y��
}�������77��Ä��L��Kԇ��Y���݊��_�������_��:ݐ�zY���ԓ�YN��"ǖ��>�������+������	��Ɉ�������n���ࣼ�R��Ħ�J5��S�����҇��i����h���ٰ�-J��庳��+��Ĝ��������h񺼞c��Qֽ��  �  �N="�M=)M=~nL=��K=e�J=�<J=��I=�H=H=�IG=r�F=��E=�E=�MD=�C=��B=�	B=�FA=7�@=��?="�>=�2>=	k==S�<=��;=y;=A:=vs9=V�8=��7=�7=�-6=�X5=_�4=X�3=U�2=X�1=)1=�/0=L/=�e.=}-=��,=i�+=-�*=��)=��(=��'=��&=�%=��$=~�#=^�"=+�!=ʉ =p=�Q=/=�=`�='�=�s=�8= �=c�=Fg=�=�=�e==�=�3=��	=�L=�=Q=��=)A=� =�;�<k
�<��<!��<�A�<��<���<�/�<h��<-T�<l��<;^�<��<FP�<���<�,�<���<���<�S�<��<��<�W�<`��<��<J>�<օ�<"ˢ<W�<�O�<���<�͓<�
�<�F�<��<���<���<baz<�r<WIk<�c<�3\<V�T<�$M<�E<�><'�6<Y#/<��'<�7 <��<�^<�	<w�<ǅ�;���;/N�;&��;�T�;O�;k��;f�;�>�;]Zj;�eN;+�2;�;�c�:��:�;�:N�+:���9���9���qu�D�����ߺW���@!��{9��fQ�� i��$��ɞ��Q��{���෻p�»�ͻJQ׻|w��r�E�������6���?{�� ��r����n ��\#�}�'���+�Ʈ/�z�3���7�pv;��G?��C���F�vnJ�N��Q��,U��X��#\���_��b��Pf�.�i���l��6p�(us��v���y�w
}�{�����/7��Ä��L��]ԇ��Y���݊�`�������_��Gݐ��Y���ԓ�|N��-ǖ��>�������+��������∟������n���ࣼ�R��Ħ�35��O�����Ƈ��T����h��zٰ�J��к���+���������o��L񺼉c��Gֽ��  �  �N=+�M=�(M={nL=��K=e�J=�<J=��I=�H=H=�IG=o�F=��E=~E=�MD=�C=��B=�	B=�FA=-�@=��?=�>=�2>=k==[�<=��;=u;="A:=ws9=a�8=��7=�7= .6=�X5=m�4=b�3=f�2=^�1=21=�/0=L/=�e.=}-=��,=]�+=/�*=��)=��(=��'=��&=�%=��$=y�#=Z�"=%�!=�� =�o=�Q=/=�=Q�=$�=�s=�8=#�=d�=Lg=�=�=�e='=�=�3=��	=�L=��='Q=��=;A=� =�;�<x
�<.��<)��<�A�<��<���<�/�<h��<0T�<W��<3^�<��</P�<���<�,�<t��<���<�S�<��<��<zW�<@��<��<1>�<˅�<!ˢ<e�<�O�<w��<�͓<�
�<�F�< ��<���<���<�az<b�r<zIk<L�c<#4\<z�T<�$M<�E<><,�6<#/<��'<�7 <��<�^<
�	<D�<���;n��;�M�;��;�T�;��;ɡ�;�e�;Q>�;Zj; eN;r�2;d;�a�:&�:);�:��+:���9f��x��)ru����7�ߺ��j@!��z9��eQ�> i�*$���������5���෻g�»iͻ�Q׻pw��r� E������7����{�� ��r����� �,]#���'���+�Ԯ/���3���7��v;��G?��C���F�gnJ�-N��Q��,U���X�V#\���_���b��Pf��i�U�l��6p��ts�Ҭv���y�f
}�c������)7��Ä��L��Oԇ� Z���݊�`�������_��_ݐ��Y���ԓ��N��Tǖ�?��˵���+��͠��2��鈟�����n���ࣼ�R��Ħ�J5��=���������D����h��hٰ�J�������+���������_��;�}c��2ֽ��  �  �N=4�M=�(M=�nL=��K=[�J=�<J=��I=�H=H=}IG=b�F=��E=yE=�MD=�C=��B=�	B=�FA=(�@=��?=�>=�2>=�j==`�<=��;=|;=)A:=xs9=i�8=��7=�7=.6=�X5=t�4=h�3=p�2=f�1=H1=�/0=L/=�e.=}-=��,=a�+=8�*=�)=��(=��'=��&=�%=��$=s�#=K�"=�!=�� =�o=�Q=/=�=H�=$�=�s=�8= �=Z�=Vg=�=�=�e=/=!�=�3=��	=�L=��=0Q=��=IA=�� =�;�<�
�<>��<1��<�A�<*��<���<�/�<Q��<1T�<N��<-^�<��<P�<���<{,�<j��<���<�S�<�<e�<nW�<0��<��< >�<ȅ�<ˢ<\�<�O�<{��<�͓<�
�<�F�<%��<Ƽ�< ��<�az<��r<�Ik<m�c<M4\<īT<�$M<)�E<D><(�6<�#/<��'<8 <��<�^<�	<"�<���;3��;�M�;���;%T�;��;o��;�e�;�=�;+Yj;odN;	�2;$;�`�:	�:x9�:��+:���9�����Xru�P����ߺ���?!�7z9��eQ���h��#��l���k���*���෻l�»$ͻ�Q׻.w�:s�1E������"7����{�� �s����� �I]#���'��+���/��3���7��v;��G?��C�,�F�BnJ�N���Q��,U��X�F#\�w�_���b��Pf���i�;�l�q6p��ts���v�H�y�Y
}�W������7�����L��@ԇ�Z���݊�(`�������_��qݐ��Y���ԓ��N��hǖ�?��浙��+��ؠ��A��戟�����n���ࣼ�R��	Ħ�E5��,���������@����h��@ٰ��I������{+��|������;��%�xc��!ֽ��  �  �N=0�M=)M=}nL=��K=_�J=�<J=��I=�H=H=zIG=^�F=��E=rE=�MD=��C=��B=�	B=�FA=#�@=��?=�>=�2>=�j==Y�<=��;=|;=(A:=�s9=o�8=��7=�7=.6=�X5=z�4=t�3=r�2=h�1=?1=�/0=L/=�e.= }-=��,=b�+=2�*=��)=��(=��'=��&=��%=��$=o�#=I�"=�!=�� =�o=�Q=�.=�=K�=�=�s=�8=$�=`�=Pg=�=�=�e=5=(�=�3=��	=�L=��=<Q=��=JA=�� =�;�<�
�<K��<E��<�A�<)��<���<�/�<^��<6T�<Q��< ^�<���<"P�<���<|,�<[��<���<�S�<譼<_�<dW�<0��<��<!>�<ʅ�<ˢ<V�<�O�<���<�͓<�
�<G�<5��<ʼ�<���<�az<��r<�Ik<�c<T4\<��T<�$M<N�E<\><K�6<�#/<��'<�7 <��<�^<�	< �<T��;!��;�M�;p��;T�;m�;c��;;e�;�=�;�Xj;ZdN;��2;�;�`�:#�:�9�:��+:ۺ�9Y��p��pu�������ߺ8���?!�@z9�-eQ�.�h��#��Y����������r෻=�»?ͻ�Q׻bw�&s�E������)7�9���{�� � s���� �W]#�؈'��+��/�ת3��7��v;��G?��C��F�]nJ�N�ĢQ��,U�ϬX�-#\�X�_���b��Pf���i��l�K6p��ts���v�W�y�5
}�K��騁�7�����L��Qԇ�Z���݊�%`�������_��oݐ��Y���ԓ��N��iǖ�?����+��⠜�B����������n���ࣼ�R��Ħ�?5��1����������1����h��Rٰ��I������b+��s������J��$�gc��ֽ��  �  ˡN=��M=S/M=�uL=��K=K=7FJ=��I=L�H=-H=|VG=V�F=��E=TE=^D=�C=��B=�B=\A=��@=A�?=�?=�L>=��==6�<=��;=*-;=Db:=�9=w�8=��7=�(7=�V6=,�5=��4=]�3='�2=�!2=�D1=#e0=5�/=�.=$�-=��,=Z�+=�*=� *=O)=�(=Z'=�&=%=�$=g #=��!=9� =!�=o�=1�=a=6==��=n�=�V=�=��=�v=!=��=�d=^�=s�=� 
=��=�-=�=%=2�=I=���<��<�q�<�*�<���<Ƃ�<�"�<��<�K�<���<�X�<���<WL�<T��<�(�<k��<��<]N�<B��<J��<�M�<���<��<h.�<�s�<K��<���<J5�<�q�<���<}�<��<%V�<���<�<��<�Zz<A�r<0k<��c<x\<^vT<b�L<vXE<�=<�D6<��.<�>'<;�<�H<��<Mf	<��<_7�;ـ�;B��;�?�;���;!A�;�ݝ;���;#S�;[\f;�AJ;YW.;y�;>:�:z��:̓�:h�:"}59��o�u;$���������2�:��E('��x?��wW��#o�u=�����j=��<�������Ż�-лQ{ڻ8��L���a��������e
�	��y�R��3?�e� ��$�o�(���,���0�X�4�t�8�(�<�&p@��+D���G��}K�BO���R��#V���Y��
]��o`���c�� g��mj���m���p�
(t��Xw��z�:�}��d��'�N}��3������������P���	������ ����������v��햼�b���י�mK�������0��٢��������S���Ye��զ��D��鳩�#��8���7��%p��E߰�=N�������,��]������|��e캼#]��]ν��  �  ¡N=��M=F/M=�uL=��K=K=FFJ=�I=M�H=%H=~VG=V�F=��E=UE=p^D=�C=��B=�B=\A=��@=C�?=?=�L>=��==8�<=��;= -;=:b:=�9=��8=��7=�(7=�V6=%�5=��4=h�3='�2=�!2=�D1=e0=;�/=��.=�-=��,=I�+=�*=� *=Z)=�(=]'=�&=%=�$=c #=��!=1� =�=u�=-�=a=6=	=��=y�=�V=�=��=�v=!=��=�d=e�=e�=� 
=�=�-=��="%=-�=D=���<��<�q�<�*�<���<���<�"�<��<�K�<���<�X�<���<ML�<S��<�(�<k��<��<?N�<B��<W��<�M�<���<��<g.�<�s�<g��<���<O5�<�q�<ᬗ<p�<��<6V�<���<�<��<�Zz<H�r<E0k<��c<C\<YvT<T�L<nXE<*�=<�D6<��.<[>'<)�<�H<��<�f	<��<l7�;���;Q��;�?�;���;2A�;�ݝ;ύ�;1S�;�\f;�AJ;�V.;��;;�:$��:I��:�:;t59t�o��=$�N���ؾ��3���c('��x?�wW��"o�n=��B�������=���;�������Ż�-л�{ڻB��6��~a�������e
����x�`��?��� ��$�W�(���,�s�0�a�4�z�8��<��o@��+D���G�~K��O��R�$V���Y��
]��o`���c�� g��mj���m���p�(t�Yw��z�f�}��d��1�c}��E��������𔉼6��ᕌ������� ��	��������v��3햼�b���י�oK������1��ۢ����ᄢ�D���Ue��զ��D������ #��&���6��2p��C߰�VN�������,��W�����|��k캼&]��Hν��  �  ��N=��M=I/M=�uL=��K=K=BFJ= �I=X�H=)H=�VG=Z�F=��E=eE=z^D=��C=��B=�B=#\A=��@=K�?=�?=�L>=��==:�<=��;='-;=Ab:=�9=��8=r�7=�(7=�V6=�5=��4=R�3=!�2=�!2=�D1=
e0=:�/=�.=�-=��,=I�+=�*=� *=R)=�(=^'=�&=%=�$=a #=��!=@� =!�=��=*�=a=6==��=q�=�V=�=��=�v=!=��=�d=d�=U�=� 
=�=�-=�=%=#�=8=���<ʯ�<�q�<{*�<���<Â�<�"�<��<�K�<���<�X�<���<WL�<Z��<�(�<h��<2��<RN�<_��<i��<�M�<ț�<��<}.�<�s�<_��<���<I5�<�q�<欗<��<��<-V�<���<�<��<�Zz<*�r<�/k<��c<$\<MvT<0�L<CXE<�=<�D6<ʿ.<h>'<9�<�H<��<yf	<��<�7�;���;���;�?�;귺;�A�;�ݝ;c��;BS�;5]f;BJ;jW.;;�;�:�:ޥ�:b��:*�:rx59��o��;$��������5�E���('�[y?�RxW�)$o��=���������/>���;������Żv-л�{ڻ��o�a�������e
����x�f���>�D� �߻$��(���,�L�0�\�4�_�8��<�p@��+D���G��}K��O��R�!$V��Y��
]�p`���c�!g��mj��m���p�8(t�6Yw��z���}��d��A�W}��2�������� ���?��알�������������������lv�� 햼�b��vי�jK��}����0��Ƣ����ꄢ�W���\e��զ��D��ݳ��,#��0���D��Hp��D߰�fN�������,��i���'�� |��|캼:]��Nν��  �  ��N=��M=A/M=�uL=��K=K=LFJ=	�I=\�H=7H=�VG=h�F=��E=jE=�^D=��C=��B=�B=+\A=��@=P�?=?=�L>=��==9�<=��;=-;=9b:=�9=u�8=r�7=�(7=�V6=�5=��4=G�3=�2=�!2=�D1=e0=1�/=�.=�-=��,=E�+=�*=� *=c)=�(=f'=�&=%=�$=r #=��!=G� =,�=��=;�=&a=6==��=z�=�V=�=��=�v=� =��=�d=W�=Q�=� 
=ө=�-=٫=%=�='=���<Ư�<�q�<i*�<���<���<�"�<��<�K�<���<�X�<���<lL�<i��<)�<���<8��<pN�<i��<w��<�M�<؛�<��<�.�<�s�<v��<���<S5�<�q�<ڬ�<n�<��<V�<���<}<���<�Zz<�r<�/k<f�c<\<vT<�L<5XE<��=<�D6<��.<C>'<&�<�H<��<�f	<�<�7�;.��;���;U@�;?��;�A�;jޝ;���;�S�;^f;�BJ;dX.;��;a<�:���:n��:��:�y59�o� =$�G��������4����)'�yy?��xW��$o��=��þ��_��@>��+<��L���Ż�-л�{ڻ��/��-a����ǽ�be
�����x����>�$� ���$��(���,� �0�4�4�9�8��<��o@��+D���G��}K��O�#�R�$$V�D�Y��
]�p`���c�L!g��mj��m��p�G(t�mYw�R�z���}��d��M�d}��O��������蔉�#��ؕ��������������������ev��햼�b��gי�KK��o����0��������Ԅ��7���Re��զ��D������,#��I���M��Xp��i߰�qN������-��w���/��D|���캼?]��gν��  �  ��N=��M=G/M=�uL=��K=K=IFJ=�I=c�H=EH=�VG=x�F=��E=yE=�^D=�C=��B=�B=7\A=��@=W�?=?=�L>=��==2�<=��;=-;=4b:=��9=d�8=f�7=�(7=�V6=�5=��4=?�3=�2=�!2=~D1=�d0=#�/=ڞ.=�-=��,=N�+=�*=� *=[)=�(=p'=�&=-%=�$=� #=�!=X� ==�=��=Q�=,a=-6= =��=}�=�V=�=��=�v=� =��=�d=E�=C�=� 
=ĩ=j-=˫=�$=�==���<���<iq�<W*�<���<���<�"�<Һ�<�K�<���<�X�<���<�L�<���<)�<���<S��<�N�<���<���<N�<曵<��<�.�<�s�<u��<���<P5�<�q�<鬗<[�<��<�U�<���<f<���<>Zz<��r<�/k<�c<�\<�uT<��L<XE<��=<�D6<r�.<V>'<(�<yH<��<�f	<I�<$8�;���;4��;�@�;︺;mB�;ߝ;��;�T�;_f;�CJ;QY.;S�;?>�:8��:���:��:U�59 �o��=$����������5뺘��
*'��z?��yW�$%o�^>��(������>���<����� �Ż.л�{ڻ:��3��_a�������?e
����~x�����>�څ �f�$���(�I�,��0���4��8�Ʀ<��o@��+D���G�~K�jO�3�R�+$V�a�Y��
]�@p`��c�z!g�nj�3�m�F�p��(t��Yw���z�̩}��d��X�m}��Q��������ꔉ�2��Õ�����������΅������Jv���얼�b��@י�'K��a����0���������ք��>���We��զ��D�����0#��a���c��op��߰��N��ͽ��-������Y��X|���캼U]���ν��  �  ��N=��M=</M=�uL=��K=!K=PFJ= �I=o�H=NH=�VG=��F=��E=�E=�^D=#�C=��B=�B=K\A=Ù@=c�?=?=�L>=��==;�<=��;=-;=,b:=�9=\�8=V�7=�(7=�V6=�5=w�4=,�3=��2=�!2=rD1=�d0=�/=О.=�-=��,=A�+=�*=� *=`)=�(=z'=�&=;%=�$=� #=�!=h� =K�=��=Y�==a=<6='=��=��=�V=�=��=�v=� =��=�d=8�=*�=� 
=��=S-=��=�$=�==}��<|��<Rq�<5*�<���<~��<�"�<ۺ�<�K�<���<�X�<���<�L�<���<?)�<Ə�<}��<�N�<���<���<!N�<��<��<�.�<�s�<���<���<f5�<�q�<Ӭ�<U�<��<�U�<n��<=<���<�Yz<i�r<J/k<Śc<j\<�uT<|�L<�WE<~�=<>D6<Z�.<(>'<�<�H<��<�f	<r�<�8�;��;���;nA�;m��;C�;�ߝ;Ώ�;�T�;W`f;EJ;Z.;C�;�?�:P��:+��:��:q}59��o��>$�ḅ�¸��7뺆���*'��{?��zW�/&o��>��������?���<�����t�Ż5.л�{ڻ.��Ĕ�3a��n�p��e
�h��+x����@>��� �+�$��(�!�,���0���4���8���<��o@��+D���G��}K��O�P�R�e$V���Y�
]��p`�>�c��!g�jnj�z�m���p��(t��Yw�΄z��}��d��r򁼀}��d��"������֔��)���������k����������s���v���얼fb��"י�	K��6����0���������Ǆ��7���Be��!զ��D�����O#��u���|���p���߰��N���:-����|��q|���캼r]���ν��  �  ��N=��M=7/M=�uL=��K=#K=_FJ=%�I=~�H=]H=�VG=��F=��E=�E=�^D=9�C=��B=B=W\A=ԙ@=p�?=%?=�L>=��==:�<=��;=-;=(b:=�9=Q�8=F�7=�(7=�V6=��5=e�4=�3=��2=�!2=`D1=�d0=
�/=Ȟ.=��-=��,==�+=�*=� *=g)=�(=�'=�&=F%=�$=� #=2�!=|� =_�=��=f�=Pa=F6=6= �=��=�V=�=��=�v=� =��=�d=%�=�=� 
=��=@-=��=�$=ט=�=X��<W��</q�<*�<z��<s��<~"�<Ӻ�<�K�<���<	Y�<���<�L�<���<c)�<��<���<�N�<ܧ�<���<AN�<6��<��<�.�<�s�<���<��<b5�<�q�<ˬ�<P�<��<�U�<L��< <���<�Yz<%�r<�.k<�c<\<>uT<<�L<}WE<O�=<D6<I�.<>'<�<�H<�<�f	<��<9�;v��;m��;�A�;��;�C�;+��;���;�U�;�af;FJ;`[.;S�;>A�:���:l��:B�:��59��o��>$�t���ø�39�7��,'��|?��{W��'o�J?��E������w?��;=��	����ŻK.л
|ڻ��ߔ��`��7�M���d
�6���w�Z���=�?� �պ$�&�(���,�c�0���4���8�x�<�yo@�s+D���G��}K��O�Y�R�w$V���Y�E]��p`���c�"g��nj�ֳm���p�.)t�+Zw��z�N�}�e���򁼇}��h��!������ޔ�����������I����������V����u���얼8b���֙��J������0��t����������-���He�� զ��D�����^#����������p���߰��N�����p-��✶�����|���캼�]���ν��  �  ��N=��M=6/M=�uL=��K=)K=cFJ=.�I=��H=mH=�VG=��F=��E=�E=�^D=I�C=�B="B=d\A=�@=y�?=,?=�L>=��==9�<=��;=	-;=b:=�9=?�8=9�7=�(7=�V6=̂5=N�4= �3=��2=�!2=LD1=�d0=��/=��.=��-=u�,=A�+=�*=� *=i)=�(=�'=�&=S%=$=� #=A�!=�� =t�=ɨ=}�=^a=P6=C=�=��=�V=�=��=�v=� =��=�d=�=�={ 
=��=%-=��=�$=��=�=)��<6��<q�<*�<V��<^��<"�<ʺ�<�K�<���<Y�<���<�L�<н�<�)�<��<���<O�< ��<��<nN�<T��<�<�.�<t�<���<��<c5�<�q�<Ϭ�<1�<��<�U�<*��<<u��<YYz<��r<�.k<�c<�\<�tT<��L<:WE<�=<�C6<�.<>'<�<�H<�<�f	<��<[9�;���;���;�B�;���;�D�;�;,��;QV�;cf;GJ;�\.;�;�B�:���:j��:�:}�59��o��A$�㹅� Ÿ��:�/���,'��}?��|W��(o��?������$���?���=��S��ҴŻ�.л�{ڻ��ה��`��'�(���d
�����w�����=�� �z�$���(���,�#�0�R�4�k�8�U�<�io@�k+D���G��}K��O���R��$V�ҜY��]��p`���c�R"g��nj�)�m�1�p�)t�gZw�R�z��}�9e���򁼣}��v��������Ք�����������*���v��`���)����u��i얼b���֙��J������u0��^����������$���He��զ��D��8���k#����������p���߰�O��<����-���������|����]���ν��  �  ��N=�M=0/M=�uL=��K=3K=hFJ==�I=��H=|H=�VG=��F=
�E=�E=�^D=Z�C=#�B=/B=y\A=�@=��?=<?=�L>=��==;�<=��;=-;=b:=ٕ9=4�8=.�7=�(7=�V6=��5=<�4=��3=��2=�!2=;D1=�d0=�/=��.=�-=r�,=6�+=�*=� *=r)=�(=�'=�&=e%=$=� #=Q�!=�� =��=ڨ=��=ja=c6=J=�=��=�V=�=��=�v=� =x�=�d=�=��=f 
=t�=-=n�=�$=��=�=���<��<�p�<�)�<<��<N��<`"�<Ǻ�<�K�<���<-Y�<���<�L�<���<�)�<-��<���<-O�<!��<*��<�N�<y��<<�<�.�<&t�<���<��<s5�<�q�<���<'�<t�<�U�<��<���<P��<'Yz<m�r<[.k<ƙc<�\<�tT<��L<WE<��=<�C6<�.<�='<��<�H<=�<g	<��<�9�;~��;���;*C�;Q��;E�;��;ʑ�;�V�;df;�HJ;�].;��;	E�:q��:D��:r�:,�59��o��B$������Ÿ�v;�b���-'��~?��}W�W)o��@���������K@���=������Ż�.л+|ڻ<��p�`��� ����rd
����_w����a=��� �4�$���(�G�,���0���4�F�8�'�<�2o@�J+D�~�G�~K��O���R��$V���Y��]�5q`��c�x"g�Noj�_�m�u�p��)t��Zw���z���}�Le���򁼶}����2�������������r���������J��H�������u��C얼�a���֙��J��ӽ��U0��N�������������9e��.զ��D��C���~#����������p��఼O��e����-��:�������|��1��]���ν��  �  ��N=��M=2/M=�uL=��K=.K=pFJ=@�I=��H=�H=�VG=ęF= �E=�E=�^D=q�C=6�B=;B=�\A=��@=��?==?=�L>=��===�<=��;=
-;=b:=Ε9=.�8=�7=�(7=pV6=��5=+�4=��3=��2=y!2=2D1=�d0=�/=��.=�-=y�,=7�+=�*=� *=s)=�(=�'=�&=p%= $=� #=i�!=�� =��=�=��=xa=l6=X=�=��=�V=�=��=�v=� =n�={d=��=�=[ 
=Z�=�,=X�=�$=��=�=���<��<�p�<�)�<4��<U��<]"�<ʺ�<�K�<���<+Y�<��<�L�<	��<�)�<L��<��<:O�<G��<Y��<�N�<���<T�< /�</t�<̶�<��<k5�<�q�<ì�<3�<Z�<�U�<���<���<5��<�Xz<1�r<
.k<��c<8\<qtT<~�L<�VE<��=<�C6<��.<�='<��<�H<*�<1g	<��<(:�;ރ�;���;�C�;��;�E�;��;���;�W�;�df;nIJ;r^.;إ;�E�:���:���:��:�59�o�DB$�л��|Ƹ�!=뺦���.'��?��~W�t*o��@����������@��L>�����_�Żu.л|ڻ��仩��t`��� �ۼ�1d
����"w�����<�j� ��$�7�(��,���0���4�	�8��<�(o@�<+D���G��}K��O�r�R��$V�(�Y��]�rq`�9�c��"g��oj���m���p�*t��Zw���z��}�[e���򁼸}��s��0������Δ�����q���v������8��-��������u��5얼�a���֙��J������>0��-�������������Be��"զ��D��7����#��Ȓ�����	q��఼HO�������-��W���
���|��B��]���ν��  �  y�N=y�M=#/M=�uL=��K=8K={FJ=B�I=��H=�H=�VG=֙F=$�E=�E=�^D=w�C=<�B=MB=�\A=�@=��?=<?= M>=��==A�<=��;=�,;=b:=Õ9='�8=�7=�(7=`V6=��5=&�4=��3=��2=i!2=&D1=�d0=؂/=��.=ַ-=j�,=,�+=�*=� *=�)=�(=�'=�&=o%=.$=� #=m�!=�� =��=��=��=�a=k6=a=�=��=�V=�=��=�v=� =a�=rd=��=ؑ=M 
=F�=�,=I�=w$=��=�=���<Ԯ�<�p�<�)�<��</��<L"�<κ�<�K�<���<&Y�<(��<M�<��<�)�<\��< ��<RO�<T��<`��<�N�<���<V�<8/�<7t�<߶�<4��<o5�<�q�<���<�<F�<�U�<㋈<���<��<�Xz< �r<�-k<r�c<
\<9tT<[�L<�VE<��=<rC6<ʾ.<�='<��<�H<P�<^g	<�<�:�;��;U��;D�;7��;F�;p�;Ӓ�;�W�;7ff;�IJ;�^.;ʦ;�E�:��:���:�:�59��o��D$�޼��Ǹ�g>�����/'��?��~W�Q+o��@���4���@���>������Ż�.лm|ڻڝ仞���_��� ����d
�����v�\���<�L� �ݹ$�(�(���,�j�0���4���8��<�o@��*D���G��}K��O���R�%V�C�Y� ]��q`�g�c�#g��oj�ߴm���p�*t�1[w�݅z��}�ke�����}�����=������Ŕ�����s���[��쏏�/���������xu��얼�a���֙�oJ������=0��������t�������>e��"զ��D��M����#��В����q��8఼aO�������-��`��� ��}��R��]���ν��  �  }�N=|�M=,/M=�uL=��K=3K=pFJ=J�I=��H=�H=�VG=ٙF=+�E=�E=_D=}�C=D�B=MB=�\A=�@=��?=B?=�L>=��==;�<=��;=-;=b:=ĕ9=�8=�7=~(7=^V6=��5=�4=��3=��2=k!2=D1=�d0=҂/=��.=ܷ-=o�,=4�+=�*=� *=x)=�(=�'=�&=~%=/$=� #=s�!=�� =��=��=��=�a=z6=`=$�=��=�V=�=��=�v=� =g�=nd=��=Ց=C 
=G�=�,=<�=g$=~�=�=���<̮�<�p�<�)�<!��<=��<X"�<���<�K�<���<-Y�<1��<M�<,��<�)�<l��<,��<}O�<o��<o��<�N�<���<q�<9/�<Gt�<϶�<(��<j5�<�q�<���<%�<M�<yU�<׋�<���<��<�Xz<��r<�-k</�c<�\<$tT<2�L<�VE<�=<~C6<׾.<�='<��<�H<=�<5g	<$�<�:�;T��;���;:D�;w��;jF�;*�;��;$X�;Cff;�JJ;]_.;/�;�F�:���:���:�:׆59
�o�'C$�����Iȸ��>뺮���/'�n�?��W��+o�xA������r��A���>��0��w�Ż�.л(|ڻ�仦��D`��� ����d
�D���v�3���<�� ���$��(���,�q�0���4���8�ǥ<�"o@�++D���G��}K��O���R��$V�O�Y�]��q`���c�#g��oj��m��p�M*t�.[w��z�%�}�~e�����}�����/������ǔ�����j���P��珏���	�������ku���떼�a��r֙�bJ������"0���������������De��$զ��D��F����#��㒬���'q��F఼eO������.������(�� }��e�^��Ͻ��  �  x�N=n�M=&/M=�uL=��K=@K=yFJ=S�I=��H=�H=�VG=ۙF=8�E=�E=_D=|�C=P�B=KB=�\A=�@=��?=L?=�L>=��==>�<=��;=�,;=�a:=9=�8=�7=y(7=`V6=��5=�4=��3=��2=k!2=D1=�d0=ւ/=��.=շ-=b�,=1�+=
�*=� *=�)=�(=�'=�&=�%=-$=� #=v�!=�� =��=��=��=�a=�6=W=%�=��=�V=�=��=�v=� =]�=jd=��=֑=; 
=I�=�,=H�=k$=w�=�=���<ծ�<�p�<�)�<��<)��<R"�<���<�K�<���<EY�<%��<�L�<A��<�)�<���<+��<hO�<f��<���<�N�<���<�<&/�<Ut�<ⶦ<?��<z5�<�q�<���<	�<B�<tU�<勈<���<��<�Xz<��r<�-k<$�c<�\<tT<.�L<�VE<t�=<lC6<��.<�='<��<�H<t�<Yg	<F�<O:�;n��;���;JD�;Ἲ;PF�;��;��;�X�;*ff;WKJ;8_.;��;�G�:e��:���:��:�59C�o�uF$�׼��+ȸ��=���r/'��?��W��*o��A���������A���>��B����Ż!/лB|ڻ��6��`��� ����%d
����v����<�+� ���$��(���,�{�0�`�4� �8�å<��n@�+D�Y�G��}K��O�͢R�%V�\�Y�]��q`���c�#g��oj�شm��p�k*t�[w�&�z��}�|e�����}�����5�������������R���]��򏏼�
���������mu��얼�a��_֙�_J������0��'���u��r�������4e��(զ��D��a����#��璬� ��'q��L఼hO�������-������/��#}��g��]��Ͻ��  �  }�N=|�M=,/M=�uL=��K=3K=pFJ=J�I=��H=�H=�VG=ٙF=+�E=�E=_D=}�C=D�B=MB=�\A=�@=��?=B?=�L>=��==;�<=��;=-;=b:=ĕ9=�8=�7=~(7=^V6=��5=�4=��3=��2=k!2=D1=�d0=҂/=��.=ܷ-=o�,=4�+=�*=� *=x)=�(=�'=�&=~%=/$=� #=s�!=�� =��=��=��=�a=z6=`=$�=��=�V=�=��=�v=� =g�=nd=��=֑=C 
=G�=�,=<�=g$=�=�=���<ͮ�<�p�<�)�<"��<>��<Y"�<���<�K�<���<.Y�<2��<M�<,��<�)�<l��<,��<~O�<o��<o��<�N�<���<q�<9/�<Ft�<ζ�<(��<i5�<�q�<���<$�<M�<xU�<׋�<���<��<�Xz<��r<�-k</�c<�\<$tT<3�L<�VE<��=<C6<ؾ.<�='<��<�H<?�<6g	<%�<�:�;V��;���;;D�;x��;jF�;*�;��;"X�;?ff;�JJ;W_.;)�;�F�:���:���:�:J�59��o�LC$�����[ȸ��>뺷���/'�v�?��W��+o�{A�� �u��A���>��2��y�Ż�.л*|ڻ�仨��E`��� ����d
�E���v�3���<�� ���$��(���,�q�0���4���8�ǥ<�#o@�++D���G��}K��O���R��$V�O�Y�]��q`���c�#g��oj��m��p�M*t�.[w��z�%�}�~e�����}�����/������ǔ�����j���P��珏���	�������ku���떼�a��r֙�bJ������"0���������������De��$զ��D��F����#��㒬���'q��F఼eO������.������(�� }��e�^��Ͻ��  �  y�N=y�M=#/M=�uL=��K=8K={FJ=B�I=��H=�H=�VG=֙F=$�E=�E=�^D=w�C=<�B=MB=�\A=�@=��?=<?= M>=��==A�<=��;=�,;=b:=Õ9='�8=�7=�(7=`V6=��5=&�4=��3=��2=i!2=&D1=�d0=؂/=��.=ַ-=j�,=,�+=�*=� *=�)=�(=�'=�&=o%=.$=� #=m�!=�� =��=��=��=�a=k6=a=�=��=�V=�=��=�v=� =b�=rd=��=ّ=N 
=F�=�,=I�=x$=��=�=���<֮�<�p�<�)�<��<1��<N"�<Ϻ�<�K�<���<(Y�<)��<M�<��<�)�<\��<!��<RO�<T��<_��<�N�<���<U�<7/�<5t�<޶�<3��<n5�<�q�<���<�<E�<�U�<⋈<���<��<�Xz< �r<�-k<r�c<\<:tT<]�L<�VE<��=<tC6<̾.<�='<��<�H<S�<`g	<�<�:�;���;X��;D�;8��;F�;o�;ђ�;�W�;0ff;�IJ;�^.;��;�E�:���:���:پ:�59��o��D$����AǸ��>����/'��?�W�_+o��@���:���@���>������Ż�.лp|ڻݝ仠���_��� ����d
�����v�\���<�L� �ݹ$�(�(���,�j�0���4���8��<�o@��*D���G��}K��O���R�%V�C�Y� ]��q`�g�c�#g��oj�ߴm���p�*t�1[w�݅z��}�ke�����}�����=������Ŕ�����s���[��쏏�/���������xu��얼�a���֙�oJ������=0��������t�������>e��"զ��D��M����#��В����q��8఼aO�������-��`��� ��}��R��]���ν��  �  ��N=��M=2/M=�uL=��K=.K=pFJ=@�I=��H=�H=�VG=ęF= �E=�E=�^D=q�C=6�B=;B=�\A=��@=��?==?=�L>=��===�<=��;=
-;=b:=Ε9=.�8=�7=�(7=pV6=��5=+�4=��3=��2=y!2=2D1=�d0=�/=��.=�-=y�,=7�+=�*=� *=s)=�(=�'=�&=p%= $=� #=i�!=�� =��=�=��=ya=l6=X=�=��=�V=�=��=�v=� =o�=|d=��=�=\ 
=[�=�,=Y�=�$=��=�=���<��<�p�<�)�<7��<X��<`"�<̺�<�K�<���<-Y�<��<�L�<��<�)�<M��<��<:O�<G��<X��<�N�<���<S�</�<-t�<˶�<��<i5�<�q�<���<1�<X�<�U�<���<���<4��<�Xz<0�r<
.k<��c<9\<stT<��L<�VE<��=<�C6<��.<�='<��<�H<.�<4g	<��<.:�;��;���;�C�;��;�E�;��;���;�W�;�df;bIJ;c^.;ǥ;`E�:ͭ�:���:$�:i�59��o��B$�����Ƹ�R=뺾���.'��?��~W��*o��@����������@��R>�����e�Żz.л"|ڻ��们��w`��� �ܼ�1d
����"w�����<�k� ��$�7�(��,���0���4�	�8��<�(o@�<+D���G��}K��O�r�R��$V�(�Y��]�rq`�9�c��"g��oj���m���p�*t��Zw���z��}�[e���򁼸}��s��0������Δ�����q���v������8��-��������u��5얼�a���֙��J������>0��-�������������Be��"զ��D��7����#��Ȓ�����	q��఼HO�������-��W���
���|��B��]���ν��  �  ��N=�M=0/M=�uL=��K=3K=hFJ==�I=��H=|H=�VG=��F=
�E=�E=�^D=Z�C=#�B=/B=y\A=�@=��?=<?=�L>=��==;�<=��;=-;=b:=ٕ9=4�8=.�7=�(7=�V6=��5=<�4=��3=��2=�!2=;D1=�d0=�/=��.=�-=r�,=6�+=�*=� *=r)=�(=�'=�&=e%=$=� #=Q�!=�� =��=ڨ=��=ka=c6=J=�=��=�V=�=��=�v=� =x�=�d=�=��=g 
=u�=-=p�=�$=��=�=���<��<�p�<�)�<?��<Q��<d"�<ʺ�<�K�<���<0Y�<���<�L�<���<�)�<.��<���<-O�<!��<)��<�N�<x��<;�<�.�<$t�<���<��<q5�<�q�<���<$�<r�<�U�<��<���<O��<&Yz<m�r<[.k<Ǚc<�\<�tT<��L<WE<��=<�C6<�.<�='<��<�H<B�<g	<��<�9�;���;���;-C�;S��;E�;��;Ǒ�;�V�;�cf;�HJ;�].;ߤ;�D�:>��:��: �:Q~59h�o�mC$�����7Ƹ��;����-'��~?��}W�p)o��@���������T@��>�����#�Ż�.л1|ڻA��t�`��� ����td
����`w����b=��� �5�$���(�G�,���0���4�F�8�(�<�2o@�J+D�~�G�~K��O���R��$V���Y��]�5q`��c�x"g�Noj�_�m�u�p��)t��Zw���z���}�Le���򁼶}����2�������������r���������J��H�������u��C얼�a���֙��J��ӽ��U0��N�������������9e��.զ��D��C���~#����������p��఼O��e����-��:�������|��1��]���ν��  �  ��N=��M=6/M=�uL=��K=)K=cFJ=.�I=��H=mH=�VG=��F=��E=�E=�^D=I�C=�B="B=d\A=�@=y�?=,?=�L>=��==9�<=��;=	-;=b:=�9=?�8=9�7=�(7=�V6=̂5=N�4= �3=��2=�!2=LD1=�d0=��/=��.=��-=u�,=A�+=�*=� *=i)=�(=�'=�&=S%=$=� #=A�!=�� =t�=ʨ=}�=_a=P6=C=�=��=�V=�=��=�v=� =��=�d=�=�=} 
=��='-=��=�$=��=�=,��<9��<q�<
*�<Z��<b��<�"�<κ�<�K�<���<Y�<���<�L�<ҽ�<�)�<��<���<O�< ��<��<mN�<R��<�<�.�<t�<���<	��<`5�<�q�<̬�</�<��<�U�<(��<<t��<WYz<��r<�.k<�c<�\<�tT<�L<>WE<�=<D6<�.<>'<�<�H<�<g	<��<c9�;��;���;�B�;���;�D�;�;(��;LV�;�bf;GJ;�\.;�;nB�:V��:.��:h�:k�59�o�GB$�(���EŸ��:�P���,'��}?��|W��(o��?������/���?���=��[��ٴŻ�.л�{ڻ��۔��`��)�*���d
� ���w�����=�� �{�$���(���,�#�0�R�4�l�8�U�<�io@�k+D���G��}K��O���R��$V�ҜY��]��p`���c�R"g��nj�)�m�1�p�)t�gZw�R�z��}�9e���򁼣}��v��������Ք�����������*���v��`���)����u��i얼b���֙��J������u0��^����������$���He��զ��D��8���k#����������p���߰�O��<����-���������|����]���ν��  �  ��N=��M=7/M=�uL=��K=#K=_FJ=%�I=~�H=]H=�VG=��F=��E=�E=�^D=9�C=��B=B=W\A=ԙ@=p�?=%?=�L>=��==:�<=��;=-;=(b:=�9=Q�8=F�7=�(7=�V6=��5=e�4=�3=��2=�!2=`D1=�d0=
�/=Ȟ.=��-=��,==�+=�*=� *=g)=�(=�'=�&=F%=�$=� #=2�!=|� =_�=��=f�=Pa=F6=6= �=��=�V=�=��=�v=� =��=�d=&�=�=� 
=��=A-=��=�$=ؘ=�=\��<Z��<3q�<!*�<~��<w��<�"�<׺�<�K�<���<Y�<���<�L�<���<d)�<��<���<�N�<ܧ�<���<@N�<5��<��<�.�<�s�<���<���<_5�<�q�<ɬ�<M�<��<�U�<J��<<���<�Yz<$�r<�.k<��c<\<AuT<@�L<�WE<T�=<D6<N�.<>'<�<�H<�<�f	<��<
9�;}��;s��;�A�;	��;�C�;*��;���;U�;�af;�EJ;K[.;;�;A�:{��:-��:��:\59��o�g?$�����fø�y9�Y��#,'��|?��{W��'o�W?��Q�������?��D=������ŻQ.л|ڻ$�����`��8�N���d
�8���w�[���=�?� �պ$�&�(���,�d�0���4���8�y�<�zo@�s+D���G��}K��O�Y�R�w$V���Y�E]��p`���c�"g��nj�ֳm���p�.)t�+Zw��z�N�}�e���򁼇}��h��!������ޔ�����������I����������V����u���얼8b���֙��J������0��t����������-���He�� զ��D�����^#����������p���߰��N�����p-��✶�����|���캼�]���ν��  �  ��N=��M=</M=�uL=��K=!K=PFJ= �I=o�H=NH=�VG=��F=��E=�E=�^D=#�C=��B=�B=K\A=Ù@=c�?=?=�L>=��==;�<=��;=-;=,b:=�9=\�8=V�7=�(7=�V6=�5=w�4=,�3=��2=�!2=rD1=�d0=�/=О.=�-=��,=A�+=�*=� *=`)=�(=z'=�&=;%=�$=� #=�!=h� =K�=��=Y�==a=<6='=��=��=�V=�=��=�v=� =��=�d=9�=,�=� 
=��=T-=��=�$=�=	=���<���<Vq�<9*�<���<���<�"�<޺�<�K�<���<Y�<���<�L�<���<@)�<Ǐ�<~��<�N�<���<���< N�<��<��<�.�<�s�<���<���<c5�<�q�<Ѭ�<S�<��<�U�<l��<;<���<�Yz<i�r<J/k<ƚc<l\<�uT<�L<�WE<��=<CD6<_�.<->'<�<�H<��<�f	<v�<�8�;���;���;rA�;o��;C�;�ߝ;ˏ�;�T�;J`f;EJ;Z.;,�;�?�:��::�:`{59��o�5?$�&���^¸��7뺧���*'��{?��zW�J&o��>��������(?���<�����{�Ż<.л�{ڻ3��Ȕ�6a��p�r��e
�i��,x����A>��� �,�$���(�"�,���0���4���8���<��o@��+D���G��}K��O�P�R�e$V���Y�
]��p`�>�c��!g�jnj�z�m���p��(t��Yw�΄z��}��d��r򁼀}��d��"������֔��)���������k����������s���v���얼fb��"י�	K��6����0���������Ǆ��7���Be��!զ��D�����O#��u���|���p���߰��N���:-����|��q|���캼r]���ν��  �  ��N=��M=G/M=�uL=��K=K=IFJ=�I=c�H=EH=�VG=x�F=��E=yE=�^D=�C=��B=�B=7\A=��@=W�?=?=�L>=��==2�<=��;=-;=4b:=��9=d�8=f�7=�(7=�V6=�5=��4=?�3=�2=�!2=~D1=�d0=#�/=ڞ.=�-=��,=N�+=�*=� *=[)=�(=p'=�&=-%=�$=� #=�!=Y� =>�=��=Q�=,a=-6= =��=~�=�V=�=��=�v=� =��=�d=F�=D�=� 
=ũ=k-=̫=�$=�==���<���<mq�<[*�<���<���<�"�<պ�<�K�<���<�X�<���<�L�<���<)�<���<S��<�N�<���<���<N�<囵<��<�.�<�s�<s��<���<M5�<�q�<笗<Y�<��<�U�<���<e<���<<Zz<��r<�/k<�c<�\<�uT<��L<XE<��=<�D6<v�.<[>'<-�<~H<��<�f	<M�<+8�;���;9��;�@�;�;mB�;ߝ;	��;�T�;�^f;�CJ;?Y.;>�;>�:��:p��:2�:{�59�o�&>$���������36뺵��&*'��z?��yW�<%o�i>��3�������>���<������Ż.л�{ڻ?��7��ca�������@e
����x�����>�څ �g�$���(�I�,��0���4��8�Ʀ<��o@��+D���G�~K�jO�3�R�+$V�a�Y��
]�@p`��c�z!g�nj�3�m�F�p��(t��Yw���z�̩}��d��X�m}��Q��������ꔉ�2��Õ�����������΅������Jv���얼�b��@י�'K��a����0���������ք��>���We��զ��D�����0#��a���c��op��߰��N��ͽ��-������Y��X|���캼U]���ν��  �  ��N=��M=A/M=�uL=��K=K=LFJ=	�I=\�H=7H=�VG=h�F=��E=jE=�^D=��C=��B=�B=+\A=��@=P�?=?=�L>=��==9�<=��;=-;=9b:=�9=u�8=r�7=�(7=�V6=�5=��4=G�3=�2=�!2=�D1=e0=1�/=�.=�-=��,=E�+=�*=� *=c)=�(=f'=�&=%=�$=r #=��!=G� =,�=��=;�=&a=6==��=z�=�V=�=��=�v=� =��=�d=X�=R�=� 
=ԩ=�-=۫=%=�=(=���<ȯ�<�q�<l*�<���<���<�"�<��<�K�<���<�X�<���<nL�<j��<)�<���<9��<pN�<i��<w��<�M�<כ�<��<�.�<�s�<t��<���<Q5�<�q�<ج�<l�<��<V�<���<|<���<�Zz<�r<�/k<f�c<\<vT<�L<8XE<��=<�D6<��.<F>'<*�<�H<��<�f	<�<�7�;3��;���;W@�;A��;�A�;iޝ;���;�S�;^f;�BJ;UX.;��;;<�:���:B��::�:%x59��o�d=$�y�����5�����)'��y?��xW��$o��=��˾��g��G>��1<��R���Ż�-л�{ڻ��3��0a����Ƚ�ce
�����x����>�$� ���$��(���,� �0�4�4�9�8��<��o@��+D���G��}K��O�#�R�$$V�E�Y��
]�p`���c�L!g��mj��m��p�G(t�mYw�R�z���}��d��M�d}��O��������蔉�#��ؕ��������������������ev��햼�b��gי�KK��o����0��������Ԅ��7���Re��զ��D������,#��I���M��Xp��i߰�qN������-��w���/��D|���캼?]��gν��  �  ��N=��M=I/M=�uL=��K=K=BFJ= �I=X�H=)H=�VG=Z�F=��E=eE=z^D=��C=��B=�B=#\A=��@=K�?=�?=�L>=��==:�<=��;='-;=Ab:=�9=��8=r�7=�(7=�V6=�5=��4=R�3=!�2=�!2=�D1=
e0=:�/=�.=�-=��,=I�+=�*=� *=R)=�(=^'=�&=%=�$=a #=��!=@� ="�=��=*�=a=6==��=q�=�V=�=��=�v=!=��=�d=d�=U�=� 
=�=�-=�=%=$�=9=���<̯�<�q�<}*�<���<ł�<�"�<��<�K�<���<�X�<���<XL�<[��<�(�<i��<3��<RN�<_��<h��<�M�<ț�<��<|.�<�s�<^��<���<H5�<�q�<嬗<��<��<,V�<���<�<��<�Zz<)�r<�/k<��c<$\<NvT<2�L<EXE<�=<�D6<Ϳ.<j>'<<�<�H<��<|f	<��<�7�;���;���;�?�;췺;�A�;�ݝ;b��;@S�;.]f;BJ;_W.;/�;�:�:���:C��:�:`w59��o��;$�0���ʾ��95�V���('�jy?�`xW�7$o��=���������4>���;������Żz-л�{ڻ��r�a�������e
����x�g���>�D� �߻$��(���,�L�0�\�4�_�8��<�p@��+D���G��}K��O��R�!$V��Y��
]�p`���c�!g��mj��m���p�8(t�6Yw��z���}��d��A�W}��2�������� ���?��알�������������������lv�� 햼�b��vי�jK��}����0��Ƣ����ꄢ�W���\e��զ��D��ݳ��,#��0���D��Hp��D߰�fN�������,��i���'�� |��|캼:]��Nν��  �  ¡N=��M=F/M=�uL=��K=K=FFJ=�I=N�H=%H=~VG=V�F=��E=UE=p^D=�C=��B=�B=\A=��@=C�?=?=�L>=��==8�<=��;= -;=:b:=�9=��8=��7=�(7=�V6=%�5=��4=h�3='�2=�!2=�D1=e0=;�/=��.=�-=��,=I�+=�*=� *=Z)=�(=]'=�&=%=�$=c #=��!=1� =�=u�=-�=a=6=	=��=y�=�V=�=��=�v=!=��=�d=e�=f�=� 
=�=�-=��=#%=-�=D=���<��<�q�<�*�<���<���<�"�<��<�K�<���<�X�<���<ML�<T��<�(�<l��<��<?N�<B��<W��<�M�<���<��<g.�<�s�<g��<���<N5�<�q�<ଗ<o�<��<6V�<���<�<��<�Zz<H�r<E0k<��c<D\<ZvT<U�L<oXE<+�=<�D6<��.<]>'<*�<�H<��<�f	<��<n7�;���;S��;�?�;���;2A�;�ݝ;ύ�;/S�;�\f;�AJ;�V.;��;�:�:��:9��:�:�s59�o��=$�`���꾸��3�!��l('��x?��wW��"o�q=��E�������=���;�������Ż�-л�{ڻD��8��a�������e
����x�`��?��� ��$�W�(���,�s�0�a�4�z�8��<��o@��+D���G�~K��O��R�$V���Y��
]��o`���c�� g��mj���m���p�(t�Yw��z�f�}��d��1�c}��E��������𔉼6��ᕌ������� ��	��������v��3햼�b���י�oK������1��ۢ����ᄢ�D���Ue��զ��D������ #��&���6��2p��C߰�VN�������,��W�����|��k캼&]��Hν��  �  ��N=P�M=�5M=�|L=��K=
K=PJ=��I=��H=�H=�cG=��F=��E=�-E=�oD=[�C=M�B=�2B=rA=Ű@=��?=�+?=�g>=�==��<=<=�M;=v�:=Թ9=��8=u 8=�Q7=,�6=,�5=t�4=�4=�.3=YU2=�y1=k�0=��/=I�.=��-=-=�#,=�6+=sF*=S)=^\(=8b'=sd&=�b%=�]$=+T#=�F"=�4!=a =R=��=�=r�=�f=�2=!�=-�=�u=�+=��=�=�*=��=�b="�=��
=�	=^�=s=&�=��=�b=���<�]�<!�<���<]{�<��<���<�L�<���<]�<��<eR�<���<W/�<c��<���<�R�<���<&��<�M�<���<��<a(�<k�<,��<��<8$�<�]�<Y��<o˗< �<�3�<�e�<���<�Ȅ<:��<�Sz<1�r<�k<Wwc<��[<�>T<C�L<�E<�x=<��5<�W.<��&<�E<�<SE<��<eZ<���;��;�S�;Y��;�	�;y~�;��;á�;c�~;�2b;��E;�);��;1��:�ŭ:{�n:��:K/�8�����:�<���ĺ)2��ޣ�Q]-��E�I�]���u����,���b��`���Ǒ��e��ɻ�ӻ?�ݻB��u�񻨦�����qX�W��\�����i�����!�+&�H*�|S.��N2�H:6��:���=� �A�.XE�u�H�ƘL�i'P���S��$W�v�Z���]��Wa���d���g��=k�2{n�űq���t��x��/{��M~������=���Ń��K��|φ��Q���щ�^P��X͌��H��Ï��;������3*�������������@���l��)ݜ��M�������,��Л��\
���x���榼PT��©��/�����q
���w��e尼�R������:.��D���^
���x���纼�V��Jƽ��  �  ��N=L�M=�5M=�|L=��K=
K=PJ=��I=��H=�H=�cG=��F=��E=�-E=�oD=`�C=P�B=�2B=rA=��@=��?=�+?=�g>=��==�<=�<=�M;=m�:=˹9=��8=j 8=�Q7=.�6=*�5=w�4= 4=�.3=WU2=�y1=b�0=��/=E�.=v�-=-=�#,=�6+=|F*=S)=e\(=;b'=qd&=�b%=�]$=/T#=�F"=�4!=Q =]=��=
�=k�=�f=�2=%�=7�=�u=�+=��=�=�*=��=�b=�=Ń
=�	=_�=t=)�=��=�b=���<�]�<,�<���<I{�<|�<���<�L�<���<1]�<��<qR�<���<N/�<n��<���<�R�<���<��<�M�<���<��<R(�<k�<0��<��<Q$�<�]�<V��<S˗<���<r3�<�e�<���<�Ȅ<J��<�Sz<D�r<�k<hwc<��[<�>T<?�L<�E<�x=<��5<�W.<��&<�E<5�<�E<�<fZ<���;��;�S�;w��;�	�;�~�;E�;硍;��~;3b;��E;��);��;V��:�ƭ:��n:�:}%�8�����:�{=��_�ĺv3����� ]-��E��]�i�u����9���b����������e��_ɻ�ӻ��ݻ9��*��C���{��gX�\��������i����&�!�Q+&��G*�pS.��N2�f:6��:���=��A�XE�R�H���L��'P���S�%W���Z���]��Wa�~�d���g��=k�({n���q���t��x��/{��M~������=���Ń��K���φ�|Q���щ�KP��U͌��H��$Ï�<������0*������!������.���l��$ݜ��M��z����,������D
���x���榼lT��
©��/�����y
���w��U尼�R������<.��;���^
���x���纼�V��Dƽ��  �  ��N=V�M=�5M=�|L=��K=
K=PJ=��I=��H=�H=�cG=��F=��E=�-E=�oD=u�C=U�B=�2B=rA=ɰ@=��?=�+?=�g>=�==�<=�<=�M;=s�:=¹9=��8=\ 8=�Q7=�6=�5=m�4=�4=�.3=BU2=�y1=T�0=��/==�.=s�-=-=�#,=�6+=sF*=S)=c\(=Ab'=�d&=�b%=�]$=1T#=�F"=�4!=a =q=��=�=t�=�f=�2=#�=3�=�u=�+=��= �=�*=��=�b=�=��
=�	=S�=`=�=��=�b=���<x]�<&�<���<J{�<��<���<�L�<���<.]�<��<�R�<���<c/�<���<���<�R�<���<E��<�M�<	��<��<`(�<,k�<7��<��<F$�<�]�<_��<\˗< �<d3�<�e�<~��<�Ȅ<2��<1Sz<$�r<Gk<Dwc<8�[<�>T<�L<�E<�x=<��5<X.<��&<�E<�<`E<
�<jZ<Q��;��;;T�;���;
�;0�;��;���;�~;4b;�E;��);��;���:Cǭ:ǲn:��:p)�8����:�b>��4�ĺ�4�����^-���E���]�f�u��������b���������Ye��qɻ��ӻ��ݻ��g��e���~��KX� ��]��>��i�x����!�+&��G*�kS.��N2�;:6��:���=��A�XE�u�H���L��'P�O�S�%W���Z���]�Xa���d�3�g��=k�n{n��q���t��x��/{�8N~������=���Ń��K���φ�Q���щ�KP��S͌��H��Ï��;������+*������ ��y�������k��ݜ��M��]����,������Q
���x���榼dT�������/������
���w��m尼�R������a.��K����
���x���纼�V��Jƽ��  �  ��N=E�M=�5M=�|L=��K=
K=PJ=��I=��H=�H=�cG=ŧF=�E=�-E=�oD={�C=f�B=�2B=rA=հ@=��?=�+?=�g>=�==�<=�<=�M;=i�:=��9=��8=W 8=|Q7=�6=�5=_�4=�4=�.3=6U2=�y1=M�0=u�/=5�.=n�-=�-=�#,=�6+=vF*="S)=m\(=Gb'=�d&=	c%=�]$=AT#=�F"=�4!=o =s=��=$�=�=�f=�2=+�=>�=�u=�+=��=�=�*=��=�b=��=��
=�	=E�=O=�=��=�b=i��<f]�<�<{��<1{�<]�<}��<�L�<���<A]�<��<�R�<���<w/�<���<���<�R�<Ī�<Y��<N�<,��<��<|(�<5k�<I��<��<[$�<�]�<]��<O˗<���<Z3�<�e�<m��<zȄ<��<�Rz<�r<k<wc<�[<~>T<�L<gE<~x=<k�5<�W.<��&<�E<&�<�E<6�<�Z<k��;)�;�T�;D��;�
�;~�;b�;ࢍ;<�~;�4b;J�E;~�);�;h��:ɭ:��n:5�:0�8�����:�?����ĺR5��u���^-�@�E�^�]�(�u�/���(��c��6�������e���ɻU�ӻ��ݻ��E������U��/X� ��)���]i�e����!��*&�G*�&S.�eN2�	:6��:���=��A��WE�h�H���L��'P���S�"%W�ɔZ���]�'Xa�Ĭd�g�g�>k��{n�%�q��t��x��/{�MN~�ɳ��>���Ń��K���φ�{Q���щ�4P��=͌��H�����;��~���*��|������e�������k���ܜ�qM��U����,������<
���x���榼rT��©��/��$����
��x���尼S������z.��f����
��y���纼�V��cƽ��  �  ��N==�M=�5M=�|L=��K=
K=PJ=ŕI=��H=�H=dG=ڧF=&�E=�-E=pD=��C=��B=�2B=.rA=�@=��?=�+?=�g>=��==�<=�<=�M;=a�:=��9=��8=D 8=dQ7=�6=��5=C�4=�4=p.3=&U2=�y1=;�0=d�/='�.=h�-=�-=�#,=�6+=}F*=#S)=q\(=Qb'=�d&=c%=�]$=_T#=�F"=�4!=� =�=��=,�=��=�f=�2=/�=<�=�u=�+=��=��=�*=t�=�b=��=��
=�	=#�=3=�=b�=�b=.��<9]�<��<a��<{�<U�<y��<�L�<���<7]�<#��<�R�<��<�/�<���<���<S�<��<���<FN�<_��<�<�(�<Qk�<_��<��<e$�<�]�<W��<U˗<���<S3�<�e�<G��<MȄ<���<�Rz<r�r<�k<�vc<��[<@>T<��L<E<3x=<U�5<�W.<��&<�E<.�<�E<2�<�Z<���;��;�T�;���;v�;-��;=�;���;2�~;6b;~�E;&�); ;	��:oɭ:��n:��:89�8r�����:�`?��"�ĺ17�����v_-���E���]�W�u��������c�����������e���ɻr�ӻ��ݻ2�������?��X����Ո����h���L�!�q*&�"G*��R.�>N2��96�W:�~�=�ϤA��WE�K�H���L��'P���S�>%W���Z�4�]�lXa��d���g��>k� |n���q��t�6x�30{��N~�賀�>���Ń��K���φ��Q���щ�7P��.͌��H�����;��g����)��U������<��������k���ܜ�AM��;����,������5
���x���榼mT��)©��/��D����
��3x���尼9S�������.�������
��$y���纼W���ƽ��  �  p�N=8�M=�5M=�|L=��K=
K=)PJ=ՕI=�H=�H= dG=�F=5�E=�-E="pD=��C=��B=�2B=GrA=��@=��?=�+?=�g>=�==�<=�<=�M;=V�:=��9=��8=4 8=QQ7=�6=�5=1�4=�4=].3=U2=�y1=#�0=\�/=�.=W�-=�-=�#,=�6+=�F*=&S)=�\(=ab'=�d&=0c%=�]$=kT#=�F"=�4!=� =�=��=D�=��=�f=�2=;�=?�=�u=+=��=��=�*=`�=}b=��=w�
=�	=
�==ς=G�=�b=���<	]�<��<2��<�z�<H�<\��<�L�<���<F]�<<��<�R�<��<�/�<��<���<IS�<!��<���<iN�<~��<4�<�(�<uk�<���<�<p$�<�]�<O��<G˗<���<.3�<�e�<2��<Ȅ<���<NRz<!�r<Nk<?vc<E�[<�=T<-�L<�E<x=<�5<zW.<��&<�E<4�<�E<f�<�Z<a��;d�;�U�;���;�;)��;	�;���;I�~;�7b;H�E;�);|;���:b˭:c�n:��:�/�8����z�:�6A��v�ĺ�8������`-���E���]���u�����1	��Nd��f�������Hf��/ɻf�ӻ��ݻ/�������������W����������h������!�*&��F*�nR.��M2�l96�:�<�=���A��WE�&�H���L��'P���S�%W�5�Z�R�]��Xa�u�d���g��>k�W|n�ݲq���t��x�~0{��N~�����9>��ƃ��K���φ��Q���щ�"P��͌��H�����;��5����)����������������k���ܜ�$M������,������,
��~x���榼}T��/©��/��[����
��`x���尼jS������.��Ŝ���
��Vy��躼W���ƽ��  �  d�N=/�M=�5M=�|L=��K=
K=6PJ=ܕI=�H=�H=8dG=�F=R�E=.E=3pD=ɱC=��B=�2B=YrA=	�@=��?=�+?=�g>= �==
�<=�<=�M;=N�:=��9=��8= 8=@Q7=π6=ˮ5=�4=�4=F.3=�T2=�y1=�0=A�/=
�.=L�-=�-=�#,=�6+=�F*=0S)=�\(=jb'=�d&=<c%=�]$=�T#=�F"=5!=� =�=��=^�=��=�f=�2=B�=F�=�u=�+=��=�=~*=M�=^b=��=_�
=g	=�=�
=��=(�=�b=Е�<�\�<��<��<�z�<)�<S��<�L�<���<U]�<D��<�R�<7��<�/�<��<.��<�S�<B��<���<�N�<���<i�<�(�<�k�<���<-�<}$�<�]�<Y��<=˗<���<3�<ue�<���<�Ǆ<���<�Qz<��r<�k<�uc<��[<t=T<�L<rE<�w=<��5<QW.<`�&<�E<;�<�E<��<[<��;��;�V�;���;��;+��;�	�;���;>�~;�9b;��E;��);�;���:�ͭ:g�n:��: =�8n���H�:�_B��щĺF;�����$b-�&�E�S�]�k�u�+����	���d��咨������f��vɻ��ӻ��ݻ������i���˟��W�-��O���Jh�+����!��)&�AF*�R.�eM2�496��:��=�i�A��WE�3�H���L��'P��S��%W�n�Z���]�Ya���d�h�g�.?k��|n�L�q�7�t� x��0{�=O~�%���T>��&ƃ��K���φ�vQ���щ�P��͌�vH����f;������~)��ߞ��_��͆��u���Uk��vܜ�M��򼟼t,��p���!
��{x���榼�T��C©��/��|������x��氼�S��;���/������ ���y��5躼KW���ƽ��  �  \�N="�M=�5M=�|L=��K=&
K=?PJ=�I=1�H=�H=IdG=�F=j�E=*.E=SpD=�C=��B=�2B=jrA=#�@=��?=�+?=�g>=�==�<=�<=�M;=C�:=��9=|�8= 8=%Q7=��6=��5=��4=�4=(.3=�T2=�y1=�0=.�/=��.=D�-=�-=�#,=�6+=�F*=:S)=�\(=vb'=�d&=Qc%=�]$=�T#=G"=)5!=� =�=�=n�=��=�f=�2=G�=N�=�u=w+=��=݅=q*=<�=Eb=��=>�
=I	=ɍ=�
=��=�=cb=���<�\�<S�<���<�z�<�<K��<�L�<���<d]�<U��<�R�<h��<�/�<?��<c��<�S�<���<&��<�N�<暹<��<)�<�k�<���<?�<�$�<�]�<O��<>˗<���<3�<Qe�<ږ�<�Ǆ<\��<tQz<>�r<{k<Zuc<g�[<�<T<{�L<%E<ew=<��5<W.<O�&<�E<-�<�E<��<Q[<���;��;0W�;P��;��;��;�
�;z��;"�~;i;b;�E;r�);;!��:|ϭ:۾n:��:D�8|�����:��B����ĺd<�����xc-���E���]�T�u�����
���e��I������g���ɻ�ӻ��ݻ�绷��������YW���������g�ʺ��!�?)&��E*��Q.�M2��86�c:���=�G�A�eWE�'�H�L��'P��S��%W���Z��]�MYa�0�d���g��?k�!}n���q���t�`x�51{�mO~�M���e>��;ƃ��K���φ��Q���щ��O���̌�VH��^�C;��ղ��G)������������D���#k��Sܜ��L��Ǽ��Y,��a���
���x���榼�T��^©� 0������)���x��:氼�S��z���9/��0���W���y��c躼mW���ƽ��  �  M�N=�M=�5M=�|L=��K=+
K=FPJ=��I=9�H= H=]dG=7�F=��E==.E=lpD=�C=��B=3B=�rA=+�@=�?=�+?=�g>=�==	�<=�<=�M;=3�:=|�9=l�8=  8=Q7=��6=��5=��4=j4=.3=�T2=fy1=�0="�/=��.=4�-=�-=�#,=�6+=�F*=;S)=�\(=�b'=�d&=dc%=^$=�T#=!G"=<5!=� =�=)�=��=ӕ=�f=�2=T�=K�=�u=s+=��=҅=]*='�=3b=��=�
=6	=��=�
=o�=��=Qb=M��<}\�<)�<���<�z�<��<7��<�L�<���<_]�<t��<�R�<s��<)0�<o��<���<�S�<���<J��<O�<��<��<<)�<�k�<֫�<T�<�$�<�]�<O��<2˗<���<�2�<.e�<Ö�<�Ǆ<,��<6Qz<Ǳr<k<�tc<#�[<�<T<�L<�E<w=<b�5<�V.<7�&<}E<H�<�E<��<�[<���;,�;�W�;#��;��;���;��;-��;կ~;M=b;��E;?�););��:BЭ:�n:��:	C�8������:�>D��X�ĺ�=��\��#d-���E�\�]���u�܃����]f������\����g��ɻ8�ӻ��ݻ��X������m��W�������p�{g�r����!��(&��E*�GQ.��L2��86�F:���=��A�eWE���H���L��'P�*�S�&W��Z�>�]��Ya���d���g�@k�}n��q� �t��x��1{��O~�m����>��\ƃ��K���φ�|Q���щ��O���̌�=H��O�;������)���������u�������j��,ܜ��L������3,��M���

��ox���榼�T��s©�0������?���x��i氼�S������f/��j���v���y���躼�W��ǽ��  �  D�N=�M=�5M=�|L=��K=*
K=MPJ= �I=J�H= H=tdG=D�F=��E=Z.E=�pD=�C=��B= 3B=�rA=>�@=�?=,?=h>=�==�<=�<=�M;=1�:=r�9=^�8=�8=Q7=��6=��5=��4=T4=�-3=�T2=\y1=ٛ0=�/=��.=-�-=�-=�#,=�6+=�F*=;S)=�\(=�b'=�d&=vc%=%^$=�T#=;G"=U5!=� = =7�=��=�=g=�2=Y�=K�=�u=v+=y�=υ=S*=�=b=n�=�
=	=��=�
=T�=��=/b=1��<J\�<�<���<�z�<��<#��<�L�<���<d]�<y��<S�<���<L0�<���<���<T�<۫�<���<6O�<3��<��<c)�<�k�<㫪<e�<�$�<�]�<S��<$˗<���<�2�<e�<���<�Ǆ<��<�Pz<w�r<�k<�tc<��[<S<T<آL<�E<�v=<6�5<�V.<�&<sE<M�<�E<��<�[<z��;��;�X�;���;e�;���;m�;3��;�~;q>b;P�E;��);d;���:�ѭ:_�n:��:\@�8I�����:�E����ĺc@�����e-�;�E���]��u�h�������f��o���ꔳ��g��Eɻ"�ӻ2�ݻ���k�����O���V�e��V���=g���T�!��(&�E*�Q.�eL2�B86�:�f�=��A�\WE��H���L�(P�*�S�&W�
�Z���]��Ya���d�|�g�i@k��}n�p�q�e�t�	x��1{�
P~������>��dƃ� L���φ�pQ���щ��O���̌�!H��+��:�������(��P������=��������j���ۜ��L������),��=���	
��nx���榼�T��p©�10��ٝ��m���x���氼%T�������/���������z���躼�W��ǽ��  �  9�N=�M=�5M=�|L=��K=6
K=\PJ=�I=V�H=! H=dG=T�F=��E=g.E=�pD=�C=��B=.3B=�rA=H�@=�?=,?=h>=�==�<=�<=�M;=(�:=j�9=Y�8=�8=�P7=}�6=y�5=��4=C4=�-3=�T2=Py1=Λ0=�/=��.="�-=�-=�#,=�6+=�F*=PS)=�\(=�b'=�d&=zc%=3^$=�T#=CG"=b5!= =	=D�=��=�=g=�2=^�=`�=�u=s+=s�=��=F*=�=b=_�=�
=�
	=��=�
=E�=��=b=��<*\�<��<���<lz�<��<��<�L�<���<�]�<���<$S�<���<Z0�<���<���<*T�<���<���<JO�<Q��<�<n)�<l�<�<~�<�$�<�]�<N��<˗<���<�2�<e�<y��<nǄ<���<�Pz<Y�r<ck<ntc<q�[<<T<��L<PE<�v=<�5<�V.<��&<dE<Q�<F<6�<�[<���;	�;Y�;)��;��;)��;��;���;��~;x?b;��E;l�);8;���:~ԭ:E�n:��:�>�8c���b�:��E���ĺ�A��P���f-���E� �]��u�x���i���f������C����g���ɻ}�ӻU�ݻ���a��@���*���V�*��?��� �g�޹��!�P(&��D*��P.�,L2�+86��:�G�=�УA� WE�	�H���L�(P�]�S�E&W��Z���]�Za��d���g�t@k�~n���q�z�t�Mx��1{�?P~������>��wƃ�L���φ�nQ���щ��O���̌�H����:��e����(��7������!��������j���ۜ��L��~���,��%����	��nx���榼�T���©�H0��۝�����
y���氼FT�������/���������'z���躼�W��ǽ��  �  8�N=�M=�5M=�|L=��K=0
K=SPJ=�I=Y�H=- H=�dG=b�F=��E=p.E=�pD=%�C=�B=93B=�rA=N�@=$�?=,?=h>=�==�<=�<=�M;=(�:=f�9=K�8=�8=�P7=y�6=n�5=��4=24=�-3=�T2=@y1=0=��/=��.=!�-=�-=�#,=�6+=�F*=ES)=�\(=�b'=�d&=�c%=6^$=�T#=OG"=p5!= ==U�=��=��=g=�2=^�=R�=�u=n+={�=��=E*=�=b=R�=��
=�
	=r�={
=0�=��=b=��<\�<��<���<kz�<��<%��<�L�<���<s]�<���<2S�<���<t0�<���<���<9T�<��<���<eO�<q��<�<�)�<l�<��<p�<�$�<�]�<W��<'˗<���<�2�<�d�<j��<SǄ<���<kPz<�r<+k<tc<T�[<�;T<s�L<7E<�v=<�5<�V.<�&<wE<E�<�E<�<�[<���;l�;KY�;���;P�;u��;��;���;b�~;E@b;��E;��);�;���:Eӭ:��n:?�:7O�8������:�F����ĺ�B��E���f-�G�E�M�]��u�%���s��pg���������:h���ɻu�ӻ�ݻ���O�񻏤��-���V�$�� ��� ��f������!�(&��D*��P.�L2��76��:� �=�ʣA�3WE��H���L��'P�U�S�C&W�B�Z���]�FZa�-�d���g��@k�^~n��q���t�Wx�02{�`P~������>��tƃ�L���φ�yQ���щ��O���̌� H����:��U����(��'��������������j���ۜ�pL��|���,��5����	��ox���榼�T���©�G0��󝬼���%y���氼PT��³��/��ȝ�����7z���躼�W��9ǽ��  �  7�N= �M=�5M=�|L=��K=:
K=YPJ=�I=V�H=5 H=�dG=]�F=��E=l.E=�pD=�C=�B=03B=�rA=P�@=$�?=,?=h>=�==�<=�<=�M;=�:=d�9=G�8=�8=�P7=u�6=c�5=��4=E4=�-3=�T2=;y1=ț0=��/=��.=�-=�-=�#,=�6+=�F*=FS)=�\(=�b'=�d&=�c%=1^$=�T#=OG"=m5!= ==V�=��=�=g=�2=h�=Q�=�u=k+=q�=��=A*=�=b=X�=�
=�
	=g�=�
=;�=��=b=��<)\�<��<���<[z�<��<��<�L�<���<v]�<���<7S�<���<�0�<���<���</T�<��<���<gO�<j��<�<�)�<l�<��<�<�$�<�]�<D��<˗<q��<�2�<�d�<t��<TǄ<���<YPz<�r<vk<tc<;�[<�;T<l�L<PE<�v=< �5<~V.<��&<WE<T�<&F<)�<\<���;��;IY�;x��;X�;X��;��;Ϩ�;a�~;�?b;#�E;�);�;5��:�ӭ:��n:��:�>�8����S�:�MF���ĺkA��m��g-���E���]���u�\���z���g��씨�f���lh���ɻ��ӻQ�ݻ���񻄤�����V�@��ӆ�� ��f������!�(&��D*��P.�4L2��76��:��=���A�5WE���H�ŘL�(P�~�S�R&W�S�Z���]�,Za�D�d���g��@k�~n���q���t�gx�=2{�7P~������>���ƃ�&L���φ�yQ��cщ��O���̌��G����:��c����(��1��������������j���ۜ�ZL�������+��%����	��fx���榼�T���©�I0��������#y���氼YT��³��/��̝�����?z���躼�W��Fǽ��  �  8�N=�M=�5M=�|L=��K=0
K=SPJ=�I=Y�H=- H=�dG=b�F=��E=p.E=�pD=%�C=�B=93B=�rA=N�@=$�?=,?=h>=�==�<=�<=�M;=(�:=f�9=K�8=�8=�P7=y�6=n�5=��4=24=�-3=�T2=@y1=0=��/=��.=!�-=�-=�#,=�6+=�F*=ES)=�\(=�b'=�d&=�c%=6^$=�T#=OG"=p5!= ==U�=��=��=g=�2=^�=R�=�u=o+={�=��=E*=�=b=S�=�
=�
	=r�=|
=1�=��=b=��<\�<��<���<mz�<��<&��<�L�<���<t]�<���<3S�<���<u0�<���<���<:T�<��<���<eO�<q��<�<�)�<l�<��<o�<�$�<�]�<V��<&˗<���<�2�<�d�<j��<SǄ<���<jPz<�r<+k<tc<T�[<�;T<t�L<8E<�v=<�5<�V.<�&<yE<G�<�E<�<�[<���;o�;MY�;���;Q�;v��;��;���;^�~;@@b;��E;��);�;��:1ӭ:��n:�:�M�8����*�:�&F����ĺ�B��P���f-�R�E�W�]��u�)���w��sg���������=h���ɻx�ӻ�ݻ���P�񻑤��.���V�%�� ��� ��f������!�(&��D*��P.�L2��76��:� �=�ʣA�3WE��H���L��'P�U�S�C&W�B�Z���]�FZa�-�d���g��@k�^~n��q���t�Wx�02{�`P~������>��tƃ�L���φ�yQ���щ��O���̌� H����:��U����(��'��������������j���ۜ�pL��|���,��5����	��ox���榼�T���©�G0��󝬼���%y���氼PT��³��/��ȝ�����7z���躼�W��9ǽ��  �  9�N=�M=�5M=�|L=��K=6
K=\PJ=�I=V�H=! H=dG=T�F=��E=g.E=�pD=�C=��B=.3B=�rA=H�@=�?=,?=h>=�==�<=�<=�M;=(�:=j�9=Y�8=�8=�P7=}�6=y�5=��4=C4=�-3=�T2=Py1=Λ0=�/=��.="�-=�-=�#,=�6+=�F*=PS)=�\(=�b'=�d&=zc%=3^$=�T#=CG"=b5!= =	=D�=��=�=g=�2=^�=`�=�u=t+=s�=��=G*=�=b=`�=�
=�
	=��=�
=F�=��=b=��<,\�<��<���<oz�<��<��<�L�<���<�]�<���<&S�<���<[0�<���<���<*T�<���<���<JO�<Q��< �<m)�<l�<�<|�<�$�<�]�<L��<˗<���<�2�<e�<x��<mǄ<���<�Pz<X�r<ck<otc<r�[<<T<��L<SE<�v=<	�5<�V.<��&<hE<T�<F<:�<�[<���;�;
Y�;,��;��;)��;��;���;��~;o?b;��E;^�);(;ַ�:Xԭ:��n:��:�;�8�����:��E���ĺ�A��f���f-���E�4�]��u�����p���f��ǔ��I����g���ɻ��ӻY�ݻ���d��B���+���V�+��@��� �g�߹��!�P(&��D*��P.�,L2�,86��:�G�=�УA� WE�	�H���L�(P�]�S�E&W��Z���]�Za��d���g�t@k�~n���q�z�t�Mx��1{�?P~������>��wƃ�L���φ�nQ���щ��O���̌�H����:��e����(��7������!��������j���ۜ��L��~���,��%����	��nx���榼�T���©�H0��۝�����
y���氼FT�������/���������'z���躼�W��ǽ��  �  D�N=�M=�5M=�|L=��K=*
K=MPJ= �I=J�H= H=tdG=D�F=��E=Z.E=�pD=�C=��B= 3B=�rA=>�@=�?=,?=h>=�==�<=�<=�M;=1�:=r�9=^�8=�8=Q7=��6=��5=��4=T4=�-3=�T2=\y1=ٛ0=�/=��.=-�-=�-=�#,=�6+=�F*=;S)=�\(=�b'=�d&=vc%=&^$=�T#=;G"=U5!=� = =7�=��=�=g=�2=Y�=K�=�u=w+=y�=υ=T*=�= b=o�=�
=	=��=�
=V�=��=1b=4��<M\�<�<���<�z�<��<'��<�L�<���<g]�<|��<S�<���<N0�<���<���<T�<۫�<���<6O�<2��<��<b)�<�k�<᫪<c�<�$�<�]�<Q��<"˗<���<�2�<e�<���<�Ǆ<	��<�Pz<w�r<�k<�tc<��[<V<T<ۢL<�E<�v=<:�5<�V.<�&<xE<S�<�E<��<�[<���;��;�X�;���;g�;���;l�;0��;��~;d>b;@�E;��);N;˶�:Pѭ:��n:m�:e<�8N����:�VE����ĺ�@������e-�W�E���]��u�t�������f��x���򔳻�g��Lɻ(�ӻ7�ݻ���o�����P���V�g��W���>g���U�!��(&�E*�Q.�eL2�B86�:�f�=��A�\WE��H���L�(P�*�S�&W�
�Z���]��Ya���d�|�g�i@k��}n�p�q�e�t�	x��1{�
P~������>��dƃ� L���φ�pQ���щ��O���̌�!H��+��:�������(��P������=��������j���ۜ��L������),��=���	
��nx���榼�T��p©�10��ٝ��m���x���氼%T�������/���������z���躼�W��ǽ��  �  M�N=�M=�5M=�|L=��K=+
K=FPJ=��I=9�H= H=]dG=7�F=��E==.E=lpD=�C=��B=3B=�rA=+�@=�?=�+?=�g>=�==	�<=�<=�M;=3�:=|�9=l�8=  8=Q7=��6=��5=��4=j4=.3=�T2=fy1=�0="�/=��.=4�-=�-=�#,=�6+=�F*=;S)=�\(=�b'=�d&=dc%=^$=�T#=!G"=<5!=� =�=)�=��=ԕ=�f=�2=U�=K�=�u=t+=��=Ӆ=^*=(�=4b=��=!�
=8	=��=�
=q�=��=Sb=R��<�\�<-�<���<�z�<�<;��<�L�<���<b]�<w��< S�<u��<+0�<q��<���<�S�<���<J��<O�<��<��<:)�<�k�<ԫ�<R�<�$�<�]�<L��</˗<���<�2�<,e�<���<�Ǆ<+��<4Qz<Ʊr<k<�tc<%�[<�<T<�L<�E<w=<h�5<�V.<>�&<�E<N�<�E<��<�[<���;4�;�W�;'��;��;���;��;*��;ɯ~;<=b;��E;'�);;ʵ�:�ϭ:�n:'�:*>�8������:��D����ĺ$>�����Hd-���E�~�]�şu�ꃆ���if�����f����g��!ɻ@�ӻ�ݻ��]������o��W�������q�|g�s����!��(&��E*�GQ.��L2��86�F:���=��A�eWE���H���L��'P�*�S�&W��Z�>�]��Ya���d���g�@k�}n��q� �t��x��1{��O~�m����>��\ƃ��K���φ�|Q���щ��O���̌�=H��O�;������)���������u�������j��,ܜ��L������3,��M���

��ox���榼�T��s©�0������?���x��i氼�S������f/��j���v���y���躼�W��ǽ��  �  \�N="�M=�5M=�|L=��K=&
K=?PJ=�I=1�H=�H=IdG=�F=j�E=*.E=SpD=�C=��B=�2B=jrA=#�@=��?=�+?=�g>=�==�<=�<=�M;=C�:=��9=|�8= 8=%Q7=��6=��5=��4=�4=(.3=�T2=�y1=�0=.�/=��.=D�-=�-=�#,=�6+=�F*=:S)=�\(=vb'=�d&=Qc%=�]$=�T#=G"=)5!=� =�=�=n�=��=�f=�2=H�=O�=�u=x+=��=ޅ=q*==�=Fb=��=?�
=K	=ˍ=�
=��=�=eb=���<�\�<X�<���<�z�<�<P��<�L�<���<h]�<Y��<�R�<k��<�/�<A��<d��<�S�<���<&��<�N�<嚹<��<)�<�k�<���<<�<�$�<�]�<L��<:˗<���<3�<Oe�<ؖ�<�Ǆ<[��<rQz<=�r<{k<[uc<i�[<=T<�L<*E<jw=<��5<W.<U�&<�E<4�<�E<��<W[<���;��;7W�;U��;��;��;�
�;v��;�~;W;b;��E;X�);�;ܲ�:2ϭ:;�n:�:�>�8������:�C���ĺ�<��$���c-���E���]�w�u�����
���e��U������)g���ɻ��ӻ��ݻ%�绽��������[W���������g�˺��!�@)&��E*��Q.�M2��86�d:���=�G�A�eWE�'�H�L��'P��S��%W���Z��]�MYa�0�d���g��?k�!}n���q���t�`x�51{�mO~�M���e>��;ƃ��K���φ��Q���щ��O���̌�VH��^�C;��ղ��G)������������D���#k��Sܜ��L��Ǽ��Y,��a���
���x���榼�T��^©� 0������)���x��:氼�S��z���9/��0���W���y��c躼mW���ƽ��  �  d�N=/�M=�5M=�|L=��K=
K=6PJ=ܕI=�H=�H=8dG=�F=R�E=.E=3pD=ɱC=��B=�2B=YrA=	�@=��?=�+?=�g>= �==
�<=�<=�M;=N�:=��9=��8= 8=@Q7=π6=ˮ5=�4=�4=F.3=�T2=�y1=�0=A�/=
�.=L�-=�-=�#,=�6+=�F*=0S)=�\(=jb'=�d&=<c%=�]$=�T#=�F"=5!=� =�=��=^�=��=�f=�2=B�=F�=�u=�+=��=�=*=N�=_b=��=a�
=i	=�=�
=��=+�=�b=Օ�<�\�<��<��<�z�</�<X��<�L�<���<Z]�<H��<�R�<:��<�/�<��<0��<�S�<B��<���<�N�<���<h�<�(�<�k�<���<*�<z$�<�]�<U��<:˗<���<3�<re�<���<�Ǆ<���<�Qz<��r<�k<�uc<��[<x=T<�L<wE<�w=<��5<WW.<g�&<�E<C�<�E<��<"[<��;��;�V�;���; �;,��;�	�;���;0�~;�9b;��E;t�);�;���:Kͭ:»n:��:7�8�����:��B��-�ĺ�;�����Nb-�N�E�y�]���u�<���
���d��򒨻�����f���ɻ��ӻ��ݻ������n���͟��W�/��P���Kh�,����!��)&�AF*�R.�eM2�496��:��=�i�A��WE�3�H���L��'P��S��%W�n�Z���]�Ya���d�h�g�.?k��|n�L�q�7�t� x��0{�=O~�%���T>��&ƃ��K���φ�vQ���щ�P��͌�vH����f;������~)��ߞ��_��̆��u���Uk��vܜ�M��򼟼t,��p���!
��{x���榼�T��C©��/��|������x��氼�S��;���/������ ���y��5躼KW���ƽ��  �  p�N=8�M=�5M=�|L=��K=
K=)PJ=ՕI=�H=�H= dG=�F=5�E=�-E="pD=��C=��B=�2B=GrA=��@=��?=�+?=�g>=�==�<=�<=�M;=V�:=��9=��8=4 8=QQ7=�6=�5=1�4=�4=].3=U2=�y1=#�0=\�/=�.=W�-=�-=�#,=�6+=�F*=&S)=�\(=ab'=�d&=0c%=�]$=kT#=�F"=�4!=� =�=��=D�=��=�f=�2=<�=?�=�u=+=��=��=�*=a�=~b=��=y�
=�	=�==т=I�=�b=��<]�<��<7��<�z�<M�<a��<�L�<���<J]�<@��<�R�<��<�/�<��<���<JS�<!��<���<iN�<}��<2�<�(�<rk�<~��<�<l$�<�]�<K��<C˗<���<+3�<�e�<0��<Ȅ<���<LRz< �r<Nk<@vc<G�[<�=T<1�L<�E<x=<	�5<�W.<��&<�E<;�<�E<l�<[<k��;m�;�U�;���;	�;*��;	�;���;<�~;�7b;1�E;��);];B��:˭:ĺn:2�:5*�8����.�:��A��χĺ9��ݦ��`-���E��]���u�����@	��\d��s���͒��Rf��8ɻn�ӻ��ݻ6�����ť������W����������h������!�*&��F*�oR.��M2�l96�:�<�=���A��WE�&�H���L��'P���S�%W�5�Z�R�]��Xa�u�d���g��>k�W|n�ݲq���t��x�~0{��N~�����9>��ƃ��K���φ��Q���щ�"P��͌��H�����;��5����)����������������k���ܜ�$M������,������,
��~x���榼}T��/©��/��[����
��`x���尼jS������.��Ŝ���
��Vy��躼W���ƽ��  �  ��N==�M=�5M=�|L=��K=
K=PJ=ŕI=��H=�H=dG=ڧF=&�E=�-E=pD=��C=��B=�2B=.rA=�@=��?=�+?=�g>=��==�<=�<=�M;=a�:=��9=��8=D 8=dQ7=�6=��5=C�4=�4=p.3=&U2=�y1=;�0=d�/='�.=h�-=�-=�#,=�6+=}F*=#S)=q\(=Qb'=�d&=c%=�]$=_T#=�F"=�4!=� =�=��=,�=��=�f=�2=/�==�=�u=�+=��= �=�*=u�=�b=��=��
=�	=%�=5=�=d�=�b=2��<=]�<��<e��<{�<Y�<~��<�L�<���<;]�<&��<�R�<��<�/�<���<���<S�<��<���<EN�<^��<��<�(�<Ok�<\��<��<b$�<�]�<T��<R˗<���<Q3�<�e�<E��<KȄ<���<�Rz<q�r<�k<�vc<��[<C>T<��L<E<8x=<[�5<�W.<��&<�E<4�<�E<8�<�Z<���;��;�T�;���;x�;-��;<�;���;&�~;6b;i�E;�);  ;ˬ�:,ɭ:�n:�:\4�8����^�:��?��r�ĺ7�����_-���E��]�v�u��������c��ő�������e���ɻy�ӻ��ݻ8�������A��X����ֈ����h���M�!�q*&�#G*��R.�>N2��96�W:�~�=�ФA��WE�K�H���L��'P���S�>%W���Z�4�]�lXa��d���g��>k� |n���q��t�6x�30{��N~�賀�>���Ń��K���φ��Q���щ�7P��.͌��H�����;��g����)��U������<��������k���ܜ�AM��;����,������5
���x���榼mT��)©��/��D����
��3x���尼9S�������.�������
��$y���纼W���ƽ��  �  ��N=E�M=�5M=�|L=��K=
K=PJ=��I=��H=�H=�cG=ŧF=�E=�-E=�oD={�C=f�B=�2B=rA=հ@=��?=�+?=�g>=�==�<=�<=�M;=i�:=��9=��8=W 8=|Q7=�6=�5=_�4=�4=�.3=6U2=�y1=M�0=u�/=5�.=n�-=�-=�#,=�6+=vF*="S)=m\(=Gb'=�d&=	c%=�]$=AT#=�F"=�4!=o =s=��=$�=�=�f=�2=,�=>�=�u=�+=��=�=�*=��=�b=��=��
=�	=F�=P=�=��=�b=m��<j]�<�<~��<5{�<a�<���<�L�<���<D]�<��<�R�<���<y/�<���<���<�R�<Ū�<Y��<N�<+��<��<z(�<3k�<G��<��<Y$�<�]�<Z��<M˗<���<W3�<�e�<k��<xȄ<��<�Rz<�r<k<wc<�[<�>T<�L<kE<�x=<o�5<�W.<��&<�E<+�<�E<;�<�Z<s��;0�;�T�;H��;�
�;�;`�;ݢ�;2�~;�4b;9�E;j�);	�;6��:�ȭ:�n:��:,�8���i�:�P?���ĺ�5������^-�\�E�z�]�B�u�;���3��c��?��� ����e���ɻ[�ӻ��ݻ
��I������W��1X���*���^i�f����!��*&�G*�&S.�fN2�	:6��:���=��A��WE�h�H���L��'P���S�"%W�ɔZ���]�'Xa�Ĭd�g�g�>k��{n�%�q��t��x��/{�MN~�ɳ��>���Ń��K���φ�{Q���щ�4P��=͌��H�����;��~���*��|������e�������k���ܜ�qM��U����,������<
���x���榼rT��©��/��$����
��x���尼S������z.��f����
��y���纼�V��cƽ��  �  ��N=V�M=�5M=�|L=��K=
K=PJ=��I=��H=�H=�cG=��F=��E=�-E=�oD=u�C=U�B=�2B=rA=ɰ@=��?=�+?=�g>=�==�<=�<=�M;=s�:=¹9=��8=\ 8=�Q7=�6=�5=m�4=�4=�.3=BU2=�y1=T�0=��/==�.=s�-=-=�#,=�6+=sF*=S)=c\(=Ab'=�d&=�b%=�]$=1T#=�F"=�4!=a =q=��=�=t�=�f=�2=#�=3�=�u=�+=��=!�=�*=��=�b=�=��
=�	=T�=a=�=��=�b=���<{]�<)�<���<M{�<��<���<�L�<���<0]�<	��<�R�<���<e/�<���<���<�R�<���<D��<�M�<	��<��<_(�<*k�<5��<��<D$�<�]�<]��<Z˗< �<c3�<�e�<}��<�Ȅ<1��<0Sz<#�r<Gk<Ewc<9�[<�>T<�L<�E<�x=<��5<X.<��&<�E<�<cE<�<mZ<V��;��;>T�;���;
�;0�;��;���;�~;�3b;t�E;u�);��;���:ǭ:u�n:{�:�&�8>�B�:��>��b�ĺ5��ң�^-���E���]�x�u��������b�������^e��vɻ��ӻ��ݻ��j��g������LX�!��^��?��i�x����!�+&��G*�kS.��N2�;:6��:���=��A�XE�u�H���L��'P�O�S�%W���Z���]�Xa���d�3�g��=k�n{n��q���t��x��/{�8N~������=���Ń��K���φ�Q���щ�KP��S͌��H��Ï��;������+*������ ��y�������k��ݜ��M��]����,������Q
���x���榼dT�������/������
���w��m尼�R������a.��K����
���x���纼�V��Jƽ��  �  ��N=L�M=�5M=�|L=��K=
K=PJ=��I=��H=�H=�cG=��F=��E=�-E=�oD=`�C=P�B=�2B=rA=��@=��?=�+?=�g>=��==�<=�<=�M;=m�:=˹9=��8=j 8=�Q7=.�6=*�5=w�4= 4=�.3=WU2=�y1=b�0=��/=E�.=v�-=-=�#,=�6+=|F*=S)=e\(=;b'=qd&=�b%=�]$=/T#=�F"=�4!=Q =]=��=
�=k�=�f=�2=%�=7�=�u=�+=��=�=�*=��=�b=�=Ń
=�	=`�=u=)�=��=�b=���<�]�<-�<���<J{�<}�<���<�L�<���<2]�<	��<rR�<���<N/�<n��<���<�R�<���<��<�M�<���<��<Q(�<k�</��<��<P$�<�]�<U��<R˗<���<q3�<�e�<���<�Ȅ<I��<�Sz<D�r<�k<hwc<��[<�>T<@�L<�E<�x=<��5<�W.<��&<�E<6�<�E<
�<hZ<���;��;�S�;y��;�	�;�~�;D�;桍;��~;3b;��E;��);��;C��:�ƭ:~�n:��:$�8����N�:��=��w�ĺ�3�����+]-��E��]�r�u����=���b���������� e��aɻ�ӻ��ݻ;��,��D���|��gX�]��������i����&�!�Q+&��G*�pS.��N2�f:6��:���=��A�XE�R�H���L��'P���S�%W���Z���]��Wa�~�d���g��=k�({n���q���t��x��/{��M~������=���Ń��K���φ�|Q���щ�KP��U͌��H��$Ï�<������0*������!������.���l��$ݜ��M��z����,������D
���x���榼lT��
©��/�����y
���w��U尼�R������<.��;���^
���x���纼�V��Dƽ��  �  ��N=�M=f<M=V�L=��K=:K=ZJ=��I=��H=^,H=�qG=T�F=��E=^>E=��D=E�C=`C=�GB=��A=��@=�@=+F?=��>=+�==��<=06<=�o;=��:=��9=M9=�H8=w{7=ܬ6=��5=�
5=K74=�a3=��2=*�1=��0=��/=�/=65.=�O-=�g,=�|+=��*=̝)=K�(=Q�'=��&=W�%=�$=��#=�"=-�!=�{ =�b=�D=�!=o�=��=.�=�`=�"=��=Z�=�E=i�= �=�3=B�=�^=��
=�r	=$�=�o=��=�V=:�=�( =��<���<�|�<�#�<���<�W�<S��<�k�<���<c�<���<:@�<��<f�<�a�<8��<f
�<SX�<~��<	�<I,�<�l�<۩�<��<�<MS�<���<��<��<w�<�H�<2v�<Ӣ�<�΄<i��<�Kz<��r<�j<�Qc<�[<hT<�aL<_�D<N!=<=�5<T�-<W&<��<�8<��<�-<�� <�r�;��;^��;`��;J�;"��;m�;��;yz;z�];�mA;�0%;�'	;3��:sv�:BrY:���9�K�6QҹvdR�fP����кJ�����3�aL�}�d��]|��뉻�z���۠�a��`��������̻,׻�MỲh�hU������S��	�Ť�1-���� �tL�5�#�r�'�ѿ+���/�q�3��7�Yk;�0?���B���F��-J���M�;DQ��T��/X�;�[���^�Hb�]�e�k�h�(l�kJo�2yr���u���x�~�{���~����������1���������N�����Y��`��	���om���Ⓖ�V��ʕ�0<������������������j���؟�(F��2������L���y���zd��kЩ�E<������������밼~W���ó��/��������xu���⺼
P�������  �  ��N=�M=_<M=X�L=��K=<K=ZJ=��I=��H=_,H=�qG=Y�F=��E=f>E=��D=N�C=bC=�GB=��A=��@=�@=!F?=��>=/�==��<=16<=�o;=��:=��9=Q9=�H8=w{7=ڬ6=��5=�
5=974=�a3=��2=.�1=��0=��/=�/=55.=�O-=�g,=�|+=��*=͝)=F�(=M�'=��&=U�%=�$=��#=$�"=.�!=�{ =�b=�D=�!=l�=�=+�=�`=�"=��=a�=�E=i�=��=�3=@�=�^=��
=�r	=$�=�o=��=�V=5�=�( =��<���<�|�<�#�<���<�W�<b��<�k�<���<�b�<���<B@�<��<n�<�a�<K��<d
�<]X�<���<�<U,�<�l�<�<��<�<PS�<���<��<��<y�<�H�<3v�<Ƣ�<�΄<n��<�Kz<��r<��j<�Qc<�[<jT<�aL<=�D<Q!=<2�5<R�-<�V&<��<�8<��<�-<e� <�r�;���;���;���;BJ�;b��;h�;p��;Kyz;��];�mA;�0%;�'	;��:�v�:�sY:)��9	��6\ҹfdR�ZP��:�к������3��`L��d��^|��뉻�z���۠����v������ƍ̻#׻N�wh�RU������S�	����7-����z �[L�.�#�h�'���+���/�Z�3��7�Ck;�0?��B���F��-J���M�JDQ��T��/X�:�[���^�/Hb�Q�e�t�h�#l��Jo�Zyr���u���x�y�{���~�	��⋂����5������񒈼F�����m��Y������om���Ⓖ�V��ʕ�1<��y���������������j���؟�7F��8������E���q����d��kЩ�J<������������밼|W���ó��/��������vu���⺼P�������  �  ��N=�M=Z<M=W�L=��K=>K=$ZJ=��I=��H=h,H=�qG=d�F=��E=x>E=��D=`�C=hC=�GB=��A=��@=�@=%F?=��>=.�==��<=-6<=�o;=��:=��9=J9=�H8=o{7=Ȭ6=��5=�
5=+74=�a3=u�2=#�1=��0=��/=�/=+5.=�O-=�g,=�|+=��*=ԝ)=O�(=U�'=ĵ&=`�%=�$=��#=.�"=>�!=�{ =�b=�D=�!=v�=�=3�=�`=�"=��=`�=�E=e�=�=�3=2�=�^=��
=�r	=�=�o=��=�V=�=�( =��<���<�|�<u#�<���<rW�<\��<�k�<���<�b�<���<V@�<'��<��<�a�<m��<�
�<�X�<���<'�<y,�<�l�<��<��<"�<ZS�<���<��<��<u�<�H�<$v�<���<�΄<R��<wKz<b�r<��j<�Qc<��[<'T<�aL<�D<0!=<��5<E�-<�V&<��<�8<��<�-<t� <;s�;B��;��;���;�J�;��;��;��;�yz;��];�nA;�1%;�(	;��:0x�: tY:��9�{�6�ҹ�dR��Q����кn��]���3��aL�T�d�\_|��뉻G{��"ܠ������������̻)׻:N�fh�_U��j���S��	�n��-����a �1L��#�&�'��+���/��3�ė7�
k;��/?���B�p�F��-J���M�_DQ��T��/X�g�[���^�`Hb�z�e���h�Ll��Jo�}yr�ơu��x���{���~����������;������򒈼I������a��C������Tm���Ⓖ�V���ɕ�<��T����������t����j���؟�0F��&������F���p����d��oЩ�_<��&���������밼�W���ó��/��/�������u���⺼3P������  �  }�N=�M=W<M=V�L=��K=@K=*ZJ=��I=��H=u,H=�qG=y�F=��E=�>E=āD=p�C=�C=�GB=��A=��@=�@=8F?=��>=1�==��<=-6<=~o;=��:=��9=:9=H8=Z{7=��6=��5=�
5=74=�a3=e�2=�1=��0=��/=�/=$5.=�O-=�g,=�|+=��*=՝)=X�(=b�'=ǵ&=o�%=,�$=ԫ#=D�"=S�!=�{ =�b=�D=�!=��=�==�=�`=�"=��=[�=�E=U�=�=�3=�=�^=��
=�r	=��=�o=��=�V=
�=f( =��<���<�|�<^#�<���<kW�<Y��<�k�<���<c�<���<e@�<E��<��<b�<���<�
�<�X�<̢�<V�<�,�<�l�<��<��<4�<`S�<���<��<��<\�<�H�<v�<���<�΄<-��<%Kz<��r<G�j<-Qc<A�[<�T<HaL<˿D<� =<ۄ5<�-<�V&<��<�8<��<�-<ð <qs�;���;���;���;aK�;���;��;���;�{z;@�];pA;�2%;�)	;٭�: y�:�uY:f��9��6�ҹ�eR�,R��T�к���k���3��bL���d�`|��쉻�{���ܠ�G��,������2�̻�׻#NỂh�1U��T��kS��	�^���,�x������K���#�Ԫ'�0�+�E�/�۴3���7��j;��/?���B�k�F��-J���M�ZDQ�C�T��/X�|�[��^��Hb�Дe��h��l�Ko��yr�'�u�[�x���{�/�~�<��������N�������@������A��2������4m��vⒼ�V���ɕ��;��/������V���W����j���؟�
F��������?���v����d���Щ�m<��=���������밼�W���ó��/��`�������u���⺼MP��$����  �  s�N=�M=V<M=S�L=��K=IK=3ZJ=��I=��H=�,H=�qG=��F=��E=�>E=�D=��C=�C=HB=��A=��@=�@=FF?=��>=<�==��<=,6<=zo;=��:=��9=#9=kH8=@{7=��6=h�5=�
5= 74=�a3=N�2=��1=~�0=��/=�/=5.=�O-=�g,=�|+=�*=ݝ)=d�(=t�'=ܵ&=��%=>�$=�#=\�"=m�!=�{ =�b=�D=�!=��='�=L�=�`=�"= �=S�=�E=I�=֔=k3=�=�^=��
=�r	=��=�o=��=iV=��=G( =c�<}��<e|�<<#�<l��<]W�<K��<�k�<���<$c�<���<�@�<r��<��<@b�<���<�
�<�X�<��<��<�,�<�l�<=��<�<I�<tS�<���<��<��<L�<�H�<�u�<h��<`΄<���<�Jz<w�r<��j<�Pc<�[<pT<�`L<o�D<� =<��5<��-<�V&<��<�8<Ѱ<�-< � <�s�;���;S��;|��;\L�;���;��;���;�}z;��];�qA;�4%;+	;P��:�z�:�yY:���9:}�6@ҹEgR��R����к�������3�OdL�F�d��a|��퉻P|��qݠ�������������̻�׻NỐh��T����6S�[	���K,�&�����jK�!�#�Y�'�ƾ+���/���3��7��j;�v/?��B�M�F�h-J���M�^DQ�b�T��/X�ǖ[�g�^��Hb�6�e�]�h�,l��Ko�Hzr���u���x�Y�{��~�k��"������Z��� ��򒈼,���$��������m��IⒼXV���ɕ��;������j��"���/����j���؟��E��������6���}����d���Щ��<��i���H��$���
찼�W��ĳ�90������	���u��㺼vP��Q����  �  ^�N=��M=M<M=Q�L=��K=PK=FZJ=ΠI=��H=�,H=�qG=��F=��E=�>E=�D=��C=�C="HB=؈A=��@=�@=SF?=ƃ>=?�==��<=&6<=uo;=��:=v�9=9=RH8=){7=z�6=I�5=q
5=�64=|a3=(�2=ذ1=h�0=��/=�/=5.=�O-=�g,=�|+= �*=�)=t�(=��'=�&=��%=`�$=�#=z�"=��!=| =�b=�D=�!=��=:�=X�=�`=�"=��=P�=�E=@�=��=Q3=��=�^=i�
=dr	=��=^o=��=DV=��=)( =!�<R��<.|�<#�<Z��<EW�<A��<�k�<���<8c�<��<�@�<���<�<ib�<��<,�<#Y�<<��<��<-�<"m�<p��<�<s�<�S�<���<��<��<:�<qH�<�u�<B��<3΄<���<-Jz<�r<5�j<:Pc<F�[<�T<l`L<�D<E =<M�5<��-<�V&<��<�8<�<K.<5� <�t�;J��;P��;���;HM�;Ĭ�;��;֤�;�z;G�];�sA;16%;�,	;���:�}�:&|Y:���9���6�ҹYiR��T����кA�����3�	fL�ϐd��c|�Am}��9ޠ����@�������̻�׻]N�uh��T������R� 	�����+�������J���#�Щ'�D�+�o�/���3���7�Cj;�6/?�A�B� �F�t-J���M��DQ�o�T�90X��[���^�QIb���e���h��l�Lo��zr�	�u�R�x���{���~����L������`�����򒈼+��΋��
���~������l��Ⓖ.V��Gɕ�i;������1��錛�����hj��T؟��E��޲�����;���~����d���Щ��<������m��O���J찼DX��Kĳ�0��ќ��c	��0v��3㺼�P��q����  �  J�N=��M=@<M=Q�L=�K=SK=OZJ=ܠI=�H=�,H=rG=ӶF= �E=�>E=�D=��C=�C=FHB=�A=��@=@=_F?=σ>=@�==��<= 6<=eo;=��:=a�9=�9=.H8={7=^�6=*�5=K
5=�64=[a3=�2=��1=F�0=��/=�/=�4.=�O-=�g,=�|+=�*=�)=}�(=��'=�&=��%=��$='�#=��"=��!=/| =c=�D=�!=��=Q�=i�=�`=�"=��=V�=�E=,�=��=83=��=q^=H�
==r	=��=,o=U�=V=��=( =��<��<�{�<�"�<.��<*W�<P��<�k�<���<Gc�<4��<�@�<Φ�<Y�<�b�<S��<^�<hY�<���<�<I-�<Km�<���<@�<��<�S�<���<��<��<!�<MH�<�u�<���<�̈́<���<�Iz<��r<~�j<�Oc<��[<iT<�_L<~�D<�=<�5<m�-<^V&<��<�8<��<m.<p� <�u�;���;U��;� �;�N�;��;��;@��;�z;��];�uA;8%;�.	;
��:}�: ~Y:��9���6�ҹfkR��V����к&��O���3��gL��d�f|�#X~���ޠ���������w�̻.׻�N�%h뻳T��i���R��	�3���+�
�����GJ��#�[�'���+���/�k�3�d�7��i;��.?��B���F�d-J�z�M��DQ���T�}0X�a�[��^��Ib��e�{�h�l��Lo�]{r���u���x��{�y�~����w�����������ْ��&����������~��N����l���ᒼ�U���ȕ�6;��p��������������Bj�� ؟��E��˲�����*���w����d���Щ��<�������������{찼�X���ĳ��0������	��bv��n㺼�P�������  �  <�N=��M=><M=F�L=�K=`K=[ZJ=�I= �H=�,H=%rG=�F=@�E=?E=J�D=��C=�C=^HB=�A=�@=)@=rF?=݃>=M�==��<=6<=ao;={�:=Q�9=�9=H8=�z7==�6=�5=*
5=�64=2a3=�2=��1=,�0=|�/=u/=�4.=�O-=�g,=�|+=�*=��)=��(=��'="�&=Զ%=��$=D�#=��"=ѐ!=W| =(c=E="=��=f�=z�= a=�"=��=E�=�E=�=��=3=��=U^=�
=r	=\�=	o=-�=�U=s�=�' =��<���<�{�<�"�<��<W�<7��<�k�<��<ac�<P��<A�<��<��<�b�<���<��<�Y�<ɣ�<D�<�-�<�m�<Ԫ�<m�<��<�S�<���<���<��<�<5H�<hu�<ѡ�<�̈́<5��<Iz<ޟr<�j<Oc<!�[<�T<i_L< �D<v=<��5<B�-<MV&<Q�<�8<&�<�.<ñ <>v�;!��;M��;��;�O�;A��;[!�;f��;o�z;��];LxA;t:%;G0	;+��:��:�Y:���9�x�6�ҹQlR�8X��s�к����V�3��iL���d�fg|�Q���B���ߠ�6�����'�����̻s׻�N�zh�dT�����~R�w	�Ԣ�+�������I�w�#���'�!�+�o�/��3�ҕ7�ti;��.?���B���F�<-J���M��DQ�ҿT��0X���[�p�^�5Jb���e���h��l�%Mo��{r�!�u�H�x���{���~��������������'��撈�����������~�����Zl���ᒼ�U���ȕ��:��&������o���w����i���ן��E���������!��������d���Щ��<��⨬����ɀ���찼�X���ĳ�1��`����	���v���㺼Q��;���  �  /�N=��M=8<M=G�L=�K=iK=hZJ=�I=/�H=�,H=<rG=�F=c�E=)?E=l�D=�C=!C=}HB=*�A=�@=:@=�F?=�>=X�==��<=6<=Yo;=h�:=D�9=�9=H8=�z7=!�6=��5=
5=x64=a3=щ2=y�1=�0=h�/=a/=�4.=�O-=�g,=�|+=�*=��)=��(=��'=0�&=�%=��$=k�#=٠"=�!=u| =Bc=@E=-"=��=r�=��=a=�"=�=@�=�E=�=��=3=��=8^=��
=�q	=5�=�n=�=�U=Q�=�' =a�<���<�{�<�"�<���<W�<*��<�k�<	��<�c�<p��<0A�<4��<��<1c�<���<��<�Y�<��<��<�-�<�m�<���<��<��<�S�<Ǉ�<���<��<��<H�<:u�<���<�̈́<���<�Hz<G�r<��j<mNc<��[<OT<�^L<ͽD<=<w�5<��-<.V&<P�<�8<G�<�.<� <�v�;ٖ�;��;��;�P�;0��;�"�;Q��;�z;�];�yA;�;%;�1	;T��:ă�:&�Y:x��9w�68ҹ�oR�(Y����к�������3�wkL���d�@i|�B�����࠻���M�������̻�׻�N�mh�!T�����<R�!	�����*�=��{��UI���#�2�'���+�Ϳ/���3�q�7�9i;�A.?���B���F�-J���M��DQ��T��0X���[���^��Jb� �e�X�h�5l��Mo�f|r���u���x�/�{��~�������3������!��ꒈ�����������l~������0l��Tᒼ^U���ȕ��:��齃�d��#���I����i���ן�]E������z����������d�� ѩ�=����� ��������X��"ų�E1������
���v���㺼2Q�������  �  !�N=��M=.<M=G�L=	�K=jK=rZJ=�I=F�H=-H=WrG=)�F=y�E=G?E=��D=/�C=7C=�HB=D�A=,�@=P@=�F?=�>=W�==��<=6<=Po;=^�:=4�9=�9=�G8=�z7=�6=��5=�	5=W64=�`3=��2=d�1=��0=Q�/=N/=�4.=�O-=�g,=�|+=�*=�)=��(=ɱ'=G�&= �%=ɳ$=�#=��"=�!=�| =^c=SE=D"=�=��=��=a=�"=��=@�=�E= �=s�=�2=u�=^=��
=�q	=�=�n=��=�U=0�=�' =�<e��<q{�<v"�<���<�V�<)��<�k�<��<�c�<���<ZA�<a��<��<\c�<��<2�<(Z�<=��<��<�-�<�m�<%��<��<��<�S�<͇�<���<��<��<�G�<u�<s��<P̈́<���</Hz<۞r<�j<�Mc<5�[<�T<�^L<P�D<�=<4�5<��-<V&<J�<�8<J�<�.<F� <�w�;���;��;��;�Q�;@��;�#�;z��;Ĉz;�];�{A;�=%;h3	;2��:s��:G�Y:���91K�6>ҹ�pR��Z����к�����B�3��lL�&�d�(k|�򉻿����ᠻ������=���{�̻�׻�N�Kh�T�����
R��	�5��U*�ם�$���H��#���'�8�+�w�/�8�3��7��h;��-?�b�B���F�-J���M��DQ��T�1X�C�[��^��Jb�q�e���h��l�)No��|r��u� �x�}�{���~�A��֌��J������2��㒈�����������C~�������k��ᒼ1U��Bȕ�a:������5����������i���ן�HE������t����������d��ѩ�=��/���8��+���0�7Y��Uų��1��ܝ��X
��w��亼lQ������  �  �N=��M=,<M=D�L=
�K=nK=~ZJ=�I=U�H=-H=jrG=9�F=��E=_?E=��D=F�C=IC=�HB=U�A=:�@=Z@=�F?=��>=W�==��<=6<=No;=V�:=!�9=�9=�G8=�z7=�6=��5=�	5=D64=�`3=��2=T�1=��0=H�/=E/=�4.=�O-=�g,=�|+=�*=�)=��(=α'=V�&=�%=߳$=��#=�"=�!=�| =uc=bE=Y"=�=��=��=a=�"=��=>�=�E=��=d�=�2=k�=^=��
=�q	=��=�n=��=�U=�=�' =��<U��<J{�<]"�<���<�V�<-��<�k�<)��<�c�<���<sA�<���<�<|c�<0��<M�<WZ�<k��<��<.�<n�<G��<��<��<�S�<·�<���<��<��<�G�<	u�<[��<1̈́<���<�Gz<��r<��j<�Mc<Ȧ[<�T<M^L<�D<�=<�5<��-<�U&<;�<�8<Z�<+/<i� <x�;���;���;7�;_R�;��;$�;L��;�z;W�];&}A;�>%;@4	;���:���:�Y:���9�L�6�ҹGrR��\����кH������3�GnL�=�d�:l|�u򉻃����ᠻ��5��z����̻׻O�Sh�T��,���Q��	���*�z�����~H�0�#�t�'�ӻ+�4�/�ݱ3��7��h;��-?�I�B�d�F�-J���M��DQ�#�T�G1X�m�[�8�^�?Kb���e�8�h��l�wNo�#}r�b�u���x���{���~�H������\������;��ْ�����g������5~�������k������U��ȕ�F:��������Ջ�������i���ן�6E��l���f����������d��ѩ�E=��?���O��I���W�kY��tų��1�������
��?w��,亼�Q��'����  �  	�N=��M=+<M=D�L=�K=tK=�ZJ=$�I=\�H= -H=rrG=J�F=��E=h?E=��D=O�C=_C=�HB=^�A=E�@=b@=�F?=��>=\�==��<=6<=Io;=M�:=�9=�9=�G8=�z7=�6=��5=�	5=464=�`3=��2=D�1=��0=<�/=:/=�4.=�O-=�g,=�|+=�*=�)=��(=۱'=`�&=�%=�$=��#=�"=&�!=�| =c=vE=b"=%�=��=��= a=�"= �=;�=�E=��=Z�=�2=[�=�]=��
=�q	=��=�n=��=�U=
�=t' =��<5��<9{�<G"�<���<�V�<'��<�k�<*��<�c�<���<�A�<���<)�<�c�<D��<j�<iZ�<���<�<!.�<(n�<T��<��<��<�S�<Շ�<���<��<��<�G�<�t�<G��<̈́<���<�Gz<K�r<k�j<lMc<��[<[T<^L<�D<n=<ς5<��-<�U&<:�<�8<q�<5/<�� <<x�;e��;���;��;S�;i��;�$�;���;��z;I�];�}A;?%;�4	;"��:!��:�Y:1��9.��6�ҹtR��\��m�к������3��nL�L�d�m|��򉻭���m⠻n����������̻E׻�N�Ih��S�����Q��	�ȡ��)�S�����OH�	�#�E�'���+��/���3���7�mh;��-?�&�B�\�F��,J���M��DQ�E�T�f1X���[�m�^�mKb��e�P�h�l��No�j}r���u���x���{���~�d�����n������7��ܒ�����d���r�� ~�������k�������T���Ǖ�):��q��������������oi��}ן�E��g���]����������d��%ѩ�N=��Z���b��g���p�vY���ų��1��!����
��Uw��L亼�Q��E����  �  �N=��M=(<M=>�L=
�K=yK=�ZJ=&�I=Z�H=(-H=srG=J�F=��E=m?E=��D=R�C=^C=�HB=c�A=K�@=b@=�F?=��>=c�==��<=6<=Ho;=P�:=$�9=�9=�G8=�z7=�6=��5=�	5=564=�`3=��2=?�1=��0=7�/=8/=�4.=�O-=�g,=�|+=�*=�)=��(=۱'=^�&= �%=�$=��#=�"=1�!=�| =~c=xE=^"=*�=��=��="a=�"=�=2�=�E=��=a�=�2=V�=�]=��
=�q	=��=�n=��={U=�=n' =��<$��<B{�<M"�<���<�V�<��<�k�<&��<�c�<���<�A�<���<$�<�c�<F��<��<uZ�<���<�<".�<9n�<N��<��<��<�S�<҇�<칛<��<��<�G�<�t�<A��<
̈́<v��<�Gz<%�r<p�j<IMc<��[<DT<�]L<�D<R=<��5<��-<�U&<$�<�8<��<5/<�� <1x�;���;���;��;S�;���;>%�;���;��z;$�];+~A;�?%;�4	;r��:��:��Y:���9�O�6�ҹ>sR�\����к�����S�3�oL���d�m|�:󉻼����⠻e���������̻̐K׻Oốh��S�����Q��	�Ρ��)�Z�����OH�܀#��'���+�ؾ/���3���7�mh;��-?��B�Z�F��,J���M��DQ�L�T�F1X���[���^�eKb��e�X�h�Bl��No�p}r���u���x��{���~�s������f����;��蒈����f���q��~�������k�������T���Ǖ�:��e��������������]i���ן�E��g���V����������d��%ѩ�9=��f���h��n���{�|Y���ų��1��1����
��`w��V亼�Q��R����  �  	�N=��M=+<M=D�L=�K=tK=�ZJ=$�I=\�H= -H=rrG=J�F=��E=h?E=��D=O�C=_C=�HB=^�A=E�@=b@=�F?=��>=\�==��<=6<=Io;=M�:=�9=�9=�G8=�z7=�6=��5=�	5=464=�`3=��2=D�1=��0=<�/=:/=�4.=�O-=�g,=�|+=�*=�)=��(=۱'=`�&=�%=�$=��#=�"=&�!=�| =c=vE=b"=%�=��=��= a=�"= �=<�=�E=��=Z�=�2=[�=�]=��
=�q	=��=�n=��=�U=�=u' =��<6��<;{�<I"�<���<�V�<(��<�k�<+��<�c�<���<�A�<���<*�<�c�<D��<j�<iZ�<���<�<!.�<'n�<S��<��<��<�S�<ԇ�<���<��<��<�G�<�t�<F��<̈́<���<�Gz<K�r<k�j<lMc<��[<\T<	^L<�D<p=<҂5<��-<�U&<=�<�8<s�<8/<�� <@x�;h��;���;��;S�;i��;�$�;���;��z;B�];�}A;u?%;�4	;
��:��:��Y:���9o��6zҹGtR�]����к������3��nL�Y�d�%m|��򉻲���r⠻r����������̻H׻�N�Lh��S�����Q��	�ɡ��)�S�����OH�	�#�F�'���+��/���3���7�mh;��-?�'�B�\�F��,J���M��DQ�E�T�f1X���[�m�^�mKb��e�P�h�l��No�j}r���u���x���{���~�d�����n������7��ܒ�����d���r�� ~�������k�������T���Ǖ�):��q��������������oi��}ן�E��g���]����������d��%ѩ�N=��Z���b��g���p�vY���ų��1��!����
��Uw��L亼�Q��E����  �  �N=��M=,<M=D�L=
�K=nK=~ZJ=�I=U�H=-H=jrG=9�F=��E=_?E=��D=F�C=IC=�HB=U�A=:�@=Z@=�F?=��>=W�==��<=6<=No;=V�:=!�9=�9=�G8=�z7=�6=��5=�	5=D64=�`3=��2=T�1=��0=H�/=E/=�4.=�O-=�g,=�|+=�*=�)=��(=α'=V�&=�%=߳$=��#=�"=�!=�| =uc=bE=Y"=�=��=��=a=�"=��=>�=�E=��=d�=�2=k�=^=��
=�q	= �=�n=��=�U=�=�' =��<Y��<M{�<a"�<���<�V�<0��<�k�<,��<�c�<���<uA�<���<�<}c�<1��<M�<WZ�<k��<��<.�<n�<E��<��<��<�S�<̇�<���<��<��<�G�<u�<Y��</̈́<���<�Gz<��r<��j<�Mc<ʦ[<�T<P^L<�D<�=<�5<��-<�U&<@�<�8<^�<0/<m� <
x�;���;���;;�;aR�;��;$�;J��;�z;K�];}A;�>%;+4	;g��:j��:��Y:���9t�6�ҹ�rR��\��,�кf������3�anL�V�d�Ql|��򉻍��� ⠻��<�������̻	׻	O�Wh�T��/���Q��	���� *�z�����H�0�#�u�'�Ի+�4�/�ݱ3��7��h;��-?�I�B�d�F�-J���M��DQ�#�T�G1X�m�[�8�^�?Kb���e�8�h��l�wNo�#}r�b�u���x���{���~�H������\������;��ْ�����g������5~�������k������U��ȕ�F:��������Ջ�������i���ן�6E��l���f����������d��ѩ�E=��?���O��I���W�kY��tų��1�������
��?w��,亼�Q��'����  �  !�N=��M=.<M=G�L=	�K=jK=rZJ=�I=F�H=-H=WrG=)�F=y�E=G?E=��D=/�C=7C=�HB=D�A=,�@=P@=�F?=�>=W�==��<=6<=Po;=^�:=4�9=�9=�G8=�z7=�6=��5=�	5=W64=�`3=��2=d�1=��0=Q�/=N/=�4.=�O-=�g,=�|+=�*=�)=��(=ɱ'=G�&=�%=ɳ$=�#=��"=�!=�| =^c=SE=D"=�=��=��=a=�"= �=@�=�E= �=t�=�2=v�=^=��
=�q	=�=�n=��=�U=2�=�' = �<i��<v{�<{"�<���<�V�<-��<�k�<��<�c�<���<]A�<c��<��<^c�<��<2�<(Z�<<��<��<�-�<�m�<#��<��<��<�S�<ʇ�<���<��<��<�G�<u�<q��<N̈́<���<,Hz<ڞr<�j<�Mc<7�[<�T<�^L<U�D<�=<:�5<��-<	V&<Q�<�8<Q�</<L� <�w�;���;��;��;�Q�;@��;�#�;v��;��z;��];�{A;�=%;J3	;��:+��:��Y:[��9���6�ҹ�qR��Z���к����i�3�mL�I�d�Ik|��̀���ᠻ�����G�����̻׻�N�Qh�T�����R��	�6��V*�؝�$���H��#���'�8�+�w�/�9�3��7��h;��-?�b�B���F�-J���M��DQ��T�1X�C�[��^��Jb�q�e���h��l�)No��|r��u� �x�}�{���~�A��֌��J������2��㒈�����������C~�������k��ᒼ1U��Bȕ�a:������5����������i���ן�HE������t����������d��ѩ�=��/���8��+���0�7Y��Uų��1��ܝ��X
��w��亼lQ������  �  /�N=��M=8<M=G�L=�K=iK=hZJ=�I=/�H=�,H=<rG=�F=c�E=)?E=l�D=�C=!C=}HB=*�A=�@=:@=�F?=�>=X�==��<=6<=Yo;=h�:=D�9=�9=H8=�z7=!�6=��5=
5=x64=a3=щ2=y�1=�0=h�/=a/=�4.=�O-=�g,=�|+=�*=��)=��(=��'=0�&=�%=��$=k�#=ڠ"=�!=u| =Bc=@E=-"=��=r�=��=a=�"=�=A�=�E=�=��=3=��=:^=��
=�q	=7�=�n=�=�U=T�=�' =g�<���<�{�<�"�<���<W�<0��<�k�<��<�c�<u��<4A�<7��<��<3c�<¹�<��<�Y�<��<��<�-�<�m�<�<��<��<�S�<Ç�<���<��<��<H�<6u�<���<̈́<���<�Hz<F�r<��j<oNc<��[<RT<�^L<ӽD<=<�5<��-<7V&<X�<�8<O�<�.<%� <�v�;��;"��;��;�P�;1��;�"�;L��;�z;��];�yA;�;%;�1	;��:l��:k�Y:���9��6�ҹ�pR��Y��c�к-��� �3��kL��d�hi|�U�����࠻���Z������"�̻�׻�N�th�'T�����>R�#	�����*�>��|��UI���#�2�'���+�Ϳ/���3�q�7�:i;�A.?���B���F�-J���M��DQ��T��0X���[���^��Jb� �e�X�h�5l��Mo�f|r���u���x�/�{��~�������3������!��ꒈ�����������l~������0l��Tᒼ^U���ȕ��:��齃�d��#���I����i���ן�]E������z����������d�� ѩ�=����� ��������X��"ų�E1������
���v���㺼2Q�������  �  <�N=��M=><M=F�L=�K=`K=[ZJ=�I= �H=�,H=%rG=�F=@�E=?E=J�D=��C=�C=^HB=�A=�@=)@=rF?=݃>=M�==��<=6<=ao;={�:=Q�9=�9=H8=�z7==�6=�5=*
5=�64=2a3=�2=��1=,�0=|�/=u/=�4.=�O-=�g,=�|+=�*=��)=��(=��'="�&=Զ%=��$=D�#=��"=ѐ!=W| =(c=E="=��=g�=z�=a=�"=��=F�=�E=�=��=3=��=V^= �
=r	=^�=o=0�=�U=v�=�' =��<���<�{�<�"�<��<W�<=��<�k�<��<gc�<T��<A�<��<��<�b�<���<��<�Y�<ȣ�<B�<-�<�m�<Ъ�<i�<��<�S�<���<���<��<�<1H�<du�<Ρ�<�̈́<2��<Iz<ݟr<�j<
Oc<$�[<�T<o_L<'�D<~=<��5<K�-<VV&<[�<�8</�<�.<˱ <Lv�;-��;W��;��;�O�;B��;X!�;a��;^�z;��];.xA;P:%;0	;ѷ�:���:�Y:?��9��6�ҹ=mR��X����к6��U���3�jL��d��g|�g���U���ߠ�F�����4���ʏ̻}׻�NỂh�kT������R�z	�֢�+���� ���I�x�#���'�"�+�p�/��3�ӕ7�ti;��.?���B���F�=-J���M��DQ�ҿT��0X���[�p�^�5Jb���e���h��l�%Mo��{r�!�u�H�x���{���~��������������'��撈�����������~�����Zl���ᒼ�U���ȕ��:��&������o���w����i���ן��E���������!��������d���Щ��<��⨬����ɀ���찼�X���ĳ�1��`����	���v���㺼Q��;���  �  J�N=��M=@<M=Q�L=�K=SK=OZJ=ܠI=�H=�,H=rG=ӶF= �E=�>E=�D=��C=�C=FHB=�A=��@=@=_F?=σ>=@�==��<= 6<=eo;=��:=a�9=�9=.H8={7=^�6=*�5=K
5=�64=[a3=�2=��1=F�0=��/=�/=�4.=�O-=�g,=�|+=�*=�)=}�(=��'=�&=��%=��$='�#=��"=��!=0| =c=�D=�!=��=Q�=j�=�`=�"=��=V�=�E=-�=��=93=��=s^=J�
=?r	=��=.o=W�=!V=��=
( =��<��<�{�<�"�<5��<0W�<V��<�k�<���<Lc�<9��<�@�<Ҧ�<[�<�b�<T��<_�<hY�<���<
�<F-�<Hm�<���<<�<��<�S�<���<	��<��<�<HH�<�u�<���<�̈́<~��<�Iz<��r<~�j<�Oc<��[<mT<�_L<��D<�=<��5<v�-<hV&<��<�8<��<v.<x� <�u�;��;_��;� �;�N�;��;��;;��;�z;��];�uA;�7%;�.	;���:�:G}Y:J��9��6yҹZlR�MW��E�кa������3��gL��d�4f|�9l~���ޠ������������̻9׻�N�.h뻺T��o���R��	�5���+������HJ��#�\�'���+���/�k�3�d�7��i;��.?��B���F�d-J�z�M��DQ���T�}0X�a�[��^��Ib��e�{�h�l��Lo�]{r���u���x��{�y�~����w�����������ْ��&����������~��N����l���ᒼ�U���ȕ�6;��p��������������Bj�� ؟��E��˲�����*���w����d���Щ��<�������������{찼�X���ĳ��0������	��bv��n㺼�P�������  �  ^�N=��M=M<M=Q�L=��K=PK=FZJ=ΠI=��H=�,H=�qG=��F=��E=�>E=�D=��C=�C="HB=؈A=��@=�@=SF?=ƃ>=?�==��<=&6<=uo;=��:=v�9=9=RH8=){7=z�6=I�5=q
5=�64=|a3=(�2=ذ1=h�0=��/=�/=5.=�O-=�g,=�|+= �*=�)=t�(=��'=�&=��%=`�$=�#=z�"=��!=| =�b=�D=�!=��=:�=Y�=�`=�"=��=Q�=�E=A�==R3=��=�^=k�
=fr	=��=`o=��=GV=��=,( ='�<Y��<5|�<#�<a��<LW�<H��<�k�<���<>c�<��<�@�<���<�<kb�<��<,�<#Y�<;��<��<-�<m�<l��<�<n�<�S�<���< ��<��<5�<mH�<�u�<>��<0΄<���<*Jz<�r<5�j<;Pc<I�[<�T<r`L<�D<L =<U�5<��-<�V&<��<�8<��<T.<=� <�t�;V��;Z��;���;LM�;Ŭ�;��;Ѥ�;�z;0�];�sA;6%;�,	;[��:*}�:U{Y:���9K&�6�ҹEjR�]U��f�кz��+�E�3�<fL���d��c|�V�}��Kޠ����O�����
�̻�׻fN�}h��T������R�"	�����+�������J���#�Щ'�D�+�p�/���3���7�Cj;�6/?�A�B�!�F�t-J���M��DQ�o�T�90X��[���^�QIb���e���h��l�Lo��zr�	�u�R�x���{���~����L������`�����򒈼+��΋��
���~������l��Ⓖ.V��Gɕ�i;������1��錛�����hj��T؟��E��޲�����;���~����d���Щ��<������m��O���J찼DX��Kĳ�0��ќ��c	��0v��3㺼�P��q����  �  s�N=�M=V<M=S�L=��K=IK=3ZJ=��I=��H=�,H=�qG=��F=��E=�>E=�D=��C=�C=HB=��A=��@=�@=FF?=��>=<�==��<=,6<=zo;=��:=��9=#9=kH8=@{7=��6=h�5=�
5= 74=�a3=N�2=��1=~�0=��/=�/=5.=�O-=�g,=�|+=�*=ݝ)=d�(=t�'=ܵ&=��%=>�$=�#=]�"=m�!=�{ =�b=�D=�!=��='�=L�=�`=�"= �=T�=�E=J�=ؔ=l3=�=�^=��
=�r	=��=�o=��=kV=��=J( =h�<���<k|�<B#�<r��<bW�<Q��<�k�<���<)c�<���<�@�<u��<��<Bb�<���<�
�<�X�<��<��<�,�<�l�<:��<��<F�<pS�<���< ��<��<H�<�H�<�u�<e��<]΄<���<�Jz<v�r<��j<�Pc<�[<tT<�`L<u�D<� =<��5<��-<�V&<��<�8<ٰ<.<� < t�;���;[��;���;`L�;���;��;���;�}z;��];�qA;�4%;�*	;���:-z�:1yY:
��9��6�ҹhR�PS���к,����3�}dL�q�d��a|��퉻a|���ݠ�������������̻�׻Nỗh��T����9S�]	���M,�'�����kK�"�#�Z�'�ƾ+���/���3��7��j;�v/?��B�M�F�h-J���M�^DQ�b�T��/X�ǖ[�g�^��Hb�6�e�]�h�,l��Ko�Hzr���u���x�Y�{��~�k��"������Z��� ��򒈼,���$��������m��IⒼXV���ɕ��;������j��"���/����j���؟��E��������6���}����d���Щ��<��i���H��$���
찼�W��ĳ�90������	���u��㺼vP��Q����  �  }�N=�M=W<M=V�L=��K=@K=*ZJ=��I=��H=u,H=�qG=y�F=��E=�>E=āD=p�C=�C=�GB=��A=��@=�@=8F?=��>=1�==��<=-6<=~o;=��:=��9=:9=H8=Z{7=��6=��5=�
5=74=�a3=e�2=�1=��0=��/=�/=$5.=�O-=�g,=�|+=��*=՝)=X�(=b�'=ǵ&=o�%=,�$=ԫ#=D�"=S�!=�{ =�b=�D=�!=��=�==�=�`=�"=��=\�=�E=V�=�=�3=�=�^=��
=�r	=��=�o=��=�V=�=i( =��<���<�|�<c#�<���<pW�<^��<�k�<���<c�<���<h@�<G��<��<b�<���<�
�<�X�<ˢ�<U�<�,�<�l�<��<��<1�<]S�<���<��<��<Y�<�H�<v�<���<�΄<,��<#Kz<��r<G�j<.Qc<C�[<�T<LaL<пD<� =<�5<�-<�V&<��<�8<��<�-<ɰ <{s�;���;���;���;dK�;���;��;���;�{z;/�];�oA;�2%;�)	;���:�x�:auY:$��9
��6Gҹ�fR��R����к(������3�#cL���d�5`|��쉻�{���ܠ�S��7�� ���:�̻�׻*NỈh�6U��X��mS��	�_���,�y������K���#�Ԫ'�0�+�F�/�۴3���7��j;��/?���B�k�F��-J���M�ZDQ�C�T��/X�|�[��^��Hb�Дe��h��l�Ko��yr�'�u�[�x���{�/�~�<��������N�������@������A��2������4m��vⒼ�V���ɕ��;��/������V���W����j���؟�
F��������?���v����d���Щ�m<��=���������밼�W���ó��/��`�������u���⺼MP��$����  �  ��N=�M=Z<M=W�L=��K=>K=$ZJ=��I=��H=h,H=�qG=d�F=��E=x>E=��D=`�C=hC=�GB=��A=��@=�@=%F?=��>=.�==��<=-6<=�o;=��:=��9=J9=�H8=o{7=Ǭ6=��5=�
5=+74=�a3=u�2=#�1=��0=��/=�/=+5.=�O-=�g,=�|+=��*=ԝ)=O�(=U�'=ĵ&=`�%=�$=��#=.�"=>�!=�{ =�b=�D=�!=v�=�=4�=�`=�"=��=`�=�E=e�=�=�3=3�=�^=��
=�r	=�=�o=��=�V=!�=�( =��<���<�|�<x#�<���<uW�<_��<�k�<���<�b�<���<X@�<)��<��<�a�<n��<�
�<�X�<���<&�<w,�<�l�<	��<��< �<WS�<���<
��<��<s�<�H�<#v�<���<�΄<Q��<uKz<a�r<��j<�Qc<��[<)T<�aL<	�D<4!=<�5<I�-<�V&<��<�8<��<�-<x� <Cs�;H��;��;���;�J�;��;��;��;�yz;��];�nA;�1%;�(	;֪�:�w�:�sY:��9�@�6�ҹ
eR��Q����к���z��3��aL�m�d�s_|�
쉻Q{��+ܠ������������̻.׻?N�kh�cU��m���S��	�o��	-����b �2L��#�&�'��+���/��3�ŗ7�
k;��/?���B�q�F��-J���M�_DQ��T��/X�g�[���^�`Hb�z�e���h�Ll��Jo�}yr�ơu��x���{���~����������;������򒈼I������a��C������Tm���Ⓖ�V���ɕ�<��T����������t����j���؟�0F��&������F���p����d��oЩ�_<��&���������밼�W���ó��/��/�������u���⺼3P������  �  ��N=�M=_<M=X�L=��K=<K=ZJ=��I=��H=_,H=�qG=Y�F=��E=f>E=��D=N�C=bC=�GB=��A=��@=�@=!F?=��>=/�==��<=16<=�o;=��:=��9=Q9=�H8=w{7=ڬ6=��5=�
5=974=�a3=��2=.�1=��0=��/=�/=55.=�O-=�g,=�|+=��*=͝)=F�(=M�'=��&=U�%=�$=��#=$�"=.�!=�{ =�b=�D=�!=l�=�=+�=�`=�"=��=a�=�E=i�=��=�3=@�=�^=��
=�r	=%�=�o=��=�V=6�=�( =��<���<�|�<�#�<���<�W�<d��<�k�<���<�b�<���<C@�<��<o�<�a�<L��<e
�<]X�<���<�<T,�<�l�<쩮<��<�<OS�<���<	��<��<w�<�H�<2v�<Ţ�<�΄<m��<�Kz<��r<��j<�Qc<�[<kT<�aL<?�D<S!=<5�5<T�-<�V&<��<�8<��<�-<h� <�r�;���;���;���;CJ�;b��;g�;o��;Fyz;��];�mA;�0%;�'	;���:�v�:[sY:���9lw�6�ҹ�dR�zP��Z�к�����3��`L��d��^|��뉻�z���۠����z������ɍ̻%׻N�yh�TU������S�	����8-����z �[L�.�#�i�'���+���/�Z�3��7�Dk;�0?��B���F��-J���M�JDQ��T��/X�:�[���^�/Hb�Q�e�t�h�#l��Jo�Zyr���u���x�y�{���~�	��⋂����5������񒈼F�����m��Y������om���Ⓖ�V��ʕ�1<��y���������������j���؟�7F��8������E���q����d��kЩ�J<������������밼|W���ó��/��������vu���⺼P�������  �  ��N=�M=2CM=�L=��K=�K=ddJ=ΫI=��H=f9H=�G=O�F=�
F=nOE=ƓD=��C=�C=�]B=��A=��@=y!@=Ha?=1�>=B�==H==HW<=<�;=�:=�:=�;9=r8=��7=��6=�6=�;5=)j4=��3=��2=[�1=
1=�50=�W/=Fw.=S�-=��,=��+=\�*=��)=L�(=�(=E
'=5&=&%=�$=��"=��!=A� =�=�=��=4b=@6=�=��=��=�M=�=p�=.`=�=
�=>;=@�=4Y=�	=_=Q�=�M=��=-&=d� =���<I��< 2�<���<Zl�<���<Є�<[�<n~�<���<V\�<���<�!�<�{�<��<�!�<�m�<ɵ�<��<�:�<~x�<��<��<( �<S�<�<в�<�ߛ<��<�5�<�^�<���<b��<7Մ<���<�Cz<;�r<U�j<�*c<�y[<��S<L<+pD<��<<C 5<�|-<�%<A<z�<�<y�<B  <���;��;��;�A�;�x�;��;`�;���;W v;VY;E�<;�Q ;�;�=�:Q��:�EC:�5�9�Q�����k�����ݺ]y���!�O�:�yNS�(�k�|���ς�����․�h���������Ż�<л��ڻ�����>����V���9�
��b�����Q�c���� �@%��<)�XH-�TB1�Y+5�C9���<���@��5D�R�G�XhK���N��kR���U��CY��\��_��@c�ۃf�S�i���l�^ p��Fs�Lgv���y���|�����X��$܂�c]���܅�IZ��)ֈ�uP��uɋ��@��G���\,��:�����Ԅ������e��}Ԙ��B��!������%�������6`��9ˢ��5��]����
���t��(ߩ�FI��e������������6\���Ƴ�1��盶�����q��fݺ�=I��x����  �  ��N=�M=4CM=�L=}�K=�K=edJ=̫I=��H=f9H=�G=W�F=�
F={OE=ғD=��C=�C=�]B=��A=��@=!@=Ea?=0�>=3�==F==MW<=<�;=�:=�:=�;9=r8=��7=��6=�6=�;5=j4=��3=��2=R�1=1=50=�W/=Kw.=U�-=��,=�+=O�*=v�)=G�(=�(=R
'=6&=,%=$=��"=��!=R� =�=�=��=4b=K6=�=��=��=�M=�=s�=,`=�=�=7;=8�=*Y=�	=_=<�=�M=��=&=[� =���<@��<2�<���<Tl�<���<Є�<=�<g~�<���<[\�<���<�!�<�{�< ��<�!�<�m�<��<*��<�:�<�x�<��<��<' �<S�<݃�<���<�ߛ<��<�5�<�^�<��<Z��<'Մ<���<�Cz<(�r<�j<�*c<�y[<��S<�L<pD<��<<D 5<�|-<�%<+A<\�<O<x�<;  <!��;��;��;7B�;�x�;���;��;��;� v;�VY;x�<;[R ;R;�=�:b��:qBC:�5�9�D��2�'k�c���ݺ�y�N�!��:��NS�k����҂�����"�����������K�Ż�<л��ڻn�什ﻥ����V���>�
�[b�����Q�?��h� ��%��<)�=H-�7B1�9+5�@9���<���@��5D�m�G��hK���N��kR���U��CY��\�/�_��@c���f���i���l�� p�$Gs�Xgv�ցy���|�����X��܂�W]���܅�AZ��&ֈ��P��yɋ�A��?���L,��7������Ȅ������be��^Ԙ��B��������%�������9`��:ˢ��5��o����
���t��ߩ�BI��_������������H\���Ƴ�C1��󛶼���r��tݺ�FI��u����  �  ��N=�M=*CM=�L=��K=�K={dJ=ӫI=��H=p9H=�G=g�F=�
F=�OE=ܓD=��C=�C=�]B=��A=��@=�!@=Ma?=E�>=<�==H==IW<=2�;= �:=�:=�;9=�q8=��7=��6=�6=�;5=j4=��3=r�2=C�1=�1=p50=�W/=<w.=I�-=��,=��+=S�*=��)=X�(=�(=_
'=?&=;%=$=��"=��!=]� =$�=�=ǈ=<b=X6=�=��=��=�M=�=h�=`=�=��=#;=+�=Y=��	=_=*�=�M=��=
&=I� =���<��<�1�<��<:l�<���<ʄ�<E�<�~�<���<j\�<���<�!�<	|�<>��<�!�<�m�<��<D��<;�<�x�<)��<�<5 �<=S�<���<ʲ�<�ߛ<v�<�5�<�^�<ꆌ<<��<Մ<o��<\Cz<��r<��j<�*c<Hy[<�S<�L<�oD<��<< 5<�|-<��%<A<g�<<Έ<U  <���;&�;B�;�B�;uy�;¦;)�;���;�!v;�WY;x�<;ES ;5;0?�:���:�EC:n8�9�F����k����ݺ^z���!�߳:�\OS�S�k�m������Q������丯������Ż=л�ڻ��仂�u����V���"�
�"b�����Q����6� ��%��<)�H-��A1��*5�9���<���@�|5D��G�|hK���N��kR���U��CY�'�\�o�_��@c�1�f�ʿi���l�� p�SGs��gv��y��|�ɦ��X��7܂�n]���܅�MZ��&ֈ��P��Pɋ��@��,���3,��!����������n���Pe��CԘ��B��𯛼����������-`��ˢ��5��g����
��	u��.ߩ�_I��w������͇���h\���Ƴ�]1��������)r���ݺ�bI�������  �  ��N=�M=.CM=��L=��K=�K=wdJ=�I=��H=�9H=�G=��F=�
F=�OE= �D=��C=C=�]B=��A=
�@=�!@=^a?=@�>=F�==H==GW<=6�;=��:=�:=�;9=�q8=�7=��6=c6={;5=�i4=��3=_�2=$�1=�1=_50=�W/=2w.=J�-=��,=��+=^�*=��)=\�(=�(=m
'=\&=P%=1$=��"=��!=z� =H�=!�=ڈ=Xb=c6=�=��=��=�M=�=g�=`=�=�=;=�=�X=��	=�^=�=~M=f�=�%=!� =���<��<�1�<_��<8l�<���<���<P�<x~�<���<�\�<��<�!�</|�<|��<
"�<*n�<@��<���<P;�<�x�<f��<'�<d �<>S�< ��<۲�<�ߛ<�<�5�<�^�<Ɔ�<��<�Ԅ<;��<�Bz<R�r<P�j<�)c<�x[<�S<,L<|oD<H�<<�5<�|-<��%<�@<r�<�<��<�  <	��;
�;�;�C�;�z�;æ;b�;���;5$v;�YY;|�<;�T ;�;�A�:���:qIC:8;�9�>��v��k�a����ݺG{���!��:�EQS�g�k�4���B������l������������ŻE=лɲڻ��仲�����V�����
��a�#��<Q�y���� �N%�<)�uG-�lA1��*5��9�S�<�D�@�^5D�4�G�LhK���N��kR���U��CY�d�\���_�8Ac���f��i�V�l�[!p��Gs�'hv�a�y�p�|���Y��N܂��]���܅�LZ��+ֈ�oP��[ɋ��@�����,��蟑����i���+���e��Ԙ�7B���������׈������`��ˢ��5��X����
��u��8ߩ�pI������������I򰼔\��ǳ��1��W���.��Wr���ݺ��I�������  �  ��N=��M=!CM=��L=��K=�K=�dJ=��I= �H=�9H=�G=��F=�
F=�OE='�D=��C=7C=�]B=۟A=$�@=�!@=ta?=L�>=P�==H==@W<=%�;=��:=w:=�;9=�q8=_�7=��6=F6=Y;5=�i4=h�3=B�2=��1=�1=D50=pW/="w.=4�-=��,=��+=g�*=��)=l�(=�(=�
'={&=n%=O$=��"=�!=�� =d�=?�=��=wb=x6=�=��=��=�M==X�=`==΢=�:=��=�X=��	=�^=��=UM=@�=�%=�� =U��<���<�1�<%��<l�<g��<���<[�<�~�<���<�\�<B��<"�<l|�<���<G"�<zn�<���<���<�;�<y�<���<S�<� �<[S�<��<벟<�ߛ<j�<�5�<�^�<���<魈<�Ԅ<���<|Bz<��r<��j<O)c<Px[<x�S<�L<oD<��<<�5<>|-<��%<�@<~�<�<�< <���;��;+�;�D�;�{�;=Ħ;��;ӎ�;�&v;
\Y;��<;�V ;V!;�E�:���:�MC:�>�9�>��3��k�������ݺ;|�W�!���:��RS�A�k����G������~���C���Q�����Ż�=лj�ڻ��们ﻻ���oV�B�Y�
��a�����P����"� ��%�u;)��F-��@1�'*5�9���<�ۇ@�5D��G�#hK���N��kR��U�FDY���\�!�_��Ac�H�f���i���l��!p�dHs��hv��y���|�o��IY��v܂��]���܅�ZZ��+ֈ�YP��Aɋ��@��ܶ���+������r��%��������d���Ә��A��z���X������}����_���ʢ��5��M����
��u��gߩ��I��г�����>������\��]ǳ��1������l���r��޺��I��鵽��  �  m�N=��M=CM=��L=��K=�K=�dJ=�I=!�H=�9H= �G=��F=F=�OE=O�D= �C=`C=^B=��A=G�@=�!@=}a?=e�>=Q�==K==AW<=�;=��:=a:=�;9=�q8=B�7=g�6=6=-;5=�i4=A�3=�2=��1=�1=50=VW/=w.=)�-=��,=��+=`�*=��)=~�(=�(=�
'=�&=�%=w$=�"=;�!=�� =��=e�=�=�b=�6==��=��=�M==J�=�_=i=��=�:=��=�X=�	=z^=��=M=�=�%=҉ =���<N��<K1�<���<�k�<S��<���<J�<�~�<���<�\�<���<P"�<�|�<��<�"�<�n�<��<,��<�;�<hy�<ೲ<��<� �<�S�<;��<鲟<�ߛ<X�<u5�<h^�<\��<���<[Ԅ<���<�Az<�r< �j<�(c<}w[<��S<%L<onD<I�<<'5<|-<|�%<�@<u�<�<F�<. <���;��;i�;.F�;F}�;�Ŧ;4!�;y��;�)v;(_Y;}�<;�Y ;�#;�G�:
��:PC:rD�9d.�����k�������ݺU~���!�]�:�RUS���k�p���Z���/��S���9���bº�r�Ż%>л��ڻ��l�����V���#�
��`�4��P�L��i� ��%��:)�GF-�D@1�z)5��9�c�<���@��4D���G�9hK���N��kR�J�U��DY��\���_�4Bc���f�^�i�~�l��"p�Is�Hiv���y�h�|����Y���܂��]���܅�_Z��!ֈ�^P��ɋ��@�������+��j�����҃������id��hӘ��A��$�����e���9����_���ʢ��5��R����
��.u��xߩ��I�����I��|�����8]���ǳ�52�������r��@޺�J��#����  �  Q�N=��M=CM=��L=��K=�K=�dJ=$�I=E�H=�9H='�G=��F=KF=(PE=|�D=R�C=�C=,^B=�A=c�@=�!@=�a?=w�>=V�==T==8W<=�;=��:=F:=�;9=yq8=�7=?�6=�
6=�:5=ii4=�3=��2=��1=s1=50=AW/=�v.="�-=v�,=�+=e�*=��)=��(=�(=�
'=�&=�%=�$=B�"=f�!=�� =��=��=E�=�b=�6= =��=��=�M=�=8�=�_=H=��=�:=��=qX=J�	=G^=j�=�L=ػ=W%=�� =���< ��<1�<���<�k�<.��<���<G�<�~�<��<]�<���<�"�<}�<[��<#�<&o�<@��<���<=<�<�y�<!��<��<� �<�S�<M��<���<�ߛ<?�<`5�<0^�<9��<U��<�ӄ<R��<�@z<^�r<�j<�'c<�v[<(�S<bL<�mD<��<<�5<�{-<<�%<�@<��<�<��<� <���;��;� �;�G�;�~�;�Ǧ;�"�;B��;�,v;>bY;.�<;�[ ;Y&;�K�:n��:}SC:%M�9�/��t�k�D���n�ݺ�����!���:��WS�=�k�����y���w��d�������ú� �Ż�>л˳ڻJ��'ﻝ����U�����
�U`����bO������ �J%�:)�xE-��?1��(5�*9���<��@�|4D�s�G�hK�}�N�lR�d�U��DY�|�\���_��Bc�Q�f��i�!�l�]#p��Is��iv�Z�y��|�����Y���܂��]��݅�uZ��ֈ�SP���ȋ�b@��e���V+��$����������,���d��
Ә�CA��ծ�����'����󟼁_���ʢ��5��E����
��Iu���ߩ��I��(������و��)󰼗]��ȳ��2��F���+��;s���޺�MJ��B����  �  7�N=��M=CM=�L=��K=�K=�dJ=@�I=T�H=
:H=S�G=�F=xF=TPE=��D=}�C=�C=S^B=N�A=��@="@=�a?=��>=c�==R==2W<=�;=��:=&:=m;9=Zq8=�7=�6=�
6=�:5=<i4=�3=��2=��1=Q1=�40=W/=�v.=�-=q�,=��+=p�*=��)=��(=(=�
'=�&=�%=�$=j�"=��!="� =��=��=g�=�b=�6=5=��=��=�M=r=+�=�_=+=e�=x:=`�=?X=�	=
^=4�=�L=��=&%=n� =4��<���<�0�<���<�k�<��<���<R�<�~�<K��<3]�<���<�"�<T}�<���<U#�<�o�<���<���<�<�<z�<w��<	�<+!�<�S�<g��<��<�ߛ<7�<;5�<�]�<<��<�ӄ<���<8@z<��r<c�j<'c< v[<r�S<�L<KmD<c�<<25<t{-<�%<�@<��<<҉< <r �;?
�;0"�;�H�;R��;ɦ;�$�;͓�;0v;eY;��<;[^ ; (;�P�:�:�XC:DP�9�+��~�� k�`���`�ݺ ���!���:�-ZS�˝k�Á�����������������ú���Ż�?л4�ڻ`��[�1����U�?�$�
�`�����N����� ��%�>9)��D-��>1�8(5�k9���<���@�4D�W�G��gK���N�lR���U�:EY� �\���_�yCc���f���i���l�$p��Js��jv��y���|�@���Y��݂�^��݅�Z��ֈ�<P���ȋ�*@��=���$+��Ğ��}��&����󕼩c���Ҙ��@������g��Շ����K_���ʢ�}5��6����
��Su���ߩ�&J��q������ ���|��]��fȳ��2����������s���޺��J�������  �  -�N=��M=�BM=�L=��K=�K=�dJ=U�I=q�H=2:H=o�G=D�F=�F=}PE=ߔD=��C=�C=t^B=n�A=��@="@=�a?=��>=n�==M==6W<=��;=��:=:=K;9=>q8=ɥ7=��6=�
6=�:5=i4=��3=��2=e�1=51=�40=W/=�v.=��-=t�,=��+=s�*=��)=��(=.(=�
'=&=�%=�$=��"=��!=N� =�=�=��=�b=�6=H=��=��=�M=f=+�=�_==L�=M:=>�=X=��	=�]=��=vL=g�=�$=<� =���<i��<�0�<T��<ak�<��<~��<\�<�~�<e��<^]�<*��<(#�<�}�<��<�#�<�o�<��<@��<�<�<Nz�<˴�<J�<Z!�<�S�<���<��<�ߛ<5�<5�<�]�<���<Ӭ�<kӄ<���<�?z<Ƌr<��j<M&c<Mu[<��S<L<�lD<��<<�5<{-<��%<�@<��<G<��<i <i�;��;-#�;PJ�;���;�ʦ;;&�;1��;�3v;�gY;�<;Xa ;%*;�S�:�Ę:O]C:PQ�9���!��#k�������ݺ{��3�!��:��\S�{�k�Nā�5���� ��ˇ��V����ĺ���Ż�?л�ڻ2��w�����U����
��_�M��PN�%��I� ��%��8)�.D-�>1��'5�� 9� �<�R�@��3D�)�G��gK���N�lR���U�pEY�F�\��_��Cc���f�O�i���l��$p�GKs�ikv���y�P�|����6Z��/݂�<^��H݅�tZ��%ֈ�&P���ȋ�@��
����*������?��������Lc��YҘ��@��*���.�������� _��pʢ�h5��9����
��Xu���ߩ�9J������	��f�����9^���ȳ�J3���������s��.ߺ��J��ɶ���  �  �N=��M=�BM=�L=��K=�K=�dJ=f�I=��H=F:H=��G=i�F=�F=�PE= �D=��C=
C=�^B=��A=��@=5"@=�a?=��>=x�==P==/W<=�;=��:=:=6;9=!q8=��7=��6=s
6=�:5=�h4=��3=k�2=E�1=1=�40=�V/=�v.=�-=h�,=��+=z�*=��)=��(=B(='=&=!%=$=��"=��!=m� =*�=�=��=c=�6=Z=��=̐=�M=b=�=�_=�=-�=.:=�=�W=��	=�]=��=ML=A�=�$=� =���<0��<J0�<)��<@k�<���<x��<g�<�~�<���<�]�<X��<X#�<�}�<V��<�#�<,p�<8��<{��<6=�<�z�<���<��<�!�<$T�<���<��<�ߛ<�<�4�<�]�<���<���<(ӄ<_��<�>z<C�r<�j<�%c<�t[<,�S<�L<FlD<y�<<�5<�z-<��%<�@<��<~<Q�<� <_�;A�;8$�;�K�;��;�˦;k'�;v��;	6v;mjY;#�<; c ;,;�V�:xȘ:�aC:�U�9��*#��%k� ����ݺ�����!���:�l^S�E�k�qŁ�����!������U����ź�>�Żd@л<�ڻ~��iﻼ���)U���p�
�	_�����M������ �G%��7)��C-��=1�2'5�g 9���<���@��3D���G��gK���N�/lR�(�U��EY���\�u�_�gDc�!�f���i��l�[%p��Ks��kv��y�˚|�%��bZ��`݂�[^��^݅��Z��"ֈ�P���ȋ��?��ڵ���*��M���������D�c��Ҙ�T@��䭛����]���Y��^��Dʢ�H5��-����
��ou���ߩ�hJ��Ѵ��<����������^��ɳ��3��F���	��&t��mߺ��J��񶽼�  �  �N=��M=�BM=�L=��K=�K=�dJ=o�I=��H=Z:H=��G=�F=�F=�PE=�D=��C=C=�^B=��A=��@=G"@=�a?=��>=u�==W==&W<=�;=��:=�:=';9=q8=��7=��6=N
6=c:5=�h4=w�3=J�2=0�1=�1=�40=�V/=�v.=�-=^�,=��+=y�*=��)=��(=N(=%'=.&=A%=)$=��"=��!=�� =R�=�==!c=7=e=�=Đ=�M=d=�=�_=�=�=:=��=�W=��	=�]=��=)L=�=�$=�� =\��<��<0�<��<<k�<���<���<X�<�~�<���<�]�<x��<�#�<~�<{��<8$�<dp�<���<���<a=�<�z�<��<��<�!�<7T�<���<"��<�ߛ<�<�4�<�]�<j��<o��<�҄<0��<j>z<Êr<y�j<B%c<$t[<��S<%L<�kD<4�<<D5<�z-<��%<}@<��<m<o�<� <��;��;E%�;QL�;��;ͦ;o(�;ٗ�;�7v;dlY;�<;�d ;�-;�X�:�ɘ:�aC:�[�9X��"�%k����I�ݺ����!�<�:��`S���k�fƁ�����"��H���-���ƺ�țŻ�@л��ڻ���@﻽���6U�}�:�
��^����9M�X��)� ��%�}7)� C-�X=1��&5� 9�F�<���@�k3D���G��gK���N�]lR��U��EY���\���_��Dc�t�f�Y�i���l��%p�CLs�xlv���y�&�|����Z���݂�a^��X݅��Z��ֈ�P���ȋ��?�������*��������Y������b���ј�@���������6���8��^��4ʢ�P5��'����
��u���ߩ��J������j��܉��@����^��>ɳ��3������]	��Ut���ߺ�0K������  �  ��N=��M=�BM=�L=��K=�K=�dJ=~�I=��H=h:H=��G=��F=�F=�PE=*�D=��C=/C=�^B=��A=��@=S"@=�a?=��>=��==Y=="W<=ޑ;=z�:=�:=;9=�p8=��7=��6=A
6=V:5=�h4=i�3=:�2=�1=�1=�40=�V/=�v.=ݓ-=X�,=��+=�*=��)=��(=[(=4'=9&=N%=9$=��"=�!=�� =]�="�=ω=)c=7=q=�=͐=�M=c=�=�_=�=	�=
:=��=�W=��	=w]=��=L=�=�$=� =C��<��< 0�<���<k�<���<~��<i�<�<���<�]�<���<�#�<-~�<���<N$�<p�<���<���<�=�<�z�<=��<��<�!�<MT�<���<+��<�ߛ<�
�<�4�<�]�<R��<X��<�҄<��<->z<��r<K�j<%c<�s[<}�S<�L<�kD<��<<#5<�z-<x�%<p@<��<�<��< <[�;f�;�%�;�L�;���;}ͦ;�(�;E��;�8v;hmY;�<;�e ;z.;�Z�:�ʘ:OeC:�]�91#��:%�R)k������ݺ����!�"�:�;aS���k��Ɓ�u���#��É��u���|ƺ��ŻAл��ڻ���5ﻄ���U�M��
��^�m��M����� ��%�G7)��B-�=1�s&5���8��<���@�63D���G��gK���N�llR�`�U�FY��\���_�Ec���f���i���l�&p�wLs��lv�نy�^�|�����Z���݂��^��{݅��Z��ֈ�P���ȋ��?������a*��������7����򕼵b���ј��?��������������^��ʢ�;5������
���u��੼�J������������b����^��]ɳ��3������y	��vt���ߺ�FK��)����  �  ��N=��M=�BM=�L=��K=�K=�dJ=}�I=��H=m:H=��G=��F=�F=�PE=>�D=��C=8C=�^B=��A=��@=O"@=�a?=��>=}�==Q==-W<=�;=|�:=�:=;9=�p8=��7=��6=;
6=F:5=�h4=_�3=4�2=�1=�1=�40=�V/=�v.=ߓ-=e�,=��+={�*=��)=��(=U(=7'=?&=V%=F$=��"=�!=�� =^�=.�=։=/c=7=j=�=ΐ=�M=[=�=�_=�=�=�9=��=�W=}�	=n]=��=L= �=�$=� =>��<˄�<0�<���<*k�<���<l��<a�<�~�<���<�]�<���<�#�<B~�<���<R$�<�p�<���<���<�=�<�z�<I��<��<�!�<BT�<���<!��<�ߛ<�<�4�<�]�<C��<Q��<�҄<���<>z<M�r<�j<�$c<�s[<\�S<�L<�kD<��<<*5<�z-<��%<�@<��<�<��< <V�;��;�%�;GM�;Ą�;�ͦ;�)�;j��;g9v;BnY;��<;f ;E.;sZ�:sʘ:�dC:cZ�9��"��(k����*�ݺ��&�!���:��aS���k�"ǁ���N#����������ƺ��Ż�@л��ڻ���Uﻥ���	U�b��
�z^�V���L����� �L%��6)��B-��<1�R&5���8���<���@�M3D���G��gK���N�7lR�L�U�FY��\��_�Ec�ӈf���i���l�H&p��Ls��lv���y�w�|�ƪ��Z���݂�~^��d݅��Z�� ֈ�P���ȋ��?������Z*���������%����򕼍b���ј��?��������������^��*ʢ�<5��)����
��uu��੼�J������������r����^��vɳ�
4�������	���t���ߺ�HK��<����  �  ��N=��M=�BM=�L=��K=�K=�dJ=~�I=��H=h:H=��G=��F=�F=�PE=*�D=��C=/C=�^B=��A=��@=S"@=�a?=��>=��==Y=="W<=ޑ;=z�:=�:=;9=�p8=��7=��6=A
6=V:5=�h4=i�3=:�2=�1=�1=�40=�V/=�v.=ݓ-=X�,=��+=�*=��)=��(=[(=4'=9&=N%=9$=��"=�!=�� =]�="�=ω=)c=7=q=�=͐=�M=c=�=�_=�=	�=
:=��=�W=��	=w]=��=L=�=�$=� =E��<��<0�<���<k�<���<���<k�<�<���<�]�<���<�#�<.~�<���<O$�<�p�<���<���<=�<�z�<<��<��<�!�<KT�<���<)��<�ߛ<�
�<�4�<�]�<Q��<W��<�҄<��<,>z<��r<K�j<%c<�s[<�S<�L<�kD< �<<&5<�z-<{�%<s@<��<�<��< <`�;k�;�%�;�L�;���;}ͦ;�(�;D��;�8v;`mY;��<;�e ;k.;�Z�:�ʘ:eC:O]�9�%���%��)k�����ݺ(����!�5�:�MaS�ɤk��Ɓ�|���&#��ɉ��{����ƺ�
�ŻAл��ڻ���8ﻆ���U�N��
��^�n��M����� ��%�G7)��B-�=1�s&5���8��<���@�63D���G��gK���N�llR�`�U�FY��\���_�Ec���f���i���l�&p�wLs��lv�نy�^�|�����Z���݂��^��{݅��Z��ֈ�P���ȋ��?������a*��������7����򕼵b���ј��?��������������^��ʢ�;5������
���u��੼�J������������b����^��]ɳ��3������y	��vt���ߺ�FK��)����  �  �N=��M=�BM=�L=��K=�K=�dJ=o�I=��H=Z:H=��G=�F=�F=�PE=�D=��C=C=�^B=��A=��@=G"@=�a?=��>=u�==W==&W<=�;=��:=�:=';9=q8=��7=��6=N
6=c:5=�h4=w�3=J�2=0�1=�1=�40=�V/=�v.=�-=^�,=��+=y�*=��)=��(=N(=%'=.&=A%=)$=��"= �!=�� =R�=�==!c=7=f=�=Đ=�M=d=�=�_=�=�=:=��=�W=��	=�]=��=+L=�=�$=�� =`��<��<0�<��<Ak�<���<���<\�<�~�<���<�]�<{��<�#�<~�<|��<9$�<dp�<���<���<`=�<�z�<��<��<�!�<4T�<���<��<�ߛ<�<�4�<�]�<g��<m��<�҄</��<h>z<r<y�j<C%c<&t[<��S<)L<�kD<9�<<J5<�z-<��%<�@<��<s<u�<� <�;��;K%�;VL�;��;ͦ;m(�;՗�;�7v;TlY;�<;�d ;o-;QX�:=ɘ:`aC:hZ�92$���"��%k������ݺ���C�!�_�:��`S��k�uƁ�#����"��S���8���(ƺ�ЛŻ�@л�ڻ���F�����8U��;�
��^����:M�Y��*� ��%�}7)� C-�X=1��&5� 9�F�<���@�k3D���G��gK���N�]lR��U��EY���\���_��Dc�t�f�Y�i���l��%p�CLs�xlv���y�&�|����Z���݂�a^��X݅��Z��ֈ�P���ȋ��?�������*��������Y������b���ј�@���������6���8��^��4ʢ�P5��'����
��u���ߩ��J������j��܉��@����^��>ɳ��3������]	��Ut���ߺ�0K������  �  �N=��M=�BM=�L=��K=�K=�dJ=f�I=��H=F:H=��G=i�F=�F=�PE= �D=��C=
C=�^B=��A=��@=5"@=�a?=��>=x�==P==/W<=�;=��:=:=6;9=!q8=��7=��6=s
6=�:5=�h4=��3=k�2=E�1=1=�40=�V/=�v.=�-=h�,=��+=z�*=��)=��(=B(='=&=!%=$=��"=��!=m� =+�=�=��=c=�6=Z=��=̐=�M=c=�=�_=�=.�=0:=�=�W=��	=�]=��=OL=D�=�$=� =���<6��<Q0�</��<Fk�<���<~��<m�<�~�<���<�]�<\��<\#�<�}�<X��<�#�<-p�<7��<z��<4=�<�z�<�<��<~!�< T�<���<��<�ߛ<�<�4�<�]�<���<���<%ӄ<]��<�>z<A�r<�j<�%c<�t[<0�S<�L<LlD<��<<�5<�z-<��%<�@<��<�<Y�<� <m�;M�;A$�;�K�;��;�˦;i'�;p��;�5v;VjY;�<;�b ;�+;�V�:Ș:�`C:)T�9���
$��&k�� ��9�ݺ0��	�!���:��^S�s�k��Ł�(����!��ǈ��e����ź�J�Żo@лF�ڻ���q�����,U���r�
�_�����M������ �H%��7)��C-��=1�2'5�g 9���<���@��3D���G��gK���N�/lR�(�U��EY���\�u�_�gDc�!�f���i��l�[%p��Ks��kv��y�˚|�%��bZ��`݂�[^��^݅��Z��"ֈ�P���ȋ��?��ڵ���*��M���������D�c��Ҙ�T@��䭛����]���Y��^��Dʢ�H5��-����
��ou���ߩ�hJ��Ѵ��<����������^��ɳ��3��F���	��&t��mߺ��J��񶽼�  �  -�N=��M=�BM=�L=��K=�K=�dJ=U�I=q�H=2:H=o�G=D�F=�F=}PE=ߔD=��C=�C=t^B=n�A=��@="@=�a?=��>=n�==M==6W<=��;=��:=:=K;9=>q8=ɥ7=��6=�
6=�:5=i4=��3=��2=e�1=51=�40=W/=�v.=��-=t�,=��+=s�*=��)=��(=.(=�
'=&=�%=�$=��"=��!=N� =�=�=��=�b=�6=H=��=��=�M=g=,�=�_==N�=O:=@�=X=��	=�]=�=yL=k�=�$=?� =���<q��<�0�<\��<ik�<��<���<c�<�~�<k��<c]�</��<,#�<�}�< ��<�#�<�o�<��<>��<�<�<Lz�<Ǵ�<F�<V!�<�S�<{��<��<�ߛ<0�<5�<�]�<���<Ь�<hӄ<���<�?z<ŋr<��j<O&c<Qu[<��S<%L<�lD<��<<5<{-<�%<�@<��<R< �<r <z�;��;9#�;XJ�;���;�ʦ;9&�;*��;�3v;�gY;��<;.a ;�);kS�:JĘ:X\C:IO�9l���"� %k�5���_�ݺ���t�!�1�:��\S���k�hā�M���� ��߇��i���ź���Ż�?л�ڻ<�什�����U�	���
��_�O��RN�&��K� ��%��8)�/D-�>1��'5�� 9� �<�S�@��3D�)�G��gK���N�lR���U�pEY�F�\��_��Cc���f�O�i���l��$p�GKs�ikv���y�P�|����6Z��/݂�<^��H݅�tZ��%ֈ�&P���ȋ�@��
����*������?��������Lc��YҘ��@��*���.�������� _��pʢ�h5��9����
��Xu���ߩ�9J������	��f�����9^���ȳ�J3���������s��.ߺ��J��ɶ���  �  7�N=��M=CM=�L=��K=�K=�dJ=@�I=T�H=
:H=S�G=�F=xF=TPE=��D=}�C=�C=S^B=N�A=��@="@=�a?=��>=c�==R==2W<=�;=��:=&:=m;9=Zq8=�7=�6=�
6=�:5=<i4=�3=��2=��1=Q1=�40=W/=�v.=�-=q�,=��+=p�*=��)=��(=(=�
'=�&=�%=�$=j�"=��!="� =��=��=h�=�b=�6=6=��=��=�M=s=-�=�_=-=g�=z:=b�=AX=�	=^=7�=�L=��=*%=r� =<��<Ʌ�<�0�<���<�k�<��<���<Z�<�~�<R��<9]�<���<�"�<X}�<���<W#�<�o�<���<���<�<�<z�<s��<�<&!�<�S�<a��<��<�ߛ<1�<55�<�]�<ꅌ<��<�ӄ<���<4@z<��r<c�j<'c<v[<x�S<�L<SmD<m�<<>5<�{-<+�%<�@<��<)<މ< <� �;O
�;="�;�H�;W��;ɦ;�$�;Ɠ�; 0v;�dY;u�<;-^ ;�';P�:+:�WC: N�965��� ��!k�������ݺk��_�!�۽:�oZS�	�k�8Á����������������ú��Ż�?лA�ڻk��e�:����U�B�'�
�`�����N����� ��%�?9)��D-��>1�9(5�l9���<���@�4D�W�G��gK���N�lR���U�:EY� �\���_�yCc���f���i���l�$p��Js��jv��y���|�@���Y��݂�^��݅�Z��ֈ�<P���ȋ�*@��=���$+��Ğ��}��&����󕼩c���Ҙ��@������g��Շ����K_���ʢ�}5��6����
��Su���ߩ�&J��q������ ���|��]��fȳ��2����������s���޺��J�������  �  Q�N=��M=CM=��L=��K=�K=�dJ=$�I=E�H=�9H='�G=��F=KF=(PE=|�D=R�C=�C=,^B=�A=c�@=�!@=�a?=w�>=V�==T==8W<=�;=��:=F:=�;9=yq8=�7=?�6=�
6=�:5=ii4=�3=��2=��1=s1=50=AW/=�v.="�-=v�,=�+=e�*=��)=��(=�(=�
'=�&=�%=�$=B�"=f�!=�� =��=��=F�=�b=�6= =��=��=�M=�=9�=�_=J=��=�:=��=tX=M�	=J^=m�=�L=ܻ=Z%=�� =���<)��<1�<���<�k�<7��<���<P�<�~�<$��<]�<���<�"�<}�<^��<#�<&o�<?��<���<;<�<�y�<��<��<� �<�S�<G��<�<�ߛ<9�<Z5�<*^�<4��<P��<�ӄ<O��<�@z<\�r<�j<�'c<�v[<.�S<jL<�mD<�<<�5<�{-<I�%<�@<��<�<��<� < �;	�;� �;�G�;�~�;�Ǧ;�"�;:��;�,v;bY;�<;�[ ;"&;�K�:还:_RC:�J�9�9��� �Mk������ݺ׀�1�!�ɻ:��WS�}�k������������|�������ú��Ż�>лٳڻV��2ﻦ����U�����
�X`����cO������ �K%�:)�xE-��?1��(5�*9���<��@�|4D�t�G�hK�}�N�lR�d�U��DY�|�\���_��Bc�Q�f��i�!�l�]#p��Is��iv�Z�y��|�����Y���܂��]��݅�uZ��ֈ�SP���ȋ�b@��e���V+��$����������,���d��
Ә�CA��ծ�����'����󟼁_���ʢ��5��E����
��Iu���ߩ��I��(������و��)󰼗]��ȳ��2��F���+��;s���޺�MJ��B����  �  m�N=��M=CM=��L=��K=�K=�dJ=�I=!�H=�9H= �G=��F=F=�OE=O�D= �C=`C=^B=��A=G�@=�!@=}a?=e�>=Q�==K==AW<=�;=��:=a:=�;9=�q8=B�7=g�6=6=-;5=�i4=A�3=�2=��1=�1=50=VW/=w.=)�-=��,=��+=`�*=��)=~�(=�(=�
'=�&=�%=x$=�"=<�!=�� =��=e�=�=�b=�6==��=��=�M=�=K�=�_=j=��=�:=��=�X=��	=}^=��=!M=�=�%=։ =���<V��<T1�<��<�k�<\��<���<R�<�~�<���<�\�<���<T"�<�|�<��<�"�<�n�<��<+��<�;�<ey�<ܳ�<��<� �<�S�<5��<㲟<�ߛ<R�<o5�<c^�<W��<���<XԄ<���<�Az<�r< �j<�(c<�w[<��S<,L<xnD<S�<<25<|-<��%<�@<��<�<R�<9 <���;�;v�;8F�;K}�;�Ŧ;2!�;r��;�)v;	_Y;V�<;~Y ;V#;IG�:���:OC:/B�9�7����k�m���O�ݺ�~��!���:��US���k�����u���H��j���N���uº���Ż4>л��ڻ��w�����V���&�
��`�6��P�M��j� � %��:)�HF-�D@1�{)5��9�d�<���@��4D���G�9hK���N��kR�J�U��DY��\���_�4Bc���f�^�i�~�l��"p�Is�Hiv���y�h�|����Y���܂��]���܅�_Z��!ֈ�^P��ɋ��@�������+��j�����҃������id��hӘ��A��$�����e���9����_���ʢ��5��R����
��.u��xߩ��I�����I��|�����8]���ǳ�52�������r��@޺�J��#����  �  ��N=��M=!CM=��L=��K=�K=�dJ=��I= �H=�9H=�G=��F=�
F=�OE='�D=��C=7C=�]B=۟A=$�@=�!@=ta?=L�>=P�==H==@W<=%�;=��:=w:=�;9=�q8=_�7=��6=F6=Y;5=�i4=h�3=B�2=��1=�1=D50=pW/="w.=4�-=��,=��+=g�*=��)=l�(=�(=�
'={&=n%=O$=��"=�!=�� =e�=?�=��=xb=x6=�=��=��=�M=�=Y�=`=�=Т=�:=��=�X=��	=�^=��=XM=C�=�%=�� =\��<���<�1�<-��<
l�<n��<���<b�<�~�<���<�\�<G��<"�<o|�<���<H"�<{n�<���<���<�;�<y�<���<O�<� �<VS�<��<岟<�ߛ<e�<~5�<�^�<���<孈<�Ԅ<���<yBz<��r<��j<Q)c<Tx[<}�S<�L<'oD<��<<�5<I|-<��%<�@<��<�<��< <���;��;7�;�D�;�{�;?Ħ;��;͎�;�&v;�[Y;��<;�V ;&!;0E�:���:�LC:�<�9EG��F��k�z���>�ݺ~|���!���:�	SS�y�k�9���`����������V���b���ϗŻ�=лv�ڻ��仵�����rV�E�[�
��a�����P����#� ��%�u;)��F-��@1�(*5�9���<�܇@�5D��G�#hK���N��kR��U�FDY���\�!�_��Ac�H�f���i���l��!p�dHs��hv��y���|�o��JY��v܂��]���܅�ZZ��+ֈ�YP��Aɋ��@��ܶ���+������r��%��������d���Ә��A��z���X������}����_���ʢ��5��M����
��u��gߩ��I��г�����>������\��]ǳ��1������l���r��޺��I��鵽��  �  ��N=�M=.CM=��L=��K=�K=wdJ=�I=��H=�9H=�G=��F=�
F=�OE= �D=��C=C=�]B=��A=
�@=�!@=^a?=@�>=F�==H==GW<=6�;=��:=�:=�;9=�q8=�7=��6=c6={;5=�i4=��3=_�2=$�1=�1=_50=�W/=2w.=J�-=��,=��+=^�*=��)=\�(=�(=m
'=\&=P%=1$=��"=��!=z� =I�="�=ۈ=Yb=c6=�=��=��=�M=�=h�=`=�=�=;=�=�X=��	=�^=�=�M=i�=�%=$� =���<���<�1�<f��<?l�<���<���<V�<}~�<���<�\�<��<�!�<2|�<~��<"�<+n�<@��<���<N;�<�x�<d��<#�<` �<:S�<���<ײ�<�ߛ<z�<�5�<�^�<Æ�<��<�Ԅ<9��<�Bz<P�r<Q�j<�)c<�x[<�S<2L<�oD<O�<<�5<�|-<��%<A<{�<�<Ȉ<�  <��;�;)�;�C�;�z�;æ;`�;���;%$v;�YY;`�<;�T ;�;�A�:2��:�HC:�9�9�E��W��k�������ݺ~{���!��:�uQS���k�I���V������}�����������*�ŻP=лӲڻ��仺�����V�����
��a�%��=Q�z���� �N%�<)�uG-�lA1��*5��9�S�<�D�@�^5D�5�G�LhK���N��kR���U��CY�d�\���_�8Ac���f��i�V�l�[!p��Gs�'hv�a�y�p�|���Y��N܂��]���܅�LZ��+ֈ�oP��[ɋ��@�����,��蟑����i���+���e��Ԙ�7B���������׈������`��ˢ��5��X����
��u��8ߩ�pI������������I򰼔\��ǳ��1��W���.��Wr���ݺ��I�������  �  ��N=�M=*CM=�L=��K=�K={dJ=ӫI=��H=p9H=�G=g�F=�
F=�OE=ܓD=��C=�C=�]B=��A=��@=�!@=Na?=E�>=<�==H==IW<=2�;= �:=�:=�;9=�q8=��7=��6=�6=�;5=j4=��3=r�2=C�1=�1=p50=�W/=<w.=I�-=��,=��+=S�*=��)=X�(=�(=_
'=?&=;%=$=��"=��!=]� =$�=�=ǈ==b=X6=�=��=��=�M=�=h�=`=�= �=$;=,�=Y=��	=_=,�=�M=��=&=K� =���<��<�1�<���<?l�<���<τ�<I�<�~�<���<m\�<���<�!�<|�<?��<�!�<�m�<��<D��<;�<�x�<'��<�<2 �<:S�<���<ǲ�<�ߛ<r�<�5�<�^�<熌<:��<Մ<n��<ZCz<��r<��j<�*c<Jy[<��S<�L<�oD<��<<	 5<�|-<��%<A<m�<�<Ԉ<[  <���;/�;I�;�B�;xy�;¦;(�;���;�!v;�WY;d�<;-S ;;�>�:A��:EC:B7�9qK��n��k�.���]�ݺ�z��!��:�OS�t�k�}���)���^������︯�&�����Ż=л�ڻ��仇�y����V���$�
�#b�����Q����7� ��%��<)�H-��A1��*5�9���<���@�|5D��G�|hK���N��kR���U��CY�'�\�o�_��@c�1�f�ʿi���l�� p�SGs��gv��y��|�ɦ��X��7܂�n]���܅�MZ��&ֈ��P��Pɋ��@��,���3,��!����������n���Pe��CԘ��B��𯛼����������-`��ˢ��5��g����
��	u��.ߩ�_I��w������͇���h\���Ƴ�]1��������)r���ݺ�bI�������  �  ��N=�M=4CM=�L=}�K=�K=edJ=̫I=��H=f9H=�G=W�F=�
F={OE=ғD=��C=�C=�]B=��A=��@=!@=Ea?=0�>=3�==F==MW<=<�;=�:=�:=�;9=r8=��7=��6=�6=�;5=j4=��3=��2=R�1=1=50=�W/=Kw.=U�-=��,=�+=O�*=v�)=G�(=�(=R
'=6&=-%=$=��"=��!=R� =�=�=��=4b=K6=�=��=��=�M=�=s�=,`=�=�=7;=9�=+Y=�	=_==�=�M=��=&=\� =���<B��<2�<���<Vl�<���<ӄ�<?�<i~�<���<]\�<���<�!�<�{�<!��<�!�<�m�<��<*��<�:�<�x�<��<��<& �<S�<ۃ�<���<�ߛ<��<�5�<�^�< ��<Y��<&Մ<���<�Cz<'�r<�j<�*c<�y[<��S<�L<pD<��<<G 5<�|-<�%</A<`�<R<{�<>  <&��;��;��;:B�;�x�;���;��;��;� v;�VY;n�<;NR ;D;~=�:@��:'BC:�4�9DG����yk�����ݺ�y�a�!�#�:��NS�ґk����ق�����(�����������P�Ż�<л��ڻq�仃ﻧ����V���?�
�\b�����Q�@��h� ��%��<)�=H-�7B1�:+5�@9���<���@��5D�m�G��hK���N��kR���U��CY��\�/�_��@c���f���i���l�� p�$Gs�Xgv�ցy���|�����X��܂�W]���܅�AZ��&ֈ��P��yɋ�A��?���L,��7������Ȅ������be��^Ԙ��B��������%�������9`��:ˢ��5��o����
���t��ߩ�BI��_������������H\���Ƴ�C1��󛶼���r��tݺ�FI��u����  �  �N=1 N=0JM=ۓL=@�K=L&K=�nJ=4�I=�H=�FH=ƍG=��F=�F=�`E=A�D=G�C=�/C=�sB=�A=��@=�;@=}?=|�>=�==�;==Iy<=�;=Y�:=�+:=�d9=��8=(�7=M7=�;6=n5=��4=Y�3=W�2=^%2=XN1=*u0=��/=��.=&�-=��,=�,=�(+=%<*=dL)=*Y(=@b'=�g&=�h%=f$=�^#=_S"=C!=	. =�=��=��=��=�u=�?=�=��=My=�*=��=z=-=ܯ= A=�=�P
=c�=�G=��=�'=��=�� =��<SJ�<���<���<��<��<"+�<���<T�<1��<g��<H�<ˡ�<���<�D�<���<���<p�<�T�<p��<Ƕ<���<�-�<{]�<Ŋ�<��<jߟ<��<%-�<�Q�<�u�<Y��<P��<�ۄ<���<u;z<5}r<��j<�c<�F[<w�S<��K<cD<ii<<'�4<�	-<_%<��<H<w<��<���;�w�;i�;7h�;�v�;���;<Ƥ;�	�;a�;��q;ءT;��7;�?;y��:Fa�:�|�:�%,:�#y9m:��B�o��l%��1@��\�B�(���A���Z���r�v��F��=圻wS��	�������sɻEԻЍ޻[���������49����Ϣ�%5�Ͱ���zg�p�"�r�&��*���.��2��6��:��>>� �A�M�E�Y&I���L��+P�9�S�4W�aZ���]��`�Ad�{g�`�j���m���p��t��2w��Dz��Q}�-������m.��*���(��Z�����F���[��}������c��`ԑ��D������Z"��㏗�����_h���ӛ�$>���������z���㢼\L��䴥�h������bV��Ͼ��B'��Ǐ��M����`���ɳ��2���������Vn�� غ�4B�������  �  �N=7 N=3JM=�L=<�K=<&K=�nJ=:�I=#�H=�FH=ύG=��F=�F=�`E=R�D=S�C=�/C=�sB=�A=��@=�;@=}?=|�>=�==�;==Oy<=�;=`�:=�+:=�d9=��8=!�7=<7=�;6=n5=��4=V�3=G�2=Q%2=NN1="u0=��/=��.=,�-=��,=�,=�(+=<*=iL)=2Y(=Ob'=�g&=�h%=#f$=_#=pS"=-C!=. =�=��=��=��=�u=�?=�=��=Ty=�*=��=z=*=ѯ=A=
�=�P
=\�=�G=��=�'=��=�� =��<>J�<���<���<��<��<%+�<f��<M�<:��<|��<�H�<ԡ�<���<�D�<Ύ�<���<��<�T�<���<&Ƕ<���<�-�<�]�<Ί�<���<`ߟ<	�<--�<�Q�<�u�<P��<D��<�ۄ<���<?;z< }r<O�j<jc<�F[<8�S<��K<@D<Li<<�4<�	-<_%<�<5<�v<��<͓�;x�;<i�;~h�;$w�;�;�Ƥ;
�;�a�;�q;��T;j�7;�@;z��:fb�:�|�:�!,:�'y9�:�UA��m���%���@�]���(���A��Z�z�r�v��*F���圻�S��T�������$sɻKԻ��޻+�軔��4���R9��������4������Sg�I�"�,�&���*���.���2�Ͱ6�~:��>>���A�;�E�r&I���L��+P�"�S�%W�aZ���]�/�`�BAd�<{g���j���m�%�p�
t��2w�3Ez�R}�-��ͮ��u.�����(��N�����k���_��}�������b��Uԑ��D������E"������d���Sh��yӛ�>���������z���㢼vL��𴥼V������lV��ؾ��O'��Տ��i���a���ɳ��2���������tn��.غ�CB�������  �  ۵N=) N=#JM=��L=D�K=G&K=�nJ=>�I=/�H=�FH=�G=��F=�F=�`E=_�D=g�C=�/C=�sB=+�A=��@=�;@=}?=��>=�==�;==Iy<=ӵ;=Q�:=�+:=�d9=��8=�7=)7=�;6=�m5=r�4=A�3=/�2=C%2=?N1=u0=��/=��.=�-=��,=�,=�(+=.<*=xL)=7Y(=^b'=�g&=i%=:f$=_#=~S"=;C!=&. ==��=��=��=�u=�?=�=��=Uy=�*=��=z==��=�@=��=�P
=C�=�G=��=s'=ǎ=�� =՚�<J�<���<���<��<���<,+�<r��<o�<G��<���<�H�<��<���<�D�<���<���<��<�T�<���<SǶ<��<.�<�]�<���<��<rߟ<	�<-�<�Q�<|u�<7��< ��<�ۄ<���<�:z<�|r<��j<c<9F[<�S<t�K<�D<i<<��4<�	-<�^%<�<Q<w<��<��;ix�;�i�;+i�; x�;���;vǤ;�
�;?b�;��q;��T;��7;�A;M��:�c�:��:�%,:�4y9�:�*D�o��:'��B��]�(�(���A�?�Z�j�r��v���F��]朻1T������<���xsɻ�Ի��޻���y������9�a������4����T��f���"���&���*�h�.�~�2�n�6�A:�G>>���A��E�$&I�ۮL��+P�S�S�VW�TaZ�ٴ]�w�`��Ad�u{g���j��m�l�p�Pt�+3w��Ez�FR}�5-����.��?���-(��_�����X���6���|�������b��6ԑ�hD��Ƴ��"������?���(h��Gӛ��=����������z���㢼ZL��ᴥ�Y��х��(�V��񾬼r'����������Aa���ɳ��2��蛶�&���n��Hغ�gB��Ь���  �  εN= N=)JM=ۓL=C�K=M&K=�nJ=S�I=G�H=�FH=�G=��F=%F=aE=��D=��C=	0C=�sB=O�A=�@=�;@=,}?=��>=�==�;==Ey<=ص;=B�:=�+:=�d9=m�8=��7=7=�;6=�m5=L�4=�3=�2=%2=N1=�t0=|�/=��.=�-=��,=�,=�(+=/<*=�L)=NY(=wb'=�g&="i%=Yf$=A_#=�S"=iC!=M. =$=��=�=��=�u=�?=�=��=Hy=�*=�=�y=�=��=�@=��=�P
=�=�G=M�=<'=��=�� =���<�I�<L��<[��<�<��<+�<y��<^�<Z��<���<�H�<7��< ��<E�<H��<.��<�<9U�<���<�Ƕ<U��<F.�<�]�<��<*��<zߟ<�<-�<�Q�<cu�<��<幈<Gۄ<K��<L:z<�{r<d�j<Jc<�E[<U�S<��K<nD<�h<<�4<r	-<�^%<�<F<w<��<���;,y�;�j�;?j�;�x�;��;�Ȥ;N�;�c�;w�q;��T;y�7;xD;M��:�f�:���:x),:"5y9:�A�0p��n(���D�|_�M�(�Q�A���Z���r�x��;H��,眻QU���������1tɻ#Ի�޻n�軡������8�9��.��:4�ݯ���mf�P�"�4�&���*���.���2��6��~:��=>�Y�A�ԐE�%&I���L��+P�X�S�_W��aZ�;�]���`�Bd�|g�l�j���m��p��t��3w��Ez��R}�s-��%����.��a���'(��f�����E���<���|��M����b���ӑ�0D��z����!��@��������g��ӛ��=������U���z���㢼QL��ݴ��c��ą��9�V��(����'��6��������a��^ʳ�+3��G���q���n���غ��B������  �  ��N= N=JM=דL=K�K=`&K=oJ=z�I=b�H=�FH=-�G=��F=TF=AaE=æD=��C=80C=#tB=w�A=�@=<@=S}?=��>=)�==�;==@y<=Ƶ;=(�:=w+:=~d9=R�8=��7=�7=;6=�m5= �4=��3=��2=�$2=�M1=�t0=c�/=~�.=��-=��,=�,=�(+=@<*=�L)=pY(=�b'=�g&=Li%=�f$=l_#=�S"=�C!=u. =S=��=5�=ԥ=�u=�?=�=��=By=�*=_�=�y=�=p�=�@=��=LP
=��=iG=�='=j�=S� =:��<wI�<��<��<H�<Ũ�<+�<���<{�<���<���<I�<���<q��<`E�<���<���<g�<�U�<_��<�Ƕ<���<~.�<^�<8��<T��<�ߟ<��<-�<�Q�<8u�<Ǘ�<���<�ڄ<���<�9z<0{r<��j< c<�D[<v�S<�K<�D<h<<�4<�-<�^%<ӷ<[<\w<G�<Е�;z�;�k�;�k�;�z�;���;`ʤ;�;4e�;�q;�T;x�7;�F;���:�l�:d��:�/,:�Cy9�:�vC�Yr��.*���G뺵`���(���A���Z���r�By���I��G蜻�V������֜���tɻ�ԻЎ޻��軒��P����8��������3�L��)��e���"�n�&� �*��.�0�2�S�6�~:�|=>���A�b�E��%I���L��+P�m�S��W��aZ���]�` a�|Bd��|g��j���m���p��t��4w��Fz��S}��-��e����.������M(��p�����(������|�����lb���ӑ��C�����x!��ߎ������wg���қ�P=��h���!��Mz��a㢼,L��д��k��߅��q�V��b����'������=����a���ʳ��3���������Bo���غ��B��E����  �  ��N=��M=JM=ٓL=K�K=i&K=+oJ=��I=��H=+GH=`�G=-�F=�F=�aE=��D=��C=t0C=YtB=��A=O�@=7<@=`}?=��>=,�==�;===y<=��;=�:=V+:=Td9=�8=��7=�7=F;6=Zm5=ݝ4=��3=��2=�$2=�M1=�t0=A�/=f�.=��-=��,=�,=�(+=T<*=�L)=�Y(=�b'=h&=�i%=�f$=�_#=T"=�C!=�. =�=%�=[�=�=�u=�?=�=��=@y=z*=J�=�y=�=5�=u@=V�=P
=��=G=ǹ=�&='�= � =���<I�<���<��<�<���<+�<x��<��<���<��<kI�<Ԣ�<���<�E�<��< ��<��<V�<ː�<Zȶ<���<�.�<A^�<i��<u��<�ߟ<
�<�,�<�Q�<u�<���<B��<�ڄ<���<�8z<9zr<��j<��b<�C[<��S<P�K<D<^g<<��4<�-<\^%<η<V<|w<��<D��;r{�;tm�;Vm�;`|�;���;�̤;�;zg�;,�q;�T;�7;XJ;���:�o�:Ԉ�:%3,:�Ry9�:��D�s��-��	L�gc���(���A��Z��r�'{�� K��ꜻ�W��퓳�L����uɻgԻ�޻���P��M���N8�r��9��3����N��d���"�|�&��*��.�C�2�x�6�[}:��<>�o�A� �E�z%I���L��+P���S��W�DbZ��]�"a�?Cd��}g��j�b�m���p��t�q5w��Gz�QT}�.������&/������j(��w��� ��(������v|���b��?ӑ�oC������� ��n������g��Cқ��<��������*z��6㢼L��д��d�������W������N(��㐯�����Ob��1˳�4�����<���o��Bٺ�@C�������  �  o�N=��M=�IM=ГL=O�K=v&K=GoJ=��I=��H=XGH=��G=d�F=�F=�aE=;�D=:�C=�0C=�tB=طA={�@=d<@=x}?=ֽ>=7�==�;==0y<=��;= �:=,+:=7d9=�8=^�7=g7=;6="m5=��4=n�3=l�2=�$2=�M1=�t0=�/=@�.=��-=��,=�,=�(+=e<*=�L)=�Y(=�b'=Ih&=�i%=�f$=�_#=MT"=
D!=�. =�=Y�=��=+�=v=�?=�=��=6y=]*=4�=�y=~=�=3@=�=�O
=F�=�F=��=v&=ڍ=�� =;��<�H�<I��<���<��<v��<�*�<}��<��<ʄ�<g��<�I�<.��<B��<?F�<���<���<i�<�V�<=��<�ȶ<W��<B/�<�^�<���<���<�ߟ<�<�,�<jQ�<�t�<@��<���<%ڄ<��<�7z<Vyr<��j<��b<�B[<��S<b�K<TD<�f<<ӵ4<^-<^%<��<\<�w<�<5��;�|�;�n�;o�;D~�;���;�Τ;I�;�i�;/�q;�T;��7;�M;���:)t�:���:�8,:<_y9K:��E��t��-1���N��e���(�0�A���Z��r��|���L���뜻�Y������.����vɻtԻX�޻N��O������7������G2�٭�h��c���"���&��*��.�m�2���6��|:��;>���A���E�+%I�u�L��+P�֝S�'W��bZ���]��a�Dd�^~g��j�H�m�� q��t�m6w��Hz�$U}�x.������x/��묄��(���������������D|��}�a���ґ��B��4���z ��퍗������f���ћ��<������i���y��㢼�K��ƴ��p������bW��鿬��(��P�������b���˳��4���������p���ٺ��C��̭���  �  S�N=��M=�IM=͓L=Y�K=�&K=[oJ=зI=��H=�GH=ɎG=��F=	F=�aE=x�D=o�C=�0C=�tB=�A=��@=�<@=�}?=�>=J�==�;==+y<=��;=��:=+:=
d9=��8=(�7=17=�:6=�l5=`�4=.�3=6�2=M$2=dM1=Ut0=�/='�.=��-=��,=�,=�(+=s<*=�L)=�Y(=c'=}h&=�i%=0g$=`#=�T"=CD!="/ =�=��=��=C�=#v=@=�=��=/y=L*=�=cy=M=ծ=�?=��=wO
=��=�F=5�=,&=��=�� =Ƙ�<DH�<���<K��<��<V��<�*�<���<��<
��<���<�I�<���<���<�F�<���<���<��<W�<���<8ɶ<���<�/�<�^�<؋�<���<�ߟ<�<�,�<6Q�<|t�<斌<���<�ل<���<�6z<Kxr<u�j<��b<�A[<��S<��K<�D<	f<<Q�4<�-<�]%<��<{<�w<^�<���;�}�;]p�;�p�;]��;;�Ф;q�;�k�;ذq;K�T;��7;�P;B��:�z�:Đ�:L@,:oy9w:�rG��v���3��(S�=h���(�!�A���Z���r��~��~N��^휻%[��䖳�j����wɻ Ի�޻���B��]����7��������1�������b���"���&�#�*�0�.�j�2���6��{:�;>�9�A�-�E��$I�%�L��+P���S�xW�7cZ�R�]�La��Dd�@g�ٱj�F�m��q��t�a7w�\Iz�V}��.��P����/������(���������ꑊ�����{��6la��oґ��B������ ��s���&���f��Vћ�<��W���/���y���⢼�K������u��4�����W��C����(������x���@c��̳�5�����.���p��ں��C��(����  �  F�N=��M=�IM=̓L=X�K=�&K=foJ=�I=��H=�GH=��G=��F=CF=3bE=��D=��C=(1C=�tB=?�A=��@=�<@=�}?=�>=U�==�;==+y<=��;=��:=�*:=�c9=��8=��7=�7=�:6=�l5='�4=��3=��2=$2=7M1="t0=Ә/=�.=��-=��,=�,=�(+=�<*=�L)=�Y(=2c'=�h&=j%=fg$=Q`#=�T"=�D!=V/ =/=��=��=m�=@v=!@=�=��="y=F*=��=Jy='=��=�?=��=0O
=��=@F=�=�%=V�=Z� =[��<�G�<���<��<p�<H��<�*�<���<��<1��<���<RJ�<��<���<3G�<o��<���<T�<�W�<#��<�ɶ<(��<�/�<"_�<���<޶�<�ߟ<��<�,�<Q�<dt�<���<8��<Zل<&��<�5z<<wr<��j<s�b<�@[<ІS<��K<�D<Pe<<�4<s-<�]%<y�<q<x<��<���;.�;r�;ar�;���;롳;�Ҥ;��;�m�;�q;r�T;��7;�T;���:U�:D��:�E,:uy9q�9�I�ux��=5��
X뺅j�v�(���A�8�Z�+s�E���OP��$�\��,���桾��xɻ}Ի��޻f��\��'���u7�/��i��1�-�����a�͝"���&��*�Q�.�{�2��6��z:��:>���A�َE��$I��L��+P��S��W�wcZ���]�a��Ed��g�ʲj�>�m��q�� t�M8w�4Jz��V}�)/�������/��C����(������ ��ؑ������{���a��ґ�=B��9������쌗������e���Л��;������Zy���⢼�K������|��;���塚�W������S)����������c���̳�w5����������p��wں�JD��{����  �  �N=��M=�IM=œL=\�K=�&K=�oJ=�I= I=�GH="�G=�F=oF=cbE=�D=��C=P1C=*uB=e�A=��@=�<@=�}?=�>=a�==�;==$y<=v�;=��:=�*:=�c9=s�8=��7=�7=a:6=wl5=��4=��3=��2=�#2=M1=
t0=��/=��.=��-=��,=�,=�(+=�<*=M)=Z(=Pc'=�h&=Aj%=�g$=|`#=�T"=�D!=�/ =X=��= �=��=Rv=1@==��=y=4*=��=%y==w�=�?=[�=�N
=~�=F=��=�%=�=%� =��<�G�<U��<ɉ�<>�<)��<�*�<���<�<V��<��<�J�<2��<`��<G�<ɑ�<���<��<�W�<���<�ɶ<a��<0�<S_�<3��<��<�ߟ<��<�,�<�P�<t�<_��<��<ل<���<�4z<�vr<��j<��b<@[<	�S<��K<CD<�d<<b�4<-<L]%<W�<~<Yx<��<E��;6��;s�;�s�;���;q��;sԤ;b�;ko�;�q;5�T;W�7;�V;h��:&��:×�:�J,:a�y9��9��K��z��)9��oZ�9l���(���A�̥Z��s�����mQ�����]��I��������yɻqԻ5�޻���[�����7�������0�����?a��"���&�\�*���.���2�K�6�{z:�F:>�R�A���E�a$I���L��+P��S�'W��cZ�:�]�wa�Fd�Àg���j���m�Zq�G!t�9w��Jz��W}�o/��㰁�.0��y����(���������ő��G���{����`���ё��A��바�=������L���Be���Л�c;���������-y���⢼�K���������^���6塚�W�������)��d���=���d���̳��5��ޞ����Kq���ں��D�������  �  
�N=��M=�IM=ǓL=a�K=�&K=�oJ=�I=: I=�GH=G�G=%�F=�F=�bE=�D=�C=r1C=QuB=��A=�@=�<@=�}?=�>=\�==�;==!y<=s�;=��:=�*:=�c9=K�8=��7=�7=7:6=Ll5=Ɯ4=��3=��2=�#2=�L1=�s0=��/=�.=��-=��,=�,=�(+=�<*=M)=Z(=kc'=�h&=ij%=�g$=�`#=U"=�D!=�/ =q=�=�=��=fv=?@==��=y=%*=��=y=�=U�=c?=9�=�N
=N�=�E=��=}%=�= � =���<HG�<��<���<.�<��<�*�<���<�<k��<7��<�J�<m��<���<�G�<2��<#��<�</X�<̒�<Bʶ<���<W0�<t_�<S��<���<�ߟ<�<�,�<�P�<�s�<.��<���<�؄<���<H4z<�ur<۷j<�b<`?[<��S<e�K<�D<jd<<�4<-<(]%<Y�<�<Ax<0�<���; ��;�s�;!u�;ӄ�;¤�;֤;��;2q�;��q;��T;��7;
Y;���:���:y��:�J,:��y9y�9��J��z��;���\�hn�k�(�U�A�+�Z�.s�����R���񜻬^��q���j���lzɻ�Ի�޻�����ο��7�������0�9��s��`�U�"�"�&���*���.�Y�2���6��y:��9>���A�<�E�[$I��L��+P�?�S� W�dZ���]��a��Fd�.�g��j���m�q��!t��9w�wKz��W}��/�����\0�������(���������ˑ��<��z{����`���ё��A���������J��������d��RЛ�;��}���f��y��d⢼�K������}��m���4塚 X�������)������t���dd��Aͳ�@6��.���T���q��ۺ��D��⮽��  �  �N=��M=�IM=��L=e�K=�&K=�oJ=#�I=H I=HH=T�G=6�F=�F=�bE= �D= �C=�1C=`uB=��A=�@=�<@=�}?=!�>=l�==�;==y<=d�;=��:=�*:=�c9==�8=��7=�7=":6=:l5=��4=��3=��2=�#2=�L1=�s0=��/=ݺ.=��-=��,=�,=�(+=�<*=)M)=&Z(=|c'=�h&=vj%=�g$=�`#=)U"=�D!=�/ =�=�=,�=��=pv=L@==��=y=*=��=y=�=B�=P?=�=�N
=5�=�E=l�=d%=،=�� =~��<"G�<	��<���<�<���<�*�<���<�<���<L��<�J�<���<���<�G�<[��<H��<6�<ZX�<�<]ʶ<���<u0�<�_�<q��<��<�ߟ<��<t,�<�P�<�s�<��<���<�؄<Y��<�3z<�ur<��j<��b<�>[<�S<�K<`D<8d<<�4<�-<�\%<9�<�<�x<m�<A��;���;�t�;�u�;q��;���;�֤;\�;�q�;=�q;!�T;��7;YZ;���:H��:���:�O,:T�y9��9�N��|��P;��2^�!o���(���A�\�Z�&s�y���7S��C�k_��ޚ��ޣ���zɻԻ��޻?��A��y����6�C�����/���;�}`���"���&�u�*�|�.��2�k�6��y:��9>���A���E�'$I�íL��+P�`�S�oW�PdZ���]�$a� Gd���g�s�j���m�Vq�8"t��9w��Kz�QX}��/��3���e0������)��ˢ���������"��Y{��ql`��jё�gA��|������%��������d��-Л��:��Y���J���x��H⢼�K�������������^塚+X������)��ђ�������d��iͳ�Z6��V�������q��5ۺ��D�������  �   �N=��M=�IM=��L=]�K=�&K=�oJ=)�I=N I=	HH=\�G=F�F=�F=�bE=/�D=$�C=�1C=muB=��A=$�@=�<@=�}?=�>=h�==�;=="y<=o�;=��:=�*:=�c9=:�8=��7=�7=:6=)l5=��4=~�3=��2=�#2=�L1=�s0=��/=غ.=��-=��,=�,=�(+=�<*=%M)=*Z(=�c'=�h&=j%=�g$=�`#=6U"=�D!=�/ =�=�=4�=��=rv=J@==��=y=)*=��=�x=�=3�=K?=�=�N
=)�=�E=Y�=Z%=͌=�� =w��<G�<���<|��<�<��<�*�<���<�<���<S��<�J�<���<���<	H�<b��<f��<J�<mX�<��<mʶ<���<�0�<�_�<b��<��<�ߟ<��<�,�<�P�<�s�<���<���<�؄<B��<�3z<Qur<^�j<~�b<�>[<�S<��K<HD<�c<<׳4<�-<A]%<A�<|<vx<V�<v��;΁�;�t�;�u�;��;女;	פ;��;r�;1�q;
�T;s�7;�Z;0��:��:��:�N,:2�y96�9�K��|��5<��$`�Mo�I�(�k�A�ͩZ�As�	����S��m��_�����8����zɻBԻ��޻���f�򻤿���6�R��o���/�Ԫ��6`��"���&�=�*�i�.���2�B�6��y:�g9>���A��E�4$I�حL��+P� �S�\W�adZ��]�\a�Gd���g���j��m��q��"t�:w��Kz�zX}��/��R���u0������)������������.��R{��j]`��Wё�MA��]��������������d��Л��:��M���=���x��V⢼�K���������^���^塚8X��,����)��ݒ�������d���ͳ�z6��t�������q��Dۺ��D������  �  �N=��M=�IM=��L=e�K=�&K=�oJ=#�I=H I=HH=T�G=6�F=�F=�bE= �D= �C=�1C=`uB=��A=�@=�<@=�}?=!�>=l�==�;==y<=d�;=��:=�*:=�c9==�8=��7=�7=":6=:l5=��4=��3=��2=�#2=�L1=�s0=��/=ݺ.=��-=��,=�,=�(+=�<*=)M)=&Z(=|c'=�h&=vj%=�g$=�`#=)U"=�D!=�/ =�=�=,�=��=pv=M@==��=y=*=��=y=�=B�=P?=�=�N
=6�=�E=m�=f%=ٌ=�� =���<%G�<��<���<�<��<�*�<���<�<���<N��<�J�<���<���<�G�<[��<H��<5�<ZX�<�<\ʶ<���<s0�<�_�<n��<��<�ߟ<��<r,�<�P�<�s�<��<���<�؄<X��<�3z<�ur<��j<��b<�>[<�S<�K<cD<;d<<��4<�-< ]%<=�<�<�x<q�<I��;���;�t�;�u�;u��;���;�֤;[�;�q�;5�q;�T;��7;IZ;i��:��:}��:OO,:��y9h�9�~N��|���;��g^�<o���(���A�s�Z�<s�����AS��L�s_��嚳�䣾��zɻ Ի��޻C��D��|����6�D������/���<�}`���"���&�u�*�|�.��2�k�6��y:��9>���A���E�'$I�íL��+P�`�S�oW�PdZ���]�$a� Gd���g�s�j���m�Vq�8"t��9w��Kz�QX}��/��3���e0������)��ˢ���������"��Y{��ql`��jё�gA��|������%��������d��-Л��:��Y���J���x��H⢼�K�������������^塚+X������)��ђ�������d��iͳ�Z6��V�������q��5ۺ��D�������  �  
�N=��M=�IM=ǓL=a�K=�&K=�oJ=�I=: I=�GH=G�G=%�F=�F=�bE=�D=�C=r1C=QuB=��A=�@=�<@=�}?=�>=\�==�;==!y<=s�;=��:=�*:=�c9=K�8=��7=�7=7:6=Ll5=Ɯ4=��3=��2=�#2=�L1=�s0=��/=�.=��-=��,=�,=�(+=�<*=M)=Z(=kc'=�h&=ij%=�g$=�`#=U"=�D!=�/ =r=�=�=��=fv=?@==��=y=&*=��=y=�=W�=d?=;�=�N
=P�=�E=��=%=��=� =���<NG�< ��<���<4�<��<�*�<���<
�<o��<;��<�J�<q��<���<�G�<3��<$��<�<.X�<ʒ�<@ʶ<���<T0�<q_�<O��<���<�ߟ<��<�,�<�P�<�s�<*��<���<�؄<���<F4z<�ur<۷j<�b<b?[<��S<j�K<�D<qd<<�4<-<1]%<b�<�<Ix<9�<ǚ�;.��;t�;*u�;ڄ�;Ƥ�;	֤;��;.q�;|�q;�T;��7;�X;M��:N��:!��:J,:��y9��9��K��z���;��]뺚n���(���A�X�Z�Xs�'����R���񜻻^�����v���wzɻ�Ի�޻����Կ��!7������� 0�:��t��`�U�"�#�&���*���.�Z�2���6��y:��9>���A�<�E�[$I��L��+P�?�S� W�dZ���]��a��Fd�.�g��j���m�q��!t��9w�wKz��W}��/�����\0�������(���������ˑ��<��z{����`���ё��A���������J��������d��RЛ�;��}���f��y��d⢼�K������}��m���4塚 X�������)������t���dd��Aͳ�@6��.���T���q��ۺ��D��⮽��  �  �N=��M=�IM=œL=\�K=�&K=�oJ=�I= I=�GH="�G=�F=oF=cbE=�D=��C=P1C=*uB=e�A=��@=�<@=�}?=�>=a�==�;==$y<=v�;=��:=�*:=�c9=s�8=��7=�7=a:6=wl5=��4=��3=��2=�#2=M1=
t0=��/=��.=��-=��,=�,=�(+=�<*=M)=Z(=Pc'=�h&=Aj%=�g$=|`#=�T"=�D!=�/ =Y=��= �=��=Sv=1@==��=y=5*=��='y==y�=�?=]�=�N
=��=	F=��=�%=�=)� =
��<�G�<]��<҉�<F�<1��<�*�<���<	�<]��<��<�J�<6��<d��<�G�<ˑ�<���<��<�W�<���<�ɶ<]��<0�<N_�<-��<���<�ߟ<��<�,�<�P�<t�<Z��<���<ل<���<�4z<�vr<��j<��b<@[<�S<��K<LD<�d<<m�4<-<X]%<c�<�<ex<	�<Z��;I��;s�;�s�;���;v��;tԤ;_�;eo�;��q;�T;2�7;�V;��:���:F��:�I,:|y95 :��L�i{���9��[뺀l��(���A��Z��s������Q�����]��\��������yɻԻA�޻���d������"7�������0�����@a��"���&�]�*���.���2�K�6�{z:�F:>�S�A���E�b$I���L��+P��S�'W��cZ�:�]�wa�Fd�Àg���j���m�Zq�G!t�9w��Jz��W}�o/��㰁�.0��y����(���������ő��G���{����`���ё��A��바�=������L���Be���Л�c;���������-y���⢼�K���������^���6塚�W�������)��d���=���d���̳��5��ޞ����Kq���ں��D�������  �  F�N=��M=�IM=˓L=X�K=�&K=foJ=�I=��H=�GH=��G=��F=CF=3bE=��D=��C=(1C=�tB=?�A=��@=�<@=�}?=�>=U�==�;==+y<=��;=��:=�*:=�c9=��8=��7=�7=�:6=�l5='�4=��3=��2=$2=7M1="t0=Ә/=�.=��-=��,=�,=�(+=�<*=�L)=�Y(=2c'=�h&=j%=fg$=Q`#=�T"=�D!=V/ =0=��=��=n�=Av="@=�=��=#y=G*=��=Ly=)=��=�?=��=3O
=��=DF=�=�%=Z�=_� =e��<�G�<���<��<{�<R��<�*�<���<��<9��<���<XJ�<���<���<6G�<q��<���<S�<�W�< ��<�ɶ<#��<�/�<_�<�<׶�<�ߟ<��<�,�< Q�<]t�<���<3��<Vل<"��<�5z<9wr<��j<u�b<�@[<׆S<��K<�D<]e<<�4<�-<�]%<��<�<*x<��<���;E�;0r�;qr�;���;�;�Ҥ;��;�m�;��q;M�T;W�7;WT;i��:�~�:���:?D,:�oy9�:�uJ�+y���5���X��j���(�K�A���Z�ts�g���nP��A�\��C��������xɻ�Ի��޻s��g��1���y7�3��m��1�/�����a�Ν"���&��*�R�.�|�2��6��z:��:>���A�َE��$I��L��+P��S��W�wcZ���]�a��Ed��g�ʲj�>�m��q�� t�M8w�4Jz��V}�)/�������/��C����(������ ��ؑ������{���a��ґ�=B��9������쌗������e���Л��;������Zy���⢼�K������|��;���塚�W������S)����������c���̳�w5����������p��wں�JD��{����  �  S�N=��M=�IM=͓L=Y�K=�&K=[oJ=зI=��H=�GH=ɎG=��F=	F=�aE=x�D=o�C=�0C=�tB=�A=��@=�<@=�}?=�>=J�==�;==+y<=��;=��:=+:=
d9=��8=(�7=17=�:6=�l5=`�4=.�3=6�2=M$2=dM1=Ut0=�/='�.=��-=��,=�,=�(+=s<*=�L)=�Y(=c'=}h&=�i%=0g$=`#=�T"=CD!=#/ =�=��=��=C�=#v=@=�=��=0y=M*=�=ey=O=׮=�?=��={O
=��=�F=:�=1&=��=�� =ј�<OH�<���<W��<��<a��<�*�<���<��<��<���<�I�<���<���<�F�<���<���<��<
W�<���<4ɶ<���<{/�<�^�<Ћ�<���<�ߟ<��<�,�<.Q�<ut�<ߖ�<���<�ل<���<�6z<Ixr<u�j<��b<�A[<��S<��K<�D<f<<`�4<�-<�]%<��<�<�w<m�<���;~�;sp�;�p�;j��;���;�Ф;n�;�k�;��q;"�T;��7;eP;���:�y�:��:�>,:(iy9�:�I��w���4���S뺟h�
�(�{�A�O�Z���r��~���N��~휻B[����������xɻ3Ի�޻���O��i����7��������1�������b���"���&�$�*�1�.�k�2���6��{:�;>�:�A�.�E��$I�%�L��+P���S�yW�7cZ�R�]�La��Dd�@g�ٱj�F�m��q��t�a7w�\Iz�V}��.��P����/������(���������ꑊ�����{��6la��oґ��B������ ��s���&���f��Vћ�<��W���/���y���⢼�K������u��4�����W��C����(������x���@c��̳�5�����.���p��ں��C��(����  �  o�N=��M=�IM=ГL=O�K=v&K=GoJ=��I=��H=XGH=��G=d�F=�F=�aE=;�D=:�C=�0C=�tB=طA={�@=d<@=x}?=ֽ>=7�==�;==0y<=��;= �:=,+:=7d9=�8=^�7=g7=;6="m5=��4=n�3=l�2=�$2=�M1=�t0=�/=@�.=��-=��,=�,=�(+=e<*=�L)=�Y(=�b'=Ih&=�i%=�f$=�_#=MT"=D!=�. =�=Z�=��=,�=v=�?=�=��=7y=^*=5�=�y=�=�=6@=�=�O
=J�=�F=��={&=ߍ=�� =F��<�H�<T��<���<��<���<�*�<���<��<ӄ�<p��<�I�<4��<G��<CF�<���<���<h�<�V�<9��<�ȶ<Q��<</�<|^�<���<���<�ߟ<��<�,�<bQ�<�t�<9��<�< ڄ<	��<�7z<Tyr<��j<��b<�B[<��S<l�K<`D<�f<<�4<o-<^%<��<n<�w<�<S��;}�;o�;%o�;R~�;���;�Τ;F�;�i�;�q;�T;��7;�M;;��:�s�:ь�:*7,:Yy9�:��G��u���1��ZO�[f�3�(���A���Z�i�r��|���L���뜻�Y������F����vɻ�Իi�޻^��\�����8������J2�ۭ�j��c���"���&��*� �.�n�2���6��|:��;>���A���E�+%I�v�L��+P�֝S�(W��bZ���]��a�Dd�^~g��j�H�m�� q��t�m6w��Hz�$U}�x.������x/��묄��(���������������D|��}�a���ґ��B��4���z ��퍗������f���ћ��<������i���y��㢼�K��ƴ��p������bW��鿬��(��P�������b���˳��4���������p���ٺ��C��̭���  �  ��N=��M=JM=ٓL=K�K=i&K=+oJ=��I=��H=+GH=`�G=-�F=�F=�aE=��D=��C=t0C=YtB=��A=O�@=7<@=`}?=��>=,�==�;===y<=��;=�:=V+:=Td9=�8=��7=�7=F;6=Zm5=ݝ4=��3=��2=�$2=�M1=�t0=A�/=f�.=��-=��,=�,=�(+=T<*=�L)=�Y(=�b'=h&=�i%=�f$=�_#=T"=�C!=�. =�=%�=[�=�=�u=�?=�=��=Ay={*=K�=�y=�=8�=x@=Y�=P
=��=G=˹=�&=,�=%� =ə�<I�<���<��<!�<���<+�<���<��<���<%��<rI�<ڢ�<���<�E�<��<��<��<V�<Ȑ�<Uȶ<���<�.�<:^�<a��<m��<�ߟ<�<�,�<�Q�<�t�<z��<<��<�ڄ<���<�8z<7zr<��j<��b<�C[<��S<Z�K<D<kg<<��4<�-<m^%<߷<g<�w<��<a��;�{�;�m�;hm�;m|�;ě�;�̤;�;qg�;�q;��T;��7;J;V��:o�:*��:�1,:�Ly9�:�#F��s���-���L��c�V�(��A�j�Z�X�r�M{��CK��%ꜻX�����d����uɻzԻ�޻���]��Y���S8�v��=��3����P��d���"�~�&��*��.�D�2�y�6�[}:��<>�o�A� �E�z%I���L��+P���S��W�DbZ��]�"a�?Cd��}g��j�b�m���p��t�r5w��Gz�QT}�.������&/������j(��w��� ��(������v|���b��?ӑ�oC������� ��n������g��Cқ��<��������*z��6㢼L��д��d�������W������N(��㐯�����Ob��1˳�4�����<���o��Bٺ�@C�������  �  ��N= N=JM=דL=K�K=`&K=oJ=z�I=b�H=�FH=-�G=��F=TF=AaE=æD=��C=80C=#tB=w�A=�@=<@=S}?=��>=)�==�;==@y<=Ƶ;=(�:=w+:=~d9=R�8=��7=�7=;6=�m5= �4=��3=��2=�$2=�M1=�t0=c�/=~�.=��-=��,=�,=�(+=@<*=�L)=pY(=�b'=�g&=Li%=�f$=l_#=�S"=�C!=u. =S=��=5�=ԥ=�u=�?=�=��=Cy=�*=`�=�y=�=r�=�@=��=OP
=��=lG=�=
'=n�=X� =D��<�I�<��<&��<R�<Ϩ�<+�<���<��<���<���<I�<���<v��<cE�<���<���<g�<�U�<\��<�Ƕ<���<x.�<^�<1��<M��<�ߟ<��< -�<�Q�<2u�<���<���<�ڄ<���<�9z<.{r<��j<� c<�D[<|�S<"�K<�D<h<<&�4<	-<�^%<�<j<kw<V�<��;#z�;�k�;�k�;�z�;ř�;bʤ;�;,e�;ʣq;��T;J�7;YF;q��:/l�:˃�:�.,:�>y9!:��D�s���*���H�a�<�(�M�A�B�Z���r�dy���I��d蜻�V������윾��tɻ�Իߎ޻��軝��Z����8��������3�N��+��e���"�o�&��*��.�0�2�S�6�	~:�|=>���A�b�E��%I���L��+P�m�S��W��aZ���]�a a�|Bd��|g��j���m���p��t��4w��Fz��S}��-��e����.������M(��p�����(������|�����lb���ӑ��C�����x!��ߎ������wg���қ�P=��h���!��Mz��a㢼,L��д��k��߅��q�V��b����'������=����a���ʳ��3���������Bo���غ��B��E����  �  εN= N=)JM=ۓL=C�K=M&K=�nJ=S�I=G�H=�FH=�G=��F=%F=aE=��D=��C=	0C=�sB=O�A=�@=�;@=,}?=��>=�==�;==Ey<=ص;=B�:=�+:=�d9=m�8=��7=7=�;6=�m5=L�4=�3=�2=%2=N1=�t0=|�/=��.=�-=��,=�,=�(+=/<*=�L)=NY(=wb'=�g&="i%=Yf$=A_#=�S"=iC!=M. =$=��=�=��=�u=�?=�=��=Hy=�*=��=�y=�=��=�@=��=�P
=
�=�G=P�=?'=��=�� =���<�I�<U��<d��<��<��<+�<���<e�<a��<���<�H�<;��<#��<E�<I��<.��<�<8U�<���<�Ƕ<Q��<A.�<�]�<���<$��<tߟ<��<-�<�Q�<^u�<���<Ṉ<Dۄ<H��<H:z<�{r<d�j<Kc<�E[<[�S<��K<wD<�h<<��4<~	-<�^%<��<R<"w<��<���;?y�;k�;Mj�;	y�; ��;�Ȥ;K�;�c�;b�q;��T;T�7;KD;��:Kf�:)��:n(,:�0y9�:�CB��p��)��eE��_���(���A���Z�&�r�&x��UH��D眻gU������#���Atɻ1Ի�޻y�軫������8�<��1��<4�߯���of�Q�"�5�&���*���.���2��6��~:��=>�Y�A�ԐE�%&I���L��+P�X�S�_W��aZ�;�]���`�Bd�|g�l�j���m��p��t��3w��Ez��R}�s-��%����.��a���'(��f�����E���<���|��M����b���ӑ�0D��z����!��@��������g��ӛ��=������U���z���㢼QL��ݴ��c��ą��9�V��(����'��6��������a��^ʳ�+3��G���q���n���غ��B������  �  ۵N=) N=#JM=��L=D�K=G&K=�nJ=>�I=/�H=�FH=�G=��F=�F=�`E=_�D=g�C=�/C=�sB=+�A=��@=�;@=}?=��>=�==�;==Iy<=ӵ;=Q�:=�+:=�d9=��8=�7=)7=�;6=�m5=r�4=A�3=/�2=C%2=?N1=u0=��/=��.=�-=��,=�,=�(+=.<*=xL)=7Y(=^b'=�g&=i%=:f$=_#=S"=;C!=&. ==��=��=��=�u=�?=�=��=Vy=�*=��=	z==��=A=��=�P
=E�=�G=��=v'=ʎ=�� =ښ�<J�<���<���<��<���<2+�<w��<t�<L��<���<�H�<��<���<�D�<���<���<��<�T�<���<QǶ< ��<.�<�]�<�<��<nߟ<�<
-�<�Q�<xu�<4��<��<�ۄ<���<�:z<�|r<��j<c<;F[<�S<y�K<�D<i<<ɷ4<�	-<�^%<�<Y<w<��<���;vx�;�i�;5i�;x�;���;wǤ;�
�;:b�;��q;r�T;��7;�A;��:{c�:��:�$,:�1y9�:��D��o���'���B�%^�X�(���A�k�Z���r�w���F��n朻@T��ɐ��I����sɻ�Ի �޻���������9�c������4����U��f���"���&���*�i�.��2�o�6�A:�G>>���A��E�$&I�ܮL��+P�S�S�VW�TaZ�ٴ]�w�`��Ad�u{g���j��m�l�p�Pt�+3w��Ez�FR}�5-����.��?���-(��_�����X���6���|�������b��6ԑ�hD��Ƴ��"������?���(h��Gӛ��=����������z���㢼ZL��ᴥ�Y��х��(�V��񾬼r'����������Aa���ɳ��2��蛶�&���n��Hغ�gB��Ь���  �  �N=7 N=3JM=�L=<�K=<&K=�nJ=:�I=#�H=�FH=ύG=��F=�F=�`E=R�D=S�C=�/C=�sB=�A=��@=�;@=}?=|�>=�==�;==Oy<=�;=`�:=�+:=�d9=��8=!�7=<7=�;6=n5=��4=V�3=G�2=Q%2=NN1="u0=��/=��.=,�-=��,=�,=�(+=<*=iL)=2Y(=Ob'=�g&=�h%=#f$=_#=pS"=-C!=. =�=��=��=��=�u=�?=�=��=Ty=�*=��=z=*=ү=A=�=�P
=]�=�G=��=�'=�=�� =��<AJ�<���<���<��<��<(+�<i��<O�<=��<~��<�H�<ա�<���<�D�<Ύ�<���<��<�T�<���<%Ƕ<���<�-�<�]�<̊�<���<^ߟ<�<+-�<�Q�<�u�<N��<B��<�ۄ<���<>;z<}r<O�j<kc<�F[<:�S<��K<CD<Pi<<�4<�	-<#_%< �<9<�v<��<Փ�;x�;Bi�;�h�;'w�;�;�Ƥ;
�;�a�;ݛq;��T;\�7;�@;U��:<b�:�|�:g!,:G&y9U:��A�n�� &��A�7]���(���A�6�Z���r��v��4F���圻�S��[���Ú��*sɻPԻ��޻/�軗��7���T9��������4�°���Sg�J�"�,�&���*���.���2�Ͱ6�~:��>>���A�;�E�r&I���L��+P�"�S�%W�aZ���]�/�`�BAd�<{g���j���m�%�p�
t��2w�3Ez�R}�-��ͮ��u.�����(��N�����k���_��}�������b��Uԑ��D������E"������d���Sh��yӛ�>���������z���㢼vL��𴥼V������lV��ؾ��O'��Տ��i���a���ɳ��2���������tn��.غ�CB�������  �  Z�N=vN=bQM=�L=(�K=0K=�yJ=��I=�I=TH=/�G=��F=c+F=arE=��D=:�C=
EC=K�B=�A=0A=�V@=u�?=p�>=�>=�\==0�<=p�;=�;=�S:=��9=p�8=� 8=�77=�m6=�5=��4=�4=�43=1b2=��1=�0=��/=x/=i$.=�C-='`,=�y+=Ï*=��)=�(=��'=��&=U�%=�$=c�#=6�"=O�!={� =��=Ke=�B==��=9�=�|=y;=��=¥=�P=p�=;�=T*=к=�D=,�
=7E	=�=�,=��=��=.\=�l�<G�<��<	L�<���<�\�<���<_L�<u��<��<�{�<I��<�&�<�s�<��<r��<�>�<1z�<��<��<�<�F�<�r�<���<"ħ<��<I�<I/�<�O�<�n�<��<5��<�ƈ<y�<���<�2z<�ir<��j<��b<5[<�LS<x�K<1�C<	<<�L4<,�,<E�$<�*<>|<`�<-<�;���;��;<��;1��;"��;_��;��;!�;Y�l;ƾO;+�2;��;���:j�:�ρ::��9x��,|4��⏺��ĺ'Y��&��R0��OI��'b���z�F\��J7��qߠ�
U��Ö��̤»�~ͻ%ػ,�⻠�� ���M^ �Q2���	�R��)�֑�H��k8 ��k$�P�(��,�ތ0�,r4�}F8��	<�ٽ?��bC���F���J�� N��rQ���T��5X���[���^�Fb�]Ie��yh�u�k�h�n�x�q���t��x�b{�$~���������������:u���뇼�a���Պ��H������a+������	���w��Q䔼TP��b����%���������,`���Ǟ�,/���������Nc���ɥ�>0������C����c��`ʬ�1��엯������e���̳�4��l�������j���Һ��:�������  �  L�N=~N=bQM=�L=-�K=0K=�yJ=��I=�I=%TH=>�G=�F=c+F=qrE=�D=J�C=	EC=T�B=�A=:A=�V@=z�?=r�>=�>=�\==.�<=t�;=�;=�S:=��9=c�8=� 8=�77=�m6=ء5=��4=�4=�43=-b2=��1=ֶ0=��/=j/=r$.=�C-=)`,=�y+=ď*=��)=��(=��'=��&=b�%=�$=k�#=B�"=Z�!=�� =��=Ve=�B==��=?�=�|=u;=��=��=�P=b�=$�=I*=ĺ=�D=�
=.E	=�=�,=��=��=&\=sl�<+�<׵�<�K�<���<�\�<���<KL�<t��<��<|�<]��<�&�<�s�<���<���<�>�<Pz�<��<��<%�<�F�<�r�<���<(ħ<��<R�<N/�<�O�<�n�<��<��<�ƈ<j�<���<�2z<lir<��j<��b<[<�LS<U�K<��C<�<<�L4<H�,<?�$<�*<M|<O�<-<��;���;O��;���;\��;)��;踢;�;�!�;a�l;t�O;�2;_�;#��:\�:OЁ:X:$�99��`z4��ᏺ��ĺ8Z��Ώ��0�>PI�(b�D�z��\��r7���ߠ�!U������»�ͻz%ػ֗⻺�����I^ �H2���	� ���������r8 ��k$��(��,���0�3r4�NF8��	<���?��bC���F���J�� N��rQ��T�^5X�Ӈ[�!�^�kb��Ie��yh���k���n���q���t��x��{�:~�������ւ������-u��쇼�a���Պ��H��~���D+�������	��{w��T䔼6P��E���}%��
�������`���Ǟ�/���������Sc���ɥ�;0������.����c��~ʬ�'1�����������e���̳�/4��}�������j���Һ��:�������  �  >�N=sN=PQM=�L=5�K=0K=�yJ=��I=�I=5TH=Z�G="�F=�+F=�rE=)�D=o�C=(EC=u�B=(�A=JA=�V@=��?=��>=�>=�\==$�<=e�;=�;=�S:=��9=H�8=� 8=�77=m6=��5=^�4=j4=�43=b2=u�1=Ƕ0=��/=]/=i$.=�C-=.`,=�y+=Ώ*=��)=	�(=��'=��&=��%=1�$=��#=`�"=u�!=�� =��=we=�B=*=��=E�=�|=u;=��=��=�P=O�=�=9*=��=�D=��
=
E	=ۻ=�,=t�=��=\=.l�<�<���<�K�<���<�\�<���<NL�<���<��<)|�<y��<�&�<"t�<7��<���<?�<�z�<`��<��<f�<G�<#s�<ɜ�<Nħ<��<c�<N/�<�O�<�n�<錐<��<eƈ<.�<���<2z<�hr<�j<M�b<�[<HLS<ՈK<��C<�<<EL4<�,<��$<�*<i|<n�<Y-<��;!��;ѿ�;���;n��;O��;��;�;�"�;��l;��O;��2;��;���:o�:�Ӂ:�:��9����|4��⏺K�ĺBZ��.��0�5RI��)b��z��]��58���࠻�U��՗��u�»�ͻ�%ػ��4������2^ �2���	�����n������7 ��j$���(�r�,��0��q4��E8��	<�]�?��bC���F�[�J�� N�wrQ�M�T��5X��[�8�^��b��Ie�0zh�8�k���n�G�q�B�t�\x�#{��~�Q�����肃�����Eu��쇼xa���Պ��H��k���(+��Ԛ���	��9w��䔼�O�����:%��Î�������_���Ǟ��.��액�����@c���ɥ�?0��ʖ��C����c���ʬ�S1��7������'f��2ͳ�w4������C���j���Һ�.;��ɣ���  �  (�N=]N=OQM=�L=3�K='0K=�yJ=��I=�I=bTH=��G=L�F=�+F=�rE=c�D=��C=\EC=��B=R�A=wA=�V@=��?=��>=�>=�\==$�<=_�;=�;=�S:=u�9= �8=� 8=�77=Om6=��5=0�4=44=z43=�a2=L�1=��0=��/=G/=V$.=�C-=-`,=�y+=ݏ*=Ƣ)=)�(=�'=��&=��%=_�$=��#=��"=��!=֚ =�=�e=�B=N=��=Z�=�|=r;=��=��=�P=2�=�=�)=n�=YD=��
=�D	=��=a,=8�=J�=�[=�k�<��<n��<�K�<���<�\�<}��<ML�<���<��<d|�<���<A'�<pt�<���<4 �<�?�<�z�<Ų�<F�<��<eG�<ps�<��<~ħ<��<f�<R/�<�O�<�n�<���<ũ�<ƈ<��<X��<N1z<hr<T�j<j�b<�[<�KS<+�K<��C<�<<�K4<��,<��$<�*<U|<��<�-<��;E��;L��;��;��;��;ǻ�;	�;�$�;k�l;��O;�2; ;d��::�:�ց:�:��9��|4��䏺n�ĺ_��1���0�kTI�g,b�ޥz�_���9���ᠻW������Ѧ»�ͻ_&ػ���������$^ ��1��	�c����������27 �?j$���(���,�Y�0��p4�E8��<���?��aC�#�F� �J�� N�|rQ�N�T��5X�[�[���^�Ub��Je��zh��k���n��q��t�!x��{�C~�����a��������Xu��쇼�a���Պ�rH��5����*��~���8	���v���㔼�O�������$��a���=����_��AǞ��.������{���(c���ɥ�@0��ʖ��m���d���ʬ��1������u����f���ͳ��4��&������Lk��7Ӻ��;������  �  �N=CN=AQM=�L=;�K=;0K=�yJ=$�I=I=�TH=��G=��F=�+F=sE=��D=��C=�EC=ߊB=��A=�A=
W@=ř?=��>=�>=�\==�<=N�;=l;=vS:=I�9=��8=R 8=^77=m6=@�5=��4=�4=<43=�a2=�1=n�0=�/=*/=@$.=�C-=%`,=�y+=��*=�)=M�(=	�'=��&=��%=��$=��#=ӻ"=�!=� ='�=�e= C=n=��=r�=�|={;=��=��=�P=�==�)=7�=D=p�
=zD	=S�=,=�=��=�[=Zk�<)�<��<IK�<T��<�\�<n��<`L�<���<�<�|�<��<�'�<�t�<(��<� �<@�<z{�<O��<��<2�<�G�<�s�<b��<�ħ<�<��<G/�<�O�<�n�<���<q��<�ň<t�<���<M0z<�fr<I�j<E�b<�[<jJS<4�K<�C<8<<RK4<,�,<��$<m*<k|<��<�-<�;d��;���;��;$��;a��;���;��;�&�;c�l;��O;r�2;z;g��:G"�:cځ:�:D9!���}4��揺��ĺPc��0��V#0��WI�0b���z��`���;���㠻Y��D�����»��ͻ%'ػ��U�������] �x1���	�Ə�i�؏����6 �4i$���(�}�,�V�0��o4�/D8��<�"�?�daC���F�΂J�{ N��rQ�v�T�6X�̈[�C�^��b�IKe��{h�ߤk���n��q��t�1x��{�G~�􉀼���`���J���~u��0쇼{a��rՊ�PH����*��.������kv�� 㔼O�����W$��ڍ������_���ƞ�W.��a���N��� c���ɥ�Q0��疨�����Kd��(ˬ��1��혯������f��&γ�M5���������k���Ӻ��;��t����  �  ߺN=(N=.QM=�L=B�K=G0K=�yJ=K�I=7I=�TH=��G=��F=G,F=SsE=��D=- D=�EC= �B=��A=�A=?W@=�?=��>=�>=�\==�<=:�;=O;=JS:=�9=��8= 8=77=�l6=�5=��4=�4=�33=ca2=ی1=5�0=T�/=/=+$.=�C-=)`,=�y+= �*=��)=|�(=C�'=7�&=#�%=��$=I�#=�"=4�!=`� =c�=f=:C=�=&�=��=�|=|;=��=u�=�P=��=��=�)=�=�C=�
=D	=�=�+=��=��=2[=�j�<��<���<�J�<��<c\�<b��<ZL�<Ը�<E�<�|�<q��<$(�<`u�<���<Q�<�@�<|�<볾<]�<��<KH�<4t�<���<�ħ</�<��<P/�<�O�<hn�<4��<��<@ň<���<G��</z<�er<�j<��b<g[<MIS<�K< �C<x<<�J4<��,<3�$<V*<||<��<o.<[�;'��;���;$��;a��;�;���; �;�)�;��l;~�O;8�2;�;���:�(�:�߁:S#:�!9���.4��菺��ĺ�g������&0�l[I�*4b��z�c���=���堻�Z��)�����»��ͻ4(ػ��⻭�컬����] �*1��	����s�َ����5 ��g$���(�H�,��0��n4�$C8��<�5�?��`C��F�}�J�T N�xrQ���T�g6X�]�[���^��b�XLe��|h���k��n�G�q�J�t�Zx��{�K~�x��������������u��E쇼oa��cՊ�H������0*������D���u���┼mN��{����#��B���0����^��hƞ��-���������b���ɥ�N0����������d��{ˬ�u2��r���} ���g���γ��5��H������Ql��-Ժ�Q<��Ǥ���  �  ��N=N=QM=ޛL=J�K=\0K=zJ=k�I=oI=UH=G�G=�F=�,F=�sE=J�D=� D=4FC=m�B=�A=A=rW@=�?=��>=�>=�\==�<=%�;=1;=S:=�9=s�8=��7=�67=nl6=��5=H�4=S4=�33=a2=��1=��0=#�/=�/=$.=�C-=(`,=�y+=�*="�)=��(=w�'=o�&=m�%=-�$=��#=s�"=��!=�� =��=Wf=pC=�=J�=��=�|={;=��=Z�=^P=��=L�==)=��=cC=��
=�C	=��=Q+=(�=F�=�Z=j�<�<��<�J�<���<9\�<P��<\L�<��<p�<N}�<���<�(�<�u�<;��<��<SA�<�|�<���<��<Z�<�H�<�t�<	��<Hŧ<g�<��<P/�<_O�<>n�<܋�<���<�Ĉ<c��<���<�-z<adr<u�j<��b<�[<�GS<�K<��C<�<<�I4<8�,<��$<7*<�|<K�<�.<g�;���;���;���;���;���;�â;#�;�,�;��l;�O;d�2;W;���:-.�:��:�*:�49M���4��ꏺ��ĺ�l����^*0��_I��8b�q�z��e��@��N蠻�\�����C�»!�ͻI)ػ?��$�컈���v] ��0�|�	�Q����������3 ��f$��(��,�Ǉ0��m4��A8��<�^�?��_C���F��J�/ N�qrQ���T��6X��[���^��b�`Me�	~h�S�k�M�n���q���t��x�#{�^~����������������u��U쇼ia��JՊ��G��j����)��L������Nu��┼�M��и��#�����������]���Ş�z-��ʔ�������b���ɥ�T0��2��������d���ˬ��2��������=h��\ϳ��6��坶�\���l���Ժ��<��/����  �  ��N=�N=QM=֛L=O�K=q0K=3zJ=��I=�I=EUH=��G=m�F=�,F=�sE=��D=� D=�FC=��B=T�A=PA=�W@=4�?=��>=�>=�\==�<=�;=;=�R:=��9=:�8=��7=~67=l6=L�5=��4=4=T33=�`2=X�1=µ0=��/=�/=�#.=yC-=%`,=�y+=/�*=A�)=в(=��'=��&=��%=��$=��#=��"=ٮ!=�� =��=�f=�C==q�=��=�|=�;=��=E�=5P=|�=�=�(=H�=C=\�
=\C	=&�=�*=Ǖ=��=�Z={i�<��<���<.J�<z��<\�<:��<nL�< ��<��<�}�<C��<)�<�v�<��<��<B�<j}�<7��<��<��<OI�<u�<t��<�ŧ<��<��<I/�<CO�<�m�<���<N��<LĈ<�߄<
��<m,z<�br<�j<8�b<�[<�FS<��K<��C<�<<"I4<��,<l�$<*<�|<��<[/<� �;���;���;İ�;���;��;~Ƣ;*�;�/�;m;��O;Z�2;�;��:t5�:��:+3:E9�
��(�4��폺Z�ĺKr����f.0�dI�1=b�S�z�h��mB��W꠻$_������լ»q�ͻ*ػ��_�����@] �L0���	������Ќ����q2 �Ze$�Ƀ(���,�z�0�8l4��@8��<�y�?�/_C�	�F���J���M�wrQ��T�97X�q�[�b�^��b�UNe�<h�t�k���n���q���t��	x�S{��~�s������c������v��f쇼ha��#Պ��G�����l)��Ԙ��;���t��Wᔼ)M��"���m"����������q]��sŞ�-��h��������b��ɥ�`0��T���E���9e��J̬�f3����������h��	г�P7����������m��?պ�C=�������  �  k�N=�N=�PM=ϛL=S�K=�0K=NzJ=��I=�I=�UH=̝G=��F=4-F=EtE=��D=D=�FC=��B=��A=�A=�W@=^�?=�>=�>=�\==��<= �;=�;=�R:=v�9=��8=>�7==67=�k6=��5=��4=�4=33=�`2=�1=��0=��/=�/=�#.=pC-=`,=�y+=C�*=a�)=��(=޾'=��&=��%=��$=/�#=�"=%�!=B� =;�=�f=�C=4=��=ݷ=�|=�;=��=2�=P=O�=ӑ=�(=��=�B=�
=�B	=˹=�*=j�=��=.Z=�h�<��<:��<�I�<D��<�[�<��<{L�<8��<��<�}�<���<�)�<�v�<r��<*�<�B�<~�<ѵ�<)�<p�<�I�<}u�<ў�<�ŧ<��<��<A/�<5O�<�m�<W��<㧌<�È<O߄<���<?+z<�ar<טj<��b<m
[<�ES<��K<��C<�<<tH4<�,<1�$<�)<�|<��<�/<N"�;��;���;��;��;��;)ɢ;��;92�;�m;S�O;E�2;o;���:U<�:�:�::XO9���E�4�����ź#x����20��gI�}Ab�лz�%j���D��G젻�`������y�»�ͻ+ػ��⻀�컔���] ��/�c�	�Ό���������_1 �+d$���(�L�,�I�0�"k4��?8��<���?�y^C�y�F�Z�J���M��rQ�4�T��7X���[�,�^��b�UOe�@�h�{�k���n�'�q�%�t�x�Z{��~�틀�h	����K���$v��z쇼oa��Պ�G��ȸ��)��b������=t�������L��}����!��h���t����\���Ğ��,�����X���fb��qɥ�n0��e��������e���̬��3�����/��di���г��7��4������	n���պ��=��	����  �  F�N=�N=�PM=țL=\�K=�0K=hzJ=��I=�I=�UH=�G=��F=s-F=�tE=2�D=bD=GC=;�B=��A=�A=�W@=z�?=-�>=>=�\==�<=��;=�;=�R:=S�9=��8=�7=�57=�k6=��5=`�4=p4=�23=O`2=ދ1=a�0=��/=v/=�#.=^C-=`,=�y+=V�*=|�)=�(=�'=�&=0�%=��$=q�#=L�"=c�!=�� =v�=g=D=Y=��=�=�|=�;=��=�=�O=%�=��=�(=��=pB=��
=�B	=z�==*=�=E�=�Y=bh�<��<ز�<�I�<��<�[�<��<�L�<V��<�<0~�<���<�)�<w�<��<��<#C�<�~�<V��<��<��<0J�<�u�<��<Ƨ<��<��<7/�<O�<�m�<��<���<�È<�ބ<���<*z<�`r<��j<��b<G	[<tDS<��K<�C<<<�G4<��,<��$<�)<�|<�<20<?#�;|��;O��;���;��;?��;�ˢ;H��;�4�;�m;4�O;"�2;�;]�:5A�:��:�@:b9�	���4���ź\{�����:50��kI�BEb�t�z�/l���F��c�b��_�����»��ͻ,ػ4����컁����\ ��/���	�;��%���s��[0 �c$�~�(�E�,�7�0�$j4��>8�3<��?��]C��F��J���M�rQ�v�T��7X�v�[���^�b�3Pe�.�h���k���n�7�q�(�t�%x�v{��~�V����	���������Nv���쇼_a���Ԋ�RG�������(�����W���s��H���L�����J!��抚���q\���Ğ�^,��Փ��#���Gb��]ɥ�|0�����������e���̬�-4��y�������i��'ѳ�p8���������n��;ֺ�>��N����  �  '�N=�N=�PM=˛L=\�K=�0K=zJ=��I=%I=�UH=,�G=�F=�-F=�tE=_�D=�D=>GC=h�B=��A=�A=X@=��?=B�>=>=�\==�<=��;=�;=�R:=/�9=��8=��7=�57=_k6=��5='�4=C4=�23=%`2=��1=7�0=w�/=[/=�#.=WC-= `,=�y+=a�*=��)=8�(=8�'=B�&=W�%='�$=��#={�"=��!=�� =��=:g=6D=�=��=�=�|=�;=��=�=�O=�=y�=O(=��=>B={�
=zB	=8�=�)=�=�=�Y=�g�<B�<���<II�<���<�[�<��<uL�<u��<?�<m~�<L��<9*�<�w�<@��<�<�C�<�~�<���<�<>�<�J�<:v�<H��<7Ƨ<��<��<C/�<O�<~m�<Ԋ�<U��<$È<}ބ<���<A)z<�_r<��j<�b<j[<�CS<�K<Z�C<r<<GG4<S�,<��$<�)<�|<�<�0<$�;���;���;B��;���;ڴ�;[͢;���;�6�;'m;}�O;�2;;�:E�:4��:�B:&j9�����4���7
ź$��%��;70�nI��Gb�W�z��m���G����c������Ȱ»��ͻ�,ػ�����U����\ �a/���	�ǋ�]�h������/ �Ib$���(���,�e�0�ti4�>8��<�,�?�r]C���F�ŀJ���M�vrQ���T�8X�ދ[�J�^��b��Pe�сh�i�k���n��q���t��x�1{�~������	��L�������kv���쇼_a���Ԋ�*G��e����(��������Ys���ߔ��K������� ��������&\��NĞ�,����������<b��]ɥ�r0����������f��Aͬ��4��͛����Xj���ѳ��8�����z���n���ֺ�l>�������  �  �N=�N=�PM=L=b�K=�0K=�zJ=�I=*I=�UH=H�G=<�F=�-F=�tE=��D=�D=aGC=��B=�A=�A= X@=��?=K�>=>=�\==�<=��;=�;=yR:=�9=��8=��7=�57=:k6=i�5=�4=4=u23=`2=��1=%�0=j�/=R/=�#.=QC-=`,=�y+=k�*=��)=?�(=?�'=]�&=p�%=M�$=��#=��"=��!=М ==Qg=QD=�=��=�=�|=�;=��=�=�O=��=h�=8(=j�=B=W�
=LB	=�=�)=��=��=�Y=�g�<�<d��<'I�<���<�[�<��<�L�<���<U�<o~�<i��<r*�<x�<���<R�<�C�<;�<���<N�<x�<�J�<Gv�<a��<OƧ<�<�<0/�<�N�<Wm�<���<1��<È<Kބ<_��<�(z<;_r<?�j<q�b<�[<2CS<q�K<�C<<<G4<�,<��$<�)<�|<d�<�0<p$�;"��;���;6��;���;��;u΢;"��;�7�;�m;��O;2�2;�;	�:>G�:���:QH:o9J���4�<���`źq���	��90��oI�Jb�4�z��n��I�����d��<���E�»T�ͻ-ػ��?�컟����\ �2/�V�	����<����c��/ ��a$�,�(��,��0��h4��=8�<��?�V]C�}�F���J�[�M��rQ���T�O8X��[�|�^�b�2Qe�\�h��k�#�n���q�y�t�zx��{��~�ӌ��#
��e�������v���쇼ca���Ԋ�G��J���}(���������&s���ߔ�dK��^���� ��E���W��[��Ğ��+����������b��Mɥ��0����������f��cͬ��4������G���j���ѳ�9��W������"o���ֺ��>�������  �  �N=�N=�PM=��L=d�K=�0K=�zJ=�I=6I=�UH=O�G=C�F=�-F=�tE=��D=�D=lGC=��B=�A=A=1X@=��?=A�>=>=�\==�<=��;=�;=rR:=�9=��8=��7=�57=6k6=[�5= �4=4=w23=�_2=��1=�0=\�/=M/=�#.=XC-=`,=�y+=d�*=��)=T�(=I�'=h�&=t�%=W�$=��#=��"=¯!=՜ =̈́=Tg=ZD=�=��=�=�|=�;=��=�=�O=��=X�=+(=a�=	B=X�
=?B	=	�=�)=��=��=�Y=�g�<��<N��<I�<���<�[�<���<�L�<j��<r�<�~�<���<�*�<x�<���<a�<�C�<T�<��<_�<��<�J�<]v�<���<DƧ<�<�<"/�<�N�<Tm�<���<��<�<0ބ<O��<�(z<�^r<��j<.�b<�[<CS<5�K<�C<�<<G4<��,<��$<~)<�|<a�<�0<�$�;���;���;w��;���;E��;�΢;���;�7�;Ym;��O;��2;�;@�:%I�:���:�H:n9���k�4�d���ź#���d���90��oI�XJb��z��n��uI����9e��������»ͻ1-ػ!���컾����\ �P/�E�	�O���ɉ�N���. ��a$��(���,�Ղ0��h4��=8��<��?� ]C�U�F�ĀJ�F�M��rQ���T�V8X��[���^�2b�NQe���h�٫k�T�n���q���t��x��{��~�ߌ��=
��y��������v���쇼ga���Ԋ�.G��,���V(��x������s���ߔ�VK��9���� ��7���F��[�� Ğ��+��i�������"b��Hɥ��0����������%f���ͬ��4�����U���j���ѳ�:9��x������.o���ֺ��>��ݦ���  �  �N=�N=�PM=L=b�K=�0K=�zJ=�I=*I=�UH=H�G=<�F=�-F=�tE=��D=�D=aGC=��B=�A=�A= X@=��?=K�>=>=�\==�<=��;=�;=yR:=�9=��8=��7=�57=:k6=i�5=�4=4=u23=`2=��1=%�0=j�/=R/=�#.=QC-=`,=�y+=k�*=��)=?�(=?�'=]�&=p�%=M�$=��#=��"=��!=М ==Qg=QD=�=��=�=�|=�;=��=�=�O=��=i�=9(=j�=B=X�
=NB	=�=�)=��=��=�Y=�g�<�<h��<+I�<���<�[�<��<�L�<���<X�<r~�<l��<t*�<x�<���<S�<�C�<;�<���<M�<w�<�J�<Ev�<_��<LƧ<�<�<-/�<�N�<Tm�<���</��<È<Jބ<^��<�(z<:_r<?�j<r�b<�[<5CS<t�K<�C<$<<G4<�,<��$<�)<�|<j�<�0<z$�;+��;���;=��;���;��;u΢;!��;�7�;�m;~�O; �2;�;��:G�:���:�G:�l9a��y�4������ź����+��=90�pI�3Jb�P�z��n��I�����d��E���M�»[�ͻ-ػ��D�컣����\ �4/�W�	����=����d��/ ��a$�,�(��,��0��h4��=8�<��?�V]C�}�F���J�[�M��rQ���T�O8X��[�|�^�b�2Qe�\�h��k�#�n���q�y�t�zx��{��~�ӌ��#
��e�������v���쇼ca���Ԋ�G��J���}(���������&s���ߔ�dK��^���� ��E���W��[��Ğ��+����������b��Mɥ��0����������f��cͬ��4������G���j���ѳ�9��W������"o���ֺ��>�������  �  '�N=�N=�PM=˛L=\�K=�0K=zJ=��I=%I=�UH=,�G=�F=�-F=�tE=_�D=�D=>GC=h�B=��A=�A=X@=��?=B�>=>=�\==�<=��;=�;=�R:=/�9=��8=��7=�57=_k6=��5='�4=C4=�23=%`2=��1=7�0=w�/=[/=�#.=WC-= `,=�y+=a�*=��)=8�(=8�'=B�&=W�%='�$=��#={�"=��!=�� =��=:g=6D=�=��=�=�|=�;=��=�=�O=�={�=Q(=��=@B=}�
=|B	=;�=*=�=�=�Y=�g�<J�<���<QI�<���<�[�<��<|L�<{��<E�<r~�<Q��<=*�<�w�<B��<�<�C�<�~�<���<�<;�<�J�<5v�<C��<1Ƨ<��<��<=/�<�N�<ym�<ϊ�<Q��< È<zބ<���<>)z<�_r<��j<	�b<m[<�CS<�K<b�C<{<<RG4<^�,<��$<�)<�|<*�<�0<$�;���;���;O��;���;ߴ�;\͢;���;�6�;m;b�O;��2;�;��:�D�:���:�A:f9�����4�P��
ź���g��{70�XnI�/Hb���z��m���G����c������ذ»�ͻ�,ػ���%��]����\ �d/���	�ɋ�^�j������/ �Jb$���(���,�f�0�ui4�>8��<�,�?�r]C���F�ŀJ���M�vrQ���T�8X�ߋ[�J�^��b��Pe�сh�i�k���n��q���t��x�1{�~������	��L�������kv���쇼_a���Ԋ�*G��e����(��������Ys���ߔ��K������� ��������&\��NĞ�,����������<b��]ɥ�r0����������f��Aͬ��4��͛����Xj���ѳ��8�����z���n���ֺ�l>�������  �  F�N=�N=�PM=țL=\�K=�0K=hzJ=��I=�I=�UH=�G=��F=s-F=�tE=2�D=bD=GC=;�B=��A=�A=�W@=z�?=-�>=>=�\==�<=��;=�;=�R:=S�9=��8=�7=�57=�k6=��5=`�4=p4=�23=O`2=ދ1=a�0=��/=v/=�#.=^C-=`,=�y+=V�*=|�)=�(=�'=�&=0�%=��$=q�#=L�"=c�!=�� =v�=g=D=Z=��=�=�|=�;=��=�=�O='�=��=�(=��=sB=��
=�B	=~�=A*=�=I�=�Y=lh�<��<��<�I�<��<�[�<%��<�L�<`��<'�<8~�<���<�)�<�w�<��<��<$C�<�~�<T��<��<��<+J�<�u�<��<�ŧ<��<��<//�<O�<�m�<��<���<zÈ<�ބ<���<*z<�`r<��j<��b<L	[<|DS<��K<(�C<<<�G4<��,<��$<�)<�|<(�<A0<\#�;���;e��;��;"��;F��;�ˢ;E��;�4�;�m;�O;��2;�;��:�@�:��:s?:R\9�����4����ź|�����50��kI��Eb���z�Sl���F����b��x�����»�ͻ,ػD���컍����\ ��/���	�>��(���u��]0 �c$��(�F�,�8�0�$j4��>8�4<��?��]C�	�F��J���M�rQ�w�T��7X�v�[���^�b�3Pe�.�h���k���n�7�q�(�t�%x�v{��~�V����	���������Nv���쇼_a���Ԋ�RG�������(�����W���s��H���L�����J!��抚���q\���Ğ�^,��Փ��#���Gb��]ɥ�|0�����������e���̬�-4��y�������i��'ѳ�p8���������n��;ֺ�>��N����  �  k�N=�N=�PM=ϛL=S�K=�0K=NzJ=��I=�I=�UH=̝G=��F=4-F=EtE=��D=D=�FC=��B=��A=�A=�W@=^�?=�>=�>=�\==��<= �;=�;=�R:=v�9=��8=>�7==67=�k6=��5=��4=�4=33=�`2=�1=��0=��/=�/=�#.=pC-=`,=�y+=C�*=a�)=��(=޾'=��&=��%=��$=/�#=�"=%�!=B� =;�=�f=�C=4=��=޷=�|=�;=��=3�=P=Q�=֑=�(=��=�B=�
= C	=й=�*=o�=��=4Z=�h�<�<G��<�I�<Q��<�[�<+��<�L�<D��<��<�}�<���<�)�<�v�<v��<,�<�B�<~�<ϵ�<%�<k�<�I�<vu�<ɞ�<�ŧ<��<��<7/�<+O�<�m�<N��<ۧ�<�È<J߄<~��<9+z<�ar<טj<��b<s
[<�ES<��K<��C<�<<�H4<�,<E�$<�)<�|<��<�/<q"�;3��;��;��;��;��;,ɢ;��;/2�;em;#�O;	�2;';��:�;�:N�:9:PH9m���4�����qźy������20�hI��Ab�.�z�Qj���D��l젻a��ݡ����»�ͻ++ػԛ⻑�컢���] ��/�h�	�Ҍ���������a1 �-d$���(�M�,�J�0�#k4��?8��<���?�y^C�z�F�Z�J���M��rQ�4�T��7X���[�,�^��b�UOe�@�h�{�k���n�'�q�%�t�x�Z{��~�틀�h	����K���$v��z쇼na��Պ�G��ȸ��)��b������=t�������L��}����!��h���t����\���Ğ��,�����X���fb��qɥ�n0��e��������e���̬��3�����/��di���г��7��4������	n���պ��=��	����  �  ��N=�N=QM=֛L=O�K=q0K=3zJ=��I=�I=EUH=��G=m�F=�,F=�sE=��D=� D=�FC=��B=T�A=PA=�W@=4�?=��>=�>=�\==�<=�;=;=�R:=��9=:�8=��7=~67=l6=L�5=��4=4=T33=�`2=X�1=µ0=��/=�/=�#.=yC-=%`,=�y+=/�*=A�)=в(=��'=��&=��%=��$=��#=��"=ٮ!=�� =��=�f=�C==r�=·=�|=�;=��=G�=7P=�=�=�(=L�=
C=a�
=aC	=+�=�*=͕=��=�Z=�i�<��<ó�<=J�<���<\�<H��<|L�<-��<��<�}�<L��<")�<�v�<��<��<B�<i}�<5��<��<��<HI�<u�<j��<ŧ<��<��<>/�<8O�<�m�<���<F��<DĈ<�߄<��<g,z<�br<�j<;�b<�[<�FS<K<��C<�<<5I4<��,<��$<*<�|<��<p/<
!�;���;���;ܰ�;���;���;�Ƣ;&�;u/�;�m;Z�O;�2;�;M��:�4�:��:M1:+=9���:�4��c źPs��r���.0��dI��=b���z�6h���B���꠻J_������»��ͻ5*ػ0��r�컏���G] �S0���	������ӌ����s2 �\e$�˃(���,�{�0�8l4��@8��<�z�?�/_C�	�F���J���M�wrQ��T�97X�q�[�b�^��b�UNe�<h�t�k���n���q���t��	x�S{��~�s������c������v��f쇼ia��#Պ��G�����l)��Ԙ��;���t��Wᔼ)M��"���m"����������q]��sŞ�-��h��������b��ɥ�`0��T���E���9e��J̬�f3����������h��	г�P7����������m��?պ�C=�������  �  ��N=N=QM=ޛL=J�K=\0K=zJ=k�I=oI=UH=G�G=�F=�,F=�sE=J�D=� D=4FC=m�B=�A=A=rW@=�?=��>=�>=�\==�<=%�;=1;=S:=�9=s�8=��7=�67=nl6=��5=H�4=S4=�33=a2=��1=��0=#�/=�/=$.=�C-=(`,=�y+=�*="�)=��(=w�'=o�&=m�%=-�$=��#=s�"=��!=�� =��=Xf=pC=�=J�=��=�|=|;=��=[�=`P=��=O�=@)=��=gC=��
=�C	=��=W+=/�=M�=�Z=j�<+�<-��<�J�<���<H\�<_��<kL�<��<|�<Y}�<���<�(�<�u�<?��<��<TA�<�|�<���<��<T�<�H�<�t�< ��<=ŧ<\�<��<D/�<TO�<3n�<ҋ�<���<�Ĉ<\��<���<�-z<]dr<u�j<��b<�[<HS<��K<��C<�<<�I4<N�,<��$<N*<�|<b�</<��;��;���;���;��;���;�â;�;�,�;��l;��O;�2;;!��:X-�:��:�(:�,9��2�4��돺��ĺn������*0�a`I�B9b�ݲz��e��K@��y蠻]��&���c�»=�ͻc)ػU��7�컙���}] ��0���	�V����������3 ��f$��(��,�ȇ0��m4��A8� <�^�?��_C���F��J�0 N�qrQ���T��6X��[���^��b�`Me�	~h�S�k�M�n���q���t��x�#{�^~����������������u��U쇼ia��JՊ��G��j����)��L������Nu��┼�M��и��#�����������]���Ş�z-��ʔ�������b���ɥ�T0��2��������d���ˬ��2��������=h��\ϳ��6��坶�\���l���Ժ��<��/����  �  ߺN=(N=.QM=�L=B�K=G0K=�yJ=K�I=7I=�TH=��G=��F=G,F=SsE=��D=- D=�EC= �B=��A=�A=?W@=�?=��>=�>=�\==�<=:�;=O;=JS:=�9=��8= 8=77=�l6=�5=��4=�4=�33=ca2=ی1=5�0=T�/=/=+$.=�C-=)`,=�y+= �*=��)=|�(=C�'=7�&=#�%=��$=I�#=�"=4�!=`� =d�=f=:C=�='�=��=�|=};=��=w�=�P=��=��=�)=�=�C= �
=$D	=��=�+=��=��=9[=�j�<��<���<�J�<!��<r\�<p��<hL�<��<Q�<}�<{��<,(�<fu�<���<T�<�@�<|�<鳾<X�<��<DH�<,t�<���<�ħ<$�<��<E/�<wO�<^n�<*��<��<8ň<���<B��<
/z<�er<�j<�b<n[<WIS<�K<�C<�<<�J4<Ñ,<J�$<m*<�|<�<�.<��;J��;���;<��;r��;���;���;�;�)�;f�l;H�O;��2;o;���:�'�:�ށ:u!:�9���?�4��鏺��ĺ�h��#��X'0��[I��4b�k�z�Pc���=���堻�Z��K�����»ۂͻL(ػ��⻿�컼����] �01��	����w�܎����5 ��g$���(�J�,��0��n4�%C8��<�6�?��`C��F�}�J�T N�xrQ���T�g6X�]�[���^��b�XLe��|h���k��n�G�q�K�t�Zx��{�K~�x��������������u��E쇼oa��cՊ�H������0*������D���u���┼mN��{����#��B���0����^��hƞ��-���������b���ɥ�N0����������d��{ˬ�u2��r���} ���g���γ��5��H������Ql��-Ժ�Q<��Ǥ���  �  �N=CN=AQM=�L=;�K=;0K=�yJ=$�I=I=�TH=��G=��F=�+F=sE=��D=��C=�EC=ߊB=��A=�A=
W@=ř?=��>=�>=�\==�<=N�;=l;=vS:=I�9=��8=R 8=^77=m6=@�5=��4=�4=<43=�a2=�1=n�0=�/=*/=@$.=�C-=%`,=�y+=��*=�)=M�(=	�'=��&=��%=��$=��#=ӻ"=�!=� ='�=�e= C=o=��=s�=�|=|;=��=��=�P=�=Ē=�)=:�=D=t�
=~D	=X�=,=�=�=�[=gk�<6�<��<VK�<b��<�\�<{��<lL�<���<�<�|�<��<�'�<�t�<,��<� �<@�<y{�<M��<��<,�<�G�<�s�<Z��<�ħ<�<x�<=/�<�O�<�n�<���<i��<�ň<n�<���<G0z<�fr<I�j<H�b<�[<sJS<?�K< �C<H<<dK4<?�,<��$<�*<|<��<.<>�;���;��;���;3��;k��;���;��;�&�;@�l;u�O;6�2;2;���:�!�:�ف:9:<9���[4�}珺��ĺ;d������#0�]XI�v0b��z��`���;���㠻/Y��b����»��ͻ;'ػ1��f�������] �~1���	�ʏ�m�ۏ����6 �6i$���(�~�,�W�0��o4�/D8��<�#�?�eaC���F�ςJ�| N��rQ�v�T�6X�̈[�C�^��b�JKe��{h�ߤk���n��q��t�1x��{�G~�􉀼���`���J���~u��0쇼{a��rՊ�PH����*��.������kv�� 㔼O�����W$��ڍ������_���ƞ�W.��a���N��� c���ɥ�Q0��疨�����Kd��(ˬ��1��혯������f��&γ�M5���������k���Ӻ��;��t����  �  (�N=]N=OQM=�L=3�K='0K=�yJ=��I=�I=bTH=��G=L�F=�+F=�rE=c�D=��C=\EC=��B=R�A=wA=�V@=��?=��>=�>=�\==$�<=_�;=�;=�S:=u�9= �8=� 8=�77=Om6=��5=0�4=44=z43=�a2=L�1=��0=��/=G/=V$.=�C-=-`,=�y+=ݏ*=Ƣ)=)�(=�'=��&=��%=_�$=��#=��"=��!=֚ =�=�e=�B=O=��=Z�=�|=s;=��=��=�P=4�=��=*=q�=\D=��
=�D	=��=e,=<�=O�=�[=�k�<��<y��<�K�<���<�\�<���<WL�<���<��<l|�<���<G'�<ut�<���<6 �<�?�<�z�<ò�<C�<��<`G�<js�<��<vħ<��<^�<J/�<�O�<�n�<���<���<ƈ<��<T��<I1z<hr<T�j<l�b<�[<�KS<5�K<��C<<<�K4<��,<��$<�*<f|<��<�-<�;_��;a��;���;��;��;ʻ�;�;�$�;O�l;��O;��2;��;���:��: ց:q:�9���}4�R叺0�ĺ�_�����R 0��TI��,b�+�z�3_���9��⠻'W������»��ͻp&ػ���(������)^ ��1��	�g�� �������47 �Aj$�(���,�Z�0��p4�E8��<���?��aC�#�F� �J�� N�|rQ�N�T��5X�[�[���^�Ub��Je��zh��k���n��q��t�!x��{�C~�����a��������Xu��쇼�a���Պ�rH��5����*��~���8	���v���㔼�O�������$��a���=����_��AǞ��.������{���(c���ɥ�@0��ʖ��m���d���ʬ��1������u����f���ͳ��4��&������Lk��7Ӻ��;������  �  >�N=sN=PQM=�L=5�K=0K=�yJ=��I=�I=5TH=Z�G="�F=�+F=�rE=)�D=o�C=(EC=u�B=(�A=JA=�V@=��?=��>=�>=�\==$�<=e�;=�;=�S:=��9=H�8=� 8=�77=m6=��5=^�4=j4=�43=b2=u�1=Ƕ0=��/=]/=i$.=�C-=.`,=�y+=Ώ*=��)=	�(=��'=��&=��%=1�$=��#=`�"=u�!=�� =��=we=�B=*=��=E�=�|=v;=��=��=�P=P�=�=:*=��=�D=��
=E	=޻=�,=w�=��=\=5l�<�<���<�K�<���<�\�<���<UL�<���<��</|�<~��<�&�<%t�<:��<���<?�<�z�<_��<��<c�<G�<s�<Ĝ�<Iħ<��<]�<H/�<�O�<�n�<䌐<��<aƈ<+�<���<2z<�hr<�j<O�b<�[<MLS<܈K<��C<�<<PL4<�,<��$<�*<u|<z�<d-<
�;3��;��;���;w��;T��;��;�;�"�;��l;��O;��2;��;���:�:Ӂ:�:��9����}4�-㏺��ĺ�Z��p��G0�rRI�*b�A�z��]��M8���࠻�U��旷���»�ͻ�%ػ��=������6^ �2���	�����o������7 ��j$���(�r�,��0��q4��E8��	<�^�?��bC���F�[�J�� N�wrQ�M�T��5X��[�8�^��b��Ie�0zh�8�k���n�G�q�B�t�\x�#{��~�Q�����肃�����Eu��쇼xa���Պ��H��k���(+��Ԛ���	��9w��䔼�O�����:%��Î�������_���Ǟ��.��액�����@c���ɥ�?0��ʖ��C����c���ʬ�S1��7������'f��2ͳ�w4������C���j���Һ�.;��ɣ���  �  L�N=~N=bQM=�L=-�K=0K=�yJ=��I=�I=%TH=>�G=�F=c+F=qrE=�D=J�C=	EC=T�B=�A=:A=�V@=z�?=r�>=�>=�\==.�<=t�;=�;=�S:=��9=c�8=� 8=�77=�m6=ء5=��4=�4=�43=-b2=��1=ֶ0=��/=j/=r$.=�C-=)`,=�y+=ď*=��)=��(=��'=��&=b�%=�$=k�#=B�"=Z�!=�� =��=Ve=�B==��=?�=�|=u;=��=��=�P=b�=%�=I*=ź=�D=�
=0E	=�=�,=��=��=(\=wl�</�<۵�<L�<���<�\�<���<OL�<x��<��<|�<_��<�&�<�s�<���<���<�>�<Pz�<��<��<#�<�F�<�r�<���<%ħ<��<O�<K/�<�O�<�n�< ��<��<�ƈ<h�<���<�2z<kir<��j<��b<[<�LS<X�K<��C<�<<�L4<N�,<E�$<�*<S|<U�<-<��;���;W��;���;a��;,��;鸢;�;�!�;W�l;e�O; �2;I�;���:%�:Ё:�:
�9O���z4�5⏺��ĺ~Z������0�^PI�#(b�`�z��\��7���ߠ�+U�����"�»�ͻ�%ػܗ⻿�����K^ �I2���	�!���������s8 ��k$��(��,���0�4r4�OF8��	<���?��bC���F���J�� N��rQ��T�^5X�Ӈ[�!�^�kb��Ie��yh���k���n���q���t��x��{�:~�������ւ������-u��쇼�a���Պ��H��~���D+�������	��{w��T䔼6P��E���}%��
�������`���Ǟ�/���������Sc���ɥ�;0������.����c��~ʬ�'1�����������e���̳�/4��}�������j���Һ��:�������  �  ��N=�N=�XM=7�L=L�K=:K=|�J=��I=FI=�aH=��G=��F= <F=!�E=��D=fD=�ZC=,�B=S�A=-A=r@=r�?=�>=�<>=�~==�<=��;=�>;=�|:=��9=X�8=�/8=�h7=��6=�5=5=Y?4=q3=נ2=��1=��0=G$0=�K/= p.=6�-=Q�,=n�+=W�*=��)=)=c(=�&'=y-&=�/%=�-$=='#=�"=!=�=��=\�=ݓ=Gg=s4=�=+�=st=�&=Q�=�v=q=�=�:=P�=hE=��	=�5=�==�o=w�=�# =w��<4��<��<��<��<(��<���<�^�<��<�<e�<C��<4��<J7�<�s�<=��<���<�<5@�<=k�<ȓ�<���<�ݫ<	��<��<�<�<�X�<xs�<Ќ�<Y��<���<Pӈ<g�<6��<�)z<NUr<k�j<�b<.�Z<�S<�<K<epC< �;<��3<6,<�W$<f�<��<�(<�v<U��;LG�;��;���;���;.��;N��;���;˂;h;��J;I|-;��;r�:2V�:�Wk:: �9=q:8�;Ź��O�'睺6JӺc� ���7�cQ�tj��W��%q���W��v	��܆��4λ��ƻ��ѻ�aܻ �滄�@��Ls��B����Q��d�������"��G&�p\*��\.��I2�j#6� �9���=��KA�o�D�*oH��K�H^O�*�R��V�;pY�.�\�l�_�n+c�Yf�vi�A�l���o��r���u��x���{���~� 瀼�`���؃�O���Æ�.7��u���j��w���J���dg��`Ԑ��@���������}���痼�O��ڶ�� ��	���C螼=M��ȱ��H���z���ޥ�MC��̧��|��q���լ��:��#���[���j��г�s5������ ���f���̺�j3��T����  �  ��N=�N=�XM=/�L=P�K=:K=��J=��I=VI=�aH=ЪG=��F=<F=0�E=�D=yD=�ZC=6�B=c�A=-A=r@=u�?=�>=�<>=�~==ܿ<=��;=�>;=�|:=��9=H�8=�/8=�h7=��6=�5=�5=P?4=�p3=٠2=��1=��0=,$0=tK/=+p.=,�-=M�,=v�+=c�*=��)=)=p(= ''=�-&=�/%=�-$=G'#=�"=�!=��=�=i�=�=Tg=y4= �=0�=nt=�&=Y�=�v=Q=ߪ=�:=O�=]E=��	=�5=r�=�=�o=u�=�# =U��<��<��<��<b�<$��<���<�^�<��<�<%e�<^��<K��<H7�<�s�<L��<���<�<5@�<^k�<ޓ�<ֹ�<�ݫ<��<��<�<�<�X�<ps�<ߌ�<*��<~��<3ӈ<^�<5��<�)z<'Ur<!�j<��b<�Z<�S<�<K< pC<��;<�3<@,<}W$<>�<��<�(<w<l��;�G�;��;G��;Ϯ�;[��;ԗ�;���;'̂;Nh;��J;�}-;t�;dt�:�V�:�Zk:t�9D�:8K@Ź��O�@睺�MӺ���u�7�)Q��j�X���q���W���	������tλ�o�ƻ��ѻEbܻ�����[��*s��B����$��/�f�����"��G&�C\*��\.�TI2��#6���9���=�UKA�6�D�oH���K�*^O�7�R�/V�pY�j�\���_��+c�QYf�ni�_�l���o�Q�r��u�"�x���{���~�B瀼a���؃�'O���Æ�I7��s���\��b���B���Bg��GԐ�i@���������X���痼�O��˶��"��ꂝ�/螼 M������9���z���ޥ�\C��֧��o��2q��#֬�;��-���[���j��г��5��,���� ���f��ͺ��3��x����  �  ��N=�N=�XM=.�L=S�K=":K=��J=��I=tI=�aH=��G=��F=7<F=d�E=&�D=�D=�ZC=f�B=��A=%-A=/r@=��?=�>=�<>=�~==ֿ<=��;=�>;=�|:=��9=!�8=�/8=�h7=y�6=��5=�5=*?4=�p3=��2=��1=�0= $0=`K/=#p.=�-=S�,=v�+=l�*=�)=!)=�(=''=�-&=0%=.$=r'#="=�!=%�=7�=��=�=hg=�4='�=+�=ot=�&=K�=�v=;=Ȫ=N:=�=E=��	=�5=;�=�=ao=A�=�# =0��<���<��<��<?�<"��<���< _�<���<L�<Re�<���<���<�7�<Kt�<���<Z��<��<�@�<�k�<��<��<�ݫ<C��<��<�<�<�X�<^s�<ӌ�< ��<m��<�҈<�<���<�(z<�Tr<W�j<V�b</�Z<�
S<<K<�oC<�;<��3<
,<HW$</�<��<�(<Lw<��;�H�;��;���;O��;��;���;<��;΂;�h;��J;m�-;��;y�:�Y�:�`k:�	�9��:8�>Ź��O��睺KOӺ'�����7�"Q�Cj�5Y���r���X��;������ϻ���ƻμѻ�bܻ������s�vB����ƕ��������o"��F&��[*��[.�kH2��"6��9��=��JA���D��nH���K�+^O��R�aV�0pY���\��_��+c�Zf��i�7�l�A�o��r���u���x���{���~��瀼"a��"ك�DO���Æ�[7��f���^��D���(���g��Ԑ� @��<�������~���痼PO��`�����������瞼�L���������z���ޥ�WC������_q��6֬�N;���������k��eг��5��x���K��-g��Yͺ��3�������  �  ��N=�N=�XM=0�L=W�K=4:K=��J=��I=�I=bH=1�G=��F=u<F=��E=p�D=�D=�ZC=��B=��A=[-A=Zr@=��?=>�>=�<>=�~==ٿ<=��;=�>;=�|:=]�9=��8=X/8=oh7=@�6=��5=�5=�>4=�p3=v�2=d�1=H�0=�#0=?K/=p.=�-=V�,=z�+=��*=(�)=J)=�(=N''=�-&=I0%=G.$=�'#=T"=�!=e�=f�=��=2�=�g=�4=<�=)�=kt=�&=$�=�v==��=:=��=�D=L�	=85=�=�=o=�=P# =���<R��<:�<���<.�<��<���</_�<:��<��<�e�< ��<��<8�<�t�<*��<���<�<A�<.l�<���<}��<ޫ<���<�<�<�<�X�<Ls�<���<���<��<�҈<��<`��<�'z<fSr<0j<-�b<6�Z<�	S<;;K<�nC<��;<�3<o,<�V$<'�<��< )<�w<0��;.J�;q	�;{��;\��;1��;���;Ϋ�;%Ђ;.h;�J;Y�-;��;��:H`�:lk:��9��:8k7Ź0�O�^ꝺ)RӺ�-�C�7�7%Q�Vj�![���t���Z���������
ѻ���ƻ�ѻ�cܻ���#����s�B�������������]"��E&�Z*��Z.��G2��!6�J�9�7�=�JA�.�D�KnH�6�K�^O�
�R�aV��pY�.�\���_��,c��Zf��i�&�l�1�o�&�r���u���x���{�]�~��瀼�a��kك��O��)Ć�U7��c���L����������f���Ӑ��?��Ҫ����w~��痼�N��굚�M��$����瞼�L��F������Zz���ޥ�SC���������q���֬��;��䠯�*���k���г��6���������g���ͺ�+4��򚽼�  �  ��N=�N=�XM="�L=c�K=O:K=ʄJ=��I=�I=ZbH={�G=S�F=�<F=��E=��D=@D=S[C=�B=�A=�-A=�r@=ʶ?=R�>==>=�~==ʿ<=��;=�>;=p|:= �9=��8=/8=h7=�6=B�5=+5=�>4=9p3="�2=!�1=�0=�#0=K/=�o.=
�-=J�,=��+=��*=A�)=r)=�(=�''=2.&=�0%=�.$=(#=�"=L!=��=��=��=d�=�g=�4=I�=6�=Wt=�&=�=gv=�=9�=�9=u�=pD=ڿ	=�4=z�==�n=��=�" =��<؃�<��<^��<��<���<���<B_�<a��<��<)f�<���<���<�8�<cu�<���<���<��<�A�<�l�<,��<<jޫ<���<D�<�<�<�X�<5s�<j��<��<���<҈<�<���<�&z<�Qr<�}j<��b<��Z<^S<�9K<�mC<��;<\�3<�,<�V$<ۘ<��<c)<x<R��;�K�;��;���;.��;L��;Ϟ�;V��;;ӂ;�h;��J;�-;��;���:2f�:uk:,�9�?;867Ź7�O��읺�UӺ�U���7��)Q�j#j��]��jw���]��K�������һ�7�ƻ��ѻ�dܻ&��~����r��A����f����օ�����"��D&��X*�4Y.�*F2�T 6��9���=�#IA���D��mH���K��]O�-�R��V��pY���\���_��-c��[f�@�i�v�l���o���r�B�u�,�x���{���~�q耼b���ك��O��PĆ�p7��d�����ۉ������]f��#Ӑ�?��4���_���}��C旼N��6�����������枼 L���������%z���ޥ�nC��!�������q��׬�/<��w������7l���ѳ�27��Ɯ��l��Ih��Sκ��4��g����  �  F�N=�N=yXM=�L=m�K=_:K=��J=<�I=I=�bH=ѫG=��F=7=F=d�E=6�D=�D=�[C=G�B=`�A=�-A=�r@=�?=y�>=#=>=�~==��<=��;=q>;=5|:=�9=`�8=�.8=�g7=}�6=��5=�
5=%>4=�o3=Ɵ2=��1=��0=�#0=�J/=�o.=��-=J�,=��+=��*=s�)=�)=5(=�''=�.&=�0%=/$=p(#="=�!=�=��=I�=��=�g=�4=V�=<�=Mt=�&=��=!v=~=�=X9=�=D=a�	=R4=�=�=An=-�=�" =k��<@��<S�<��<��<��<��<n_�<���<W�<�f�<0��<L��<�9�<=v�<���<e��<��<�B�<m�<͕�<���<�ޫ<. �<r�<�<�<�X�<s�<"��<��<+��<�ш<X�<���<�$z<2Pr<|j<�b<�Z<�S<k8K<DlC<��;<Q�3<.,<.V$<��<�<�)<�x<c��;N�;>�;���;:��;ͤ�;v��;���;ׂ;� h;��J;z�-;W�;��:	p�:b�k:Q=�9��;8?5Ź�O�W�A[Ӻ����j�7��.Q�.)j��`��?z��P`����������ջ��ƻ�ѻfܻ������Or�:A����N�������K��~"��B&�`W*��W.�hD2��6���9���=�HA�t�D�mH�|�K�p]O� �R��V�iqY���\�h�_��.c�%]f���i��l�J�o�&�r���u���x�Y�{��~�逼�b��6ڃ�%P���Ć��7��W����������+����e���Ґ�t>����������|���嗼MM��b������䀝�`枼�K��w���K��z���ޥ�vC��M���>��Zr��y׬��<��(�������l��tҳ��7������7��i��Ϻ�B5��ԛ���  �  �N=cN=`XM=�L=v�K=x:K='�J=m�I=`I=�bH=8�G=�F=�=F=ׅE=��D=D=\C=��B=��A=1.A=s@=7�?=��>=6=>=�~==��<=��;=M>;=�{:=��9=�8=X.8=Vg7=�6=n�5=Q
5=�=4=lo3=i�2=s�1=o�0=C#0=�J/=�o.=�-=K�,=��+=��*=��)=�)=�(=;('=�.&=_1%=o/$=�(#=}"=!=v�=e�=��=�=h=5=t�=;�=Et=j&=��=�u=,=~�=�8=��=C=�	=�3=z�==�m=��=-" =���<���<��<���<�<Ҍ�<��<�_�<��<��<)g�<ڲ�<��<W:�<w�<���<O��<s�<]C�<Zn�<w��<#��<j߫<� �<��<=�<�X�<�r�<勔<���<���<�Ј<��<)��<#z<eNr<zj<�b<.�Z<S<�6K<�jC<G�;<Z�3<�,<�U$<��<&�<�)<�y<���;dP�;��;A��;׻�;h��;m��;���;ۂ;q(h;y�J;��-;?�;S��:wx�:��k:P�9�<8r0Źy�O���f`Ӻ��$���7��4Q�6/j��c���}��^c��$��3����׻���ƻ��ѻcgܻ���N���r��@����d����0������"�!A&��U*��U.��B2�66���9�R�=��FA���D�:lH���K�A]O��R� V��qY�7�\�i�_�0c�q^f��i���l���o���r���u�{�x��{�q�~��逼(c���ڃ�rP���Ć��7��J������>�������Re��Ґ��=���������|���䗼gL������������垼K���������y���ޥ�{C��y������r��ج�t=��Ϣ��M���m��Nӳ��8��f������i���Ϻ��5��g����  �  �N=4N=IXM=�L={�K=�:K=K�J=��I=�I=HcH=��G={�F=>F=F�E=�D=�D=�\C=�B=�A=�.A=Vs@=i�?=��>=I=>=�~==��<=b�;=>;=�{:=N�9=��8=�-8=�f7=��6=��5=�	5=I=4= o3=��2=�1="�0=#0=�J/=�o.=ב-=D�,=��+=��*=��)=$)=�(=�('=F/&=�1%=�/$=L)#=�"=�!=��=��=�=4�=Qh=$5=��=:�=2t=P&=o�=�u=�=�=�8=�=�B=]�	=F3=�=�
=@m=A�=�! =���<��<U�<>��<J�<���<��<�_�<T��<8�<�g�<u��<���<1;�<�w�<��<4��<R�<2D�<o�<,��<ɼ�<�߫<� �<��<$=�<�X�<�r�<���<K��<��<6Ј<��<I��<d!z<�Lr<Dxj<%�b<h�Z<IS<=5K<jiC<�;<v�3<�,<;U$<P�<+�<Q*<z<���;�R�;��;��;;��;%��;G��;���;�ނ;_0h;��J;��-;ܞ;c��:��:�k:c�9T[<8�,ŹD�O�����dӺh�B(���7�g:Q�"5j��f�������f��=��_���tڻ���ƻ��ѻ�hܻ��滔�����q�@�%��a��B�ځ�,��"�n?&��S*�
T.��@2�{6���9��=�{EA���D��kH�W�K�]O� �R�P V��rY���\�X�_�B1c��_f�Ɇi�K�l���o���r�_�u�%�x���{��~�fꀼ�c��ۃ��P��ņ��7��L����������j����d��Tѐ�=��꧓����4{���㗼�K������L��h��垼fJ����������y���ޥ��C���������!s���ج�>������&	���n��4Գ��9��L�������j��wк��6����  �  ��N=N=9XM=�L=��K=�:K=u�J=��I=�I=�cH=�G=��F=s>F=��E=�D=�D=�\C=o�B=l�A=�.A=�s@=��?=��>=_=>=�~==��<=P�;=�=;=�{:=	�9=n�8=�-8=�f7=<�6=��5=�	5=�<4=�n3=��2=��1=��0=�"0=MJ/=`o.=Ñ-=>�,=��+=	�*=��)=[)=(=�('=�/&=!2%=;0$=�)#=K"=�!=3�=�=2�=h�=h=P5=��=C�="t=1&=G�=_u=�=˨=#8=��=�B=ڽ	=�2=x�=
=�l=��=b! =,��<c��<��<���<�<���<��<`�<���<��<Gh�<��<���<�;�<�x�<H��<���<%�<�D�<�o�<ؗ�<B��<e�<R�<0 �<C=�<�X�<�r�<>��<Ѣ�<���<�ψ<1�<���<�z<�Jr<�vj<^�b<��Z<�S<�3K<,hC<֞;<V�3<�,<�T$<�<>�<�*<�z<���;�T�;S�;��;f¾;���;���;=��;l�;g7h;?�J;��-;v�;J��:o��:��k:sv�9��<8z*Ź�O�i���wkӺ��>,�s�7�A?Q�,;j��i��~����i�����򖰻�ܻ���ƻ��ѻMjܻ��������q��?�P��t��S�w������"��=&�.R*�rR.�]?2�6�"�9���=��DA���D��jH���K��\O�.�R�� V��rY�ѻ\�h�_�I2c�af�1�i���l�l�o�:�r���u���x��{�{�~�뀼Id���ۃ�<Q��.ņ��7��J��������������_d���А�b<��2���4��qz���◼�J��籚�����~��s䞼�I��+���G��ay��uޥ��C������.���s��٬��>��?����	��po��ճ��:��!������Qk��#Ѻ�7������  �  |�N=�N=XM=��L=��K=�:K=��J=�I=I=�cH=2�G=,�F=�>F=	�E=��D=ND=C]C=ģB=��A=/A=�s@=ķ?=�>=o=>= ==��<=6�;=�=;=`{:=շ9="�8=N-8=;f7=�6=9�5=	5=�<4=Fn3=S�2=w�1=��0=�"0=/J/=Ko.=��-=@�,=��+=�*=�)=�)=F(=)'=�/&=q2%=�0$=*#=�"=B!=��=\�=n�=��=�h=i5=��=H�=t=&=%�=5u=R=��=�7=P�=%B=s�	=[2=
�=�	=hl=z�=! =���<���<}�<���<��<���<(��<`�<��<��<�h�<���<$��<�<�<xy�<���<���<��<�E�<op�<[��<ý�<��<��<\ �<h=�<�X�<}r�<��<���<*��<ψ<��<���<Cz<IIr<�tj<�b<+�Z<] S<z2K<�fC<��;<��3<x,<eT$<�<o�<�*<#{<͠�;�V�;d�;���;?ž;���;��;Y��;��;�=h;]�J;ީ-;;�;��:g��:�k:+��9�=8�+ŹD�O������nӺx�`0�i�7�8DQ�@@j�l��_���Gl�����6���#߻���ƻ��ѻkܻ\�滹���>q�7?�������V�j�`��J"�B<&��P*��P.��=2��6���9���=��CA���D�4jH���K��\O��R�� V�JsY�F�\��_�53c�Qbf�_�i�#�l���o���r�l�u�:�x�|�{���~��뀼�d���ۃ�nQ��\ņ��7��1���g�����������c��PА��;����������y��>◼J��2������~���㞼~I��ڮ����=y��Vޥ��C������W���s��x٬�%?��٤��|
��+p���ճ�P;��Ѡ��e���k���Ѻ��7��᝽��  �  U�N=�N=XM=��L=��K=�:K=��J=%�I=SI=dH=d�G=g�F=?F=N�E=�D=�D=|]C=��B=��A=C/A=�s@=�?=#�>=x=>=�~==��<=!�;=�=;=6{:=��9=��8=-8=�e7=��6=��5=�5=L<4=n3=�2=B�1=i�0=h"0=J/=,o.=��-=>�,=��+=4�*=9�)=�)=(=K)'=!0&=�2%=�0$=H*#=�"=y!=��=��=��=ҕ=�h=�5=��=@�=t=�%=��=u==A�=�7=�=�A=0�	=2=��=c	=l=:�=�  =$��<���<$�<g��<��<���<$��<M`�<��<F�<i�<���<���<=�<�y�<���<H��<S�<F�<�p�<���<8��<�<��<� �<e=�<�X�<ar�<ي�<?��<Ѹ�<�Έ<)�<o��<3z<QHr<�sj<�b<�Z<\�R<�1K< fC<2�;<�3<�,<T$<ȗ<`�<&+<�{<��;TX�;�;a��;?Ǿ;���;m��;�Ñ;>�;�Ah;r�J;n�-;�;���:㕮:��k:Î�9c1=8k)ŹG�O������rӺ!�c3�D�7��GQ�yCj�Wn��{����m����������໻�ƻ�ѻ/lܻ9������?q��>�=����e��~����T"�Y;&��O*��O.��<2��6���9���=��BA�>�D��iH�"�K��\O��R�!V��sY�׼\���_�4c�cf�-�i�2�l���o���r�u�u��x���{�p�~�쀼e��B܃��Q���ņ�8��9���\��O���u����c���ϐ�};�������+y���ᗼxI������r���}���㞼I���������y��]ޥ��C��������.t���٬��?��>����
���p��/ֳ��;��J������nl��#Һ�8��:����  �  D�N=�N=XM=��L=��K=�:K=��J=;�I=[I='dH=��G=��F=5?F=u�E=M�D=�D=�]C=*�B=�A=\/A= t@=��?=+�>=�=>=�~==��<=�;=�=;="{:=��9=��8=�,8=�e7=q�6=��5=�5=<4=�m3=�2=�1=N�0=N"0=�I/=o.=��-=6�,=��+=<�*=H�)=�)=�(=u)'=J0&=�2%=�0$=t*#="=�!=��=��=��=ܕ=�h=�5=��=G�=t=�%=��=�t= =�=`7=ٿ=�A=�	=�1=��=#	=�k=�=�  =���<R��<��<K��<��<j��<3��<S`�<<��<V�<Ai�<L��<���<i=�<Dz�<��<���<��<�F�</q�<��<K��<4�<��<� �<p=�<�X�<ar�<���<!��<���<tΈ<��<��<rz<oGr<'sj<�b<K�Z<��R<�0K<�eC<��;<��3<�,<T$<��<c�<I+<�{<���;�X�;'�;���;�Ⱦ;H��;Ǵ�;oő;��;NEh;��J;��-;�;���:h��:h�k:��9�;=8�'Źg�O�� ���tӺ�"��4���7�GJQ��Fj��o�������o��� ��%����ỻ��ƻ��ѻ�lܻ��������q��>����ʎ�8�~����z"��:&��N*�%O.�H<2��6�N�9�+�=�wBA���D�qiH��K�T\O�8�R�!V��sY��\��_�|4c��cf��i�תl���o���r�.�u���x�-�{�2�~�A쀼Se��m܃��Q���ņ�8��E���E��@���K���~c���ϐ�";��¥������x��Sᗼ'I��b�����]}��M㞼�H��m������y��Tޥ��C��������Lt��ڬ��?������I��q���ֳ�*<������F���l��wҺ�H8��w����  �  A�N=�N=XM=�L=��K=�:K=��J=X�I=lI=7dH=��G=��F=>?F=}�E=^�D=�D=�]C=)�B=�A=k/A=t@=�?=$�>=�=>= ==��<=�;=�=;={:=y�9=��8=�,8=�e7=h�6=��5=�5=<4=�m3=��2=�1=A�0=="0=�I/=o.=��-=6�,=��+=5�*=S�)=�)=�(=�)'=H0&=�2%=�0$=~*#="=�!=��=��=ϼ=�=�h=�5=��=S�=t=�%=��=�t=�=�=P7=ȿ=�A=ݼ	=�1=x�=	=�k=��=�  =���<>��<��<2��<��<s��<F��<@`�<c��<��<[i�<]��<���<~=�<Xz�<
��<���<��<�F�<.q�</��<i��<q�<��<� �<�=�<�X�<Pr�<���<��<t��<^Έ<��<���<gz<"Gr<sj<��b<:�Z<�R<�0K<meC<n�;<��3<|,<�S$<��<��<K+<�{<���;2Y�;��;���;�Ⱦ;���;��;Ƒ;��;Fh;��J;�-;�;���:u��:��k:ߛ�9�Y=8m*Ź��O����tuӺi#�T5���7�JQ�7Gj�6p��Ӊ��p��� ������⻻E�ƻ`�ѻ�lܻ���������p��>����J����}����q"��:&��N*��N.�(<2��6�V�9��=�CBA���D�:iH�'�K�\O�2�R�%!V�$tY�"�\�U�_��4c��cf�-�i�êl���o���r�\�u�(�x��{�r�~�X쀼me��܃��Q���ņ�8��;���1��S���#���Mc���ϐ�;��ƥ������x��2ᗼI��R�����^}��+㞼�H��0������y��<ޥ��C��%������Qt��)ڬ��?������\��q���ֳ�:<��ӡ��M���l���Һ�[8�������  �  D�N=�N=XM=��L=��K=�:K=��J=;�I=[I='dH=��G=��F=5?F=u�E=M�D=�D=�]C=*�B=�A=\/A= t@=��?=+�>=�=>=�~==��<=�;=�=;="{:=��9=��8=�,8=�e7=q�6=��5=�5=<4=�m3=�2=�1=N�0=N"0=�I/=o.=��-=6�,=��+=<�*=H�)=�)=�(=u)'=J0&=�2%=�0$=t*#="=�!=��=��=��=ܕ=�h=�5=��=H�=t=�%=��=�t== �=b7=ڿ=�A=�	=�1=��=%	=�k=�=�  =���<X��<�<P��<��<o��<8��<X`�<@��<Z�<Di�<O��<���<j=�<Ez�<��<���<��<�F�<-q�<��<H��<1�<��<� �<l=�<�X�<]r�<���<��<���<qΈ<��<��<oz<nGr<'sj<�b<M�Z<��R<�0K<�eC<��;<��3<�,<T$<��<k�<Q+<�{<���;�X�;2�;���;�Ⱦ;L��;ȴ�;nő;��;@Eh;��J;�-;��;s��:��:��k:���9�0=8)Ź!�O�T��)uӺ�"��4��7�pJQ��Fj��o�������o��� ��2����ỻ��ƻ��ѻ�lܻ��������q��>����̎�9�~����{"��:&��N*�%O.�H<2��6�O�9�+�=�wBA���D�riH��K�T\O�8�R�!V��sY��\��_�|4c��cf��i�תl���o���r�.�u���x�-�{�2�~�A쀼Se��m܃��Q���ņ�8��E���E��@���K���~c���ϐ�";��¥������x��Sᗼ'I��b�����]}��M㞼�H��m������y��Tޥ��C��������Lt��ڬ��?������I��q���ֳ�*<������F���l��wҺ�H8��w����  �  U�N=�N=XM=��L=��K=�:K=��J=%�I=SI=dH=d�G=g�F=?F=N�E=�D=�D=|]C=��B=��A=C/A=�s@=�?=#�>=x=>=�~==��<=!�;=�=;=6{:=��9=��8=-8=�e7=��6=��5=�5=L<4=n3=�2=B�1=i�0=h"0=J/=,o.=��-=>�,=��+=4�*=9�)=�)=�(=K)'=!0&=�2%=�0$=H*#=�"=y!=��=��=��=ӕ=�h=�5=��=@�=t= &= �=u= =C�=�7=�=�A=3�	=2=��=g	=l=?�=�  =.��<���</�<r��<��<���<.��<U`�<!��<M�<!i�<���<���<=�<�y�<���<H��<Q�<F�<�p�<���<2��<�<��< �<^=�<�X�<Zr�<Ҋ�<8��<˸�<�Έ<$�<l��<.z<NHr<�sj<�b<!�Z<b�R<�1K<fC<>�;<�3<�,<'T$<ؗ<p�<6+<�{<���;lX�;�;r��;KǾ;���;p��;�Ñ;7�;�Ah;N�J;@�-;ެ;'��:V��:��k:7��9 =8-,Ź��O�V ���sӺg!��3���7�HQ��Cj�{n�������m�����К���໻/�ƻ-�ѻ?lܻG������Cq��>�@����g��~����U"�[;&��O*��O.��<2��6���9���=��BA�>�D��iH�"�K��\O��R�!V��sY�׼\���_�4c�cf�-�i�2�l���o���r�u�u��x���{�p�~�쀼e��B܃��Q���ņ�8��9���\��O���u����c���ϐ�};�������+y���ᗼxI������r���}���㞼I���������y��]ޥ��C��������.t���٬��?��>����
���p��/ֳ��;��J������nl��#Һ�8��:����  �  |�N=�N=XM=��L=��K=�:K=��J=�I=I=�cH=2�G=,�F=�>F=	�E=��D=ND=C]C=ģB=��A=/A=�s@=ķ?=�>=o=>= ==��<=6�;=�=;=`{:=շ9="�8=N-8=;f7=�6=9�5=	5=�<4=Fn3=S�2=w�1=��0=�"0=/J/=Ko.=��-=@�,=��+=�*=�)=�)=F(=)'=�/&=q2%=�0$=*#=�"=B!=��=]�=o�=��=�h=j5=��=I�=t=&='�=7u=U=��=�7=T�=)B=w�	=`2=�=�	=nl=��=! =���<��<��<���<��<���<6��<&`�<��<��<�h�<���<*��<�<�<{y�<���<���<��<�E�<ip�<T��<���<��<��<Q �<]=�<�X�<rr�<��<���<!��<ψ<��<���<<z<FIr<�tj<�b<2�Z<g S<�2K<�fC<	�;<��3<�,<{T$<��<��<�*<8{<��;�V�;��;���;Qž;���;��;V��;��;b=h;*�J;��-;�;e��:���:g�k:���9��<8�/ŹA�O������oӺ���0���7��DQ��@j��l������ql�����Y���C߻���ƻ�ѻ,kܻp������Eq�=?�������Z�m�b��L"�C<&��P*� Q.��=2��6���9���=��CA���D�5jH���K��\O��R�� V�JsY�F�\��_�53c�Qbf�_�i�#�l���o���r�l�u�:�x�|�{���~��뀼�d���ۃ�nQ��\ņ��7��1���g�����������c��PА��;����������y��>◼J��2������~���㞼~I��ڮ����=y��Vޥ��C������W���s��x٬�%?��٤��|
��+p���ճ�P;��Ѡ��e���k���Ѻ��7��᝽��  �  ��N=N=9XM=�L=��K=�:K=u�J=��I=�I=�cH=�G=��F=s>F=��E=�D=�D=�\C=o�B=l�A=�.A=�s@=��?=��>=_=>=�~==��<=P�;=�=;=�{:=	�9=n�8=�-8=�f7=<�6=��5=�	5=�<4=�n3=��2=��1=��0=�"0=MJ/=`o.=Ñ-=>�,=��+=	�*=��)=[)=(=�('=�/&=!2%=<0$=�)#=L"=�!=3�=�=3�=h�=�h=Q5=��=E�=$t=3&=I�=bu=�=Ϩ='8=��=�B=�	=�2=�=
=�l=��=k! =>��<t��<��<��<!�<���<.��<`�<���<��<Sh�<'��<���<�;�<�x�<I��<���<"�<�D�<�o�<ϗ�<8��<Z�<E�<# �<5=�<�X�<�r�<2��<Ţ�<}��<�ψ<*�<���<�z<�Jr<�vj<b�b<��Z<�S<�3K<?hC<�;<n�3<�,<U$<4�<Y�<�*<�z<ǟ�;�T�;v�;2��;{¾;���;���;9��;^�;:7h;�J;3�-;�;p��:|��:��k:
r�9��<8B/Ź��O������lӺ���,��7��?Q��;j�+j������j�������ݻ���ƻ��ѻhjܻ��������q��?�V��y��W�z������"��=&�0R*�sR.�^?2�6�#�9���=��DA���D��jH���K��\O�.�R�� V��rY�һ\�h�_�I2c�af�1�i���l�l�o�:�r���u���x��{�{�~�뀼Id���ۃ�<Q��.ņ��7��J��������������_d���А�b<��2���4��qz���◼�J��籚�����~��s䞼�I��+���G��ay��uޥ��C������.���s��٬��>��?����	��po��ճ��:��!������Qk��#Ѻ�7������  �  �N=4N=IXM=�L={�K=�:K=K�J=��I=�I=HcH=��G={�F=>F=F�E=�D=�D=�\C=�B=�A=�.A=Vs@=i�?=��>=I=>=�~==��<=b�;=>;=�{:=N�9=��8=�-8=�f7=��6=��5=�	5=I=4= o3=��2=�1="�0=#0=�J/=�o.=ב-=D�,=��+=��*=��)=$)=�(=�('=F/&=�1%=�/$=L)#=�"=�!=��=��=�=5�=Rh=%5=��=<�=4t=R&=r�=�u=�="�=�8=�=C=c�	=M3=��=�
=Hm=J�=�! =���<��<i�<R��<^�<Č�<��<�_�<c��<F�<�g�<��<���<7;�<�w�<���<2��<O�<,D�<o�<"��<���<�߫<� �<��<=�<�X�<�r�<��<>��<��<+Ј<��<B��<[!z<|Lr<Dxj<*�b<q�Z<WS<N5K<iC<.�;<��3<�,<YU$<n�<I�<o*<-z<��; S�;��;?��;S��;4��;L��;���;�ނ;-0h;=�J;��-;s�;p��:��:˝k:'^�92<8�1Ź��O�`���HfӺ��(�V�7� ;Q��5j�Ag��򀍻�f��s�������ڻ���ƻ��ѻ�hܻ�滬�����q�@�,��g��G�݁�/��"�p?&��S*�T.� A2�|6���9��=�|EA���D��kH�W�K�]O� �R�P V��rY���\�X�_�B1c��_f�Ɇi�K�l���o���r�_�u�%�x���{��~�fꀼ�c��ۃ��P��ņ��7��L����������j����d��Tѐ�=��꧓����4{���㗼�K������L��h��垼fJ����������y���ޥ��C���������!s���ج�>������&	���n��4Գ��9��L�������j��wк��6����  �  �N=cN=`XM=�L=v�K=x:K='�J=m�I=`I=�bH=8�G=�F=�=F=ׅE=��D=D=\C=��B=��A=1.A=s@=7�?=��>=6=>=�~==��<=��;=M>;=�{:=��9=�8=X.8=Vg7=�6=n�5=Q
5=�=4=lo3=i�2=s�1=o�0=C#0=�J/=�o.=�-=K�,=��+=��*=��)=�)=�(=;('=�.&=_1%=o/$=�(#=}"=!=w�=f�=��=�=h=5=v�=<�=Gt=m&=��=�u=0=��=�8=��=�C=�	=�3=��==�m=��=6" =���<���<��<���<��<��<��<�_�<��<��<6g�<��<&��<]:�<#w�<���<M��<o�<WC�<Rn�<m��<��<]߫<� �<��<�<�<�X�<�r�<׋�<���<���<�Ј<��<"��<#z<`Nr<zj<�b<7�Z<)S<7K<�jC<`�;<u�3<�,<�U$<��<E�<*<�y<,��;�P�;��;b��;�;x��;r��;���;ۂ;=(h;0�J;?�-;ї;W��:_w�:�k:�J�9	�;8�5ŹI�O�?����aӺ^��$���7�05Q��/j�d���}���c��\��e���ػ���ƻ�ѻ�gܻ���f����r��@����j����4������"�#A&��U*��U.��B2�76���9�S�=��FA���D�:lH���K�B]O��R� V��qY�7�\�i�_�0c�q^f��i���l���o���r���u�{�x��{�q�~��逼(c���ڃ�rP���Ć��7��J������>�������Re��Ґ��=���������|���䗼gL������������垼K���������y���ޥ�{C��y������r��ج�t=��Т��M���m��Nӳ��8��f������i���Ϻ��5��g����  �  F�N=�N=yXM=�L=m�K=_:K=��J=<�I=I=�bH=ѫG=��F=7=F=d�E=6�D=�D=�[C=G�B=`�A=�-A=�r@=�?=y�>=#=>=�~==��<=��;=q>;=5|:=�9=`�8=�.8=�g7=}�6=��5=�
5=%>4=�o3=Ɵ2=��1=��0=�#0=�J/=�o.=��-=J�,=��+=��*=s�)=�)=5(=�''=�.&=�0%=/$=p(#="=�!=�=��=I�=��=�g=�4=X�==�=Ot=�&=��=$v=�=�=]9=�=D=g�	=Y4=	�=�=In=6�=�" =~��<S��<g�<��<��<���<��<_�<Ͻ�<e�<�f�<:��<T��<�9�<@v�<���<d��<��<|B�<wm�<Õ�<{��<�ޫ<  �<d�<�<�<�X�<s�<��< ��< ��<yш<P�<���<�$z<-Pr<|j<�b<�Z<�S<}8K<YlC<��;<l�3<K,<LV$<˘<2�<�)<�x<���;NN�;f�;���;R��;ܤ�;{��;���;�ւ;� h;V�J;"�-;�;��:�n�:�k:f8�9nz;8�:Ź��O��񝺝\ӺQ�N �
�7�k/Q��)j��`��~z���`��#�������ջ�D�ƻ2�ѻ>fܻ�����Xr�BA����S�������N���"��B&�bW*��W.�iD2��6���9���=�HA�u�D�mH�|�K�p]O� �R��V�iqY���\�h�_��.c�%]f���i��l�J�o�&�r���u���x�Y�{��~�逼�b��6ڃ�%P���Ć��7��W����������+����e���Ґ�t>����������|���嗼MM��b������䀝�`枼�K��w���K��z���ޥ�vC��M���>��Zr��y׬��<��(�������l��tҳ��7������7��i��Ϻ�B5��ԛ���  �  ��N=�N=�XM="�L=c�K=O:K=ʄJ=��I=�I=ZbH={�G=S�F=�<F=��E=��D=@D=S[C=�B=�A=�-A=�r@=ʶ?=R�>==>=�~==ʿ<=��;=�>;=p|:= �9=��8=/8=h7=�6=B�5=+5=�>4=9p3="�2=!�1=�0=�#0=K/=�o.=
�-=J�,=��+=��*=A�)=r)=�(=�''=2.&=�0%=�.$=(#=�"=L!=��=��=��=e�=�g=�4=J�=8�=Yt=�&=�=iv=�=<�=�9=z�=uD=�	=�4=��==�n=��=# =��<��<��<p��<	�<��<��<Q_�<p��<��<5f�<���<���<�8�<fu�<���<���<��<�A�<�l�<$��<㺯<^ޫ<���<7�<�<�<�X�<(s�<]��<s��<���<҈<�<���<&z<�Qr<�}j<��b<��Z<jS< :K<�mC<��;<t�3<,<�V$<��<�<~)<1x<���;�K�; �;��;C��;Z��;Ӟ�;R��;.ӂ;�h;��J;̉-;��;��:?e�:sk:�'�9�;8�;Ź��O��흺�VӺ�����7�H*Q��#j�^���w���]��{�����ӻ�Z�ƻ��ѻ�dܻ>�滓�,���r��A����k����څ�����"��D&��X*�5Y.�+F2�U 6��9���=�#IA���D��mH���K��]O�-�R��V��pY���\���_��-c��[f�@�i�v�l���o���r�B�u�,�x���{���~�q耼b���ك��O��PĆ�p7��d�����ۉ������]f��#Ӑ�?��4���_���}��C旼N��6�����������枼 L���������%z���ޥ�nC��!�������q��׬�/<��w������7l���ѳ�27��Ɯ��l��Ih��Sκ��4��g����  �  ��N=�N=�XM=0�L=W�K=4:K=��J=��I=�I=bH=1�G=��F=u<F=��E=p�D=�D=�ZC=��B=��A=[-A=Zr@=��?=>�>=�<>=�~==ٿ<=��;=�>;=�|:=]�9=��8=X/8=oh7=@�6=��5=�5=�>4=�p3=v�2=d�1=H�0=�#0=?K/=p.=�-=V�,=z�+=��*=(�)=J)=�(=N''=�-&=I0%=G.$=�'#=U"=�!=f�=f�=��=2�=�g=�4==�=*�=lt=�&=&�=�v==��=:=��=�D=Q�	==5=�=�=o=�=W# =���<a��<H�<���<=�<��<���<;_�<E��<��<�e�<��<��<8�<�t�<+��<���<�<A�<(l�<���<t��<ޫ<���<��<�<�<�X�<Bs�<���<���<���<�҈<��<[��<�'z<cSr<0j<0�b<=�Z<�	S<H;K<�nC<��;<�3<�,<W$<>�<��<)<�w<V��;PJ�;�	�;���;n��;<��;ě�;ʫ�;Ђ;	h;�J;�-;O�;L�:�_�:Tjk:-�9��:8Q;Ź-�O�^띺(SӺ������7��%Q��j�S[��
u���Z��
������*ѻ���ƻ1�ѻ�cܻ���4����s�B� �����������_"��E&��Z*��Z.��G2��!6�K�9�7�=�JA�/�D�LnH�6�K�^O�
�R�aV��pY�.�\���_��,c��Zf��i�&�l�1�o�&�r���u���x���{�]�~��瀼�a��kك��O��)Ć�U7��c���L����������f���Ӑ��?��Ҫ����w~��痼�N��굚�M��$����瞼�L��F������Zz���ޥ�SC���������q���֬��;��䠯�*���k���г��6���������g���ͺ�+4��򚽼�  �  ��N=�N=�XM=.�L=S�K=":K=��J=��I=tI=�aH=��G=��F=7<F=d�E=&�D=�D=�ZC=f�B=��A=%-A=/r@=��?=�>=�<>=�~==ֿ<=��;=�>;=�|:=��9=!�8=�/8=�h7=y�6=��5=�5=*?4=�p3=��2=��1=�0= $0=`K/=#p.=�-=S�,=v�+=l�*=�)=!)=�(=''=�-&=0%=.$=r'#="=�!=%�=7�=��=�=hg=�4=(�=,�=pt=�&=M�=�v===ʪ=Q:=�=!E=��	=�5=?�=�=eo=F�=�# =:��<���<��<���<I�<,��<���<	_�<��<S�<Xe�<���<���<�7�<Mt�<���<Z��<��<�@�<�k�<��<��<�ݫ<<��<��<�<�<�X�<Ws�<̌�<���<g��<�҈<�<���<�(z<�Tr<W�j<Y�b<3�Z<�
S<"<K<�oC<��;<��3<,<XW$<?�<��<�(<[w<��;�H�;��;���;\��;��;���;9��;΂;jh;ٯJ;?�-;L�;�x�:;Y�:�_k:l�9��:8�AŹC�O��蝺�OӺ��2��7�S"Q��j�XY��s��Y��W��&����ϻ��ƻ�ѻ�bܻ���,� ��#s�yB����ɕ���������p"��F&��[*��[.�lH2��"6��9��=��JA���D��nH���K�+^O��R�aV�0pY���\��_��+c�Zf��i�7�l�A�o��r���u���x���{���~��瀼"a��"ك�DO���Æ�[7��f���^��D���(���g��Ԑ� @��<�������~���痼PO��`�����������瞼�L���������z���ޥ�WC������_q��6֬�N;���������k��eг��5��x���K��-g��Yͺ��3�������  �  ��N=�N=�XM=/�L=P�K=:K=��J=��I=VI=�aH=ЪG=��F=<F=0�E=�D=yD=�ZC=6�B=c�A=-A=r@=u�?=�>=�<>=�~==ܿ<=��;=�>;=�|:=��9=H�8=�/8=�h7=��6=�5=�5=P?4=�p3=٠2=��1=��0=,$0=tK/=+p.=,�-=M�,=v�+=c�*=��)=)=p(= ''=�-&=�/%=�-$=G'#=�"=�!=��=�=i�=�=Tg=y4= �=1�=nt=�&=Z�=�v=Q=�=�:=Q�=^E=��	=�5=t�=�=�o=w�=�# =Z��<��<��<��<g�<)��<���<�^�<��<#�<)e�<a��<M��<J7�<�s�<L��<���<�<3@�<\k�<ܓ�<ӹ�<�ݫ<��<��<�<�<�X�<ls�<܌�<'��<{��<0ӈ<[�<3��<�)z<&Ur<!�j<��b<�Z<�S<�<K<&pC<��;<�3<H,<�W$<F�<��<�(<w<z��;�G�;��;P��;ծ�;_��;֗�;���;#̂;Ah;��J;k}-;X�;#t�:�V�:;Zk:"�92x:8�AŹw�O��睺NӺA����7�RQ��j� X���q���W���	��ˆ���λ�z�ƻ��ѻMbܻ�����a��,s��B����&��1�g�����"��G&�C\*��\.�TI2��#6���9���=�UKA�6�D�oH���K�*^O�7�R�/V�pY�j�\���_��+c�QYf�ni�_�l���o�Q�r��u�"�x���{���~�B瀼a���؃�'O���Æ�I7��s���\��b���B���Bg��GԐ�i@���������X���痼�O��˶��"��ꂝ�/螼 M������9���z���ޥ�\C��֧��o��2q��#֬�;��-���[���j��г��5��,���� ���f��ͺ��3��x����  �  ��N=�N=R`M=��L=��K=DDK=��J=��I=%I=noH=i�G=4G=�LF=�E=��D=�'D=0pC=G�B=��A=4GA=Ѝ@=��?=1?=�]>=��==f�<=>&<=g;=��:=��9=W#9=�_8=�7=�6=�6=�D5=�z4=�3=B�2=�2=f@1=�l0=͖/=P�.=2�-=+-='$,=�?+=]X*=Km)=�~(=��'=J�&=��%=B�$=r�#=Ԏ"=$�!=:n =�U=v7=)=��=��=�=A=M�=p�=>Z=��=�=�1=��=1H=��=�B
=t�=�!=�=��=�A=Q� =*��<O]�<5��<�e�<���<I�<J��<��<b�<|��<���<n>�<�|�<M��<d��<��<9J�<�t�<���<���<��<Q�<��<g;�<U�< m�<N��<*��<���<!��<�ό<e��<���<� �<� z<�@r<aj<C�b<�Z<��R<j�J<bC<N@;<�l3<�+<n�#<�<�<<�y<c�<�;s��;�?�;���;��;-��;�b�;�W�;"`�;��b;RhE;Q(;��
;y��:E#�:NR:��9�s������9l�Ȁ���D�|��"�%���?�5GY��cr����浑������d���괻8���M˻�+ֻz���?�gv���v�����jk	�������0���� ��$��8(��B,�p70�s4�4�7�;�;��L?���B��sF���I�lbM���P�S T��nW���Z���]�x"a�DMd�pg���j�h�m�k�p�`�s�u�v��y���|���<G��޼���0�������΃����p`��g͌�S9���������nx��ᓼ�H��ܯ�����/{���ߚ�tC��Ʀ��y	���k��Ρ�70��;���P����V����������~���ᬼ�D��K������To��ӳ��6�����������b��Ǻ��+�������  �  ��N=�N=H`M=��L=��K=QDK=��J=��I=$%I=xoH=y�G=@G=�LF=�E=	�D=�'D=;pC=T�B= B==GA=��@=��?=H?=�]>=��==\�<=;&<=g;=�:=��9=D#9=�_8=��7=��6=�6=�D5=�z4=Ԯ3=C�2=�2=Z@1=�l0=/=O�.='�-=(-=*$,=�?+=hX*=Vm)=�~(=��'=^�&=��%=V�$=��#=�"=9�!=An =�U=�7=4=��=��=�=A=M�=c�=;Z=��=��=�1=��=.H=��=fB
=^�=�!=�=��=�A=:� =��<"]�<��<ze�<���<I�<Z��<��<b�<���<���<}>�<�|�<^��<���<��<aJ�<�t�<��<���<��<{�< �<�;�<2U�<m�<D��<��<���<���<�ό<J��<���<| �<� z<[@r<�`j<��b<y�Z<��R<N�J<C<@;<�l3<��+<=�#<�<�<<*z<��<O�;���;@�;K��;���;���;tc�;�W�;�`�;��b;\iE;9(;��
;��:%�: &R:���9��r�7����9l�	����F⺯���%���?��GY��dr�s���^���	���We���괻L8��:N˻�+ֻ��໿?뻷v���v�����2k	������D0�|������$�c8(�=B,�*70�4��7��;��L?���B��sF�[�I�3bM���P�M T�oW���Z���]��"a�pMd�Xpg���j���m�®p���s���v�T�y��|���aG�����0�������ト���Y`��>͌�A9��������[x�������H���������{���ߚ�_C������_	���k���͡�0�����L����V���������~���ᬼ�D��X�������o��0ӳ��6��Ú�������b��Ǻ��+��͐���  �  z�N=�N=<`M=��L=��K=VDK=��J=��I=O%I=�oH=��G=vG=�LF=I�E=@�D=(D=rpC=��B=6 B=fGA=	�@=�?=V?=�]>=��==Z�<=.&<=g;=Ʀ:=��9=#9=�_8=7=��6=k6=�D5=qz4=��3=�2=�2=3@1=�l0=��/=B�.=�-=/-=,$,=@+=|X*=sm)=�~(='�'=��&=��%=��$=��#=�"=y�!=tn =�U=�7=W=��=��=�=A=N�=S�=$Z=��=ϛ=�1=Z�=�G=q�= B
=�=�!=��=��=�A=�� =���<�\�<���<Je�<���<I�<N��<��<0b�<ڱ�<7��<�>�<H}�<Ŷ�<��<0�<�J�<7u�<���<��<�<��<C �<�;�<JU�<m�<X��<��<���<̽�<Oό<�߈<%��< �<�z<{?r<�_j<�b<f�Z<��R<m�J<:C<�?;<l3<��+<��#<�<�<<4z<�<��;R��;pA�; ��;V��;���;�e�;�Y�;Cc�;�c;�mE;-(;��
;y��:�(�:c,R:���9��r�����&:l�Ձ��6I�ܳ���%��?��JY�zhr������������$g��촻�9��PO˻�,ֻi��
@��v���v��}���j	�Q����/�˔����$�[7(�PA,�C60�4�;�7��;�L?��B��rF��I��aM���P�, T�;oW�6�Z��]�&#a��Md�8qg�Ìj���m���p���s���v�K�y�֭|�����G��(���1��<���*��냈���S`��#͌�9��1�������w������]H��*���X���z��ߚ��B��1���	��k���͡��/�����B����V��%�������~���ᬼSE��¨��J���o���ӳ�m7��/���3���5c���Ǻ�&,������  �  R�N=fN=#`M=��L=��K=oDK=яJ=��I=�%I=�oH=��G=�G=RMF=��E=��D=c(D=�pC=ݸB=� B=�GA=?�@=9�?=y?=�]>=��==S�<=&<=�f;=��:=F�9=�"9=<_8=p�7=g�6=6=MD5=z4=C�3=��2=[2=�?1=dl0=��/=�.=�-=+-=7$,=@+=�X*=�m)=�~(=n�'=ݕ&=�%=�$=�#=y�"=ǁ!=�n =AV=�7=�=��=��=�=A=@�=<�=�Y=l�=��=h1=�=�G=�=�A
=��=!=9�=4�=LA=�� =��<I\�<x��<�d�<T��<�H�<Z��<�<�b�<3��<���<e?�<�}�<u��<���<��<�K�<�u�<2��<���<��<P�<� �<<�<�U�<4m�<X��<䗘<F��<���<�Ό<s߈<��<h��<7z<�=r<7^j<�b<�Z<6�R<&�J<'C<�>;<Vk3<��+<�#<�<=<�z<�<��;��;�C�;���;��;���;�h�;l]�;Mf�;�c;esE;�(;��
;>��:R1�:C9R:\�9�Or�9��.>l�����GM� ����%�?�?�MOY��lr������������si��\�;��Q˻S.ֻs��
A�7w���v��A��mj	���+���.��������$�6(��?,��40��4���7�۟;��J?��B�*rF�Q�I�yaM���P�8 T�foW�ǴZ���]��#a��Nd�-rg���j��m���p��s��v���y�$�|���GH������d1������n��������.`���̌��8��ǣ����aw���ߓ��G����������y��gޚ�JB���������k��a͡��/��ܑ��2����V��P�����,��g⬼�E��P�������p��PԳ�8��盶������c��Ⱥ��,������  �  �N==N=`M=��L=��K=�DK=��J=�I=�%I=CpH=^�G=<G=�MF=�E=$�D=�(D=HqC=J�B=� B= HA=��@=u�?=�?=^>=��==I�<=�%<=�f;=a�:=��9={"9=�^8=�7=��6=�6=�C5=�y4=ԭ3=Q�2=�2=�?1= l0=V�/=��.=�-=%-=K$,=?@+=�X*=�m)=F(=Ќ'=B�&=��%=U�$=��#=�"=4�!==o =�V=K8=�=%�=�=�=A=.�=!�=�Y=/�=8�= 1=��=G=��=(A
=�=� =��=��=�@=6� =H��<�[�<���<�d�<��<�H�<q��<<�<�b�<���<H��<@�<�~�<i��<���<��<�L�<�v�<&��<�·<��<��<O!�<�<�<�U�<Ym�<Q��<ϗ�<���<!��<EΌ<�ވ<��<���<_z<�;r<[\j<{}b<�Z<T�R<`�J<�C<'=;<^j3<6�+<�#<S<=<�z<"�<��;w��;�F�;���;���;Ɗ�;�l�;�a�;Tj�;�c;[{E;#(;��
;���:W;�:HHR:(�9��q�Uz���>l������Q���J�%���?�)UY��sr�����ؽ�������l���񴻎>��wS˻40ֻ����A�ow���v��ٟ��i	�����X-������$�44(��=,��20��4���7�/�;�SI?���B�qF��I��`M�0�P�F T��oW�>�Z�W�]��$a�KPd��sg���j���m��p�̺s��v�w�y�Ұ|�����H��L����1��ۣ�����������_���̌�H8��9���P���v��ߓ��F����������x��uݚ�^A��֤�����yj���̡�D/����������V��m���k������⬼uF���������q��Hճ��8��ܜ��� ���d���Ⱥ�I-������  �  ��N=	N=�_M=��L=��K=�DK=0�J=\�I=*&I=�pH=ӺG=�G=TNF=��E=��D=e)D=�qC=ƹB=SB=cHA=ߎ@=��?=�?=%^>=��===�<=�%<=zf;=�:=��9="9=_^8=��7=i�6=6=LC5=y4=O�3=��2=�2=D?1=�k0=�/=ν.=��-=&-=[$,=c@+=Y*=8n)=�(=5�'=��&=�%=�$=�#=t�"=��!=�o =W=�8=,=l�=�=�=A="�=��=�Y=��=Ӛ=�0=�=}F=��=�@
=x�=�=�=�=9@=�� =j��<�Z�<I��<d�<���<�H�<u��<s�<Cc�<A��<���<�@�<��<a��<���< �<�M�<�w�<(��<�÷<Y�<��<�!�<�<�<$V�<�m�<S��<���<���<���<�͌<�݈<��<���<7z<�9r<�Yj<3{b<ٝZ<7�R<g�J<�C<�;;<i3<?�+<��#<<5=<\{<�<�
�;d��;J�;���;,��;f��;�q�;�f�;no�;;c;d�E;�(;j�
;���:{F�:�YR:"?�9�mq�Nu���Al�����HY����%��?�\Y�{r�ʙ����������kp�������A��V˻m2ֻ���C��w��dv�����1i	�������+�Y��#���$��1(��;,��00��4���7�D�;��G?�?�B��oF�z�I�U`M���P�2 T��oW�ڵZ�q�]�:&a��Qd�yug���j���m��p���s��v���y�ʲ|�i���I������u2��[������/������_��>̌��7����������u��ޓ��E��~�������w��bܚ�g@��裝�����i��N̡��.��]����󥼳V���������%����㬼=G���������r��Zֳ� :��흶�����e���ɺ�.�������  �  ��N=�N=�_M=��L=��K=�DK=j�J=��I=�&I=qH=V�G=@G=�NF==�E=@�D=�)D=TrC=O�B=�B=�HA=7�@=��?=?=@^>=��==&�<=�%<=Cf;=å:=@�9=�!9=�]8=��7=��6=v6=�B5=�x4=��3=X�2=2=�>1=xk0=̕/=��.=��-= -=j$,=�@+=LY*=}n)=�(=��'==�&=��%=n�$=��#=�"=L�!=4p =�W=9=�=��=K�=/�="A=�=ʭ=NY=��=f�=0=��=�E=A�=�?
=��=3=Z�=i�=�?="� =i��< Z�<���<�c�<m��<�H�<���<��<�c�<г�<���<�A�<���<l��<���<3!�<�N�<y�<C��<�ķ<C�<��<�"�<�=�<xV�<�m�<I��<f��<J��<��<�̌<݈<��<o��<�z<D7r<VWj<�xb<_�Z<�R<_�J<�C<:;<�g3<P�+<��#<�<L=<�{<Ҿ<��;v��;�M�;.�;�¼;;��;�v�;�k�;�t�;$%c;j�E;�&(;��
;���:�Q�:�mR:�X�9��p��u���El������`���� &���?�	dY�%�r����eƑ������t������E��Y˻�4ֻs�� D뻻x��_v��*��qh	������(*�}������$��/(�=9,�5.0�Q4���7��;��E?���B��nF���I��_M���P�7 T�_pW�|�Z�j�]��'a�LSd�9wg���j��m�K�p�o�s�k�v�սy��|�R���J������3��Τ��0��e���u򉼞_���ˌ�E7��塏�����t��ݓ��D��O���[���v��Eۚ�V?��ܢ�����h���ˡ�`.��������V��깨�-������T䬼H��髯�����s���׳�Z;���������f���ʺ��.��w����  �  C�N=�N=�_M=v�L=��K=�DK=��J=��I=�&I=�qH=ͻG=�G=sOF=јE=��D=�*D=�rC=ԺB=DB=:IA=��@==�?=3?=c^>=��==�<=�%<=	f;=}�:=��9=/!9=_]8=m�7=I�6=�
6=B5=�w4=4�3=��2=�2=n>1=%k0=��/=n�.=��-=-=�$,=�@+=�Y*=�n)=k�(=�'=��&=�%=��$=?�#=��"=Ճ!=�p =X=}9=�=��=|�=I�=/A=��=��=Y=/�=�=�/=��=CE=��=)?
=�=~=��=��=�>=�� =e��<AY�< ��< c�<"��<�H�<���<��<d�<l��<}��<�B�<���<���<��<k"�<P�<Fz�<k��<�ŷ</�<a�<3#�<�=�<�V�<�m�<D��<7��<ᩔ<���<8̌<I܈<��<P��<�z<�4r<�Tj<-vb<�Z<��R<'�J<C<h8;<sf3<A�+<4�#<<y=<X|<��<i�;���;LQ�;)�;|Ǽ;?��;|�;3q�;�y�;�/c;�E;�/(;��
;^��:�]�: R:v�9Jmp�7q��Il�L����f�1���&���?��kY�0�r�y����ʑ������x�������H��'\˻;7ֻ,�໌E�Hy��Uv������g	���&��}(�������6$�T-(��6,��+0�4�t�7�!�;�D?���B�9mF���I��^M�)�P�8 T��pW�C�Z�[�]��(a��Td�yg���j��m���p���s���v��y�5�|�v���K�������3��A����������g�\_��~ˌ��6��2����
���s��
ܓ�yC��/���$��mu��#ښ�:>��록�=��9h��'ˡ��-��ʐ�����V��!������8���嬼�H��謯�����t���س�|<��F������g���˺��/��1����  �   �N=kN=�_M=h�L=��K=EK=ҐJ=9�I=:'I=�qH=@�G=HG=�OF=Y�E=n�D=+D=ksC=O�B=�B=�IA=�@=��?=d?=}^>=��==�<=n%<=�e;=5�:=��9=� 9=�\8=�7=��6=P
6=�A5=\w4=��3=R�2=+2=>1=�j0=J�/=C�.=��-=-=�$,=�@+=�Y*=o)=��(=�'=(�&=��%=~�$=Ě#=!�"=X�!=9q ={X=�9=6=9�=��=a�=4A=��=��=�X=��=��=/=t�=�D=�=>
=m�=�=�=.�=m>=� =~��<yX�<X��<�b�<���<[H�<���</�<�d�<���<%��<~C�<|��<���<��<�#�<(Q�<Y{�<o��<�Ʒ<�<�<�#�<}>�<W�<n�<1��<��<���<��<�ˌ<}ۈ<��<O��<`z<e2r<�Rj<�sb<��Z<t�R<*�J<SC<�6;<@e3<S�+<��#<+<�=<�|<m�<��;?��;�T�;	�;�˼;͝�;ˀ�;Lv�;�~�;#9c;	�E;8(;_;��:�i�:�R:��9Zp��n��LLl�%����m����&�y�?�lrY��r�v����Α�3���3|��- ���K���^˻�9ֻ�໮F뻪y��jv��L��g	���٪�'�����/$�)+(��4,��)0��
4�h�7�>�;�EB?���B��kF�z�I�V^M���P�J T��pW��Z�]�]�*a�oVd��zg���j��m��p���s���v�O�y�$�|�S��jL��G���@4�������������i�._��#ˌ�.6������'
�� s��ۓ�qB�������^t��ٚ�>=�����d���g���ʡ��-���������V��S�����������嬼�I��̭������u���ٳ��=��f������h���̺��0��唽��  �  ��N=AN=y_M=a�L=��K=EK=��J=n�I=�'I=CrH=��G=�G=lPF=ԙE=��D=�+D=�sC=��B=B=�IA=*�@=��?=�?=�^>=��==��<=L%<=�e;=�:=4�9=g 9=�\8={�7=F�6=�	6=A5=�v4=9�3=��2=�2=�=1=�j0=�/= �.=��-=-=�$,=�@+=�Y*=Wo)=�(=ڎ'=��&=��%=�$=6�#=��"=̈́!=�q =�X==:=�=n�=ָ=s�=4A=��=Y�=�X=��=C�=�.=��=3D=y�=�=
=ڰ=I=y�=��=�==�� =���<�W�<���<Jb�<���<GH�<���<^�<�d�<l��<���<;D�<N��<h��<��<r$�<R�<K|�<O��<kǷ<��<��<S$�<�>�<QW�<$n�<5��<ז�<9��<���<�ʌ<�ڈ<.�<j��<Zz<�0r<�Pj<�qb<��Z<��R<|�J<�	C<�5;<#d3<��+<�#<�<�=<}<�<��;ǯ�;�W�;|�;pϼ;���;��;;z�;)��;5Ac;��E;�?(;�;V	�: r�:�R:��9b�o�Km��sPl�񝬺Rt⺵��P&��?�yY��r�䩅�.ґ�tĝ����M���N��ua˻�;ֻ��໛G�Wz��+v�����f	������%�j��Z��x
$�>)(��2,��'0��4���7���;��@?�;�B��jF���I��]M���P�; T�WqW�g�Z�2�]�*+a��Wd�M|g�>�j��m���p���s���v�'�y��|���1M�������4�����
��˄��^�_���ʌ��5��
���~	��7r��=ړ��A��$��� ��js��+ؚ�g<��4�������f�� ʡ�.-��c������V������L��6���I欼jJ����������v���ڳ��>��K������i��fͺ�P1��w����  �  ��N=N=a_M=\�L=��K=9EK="�J=��I=�'I=rH=�G=G=�PF=0�E=6�D=�+D=.tC=�B=bB=.JA=f�@=��?=�?=�^>=¡==��<=2%<=xe;=��:=��9=! 9=9\8=&�7=��6={	6=�@5=�v4=ߪ3=��2=~2=v=1=Tj0=ߔ/=��.=p�-=-=�$,=A+=Z*=�o)=N�(=�'=ߘ&=L�%=D�$=��#=�"=�!=�q =+Y=u:=�=��=��=��=5A=��=>�=qX=X�=�=g.=��=�C=�=�=
=g�=�=�=9�=�==D� =#��<>W�<b��<�a�<f��<;H�<���<��<e�<ӵ�<0 �<�D�<��<
��<���<&%�<�R�<�|�<���<ȷ<O�<E�<�$�<.?�<�W�<6n�<1��<���<�<��<�ʌ<=ڈ<��<���<�z</r<�Nj<epb<?�Z<&�R<6�J<�C<�4;<3c3<�+<��#<�<�=<h}<��<��;ڱ�;�Y�;�;4Ҽ;���;5��;Q}�;Y��;Gc;ԮE;�D(;{;��:�x�:ثR:ɮ�99^o��k��Tl������y⺖��&��?��}Y���r�����Ց��Ɲ�w���u���P��Ec˻/=ֻ�໎H��z��v��ޝ�f	�J����$�t����#	$��'(�B1,�;&0��4�^�7�H�;��??�9�B�&jF�1�I�O]M�z�P�2 T��qW��Z���]��+a��Xd�r}g�c�j�V�m��p�b�s�^�v�n�y�_�|����M��Z�65��q���D������T��^���ʌ��5������	���q���ٓ��@��t���m���r���ך��;������<��uf���ɡ��,��(���~�W��������������欼�J��&���Q��vw��^۳�Y?���������Oj���ͺ��1��啽��  �  w�N=
N=]_M=U�L=��K=EEK=.�J=��I=�'I=�rH=$�G==G=�PF=f�E=u�D=$,D=ltC=B�B=�B=ZJA=��@=��?=�?=�^>=��==��<=(%<=ee;=��:=��9=�9=\8=�7=��6=>	6=z@5=Tv4=��3=`�2=M2=O=1=.j0=Δ/=�.=m�-=	-=�$,=A+=&Z*=�o)=k�(=K�'=�&=��%=�$=ƛ#=!�"=V�!=*r =[Y=�:=�=��=�=��=6A=��=5�=[X=>�=֘=7.=l�=�C=��=J=
=%�=�=͂=��=U==� =���<�V�<(��<�a�<S��< H�<���<��<3e�<��<| �<!E�<P��<���<(��<�%�<JS�<t}�<n��<rȷ<��<��<�$�<P?�<�W�<9n�<$��<���<֨�<���<1ʌ<�و<#�<L��<�z<�-r<�Mj<Job<F�Z<;�R<G�J<�C<�3;<�b3<��+<��#<�<�=<�}<��<��;ò�;Q[�;��;Լ;���;��;�;>��;yKc;��E;�H(;�;�:�|�:��R:��9�Zo��i���Tl�/���|⺵��P&�>�?��Y�(�r�W����֑��ȝ����;��2R��gd˻D>ֻw���H��z��Pv����e	������9$����G��,$��&(�^0,�Q%0��4�f�7�y�;��>?���B��iF���I�]M�[�P�S T��qW� �Z�9�]��,a�VYd�,~g�N�j�-�m���p�C�s�J�v�n�y�9�|����N����m5������^��儈�b��^��zʌ�T5��]������Eq��3ٓ�q@��������Dr��	ך�Q;��6������>f���ɡ��,�����}�W���������Ă��笼@K����������w���۳��?��~���$���j��kκ�)2��:����  �  n�N=�N=P_M=S�L=�K=NEK=4�J=��I=�'I=�rH=)�G=FG=QF=v�E=��D=4,D=�tC=F�B=�B=gJA=��@=
�?=�?=�^>=��==��<=%<=Te;=��:=��9=�9=�[8=�7=��6=+	6=m@5=>v4=��3=O�2=C2=F=1=j0=Ɣ/=ݼ.=b�-=-=�$,=A+=,Z*=�o)=t�(=\�'=�&=��%=��$=֛#=1�"=l�!=7r =XY=�:=�=��=
�=��=>A=��=,�=JX=2�=Ƙ=*.=^�=�C=��=1=
=�=�=��=��=?==� =���<�V�<��<�a�<K��<$H�<֮�<��<Le�<��<� �<4E�<R��<���<K��<�%�<hS�<�}�<���<yȷ<��<��<%�<[?�<�W�<Jn�<��<���<���<㹐<ʌ<�و<	�<0��<�z<�-r<�Mj<�nb<�Z<�R<�J<�C<�3;<�b3<G�+<Y�#<�<�=<�}< �<��;��;�[�;��;iԼ;���;���;3��;ӈ�;�Lc;�E;.I(;�;��:L�:�R:���9�Ao�tj�� Xl�7���v}����.&�h�?���Y�<�r�뮅�ב��ɝ�I������|R���d˻�>ֻ���xI�{��`v������e	���L��$�F��H���$��&(�0,�%0�S4�.�7���;��>?���B�riF���I�]M�5�P�] T��qW�]�Z�^�]��,a��Yd�Y~g���j�M�m�Y�p���s���v���y�Z�|�E��2N�����5������x��너�]��^��uʌ�:5��F������3q��1ٓ�M@��⦖����&r���֚�=;��0������.f��dɡ��,�����k�W��ں�����؂��)笼PK����������w��ܳ��?������B���j���κ�:2��[����  �  w�N=
N=]_M=U�L=��K=EEK=.�J=��I=�'I=�rH=$�G==G=�PF=f�E=u�D=$,D=ltC=B�B=�B=ZJA=��@=��?=�?=�^>=��==��<=(%<=ee;=��:=��9=�9=\8=�7=��6=>	6=z@5=Tv4=��3=`�2=M2=O=1=.j0=Δ/=�.=m�-=	-=�$,=A+=&Z*=�o)=k�(=K�'=�&=��%=�$=ƛ#=!�"=V�!=*r =[Y=�:=�=��=�=��=7A=��=6�=\X=?�=ט=9.=n�=�C=��=L=
='�=�=Ђ=��=X==� =���<�V�</��<�a�<Z��<'H�<Ʈ�<��<9e�<	��<� �<%E�<S��<���<)��<�%�<JS�<s}�<l��<pȷ<��<|�<�$�<K?�<�W�<4n�<��<���<Ѩ�<���<-ʌ<�و< �<J��<�z<�-r<�Mj<Lob<I�Z<@�R<M�J<�C<�3;<�b3<��+<��#<�<�=<�}<��<��;Ӳ�;_[�;��;Լ;���;��;}�;9��;gKc;��E;}H(;�;��:�|�:دR:$��9aio��k���Ul������|�����&�v�?�9�Y�Z�r�o����֑��ȝ����L��AR��td˻P>ֻ����H��z��Wv��ŝ��e	������:$����H��-$��&(�^0,�R%0��4�f�7�z�;��>?���B��iF���I�]M�[�P�S T��qW� �Z�9�]��,a�VYd�,~g�N�j�-�m���p�C�s�J�v�n�y�9�|����N����m5������^��儈�b��^��zʌ�T5��]������Eq��3ٓ�q@��������Dr��	ך�Q;��6������>f���ɡ��,�����}�W���������Ă��笼@K����������w���۳��?��~���$���j��kκ�)2��:����  �  ��N=N=a_M=\�L=��K=9EK="�J=��I=�'I=rH=�G=G=�PF=0�E=6�D=�+D=.tC=�B=bB=.JA=f�@=��?=�?=�^>=¡==��<=2%<=xe;=��:=��9=! 9=9\8=&�7=��6={	6=�@5=�v4=ߪ3=��2=~2=v=1=Tj0=ߔ/=��.=p�-=-=�$,=A+=Z*=�o)=N�(=�'=ߘ&=L�%=D�$=��#=�"=�!=�q =+Y=u:=�=��=��=��=6A=��=@�=rX=Z�=�=i.=��=�C=�=�=
=k�=�=�=?�=�==J� =0��<KW�<p��<b�<s��<HH�<Į�<��<e�<ܵ�<8 �<�D�<��<��<���<'%�<�R�<�|�<���<ȷ<H�<=�<�$�<$?�<�W�<,n�<&��<���<ꨔ<��<~ʌ<6ڈ<��<���<�z</r<�Nj<hpb<F�Z</�R<B�J<�C<�4;<Fc3<��+<��#<�<�=<}}<��<�;���;�Y�;�;DҼ;���;8��;N}�;N��;�Fc;��E;~D(;3;��:�w�:E�R:n��9dzo�"o���Ul������z�
���&�x�?�I~Y���r�����>Ց�ǝ���������P��^c˻F=ֻ�໠H��z��!v����f	�N����$�v����%	$��'(�C1,�<&0��4�_�7�I�;��??�:�B�&jF�1�I�O]M�z�P�2 T��qW��Z���]��+a��Xd�r}g�c�j�V�m��p�b�s�^�v�n�y�_�|����M��Z�65��q���D������T��^���ʌ��5������	���q���ٓ��@��t���m���r���ך��;������<��uf���ɡ��,��(���~�W��������������欼�J��&���Q��vw��^۳�Y?���������Oj���ͺ��1��啽��  �  ��N=AN=y_M=a�L=��K=EK=��J=n�I=�'I=CrH=��G=�G=lPF=ԙE=��D=�+D=�sC=��B=B=�IA=*�@=��?=�?=�^>=��==��<=L%<=�e;=�:=4�9=g 9=�\8={�7=F�6=�	6=A5=�v4=9�3=��2=�2=�=1=�j0=�/= �.=��-=-=�$,=�@+=�Y*=Wo)=�(=ڎ'=��&=��%=�$=6�#=��"=̈́!=�q =�X=>:=�=o�=׸=t�=5A=��=[�=�X=��=F�=�.= �=7D=~�=�=
=�=P=��=��=�==�� =���<�W�<���<]b�<���<ZH�<���<n�<�d�<y��<���<ED�<V��<n��<��<s$�<R�<H|�<J��<cǷ<��<��<G$�<�>�<CW�<n�<&��<Ȗ�<+��<|��<�ʌ<�ڈ<&�<d��<Qz<�0r<�Pj<�qb<��Z<��R<��J<�	C<�5;<=d3<��+<1�#<<�=<!}</�<��;���;�W�;��;�ϼ;Ρ�;��;6z�;��;Ac;��E;4?(;\;k�:�p�:ӜR:V��92�o�nr��Sl�A����u�Y���&���?��yY�m�r�%���iґ��ĝ����z���N���a˻�;ֻ��໴G�lz��=v�����f	������%�m��]��{
$�@)(��2,��'0��4���7���;��@?�;�B��jF���I��]M���P�; T�WqW�g�Z�2�]�*+a��Wd�M|g�>�j��m���p���s���v�'�y��|���1M�������4�����
��˄��^�_���ʌ��5��
���~	��7r��=ړ��A��$��� ��js��+ؚ�g<��4�������f�� ʡ�.-��c������V������L��6���I欼jJ����������v���ڳ��>��K������i��fͺ�P1��w����  �   �N=kN=�_M=h�L=��K=EK=ҐJ=9�I=:'I=�qH=@�G=HG=�OF=Y�E=n�D=+D=ksC=O�B=�B=�IA=�@=��?=d?=}^>=��==�<=n%<=�e;=5�:=��9=� 9=�\8=�7=��6=P
6=�A5=\w4=��3=R�2=+2=>1=�j0=J�/=C�.=��-=-=�$,=�@+=�Y*=o)=��(=�'=(�&=��%=~�$=Ś#=!�"=X�!=9q =|X=�9=6=:�=��=b�=6A=��=��=�X=��=��=/=y�=�D=�=�>
=u�=�=�=8�=w>= � =���<�X�<o��<�b�<���<qH�<®�<C�<�d�<��<4��<�C�<���<���<��<�#�<&Q�<U{�<h��<�Ʒ<
�<�<�#�<m>�<W�<�m�<��<���<u��<�<vˌ<qۈ<��<H��<Vz<`2r<�Rj<�sb<ʖZ<��R<?�J<lC<�6;<`e3<u�+<��#<P<�=<�|<��<�;w��;�T�;(	�;�˼;ޝ�;р�;Fv�;�~�;�8c;��E;�7(;� ;���:Xh�:0�R:C��9>p�u��Ol�����Fo⺕���&�5�?�sY���r�Ŧ���Α�w���q|��e ���K��_˻�9ֻ(���F��y���v��U��'g	���ߪ�'�����2$�,+(��4,��)0��
4�i�7�?�;�FB?���B��kF�z�I�V^M���P�K T��pW��Z�^�]�*a�oVd��zg���j��m��p���s���v�O�y�$�|�S��jL��G���@4�������������i�._��#ˌ�.6������'
�� s��ۓ�qB�������^t��ٚ�>=�����d���g���ʡ��-���������V��S�����������嬼�I��̭������u���ٳ��=��f������h���̺��0��唽��  �  C�N=�N=�_M=v�L=��K=�DK=��J=��I=�&I=�qH=ͻG=�G=sOF=јE=��D=�*D=�rC=ԺB=DB=:IA=��@==�?=3?=c^>=��==�<=�%<=	f;=}�:=��9=/!9=_]8=m�7=I�6=�
6=B5=�w4=4�3=��2=�2=n>1=%k0=��/=n�.=��-=-=�$,=�@+=�Y*=�n)=k�(=�'=��&=�%=��$=?�#=��"=փ!=�p =X=}9=�=��=}�=K�=0A= �=��=Y=3�=�=�/=��=IE=��=1?
=�=�=��=��=	?=�� =~��<[Y�<��<:c�<;��<�H�<���<�<!d�<~��<���<�B�<���<���<��<m"�<P�<Az�<c��<�ŷ<"�<R�<"#�<�=�<�V�<�m�<0��<#��<Ω�<r��<(̌<;܈<��<G��<~z<�4r<�Tj<3vb<�Z<��R<?�J<1C<�8;<�f3<h�+<\�#<�<�=<�|<��<��;٪�;�Q�;U�;�Ǽ;S��;|�;-q�;�y�;n/c;��E;/(;W�
;��:\�:|R:�o�9��p�;x���Ll�����h����&���?�alY��r�Ѣ���ʑ�K����x�������H��Y\˻g7ֻS�໮E�fy��nv������g	���-���(�������9$�W-(��6,��+0�4�u�7�"�;�D?���B�:mF���I��^M�)�P�9 T��pW�C�Z�[�]��(a��Td�yg���j��m���p���s���v��y�5�|�v���K�������3��A����������g�\_��~ˌ��6��2����
���s��
ܓ�yC��/���$��mu��#ښ�:>��록�=��9h��'ˡ��-��ʐ�����V��!������8���嬼�H��謯�����t���س�|<��F������g���˺��/��1����  �  ��N=�N=�_M=��L=��K=�DK=j�J=��I=�&I=qH=V�G=@G=�NF==�E=@�D=�)D=TrC=O�B=�B=�HA=7�@=��?=?=@^>=��==&�<=�%<=Cf;=å:=@�9=�!9=�]8=��7=��6=v6=�B5=�x4=��3=X�2=2=�>1=xk0=̕/=��.=��-= -=j$,=�@+=LY*=}n)=�(=��'==�&=��%=n�$=��#=�"=M�!=4p =�W=9=�=��=M�=1�=$A=�=ͭ=RY=��=j�=0=��=�E=I�=�?
=Ȳ===e�=t�=�?=/� =���<Z�<���<�c�<���<�H�<���<��<�c�<��<���<�A�<���<t��<���<4!�<�N�<y�<;��<�ķ<5�<}�<u"�<o=�<dV�<�m�<4��<Q��<7��<�<�̌<݈<��<e��<�z<>7r<VWj<�xb<l�Z<�R<w�J<C<,:;<�g3<x�+<��#<�<v=<�{<��<=�;���;�M�;[�;�¼;P��;�v�;�k�;�t�;�$c;�E;i&(;��
;t��:8P�:{jR:�Q�9)q��|��IIl������b�����&�n�?��dY��r�q����Ƒ�򸝻�t������PE��IY˻5ֻ���CD��x��yv��5��zh	������.*��������$��/(�@9,�7.0�S4���7��;��E?���B��nF���I��_M���P�8 T�_pW�|�Z�j�]��'a�LSd�:wg���j��m�K�p�o�s�k�v�սy��|�R���J������3��Τ��0��e���u򉼞_���ˌ�E7��塏�����t��ݓ��D��O���[���v��Eۚ�V?��ܢ�����h���ˡ�`.��������V��깨�-������T䬼H��髯�����s���׳�Z;���������f���ʺ��.��w����  �  ��N=	N=�_M=��L=��K=�DK=0�J=\�I=*&I=�pH=ӺG=�G=TNF=��E=��D=e)D=�qC=ƹB=SB=cHA=ߎ@=��?=�?=%^>=��===�<=�%<=zf;=�:=��9="9=_^8=��7=i�6=6=LC5=y4=O�3=��2=�2=D?1=�k0=�/=ν.=��-=&-=[$,=c@+=Y*=8n)=�(=5�'=��&=�%=�$=�#=t�"=��!=�o =W=�8=-=m�=�=�=!A=%�=��=�Y=��=ؚ=�0=�=�F=��=�@
=��=�=�="�=E@=�� =���<�Z�<d��<9d�<���<�H�<���<��<Xc�<S��<��<�@�<��<i��<���< �<�M�<�w�< ��<}÷<L�<��<�!�<�<�<V�<qm�<?��<���<���<~��<�͌<�݈<��<}��<+z<�9r<�Yj<9{b<�Z<I�R<~�J<�C<�;;<(i3<e�+<��#<B<^=<�{<�<�;���;HJ�;���;M��;z��;�q�;�f�;Zo�;�c;�E;(;��
;o��:E�:�VR:�8�93�q�Q|��El�V���[�����%���?��\Y��{r�"���B�״���p��;���B��:V˻�2ֻ���3C�x��~v�����;i	�������+�]��'���$��1(��;,��00��4���7�E�;��G?�@�B��oF�{�I�U`M���P�2 T��oW�ڵZ�q�]�:&a��Qd�yug���j���m��p���s��v���y�ʲ|�i���I������u2��[������/������_��>̌��7����������u��ޓ��E��~�������w��bܚ�g@��裝�����i��N̡��.��]����󥼳V���������%����㬼=G���������r��Zֳ� :��흶�����e���ɺ�.�������  �  �N==N=`M=��L=��K=�DK=��J=�I=�%I=CpH=^�G=<G=�MF=�E=$�D=�(D=HqC=J�B=� B= HA=��@=u�?=�?=^>=��==I�<=�%<=�f;=a�:=��9={"9=�^8=�7=��6=�6=�C5=�y4=ԭ3=Q�2=�2=�?1= l0=V�/=��.=�-=%-=K$,=?@+=�X*=�m)=F(=Ќ'=C�&=��%=V�$=��#=�"=4�!==o =�V=K8=�=&�=�=�=A=0�=$�=�Y=2�=<�=1=��=G=��=/A
=&�=� =��=��=�@=A� =^��<�[�<��<�d�</��<�H�<���<P�<�b�<���<W��<)@�<�~�<p��<���<��<�L�<�v�< ��<�·<u�<��<@!�<o<�<�U�<Gm�<?��<���<<��<7Ό<�ވ<��<}��<Uz<�;r<[\j<�}b<!�Z<d�R<t�J<�C<D=;<~j3<Y�+<>�#<x<4=<{<D�<��;���;�F�;��;��;؊�;�l�;�a�;Bj�;�c;{E;�(;L�
;���::�:�ER:8"�9�.r�����Bl�4����S�λ��%���?��UY�2tr�F���!���ܰ���l�����>���S˻[0ֻ���B뻊w���v�����i	���	��]-������$�64(��=,��20��4���7�0�;�TI?���B�qF��I��`M�0�P�F T��oW�>�Z�W�]��$a�KPd��sg���j���m��p�̺s��v�w�y�Ұ|�����H��L����1��ۣ�����������_���̌�H8��9���P���v��ߓ��F����������x��uݚ�^A��֤�����yj���̡�D/����������V��m���l������⬼uF���������q��Hճ��8��ܜ��� ���d���Ⱥ�I-������  �  R�N=fN=#`M=��L=��K=oDK=яJ=��I=�%I=�oH=��G=�G=RMF=��E=��D=c(D=�pC=ݸB=� B=�GA=?�@=9�?=y?=�]>=��==S�<=&<=�f;=��:=F�9=�"9=<_8=p�7=g�6=6=MD5=z4=C�3=��2=[2=�?1=dl0=��/=�.=�-=+-=7$,=@+=�X*=�m)=�~(=n�'=ݕ&=�%=�$=�#=z�"=ǁ!=�n =AV=�7=�=��=��=�=A=B�=>�=�Y=o�=��=l1=�=�G=�=�A
=��="!=A�=<�=TA=�� =)��<\\�<���<�d�<g��<I�<l��<�<�b�<A��<���<o?�<�}�<{��<���<��<�K�<�u�<,��<���<��<D�<� �<	<�<zU�<%m�<I��<՗�<9��<t��<�Ό<h߈<��<a��<.z<�=r<7^j<�b<�Z<C�R<7�J<;C<�>;<qk3<�+<��#<�<!=<�z<��<��;D��;�C�;���;5��;���;�h�;g]�;?f�;�c;"sE;s(;��
;S��:L0�:	7R:�
�9�wr�\����@l�����N�ķ�\�%���?��OY�qmr�Ӓ��ẑ�D����i����;��4Q˻s.ֻ���#A�Mw���v��I��sj	���0���.��������$�6(��?,��40��4���7�ܟ;��J?��B�+rF�R�I�zaM���P�8 T�goW�ǴZ���]��#a��Nd�-rg���j��m���p��s��v���y�$�|���GH������d1������n��������.`���̌��8��ǣ����aw���ߓ��G����������y��gޚ�JB���������k��a͡��/��ܑ��2����V��P�����,��g⬼�E��P�������p��PԳ�8��盶������c��Ⱥ��,������  �  z�N=�N=<`M=��L=��K=VDK=��J=��I=O%I=�oH=��G=vG=�LF=I�E=@�D=(D=rpC=��B=6 B=fGA=	�@=�?=V?=�]>=��==Z�<=.&<=g;=Ʀ:=��9=#9=�_8=7=��6=k6=�D5=qz4=��3=�2=�2=3@1=�l0=��/=B�.=�-=/-=,$,=@+=|X*=sm)=�~(='�'=��&=��%=��$=��#=�"=y�!=tn =�U=�7=W=��=��=�=A=O�=T�=&Z=��=ћ=�1=]�=�G=u�=$B
=�=�!=��=��=�A=�� =���<�\�<���<We�<���<I�<Z��<��<;b�<��<@��<�>�<N}�<ɶ�<��<1�<�J�<4u�<~��<��<�<��<: �<�;�<@U�<m�<N��<���<���<ý�<Gό<�߈<��<	 �<�z<x?r<�_j<�b<m�Z<��R<y�J<IC<�?;<+l3<Û+<�#<�<=<Iz<��<�;r��;�A�;6��;g��;ƃ�;�e�;�Y�;9c�;vc;dmE;�(;��
;ӱ�:�'�:�*R:p��9��r�2����;l�Â��!J�P��8�%���?�BKY��hr�'���B���Ī��Gg��;촻:��jO˻�,ֻ}��@��v���v������j	�U����/�͔����
$�\7(�QA,�D60�4�;�7��;�L?��B��rF��I��aM���P�, T�;oW�6�Z��]�&#a��Md�8qg�Ìj���m���p���s���v�K�y�֭|�����G��(���1��<���*��냈���S`��#͌�9��1�������w������]H��*���X���z��ߚ��B��1���	��k���͡��/�����B����V��%�������~���ᬼSE��¨��J���o���ӳ�m7��/���3���5c���Ǻ�&,������  �  ��N=�N=H`M=��L=��K=QDK=��J=��I=$%I=xoH=y�G=@G=�LF=�E=	�D=�'D=;pC=T�B= B==GA=��@=��?=H?=�]>=��==\�<=;&<=g;=�:=��9=D#9=�_8=��7=��6=�6=�D5=�z4=Ԯ3=C�2=�2=Z@1=�l0=/=O�.='�-=(-=*$,=�?+=hX*=Vm)=�~(=��'=^�&=��%=V�$=��#=�"=9�!=An =�U=�7=4=��=��=�=A=M�=d�=<Z=��=��=�1=��=0H=��=hB
=`�=�!=�=��=�A==� =��<)]�<&��<�e�<���<I�<a��<��<"b�<���<���<�>�<�|�<`��<���<��<aJ�<�t�<��<���<��<w�< �<�;�<-U�<m�<?��<��<���<���<~ό<F��<���<z �<� z<Y@r<�`j<��b<|�Z<��R<T�J<C<#@;<�l3< �+<G�#<�<�<<5z<��<b�;��;'@�;V��;���;Á�;vc�;�W�;�`�;�b;CiE;(;��
;���:�$�:O%R:��9*�r�����:l�����!G���@�%���?��GY�,er�����t������je���괻Z8��GN˻ ,ֻ����?뻿v�� w�����5k	������F0�}������$�c8(�=B,�*70�4��7��;��L?���B��sF�[�I�3bM���P�M T�oW���Z���]��"a�pMd�Xpg���j���m�®p���s���v�T�y��|���aG�����0�������ト���X`��>͌�A9��������[x�������H���������{���ߚ�_C������_	���k���͡�0�����L����V���������~���ᬼ�D��X�������o��0ӳ��6��Ú�������b��Ǻ��+��͐���  �  ��N=�N=hM=M�L=-L=�NK=��J=��I=�1I=+}H=�G=�G=W]F=��E=��D=<D=�C={�B=�B=�aA=�@=��?=�8?=f>=��==�	==sM<=5�;=��:=�:=cR9=��8=d�7=�
7=�E6=X5=��4=f�3={#3=�V2=,�1=m�0=f�/=�/=�6.=�[-=�},=x�+=�*=��)=�(=r�'=� '=�&=�%=�$=5#=p�!=Q� =��=�=�=�o=�@=�
=a�=��=�<=��=y�=f*=��=qM=��=�R=m�
==;	=?�=�=�e=ϼ=�=���<�>�<���<t8�<ئ�<v�<�i�<���<�<lT�<���<���<.�<�8�<2f�<׏�<��<Nٿ<���<��<=3�<�L�<�c�<:y�<֌�<���<�<ν�<U˔<�א<!�<��<+��<�<�z<�+r< @j<RUb<*lZ<=�R<A�J<+�B</�:<��2<�+<�A#<�j<ߖ<��<��<g�;���;�j�;$��;A��;�U�;e�;.�;˼{;��];��?;ZV";��;�q�:�{�:��7:��9�;,�����℺ ������ ��l.�� H�
�a��{����+��!,��h�ہ����Ļ'�ϻ��ڻ/u廃����~�U��Ӭ�TW�J��b]�����!�*&��>*�=.��%2� �5�ߺ9�.i=�A� �D��H���K���N��:R���U���X�� \�/0_�;Wb�ive��h���k���n�4�q�˩t��w���z���}�D6��)���a������K���he���ш��<������t���z���⏼�J���������$}���ᖼE��ͧ���	���j��h˝�w+��O����꡼oJ������	���i��1ʨ��*��拫�2��N��K���"���s��ֳ��7��������_^�������#��Æ���  �  ��N=tN=hM=M�L=,L=�NK=њJ=��I=2I=6}H='�G=�G=t]F=ۧE=�D='<D=��C=��B=�B=�aA=�@=��?=9?=g>=��==�	==fM<=*�;=��:=�:=LR9=ܐ8=A�7=�
7=�E6=;5=��4=D�3=d#3=�V2=�1=k�0=[�/=�/=�6.=�[-=�},=�+=�*=��)=�(=}�'=� '=	&=�%=$=T#=��!=n� =��=��= �=�o=�@=�
=Z�=��=�<=��=j�=_*=��=WM=��=�R=I�
=;	=�=�=�e=��=�=���<�>�<i��<K8�<Ʀ�<i�<�i�<��<,�<T�<���<
��<b�<9�<of�<��<[��<�ٿ<���<��<Y3�<�L�<d�<ey�<猤<���<���<���<@˔<�א<#�<��< ��<��<Qz<!+r<�?j<�Tb<�kZ<��R<؝J<йB< �:<��2<�+<�A#<�j<ϖ<��<��<fg�;C��;�j�;���;9��;�V�;x�;,�;��{;��];�?;�W";�;ft�:"~�:��7:�904,�D���ㄺ����������~.�%"H���a��{�;����,���,��_���������Ļz�ϻ��ڻuu����K��e�]�����W���]�Ź���!��)&�O>*��<.�]%2���5�g�9��h=��A���D��H���K�|�N��:R���U���X�� \�X0_�DWb��ve�R�h��k��n���q�A�t�T�w�4�z�N�}�q6��S���k�����_����e���ш��<������J��qz���⏼�J����������|��Tᖼ�D������t	���j��=˝�`+��+����꡼KJ�������	���i��Gʨ��*������3��N��w���Y��:t��0ֳ�"8��6���U����^�������#��Æ���  �  `�N=`N=�gM=M�L=6L=�NK=�J=��I=A2I=s}H=j�G=,G=�]F='�E=`�D=s<D=E�C=��B=B=�aA=J�@=�?=$9?=r>=��==�	==TM<=�;=��:=w:=R9=��8=�7=A
7=@E6=�~5=;�4=��3=&#3=~V2=�1=9�0=7�/=�/=�6.=�[-=�},=��+=�*=�)=U�(=��'=$'=S	&=%=I$=�#=��!=�� =��=5�=Y�=�o=�@=�
=^�=��=�<=��==�= *=[�=
M=J�=0R=��
=�:	=Ť=>=[e=f�=�=��<:>�<��<	8�<���<\�<�i�<;��<^�<�T�<��<���<��<�9�<g�<���<���<ڿ<���<b�<�3�<1M�<Xd�<�y�<��<Ӟ�<��<���<˔<Wא<��<N�<���<U�<2z<�)r<?>j<�Sb<njZ<��R<J<��B<5�:<��2<@+<@A#<uj<�<�<j�<{h�;��;�l�;��;���;�X�;�;���;b�{;��];7�?;p\";��;�|�:��:N8:���9\,����䄺1�����񺙱��.�0%H�.�a�+{�8����.���.��L���<���W�Ļ,�ϻ2�ڻnv�x��u��C�!��F���V�\��\�Ǹ���!�z(&�*=*�e;.�4$2���5�K�9��g=��A�ÑD��H��K��N��:R���U���X�4\��0_�Xb�wwe�Q�h��k��n���q�z�t�x�w�>�z�L�}��6��ѩ�����e��������e���ш��<��p�����-z��|⏼J�������b|������HD���������j���ʝ��*������v꡼J��Щ���	���i��aʨ�+��I�����DO����������t���ֳ��8����������_��x���6$��*����  �  )�N=6N=�gM=A�L=CL=�NK=�J=��I=�2I=�}H=��G=�G=9^F=��E=��D=�<D=C=I�B=�B=IbA=��@=D�?=G9?=�>=�==�	==9M<=�;=��:=):=�Q9=3�8=��7=�	7=�D6=p~5=��4=��3=�"3= V2=��1=�0=�/=�/=�6.=�[-=�},=��+=B�*=G�)=��(=�'=�'=�	&=�%=�$=#=M�!=$� =M�=��=��=*p=�@=�
=p�=��=c<=��=��=�)=��=�L=��=�Q=`�
=(:	=.�=�=�d=޻==D��<�=�<���<�7�<]��<;�<�i�<^��<��<JU�<���<K��<��<z:�<�g�<���<���<$ۿ<|��<=�<�4�<�M�<�d�<z�<p��<��<���<���<�ʔ<�֐<.�<��<���<l �<Hz<�'r<<<j<�Qb<lhZ<��R<��J<X�B<��:<��2<q+<�@#<#j< �<��<�<�j�;Q��;�o�;e�;[��;<]�;h"�;_��;2�{;��];@;Pd";h�;���:���:r8:H�9,�[��儺o���]��f���.�+H�9�a��{�����^2��m2������������ĻC�ϻ-�ڻ�w�[�����W��������U�B���Z�����!��&&�#;*�Z9.�("2�}�5�`�9�f=�;A���D��H�K���N�:R���U���X��\��1_� Yb��xe���h�ˡk�߫n���q�i�t�r�w�+�z��}��7��x���s��䊄������e���ш��<��&�������y���ᏼwI��9���F��i{���ߖ�GC���������0i���ɝ�#*��&����顼�I�������	���i���ʨ�q+������-�O����������u���׳��9��Û�������_��Fº��$��Ç���  �  ��N=�N=�gM=<�L=KL=OK=Q�J=V�I=�2I=J~H=X�G=1G=�^F=A�E=��D=�=D=`�C=��B=B=�bA=�@=��?={9?=�>=�==�	==M<=��;=8�:=�:=HQ9=��8=�7=)	7= D6=�}5=�4=��3=)"3=�U2=&�1=��0=��/=i/=�6.=�[-=�},=ݜ+=��*=��)=�(=��'='=]
&=-%=_$=�#=��!=�� =��=�=��=}p=5A=�
=x�=��=?<=:�=��=Z)=r�=L=�=�P=��
=p9	=q�=�=%d=6�=�=1��<�<�<о�<7�<��<�<�i�<���<@�<�U�<r��<@��<�	�<�;�<.i�<���<9��<hܿ<���<]�<�5�<�N�<�e�<�z�<ȍ�<.��< ��<e��<aʔ<g֐<h�<��<���<H��<�z<=%r<�9j<�Nb<�eZ<M~R<��J<Q�B<�:<m�2<=+<'@#<�i<�<��<��<dm�;���;�s�;�	�;U��;�b�;�'�; �;�{;�];�@;En";X;���:���:))8: 0�9��+�2���愺˺����񺡺��$.�t2H��a��"{�W����6���6������}�����Ļ��ϻ��ڻ�y����7��H�<������T����1Y�����!�"$&��8*��6.��2��5��9��c=�:A�ߎD�OH��}K���N��9R���U�9�X��\��2_�~Zb�dze���h��k�#�n�4�q�үt��w���z�H�}��8��d���L������x���:f���ш��<��馋�p��y��3ᏼ�H��2���(��0z���ޖ�B���������h���ȝ�-)��\���5顼?I��B����	���i���ʨ��+��C�����P����������v���س��:���������a��Mú��%�������  �  ��N=�N=�gM=1�L=bL=2OK=��J=��I=c3I=�~H=��G=�G=�_F= �E=F�D=I>D=�C=��B=�B=DcA=`�@=��?=�9?=�>=�==x	==�L<=a�;=��:=J:=�P9=�8=W�7=v7=eC6=}5=h�4=E�3=�!3=U2=��1=)�0=q�/=2/=^6.=�[-=�},=�+=˸*=�)=��(= �'=�'=&=�%=$=k#=��!=]� =q�=��=w�=�p=qA==|�=��=<=��=>�=�(=ֽ=UK=d�=&P=��
=�8	=��==Rc={�=�=���<�;�<��<{6�<���<�<�i�<���<��<�V�<f��<N��<�<=�<�j�<z��<���<�ݿ<��<��<�6�<�O�<}f�<D{�<B��<p��<��< ��<�ɔ<�Ր<���<��<{�<���<�z<>"r<j6j<�Kb<�bZ<x{R<�J<�B<�:<��2<+<C?#<�i<A�<��<��<p�;j��;qx�;%�;&��;�h�;Z.�;��;��{;��];4@;wy";�;e��:[��:B8:Q�9�+����c鄺����%��y��},.��:H���a��,{����a<��<�����������Ļ,�ϻ��ڻ�{�\�����������US�#��W����!�[!&��5*��3.��2��5�/�9�'a=��@���D��H��|K���N�E9R���U���X�a\��3_�\b�`|e��h�V�k��n���q��t��w�q�z��}�
:������>��K�������f��҈��<���������ux��]����G���������x��ݖ��@��?���F���f���ǝ�(��a����衼�H��ۨ��P	��j��˨�b,����לּ�Q��鳯���Bx��hڳ�{<��t���a ��ab��yĺ��&��k����  �   �N=yN=ugM=#�L=pL=ZOK=�J=�I=�3I=eH=��G=�G=K`F=ΪE=�D=?D=ˈC=8�B=?B=�cA=ݫ@=I�?=:?=�>=#�==a	==�L<=�;=n�:=�:=P9=i�8=��7=�7=�B6=I|5=��4=��3=� 3=hT2=!�1=��0=�/=�/=66.=�[-=~,=K�+=#�*=n�)=�(=��'=]'=�&=�%=�$=.	#=X�!=� =�=�=��=5q=�A===��=q�=�;=��=ɋ=G(=8�=�J=��=@O=��
=�7	=��=0=lb=��==ĭ�<�:�<$��<�5�<B��<��<�i�<Z��<P�<wW�<k��<~��<c�<k>�<Cl�<
��<_��<o߿<���<�<8�<�P�<eg�<|�<���<���<���<ۼ�<�ɔ<Ր<�ߌ<��<$�<y��<�z<r<3j<�Hb<�_Z<OxR<:�J<b�B<��:<��2<�+<m>#<9i<Y�<+�<6�<As�;���;A}�;��;)��;Mo�;q5�;��;�{;*�];&@;��";�; ��:���:0]8:Tq�9�+����.넺�Ż�V��X���4.��CH�I�a��7{�3
��B���A�����.�����Ļ��ϻ�ڻi~建�������P������Q�O���T�g��C�!��&��2*��0.�d2���5�\�9�e^=���@���D��	H�Y{K���N��8R���U�:�X�#\�:5_��]b�[~e��h��k��n���q���t���w�v�z�	�}�c;��í��.��&��������f��Q҈��<��s���]���w��mߏ�fF��ά��j��aw��tۖ��>���������Ee��EƝ��&��P����硼H������1	��j��a˨��,���������R��8�������y���۳�
>����������c���ź��'��V����  �  ��N=(N=NgM=�L=�L=�OK=-�J=w�I=`4I=�H=F�G=KG=aF=��E=��D=�?D=��C=��B=�B=`dA=Q�@=��?=E:?="�>=+�==O	==�L<=��;=�:=J:=�O9=��8=��7=�7=�A6=�{5=ڳ4=��3=' 3=�S2=��1=>�0=��/=�/=6.=�[-=,~,=w�+=u�*=��)=��(=R�'='=r&=c%=�$=�	#=�!=�� =��=��=d�=�q=B=Z=��=X�=�;=L�=R�=�'=��=�I=��=iN=��
=�6	=��=C=�a=ڸ=O
=j��<m9�<2��<B5�<ޤ�<��<j�<���<��<AX�<_��<���<��<�?�<�m�<���<��<�<�<{�<W9�<�Q�<Oh�<�|�<��<ܟ�<���<���<�Ȕ<?Ԑ<�ތ<x�<��<
��<�z<�r<�/j<)Eb<D\Z<HuR<f�J<ۭB<��:<,�2<i+<�=#<�h<|�<��<8 <�v�;���;��;W�;v��;�u�;*<�;��;�|;=^;R3@;�";W";���:�ʕ:�s8:#��9Lg+����i턺"ͻ�p	�_��l<.�MH�*�a��B{����G���G�����M���A�Ļлv�ڻ�廍�ﻐ�������/��pP�����R�ڭ�}�!�p&�w/*�x-.�E2���5�G�9��[=��@���D�*H��yK�9�N�M8R���U���X�\��6_��_b���e���h�۫k�Ѷn�/�q��t�$�w���z�ѐ}��<��󮁼C�����W���]g��|҈��<��$�������v���ޏ�YE���������u���ٖ�d=�����7���c���ĝ��%��c����桼qG��,���	��3j���˨�t-��z�����T��������G{���ݳ��?������l��8e��Ǻ�)��_����  �  i�N=�N="gM= �L=�L=�OK=j�J=��I=�4I=��H=��G=�G=�aF=H�E=��D=�@D=D�C=��B=yB=�dA=��@=��?=}:?=J�>=.�==8	==RL<=u�;=��:=�:= O9=�8=8�7=97=A6=�z5=�4=�3=y3=9S2=
�1=մ0=f�/=u/=�5.=�[-=@~,=��+=��*=:�)=��(=��'=�'=&=%=V$=�
#=��!=k� =K�=;�=֚=�q=<B=}=��=8�=o;=��=�=7'=�=)I=��=�M=�
=�5	=՟=h=�`=�=�	=#��<v8�<f��<�4�<~��<w�<1j�<���<h�<�X�<K��<���<��<OA�<'o�<-��<h��<q�<~�<��<�:�<�R�<i�<=}�<���<��<߮�<_��<qȔ<�Ӑ<�݌<d�<���<���<�z<�r<�,j<�Ab<HYZ<[rR<��J<�B<��:<��2<+<�<#<gh<��<o�<-<my�;:��;���;_�;%ƺ;|�;�B�;��;�|;^;"?@;�";w,;���:�ؕ:�8:(��9�G+��������ӻ�������C.�&VH��b�=M{����^M�� M����Y���_�Ļ�лt�ڻ/��^��/���G��M��BO�����P�}���!��&��,*�q*.�12��5�r�9�/Y=���@���D��H��xK�f�N��7R�ĆU��X�\��7_�Eab���e�!�h���k���n�#�q��t�"�w�z�z���}�>�����J �����������g���҈��<��ݥ�����Zv���ݏ�VD��\������nt���ؖ��;������� ��tb���Ý��$��|���&桼�F��˧�����Yj���˨� .�������U������C���|��߳�A���������f��MȺ�"*��K����  �  �N=�N=gM=��L=�L=�OK=��J=�I=55I=��H=a�G=�G=]bF=�E=2�D=-AD=ڊC=�B=�B=WeA= �@=F�?=�:?=_�>=2�==*	==-L<=7�;=M�:=d:=�N9=��8=��7=�7=w@6=z5=��4=~�3=�3=�R2=��1=t�0=�/=E/=�5.=�[-=M~,=֝+=��*=��)=h�(=V�'=!'=�&=�%=�$=>#=S "=�� =��=��=<�=9r=rB=�=��=&�=C;=��=��=�&=c�=�H=N�=�L=h�
=5	=�=�=`=l�=	=��<�7�<���<4�<0��<U�<3j�<<��<��<�Y�<��<���<��<sB�<dp�<_��<���<��<��<� �<�;�<�S�<�i�<�}�<ߏ�<*��<ᮜ<)��<Ȕ<�Ґ<�܌<s�<��<u��<z<�r<�)j<a?b<�VZ<�oR<l�J<i�B<��:<�2<+<)<#<3h<��<��<3<�{�;���;���;�#�;�ʺ;b��;H�;� �;�|;�^;ZI@;�";5;3��:	�:|�8:�͌9B-+������6ػ���4��WJ.��]H�Zb�!V{���R���Q�����~���+�Ļ:
л5�ڻn�廣���������z��N����O������!�O&�**��'.��2���5�(�9�W=���@�ЄD�2H��wK���N��7R�ÆU�g�X��\� 9_��bb�a�e�"�h���k���n���q���t���w��z��}�?�� ���!��y���j���"h���҈��<���������u���܏�rC��[������Es��Oז��:��h�������Va�����#�������塼mF���������aj��1̨�i.��ǐ��`�V������e���}��:೼]B��H������g��Zɺ�+������  �  ��N=�N=�fM=�L=�L=�OK=לJ=V�I=�5I=F�H=��G=�G=�bF=k�E=��D=�AD=N�C=��B=]B=�eA=j�@=z�?=�:?=v�>=>�==	==
L<=
�;=	�:=:= N9=+�8=.�7=7=�?6=�y5=�4=�3=�3=KR2=I�1=1�0=��/=%/=�5.=�[-=\~,=�+=(�*=��)=��(=��'=�'=&=$%=j$=�#=� "=_� =6�=��=~�=sr=�B=�=��=�=;=��=D�=m&=�=H=��=VL=��
=}4	=��==�_=�=�=e��<�6�<.��<�3�<ޣ�<N�<Aj�<n��<(�<"Z�<���<r��<��<TC�<cq�<T��<���<��<��<�!�<*<�<cT�<Kj�<4~�<��<O��<خ�<㻘<�ǔ<wҐ<r܌<��<��<���<z<�r<�'j<H=b<~TZ<�mR<��J<ۧB<��:<��2<[+<|;#<�g<Ɨ<5�<�<�}�; �;8��;Z'�;�κ;x��;�L�;%�;�"|;$^;zQ@;��";�:;���:��:��8:�9�+����&���ܻ��!�����O.�dcH��b�}]{�����U��DU��3������I�Ļ�л!�ڻ��x�������������[M�s���M�7���!��&�"(*��%.��2���5�d�9�=U=�c�@���D�$H� wK��N�b7R���U���X�D\��9_��cb���e�˟h�W�k��n���q���t���w��z�ŗ}��?��ͱ���!���������dh���҈��<���������ku��`܏��B���������`r��N֖��9��h�������w`������#�����塼F��Q������pj��}̨��.��G����󬼴V������?���~��4᳼cC��D���	���h��+ʺ��+�������  �  ��N=eN=�fM=�L=�L=�OK=�J=��I=�5I=��H=�G=0G=cF=��E= �D=�AD=��C=��B=�B=�eA=��@=��?=�:?=��>=;�==	==�K<=�;=��:=�:=�M9=�8=��7=�7=�?6=Sy5=��4=��3=<3=	R2=
�1=��0=��/=	/=�5.=�[-=`~,=�+=D�*=��)=��(=��'=�'=V&=e%=�$= #="=�� =p�=8�=��=�r=�B=�=��=�=�:=a�=�=0&=��=�G=��=L=~�
=&4	=.�=�=1_=��=I=ը�<n6�<׹�<t3�<���<5�<Hj�<���<g�<~Z�<��<���<O�<�C�<�q�<���<E��<6�<�<3"�<�<�<�T�<�j�<g~�<E��<W��<ʮ�<ʻ�<�ǔ<3Ґ<܌<A�<#�<���<��y<�r<~&j<<b<SSZ<�lR<��J<ҦB<��:<\�2<�+<2;#<�g<Ɨ<w�<7<�;��;R��;s)�;�к;ˇ�;�N�;�'�;�'|;)^;�U@;H�";�?;O�:��:P�8:(�9^	+���������޻�a%�)��/S.�(gH�b��a{����X��vW��?������9�Ļ]л��ڻ��9�������������L�����L�2���!��&�'*��$.��2�o�5�[�9�BT=�a�@���D�WH�|vK���N�H7R���U��X��\�h:_��db���e�ˠh�m�k���n���q���t�ùw��z���}�o@��F���$"��V�������h��ӈ��<��{������!u���ۏ�cB�� ���Q���q���Ֆ�9��ٛ������_��d����"�������䡼�E��.�������j���̨��.������U���0W��������j���᳼�C��ܥ�����"i���ʺ�D,������  �  ��N=ON=�fM=�L=�L=PK=��J=��I=�5I=��H=�G=OG=:cF=ǭE=�D=BD=��C=��B=�B=�eA=��@=��?=;?=��>=8�==	==�K<=ۍ;=��:=�:=�M9=ҋ8=��7=�7=�?6=3y5=��4=��3=!3=�Q2=��1=�0=��/=�/=�5.=�[-=d~,=�+=M�*=��)=��(=��'=�'=z&=�%=�$=#=+"=�� =��=J�=��=�r=�B=�=��=�= ;=Q�=	�=!&=��=�G=d�=�K=]�
=4	=	�=�=_=��=;=���<R6�<���<b3�<���<*�<Vj�<���<z�<Z�<4��<��<��<"D�< r�<5��<u��<{�<S�<e"�<�<�<�T�<�j�<}~�<`��<V��<Ȯ�<ǻ�<_ǔ<Ґ<�ی<$�<�<���<n�y< r<&j<;b<�RZ<SlR<9�J<��B<n�:<$�2<�+<$;#<�g<ė<��<l<^�;��; ��;>*�;�Ѻ;�;�O�;�(�;h)|;g+^;�W@;ݳ";�@;��:{��:x�8:@�9
+���� ����໺�&�A���S.��hH��b�_c{�� �� Y��lX����n�����Ļ�л�ڻj���������}��e���L�����L�����!��&��&*�V$.�2���5�Σ9��S=��@���D�KH�VvK��N�47R���U��X��\��:_��db�Ȇe���h�سk�k�n�%�q�M�t�G�w�y�z�V�}��@��^���I"��l���(����h��ӈ��<��j���{��u���ۏ�FB���������q���Ֆ��8�����������_��2���t"�������䡼�E���������j���̨�/������t���KW��0��������⳼2D��������]i���ʺ�],��/����  �  ��N=eN=�fM=�L=�L=�OK=�J=��I=�5I=��H=�G=0G=cF=��E= �D=�AD=��C=��B=�B=�eA=��@=��?=�:?=��>=;�==	==�K<=�;=��:=�:=�M9=�8=��7=�7=�?6=Sy5=��4=��3=<3=	R2=
�1=��0=��/=	/=�5.=�[-=`~,=�+=D�*=��)=��(=��'=�'=V&=e%=�$= #="=�� =p�=8�=��=�r=�B=�=��=�= ;=b�=�=2&=��=�G=��=L=��
=)4	=1�=�=5_=��=M=ި�<w6�<��<}3�<���<>�<Pj�<���<o�<�Z�<��<���<S�<�C�<�q�<���<D��<5�<�</"�<�<�<�T�<�j�<`~�<>��<P��<î�<û�<�ǔ<-Ґ<�ی<<�<�<���<��y<�r<~&j<<b<WSZ<�lR<��J<ܦB<��:<h�2<�+<@;#<�g<ԗ<��<D<4�;��;f��;�)�;�к;҇�;�N�;�'�;�'|;�(^;�U@;�";_?;��:s�:=�8:��9*+���4���m߻�&�x��{S.�qgH�Kb��a{� ��X���W��W������L�Ļnл��ڻ ��E��%�����������L�����L�3���!��&�'*��$.��2�o�5�\�9�CT=�a�@���D�WH�}vK���N�H7R���U��X��\�h:_��db���e�ˠh�m�k���n���q���t�ùw��z���}�o@��F���$"��V�������h��ӈ��<��{������!u���ۏ�cB�� ���Q���q���Ֆ�9��ٛ������_��d����"�������䡼�E��.�������j���̨��.������U���0W��������j���᳼�C��ܥ�����"i���ʺ�D,������  �  ��N=�N=�fM=�L=�L=�OK=לJ=V�I=�5I=F�H=��G=�G=�bF=k�E=��D=�AD=N�C=��B=]B=�eA=j�@=z�?=�:?=v�>=>�==	==
L<=
�;=	�:=:= N9=+�8=.�7=7=�?6=�y5=�4=�3=�3=KR2=I�1=1�0=��/=%/=�5.=�[-=\~,=�+=(�*=��)=��(=��'=�'=&=$%=j$=�#=� "=_� =7�=��=�=tr=�B=�=��= �=;=��=G�=o&=�=H=��=ZL=��
=�4	=��=#=�_=��=�=v��<�6�<@��<�3�<��<_�<Rj�<~��<6�</Z�<���<{��<��<ZC�<fq�<U��<���<��<��<�!�<!<�<XT�<?j�<'~�<��<A��<ˮ�<ջ�<�ǔ<kҐ<g܌<��<��<���<z<�r<�'j<L=b<�TZ<nR<��J<�B<��:<�2<u+<�;#<h<�<Q�<�<�}�;K �;]��;x'�;�κ;���;�L�;%�;�"|;�#^;;Q@;h�";�:;���:��:�8:�݌95+����]���=ݻ��"�}��eP.��cH�wb��]{����V��vU��a������n�Ļ�л>�ڻ3�廎�������������`M�x���M�:���!��&�#(*��%.��2���5�e�9�=U=�c�@���D�%H� wK��N�b7R���U���X�D\��9_��cb���e�˟h�W�k��n���q���t���w��z�ŗ}��?��ͱ���!���������dh���҈��<���������ku��`܏��B���������`r��N֖��9��h�������w`������#�����塼F��Q������pj��}̨��.��G����󬼴V������?���~��4᳼cC��D���	���h��+ʺ��+�������  �  �N=�N=gM=��L=�L=�OK=��J=�I=55I=��H=a�G=�G=]bF=�E=2�D=-AD=ڊC=�B=�B=WeA= �@=F�?=�:?=_�>=2�==*	==-L<=7�;=M�:=d:=�N9=��8=��7=�7=w@6=z5=��4=~�3=�3=�R2=��1=t�0=�/=E/=�5.=�[-=M~,=֝+=��*=��)=h�(=V�'=!'=�&=�%=�$=>#=T "=�� =��=��==�=:r=tB=�=��=(�=E;=��=��=�&=h�=�H=T�=�L=o�
=5	=#�=�=`=w�=	=5��<�7�<˺�<04�<I��<m�<Jj�<R��<��<�Y�<-��<���<�<zB�<hp�<`��<���<��<��<� �<s;�<�S�<�i�<�}�<̏�<��<ͮ�<��<�ǔ<�Ґ<�܌<e�<z�<l��<z<�r<�)j<g?b<�VZ<�oR<��J<��B<��:<<�2<7+<P<#<[h<×<��<X<|�;���;Ί�;�#�;˺;v��;H�;� �;�|;�^;I@;�";�4;���:��:��8:zǌ9_:+����k��ٻ�����'K.�o^H�b��V{�e��`R���Q���������_�Ļh
л^�ڻ��������������&N����O������!�R&� **��'.��2���5�)�9�W=���@�ЄD�2H��wK���N��7R�ÆU�g�X��\� 9_��bb�a�e�"�h���k���n���q���t���w��z��}�?�� ���!��y���j���"h���҈��<���������u���܏�rC��[������Es��Oז��:��h�������Va�����#�������塼mF���������aj��1̨�i.��ǐ��`�V������e���}��:೼]B��H������g��Zɺ�+������  �  i�N=�N="gM= �L=�L=�OK=j�J=��I=�4I=��H=��G=�G=�aF=H�E=��D=�@D=D�C=��B=yB=�dA=��@=��?=}:?=J�>=.�==8	==RL<=u�;=��:=�:= O9=�8=8�7=97=A6=�z5=�4=�3=y3=9S2=
�1=մ0=f�/=u/=�5.=�[-=@~,=��+=��*=:�)=��(=��'=�'=&=%=W$=�
#=��!=k� =L�=<�=ך=�q==B=~=��=:�=r;=��=�=;'=�=0I=��=�M='�
=�5	=��=t=�`=�=�	=A��<�8�<���<�4�<���<��<Nj�<���<��<Y�<_��<���<��<YA�<-o�</��<f��<k�<u�<��<x:�<�R�<	i�<'}�<t��<���<Ǯ�<H��<ZȔ<�Ӑ<�݌<T�<���<���<�z<zr<�,j<Bb<VYZ<prR<ՍJ<��B<��:<��2<H+<�<#<�h<ʗ<��<Z<�y�;���; ��;��;Lƺ;/|�;�B�;��;Y|;�^;�>@;\�";�+;W��:Bו:[�8:|��9�W+������"ջ������D.�WH��b�N{�����M��wM��P��������Ļ,л��ڻ[�廄��P��%�S��W��KO�����P�����!��&��,*�t*.�32��5�t�9�0Y=���@���D��H��xK�f�N��7R�ĆU��X�\��7_�Eab���e�!�h���k���n�#�q��t�"�w�z�z���}�>�����J �����������g���҈��<��ݥ�����Zv���ݏ�VD��\������nt���ؖ��;������� ��tb���Ý��$��|���&桼�F��˧�����Yj���˨� .�������U������C���|��߳�A���������f��MȺ�"*��K����  �  ��N=(N=NgM=�L=�L=�OK=-�J=w�I=`4I=�H=F�G=KG=aF=��E=��D=�?D=��C=��B=�B=`dA=Q�@=��?=E:?="�>=+�==O	==�L<=��;=�:=J:=�O9=��8=��7=�7=�A6=�{5=ڳ4=��3=' 3=�S2=��1=>�0=��/=�/=6.=�[-=,~,=w�+=u�*=��)=��(=R�'='=r&=c%=�$=�	#=�!=�� =��=��=e�=�q=B=\=��=[�=�;=P�=V�=�'=��=�I=��=sN=�
=�6	= =P=�a=�=_
=���<�9�<T��<d5�< ��<��<6j�<���<�<ZX�<u��<���<��<�?�<�m�<���<��<��<�<m�<F9�<�Q�<9h�<�|�<���<���<ޮ�<���<�Ȕ<'Ԑ<�ތ<f�<��<���<�z<�r<�/j<1Eb<T\Z<`uR<��J<�B<��:<[�2<�+<�=#<i<��<��<k <�v�;���;c��;��;���;v�;4<�;��;�|;�^;�2@;J�";�!;���:�ȕ:�o8:���95y+�4���}ϻ������=.�&NH�-�a��C{����<H���G��M��������ĻKл��ڻ9�廷�ﻵ������:��zP�����R�����!�t&�z/*�{-.�G2���5�I�9��[=��@���D�+H��yK�9�N�N8R���U���X�\��6_��_b���e���h�۫k�Ѷn�/�q��t�$�w���z�ѐ}��<��󮁼C�����W���]g��|҈��<��$�������v���ޏ�YE���������u���ٖ�d=�����7���c���ĝ��%��c����桼qG��,���	��3j���˨�t-��z�����T��������G{���ݳ��?������l��8e��Ǻ�)��_����  �   �N=yN=ugM=#�L=pL=ZOK=�J=�I=�3I=eH=��G=�G=K`F=ΪE=�D=?D=ˈC=8�B=?B=�cA=ݫ@=I�?=:?=�>=#�==a	==�L<=�;=n�:=�:=P9=i�8=��7=�7=�B6=I|5=��4=��3=� 3=hT2=!�1=��0=�/=�/=66.=�[-=~,=K�+=#�*=n�)=�(=��'=]'=�&=�%=�$=.	#=Y�!=� =�=�=��=6q=�A=?=��=t�=�;=��=͋=L(=?�=�J=��=IO=��
=�7	=��=>={b=��==��<�:�<H��<6�<e��<��<j�<y��<m�<�W�<���<���<r�<v>�<Jl�<��<]��<i߿<���<�<8�<�P�<Mg�<�{�<���<���<㮜<���<oɔ<�Ԑ<�ߌ<��<�<m��<�z<r<3j<�Hb<�_Z<hxR<Z�J<��B<*�:<-�2<+<�>#<ri<��<b�<k�<�s�;��;�}�;��;V��;io�;{5�;��;��{;��];�%@;�";�;j��:���:Y8:yh�9n�+�����턺Ȼ������5.��DH�V�a��8{��
���B��B��
	��������Ļ5�ϻV�ڻ�~�������^�����Q�X���T�m��H�!��&��2*��0.�f2���5�^�9�f^=���@���D��	H�Z{K���N��8R���U�:�X�#\�:5_��]b�[~e��h��k��n���q���t���w�v�z�	�}�c;��í��.��&��������f��Q҈��<��s���]���w��mߏ�fF��ά��j��aw��tۖ��>���������Ee��EƝ��&��P����硼H������1	��j��a˨��,���������R��8�������y���۳�
>����������c���ź��'��V����  �  ��N=�N=�gM=1�L=bL=2OK=��J=��I=c3I=�~H=��G=�G=�_F= �E=F�D=I>D=�C=��B=�B=DcA=`�@=��?=�9?=�>=�==x	==�L<=a�;=��:=J:=�P9=�8=W�7=v7=eC6=}5=h�4=E�3=�!3=U2=��1=)�0=q�/=2/=^6.=�[-=�},=�+=˸*=�)=��(= �'=�'=&=�%=$=k#=��!=]� =q�=��=x�=�p=rA==�=��=<=��=B�=�(=ܽ=\K=l�=0P=��
=�8	=��=$=`c=��=�=��<�;�<+��<�6�<ץ�<"�<j�<��<��<�V�<|��<a��<�<=�<�j�<|��<���<�ݿ<��<��<�6�<�O�<ff�<+{�<(��<U��<鮜<��<�ɔ<�Ր<z��<��<k�<���<�z<6"r<i6j<�Kb<�bZ<�{R<=�J<�B<>�:< �2<G+<x?#<�i<x�<��<(�<_p�;���;�x�;`�;Q��;�h�;d.�;��;Y�{;^�];�@;�x";�;���:���:>8:�H�9��+�8���넺����z�����-.��;H���a��-{����<��z<��S��H����Ļk�ϻ	�ڻ�{廆��$��+�������_S�,��W���
�!�_!&��5*��3.��2��5�1�9�(a=��@���D��H��|K���N�E9R���U���X�a\��3_�\b�`|e��h�V�k��n���q��t��w�q�z��}�
:������>��K�������f��҈��<���������ux��]����G���������x��ݖ��@��?���F���f���ǝ�(��a����衼�H��ۨ��P	��j��˨�b,����לּ�Q��鳯���Bx��hڳ�{<��t���a ��ab��yĺ��&��k����  �  ��N=�N=�gM=<�L=KL=OK=Q�J=V�I=�2I=J~H=X�G=1G=�^F=A�E=��D=�=D=`�C=��B=B=�bA=�@=��?={9?=�>=�==�	==M<=��;=8�:=�:=HQ9=��8=�7=)	7= D6=�}5=�4=��3=)"3=�U2=&�1=��0=��/=i/=�6.=�[-=�},=ݜ+=��*=��)=�(=��'='=^
&=-%=`$=�#=��!=�� =��=�=��=~p=6A=�
=z�=��=B<=>�=��=_)=x�=L=&�=Q=��
=z9	=|�=�=2d=D�=�=N��<�<�<��<:7�<2��<.�<�i�<���<Y�<V�<���<P��<�	�<�;�<3i�<���<7��<bܿ<���<P�<�5�<�N�<�e�<�z�<���<��<箜<M��<Kʔ<R֐<U�<��<���<>��<�z<5%r<�9j<�Nb<�eZ<b~R<ИJ<s�B</�:<��2<k+<W@#<j<5�<&�<�<�m�;���;5t�;
�;|��;�b�;�'�;���;��{;��];1@;�m";�;��:��:�%8:U(�9��+�V���脺缻���񺨻��%.�i3H��a��#{�����7��M7�����ċ����Ļ��ϻ��ڻ�y���X��V�H�����T����7Y�����!�&$&��8*��6.��2��5��9��c=�;A���D�OH��}K���N��9R���U�9�X��\��2_�~Zb�dze���h��k�#�n�4�q�үt��w���z�H�}��8��d���L������x���:f���ш��<��馋�p��y��3ᏼ�H��2���(��0z���ޖ�B���������h���ȝ�-)��\���5顼?I��B����	���i���ʨ��+��C�����P����������v���س��:���������a��Mú��%�������  �  )�N=6N=�gM=A�L=CL=�NK=�J=��I=�2I=�}H=��G=�G=9^F=��E=��D=�<D=C=I�B=�B=IbA=��@=D�?=G9?=�>=�==�	==9M<=�;=��:=):=�Q9=3�8=��7=�	7=�D6=p~5=��4=��3=�"3= V2=��1=�0=�/=�/=�6.=�[-=�},=��+=B�*=G�)=��(=�'=�'=�	&=�%=�$=#=M�!=$� =M�=��=��=+p=�@=�
=r�=��=f<=��= �=�)=�=�L=��=�Q=g�
=1:	=7�=�=�d=�=!=\��<�=�<���<�7�<v��<S�<�i�<t��<��<\U�<���<X��<��<�:�<h�<���<���<ۿ<u��<3�<�4�<�M�<�d�<z�<]��<�<宜<s��<�ʔ<�֐<�<��<���<d �<<z<�'r<<<j<�Qb<whZ<ʀR<�J<s�B<��:<��2<�+<�@#<Kj<(�<��<&�<�j�;���;+p�;��;{��;P]�;p"�;Y��;�{;��];�@;�c";��;Ɇ�:E��:�8:�99,�����愺(�����=���.��+H���a��{�"����2���2����������3�Ļq�ϻV�ڻ�w�{�����c��������U�H���Z�!����!��&&�%;*�\9.�)"2�~�5�a�9�f=�;A���D��H�K���N�:R���U���X��\��1_� Yb��xe���h�ˡk�߫n���q�i�t�r�w�+�z��}��7��x���s��䊄������e���ш��<��&�������y���ᏼwI��9���F��i{���ߖ�GC���������0i���ɝ�#*��&����顼�I�������	���i���ʨ�q+������-�O����������u���׳��9��Û�������_��Fº��$��Ç���  �  `�N=`N=�gM=M�L=6L=�NK=�J=��I=A2I=s}H=j�G=,G=�]F='�E=`�D=s<D=E�C=��B=B=�aA=J�@=�?=$9?=r>=��==�	==TM<=�;=��:=w:=R9=��8=�7=A
7=@E6=�~5=;�4=��3=&#3=~V2=�1=9�0=7�/=�/=�6.=�[-=�},=��+=�*=�)=U�(=��'=$'=S	&=%=I$=�#=��!=�� =��=6�=Y�=�o=�@=�
=_�=��=�<=��=@�=#*=^�=M=O�=5R=��
=�:	=ˤ=E=ce=n�=�=��<L>�<&��<8�<���<m�<�i�<J��<l�<�T�<��<���<��<�9�<g�<���<���<ڿ<���<[�<�3�<&M�<Md�<�y�<��<Ş�<���<���<˔<Jא<��<E�<y��<O�<*z<�)r<?>j<�Sb<vjZ<��R<ҜJ<˸B<K�:<��2<[+<\A#<�j<��<�<��<�h�;<��;m�;�;���;�X�;�;���;G�{;��];��?;!\";q�;�{�:��::8:w�9�',�	��G儺i���"��0��R.��%H���a��{�s��� /���.��z���e���|�ĻM�ϻO�ڻ�v廎�ﻈ��L�(��L���V�`��\�ʸ���!�|(&�+=*�f;.�5$2���5�L�9��g=��A�ÑD��H��K��N��:R���U���X�4\��0_�Xb�wwe�Q�h��k��n���q�z�t�x�w�>�z�L�}��6��ѩ�����e��������e���ш��<��p�����-z��|⏼J�������b|������HD���������j���ʝ��*������v꡼J��Щ���	���i��aʨ�+��I�����DO����������t���ֳ��8����������_��x���6$��*����  �  ��N=tN=hM=M�L=,L=�NK=њJ=��I=2I=6}H='�G=�G=t]F=ۧE=�D='<D=��C=��B=�B=�aA=�@=��?=9?=g>=��==�	==fM<=*�;=��:=�:=LR9=ܐ8=A�7=�
7=�E6=;5=��4=D�3=d#3=�V2=�1=k�0=[�/=�/=�6.=�[-=�},=�+=�*=��)=�(=}�'=� '=	&=�%=$=T#=��!=n� =��=��= �=�o=�@=�
=[�=��=�<=��=l�=a*=��=YM=��=�R=L�
=;	=!�=�=�e=��=�=���<�>�<r��<T8�<Ϧ�<r�<�i�< ��<3�<�T�<���<��<f�<9�<qf�<��<[��<�ٿ<���<��<T3�<�L�<�c�<^y�<���<���<ﮜ<���<9˔<�א<�<��<���<��<Mz<+r<�?j<�Tb<�kZ<R<��J<ڹB<+�:<��2<�+<�A#<�j<ݖ<��<�<g�;Y��;	k�;���;E��;�V�;{�;*�;�{;��];��?;jW";��;�s�:�}�:��7:��9�8,����-䄺\���{��D���.�n"H�+�a��{�Y����,���,��w���������Ļ��ϻ��ڻ�u���U��i�a�����W���]�ǹ���!��)&�P>*��<.�^%2���5�h�9��h=��A���D��H���K�|�N��:R���U���X�� \�X0_�DWb��ve�R�h��k��n���q�A�t�T�w�4�z�N�}�q6��S���k�����_����e���ш��<������J��qz���⏼�J����������|��Tᖼ�D������t	���j��=˝�`+��+����꡼KJ�������	���i��Gʨ��*������3��N��w���Y��:t��0ֳ�"8��6���U����^�������#��Æ���  �  ��N=�!N=pM=4�L=�L=;YK=�J=��I=�>I=׊H=��G=@"G=�mF=X�E=�E=9PD=��C=��B=�1B=F|A=��@=4@=:Y?=��>=�==�/==su<=4�;=��:=�@:={�9=<�8=�8=qA7=�~6=�5=��4=�/4=ig3=��2=��1=61=D40=�a/=̌.=�-=�,=��+=z+=�5*=�L)=g`(=�o'=3{&=*�%=�$= �#=iz"=`m!=�Z =�A=�"=��= �=�=o`==��=�~=J#=�=�T=7�=f=M�=�X=l�	=�.=h�=��=9==ފ=m��<*�<	��<��<z�<]��<,�<�x�<$��<���<�4�<�g�<a��<���<���<��<-$�<�?�<DY�<Qp�<A��<+��<5��<Q��<�Ť<�Ѡ<�ۜ<u�<��<"�<d��<���< �<��<�z<#r<�j<�'b<]2Z<n>R<ZLJ<\B<n:<V�2<��*<�"<��<��<<�4<ž�;A�;��;k��;"��;!�;���;?w�;3�v;�SX;K:;�t;4��:S��:_�:��:i�'9��V�8�5;���w˺�������6��P���j�k������Ԛ��㦻ն���N���ɻ��Ի?�߻O껡���:����k�5H	�;�U���4�ۢ�c���0$��Q(��Z,��L0��(4�3�7�ʡ;�sA?�X�B�DMF���I��M��pP�9�S� �V�C+Z�V]��x`�Q�c�c�f�K�i�|�l�:�o�\�r�5�u��x��x{��\~�W������Cy���䄼�N��㷇�| ��M����vV������~"��ˇ��2쒼�O��ײ������u���ՙ��4��e����WN��H������d������W��!}��Lۨ��9���������<X��"���@��gx���س��8��;���Z����Y��<�����O|���  �  ��N=�!N=pM=<�L=�L=9YK=%�J=��I=�>I=�H=��G=l"G=�mF=��E=�E=cPD=��C=��B=�1B=b|A=��@=:@=FY?=��>=�==�/==eu<=%�;=��:=�@:=`�9=�8=�8=NA7=�~6=�5=��4=P/4=;g3=~�2=��1=11=840=�a/=ʌ.=��-=�,=��+=�+=�5*=�L)=y`(=p'=^{&=P�%=��$=*�#=�z"=�m!=�Z =�A=�"=�='�=�=f`==��=�~=9#=޿=oT=�=�e=�=�X=<�	=�.=>�=F�===��=>��<�)�<ݣ�<��<z�<]��<�+�<�x�<"��<���< 5�<�g�<���<��<3��<��<�$�<Q@�<�Y�<�p�<q��<T��<K��<u��<�Ť<�Ѡ<�ۜ<n�<��<�<_��<���<���<n�<4z<�r<�j<'b<�1Z<�=R<�KJ<�[B<�m:<�2<��*<ر"<��<��<<"5<��;��;���;y��;���;x�;��;�x�;&�v;�VX;XN:;�v;���:���:�`�:�:ȼ'9Pꏹ��8��;��`x˺�������6��P�#�j�S������֚��䦻G���	P���ɻ�ԻK�߻SO����<����k�:H	�����4�����0$�*Q(�VZ,�KL0�	(4���7��;��@?��B��LF���I��M��pP�P�S��V�D+Z�NV]��x`�d�c���f�Ųi�/�l��o�دr�բu���x�.y{�]]~��������_y���䄼�N�����s ��>����[V������k"�������뒼�O�����g��hu��uՙ��4�������.N��&������d������T��}��[ۨ�:���������jX��f�������x��ٳ�19��{�������Z������K��Y|���  �  }�N=s!N=pM=5�L=�L=QYK=T�J=��I=<?I=>�H=�G=�"G=XnF=�E=`E=�PD=�C=<�B=2B=�|A=��@=q@=tY?=��>=�==�/==Ou<= �;=��:=b@:=�9=��8=`8=�@7=P~6=��5=x�4=�.4=�f3=5�2=��1=�1=40=�a/=��.=�-=�,=�+=�+=�5*=@M)=�`(=\p'=�{&=��%=�$=��#=�z"=�m!=![ =HB= #=6�=R�=-�=l`=	=��=b~=�"=��=T=��=�e=��=[X=��	=&.=Ў=��=�<=[�=~��<:)�<f��<k�<�y�<F��<,�<y�<y��<4��<�5�<�h�<b��<���<���<��<T%�<A�<dZ�<Tq�<��<���<ҩ�<渨<!Ƥ<�Ѡ<�ۜ<T�<��<��<���<7��<7��<��<�z<r<)j<e%b<0Z<8<R<jJJ<NZB<�l:<��2<�*<n�"<��<��<O<�5<���; �;+��;=�;���;��;�;X|�;	�v;_]X;'U:;�|;��:���:j�:@�:��'9_ޏ���8�s<���z˺����c�6���P�̱j����ǐ��ٚ�E离Ӻ��=R����ɻJ�Ի<�߻�P껯��������k��G	�x�G���3�1������.$��O(��X,��J0�_&4��7���;�e??���B��KF���I��M�pP��S�	�V�|+Z��V]��y`�o�c�ܧf��i�b�l�r�o�7�r�t�u�#�x��z{��^~�A���d���y�� 儼O��5���� ��5���zV��E����!������`뒼�N��Ʊ������t���ԙ��3��S���-𝼎M����������d������B��}���ۨ�B:����������X������=��|y���ٳ�:��;���i����Z���������|���  �  9�N=;!N=�oM=&�L=L=�YK=��J=?�I=�?I=��H=��G=e#G=oF=��E=	E=oQD=��C=��B=�2B='}A=8�@=�@=�Y?=ԡ>='�==�/==2u<=Ĺ;=f�:=@:=��9=4�8=�8=I@7=�}6=�5=��4=[.4=Tf3=��2=)�1=�1=�30=�a/=��.=�-=:�,=A�+=�+=*6*=�M)=Na(=�p'=W|&=V�%=��$=3�#=�{"=�n!=�[ =�B=}#=��=��=D�=�`=�=��=&~=�"=!�=�S=�=�d=��=�W=�	=c-=�=!�=�;=��=���<m(�<���<��<�y�<��<9,�<9y�<���<���<y6�<�i�<{��<���<G��<�<�&�<wB�<�[�<�r�<7��<ԙ�<���<n��<�Ƥ<Ҡ<�ۜ<1�<@�<%�<$��<b��<��<��<
z<Jr<�j<�"b<T-Z<�9R<�GJ<\XB<�j:<�2<��*<ΰ"<I�< �<�<�6<`��;##�;E��;��;㋸;y!�;Sș;3��;�v;�iX;`:;W�;���:%��:�w�:��:)0(94̏���8��<��]˺�F���6��P�<�j����t����ݚ�P즻>����V��Ѱɻ+�Ի��߻zR�Թ������k�AG	�����+2�������L,$�M(�V,��G0��#4�U�7�
�;�=?���B��IF��I��M�loP�_�S��V��+Z�NW]��z`���c�k�f���i���l�Һo��r���u���x�F}{� a~�p���\���z���儼�O��t���� ��/����U������*!�����F꒼�M��s���N��Ds��Uә��2������L��ʩ�����d��`�����3}���ۨ��:����������Y�����o���z��۳�E;�����������[��6�������}���  �  ��N=� N=�oM= �L=L=�YK=٦J=��I=$@I=a�H=U�G=$G=�oF=h�E=�E=GRD=��C=��B=Z3B=�}A=��@=2@=�Y?=��>=/�==�/== u<=j�;=��:=t?:=�9=��8=8=�?7=�|6=�5=��4=�-4=�e3=�2=��1=1=d30=Ba/=��.=�-=S�,={�+=Y+=�6*=2N)=�a(=�q'=}&="�%=��$=�#=\|"=9o!=R\ =iC=$=��=��=p�=�`=�=^�=�}=+"=��=�R=T�=�c=�=�V=�	=k,=�=<�=;=��=��<@'�<���<E�<1y�<���<P,�<�y�<���<���<�7�<�j�<ۘ�<u��<���<�	�<i(�< D�<9]�<�s�<���<��<���<3��<Ǥ<@Ҡ<�ۜ<�<��<m�<��<)��<���<
 �<�z<�r<�j<	b<�)Z<k6R<�DJ<�UB<~h:<�}2<n�*<�"<�<�<�<�7<��;'�;���;��; ��;n(�;�ϙ;���;N�v;xX;lm:;��;8��:'��:)��:9:|(9�m�8�?����˺}�j�Ƭ6���P���j�1��^����㚻]��Ĳ��[����ɻs�Ի!�߻U�ʻ��q����k��F	������0�2�����p)$�	J(��R,��D0�< 4��7���;�J:?���B��GF��I��M�inP��S��V�,Z�]X]�|`���c���f���i���l�ܽo�4�r�?�u��x�r�{�d~�١������{���愼MP��⸇�� ��&����)U��κ��$ ��ل���蒼[L��㮕�����q���љ��0�������흼<K���������bc���������<}���ۨ�F;��Ӛ������
[��j������E|���ܳ��<��2���:���`]����������~���  �  [�N=� N=�oM=�L=2L=�YK=;�J=*�I=�@I=�H=*�G=%G=�pF=e�E=�E=@SD=s�C=y�B=#4B=y~A=T�@=�@=IZ?=.�>=@�==t/==�t<=�;=v�:=�>:=J�9=��8= 8=�>7=�{6=�5=�4=�,4=�d3=D�2=��1=�1= 30=�`/=Z�.=�-=p�,=��+=�+= 7*=�N)=�b(={r'= ~&=�%=��$= �#=I}"=p!=2] =D=�$=h�=.�=��=�`=�=�=b}=�!=ܽ=R=l�=�b=��=�U=��	=?+=�=�=:=�=t��<�%�<���<m�<�x�<���<k,�<z�<F��<���<�8�<Dl�<���<J��<���<��<n*�<F�<1_�<�u�<��<l��<���<��<�Ǥ<�Ҡ<�ۜ<��<(�<��<��<���<$��<7��<�z<�	r<�j<�b<�%Z<�2R<~AJ<wRB<�e:<�{2<��*<Ѯ"<�<N�<t<D9<���;�,�;���;��;B��;�0�;vؙ;���;��v;7�X;�~:;z�;T��:�:���:H<:��(9���Ի8��B��c�˺��r�~�6���P���j�
!��|���+뚻 ���
̲�4b��9�ɻm�Ի'�߻�W껢�������|k�F	�U���.�^������%$�2F(��N,�t@0�/4��7�-�;��6?���B��DF��I�mM�mP�^�S��V��,Z�qY]�|}`�c�\�f���i���l���o��r�W�u��x�1�{��g~�t�����}���焼�P��l���!�����xmT��������s���^璼zJ���������o���ϙ�/�������라�I��g�������b��t������Y}��dܨ��;������ ���n\���������3~���޳��>�����(���,_��!���^������  �  ��N=@ N=IoM= �L=IL=#ZK=��J=��I=sAI=׍H=�G=&G=�qF=v�E=�E=TTD=s�C=f�B=�4B=8A=��@=@=�Z?=[�>=R�==[/==t<=��;=��:=5>:=v9=ӿ8=*�7=�=7=�z6=��5=�4=�+4=�c3=b�2=3�1=�1=20=�`/=(�.=�-=��,=�+='+=�7*=�O)=qc(=[s'=�~&=�%=��$= �#=O~"=q!=^ =�D=L%=��=��=�=�`=�=��=�|=!="�==Q=c�=�a=��=JT=��	=*=��=��=9=
�=О�<f$�<���<��<x�<���<~,�<�z�<��<� �<5:�<�m�<n��<:��<��<��<�,�<>H�<*a�<�w�<ȋ�<ꝰ<ڭ�<��<EȤ<�Ҡ<�ۜ<C�<��<��<��<=��<S��<S��<��y<�r<$j<�b<p!Z<|.R<�=J<OB<	c:<2y2<5�*<��"<�<~�<.<�:<���;N2�;���;Q�;d��;�9�;��;��;7�v;~�X;
�:;t�;v�:%,�:���:�]:�*)9�}���8�F��̔˺k �c���6�"Q�b�j�r(�����󚻶 ��pӲ��h����ɻ��Իe�߻u[껾�������Ek�}E	�"�����+�w�����"$�NB(��J,�6<0��4���7�D�;��2?���B��AF���I��M��kP�ӶS���V�o-Z��Z]�g`��c��f��i�~�l���o���r���u��x�N�{��k~�:������f~���脼�Q��򹇼J!��퇊�'�S�������������咼�H��
������{m���͙��,��׋��3ꝼFH���������a��������f}���ܨ��<��˜��/����]������x��6����೼A��*���-��a������� ������  �  P�N=�N=oM=�L=XL=`ZK= �J=7�I=BI=��H=��G=�&G=�rF=��E= 
E=[UD=t�C=N�B=�5B=�A=��@=�@=�Z?=��>=V�==@/==@t<=F�;=]�:=�=:=�~9=�8=8�7=|<7=�y6=�5=��4=�*4=�b3=��2=x�1=U1=20=X`/= �.=ִ-=��,=O�+=�+=B8*=0P)=Hd(=9t'=�&=�%=��$=�#=M"=�q!=�^ =�E=�%=q�=��=�=�`=�=��=�|=s =`�=]P=k�=�`=��=	S=_�	=�(=}�=��=�7=�=��<�"�<S��<��<�w�<U��<�,�<�z�<���<��<~;�<|o�<)��<1��<��<�<�.�<VJ�< c�<�y�<���<@��<��<켨<�Ȥ<Ӡ<�ۜ<��<��<��<x�<��<���<d��<k�y<� r<�j<�b<Z<e*R<�9J<�KB<`:<�v2<`�*<��"<��<��<	<E<<@��;R7�;���;�!�;g��;pB�;�;���;��v;֭X;��:;)�;1�:@D�:�ǈ:c}:2�)9�g��W�8�1I���˺�&�w'�f�6�{Q���j�0��豎���������ڲ��o����ɻ��Ի��߻�^���������Uk��D	�����8)�Ȕ���w$�[>(�cF,��70��4���7�L�;�\/?�)�B�:?F�G�I��M��jP�(�S�	�V��-Z��[]�D�`���c��f�:�i��l���o�H�r���u�P�x���{��o~����S������鄼�R��v����!�������틼"S�������������㒼�F��
���{
��Xk��q˙��*������k蝼�F��̤����� a������T���}��0ݨ�F=��Ɲ�����n_��o���U!��:����⳼/C��O���7���b���º�o"��o����  �  ��N=|N=�nM=ֽL=nL=�ZK=M�J=��I=�BI=V�H=��G=�'G=�sF=u�E=E=JVD=l�C=-�B=�6B=��A=%�@=@=B[?=Ȣ>=a�==%/==�s<=�;=��:=�<:=�}9=�8=F�7=�;7=�x6=��5=��4=�)4=b3=И2=��1=� 1=�10=�_/=֋.=ʴ-=��,=��+=�+=�8*=�P)= e(=u'=π&=�%=��$=�#=0�"=�r!=�_ =UF=~&=��=8�=C�=�`=j=H�=|=�=��=�O=��=�_=~�=�Q=3�	=�'=\�=��=�6=/�=b��<�!�<H��<��<w�<!��<�,�<P{�<���<��<�<�<�p�<ϟ�<��<���<�<�0�<ML�<e�</{�<
��<���<0��<���<wɤ<jӠ<�ۜ<��<�<��<C��<N�<���<o��<{�y<��q<�j<�b<�Z<L&R<46J<�HB<?]:<�t2<��*<~�"<
�<��<�<r=<D��;`<�;���;�(�;=��;�J�;s�;���;��v;i�X;!�:;��;�K�:�[�:pڈ:T�:��)9�O��;�8��M��-�˺�,�R0��6��Q���j�	7��A���������᲻�v��i�ɻ�Ի�߻�a�~�������\k�D	�� ����'�����)$�~:(��B,��30��4���7�p�;�,?�&�B��<F� �I�=M��iP�~�S� �V��.Z�(]]�ɂ`���c���f�0�i���l�H�o�$�r���u�R�x�Y�{�Gs~�˨�����&����ꄼqS������!��懊�\틼�R��8���q��4��kⒼ$E��������Oi���ə�	)������杼7E���������b`�� ������}���ݨ�>�����������`��¯�9#������䳼'E��G������d��Gĺ��#�������  �  j�N=.N=�nM=ǽL=uL=�ZK=��J=�I=2CI=�H=c�G=�(G=�tF=G�E=�E=WD=1�C=��B=M7B=>�A=��@=p@=�[?=�>=e�==/==�s<=��;=j�:=O<:=R}9=`�8=��7=�:7=�w6=�5=#�4=�(4=La3=�2=(�1=D 1=410=�_/=��.=ƴ-=��,=��+=D+=69*=`Q)=�e(=�u'=��&=Ɉ%=M�$=̈#=��"=�s!=T` =�F='=P =��=q�=�`=S=�=�{=m=�=�N=��=�^=��=�P=2�	=�&=g�=��=
6=b�=���<h �<K��<1�<�v�<���<�,�<�{�<��<��<�=�<+r�<6��<���<���<��<^2�<�M�<�f�<�|�<Y��<ġ�<��<f��<�ɤ<�Ӡ<�ۜ<S�<��<��<6�<�<��<���<&�y<H�q<� j<
b<�Z<*#R<*3J<�EB<�Z:<�r2<0�*<��"<��<��<|<�><���;�@�;ȱ�;z.�;���;�Q�;���;���;�w;��X;��:;e�;*c�:�o�:[�:��:�#*9?���8��P����˺�2��7�0�6��%Q�5k��<������u��)���粻�{����ɻ��Ի��߻�d�N�������Hk��C	������&%�Ə����?$�u7(�\?,��00�J4���7�c�;�)?���B�F:F�?�I��M��hP�<�S��V�/Z�*^]�e�`���c��f���i���l�W�o�o�r�#�u���x���{�Iv~�0�����D����넼.T�������!��ᇊ�,틼�Q��z���t��~��ᒼ�C����������g���Ǚ�y'������t坼�C��w���� ���_���������}���ݨ��>������� ��b��jï��$������z泼�F���������:f���ź�%�������  �  �N=�N=}nM=��L=�L=�ZK=ڨJ=^�I=�CI=b�H=��G=+)G=0uF=��E=yE=�WD=ϢC=��B=�7B=��A=��@=�@=�[?=��>=o�==�.==�s<=P�;=�:=�;:=�|9=Ѽ8=��7=	:7=Cw6=n�5=u�4=F(4=�`3=��2=��1=��0=�00=�_/=��.=Ŵ-=��,=��+=�+=9*=�Q)=f(=Jv'=�&=s�%=�$=h�#=��"=-t!=�` =dG=Z'=� =��=��=�`=E=��=~{==��=NN=�=;^=��='P=n�	=�%=��=�=_5=��=��<~�<���<��<9v�<���<�,�<�{�<���<@�<�>�<.s�<^��<���<���<�<�3�<AO�<�g�<�}�<O��<���<���<쾨<.ʤ<�Ӡ<�ۜ<��<7�<3�<u�<�<_�<���<Y�y<w�q<�i<Jb<�Z<� R<�0J<�CB<5Y:<?q2<=�*<��"<H�<��<�<�?<���;�C�;��;S3�;���;7W�;{ �;���;�w;��X;��:;��;Ls�:�}�:���:��:!R*9=.���8��S���˺7��<��6��-Q�Pk��A��pĎ�d��A��{첻?�����ɻ��Ի}�߻�f�T�������5k�dC	������#�0�����$�5(��<,�.0��	4���7� �;��&?���B��8F���I��M�	hP��S��V��/Z��^]���`��c���f��i���l���o�*�r���u�^�x�[�{��x~�N���'������센�T��׻��8"��ч���싼�Q���������7}������B��]������ef���ƙ�*&��t���L䝼C������o ��<_��i�������}��Oި��>��*���|�� c���į��%��
����糼8H��L�����ng���ƺ�&��z����  �  ��N=�N=hnM=��L=�L=�ZK=��J=��I=�CI=��H=?�G=�)G=�uF=P�E=�E=%XD=+�C=��B=!8B=�A=F�@=�@=�[?=�>=u�==�.==zs<=�;=��:=�;:=}|9=z�8=��7=�97=�v6=�5=�4=�'4=^`3=C�2=i�1=��0=�00=d_/=p�.=��-=��,=�+=�+=�9*=
R)=af(=�v'=t�&=ɉ%=P�$=̉#=�"=�t!=+a =�G=�'=� =��=��=�`=:=��=J{=�=X�=�M=��=�]=j�=�O=��	=]%=.�=��=�4=`�=E��<��<��<Y�<	v�<���<�,�<|�<���<��<?�<�s�<���<~��<���<��<{4�<�O�<�h�<u~�<鑴<.��<7��<:��<\ʤ<�Ӡ<�ۜ<��<��<��<��<i��<��<��<��y<��q<J�i<�b<Z<�R<[/J<BBB<�W:<Cp2<p�*<G�"<&�<�<1<0@<���;WF�;���;�5�;���;lZ�;��;9��;w;S�X;��:;�;c~�:���:���:s�:�p*9@%����8�4V���˺F:��@���6��2Q��k��D��uǎ�z����3ﲻ���� �ɻ3�Իf�߻}h껒���?���8k�,C	����`���"����Q���$��3(�2;,�b,0�4��7���;��%?�e�B��7F��I�M��gP���S��V��/Z�^_]�`�`�
�c���f�N�i�V�l�^�o���r�j�u���x�ɗ{�?z~� ����������턼U�����R"��Ǉ���싼nQ������>���|��zߒ��A����������e���ř�r%��Ǆ���㝼�B��$��������^��A�������}��wި�U?������
���c��&ů��&�������購	I��������)h��jǺ��&������  �  ��N=�N=knM=��L=�L=�ZK=
�J=��I=�CI=ŐH=c�G=�)G=�uF=q�E=E=DXD=Z�C=��B=C8B=	�A=K�@=�@=�[?=�>=l�==�.==vs<=�;=��:=�;:=i|9=W�8=a�7=�97=�v6=ܲ5=��4=�'4=3`3=+�2=N�1=��0=�00=U_/=v�.=��-=��,=�+=�+=�9*=R)=}f(=�v'=��&=�%=u�$=�#=�"=�t!=Va =�G=�'=� =��=��=�`=0=��=9{=�=L�=�M=��=�]=9�=�O=Ž	=.%=�=u�=�4=I�=��<��<���<C�<	v�<���<�,�<<|�<���<��<E?�<�s�<T��<���<���<1�<�4�<IP�<�h�<�~�<��<A��<J��<X��<uʤ<�Ӡ<�ۜ<��<��<��<��<0��<s�<��<!�y<&�q<��i<�b<kZ<AR<�.J<�AB<�W:<(p2<6�*<U�"<�<��<]<n@<��;�F�;ٸ�;7�;(¸;�[�;��;���;Cw;�X;��:;Z�;���:��:C �:��:�z*9�(��W�8��V��j�˺�:��A��6��4Q�Jk��E���Ȏ����Q����D�����ɻ�Ի��߻�h��������Rk�7C	�h��)���"��������$��2(��:,��+0�{4��7�;��$?��B�=7F�٩I��M�ZgP���S�.�V��/Z��_]���`�-�c�i�f���i���l��o�B�r��u���x�f�{��z~�K������Ӄ��턼0U��'���M"��؇���싼NQ��w���6��x|��9ߒ��A��D������Be���ř�(%��j���k㝼MB����������^��&�������}��jި�o?������$���c��dů��&������購_I��g���	���h���Ǻ��&��,����  �  ��N=�N=hnM=��L=�L=�ZK=��J=��I=�CI=��H=?�G=)G=�uF=P�E=�E=%XD=+�C=��B=!8B=�A=F�@=�@=�[?=�>=u�==�.==zs<=�;=��:=�;:=}|9=z�8=��7=�97=�v6=�5=�4=�'4=^`3=C�2=i�1=��0=�00=d_/=p�.=��-=��,=�+=�+=�9*=
R)=af(=�v'=t�&=ɉ%=P�$=̉#=�"=�t!=+a =�G=�'=� =��=��=�`=;=��=K{=�=Z�=�M=��=�]=n�=�O=��	=b%=3�=��=�4=e�=Q��<��<%��<e�<v�<���<�,�<)|�<���<��<'?�<�s�<���<���<���<��<z4�<�O�<~h�<p~�<㑴<'��<.��<1��<Rʤ<�Ӡ<�ۜ<��<��<��<��<b��<��<��<��y<��q<J�i<�b<Z<R<f/J<OBB<X:<Tp2<��*<Z�"<9�<'�<D<B@<���;uF�;��;�5�;���;vZ�;��;6��;w;4�X;Y�:;��;�}�:��:���:�:�j*9k(��S�8�W����˺�:�QA�Y�6�3Q��k��D���ǎ����/��Rﲻ����ɻI�Իy�߻�h껠���L���=k�0C	����c���"����S���$��3(�3;,�c,0�4���7���;��%?�e�B��7F��I�M��gP���S��V��/Z�^_]�`�`�
�c���f�O�i�V�l�^�o���r�j�u���x�ɗ{�?z~� ����������턼U�����R"��Ǉ���싼nQ������>���|��zߒ��A����������e���ř�r%��Ǆ���㝼�B��$��������^��A�������}��wި�U?������
���c��&ů��&�������購	I��������)h��jǺ��&������  �  �N=�N=}nM=��L=�L=�ZK=ڨJ=^�I=�CI=b�H=��G=+)G=0uF=��E=yE=�WD=ϢC=��B=�7B=��A=��@=�@=�[?=��>=o�==�.==�s<=P�;=�:=�;:=�|9=Ѽ8=��7=	:7=Cw6=n�5=u�4=F(4=�`3=��2=��1=��0=�00=�_/=��.=Ŵ-=��,=��+=�+=9*=�Q)=f(=Jv'=�&=s�%=�$=h�#=��"=-t!=�` =eG=['=� =��=��=�`=G=��=�{==��=RN=�=A^=��=-P=u�	=�%=��=�=i5=Ƀ=��<��<���<��<Pv�<���<�,�<|�<���<Q�<�>�<:s�<h��<���<���<�<�3�<=O�<�g�<�}�<C��<���<���<ھ�<ʤ<�Ӡ<�ۜ<��<&�<#�<g�<�<T�<���<M�y<q�q<�i<Ob<�Z<� R<�0J<�CB<SY:<`q2<a�*<ҩ"<n�< �<<�?<���;!D�;���;|3�;ؽ�;JW�;� �;���;`w;��X;O�:;*�;Pr�:�|�:z�:7�:sF*9Z4��@�8��U����˺�7�`=�?�6�h.Q��k�NB���Ď��������첻t�����ɻ��Ի��߻g�p�������?k�mC	�&�����#�4������$�5(��<,�.0��	4���7��;��&?���B��8F���I��M�	hP��S��V��/Z��^]���`��c���f��i���l���o�*�r���u�^�x�[�{��x~�N���'������센�T��׻��8"��ч���싼�Q���������7}������B��]������ef���ƙ�*&��t���L䝼C������o ��<_��i�������}��Oި��>��*���|�� c���į��%��
����糼8H��L�����ng���ƺ�&��z����  �  j�N=.N=�nM=ǽL=uL=�ZK=��J=�I=2CI=�H=c�G=�(G=�tF=G�E=�E=WD=1�C=��B=M7B=>�A=��@=p@=�[?=�>=e�==/==�s<=��;=j�:=O<:=R}9=`�8=��7=�:7=�w6=�5=#�4=�(4=La3=�2=(�1=D 1=410=�_/=��.=ƴ-=��,=��+=D+=69*=`Q)=�e(=�u'=��&=ʈ%=M�$=̈#=��"=�s!=U` =�F='=Q =��=r�=�`=V=�=�{=r=�=�N=��=�^=��=�P==�	=�&=s�=��=6=q�=��<� �<l��<R�<�v�<��<�,�<�{�<6��<��<�=�<=r�<D��<���<���<��<\2�<�M�<�f�<�|�<H��<���<��<N��<�ɤ<oӠ<�ۜ<9�<y�<��<!�<��<r�<���<�y<?�q<� j<%
b<�Z<A#R<H3J<�EB<[:<�r2<b�*<ɪ"<��<�<�<�><���;*A�;��;�.�;���;�Q�;���;�;Zw;6�X;"�:;��;�a�:?n�:��:��:*9�G����8�)S��8�˺�3��8�@�6��&Q�,k�b=��򿎻�������粻A|����ɻ��Ի �߻�d�v�������Vk��C	����#��.%�̏����C$�y7(�^?,��00�K4���7�d�;�)?���B�G:F�?�I��M��hP�<�S��V�/Z�+^]�e�`���c��f���i���l�W�o�o�r�#�u���x���{�Iv~�0�����D����넼.T�������!��ᇊ�,틼�Q��z���t��~��ᒼ�C����������g���Ǚ�y'������t坼�C��w���� ���_���������}���ݨ��>������� ��b��jï��$������z泼�F���������:f���ź�%�������  �  ��N=|N=�nM=ֽL=nL=�ZK=M�J=��I=�BI=V�H=��G=�'G=�sF=u�E=E=JVD=l�C=-�B=�6B=��A=%�@=@=B[?=Ȣ>=a�==%/==�s<=�;=��:=�<:=�}9=�8=F�7=�;7=�x6=��5=��4=�)4=b3=И2=��1=� 1=�10=�_/=֋.=ʴ-=��,=��+=�+=�8*=�P)= e(=u'=π&=�%=��$=�#=0�"=�r!=�_ =VF=&=��=:�=E�=�`=m=L�=|=�=��=�O=��=�_=��=�Q=@�	=�'=l�=��=�6=A�=���<�!�<p��<	�<;w�<H��<�,�<s{�<���<��<�<�<q�<���<#��<���<�<�0�<EL�<�d�<{�<���<~��<��<���<Xɤ<JӠ<�ۜ<�<��<��<*��<8�<���<a��<g�y<��q<�j<�b<
Z<i&R<Y6J<�HB<s]:<u2<؎*<��"<L�<�<+<�=<���;�<�;��;�(�;r��;�J�;��;���;g�v;�X;��:;�;4J�:�Y�:A؈:��:��)9�Z����8�}P���˺�-��1�i�6�Q���j��7��ƹ��}��g�� ⲻ�v����ɻc�ԻM�߻�a껮�������nk� D	�� ����'�!����/$��:(��B,��30��4���7�r�;�,?�'�B��<F�!�I�>M��iP�~�S� �V��.Z�(]]�ɂ`���c���f�0�i���l�H�o�$�r���u�R�x�Y�{�Gs~�˨�����&����ꄼqS������!��懊�\틼�R��8���q��4��kⒼ$E��������Oi���ə�	)������杼7E���������b`�� ������}���ݨ�>�����������`��¯�9#������䳼'E��G������d��Gĺ��#�������  �  P�N=�N=oM=�L=XL=`ZK= �J=7�I=BI=��H=��G=�&G=�rF=��E= 
E=[UD=t�C=N�B=�5B=�A=��@=�@=�Z?=��>=V�==@/==@t<=F�;=]�:=�=:=�~9=�8=8�7=|<7=�y6=�5=��4=�*4=�b3=��2=x�1=U1=20=X`/= �.=ִ-=��,=O�+=�+=B8*=0P)=Hd(=9t'=�&=�%=��$=�#=M"=�q!=�^ =�E=�%=r�=��=�=�`=�=��=�|=y =f�=eP=t�=�`=��=S=m�	=�(=��=��=8='�==��<#�<���<��<�w�<���<�,�<{�<��<��<�;�<�o�<<��<?��<��<�<�.�<MJ�<c�<qy�<j��<%��<���<˼�<�Ȥ<�Ҡ<�ۜ<��<��<o�<[�<��<��<T��<V�y<� r<�j<�b<!Z<�*R<�9J<�KB<@`:<w2<��*<ެ"<��<��<P<�<<���;�7�;��;6"�;���;�B�;�;{��;|�v;d�X;V�:;_�;+/�:B�:ň:x:�r)9�s��l�8�HL���˺w(��(���6��Q�0�j��0��|���2���9	��.۲�p��+�ɻ8�ԻF�߻_�$�������ik��D	���#��B)�Д�$��}$�`>(�gF,��70��4���7�N�;�]/?�*�B�;?F�G�I��M��jP�)�S�
�V��-Z��[]�D�`���c��f�:�i��l���o�H�r���u�P�x���{��o~����S������鄼�R��v����!�������틼"S�������������㒼�F��
���{
��Xk��q˙��*������k蝼�F��̤����� a������T���}��0ݨ�F=��Ɲ�����n_��o���U!��:����⳼/C��O���7���b���º�o"��o����  �  ��N=@ N=IoM= �L=IL=#ZK=��J=��I=sAI=׍H=�G=&G=�qF=v�E=�E=TTD=s�C=f�B=�4B=8A=��@=@=�Z?=[�>=R�==[/==t<=��;=��:=5>:=v9=ӿ8=*�7=�=7=�z6=��5=�4=�+4=�c3=b�2=3�1=�1=20=�`/=(�.=�-=��,=�+='+=�7*=�O)=qc(=\s'=�~&=�%=��$= �#=P~"=q!=^ =�D=M%=��=��=�=�`=�=��=�|=!=)�=EQ=l�=�a=��=WT=��	=*=͊=�=9=�=���<�$�<���<��<Dx�<���<�,�<�z�<-��<� �<R:�<�m�<���<H��<��<��<�,�<5H�<a�<�w�<���<Ν�<���<仨<!Ȥ<�Ҡ<�ۜ<�<b�<c�<��<$��<>��<B��<��y<ur<$j<�b<�!Z<�.R<�=J<:OB<Ec:<ty2<|�*<�"<c�<��<x<;<\��;�2�;X��;��;���;�9�;��;���;��v;	�X;e�:;��;�:�)�:��:0X:�)9���_�8�8I�� �˺"���O�6��Q���j�)��������7���Ӳ�>i��)�ɻ��Ի��߻�[����� ���Yk��E	�1����+�������"$�SB(��J,�9<0��4���7�F�;��2?���B��AF���I��M��kP�ӶS���V�o-Z��Z]�g`��c��f��i�~�l���o���r���u��x�N�{��k~�:������f~���脼�Q��򹇼J!��퇊�'�S�������������咼�H��
������{m���͙��,��׋��3ꝼFH���������a��������f}���ܨ��<��˜��/����]������x��6����೼A��*���-��a������� ������  �  [�N=� N=�oM=�L=2L=�YK=;�J=*�I=�@I=�H=*�G=%G=�pF=e�E=�E=@SD=s�C=y�B=#4B=y~A=T�@=�@=IZ?=.�>=@�==t/==�t<=�;=v�:=�>:=J�9=��8= 8=�>7=�{6=�5=�4=�,4=�d3=D�2=��1=�1= 30=�`/=Z�.=�-=p�,=��+=�+= 7*=�N)=�b(={r'= ~&=�%=��$= �#=I}"=p!=2] =D=�$=j�=0�=��=�`=�=�=g}=�!=�=R=u�=�b=��=�U=��	=O+=�=/�=+:='�=���<&�<��<��<�x�<���<�,�<?z�<j��<���<�8�<\l�<���<W��<���<��<k*�<F�<#_�<�u�<��<Q��<���<���<�Ǥ<hҠ<�ۜ<}�<�<l�<��<���<��<'��<�z<�	r<�j< b<�%Z<�2R<�AJ<�RB<�e:<�{2<:�*<�"<��<��<�<�9<7��;&-�;��;7�;|��;�0�;�ؙ;���;��v;ňX;*~:;��;n��:��:D��:�6:�(9����8��E��{�˺+����6��P�&�j��!������뚻����{̲��b����ɻ��Իn�߻X�ؽ�������k�-F	�c����.�f������%$�7F(��N,�w@0�14� �7�/�;��6?���B��DF��I�nM�mP�_�S��V��,Z�qY]�}}`�c�\�f���i���l���o��r�W�u��x�1�{��g~�t�����}���焼�P��l���!�����xmT��������s���^璼zJ���������o���ϙ�/�������라�I��g�������b��t������Y}��dܨ��;������ ���n\���������3~���޳��>�����(���,_��!���^������  �  ��N=� N=�oM= �L=L=�YK=٦J=��I=$@I=a�H=U�G=$G=�oF=h�E=�E=GRD=��C=��B=Z3B=�}A=��@=2@=�Y?=��>=/�==�/== u<=j�;=��:=t?:=�9=��8=8=�?7=�|6=�5=��4=�-4=�e3=�2=��1=1=d30=Ba/=��.=�-=S�,={�+=Y+=�6*=2N)=�a(=�q'=}&="�%=��$=�#=\|"=9o!=R\ =jC=$=��=��=s�=�`=�=b�=�}=0"=��=�R=\�=�c=�=�V=�	=y,= �=M�=%;=�=;��<g'�<ܡ�<m�<Yy�<��<v,�<�y�<ƿ�<���<�7�<�j�<��<���<���<�	�<f(�<D�<,]�<�s�<���<隰<���<��<�Ƥ< Ҡ<�ۜ<��<��<Q�<��<��<���<���<�z<�r<�j<b<*Z<�6R<EJ<�UB<�h:< ~2<��*<C�"<F�<]�<�<8<���;�'�;��;�;U��;�(�;�ϙ;퉊;�v;�wX;�l:;ϓ;���:2��:���:y:�g(9������8��A��~�˺�����6���P���j����㛎�#䚻��EŲ�S\���ɻ��Ի`�߻UU����������k��F	������&0�:�����v)$�J(��R,��D0�? 4��7���;�K:?���B��GF��I��M�jnP��S��V�,Z�]X]�|`���c���f���i���l�ܽo�4�r�?�u��x�r�{�d~�١������{���愼MP��⸇�� ��&����)U��κ��$ ��ل���蒼[L��㮕�����q���љ��0�������흼<K���������bc���������<}���ۨ�F;��Ӛ������
[��j������E|���ܳ��<��2���:���`]����������~���  �  9�N=;!N=�oM=&�L=L=�YK=��J=?�I=�?I=��H=��G=e#G=oF=��E=	E=oQD=��C=��B=�2B='}A=8�@=�@=�Y?=ԡ>='�==�/==2u<=Ĺ;=f�:=@:=��9=4�8=�8=I@7=�}6=�5=��4=[.4=Tf3=��2=)�1=�1=�30=�a/=��.=�-=:�,=A�+=�+=*6*=�M)=Na(=�p'=W|&=V�%=��$=3�#=�{"=�n!=�[ =�B=~#=��=��=E�=�`=�=��=)~=�"=&�=�S=!�=�d=��=�W=�	=o-=�=/�=�;=ω=���<�(�<Ӣ�<�<�y�<<��<X,�<Vy�<��<���<�6�<�i�<���<���<M��<�<�&�<qB�<�[�<ur�<&��<���<���<V��<{Ƥ<�Ѡ<�ۜ<�<(�<�<��<O��<
��<�<
z<Ar<�j<�"b<d-Z<�9R<HJ<�XB<k:<�2<'�*<�"<�<6�<1<�6<���;v#�;���;%�;��;�!�;]ș;,��;�v;6iX;�_:;;z��:���:v�:��:�(9�ԏ���8�-?����˺��_���6��P�3�j�	��ᕎ��ݚ��즻�����V���ɻf�Իή߻�R�����-����k�MG	���'��22�������P,$�!M(�V,��G0��#4�V�7��;� =?���B��IF��I��M�moP�`�S��V��+Z�NW]��z`���c�k�f���i���l�Һo��r���u���x�F}{� a~�p���\���z���儼�O��t���� ��/����U������*!�����F꒼�M��s���N��Ds��Uә��2������L��ʩ�����d��`�����3}���ۨ��:����������Y�����o���z��۳�E;�����������[��6�������}���  �  }�N=s!N=pM=5�L=�L=QYK=T�J=��I=<?I=>�H=�G=�"G=XnF=�E=`E=�PD=�C=<�B=2B=�|A=��@=q@=tY?=��>=�==�/==Ou<= �;=��:=b@:=�9=��8=`8=�@7=P~6=��5=x�4=�.4=�f3=5�2=��1=�1=40=�a/=��.=�-=�,=�+=�+=�5*=@M)=�`(=\p'=�{&=��%=�$=��#=�z"=�m!=![ =HB=!#=7�=S�=.�=n`==��=e~=#=��=T=��=�e=��=bX=��	=/.=َ=��=�<=f�=���<Q)�<}��<��<�y�<]��<,�<#y�<���<E��<�5�<�h�<l��<���<���<��<R%�<A�<]Z�<Jq�<��<<©�<ո�<Ƥ<�Ѡ<�ۜ<B�<��<��<���<*��<,��<��<�z<r<)j<j%b<0Z<H<R<JJ<hZB<�l:<�2</�*<��"<��<��<t<�5<���;M �;]��;f�;Ά�;��;�;S|�;�v;$]X;�T:;~|;���:���:�h�:��:�'9|䏹�8�>���|˺j�m�#�6���P�{�j�#�����Oٚ��离���rR��'�ɻt�Իa�߻�P�ʸ�������k��G	��M���3�6������.$��O(��X,��J0�a&4��7���;�f??���B��KF���I��M�pP��S�	�V�|+Z��V]��y`�o�c�ܧf��i�b�l�r�o�7�r�t�u�#�x��z{��^~�A���d���y�� 儼O��5���� ��5���zV��E����!������`뒼�N��Ʊ������t���ԙ��3��S���-𝼎M����������d������B��}���ۨ�B:����������X������=��|y���ٳ�:��;���i����Z���������|���  �  ��N=�!N=pM=<�L=�L=9YK=%�J=��I=�>I=�H=��G=l"G=�mF=��E=�E=cPD=��C=��B=�1B=b|A=��@=:@=FY?=��>=�==�/==eu<=%�;=��:=�@:=`�9=�8=�8=NA7=�~6=�5=��4=P/4=;g3=~�2=��1=11=840=�a/=ʌ.=��-=�,=��+=�+=�5*=�L)=y`(=p'=^{&=P�%=��$=+�#=�z"=�m!=�Z =�A=�"=�='�=�=g`==��=�~=:#=�=qT=�=�e=�=�X=@�	=�.=C�=K�===��=J��<�)�<��<��<"z�<h��<
,�<�x�<,��<���<'5�<�g�<���<��<5��<��<�$�<N@�<�Y�<�p�<j��<M��<C��<l��<�Ť<�Ѡ<�ۜ<e�<��<�<X��<���<���<j�<.z<�r<�j<'b<�1Z<�=R<�KJ<�[B<�m:<.�2<*<�"<��<��<<45<��;��;���;���;���;��;��;�x�;�v;�VX;.N:;�v;��:H��:%`�:��:��'9z폹Y�8��<��4y˺	�S���6�w�P�}�j�~��"���<֚��䦻e���$P�� �ɻ1�Ի^�߻dO� ���H����k�>H	��!���4������0$�+Q(�WZ,�LL0�	(4���7��;��@?��B��LF���I��M��pP�P�S��V�D+Z�NV]��x`�d�c���f�Ųi�/�l��o�دr�բu���x�.y{�]]~��������_y���䄼�N�����s ��>����[V������k"�������뒼�O�����g��hu��uՙ��4�������.N��&������d������T��}��[ۨ�:���������jX��f�������x��ٳ�19��{�������Z������K��Y|���  �  6�N=)N=uxM=d�L=�L=�cK=��J=��I=�KI=d�H=��G=v1G=~F=��E=YE=dD=��C=��B=�JB=�A=6�@=�.@=�y?=P�>=�>=�V==J�<=�;=�*;=�o:=��9=��8=}88=oy7=W�6=/�5=�55=r4=�3=>�2=�2="S1=e�0=A�/=v�.=�.=09-=X^,=�+=l�*=�)=��(=��'=1�&=��%=J%=;$=�"=m�!=�� =��=^�=s�=$f=H4=��=��=on=�=��=�\=��=f|=��=�z=g�=VZ
=�=d=&s=Y�=Z=SQ =;�<��<L��<�U�<��<���<9�<�t�<(��<	��<��<'�<{G�<
d�<�}�<��<=��<;��<<ʸ<uش<��<��<���<���<~�<�	�<@�<q�<f�<n�<�
�<e�<��<z<� r<��i<A�a<��Y<7�Q<��I<��A< :<�	2<�*<�"<.<�><S
<Ej<H�;�J�;Δ�;~��;WP�;UŦ;�K�;&�;�)q;b�R;To4;�\;.��:�:��u:�� :�kN8�˹��W�'&����ۺt	���$��t?�I�Y�!�s��Æ��X�������ѫ������Sû!�λF�ٻռ�aﻕ���>�����M��i~��������K"��{&�l�*�K�.��r2��@6���9���=��+A��D��H��tK�g�N��	R�uBU�TqX���[���^���a�1�d���g��j�+�m�b�p�/�s��v��y�M`|�:���Tq��Rك� @�����8���o��vԊ��8��d�������6c��Ƒ�'(������ꕼ�I��駘�S���a��4������%r��̠��%�����ڤ��4��,���쨼�H��ץ��s��ia������7���|��B۳��9�����Z����T��I�����Mq���  �  &�N=�(N=fxM=i�L=�L=�cK=��J=��I=�KI=��H=#�G=�1G=8~F=��E=~E=NdD=-�C=��B=�JB=-�A=L�@=�.@=z?=Y�>=�>=�V===�<=�;=�*;=�o:=|�9=`�8=N88=Fy7=*�6=��5=�55=�q4=Ƭ3=�2=�2=S1=U�0=4�/=p�.=�.=89-=k^,=0�+=z�*=�)=��(=��'=b�&=��%=q%=`$=:�"=��!=0� =��=��=��=1f=X4=��=��=gn=�=��=�\=��=2|=t�=�z=7�=Z
=��=2=�r="�=$=1Q =�<���<��<�U�<���<���<9�<u�<F��<P��<��<r'�<�G�<sd�<�}�<s��<���<���<�ʸ<�ش<#�<��<���< �<��<�	�</�<_�<P�<R�<p
�<�<U�<Zz<( r<��i<��a<��Y<l�Q<-�I<��A<�:<G	2<A*<["< .<?<%S
<}j<|�;fK�;��;���;�Q�;Ǧ;uM�;z�;o-q;�R;�r4;�_;h �:��:��u:�� :�N8��˹�W�x&����ۺ]t	���$�zv?�x�Y���s��Ć��Y��d����ҫ����UûS�λ�ٻ8��ua�����K����� ��~�h�>��p�OK"��z&���*�m�.�Hr2��?6���9�Κ=��*A���D�H�dtK�#�N�8	R�XBU�qX���[���^���a�t�d�)�g�-�j���m�.�p�Ƿs�۟v�˂y��`|��:�c���q���ك�>@�����R���o��UԊ�r8��C�������
c���ő��'��9����镼%I���������Ka��м������q���ˠ��%������٤��4�����'쨼�H����������a��	������}���۳��9��k�������,U������\��pq���  �  ��N=�(N=MxM=`�L=�L=dK=ڱJ='�I=1LI=�H=��G= 2G=�~F=a�E=E=�dD=��C=r�B=KB=��A=��@=8/@==z?=s�>=�>=zV==#�<=��;=�*;=Mo:=�9=��8=�78=�x7=��6=m�5=55=kq4=\�3=��2=02=�R1=�0=�/=X�.=�.=G9-=�^,=o�+=ɞ*=z�)=K�(=)�'=��&=;�%=%=�$=��"=�!=�� =�=�=Ȑ=if=y4=��=��=An=�=@�={\=C�=�{=��=&z=��=qY
=�=�=Qr=��=�=�P =5�<+��<���<bU�<��<���<Z9�<vu�<ߪ�<��<��<[(�<�H�<�e�<�~�<���<���<���<�˸<�ٴ<��<y�<Q��<h �<��<�	�<�<"�<��<��<�	�<C�<p�<4z<��q<z�i<9�a<�Y<r�Q<e�I<�A< :<�2<s*<�"<�-<)?<�S
<dk<��;xN�;]��;���;�U�;l˦;�R�;��;�7q;��R;�{4;�g;�:���:l�u:I� :ۇO8��˹�W��&����ۺ�w	��$��{?���Y�<�s�pȆ��]��o���s֫�˶��Xû"�λ��ٻ���cﻼ������������Y}�T�������I"�y&���*�A�.��o2��=6�{�9��=��(A��D�sH�sK��N��R�BU�qX�
�[�9�^���a���d���g���j�z�m�8�p�޹s��v� �y��b|��<�.	��nr��5ڃ��@��������!p��AԊ�C8��؛��V���Xb���đ�'��E����蕼H��r������E`��⻜����q��
ˠ�%��.���٤��4��)���Z쨼I��z���?��vb������p��~���ܳ�;��|�������V��j���"��r���  �  ��N=�(N=$xM=V�L=L=SdK=&�J=��I=�LI=��H=R�G=�2G=�F==�E=�E=�eD=��C=I�B=�KB=0�A=*�@=�/@=z?=��>=�>=gV==�<=�;=#*;=�n:=v�9=<�8=78=�w7=Ƿ6=��5=545=�p4=��3=��2=�2=MR1=��0=̶/=9�.=�.=o9-=�^,=ɀ+=>�*=�)=��(=��'=��&=�%=�%=�$=��"=��!=f� =��=e�=4�=�f=�4=��=��=n=,=˿=�[=��=�z=�=5y=��=vX
=�=�=^q=��=�=
P =�<0��<���<�T�<���<���<�9�<v�<���<��<��<�)�<J�<Cg�<���<f��<���<n��<7͸<۴<*�<�<��<� �<)�<�	�<��<��<(�<�
�<}�<��<��<��y<R�q<�i<��a<��Y<�Q<(�I<W�A<��9<E2<�*<�"<S-<\?<@T
<~l<e�;�R�;���;���;:]�;�Ҧ;Z�;d�;Gq;��R;b�4;�u;-(�:bѵ:y�u:�� :c�P8I�˹�W�)����ۺ�{	���$� �?��Y�C t��Ά�d��a����ܫ������]ûO�λ��ٻ��仌eﻘ������`��	��\|������y���F"��u&�3�*�ć.�kl2�:6��9�g�=��%A��D�)H�+qK���N��R�[AU��pX�}�[�B�^��a�e�d���g�u�j���m�c�p�X�s�b�v�W�y�hf|��?��
���s��Iۃ��A��1������Pp��/Ԋ��7��Y�������Ya���Ñ��%�������敼QF���������^��)���.���o���ɠ�,$���~��@٤�n4��6����쨼�I��/���4���c��F¯�!�����Z޳��<��0���j����W��⵺�X��s���  �  �N=(N=�wM=J�L=,L=�dK=��J=1 J=kMI=u�H=A�G=�3G=��F=c�E=E=�fD=��C=B C=�LB=�A=��@=50@=�z?=��>=>=XV==��<=�;=�);=n:=��9=N�8=68=�v7=��6=v�5=35=�o4=��3=!�2=�2=�Q1=E�0=u�/=�.=�.=�9-=_,=H�+=ݟ*=ź)=��(=��'=��&=,�%=�%=�$=� #=��!=L� =��=�=ő=(g=�4=��=k�=�m=�=0�=)[=��=�y=��=x=I�=W
=��=E=/p=��=�
=O =��<��<��<}T�<���<���<*:�<w�<߬�<���<��<�+�<�L�<�i�<��<���<ԭ�<���<4ϸ<�ܴ<��<��<��<��<��<�	�<��<��<1�<h	�<��<��<� �<��y<��q<"�i<��a<k�Y<��Q<,�I<��A<��9<�2<�*<�"<�,<�?<5U
<+n<!�;�X�;��;���;�e�;uܦ;-d�;���;�[q;��R;��4;G�;�H�:��:xv::�R8��˹!�W��+��p�ۺ^�	��$��?��Z�
t�7ֆ�Jl���Ɵ��䫻ķ��dû��λ��ٻ\���h�����7��A��A���z���W��Q��(C"��q&��*�3�.��g2�m56�p�9��=��!A�p�D� H��nK�t�N�?R��@U��pX���[�v�^���a���d���g���j�X�m�\�p���s���v��y��j|��C����du���܃��B��������pp��Ԋ�n7������h���`��!��#�������䕼D��a�������R\�����N���m���Ƞ��"���}���ؤ�.4��I����쨼fJ��1������9e��	į��"�������೼
?��p���}����Y���������~t���  �  [�N=�'N=�wM=4�L=HL=�dK=�J=� J=BNI=f�H=]�G=75G=��F=��E=rE=1hD=ߴC=|C=�MB=�A=��@=�0@=^{?="�>=>=6V==g�<=��;=�(;=Am:=��9=5�8=�48=�u7=]�6=%�5=�15=Pn4=v�3=�2=�2=�P1=��0=�/=��.=�.=�9-=x_,=Ё+=��*=��)=��(= �'=��&=m�%=G%=3$=�#=�!=l� =r�=�=j�=�g=*5=��=K�=ym=<=|�=>Z=��=�x=��=�v=��=�U
=)�=�=�n=<�=�	=N =��<���<��<�S�<H��<��<�:�<�w�<:��<C��<��<&.�<O�<'l�<Ʌ�<|��<w��<%¼<�Ѹ<
ߴ<��<U��<L��<p�<��<�	�<1�<6�< 
�<��<�<��<\��<�y<K�q<��i<T�a<��Y<{�Q<}�I<��A<�9<� 2<*<p"<@,<�?<;V
<p<H�;n_�;׭�;P�;up�;��;�o�;�
�;Ssq;q�R;9�4;w�;�l�:�:�:v:�F:�YT8^i˹S�W�'/����ۺ��	�A�$�̛?�UZ��t��߆��u���П�>�ͷ��mû+�λ�ٻ����l�?��������d��Iy�V�Y�����?"�.m&��*��}.�Sb2�06�6�9� �=��A�h�D�dH��kK�8�N��R��?U��pX���[�ҷ^��a���d�I�g���j���m�~�p���s�.�v��y��o|��H����Ow��`ރ�5D��������p�� Ԋ��6������<���w^��M����!��B���J╼hA����������Y������
��l���Ơ��!���|��ؤ��3��e���w�&K��m�����g��!Ư�R%��V���㳼�A��������� \��͹�����	v���  �  ��N=:'N=^wM=&�L=mL=3eK=��J=�J=)OI=m�H=��G=~6G=P�F=#�E=�E=�iD=6�C=�C=�NB=�A=��@=o1@=�{?=e�>=;>=V==	�<=�;=)(;=bl:=��9=
�8=�38=1t7=�6=��5=w05=�l4=G�3=��2=2=#P1=�0=��/=��.=�.=�9-=�_,=Z�+=M�*=��)=��(=2�'=4�&=� &=�%=�$=D#=Y�!=�� =r�=̶=�=h=n5=��=3�=m=�=��=KY=y�=Sw=*�=�t=1�=�S
=~�=&=+m=ѽ=E=�L =��<��<���< S�<��<;��<];�<�x�<���<��<�
�<�0�<�Q�<�n�<���<a��<I��<�ļ<Ը<A�<��<���<{��<;�<_�<�	�<�
�<Q
�<��<J�<
�<t��<���<~�y<k�q<W�i<U�a<�Y< �Q<^�I<�A<X�9<��1<�
*<�"<�+<!@<LW
<r<� �;�f�;o��;A�;n{�;N�;N|�;�;ǌq;�S;��4;�;p��:�/�:5pv:q:BV8�@˹	�W��4��� ܺ��	���$�Ϫ?��"Z��1t�v醻���F۟������׷�Uvû��λ�ٻp�仝q�J���������w���w���4������:"�4h&��|*�Vx.��\2�Q*6���9�Ԇ=��A��D��H�vhK��N�	R�?U��pX�|�[�}�^���a���d��g�k�j���m���p�=�s��v���y�Du|��M����y��*����E��$������q���ӊ�6��՘������\��R���g������ߕ��>��眘�H���W���������i���Ġ�< ���{��bפ��3��s���L��ͪ���	��i��tȯ��'������峼�D��â��� ��s^��!�������w���  �  �N=�&N=wM=�L=L=�eK=�J=7J=�OI=z�H=��G=�7G=��F=��E=ME= kD=��C=�C=#PB=�A=N�@=2@=I|?=��>=?>=�U==��<=��;=t';=uk:=��9=��8=D28=�r7=��6=J�5=/5=�k4=�3=��2=2=NO1=t�0==�/=d�.=�.=:-=5`,=�+=	�*=t�)=��(=Y�'=v�&= &=%=�$=�#=��!=�� =��=��==�h=�5=��=��=�l==�=NX=N�=v=��=os=��=@R
=ն=�=�k=\�=�=�K =��<���<���<eR�<���<k��<�;�<�y�<��<���<��<�2�<HT�<�q�<���<B��<��<rǼ<�ָ<��<{�<���<���<�<��<�	�<:
�<v	�<p�<��< �<��<8��<��y<r�q<_�i<E�a<.�Y<��Q<C�I<��A<U�9<��1<M*<K"<�*<5@<}X
<t<j&�;�m�;L��;0�;��;��;���;�#�;Υq;M-S;�4;��;��:P�:f�v:��:�:X8�$˹
�W�W9���ܺf�	���$��?��3Z��Dt�}�y����埻���᷻�û�λb�ٻ����u�(���Q���������u�������*6"�gc&�[w*��r.��V2��$6���9���=�>A�w�D��H�meK�|�N�aR�?>U��pX�O�[��^���a�
�d���g���j���m��p���s���v�c�y��z|�)S�����{��	⃼+G��9������gq���ӊ��5�������9[��c�����_}���ܕ��;�����v���ST������T���g��Cà����~z���֤�g3�������M�����p��k���ʯ�G*�������購gG������{���`��t������xy���  �  ^�N=?&N=�vM=��L=�L=�eK=��J=�J=�PI=f�H=��G=�8G=��F=��E=�E=BlD=ظC=#C=.QB=֜A=�@=�2@=�|?=��>=I>=�U==`�<=	�;=�&;=�j:=��9=��8=18=�q7=2�6=��5=�-5=kj4=Х3=��2=2=�N1=߂0=ʴ/=,�.=�.=>:-=�`,=d�+=��*=C�)=��(=r�'=��&=\&=N	%=9
$=�#=��!=�� =o�=g�=g�=�h=�5=��=ٷ=hl=�=4�=bW=9�=�t=O�=�q=	�=�P
=F�==)j=��=�=�J =�<��<���<�Q�<x��<���<r<�<�z�<^��<w��<��<!5�<�V�<@t�<8��<ܤ�<���<ʼ<�ظ<��<1�<���<���<��<�<�	�<�	�<��<;�<��<��<���<���<��y<��q<��i<��a<��Y<@�Q<t�I<[�A<��9<��1<�*<�"<D*<h@<nY
<�u<�+�;Dt�;��;Q%�;���;T
�;ғ�;�/�;��q;�DS;��4;��;���:�n�:��v:��:v�Y8_˹D�W�^>��8ܺɤ	�K�$�4�?��CZ��Vt�����_��������귻Ɉû��λ"ڻ-��z�K���������˾�t�r������/2"��^&�5r*��m.��Q2�B6���9�h|=��A�x�D�h H�ybK�e�N� R�x=U��pX��[���^��a��d�x�g���j�X�m���p��s��v���y��|�X�����}���ー�H��K���R���q���ӊ��5��8��������Y������	��{��`ڕ�J9��`��������Q�����(
���e������l���y��֤�+3��ڐ��屮�M��K������l���̯��,��:���`볼J��@�����vc���������${���  �  ��N=�%N=�vM=��L=�L=fK=�J=fJ=zQI=3�H=��G=�9G=�F=��E=� E=_mD=ݹC=C=RB=��A=��@=63@=}?=�>=P>=�U==�<=��;=)&;=�i:=��9=��8=08=np7=
�6=��5=�,5=Yi4=ۤ3=��2=O2=�M1=S�0=l�/=��.=�.=N:-=�`,=Ӄ+=Q�*=��)=��(=`�'=��&=j&=j
%=U$=�#=��!=�� =7�=�=�=\i=%6=��=��=l==��=�V=F�=�s=0�=�p=��=ZO
=�=�=�h=ڹ=�=�I =w�<���<���<%Q�<>��<���<�<�<�{�<���<���<��<�6�<�X�<sv�<���<+��<��<̼<�ڸ<J�<��<0��<� �<Y�<B�<�	�<Y	�<��<�<��<d��<���<��<�y<�q<��i<��a<�Y<��Q<b�I<��A<t�9<��1<�*<�"<�)<z@<3Z
<6w<0�;z�;���;-�;��;t�;���;�9�;��q;uWS;�	5;�;'��: ��:�w:I�:8[8��ʹj�W�}C��"ܺ��	�K�$���?�QQZ�ret���󜓻N���^�����û��λ'ڻ
��	~�����������_��Hs����������."��Z&�7n*�@i.��L2��6���9�jx=��
A��D�f�G�`K���N���Q�=U�	qX�ܛ[��^�+�a���d���g�s�j�%�m�8�p���s���v�[�y�k�|�D\����e��O僼�I��J������r���ӊ�F5����������nX�����S��y��\ؕ�7������򙼢O��'���P��Rd��@���W���x���դ�3�� ����屮�N��p���n���n���ί��.��e�����eL������4��te���º�z���|���  �  W�N=�%N=RvM=��L=�L=,fK=;�J=�J=�QI=ϟH=i�G=�:G=ևF=��E=�!E=;nD=��C=�C=�RB=4�A=2�@=�3@=R}?=6�>=V>=�U==ۛ<=>�;=�%;=Si:=�9= �8=$/8=�o7=.�6=��5=�+5=wh4=�3=+�2=�2=aM1=�0=-�/=��.=�.=g:-=a,=*�+=��*=��)=`�(=�'=o�&=B&=9%=!$=�#=��!=c� =��=��=L�=�i=S6=�=��=�k=�=
�=�U=��=�r=?�=�o=��=XN
=�=�=�g=�=�=I =K�<ͅ�<"��<�P�<��<���<V=�<B|�<O��<���<��<�8�<iZ�<-x�<1��<��<���<�ͼ<[ܸ<��<��<��<e�<��<u�<�	�<��<C�<A�<� �<��<t��<��<c�y<p�q<�i<�a<G�Y<C�Q<�I<��A<'�9<��1<�*<�"<>)<�@<�Z
<~x<3�;Y~�;��;g3�;Ο�;��;8��;(A�;��q;9fS;15;y�;��:��:h%w:��:H<\8��ʹ��W�G��6)ܺh�	�k�$��?�M\Z�*rt�m��\��������������%�û�λ�ڻ�����ﻊ���Q�������>r�
���M��,"��W&�k*��e.��I2�M6��9�8u=��A�Y�D�&�G�U^K�,�N���Q��<U�qX���[��^���a���d���g�H�j�a�m���p��s��v�ͪy�܇|��_�M������e惼�J������`��Tr���ӊ�5�����������W�������w���֕�]5��q������M���������c��7������#x��Dդ��2�� ����WO��J���r���o��;Я�c0��'���`ﳼN��C����	��'g��ĺ�� ���}���  �  
�N=K%N=2vM=��L=�L=EfK=c�J=	J=RRI=3�H=��G=';G=\�F=Q�E=&"E=�nD=1�C=OC=*SB=��A=��@=�3@=v}?=O�>=[>=zU==��<=��;=d%;=�h:=��9=��8=�.8=o7=��6=U�5=1+5=�g4=��3=��2=P2=
M1=��0=��/=��.=�.=z:-=a,=[�+=�*=޿)=��(=~�'=��&=�&=�%=�$=2#=�!=�� =4�=�=��=�i=g6=�=��=�k=v=��=�U=�=pr=��=/o=�=�M
=A�==`g=d�=j=�H =��<*��<���<fP�<���<���<�=�<�|�<��<���<��<R9�<m[�<:y�<Q��< ��<���<�μ<1ݸ<q�<��<���<��<�<��<p	�<��<��<��<���<L��<���<��<U�y<�q<��i<��a<%�Y<:�Q<C�I<�A<��9<��1<�*< "<�(<�@<5[
<&y<^5�;B��;g��;�6�;ȣ�;M�;�;!F�;t�q;�oS;* 5;��;l �:��:`:w::��\8�ʹ
�W��I��n/ܺ��	� �$���?��bZ��xt�N��ǧ��T��
 �����Ùû�λ�ڻC�����������������q�=	�������|*"�LV&��h*��c.�[G2�6���9�+s=�*A�̇D���G�]K�P�N�V�Q�Q<U�/qX�ߜ[���^���a���d���g���j�I�m���p�7�s�^�v�%�y���|��a�;������4烼`K��z������qr���ӊ��4������j����V��,��� ���v���Օ�P4��T�����L������
��Jb���������w��դ��2��:���>��O��⯫�.���p��ѯ�U1�� �����NO��n����
��h���ĺ��!��S~���  �  �N=9%N=&vM=��L=�L=TfK=r�J=J=dRI=[�H=��G=U;G=��F=}�E=Y"E=�nD=a�C=|C=VSB=��A=��@=�3@=�}?=Z�>=Q>=mU==��<=��;=X%;=�h:=�9=Y�8={.8=�n7=n�6=1�5=�*5=�g4=Z�3=��2='2=�L1=��0=�/=��.=�.={:-=)a,=g�+=�*=��)=��(=��'=�&=�&=�%=�$=U#=1�!=�� =]�=�=��=�i=p6=
�=w�=�k=^=��=�U=��=Cr=w�=�n=��=�M
=�=�=)g=,�=>=rH =b�<���<���<MP�<ާ�<���<�=�<�|�<��<���<��<�9�<�[�<�y�<���<\��<��<ϼ<�ݸ<��<��<���<��< �<��<M	�<��<��<��<���<���<8��<y�<��y<2�q<��i<��a<N�Y<j�Q<��I<]�A<�9<��1<J*<�"<�(<�@<x[
<iy<�5�;���;���;Z8�;Z��;� �;{��;�G�;L�q;�rS;J#5;�;`%�:���:�>w::_]8o�ʹ��W�qK��j1ܺD�	���$�:�?�fZ�|t������o���!������b�ûH�λ�ڻ���d�ﻁ������8��u���q�		�f��r���)"��U&�6h*�c.��F2�K6�S�9�ar=�sA��D�C�G��\K��N�$�Q�H<U�iqX���[��^��a��d�*�g�u�j��m�]�p��s���v�ʭy�׊|�_b����ց��y烼{K����������r���ӊ��4������K����V�������^v��YՕ�4��푘���L��H�������a��^�������w���Ԥ��2��[���R��O������\���p��gѯ��1�������𳼙O��ϭ��U��{h��7ź��!���~���  �  
�N=K%N=2vM=��L=�L=EfK=c�J=	J=RRI=3�H=��G=';G=\�F=Q�E=&"E=�nD=1�C=OC=*SB=��A=��@=�3@=v}?=O�>=[>=zU==��<=��;=d%;=�h:=��9=��8=�.8=o7=��6=U�5=1+5=�g4=��3=��2=P2=
M1=��0=��/=��.=�.=z:-=a,=[�+=�*=޿)=��(=~�'=��&=�&=�%=�$=2#=�!=�� =4�=�=��=�i=h6=�=��=�k=w=��=�U=�=sr=��=3o=�=�M
=F�==fg=k�=q=�H =��<:��<���<vP�<	��<���<�=�<�|�<��<���<��<Y9�<r[�<=y�<R��<���<���<�μ<*ݸ<i�<��<���<��<��<��<c	�<��<��<��<���<C��<���<��<M�y<�q<��i<��a<,�Y<F�Q<R�I<�A<��9<��1<�*<"<)<�@<N[
<>y<�5�;k��;���;�6�;ݣ�;Z�;���;F�;\�q;doS;�5;��;��:K��:�8w:?	:�\8J�ʹ0�W��J���0ܺ.�	���$�?�?�kcZ�syt�����������4 ��3����û#�λ�ڻ[����������������q�A	�������~*"�MV&��h*��c.�\G2�6���9�,s=�*A�̇D���G�]K�P�N�V�Q�Q<U�/qX�ߜ[���^���a���d���g���j�I�m���p�7�s�^�v�%�y���|��a�;������4烼`K��z������qr���ӊ��4������j����V��,��� ���v���Օ�P4��T�����L������
��Jb���������w��դ��2��:���>��O��⯫�.���p��ѯ�U1�� �����NO��n����
��h���ĺ��!��S~���  �  W�N=�%N=RvM=��L=�L=,fK=;�J=�J=�QI=ϟH=i�G=�:G=ևF=��E=�!E=;nD=��C=�C=�RB=4�A=2�@=�3@=R}?=6�>=V>=�U==ۛ<=>�;=�%;=Si:=�9= �8=$/8=�o7=.�6=��5=�+5=wh4=�3=+�2=�2=aM1=�0=-�/=��.=�.=g:-=a,=*�+=��*=��)=`�(=�'=o�&=B&=9%="$=�#=��!=c� =��=��=M�=�i=U6=�=��=�k=�=�=V=��=�r=F�=�o=��=bN
=��=�=�g=��=�="I =i�<��<A��<�P�</��<���<q=�<[|�<e��<��<��<�8�<rZ�<2x�<2��<��<���<�ͼ<Mܸ<��<��<���<N�<��<\�<l	�<��<,�<+�<o �<��<f��<��<T�y<h�q<�i<�a<V�Y<Y�Q<;�I<��A<O�9<+�1<�*<�"<q)<�@<[
<�x<i3�;�~�;U��;�3�;���;��;B��;"A�;��q;�eS;�5;��;��:���:"w:$�:��[8��ʹۖW�(I��Q+ܺs�	�o�$��?�=]Z�st��������1���$������h�ûA�λ�ڻ���'�ﻭ���`�������Hr�
���R��,"��W&�k*��e.��I2�O6��9�:u=��A�Y�D�&�G�V^K�,�N���Q��<U�qX���[��^���a���d���g�H�j�a�m���p��s��v�ͪy�܇|��_�M������e惼�J������`��Tr���ӊ�5�����������W�������w���֕�]5��q������M���������c��7������#x��Dդ��2�� ����WO��J���r���o��;Я�c0��'���`ﳼN��C����	��'g��ĺ�� ���}���  �  ��N=�%N=�vM=��L=�L=fK=�J=fJ=zQI=3�H=��G=�9G=�F=��E=� E=_mD=ݹC=C=RB=��A=��@=63@=}?=�>=P>=�U==�<=��;=)&;=�i:=��9=��8=08=np7=
�6=��5=�,5=Yi4=ۤ3=��2=O2=�M1=S�0=l�/=��.=�.=N:-=�`,=Ӄ+=Q�*=��)=��(=`�'=��&=j&=j
%=U$=�#=��!=�� =8�=�=�=^i='6=��=��=l==��=�V=M�=�s=9�=�p=��=hO
=��=�= i=�=�=�I =��<��<���<PQ�<h��<���<=�<�{�<���<���<��<7�<�X�<{v�<���<(��<��<̼<�ڸ<3�<��<��<� �<7�<�<u	�<7	�<��<��<m�<K��<���<��<��y<�q<��i<��a<�Y<
�Q<��I<��A<��9<=�1<>*<�"<�)<�@<yZ
<yw<�0�;�z�;?��;h-�;E��;��;ɝ�;�9�;O�q;WS;.	5;>�;P��:��:8w:*�:��Z8`�ʹG�W�wF��%ܺ�	���$�5�?��RZ��ft��������������F�L�û��λrڻK��B~����������n��Ts����������."��Z&�;n*�Di.��L2��6���9�kx=��
A��D�g�G�`K���N���Q�=U�	qX�ܛ[��^�+�a���d���g�s�j�%�m�8�p���s���v�[�y�k�|�D\����e��O僼�I��J������r���ӊ�F5����������nX�����S��y��\ؕ�7������򙼢O��'���P��Rd��@���W���x���դ�3�� ����屮�N��p���n���n���ί��.��e�����eL������4��te���º�z���|���  �  ^�N=?&N=�vM=��L=�L=�eK=��J=�J=�PI=f�H=��G=�8G=��F=��E=�E=BlD=ظC=#C=.QB=֜A=�@=�2@=�|?=��>=I>=�U==`�<=	�;=�&;=�j:=��9=��8=18=�q7=2�6=��5=�-5=kj4=Х3=��2=2=�N1=߂0=ʴ/=,�.=�.=>:-=�`,=d�+=��*=C�)=��(=r�'=��&=]&=N	%=:
$=�#=��!=�� =p�=h�=i�= i=�5=�=ݷ=ml=�=;�=jW=B�=�t=[�=
r=�=�P
=X�==>j=�=�=�J =C�<B��<���<�Q�<���<���<�<�<{�<���<���<�<75�<�V�<It�<:��<ؤ�<���<�ɼ<�ظ<s�<�<���<���<��<��<�	�<�	�<d�<�<��<���<���<���<��y<��q<��i<��a<��Y<f�Q<��I<��A<��9<��1<J*<3"<�*<�@<�Y
<�u<T,�;�t�;���;�%�;쐶;�
�;㓗;�/�;=�q;GDS;7�4;��;���: l�:��v:��:��Y8U˹s�W�B���ܺ��	��$���?��EZ�Xt�����
���=�c��Q뷻>�û$�λ~ڻ~��Qzﻇ����� ��޾��t�������72"��^&�;r*��m.��Q2�E6���9�j|=��A�y�D�i H�zbK�f�N� R�x=U��pX��[���^��a��d�x�g���j�X�m���p��s��v���y��|�X�����}���ー�H��L���R���q���ӊ��5��8��������Y������	��{��`ڕ�J9��`��������Q�����(
���e������l���y��֤�+3��ڐ��屮�M��K������l���̯��,��:���`볼J��@�����vc���������${���  �  �N=�&N=wM=�L=L=�eK=�J=7J=�OI=z�H=��G=�7G=��F=��E=ME= kD=��C=�C=#PB=�A=N�@=2@=I|?=��>=?>=�U==��<=��;=t';=uk:=��9=��8=D28=�r7=��6=J�5=/5=�k4=�3=��2=2=NO1=t�0==�/=d�.=�.=:-=5`,=�+=
�*=t�)=��(=Y�'=v�&= &=%=�$=�#=��!=�� =��=��=ē=�h=�5=��=�=�l==��=WX=X�=v=��=~s=��=RR
=�=�=�k=v�==�K =�<���<��<�R�<���<���</<�<)z�<:��<���<�<�2�<YT�<�q�<���<=��<��<_Ǽ<yָ<n�<W�<X��<���<��<��<�	�<

�<I	�<F�<e�<� �< ��<#��<��y<c�q<^�i<S�a<K�Y<��Q<{�I<��A<��9<��1<�*<�"<N+<�@<�X
<ft<'�;en�;ο�;��;f��;K��;���;�#�;w�q;�,S;2�4;��;���:6M�:��v:��:�W8$4˹�W�g=���ܺh�	���$��?�~5Z�\Ft�K�8���j査���ⷻ.�ûw�λ��ٻ���1v�k���n��������u�������36"�nc&�aw*��r.��V2��$6��9���=�@A�x�D��H�neK�}�N�aR�?>U��pX�O�[��^���a�
�d���g���j���m��p���s���v�c�y��z|�)S�����{��	⃼+G��9������gq���ӊ��5�������9[��c�����_}���ܕ��;�����v���ST������T���g��Cà����~z���֤�h3�������M�����p��k���ʯ�G*�������購gG������{���`��t������xy���  �  ��N=:'N=^wM=&�L=mL=3eK=��J=�J=)OI=m�H=��G=~6G=P�F=#�E=�E=�iD=6�C=�C=�NB=�A=��@=o1@=�{?=e�>=;>=V==	�<=�;=)(;=bl:=��9=
�8=�38=1t7=�6=��5=w05=�l4=G�3=��2=2=#P1=�0=��/=��.=�.=�9-=�_,=Z�+=M�*=��)=��(=2�'=5�&=� &=�%=�$=E#=Y�!=�� =s�=Ͷ=�=h=q5=��=8�="m=�=��=TY=��=_w=8�=u=B�=�S
=��=>=Dm=�=a=M =�<C��<,��<]S�<Y��<t��<�;�<y�<��<:��<�
�<�0�<�Q�<o�<���<\��<=��<�ļ<Ը< �<w�<���<M��<�<-�<�	�<
�<"
�<�<"�<��<X��<���<`�y<[�q<W�i<d�a<"�Y<L�Q<��I<R�A<��9<��1<�
*<1"<#,<�@<�W
<cr<X!�;}g�;���;��;�{�;��;b|�;�;m�q;KS;��4;ݯ;א�:�,�:�iv:�i:��U8�P˹U�W��8���ܺՕ	���$�Ŭ?��$Z��3t�Kꆻ΀���۟�/���5ط��vû4�λ�ٻ����qﻐ�������������w��A������:"�;h&��|*�[x.��\2�T*6���9�ֆ=� A��D��H�whK��N�
R�?U��pX�}�[�}�^���a���d��g�k�j���m���p�=�s��v���y�Du|��M����y��*����E��$������q���ӊ�6��՘������\��R���g������ߕ��>��眘�H���W���������i���Ġ�< ���{��bפ��3��s���L��ͪ���	��i��tȯ��'������峼�D��â��� ��s^��!�������w���  �  [�N=�'N=�wM=4�L=HL=�dK=�J=� J=BNI=f�H=]�G=75G=��F=��E=rE=1hD=ߴC=|C=�MB=�A=��@=�0@=^{?="�>=>=6V==g�<=��;=�(;=Am:=��9=5�8=�48=�u7=]�6=%�5=�15=Pn4=v�3=�2=�2=�P1=��0=�/=��.=�.=�9-=x_,=Ё+=��*=��)=��(= �'=��&=m�%=G%=3$=�#=�!=m� =s�=�=l�=�g=,5=��=O�=~m=B=��=GZ=��=�x=��=�v=��=�U
=>�=�=�n=U�=�	=/N =��<ӌ�<W��<	T�<���<H��< ;�<!x�<e��<i��<��<?.�<O�<2l�<̅�<x��<k��<¼<�Ѹ<�޴<z�<,��< ��<A�<��<�	�<�<	�<�	�<��<��<��<G��<��y<<�q<��i<c�a<��Y<��Q<��I<��A<f�9<(2<d*<�"<�,<)@<�V
<up<��;`�;Y��;��;�p�;��;�o�;�
�;�rq;��R;f�4;l�;j�:+
�: 4v:�?:��S8�x˹V�W�83����ۺ��	�8�$���?�%Z��!t�\���ev��<џ��Tη�nû��λm�ٻ(��Cmﻂ������3��y��Zy�e�f�����&?"�5m&��*�~.�Wb2�06�9�9�"�=��A�i�D�eH��kK�9�N��R��?U��pX���[�ҷ^��a���d�I�g���j���m�~�p���s�.�v��y��o|��H����Ow��`ރ�5D��������p�� Ԋ��6������<���w^��M����!��B���J╼hA����������Y������
��l���Ơ��!���|��ؤ��3��e���w�&K��m�����g��!Ư�R%��V���㳼�A��������� \��͹�����	v���  �  �N=(N=�wM=J�L=,L=�dK=��J=1 J=kMI=u�H=A�G=�3G=��F=c�E=E=�fD=��C=B C=�LB=�A=��@=50@=�z?=��>=>=XV==��<=�;=�);=n:=��9=N�8=68=�v7=��6=v�5=35=�o4=��3=!�2=�2=�Q1=E�0=u�/=�.=�.=�9-=_,=H�+=ݟ*=ź)=��(=��'=��&=,�%=�%=�$=� #=��!=L� =��=�=Ƒ=+g=�4=��=o�=�m=�=6�=1[=��=�y=��=x=X�=0W
=��=Y=Ep=��=�
=5O =��<(��<T��<�T�<���<��<X:�<-w�<��<���<��<�+�<�L�<�i�<��<���<ɭ�<���<ϸ<�ܴ<��<��<���<~�<]�<�	�<g�<��<�<F	�<��<��<� �<h�y<��q<"�i<��a<��Y<��Q<^�I< �A<��9<2<J*<!"<9-<�?<�U
<|n<��;
Y�;g��;E��;&f�;�ܦ;>d�;���;P[q;�R;М4;W�;FF�:2�:� v:�:@$R8��˹P�W�]/���ۺ+�	�Ϲ$���?��Z��t��ֆ��l��wǟ�~嫻�ķ�aeû�λ��ٻ���4i����Q��X��T��{���c��Z��0C"��q&���*�7�.��g2�p56�s�9� �=��!A�q�D�H��nK�t�N�@R��@U��pX��[�w�^���a���d���g���j�X�m�\�p���s���v��y��j|��C����du���܃��B��������pp��Ԋ�n7������h���`��!��#�������䕼D��a�������R\�����N���m���Ƞ��"���}���ؤ�.4��I����쨼fJ��1������9e��	į��"�������೼
?��p���}����Y���������~t���  �  ��N=�(N=$xM=V�L=L=SdK=&�J=��I=�LI=��H=R�G=�2G=�F==�E=�E=�eD=��C=I�B=�KB=0�A=*�@=�/@=z?=��>=�>=gV==�<=�;=#*;=�n:=v�9=<�8=78=�w7=Ƿ6=��5=545=�p4=��3=��2=�2=MR1=��0=̶/=9�.=�.=o9-=�^,=ɀ+=>�*=�)=��(=��'=��&=�%=�%=�$=��"=��!=g� =��=f�=5�=�f=�4=��=��=n=0=п=�[=��=�z=�=@y=��=�X
=�=�=pq=��=�=P =I�<[��<)��<U�<��<���<�9�<?v�<٫�<8��<�<*�<�J�<Kg�<À�<c��<���<a��<$͸< ۴<�<a�<���<� �<�<�	�<��<w�<	�<�
�<e�<��<��<��y<G�q<�i<��a< �Y<%�Q<P�I<��A<��9<�2</*<-"<�-<�?<�T
<�l<��;S�;
��;E��;s]�;Ӧ;%Z�;[�;�Fq;_�R;Ȋ4;u;W&�:Eϵ:��u:�� :2�P8��˹��W�,����ۺb}	��$�c�?�d�Y��t�'φ��d��⾟�Gݫ����/^û��λI�ٻ����e��������s����i|���������F"��u&�7�*�Ǉ.�nl2�!:6��9�h�=��%A��D�)H�+qK���N��R�[AU��pX�}�[�B�^��a�e�d���g�u�j���m�c�p�X�s�b�v�W�y�hf|��?��
���s��Iۃ��A��1������Pp��/Ԋ��7��Y�������Ya���Ñ��%�������敼QF���������^��)���.���o���ɠ�,$���~��@٤�n4��6����쨼�I��/���4���c��F¯�!�����Z޳��<��0���j����W��⵺�X��s���  �  ��N=�(N=MxM=`�L=�L=dK=ڱJ='�I=1LI=�H=��G= 2G=�~F=a�E=E=�dD=��C=r�B=KB=��A=��@=8/@==z?=s�>=�>=zV==#�<=��;=�*;=Mo:=�9=��8=�78=�x7=��6=m�5=55=kq4=\�3=��2=02=�R1=�0=�/=X�.=�.=G9-=�^,=o�+=ɞ*=z�)=K�(=)�'=��&=<�%=%=�$=��"=�!=�� =�=�=ɐ=jf=z4=��=��=Dn=�=D�=�\=I�=�{=��=.z=��={Y
=�=�=]r=��=�=�P =S�<J��<���<�U�<��<���<u9�<�u�<���<��<��<h(�<�H�<�e�<�<���<���<���<�˸<�ٴ<��<d�<:��<P �<��<�	�<��<
�<��<��<�	�<5�<e�<$z<��q<z�i<@�a<��Y<��Q<��I<6�A<7 :<+2<�*<�"<�-<\?<�S
<�k<0�;�N�;���;���;V�;�˦;�R�;��;�7q;��R;x{4;=g;��:8��:�u:�� :/JO8��˹4�W��(����ۺ�x	��$��|?���Y��s��Ȇ�H^��ʸ���֫����UXû]�λ�ٻ���Gc��������������b}�\��������I"�y&���*�C�.��o2��=6�}�9��=��(A��D�tH�sK��N��R�BU�qX�
�[�9�^���a���d���g���j�z�m�8�p�޹s��v� �y��b|��<�.	��nr��5ڃ��@��������!p��AԊ�C8��؛��V���Xb���đ�'��E����蕼H��r������E`��⻜����q��
ˠ�%��.���٤��4��)���Z쨼I��z���?��vb������p��~���ܳ�;��|�������V��j���"��r���  �  &�N=�(N=fxM=i�L=�L=�cK=��J=��I=�KI=��H=#�G=�1G=8~F=��E=~E=NdD=-�C=��B=�JB=-�A=L�@=�.@=z?=Y�>=�>=�V===�<=�;=�*;=�o:=|�9=`�8=N88=Fy7=*�6=��5=�55=�q4=Ƭ3=�2=�2=S1=U�0=4�/=p�.=�.=89-=k^,=0�+=z�*=�)=��(=��'=b�&=��%=q%=`$=:�"=��!=1� =��=��=��=1f=Y4=��=��=hn=�=��=�\=��=5|=w�=�z=;�=Z
=��=8=�r=)�=+=8Q =�<ϐ�<-��<�U�<��<���< 9�<u�<R��<Z��<��<y'�<�G�<vd�<�}�<r��<���<���<�ʸ<�ش<�<��<���< �<��<�	�<#�<R�<E�<H�<g
�<�<O�<Rz<$ r<��i<��a<��Y<x�Q<<�I<��A<�:<^	2<Z*<t"<.</?<?S
<�j<��;�K�;3��;��;R�;Ǧ;zM�;w�;X-q;ƸR;�r4;�_;���:G��:�u:�� :�N8�˹�W��'����ۺ�t	�*�$��v?���Y�
�s��Ć�0Z�������ҫ�7���?Uûr�λ0�ٻP�今a�����R�����%��~�l�B��s�RK"��z&���*�o�.�Ir2��?6���9�Κ=��*A���D�H�dtK�#�N�8	R�YBU�qX���[���^���a�t�d�)�g�-�j���m�.�p�Ƿs�۟v�˂y��`|��:�c���q���ك�>@�����R���o��UԊ�r8��C�������
c���ő��'��9����镼%I���������Ka��м������q���ˠ��%������٤��4�����'쨼�H����������a��	������}���۳��9��k�������,U������\��pq���  �  �N=�0N=$�M=��L=$ L=�nK=�J=�
J=aXI=��H=��G=3@G=��F=Q�E=_)E=swD=��C=�C=/cB=��A=��@=�M@=�?=��>=N3>=+~==��<=�<=�X;=��:=��9=�*9=7o8=��7=�6=�66=�v5=H�4=6�3=�03=]k2=0�1=��0=0=�@/=po.=+�-=��,=��+=]
+=>(*=iB)=�X(=�j'=�x&=�%=��$=4�#=p�"=�t!=�b =J=Y*=�=��=�=�[=�=��= f=	=�=o= �=3=2�=P�
=�U	=��==�O=��=c� =��<���<���<:�<���<R��<���<�1�<�\�<���<��<��<���<3��<'��<K�<~�<�<%�<�,�<p2�<�6�<�9�<;�<�:�<�8�<%5�<0�<�)�<_"�<"�<\�<$�<��y<��q<��i<{�a<�Y<[�Q<��I<��A<}�9<��1<A�)<�!<��<�<%�	<��<�L�;k�;6��;���;��;�^�;�Ô;�=�;!�k;�L;{].;n;D��:��:8xY:�Z�9 �����s�w�B������E0�I�-�۩H�tRc�ۏ}�4����Y���Ǥ����e弻G�ȻF�ӻ�$߻�	����D��p���	�`\�d����i��{ �»$���(��,��0�A�4��n8�<�#�?��'C��F���I��;M��zP���S���V�n�Y�(
]�o`�5c�>f��i�l���n�1�q�K�t� �w��wz�K}����r��ׂ�H:��Y�������	_��￉�!������ ㍼D���������e���Ĕ�#��]����ۘ��6��L����蜼$@��������D��㚣�"�J��ˢ��_����V���������.j���Ư��#������`ݳ��9��������SO������{���e���  �  ��N=�0N=�M=��L=0 L=�nK=/�J=J=�XI=�H=%�G=q@G=�F=��E=})E=�wD=4�C=�C=icB=�A=$ A=�M@=*�?=��>=X3>=~==��<=�<=�X;=��:=��9=�*9=o8=`�7=��6=Z66=�v5=�4=�3=u03=3k2=�1=��0=�0=�@/=uo.=8�-=��,=��+=}
+=k(*=�B)=�X(=k'=�x&=>�%=�$={�#=��"=�t!=�b =EJ=y*==��=�=�[=�=��=�e=�=�='=Ġ=�=�=�
=�U	=��=�=MO=O�=5� =��<\��<���<�9�<���<Y��<���<�1�<�\�<��<���<b��<T��<���<j��<��<�<��<�%�<�,�<�2�<E7�<:�<G;�<�:�<�8�<5�<�/�<�)�<("�<��<��<��<�y<��q<��i<��a<)�Y<k�Q<��I<��A<�9<ݎ1<ɋ)<v�!<J�<�<Z�	<>�<rM�;il�;���;���;��;a�;�Ŕ;�>�;��k;��L;#b.;�;���:��:��Y:hp�9�Ј������w� ������[1�]�-���H��Tc���}����� [��Qɤ�n����漻��Ȼ�ӻ�%߻�
�ӭ���������	�!\� �����{ ��$�|�(��,���0���4�2n8��<�9�?��&C��F���I�>;M�RzP�I�S���V�M�Y�{
]��`��c��f��i��l�_�n���q��t�ޠw��xz��K}����Cs���ׂ��:���������3_������ ��ہ���⍼�C������D��2e��mĔ��"������ۘ�]6������蜼�?������@��C���������I��Т�������V��?������j��9ǯ�$�������ݳ�q:������^󷼼O��,�������e���  �  ��N=�0N=�M=��L=B L=oK={�J=iJ=
YI=n�H=��G=AG=��F=X�E=G*E=�xD=��C=pC=dB=n�A=� A=MN@=p�?=��>=h3>=~==��<=�<=JX;=0�:=�9=,*9=Xn8=��7=�6=�56=v5=a�4=h�3=�/3=�j2=��1=g�0=�0=�@/=}o.=L�-=��,=/�+=�
+=�(*=&C)=yY(=�k'=�y&=�%=��$=A�#=E�"=�u!=~c =�J=�*=Y=��=�=�[=�=��=ve=`=\�={=�=#=�=(�
=�T	=׮==�N=��=�� =t�<���<��<s9�<h��<^��<4 �<^2�<�]�<ւ�<���<���<���<]��<��<^�<��<��<�&�<%.�<�3�<%8�<�:�<�;�<;�<�8�<�4�<�/�<�(�<d!�<��<��<r�<�y<��q<j�i<��a<!�Y<��Q<�I<Z�A<��9<-�1<��)<ɉ!<��<4�<ۓ	<T�<KP�;Vp�;��;��;{�;Eg�;�̔;�E�;R�k;S�L;yn.;Q;|��:�.�:��Y:ƣ�9�Q�������w�头���캶5�f�-���H��\c�ԛ}�����b`���Τ������뼻�ȻԻ�(߻i������������	��[��¤�#��x ���$���(�z�,���0�W�4��j8��<���?�9$C�ՐF���I��9M�yP�_�S�2�V�(�Y��
]�<`�� c�V!f�Ii�6l���n���q���t��w��{z��N}����qt���؂�Z;��_�������j_��2���� ������a⍼5C��֣��<��d��Ô�F!��/~��ژ��4��@����朼c>������@젼C��������I��Т������ZW��������k��Xȯ�S%��W���4߳��;��g�������Q��O����	���f���  �  �N=-0N=M=��L=c L=ioK=�J=J=�YI=N�H=��G=6BG=��F=~�E=w+E=�yD=�C=�C=�dB=I�A=QA=�N@=ۛ?=�>=�3>=~==��<=!<=�W;=x�:=D�9=6)9=Lm8=��7= �6={46=�t5=N�4=b�3=/3=�i2=	�1=��0=0=h@/=~o.=|�-=P�,=��+=�+=�)*=D)=|Z(=�l'=�z&=,�%=Ј$=P�#=\�"=�v!=Zd =�K=p+=�=3�=;�=�[=i=)�=�d=� =n�=s=ٞ=�=ш=��
=VS	=��=� =bM=��=�� =��<_��<7��<�8�<<��<���<� �<=3�<�^�<d��<e��<���<���<���<i��<�	�<��<Y �<)�<0�<�5�<�9�<�;�<�<�<�;�<�8�<�4�</�<(�< �<C�<��<Q�<��y<*�q<��i<��a<r�Y<�Q<�I<ϔA<ˎ9<��1<҈)<��!<��<}�<ݔ	<�<U�;`v�;a��;a��;��;�p�;�֔;ZP�;��k;�M;�.;�.;��:bK�:G�Y:���9Ym��[��]�w�G�������;���-�M�H�>jc���}�j����h���֤�����󼻭�Ȼ�Ի�.߻��<������I��m�	��Z�v����l��u ���$���(���,�D�0���4�4f8�J<��?� C�#�F�]�I��6M��vP�ЪS�T�V��Y�:]��`��"c��#f�Vi��l�� o��q�L�t�M�w��z�
S}����fv��Aڂ��<������n����_��W���� ��&����፼B��u������!b���������{���ט�o2��	����䜼d<�������꠼�A��!����𤼌I��ע�����X��峫�@��m��*ʯ�d'��~���q᳼/>����������S��+���p��h���  �  o�N=�/N=z�M=��L=� L=�oK=|�J=�J=�ZI=u�H=��G=�CG=@�F=
�E=-E=/{D=��C=�C=3fB=e�A=7A=�O@=^�?=j�>=�3>=�}==7�<=�<=W;=��:=1�9=�'9=�k8=!�7=u�6=�26=ws5=�4=�3=�-3=�h2=5�1=W�0=0=3@/=xo.=��-=��,=J�+=U+=�**=9E)=�[(=,n'=5|&=��%=V�$=̉#=Ń"=�w!=}e =sL=*,=S=��=]�=�[==��=d=��=8�==V�=E=�=�
=�Q	=ѫ=+�=�K=>�=|� =��<Ѓ�<��<@8�<���<���<h�<a4�<o`�<_��<���<B��<���<���<���<��<�<L#�<�+�<�2�<�7�<J;�<2=�<|=�<<�<�8�<F4�<'.�<�&�<S�<0�<��<��<��y<��q<=�i<*�a<>�Y<F�Q<��I<�A<��9<��1<X�)<!�!<�<َ<&�	<!�<([�;~�;���;���;�(�;	~�;v�;1^�;!�k;#M;`�.;�E;�H�:�o�:qZ:�P�9;H����@�w�>���U��oD��-���H��{c�ɽ}�ǋ��s��P⤻	�����=�Ȼ�Ի6߻�껂���������J�	��Y������	�pq ��$�h�(���,��0�C�4��_8�<�"�?��C�?�F�8�I��3M�ItP��S�A�V���Y��]�(`��$c��&f�R"i�!l��o�v�q�R�t�w�w�E�z��X}�����x��r܂��>������� ���`������� �����������@������\ ���_��R������x���Ԙ�T/�������᜼�9��b����蠼:@������2�+I����������Y��3�����$o���̯�*��R���|䳼:A�����������U����������i���  �  ��N=/N=#�M=��L=� L=.pK=&�J=�J=�[I=��H=~�G=0EG=�F=��E=�.E=�|D=.�C=rC=�gB=��A=CA=pP@=��?=��>=�3>=�}==��<=�<=#V;=u�:=��9=}&9=]j8=o�7=��6=816=�q5=F�4=��3=~,3=�g2=;�1=��0=�0=�?/=so.=��-=.�,=�+=J+=�+*=�F)=?](=�o'=�}&=p�%=�$=�#=T�"=;y!=�f =�M=-=�=��=z�=r[=�=�='c=n�=ِ=y=��=X=�=�
=�O	=Ω=A�=J=��=� =��<��<���<f7�<���<��</�<�5�<=b�<���<k��<M��<��<3��<.�<��<��<�&�<�.�<h5�<(:�<T=�<�>�<�>�<�<�<�8�<�3�<.-�<@%�<X�<��<��<b��<��y<��q<��i<߳a<�Y<o�Q<5�I<w�A<�9<��1<��)<S�!<�</�<��	<��<@b�;��;˵�;���;�6�;���;��;n�;0�k;bAM;��.;8a;y�:왨:eVZ:ۿ�9W��0����w�˯�����4O���-���H�q�c���}�tӋ�[���碌���v
����ȻRԻ�>߻�����7������	�fX��	�Ü����l �n�$�&�(�c�,���0��4��X8�� <���?��C���F�~�I�}/M�$qP��S�&�V���Y��]��`��'c��*f��&i��l��o��q�+�t�W�w��z��_}�����{��߂��@��Ρ�����~a�����f �����yߍ�?�����������\��,������Su��ј��+�������ޜ��6�������格f>������W祿�H�����8���Z��ж�����q��aϯ� -�������糼�D�����#����X��v������k���  �  ��N=t.N=�M=��L=� L=�pK=տJ=�J=]I=�H=�G=�FG=ǔF=��E=�0E=�~D=��C=(C=,iB=��A=fA=OQ@=��?=�>=�3>=�}==b�<=B<=4U;=H�:=y�9=�$9=�h8=��7=��6=J/6=�o5=|�4=��3=+3=�f2=/�1=��0=0=�?/=oo.=-�-=��,=��+=I+=-*=�G)=�^(=�q'=�&=L�%=�$=M�#=�"=�z!=$h =�N=�-=�=F�=��=I[=-=)�=$b=+�=R�=�=��=E=�=��
=JM	=��=1�=/H=ߎ=�� =�<��<6��<�6�<_��<L��<	�<7�</d�<���<<��<���<���<���<�<v�<i �<S*�<B2�<Y8�<�<�<v?�<m@�<�?�<#=�<�8�<-3�<	,�<�#�<)�<��<��<���<'�y<��q<��i<׫a<�Y<�Q<|�I<\�A<�9<�1<m�)<F�!<V�<z�<��	<S�<�i�;��;��;���;yE�;���;��;�~�;l;ZbM;B�.;�};F��:uǨ:��Z:6�9�у���w�C���u	�Z�1�-�-�H�G�c�s�}�����a���{����+�������Ȼf&Ի9H߻�&����������ވ	�BW�:������yg ���$�r�(�&�,�q�0�Y�4��P8�u�;�\�?��C��|F�V�I�H+M��mP�ΤS��V���Y��]� `��*c��.f��+i�r"l�bo� �q���t��w���z�$g}�Y�����ႼVC������Q��ub��e���B ��?��?ލ�`=��m���R����Y��Ʒ�����q��A͘��'��せ�ۜ��3�����!䠼|<��+���rrH��@�������\[������7��It��hү�s0��J����볼�H��ޤ��� ��=\���������)n���  �  ��N=�-N=ZM=p�L=� L=�pK=~�J=�J='^I={�H=��G=�HG=��F=��E=�2E=��D=��C=�C=�jB=I�A=|A=*R@=5�?=s�>=�3>=_}==��<=�<=;T;=�:=�9=T#9=�f8=��7=��6=b-6=n5=��4=@�3=�)3=5e2=�1=��0=g0=O?/=_o.=`�-=,�,=��+=>+=I.*=aI)=h`(=7s'=��&=*�%=ɏ$=�#=��"=T|!=�i =�O=�.=B=��=��=[=�=`�=a=��=ƍ==��=.=��=��
=K	=y�=�=<F='�=� =w�<�}�<���<�5�<���<���<��<h8�<f�<b��<��<���<��<���<�	�<U�<4$�<�-�<�5�<Z;�<[?�<�A�<B�<�@�<�=�<�8�<�2�<�*�<�!�<��<N�<[�<b��<��y<��q<��i<��a<;�Y<��Q<��I<f~A<�{9<K{1<9})<@�!<g�<��<d�	<�<q�;W��;���;�	�;T�;���;P�;��;�<l;?�M;��.;I�;���:3�:L�Z:;��9 ���}w���w�b���'�f���-�DI�8�c�(~�q�������9��]%��q�Ȼm1Ի�Q߻�.�����N!�����؈	�0V��\���
�nb ���$��(��,��0���4�6I8��;�?�?�sC��vF�N�I�?'M��jP���S��V���Y�]�]"`�$.c�3f�1i�B(l�o�Mr���t���w�X�z��n}����H����䂼�E���������vc������8 ���~��ݍ��;��P��������V����������m��eɘ�($��8~���ל��0��5����ᠼ�:��̓����)H��x��������\��R�������v��wկ��3��푲�fﳼ]L������s���_������v���p���  �  ��N="-N=�~M=K�L=!L=XqK=�J=YJ=-_I=��H=
�G=3JG=I�F=O�E=c4E=l�D=x�C=\C=lB=��A=zA=�R@=��?=��>=�3>=+}==z�<=�<=MS;=�:=��9=�!9=Fe8=	�7=)�6=�+6=@l5=�4=��3=(3= d2=�1=�0=�0=�>/=No.=��-=��,=/�+=(+=[/*=�J)=�a(=�t'=4�&=Ԍ%=s�$=��#=N�"=�}!=�j =�P=�/=�=��=��=�Z=<=��=`=��=Y�=X=��=F=�~=��
=�H	=q�=1�=kD=��=�� =�<�{�<F��<�4�<���<���<z�<�9�<�g�<���<���<���<f��<��<q�<��<�'�<61�<�8�<>�<�A�<uC�<pC�<�A�<>�<�8�<�1�<�)�<. �<��<�
�<V��<�<��y<5�q<��i<�a<��Y<��Q<!}I<�xA<�v9<Kw1<*z)<S!<~�<ޏ<��	<,�<�w�;آ�;j��;A�;�a�;'��;K$�;z��;![l;��M;|/;��;��:5�:u,[:L
�9�w��8d��w�lĴ�3)�`r���-��I���c�c~����ĩ������F���1��=�Ȼ#<Ի�Z߻b6껱���4%�����و	�)U�.�i�����] �:�$��(�v�,��0���4�HB8�#�;��?�dC�|qF���I�k#M��gP��S�)�V��Y�']�q$`�L1c�7f��5i��-l�Po��	r��t���w�w�z��u}� !��V���y炼 H������J��cd��I�) ��~��܍�0:��[���Y���T��q���4��sj���Ř�� ���z��qԜ��-�������ߠ��8�������줼�G������b ���]��������ty��hد�7��F������O��?�������b���������r���  �  )�N=�,N=�~M=&�L=.!L=�qK=��J=J=`I=ͮH=B�G=�KG=��F=��E=�5E=�D=��C=�C=DmB=��A=YA=�S@=3�?=��>=�3>=�|==�<==<=�R;=�:=��9=� 9=�c8=��7=��6=	*6=�j5=��4=_�3=�&3=�b2=1�1=k�0=_0=�>/=<o.=��-=��,=��+=�+=Q0*=�K)=c(=!v'=��&=W�%=��$=.�#=��"=�~!=�k =�Q=_0=P=;�=Ü=�Z=�=�=C_=��=�=�=]�=�=�|=��
=.G	=��=��=�B=�=f� =��<6z�<��<�3�<T��<���<�<�:�<<i�<o��<��<?��<!��<��<��<��<�*�< 4�<8;�<f@�<�C�<	E�<�D�<gB�<h>�<�8�<\1�<�(�<��<��<u�<���<H�<A�y<��q<X�i<~�a<v�Y<�~Q<�wI<�sA<�r9<�s1<�w)<�}!<��<�<��	<0�<}}�;z��;Q��;� �;m�;�Ǥ;�1�;���;Mvl;$�M;�+/;�;~6�:>�:�c[:*b�9�����S�^�w�˴�c6�c|��.�|(I���c�3~�]��d����$��}R���<���ȻWEԻ�b߻�<�����}(������	�^T�}������Y ���$�ȴ(���,��0�l}4�<8��;�+z?�F�B��lF���I�L M��eP�F�S�w�V��Y�@]�/&`��3c�l:f��9i��2l�v$o��r�3�t��w���z��{}�$�������邼J��>������3e���� ���}��8ۍ��8������R����Q��ٮ��o��mg��������w���ќ�1+��}����ݠ�x7������1줼�G������^������t���{���گ��9��I������S��T����
���e�����O���t���  �  ��N=&,N=R~M=�L=6!L=�qK=��J=�J=�`I=��H=2�G=�LG=ΚF=��E=7E=�D=��C=� C=+nB=M�A=A=T@=��?=(�>=�3>=�|==��<=�<=�Q;=-�:=��9=�9=�b8=h�7=q�6=�(6=�i5=i�4=M�3=�%3=b2=��1=��0=�
0=r>/=,o.=ʜ-=9�,=#�+=t+=1*=�L)=d(=)w'=��&=l�%=�$=7�#=��"=�!=�l =sR=�0=�=s�=Ü=�Z=v=��=�^=��=�=�=$�=B=�{=U�
=�E	=c�=/�=�A=�=o� =Y�<�x�<��<43�<��<���<��<j;�<_j�<ݒ�<���<=��<?��<O�<��<A!�<�,�<+6�<;=�<B�<6E�<5F�<�E�<�B�<�>�<�8�<�0�<�'�<��<x�<��<���<�<��y<��q<N�i<��a<��Y<�yQ<rsI<�oA<Bo9<)q1<�u)<*|!<��<�<v�	<��<���;f��;��;�(�;v�;$Ѥ;�;�;Զ�;Z�l;��M;�>/;�;�T�:eX�:5�[:)��9����I���w�\Ѵ��A���o.�5I�~�c��C~��������-���Z���E��$�ȻqLԻ<i߻�A껹���\+��Q����	��S�; �C��F��V �T�$���(���,���0��x4��78���;��u?�7�B��iF���I��M��cP��S��V�B�Y� ]��'`�6c�=f�:=i�p6l��(o�@r���t���w�c�z��}�G&��쉁��낼�K����������e��É� ��X}���ڍ�8��f������O��ά��K	��7e������o���u���Ϝ�H)��炟�dܠ�g6�������뤼�G��#�������_���������i}���ܯ��;������Q���uU���������g��º���v���  �  4�N=�+N=+~M=��L=>!L=�qK=1�J=�J=4aI=�H=��G=6MG=��F=��E=�7E=ƅD=��C=P!C=�nB=ƻA=hA=hT@=��?=B�>=�3>=�|==��<=t<=~Q;=��:=&�9=�9=b8=��7=��6=(6=�h5=��4=��3=Z%3=�a2=�1=��0=�
0=X>/=o.=ٜ-=T�,=f�+=�+=v1*= M)=�d(=�w'=g�&=$�%=��$=�#=J�"={�!=m =�R=?1=�=��=Ɯ=qZ=K=6�=.^=@�=�=)=`�=�
=�z=l�
=�D	=��=o�=�@=\�=�� =X�<x�<{��<�2�<���<���<��<�;�<k�<���<���<n��<���<��<Q�<�"�<_.�<�7�<p>�<4C�<F�<G�<F�<:C�<�>�<r8�<�0�<M'�<��<�<��<���<��<��y<��q<��i<$�a<��Y<wQ<�pI<�mA<"m9<�o1<Et)<q{!<��<�<�	<��<���;ٳ�;X��;�-�;�{�;=פ;�A�;���;8�l;Y�M;�I/;~�;�f�:5h�:��[:���9V�$E���w�մ�LI�����.��<I���c�cM~�-��3Ę��3�� a��~J��5�Ȼ�PԻ'm߻9E�:���1-������	��S���� �����U ��$�V�(��,�Р0��u4��48���;�s?���B�TgF��I�KM��bP���S���V�j�Y�]��(`�`7c��>f�P?i��8l�S+o��r���t���w���z��}��'��9����삼�L��X���"	��Qf��EÉ�) ��'}��5ڍ�f7���������N����������c��"������_t��_Μ� (��ف���۠��5��<����뤼uG��D������X`��[������v~��ޯ�D=��雲�����W��@�����*i��Dú����v���  �  �N=�+N=~M=��L=F!L=	rK=G�J=J=RaI=L�H=��G=kMG=��F=��E=8E=��D=��C=�!C=�nB=��A=�A=�T@=ϟ?=V�>=�3>=�|==z�<=X<=bQ;=�:=��9=�9=�a8=^�7=q�6=�'6=�h5=��4=b�3="%3=`a2=�1=k�0=�
0=H>/=o.=�-=i�,=��+=�+=�1*=]M)=�d(=x'=��&=Z�%=��$=�#=y�"=��!=Zm =�R=\1==��=ל=bZ=6=�=	^=�=J�=�=�=@
=gz=@�
=�D	=/�=/�=�@="�=�� =�<�w�<G��<�2�<ҁ�<��<��</<�<Tk�<��<"��<���<��<&�<��<$#�<�.�<�7�<�>�<�C�<TF�<@G�<9F�<aC�<�>�<X8�<}0�<'�<��<#�<5�<��<�<��y<x�q<t�i<2�a<�Y<vQ<�oI<�lA<nl9<o1<�s)<+{!<r�<B�<?�	<�<���;��;&��;�/�;�}�;+٤;�C�;���;Úl;8�M;�M/;��;$m�:�l�:��[:��9��~�;D�ދw�s״�rL�j��H.��?I�� d� Q~�w���Ř��4��8c��YL��7�Ȼ�RԻ�n߻sF�&���.��ݟ�>�	�BS�a����� ���T ��$���(��,��0�u4��38��;�Mr?��B�ZfF�|�I��M�MbP�;�S�i�V���Y��]�)`��7c�c?f�
@i��9l�Z,o��r���t���w�L�z�B�}�(������)킼M������[	��}f��^É�1 ���|��ڍ�)7��\�����eN��.���y��bc����������s���͜��'��k���V۠�j5�����Y뤼ZG��Z��� ���`������+���~��xޯ��=��l���s���BW���������i���ú���Sw���  �  4�N=�+N=+~M=��L=>!L=�qK=1�J=�J=4aI=�H=��G=6MG=��F=��E=�7E=ƅD=��C=P!C=�nB=ƻA=hA=hT@=��?=B�>=�3>=�|==��<=t<=~Q;=��:=&�9=�9=b8=��7=��6=(6=�h5=��4=��3=Z%3=�a2=�1=��0=�
0=X>/=o.=ٜ-=T�,=f�+=�+=v1*= M)=�d(=�w'=g�&=$�%=��$=�#=J�"={�!= m =�R=@1=�=��=Ȝ=rZ=M=8�=0^=C�=��=-=d�=�
=�z=r�
=�D	=��=w�=�@=f�=�� =l�<,x�<���<�2�<��<��<��<<�<'k�<œ�<���<w��<���<��<R�<�"�<Z.�<�7�<g>�<(C�<F�<�F�<�E�<)C�<�>�<a8�<�0�<='�<��<q�<��<���<��<��y<|�q<��i<)�a<��Y<wQ<�pI<�mA<>m9<�o1<ft)<�{!<<;�<�	<��<���;��;���;�-�;�{�;Oפ;�A�;���;�l;$�M;�I/;�;�e�:/g�::�[:���9{H��G�^�w�~ִ��J�v��:.�d=I���c��M~�u��uĘ��3��7a���J��a�Ȼ�PԻJm߻WE�T���H-�����#�	��S����$�����U ��$�X�(��,�Ҡ0��u4��48���;�s?���B�TgF��I�LM��bP���S���V�j�Y�]��(`�`7c��>f�P?i��8l�S+o��r���t���w���z��}��'��9����삼�L��X���"	��Qf��EÉ�) ��'}��5ڍ�f7���������N����������c��"������_t��_Μ� (��ف���۠��5��<����뤼uG��D������X`��[������v~��ޯ�D=��雲�����W��@�����*i��Dú����v���  �  ��N=&,N=R~M=�L=6!L=�qK=��J=�J=�`I=��H=2�G=�LG=ΚF=��E=7E=�D=��C=� C=+nB=M�A=A=T@=��?=(�>=�3>=�|==��<=�<=�Q;=-�:=��9=�9=�b8=h�7=q�6=�(6=�i5=i�4=M�3=�%3=b2=��1=��0=�
0=r>/=,o.=ʜ-=9�,=#�+=t+=1*=�L)=d(=)w'=��&=l�%=�$=7�#=��"=�!=�l =tR=�0=�=u�=Ŝ=�Z=y=��=�^=��=$�=�=-�=L=�{=a�
=�E	=r�=@�=�A=�=�� =��<y�<6��<\3�<9��<	��<��<�;�<}j�<���<���<N��<K��<V�<��<>!�<�,�<6�<)=�<B�<E�<F�<nE�<�B�<t>�<j8�<�0�<�'�<v�<]�<��<���<��<{�y<�q<N�i<��a<��Y<zQ<�sI<	pA<wo9<dq1<�u)<l|!<A�<J�<��	<��<5��;ϰ�;_��;)�;Jv�;GѤ;�;�;̶�;�l;D�M;>/;N�;�R�:lV�:χ[:���9���+O�.�w�!Դ�hD����.�V6I���c��D~�������.��6[���E��z�Ȼ�LԻi߻B������+��c���	��S�F �L��N��V �Y�$�İ(���,���0��x4��78���;��u?�8�B��iF���I��M��cP��S��V�B�Y� ]��'`�6c�=f�:=i�q6l��(o�@r���t���w�c�z��}�G&��쉁��낼�K����������e��É� ��X}���ڍ�8��f������O��ά��K	��7e������o���u���Ϝ�H)��炟�dܠ�g6�������뤼�G��#�������_���������i}���ܯ��;������Q���uU���������g��º���v���  �  )�N=�,N=�~M=&�L=.!L=�qK=��J=J=`I=ͮH=B�G=�KG=��F=��E=�5E=�D=��C=�C=DmB=��A=YA=�S@=3�?=��>=�3>=�|==�<==<=�R;=�:=��9=� 9=�c8=��7=��6=	*6=�j5=��4=_�3=�&3=�b2=1�1=k�0=_0=�>/=<o.=��-=��,=��+=�+=Q0*=�K)=c(=!v'=��&=X�%=��$=.�#=��"=�~!=�k =�Q=a0=R=>�=Ɯ=�Z=�=�=I_=��=#�=�=i�=�=�|=��
=AG	=��=��=C=-�=�� =/�<oz�<H��<4�<���<	��<K�<�:�<fi�<���<��<W��<3��<"��<��<��<�*�<�3�<;�<H@�<�C�<�D�<wD�<9B�<9>�<�8�<.1�<~(�<��<��<U�<���<3�<$�y<��q<X�i<��a<��Y<�~Q<�wI<�sA<�r9<)t1<�w)<�}!<�<e�<�	<��<"~�;��;���;!�;am�;�Ǥ;�1�;�;�ul;��M;�*/;�;4�:J;�:_][:�T�9�ˀ�E[��w��δ�M:�Q~��.�L*I���c��4~�!�����]%��S��s=����Ȼ�EԻ@c߻ =�����(�������	�qT��������Y ���$�δ(��,��0�p}4�
<8��;�-z?�G�B��lF���I�M M��eP�G�S�w�V��Y�@]�/&`��3c�l:f��9i��2l�w$o��r�3�t��w���z��{}�$�������邼J��>������3e���� ���}��8ۍ��8������R����Q��ٮ��o��mg��������w���ќ�1+��}����ݠ�x7������1줼�G������^������t���{���گ��9��I������S��T����
���e�����O���t���  �  ��N="-N=�~M=K�L=!L=XqK=�J=YJ=-_I=��H=
�G=3JG=I�F=O�E=c4E=l�D=x�C=\C=lB=��A=zA=�R@=��?=��>=�3>=+}==z�<=�<=MS;=�:=��9=�!9=Fe8=	�7=)�6=�+6=@l5=�4=��3=(3= d2=�1=�0=�0=�>/=No.=��-=��,=/�+=(+=[/*=�J)=�a(=�t'=4�&=Ԍ%=s�$=��#=O�"=�}!=�j =�P=�/=�=��=��=�Z=A=��=$`=��=e�=e=�=W=�~=��
=I	=��=M�=�D=��=�� =I�<!|�<���<�4�<���<���<��<�9�<�g�<���<۱�<���<{��<��<t�<��<�'�<1�<|8�<�=�<uA�<DC�<;C�<gA�<�=�<�8�<�1�<t)�<��<��<�
�<5��<��<h�y<#�q<��i<%�a<�Y<ׄQ<c}I<yA<w9<�w1<�z)<�!<�<T�<�	<��<�x�;���;��;��;b�;c��;c$�;m��;�Zl;�M;�/;��;��:��:�$[:���9J���mm�_�w�8ɴ��-�t���-��I�	�c�d ~� �����������G��[2����Ȼ�<ԻL[߻�6�	����%�������	�@U�B�y�����] �C�$���(�}�,��0���4�LB8�&�;��?�fC�}qF���I�l#M��gP��S�*�V��Y�(]�q$`�L1c�7f��5i��-l�Po��	r��t���w�w�z��u}� !��V���y炼 H������J��cd��I�) ��~��܍�0:��[���Y���T��q���4��sj���Ř�� ���z��qԜ��-�������ߠ��8�������줼�G������b ���]��������ty��hد�7��F������O��?�������b���������r���  �  ��N=�-N=ZM=p�L=� L=�pK=~�J=�J='^I={�H=��G=�HG=��F=��E=�2E=��D=��C=�C=�jB=I�A=|A=*R@=5�?=s�>=�3>=_}==��<=�<=;T;=�:=�9=T#9=�f8=��7=��6=b-6=n5=��4=@�3=�)3=5e2=�1=��0=g0=O?/=_o.=`�-=,�,=��+=>+=I.*=aI)=h`(=8s'=��&=+�%=ɏ$=�#=��"=U|!=�i =�O=�.=E=��=��=[=�=h�=&a=��=ҍ==ė=A=Ҁ=��
=+K	=��=8�=^F=K�=1� =��<&~�<���<�5�<B��<���<�<�8�<Af�<���<9��<���<7��<���<�	�<O�<$$�<�-�<c5�<1;�<*?�<OA�<�A�<v@�<Y=�<�8�<S2�<�*�<�!�<��<!�<6�<E��<g�y<��q<��i<ˣa<a�Y<ËQ<�I<�~A<�{9<�{1<�})<��!<�<%�<�	<[�<�q�;!��;d��;{
�;~T�;Ѭ�;l�;�;<l;{�M;��.;�;n��:c�:��Z:���9����Á�;�w��´��Pi�N�-��I���c�d	~�|w������[:��&���Ȼ 2ԻbR߻A/�(����!�������	�JV��n���
�zb ���$��(��,�
�0���4�9I8��;�A�?�uC��vF�O�I�@'M��jP���S��V���Y�]�]"`�$.c�3f�1i�B(l�o�Mr���t���w�X�z��n}����H����䂼�E���������vc������8 ���~��ݍ��;��P��������V����������m��eɘ�($��8~���ל��0��5����ᠼ�:��̓����)H��x��������\��R�������v��wկ��3��푲�fﳼ]L������s���_������v���p���  �  ��N=t.N=�M=��L=� L=�pK=տJ=�J=]I=�H=�G=�FG=ǔF=��E=�0E=�~D=��C=(C=,iB=��A=fA=OQ@=��?=�>=�3>=�}==b�<=B<=4U;=H�:=y�9=�$9=�h8=��7=��6=J/6=�o5={�4=��3=+3=�f2=/�1=��0=0=�?/=oo.=,�-=��,=��+=I+=-*=�G)=�^(=�q'=�&=M�%=�$=N�#=�"=�z!=&h =�N=�-=�=J�=��=N[=4=1�=-b=6�=_�=�=��=Y= �=��
=eM	=ħ=R�=RH=�=�� =[�<6��<���<�6�<���<���<Q�<T7�<jd�<1��<g��<���<���<��<�<o�<Y �<9*�<2�<.8�<�<�<>?�<0@�<b?�<�<�<�8�<�2�<�+�<W#�<��<��<Z�<���<��y<��q<��i<�a<F�Y<N�Q<ȊI<��A<K�9<�1<�)<˃!<ވ<�<y�	<ѥ<�j�;���;���;v��;�E�;;��;�~�;�l;�aM;"�.;m|;ר�:�è:ΗZ:�"�9#��d���w�ͻ����T]���-���H���c���}��ዻa���e���U,�����j�Ȼ�&Ի�H߻5'�3���p�������	�]W�Q�������g ���$�{�(�.�,�w�0�]�4��P8�x�;�^�?��C��|F�W�I�I+M��mP�ϤS��V���Y��]� `��*c��.f��+i�r"l�bo�!�q���t��w���z�$g}�Y�����ႼVC������Q��ub��e���B ��?��?ލ�`=��m���R����Y��Ʒ�����q��A͘��'��せ�ۜ��3�����!䠼|<��+���rrH��@�������\[������7��It��hү�s0��J����볼�H��ޤ��� ��=\���������)n���  �  ��N=/N=#�M=��L=� L=.pK=&�J=�J=�[I=��H=~�G=0EG=�F=��E=�.E=�|D=.�C=rC=�gB=��A=CA=pP@=��?=��>=�3>=�}==��<=�<=#V;=u�:=��9=}&9=]j8=o�7=��6=816=�q5=F�4=��3=~,3=�g2=;�1=��0=�0=�?/=so.=��-=.�,=�+=J+=�+*=�F)=?](=�o'=�}&=p�%=�$=��#=T�"=<y!=�f =�M=-=�=��=~�=w[=�=�=0c=y�=�=�=��=k=#�= �
=�O	=�=`�=4J==D� =��<:��<��<�7�<���<^��<t�<�5�<vb�<ʈ�<���<n��<��<A��<1�<��<��<�&�<�.�<>5�<�9�<=�<�>�<L>�<[<�<�8�<�3�<�,�<%�<%�<��<t�<F��<��y<��q<��i<�a<'�Y<��Q<�I<ЊA<i�9< �1<�)<Ӆ!<��<��<	�	<)�<"c�;߇�;y��;��;�6�;���;8��;n�;��k;�@M;��.;�_;�u�:��:�MZ:`��9�a��v��F�w�$�������Q�O�-�6�H�ϒc���}�ԋ�S���𤻏��0��E�Ȼ�Ի%?߻��[������ٚ�8�	�X��	�՜�	��l �x�$�.�(�j�,� �0��4��X8�<���?��C���F��I�~/M�%qP��S�'�V���Y��]��`��'c��*f��&i��l��o��q�+�t�W�w��z��_}�����{��߂��@��Ρ�����~a�����f �����yߍ�?�����������\��,������Su��ј��+�������ޜ��6�������格f>������W祿�H�����8���Z��ж�����q��aϯ� -�������糼�D�����#����X��v������k���  �  o�N=�/N=z�M=��L=� L=�oK=|�J=�J=�ZI=u�H=��G=�CG=@�F=
�E=-E=/{D=��C=�C=3fB=e�A=7A=�O@=^�?=j�>=�3>=�}==7�<=�<=W;=��:=1�9=�'9=�k8=!�7=u�6=�26=ws5=�4=�3=�-3=�h2=5�1=W�0=0=3@/=xo.=��-=��,=J�+=U+=�**=9E)=�[(=,n'=5|&=��%=V�$=̉#=Ń"=�w!=e =uL=,,=V=��=`�=�[==��=#d=��=D�=&=e�=V="�="�
=�Q	=�=H�=�K=^�=�� =;�<��<M��<�8�<B��<��<��<�4�<�`�<���<ئ�<`��<���<���<���<��<�<5#�<�+�<p2�<�7�<;�<�<�<E=�<�;�<�8�<4�<�-�<�&�<%�<�<c�<��<��y<��q<=�i<<�a<a�Y<y�Q<їI<h�A<�9<�1<Ɔ)<��!<b�<N�<��	<��<�[�;�~�;���;]��;;)�;E~�;��;$^�;��k;R"M;g�.;�D;�E�:@l�:�Z::@�9����K����w�	��� ���F�g�-��H��}c�ʿ}�
ȋ��t��㤻�������ҩȻ�Ի�6߻b�ڷ��=�� ��e�	��Y������|q ��$�o�(���,��0�G�4��_8�<�$�?��C�@�F�9�I��3M�JtP��S�A�V���Y��]�(`��$c��&f�R"i�!l��o�v�q�R�t�w�w�E�z��X}�����x��r܂��>������� ���`������� �����������@������\ ���_��R������x���Ԙ�T/�������᜼�9��b����蠼:@������2�+I����������Y��3�����$o���̯�*��R���|䳼:A�����������U����������i���  �  �N=-0N=M=��L=c L=ioK=�J=J=�YI=N�H=��G=6BG=��F=~�E=w+E=�yD=�C=�C=�dB=I�A=QA=�N@=ۛ?=�>=�3>=~==��<=!<=�W;=x�:=D�9=6)9=Lm8=��7= �6={46=�t5=N�4=b�3=/3=�i2=	�1=��0=0=h@/=~o.=|�-=P�,=��+=�+=�)*=D)=|Z(=�l'=�z&=,�%=Ј$=P�#=\�"=�v!=[d =�K=q+=�=6�=>�=�[=n=.�=�d=� =x�=}=�=�=�=��
=jS	=��=� ={M=��=�� =&�<���<p��<09�<t��<���<� �<l3�<_�<���<���<ѿ�<���<���<l��<�	�<��<F �<�(�<�/�<y5�<`9�<�;�<[<�<Q;�<�8�<{4�<�.�<�'�<��<"�<��<<�<��y<�q<��i<��a<��Y<6�Q<�I<�A<�9<�1<,�)<�!<��<ݎ<;�	<[�<�U�;�v�;��;���;F�;q�;ה;OP�;<�k;9M;��.;�-;F�:�H�:�Y:'��9������w�1�������=���-��H��kc�J�}�.���9i���פ�k��o���&�Ȼ�Ի�.߻J껃���5��d����	��Z������w��u ��$���(���,�H�0���4�7f8�L<��?� C�$�F�^�I��6M��vP�ЪS�T�V��Y�:]��`��"c��#f�Vi��l�� o��q�L�t�M�w��z�
S}����fv��Aڂ��<������n����_��W���� ��&����፼B��u������!b���������{���ט�o2��	����䜼d<�������꠼�A��!����𤼌I��ע�����X��峫�@��m��*ʯ�d'��~���q᳼/>����������S��+���p��h���  �  ��N=�0N=�M=��L=B L=oK={�J=iJ=
YI=n�H=��G=AG=��F=X�E=G*E=�xD=��C=pC=dB=n�A=� A=MN@=p�?=��>=h3>=~==��<=�<=JX;=0�:=�9=,*9=Xn8=��7=�6=�56=v5=a�4=h�3=�/3=�j2=��1=g�0=�0=�@/=}o.=L�-=��,=/�+=�
+=�(*=&C)=yY(=�k'=�y&=�%=��$=A�#=F�"=�u!=c =�J=�*=Z=��=!�=�[=�=��={e=e=c�=�=�=-=#�=5�
=�T	=�==�N=��=�� =��<���<G��<�9�<���<���<X �<2�<�]�<���<���<���<���<d��<��<Z�<��<��<�&�<.�<�3�<	8�<�:�<�;�<�:�<�8�<�4�<�/�<�(�<I!�<��<��<c�<�y<��q<j�i<��a<4�Y<��Q</�I<��A<3�9<h�1<��)<�!<A�<x�<�	<��<�P�;�p�;x��;]��;��;hg�;�̔;�E�;�k;��L;�m.;�;���:�,�:��Y:4��9Cz����r�w��������7���-��H�^c���}�C����`��VϤ�!���X켻m�ȻfԻ8)߻��5����������	��[��ˤ�+��x ���$���(�}�,���0�Y�4��j8��<���?�:$C�֐F���I��9M�yP�_�S�2�V�(�Y��
]�<`�� c�V!f�Ii�6l���n���q���t��w��{z��N}����qt���؂�Z;��_�������j_��2���� ������a⍼5C��֣��<��d��Ô�F!��/~��ژ��4��@����朼c>������@젼C��������I��Т������ZW��������k��Xȯ�S%��W���4߳��;��g�������Q��O����	���f���  �  ��N=�0N=�M=��L=0 L=�nK=/�J=J=�XI=�H=%�G=q@G=�F=��E=})E=�wD=4�C=�C=icB=�A=$ A=�M@=*�?=��>=X3>=~==��<=�<=�X;=��:=��9=�*9=o8=`�7=��6=Z66=�v5=�4=�3=u03=3k2=�1=��0=�0=�@/=uo.=8�-=��,=��+=}
+=k(*=�B)=�X(=k'=�x&=>�%=�$={�#=��"=�t!=�b =FJ=y*==��=�=�[=�=��=�e=�=�=*=ɠ=�=��=�
=�U	=��=�=VO=X�=?� =��<q��<���<�9�<���<m��<���<�1�<]�<���<���<k��<[��<���<k��<��<�<��<�%�<�,�<�2�<67�<�9�<6;�<�:�<�8�<�4�<�/�<�)�<"�<��<��<��<��y<��q<��i<��a<3�Y<z�Q<��I<��A<��9<��1<�)<��!<m�<?�<|�	<_�<�M�;�l�;��;���;��;)a�;�Ŕ;�>�;��k;��L;�a.;};���:��:i�Y:uk�9戸n����w�����J��2��-�P�H��Uc�&�}�����b[���ɤ������漻ӓȻ)�ӻ�%߻�
�����������	�(\��#����{ ��$�~�(��,���0���4�3n8��<�:�?��&C��F���I�>;M�RzP�I�S���V�N�Y�{
]��`��c��f��i��l�_�n���q��t�ޠw��xz��K}����Cs���ׂ��:���������3_������ ��ہ���⍼�C������E��2e��mĔ��"������ۘ�]6������蜼�?������@��C���������I��Т�������V��?������j��9ǯ�$�������ݳ�q:������^󷼼O��,�������e���  �  `�N=9N=@�M=��L=�*L=zK=��J=�J=�dI=��H=P H=@NG={�F=#�E=d:E=�D=5�C=�*C=p{B=;�A=�A=�l@=��?=~?=vY>=��==��<=�=<=��;=��:=:=e`9=�8=��7=27=Nv6=��5=�4==4=�|3=�2=Z�1=�11=Ni0=��/=��.=��-=�+-=`T,=Uy+=��*=>�)=��(=��'=S�&=�&=Q%=�$=I#=�	"=�� =�=��=�=�z=qE=1=��=�n=�=��=�A=��=J=r�=�/=ԕ=��	=�J=��=�=�#=)_=1)�<}��<���<�&�<-g�<h��<��<+��<7�<Z.�<C�<hS�<4`�<�i�<�q�<w�<D{�<O~�<��<��<���<�~�<�{�<Cw�<�p�<�h�<?_�<�S�<LG�<U9�<�*�<�<4�<��y<Y�q<	�i<�a<��Y<�fQ<^OI<�9A<�%9<�1<D)<B� <��<D�<��<-� <A��;
�;���;��;峱;��;$�;�z�;��e;`�F;t(;7�	;oP�:��:�e<:�?�9��@�!%�Kb����ź�m���>�!�6��:R��!m�̃� ͐�������@V���S»�λٻK��g�ﻁ5���I�vW��D���-�� N����m#� G'�i`+�0]/�N?3��7��:��K>���A��7E� �H���K��O��<R��\U��rX�!�[�d�^��a�|d��mg�*Zj�`@m�}!p���r���u��x�lp{�:8~�9~���ށ��=����������V��	���,���m���ˌ�b*�����萼�F��Ӥ��:��f^��j�������j����������i���������b������	���^��㴧���Ud��x������8r��Dͯ��(�������޳��9��s����9I���������$Y���  �  2�N=�8N=2�M=��L=�*L=zK=��J=,J=eI=زH=� H=�NG=ϜF=x�E=�:E=Y�D=��C=+C=�{B=r�A=�A=.m@=��?=�?=�Y>=�==|�<=y=<=y�;=��:=�:=+`9=Ȧ8=��7=�17=v6=^�5=��4=�<4=�|3=ֺ2=,�1=c11=<i0=n�/=��.= .=�+-=�T,=�y+=�*={�)=:�(=�'=��&=�&=�%=A$=�#=�	"=� =L�=%�=�=�z=|E=.=��=cn=�=[�=�A=p�=3J=�=f/={�=��	=J=a�=��=x#=�^=�(�<��<���<�&�< g�<s��<<��<o��<��<�.�<�C�<�S�<�`�<�j�<r�<�w�<�{�<�~�<���<���<��<p�<=|�<�w�<q�<�h�<-_�<�S�<�F�<9�<*�<��<�
�<x�y<$�q<Ƿi<��a<6Y<�eQ<:NI<�8A<�$9<1<�)<�� <a�<G�<��<�� <̄�;��;o��;]��;b��;��;�&�;A}�;��e;�F;N(;��	;tY�:n�:`v<:�\�9��@���$��a��еź#o���@���6�>R�?$m��̓�Gϐ�풝����WX���U»nλ�ٻ��仡�ﻏ6��2J��W��D�A����EM�����#�F'�%_+�\/��=3�t7�̳:�SJ>���A�@6E��H�#�K�O��;R�N\U��rX��[�Ʌ^�h�a��|d��ng��Zj�Am�p"p���r�&�u�)�x��q{��9~��~�� ߁�>�����]���IV��2���O���m���ˌ�*�������琼)F��I�������]���������i��D���S��Zi������|��cb��Ƶ���	���^��촧�)��{d��ҽ������r���ͯ�)��a���}߳�\:�����|﷼�I���������~Y���  �  ��N=�8N=�M=��L=�*L=[zK==�J=�J=�eI=��H=wH=wOG=ɝF=��E=�;E=h�D=w�C=�+C=�|B=%�A=�A=�m@=�?=�?=�Y>=v�==Q�<=*=<=�;=�:=:=f_9=�8=��7=�07=u6=k�5=��4=<4=�{3==�2=��1=11=i0=P�/=��.=- .=D,-=�T,=z+=��*==�)=!�(=��'=��&=�&=�%=F$=n#=�
"=�� =��=��=p�=�z=�E=*=S�=n=-=��=�@=��=?I=�=G.=L�=n�	=�H=Q�=��=�"=0^=d'�<��<���<O&�<g�<���<���<��<��<�/�<E�<�U�<�b�<�l�<!t�<�y�<
~�<܀�<���<"��<���<���<&}�<+x�<q�<(i�<_�<fS�<8F�<8�<�(�<�<��<��y<"�q<s�i<��a<{Y<�aQ<�JI<�5A<�"9<�1<O)<�� <�<��<��<� <i��;��;Z��;���;-��;��;/0�;@��;��e;y�F;Q)(;v�	;�t�:�)�:��<:3��9O3@���$��]��s�ź^t��
F�d�6��GR��.m�ԃ�֐������R_���\»_λ��ٻ��#��=9���J�X�(D���n���K�����#��B'�k[+�[X/��93�97���:�F>���A��2E��H�s�K��O�E:R�[U��qX��[�,�^�*�a�~d��pg�@]j�{Dm��%p��s���u�3�x�zu{�_=~����������?��)���K����V������j���m��Pˌ�m)��݇��_搼�D�����������[���������g��F���}���g�����2��ka�����P	���^��ߴ��q���d����������s��Mϯ��*��?���e᳼g<������_�wK�����������Z���  �  �N=58N=ĉM=��L=+L=�zK=��J=wJ=�fI=´H=�H=�PG=K�F=�E=N=E=�D=��C=V-C=�}B=L�A=�A=dn@=��?=!?=�Y>=`�==��<=�<<=M�;=�:=�:= ^9=��8=C�7=?/7=}s6=��5=d�4=�:4=�z3=6�2=��1=e01=�h0="�/=��.=h .=�,-=�U,=�z+=��*=r�)=t�(=h�'=(�&=�	&=)%=�$=�#=$"=�� =��=q�=
�=J{=�E=
=�=~m=f=��=�?=5�=�G=_�=�,=��=��	=EG=��=5�=5!=�\=d%�<���<���<�%�<�f�<؞�<���<N��<>�<2�<uG�<mX�<�e�<�o�<jw�<}�<*��<���<u��<���<τ�<u��<�~�<Dy�<r�<Ai�<�^�<�R�<E�<R6�<�&�<��<0�<��y<��q<�i<�a<�tY<\Q<ZEI<�0A<[9<�1<��(<\� <{�<��<3�<|� <��;!��;;��;���;�ʱ;���;�=�;���;Of; 
G;VC(;��	;x��:�P�:e�<:��97�?���$�Y���źr~��QN��7��UR��@m��݃�^���&���F)��j��g»-λ�ٻ���<�ﻉ=��WL��X��C�b�@���H�ӷ�Y	#��='��U+�>R/��33���6� �:��?>���A�-E���H��K�F
O�i7R��XU��pX��[���^�҆a�`�d��sg�Iaj��Hm��*p�+s���u�J�x��{{�C~�X���Cぼ�A���������X��G������lm���ʌ�D(��X���{䐼�B��$��������X����������d��C�������d������#���_������j��1^��񴧼����e��񿫼���v���ѯ�q-�����]䳼o?������/���+N�������U\���  �  :�N=�7N=q�M=��L=F+L=B{K=��J=�J=�gI=F�H=uH=�RG=V�F=*�E=l?E=�D=�C=2/C=|B=��A=�A=bo@=T�?=�?=�Y>=>�==��<=�;<=^�;=��:=�:=v\9=��8=M�7=>-7=�q6=�5=��4=�84=7y3=�2=��1=�/1=h0=�/=��.=� .=N--=tV,=|+=�*=�)=*�(=V�'=(�&=�&=7%=�$=�#=�"=~� =2�={�=˨=�{=�E=�=��=�l=d=p�=>=f�=�E=/�==*=/�=K�	=�D=v�=-�=k=Y[=�"�<y��<:��<�$�<~f�<0��<Z��<���<X�<�4�<�J�<�[�<�i�<�s�<�{�<a��<e��<���<��<��<���<ㄭ<x��<�z�<�r�<]i�<B^�<Q�<iC�<4�<�#�<V�<��<��y<Z�q<��i<v�a<�lY<)TQ<.>I<�*A<�9<�	1<��(<�� <��<W�<��<B� <B��;y��;ע�;ݷ�;�ڱ;��;�O�;O��;$'f;�.G;�e(;��	;��:끚:�1=:͇�9��>���$�*T��#�ź����TY��7�9iR��Wm�냻�볝��7��3y��7u»H+λ��ٻv��	��+C��:N�&Y��C���ʸ�E����#�j7'��N+�EJ/�V+3�G�6���:��7>���A��%E�u�H�z�K��O��3R��VU�WoX�l[���^��a�l�d��wg��fj��Nm��1p��s���u�<�x���{��J~�����恼�D����������rY��(������7m���Ɍ� '��m���␼�?��՜��S����T��o�������`��-�������a�������	���]��(���j���]�������g����������x���ԯ�1��ጲ�j購dC����������Q��B�������^���  �  �N=�6N= �M=��L=�+L=�{K={�J=�J=siI=�H=xH=�TG=��F=��E=�AE=c�D=A�C=N1C=q�B=s�A=0!A=p@=�?=?=
Z>=�==�<=;<=1�;=i�:=�:=�Z9=��8=
�7=�*7=$o6=��5=U�4=�64=]w3=U�2=}�1=�.1=^g0=��/=��.=.=�--=lW,=Q}+=n�*=׽)=3�(=x�'=w '=�&=�%=$=�#=�"=C!=��=��=��=7|=F=�=�=�k=#=�=3<=:�=OC=��=�'=s�=��	=FB=��=��=@=�Y=��<��<��<�#�<5f�<���<c��<���<��<�7�<@N�<
`�<�m�<�x�<���<H��<2��<{��<b��<挵<䊱<���<���<�{�<�s�<si�<�]�<P�<UA�<q1�<� �<}�<E��<��y<��q<��i<|}a< cY<#KQ<�5I<#A<�9<c1<��(< � <��<��<��<�� <���;q��;w��;���;�;| �;�d�;v��;�Qf;�WG;��(;��	;H�:��:�=:+�9r>�F�$��O��A�ź�����g�h%7�3�R�Ysm�'���9���,ŝ��I��p���n�»W:λX�ٻ���j��vJ��}P�-Z�5C�"����@����t�"��/'�kF+�tA/��!3���6���:�6.>��A��E��xH�%�K�R O��/R��SU��mX�*[���^�K�a�O�d��|g��lj�MVm��9p�=s���u���x��{�T~�<����ꁼ/H������ ��D[��8���d���l���Ȍ��%��C���Sߐ�V<������ ���iP����������[������h��u]��
������![��W���?��]��)���T���h���ë����|���د�5��M����H�����������U�������ga���  �  ��N=�5N=��M=k�L=�+L=^|K=g�J=�J=kI=عH=�H=BWG=�F=�E=_DE=�D=��C=�3C=x�B=8�A=�"A=�q@=��?=�?=$Z>=ϥ==��<=/:<=�;=��:=�:=nX9=E�8=��7=\(7=�l6=&�5=��4=�44=gu3=��2=�1=�-1=�f0=&�/=��.=W.=�.-=jX,=�~+=�*=��)=X�(=��'=�'=i&=%=q$=2#=�"=!=5�=��=��=�|=/F=|=t�=�j=�=1�=+:=��=�@=�=�$=t�=��	=d?=,�=J�=�=~W=Q�<R~�<���<{"�<�e�<���<���<o��<K�<�:�<R�<dd�<�r�<�}�<���<���<N��<Y��<���<ݐ�<d��<j��<ń�<p}�<Kt�<li�<�\�<�N�<&?�<�.�<�<a�<���<a�y<�q<��i<�ra<�XY<3AQ<�,I<
A<�9<��0<��(<z� <��<9�<��<"� <~��;O��;���;���;� �;�5�;@{�;!ӂ;Of;��G;z�(;�
;�_�:���: �=:B��9�0=�#y$��L��S�ź����w�d:7��R��m���:��؝��\������w�»�Jλ�ٻ���ѹ�R���R�h[�C��
����<�6����"�('��=+��7/��3�E�6���:�$>�K�A��E�&qH�J�K���N��+R��PU�llX�6[�&�^��a�e�d�t�g�Rsj�^m�uBp�� s���u���x�)�{��]~�������K��ɧ�����&]��r�������l��Ȍ��#�����oܐ��8�������𔼕K�����������V���������7Y��Z���b���X��p���	���\��i���@��3j��ƫ��"������ܯ��9��'����MM������]��tZ��������md���  �  ��N=5N=��M=A�L=�+L=�|K=>�J=J=�lI=��H=�
H=�YG=��F=��E=�FE=o�D=�C=�5C=x�B=��A="$A=�r@=��?=�?=?Z>=��==��<=89<=��;=5�:=:=LV9=�8=�7=�%7=�i6=��5=��4=�24=os3=ݲ2=��1=l,1=�e0=��/=��.=�.==/-=\Y,=�+=��*=��)=p�(=�'=S'=�&=�%=�$=|#=�"=�!=��=�=Y�==}=PF=@=ؼ=�i=u=~�=8=��=->=�=�!=}�=��	=|<=h�=��=�=pU=��<�{�<���<M!�<Ee�<*��<���<-��<� �<>�<�U�<�h�<xw�<���<���<���<]��<4��<G��<Ԕ�<͑�<(��<φ�<�~�<�t�<ci�<\�<M�<�<�<�+�<��<-�<��<5�y<H�q<��i<�ga<�MY<17Q<�#I<�A<�9<Y�0<��(<�� <c�<��<��<a� <��;��;���;��;��;�J�;`��;�;�f;��G;��(;�?
;���:F0�:�P>:�G�9}c<�S\$��I��N�ź����߆�&P7���R���m���t#��띻�o�������»�[λ��ٻ���V��Z���U��\��B�)	���{8�â���"�U '��4+�>./��3���6�8�:�">���A�E�riH���K�b�N�y'R�/NU�kX�4[���^��a���d���g�+zj��em�PKp�Y*s��v�1�x�a�{��g~�����󁼶O�����O��#_��ɸ������l��Bǌ�d"���}���ِ�]5�����2씼�F�����������Q���������U������B ��*V���������;\������9���k��eȫ��%��(����௼,>�����*���lR��Ȭ��B��_��H���T���g���  �  ��N=64N=n�M=�L=,L=X}K=�J=<J=�mI=Y�H=�H=�[G=��F=��E=TIE=��D=M�C=�7C=V�B=��A=t%A=�s@=y�?=[?=JZ>=F�==F�<=J8<=p�;=��:=M:=AT9=ș8=��7=h#7=�g6==�5=N�4=o04=�q3=9�2=I�1=Z+1=e0=L�/=��.=�.=�/-=EZ,=�+=#�*=U�)=`�(=3�'=�'=5&=�%=!$=�#=�"=�!=�=%�=%�=�}=eF=�=4�=�h=&=ޥ=66=m�=�;=��=	=��=��	=�9=ۉ=F�=w=�S=��< y�<���< �<�d�<f��<x��<���<#�<�@�<IY�<�l�<�{�<D��<���<���<��<���<\��<���<���<���<ƈ�<��<�u�<*i�<-[�<�K�<�:�<�(�<�<!�<|��<Ƽy<@�q<�zi<�]a< DY<�-Q<�I<LA<a�8<�0<�(<	� <�<��<�<�� <5��;]��; ��;V��;j&�;O^�;ҥ�;���;��f;~�G;s);�b
;*��:ke�:{�>:mЎ9�;�RE$��I��f�ź�������Zd7�
�R���m��+���4������⁪�����A�»xkλ9�ٻ���o���a��dX�^�#C�������4������"��'��,+��%/�x3�i�6��x:��>��A��E�bH���K�f�N��#R��KU��iX��[�'�^�ԓa���d�D�g���j�Rmm��Sp� 3s�ev���x���{�Dq~�����:���aS��&������a�����,���l���ƌ�!���{�� א�<2��V���(蔼iB����������L��8�������4Q��7���q����S����������[�����?���m���ʫ�u(�������䯼gB����������3W�������
��Oc��I������gj���  �  ��N=�3N=��M=��L=,L=�}K=��J=J=oI=��H='H=n]G=��F=��E=NKE=ǚD=6�C=�9C=�B=��A=�&A=�t@=�?=�?=RZ>=�==��<=�7<=W;=h�:=�:=�R9=ؗ8=��7=R!7=|e6=/�5=L�4=�.4=�o3=ί2=�1=g*1=yd0=�/=��.=	.=80-=�Z,=�+=e�*=��)=
�(=�'=�	'='&=�%=�"$=S #=}"=�!=N�=
�=¬=�}=lF=�=��=h= =r�=�4=��=�9=D�=�=K�=l�	=e7=��=9�=�=�Q=��<�v�<��<��<Jd�<z��<>��<* �< %�<uC�<B\�<p�<��<T��<Ɠ�<���<��<_��<ٝ�<���<���<Ǒ�<P��<���<�u�<�h�<hZ�<CJ�<�8�<2&�<
�<���<��<C�y<��q<�qi<�Ta<];Y<�%Q<�I<�A<��8<J�0< �(<�� <��<��<P�<� <l��;=��;���;@
�;�5�;-o�;z��;��;��f;#�G;8&);��
;o�:c��:��>:[?�94;��2$�4J��+�ź�������v7���R���m�:���C�����ؑ��dѶ�s�»7yλ��ٻ���U���h���Z�h_�?C������t1����y�"��'��%+�!/�l�2�[�6��p:��>���A��D�\H�I�K�M�N�� R��IU�iX��[���^�3�a�`�d��g��j��sm��Zp�;s��v�2�x�V�{�my~�圀������V��а��
���b��$�������l��ƌ����7z���Ԑ��/��8����䔼�>���������H��O���N����M��f��� ���R������0���[��`��� ���n���̫��*������	诼%F������ ��p[���������g����������l���  �  ��N=�2N=��M=��L=,,L=�}K=1�J=�J=pI=̿H=bH=�^G=�F={�E=�LE=A�D=��C=�:C=�B=��A=r'A=Iu@=��?=�?=XZ>=ͤ==M�<=�6<=}~;=]�:=�:=7Q9=_�8==�7=�7=�c6=��5=��4=;-4=�n3=��2=&�1=�)1=�c0=��/=o�.=".=�0-=�[,=т+=]�*=��)=P�(=a�'=�
'=�&=>!%=`$$=�!#=�"=�!=9�=��=;�=G~=lF=�=2�=gg=
=X�=>3=�=8=��=�=r�=��	=�5=م=��==�P=��<u�<���<$�<�c�<���<���<,�<�&�<aE�<x^�<�r�<I��<D��<ٖ�<���<��<<��<���<ѝ�<���<S��<|��<���<7v�<�h�<�Y�<I�<7�<9$�<��<��<��<�y<
�q<�ji<Na<�4Y<�Q<�I<v�@<L�8<��0<B�(<�� <�<��<b�<� <���;���;���;��;�A�;�{�;�Ē;�;vg;�H;�>);Җ
;�>�:$��:�'?:9�:��$$��J��]�ź������g�7�B�R���m��D��O��t������ܶ���»��λ�ٻ�S��Sn���\�w`�QC�c���/�i��i�"��'�� +�w/���2�/�6��j:�>��A���D��WH�?�K��N�@R�,HU��hX��[���^�a�a�@�d���g���j��xm�B`p�*As��v���x���{�r~�㟀�]����X��񲄼���d�����<���l���Ō����x��!Ӑ��-��臓��ᔼ�;������혼�E��w�������bK��C�������P����������[���������#p��AΫ��,��ً���꯼�H������%���^��ϸ������i��=���-���n���  �  E�N=�2N=S�M=��L=-,L="~K=y�J== J=�pI=z�H='H=�_G=�F=t�E=�ME=4�D=��C=�;C=ފB=��A=�'A=�u@=��?=�?=OZ>=��==
�<=s6<=�};=��:=�
:=PP9=s�8=;�7=�7=�b6=��5=��4=O,4=�m3=��2=��1=<)1=�c0=f�/=V�.=1.=�0-=�[,=G�+=�*=��)=�(=@�'=�'=�&=9"%=M%$=�"#=|"=�	!=��=)�=��=d~=mF=[=�=�f=�	=��=r2=%�=7=t�=�=E=f�	=z4=ʄ=��=9=�O=j�<�s�<���<��<�c�<���<*��<��<i'�<�F�<�_�<>t�<��<,��<��<���<���<
��<��<M��<���<P��<(��<(��<Rv�<�h�<UY�<^H�<;6�<�"�<5�<K��<��<�y<��q<Zfi<�Ia<�0Y<�Q<-
I<W�@<��8<��0<��(<�� <g�<��<��</� <���;Z��;���;t�;+I�;���;;͒;'�;r%g;i$H;N);��
;�V�:ɛ:�I?:Ï9�r:��$��K����ź��������7�
 S�Qn��K���V��x ��ᥪ�	嶻0�»��λF�ٻT廯��iq���]�a��C�����-�t��#�"��'�r+��/���2�)�6��f:�'�=�N�A���D��TH���K�,�N��R�kGU�4hX�3�[�e�^���a��d�ԗg�:�j��{m��cp��Ds��v���x��{���~�����/����Z��?�������d����������l��oŌ����4x��$Ґ�H,��f���Z����9��"����똼�C���������I��ܠ������O�����6��u[��ض��L���p��!ϫ�.��@���J쯼�J������D���`�������k���º����)p���  �  �N=W2N=A�M=��L=3,L=0~K=��J=l J=�pI=��H=dH=�_G=a�F=��E="NE=~�D=��C=<C= �B=��A=(A=�u@=��?=?=SZ>=��==��<=H6<=�};=z�:=�
:=P9=+�8=��7=^7=�b6=@�5=��4= ,4=�m3=ǭ2=X�1=)1=oc0=P�/=K�.=E.=�0-=�[,=u�+=�*=��)=N�(=��'=+'=�&=~"%=�%$=�"#=�"=�	!=��=Q�=��=s~=F=L=Ժ=�f=`	=i�=22=ڸ=�6=#�=X=�~=�	=4={�=D�=�=�O=��<�s�<���<��<�c�<Ϡ�<L��<&�<�'�<�F�<z`�<�t�<���<Đ�<��<G��<���<���<���<џ�<��<���<]��<H��<av�<�h�<(Y�<H�<�5�<t"�<��<���<�<��y<�q<1ei<*Ha<\/Y<TQ< 	I<m�@<��8<��0<��(<l� <I�<��<E�<�� <Q��;���;���;��;�K�;���;�ϒ;�)�;�*g;*H;�R);��
;_�:�ϛ:�V?:1Ϗ9�Z:��$��L��@�ź���ع�G�7��S��
n�N��[Y���"�������綻r�»,�λ[�ٻ��n���r��[^�]a��C���Ǩ� -����g�"�o
'��+��/�m�2��6�be:���=�#�A���D��SH�4�K�x�N�JR�GU��gX�P�[���^��a���d���g��j��|m�.ep��Es�B v���x��{��~�C��������Z������K��9e��Ἀ�����l��@Ō�o���w���ѐ��+��م���ߔ�\9������,똼SC��蚛�B�bI��Y�������UO��ʧ����a[����s��-q���ϫ��.�������쯼nK��*������Da���������gl���ú�	���p���  �  E�N=�2N=S�M=��L=-,L="~K=y�J== J=�pI=z�H='H=�_G=�F=t�E=�ME=4�D=��C=�;C=ފB=��A=�'A=�u@=��?=�?=OZ>=��==
�<=s6<=�};=��:=�
:=PP9=s�8=;�7=�7=�b6=��5=��4=O,4=�m3=��2=��1=<)1=�c0=f�/=V�.=1.=�0-=�[,=G�+=�*=��)=�(=@�'=�'=�&=9"%=M%$=�"#=|"=�	!=��=*�=��=e~=oF=]=�=g=�	=��=v2=*�=7=z�=�=N=o�	=�4=Մ=��=E=�O=��<t�<��<��<�c�<���<B��<��<}'�<�F�<�_�<Jt�<(��<1��<��<���<��<��<��<>��<���<=��<��<��<;v�<�h�<>Y�<HH�<&6�<�"�<%�<>��<��<کy<��q<Zfi<�Ia<�0Y<�Q<G
I<w�@<��8<��0<��(<�� <��<�<)�<Z� <���;���;���;��;QI�;ڃ�;E͒;'�;K%g;#$H;�M);}�
;�U�:�Ǜ:�F?:���9r�:��#$��M��m�źk	��w��r�7�� S�%n�3L��W��� ��/���P嶻p�»�λx�ٻ����ﻊq���]�a��C��%���-�y��'�"��'�u+��/���2�*�6��f:�'�=�O�A���D��TH���K�,�N��R�kGU�4hX�3�[�e�^���a��d�ԗg�:�j��{m��cp��Ds��v���x��{���~�����/����Z��?�������d����������l��oŌ����4x��$Ґ�H,��f���Z����9��"����똼�C���������I��ܠ������O�����6��u[��ض��L���p��!ϫ�.��@���J쯼�J������D���`�������k���º����)p���  �  ��N=�2N=��M=��L=,,L=�}K=1�J=�J=pI=̿H=bH=�^G=�F={�E=�LE=A�D=��C=�:C=�B=��A=r'A=Iu@=��?=�?=XZ>=ͤ==M�<=�6<=}~;=]�:=�:=7Q9=_�8==�7=�7=�c6=��5=��4=;-4=�n3=��2=&�1=�)1=�c0=��/=o�.=".=�0-=�[,=т+=]�*=��)=P�(=a�'=�
'=�&=?!%=`$$=�!#=�"=�!=:�=��==�=I~=nF=�=6�=kg= 
=_�=G3=�=8=��=�=��=��	=�5=�=��=6=�P=��<9u�<���<Y�<.d�< �<��<X�<�&�<�E�<�^�<�r�<Y��<M��<ܖ�<���<���<+��<h��<���<o��<-��<S��<���<v�<�h�<�Y�<�H�<�6�<$�<��<���<��<ѭy<��q<�ji<&Na<�4Y<�Q<I<��@<��8<��0<��(<� <^�<D�<��<[� <���;���;W��;7�;�A�;�{�;�Ē;��;)g;H;>);��
;J<�:���:�!?:H��9��:��+$�`N���ź������%�7���R���m��E���O��������wݶ�x�»�λu�ٻo廝�ﻒn���\��`�eC�t����#/�r��q�"��'�� +�|/���2�1�6��j:�>��A���D��WH�@�K��N�AR�,HU��hX��[���^�a�a�@�d���g���j��xm�B`p�*As��v���x���{�r~�㟀�]����X��񲄼���d�����<���l���Ō����x��!Ӑ��-��臓��ᔼ�;������혼�E��w�������bK��C�������P����������[���������#p��AΫ��,��ً���꯼�H������%���^��ϸ������i��=���-���n���  �  ��N=�3N=��M=��L=,L=�}K=��J=J=oI=��H='H=n]G=��F=��E=NKE=ǚD=6�C=�9C=�B=��A=�&A=�t@=�?=�?=RZ>=�==��<=�7<=W;=h�:=�:=�R9=ؗ8=��7=R!7=|e6=/�5=L�4=�.4=�o3=ί2=�1=g*1=yd0=�/=��.=	.=80-=�Z,=�+=e�*=��)=
�(=�'=�	'=(&=�%=�"$=T #=}"=�!=O�=�=Ĭ= ~=pF=�=��=$h=	=|�=�4=��=�9=V�=�=b�=��	=�7=��=Y�=�=R=*�<w�<S��<<�<�d�<���<���<h �<8%�<�C�<k\�</p�<��<a��<ɓ�<���<��<F��<���<`��<W��<���<��<���<�u�<�h�<+Z�<J�<w8�< &�<��<���<�<�y<��q<�qi<�Ta<�;Y<�%Q<�I< A<!�8<��0<��(<9� <]�<R�<��<�� <J��;��;���;�
�;`6�;po�;���;��;y�f;f�G;,%);.
;:�:���:��>:z-�9:E;�r<$�MO��S�ź
���A��}x7�[�R���m�;���D��q������&Ҷ�!�»�yλ/�ٻ 廽��(i���Z��_�[C������1������"�'��%+�'/�q�2�_�6��p:��>���A��D�\H�J�K�N�N�� R��IU�iX��[���^�3�a�`�d��g��j��sm��Zp�;s��v�2�x�V�{�my~�圀������V��а��
���b��$�������l��ƌ����7z���Ԑ��/��8����䔼�>���������H��O���N����M��f��� ���R������0���[��`��� ���n���̫��*������	诼%F������ ��p[���������g����������l���  �  ��N=64N=n�M=�L=,L=X}K=�J=<J=�mI=Y�H=�H=�[G=��F=��E=TIE=��D=M�C=�7C=V�B=��A=t%A=�s@=y�?=[?=JZ>=F�==F�<=J8<=p�;=��:=M:=AT9=ș8=��7=h#7=�g6==�5=N�4=o04=�q3=9�2=I�1=Z+1=e0=L�/=��.=�.=�/-=EZ,=�+=#�*=U�)=`�(=3�'=�'=6&=�%=!$=�#=�"=�!=�=(�=(�=�}=jF=�=;�=�h=0=�=D6=~�=�;=��="=Մ=��	=�9= �=m�=�=�S=�<\y�< ��<g �<e�<���<���<)��<Z#�<9A�<{Y�<�l�<�{�<T��<ď�<x��<��<v��<3��<R��<���<z��<��<��<;u�<�h�<�Z�<@K�<f:�<p(�<��<��<Z��<��y<(�q<�zi<�]a<NDY<6.Q<AI<�A<��8<��0<�(<�� <��<\�<��<� <E��;P��;���;��;�&�;�^�;���;���;#�f;��G;+);a
;<��:�`�:g�>:���9��;�zQ$��O����ź,������`g7���R���m�-���5��
���肪��¶��»6lλ��ٻ������Lb���X�B^�EC��í��4�Ɲ���"�	'��,+��%/�~3�n�6��x:��>��A��E�bH���K�g�N��#R��KU��iX��[�'�^�ԓa���d�D�g���j�Rmm��Sp� 3s�ev���x���{�Dq~�����:���aS��&������a�����,���l���ƌ�!���{�� א�<2��V���(蔼iB����������L��8�������4Q��7���q����S����������[�����?���m���ʫ�u(�������䯼gB����������3W�������
��Oc��I������gj���  �  ��N=5N=��M=A�L=�+L=�|K=>�J=J=�lI=��H=�
H=�YG=��F=��E=�FE=o�D=�C=�5C=x�B=��A="$A=�r@=��?=�?=?Z>=��==��<=89<=��;=5�:=:=LV9=�8=�7=�%7=�i6=��5=��4=�24=os3=ݲ2=��1=l,1=�e0=��/=��.=�.==/-=\Y,=�+=��*=��)=p�(=�'=T'=�&=�%=�$=|#=�"=�!=��=�=\�=A}=UF=F=�=�i=�=��=.8=��=B>=5�=�!=��=��	=�<=��=��=�=�U=T�<|�<���<�!�<�e�<���<���<���<!�<\>�<�U�<�h�<�w�<���<���<���<H��<��<��<���<���<ߌ�<���<~�<�t�<i�<�[�<�L�<�<�<=+�<E�<��<��<�y<.�q<��i<�ga<(NY<}7Q<$I<vA<i9<��0<,�(<d� <�<E�</�<� <>��;���;���;���;�;9K�;���;��;��f;��G;t�(;�=
;���:;+�:�E>:/�9o�<��i$��P��Y�ź����U���S7��R���m�����$��T읻#q�������»�\λy�ٻa����ﻋZ��V��\�C�I	�1���8�֢���"�b '��4+�F./��3���6�=�:�&>���A�E�tiH���K�c�N�z'R�0NU�kX�5[���^��a���d���g�+zj��em�PKp�Y*s��v�1�x�a�{��g~�����󁼶O�����O��#_��ɸ������l��Bǌ�d"���}���ِ�]5�����2씼�F�����������Q���������U������B ��*V���������;\������9���k��eȫ��%��(����௼,>�����*���lR��Ȭ��B��_��H���T���g���  �  ��N=�5N=��M=k�L=�+L=^|K=g�J=�J=kI=عH=�H=BWG=�F=�E=_DE=�D=��C=�3C=x�B=8�A=�"A=�q@=��?=�?=$Z>=ϥ==��<=/:<=�;=��:=�:=nX9=E�8=��7=\(7=�l6=&�5=��4=�44=gu3=��2=�1=�-1=�f0=&�/=��.=W.=�.-=jX,=�~+=�*=��)=X�(=��'=�'=i&=%=q$=3#=�"=!=7�=��=��=�|=4F=�=|�=�j=�=?�=<:=�=�@=��=�$=��=��	=�?=V�=w�=&=�W=��<�~�<���<�"�<"f�<D��<���<���<��<+;�<=R�<�d�<�r�<�}�<���<|��<8��<6��<���<���<!��<��<s��<}�<�s�<i�<�\�<[N�<�>�<:.�<��<-�<s��<+�y<�q<��i<�ra<�XY<�AQ<9-I<�A<l9<��0<��(<,� <E�<��<b�<�� <���;h��;���;t��;j�;6�;g{�;ӂ;�~f;��G;��(;�
;C[�:p�:\�=:���9�f=�,�$��S����źʸ���z��=7�>�R�K�m�������[ٝ�^�����m�»�Kλķٻk��d�ﻞR��0S��[�=C��
�����<�I����"�('��=+��7/��3�K�6���:�$>�N�A��E�(qH�L�K���N��+R��PU�llX�7[�&�^��a�e�d�t�g�Rsj�^m�vBp�� s���u���x�)�{��]~�������K��ɧ�����&]��r�������l��Ȍ��#�����oܐ��8�������𔼕K�����������V���������7Y��Z���b���X��p���	���\��i���@��3j��ƫ��"������ܯ��9��'����MM������]��tZ��������md���  �  �N=�6N= �M=��L=�+L=�{K={�J=�J=siI=�H=xH=�TG=��F=��E=�AE=c�D=A�C=N1C=q�B=s�A=0!A=p@=�?=?=
Z>=�==�<=;<=1�;=i�:=�:=�Z9=��8=
�7=�*7=$o6=��5=U�4=�64=]w3=U�2=}�1=�.1=^g0=��/=��.=.=�--=lW,=Q}+=n�*=׽)=3�(=x�'=w '=�&=�%=$=�#=�"=D!=��=��=��=;|=F=�=�=�k=.=�=C<=M�=dC=ù=�'=��=��	=kB=�=��=n=�Y= �<Y��<���<$�<�f�<���<���<���<�<�7�<xN�<6`�<n�<�x�<���<@��<��<Y��<4��<���<���<Q��<D��<�{�<Fs�<i�<F]�<�O�<	A�<,1�<y �<L�<��<O�y<w�q<��i<�}a<3cY<oKQ<,6I<�#A<F9<�1<��(<�� <t�<��<g�<:� <��;���;a��;���;��;� �;e�;d��;0Qf;�VG;'�(;��	;��:��:Є=:��9g9>�գ$��V��L�ź����)k��(7�q�R�nvm������ ��lƝ��J��x���\�»*;λ�ٻ�������J���P�ZZ�[C�B����@�ҭ���"��/'�uF+�|A/��!3���6���:�:.>��A��E��xH�&�K�S O��/R��SU��mX�*[���^�K�a�O�d��|g��lj�MVm��9p�=s���u���x��{�T~�<����ꁼ/H������ ��D[��8���d���l���Ȍ��%��C���Sߐ�V<������ ���iP����������[������h��u]��
������![��W���?��]��)���T���h���ë����|���د�5��M����H�����������U�������ga���  �  :�N=�7N=q�M=��L=F+L=B{K=��J=�J=�gI=F�H=uH=�RG=V�F=*�E=l?E=�D=�C=2/C=|B=��A=�A=bo@=T�?=�?=�Y>=>�==��<=�;<=^�;=��:=�:=v\9=��8=M�7=>-7=�q6=�5=��4=�84=7y3=�2=��1=�/1=h0=�/=��.=� .=N--=tV,=|+=�*=�)=+�(=W�'=(�&=�&=7%=�$=�#=�"=� =3�=}�=Ψ=�{=�E=�=��=�l=n=|�=>=w�=�E=E�=V*=K�=j�	=E=��=U�=�=�[=&#�<Ճ�<���<&%�<�f�<���<���<)��<��<�4�<�J�<!\�<�i�<�s�<�{�<Y��<R��<ڇ�<눹<܈�<i��<���<1��<8z�<~r�<i�<�]�<7Q�<%C�<�3�<�#�<*�<^�<��y<B�q<��i<��a<�lY<mTQ<�>I<�*A<u9<
1<Q�(<� <Q�<��<l�<�� <Q��;m��;���;���;=۱;��;P�;?��;�&f;�-G;Vd(;B�	;+��:e}�:�'=:�q�9�
?���$�hZ��s�źB���n\��7�!lR��Zm�Y샻�
���9�� z��v»,λ2�ٻ	�仉�ﻚC��iN�OY��C�����E�'���#�u7'��N+�LJ/�\+3�L�6���:��7>���A��%E�v�H�{�K��O��3R��VU�XoX�l[���^��a�l�d��wg��fj��Nm��1p��s���u�<�x���{��J~�����恼�D����������rY��(������7m���Ɍ� '��m���␼�?��՜��S����T��o�������`��-�������a�������	���]��(���j���]�������g����������x���ԯ�1��ጲ�j購dC����������Q��B�������^���  �  �N=58N=ĉM=��L=+L=�zK=��J=wJ=�fI=´H=�H=�PG=K�F=�E=N=E=�D=��C=V-C=�}B=L�A=�A=dn@=��?=!?=�Y>=`�==��<=�<<=M�;=�:=�:= ^9=��8=C�7=?/7=}s6=��5=d�4=�:4=�z3=6�2=��1=e01=�h0="�/=��.=h .=�,-=�U,=�z+=��*=r�)=t�(=h�'=(�&=�	&=)%=�$=�#=%"=�� =��=s�=�=M{=�E==�=�m=n=ŭ=�?=C�=�G=q�=�,=��=��	=`G=Ö=U�=W!=]=�%�<υ�<���<�%�<g�<��<���<���<v�<62�<�G�<�X�<�e�<�o�<nw�<}�<��<׃�<T��<���<���<@��<s~�<y�<�q�<i�<k^�<TR�<�D�< 6�<�&�<t�<�<��y<��q< �i<+�a<%uY<?\Q<�EI<!1A<�9<-1<R�(<�� <��<b�<��<�� <�;��;��;*��;�ʱ;@��;�=�;���;�f;B	G;JB(;3�	;B��:M�:*�<:���9@�?�m�$�+^��>�ź�����P�+7�LXR��Bm�
߃�[ᐻ���*���j���g»�λ��ٻ�令���=��~L��X�	D�y�S���H���d	#��='��U+�DR/��33���6�$�:� @>���A�-E���H��K�F
O�i7R��XU��pX��[���^�҆a�`�d��sg�Iaj��Hm��*p�+s���u�J�x��{{�C~�X���Cぼ�A���������X��G������lm���ʌ�D(��X���{䐼�B��$��������X����������d��C�������d������#���_������j��1^��񴧼����e��񿫼���v���ѯ�q-�����]䳼o?������/���+N�������U\���  �  ��N=�8N=
�M=��L=�*L=[zK==�J=�J=�eI=��H=wH=wOG=ɝF=��E=�;E=h�D=w�C=�+C=�|B=%�A=�A=�m@=�?=�?=�Y>=v�==Q�<=*=<=�;=�:=:=f_9=�8=��7=�07=u6=k�5=��4=<4=�{3==�2=��1=11=i0=P�/=��.=- .=D,-=�T,=z+=��*==�)=!�(=��'=��&=�&=�%=F$=o#=�
"=�� =��=��=q�=�z=�E=-=W�=n=3=Ů=�@=��=JI=�=U.=\�=��	=I=f�=��=�"=I^=�'�<N��<��<�&�<@g�<���<���<?��<��<0�<6E�<�U�<�b�<�l�<$t�<�y�<�}�<ʀ�<���<��<j��<j��<�|�<�w�<Sq�<�h�<�^�<<S�<F�<�7�<�(�<��<��<|�y<�q<s�i<��a<9{Y<bQ<�JI<�5A<�"9<<1<�)<D� <u�<��<�<k� <��;���;ӌ�;��;w��;#�;B0�;6��;Q�e;��F;�((;��	;�r�:_'�:�<:���94N@���$�1a���źx���G�"�6�6IR�\0m��ԃ��֐���������_��?]»�λ��ٻk��m��}9���J�-X�;D���|���K�����#��B'�p[+�_X/��93�<7���:�F>���A��2E��H�t�K��O�F:R�[U��qX��[�,�^�*�a�~d��pg�@]j�{Dm��%p��s���u�3�x�zu{�_=~����������?��)���K����V������j���m��Pˌ�m)��݇��_搼�D�����������[���������g��F���}���g�����2��ka�����P	���^��ߴ��q���d����������s��Mϯ��*��?���e᳼g<������_�wK�����������Z���  �  2�N=�8N=2�M=��L=�*L=zK=��J=,J=eI=زH=� H=�NG=ϜF=x�E=�:E=Y�D=��C=+C=�{B=r�A=�A=.m@=��?=�?=�Y>=�==|�<=y=<=y�;=��:=�:=+`9=Ȧ8=��7=�17=v6=^�5=��4=�<4=�|3=ֺ2=,�1=c11=<i0=n�/=��.= .=�+-=�T,=�y+=�*={�)=:�(=�'=��&=�&=�%=A$=�#=�	"=� =M�=&�=�=�z=}E=0=��=fn=�=^�=�A=t�=9J=�=n/=��=��	=$J=l�=��=�#=�^=�(�<1��<���<�&�<;g�<���<U��<���<��<�.�<�C�<T�<�`�<�j�<r�<�w�<�{�<�~�<���<x��<��<]�<(|�<nw�< q�<�h�<_�<�S�<�F�<�8�<
*�<��<�
�<j�y<�q<Ƿi<��a<DY<�eQ<TNI<�8A<%9<51<�)<
� <��<v�<,�<�� <��;5��;���;���;���;��;'�;<}�;��e;��F;�(; �	;GX�:�:\s<:V�9��@���$�fc����źq���A���6��>R�%m�Z΃��ϐ�C�������X��9V»�λE�ٻ��ǔﻰ6��AJ��W��D�J����KM�����#�!F'�(_+�\/��=3�u7�ͳ:�TJ>���A�A6E��H�#�K�O��;R�N\U��rX��[�Ʌ^�h�a��|d��ng��Zj�Am�p"p���r�&�u�)�x��q{��9~��~�� ߁�>�����]���IV��2���O���m���ˌ�*�������琼)F��I�������]���������i��D���S��Zi������|��cb��Ƶ���	���^��촧�)��{d��ҽ������r���ͯ�)��a���}߳�\:�����|﷼�I���������~Y���  �  9�N=�AN=�M=8�L=�5L=r�K=o�J=�"J=�pI=�H=�H=B[G=(�F=��E=JE=^�D=a�C=�?C=�B=I�A=`9A=<�@=s�?=�/?=U�>=��====Jk<=��;=�;=QM:=��9=�8=|(8=?p7=f�6=��5=VC5=��4=��3=�3=�L2=��1=�0=��/=�4/=�g.=��-=��,=6�+=�+=1*=QN)=�g(=^}'=��&=��%=�$=Ѧ#=�"=��!=a� =qr=QR=Z)= �="�=<u=%=��=>f=��==��=Cq=��=U?=ę
=V�=a7=5{=P�=��=a =œ�<���<��<"R�<~�<��<S��<���<���<���<���<���<4��<���<���<���<�߽<�ڹ<<յ<�α<Dǭ<���<O��<J��<m��<���<&y�<*f�<�Q�<+<�<�%�<3�<?�y<-�q<^�i<�ma<mEY<�Q<	�H<��@<ض8<��0<y(<�\ <
@<@$<Y	<$��;���;��;Fe�;�N�;�F�;�N�;rj�;?7;��_;��@;o�!;3�;RC�:�}�:�X:_[9ix���F�3z��-Z׺�P���$�ѕ@�Z(\��Qw�����!��h ��^������ǻ��ӻ�@߻�r��[��r���R+�V5
��������*�g{!���%���)���-���1��5��w9��=�#�@�eD�7[G���J���M�p�P��
T��W��Z��]��`���b��e�P�h�y�k��xn��Lq�Rt�d�v���y�k|�S'���J��f���4����U��������>`����������q���Ώ�,��=���擼�A��v���_���yL��d���Z����E�������䟼n3�����cѣ��!��,s��1Ƨ�����p���ǫ�E ��Gy���ү��,��'����߳��8�������鷼:B��n����򻼆K���  �  �N=�AN=�M=5�L=�5L=��K=��J=&#J=BqI=9�H=DH=�[G=��F=;�E=�JE=ۛD=��C=`@C=^�B=��A=�9A=|�@=��?= 0?=c�>=��====-k<=S�;=�;=M:=��9=��8=(8=�o7=��6=X�5=�B5=i�4=��3=w3=rL2=h�1=��0=��/=�4/=�g.= �-= �,=��+=H+=W1*=�N)=3h(=�}'=:�&=3�%=W�$=0�#=M�"=��!=�� =�r=�R=|)=(�=�=&u=�$=��=�e=B�=�~=^�=�p=�=�>=B�
=��=�6=�z=�=��= =S��<c��<��<R�<~�<F��<���<��<[��<���<���<���<#��<���<���<s��<��<�۹<�յ<vϱ<�ǭ<��<���<���<���<���<y�<�e�<1Q�<�;�<=%�<��<z�y<i�q<��i<la<�CY<Q<��H<F�@<��8<��0<�x(<\ <�?<H$<�	<���;���;���;�g�;�Q�;�I�;aR�;�n�;�@;��_;ۗ@;�!;!�;P�:1��:�n:��9#_��6F��w���X׺�P�b�$���@�,\��Uw�=���$��<��n���'���ȻC�ӻ�B߻�t껚]������z+�p5
������<��/�$z!�U�%�^�)�b�-�E�1�M�5��u9��=�Q�@��D��YG�J�J���M�9�P��	T��W��Z��]��`���b���e�L�h���k��yn�Nq�t��v�5�y��l|�)������K���������V��S������H`����������q��OΏ�|+������c哼%A������m���cK��[������D��𔞼䟼�2�������У�X!��s��4Ƨ�����p��Sȫ�� ���y���ӯ�H-������೼�9��m����근�B�����D�
L���  �  y�N=mAN=��M=9�L=�5L=�K=)�J=�#J=rI=9�H=lH=�\G=�F=��E=�KE=4�D=�C=�AC=~�B=��A=�:A=�@=�?=M0?=��>=��==�==�j<=��;=�;=L:=��9=��8=�&8=�n7=��6=�5=�A5=S�4=��3=�3=�K2=�1=��0=��/=�4/=�g.=��-=��,==�+=0+=`2*=�O)=wi(='=��&=��%=��$=p�#=u�"=��!=�� =hs=S=�)=L�=�=�t=�$=��=%e=D�=w}=�=Uo=��=Q==ė
=Z�=u5=~y=��=��=6 =��<p��<4�<�Q�<>~�<��<���<j��<��<���<��<��<���<���<h��<9��<}�<0޹<'ص<jѱ<}ɭ<\��<���<"��<ƚ�<{��<�x�<�d�<�O�<�9�<0#�<9�<[�y<2�q<�i<�fa</>Y<	Q<�H<)�@<^�8<��0<w(<�Z <p?<�$<�
<M��;���;n��;�o�;w[�;�T�;�]�;�z�;BX;��_;ï@;�!;Y�;�u�:���:c�:_X9y����E��r��RZ׺T���$���@��8\��cw�f���-��W��ާ��:���$ȻL�ӻ@J߻�z�%b���  �w,��5
��q��s����w!���%��)���-��1��5�:p9� =��@���C��TG���J���M�$�P��T�W��Z�]�$`��b���e���h�ʣk��}n�KRq��!t��v�N�y��q|��-�"󀼘M��馃�>���>W��!���|��r`��;������p��͏��)������*㓼�>������񗼺H��������`B������
⟼ 1��4����ϣ�� ���r��Ƨ�/���q��\ɫ�"���{���կ��/��{���㳼:<��锶�C�6E��������cM���  �  ��N=�@N=Y�M=2�L=66L=u�K=��J=�$J=rsI=��H=.H=�^G=��F=��E=&NE=W�D=(�C=CC==�B=�A=�;A=&�@=��?=�0?=��>=��==\==j<=ϵ;=� ;=�J:=��9=��8=�$8=�l7=��6=�5=�?5=��4=%�3=L
3=�J2=!�1=#�0=��/=�4/==h.='�-=��,=d�+=�+=
4*=�Q)=pk(=2�'=��&=��%=��$=e�#=0�"=��!=�� ={t=�S=S*=��=�=�t=�#=��=�c=��=�{=�=%m=O�=�:=Y�
=�=E3=tw=�=��=� = ��<���<e�<�Q�<�~�<��<E��<���<���<���<���<(��<��<��<���<���<��<��<�۵<gԱ<̭<Y©<	��<�<���<��<xw�<Bc�<�M�< 7�<��<��<e�y<��q<;�i<�]a<�5Y<+Q<��H<��@<�8<��0<�s(<�X <�><D%<�<p��;e��;.��;'}�;?j�;�d�;�o�;Z��;;`;Z�@;��!;.�;.��:�ߋ:��:�m9:���|�E��k��^׺�Z���$���@�&L\�{w�f���;�����9���9��ȻR�ӻ�U߻����i��_ �R.�d6
�����������7r!�ȹ%�-�)�7�-���1�J�5�eg9�I=�Y�@�s�C�wMG�&�J� �M�S�P��T�rW��Z��]��`��b���e���h��k�уn�4Yq�Q)t��v���y�
z|��5������P��٩�����1Y������]���`��񹋼��;o��ˏ�\'�������ߓ��:��󔖼v헼UD��T����웼x>������ޟ�J.���}��.Σ�w��r�� Ƨ�����r��˫�`$��`~���د�3��L���糼`@�������H��N��������O���  �  m�N=�?N=�M=�L=�6L=#�K=��J=R&J=%uI=��H=�H=daG=��F=~ F=QE=�D=��C=�EC=��B=�A=q=A=z�@=��?=d1?=�>=y�==�==4i<=��;=�:=�H:=Ñ9=F�8=G"8=�i7=��6=r�5=M=5=@�4=�3=�3=RI2=�1=s�0=9�/=�4/=�h.=�-=��,=��+=Y+=$6*= T)=n(=ك'=m�&=d�%=W�$=�#=��"=��!=�� =�u=�T=�*=��=պ=�s=�"=��=%b=��=Hy=]�=@j==�=�7=?�
=��=]0=�t=��=��=3 =P��<��<U�<[Q�<5�<*��<]��<l��<W��<��<n��<b��<���<���<���</��<��<��<�<5ر<Hϭ<�ĩ<θ�<瑱<,��<���<v�<"a�<�J�<�3�<��<��<��y<e�q<�|i<�Ra<�*Y<�Q<S�H<��@<ڥ8<,�0<�o(<rV <�=<�%<�<��;���;��;��;�}�;�z�;��;o��;h�;�B`;�A;��!;�!;(��:1!�:k:-�96���E�=d���b׺�c�^�$�n�@�$f\�H�w��,���N��2/���ʯ� ���+Ȼ��ӻ�d߻���Ot�� ��0�+7
�����@����k!�]�%�u�)��-�J�1�Z�5�\9���<�i}@���C��CG�m�J���M��P���S�!W�Z�]��	`���b���e�`�h�֯k�͋n�dbq�;3t���v�3�y���|�K@�����rU������
���[��q���n	��a���������qm���ȏ�$$�����=ۓ�6������ 藼�>��ʓ��C盼S9��a����ڟ��*��{��̣���`q��5Ƨ�~��St��Oͫ�['�������ܯ��7��\���k쳼�E��U���7����M�����������R���  �  ��N=�>N=[�M= �L=�6L=��K=*�J=�'J=#wI=)�H=$H=JdG=ʳF=�F=ATE=M�D=��C=�HC=�B=M�A=W?A=��@=��?=2?=(�>=<�==4==h<=�;="�:=sF:=1�9=o�8=>8=�f7=ĭ6=]�5=^:5=�4=��3=�3=�G2=Ɇ1=��0=��/=5/=i.=͙-=��,=��+=n+=�8*=�V)=�p(=��'=��&=��%=q�$=ѯ#=(�"=�!=�� =tw=�U=�+=�=��=Is=�!=�=`=4�=wv=A�=�f=��=4=��
=d�=�,=�q=��=w�=, =��<���<��<�P�<��<���<���<���<n��<���<���<f�<��<t �<.��<���<!�<��<3�<�ܱ<�ҭ<�ǩ<���< ��<Y��<Ĉ�<ct�<{^�<JG�<0/�<��<���<b�y<F�q<joi<Ea<�Y<��P<8�H<��@<��8<n�0<�j(<LS <�<<�&<�<��;��;L��;?��;��;t��;���;���;��;�|`;=A;.";�Q;S�:m�:��:wQ9թ��ϋE�=^���j׺/o���$��@���\���w��A��:e���F���⯻%7���AȻ�Ի�v߻͠껭���� ��3��8
������\����d!���%���)�E�-�?�1�{�5��N9���<��p@���C��8G��J��M���P���S�W
W�Z�]�j`���b���e���h�Էk�Q�n��lq��>t��
w���y�e�|�wL�j���Z��V�������^�������
���a��=������[k���ŏ�p ��o{��1֓�[0�������ᗼ#8��L�������y3������՟��&���w���ɣ�v���p��UƧ����;v��Ы��*��B����᯼M=��R�����L������8���"S����������eV���  �  l�N=�=N=��M=��L=7L=��K=c�J=�)J=7yI=��H=�H=[gG=�F=.F=�WE=��D="�C=�KC=ʝB=��A=OAA=}�@=�?=�2?=S�>=��==s==�f<=a�;=�:=�C:=]�9=L�8=�8=Oc7=Z�6=�5=%75=�|4=�3==3=�E2=[�1=��0=>�/=�4/=|i.=��-=R�,=T�+=�+=;*=�Y)=t(=G�'=��&=�%=��$=ݲ#=��"=h�!=�� =y=(W=`,=2�=\�={r=� =E�=�]=��=fs=��=(c=��=-0=��
=��=F)==n=��=��=� =���<K��<S�<qP�<��<%��<#��<��<���<��<��<��<��<x�<D�<���<���<��<��<N�<�֭<�ʩ<���<���<V��<ɇ�<�r�<�[�<iC�<q*�<
�<���<ٽy<2�q<�`i<�6a<�Y<,�P<�H<�@<��8<|0<ue(<�O <;<'<<6 <��;a��;ȵ�;ϫ�;���;y��;�ߏ;��;�`;�wA;�e";�;��:Ի�:ki :L� 9���kcE�~Z���u׺
|���$���@��\�2�w�]X��_}���_��R���*P��ZȻ&Ի��߻���t���� ��6�!:
�H����b{����d]!���%��)�l�-���1�ۊ5��@9���<��b@��C��,G�uJ��M���P���S�wW�6Z��]�K`�Wc� �e�(�h���k���n��xq��Kt�#w���y��|��Y����]`��\���#��Ob��?���r��Xb���������7i��������v���Г�Z*�� ����ڗ�71��c���Xڛ�N-��W���П��"��zt��ǣ����
p���Ƨ����Lx��ӫ��.��􊮼K篼_C��͞��T����R��P������EY��������aZ���  �  ��N=�<N=��M=��L=S7L=I�K=��J=+J=;{I=�H=�H=pjG=X�F=�
F="[E=�D=^�C=�NC=|�B=�A=>CA=��@=�?==3?=s�>=��==�==�e<=��;=��:=xA:=��9=4�8=�8=�_7=�6=��5=�35=�y4=_�3=�3=�C2=�1=��0=��/=�4/=�i.=~�-=��,=�+=�+=�=*=k\)=#w(=��'=P�&=A�%=�$=�#=��"=֦!=�� =�z=HX=�,=_�=�=�q=)=u�=�[=��=Np=d�={_=��=0,=��
=��=�%=�j=��=�=� =���<���<��<�O�<}��<s��<���<b��<���<�<�	�< �<��<e�<-�<Z�<  �<���<��<��<_ڭ<Jͩ<���<ୡ<<��<���<^p�<�X�<o?�<�%�<g�<j�<>�y<�q<3Ri<�'a<�Y<��P<׿H<$�@<7�8<�t0<�_(<+L <m9<�'<i<� <���;���;��;Sÿ;.ȯ;�ڟ;=��;$2�;��`;��A;<�";��;��:,	�:�� :j"9ᖝ��>E�-W����׺��� �$��A��\�6x��n������y��R���i��>rȻ�.ԻӞ߻��t���L ��:��;
�B�����w�e��V!���%���)���-���1��}5�E39��<��U@�2�C�� G��jJ��M�t�P�~�S��W�bZ�%]�,`�Fc���e���h���k�=�n���q�^Xt��%w�f�y�Ĭ|�g����%f��r�������e��빇�3��c��ݸ�����Kg��¿�����-r��~˓�c$���|��ԗ�b*������ӛ�'���y��̟�d��&q���ģ�m��so��ǧ� ���z��:֫��2�����쯼rI��P���7 ���Y��4���J	��b_�������	��~^���  �  G�N=�;N=H�M=@�L=y7L=�K=��J=�,J=}I==�H=<H=<mG=[�F=�F=Q^E=/�D=W D=�QC=�B=!�A=�DA=Y�@=��?=�3?=|�>=3�==�==bd<=�;=��:=?:=Ά9=D�8={8=�\7=��6=h�5=�05=�v4=ݻ3=��2=B2=v�1=��0="�/=�4/=-j.=5�-=��,=��+=�+=�?*=�^)=�y(=��'=o�&=]�%=�$=��#=D�"=�!=�� =|=LY=�-=}�=��=�p=�=��=zY==�=hm=&�=\=@�=s(=��
=��=("=�g=��=��=� =��<��<�<O�<ǀ�<���<���<b��<���<��<��<��<��<��<��<��<�<��<���<��<�ݭ<�ϩ<��<���<���<���<In�<�U�<�;�<� �<�<{�<[�y<!rq<sDi<+a<6�X<U�P<Y�H<�@<Y�8<�m0<>Z(<�H <�7<�'<{<w
 <���;��;���;�ؿ;9�;���;��;KN�;5-a;d�A;��";	�;�Z�:"O�:\!:�#9���"E��V����׺���%��3A�x�\�I7x�����z�������.��#���0�ȻDԻ��߻������{ �)>��=
�������t�k���O!���%�'�)��-��1�1q5�b&9�:�<�8I@���C�TG�"aJ�%�M���P���S���V��Z��]�<`� 
c�%�e���h���k��n���q�cdt��2w�f�y�ù|��s�����k��C������)i��w�������c��帋�����e�� ���p��n���Ɠ�����v���͗�$��Ry���͛�j!���t���ǟ����-n���£�%��
o���ǧ�h!���|��;٫��6��L�����+O��{������N`���������'e��깺�,��ob���  �  ��N=�:N=��M=��L=�7L=Q�K=\�J=�-J=�~I=�H=dH=�oG=�F=YF=�`E=رD=�D=�SC=
�B=��A=sFA=q�@=��?=4?=��>=��====Mc<=��;=�:==:=s�9=��8=�8=�Y7=ˠ6=��5=B.5=St4=��3=��2=r@2=3�1=��0=��/=�4/=[j.=��-=��,=��+=H+=�A*=5a)=`|(=�'=�&=�%=v�$=�#=q�"=�!=� =M}=Z=�-=��=H�=p=�=7�=�W=
�=�j=V�=�X=!�=4%=�
=��=!=�d=*�=[�=� =�|�<���<��<uN�<ހ�<���<_��<���<��<�	�<\�<��<�<=�< �<��<�<��<���<W�<i�<�ѩ<X��<��<���<���<~l�<�R�<H8�<��<l�<E�<5�y<�fq<R8i<ia<��X<Z�P<G�H<�@<�z8<7g0<�U(<VE <6<�'< <� <C�;���;+��;9�;���;�;"0�;�e�;�\a;$B; �";];��:6��:�!:��$9GŜ��
E� X��:�׺P��Q'%��KA��	]�~Yx�����~���ۦ��DD��ǖ��F�Ȼ�VԻz�߻�������  �LA�w?
������r�[��J!�ۈ%�/�)��-�	�1��f5��9���<��>@���C�$G�,YJ�Y�M���P���S�\�V��Z��]�7`�zc��f���h���k�ּn�p�q��nt�^=w��z���|��~���`p��|Ń�H��0l������w���d������$d���������j����T���q���ȗ�����s���ț����=p���ß�����k������0���n���ǧ��"���~���۫��9��8�������2T��Ѱ��'��	f��.������:j������+���e���  �  ��N=�9N=�M=��L=�7L=��K=�J=�.J=�I=�H=!H=oqG=��F=gF=cE=�D=�D=�UC=��B=G�A=�GA=H�@=L�?=^4?=��>=��==}==ob<=p�;=��:=_;:=��9=��8=�8=�W7=��6=��5=5,5=zr4=�3=S�2=4?2=4�1=��0=!�/=g4/=zj.=3�-=d�,=��+=�+=:C*=�b)=/~(=�'=�&=��%=i�$=�#=�"=S�!=?� =1~=�Z=M.=��=�={o=�=�=V=U�=�h=:�=�V=��=�"=,}
=m�=�=�b=0�=��=8 =Ez�< ��<��<�M�<���<_��<���<���<���<��<��<��<�<r�<W�<�<��<!�<���< �<|�<^ө<H¥<[��<x��<���<k�<�P�<�5�<��<���<V�<x�y<�]q< /i<>a<��X<�P<��H<�@<�t8<Mb0<�Q(<�B <�4<�'<7<N <��;���;+��;$��;p�;��;$B�;0x�;3�a;�8B;�#;�*;|��:F��:�":��%9������D�Z���׺د�Y6%��^A��!]�Qsx�4���hі�<����T�������Ȼ�dԻ��߻��I����# ��C�A
��-���o�C��F!���%�!�)���-���1��^5�K9�)�<��6@��C�7G�"SJ��M�p�P���S�_�V�@Z�U]��`�/c��f���h���k���n���q�wt��Ew��z���|� �����s���ȃ����n���������re���������c��i���d���g��p������n���ė�����o���ě�����l���������i������n���n��_ȧ��#��C���ޫ�<��T�������W������q��pj��{¶���n��
º�V��lh���  �  '�N==9N=M=��L=�7L=�K=_�J=//J=x�I=i�H=
"H=�rG=�F=�F=TdE=�D=�D=�VC=��B=$�A=;HA=˗@=��?=�4?=q�>=O�====�a<=��;=��:=Y::=��9=p�8=V8=NV7=C�6=2�5=�*5=@q4=Ҷ3=]�2=e>2=�1=��0=��/=D4/=�j.=x�-=��,=q�+=L +=-D*=�c)=V(=8�'=K�&=5�%=��$=�#=�"=@�!=�� =�~=[=.=��=Ǹ=o=G=K�=0U=;�=�g=��=+U=,�=.!=�{
=��=[=Ra=��=��=V =�x�<��<��<�M�<��<Ϋ�<���<��<$��<��<��<�<�!�<!�<��<��<I�<M�<���<��<��<6ԩ<�¥<��<2��<��<j�<�O�<�3�<��<w��<�߀<�y<�Wq<c)i<�`<�X<��P<��H<ȅ@<9q8<p_0<�O(<9A <�3<w'<<� <8�;��;���;��;N�;�&�;M�;���;c�a;�NB;�/#;�=;h��:Hэ:`,":�;&9�V����D��\���׺~���?%�nkA��0]�܄x�ɯ���ۖ�����_��S����Ȼ%nԻ�߻a��]���& ��E��A
�t�����n�z���C!�m�%�4�)���-�Ӌ1��Y5�19�
�<��1@�Q�C��G�/OJ��M���P���S�3�V��
Z��]��`��c�-f���h�z�k���n���q�C|t�?Kw��z��|�W�����Sv���ʃ�����o����������e��*���F��fb��j�����(f��m�������k������bm��:�����j���������h��þ������n���ȧ�G$��<���N߫�->��I���E���yZ������#��m��.Ŷ�����p��Wĺ�S��!j���  �  ��N=9N=��M=��L=�7L=�K=w�J=i/J=��I=��H=Y"H=�rG=��F=F=�dE=��D=mD=2WC=�B=o�A=zHA=��@=��?=�4?=q�>=@�==�==�a<=u�;=��:=	::=�9=�8=�8=�U7=��6=��5=�*5=�p4={�3=�2=>2=[1=V�0=��/=94/=�j.=��-=��,=��+=� +=yD*==d)=�(=��'=��&=��%=�$=w�#=i�"=��!=9� =�~=8[=�.=��=��=�n==�=�T=��=?g=e�=�T=��=� ={
=n�=�=�`=��=9�= =Wx�<���<��<�M�<#��<��<���<���<���<!�<��<��<w"�<�!�<��<k�<�<��<b��<
�<1�<lԩ<�¥<���<��<Ƃ�<�i�<
O�<E3�<!�<���<�ހ<G�y<�Uq<'i<]�`<^�X< �P<�H<w�@<�o8<X^0<�N(<�@ <�3<�'<d<> <<�;�;��;��;��;z*�;�P�;r��;�a;uVB;�5#;1C; �:dڍ:~;":U&9NL��:�D�V^���׺��&D%��pA�d5]��x�粉��ޖ��ţ�_c�� �����Ȼ@qԻ��߻��������& �8F�BB
�������n����}B!�U%���)�\�-��1��W5��9�[�<��/@���C�� G��MJ�ыM���P�$�S� �V��
Z��]�'`��c�#	f��h���k�S�n�(�q��}t�Mw��z�#�|���p ��w���˃�����p������f��/���,��Eb���������e��Ҽ������j��6������l��_������>j��q��� ��Jh����������n���ȧ�|$�������߫��>��睮�����B[��h�����/n��1ƶ����\q��ź�����j���  �  '�N==9N=M=��L=�7L=�K=_�J=//J=x�I=i�H=
"H=�rG=�F=�F=TdE=�D=�D=�VC=��B=$�A=;HA=˗@=��?=�4?=q�>=O�====�a<=��;=��:=Y::=��9=p�8=V8=NV7=C�6=2�5=�*5=@q4=Ҷ3=]�2=e>2=�1=��0=��/=D4/=�j.=x�-=��,=q�+=L +=-D*=�c)=V(=8�'=K�&=5�%=��$=�#=�"=@�!=�� =�~=[=�.=��=ɸ=o=J=O�=5U=@�=�g=��=4U=5�=9!=�{
=��=i=aa=�=��=h = y�<0��<��<�M�<2��<��<���<��<<��<��<�<$�<�!�<!�<��<��<=�<=�<���<l�<��<ԩ<�¥<a��<��<備<�i�<|O�<�3�<��<e��<�߀<܉y<�Wq<c)i<��`<�X<ùP<˝H<�@<jq8<�_0<�O(<vA <4<�'<Q< <��;�;H �;A�;��;�&�;!M�;���;0�a;qNB;n/#;�<;���:ύ:d(":�*&9�_����D�p_��a�׺����@%��lA��1]���x�J����ۖ�����_������A�ȻnnԻC�߻��껍���"& ��E�B
�������n�����C!�r�%�8�)���-�Ջ1��Y5�39��<��1@�R�C��G�/OJ��M���P���S�3�V��
Z��]��`��c�-f���h�z�k���n���q�C|t�?Kw��z��|�W�����Sv���ʃ�����o����������e��*���F��fb��j�����(f��m�������k������bm��:�����j���������h��þ������n���ȧ�G$��<���N߫�->��I���E���yZ������#��m��.Ŷ�����p��Wĺ�S��!j���  �  ��N=�9N=�M=��L=�7L=��K=�J=�.J=�I=�H=!H=oqG=��F=gF=cE=�D=�D=�UC=��B=G�A=�GA=H�@=L�?=^4?=��>=��==}==ob<=p�;=��:=_;:=��9=��8=�8=�W7=��6=��5=5,5=zr4=�3=S�2=4?2=4�1=��0=!�/=g4/=zj.=3�-=d�,=��+=�+=:C*=�b)=/~(=�'=�&=��%=i�$=�#=�"=T�!=@� =3~=�Z=O.=��=�=�o=�=�=(V=_�=�h=I�=�V=��=�"=C}
=��=�=�b=O�=��=Z =�z�<f��<��<;N�<:��<���<���<��<���<��<��<��<(�<v�<Q�<��<��<�<���<��<J�<'ө<¥<��<=��<]��<�j�<�P�<�5�<��<���<<�<T�y<x]q< /i<Oa<��X<D�P<�H<o�@<Uu8<�b0<SR(<=C <E5<
(<�<� <|�;� �;���;���;��;9�;>B�;$x�;πa;�7B;�#;�);{��:ѳ�:��!:&�%9t���@E��^��ޮ׺<���8%�aA��#]�gux�.���PҖ�����U�������ȻCeԻ�߻|�껦����# �D�"A
�+�A��	p�Q��F!���%�)�)��-���1��^5�N9�+�<��6@��C�8G�#SJ��M�q�P���S�_�V�@Z�U]��`�/c��f���h���k���n���q�wt��Ew��z���|� �����s���ȃ����n���������re���������c��i���d���g��p������n���ė�����o���ě�����l���������i������n���n��_ȧ��#��C���ޫ�<��T�������W������q��pj��{¶���n��
º�V��lh���  �  ��N=�:N=��M=��L=�7L=Q�K=\�J=�-J=�~I=�H=dH=�oG=�F=YF=�`E=رD=�D=�SC=
�B=��A=sFA=q�@=��?=4?=��>=��====Mc<=��;=�:==:=s�9=��8=�8=�Y7=ˠ6=��5=B.5=Rt4=��3=��2=r@2=3�1=��0=��/=�4/=[j.=��-=��,=��+=H+=�A*=5a)=`|(=�'=�&=�%=w�$=�#=r�"=�!=� =O}=Z=�-=��=N�=p=�=A�=�W=�=�j=j�=Y=;�=Q%=�
=�=H=�d=V�=��=� =�|�<C��<
�<�N�<<��<��<���<6��<O��<�	�<��<
�<�<B�<�<��<�
�<y�<��<�<"�<�ѩ<��<���<e��<2��</l�<�R�<8�<��<<�<�<�y<xfq<R8i<�a<��X<��P<��H<��@<X{8<�g0<8V(<�E <�6<P(<�<Z <l�;���;��;��;s��;u�;H0�;�e�;M\a;*B;��";�;���:T��:,�!:X�$9gޜ��E��^���׺����*%�OA�]�p\x� �����
���XE������%�Ȼ}WԻ'�߻o�����V  �|A��?
�����r�n��.J!��%�:�)��-��1��f5��9���<��>@���C�&G�-YJ�[�M���P���S�]�V��Z��]�7`�zc��f���h���k�ּn�p�q��nt�^=w��z���|��~���`p��|Ń�H��0l������w���d������$d���������j����T���q���ȗ�����s���ț����=p���ß�����k������0���n���ǧ��"���~���۫��9��8�������2T��Ѱ��'��	f��.������:j������+���e���  �  G�N=�;N=H�M=@�L=y7L=�K=��J=�,J=}I==�H=<H=<mG=[�F=�F=Q^E=/�D=W D=�QC=�B=!�A=�DA=Y�@=��?=�3?=|�>=3�==�==bd<=�;=��:=?:=Ά9=D�8={8=�\7=��6=h�5=�05=�v4=ݻ3=��2=B2=v�1=��0="�/=�4/=-j.=5�-=��,=��+=�+=�?*=�^)=�y(=��'=o�&=^�%=�$=��#=E�"=�!=�� =|=OY=�-=��=��=�p=�=��=�Y=O�=}m=?�=\=`�=�(=�
=(�=X"=�g=�=��=� =��<���<��<�O�<:��<��<��<���<��<��<�<�<��<��<��<��<��<���<h��<��<\ݭ<fϩ<���<-��<���<2��<�m�<?U�<F;�<� �<��<M�<�y<rq<sDi<Ja<t�X<��P<ϴH<x�@<��8<Dn0<[(<]I <l8<u(<H<: <��;J��;���;�ٿ;��;G��;��;7N�;�,a;2�A;��";��;�U�:&I�:�N!:��#9�=��2E�_��٘׺Μ�+%��7A�E�\��:x�7������u���0��T���A�Ȼ�DԻ��߻d�껰���� �d>��=
������t�����O!���%�4�)��-�
�1�8q5�h&9�?�<�<I@���C�WG�$aJ�&�M���P���S���V��Z��]�<`�!
c�&�e���h���k��n���q�cdt��2w�f�y�ù|��s�����k��C������)i��w�������c��帋�����e�� ���p��n���Ɠ�����v���͗�$��Ry���͛�j!���t���ǟ����-n���£�%��
o���ǧ�h!���|��;٫��6��L�����+O��{������N`���������'e��깺�,��ob���  �  ��N=�<N=��M=��L=S7L=I�K=��J=+J=;{I=�H=�H=pjG=X�F=�
F="[E=�D=^�C=�NC=|�B=�A=>CA=��@=�?==3?=s�>=��==�==�e<=��;=��:=xA:=��9=4�8=�8=�_7=�6=��5=�35=�y4=_�3=�3=�C2=�1=��0=��/=�4/=�i.=~�-=��,=�+=�+=�=*=k\)=#w(=��'=P�&=A�%=�$=�#=±"=צ!=�� =�z=KX=-=e�=�=�q=5=��=�[=��=ep=�=�_=�=X,=ˆ
=��=�%=	k=Щ=Z�=� =���<,��<@�<RP�<���<��<���<���<P��<[�<�	�<J�<��<l�<"�<=�<���<]��<��<y�<�٭<�̩<��<m��<Ț�<H��<�o�<$X�<?�<E%�<$�<7�<��y<�q<2Ri<(a<�Y<B�P<\�H<Ĥ@<�8<wu0<�`(<M <X:<p(<N<\ <���;i��;A��;SĿ;�ȯ;2۟;p��;2�;��`;/�A;Y�";C�;��:�:�� :})"96���qPE�\`���׺2���%�<A�?�\�<x��p��ɗ��J{�����:k��osȻ�/Ի��߻���'���� ��:�<
�q�����w����/V!���%�»)���-���1��}5�K39��<��U@�5�C�� G��jJ��M�v�P��S��W�cZ�%]�,`�Gc���e���h���k�=�n���q�^Xt��%w�f�y�Ĭ|�g����%f��r�������e��빇�3��c��ݸ�����Kg��¿�����-r��~˓�c$���|��ԗ�b*������ӛ�'���y��̟�d��&q���ģ�m��so��ǧ� ���z��:֫��2�����쯼rI��P���7 ���Y��4���J	��b_�������	��~^���  �  l�N=�=N=��M=��L=7L=��K=c�J=�)J=7yI=��H=�H=[gG=�F=.F=�WE=��D="�C=�KC=ʝB=��A=OAA=}�@=�?=�2?=S�>=��==s==�f<=a�;=�:=�C:=]�9=L�8=�8=Oc7=Z�6=�5=%75=�|4=�3==3=�E2=[�1=��0=>�/=�4/=|i.=��-=R�,=T�+=�+=;*=�Y)=t(=G�'=��&=�%=��$=޲#=��"=j�!=�� =y=,W=d,=8�=d�=�r=� =S�=�]=��=~s=��=Hc=��=W0=̊
=��=})=yn=�=�=3 =(��<���<��<�P�<���<���<���<v��<��<N��<��<��<��<~�<8�<u��<i��<g�<B�<��<B֭<"ʩ<@��<~��<ߚ�<T��<r�<#[�<
C�<*�<��<��<��y<�q<�`i<�6a<Y<��P<��H<��@<E�8<�|0<Xf(<�P <<<(<�< <���;���;��;٬�;���;���;��;��;�`;�vA;�c";��;��:봌:Z :g� 9|A���uE��c��׺Ӏ���$���@�M�\�\�w�QZ��0���a�������Q��U[Ȼ=Ի��߻���-���@ �7�[:
�x�����{����{]!���%��)�y�-���1��5��@9���<��b@��C��,G�uJ���M���P���S�xW�7Z��]�K`�Xc� �e�(�h���k���n��xq��Kt�#w���y��|��Y����]`��\���#��Ob��?���r��Xb���������7i��������v���Г�Z*�� ����ڗ�71��c���Xڛ�N-��W���П��"��zt��ǣ����
p���Ƨ����Lx��ӫ��.��􊮼K篼_C��͞��T����R��P������EY��������aZ���  �  ��N=�>N=[�M= �L=�6L=��K=*�J=�'J=#wI=)�H=$H=JdG=ʳF=�F=ATE=M�D=��C=�HC=�B=M�A=W?A=��@=��?=2?=(�>=<�==4==h<=�;="�:=sF:=1�9=n�8=>8=�f7=ĭ6=]�5=^:5=�4=��3=�3=�G2=Ɇ1=��0=��/=5/=i.=̙-=��,=��+=n+=�8*=�V)=�p(=��'=��&=��%=r�$=ү#=*�"=��!=�� =vw=�U=�+=�=��=Rs=�!=�=0`=H�=�v=]�=�f=��=F4=��
=��=1-=�q=�=��=n =���<W��<v�<�Q�<2��<��<&��<��<���<-��<(��<��<�<z �<#��<���<��<d�<��<Rܱ<�ҭ<4ǩ<N��<���<嚝<S��<�s�<^�<�F�<�.�<V�<���<�y<"�q<ioi<2Ea<Y<��P<��H<T�@<Q�8<:�0<�k(<2T <�=<�'<k<���;���;���;y��;��;5��;s��;���;}�;�{`;�;A;%,";TO;@M�:Yf�:�:�9)̞���E�lg��#t׺�s�L�$���@���\���w�dC���f��_H��:䯻y8��CȻ�Ի�w߻���`��� ��3��8
������|����d!���%���)�Q�-�I�1���5��N9���<��p@���C��8G��J��M� �P���S�W
W�Z�]�k`���b���e���h�շk�Q�n��lq��>t��
w���y�e�|�wL�j���Z��V�������^�������
���a��=������[k���ŏ�p ��o{��1֓�[0�������ᗼ#8��L�������y3������՟��&���w���ɣ�v���p��UƧ����;v��Ы��*��B����᯼M=��R�����L������8���"S����������eV���  �  m�N=�?N=�M=�L=�6L=#�K=��J=R&J=%uI=��H=�H=daG=��F=~ F=QE=�D=��C=�EC=��B=�A=q=A=z�@=��?=d1?=�>=y�==�==4i<=��;=�:=�H:=Ñ9=F�8=G"8=�i7=��6=r�5=M=5=@�4=�3=�3=RI2=�1=s�0=9�/=�4/=�h.=�-=��,=��+=Y+=$6*= T)=n(=ڃ'=m�&=e�%=X�$=�#=��"=��!=�� =�u=�T=�*=��=ۺ=t=�"=��=4b=��=]y=u�=]j=]�=�7=g�
=�=�0=�t=��=�=n =ɍ�<���<��<�Q�<��<���<���<���<���<\��<���<���<���<���<|��<��<��<��<�ߵ<�ױ<�έ<pĩ<j��<���<Ś�<2��<�u�<�`�<qJ�<;3�<n�<}�<��y<E�q<�|i<�Ra<+Y<Q<��H<�@<�8<�0<{p(<@W <�><�&<�<���;��;H��;��;�~�;\{�;r��;���;@�;QB`;UA;��!;r;���:5�:�]:>�9�T��'�E�yl���j׺�g�q�$�c�@��i\��w��.��~P���0��E̯�>!���,Ȼ��ӻ�e߻E���t��] ��0�]7
�H����^��0��k!�m�%���)���-�S�1�a�5�\9���<�m}@���C��CG�o�J���M��P���S�"W�Z�]��	`���b���e�`�h�֯k�΋n�dbq�;3t���v�3�y���|�K@�����rU������
���[��q���n	��a���������qm���ȏ�$$�����=ۓ�6������ 藼�>��ʓ��C盼S9��a����ڟ��*��{��̣���`q��5Ƨ�~��St��Oͫ�['�������ܯ��7��\���k쳼�E��U���7����M�����������R���  �  ��N=�@N=Y�M=2�L=66L=u�K=��J=�$J=rsI=��H=.H=�^G=��F=��E=&NE=W�D=(�C=CC==�B=�A=�;A=&�@=��?=�0?=��>=��==\==j<=ϵ;=� ;=�J:=��9=��8=�$8=�l7=��6=�5=�?5=��4=%�3=L
3=�J2=!�1=#�0=��/=�4/==h.='�-=��,=d�+=�+=
4*=�Q)=pk(=2�'=��&=��%=��$=e�#=1�"=��!=� =}t=�S=W*=��=�=�t=�#=��=�c=��=�{="�=<m=i�=;=z�
='�=l3=�w=�=#�= =c��<T��<��<R�<�<C��<���<���<��<��<���<F��<*��<��<���<���<v�<��<v۵<'Ա<�˭<©<���<���<���<Ɖ�<)w�<�b�<oM�<�6�<��<i�<1�y<��q<:�i<^a<6Y<uQ<5�H<?�@<r�8<M�0<mt(<�Y <v?<�%<L<���;���;8��;~�;�j�;�e�;@p�;���;�~;}`;`�@;+�!;i�;��:�ڋ:�:�>9]Ο���E��r���d׺'^��$�Ǵ@�@O\� ~w����;=�����M���2���Ȼ�ӻSV߻@��sj��� ��.��6
������ǆ��Gr!�ֹ%�8�)�@�-���1�P�5�jg9�M=�\�@�v�C�yMG�(�J�!�M�T�P��T�sW��Z��]��`��b���e���h��k�уn�4Yq�Q)t��v���y�
z|��5������P��٩�����1Y������]���`��񹋼��;o��ˏ�\'�������ߓ��:��󔖼v헼UD��T����웼x>������ޟ�J.���}��.Σ�w��r�� Ƨ�����r��˫�`$��`~���د�3��L���糼`@�������H��N��������O���  �  y�N=mAN=��M=9�L=�5L=�K=)�J=�#J=rI=9�H=lH=�\G=�F=��E=�KE=4�D=�C=�AC=~�B=��A=�:A=�@=�?=M0?=��>=��==�==�j<=��;=�;=L:=��9=��8=�&8=�n7=��6=�5=�A5=S�4=��3=�3=�K2=�1=��0=��/=�4/=�g.=��-=��,=<�+=0+=`2*=�O)=wi(='=��&=��%=��$=p�#=v�"=��!=�� =is=S=�)=O�=!�=�t=�$=��=.e=O�=�}=&�=eo=��=f==ۗ
=s�=�5=�y=ض=��=Y =[��<���<z�<:R�<�~�<#��<۽�<���<G��<���<-��<0��<���<���<b��<*��<e�<޹< ص<<ѱ<Jɭ<%��<a��<模<���<A��<Rx�<�d�<�O�<�9�<#�<�<7�y< �q<�i<�fa<S>Y<=Q<F�H<|�@<��8<d�0<xw(<6[ <�?<7%<=<0��;���;*��;�p�;�[�;�T�;^�;�z�;+X;t�_;�@;�!;�;�r�:7��:��:�69>/���F�]w��_׺iV���$�Σ@��:\��ew�`���.��-�����������Ȼ��ӻ�J߻>{껂b���  ��,��5
�'���������w!���%��)���-��1��5�>p9�#=��@���C��TG���J���M�$�P��T�W��Z�]�$`��b���e���h�ʣk��}n�KRq��!t��v�N�y��q|��-�"󀼘M��馃�>���>W��!���|��r`��;������p��͏��)������*㓼�>������񗼺H��������`B������
⟼ 1��4����ϣ�� ���r��Ƨ�/���q��\ɫ�"���{���կ��/��{���㳼:<��锶�C�5E��������cM���  �  �N=�AN=�M=5�L=�5L=��K=��J=&#J=BqI=9�H=DH=�[G=��F=;�E=�JE=ۛD=��C=`@C=^�B=��A=�9A=|�@=��?= 0?=c�>=��====-k<=S�;=�;=M:=��9=��8=(8=�o7=��6=X�5=�B5=i�4=��3=w3=rL2=h�1=��0=��/=�4/=�g.= �-= �,=��+=H+=W1*=�N)=3h(=�}'=:�&=3�%=W�$=1�#=M�"=��!=�� =�r=�R=})=)�= �=(u= %=��=�e=G�=�~=e�=�p="�=�>=N�
=��=�6=�z=��=��= =w��<���<��<1R�<(~�<g��<˼�<��<r��<���<���<���<)��<���<���<l��<��<�۹<�յ<_ϱ<�ǭ<���<���<d��<d��<���<�x�<�e�<Q�<�;�<+%�<v�<h�y<`�q<��i<la<�CY<"Q<��H<q�@<ĵ8<Ԗ0<%y(<I\ <@<�$<�	<��;��;��;h�;R�;J�;�R�;�n�;�@;��_;��@;c�!;{�;�N�:g��:�j:Q�9Vh��F��y��6[׺*R���$��@�@-\��Vw����U%�����Ӟ������jȻ��ӻC߻�t��]�������+�5
������E��6�*z!�Z�%�b�)�f�-�H�1�O�5��u9��=�R�@��D��YG�J�J���M�9�P��	T��W��Z��]��`���b���e�L�h���k��yn�Nq�t��v�5�y��l|�)������K���������V��S������H`����������q��OΏ�|+������c哼&A������m���cK��[������D��𔞼䟼�2�������У�X!��s��4Ƨ�����p��Sȫ�� ���y���ӯ�H-������೼�9��m����근�B�����D�
L���  �  ��N=dKN=P�M=A�L=<AL=*�K=<�J=�.J=�|I=R�H=JH=�fG=,�F=�F=XE=��D=��C=�SC=��B=��A=�UA=��@=� @=�T?=�>=��==�J==�<=��;=6;=��:=��9=F9=>e8=֯7=��6=XC6=0�5=�4=�4=u`3=A�2=	�1=[%1=b0=��/=�.=�.=I4-=�_,=�+=y�*=X�)=��(=A(=�'=�+&=�8%=�@$=:C#=>?"=4!=%! =~=u�=��=Rx=S4=^�=��=�&=�=�<=y�=,*=L�=s�=�G=��	=e�=g=jS=ڄ=�� =��<���<g�<�E�<;e�<�{�<"��<^��<���<���<���<�}�<r�<Re�<�X�<NL�< @�<=4�<x(�<`�<��<��<+�<��<^͝<̷�<��<���<�k�<?O�<2�<��<��y<��q<�yi<CAa<Y<4�P<c�H<�u@<�G8<�0<��'<K�<��<�l<v@<�(�;���;+��;/5�;e��;���;���;��;�<y;}�Y;�:;s�;v_�:���:��x:|��9���7����<h�S��E��|���R.�W�J�{sf��Co����������E]��������ͻF�ٻC��z�e��)��,��2�B�[���w�7���V$��(�S�,���0��4��^8��<���?���B�UF���I�P�L���O���R���U�b�X�<�[��^�Q�a�ld�!Dg�?j�(�l���o�Izr�B<u���w�$�z��f}�����a�������m^������a���Y���������|_��˹����[q���͒��)������ޖ�,5������ۚ�b+���x��Ğ�W��X��㡢��주�8��r���G֧�	(���{���Ы��'��'��9ׯ�p/������d߳��6������䷼:�����滼�<���  �  ��N=CKN=>�M=B�L=OAL=T�K=|�J=�.J=�|I=��H=�H=hgG=��F=AF=�XE=��D=��C=�TC=�B= B=VA=ѫ@=� @=U?=�>=��==�J==�<=H�;=�5;=T�:=P�9=�9=�d8=1�7=>�6=�B6=��5=��4=�4=`3=�2=��1=C%1=b0=��/=,�.= .=�4-=I`,=p�+=�*=��)=0�(=�(=�'=P,&=^9%=^A$=�C#=�?"=�4!=n! =�=��=��=Lx=?4=:�=A�=P&=��=e<=�=�)=��=��=G=G�	=��=�=�R=a�=�� ={��<Q��<+�<�E�<?e�<�{�<��<��<d��<ۏ�<���<�~�<Ds�<�f�<9Z�<�M�<_A�<n5�<�)�<Z�<j�<V�<��<0�<�͝<̷�<<C��<�j�<�N�<I1�<��<��y<|�q<�vi<�>a<�Y<��P<a�H<�s@<EF8< 0<��'<��<d�<�l<�@<O*�;���;9��;�8�;���;�Ƭ;`��;癌;�Iy;:�Y;g:;�;,s�:�Ĺ:f
y:��9(��7v��0h�D�����=���U.��J��wf����r������)���.b��������ͻ��ٻ�E�L}�g����
-��2������v�.���U$��(�v�,�R�0���4�e\8��<���?�	�B��RF�c�I�t�L���O���R��U���X���[��^�^�a�ald��Dg�yj���l�#�o�$|r��>u��w��z�3i}����c������_��E������Z���������B_��Q�������p���̒��(�������ܖ��3�������ښ�<*��{w��Þ�k��?W��O���*주c8��J���@֧�)(��|��yѫ�F(�����د�i0�������೼�7��ӎ��!巼;��ܐ���滼>=���  �  ��N=�JN=��M=F�L=�AL=ёK=;�J=�/J=~I=�H=XH=iG=��F=	F=�ZE=p�D=OD=,VC=��B=gB=8WA=��@=�@=uU?=H�>=��==9J==o�<=��;=�4;="�:=��9=19=c8=��7=��6=,A6=�5=1�4=C4=_3= �2=/�1=�$1=�a0=Л/=z�.=�.=Q5-=Ga,=��+=L�*=t�)=��(=�(=j'=.&=;%=C$=ME#=A"=�5!=\" =i= �=ޱ=Ex=�3=��=t�=K%=[�=�:=5�=�'=��=��=E=^�	=��==aQ=�=�� =ԧ�<��<}�<sE�<�e�<�|�<��<Γ�<���<���<��<3��<�v�<{j�<�]�<=Q�<�D�<�8�<x,�<��<��<&�<��<��<�͝<���<=��<
��<Pi�<WL�<�.�<��<��y<��q<�oi<�7a<�Y<6�P<F�H<�n@<B8<�0<G�'<�<�<im<B<�/�;���;���;�C�;`�;լ;´�;]��;;iy; �Y;�1:;��;��:c��:Ocy:�i�9��7��dh����Y��{���].���J��f������}�� ���=���tn��~���r�ͻj�ٻvO�+��m���V.�_3�l����Wt����YQ$��(�ï,��0���4�5U8�^�;�l�?���B��KF��I�øL���O�n�R���U��X���[�c�^��a��md�]Gg��j���l�7�o��r��Du�dx���z��o}����+f������>��a��ȳ������Z��˯��R��r^���������{n��Rʒ��%��O���aٖ�S0�������֚��&��t��򿞼�
���T��f����꣼Y7������(֧��(���|���ҫ�*��!����گ�h3�������㳼V;�����U跼>������黼?���  �  ��N=JN=��M=L�L=�AL=��K=R�J=`1J=�I=C�H=�H=�kG=f�F=�F=�]E=b�D= D=�XC=�B=uB=�XA=$�@=�@=!V?=��>=��==�I==��<=S�;=,3;=B:=��9=�9=g`8=Ȫ7=��6=j>6=��5=��4=>4=S]3=��2=.�1=B$1=�a0=�/=��.=�.=�6-=�b,=��+=��*=��)=��(=v	(=['=�0&=�=%=�E$=�G#=6C"=~7!=�# =�=��=8�=4x=}3=��=/�=�#=T�=�8=��=�$=��=|�=�A=3�	=��=f= O=�=Ϭ =>��<e��<��<CE�<Cf�<2~�<*��<ɖ�<h��<
��<���<���<�|�<�p�<�c�<>W�<�J�<�=�<61�<$�<�<��<���<*�<FΝ<?��<��<��<vf�<�H�<Z*�<��<�y<�q<�ci<�+a<K�X<��P<֓H<of@<;8<'0<]�'<��<I�<Kn<�D<�7�;���;��;jU�;`�;��;^͜;Ì;�y;��Y;�d:;a;W�:|F�:f�y:�+ :���7r��u�g������� ��l.��J�[�f����F����Л��ͨ��������Tλ��ٻy^��w����T0��3������p�����J$�I�(�v�,��0���4�hI8�G�;�Qy?��B��@F��I�y�L��O���R�}�U�~�X�9�[���^���a�pd�,Kg�"j�Z�l�.�o��r��Nu�]x���z��z}�P��k��1�����Bd��J�������[���������)]�������k��Nƒ�:!��K{���Ӗ�r*���~��	њ�� ���n��!���R��;Q��L���W裼�5��鄦�֧�+)��F~���ԫ��,�������ޯ�$8�����Y鳼�@���������B��̗���컼B���  �  ,�N=IN=�M=8�L=`BL=��K=��J=<3J=/�I= �H=�H=oG=��F=�F=taE=�D=�D=\C=��B=B=)[A=�@=�@=�V?=�>=��==%I==q�<=��;=1;=�|:=��9=�9=�\8=;�7=;�6=�:6=8�5=��4=�4=[3=�2=��1=^#1=<a0=�/=��.=�.=8-=�d,=�+=d�*=�)= �(=
(=#'=�4&=�A%=I$=�J#=�E"=�9!=�% =�=��=��=x=�2=��=v�=b!=��=\5=�=� =��=V�=�==-�	=�=�=�K=T~=�� =���<���<"�<�D�<g�< ��<���<���<3��<Ɯ�<.��<���<��<Px�<�k�<�^�<�Q�<�D�<77�<+)�<c�<+
�<e��<��<�Ν<���<I��<>��<�b�<�C�<�$�< �<$�y<;�q<�Ti<�a<��X<εP<-�H<k[@<�18<�	0<�'<��<�<_o<`H<pB�;v��;���;l�;�3�;	�;R�;��;`�y;{)Z;�:;�T;�u�:���:C�z:�� :���7���հg����2�麻���.�l�J��f��"�������電�稻����M» %λ��ٻ�r�̢�[�����V3��4���4���k���@B$�=~(���,�̘0�{x4��:8��;�j?�X�B�w2F��tI���L���O�x�R��U���X�}�[��^��a�Xsd�oPg�7)j�S�l���o�H�r��[u�Dx���z��}�-���q��'ł�9���h�������
��]��r���L���[����������f�����0���t���̖�#��Lw���ɚ�����g��ƴ��� ���L��z���w壼�3��惦�֧�.*��F����׫��0��u����䯼o>������c�H������M���6I�������F���  �  Y�N=�GN=^�M=�L=�BL=�K=J�J=O5J=ބI=�H=e#H=
sG=5�F=F=�eE=n�D=�D=�_C=e�B=	B=�]A=ر@=S@=�W?=5�>=`�==HH==�<=��;=�.;=�y:=d�9=�9=�X8=��7=��6=�66=>�5=2�4=Q4=BX3=��2=*�1=F"1=�`0=�/='�.=�.=�9-=g,=��+=��*=��)=��(=?(=Z''=�8&=�E%=M$=^N#=I"=�<!=�' =l
=��=�=�w=�1=(�=k�=�=`�=�1=ѫ=\=ƃ=f�=�8=l�	=��=�=H={=� =���<���<d�<nD�<�g�<��<��<��<���<&��<���<��<͌�<0��<�t�<�g�<Z�<7L�<�=�<//�<3�<��<���<��<�Ν<���<)��<�|�<^�<7>�<��<���<_�y<�}q<hBi<�
a<H�X<��P<pxH<EN@<�&8<<0<��'<��<��<Ap<�K<kN�;��;���;Յ�;�Q�;�)�;��;�	�;].z;�vZ;D�:;��;���:��:�g{:pb:?�8�)�oxg���2�����l�.���J��f�;��`�������޽��o'»Cλ�ڻ׊�u��}���~�7��6���v���f�����8$��r(���,�ԉ0�h4�d)8�^�;�fX?��B�"F��eI���L�L�O��R���U���X���[�y�^�ԓa�|wd��Vg��1j�%m�r�o�f�r��ku��+x���z�(�}�U$��?y��̂�]���m����������^��������Z��°������a��$���{��m��kĖ�f���n������0���_����������G��3���3⣼�1������0֧��+������p۫�u5��2���민�E��ş�������P�����[����P��&���l����J���  �  =�N=RFN=��M=��L=/CL=u�K=��J=t7J=��I=]�H=-'H=,wG=��F=�F=|jE=�D=1D=�cC=�B=FB=Q`A=�@=�@=�X?={�>= �==PG==|�<=��;=�+;=jv:=��9=�
9=�T8=m�7=Z�6=G26=�{5=H�4=�4=HU3=;�2=E�1=
!1=�_0=�/=��.=�	.=�;-=li,=��+=��*=��)=�(=�(=�+'=�=&=J%=!Q$=+R#=aL"=C?!=�) ==��=5�=�w=�0=��=�=�=�=�-=Q�=p=�~= �=�3=B�	=��=8
=D=�w=�� =��<���<`�<�C�<Bh�<���<M��<���<n��<��<w��<d��<���<���<*~�<�p�<�b�<\T�<*E�<P5�<*$�<��<���<^�<ϝ<C��<���<�x�<�X�<�7�<��<?��<2�y<�jq<�.i<(�`<]�X<�P<RhH<@@<�8<a�/<��'<��<<q<�N<�Z�;�;���;'��;tq�;�L�;�6�;�1�;��z;��Z;�>;;S�;��:���:#8|:�:�8�p߹C@g�m뮺������R�.�8K�#g��U�������(���)��^ൻiI»�cλk,ڻ<�廮�𻤧��\�_;��8�Y����{a���/$��f(�~,��y0�W4�8���;��E?���B�F��UI�}�L�X�O�[�R�\�U���X�Y�[��^�6�a�|d��]g�F;j��m�E�o�ܴr��|u��=x�J�z�a�}�9-�������ӂ�$��Is��A�1�� a�����X���X����������\��򴒼:���d��ֻ��<��;e������E���W��������wA��ʏ���ޣ��/�����|֧� -��f����߫��:��e���I��M��z�������Y��'������X��s�������P���  �   �N=�DN=��M=��L=sCL=X�K=a�J=�9J==�I=��H=�*H=A{G=�F=BF=oE=��D=�D=�gC=��B=WB=�bA=�@="@=hY?=��>=��===F==Œ<=H�;=);=
s:=̼9=j9=P8=Ǚ7=��6=�-6=�w5=B�4=5
4=6R3=��2=P�1=�1=@_0=�/=/�.=�
.=<=-=�k,=i�+=N�*=O�)=D�(=(=e0'=�A&=xN%=<U$=�U#=�O"=�A!=, =�=n�=k�=w=�/=��=��=�=T�=m)=��=�=`y=��=-.=
}	=��=�=�?=t=� =G��<;��<+�<�B�<�h�<���<t��<��<���<ǰ�< ��<��<
��<���<���<�y�<rk�<?\�<1L�<?;�<)�<x�<���<�<�Ν<ܲ�<ޔ�<�t�<�S�<�1�<��<��<�y<*Wq<i<h�`<i�X<��P<�WH<�1@<�8<��/<�'<+�<[�<aq<R<f�;4)�;���;��;���;�o�;�\�;�Y�;��z;�[;�;;�/;��:�:6}:��:�8��޹�g�6鮺��d���.�o@K��Kg��q��[����I��wL������k»߃λ�Jڻg�廲��Y����!�4@�	;���:���\�����%$��Z(��q,�ej0��E4�8�!�;�$3?���B���E�rFI��zL�ÞO�ܴR�<�U�$�X��[���^���a�4�d��eg�Ej��m�k�o���r���u��Ox��
{��}�?6�����fۂ��*��y���Ɔ����Ic�����H��W��q������W��񮒼-��]��7���7��	\��g���q���mO������M퟼<��f����ۣ��-��_���ק��.��k����㫼�?��Ĝ�������U��.����� c��f�������`��󲺼>��hU���  �  �N=3CN=��M=�L=�CL=�K=��J=s;J=��I=��H=0.H=�~G=�F=y!F=asE=��D=�D=�kC=�B=/B="eA=��@=K	@=Z?=��>=�==(E==�<=�;=<&;=�o:=3�9=n9=�K8=g�7=P�6=_)6=�s5=u�4=�4=?O3=C�2=q�1=I1=�^0=��/=��.=�.=�>-=�m,=��+=\�*=��)=)=(=�4'=,F&=vR%=Y$=3Y#=�R"=dD!=�- =�='�=��=xv=�.=�=r~=�=�=�%=^�=�=qt=��=))=x	=�=R=<=�p=3� =���<���<�<�A�<i�<1��<+��<˫�<&��<���<'��<ԯ�<`��<���<3��<W��<^s�<nc�<�R�<�@�<l-�<��<�<W�<uΝ<o��<��<q�<�N�<Y+�<��<��<��y<�Dq<�i<��`<S�X<�pP<}HH<�#@<�8<#�/<��'<v�<��<Vq<�T<�o�;48�;��;���;��;돭;��;~~�;�{;1d[;��;;�r;��:�}�:ʺ}:K:�8t&޹��f��论@�麥���.��fK�&xg�ً������i��_m���$��Ԍ»<�λ�gڻ��������^(�'E�b=��I���X�����$�,P(�e,�P\0�G64���7���;��!?� �B�%�E�V8I�
nL��O�e�R��U��X�D�[�?�^�{�a�m�d��lg��Nj�r+m��p���r��u�ax�q{���}��>������₼K1���~��Tˆ�)���e��4���c���U��8�������LS��]��������U��>�������vS��讀�X����G��Ǘ��M矼7������٣�,����ק��0��e����竼E��آ��� ���]����������k��!¶�R���h��񹺼c
���Z���  �  ?�N=�AN=��M=��L=�CL=��K=��J=�<J=��I=��H=1H=*�G=n�F=%F=�vE=<�D=�D=�nC=��B=�B=gA=�@=D
@=�Z?=��>=|�==D==��<=,�;=�#;=m:=�9=��8=*H8=��7=��6=�%6=�o5=&�4=�4=�L3=�2=��1=1=�]0=f�/=��.=�.=�?-=ho,=!�+=��*=��)=H)={!(=8'=�I&=�U%=.\$=\#=U"=qF!=�/ =�=��=��= v=�-=��=m|=t=�=+"=��=�	=Ap=k�=�$=�s	=�=��=�8=�m=�� =Ë�<���<�<�@�<<i�<j��<p��<!��<u��<,��<7��<g��<i��<���<|��<e��<z�<�i�<	X�<7E�<1�<H�<��<��<Ν<گ�<���<�m�<J�<�%�<��<�݀<�vy<=5q<_�h<��`<�X<JbP<�:H<�@<|�7<��/<W�'<֥<��<?q<�V<Qx�;�D�;|�;m��;�Ž;W��;!��;���;�\{;�[;<;d�;4��:ټ:�U~:}�:� 8�ݹ�f�쮺���&�/�@�K�B�g�6���P6����������tA��è»9�λπڻQ�廁������.��I�@������@U�]���$�8G(�nZ,�P0�)4���7�{�;�|?�(�B���E�,I�pcL��O�<�R�ӳU�ָX��[��^�G�a�&�d�6sg��Vj��5m�Rp���r�#�u��ox��+{���}�
F�����&邼 7������Qφ�0���g��d������$U��e��������O������@����O����������NL��֞����rA��𑞼L⟼�2��\����֣��*������xا�V2�����(뫼}I��-������qd������&���s���ɶ�}���o��2������B_���  �  ��N=�@N=��M=[�L=�CL=�K=��J=$>J=1�I=��H=13H=��G=�F=�'F=�yE=��D=pD=qC=��B=NB=�hA=�@=�
@=�Z?=��>=
�==RC=={�<=��;=";=�j:=��9=W�8=CE8=��7=�6=�"6=9m5=��4=�4=�J3=k�2=e�1=1=]0=(�/=��.=".=�@-=�p,=��+=��*=��)=�)=&$(=�:'=XL&=}X%=�^$=G^#=�V"=�G!=�0 =�=	�=��=�u=�,=X�=�z=y=��=}=��=�=�l=�=q!=�p	=��=��=6=qk=�� =���<u��<x�<4@�<5i�<;��<��<���<���<��<ƿ�<q��<��<���<$��<��<)�<4n�<\�<�H�<�3�<+�<��<A�<�͝<���<���<�j�<�F�<�!�<���<�؀<�jy<�(q<��h<O�`<��X<.WP<{0H<�@<��7<	�/<h�'<_�<��<�p<�W<\~�;)N�;3!�;���;�׽;��;��;���;��{;*�[;�@<;��;�6�:�:��~:�!:��$8S`ݹ��f�]����k4�/��K�D�g������I��s���D���SX��0�»W�λؓڻ)滋�t����3��L�-B�#�#��S�����$��@(�~R,� G0�!4���7�e~;�f?�#{B���E��"I�z[L�i�O���R��U���X�_�[���^���a���d�vxg��]j�F=m��p���r��u�|{x��7{���}��K��V����;��G����҆����qi��b�������T��$��������L��I���0���K������h��F��T���8뛼�<�������ޟ��/������.գ��)������٧��3������L��T���v���i��YƲ�!���y��|϶�3#���t���ĺ����b���  �  ��N=@N=��M=�L=�CL=O�K=��J=�>J=�I=��H=�4H=�G=��F=i)F=b{E=��D=	 D=�rC=�B=jB=[iA=ĺ@=[@=�Z?=w�>=��==�B==��<=��;=� ;=�i:=
�9=��8=zC8=�7=��6=� 6=pk5=�4= 4=gI3=Z�2=��1=t1=�\0=��/=��.=x.=TA-=kq,=��+=
�*=H�)==
)=�%(=g<'=�M&=
Z%=`$=�_#=X"=�H!=k1 ==G�=��=Iu=^,=��=�y=<=)�=�=�=�=�j=��=m=�n	=�=��=x4=�i=�� =���<���<��<�?�<Ni�<͉�<-��<#��<���<���<���<���<1��<���<���<<��<^��<q�<�^�<�J�<I5�<I�<m�<n�<;͝<ĭ�<>��<�h�<ND�<��<���<Հ<Dcy<O!q<�h<��`<{X<�OP<�)H<�@<��7<��/<"�'<1�<��<�p<�X<"��;T�;�(�;��;��;Fͭ;;č;C�{;.�[;b]<;��;Yh�:�G�::*Y:�5'8�,ݹ�f�����}>�e'/��K�D�g������V�����ƭ���e����»�λj�ڻ6�C'�����6�eO��C�������Q�/��V$�{<(�wM,�<A0��4� �7��w;��?��tB���E�0I�nVL�M�O�ƜR���U�:�X�ִ[�4�^��a�9�d��{g��aj�QBm�Mp�@�r�$�u���x��>{���}�kO��ӡ��'�I>�������Ԇ�9���j���������OT��V�������K�������H��\���1�rC�����蛼�9��׊��8ܟ�.������3ԣ�g)��{����٧��4��}����﫼:O������s���l���ɲ��$��}��Ӷ��&��x���Ǻ����e���  �  ��N=�?N=[�M=�L=�CL=b�K=�J="?J=m�I=S�H=�4H=��G=8�F=*F=|E=3�D=� D=sC=��B=�B=�iA=�@=y@=[?=t�>=��==�B==t�<=W�;=h ;=i:=}�9=�8=�B8=.�7=��6=V 6=�j5=s�4=��3=�H3=��2=D�1=71=�\0=�/=��.=�.=�A-=�q,=	�+=i�*=��)=�
)=D&(=='=�N&=�Z%=�`$=`#=vX"=6I!=�1 =C=O�=y�=3u=;,=B�=}y=�=��=O=H�==8j=*�=�=�m	=Z�=M�=�3=�i=0� =��<���<T�<�?�<Xi�<���<���<���<m��<k��<���<���<^��<]��<ѡ�<]��<q��<r�<Q_�<MK�<�5�<��<��<j�<͝<t��<���<Vh�<}C�<�<}��<�Ӏ<�`y<�q<��h<�`<�xX<|MP<�'H<�@<��7<��/<�'<��<V�<�p<IY<r��;�V�;�+�;-�;q�;�ѭ;�Ɲ;�ɍ;<�{;��[;g<;��;fw�:�T�:�%:�l:��'8-!ݹ�f�����)	�5B��+/���K��g��ā��[������{���l����»��λ�ڻ��*�C����7�LP��C������>Q�c��$�;(��K,�X?0��4���7��t;���>�prB�b�E�PI��TL��~O���R��U���X�ϴ[�Y�^�i�a��d��|g�cj�Dm�.p�~�r�{�u��x��A{���}��P�����C�1?������Ն�����j��"������;T��#���*���qJ��f�����"G��A���
B�����曼{8��󉞼u۟�S-������ӣ�A)��{����٧��4������h��O��ݯ��z��n��˲��%���~��fԶ��'��Cy��ɺ�����e���  �  ��N=@N=��M=�L=�CL=O�K=��J=�>J=�I=��H=�4H=�G=��F=i)F=b{E=��D=	 D=�rC=�B=jB=[iA=ĺ@=[@=�Z?=w�>=��==�B==��<=��;=� ;=�i:=
�9=��8=zC8=�7=��6=� 6=pk5=�4= 4=gI3=Z�2=��1=t1=�\0=��/=��.=x.=TA-=kq,=��+=
�*=H�)==
)=�%(=h<'=�M&=
Z%=`$=�_#=X"=�H!=l1 ==I�=��=Ku=a,=��=�y=B=0�=�=�=�=�j=�=|=�n	=�=��=�4=j=�� =ц�<%��<��<�?�<{i�<���<U��<G��<ս�<���<���<���<9��<���<���<1��<N��<q�<n^�<}J�<&5�<#�<E�<E�<͝<���<��<�h�<-D�<��<~��<�Ԁ<+cy<B!q<�h<Ƭ`<{X<
PP< *H<	@<��7<:�/<q�'<��<�<q<8Y<���;�T�;c)�;@�;��;�ͭ;4;.č;4�{;��[;�\<;N�;�f�:sE�:Y	:�S:&�&8(9ݹ]�f�(���$�@��(/���K���g�8����W������U���yf��]�»t�λƠڻ�滉'�����6�{O��C�������Q�8��^$��<(�|M,�@A0��4�#�7��w;��?��tB���E�1I�nVL�M�O�ƜR���U�:�X�״[�4�^��a�9�d��{g��aj�QBm�Mp�@�r�$�u���x��>{���}�kO��ӡ��'�I>�������Ԇ�9���j���������OT��V�������K�������H��\���1�rC�����蛼�9��׊��8ܟ�.������3ԣ�g)��{����٧��4��}����﫼:O������s���l���ɲ��$��}��Ӷ��&��x���Ǻ����e���  �  ��N=�@N=��M=[�L=�CL=�K=��J=$>J=1�I=��H=13H=��G=�F=�'F=�yE=��D=pD=qC=��B=NB=�hA=�@=�
@=�Z?=��>=
�==RC=={�<=��;=";=�j:=��9=W�8=CE8=��7=�6=�"6=9m5=��4=�4=�J3=k�2=e�1=1=]0='�/=��.=".=�@-=�p,=��+=��*=��)=�)=&$(=�:'=XL&=}X%=�^$=H^#=�V"=�G!=�0 =�=�=��=�u=�,=_�=�z=�=��=�=ї=�=m=�=�!=�p	= �=��=>6=�k=� =���<���<��<�@�<�i�<���<g��<��<��<C��<��<���<��<���<��<Ԏ�<
�<
n�<�[�<_H�<l3�<��<k�<��<D͝<M��<W��<zj�<ZF�<z!�<���<^؀<�jy<�(q<��h<g�`<��X<tWP<�0H<@<�7<��/< �'<��<d�<�q<�X<��;AO�;/"�;���;xؽ;���;Y��;ӵ�;��{;��[;�?<;n�;l3�:#�:��~:�:�	$8�wݹ�f�����2�麑7�+/��K�"�g�W���?K������Y���NY���» �λ��ڻ��������3�M�QB�A�<��(S�����$��@(��R,�G0�'4���7�i~;�j?�&{B���E��"I�|[L�j�O���R��U���X�_�[���^���a���d�vxg��]j�G=m��p���r��u�|{x��7{���}��K��V����;��G����҆����qi��b�������T��$��������L��I���0���K������h��F��T���8뛼�<�������ޟ��/������.գ��)������٧��3������L��T���v���i��YƲ�!���y��|϶�3#���t���ĺ����b���  �  ?�N=�AN=��M=��L=�CL=��K=��J=�<J=��I=��H=1H=*�G=n�F=%F=�vE=<�D=�D=�nC=��B=�B=gA=�@=D
@=�Z?=��>=|�==D==��<=,�;=�#;=m:=�9=��8=*H8=��7=��6=�%6=�o5=&�4=�4=�L3=�2=��1=1=�]0=f�/=��.=�.=�?-=ho,=!�+=��*=��)=H)={!(=8'=�I&=�U%=/\$=\#=U"=rF!=�/ =�=��=��=v=�-=��=z|=�=��=@"=��=�	=bp=��=%=t	=C�=��=�8=�m=�� =E��<G��<��<}A�<�i�<���<ݟ�<���<˸�<t��<o��<���<���<���<q��<I��<�y�<ci�<�W�<�D�<�0�<��<F�<��<�͝<k��<(��<;m�<�I�<�%�<L�<�݀<\vy<5q<^�h<�`<-�X<�bP<W;H<�@<0�7<��/<.�'<��<��<%r<�W<�y�;;F�;��;���;�ƽ;��;���;���;�\{;U�[;�<;��;���:~Ӽ:�H~:�:��8C�ݹ[�f��������y*�b	/�|�K�Q�g�"���8��<���C����B���»U�λˁڻ-��@�e����.��I�5@�����]U�u���$�IG(�{Z,�&P0� )4���7���;��?�,�B���E�,I�rcL��O�>�R�ԳU�׸X��[��^�G�a�&�d�6sg��Vj��5m�Rp���r�#�u��ox��+{���}�
F�����&邼 7������Qφ�0���g��d������$U��e��������O������@����O����������NL��֞����rA��𑞼L⟼�2��\����֣��*������xا�V2�����(뫼}I��-������qd������&���s���ɶ�}���o��2������B_���  �  �N=3CN=��M=�L=�CL=�K=��J=s;J=��I=��H=0.H=�~G=�F=y!F=asE=��D=�D=�kC=�B=/B="eA=��@=K	@=Z?=��>=�==(E==�<=�;=<&;=�o:=3�9=n9=�K8=g�7=P�6=_)6=�s5=u�4=�4=?O3=C�2=q�1=I1=�^0=��/=��.=�.=�>-=�m,=��+=\�*=��)=)=(=�4'=-F&=vR%=Y$=4Y#=�R"=gD!=�- =�=,�=��=�v=�.=�=�~==��=�%=|�=�=�t=��=\)=Xx	=U�=�=f<=�p=�� =[��<y��<��<zB�<�i�<���<���<C��<���<L��<l��<��<|��<���<%��<4��<'s�<$c�<MR�<D@�<�,�<"�<��<��<�͝<簙<���<�p�<(N�<�*�<��<��<7�y<�Dq<�i<��`<��X<xqP<IH<�$@<�8<�/<��'<��<�<pr<�U<�q�;:�;[�;*��;?��;Ӑ�;Z��;�~�;S{;Nc[;�;;�p;*{�:�v�:�}:j9:�8&O޹�g�v�6�����.��kK�}g�3�������k��>o��B&��[�»��λ�hڻ������i����(�pE��=�6�t���X����$�@P(�e,�]\0�Q64���7��;��!?�$�B�(�E�Y8I�nL��O�f�R��U��X�E�[�?�^�|�a�m�d��lg��Nj�r+m��p���r��u�ax�q{���}��>������₼K1���~��Tˆ�)���e��4���c���U��8�������LS��]��������U��>�������vS��讀�X����G��Ǘ��M矼7������٣�,����ק��0��e����竼E��آ��� ���]����������k��!¶�R���h��񹺼c
���Z���  �   �N=�DN=��M=��L=sCL=X�K=a�J=�9J==�I=��H=�*H=A{G=�F=BF=oE=��D=�D=�gC=��B=WB=�bA=�@="@=hY?=��>=��===F==Œ<=H�;=);=
s:=̼9=j9=P8=Ǚ7=��6=�-6=�w5=B�4=5
4=6R3=��2=P�1=�1=@_0=�/=/�.=�
.=<=-=�k,=i�+=N�*=O�)=D�(=(=e0'=�A&=xN%==U$=�U#=�O"=�A!=, =�=s�=s�=w=�/=��=Ȁ=�=m�=�)=ע=�=�y=��=g.=I}	=�=�=?@=et=]� =���<���<��<�C�<ni�<T��<	��<i��<p��<)��<m��<$��<*��<��<r��<�y�<5k�<�[�<�K�<�:�<�(�<��<^��<��</Ν<E��<M��<pt�<DS�<1�<��<��<��y<�Vq<i<��`<İX<��P<�XH<t2@<�8<��/<<�'<_�<��<�r<8S<Yh�;R+�;���;���;�;�p�;w]�;�Y�;��z;�[;[�;;%-;���:Y�:��|:��:�8�޹C+g�S���K��x���.�8FK�;Qg�ft�����L���N��f���m»d�λ2Lڻ��廷��:����!��@�N;���j���\����%$��Z(��q,�tj0�F4�8�)�;�+3?���B���E�uFI��zL�ŞO�ݴR�>�U�%�X��[���^��a�4�d��eg�Ej��m�k�o���r���u��Ox��
{��}�?6�����fۂ��*��y���Ɔ����Ic�����H��W��q������W��񮒼-��]��7���7��	\��g���q���mO������M퟼<��f����ۣ��-��_���ק��.��k����㫼�?��Ĝ�������U��.����� c��f�������`��󲺼>��hU���  �  =�N=RFN=��M=��L=/CL=u�K=��J=t7J=��I=]�H=-'H=,wG=��F=�F=|jE=�D=1D=�cC=�B=FB=Q`A=�@=�@=�X?={�>= �==PG==|�<=��;=�+;=jv:=��9=�
9=�T8=m�7=Z�6=G26=�{5=H�4=�4=HU3=;�2=E�1=
!1=�_0=�/=��.=�	.=�;-=li,=��+=��*=��)=�(=�(=�+'=�=&=J%="Q$=,R#=cL"=E?!=* ==��=<�=�w=�0=��=/�=�=��=�-=u�=�=�~=U�=�3=��	=��=�
=aD=�w=U� =͙�<l��<�<�D�<�h�<���<��<��<��<t��<Ǧ�<���<��<���<~�<�p�<�b�<T�<�D�<�4�<�#�<H�<���<��<dΝ<���<��<fx�<}X�<�7�<.�<��<Ѩy<[jq<�.i<W�`<��X<q�P<	iH<�@@<�8<{�/<��'<>�<�<Tr<7P<]�;A�;���;ڢ�;�r�;�M�;|7�;C2�;M�z;��Z;�<;;��;y�:���:�%|:s�:Š
8ğ߹�Xg�����X��I����.�5 K��!g��X��9㎻�*���+��U⵻-K»eλ�-ڻs�廼�𻌨�����;��8�������a�9��9/$��f(��,��y0�W4�!8���;��E?���B�
F��UI���L�Z�O�]�R�]�U���X�Z�[��^�7�a�|d��]g�F;j��m�E�o�ܴr��|u��=x�J�z�a�}�9-�������ӂ�$��Is��A�1�� a�����X���X����������\��򴒼:���d��ֻ��<��;e������E���W��������wA��ʏ���ޣ��/�����|֧� -��f����߫��:��e���I��M��z�������Y��'������X��s�������P���  �  Y�N=�GN=^�M=�L=�BL=�K=J�J=O5J=ބI=�H=e#H=
sG=5�F=F=�eE=n�D=�D=�_C=e�B=	B=�]A=ر@=S@=�W?=5�>=`�==HH==�<=��;=�.;=�y:=d�9=�9=�X8=��7=��6=�66=>�5=2�4=Q4=BX3=��2=*�1=F"1=�`0=�/='�.=�.=�9-=g,=��+=��*=��)=��(=?(=Z''=�8&=�E%=M$=`N#=I"=�<!=�' =p
=��=�=�w=�1=6�=|�=�=y�=�1=�=�=�=��=9=��	=��==lH=m{=D� =\��<���<�<E�<Uh�<���<���<���<)��<���<��<��<��<8��<�t�<`g�<�Y�<�K�<�=�<�.�<��<g�<f��<`�<LΝ<�<���<X|�<�]�<�=�<��<G��<�y<k}q<gBi<�
a<��X< �P<!yH<O@<�'8<M0<��'<й<�<|q<�L<�P�;	�;���;y��;�R�;�*�;N�;�	�;&.z;�uZ;��:;-�;���:J�:9V{:�N:I<8W��g�����k����d�.�y�J���f��=���Ď�
���	��ÿ��$)»�Dλ;ڻ��z��^�����j7��6�!�����f�����8$��r(���,��0�#h4�m)8�e�;�lX?��B�"F��eI���L�M�O��R���U���X���[�y�^�ԓa�}wd��Vg��1j�%m�r�o�f�r��ku��+x���z�(�}�U$��?y��̂�]���m����������^��������Z��°������a��$���{��m��kĖ�f���n������0���_����������G��3���3⣼�1������0֧��+������p۫�u5��2���민�E��ş�������P�����[����P��&���l����J���  �  ,�N=IN=�M=8�L=`BL=��K=��J=<3J=/�I= �H=�H=oG=��F=�F=taE=�D=�D=\C=��B=B=)[A=�@=�@=�V?=�>=��==%I==q�<=��;=1;=�|:=��9=�9=�\8=;�7=;�6=�:6=8�5=��4=�4=[3=�2=��1=^#1=<a0=�/=��.=�.=8-=�d,=�+=d�*=�)= �(=
(=#'=�4&=�A%=I$=�J#=�E"=�9!=�% =�=��=��=x=�2=��=��=u!=��=v5=�=!=��=��=�==f�	=W�== L=�~=� =a��<���<��<�E�<�g�<���<|��<��<���<��<t��<��<5��<Wx�<�k�<�^�<�Q�<VD�<�6�<�(�<��<�	�<���<�<Ν<��<Ǜ�<��<2b�<�C�<T$�<��<��y<�q<�Ti<�a<�X<G�P<̇H<+\@<�28<�
0<�'<ý<1�<yp<tI<}D�;\��;k��;�m�;5�;��;��;��;/�y;�(Z;n�:;�R;p�:��:i�z:ެ :b6�7��	�g����(��.��݄.���J��f�+%��ި���뛻�騻j����	»|&λ#�ٻ�s延��$������3�,5���_���k�*��YB$�Q~(�ǚ,�٘0��x4��:8��;�j?�\�B�{2F��tI���L���O�y�R��U���X�~�[��^��a�Xsd�pPg�7)j�S�l���o�H�r��[u�Dx���z��}�-���q��'ł�9���h�������
��]��r���L���[����������f�����0���t���̖�#��Lw���ɚ�����g��ƴ��� ���L��z���w壼�3��惦�֧�.*��F����׫��0��u����䯼o>������c�H������M���6I�������F���  �  ��N=JN=��M=L�L=�AL=��K=R�J=`1J=�I=C�H=�H=�kG=f�F=�F=�]E=b�D= D=�XC=�B=uB=�XA=$�@=�@=!V?=��>=��==�I==��<=S�;=,3;=B:=��9=�9=g`8=Ȫ7=��6=j>6=��5=��4=>4=S]3=��2=.�1=B$1=�a0=�/=��.=�.=�6-=�b,=��+=��*=��)=��(=v	(=['=�0&=�=%=�E$=�G#=7C"=�7!=�# =�=��=>�=;x=�3=��=<�=�#=f�=�8=��=�$=��=��=B=a�	="�=�=:O=I�=� =���<���<�<�E�<�f�<�~�<���<+��<���<R��<���<ه�<�|�<�p�<�c�<"W�<VJ�<�=�<�0�<�#�<��<j�<w��<��<�͝<ж�<���<���<f�<~H�<*�<n�<��y<�q<�ci<�+a<��X<�P<W�H<g@<�;8<�0<4�'<��</�<1o<�E<�9�;J��;h��;�V�;\�;��;�͜;HÌ;�y;��Y;Qc:;�;���:�@�:t�y:A :��7�����g����z�麓��jp.�'�J�i�f�������dқ�Ϩ�_���Z���pλ��ٻU_廁��_x�����0�4���=���p�����J$�Y�(���,���0���4�nI8�L�;�Vy?��B��@F�	�I�{�L��O���R�~�U��X�9�[���^���a�pd�,Kg�"j�Z�l�.�o��r��Nu�]x���z��z}�P��k��1�����Bd��J�������[���������)]�������k��Nƒ�:!��K{���Ӗ�r*���~��	њ�� ���n��!���R��;Q��L���W裼�5��鄦�֧�+)��F~���ԫ��,�������ޯ�$8�����Y鳼�@���������B��̗���컼B���  �  ��N=�JN=��M=F�L=�AL=ёK=;�J=�/J=~I=�H=XH=iG=��F=	F=�ZE=p�D=OD=,VC=��B=gB=8WA=��@=�@=uU?=H�>=��==9J==o�<=��;=�4;="�:=��9=19=c8=��7=��6=,A6=�5=0�4=C4=_3= �2=/�1=�$1=�a0=Л/=z�.=�.=Q5-=Ga,=��+=L�*=t�)=��(=�(=j'=.&=;%=C$=ME#=A"=�5!=^" =k=#�=�=Ix=�3=��=}�=V%=h�=�:=G�=�'=Տ=��=4E=�	=��=<=�Q=E�=�� =0��<y��<��<�E�<�e�<5}�<4��<��<���<ʒ�<��<O��<�v�<j�<�]�<)Q�<�D�<�8�<D,�<��<U�<��<��<��<�͝<>��<�<Ą�<i�< L�<e.�<]�<��y<��q<�oi<�7a<�Y<|�P<��H<o@<�B8<:0<��'<��<��<n<C<�0�;���;���;�D�;�;�լ;��;���;iy;��Y;�0:;��;���:i�:(Zy:rU�9�<�7z2⹢h������麡���`.���J�ˊf�������M���Q���oo��`���;�ͻ�ٻP廲��n��O��.��3������kt����gQ$��(�̯,��0���4�:U8�a�;�o�?���B��KF��I�ĸL���O�o�R���U��X���[�c�^��a��md�]Gg��j���l�7�o��r��Du�dx���z��o}����+f������>��a��ȳ������Z��˯��R��r^���������{n��Rʒ��%��O���aٖ�S0�������֚��&��t��򿞼�
���T��f����꣼Y7������(֧��(���|���ҫ�*��!����گ�h3�������㳼V;�����U跼>������黼?���  �  ��N=CKN=>�M=B�L=OAL=T�K=|�J=�.J=�|I=��H=�H=hgG=��F=AF=�XE=��D=��C=�TC=�B= B=VA=ѫ@=� @=U?=�>=��==�J==�<=H�;=�5;=T�:=P�9=�9=�d8=1�7=>�6=�B6=��5=��4=�4=`3=�2=��1=C%1=b0=��/=,�.= .=�4-=I`,=p�+=�*=��)=0�(=�(=�'=P,&=^9%=^A$=�C#=�?"=�4!=o! =�=��=��=Nx=B4=>�=F�=U&=��=m<=�=�)=��=��=G=X�	=��=�=�R=w�=�� =���<���<[�<�E�<le�<|�<���<��<���<���<̈�<�~�<Ls�<�f�<5Z�<zM�<OA�<X5�<i)�<;�<G�<0�<��<�<^͝<���<ǟ�<��<�j�<rN�<11�<��<l�y<o�q<�vi<�>a<�Y<�P<��H<,t@<�F8<i0<�'<�<��<2m<4A<�*�;8��;���;89�;��;�Ƭ;���;���;�Iy;��Y;�:;p�;vq�:�¹:�y:���9��77��7h������޸�EW.���J�wyf������s��"��������b������ͻ��ٻ F廒}��g��	�-�3�����v�6���U$��(�{�,�U�0���4�g\8��<���?��B��RF�d�I�t�L���O���R��U���X���[��^�^�a�ald��Dg�yj���l�#�o�$|r��>u��w��z�3i}����c������_��E������Z���������B_��Q�������p���̒��(�������ܖ��3�������ښ�<*��{w��Þ�k��?W��O���*주c8��J���@֧�)(��|��yѫ�F(�����د�i0�������೼�7��ӎ��!巼;��ܐ���滼>=���  �  :O=�UN=��M=	�L=SML=Q�K=!�J=:J=Y�I=��H="H=mpG=�F=�F=�cE=;�D=gD= fC=��B=B=�qA=��@=##@=�z?=��>=%>=Lx==�<=�<=|j;=g�:=�:=�U9=\�8=��7=�=7=��6=��5=L"5=�l4=R�3=�2=�C2=W�1=��0=^0=l?/=�u.=h�-=H�,=|,==*+=�N*=�o)=k�(=��'=m�&=�%=��$=Q�#=w�"=T�!=� =��=c�=}u=O?=��=$�=�V=��=�=%=O~=��=�Q=��=��=�G
=C�=��=��=_!=�F=���<j��<�%�<B�<HT�<�\�<b]�<@V�<%I�<q7�<p"�<��<���<n��<��<
��<���<.��<�y�<�h�<wW�<�D�<�0�<��<��<��<�ȕ<7��<}��<]d�<?@�<��<��y<ڤq< ]i<�a<��X<+�P<�QH<@<�7<(�/<rf'<�,<(�<��<v<.l�;���;ql�;n��;���;�"�;ԙ;��;��r;6�R;v33;ϩ;̹�:[��:l�Y:ɂ�9��ӸyX�]���@A���O���g��V8�<�T��q�Ym�����q�������\����ǻ=Ի�߻���h���v� ��'�cO�cQ��/�n��Ճ���"�5S'�+�+�4�/���3�0j7�[;��>��(B�A�E�b�H��K�d�N���Q�)�T��W���Z�@}]�oN`��c���e�7�h��qk��2n���p�8�s�^v��y�V�{�@b~�C����Ӂ��"���p����������[����������R������z��\�� �������p��˕�$���y���̙����g����������l:��j~��~¢����O�������䧼�3���9ث�7-��J����ٯ��0��s����ݳ�'3��#����ܷ�k0��
����׻��+���  �  � O=�UN=��M=�L=vML=��K=r�J=r:J=�I=7�H=�"H=4qG=��F=�F=�dE=�D=5D=�fC=b�B=�B=rA=�@=q#@=�z?=��>=(%>=;x==��<=v<=j;=�:=.:=
U9=��8=��7=�<7=ŉ6=�5=�!5=\l4=۵3=��2=�C2=:�1=��0=y0=�?/=v.=��-=��,=,=�*+=NO*=lp)=<�(=��'=W�&=��%=��$=�#=�"=��!=}� =�=��=�u=Z?=��=�=}V=@�=��=z=�}=!�=�P=��=��=G
=g�=4�=��=� =6F=��<���<\%�<�A�<YT�<Q]�<�]�<W�<DJ�<�8�<�#�<�<���<P��<���<ǲ�<-��<ƌ�<V{�<j�<oX�<�E�<~1�<�<)�<��<�ȕ<¨�<Ά�<|c�<'?�<M�<��y<��q<dYi<ka<��X<!�P<POH<�@<��7<}�/<je'<�+<�<��<�v</n�;Y��;�p�;i��;z��; )�; ۙ;ݣ�;@s;�	S;:B3;W�;���:���:��Y:�ž9s�Ҹ�A�B���w:���L��Lh��Y8���T�� q��p�����v�������b��g�ǻ�Ի��߻v�뻷����� ��(��O�KQ� /�������T�"�lQ'���+�~�/���3��f7�;�'�>��$B��}E�1�H�n�K���N�2�Q�V�T���W�v�Z��|]��M`��c�M�e�'�h�sk�t4n�(�p���s��`v�}y�Խ{��e~������ԁ��#���q������]���[��竉������Q��>���� ��][��"���Y��Po���ɕ��"��.x���ʙ����qe�����r���"9��C}������7���N��X����䧼�3��3����ث��-��<���ۯ� 2��눲�/߳��4��ĉ��	޷��1��,����ػ��,���  �   O=#UN==�M=2�L=�ML=?�K=|�J=�;J=z�I=�H=�$H=zsG=+�F=TF=gE=��D=�D=iC=a�B=mB=�sA=T�@=l$@=Z{?=��>=(%>=�w==J�<=�<=�h;=S�:=^:=S9=z�8=��7=�:7=��6=��5=�5=�j4=u�3=��2=�B2=��1=��0=�0=@/=�v.=ש-=�,=�,=�,+=lQ*=�r)=��(=�'=��&=A�%=��$=#�#=��"=�!=�� =�=V�=�u=c?=6�=D�=~U=��=�~==U{=��=%N=	�=��=}D
=�=��=��==�D= ��<o��<�$�<�A�<�T�<�^�<�_�<�Y�<vM�<f<�<.(�<��<���<Z��<��<׷�<��<A��<W�<�m�<n[�<OH�<]3�<<�<��<��<ȕ<@��<���<�`�<�;�<I�<��y<@�q<�Oi<�	a<6�X<^�P<XGH<�@<c�7<�/<Db'<�)<��<��<�x<�u�;?��;.}�;0�;���;R<�;��;I��;�7s;�5S;;m3;Y�;��:��:�kZ:o��9}и� ����e/��_M���m��c8�p�T��5q��}��#������⡮��s����ǻ1*Ի�
���������� �G+�>Q��Q��-�o�����"��K'�؀+�ɕ/��3��]7�#;�)�>��B�tE�ĲH���K�
�N�c�Q���T�,�W���Z�pz]�M`�c��e��h�'wk��9n���p�A�s�Niv�>y���{��n~�
���ف��'��u���D��H]����������@Q����� ����X��0������`k���ŕ����Gs���ř�����`������C�v5��z�������M��~���䧼/4��I���yګ�D0��+����ޯ�
6��*����㳼h9��4���Mⷼ�5�������ۻ�/���  �  ��N=9TN=بM=A�L=jNL=C�K=��J=�=J=�I=��H=!(H=wG=��F=NF=%kE=��D=_D=lC=��B=2B=�uA==�@=�%@=D|?=j�>=%>=`w==D�<=�<=�f;=ִ:=x:=�O9=�8=�7=77=�6=��5=�5=h4=3�3=��2=�A2=�1=��0=�0=�@/=�w.={�-=:�,=A,=�/+=�T*=Sv)=}�(=�'=��&=�%=��$=h�#=��"=��!=�� =��=D�=ov=Z?=��=:�=�S=��=,|=b�=�w=��=�I=Ǥ=��=L@
=�=m�=��=a=�B=���<G��<k#�<�A�<�U�<�`�<�b�<�]�<tR�<cB�<�.�<1�<w�<���<8��<ؿ�<���<M��<���<s�<`�<�K�<�5�<��<U�<>�<�ƕ<���<�<�[�<6�<��<��y<ňq<9@i<�`<+�X<�wP<�:H<� @<;�7<�/<\]'<H'<��<�<c|<���;�;���;��;���;]Z�;u�;�ۉ;s;�{S;Q�3;6!;��:!^�:U%[:��9�J̸ǣ�<s��� ��N���v��u8��U��Wq�����*:������4����3ȻTCԻ�!��뻮���#� ��/��S�R��,�(��z���"��B'�_v+�l�/�<|3��N7�Y;���>��
B�@dE��H��K���N���Q���T�9�W�3�Z�[w]��K`��c���e��h�~k��Bn�Eq�I�s��vv��(y�v�{�C}~�6����߁�k-��)z��Mƅ�}��s_��ǭ��
���~P��N���k���CU������m
��e������B��bk����������X��Z����鞼�/�� u�������J��C���E䧼�4������1ݫ�4������䯼C<������과�@������:鷼<��O���y໼�2���  �  ��N=�RN=/�M=?�L=OL=��K=��J=B@J=��I=��H=R,H=�{G=��F=cF=HpE=��D=>D=qC=��B=� B=�xA=��@=�'@=q}?=��>=�$>=�v==��<=�<=d;=��:=��9=�K9=Y�8=?�7=B27=;6=$�5=�5=sd4=;�3=��2=�?2=�1=�0=0=�A/=uy.=��-=��,=�
,=�3+=
Y*=�z)=c�(=�'=��&=��%=(�$=��#=��"=�!=V� =k�=��=w=<?=��=��=�Q=��=�x=D�=s=��=�D=8�=(�=�:
=�|=��=��=�=�?=H��<,��<�!�<yA�<W�<c�<�f�<�b�<�X�<J�<�7�<�"�<��<��<���<��<T��<X��<���<z�<�e�<sP�<X9�<��<��<|�<aĕ</��<|�<�U�<�.�<6�<��y<�tq<�+i<��`<��X<�dP<*H<�?<?�7<��/<�V'<B#<��<��<�< ��;��;ש�;8=�;(ٺ;���;�:�;��;J�s;g�S;�4;t;�/�:��:�\:�Y�9t\Ǹ�,�N��u���T�������8�c=U���q�����}Y�������஻
���i5Ȼ�dԻ�@ໄ�������� ��5�nW�FS�7+����s���"�v7'��h+��y/��j3��;7�B�:�C�>��A�,PE���H�l�K���N�|�Q���T��W�חZ��s]��J`�Jc���e���h�/�k�LNn�/q�}�s��v�i;y���{�u�~�i���>聼N5��ۀ���˅�����b������|����O����� ����P��©��}�� ]���������Ya��S�������N�����)ូ&(���n��ĵ�����:H��͔��#䧼	6�������ૼ9�����z민�D������l���bJ�����E�zD��ҕ���滼8���  �  N�N=LQN=P�M=*�L=�OL=�K=��J=CJ=��I=��H=1H=�G=��F=N#F=:vE=q�D=�D=/vC=E�B=�$B=?|A=<�@=�)@=�~?=]�>=�$>=�u==	�<=_<=�`;=��:=�9=fF9=�8=��7=�,7=�y6=��5=�5=4`4=��3=��2=�=2=��1=x�0=40=hB/=
{.=ݯ-=��,=D,=�7+=�]*=X�)=�(=�'=��&=��%=v�$=k�#=��"=��!=)� =|�=ڤ=zw=�>=��=ݪ=O=��=rt=Y�=�m=��=5>=��=��=�4
=�v==�=��=�=`<=���<p��<��<�@�<�W�<�e�<�j�<�h�<9`�<�R�<�A�<�-�<K�<�<���<���<���<���<ؖ�<��<cl�<�U�<�<�<�!�<��<]�<���<͜�<!v�<N�<�%�<��<��y<P]q<ki<��`<5�X<2OP<{H<7�?<��7<R~/<nN'<A<�<�<]�<'��;2�;���;�_�;�;}��;uk�;R;�;�At;�=T;�m4;��;��: ��:�]:E�9~������'������`��8����8��hU���q�4Ά��~���须5�� ޻�A_Ȼ��Ի�d�u�����?� ��=�\��T��)�a���l��"��*'�EY+�h/��V3��%7���:�Ph>��A��8E��zH�Z�K�6�N���Q� �T�ثW���Z��o]��I`�O c���e���h�1�k�i\n��!q�Y�s�!�v�{Qy���{�'�~�\�����~>�������҅���6f��̱��%����N�����=����K��(��������S��p������U��q��������C��e����מ�����g���������kE������$䧼�7�������嫼?������2���sN�����������U��I������kN������u>>���  �  ��N=nON=2�M=��L=/PL=-�K=�J=�EJ=4�I=�H=!6H=x�G=��F=�)F=�|E=��D=�%D=�{C=1�B=�(B=�A=��@=n+@=�?=��>=5$>=?t==��<=u<=,];=3�:=�9=�@9=�8=o�7=T&7=�s6=�5=�5=�[4=��3=r�2=N;2=�1=��0=-0=-C/=�|.=2�-=��,=,=i<+=c*=�)=	�(=�'=��&=��%=�$=��#=1�"=W�!=� =��=�=�w=�>=��=��=L=��=�o=��=�g=�=I7=��=��=�-
=jp=F�=U�==�8=��<*��<�<@�<�X�<Wh�< o�<�n�<�g�<�[�<"L�<@9�<�$�<��<���<Y��<K̾<}��<s��<D��<s�<�Z�<M@�<�#�<��<��<}��<���<qo�<�E�<��<��<�y<�Cq<�h<��`<�rX<�7P<H<X�?<�7<sq/<-E'<4<��<�<͉<$��;�H�;���;!��;�+�;�ݪ;���;|q�;S�t;׫T; �4;�6;Փ�:�!�:R3^:���9�M��L7�6�������r�����i�8�^�U���q�򆻏���Z��`9������ȻR�ԻI�໕
�l3��I��F��a��W�R)�����e��"��'�VI+�1U/�'A3��7�w�:�O>���A�C E��cH��K�[�N��Q��T��W�Q�Z�sl]�yI`�n#c��e�!�h�؞k��kn�B4q���s��v��iy�Q|�ѿ~�V��������H��ّ���م�"���j������Y ��XN�����]F��]���K�9J����������OI��ߚ��>ꚼ�7��0���H͞����`��&���T����B��C����䧼�9������꫼�E��ա������+Y��m������Eb���������@Y��Y�������'E���  �  ��N=^MN=�M=\�L=�PL=V�K=��J=�HJ=��I=V�H=;H=�G=j�F=�/F=��E=��D=�+D=��C=��B=-B=�A=��@=)-@=��?=��>=�#>=�r==��<=x<=hY;=��:=��9=;;9=��8=1�7= 7=zm6=J�5=(	5=�V4=��3=�2=�82=�1=��0=�0=�C/=�}.=a�-= �,=�,=�@+=h*=~�)=�(= �'=��&=l�%=��$=v $=��"=��!=�� =��=.�=3x=�==�=u�=�H=��=k=w�=ma=��=J0=_�=Y�=�&
=�i=�=��=[=�4=���<���<�<�>�<vY�<�j�<;s�<�t�<Ao�<�d�<eV�<�D�<�0�<z�<L�<���<�׾< ��<˩�< ��<�y�<o_�<sC�<F%�<a�<���<ۺ�<s��<sh�<1=�<��<��<�yy<�)q<n�h<��`<SYX<sP<��G<�?<7<Zd/<9;'<�<6�<q�<��<½�;_�;r�;���;/U�;��;�њ;ئ�;�u;AU;V@5;И;4F�:��:9?_:`��9�4��Y���儺����\�������8���U��9r����є�C��Uh��t<����ȻJ�Իi���.�#R����P�h�[��)�[���_���"�I'�:+��B/��,3���6�4�:�#6>�ثA� E��LH�E|K�
�N���Q�}�T���W�b�Z�ri]��I`�'c�� f�	�h��k��{n�)Gq�mt���v��y�n1|���~�i���	��S�������ᅼ+(��.o���������:N�����GZA��Е��M뒼�@��
���Oꖼ.=��x����ݚ��+��,x��hÞ�,���X��g���L�-@��]���\姼<�����L��L��S������+d��*���*���n���¶����Vd��k�������[L���  �  �N=HKN=��M=��L=�PL=?�K=��J=KJ=֜I=5�H=t?H=�G=��F=E5F=s�E=H�D=�0D=܅C=F�B=�0B=�A=��@=�.@=n�?=��>=�">=]q==��<=�
<=�U;=x�:=�9=�59=9�8=D�7=7=�g6=õ5=5=8R4=��3=��2=<62=B~1=��0=�0=*D/=.=?�-=��,=%,=�D+=�l*=��)=W�(=��'=X�&=��%=��$=�$=o#=�!=M� =/�=�=@x====��=(�=�E=��=�f=N�=�[==�=�)=��=��= 
=�c=a�=��=�=�0=���<��<E�<}=�<�Y�<il�<�v�<�y�<v�<m�<�_�<AO�<<�<!'�<��<���<��<�ʺ<Q��<9��<*�<�c�<F�<:&�<��<�ޙ<��<F��<�a�<�4�<!�<�ۀ<4by<�q<D�h<�`<AX<�P<D�G<��?<�~7<�W/<Q1'<=<��<�<̐<W��;�r�;`�;��;�z�;�7�;| �;�׊;��u;�{U;ߠ5;L�;���:�N�:t.`:��9�²�Zf��Є��������v��h9���U��ur��:�������m������i��8�Ȼ]ջ��8Q��o���MY��n�Q^�>*�I���Z���"�C'�,+�62/��3���6��:�4>�ޔA���D��7H�kiK�X�N���Q���T���W�`Z��g]��J`��*c��f���h���k�f�n��Xq�� t���v�W�y�/I|���~��ǀ�����\������%酼'.���s������X��uN��͛��{뎼=�����䒼N8��m����ߖ�2������Қ�� ��n��b���F��yR��f�����.>������T槼\>����������S��q�������n��^ʲ��#���z���ζ�����n��ջ�����jS���  �  ��N=kIN=h�M=4�L=�PL=�K=��J=MJ=q�I=e�H==CH=-�G=^�F=:F=D�E= �D=R5D=�C=��B=�3B=~�A=��@=�/@=��?=��>=">=�o==��<=�<=�R;=��:=��9=519=E|8=&�7=�7=�b6=�5=��4=6N4=-�3=��2=�32=�|1={�0=.0=gD/=�.=ɷ-=��,=�,=5H+=�p*=�)=�(=l�'=�&=M�%=�%=�$=�#=��!=L� =��=��=:x=�<=8�=�=-C=��=�b=��=�V=��=�#=�}=��=h
=&^=Y�=6�=�=}-=I��<���<�<'<�<�Y�<�m�<�y�<�}�<�{�<�s�<�g�<X�<uE�<�0�<��<z�<��<�Һ<T��<��<̓�<�f�<H�<�&�<,�<�ܙ<���<���<�[�<�-�<���<rҀ<�My<��p<��h<%j`<�+X<��O<�G<��?<q7<`L/<�('<<��<��<#�<���;���;1�;���;C��;\�;�'�;��;��u;�U;��5;�>;.r�:�Ů:v�`:�N�9��!�:�������V������
A9�,V��r�BZ�����!���ɻ������eɻ-3ջ�໶o�����'��a��t�
b�O+����TV���"�'�&�x +�f$/��	3�8�6�c|:��>�w�A�&�D�/&H�7YK�yzN��Q���T� �W�M{Z�2f]�9L`��.c�6f���h���k��n��hq�2t��v�P�y��]|���р�M��xe��>�����3���w������	���N��ؚ��,鎼r9��I���ޒ�#1��-����֖��(��by��ɚ����te���������� M��M����꣼�<������h秼�@������p����Y������3���w��#Բ�.������ض��)��x��)ĺ�	���Y���  �  ��N=�GN=i�M=��L=�PL=^�K=��J=�NJ=k�I=��H=FH=U�G=��F=�=F=�E=��D=�8D= �C=��B=*6B=\�A=��@=�0@=J�?=��>=t!>=�n==�<=�<=
P;=��:={�9=�-9=hx8='�7=�7=�^6=2�5=.�4=K4=}�3=��2=22=M{1=��0=�0=�D/=��.=�-=d�,=,=�J+=�s*=�)=m�(=	�'=��&=��%=�%=�$=#	#=��!=�� =~�=!�=x=�;=�=��=A=��=�_=/�=�R=��=�=3y=0�=�
=�Y=z�=��=��=�*=!��<���<R�<;�<�Y�<�n�<�{�<��<��<y�<�m�<�^�<�L�<d8�<I"�<�
�<3�<�غ<���<���<3��<Ci�<aI�<?'�<�<ۙ<��<���<�V�<(�<��<-ˀ<�=y<��p<V�h<AY`<�X<��O<�G<�?<pf7<gC/<�!'<J <��<��<��<D��;n��;�A�;���;n��;]w�;F�;�!�;�v;�V;�/6;�w;��:��:�a:�5�9�x������������������]9�	OV���r��r��j6��X���2گ������,ɻ�OջZử��n���y0��h�qy��d�R,�����S�2�"�L�&��+��/���2���6��m:���=��rA���D��H�0MK�pN�T�Q���T�c�W��xZ��e]�hM`��1c�
f���h���k�e�n�uq��?t��w�	�y��m|���ـ��$��)l��?������7��*{��ӿ��k��/O��V����玼�6������sْ��+��~��Ж�[!��
r���������_��򬞼����I��J��� 飼�;������U觼�B��f���R���|^��.�������~���۲��5��!����඼f1�����ʺ����Z^���  �  E�N=�FN=��M=L�L=�PL=��K=��J=jOJ=��I=X�H=�GH=S�G=��F=�?F=.�E=��D=�:D=�C=d�B=�7B=z�A=��@=51@=��?=w�>=!>=n==޹<=�<=kN;=�:=`�9=O+9=�u8=��7=m7=:\6=ժ5=��4=I4=��3=1�2=�02=_z1=
�0=�0=�D/=�.=��-=X�,=N,=UL+=Tu*=$�)=��(=8�'=��&=��%=	%=x$=�
#= "=�� =�=h�=x=|;=Z�=e�=�?=6�=�]=��=;P=�=�=hv=e�=7
=ZW=
�=��=��=8)=g��<���<��<L:�<�Y�<�o�<
}�<���<���<j|�<�q�<�b�<HQ�<�<�<�&�<>�<i��<�ܺ<���<9��<9��<�j�<9J�<Y'�<��<�ٙ< ��<<��<�S�<X$�<��<�ƀ<�3y<��p<ϓh<�N`<[X<��O<�G<G�?<�_7<�=/<f'<�<��<��<��<��;ڕ�;�K�;��;�»;���;�X�;T5�;q@v;�8V;�U6;}�;h�:W�:w�a:��9�⪸��������������'��o9�nfV�'�r������G���¢�!��¼�r?ɻ	bջN)Ử������6�m��|�g�<-�t���Q�B�"�D�&�R+�V/��2���6�e:���=��iA���D��H��EK�fiN��}Q���T�{�W��vZ�
e]�eN`��3c��f�,�h�s�k�;�n��|q�xHt�7w���y��w|����ހ�4)��lp�� �������:��_}��w���_���O��񙍼�掼Q5��~����֒�[(��4z���˖�����m��M���i��[��V��������F��w����磼;������
駼�C��e���� ���a���®��#��#����಼�:������嶼86�������κ�X��va���  �  ��N=�FN=��M=+�L=�PL=��K=��J=�OJ=�I=��H=jHH= �G=��F=�@F=�E=��D=�;D=��C=��B=8B=܋A=�@=U1@=��?=_�>=� >=�m==��<=<=�M;=A�:=��9=�*9=$u8=��7=7=_[6=�5=3�4=nH4=�3=��2=�02=z1=��0=i0=�D/=	�.=Ź-=��,=�,=�L+=�u*=Ԛ)=F�(=�'=��&=��%=�	%=$=5#=q "=� =C�=u�=x=P;=�=�=:?=��=�\=:�=`O=	�=�=du=c�=O
=}V=8�=��=:�=�(=���<%��<��<:�<�Y�<�o�<�}�<���<s��<�}�<�r�<|d�<�R�<�>�<�(�<��<���<�ݺ<�¶<��<߉�<k�<RJ�<5'�<��<_ٙ<s��<q��<�R�<�"�<e�<�Ā<�0y<��p<�h<�J`<�X<��O<�G<��?<Z]7<8</<'<J�<��<R�<��<���;���;XO�;��;�ǻ;���;>_�;�<�;�Ov;�FV;�b6;S�;�-�:Ph�:Lb:M��9Ǉ��C��~���7�������� v9��oV�o�r�]���N���ɢ�p���ʼ�<Fɻdhջr/���ʰ���7�]n�~��g��-�w��wQ�[�"���&��+�1/���2�Ӹ6�b:���=�)fA���D��H�/CK�8gN�|Q�0�T���W��vZ�
e]��N`��4c��f���h�Q�k���n�nq��Kt�gw�-�y�}{|��"�)����*���q��R���6���`;��~�������O��虍�p掼�4�������Ւ�@'���x��dʖ�l���k�������
���Y��2��������E��ӕ��f磼�:��֐��H駼^D���������b��Į�%������Ⲽ�<�������綼�7��(���-к�����b���  �  E�N=�FN=��M=L�L=�PL=��K=��J=jOJ=��I=X�H=�GH=S�G=��F=�?F=.�E=��D=�:D=�C=d�B=�7B=z�A=��@=51@=��?=w�>=!>=n==޹<=�<=kN;=�:=`�9=O+9=�u8=��7=m7=:\6=ժ5=��4=I4=��3=1�2=�02=_z1=
�0=�0=�D/=�.=��-=X�,=N,=UL+=Tu*=$�)=��(=8�'=��&=��%=	%=x$=�
#= "=�� =�=j�=x=;=]�=j�=�?==�=�]=�=FP=��=�=yv=y�=M
=rW=$�=��= �=V)=���<��<,�<�:�<�Y�<�o�<?}�</��<���<�|�<�q�<c�<SQ�<�<�<�&�<0�<S��<�ܺ<���<��<
��<�j�<J�<"'�<��<�ٙ<쮕<��<�S�<2$�<��<gƀ<�3y<��p<ϓh<�N`<|X<	�O<U�G<��?<�_7<)>/<�'<��<n�<��<$�<���;���;TL�;3�;Eû;��;Y�;n5�;^@v;�8V;U6;��;$�:ST�:1�a:��9C�����ϸ�����@���L�r9�vhV��r�w����H���â���Gü�@ɻ�bջ�)������)6�+m��|�,g�O-�����Q�M�"�L�&�Y+�\/�"�2���6�
e:���=��iA���D��H��EK�giN��}Q���T�|�W��vZ�
e]�fN`��3c��f�,�h�s�k�;�n��|q�xHt�7w���y��w|����ހ�4)��lp�� �������:��_}��w���_���O��񙍼�掼Q5��~����֒�[(��4z���˖�����m��M���i��[��V��������F��w����磼;������
駼�C��e���� ���a���®��#��#����಼�:������嶼86�������κ�X��va���  �  ��N=�GN=i�M=��L=�PL=^�K=��J=�NJ=k�I=��H=FH=U�G=��F=�=F=�E=��D=�8D= �C=��B=*6B=\�A=��@=�0@=J�?=��>=t!>=�n==�<=�<=
P;=��:={�9=�-9=hx8='�7=�7=�^6=2�5=.�4=K4=}�3=��2=22=M{1=��0=�0=�D/=��.=�-=d�,=,=�J+=�s*=�)=m�(=	�'=��&=��%=�%=�$=%	#=��!=�� =��=%�="x=�;=!�=��=A=��=�_=B�=�R=��=�=Uy=W�=$
=+Z=��=��= =+=���<^��<��<�;�<Z�<Oo�<|�<g��<)��<by�<n�<�^�<�L�<j8�<>"�<�
�<�<�غ<^��<<��<ن�<�h�<�H�<�&�<�<�ڙ<���<\��<|V�<�'�<���<�ʀ<�=y<��p<U�h<`Y`<�X<��O<m�G<��?<g7<%D/<�"'<<��<Ѻ<e�<���;��;�B�;���;\��;x�;�F�;�!�;�v;�V;Q.6;/v;���:_�:�a:��9��Q��3�����������a9��RV���r��t��8��߱���ۯ�Ѱ���-ɻ�Pջ;�r������0��h��y�'e�v,����S�F�"�]�&��+�/���2��6��m:���=��rA���D��H�2MK�
pN�U�Q���T�d�W��xZ��e]�hM`��1c�
f���h���k�e�n�uq��?t��w�
�y��m|���ـ��$��)l��?������7��*{��ӿ��k��/O��V����玼�6������sْ��+��~��Ж�[!��
r���������_��򬞼����I��J��� 飼�;������U觼�B��f���R���|^��.�������~���۲��5��!����඼f1�����ʺ����Z^���  �  ��N=kIN=h�M=4�L=�PL=�K=��J=MJ=q�I=e�H==CH=-�G=^�F=:F=D�E= �D=R5D=�C=��B=�3B=~�A=��@=�/@=��?=��>=">=�o==��<=�<=�R;=��:=��9=519=E|8=&�7=�7=�b6=�5=��4=6N4=-�3=��2=�32=�|1={�0=-0=gD/=�.=ɷ-=��,=�,=5H+=�p*=�)=�(=l�'=�&=N�%=�%=�$=�#=��!=O� =��=��=@x=�<=B�=�==C=��=�b=��=�V=��=%$=�}=��=�
=h^=��=��=*=�-=���<���<,�<�<�<cZ�<�n�<6z�<Q~�<|�<Rt�<$h�<IX�<�E�<�0�<��<T�<H�<vҺ<�<���<M��<[f�<�G�<Q&�<��<*ܙ<)��<��<[�<O-�<V��</Ҁ<qMy<l�p<��h<Qj`<X,X<S�O<��G<x�?<r7<kM/<�)'<9<��<��<P�<��;���;�2�;���;���;]�;�(�;��;��u;�U;,�5;z<;�k�:��:S�`:c(�9����2��̄����#���|���F9��1V�Z�r��\�����I���½��]����ɻ�4ջF���p�����:(�b�u�Hb��+����wV��"�?�&�� +�u$/��	3�C�6�k|:��>�|�A�*�D�2&H�:YK�{zN��Q���T�!�W�M{Z�2f]�:L`��.c�7f���h���k��n��hq�2t��v�P�y��]|���р�M��xe��>�����3���w������	���N��ؚ��,鎼r9��I���ޒ�#1��-����֖��(��by��ɚ����te���������� M��M����꣼�<������h秼�@������p����Y������3���w��#Բ�.������ض��)��x��)ĺ�	���Y���  �  �N=HKN=��M=��L=�PL=?�K=��J=KJ=֜I=5�H=t?H=�G=��F=E5F=s�E=H�D=�0D=܅C=F�B=�0B=�A=��@=�.@=n�?=��>=�">=]q==��<=�
<=�U;=x�:=�9=�59=9�8=D�7=7=�g6=õ5=5=8R4=��3=��2=<62=B~1=��0=�0=)D/=.=?�-=��,=%,=�D+=�l*=��)=W�(=��'=X�&=��%=��$=�$=q#=!�!=Q� =3�=�=Gx=F==��=8�=�E= �=�f=o�=�[=j�=�)=Ճ=��=` 
=�c=��=�=*=81=w��<���<�<M>�<xZ�<'m�<tw�<6z�<�v�<�m�<#`�<�O�<(<�<*'�<��<���<;�<6ʺ<ر�<���<�~�<�b�<YE�<�%�<(�<*ޙ<n��<���<a�<w4�<��<�ۀ<�ay<�q<B�h<�`<�AX<R	P<�G<��?<�7<�X/<�2'<�<_�<��<<�<��;u�;��;��;�|�;�8�;G�;P؊;~�u;�zU;̞5;W�;B��:�E�:v`:���9����E���ބ�J��^������o%9�wV�||r��=�������p��z����k��-�Ȼջ��ໍR�#q�����Y�o��^�~*�~���Z���"�`'�,+�I2/��3���6��:�<>��A���D��7H�niK�Z�N���Q���T���W�aZ��g]��J`��*c��f���h���k�f�n��Xq�� t���v�W�y�/I|���~��ǀ�����\������%酼'.���s������X��uN��͛��{뎼=�����䒼N8��m����ߖ�2������Қ�� ��n��b���F��yR��f�����.>������T槼\>����������S��q�������n��^ʲ��#���z���ζ�����n��ջ�����jS���  �  ��N=^MN=�M=\�L=�PL=V�K=��J=�HJ=��I=V�H=;H=�G=j�F=�/F=��E=��D=�+D=��C=��B=-B=�A=��@=)-@=��?=��>=�#>=�r==��<=x<=hY;=��:=��9=;;9=��8=1�7= 7=zm6=J�5=(	5=�V4=��3=�2=�82=�1=��0=�0=�C/=�}.=a�-=��,=�,=�@+=h*=~�)=�(= �'=��&=m�%=��$=x $=��"=��!=�� =��=4�=<x=>=�=��= I=��=<k=��=�a=��=�0=��=��='
=-j=��=C�=�=5=���<���<��<�?�<VZ�<ek�< t�<3u�<�o�<ne�<�V�<E�<1�<��<7�<}��<�׾<���<D��<���<�x�<�^�<�B�<y$�<��<��<��<���<�g�<�<�</�<B�<yy<a)q<l�h<8�`<�YX<( P<��G<$�?<�7<�e/<�<'<D<��<�<Y�<���;�a�;��;ϩ�;�V�;��;�Қ;:��;gu;�U;>5;��;�=�:�:�'_:7X�9���_��f������z�����f 9�>�U��@r���EԔ�F��k���>���Ȼ:�Ի��w0�kS��]��P�}h�V[��)�����_���"�j'�:+��B/��,3���6�?�:�,6>�߫A�E��LH�I|K��N���Q��T���W�c�Z�si]��I`�'c�� f�	�h��k��{n�*Gq�mt���v��y�n1|���~�i���	��S�������ᅼ+(��.o���������:N�����GZA��Е��M뒼�@��
���Oꖼ.=��x����ݚ��+��,x��hÞ�,���X��g���L�-@��]���\姼<�����L��L��S������+d��*���*���n���¶����Vd��k�������[L���  �  ��N=nON=2�M=��L=/PL=-�K=�J=�EJ=4�I=�H=!6H=x�G=��F=�)F=�|E=��D=�%D=�{C=1�B=�(B=�A=��@=n+@=�?=��>=5$>=?t==��<=u<=,];=3�:=�9=�@9=�8=o�7=T&7=�s6=�5=�5=�[4=��3=r�2=N;2=�1=��0=-0=-C/=�|.=2�-=��,=,=i<+=c*=�)=	�(=�'=��&=��%=�$=��#=3�"=Z�!=� =��="�=�w=�>=��=Ө=!L=��=�o= �=�g=P�=�7=ё=��=�-
=�p=��=��=�=�8=���<��<��<A�<�Y�<3i�<�o�<no�<zh�<\�<�L�<�9�<�$�<��<���<#��<�˾<��<矶<���<Qr�<�Y�<~?�<�"�<��<��<���<���<�n�<3E�<R�<��<��y<gCq<�h<ĳ`<FsX<I8P<H<��?<t�7<�r/<�F'<�<5�<��<w�<O��;�K�;_��;h��;�-�;`ߪ;��;�q�;�t;�T;��4;�3;��:,�:^:ڞ�9H8��aV�d�� ��|��������8�8�U�|r�����ݪ��g��+<��m��Y�ȻS�Ի����4����+G�b�X��)�����e�7�"�'�rI+�GU/�9A3��7���:�O>���A�I E��cH��K�^�N�
�Q��T�	�W�R�Z�tl]�zI`�o#c��e�"�h�؞k��kn�B4q���s��v��iy�Q|�ѿ~�V��������H��ّ���م�"���j������Y ��XN�����]F��]���K�9J����������OI��ߚ��>ꚼ�7��0���H͞����`��&���T����B��C����䧼�9������꫼�E��ա������+Y��m������Eb���������AY��Y�������'E���  �  N�N=LQN=P�M=*�L=�OL=�K=��J=CJ=��I=��H=1H=�G=��F=N#F=:vE=q�D=�D=/vC=E�B=�$B=?|A=<�@=�)@=�~?=]�>=�$>=�u==	�<=_<=�`;=��:=�9=fF9=�8=��7=�,7=�y6=��5=�5=4`4=��3=��2=�=2=��1=x�0=40=hB/=
{.=ݯ-=��,=D,=�7+=�]*=X�)=�(=�'=��&=��%=v�$=l�#=��"=��!=-� =��=�=�w=
?=��=�=#O=��=�t=~�=�m=��=o>=�=��=�4
=Kw=��=�==�<=��<^��<� �<�A�<�X�<�f�<�k�<ci�<�`�<<S�<�A�<.�<u�<#�<���<���<3��<%��<Q��<w��<�k�<�T�<<�<!�<��<��<���<��<}u�<�M�<"%�<���<�y<]q<ii<��`<��X<�OP<gH<U�?<=�7<�/<�O'<�<��<��<��<6��;�4�;z��;�a�;��;ٯ�;Wl�;�;�;wAt;�<T;4k4;8�;���:�u�:�]:��9ڹ¸��k7��~���p��8����8�rpU���q��ц�����졻����໻paȻ��Իlf�������� �*>��\�RU�:*�����l�-�"��*'�_Y+�h/��V3��%7� �:�Xh>��A��8E��zH�^�K�8�N���Q��T�٫W���Z� p]��I`�O c���e���h�2�k�j\n��!q�Z�s�!�v�{Qy���{�'�~�\�����~>�������҅���6f��̱��%����N�����=����K��(��������S��p������U��q��������C��e����מ�����g���������kE������$䧼�7�������嫼?������2���sN�����������U��I������kN������u>>���  �  ��N=�RN=/�M=?�L=OL=��K=��J=B@J=��I=��H=R,H=�{G=��F=cF=HpE=��D=>D=qC=��B=� B=�xA=��@=�'@=q}?=��>=�$>=�v==��<=�<=d;=��:=��9=�K9=Y�8=?�7=B27=;6=$�5=�5=sd4=;�3=��2=�?2=�1=�0=0=�A/=uy.=��-=��,=�
,=�3+=
Y*=�z)=c�(=�'=��&=��%=)�$=��#=��"=�!=Y� =p�=��=w=F?=��=ì=�Q=�=�x=e�=;s=��=�D=s�=k�=7;
=O}=�=��=>=6@=��<��<�"�<JB�<�W�<�c�<^g�<tc�<gY�<�J�<�7�<#�<��<��<���<���<��<���<E��<�y�<Pe�<�O�<�8�<>�<>�<��<�Õ<���<|{�<,U�<.�<��<q�y<�tq<�+i<��`<��X<�eP<�*H<�?<f�7<��/<�W'<�$<-�<+�<T�<���;m�;!��;1?�;�ں;΂�;�;�;:�;�s;=�S;�4;q;(�:|ܫ:��[:�*�9j'ȸ�G� \�����Xc��)����8�0DU�t�q�����Z\��/ġ�K㮻:���^7Ȼ`fԻ1B��������E� �j6��W��S�v+�R���s��"��7'��h+��y/��j3��;7�K�:�J�>��A�1PE�ĐH�o�K���N�~�Q���T���W�ؗZ��s]��J`�Kc���e���h�0�k�MNn�/q�~�s��v�i;y���{�u�~�i���>聼N5��ۀ���˅�����b������|����O����� ����P��©��}�� ]���������Ya��S�������N�����)ូ&(���n��ĵ�����:H��͔��#䧼	6�������ૼ9�����z민�D������l���bJ�����E�zD��ҕ���滼8���  �  ��N=9TN=بM=A�L=jNL=C�K=��J=�=J=�I=��H=!(H=wG=��F=NF=%kE=��D=_D=lC=��B=2B=�uA==�@=�%@=D|?=j�>=%>=`w==D�<=�<=�f;=ִ:=x:=�O9=�8=�7=77=�6=��5=�5=h4=3�3=��2=�A2=�1=��0=�0=�@/=�w.={�-=:�,=A,=�/+=�T*=Sv)=}�(=�'=��&=�%=��$=i�#=��"=��!=�� =��=I�=uv=b?=��=G�=�S=��=C|=}�=�w=��=J=��=��=�@
=Z�=��=�=�=C=e��<���<$�<lB�<�V�<!a�<kc�<1^�<�R�<�B�<+/�<f�<��<���<)��<���<P��<���<L��<�r�<�_�<XK�<j5�<Y�<��<��<ƕ<5��<|��<y[�<�5�<��<E�y<��q<7@i<B�`<��X<xP<z;H<�@<,�7<(�/<|^'<u(< �<C�<�}<���;$
�;���;� �;O��;[[�;�;	܉;�~s;�zS;��3;�;Ӑ�:�V�:/[:ݨ�9��̸¹��~��H,���Y���|�^{8�yU�]q�}����<��顡�-��������Ȼ�DԻ�"���뻟����� �0��S�]R��,�S��;z���"��B'�sv+�|�/�I|3��N7�a;��>��
B�DdE���H��K���N���Q���T�:�W�4�Z�\w]��K`��c���e��h�~k��Bn�Eq�I�s��vv��(y�v�{�C}~�6����߁�k-��)z��Mƅ�}��s_��ǭ��
���~P��N���k���CU������m
��e������B��bk����������X��Z����鞼�/�� u�������J��C���E䧼�4������1ݫ�4������䯼C<������과�@������:鷼<��O���y໼�2���  �   O=#UN==�M=2�L=�ML=?�K=|�J=�;J=z�I=�H=�$H=zsG=+�F=TF=gE=��D=�D=iC=a�B=mB=�sA=T�@=l$@=Z{?=��>=(%>=�w==J�<=�<=�h;=S�:=^:=S9=z�8=��7=�:7=��6=��5=�5=�j4=u�3=��2=�B2=��1=��0=�0=@/=�v.=ש-=�,=�,=�,+=lQ*=�r)=��(=�'=��&=B�%=��$=$�#=��"=��!=�� =	�=Y�=�u=i?==�=M�=�U=�=�~=�=k{=��=CN=+�=%�=�D
="�=+�=�=K=E=y��<���<%�<cB�<qU�<_�<.`�<�Y�<�M�<�<�<b(�<��<���<`��<���<���<ۣ�<��<�<Ym�<[�<�G�<�2�<��<E�<&�<�Ǖ<⦑<O��<L`�<f;�<�<��y<�q<�Oi<�	a<u�X<��P<�GH<e@<�7<ښ/<c'<�*<��<��<�y<cw�;���;�~�;T�;���;=�;�;|��;�7s;�4S;l3;��;��:��:�_Z:nw�9��и������7���U���q��g8�\U��9q�N���$��8���G����t����ǻ2+Ի�໽�뻠����� ��+�rQ��Q�.�������"��K'��+�ԕ/��3��]7�(;�.�>��B�tE�ƲH���K��N�d�Q���T�-�W���Z�qz]�M`�c��e��h�'wk��9n���p�A�s�Niv�>y���{��n~�
���ف��'��u���D��H]����������@Q����� ����X��0������`k���ŕ����Gs���ř�����`������C�v5��z�������M��~���䧼04��I���yګ�D0��+����ޯ�
6��*����㳼h9��4���Mⷼ�5�������ۻ�/���  �  � O=�UN=��M=�L=vML=��K=r�J=r:J=�I=7�H=�"H=4qG=��F=�F=�dE=�D=5D=�fC=b�B=�B=rA=�@=q#@=�z?=��>=(%>=;x==��<=v<=j;=�:=.:=
U9=��8=��7=�<7=ŉ6=�5=�!5=\l4=۵3=��2=�C2=:�1=��0=y0=�?/=v.=��-=��,=,=�*+=NO*=lp)=<�(=��'=W�&=��%=��$=�#=�"=��!=~� =	�=��=�u=\?=��=��=�V=G�=��=�=�}=.�=�P=��=��=$G
=�=N�=��=� =UF=W��<*��<�%�<.B�<�T�<�]�<^�<=W�<mJ�<�8�<$�<1�<���<S��<���<���<��<���<2{�<�i�<@X�<�E�<H1�<��<��<��<�ȕ<���<���<Vc�<?�<5�<��y<{�q<dYi<|a<��X<R�P<�OH<@<U�7<ޞ/<�e'<b,<��<�<�v<o�;��;Rq�; ��;���;~)�;<ۙ;���;.s;�	S;�A3;u�;w��:���:��Y:Ϸ�9	Ӹ�I�r����>���P��qj��[8���T��"q��q��h���v��M����c����ǻ	Ի%�߻ی������ ��(��O�bQ�/�������_�"�uQ'���+���/���3�g7�;�)�>��$B��}E�2�H�o�K���N�2�Q�W�T���W�v�Z��|]��M`��c�M�e�'�h�sk�t4n�(�p���s��`v�}y�Խ{��e~������ԁ��#���q������]���[��竉������Q��>���� ��][��"���Y��Po���ɕ��"��.x���ʙ����qe�����r���"9��C}������7���N��X����䧼�3��3����ث��-��<���ۯ� 2��눲�/߳��4��ĉ��	޷��1��,����ػ��,���  �  �O=paN=�M=�M=JZL=��K=�J=	EJ='�I=<�H=�)H=UwG=��F=F=�kE=�D=�D=�uC=��B=�.B=u�A=��@=�E@=�?=�>=�Q>=H�=={�<=`N<=G�;=w�:=+B:=��9=�8=@38=k�7=m�6=+#6=hr5=��4=j4=gZ3=u�2=�1=�01=r0=Ư/=v�.=&.=�P-=,=ҩ+=a�*=$�)=)=?7(=dS'=�k&=��%=ҏ$=�#=�"=��!=o� =�i={C==
�=.�=�-=9�=|V=��=2O=��=H=�q=�=�=�>	={r=�=��=��=���<)�<#9�<�G�<oK�<E�<�5�<��<��<M��<��<��<r�<#O�<�.�<��<V��<>޺<1ȶ<���<
��<���<'p�<�U�<;8�<��<?��<4Α<�<|�<�P�<0%�<��y<�q<�Di<��`<��X<NP<� H<��?<�m7<�&/< �&<K�<,K<��<ͪ<e��;.��;7J�;ԝ�;���;�d�;+�;}�;�hl;�L;D	,;
@;ps�:�:v�9:v�x9(�q��\6�������Ӻ)���b%���B�P�_�{|�����䙻*l�����A���9λl�ڻ�w���bX��K#�:p	�������j���-�!�N"&�.r*���.���2�0�6� ^:�r>�ăA���D��#H��FK��ON��BQ�%#T�U�V��Y�d}\�P9_��a�תd��ag��j���l��}o��,r���t�w�P"z�O�|�U\����� D�����DՄ�\���e��ӯ������J�����������H������� ��=^������F��p��NŘ�����a������일	,���i��Φ��䢼�"��Vd��
���C��<��͋��3ݫ��0��D����گ�0��:����ٳ��-��ʀ��ӷ��$��v��@ǻ����  �  lO=HaN=�M=	M=xZL=F�K=��J=�EJ=�I=�H=�*H=]xG=��F=/F=mE=N�D=�D=�vC=��B=�/B=8�A=C�@=[F@=!�?=@�>=�Q>=8�==H�<=�M<=��;=��:=fA:=Ǒ9=�8=>28=b�7=q�6=6"6=�q5=/�4=�4=�Y3=(�2=��1=�01=?r0=��/=��.=�.=�Q-=�,=��+=]�*=+�)=,)=_8(=�T'=m&=��%=͐$=��#=ʛ"=*�!=� =�i=�C==��=��=&-=��=�U=��=6N={�==�p=��=�=�=	=yq=#�=��=B�=���<��<�8�<�G�<�K�<�E�<�6�<��<.�<���<���<��<ft�<lQ�<�0�<H�<���<\�<ʶ<ϴ�<���<1��<q�<OV�<�8�<��<,��<�͑<��<�z�<hO�<q#�<��y<Җq<*@i<��`<l�X<JP<P�G<T�?<Ok7<�$/<��&<��<K<�<��<h��;���;1P�;|��;��;gm�;��;#��;3|l;�*L;�,;PS;��:�:��9:Yy9�Sq��>6�j���}�Ӻ����b%�8�B�;�_��&|����뙻�r��(�������'@λY�ڻ�}�@��\���$�1q	�Ӕ����Zi�����!� &�]o*�V�.�_�2�%�6��Y:���=�'A��D�LH�kBK��KN��>Q��T���V�ǺY��{\�m8_�_�a��d�jbg��j���l�"�o��/r�/�t�؂w�6&z�i�|�e`������E�������ք�}���f��G�������J��j������H������#����\������;���m�������i_������ꝼ*��h��6����⢼�!���c��������<������ݫ��1������,ܯ��1��-����۳��/��ǂ���Է�t&���w���Ȼ����  �  X
O=�`N=��M=2	M=[L=F�K=��J=^GJ=�I=��H=~-H=p{G=�F=�F=wpE=��D=/D=�yC=v�B=62B=B�A=��@=�G@=
�?=��>=�Q>=�==��<=�L<=+�;=��:=	?:=�9=�8=8/8=T7=v�6=e6=o5=�4=4=�X3=5�2=k�1=�01=�r0=��/=��.=(!.=vS-=�,==�+=B�*=F�)=�)=�;(=�W'=tp&=��%=��$=s�#=�"=�!=F� =�j=&D=5=��=0�=�+=��=�S=<�=MK=8�=�=m=!�=L�
=<:	=�n=��=��=��=��<��<�7�<�G�<�L�<jG�<?9�<u#�<z�<	��<���<X��<B{�<mX�<8�<7�<��<��<�϶<���<���<���<�s�<X�<�9�<��<:�<�ˑ<\��<(w�<�J�<!�<��y<1�q<+3i<��`<ՌX<V>P<��G<q�?<.d7<�/<��&<n�<�J<��<ٮ<���;��;a�;}��;��;M��;�	�;आ;��l;�gL;�W,;ӊ;%��:�^�:qf::�}{9σo���5�ߓ��i�ӺT��Ph%���B���_�}A|�E/������B���tǴ�T���lVλl�ڻN��E)�i���)��t	�t������g�v�۪!��&��g*�&�.��2�F�6�0M:�#�=�,qA��D��H��5K��?N�m4Q��T���V���Y�-w\�d5_���a�"�d�Ddg�nj���l��o�8r��t��w�2z���|��l����`K��s����ڄ��!��2i��㱈������I��u���`qE��Y���(����W��S���6���g��������X������㝼a$��c��ߠ��7ߢ����a��a�����m=��P����߫�r4��D����௼�6��録��᳼�5��ˈ���ڷ��+��|��b̻����  �  �O=�_N=9�M=h	M=�[L=��K=�J=JJ=`�I=q�H=�1H=K�G=1�F=�!F=�uE=�D=K$D=[~C=��B= 6B=m�A={�@=�I@=\�?=u�>=�Q>=T�==E�<=�J<=��;=��:=3;:=Ȋ9=u�8=R*8=oz7=��6=�6=�j5=��4=	4=\V3=��2=��1=x01=�r0=��/=��.=g#.=ZV-=��,=E�+=��*=2�)=�!)=A(==]'=�u&=|�%=�$=e�#=N�"=��!=U� =gl=�D=H=	�=�=�)=F�=2P='�=�F=�=-=pg=s�=��
=!5	=�i={�=[�=��=���<@�<�6�<�G�<�M�<,J�<d=�<�(�<]�<��<���<d��<��<�c�<C�<%�<h	�<�<"ض<��<ݩ�<���<Ww�<�Z�<�:�<��<��<�ȑ<���<q�<|C�<��<��y<�uq<[i<��`<�xX<�+P<\�G<*�?<�X7<0/<��&<X�<BJ<� <׳<	��;"�;�{�;���;�=�;X��;�5�;8ӆ;3m;��L;s�,;��;6��:�:>`;:F�~9S�l��c5��g��ʵӺ<���r%���B�O�_��m|�~J����������봻���tzλ��ڻٮ滕C�Q���1��y	�A��ˑ�ve�����!�Q&��[*���.�R�2��t6�9:���=�d[A�<�D�n�G��!K�p-N��#Q�KT���V�+�Y�.p\��0_���a���d�dgg�E"j�t�l�M�o��Er��t���w�Ez�0�|�!�����S��?���]ᄼ'��/m�����������I��9����덼�A��\�������tP��ԫ�����W]��|�������M������ڝ�w��&[�� ����٢�����^������
�>��[���J㫼99��[����篼K?�������볼�?�������㷼4�������һ��!���  �  'O=�]N=��M=�	M=�\L=��K=��J=�MJ=��I=c�H=�7H=��G=��F=�(F=�|E=��D=�*D=t�C==�B=�:B=n�A=��@=L@=��?=<�>=�Q>=j�==~�<=GH<=�;=@�:=6:=�9=I�8=�#8=�s7=W�6=6=�e5=ݵ4==4=QS3=��2=;�1= 01=Us0=��/=��.=?&.=�Y-=�,=k�+=��*=�*=_()=�G(=d'=@|&=ȏ%=͝$=l�#=��"=�!=� =n=�E=A=�=�=6'=��=�K=��=h@=Q�=�	=�_=��=��
=[.	=�c=�=ƹ=!�=j��<�<�4�<�G�<�O�<�M�<�B�<�/�<�<q��<���<l��<���<�q�<SQ�<�2�<��<��<�<wʲ<ñ�<ɗ�<�{�<d]�<�;�<�<�<cđ<f��<�h�<�9�<$
�<��y<�Zq<�i<O�`<�^X<GP<u�G<h�?<�H7<9
/<y�&<��<I<^<��<���;�<�;���;r�;�l�;6�;_o�;4�;��m;�?M;8*-;�P;i�:��:�<:�z�9�i�t�4��3����Ӻg����%���B�� `��|��n��UG��Dا�:���»B�λ��ڻ���sf�>���=���	����Ւ�3c���!�E&�{L*��s.�$y2�]6�:���=�9?A��D��G��K��N��Q�/�S���V�E�Y��g\�o+_���a���d�8lg�q*j�*�l�v�o��Wr�p
u�+�w�K^z��|��������_������!ꄼR.���r��B�������AJ��ߗ���荼=�����푼G���������/P��ţ�����?��=���p͝���Q�������Ң�}���Z��p����識N?��U����竼�?��k�����^J�����P����L��Z����M?��X����ڻ��(���  �  O=�[N=s�M=q	M=�]L=Y�K=iK=8QJ=?�I=��H=�=H=��G=��F=�0F=�E=��D=j2D=e�C=��B=,@B=�A==�@=�N@=��?=��>=nQ>='�==9�<=E<=ɓ;=�:=0:=O~9= �8=J8=Hl7=�6=�6=5_5=@�4=� 4=�O3=Ĝ2=��1=C/1=�s0=�/=��.=X).=�]-=�,=@�+=�*=�*=0)=�O(=l'=�&=�%=H�$=#�#=S�"=�!=�� =�o=�F==��=�=�#=,�='F=L�=9=N�=n=:W=A�=!�
=\&	=h\=��=P�=��=���<��<"2�<�F�<Q�<2Q�<SH�<�7�<� �<C�<"��</��<���<*��<�a�<�B�<�%�<�	�<Z�<ղ<b��<���<���<1`�<�<�<��<��<ž�<���<_�<�-�<���<̘y<N;q<4�h<
�`<�?X<S�O<U�G<�r?<667<��.<��&<L�<G<f<E�<���;bZ�;���;�/�;ݢ�;�!�;Ű�;uT�;6 n;��M;�-;��;�R�:�s�:��=:FŃ9��e� 4�e���?�Ӻ����%��C�9`�w�|�g���y����%U���G»��λ#ۻ��Ɛ�i����J��	�n��Ӕ�[a��
���!�!�%��;*�_.�a2�B6��:�0�=��A��~D���G�	�J���M���P���S��V�C�Y��^\�?&_�}�a�b�d��rg��4j���l���o�nr��#u��w��{z��}�d��.&��4m��Ա����7��dy��������	K��Ŗ���卼 8��6���M䑼x<�������땼JA�������㙼�/���x�� ������E�� ���ˢ�����V��|����識6A��0������G��B���*���pW��K���S��	\��k���l����L������仼�0���  �  ��N=xYN=�M=	M=h^L=�K=)K=UJ=�I=��H=�DH=�G=��F=O9F=~�E==�D=]:D=��C=�B=�EB=��A=��@=$Q@=�?=T�>=�P>=��==��<=AA<=�;=9�:=h):=�v9=�8=�8=�c7=��6=C6=.X5=�4=M�3=gK3=��2=p�1=0.1=�s0=�/=��.=_,.=b-=�,=E�+=�*=U*=!8)=5X(=Nt'=�&=t�%=�$=�#=@�"=��!=y� =�q=G=v=1�=}=�=1�=@=/�=1=��=/�=�M=��=��
=�	=pT=��=F�=��=���<A�<�.�<�E�<6R�<�T�<�M�<�?�<	+�<|�<L��<���<F��<k��<"s�<�S�<�5�<��<��<�߲<<î<O��<S��<�b�<�<�<��<��<H��<���<T�<� �<��<xy<�q<��h<�j`<sX<��O<��G<�Y?<j!7<��.<�&<�}<�C<�<�<��;�x�;i��;�_�;{۸;_a�;��;���;9�n;�`N;@.;V;�E�:�I�:eo?:�9�Eb��y3��Ж��}Ӻ����%�-FC�^y`�:D}��ʌ�鯚�-J�������»| ϻ�]ۻK=绱������\Z��	�������`�����!�4�%��**��I.�LH2��%6�s�9�=���@��\D�c�G���J�&�M���P�n�S��V�w�Y��U\��!_��a�%�d�_zg�Aj��m�+�o�n�r�O?u���w�V�z�'?}����;6��4|��W���� ���@��"�������}L�����㍼G3��[���Mۑ��1��և��uݕ��1��R����ҙ�����h�����t����9��~��.â��	��OS��ퟦ���C��Ț������WP��.����	���e����������l��ྶ�6��[�����𻼲9���  �  ��N=�VN=f�M=vM=�^L=��K=�K=�XJ=��I=e�H=+KH=i�G=z�F=�AF=��E=k�D=,BD=�C=X�B=&KB=�A=�@=bS@=I�?=��>=�O>=��==��<=H=<=�;=L�:=�":=Ho9=�8=�8=m[7=r�6=e�5=�P5=��4=��3=�F3=;�2=�1=�,1=9s0=ܵ/=��.=./.=�e-=�,=&�+=��*=�*=@)=l`(=�|'=Փ&=إ%=��$=Ŷ#=�"=`�!=�� =�r=mG=�=O�=
z=�=��=�9=�=�(=��=��=D=�=��
=�	=HL=U}=�=x�=���<>�<�*�<TD�<�R�<�W�<3S�<CG�<�4�<l�<�<:��<���<w��<+��<[d�<!E�<�&�<{�<Z�<�ˮ<z��<c��<�d�<�<�<H�<��<T��<�}�<�H�<Y�<�ހ<�Vy<��p<��h<�F`<��W<.�O<fxG<	@?<�7<w�.<֧&<�t<�?<�<��<k�;
��;�;���;��;ҟ�;n:�;]�;�Ho;f�N;��.;�;�2�:��:�@:%Q�9w�^���2���� zӺ�����%�VyC��`�{�}�����6蚻���zӵ���»�_ϻ��ۻ;t�������j�d�	�/��a���`�����!�(�%�9*��5.�02�
6���9��^=��@��:D��G�%�J�p�M�Z�P�%�S���V��yY��M\�_���a�طd�W�g��Mj�!m�r�o�e�r��[u��x�a�z�a}�����F������A̓����K��P����Ȉ�
��cN�������/������ґ��&��Y{��Rϕ�"��s������m���X��:���9螼s.���t��˻�����*P��Ԟ����F�����������Y��o������t���ϲ�u(���}���϶�F���i��^���z���IC���  �  /�N=TN=��M=�M=�^L=��K=�K=�[J=��I=y�H=QH=�G=��F=IF=��E=��D=HID=`�C=�B=PB=ħA=�@=@U@=.�?=p�>=�N>=��==��<=h9<=)�;=��:=�:=h9=-�8=�8=]S7=��6=��5=J5=��4=��3=�B3=Ւ2=��1=j+1=�r0=H�/=��.=�1.=`i-=C�,=y�+=��*=�"*=OG)=�g(= �'=�&=��%=��$=��#=%�"=��!=#� =
t=sG=�=S�=w=�=�=�3=�=,!=?�=��=�:=��=��
=h	=�D=hv=��=x�=���<4 �<'�<[B�<S�<�Y�<�W�<�M�<�=�<?(�<��<?��<���<��<���<ts�<HS�<c3�<��<��<�Ү<ư�<���<�e�<�;�<x�<�ݕ<d��<�t�<�=�<g�<Ѐ<j7y<9�p<�xh<�$`<B�W<��O<^\G<a'?<��6<��.<��&<�k<�:<G<��<p'�;��;�2�;���;�D�;�ب;�x�;0'�;�o;�wO;&M/;TP;�
�:֟:mB:F�9$\��q2�����JӺ���\�%��C�la��}��,��������:���û�ϻ?�ۻf�给�7��N{��	���J��b�L��Nz!���%��*�r#.�2���5��9��@=�Y�@�D�bG�=�J�T�M�X�P���S�u�V�,oY��G\��_�;�a�(�d���g�[j�(m��o���r��vu�@.x���z�9�}����V��	����ڃ�X���T��K����Έ�T���P��U���Oߍ��+��Xz��Kˑ�r��p�������d��w���J���;J��Ɠ��9ܞ�$��Sl��_���S ���M��[���}�.J��F������b��Uî��#�������޲�^8��捵��߶�p-��x��'�������L���  �  ��N=yQN=�M=�M=�^L=b�K=`
K=.^J=!�I=�I=VH=��G=��F=�OF=
�E=I�D=JOD=�C=��B=TB=�A=OA=�V@=ê?=1�>=�M>=��==��<=�5<=܀;=w�:=G:=�a9=n�8=��7=[L7=��6=k�5=D5=+�4=��3=�>3=��2=X�1=�)1=r0=y�/=��.={3.=l-=ߠ,=��+=�*=G(*=tM)=En(=X�'=/�&=?�%=ּ$=<�#=��"=�!=Ȗ =�t=OG=�=]�=;t=$=i�=t.=ة=f=߀=(�=�2=	�=��
=	=�==Wp=��=��=S��<���<1#�<c@�<�R�<q[�<:[�<YS�<�D�<91�<M�<��<{��<J��<���<;��<9_�<>�<��<K��<�خ<�<��<if�<�:�<��<6ٕ<���<�l�<�3�<��<_À<�y<?�p<�Zh<�`<��W<�|O<DG<�?<�6<&�.<Վ&<�c<�5<<��<4�;0��;�N�;���;o�;	�;���;O_�;.Bp;v�O;��/;��;Y��:.q�:�C:׋9,�Y�o2����ՋӺ��!&���C��=a�o4~��V��M�����E��X:ûC�ϻvܻO�继G��Z�������	�?������c����yu!���%�_ *�i.��2���5���9��'=�C�@� D��HG��xJ��M�3�P��S���V�gY�C\��_�U�a���d�B�g� gj�67m�Fp���r���u�EHx��z�;�}�����c��Φ��惼�"���]������rԈ�S��S�����Oލ��(���u��!ő�����f���������eW������g��=��i���&Ҟ����_e��0�������L��O���"���|M��*����	���j���̮��.��ˎ��B첼*F��웵�u��:��z���M˺�c���T���  �   �N=rON=u�M=�M=�^L=еK=�K=�_J=��I=�I=�YH=�G=` G=eTF=�E=�D=�SD=�C={ C=WB=L�A=�A=�W@=
�?=��>=�L>=)�==��<=3<=r};=z�:=�:=�\9=<�8=1�7=�F7=j�6=Y�5=l?5=�4=F�3=�;3=E�2=��1=�(1=yq0=y�/=��.=�4.=n-=��,=$�+=�+=�,*=R)=s(=$�'=ͥ&=}�%=��$=u�#=8�"=��!=� =<u=
G=�=��=�q=D=ܣ=A*=�=!=/{=6�=�,=�y=�
=n�=�8=�k=��=|�=���<M��<! �<�>�<rR�<�\�<�]�<`W�<wJ�<8�<Q!�<��<+��<A��<��<ډ�<(h�<7F�<�#�<� �<ݮ<෪<���<�f�<�9�<	�<sՕ<Ӟ�<f�<,�<0�<q��<Ry<۠p<�Ch<��_<��W<�gO<�0G<� ?<��6<�.<��&<�\<�1<�<U�<�<�;���;�c�;C��;��;�-�;�՘;뉈;��p;�?P;50;c;#F�:�:�C:c��9`>X�@�1�bw��p�Ӻ�#�k9&��D�0na��n~�Ax��r��r��n��-dû��ϻd+ܻL���g��v�������	���ڪ��e�L��[r!���%���)�&	.�_�1���5�9��=�~�@�E�C��5G�gJ��M���P���S�]{V�[aY�@\�4_�S�a�Q�d�S�g��pj�?Cm��p�m�r�(�u�d\x�{���}��&��n������&�*���d��P����؈����U�������ݍ� '���r����������_��r�������M�������蚼�4������ʞ�-��5`��s���p����J����������4P��������Jq���Ԯ�U7��^��������P��ߦ��'���E��%���Ժ�"��b[���  �  l�N=NN={�M=YM=�^L=�K=3K=aJ= �I=�I=\H=��G=FG=iWF=��E=E=�VD=��C=�C=�XB=��A=�A=FX@==�?=��>==L>=�==S�<=B1<=B{;=��:=�:=�Y9=�8=��7=qC7=��6=(�5=l<5=E�4=��3=�93=��2=<�1=�'1=q0=t�/= �.=�5.=To-=/�,=.�+=F+=I/*=�T)=v(= �'=��&=2�%=�$=q�#=��"=�!=�� ={u=�F==��=~p=d=��=�'=�=�=�w=d�=�(=v=8�
=��=N5=�h=��=J�=��<o��<(�<�=�<FR�<7]�<Y_�<�Y�<�M�<E<�<N&�<��<6��<|��<D��<��<�m�<*K�<(�<X�<�߮<���<b��<�f�<�8�<Z�<�ҕ<|��<�a�</'�<~�<��<��x<h�p<?5h<2�_<��W<�ZO<�$G<�><W�6<��.<T&<RX</<�<X�<B�;��;Vp�;��;�;�D�;��;Y��;��p;uP;�>0;h0;4��:�,�:�8D:��9|KW�P�1�|u��)�Ӻ�0��L&��D��a�ԓ~���������5�������~ûMлDܻr軎|�Ո������	����ܭ�9g����p!�7�%���)�p.���1��5��s9��=�>�@� �C��)G��[J�#zM��P�܄S�KvV��]Y�P>\�_���a�j�d�.�g��vj��Jm��p���r�
�u�ix��{���}�}-���t���������/��i�������ۈ����|V��[����ݍ��%���p��㽑�+��9[��e���d����G�������⚼�.���z���Ş�:��"]��+�������[J����������R��ǰ��#��ju��gٮ��<��v��������W��ŭ��
����K��F����ٺ����_���  �  ��N=�MN=5�M=-M={^L=$�K=^K=oaJ=��I=]	I=�\H=s�G=>G=gXF=�E=E=�WD=r�C=rC=|YB=2�A=HA=eX@=B�?=��>=L>=ș==��<=�0<=uz;=�:=�:=�X9=��8=��7=PB7=ϓ6=�5=f;5=_�4=�3=�83=�2=��1=�'1=�p0=q�/=�.=�5.=�o-=��,=��+=+=40*=�U)=w(=!�'=��&=�%=��$="�#=N�"=}�!=٘ =�u=�F=�=q�=	p=�=͠=�&=�=�=pv=�=�'=�t=��
=��=;4=�g=�=��=��<���<��<;=�<DR�<g]�<�_�<�Z�<O�<�=�<	(�<��<9��<���<Q��<��<�o�<�L�<q)�<p�<s�<���<y��<pf�<<8�<��<�ѕ<:��<C`�<d%�<��<簀<��x<g�p<�0h<<�_<הW<rVO<� G<��><�6<�.<}&<<W<e.<�<��<FD�;~��;u�;��;���;pL�;O��;$��;��p;��P;�O0;�?;-��:�C�:�]D:�ۍ9�W�Y�1�x��A�ӺA5�ST&��$D���a�h�~�����ᑛ�>��󑶻Їû�л�Lܻ�軪��9�������	�3������g�	��p!�1�%� �)� .�	�1�Ҿ5�p9��=�#~@���C��%G�XJ��vM��P�y�S�}tV��\Y��=\��_���a�Q�d���g�	yj��Mm�5p���r��u�Tmx�k{�^�}��/��w����������1���j��Q����܈�y���V�������ݍ��%��Gp��鼑��
���Y������x����E�����������,���x��QĞ����\��h�������?J��ݞ�������R������N���v��ۮ��>������=���Z�����d���M��V����ۺ����(a���  �  l�N=NN={�M=YM=�^L=�K=3K=aJ= �I=�I=\H=��G=FG=iWF=��E=E=�VD=��C=�C=�XB=��A=�A=FX@==�?=��>==L>=�==S�<=B1<=B{;=��:=�:=�Y9=�8=��7=qC7=��6=(�5=l<5=E�4=��3=�93=��2=<�1=�'1=q0=t�/= �.=�5.=To-=/�,=.�+=F+=I/*=�T)=v(= �'=��&=2�%=�$=r�#=¿"=�!=�� =}u=�F==��=�p=k=��=�'= �=�=�w=x�=)=(v=U�
=�=p5=�h=$�=r�=W��<���<|�<�=�<�R�<�]�<�_�<Z�<N�<s<�<s&�<��<D��<���<<��<ҏ�<�m�<K�<�'�< �<o߮<Z��<��<Jf�<P8�<�<�ҕ<;��<�a�<�&�<S�<���<��x<Q�p<?5h<G�_<ęW<[O<3%G<~�><��6<�.<�&<�X<�/<l<��<�C�;��;@q�;��;���;E�;�;}��;z�p;�tP;�=0;</;4��:)�:q0D:��9�sW���1�{��ҪӺ�3��O&��D���a�^�~�*���Њ��6�������ûл�Dܻ�}�D���I����	�������Qg�#���p!�D�%���)�x.���1��5��s9��=�@�@��C��)G��[J�$zM��P�܄S�KvV��]Y�P>\�_���a�j�d�.�g��vj��Jm��p���r�
�u�ix��{���}�}-���t���������/��i�������ۈ����|V��[����ݍ��%���p��㽑�+��9[��e���d����G�������⚼�.���z���Ş�:��"]��+�������[J����������R��ǰ��#��ju��gٮ��<��v��������W��ŭ��
����K��F����ٺ����_���  �   �N=rON=u�M=�M=�^L=еK=�K=�_J=��I=�I=�YH=�G=` G=eTF=�E=�D=�SD=�C={ C=WB=L�A=�A=�W@=
�?=��>=�L>=)�==��<=3<=r};=z�:=�:=�\9=<�8=1�7=�F7=j�6=Y�5=l?5=�4=F�3=�;3=E�2=��1=�(1=yq0=y�/=��.=�4.=n-=��,=$�+=�+=�,*=R)=s(=$�'=ͥ&=}�%=��$=v�#=9�"=��!=� =@u=G=�=��=	r=Q=�=U*=+�===P{=\�=-="z=:�
=��=�8=�k=�=ɿ=N��<���<� �<U?�<S�<]�<E^�<�W�<�J�<f8�<�!�<1�<H��<H��<���<���<�g�<�E�<v#�<� �<�ܮ<\��<���<	f�<�8�<��<�ԕ<V��<�e�<�+�<��<2��<�y<��p<�Ch<��_<�W<ihO<�1G<|?<x�6<�.<��&<�]<�2<�<r�<�>�;���;ke�;���;X��;r.�;!֘;0��;n�p;�>P;�	0;!�;W@�:ߠ:��C:�Ռ9�X���1����`�Ӻs)��>&�JD�Vsa��s~��z��)t��l���o���eûN�ϻ�,ܻj���h��w�����	�B�����e�q��yr!���%���)�6	.�l�1���5� 9��=���@�I�C��5G�gJ��M���P���S�^{V�\aY�@\�4_�S�a�Q�d�T�g��pj�?Cm��p�m�r�(�u�d\x�{���}��&��n������&�*���d��P����؈����U�������ݍ� '���r����������_��r�������M�������蚼�4������ʞ�-��5`��s���p����J����������4P��������Jq���Ԯ�U7��^��������P��ߦ��'���E��%���Ժ�"��b[���  �  ��N=yQN=�M=�M=�^L=b�K=`
K=.^J=!�I=�I=VH=��G=��F=�OF=
�E=I�D=JOD=�C=��B=TB=�A=OA=�V@=ê?=1�>=�M>=��==��<=�5<=܀;=w�:=G:=�a9=n�8=��7=[L7=��6=j�5=D5=+�4=��3=�>3=��2=X�1=�)1=r0=y�/=��.={3.=l-=ߠ,=��+=�*=G(*=tM)=En(=X�'=/�&=?�%=׼$=>�#=��"=�!=̖ =�t=VG=�=i�=Jt=7=��=�.=��=�=�=^�=83=N�==�
=k	=4>=�p=#�=k�=5��<���<$�<EA�<�S�<@\�<�[�<T�<�E�<�1�<��<`��<���<S��<��<��<�^�<�=�<d�<���</خ<9��<B��<�e�<�9�<�
�<xؕ<G��<�k�<Y3�<���<À<;y<��p<�Zh<�`<�W<t}O<�DG<�?<_�6<��.<U�&<e<m7<�<��<7�;���;.Q�;���;�p�;s
�;z��;�_�;�Ap;7�O;~�/;T�;&��:Qg�: �B:w��9�BZ��62�����L�Ӻ���%&�+�C�Ea�_;~�:Z��P�������G���<ûO�ϻEܻ���I��[��q���	����Ц� d����u!���%�{ *��.�2���5���9��'=�J�@�D��HG��xJ��M�5�P��S��V�gY�C\��_�U�a���d�B�g� gj�67m�Gp���r���u�EHx��z�;�}�����c��Φ��惼�"���]������rԈ�S��S�����Oލ��(���u��!ő�����f���������eW������g��=��i���&Ҟ����_e��0�������L��O���"���|M��*����	���j���̮��.��ˎ��B첼*F��웵�u��:��z���M˺�c���T���  �  /�N=TN=��M=�M=�^L=��K=�K=�[J=��I=y�H=QH=�G=��F=IF=��E=��D=HID=`�C=�B=PB=ħA=�@=@U@=.�?=p�>=�N>=��==��<=h9<=)�;=��:=�:=h9=-�8=�8=]S7=��6=��5=J5=��4=��3=�B3=Ւ2=��1=j+1=�r0=H�/=��.=�1.=`i-=C�,=y�+=��*=�"*=OG)=�g(=�'=�&=��%=��$=��#=(�"=��!=(� =t=|G=�=a�=w=�=�=�3=�=]!=y�="�=1;=E�=�
=�	=E=�v=�=��=���<M�<(�<oC�<T�<�Z�<�X�<�N�<e>�<�(�<�<���<���<'��<���<5s�<�R�<�2�<�<��<Ү<⯪<���<�d�<�:�<��<�ܕ<���<�s�< =�<��<�π<�6y<��p<�xh<E%`<��W<j�O<y]G<�(?<(�6<:�.<��&<�m<�<<@<�<+�;k��;�5�;6��;G�;qڨ;�y�;�'�;��o;dvO;hJ/;iL;� �:�ɟ:��A:&�9��\�'�2�x���;�Ӻo��&�Q�C�V
a���}��0��r!���Ĩ�X���ûc�ϻu�ۻV��G � 9���{�x�	�q�����Xb�����z!���%�*��#.�(2��5�(�9��@=�b�@�D�bG�B�J�X�M�[�P���S�w�V�-oY��G\��_�<�a�)�d���g�[j�(m��o���r��vu�@.x���z�9�}����V��	����ڃ�X���T��K����Έ�T���P��U���Oߍ��+��Xz��Kˑ�r��p�������d��w���J���;J��Ɠ��9ܞ�$��Sl��_���S ���M��[���}�.J��F������b��Uî��#�������޲�^8��捵��߶�p-��x��'�������L���  �  ��N=�VN=f�M=vM=�^L=��K=�K=�XJ=��I=e�H=+KH=i�G=z�F=�AF=��E=k�D=,BD=�C=X�B=&KB=�A=�@=bS@=I�?=��>=�O>=��==��<=H=<=�;=L�:=�":=Ho9=�8=�8=m[7=r�6=e�5=�P5=��4=��3=�F3=;�2=�1=�,1=9s0=ܵ/=��.=./.=�e-=�,=&�+=��*=�*=@)=l`(=�|'=֓&=٥%=��$=Ƕ#=��"=d�!=� =s=wG=�=`�=z=�=�=�9=�=!)=��=�=]D=q�=��
=8	=�L=�}=��=�=���<w�<6,�<�E�<T�<�X�<8T�</H�<�5�<�<��<���<���<���<��<d�<�D�<&�<��<��<�ʮ<|��<W��<{c�<y;�<9�<��<b��<�|�<�G�<��<ހ<&Vy<K�p<��h<NG`<�W< �O<�yG<�A?<R7<`�.<�&<w<�A<(	<�<��;ט�;r�;��;�;���;�;�;��;GHo;��N;��.;��;�'�:o�:�@:�9Z�_�3�Ⱦ��@�Ӻ���r�%���C��`���}�7��]욻芨��ֵ���»ybϻ�ۻdv绳��H���k���	����ʜ�/a���!�X�%�_*��5.�&02�
6� �9��^=��@��:D��G�*�J�t�M�^�P�'�S���V��yY��M\�_���a�طd�X�g��Mj�!m�r�o�e�r��[u��x�a�z�a}�����F������A̓����K��P����Ȉ�
��cN�������/������ґ��&��Y{��Rϕ�"��s������m���X��:���9螼s.���t��˻�����*P��Ԟ����F�����������Y��o������t���ϲ�u(���}���϶�F���i��^���z���IC���  �  ��N=xYN=�M=	M=h^L=�K=)K=UJ=�I=��H=�DH=�G=��F=O9F=~�E==�D=]:D=��C=�B=�EB=��A=��@=$Q@=�?=T�>=�P>=��==��<=AA<=�;=9�:=h):=�v9=�8=�8=�c7=��6=C6=.X5=�4=M�3=gK3=��2=p�1=0.1=�s0=�/=��.=_,.=b-=�,=E�+=�*=U*=!8)=6X(=Ot'=�&=u�%=�$=
�#=C�"=¤!=� =�q=%G=�=B�=#}= =R�==@=_�=V1=͙=|�=N=�=P�
=	=�T=�=ۮ=G�=��<��<0�<G�<jS�<�U�<O�<�@�<�+�<.�<���<<��<��<y��<s�<�S�<%5�<��<W��<߲<I®<H��<>��<�a�<�;�<��<w�<N��<��<NS�<! �<G�<lwy<|q<��h<.k`<X<��O<��G</[?<2#7<��.<�&<�<�E<�<H�<��;x|�;���;c�;�ݸ;Cc�;Z��;��;�n;'_N;�<.;�Q;:�:�;�:DO?:�҅9��b���3��喺��Ӻ����%��PC���`�	N}�Wό�6���"N��G���]�»`#ϻA`ۻ�?绡��o���[���	�6������`��ڈ!�e�%��**��I.�fH2��%6���9�"=���@��\D�i�G���J�*�M���P�p�S��V�x�Y��U\��!_��a�&�d�_zg�Aj��m�+�o�n�r�P?u���w�V�z�'?}����;6��4|��W���� ���@��"�������}L�����㍼G3��[���Mۑ��1��և��uݕ��1��R����ҙ�����h�����t����9��~��.â��	��OS��ퟦ���C��Ț������WP��.����	���e����������l��ྶ�6��[�����𻼲9���  �  O=�[N=s�M=q	M=�]L=Y�K=iK=8QJ=?�I=��H=�=H=��G=��F=�0F=�E=��D=j2D=e�C=��B=,@B=�A==�@=�N@=��?=��>=nQ>='�==9�<=E<=ɓ;=�:=0:=O~9= �8=J8=Hl7=�6=�6=5_5=@�4=� 4=�O3=Ĝ2=��1=C/1=�s0=�/=��.=W).=�]-=�,=@�+=�*=�*=0)=�O(=l'=�&=�%=J�$=%�#=V�"=�!=č =�o=�F==��=�=�#=L�=MF={�=U9=��=�=�W=��=��
=�&	=�\=*�=�=B�=���<�<Z3�<-H�<BR�<LR�<XI�<�8�<�!�<��<���<���<ã�<7��<�a�<�B�<D%�<j	�<��<9Բ<x��<���<��<_�<�;�<��<��<ӽ�<֎�<X^�<1-�<'��<$�y<�:q<1�h<[�`<(@X<E�O<��G<,t?<�77<i�.<�&<s�<6I<�<k�<���;/^�;3��;�2�;H��;S#�;���;�T�;�n;��M;��-;x�;�G�:Df�:��=:&��9�|f��C4���^�Ӻ2��l�%�(!C��B`���|�ݞ��4}��Q���X���J»��λ%ۻ
绦�����tK��	���;���a��
�ב!�Q�%��;*�-_.�6a2�*B6��:�=�=��A��~D���G��J���M���P���S��V�E�Y��^\�@&_�}�a�b�d��rg��4j���l���o�nr��#u��w��{z��}�d��.&��4m��Ա����7��dy��������	K��Ŗ���卼 8��6���M䑼x<�������땼JA�������㙼�/���x�� ������E�� ���ˢ�����V��|����識6A��0������G��B���*���pW��K���S��	\��k���l����L������仼�0���  �  'O=�]N=��M=�	M=�\L=��K=��J=�MJ=��I=c�H=�7H=��G=��F=�(F=�|E=��D=�*D=t�C==�B=�:B=n�A=��@=L@=��?=<�>=�Q>=j�==~�<=GH<=�;=@�:=6:=�9=I�8=�#8=�s7=W�6=6=�e5=ݵ4==4=QS3=��2=;�1= 01=Us0=��/=��.=?&.=�Y-=�,=k�+=��*=�*=_()=�G(=d'=@|&=ɏ%=Ν$=n�#=��"=�!=� =%n=�E=M=*�=*�=M'=��=�K=��=�@=��=2
=K`=T�=��
=�.	=d=��=F�=��=��<��<�5�<�H�<�P�<�N�<�C�<�0�<��<��<4��<ö�<ۓ�<�q�<9Q�<�2�<B�<���<d�<�ɲ<�<喪<�z�<n\�<�:�<�<�<�Ñ<���<Rh�<9�<�	�<��y<�Zq<�i<��`</_X<P<��G<��?<lJ7<�/<Q�&<��<K<W<�<1��;^@�;���;�;�n�;��;pp�;��;��m;R>M;z'-;M;_�:���:-�<:�<�9�j��4�	F����Ӻ���,�%��B��	`���|��r��K���ۧ�X���»ìλ��ڻ���!h򻰝���=��	���2���c�O�"�!�p&��L*��s.�;y2�.]6�$:���=�B?A��D��G��K��N��Q�1�S���V�F�Y��g\�p+_���a���d�9lg�q*j�*�l�w�o��Wr�p
u�+�w�K^z��|��������_������!ꄼR.���r��B�������AJ��ߗ���荼=�����푼G���������/P��ţ�����?��=���p͝���Q�������Ң�}���Z��p����識N?��U����竼�?��k�����^J�����P����L��Z����M?��X����ڻ��(���  �  �O=�_N=9�M=h	M=�[L=��K=�J=JJ=`�I=q�H=�1H=K�G=1�F=�!F=�uE=�D=K$D=[~C=��B= 6B=m�A={�@=�I@=\�?=u�>=�Q>=T�==E�<=�J<=��;=��:=3;:=Ȋ9=u�8=R*8=oz7=��6=�6=�j5=��4=	4=[V3=��2=��1=x01=�r0=��/=��.=f#.=ZV-=��,=E�+=��*=2�)=�!)=A(==]'=�u&=|�%=�$=f�#=Q�"=��!=Z� =ll=�D=R=�=��=*=]�=NP=I�=�F=K�=c=�g=��=#�
=w5	=8j=ߗ=ž=:�=���<%�<�7�<�H�<�N�<�J�<#>�<�)�<��<���<]��<���<��<�c�<�B�<�$�<	�<��<�׶<{��<2��<ϐ�<�v�<�Y�<�9�<��<��<ȑ<��<�p�<C�<9�<C�y<�uq<Yi<�`<jyX<�,P<C�G<B�?<�Y7<�/<d�&<�<�K<r<j�<	��;�$�;>~�;���;�?�;���;�6�;�ӆ;�m;��L;5�,;��;��:9�:�I;:f~9Im���5��v��A�Ӻ���z%�
�B���_��t|��M��� ��O���yM���|λ��ڻm���D�~���e2�Wz	�������e���ޣ!�t&��[*�Ӆ.�e�2��t6�9:��=�k[A�B�D�s�G��!K�s-N��#Q�MT���V�-�Y�/p\��0_���a���d�egg�E"j�t�l�N�o��Er��t���w�Ez�0�|�!�����S��?���]ᄼ'��/m�����������I��9����덼�A��\�������tP��ԫ�����W]��|�������M������ڝ�w��&[�� ����٢�����^������
�>��[���J㫼99��[����篼K?�������볼�?�������㷼4�������һ��!���  �  X
O=�`N=��M=2	M=[L=F�K=��J=^GJ=�I=��H=~-H=p{G=�F=�F=wpE=��D=/D=�yC=v�B=62B=B�A=��@=�G@=
�?=��>=�Q>=�==��<=�L<=+�;=��:=	?:=�9=�8=8/8=T7=v�6=e6=o5=�4=4=�X3=5�2=k�1=�01=�r0=��/=��.=(!.=vS-=�,==�+=B�*=F�)=�)=�;(=�W'=tp&=��%=��$=t�#=�"=�!=I� =�j=+D=<=��=:�=�+=�=�S=T�=jK=Y�=�=Dm=S�=��
=x:	=�n=כ=�=��=���<��<�8�<KH�<M�<�G�<�9�<�#�<��<c��<��<���<_{�<tX�<�7�<�<���<5�<2϶<6��<��<��<s�<~W�<9�<I�<��<^ˑ<롍<�v�<�J�<��<E�y<�q<*3i<��`<*�X<�>P<��G<6�?<e7<�/<��&<��<�K<��<��<̹�;��;�b�;��;5�;?��;b
�;%��;X�l;�fL;V,;��;X��:�W�:_V::H6{9k�o�4�5�����Y�Ӻ����m%��B���_�dF|��1��� ��<���Aɴ�����Wλ��ڻl��=*�oj��*��t	�������g�����!��&��g*�6�.���2�Q�6�8M:�*�=�1qA��D��H��5K��?N�n4Q��T���V���Y�.w\�e5_���a�"�d�Edg�nj���l��o�8r��t��w�2z���|��l����`K��s����ڄ��!��2i��㱈������I��u���`qE��Y���(����W��S���6���g��������X������㝼a$��c��ߠ��7ߢ����a��a�����m=��P����߫�r4��D����௼�6��録��᳼�5��ˈ���ڷ��+��|��b̻����  �  lO=HaN=�M=	M=xZL=F�K=��J=�EJ=�I=�H=�*H=]xG=��F=/F=mE=N�D=�D=�vC=��B=�/B=8�A=C�@=[F@=!�?=@�>=�Q>=8�==H�<=�M<=��;=��:=fA:=Ǒ9=�8=>28=b�7=q�6=6"6=�q5=/�4=�4=�Y3=(�2=��1=�01=?r0=��/=��.=�.=�Q-=�,=��+=]�*=+�)=,)=_8(=�T'= m&=��%=ΐ$=��#=˛"=+�!=� =�i=�C==��=��=--=��=�U=��=DN=��=2=�p=Ž=�=�=	=�q=G�=�=j�=���<��<9�<�G�<�K�<�E�<�6�<8 �<e�<"��<!��< ��<tt�<pQ�<�0�<5�<o��<5�<�ɶ<���<O��<툪<�p�<V�<k8�<��<��<t͑<פ�<�z�<>O�<P#�<Y�y<��q<)@i<��`<��X<DJP<��G<��?<�k7<%/<U�&<$�<�K<��<�<���;� �;Q�;F��;2�;�m�;�;G��;|l;`*L;�,;$R;��:y��:P�9:�3y9|q�aI6�����&�Ӻ���te%���B��_�X)|� ��5왻�s�����y����@λ�ڻ/~���>]��)%�Yq	�������qi���ȯ!�+ &�ho*�^�.�f�2�*�6��Y:���=�)A��D�NH�mBK��KN��>Q��T���V�ǺY��{\�m8_�_�a��d�jbg��j���l�"�o��/r�/�t�؂w�6&z�i�|�e`������E�������ք�}���f��G�������J��j������H������#����\������;���m�������i_������ꝼ*��h��6����⢼�!���c��������<������ݫ��1������,ܯ��1��-����۳��/��ǂ���Է�t&���w���Ȼ����  �  �O=rnN=��M=M=EhL=N�K=-K={OJ=��I=��H=S.H=�zG=�F=wF=ioE=��D=)#D=��C=�B=DB=\�A=LA=i@=	�?=�$?=u>=��==l.==��<=��;=+;=6~:=L�9=l$9=�w8=�7=Y7=�q6=��5=25=�h4=8�3=�3=�S2=��1=��0=&#0=	`/=q�.=��-=K�,=�*,=�T+=�|*=��)=9�(=F�'=�'=�$&=<%=�M$=X#=�Y"=Q!=�< =G=<�=s�=�h=�=>�=P8=��=2,=�=t�=&B=��=��=*�	=|*=rP=ao=ه=� =�K�<YW�<�V�<�J�<�3�<P�<{��<c��<���<�R�<e�<��<���<Z��<Ji�<,H�<F+�<��< ��<��<gʪ<��<0��<�p�<wK�<o"�<U��<�Ǎ<疉<�d�<2�<��y<��q<�2i<��`<zmX<�P<{�G< [?<�7<��.<�Z&<<��<�F<��<0��;�;%�;�1�;�Q�;Ӂ�;1ɓ;.�;�ne;��D;�w$;�r;'r�:���:Q:���8����UZ�.F���Ͳ�w�/�4IM��j�G���)���|螭����*Ȼq�Ի 6��=�q�����������c����D��nu �K%�>l)�w�-���1�4�5�j�9��{=��A�k}D���G���J�#�M�/�P���S�#dV�yY�˹[��Z^�i�`�U�c�`;f�v�h��k�o%n���p��gs��v���x��2{�N�}�%)���n��w���\���{7���y������p���H������%㌼�6��o����됼K��y�������i��ė�i��7h�����D��/��,h��j����ѡ�����=��5x��L�������=C������/߫�.1�������د��,��F���5ӳ�/%��wv���Ʒ�T��Xe��%�������  �  SO=BnN=��M=9M=�hL=ƷK=�K=XPJ=��I=��H=�/H=�{G=��F=	F=�pE=�D=�$D=�C=`�B= EB=`�A=!	A=�i@=y�?=%?=�>=��==,.==�<=��;=,*;=)}:=�9=$#9=\v8=��7=7=hp6=��5=55=h4=��3=_3=�S2=��1=*�0=�#0=�`/=0�.=��-=W�,=�+,=7V+=j~*=��)=��(=��'=#
'=&&=g=%=�N$=Y#=�Z"=�Q!=j= =�=\�=Q�=Hh=G=�=\7=U�=�*=��=��=�@=�=5�=��	=#)=3O=an=�=[� =�J�<�V�<�V�<@K�<�4�<��<)��<G��<F��<,U�<B �<0��<���<���<�l�<?K�<8.�<^�<i��<��<+̪<O��<3��<kq�<�K�<Z"�<���<uƍ<J��<�b�<�/�<��y<=�q<�,i</�`<�gX<�	P<��G<�V?<�7<s�.<�X&<<}�<IG<�<���;0�;� �;�:�;_\�;���;֓;�;�;ވe;��D;0�$;�;��:)��:i:���8x���A'Z�q3�����Ư�T�/�)MM�a�j�ă�����q���Χ�����Ȼ��Ի�>ỤE������ʓ����������2���s �%�$�i)���-���1�^�5�޻9��u=��	A�NwD���G���J�D�M���P�#�S��_V��Y���[��X^���`�^�c�c;f���h�=�k��'n���p��ks��v�y�x�8{���}��+��q��ش��w���a9��2{���������I�������⌼#6��A���1ꐼ�H��O���1	��g�����7��:e��孛�1�	-��{e������ϡ����R<��Dw����������YC������ૼm2��=����گ��.��Ȃ���ճ��'��y��Rɷ����fg��굻�����  �  O=�mN=��M=�M=�iL=-�K=�K=�RJ=��I=2�H=�3H=#�G=�F=� F=�uE=��D=)D=�C=!�B=\HB=!�A=aA=zk@=��?=�%?=�>=��==W-==��<=��;=�';=z:=��9=?9=>r8=��7=7=�l6=C�5=i5=�e4=��3=A3=S2=��1=��0=�$0=b/=;�.=4�-=X-=,/,=0Z+=��*=�)=e�(=i�'=�'=E*&=RA%=YR$=\#=�\"=�S!=�> =d=��=�=xg=�=n�=�4=�='=G�=O�=�;=J�=��=h�	=V%=�K=�k=߄=ϗ =I�<V�<NW�<�L�<Z7�<0�<���<��<H��<*]�<�(�<���<E��<S��<�u�<-T�<�6�<��<��<]�<�Ъ<䴦<Õ�<�r�<�K�<�!�<��< Í<���<]�<�(�<��y<7�q<i<��`<#WX<i�O<J�G<�K?<��6<��.<�T&< <��<�I<��<���;+�;�7�;�U�;A|�;ڰ�;8��;Qd�;;�e;9E;8�$;��;�.�:�+�:�B:Î�8�X��+�Y�������֪�3�/�W\M�(�j��ԃ�E�����Zĭ��*��>Ȼ��Ի�Z�>^�d���$����������^��l��o �j�$��`)�?�-�+�1��5���9�xd=��@�1dD���G���J���M�g�P�S��SV�PY�A�[�"R^�[�`�Жc�;f���h�h�k�.n�f�p�pvs��v�=�x�H{�Y�}�4���x����������>��2����������I��G���ጼ�3�������吼�C��󢓼����^��]�������[��h���&眼�$���]��S����ɡ�����b8��Xt�����������C��8����⫼�5���i௼�5��c����ݳ�J0��8����з����Hm������r���  �  �O=MlN=-�M=M=�jL=E�K=�	K=bVJ=�I=}�H=q9H=��G=�F=(F=}E=�D=0D=��C=��B=�MB=u�A=�A=6n@=��?='?=�>=��==�+==N<=��;=w#;=u:=��9=9=�k8=��7=�7=�f6=�5=�5=#b4=8�3=f3=R2=��1=u�0=&0=zd/=]�.=#�-=-=�4,=K`+=^�*=!�)=��(=��'=�'=�0&=[G%=�W$=�`#=�`"=�V!=�@ =�=��=��=�e=b=�=V0=Ů=� =��=�=54=�{=b�=��	=-=�F=Jg=w�=R� =�E�<�T�<�W�<�N�<e;�<��<s��<���<.��<�i�<�6�<�<[��<i��<���<7b�<nC�<k'�<�<��<�ת<4��<]��<�t�<.L�<��<��<a��<<YS�<n�<��y<<fq<6�h<��`<�<X<��O<t�G<9?<��6<��.<SM&<��<ۧ<sM<�<k�;7�;"\�;&��;���;��;[8�;W��;�\f; �E;�^%;)N;i�:�:_�:l��8������X�%Ʃ�k�溝��'�/�3vM�a�j���7��r9����[��DoȻ�)ջ��Ỳ��%���2����K���������5h �6�$�SS)��-�x�1���5���9�I=�Z�@�rFD�ÎG�:�J�r�M�X�P�[}S��?V��X�5�[�H^���`�w�c��:f��h�e�k��8n���p�E�s��*v���x�'a{�~�}�A��W����ǂ����G������Ň�����J��˒��ߌ�0��n����ސ�!;��̘��\���R������j����L�������؜�>���Q����������h���h2���o��򱦼�����C�������櫼�;�������鯼�@��j����과c=�����ݷ��*���v���»�����  �  �O=qjN=p�M=nM=7lL=��K=/K=[J=��I=.�H=AH=.�G=0�F=�1F=��E=w�D=9D=ȕC=O�B=�SB=ٳA=GA=wq@=��?=7(?=4�>=��==�)==|<=.�;=�;=dn:=H�9=�9=c8=E�7=4
7=�^6=ɳ5=�5=!]4=`�3=�3=�P2=G�1=$�0=�'0=5g/=6�.=�-=-=�;,=h+=��*=E�)=�(= (=�'=�9&=O%=~^$=ef#=\e"=Z!=>C =�=)�=��=�c=	=n�=r*=��=�={~=\�=D*=�q=��=��	==�?=_a=�|=� =vA�<�R�<�W�<hQ�<@�<%�<��<H��< ��<�y�<RH�<��<���<��<���<-t�<�S�< 6�<��<���<,�<q��<}��<�v�<�K�<��<��<W��<j~�<yF�<_�<�y<Bq<Q�h<w`<pX<G�O<�nG<� ?<��6<��.<C&<4�<��<YQ<}�<�'�;^[�;��;R��;>�;0�;*��;��;fg;�^F;��%;V�;��:/�:�<:W��8�F���X�;|�����E����/�l�M��k�e��g��4q���/��'����Ȼjջ���{��FS��@E�ױ������)����C` �g�$�C)�v�-��1��5��r9��%=��@� D�DhG�ߏJ��M�K�P��`S�\'V���X��[��<^�&�`�&�c��;f�f�h�>�k�iGn�U�p��s��Fv��x��{�4~�qR������ւ�����R��J���ḋ�[��0M��Ғ���܌��+��.��m֐��0��&����甼�A�������똼�9��ł���Ɯ�,��FB���{������#+���j��ݮ������5E�����G쫼!D��0�������PO�����������N��V���f�w9��߃��nͻ����  �  	O=�gN=<�M={M=�mL=?�K=�K= `J=��I=��H=�IH=ɘG=�F=T<F=��E=0�D=0CD=5�C=��B=0[B=ԹA= A=�t@=,�?=@)?=�>=��==�&==�w<=��;=
;=df:=D�9=9=�X8=��7=* 7=rU6=J�5=a5=W4=��3=\�2=�N2=q�1=��0=�)0=j/=Z�.=l�-=�-=tC,=q+=��*=��)=��(=�
(=$)'=+C&=�W%=:f$=�l#=tj"=�]!=�E =!=�=�= a=�=��=]#=A�= =�s=��=�=f=Y�= �	=t=%7=MZ=w=�� =�;�<�O�<W�<�S�<�D�<�,�<K�<r��<��<���<^\�<[-�< �<,��<O��<���<�f�<�F�<�'�<.	�<=�<�Ʀ<���<x�<iJ�<��<��<p��<�q�<�6�<^��</�y<�q<��h<�K`<��W<��O<LG<�?<m�6<�y.<6&<��<ͤ<�T<'�<�C�;؂�;R��;���;E6�;���;�ޔ;�R�;�g;�G;�&;��;"R�:���::��9m޶�Q7W��2��Aw�ī��/�[�M��dk�JH����������x��4黻��Ȼc�ջ����-����[�w�������G����YX ���$��1)�l-�Ԅ1��z5�N9��<���@�=�C�s<G�OeJ�5qM��cP�S@S�V�S�X��[�[0^���`���c�n>f���h�S�k��Yn��q��s�fhv�/y���{�W@~��f��ʩ��邼�%��`������Շ�L��iP������#ی��'���x��=͐��$���}��ה�/��t���W֘��#��!m��걜��򝼨0���l��O����䢼d#���e��򫦼I���ZG��������6N��﩮�����`������"��ec������� ��K��j���yڻ�|!���  �  �O=�dN=��M=M=qnL=��K=�K=eJ=h�I=bI=�RH=עG=g�F=�GF=�E=��D=�MD=�C=nC=�bB=�A=�A=@x@= �?=�)?=N>=w�==�#==s<=x�;=c;=]:=Q�9=H�8=�M8=��7=1�6=K6=�5=&�4=*P4=-�3=R�2=�K2=-�1=��0=�*0=�l/=a�.=��-=p-=wK,=Cz+=��*=��)=�(=(=4'=`M&=a%=n$=[s#=�o"=~a!=�G =�!=j�=�=�]=��=M�=e=ٕ=x=h=��=�=@Y=��=Z�	=�=�-=bR=�p=�� =�4�<|K�<0V�</U�<pI�<34�<��<��<e��<���<�q�<	D�<y�<���<%��<�<�y�<�W�<]6�<��<)�<%ͦ<֤�<�x�<"H�<z�<;ۑ<��<c�<~%�<��<gZy<��p<r~h<
`<�W<<pO<�%G<��><1�6<wd.<R&&<��<ޠ<QV<�<I_�;���;���;s6�;|��;.ץ;M<�;V��;��h;��G;�v';[C;	��:��:�:� 
9y{��+aV��󨺪c�U���0��N�Q�k��~���ᒻy���Eɮ��=��Uɻ�	ֻ�Y�fD����u������/�������Q ���$�s )�TU-��h1��Y5�@(9��<��]@��C�7G�^8J�GM��=P�BS���U���X��n[��$^���`���c��Bf���h���k��nn��'q�j�s�t�v�+6y���{��m~�i}��Z���9����7��p��P����އ�e���T��0���"ڌ��#��.r��1Đ����eo��Ɣ���� o��Ϳ�����HV������yޝ����]��(���Rڢ�����`��٩������zJ������f����Y��R�������s���β�D&��z���ɶ�����^������+黼H-���  �  �O=FaN=R�M=GM=�nL=P�K=�K=�iJ=c�I=�
I=Y[H=��G=�F=�RF=e�E=��D=dXD=��C=�C=�iB=��A=� A=#{@=��?=
*?=/~>=��==�==�m<=Ѻ;=;=[T:=�9=D�8=8B8=%�7=��6={@6=B�5=��4=�H4=K�3=��2=�H2=p�1=1�0=�+0=o/=��.=��-=�-=BS,=@�+=��*=O�)=1�(=-!(=�>'=LW&=�i%=�u$=�y#=Gt"=�d!=�I =!"=Q�=��=�Y=u�=l�===�=��=%\=ݴ=�=;L=Q�=r�	=�=9$=J=�i==� =�,�<~F�<�S�<�U�<M�<�:�<� �<���<E��</��<,��<.Z�<�.�<��<b��<Ĳ�<Ō�<h�<�C�<��<%��<PҦ<#��<6x�<�D�<@�<ґ<ד�<�S�<��<Ԁ<p-y<[�p<�Mh<��_<C�W<�DO<��F<¿><B�6<[M.<�&<@�<'�<3V<�<\w�;��;�!�;gt�;�ʶ;�*�;���;�;�Si;��H;3(;5�;5��:�&�:��!:��9cU��ͪU��Ĩ�`����30��ON�l�춄��$���I��7��������ɻ�_ֻ������	��M�������^"����>��oM ���$�)�v@-�N1��95�a9�+�<�2@���C���F��J�	M��P��R�5�U�ϞX��_[��^�m�`�Սc�If��i���k�n�9Dq���s���v�L`y�b|���~�T����Ձ����VJ��"���괆��釼b ��"Z������ڌ�B!���l���������ya��w������`Z��ϩ��E����?�������ʝ�����M��܎���Т�,���\������$����N��|������f��MǮ�D(������B䲼�<������඼�+���r��a���h����9���  �  ��N=�]N=ݺM=M=�nL=��K=NK=�mJ=��I=hI=-cH={�G=�G=]F=��E=�	E=�aD=>�C=pC=pB=��A=�$A=i}@=��?=�)?=�|>==�==�==�h<=\�;=��:=}K:=`�9=��8=b78==�7=I�6=k66=��5=j�4=�A4=��3=S�2=E2=Z�1=Y�0=),0=�p/=��.=-�-=y%-=:Z,=X�+=�*=�)=I	)=C+(=tH'=K`&=�q%=�|$=�~#=Zx"=]g!=�J ="=��=ͧ=�U=�=��==݂=�=�P=�=Z�=�?=a�=3�	=��=�=B="c=�} =�$�<�@�<Q�<�U�<�O�<z@�<)�<T�<���<���<��<sn�<�C�<��<���<�ſ<���<�v�<P�<)�<� �<?֦<{��<�v�<�@�<��<�ȑ<χ�<1E�<+�<{��<�y<=�p<�h<��_<gW<IO<��F<��><Ni6<�6.<�&<��<�<�T<�<֊�;���;&M�;���;Y�;�v�;]�;�n�;�j;�\I;��(;�;���:�:-V#:��9����U�����'m溘���b0���N�#ol��f��D����j��缻��ɻq�ֻ��
��I����q��-�".�������J �]�$�")�0.-��61��5�(�8��<�
@�IoC�d�F���I���L�5�O�'�R���U���X��R[��^���`���c��Pf�5i�t�k�G�n��_q�5t�:�v�)�y��-|��~�
���ꁼz%��G\��揅��t􇼖(���_������ڌ���th������P��1U�����������G�������ᙼ�+��s��ĸ������b@������Ȣ�����Y��Z���Z���3S���������+r���ծ�V9����������mR��禵�.���$@�������Ǻ�N��XF���  �  �N=,ZN=v�M=�M=�nL=c�K=:K=�pJ=��I=�I=�iH=�G=�G=�eF=f�E=6E=�iD=}�C=�C=5uB=��A=a'A=@=-�?=@)?={>=��====�c<=��;=��:=�C:=ˏ9=��8=�-8=��7=��6=�-6=چ5=(�4=�;4=F�3=�2=lB2=B�1=T�0=6,0=�q/=9�.=��-=!*-=�_,=�+=��*=]�)=�)=�3(=�P'=�g&=�x%=$�$=w�#=�{"=Pi!=�K =�!=X�=!�=�Q=$�=��=�=�z=��=�F=g�=��=45=�u=O�	=��=�=;= ]=�x =/�<�;�<N�<U�<{Q�<�D�< 0�<��<Q��<���<Ȩ�<��<CU�<�*�<���<�տ<⫻<΂�<�Y�<�0�<��<�ئ<���<u�<�<�<y �<��<�|�<�7�<��<O��<L�x<�dp<�g<i�_<B@W<�N<�F<]�><iP6<�!.<t�%<R�<�<BR<�<s��;;�;�p�;q��;�D�;���;"2�;���;�j;�I;�o);E	;���:�:��$:��9_,��-�T�q���y��S��0�z�N���l�� ��\����ҡ������/��dIʻ(�ֻe<�Fﻃ������9��=�c9�G�����I ���$�N�(��-�O#1�b5�a�8��f<�1�?�NLC�p�F���I�w�L�C�O�w�R�R�U��}X��H[�[^�'�`��c��Xf��i���k���n�/xq��;t�R�v�z�y�S|�`�~���������6���k��Ν���͆�@���<0��:e�����8܌����_e���������K��K���`镼�7������IЙ�3���b�������K5��({��O¢����X�����������W��'���d��}���⮼6H��F����
��?e�����	��IR��q����ֺ����uQ���  �  v�N=OWN=j�M=nM=0nL=��K=�K=�rJ=�I=�I=�nH=��G=�G=lF=��E=�E=�oD=��C=e C=yB=��A=^)A=5�@=X�?=�(?=�y>=d�====�_<=�;=��:=�=:=�9=��8=�&8=9y7=��6=�&6=��5=y�4=�64=�3=��2=�?2=z�1=Z�0=�+0=�r/=ʴ.=�-=�--=5d,=8�+=]�*=~�)=?)=1:(=�V'=�m&=�}%=R�$=#=�}"=�j!=L =!=��=�=�N=4�=�{==�=Gt=��=+?=]�=E�=�,=�m=��	=��=q=t5=dX=u =�<K7�<{K�<T�<�R�<�G�<�4�<��<.��<���<���<|��<�b�<�7�<��<w�<���<���<a�<�5�<[	�<�ڦ<Ө�<As�<U9�<&��<��<&t�<n-�<��<ס�<%�x<JFp<��g<qv_<9"W<��N<l�F<Rj><�<6<h.<]�%<��<Ԇ<�O<<���;�;8��;���;�n�;��;�f�;j�;�k;�fJ;�);�z	;���:�z�:ӑ%:σ9U6���xT������)��0�1
O��m�7H���̓�c���毻�g��e�ʻ�0׻�q�#D������('�IJ�C�������I ���$�n�(�O-�1���4�c�8�yO<��?�2C�"zF�\�I��L�)�O���R��U��sX�!B[��
^���`�z�c�@_f�)i���k�"�n��q�?Rt�gw���y��o|� ��ˀ�+��SD��/x������l׆���x6���i�������݌�}��Oc��ૐ������C������ޕ��+���w��/Ù�=��LV��V����垼-���t��ý�����"W��b���! ���[���������΅��M��S��G�������s���ȵ����U`�������⺼��aZ���  �  $�N=mUN=
�M=�M=�mL=��K=CK=tJ=��I=MI=�qH=�G=�G=3pF=%�E=�E=�sD=V�C=E#C=[{B=D�A=�*A=ˀ@=h�?='(?=�x>=��==
==�]<=�;=�:=�9:=ل9=�8=�!8=t7=�6=@"6=d|5=��4=r34=h�3=��2=>2=D�1=��0=�+0=�r/=��.=��-=�/-=�f,=T�+=��*=`�)=T)=G>(=�Z'=q&=��%=��$=��#=;"=tk!=DL =� =�=h�=�L=��=�x=��=/p=U�=P:=.�=��=�'=�h=գ	=�=p=�1=qU=�r =�<p4�<�I�<�S�<S�<xI�<�7�<��<��<��<'��<���<)k�<U@�<��<��<<(��<Xe�<�8�<N�<aۦ<���<�q�<�6�<���<���<}n�<�&�< ߄<1��<��x<|2p<��g<jb_<2W<��N<�F<�[><06<$.<��%<{�<��<�M<�<|��;s$�;��;��;W��;��;���;(�;t_k;ʮJ;D *;��	;���:�Ԓ:? &:�49�����XT�q���խ�s1���0�\,O��.m��a��Lꓻ�%��l	��y�����ʻ�T׻Z���c�w���,��[1��R��I��^��J �߭$�[�(��-��1� �4���8��@<�2�?�O!C�^iF�e�I�E�L�F�O�߭R���U�:mX�>[�a	^���`� �c��cf��/i�^�k���n�j�q��`t��!w�<�y�B�|���QՀ�S���L��(�������p݆����:��m�������ތ�w��Fb��������?��p����ו�7$���o��к�����N��K����ߞ�(���p��ﺢ�8���V���������V^��`���$��a�����l[�������!��3}��kҵ�!��Ci������3꺼�%��`���  �  J�N=�TN=��M=7M=�mL=�K=wK=�tJ=��I=3I=�rH=*�G=G=�qF=~�E=�E=�tD=q�C=G$C=3|B=��A=�*A=�@=u�?=�'?=Mx>=l�==R==�\<=�;=��:=k8:=j�9={�8== 8= s7=v�6=� 6= {5=��4=^24=i�3=��2=|=2=ې1=V�0=�+0=�r/= �.=�-=C0-=�g,=_�+=�*=��)=�)=�?(=�['=Dr&=Á%=ˉ$=b�#=�"=�k!=FL =� =��=�=�K=��=�w=x�=�n=��=�8=o�=Z�=�%=g=C�	=��=(=�0=mT=�q =��<�3�<8I�<�S�<OS�<1J�<%9�<�!�<��<W��<���<>��<�m�<C�<P�<?�<��<��<�f�<�9�<��<�ۦ<P��<q�<�5�<-��<���<Ml�<`$�<a܄<2��<E�x<�+p<��g<�[_<�W<��N<h�F<5W><�+6<�.<9�%<��<��<�M<<���;�(�;��;��;���;:�;���;�!�;Hwk;��J;h6*;��	;7�:��:�N&:��9đ��0QT����A��t8���0�q:O�B?m��j�����-1�����Ҙ���ʻ�a׻���n�Q���f��?5��U��K���^��J �u�$��(��-��	1��4�V�8��;<���?��C��cF�0�I�f�L���O���R���U��jX��<[�	^���`��c�cef��1i� l�h�n���q��et�/'w��y���|��#�^؀�v���O����������߆����<��n��Q���ߌ�h��b��ר��V�t=��q����Օ��!��Pm��!���e���K�������ݞ�.&��~o����������V��!���n��<_�������%��m������^��kñ��$��_���bյ�F$��Pl��ή���캼�'��(b���  �  $�N=mUN=
�M=�M=�mL=��K=CK=tJ=��I=MI=�qH=�G=�G=3pF=%�E=�E=�sD=V�C=E#C=[{B=D�A=�*A=ˀ@=h�?='(?=�x>=��==
==�]<=�;=�:=�9:=ل9=�8=�!8=t7=�6=@"6=d|5=��4=r34=h�3=��2=>2=D�1=��0=�+0=�r/=��.=��-=�/-=�f,=T�+=��*=`�)=T)=H>(=�Z'=q&=��%=�$=��#=="=vk!=GL =� =�=n�=�L=��=�x=��=?p=h�=f:=G�=�=�'=�h=��	=4�=�=&2=�U=�r =��<�4�<#J�<�S�<|S�<�I�<I8�<= �<��<N��<I��<���<.k�<J@�<��<��<���<琷<e�<�8�<�
�<ۦ<!��<eq�<u6�<2��</��<.n�<z&�<�ބ<��<i�x<\2p<��g<�b_<lW<�N<]�F<u\><�06<�.<��%<A�<|�<�N<J<���;�%�;R��;��;5��;��;���;Y�;Y_k;1�J;0*;/�	;���:В::&:�9A˭��fT�Ğ��P��55���0��/O�72m�ic���듻6'���
������
�ʻ�U׻1�㻤d����q���1��R��I�3�{��J ��$�j�(��-��1��4���8��@<�6�?�R!C�`iF�g�I�F�L�G�O��R���U�;mX�>[�b	^���`� �c��cf��/i�^�k���n�j�q��`t��!w�<�y�B�|���QՀ�S���L��(�������p݆����:��m�������ތ�w��Fb��������?��p����ו�7$���o��к�����N��K����ߞ�(���p��ﺢ�8���V���������V^��`���$��a�����l[�������!��3}��kҵ�!��Ci������3꺼�%��`���  �  v�N=OWN=j�M=nM=0nL=��K=�K=�rJ=�I=�I=�nH=��G=�G=lF=��E=�E=�oD=��C=e C=yB=��A=^)A=5�@=X�?=�(?=�y>=d�====�_<=�;=��:=�=:=�9=��8=�&8=9y7=��6=�&6=��5=y�4=�64=�3=��2=�?2=z�1=Z�0=�+0=�r/=ʴ.=�-=�--=5d,=8�+=\�*=~�)=?)=1:(=�V'=�m&=�}%=S�$=Ć#=�}"=�j!=$L =!!=�=�=�N=D�=�{=V�=et=�=U?=��=~�=+-=/n=��	=��=�=�5=�X=�u =��<!8�<NL�<�T�<WS�<SH�<�5�<G�<���<���<��<���<�b�<�7�<q�<+�<��<B��<�`�<!5�<��<�٦<��<�r�<�8�<r��<i��<�s�<�,�<��<���<��x<Fp<��g<�v_<�"W<\�N<F�F<[k><�=6<�.<��%<4�<Z�<.Q<�<w��;��;���;���;^p�;�;�g�;��;Vk;�eJ;��);�w	;H��:�q�:�|%:�$9�i���T�*���x��l&�M�0�4O�B
m�mK���ϓ�.��鯻)j��z�ʻY2׻6s㻍E�V�������'��J�nC������I ���$���(�g-�(1���4�o�8��O<��?�2C�&zF�`�I�
�L�+�O���R��U��sX�"B[��
^���`�z�c�@_f�)i���k�"�n��q�?Rt�gw���y��o|� ��ˀ�+��SD��/x������l׆���x6���i�������݌�}��Oc��ૐ������C������ޕ��+���w��/Ù�=��LV��V����垼-���t��ý�����"W��b���! ���[���������΅��M��S��G�������s���ȵ����U`�������⺼��aZ���  �  �N=,ZN=v�M=�M=�nL=c�K=:K=�pJ=��I=�I=�iH=�G=�G=�eF=f�E=6E=�iD=}�C=�C=5uB=��A=a'A=@=-�?=@)?={>=��====�c<=��;=��:=�C:=ˏ9=��8=�-8=��7=��6=�-6=چ5=(�4=�;4=F�3=�2=lB2=B�1=T�0=5,0=�q/=9�.=��-=!*-=�_,=�+=��*=\�)=�)=�3(=�P'=�g&=�x%=&�$=z�#=�{"=Ui!=�K =�!=c�=/�=�Q=;�=ˀ==�z=2�=G=��=��=�5=Qv=��	=�=M=�;=�]=�y =^�<�<�<FO�<1V�<�R�<�E�<�0�<��<���<v��<&��<��<OU�<m*�<���<տ<R��<��<Y�<�/�<��<�צ<맢<t�<�;�<{��<,��<|�<B7�<O�<׮�<��x<mdp<�g<��_<�@W<��N<D�F<ӂ><R6<�#.<w�%<m�<�<jT<<v��;�
�;Pt�;U��;"G�;K��;N3�;��;��j;`�I;�l);
	;���:ؑ:��$:�.9u����T�u����溘��0�d�N�@�l�%�������֡�.����2��VLʻ��ֻ�>�F�=��������>��9������I �1�$�x�(��-�j#1�w5�r�8��f<�<�?�WLC�w�F���I�{�L�F�O�z�R�T�U��}X��H[�\^�(�`��c��Xf��i���k���n�/xq��;t�R�v�z�y�S|�`�~���������6���k��Ν���͆�@���<0��:e�����8܌����_e���������K��K���`镼�7������IЙ�3���b�������K5��({��O¢����X�����������W��'���d��}���⮼6H��F����
��?e�����	��IR��q����ֺ����uQ���  �  ��N=�]N=ݺM=M=�nL=��K=NK=�mJ=��I=hI=-cH={�G=�G=]F=��E=�	E=�aD=>�C=pC=pB=��A=�$A=i}@=��?=�)?=�|>==�==�==�h<=\�;=��:=}K:=`�9=��8=b78==�7=I�6=k66=��5=j�4=�A4=��3=S�2=E2=Y�1=Y�0=),0=�p/=��.=-�-=y%-=:Z,=X�+=�*=�)=I	)=C+(=tH'=K`&=�q%=�|$=#=^x"=cg!=�J ="=��=ާ=�U=-�=چ=:=�=Z�=!Q=5�=��=_@=܀=��	=/�=�=�B=�c=�~ =	&�<bB�<�R�<W�<Q�<�A�<8*�<J�<[��<���<f��<�n�<�C�<��<^��<"ſ<��<�u�<
O�<(�<���<�Ԧ<1��<�u�<�?�<��<�Ǒ<Ȇ�<LD�<m�<迀<y<Ջp<�h<��_<�gW<kO<u�F<s�><^k6<�8.<&<��<��<JW<:<���;"��;?Q�;F��;A�;�x�;��;So�;�j;�ZI;<�(;��;���:�:J1#:H*9氹�IU�D���.��+��$o0��N��zl�K�Ok�����`o��"뼻zʻ��ֻ���}��"K��Ϭ�5�y.��.�[����J ���$�U)�Y.-��61�5�=�8�.�<�)
@�ToC�l�F���I���L�9�O�*�R���U���X��R[��^���`���c��Pf�6i�t�k�G�n��_q�5t�:�v�)�y��-|��~�
����ꁼz%��G\��揅��t􇼗(���_������ڌ���th������P��1U�����������G�������ᙼ�+��s��ĸ������b@������Ȣ�����Y��Z���Z���3S���������+r���ծ�V9����������mR��禵�.���$@�������Ǻ�N��XF���  �  �O=FaN=R�M=GM=�nL=P�K=�K=�iJ=c�I=�
I=Y[H=��G=�F=�RF=e�E=��D=dXD=��C=�C=�iB=��A=� A=#{@=��?=
*?=/~>=��==�==�m<=Ѻ;=;=[T:=�9=D�8=8B8=%�7=��6={@6=B�5=��4=�H4=K�3=��2=�H2=p�1=1�0=�+0=o/=��.=��-=�-=AS,=@�+=��*=O�)=1�(=-!(=�>'=MW&=�i%=�u$=�y#=Kt"=�d!=�I =-"=`�=��=�Y=��=��=@=v�=��=w\=;�==�L=ڌ=	�	=��=�$=�J=�j=� =E.�<H�<�U�<XW�<�N�<9<�<�!�<�<*��<��<���<wZ�<�.�<��<��<1��<��<&g�<�B�<�<���<�Ц<���<�v�<tC�<��<�Б<���<�R�<��<oӀ<�,y<�p<�Mh<��_<�W<FO<� G<��><��6<�O.<�&<"�<�<%Y<�<�|�;#��;U&�;Zx�;-ζ;-�;S��;��;:Si;��H;/(;m�;\��:��:o�!:I 9����l�U�P਺�{�����@0�X]N�!"l�����*��O��)!��5�����ɻqcֻ)�⻷�� ��O��������"�: �����M �;�$�T)��@-�8N1��95�y9�>�<�2@���C���F��J�M��P��R�8�U�ўX��_[��^�n�`�֍c�If��i���k�n�9Dq���s���v�L`y�b|���~�T����Ձ����VJ��"���괆��釼b ��"Z������ڌ�B!���l���������ya��w������`Z��ϩ��E����?�������ʝ�����M��܎���Т�,���\������$����N��|������f��MǮ�D(������B䲼�<������඼�+���r��a���h����9���  �  �O=�dN=��M=M=qnL=��K=�K=eJ=h�I=bI=�RH=עG=g�F=�GF=�E=��D=�MD=�C=nC=�bB=�A=�A=@x@= �?=�)?=N>=w�==�#==s<=x�;=c;=]:=Q�9=H�8=�M8=��7=1�6=K6=�5=&�4=*P4=-�3=R�2=�K2=-�1=��0=�*0=�l/=a�.=��-=o-=wK,=Cz+=��*=��)=�(=(=4'=aM&=	a%=n$=^s#=�o"=�a!=�G =�!=y�=�=�]=��=u�=�=�=�=sh=��==�Y=��=��	=�=�.=%S=wq=q� =J6�<(M�<�W�<�V�<�J�<�5�<'�<��<R��<s��<r�<UD�<��<���<���<Y��<$y�<�V�<;5�<��<��<�˦<Y��<$w�<�F�<�<�ّ<<b�<�$�<��<~Yy<��p<n~h<y`<��W<�qO<�'G<��><��6<g.<*)&<��<�<^Y<�<�d�;ۯ�;t��;�:�;ք�;�٥;�=�;��;/�h;��G;�r';^=;���:�:q�:6c	9Mⴹ��V����������0��N���k������璻��cή��B��:Yɻ�ֻ]�:G�����v����U��������IR �B�$�� )��U-��h1��Y5�X(9� �<��]@��C�AG�f8J�GM��=P�ES���U���X��n[��$^���`���c��Bf���h���k��nn��'q�j�s�t�v�+6y���{��m~�i}��Z���9����7��p��P����އ�e���T��0���"ڌ��#��.r��1Đ����eo��Ɣ���� o��Ϳ�����HV������yޝ����]��(���Rڢ�����`��٩������zJ������f����Y��R�������s���β�D&��z���ɶ�����^������+黼H-���  �  	O=�gN=<�M={M=�mL=?�K=�K= `J=��I=��H=�IH=ɘG=�F=T<F=��E=0�D=0CD=5�C=��B=0[B=ԹA= A=�t@=,�?=@)?=�>=��==�&==�w<=��;=
;=cf:=D�9=9=�X8=��7=* 7=rU6=J�5=a5=W4=��3=\�2=�N2=q�1=��0=�)0=j/=Z�.=l�-=�-=sC,=q+=��*=��)=��(=�
(=$)'=,C&=�W%=<f$=�l#=yj"=�]!=�E =!=�=�=a=�=�=�#={�=e=#t=U�=�=�f=�=��	==�7=
[=�w=a� =M=�<2Q�<Y�<9U�<_F�<.�<��<���< ��<t��<�\�<�-�<" �<��<��<���<�e�<�E�<�&�<��<��<�Ŧ<��<�v�<�H�<g�<A�<K��<�p�<6�<���<N�y<q<��h<�K`<��W<�O<�MG<�?<��6<�|.<�8&<w�<��<�W<<[I�;��;���;���;�9�;��;6��;@S�;��g;NG;�&;6�;GC�:	�:��:qB9�A���kW��M��*��ɹ���/���M��qk�{N��Ѧ������}���� ɻ��ջ(⻲�����]�Q�����p����p���X �,�$��1)�;l-���1��z5�1N9��<���@�I�C�|<G�VeJ�;qM��cP�V@S�V�V�X��[�\0^���`���c�o>f���h�T�k��Yn��q��s�fhv�/y���{�W@~��f��ʩ��邼�%��`������Շ�L��iP������#ی��'���x��=͐��$���}��ה�/��t���W֘��#��!m��걜��򝼨0���l��O����䢼d#���e��򫦼I���ZG��������6N��﩮�����`������"��ec������� ��K��j���yڻ�|!���  �  �O=qjN=p�M=nM=7lL=��K=/K=[J=��I=.�H=AH=.�G=0�F=�1F=��E=w�D=9D=ȕC=O�B=�SB=ٳA=GA=wq@=��?=7(?=4�>=��==�)==|<=.�;=�;=dn:=H�9=�9=c8=E�7=4
7=�^6=ɳ5=�5=!]4=`�3=�3=�P2=G�1=$�0=�'0=5g/=6�.=�-=-=�;,=h+=��*=E�)=�(= (=�'=�9&=O%=�^$=hf#=`e"=Z!=FC =�=7�=��=�c=(	=��=�*=��==�~=��=�*=:r=0�=&�	=�=8@=b=�}=�� =�B�<4T�<XY�<�R�<`A�<M&�<��<=��<��<&z�<�H�<"�<���<Ⱦ�<a��<�s�< S�<H5�<��<w��<�ު<0��<3��<Wu�<rJ�<��<f�<P��<�}�<�E�<��<V�y<�Aq<M�h<hw`<4X<i�O<pG<W"?<��6< �.<�E&<��<��<�S<�<�,�;�_�;���;ݻ�;&�;>2�;���;���;
g;�\F;�%;&�;M
�:'Ԍ::�p�8�����KX��������ײ�[�/���M�Q'k����Tl��
v��4��,����ȻLmջp����cU��(F����&��k����_���` ���$�LC)���-�6�1�:�5��r9��%=��@� D�LhG��J� �M�O�P��`S�^'V���X��[��<^�'�`�'�c��;f�g�h�?�k�jGn�V�p��s��Fv��x��{�4~�qR������ւ�����R��J���ḋ�[��0M��Ғ���܌��+��.��m֐��0��&����甼�A�������똼�9��ł���Ɯ�,��FB���{������#+���j��ݮ������5E�����G쫼!D��0�������PO�����������N��V���f�w9��߃��nͻ����  �  �O=MlN=-�M=M=�jL=E�K=�	K=bVJ=�I=}�H=q9H=��G=�F=(F=}E=�D=0D=��C=��B=�MB=u�A=�A=6n@=��?='?=�>=��==�+==N<=��;=w#;=u:=��9=9=�k8=��7=�7=�f6=�5=�5=#b4=7�3=f3=R2=��1=u�0=&0=zd/=]�.=#�-=-=�4,=J`+=^�*=!�)=��(=��'=�'=�0&=\G%=�W$=�`#=�`"=�V!=�@ =�=
�=��=
f=y=,�=y0=�="!=��=U�=�4=|=Ǻ=�	=�=G=�g=�=� =G�<V�<�X�<P�<v<�<��<X��<P��<֜�<j�<�6�<G�<g��<L��<h��<�a�<�B�<�&�<P�< �<�֪<.��<O��<�s�<$K�<��<��<���<3��<�R�<��<!�y<�eq<3�h<K�`<^=X<��O<��G<�:?<l�6<y�.<VO&<��<�<�O<#�<o�;�:�;{_�;��;��;c�;�9�;ݣ�;q\f;]�E;�[%;�I;���:�:<w: z�8bɻ�FY�(ک������O�/��M���j����[;��d=��z���\^��6rȻ),ջ�Ỳ��M'��P3�^�����}�
��	��th �j�$�}S)�	�-���1���5���9�I=�e�@�{FD�ʎG�@�J�v�M�\�P�^}S��?V��X�7�[�H^���`�x�c��:f��h�e�k��8n���p�E�s��*v���x�'a{�~�}�A��W����ǂ����G������Ň�����J��˒��ߌ�0��n����ސ�!;��̘��\���R������j����L�������؜�>���Q����������h���h2���o��򱦼�����C�������櫼�;�������鯼�@��j����과c=�����ݷ��*���v���»�����  �  O=�mN=��M=�M=�iL=-�K=�K=�RJ=��I=2�H=�3H=#�G=�F=� F=�uE=��D=)D=�C=!�B=\HB=!�A=aA=zk@=��?=�%?=�>=��==W-==��<=��;=�';=z:=��9=?9=>r8=��7=7=�l6=C�5=i5=�e4=��3=A3=S2=��1=��0=�$0=b/=;�.=4�-=X-=,/,=0Z+=��*=�)=e�(=i�'=�'=E*&=SA%=ZR$=\#=�\"=�S!=�> =j=��=�=�g=�=��=�4=.�=='=q�=��=�;=��=��=��	=�%=DL=l=E�=9� =�I�<�V�<!X�<�M�<8�<��<���<���<���<�]�<')�<���<N��<?��<�u�<�S�<26�<K�<a�<��<Ъ<+��<��<&r�<=K�<� �<��<�<)��<�\�<w(�<f�y<��q<i<�`<�WX<�O<$�G<�L?<��6<٧.<V&<�<D�<^K<M�<���;��;>:�;�W�;�}�;��;��;�d�;�e;�7E; �$;��;�&�:�"�:u-:���8>���i�Y����_����b�/�XcM��j�3؃�G������ƭ��,��@Ȼ��Ի�\ứ_���W%�*��/��F��������;o ���$��`)�W�-�?�1��5���9��d=��@�7dD���G���J���M�i�P�ēS��SV�QY�B�[�#R^�[�`�Жc�;f���h�i�k�.n�f�p�pvs��v�=�x�H{�Y�}�4���x����������>��2����������I��G���ጼ�3�������吼�C��󢓼����^��]�������[��h���&眼�$���]��S����ɡ�����b8��Xt�����������C��8����⫼�5���i௼�5��c����ݳ�J0��8����з����Hm������r���  �  SO=BnN=��M=9M=�hL=ƷK=�K=XPJ=��I=��H=�/H=�{G=��F=	F=�pE=�D=�$D=�C=`�B= EB=`�A=!	A=�i@=y�?=%?=�>=��==,.==�<=��;=,*;=)}:=�9=$#9=\v8=��7=7=hp6=��5=55=h4=��3=_3=�S2=��1=*�0=�#0=�`/=0�.=��-=W�,=�+,=7V+=j~*=��)=��(=��'=#
'=&&=g=%=�N$=Y#=�Z"=�Q!=l= =�=`�=W�=Oh=P=��=i7=d�=�*=��=�=�@=7�=Y�=��	=O)=cO=�n==�=�� =SK�<RW�<LW�<�K�<5�<��<}��<���<���<\U�<d �<D��<���<���<ol�<K�<.�<�<��<��<�˪<ﰦ<В�<q�<EK�<�!�<a��<&ƍ<��<�b�<�/�<m�y<�q<�,i<L�`<hX<
P<�G<_W?<7<!�.<�Y&<�<G�<H<��<4��;�	�;7"�;�;�;>]�;:��;z֓;�;�;e;b�D;�$;��;��:^��:^:�a�8���[5Z��:��l纇���/��PM�ߡj��Ń���������!���8���Ȼ��Ի�?�`F�=�������,�������N���s �8�$�)i)���-���1�f�5��9��u=��	A�QwD���G���J�F�M���P�$�S��_V��Y���[��X^���`�_�c�c;f���h�=�k��'n���p��ks��v�y�x�8{���}��+��q��ش��w���a9��2{���������I�������⌼#6��A���1ꐼ�H��O���1	��g�����7��:e��孛�1�	-��{e������ϡ����R<��Dw����������YC������ૼm2��=����گ��.��Ȃ���ճ��'��y��Rɷ����fg��굻�����  �  I%O=}N=5�M=�&M=�wL=��K=�K=8YJ=m�I=K�H=�.H=�xG=��F=�F=[lE=��D=�%D=��C=��B=^VB=��A=t&A=��@=;�?=Q?=�>='
>=
c==[�<=�<=zf;=$�:=�:= h9=x�8=8=�k7=��6=O6=�o5=��4=�4=�m3=q�2=�2=U1=��0=�/=8/=^J.=w|-=c�,=��+=�+=�,*=�U)=O~(=Q�'=�&=�%=�%=H$=�&#='"=�!=�  =��=�=JX=x=ś=�'=ܥ=�=�z=q�=�=`=��=��
=��=&
=�!=�2=�==:��<���< p�<S�<�)�<���<���<�t�<�,�<s��<���<aX�< �<���<���<���<�o�<�T�<'<�<�$�<��<O�<SТ<���<4��<�S�<�!�<��<���<}�<_C�<�z<��q<�)i</�`<�DX<�O<:kG<�?<J�6<�<.<��%< t<�<ӓ<�<��;f �;���;���;E��;q�;�x�;ZF;��];U�<;�g;A]�:���:�r:x��98(���~5�V<��F�������(:��4X���u�򙉻���v*���������:�λW�ۻ�,�OL�� ����&��o�X���|�0H���#�hu(���,��1��B5�A9�j=���@��MD�.�G��J���M��P��S��&V���X�qA[��]��>`���b��Be�w�g�cYj�x�l�}o�=r�6�t��,w���y�\=|���~������߁����|Z������?ӆ�y���O������ڋ�y'��{���ԏ�Z4��엒������b��}Ŗ��"��py��\ǚ�����H���}��6����֠�* ��d*���W��8����¦�U���E�� ����ݫ��.������ӯ��%��Cw��lȳ����h������]��HQ�������꼼�  �  �$O=�|N=2�M='M=+xL=@�K=zK=`ZJ=ѡI=��H=�0H=�zG=��F=�F=�nE=��D=�'D=��C=_�B=�WB=�A=�'A=y�@=��?=�Q?=,�>=
>=�b==ֹ<=�<=Re;=ú:=n:=if9=��8=@8=	j7=��6=�6=�n5=��4=�4=am3=O�2=�2=zU1=[�0=L�/=A/=�K.=�}-=�,=��+=�+=�.*=X)=t�(=w�'=�&=��%=o%=�$=�'#=("=�!=Q ==�=֟=X=� =�=�&=\�=�=�x=`�=�=�]=k�=��
=��=�=h =�1=�<=b��<P��<rp�<�S�<'+�<���<ں�<_w�<�/�<��<���<�\�<~�<r��<9��<A��<�s�<)X�<m?�<�'�<a�<P�<�Ѣ<Ϭ�<���<�S�<@!�<��<���<�z�<f@�<�z<��q<�!i<t�`<c=X</�O<�dG<~�><p�6<�9.<�%<s<.<3�<�<T%�;��;b��;A��;퓲;Z��;1��;�k;,^;"#=;2�;��:�ڸ:Cs:��9p9��2��~����U�������':��7X��u���������4�����a���[�λ �ۻ�8軽V��� �N��)��p����9|�PF���#��q(���,��1��<5�c:9��=���@��DD�]�G�J�J���M�ٵP�xS�$ V�ɴX�H<[�ռ]�d;`��b��@e��g��Yj���l�so��r�)�t��2w�1�y�XD|��~�R���"ぼ� ��F]������Ԇ����qP�������ً�z&���y��ӏ�*2��B���{���b_���������u��Ú�9���D���y�������Ӡ�T���(���U����������� ���E��_����ޫ��/�������կ��(���z���˳�D���k��칷�e���S�����_켼�  �  Z#O=O|N=K�M=�'M=�yL=?�K=%K=�]J=ѥI=u�H=�5H=]�G=��F=HF=uE=U�D=�-D=<�C=w�B=^\B=��A=�*A=��@=��?=�R?=ɯ>=
>= b==0�<=h<=b;=ʶ:=�:=9a9=;�8=�8=�d7=�6=�6=k5=�4=�4=4l3=��2=72=uV1=��0=��/=/=O.=�-=̱,=�+=�
+=5*=w^)=؆(=��'=��&=<�%=$%=� $=4+#=�*"=�!=� =��=��=@W=J�=r�=8#=%�=�=s=I�=6=�W=P�=$�
=��=Q==0/=%;=���<��<pq�< V�<�.�<���<���<y�<m9�<���<˫�<�i�<�,�<���<��<n��<�<Pb�<tH�<(/�<��<Y��<�բ<B��<���<pS�<��<��<孉<�r�<P7�<��y<
�q<e
i<=�`<"'X<!�O<ySG<��><:�6<�1.<��%<vq<~	<T�<�<�8�;�!�;�;���;��;P��;��;��;�^;�=;��;Jq�:e��:ϕt:���9�@��~[��D~�hݼ�4]�����):��GX�Xv������(���V��9�������ϻ�ۻ:^��v�� ����0��t�(��Zz��A���#��h(���,�1�d+5��&9���<��@��+D�=�G�3�J���M�#�P�bS��V���X��-[��]�/2`�O�b��<e���g��Zj�+�l��o��r�>�t�YCw���y�uY|��~�>����큼.*��^e��ȟ���ن���/R��뒊��؋�$��v��9Ώ�,��������VU��~������Kh�����D���T8��n������Mʠ�1���M!��oP���������������E��Z����᫼=4������5ݯ�n1�������ֳ�Q'��gv��ķ�e���[��@������  �  � O=�zN=)�M=�(M=�{L=H�K=0K=�bJ=�I=��H=>H=d�G=��F=H)F=$E=E�D=n7D=�C=`�B=RcB=��A=�/A=ѓ@=��?=�T?=��>=�	>=q`==m�<=O	<=�\;=A�:=7:=�X9=��8=�8=5\7= �6=�6=&e5=Z�4=�4=!j3=�2=w2=�W1=C�0=��/=v/=}T.=��-==�,=p�+=�+=�>*=rh)=ѐ(=I�'=��&=��%=r%= '$=Y0#=�."=� != =��=l�=�U=|�=P�=�=V�=�=
j=��="=�M=��=#�
=��=��=r= +=98=~�<�~�<�r�<�Y�<�4�<��<���<1��<TH�<��<���<r}�<OA�<m�<8��<���<���<r�<9V�<�:�<g�<���<*ۢ<s��<���<�Q�<��<���<��<zf�<`(�<M�y<�[q<��h<r`<�X<��O<7G<_�><�}6<�$.<G�%<&n<�
<I�<*<W�;�I�;>2�;m�;��;S��;:�;�C�;h:_;�B>;�;s��:���:P�v:r�9�Q���dC}�z���!�����_2:��eX�wBv�Lۉ�XW��⍦��v��2» Fϻ�!ܻ�����+ ����?<��{�Ў�Ox��;���#�YZ(��,���0��5�Y9���<�w�@�;D��[G�|�J��M��xP��?S��U�4�X��[���]�9$`��b��6e���g��]j���l�Гo��/r�)�t��^w���y�Y{|�2�����J���|9���r������^↼����U������e׋�� ���p���Ə��"��1���䓼�E���������}T��̡��0盼�$���[�����������衼���H��B~��X��������E������6櫼�;��t���}鯼�?��ޔ���糼�8������cԷ���(h��a���m����  �  LO=�xN=��M=�)M=�}L=��K= K=�hJ=��I=��H=eHH=ڔG=��F=16F=>�E=�D=�CD=J�C=jC=lB=�A=|5A=S�@=��?=qV?=�>=�>=^==}�<=�<=}U;=�:=1�9=�M9=�8=6�7=�P7=��6=26=2]5=��4=�4=g3=r�2=c2=Y1=ܠ0=��/=�!/=![.=��-=��,=
�+=y+=)K*=Ku)=��(=��'=��&=&=�%=�.$=�6#=�3"=�#!=� =A�=��=;S=v�=��=6=/�=2�=^=��=��=7@=�x=D�
=H�=h�=�=A%=4=y�<�|�<�s�<h]�<J;�<l�<���<'��<O[�<��<���<��<�[�<&�<��<�˿<僚<���<Hg�<?I�<�)�<��<:�<���<τ�<�N�<��<�֍<���<�U�<|�<��y<^+q<�h<�@`<��W<�oO<:G<��><�d6<.<:�%<�h<L<��<46<={�;uz�;ho�;�a�;�X�;)^�;�y�;ʲ�;`;�$?;�|;&H�:�.�:�7y:���9�?&�$���|����4���ش�KE:���X�ǋv����w����צ�,ɴ�c»
�ϻ*xܻ������I ����qM�������Bw�O5�1�#��I(�t�,�9�0���4���8�w�<��S@�j�C�''G�VJ�'`M��HP�QS�e�U�hX�%�Z��]��`�_�b�+1e�~�g��cj�}m�ѥo�WHr�5�t�փw��z���|�0�؀�����M�����������톼#���Z������֋�S���j��������s���ғ��1��Վ���痼�:������I͛����D���x��^���<١�%
��.>���v����������ZF��������E��ޟ�����-S��V�������iP��̞��근�2��y��$�������  �  |O=�uN=Y�M=�)M=�L=8�K="K=�oJ=�I=�I=
TH=١G=��F=�DF="�E=��D=uQD=�C=�C=�uB=�A=�;A=�@=��?=�W?=�>=+>=�Z==C�<=��;=�L;=�:=�9=�@9=�8=W�7=VC7=��6=��5=�S5=-�4=�	4=�b3=�2=�2=�Y1==�0=��/=A'/=Tb.=d�-=%�,=�+=�,+=QY*=�)=K�(=��'=��&=�&=(%=f7$=�=#=�8"=Z'!== =I�=�=�O=/�=_�==�=e�=�O=i�=�=t0=�i=�
=��=l�=�=�=�.=!r�<Ny�<ks�<�`�<�A�<��<���<̭�<�p�<G1�<���<g��<Az�<uD�<��<��<$��< ��<8z�<�X�<,6�<��<��<��<���<&J�<��<ʍ<#��<A�<���<�ry<"�p<8xh<	`<��W<<O<��F<O�><lE6<��-<B�%<�_<D	<c�<B<6��;��;m��;���;[��;S̢;��;�1�;B"a;T&@;�s;r�:�ѽ:�|:���99������E�z�����ӳ��8��e:���X�t�v��K��W㘻*1�� ,��X�»�л��ܻ>J��H���m ����c�Ǖ�����x��0�M�#��8(��,�D�0�g�4���8�6}<��@���C�n�F�?J�E&M��P���R��U��CX�F�Z��q]�-`��b�-e���g�)lj�_m��o��fr�u�?�w�vKz�3�|�|g���	/��3f������˅�a����-���a������׋�����d������
��Qd��󿓼����u��-̗�����i�������t*���`��씠�ȡ�S����3���o�����������H��	���9����R��G�����`j��	Ĳ�!��,l��#�����%J��s����λ�/���  �  �O=rN=6�M=�)M=�L=/�K=�&K=3vJ=S�I=�I=`H=a�G=� G=`TF=ȪE=E=�_D==�C=QC=�B=�A=�AA=U�@=z�?=�X?==�>=�>=dV==�<=��;=�B;=�:=��9=F29=�8=	�7=�47=�6=c�5=�H5=0�4=�4=�]3=��2=
2=�Y1=�0=.�/=�,/=ii.=_�-=��,=�
,=�:+=/h*=P�)=��(=��'=�'=E&=�2%=@$=AD#=v="=C*!=M	 =��=f�=|K=��==�=�x=<�=/@=��=��=6=�X=��
=~�=�=��=�=n(=/i�<t�<�q�<�b�<�G�<t"�<x��<ο�<���<�J�<}�<1��<!��<^d�<i2�<m�<#ڻ<β�<Z��<1h�<�A�<��<d�<��<��<�C�<_�<q��<'s�<*�<��<�7y<<�p<J7h<��_<_W<5O<��F<�f><�!6<�-<[�%<CS<R<��<�K<���;���;��;�	�;4�;R?�;6p�;���;�3b;�5A;uw ;A��:Ɂ�:*
:��9��6t���C�y�aZ��:������:�RY��Ww�P����9������똵�K>ûB}лOPݻ���h���� ��#��}�t����}}�|.���#�>)(��t,���0�P�4���8�eJ<�D�?�[C���F�n�I�y�L���O�ǯR��oU�LX���Z��[]�!�_��b��+e�1�g��xj��&m�?�o���r��8u���w���z�,}������'L��1���
���(������:���j�����ً�&���_��̬�������T����������[��n���L����J������Ҝ����H�����Զ����)��ni������P���oL��m���J��ha�� î��$�����Q಼8��֊��2ض�� ��3d��]���;⻼����  �  ZO=zmN=X�M=h(M=d�L=k�K=�*K=
|J=�I=�I=�kH=|�G=�G=ocF=�E=�E=nD=�C={)C=��B=g�A=[GA=�@=Q @=�X?=��>=c>=bQ==K�<=��;=8;=Ԅ:=�9=a#9=nv8=c�7=@%7=ŀ6=e�5=X=5=��4=*�3=�W3=��2=�2=NY1=�0=��/=1/=�o.=��-=&�,={,=�G+=�v*=Q�)=��(=�'=�'=!)&=�<%=8H$=QJ#=�A"=s,!=�	 =�=(�=`F=��=v=��=�k=��=!0=��=�=�=�G=�{
= �=`�=��=�=i!=�^�<wm�<�n�<Qc�<GL�<�*�<�<���<���<�c�<F*�<&��<W��<���<jP�<` �<5�<uȷ<'��< v�<L�<B�<N�<_��<�|�<�;�<|��<e��<_�<&�<rƀ<V�x<�rp<�g<
�_<�W<��N<�|F<G9><��5<��-<��%<
D<m�<0�<
S<���;U�;�7�;[�;���;��;:�;\:�;)@c;�=B;[t!;�� ;J#�:��:�5:9;R7����x�� �����%����:��wY���w�ߊ����t����	��x�û��л)�ݻ:"����� �H�˚�߽�������/�1�#��(�=a,�ԃ0���4�l`8�a<�g�?� C�goF��I�Z�L���O�~~R�[EU���W�åZ�kH]� �_�҈b�U-e�~�g��j�[=m�(�o�;�r�eu��x�A�z��U}���31��"j������ʄ���������H��8u�����p܋�S���\������v���uF��k����JB�������ᘼ�+���r��G�������+1�� l��ڦ���⢼�!���d��T���L����Q��C�������q��׮�<������l����V��#�������=����'�������"0���  �  �O=�hN=��M=�&M=,�L=��K=�-K=��J=��I=5$I=�uH=S�G=�G="qF=��E=� E=�zD=��C=j3C=��B=��A=�KA=��@=V@=lX?=��>=��==L==K�<=,�;=�-;=�x:=��9=09=�g8=��7=�7=s6=��5=J25=7�4=p�3=�Q3=E�2=�2=�W1=W�0=��/=�4/=Iu.=��-=6�,=8!,=T+=��*=��)=M�(=0�'=�'=�3&=�E%=5O$=qO#=�D"=�-!=C	 =
�=f�=�@=��=*m=�=u_=��=� =]r=h�=��=�7=\l
=�=�=�=�=A=�S�<�e�<�j�<�b�<O�<�1�<��<[��<:��<�y�<�C�<i�<���<ޟ�<�k�<�9�<�	�<�۷<���<	��<%T�<�#�<��<L��<[w�<�2�< �<K��<UK�<���< ��<��x<@5p<.�g<{E_<��V<��N<�IF<><a�5<X�-<m%<?3<f�<�<�V<H��;�8�;o�;f��;ش;^�;~[�;z��;�3d;/C;�Z";��;���:j(�:;:��7���4x���������;�R�Y�NJx��)��D왻v^��!u��V%Ļ�fѻ�4޻*���k��V� ��k�����������a3���#�(��Q,��l0��e4�;8�]�;��|?�y�B��7F�FfI��xL��pO�5RR��U�d�W�ƎZ��8]���_���b��1e�2�g�˘j��Tm�Ap��r���u�hFx�l�z���}�A���N����������ㄼ�
���0��W��:���ȭ��ዼ����Z������됼9:������g۔��+��(z���Ƙ�,���V������ܝ�2���Z������آ����a��h�������)X��Ҷ�����Ӂ���ꮼ�R��O���1��t���ǵ�x���Y������EӺ�l
���@���  �  ��N=�cN=��M=�$M=f�L=f�K=�/K=��J=(�I=-+I=d~H=(�G=�&G=�|F=��E=
,E=��D=�C=�;C=��B=��A=,OA=d�@=�@=\W?=)�>=��==G==ԑ<=[�;=|$;=hn:=0�9=�9=�Z8=k�7=�	7=
g6=��5=r(5=��4=a�3= L3=��2=�2=SV1=��0=��/=J7/=vy.=ʷ-=��,= *,=7^+=ʎ*={�)=��(=7(=%'=�<&=�L%=�T$=YS#=�F"=g.!=X =��=��=�;=�=e=v�=kT=H�=h=&d=ɬ=W�=�)=_
=׎=�=��=��=�=�I�<d^�<�e�<�`�<�P�<r6�<(�<M��<���<R��<�X�<v#�<���<ѷ�<���<�N�<>�<�<��<��<Z�<�&�<y�<\��<�q�<*�<Kݑ<���<�9�<#�<���<��x<m�o<�~g<�_<2�V<o_N<DF<��=<ȴ5<T�-<W%<�"<��<@�<@X<p	�;<V�;y��;+��;� �;�h�;���;X�;e;�C;M#;�h;L��:,�:�:�G�7�H�3�w��������� 2��M;�m-Z�g�x�nm���:��Q���1Զ���Ļv�ѻ��޻�껨����3�����������ϙ��8��#��(�F,�-[0�pM4��8���;�rS?�d�B��F�27I�JKL�CGO�o-R�� U���W�}Z�x-]�T�_�W�b��7e���g�\�j��jm��/p�N�r�^�u��qx�F!{�U�}�_)���h��џ��σ�Z���m���@��Od������~���.拼6���Z��˝���吼�0���}��V˔����e�����������?������ȝ��
��cL�������Т�b���_������q���^�������&������$���g���α��1��ʍ��"⵼?.��yr��ǯ���纼P���O���  �  ��N=�_N=��M=�"M=~L=��K=S1K=+�J=�I=O0I=��H=��G=/G=^�F=��E=�4E=��D=K�C=�AC=v�B=E�A=qQA=��@=�@=:V?=��>=��==�B==��<=�;=#;=!f:=	�9=��8=�P8=G�7= 7=�]6=%�5=� 5=��4=��3=qG3=L�2=6�1=�T1=e�0=|�/=9/=e|.=�-=�,=�0,=�e+=�*=�)=o�(=}(=�,'=1C&=@R%=�X$=V#=hH"=�.!=R =��=n�=~7=��=�^=��=�K=��=�=(Y={�=�=�=�T
=I�=|�=��=_�=U=%A�<X�<�a�<_�<XQ�<�9�<#�<��<��<>��<uh�<�4�<���<���<ғ�<^�<*�<���<ĳ<s��<	^�<2(�<��<Z��<Rl�<�"�<�ӑ<���<>+�<�Մ<J��<�fx<��o<)Tg<^�^<�V<�8N<<�E<c�=<�5<�o-<�D%<<m�<u�<UX<��;k�;��;��;�V�;���;� �;�a�;I�e;�D;7�#;'�;��:3�:v:z�7�1�k�w�����7���-X�c�;�uvZ�Ay������x������s����Ļ�һ��޻1뻽���/�2��{�����8��e��c>�o�#��(�~>,��N0��;4��8���;�M4?���B�Q�E��I�N)L��'O��R�)�T��W�{pZ��%]�O�_�"�b��=e���g�|�j�(}m�=Fp��s���u�J�x��F{���}��=��}��U����ჼ	��P,��mM��o��J�������ꋼ���[��ʛ��Pᐼ�)��Ft��z����
��!U������發b.���t�����������A��녡�~ˢ�e��B_��=�����qd���Ǫ�b0��m���,
���v���౼�D������h���6B���������������*���[���  �  I�N=)]N=��M=2!M=�~L=��K=�1K=��J=M�I=m3I=��H=�G=(4G=ŊF=�E=�9E=��D=��C=cEC=e�B=a�A=�RA=��@=^@=ZU?=z�>=��==@==-�<=��;=p;=�`:=A�9=��8=!J8=ʟ7=��6=�W6=��5=�5=�4=��3=gD3=�2=p�1=�S1=�0=��/=�9/=%~.=��-=w�,=�4,=�j+=?�*=��)=��(=�(=T1'=4G&=�U%=j[$=�W#=&I"=�.!=� =�=I�=�4=6�=]Z=��=2F=s�=M=%R=I�=��=�=N
=7=�=/�=H�=�
=�;�<�S�<_�<�]�<gQ�<�;�<��<s��<��<̢�<nr�<�?�<�
�<���<���<3h�<r2�<���<Yɳ<,��<�_�<�(�<��<��<�h�<��<B͑<�x�<"�</˄<�v�<bMx<��o<�8g<�^<1lV<k N<��E<��=<��5<va-<-9%</<)�<�<�W<�;�w�;y��;�#�;Fx�;�Ϥ;!-�;=��;��e;$�D;�$;�=;~?�:*^�:�:��7���4ww��
�����r�B�;���Z��Py��Ƌ�����
(��N��Ż�Kһk߻m_��.��4C�������'�H�����B��#�w
(�k:,�CG0�14��7���;�!?�f�B�G�E���H�"L��O�/R�+�T�W�W��hZ��!]�a�_���b��Ae�R�g���j��m��Tp�!s���u�S�x��^{��~��J������ǿ��<탼����5���U�� v������{����틼�!���[������ސ��%���n��5������-K������ܙ��#��>j��h���	���j;��0���KȢ����=_�������	��8h���̪��6��/���*��2����뱼�P������h��O��摸�"͹�D���3���c���  �  $�N=4\N=�M=� M=|~L=��K=-2K=)�J=�I=�4I=�H=��G=�5G=��F=��E=�;E=<�D=(�C=�FC=e�B=
�A=3SA=$�@=W@=U?=ߥ>=��==?==��<=��;=�;=�^:=>�9=��8=�G8=��7=��6=�U6=��5=�5=~4=��3=QC3=�2=��1=S1=��0=��/=4:/=�~.=h�-=��,=56,=l+=��*=F�)=��(=X(=�2'=�H&=�V%=5\$=2X#=eI"=�.!=P =��={�=�3=��=�X=E�=PD=b�= =�O=�=z�=S=�K
=2}=C�=��=��=�	=�9�<�R�<(^�<�]�<�Q�<R<�<��<]��<���<���<�u�<C�<��<���<��<_k�<F5�<���<�ʳ<5��<{`�<�(�<-�<嬞<9g�<��<�ʑ<�u�<��<hǄ<pr�<�Dx<�o<�/g<ѿ^<hcV<*N<J�E<�=<�5<�\-<F5%<H	<�<�<2X<��;�|�;,��;�-�;f��;�ݤ;2<�;���;�f;gE;�$$;IX;�n�:D��:I�:74�7��sw����i-��b~�Ǻ;�ǹZ�4gy��Ӌ�ɯ��8��:_���Ż ]һ�%߻�o��=��J�������]�������[D�v�#�#
(�9,��D0��-4�'�7�F�;��?�mB��E���H�!L�O�{�Q�9�T��W��fZ�m ]��_�>�b��Ce�� h�.�j�N�m�Zp�'s�m�u�ѱx��f{��~��N��]���Ă�D񃼙��$9���X��wx��	����&a"���[��Ú��
ސ�{$���l����������G��t���nؙ�����f��R���I�$9�����IǢ�q��,_��
����
���i���Ϊ��8��䦭�@��Ä���ﱼU��񲴼����S�����ѹ�����6���f���  �  I�N=)]N=��M=2!M=�~L=��K=�1K=��J=M�I=m3I=��H=�G=(4G=ŊF=�E=�9E=��D=��C=cEC=e�B=a�A=�RA=��@=^@=ZU?=z�>=��==@==-�<=��;=p;=�`:=A�9=��8=!J8=ʟ7=��6=�W6=��5=�5=�4=��3=gD3=�2=p�1=�S1=�0=��/=�9/=%~.=��-=w�,=�4,=�j+=?�*=��)=��(=�(=U1'=4G&=�U%=k[$=�W#=(I"=�.!=� =�=O�=�4=@�=jZ=�=EF=��=h=ER=o�=�=�=BN
=q=I�=q�=��=1=E<�<�T�<�_�<M^�<�Q�<�;�<-�<���<p��<��<�r�<�?�<�
�<���<l��<�g�<,2�<:��<�ȳ<���<�_�<((�<1�<���<?h�<2�<�̑<gx�<�!�<�ʄ<Rv�<Mx<��o<�8g<7�^<lV<� N<v�E<N�=<p�5<`b-<):%<7<7�<�<�X<�;�y�;��;%�;oy�;�Ф;�-�;��;s�e;[�D;S$;�;;8:�:�W�:G�:M��79���w�����%���w�)�;���Z�&Uy�ɋ�����)���O���	ŻXMһ�߻~`��/���C�T��
��d�{�����B��#��
(�}:,�RG0�!14��7� �;�!?�k�B�J�E���H�$L��O�0R�,�T�X�W��hZ��!]�a�_���b��Ae�R�g���j�	�m��Tp�!s���u�T�x��^{��~��J������ǿ��<탼����5���U�� v������{����틼�!���[������ސ��%���n��5������-K������ܙ��#��>j��h���	���j;��0���KȢ����=_�������	��8h���̪��6��/���*��2����뱼�P������h��O��摸�"͹�D���3���c���  �  ��N=�_N=��M=�"M=~L=��K=S1K=+�J=�I=O0I=��H=��G=/G=^�F=��E=�4E=��D=K�C=�AC=v�B=E�A=qQA=��@=�@=:V?=��>=��==�B==��<=�;=#;=!f:=	�9=��8=�P8=G�7= 7=�]6=%�5=� 5=��4=��3=qG3=L�2=6�1=�T1=e�0=|�/=9/=e|.=�-=�,=�0,=�e+=�*=�)=o�(=}(=�,'=2C&=AR%=�X$=V#=lH"=�.!=X =��=z�=�7=��=�^=��=�K=ʯ=	=fY=á=a�=�=�T
=��=��=�=��=�=?B�<0Y�<�b�<!`�<YR�<�:�<��<���<���<���<�h�<�4�<���<���<���<^�<�)�<���<Só<���<]�<;'�<��<Z��<Wk�<�!�<�ґ<��<�*�<3Մ<؁�<	fx<`�o<&Tg<��^<��V<�9N<`�E<��=<��5<�q-<�F%< <x�<�<SZ<��;�n�;��;��;5Y�;C��;��;ub�;�e;|�D;t�#;1�;���:�ރ:9�:`*�7v񹀲w����R���a�ێ;��Z�y�ۧ���|��a����!����ĻFһW�޻*3뻆���0�ئ������������>���#��(��>,��N0��;4�8���;�Y4?���B�X�E��I�S)L��'O��R�+�T��W�|pZ��%]�P�_�#�b��=e���g�}�j�(}m�=Fp��s���u�J�x��F{���}��=��}��U����ჼ	��P,��mM��o��J�������ꋼ���[��ʛ��Pᐼ�)��Ft��z����
��!U������發b.���t�����������A��녡�~ˢ�e��B_��=�����qd���Ǫ�b0��m���,
���v���౼�D������h���6B���������������*���[���  �  ��N=�cN=��M=�$M=f�L=f�K=�/K=��J=(�I=-+I=d~H=(�G=�&G=�|F=��E=
,E=��D=�C=�;C=��B=��A=,OA=d�@=�@=\W?=)�>=��==G==ԑ<=[�;=|$;=hn:=0�9=�9=�Z8=k�7=�	7=
g6=��5=r(5=��4=`�3= L3=��2=�2=SV1=��0=��/=J7/=vy.=ʷ-=��,= *,=7^+=ʎ*={�)=��(=8(=%'=�<&=�L%=�T$=\S#=�F"=n.!=b =��=��=�;=4�=4e=��=�T=��=�=~d=.�=��=*=�_
=u�=��=<�=��=o=9K�<�_�<yg�<eb�<R�<�7�<X�<W��<���<��<Y�<�#�<���<���<H��<N�<~�<.�<���<䉯<�X�<J%�<�<�<*p�<�(�<ܑ<���<�8�<R�<��<��x<��o<�~g<$_<�V<�`N<�F<��=<	�5<Ԉ-<�Y%<�%<��<"�<[<��;8[�;���;
��;�#�;/k�;D��;�;�e;��C;e#;Nc;��:��:,�:��7K��<�w�=�������?�Y[;�v:Z���x�\s��@��s����ض�ߌĻ<�ѻ �޻���/���*���w�������A��59�5�#��(�NF,�T[0��M4��8���;��S?�q�B��F�:7I�PKL�HGO�s-R�� U���W�}Z�z-]�U�_�X�b��7e���g�\�j��jm��/p�N�r�_�u��qx�F!{�U�}�_)���h��џ��σ�Z���m���@��Od������~���.拼6���Z��˝���吼�0���}��V˔����e�����������?������ȝ��
��cL�������Т�b���_������q���^�������&������$���g���α��1��ʍ��"⵼?.��yr��ǯ���纼P���O���  �  �O=�hN=��M=�&M=,�L=��K=�-K=��J=��I=5$I=�uH=S�G=�G="qF=��E=� E=�zD=��C=j3C=��B=��A=�KA=��@=V@=lX?=��>=��==L==K�<=,�;=�-;=�x:=��9=09=�g8=��7=�7=s6=��5=J25=7�4=p�3=�Q3=E�2=�2=�W1=W�0=��/=�4/=Iu.=��-=6�,=8!,=T+=��*=��)=M�(=0�'=�'=�3&=�E%=8O$=uO#=�D"=�-!=N	 =�=z�=A=��=Tm=C�=�_=��=5!=�r=�=z�=X8=m
=ϛ=��=��=�=1=�U�<�g�<tl�<rd�<�P�<@3�<B�<���<K��<�z�<D�<��<���<���<Mk�<�8�<��<^ڷ<Q��<���<�R�<&"�<��<���<�u�<1�<{�<뙍<#J�<���<;��<s�x<�4p<)�g<�E_<��V<,�N<�KF<�><#�5<g�-<`p%<�6<��<��<[Z<���;�>�;�t�;$��;�۴;P�;m]�;Y��;Z3d;g,C;�U";�;��:*�:%
:�7�7^��7sx��!�����A�A;�I�Y��Yx�1��󙻾d���z���*Ļ�kѻ�8޻����n���� ��l���N��W������3��#�h(��Q,�
m0��e4�;;8�v�;��|?���B��7F�PfI��xL��pO�:RR��U�g�W�ȎZ��8]���_���b��1e�3�g�˘j��Tm�Ap��r���u�hFx�l�z���}�A���N����������ㄼ�
���0��W��:���ȭ��ዼ����Z������됼9:������g۔��+��(z���Ƙ�,���V������ܝ�2���Z������آ����a��h�������)X��Ҷ�����Ӂ���ꮼ�R��O���1��t���ǵ�x���Y������EӺ�l
���@���  �  ZO=zmN=X�M=h(M=d�L=k�K=�*K=
|J=�I=�I=�kH=|�G=�G=ocF=�E=�E=nD=�C={)C=��B=g�A=[GA=�@=Q @=�X?=��>=c>=bQ==K�<=��;=8;=Ԅ:=�9=a#9=nv8=c�7=@%7=ŀ6=e�5=X=5=��4=*�3=�W3=��2=�2=MY1=
�0=��/=1/=�o.=��-=&�,=z,=�G+=�v*=Q�)=��(=�'=�'=")&=�<%=;H$=UJ#=�A"=},!=�	 =.�=?�=~F=�=Ev=��=2l=��=�0=�=��=;=�H=Q|
=ة=H�=��=�=u"=�`�<�o�<�p�<\e�<7N�<�,�<��<��<���<d�<�*�<���<m��<M��<�O�<��</�<3Ƿ<���<|t�<@J�<c�<a�<p��<�z�<�9�<��<ܩ�<�]�<	�<�ŀ<(�x<rp<�g<��_<!!W<d�N<�~F<�;><��5<h�-<`�%<�G<^ <"�<�V<���;#�;�=�;Q`�;��;_��;b�;T;�;�?c;;B;o!;� ;��:�Ԁ:8�:Z
C7�����#y��D��������8�:���Y���w�犻����v�����?�û	�л��ݻ6&�A���� �ZI�ڛ�¾�J�����0���#�(��a,��0�߃4��`8�}<�}�?�+ C�uoF��I�b�L���O��~R�_EU���W�ťZ�mH]��_�Ԉb�V-e��g��j�\=m�(�o�<�r�eu��x�A�z��U}���31��"j������ʄ���������H��8u�����p܋�S���\������v���uF��k����JB�������ᘼ�+���r��G�������+1�� l��ڦ���⢼�!���d��T���L����Q��C�������q��׮�<������l����V��#�������=����'�������"0���  �  �O=rN=6�M=�)M=�L=/�K=�&K=3vJ=S�I=�I=`H=a�G=� G=`TF=ȪE=E=�_D==�C=QC=�B=�A=�AA=U�@=z�?=�X?==�>=�>=dV==�<=��;=�B;=�:=��9=F29=�8=	�7=�47=�6=c�5=�H5=0�4=�4=�]3=��2=
2=�Y1=�0=-�/=�,/=ii.=^�-=��,=�
,=�:+=/h*=P�)=��(=��'=�'=F&=�2%="@$=FD#=}="=M*!=Z	 =��=~�=�K=	�=B=�=	y=��=�@=1�=K�=�=�Y=O�
=]�=�=��=�=�)=dk�<Pv�<t�<�d�<�I�<P$�<&��<G��<�<�K�<,�<���<8��<'d�<�1�<��<ٻ<���<Ջ�<~f�<@�<��<f�<��<�<�A�<���<۹�<�q�<�(�<
�<�6y<��p<C7h<i�_<E`W<�O<B�F<�i><%6<��-<)�%<@W<g<԰<�O<5��;���;b��;C�;�#�;�B�;rr�;���;;3b;x2A;�q ;e��:em�:�~:�X�9u�6�T��sz����n���6����:��1Y�]iw������A��������FDû��лUݻ�������o� �%��~�_��ԧ�~� /�*�#��)(�u,��0�}�4�ʊ8��J<�[�?�[C���F�y�I���L���O�̯R��oU�OX���Z��[]�#�_��b��+e�2�g��xj��&m�@�o�r��8u���w���z�,}������'L��1���
���(������:���j�����ً�&���_��̬�������T����������[��n���L����J������Ҝ����H�����Զ����)��ni������P���oL��m���J��ha�� î��$�����Q಼8��֊��2ض�� ��3d��]���;⻼����  �  |O=�uN=Y�M=�)M=�L=8�K="K=�oJ=�I=�I=
TH=١G=��F=�DF="�E=��D=uQD=�C=�C=�uB=�A=�;A=�@=��?=�W?=�>=+>=�Z==C�<=��;=�L;=�:=�9=�@9=�8=W�7=VC7=��6=��5=�S5=-�4=�	4=�b3=�2=�2=�Y1==�0=��/=A'/=Tb.=d�-=%�,=�+=�,+=QY*=�)=K�(=��'=��&=�&=
(%=j7$=�=#=�8"=c'!=K =[�=��=�O=U�=��=T=f�=��=@P=�=��=1=Cj=ܛ
=f�=T�=�==�/=Bt�<q{�<�u�<�b�<�C�<��<5��<7��<�q�<62�<���<ȴ�<Wz�<AD�<
�<��<��<ݚ�<�x�<>W�<f4�<��<��<��<ځ�<UH�<0
�<�ȍ<΄�< @�<���<�qy<��p<2xh<�`<��W<�=O<��F<��><~H6<)�-<�%<�c<5<T�<�E<���;N��;���;��;���;�Ϣ;��;�2�;�!a;d#@;�n;�:㽽:0�{:�b�9�gJ��j�� %{��һ��������ew:���X���v��S���꘻*8��e2���»�л��ܻ;N�=L��o �&��d����@��yy�'1���#��8(�P�,�{�0���4�ڶ8�Q}<��@���C�{�F�JJ�M&M��P���R��U��CX�H�Z��q]�.`��b�-e���g�)lj�_m��o��fr�u�?�w�vKz�3�|�|g���	/��3f������˅�a����-���a������׋�����d������
��Qd��󿓼����u��-̗�����i�������t*���`��씠�ȡ�S����3���o�����������H��	���9����R��G�����`j��	Ĳ�!��,l��#�����%J��s����λ�/���  �  LO=�xN=��M=�)M=�}L=��K= K=�hJ=��I=��H=eHH=ڔG=��F=16F=>�E=�D=�CD=J�C=jC=lB=�A=|5A=S�@=��?=qV?=�>=�>=^==}�<=�<=}U;=�:=1�9=�M9=�8=6�7=�P7=��6=26=2]5=��4=�4=g3=r�2=c2= Y1=ܠ0=��/=�!/= [.=��-=��,=	�+=y+=(K*=Ku)=��(=��'=��&=&=�%=�.$=�6#=�3"=$!=� =Q�=��=VS=��=Î=k=o�=��=v^=�=D�=�@=fy=��
=	�=8�=�=*&=
5=�z�<�~�<tu�<<_�<=�<	�<��<n��<`\�<|�<>��<u��<\�<�%�<���<K˿<��<؄�<�e�<�G�<W(�<�<�ߢ<�<��<"M�<��<TՍ<p��<�T�<��<w�y<�*q<�h<A`<��W<#qO<2G<�><Ug6<�.<��%<l<�<�<�9<ҁ�;���;�t�;of�;�\�;a�;�{�;���;`;�!?;�w;g:�:�:y:��9��3�2���]S|�m5��I��p���U:���X��v����B���ަ��δ�0h»��ϻ@|ܻ������dJ ����dN����Z���w��5���#��I(���,�j�0��4���8���<��S@�y�C�4'G�VJ�/`M��HP�VS�i�U�!hX�'�Z��]��`�`�b�,1e�~�g��cj�}m�ҥo�WHr�5�t�փw��z���|�0�؀�����M�����������톼#���Z������֋�S���j��������s���ғ��1��Վ���痼�:������I͛����D���x��^���<١�%
��.>���v����������ZF��������E��ޟ�����-S��V�������iP��̞��근�2��y��$�������  �  � O=�zN=)�M=�(M=�{L=H�K=0K=�bJ=�I=��H=>H=d�G=��F=H)F=$E=E�D=n7D=�C=`�B=RcB=��A=�/A=ѓ@=��?=�T?=��>=�	>=q`==m�<=O	<=�\;=A�:=7:=�X9=��8=�8=5\7= �6=�6=&e5=Z�4=�4=!j3=�2=v2=�W1=C�0=��/=u/=}T.=��-=<�,=o�+=�+=�>*=rh)=ѐ(=J�'=��&=��%=t%='$=]0#=�."=� !=� =��=}�=�U=��=s�=�=��="=Uj=��=�=N=�=��
=��=+�='=�+=�8=��<u��<:t�<[�<6�<��<��<<��<3I�<��<��<�}�<_A�<G�<���<��<鏻<1q�<&U�<�9�<�<���<�٢<	��<#��<mP�<��<tߍ<��<�e�<�'�<q�y<\[q<��h<�r`<�X<ޛO<�8G<R�>< �6<O'.<��%<�p<�<+�<�,<v\�;�N�;�6�;M�;��;���;��;8D�;:_;�@>;�;:��:��:��v:"�9�ᔷMG�qv}������<��&���?:��rX��Nv�9ቻ�\�����_{��m»�Iϻ�$ܻ���v���), ����=��|�Z���x��;��#��Z(���,���0�5�s9���<���@�GD��[G���J��M��xP��?S��U�6�X��[���]�:$`���b��6e���g��]j���l�Гo��/r�*�t��^w���y�Y{|�2�����J���|9���r������^↼����U������e׋�� ���p���Ə��"��1���䓼�E���������}T��̡��0盼�$���[�����������衼���H��B~��X��������E������6櫼�;��t���}鯼�?��ޔ���糼�8������cԷ���(h��a���m����  �  Z#O=O|N=K�M=�'M=�yL=?�K=%K=�]J=ѥI=u�H=�5H=]�G=��F=HF=uE=U�D=�-D=<�C=w�B=^\B=��A=�*A=��@=��?=�R?=ɯ>=
>= b==0�<=h<=b;=ʶ:=�:=9a9=;�8=�8=�d7=�6=�6=k5=�4=�4=4l3=��2=72=uV1=��0=��/=/=O.=�-=̱,=�+=�
+=5*=w^)=؆(=��'=��&==�%=%%=� $=6+#=�*"=�!=� =��=˟=OW=]�=��=V#=J�==Cs=��=~=�W=��=��
=]�=�=�=�/=�;=���<��<�r�</W�<�/�<���<[��<6��<:�<h��<#��<�i�<�,�<���<���<��<�~�<�a�<�G�<O.�<��<a��<�Ԣ<B��<���<R�<�<��<4��<cr�<�6�<T�y<�q<b
i<��`<�'X< �O<�TG<V�><ё6<�3.<y�%<us<�<^�<�!<�<�;�%�;I�;J��;W��;��;5��;��;Չ^;n�=; �;Yi�:1��:>}t:+��9&0ķ�}��h~�$�Mp��x���2:�QX�0v�溉��,��:Z��m<������Wϻn�ۻJ`軬x��� �@���0�Lu�����z�B�$�#��h(���,�11�{+5��&9��<���@��+D�D�G�9�J���M�'�P�bS��V���X��-[��]�/2`�P�b��<e���g��Zj�+�l��o��r�>�t�YCw���y�uY|��~�>����큼.*��^e��ȟ���ن���/R��뒊��؋�$��v��9Ώ�,��������VU��~������Kh�����D���T8��n������Mʠ�1���M!��oP���������������E��Z����᫼=4������5ݯ�n1�������ֳ�Q'��gv��ķ�e���[��@������  �  �$O=�|N=2�M='M=+xL=@�K=zK=`ZJ=ѡI=��H=�0H=�zG=��F=�F=�nE=��D=�'D=��C=_�B=�WB=�A=�'A=y�@=��?=�Q?=,�>=
>=�b==ֹ<=�<=Re;=ú:=n:=if9=��8=@8=	j7=��6=�6=�n5=��4=�4=am3=O�2=�2=zU1=[�0=L�/=A/=�K.=�}-=�,=��+=�+=�.*=X)=t�(=w�'=�&=��%=p%=�$=�'#=("=�!=U =B�=ܟ=X=� = �=�&=p�=�=�x=��=�=^=��=��
=�=�=� =2="==��<��<q�<aT�<�+�<��<I��<�w�<40�<T��<$��<�\�<��<d��<��<��<�s�<�W�<?�<'�<��<��<uѢ<K��<!��<bS�<� �<:�<d��<4z�<+@�<�z<k�q<�!i<��`<�=X<��O<yeG<4�><C�6<�:.<�%<t<=	<B�<�<L'�;~
�;��;���;��;<��;Ŋ�;yl;
^;Y"=;Ë;̠�:}ո:P6s:�h�9�B�qD���\)��8������u,:�}<X���u�%�������6����������λY�ۻ:軪W�� ����K)�0q����c|�rF��#�r(���,��1��<5�l:9��=���@��DD�`�G�L�J���M�۵P�xS�% V�ʴX�I<[�ռ]�e;`��b��@e��g��Yj���l�so��r�*�t��2w�1�y�XD|��~�R���"ぼ� ��F]������Ԇ����qP�������ً�z&���y��ӏ�*2��B���{���b_���������u��Ú�9���D���y�������Ӡ�T���(���U����������� ���E��_����ޫ��/�������կ��(���z���˳�D���k��칷�e���S�����_켼�  �  �4O=��N=��M=�8M=ȈL=��K=$K=$bJ=ߤI=��H=*H=�oG=H�F=1
F=�`E=i�D=� D=>�C=��B=#eB=�A=DA=��@=�@=?=k�>=l>>=��==�<=iK<=��;=H�:=GU:=��9=y9=tb8=n�7=�7=�p6=(�5=5%5=�~4=��3=[,3=Z~2=��1=�1=�U0=]�/=a�.=��-=;+-=�X,=��+=ղ*=�)=[)=@(=�n'=�&=g�%==�$=��#=�#=N"=3� =j�=��=�V=� =#�=�%=�=�=p=��=O	=�C=rs=a�=��	=��=��=��=��=Y��<���<M��<�d�<''�<)��<���<4,�<���<xk�<��<���<l�<j*�<v��<�ɿ<!��<ō�<�w�<�b�<�K�<1�<��<��<E��</��<�Q�<d�</ى<���<�Z�<�4z</�q<�.i<*�`<'X<�O<�)G<��><y>6<��-<m^%<p�<(n<��<�P<�Y�;���;ԁ�;#�;���;c&�;��;��w;��U;��4;÷;��:䷦:�N:;E�9u�/�k�(�&w����к;M��2&��D�kgc��ŀ�.���i>��ӕ��E���p[ȻI�ջ>�⻳h�ˤ��ҹ��j	�����*�_@��*���"���'�e,�=p0��4��8��<�/�@�uMD���G��	K�cN��Q�̺S�OV�A�X��([�Z]��_�j'b�e�d�7�f��Xi��k�HOn���p�URs���u� Nx�(�z��=}�������K��ȃ��U���.��(��Y`��!���؊����g���������A}���璼�U��VÕ�e-��r����陼x7���x��)����؞��������3���O��Fq������&ʦ�k��yD��-����ث�/(���x��dɯ�����h����������S��样���9������μ��  �  14O=��N=��M=9M=��L=��K=�K=�cJ=��I= �H=�,H=�rG=4�F=9F=�cE=n�D=�#D=�C=e�B=CgB=��A=�EA=ޱ@=�@=�?=��>=�>>=[�==w�<=�J<=d�;=��:=0S:=e�9=�9=�_8=�7=c7=�n6=��5=$$5=
~4=\�3=I,3=�~2=p�1=�1=/W0=Ɠ/=�.=��-=--=>[,=Y�+=ȵ*=�)=_)=�B(=�q'=�&=��%=/�$=*�#=E#=g"=�� =��=��=]V=T =;�=�$=.�=�=nm=�=X=�@=�p==m�	=��=O�=��=�=y��<���<��<�e�<)�<s��<s��<�/�<^��<�p�<0�<���<,r�<�0�<���<rϿ<���<���<|�<�f�<XO�<�3�<��<Y�<@��<c��<Q�<B�<׉<{��<�V�<�+z<��q<�#i<��`<�X<�O<�!G<h�><�96<>�-<M\%<��<o<��<CT<�b�;��;���;*�;���;�<�;��;H�w;9V;߿4;��;��:��:�pO:[i�9��-�(�JF���mк�=�*&���D��ic��ɀ�����I�� �������[mȻ��ջ���	yﻔ���t��qn	�����+�A@��(���"�щ'�Q	,�Zj0�_�4���8���<�ɛ@�BD���G�y�J�N���P�f�S��DV���X�� [��x]�S�_�m"b��d���f��Wi�$�k��Pn�>�p�`Vs���u��Ux���z�aG}�9�����CP�����꾄����*���a�������׊�5��f��������Kz��[䒼�Q������(�������㙼h1���r��J���9Ӟ�������</���L��~n��`���pȦ�>��D��t����٫��)��+{���̯����ym�������
���X��~�����z<������Qм��  �  �2O=/�N=g�M=~:M=ˋL=��K=R"K=RhJ=A�I=p�H=�3H=�zG=��F=F=ulE=,�D=�+D=��C=S�B=gmB=/�A=�IA=~�@=�@=ہ?="�>=�>>===��<=�G<=T�;=d�:=M:=��9=��8=�X8=��7=�7=Wi6=�5=� 5=�{4=:�3=A,3=�2=�1=-1=iZ0=ԗ/=��.=�.=4-=�b,=Y�+=D�*=��)=)=rK(=�y'=L�&=�%=��$=�$=#=W"=� =&�=�=�U=��=L�=s =ך=3=f=�=��=p8=�h=a�=�	=T�=�=��=?�=���<��<��<�i�<�.�<���<�<;�<d��<^�<�$�<���<B��<�B�<G�<-�<��<���<{��<8q�<bX�<K;�<��<f�<|��<���<�N�<��<�ω<͍�<K�<	z<�q<�i<��`<��W<��O<G<�><H,6<'�-< X%<^�<_r<��<t^<�~�;&&�;���;PH�;Nگ;�~�;[B�;bx;P�V;1Y5;�;}'�:|�:�?Q:Q��9+�'�\�&��ʑ�к@�&�w�D�yc��ڀ�ď��m��iЬ�5亻o�Ȼ�ֻ����k���x��{	���_/�n?��$��"�]'���+�xY0�4�4�^�8��<��}@��!D��G���J�r�M��P�ĎS��&V�2�X�5	[��d]���_�b��ud�i�f��Si���k��Tn���p��cs�Q�u�]kx���z�Sc}����,&��^��x���eɄ�Z����0��Pe��.���]׊����6b��Z�������q���ْ�tE��谕����-z��^ҙ����+a��[���`Þ��矼���$��)C���f��E����æ�9����B���[ܫ��.������I֯�,)���z���ʳ�����f��첷�[���MF��/����ռ��  �  �/O= �N=��M=U<M=��L=g�K=�'K=ToJ=��I=2�H=�>H=�G=��F=�#F=vzE=��D=�8D=��C=*
C=�vB=6�A=�PA=ܺ@=�!@=��?=��>=?>=Y�==��<=�B<=��;=��:=C:=p�9= �8=�L8=��7=e7=)`6=��5=5=�w4=�3=�+3=k�2=b�1=�1=1_0=�/=M�.=O.=5>-=
n,=�+=��*=��)=�))=�X(=B�'=��&=�%=G�$=�$=�#=�"=� =��=6�=gT=��=c�=�=.�=��=Z=�=f�=�*=�[=��=��	=��=P�=��=�=���<ŵ�<���<.o�<�6�<��<��<]L�<���<���<J>�<���<���<^_�<(�<i��<ջ<.��<&��<R��<�e�<F�<� �<���<���<Ј�<~J�<Q�<�É<�}�<{7�<%�y<BYq<�h<�N`<�W<�WO<w�F<�{><�6<�-<�O%<h�<iv<m�<n<��;�\�;*��;��;�6�;L�;��;7Oy;�W;�I6;h;u��:꠩:hT:�y�9D��� %�q��ϺR��f�%���D���c�m�����-������47����Ȼ�aֻc�����!�����	���I6�=@�����"��o'�{�+�*@0��y4���8�x�<�-O@�Q�C��_G�ΡJ�T�M��P�l[S���U�txX�l�Z�F]���_�)b�sfd���f�VOi�G�k�p\n���p�sys�^v�\�x�{�ݐ}�t���=��xt�������ڄ���;���k��W���q׊����\��=������yd��'ʒ��2������� ��5`���������sE���|��r����П������4��[��"���C���A���{A������T᫼O7������毼)<��J���	⳼[1��C~���ȷ����jV�������޼��  �  �+O=�N=��M=>M=J�L=j�K=�.K=�wJ=�I=tI=�LH=��G=��F=�5F=]�E=r�D=�ID=��C=�C=��B=�A=�XA=#�@=a&@=��?=	�>=�>>=ה==��<=�;<=d�;=�:=�5:=��9=a�8=�<8=P�7=g�6=�S6=G�5=5=2r4=��3=G*3=��2=��1=�1=�d0=�/=Q�.=:.=�J-=�|,=۬+=��*=B*=;)=�i(="�'=�&=��%=��$=�$=y#=�"=-� =�=ɛ=�Q=��=p�=D=Y�=��=GJ=�=�==�J=�s=��	=��=��=��=I�=w��<u��<ޛ�<u�<M@�<b��<b��<b�<��<M��<_�<��<$��<ԃ�<iK�<��<e�<&ѷ<h��<ה�<�u�<�R�<�)�<B��<�Ú<B��<yC�<k��<���<�g�<3�<}�y<xq<�h<?`<\�W<�O<��F<�R><��5<0�-<eB%<��<Cy<i<�<��;��;zQ�;���;���;�i�;�B�;�~z;��X;�}7;ڏ;P�:��:>�W:�|�9[l�m#��=����κ��A�%���D���c�7&��2�������{������8rɻ�ֻ��ud���S���	��� B�D���O�"��^'���+�"0�NT4��d8�.P<�5@�|�C�NG�'ZJ��mM�WP�MS���U��CX�m�Z�� ]���_��a�Vd���f�8Li���k�9in�$ q�L�s�y.v�пx�IJ{�>�}��#��]��,����Ã��%��nI���u��Τ���؊����1W��Y���W����T��Ŷ����������▼3?������ߚ�"���Z�����������٠�����#��fM���}��>���x��� A��c���髼�C�����������U��㬲�� ���P��8����巼{*��hl��7���n뼼�  �  &O=ÆN=��M=�>M= �L=5�K=v5K=��J= �I=�I=�\H=+�G=��F=�IF=��E=n�D=k\D=@�C='C=��B=��A=.aA=��@=�*@=�?=v�>=�<>=�==��<=�2<=�;=��:=�%:=z9=��8=*8= �7=z�6=�D6=��5= 	5=�j4=��3=�'3={�2=�1="1=)j0=��/=��.="#.=Y-=Č,=�+=�*=T *=�O)=)}(=$�'=.�&=��%=�
%=�$=Z#=D"=�� =��='�=N=��=w�=�=�w=��==7=j�=:�=�="6=�`=��	=��=S�=��=��=`��<ư�<~��<�y�<�I�<4�< ��<�y�<a(�<���<V��<�6�<���<h��<�s�<'A�<a�<��<�˳<���<$��<�^�<2�<N��<WÚ<Z��<N9�<��<q��<M�<f��<�_y</�p<?h<3�_<FW<T�N<yF<!><<�5<$�-<�/%<��<Ox<#<�<P�;H��;R��;�k�;�.�;?��;g�;��{;1Z;[�8;$�;St�:gɭ:.Z[:�9��
��� �kj���Qκ�����%��E��d�?a��Ђ��|b����+����ɻ�i׻<b����;���C�o�	��,��S�FL���k�"�gO'���+��0�k,4��38��<���?��cC�w�F�pJ��M��P�b�R��yU�
X�K�Z���\��e_�.�a�KGd���f�#Mi�)�k��{n��q�B�s��_v�n�x�7�{��~��I�����׵��;䃼\���5���[��Ђ�������܊�d���R�� ���쏼XD��ۡ��6���b���������Bl��%�������4��;g����������硼)��I?���s��&���J���C��}�������S��ܴ�����ct��dϲ��%���v��+¶�g���I��1�����������  �  �O=�N=%�M=�>M=�L=
�K=�;K=.�J="�I=� I=�lH=l�G=�
G=�^F=�E=GE=pD=�C=�6C=��B=AB=iA=�@=.@=t�?=��>=�9>=��==��<=�(<=�u;=��:=�:=pf9=-�8=S8=r7=��6=;46=d�5=Z�4=�a4=P�3=�#3=�~2=��1={$1=�n0=[�/=$�.=�..=cg-=�,=��+=>+=E5*={d)=S�(=ú'=��&=��%= %=�#$=�%#=
"=<� =��=%�=�H=��=�w=#�=�g=�=A"=�n=�=��=�=L=Zr	=��=��=(�=��=[��<q��<Ț�<�|�<Q�<��<-��<���<�E�<.��<���<�`�<��<���<q��<h�<O8�<�<��<���<d��<ui�<:8�<! �<i��<�y�<!,�<�ٍ<Ʉ�<�.�<�ـ<y<�up< �g< f_<�V<E�N<6F</�=<J�5<�\-<�%<��<�r<�<��<�;�;(�;��;���;�;)��;*��;�D};<�[;�L:;d>;f��:b�:�?_:j��9� ���������ͺ {���%�+PE��wd�b�������P՟�<y��#�����ʻ�ػ[��~u��p��|y�h�	�gN��j�Z�� ���"��C'�ɤ+���/� 4�08���;���?��C�CyF�#�I�{�L�u�O���R�5U���W�zVZ�u�\��H_�ʿa�u<d��f�/Si���k�;�n�m?q���s���v�&<y�L�{�ze~��r������H݂�l��(.���P��9q��	���!���㊼p���P��ה��[ᏼ5�������蓼*D��h������B������rϛ����MB��t��Ţ��vС������2���k�����_����G��y������f��Zͮ�r3����������6N��O����궼�.���l��h���ۻ�����  �  �O=|N=n�M=�<M=T�L=��K=t@K=��J= �I=2-I=�{H=��G=8G=sF=��E=�%E=�D=!�C=AEC=¨B=�B=�oA=x�@=80@=`�?=��>=�5>=9�==��<=<=�g;=s�:=I:=@R9=�8= 8=S]7=l�6=�"6==�5=��4=�W4=ļ3=|3=�{2=v�1=�%1=�q0=�/=S�.=�9.=�t-=d�,=��+=�+=�I*=�x)=�(=��'=��&=&= %=R+$=�*#=�"=r� =��=ے=B=��=.l=��=�V=x�=�=�W=�=��=�=�6=�^	=��=��=��=��=��<���<N��<�|�<4V�<A$�<8��<���<fa�<'�<x��<<��<ZD�<�<��<���<�Y�<n)�<���<�ϯ<'��<tq�<�;�<��<�<=o�<��<ō<8j�<��<㴀<	�x<Hp<
�g<�_<��V<a?N<��E<ҫ=<lo5<e5-<�$<��<�g<�<��<@`�;�b�;�W�;wF�;�6�;~/�;87�;��~;�];Ȳ;;�;,k�:�1�:�b:��9J��0&��#����ͺ�{��&�h�E��d����� F��/O�����WX���=˻��ػj��
�)���]��;/
�t�Ն��l��*��"��='�ߕ+���/���3���7���;��L?�,�B�w)F�`I�<sL�_eO��9R���T�:�W��)Z�'�\��0_�R�a��6d�!�f�V^i��l�H�n�Ffq��t�*�v� �y��#|�˷~�~���ց�����-���O��m������W����ŉ��늼#��)Q�����'ُ��'��W{��(ѓ�K'���{��J͗�w��c��g����䜼���U��ƈ��⻡�Q�:(���e��Ϊ��L���~N��謪����{���箼�R����������w���ʵ�����V��ߐ��Lź�����m%���  �  �O=NuN=��M=7:M=��L=��K=�CK=x�J=��I=:8I=[�H=��G=�/G=��F=��E=�7E=0�D=e�C=<RC=6�B=�B=FuA=e�@=1@=-�?=g�>=�0>=~==��<=u<=�Y;=h�:=V�9=�>9=Ԓ8=��7=xI7=ū6=�6=qz5=!�4=hM4=��3=l3=�w2=V�1=u%1=�s0=-�/=�/=�B.=��-=��,=��+=�)+=-\*=b�)=��(=��'=��&=�&=t)%=�1$=I.#=�"=w� =��=��=�:=�=O`=t�=F=��=��=�A=H�=��=��=
"=7L	=1q=y�=��=;�=5��<��<���<�z�<�X�< ,�<p��<Z��<�y�<�6�<_��<��<�j�<z)�<���<N��<w�<:B�<��<(ޯ<���<�v�<m<�<���<Y��<3c�<"�<���<�O�<_�<��<3ox<d�o<!7g<_�^<�KV<[�M<��E<�p=<==5<�-<�$<q�<�X<�<��<xy�;���;"��;���;C��;��;�͐;�;�Y^;��<;��;��:��:�f:ş�9�H޸\���č�Iͺʏ��O&�!�E�ohe��I�������Ơ�"����뽻��˻xHٻY4滫��ny����T_
���$����9���"�d<'���+�i�/���3�J�7�t;��?�ŋB�J�E��I��'L��O�	�Q�/�T�efW��Z���\��_�p�a�16d���f�jmi��l���n���q�7Ot�Hw��y��m|���*ƀ������,��9R��2p��7���j���p���iԉ������ ��T��ݏ���ӏ����,l��ϼ������]��H�������Y=��3�����������j9��$r��r����㢼� ���b��᫦�W���eW��蹪�F#���������kq��Rݱ��B�������=���|�� ���g亼����;���  �  [O=�nN=��M=�6M=�L=�K=FK=��J=�I=AI=v�H=��G=4>G="�F=x�E=9GE=i�D=�C=�\C=��B=�B=yA=�@=�0@=1�?=��>=J+>=w==�<=�<=`M;=�:=��9=�-9=�8=��7=	87=T�6=�6=m5=��4=�C4=�3=e3=;s2=��1=^$1=�t0=��/=�/=+J.=1�-==�,=U,=I8+=�k*=��)=S�(=a�'=E	'=!&=|0%=36$=�0#="=�� =$�=V�=�3=#�=bU={�=7=�=��=X.=do= �=�=�=�;	=gb=��=۞=J�=؀�<F��<Ĉ�<Lw�<�Y�<#1�<[ �<S��<���<O�<u�<���<��<�I�<c	�<*��<w��<HV�<�< �<O��<�x�<;�<���<<1W�<=��<���<�7�<1ӄ<Sq�<�)x<ʀo<��f<�l^<�V<j�M<�nE<�:=<�5<��,<��$<�<�H<��<��<L��;��;w��;���;��;�%�;K�;{�;lo_;]>;�;�k�:ǭ�:�h:6��9S�Ҹ����ۈͺU���&��MF��e�E�������1����n��/a̻G�ٻ�滗�D������
����Y��G���H� �"�J?'��+��/���3�)�7��L;���>� UB�#�E�`�H�d�K��N�޿Q��T��>W�~�Y��~\�;_��a��9d���f�~i�J1l���n��q�{|t�Bw�`�y��|�L��逼3"��8O��0r��)���¢��,���aʈ��≼���t(��QX��Ӑ���Џ�����`����������D��#���uט����b��G���o䝼�"���_��ݜ���ڢ���b��Ů��l���`���ƪ��3���������񌰼
���7d��3ô�n��d`��s���ӹ�J ���(��P���  �  k�N=+iN=r�M=�3M=,�L=��K=3GK=��J=��I=yGI=��H=p�G=)IG=͠F=Y�E=�RE=�D=oD=�dC=��B=�B=o{A=��@=0@="�?=g�>=�&>=;q==��<=B�;=]C;=��:=��9=m 9=4s8=��7=a*7=d�6=��5=lb5=j�4=�;4=f�3=:3=;o2=��1=#1=�t0=��/=C
/=KO.=�-=��,=f,=kC+=Qw*=��)=s�(=o�'=�'=�'&=p5%=N9$=�1#=�"=�� =��=��=�-=��=�L=:�=M+=��=j�===�_=��=t�=�=�.	=�V=~y=�=�=�t�<��<=��<�s�<"Y�<#4�<9�<��<K��<>a�<�#�<#��<Q��<�a�<x �<��<f��<�d�<	*�<P�<;��<�y�<�8�<��<��<�L�<��<Z��<D$�<μ�<6X�<�w<6Go<��f<2^<��U<�{M<�>E<�=<	�4<��,<`�$<�r<O:<9�<;�<���;���;)��;;$�;�M�;�y�;��;���;g@`;��>;5�;���:�Զ:j:�p�9�A˸
k�����U�ͺF��/�&�S�F��Ff�5Ԃ�RQ��*����c���Ծ�0�̻s>ڻ�$绾|�GI���H���
�y���������W���"��C'���+�m�/�g�3��|7�G0;�W�>��+B��wE�إH�ȸK��N�j�Q� eT��!W���Y�[p\��
_��a�,>d���f�^�i�REl�!o���q�v�t��kw�l.z�F�|�������>��-j��u���&�������Ǉ�&و�����/���\�������Ϗ�R���X������锼a2���y��}������J��$����Н����R��I���բ�l��{b�����X	��ai���Ѫ�'A�������,��â��U��{~���޴�o3���{��츸��빼g��Q<���`���  �  ��N=geN=��M=�1M=̑L=3�K=�GK=�J=f�I=[KI=��H=b�G=�OG=��F=� F=�YE=��D=)D=biC=*�B=5!B=�|A=�@=\/@=��?=�>=�#>=Im==�<=��;=�<;=��:=�9=�9=]j8=��7=�!7=+�6=I�5=�[5=h�4=�64=�3=�	3=�l2=
�1=�!1=�t0=c�/=4/=[R.=M�-=�,=�,=AJ+=�~*=��)=F�(=��'='=�+&=g8%=;$=}2#=$"=N� =��=x�=�)=��=�F=��=�#=^~=^�=�=V=�=��=��
=k&	=TO=�r=k�=&�=m�<�|�<�}�<q�<eX�<�5�<X�<���<H��<_l�<�0�<p��<X��<�p�<�.�<���<A��<ym�<s0�<u��<���<�y�<�6�<�<���<�E�<��<{��<��<k��<'H�<Y�w<�"o<J�f<�^<�U<OZM<� E<}�<<C�4<�,<��$<�e<�0<	�<ס<(��;h��;��;�E�;�x�;C��;��;��;��`;T?;0 ;���:���:�k:��9�Ƹ�,�����ͺ!����&��F�|�f�����Ӂ��Y�����������ͻ��ڻQh绻��7����b���
�V��k�����a�}�"�[G'���+���/��3��o7��;�ܩ>��B��[E�z�H�Z�K��N��|Q�lOT�2W���Y��g\�	_�_�a�-Bd���f���i��Rl��o���q��t�w�oLz��}�������O��B{������β��)Ć�Ӈ��∼����x��T4��`��%���\Ϗ�����S���������#'���l��a���R���$<�������ĝ�����J�������Ѣ�Z��Rc������t��
o���ت�J��x���%9�������#��)���:�;E�������ɸ�6����$���H��uk���  �  M�N=dN=s�M=�0M=C�L=�K=�GK=��J=2�I=�LI=H�H=j�G=6RG=s�F=<F=O\E=��D=D=kC=O�B=�!B=7}A=;�@=/@=��?=9�>=i">=�k==K�<=��;=�:;=�:=;�9=�9=Sg8=�7=�7=K�6=��5=CY5=T�4=54=��3=o3=�k2=Q�1=}!1=}t0=��/=�/=IS.=��-=��,=�,=�L+=��*=7�)=��(=��'=�'=g-&=M9%=�;$=�2#="=�� =��=X='(=-�=�D=A�=2!=�{=C�=o=�R=��=��=��
=�#	=�L=�p=��=��={j�<�z�<f|�<ep�<~X�<�6�<��<���<}��<Dp�<B5�<c��<���<�u�<i3�<��<֯�<7p�<:2�<���<p��<Jy�<�5�<n�<|��<�B�<��<�|�<�<H��<mB�<�w<�o<�~f<9 ^<��U<�NM<HE<o�<<��4<%�,<4�$<�a<�-<%�<��<���;���;X�;hQ�;(��;J��;$��;]5�;j�`;	?;d(;���:�÷:�l:���9��Ÿ �ꃍ�"�ͺ��� '���F���f�g�������ҡ����(.��)ͻӛڻ?�绎��.���,l��
���"��߾�[e�3�"��H'���+�M�/���3�l7�;���>��	B�KRE�Y~H�/�K�L�N�$tQ�HT�<
W��Y�ye\��_�M�a��Cd���f�c�i��Wl��o���q�N�t��w��Vz�P}�������U��.���#���귅��Ȇ��և�戼�������6��Ha������1Ϗ����R��◓��ݔ�Q#��yh������C�07���{��g���k��H��狡��Т�����c������ �� q���۪�$M��ĭ�n=������<)������D���JK�������ϸ�� ��u)��0M��-o���  �  ��N=geN=��M=�1M=̑L=3�K=�GK=�J=f�I=[KI=��H=b�G=�OG=��F=� F=�YE=��D=)D=biC=*�B=5!B=�|A=�@=\/@=��?=�>=�#>=Im==�<=��;=�<;=��:=�9=�9=]j8=��7=�!7=+�6=I�5=�[5=h�4=�64=�3=�	3=�l2=
�1=�!1=�t0=c�/=4/=[R.=M�-=�,=�,=AJ+=�~*=��)=F�(=��'='=�+&=h8%=;$=2#=&"=R� =��=�=�)=��=�F=��=�#={~=��=�=EV=�=9�=�
=�&	=�O=Cs=ǐ=��=�m�<�}�<�~�<�q�<Y�<n6�<��<��<���<�l�<�0�<���<_��<�p�<v.�<���<㫼<m�<�/�<��<V��<�x�<6�<a�<��<�D�<P�<��< �<��<�G�<��w<P"o<H�f<%^<M�U<�ZM<e!E<r�<<]�4<��,<�$<Zg<#2<s�<8�<ɗ�;���;��;�G�;xz�;q��;��; �;��`;S?;L�;5��:���:�k:���9ƟǸbD�{�����ͺ����&���F�f�� ����������*�������ͻb�ڻ�i���b���[c�U�
����������a���"�|G'��+�ɣ/�#�3�p7��;��>��B��[E�~�H�]�K��N��|Q�mOT�3W���Y��g\�
_�_�a�-Bd���f���i��Rl��o���q��t�w�oLz��}�������O��B{������β��)Ć�Ӈ��∼����x��T4��`��%���\Ϗ�����S���������#'���l��a���R���$<�������ĝ�����J�������Ѣ�Z��Rc������t��
o���ت�J��x���%9�������#��)���:�;E�������ɸ�6����$���H��uk���  �  k�N=+iN=r�M=�3M=,�L=��K=3GK=��J=��I=yGI=��H=p�G=)IG=͠F=Y�E=�RE=�D=oD=�dC=��B=�B=o{A=��@=0@="�?=g�>=�&>=;q==��<=B�;=]C;=��:=��9=m 9=4s8=��7=a*7=d�6=��5=lb5=j�4=�;4=f�3=:3=;o2=��1=#1=�t0=��/=C
/=KO.=�-=��,=f,=kC+=Pw*=��)=s�(=o�'=�'=�'&=r5%=Q9$=�1#=�"=�� =��=��=�-=��=�L=`�={+=�=��=�=>`=�=��=N=7/	=YW=&z=Ŗ=��=Qv�<[��<���<"u�<wZ�<_5�<W�<���<��<�a�<$�<e��<`��<�a�<! �<���<���<�c�<)�<.�<��<yx�<�7�<o�<š�<�K�<��<K��<W#�<	��<�W�<N�w<�Fo<��f<~2^<W�U<�|M<�@E<{=<*�4<��,<�$<�u<=<��<�<Ŗ�;��;f��;�'�;�P�;�{�;���;��;@`;��>;��;7��:cǶ:8kj:�%�9I�̸:������$�ͺ�����&�ΨF��Rf�ڂ��V��H���:h��Aپ�
�̻�Aڻ�'�[�K��yI���
�'�������X���"��C'�ֆ+���/���3��|7�\0;�h�>��+B��wE��H�θK��N�n�Q�#eT��!W���Y�\p\��
_��a�->d���f�_�i�REl�!o���q�w�t��kw�l.z�F�|�������>��-j��u���&�������Ǉ�&و�����/���\�������Ϗ�R���X������锼a2���y��}������J��$����Н����R��I���բ�l��{b�����X	��ai���Ѫ�'A�������,��â��U��{~���޴�o3���{��츸��빼g��Q<���`���  �  [O=�nN=��M=�6M=�L=�K=FK=��J=�I=AI=v�H=��G=4>G="�F=x�E=9GE=i�D=�C=�\C=��B=�B=yA=�@=�0@=1�?=��>=J+>=w==�<=�<=`M;=�:=��9=�-9=�8=��7=	87=T�6=�6=m5=��4=�C4=�3=e3=;s2=��1=^$1=�t0=��/=�/=+J.=1�-==�,=U,=H8+=�k*=��)=S�(=a�'=F	'=!&=0%=66$=�0#="=�� =3�=j�=�3=E�=�U=��=]7=3�=�=�.=�o=��='�=�=z<	=Ec=��=՟=L�=��<Y��<ϊ�<Gy�<b[�<�2�<��<���<��<�O�<�<E��<"��<oI�<��<j��<v��<U�<��<e�<���<(w�<+9�<���<��<jU�<���<��<A6�<҄<{p�<�(x<1�o<��f<m^<V<�M<qE<�==<�5< �,<J�$<�<�L<�<��<|��;���;u��;��;,�;�(�;=M�;|�;�n_;�>;��;�\�:���:�h:22�9Y�Ը�6������ͺ4����&�h_F�5�e�{�������8���
��$t���f̻�ٻ.��I�r���� ���
����%����yI�p�"��?'�Q�+�$�/��3�N�7��L;���>�UB�2�E�k�H�m�K���N��Q��T��>W���Y��~\�<_��a��9d���f�~i�K1l���n��q�{|t�Bw�`�y��|�L��逼3"��8O��0r��)���¢��,���aʈ��≼���t(��QX��Ӑ���Џ�����`����������D��#���uט����b��G���o䝼�"���_��ݜ���ڢ���b��Ů��l���`���ƪ��3���������񌰼
���7d��3ô�n��d`��s���ӹ�J ���(��P���  �  �O=NuN=��M=7:M=��L=��K=�CK=x�J=��I=:8I=[�H=��G=�/G=��F=��E=�7E=0�D=e�C=<RC=6�B=�B=FuA=e�@=1@=-�?=g�>=�0>=~==��<=u<=�Y;=h�:=V�9=�>9=Ԓ8=��7=xI7=ū6=�6=qz5=!�4=hM4=��3=l3=�w2=V�1=u%1=�s0=-�/=�/=�B.=��-=��,=��+=�)+=-\*=b�)=��(=��'=��&=�&=v)%=�1$=P.#=�"=�� =��=ʍ=�:=D�=�`=��=\F=��=_�=6B=�=��=��=�"=3M	=Br=��=�=x�=���<���<x��<J}�<[�<$.�<`��<��<1{�<�7�<)��<���<�j�<:)�<5��<b��<�u�<�@�<��<1ܯ<���<Qt�<:�<H��<��<a�<
�<���<(N�<
�<��<�mx<��o<7g<�^<3MV<`�M<F�E<�s=<�@5<�-<y�$<�<�]<�<Y�<F��;���;y��;T��;y��;��;DА;r�;TY^;;�<;8�;��:D�:7�e:��9Ǌฦ*�#B�ͺ����e&��	F�m}e��S�����hϠ�J���I󽻁�˻dNٻ�9�2��S}������`
�I��������9�A�"��<'��+���/���3�x�7�Ct;��?�ۋB�\�E��I��'L��O��Q�5�T�ifW��Z���\��_�q�a�36d���f�kmi��l���n���q�7Ot�Iw��y��m|���*ƀ������,��9R��2p��7���j���p���iԉ������ ��T��ݏ���ӏ����,l��ϼ������]��H�������Y=��3�����������j9��$r��r����㢼� ���b��᫦�W���eW��蹪�F#���������kq��Rݱ��B�������=���|�� ���g亼����;���  �  �O=|N=n�M=�<M=T�L=��K=t@K=��J= �I=2-I=�{H=��G=8G=sF=��E=�%E=�D=!�C=AEC=¨B=�B=�oA=x�@=80@=`�?=��>=�5>=9�==��<=<=�g;=s�:=I:=@R9=�8= 8=S]7=l�6=�"6==�5=��4=�W4=ļ3={3=�{2=u�1=�%1=�q0=�/=R�.=�9.=�t-=c�,=��+=�+=�I*=�x)=�(=��'=��&=&=� %=W+$=�*#=�"=�� =��=��=@B=��=hl=�=�V=�=-=[X=��=��=�	=�7=
`	=ւ=�=ܶ=)�=Ԡ�<b��<��<��<�X�<�&�<a��<e��<�b�<e�<Z��<���<wD�<��<h��<���<&X�<�'�<��<^ͯ<ǟ�<�n�<9�<q��<g��<�l�<q�< Í<nh�<0�<���<v�x<xp<�g<�_<0�V<�AN<��E<c�=<�s5<�9-<��$<ٺ<�l<<ϩ<j�;�k�;�_�;�M�;^<�;�3�;:�;5�~;�];�;;݋;�V�:~�:.�b:"��9a�}��Q��{�ͺ+��2&���E��e�"���P��Y������`��HE˻��ػ8������7���0
�Su����m��+���"�>'�C�+���/���3���7���;��L?�E�B��)F�`I�HsL�ieO��9R���T�?�W��)Z�)�\��0_�T�a��6d�"�f�W^i��l�I�n�Ffq��t�*�v� �y��#|�̷~�~���ց�����-���O��m������W����ŉ��늼#��)Q�����'ُ��'��W{��(ѓ�K'���{��J͗�w��c��g����䜼���U��ƈ��⻡�Q�:(���e��Ϊ��L���~N��謪����{���箼�R����������w���ʵ�����V��ߐ��Lź�����m%���  �  �O=�N=%�M=�>M=�L=
�K=�;K=.�J="�I=� I=�lH=l�G=�
G=�^F=�E=GE=pD=�C=�6C=��B=AB=iA=�@=.@=t�?=��>=�9>=��==��<=�(<=�u;=��:=�:=pf9=-�8=S8=r7=��6=;46=d�5=Z�4=�a4=P�3=�#3=�~2=��1={$1=�n0=[�/=$�.=�..=bg-=�,=��+=>+=E5*={d)=S�(=ú'=��&=��%=%=�#$=�%#="=K� =�=@�=�H=��=x=n�=h=}�=�"=~o=��=[�=� =!M=|s	=ϓ=I�=��=T�=F��<_��<���<S�<�S�<F�<i��<���<WG�<w��<��<a�<�<���<�<�f�<�6�<O�<��<k��<<�f�<�5�<t��<ɽ�<w�<�)�<�׍<<3-�<�؀<fy<up<��g<�f_<��V<��N<9F<��=<��5<�a-<�%<��<x<<�<(F�;�1�;f�;���;���;���;+��;WG};��[;�H:;7;a��:W�:��^:^��9�i�h3�l⎺�κE��&�iE��d������됻�ߟ������Ǽ�8�ʻ�ػ^廸z�{u��g{�
��O�l��Z��!�y�"�ZD'�0�+�(�/�B4�e8��;���?��C�WyF�3�I���L��O��R�5U���W�~VZ�w�\��H_�̿a�v<d��f�/Si���k�<�n�n?q���s���v�&<y�L�{�ze~��r������H݂�l��(.���P��9q��	���!���㊼p���P��ה��[ᏼ5�������蓼*D��h������B������rϛ����MB��t��Ţ��vС������2���k�����_����G��y������f��Zͮ�r3����������6N��O����궼�.���l��h���ۻ�����  �  &O=ÆN=��M=�>M= �L=5�K=v5K=��J= �I=�I=�\H=+�G=��F=�IF=��E=n�D=k\D=@�C='C=��B=��A=.aA=��@=�*@=�?=v�>=�<>=�==��<=�2<=�;=��:=�%:=z9=��8=*8=�7=z�6=�D6=��5= 	5=�j4=��3=�'3=z�2=�1="1=(j0=��/=��.=!#.=Y-=Ì,=�+=�*=S *=�O)=)}(=$�'=/�&=��%=�
%=�$=a#=O"=�� =��=B�=3N=��=��=�=Qx=B�=�7=�=��=�=7=�a=�	=�=��= �=H�=2��<���<I��<�|�<&L�<��<I��<�{�<�)�<���<7��<E7�<���<!��<�r�< @�<�<*�<�ɳ<u��<Ã�<p\�<o/�<���<���<�~�<
7�<��<���<�K�<@��<�]y<_�p<�>h<�_<�GW<��N<|F<�$><X�5<��-<l4%<��<�}<j<9�<#�;e��;���;�r�;�4�;��;N�;[�{;u0Z;~�8;�;`�:E��:9[:$}�9���4!�����|�κ��n�%��0E��,d�tl��g���\l������R3��Iʻlp׻
h��������D� �	�K.��T�,M�r��"��O'���+�0��,4��38��<���?� dC���F��J��M��P�i�R��yU�
X�O�Z���\��e_�/�a�MGd���f�$Mi�*�k��{n��q�B�s��_v�n�x�7�{��~��I�����׵��;䃼\���5���[��Ђ�������܊�d���R�� ���쏼XD��ۡ��6���b���������Bl��%�������4��;g����������硼)��I?���s��&���J���C��}�������S��ܴ�����ct��dϲ��%���v��+¶�g���I��1�����������  �  �+O=�N=��M=>M=J�L=j�K=�.K=�wJ=�I=tI=�LH=��G=��F=�5F=]�E=r�D=�ID=��C=�C=��B=�A=�XA=#�@=a&@=��?=	�>=�>>=ה==��<=�;<=d�;=�:=�5:=��9=a�8=�<8=P�7=g�6=�S6=G�5=5=2r4=��3=F*3=��2=��1=�1=�d0=�/=P�.=9.=�J-=�|,=ڬ+=��*=A*=;)=�i(="�'=	�&=��%=��$=�$=�#=�"=:� =+�=�=R=�=��=�=��=�=�J=l�=�=�=TK=�t=��	=�=�=��=��=���<���<_��<tw�<�B�<��<R��<�c�<)�<k��<�_�<"�<=��<���<�J�<��<*�<�Ϸ<���<ߒ�<ys�<WP�<~'�<���<j��<��<qA�<���<!��<�f�<,�<�y<�q<�h<�`<��W<� O<��F<*V><]�5<G�-<�F%<G�<�}<$<7�<���;5��;�X�;,�;ర;�m�;gE�;Q�z;T�X;pz7;��;��:���:�HW:���9����Y#�g���Ϻ���* &�}E���c�C0��~;�����ڃ�� ����xɻ�ֻM���h�v�����%�	���C��D�]���"�H_'�A�+�V"0��T4��d8�RP<�R@���C�_G�5ZJ��mM�WP�TS���U��CX�p�Z�� ]���_��a�Vd���f�9Li���k�9in�$ q�L�s�z.v�ѿx�IJ{�>�}��#��]��,����Ã��%��nI���u��Τ���؊����1W��Y���W����T��Ŷ����������▼3?������ߚ�"���Z�����������٠�����#��fM���}��>���x��� A��c���髼�C�����������U��㬲�� ���P��8����巼{*��hl��7���n뼼�  �  �/O= �N=��M=U<M=��L=g�K=�'K=ToJ=��I=2�H=�>H=�G=��F=�#F=vzE=��D=�8D=��C=*
C=�vB=6�A=�PA=ܺ@=�!@=��?=��>=?>=Y�==��<=�B<=��;=��:=C:=p�9= �8=�L8=��7=e7=)`6=��5=5=�w4=�3=�+3=k�2=a�1=�1=1_0=�/=M�.=O.=5>-=
n,=�+=��*=��)=�))=�X(=B�'=��&=�%=I�$=�$=�#=�"=� =��=J�=�T=��=��=�=o�=�=wZ=��=��=�+=D\=>�=j�	=��==�=��=�=���<ط�<���<)q�<�8�<���<���<�M�<	��<���<�>�<���<Р�<*_�<�'�<���<Ի<�<���<��<d�<JD�<��<��<��<	��<�H�<��<g<�|�<�6�<��y<�Xq<�h<)O`<-�W<sYO<��F<(~><�6<h�-<BS%<.�<Fz<J�<�q<K��;gc�;+�;K��;�:�;��;?��;&Qy;��W;!G6;�b;���:ō�:J�S:��9� ��`%�H3��*�Ϻ/��J&�l�D�ިc����^���f���4 ��B=��`ɻ�fֻCg�u��%�����&�	����7��@�/ �8�"�*p'���+�e@0��y4�Ǒ8���<�DO@�d�C��_G�ڡJ�]�M���P�q[S���U�wxX�o�Z�F]���_�+b�tfd���f�WOi�G�k�q\n���p�sys�_v�\�x�{�ݐ}�t���=��xt�������ڄ���;���k��W���q׊����\��=������yd��'ʒ��2������� ��5`���������sE���|��r����П������4��[��"���C���A���{A������T᫼O7������毼)<��J���	⳼[1��C~���ȷ����jV�������޼��  �  �2O=/�N=g�M=~:M=ˋL=��K=R"K=RhJ=A�I=p�H=�3H=�zG=��F=F=ulE=,�D=�+D=��C=S�B=gmB=/�A=�IA=~�@=�@=ہ?="�>=�>>===��<=�G<=T�;=d�:=M:=��9=��8=�X8=��7=�7=Wi6=�5=� 5=�{4=:�3=@,3=�2=�1=,1=hZ0=ӗ/=��.=�.=4-=�b,=X�+=D�*=��)=)=rK(=�y'=L�&=�%=��$=�$=#=\"=� =0�=�=�U=��=j�=� =�=k=Kf=a�=H�=�8=
i=�=��	=��=��=l�=��=a��<Z��<X��<�j�<�/�<��<��<<�<6��<��<�$�<A��<Q��<�B�<��<�߿<T��<͟�<v��<p�<'W�<�9�<T�<�<,��<c��<�M�<v�<�Ή<��<xJ�<9z<��q<�i<�`<N X<ǃO<�G<��><h.6<��-<�Z%<	�<u<B�< a<��;�*�;ο�;�K�;Rݯ;뀞;�C�;ccx; �V;1W5;|;��:��:+Q::U�9I�(��'��⑺�$к�&��!&���D�,�c������ɏ��r��լ�}躻H�Ȼdֻ�㻁�ﻬ���n���{	�����/��?��$�m�"��'���+��Y0�V�4�x�8�(�<�~@��!D��G���J�x�M��P�ȎS��&V�5�X�7	[��d]���_�b��ud�j�f��Si���k��Tn���p��cs�Q�u�]kx���z�Sc}����,&��^��x���eɄ�Z����0��Pe��.���]׊����6b��Z�������q���ْ�tE��谕����-z��^ҙ����+a��[���`Þ��矼���$��)C���f��E����æ�9����B���[ܫ��.������I֯�,)���z���ʳ�����f��첷�[���MF��/����ռ��  �  14O=��N=��M=9M=��L=��K=�K=�cJ=��I= �H=�,H=�rG=4�F=9F=�cE=n�D=�#D=�C=e�B=CgB=��A=�EA=ޱ@=�@=�?=��>=�>>=[�==w�<=�J<=d�;=��:=0S:=e�9=�9=�_8=�7=c7=�n6=��5=$$5=
~4=\�3=I,3=�~2=p�1=�1=/W0=œ/=�.=��-=--=>[,=Y�+=ȵ*=�)=_)=�B(=�q'=�&=��%=0�$=+�#=G#=j"=�� =��=��=fV=` =K�=�$=F�=�=�m=F�=�=A=�p=�=��	=��=��=!�=s�=;��<V��<���<�f�<�)�<��<��<j0�<���<�p�<l�<���<4r�<�0�<u��<,Ͽ<B��<L��<�{�<�e�<�N�<O3�<K�<��<���<���<hP�<��<�։<��<�V�<;+z<Ƨq<�#i<��`<MX<��O<n"G<\�><;6<w�-<�]%<$�<}p<D�<�U<fe�;
�;+��;�;=��;'>�;���;��w;V;־4;��;}�:��:�_O:{B�9;�-�'(��R���zк�D��0&�o�D��oc��̀�����uL����������XoȻ��ջq��cz﻿������n	�G��&,�~@� )���"��'�l	,�oj0�p�4���8���<�қ@�BD���G�}�J�N���P�h�S��DV���X�� [��x]�S�_�n"b��d���f��Wi�$�k��Pn�>�p�aVs���u��Ux���z�aG}�9�����CP�����꾄����*���a�������׊�5��f��������Kz��[䒼�Q������(�������㙼h1���r��J���9Ӟ�������</���L��~n��`���pȦ�>��D��t����٫��)��+{���̯����ym�������
���X��~�����z<������Qм��  �  �EO=@�N=N�M=�LM=�L=��K=B*K=�iJ=@�I=f�H=�H=�]G=�F=��E=�HE=c�D=�D=ӀC=a�B="oB=��A=�`A=6�@=�D@=2�?= ?=�t>=��==P-==�<=.�;=?;=�:=9�9=�V9==�8=[8={n7=��6=P)6=L�5=G�4=fB4=O�3=a�2==F2=��1=��0=�0=(I/=hz.=g�-=#�,=�,=`2+=re*=�)=��(=�(=EK'=/�&=M�%=i�$=:�#=.�"=}�!=�� =��=�d=-=l�=S4=��=�=9v=�==�6=Z]=wy=��
=c�=��=�=��=p� =���<���<$��<#,�<���<�X�<���<�b�<��<�o�<'�<n��<�X�<)�<!�<�ϻ<㹷<�<I��<ȉ�<Sr�< S�<�*�<���<C<5��<�D�<w�<��<�z�<�iz<;�q<LGi<k�`<�X<g�O<��F<�e><;�5<Bd-<��$<g<��<�@<@�<���;��;t�;�5�;=X�;���;�;&o;"�L;�B+;�;
;���:�:�(:�-9�P��6{N������N�"}�^�0�?�O��n�|����ѕ�����8,���g��0Qϻ[�ܻ�����������R�.��������!���&��P+��/��-4�=s8���<���@��pD��H��K���N�ɨQ��eT���V��MY�[��]���_�>�a��d��Ff� �h���j�aDm�6�o� r���t�	�v�ey���{��.~�_I��|������ーp���H��}z��[���G�������X������.����Y���Ƒ��;��4���|0��������p��"���X����(��KF��PX��Nc���k��Pw����������ͦ�y ��(>������ϫ�����l������W��S������c괼7��ǃ��Rи�����e��鮼��  �  qEO=\�N=��M=�MM=T�L=��K=;,K=lJ=ݨI=k�H=>!H=�aG=�F=�E=�LE=��D=�D=��C=��B=rB=>�A=�bA=$�@=wF@=j�?=?=+u>=��==�,==�<=��;=�<;=!�:=�9=qS9=ٰ8="8=�k7=6�6=j'6=�5=��4=3B4=��3=�2=OG2=��1=z�0=�0=pK/=&}.=��-=��,=s,=n6+=�i*=M�)=��(=�(=�N'=F�&=��%=��$=�#=��"=��!=�� =)�=�d=�=q�=�2=^�=�=�r=]�= =�2=�Y=v=��
=
�=:�=�=�=1� =(��<���<��<�.�<N��<]�<���<�h�<��<�w�<q�<��<�a�<�$�<O��<#׻<���<��<���<���<�v�<pV�<f-�<���<5Ö< ��<�C�<���<2��<xu�<L]z<��q<�8i<&�`< X<]vO<��F<0^><��5<�`-<=�$<wg<��<VD<u�<%��;���;!*�;fM�;�s�;¯�;��;�fo;�-M;[�+;p�
;��:�:Z�):?09t꡹h�M��p��Q亙d���0�,�O�)�n���ە�����2?��~��miϻ7�ܻT0�������{��&W�@���4���!�G�&�&K+���/��%4��i8�h�<�7�@�obD��H�rpK���N���Q�jUT���V�_?Y��}[�ͦ]�v�_��a�@d�Af���h���j�)Cm�̰o�y"r�b�t�[w��ny�*�{��;~�(P��ۂ��ܵ���胼���(L���|��d���a������ W��F���/���$V��c�7��q����)������
��Dh�������󜼘 ���>��iQ��1]���f���r������4���rʦ�s����<��σ��BЫ����ro������u��Y��:���1񴼙=��㉷��ո�����h�������  �  0DO=��N=a�M=+PM=�L=�K=�1K=�rJ=�I=-�H=+H=�lG=��F=9F=YE=��D=\ D=-�C=GC=�zB=��A=&iA=e�@=�J@=ʳ?=l?=fv>=��==7+==��<=��;=L6;=)�:=�9=�I9=��8=�8=c7=��6=�!6=�5==�4=tA4=:�3=��2=@J2=ܖ1=N�0=~0=JR/=!�.=��-=��,=�,=)B+=�u*=k�)=��(=�(=�X'=3�&=ϼ%=:�$=��#=C #=�!= � =p�=�d=7=C�=�-=��=�=i=��=��=�'=�N=al=c�
=R�=6�=��=W�=� =��<���<2��<97�<���<j�<���<�z�<��<+��<�$�<��<�z�<=�<c�<k�< Է<4��<���<|��<s��<T_�<E4�<l �<�Ė<���<�>�<D��<鮅<�e�<�8z<q�q<�i<�x`<o�W<�SO<��F<�G><�5<�W-<Z�$<�i</�<�O<C�<���;�(�;�f�;A��;kĬ;2
�;w�;�5p;N;�^,;�N;%��:�o�:K,:�99���r(L�&����{㺮)�o�0���O�L�n�gՆ������ߤ�y������d�ϻ�Fݻow�J=��?��ص��e�X����[���!�u�&��:+�\�/��4��M8��m<�Xi@�O9D��G��@K�KpN�rfQ��%T�޲V�Y�Y[��]�U�_�=�a�b�c�1f�]{h���j��?m�	�o�-+r��t��w�Ԋy���{��`~��c��b���Ȃ�����s(���V�����������������R�������쎼�K������(������������L�KP������ۜ�1	���(���=��sK��*W���e��Zz������æ������9��	���lҫ��$��Vx���ʯ�����j��O������P�������丼},��"r������  �  �AO=M�N=�M=�SM=��L=��K=�9K=`|J=�I=��H=R:H=y}G= �F=RF=xlE=��D=^2D=��C=$C=��B=��A=�rA=�@=Q@={�?=w?=�w>=�==#(==!~<=O�;=k+;=�:=>�9=�99=��8=Y�7=U7=�6=:6=-{5=�4=�?4=��3=>�2=3N2=o�1=E�0=#0=�\/=�.=��-=��,=�",=�T+=؈*=�)=��(=�0(=xh'=��&=��%=!�$=� $=�#=��!=� =��=�c=G= =�%=��==[Y=Q�=��=o=�==�\=�s
=y�=�=�=8�=� =���<c��<(��<NC�<���<�}�<P�<ǖ�<�!�<���<�J�<x��<��<Uc�<O2�<W�<l�<�ڳ<�ů<L��<(��<�k�<f=�<��<#Ɩ<��<�5�<��<���<aL�<F�y<�bq<��h<r5`<G�W<�O<��F<�"><ݲ5<�G-<��$<vk<`�<N`<�<�
�;�t�;���;V�;�B�;闛;��;|q;�PO;+�-;?�;��:���:(�/:r]F9�A��6�I�ׯ��q����`0�!�O��o�;����3���-���ٳ�0»*л��ݻ��껈������S���~�5�����A�!��&��"+��/��3�P#8��<<�m0@�a�C��G���J��"N��Q�s�S�blV���X��[��T]� _���a���c��f��jh���j�a=m��o��:r���t�,>w���y��.|�ޝ~�ƃ��$���悼����>���g��r��������≼����L�����������<���������9��������h���Ϙ�|*��Pw��;���a䝼������B0���?���Q���i�������������5��-����֫��.������ޯ�[4��6���z׳�%��$p������7���A��l��������  �  ==O=��N=�M=�VM=(�L=��K=CK=��J=��I=%I=jMH=ԒG=+�F=�-F=�E=��D=1ID=��C=�$C=��B=,B=�}A=��@=�W@=:�?=A?=*x>=��==#==�u<=��;=�;=or:=k�9=�$9=��8=��7=cB7=�6=&6=fq5=��4=C<4=�3=�2=R2=>�1=�0=	-0=�h/=�.=��-=C-=�8,=l+=�*=��)=^)=�F(= |'='�&=�%=��$=
$=�#=��!=�� =B�=�a=R=��= =��=��=TD=E�=��=s�=�&=�G=�a
=�u=��=ڋ=�=�� =[��<��<H��<�P�<V��<���<�)�<��<J�<���<�z�<�!�<G��<ؓ�<�_�<�6�<��<i��<��<Rī<բ�<Yy�<�F�<Z
�<%Ŗ<�x�<�'�<�Ӊ<m~�<�)�<]�y<�q<@ph<�_<QW<y�N<�ZF<��=<�5<�.-<��$<ti<��<�p<��<�P�;���;
3�;���;��;�K�;�֊;!s;��P;�O/;�!;���:#8�:��4:��V9ZU����F�����A����T50�g�O�f:o�=,������2���|\��g�»�л�b޻���^6���2��
�1�����$�f���!���&��	+��r/�j�3���7� <���?���C�
9G���J�=�M�4�P�{S�"V���X���Z�]�`L_��a��c��f�?Zh�J�j��>m�\�o�dSr�W�t�qw���y�Vx|�4�~�=���`�����e7��]�����Ϡ�����牼:���G������ӎ��+�����Y����f��"Օ��?��N���}���F��v�������t۞�����x��:#���9���V���|��ȭ���ꧼH3������߫��<��
���\����U������� ���O��ՙ��Q߷�P ��W]��*����ϼ��  �  �6O=e�N=u�M=�XM=~�L=� L==LK=֓J=��I=-I=�bH=٪G=[�F=@IF=�E=�D=�bD=�C=&9C=�B=kB=ڈA=��@=�]@=�?=�?=�v>=��==�==�j<=�;=`
;=�\:=��9=�9="h8=K�7=�+7=.�6=��5=�d5=��4=�64=y�3=C�2=�T2=J�1=��0=70=�u/=ϯ.=��-=I-=MQ,=��+=��*=T�)=�))=b_(=�'=ۿ&=��%=C%=S$=7#=�"=I� =�=�]=�=Ǎ=I=y=��=�*=�q=�=��=e=�.=�K
=9c=�t=�=��=@� ==��<@��<���<�]�<��<���<�I�<���<�w�<��<ֱ�<�Z�<W�<���<��<�d�<�=�<M�<C��<�ګ<߳�<c��<�M�<��<���<�m�<��<���<�[�<���<�Ly<!�p<�h<q_<��V<4uN<wF<��=<J\5<�-<��$<�_<��<�|<�<���;�,�;ի�;1�;���;`�;ɵ�;��t;9�R;01;��;�!�:�*�:��9:�h9�#��4�C��`����ງH��!0���O��o�Ut��얻��������yû��ѻ�&߻"F�0���b~��H�x��% �7���s�!�;w&�_�*�S/�s�3���7���;�G�?�AOC���F��*J�.PM�FP��S�_�U��*X�ڊZ�s�\�P_�Va�c��e��Mh��j�GGm���o�Gur�u���w�0Fz���|��P�Aြ��&>���b��D�������y��� ҈�����G���E�������ǎ����.x���ܒ��D��謕�O��-o���Ù�$��M��􀝼ժ���̟��頼����!���C���n������b槼�3��Ƌ��u뫼NP��붮�����~���۲��2�������˶� ���I��H���߲���㼼�  �  �-O=ǕN=��M=�XM=��L=�L=!TK=ӞJ=Q�I=&/I=xH=x�G=wG=�eF=9�E=�E=�}D=�C=�MC=�B='B="�A=��@=Xb@=�?=	?=�s>=��====�]<=�;=��:=�D:=�9=��8=�K8= �7=w7=�{6=�5=�U5=U�4=�.4=ږ3=i�2=�U2=��1=q�0=�?0=��/=G�.=��-=�2-=�j,=%�+=`�*=*=uE)=�x(=g�'=��&=��%=�%=f$= #=�"=�� =��=]W=R�=`�=�=�c=��=�=LS=Q�=A�=�=�=53
=/N=�c=�s=�|=�~ =���<p��<��<Yg�<�<"��<�h�<��<��<F�<���<���<�H�<��<u��<]��<�e�<R=�<q�<o�<���<���<�P�<	�<·�<�]�<'��<ǘ�<�3�<Ѐ<[�x<e/p<;�g<��^<�{V<=N<��E<�e=<�!5<[�,<1�$<N<��<�<L�<9��;G��;� �;��;�F�;�;k��;��v;��T;�$3;��;��:
-�:�>::y9dT���GA�p���M�(&��-0��*P��p��·��f������*���>CĻu`һ��߻�h������A��+� J�fS�'.�(�!��q&���*�X9/�q3���7��~;�HN?���B��mF��I���L�Q�O�i�R��FU�p�W�6<Z�R�\�R�^��0a���c���e�qIh��j�IXm�^�o�ɠr�ENu��w�Νz��5}�H�����,K���s���������������҇�/戼�������]G��"}������'��Rd���'#��/��� ▼{:��O����Ӛ�[��CJ���x������Ġ�硼�
��e3��(d������姼�8��P�������kh���֮��C������w���i��l���N��9B���x��9���fӻ������  �  �"O=�N=��M=dVM=)�L=[L=�YK=��J=��I=�?I=?�H=��G=�,G=��F=}�E=7E=<�D=��C=GaC=��B=�2B=��A=�A=�d@=��?=!?=)n>=6�==}==�N<=Q�;=��:=�+:=�|9=��8=�.8=��7=>�6=hd6=��5=3E5=K�4=1%4=�3=e�2=T2=��1=,�0=�F0=݋/=�.=|.=�G-=�,=��+=,�*=�+*=`)=�(=�'='�&=&&=c%={!$=�#=�"=�� =��=�N=��=9q=#�=M=\�=��=�3=�m=נ=��=�=H
=�7=&Q=~d=q=�u =���<��<x��<�l�<�(�<9��<��<+,�<��<�x�<>"�<���<A��<�:�<���<{��<���<�Z�<�,�<��<#˧<���<�N�<	�<���<�I�<��<�u�<��<>��<rx<ɷo<7g<�^<�V<�M<�UE<=<0�4<�,<�u$<�3<3�<~<V<���;}��;p��;j<�;�;��;�}�;��x;��V;�	5;�;.��:$�:��C:0%�9��z�5?�Ɵ�V�ߺP)��\0��P���p�G7��v헻�[��Rn��Ż�=ӻ������zp��".�}��.J�"{�|w�LF���!�Qu&�v�*�7(/��S3��^7��E;�?�D�B��
F��NI��jL�`O��1R�2�T�:wW�:�Y��\\�g�^��a� qc�	�e�aNh���j��qm��p�Q�r��u�'Ix�_�z�p�}�����S���������_Ƅ�rم��憼������V��)���M���~���������QT��)������2^���������T��e����ۛ�m��EI�� x��+����̡�����'���]��$���ꧼ�A�����������Y����m���ܱ��D�����������<��2x�������Һ�����<���  �  >O=��N=\�M=.RM=W�L=$	L=q]K=��J=C�I=�MI=�H=��G='DG=֚F=�E=�OE=I�D=D=(rC=��B=\<B=��A=�A=�d@=<�?=j?=g>=��==!�<=)?<=ȃ;=��:=k:=b9=�8=�8=�u7=��6=fM6=�5=S45=��4=c4=ه3=��2=�P2=��1=��0=&K0=��/=��.=�.=�Z-=��,=��+=F+=�D*=�w)=��(=�'=#�&=P&=�%=M%$=�#=�"=�� =��=�D=��=a=�=�6=ދ=}�=�=�N=с=�=�= 
=�!=C>=�T=Ld=�k =��<&��<%��<an�<�0�<���<Ĝ�<�K�<��<3��<T�<��<=��<Dl�<�&�<M�<٪�<Is�<+>�<��<Ч<��<DI�<A��<>��<�3�<Iō<`R�<�ބ<�m�<�x<�Do<G�f<�^<�U<�=M<��D<��<<R�4<�v,<�J$<�<0�<�r<�<��;� �;1��;b��;Ά�;b�;�G�;Xyz;}�X;��6;�.;��:�:U�G:�k�9H�q���=�`f����ߺUM���0��Q��Dq�4���-u�������'����ŻcԻ�����5��І�*	����7�����d�"�݀&�Y�*��/��?3��=7�x;���>�QB�S�E���H�[L���N�%�Q�։T�;*W�J�Y��,\��^� a�ic���e�[h���j���m��Fp��s� �u�n�x�U{�N~��L����������W�������z�����G��a��1#���7���W��σ��Ż��t���I�����듼<=��G���ڗ�D#��7h��*����圼����S��@��������颼e���[��8�����tN������D(��ᠭ�e��Ԗ��0���x���ٴ��-���s��a���Eٹ���������6���  �  �O=�{N=?�M=MM=7�L=;L="_K=H�J=J=�XI=4�H=$H=�WG=��F=c	F=�dE=S�D=�D=�C=<�B=eCB=h�A=�A=\c@=��?=�?=�_>=�=="�<=�0<=�r;=]�:=��9=�J9=��8=6�7=�]7=>�6=�86=ɭ5=�$5=v�4=�4=X3=)�2=L2=�1=��0=�M0=6�/=K�.=�&.=�i-=��,=��+=0#+=�Y*=܋)=��(=:�'=�&=�&=�$%=O'$=�#=# "=b� =��=;=��=�R=��=�"=.u=��=j�=�3=�f=Õ=m�=��	=�=�,=F=X=�a =x��<շ�<X��<�l�<X5�<��<��<1e�<�<���<�}�<S/�<���<r��<�K�<��<)ĸ<��<�J�<-�<"ѧ<^��<OA�<��<]��<��<"��<�1�<Q��<;B�<N�w<��n<�3f<+�]<{5U<6�L<L�D<*~<<5_4<�B,<9 $<0�<��<�b<� <��;�%�;��;��;� �;���;U��;��{;��Y;/8;��;a�:ˆ�:+�J:�<�9.�k�Z�<��I��w!�τ��1��Q�k�q����(�2����̷�{�ƻ��Ի�u�_}ﻓ���$��p	�y����_��w���"���&�e�*�`/�43�$&7���:�,�>�B�miE���H�7�K�b�N��~Q�T@T�k�V��Y��\�(�^�;�`�hc�j�e��kh��k���m��pp� <s�1v���x�*�{��[~�{|��Ǽ���킼o���#���,��5/���.���/��7��]G��c��Y���)��������A������5ד��"���l������0����=��-�����������6��co��@����ߢ�e���\���������;\���Ȫ��>��#����<��2���16������0
���^��P����ڸ�����"���;���R���  �  O=�sN=��M="HM=�L=�L=�_K=�J=7J=�`I=��H=�H=;fG=p�F=fF=tE=��D=,D=��C=o�B=HB=��A=�A=aa@=��?=�?=�X>=��==�<=�$<=	e;=Ӧ:=��9=:89=c�8=��7=�J7=s�6=�(6=7�5=!5=��4=�4=�w3=!�2=�G2=N�1=��0=�N0=��/=B�.=N/.=�t-=ѷ,=r�+=�2+=�i*=̚)=��(=f�'=�'=�&=(%=�'$=>#=��!=� =��=~2=b�=�F=��=�=Bc=�=��=:=ZQ="�=�=��	=��==:=�M=ZY =p��<T��<���<Ij�<F7�<N��<ǻ�<�w�<�0�<���<ܜ�<P�</�<<��<\g�<	�<%ָ<ْ�<?R�<7�<Ч<���<�8�<0ߚ<�z�<5�<˓�<4�<���<��<*\w<p�n<D�e<�T]<��T<�L<�eD<ED<<%-4<�,<�#<��<��<sS<�<>!�;�;�;�I�;�R�;�Z�;�c�;�n�;2�|;[;C9;��;���:�:�/M:���9��g��l<�R���d�i��2[1���Q�6zr�Pc��uY������O��� ǻdջ����m��A�T�	����v
�	��q��h1"���&��*�!/��.3�)7���:��r>�3�A�43E��_H�2oK�CdN��AQ��	T���V��]Y�,�[��q^���`��jc���e��|h��k�t�m�'�p�qfs��?v�Uy���{�/�~����iぼ-���4��GF��pL��K���F��]D��H��9U��#n������Î�e���&>������fɓ�����T��o���Kۘ�����_������᝼*!��1_��S����٢����_��M���>���h��ت��Q��sҭ��V�� ڰ�zW���ʳ�40������sʷ�����^%��A��V��Di���  �  ��N=tnN=O�M=�DM=S�L=:L=a_K=J�J=<J=BeI=��H=�H=oG=�F=O#F=�}E=:�D=v3D=��C=��B=�JB=��A=UA=�_@=.�?=�?=T>=�==c�<= <=\;=ќ:=��9=},9=28=��7=�>7=�6=6=͕5=�5=u�4=x 4=�r3=��2=hD2=�1=��0=O0=��/=��.=�4.=�{-=�,=� ,=�<+=Cs*=�)=��(='�'=�'= &=�)%= ($=�#=��!=T� =6�=�,=��=�>=l�=H=�W=��=��=�=�C=t=ɡ=��	=��==22=G=�S =��<��<���<�g�<�7�<v �<���<��<T?�<��<���<Ld�<4�<���<	x�< +�<��<H��<GV�<�<=Χ<W��<�2�<�֚<p�<���<���<��<ą�<�	�<@,w<�]n<��e<v!]<жT<lL<�;D<�<<>4<[�+<��#<.�<�<>H<��<��;�G�;Xd�;�{�;���;��;໏;��};P�[;�9;#;���:E�:,�N:�g�9(ne��G<�ri��R�����3�1��DR���r��������{R��ä���{ǻ�ջ�k�+m�.����=���	�K�7&�s���
A"��&�$�*�g$/��,3��7��:�]>�s�A�E��:H��GK��<N�kQ�"�S��V��GY���[�pi^���`�}nc���e�0�h�-k�s�m��p���s��`v�n=y��|�D�~�޹�������,��6L��u\���`��&]���V��R���S���^���u��똍�)ǎ�����<��~���������E��M���pȘ��	��8L������ѝ�'��]U��啡��֢�$��Db��4������q���⪼T^��V᭼�g��n��l���᳼TH��L����ⷼ(���:���T��~g��gx���  �  v�N=~lN=��M=VCM=[�L=�L=L_K=��J=#J=�fI=�H=OH=/rG=`�F=�&F=ـE=:�D=�5D=��C=&�B=mKB=ѨA=(A=
_@=&�?=�?=TR>=�==#�<=p<=Y;=V�:=��9=m(9=�z8=P�7=�:7=�6=r6=��5=�5=�4=_�3=�p3=��2=<C2=:�1=D�0=#O0=�/=��.=<6.=�}-=��,=�,=�?+=�v*=�)=��(=i�'=�'=)!&=7*%=�'$=Y#=��!=�� =��=�*=/�=�;=J�=�=�S=c�=�=)=Y?=�o=��=��	=Z�==�/=�D=�Q =*��<���<��<cg�<^8�<��<3��<چ�<aD�<"��<���<Ak�<�<[��<�}�<w/�<C�<Z��<>W�<�<Aͧ<g��<0�<�Ӛ<l�<���<]�<j��<�~�<��<Xw<cLn<��e<�]<�T<B\L<�-D<+<<~4<Z�+<��#<��<��<�D<.�<� �;iL�;Rm�;���;���;���;�֏;��};��[;�%:;UX;�F�: /�:%�N:��9D�d��F<��x��A��k�}�1��cR�2�r���������Kn��{ø�I�ǻ��ջ���3�������L���	��"��/��
�+���F"�t�&�O�*��%/�&,3��7�e�:� V>�9�A��E�.H�::K� /N��Q���S�|�V��@Y�%�[�g^�+�`��oc��e���h��2k���m�W�p�"�s��kv�?Jy�u|��~��u��5��\T��6d���g��dc��
\���V���W��Wb���x��	����Ȏ����<���|��v��� ��A��[����������E�������̝����5R����բ�2��:c���������t���檼�b��c歼�m�����Rt���鳼�P��զ��뷼:���B��\[��m���}���  �  ��N=tnN=O�M=�DM=S�L=:L=a_K=J�J=<J=BeI=��H=�H=oG=�F=O#F=�}E=:�D=v3D=��C=��B=�JB=��A=UA=�_@=.�?=�?=T>=�==c�<= <=\;=ќ:=��9=},9=28=��7=�>7=�6=6=͕5=�5=u�4=x 4=�r3=��2=hD2=�1=��0=O0=��/=��.=�4.=�{-=�,=� ,=�<+=Cs*=�)=��(='�'=�'= &=�)%=($=�#=�!=Z� =>�=�,=��=�>=��=e=�W=ٜ=��=�=/D=mt="�=��	=$�=�=�2=�G=%T =��< ��<���<�h�<�8�<:�<7��<~��<�?�<^��<*��<Vd�<�<���<�w�<�*�<^�<���<~U�<=�<Wͧ<j��<�1�<�՚<=o�<���<���<�<;��<Q	�<�+w<�]n<��e<�!]<[�T<�lL<�<D<�<<�4<��+<w�#<�<d�<"J<��<�#�;K�;Gg�;M~�;���;���;꼏;��};�[;��9;� ;���:�ܩ:�yN:y4�9��e��f<��y��V�ຝ��ܢ1�MR���r�����à���U����~ǻ��ջ�m�&o������>�~�	����&���+��GA"�5�&�L�*��$/��,3�7��:�]>�}�A�&E��:H��GK��<N�nQ�$�S��V��GY���[�pi^���`�}nc���e�0�h�-k�s�m��p���s��`v�n=y��|�D�~�޹�������,��6L��u\���`��&]���V��R���S���^���u��똍�)ǎ�����<��~���������E��M���pȘ��	��8L������ѝ�'��]U��啡��֢�$��Db��4������q���⪼T^��V᭼�g��n��l���᳼TH��L����ⷼ(���:���T��~g��gx���  �  O=�sN=��M="HM=�L=�L=�_K=�J=7J=�`I=��H=�H=;fG=p�F=fF=tE=��D=,D=��C=o�B=HB=��A=�A=aa@=��?=�?=�X>=��==�<=�$<=	e;=Ӧ:=��9=:89=c�8=��7=�J7=s�6=�(6=7�5=!5=��4=�4=�w3=!�2=�G2=N�1=��0=�N0=��/=B�.=N/.=�t-=ѷ,=r�+=�2+=�i*=˚)=��(=f�'=�'=�&=(%=�'$=D#=��!=$� =�=�2=~�=�F=մ=�=�c=o�=�=�=�Q=��=��=��	=��=�=�:=�N=QZ =a��<>��<g��<l�<�8�<���<��<�x�<�1�<s��<3��<P�<��<ǳ�<�f�<�<�Ը<~��<�P�<��<GΧ<���<,7�<nݚ<�x�<�	�<_��<��<���<�<[w<ߏn<=�e<U]<�T<��L<�gD<�F<<�/4<�,<��#<b�<��<W<��<(�;*B�;�O�;�W�;�^�;�f�;�p�;�|;�[;z@9;��;���:�:�M:6!�9ah�z�<��q��`��"���k1�uR�*�r��j���`�����V��J&ǻiջ:㻰��p������	����K�������1"�X�&�d�*�>!/��.3�P7��:��r>�F�A�C3E��_H�;oK�JdN��AQ��	T��V��]Y�.�[��q^���`��jc���e��|h��k�u�m�'�p�qfs��?v�Uy���{�/�~����iぼ-���4��GF��pL��K���F��]D��H��9U��#n������Î�e���&>������fɓ�����T��o���Kۘ�����_������᝼*!��1_��S����٢����_��M���>���h��ت��Q��sҭ��V�� ڰ�zW���ʳ�40������sʷ�����^%��A��V��Di���  �  �O=�{N=?�M=MM=7�L=;L="_K=H�J=J=�XI=4�H=$H=�WG=��F=c	F=�dE=S�D=�D=�C=<�B=eCB=h�A=�A=\c@=��?=�?=�_>=�=="�<=�0<=�r;=]�:=��9=�J9=��8=6�7=�]7=>�6=�86=ɭ5=�$5=v�4=�4=X3=)�2=L2=�1=��0=�M0=6�/=K�.=�&.=�i-=��,=��+=/#+=�Y*=܋)=��(=:�'=�&=�&=�$%=U'$=�#=. "=r� =�=";=��=�R=��=#=�u=�=��=24=^g=��=`�=��	=�=*.=gG=]Y=Cc =6��<���<���<}o�<�7�<,��<��<�f�<P�<���<~�<o/�<Q��<̔�<�J�<��<�¸<*��<fH�<��<�Χ<؊�<�>�<g�<���<��<��<�/�<ݶ�<A�<åw<�n<�3f<�]<�6U<j�L<,�D<��<<<c4<#G,<%$<>�<�<h<�<�(�;�.�;�%�;��;o�;��;.�;*�{;:�Y;e+8;�~;���:sm�:�J:���9}�l�*2=��v���O�u��-1�8�Q��r�]��M�������Zշ�O�ƻ��Ի�{�ǂ�?���#���q	����C��Y��C���"�<�&���*��/�[43�[&7��:�N�>� B��iE���H�D�K�l�N��~Q�Z@T�o�V��Y��\�*�^�=�`� hc�k�e��kh��k���m��pp� <s�1v���x�*�{��[~�{|��Ǽ���킼o���#���,��5/���.���/��7��]G��c��Y���)��������A������5ד��"���l������0����=��-�����������6��co��@����ߢ�e���\���������;\���Ȫ��>��#����<��2���16������0
���^��P����ڸ�����"���;���R���  �  >O=��N=\�M=.RM=W�L=$	L=q]K=��J=C�I=�MI=�H=��G='DG=֚F=�E=�OE=I�D=D=(rC=��B=\<B=��A=�A=�d@=<�?=j?=g>=��==!�<=)?<=ȃ;=��:=k:=b9=�8=�8=�u7=��6=fM6=�5=S45=��4=c4=ه3=��2=�P2=��1=��0=%K0=��/=��.=�.=�Z-=��,=��+=F+=�D*=�w)=��(=�'=$�&=S&=�%=T%$=�#=�"=	� =Ә=E=#�=�a=j�=A7=V�=�==�O=��=�=9�=Y
=%#=�?=iV=�e=�m =k��<y��<^��<qq�<�3�<c��<��<�M�<���<?��<�T�<��<��<zk�<�%�<��<Ө�<�p�<�;�<��<ͧ<��<*F�<5��<S��<1�<�<;P�<�܄</l�<�x<�Co<;�f<�^<әU<[@M<S�D<��<<@�4<,|,<tP$<�<��<�x<�<f�;��;��;��;Ǎ�;dg�;{K�;�|z;҆X;�6;I&;��:�a�:z_G:Z��9{s��(>�S����.�Kj���0�h!Q�I`q�e�������)	��12����Ż�Ի"�ỡ���:��C��*,	�a��������e��"���&���*� /�P@3�>7��;���>�:QB�m�E���H�kL���N�/�Q�މT�A*W�N�Y��,\��^� a� ic���e�[h���j���m��Fp��s� �u�n�x�U{�N~��L����������W�������z�����G��a��1#���7���W��σ��Ż��t���I�����듼<=��G���ڗ�D#��7h��*����圼����S��@��������颼e���[��8�����tN������D(��ᠭ�e��Ԗ��0���x���ٴ��-���s��a���Eٹ���������6���  �  �"O=�N=��M=dVM=)�L=[L=�YK=��J=��I=�?I=?�H=��G=�,G=��F=}�E=7E=<�D=��C=GaC=��B=�2B=��A=�A=�d@=��?=!?=)n>=6�==}==�N<=Q�;=��:=�+:=�|9=��8=�.8=��7=>�6=hd6=��5=3E5=K�4=1%4=�3=e�2=T2=��1=,�0=�F0=܋/=�.={.=�G-=�,=��+=+�*=�+*=
`)=�(=��'=(�&=)&=g%=�!$=�#=�"=�� =�=O=��=~q={�=�M=�=J�=�4=�n=ܡ=�=M�=�
=R9=�R=>f=�r=�w =���<���<��<Bp�<�+�<��<���<E.�<���<�y�<�"�<���<��<�9�<t��<���<���<7X�<�)�<���<�ǧ<5��<�K�<���<A��<�F�<"ߍ<^s�<��<���<px<��o<*g<�^<�	V<�M<�YE<�=<��4< �,<@|$<�:<C�<�<<<��;���;f��;�E�;���;���;���;D�x;�V;�5;��;F��:~�:vBC:�d�9!�|���?�e���=ພI�}0��P�S�p��E��P���ch�� z��/ŻvGӻK��_���v���0����L��|��x�dG�l�!�	v&�
�*��(/�1T3�,_7�/F;�2?�i�B�F��NI��jL�#`O��1R�;�T�@wW�?�Y��\\�j�^��a�"qc�
�e�bNh���j��qm��p�R�r��u�'Ix�_�z�p�}�����S���������_Ƅ�rم��憼������V��)���M���~���������QT��)������2^���������T��e����ۛ�m��EI�� x��+����̡�����'���]��$���ꧼ�A�����������Y����m���ܱ��D�����������<��2x�������Һ�����<���  �  �-O=ǕN=��M=�XM=��L=�L=!TK=ӞJ=Q�I=&/I=xH=x�G=wG=�eF=9�E=�E=�}D=�C=�MC=�B='B="�A=��@=Xb@=�?=	?=�s>=��====�]<=�;=��:=�D:=�9=��8=�K8= �7=v7=�{6=�5=�U5=U�4=�.4=ٖ3=i�2=�U2=��1=q�0=�?0=��/=F�.=��-=�2-=�j,=$�+=_�*=*=tE)=�x(=g�'=��&=��%=�%=m$=,#=�"=�� =��=�W=��=��=^�=9d=�=o=T=;�=O�=P�=9=�4
=�O=�e=pu=�~=�� =���<F��<Ѩ�<�j�<X�<��<~k�<�	�<���<MG�<���<��<XH�<��<��<w��<�c�<�:�<g�<$�<6��<O��<M�<��<e��<�Z�<P��<M��<t1�<�΀<-�x<D.p<.�g<��^<�}V<YN<÷E<�j=<H'5<��,< �$<8U<��<S�<q<���;��;+,�;��;O�;%�;t��;n�v;9�T;r3;-�;l�:&	�:��>:��w9 2����A�|�����ບG�EO0��KP��&p�އ�u���Ħ�b���NNĻ[jһ�໽����������.��K��T�H/��!�Gr&���*��9/�wq3��7�8;�xN?���B��mF��I���L�_�O�t�R��FU�v�W�;<Z�W�\�U�^��0a���c���e�rIh��j�JXm�_�o�ɠr�ENu��w�Νz��5}�H�����,K���s���������������҇�/戼�������]G��"}������'��Rd���'#��/��� ▼{:��O����Ӛ�[��CJ���x������Ġ�硼�
��e3��(d������姼�8��P�������kh���֮��C������w���i��l���N��9B���x��9���fӻ������  �  �6O=e�N=u�M=�XM=~�L=� L==LK=֓J=��I=-I=�bH=٪G=[�F=@IF=�E=�D=�bD=�C=&9C=�B=kB=ڈA=��@=�]@=�?=�?=�v>=��==�==�j<=�;=`
;=�\:=��9=�9="h8=K�7=�+7=.�6=��5=�d5=��4=�64=x�3=C�2=�T2=I�1=��0=
70=�u/=ί.=��-=H-=MQ,=��+=��*=S�)=�))=a_(=�'=ܿ&=��%=G%=Z$=B#=�"=`� =$�=�]=H�=�=�=|y=�=�+=~r=Ү=��=�=0=RM
=�d=�v=Ă=��=� =���<���< ��<%a�<��<���<'L�<���</y�<��<���<�Z�<��<���<���<�b�<�;�<��<S��<g׫<���<�<J�<^�<l��<�j�<�<F��<�Y�<	��<�Jy<
�p<�h<r_<��V<4xN<cF<��=<�a5<�-<�$<�f<��<�<��<���;�8�;ζ�;�'�;P��;J�;���;`�t;z�R;+1;=�;��:;�:%`9:єf9����*YD�ٝ��}*��h�&B0�ZP��o��������^+�����g�û&�ѻZ/߻�M컓������J�i���!�k8���W�!��w&���*�{S/�і3�ѻ7��;�u�?�fOC���F��*J�?PM�FP��S�g�U��*X�ߊZ�w�\�S_�Va�Ěc��e��Mh��j�GGm���o�Gur�	u���w�1Fz���|��P�Aြ��'>���b��D�������y��� ҈�����G���E�������ǎ����.x���ܒ��D��謕�O��-o���Ù�$��M��􀝼ժ���̟��頼����!���C���n������b槼�3��Ƌ��u뫼NP��붮�����~���۲��2�������˶� ���I��H���߲���㼼�  �  ==O=��N=�M=�VM=(�L=��K=CK=��J=��I=%I=jMH=ԒG=+�F=�-F=�E=��D=1ID=��C=�$C=��B=,B=�}A=��@=�W@=:�?=A?=*x>=��==#==�u<=��;=�;=or:=k�9=�$9=��8=��7=cB7=�6=&6=fq5=��4=C<4=�3=�2=R2==�1=�0=-0=�h/=�.=��-=B-=�8,=l+=�*=��)=])=�F(= |'=(�&=�%=��$=
$=�#=��!=�� =]�=�a=�=٘=N=�=3�=�D=�=v�=\�=�'=I= c
=�v=	�=m�=��=M� =���<c��<���<T�</��<>��<,�<̻�<�K�<���<{�<�!�<���<��<|^�<�4�<��<��<�ݯ<x��<ӟ�<Bv�<|C�<O�<;<Gv�<6%�<�щ<�|�<k(�<z�y<�
q<5ph<��_<�RW<)�N<O^F<:�=<��5<g4-<��$<�o<5�<�v<!�<Y\�;���;�<�;��;��;�P�;0ڊ;W s;&�P;`K/;I;���:�:�E4:TKU9}���;G�����6����FR0���O��Uo�j9���������g����»��л�j޻+��<��k5������B%�a���!�B�&�J
+�_s/���3���7�7 <���?��C�$9G�J�M�M�@�P� {S�*V��X���Z�]�cL_��a��c��f�@Zh�K�j��>m�]�o�eSr�W�t�qw���y�Vx|�4�~�=���`�����e7��]�����Ϡ�����牼:���G������ӎ��+�����Y����f��"Օ��?��N���}���F��v�������t۞�����x��:#���9���V���|��ȭ���ꧼH3������߫��<��
���\����U������� ���O��ՙ��Q߷�P ��W]��*����ϼ��  �  �AO=M�N=�M=�SM=��L=��K=�9K=`|J=�I=��H=R:H=y}G= �F=RF=xlE=��D=^2D=��C=$C=��B=��A=�rA=�@=Q@={�?=w?=�w>=�==#(==!~<=O�;=k+;=�:=>�9=�99=��8=Y�7=U7=�6=:6=-{5=�4=�?4=��3==�2=3N2=n�1=E�0=#0=�\/=�.=��-=��,=�",=�T+=׈*=~�)=��(=�0(=yh'= �&=��%=%�$=� $=�#=��!=)� =ͩ=d=o=��=�%=�=e=�Y=ޤ=Y�=-=�>=�]=�t
=��=H�=T�=��=Q� =���<��<ʓ�<�E�<��<��<'�<R��<�"�<���<K�<���<ԡ�<�b�<M1�<��<��<�س<�ï<���<���<oi�<�:�<Q�<�Ö<�}�<�3�<��<��<BK�<��y<bq<��h<,6`<��W<�O<��F<x&><�5<QL-<h�$<�p<��<ze<��<R�;�}�;���;J�;{H�;>��;��;q;PO;q�-;d�;O��:?v�:�/:dCE9�ޘ� 
J��ܣ���⺪���w0�`�O�o����>��D7��-⳻�7»1л��ݻB��5��������A��d��������!���&�Y#+�q�/�J�3��#8��<<��0@�|�C���G���J��"N��Q�{�S�ilV���X��[��T]�#_���a���c��f��jh���j�b=m��o��:r���t�,>w���y��.|�ޝ~�ƃ��$���悼����>���g��r��������≼����L�����������<���������9��������h���Ϙ�|*��Pw��;���a䝼������B0���?���Q���i�������������5��-����֫��.������ޯ�[4��6���z׳�%��$p������7���A��l��������  �  0DO=��N=a�M=+PM=�L=�K=�1K=�rJ=�I=-�H=+H=�lG=��F=9F=YE=��D=\ D=-�C=GC=�zB=��A=&iA=e�@=�J@=ʳ?=l?=fv>=��==7+==��<=��;=L6;=)�:=�9=�I9=��8=�8=c7=��6=�!6=�5==�4=tA4=:�3=��2=@J2=ܖ1=M�0=~0=JR/=!�.=��-=��,=�,=)B+=�u*=j�)=��(=�(=�X'=3�&=м%=<�$=��#=I #=�!=� =��=�d=S=g�=�-=ޥ=�=pi=�=O�=(=�O=m= �
=�=�=��=H�=� =��<���<��<�8�<���<�k�<���<�{�<x�<Ǝ�<�$�<)��<�z�<�<�<��<w�<�ҷ<ؿ�<��<֙�<��<�]�<{2�<���<LÖ<&��<,=�<��<⭅<3e�<�7z<�q<�i<Cy`<z�W<~UO<��F<J><��5<�Z-<��$<pm<��<�S<֩<f��;%/�;5l�;,��;tȬ;C�;y�;�7p;�N;"\,;�I;/��:�]�:��+:GQ89�z��~dL��٤�ʜ�e:�$�0�j�O�8�n�݆�$���椻4��h���V�ϻAKݻB{껙@��������f�/��f���o�!�ԧ&�;+���/��4��M8��m<�qi@�b9D��G��@K�TpN�zfQ��%T��V�Y�
Y[��]�W�_�>�a�c�c�1f�^{h���j��?m�	�o�-+r��t��w�Ԋy���{��`~��c��b���Ȃ�����s(���V�����������������R�������쎼�K������(������������L�KP������ۜ�1	���(���=��sK��*W���e��Zz������æ������9��	���lҫ��$��Vx���ʯ�����j��O������P�������丼},��"r������  �  qEO=\�N=��M=�MM=T�L=��K=;,K=lJ=ݨI=k�H=>!H=�aG=�F=�E=�LE=��D=�D=��C=��B=rB=>�A=�bA=$�@=wF@=j�?=?=+u>=��==�,==�<=��;=�<;=!�:=�9=qS9=ٰ8="8=�k7=6�6=j'6=�5=��4=3B4=��3=�2=OG2=��1=z�0=�0=oK/=&}.=��-=��,=s,=m6+=�i*=M�)=��(=�(=�N'=F�&=��%=��$=!�#=��"=��!=�� =2�=�d=�=��=�2=|�==�r=��=\ =3=�Y=\v=�
=u�=��=\�=}�=�� =)��<���<��<�/�<(��<�]�<���<i�<���<�w�<��<��<�a�<s$�<���<�ֻ< ��<^��<П�<ʍ�<�u�<�U�<y,�<��<V<P��<�B�<S��<���<u�<�\z<I�q<�8i<j�`<�X<*wO<��F<v_><Y�5<~b-< �$<Pi<��<;F<O�<���;��;-�;�O�;�u�;X��;��;�go;�-M;��+;�
;Y
�:��:�):��/9�#��}�M�L���V$�@m�=�0���O�g�n��Ɔ��ޕ�"���[B������kϻ{�ܻO2껜���ȭ����W����`�����!�x�&�NK+���/��%4��i8�w�<�D�@�ybD��H�xpK���N���Q�mUT���V�a?Y��}[�Φ]�w�_��a�@d�Af���h���j�)Cm�̰o�y"r�b�t�[w��ny�*�{��;~�(P��ۂ��ܵ���胼���(L���|��d���a������ W��F���/���$V��c�7��q����)������
��Dh�������󜼘 ���>��iQ��1]���f���r������4���rʦ�s����<��σ��BЫ����ro������u��Y��:���1񴼙=��㉷��ո�����h�������  �  lXO=��N=:N=TcM=��L=��K=8K=SpJ=��I=��H=�H="?G=�~F=3�E=�E=,�D=��C=(lC=\�B=�rB=��A=�|A=��@=,r@=��?=NJ?=�>=�>=�h==�<=�$<=��;=��:=EI:=Q�9=\9=Pl8=u�7=x*7=^�6=��5=�M5=C�4=�4=�m3=��2=a2=�X1=&�0=�/=��.=� .=+J-=v,=�+=U�*=�*=#b)=��(=��'=QA'=��&=�%=��$=��#= #=L�!=}� =I�=)0=��=T=+�=s6=�=
�= =�;=�W=�g=$n=�m	=�g=�]=�O=&<=�C�<���<7��<o9�<H��<�(�<̌�<���<KM�<��<p2�<��<g�<�$�<���<�߻<"Է<�ϳ<�̯<�ī<���<���<�n�<*;�<���<���<�w�<�1�<��<"��<Ÿz<�r<}i<��`<#!X<DoO<[�F<�><%�5<��,<�t$<"�<�R<٤
<\�<���;���;А�;�5�;�٨;���;��;\�e;��B;�� ;
g�:��:�}:{ :��_7(��;du�aS���Z�� ��+�;��A[���z��ጻ`,��0��9湻MOȻ�iֻ�0�D�������ե��j�=���)��-!� &��*�0:/��3�k8�Uc<��@���D�t�H�I-L�ٓO���R�>�U�?X��jZ�	�\�|^�-Z`��0b�Gd���e�yh�~(j�dl��n�*q�ks��u��x�nz���|�'�謀��؁�����8��Wj��<��� ȇ���q"���T�������׍�//��җ��A��B����!�������5��T������Kg��ʟ������͟��ɠ�z���׬��g���������=ʦ������2��'x��Lë�B��?\��ԥ���찼�2��@y��7´�����[�����������C��ꋼ��  �  dXO=7�N=sN=eM=	�L=o�K=�:K=�sJ=R�I=�H=FH=SDG=p�F=�E=�%E=��D=�C=CqC=��B=�vB=��A=�A=��@=�t@=��?=�K?=�>=L>=�h==�<=�"<=E�;=F�:=E:=�9=�9=h8=��7=]'7=�6=4�5=WM5=~�4=�4=Lo3=|�2=�2=�[1=%�0=v�/=��.=%.=	O-=c{,=��+=1�*=�"*=�g)=H�(=|�'=�E'=R�&=I�%=]�$= $=�#=��!=�� =ڃ=0=��=7R=u�=�2=j�=�=�=�6=�R=5c=j=�j	=f=�\=FO=\<=HE�<�<w��<�=�<U��<�.�<���<]��<�V�<���<�=�<0��<=s�<�0�<2�<+�<�ݷ<[س<Kԯ<�˫<<��< ��<�s�<�>�<� �<n��<�v�</�<�<���<Y�z<sr<
ji<�`<X<�_O<�F<�><1�5<��,< u$<��<�V<��
<s�<���;���;���;BV�;��;;o��;��e;�;C;XD!;u ;�=�::0M:!\�7����xt�c븺����o���x;�%-[���z�y䌻�6��[A������mȻ��ֻ�Q�������z��ݭ��o����U(��)!���%�	�*��0/��3�	8��U<�s�@�:�D��qH��L��|O�՛R�rrU�NX�jUZ�(s\�pj^��J`�#b�d���e�q�g�� j�L^l�!�n��q�ms�K�u�#&x�zz���|�&�ȵ���ၼ!�� @���o��,���]ʇ�V����!���R�������Ӎ�~*��F���
��3����������v+��j����
��f[�����~�����������_���ޚ��=�������Ʀ����70���v��+ë����u_������V󰼐:��쁳�#˴�����c��v�������G�������  �  �WO=��N=�N=�iM=ֹL=KL=�BK=�|J=��I=.�H=�H=[SG=��F=��E=�6E=ęD= D=�C=2�B=��B=�B=��A=\A=0{@=h�?=AP?=�>=d>=�g==��<=�<=�y;=��:=�8:=ƙ9=��8=b[8=H�7=7=-�6=��5=TK5=��4=�4=�r3=��2=�2=�b1=w�0=�/=�/=�1.=]-=��,=�+=�*=�3*=!x)=��(=v
(=�Q'=2�&=��%=J�$=�$=�#=:�!=�� =�=T/=��=�L=I�=5(=�~=��=��=�'=�D=�V=�_=�b	=g`=�Y=GN=>==AJ�<��<���<5J�<���<#A�<���<j�<ls�<#��<�_�<���<��<�R�<*$�<��< ��<+�<T�<Bޫ<eʧ<㪣<�~�<G�<��<���<Xr�<N%�< ؅<q��<�wz<\�q<I1i<9�`<<�W<�2O<��F< �=<qr5<f�,<�u$<��<e<c�
<��<�/�;�.�;� �;���;�n�;8?�;�B�;,g;VbD;Lh";h.;;M�:�f�:��:�K�7�(�Or�dܷ�����R��1;�2[���z�X����\��j{��iK��p�Ȼ��ֻ����p��z����������%��!���%���*�9/��3���7�.<�8Y@�D`D��8H���K��:O�LWR��-U���W��Z��9\�N7^�H`���a�
�c�t�e�Z�g�!j��Nl��n�
q��ss���u��@x�/�z�J�|�HK�bЀ�����(���U�����t����ч��������#M��$����ȍ�v�����w����y��b��y���P��Ʉ���隼.9��r���F���~����������������� ���/����ꧼp)��9s���ë����~i����������Q�������崼z0���{��~Ÿ����Q��;����  �  DVO=,�N=�N=�oM=��L=L=�NK=p�J=��I=��H=�.H=�jG=߭F=g�E=�QE=�D=� D=ӖC=�C=o�B="B=ƕA=�A=��@=�?= V?=s�>=/>=Ke==��<=�<=)l;=��:=.%:=q�9=�8=�F8=ة7=�7=ru6=��5=SG5=�4=Q4=�w3=R�2=[$2=m1=��0=d�/==/=�D.=�r-=��,=��+=�+="N*=��)=��(=
 (=e'=��&=q�%=��$=P$=4#=��!=� =�=@-=�=C=��=�=�i=��=k�=@=-=B=�N=UU	=�V=�S=�K=�==QP�<�<���<c\�<>��<�\�<���<04�<���<U�<4��<�&�<���<{��<�U�<�4�<� �<��<X�<��<��<V��<S��<�Q�<�<���<qi�<+�<e��<,i�<�(z<"q<x�h<�,`<+�W<'�N<�UF<��=<vU5<��,<)t$<��<�w<��
<<Ȇ�;��;N�;)N�;O�;g�;��;�h;�/F;31$;~�;~�:kN�:��	:M�C8� ��n�W������%��I�:��Z���z����h���ޫ�Bʺ�U\ɻ��׻�[�'��E��������#��� ��%��!�`�%�Yq*���.��]3�H�7�V�;�W@�D���G��xK��N�3�Q���T��XW�v�Y�s�[���]�3�_�+�a���c��e�¿g���i�z:l�:�n��
q�_�s�V�u��mx�3�z��>}���s����&���P��}x��v���:����އ�n�������F��y��Ĺ���
��"m���ޑ��[��Cߔ�(c��&ᗼPS��>������=��b�� u���y��v���o��Sl��rr�����������ݧ�� ���o��:ƫ�~ ���z���ү�'���w���ų����Z�����m渼'���c�������  �  RRO=*�N=
N=�uM=P�L=�L=�[K=k�J=��I=7I=�HH=�G=��F=F=�sE=[�D=e@D=~�C=�,C=B�B=�(B=�A=!A=֎@=��?=z[?=�>=[>=g`==1�<=�<=Y;=V�:=�
:=�g9=�8=
+8=�7=��6=�d6=R�5=f@5=��4=u4=|3=�2={-2=�x1=��0=M�/=c*/=r\.=΍-=��,=��+=.1+=�o*=�)=��(=;(=u|'=I�&=��%=
%=�$=#=>�!=�� =o�=�(=�=05=��=��=�M=��=��=��=�=z&=T7=�B	=:I= K=>G=�<=~T�<v�<{��<Wp�<E��<M}�<���<=d�<;��<vQ�<��<�k�<�<o��<3��<Lm�<^R�<�>�<�,�< �<5��<ӣ<���<�[�<��<��<MZ�<���<���<�;�<��y<	q<�Zh<��_<TW<�N<�F<��=<�)5<r�,<�j$<�<w�<�
<+D<���;�;��;>�;���;���;�&�;�k;�|H;Uv&;	;��:��:PG:��8a�ع��j�C����i��)H�X~:�ιZ���z��R��*���h���w���%ʻ�hػ9�ʏ�+1 �,U��1�;�����,�h!���%��S*���.��-3�z7���;���?���C��rG�]�J��ON��cQ��9T�!�V��:Y��r[���]�q�_��{a�:tc��{e���g���i�	(l��n�dq��s��&v���x�`,{��}�w��5��-`������진��ą��܆���.��Q!�� B���n����������T��|����7��e���B1����������r��a��������!���9��E��H���H���K��|W��p��P���-ѧ�����n��.ͫ�^0��*�������
S��&��������J��5���ַ�E��"K��6~�������  �  @KO=f�N=�N=�yM=��L=< L=+hK=N�J=��I=t&I=�eH=ƨG=��F=BF=d�E=�D=�cD=c�C=�HC=��B=�;B=-�A=�(A=��@=�?=�^?=+�>=�	>=JX==�<=)�;=LA;=̓:=h�9=�E9=E�8=�	8=�r7=��6=P6=��5=65=��4=�4=�}3=��2=52=Ԃ1=&�0=a0=�?/=v.=��-=s�,=`,=5W+=ו*=��)=G)=�X(=ԕ'="�&=:�%=�%=�#$=,#=g "=�� =́=� =M�=#=݉=��=%,={j=��=�=��==�=A+	=M7=C>=/?=�8=ZS�<�!�<���<���<�<���<��<���<�<��<�"�<���<�`�<��<���<���<��<�k�<R�<6�<��<��<�<a�<r�<��<CD�<Gى<�m�<��<<y<6{p<�g<C"_<E�V<�N<ŝE<�?=<l�4<3�,<�U$<��<"�<	<�d<G�;���;��;�ν;�;��;X�;��m;�K;[);��;,��:y�:�&:`^�81	Ϲ �f�U���2� ��J:���Z�+{� ���儝�i���M���˻�oٻ�D�K���˥ ����V��=�4>��?�!��%�/=*�ʪ.��3��A7�)g;��k?�\IC�&�F��uJ�߻M���P���S��@V��X�-�Z��]��._��4a�v<c��Pe�Pzg���i�	l�\�n��'q���s�Gbv���x�d�{��~��G���z��6���~ǃ��ᄼW���-����u���)���B���h������掼�=��+������ˆ�������i��Ϙ��'��Ar��M���<ٝ�t����
��������+���=���\��Z����ȧ�"���s��Jګ�G�������!��,���X鲼UA������5׶����dJ��nx��Ӡ��wƼ��  �  �@O=*�N=:N=BzM=k�L=�&L='rK=I�J=��I=>I=R�H=�G=�G=oiF=n�E="E=��D=��C==dC=�B=MB=8�A=2A=l�@=�@=�^?=ɳ>=�>=�L==d�<=�;=�%;=zs:=`�9=V9=�~8=��7=tP7=��6=�76=��5=A(5=۞4=�4=O|3=[�2=]92=c�1=P�0=�0=�S/=4�.=��-=�-=A,=�~+=J�*=b�)=�:)=�v(=Ԯ'=��&=�&=� %=4*$=�#= "=�� =�z=K=��==+n=��=D=;A=�r=!�=��=��=��
=�	=�!=�-=q3=1=�J�<��<V��<��<�+�<��<|F�<���<�S�<���<�p�<'�<��<�c�<$!�<(�<���<疴<�s�<xO�<%�<w�<���<o_�<�<���<�&�<l��<�8�<IĀ<��x<q�o<�#g<�^<3�U<��M<�(E<�<<q�4<[m,<2$<��<��<<�y<Ő�;9 �;=Q�;t��;�Ԭ;R&�;���;Np;��M;��+;�
;A��:l�:��:�q�8Qƹ�;c��ӱ��^���"K:�U[�r�{�����#��㭻�A���,̻�ڻ`n�4���k)�5+���jI��q�!`�J!�ٸ%�N4*�^�.���2��7�G';��?�n�B��~F���I��"M�u)P�>�R���U�8$X�q|Z���\�#�^���`��c��0e�<gg�t�i��#l�o�n��Iq���s�-�v��^y�|�W�~�^����ǁ���1���#��{-���0���0���1���8��9J���i�����1ێ�,���������Z���ĕ��)��3���Lڙ�9"��&^��~���ﳞ�GП�6格J���&��)���N��؂��ǧ����0��~e��,ޮ�oU���Ʊ�:/������޵��"���[���������ʻ��弼�  �  �2O=b�N=�N=�vM=!�L=�)L=�xK='�J=WJ=SSI=�H=��G=G:G=^�F=�E=�GE=��D=@D=�}C=�B=�[B=�A=�7A=��@=� @=�Z?=��>=��==�===�<=��;=F;=}Q:=Ԡ9=��8=�V8=ѽ7=�,7=D�6=�6=�5=w5=v�4=U4=w3=�2=:2=C�1=�0= "0=>e/=�.=��-=�%-=Me,=��+=V�*=� *=�[)=�(=��'=��&=�&=�'%=�,$=#=��!=�� =�o=d=?�=e�=;P=��=��=v=�F=�p=��=��=J�
=i�=.	=K=]$=�%=M;�<��<���<��<�9�<j��<jj�<V��<|��<?#�<Q��<�Z�<� �<Z��<�d�<�$�<�<C��<,��<�a�<�/�<f��<{��<DV�<]�<��<��<��< �<��<x<�9o<{f<��]<&XU<c�L<�D<�v<<aO4<U+,<� $<%�<�t<�<��<��;�U�;���;aC�;��;�2�;eÊ;��r;$nP;�H.;�r;���:���:�$:S9s9����`������X��L�:���[��y|�����֞�&��� C���Kͻ�ۻK�黤���n�����E������׍�">!���%�h:*���.���2���6�K�:���>���B��F��dI�яL��O��dR��U�ȝW�kZ��W\�)�^�o�`���b�$e��bg�2�i�f7l�/�n��yq��8t�� w�p�y�w�|��,�Iހ����eA���[��fh���i���b���X��RP���N��Y��ar�������׎��!��Jw��?Ԓ�4������햼�B������ ՚�����F���s��ڙ�������ء�W���<��mH��ł���̧��'������	���������.������/x���ڴ�,.���q��O���$˹��庼d���D
���  �  7#O=�N=�N=vpM=Y�L=�(L=�{K=}�J=�J=�dI=�H=rH=�YG=v�F=�F=CiE=��D=-D=x�C=q�B=�fB=]�A=�9A='�@=p�?=�S?=Ӣ>=��==_-==Cl<=��;=��:=)0:=z|9=x�8= 08=v�7=�	7=�6=�6=r�5=!5=��4=�3=�n3=X�2=572=��1=]�0=�*0=s/=_�.=s�-=�B-=��,=��+=�+=A*=�x)=��(=��'=��&=�&=5+%=-,$=�#=~�!=N� =3b=��=]r=�=H2={=��=Y�==[F=�m=��=B�
=��=�=|=T= =�%�<�<��<Ñ�<AA�<"��<m��<�$�<.��<4`�<���<5��<qG�<!��<נ�<oW�<��<ڴ<��<�l�<�2�<��<��<�F�<Pۖ<b�<�ݍ<S�<�Ƅ<�>�<�w<՛n<��e<K9]<O�T<�gL<�.D<%<<�3<��+<Y�#<�<�S<��
<�y<l��;���;�7�;e׿;�w�;��;(Ӌ;�)u;��R;�0;K�;h��:Kۖ:� ):#{9���_L_��ǰ��#�E��u�:�U&\��Z}�:5��������@���bλ��ܻ������:������S��J��3���g!���%�N*�+�.�;�2�O�6���:��>��5B��E���H��L��O��Q�ގT��&W� �Y�?\��W^�q�`�{�b�ge�zlg�|�i��Wl���n�߱q�D�t��Xw�Q1z���|�>���(���d�����-���ϫ��D�������悈�:r���i���m��=������#ێ�`���k��.�������h��K���u���L��A���b͛����5;���j�����ྡ��碼`�� I������l٧��9��ѩ���'��0����:��Ű�%H�����j&��[{��e����츼.�����a)���1���  �  dO=�N=�M=4hM=x�L=�%L=�{K=��J=G J=lrI=(�H=H=tG=��F=�(F=A�E=�D=�BD=��C=�C=�nB=��A=09A=[�@=�?=�J?=��>=Q�==�==�X<=V�;=;�:=G:='\9=��8=8=\w7=��6=�f6=��5=4n5=?�4=u4=��3=�d3=��2=22=��1=��0=y00=P}/=[�.=.=cZ-=q�,=W�+="+=�[*=v�)=>�(=��'=�'= &=�+%=)$=�#=��!=ϫ =!T=��=C^=l�=�=%\=|�=	�=|�=� =�I=�p=��
=ʹ=��=q�=R=�	=x�<���<S��<��<|C�<���<$��<E�<���<]��<'8�<P��<G��<v(�<���<)��<�4�<��<ȯ�<Bq�<j0�<��<n��<4�<;Ö<�C�<���<�&�<˒�<s�<��v<^n<OIe<o�\<�7T<p�K<5�C<��;<��3<&�+<��#<�g<-<��
<_j<���;-��;���;�I�;��;J�;���;?w;�T;��2;�g;���:�p�:�-:˘!9;ɶ�Y�^��ް�Z��!N�;���\�GB~�ď�u:��Fe���$���[ϻ[�ݻ��������Ɗ�6��C��:������!�q&��i*�&�.���2���6���:��l>���A��WE��H�~�K�p�N�YeQ�!T���V��QY�]�[��+^���`���b�5"e�cg�>�i��}l�L'o��q�K�t�H�w�ǒz��m}����aj�������у�>愼4腼Yۆ��ć����ޓ��o���B���S���w���^㎼R ��f��ذ������;G��Ď��Fӗ�<��qU��l����ќ�	��;E��z��g���Xޢ�%���N��㔦�n駼/N��Kê��F��Wԭ��f�����Ձ��D���:i������ ���,���F���R��0V���W���  �  �O=��N=T�M=7`M=a�L=�!L=�zK=}�J=�%J=�{I=_�H=�,H=y�G=��F=�>F=&�E=��D=�RD=�C=KC='sB=��A=E7A=�@=��?=TB?=��>=f�==�==PH<=x�;=غ:=��9=�B9=�8=@�7=B]7=?�6=iP6=��5=�\5=I�4=;h4=��3=�[3=u�2=�,2=k�1=l�0=k30=�/=��.=g .=�k-=e�,=��+=P7+=�o*=	�)=��(='�'='=�"&=+%=@%$==#=�!=V� =�G=+�=�M=-�=� =�C=�{=��=#�=�=H-=]V=o~
=�=��=��=��=u� =^��<���<���<���<�B�<1��<���<�[�<�
�<���<+b�<{	�<D��<�Q�<���<���<�J�<.��<���<�q�<M+�<�ޣ<���<F"�<���<�)�<ř�<�<�h�<2�<��v<��m<��d<<\<��S<�K<8dC<�Y;<q\3<_+<]W#<Y<<4	<��
<�X<1��;���;=��;��;���;�q�;�\�;��x;DV;=�3;@�;N2�:*O�:�/: �(9;�����^��%��["�r��T<�ρ]�5��;��Ƞ��������� лp�޻M��-���~�����Z�6��t��-��!�%0&�"�*��.�k�2�k�6�s�:��P>�y�A�!E��FH�WNK�":N��Q�R�S��|V�Y��[�G^��s`�j�b�Z-e��g��j�{�l��Qo�ur�u���w���z�l�}��I��N���ނ�����������>뇼̈�V�������ݘ�����������쎼�$���d��t����쓼Y/���o������똼F*���i������라�)���f�������٢����U����������Ja���٪�.a��@�֊��:!������K0��֝��A���J5���^���t��H|���z��w���  �  ��N=�xN=��M=yZM=οL=�L=yK=�J=�(J=)�I=B�H=�6H=`�G=��F=�KF=��E=E=a\D=k�C=+C=�uB=��A=s5A=n�@=��?=]<?=��>=>�==n==l=<=t;=��:=X�9=N29= �8=%�7=�L7=}�6=�A6=��5=>Q5=7�4=�_4=q�3=&U3=�2=�(2=͆1=��0=�40=��/=�.=�(.=�v-=��,=�,=lD+=7|*=ɬ)=3�(=V�'=�'=�#&=�)%=4"$=�	#=��!=� =^?=y�=rB=~�=��=�3=pj=[�=v�=�=C=lE=�n
=�=#�=��=^�=� =
��<���<���<�< A�<z��<��<�i�<R�<r��<�{�<�$�<U��<�j�<��<R��<�W�<��<¹�<�p�<�&�<�֣<}�<y�<O��<��<Ȅ�<��<6M�<�j<�Rv<m\m<�d<��[<s�S<lGK<E*C<&;<�.3<?7+<�4#<�<]�<�
<�K<���;���;���;���;�ʯ;ʞ;9č;�hy;~.W;��4;�; ��:�k�:0u1:R�,9�4��آ^��k��4�����h<�{�]�G�������%���r���P���л�D߻�+�|J��P��	�a���� ��[O���!��H&���*���.���2���6�>�:��@>�̲A���D�%H��K��N�|�P�1�S��PV�I�X���[��]�sm`���b��6e�ѣg��"j�ĺl��oo��@r��(u�;x�{���}��h�����G ��!)��p:���6���"��A��7∼�É�H���)��������ʍ�
��(���d��*����㓼3!���\��]���\Ҙ�����O��n���S֝����[��G���0آ�t���[��y���?���n��k骼3s���������;��]Ͳ�GP��w�����
W����钺�W���В������  �  �N=�uN=�M=kXM=&�L=�L=xxK=+�J=�)J=�I=��H=Q:H=w�G=Y�F=RPF=G�E=zE=�_D=˺C=�C=IvB=��A=�4A= �@=��?=::?= �>=M�==#==�9<=�o;=.�:=�9=�,9==~8=3�7=�F7=�6=�<6={�5=DM5=��4=j\4=��3=�R3=�2='2=Ņ1=+�0=50=̈/=�.=�+.=Cz-=��,=
,=�H+=a�*={�)=�(=Q�'=�'=$&=j)%=!$=�#=��!=� =P<=�=�>=*�=��=X.=�d=.�=�=��=0=�?=�i
=w�=	�=G�=+�=Q� =a��<���<ί�<N}�<�@�<���<��<Pn�<�#�<w��<Ä�<�-�<\��<Is�<%�<ش�<�[�<�<#��<}o�<8$�<�ӣ<�x�<m�<^��<�<)}�<@�<�C�<]U<Q;v<�Cm<"xd<}�[<1qS<�1K<�C<�;<�3<*+<@)#<�<a�<�
<hG<t��;|��;��;c��;��;��;H�;��y;�|W;�,5;��;��:]Ĝ:|�1:h�-9���$�^� ������$�d�<��$^�z�������G������{��&�л	t߻s[�ux���e�|.	���������n[���!��Q&��*�U�.���2�*�6���:�<>���A�s�D�1H��K��M���P�.�S�UAV�u�X�1y[���]��k`���b��:e���g�]*j���l�izo��Lr��6u��-x��&{��~��s���ʁ�$���4���E��oA��q,������鈼=ʉ�?���i�������΍�����z*��7e��ꢒ���������V�������ɘ�����F��'���=ϝ�b��uW��W����ע����^������H��ys��謁�y��=������"E���ײ�P[�� ˵�d#���b��;���>����������o����  �  ��N=�xN=��M=yZM=οL=�L=yK=�J=�(J=)�I=B�H=�6H=`�G=��F=�KF=��E=E=a\D=k�C=+C=�uB=��A=s5A=n�@=��?=]<?=��>=>�==n==l=<=t;=��:=X�9=N29= �8=%�7=�L7=}�6=�A6=��5=>Q5=7�4=�_4=q�3=%U3=�2=�(2=͆1=��0=�40=��/=�.=�(.=�v-=��,=�,=kD+=6|*=ɬ)=3�(=V�'=�'=�#&=�)%=7"$=�	#=��!=� =j?=��=�B=��=��=�3=�j=��=��=^�=�=�E=\o
=��=��=}�=�=�� =^��<!��<���<R��<AB�<���<��<cj�<��<���<1|�<�$�<3��<pj�<S�<���<�V�<	�<���<ro�<P%�<�գ<�{�<A�<$��<��<̃�<��<L�<�i<�Qv<	\m<�d<Y�[<,�S<�HK<�+C<�';<�03<o9+<>7#<;!<��<��
<	N<���;Q��;���;E��;Jͯ;.̞;�ō;*jy;?.W;��4;��;���:j_�:�W1:�!,9󀴹�^�����®�A� t<��^�&�������*��w���T����л<H߻�.��L��Q�t	�&���������O�?�!�I&�Й*���.���2���6�U�:� A>�ڲA��D�.H��K��N���P�4�S��PV�K�X���[��]�tm`���b��6e�ѣg��"j�ĺl��oo��@r��(u�;x�{���}��h�����G ��!)��p:���6���"��A��7∼�É�H���)��������ʍ�
��(���d��*����㓼3!���\��]���]Ҙ�����O��n���S֝����[��G���0آ�t���[��y���?���n��k骼3s���������;��]Ͳ�GP��w�����
W����钺�W���В������  �  �O=��N=T�M=7`M=a�L=�!L=�zK=}�J=�%J=�{I=_�H=�,H=y�G=��F=�>F=&�E=��D=�RD=�C=KC='sB=��A=E7A=�@=��?=TB?=��>=f�==�==PH<=x�;=غ:=��9=�B9=�8=@�7=B]7=>�6=iP6=��5=�\5=I�4=;h4=��3=�[3=u�2=�,2=k�1=k�0=j30=�/=��.=f .=�k-=e�,=��+=O7+=�o*=	�)=��(='�'='=�"&=+%=F%$=E#=�!=h� =�G=K�=�M=c�=6=�C=�{= �=��=R=.=<W=f
=!�=��=�=,�=�� =���<N��<,��<���<�D�<+��<f��<a]�<��<a��<�b�<�	�<��<�P�<���<q��<GI�<^��<���<�o�<�(�<cܣ< ��<��<M��<�'�<ߗ�<c �<Og�<�<��v<ڡm<��d<�<\<�S<-�K<�fC<1];<@`3<Xc+<�[#<!A<<��
<�]<K��;��;Ҷ�;���;��;v�;]_�;2�x;�CV;��3;ܵ;��:e7�:��/:�'9K���S�^��O���M���p<���]�5 ��E��rѠ��������(л��޻����������G\�s��"u��.���!��0&���*�t�.���2���6���:��P>���A�7E��FH�dNK�,:N��Q�X�S��|V�Y��[�I^� t`�l�b�[-e��g��j�{�l��Qo�ur�u���w���z�l�}��I��N���ނ�����������>뇼̈�V�������ݘ�����������쎼�$���d��t����쓼Y/���o������똼F*���i������라�)���f�������٢����U����������Ja���٪�.a��@�֊��:!������K0��֝��A���J5���^���t��H|���z��w���  �  dO=�N=�M=4hM=x�L=�%L=�{K=��J=G J=lrI=(�H=H=tG=��F=�(F=A�E=�D=�BD=��C=�C=�nB=��A=09A=[�@=�?=�J?=��>=Q�==�==�X<=V�;=;�:=G:='\9=��8=8=\w7=��6=�f6=��5=4n5=?�4=u4=��3=�d3=��2=22=��1=��0=y00=O}/=[�.=.=bZ-=p�,=V�+="+=�[*=u�)=>�(=��'=�'= &=�+%= )$=�#=��!=� =DT=��=�^=��=S=�\=�=��=O�=�!=�J=/r=�
=G�==�="�==�=�<]��<���<7��<�F�<���<���<G�<���<���<�8�<s��<��<�'�<z��<^~�<�2�<g�<鬰<%n�<"-�<,�<
��<�0�<��<�@�<��<3$�<ؐ�<��<��v<Kn<BIe<h�\<�9T<`�K<�C<F�;<�3<"�+<#�#<�n<�3<��
< q<���;��;C��;AS�;v�;�;u��;�w;\�T;��2;�^;���:'O�:��,:�" 9E����_�~�����rm��;�~�\��_~�>ҏ��G���q��!0���eϻY�ݻ���������F��Q��E�<������!�9&�1j*���.���2���6��:��l>���A��WE�)�H���K��N�deQ�$!T���V��QY�a�[��+^���`���b�6"e�dg�?�i��}l�M'o��q�K�t�H�w�ǒz��m}����aj�������у�>愼5腼Zۆ��ć����ޓ��o���B���S���w���^㎼R ��f��ذ������;G��Ď��Fӗ�<��qU��l����ќ�	��;E��z��g���Xޢ�%���N��㔦�n駼/N��Kê��F��Wԭ��f�����Ձ��D���:i������ ���,���F���R��0V���W���  �  7#O=�N=�N=vpM=Y�L=�(L=�{K=}�J=�J=�dI=�H=rH=�YG=v�F=�F=CiE=��D=-D=x�C=q�B=�fB=]�A=�9A='�@=p�?=�S?=Ӣ>=��==_-==Cl<=��;=��:=)0:=z|9=x�8= 08=v�7=�	7=�6=�6=r�5=!5=��4=�3=�n3=X�2=572=��1=\�0=�*0=s/=^�.=r�-=�B-=��,=��+=�+=A*=�x)=��(=��'=��&=�&=;+%=7,$=�#=��!=m� =]b=��=�r=j�=�2=�{=@�=3�==�G=o=6�=�
=��=�=�=|=U=f*�<}�<L��<Օ�<
E�<���<l��<'�<&��<�a�<� �<`��<�F�<��<2��<<U�<��<�ִ<���<�h�<�.�<��<ߞ�<�B�<iז<t^�<`ڍ<-P�<�Ą<=�<a}w<��n<��e<{:]<��T<�kL<o3D<�<<��3<��+<>�#<7�<\<Z�
<8�<0��;X��;�D�;��;���;'�;�׋;.u;�R;�0;7�;p��:��:P�(:"�9���T�_�s��ho���;��K\�C}��F��-���Ȫ��QN��Doλ��ܻK��s���=�� �+��x��������h!���%��N*�ș.���2���6��:�X�>��5B��E���H��L�O�$�Q��T��&W�&�Y�D\��W^�t�`�}�b�ie�{lg�}�i��Wl���n��q�D�t��Xw�R1z���|�?���(���d�����-���ϫ��D�������悈�:r���i���m��=������#ێ�`���k��.�������h��K���u���L��A���b͛����5;���j�����ྡ��碼`�� I������l٧��9��ѩ���'��0����:��Ű�%H�����j&��[{��e����츼.�����a)���1���  �  �2O=b�N=�N=�vM=!�L=�)L=�xK='�J=WJ=SSI=�H=��G=G:G=^�F=�E=�GE=��D=@D=�}C=�B=�[B=�A=�7A=��@=� @=�Z?=��>=��==�===�<=��;=F;=}Q:=Ԡ9=��8=�V8=ѽ7=�,7=D�6=�6=�5=w5=u�4=T4=w3=�2=:2=B�1=�0="0==e/=�.=��-=�%-=Le,=��+=U�*=� *=�[)=�(=��'= �&=�&=�'%=�,$=*#=��!=�� =�o=�=��=��=�P=)�=��=j=�G=&r=	�=N�=&�
=p�=\=�=�&=K(=D@�<q�<���<���<�=�<;��<�m�<"��<���<�$�<2��<)[�<- �<,��<c�<7"�<�<���<?��<�]�<,+�<��<٧�<�Q�<�<t{�< �<L�<[��<�<>x<#8o<�zf<L�]<�ZU<f�L<N�D<1}<<�V4<�3,<z	$<a�<,~<�<��<���;f�;4��;P�;���;u:�;�Ȋ;��r;9mP;B.;�f;���:�r�:�#:�S9�U���ca�b���X� ���:�w�[�5�|�񴎻1螻�Ϯ�PR���YͻW�ۻ�����u��n���H�S�����v��s?!���%�C;*�n�.� �2�G�6���:��>��B�F��dI��L� �O��dR�U�ѝW�sZ��W\�.�^�r�`���b�&e��bg�4�i�g7l�/�n��yq��8t�� w�q�y�x�|��,�Iހ����eA���[��fh���i���b���X��RP���N��Y��ar�������׎��!��Jw��?Ԓ�4������햼�B������ ՚�����F���s��ڙ�������ء�W���<��mH��ł���̧��'������	���������.������/x���ڴ�,.���q��O���$˹��庼d���D
���  �  �@O=*�N=:N=BzM=k�L=�&L='rK=I�J=��I=>I=R�H=�G=�G=oiF=n�E="E=��D=��C==dC=�B=MB=8�A=2A=l�@=�@=�^?=ɳ>=�>=�L==d�<=�;=�%;=zs:=`�9=V9=�~8=��7=tP7=��6=�76=��5=A(5=۞4=�4=N|3=[�2=]92=b�1=O�0=�0=�S/=3�.=��-=�-=A,=�~+=H�*=a�)=�:)=�v(=Ԯ'=��&=�&=� %=@*$= #= "= � =�z=�=�=r=�n==�==7B=!t={�=��=a�=��
=	=�#= 0=�5=�3=P�<�$�<G��<ʒ�<�/�<���<�I�<���<�U�<P��<�q�<Z�<���<\b�<=�<��<߹�<E��<�o�<K�<b �<��<4��<�Z�<���<���<*#�<��<56�<(<ȧx<��o<�#g<m�^<��U< �M<�-E<��<<�4<�u,<-;$<8�<x�<�<`�<���; �;n`�;���;r߬;�.�;��;Sp;�M;í+;��	;Kl�:ȶ�:�r:�N�8�wǹ�c�!(����.��Ww:��2[�e�{�}-���6��Z���iQ��;̻��ڻ�y�����-��.����K��s��a�� !��%�15*��.�t�2��7��';�?���B��~F��I��"M��)P�N�R���U�A$X�x|Z���\�(�^���`��c��0e�=gg�u�i��#l�p�n��Iq���s�-�v��^y�|�W�~�^����ǁ���1���#��{-���0���0���1���8��9J���i�����1ێ�,���������Z���ĕ��)��3���Lڙ�9"��&^��~���ﳞ�GП�6格J���&��)���N��؂��ǧ����0��~e��,ޮ�oU���Ʊ�:/������޵��"���[���������ʻ��弼�  �  @KO=f�N=�N=�yM=��L=< L=+hK=N�J=��I=t&I=�eH=ƨG=��F=BF=d�E=�D=�cD=c�C=�HC=��B=�;B=-�A=�(A=��@=�?=�^?=+�>=�	>=JX==�<=)�;=LA;=̓:=h�9=�E9=E�8=�	8=�r7=��6=P6=��5=65=��4=�4=�}3=��2=52=Ԃ1=%�0=`0=�?/=v.=��-=r�,=_,=3W+=֕*=��)=F)=�X(=Օ'=$�&=>�%=�%=�#$==#= "=�� =��=!=��=m#=c�=_�=�,=nk=�=U�=t�=�=n=I-	={9=�@=�A=:;=PX�<u&�<\��<{��<N�<~��<� �<l��<;�<���<}#�<���<`�<��<��<��<��<Uh�<.N�<�1�<f�<X�<K��<�\�<�<q��<�@�<։<�j�<��<L9y<�yp< �g<�#_<��V<�N<�E<(F=<��4<[�,<l^$<<��<�<n<�X�;֢�;���;q۽;o�;��;H]�;��m;�K;�);Mu;q��:l��:��:)_�8�%й2g��`��Ԇ����t:���Z��S{�h�������)(��(]���'˻ |ٻ�O绫���ҩ �g��8����/@�2A�i!���%�
>*�y�.�y3�?B7��g;�l?��IC�P�F��uJ���M���P���S��@V��X�4�Z��]��._��4a�x<c��Pe�Qzg���i�
l�]�n��'q���s�Gbv���x�d�{��~��G���z��6���~ǃ��ᄼW���-����u���)���B���h������掼�=��+������ˆ�������i��Ϙ��'��Ar��M���<ٝ�t����
��������+���=���\��Z����ȧ�"���s��Jګ�G�������!��,���X鲼UA������5׶����dJ��nx��Ӡ��wƼ��  �  RRO=*�N=
N=�uM=P�L=�L=�[K=k�J=��I=7I=�HH=�G=��F=F=�sE=[�D=e@D=~�C=�,C=B�B=�(B=�A=!A=֎@=��?=z[?=�>=[>=g`==1�<=�<=Y;=V�:=�
:=�g9=�8=
+8=�7=��6=�d6=R�5=f@5=��4=t4=|3=�2={-2=x1=��0=L�/=b*/=q\.=͍-=��,=��+=,1+=�o*=�)=��(=;(=v|'=K�&=��%="
%=�$=##=U�!=�� =��=�(=X�=�5=,�=��=�N=q�=��=�==�'=�8=�D	=.K=M=fI=?=�X�<� �<���<jt�<�<���<���<�f�<4��<�R�<���<#l�<��<_��<���<k�<�O�<c;�<s)�</�</��<�Σ<֙�<�W�<
�<}��<W�<���<J��<�9�<+�y<�q<�Zh<��_<�W<{�N<jF<;�=<#05<��,<�r$<<�<��
<tL<���;�$�;
&�;��;T��; �;�+�;�!k;�{H;Rp&;�;�a�:�:��:�X�8��ٹk�<�Q����n���:�^�Z�&�z��c��b���w������'2ʻ�sػ�B�2���4 �>X�i4�b����_.��!���%�_T*�]�.�^.3�xz7��;�%�?��C��rG�z�J��ON��cQ�:T�,�V��:Y��r[�Ƈ]�u�_��{a�=tc��{e���g���i�
(l��n�dq��s��&v���x�`,{��}�w��5��-`������진��ą��܆���.��R!�� B���n����������T��|����7��e���B1����������r��a��������!���9��E��H���H���K��|W��p��P���-ѧ�����n��.ͫ�^0��*�������
S��&��������J��5���ַ�E��"K��6~�������  �  DVO=,�N=�N=�oM=��L=L=�NK=p�J=��I=��H=�.H=�jG=߭F=g�E=�QE=�D=� D=ӖC=�C=o�B="B=ƕA=�A=��@=�?= V?=s�>=/>=Ke==��<=�<=)l;=��:=.%:=q�9=�8=�F8=ة7=�7=ru6=��5=SG5=�4=P4=�w3=R�2=Z$2=m1=��0=d�/=</=�D.=�r-=��,=��+=�+=!N*=��)=��(=
 (=e'=��&=u�%=��$=X$=@#=��!=)� =5�=o-=M�=kC=
�=/=rj=E�==�=4=�.=@C=P=�V	=�X=�U=�M=�?=�S�<��<]��<�_�<V��<Z_�<��<=6�<H��<y�<ڔ�<�&�<G��<���<aT�<3�<`�<�<w�<���<;ާ<���<<�N�<��<���<�f�<��<t��<�g�<�&z<~q<k�h<�-`<"�W<�N<�YF<>�=<�Z5<��,<�z$<�<�~<��
<�$<���;��;��;wW�;�#�;6�;��;��h;?/F;J,$;j�;�c�:�,�:��	:��=8q���o�����y
��s����:���Z�2�z��%�������꫻sպ�kfɻ��׻oc���+���i���������&��!�)�%��q*�2�.�K^3���7���;��@�@D���G��xK�0�N�A�Q���T��XW�}�Y�y�[���]�6�_�-�a���c��e�ÿg���i�{:l�:�n��
q�_�s�W�u��mx�3�z��>}���s����&���P��}x��v���:����އ�n�������F��y��Ĺ���
��"m���ޑ��[��Cߔ�(c��&ᗼPS��>������=��b�� u���y��v���o��Sl��rr�����������ݧ�� ���o��:ƫ�~ ���z���ү�'���w���ų����Z�����m渼'���c�������  �  �WO=��N=�N=�iM=ֹL=KL=�BK=�|J=��I=.�H=�H=[SG=��F=��E=�6E=ęD= D=�C=2�B=��B=�B=��A=\A=0{@=h�?=AP?=�>=d>=�g==��<=�<=�y;=��:=�8:=ƙ9=��8=b[8=H�7=7=-�6=��5=TK5=��4=�4=�r3=��2=�2=�b1=v�0=�/=�/=�1.=]-=��,=�+=�*=�3*=!x)=��(=u
(=�Q'=3�&=��%=N�$=�$=�#=G�!=�� =/�=u/=��=�L=��=�(=	=F�=a�=D(=GE=dW=�`=�c	=�a=�Z=�O=�>=�L�<C�<	��<�L�<���<C�<a��<��<�t�<���<`�<��<ڕ�<R�<6#�<X�<���<Y�<K�<ܫ<ȧ<���<�|�<�D�<��<ۻ�<sp�<�#�<�օ<a��<nvz<��q<?1i<�`<��W<�4O<m�F<I�=<<v5<��,<dz$<T�<�i<H�
<��<�8�;\7�;H�;���;Bt�;SC�;AE�;�g;�aD;�d";�';�:�:�N�:e:��7B��ar����y@��i��G;��[���z�Q����e�����RS����Ȼ��ֻV���!���@��%�����%���&�^ !�X�%���*��/�\�3���7�..<�\Y@�``D��8H���K��:O�VWR��-U���W��Z��9\�Q7^�J`���a��c�u�e�Z�g�"j��Nl��n�
q��ss���u��@x�/�z�J�|�HK�bЀ�����(���U�����t����ч��������#M��$����ȍ�v�����w����y��b��y���P��Ʉ���隼.9��r���F���~����������������� ���/����ꧼp)��9s���ë����~i����������Q�������崼z0���{��~Ÿ����Q��;����  �  dXO=7�N=sN=eM=	�L=o�K=�:K=�sJ=R�I=�H=FH=SDG=p�F=�E=�%E=��D=�C=CqC=��B=�vB=��A=�A=��@=�t@=��?=�K?=�>=L>=�h==�<=�"<=E�;=F�:=E:=�9=�9=h8=��7=]'7=�6=4�5=WM5=~�4=�4=Lo3=|�2=�2=�[1=%�0=v�/=��.=%.=	O-=b{,=��+=1�*=�"*=�g)=H�(=|�'=�E'=R�&=J�%=_�$= $=#=��!=�� =�=0=��=SR=��=3=��=Y�=A=7='S=�c=�j=fk	=�f=u]=�O===�F�<S�<���<�>�<w��<�/�<ܔ�<��<�W�<1��<8>�<>��<s�<o0�<��<��<�ܷ<j׳<>ӯ<�ʫ<��<Û�<Cr�<z=�<���<X��<�u�<5.�<c�<���<��z<r<ji<o�`<�X<�`O<l�F<a><(�5<��,<[w$<��<dY<��
<��<C��;E��;���;�Y�;��;>Ė;׻�;��e;�;C;�B!;" ;74�:Q�~:c/:�7���J�t�2��>����O�;�]8[�[�z��錻|;���E�����pȻՌֻ�T�u������e�����pp�T���(��)!�H�%�D�*�1/��3�*	8��U<���@�I�D��qH��L�}O�ڛR�wrU�QX�lUZ�*s\�qj^��J`�#b�d���e�q�g�� j�L^l�!�n��q�ms�K�u�#&x�zz���|�&�ȵ���ၼ!�� @���o��,���]ʇ�V����!���R�������Ӎ�~*��F���
��3����������v+��j����
��f[�����~�����������_���ޚ��=�������Ʀ����70���v��+ë����u_������V󰼐:��쁳�#˴�����c��v�������G�������  �  !lO=f�N=�&N=D}M=\�L=�L=�FK=/uJ=ЛI=
�H=��G=�G=�DF=މE=��D=�GD=�C=�FC=o�B=�mB=�B=3�A=�!A=M�@=�@=N�?=&�>=�F>=D�==X==�h<=+�;=8;=D�:=	:=)n9=�8=�/8=Ȏ7=�6=R6=��5=�5=.�4=��3=uG3=ə2=��1=�1=�H0=�n/=(�.=��-=��,=g
,=\E+=��*=.�)=E;)=��(=��'=�Y'=P�&=��%=�%=�$=�#=��!=� =b=�=��= =i=��=�="8=�W=f=�f=7]=>M
=�9=$=/=��=9��<�F�<a��<�O�<6��<���<�/�<2b�<���<���<Q7�<G��<H�<��<Qܿ<�ϻ<�շ<�<���<��<<��<Gߣ<���<��<$>�<5��<��<�h�<�#�<%߁<�-{<�r<��i<6a<�JX<htO<�F<�=<R15<=�,<�$<t<e�<�
<W0<�6�;��;J��;���;=��;��;�;��Z;	H7;��;X��:��:\P:Ǎ�9�1�ol!����P8ͺPR��^&���F��f��h��n/��ج��ڱ�����`FϻK�ݻ����B��^J�׷	�T�� ���?�$y ��n%��-*�W�.��H3�&�7�7(<��@�#�D���H���L�$�P�FT��%W�p�Y�&6\��@^��
`�S�a�}'c�Ǧd��6f�/�g�,�i�|�k���m��p�Wfr�²t���v��1y��a{�ۍ}�Ͻ�m����!���N��k���ӳ���䆼���:���`��A���l���V���^��ѐ��Y��T�������mD���䘼s���盼�<���o�������v��:V���(��)����Σ�`���t���俦��秼�!��ah��N�������:G��򈯼8ư����pA��$���#ҵ�$���x���̹����yf���  �  �lO=�N=�(N=7�M=��L=�L=:KK=�yJ=�I=��H=>�G=�G=�LF=��E=!�D=�OD=��C=�MC=��B=�sB=�	B=͛A=�%A=�@=@=�?=i�>=6H>=��==�==vf<=��;=u3;=қ:=0:=h9=Q�8=�*8=Պ7=Y�6=�P6=ͷ5=� 5=$�4=��3=�J3=`�2=��1=1=fM0=jt/=@�.=V�-=�,=J,=rM+=��*=�)=�B)=K�(=(=�^'=�&=��%=�%=�"$=�#=��!=�� =�b=Y�=��=��=�d= �=j�=,1=�P=�_=�`=�X=�I
=�7=#=i=��=���<K�<���<uV�<ʵ�<d��<�9�<%n�<��<���<jG�<��<�X�<��<��<o޻<�<(�<���<D�<���<��<q��<��<�B�<���<�<�e�<�<�ց<}{<�wr<��i<�a<93X<Q`O<t�F<��=<�+5<X�,<
$<Rz<�<�!
<*=<�T�;E��; �;�"�;<+�;�S�;l�;�/[;T�7;>�;ޕ�:M�: �Q:���9���l����9�̺�� &�iF�6�f��^���/��;����ﱻ~���umϻ��ݻS�뻆m��]�Y�	�	��Ǽ�S?�9t �#f%��"*��.��93���7�	<�s@���D� �H�2�L�e�P�^�S��W���Y�\� #^���_�p�a�Mc�͒d��$f��g���i���k�N�m�dp��ar���t��v�#<y�	q{���}�x��p���-���Y��ȉ��庅��醼����9��0^��݆��칌�����LW���Ȑ��P��듼�����7���֘��c���כ�#,��i_��r��Qh���H�������ţ���������⸦��᧼����d������� ���J��򎯼�ΰ����M��K����ݵ��.������9ӹ�d ���g���  �  nO=:�N=a/N=a�M=M�L=HL=WK='�J=�I=��H=9�G=�*G=HcF=��E= E=.gD=��C=DbC=f�B=��B=TB=��A=�1A=i�@=T$@=�?=f�>=�K>=6�==�==�_<=n�;=�%;=��:=]�9=�U9=,�8=�8=�~7=�6=$L6=�5=#5=�4=��3==S3=4�2=��1=d*1=$[0=��/=��.=��-=��,=7),=e+=C�*=�)=X)=׶(=c(=6n'=t�&=��%=�%=�+$=f#=��!=u� =�c=1�=�~=��=�V=&�=$�=�=.<=jL=YP=4K=@
=�1=� =/=�=[��<
Y�<���<�i�<G��<��<2X�<+��<���<~�<�v�<���<���<3B�<V�<h�<�<y�<��<[!�<��<���<�џ<���<�M�<Y��<���<X[�<��<���<��z<g.r<�xi<2�`<��W<�%O<7fF<D�=<*5<#�,<�$<x�<��<qB
<\c<v��;R>�;Y��;���;�ƥ;��;g��;4�\;n9;�;���:ߪ:�1W:�m�9�����!2���˺�R��%���E�MXf�L��h9���ᢻ8���9��u�ϻ�A޻�G�j�����]�	���_���@�i �RP%�*��.�	3�|7���;��:@��|D�!�H�ƉL��7P���S�5�V��YY��[���]���_�Ea��b��Zd���e���g���i�s�k�O�m�b�o�lWr���t�Dw��[y�)�{�&�}�&���,��Q���z��ץ��aЅ�����7��19���W��^{�������덼�B�����T7��[Γ�p�� ��󭘼�7������L����/���D��>��g"��s���)Ϣ�/�������5��������Ч�����[��������\U��1����簼,���o������� ��;N������G湼�+���k���  �  �nO=%�N=�7N=Q�M=J�L=2,L=#hK=��J=F�I=T�H=3H=AKG=]�F=��E=o%E=��D=� D=�C=�C=ÜB=�-B=��A=BA=�@=�0@=]�?=�>=�O>=��==��<=1T<=��;=+;=�p:=|�9=�89=e�8=/8=k7=��6=�C6=�5=6%5==�4=��3=�^3=δ2=o�1=<1=Lo0=%�/=N�.=��-=�-=�L,=�+=1�*=�!*=6y)=��(=�/(=�'=�&=e&=�,%=28$=�)#=k "=ؽ =�c=c�=Ht=P�=j@=��=�=��=Y=�-=Q5=25=�/
=T'=�=$=��=/��<�k�<��<���<��<a@�<;��<���<=�<�[�<���<�<�<���<���<]�<�E�<@�<�C�<6I�<3H�<m:�<�<{�<穛<�Z�<=�<���<)H�<�<p��<nz<u�q<
�h<�<`<f}W<m�N<�F<�=<��4<̉,<)$<��<A<lo
<�<�-�;���;�:�;Oz�;Ե�;��;槁;�3_;m�;;��;�_�:-E�:�-_:N��9m�Ҹ�{�;����ȺT���$�?E���e�{<���V���.�����W���(�л�߻Y(��������>
�A=�����H��] ��4%��)��d.�8�2�?7�Ӛ;�Y�?�$D�+0H�$L�]�O��S��V�B�X��([��D]��$_���`�(sb�xd���e�ig�Mi��Zk���m�.�o��Lr���t�l,w�-�y�5�{�j<~�'C��g������t���Ԅ���W��C'��S;���P���l��N����ҍ�G&��b���F������B?��mۖ�jo��.�`�������坼���������砼�ơ����炣�*q���r��B�������B���GQ��V������h��I�������^������`��9��с���Ƹ�����@���t���  �  �lO=U�N=?N=�M=��L=$<L=�zK=��J=j�I=4I=�=H=�sG=��F=D�E=�TE=�D=,D=V�C=K/C=��B=GB=��A=$TA=>�@=�=@=R�?=��>=�Q>=G�==��<=�B<=v�;=-�:=M:=��9=H9=�w8=��7=�O7=@�6=o66=ͭ5=�$5=�4=\4=cj3=��2=22=�O1=��0=��/=��.=.=XB-=�y,=�+= +=�N*=�)=��(=�O(=/�'=��&=&=�;%=�D$=73#=�"=2� =La=m�=(d=��=q!=hi=U�=��=k�=W=�=�=�
=�="=)
=��=K��<}�<��<ޢ�<��<lm�<N��<��<�W�<���<��<G��<6�<O��<��<+��<�<�~�<�{�<�s�<`�<<�<��<켛<�d�<J�<��<}*�<ɾ�<�U�<n�y<Eq<�Th<e�_<��V<�AN<��E<�6=<��4<Xt,<�$<ȷ<�;<��
<��<��;Y��;4�;�v�;"ާ;Jb�;�;Pb;u ?;t�;�Z�:�Ŵ:�i:i
�9�ܖ�^��1Ԇ�FJƺhD���#�0�D���e��?������6���pg��<�»��ѻ�G�tW���tt�2�
����V��]�nZ �v%�x�)�\3.���2�"�6�WI;���?���C���G�syK��O��RR�RU�.X��qZ��\���^�T`� b��c��Ye�h$g�i�B+k�lm���o�KKr�
�t�D^w���y�dW|�ٿ~�n��������ق����O��'���4��=���C��lM���`�����鹍�-���m��l葼�r�����(����!��ۜ������R���������ê�����Ň���l���U��K��tR���o��������I��8������y����쯼�K����������O@��Ȇ���Ƿ�����4���_�������  �  �eO=c�N=�BN=E�M=�L=�IL=ӋK=��J=��I=�.I=�dH=g�G=,�F=�1F=j�E=$�D=�\D=��C=�TC=��B=b`B=�A=AdA=�@=nG@=�?=] ?=�O>=�==r�<=�+<=_x;=�:=y!:=�~9=��8=~J8=�7='-7={�6=�#6=��5=H 5=��4=O4=�r3=S�2=�2=b1=v�0=	�/=!/=�9.=�p-=5�,=��+=�4+=0�*=+�)=�")=4r(=�'=��&=#,&=�H%=5N$=V9#=I	"=6� =�Y=�=N=C�=	�=;<=	q=��=��=��=*�=A�=$�	=�=�=F=�=���<n��<�-�<h��<73�<��<x��<�O�<���<��<.��<
�<���<3P�<]�<��<≠<��<���<|��<K��<�V�<��<ɛ<g�<<��<j~�<a�<���<\�<�/y<�Up<G�g<]�^<�-V<��M<�,E<��<<L�4<�J,<�	$<�<.N<9�
<�<�9�;4(�;o��;.��;�!�;7ږ;���;��e;f�B;oH ;��:޺:��s:Mg�9-2���	��'���ĺ�\�m#�L/D��{e��e���򓻌H��:L���ûVӻ��Ứ��`E����$,�u��2a�����h �8%���)�5.�pk2���6�h�:�_*?��9C�. G�M�J��MN�u�Q��|T�j0W���Y���[��]�J�_�E�a�qJc��e���f���h�Ok�bVm�_�o�N[r���t���w�oHz���|�4`�j瀼����7��PQ���`���f���d��>]��^U���R��\���v�����BN������A���ǔ��M���˗��<��(����盼����@��)P��	P��FE��N6��*��4(���6��sZ��]���{樼�J��K���E5��u����%�����������P�������㶼���/K��?o������*����  �  �YO=��N=�@N=��M=�M=RL=U�K=��J=�J=�MI=�H=��G=�G= hF=��E=�#E=O�D=� D=qyC=�B=�vB={�A=�oA=��@=�K@=٩?={�>=H>=o�==��<=E<=%T;=��:=`�9=;J9=��8=�8=Ȋ7=�7=��6=�6=ܑ5=5=��4=�
4=wu3=H�2=L'2=�o1=�0=�/=V'/=Ab.=v�-=	�,=$,=bk+=&�*=@ *=!K)=K�(=��'=g'=�8&=�P%=)R$=�9#=�"=[� =HL=��=<2=I�=!�=8	=�8=�_=�=�=�=*�=��	=��=��=��=��=��<J��<F4�<k��<�L�<^��<�+�<���<� �<�s�<���<�z�<	�<��<&s�<|;�<��<��<qذ<ü�<㘨<�f�<h"�<�ɛ<$^�<�<�Z�<f͉<�?�<e��<ajx<�}o< �f<z�]<8_U<`�L<��D<�V<<�,4<Y
,<��#<J�<�I<��
<�<-��;	��;5��;��;qb�;�W�;pq�;�ti;�tF;��#;��;�
�:*f~:A�9ɲ��������rº���"��D��e�۶��'����EY��1Ż2�Ի�D�#a�l���P������j�W��N���� �!&%��)��-��O2�ґ6�&�:�_�>���B���F��/J�B�M�{�P��S�ESV�j�X�k[�~?]�=_�!a���b���d�ǿf��h���j�SWm���o�r�r�W=u��x���z��x}�D��jL���~��8���z���?������Y���b���6r��|c���b���u��]�������Y8��N��������������u���ژ�f1��Fy��t���1ڝ�d���������������+��.%���O��>����騼�V��fӫ��Y��*㮼�h���屼{V��2���
��pK���|�����Q������VǼ��  �  DHO=��N=�8N=8�M=} M=1TL=�K=(�J=b&J=�hI=�H=��G=9GG=2�F=��E=KWE=w�D=V)D=��C=vC=��B=� B=vuA=��@=dI@=b�?=l�>=�:>=�y==��<=�;=�,;=bp:=ݼ9=�9=bu8=a�7=�Y7=��6=c6=`�5=~|5=�5=ω4=�4=�q3=��2=�*2=x1=��0=�0=�D/=~�.=��-=�-=eX,=��+=��*=�,*=�p)=Ұ(=8�'=^'=S@&=�R%=�O$=�3#=)�!=w� =9=�=O=�`=�=��=r�=�"=HC=�`=}=��=�	=�=�=�=�=���<ix�<5.�<���<�[�<���<Y�<���<!O�<���<,X�<8��<�~�<� �<J��<���<�O�<~!�<Q��<�Ѭ<루<�i�<1�<$��<mI�<�<�-�<���<��<w[�<��w<��n<Y�e<�]<��T<�&L<f�C<��;<]�3<J�+<Ţ#<x<*,<�
<<���;��;�C�;kd�;��;��;��;��l;�J;y';n>;Z��:��:�V:,q�6Ƀ��������~����"��fD�vOf�0���.��	 ��s�����ƻ�ֻ����6 �_��Si����'����� ��L%���)��	.��M2�'�6�؜:���>�VtB��F�#�I���L���O���R��~U��X��hZ���\���^�I�`���b���d�1�f���h��k��qm�Ep� �r��u�*px�ZO{�. ~��k������삼���l�������Sᇼ����������u��<�������ߎ�.��=���u󒼐]��ŕ��%��q}��;˙�	���H���x��6���(����͠�[ܡ��ꢼj������'R�����!���n������g���������*>��`����#���x��Ʒ���Ḽ����# ��,���d����  �  13O=߳N=Z+N=��M=V�L=�PL=[�K==�J=a4J=�~I=��H=�H=rG=��F=�&F=7�E=�D=�LD=��C=�$C=�B=bB=�uA=��@=�A@=v�?=r�>=4)>=�c==#�<=~�;=�;=�B:=��9=��8=@8=��7=(*7=[�6=�>6=8�5=d5=��4=Iz4=>�3=qh3=��2=�(2=w{1=��0=O0=G]/=��.=��-=�=-=>�,=��+=�+=�S*=Ȑ)=3�(=]�'=�$'=KB&=RO%=�G$=(#=I�!=� =�"=Q�=��=�8=eq=V�=��=W�=�=�(=XI=�i=X�	=��=O�=��=&�=���<6`�<��<���<m`�<t��<�{�<��<v��<�"�<X��<�H�<���<[{�<T�<˽<ʂ�<�D�<��<�ڬ<��<�`�<n�<���<@+�<��<��<�Q�<ʦ�<G�<��v<��m<��d<�1\<��S<[gK<CC<y=;<>H3<�T+<lS#<�7<��<�
<�<���;L�;m��;W�;�;���;}�;*p;�LM;��*;N(;R��:�B�:.�
:�H�70
���������O���:#�m	E��1g�Ȅ�F�������.����ǻJ�׻/��_����� ��:��n�2���p�%!���%���)�+.�!b2�O�6��:�,t>�&0B���E�.I��=L�9O��R�a�T��SW�C�Y�� \��[^�d`�.�b���d�.�f��h�@,k�_�m��Ap�(	s�E�u��x�"�{���~�.ʀ����oW�� y������cs���R���%��V�(Ɖ�@���j������������莼�.��5���Dܒ�=7������U���Y+��p��ʯ��*뛼�!���R���|��A�������Zۢ������%���_��ۭ����������������]�������������_����㶼� ��ZD���Q��"M���=���*���  �  MO=Q�N=�N=��M=��L=�IL=m�K=��J=O=J=��I=2�H=�:H=4�G=C�F=�MF=4�E=P	E=|iD={�C=�2C=|�B=�B=�qA=��@=o6@=��?=�>=�>=�L==?~<=ͭ;=/�:=�:=�]9=��8=�8=��7=0�6=��6=�6=7�5=�K5=>�4=�h4=N�3=\3=R�2=�"2=z1=)�0=z0=�o/=�.=G.=�a-=�,=w�+=_7+=�s*=s�)=��(=](=�('=@&=9H%=�<$=�#=)�!=� =u=�y=��=`=-G=�p=��=e�= �=�==1@=�d	=�=�=��=��=�g�<�B�<�<���<]�<4��<���<�.�<U��<�e�<� �<)��<�/�<���<}_�<���<��<�\�<k�<�ڬ<ߙ�<vP�<���<;��<��<%q�<�ȍ<M�<p_�< _<Jv<,m<�d<m[<!�R<�J<7�B<�:<�2<�*<�"<��<U�<Ee
<�<��;-_�;�;|��;�M�;<��;���;E�r;k�O;�@-;k�
;��:X��:�x:@8_B��H��Hº�I��#�$�E�98h�Ki��Ҹ��t姻�ø��(ɻ��ػ�绪��˱���4��~��
�v��-^!�F�%��*�CY.��2��6���:�'`>�1B�pE��H��K�^�N��pQ��"T�j�V��FY�}�[�^^��N`�}b�7�d���f�Bi�K\k���m���p��Zs�rOv��Wy�]c|�F`�C��'x��:���Wׄ��ۅ��Ɔ����cf��&+��~�xʊ�ȳ��߳���ˍ�X����7��-����Β�����d�������痼�$���`�������ڜ�i���L���~��H���1բ�� ��Z3���s���ǧ�2��,����H����ę���D��%岼|s��J鵼�B���}������𡺼����z���^���  �  
O=h�N=�N=�}M=�L=\AL=��K=U�J=ABJ=c�I=��H=�PH=1�G=�G=UkF=^�E={"E=+~D=��C=X<C=.�B=*B=lA=��@="+@=Z~?=��>=�>=)9==|g<=��;=��:=��9=k:9=��8=/�7=t\7=�6=�j6=6=��5={65=��4=oX4=�3=�O3=<�2=�2=�v1=p�0=9%0=|/=W�.=q).=�|-=��,=N,=SR+=�*=ռ)=(�(=(=�)'=<&=-@%=�1$="#=G�!=�o =��=�b=�=&�=\%=oK=Xl=��=b�=��=a�=�=�F	=�k==o�=t�=�G�<,'�<��<���<4V�<���<��<�J�<��<���<39�<+��<?k�<��<���< %�<ù<zk�<B�<6լ<&��<�=�<���<�o�<��<�K�<0��<��<\%�<�~<��u<�hl<�}c<+�Z<�dR<�1J<>-B<�H:<et2<S�*<B�"<J�<��<6
<��<��;�]�;�.�;&�;Pܭ;]��;ό�;`�t;.�Q;�3/;�U;�:��:��:qa18:J���<����º���Ќ$�f�F�>-i������a����������`&ʻm ڻl��?��5?�7g�-��m��h�}�פ!�_&�Q*�ʇ.��2���6�J�:�/Y>�r�A�s<E��bH��^K�h9N���P�~�S��QV���X�Qj[��]��0`�Hub���d�k�f�J+i�9�k��n���p��s�7�v�D�y�w�|����b��D���� ���!��0#��	���؇�a���dY������튼�ҋ��Ό��⍼����C��儑��Ȓ�p
���G��J��������옼X&��d��ȥ���蝼U*���g��#����Ԣ�	��C�����᧼5O���Ԫ��n������˯�m}���$��ݸ���2��n����Ǹ�|⹼E⺼�ͻ�}���Ҋ���  �  ��N=��N=5N=ntM=��L=	;L=��K=:�J=wDJ=]�I=k�H=�]H=�G=G=�}F=��E=�1E=��D=��C=tAC=��B=`B=gA=�@=�"@=�t?=�>=y�==�+==5X<={�;=E�:=~�9=�#9=�r8=D�7=E7=�6=\V6=��5=ދ5=1(5="�4=M4=��3=�F3=��2=�2=�s1=Y�0=�(0=R�/=0�.=�7.=�-=��,=-$,=�b+=3�*=��)=j�(=U(=�)'=�8&=�9%=E)$=2#=	�!=jc =��=�R=N�=m�=m=�3=S=�q=z�=۶=��=;	=f3	=0Z=Jz=��=��=:1�<s�<V��<T��<MP�<���<���<C[�<
�<ߵ�<1\�<g��<���<��<���<;�<�ѹ<�r�<��<�Ϭ<��<�/�<Aϟ<�[�<�і<2�<��<��<"��<̆~<�.u<�l<�c<�nZ<�R<��I<��A<� :<-42<Fd*<+�"<�<`\<�
<q�<d�;�V�;,D�;�7�;�1�;+�;?�;��u;>S;�g0;ok;��:�@�:pw:m?8�:��'����púA�9%�+EG���i�&]���ԗ�.���:��j�ʻ��ڻS��2������A��=l����;���V���!�3&�!x*�]�.���2���6���:�fX>���A��E�66H�Z%K�Z�M�r�P��dS��V���X��<[��]�>!`��sb���d���f��Hi���k��;n�5�p�!�s���v���y�}����������0��AQ��+Q���3�� ��B���Zx��8��2���苼�⌼
􍼗��qM��$����ƒ����6��h��Q���|ʘ� ���@��n����͝���[��隡�<֢�z��KO��蘦���d���몼����L6���쯼����N���崼�a��B�������������c��μ������  �  <�N=^�N=c�M= qM=�L=�8L=�K=��J=EJ=T�I=� I=FbH=r�G=[%G=��F=��E=7E=ƎD=��C=CC=��B=�B=�eA=��@=�@=(q?=�>=�==�&==�R<={|;=��:=1�9=�9=�j8=�7=	=7=��6=SO6=��5=8�5=#5=��4= I4=:�3=�C3=��2=�2=Gr1=*�0=�)0=��/=��.=9<.=��-=��,=*,=xh+=��*=n�)=��(=\(=K)'=:7&=�7%=N&$=��"=��!=�^ =��=qM=1�=��=�=�+=tJ=�h=ǉ=k�=�=�=�,	=dT=u=ڋ=̖=�)�<��<��<\��<XN�<%��<���<�`�<>�<C��<h�<��<��<*�<��<B�<?ֹ<Yt�<��<�̬<�}�<�)�<Lȟ<�S�<ɖ<N(�<�t�<ٴ�<r�<�h~<�u<��k<��b<�LZ<��Q<�I<0�A<��9<�2<Q*<p"<�q<�N<�
<٤<&Y�;�T�;^L�;�J�;"O�;fR�;OF�;�=v;��S;�0;`�;�y�:{��:� :KB8vu���ŀ���ú�n�UG%�A�G��!j�U�������^���p���˻w�ڻd껓<��к�4�������t���j���!��B&�w�*��.�M�2�#�6�a�:��X>�o�A��E��'H�4K���M���P��LS�>�U��X��-[��]�b`��sb�1�d�/g�+Si���k�QJn�bq�#�s���v�z�1}�}#��y��������@���a���`���B�����iʈ�4����A��������錼H������JQ�����$ƒ����1��`��.������������4���z���ĝ�e���V��_��� ע�����S������j����k��1��������@��Z�������^\�������q���ͷ������`��� ���ڼ�����  �  ��N=��N=5N=ntM=��L=	;L=��K=:�J=wDJ=]�I=k�H=�]H=�G=G=�}F=��E=�1E=��D=��C=tAC=��B=`B=gA=�@=�"@=�t?=�>=y�==�+==5X<={�;=E�:=~�9=�#9=�r8=D�7=E7=�6=\V6=��5=ދ5=1(5="�4=M4=��3=�F3=��2=�2=�s1=X�0=�(0=R�/=0�.=�7.=�-=��,=-$,=�b+=3�*=��)=j�(=U(=�)'=�8&=�9%=J)$=9#=�!=xc =�=S=p�=��=�=�3=^S=r=�=_�=y�=�	=4	=�Z={=c�=ܛ=�2�<2�<	��<��<�Q�<���<���<B\�<�
�<l��<�\�<x��<ɏ�<��<��<5:�<�й<Wq�<1�<ά<䀨<�-�<�͟< Z�<0Ж<�0�<A~�<࿈<.��<R�~<�-u<	l<�c<RoZ<�R<f�I<��A<>:<�62<4g*<S�"<7�<�_<b
<��<gj�;s\�;lI�;<�;i5�;�-�;�;Q�u;�=S;Pe0;g;_��:�0�:P:�4<8����������úP�i %�OTG���i�Nd���ۗ�f4���@����ʻj�ڻ�������V�����am������wW�Z�!�n3&�xx*���.��2��6���:��X>���A��E�C6H�d%K�b�M�x�P��dS��V���X��<[��]�?!`��sb���d���f��Hi���k��;n�5�p�!�s���v���y�}����������0��AQ��+Q���3�� ��B���Zx��8��2���苼�⌼
􍼗��qM��$����ƒ����6��h��Q���|ʘ� ���@��n����͝���[��隡�<֢�z��KO��蘦���d���몼����L6���쯼����N���崼�a��B�������������c��μ������  �  
O=h�N=�N=�}M=�L=\AL=��K=U�J=ABJ=c�I=��H=�PH=1�G=�G=UkF=^�E={"E=+~D=��C=X<C=.�B=*B=lA=��@="+@=Z~?=��>=�>=)9==|g<=��;=��:=��9=k:9=��8=/�7=t\7=�6=�j6=6=��5={65=��4=oX4=�3=�O3=<�2=�2=�v1=p�0=9%0=|/=V�.=p).=�|-=��,=M,=QR+=�*=Լ)=(�(=(=�)'="<&=3@%=�1$=0#=Z�!=
p =�=�b='�={�=�%=�K=�l=j�=?�=��=��= =)H	=m=V�=�=$�=
K�<�*�<���<��<Y�<w �<i��<�L�<���<���<�9�<L��<�j�<M��<���<O#�<���<i�<��<EҬ<��<�:�<�ݟ<�l�<��<I�<���<}��<�#�<?�~<��u<�gl<�}c<�Z<�fR<Q4J<�0B<[M:<|y2<��*<\�"<��<%�<�<
<�<B��;�h�;�8�;�
�;��;ֽ�;n��;��t;��Q;X//;LM;���:���:�a:��+8���}q���ú���(�$���F��Ii�����n��Ѷ��鰹��0ʻ�	ڻ���F��HB��i�b��o�;j�� �ڥ!�0&��Q*�P�.�q�2��6���:�bY>���A��<E��bH��^K�w9N���P���S��QV���X�Uj[��]��0`�Jub���d�l�f�K+i�:�k��n���p��s�7�v�D�y�w�|����b��D���� ���!��0#��	���؇�a���dY������튼�ҋ��Ό��⍼����C��儑��Ȓ�p
���G��J��������옼X&��d��ȥ���蝼U*���g��#����Ԣ�	��C�����᧼5O���Ԫ��n������˯�m}���$��ݸ���2��n����Ǹ�|⹼E⺼�ͻ�}���Ҋ���  �  MO=Q�N=�N=��M=��L=�IL=m�K=��J=O=J=��I=2�H=�:H=4�G=C�F=�MF=4�E=P	E=|iD={�C=�2C=|�B=�B=�qA=��@=o6@=��?=�>=�>=�L==?~<=ͭ;=/�:=�:=�]9=��8=�8=��7=0�6=��6=�6=7�5=�K5==�4=�h4=N�3=\3=R�2=�"2=z1=)�0=y0=�o/=�.=F.=�a-=�,=v�+=]7+=�s*=q�)=��(=](=�('=#@&=AH%=�<$=�#=E�!=2� =�=/z=��=�=�G==q=��=p�=9�=}�=�=�A=�f	=��=(�=S�=�=�l�<�G�<��<���<+a�<���<ɗ�<�1�<x��<lg�<|�<X��<3/�<���<�]�<6��<(��<}Y�<��<V֬<{��<�K�<N�<Ɔ�<x�<+m�<�č<*�<�\�<[<�v<��l<td<Nn[<��R<ҾJ<Y�B<[�:<;�2<�*<�#<��<��<�n
<�< ��;$o�;l�;㱾;�W�;��;��;�r;��O;e:-;t�
;���:�_�:':E8�V��o:��R`º�r��	$��F��`h��|��a˖������Ӹ�7ɻ��ػ��综&��#�����S����9���_!�n�%��*� Z.���2���6��:�p`>�jB�KpE�A�H��K�s�N��pQ��"T�s�V��FY���[�c^��N`�}b�9�d���f�Di�L\k���m���p��Zs�sOv��Wy�^c|�F`�C��'x��:���Wׄ��ۅ��Ɔ����cf��&+��~�xʊ�ȳ��߳���ˍ�X����7��-����Β�����d�������痼�$���`�������ڜ�i���L���~��H���1բ�� ��Z3���s���ǧ�2��,����H����ę���D��%岼|s��J鵼�B���}������𡺼����z���^���  �  13O=߳N=Z+N=��M=V�L=�PL=[�K==�J=a4J=�~I=��H=�H=rG=��F=�&F=7�E=�D=�LD=��C=�$C=�B=bB=�uA=��@=�A@=v�?=r�>=4)>=�c==#�<=~�;=�;=�B:=��9=��8=@8=��7=(*7=[�6=�>6=8�5=d5=��4=Iz4==�3=qh3=��2=�(2=v{1=��0=N0=F]/=��.=��-==-=<�,=��+=�+=�S*=Ɛ)=2�(=^�'=�$'=PB&=[O%=�G$=2(#=k�!=M� =$#=��=�= 9=r=8�=��=��=I
=�*=KK=	l=��	=<�=	�=v�=�=��<f�<E#�<��<ve�<��<��<?
�<��<b$�<d��<�H�< ��<�y�<!�<#Ƚ</�<�@�<�	�<�լ<���<\[�<��<��<&�<&��<���<'N�<���<��<-�v<�m<��d<u3\<�S<)lK<cIC<E;<Q3<p^+<�]#<C<<Z�
<�<���;�_�;��;�+�;m��;b�;P��;p;�KM;ə*;�;���:=�:/1
:E�7�\��U��a���g��m#�<E��cg�����
�����������ǻ@�׻N�滴�����?������՝��r��!� �%���)��+.��b2���6�Y�:��t>�l0B�ۻE�XI��=L��9O�R�p�T��SW�L�Y�� \��[^�i`�1�b���d�0�f��h�A,k�`�m��Ap�)	s�E�u��x�"�{���~�.ʀ����pW�� y������cs���R���%��V�(Ɖ�@���j������������莼�.��5���Dܒ�=7������U���Y+��p��ʯ��*뛼�!���R���|��A�������Zۢ������%���_��ۭ����������������]�������������_����㶼� ��ZD���Q��"M���=���*���  �  DHO=��N=�8N=8�M=} M=1TL=�K=(�J=b&J=�hI=�H=��G=9GG=2�F=��E=KWE=w�D=V)D=��C=vC=��B=� B=vuA=��@=dI@=b�?=l�>=�:>=�y==��<=�;=�,;=bp:=ݼ9=�9=bu8=a�7=�Y7=��6=c6=`�5=~|5=�5=ω4=�4=�q3=��2=�*2=x1=��0=�0=�D/=}�.=��-=~-=cX,=��+=��*=�,*=p)=Ұ(=9�'=a'=Z@&=�R%=�O$=�3#=O�!=�� =�9=x�=�=ka=�=��=��=h$=�D=�b=0=L�=��	=��=�=��=K�=���<�~�<�4�<���<_a�<���<s]�<���<R�<���<WY�<x��<E~�<7�<���<a��<�K�<��<��<�ˬ<Ꝩ<�c�<��<��<�C�<*��<�(�<>��<h��<�X�<4�w<��n<?�e<�]<��T<=,L<f�C<#�;</�3<6�+<��#<p�<�8<��
<^+<m��;q*�;"W�;bu�;���;�ə;��;h�l;�J;<p';.;
��:�׃:��:ь�6�~ �X���º_��6#�G�D�цf��J���G�����H�����ƻ�"ֻ������; �o���m�����*����� �{N%�ض)��
.�ON2�ɀ6�X�:��>��tB��F�S�I���L��O��R��~U��X��hZ���\���^�M�`���b���d�4�f���h��k��qm�Fp�!�r��u�*px�ZO{�. ~��k������삼���l�������Sᇼ����������u��<�������ߎ�.��=���u󒼐]��ŕ��%��q}��;˙�	���H���x��6���(����͠�[ܡ��ꢼj������'R�����!���n������g���������*>��`����#���x��Ʒ���Ḽ����# ��,���d����  �  �YO=��N=�@N=��M=�M=RL=U�K=��J=�J=�MI=�H=��G=�G= hF=��E=�#E=O�D=� D=qyC=�B=�vB={�A=�oA=��@=�K@=٩?={�>=H>=o�==��<=E<=%T;=��:=`�9=;J9=��8=�8=Ȋ7=�7=��6=�6=ܑ5=5=��4=�
4=vu3=H�2=K'2=�o1=�0=�/=T'/=@b.=t�-=�,=$,=_k+=$�*=> *=K)=J�(=��'=j'=�8&=�P%=;R$=�9#="=�� =�L=V�=�2=�=��==
=:=`a=Ł=�=(�=��=��	=��=��=��=��=���<��<�:�<���<uR�<���<E0�<x��<��<�u�<(��<
{�<W�<L��<�p�<8�<��<��< Ӱ<޶�<���<g`�<��<�Û<X�<�ܒ<�U�<�ȉ<<�<���<zfx<�{o<�f<L�]<�bU<��L<��D<a_<<&74<�,<��#<�<�V<��
<c)<���;���;���;���;�p�;�b�;�x�;G{i;�sF;��#;��;���:��}:���9��������m����º����"�[SD�c�e�w҃�[����-���o���EŻ��Ի�T�ao����������kn�d������� ��'%�8�)� .��P2�z�6���:���>���B��F��/J�h�M���P��S�WSV�x�X�v[��?]�=_�!a���b���d�ɿf��h���j�TWm���o�s�r�W=u��x���z��x}�D��jL���~��8���z���@������Y���b���6r��|c���b���u��]�������Y8��N��������������u���ژ�f1��Fy��t���1ڝ�d���������������+��.%���O��>����騼�V��fӫ��Y��*㮼�h���屼{V��2���
��pK���|�����Q������VǼ��  �  �eO=c�N=�BN=E�M=�L=�IL=ӋK=��J=��I=�.I=�dH=g�G=,�F=�1F=j�E=$�D=�\D=��C=�TC=��B=b`B=�A=AdA=�@=nG@=�?=] ?=�O>=�==r�<=�+<=_x;=�:=y!:=�~9=��8=~J8=�7=&-7={�6=�#6=��5=H 5=��4=N4=�r3=S�2=�2=b1=u�0=�/= /=�9.=�p-=3�,=��+=�4+=.�*=)�)=�")=4r(=�'=��&=),&=�H%=FN$=p9#=o	"=l� =�Y=w�=�N=�=��=8==;r= �=O�=t�=V�=��=��	=�=�=r=E�=��<��<H4�<s��<�8�<��<���<ES�<��<��<Y��<Y
�< ��<�N�<��<H�<5ȸ<O��<C��<ʖ�<I{�<�P�<T�<�<2a�<��<�y�<��<���<��<�+y<�Sp<-�g<�^<r1V<��M<�3E<!�<<�4<�U,<�$<f�<�Z<��
<<8Q�;>�;��;,��;�/�;��;�Ȅ;��e;F�B;�? ;���:���:�Is:*@�9|�<��C
����� |ĺe��R#��gD�%�e�s���@��4`��	b����ûӻ<��h��?Q����j0���&d����j ��%�͠)�9.�>l2���6���:��*?��9C�k G�}�J��MN���Q��|T�{0W���Y���[�	�]�P�_�J�a�tJc��e���f���h�Pk�cVm�_�o�O[r���t���w�oHz���|�5`�j瀼����7��PQ���`���f���d��>]��^U���R��\���v�����BN������A���ǔ��M���˗��<��(����盼����@��)P��	P��FE��N6��*��4(���6��sZ��]���{樼�J��K���E5��u����%�����������P�������㶼���/K��?o������*����  �  �lO=U�N=?N=�M=��L=$<L=�zK=��J=j�I=4I=�=H=�sG=��F=D�E=�TE=�D=,D=V�C=K/C=��B=GB=��A=$TA=>�@=�=@=R�?=��>=�Q>=G�==��<=�B<=v�;=-�:=M:=��9=H9=�w8=��7=�O7=@�6=o66=̭5=�$5=�4=\4=bj3=��2=12=�O1=��0=��/=��.=.=WB-=�y,=�+= +=�N*=�)=��(=�O(=0�'=��&=&=�;%=�D$=O3#=�"=b� =�a=��=�d=D�=)"=Kj=g�=��=��==�==?
=%=�==��=1��<��<n"�<I��<��<�q�<L��<�<XZ�<���<��<���<{5�<���<а�<:��<U��<Uz�<�v�<�n�<�Z�<�6�<���<y��<�_�<n��<���<�&�<���<S�<�y<�q<�Th<��_<��V<�FN<�E<I>=<��4<~,<&$<��<#G<�
<��<��;���;��;ꅺ;��;�k�;h$�;�Ub;r?;��;o=�:��:�h:��9נ�����/��3�ƺ�v�z�#���D��e��W��9���i����z����»��ѻ�U��c�e����x��
������_�2\ ��%���)�E4.�<�2���6��I;��?��C�׬G��yK��O��RR�*RU�>X��qZ��\���^�T`�%b��c��Ye�j$g�i�C+k�lm���o�LKr��t�E^w���y�dW|�ٿ~�n��������ق����O��'���4��=���C��lM���`�����鹍�-���m��l葼�r�����(����!��ۜ������R���������ê�����Ň���l���U��K��tR���o��������I��8������y����쯼�K����������O@��Ȇ���Ƿ�����4���_�������  �  �nO=%�N=�7N=Q�M=J�L=2,L=#hK=��J=F�I=T�H=3H=AKG=]�F=��E=o%E=��D=� D=�C=�C=ÜB=�-B=��A=BA=�@=�0@=]�?=�>=�O>=��==��<=1T<=��;=+;=�p:=|�9=�89=e�8=/8=k7=��6=�C6=�5=6%5==�4=��3=�^3=δ2=n�1=<1=Ko0=$�/=M�.=��-=�-=�L,=�+=/�*=�!*=4y)=��(=�/(=�'=�&=j&=�,%=?8$=�)#=� "=�� =3d=��=�t=��= A=d�=��=��=�=/=�6=�6=�1
=l)=4=v=?�=���<lp�<(
�<��<$��<D�<~��<���<b�<=]�<���<�<�<��<g��<6[�<C�<=�<{@�<\E�<D�<6�<��<��<t��<XV�<F��<���<	E�<i�<n��<Qkz<�q<��h<>`<�W<T�N<�F<9�=<�5<Ƒ,<�#$<Ȯ<�$<�x
<��< ?�;���;�H�;Ć�;��;`�;��;U8_;��;;)�;�G�:i"�:��^:���9?�ָ5�/���-ɺ�|��$�VhE�f��O��'i��@���Ĳ�����)�лe)߻j2�j������B
��?����SJ��^ �6%���)��e.���2��?7�1�;���?�]D�X0H�GL�x�O��S��V�N�X��([��D]��$_���`�+sb�{d���e�
ig�Mi��Zk���m�/�o��Lr���t�l,w�-�y�5�{�j<~�'C��g������t���Ԅ���W��C'��S;���P���l��N����ҍ�G&��b���F������B?��mۖ�jo��.�`�������坼���������砼�ơ����炣�*q���r��B�������B���GQ��V������h��I�������^������`��9��с���Ƹ�����@���t���  �  nO=:�N=a/N=a�M=M�L=HL=WK='�J=�I=��H=9�G=�*G=HcF=��E= E=.gD=��C=DbC=f�B=��B=TB=��A=�1A=i�@=T$@=�?=f�>=�K>=6�==�==�_<=n�;=�%;=��:=]�9=�U9=,�8=�8=�~7=�6=$L6=�5=#5=�4=��3==S3=3�2=��1=d*1=$[0=�/=��.=��-=��,=6),=e+=B�*=�)=X)=ֶ(=c(=7n'=v�&=��%=�%=�+$=t#=��!=�� =�c=d�=(=I�=SW=��=��=b=
==hM=xQ=tL={A
=/3=`"=�=��=®�<k\�<���<�l�<0��<<�<�Z�<��<f��<��<w�<���<7��<aA�<�<��< �<
�<��<g�<��<���<pΟ<[��<�J�<���<��<"Y�<�	�<Q��<��z<d-r<�xi<�`<��W<b(O<�iF<��=<;!5<Ǘ,<�$<ܓ<J�<�H
<�i<���;�I�;���;q��;Υ;D�;��;��\;�m9;�;��:nƪ:M�V:�Դ9\-�Ӂ�#g���;˺�o�e�%��F��tf��Y��|F��[C��D����ϻ�I޻�N컐��������	��	�����A�j �%Q%��*�h�.�t3��7���;�;@��|D�@�H�߉L��7P���S�A�V��YY��[���]���_�!Ea��b��Zd���e���g���i�t�k�O�m�b�o�lWr���t�Dw��[y�)�{�&�}�&���,��Q���z��ץ��aЅ�����7��19���W��^{�������덼�B�����T7��[Γ�p�� ��󭘼�7������L����/���D��>��g"��s���)Ϣ�/�������5��������Ч�����[��������\U��1����簼,���o������� ��;N������G湼�+���k���  �  �lO=�N=�(N=7�M=��L=�L=:KK=�yJ=�I=��H=>�G=�G=�LF=��E=!�D=�OD=��C=�MC=��B=�sB=�	B=͛A=�%A=�@=@=�?=i�>=6H>=��==�==vf<=��;=u3;=қ:=0:=h9=Q�8=�*8=Պ7=Y�6=�P6=ͷ5=� 5=$�4=��3=�J3=`�2=��1=1=fM0=jt/=@�.=U�-=�,=J,=qM+=��*=�)=�B)=J�(=(=�^'=�&=��%=�%=�"$=�#=��!=�� =�b=t�=�=��=�d=D�=��=�1=Q=`=�a=6Y=�J
=G8=�#=B=��=\��<�L�<���<X�<L��<� �<;�<%o�<��<8��<�G�<���<�X�<v�<.�<�ݻ<
�<��<9��<��<���<$�<ȼ�<f��<QA�<E��<���<wd�<#�<�Ձ<{{< wr<��i<Ca</4X<�aO<R�F<��=<>.5<C�,<0$<�}<i�<%
<{@<[�;"��;f�;D'�;�.�;�V�;2�;z1[;�7;ޅ;��:���:#�Q:���9=��-0 �i��1�̺��/&�5xF��f��e��K6��������������7rϻ��ݻ�뻴p��_^��	��������?��t ��f%�R#*�_�.�:3��7�+<�"s@�	�D�1�H�?�L�o�P�f�S��W���Y�\�#^���_�r�a�Nc�Βd��$f��g���i���k�O�m�ep��ar���t��v�#<y�	q{���}�x��p���-���Y��ȉ��庅��醼����9��0^��݆��칌�����LW���Ȑ��P��듼�����7���֘��c���כ�#,��i_��r��Qh���H�������ţ���������⸦��᧼����d������� ���J��򎯼�ΰ����M��K����ݵ��.������9ӹ�d ���g���  �  �wO=��N=;N=j�M=��L=�'L=6XK=�xJ=��I=��H=��G=�F=<�E=�*E=�D=��C=�qC=�	C=�B=�]B=B=~�A=:KA='�@=�N@=t�?=s?=Jz>=k�==�===�<=�<=�;=J;=Pv:=��9=�A9=G�8=��7=kR7=/�6=�6=��5=��4=�e4=L�3=�#3=rk2=R�1=#�0=,�/=��.=m.=+)-=;T,=�+=b�*=^D*=D�)==4)=t�(=�/(=��'=�&=�2&=HP%=�M$=�,#=��!=�� =r:=��=BD=ұ=�=�Q=~=]�=ˍ=lx=�W=j1=�
	=��=8�=,�=6| =���<��<�q�<���<���< ��<e��<w��<C��<��<$^�<��<���<��<�<���<�<��<F0�<]8�<�%�<S��<J��<�p�<�#�<�ڎ<.��<U`�<�(�<��{<Es<ŋj<Ψa<��X<&�O<�F<O�=<�4<�	,<�u#<s�<�Q<��	<�� <ک�;,��;;"�;_�;`��;{�;�3s;��M;�);�;���:o-�:\:��9d��!�K�!颺�u�p��EV1��GR��8s��艻3登z���9���6�ǻ5.ֻN�仦��s �/X�W��^��\�?��L(%��*�=�.��3��7�b�;��c@���D��UI�	�M�m�Q��U�=&Y�g-\��^���`���b�R�c�e�� f�0g��_h�m�i�<ik��Lm�/co�Z�q�<�s�#v�?x�eLz��F|��;~�����*���I���z��H�������64���f��ꍉ�����nʋ����-��1���X��ա���\���)���������Xl��D���`Q���}���{��6Q��v��$����P��+����ä���������ا�t���d�����������:��!l��ٔ�����벼)���w���ն�;��x�������O���  �  OzO=l�N=�?N=ɛM=y�L=�-L=�^K=�J=9�I=��H=O�G=+�F="�E=P6E=�D="�C=Q|C=�C=2�B=�eB=mB=B�A=�QA=3�@={T@=��?=!?=�}>=V�==�===�<=�<=V�;=�:=3n:=��9=�99=ږ8=7�7=�O7=u�6=�6=ъ5=�4=�j4=��3=�)3=�q2=ۧ1=6�0=��/=O�.=�.=�3-=W_,=��+=��*={O*=��)=�=)=�(=n7(=}�'=P�&=�8&=�U%=�R$="1#=n�!=� =;=_�=�@=F�=?=�H=�t=�=�=q=�Q=�-=a		=2�=�=.�=� =���<2�<5|�<��<���<���<O��<s��<��<M�<tu�<� �<���<؟�<]��<Uɷ<K��<�!�<R?�<�F�<�3�<�<�ƛ<�y�<�)�<eݎ<t��<-Z�<��<@�{<@$s<Thj<D�a<ӅX<yO<�qF<�=<˶4<|,<S�#<��<�b<*�	<�� <z��;���;�[�;d��;�֠;�5�;O�s;�|N;k*;1�;)Q�:C��:W�:�t9&����oI�����I���0���Q��r�Љ�{ݙ�����Ѹ���ǻFbֻ+�仓�x� �p����h�*^�D���%�$�)���.��3�uk7��;��H@�!�D�O6I��M���Q�D�U�a�X�e�[��^���`�
db�w�c���d�� f�Ng�(Eh���i�XQk�:6m�6Oo�C�q�)�s��v�Ax��Vz��X|��T~��,��#;��.Z��R���Ä� ���8��g��p�����������a猼X"��&{������l���ON��t��藼ԫ��W���ޜ�i:��g���e���<������"���4A��>𣼦�������夦�'ͧ����]������0���c=���r�����nʱ�y����9��̇���㶼�E��n���� ���M���  �  S�O=i�N=�LN=��M=��L=�>L=�pK=�J=u�I=��H=��G=w�F=�F=�WE=��D=5D=��C=�0C=�B=�|B=0'B=-�A=LcA=��@=Ud@=�?=H-?=��>=W�==�===��<=�
<=�x;=T�:=�U:=�9=�"9=b�8=��7=�F7=��6=�6=;�5=%5=1x4=�3=�93=ւ2=(�1=�0=��/=�/=a0.=�Q-=�,=ֽ+=+=�o*=��)=%Y)=u�(=
M(=η'=�'=I&=e%=�`$=^=#=�!=�� =T<=�=06=��=i�=/=�X=7l=�k=�[=�A=�#=>	=Y�=��=�=9� =s��<i;�<֚�<���<W��<���<z��<�<�!�<�Z�<��<2E�<���<�ݿ<��<��<A%�<�L�<�g�<�l�<�W�<q(�<��<��<�8�<�<�<�E�<Q��<Lg{<�r<��i<�a<*X<�.O<x=F<Yf=<B�4<�,<̞#<"$<��<{�	<�� <u^�;3f�;=�;&_�;ǯ�;�(�;��u;j�P;��,;t

;���:K��:�&:��59�敹f�C��N��:޺H���/��P�A3r�F���4Ι�ݫ��Z$��k=Ȼ�׻ˈ����� �m��QJ�a��f�-����$�r�)�@W.���2�$(7�Z�;���?�mrD�6�H�})M��?Q�U�OwX��x[�!	^��*`��a��Wc���d�ӧe���f�#�g��ei�sk�r�l�o��\q���s��v�=Ix��vz�a�|���~�AZ��yl���������焼S���E���h��~���q��������ʌ�����Y���Ӑ��n��>%���땼鴗��r��5��˜�����R$��&�����鿡�!m��>��Yɣ�y���nz������<�����PH����������oE����������:󱼰*��gk��}���L��Vf��Լ��(
���K���  �  �O=P�N=�]N=ҾM=�M=zVL=�K=خJ=��I=G�H=0�G=�G=�IF=>�E=%�D=cLD=��C=�\C=[�B=g�B=�EB=V�A=3|A=,A=z@=��?=�=?=��>=��==�:==^�<=�;=�[;=��:=a.:=��9=�8=5c8=.�7=I77=�6=o 6=8�5=�5=��4=��3=P3=�2=$�1=��0=f0=�;/=0Z.=�-=P�,=��+=�A+=��*=*=��)=C�(=m(=��'=�&'=�_&=�y%=�s$=�M#=`
"=�� =�;=��=�#=�=��=&=�+=l?=TB=�8='=�=u�=��=��=��=c� =���<@b�<���<��<�+�<�=�<PJ�<�\�<��<��<~$�<���<gc�<�=�<\8�<�J�<uj�<Պ�<���<ա�<]��<V�<>�<G��<J�<g�<��<�!�<�ǁ<6�z<�r<�Si<�x`<d�W<�N<k�E<<1=<�4<�),<��#<]<��<>,
<S?<Q�;o>�;F��;��;���;���;�1y;�T;�)0;�};�'�:��:8	2:�p]9�+����;�ؗ��{�ںN{��[.�ŶO��@q�FS���͙�F�������;ɻ�ػ��k��hz�6����M��d|������$���)��	.��n2��6�\+;�{�?��C�YH�m�L���P��OT�C�W�V�Z�^7]�a_��-a���b��c�D#e��Mf���g��i�j�j�ףl���n�c q���s�2�u��_x�h�z���|�m�Ȥ��Ӽ���ڂ������"���D��/_��p���x��S~��k�������׍��+��#���*9��3铼����og����������6��E�������Kß�h���n���$���֢����\_���J��X��>���?Ш�^-��q��������V�����J�c6���w��6���\���Q��霸�,⹼[��|M���  �  �O=��N=gnN=��M=;)M=HoL=^�K=�J=��I=�
I=�*H=�RG=~�F=��E=�#E=�D=WD=@�C=@*C=��B=�hB=�B=��A=�A=%�@=(�?=LM?=y�>=��==3==��<=��;=�3;=F�:=��9=/`9=��8=�68=J�7=}7=y�6=86=͡5=�"5=j�4=�	4=�g3=c�2=��1=Y1=�E0=�h/=��.=��-=�,=63,=��+=��*=H*=p�)=�&)=��(=|�'=�A'=\w&=�%=4�$=�\#=�"=� =)6=��==�X=t�=��=@�=8=�
=�=A=q�
=�=��=�=��=� =J��<k��<���<O;�<�j�<R��<r��<���<���<�B�<���<\6�<v��<���<��<q��<c��<�Ѱ<M߬<�ڨ<p��<r��<�1�<�ʗ<jV�< ܎<b�<�<�z�<"z<rCq<�lh<�_<��V<�	N<3dE<��<<�v4<k',<�#<Ǐ<�<m{
<��<���;�1�;!�;�۷;���;t�;�@};�nX;��4;��;�p�:�;�:��?:]{�9��^��2�)}����ֺ�����,�tN��_p��$����,q��z���Dʻg�ٻT�#����@����F-���J��^��3�$�	O)�>�-��2��i6���:�h?��wC���G���K�T�O��eS�y�V�|�Y�.\�b^�B`�f�a�!@c��d���e��g��h��Uj��Nl�ǃn��p��ms���u��x�{��u}�����	��j)��PF��[`���u��=���)�������v��@l��|k�� ~��/�������5m������s����V��$	�� ����A��A����	���9���F���4���	��6Ρ�����Q���'�����X*���]��X������ȉ������t���ޯ��=������y೼^)���n������^鸼;���=���X���  �  5�O=�O=yN=a�M=u:M=$�L=ҼK=��J=�J=�6I=�_H==�G=9�F=�F=nE=��D=�KD=�C=A]C=��B=��B=�B=��A=�.A=֠@=�@=�V?=�>=��==�#==jg<=��;=� ;=�X:=��9=N9=��8=��7=�{7=��6=��6=�6=ʡ5=�)5=��4=\4=�y3=;�2={	2=�=1=�k0=M�/=e�.=��-=E6-=�|,=/�+=�&+=-�*=Y�)=wU)=g�(=((=LY'=(�&=z�%=��$=�e#=."=_� =�(=�=��=4'=�]=�=d�=��=��=��=�=y�
=[�=��=��=��=v� =��<!��<��<i�<\��<���<��<�:�<s}�<$��<IC�<���<�t�<;8�<e�<A
�<��<o�<H�<�
�<|�<d��<�M�<Rڗ<~U�<6Ǝ<�3�<���<��<J.y<�9p<;Vg<a�^<��U<�4M<ƼD<g<<�.4<O,<T�#<��<�I<
�
<��<��;��;�<�;�D�;<M�;y�;7�;M];q�9;>�;���:5��:%N:�/�9x�5�=*��Γ�t�Ӻ�T
�Ɯ+�S�M�G�o��(��cK���.��{�����˻kMۻ�H�c���%2�x�	���������?��M�$�-)�s�-��1�X6�j:��>���B��!G��K�V�N�lcR�ݔU�MuX�E[��D]�@=_���`��b���c�DJe�G�f��Gh�ej�Kl�:Qn���p�@js�/ v� �x�߈{��"~��Q��o���֬���ȃ��؄�݅��Ԇ�W����������g��pY��9c��]����Վ��@��ȑ�Fb�����!���6:��M���5&���t������+���緟�����=t��D��������j�\���?������&
��v���������\%������Y��q_��m����A#���I���b���n��r���  �  B|O=5 O=zN=��M=�AM=��L=��K=B K=�/J=X_I=�H=��G=JG='aF=�E= E=�D=�
D=7�C=�C=¦B=�3B=]�A=l8A=��@=�@=�V?=�>=��==�==�C<=��;=!�:=E:=Co9=}�8=4E8=��7=�F7=��6=�j6=�6=��5=�'5=��4=�4=��3=��2=J2=-V1=�0=$�/=�.=�9.=~-=��,=,=�n+=��*=R%*=Y�)=o�(={((=�h'=Ó&=��%=�$=<d#=�"=� =~=Hm=д=�=�=�:=-U=�i=�z=��=M�=��
=��=m�=<�=>�=�� =�<4��<'�<)��<9��<Y�<�a�<���<Z�<�i�<���<�i�<�<���<J��<�e�<�S�<J�<�>�<�(�<���<z��<�U�</ח<-B�<���<$�<�J�<���<� x<o<�f<1U]<B�T<>L<j�C<��;<�3<��+<н#<�<�L<��
<� <,	�;r��;U2�;%��;��;��;�7�;�Ub;p�>;"�;= �:���:�Q\:!*�9���86#�)���{Ѻ9�	�k�*��.M�J�o��s���ꚻ�.����=�ͻTݻ-{�=���)C�ݩ
�>���4��a�)9 ���$�x0)��y-��1���5��6:�~o>��B�ŘF�mJ�TN��^Q�arT��BW���Y�q \��5^��`��a��^c���d��pf�Kh���i�%�k��Fn���p�k�s�;dv��Hy�d'|���~��̀����
@���Z��ya���T��o6��A
���Ո�k���Bt���Z��N\���~��Î�\&��⡑��+�������E��^ŗ�/5�����ۛ�����.��j:��}4��� ��L��ꢼ�أ��ڤ�0���,6��.���b������}A��;⮼�|��
��/���?hA���~��ئ��ź����������6����  �   gO=}�N=�oN=��M=d=M=�L=��K=�K=
FJ=�I=��H=�H=�TG=?�F=�F=9gE=��D=,AD=,�C=�7C=��B=_>B=��A=�6A=��@=�?=�K?="�>=ٽ==��<=�<=�K;=݆:=�9=M#9=��8=h�7=�}7=7=��6=�F6=��5=Ӆ5=u5=��4=|4=�~3=��2=5!2=re1=��0=��/=\-/=v.=G�-=9-=�a,=��+=v+=�V*=�)=��(=�6(='n'={�&=��%=u�$=uW#=� "=$� =A�=D=��=��=��=[�=� =�=+=�A=!Z=�s
=�=\�=��=�=v� =9��<��<<#�<���<*��<�R�<ȱ�<��<D��<h��<�v�<��<��<�7�<��<ճ�<!��<@m�<R�<0�<��<��<�F�<ƾ�<�</f�<=��<P�<�+�<w<��m<��d<�\<a�S<x5K<0C<�;<73<n[+<fp#<b<�!<ǧ
<"�<$�;r�;���;���;t{�;d�;�k�;�)g;��C;�� ;.�:ܸ�:w�h:ۇ�9�S츿��y؏�G�к�k	��+���M�	�p����nʛ�Rd��X����dϻ&y߻���:��0b����D��������� �J%��^)�֘-���1�" 6�/:��O>� TB��.F��I�>M�(kP�d^S��V���X�=
[��>]��I_��-a���b���d��Pf�jh�4�i��l�qin��q�C�s�Z�v���y���|����<R��.���Xك�T�K�\Ն�9���-a�����"Љ�q����q��ql��:���!ǎ�!������_��s��e򕼪Z��$������@G���}��]���ƞ��֟�۠��֡�VϢ��ͣ��ڤ�+ ���C�������-��̫�{���/���߰�H������׃��,۶���12��5��*"��t ���ؼ��  �  �JO=F�N=\N=��M=/M=��L=��K=�K=mSJ=�I=�H=�7H=ȎG={�F=�FF=o�E= 	E=�oD=��C=NC=��B=�?B=��A=^+A=|�@=m�?=R7?=�q>='�==��<=�;=?;=�G:=]�9=��8=K=8=��7=�;7=��6= u6=�6=L�5=Vk5=�5=��4=+4=Jq3=��2=�2=�k1=��0=�0=uV/=�.=��-=R-=�,=.�+=�9+=��*=E�)=�)=�<(=�j'=��&=>�%=-x$=?A#==�!=�j =I�=�=4J=�m=��=9�=��=��=��=��=y=#>
=d_=b{=��=r�=� =Q��<�}�<��<z��<�<�x�<���<o�<'��<!w�<r��<���<s�< ��<A�<S�<��<�}�<�Q�<]#�<j�<ꔠ<�$�<���<��<I"�<�P�<C|�<�_<��u<L�l<i�c<��Z<2gR<.J<�-B<�W:<~�2<5�*<�#<}<��<7d
<#�<���;�1�;�W�;ր�;��;�;�^�;�zk;�=H;M%;��;Cf�:�ts:3_�9�ȸϛ��ď�GyѺ5�	�r�+���N��q�gՊ�x՜������C���Gѻ��&�v~���y�X��g�T�����!�/u%���)���-�	2��06��M:��T>�7B�4�E��\I���L�@�O�EjR��U���W��Z��h\���^���`���b���d��Uf��0h�b(j�hOl�8�n��Xq��:t��Jw��tz��}��\�� Ձ��1���m�� ����}���T��D��$���Bc������Ɗ�B���@���駍��ގ��.��������/U������8 ��9G������eÚ����� 2���a��3�������L����Ƣ�nգ��3��ue���Ϩ�-[��s�����������F������K���#��Gp��)�������v���2���wW��2���  �  �+O=�N=VCN=,�M=)M=DrL=�K=�K=�YJ=��I=*I=�^H=�G=uG=x}F=�E=�6E=8�D=��C=�\C=e�B=s:B=W�A=2A=�~@=o�?=#?=�U>=9�==��<=Q�;=��:=�:=�I9=��8=��7=js7=��6=�6=XF6=��5=2�5=�M5=.�4=�v4=o�3=u^3=*�2=-2=>k1='�0=0=!v/=��.=�/.=��-=��,=�!,=d+=��*=
�)=;)=�;(=�`'=�w&=Xy%=�_$=K&#=��!=�I =h�=��=%=�3=�F=�V=�g=�|=��=Ϻ=+�=�
=�3=tU=,l=t=/k ==��<�R�<���<Xz�<��<O��<��<9��<�K�<���<�l�<���<t�<���<Ɓ�<��<�ĵ<�<�C�<�	�<�Ť<�l�<v��<la�<���<1܍<���<��<�}~<��t<��k<��b<;�Y<�bQ<�?I<�YA<��9<`�1<�M*<c�"<Õ<�l<�
<�}<���;!�;���;��;ګ�;0R�;���;o;1�K;(;�.;϶�:�c{:���9_Q���v�������Һ��
�3-�\�O�bZs�]���o睻L���*���*�һx�\��� �Xt���l7��^�d#��!�Y�%�!*�:.��[2�x6�_�:��t>�&6B���E�@I�dL�4�N�ޢQ�=T���V�JY���[��^��Z`�"|b�A�d�uf��hh��qj��l�o���q�-�t���w��{��X~�aƀ�@K��k���L��
������zȇ��x��������M������#΋������э�.��bH�����>풼�:���~��O����헼� ��hV��ܑ���ќ�J��_N��ā��̪���ˢ��飼E��;C���� �����a@��>���ׯ�S����h����Ֆ�����w)���5�����D�뫼��f���  �  8O=ɥN=�+N=2�M=M=aL=i�K='K=�ZJ=�I=XI=OzH=��G=�EG=ۥF=� F=�WE=&�D=�D=�dC=��B=�2B=��A=@A=^j@=�?=L?=G<>=�c==Ł<=�;=��:=��9=b9=
d8=��7=�@7=+�6=�q6=�6=��5=]�5=35=��4=�_4=��3=K3=O�2=_2=)g1=D�0=	'0= �/=��.=�S.=;�-=O -=UF,=��+=)�*=L�)=f)=d7(=vU'=�f&=sd%=�H$=#=}�!=, =��=��=^�=�=z=�=�.=LD="b=�=��=��	=0=�4=kN=xX=]Q =zs�<�(�<���<�d�<���<��<�>�<���<���<,�<���<jD�<���<4�<y��<�5�<@ε<sx�<"0�<<�<��<nD�<I˛<!1�<�u�<���<R��<Ƀ<v�}<�&t<G�j<�a<��X<N�P<��H<��@<�9<�p1<��)<�"<i/<�<�	<R5<�1�;���;���;Xm�;LS�;MB�;� �;�q;i�N;�D+;��;i��:�h�:{��97���Z�͑��Ժ@��8.�U!Q���t�Ɖ���՞�7��%û�aԻe�仠�������:�4S�M��N��z��R"�cM&��s*���.�E�2�s�6���:�.�>�!DB��E�G�H�m�K�uN��Q���S��'V���X��?[�ļ]��!`�gb���d�2�f���h���j���l�Lmo�7"r��u��Fx�;�{���~��������f���Z��s��l_�� %��K̈��`���"���o3��*����댼0����&���d��X����|,���^��I��������Ԙ����C��s���ٝ��%���k��/����֢�����/���j������E/��ê�w���C��n��m��������q��o����]������o����x��n=��������  �  �N=�N=�N=,�M=W�L=kTL=��K=b K=ZJ=�I=_ I=�H=��G=�]G=��F=\F=lE=��D=cD=[hC=��B=�+B=�A=�@=R[@=�?=3�>=!*>=`P==)l<=˃;=��:=?�9=V�8=�B8=�7=�7=V�6=zU6=v6=X�5=�r5=N 5=�4=O4=K�3=�<3=k�2=�2=�b1=E�0= .0=�/=�/=j.=��-=�-=�\,=�+=A�*=w�)=x)=�2(=rL'=	Z&=ZU%=�7$=��"=W�!=� =eq=V�=��=h�=O�=l�=i
= =#?=Cg=�=��	=��=�=�9=AE=2? =�Q�<�
�<1��<]T�<���<ߟ�<�O�<��<���<�[�<L��<ev�<��<�X�<JȾ<�C�<oе<qp�<��<�ը<T��<&�<˪�<7�<�O�<�t�<"��<���<sP}<ۤs<�;j<�%a<slX<TP<)H<K=@<��8<1<�)<'�!<��<t�<�y	<Y<,��;���;@��;���;i��;Sӛ;9؊;�Ts;�fP;^�,;p�;(��:}��:5�9몸�g��Ғ��ֺ����/�2R�i�u�%��z���̱�f�û�Iջ"��Ξ����ϻ����N�qW�����_"�ו&�Ƿ*���.���2�#�6���:���>��SB���E�!�H��K�|+N�;�P�:S��U��ZX���Z�\�]��`�`b�)�d���f��h�:�j��7m�H�o��gr�cu�F�x���{��T��S���悼�W��+����������a�����ʑ����������W��� ��T������A���z���������n&���L���i��;���.���0ԙ����]`��˶�����%`������]ᢼ����H������\ݧ��P���檼���Fm���K���*��>��������?��V���ӹ��ֺ�ܲ��)r���!��QϽ��  �  0�N=z�N=�N=V�M= �L=�OL=�K=*�J=�YJ=��I=�#I=U�H=��G=�eG=�F=- F=�rE=��D=�D=riC=�B=9)B=�A=?�@=�U@=�?=�>=�#>=bI==wd<=={;=	�:=��9=K�8='78=t�7=~7=æ6=�K6=�5=P�5=�k5=�5=��4=I4=��3=�73=��2=~�1=:a1=j�0==00='�/=�	/=vq.=��-=� -=d,=�+=��*=��)=�)=91(=I'=[U&=�O%=�1$=v�"=��!=U =�i=��=P�=��=
�=i�=.�=�=O3=D\=ۋ=T�	=��=<=3=�>=9 =TF�<� �<ت�<�N�<���<���<�U�<��<���<�k�<^�<
��<���<fd�<\о<�G�<;е<�l�<��<X̨<�{�<>�<P��<� �<�A�<Re�<�u�<s��<�&}<�ws<j<��`<�<X<�O<'�G<�@<%~8<��0< f)<5�!<E�<�<0e	<�� <<��;���;���;#��;;׬;Y�;�;�s;��P;n-;Qk	;s��:s�:��9ቫ�:���D��Φֺ,��z/�'yR�*=v��S������W��jĻ͛ջ�L�p����@�������u��z�4�|"��&�Y�*�j�.�93�7�;���>��YB���E�ūH��uK�:N�r�P�1S��U��<X���Z�t]���_��^b��d���f�h�h�W	k�UNm�1�o�Ԁr��}u��x��|�_x�Wg������8n������̆�5����u�������+������e���,��)���$��fK���;���F����$���F��`��<x�������Ù����R���������\�����f墼����Q�������觼�\��_󪼙���+|��F\���<��<��Ƶ�uV��T����鹼F캼ǻ�����Y2��b޽��  �  �N=�N=�N=,�M=W�L=kTL=��K=b K=ZJ=�I=_ I=�H=��G=�]G=��F=\F=lE=��D=cD=[hC=��B=�+B=�A=�@=R[@=�?=3�>=!*>=`P==)l<=˃;=��:=?�9=V�8=�B8=�7=�7=V�6=zU6=v6=X�5=�r5=N 5=�4=O4=K�3=�<3=k�2=�2=�b1=E�0= .0=�/=�/=j.=��-=�-=�\,=�+=@�*=w�)=x)=�2(=sL'=Z&=^U%=�7$=��"=f�!=� =�q=�=�=��=��=��=�
=� =�?=h=ߖ=v�	=��=�=;=iF=]@ =T�<@�<W��<]V�<���<s��<$Q�<��<e��<\�<b��<(v�<���<�W�<Ǿ<B�<�ε<�n�<��<eӨ<��<�#�<���< �<N�<)s�<���<f��<yN}<�s<�:j<�%a<mX<�P<H<�?@<ģ8<�1<�)<a�!<��<��<V~	<�<���;ǿ�;C��;��;c��;כ;�ڊ;Ws;?fP;D�,;��;e��:��:i��9|ͬ�ݪ� ���>ֺ����3/�<-R��u��%������ձ��ûxPջI��7����ѽ����YP��X����_`"�x�&�G�*�X�.�G�2�c�6�
�:�&�>��SB���E�4�H���K��+N�C�P�%:S��U��ZX���Z�^�]��`�`b�*�d���f��h�:�j��7m�H�o��gr�cu�F�x���{��T��S���悼�W��+����������a�����ʑ����������W��� ��T������A���z���������n&���L���i��;���.���0ԙ����]`��˶�����%`������]ᢼ����H������\ݧ��P���檼���Fm���K���*��>��������?��V���ӹ��ֺ�ܲ��)r���!��QϽ��  �  8O=ɥN=�+N=2�M=M=aL=i�K='K=�ZJ=�I=XI=OzH=��G=�EG=ۥF=� F=�WE=&�D=�D=�dC=��B=�2B=��A=@A=^j@=�?=L?=G<>=�c==Ł<=�;=��:=��9=b9=
d8=��7=�@7=+�6=�q6=�6=��5=]�5=35=��4=�_4=��3=K3=O�2=_2=(g1=D�0='0=�/=��.=�S.=9�-=M -=SF,=��+=(�*=J�)=e)=d7(=xU'=�f&=|d%=�H$=#=��!=., =�=B�=��=c==� =�/=gE=jc=i�=��=T�	=$=�6=�P=�Z=�S =�w�<3-�<���<�h�<1�<"��<A�<���<i��<L-�<���<�C�<��<]2�<7��<�2�<˵<�t�<3,�<�<8��<"@�<Ǜ<-�<r�<���<Z��<�ƃ<��}<�#t<��j<k�a<��X<ʖP<]�H<|�@<h9<�w1<"�)<""<�7<�<��	<�=<�A�;���;���;y�;�\�;�I�;_%�;��q;��N;�>+;R|;d�:?�:T5�9}ۯ����W��&պ�.��_.�HQ���t�����9瞻H#���ûNoԻH����1���>�|V������V���"��N&��t*�d�.��2���6�_�:�y�>�[DB��E�j�H���K�$uN�Q���S��'V���X��?[�ɼ]��!`�gb���d�4�f���h���j���l�Mmo�7"r��u��Fx�<�{���~��������f���Z��s��l_�� %��K̈��`���"���o3��*����댼0����&���d��X����|,���^��I��������Ԙ����C��s���ٝ��%���k��/����֢�����/���j������E/��ê�w���C��n��m��������q��o����]������o����x��n=��������  �  �+O=�N=VCN=,�M=)M=DrL=�K=�K=�YJ=��I=*I=�^H=�G=uG=x}F=�E=�6E=8�D=��C=�\C=e�B=s:B=W�A=2A=�~@=o�?=#?=�U>=9�==��<=Q�;=��:=�:=�I9=��8=��7=js7=��6=�6=XF6=��5=2�5=�M5=.�4=�v4=o�3=t^3=)�2=,2==k1=&�0=0=v/=��.=�/.=��-=��,=�!,=d+=��*=�)=:)=�;(=�`'=�w&=dy%=�_$=h&#=��!=�I =��=L�=�=o4=�G=�W=�h=~=a�=�={�=P
=�6=cX=>o==w=an =���<Y�<���<��<��<���<�#�<��<�M�<���<(m�<9��<�r�<���<�~�<��<b��<�y�<%>�<��<���<�f�<�<�[�</��<a׍<���<S�<{x~<:�t<��k<��b<��Y<BfQ<�DI<�`A<��9< 2<eX*<�"<�<4y<,
<��<���;{+�;��;�#�;u��;�\�;j��;to;.�K;G�(;�;���:a�z:���9�x��\.�����^Ӻ.�:?-� 
P���s�ԋ������� ���ӻۈ�!�F� ��y����M;��a�&�7�!��%��*�.;.��\2��x6��:��t>�y6B�ɾE�rI��L�R�N���Q�=T���V�)JY���[��^��Z`�%|b�D�d�uf��hh��qj��l�o���q�-�t���w��{��X~�aƀ�@K��l���L��
������zȇ��x��������M������#΋������э�.��bH�����>풼�:���~��O����헼� ��hV��ܑ���ќ�J��_N��ā��̪���ˢ��飼E��;C���� �����a@��>���ׯ�S����h����Ֆ�����w)���5�����D�뫼��f���  �  �JO=F�N=\N=��M=/M=��L=��K=�K=mSJ=�I=�H=�7H=ȎG={�F=�FF=o�E= 	E=�oD=��C=NC=��B=�?B=��A=^+A=|�@=m�?=R7?=�q>='�==��<=�;=?;=�G:=]�9=��8=K=8=��7=�;7=��6= u6=�6=L�5=Vk5=�5=��4=*4=Jq3=��2=�2=�k1=��0=�0=sV/=�.=��-=R-=�,=+�+=�9+=��*=C�)=�)=�<(=�j'=�&=M�%=Ex$=cA#=r�!=�j =��=u=�J=�n=��=��=P�=��=��=(�=N=AA
=�b=�~=~�=Q�=� =��<Z��<��<,��<	�<�}�<���<�r�<���<�x�<���<̓�<��<��</=�<��<q��<Lw�<K�<*�<�<x��<q�<���<W��<d�<jK�<�w�<VY<+�u<�l<G�c<��Z<~kR<�4J<U6B<�a:<F�2<Q�*<#<T<�<gs
<��<�; L�;3o�;'��;-ʪ;��;g�;؂k;M<H;��$;q�;.�:��r:� �9gθ�|��>����Ѻ�@
��#,��N��r���L�XҮ�&]���^ѻ���;�'���������k�D������!�Kw%�a�)��-�
2��16��N:�qU>��7B���E��\I�ٖL�e�O�bjR��U���W��Z��h\���^���`���b���d��Uf��0h�d(j�iOl�8�n��Xq��:t��Jw��tz��}��\�� Ձ��1���m�� ����}���T��D��$���Bc������Ɗ�B���@���駍��ގ��.��������/U������8 ��9G������eÚ����� 2���a��3�������L����Ƣ�nգ��3��ue���Ϩ�-[��s�����������F������K���#��Gp��)�������v���2���wW��2���  �   gO=}�N=�oN=��M=d=M=�L=��K=�K=
FJ=�I=��H=�H=�TG=?�F=�F=9gE=��D=,AD=,�C=�7C=��B=_>B=��A=�6A=��@=�?=�K?="�>=ٽ==��<=�<=�K;=݆:=�9=M#9=��8=h�7=�}7=7=��6=�F6=��5=҅5=t5=��4=|4=�~3=��2=4!2=qe1=��0=��/=Z-/=v.=E�-=6-=�a,=��+=r+=�V*=�)=��(=�6(=+n'=��&=�%=��$=�W#=*"=w� =��=�D=[�=��=��=��=�==�-=uD=H]=w
=я=^�=�=o�=Ԣ =��<U��<E+�<��<���<�X�<���<v�<��<���<w�<4��<Α�<_4�<V�<t��<܄�<;f�<{J�<(�<���<���<�>�<���<��<�_�<���<���<F(�<�v<L�m<��d<\<*�S<�<K<�C<($;<;D3<j+<)�#<�r<�2<��
<�<�C�;�6�;��;P»;��;<r�;Fu�;V2g;D�C;� ;���:z�:]Zh:e �91a����k`���cѺ޵	��g+��M�%�p�
+���뛻J����¾�=~ϻ�߻-��{L���i������g��4���� ��%��`)�V�-���1�6��/:�8P>�rTB��.F�\�I�B>M�QkP��^S��V��X�L
[� ?]��I_��-a���b���d��Pf�lh�5�i��l�rin��q�D�s�Z�v���y���|����<R��.���Xك�T�K�\Ն�9���-a�����"Љ�q����q��ql��:���!ǎ�!������_��s��e򕼪Z��$������@G���}��]���ƞ��֟�۠��֡�VϢ��ͣ��ڤ�+ ���C�������-��̫�{���/���߰�H������׃��,۶���12��5��*"��t ���ؼ��  �  B|O=5 O=zN=��M=�AM=��L=��K=B K=�/J=X_I=�H=��G=JG='aF=�E= E=�D=�
D=7�C=�C=¦B=�3B=]�A=l8A=��@=�@=�V?=�>=��==�==�C<=��;=!�:=E:=Co9=}�8=4E8=��7=�F7=��6=�j6=�6=��5=�'5=��4=�4=��3=��2=J2=+V1=�0="�/=�.=�9.=~-=��,=,=�n+=��*=N%*=W�)=n�(=|((=�h'=͓&=�%=�$=gd#=6"=n� =�=�m=��=�==r<=W=l=Q}=��=��=U�
=m�=��=��=��=*� =�<��<^/�<��<;��<z"�<g�<���<2�<Qk�<@��<�h�<��<(��<���<F`�<uM�<�B�<7�<i �<i��<ᯠ<9M�<ϗ<�:�<ᗎ<9�<�E�<䣀<ex<Ko<�f<�W]<5�T<�EL<�C<L�;<��3<�+<�#<�<>^<H�
<�<�)�;���;�M�;���;b�;���;\A�;�^b;�>;�;O��:嵯:ũ[:i��9�[��:$�յ���Һ�	�@M+�K|M��4p�,���'���N��r3��՛ͻ�kݻ
��Z����J�o�
����69��e�2< �<�$�m2)�}{-�O�1���5�d7:�p>�e�B�!�F�ZmJ��N��^Q��rT��BW��Y�� \��5^��`�!�a��^c���d��pf�Nh���i�&�k��Fn���p�k�s�<dv��Hy�d'|���~��̀����
@���Z��ya���T��o6��A
���Ո�k���Bt���Z��N\���~��Î�\&��⡑��+�������E��^ŗ�/5�����ۛ�����.��j:��}4��� ��L��ꢼ�أ��ڤ�0���,6��.���b������}A��;⮼�|��
��/���?hA���~��ئ��ź����������6����  �  5�O=�O=yN=a�M=u:M=$�L=ҼK=��J=�J=�6I=�_H==�G=9�F=�F=nE=��D=�KD=�C=A]C=��B=��B=�B=��A=�.A=֠@=�@=�V?=�>=��==�#==jg<=��;=� ;=�X:=��9=N9=��8=��7=�{7=��6=��6=�6=ɡ5=�)5=��4=\4=�y3=:�2=z	2=�=1=�k0=K�/=c�.=��-=C6-=�|,=,�+=�&+=*�*=V�)=uU)=f�(=)(=QY'=2�&=��%=Ғ$=�e#=j"=�� =i)=��=��=/(=#_=o�=1�=ʼ=`�=X�=;�=��
=�=��=�=��=ӳ =��<���<��<�p�<"��<x��<�
�<�>�<3��<���<�C�<���<�r�<�4�<�<��<S�<f�<��<��<7ߤ<��<dE�<�җ<=N�<���<�-�<랅<��<B)y<�6p<Vg<��^<��U< <M<�D<]r<<�;4<�,<�#<�<�Z<��
<Z�<q��;�.�;W�;E[�;�_�;D��;��;�U];�9;��;��:LW�:��M:���9�H9��+��V��" Ժ�
���+��M�O%p�L���l���M���ϻ�c�˻Pdۻ�\�����9�һ	���[��`��/����$� /)���-�2�1�H6��j:�|�>���B�?"G� K���N��cR���U�fuX�X[��D]�K=_���`��b���c�HJe�J�f��Gh�gj�Ll�;Qn���p�@js�/ v� �x�߈{��"~��Q��o���֬���ȃ��؄�݅��Ԇ�W����������g��pY��9c��]����Վ��@��ȑ�Fb�����!���6:��M���5&���t������+���緟�����=t��D��������j�\���?������&
��v���������\%������Y��q_��m����A#���I���b���n��r���  �  �O=��N=gnN=��M=;)M=HoL=^�K=�J=��I=�
I=�*H=�RG=~�F=��E=�#E=�D=WD=@�C=@*C=��B=�hB=�B=��A=�A=%�@=(�?=LM?=y�>=��==3==��<=��;=�3;=F�:=��9=/`9=��8=�68=J�7=|7=y�6=86=͡5=�"5=i�4=�	4=�g3=c�2=��1=X1=�E0=�h/=��.=��-=�,=33,=��+=��*=H*=n�)=�&)=��(=}�'=�A'=ew&=�%=M�$=�\#=�"=g� =�6=�=�=�Y=��=��=��= =�=M==��
=x�=0�=��=��=� =�<���<���<B�<�p�<���<��<J��<���<7D�<ݫ�<�5�<���<Ʊ�<"��<���<���<1˰<vج<�Ө<��<}�<�*�<�×<�O�<!֎<�\�<��<�w�<�z<Aq<�lh<%�_<��V</N<�lE<��<<D�4<|4,<*�#<��<�-<��
<��<
�;L�;�5�;��;M��;Ѐ�;�Q};�vX;^�4;�;�I�:}�:�?:B�92)b�Ǚ3�;����J׺:�-��N�g�p�ED��I��ߌ��窺�[ʻ�ٻf�Һ��@G����2��������S�$��P)���-��2��j6�^�:��?�xC��G�<�K���O�fS���V���Y�.\�b^�"B`�n�a�'@c��d���e��g��h��Uj��Nl�ȃn��p��ms���u���x��{��u}�����	��j)��PF��[`���u��=���)�������v��@l��|k�� ~��/�������5m������s����V��$	�� ����A��A����	���9���F���4���	��6Ρ�����Q���'�����X*���]��X������ȉ������t���ޯ��=������y೼^)���n������^鸼;���=���X���  �  �O=P�N=�]N=ҾM=�M=zVL=�K=خJ=��I=G�H=0�G=�G=�IF=>�E=%�D=cLD=��C=�\C=[�B=g�B=�EB=V�A=3|A=,A=z@=��?=�=?=��>=��==�:==^�<=�;=�[;=��:=a.:=��9=�8=5c8=.�7=I77=�6=o 6=8�5=�5=��4=��3=P3=�2=#�1=��0=e0=�;/=/Z.=�-=N�,=��+=�A+=��*=*=�)=B�(=m(=��'=�&'=�_&=�y%=�s$=�M#=�
"=� =�;=�=5$=��=s�=?=-=�@="D=�:=_)=p=4�=��=��=��=�� =���<nh�<���<-�<�0�<UB�<�M�<�_�<��<8��<�$�<���<�a�<>;�<%5�<�F�<�e�<���<���<�<P��<	P�<J�<���<�D�<�ގ<�{�<e�<Ł<��z<
r<�Si<Uz`<�W<?�N<;�E<�9=<��4<64,<U�#<+i<>�<�8
<rK<n5�;�S�;��;���;�	�;i��;�?y;x T;�(0;@u;��:�w�:�1:!1[9Gw��L�<�������ں����.�l�O�Vvq��l��晻�
��J̹� (ɻk$ػ���9�����:�������� ��d�$��)�.��o2���6��+;��?�e�C�EYH���L�ߖP��OT�[�W�h�Z�l7]�a_��-a���b��c�H#e��Mf���g��i�k�j�أl���n�d q���s�2�u��_x�h�z���|�m�Ȥ��Ӽ���ڂ������"���D��/_��p���x��S~��k�������׍��+��#���*9��3铼����og����������6��E�������Kß�h���n���$���֢����\_���J��X��>���?Ш�^-��q��������V�����J�c6���w��6���\���Q��霸�,⹼[��|M���  �  S�O=i�N=�LN=��M=��L=�>L=�pK=�J=u�I=��H=��G=w�F=�F=�WE=��D=5D=��C=�0C=�B=�|B=0'B=-�A=LcA=��@=Ud@=�?=H-?=��>=W�==�===��<=�
<=�x;=T�:=�U:=�9=�"9=b�8=��7=�F7=��6=�6=;�5=%5=0x4=�3=�93=ւ2=(�1=�0=��/=�/=`0.=�Q-=�,=Խ+=+=�o*=��)=#Y)=t�(=	M(=η'=�'=	I&=e%=�`$=s=#=5�!=)� =�<=P�=�6=<�=�=�/=�Y=Pm=�l=.]=�C=n%=/	=j�=��=O�={� =��<�?�< ��<���<���<� �<�<!	�<#�<U[�<��<�D�<���<Gܿ<9߻<P��<�!�<I�<�c�<�h�<hS�<&$�<�ߛ<��<�4�<�ގ<���<tC�<l��<�d{<��r<��i<� a<z,X<�2O<IBF<3l=<�4<7$,<�#<�,<��<@�	<+� <�n�;]u�;��;�j�;y��;�/�;zv;�P;�,;h
; |�:�k�:��&:�;49і��aD�����R޺�B���/��!Q��Xr�i���[ߙ�׻��3���JȻ�׻7������ ����M�����g������$�n�)�	X.�7�2��(7���;�G�?��rD�e�H��)M�@Q�U�`wX��x[�+	^��*`��a� Xc���d�էe���f�$�g��ei�tk�s�l�o��\q���s��v�=Ix��vz�a�|���~�AZ��yl���������焼S���E���h��~���q��������ʌ�����Y���Ӑ��n��>%���땼鴗��r��5��˜�����R$��&�����鿡�!m��>��Yɣ�y���nz������<�����PH����������oE����������:󱼰*��gk��}���L��Vf��Լ��(
���K���  �  OzO=l�N=�?N=ɛM=y�L=�-L=�^K=�J=9�I=��H=O�G=+�F="�E=P6E=�D="�C=Q|C=�C=2�B=�eB=mB=B�A=�QA=3�@={T@=��?=!?=�}>=V�==�===�<=�<=V�;=�:=3n:=��9=�99=ږ8=7�7=�O7=u�6=�6=ъ5=�4=�j4=��3=�)3=�q2=ۧ1=5�0=��/=N�.=�.=�3-=V_,=��+=��*={O*=��)=�=)=�(=m7(=}�'=R�&=�8&=�U%=�R$=-1#=~�!=!� =.;=��=�@=��=�=AI=u=v�=��=�q=�R=�.=b
	=D�=2�=V�= � =ؠ�<u!�<]~�<��<w��<H��<���<��<���<��<�u�<^ �<��<���</��<�Ƿ<���<��<G=�<�D�<`1�<��<pě<�w�<�'�<�ێ<햊<�X�<��<�{<�#s<Jhj<�a<�X<�zO<YtF<�=<K�4<b,<��#<1�<kg<��	<� <���;���;�b�;���;�۠;�9�;a�s;4N;�j*;�;vE�:W��:��:�9�n��&�I����,�ຶ]�� 1���Q�� s�nى�[晻Z���!ٸ���ǻghֻ���B�{� ��q���i�"_���{%���)��.�3��k7�>�;��H@�@�D�g6I���M�ŮQ�O�U�i�X�k�[��^���`�db�y�c���d�� f�Og�)Eh���i�YQk�;6m�6Oo�C�q�)�s��v�Ax��Vz��X|��T~��,��#;��.Z��R���Ä� ���8��g��p�����������a猼X"��&{������l���ON��t��藼ԫ��W���ޜ�i:��g���e���<������"���4A��>𣼦�������夦�'ͧ����]������0���c=���r�����nʱ�y����9��̇���㶼�E��n���� ���M���  �  �`O=��N=3N=��M=E�L=�7L=8cK=kvJ=�uI=�iH=a]G=�[F==oE=��D=��C=YfC=��B=�B=�qB=�>B=�B=��A=�mA=l�@=5u@=�?=�3?=x�>=��==�T==e�<=U<=��;=�m;=8�:=�]:=&�9=�
9=vS8=&�7=��6=�Z6=F�5=I5=��4=k<4=��3=��2=X$2=]@1=�I0=~I/=4J.=�V-=Dx,=�+=u+=��*=�*=)�)='`)=�)='�(=�(=`\'=��&=�%=�a$=�!#=��!=j =�=M�=�=�k=޷=��=w�==�=�=7L=�=��	=*�=W_=6:=&=���<_B�<���<��<��<,D�<���<A��<lz�<�y�<ó�<E0�<$��<f�<��<l�<�Ƴ<��<�N�<0`�<`I�<
�<���<a�<|�<BƎ<P��<'{�<h�<#�|<j-t<Btk<�eb<�Y<G�O<�F<��<<�3<1�*<1]"<��<Pw<��<���;E��;�i�;�!�;H^�;Qp�;���;o�d;>;�#;���:y�:�Y:�0�9񑃸��i�x��ٸ�������G>�'`�������ء�e��G^���λ	Dݻ���)$���`����������{%�}�*�-c/���3���7��+<�u@�a�D�(�I��/N���R�EW��[[���^���a��gd��6f��zg�Ph�'�h��Qi���i���j���k�
Im��)o��Nq���s�0�u��	x�� z���{�D\}���~��K��;?��uY��V�����X��Դ�����z&��j;���D��XR��qw���Ï��A����[Ӕ��і�Aژ��֚�ﰜ��W��ÿ��䠼Rơ�eo��j��T��Z����9��ޤ��������;��C��O���u���.?��$h��w���t��Vr��v���ò��	������/������H���z���  �  �fO=��N=�<N=%�M=��L=�AL=�mK= �J=�I=�uH=�jG=jF=�~E=ԯD=�D=lvC=4C=1�B=g~B=VJB=�B=6�A=xA=�A=�@=�?=�<?=�>=2�==HW==��<=`Q<=��;=�d;=��:=�R:=T�9=�9=bN8=@�7=�6=�^6=��5=�Q5=P�4=�F4=�3=L�2=�.2=/K1=/U0=�U/=�W.=ye-=��,=��+=�+=B�*=5$*=��)=hl)=?)=��(=�(=If'=�&=��%=�j$=�)#=��!=�m =��=��=��=�b=��=J�=�=*�=/�=;F=� =0�	=9�=�d=UA=@=��<�S�<j��<���<���<�Y�<��< ��<��<���<
��<�Q�<��<"�<e9�<���<�߳<0�<]f�<�w�<�`�<
&�<қ<�s�<m�<�Ύ<x��<`v�<�\�<�v|<t<"Fk<+9b<��X<�uO</F<��<<λ3<#�*<�v"<^<'�<��<���;�D�;!��;3w�;뻰;ٛ;A'�;��e;�&?;�:;���:���:��]:f��9w[P��L ��u�M���<������`=��x_�=����{��ݸ���^��s���ϻ��ݻ����t��������A����J���i%���*��?/���3�g�7�^<��J@���D�3UI��N���R�sW�� [���^��a��%d��e�e?g�(h�)�h�Z#i��i��yj�Y�k��m�P o��'q�
us���u���w�4�y��{�?o}�+
��^���T���n��쫃� ���`��t���c���i���,��u2��l>���b�����(-���ޒ�P����������ֺ�������7������à�+���qR���Ң��<������$��ɤ�$���˧���ܧ��0������E�7���f��]|��.����������pȳ����ˑ��U���������nt���  �  �vO=��N=&VN=��M=kM=�^L=׊K=�J=��I=,�H=?�G=n�F=^�E=��D=�1D=��C=?7C=��B=V�B=�kB=�2B=��A=:�A=�$A=@�@=��?=�U?=ۧ>=��==�]==��<=�E<=e�;=I;=[�:=�2:=Г9=��8=�>8=��7=��6=j6=�5=�h5=��4=�b4=��3=J3=
L2=Yi1=ku0=y/=�~.=�-=[�,=��+=�M+=��*=�N*=��)=|�)=/)=/�(=�1(=
�'=�&=E�%=y�$=?#=O�!=�v =[�=�z=}�=�G=ǋ=I�=R�=ٝ=Oo=�4=�=w�	=��=�t=�U=�3=�
�<چ�<���<3��<���<���<^R�<�<��<���<�5�<j��<�m�<�c�<W��<ѷ<�$�<vq�<@��<���<���<�b�<�	�<���<�=�<��<���<�d�<�7�<�|<G�s<P�j<��a<"vX<�O<,�E<a�<<��3<I0+<��"<�g<��<e_	<k <D"�;���;�o�;ϱ;��;R}�;#�h;=B;�b;���:���:��h:��9dxb� ��m�� ��򺦽��n;���]���"𐻊n��5_�����g�ϻPS޻t���j����C���H������8%��B*�V�.��03��]7�s�;���?��ED���H��~M�R�hqV�8uZ���]���`��gc�I?e��f�5{g��h���h�P6i� j�'k���l���n�w�p�s�yu���w��y�
�{���}��f��������߭���ー�,���z��Q����ꈼ� ��K��_������)��9u����ţ������w���w��[j��R;��۝��?��Se��4M����������Y���7f��A裼����e��n��Ϥ������e���̫��$��xe��΍��ģ��統�kӲ����[���Ŷ��=��7���X��%c���  �  ܋O=�O=�yN=��M=�AM=a�L=��K=e�J=��I=l�H=��G=�F=��E=�'E=�{D=h�C=z{C=�!C=��B=՜B=�^B=�B=ټA=LA=��@=�%@=�x?=�>=�>=�d==l�<=�/<=e�;=�;=��:=��9=�b9=��8=�"8=;�7=��6=�w6=x�5=�5=�5=ى4=J�3=�>3=%t2=��1=ߣ0=4�/=j�.=j�-=��,==,=,�+=o	+=m�*=m&*=t�)=�\)=��(=�X(=i�'=��&=��%=��$=^\#=��!=�� =��=�i=��==�U=4v=�{=�h=:D=�=��='�	=آ=ĉ=�q=�S=�N�<��<�<52�<�!�<]��<��<���<�u�<��<	��<�H�<���<��<.�<S>�<���<Ͱ<���<U�<J��<M��<�W�<y�<sm�<���<���<YB�<���<�[{<�r<��i<+�`<A�W<��N<,uE<܎<<��3<�q+<'#<��<��<��	<]� <�Q�;���;���;�e�;�ޞ;䌊;]hm;G;�N";��:8�:E�y:{ :��%8_�չJ,a�Vc���l캇��"�8�t:[�q�}��8��"��:~��EW��Űл�߻^m������Y���u����#����$��)��Y.���2�ؽ6�0�:��3?�"�C�:.H�[�L��?Q�ʃU��lY��\�u�_��?b��!d��e���f��Gg���g���h��bi��j�<l�]�m�O'p�v�r�eu�y�w���y��|��~���_���)���?���@���u������·�P����݉��͊����'���ۍ�[&��ף��ER��`(������
�������J�������ҟ�k���~�����}���-�������>��M��^��pW�������'��������� j��:���D᰼�
���7��s���������-~��ع�+���O���  �  I�O=5!O=˝N=-N=iM=ѭL=�K=��J=��I=I=�H=� G=SGF=�E=��D=�HD=a�C=�mC=�C=g�B=��B=]AB=��A=�sA=��@=�K@=e�?=��>=E!>=�f==;�<=�<=wr;=��:=�I:=M�9=�9=f�8=��7=r7=�6=,�6=�6=9�5=�45=Ӱ4=�4=*f3=7�2=��1=��0=��/=C /=/".=RT-=�,="�+=/b+=��*=�m*= *=�)=R)=�(=d�'=�&=�%=��$=�x#=/"=� =-�=N=��=��=i=�%=�+= ==
�=��=�	=ש=��=ь=�r=W��<��<N]�<t}�<Wx�<�[�<.8�<��<h�<�>�<4��<��<��<@��<g��<��<|��<�.�<�X�<�e�<uL�<��<Ӧ�<�'�<���<��<��<a
�<��<|dz<�q<ڧh<��_<r�V<N�M<��D<�H<<{�3<��+<�#<�`<�<�}
<�<<��;Q6�;�_�;=;�;$�;p�;bs;9$M;Ǒ(;=y;���:�g�:��:���8�p���uT��c����J	���5��X���{������蠻 ر��D»'һ!��_���5���������D!�b����$�?x)��-�~�1��6�H:�	�>���B�_vG�R�K�JP�EeT��&X�;~[� `^�c�`���b��?d�$je�+Of��g�e�g�\�h�%�i��pk��Um�L�o��r�9�t��Zw���y�sc|���~��n��!~������L���5����܅��(�,���Q���1����x��p�������׎�T������:ʓ�ĩ��G����Z����u���𝼜�����࠼񉡼#������<����YǤ��Х��	���k���ꩼlv��� ���|���导�:�������������/L��󕷼%۸�h���5��E���  �  n�O=�5O=ͷN=s)N=υM=��L==�K=%K=�+J=�<I=�RH=�tG=��F=��E=�BE=j�D=_-D=s�C=�^C=
C=$�B='dB=sB=p�A=�A=�g@=}�?=O�>=�(>=�^==��<=��;=!2;=��:=��9=	\9=��8=�B8=5�7=�N7=��6=�6=�#6=ݿ5=�O5=O�4=;44=��3=��2=@�1=�1=&0=�J/=�y.=E�-=�-=,\,=��+=�9+=��*=�<*=��)=�8)=�(=	�'=5'=u	&=��$=��#=p"=� =��=K%=`=}�=ԯ=��=	�=�=�=.�=r�=R�	=j�=T�=�=߆=)��<q;�<��<���<���<���<z��<׺�<���<�
�<ea�<���<�{�<JC�<q/�<v;�<o\�<��<�<l��<p��<�L�<��<vW�<[��<��<4\�<��<�!�<�-y<!(p<\.g<@^<fU<��L<s%D<��;<W�3<v�+<F�#<۱<o<�
<��<�l�;�O�;���;{
�;�R�;�ӏ;R\y;��S;Ǚ/;�V;��:��:�&:��(9FT���gI�Vp�����s��%�3��V��[z��%�����߉����û�Իp�㻻7�� ����|�����������$��8)�Eq-���1�3�5���9��>�UsB���F�s+K��SO��7S�-�V���Y�ż\�'$_�),a�9�b�8d�%Ue��If��4g�8h��ri�q�j�D�l��#o�1�q�Gtt�(Pw�)z���|���.���M#���@���U���a��:a���O���*��_�˳��Nu��`G��g8��7S��ߝ��z������+w��A��n��Ի��tT��b˛����hJ���Q���5������J���K����x���ό��F���Ѧ�7��>���n_����������4��ԯ��G���l����������:.��1T���e���b���M���  �  ��O=�9O=�N=�3N=d�M=c�L=	L=9.K=MJ=�lI=�H=}�G=iG=�SF=v�E=�E=b�D=�D=E�C=�6C=��B=ExB=BB=��A=A=r@=z�?=��>=)!>=�H==2s<=F�;=��:=�2:=��9=n�8=l8=?�7=��7=�7=��6=�u6=a"6=��5=@Y5=��4=�>4=��3=>�2=� 2=�-1=�[0=X�/=�.==.=�k-=X�,=B(,=��+=��*=�r*=_�)=�P)=��(=-�'=	'=x&=�$=��#=�"=cq =�=N�=�=D3=rG=CT=\[=L_=@c=^j=�u=��	=�=��=ћ=��=��<�C�<m��<`��<���<��<�(�<cQ�<���<���<�<�<���<F�<���<D��<ͪ�<�<��<Gͭ<�̩<���<2j�<���<�f�<ޱ�<��<��<�N�<���<�w<�n<$�e<�\<��S<oK<�/C<1);<BN3<��+<��#<;�<*�<��
<�<��;���;L��;Q��;)u�;���;ʲ;#�Z;��6;�X;�M�:ɳ�:G�7:w�_9効&�A�����Yߺ����2�U�U�Z�y��2��?���؟��5GŻ�Tֻ@��g?�����r	����=��\��X �9�$��5)�SQ-�t^1��s5�̞9���=�g+B��mF���J��yN�[R��gU�cX��[�w]�٘_��wa�c�2vd�g�e���f���g�Y@i�4�j� �l���n���q��ut��~w���z���}�?B��4�������_��������!����ȇ��}��1#��Lŉ�$r��?8��W$��>��쇎���������<��딼�����"��_���Q����F��Sw����������[t��)D��9��JĢ������u�����=���%�������f��w&���箼�=���ó�_0��h���ٽ���޸�|幼.Һ�娻��q���  �  �O=+O=%�N=9)N=�M=��L=gL=�3K=�_J=�I=)�H=!H=v_G=ѶF=KF=wE=q�D=aRD=H�C=�VC=J�B=K{B=#B=l�A=�A=�g@=��?=��>=v	>=9%==8@<=#b;=7�:=�9=$9=�8=�8=t�7=�47=N�6=��6=GY6=�6=��5=JN5= �4=�44=O�3=��2=�	2=�E1=B�0=��/=/=�u.=��-=�*-=��,=��+=&>+=��*=��)=GY)=��(=��'=N'=g &=(�$= y#=Q�!=O =�=��=0�=��=��=D�=��=,�==0=�6=�U	=�q=8�=;�=v=[��<i#�<���<���<�<�B�< ��<m��<r4�<���<"�<W��<��<��<F=�<t�<��<�ֱ<�ҭ<�Ʃ<���<p]�<y�<�O�<$��<p��< ��<τ<��<�@v<��l<�c<k�Z<CTR<�J</B<3O:<t�2<�+<wb#<uy<�F<��
<�<��; �;{r�;�ʹ;bH�;@��;?ς;<�a;�=;�;>�:��:�CG:�%�9��{�@�>������]ߺ�����2�	V� ez�Ï��z�����DHǻ��ػk�黙v���#���M�-
�B=�_� ��V%��x)�~-�ւ1��5���9���=�+B��CF��*J�i�M�� Q�(T��V�x|Y�(�[��^�<2`��b���c�Ae���f���g��[i�&�j��l�(o�}�q�E�t���w��7{�-�~��Հ��P������ᄼV�^�������T��[爼�m���������UP���9��S������J��H���� �������.��|���d����=��K{������ڝ�������������ۡ�ݶ��T�����������bѦ�l;���ҩ�ӏ��e���B�����v۲�h�������Z��󎸼,���]����R�����H����  �  8kO=O=�N=N=�iM=�L=��K=1*K=@eJ=r�I=��H=�MH=Q�G=vG=�mF= �E=N*E=�D=��C=1jC=��B=$oB=��A=�wA=7�@=�J@=[�?=3�>=�==��<=�<=�;=^;:=/p9=F�8=�!8=R�7=F97=B�6=��6=�i6=906=��5=��5=h15=a�4=4=�o3=��2=�2=�P1=�0=]�/=�a/=&�.=�'.=͂-=��,=�$,=p+=!�*=�*=�S)=�(=�'=%�&=��%=��$=�U#=�!=i  =tP=�g=�n=ln=l=<m=[u=ֆ=c�=��=��
=B	=�B=�[=�a=R=�V�<x��<�M�<̨�<G �<0_�<���<eC�<��<�F�<���<�6�<���<]�<���<�?�<���<cѱ<嶭<���<#t�<�+�<���<�<�H�<[W�<�P�<
E�<f�~<��t<7k<�b<�3Y<��P<��H<��@<[V9<_�1<'n*<4�"<R�<��<B
<�y<��;C��;���;��;)��;!�;*a�;�`g;��C;��;&��:�:�FS:���9��p�U_?�*�����&��}4��xW�|�GŐ�`ʣ�gȶ��nɻ�oۻ,�����C��=��{���;�=7���!���%�c�)�L�-�Y�1��6��):��S>�MjB��SF���I�RM��YP��S��U�aX��|Z���\��_�9Ga�Bc�%e��f��0h��i��fk�nUm��o�Ar�\Bu��x�� |��}��o��j���r��j����Æ�;����X���舼�_��A͉�uC���ӊ�T���s�����{Ў��4��!���� ��u����啼�,���c��g����Ț�p��A>���x��姟�ZĠ�͡��Ƣ�;��������Υ��
��\u��-��֫�?�����������~���:��4̶�V-��x\���Z��b-��Jݻ�/w������  �  �?O=��N=�pN=3�M=ECM=]�L=Q�K=tK=�`J=��I=I=�|H=~�G=�SG=��F=�F=�dE=��D=�D=�rC=�B=�YB=��A=@SA=V�@=r#@=�k?=p�>=��==*�<=V�;=Y�:=��9=j9=x_8=�7=�F7=��6=8�6=�c6=�36=y6=��5=�r5=�	5=!�4=�3=�M3=��2=8�1=EQ1=�0=b#0=ו/=�/=�n.=N�-=�-=�Y,=*�+=��*=�	*=�D)=�{(=�'=X�&=ô%=�$=Q)#=8�!=��=%=�"==�=�
=�=L=`&=�I=}x=��
=t�=�=�+=�3=�$=���<���<2�<�s�< ��<dg�<��<ϕ�<:7�<B��<tW�<��<�)�<���<�<�d�<���<x��<Ɇ�<_�<r.�<�<�n�<bʗ<`��<���<x߈<���<Q}<2]s<Q�i<7~`<��W<GUO<n`G<��?<�\8<1<<�)<�"<�C<�<��	<�� <
�;K:�;=��;O�;�;
��;8p�;�l;{�H;��$;���:9y�:��[:��9[�p�1�B�8����]废�76��Y�F~����?@��b�����˻��ݻ�:ﻂt��-������c\�m.���"���&���*�X�.��2��6���:��>�G�B���F���I��M�t�O�?FR�@�T�*�V�)[Y���[�2E^�ŭ`���b�� e���f� �h��>j�N�k���m�m8p���r���u�ADy���|��;���������R&���n��+~��:U�������u��@؉��3��)����%��wڋ�����ڍ�h��wt���ב��3��z�������ؖ������X7���s��Z������tg������ӡ��颼������{��aY��.Ĩ�x`���+���������$��F��=嵼/���l鸼`�����3Ȼ�mc��\鼼{m���  �  �O=�N=9IN=ٽM=�M=�lL=ǶK=�K=�WJ=g�I=Y'I=ܝH=|H=��G=��F=�BF=��E=��D=�D= tC=L�B=�BB=��A=�.A=��@=�?=pD?=vt>=ɍ==b�<=�;=y�:=�9=F�8=8=z7=��6=c�6=S_6=�-6=�6= �5=��5=K5=��4=�a4=9�3=�+3=��2=�1=�L1=@�0=5;0=��/=5/=٢.={�-=�F-=S,=ح+=�*=o*=�3)=�_(=��'=z�&=ߊ%=Z$=J�"=�s!=L�=�=+�=��=F�=s�=�=��=��=�=8=t
=��=^�=��=�=�� =:��<�<�<,��<�>�<R��<d�<k�<���<Ј�<C4�<3��<�3�<a��<���<��<�w�<!��<ϖ�<�S�<��<��<���<\#�<w}�<���<W��<�{�<TM�<�P|<[Br<F�h<�I_<X�V<�1N<TF<��><C�7<�J0<��(<�p!<��<q<�<�P <W�;��;�C�;d8�;k�;H��;��;r�o;PLL;��';��;]��:K\a:|��9p}v��G������E麚#��h8�0�[�pG��,=����������?ͻ�߻=^�S� �1O���q��=J�L�=J#�$O'�/7+��!/�+ 3��37��O;�[?��7C���F��J���L��dO��Q�{�S��&V���X��[���]�G`���b��e��g�`�h���j��l�.�n��p��}s���v�g�y�9�}������y���.��O������K��t∼�|��뉼*@���������u��I)������'���c��#���M��9N��������r���r���I���A͙����Qg���ѝ��=��Q���⡼���-���D���g�������ɯ���}��'t��X���0������Kn��Z���}��"���%����F��+Լ�4M��ǽ��  �  ��N=ɞN=:,N=�M=M=tSL=-�K=�J=�OJ=9�I=�1I=�H=�/H=��G=�G=�`F=��E=�D=(D=�rC=H�B=�1B=ݡA=�A=��@=6�?=k'?=AW>=�o==~v<=Ft;=t:=�9=!�8=��7=�J7=��6=�v6=H76=x	6=��5=J�5=�}5=�-5=��4=TE4=�3=�3=�r2=��1=AG1=�0=mH0=J�/='Q/=D�.=.=Nc-=��,=��+=R�*=_ *=
&)=�K(=yj'=y&=�l%=�;$=��"=�S!=�=S�=�=��=��=�=�=�=ƨ=��=�=�M
=L�=9�=��=C�=�� =qk�<;�<���<��<B��<�]�<��<A��<ǹ�<�p�<�<�t�<>��<��<�2�<�~�<Q�<P|�<�,�<{�<a��<\a�<��<"D�<�i�<�`�<}7�<`�<ը{<��q<��g<��^<��U<wM<�E<J1><�6<��/<
{(<{� <� <��<։<���;(l�;��;��;�H�;Oʪ;	e�;mԉ;�q;3�N;�*;8�;���:�Sd:��9&�|���J��&���+����:�9�]��"��J ��񌧻	��jλ��G�򻞒��		�t��_����\��R�#���'�ܩ+��/�$�3�Q�7��;�t�?�O�C�w�F�9J���L�W.O��XQ��tS���U��X�[�Z�dP]�j`�ѯb��e��Ng� Ii�f#k�y�l���n��Iq� �s�& w�bjz�P~��0ɂ�U���E��ma���o��T=��eщ��8��y����Њ�.��I���Wc��TJ��;`������U␼+���c�����ߊ���~���o���o�����zΚ�91��˩��'�������|.��5W��
w�����o᧼�L��ꪼ+���g����Ű�q޲��崼�ƶ��q���ܹ����*껼���8��V�������  �  )�N=V�N=�!N=��M=��L=JL=B�K=[�J=}LJ="�I=�4I=J�H=�8H=�G=�G=�jF=�E=��D=�*D=rC=��B=q+B=��A=6A=Ew@=��?=?=�L>=e==$k<=h;=�f:=�r9=��8=��7=*:7=��6=�g6=i)6=��5=��5=O�5=�r5=�#5=B�4=�:4=�3=�
3=�k2=��1=E1=�0=�L0=j�/=yZ/=��.=�(.=�l-=�,=�+=q�*=F�)=!)=;D(=9a'=�n&=�a%=�0$=��"=�H!=N�=Ͱ=��=��=��=	{=�s=�|=�=�=z�=�@
=>=ܲ=��=��=� =yV�<���<m|�<�
�<-��<�[�<�#�<��<:��<"��<M�<5��<���<��<|:�<��<4�<�q�<h�<ݨ<��<WL�<�՛<�.�<�S�<�I�<��<[�<�m{<�Kq<��g<E?^< yU<�6M<�jE<�=<��6<̖/<mO(<G� <��<��<Gb<���;�0�;���;��;�M�;P�;1��;5"�;�br;>>O;��*;B;l�:{.e:��9$����K�l���P�"Y���:��&^��u��[v���移�|��_�λ��Ỏ=����sK	������Y��S�#���'�K�+�ѻ/���3��7��;���?�ڡC��G�c J�g�L�O��;Q�OS��|U���W��sZ�o2]��_�U�b��$e�"ag�0ei��Fk��%m�@)o��rq�|t�=*w��z��D~�����䂼&���1��4��������\����S������犼�C��>ŋ��w��_���t�����L�8��l��K�������Pt���_��\��xw������A������ ��	������V9���f������@���(����a������xά��Ȯ��ݰ�L�����A嶼摸�t���2$���������X9��B���/���  �  ��N=ɞN=:,N=�M=M=tSL=-�K=�J=�OJ=9�I=�1I=�H=�/H=��G=�G=�`F=��E=�D=(D=�rC=H�B=�1B=ݡA=�A=��@=6�?=k'?=AW>=�o==~v<=Ft;=t:=�9=!�8=��7=�J7=��6=�v6=H76=x	6=��5=J�5=�}5=�-5=��4=TE4=�3=�3=�r2=��1=AG1=�0=mH0=I�/=&Q/=C�.=.=Mc-=��,=��+=Q�*=^ *=
&)=�K(={j'=y&=�l%=�;$=�"=T!=;�=��=[�=�=�=u�=��=��=��=��=�=�N
=��=��=D�=��=D� =�n�<;�<q��<��<���<�_�<F!�<���<���<Wq�<0�<=t�<~��<���<51�<
}�<�<�y�<�)�<��<k��<b^�<�<VA�<�f�<^^�<n5�<���<0�{<��q<��g<��^<W�U<�xM<��E<�4><'�6<��/<J�(<$� <�&<��<�<���;lw�;F%�;�;�P�;�Ъ;j�;�׉;�q;�N;�*;��;ɂ�:d:�_�9~:~���J��V���^�B���+:�Ğ]�w/���,�������%��tλ��3�����	����}�����̐�|�#���'���+���/���3���7�_�;���?�{�C���F�TJ���L�g.O��XQ��tS���U��X�_�Z�gP]�l`�ӯb��e��Ng� Ii�g#k�y�l���n��Iq��s�& w�bjz�P~��0ɂ�U���E��ma���o��T=��eщ��8��y����Њ�.��I���Wc��TJ��;`������U␼+���c�����ߊ���~���o���o�����zΚ�91��˩��'�������|.��5W��
w�����o᧼�L��ꪼ+���g����Ű�q޲��崼�ƶ��q���ܹ����*껼���8��V�������  �  �O=�N=9IN=ٽM=�M=�lL=ǶK=�K=�WJ=g�I=Y'I=ܝH=|H=��G=��F=�BF=��E=��D=�D= tC=L�B=�BB=��A=�.A=��@=�?=pD?=vt>=ɍ==b�<=�;=y�:=�9=F�8=8=z7=��6=c�6=S_6=�-6=�6= �5=��5=K5=��4=�a4=9�3=�+3=��2=�1=�L1=?�0=4;0=��/=5/=ע.=x�-=�F-=P,=խ+=��*=m*=�3)=�_(=��'=��&=�%=�Z$=j�"=t!=��=_�=��=B�=�=k�=4�=0�=o�=k=%:=]v
=4�=�=�=�
=�� =/��<�B�<���<�C�<���<h�<��<���<���<S5�<m��<N3�<��<���<��<�s�<��<���<>N�<$�<A�<���<��<x�<y��<Ț�<�w�<J�<�K|<�>r<r�h<{I_<��V<O5N<YF<�><$�7<�S0<�)<�{!<�<�|<�	</\ </�;��;�U�;H�;�w�;ř;1�;��o;pKL;��';1�;sϺ:J�`:'��9��x�L�G���;�麎V�^�8�y\�w`��.U�������#���Rͻ^�߻�m�� ��T��
����M��}L#��P'��8+��"/�!3�\47�hP;��[?�8C���F��J���L��dO��Q���S��&V�ȇX��[���]�G`� �b��e��g�a�h���j��l�/�n��p��}s���v�g�y�9�}������y���.��O������K��t∼�|��뉼*@���������u��I)������'���c��#���M��9N��������r���r���I���A͙����Qg���ѝ��=��Q���⡼���-���D���g�������ɯ���}��'t��X���0������Kn��Z���}��"���%����F��+Լ�4M��ǽ��  �  �?O=��N=�pN=3�M=ECM=]�L=Q�K=tK=�`J=��I=I=�|H=~�G=�SG=��F=�F=�dE=��D=�D=�rC=�B=�YB=��A=@SA=V�@=r#@=�k?=p�>=��==*�<=V�;=Y�:=��9=j9=x_8=�7=�F7=��6=8�6=�c6=�36=y6=��5=�r5=�	5= �4=�3=�M3=��2=6�1=DQ1=ߵ0=`#0=Օ/=�/=�n.=J�-=�-=�Y,=&�+=��*=�	*=�D)=�{(=�'=b�&=ִ%=2�$=)#={�!=�=�=@#=�=�==l	=J=�(=�L={=��
=�=�=0=/8=�(=g�<���<�<{�<���<$m�<���<���<�9�<���<�W�<2��<�'�<���<��<�_�<���<���<X�<2W�<Z&�<�ڠ<�f�<�<@�<X�<�و<��<�I}<>Xs<��i<~`<��W<�YO<lgG<�?<�g8<�1<��)<?,"<�S<|(<��	<�� <�(�;�V�;ڞ�;p�;ѩ;۩�;dy�;]$l;>�H;�|$;���:z<�:}>[:!g�9�#t�?�C�S���庵J��6���Y��~��'��A`�����ۜ˻1�ݻ�P�e����5�������0a�\2��"�<�&�Ǜ*���.�:�2��6�b�:���>���B�S�F���I��M���O�`FR�Z�T�>�V�8[Y���[�;E^�̭`���b�� e���f��h��>j�P�k���m�n8p���r���u�ADy���|��;���������R&���n��+~��:U�������u��@؉��3��)����%��wڋ�����ڍ�h��wt���ב��3��z�������ؖ������X7���s��Z������tg������ӡ��颼������{��aY��.Ĩ�x`���+���������$��F��=嵼/���l鸼`�����3Ȼ�mc��\鼼{m���  �  8kO=O=�N=N=�iM=�L=��K=1*K=@eJ=r�I=��H=�MH=Q�G=vG=�mF= �E=N*E=�D=��C=1jC=��B=$oB=��A=�wA=7�@=�J@=[�?=3�>=�==��<=�<=�;=^;:=/p9=F�8=�!8=R�7=F97=B�6=��6=�i6=906=��5=��5=g15=a�4=4=�o3=��2=�2=�P1=�0=[�/=�a/=#�.=�'.=ɂ-=��,=�$,=p+=�*=�*=�S)=�(=�'=2�&=��%=��$=�U#=Z�!=�  =Q=�h=�o=�o=�m=Fo=�w=��=��=��=��
=�!	=�G=�`=g=CW=La�<���<*W�<���<V�<<f�<���<H�<H��<�H�<,��<�5�<��<t�<W��<d9�<��<�ȱ<ƭ�<擩<9j�<�!�<쮜<��<@�<xO�<�I�<V?�<��~<��t<�3k<wb<�6Y<��P<��H<��@<�c9<�1<�*<�"</<��<fV
<��<�!�;@��; ��;$��;oͨ;�;jl�;1kg;/�C;�;�`�:��:Q�R:ˑ9Uu���@�2��T�xS��x4���W��\|���񣻿춻��ɻ��ۻ���
���8���������A�<�q�!���%���)�K�-���1��6��*:�YT>��jB�oTF�A�I�GRM��YP��S� �U�yX��|Z���\��_�BGa�Bc�*e���f��0h��i��fk�oUm��o�Ar�\Bu��x�� |��}��o��j���r��j����Æ�;����X���舼�_��A͉�uC���ӊ�T���s�����{Ў��4��!���� ��u����啼�,���c��g����Ț�p��A>���x��姟�ZĠ�͡��Ƣ�;��������Υ��
��\u��-��֫�?�����������~���:��4̶�V-��x\���Z��b-��Jݻ�/w������  �  �O=+O=%�N=9)N=�M=��L=gL=�3K=�_J=�I=)�H=!H=v_G=ѶF=KF=wE=q�D=aRD=H�C=�VC=J�B=K{B=#B=l�A=�A=�g@=��?=��>=v	>=9%==8@<=#b;=7�:=�9=$9=�8=�8=t�7=�47=N�6=��6=FY6=�6=��5=IN5= �4=�44=N�3=��2=�	2=�E1=@�0=��/=	/=�u.=��-=�*-=�,=��+=!>+=��*=�)=EY)=��(=��'=]'=� &=R�$=@y#=��!=�O =��=p�=`�=]�=��=��=��=Y�=�=K=~;=�Z	=w=É=�=�{=ި�<�.�<���<���<�<kJ�<���<���<8�<���<��<$��< �<���<q7�<G��<fڵ<�ͱ<xȭ<<���<RR�<��<WE�<k��<���<Y��<�Ȅ<��<�9v<�l<��c<��Z<�ZR<J<�B<^^:< �2<)+<�w#<��<9]<H�
<)<��;G�;���;�;Ca�;,�;�ۂ;�a;>�=;��;��:�S�:�lF:��9PW��T�?�F����� ��'3�lV���z�Y�&���)<��?mǻ�ػ��^����.��
��U����B��� �WZ%��{)�I�-���1���5���9�Z�=��+B�qDF�+J���M�� Q�K(T�%�V��|Y�=�[��^�I2`��b���c� Ae���f���g��[i�(�j��l�(o�~�q�F�t���w��7{�.�~��Հ��P������ᄼV�^�������T��[爼�m���������UP���9��S������K��H���� �������.��|���d����=��K{������ڝ�������������ۡ�ݶ��T�����������bѦ�l;���ҩ�ӏ��e���B�����v۲�h�������Z��󎸼,���]����R�����H����  �  ��O=�9O=�N=�3N=d�M=c�L=	L=9.K=MJ=�lI=�H=}�G=iG=�SF=v�E=�E=b�D=�D=E�C=�6C=��B=ExB=BB=��A=A=r@=z�?=��>=)!>=�H==2s<=F�;=��:=�2:=��9=n�8=l8=?�7=��7=�7=��6=�u6=a"6=��5=@Y5=��4=�>4=��3=<�2=� 2=�-1=�[0=V�/=�.=9.=�k-=T�,==(,=�+=��*=�r*=[�)=�P)=��(=4�'='=�&=G�$=ċ#="=�q =Ѻ=A�=�=�4=bI=�V=+^=�b=g=�n=vz=�	=~�=i�=��=��=��</O�<���<���<���<�<�/�<�V�<W��<���<�<�<���<*C�<��<8��<[��<B��<U��<�­<e��<��<�^�<��<�[�<Ч�<n��<��<�G�<䊀<�w<e�n<�e<L�\<+�S<�xK<�<C<�8;<f`3<��+<|�#<%�<��<<�/<���;<"�;���;���;���;/��;��;q�Z;��6;�H;7�:�]�:+7:�[9�R��b9C�G>��������2��"V�F1z��b��a����ɳ�smŻ&wֻ���Z������|	������b�.] ���$��8)��S-�G`1�u5��9�l�=�,B�wnF��J�zN��R��gU�0cX�[�#w]��_��wa�'c�9vd�l�e���f���g�\@i�6�j��l���n���q��ut��~w���z� �}�?B��5�������_��������!����ȇ��}��1#��Lŉ�$r��?8��W$��>��쇎���������<��딼�����"��_���Q����F��Sw����������[t��)D��9��JĢ������u�����=���%�������f��w&���箼�=���ó�_0��h���ٽ���޸�|幼.Һ�娻��q���  �  n�O=�5O=ͷN=s)N=υM=��L==�K=%K=�+J=�<I=�RH=�tG=��F=��E=�BE=j�D=_-D=s�C=�^C=
C=$�B='dB=sB=p�A=�A=�g@=}�?=O�>=�(>=�^==��<=��;=!2;=��:=��9=	\9=��8=�B8=4�7=�N7=��6=�6=�#6=ݿ5=�O5=N�4=:44=��3=��2=?�1=�1=}&0=�J/=�y.=B�-=�-='\,=��+=�9+=��*=�<*=��)=�8)=	�(=�'=C'=�	&=��$=�#=�"=�� =��=6&=Ba=��=��=��=��=:�=��=F�=��=@�	=��=ݪ=��=��=���<�F�<���<���<���<���<��<��<Y��<��<�a�<���<#y�<�>�<�)�<B4�<
T�<�z�<���<���<_��<�A�<�ל<M�<���<���<�T�<ò�<��<�&y<�$p<&.g<%C^<nlU<�L<�1D<�;<��3<��+<S�#<��<ą<��
<�<Ֆ�;w�;���;�(�;�k�;��;�uy;�T;�/;�G;�E�:�X�:�0%:��$9ƭ����J�\%��ѝ� ��4��W�F�z�#T��r-��E����û�.Ի�
�yQ� �L�l��|��z��|����$�h;)��s-�Y�1���5���9��>��sB�U�F��+K�TO��7S�[�V���Y��\�<$_�9,a�E�b�"8d�,Ue��If��4g�8h��ri�s�j�E�l��#o�2�q�Gtt�(Pw�)z���|���.���M#���@���U���a��:a���O���*��_�˳��Nu��`G��g8��7S��ߝ��z������+w��A��n��Ի��tT��b˛����hJ���Q���5������J���K����x���ό��F���Ѧ�7��>���n_����������4��ԯ��G���l����������:.��1T���e���b���M���  �  I�O=5!O=˝N=-N=iM=ѭL=�K=��J=��I=I=�H=� G=SGF=�E=��D=�HD=a�C=�mC=�C=g�B=��B=]AB=��A=�sA=��@=�K@=e�?=��>=E!>=�f==;�<=�<=wr;=��:=�I:=M�9=�9=f�8=��7=r7=�6=,�6=�6=9�5=�45=Ұ4=�4=)f3=6�2=��1=�0=��/=@ /=,".=OT-=�,=�+=+b+=��*=�m*= *=��)=P)=�(=j�'='�&=%�%=!�$=�x#=�"=�� =��=�N=��=5�==�'=7.=�"=S=��=��=N�	=��=��=�=x=���<�<�f�<d��<p��<�b�<>�<*#�<� �<�@�<���<��<[��<Q��<%��<���<��<�&�<�O�<�[�<�B�<��<��<J�<呓<��<3~�<��<���<x^z<�q<��h<Z�_<!�V<��M<�D<kV<<&�3<�+<�#<~t<Q&<�
<��<��;qY�;F�;�V�;�#�;~'�;	-s;�.M;?�(;rk;��:��:�#:5��8����C�U����8:级a�D6��Y�<|�䵏����.���f»�Dһ���q��I��d��֙��� &�V����$��z)�"�-� 2��6�I:�ˑ>�@�B��vG���K�RJP�{eT��&X�[~[�`^�v�`���b�@d�,je�1Of��g�i�g�_�h�(�i��pk��Um�L�o��r�9�t��Zw���y�sc|���~��n��"~������L���5����܅��(�,���Q���1����x��p�������׎�T������:ʓ�ĩ��G����Z����u���𝼜�����࠼񉡼#������<����YǤ��Х��	���k���ꩼlv��� ���|���导�:�������������/L��󕷼%۸�h���5��E���  �  ܋O=�O=�yN=��M=�AM=a�L=��K=e�J=��I=l�H=��G=�F=��E=�'E=�{D=h�C=z{C=�!C=��B=՜B=�^B=�B=ټA=LA=��@=�%@=�x?=�>=�>=�d==l�<=�/<=e�;=�;=��:=��9=�b9=��8=�"8=:�7=��6=�w6=w�5=�5=�5=ى4=I�3=�>3=$t2=��1=ޣ0=3�/=h�.=h�-=��,==,=(�+=k	+=i�*=i&*=p�)=�\)=��(=�X(=n�'=��&=��%=��$=�\#=
�!=� =w�=�j=��=(=�V=�w=�}=k=�F=�=��=��	=��=Ѝ=#v=X=NW�<Q��<��<�9�<n(�<'��<���<c��<�x�<v��<[��<�G�<���<T�<���<
9�<k��<ư<q��<t�<0�<+��<�O�<�ݗ<\f�<N��<���<�=�<Z�<�V{<]�r<��i<n�`<�W<��N<?~E<�<<��3<�+<n6#<��<.�<� 
<�<�p�;x��;���;M|�;#�;ך�;�zm;�G;tM";V��:��:�by:��9Ŧ8�@׹�!b��筺��캪6�9�ʂ[��?~��Z���:������<r���л��߻3��	��Ѻ�+���z����^��6�$��)��[.��2�ݾ6���:�Y4?���C��.H���L�5@Q���U�mY�.�\���_��?b��!d�
�e�Ƌf��Gg���g���h��bi��j�>l�^�m�P'p�v�r�eu�y�w���y��|��~���_���)���@���@���u������·�P����݉��͊����'���ۍ�[&��ף��ER��`(������
�������J�������ҟ�k���~�����}���-�������>��M��^��pW�������'��������� j��:���D᰼�
���7��s���������-~��ع�+���O���  �  �vO=��N=&VN=��M=kM=�^L=׊K=�J=��I=,�H=?�G=n�F=^�E=��D=�1D=��C=?7C=��B=V�B=�kB=�2B=��A=:�A=�$A=@�@=��?=�U?=ۧ>=��==�]==��<=�E<=e�;=I;=[�:=�2:=Г9=��8=�>8=��7=��6=j6=�5=�h5=��4=�b4=��3=I3=
L2=Yi1=ju0=y/=�~.=��-=Y�,=��+=�M+=��*=�N*=��)=z�)=/)=.�(=�1(=�'=�&=S�%=��$='?#=�!=4w =��=R{=�=xH=��=v�=��=|�=/q=7=e�=�	=[�=�w=�X=�6=��<���<��<^��<k��<���<�U�<��<���<���<�5�<ɱ�<zl�<�a�<L��<Gͷ<] �<�l�<���<g��<͙�<�\�<Q�<E��<�8�<ߎ<���<oa�<L5�</	|<x�s<4�j<2�a<iyX<�#O<��E</�<<��3<Y:+<~�"<'s<W
<"k	<�v <'8�;ϳ�;���;�ޱ;��;2��;B�h;5CB;�a;���:�ײ:wh:"8�9�+��U𹳸m��~���}����;���]����������t��'�����ϻ�b޻���Av�����`#�������:%��C*���.��13�h^7��;��?�FD���H�M�>R��qV�PuZ���]��`��gc�R?e��f�9{g�h���h�R6i�!j�'k���l���n�x�p�s�yu���w��y�
�{���}��f��������߭���ー�,���z��R����ꈼ� ��K��_������)��9u����ţ������w���w��[j��R;��۝��?��Se��4M����������Y���7f��A裼����e��n��Ϥ������e���̫��$��xe��΍��ģ��統�kӲ����[���Ŷ��=��7���X��%c���  �  �fO=��N=�<N=%�M=��L=�AL=�mK= �J=�I=�uH=�jG=jF=�~E=ԯD=�D=lvC=4C=1�B=g~B=VJB=�B=6�A=xA=�A=�@=�?=�<?=�>=2�==HW==��<=`Q<=��;=�d;=��:=�R:=T�9=�9=bN8=@�7=�6=�^6=��5=�Q5=P�4=�F4=�3=K�2=�.2=/K1=/U0=�U/=�W.=xe-=��,=��+=�+=@�*=4$*=��)=gl)==)=��(=�(=Kf'=��&=��%=�j$=�)#=�!=�m =��=ԃ="�=�b=7�=��=��=�=(�=SG=0=��	=��=Af=�B=�=��<�V�<H��<5��<��<�[�<��<���<��<��<(��<vQ�<��<�
�<�7�<Ʉ�<�ݳ<�-�<�c�<�t�<�]�<#�<+ϛ<�p�<��<|̎<n��<�t�<V[�<�t|<t<Fk<�9b<L�X<wxO<�	F<�<<z�3<X+<�|"<G<8�<��<� <5P�;���;���;İ;�ߛ;^,�;��e;*?;;:;���:Q�:�t]:&�9*�T��� ���u��}��.p��*��={=���_� ΀�����ġ�|i���|��� ϻ|�ݻ����z��6������\��y���j%�f�*�F@/�6�3���7��<�#K@��D�VUI��N���R��W�� [���^��a��%d��e�h?g�*h�+�h�\#i��i��yj�Y�k��m�P o��'q�us���u���w�4�y��{�?o}�+
��^���T���n��쫃� ���`��t���c���i���,��u2��l>���b�����(-���ޒ�P����������ֺ�������7������à�+���qR���Ң��<������$��ɤ�$���˧���ܧ��0������E�7���f��]|��.����������pȳ����ˑ��U���������nt���  �  J�N=�hN=�M=peM=�L=&L=�SK=W\J=hEI=�H=�F=�E=R�D=��C=3#C=g�B=;PB=)$B=B=OB=��A=s�A=tA=�A=�l@=8�?=�?=�M>=ި====f�<=h[<=P<=r�;=dI;=y�:=�:=�R9=C�8=��7=Q�6=�J6=��5=�O5='�4=�y4=8�3=yV3=:�2=d�1=B�0=�/=�c.=�U-=we,=Ɯ+=� +=e�*=H*=r*=��)=��)=2�)=)=.w(=��'=�&=Ak%=�$=_�"=�`!=s =/�=<=��=�=�==C1=�=�=�=��=m3
=��=�=��=�q=E��<�*�<�r�<�m�<��<��<���<uH�<���<|�<��<���<���<��<P�<�ٶ<)i�<w�<,�<�;�<��<���<{4�<^��<�S�<��<a�<�.�<�X�<��|<:�t<��k<�b<]�X<��N<��D<;�:<�r1<�(<�	 </�<(�<�e<�?�;&��;��;M{�;~��;�L�;(S~;�^S;��*;o�;>�:���:�:���8.����;�X����1Ӻ�	�8�+�>�N�C�r�R���1���]��������ɻw�׻[�����b��	����%�������&�Ò,���1��56��0:�L�=���A�Q�E��J��N�?�S�K�X��r]�e�a���e���h�g k�e�l�i=m�X]m��,m�9�l�&�l��Lm��=n���o�E�q��5t���v�� y�&8{�4�|�{'~��,�;��u���􈁼�������}��K��`���t#���^���f��L���)������G�������t���w��W�������B���]��42������QƢ�‣��꣼k��6���X��墤�`+������w��w��E����w���ᬼK�� ��/񯼕���!m��.S��~r��}Ӵ�Ho��02����������B���  �  SO=�xN=�M=�wM=��L=s6L=wcK=�kJ=~UI=-+H=��F=��E=��D=*�C=�:C=��B=ofB=�8B=l"B=:B=��A=��A=��A=hA=z~@=��?=�?=&]>=�==�&==g�<=OY<=�<=b�;=$=;=˲:=�
:=vJ9=}8=v�7=$�6=�T6=��5=e`5=i�4=�4=K	4=�f3=͞2=�1=��0=��/=Nw.=Xk-=,|,=/�+=^+='�*=�]*=�,*=�*=��)=��)=%)=��(=E�'=(�&=�|%=.$=��"=�j!=p =��=�6=�==�.=�"=R�=��=�=i�=F8
=��=Ź=��=m�='��<�G�<���< ��<m;�<��<�<xo�<���<���<���<�(�<���<6�<y�<���<��<\�<4O�<`�<�4�<|ן<�[�<ܖ<q�<�.�<�<�.�<�N�<.�|<�t<��k<��b<��X<'�N<o�D<��:<��1<��(<�A < <=�<T�<O��;���;��;���;��;��;�;'�T;f,;�";�+�:�Ņ:�l:� 9{���/7����к���h*���M�(�q�����V�������b���ɻ�׻���U�����J2	�p��u�����F&��f,�H�1���5�6�9�դ=�lA��mE���I��nN�WS�QX��#]�S�a�)ke���h��j��1l���l�Bm�0�l��l�&�l��m���m���o�_�q���s�Auv���x�l{���|�M"~�T;�'��Pˀ�4���ݷ���
��ڋ���!���������6G��5H��)��N��c���<&������qU���W��Ō��#ؙ�����1�� ���}������S������C���g��h8��������ޥ������R���Щ��V��Ǭ� 
����������@���j�� ���?봼����=��x�������0���  �  d)O=ȤN=�(N=�M=dM=cL=3�K=8�J=y�I=�ZH=�0G=WF=^E=d0D=CC=�B=�B=�qB=�UB=�BB=8)B=9�A=�A=v?A=ƭ@=@=�D?=��>=��==3<==e�<=�Q<=�;=��;=p;=�:=��9=�09=wo8=��7=97=�q6=�5=��5=�)5=�4=R74=l�3=!�2=��1=��0=��/=ͭ.=v�-=�,=��+=.\+=�*=�*=�c*=�7*=D*=(�)=N)=��(=)�'=��&=��%=WY$=��"=��!== =�=#&=�=��=�=�=�=�k=�=ם=F
=�=��=I�=ͬ=��<���<��<u��<ۋ�<��<�t�<���<`i�<�/�<�E�<$��<Nz�<ݒ�<�<�f�<��<�`�<٫�<࿨<嘤<J>�<���<�9�<Ⱦ�<�d�<	5�<�(�<�+�<QF|<��s<$k<��a<�LX<wN<_�D<�
;<��1<�,)<J� <&�<�<�R<Q�;VA�;xM�;�P�;ߗ�;n��;��;��X;��0;W�
;�:�7�::$:JI9Kvp�Z�*�������ʺ�Z�"'�'YJ��Pn���5���}K�����1ʻg�ػ��滻l���"�6�	�yN���L���>&�K�+���0�Y65�V!9�u�<�ް@���D��I��M�A�R���W�#H\��`�Qfd�pg���i��+k���k��0l��l�E�k���k�Fel��Nm�l�n���p��*s���u�\Fx���z�(�|��~��k��W�����~큼���I�������3��Ӣ��<퉼A����ˌ�N���e����ˏ�BA��� �����D0��Fr�����������������w���Ӣ�~J����������ߣ��.��ܶ��z�������#��p�������|��b֭����������ְ�Ƕ��򰲼	س��2������aa��9
��!��������  �  2ZO=a�N=�iN=��M=�RM=��L=}�K=��J=ҽI=&�H=N}G=^iF==oE=/�D=�C=�bC=�C=v�B=n�B=m�B=wdB=�3B=��A=�zA=��@=B@=�?=v�>=^>=�W==;�<=$A<=-�;=X;=��:=bM:=9�9=_9=nU8=��7=x7=ח6=$,6=��5=�j5=��4=<t4=��3="3=	2=�1=�0=��.=�.=5 -=u`,=��+=�L+=��*=��*=�}*=�B*=6�)=�)=h�(=�(= '=��%=S�$=%#=��!=�" =��=k=�b=t�=^�=�=M�=<=��=>�=�V
=�)=l=��=��=&��<��<YC�<=�<��<o��<��<��<Q$�<��<s�<��<�D�<rK�<���<���<rq�<\ݰ<�&�<�>�<��<Ƞ<nJ�<g��<�'�<ɫ�<�P�<q�<��<w|{<��r<rj<z�`<moW<~�M<dYD<�;<�C2<��)<ڵ!<��<Ɲ<�9	<_ <���;��;�/�;��;��;���;�B_;�W7;��;��:�	�:�M;:-�9#:&�V���|��_�º�%�r�"���E���i�)��	���^H���º�uvʻ�ٻot�G����b�
����
!�t����%��P+�0��84�m8���;�L�?��C��3H���L�=�Q�KoV��[�w6_�Z�b���e��
h���i�΃j�n�j�0 k���j��k���k�ril���m�w�o�1&r���t��lw���y��4|�� ~����<����~��l���~��򵄼����Y��K���z�������A����K���!�����T���ϐ�r����������tߘ�������ǳ���!���?���������*���e������wF�����(!���p��C屮턪�"��ّ���⮼�	��������(���W��������������!��N���U����  �  �O=�O=��N=�(N=��M=��L=��K=-K=��I=�H=��G=��F=��E=�E=ZlD=��C=�wC=#+C=f�B=w�B=i�B=kB=B=�A=�)A=s�@=��?=�>=�0>=�o==�<=�"<=��;=�;=�:=��9=�]9=0�8=]+8=��7=�#7=��6=�`6=�	6=m�5=�:5=�4=4=q73=�P2=�W1=W0=�Z/=�n.=*�-=�,=�F,=��+=�b+=�+=��*=�*=b,*=��)=�)=O(=Q'=+#&=��$=WT#=a�!=P* =��=,�=>=[G=iY=�N=J+=��=F�=Ї=�`
=sI=�<=�1=�=[��<�g�<���<*��<Gg�<�<��<�E�<p�<���<?'�<���<_=�<�)�<�N�<؜�<,��<#\�<��<Ѻ�<ᠥ<cQ�<PԜ<8�<���<�<^�<��<6��<Yz<<�q<��h<�u_<V4V<j�L<�C<5	;<��2<�t*<��"<l�<��<�
<�/<���;&��;�$�;?�;�ݜ;;�;wg;��?;�`;��:�ª:� W:.(�9,�����mi|�����f���dW�LA�Rqe�5���j��p\������D˻�5ۻ�������o������� ��j	 ��%�ʸ*��-/�~93�(7���:�)�>���B�.UG���K���P��2U�ǌY��~]���`���c���e�1�g���h�#mi���i���i�-,j��j�t�k���l���n�7#q���s� �v��[y��{�O~��3��+���������-���O���y��c���ʦ��J���Z��d��͋������#Ꮌ�b��>"������#���8���;��������:���=�� ��ơ��;��ɓ��S梼�K���٣�:���������n��(��+���XS��}ծ��3��Hs�������ϳ��	��nU��ҭ��s���Q���}�������  �  x�O=|HO=D�N=�WN=I�M=��L=�"L=F1K=�0J=),I=�-H=�>G=veF=~�E=��D=xkD=��C=ȓC=�HC=�C=��B=��B=�CB=@�A=rUA=�@=��?=�%?=qN>=�x==I�<=��;=JI;=ȫ:=�:=0�9=��8=,m8=�7=,�7=�!7=D�6=��6=-86=��5=0h5=��4=�(4=�]3=v}2=W�1=�0=��/=�.=V.=�o-=��,=�L,=;�+=�q+=x+=U�*=uW*=W�)=�<)=s(=�x'=4M&=�$=t#=��!=�! =(`=��=��=*�=H�=��=��=ț=�|='f=�Z
=VY=�Z=�V=UC== =ۥ�<���<���<���<!��<@�<S�<)��<��<AK�<��<EJ�<��<��<�7�<�x�<��<~��<��<��<���<�>�<<��<�ړ<��<�M�<��<���<�x<��o<w�f<�]<@�T<g�K<�C<��:<h�2<��*<(#<�=<�$<��
<�<���;/�;m��;�@�;���;�z�;�ko;I;��#;P+ ;��:I^t:Z)�9��޶4���$o��`����q��f�=���a�l���~B��kߨ�����̻zlݻ^��46��N$��a��@����z �a�%�?X*���.�#v2��C6��:��>�OPB�޴F��4K�K�O�~T�?X���[���^��a���c�I�e���f�2�g���h��i�%ti�fj���j�	Kl�	n��bp�os���u�B�x���{�
�~�襀�ҁ��낼����*��������m���Ј�:���4"��㾊�wm��mA��tJ���������ґ�R���̦��Ė��o��v!��n���w���1$��-��4砼
���l���z����������\T���U�����n������ o��1��&殼�~��[���W��R����뵼O-���g������#��������h���  �  ϴO=[O=#�N=�iN=H�M=9M=P.L=�CK={QJ=�`I=a{H=��G=m�F=Z/F=ˊE=�D=6lD=|�C=��C=�;C=��B=�B=�NB=e�A=vdA=5�@=�	@=�6?=�T>=�l==�<=��;=��:=8:=�9=� 9={8=�8=r�7=,N7=!7=8�6=ړ6=*L6=�5=2y5=^�4=D34=k3=��2=ö1=��0=�0=�P/=W�.= �-=�a-=��,=HG,=3�+=�S+=��*=Tl*=��)=C)=7z(=��'=�Z&=� %=z#=��!= =�&=�<=�I=�O=kM=�D=m8=�-=+*=B0=-?
=RQ=_=�_=<L=� =���<���<���<W��<��<-��<���<���<V �<Yn�<��<�R�< ��<n��<���<�͵<n��<�"�<?9�<*�<T�<�q�<Ș<���<�	�<�<O(�<sN�<�w<�m<�d<!�[<J�R<4J<��A<O:<�e2<��*<�=#<�q<cS<��
<=�<���;���;���;m��;6F�; �;W�w;IKR;0�-;�m	;�[�:
�:�|:|Z8�e۹�g�mp��W��V�"�;�]`�Զ���ԕ����:���{λ�3�k񻁏 ��#�@�H��;���6!��&�DQ*�<L.��2�]�5���9���=��B�zF���J�O��S�{�V��Y��\��N_�g�a��|c��&e�b�f��g��^h�	i�|�i���j�l���m�p��r��u�a�x�9C|�Px��<������ރ����~��� ���և������!���������E����C��$��[+���z��������}���K��w��6����4��ۗ��ߜ����G������堼�����5��΢��u��V?���:��q���㧼=����Y���;�����Vﰼ����n1��h������*���F���A��-��ӻ��w���  �  ͢O=�OO=a�N=�[N=��M=T�L=L=;;K=ZJ=��I=�H=�G=�RG=��F=pF=�pE=8�D=�HD=k�C=eVC=��B=��B=[;B=��A=�RA=�@=B�?=�*?=N@>=CI==-P<=�_;=��:=5�9=�9=Ir8=q�7=��7=�B7=n
7=��6=�6=��6=�A6=X�5=Pi5=w�4=q4=[3=ȏ2={�1=Q1=V0=�/=B/=d}.=R�-=�F-=e�,=a,= +=��*=^g*=�)=I*)=a(=m'=NH&=�$=�c#=��!=&�=
�=��=�=��=Z�=r�=R�=��=��=��=�
=;/=WF=HJ=�4=� =�o�<{��< ��<<��<���<d%�<1g�<���< �<�z�<9��<�B�<��<0O�<Y�<�<���<��<��<��<&ס<Te�<0��<vؓ<XЎ<N��<��<3<	u<Q�k<�9b<XDY<��P<	xH<l�@<�9<-�1<k*<��"<�(<l <�j
<�n<�A�;�>�;��;-�;�O�;�ؑ;�/;��Z; g6;��;�n�:��:��:SW�8��ҹQg�*N�����=��g<�o`�^؂��=��H���W�����л�h�2���ӱ��P
��M����A?��9"��&��*��}.�2<2�e6�t:�@)>��kB�`�F�Z�J���N�obR�B�U�dX���Z��D]�:}_�r�a���c��We�Z�f�h�8i��j�Qk�Ljl��n�SAp���r��u�[y� �|��=��9����1脼 ���(��g��7����5��{����뉼xD������X���3���M��ݣ��7)��Z̑�y�����W�������a��젚�؛�����9��D[��e���P�����>ܢ�����$i���`����������]���l{��]w��ۀ��<����g���$��ղ������?��r>�����᲻�2:�������  �  yO=�)O=��N=�0N=��M=�L=��K=�K=�LJ=��I=��H=FH=�G=-G=+F=�E=�1E=��D=+�C=(]C=��B=�tB=�B=S�A=z$A=*�@=��?=b?=�>=�==�<=;=�:=�59=�{8=�7==l7=�7=��6=��6=W�6=9�6=�\6=�6=[�5=�<5=��4=��3=�13=�t2="�1=�1=�0=� 0=�y/=��.=,R.=��-=@�,=6G,=ߖ+=�*=�K*=��)=�(=g,(=E;'=�&=J�$=�4#=�t!=.�=^�=9i=�H=�+=�=b==t3=�]=h�=��	=��==
=;=���<|��<�A�<Au�<7��<!��<�`�<@��<8j�<f��<ra�<
��<�<`Y�<h��<�:�</�<dʱ<3ƭ<Oʩ<콥<���<X�<�s�<���<�m�</�<��<%Q}<�s<Ei<�_<��V<��N<Q�F<&?<��7<��0<�)<b9"<�r<>><e�	<� <���;�4�;;��;o��;(¥;�<�;E��;* b;7>;�E;��:�Ɲ:��):�]�8+^չAm�Ғ��ސ����$>���a�Jσ�Od���z�������ӻ���
�������yb�"w�f���m#�ӑ'��b+��/���2�1�6���:�^�>��#C�sRG�/FK� �N��R���T��#W��ZY���[��]��`��Ib�?yd�Upf��h�h~i�Z�j��k�S*m���n���p�|s��v��z���}�<ـ�����q�������<��SD��P����|�+��G\��$�����뤋�J������s������������v��rd��2������dϙ�	����0���y���Ǟ��	���0���4�����,bɤ�����:妼@H���nͫ��ۭ�A��+��t;������Ƿ�0���V���;���廼Z`����� ���  �  AO=w�N=�N=w�M=�EM=��L=ӴK=��J=?1J=i�I=s�H=�yH=b�G=�pG=B�F=T.F=7vE=�D=��C=�TC=\�B=�BB=��A=�`A=�@=�R@=C�?=�>=��==M�<=׼;=�:=�9=P�8=@�7=�_7=��6=�6=�{6=h6=?\6=zJ6=�%6= �5=��5=��4=�_4=^�3=��2=KK2=B�1=,$1=W�0=�;0=��/=�B/=��.=��-=�7-=�k,=&�+=%�*=	"*=9n)=ڴ(=��'=a�&=n�%={�$=!�"=h2!=^?=�)=��=m�=W�=��=�=ɔ={�=��=�:=�}	=��=��=E�=a�=4�<�p�<��<��<z_�<���<@}�<5�<���<���<��<7r�<��<���<���<�G�<�ŵ<�{�<z]�<�T�<G�<�<���</�<q�<��<���<�6�<A�{<:q<�5g<�]<�T<V�L< �D<V�=<|�6<Ƽ/<��(<�G!<�{<:<̍<�(�;N��;/��;��;��;߫�;��;5�;��g;�'D;$;b��: �:�A1:��8�@�~Bw���������_y�.bA�	e��P��� ��nV��9����Tֻ�M���c��Ƃ��M�<3��F ��$�w�(��H,���/��3��7��;�d�?�D��,H���K�)O�.�Q��0T�4V�;"X�K&Z��Z\���^�9Ra���c��Gf��_h��j�X�k���l��,n���o���q�@Wt��nw�� {���~��z��Jx���P��vzB��/H�������p������fƊ�ߊ�U���q�����J����'��⅏�� ���~��m瓼�*���C��>>���.��I+��6E��K���C圼�Z��pП�I/��g��$t��Wc��uI���?��_��׹���Y���<���V�������ֲ�������7Ƹ��6���V���'��R���]���R�������  �  tO=�N=GJN= �M=�M=KAL=�yK=��J=J=��I=\	I=��H=�+H=a�G=G=tiF=S�E=M�D=�D=XFC=�B=�B=�A=�A=��@= @=(g?=�>=͢==�<=x;=�Z:=QL9=�Z8=��7=Q�6=;�6=�G6=�(6=6=6=�6=��5=	�5=�F5=��4=�4=�o3=��2=; 2=�1=�!1=O�0=qc0=#�/=�/=+�.=1.=�`-=�,=W�+=��*=�)= 5)=gs(=u�'="�&=��%=�G$=�"=�� =��=��=�= l=�8=n=n=�)=�Z=��=r�
=�8	=et=)�=^�=�|=D��<q��<�7�<���<�<��<>��<j�<J�<8�<֚�<g��<@�<�<�"�<B�<	��<�'�<N�<Eܨ<�ˤ<}��<�B�<���<v��<?}�<��<��<Rz<�o<��e<?\<�0S<�	K<l~C<�e<<�5<A�.<�'<U <��<4<g�<��;w�;�;�;��;�N�;�*�;�.�;��;�l;��H;5#;k��:���:XM5:!��8�������úDd��#�6�D�
[h�rG���2%��5�û�ػ���r���Im��!�������׊!���%���)�~+-�|�0�9y4�,m8�&�<�5�@�E��	I�H�L��O���Q��S��U� FW�e*Y�b][�	�]���`���c�zEf���h�þj�fl���m�p1o�o�p�^�r��;u�\Ox��{�����
�����@	��1���]�����iƊ��$���I���Q��[�����⋼)����v���������{��}璼�1���L���8������ӗ�����ř�3	��v}��?�������=��Ƞ���У��פ��ɥ�¦��ܧ�O0���ʪ������ͮ�����l��(���oƷ�+���O
���%��m輼8a������vؽ�����  �  &�N=K�N=�N=*�M=I�L=�L=NK=*�J=��I=GyI=�I=(�H=IH=c�G=>G=]�F=��E=�D={D=�9C=�B=��A=BgA=��@=]t@=��?=�:?=fk>=Yx==�h<=�G;=%:=�9=�8=N7=�6=JG6=

6=}�5=y�5=��5=��5=r�5=��5=-5=��4=�3=&A3=�2=L 2=�1=T1=�0=�y0=�0=
�/=R/=}Q.=�w-=��,=��+=R�*=>�)=)=cC(=q'= �&=�i%=L$=c�"=B� =]�=X�=k=S*=��=}�=��=F�=%=�d=#�
=�	=�E=
i=�j=*K=[�<��<���<�B�<��<(��<u��<@��<�~�<)Q�<���<~>�<�X�<YK�<'5�<\7�<n�<�<�<i��<bn�<�E�<�<�I�<r[�<�%�<]��<C4�<Kfy<��n<�wd<��Z<�R<� J<��B<��;<|�4<��-<W '<��<c�<�q<:�<��;���;#�;=<�;��;�d�;�ؗ;q�;s�n;1.K;��%;<��:�&�:%7:�6�8q���3��N�Ⱥ�)���%���G���j��/��o훻�z��tŻ�Tڻ�� ��w	��.�B��@��og"��&��I*�p�-�Rd1��"5�%9�(R=�#�A�z�E�ɬI��M��O�v�Q�B�S��7U�>�V���X���Z�F`]��J`�Yc��Pf��h��8k�m�3�n��o�r�q��rs���u�w�x���|��N���n���������Y;��ܝ�������G����������ڳ������;؋��6��ߌ�Ӎ�5��ph���֑��4���i��Zi��S8��B떼����wr��z��<��� A��M라(���,M���̢�����-���(��#���:��.���� �����$��rt��mԳ�3$��$D�����[�������%g���ս�w��I7��_j���  �  ��N=��N=N=�uM=
�L=��K=>K=U�J=��I=guI=�I=�H=�RH=]�G=�JG=�F=n�E=�D=�D=�4C=�yB=I�A=�VA=v�@=5b@=f�?=�*?=�[>=�h==NX<=86;=�:=��8=8=�67=]�6=:06=�5=i�5=]�5=@�5=�5=�5=�p5=d5=~4=��3=�/3=��2=��1=�z1=%1=��0=�0=U'0=j�/=�/= \.=y-=�,=��+=W�*=��)=��(=�1(= ^'=rp&=�W%=P$=�{"=V� =��=�=�U=7=i�=��=�=R�=�=3P=��
=[�=�5=�X=GZ=�9=���<�Z�<���<z&�<���<>��<��<���<W��<�h�<4�<�W�<Om�<Y�<�9�<�1�<6^�<�ϰ<Ѐ�<�]�<�I�<f"�<Kɛ<�)�<g;�<��<��<��<�y<nQn<^d<��Z<8�Q<ģI<�3B<:;<�{4<��-<��&<�`<��<�,<~r<	�;a2�;_��;���;���;�w�;��;BI�;�do;LL;}z&;�:-�:�`7:4��8�3��NɆ��ʺ�C�F'��H���k�F���<j��������Ż��ڻ�6�$#�j�	���<�q���"���&�|�*��.�Y�1�Ja5�-a9���=�f�A�PF�[�I�j:M�-�O��R�4�S�(U��V��bX�)�Z��4]��+`�<Kc�Wf��i��ek��Bm��n�C<p�!�q���s�*v��6y���|��o������ǲ�����Fi���̉��Њ�iu��eǋ�u݋��֋�[Ջ�����V�����L���`,��판�*����P��f~��qt��89��f▼�����[���`��駚�2-���ޝ������S��@ݢ�q.��M��EL���G��&^��T���W@��!���D��k���y���6M���p���G��x»�Wڼ�铽������5���Y��t����  �  &�N=K�N=�N=*�M=I�L=�L=NK=*�J=��I=GyI=�I=(�H=IH=c�G=>G=]�F=��E=�D={D=�9C=�B=��A=BgA=��@=]t@=��?=�:?=fk>=Yx==�h<=�G;=%:=�9=�8=N7=�6=JG6=

6=|�5=y�5=��5=��5=r�5=��5=-5=��4=�3=&A3=�2=L 2=�1=S1=�0=�y0=�0=	�/=Q/={Q.=�w-=��,=��+=P�*==�)=
)=dC(=q'=&�&=�i%=]$=~�"=h� =��=��=|k=�*=\�=B�=��=^�=i=f=��
=F		=�G=k=�l=9M=s!�<̓�<O��<F�<N��<��<ʆ�<��<��<�Q�<��<>�<�W�<�I�<3�<�4�<k�<��<O��<�}�<mj�<B�<�<.F�<�W�<�"�<���<�1�<�by<��n<�vd<��Z<R<�J<�B<,�;<��4<�.<Z'<�<R�<
z<V�<���;���;1�;�H�;��;�m�;kߗ;���;��n;�-K;��%;��:?	�:�6:�V�8����Tn��t�Ⱥ�K��&��G�k��@���������R�Ż�aڻ��� �|	��2�m������i"�&�K*���-�3e1�M#5��9��R=�v�A���E���I��M�$�O���Q�T�S��7U�H�V�ĔX���Z�K`]��J`�Yc��Pf��h��8k�m�4�n��o�r�q��rs� �u�w�x���|��N���n���������Z;��ܝ�������G����������ڳ������;؋��6��ߌ�Ӎ�5��ph���֑��4���i��Zi��S8��B떼����wr��z��<��� A��M라(���,M���̢�����-���(��#���:��.���� �����$��rt��mԳ�3$��$D�����[�������%g���ս�w��I7��_j���  �  tO=�N=GJN= �M=�M=KAL=�yK=��J=J=��I=\	I=��H=�+H=a�G=G=tiF=S�E=M�D=�D=XFC=�B=�B=�A=�A=��@= @=(g?=�>=͢==�<=x;=�Z:=QL9=�Z8=��7=Q�6=;�6=�G6=�(6=6=6=�6=��5=	�5=�F5=��4=�4=�o3=��2=: 2=�1=�!1=M�0=oc0=!�/=�/=(�.=1.=�`-=��,=S�+=��*=�)=�4)=hs(=y�'=-�&=
�%=�G$=�"=�� =4�=�=§=�l=$:=�=9=�+=8]=F�=��
=�;	= x=��=H�=|�=+��<$��<?�<h��<3�<i��<���<�m�<�L�<��<"��<���<R�<�<��<"=�<G��<c!�<I�<�Ԩ<3Ĥ<ϙ�<1;�<K��<���<'w�<8�<���<�Kz<l�o<I�e<\<�2S<fK<�C<kn<<��5<k�.<��'<�c <M�<�C<�<,6�;�(�;�V�;B	�;cc�;�;�;�;�;���;�l;��H;�*#;Y��:�W�:L�4:�T�8���~���#ĺ���nb#��&E�ڞh�y���ɚ��B���Ļ�ػ��� ����u��(��������!�H�%���)��--�0�0��z4�8n8���<���@��E��	I���L�S�O� �Q�5�S��U�4FW�t*Y�n][��]���`��c�~Ef���h�ƾj�fl���m�q1o�p�p�_�r��;u�\Ox��{�����
�����A	��1���]�����iƊ��$���I���Q��[�����⋼)����v���������{��}璼�1���L���8������ӗ�����ř�3	��v}��?�������=��Ƞ���У��פ��ɥ�¦��ܧ�O0���ʪ������ͮ�����l��(���oƷ�+���O
���%��m輼8a������vؽ�����  �  AO=w�N=�N=w�M=�EM=��L=ӴK=��J=?1J=i�I=s�H=�yH=b�G=�pG=B�F=T.F=7vE=�D=��C=�TC=\�B=�BB=��A=�`A=�@=�R@=C�?=�>=��==M�<=׼;=�:=�9=P�8=@�7=�_7=��6=�6=�{6=h6=?\6=zJ6=�%6= �5=��5=��4=�_4=]�3=��2=IK2=@�1=*$1=U�0=�;0=��/=�B/=��.=��-=�7-=k,=�+=�*="*=6n)=۴(=��'=q�&=��%=��$=i�"=�2!=�?=�*=� =��=
�=��=��=Ɨ=�=��=?=s�	=ƹ=)�=��=��=_�<�{�<}��<=�<7h�<@��<���<:�<{��<��<W�<q�<T��<���<;��<�@�<ս�<�r�<�S�<lJ�<@<�<7�<ੜ<��<��<B�<��<�0�<��{<u3q<h2g<Ѿ]<(�T<��L<T�D<��=<Y�6<��/<��(<�\!<5�<<P<�<�S�;r�;F��;@�;���;Ħ;'�;MA�;b�g;:&D;t;��:���:�q0:��8,�⹉�x�S���<�������A��he�A��`-��k���»xֻ(����p����uV�m:�xL ���$�O�(��K,���/�ȝ3���7�2�;�I�?��D�^-H�0�K�c)O�m�Q�1T�@4V�W"X�`&Z��Z\���^�BRa���c��Gf��_h��j�[�k���l��,n���o���q�AWt��nw�� {���~��z��Jx���P��vzB��/H�������p������fƊ�ߊ�U���q�����J����'��⅏�� ���~��m瓼�*���C��>>���.��I+��6E��K���C圼�Z��pП�I/��g��$t��Wc��uI���?��_��׹���Y���<���V�������ֲ�������7Ƹ��6���V���'��R���]���R�������  �  yO=�)O=��N=�0N=��M=�L=��K=�K=�LJ=��I=��H=FH=�G=-G=+F=�E=�1E=��D=+�C=(]C=��B=�tB=�B=S�A=z$A=*�@=��?=b?=�>=�==�<=;=�:=�59=�{8=�7==l7=�7=��6=��6=V�6=9�6=�\6=�6=Z�5=�<5=��4=��3=�13=�t2= �1=�1=�0=� 0=�y/=��.='R.=��-=9�,=/G,=ؖ+=��*=�K*=��)=�(=o,(=X;'=�&=��$=�4#=<u!=�=U�=�j=�J=�-==z=�=�7=~b=��=��	=��=�=� =	=g��<��<�N�<��<��<�<�h�<e��<�n�<���<�a�<���<�	�<,T�<s��<�1�</�<.��<��<u��<���<V}�<M�<_g�<�~�<c�<�%�<ރ<[E}<�s<�@i<��_<>�V<'�N<��F<�4?<��7<��0<u�)<�R"<P�<_Y<��	<�� <�;�c�;"��;���;�ߥ;�S�;Hς;j.b;[>;�3;���:�c�:K�(:\��8D'ع<�n��i���s���}�b�>�$qb�d������	࿻:�ӻ[����������m�������s#���'��f+��/��2��6�)�:�w�>��$C�SG��FK�d�N��R���T��#W�[Y���[���]��`� Jb�Hyd�\pf��h�l~i�]�j��k�U*m���n���p�|s��v��z���}�<ـ����� q�������<��SD��P����}�+��G\��$�����뤋�J������s������������v��rd��2������dϙ�	����0���y���Ǟ��	���0���4�����,bɤ�����:妼@H���nͫ��ۭ�A��+��t;������Ƿ�0���V���;���廼Z`����� ���  �  ͢O=�OO=a�N=�[N=��M=T�L=L=;;K=ZJ=��I=�H=�G=�RG=��F=pF=�pE=8�D=�HD=k�C=eVC=��B=��B=[;B=��A=�RA=�@=B�?=�*?=N@>=CI==-P<=�_;=��:=5�9=�9=Ir8=q�7=��7=�B7=n
7=��6=�6=��6=�A6=W�5=Oi5=v�4=p4=[3=Ǐ2=y�1=O1=V0=�/=>/=_}.=L�-=�F-=]�,=Y,=�~+=��*=Xg*=�)=J*)=(a(=�m'=vH&=V�$=�c#=Q�!=��=�=
�=��=N�=7�=�=d�=D�=2�=��=A
=-6=�M=�Q=�<=| =�~�<���<V��<2��<�<$.�<n�<���<��<�{�<���<)?�<��<jG�<��<��<E�<j�<Q�<"�<Tȡ<�V�<F��<~˓<�Ď<��<���<�~<u<�k<�9b<yHY<v�P<��H<�@<19<��1<'�*<�
#<wF<�<�
<?�<�y�;s�;�H�;�9�;�p�;��;gQ;��Z;e6;��;#�:���:Bv:Ď�8��չqi��=�����G�C�<�-�`����z��}-��8ս��ѻ����B���^
�~Y�o��YG�@"�^�&�R�*��.��>2�o6�
:�{*>��lB��F���J�.�N��bR���U�7dX���Z��D]�P}_���a���c��We�b�f�$h�=i��j�Tk�Njl��n�TAp���r��u�[y�!�|��=��9����1脼 ���(��g��7����5��{����뉼xD������X���3���M��ݣ��7)��Z̑�y�����W�������a��젚�؛�����9��D[��e���P�����>ܢ�����$i���`����������]���l{��]w��ۀ��<����g���$��ղ������?��r>�����᲻�2:�������  �  ϴO=[O=#�N=�iN=H�M=9M=P.L=�CK={QJ=�`I=a{H=��G=m�F=Z/F=ˊE=�D=6lD=|�C=��C=�;C=��B=�B=�NB=e�A=vdA=5�@=�	@=�6?=�T>=�l==�<=��;=��:=8:=�9=� 9={8=�8=r�7=,N7= 7=8�6=ٓ6=)L6=�5=1y5=]�4=C34=k3=��2=��1=��0=�0=�P/=R�.=�-=�a-=��,=@G,=*�+=�S+=��*=Nl*=��)=C)=Az(=��'=	[&=C%=�z#=-�!=� =�'='>=�K=�Q=aP=:H=�<=�2=�/=e6=�E
=�X=�f=�g=*T=�& =��<���<� �<���<���<A��<��<���<-#�<�n�<o��<O�<���<]��<���<µ<v�<��<g*�<��<�١<�b�<���<'�<���<�
�<��<�G�<�w<'�m<Ðd<d�[<�R<.AJ<�B<5&:<~2<��*<�Z#<��<�r<4�
<��<+"�;���;k �;Z"�;�h�;Q��;*�w;�[R;�-;�X	;"�:���:�T:cD8S�޹�i��h��@�����l<���`���������F���>��Y�λR`໗=񻁠 �n2�_L�~�����T=!�&��U*��O.��2�|�5���9��=�� B��zF�G�J��O�S���V�5�Y�6�\��N_��a��|c��&e�l�f��g�_h�i���i���j�l���m��p��r��u�b�x�9C|�Qx��<������ރ����~��� ���և������!���������E����C��$��[+���z��������}���K��w��6����4��ۗ��ߜ����G������堼�����5��΢��u��V?���:��q���㧼=����Y���;�����Vﰼ����n1��h������*���F���A��-��ӻ��w���  �  x�O=|HO=D�N=�WN=I�M=��L=�"L=F1K=�0J=),I=�-H=�>G=veF=~�E=��D=xkD=��C=ȓC=�HC=�C=��B=��B=�CB=@�A=rUA=�@=��?=�%?=qN>=�x==I�<=��;=JI;=ȫ:=�:=0�9=��8=+m8=�7=,�7=�!7=D�6=��6=,86=��5=0h5=��4=�(4=�]3=t}2=U�1=�0=��/=�.=R.=o-=��,=�L,=3�+=�q+=p+=N�*=oW*=T�)=�<)=s(=�x'=\M&=N�$=ot#=Q�!=�" =>a=��=q�=~�=%�=�=��=y�=4�=l=ba
=D`=b=^=�J=�  =���<���<��<���<���<�H�<9�<	�<��<�K�<{��<�F�<��<	�<�-�<�m�<���<��<Q�<�<���<0�<W��<	Γ<��<�C�<���<@��<$�x<O�o<,�f<'�]<��T<�K<s C<��:<��2<��*<:2#<n[<C<��
<q�<G��;i5�;Y��;$i�;ڟ;��;��o;
I;��#; ;�i�:πs:<��9��E�����p��P��,����x�8>>�4gb�����<��}��OA���̻]�ݻ)��W��Y2��m��J������ ���%�|\*��.��x2��E6�X:�)>�DQB���F�B5K���O��T��X��[���^�&�a���c�Z�e���f�<�g���h��i�)ti�ij���j�Kl�n��bp�ps���u�B�x���{�
�~�襀�ҁ��낼����*��������m���Ј�:���4"��㾊�wm��mA��tJ���������ґ�R���̦��Ė��o��v!��n���w���1$��-��4砼
���l���z����������\T���U�����n������ o��1��&殼�~��[���W��R����뵼O-���g������#��������h���  �  �O=�O=��N=�(N=��M=��L=��K=-K=��I=�H=��G=��F=��E=�E=ZlD=��C=�wC=#+C=f�B=w�B=i�B=kB=B=�A=�)A=s�@=��?=�>=�0>=�o==�<=�"<=��;=�;=�:=��9=�]9=0�8=]+8=��7=�#7=��6=�`6=�	6=l�5=�:5=�4=4=o73=�P2=W1=�V0=�Z/=�n.=&�-=�,=�F,=��+=�b+=�+=��*=�*=\,*=��)=�)=O(=Q'=O#&="�$=�T#=��!=+ =��=u�=�=qI=�[=�Q=�.=��=	�=�=�f
=�O=&C=|8=�$=��<(u�<B��<��<
r�<w�<ӫ�<L�<��<Y��<�'�<B��<�9�<�$�<�G�<7��<��<�P�<J��<�<���<D�<Jǜ<�+�<��<��<bU�<��<^��<
Qz<�q<A�h<y_<�;V<��L<��C<?;<ڪ2<4�*<��"<޵<��<�0
<J<���;��;�N�;�5�;���;��;�$g;�?;�^;���:M~�:�YV:2%�9�α�3E	�0�}�n��v���l��@�A�l�e�(Q����������Iۺ��o˻@\ۻk��m ��4|�A�����k��Y �۸%���*��0/��;3�7�3�:�F�>���B��UG�l�K��P��2U��Y��~]���`���c���e�@�g���h�-mi���i���i�1,j���j�w�k���l���n�8#q���s� �v��[y��{�O~��3��+���������-���O���y��c���ʦ��J���Z��d��͋������#Ꮌ�b��>"������#���8���;��������:���=�� ��ơ��;��ɓ��S梼�K���٣�:���������n��(��+���XS��}ծ��3��Hs�������ϳ��	��nU��ҭ��s���Q���}�������  �  2ZO=a�N=�iN=��M=�RM=��L=}�K=��J=ҽI=&�H=N}G=^iF==oE=/�D=�C=�bC=�C=v�B=n�B=m�B=wdB=�3B=��A=�zA=��@=B@=�?=v�>=^>=�W==;�<=$A<=-�;=X;=��:=bM:=9�9=_9=nU8=��7=w7=ח6=$,6=��5=�j5=��4=<t4=��3=!3=2=�1=�0=��.=�.=1 -=r`,=��+=�L+=��*=��*=�}*=�B*=1�)=�)=i�(=�(=1'=��%=��$=K%#=��!=k# =k�=x=d=)�=w�=��=D�=�?=��=��=q[
=�.=�=�=%�=R��<m�<�M�<�F�<��<$��<>	�<��<�'�< ��<��<���<	B�<%G�<:��<t�<9i�<(԰<��<4�<�<'��<�?�<<��<F�<?��<-I�<G�</�<�u{<R�r<;j<x�`<�uW<��M<weD<[*;<�T2<��)<b�!<)�<�<�O	<�t <A�;?-�;6R�;�կ;Z�;j��;�[_;\c7;��;���:�њ:�::���9�3*�}����p`ú���#�c:F�zKj��K��o+��r���麻v�ʻp�ٻ��_��"��
� � '�N����%��S+�
0��:4��8��;�6�?���C�74H�#�L���Q��oV�[��6_�v�b���e��
h��i�؃j�v�j�6 k���j��k���k�til���m�x�o�2&r���t��lw���y��4|�� ~����<����~��l���~��򵄼����Y��K���z�������A����K���!�����T���ϐ�r����������tߘ�������ǳ���!���?���������*���e������wF�����(!���p��C屮턪�"��ّ���⮼�	��������(���W��������������!��N���U����  �  d)O=ȤN=�(N=�M=dM=cL=3�K=8�J=y�I=�ZH=�0G=WF=^E=d0D=CC=�B=�B=�qB=�UB=�BB=8)B=9�A=�A=v?A=ƭ@=@=�D?=��>=��==3<==e�<=�Q<=�;=��;=p;=�:=��9=�09=wo8=��7=97=�q6=�5=��5=�)5=�4=R74=l�3= �2=��1=��0=��/=˭.=t�-=�,=��+=+\+=�*=��*=�c*=�7*=@*=%�)=N)=��(=.�'=��&=��%=yY$=��"=B�!=� =y�=�&=֕=�=U=��= �==n=y=�=iI
=
=��=0�=İ=n�<D��<r��<T��<��< �<$y�<$��<�k�<1�<�E�<M��<Wx�<я�<�<�a�< �<#Z�<ʤ�<n��<?��<�6�<���<q2�<��<�^�<�/�<�$�<�(�<�A|<p�s<�#k<��a<QX<�}N<�D<O;< �1<E:)<�� <j�<��<pb<�#�;�^�;�h�;�h�;���;ɡ�;:��;tY;�0;?�
;���:��:Ɲ#:'�F9
Gs��+�Z��RI˺|���e'�k�J�-�n��9�������h��,.���'ʻ��ػ+�滳}��*�Z�	��S�L�����JA&���+�p�0��75�i"9�K�<���@��D�I�g�M�|�R��W�FH\�,�`�efd�pg�ưi��+k���k��0l��l�H�k���k�Hel��Nm�m�n���p��*s�¼u�\Fx���z�(�|��~��k��W�����~큼���I�������3��Ӣ��<퉼A����ˌ�N���e����ˏ�BA��� �����D0��Fr�����������������w���Ӣ�~J����������ߣ��.��ܶ��z�������#��p�������|��b֭����������ְ�Ƕ��򰲼	س��2������aa��9
��!��������  �  SO=�xN=�M=�wM=��L=s6L=wcK=�kJ=~UI=-+H=��F=��E=��D=*�C=�:C=��B=ofB=�8B=l"B=:B=��A=��A=��A=hA=z~@=��?=�?=&]>=�==�&==g�<=OY<=�<=b�;=$=;=˲:=�
:=vJ9=}8=v�7=#�6=�T6=��5=e`5=i�4=�4=K	4=�f3=͞2=�1=��0=��/=Mw.=Wk-=*|,=.�+=\+=%�*=�]*=�,*=�*=��)=��)=%)=��(=H�'=.�&=�|%=&.$=��"=�j!=� =A�=#7=��=�=�/=�#=h�=܈=.=��= :
=��=��=��=z�=?��<�K�<m��<���<�>�<���<}�<Uq�<D��<p��<ݺ�<T(�<���<��<�v�<��<
��<� �<�K�<&\�<�0�<�ӟ<X�<Mؖ<�m�<q+�<h�<s,�<�L�<˸|<�~t<��k<ˆb<�X<��N<��D<=�:<�1<��(<_I <�"<Y<s�<1��;�;��;w�;�$�;��;��;F�T;�#,;.";� �:簅:�0::�9�5��^�7��ה�t#Ѻ����*���M�%�q������Л�����p����ɻ�ػ�滧^�����x5	�����������&�"h,�0�1�j�5���9�D�=�qlA��mE���I��nN�!WS�5QX�
$]�a�a�3ke���h�
�j��1l���l�Em�3�l��l�'�l��m���m���o�_�q���s�Auv���x�l{���|�M"~�T;�'��Pˀ�4���ݷ���
��ڋ���!���������6G��5H��)��N��c���<&������qU���W��Ō��#ؙ�����1�� ���}������S������C���g��h8��������ޥ������R���Щ��V��Ǭ� 
����������@���j�� ���?봼����=��x�������0���  �  ��M=PfM=TM=d�L=�JL=G�K=�J=�J=�H=��G=)1F=1�D=s�C=^�B=��A=��A=%VA=&SA=�kA=�A=��A={A=�.A=��@=��?=�?=�;>=Ui==Ͻ<=4E<="�;=��;=x�;=;�;=9;='�:=�:="9=/)8=�.7=K6=1�5=*5=y�4=4z4=�>4=I�3=�k3=[�2= �1=��0=�w/=O:.=�-=�,=�0+=ğ*=�O*=�5*=�=*=-R*=�Y*=�=*= �)=�Q)=�q(=�P'=��%=d�$=�&#=��!=�� =�H=f	=_�=T=�E=�%=�=�!=�f=O�=
=��=TV=�D=�I=���<�]�<��<���<�G�<	x�<.s�<�c�<�x�<1��<���<��<���<]J�<�<.��<�~�<b�<�i�<�]�<���<eM�<}��<˔<�L�<L'�<\[�<̈́<�P�<�g{<��s<��j<ka<�W<FL<-NA<b�6<�,<�k#<� <^t<��<�T<�#�;���;���;m�;F��;_6�;��j;��<;z�;���:��:� :�OA9��_�2��r􂺎Ϻ����l���1B���h�����#����(���/��&�ʻfػ����$�5 ��������'� � ��(�]D0�ס6���;���?�KC�VF�*I�\lL�YiP�9U�?$Z���_���d�O�i�{�m��2q��Is�J<t�9t�#�s�ۄr�Ԋq���p�|q���q�G�s��Lv�\Fy�uN|��~�@����!���l��݉��L��������������:2������s�*܊�Վ��a獼Rݎ�_����������샑�Œ�{x��Ӗ��J��ݠ��:������$���]J��>U��Zۥ�`���ҥ�f����o��������3�kK��L���ɫ�w������F��v��؊��P汼�R������&��au��bF��YY��:���0����T���  �   N= �M=#M=\�L=�aL=��K=�K=LJ=[�H=��G=PHF=��D=��C=q�B=�B=��A=�sA=$mA=,�A=��A=��A=��A=lAA=��@=�@=8?=�W>=��==g�<=YX<=�<=V�;=$�;=b�;=�,;=b�:=i�9=9=�)8=�67=�Z6=��5=�'5=c�4=~�4=�W4=4=H3=O�2=��1=��0=��/=�R.=h(-=�",=_R+=N�*=so*=�Q*=VV*=2g*=�l*=O*=l�)=�d)=ֆ(=�h'=�&=�$=
@#=0�!=�� =�O=�=��=�=�6=X=��=�=]f=��=
=3�=n=S]=1a=���<���<���<6��<Rg�<s��<���<]��<��<��<9��<>U�<�5�<���<!�<��<Z��<�A�<E��<��<y*�<���<
��<h�<˃�<�T�<�y�<�ڄ<xN�<ZI{<8fs<��j<+6a<��V<�5L<"ZA<��6<��,<��#<Q�<-�</]<ȧ<��;s�;�Z�;���;Õ�;l�;ܥl;g�>;��;�M�:��:ȏ(:e*^9MPF����D���*��'N��c6��~@��f���������O��ă��@;ʻ��׻E��_�; �8�����<�N� �N�(�0��E6��^;��f?�P�B�L�E�حH�|L�` P�R�T� �Y�'._��qd�Pi��xm�h�p���r�A�s���s��%s�\/r��>q���p���p���q��ls���u���x���{�7�~�!T��( ��[��Y������K������σ��D������눼�Ɗ�*j��&���򦎼�M��0׏��v��OY�����U���r��iߘ��t�����fi��ts��������
���¥����xl���J���g��7⥼�ʦ�����©�ݑ���X��o箼1��� ~���豼a��8����������U��]��0w���t��5+���  �  �DN=��M=�nM=FM=a�L=�	L=~@K=�CJ=3I=��G=A�F=yHE=$&D=�3C=�|B=�B=�A==�A=��A=	�A=��A=y�A=�tA=B�@=N@=`�?=أ>=v�==c==��<=.'<=��;=�;=�e;=�;=s�:=��9=T9=�(8=fK7=�6=��5=:o5=�5=�4=x�4=R>4=*�3=��2=�
2=&�0=5�/=��.=Bx-=�{,=��+=�+=��*=0�*=�*=�*=��*=�~*=�**=ݗ)=x�(=��'=k`&=��$=��#=="=� =�a==��=a�=	=^�=΍=�=zd=��=�?
=2�=�=��=b�=07�<���<KE�<�5�<���<0�<`�<a$�<�W�<���<O��<7�<p��<�&�<���<�b�<�<x��<��<��<��<^�<d^�<c��<��<�Ȍ<lƈ<0��<\A�<�z<��r<Qj<ߕ`<|V<9 L<�wA<}=7<[�-<��$<e�<��<e<6�<dY�;��;���;o'�;�]�;��;
�q;�D;�;���:�2�:R?:���93����r�������)�@�;��a����������%̹�(ɻy|׻5L�l)��� ��]�?U����� ��[(��T/��P5�E;:��0>�|�A��D���G�bAK�wWO��S��Y��=^��Zc�uh�l��1o�!Gq�Ur�1�r��r�a<q��ip���o���o���p�c|r���t���w�$�z��q}�
��|����,������ׁ��N��V
��7��g��"���߈�����	���5�����Ĵ��WE����}䐼�6��L󓼍��Tr��f���u��������`H��SW��Q祿�&���������#䤼_���}��+\�������6���������3\��K���Φ���^����x����X��`l��Ե������l���\���-�������  �  ��N=y4N=q�M=IsM=�L=�UL= �K=نJ=�cI=*H=��F=��E=��D=�C=C=W�B=vFB=�%B=�B=\#B=�B=< B=غA=�GA=,�@=T�?=?=5>=6q==��<=�L<=��;=�;=3;=��:=�?:=8�9=e�8=28=vb7=m�6=�46=^�5=��5=�E5=/�4=2�4="�3=<3=1N2=S?1=�0=��.=��-=� -=A=,=��+=�N+=�+=�+=��*=�*=��*=Lk*=��)=`)=�(=��&=FZ%=��#=�c"=�� =t=E�=�_=��=>�=n�=�M=�=Z=�=t
=�-=�
=� =}�=���<�y�<`��<��<B�<���<?��<c��<�P�< ��<5��<q4�<:��<7�<���<��<��<MB�<���<���<�h�<��<�6�<A{�<֑<jb�<L'�<��</�<'+z<;�q<Q�h<�_<M�U<�K<ׄA<��7<��.<u&<�<Oq<��<0�<E��;���;���;B\�;]��;F%�;R�x;;�L;,#;R��:���:'ya:�s�9R�������]��W����]����5���Z������0��Y���&�ǻ�.׻������t���`	� 4�y��� �]�'�s.�P4���8��<�Z�?�;C��dF��J�YEN���R�.�W���\�&�a��-f���i��l�/o��9p���p�gp���o��;o�L�n�)�n�޲o�R5q�,hs�Zv��y���{�=h~�s4��J�������*��꿂�Đ�������腼b\��݈��J������Z���TI���㍼�}���=���E��é���m��9���W֗�g?������ɞ�5���,��"?���飼b>��BV��YQ���S��?�������.ƥ������v���,��[�����D��;G���>����沼�ӳ�����}Q��:㷼����9D��ռ�?-���  �  ��N=ݜN=R?N=W�M=�LM=�L=��K==�J=@�I=ӃH=:[G=#AF=�AE=VfD=j�C=t4C=��B=B�B=7�B=�xB=�eB=�@B=��A=��A=��@=�F@=�u?=�>=��==�==5i<=��;=_;=�:=�g:=��9=�E9=̤8=?8=n7=��6=�6=|26=Y�5=�5=ZW5=��4=�C4=n|3=9�2=T�1=X0=�u/=�|.=��-=b�,=5V,=�+=�+=�{+=�Z+=�7+=�+=,�*=u*=�X)=�W(=0 '=��%=�;$=_�"=�!=y=��=�=*D=�K=G.=��=��=
==��=�
=v=Pc=�]=�U=�: =��<�7�<;�<���<r2�<��<O��<�x�<�2�<�5�<��<=�<�9�<w�<�<,`�<+ذ<�,�<sH�<��<���<<�<�V�<V��<���<|y�<g�<`р<�y<�Fp<�?g<��]<�aT<^�J<9SA<W08<˃/<�V'<��<��<�0<�<5��;���;��;s��;Ь;R��;�؀;zW;�2.;$�;���:�+�:�:|S�8����
LH��x��8�ٺ�x�/��T���y�},����lT��D�ƻTO׻�H�^����(��
�Ł����"!��'���-���2�k7���:��<>���A�HE���H�=M�z�Q�ҙV�IX[���_���c��{g��Qj��cl�w�m�_[n��~n�oLn�3�m���m��m�՞n���o�`�q�K�t�5dw�iYz��#}�H��o׀����T����h��T���^��쇆�����z���������ۋ��}��6��㴍����<���#���쒼:���
/��Oo��˝������{c���ՠ��˱���,��
r��4���[���u���[s��T6���N�����\��o ��s⬼��������8��nZ��kn�����������	���q��⹼�F������H����  �  EO=!�N=�N=�N=8�M=G�L=��K=-�J=>�I='�H=m�G=�F=%�E=RE=�lD=��C=NxC=)C=��B=��B=�B=\kB='B=��A=A=A=��@=g�?=��>=�>=e5==�n<=�;=;=|:=~�9=i\9=�8=UK8=q�7=�a7=�7=��6=�~6=�C6=$�5=��5=�5=Qp4=N�3=4�2=��1=0�0=�/=�/=F.=��-=�	-=Q�,=;,=+�+=ܳ+=�v+=�.+=0�*=ID*=r�)=�(=�f'="&=y$=��"=�&!=zd=�=Y�=��=��=N�=r=�;=�=
�=��
=ܦ=,�=��=��=Gn =N�<vx�<Za�<-�<<��<fK�<\��<2��<F��<K��<���<L��<`�<f�<���<r�<DF�<���<��<i��<Q�<<X�<�3�<�`�<���<��<�O�<�rw<�Hn<�e<k�[<��R<a�I<	�@<�48<"0<�C(<Ū <<�.<��<���;��;��;&n�;�[�;�9�;�L�;|�a;��9;��;�G�:=��:�2:��X9�5����6�!"����Һ	�P�*��N��t�|S��絠�>̳�TSƻ�1ػ^j黨���C���D��U���!���'��1-��1���5��~9���<��x@�|5D�??H�ؑL��Q���U�0�Y�G^�p�a���d��g�t�i��k��l��l���l���l�2m��Gm�_�m�^!o��p��Is��v��"y��5|�!�瀼����=��#M��'U��<\���a���]��&H����9Ȋ��Z���݋�:j��s�����hF��	ΐ�Ԙ��!���נ����������n��"
��	j��D���#l�����$�������GG������-!���٤�'ۥ��(��?����z��2P�����*ү�bc��_ղ�0/���y������k���.9��{e��Kz��)p��C���  �  �gO=�O=ƹN=7;N=?�M=�L=��K=9�J=T J=0	I=H=�BG=�xF=L�E=GE=��D=<	D=Y�C=�>C=��B=�B=qB=P)B=}�A=IQA=�@=��?=C?=�+>=<==�S<=�x;=`�:=��9=�Q9="�8=eA8=��7=}7=
67=d�6=!�6=�6=:o6="6=z�5=I%5=�s4=��3=��2=��1=�1=�L0=��/=��.=AF.=8�-=�5-=��,=W,=��+=�+=s9+=��*=�A*=��)=)�(=R�'=,)&=��$=!�"=0!=&/=8=�3=^%==�=�=(�=T�=a�=E�
=�=2�=��=E�=�v =jH�<rg�<_X�<q/�<0�<���<B��<���<���<��<�^�<���<�k�<{0�<� �<Z9�<�n�<3��<kթ<{ե<���<O�<�g�<܂�<;��<��<@��<K%<�ju<��k<�~b<�ZY<�yP<��G<7�?<��7<i0<�(<I*!<��<ԃ<�	<s��;���;O�;�A�;5!�;��;]S�;��k;YGE;�;�	�: ��:ĒS:�_�9�"E��-�WD���Lкϟ���(���K��p� ����r��?R���ƻ
ڻp컺	���[��.�_s����"#��(�[@-��o1��45���8�QP<�B@���C��(H��L��P��U���X�|s\���_�%`b�+�d���f���h���i���j�u�k��[l�N�l��:m���m�c�n���p�޵r��hu�Ղx�m�{�d/�6������!���g������
���&r��3��cӉ�?V��q���E!��������d׌�����s4���ɐ�~����l��I�����FÙ��R��.������3��D9��o��ޡ������������q���Ϥ�����7j���#�� �������ﯼ̱�Ɗ���'��i���9����)��(8��#���뻼̕��)���  �  (`O=�O=��N=q)N=zM=ΪL=`�K=��J=��I= I=�XH=r�G=��F=�WF=	�E=VE=�D=��C=!qC=��B=��B==LB=��A=�A=5A=�@=,�?=C?=O!>=�==0<=";=l/:=�[9=ϥ8=�8=e�7=nI7=D7=��6=�6=r�6=:�6=�l6={6=�5=5=oH4=!~3=Ѱ2=��1=�81=�0=t�/=�l/=��.=iQ.=��-=R/-=�,=�,=��+=_+=֞*=*=�b)=	�(=p'=�&=��$=��"=!� =��=D�=5�=As=�O=�5=>)=+=�:=U=ev
=�=t�=)�=*�=pO =?��<f��<N��<x��<	�<j/�<k�<��<�<�O�<>��<i��<qF�<���<�f�<�=�<�C�<�i�<���<ʥ�<���<j�<Bn�<}�<�Z�<m�<.ڃ<�D}<*
s<Ci<5�_<ҋV<H�M<�E<X><c�6<G{/<�N(<� <gE<�<9j<܄�;?��;6�;1��;߱;t�;蔌;Lt;�jO;�[*;�';(�:�!n:�|�9�&�b�,�^���s�Ӻ�$	�&�)�|�K��Fp�Df���y������Ȼ.�ܻ�8��Z���	�������>�>�$���)�"�-���1�T75�t�8�4j<�8S@�
{D��H��M�$@Q��U�waX�_P[�h�]��6`�7[b��dd��Wf��*h���i�#5k�Tl�.m�Z�m��n���o���p���r��ru���x��|������ ���4������(ꇼBꈼ�����7������JԊ�����8��������I�^������l!���ے�唔��6�����G��7d������
Ҝ����+1���R���_���O��T��Wϣ�s���#�����z���x��$'�����3+���Q���o��s���L�����V��7|���b��������_����Z���  �  �4O=u�N=��N=l�M=�0M=�XL=dtK=D�J=��I=RI=�tH=A�G=%_G=��F=�:F=��E=��D=N/D=�C=��B=KjB=>B=��A=cTA=��@=k@=K�?=:�>=��==��<=��;=�:=��9=�8=$�7=6[7=��6=��6=2�6=��6=K�6=��6=�w6=B6=��5=w^5=&�4=1�3=�.3=Rq2=2�1=d91=M�0=�K0=;�/=#^/=|�.=0.=��-=.�,=�,=u+=�*=QL*=��)=9)='=(=b3'=��%=5[$=W�"=ƒ =�p=�8=��=�=�=8r=�r=��=�=��=�(
=�Y=fu=�q=!J=��<�/�<dB�<S�<�|�<���<HE�<U��<Dj�<���<yY�<H��<���<^��<��<�j�<���<�ΰ<�٬<�<� �<0�<�Ɯ<V#�<&-�< �</��<	�<.({<��p<]Gf<ؠ\<�S<�NK<-�C<�D<<uJ5<n.<lu'<Z) <�a<�
<�,<@��;��;Y��;
��;J��;�&�;�;�1{;��W;�D3;�;��:Չ�:4l�9�)���5�����S6ܺ�L�*+-���N��zr�>b��)��������ʻI�r�������&��*����!���&��+���.�Dd2�o�5��\9��,=��JA���E�J�!TN�7R�&�U�"XX�1�Z�K�\��{^�R\`�wbb���d���f�[i��k�F�l�� n�'o���o���p���q�7�s�� v��5y���|�Fl���|������^������*T��mQ�������V���|������N����������v���a��F���!���Ǒ��r��\���f�����O�����������Bϛ�
��Y`��������^��vs���W������ȥ����������ڨ��z��j��{����簼�<���y��a����N��Oú��ܻ�g���m��@j��;����ʽ��  �  w�N=��N=�9N=ŗM=T�L=��K=VK=�8J=��I=��H=WxH=dH=�G=�/G=h�F=~�E=-%E=oPD=�~C=Q�B=, B=��A=tAA=[�@=r�@=<@=�x?=H�>=��==�<=Kg;=�7:=�9=�8=gJ7=!�6=YN6=�6=�6=�$6=�;6=-G6= 76=[�5=r�5=�5='P4=#�3=
�2=&2=W�1=�"1=K�0=�0=�*0=�/=�0/=K�.=�-=�,=�,=�<+=��*=z�)=sJ)=T�(=�'=��&=f�%= $=GB"=v7 =,=r�=.Z=e=��=/�=��=q�=�3=ށ=x�	=�
=�(=v =`�= /�<�O�<�_�<��<���<Jh�<l,�<Y�<���<E��<|$�<�c�<�i�<N�<s3�<�=�<��<�+�<��<_<�<h�<?s�<:�<���<䯒<>c�<�ׇ<�-�<�y<�n<h�c<��Y<M�P<��H<TA<te:<�3<x$-<M&<P<�<:�<�<8j�;y��;��;�l�;=��;Zf�;*g�;�;�5^;� :;��;u��:dr�:X�9i<E���D�F?�����^��o2�P<S��bv�5*��'z���ҷ�g�ͻa��x����;�mF��?�����#��(�
�,�o 0��m3�{�6��`:��W>�	�B�0G���K�Q�O���S�rV�z�X��aZ�>�[��5]���^���`�[Dc���e��h��ek���m�jo���p�l�q��Rr��^s���t��2w��7z�y�}����UE���v�����MC������k���$6��fo���h���@�������b�����M��\���򚒼�5��q����Ö����Jr��//��4��p
���M��ɝ��h��:����������
��7䥼�����W���>���p��d����물�&��5����� ��ڴ�� ��� ���*���ӽ��)���F���K���\���  �  ��N=�hN=Z�M=�@M=�mL=��K=��J=��I=<I=��H=�mH=�%H=��G=(oG=j�F=,*F=%OE=�^D=ImC=ݎB=��A=�CA=��@=|�@=0@=q�?=j.?=]g>=�n==$M<=�;=^�9=�8=��7=��6="6=�5=��5=��5=��5=7�5=L6= �5=i�5=rG5=��4=��3=�"3=�d2=A�1=�P1=r1=n�0=c�0=�_0=��/=(s/=�.=�-=��,=��+=��*=�0*=�~)=��(=};(=m{'=��&=�N%=z�#=��!=V�=�=T>=M�=Yz=;=�#=�7=bp=E�=�!={	=��=��=��==�=�d�<�v�<���<���<�1�<���<���<k �<�7�<�<߰�<���<���<��<B1�<=��<��<σ�<�Y�<}v�<N��<,ʟ<��<0�<(-�<�׌<x6�<�l�<uFw<l<]a<��W<ͣN<��F<�r?<��8<_2<)�+<�'%<��<��<�,<�<��;�O�;�;�;q>�;X�;1�;�8�;�ȁ;��b;��>;�I;�y�:!��:q��9{�k��OU�ױ��������7�-X�Ԣz�b���j�������7л��滶.��>��m�Rn��) �ճ%�%:*�S�-��K1�vw4���7��s;�ߏ?��D�h�H��LM�9oQ�t�T�BgW�+Y�a]Z�oP[�O]\�)�]���_��db��pe�p�h��k���n��p��1r��&s�i�s���t�>3v�`Qx�}C{���~����$����J���t���Q��Iŋ�t����?��]���4���쌼��������錼Ǖ��g������T����j������;��-���ؗ�9\������􍙼ق���̛�xf��8�����|ꢼ�|��x�������k������屮��q���<q��E���95��vѴ�&^��%���k����6��z@��վ�y�������꾼�  �  �N=�5N=�M=� M=�&L=<K=TZJ=�I=^I=ˢH=�aH=q.H=��G=F�G=�G=�LF=�eE=icD=G\C=hB=��A=��@=܍@=>:@=D�?=J�?=p�>=^5>=�===�<=|�:=��9=�U8=�?7=	`6=��5=k5=�O5=ja5=��5=
�5=��5=+�5=��5=�5=g4=��3=5�2=�2=O�1=W!1=l�0=��0=@�0=n}0=F%0=/�/=��.=j�-=��,=1�+=��*=��)=�3)=N�(=D�'=F5'=�H&=%=1�#=��!=٨=�\=��=�~=�= �=l�=��=�=�x=��
=UA	=Ӈ=�=��=�Q=���<7��<|��</%�<���<���<���<*$�<}a�<�`�<�<x9�<v�<%��<�$�<�¸<Z��< �<%ʪ<��<&!�<�L�<�5�<���<�̑<�r�<�ņ<]�<�v<&�j<��_<��U<� M<�AE<�2><��7<�l1<
+<�V$<��<��<$<w�<���;z��;L �;���;?V�;��;���;ж�;)1e;R�A;��;Q�:���:��9_����b��ݹ��W���T���;���[���}�����ۥ��~����ѻ���p�����	�����s�!�~�&�=U+���.�r2��75�Ά8�@<�=v@��E�N�I��zN�V�R�J�U�-#X���Y��nZ��[���[�-5]�84_���a�,e�W�h��8l�Ko�I�q��Us�Xt�eu���u��!w�L%y��|������ur���؆�(��4������{�������l���Uc����n��`L��S���%�������Q��+��Ԅ��:���)�������W��R���+K���4�����/0��"���/���)��B䤼�C��F��M������Iq���~��񫼯ҭ��������R����]��g�����Z����G��������_���O���  �  TnN=r#N=L�M=5�L=kL=E K=�>J=�I=�H=�H=�\H=�0H=��G=�G=yG=�WF=qlE=dD=UC=wYB=�A=��@=r@=�@=��?=�n?=d�>=1#>=,==�<=��:=x9=7:8=� 7=�>6=$�5=�J5=�25=H5=�u5=��5=־5=i�5=�o5=%�4=�N4=ч3=A�2=��1=ln1=_1=5�0=�0=��0=�0=�10=��/=x�.=A�-=��,=��+=^�*=��)=E)=�s(=f�'=�'=�1&=|%=�#=c�!=�=PE=��=:`=G�=|�=5�=��=y�=�^=��
=r-	=u==�=j=�:=���<��<V��<i��<T��<݄�<���<�$�<�n�<!w�<��<�R�<�"�<o��<~�<㫸<I��<;Ԯ<���<��<J�<��<9�<<��<	��<7M�<:��<>��<��u<�+j<�W_<TpU<\�L<��D</�=<%Q7<51<y�*<5$<��<�<�<{s<���;��;�]�;�;O��;ȟ;���;��;%	f;��B;m�;�(�:4M�:��9T~��H g�E������"���=��]���#��>h������һ�U�p��,
�de�5l��"�:l'���+��E/�Bj2��}5�8�8�ڊ<���@��rE�TEJ�V�N���R��3V�0jX�üY�xZ�� [���[�5]��_���a��e���h��]l���o��r�P�s���t�wyu�C>v��xw��ry�>O|���J7��|����
��4Q���E��tƌ����r/���3��� ����<���'��sp���)���R��Ր������:��t����ݖ��������W�������5��'��k�����0��j8���A��X��iu��}��<��=ᨼ����F���j�������;��3̲�:���'��o��������8��U<�����nٿ���������Tt���  �  �N=�5N=�M=� M=�&L=<K=TZJ=�I=^I=ˢH=�aH=q.H=��G=F�G=�G=�LF=�eE=icD=G\C=hB=��A=��@=܍@=>:@=D�?=J�?=p�>=^5>=�===�<=|�:=��9=�U8=�?7=	`6=��5=k5=�O5=ja5=��5=	�5=��5=+�5=��5=�5=g4=��3=4�2=�2=N�1=V!1=k�0=��0=?�0=m}0=D%0=-�/=��.=g�-=��,=-�+=��*=��)=�3)=L�(=D�'=J5'=�H&=%=K�#=��!=�=�\=�=.=�=��=��=1�=i=ez=��
=�C	=E�=��=��=fT=S��<{��<���<�)�<���<K��<���<�&�<3c�<�a�<5�<�8�<#�<��<�!�<;��<c��<� �<OŪ<�ަ<��<VG�<�0�<���<�Ǒ<�n�<���<Q�<v<�j<��_<��U<s"M<�DE<%7><��7<�s1<e+<�_$<�<2�<�.<<�<���;��;�2�;a��;�d�;p�;|��;¼�;�6e;��A;��;���:+Պ:���9$���u�b�H,����������(<��[��~�����q����#һ˧�i��� �	�������g�!���&��W+��.� 2��85�ԇ8��@<��v@�eE���I��zN���R�u�U�M#X�̔Y��nZ��[���[�65]�?4_���a�,e�Z�h��8l�Ko�J�q��Us�Xt�eu���u��!w�L%y��|������ur���؆�(��4������{�������l���Uc����n��`L��S���%�������Q��+��Ԅ��:���)�������W��R���+K���4�����/0��"���/���)��B䤼�C��F��M������Iq���~��񫼯ҭ��������R����]��g�����Z����G��������_���O���  �  ��N=�hN=Z�M=�@M=�mL=��K=��J=��I=<I=��H=�mH=�%H=��G=(oG=j�F=,*F=%OE=�^D=ImC=ݎB=��A=�CA=��@=|�@=0@=q�?=j.?=]g>=�n==$M<=�;=^�9=�8=��7=��6="6=�5=��5=��5=��5=7�5=K6= �5=i�5=rG5=��4=��3=�"3=�d2=@�1=�P1=q1=m�0=`�0=�_0=��/=$s/=�.=�-=��,=��+=��*=�0*=�~)=��(=~;(=t{'=��&=�N%=��#=��!=��=��=2?=s�=�{=�<=7&=`:=�s=��=�%=�	=��=��=��=v�=�n�<׀�<���<���<+:�<���<��<%�<;�<��<C��<z��<a��<$��<�+�<���<#�<7{�<�P�<�l�<,��<���<��<��<<$�<�ό<i/�<�f�<W=w<��k<�Ya<j�W<��N<f�F<�{?<n�8<�l2<I�+<�9%<2�<��<UA<�<UA�;uv�;�_�;�^�;�s�;�G�;�I�;xԁ;��b;��>;1<;6F�:$O�:q:�9�lo��_V��n���*��EG��?8�oX���z��F��������x[л�滘K���J��x��w��1 ��%�8?*�d.�O1��y4���7�Bu;��?�kD��H�MM��oQ���T��gW�6+Y��]Z��P[�d]\�9�]���_�eb��pe�v�h� �k���n��p��1r��&s�j�s���t�?3v�`Qx�}C{���~����$����J���t���Q��Iŋ�t����?��]���4���쌼��������錼Ǖ��g������T����j������;��-���ؗ�9\������􍙼ق���̛�xf��8�����|ꢼ�|��x�������k������屮��q���<q��E���95��vѴ�&^��%���k����6��z@��վ�y�������꾼�  �  w�N=��N=�9N=ŗM=T�L=��K=VK=�8J=��I=��H=WxH=dH=�G=�/G=h�F=~�E=-%E=oPD=�~C=Q�B=, B=��A=tAA=[�@=r�@=<@=�x?=H�>=��==�<=Kg;=�7:=�9=�8=gJ7=!�6=XN6=�6=�6=�$6=�;6=-G6= 76=[�5=r�5=�5=&P4="�3=	�2=%2=U�1=�"1=H�0=
�0=�*0=޽/=�0/=D�.=w�-=�,=�,=�<+=��*=r�)=nJ)=U�(=�'=�&=��%=j$=�B"=8 ==��=�[=~=��=e�=��=��=�8=��=��	=B=�/=�'=��=�=�<1^�<�m�<���<��<kr�<�4�<��<���<��<
%�<9b�< f�<gH�<�+�<�4�<0��<d�<o�<w.�<�Y�<�d�<�+�<��<J��<�W�<�͇<N%�<�y<�n<Ɠc<w�Y<X�P<��H<s`A<�u:<��3<;;-<_f&<�<�:<��<A�<���;��;sK�;F��;{��;���;��;b/�;vE^;:;��;���:1�:���9�qJ��eF�p����b����2�E�S�O�v�Sg�������	����ͻ)��<���XM��U��L�����#�D�(�Ϡ,�%0�Aq3�K�6��b:��Y>�W�B�1G�`�K���O�
�S�erV���X��aZ�f�[��5]���^���`�hDc���e��h��ek�©m�jo���p�n�q��Rr��^s���t��2w��7z�z�}����UE���v�����MC������k���$6��fo���h���@�������b�����M��\���򚒼�5��q����Ö����Jr��//��4��p
���M��ɝ��h��:����������
��7䥼�����W���>���p��d����물�&��5����� ��ڴ�� ��� ���*���ӽ��)���F���K���\���  �  �4O=u�N=��N=l�M=�0M=�XL=dtK=D�J=��I=RI=�tH=A�G=%_G=��F=�:F=��E=��D=N/D=�C=��B=KjB=>B=��A=cTA=��@=k@=K�?=:�>=��==��<=��;=�:=��9=�8=$�7=6[7=��6=��6=1�6=��6=K�6=��6=�w6=B6=��5=v^5=%�4=/�3=�.3=Pq2=/�1=a91=J�0=�K0=6�/=^/=u�.=0.=��-=#�,=�,=u+=�*=GL*=��)=;)=3=(=�3'=��%=�[$=�"=�� =�q=:=��=��=+�=%v=�w=��=L�=��=U0
=�a=�}=�z=(S=� =rA�<+S�<�b�<֊�<=��<�O�<{��<p�<��<&Z�<b��<V��<u��<��<�_�<��<῰<�ɬ<��<3�<��<W��<��<��<�<z�<���<{{<vp<�Af<y�\<�S<YK<P�C<�X<<�b5<ډ.<^�'<�J <ׄ<�.<�P<a�;�"�;K9�;���;cɱ;(N�;
�;�Y{;��W;EB3;\p;���:��:���9�v/��7������Qݺ�����-�IO��s������蠻 鵻�3˻=F�ߣ�������
��l��g�!�c�&��+�5�.��h2���5��_9��.=�\LA�ݥE�J��TN��7R���U�vXX�q�Z�|�\��{^�n\`��bb��d��f�di�k�K�l�� n�+o���o���p���q�8�s�� v��5y���|�Fl���|������^������*T��mQ�������V���|������N����������v���a��F���!���Ǒ��r��\���f�����O�����������Bϛ�
��Y`��������^��vs���W������ȥ����������ڨ��z��j��{����簼�<���y��a����N��Oú��ܻ�g���m��@j��;����ʽ��  �  (`O=�O=��N=q)N=zM=ΪL=`�K=��J=��I= I=�XH=r�G=��F=�WF=	�E=VE=�D=��C=!qC=��B=��B==LB=��A=�A=5A=�@=,�?=C?=O!>=�==0<=";=l/:=�[9=ϥ8=�8=e�7=nI7=D7=��6=�6=r�6=:�6=�l6={6=�5=5=nH4=~3=ϰ2=��1=�81=�0=p�/=�l/=��.=aQ.=w�-=G/-=��,=�,=��+=R+=˞*=*=�b)=�(=?p'=<&=��$=K�"=� =��=��=r�= v=S=:=t.=.1=kA=�\=�~
=.�=�=�=9�=uY =���<�<��<H�<��<;�<4t�<[��<��<JP�<��<p��<�>�<���<IZ�<�.�<93�<�W�<���<H��<�o�<1
�<�[�<�k�<LK�<��<�΃<Z3}<,�r<�i<˚_<J�V<�N<S�E<e/><2�6<C�/<
q(<2!<ql<�A<:�<��;���;{�;G)�;��;�J�;}��;�xt;�O;fY*;e;�ÿ:X�l:+��9�0-�/��ۖ�M�Ժ�	��?*���L�Y�p�����fɟ�-L����Ȼy�ܻEp�1s�z
�������J�$�$���)�s�-���1�7;5�y�8��l<�U@�l|D��H��M��@Q�>U��aX��P[���]�7`�W[b��dd��Wf��*h���i�+5k�Tl�.m�]�m��n���o���p���r��ru���x��|������ ���4������(ꇼBꈼ�����7������JԊ�����8��������I�^������l!���ے�唔��6�����G��7d������
Ҝ����+1���R���_���O��T��Wϣ�s���#�����z���x��$'�����3+���Q���o��s���L�����V��7|���b��������_����Z���  �  �gO=�O=ƹN=7;N=?�M=�L=��K=9�J=T J=0	I=H=�BG=�xF=L�E=GE=��D=<	D=Y�C=�>C=��B=�B=qB=P)B=}�A=IQA=�@=��?=C?=�+>=<==�S<=�x;=`�:=��9=�Q9="�8=eA8=��7=}7=
67=c�6=!�6=�6=9o6="6=y�5=H%5=�s4=��3=��2=��1=�1=�L0=��/=��.=:F.=0�-=�5-=��,=W,=��+= �+=f9+=��*=�A*=��)=8�(=u�'=m)&='�$=��"=!=r0=�9=+6=X(=�=��=o�=m�=z�=\�=�
=��=�=��=��=>� =�\�<�z�<mj�<�?�<��<���<���<E��<���<��<�\�<���<�c�<�%�<��<*�<V]�<���<���<J��<���<j�<�T�<q�<*t�<�q�<�v�<E<~^u<]�k<^~b<?`Y<G�P<L�G<��?<W�7<s00<��(<�P!<	�<6�<�,	<�% <�J�;���;���;�X�;�L�;8v�;��k;|]E;_�;���:/U�:qdR:Q�9��L�d5/�s����Ѻ
L�pb)��lL�qjq�/ ���ğ�f���$5ǻlFڻ`���;��Dq�>A�����)�-#�\�(��F-�u1��85�"�8��R<�"@���C��)H�׀L���P�1U�[�X��s\��_�P`b�M�d���f��h���i���j�~�k��[l�S�l��:m���m�e�n���p�ߵr��hu�ւx�n�{�e/�6������!���g������
���&r��3��cӉ�?V��q���E!��������d׌�����s4���ɐ�~����l��I�����FÙ��R��.������3��D9��o��ޡ������������q���Ϥ�����7j���#�� �������ﯼ̱�Ɗ���'��i���9����)��(8��#���뻼̕��)���  �  EO=!�N=�N=�N=8�M=G�L=��K=-�J=>�I='�H=m�G=�F=%�E=RE=�lD=��C=NxC=)C=��B=��B=�B=\kB='B=��A=A=A=��@=g�?=��>=�>=e5==�n<=�;=;=|:=~�9=i\9=�8=UK8=q�7=�a7=�7=��6=�~6=�C6=#�5=��5=�5=Pp4=M�3=2�2=��1=-�0=�/=�/=�E.=��-=�	-=H�,=;,= �+=ϳ+=�v+=�.+=%�*=DD*=t�)=�(=�f'=a&=�$=|�"=�'!=�e=��=��=��=2�=��=<w=�A=�=��=p�
=�=��=��=˞=Mx =�a�<+��<�r�<)�<��<	W�<���<���<��<��<���<J��<KX�<�[�<A��<�۴<�5�<À�<��<琥<w=�<ή�<��<�"�<RQ�<��<��<�F�<�fw<�Bn<-e<��[<ϱR<�I<��@<UO8</0<f(<�� <4<�V<�	<�$ <Z�;�b�;X��;���;f�;[n�;{�a;Y:;%�;9�:~'�:,x1:��R9<Ȇ���8��F����Ӻ��	�Ł+��KO� �t�����Y������ƻ�oػ���9��� �����S�!b���!���'�S8-��1��5���9� �<�[z@��6D�R@H���L�DQ�	�U���Y��^���a��d��g���i��k��l��l���l���l�7m��Gm�b�m�`!o��p��Is��v��"y��5|�!�瀼����=��#M��'U��<\���a���]��&H����9Ȋ��Z���݋�:j��s�����hF��	ΐ�Ԙ��!���נ����������n��"
��	j��D���#l�����$�������GG������-!���٤�'ۥ��(��?����z��2P�����*ү�bc��_ղ�0/���y������k���.9��{e��Kz��)p��C���  �  ��N=ݜN=R?N=W�M=�LM=�L=��K==�J=@�I=ӃH=:[G=#AF=�AE=VfD=j�C=t4C=��B=B�B=7�B=�xB=�eB=�@B=��A=��A=��@=�F@=�u?=�>=��==�==5i<=��;=_;=�:=�g:=��9=�E9=̤8=?8=n7=��6=�6=|26=X�5=�5=YW5=��4=�C4=m|3=7�2=R�1=V0=|u/=�|.=��-=\�,=.V,=w�+=�+=�{+=�Z+=�7+=�+=#�*=p*=�X)=�W(=O '=޼%=<$=�"=�!=8z=f�=�=�F=O=/2=;�=��=7C=��=��
=3~=�k=�f=�^=�C =��<�H�<�.�<���<�>�<���<���<e~�<�5�<Z6�<.��<�8�<�2�<�m�<�շ<�R�<Cɰ<��<m7�<�<���<��<$F�<�<��<`m�<[�<�ɀ<Q�x<WAp<�?g<��]<�kT<W�J<�fA<IH8<��/<du'<�<�<�T<�2<\��;�(�;�;K��;` �;"�;��;�3W;#F.;Բ;���:�Є:-:)��8�ȳ��$J������ںo��T.0�ѱT�L�z�(w��W^��,�����ƻ��׻z绵��Y;���
�����+!��'�d�-�9�2��7���:�?>�L�A��E���H��=M��Q�A�V��X[��_���c�|g�Rj�dl���m�l[n��~n�vLn�9�m���m��m�מn���o�a�q�L�t�6dw�jYz��#}�H��p׀����U����h��T���^��쇆�����z���������ۋ��}��6��㴍����<���#���쒼:���
/��Oo��˝������{c���ՠ��˱���,��
r��4���[���u���[s��T6���N�����\��o ��s⬼��������8��nZ��kn�����������	���q��⹼�F������H����  �  ��N=y4N=q�M=IsM=�L=�UL= �K=نJ=�cI=*H=��F=��E=��D=�C=C=W�B=vFB=�%B=�B=\#B=�B=< B=غA=�GA=,�@=T�?=?=5>=6q==��<=�L<=��;=�;=3;=��:=�?:=8�9=d�8=28=vb7=m�6=�46=^�5=��5=�E5=.�4=1�4=!�3= <3=/N2=Q?1=�0=��.=��-=� -===,=��+=�N+=�+=�+=��*=�*=��*=Ek*=��)=b)=�(=��&=uZ%=��#=�c"=o� =u=��=�a=ѧ=ݽ=��=�Q=w�=#_=��=<z
=u4=�==�=o��<Q��<��<��<�M�<���<���< �<�U�<���<���<�2�<���<}�<[{�<y�<.��<6�<���<���<�Z�<�ן<�(�<�m�<qɑ<W�<k�<h�<��<w"z<��q<�h<܃_<r�U<��K<ޔA<]�7<<�.<�'&<�0<�<��<��<���;70�;��;��;��;�E�;&y;mM;�;#;���:7l�:��`:��9��ѷB]��>_�l.����{��O6��|[��ڀ��铻^W��ּ��KȻ�[׻�"�C�������m	��>�r��� �C�'��w.�4�|�8�%�<��?��C��eF��J��EN���R���W�:�\�[�a��-f��i�*�l�Ao��9p�Ûp�gp���o��;o�P�n�,�n��o�T5q�-hs�[v��y���{�=h~�s4��J�������*��꿂�Đ�������腼b\��݈��J������Z���TI���㍼�}���=���E��é���m��9���W֗�g?������ɞ�5���,��"?���飼b>��BV��YQ���S��?�������.ƥ������v���,��[�����D��;G���>����沼�ӳ�����}Q��:㷼����9D��ռ�?-���  �  �DN=��M=�nM=FM=a�L=�	L=~@K=�CJ=3I=��G=A�F=yHE=$&D=�3C=�|B=�B=�A==�A=��A=	�A=��A=y�A=�tA=B�@=N@=`�?=أ>=v�==c==��<=.'<=��;=�;=�e;=�;=s�:=��9=T9=�(8=fK7=�6=��5=:o5=�5=�4=w�4=Q>4=*�3=��2=�
2=%�0=3�/=��.=@x-=�{,=��+=�+=��*=*�*=��*=ۢ*=|�*=�~*=�**=ڗ)=y�(=��'=~`&=��$=Ä#=�"=� =kb=�=̍=��=�
=��=|�=�=h=��=6D
=��=ֵ=ŧ=��=�A�<���<O�<�>�<���<j	�<q�<()�<X[�<���<���<�<���<�"�<N��<\�<Y�<֤�<���<���<覣<0�<iT�<֚�<�
�<���<p��<g�<�<�<��z<��r<j<��`<ہV<�L<��A<KK7<\�-<��$<��<�<�y<��<��;��;���;�G�;�y�;��;U�q;��D;!;���:�:��>:���9� �	�)(s�㳱����8��SX<��b�7L���?���B����xKɻ��׻�h�hB�� ��f��\�p��(� �"`(��W/�_S5�T=:�s2>���A�܏D�X�G��AK��WO�g�S�;Y��=^�[c��h�3l��1o�.Gq�Ur�9�r��r�f<q��ip���o���o���p�d|r���t���w�%�z��q}�
��|����,������ׁ��N��V
��7��g��"���߈�����	���5�����Ĵ��WE����}䐼�6��L󓼍��Tr��f���u��������`H��SW��Q祿�&���������#䤼_���}��+\�������6���������3\��K���Φ���^����x����X��`l��Ե������l���\���-�������  �   N= �M=#M=\�L=�aL=��K=�K=LJ=[�H=��G=PHF=��D=��C=q�B=�B=��A=�sA=$mA=,�A=��A=��A=��A=lAA=��@=�@=8?=�W>=��==g�<=YX<=�<=V�;=$�;=b�;=�,;=b�:=i�9=9=�)8=�67=�Z6=��5=�'5=c�4=~�4=�W4=4=H3=N�2=��1=��0=��/=�R.=g(-=�",=]R+=K�*=qo*=�Q*=SV*=.g*=�l*=O*=i�)=�d)=׆(=�h'=�&=$�$=&@#=Z�!=֑ =6P=	=J�=m=�7=�=�=@=4h=��=G
=��=�p=�_=�c=&��<���<���<���<�k�<2��<���<ח�<ʳ�<��<n��<�T�<?4�<߁�<5�<�<Y��<I=�<l��<�<9%�<?��<ݺ�<u�<0�<`P�<�u�<�ׄ<(L�<.F{<�ds<v�j<�7a<�V<	:L<�_A<��6<��,<6�#<N�<��<�g<��< ��;��;�m�;^��;N��;h��;,�l;��>;��;L�:_�:Y(:��\9"�G��W�ۋ���y��D���3c��@�s�f��ǆ�i���	e�������Mʻs�׻��l�"A ��������?��� �x�(�90��F6�`;��g?���B�˥E�:�H��L�� P�~�T�B�Y�@._��qd�Pi��xm�q�p���r�F�s���s��%s�^/r��>q���p���p���q��ls���u���x���{�8�~�!T��( ��[��Y������K������σ��D������눼�Ɗ�*j��&���򦎼�M��0׏��v��OY�����U���r��iߘ��t�����fi��ts��������
���¥����xl���J���g��7⥼�ʦ�����©�ݑ���X��o箼1��� ~���豼a��8����������U��]��0w���t��5+���  �  �zK=9K=��J=U�J=�J=UkJ=8�I=��H=��G=�hF==�D=JrC=b B=�A=P@=��?=��?=Q�?=�7@=hz@=I�@=́@=�@=�a?=�g>=�F==`%<=B,;=�w:=:=��9=�:=�<:=iS:=�/:=p�9=��8=��7={�6=�b5=P4=T3=�2=>�2=0�2=,�2=��2=�2=�2=G1=�*0=z�.=$�-=09,=�+= D*=��)=��)=��)=��)=�'*=F_*=�`*=�*=oc)=bV(=�&=�l%=��#=�N"=D� =��=��=��=V�=:=�r=N9=��=�=Ԅ=�p=�=#�=R�=J�=Y��<�]�<���<�}�<���<2<�<�=�<i��<�q�<�#�<55�<=��<T�<�	�<&��<�]�<_�<J�<2�<N	�<���<���<���<�A�<}1�<���<J��<�
�<��<��{<��u<��n<�,f<f=\<�Q<��D<t�8<2-<I"<�<��<�	<E�<�'�;���;�7�;���;��;K�;6݀;T O;�6;w{�:���:��:S��8����|5�Za���8��g����TkA���j�Q銻����ܴ��ǻ|�ֻQ{��g�s���{��E
����մ��?$�.��[7��?�*|F�+�K��%O�jQ�US���T�s�V�[ Z��)^��8c�^�h�0�n�Z�s�z]x�֩{���}��~��j}�8�{��"z��x�7�w��w��y���{�cH���������������iz��UX���煼�p��UD�����;���!|��2���%;������॑�"������Z���^���^��'���uu���䖼���� ����b���K�������B��	5�~G���������R�����{ǧ�j����������˭�d)��T������!���������x|���]������&}��m���=��Gּ�8����	¼|ļ�  �  ��K=�6K=K=��J=w�J=��J=��I=I=��G=$F=nE=Z�C=FB=�7A=�y@=�@=��?=B@=�Q@=�@=��@=`�@=�/@=4|?=�>=k==�M<=�U;=x�:=6:=>:=>":=(C:=�P:=�':=��9=��8=��7=�6=z5=�o4=b�3='3=3�2=u�2=� 3=��2=��2=�12=8Z1=�>0=A�.=B�-=�[,=�B+=m*=��)=��)=��)=p�)=�?*=xs*=ds*=?%*=�y)=cq(=�'=`�%=��#=Kv"=�!=%�=��=��=��=52=�f=-=��=D�=��=��=�==A�=Q�=l
 =���<���<���<���<Z]�<�c�<��<ͭ�<:k�<��<y)�<�p�<�Y�<�˹<���<Ò�<xx�<z�<U:�<Iۤ<��<�՚<���<)��<��<�؇<�I�<��<J|<��u<�n<hf<5\<��P<�E<s�8<�i-<��"<dr<�i<tr
<b<�;t��;l��;�p�;���;���;洁;�7Q;=� ; ��:�r�:�:��9O���|-�h!��%:��b�'e�I}?�6Lh�V���J"���s����Ż�ջ<��*�ﻴ]��Ѭ��]
��H��3$���-�o�6��&?�*�E�o�J�vN���P�!R��6T�o~V�_�Y�+�]���b�@uh��n��Ss�:�w�v{���|�Qx}���|��z{��y�/x�gBw�D^w�=�x��E{���~�E[��B���̄��̅� 9��(��I̅�_j���M��M���qʆ������������Bj��Ra��:Ӓ�����	�������Wr��aH��8���Θ�g[��30����T���������X���7���zڨ�l���駼/������ @��g��:P������,ۯ���������״��f�������h��i]������
���C��%?���ļ�ob�������ü�  �  �L=ҩK=stK=�TK=�&K=~�J=E+J=[BI=�H=ھF=XSE=��C=2�B=f�A=��@=7�@=#^@=Sn@=-�@=1�@=��@==�@=�l@=�?=��>=�==ƽ<=��;=V;=��:==\:=�N:=�Q:=TF:=::=�9=�8=/�7=��6=Ͷ5=��4=	4= �3=�d3=�\3=7_3=�H3=~�2=�i2=%�1=x0=(;/=.�-=��,=��+=��*=�\*=�!*=�#*=VM*=R�*=�*=��*=�Z*=��)=��(=�s'=+�%=0g$=y�"=-!=�< =�=��=6�=�=�A=x	=�v=��=��=e�=P�=�t=�6=�:=i =8�<�_�<��<91�<%��<X��<Y��<�Z�<�7�<fi�<*�<D_�<�:�<F��<�E�<�!�<_��<���<Ի�<�q�<��<���<�z�<�w�<~ӌ<.��<�<���<�y|<w�u<>n<�{e<�[<I�P<�CE<H�9<��.<"9$<=<<\<ny<9u�;��;���;;�;�7�; ��;�.�;�:W;��';B��:	�:�;:7w9~�F��\��i|��0��d`�c��TX:�wBb��1��Oc�������"»3�һ��@����� ���
�w���!$��L-��6�y�=��7D�N+I���L�_O�� Q���R��sU�G�X��]���a��bg�l�l���q��v��.y��{��{�ZM{��&z�D�x��Fw��mv�r�v���w�z��P}����A^���烼y���񆅼7��������_��\o��v����@��������Ȍ�2ގ�-��������ɒ�$(��!F���k���ݓ��̔��P���b��O㚼n���U\��u碼������ʲ��x"��@���̧�Pg���"���6���̧����������¬�j ��y��vղ����ô�����7���c��[ص�ɶ��I���J��q�������1��uü�  �  ^�L=NL=L=��K=��K=s*K=�zJ=��I=4dH=>G=4�E=y{D=VPC=�WB=�A=S-A=K�@=��@=�	A=f%A=L0A=A=ھ@=�)@=!Z?==b>=^==m<=��;=�;=;�:=\�:=\:=|+:=��9=o]9=��8=��7=��6=�6=;5=a�4=U:4=�4=A�3=��3=�3=�U3=��2=U�1=��0=H�/=�n.=�O-=�T,=�+=`+=��*=�*=g�*=J�*=;�*=��*=�*=2*=#)=��'=��&=~%=w}#=�	"=C� =�X=H =��=Y�=��=Q�=�I=
�=��=�=�l	=��=}�=��=�� =f�<��<��<���<LC�<Ft�<n�<�[�<�h�<���<[�<8��<K��<꽻<>B�<��<¤�<�/�<�k�<!@�<�<=ɜ<���<K˒<��<�ŉ<�ʅ<A�<��|<tWu<�Rm<N�d<��Z<8LP<:eE<oz:<��/<w-&<3Y<!}<`]<v�<�s <�\�;��;�-�;���;n��;m܇;U4`;%�1;\J;/i�:D�h:���9/vJ�Dd򹢄b��򦺶f�>���33�ĿY��J����W3�� ��=λz�ݻ�`�^I��� ��o��B�����3$���,�|�4�<�;�1�A���F�mJ��L���N��3Q�GT�̔W���[�<�`���e���j��}o��qs��qv�@Vx�! y�w�x��/x�@w�:�u��Ju�Uu��Wv�W_x�
E{�#�~����!����Ѓ�j���a���9��%f������I[��/g���؈�U���g��'��Y���Eɐ������呼����o������$�����8ϗ��6��Ȝ�wV��e�������N��LX��o়����ᦼ���B��������0��?;���é�%���#ȭ�Jӯ�l������t과s����������t1���7��/����q��:s��U}��p`��=����  �  9WM=?�L=�L=muL=�L=
�K=��J=K�I=��H=>~G=sGF=#E=1D=#C=pB=��A=�A=ʍA=��A=v�A=#yA=�VA=NA=��@=��?=��>=
>=�==�I<=n�;=�;=��:='Q:=��9=�9=�9=�f8=��7=	�6=0I6=u�5=�65=@�4=R�4=?�4=ao4=K%4=��3=��2=22=�1=�
0=L�.=u�-=�-=�],=j�+=�+=�b+=�V+=�U+=.N+=�-+=��*=xX*=�)=pq(= '=ߧ%=�$=+�"=9!=̔=.=�a=%�=��=`=��=Nu=��=�P=��	=Z�==j=�k=N|=��<���<�*�<=$�<���<�<�Q�<x��<���<&O�<C'�<ih�<��<��<na�<sյ<�Y�<{ή<��<�
�<���<#��<�<u8�<�t�<�<���<�~�<y�|<y�t<�l<��b<,_Y<�_O<2-E<;<L1<'%(<q�<<~�<Z�	<=.<��;���;"*�;��;��;y�;(�j;5;>;л;�-�:mh�:Ƹ:˭�8�����cF��n��,�պ�	
�� ,�[�P��x�bB���W��������ɻ��ڻ���Vj�����S��ȑ���m�$��g,�$�3�:��}?�?�C�LMG��J��L�CpO��R�xV���Z�sg_��d�/�h�t�l�vhp�&6s�#u�$v�Dv���u��Qu���t�M6t�Ct�*u�5�v��%y�_/|�Ou��H��3���o����n����˛��]=��t
������N�����L"���|��ץ��l���K$��󊐼j琼�l��E��(����7��@��f����ڛ�~)��[O���/������;����e��۹��إ��ݥ��ꥼ� ��j���s���|ڨ�?���z��s���E��-Ա�����������յ��ȶ�n근�C���ͺ�s�����䖿������  �  ��M=ΓM=�FM=��L=�hL=��K='�J=�I=��H='�G=L�F=��E=y�D=��C=�FC=�B=�cB= B=�A=��A=n�A=�vA=�1A=y�@=�3@=�u?=��>=�==��<=�<=R;=��:=":=�9=D9=g�8=��7=�o7=+�6=�m6==6=d�5=�w5=�K5=j5=��4=�n4==�3=3=
?2=`S1=/d0=�z/=R�.=$�-=�0-=d�,=N,=,=��+=�+=��+=0O+=��*=�~*=��)=��(=И'=Q0&=�$=E	#=�a!=��=��=�=�=�=(�=�=i*=	�=ep=�)
= �=Q�=��=��=��<�)�<)a�<UL�<���<x��<��<ޙ�<�/�<���<f��<C�<���<l�<qj�<r��<hڲ<-�<Tr�<���<�c�<9�<TD�<Nq�<q��<�ڋ<�7�<��<�S|<�Es<�j<}�`<HVW<��M<�^D<�;<E"2<_�)<��!<�"<S�<�I<V<{�;���;��;rm�;�=�;uҏ;"�t;��J;�!;��:b[�:��K:�͐9�#V�`:/�E��NϺ�[��'��J�guo�P��E������0ƻ�ػ�j껥����;�<u��z�Z;�M�%�)�,��2�;�8��}=�b�A�O�D�T�G�N�J�s>N���Q���U��/Z��}^�+�b�H�f��3j�kUm��o�H�q�'�r���s���s��s�D�s�i�s�|�s�	[t�K�u�Ӎw��$z�5&}��"��ם����������#����������
��w������!��b���ݍ�(�����mh��q폼2����ő�q7��b�������t��F��l잼������f��<飼�|���礼:�����]ݥ��\������9��۫��Of��H��)���갼����과7���s�������븼.��Cu��B�����S
�������  �  �;N=��M={�M=�M=�|L=�K=�J=`�I=��H=��G=�
G=B4F=�kE=ٲD=�D=~C= C=��B=94B=�A=��A=�\A=A=��@=�N@=z�?=��>=I>=�%==v<<=�\;=�:=��9=�9=�m8=��7=�e7=��6=�6=Ib6=�(6=>�5=��5=_�5=�e5=z5=�w4=;�3=@�2=B,2=�[1=��0=��/=y*/=�.=��-=q-=8�,=c�,=�;,=��+=b�+=5:+=��*=/e*=��)=��(=��'=Q~&=K�$=�E#=Qz!=,�=k�=��=�q=�E=+=��=s�=ӄ=_=sE
=�8=5=.=�=��<D	�<��<��<��<���<���<q�<Ya�<a_�<at�<���<��<���<�-�<i��<���<7�<iX�<���<ӛ�<�j�</�<A:�<"X�<@d�<�m�<)z�<&{<hCq<��g<��]<ʩT<}�K<:�B<�^:<�22<�[*<��"<^<��<W�<�{<R��;`��;?E�;�]�;�i�;��;�D};�U;X�.;R;t:�:ƾx:�!�9���N�"�g���zϺǁ��&��9G���j�f.��2䛻����$Ļp�׻zd�A���8�a������y �2R'�/�-�3�88�UG<��@�lC���F�ZCJ��N��R�oQV��qZ�5T^���a��e�z h���j��l��n�''p��Vq�Gr���r��s�7�s�@0t�5�t���u���v��y�K�{�j�~����g����%�����������1��OS���N��%���݋�\}��B��y��G܍��>������Ao���q��lǑ�!d���-�����Ә�c���0��8����(��u��+��������w���=���뤼�����	��F���&8�����iI��@ʪ���� v��yf��hJ�����J̵�yf���⸼�:���h���p���Z���)��'߾�}���  �  �SN=�N=��M=LM=�EL=VbK=�nJ=_I=��H=��G='*G=@�F=��E=BQE=�D=ND=$xC=��B=�GB=��A=XA=tA=�@=�w@=M@=C�?=�>=b+>=�:==`9<=u3;=�3:=B9=g8=��7=o7=��6=�h6=�=6=�$6=�6=�6=��5=ݼ5= e5=��4=�64=Kp3= �2=��1=Z+1=i�0=�	0=�/=E/=ݖ.=&.=U�-=��,=�o,=d�+=�_+=&�*=�x*=*=�x)=!�(=��'=��&=�%=�E#=�Z!=�L=^$=.�=E�=�j=l;=�=�=E==�(
=v7=s<=�*=o�=�C�<UW�<�E�<�0�<	3�<*X�<X��<w��<BE�<���<h��<���<�#�<P�<���<��<���<I��<���<T��<�>�<�L�<��<Jx�<Ǔ�<�v�<#6�<��<�)y<��n<Ipd<�Z<ryQ<��H<ƭ@<a�8<�n1<?(*<@�"<.�<Y�<�g</{<�&�;���;�{�;(~�;��;���;K��;<z^;L^9;	�;���:O��:�:q��TL$�K�����׺ �t�)��I���j�,K������#�����û%�ػ�����7�
���� �A#�ƙ)�p$/� �3��88�(<�)�?�=C�e�F�,�J��O��qS�N�W��[�a_��a�{Sd��of��_h��<j�;l�K�m�޳o��kq���r��1t�Bu�Q�u��v���v��w�0y��m{��c~��瀼����T���~d����5���Pފ�oՋ���������6��c������6�������������*ɐ�H[��d���䕼@���D��Fq��׫���՜�����'���W������Ƣ���+���󥼣���"O���ߧ������{������-\��FC���X��t���c����������8[���Ȼ�T弼Y����P���þ�N��qu���  �  3N=D�M=�gM=�L=��K=Y�J=?�I=��H=3H=��G=�G=ǭF=�AF=��E=�5E=0�D=��C=W�B={,B=�vA=y�@=s@=�'@=�?=ʰ?=�T?=��>=�	>=�== <=��:=�9=Z�8=3�7=�6=5B6=��5=5�5=Ա5=)�5=��5=��5=-�5=�5=�#5=�4=&�3=1�2=�2=�W1=<�0=-^0=0=��/=hu/=\/=֑.=��-=�:-=Cv,=^�+=D�*=c*=��)=�k)=�(=QQ(=`v'=O&=�$=�#=�!=x�=��=>+=��=ɀ=�R=�F=X=F}=a�=v�	=� =	=��=�=9O�<�.�<E�<`��<�,�<���<�N�<��<���<�p�<���<G��<��<6��<��<���<�<Җ�<���<���<c�<W��<��<y8�<�[�<@!�<�<��<��v<�k<)a<&W<iN<2�E<)><n�6<� 0<�0)<72"<��<�<=�	<�� <���;��;��;��;d�;qc�;�;\�d;7�A;��;^�:��:��:�ꥸ�G2�M���D�,��0�3�N��}n��q���L�������;Ż�Vۻ�p�q{�A��v��D��U&�E,��@1��y5�)9��<���?���C���G��+L��P�ŮU�Z�ǰ]��`��b�Dd���e���f�JHh�xj��Il���n�_Gq�Y�s�k�u��w�v�w�*Xx��x�Ay�0z�5|���~�M4���6���V���s��Jn���)��z����|��H���9��V4�������������I�������[���4h��YF���������ݽ�����$����F��X ��!'���f��ڠ�<n�����e���ɦ��ŧ��y������[~���.���5����������m������񁵼d᷼��:���+v�������*������ܦ��C���"ӿ��  �  ��M=j�M=�	M=�8L=n;K=�+J=$)I=*NH=5�G=�5G=��F=r�F=�qF=7F=��E=v�D=��C=��B=9�A=|
A=HO@={�?=�w?=�H?=T!?=w�>=�p>=��==��<=ص;=�w:=l29=��7=��6=6=`r5=W5=�5=5=K5=�{5=�5=��5=D5=�4=��3=�3=A02=�]1=!�0=^J0=h0=�/=a�/=��/=g/=��.=�1.=XQ-={Z,=�c+=�*=��)=�-)=j�(=�I(=��'= '=��%=Ն$=�"=�� =([=��=7l=��=�==s=]t=O�=<�=�0={	=��=��=Ǆ=O=�<���<\��<$��<���<��<���<���<��<2�<Z��<(��<d�<��<BU�<��<�<'e�<jY�<U��<�C�<���<��<Ϊ�<vܐ<���<��<��<0Et<o�h<��]<��S<��J<��B<&b;<�4<rG.<��'<9� <�n<c<��<�&�;��;Bj�;���;���;D��;g	�;�U�;�<h;�hG;�0#;��:Y:�:3x:���ՎH�����@����Vg:�V�V���t�!ڊ��1�������tǻ;Z޻�q��������%�r"�%])�[�.�{�3��<7�,{:��=�e�@�0�D�%8I��+N� \S��\X�ܹ\�@$`���b���c�"�d�]>e���e���f���h��Ek�z\n�\�q���t���w�V�y�[�z��{��{�,/{���{��`}���<���Nー3:��F����ˊ�㲌�9(���������B����H���莼엎�o���IՎ�2�������6���\�������"]������矚��7�������������u�����p���]���\���=���֧�����٩�0T������(��/����>��{���D���γ��y�����(���牽�������������Х��6z���i���  �  ��M=rMM=��L=r�K=��J=K�I=ׄH=N�G=� G=C�F=ѬF=3�F=U�F=�FF=��E=��D=w�C=��B=��A=ʛ@=��?=�)?=��>=��>=F�>=1o>=^>=8u=={�<=Mg;=:=��8=Fm7=�F6=^^5=q�4=+v4=�o4=p�4=l�4=�&5=bO5=B5=O�4=�T4=�~3=l�2=v�1=J�0=�!0=��/=ڱ/=��/=��/=�/=њ/=k/=�S.=3Q-=�/,=.+={*=�+)=w�(=�(=�'=<'=��&=t�%=�3$=l"=�K =��=�^=�=�C=d�=k�=1�=��=6Z=��
=@	=;X=�[=Y=s� =��<���<J9�<�B�<��<L��<)&�<���<E+�<�W�<p�<K�<��<���<x��<�A�<���<�>�< �<΃�<O0�<C؜<�3�<N�<HO�<���<�2�<�M~<�r<`:f<�[<��P<�G<x@<9<t�2<޳,</{&<ղ<�<n<l�<Α�;�;�8�;N�;A��;�ٝ;�F�;���;Qj;~�J;X';U��:���:�X:�4�%�`���º�E���&�KeC��^�wo{��{��`��;���u�ɻ�.�P���#��
�c���$%���+��L1�`{5�q�8�{�;���>�t
B��F�i�J�EP�E�U�*�Z�)A_��{b��td�TUe�te�/Ie��Xe��f�o�g��j�Wn�Rr��,v��uy���{��3}��}��m}��5}�.�}��~�/���Q�����o��+���(���Y ��S����u���ΐ�����;��1����7������m��6\��Jڑ�tœ��㕼�염ƞ���Қ�����Λ��ݛ��@������_���>���v���̤�����ߨ�BC���!�������Ϋ�O������᭼�����ڱ�J����W��U&������O߾�Pw���q��`�����������0������  �  !sM=JM=�aL=ElK=�IJ=ZI=�H=�AG=�F=�F=J{F=��F=X�F=�^F=��E=�E=)�C=�B=�qA=�H@=�[?=޸>=�`>=�@>=�7>=j>=��==�;==oX<=R/;=9�9=k8=S7=��5=��4=�L4=4=k	4=�C4=_�4=5�4=�5=}5=ڰ4=w	4=n$3=l2=I1=<G0=��/=�o/=+m/=�/=i�/=��/=y�/=�7/=*c.={I-=�
,=}�*=ȩ)=�(=�(=��'=�B'=��&=�A&=�P%=X�#=D1"=�
 =)�=�=�]=��=�e=A:=�L=�=��=xv
=�==�=��=�O =Z4�<���<�K�<\X�<���< �<ʬ�<�t�<y)�</��<�@�<2O�<��<s��< ��<S��<h@�<�j�<�A�<���<(l�<�/�<���<���<G�<3��<���<w}<�p<�d<2Y<E�N<}F<4G><?�7<�z1<g�+<�%<k�<�<@D< �<�_�;���;z��;�{�;���;���;�Ԏ;���;|�j;��L;X�);n� ;"�:�
:�?c��"s���κ����E-���I���d����s��
�����.`˻'��s���	����3����&���-���2��6�&�9�"�<�d?���B�9G���K��Q��>W��\�/	a��(d���e�ef��f�roe��e�;�e�rtg��wj�*rn���r�c2w�"�z��}�/�~��b�����~�J�~����]���x������@����?�����������r���_��쪑�Cp��J����3��n����}���ޏ�����wz��������� Ҙ����������/��E�������%��`Μ��-���+������[)��ۖ��8��� �����Js��}���ʬ�<N��Z����/G������^)ܺ������Ŀ�gc��eX¼>�¼��¼�"¼���Wo���  �  �_M=��L=aHL=�MK=&J=��H=*�G=�G=�F=(eF=�gF=}�F=��F=�eF=��E=E=}�C=Y�B=\A=b*@=S6?=�>=t7>=�>=�>=��==$�=='==;E<=E;=�9=�N8=m�6=��5=��4=#4=H�3=b�3=%4==�4=�4=�5=��4=�4=H�3=3==�1=��0=�0=O�/=�M/=gS/=K�/=��/=�/=��/=@/=Fg.=�E-=��+=g�*=&�)=��(=��'=�r'=�'=~�&=�$&=08%=�#="=��=A�=�=�7=�=�9=�=$=�p=*�= ]
=.�=�=�=ý=�1 =���<�\�</��<*�<Ԧ�<b��<
��<�]�<'�<���<T�<`�<��<\��<�~�<x��<��<�<u�<�[�<�#�<��<�r�<�k�<���<Ef�<���<O�|<�p<�c<h�X<�JN<�XE<8�=<�7<
1<D+<�8%<%y<�<)�<�<�D�;WK�;�U�;CC�;Zn�;m��;H�;&R�;k;zvM;�M*;Z/;�!�:��:Sjv�?z��Ӻ�J���/��(L�]�f�����5���������� ̻����U���"
�P�3=�o�'�L.��l3��J7��O:�q�<�)�?��)C�ZG�M_L��R���W��<]�D�a���d��jf�)�f�VMf��e��e���e�Rg�Bfj���n��s��w�}b{��~�!��������(�8#�/��i$���Ⴜ�(��nƇ�|������/���Ő�,���n���,�������b���я�:���������D����ǔ���$���Ӛ�G�n��6r��50��H��������������'�������M��iΧ��穼�o��~[��Nì�⬼~����������,��4n��y(���"������Խ�m��������¼@�¼��¼�X¼`��������  �  !sM=JM=�aL=ElK=�IJ=ZI=�H=�AG=�F=�F=J{F=��F=X�F=�^F=��E=�E=)�C=�B=�qA=�H@=�[?=޸>=�`>=�@>=�7>=j>=��==�;==oX<=R/;=9�9=k8=S7=��5=��4=�L4=4=j	4=�C4=_�4=5�4=�5=}5=ڰ4=w	4=n$3=l2=H1=<G0=��/=�o/=*m/=�/=g�/=��/=v�/=�7/='c.=wI-=
,=x�*=©)=��(=�(=��'=�B'=��&=�A&=Q%=q�#=m1"=�
 =��===?^=��=�f=�;=�N=.�=Y='y
=��=D= =J�=S =`;�<���<sR�<�^�<��<�<��<�w�<�+�<v��<'A�<sN�<C��<���<{��<Ա�<*;�<e�<7;�<ۤ�<Ge�<)�<ޠ�<D��<<ߏ<���<İ�<t}<Οp<Ʉd<�/Y<�N<vF<AK><C�7<p�1<�+<�%<��<<�Q<�<)|�;#��;ҳ�;^��;���;���;2�;Џ�;A�j;+�L;��);6� ;ĥ:K�	:cRe�f�s�WϺb�}-�gJ���d�V:������'���6��z˻�>�u�����	���W����&���-���2�,�6���9��<��?��B�G�O�K���Q�D?W�h�\�l	a�)d��e�.ef��f��oe��e�D�e�ytg��wj�.rn���r�e2w�#�z��}�0�~��b�����~�J�~����]���x������@����?�����������r���_��쪑�Cp��J����3��n����}���ޏ�����wz��������� Ҙ����������/��E�������%��`Μ��-���+������[)��ۖ��8��� �����Js��}���ʬ�<N��Z����/G������^)ܺ������Ŀ�gc��eX¼>�¼��¼�"¼���Wo���  �  ��M=rMM=��L=r�K=��J=K�I=ׄH=N�G=� G=C�F=ѬF=3�F=U�F=�FF=��E=��D=w�C=��B=��A=ʛ@=��?=�)?=��>=��>=F�>=1o>=^>=8u=={�<=Mg;=:=��8=Fm7=�F6=^^5=q�4=+v4=�o4=p�4=l�4=�&5=bO5=B5=N�4=�T4=�~3=k�2=u�1=I�0=�!0=�/=ر/=��/=��/=�/=̚/=e/=�S.=+Q-=�/,=$+=p*=�+)=l�(=�(=�'=<'=��&=��%=4$=�l"=4L =h�=�_=j�=�E=��=K�=��=�=�^=��
=�#	=U^=Zb=&==� =�
�<͘�<�E�<oN�<���<���<.�<��<�/�<oZ�<��<��<���<���<m�<69�<l�<n3�<��<�v�<
#�<�ʜ<�&�<��<�C�<7�<�)�<`>~<�r<2f< [<A�P<��G<B@<�"9<��2<-�,<G�&<A�<�'<��<�<<��;@<�;Tk�;{"�;���;���;�d�;��;�1j;K;yV';���:�`�:0�:�8�F�a���ú����&��C� \_�C�{�I���"����ĳ���ɻ�\�-��X6���)��0%�E�+��T1��5�G�8�D�;���>��B�mF���J�J P��U���Z��A_�|b�ud��Ue�Gte�MIe��Xe��f�|�g��j�Wn�Rr��,v��uy���{��3}��}��m}��5}�/�}��~�/���Q�����o��+���(���Y ��S����u���ΐ�����;��1����7������m��6\��Jڑ�tœ��㕼�염ƞ���Қ�����Λ��ݛ��@������_���>���v���̤�����ߨ�BC���!�������Ϋ�O������᭼�����ڱ�J����W��U&������O߾�Pw���q��`�����������0������  �  ��M=j�M=�	M=�8L=n;K=�+J=$)I=*NH=5�G=�5G=��F=r�F=�qF=7F=��E=v�D=��C=��B=9�A=|
A=HO@={�?=�w?=�H?=T!?=w�>=�p>=��==��<=ص;=�w:=l29=��7=��6=6=`r5=W5=�5=5=K5=�{5=�5=��5=D5=�4=��3=�3=@02=�]1=�0=\J0=f0=�/=]�/=��/=g/=��.=�1.=MQ-=oZ,=�c+=�*=u�)=�-)=\�(=�I(=��'='=��%=�$=y�"=R� =.\=]�=+n=�=c�=Kw=?y=�=��=78=
�	=L�=ͼ=5�=�(=+0�<��<J��<��<)�<@��<���<���<!�<��<��<��<R_�<���<LK�<��<��<+U�<H�<��<B1�<��<eߙ<%��<�ː<���<�م<�<94t<��h<n�]<%�S<�J<��B<zr;<T�4<Ia.<[�'<R!<��<�4<K<�s�;�`�;���;d�;���;*�;�3�;v�;%hh;G}G;o.#;Y~�:nڠ:�`:U���DJ�T��GY�����;��W��u��+�����{ϱ�X�ǻ\�޻{�����Ѩ��8�P�"��j)�?/�0�3�dC7���:��=���@���D�:I�q-N�<]S�|]X���\��$`���b�"�c�Z�d��>e���e���f���h��Ek��\n�e�q���t�Íw�Z�y�^�z��{��{�-/{���{��`}�	��<���Nー3:��F����ˊ�㲌�9(���������B����H���莼엎�o���IՎ�2�������6���\�������"]������矚��7�������������u�����p���]���\���=���֧�����٩�0T������(��/����>��{���D���γ��y�����(���牽�������������Х��6z���i���  �  3N=D�M=�gM=�L=��K=Y�J=?�I=��H=3H=��G=�G=ǭF=�AF=��E=�5E=0�D=��C=W�B={,B=�vA=y�@=s@=�'@=�?=ʰ?=�T?=��>=�	>=�== <=��:=�9=Z�8=2�7=�6=5B6=��5=4�5=ӱ5=)�5=��5=��5=-�5=�5=�#5=�4=%�3=/�2=�2=�W1=9�0=)^0=0=��/=bu/=U/=̑.=��-=�:-=4v,=M�+=1�*=�b*=��)=~k)=�(=RQ(=rv'=5O&=g�$=�#=e!=��=��=�-=�=˄=�W=�L=_=F�=T�=F�	=P=7=�=��=�f�<�E�<0�<��<�?�<��<c\�<��<6��<�t�<���<���<2��<��<ъ�<���<�ױ<H��<b��<g�<,L�<W��<���<�"�<�G�<��<���<r��</�v<��k<�a<�%W<�N<��E<$><y�6<� 0<U)<�Z"<o�<��</
<�� <}��;�[�;�d�;�W�;�,�;���;�(�;[�d;��A;��;��:;��:H�:�ȳ��_4��G�����#����1�m�O��Go�WՈ�l�����=�Ż)�ۻ��a����<��X�f&�vR,��K1�[�5��/9�3�<���?���C�Q�G�Q-L�~�P�ѯU��Z�c�]�j�`�J�b�XDd��e���f�hHh��j��Il���n�jGq�a�s�q�u��w�z�w�-Xx��x�By�0z�6|���~�M4���6���V���s��Jn���)��z����|��H���9��V4�������������I�������[���4h��YF���������ݽ�����$����F��X ��!'���f��ڠ�<n�����e���ɦ��ŧ��y������[~���.���5����������m������񁵼d᷼��:���+v�������*������ܦ��C���"ӿ��  �  �SN=�N=��M=LM=�EL=VbK=�nJ=_I=��H=��G='*G=@�F=��E=BQE=�D=ND=$xC=��B=�GB=��A=XA=tA=�@=�w@=M@=C�?=�>=b+>=�:==`9<=u3;=�3:=B9=g8=��7=o7=��6=�h6=�=6=�$6=�6=�6=��5=ܼ5=�d5=��4=�64=Jp3=�2=��1=W+1=f�0=�	0=��/=>/=Ԗ.=.=H�-=��,=�o,=Q�+=�_+=�*=�x*=�*=�x)=#�(=�'=�&=D%=qF#=�[!=2N=[&=��=ʫ=o=�@=W%=�=-=$=�3
=8C=�H=�7=�=�]�<�p�<*^�<cG�<�G�<Xj�<���<x��<�M�<���<i��<	��<I�<�E�<c��<��<��<�y�<��<�<\%�<23�<���<3`�<K}�<-b�<V$�<�ց<�y<�n<�gd<[�Z<��Q<��H<��@<^9<��1<�P*<b#<Թ<i�<I�<��<���;^2�;G��;�ϸ;f4�;��;���;y�^;�z9;�;o��:�y�:N:�誸ѡ&�3P���rٺ��=m*��I��fk�g������a��GHĻ�Uٻ+�W8�,�
����7��S#���)�w0/��4� @8��<���?��C�
�F�0�J�/O��rS�3�W���[��_���a��Sd��of��_h��<j�Ul�_�m��o��kq���r��1t�Gu�U�u��v���v��w�1y��m{��c~��瀼����T���~d����5���Pފ�oՋ���������6��c������6�������������*ɐ�H[��d���䕼@���D��Fq��׫���՜�����'���W������Ƣ���+���󥼣���"O���ߧ������{������-\��FC���X��t���c����������8[���Ȼ�T弼Y����P���þ�N��qu���  �  �;N=��M={�M=�M=�|L=�K=�J=`�I=��H=��G=�
G=B4F=�kE=ٲD=�D=~C= C=��B=94B=�A=��A=�\A=A=��@=�N@=z�?=��>=I>=�%==v<<=�\;=�:=��9=�9=�m8=��7=�e7=��6=�6=Ib6=�(6=>�5=��5=_�5=�e5=y5=�w4=9�3=>�2=?,2=�[1=��0=��/=s*/=�.=��-=q-=+�,=T�,=�;,=��+=M�+=:+=��*=e*=��)=��(=��'=�~&=��$=�F#=U{!=��=~�=��=4u=J=�=s�=}�=�=Si=�P
=(E=�A=g;=m"=���<�#�<-2�<��<���<���<ę�<�}�<(j�<]d�<lu�<���<� �<a}�<��<�<d�<��<	@�<t�<i��<LP�<&ؚ<P!�<�@�<*O�<[�<�j�<]�z<	3q<g<a�]<9�T<ͯK<�B<�|:<W2<��*<W�"<i�<�<{"<%�<2Y�;[O�;��;#��;;'��;Ԡ};��U;٢.;;a��:Эw:�9�F��^%��ʒ�Ѻ�V���&�{ H�a�k������S���o����Ļ9Yػ\�뻌����X�������� ��a'���-��"3�	8�gM<��	@��oC�_�F�uEJ�aN�6R�_RV�irZ��T^�8�a��e�� h���j�&�l��n�<'p��Vq�*Gr���r��s�<�s�D0t�8�t���u���v��y�L�{�k�~����h����%�����������1��OS���N��%���݋�\}��B��y��G܍��>������Ao���q��lǑ�!d���-�����Ә�c���0��8����(��u��+��������w���=���뤼�����	��F���&8�����iI��@ʪ���� v��yf��hJ�����J̵�yf���⸼�:���h���p���Z���)��'߾�}���  �  ��M=ΓM=�FM=��L=�hL=��K='�J=�I=��H='�G=L�F=��E=y�D=��C=�FC=�B=�cB= B=�A=��A=n�A=�vA=�1A=y�@=�3@=�u?=��>=�==��<=�<=R;=��:=":=�9=D9=g�8=��7=�o7=+�6=�m6==6=d�5=�w5=�K5=i5=��4=�n4=;�3=3=?2=]S1=+d0=�z/=L�.=�-=�0-=Y�,=N,=,=��+=��+=��+=O+=��*=�~*=��)=��(=�'=�0&=h�$=�	#=�b!=��=��=z=�==��=��=+2=��=\z=q4
=�=��=i�=�="��<)C�<�y�<c�<_�<���<%$�<��<p8�<���<i��<m�<
��<�a�<�\�<���<�Ʋ<U�<�Z�<&s�<VJ�<�ٞ<*+�<1Y�<���<�Ƌ<&�<4��<�<|<�5s<oj<��`<o]W<��M<�tD<�2;<lE2<��)<��!<pS<j�<~<g�<X��;LG�;jr�;��;F��;��;D3u;�J;��!;��:��:0�J:u͍9��]�R�1�㜔��к�)���'���J�jVp�Z���"����l���ƻ��ػ��껎���{Z��������M�Z�%�H�,��3�Э8�~�=��A���D��G�\�J�@N���Q���U��0Z��~^���b���f�4j��Um���o�b�q�;�r�Йs���s�%�s�J�s�n�s���s�[t�M�u�Սw��$z�6&}��"��ם����������#����������
��w������!��b���ݍ�(�����mh��q폼2����ő�q7��b�������t��F��l잼������f��<飼�|���礼:�����]ݥ��\������9��۫��Of��H��)���갼����과7���s�������븼.��Cu��B�����S
�������  �  9WM=?�L=�L=muL=�L=
�K=��J=K�I=��H=>~G=sGF=#E=1D=#C=pB=��A=�A=ʍA=��A=v�A=#yA=�VA=NA=��@=��?=��>=
>=�==�I<=n�;=�;=��:='Q:=��9=�9=�9=�f8=��7=�6=0I6=t�5=�65=@�4=Q�4=?�4=`o4=I%4=��3=��2=02=�1=�
0=G�.=p�-=�-=�],=a�+=��+=�b+=�V+=�U+=N+=�-+=��*=iX*=�)=sq(=# '=�%=7 $=��"=!=�=�	=cd=Q�=��=�d=�=A|=��=vY=y�	=�=du=Uw=�=#�<���<�@�<�8�<!��<b+�<�_�<K��<}��<S�<,(�<�e�<��<��<+U�<kƵ<H�<���<���<���<���< �<x�<�"�<�`�<�ي<���<^q�<��|<[�t<^�k<�b<�eY<�lO<�@E<(;<l1<�I(<��<�3<\�<P�	<3]<ga�;`M�;e{�;8�;���;�<�;Q�j;�p>;��;(�:)�:��:��8 )���|H�a����׺a�
�c�,���Q���x�O�������-���* ʻۻ�)�ܩ���������������$��r,�ө3��:��?�_�C�xPG�J���L��qO��R��xV�x�Z��g_�d�v�h���l��hp�E6s�;u�6v�"Dv���u��Qu���t�R6t�Ct�,u�7�v��%y�`/|�Pu��H��3���o����n����˛��]=��t
������N�����L"���|��ץ��l���K$��󊐼j琼�l��E��(����7��@��f����ڛ�~)��[O���/������;����e��۹��إ��ݥ��ꥼ� ��j���s���|ڨ�?���z��s���E��-Ա�����������յ��ȶ�n근�C���ͺ�s�����䖿������  �  ^�L=NL=L=��K=��K=s*K=�zJ=��I=4dH=>G=4�E=y{D=VPC=�WB=�A=S-A=K�@=��@=�	A=f%A=L0A=A=ھ@=�)@=!Z?==b>=^==m<=��;=�;=;�:=\�:=\:=|+:=��9=o]9=��8=��7=��6=�6=;5=a�4=U:4=�4=A�3=��3=�3=�U3=��2=S�1=��0=E�/=�n.=�O-=�T,=�+=Y+=��*=�*=[�*=<�*=-�*=��*=ڡ*=&*=#)=��'=��&=�%=�}#=O
"=�� =�Y=�=��=��='=W�=�N=��=`�=�=�t	=9=��=j�=1� =�/�<�*�<���<Y��<zR�<���<Qy�<�d�<o�<$��<��< ��<h��<\��<48�<��<z��<��<=Z�<�-�<:��<k��<S��<���<[	�<���<x��<k�<.�|<�Ku<�Lm<�d<��Z<�VP<XuE<��:<Q0<FK&<^z<�<�<ݭ<@� <ק�;� �;�o�;�ζ;cȟ;S�;v`;$$2;�_;�d�:�Kh:iY�9�%\��=���;d�%狀�~�:����3�tcZ�g����\�������V��كλn#޻=��2}��T7�7���R����>$���,���4���;���A��F�J��L��N��4Q�*T�y�W�!�[���`��e��j�
~o�	rs��qv�TVx�/ y���x��/x�Fw�>�u��Ju�!Uu��Wv�Y_x�E{�$�~����!����Ѓ�j���a���9��%f������I[��/g���؈�U���g��'��Y���Eɐ������呼����o������$�����8ϗ��6��Ȝ�wV��e�������N��LX��o়����ᦼ���B��������0��?;���é�%���#ȭ�Jӯ�l������t과s����������t1���7��/����q��:s��U}��p`��=����  �  �L=ҩK=stK=�TK=�&K=~�J=E+J=[BI=�H=ھF=XSE=��C=2�B=f�A=��@=7�@=#^@=Sn@=-�@=1�@=��@==�@=�l@=�?=��>=�==ƽ<=��;=V;=��:==\:=�N:=�Q:=TF:=::=�9=�8=/�7=��6=Ͷ5=��4=	4= �3=�d3=�\3=7_3=�H3=~�2=�i2=$�1=x0=&;/=,�-=�,=��+=��*=�\*=�!*=�#*=NM*=H�*=�*=��*=Z*=��)=��(=�s'=7�%=Mg$=��"=�!=r= =�=��=��=�=�C=P=_z=��=(�=��=�	={=A==�A=�o =�E�<�l�<��<=�<���<���<O��<a�<U<�<�k�<��<�]�<97�<鎺<�>�<*�<C�<g��<���<�d�<Ŧ�<d��<�m�<Zk�<�ǌ<���<��<O�<�m|<W�u<�n<A{e<��[<��P<OE<@�9<��.<?N$<�(<^1<�)<��<���;���;���;<4�;Ub�;�Ϝ; M�;?iW;�';Z�:��:�::T�t9��I�D_���}�;㲺�&�?f���:�[�b�|l��3����ٯ�/X»K�һ�H�li�u�������
����H��($�S-��6�r�=�;D��-I�e�L��O��Q���R��tU���X�O]���a��bg���l���q��v��.y��{�"�{�aM{��&z�I�x��Fw��mv�t�v���w�z��P}�����A^���烼z���񆅼7��������_��\o��v����@��������Ȍ�2ގ�-��������ɒ�$(��!F���k���ݓ��̔��P���b��O㚼n���U\��u碼������ʲ��x"��@���̧�Pg���"���6���̧����������¬�j ��y��vղ����ô�����7���c��[ص�ɶ��I���J��q�������1��uü�  �  ��K=�6K=K=��J=w�J=��J=��I=I=��G=$F=nE=Z�C=FB=�7A=�y@=�@=��?=B@=�Q@=�@=��@=`�@=�/@=4|?=�>=k==�M<=�U;=x�:=6:=>:=>":=(C:=�P:=�':=��9=��8=��7=�6=z5=�o4=b�3='3=3�2=u�2=� 3=��2=��2=�12=8Z1=�>0=@�.=@�-=�[,=�B+=m*=��)=��)=��)=l�)=�?*=ss*=_s*=:%*=�y)=aq(=�'=g�%=��#=fv"=�!=j�=�=?�=R�=(3=�g=�.=R�=W�=�=N�=ի=?=��=��=� =���<���<���<��<�b�<�h�<��<��<�m�<q��<�)�<�o�<�W�<ɹ</��<?��<;s�<��<4�<�Ԥ<��<Ϛ<᎕<���<��<9Ӈ<�D�<��<)|<̷u<�n<Af<\<��P<�E<39<s-<��"<�~<�v<:�
<z<8�;��;���;+��;���;��;�ā;PQ;~� ;���:�p�:�m:)�9�畹�.��q��������󺀜���?�@�h���K@�������Ż��ջ
�㻘�ﻨp�����d
�s�:��!7$�C�-��6��(?���E���J�l�N�g�P��R��6T��~V���Y�[�]��b�\uh��n��Ss�F�w�{���|�Vx}���|��z{��y�/x�iBw�E^w�>�x��E{���~�E[��B���̄��̅� 9��(��I̅�_j���M��M���qʆ������������Bj��Ra��:Ӓ�����	�������Wr��aH��8���Θ�g[��30����T���������X���7���zڨ�l���駼/������ @��g��:P������,ۯ���������״��f�������h��i]������
���C��%?���ļ�ob�������ü�  �  `~F=�+F=�BF=ƛF= G=W5G=G=H{F=JxE=nD=�B=0�@=Δ?=Bt>=�==�R==O==ǎ==��==�;>=P>=b>=�L==i'<=�:=29=Õ7=1c6=��5=SZ5=W�5=�6=P�6=�7=�47=2�6=��5=�w4=s�2=�91=g�/=��.=�^.=)X.=�.=�>/=J�/=b	0=��/=5_/=pi.=r'-=V�+=�f*=�>)=g(=��'=��'=1(=Dv(=��(=5)=�.)=x�(=�'=�J&=��$=ߎ"=@� =�=U�=W�=E�=8[=3�=�|=d�=�w=x=�=bl=�=ڏ=��=���<[<�<�X�<���<6�<���<��<v��<��<�7�<,��<���<��<O�<>�<�"�<驴<�<���<sp�<p��<~G�<��<vH�<g%�<�<Ɗ�<>ā<��{<۸u<d�p<��l<��g<|�a<��Y<�SO<��B<S�4<��&<*�<?�<�<��;���;�;[��;V��;:U�;eu�;6Н;��;�cX;Jx#;�3�:�#�:a�9�U_�g2�1���+5���k�ټ�o�1��>X�;c������ƍ���Mͻѱ�3�������������H��-���P$��-�9���D���O��mY�K�`��f���h��i�1[i���h�`�h��4j��m�coq���v�l�|�#��A[��d���\ׅ��酼P��E��$���0���ׁ� O��E����م������r��v���Z؏�ː��̐�B������4d��ʁ��G��9����ď��������Q.������Fy���>���#��{h���r��߸����P]��� ���i��vT���j��"Q��к��At���j������1G��|���0䬼P����䬼����(��Q����4���h��Z$��F����$"���w���o��Ⴜ�},��Vͼ�����PH��b�ļV1ȼrh˼�ͼ�  �  9�F=
kF=�~F=]�F=P-G=�YG=O-G=�F=z�E=9D=��B=%A=ӿ?=+�>=��==a�==2y==�==Z>=OV>=h>=�>=�k==�M<=�:=UM9=��7=��6=��5=ғ5=?�5=D)6=F�6=�$7=�97=g�6=�5=7�4=��2=�e1=�0=�/=�.=��.='�.=xq/={�/=:+0=�0=Mw/=L�.=�D-=��+=��*=�j)=J�(=�(=Y(=d4(=+�(=M)=�M)=F)=z�(=�'=�r&=��$=z�"=n� =�D=��=��=�'=Ty=a�=T�=e�=Hw=��=�"=�==��=��=�P�</��<ƽ�<{�<BT�<���<���<y��<���<`q�<%��<:3�<L�<�u�<`��<Z~�<���<��<�<���<`�<ω�<�g�<���<8��<���<��<9H�<,�|<`�v<�q<"m<�>h<yb<?�Y<�`O<��B<i[5<Lx'<�M<U�<o�<ބ�;
��;�'�;��;���;i&�;�'�;;�׆;pkZ;��%;��:�%�:̵�9g.���&��O�������e�l���/���U�����Y��Z����=˻���\������!�c�Wu�!S��j��<$�=�-��8��%D�O���X�D`�e���g���h� �h��h�Oh�{�i�ͷl��
q�wVv�	|�廀�}������Rz��j�������q���6������ާ��Q��+j��R����0�� �����iY���P���^�������u��w:���n��hx��Ə��`���b���;����Θ�}O��i��������������a��Cj���_��i)���Н�R5��_���!������Y`��"������M��t����Q�������^��ճ���ܭ��᯼꠲�q˵��<���&���񚾼˹��|$��X5��Ga�����dǼ�����)���pļ��Ǽ-˼:wͼ�  �  �nG=�G=�&G=fG=ĨG=]�G=�yG=`�F=!�E=8�D=�
C= �A=C9@=^%?=�f>=>=��==�>=�a>=��>=̦>=�a>=+�==Ҵ<=K`;=��9=.~8=�U7=��6=�46=p>6="�6=-�6=�C7=�B7=��6=��5=b�4=-M3=
�1=7�0=�/=#Q/=�F/=��/=�/=�_0=؄0=O0=ص/=��.=��-=�C,=d�*=��)=�)=��(=>(=#�(=!�(=�T)=��)=Q�)=�)=00(=��&=X6%=�a#=��!=~�=��=�}=��=��=\�=ߍ=�=�r=P�=�R=��=�x=7T=��=vO =9��<X��<��<��<���<�@�<^(�<�[�<@�<+��<;�<4	�<c��<3��<�< �<ȩ�<p��<'<�<���<o1�<�7�<���<�ʓ<�<�<ϵ�<�g<.�x<bs<iRn</�h<�0b<�Y<0uO<�pC<�X6<�)<�Y<<x�<F��;x��;U��;Y��;dc�;Db�;��;2q�;�;�`;��,;��:|j�:	:�G	�"O���s��O���޺��q�*�4#P���z�T���X����Żt�ۻ���c���h���U�|\�<���6�M$��z-�7�7�-�B��!M�\.V��S]�QIb��e��;f�Tf��Hf��f��h�R�k� p��u�!�z�
�����	���5o������5���;���@��gx���*����������(�����X����#���򍼹����+������C��Ќ�SB��$n��ဍ�u���������@Ǘ�q��!����X���O������%
����������(����S��M����o���W��$���^��������X��� ��6���?��ޫ��4��LG��$�����J���S����B���1���L�����)A���������.��ο��f��L�����üǼ��ɼ�,̼�  �  }qH=8!H=�H=�7H=QH=>:H=��G=P!G=F=��D=C�C=�'B=�@=��?=K/?=��>=��>=�>=m�>==�>=��>=�>=� >=y<==)<=��:=�u9=-[8=��7=�7=:�6=�7=&H7=�b7=�A7=��6=�6=��4=A�3=�2=�{1=$�0=QV0={F0=w0=8�0=��0=V�0=e�0=0=�/=��-=��,=S�+=\�*=��)=0h)=]9)= H)=8~)=Ȼ)=��)=%�)=�b)=��(=�m'=��%=i>$= �"=r� =i�=?L=�:=v0=�=�=/�=�\='�=��=�M=	=*$=ف=C=߿�<�z�<�`�<E�<�A�<���<��<��<���<*��<�m�<?��<+�<^C�<8��<�.�<M��<yd�<t��<�5�<}�<!F�<3
�<�z�<��<���<Ʌ<\��<�|<,�u<��o<!}i<`0b<��Y<2WO<��C<�7<!+<t;<J�<�W<Z�<���;9��; ��;��;y �;IT�;�Ң;��;c�g;ݡ6;bw;�G�:�?:L.9pA��t�J�|~���?Ѻ����$���H��>q��Ꮋ�>��i��) ӻy�滝M��F��7	����j-�3#�_&$��1-���6��@��xJ���R�1jY�_'^�ca���b�)8c�g�c�>e�Cg���j��n�\}s�sxx�v-}�$�����a߂�}���т��-��Nm���Ѐ����值�݁��}������B����'���狼����u��9S��z׌�T��{��5z������o@���~��l����V���K��/����M���[��b��7���^~��-뙼���W���U���_���<�������਼�z��"}���o꫼ҡ��HT���?��F��������.��i�����'ǵ�_=��$*���i������/���ջ�C�����#м��]�������%üN�ż5VȼSPʼ�  �  T�I=iBI=�!I=nI=��H=ȪH=_ H=,WG=pXF=�3E=��C=R�B= �A=2�@=@=��?=�_?=�F?=�D?=�B?=~*?=,�>=Ap>= �==��<=�;=�:=�~9=��8=�8=��7=g�7=m�7=�h7=i#7=w�6=Z�5=Z5=""4=�03=?c2=�1='z1=b1=�r1=��1=�1=oX1=��0=�50=V/=IW.=N-=�P,=�t+=��*=Q*=�*=��)=A*=�*=$*=��)=��)=��(=X�'=~�&=�*%=��#=�"=^� =�(=2�=ފ={=3p='u=$=�=c�=d�=��	=�=K�=�P=N^ =-�<��<��<���</$�<K�<#|�<���<���<���<oI�<U �<e�<ꪼ<>��<SӴ<�1�<���<(��<��<Z;�<�e�<
B�<��<m�<i�<L��< �<�6x<�q<пi<ϳa<��X<�N<��C<��8<�-<�@"<�R<�<��<{K<S)�;Yk�;pK�;c)�;�߸;��;���;��o;ynA;��;��:[�~:d�9A� ����S����ĺ� ����]CB�k&h������j���`���ɻ�3ݻ2ﻉ��k�����O������$��Q-��X6�<R?�O�G�qO�U���Y�D�\��^���_��}a�I�c��:f�F�i�n�m�7�q�JUv��`z�H�}�A4��8
���j��d��>��Ԧ���I���)��(j���$��c������l������ ۊ�e����?��������0��g�'ȍ�?�����$���ZՔ��[��n��q���4���*���+���{���C��Ɏ��tO��$j����������A���%���������*R��C���¥��h���[Ǫ��1��2��=X���)��/_�����*����巼�T���F��XӺ�c(�����m�����4����h����¼��ļ?�Ƽ�Cȼ�  �  ��J=�EJ=�J=��I=�gI=%�H=�+H=�QG=]F=RZE=�UD=k[C=�uB=5�A=~A=�|@=s@=��?=Ӑ?=�_?=�*?=��>=��>=��==�C==�f<=�s;=�:=>�9=��8=�i8=��7=M�7=u@7=��6=eT6=��5=�5=_4=��3=�+3=��2=
�2=Q^2=^H2=�(2=��1=�|1=D�0=\00=gc/=��.=�-=��,=�?,=i�+=�5+=�*=��*=v*=�S*=,*=J�)=��)=�)=W?(=�4'=W�%=�~$=��"=�o!=1�=&U=��==�=�=7�=�9=И=j�=�F
=��=j=�>=�8=��<Ő�<�[�<g��< �<���<��<g-�<p��<�I�<Y��<*��<0��<�J�<T�<���<ī�<���<eک<��<K��<�X�<���<ٓ<���<�4�<T��<�=�<f
z<ɹq<VFi<�s`<D#W<�SM<� C<��8<��.<7�$<�<Q<��<l�<�.�;��;���;^F�;3��;���;�
�;��u;�K;޲ ;x��:��:�"%:�m�8�t�mVz��6������J�,w?���b�M���Zח�
Z������ޭԻ����s��L2��]�s����t�%�R+.��c6�^H>�v�E���K�$Q��QU�َX�y%[�Z~]��_���b�d%f�ϴi��jm�kq���t��w���z�\�|�sy~������=2���/��='���1��'i��L值����4ꂼ�f�����ʎ��R舼�����Њ��q��� �����%j���h�����:򐼔R��s���Ѧ��+p������]P����������뗼���Ҕ���R��8��,�����ࣼx���Ӧ��`ʨ�2n��@驼�O������==��%���,���-V���������{����ص��x��!и��幼 Ϻ�0�������rɽ�C��ڡ��}>¼F�üHCż�pƼ�  �  2SK=l�J=P�J==J=�zI=��H=��G=��F=�F=:E=}qD=Q�C=C=�fB=��A=�0A=�@=�@=R�?=14?=2�>=M�>=F8>=e�==�e==3�<=�<=�=;=Hf:=�9=��8=(8=Vu7=��6=�M6=��5=�D5=��4=L^4=L�3=��3=Es3=�>3=�	3=~�2=�h2=�1=fC1=׎0=�/=�#/=�~.=�-=oa-=_�,=kk,=��+= �+=)+=�*=�H*=��)=3�)=�3)=��(=�+(=�a'=�Y&=!%=o�#=�"=�Z =Z�=��=b�=�=�\=�=��=�J=��=��
=J<=i=��=�=]1�<k��<W�<�$�<�(�<#$�<7#�<|+�<�<�<~Q�<�c�<�r�<��<��<�Ǻ<�<8��<�W�<H�<"^�<�<���<Lk�<��<yp�<ĺ�<j��<�1�<
�z<�_q<?�g<G^<}�T<�K<boA<,8<��.<�)&<��<)�<�8<đ<ha�;c��;K�; ��;���;�^�;�$�;K�w;h�Q;�+;6;;�s�:��X:��u9���7o��ľ�oq��="��_B���b��-�����r覻4���gλ7J�����<��������)����'�g�/��\7�W2>��SD�r�I��NN��GR�W�U�Y��j\���_�ȷc��yg��k�]_n��Mq�0�s�Xv��x�'�y��k{�n�|�0L~�^��=��[���7‼��� a��\ˁ��x���t������2�������戼�2��(c���|��?���\���}��
m��Q��u#���ܒ�z�����?������}˕��˖�Y�������L������Ꙟ���冡�ע�H���I��nt��ݔ��l���?�������G����������PW���>���m��z簼v���`��(��^ݷ�v��~�S��=���"龼�#��R���o¼�uü�]ļ�'ż�  �  �K=�IK=ȽJ=�J=� I=w#H=�$G=�9F=�oE=��D=�ED=��C=+fC=m�B=�XB=حA=��@=Q%@=�b?=��>=�.>=��==��==T==|==�<=w@<=��;=
�:=��9=��8=~�7=�7=w?6=S�5='5=��4=kJ4=i4=0�3=�3=��3=B�3=5N3= �2=n;2=�v1=��0=��/=�/=��.=�#.=��-=ȓ-=�M-=_�,=K�,=[�+=N+=��*=#�)=�Y)=��(=q(=d(=p�'=!'=�X&=�G%=6�#=�R"=�} =z=pS=G=��=}=.3=��=̾=̗=sz
=>a=�D=�=p�=x�<��<���<���<w��<���<	�<Ε�<6>�<u��<�[�<��<��<�u�<�.�<��<|�<�A�<���</�<	r�<��<�I�<�^�<_�<���<ᝇ<��<I�z<M�o<�e<=[<�SQ<S�G<��><bL6<y-.<�\&<{�<`<5(<��<w0�;u�;N�;��;g��;�N�;3ɋ; �u;�
T;2�1;��;I�:�m~:9��9"����_v��rʺ�-
�k3,��K�ץi��̓�U��������M��&˻�߻�������"H�
,��m"���*�ˊ2��G9��'?�1FD���H���L���P�:�T�r�X�)]��a��/f�LYj�_�m���p�4�r�'!t��=u��Rv� �w�g5y�*{�7a}�����‼����BI��/�������j���a₼�Z��w2��a���Ԇ��u��0+��R܋�s��8܎�A������Q���[-��c���������eL���ӓ�����\͕��S�����S���jƜ�]V��r�������h}���F��"$���+��@g��Ӧ�^���ꩼ1U�����Bi��|������� ���������+���������������������m��V��"t��ѕ���w¼S"ü�ü<ļ�ļ�  �  `�K==K=k�J=�I=#mH=<G=z F=T5E=l�D=�D=#�C=�C=��C=4C=��B=��A=nA=��?=��>=��==�>==��<=�<=~v<=Gt<=�\<=�<=&�;=��:=��9=��8=,�7=v6=`y5=�4=�4=S�3=5�3={�3=��3=�3=��3=��3=�53=��2=�1=��0=[�/=��.=�!.=��-=-=Ђ-=��-=�}-=�E-=��,=G',=�I+=cQ*=�[)=`�(=��'=�b'=�'=��&=��&=B�%=�%=�#=�C"=BV =O&=��=T=��=#|=/4=�=Q=�=5,
=�:=�0= ={�=9�<ӟ�<��<;��<�d�<���<Ok�<��<���<b��<���<1U�<wN�<���<��<�N�<ν�<���<i�<w'�<���<T��<�j�<8��<
	�<z��<���<�D�<�Fy<��m<�{b<��W<TyM<�D<��;<��3<��,<�z%<�V<Z�<ǭ<��<y�;���;]��;�P�;za�;��;�b�;�wo;!�R;̒4;�l;���:���:�]�9֪��톺G�޺�i���:�QZ�Qv��R���2��ٙ�����pʻE�߻����wN����R"�]�%��k.���5���;���@�1;E�lI���L�P�P�%�T���Y��#_�۰d�*�i��kn���q���s��u��au�'_u�?�u��Qv�q�w�Qz��g}��g������[���>�����������P�����_����l���_��F͆���������Ì��Ď�����ّ��Œ��E���h��FN��@!�����A��fۓ�H�'���3����Κ������՞��>��D*��%����.��}�������#Τ���������6��������G��nn������_���u�������#�� ��#���z����ʷ�}6��<���;޾�����E¼tQü��ü�:ļOPļ_ļ�ļ�  �  K=��J=(J=��H=��G=\1F=��D=HD=X�C=�GC=�JC=�hC=(wC=fNC=��B=%B=��@=1�?=�G>=M==Y2<=��;=�h;=t;=w�;=L�;=�;=sH;=��:=�9= _8=�7=��5=Y�4=6�3=K.3=�2=U�2=�3=O3=l�3=ה3=b3=��2=Y2=[�0=��/=)�.=t�-=�-=��,=I�,=	-=vS-=�~-=Ef-=�,=w,,=*+=r�)=��(=��'=&�&=�8&=F�%=�%=r�%=�d%=��$=K�#=�!=��=E�=�%=��=��=/{=�4="=�==x=Y�	=#�=��=̪=�(=���<���<u��<�6�<��<Iz�<D��<`(�<���<9��<��<��<͘�<���<��<uX�<TD�<���<���<���<&��<�ߙ<��<�<�y�<�-�<64�<�<�qw<{Dk<�I_<��S<��I<Z@<�68<�1<Ng*<4�#<%-<J�<J<_�<y�;y>�;�;�;�R�; �;��;�f;��N;�y4;V;���:���:���9g�˹���Z���&�Z�K���j��u��_��V����h��T���b�˻�%�mV���-����E��X)�1 2��9�g�>�.C�V�F��J��~M�rsQ��0V��[�pb�bh�M:n�g�r�D+v�S�w�.x�Bw�.1v�q�u�9�u��Vw�H4z�� ~�:J��7s���;��l��q솼Yˆ�:��J������6!��]؅��7��%��aq���፼+6���2������q����씼�Ȕ��X���ړ�
���c���G]�����������-���ʜ�,3������^��\󢼅���.����p��L���R5������������������>���F��٪���^���|��2@��> ��2��������������f��V���۽�h����¼�ļ�ż}�ż�~żR>żPż%ż�  �  �1K=:�J=�I=8<H=ɹF=�=E=m�C=)C=B=@�B=�B=�C=�PC=�KC=��B=E�A=C�@=�4?=�==�J<=k?;=��:=�f:=��:=g�:=7;={2;=b�:=�F:=�C9=��7=Y�6=�-5=x�3=� 3=�e2=�%2=k62=��2= �2=�/3=XI3=�3=4v2=�|1=�<0=�.=�-=��,=�
,=O�+=�,=̉,=	-=f-=Oi-=�,=R,=��*=�b)=��'=}�&=޿%=�.%=�$=��$=��$=x�$=�=$=�4#=R�!=��=�4=��=��=�#=I�=�\=+X=�=��
=�A	=I�=�=D=�� =Ht�<�<�<t �<s!�<]��<��<��<��<$�<H�<��<3��<h��<��<��<�U�<�ج<� �<#
�<��<�ښ<@�<�Ε<��<式<��<�<���<u<�h<+x\<��P<cQF<�#=<D5<Zy.<�U(<�H"<L�<�S<_�<Ԗ<���;�j�;VH�;��;Y;�;���;��s;^;��I;��2;l�;r��:%��:1L�9�F��� ���w��4�g�Z���y�k���K��:���֫��:����ͻ7f�2��+
��l��"�'[,��5��<��UA��LE�\pH�AZK�ߚN�/�R���W�}�]� �d���k��r� w�Qz�J{���z��9y��Iw�x�u���u��?w���z��#��:��l҄�����Xa������%ň�p ������8������~��g·�Ή�PG�������p���R>��)#���\��f��M\��!���T0��_B��o������a�����A��� 4���&��SJ��뛤��B������ܢ��G&��c���%ܦ������׬�v������(����h��i��=�G_�� ��9�������ؓ��#��+��u�������ļ��ż͝Ƽu�Ƽ�Ƽ�-Ƽ��ż�ż�  �   �J=�EJ=;.I=B�G=�#F=ŔD=�GC=bB=��A=�A=	MB=x�B=�,C=�?C=�B=>�A=��@=�>=Q6==S�;=d�:=A�9=\�9=$�9=�D:=B�:=��:=��:=q:=9=L�7=76=��4=�w3=�|2=?�1=��1=K�1=�2=��2=��2=�
3=��2=n"2=�1=��/=�B.=��,=!�+=}\+=�B+=A�+=�),=��,=K-=b-=I�,=��+=��*=)=�p'=�&=�%=zx$=?A$=�L$=�g$=�U$=��#=��"= `!=�Q=��=�!=T=)�=Z=��=��=J=�{
=��=8=�B=K�=�B =/}�<�<���<��<�z�<�$�<H��</��<�t�<���<���<���<?��<�p�<���<��<Oӫ<ɥ<W��<C��<S��<��<֔<�O�<�!�<��<��<t`�<4t<6<g<�Z<��N<A"D<Y�:<�D3<��,<��&<
!<Ĭ<<7<�R
<W��;���;A��;��;�G�;:��;1��;1.k;Z�W;VlE;��0;�o;�_�:g�:m	�9������(����>�1\e��$���R��Ӕ���������;_��,�ϻmK� q��r�,���#�~a.�s7���=��C���F���I�>`L�a�O�~�S��Y���_�E�f��Bn�B�t���y�=�|���}���|���z�J3x�QHv���u�Uw���z����-�Oυ�+������C^��7"���>��������������:K���T���茼���g��ѩ��>I���,��~V���於���`?��)�����������X��Uٙ��֜�"柼h�������ʝ���ƥ�=1��A2��#;���Ģ��.��������C������:Ѱ��\����� ϵ�w���?!��_��d볼% ��,������������ѿ�[�¼żo�Ƽ{�Ǽ��ǼW~Ǽ�ƼWMƼ�!Ƽ�  �  �J=!(J=C	I=��G=��E=�XD=]C=P#B=�A=}�A=T%B=b�B=�C=:C=
�B=�A=*y@='�>===��;=�[:=�9=jv9=�9=i:=�|:=ϱ:=V�:=�9=��8=��7=h6=l�4=FL3={N2=��1=�x1=��1=j�1=�o2=��2=��2=��2=�2=��0=g�/=�
.= �,=��+=�+=�
+=d+=,=�,=�?-=�]-=z�,=��+=͈*=m�(=B'=��%=��$=	8$=$=*$=�4$=c+$=�#=��"=[E!=r5=��=-�=(=Cj=��=\�=��=��=�V
=.�=H=�(=�= =�%�<���<�6�<�6�<���<���<B�<p��<�6�<���<E��<���<X��<'X�<�j�<�G�<�r�<6W�<�9�<F-�<%�<婖<<x�<��<<�<�ߊ<)�<�'�<�s<P�f<�Y<v�M<�_C<?:<Α2<`,<-N&<�� <�G<��<�	<���;�j�;���;��;V�;�Ɏ;��;�$h;�GU;��C;y0;C;uc�:�t�:�9iL���w��B�p-i����� ��S/��}������@���lл*��U����β�&�$��/���7��>�D�C�=`G��&J�o�L���O��T�H�Y��3`��g��!o���u�A�z���}���~���}�+D{�3�x�tv�L�u�
cw�{�o*��w6��1+������K5��9݊�@���Ұ���v��1f��a膼)>��5{�������$��<�������_��/�����������5��U]���y���䔼z��ӕ�0����.���=���Z�����K������1��T��� q���`���Ԣ��4��H����8���v��H���04���г������M��	8��ˎ��E���07���\���^���A���߹�}�	��üNkż�Ǽ�Ǽz,ȼi�Ǽ Ǽ�Ƽ�QƼ�  �   �J=�EJ=;.I=B�G=�#F=ŔD=�GC=bB=��A=�A=	MB=x�B=�,C=�?C=�B=>�A=��@=�>=Q6==S�;=d�:=A�9=\�9=$�9=�D:=B�:=��:=��:=q:=9=L�7=76=��4=�w3=�|2=?�1=��1=K�1=�2=��2=��2=�
3=��2=n"2=�1=��/=�B.=��,= �+=|\+=�B+=@�+=�),=��,=K-=b-=E�,=��+=��*=)=�p'=�&=�%=px$=6A$=}L$=�g$=�U$=��#=��"='`!=R=)�=�"=�T=K�=�=��=��=�=�~
=�=�;=G=��=G =3��<!�<յ�<���<ق�<�+�<���<���<y�<���<���<T��<C��<5n�<��<:��<nͫ<G¥<���<��<���<��<9͔<�F�<>�<��<��<AZ�<�)t<4g<L�Z<��N<
"D<� ;<J3<��,<�&<Y!<ۺ<�F<�c
<Z <��;���;0�;�i�;�Ӑ;֮�;�_k;Q�W;��E;z�0;�y;�]�:Nڏ:�Q�9�$�uv��s���>���e��H��,x��[����⢻ ���N���|�ϻl廐�����\"�<�#�wj.��#7��>�� C���F���I�}bL��O�έS��Y�W�_���f�Cn���t��y�o�|�ڻ}���|���z�[3x�^Hv���u�Uw���z����/�Qυ�+������C^��7"���>��������������;K���T���茼���g��ѩ��>I���,��~V���於���`?��)�����������X��Uٙ��֜�"柼h�������ʝ���ƥ�=1��A2��#;���Ģ��.��������C������:Ѱ��\����� ϵ�w���?!��_��d볼% ��,������������ѿ�[�¼żo�Ƽ{�Ǽ��ǼW~Ǽ�ƼWMƼ�!Ƽ�  �  �1K=:�J=�I=8<H=ɹF=�=E=m�C=)C=B=@�B=�B=�C=�PC=�KC=��B=E�A=C�@=�4?=�==�J<=k?;=��:=�f:=��:=g�:=7;={2;=b�:=�F:=�C9=��7=Y�6=�-5=x�3=� 3=�e2=�%2=k62=��2= �2=�/3=XI3=�3=4v2=�|1=�<0=�.=�-=��,=�
,=M�+=,=ɉ,=-=�e-=Ji-=x�,=J,=��*=�b)=��'=m�&=Ϳ%=�.%=
�$=��$=��$=w�$=�=$=�4#=��!=A�=k5=َ=)�=�%=&�=�`=�\=@�=|�
=�H	=��=�=KL=J� =���<aN�<��<�1�<���<��<^��<h��<G&�<�M�<N��<���<���<n��<��<�L�<dͬ<��<p��<���<7ʚ<�.�<���<��<Ȭ�<��<I��<��<��u<m�h<Wm\<!�P<�PF<�(=<%N5<`�.<?i(<�`"<��<+r<��< �<�'�;9��;&��;h'�;�x�;�ކ;n$t;k^;��I;��2;ž;���:�|�:��9�K���ǩ�����(5��W[��Qz��������焟�� ��e���;λ���l���(
�D���"�wl,��5�|<��^A��SE�vH��^K�8�N���R���W���]��d�^�k�Wr�~w��z�UJ{���z��9y� Jw���u��u��?w���z��#��:��n҄�����Ya������%ň�p ������8������~��g·�Ή�PG�������p���R>��)#���\��f��M\��!���T0��_B��o������a�����A��� 4���&��SJ��뛤��B������ܢ��G&��c���%ܦ������׬�v������(����h��i��=�G_�� ��9�������ؓ��#��+��u�������ļ��ż͝Ƽu�Ƽ�Ƽ�-Ƽ��ż�ż�  �  K=��J=(J=��H=��G=\1F=��D=HD=X�C=�GC=�JC=�hC=(wC=fNC=��B=%B=��@=1�?=�G>=M==Y2<=��;=�h;=t;=w�;=L�;=�;=sH;=��:=�9= _8=�7=��5=Y�4=6�3=K.3=�2=U�2=�3=O3=l�3=ה3=b3=��2=Y2=Z�0=��/='�.=s�-=�-=��,=E�,=	-=qS-=�~-==f-=�,=k,,=+=a�)=��(=v�'=�&=w8&=-�%=�%=c�%=�d%=Ĵ$=��#=��!=�  =d�=k'=�=��=<=�9=9(=E=h�=��	=c�=��=t�=�4=I��<k��<��<�M�<�<��<���<�6�<��<Z��<x�<���<��<h��<O��<oK�<W4�<��<��<O�<���<�Ǚ<��<2��<&c�<��<� �<��<bUw<o.k<�:_<��S<�I< a@<�D8<�1<�*<�$<�S<�<x<��<%��;ɡ�;Ol�;�z�;m��;P�;�7�;�Mg;��N;f�4;�-;$��:
x�:\��9	�ι®��Pw��O'��^L��nk�f܂�NȎ�A���LѨ�����̻��w����R��1��b�q)��2�/9���>�z8C�s�F�J���M�wQ�|3V�*�[�b�Lch�8;n��r��+v���w�}x�@Bw�\1v���u�S�u��Vw�W4z�� ~�?J��;s���;��l��s솼Zˆ�:��J������6!��]؅��7��%��aq���፼+6���2������q����씼�Ȕ��X���ړ�
���c���G]�����������-���ʜ�,3������^��\󢼅���.����p��L���R5������������������>���F��٪���^���|��2@��> ��2��������������f��V���۽�h����¼�ļ�ż}�ż�~żR>żPż%ż�  �  `�K==K=k�J=�I=#mH=<G=z F=T5E=l�D=�D=#�C=�C=��C=4C=��B=��A=nA=��?=��>=��==�>==��<=�<=~v<=Gt<=�\<=�<=&�;=��:=��9=��8=,�7=v6=`y5=�4=�4=S�3=5�3=z�3=��3=�3=��3=��3=�53=��2=�1=��0=Z�/=��.=�!.=��-=��-=ʂ-=��-=�}-=�E-=��,=9',=�I+=OQ*=�[)=E�(=e�'=db'=�'=��&=��&=A�%=�%=_�#=D"=*W =�'=��=�V=��=�=e:=e=0=�=�7
=�G=P>=d=L�=e6�<���<s#�<���<G�<���<���<��<��<T�<���<_V�<*K�<���<��<?�<G��<ֈ�<��<�<Л�<�u�<�L�<ٔ<�<bz�<��<0�<$y<��m<Mib<��W<�xM<'D<�;<��3<~�,<k�%<ƅ<�<2�<��<ܕ�;��;O�;5º;˧;�y�;W��; p;>S;t�4;s�;��:�O�:���9dR������ຈ1�5�;�
[� w�oӈ�d���������T�ʻ��߻�A��I|���|E�@�%���.�>�5���;��A�>EE�,I�q�L�ԣP���T�`�Y��%_�Z�d�M�i��ln�g�q�=�s�0u�<bu�__u�j�u��Qv���w� Qz��g}��g������[���>�����������P�����_����l���_��G͆���������Ì��Ď�����ّ��Œ��E���h��FN��@!�����A��fۓ�H�'���3����Κ������՞��>��D*��%����.��}�������#Τ���������6��������G��nn������_���u�������#�� ��#���z����ʷ�}6��<���;޾�����E¼tQü��ü�:ļOPļ_ļ�ļ�  �  �K=�IK=ȽJ=�J=� I=w#H=�$G=�9F=�oE=��D=�ED=��C=+fC=m�B=�XB=حA=��@=Q%@=�b?=��>=�.>=��==��==T==|==�<=v@<=��;=
�:=��9=��8=~�7=�7=v?6=S�5='5=��4=kJ4=i4=0�3=�3=��3=B�3=4N3=��2=m;2=�v1=��0=��/=�/=��.=�#.=��-=��-=�M-=T�,=>�,=K�+=�M+=x�*=�)=oY)=��(=�p(=B(=S�'=� '=�X&=�G%=��#=!S"=�~ =�{=�U=~=*�=��=:=�=��=%�=0�
=>o=�S=�+=��=#�<h'�<���<|��<���<���<� �<���<�M�<���<b�<Z��<4��<�l�<Y!�<�<�ٰ<�(�<_ݧ<��<�Q�<�˜<�(�<q>�<0��<ec�<y��<�l�<�hz<U�o<ke<�2[<�RQ<��G<��><)i6<S.<m�&<�<�B<)g<'<Է�;��;ҝ�;o�;��;︝;"%�;�>v;�~T;��1;�;�A�:��}:��9W�����x�f�˺�*-�ܹL�M�j�Y]��-���O��7ط��˻X*��8���%�Hu�2S�َ"��+���2�Z9�%6?��QD���H���L���P��T�b�X�c]���a��0f�EZj��m�C�p���r�z!t�->u��Rv�D�w��5y�%*{�Ga}�����‼����EI��1�������k���b₼�Z��x2��a���Ԇ��u��0+��R܋�s��8܎�A������Q���[-��c���������eL���ӓ�����\͕��S�����S���jƜ�]V��r�������h}���F��"$���+��@g��Ӧ�^���ꩼ1U�����Bi��|������� ���������+���������������������m��V��"t��ѕ���w¼S"ü�ü<ļ�ļ�  �  2SK=l�J=P�J==J=�zI=��H=��G=��F=�F=:E=}qD=Q�C=C=�fB=��A=�0A=�@=�@=R�?=14?=2�>=M�>=F8>=e�==�e==3�<=�<=�=;=Hf:=�9=��8=(8=Vu7=��6=�M6=��5=�D5=��4=K^4=L�3=��3=Es3=�>3=�	3=}�2=�h2=�1=dC1=Վ0=	�/=�#/=�~.=�-=ha-=V�,=`k,=��+=�+=+=�*=�H*=|�)=�)=�3)=l�(=�+(=�a'=�Y&=D%=ǥ#=_"=�[ =�=��=��=x�=�b=�=2�=,U=h�=(�
=�J=	=E�=9�=5T�<3��<`(�<;E�<%G�<�?�<�;�<�?�<)M�<�\�<Tj�<#t�<1~�<��<��<��<���<�=�<�*�<�>�<�_�<�m�<�H�<��<+P�<���<܆<��<(�z<�@q<��g<�;^<��T<oK<T�A<�$8<�/<�X&<z<�%<�y</�<���;�A�;]��;��;I�;̢;��;0�x;~ R;�Q+;b;-l�:��W:0qp9���A�q��T��cW��<#��rC���c�R�����~|�����7�λ��JZ����y�x�����(��0��o7�oA>�{_D���I��UN�)MR�h�U�&Y�9m\���_��c��zg�Gk��_n�%Nq���s��v��x�L�y��k{���|�@L~�j��=��^���:‼���"a��]ˁ��x���t�� ���2�������戼�2��(c���|��?���\���}��
m��Q��u#���ܒ�z�����?������}˕��˖�Y�������L������Ꙟ���冡�ע�H���I��nt��ݔ��l���?�������G����������PW���>���m��z簼v���`��(��^ݷ�v��~�S��=���"龼�#��R���o¼�uü�]ļ�'ż�  �  ��J=�EJ=�J=��I=�gI=%�H=�+H=�QG=]F=RZE=�UD=k[C=�uB=5�A=~A=�|@=s@=��?=Ӑ?=�_?=�*?=��>=��>=��==�C==�f<=�s;=�:=>�9=��8=�i8=��7=M�7=u@7=��6=eT6=��5=�5=_4=��3=�+3=��2=
�2=P^2=]H2=�(2=��1=�|1=B�0=Y00=cc/=��.=�-=��,=�?,=^�+=�5+= �*=��*=v*=jS*=�+*=*�)=x�)=�)=;?(=�4'=Z�%=$=�"=wp!=@�=�V=�=A=#=K=�=�A=��=��=�S
=��=y=�N=5I=���<_��<�|�<���<��<��<���<7A�<��<�T�<��<}��<��<:B�<Թ<ߞ�<��<���<<��<L¥</��<�7�<Ϗ�<븓<�ڎ<��<ބ�<�&�<��y<ӛq<�1i<�h`<{"W<�\M<�3C<F�8<+�.<��$<��<��<��<��<e��;^�;&�;���;��;u#�;�f�;Kv;�wK;� !;��:��:�m$:緓8�W��|�︾��B���@���@�ϙc��!h��)鬻�\��2ջ<�_���\e�����Ź�6�%�B.�4v6�W>���E���K��*Q�1WU�ӒX�|([���]�� `���b�b&f���i�vkm��q��t�S�w�Ěz���|��y~�-�����C2���/��A'���1��)i��N值����5ꂼ�f�����ʎ��R舼�����Њ��q��� �����&j���h�����:򐼔R��s���Ѧ��+p������]P����������뗼���Ҕ���R��8��,�����ࣼx���Ӧ��`ʨ�2n��@驼�O������==��%���,���-V���������{����ص��x��!и��幼 Ϻ�0�������rɽ�C��ڡ��}>¼F�üHCż�pƼ�  �  T�I=iBI=�!I=nI=��H=ȪH=_ H=,WG=pXF=�3E=��C=R�B= �A=2�@=@=��?=�_?=�F?=�D?=�B?=~*?=,�>=Ap>= �==��<=�;=�:=�~9=��8=�8=��7=g�7=m�7=�h7=i#7=w�6=Z�5=Z5=""4=�03=?c2=�1='z1=b1=�r1=��1=�1=nX1=��0=�50=V/=EW.=N-=�P,=�t+=��*=�P*=�*=��)=-*=�*=
*=��)=|�)=��(=?�'=o�&=�*%= �#=0"=� =�)=��=��=d=t=z=P*=��==�=��=1�	=�=ޒ=#_=)m =�K�<)��<��<���<�>�<I�<@��<���<���<���<O�<��<�<,��<E��<kô<%�<�v�<맩<���<��<9H�<F$�<��<`Ȍ<1 �<���<n`<!x<� q<G�i<�a<G�X<p�N<��C<Y�8<�@-<�i"<��<��<30<׆<ˢ�;���;��;���; I�;���;��;�Qp;��A;�";���:�~~:��9���p��s��*�ź�� ��� �N1C�� i�d-���잻ᴻ�ʻE�ݻ4q�`l��@�,�\����}�$�lf-�Ii6�l_?���G��O�EU�J�Y�ޗ\�Б^�� `�ka�y�c��;f���i��m���q��Uv�7az�t�}�Q4��E
���j��#d��D��ئ���I���)��*j���$��c������l������!ۊ�e����?��������0��g�'ȍ�?�����%���ZՔ��[��n��q���4���*���+���{���C��Ɏ��tO��$j����������A���%���������*R��C���¥��h���[Ǫ��1��2��=X���)��/_�����*����巼�T���F��XӺ�c(�����m�����4����h����¼��ļ?�Ƽ�Cȼ�  �  }qH=8!H=�H=�7H=QH=>:H=��G=P!G=F=��D=C�C=�'B=�@=��?=K/?=��>=��>=�>=m�>==�>=��>=�>=� >=y<==)<=��:=�u9=-[8=��7=�7=:�6=�7=&H7=�b7=�A7=��6=�6=��4=A�3=�2=�{1=$�0=PV0=zF0=w0=8�0=��0=U�0=d�0=
0=�/=��-=��,=N�+=U�*=��)=&h)=R9)=H)='~)=��)=o�)=�)=�b)=��(=�m'=��%=l>$=<�"=�� =�=M=<=12=?=/�=>�=�a=G�=Ώ=�U=j&	=z.=�=�N=)��<e��<qy�<Q)�<�X�<h��<���<P�<4��<���<%v�<��<% �<�@�<��<�$�<I��<�T�<��<V!�<3�<�.�<�<�b�<�ʏ<�|�<���<劁<��{<ԯu<��o<�mi<m(b<�Y<^O<��C<�7<�6+<	]<
�<��<��<�3�;s�;F�;Zw�;�|�;��;��;�[�;�Rh;F�6;��;+�:�?:�6,9m:��B8L�j���ZҺ���%��uI�1r� K�����ҽ�!�ӻ���u�������8	� �	J��;��:$�MB-�h7��A��J���R�KoY�F+^�Za���b��9c���c�7e��Cg�6�j���n��}s��xx��-}�6������k߂�����т��-��Qm���Ѐ����值�݁��}������C����'���狼����u��9S��z׌�T��{��5z������o@���~��l����V���K��/����M���[��b��7���^~��-뙼���W���U���_���<�������਼�z��"}���o꫼ҡ��HT���?��F��������.��i�����'ǵ�_=��$*���i������/���ջ�C�����#м��]�������%üN�ż5VȼSPʼ�  �  �nG=�G=�&G=fG=ĨG=]�G=�yG=`�F=!�E=8�D=�
C= �A=C9@=^%?=�f>=>=��==�>=�a>=��>=̦>=�a>=+�==Ҵ<=K`;=��9=.~8=�U7=��6=�46=p>6="�6=-�6=�C7=�B7=��6=��5=b�4=-M3=
�1=6�0=�/=#Q/=�F/=��/=�/=�_0=ׄ0=O0=׵/=��.=��-=�C,=`�*=��)=�)=��(=6(=�(=�(=�T)=��)=A�)=�)= 0(=��&=Q6%=�a#=��!=��=�=�~=��=��=�=�=��=v=��=�W=j�===�[=~�=�W =k��<���<K#�<�%�<ϛ�<�O�<66�<"h�<��<S��<!�<��<��<C��<�z�<ݵ<���<,~�</�<lt�<�!�<�&�<u��<Ź�<!�<�n�<���<L<�x<�Ms<�Bn<z�h<V+b<��Y<zO<�zC<�g6<X)<�q<�(<��<� <#��;���;r��;ӧ�;���;�J�;맠;�N�;�f`;2-;���:���: w	:�3�i�Y�t�\���w�ߺ����s+�w�P�ic{��>��lӭ�q�Ż��ۻ�(�������p��s�y���G��+$���-���7���B��'M�3V�BW]�Lb�� e�A=f�8Uf��If���f���h���k�O p�u�M�z�+��������<o��Ò��9���;���@��ix���*����������)�����Y����#���򍼹����+������C��Ќ�SB��$n��ဍ�u���������@Ǘ�q��!����X���O������%
����������(����S��M����o���W��$���^��������X��� ��6���?��ޫ��4��LG��$�����J���S����B���1���L�����)A���������.��ο��f��L�����üǼ��ɼ�,̼�  �  9�F=
kF=�~F=]�F=P-G=�YG=O-G=�F=z�E=9D=��B=%A=ӿ?=+�>=��==a�==2y==�==Z>=OV>=h>=�>=�k==�M<=�:=UM9=��7=��6=��5=ғ5=?�5=D)6=F�6=�$7=�97=g�6=�5=7�4=��2=�e1=�0=�/=�.=��.='�.=xq/=z�/=9+0=�0=Mw/=K�.=�D-=��+=��*=�j)=G�(=�(=U(=_4(=%�(=F)=�M)=�E)=q�(=�'=�r&=��$=|�"=x� =�D=�=��=�'=�y=A�=|�=��=!y=3�=�%=�=�=��=��=3Y�<��<���<|'�<]�<, �<���<���<���<�v�<`��<?6�<�<Pv�<^��<|�<���<�ޱ<8ݮ<բ�<��<���<]_�<٠�<Q��<���<X�<X@�<ݯ|<܃v<��q<�m<49h<�b<	�Y<(cO<� C<'c5<v�'<Z<��<<�<ئ�;���;L�;74�;Y��;,H�;G�;A��;4��;R�Z;B&;T��:):�:���9@�.��%'�Ԓ��/�h�����'0��<V��'��E���9Ѳ�Md˻���	�����81�%�v���]�ys�0D$�[�-���8��)D�-O�#�X�&`��e���g���h���h�Ch�^Oh���i��l��
q��Vv�&	|���������Uz��m�������r���7������ߧ��R��+j��R����0�� �����iY���P���^�������u��w:���n��hx��Ə��`���b���;����Θ�}O��i��������������a��Cj���_��i)���Н�R5��_���!������Y`��"������M��t����Q�������^��ճ���ܭ��᯼꠲�q˵��<���&���񚾼˹��|$��X5��Ga�����dǼ�����)���pļ��Ǽ-˼:wͼ�  �  ��<=ױ<='G==�Y>=��?=³@=�ZA=	hA=��@=��?=�W>=��<=eZ;=0:=k9=9=�9=�c9=��9=o�9=�9=��8=��7=	�5=03=9�0=��.=M�,=3,=,=��,=��-=�R/=yh0=��0=y�0=�h/=��-=<+=�(=��&=�%=%=�\%=�P&=�'=�)=�D*=��*=��*=�q*=nr)=�-(=P�&=Ӷ%=��$=	y$=Tw$=�$=�G%={�%=��%=1�%=�$=�#=6� =�7=d�=�#=8=�=�N=�-=�@=�&==N�=��==��=�q=d =*"�<��<��<,�<X��<#��<���<��<|:�<�-�<��<x��<c�<�I�<�ؾ<c�<#�<Nد<eG�<�
�<K��<��<9T�<\��<���<�r�<���<�wt<�{g<R:]<�V<%�Q<��O<�{N<ZL<��G<�[@<�5<��&<<�<!H�;ʲ�;�¸;Vܪ;."�;᭟;��;���;U�;���;�$o;þC;��;���:)�:�� �cW��o���#��e���C/�P�J�6rk��ቻ�����t��)5߻�x��������#�%�M�,�4�0�y03��4�_�7�zk<��ID��;O�^�\�v"k�Ly�����4F���ቼw����ĉ�釼�����߃�zꂼB��AT��9m��R�������獼{}���;��~!���W��,0�����Z}��8̌��H��	��Yޔ��P��ٷ��;k���᣼iȤ����	���A��J�������G��r坼��������A��$ꮼ&��P����հ�	Ȯ�V(��Q���Tا��2��^Ч�(���������j��(���
J��l8��N[��X趼�9�����,쵼������  ��@����Ƽ�V˼ϼ|Ѽ�<Ҽ
kѼalϼ6�̼k�ʼnɼR�ɼ!�˼�Lϼt�Ӽ��ؼ{�ݼ����  �  �>==$==��==��>=��?=��@=E�A=�A=��@=��?=�y>=@�<=;=�a:=�9= D9=�G9=׉9=R�9=�9=D�9=�9=�7=��5=�{3=C1=!�.=4d-=��,=t,=�-=�A.=��/=ݏ0=�1=)�0=�/=��-=�z+=�5)=�G'=��%=~%=��%=O�&=��'=�Z)=Qv*={+=�+=��*=�)=oQ(=�'=��%=�%=Z�$=��$=��$=�k%=�%=K&=Y�%=o�$=�6#=�!=؆=��=i�=3�=U=��=.z=�|=�R=t�=�=��=z4=�	=Ϯ=�Q =���<ރ�<r��<	��<"/�<N�<z�<BJ�<�s�<�^�<� �<��<�W�<���<�9�<�s�<�s�<
:�<z��<�X�<��<+4�<��<��<�j�<�	�<�`�<�v<9i<��^<�W<�WS<�Q<_iO<#M< vH<��@<N�5<�B'<(�<��<���;1��;��;��;i�;�?�;���;���;Zy�;q�;�p;�}E;?�;/��:J):|�ظW�I�$���Y�����,��H��9i�������8h���ܻ�k���&����2$�rD+��/�a2�o�3���6�j�;���C�٩N���[��!j�Cx�Q���t�����Ɖ�q���A��1��8{��#����؂����S/��U����O�����z��@֏�&�D��L獼J׌�$E�������� ���^����������$����	�������U��Hh���������>��]����ښ�\���񔡼�+������'���R��7谼����������)���~���寮M���^U���ޫ�Qͮ�I���$��u䵼�Զ�b�����������~���N���6ܶ��1��۵��i&��k�ż4�ʼ^Eμ��м2qѼ��м�μ't̼�Tʼ/-ɼ�~ɼ�y˼��μ
Ӽ�]ؼC�ܼL+��  �  m>=/I>=��>=��?=�@=�yA=5�A=�A=�6A=)@=J�>=^==�<=��:=�,:=j�9=��9=4�9=,:=,D:=�:=�T9=8=Y^6="G4=�2=�0=y�.=I�-=k�-=�.=�/=0=��0=�Q1=k�0=�/=y6.=d(,=�*=�N(=�!'=��&=Q�&=�'={�(=l
*=M�*=�n+=�_+=��*=��)=ح(=�v'=�g&=��%=�8%=�)%=qe%=R�%=�$&=C&=��%=%=�#=6�!=�\=��=�=s�=7r=C�=�P=�#=*�=��=P=��=��=%�	=H[=�,=^��<��<�(�<q�<��<��<�.�<E�<O�<���<
��<��<��<Չ�<qI�<���<���<�E�<戭<q�<��<�Т<�G�<n��<"��<<�J�<(�z<en<��c<tI\<�[W<OT<��Q<>�N<ԲI<?�A<�6<��(<�)<x�<�>�;��;���;���;�e�;�i�;���;���;Rw�;���;�t;P�I;�B;.g�:�J:��8�D#������ݺƍ�F�&��C��c�ɞ�����Y"����ջ�5����h*�0Z���&�z�+��.�e�1�F5�I�:���B��.M���Y��^g���t�����&������s��$熼�{��΃��w���恼�G������y��������m��Y������������������X)���;��I�����!Q��{����	�������뚼P��P���Ϊ���?��\���[�����R���'��C��Μ� x��Y���B¨����'���<���Pȭ�����멼]맼%���*J������ʨ��<������°�����ƴ� ����������	D����e.���G��1m��ǡ������,&ļ3kȼX�˼DGμ�2ϼӹμ�0ͼ.˼�gɼR�ȼ�ȼz�ʼ�μ�CҼ��ּ<�ڼ��ݼ�  �  )&@=��?=�J@=��@=��A=�*B=�[B==B=�vA=t@=7?=��=={�<=z�;=��:=�:=wg:=�q:=��:=��:=rH:=B�9=��8=�7=*V5=�p3=�1=�G0=�g/=3"/=_l/=�0=��0=C�1=߲1=�Q1=�Y0=��.=f-=;R+=��)=m�(=sg(=��(=)2)=�*=Z�*=�+=m�+=��+=+=U/*=�)=Y(=�'=�m&=|&=9�%=��%=i=&=�w&=��&=$5&=�v%=8:$="�"=�| =�P=�==Zt=	=:!=��='=�h=�P=ʓ=5=�=�C
=O=yj=���<���<�h�<��<[��<���<g��<!�<+��<5B�<t�<W@�<��<���<^��<0>�<S7�<彲<���<u�<e�<�r�<���<ܙ<E�<r��<�<]a�<q�t<�j<0�b<�6]<CY<PoU<�.Q<�:K<��B<8<�*<�I<�7<��;Ă�;��;��;Z%�;�>�;�7�;)�;i˛;V��;�x;B�N;��;���:]Ix:�`|9{uֹ�6��\ƺV����J=�0[^�@H���\��%i��M�̻���j��K��E�?2 ��&��X*�R@.���2���8��A�HK��W��{c��{o�}�y�&ŀ�%'�����g���� ��2?��}���������Y턼���1>��a��/d�����<C��猼P<��񏋼F8���~��z���k���
U��D������R���7���K��w1��-��b��(��������q�������ƛ�W�:�������ݨ�ߔ��v�����P��Ӽ��vX��Q������[����@��I���'
���|��~���	*��a+��.�������n��/W�����̴������O��uǽ�����"eż��ȼ��ʼ�˼z�˼��ʼ�gɼ!-ȼ��Ǽy?ȼ.ʼ��̼��м�tԼ�ؼ-�ڼ�  �  zB=��A=g�A=�>B=R�B=U�B=��B=L4B=ʀA=k�@=��?=�i>=+h==��<=�;=8c;=j;=�:=k�:=��:=4R:=\�9=��8=��7=�[6=��4=f3=k02=PY1=��0=E�0=
H1=D�1=�2=_2=e�1=��0=6�/=u.=��,=X�+=Ե*=[Y*=�e*=��*=�A+=E�+=*,=^ ,=g�+=�+=�Y*=�z)=K�(==�'=�M'=��&=�&=�&=B�&=�&=P�&=�;&=��%=ʚ$=v?#=8�!=��=��=_S=u�=�=��=?=��=I�=�=�H=iK=��
=�P=��=� =b��<��<�^�<b[�<��<���<���<���<f9�<'�<��<}��<J�<�s�<��<��<O�<��<�ի<�ҧ<��<�K�<.|�<7�<k��<���<޾�<��|<d�r<׈j<T�c<�<^<�Y<cS<rL<`�C<�9<d�,<�s<�<�<���;���;�>�;���;[B�;/�;��;��;3o�;:+y;��P;��$;�:���:��9�0���H��W��O��d�9�=�[�,n����z��ȾûD�ܻ^n��4%�99�����In%�v�*�3�0��7��?�ǗI�cMT�rZ_��i���r�*�y��p~��o�� ̀�V����_��vU��M���Q���3킼6����^�����釉�l���1X��氋����Ex��m0��h�� f���@��黍��Џ��W������r���V�� v�������;��RH��N������u㗼��ך��k��"P������J��U����D����&l������1���4़�]��x��r��M���-��H2��<���D`���q���)������|ϳ����뗴�h������H��� ����y$¼�ļ��Ƽ<)ȼ�ȼ�6ȼ�Ǽ`Ǽ��Ƽt�ǼIZɼ`�˼�μ��Ѽ��Լ��ּ�  �  �C=�C=�eC=HKC=�'C=3�B=�vB=j�A=^(A=�Z@=`�?=Q�>=��==iN==��<= <=�;=F$;=��:=�`:=]�9=�u9=f�8=�8=�7=��5=h�4=��3=X-3=W�2=�`2=O2=T2=�L2=�2=�1=I�0=��/=��.=�-=m-=��,=*,=�,=,=D(,=�,,=�,=��+=BX+=��*=�3*=��)=8)=$�(=�(=Y�'=nR'=�'=��&=��&=$:&=��%=R%=9�$="�#=�d"=2!=8�=,=��=4O=&=/�=3`=U�=��=�9=2j=�V=%'=�=�=C��<V�<N>�<���<���<9�<aC�<���<�a�<��<�k�<�=�<X�<���<Կ�<k��<Q��<nİ<��<���<�6�<�Ϟ<�O�<���<�Ȑ<j��<殆<���<�7z<��q<��i<��b<d�[<��T<��L<�C<�D9<+�-<�!<��<�
<�S <t��;�;�;���; �;�h�;��;�;9��;Q�s;�rM;�%;Zt�:'�:0:�b86������� �y\�P;�	_�﹁�ʚ���k���@����һR�������w�����U!��$(��T/�7�l�?���H��RR���[�+�d��hl���r�zw�	.z��2|���}��~�#4��&��G��Ȋ��hۄ�� ��]D���;����C����Z��Պ�O,���m����q�� ���۵��z���"q��W5��J���Tؖ��y��򤗼����?M��P�����Ę��P���A���Y���Q��������������	�����)c��`���O𥼲.��ã���3������A7��O����į��鰼�����岼ܴ��Mv���D��"=��cx�� ��麼���S��qu��8EüȠļ1zż�ż�Ƽ�8Ƽ�Ƽ�Ǽ�ɼq˼4]ͼ3�ϼ��Ѽ�{Ӽ�  �  �XE=��D=(^D=��C=m5C=<�B=��A=�A=�O@=�?=G+?=`�>=�G>=��==n@==�<=��;=�;=tR:=B�9=�9=P�8=1+8=�7=c77=s�6=��5=G5=��4=��3={r3=?3=G�2=OI2=S�1=zg1=
�0=1'0=�|/=��.=�W.=!�-=S�-=4=-=��,=��,=B,=��+=��*=�v*=� *=��)=sY)=�)=X�(=�(=�:(=��'=�"'=t�&=�%=�l%=��$=�|$=��#=�f#=z�"=�!=�� =X=��=�v=\�=X:=�o=�x=!I=~�=|8=Zt=�=u�=E=�� =��<�+�<ݩ�<*"�<���<7��<~(�<��<���<�h�<���<t�<8��<���<�Ȼ<k�<��<���<���<T��<BC�<��<���<��<?݌<֨�<[�<� �<Lw<��n<�"f<
�]<��T<��K<�VB<�28<��-<d#<�</�<�T<p0�;���;˝�;W��;�F�;_`�;F�;���;W�e;}C;�� ;,��:�7�:i�V:�_f9l�عKF��[�⺴��`1D��lj�GM������>��������̻9T߻�4�-�����+����&��//��7��U@�^I���Q��Y���`��\g�x�l�Bdq�tKu� �x�� |��6��/���������������ԗ��G���t��E�_���n�������o���|��[C��ݍ�QY���͎�,R������Eݐ�㑼<���,��#��������]��S떼h����<��<5��Nf��뷛��	���A���P���7������̡�h�������㤼6:��Ś��#�t��8"��� ���̬�����6����߯��N���ֲ��W��4��������"��Ṽ-麼r��$y������r������}"ü�9ļ(,ż�Ƽ��Ƽoȼ�tɼ8�ʼ��̼μ��ϼR�м�  �  �5F=$�E=��D=M�C=��B=��A=�v@=D�?=]�>=ْ>=Cg>=W>=Y?>=a�==c�==D�<=
�;=��:=�x9=`z8=��7=�47=�6=U�6=M�6=�6=�k6="6=zy5=��4=4=�N3=2=�1=�]1=��0=�^0=9�/=�/=�Z/=h/=��.=�a.=��-=�#-=�J,=[+=o*=Ƣ)=)=Z�(=ҝ(=r�(=-�(=��(=V�(=�t(=k�'=��&=��%=L�$=^!$=b�#=M#=��"=ǖ"=N"=��!=G!=� =��= !=�K=xI=l&=Q�=`�=,=ٲ=�7=��=�W=/�=�=�	�<Y��<��<W�<u��<�@�<N4�<ڐ�<�^�<,��<w��<h,�<��<�<2I�<Y��<�z�<�a�<<��<�B�<9��<ᖖ<1�<,�<���<pj�<�ƅ<�Ł<s�z<}q<S�g<�]<,�S<��I<��?<��5<�,<�"<̤<��<vH<)8�;�b�;���;_�;@�;�	�;�o�;�r;�1P;�r1;(�;���:���:��h:ڡ9�
���䊺Ҟ캙�&�8�T�\'~�,`��sx����������-�˻r�ڻ��뻜����j��r�>���&�y^0� 9��iB�ץJ��0R���X��^�=d��/i�h�m���r�*�w���|������]��o[��ӆ�?��������؇������U���~���*��)]��s�������gq��Ώ�\���1�����\ِ�������������Z���C��dj��������;��}W��*Y���H��i$���㛼�������Ų��v���z���Ѡ�����?|���-���uf����������h물���#���a���%���x��fO�����1ɵ��巼����Ժ�f�����W#��=^��[ռ�Ɵ��S����$��»��güżΑƼ�Ǽ�?ɼ�sʼ"�˼,�̼A_ͼ�-μ�ϼ�  �  �F=J�E=�D=!C=��A=;@=�>=��==j7==�==�N==��==!�==d�==s==�<=VR;=��9=�H8=��6=)�5=�a5=�=5=m5=��5=�"6=�O6=C76=��5="#5=�>4=N=3=�;2=U1=�0=v
0=��/=^|/=&o/=lo/=�_/=P$/=��.=n�-=��,=S�+=�#*=n�(=�'=�8'=<	'=B'=g�'=�N(=��(=W�(=�a(=/�'=�a&=��$=R�#=rx"=Ϫ!=�@!=�*!=�H!=�l!=�e!=)!=�= =D�=�S=L=v=�=�=K�=�@=�=��
=m�=�]=�=��=@:�<ŉ�<�m�<n�<?��<"��<lk�<w��<�<�<�6�<sF�<���<�r�<�,�<a�<FU�<1q�<�ۡ<H�<! �<�?�<�:�<YǍ<D��<��<q�<�r�<�J|<�{r<��g<�\<9pQ<��F<ZB<<*�2<[�)<S!<�4<c<	D	<�� <���;���;���;�0�;��;$�z;&|T;f4;U';��;B��:��:'�f:l
�9����L���v �t7��k���������񭻇���Ļ'2ϻ:"ۻ�b�LG�����{�Z����'�$�2��<��wE�OIM�;�S���Y��p^���b��g�C�l�~r���x�I���b���y���戼q�����;����������KӇ�^����K��'Ή�d��C���E�����Q��{����K��l^��M<��oB����� Ր�K����ђ��{��kT��Y ������O��؛��h��\���z����Ĝ�N���Ý��������^r��7V��WL��/����	��
N�������`��l����������B������d� ʴ��ⷼ�ĺ�}���|��h��s�va�������N���h������o��J=���Zü��ż8�Ǽ	lɼ��ʼ��˼?�̼1ͼQbͼK�ͼ#Zμ�  �  YqF=kE=s�C=�,B=Q:@=�_>=��<=��;=I_;=�;=<=��<=a^==x�==�.==7<=4�:=x�8=�6=.F5=�4=rn3=�c3=�3=܅4=�D5=��5=C�5=��5=�5=�4=��2=��1=ė0=�/=�%/=��.=��.=/=|8/=XL/=�/=4�.=K�-=�,=�m*=��(=�'=��%=�I%=�B%=��%=��&=�'=�>(=�v(=�(=� '=2�%=��#=�*"=b� =��=!J=�X=��=!? =�� =X� =� =8�=v,=G=_�=��=�5=ܧ=�B=�=�
=c===�=^�=��<�l�<I��<�t�<)m�<��<�f�<'��<��<�8�<�4�<��<�	�<B��<��<�"�<Cϭ<�.�<�<�<a�<%��<��<1�<��<��<���<�H�<.|<r<��f<��Z<ӓN<�C<�n8<q�.<fd&<a�<�<n�<�<l��;��;�|�;9��;[�;QA�;�\;Y5;V�;�� ;�I�:Q|�:}�:�W:�9�ٹ.4����k�J��Ł��0����I任"0ƻ�
λyջD�޻���V��������_���)�3n5��?�7�H��dP�aV��"[�6/_�^+c���g��(m���s���{�����G�����������H����������H���� ��k���.7��tڈ�c���k��*���F���w���.)��@���Qޗ��_���������چ���#��.����󒼅ߔ� ���Y��>G�����&����일�ʝ��h��"��D'��᝼�o���ࡼ����Ũ��r��J����:��������ܟ���;���~��̮��L�����o���H���ὼа��a¼��¼W\¼V'������c������DT��`����o����ü�~Ƽ��ȼ�˼��̼2�ͼdμ�μt�ͼ{�ͼ	nμ�  �  �#F=��D=�BC=�*A=T�>=��<=�%;=�:=J�9=+:=B�:=��;=3�<=�'==_�<=��;=�:=�7=��5=��3=Eg2=��1=ҷ1=Q2=-H3=�T4=�+5=֔5=�w5=!�4=��3='~2=� 1=��/=]�.=�W.=.= 9.=��.=��.=/=�.=8..=�,=�O+=�Q)=�G'=�}%=�3$=��#=y�#=Fr$=�%=�&=�'=�(=ϻ'=�&=��$=��"=�� =�&=�=��=8�=J=�=Ĺ=��=V�=B�=�=~�=��=m,=kd=u�=a=�?=�U	=f�=˯=֟=�4=��<��<���<���<]�<!��<C��<j��<��<��<�N�<l��<+�<�N�<V�<��<4J�<C�<�:�<�h�<��<�F�<j�<z��<���<?{�<��<���<B1{<	�p<>#e<~X<<�K<��?<�5<��+<lx#<p<5�<�.<�<���;L��;�t�;�U�;bW�;Q]q;�@;	{;�$�:�2�:�̽:��:"!�:ӚA:�W`9_��zh��f��7K\�i���߭��������Ȼ �ѻ�n׻v�ܻuB�ǐ�OD��������w[�A,��8�,�B��L��HS���X��\��`��$d���h�dqn�>�u��~�&B���	���(���$������̥���E�����򛋼����񈼩���X����׎�/�������������� �����`7��#Ȗ��g�������ۑ��)���y�����������������R��l/���X��p���jI��Ÿ��2���zm��n:�����V榼�0���e�����b�� o���������s��I���Xb��~�����C�����I}������]�ü��ż�IƼ{ż�ü����z�������������%�����ļڇǼzNʼ>�̼�Eμ"/ϼ~jϼ4(ϼW�μ�μ�μ�  �  ��E=��D=��B=dg@=��==ƻ;='�9=M�8=w�8=o 9=`#:=�W;=4[<=��<=ˎ<=Us;=��9=bS7=D�4=�2=�F1=]�0=(�0=v@1=�_2=��3=+�4=y45=D.5= �4= �3=�$2=��0=	e/=d.=*�-=��-=-�-=�%.=ۍ.=*�.=v�.=-�-=��,=&�*=1~(=mG&=�\$=�#=xl"=��"=��#=��$=�C&=�X'=��'=]q'=�B&=�i$=u0"=@�=�=^�=Y=͊=~@=�2=�=�v=\9=�<=߈=_>=��=�=}�=�(=K�=+�
=��=\=zW=PP=y� =m��<G��<�1�<�<Y3�<�+�<Oo�<[;�<ׇ�<$��<m��<w��<�{�<Tſ<�W�<�R�<o,�<r��<8d�<tI�<�Í<��<�<���<��<�S�<gɃ<�<�!z<�o<��c<�V<(�I<x�=<�2<hG)<�d!<��<n<��<{V<��;�l�;���;P�;á�;��_;"�-;ܢ;{��:��:��:ER�:E0�:�/:;�$9d+�����o�#�u�h��N��wB���û��ѻ��ٻ0g޻8��jD�Ma��b��������� �Ŭ-��:��E��4N��TU���Z�6x^��a��(e�k�i���o���w�/����ㅼ����f����������ē�����{��������������#���]��X叼"���T�������ٝ��_��%e��z@���y��5�������*���˴������*��kΘ��z��_ɝ�do���I��\��ӟ�� ���O���/�� ���W���� ��;K��i���T��[B������-�������G��lճ�8�����������ⴼ�8�����¼�Ƽ�(ȼu�ȼ��Ǽ��ż�]ü�0���п�+���ϊ��>�¼�Gż�TȼYB˼Z�ͼ�cϼ�CмZbм��ϼeeϼ<ϼPtϼ�  �  V�E=�dD=�xB=�@=�==�V;=��9=D~8=TA8=��8=��9=a;=�1<=[�<=�s<=cR;=r9=p7==�4=s2=��0=�0=�#0=��0=.
2=�W3=�o4=�5=(5=0x4=d3=�2=ߊ0=�6/=2.=j�-=Uh-=�-=O .=�m.=ݦ.=�v.=,�-=�Z,=�p*=�/(=�%=�#=o�"="=$A"=�5#=��$=�&=O3'=ɯ'=�T'=x&=�7$=��!=g�=��=�o=��=� =�=��=��=�D=2=(=�h=#=�c=�}=��=)�=�=�}
=«=��=6=�1=�� =-��<9��<��<�h�<�n�<qV�<t��<�l�<���<�_�<�z�<FX�<v9�<���<��<��<�ª<0�<���<܅�<W��<�"�<i�<��<�{�<�ބ<�q�<�̀<9�y<�Wo<~=c<�1V<�I<T�<<��1<{w(<~� <<R�<�o<��<��;��;y��;6˨;���;�sY;!)';N ;���:3��:([�:Ь�:��x:"):}p9�X���ƺ�{'�3m�	���Z���ƻ,�Ի��ܻ�ở他������S��&	����;!�O.���:���E���N�!V�B[�X
_��/b���e�j��5p��Ux�����~�����5��(W���͔����ܻ�����p���ʊ�����[�����%H������
���A��0����7��n6������(���4������/ϒ��:���i�����Л�)���ԟ���������%��G��]����g��X8���>������>Ѩ�˞��=B��|������c���LԸ�T㶼�P���ⱼ Y��E���챼3�����𕾼�9ü��Ƽ��ȼ}ɼ��ȼFvƼ��ü�����%��tԿ�<�����¼�ż�ȼO�˼�μ}�ϼ��м~�мHм��ϼ�Oϼd�ϼ�  �  ��E=��D=��B=dg@=��==ƻ;='�9=M�8=w�8=o 9=`#:=�W;=4[<=��<=ˎ<=Us;=��9=bS7=D�4=�2=�F1=]�0=(�0=v@1=�_2=��3=+�4=y45=D.5= �4= �3=�$2=��0=	e/=d.=*�-=��-=-�-=�%.=ۍ.=*�.=v�.=-�-=��,=&�*=1~(=lG&=�\$=�#=wl"=��"=��#=��$=�C&=�X'=��'=Yq'=�B&=�i$=m0"=6�=�=Q�=�X=��=o@=�2=�=�v=f9=�<=�=�>=6�=�=��=�*=��=��
=��=3#=�[=U=�� =7��<{��<"=�<�<�>�<�6�<oy�<�D�< ��<�<���<W��<�}�<�ſ<bV�<�O�<�'�<G��<�\�<�@�<���<��<겇<N��<`�<kH�<Ⱦ�<�<�z<��o<s�c<��V<�I<��=<Ū2<�J)<ak!<��<�z<E�<th<�C�;u��;���;|>�;Ќ;�`;".;��;���:�$�:fz�:Y��:�f�:�0:��$9�i�x����*$��h��o���h��?�û%�ѻx�ٻ�޻P/��t�2�𻓏��ݳ����� ���-��:��E��=N�`\U���Z��|^�n�a�t+e�S�i��o���w�����4䅼-���f��1��������ē����	|������%��������#���]��Z叼"���T�������ٝ��_��%e��{@���y��5�������*���̴������*��kΘ��z��_ɝ�do���I��\��ӟ�� ���O���/�� ���W���� ��;K��h���T��[B������-�������G��lճ�8�����������ⴼ�8�����¼�Ƽ�(ȼu�ȼ��Ǽ��ż�]ü�0���п�+���ϊ��>�¼�Gż�TȼYB˼Z�ͼ�cϼ�CмZbм��ϼeeϼ<ϼPtϼ�  �  �#F=��D=�BC=�*A=T�>=��<=�%;=�:=J�9=+:=B�:=��;=3�<=�'==_�<=��;=�:=�7=��5=��3=Eg2=��1=ҷ1=Q2=-H3=�T4=�+5=֔5=�w5=!�4=��3='~2=� 1=��/=]�.=�W.=.=�8.=��.=��.= /=�.=7..=�,=�O+=�Q)=�G'=�}%=�3$=��#=w�#=Cr$=�%=�&=�'=�(=ƻ'=ݣ&=��$=q�"=p� =�&=�=�=�=�I=l=��=��=j�=�=��=S�=��=Y.=g=��=�e=�D=\	=Ώ= �=��=�>=���<N#�<���<� �<�r�<���<���<B��<ש�</��<Y�<��<A/�<�O�<��<��<AA�<_�<�+�<#X�<���<2�<#҉<�r�<���<�e�<���<���<\{<p�p<�	e<�jX<u�K<v�?< 5<��+<:�#<�<'<(M<Ĩ<��;D9�;���;뮱;䰔;�r;�TA;p;h?�:�(�:E��:�|�:���:c B:$2`9 `�۴����w�\���������n���i�Ȼ3�ѻf�׻f�ܻ��z�����������|��%,�78��C��L�CWS� �X�-]���`��)d�F�h�0tn�Y�u���~��B��e
��?)��%��򫑼󥑼�E������������"񈼰���^����׎�2�������������� �����a7��#Ȗ��g�������ۑ��)���y�����������������R��l/���X��p���jI��Ÿ��2���zm��n:�����V榼�0���e�����b�� o���������s��I���Xb��~�����C�����I}������]�ü��ż�IƼ{ż�ü����z�������������%�����ļڇǼzNʼ>�̼�Eμ"/ϼ~jϼ4(ϼW�μ�μ�μ�  �  YqF=kE=s�C=�,B=Q:@=�_>=��<=��;=I_;=�;=<=��<=a^==x�==�.==7<=4�:=x�8=�6=.F5=�4=rn3=�c3=�3=܅4=�D5=��5=C�5=��5=�5=�4=��2=��1=ė0=�/=�%/=��.=��.=/=|8/=XL/=�/=4�.=K�-=�,=�m*=��(=�'=��%=�I%=�B%=��%=��&=��'=�>(=�v(={(=� '=�%=p�#=�*"=C� =ٸ=�I=�X=z�=�> =�� =S� =� =��=+-=|=A�=~�=�9=Ԭ=I=S=�

=�=#==W�=���<Y��<���<��<܋�<��<B��<[�<A��<KK�<RC�<�	�<��<���<���<��<�­<��<�Ϟ<�i�<�F�<�x�<�Ԍ<L �<�<�ȇ<wl�<�-�<��{<��q<ؐf<��Z<]�N<eC<'n8<3�.<}v&<^�<��<�<J�<�
 <�t�;��;�6�;��;m��;Q�\;X�5;�;7�;�h�:[X�:3}�:ڪW:y�9�۹�գ�^��4K�� ��?���@���~`��o�ƻ<�λ��ջ�
߻��������v���*��5�m�?�KI�yP�qV�/[��8_��2c���g��,m���s�ӣ{����TH��'���
���8I��׉��ޡ��h���	!��}���;7��~ڈ�k���k��/���I���z���0)��B���Rޗ��_���������ۆ���#��.����󒼅ߔ� ���Y��>G�����&����일�ʝ��h��"��D'��᝼�o���ࡼ����Ũ��r��J����:��������ܟ���;���~��̮��L�����o���H���ὼа��a¼��¼W\¼V'������c������DT��`����o����ü�~Ƽ��ȼ�˼��̼2�ͼdμ�μt�ͼ{�ͼ	nμ�  �  �F=J�E=�D=!C=��A=;@=�>=��==j7==�==�N==��==!�==d�==s==�<=VR;=��9=�H8=��6=)�5=�a5=�=5=m5=��5=�"6=�O6=C76=��5="#5=�>4=N=3=�;2=U1=�0=u
0=��/=^|/=&o/=lo/=�_/=O$/=��.=m�-=��,=R�+=�#*=m�(=�'=�8'=9	'=�A'=a�'=�N(=��(=K�(=�a(=�'=�a&=��$=2�#=Mx"=��!=Y@!=Z*!=NH!=�l!=ie!=$!=�= =��=�T=�M=�=k�=5!=c�=�H=s�=ӻ
=;�=l=�/=��=�^�<j��<��<�5�<���<;��<=��<F��<'8�<��<�H�<ES�<���<Ft�<�(�<p�<�E�<�\�<�¡<7�<���<��<��<{��<E^�<[�<��</Q�<|<�Fr<��g<�z\<kXQ<�F<hA<<ߔ2<z�)<V@!<�_<h�<N�	<r� <�Q�;�2�;�n�;H̪;Չ�;��{;y�U;�Y5;C�;�;���:Ǯ:ͨg:��9����_q����,8� �k�l���n�����2���mRŻ�ϻ��ۻB �%���t�-������(��2�5�<���E�4bM��T�Y�Y��|^��c�̨g�F�l�݁r���x�i��Sc���z��B爼`q�����n���<���å��aӇ�o����K��0Ή�k��I���I����� Q��}����K��m^��N<��oB�����!Ր�K����ђ��{��lT��Z ������O��؛��h��\���z����Ĝ�N���Ý��������^r��7V��WL��/����	��
N�������`��l����������B������d� ʴ��ⷼ�ĺ�}���|��h��s�va�������N���h������o��J=���Zü��ż8�Ǽ	lɼ��ʼ��˼?�̼1ͼQbͼK�ͼ#Zμ�  �  �5F=$�E=��D=M�C=��B=��A=�v@=D�?=]�>=ْ>=Cg>=W>=Y?>=a�==c�==D�<=
�;=��:=�x9=`z8=��7=�47=�6=U�6=M�6=�6=�k6="6=zy5=��4=4=�N3=2=�1=�]1=��0=�^0=9�/=�/=�Z/=h/=��.=�a.=��-=�#-=�J,=[+=o*=â)=)=U�(=̝(=k�(=$�(=}�(=I�(=�t(=W�'=��&=��%=(�$=5!$=3�#=#=��"=��"=�M"=��!=E!=� =3�="=�M="L==*=��=.�=�4=N�=�C=��=h=� =2�=2�<e�<���<)G�<k��<�h�<�Y�<&��<�|�<���<���<�:�<�"�<3��<wD�<L��<�i�<�J�<bs�<�"�<x�<�o�<�<붏<���<�@�<��<���<׍z<�Aq<��g<��]<��S<��I<��?<��5<T3,<��"<��< <��<���;��;�w�;*�;h�;R��;��;3s;BAQ;�^2;�;	�:�h�:�^i:���9�׶� ��� ��ޢ'�i�U�]C������!��訰��u��K�̻)�ۻ�<��:��Ÿ�]�������&�o�0�2�9�H�B���J��FR��X�d�^�)Gd�^7i��m��r�^�w� �|������^���[���ӆ���������؇�����U���~���*��4]��{�������lq��
Ώ�^���3�����^ِ�������������Z���C��dj��������;��}W��*Y���H��i$���㛼�������Ų��v���z���Ѡ�����?|���-���uf����������h물���#���a���%���x��fO�����1ɵ��巼����Ժ�f�����W#��=^��[ռ�Ɵ��S����$��»��güżΑƼ�Ǽ�?ɼ�sʼ"�˼,�̼A_ͼ�-μ�ϼ�  �  �XE=��D=(^D=��C=m5C=<�B=��A=�A=�O@=�?=G+?=`�>=�G>=��==n@==�<=��;=�;=tR:=B�9=�9=P�8=1+8=�7=c77=s�6=��5=G5=��4=��3={r3=?3=G�2=OI2=S�1=zg1=
�0=1'0=�|/=��.=�W.=!�-=S�-=3=-=��,=��,=@,=�+=��*=�v*=� *=��)=lY)=�)=M�(= �(=�:(=��'=�"'=U�&=��%=jl%=��$=�|$=��#=�f#=I�"=Ź!=�� =>X=T�=�w=4�="==�s=c~=/P=`�=OC=-�=��=�=xW=�� =���<�W�<=��<N�<a��<��<qO�<k��<	�<Ԃ�<��<Ղ�<���<O��<Ļ<�_�<l�<��<�n�<㝡<��<\��<d͔<1ǐ<N��<�}�<�1�<K�<kw<pnn<��e<@u]<)�T<�K<�UB<�>8<?�-<�(#<��<��<P�<\��;�J�;�L�;�V�;��;��;���;>!�;�	g;D;�a!;�*�:��:�OW:@f9��ڹ�(���Ԏ��0E���k����\���y��Ļ�I�ͻ�������oP�0u��O���&�b/���7��y@�H%I���Q��Y��a��gg���l�Ijq��Ou���x�Z|��8��0��2�����S��6������i���t��Y�n���y�������v������_C��ݍ�SY���͎�-R������Eݐ�㑼<���,��#��������]��S떼h����<��<5��Nf��뷛��	���A���P���7������̡�h�������㤼6:��Ś��"�t��8"��� ���̬�����6����߯��N���ֲ��W��4��������"��Ṽ-麼r��$y������r������}"ü�9ļ(,ż�Ƽ��Ƽoȼ�tɼ8�ʼ��̼μ��ϼR�м�  �  �C=�C=�eC=HKC=�'C=3�B=�vB=j�A=^(A=�Z@=`�?=Q�>=��==iN==��<= <=�;=E$;=��:=�`:=]�9=�u9=f�8=�8=�7=��5=h�4=��3=X-3=W�2=�`2=O2=T2=�L2=�2=�1=I�0=��/=��.=�-=l-=��,= *,=�,=,=C(,=�,,=�,=��+=?X+=��*=�3*=��)=/)=�(=~(=H�'=ZR'=�'=h�&=��&=�9&=d�%=�Q%=�$=�#=Yd"=!==�=j=D�=OP=�=��=d=��=ɱ=~B=�t=(c=t5=�=f-=��<�~�<jh�<y��<X�<�b�<�k�<�!�<���<���<?��<�Q�<��<���<���<���<N��<b��<�<؁�<��<x��<�(�<�|�<���<���<5��<���<3�y<�lq<F�i<?�b<��[<9�T<ҼL<��C<�P9<��-<�"<�<��
<l� <IR�;7��;�D�;0��;!�;��;���;^6�;�t;�]N;�&;���:��:��0:��`8��2_���=�5)��F<�Q-`�W��D��~�������ӻR:�{3��������@���W!��](�݅/��67�ӧ?���H��hR� �[���d�-sl���r�fw�x2z�36|��}���~��4���&��G������ۄ�� ��~D���;��(��Q����Z��Պ�U,��n��񳋼t��"���ݵ��{��𣐼#q��X5��K���Tؖ��y��򤗼����?M��P�����Ę��P���A���Y���Q��������������	�����)c��`���O𥼲.��ã���3������A7��O����į��鰼�����岼ܴ��Lv���D��"=��cx�� ��麼���S��qu��8EüȠļ1zż�ż�Ƽ�8Ƽ�Ƽ�Ǽ�ɼq˼4]ͼ3�ϼ��Ѽ�{Ӽ�  �  zB=��A=g�A=�>B=R�B=U�B=��B=L4B=ʀA=k�@=��?=�i>=+h==��<=�;=8c;=j;=�:=k�:=��:=4R:=\�9=��8=��7=�[6=��4=f3=k02=PY1=��0=E�0=
H1=D�1=�2=_2=e�1=��0=6�/=u.=��,=X�+=Ե*=[Y*=�e*=��*=�A+=C�+=(,=\ ,=d�+=|+=�Y*=�z)=C�(=3�'=�M'=��&=�&=��&=(�&=ͣ&=+�&=�;&=��%=��$=G?#=�!=��=��=�S=�=�=J�=�='=��=4�=ZP=�T=�
=�]=U�=� =ѷ�<,�<���<΁�<A��<>��<}��<@��<X�<B�<���<o��<
!�<�z�<j�<a�<#E�<��<���<Ĺ�<���<�+�<FY�<M�<�b�<�u�<}��<�9|<J�r<�Kj<�c<Y^<��X<KS<heL<l�C<�&9<��,<�<e<B<��;
y�;���;[Z�;�ݽ;-ʴ;���;��;���;�z;D�Q;��%;�:�_�::�9��0���I�����k�E��Wr:���\��������6���bĻiyݻ���Ut����c��O��)�%�q+�6�0�=�7��@��I�zaT�Ej_�P�i��r�Q�y��u~��q���̀�y����`��V��ʸ������y킼k����^����� ���~���>X��𰋼���Jx��q0��k��#f���@��껍��Џ��W������r���V�� v�������;��RH��N������u㗼��ך��k��"P������J��U����D����&l������1���4़�]��x��r��M���-��H2��<���D`���q���)������|ϳ����뗴�h������H��� ����y$¼�ļ��Ƽ<)ȼ�ȼ�6ȼ�Ǽ`Ǽ��Ƽt�ǼIZɼ`�˼�μ��Ѽ��Լ��ּ�  �  )&@=��?=�J@=��@=��A=�*B=�[B==B=�vA=t@=7?=��=={�<=z�;=��:=�:=wg:=�q:=��:=��:=rH:=B�9=��8=�7=*V5=�p3=�1=�G0=�g/=3"/=_l/=�0=��0=C�1=߲1=�Q1=�Y0=��.=f-=;R+=��)=l�(=rg(=��(=(2)=�*=Y�*=�+=k�+=�+=+=Q/*=�)=S(=�'=�m&=p&=*�%=��%=T=&=�w&=�&=5&=�v%=:$=��"=z| =�P=>=�t=}="=6�=(=�k=�T=ɘ=�"=��=�L
=�Y=Uv=��<��<���<�4�<���<���<���<m!�<���<1[�<w+�<�R�<l�<��<H��<o?�<�3�<ѵ�<[��<���<�P�<O[�<j�<���<K�<�}�<ˆ<�B�<פt<>�j<[�b<R]<��X<�RU<�Q<30K<��B<�8<U+<�d<l[<�\�;���;���;Rb�;-��;d��;W��;�l�;JA�;�b�;�ny;FeO;�~ ;���:\ny:F�~9֏ֹ���M�ƺ�V�ޣ���=�.*_�ﺂ�wؘ�뱻�>ͻ�W�	0��V�J���k ��6&�Q�*�j.���2�99��7A��\K��W���c��o�<�y�Ȁ�])��x �����������?��������4���턼��J>��t��=d�����EC��%猼U<������I8���~��{���l���U��E������S���7���K��w1��-��b��(��������q�������ƛ�W�:�������ݨ�ߔ��v�����P��Ӽ��vX��Q������[����@��I���'
���|��~���	*��a+��.�������n��/W�����̴������O��uǽ�����"eż��ȼ��ʼ�˼z�˼��ʼ�gɼ!-ȼ��Ǽy?ȼ.ʼ��̼��м�tԼ�ؼ-�ڼ�  �  m>=/I>=��>=��?=�@=�yA=5�A=�A=�6A=)@=J�>=^==�<=��:=�,:=j�9=��9=4�9=,:=,D:=�:=�T9=8=Y^6="G4=�2=�0=y�.=I�-=k�-=�.=�/=0=��0=�Q1=j�0=�/=y6.=d(,=�*=�N(=�!'=��&=P�&=�'=z�(=k
*=L�*=�n+=�_+=��*=��)=խ(=�v'=�g&=��%=�8%=�)%=de%=C�%=�$&=�B&=��%=e%=ӭ#=�!=�\=��=��=��=�r=ڪ=�Q=%=*�=��=�S=:�=�=��	=�b=5=���<��<�=�<;$�<�%�</��<�D�<�-�<��<���<���</��<"�<7��<�M�<l��<K��<@�<��<��<���<)��<5�<X̘<��<'�<�4�<
[z<��m<Ĥc<)&\<�<W<&5T<��Q<O�N<{�I<��A<M�6<��(<3=<�	<|�;#a�;�<�;�Q�;Z��;é;K�;��;�ʘ;�
�;�Wu;�uJ;��;��:Z�J: #8N#�,O��#q޺��_'�b�C�A�d���b��~���3ֻ������ X����H�&���+���.���1��85�ѱ:�d�B�I=M�~�Y�hg���t����(�������t��膼�|���΃�6x���恼-H��
������������m��f������������������[)���;��K�����"Q��{����	�������뚼P��P���Ϊ���?��\���[�����R���'��C��Μ� x��Y���B¨����'���<���Pȭ�����멼]맼%���*J������ʨ��<������°�����ƴ� ����������	D����e.���G��1m��ǡ������,&ļ3kȼX�˼DGμ�2ϼӹμ�0ͼ.˼�gɼR�ȼ�ȼz�ʼ�μ�CҼ��ּ<�ڼ��ݼ�  �  �>==$==��==��>=��?=��@=E�A=�A=��@=��?=�y>=@�<=;=�a:=�9= D9=�G9=׉9=R�9=�9=D�9=�9=�7=��5=�{3=C1=!�.=4d-=��,=t,=�-=�A.=��/=ݏ0=�1=)�0=�/=��-=�z+=�5)=�G'=��%=~%=��%=N�&=��'=�Z)=Pv*=z+=�+=��*=�)=mQ(=�'=��%=�%=V�$=��$=��$=�k%=�%=@&=L�%=b�$=t6#=�!=̆=��=m�=F�=CU=��=�z=�}=�S=۞=�=��=M7=!	=��=/V =g��<0��<V��<O��<�:�<�(�<��<�T�<�}�<�g�<�(�<��<]�<j��<�;�<Vt�<�r�<7�<䚬<oR�<D��<�+�<���<���<�_�<v��<sU�<kv<�#i<��^<��W<�GS<a�P<�^O<��L<0rH<w�@<��5<kI'<.�<��<H��;���;1�;
0�;�B�;�m�;,�;���;^��;u��;Xq;�E;c�;3��:��):R׸,�I�ۯ�'�(	��-�	�H�F�i��̈�)&��������ܻ1���F?�`(�xI$��Y+�q�/��2��
4��6���;���C�^�N���[��&j��x�����u��{���Ɖ����BB��]1��k{��I����؂����c/��b����O��"�����D֏�)�G��N獼K׌�%E�� ������ ���^����������$����	�������U��Hh���������>��]����ښ�\���񔡼�+������'���R��7谼����������)���~���寮M���^U���ޫ�Qͮ�I���$��u䵼�Զ�b�����������~���N���6ܶ��1��۵��i&��k�ż4�ʼ^Eμ��м2qѼ��м�μ't̼�Tʼ/-ɼ�~ɼ�y˼��μ
Ӽ�]ؼC�ܼL+��  �  �+=�J+=��,=l)/=��1=�4=��6=8=O~8=�8=s7=�5=�l4=�M3=��2=�12=6.2=S2=d2=B2=}-1=Rg/=��,=�9)=#H%=	[!=��=�=�=��=f�=�=��!=��#=f2%=�%=i#=�� =�=�_=9G=I=ٴ=�=Ζ=�_=0i=�1=gP!=��"=��"=}"=��!='� =��=��=`k=�u=�=�(=y\=�=�==Z-=_|=Of=6e=�	=�=?H=�M=�E=U�=��	=�
=%�=QQ=�=]o�<kw�<+��<���<��<�Z�<]��<ha�<^�<��<��<��<�"�<[�<*�<��<�F�<�ʱ<)ԫ<잦< &�<,�<_P�<5�<���<��<ki�<!�q<�d\<��F<�2<kT"<l�<ŧ<^�</�<I�<g\<�I<��<5<<O��;�I�;`��;��E;�Y ;��:q�k:�Th:��:�m�:�:�b�:ZL�:.��:��:��9?����[��n���.�+�	�R�4�t�6����a���H��ğ���޻a� �6�0r+�H�A�~�U�.�e���p��Rv�I�v��at�Q#q�.�o�Dr�#z�����}S���C�����^{��`X��@��ݡ��?���'���<=���������ȗ�0��<�������ٛ�HΝ��7���֟����잼���{���ܝ�����Y��
Ө����>M������u_ļ��Ǽ�ȼ��ƼR�¼�������
������HJ���Y�������ļd̼v�ѼT�Լ�Bռ��Ҽ�lμ��ȼü�0��eں��[�������5��9����6����¼ZPļ�=żDoż�0żd�ļ<ż7�Ƽ�ɼlpμ��Լ^�ܼ���b/���x���T��D�򼆃�]L�ۗ�p�ἶ>ἄ���輟�����m�������  �  u�+=H,= q-=~�/=2h2=��4=�7=[@8=�8=�$8=%7=��5=�4=�{3=
�2=�^2=�S2=�o2=�z2=a/2=�G1=[�/=��,=��)=��%=Q�!=&�=�K=�>=O�=0=2�=)-"=mS$=�z%=xL%=��#=P� =�|=��=�=� =�q=�D=i9=�=��=4{=�!=�"=&�"=6�"=r�!=�� =��=��=��=�=�=�B=3q=$+=d+=E=�q=��=��=v= �
=i9=��=*�=/�=j	=�(
=�]
=?	=k�=e=]'�<-`�<z��<��<xK�<D��<)
�<���<�H�<�J�<���<$Z�<<O�<�|�<<<�<Z�<Ҍ�<�"�<	7�<�<\}�<Ut�<ɋ�<jN�<�7�<�Ҋ<�<�r<;<^<�'I<q�5<8L%<<�<8�<�^<��<�e<�<�m<1�<dR<
$�;�z�;؅�;�>O;�;wx�: �:�y�:�R�:��:���:�� ;�X�:�W�:z�:��9D����4������`(��O���q�Y����j���Y��	���]�ܻN��@���j)�3?�%�R���b���m��{s�rit��Jr��ro��Xn�Eq���x���p����U������*��u欼����O4���I��а��l���|��c���%�����7ؗ�쌙�I���3z���؞��v��rS�����Wҝ��P��v���"x��.����F������{E���D��J�¼	�Ƽ�`Ǽ��ż�n��P)������E��
~��H���⵶�Mм���ü��ʼ�_м�xӼ��Ӽ�Ѽ
8ͼ��Ǽ�[¼����C����$���q���	��fa��<;¼��ü��ļż��ļ��ļ/ż�pƼ�Wɼ�μ;`Լ��ۼ3�����Ji𼯎�u��S��:q�m���1	Ἲ��62�RG�g&２����v���:��  �  �-=	.=�G/=H1=C�3=��5=��7=\�8=K�8=�Q8=G\7=C,6=(�4=�3=�;3=��2=$�2= �2=K�2=^\2=H�1=��/=��-=��*='=��#=� =�V=�L=�=��=� !=�O#=�;%=�@&=�&=��$=��!=��=g�=P�=�=��=�==L�=X=9�=�9 =|�!=��"=%*#=��"=�!=Z !=� =�s=J=�=�?=x�=��=�W=Ol=`�=)#=�=UH=�=o�=?
=��=��=o`	=5]
=�$=i%=w�	=�@=�2=�2�<���<P �<�u�<�;�<��<���<E��<���<<�<���<Q�<��<@��<��<%��<bG�<��<@?�<��<0b�<�*�<;�<�Ö<纑<ُ�<�	�<]uv<c<liO<T =<1y-<"<�<�<��<$G<�<��<ȡ<�M	<L�;܍�;��;�Vj;�z);+i�:��:zs�:pQ�:��:dg; <	;�;-��:��:w��9n���R����库~��8G���j�����"*��BL�������ػ����Ѫ�P$�2U8�D�J�5eZ�Wge�	�k��lm�4tl�@�j���j�L�m��u�a=���|��
����ě�gt��(ר��l���;��|¨��ɤ��:��	���������X��� y������蚼�E۝��w��q��f���hQ��y�@R�������ڦ�Pܬ��v���ҹ� ���c¼�Qü����f5��D���@ڴ��^�������2���ﴼ�����2��ЍǼ �̼?`ϼ��ϼ �ͼU�ɼ�0żYk���f��E���R�����|����ּ��0���P��=�¼��ü�Kļ�PļYOļ��ļ�	Ƽo�ȼj�̼��Ҽ�ټ���@��e�Yl�	��zh�Y��&��hl߼�4߼˛ἢ`����e����������  �  ;�0=��0=��1=|l3=�65=��6=�+8=��8=�8=�d8=�7=��6=X{5=M�4=w�3=�o3=b,3=j3=��2=�m2=:�1=�A0=�@.=ή+=T�(=�%==7#=�H!=
L =�^ =h!=�#=_�$=Ѓ&=P'=Y'=K�%=s#=
� =�=�{=D�=O�=�=�p=cO=*Q= !=�o"=�##=<#=��"=#+"=�c!=�� =� =��=d�=��=�=��=�d=A�=�=*�=Z6=`%=X=�M=�*=r�=1m=s�=R4=��=�9=��
=R-=fR='$�<���<��<=��<s��<5h�<��<g �<�3�<*l�<��<���<���<Q��<'��<&�<�(�<�A�<R��<�\�< ��<A �<���<��< �<�3�<%M�<J�z<
�i<�X<�wG<�19< J.<qX'<k/$<��#<�^$<y$<r� <'m<�a<�p�;���;˒�;�$�;x#V;/6+;�Y;��;�9
;^;Ђ;�;V{;I�:_��:s
:z�.�
:g���Ϻ���<�qa�q���
��ZĦ�%��Mpջ�;󻟌
�����.���?�VON�q!Y�E�_�f c�K�c���c�He�^yi�=�q��}�^}��\䎼���%���$墼
e��&����̣�~Ҡ�1_��J,��Η�}���w���D��˛����<��������)���O���!���֜�ź��./������G?��s-��a'������{���qx��k���b��H���s�������ӱ�����_�Z��p��&f�������¼��Ƽ�eɼ��ɼ=:ȼmIż����󽼴�����f��S���ic��WI��^K���"��|����¼�Bü[�ü��ü��ļ�ż>>ȼ��˼̼м�zּ��ܼ#�~��Oj� ���C��Le��)߼�1ݼ�/ݼ|k߼��㼭F�4M�̾��H����  �  �N4=�-4=��4=��5=�6=��7=0h8=ǰ8=ێ8=�8=�j7=��6=�5=n(5=k�4=�3=ބ3=B3=��2=�2=0P1==+0=J�.="�,=cl*=*,(=$&=[�$=	�#=�#=N$=ey%=��&=�'=Ie(=z(=��&=^%=��"=�� =j�=WZ=�=�/=S=�G=� =C�!="=��"=��"=��"=q""=�!=H !=�� =�Z =� =��=��=w==�H==�q=�Y=��=a�=�M=�s=�*=N}=J=�G=\=�U=ط=�	=�}=0=�<��<9�<ق�<���<��<}��<yr�<CH�<f��<9_�<d�<K	�<8M�<�&�<�Ǻ<�U�<2�<_��< ��<4��<A��<���<���<�	�<]߅<%"~<ϗo<��`<��R<>F<o<<��4<�i0<�.<X,<R�)<�.%<�.<��<��<]q�;���;��;��;�_;OQD;vK4;�+;��&;�} ; ';,�;F�:w/�:$�:-N���FI��|������<1�N�Y�f����������`����Ի�Hﻔ.�����%���3���@�K�s�R�<W��Z��^\�ؑ_� �d�lIm�'�x��/������U���e������呞�aA��ր��;֜�Ϛ������H���!��6�����������f����V��+훼6T��G���>ל��0���ݝ����n,��(��\ȧ��ݫ��᯼�Q��ޭ��ϗ��K������=���}���|��Zݫ�J���Jǯ��ֳ��y���뼼�s����¼�ü�E¼�r��K&��i⻼k���������#����ú��,��1�������]��y���j¼�Bü!ļ� ż�Ƽ�ȼl�˼�Aϼn�Ӽ�Cؼ]�ܼ4<���>l� ��f�༝\޼�#ܼ<�ڼ&ۼ�)ݼ����\��I�J����  �  k�7=�17=q+7=]7=С7=��7=��7=��7=�7=F+7=��6=7e6=��5=b5=9�4=zG4=J�3=%�2=��1=�"1=(H0=wU/=�:.=��,=��+=W*=��(=��'=	'=c�&=�'={�'=c{(=m)='A)=��(=��'=��&=&�$=�#=Ψ!=5� = =T =�O = � =�:!=͟!=B�!=7�!=��!=��!=u�!=�|!=�P!=!=� =�O =C�=m<=Ţ=��=�A=�[=;=��=�K=R�=x=�=�X=tt=��=6=�n=�6=$Z=7�	=�o=��=b)�<@8�<^��<���<G��<���<�p�<ۓ�<���<0��<֕�<���<���<��<�R�<ּ�<��<'Ұ<�x�<`�<H�<���<�'�<�Ï<�k�<���<`�~<�Rs<Z�g<Я\<�_R<\I<t�A<�P<<2�7<��3<��.<B�(<��<��<B<��;X��;�H�;�b�;��;�}r;EZ;� F;�$4;[�!;�^;� �:1��:��a:��9:e/�/�=��"����*�B�V��́�U:��&L���$Ļ�-ڻ/���Y�Z�������(�E�3�(�=��qE���K�ѫP��YU�F�Z�jFa�s�i�|st�7��r��y`�������q��H���w��\��י��u����O昼���(��$k�����G㙼�)��,���� ������nǜ��ŝ��Ξ�M埼a��R���p��9������K�������H������ů�ȭ����Q}��e���?���L��9���ۗ��`���e��?$��4���ؼ�`輼^r��F»�������M���W��m����?����z���ׇ������=����'¼	�ühJż�Ƽ��ȼ�zʼ��̼�#ϼ��Ѽ��Լ��׼�Lڼsܼ��ܼ��ܼx�ۼ��ڼ�zټeټ��ټWXۼ�0޼%��>{�&��g���  �  �C:=Ӊ9=w�8=}E8=�7=�7=�v6=m�5=��5=�|5=�5=��5=T�5=�s5=��4=�.4=�3=��1=o�0=c/=[a.=đ-=��,=eP,=�+=�/+=[�*=� *=��)=�|)=�s)=��)=��)=��)=��)="K)=�(=O�'=Zc&=�<%=94$=�\#=ͷ"=�6"=��!=&]!=�� =� =S@ =�	 =  =/ =N =x� =T!=�!=�� =� =�2=&=.=)#=�U=P�=�=�p=g�=��=N=�=C�=�=��=��=5Z=�=��=��	=%�=%�=�% =	f�<���<4��<	`�<�O�<s��<���<X{�<�!�<���<���<R8�<z��<�U�<���<��<X��<H��<�x�<u��<�o�<N�<C�<���<3>�<�{<�us<Rpk<��c<k�[<�1T<��L<�:F<V�?<Vh9<�w2<��*<(!<�O<r9
<���;T�;�y�;yȱ;^�;�;��s;�R;�3;�;���:�ԫ:��c:�d�9 Nq8�z���[N��ĩ�����z�(���Z�.������ި����ѻ���@��M5��$�%���� ���)��I2��l:���A��I�k P��=W��+_�g
h�|�q��|�5����V���鏼Bǒ�0��^����������������Ԝ�V���c㛼�'��᜚�a�������B��V���蟼�ء�ጣ��䤼�㥼_���-_��V���ʨ�6���L$��a���`����R��\Щ��P��1���k��fi����u/������#ղ�޴����cܷ�M���$�����0���<��
,���ؾ��&�����ܾ������Ⱦ�iu�������¼�-ż_�Ǽ7ʼb̼�*μ ϼQ�м� Ҽ�WӼ:�Լ)�ռ��ּ�}׼\�׼��׼k�׼��׼��׼��ؼ�Qڼ�rܼ��޼I��\�C8��  �   <=|�:=ۦ9=�28=$�6=DH5=�4=�F3=�2=�3=1�3=v=4=��4=��4=h�4=ȟ3=�&2=�^0=+�.=�,=i�+=��*=c�*=�*=��*=�N+=�+=K�+=F�+=@\+=�+=e�*=w*=� *=D�)=�@)=��(=:(=A`'=r�&=��%=C%=�m$=�o#=�E"=�� =&�=S�=˼=�O=�b=��=$�=ܩ=�] =�� =�T =�n=�=�v=q�=;�=H�=�=g�=9=j3=)B=v=��=M�=g�=�1=��=-�=ݮ=]=��	=)=�=�=j/�<15�<�=�<3�<| �<���<:U�<4�<̀�<�w�<�J�<�<�s�<D/�<2��<抴<4E�<A��<�
�<��<��<E��<h+�<TӁ<�G{<��t<�o<�k<��f< ua<�~[<��T<2M<4E<��<<��3<��*<%� <�<7<�, <�f�;&��;�ſ;���;37�;��};�!P;wf";ǚ�:�X�:��):
�\9���ѹ{-��Y~��ߵ������9/�o�f��ɑ��R���̻E��j���]�Z��|��o������#�/y*�ڐ2�s!;���C���L���U���^�X�g�Fq��y�$�����Ϋ�����DG�������㕼:���\��������)�����w���U���}��&��c��盼,���q.���=���@������	Z�����J̪�	���������3���̦�zæ�
����S��ͺ���/������{���k��/���ڬ�K<��ҩ���&���ɲ�s�������)���/s��06�����jiü�Lļ�4ļKü���i���e���XB��]���_ļ��Ǽ�u˼��μ=�ѼΔӼ�xԼ�Լu;Լ��ӼJ4Ӽ$Ӽ1Ӽ��Ӽ�`Լ�%ռ��ռ;�ּ)�׼T�ؼ=4ڼ��ۼOݼ��޼"��n��  �  �<=?l;="y9=�;7=m�4=J�2=�1=D�/=��/=,10= 81=du2=]�3=�4=`�3=B�2=8�0=�u.=�	,=��)=zf(=ߪ'=�'=VZ(=�`)=߅*=��+=y=,=�,=Ie,=��+=[X+=K�*=�)=�])=f�(=�l(=@(=��'=�r'=��&=�G&=i4%=̵#=E�!=�=�=\�=v�=�=�>=!0=��==�@=��=C�=![=̆=�V=�+=�b=�?=��=� =�=��=ը=�0=\4=�=�x=;�=��=��=nH=��=5>	=m�=�=zs=��<���< ��<�)�<���<� �<]�<}e�<Ɂ�<Qο<��<�Ӹ<	<�<+,�<�<���<#®<��<Hˡ<4[�<6��<r/�<k �<b�v<!fo<�j<M�h<D5g<�e<�Ic<J_<��X<5Q<��G<\�=<a�3<)<j�<�Y</n
<}� <ډ�;�M�;K�;tΰ;��;�\y;�4?;�;�O�:�0�9��'�WF�KY���}�0d��fF����κ�a
��<���y�,�����»�M������	��y����Rw�>���M��e ��V&�T.��H7��]A��K��'V��`��ci�u�q�y�7?���u��䙆��뉼'���E쑼����ज़�e��r��8S������pN��!w���������9���	��T�������=���t��ך���Pﰼ�[��1Y��SI��V��� ��V˦��U��H���1�������[֦����9���H��.��t꫼����9-��?󭼱���ڰ��m��W߶�$��{����ü�iǼg�ɼ��ʼ�BʼviȼL�żü���������~üO�Ƽ�3˼rмk�Լ�ؼx)ڼ��ڼ��ټ��׼D�ռ�ӼM3ҼF|Ѽ�Ѽ?vҼ��Ӽ�Nռx�ּ�_ؼf�ټM�ڼ�ۼi�ܼ9�ݼ��޼�Z��  �  �==�(;=�8= �5=��2=�/=��-=j�,=g,=8-=�.=�0=�2=��2=I�2=�1=�A/=]i,=;q)=�&=�
%=PC$=M�$=�%=�J'=�$)=Y�*=c,=j�,=��,=�=,=&k+=�w*=��)=��(=�8(=��'=,�'=�'=��'=eS'=ޑ&=�;%=�D#=�� =��=�9=S�=�>=*�=�=�]=�I=+P=��=��=�u=�=��=)=qc=�-=��=.v=	=�J=�=,q=ݚ=]=$�=Q�=.�=*�=�A=�=�=C}=m=Բ=�X=B��<�T�<�	�<��<�O�<-�<?��<���<{
�<N۸<���<X�<ر<4�<(��<(9�<�Ƭ<�<f#�<IǕ<<�<��<�>u<ͤi<N�b<��_<�_<��`<�Ob<�)b<��_<�;Z<�QR<zsH<;k=<R�1<��&<�<g�<�<=��;���;���;&��;!�;|*�;�sj;8r%;ҷ�:z��9r����؂�n����(˺��̺	ɺ�Ϻ�J�T��<�L���������Cֻd���5�R��@���(�$Z�Ź����i� �>%��v,���5���@�!WL���W�wGb�R�k�!�s���z�A��*����ۅ�<D��.���˼��Ø��$�� B���i�����t��T�������=��'��5ՠ��$��Ϛ��@��s����꫼p"���P��Ｗ�����s��hU��Xa��dP���ͧ��\���5���G��/L��\ܦ�H����8������c��hԬ���������m���g���e��~���r%��0����ü/ɼ��ͼ��мڙѼ(zм�ͼ�ʼ,�ƼuXļv�ü��ż�ɼ�μf�Լ�uڼ��޼����3�D�߼(�ܼ ټ��ռ��Ҽ&FѼ��мW�Ѽ�wӼ��ռ;�׼�zټ��ڼ ܼ
�ܼݼJlݼ�.޼o�߼�  �  ��<=ۊ:=��7=�4=�0=�N-=��*=w�)=م)=@�*=֔,=��.=�0=2�1=l�1=�_0=��-=�*=�.'=�0$=U"=�B!=o�!=F#=�<%=�'=�)=�+=,=�,=(,=9+=�*=n)=h#(=��'=�R'=�V'=�x'=|�'=�B'=�m&=��$=Ɂ"=y�=�)=��=� =�F=ڝ=�9=��=tF=��=�=��=�l=��=G=M=d�=	f=D�=�t=�:=��=�=�=��=�=��=��=��=qg=μ=��=�C
=��=�f=4=�=�_�<��<q�<&��<M�<-�<ث�<���<;�<���<R��<p�<?+�<�%�<�Ǯ<�<̪<m��<ʣ�<䎒<�̇<�.{<uj<_�]<8!W<�9U<��V<�eZ<u�]<8�_<Zi^<6�Y<CR<��G<�<<��/<�#<��<��<�<<�t�;���;��;d�;�P�;-��;�X;Q�
;�q:F8�6R���<�i�����	�����il��Ѽ��x'���\�Fq��XH���Z�g�@G� "�7�'���(��<'�'u$��f"�\�"�B�%�٘,�F6�uA���M��Y��d��1n� �u�B?|�����-����|���5��E4��>=��?���䩼 ݯ�T᳼�f��YM�������@���L��3K���7��e�������	���W֯�Tﵼ�׺������	��� ��f���!�������m��s.������j��.���R[��1p���\���Ӭ������魼F�������ݜ������B̰�ٝ������
����}ǼFμ�_Ӽ��ּ�|׼��ռBUҼh�ͼ��ɼD�Ƽ��ż'�Ǽn)̼�FҼq ټx�߼�f������d��Cἱjܼ-�׼@+Լ��Ѽ`4ѼZ�Ѽ=�Ӽ�ּG�ؼk�ڼ�Jܼ�;ݼ
�ݼ��ݼ�ݼ�S޼��߼�  �  J{<=��9=�6=t�2=��.=9t+=��(=J�'=Ï'=��(=�+=M�-=��/=s1=�1=x�/=$�,=�Z)=j�%=�c"=� =Y1=��=�L!=)�#=h}&=~)=�+=1,=�u,=��+=��*=�)=y�(=Ԧ'=n'=k�&=�&=�4'=U'=�'=/&=�s$=��!=`�=V�=7=�3=8=��=	S=B=6�=y�=��=�=ê=� =$5=��=�V=ɂ=:�=�`=dC=�"=]�=� =��=Q$=j?=Q=V�=�=fR=2u=�	=�,=��=��=4� =w��<�y�< ��<qx�<���<'��<_��<�&�<+1�<���<�<�R�<��<ɔ�<���<�N�<NV�<�t�<�ݚ<�S�<� �<Hwt<�~b<��U<DO<��M<��P<�iU<GZ<�@]<��\<��X<�KQ<J�F<��:<�=.<��!<5�<!�<y<���;��;f��;0Y�;�E�;�;��I;�
�:�:�%��cϺ����(�M9*�^��2���
���8o2���h�!ř�2�Ż��Q�U���*��s/�U�/�#-���(��u%���$�'��J-���6�IB���N�:[���f��p�"�w�)�}��:�������@������{���a}��>/���d��W7����������y��q���F�������z��������F*���^���ѫ�G���e0��t���.���}(¼�俼%���3浼����Ъ�d
��!��Ǥ�p奼jާ�I%���@���ҭ����YĮ��i���������[﮼�_�� ���k����¼�iʼߛѼW׼��ڼ��ۼ��ټ{vռ�dмȘ˼�Lȼ#kǼ[_ɼ�ͼ�Լ��ۼ6��I輷�&����C�k�޼�ټ�\ռ4�Ҽi�ѼPҼE-Լ��ּMRټl�ۼ�KݼY/޼�g޼B޼�,޼L�޼�Q��  �   V<=��9=ZU6=+b2=].=��*=�!(=��&=��&=�F(=$�*=7-=;y/=��0=W�0=�C/=��,=-�(=�%=_�!=%j=\t=��=z� =�0#=B&=k�(=��*=R,='^,=��+=)�*=�)=�q(=�w'=C�&=��&=��&=D'=+?'=U�&=&=�H$=��!=f%=�R=K�=]�=/|=)�=��=�=k=�?=��=�=c=Ѱ=r�=1M=��=��=�=Т=e�=+�=�=$�=��=��=�=	7=i=D�={*=E=�}	=a�=l�=}�=� =��<
F�<{�<��<H�<��<��<�ܼ<�³<�</�<��<��<���<�	�<L��<�˨<Q�<�8�<x��<"�<�r<l�_<d�R<�5L<�!K<�:N<��S<.�X<MK\<�U\<yX<��P<�F<�`:<��-<�1!<@�<G+<M�<���;���;]-�;���;m�;��;]D;���:;T�9N�O��m��C��3���3�ï'������Q��`�6�C:m��m����Ȼ63������!���,��G2��v2�6/��*���&��P%���'���-�&
7�;�B��SO���[�"Dg���p�.gx��.~��o��)���i���%��tN�������ꝼ`���l�����Gp��b�Mo���q��'���tA��鬥��K��ϸ���������|u���V���쿼�2üܡüK��7¼��궼�Ȱ��Y���d���E���򤼃�����k��ޖ���2�����6��ث��a.��F#�������_������üx{˼��Ҽ��ؼ�Eܼ[�ܼ��ڼv�ּ�KѼR̼z�ȼ��ǼB�ɼ�μTeռZݼ.�֩�d�������Ho��߼Y_ڼ��ռO�ҼC�Ѽ1zҼ�ZԼ�ּ�ټ��ۼ��ݼ��޼��޼I~޼<[޼*�޼����  �  J{<=��9=�6=t�2=��.=9t+=��(=J�'=Ï'=��(=�+=M�-=��/=s1=�1=x�/=$�,=�Z)=j�%=�c"=� =Y1=��=�L!=)�#=h}&=~)=�+=1,=�u,=��+=��*=�)=y�(=Ԧ'=n'=k�&=�&=�4'=U'=�'=/&=�s$=��!=`�=V�=7=�3=8=��=S=B=4�=w�=��=�=��=� =5=��=�V=��=(�=�`=LC=�"=C�=� =��=J$=z?=�Q=ʃ=�=�S=�v=�	=�/=�=�=� =0��<̅�<���<���<���<���<���<�4�<�>�<M��<���<]�<�
�<���<�Ƭ<kQ�<�V�<�r�<�ٚ<�M�<��<Mdt<�hb<��U<�O<9�M<vP<#MU<+Z<#&]<��\<��X<�7Q<��F<��:<�4.<�!<ظ<�<��<S��;O��;��;���;Dx�;(�;PJ;���:��:��#��κ�:�p�'���)��Y��j�*m
�w��p2���h��י�u�Ż�)�f�Z�l4*�|�/�?0��)-��)�B�%��$�)'��d-���6�h^B�@�N�J[���f��)p��w�(�}�I=������;B����>����}���/��Ee���7������<��� z������F�������z��#������J*���^���ѫ�H���f0��u���/���~(¼�俼%���3浼����Ъ�d
��"��Ǥ�p奼jާ�I%���@���ҭ����YĮ��i���������[﮼�_�� ���k����¼�iʼߛѼW׼��ڼ��ۼ��ټ{vռ�dмȘ˼�Lȼ#kǼ[_ɼ�ͼ�Լ��ۼ6��I輷�&����C�k�޼�ټ�\ռ4�Ҽi�ѼPҼE-Լ��ּMRټl�ۼ�KݼY/޼�g޼B޼�,޼L�޼�Q��  �  ��<=ۊ:=��7=�4=�0=�N-=��*=w�)=م)=@�*=֔,=��.=�0=2�1=l�1=�_0=��-=�*=�.'=�0$=U"=�B!=o�!=F#=�<%=�'=�)=�+=,=�,=(,=9+=�*=n)=h#(=��'=�R'=�V'=�x'=|�'=�B'=�m&=��$=Ɂ"=y�=�)=��=� =�F=؝=�9=��=pF=��=�=��=�l=��=G=9=K�=�e="�=et=T:=��=��=a=��=�=��=�=��=�h=�=�=�G
=a�=>m=�;=�=�t�<��<҉�<V��<Oh�<�:�<���<���<8U�</ֲ<�Ǯ<;�<�;�<�2�<eѮ<|��<<ͪ<E�<p��<���<���<�	{<�i<#�]<6�V<�U<��V<�.Z<R�]<Qg_<�8^<&�Y<��Q<��G<� <<��/<��#<��<�<�L<���;/��;��;���;��;��;��X;�n;ku:�s*�J������\�}��g ���������>��p{'��]������|��|�绑���u�TK"�b�'��$)�
x'�Ű$�E�"�:�"�K%&�:�,�TD6�F�A�+�M�
�Y��d�{Gn�nv��L|�)����1�����~��7��`5��>��߻���䩼{ݯ��᳼ g���M�������@���L��@K���7��l����������[֯�Wﵼ�׺������	��� ��g���!�������m��s.������j��.���R[��1p���\���Ӭ������魼F�������ݜ������B̰�ٝ������
����}ǼFμ�_Ӽ��ּ�|׼��ռBUҼh�ͼ��ɼD�Ƽ��ż'�Ǽn)̼�FҼq ټx�߼�f������d��Cἱjܼ-�׼@+Լ��Ѽ`4ѼZ�Ѽ=�Ӽ�ּG�ؼk�ڼ�Jܼ�;ݼ
�ݼ��ݼ�ݼ�S޼��߼�  �  �==�(;=�8= �5=��2=�/=��-=j�,=g,=8-=�.=�0=�2=��2=I�2=�1=�A/=]i,=;q)=�&=�
%=PC$=M�$=�%=�J'=�$)=Y�*=c,=j�,=��,=�=,=&k+=�w*=��)=��(=�8(=��'=+�'=�'=��'=dS'=ޑ&=�;%=�D#=�� =��=�9=R�=�>='�=�=�]=�I=$P=��=��=�u=�=��==Oc=�-=��=�u=�=�J=��=�p=��=S=_�=��=z�=R�=1E=k�=�=�=�=�=�e=���<9u�<�,�<��<{v�<RT�<���<7	�<�/�<��<iδ<N��<��<���<x��<�@�<Ȭ<� �<�<X��<ϋ</l�<�u<�ai<Ub<�Y_<J_<��`<	b<�a<Q_<{�Y<YR<�EH<�G=<��1<߂&<�<H�<-�<���;C�;iK�;0F�;ަ�;վ�;��k;P�&;F7�:(� :�0��=���	����rɺ�}˺.Ⱥ)Ϻ~��@����L��E�����9�ֻ�����O����Y��uz�+��7����!���%��,��-6�YA�e�L��W��lb���k���s�ίz�sH������߅�0G��X���c���IĘ��%���B��Ij��~���ht����������=��$'��Hՠ��$��ښ��@��y����꫼t"���P��񼷼����s��iU��Ya��eP���ͧ��\���5���G��/L��]ܦ�H����8������c��hԬ���������m���g���e��~���r%��0����ü/ɼ��ͼ��мڙѼ(zм�ͼ�ʼ,�ƼuXļv�ü��ż�ɼ�μf�Լ�uڼ��޼����3�D�߼(�ܼ ټ��ռ��Ҽ&FѼ��мW�Ѽ�wӼ��ռ;�׼�zټ��ڼ ܼ
�ܼݼJlݼ�.޼o�߼�  �  �<=?l;="y9=�;7=m�4=J�2=�1=D�/=��/=,10= 81=du2=]�3=�4=`�3=B�2=8�0=�u.=�	,=��)=zf(=ߪ'=�'=VZ(=�`)=߅*=��+=y=,=�,=Ie,=��+=[X+=K�*=�)=�])=f�(=�l(=?(=��'=�r'=��&=�G&=h4%=̵#=D�!=�=�=Z�=t�=�=�>=0=��=v=�@=��=0�=
[=��=�V=�+=�b=N?=}�=� =,�=k�=��=�0=X4=j�=�y=��=��=��=N=�=�G	=�=�=\�=��<8�<�<]W�<��<91�<�<�<ٔ�<@��<���<߹�<��<�X�<�B�<7�<ǡ�<Į<d�<���<�G�<hr�<��<�ۀ<��v<�o<�j<�+h<U�f<�ke<��b<��^<:�X<S�P<ӮG<�=<~n3<U�(<1�<+g<��
<�� <k��;���;`��;hw�;弘;��z;b�@;5*;`O�:���9^�dv�*U�dz�f���a���eκOf
��B<�*lz�Z���E@ûq�㻞$��
�	�>��).�d�������� ���&��o.���7�i�A��L��]V�GG`��i���q�n�y�KH���|��󞆼Dߨ��F(��������e���r���S��쨨��N��Ww��?������49���	��b�������=���t��ܚ���Sﰼ�[��3Y��TI��W���!��W˦��U��H���1�������[֦����9���H��.��t꫼����9-��?󭼱���ڰ��m��W߶�$��{����ü�iǼg�ɼ��ʼ�BʼviȼL�żü���������~üO�Ƽ�3˼rмk�Լ�ؼx)ڼ��ڼ��ټ��׼D�ռ�ӼM3ҼF|Ѽ�Ѽ?vҼ��Ӽ�Nռx�ּ�_ؼf�ټM�ڼ�ۼi�ܼ9�ݼ��޼�Z��  �   <=|�:=ۦ9=�28=$�6=DH5=�4=�F3=�2=�3=1�3=v=4=��4=��4=h�4=ȟ3=�&2=�^0=+�.=�,=i�+=��*=c�*=�*=��*=�N+=�+=K�+=F�+=@\+=�+=e�*=w*=� *=C�)=�@)=��(=:(=@`'=r�&=��%=C%=�m$=�o#=�E"=�� =$�=Q�=ȼ=�O=�b=��=�=ҩ=�] =y� =�T =|n=�=�v=B�=�=�=<=�=�=3=�A=A=��=��=o�=n3=˗=��=�=Ye=	�	==�(=�+=W�<a�<�m�<�e�<S5�<p��<!��<[i�<���<V��<�u�<+�<ۓ�<�H�<*ɷ<��<]G�<P��<��<z��<+ה<��<��<���<9�z< lt<Y?o<ӳj<y(f<-a<� [<BYT<l�L<��D<z�<<y�3<	x*<Ƒ <w%<	V<D[ <���;Pv�;~o�;]t�;��;��;��Q;K$;���: ��:7�/:�r9,{�K ʹ�$*��^|��d��B�����/�/�g��-�� ԰�A�ͻ:��}0��Y��x`��
�-l����#���*�u�2��z;�p>D�M�V��_�I#h�(q���y�R.������������dJ��􍒼N啼R;���]�����"������������U���}��@��.c��盼7���z.���=���@������Z�����L̪� 	���������3���̦�zæ�����S��ͺ���/������{���k��/���ڬ�K<��ҩ���&���ɲ�s�������)���/s��06�����jiü�Lļ�4ļKü���i���e���XB��]���_ļ��Ǽ�u˼��μ=�ѼΔӼ�xԼ�Լu;Լ��ӼJ4Ӽ$Ӽ1Ӽ��Ӽ�`Լ�%ռ��ռ;�ּ)�׼T�ؼ=4ڼ��ۼOݼ��޼"��n��  �  �C:=Ӊ9=w�8=}E8=�7=�7=�v6=m�5=��5=�|5=�5=��5=T�5=�s5=��4=�.4=�3=��1=o�0=c/=[a.=đ-=��,=eP,=�+=�/+=[�*=� *=��)=�|)=�s)=��)=��)=��)=��)="K)=�(=O�'=Zc&=�<%=94$=�\#=̷"=�6"=��!=$]!=�� =� =P@ =�	 =� =/ =F =m� =F!=�!=m� =� =�2=X&=�=�"=ZU=�=a=dp=�=3�==�=��=,�=��=�=�^=��=*�=�	
=z=�=�7 =���<�
�<��<���<���<H��<d'�<��<V�<��<��<�_�<���<p�<FϹ<���<���<(��<4j�<:�<7R�<���<��<�͆<$�<�S{<?s<Jk<�$c<�a[<R�S<k�L<`�E<ȓ?<#69<
U2<hp*<�&!<m_<�Y
<�:�;��;b�;�x�;�!�;迋;�\u;&�T;��4;JX;k�:D�:�Qi:=�9�i�8�e��QL��E�������=)��B[��燻�,���I���zһ$��;���\��כ�v�O!�v*�w�2���:�]TB�w`I�.IP�t|W��`_��5h���q��9|��?��,�� \��2�ʒ����/���]����𙼻���������S՜������㛼(������v�������B��_���
蟼�ء�匣��䤼�㥼`���._��W���ʨ�6���L$��a���`����R��\Щ��P��1���k��fi����u/������#ղ�޴����cܷ�M���$�����0���<��
,���ؾ��&�����ܾ������Ⱦ�iu�������¼�-ż_�Ǽ7ʼb̼�*μ ϼQ�м� Ҽ�WӼ:�Լ)�ռ��ּ�}׼\�׼��׼k�׼��׼��׼��ؼ�Qڼ�rܼ��޼I��\�C8��  �  k�7=�17=q+7=]7=С7=��7=��7=��7=�7=F+7=��6=7e6=��5=b5=9�4=zG4=J�3=%�2=��1=�"1=(H0=wU/=�:.=��,=��+=W*=��(=��'=	'=c�&=�'={�'=c{(=m)='A)=��(=��'=��&=&�$=�#=Ψ!=4� = =T =~O =�� =�:!=˟!=>�!=3�!=��!=�!=m�!=�|!=�P!=!=ӽ =�O =$�=G<=��=��=�A=�[=�:=H�=UK=�=N=-�=6Y=�u=��=<9=;s=G==sb=��	=�|=��=�L�<s`�<�"�<���<5��<���<���<���<��<��<8��<��<��<���<�k�<�κ<��<K԰<�r�<�ޥ<�2�<#��<��<��<>�<_΄<�h~<(�r<"fg<zF\<��Q<��H<˩A<�<<��7<�3<M�.<��(<��<��<Aa<$?�;5�;7ܶ;��;�͉;�t;��[;L�G;�5;A#;�;��:]�:�f:���9��#�ͼ;�V�������N*�)W�41�����`箻U�Ļv�ڻY�����m��c�:P)��V4�?�=�i�E��K���P�=�U���Z��ya��j���t��D���|��oh������Vv�����Mz��(���Aٙ��v������昼���O)��ck��5���j㙼�)��@���� ��᛼vǜ��ŝ��Ξ�Q埼d��T���p��;������L�������H������ů�ȭ����Q}��e���?���L��9���ۗ��`���e��?$��4���ؼ�`輼^r��F»�������M���W��m����?����z���ׇ������=����'¼	�ühJż�Ƽ��ȼ�zʼ��̼�#ϼ��Ѽ��Լ��׼�Lڼsܼ��ܼ��ܼx�ۼ��ڼ�zټeټ��ټWXۼ�0޼%��>{�&��g���  �  �N4=�-4=��4=��5=�6=��7=0h8=ǰ8=ێ8=�8=�j7=��6=�5=n(5=k�4=�3=ބ3=B3=��2=�2=0P1==+0=J�.="�,=cl*=*,(=$&=[�$=	�#=�#=N$=ey%=��&=�'=Ie(=z(=��&=^%=��"=�� =j�=VZ=�=�/=R=�G=� =A�!=��"=��"=��"=�"=i""=�!== !=� =nZ =k =e�=׷=�v=�=PH=�=�q=uY=J�="�=�M=�s=O+=X~=�K=�J=w=R[=O�=7	=.�=�==>�<�3�<)�<���<^��<���<���<���<�w�<���<���<F�<G+�<�i�<N=�<�׺<�^�<�<��<�t�<q�<���<B��<
t�<#�<J��<I�}<O8o<�x`<�dR<��E<��;<ʎ4<a&0<k�-<2,,<�)<�%<�-<7�<�</��;x�;w��;�@�;�;a;��E;n�5;�y-;[V(;K�!;e�;��;R��:C�:�:�O�J�G����e���|1��Z��߀�ކ������� ���ջ��В�����%�34�6A�izK�V�R�{�W�ZZ��\�a�_�e�Qom���x��;��(�������ְ�����甞��C��|���uל��Ϛ��	������)"��o�������У��~����V��8훼AT��N���Cל��0���ݝ����p,��*��]ȧ��ݫ��᯼�Q��߭��ϗ��K������=���}���|��Zݫ�J���Jǯ��ֳ��y���뼼�s����¼�ü�E¼�r��K&��i⻼k���������#����ú��,��1�������]��y���j¼�Bü!ļ� ż�Ƽ�ȼl�˼�Aϼn�Ӽ�Cؼ]�ܼ4<���>l� ��f�༝\޼�#ܼ<�ڼ&ۼ�)ݼ����\��I�J����  �  ;�0=��0=��1=|l3=�65=��6=�+8=��8=�8=�d8=�7=��6=X{5=M�4=w�3=�o3=b,3=j3=��2=�m2=:�1=�A0=�@.=ή+=T�(=�%==7#=�H!=
L =�^ =h!=�#=_�$=Ѓ&=P'=Y'=K�%=s#=
� =�=�{=C�=O�=�=�p=bO=(Q=�!=�o"=�##=<#=��"=+"=�c!=w� =� =x�=R�=ަ=�=��=�d=�=�=��=6=#%=&=�M=+=��=n=�=�6=��=S>=��
=5=�[=�:�<���<o��<���<��<w��<��<�G�<[�<���<�8�<L��<~��<��<{��<�*�<�5�<I�<ᝮ<>X�<|�<��<���<0��<?�<M�<9)�<�{z<4@i<r�W<�*G<��8<�.<�'<X�#<}�#<�:$<��#<E� <l<m<؞�;c �;�;J��;bW;TK,;��;5
;y;�Z;��;/H;$�;o<�:>�:b�:�8&��e��xϺ�+:<���a�ǹ�� i���5��T���� ֻm��P�
���kI/�C=@�R�N�pnY�9`�%bc�Md��,d��te���i�>�q���}�E���쎼���� ��袼�g������Σ��Ӡ��_���,��yΗ�ϑ��Jw���D���3��P��������)���O���!���֜�ɺ��1/������I?��t-��b'������{���qx��k���b��H���s�������ӱ�����_�Z��p��&f�������¼��Ƽ�eɼ��ɼ=:ȼmIż����󽼴�����f��S���ic��WI��^K���"��|����¼�Bü[�ü��ü��ļ�ż>>ȼ��˼̼м�zּ��ܼ#�~��Oj� ���C��Le��)߼�1ݼ�/ݼ|k߼��㼭F�4M�̾��H����  �  �-=	.=�G/=H1=C�3=��5=��7=\�8=K�8=�Q8=G\7=C,6=(�4=�3=�;3=��2=$�2= �2=K�2=^\2=H�1=��/=��-=��*='=��#=� =�V=�L=�=��=� !=�O#=�;%=�@&=�&=��$=��!=��=g�=O�=�=��=�==L�=X=8�=�9 =z�!=��"="*#=��"=��!=U !=� =ys=?=�=�?=d�=��=�W=.l=;�= #=��=+H=]�=`�= ?
=��=>�=~a	=�^
=Q'=�(=��	=oF=�9=�B�<P�<<�<���<�T�<E��<���<��<���<i9�<���<�%�<V��<���<m��<!��<�P�<��<Y@�<��<[�<��<}�<۱�<॑<dx�<���<�?v<)�b<&2O<��<<�D-<%�!<�g<m<�<�-<ŀ<��<�<�U	<�l�;���;��;��j;�+*;���:Qa�:�,�:n�:���:�C; 
;]m;�:D?�:���9.����Є�а�I���]G��j�򅻙l��d����j���]ٻE��|���<$��8�M6K�o�Z�ǝe���k��m��l��j�a�j���m��u�;F�����������ț��w���٨�Tn���<��vè�Eʤ�D;��q�������������By������蚼����O۝�x��q��j���kQ��|�BR�������ڦ�Qܬ��v���ҹ� ���c¼�Qü����f5��D���@ڴ��^�������2���ﴼ�����2��ЍǼ �̼?`ϼ��ϼ �ͼU�ɼ�0żYk���f��E���R�����|����ּ��0���P��=�¼��ü�Kļ�PļYOļ��ļ�	Ƽo�ȼj�̼��Ҽ�ټ���@��e�Yl�	��zh�Y��&��hl߼�4߼˛ἢ`����e����������  �  u�+=H,= q-=~�/=2h2=��4=�7=[@8=�8=�$8=%7=��5=�4=�{3=
�2=�^2=�S2=�o2=�z2=a/2=�G1=[�/=��,=��)=��%=Q�!=&�=�K=�>=O�=0=2�=)-"=mS$=�z%=xL%=��#=P� =�|=��=�=� =�q=�D=h9=�=��=3{=�!=�"=%�"=4�"=p�!=}� =��=��=�=�=�=�B=&q=+=S+=E=�q=��=��=e=��
=t9=!�=|�=��=C	=�)
=`_
=MA	=E�=�h=�/�<�i�<R��<���<XX�<���<I�<��<�V�<�X�<���<�f�<�Z�<���<�D�<�<���<�%�<�7�<v��<�y�<�n�<)��<E�<�,�<{Ɗ<�Ԃ<o�r<�^<�
I<Tx5<71%<�<7s<�J<ҭ<�X<͵<�h<��<�V<!5�;��;Ԧ�;=�O;hg;)C�:���:�]�:�;�:���:#��:.N;+#�:#�:��:�9�e���񒺱y��Fb(��O�r�浈����@��������ܻW����F�)�2?���R���b���m��s���t��`r���o�Oin�!q���x�/�������X��M���2,���笼�����4��xJ��1���Jl���|������D���-��Hؗ�����S���;z���؞��v��vS�����Xҝ��P��w���#x��/����F������{E���D��J�¼	�Ƽ�`Ǽ��ż�n��P)������E��
~��H���⵶�Mм���ü��ʼ�_м�xӼ��Ӽ�Ѽ
8ͼ��Ǽ�[¼����C����$���q���	��fa��<;¼��ü��ļż��ļ��ļ/ż�pƼ�Wɼ�μ;`Լ��ۼ4�����Ji𼯎�u��S��:q�m���1	Ἲ��62�RG�g&２����v���:��  �  A]= "=(=��=�E=d�=3$=(=�G*=�++=�+=;W*=re)=�(=9�'=�\'=7'=��&=C&= %=�"=��=��=�=�=�=�=;��<��<z*�<se =d=�&
=�]=��=��=[x=^�	=54=�x�<Qq�<�-�<���<�P�<��<<E =s=��=�H=�=�=��=�u=]�=VM=H�=�=�s=A�=��=�=��=�?=_O=�=�� =��<�?�<���<��<��<e��<���<�	�<���<~��<�<�<�<�>�<�G�<�J�<}��<븝<8'�<"͏<��<
2�<�N�<��<p�<�ݯ<��<A�<fӭ<ۨ<��<8ڜ< �<a�<>C�<!X�<�,�<�,x<̧h<t�T<U|;<|<�%�;��;�;�;��);|��:���:���:��;��U;�S�;��;��;@_I;��:�Ny���� ��_����SϻQֻ� ʻ��������0�^���(�V���-�����M['��oQ�<~��裘�#���&�Ļ��ػ�u�S� ��"�:1�N35��GP��jo�]L��煘��˦�阱�ٷ�B��K{����������������)X��鵱�e����̼�ۼ�R��x４l�K�|?�Jg߼~@Լmjɼ2��7m���Z��3�������&����ȵ�L����1���3�������;ŷ�L��<����Ƽ[Ѽ��ݼӟ�ؿ���, �c���U�6C�F���^�g�:�޼�Yۼ��ܼI�����SY�����N	�B	�������^R��7����Q�ܼ8(׼qԼ��Ӽ&ռ�ּS�ؼ�ڼuۼ&�ۼ�ܼ��ܼ�޼��⼕_�k��`b�����ω�I��� ��C����t�@1��:���������������
��N���� ��& ��  �  �=+^=�F=��=�=!A =��$=�C(=�[*=;2+=7+=�a*=�w)=��(=o�'=t'=�)'=��&=:G&=�%=��"=�-=DI=^V=��=�=m/=d�<�l�<���<\y==��
=��=�Z=~i=I=I�
=�
=r|�<��<��<`L�<���<`/�<�%=��=s=��=Q�=��=+�=`{=I�=�a=��=��=�=��=s�=8=7�=�_=��=Gq=Y=\��<�Q�<��<�z�<t5�<�C�<���<M��<7!�<��<�#�<AD�<�d�<���<d��<���<��<ژ�<�:�<���<c"�<�؝<�8�<���<�C�<O�<M �<�ҭ<��<[�<��<] �<���<rr�<�y�<�C�<'bx<li<�_U<i�<<75 <<<��;�K�;��=;�;Q��:��;2v/;Ĝb;ړ�;|j�;�9�;oR;�i�:iac�F.���x��*���vŻ �̻Vv��;���]��j�V���#�\�!��۬�J'���P�z��뿗�����Ļlػ����� ����ա��.4�_�N��l������x���k��Y���>���ȶ��D���%��p���K��j���d8��؀��L�����ʼ�ټ&��;�� �����;�ݼs�Ҽ�~ȼR���s#��~=��0������y������䄶���������ڶ��඼�����2������_sƼ�{м�]ܼ���#���b���V����� �kr�����_ ��ݼZAڼ��ۼ�἟��&M���I����
�j �K��W���������H ��(ܼO�ּ�]Լ�Ӽ[�Լz�ּ�aؼF�ټ��ڼ��ۼtܼ��ܼ.�޼ɽ⼩	�A�Ib��������o����H��Y��XT��8��m���t(��k���
�������5�����  �  �5=�=�d=BZ=n�=�!=	�%=W�(=Uv*=�*+=�+=o*=��)=��(=)(=��'= L'=[�&=j=&=�%=<�"=�=�8=��=��=�C
=	e=b=%� =�=�=��=�=W�=��={�=V�=��=�i=2=nF�<'��<,k�<4u�<�<��=�=�==Z9==��=I~=�x=7=��=?=L�=l�=��=��=�=�=i�=�(=�=�=FM�<��<G��<�z�<*�<���<�S�<_b�<��<���<� �<�(�<���<���<	��<�|�<t��<���<|�<��<���<
�<�;�<Ԟ�<51�<�Y�<=�<̭�<��<R�<�u�<|��<� �<�܌<.��<�V�<��x<�i<9W<9@<R�%<�<ހ�;�@�;�-u;��?;��,;��8;In[;od�;{V�;���;}��;�j;��;���9�䲺pH��8������%������������u�ŢA�bl�r��qG���,	��k'�ǁO�f�|��~��^#������nOֻ��� ��{�؟���1�#�J�F�f�>��mߐ�xݝ��䧼���4߯�����੼G��J���$V����#������SƼ�FӼp޼g�弎��R��l(�'�ؼ�WϼfƼ�J��L����$�����\���4V��;?��#���~�� �������'඼ҷ�%��
}��@9ż/Aμ��ؼo?�����L���P��M������h����l�YIڼ@2׼O�ؼ�_޼��`=�����P��{��z��h�i{���P�����]�Iۼ[�ּ^Լ�Լ'�Լ�aּY�׼�Xټ}fڼ-ۼ��ۼ��ܼ��޼��gV�g~�����1��	��^��X��k��O�Z&��z��(
��2�k��8��Ӈ��6��M����J��ox��  �  �l=~�=�=��=d�=L#=!x&=m�(=�9*=��*=i�*=�K*=��)=�)=i(=S�'=~Q'=��&=�%=.�$=̼"=��=�6=@�=��=�=I�	=$$=��=�=�	=�o=R*=�U=�(=	=?=|=(�
=�M=�q=| =���<� =K<=j�=��
=�=��=:=�~==c4==��=�Y=5=��=��=�G=��=�z=��=�=c�	=r0=�H =��<�!�<��<3X�<y@�<���< S�<���<���<��<J�<�a�<'i�<��<��<�(�<
��<!	�<O$�<��<�Ч<�<1��<���<��<�5�<��<n�<_M�<�ѝ<�8�<���<�(�<��<�<�^w<�i<��W<�C<)Z,<�s<�0�;���;���;K �;Y�~;/�;8�;�$�;���;q#�;��;3�;c49;��:$Mݹ�����DO��Ҁ�|���}��ȴq�k�L�{�'��������L���3��",��Q�^�z��(��=M���?��ջj3��J��X���Y.0��F��^���x�q��]~��0��� d�����Xꤼ���G���Yg������?���@���ϲ�羼d�ʼ��Լ�ۼ�O޼�(ݼ0�ؼ�0Ҽ�ʼ�Zü���؋��{���r��^+���v��o����������l]��&����]�������ͺ�K���,:ļϵ˼��Լ��ݼ[�����I��<��m�� ���(ۼ�hռ��Ҽ�%Լ�PټD[����S��"���_���S���̀������`���漦�߼Hiڼ��ּ�ռ޾Լ�Rռbּ�׼��ؼc�ټVۼT"ܼ�ݼu�߼l㼝�&％���� ����
�Fe�n6�G4�u�}j
�����s��8�V� �
<�ۆ��
�q���?��d��  �  �a=l=��=r�=�"=��$=��&=�/(=_*)=o�)=��)=ګ)=�f)=_�(=lp(=��'=��&=~&=��$=Ā#=s�!=Lt=��=�6=L�=0= =��=��=�z="C=��=��=uE=g�=M�=��=��==�8=�=a�=�G=��=0�=h%
=��=�s=��=�I=�^==Y=�~=}=�X=9=g�=�%=rr=�=�Q=��=�Z=�q
=b=�a=S��<&��<o&�<�<�F�<d�<�b�<���<e��<���<q��<���<J�<@Y�<���<wC�<=9�<;:�<��<^
�<P�<t�<Z�<s��<�ٯ<�í<��<O�<;�<���<�Y�<;��<`ӌ<9��<�M�<RYs<�1e<�U<'DD<o71<�.<�R	<�;w��;^�;T�;��;��;87�;���;�^�;N�;!��;>=h;Z>;<1:-&1������$�k�=��B��8�@'�ǋ�œ	���\�T!�G�:��Z�ݳ}�⚒�����E���Bxֻ�L�}���%��� ��a1���C���W�bm��Ѐ�3��q㑼b9���뙼�<��S���O;���`��@������U�����@���'����ɼ[�ϼxҼVҼ��ϼ��˼_�Ƽ\����_��g&������졶��ܵ��v���]��n���1���!���k���i���C�������P����ļPDʼF�мL�׼��ݼ� ��G�b�����༃=ڼ�bԼC�ϼ��ͼI6ϼ�ӼF?ڼo�἞c��7＾��3��C�"u�*��T��k�޼�9ۼ��ؼb׼�ּ��ּ�*׼<�׼��ؼڼ��ۼ�Mݼyo߼��YG���C���q��C���l��BO����E	�5N	�b��������M ��:��V����V���s��1��9
����͆��  �  6*"=N�!==�!=�"=��#=!�$=Z�%=C@&=*�&=`'=Y�'=`F(=փ(=lu(=u(=.'=��%=O~$=��"=�0!=�x="�=�=�=ee=oN=v�=6F=5�=l9==�Z=a=�=H�=ܾ=VZ=��=�=*!=�=e�=��
=.�
=��=��=�=�=H7=-=�=��=]�=�E=Z�==�=`�=,�=f�=��=�_=��=�p=`�=	�	=��=�=�r=��=L =(x�<4�<�
�<$* =� =K@ ="��<���<T��<5��<���<n��< ;�<R}�<!͸<��<Z��<C�<�į<���<x�<�)�<u�<rp�<���<�`�<lk�<��<���<�Y�<�=�<	�y<�j<�}\<K;N<��?<x{1<��"<��<'�<D��;'��;���;��;p��;{��;\��;�#�;���;H��;0��;��E;�0�:�P:��ϹL%��yغ"6 �C���y��Tp��&��4�$yE���X�Y=o����������������8�ܻ���!��ft�)�Ϩ7�(�F���U��e�p�s�a���ˆ�cQ���3������܏��揼����bҒ�/��˃��𐥼ec����zL����ü�Ǽ�Qȼ;�ǼF�Ƽ��ļbI¼93���V��U��������W��NⷼB׶�Et��wܶ�U������a��9�������ļB�Ǽ�?˼�ϼ��Ҽb�ּ�eټCۼCۼ�Yټ1ּq�Ѽ�ͼʲʼt~ɼ��ʼ�μ�JӼkHټ=߼����漗:���w����iu��a�Ǥ޼[<ݼ>	ܼ��ڼ��ټ?Bټ�ټ�ټ�ۼy/ݼ�߼�'㼪��%�鼓��`�8����
��Im��:.�������z������ ��
��
����[��LD�����k����m�;���z���
��  �  |'=��%=��$=�,$=��#=#=H�"=)�"=#=��#=��$=��%=��&=�H'=%�&=�%=�0$=�"=T�=�=�=Q===�f=I�={4=��=ʣ=<�=�5=�=�6=�g=�Y=��=r=�_=��=��=Kj=�r=)�=Ġ=��=�=�=�Q=�'=*3=�=L=ml=z�=W0=�F= �=�=Q�=��=W=�=45=Խ	=��=��=�=�_=i�=�=Ћ=3=O�=6�=��=�=o=B =���<[��<G��<���<U�<:��<���<7I�<�s�<E�<���< f�<��<�?�<Y��<#l�<4۟<r�<Ҥ�<<ۙ<���<j��<2h�<P�<r�n<��]<8)N<�@<�U5<�{+<��"<��<'�<b<��<�9<���;���;���;7�;ܶ�;KN�;*X�;ڟ�;.Mv;�*1;?��:�,M:�y���1��ۤ���躒��6/���H�K
_�[�p��~�a%�������[��Y����Ұ��5ʻB"�p���A�
�'���6��D��}O���Y�#�b�ѵk�@�s���{�g/��y����-��eU���;܋����!����S��(���H���D���}��������Ӓ��m�¼Fcļ{}ż�Ƽ�.Ƽ��ż�ļ���R澼���!������`���3ߺ�����e����ż,ɼ��˼��ͼTgϼdsмj8Ѽ4�Ѽ��Ѽ��Ѽ�ѼD�ϼ[ͼ��ʼ�Gȼ�Ƽ�Ƽ�Ǽ!�ɼ�kͼv�Ѽ�ּ��ټ5�ܼ�Q߼w�Y�⼉����伒��0�!��/[�a�Z߼8�ܼV�ۼ$�ۼ�Mݼ�W��r�	�C���l����� ������li���������oE��%o��{���
�������0n������)������������#���n��Ɍ�x������  �  �w*=~(=�W&=�$=��!=� =ܕ=�=�=�'=�� =0�"=Q{$=�n%=iM%=�#=��!=��=O�=��=��=��=�;=n�=�n=�y=��=T�=�J=3�=1�=�=9�=�=��=`}=��=_�=�+=��= =��=��=�=�=�=�+=��	=��=g�=Y	=x�
=R=K=�=c=��= p=�#=�Z=��=GC=��=8�=}=��=Ղ=�i=�%=-�=�=`^=P�=�=J�=�@==5��<E�<��<)��<��< ��<E��<���<�ʾ<�ȶ<��<�Χ<���<抜<.7�<|��<8�<8w�<p[�<'�<�T�<�J�<���<�Gt<�_<��K<T�:<S�-<r�$<�<�<�j<�G<3�<��<sQ<�a<u�	<'�<}z�;���;��;/��;¨;k��;�_;\%;���:�P:;���fx��L��*/��b������ߖ�雠��<������U(��Ć��Ύ��ܼ�-ػ����$�	�&��:�0J��:V���^���c�9qg���i�1ml�:�o�ˤs�p�x�p~��끼�����a����M��͈��O-������z����	��� ���
��l컼	���4�ż;�ɼ�ͼ!ϼ=xϼ<�ͼ��ʼ�SƼ���������m�����+�ü�ɼ�~μ$�Ҽ��ռ�׼*�ּ�ռ{�Ҽ�/м�ͼ+�˼��ɼ)ȼ��Ƽgiż�YļD�ü@�üV�ļ�Ƽ!/ɼ�̼�3ϼ�iҼ��ռ�bټH]ݼ����c��M��G��|�������q�弰9��߼�߼������F��b��(���ak���k��أ��U[��4
��%'�����}6��X����n���_���g�z��s������m���������R ���5 ����  �  �^,=��)=�2&=\�"=e�=έ=�I==�L=��==C=�=��!=�#=^#=�!=ڐ=F�=��= N=��=��=�=�=��=�<=��=��=WR=qI=��=�=��=�=`=��=�V=K�=��=�=t=��=)�=7�=�t=j�
=��=*�=K.=t�=��=��=��=��=�d=P�=>�=_�=�
=R!=��=�� =��<��<�`�<�� =55=ƍ=P�=L	=9�	=��	=��=�=��=5�=�K=&#�<�'�<ݵ�<v��<:��<#��<V��<0�<j�<�J�<��<^��<91�<��<�L�<�O�<�Z�<�]�<��<��<� �<�Ǉ<}<�Ef<>N<6A7<
[$<-< �<h�<��<'�<�m<N�<h<��<��<��<*[
<�<��;��;D
�;��;`��;�a{;��F;�~;�ݟ:IK 9��J~�Ya�pH��2����Ż� ϻz�λ�Ȼ�:��J𹻡Z��Zͻ�,�D	��� �}9���N��v`�o?l��>r�(ys��q�\Mn��Nk���i�k���n���t��#|�F���Ɇ�+���ZM�����e發����c���E��薭������s������ɼ)�м�hּڼ�!ۼ�@ټ��Լ��μ �ȼ�uü!���A����Wļ�Bʼ�vѼ�ؼzF޼��&I⼱N�$Wܼ�3׼J�Ѽ�̼�_ȼ]\ż0{ü&|¼�¼¼n¼aüZ�ü�/ż��Ƽ��ȼ=�ʼ��ͼʘѼ��ּ��ܼ���$����`�������|h��������$���輼�伪��o��]�꼧��s����� ��x���2�B"��2�u���1���V��\�`�����m�p�％�S��� ��X�j����������3����N���  �  t�,=�W)=J�$=" =^=Q�=�=%"=s=�t=�=#M=߆=�� =;� =�=a=��=p�=��=Y�
=��	=ߝ
=c�=�7=��=��=��=�=1b=��=��=\y=F�=�d=��=ju=P
=��=O�=��=�=��=0.=��=�=�= ��<g��<�{�<B��<,� =�o=�W=�=-K==h =uX=��=a��<���<ם�<���<D��<�,�<�	 =W�=L�=�.	=ko
=�
=��	=�'=�=G�=5=���<�,�<c`�<=�<փ�<���<��<��<C�<˯<���<�X�<��<z�<>�<?�<p~�<n2�<�v�<Ә�<�E�<o�<�xq<��W<�p<<ʚ"<~�<�1�;���;��;Ȃ <i�	<n�<��<�?<�<m9<T�<7�<��<��;��;И�;�S�;�ؚ;�]�;%W;�;���:x��8����o<��`��X�����޻h��>���c{���{���ܻ�qѻ˵л)߻s����B���/�OWK�d�RNw�������N���>�n�v��n�0�i���g��j���o�7x������-��ST���8��.�����_���0��g㥼�����ʲ��s���:ż`ϼ��ؼ ��-�弲�v��C߼�׼��ϼ"ɼ$�ż��żV�ɼ-Ѽ8�ټ���o��R��e��v����/eݼ^ռ��ͼ��Ǽ.�ü33��	V��u|���1��	#¼zü��ü<�ļS�żf�Ƽ(�ȼ~�˼м�lּ��޼��缴������ �L���#����Y��2�����꼄X�P����5���n�����H	�3�L�
�+	�t�0z��������������3x�n�C8��l�{���T=��Z������;/��1����6���  �  ��,=�{(=�.#=%O=v=�U=.�=��=d=u�=��=�=��=�<=�=!�=U�=e=��=�	=��=��=��=[�=)�=�=�$=~=��=*�=�I=�%=��=k�=4,=��=L=<=��=�(=�=��=�=�=�
=�=��<�,�<ޅ�<��<` �<՚�<'� =�M=�		==��
=��=@^=�v�<Q<�</��<�0�<��<q-�<���<D��<�j=��=�=�h
=y�
=��	=F=��=�i=?� =N�<���<@�<���<��<�+�<�u�<B��<�ٹ<�۪<7��<+��<Q3�<÷t<r�m<��n<�v<h1�<Ǆ<�݆<��<�|<�Lg<F�K<�K-<�<)��; (�;��;/��;x�;��;��<�<�K<w <�<P�<�<Ԩ<K��;�}�;TV�;�.�;F�;�-�;��[;"!;{�: �"���[�h������߻W��f���������c_�����*������I����<�F[��^v�&�����Y������7��|+��g�t��l�3�g���h�w#n���v�j����C��Ŭ��C�������^ߘ�����e�����ST���������?ɼ]ռ��༹���8l�E��缱�޼G�ռ�"μP�ɼ|)ʼ��μ�
׼�2�K뼏b�S����A��QT����C��%�ټ:Xм׻ȼpüޅ��ؘ����� ���m¼��üfpļu ższż�=Ƽ��Ǽk�ʼ�м�׼�p�i�켭i�������G��I�?a��������������`�$���A���XM�0s
� N��8�f������	�<H�� �����z��v�켞��u��m}�K%�e��S��v��wH��ʈ�����������  �  �\,=�'=��!=KI=�=�1=+=<X	=�	==�=�=��=�=^�=S=��=9�=r=t=��=�Z=�=�F=�=�C
=��=�=�Y=٣=�=S=�*=ҁ=̮=h�=e=P=l�=�=y3=��=]�=Z�=�=�	=:�=}�<��<ov�<P��<PL�<!��<to�<�?=WQ=^�	=a	=��=7Z=͋�<_^�<�R�<��<e~�<���<�,�<��<Le�<�c=��=�
=/�
=�	=2=-�=�!=�` =�[�<� �<���<%_�<���<���<ڻ�<3�<zP�<u�<B��<��<Ʈv<�Jf<�n_<��a<Ͻj<��v<0�<���<���<S�v<^T`<!C<:#<)�<J��;���;�k�;��;[)�;�}�;e<.�<��<��<�<�<�E<X�<���;f�;� �;K��;�s�;^��;�[;�r;wI�:�fù���[���F»��������N� ��m�Og����{)���O�Y�������&��E���e� f���d������6��A��a��Dփ�R�y���n��i���h��m���v�ƀ�����I������Z�����b���xE�����!�����������ej̼_�ټ>\����������z4�������ټ��Ѽ	ͼ�9ͼ�2Ҽ7ۼI漦#�>��5��DX�����O��B�rݼ,�Ҽ\�ɼ1�ü����󂿼4���U���¼�ļ0�ļ�\ż+�żH7Ƽ�Ǽ˼��м�ټ|�㼝[��H������	����
����	�$��6� �%���T򼀾��A�T\�����������޷���jp�������`���Ĭ��~a󼡾�����������&���e������q`��sx������� ���  �  `,,=J'=�>!=&�=v�=�=��	=�=V�=�=�=�=@i=�=�v=vZ=�=J=�#
=F�=m=s��<�=�s=BZ	=-�=�a=�=�z=	�=�M=�%=v=0�=c�=nK=� =�=b�=a/=S�=�=�=G�=��=��=rs�<<H�<���<%q�<���<`��<~��<��=��=��=*�=<=�=V��< K�<s��<��<���<*�<��<+P�<��<��=�=��	=��
="�	=;%=m�=m=I@ =A�<���<R��<�I�<6��<���<�i�<���<�\�<�¥<y��<Ty�<��q<�1a<�nZ<�]<��f<��s<�#<�q�<>�<Z�t<�]<�@<�d<Ep <L0�;�; z�;"��;-V�;}L�;��<�<B�<�{<�<V�<�<��<]��;�-�;�@�;��;T�;ž�;�yZ;I�;��:ط�C�x�����ɻ��t�,�"�U�%������������:��>��G�Q�)���H���i�����rԎ��3��q��:8��<ꌼ�9����{��p���i�-i���m�Z�v��܀�u���GH���C��6����*�������J��/&��!㫼 ����n��B�ͼ!jۼ#c�b���n����������Ｄ�弍Aۼg�Ҽn#μ�Rμ�fӼ@zܼ3��5�?^��k� ��� �uS���������D޼�\Ӽejʼ�#ļ���\�������r����¼pIļ�ż]�żd�żvBƼx�Ǽ	˼b�м��ټ���ٴ�������U
����B��
����>��_���0C���`�f���{�����ƚ���.����������J%� ���f���������K�����k��1F�H������Gt��;���b���#+���  �  �\,=�'=��!=KI=�=�1=+=<X	=�	==�=�=��=�=^�=S=��=9�=r=t=��=�Z=�=�F=�=�C
=��=�=�Y=٣=�=S=�*=ҁ=̮=h�=e=P=k�=�=y3=��=\�=Z�=�=�	=:�=}�<��<nv�<N��<ML�<��<oo�<�?=SQ=Y�	=a	=��=,Z=���<>^�<�R�<^�<+~�<���<{,�<[�<�d�<�c=y�=�
=d�
=��	= 3=��=�#=`c =�b�<0)�<���<�j�<���<��<���<.�<�a�<U1�<*Ж<���<��v<>jf<��_<)�a<D�j<�w<H�<���<O��<F�v<�J`<�
C<��"<��<���;���;�)�;�h�;:��;X6�;f�<�`<Za<��<S�<�<�5<z�<5��;}�;�*�;c��;%��;<#�;t[;��;�D�:G,������d�����)����e�%���� ��T��R�������E�/�����r'���E�N�e�s��ts��0�������}.��s郼�y�uo��5i��i�I�m���v�mр�v���l ����P`����������G��l��E���g���=����j̼��ټ|\�#�����5����4�������ټ�Ѽ$	ͼ�9ͼ�2Ҽ9ۼK漨#�?��6��EX�����P��B�rݼ,�Ҽ\�ɼ1�ü����󂿼4���U���¼�ļ0�ļ�\ż+�żH7Ƽ�Ǽ˼��м�ټ|�㼝[��H������	����
����	�$��6� �%���T򼀾��A�T\�����������޷���jp�������`���Ĭ��~a󼡾�����������&���e������q`��sx������� ���  �  ��,=�{(=�.#=%O=v=�U=.�=��=d=u�=��=�=��=�<=�=!�=U�=e=��=�	=��=��=��=[�=)�=�=�$=~=��=*�=�I=�%=��=k�=4,=��=L=;=��=�(=�=��=�=�=�
=�=��<�,�<ۅ�<��<Z �<͚�<"� =�M=�		==��
=��=,^=�v�<<�<���<c0�<���<�,�<&��<���<Hj=F�=��=�h
=��
=��	=�G=�=Sm=R� =?�<}��<*S�<��<F�<�G�</��<þ�<_��<���<�ڛ<$؍<�S�<��t<%�m<��n<CGv<�A�<�҄<P�<y��<>�|<e:g<<fK<�&-<��<�P�;���;���;OX�;���;�~�;8�<��<><7@ <�<��<Qc<��<$��;*|�;
i�;�U�;���;�z�;�J\;�;�Ч:oZ�����lg��{���D߻d]�`�t��������!���廌⻪�ﻗ�����t=�H[�ʐv������؋�.|���>���\���P��nu�uTl�#h���h��[n�%w�aƀ�zV������0������r瘼:���Pj��/ ���V����������?ɼ�]ռ ��	�H��nl�n�����޼Y�ռ�"μZ�ɼ�)ʼ��μ�
׼�2� K뼐b�T����A��RT����D��%�ټ:Xм׻ȼpüޅ��ؘ����� ���m¼��üfpļu ższż�=Ƽ��Ǽk�ʼ�м�׼�p�i�켭i�������G��I�?a��������������`�$���A���XM�0s
� N��8�f������	�<H�� �����z��v�켞��u��m}�K%�e��S��v��wH��ʈ�����������  �  t�,=�W)=J�$=" =^=Q�=�=%"=s=�t=�=#M=߆=�� =;� =�=a=��=p�=��=Y�
=��	=ߝ
=c�=�7=��=��=��=�=1b=��=��=[y=F�=�d=��=ju=P
=��=O�=��=�=��=0.=��=�=߃=���<a��<�{�<:��<&� =�o=�W=�=K= =Q =YX=��=��<p��<T��<#��<���<%,�<	 =�=��=@.	=~o
=��
=f�	=E*={=��=g=��<}C�<}{�<�\�<§�<���<\��<�?�<%�<���<�ʢ<���<L�<��<pe�<�.�<���<�I�<6��<4��<�G�<�܂<6_q<R�W<<<<�Z"<�L<���;� �;i��;�! <�$	<��<%h</�<Ub<��<n<��<��<���;Q�;k��;��;�+�;˄;�X;Q;��:H��8���:�#������(޻l����4��,����W�ܻ�7ѻR�лl߻����}b��0�\�K�bd�۟w��Ɓ���Eꂼ�t�g5w�odo�	�i�2-h��lj��2p�a~x�����H���j��FK���Д�Q��
��"7���祼�����̲�'u��<ż�`ϼ��ؼ��༒���缱��p߼�׼��ϼ$"ɼ2�ż��ż^�ɼ3Ѽ=�ټ���r��T��f��w����/eݼ^ռ��ͼ��Ǽ.�ü33��
V��u|���1��	#¼zü��ü<�ļS�żf�Ƽ(�ȼ~�˼м�lּ��޼��缴������ �L���#����Y��2�����꼄X�P����5���n�����H	�3�L�
�+	�t�0z��������������3x�n�C8��l�{���T=��Z������;/��1����6���  �  �^,=��)=�2&=\�"=e�=έ=�I==�L=��==C=�=��!=�#=^#=�!=ڐ=F�=��= N=��=��=�=�=��=�<=��=��=WR=qI=��=�=��=�=`=��=�V=J�=��=�=t=��=(�=6�=�t=i�
=��=(�=H.=p�=�=��=��=��=�d=>�='�=C�=��
='!=Y�=z� =z��<-��<�_�<>� =�4=<�=ז=		=_�	=Ŏ	=u�=��=O�=׿=�T=�9�<�C�<*��<@�<K��<"�<f��<sh�<"<�<}��<'٩<K�<�i�<�<�|�<|z�<�~�<�y�<��<��<S�<>��<��|<�f<*�M<��6<��#<;�<�J<K\<�T<tp<��<�d<]�<�/<�L<os<�%
<2�<��;��;
+�;�&�;�"�;an|;�8H;��;w'�:q�<9�Q����%_�Y������k�Ļ
Aλ�*λ�yǻ:Ѿ�V���8��ͻU�mj	��!��M9�MO���`��l��r��s�r��n�g�k�soj��k��8o��u�K{|�Zl���ꆼ�����c���/��t���,����j���K������ݟ���u�������ɼ�м�iּ�ڼ�!ۼ�@ټ��Լ��μ@�ȼ�uü3���N����Wļ�Bʼ�vѼ�ؼ}F޼���(I⼲N�%Wܼ�3׼J�Ѽ�̼�_ȼ]\ż1{ü&|¼�¼¼n¼aüZ�ü�/ż��Ƽ��ȼ=�ʼ��ͼʘѼ��ּ��ܼ���$����`�������|h��������$���輼�伪��o��]�꼧��s����� ��x���2�B"��2�u���1���V��\�`�����m�p�％�S��� ��X�j����������3����N���  �  �w*=~(=�W&=�$=��!=� =ܕ=�=�=�'=�� =0�"=Q{$=�n%=iM%=�#=��!=��=O�=��=��=��=�;=n�=�n=�y=��=T�=�J=3�=1�=�=9�=�=��=`}=��=_�=�+=��==��=��=�=�=�=�+=��	=��=b�=Y	=p�
=H=K=�=O=��=�o=h#=lZ=e�=�B=��=��==
�=@�=Bi=)%=�=!�=\_=]�==��=�G=�={��<l4�<G��<���<K��<���<���<��<b�<��<�G�<Q�<�¡<�Ŝ<�l�<Ͽ�<�_�<���<�q�<���<�W�<hC�<��<t<�9_<~mK<�k:<�E-<j2$<Q�<o�<��<z�<zS<P<�<�<(�	<.U<�'�;��;���;���;]�;�	�;a0`;�&;���:LpW:ei%��p��	��-���_�������.Ɵ�������!���!8���h��#߼��=ػ)����b�M2'��h:�s�J�N�V�� _�;�d�H h�c�j���l�p�i&t��y� o~�����:������+��f�����=�����j���R��U%������������ż:�ɼ�ͼ�!ϼ�xϼ��ͼ;�ʼ�SƼ����5��&���m�����3�ü�ɼ�~μ(�Ҽ��ռ�׼+�ּ�ռ{�Ҽ�/м�ͼ+�˼��ɼ)ȼ��Ƽgiż�YļD�ü@�üV�ļ�Ƽ!/ɼ�̼�3ϼ�iҼ��ռ�bټH]ݼ����c��M��G��|�������q�弰9��߼�߼������F��b��(���ak���k��أ��U[��4
��%'�����}6��X����n���_���g�z��s������m���������R ���5 ����  �  |'=��%=��$=�,$=��#=#=H�"=)�"=#=��#=��$=��%=��&=�H'=%�&=�%=�0$=�"=T�=�=�=Q===�f=I�={4=��=ʣ=<�=�5=�=�6=�g=�Y=��=r=�_=��=ߓ=Kj=�r=(�=à=��=�=ߤ=�Q=�'=&3=�=�K=fl=p�=J0=�F=�=ڌ=1�=��=%=q=�4=z�	=�=%�=i=V_=׼=_=��=�=g�=g�=?�=
$=,"=]L =��<���<��<���<#��<���<f7�<���<��<o��<h�<��<`٩<}�<���<��<J�<q��<���<8�<U��<߹�<|V�<��<�@n<0:]<�M<�K@<F�4<��*<$="<Xh<0M<��<�E<;�<&�;.�;�{�;P��;���;�J�;[~�;8�;#;w;
c2;h��:�T:�2�7�(������T�1���-���F��]��o�l�|�e�������
���Ν��հ��cʻ�y�o�����T(��l7�4�D�P��:Z�J�c��Jl�}t��|��r���;��jf��7!���҉�\���/��b����h���'���U��"N������#�������p���V�¼�dļ�~ż�Ƽ�/ƼT�żļ\����澼���>���(���p���?ߺ�����l���
�ż
,ɼ��˼��ͼUgϼfsмk8Ѽ5�Ѽ��Ѽ��Ѽ�ѼD�ϼ[ͼ��ʼ�Gȼ�Ƽ�Ƽ�Ǽ!�ɼ�kͼv�Ѽ�ּ��ټ5�ܼ�Q߼w�Y�⼉����伒��0�!��/[�a�Z߼8�ܼV�ۼ$�ۼ�Mݼ�W��r�	�C���l����� ������li���������oE��%o��{���
�������0n������)������������#���n��Ɍ�x������  �  6*"=N�!==�!=�"=��#=!�$=Z�%=C@&=*�&=`'=Y�'=`F(=փ(=lu(=u(=.'=��%=O~$=��"=�0!=�x="�=�=�=ee=oN=v�=6F=5�=l9==�Z=a=�=H�=ܾ=VZ=��=�=*!=�=d�=��
=-�
=��=��=�=�=E7=�,=�=}�=T�=�E=K�=*�=G�=�=?�=W�=�_=��=;p=��=��	=?�=c�=-r=��=. =�x�<\6�<��<�- =H� =�G =��<J�<���<���</��<���<�q�<���<;�<�7�<YŲ<G3�<��<�Ү<jK�<�_�<��<��<�ã<w�<�w�<���<cّ<�H�<0#�<=py<�j<t\<��M<�y?<�0<�t"<�f<�o<G��;���;T�;M��;�L�;�\�;�3�;���;K��;\��;5ъ;U�F;���:�!:D¹/v��րԺYB�����.����ps���$�K�2��D���W��Tn��τ��������� »�ݻ���������~)��#8��G�LV���e�R�t�Q'�����h���Yp��1ŏ�����������i񒼨5��;���󠥼�o��
���JS����ü#ǼsTȼ$�Ǽ��Ƽ��ļ.J¼�3��W����������W��sⷼ]׶�Zt���ܶ�a������a��>��"�����ļD�Ǽ�?˼�ϼ��Ҽc�ּ�eټCۼCۼ�Yټ1ּr�Ѽ�ͼʲʼt~ɼ��ʼ�μ�JӼkHټ=߼����漗:���w����iu��a�Ǥ޼[<ݼ>	ܼ��ڼ��ټ?Bټ�ټ�ټ�ۼy/ݼ�߼�'㼪��%�鼓��`�8����
��Im��:.�������z������ ��
��
����[��LD�����k����m�;���z���
��  �  �a=l=��=r�=�"=��$=��&=�/(=_*)=o�)=��)=ګ)=�f)=_�(=lp(=��'=��&=~&=��$=Ā#=s�!=Lt=��=�6=L�=0= =��=��=�z="C=��=��=uE=g�=M�=��=��==�8=�=`�=�G=��=/�=g%
=��=�s=��=�I=�^==Y=�~=}=�X=#=K�=�%=Gr=͉=~Q=7�=QZ=�q
=�=ia=m��<��<N&�<��<�H�<h�<$i�<;��<���<ܝ�<`��<���<<�<m��<Q!�<�t�<�n�<�r�<�I�<cF�<��<A>�<l��<6�<�	�<��<uӪ<&��<꒢<Ь�<U\�<´�<+Č<���<C.�<ss<�d<�9U<D�C<��0<x�<��<�"�;���;;.�;�.�;:�;ۓ�;bʼ;}t�;7�;�;���;7�h;6;ED5:�+�}���##���;�'+@��66��%�P��T��u�����	 �K�9�=Y��(}�y��p����̾���ֻ������|��L!���1�lKD�R|X�|�m�k���r��� ���s��7"��Yn���!��b�����1���ț��͢��'��T�������5�ɼ�ϼi{ҼoXҼc�ϼ�˼Y�Ƽ���e`���&������'����ܵ��v���]������?���+���s���o���H�������P����ļRDʼG�мM�׼��ݼ� ��G�b�����༃=ڼ�bԼC�ϼ��ͼI6ϼ�ӼF?ڼo�἞c��7＾��3��C�"u�*��T��k�޼�9ۼ��ؼb׼�ּ��ּ�*׼<�׼��ؼڼ��ۼ�Mݼyo߼��YG���C���q��C���l��BO����E	�5N	�b��������M ��:��V����V���s��1��9
����͆��  �  �l=~�=�=��=d�=L#=!x&=m�(=�9*=��*=i�*=�K*=��)=�)=i(=S�'=~Q'=��&=�%=.�$=̼"=��=�6=@�=��=�=I�	=$$=��=�=�	=�o=R*=�U=�(=	=?=|='�
=�M=�q={ =���<� =J<=i�=��
=�=��=7=�~==]4==��=�Y=#=��=��=�G=��=�z=p�=��=�	=0=sH =��<<!�<��<�X�<?B�<��<TX�<���<���<v$�<O]�<y�<ʄ�<�"�<9,�<Q�<�ϧ<I7�<ST�<�P�<��<3�<)ʯ<��<��<TX�<���<���<^]�<�ڝ<�:�<M��<A�<ۏ�<�Ё<�w<�h<�W<U4C<��+<e<jm�;���;I��;�S�;��};;��;�ō;�˝;澪;��;v��;�	�;��9;�H�:Xֹy����N�&��:�ú��*&p��LK�2a&�L�	����q����&��E+��YP�rz�g��uO���_��NKջ��ք�������0�DdF�� _�t�x�@��A���b�������o᥼���7��Ξ������Ӝ����O��p۲�4�B�ʼ��Լ܇ۼWR޼�*ݼ��ؼ�1ҼïʼQ[ü��0�������3r���+���v������������u]��-����]�������ͺ�M���-:ļе˼��Լ��ݼ\�����J��<��m�� ���(ۼ�hռ��Ҽ�%Լ�PټD[����S��"���_���S���̀������`���漦�߼Hiڼ��ּ�ռ޾Լ�Rռbּ�׼��ؼc�ټVۼT"ܼ�ݼu�߼l㼝�&％���� ����
�Fe�n6�G4�u�}j
�����s��8�V� �
<�ۆ��
�q���?��d��  �  �5=�=�d=BZ=n�=�!=	�%=W�(=Uv*=�*+=�+=o*=��)=��(=)(=��'= L'=[�&=j=&=�%=<�"=�=�8=��=��=�C
=	e=b=%� =�=�=��=�=W�=��={�=V�=��=�i=2=nF�<'��<+k�<3u�<�<��=�=�==Y9==��=F~=�x=1=��=5=?�=\�=��=��=�=��=>�=�(=��=^=�L�<\�<��<�z�<�*�<���<BV�<'f�<���<`�<*�<6�<$��<X��<���<���<թ�<O��<7�<�6�<6��<�:�<c]�<O��<�O�<Su�<�#�<#­<���<^]�<M|�<ԫ�<�<�ӌ<���<zD�<�Tx<�ui<��V<��?<�n%<n�<���;��;)t;$�>;ҩ+;��7;6�Z;%�;*�;��;���;9�j;A7;z��9p����EG��ʎ�������ؕ���g��*�t�Ə@�f��*������n���&��
O��F|��k���$������zֻ�&뻹� �h�����$(2�|�J��f�c�����$��m���������.��J����/���¡�if��Y(���-��	����Ƽ�KӼ�s޼�弆�����z)���ؼXϼ�Ƽ	K�������$��:���v���GV��J?��.���~���������+඼ҷ�%��}��A9ż0Aμ��ؼo?�����L���P��M������h����l�YIڼ@2׼O�ؼ�_޼��`=�����P��{��z��h�i{���P�����]�Iۼ[�ּ^Լ�Լ'�Լ�aּY�׼�Xټ}fڼ-ۼ��ۼ��ܼ��޼��gV�g~�����1��	��^��X��k��O�Z&��z��(
��2�k��8��Ӈ��6��M����J��ox��  �  �=+^=�F=��=�=!A =��$=�C(=�[*=;2+=7+=�a*=�w)=��(=o�'=t'=�)'=��&=:G&=�%=��"=�-=DI=^V=��=�=m/=d�<�l�<���<\y==��
=��=�Z=~i=I=I�
=�
=r|�<��<��<`L�<���<_/�<�%=��=r=��=P�=��=)�=]{=F�=�a=��=��=��=��=f�=)=$�=�_=q�=(q=�X=��<�Q�<��<�z�<�5�<cD�<˭�<B��<$�<(��<)�<0K�<m�<��<(	�<���<i�<���<�K�<Kђ<I4�<��<mJ�<�ѫ<CS�<�#�<�,�<-ݭ<��<*�<�
�<!�<���<�m�<�r�<�:�<�Jx<b�h<`AU<��<<� <�� <	y�;��;�
=;��;}��:E-;<"/;[b;�|�;U^�;�8�;�1R;O��:m�S�����qx�򩻆7Ż.H̻/��&���"EV�-w#�W���=���J���&�-P��������Ļ�&ػ^��� �a��f���O4���N�4!m�ź��:����~�����RP��+ٶ��S��13���{���U��ݐ��P?��a���������ʼQټ弡���Ｌ��D缣�ݼ��Ҽȼ~����#���=��B���(����������ꄶ���������ڶ��඼�����2������`sƼ�{м�]ܼ���#���b���V����� �kr�����_ ��ݼZAڼ��ۼ�἟��&M���I����
�j �K��W���������H ��(ܼO�ּ�]Լ�Ӽ[�Լz�ּ�aؼF�ټ��ڼ��ۼtܼ��ܼ.�޼ɽ⼩	�A�Ib��������o����H��Y��XT��8��m���t(��k���
�������5�����  �  lH�<���<���<��<X5�<���<0�=��=	K='�=�<=Q�=B�=N=�v=��=|=��=�#=��=f=|=t�<���<��<�޳<j��<���<8ő<���<\�<��<}��<?�<C�<��<���<���<ݵ<��<�W�<��<F,�<�Ջ<�Й<��<a��<'G�<�:�<�]�<�# =v,=7�=2@=`L=M)=��=^�=�C=a^=��=�r�< �<C�<���<��<�E�<�1�<�|<��h<��d<��p<ҫ�<?�<JA�<���<r9�<¡�<Jv�<_��<�R<� !<�(�;�;�.�;��;8��;��<��:<��Z<u<�k�<��<f��<O"�<�ׁ<�y<ٝm<�a<~YU<|-H<q�8<S�%<��<},�;Iч;� �:���0F��^Y�������/�E(1���"�_	���׻�u��Ԇ��f��{����D�E�$���U�B_���,��$暼����o���(��pe�E�A��}"��`
�&L���=����q�����r��u0��"'�i�3��'A��{Q��f�"�������1��������ڼ���¸��h���,��v��^,���������3�W𼒤��������)?���&���,��|.��+��%����t���S�׫��m�4Z�}޼��ڼ�ټ/Tټ�xټ2�ټ�=ڼ�ۼ��ܼ&��U9缼���; �Z�	��Z�͈���)���1��]6�9�6�ɵ2�>t+��n"�;��������8m��r�ů�'�'�4=1���8��<�L5<�)�7���/��&� �����s�	����K������u9���3�����������+�������f��J?�����4�������H,!�
�,�.�7�B�A��I�W�L��K���F�V�>���5��-��3(��s&��(��[/���8��B�n�K��R��  �  ��<��<*��<�K�<m��<Q�<�=�/=MU=��=�!=�=m=L�=h==�==��=�	=��=�(=�b=AB�<<��<:��<;;�<|�<�ۙ<7$�<�ɚ<^��<M,�<���<a\�<��<\�<h��<$s�<�޸<��<�^�<6j�<���<E��<�t�<���<���<���<��<O��<�" ==ޘ=I(=�9=�=L�=ޟ=&,=�B=�o=<g�<oC�<�<���<!��<%#�<���<g|�<zjq<�{m<r�x<�8�<H�<��<�<}�<Ɇ�<Q��<�*�<��X<{[(<� <���;C�;4��;v6�;D'<+\><�C]<5v<���<Ƈ<�D�<��<ϧ�<��x<�im<�|a<� U<��G<�8<�}%<��<�,�;S��;+��:�ĺo�����3�8	'��(�f��u��1̻�ޚ��<}����������0|�.JO�1){�z���������J������f�`���>��� �D�	�Q��u�黭����������P�:C'�(�3�vbA���Q�\f�rĀ������림�Ⱦ��ؼ?r𼍵��8
����%��y�	�����������#��U��w����ju�4u��$�1�*��L,�6�)�TK#�l��k��������[�
F޼�ۼ��ټ�xټ�ټ�ټ�aڼ�Aۼ�ݼ���mB�go����u���I����(��/��04� w4�Ӭ0���)� � �Q�=��]���m�T�:[���%�*`/���6��k:�::�L�5�-#.�?�$�q���S��v	�f���_��U���n���_��+�����WK��Я��g���pZ����y.�SL�?s��Z ��R+�BM6���?��G�ORJ� tI�T�D��!=�+q4���,��)'��y%�'�'�{-.��7��A�J�|`P��  �  ���<���<u�<��<�L�<L^ =�;=N�=W6=� =a�=w,=�=��=F1=�=�=br=�=�=�"=�=^�<"��<T��<�x�<-r�<�<8u�<ś�<	^�<�`�<h[�<b��<j��<��<���<���<�b�<��<7��<뙗<�ʕ<�}�<_��<�̷<?��<�y�<��<��<>��<J�==��=R�=��=۬=nV=c�=M�=�� =��<��<���<�V�<��<a�<z��<~ȍ<?΄<nւ<]Ӈ<D�<�c�<���<��<�m�<��<��<�m�<Pj<a�<<x�<L"�;U��;KQ�;�#<&�+<�RH<�c<�x<�|�<M��<Y=�<��<��<��w<��l<��`<�T<�{F<��6<�$<�t<��;���;�;lF7��:_�������H9��=�7����ݻ���������N�0*V��퍻u ͻ/���<��e��?������ 늼=@����p���S�Y6��������>���)�nvﻦ����-�m�����{�'�O�4�зB�#S��vg����隐��ܣ�'�����м�缽K��^!�S����05�N�����	��T�^��^T���*��f����;�$�;'&���#�p>�]�x�J������۩����`*߼;ܼ?�ڼ�ڼ�ڼ�TڼF�ڼ@ܼ�޼���`���#�/
���%��x�*�-#��*�7.�IY.�V�*�7�$�����������֙�(�Ė��{!��*���0�yE4���3�k0��h)�� !�q���3�����c �����W��������Ŋ��G���+P���6 ����Wi��X�s���U�KC��"(�U2��:�� A�[*D�kC�?"?�E8�"Z0��")��7$��"�%���*��3�c=<���D�baJ��  �  ��<���<��<�7�<���<F�=�P	=�~=(S=��=�_=�=�J=�!=��=��=c�=vO=�C=,a=+b
=�= ��<r��<m�<�P�<|�<�Y�<���<��<6�<��<{��<�a�<�@�<F��<M��<S�<�	�<���<���<و�<欧<W�<���<��<�a�<��<)/�<ID�<	��<iW= �=��=13= P=�=��=��=��=�L�<���<s�<���<��<%��< l�<�>�<s��<Zj�<7��<L��<�#�<���<�$�<l��<}J�<�߶<x��<P4�<%(�<Y[<�t9<L�"<��<�X<�*<F�><�T<#�h<#(y<9��<���<1��<���<�0~<�<u<��j<��^<�EQ<�B<e\2<#�<*	<!��;_�;n�-;���9���޺���1����ӻP�ػ�ƻD���Kv�us/�eH
�9�&�X��W��p9��� ��E���a���q�t�+�j�=Y�.�B���+�X��}��)����#���r��Й�/	����v��)�5�7�*�F�}�W���k����L��ᾠ�zi����Ƽ!�ټGl�O������qi��v`��n��t�NM߼��ܼYP�p=��i�����a��������.����� ����g�	�_��@���Ey����̺ἃr޼l�ܼ�~ۼ@#ۼ�jۼTWܼ��ݼ�n�&D�J�p(���?������0��!��.%��Z%�[k"�,��X��S��
�˜�8k��t������{K"�N (��>+��4+�o,(�!�"�c�%��J<�(���6�C2�1�������x���A���s�������A���TD���ӭ�!K	�u+�Wg�@��r�#��#,��Z3��8��);�v�:�W�6��1��F*��$����=���� ���%��"-��&5�[d<���A��  �  ���<�2�<���<���<� =��=�<	==�=�=�2=�=��=�=
�=��=Z�=�=�=,�=��=�'='�=i��<��<'�<��<8�<��< E�<EX�<���<n�<R1�<���<<�<yX�<f,�<=i�<���<"�<=�<B�<=�<���<Q��<���<���<���<8��<��<y��<S�<�v =�=��=� =�=k/=�� =JT�<���<�b�<�s�<K��<���<҂�<]��<�θ<��<`�<��<��<��<���<_L�<��<�_�<��<
�<�ͣ<�b�<x�~<\�`<̖K<y�@<χ?<��E<�/Q<*&^<$ij<�Gt<S�z<}~<AG~<��{<��v<��o<�Kf<q	Z<_fK<��:<��(<�f<= <_�;7!�;��I;b��:��m��k�R�����*��3�s��A����d���lj��g��� �Nur�;˺��` �W| ���9��I��XN���J��@��3�
�$��`�������Y@����i�	�--�����R!��S.�}�=�3�N�a�L-u�߲��)�������m������5̼}�ؼ��O輣�輱��+�߼��ؼ#�ӼE�Ҽ�ּ~�߼��켳���Z�֨���>���J�Y���I��b�Zq������(�I��k��F�ci�{o޼�{ݼ��ݼ�2߼_��q/�5��%���1����O���	���Q���������V��d���@	�K�����3��*��m���S%�D�	� �<D!��n�����L��d�%��M�	��\�>��"��)� �v����������?/ ����U�5���\�.�����ݪ��:��6 �p#&��Z+�j$/�C�0�{:0�&G-��(��##�7&�J��2������ �j%&���,�\�2�H7��  �  ��<�F�<�~�<�Q =�o=��= =�T	=Q�=��=�=P~=��=�=�}=@G=�+=�n==Y
=�=z�=v =+�<��<!�<���<T��<���<���<���<�x�<Q[�<]��<��<�� =6� =P��<���<���<��<M��<���<���<"��<� �<m�<Q�<�N�<�~�<���<�x�<NP�<���<�+�<J1 =E=�� =�n�<��<��<���<�#�<,�<�<ԓ�<h��<yL�<�0�<�S�<y�<.1�<(��<x�<��<x�<r��<�G�<�<v�<Bn�<ü�<�Y�<<��<�Ds<��e<:a^<�I\<\�]<�e`<Y�c<4�f<Oi<E?k<Bzl<�l<Wk<��f<�V^<��Q<�AA<b�-<�<3�<��;PX�;Ë;֋G;  �:9n?:6߇�d��t�º��Ϻ�����:`�����C9q��9��V��x�!g�����B&��5�������!��+�iW.��`-���)�H�%��M!�O�����f���H�)[�q�����(���6�lH��\��q��:��wύ�gF��������-4������b4ɼJ�ϼkuӼ�[Լ��Ҽ�ϼ0˼b|ȼ��ȼ)�̼�
ռ_Z��h�\��3������	�/�	�e��r�.���8��?��������	��2���+v�e�Ἦ�Ἵ伭��M�켇��R��*F���2�G\�f��%�����ۇ�Ba� ��̒������W��1���&��,~���z�-����
����a��y������~�m�
�����;������
�Up�<R��X�������}��X�+�D����	�`��9������e�����q!��O$�~C&�[�&��&�%�#� ���
4���=+���<�;��g$��M)�'-��  �  �U=XT=��=^�=�_=6 =W=�)=�=_�=��	=c�=�=�b=�d=C�=��=�>=�0=V[ =�.�<v�<^e�<B��<)6�<�?�<��<���<���<N�<Y(�<&��<�d=
�=G=��=7U=�h =�g�<E��<]a�<�e�<���<9��<<��<��<)�<��<��<S��<���<|T�<���<���<u��<B��<�k�<*�<z�<d�<��<�h�<:��<)��<�#�<�B�<���<u%�<���<)&�<�n�<J��<���<���<�/�<h��<���<���<�q�<.��<�g�<\:�<�<Ky�<ѭ�<�u<�i<6`<ZX<��R<E�N<pN<p�O<�S<�7W<a�Y<f�X<�'R<�'E<fI2<_:<�b<CT�;���;���;�K;�;ſ�:^�:�:�-::9c:Q�:�,F:3c�:UJ�:N�:���:+Dm:���8x�����&�z��������3޻�� ���Sf��n#�"�*�2�0���4�P�6�Z�5��*3���.���*�}�(�n�+��-4�#+C���W�،o�)?��2������녣��Ȫ�=���ȫ��>鹼�z���7�������S¼���9-��'����e�����F�ļ*�˼l,ռ��߼�^��������� �i�+{��Q����Ж��������V�R����u������Q輍(�cV������W�����������	���	��G
��h
��'
��a	����M��g������������ ��j#���S��H����������%���!������.�nw��W�����M��:����	�L�� !�]�����l�R���������
����p���o�Aq����d�hC���L"����V�dy�����W��If����������� ��4$��  �  �q=r�	=m=��=$�<"��<z�<P�<���<`��<c1=�L=^�	=�=�R=�o
=]�=,�=���<3v�<�o�<8x�<���<�L�<���<�D�<��<���<6y�<���<�*=�E=�+=��=�V==~�=�=�=�,�<���<U��<�J�<*��<��<��</��<m�<Q�<T%�<R$�<|��<߁�<�H�<?l�<X�<q&�<���<��<�t�<@��<���<@U�<w��<�v�<q(�<,�<Z��<m	�<c��<v<�<_��<��<�R�<F��<��<���<���<�J�<�B�<�-�<鬭<e&�<Ȗ<��<���<��k<y�W<J}E<��6<��-<��)<U,<�E3<R<<+D<]�F<B<S�4<��<ly<vc�;�ɒ;�F;�-;���:w!�:vώ:���:���:�=�:��;��;&�;	?$;��%;��;�
;���:��Z:��E��ĳ�x�,��A��ξ��ŀһ2��� �\l$�T�6��;F��R���X���Y���T���L��WC��<��<�[�C�w�S�a�k�Z2����%���1���h������Mƹ�c����{�����"ѵ�:촼hc��`,��pL����|��l�����4�ļnU̼��Լd�ݼ*0��j�MY��%��:��*D��S	�r�� ��x4�N%
�e��(M�����]��P��e𼍭���Z��������i��v� ���D�����=	��c���s]������Z��� ��>�������� ��~���#��l#�hP������
�:L������=��J
�t���'���o��O�'i�e�	������	��(�����<�����s"��j#�E�"�)�!�uz��)��������b�(E�C:��X�Y������v������_��B��k��  �  ==�=�Y=�S =���<\��<���<-�<�I�<t��<K��<���<�=$=7�=M[=
� =���<j��<��<���<+��<� �<s�<@��<}I�<���<w��<��=e=�=I[=�	=�>
=�{
=E%
=�5	=F�=��= {=�� =A%�<1��<h��<�Y�<���<|��<8W�<\C�<ҿ�<��<H��<m��<�,�<���<Y��<���<��<�3�<>��<[��<m��<�α<��<�ֳ<u��<)��<��<E�<��<�-�<��<w{�<	��<8�<mo�<� �<p7�<���<5�<���<�,�<
��<�0�<k�<j��<,1d<�E<*<p�<�<-~ <(�<��<~R<�i+<9M2<@x/<�f!<?�<o�;�;`�;Ԋ:��h���D�ÇF�6�!:�@�:��;*�>;f1Z;~�g;�xh;�^;��K;��/;��;�8�:u��9v��ڦغ�B:�T뇻Q���뻜��7/��kK��.d��v�i����*��" {�,�m�H�^��.S��O��}U��-g�LS��r0��Y£�\��������Ƽɼ�%Ǽ�O¼|���ܵ����/������Ԫ�嫼��� ���괼D˹�ϛ��m%Ƽ2ͼ�Լ	�ܼ��弒���#�������	��2���&��`��(�q���0
��^��8������U���X��=����
����������K=���2��OH��+
�89�`� ��q�������x�TK�a���鼍�鼨��׻켁�����h<��v������>�����v�T[�c���"���$�2c$���!�7�N�����*���b�a��
��	���#�Y%��*�@�,��,��*���&�S"�~�����@�?������\��n�����o�����N�_=�����m���  �  .z=�=�g=�[�<J5�<�F�<���<�~�<:��<���</�<���<]��<�(=t�=? =�a�<�r�<���<w��<Z�<��<�%�<5��<G��<���<���<�t�<D={�=g	=��
=��=�=k�=�I=J�
=$�	=F$=�=R8=DZ�<à�<O�<q�<���<3�<���<�J�<���<���<�f�<��<�+�<���<��<���<�]�<r�<<4��<�ƣ<\��<�V�<���<��<~�<��<3�<��<���<~��<�q�<���<$��<���<v��<��<}S�<Ư�<��<��<CU�<�f�<��<l^}<��U<ق.<t�
<Z#�;EC�;7�;�0�;Ʉ�;`� <��<��<M�<-<=a�;>=�;��;�������"LA���T�-�6�)"�cY��:m;q�T;��~;<�;Rʈ;���;\f;��B;{1;jm�:�XT:x9�����h�sm�����W�컰V��<@�}6e��Ђ������W��<����[���I��H7z�a�i�ab�t�g���z�Ҍ�����O���^ƼK�Ӽ?�ڼ7�ۼ��ּ��ͼ�ü���ய��`��M����C��������������P���U������0`¼hsȼyOϼ~׼��Ἀ���C��W0�l|��4��b�O �|� �.��������
���=��e������
��Z�P��g���#�dN#�� ��;��m����������k��p�Ｍ'뼒���R���漌8缊'���D��:���z�����������&�����[&��+�9�.�ļ.�s�+���%�����3��>&�ҧ��N�~F��='���.�N:4���6�$x6��3�"�-�ڸ&� ���2������c ��Z���
��G
��f
���
�W�����\���3��&���  �  w�=�
=��=ex�<���<�
�<�I�<�q�<�1�<n��<~"�<� �<>��<���<c��<��<8)�<,�<���<�<Ն�<,�<�A�<� �<�Z�<���<*K�<���<K�=�=W�
=�=+�=��=LD=��=�>=xy
=�P	=Hk=�_=[��< �<��<�x�<z�<��<���<ɤ�<�<��<�<G˲<�<Q�<ȴ�<հ�<.�<���<���<rf�<F��<v�<S��<c�<�!�<�~�<w��<�`�<���<��<���<���<� �<+�<���<��<���<2q�<�W�<0�<�T�<��<_١<�f�<32t<~�E<��<X��;��;��_;��I;�2m;p�;��;V�;��<�Z<l��;~a�;'�];K�(:j���h������� ��
����*X��@˺��9���:uT;�Ʌ;SÒ;`�;�b�;\�r;w�K;F ;���:��:G�-9�M�s, �,,a�-b��+�����%�BLR��~�.$��v-���k��YB��-y��s=��������|�s�܋w��҅��������Av¼�ּd*��y��켘��r
ټ��ʼ����:��:���X⣼t���O��׈��������#���A��o��� Ƽ`�̼*ռG+�P��w��Ul	��y���_$���(���)���&��� �U���d�ٳ	����G���	��^�t��,e!�~=(��,��.,���(��"������5��2j ��P���\�'�輦0�sn�׎�@#�I�A�o����aM�as���n�}m�s	������$���-��K4���7��7�V�3��J-��_%�\���l��@�����"�3%��#.���6��<���?��)?���:���3�t\+���"�����V��3���
��i	��l	���	�OO
�`�
�a�������������  �  A=�	=��<5��<���<�S�<�a�<�<�=�<��<j��<��<�D�<��<��<2��<?F�<���<J-�<��<Em�<�Ν<w��<���<��<ڢ�<�9�<���<u9=�=�=͓=�=J�=�=0
=E�=	�
=T�	=a�=��=���<��<��<�5�<�p�<��<�y�<́�<��< �<m�<�ة<ʟ�<[�<��<=�<���<�>�<��<��<��<�3}<��|<���<I�<Z��<`_�<P��<�B�< j�<	�<��<���<��<=1�<p��<,�<��<P��<���<��<�X�<�1�<�M�<G;l<�9<��<^ͱ;ZS;��:�z�:��;�k;�.�; ��;���;�Y<���;<��;@S ;�u���T�ʗ�� �ػ��޻(�û�J����Q���q�:��K;�+�;K��;|��;.��;X�w;��N;8�";P��:Ў�:mx�9dE3�{�����`�s����� ���.���_������䜼P�������0���W������咐�����zD~�� ��苋��W������̼�|���o���ݑ��$）W��Ѽ:��dF���:��cp��𣡼��������^���~��J�������񢿼ż�˼'fԼ�;����I����1��!�/�)���.���/�J�,�{�%��/�;��q��|��б���$A�Ћ&�).�#12�>G2�.K.���&�>���L���	�4�H����켋���A�J���;��`����r1���_i�C ��G��0f	����ø�T�(���2�A:�5>���=���9��G2��)�6a!��m�h���d ���(���2�l<���B�!F�)E��G@�Ri8���.�3�$����Lf����2i�v�	����E	���	��
��
�΀�'��lK�]/����  �  ��=�	=�<]6�<��<(x�<�!�<���<\�<��<S�<JE�<���<���<8�<���<���<��<쵺<N�<�#�<9o�<)^�<��<�м<!K�<Q��<��<K=l=�/=�==��=�==��=M�
=�	=N�=ʻ=�L�<2��<���<�3�<U��<D{�<�u�<�.�<iH�<��<۹�<4��<3��<���<��<��<S��<֨�<<��<9l�<�<�|t<��s<$�<ⷐ<ˣ<->�<Iw�<�|�<�<N�<��<���<���<MD�<���<^'�<���<��<`�<z'�< N�<�Ѡ<�k�<�(i<�+5<�� <��;�2;��:Ua�:��:jDO;I�;u�;�r�;���;���;��;��
;9�d�{[r��O���E�
��s{ӻٙ��r�1�i\	����:T�F;B��;��;-Z�;!d�;^�x;u�O;�v#;���:��:��9+�-�B2���a�6������@F2���d�;�������T������c���*��B&S���D�����m��ǒ��B����ݶ�rmϼ|b�!D���������M��j��mӼ��¼�2��D����x��i{��Oբ��o���5��9\��������>r����ļei˼)PԼtm�TO���0�|���X#���+�1�p2�.�.�e�'����n���Ϳ	�L�	�Q��<P�����](��0�/]4��r4�&S0�ϼ(����?X��<
�H������ǹ켏p��弍�a��9�弫u�x��\鼒��5>�)��9����	��������4*�s4�*<��/@��?�$�;��
4��+���"�m}�I����H�!��M*�Pm4���=��E��PH��LG��<B��:��'0���%��s�Ȭ����[�.{	����1 	�v	��	
���
�Ol��v��0�������  �  A=�	=��<5��<���<�S�<�a�<�<�=�<��<j��<��<�D�<��<��<2��<?F�<���<J-�<��<Em�<�Ν<w��<���<��<ڢ�<�9�<���<u9=�=�=͓=�=J�=�=0
=E�=	�
=T�	=a�=��=���<��<��<�5�<�p�<��<�y�<ʁ�<��<��<m�<}ة<�<Q�<��<-�<���<�>�<���<��<��<|3}<��|<0��<�H�<۫�<�^�<���<�B�<j�<�	�< ��<���<V��<�5�<���<!�<���<��<���<w�<^j�<E�<0b�<Sfl<��9<!<$�;� T;�2�:}��:(u;��k;X�;y�;N��;r[<���;w��;� ;Re���T��ڰ�&"ٻ6�޻�-Ļ����%���d��1&�:��J;W�;t�;�s�;ۍ�;Ύw;�N;��";ɯ�:��:��9�1������`�c6��ѓ ��.���_��燼~Μ�:��e������pH�����-������>~�!�������^�����̼Č�2�ɤ��ǧ��!.�o�j0Ѽq���\���O��ۃ������k������yj��k���0���׬��৿��	żԡ˼hԼ�<���"J����1�!�!�F�)���.���/�U�,���%��4�>��s��~��ѱ���%A�Ћ&�*.�$12�>G2�.K.���&�>���L���	�4�H����켋���A�J���;��`����r1���_i�C ��G��0f	����ø�T�(���2�A:�5>���=���9��G2��)�6a!��m�h���d ���(���2�l<���B�!F�)E��G@�Ri8���.�3�$����Lf����2i�v�	����E	���	��
��
�΀�'��lK�]/����  �  w�=�
=��=ex�<���<�
�<�I�<�q�<�1�<n��<~"�<� �<>��<���<c��<��<8)�<,�<���<�<Ն�<,�<�A�<� �<�Z�<���<*K�<���<K�=�=W�
=�=+�=��=LD=��=�>=wy
=�P	=Hk=�_=[��<�<��<�x�<x�<��<���<Ĥ�<z�<���<��<<˲<�<�P�<���<���<�-�<d��<d��<"f�<䣒<��<���<fb�<� �<�}�<m��<�_�<���<���<s��<��<��<�"�<���<��<��<!��<�n�<�J�<us�<�5�<���<���<W�t<�TF<��<ӡ�;�"�;��`;Y�J;�#n;�I�;�[�;)L�;��<o^<���;�5�;�];��%:�����#����������`X���~Y�~�ͺ��9Z[�:��R;�C�;�N�;��;��;t{r;�{K;�A ;���:�́:w69q�J������!`�Dͬ�Q���.%�X�Q�Ⱥ}���������E��D ���[��%��髈�a�|���r�Čw�څ�����X��Ϗ¼�ּ�M���%9����7ټi%˼�<���e���ר���������3�����R&��z��i2��N���x���Ƽ��̼�ռ�-��Q�y���l	�9z�S��0_$�
�(�ҿ)���&�� �a���d�߳	����K���	��^�v��-e!�=(��,��.,���(��"������5��2j ��P���\�'�輦0�sn�׎�@#�I�A�o����aM�as���n�}m�s	������$���-��K4���7��7�V�3��J-��_%�\���l��@�����"�3%��#.���6��<���?��)?���:���3�t\+���"�����V��3���
��i	��l	���	�OO
�`�
�a�������������  �  .z=�=�g=�[�<J5�<�F�<���<�~�<:��<���</�<���<]��<�(=t�=? =�a�<�r�<���<w��<Z�<��<�%�<5��<G��<���<���<�t�<D={�=g	=��
=��=�=k�=�I=J�
=$�	=E$=�=R8=CZ�<���<O�<o�<���<0�<���<�J�<���<���<�f�<��<�+�<s��<��<t��<�]�<�q�<���<ŵ�<nƣ<���<�U�<���<�<*�<��<�1�<��<o��<���<"u�<���<��<t��<k�<:1�<an�<��<�4�<�A�<���<���<>R�<��}<7cV<q�.<�<��;�;���;�ں;��;�� <�<L�<*�<�<b#�;/ݛ;;�;׈�������B�3=V���8����i�gx:��;\�R;�R};�m�;|A�;
J�;^�e;��B;I+;���:�oV:{��_�T���k��%���������?�S�d�|���P���"��s��+2��y'��dz�Ԏi��Ob���g���z�D匼�5���s��x�Ƽ^�Ӽ�ۼ�ۼb�ּ�ͼ>Vü�и��민|����/���s���妼a䩼�ۭ�Sk���k���Ƽ��m¼�}ȼ�Vϼ;�׼u�����E���0��|�5�	c�� ��� �(.�������$�
���E��j������
��Z�R��i���#�eN#�� ��;��m����������k��p�Ｍ'뼒���R���漌8缊'���D��:���z�����������&�����[&��+�9�.�ļ.�s�+���%�����3��>&�ҧ��N�~F��='���.�N:4���6�$x6��3�"�-�ڸ&� ���2������c ��Z���
��G
��f
���
�W�����\���3��&���  �  ==�=�Y=�S =���<\��<���<-�<�I�<t��<K��<���<�=$=7�=M[=
� =���<j��<��<���<+��<� �<s�<@��<}I�<���<w��<��=e=�=H[=�	=�>
=�{
=E%
=�5	=F�=��= {=�� =@%�</��<f��<�Y�<���<x��<2W�<UC�<ȿ�<v�<8��<Y��<�,�<c��</��<_��<��<�3�<���<ө�<Ŀ�<�ͱ<��<gճ<��<���<9�<��<ח�<�-�<��<b�<��<C�<�~�<�5�<+R�<���<�\�<@��<b�<e��<Qq�<��<t؁<��d<�IF<�*<�\<7<�� <J<& <n�<��+<�h2<(~/<�V!<��<���;n�;DY;��:���=q�^�M��Kk�#v:���:��;��<;�^X;5�e;�'g;��];�<K;�4/;/�;�֯:q��93��fֺ�8�����N������{���.���J� �c�0Iv��X���ڙz��zm���^�lS�n�N�!U��Eg��j���R��}����H׿��ǼM`ɼ�rǼ��¼�g���*��	찼�A��$Z��e������0��&+��`���幼����5Ƽ�>ͼ�Լ��ܼ#�弪���%������	�A3�9��N&��`��(�����0
��^��8������c���X��A����
����½����L=���3��OH��+
�89�a� ��q�������x�TK�a���鼍�鼨��׻켁�����h<��v������>�����v�T[�c���"���$�2c$���!�7�N�����*���b�a��
��	���#�Y%��*�@�,��,��*���&�S"�~�����@�?������\��n�����o�����N�_=�����m���  �  �q=r�	=m=��=$�<"��<z�<P�<���<`��<c1=�L=^�	=�=�R=�o
=]�=,�=���<3v�<�o�<8x�<���<�L�<���<�D�<��<���<6y�<���<�*=�E=�+=��=�V==~�=�=�=�,�<���<S��<�J�<(��<��<��<*��<m�<Q�<J%�<D$�<k��<Ɂ�<pH�<l�<�W�<6&�<���<Q�</t�<���<���<ZT�<`��<vu�<�&�<b*�<���<��<T��<�<�<;��<W�<�Z�<���<�-�<Z��<���<�o�<�o�<�a�<�<�h�<S�<!�<��<	}l<B9X<�F<�7<�.<�*<��,<ߦ3<��<<aAD<�F<�B<��4<�<L8<E��;4�;��D;c��:�թ:%�:��:�Ԣ:���:h�:��;Ѯ;;�;K�";��$;��;Ҡ;Z��:��[:�V:�����0+��~������_ѻHl��8|�V�#��5�0�E��yQ��0X�2Y���T��DL�<C�~<���;��C�r�S�2�k�8X��#G��r�q��$Գ�YX�����E���0Ը�gg���$��T;�������n������+$��k��������7���ļ�g̼��Լ��ݼ7�p��\�����!���D�HT	�Ԗ�J���4�x%
����@M�(���^�� P�f𼘭���Z��������k��v�!���D������=	��c���s]������Z��� ��>�������� ��~���#��l#�hP������
�:L������=��J
�t���'���o��O�'i�e�	������	��(�����<�����s"��j#�E�"�)�!�uz��)��������b�(E�C:��X�Y������v������_��B��k��  �  �U=XT=��=^�=�_=6 =W=�)=�=_�=��	=c�=�=�b=�d=C�=��=�>=�0=V[ =�.�<v�<^e�<B��<)6�<�?�<��<���<���<N�<Y(�<&��<�d=
�=G=��=6U=�h =�g�<D��<\a�<�e�<���<7��<9��<��<)�<��<��<H��<���<kT�<���<s��<P��<��<�k�<�)�<�y�<�c�<$�<3h�<O��<��<w"�<_A�<��<�#�<��<;%�< o�<a��<`��<D��<k<�<���<&��<���<n��<���<��<?x�<�R�<AĊ<���<`�u<Y/j<϶`<cY<J+S<P�O<ӋN<-P<�S<ÆW<4Z<��X<w.R<LE<R2<F�<.	<w�;��;-��;�I;C�;#q�:c��:��t:'0: 	:/�:��>:[Q�:o�:>b�:���:�m:��8$w��Mv%��ۃ�.���&ݻ= �v������"��*���/�m�3���5��q5�x�2�)�.�~*�	�(�]u+��/4��FC���W���o��q��hZ��@뚼2ԣ����������D���Խ�V����4¼��¼%����j������<����C��m�ļ��˼�?ռQ�߼�i꼲������� ���'|��R�A��9��������V������u����0��g輝(�oV������W�����������	���	��G
��h
��'
��a	����M��g������������ ��j#���S��H����������%���!������.�nw��W�����M��:����	�L�� !�]�����l�R���������
����p���o�Aq����d�hC���L"����V�dy�����W��If����������� ��4$��  �  ��<�F�<�~�<�Q =�o=��= =�T	=Q�=��=�=P~=��=�=�}=@G=�+=�n==Y
=�=z�=v =+�<��<!�<���<T��<���<���<���<�x�<Q[�<]��<��<�� =6� =P��<���<���< ��<L��<���<���< ��<� �<j�<L�<�N�<�~�<}��<�x�<=P�<���<p+�<81 =.=�� =Zn�<��</�<1��<�"�<:+�< �<���<���<�J�<,/�<:R�<^x�<�1�<V��<4�<��<���<��<�_�<]6�<���<I��<_�<���<�7�<��s<�-f<<_<��\<)^<Ra< Qd<�Ug<{�i<��k<��l<��l<�Dk<�f<]^<,�Q<�A<�-<h�<�q<y��;�A�;���;tE;��:!5:����<���Ǻ�Ժo3���.f�^>��L�69�T�9��X��w�����q��0m���S��w/��0!�we*�O�-���,��I)��$��� ��"1�`����@��i����ݭ(�A�6��FH��Q\�J�q��u��_��ݑ�������]�����N&��^�ɼ>�ϼ��Ӽb�Լ��ҼACϼ*I˼¨ȼ��ȼrͼ�"ռ'm�w�f��������!	���	�d��/�����8�M@��k��a��
�3�D��Gv�z�Ἶ���伵��T�켌��R��-F���2�H\�f��%�����ۇ�Ba���̒������W��2���&��,~���z�-����
����a��y������~�m�
�����;������
�Up�<R��X�������}��X�+�D����	�`��9������e�����q!��O$�~C&�[�&��&�%�#� ���
4���=+���<�;��g$��M)�'-��  �  ���<�2�<���<���<� =��=�<	==�=�=�2=�=��=�=
�=��=Z�=�=�=,�=��=�'='�=i��<��<'�<��<8�<��< E�<EX�<���<n�<R1�<���<;�<yX�<e,�<=i�<���<!�<=�<B�<;�<���<N��<���<���<���<1��<��<m��<S�<�v =�=�=� =��=J/=X� =�S�<	��<�a�<�r�<Z��<���<���<���<�͸<\�<�_�<$�<�<z��<aú<�W�< ��<Iu�<-�<�;�<��<"��<X<@a<�L<�<A<0@<k�F<<�Q<ն^<��j<y�t<�Z{<{�~<q�~<K|<M/w<�p<{Qf<��Y<�AK<H�:<��(<�<dJ�;B�;��;̕G;�#�:�������!U����L���,u�GpB����Ӥ�K�k��w��[�
�I�q�rL��T �% ��9�҅H���M�w#J�B@�#|2��X$�t���N��Y�p���h�C�	���R��DT!��k.��=���N��\a���u���P�����5����潼�̼�MټF�⼛S��!���弾�߼�ټԼ��ҼX�ּL�߼��켓���"�S��]�	��'L�F���J�3c��q�����a)��뼨��F㼄i༔o޼|ݼ��ݼ�2߼g��w/�:��%���2����O���	���Q���������W��d���@	�K�����3��*��m���S%�E�	� �<D!��n�����L��d�%��M�	��\�>��"��)� �v����������?/ ����U�5���\�.�����ݪ��:��6 �p#&��Z+�j$/�C�0�{:0�&G-��(��##�7&�J��2������ �j%&���,�\�2�H7��  �  ��<���<��<�7�<���<F�=�P	=�~=(S=��=�_=�=�J=�!=��=��=c�=vO=�C=,a=+b
=�= ��<r��<m�<�P�<|�<�Y�<���<��<6�<��<{��<�a�<�@�<F��<M��<S�<�	�<���<���<؈�<嬧<U�<���<��<�a�<��<#/�<AD�<���<bW=��=��=$3=P=n=��=^�=o�=|L�<��<xr�<;��<��<��<�j�<�=�<���<�i�<���<��<�'�<�<).�<���<�[�<���<(é<{U�<�N�<��[<��9<�_#<:<x�<vo+<�7?<U<9Zi<őy< &�<���<6��<��<pW~<gRu<^�j<ܐ^<(Q<xzB<�2<�8<��<�;�$�;�,;j��9�h�󧃻����Ի��ٻ6�ǻ%Ф��%w��	0���
��?�|�X�3�����Û �7fE�ea�S#q�u�s��^j�<�X�<5B��d+�U��-������������f�����n�	x�U�)�(�7�W�F��W��k��聼Z<��R�������<Ǽ�1ڼ������BI��~�������B����n߼�ܼ�f�VO��w��%��Q��������^0����n!�=��հ	���������y�*����Ἡr޼��ܼ�~ۼP#ۼ�jۼ\Wܼ��ݼ�n�)D�M�s(���?������0��!��.%��Z%�[k"�,��X��S��
�˜�8k��t������{K"�N (��>+��4+�o,(�!�"�c�%��J<�(���6�C2�1�������x���A���s�������A���TD���ӭ�!K	�u+�Wg�@��r�#��#,��Z3��8��);�v�:�W�6��1��F*��$����=���� ���%��"-��&5�[d<���A��  �  ���<���<u�<��<�L�<L^ =�;=N�=W6=� =a�=w,=�=��=F1=�=�=br=�=�=�"=�=^�<"��<T��<�x�<-r�<�<8u�<ś�<	^�<�`�<h[�<b��<j��<��<���<���<�b�<��<6��<뙗<�ʕ<�}�<^��<�̷<=��<�y�<��<��<7��<E�==��=I�=��=ˬ=ZV=K�=/�=�� =���<���<2��<�U�<f��<��<���<�Ǎ<΄<�ւ<�ԇ<�F�<>h�<,ū<;��<Az�<���<���<1��<ֆj<�&=<��<���;U*�;��;�x<V�+<%�H<�fc<��x<��<��<V�<!�<���<E�w<ܧl<ت`<��S<�ZF<��6<R�#<�4<h�;���;5�;`�<��`��O���_��`���������]޻#ޫ�&��VO��.V�'֍�B�̻b���i<�oce����(\��y�����wp��XS�~�5�+�����{����컫ﻝ������z������'�I�4���B��TS�X�g������������^ܹ�!�м�6��x��%7���8���F�U���5�� �`h�P��a�o��.�vi������$�N(&�Z�#� ?��]�nx����������伄*߼VܼS�ڼ�ڼ�ڼ UڼM�ڼDܼ�޼���b���#�0
���%��x�*�-#��*�7.�IY.�V�*�8�$�����������֙�(�Ė��{!��*���0�yE4���3�k0��h)�� !�q���3�����c �����W��������Ŋ��G���+P���6 ����Wi��X�s���U�KC��"(�U2��:�� A�[*D�kC�?"?�E8�"Z0��")��7$��"�%���*��3�c=<���D�baJ��  �  ��<��<*��<�K�<m��<Q�<�=�/=MU=��=�!=�=m=L�=h==�==��=�	=��=�(=�b=AB�<<��<:��<;;�<|�<�ۙ<7$�<�ɚ<^��<M,�<���<a\�<��<\�<h��<$s�<�޸<��<�^�<6j�<���<D��<�t�<���<���<���<��<M��<�" ==ۘ=E(=�9=�=D�=ԟ=,=�B=�o=g�<4C�<��<n��<���<�"�<C��<|�<Bjq<X|m<��x</:�<��<y��<��<��<��<���<�6�<7�X<�{(<�� <l4�;X�;��;���;_S<a�><Jm]<�[v<z��<OՇ<xQ�<~�<Ю�<��x<�km<Nxa<�U<��G<7�8<�a%<ƥ<;��;���;K�:�pźmǒ�oQ��G�0'��(�.������Y̻E���.Z}�N���p���&��i�;1O��
{���*�����E���>�fz`�v>��c ��b	��������Á����/�����P�0J'���3�vA�^�Q���f��ր��������߾�iؼ��;��>D
�4����y�	����.���Ŧ��-�^�x~�����\w��v���$���*�TM,���)��K#�Il��k�ؕ�5����[�F޼�ۼ�ټ�xټ�ټ�ټ�aڼ�Aۼ�ݼ���nB�ho����u���I����(��/��04� w4�Ӭ0���)� � �Q�=��]���m�T�:[���%�*`/���6��k:�::�L�5�-#.�?�$�q���S��v	�f���_��U���n���_��+�����WK��Я��g���pZ����y.�SL�?s��Z ��R+�BM6���?��G�ORJ� tI�T�D��!=�+q4���,��)'��y%�'�'�{-.��7��A�J�|`P��  �  	@�:��;"ܛ;�G
<��Q<�=�<:��<���<���<\��<���<,	�<�L�<j��<���<��<6�<���<���<D��<9P�<�F�<"��<�`<G<���;�U*:H�亏��D���ӱ:�p�;�<��E<S�f<�Ck<��R<��!<���;[��:����,h���~�r ��*:1�;�<s�]<e�<�ũ<�v�<��<|��<�}�<���<&��<�v�<�<�<���<f�<I��<o!�<�~�<m�<��Z<�<��;n���d�Rذ��ƶ�K���B���$;�l�;��<��<�<�!�;ݘ:Ѧl�����D�"Ri�@�o��PX�Z)���ֻ�!�~�:<�;�|�;H�<W<��#< !!<�<��<>�<Z��;Vf�;$��;��!;��=��$W����C��銼v����ּ������ ���mu켆�Ӽ���df��o0���A���@������s|Ӽ�����0����7� �9!�.�������r�μ���������S����q���f���d��i�y�q��E}��q��
�����������HƵ�aJ̼*���[���.�'�B���S�+g_�`d�h�a���X��JL�k�>��4��4.�	:/��b7�wE�	W���h��x������΁��/~��Hr�o�a��vO�V2=�$�,���w��x��h'
����$I�y�����hs�����j
�^��޲�z����,�{U=���O�.c�w�t�~��J�������";��E�u�b f�^�V���J���D��F��ZN��&\�[�l���|������͇�)S��.K��T�x��g��"U���C�`�4���(��W �(��_��z���q�,���W�<��m���]�G�"�l/+�ؚ6�aE�
W�gcj��}��$��`���Ï�޸���D���b���w��h�~�^��A[��&_�s�i���x��c���z���  �  ��;�P;���;�<*�Y<��<�3�<u�<۔�<_��<��<bE�<X��<��<MU�<~��<xS�<��<���<a?�<�B�<!��<y�<�f<��<�>�;��:�a_��Rƺ�WṠ�;9�;�<H�M<S�m<2r< HZ<��*<���;_�/;�"�'-�,aC���Ϻ�P�:�;J<�b<u��<��<D�<D[�<���<���<�7�<��<���<���<��<���<� �< ��<���<M%�<�6_<�<�>�;՞:w�-��^���Q��":S�Ju��0<;���;n[
<+|<L	<�N�;�F�:}hA������6�R�Z�za�~K�C��?Ż�����:,�;o?�;�w<F�<U$"<Ш<XK<4�<w� <*X�;1��;'׌;Z�;�\��8�R���=(>�V↼� ��c}м.��9��T�����)�ͼG����/��(���f懼Ĺ��槬�:�μ��q�
��R���֕�_��-�e��p�˼�2��������� "s�9Lh�2f�Ujj�r�r��C~�����O%���@���9���,���7̼1輵�W���,��@�~P�U�[�J`���]���U��mI���<���1��i,�2|-��|5��>C�(gT�m�e���t���}�T����z�35o�ym_���M��<�pH,�%g���|���
����9����$�;���/��
��,����ɇ��b,��><�(4N�ѭ`�̏q�u�~��؂��悽
�~�&�r�@tc���T�d�H��C��ED��cL���Y���i�Ȕy�J؂�
����|��A���x�u��Ke��S��B�j44���(�ԕ ��%����%K������ܢ�l���,����xB#�VN+�^d6���D�e�U�?lh���z������Q��z卽`䌽���m恽t��f���\�~�Y��Z]�w�g�hzv��y�����/���  �  �;�׸;^��;/�2<�o<�<S˳<6��<�\�<��<]�<���<�C�<��<�i�<bi�<9��<�c�<��<��<�f�<N�<�̚<=�u<��2<S�;�Et;���:�^�:1;#P�;�;�5<��d<Mƀ<̂< �o<��C<V=
<��;���:K�ĸ���	�Q:�m\;"�;Ӣ/<qKn<	�<g�<�n�<?��<��<*�<���<�#�<��<�b�<+8�<z��<�d�<�<`�<�S�<�j<��)<�R�;D�*;�>��c�Z���QZ����:���;Z��;|T<�d+<
q<���;�W;օ���j��'_�31��k8���%�:[�����Q�����;���;v�;� <�<@�<��<<<��	<���;��;���;���;P�;�BY��^M��ڻ_0��Qx�蜟� ���Y}ռ!���߼�pҼ�＼�?���A���Y����|�q������9�����㼁���-�d��.���
�����b��+�ļ����0`��b҅�D�w�Էm��dk�:�n���v��܀�
ׇ�@S������	���B	����̼6��y��?��&��A8�B!G�&aQ�S�U�o�S��:L��UA���5��;,��V'���(�50�e�<�z�L�F+]�_�j�cVs��ku���p�Ĵf���X���H��9�.�*�Qe����/�����<	�%��(������	u	��-�(w��������D+�׀9�'�I��Z�@i�y�t�>I{�V{�u���i�)�[��%N��~C�=(>�YP?���F�C4S�tb��zp�o�{������V��M�y���m�b*_� ZO��X@�f3�K#)��!��z��G�7�����m�����3�i~���Vv$�[�+��%6�"C�	dR�"'c���s��$��2T�� ���+����Ƀ��]{� fm��`���W� �T��>X�P�a�/uo�p�~�6�����  �  <<c�<��1<�U[<�R�<X��<c�<έ�<�X�<�<+~�<�!�<���<���<k��< 2�<7��<h��<=�<���<`��<��<��<xʄ<�4R<]p<f��;v��;{ �;���;��;��,<�\]<�@�<{��<�^�<u��<��h<՚6<��<�
�;��o;hW;���;���;�<�H<~{<W��<h��<ƶ<f�<D�<���<.y�<(�<���<&��<t�<&�<��<���<���<�L�<��u<|DA<k<+�;�%H;�M�:50�:B1;9��;	��;�!<ܜ><3�G<	9<n<b��;�R�:_T�ލ��������Ӕớ����Q(��9#9�%4;肢;RP�;$z <�<�<H�<W�<�Q<��;o��;��;u]X;���:1�4��FW��uϻ� ��+\�ȗ��2y��i}���¼�����󵼕ϣ��􎼙�x��'b�0(`��lu��܏��C��=2˼�r�j��b��U@����8�鼺yӼR�����������≼`i��;Uy�qv�nx�	`~��r�������֔��ߟ����r༼%�ϼM���u ��-�(���K-���9�okB��!F���D�6e>�G5�j�+��#����W(!�4(�ɔ3�2�A�D'P��:\�*�c�)f�l�b�;�Z�raO�B�t�5�,4*�*� �\���
�%��Y����	�q	�Q	�
�O	�G��[�r8�@� ��*�6�6���C��4Q�#�]�}g�G#l�6�k��pf���\�БP�M�D�o;���6���7��|>�WI��VV���b��l���q���q�~Xl�~�b�L�V��J���=�	W3�P�*�;/$�Oh����s��r����eq��1�%"��B'��.���6�(�A��vN��>\���i�7�u��@~��������]y���n���b�-�W��P��rM���P���X���d��Mr��^~�;v���  �  �U<�+X<�{i<�ӂ<oܓ<��<�&�<���<�L�<8��<�*�<���</��<J�<���<�<6��<L6�<���<���<kf�<n�<���<�\�<C�p<��J<i7,<�_<�<�[#<�u?<`+e<J|�<@L�<wn�<L��<r�<Wb�<�k<h�?<Q�<%�<-��;�<�<�X:<�u^<�N�<���<=��<��<���<E4�<��<���<�n�<lM�<�<N�<��<z��<R�<a �<w��<,,{<W$U<�U.< �
<c�;�K�;���;Q��;.�<��-<��M<k�c<�i<��Z<:�9<#�	<*��;�_�:6)���Z9���j�Y�iv���)�@�:�'<;��;�|�;Dt�;6y�;"��;���;���;I��;�n�;^{�;Gu;�	;:��9�躺H����ӻ�&�^,B�\�m������$����o�������/��h�k�?�N�/
>��f>��R�-w���������)�Ƽ��ټ�A��0��`�y�Լ:Ƽ�涼T���ϓ��x����Ћ��冼�)������ą�����S������⨼��Ƽ��׼��꼖����+�M��C�!��
+��}1��84�6�2�� .�%'�"{�{�X���f�����z(�ܐ4���@��0K��R���T�3S�I�M�F��=��3�J�+��$�M���K�h���D����d��g�����a�����t'�[�$��[,��5�}�>�lJH��Q�Y�W���Z��&Z�HRU��*M�]6C�Ir9���1�i,.�/���4���=��}H��S��`[�'`���`�}]��W�w�N���E��H=��5���.��B)�~�$��� �9�����!����Y�@�"��,'��,�M�2��:�ozB�5�K���U��_�`2h�n��_p���n��h���_�vV��M�y�F�X�D�x�G���N���X�b�c�G�m��Iu��  �  rJ�<�
�<���< ړ< �<n'�<gt�<"ҷ<J�<{��<bT�<F��<���<F��<��<!��<�}�<���< ��<ü<9ڰ<��<�i�<#Ӎ<���<�p<f"a<�NY<)�[<T9i<D^�<�Y�<�ٞ<�Ϋ<���<f?�<$��<��<xU�<)�}<:E_<+iI<0~><	v><8vG<D�V<�i<Ý|<�F�<'X�<���<��<��<�ݹ<
��<�g�<�U�<�o�<,S�<=��<�`�<_^�<=c�<�}�<�/s<�_]<�1H<5f5<ݳ'<��!<��%<,�3<��I<�&c<�Mz<���<�u�<=}<D`<��7<�d	<���;a�N;�߲:ɠ9`y�ޥ9��-:+�:�j;�A;�:t;'`�;r�;���;Vx�;���;��;U��;;�x;-�
;��q9R�byr��d��z����b�2��M�2c�9�r���x�E0t��e�C
P��8���#�h.�!� �-�oM��Vv��b���8����\Y¼m�Ǽ��Ǽ�:ļ�U��!���o���J����
��9���W����ڑ��6��/���w����P��/������hƼ�ּ[��3?�����},
�=e���`��6R!�n�"��L!�Z���y�� ���@��or������'��21��:��q@�x�C��kD���B���>�&Z:�gi5��T0��*+��%�9� �Qp�5��U��d�n_��K����K��^� �	u&��,��1�Q7�|<�h�A��;F��UI��GJ�̐H��D�\n=���5�"�-�r$(��R%�(&���*���1�WY:�]�B�o�I���N�Q�P��O��4M��AI�ָD�E@��B;��z6���1�X�,�9D(��u$�b�!�:!��,"��&%�ݘ)�r /���4���:���@�E�F�ˇL�KR�"�W�"\�g�^��F_�!�\�w�W���P��0I�=?B��=��<�wW>��C���K�F�T�:8]���c��  �  @x�<*У<���<��<�՛<) �<���<�Y�<uy�<+2�<���<�2�<���< ��<��<�g�<��<�h�<�]�<Tۤ<�T�<��<Xa�<H��<h�<'��<�$�<��<|��<nb�<}��<�q�<N�<g��<v�<!O�<�/�<<t�<���<��<&�<C�<�v<r�k<p�e<M�b<eYb<��d<�k<Ȗw<1��<C��<�(�<�#�<.��<���<��<���<�<�y�<�S�<Y?�<2�p<��b<$�Y<WHT<�Q<!Q<��R<BX<��a<S�o<��<gƉ<Pk�<���<�ϔ<g�<K��<��a<J&;<"�<�`�;+&�;�c;<�;#��:h�z:�: ��9d�9��Z:m�:�� ;;�`;cQ�;���;���;�c;9��:�T������_����ֻsv��"��!*�>�4�3<�,�@�?�A���>��m6�Ԇ)��|��J	������L����z$���'��KI�)n�� ���ژ�����y��u����w��0뾼i���x@���Q��躼�8��G.��G]��V���R��L����ԩ�z跼�Eɼ�ۼ��p�����	�#��E5��<�֜��!�͋�������?���X���'�wC�.��Ǵ�����#��*�Q1�s�5�� 9�S�:��;���;�G;�8�9��i6�f�1�,,��%�������S�b	����É�8�%��a,�6y2��n7��;�gZ=�٦>�`6?��'?�Y>��<��[9�~�4��>/��&)��|#��>��A�����\!���&��-��e4�F�:���?�	MC���E��G��G���G��$G��NE��$B�ɟ=��8��&2���,�f)���'�$)�+�,���2�_�9�g�@���F�ڹK��AO�ƏQ���R�B�S�"�S���R���P� �M�[�H�9CC��o=�Y\8�b 5��4���5�AB:�qh@�ikG�:QN�2ST��  �  8��<�<�7�<���<�(�<���<��<`�<E��<���<��<�W�<ɴ�<�5�<#��<?�<��<���<��<^��<<>u<Q�g<[4e<�l<#�y<�]�<2��<��<ڪ�<6V�<' �<	��<�G�</��<(��<r��<��<�X�<���<���<4�<|z�<�<҃<ARq<e�[<�H<^;<�6<%P;<��K<h�e<��<V��<i�<5��<pŦ<��<���<Ic�<�qc<�&G<��3<��+<`�-<W�8<T;H<�3Z<�ol<~<;v�<�<!��< p�<��<ے�<�X�<�Ě<L�<��<�vc<��@<WR<��;Է;�[q;���:�k�8_���Ո$�AH��BA���y�����9���:ī";J ;;��:�M��.O5����g���(�=�@���M�ٖO�`XI��>���0���"�������Xo�8�ڻƻ�9���7��}9ƻd{���w�$���C�'�c��������Vӟ��>�� ����ȼ�Ӽƈڼ��ܼ5�ټ��Ѽ_�Ƽ����B���vS�����X��/&˼�:������L�����v��v�x����I%��1��W����V��u �=!���R���d���} �����"
���ի�����g%��+���1��7�&y=��BB�^�E�#�F�%sE��7A�:���2��w*�V�#��; �� �/�#�f*�I2�2�:���A���F��H��%H��|E��rA��<��7��2�<�-���(���#�S������'���>��������#���(�J�.��t4��=:�E @���E�)K�ȪO�k�R�zlS�asQ���L�f�E�L<>�F 7�\�1��/��I1��\6�|>���F�q]O��6V�ًZ�\��#[��GX�tGT���O��!K��sF�j�A�?�<�T38���3��90���-�-�K�.�F2��6�u<��pB��rH��  �  ���<lG�<q"�<��<���<G�`<VK<��D<�(O<7�h<br�<�@�<ᡫ<Mض<@]�<�m�<�9�<���<�p<��I<:�.<#�#<W�(<1�<<FhZ<@}<[�<Pܠ</Y�<#��<<��<G?�<E��<cl�<r��<|l�<�g�<���<Q`�<���<ᾶ<���<�P�<�߈<@�k<��D<�n <AH<���;jp�;L<��%<HM<��u<�h�<:Ɣ<���<���<��v<0�M<��#<��<@�;]��;�d�;Q�<�g.<��Q<Ht<�O�<Rܕ<��<���<�ϫ<,�<|ڭ<���<��<k��<Ƌ�</f�<��`<��=<ǒ<�B�;-�;k��:�X庉~���ʻB�컐��u�ѻ�C����7�@2����%9%�9�8��8�y�������RE�X(m����?��W~��хm�[�P��2����Bw����λ�)��Mq���p��bn���O���8��~����h�j	��$���B�nd������瘼����*ż	�ڼ�����js���������E�k�ӼqTƼB�����{�̼9X�����
���K���#��2$��!��H�@���(���W�����X���I��H�-��2�������������7	�!e��8���'&��g/�.K9�z@C��VL��[S��(W�C�V�[�R�ՙJ���@�I6�v�-��()�(�(��w-���5��@��|J�ZS��)X�p6Y��BV�7P���G�¦>�d�5�%�-��w&� ������lw��q�ݥ�X8��#�>��]�=k ��g&��i-�|�5�Q�>�9�H��gR��[�Zpa��Ld��c�t�]��hU�X�K��'B�3O;��{8��_:�G�@��NJ�vZU��_�\�g�M�k�"�k��.h��~a�!Y��FP���G��N@�'�9�\�4�M(0���,��(*�ػ(�4�(���)��P,���/�H�4�:��~@��  �  ��<���<�ˡ<��<2V<�l(<�i	<_�;��<c'<iS<��<
�<�ߤ<,�<��<�؍<�=j<_B5<�<��;_�;���;*�<[�2<�d<b��<_��<�ڵ<��<�Z�<�r�<���<|+�<��<N�<���</h�<<$�<ex�<���<���<d�</�<)�Y<<e#<�,�;&��;��B;�/8;��;���;�\<�G<6�o<�D�<4��<|qq<��I<G�<���;]t;2�;��;�_;X�;V&<�><��n<��<�1�<0@�<a�<�7�<�D�< ��<]��<�8�<1��<�ޖ<��<��t<�"P<
w$<���;�^;J'Ĺ�K������$���<��,?���,��,�SĻVp� �
���躢�:����L9��$K������9���ɥ�S������*ڌ��n��@�d+�c��)!��V熻��a�^�O���R��h��������Ļ���F��^�.��[S���~� Ҙ�#U���bӼx������#q����	�Up ��%���ڼ��м5�Ѽaj޼s ���4	����lx&��Q0���4��3�Y4.��%��/��N�ަ��������'�z��\��˅�{����６��������>��
�"�֯�P$� 00�J�=��xK��?X��Qb��%h�P�h���c�DeZ��>N���A�q�7��1�V�1��7�^A��M�{Z�23d���i�)bj�܊e��f\��{P��|C���6���+�*�"�b���L�z���'�����S���U� ��P��'���!���)��^4�ʰ@��DN��[�-h�C>q�8�u�$�t���n�ϐd�Z�X�M�p�D�;A��DC���J�TV���c��o�1:y��}�G�|��v���l���`���S�&�G���=���5��d/���*�]�'�u&�6%�ZK%�S&�8M(�xB+��Z/���4�0	<��  �  {�<xP�<��<�un<�,<���;Ý;@)�;?~�;*t�;2"<�Z<���<��<{��<�w�<��w<�!?<V�<���;�G+;+� ;%>;��;��<n�I<��<�E�<ɔ�<-_�<���<iK�<AA�<Z��<���<U��<��<�q�<Q��<�O�<���<���<�<��<�XD<��<��;�7�:_75�(\z��Ϸ92	B;ݿ�;w <�N<�h<q�i<��P<�5#<A��;oA;h�	9�����_��7}56;���;
�&<e	c<�u�<Ű�<��<N��<L��<���<���<��<s��<���<<��<jR�<_�<߀X<6�'<�Y�;�%;�J�O�ӻ��+�� ^��Uz���|�n!g��>��L������>���h����`�ﻕe5�'�z�������\ļ�eļ����6 ��Sd����R�~��;8�,z��xc��J3�9�#�y�,�d�G�@�p����������ٻ���$�@L��k}��m��Y��b��� ��--�b� �
,�t�����~Y ����z�߼�߼D��l^�߼��%�q�4�/Y?�6 D�VB��d:�?�.�� ����`�����e�@8�v��3k�۸�k�漶���(�#����T�@�[���=-$�ɮ2��B�3�S�yc���o�� w�0x���r���g���Y��K���?��G9��9��2?�E�J��X��Ug���r�']y��|y�2Os�E�g�<Y��6I���9��-,��>!�p��d���������]�w��Q��#�6g�^M��R�U�(�^D5�?%D�^�T�s\e��Ht�hd�-~�����~#}�smq��}c��BV���L��_H���J��]S��}`� �o���}�"�����������ف��Xw��Kh���X��I�Z{=��3�Z�,�(��#%�d�#�U#��Y#�!C$���%�h�(�k,�_2��:��  �  .�<���<���<zX<��<n�;z�;��:�;v0�;,<f4><f�s<k��<�<m�<T_<#7"<�3�;��;���8,����9''J;��;�*5<�/{<�4�<8�<,��<�n�<��<(��<��<ʎ�<%��<�<���<Ց�<���<���<�B�<AH�<�cz<w'3<	��;@r;�&�R���f��`	�o�E:o]�;FA<��8<�3U<h-V<;<�|	<�n�;�J:Q��!A�����O�ןG:���;+~<S-X<<�<�ޟ<���<��<��<<E�<ه�<�µ<~s�<���<��<ӑ<��<lI[<QO'<���;:�:��Q�O��`N�����Q=��Tn��E'����a���+��l��^�����{�����aP��e��<p��W8˼UBټ��ؼ�Fʼ�<���𑼟b�%�?��M���~�Q����q���P��.8��Db�\犻ʩ�.�ϻ�h ��f ��)J�\z��R��E�ż¦�E*
�����M&��a+�6h)��.!����0=��J����鼆t�G����H	���!u-�7�=���I�T[N�<�K�gC���5���%��$�/��E��Y�꼳���ݼL�ݼ�S�$��c��n��r������ҷ��{�����%�F5��@G��Z��|k��Ly�/����L��S�|�P�p��a��"R��vE�G7>�i�=� �D��Q� �`��=p�|�|��끽-��|�--p�X�_��M�fc<��6-�y!�m$�5��Z�DU�{��d��������~�������(�#�6�0G�T�Y�:l���|�s�������OH��Op��\z���j�qo\���Q�p<M�c�O��Y�?Ng���w�K���9���̋��͊�s����
n��u\�� L��>�G3��+�f�&���#��n"��"�nd"�f=#�|�$�w*'��+��0�υ9��  �  ��<,��<�׎<�O<��<�U�;ڎ�:�,�9+�:�Bq;*�;g4<2�k<���<N��<�d�<��V<o<I:�;M�:�U��kź��ιߪ;!�;nt-<�!v<�ߛ<�ֶ<:�<l�<���<���<���<�#�<+n�<ܻ�<8��<�X�< ��<�^�<5�<�h�<�qv<k�,<| �;���:]���Æ��"��%B��[̷f�v;��;��0<�@N<�EO<�r3<�l <0Ӏ;e�6��N����4���O���7"d�;��<W�S<�2�<V��<��<4��<�ѽ<.�<m�<�>�<��<>�<<e��<̦�<b�[<̥&<"��;_|�:}�o�+����Z�<�\����Қ����t�m��E6��f��+���N����λ��	�Y���������dҼ���K�߼h�мmѶ��A���h���(�ҕ��n��ۜM��I�?��e�ح3�!%^�ﱈ�[4���ͻ�����P���I�TR��顼��ȼ������ ����)�/��-�8{$�����	��U���/�7���I��:`�TR�hi0��XA��2M�9R��lO��)F�))8���'��g����1����꼽�/�ܼc�ܼ�߼� �lI�]EＡC���
��tY�>�6��t%��6���H��V\�\en�J�|����*)������	t��cd�JqT��hG���?���?�l�F�>JS��Jc��as�},���ǃ��ȃ�x-��(s�vb�)nO�8q=���-�#!�������{������)�W�W�����w����ø��[��)�\<7�qaH��w[�Ƚn���o_��p���h ���(��}��um�|�^�b�S���N�ߒQ�C[�E�i��z��,�����Z����������8怽�Ap���]���L��e>��;3��Y+�@H&�(g#�"�R�!��"��"�.a$�@�&�D�*���0�hr9��  �  .�<���<���<zX<��<n�;z�;��:�;v0�;,<f4><f�s<k��<�<m�<T_<#7"<�3�;��;���8-����9''J;��;�*5<�/{<�4�<8�<,��<�n�<��<(��<��<ʎ�<%��<�<���<Ց�<���<���<�B�<AH�<�cz<u'3<��;5r;�9�R���f��`	�ǣE:T]�;5A<~�8<�3U<B-V<�;<�|	<Yn�;ʻJ:S��dB��U���hS���G:�;�|<�+X<n;�<�ޟ<X��<���<2 �<I�<4��<ʵ<�|�<f��<��<R�<{�<ts[<�}'<��;n��:��P��n�5+N�'ǂ��%���X��a����a���+��I��J����������s��#vP��s�������L˼0YټS�ؼ�`ʼdW�����ELb�FF%�I0������AR�Jm���K���O8�yGb��ي�6�����ϻ�K �C �D J��K��9����żR��
�9��A&��U+�v])��%!���Y7��B������t鼢���M	�*��}-��>���I��gN���K�gC�֤5���%�3��<��^����꼖�Ἂ�ݼ?�ݼ#a�j�伔�����'������e��}�o��=%��5��@G��Z��|k��Ly�7����L��]�|�X�p��a��"R��vE�I7>�k�=�"�D��Q�!�`��=p�|�|��끽-��|�--p�X�_��M�fc<��6-�y!�m$�5��Z�DU�{��d��������~�������(�#�6�0G�T�Y�:l���|�s�������OH��Op��\z���j�qo\���Q�p<M�c�O��Y�?Ng���w�K���9���̋��͊�s����
n��u\�� L��>�G3��+�f�&���#��n"��"�nd"�f=#�|�$�w*'��+��0�υ9��  �  {�<xP�<��<�un<�,<���;Ý;@)�;?~�;*t�;2"<�Z<���<��<{��<�w�<��w<�!?<V�<���;�G+;+� ;%>;��;��<n�I<��<�E�<ɔ�<-_�<���<iK�<AA�<Z��<���<U��<��<�q�<Q��<�O�<���<���<�<��<�XD<��<��;h7�:�75��\z��ͷ9�B;���;�v <լN<��h<)�i<v�P< 5#<��;
lA;��	9d����������7k,6;$��;�&<wc<�t�<n��<��<⎶<��<�<��<�%�<Cӭ<ƥ<�ϛ<�q�<��<=�X<�J(<��;ɭ&;LZ����һ�`+�&�]�L�y���|���f��>���4���B��ch�5�����Q�5���z��'��-����ļ��ļ1��4��E���ES��>�,�໻���5d��04�T�$��`-�4(H���p��e��&m��~�ٻ=Q�fb$��K��}��<��~%��-�����X�T� �N������9N �����߼��߼���f����g+%��4��n?�D�.B��:��.��� ���p���2���켸`�,������@�漀���6�*����X�J�z��v�%.$�^�2�j�B�}�S�<yc��o�� w�Kx���r���g���Y��K���?��G9��9��2?�G�J��X��Ug���r�(]y��|y�2Os�F�g�<Y��6I���9��-,��>!�p��d���������]�w��Q��#�6g�^M��R�U�(�^D5�?%D�^�T�s\e��Ht�hd�-~�����~#}�smq��}c��BV���L��_H���J��]S��}`� �o���}�"�����������ف��Xw��Kh���X��I�Z{=��3�Z�,�(��#%�d�#�U#��Y#�!C$���%�h�(�k,�_2��:��  �  ��<���<�ˡ<��<2V<�l(<�i	<_�;��<c'<iS<��<
�<�ߤ<,�<��<�؍<�=j<_B5<�<��;_�;���;*�<[�2<�d<b��<_��<�ڵ<��<�Z�<�r�<���<|+�<��<N�<���</h�<;$�<dx�<���<���<
d�</�<%�Y<6e#<�,�;��;o�B;n/8;��;w��;�\<֋G<��o<�D�<��<�pq<�I<o�<~��;�Wt;^�;f�;{_;��;�"<u><��n<���<d1�<oA�<��<�>�<�N�<���<��<!R�<���<��<��<�Zu<+�P<��$<P��;�a;�ⱹK&��q���r$��D<���>���,���
�{�û��o��.
����//;��g���r�rK�䂼q��/���^���C��]#����n���@����O��^��­��,c�s�P��zS��bh�b���须�jĻ�n��f�ܝ.�1�R�7O~�Ռ��7��Ӽ-�E���^��P����I�	�~[ ��켪�ڼ�м��ѼFv޼[7��ME	�v��Ȓ&�p0�\
5�|4��Z.��/%��V�u����0��s,�A�<��M"���}	�𼮷��B����D��
��ױ��$��00��=��xK�@X�6Rb�&h�v�h���c�ZeZ��>N���A�{�7��1�[�1��7�aA��M�}Z�33d���i�*bj�܊e��f\��{P��|C���6���+�*�"�b���L�z���'�����S���U� ��P��'���!���)��^4�ʰ@��DN��[�-h�C>q�8�u�$�t���n�ϐd�Z�X�M�p�D�;A��DC���J�TV���c��o�1:y��}�G�|��v���l���`���S�&�G���=���5��d/���*�]�'�u&�6%�ZK%�S&�8M(�xB+��Z/���4�0	<��  �  ���<lG�<q"�<��<���<G�`<VK<��D<�(O<7�h<br�<�@�<ᡫ<Mض<@]�<�m�<�9�<���<�p<��I<:�.<#�#<W�(<1�<<FhZ<@}<[�<Pܠ</Y�<#��<;��<G?�<E��<cl�<r��<|l�<�g�<���<P`�<���<ྶ<���<�P�<�߈<:�k<��D<�n <5H<���;@p�;�K<l�%<�GM<��u<�h�<	Ɣ<���<u��<�v<)�M<��#<��<�;4��;D^�;{�<gc.<�Q<rCt<N�<�ە<���<���<�׫<�8�<w�<ç�<7�</��<���<M��<"|a<�><K.<���;AH�;$�:P�ߺ)����Ȼf�뻭��ֱл�p��~z6��]���/.9���9]$:�jF9�.��"^��E��m� ����l��oՁ��8n�:�Q���2�0��"����л���:;�����%ى�쇏��=��jj��G��	��C$�ՅB�C�c�pW������HZ��T�ļ"Uڼ���V����#��~���˼�Y�㼋�Ӽe:Ƽc5������̼7t�����5
��.�j�]�#�I_$�;7!��x�p��H�l�������#���K��~�'��g������4�����>	�Yj�a<�����(&��h/��K9�	AC�WL�?\S��(W�s�V���R��J��@� I6���-��()�/�(�x-���5��@��|J�[S��)X�q6Y��BV�8P���G�¦>�d�5�%�-��w&� ������lw��q�ݥ�X8��#�>��]�=k ��g&��i-�|�5�Q�>�9�H��gR��[�Zpa��Ld��c�t�]��hU�X�K��'B�3O;��{8��_:�G�@��NJ�vZU��_�\�g�M�k�"�k��.h��~a�!Y��FP���G��N@�'�9�\�4�M(0���,��(*�ػ(�4�(���)��P,���/�H�4�:��~@��  �  8��<�<�7�<���<�(�<���<��<`�<E��<���<��<�W�<ɴ�<�5�<#��<?�<��<���<��<^��<<>u<Q�g<Z4e<�l<#�y<�]�<2��<��<ڪ�<6V�<' �<	��<�G�</��<'��<r��<��<�X�<���<���<3�<zz�<�<҃<:Rq<]�[<��H<�];<�6<P;<o�K<A�e<���<6��<�h�<���<*Ŧ<���<"��<�b�<Npc<%G<��3<��+<��-<%}8<�6H<�.Z<7kl<�~<�u�<߀�<�<y�<,�<���<�s�<��<�2�<�+�<n�c<ɆA<B�<�y�;H�;�ft;���:�9�w��7�!���E�D�>�CR��Jx�l]�9ɾ�:�>#;�! ;���:8�����6�}����Ǫ(��pA��PN��XP� J�5�>�1U1��?#�pH�Z������-~ۻ;�ƻ!����v���>ƻZF仾t�2$�tC�ac��V������t���ڭ�ι��Y�ȼ�Ӽ`)ڼ=qܼ�oټ-�ѼʇƼWк�Xy��^E�����Dh��FE˼Th�.����������0�F��������nO��Y��d�]��u���&� �%^������ȏ��� �t���-
� �����Ү�Xj%���+�2���7��y=�UCB���E�m�F�]sE��7A��:���2��w*�d�#��; �� �5�#�j*�I2�4�:���A�F��H��%H��|E��rA��<��7��2�<�-���(���#�S������'���>��������#���(�J�.��t4��=:�E @���E�)K�ȪO�k�R�zlS�asQ���L�f�E�L<>�F 7�\�1��/��I1��\6�|>���F�q]O��6V�ًZ�\��#[��GX�tGT���O��!K��sF�j�A�?�<�T38���3��90���-�-�K�.�F2��6�u<��pB��rH��  �  @x�<*У<���<��<�՛<) �<���<�Y�<uy�<+2�<���<�2�<���< ��<��<�g�<��<�h�<�]�<Tۤ<�T�<��<Xa�<H��<h�<'��<�$�<��<|��<nb�<}��<�q�<N�<g��<v�<!O�<�/�<<t�<���<��<$�<C�<�v<m�k<i�e<D�b<ZYb<��d<	�k<��w<!��<.��<�(�<�#�<��<���<���</��<��<.y�<S�<j>�<��p<�b<��Y<DT<4�Q<Q<�R<�>X<W�a<I�o<D��<�ω<�y�<���<��<�:�<�ށ<y/b<3�;<�q<���;䎣;��f;�;3W�:�ă:r: M�9V��9�.e:G��:�";Db;&׊;Y�;���;z}c;� �:ѐ͸�;�Qj��K.ػ`%������*���5���<��rA��B�	O?��7�x*����.�	�P����ﻋ������i'�u�H�X�m�t���B����]�����/����1������������������������0����������X���;婼q��ttɼ�!ܼ������&?�2
����l�Kt�U��3V�?���������d����O��>��U����������#�U�*�M1���5�-9�S�:���;�T�;��G;���9��i6���1�9,,�*�%��� ��^�j	����ǉ�;�%��a,�8y2��n7��;�hZ=�ڦ>�`6?��'?�Y>��<��[9�~�4��>/��&)��|#��>��A�����\!���&��-��e4�F�:���?�	MC���E��G��G���G��$G��NE��$B�ɟ=��8��&2���,�f)���'�$)�+�,���2�_�9�g�@���F�ڹK��AO�ƏQ���R�B�S�"�S���R���P� �M�[�H�9CC��o=�Y\8�b 5��4���5�AB:�qh@�ikG�:QN�2ST��  �  rJ�<�
�<���< ړ< �<n'�<gt�<"ҷ<J�<{��<bT�<F��<���<F��<��<!��<�}�<���< ��<ü<9ڰ<��<�i�<#Ӎ<���<�p<f"a<�NY<(�[<T9i<D^�<�Y�<�ٞ<�Ϋ<���<f?�<$��<��<wU�<'�}<8E_<(iI<,~><v><1vG<<�V<�i<��|<�F�<X�<���<��<��<�ݹ<��<tg�<�U�<mo�<�R�<���<D`�<y]�< b�<�|�<�,s<�[]<f-H<�a5<ï'<=�!<��%<V�3<��I<9c<djz<'��<n��<*c}<X�`<B8<	�	<�޷;�7Q;�S�:}�9x�Y��39�W::�:�Y;��C;|�v;�u�;�Y�;]��;^��;�2�;z��;mh�;��w;ݥ	;��W9�R�C�t������������
�3�P�M���c��Js��Xy��t�[>f�}P�ut8�($��N���
�-�:7M�Ov��*������/���s¼s\Ǽ�Ǽ��ü�ｼ6$��Z2��D`��»��N��xe��/���Z��[���y����`���M��xö���Ƽ��ּb�漐������l`
����,H�����!�P�"��x!�n��f���?��)�
��!������$��'��81�	:��t@���C�]mD���B�e�>��Z:��i5��T0�++�A�%�[� �kp�H��-U��d�v_��K����N��`� �u&��,��1�Q7�|<�h�A��;F��UI��GJ�̐H��D�\n=���5�"�-�r$(��R%�(&���*���1�WY:�]�B�o�I���N�Q�P��O��4M��AI�ָD�E@��B;��z6���1�X�,�9D(��u$�b�!�:!��,"��&%�ݘ)�r /���4���:���@�E�F�ˇL�KR�"�W�"\�g�^��F_�!�\�w�W���P��0I�=?B��=��<�wW>��C���K�F�T�:8]���c��  �  �U<�+X<�{i<�ӂ<oܓ<��<�&�<���<�L�<8��<�*�<���</��<J�<���<�<6��<L6�<���<���<kf�<n�<���<�\�<C�p<��J<i7,<�_<�<�[#<�u?<`+e<I|�<@L�<wn�<L��<r�<Vb�<�k<g�?<O�<"�<&��;�<�<�X:<�u^<�N�<���<3��<��<���</4�<��<��<�n�<.M�<�~�<�M�<M�<���<��<d�<@�<;){<� U<�Q.<�
<G\�;QG�;:��;f�;��<��-<��M<`�c<f3i<�
[<��9<��	<��;�d�:QX���6��h�cV���T�;��:d�>;V)�;3��;�k�;�G�;���;g��;���;���;�I�;�#�;�5t;��;��j97 �<v����ԻU��c�B�j�n�/_��*E��
��M����˔�/c��j�k�P O�<'>�Zi>�x�Q���v��ғ��W����Ƽ�]ټ��㼩��_༯�ԼQ�ż*���4X��E������%���𳆼��͛����������0a��5����
��$��U�Ƽ�ؼS+�} �IZ�%��[�!�
:+�>�1��c4� 3��D.�('���������v�M��{�(�:�4���@��4K�X R���T��S�?�M��F�P=��3���+��$�x���K����D�%���d��g�����a�����u'�\�$��[,��5�}�>�mJH��Q�Y�W���Z��&Z�HRU��*M�]6C�Ir9���1�i,.�/���4���=��}H��S��`[�'`���`�}]��W�w�N���E��H=��5���.��B)�~�$��� �9�����!����Y�@�"��,'��,�M�2��:�ozB�5�K���U��_�`2h�n��_p���n��h���_�vV��M�y�F�X�D�x�G���N���X�b�c�G�m��Iu��  �  <<c�<��1<�U[<�R�<X��<c�<έ�<�X�<�<+~�<�!�<���<���<k��< 2�<7��<h��<=�<���<`��<��<��<xʄ<�4R<]p<f��;v��;{ �;���;��;��,<�\]<�@�<z��<�^�<u��<��h<Ԛ6<��<�
�;��o;hW;��;���;�<�H<�}{<Q��<`��<	ƶ<X�<�C�<���<y�<�'�<V��<���<"�<��<e��<I��<۵�<�K�<��u<�AA<a	<%�;{H;�A�:�3�:P1;��;˴�;��!<O�><�G<�=9<��<'>�;D2�:���뢨�4��R����v������&�NG9�J6;w��;)7�;�� <ic<S<F�<J�<)W<m��;�v�;���;�2W;�ǿ:j;��1Y���лP� ��\�Vዼs����¸�hO¼�1��&������|���!y�`?b�7*`�Yu��Ǐ��$��3	˼�@�0��i�s�ފ��:c��.ӼDQ��3|���_������8���y�K�u���w�3L~�Vs��񾋼�씼I ��;������м����� ��S�<��1s-�c�9���B��DF��D���>�4a5�+�+�N�#����|5!��(�؜3�B�A��+P��=\�o�c��*f���b�
�Z�bO�7�B���5�n4*�Z� ����8��h����	�x	�W	�
�R	�J��[�t8�A� ��*�7�6���C��4Q�#�]�}g�H#l�6�k��pf���\�БP�M�D�o;���6���7��|>�WI��VV���b��l���q���q�~Xl�~�b�L�V��J���=�	W3�P�*�;/$�Oh����s��r����eq��1�%"��B'��.���6�(�A��vN��>\���i�7�u��@~��������]y���n���b�-�W��P��rM���P���X���d��Mr��^~�;v���  �  �;�׸;^��;/�2<�o<�<S˳<6��<�\�<��<]�<���<�C�<��<�i�<bi�<9��<�c�<��<��<�f�<N�<�̚<=�u<��2<S�;�Et;���:�^�:0;#P�;�;�5<��d<Mƀ<̂< �o<��C<V=
<��;���:	�ĸ����Q:�m\;�;͢/<jKn<�<a�<�n�<5��<��<*�<���<�#�<���<�b�<�7�<0��<}d�<��<�_�<@S�<?j<��)<�N�;ކ*;ow��g�����(Z����:�ԙ;���;+j<�+<F�<���;��X;6}���խ���H�0��
8�a|%�*����3���Z���L;*��;<��;~g<xC<.�<��<v&<j�	<{��;<h�;�`�;$�;��
;[pl�0�N�L�ۻ=�0�X�x��П�G徼b�ռ��A�߼��Ҽ����V���Q��Ub��0�|�n����	��'����f�Ł��~��y��h
�ǚ��e�ἆ�ļ�����2������w�8m��9k���n���v��݀�߇��b��7Ț�����g-����̼4������Y���&��]8��<G��{Q�G�U���S��OL�hA���5��I,�!b'��(��#0��<���L�q.]���j�Xs��lu���p�Z�f���X��H��9�^�*�te����+/�����<	�,��.������u	��-�*w��������D+�׀9�'�I��Z�@i�y�t�?I{�V{�u���i�)�[��%N��~C�=(>�YP?���F�C4S�tb��zp�o�{������V��M�y���m�b*_� ZO��X@�f3�K#)��!��z��G�7�����m�����3�i~���Vv$�[�+��%6�"C�	dR�"'c���s��$��2T�� ���+����Ƀ��]{� fm��`���W� �T��>X�P�a�/uo�p�~�6�����  �  ��;�P;���;�<*�Y<��<�3�<u�<۔�<_��<��<bE�<X��<��<MU�<~��<xS�<��<���<a?�<�B�<!��<y�<�f<��<�>�;��:�a_��Rƺ�WṠ�;9�;�<H�M<S�m<2r< HZ<��*<���;]�/;(�"�*-�0aC���Ϻ�P�:�;J<�b<s��<��<@�<?[�<���<��<�7�<��<���<���<���<���<� �<Ÿ�<[��<�$�<�5_<��<�<�;��:�-��_��OQ���4S��E�rE<;��;�f
<C�<`_	<�~�;�,�:��@�g�����6�AzZ�;�`��J������Ļ��I��:l��;���;6�<��<<"<y�<�T<3�<� <w>�;x�;	��;�;&,��f�S���\>�����;���м�������i����弭�ͼI����7�������懼$���P���̖μ���@�
�"H������Q� ��m켴�˼b�������x��Z�r�/h��f��[j�B�r�D~����E-���L��&I��e?���M̼[I����d��,��+@�9�P��[�W`���]�_�U�,wI��<��2��o,��-���5��AC�diT��e��t���}�����z��5o��m_���M��<��H,�7g������� �
����=����$�<���/��
��,����ɇ��b,��><�)4N�ѭ`�̏q�v�~��؂��悽
�~�&�r�@tc���T�d�H��C��ED��cL���Y���i�Ȕy�J؂�
����|��A���x�u��Ke��S��B�j44���(�ԕ ��%����%K������ܢ�l���,����xB#�VN+�^d6���D�e�U�?lh���z������Q��z卽`䌽���m恽t��f���\�~�Y��Z]�w�g�hzv��y�����/���  �  8-���U�˼秗�O�4�V]�c	t;h�<��l<l��<�ե<�<���<*j�<�9�<	�<���<���<ީ�<�T�<�2A<��;�S�������������������������@ǰ� �u����\ûu����\ �|�Q��a����ռ++�~V�����P���漾O��u?^�t`»"�t:���;�54<��g<�^�<+m�<$��<eJ�<�K�<���<ˮ�<i��<�j<U�7<k��;/+�:
t����V�����F漏�	�eH�ש��4�-�
t��M���H�H�(�;��S~�����+����H/�a�<��R=�D�1��,��Y ���ļ�!��z�2�֦Ȼ�/�P��,G:1O�: u�:�J:�I����к�lW�x0���Z���Q��|��h=ʼrN���%��F�-�c��Px�gွ��~�Uzp��/Z�1�@�'�)�-}�+F�?���U2���M��dl��	�������1��#��^���}w��Z���;����\��q�K�Լ`ż����Ð��V߽�SüIk˼��ּ���ƺ���R����S5���Q��[r��<��!}�����P���i��
��ߨ�vf��=�����wQ���W��rn��V����Ǡ�#W��l����ý[}Ľ@���a;���%��R�����-�r�U[��(I��<�73�b-��#*��(���(���)���,�n2��;�s�G�;iY�1�p�rM��.���.��/ݴ���G6ƽ�"ƽ����%���ǧ�b���=]��q!����k쒽	q��$J��ƹ���ĽpYɽ�iȽ�p��@���,צ�c��4ꇽxu�,A`��iP��_E��2>�n�9���7�ə7�.�8�P�:��?��F��TP��_�p�r��������J���T��;Bý�ͽ[_ѽZϽ�ǽм���@���塽 ;�����(��M䡽��������.oɽ\ҽ�  �  C���6⼏���o���z'��}9�>s�;e� <I�k<|C�<��<�+�<3�<6��<�߹<�<���<���<;��<4�<�q@<C��;���9�O�Qq�O������r������;��n�ؼ?0��P�e����W��4B��O@�9C��{���a˼	���
�cF�o�7�ܼZ��/ZR�E���*�:խ�;fZ2<Q�d<Z��<���<��<;�<��<�/�<���<;)�<��f<�5<���;��:A���R<K�7���Iܼq�����g�N����w~���Ձ�cB<�W��w/��Sq�����B��ӳ��)�zC6��37�%,��o��Y��t����8����0�� ʻ�9�}�1�'e:�/�:��m:R:�9���K����d�w彻��vS�䓼5�Ǽ�%�/�"�s�B�`V^��Br�	g{���x���j�'U�އ<�~M&��h��c����w�.���I�U~g�|;��ꊽ�������f�� s���V��9����H��ּ�#Ǽ`Y��$���<����ļ��̼�&ؼ �缡L�������l�4�cmP���o��f��7���1��iޭ��尽���u������2��Za����^��m҅����c�������䖸��뿽*X��h�����������ԕ������r�Y>[���I���<���3�/?.�#�*�g)��W)���*���-��S3��;��:H�fY���o��n�������0��d[���6��MýB�½^
����O���W����������㊊�MA��_w���墳�������z0ƽQŽ!����<��5���O���)����t��``��Q�6F�J?���:�C�8�G8��69��;�g@��F�sQ��j_��r����� ������r(��*����ʽ7ν�>̽��Ľ6�� �����&���韔�c����!�� w���.����ƽEϽ�  �  ��ɼ�N��렢��?l����q���$�;�w"<�<f<�e�<�Y�<\x�<�ݱ<fK�<�X�<s?�<��<���<(S�<w<B<<���;�đ:����R�I�����X�Ƽ��ۜ��ڼ�U��1���s�7��˻�M��-�����N��mgx�sŭ�RT׼����L��X伷#�������X2�4=�����:�m�;� +<MZ<׋{<��<'�<�N�<�W�<Z6�<�o�<Ī|<��[<�.<���;x�:&U��0�,�J卼��������-��E����F���ļz	��.Y��B�)b���o�;AL�#����6μ�o�%.�e�$��&��~�fF
�R/��챼�ڀ�0�,�8�ѻ
�]�@���l�;����9xz�9T�9�4���v��^���#Ի̧��X��V����¼�������}6��wO�zba��i�p�f�dZ���F�Rb0�&���P-�����$��
>� �Y��r��H��"D�������{�R�f���M�G�3������z���ڼ\�̼��ļ�8¼o�ü%�ȼOѼ�0ݼ��� �������g�3��L��%i��l������^��w3���󧽆Z��y.�����-j�������v�Hw��?���b��/2��
L���B��_��:����h�����is���ґ�rG��Ip�z�[��jK��p?��6�i1��i-���+� �+�.-��0��:6���>�)J��Y�8n��5��uѐ�ƻ��g�����O���!���������,��S��j&��y��oM�����_ٖ��?��UB��/���M��裼����뗬��ߟ�iF���D���s�F?a��)S���H���A�>�=��";�Ƌ:�j�;��6>���B�B�I��S���`�-�r�0R��C��FO��-��7��Z���YŽt|ýے���
��������`D���x���C��!��…��!��猾�Ďƽ�  �  ����>���ao���'�S��r��9��;��<,W<>�<*�<�<�<�Q�<���<��<���<��<�0�<Oc<e/<���;P�:DSa������l��#��b���V���e���ʊ���F�MZ�W0�E�����9&Ⱥp��Q�,�U����,��N�V��������ڗ�[a�`��,JC�C��:3��;��<=|D<�<e<tM}<N��<}�<���<�̆<e~<af< F<]�<�y�;_
;��4�
��<`�xo���3���_ʼd�ɼ��������d�;���Ļ�q��ι�5��j�?���5�׼o���[�
�g
�"�a���ɼ�ʠ���r��{-�\��[4��~�3�ɺn�j��;R�������b9h���.����/�
�g�v��mM��!��[���%��K:�� I�R�O��!M� AB��g1��;����$��w���H��5��p,�t�D�U�Z��+k���r�H�p�J�f���U�d�A�z�,����67	����MQ�4�׼��ϼ��˼�r̼u?Ѽ�ڼ����z�������#�!�K�3�P.I���`��ey�Bg�� (��`���ݚ�ș��x���ች��q]r���i���j���t��f�������?����������(y��𬗽����󊁽|�n�̰]�8�O�7�D��p<�@6�'2��0�00�c�1�p�5�"�;���C�a�N�`\��_m�~���1䋽�?������cl��.���h#��.@��Ο�8s��:=��HA��`~����}d��3q���E���ţ�O�H��h
���c���>�����鍽_O��M�s��Jd���W�?�N�z|G�'�B�5�?���>���?��C�?+H�K_O���X���d�� t��P����͆��Pޤ�����:����g���������<]�����^������ =������������������;���;����  �  �5���/�Hf�����|��[��:6�;|�<
7<��^<�h�<FT�<�}�<x*�<^�<d��<#��<+E�<Y�f<m�><j�<�b�;�q;������»����R�#�o��Ks�})Z�w6(�Nͻ�A��0�:�Dt;��;Ca;�Z�Ab��P���iY������\���z�V�X��"���ǻ�L��a�:�}�;�i�;��<wh@<n�[<�o<0y<ty<��o<$�\<$�A<* <��;��;?��:�F��QȻ��$��^��w�������H���:}���H�/
��򛻅P�ZP�����b1�����(q�SM���ļ`mڼ���|ڼ8Lȼ2��f��Eo�ޜ=����߻�f��{u��S<�,}(�{,=��{�bn���9��"R$�íS�;����Š��|��L���4��g�5#���-��1�%+/���%�-�ݫ���������V�mb������A,��R?���M�2UU��U�Q\O��HD�֊6�b(��z�Xr��N�L����꼝��ۼ�5ڼ�x޼���Z���I��6�Wz��)�x�7�dyH��2Z��Ql��h}��ǅ�6e��4̋�����r�����{���l�|�`��tZ�o�[��hd�l�s��q��d7��ቕ����z����M��S���<ɏ���������?q�F�c��[X�zFN���E�\�>�x�9��7��6�3K9�8>�+�D��sM� wW��c�~Cp��2��������# ��j���������Mř������	��כ��kv�zao���p���y�Zo���s��GC��=E���G��9���\ڞ��Q��)���c��=˂�T�w�U�k��a�^X�otP�>�J�JG���E�1G�o�J���P��X��5b�O)m�B�y�����ދ�2���J���:��d���e�������si������_$���D�������͂�;ꄽv������x5������(ت��  �  ^j��������t�׋�H��H��:��e;F
�;n��;p$<
�H<~j<NT�<�R�<+Ӌ<T{�<�u<ΓT<Pj-<=<��;��L;�VB:jҺ}�|�	���I����$��H�ǻe���{��J;�;D��;%d <��;x.�;w�:W�F��4˻O�
�:�A��j��J�仏m���>�c?����:�w;�`�;{�	<cE+<!�D<�ZR<[�R<��E<-<޵<X�;��y;*��:5\S���G��}�������'+��1��&��	�J˽�s�6�0L�6�T;9+;��:C)d�Y�����7�X���������i���.��up���Μ�L�������f���H���*�TC�m�C���祻⊪��/˻�1��+��[�����:���X���tμĜ�������d�����<���S�sh	����� �伯)м�Oü���J�ͼ������1�cc#��Q0���8���;�P�:�*6�Z�/���(�9!�����<���
��I�����S������dm��P�������)��6�[�A�3�M���X�${c�y<m�Y�t�b�y��y�ͻu��qm�\�b�r�W���N�MbJ��K�umS�4`��o��������"���Ď���������ω������W��4�y�Gp�G�f���\��AS��J�]ED���@��@���C���I��dR�� \���e�ƫo�Q+y�'C��>ۅ��2��䍽<Z������D���3��x;��Ŝ|��Ko��e���_�-�`�b9h��0t�fS��C���?���׀��/���_�������t��dg��l%���π���x�n�o�{ef�u�]��=V�^>Q�^WO�[�P���U��9]���f�t�p��<{�ͨ������(p���)����������%��ʘ�S&���ݍ����׀��"y��4v�Χy��o�����ρ��˄�������  �  	;tI:��X�0���Ӥ$�ק����8w�:	o7;[��;���;=^'<�"K<F�a<��f<��X<�A:<��<%�;��F;�':ĵ��.��L��(d��i���Y��a/��]ĺD5�9�u+;cq�;�� <1#<~7<K�9<#�)<@	<i��;�):;��8�v���x��ȟ�%���I=���2���{��`��� �R�뽥�[c�:���;�m�;Ş<� <�y!<6�<���;�I�;2�:�=���Y��Ɯ��񺻽˻`ѻ��λ�ûI��F����t��u}8�;b�;�ͻ;E>�;F�;i7D;���Sl��|S.���[��I~�?Q���u��艘���N��Gӕ�*Ì��+~��\��|8�,�J����}`�X;��Ql�Oo���Ʈ�A
ȼNܼ�'�E;�������9��h' ��b��E����H�X�߼��ͼ����f���0���������2�¼MXܼ5����P
�����# ��'��+��.��D0�L�0�G`/�X*,��&���='��q�ޟ��>�[a�.V
�ʅ���!�*�/���=�{�I��"S���Y���^��a�Ćc��3d��Vc��{`��\[��0T��K���C���=�/g;�|>=���C��M�]YZ���g��t�[>~��ڂ�5J��I���=��'&��QX��ٟ��3��H{���p�ze���Z��Q�M���L�#LQ���Y��`d���o�u�z�����ް������������Dꇽ	��H��p\��&n|��&r��g��\�0(U��fQ�WR�'�W�@a��pl��Ex�0~���ą�cψ�����nы�2?��:���7��b��"^��}"����y��o��Ye��g^�*�[�5t]���c���m�VWy�h����އ�.����䎽����O�����%ᑽ�琽�쎽����nZ��!��Ȅy��0p���i���g�+�j�ĭq�q�{��냽�Ή�ꎽ�  �  ���;:�;8��:Z���+���R`�����yk��̗���;bݮ;�<�%<�-<�<�Q�;�t;\��8��S������h��'ﻞ�ջ�[��QP�;M���|:�+K;M��;���;4� <ްA<�2[<z�i<��j<5�^<�F<B$<'L�;RϨ;�^1;�t�9Ȥ�����)ӻ�r�&���%� ��.��󱝻����J�:�c�;��;���;�_�;�;�}��z���� t��S+�j�&��2��T��M��=yW��ߡ�H�P:�9;e�;���;Sz<h�<'�<�5<��;�	v;�-G:��!��)��#����A�.q��<���-��ӵ������3Ƽ�4�����Q,������� b�0�E��>�R��:}�>��I��x�C�������
����3� �������Լ�żKh���b�� ���(�������͍�O�ʓ���X��KӼ(Y��|�XJ�ܢ�n�$�U/��8��6@�{�D�|E�_�@�"\8��-�ZJ!�nw� ��a��D���%���5�� G��W��bc�u�j��m��(l��g���a��[��7T�RpM�,�F�߶?��9�pi3��/��.���0��*6��[>�	�H�p�S��O_�)Hj���t���~�A&��!���Cy��2�������������Ʉ�=�{�A�m��2b���[�xX[��Da��8l��z��,���J���w��$D���Ǐ��y�������څ�~~��>z��q��g��R^�l6U�^ZM�#�G�;E�f�E�`J�fQ��Z��#d�cn�gx�q���慽K����������t���nY���\���	�������Pw�W�m���i��Fl��t�Y���U���,��� ����ƙ�ј��:��z���Ȕ���X���	��/���8)z���p�Wph�*ta���\��[�Q�]�W.c�%k�y�t��$�`����  �  ��<��;���:>O�T�˻���1=���E�'�1�n��|;��&uI8�/v;��;+��;���;�G;����̻��'��T��Gg�BW]���:��6��V��f�I�Eg7;� �;!p<͘6<KX<�0s<�J�<�k�<��<�߃<��t<R;Y<�6<��<|�;�{0;�s�������/�L�I0{���������o�r��<�~(ﻚaH��2�9_�;�$;l�.:�S2�Y#�68���q�F9������]���\��`#�ʻ����$y:Pe};�h�;��<!<uN2<��9<ߕ6<nO(<N<W�;�5�;D��:���Z�»��"��\i��p��P[����ܼtP������2��X5��Ӽ�o���痼���U|�嗈�#K��� Ǽ-p�|��?7�?$��%�j] �����{����nDؼ~{��;n�����%����T��%vs��o�+v�vw��\Ő�Sq�����"�ϼ.�������[�$�P�6���G�r�U��5_�1_b�{�^��|T�R;F�]�6�Z�)���!�Ew!��Z)�uT8���K�l�`�40s��X��J����Y��A����t�\g�EIY�1~L��nA��F8�M�0�o+�<�&���$���$�'��+�h�2�7;��UE���P��]��j��?z�PL����������.�������
O��gX��al���ŉ�^��.�s�uWk���j�Ipr��)��߈�i����昽QO��*9������(f���M���q��QO���p��Ad�]FY���O�X�G�łA�;N=�U|;��+<��X?��D��]L�z�U��`�5:l��z��Ƅ�(���*���S���s��+����>��w������|��8X����~�n^y��3|�{O��CE��Lp�����A����>���-��dԣ�����ݷ������������j�u�|k� �b�ʈ[�� V�7�R�"R���S�X�/j^�f�f�\sp��{��  �  ��*<$C�;���9"9���.�P"z�5��Bt��S3����r�=�&�ui���,�t�;�Q;l��:ƶ���\�K��y��NE���î�VФ�w���$lJ�ȷ���⺎�P;(#�;��0<�9\<�=}<���<���<l�<�_�<�|�<���<�F}<��\<��2<zK�;�kj;�|���Kڻ��H�]Ď��:���hü��ļ�ѳ�F���WU�h�d�q�����U���]�����[IN�� ��0���dƼ��Ǽ���~䗼��^�i�~�A��#�:�e�;��	<��,<DND<�Q<��U<�P<
�B<��+<��<cJ�;ӢS;����8��3Z�4kw�����޼�����ry�?���d��y�m� m��B���כ����E�ļ����<�)'�B�8�S�A��A�|8���(����	����Xؼ�L��4��U���4Mp�ݔ]�W T�M�S��k[�Ek�'���sj���J��3m����ڼ����I��L*�$�B���Y��m�l{�����K|��Bp�y�^���K�*;��1�a0��8��TJ�]Aa���y�󐇽����?�����M��揂� ,q��]���J��;���/�L'�M�!�l!�����z����=$�ZC*�R2�n�;�,�G�J�U�&Ag���{�����s�����Z�����EM�������֟��{��?銽
;��vz��y�+���b≽�b��8ꞽo��%S��˴�������Π�!������ʣ��'�m�Yv]�ukP�>TF���>�cF9���5���4�|65�4�7�:j<�!!C��L���W��f���w��h���͑�p7���Y��Qɮ�M��9<���ū�{���#���z����[���#���Ʌ�������n���}ݪ������3���>������n��t�����������6�|�Cn�nGb��RY�O�R�62N�k�K��HK�{�L��/P���U�IE]�v)g�O�s��  �  ��.<:��;�s������Lt�gk����Ǽ\kҼ\Ǽ˨�lz����T��� J�G�9buغ�0���y=����$뼼��ټ�q�Lռ�_���慼�� ��TU�4"4;5��;�A<�jq<�͉<�K�<�8�<�M�<��<���<�ϔ<���<��r<@�E<o�<�h;��6*� ���.���}�ݼx�������R�_���:���D�k���E�������޻�;����Z2������~������Ǣ�ﾼߌ���,�>L����:!=�;(e<V�A<�Y<T�e<9�g<
a<�&S<x�=<M� <w��;ْ;Z3:	����}!������¼�����R��-� `7��6�"�+��p�)M���ܼ�9���������� ��L	�J�$��X>��Q�I�[�JZ��nN�Mw:�H�!�(���޼ⴼ-���5y��Z��H��|@��A���J���Y���o������r��B����Ӽy���w �?�1��O��Qk�����䉽T�������	�s��?]���I�z�=��O<�`�E��uY��Ls�lg������ڛ�]������b��v���lJ|��#c�siL��9���+���!����������i��������%��y,�Y&6���B���R��Jg����&p��}���}���������gN��g���+>���]��Q;���H�������D��Ts������D+��#⳽0T���o��@0����������I�������Ln�k�Z���K�f�@��+9�U4��?1��70�R�0��3�(7�6�=���F�%KS��d��Ny�ND���(���������ֳ��5+��/��� ���譽��v�������c��~;��mP��:���ͪ�ʒ���C���6ý��������e���u��镽�'���E|�#�j�4E]��S��AM��5I��4G���F�R>H�vAK�FP�G�W�lb��p��  �  ��,<���;KU7���+� ���Ƽ��� ���9�$�ȼ����SI�A�ػ�U=�
��7Vz�f����n�n���8�ݼ�����{��;�Ѽy|��#1C����Q�;��;'�G<��{<3��<2�<�U�<`�<㣣<���<<�<�u�<��}<� N<��<�T;�T���-��X����ϼd����g��.�;�g༝�����p�Z����һ�2λl(�"yg������ܼ�S�J�	��\��U�ڼ${��S�J�&,����:�"�;�"<�L< �d<��o<��p<p�i<�[<5_G<�A+<|h<���;8�:����K*�Н��LeӼQ�
��'�U�=�� I���H�Z�<�R0(�����&4ѼPż�ѼQ��;���12��N���b�@Vm�}`k���]�7G��Y+����*��\���鑼p���N�U�<��6��8���A�_�P�e�e�
j���피���'ѼZ����/���7��\X�9�w��C��j�������������ڿ����h�ɳS�vF��zD�x�N��c�uc�����t������l˧��줽>����z���`��s^h�
�N���9���)�aI�������4=���� )�{���H"�\�)�V3��@��R�S�h�Ł�j��������2��¯��yb��^.½t����벽����eʘ������ʇ�1w��J�������������P��2½`0½�?���f���Y����������o��=Z��I�\ >��D6�ea1���.��-�*~.�e0�c\4��:�wD�֍Q���c�cf{�����P@���֪������½[�ǽ��ƽ�E���@��q5��Λ�����e���손�A/��������fw��N�ǽu̽8Fʽ��½W̶�EI������Ί��}�=ti�o�Z��P��aJ�ɎF��D�X�D���E���H��iM��T��_�n�n��  �  �~+<%ׅ;��[�ڡ9�"��;�Ѽ\���,P��m��Լ Ң���Y� ���>n�y�)� !���;����E'���7���>	��7�-ܼg���O��b���@�:V��;dI< �~<v[�<_��<<�<�W�<,��<7�<{�<�A�<h��<�lP<BD<��J;� m��$8���sBټ{����p�C	
����;��[��K�'���)���1!�G�v��8���6缞M	��Q��,�h�����^��4V�Vٷ���u:*�;��$<R1O<xh<j"s<S�s<l<W>^<�EJ<��.<��<�x�;]h�:g=���
.��z�� ټ���!�,��C��nO�<�N��vB�!`-��D�NH��-�׼"˼R�׼�������h7���S��i�Ȧs�f�q�jTc�0�K�v�.�{x�y��KJ�����مm���K��.9���2�v�5�9,?�$�M�0�b��]�;��ܘ���м����Hl�~:�H�[��U|������r��**��[�������q2���m�:&W��vI��XG���Q�/"g��Ӂ����kw���������姽FB��������Igj�u�O���9���)�I��� �J��pp�����v� <��l!�6�(��}2���?�vR��#i�����H��ǌ������p����|Ľ�UŽ���&����Q��Ͼ�����MF��p�������j���⦽qi��L���XŽ�OŽw#���᳽�O��h������p��7Z��JI��P=��^5�[�0�(.��A-�/�-��/��}3���9��OC�NQ�`d��Q|���� Ŝ��묽L��*�Ž�$˽� ʽ�2ý�׷�Xi��(���Q0�����	���噽��L��A����ʽhEϽ.Wͽ��Žv�����K��dz���x}�!<i�QZ�!P��|I���E�JD���C�+E���G�F�L��S�.�^��n��  �  ��,<���;KU7���+� ���Ƽ��� ���9�$�ȼ����SI�A�ػ�U=�
��7Vz�f����n�n���8�ݼ�����{��;�Ѽy|��$1C����Q�;��;'�G<��{<3��<2�<�U�<`�<㣣<���<<�<�u�<��}<� N<��<�T;�T���-��X����ϼf����g��.�=�m༥�����p�t��1�һ�2λ�(�lyg����Ʉܼ�S�|�I������ڼ|��m�J�#0����:"�;�"<�L<��d<"�o<��p<��i<�[<{yG<`a+<*�<��;/:�����*��~��@EӼ1w
�+�'��=�cI��H��<��&(�������U.Ѽ�Nż@�Ѽ?��w��:2�9N��
c��cm�fok���]�:GG�j+�j��H�sx��g���6p��O��<�+(6���8���A�L�P���e�I]���ܔ��خ�lѼ����� ���7�ALX���w�s;��Ub������!���k닽I�����h�+�S��sF��zD��N���c��j�R���A��������ҧ�������������/i��:oh��N���9�)�)��U�]�����E���@.��� L"�χ)��W3�T�@��R�؅h�<Ł����������2��̯���b��d.½y����벽����gʘ������ʇ�2w��J�������������P��2½`0½�?���f���Y����������o��=Z��I�\ >��D6�ea1���.��-�*~.�e0�c\4��:�wD�֍Q���c�cf{�����P@���֪������½[�ǽ��ƽ�E���@��q5��Λ�����e���손�A/��������fw��N�ǽu̽8Fʽ��½W̶�EI������Ί��}�=ti�o�Z��P��aJ�ɎF��D�X�D���E���H��iM��T��_�n�n��  �  ��.<:��;s������Lt�gk����Ǽ\kҼ\Ǽ˨�lz����T��� J�G�9buغ�0���y=����$뼼��ټ�q�Lռ�_���慼�� ��TU�4"4;5��;�A<�jq<�͉<�K�<�8�<�M�<��<���<�ϔ<���<��r<?�E<m�<�h;!��9*����1�����ݼ}�������Z�_���:���D����[F��Y����޻��;�����2���伦��������弓�������,��S��֪�:b;�;(g<*�A<��Y<֡e<��g<�1a<VOS<]&><� <�n�;���;�Q9:𸄻�!��C����¼i���4�{�,��D7�#�6�X�+�n^��>���ܼ�.������(���W��V	���$��l>���Q�ľ[��fZ��N�w�:���!������޼����\��W�y��_Z��8H��@���A�=�J���Y���o�2؆�&R���]���cӼ���D�U�1���N��1k�k����Չ�y��)㊽�냽m�s�T2]���I�!�=�P<�Q�E�Y��Zs��p��>����盽��������r������k|�CDc�o�L��9��+���!�d������������������%��~,��)6� �B���R��Kg�;��Wp��0}��~���������tN��q���3>���]��U;���H�������D��Vs������E+��#⳽1T���o��A0����������I�������Ln�l�Z���K�f�@��+9�U4��?1��70�R�0��3�(7�6�=���F�%KS��d��Ny�ND���(���������ֳ��5+��/��� ���譽��v�������c��~;��mP��:���ͪ�ʒ���C���6ý��������e���u��镽�'���E|�#�j�4E]��S��AM��5I��4G���F�R>H�vAK�FP�G�W�lb��p��  �  ��*<$C�;���9"9���.�P"z�5��Bt��S3����r�=�&�ui���,�t�;�Q;l��:ƶ���\�K��y��NE���î�VФ�w���$lJ�ȷ���⺎�P;(#�;��0<�9\<�=}<���<���<l�<�_�<�|�<���<�F}<��\<��2<uK�;�kj;}���Kڻ��H�aĎ��:���hü��ļ�ѳ�V����WU�Oh�}�q����AY��K�]�j���\JN�Q!�����eƼ�Ǽ�!���旼��^��!��A���:Fc�;��	<��,<@]D<g	R<�V<��P<��B<H,<i#<1�;9�U;���\������v� �����ݼ|��X���R�%��1F�`�N���P��$2��7ԛ�&!����ļ����S��7'�x�8���A���A�צ8���(���- ��ؼ����5Q���ֆ���p���]��RT��S�5n[��.k��o��9G��0���3��kMڼ�A��� �� *�UB�X�Y��jm�G�z�.��q(|��$p���^���K�q;��1��0��8�UbJ�@Ua���y������,��T���̐�8-��^���[q��5]���J�&�;�@�/��m'�ݫ!��:������d
 ��H$�:L*�2�J�;���G���U��Bg���{�_���t�����=Z�����XM�������֟��{��E銽;��$vz�
�y�-���d≽�b��9ꞽo��&S��˴�������Π�!������ʣ��'�m�Zv]�ukP�>TF���>�cF9���5���4�|65�4�7�:j<�!!C��L���W��f���w��h���͑�p7���Y��Qɮ�M��9<���ū�{���#���z����[���#���Ʌ�������n���}ݪ������3���>������n��t�����������6�|�Cn�nGb��RY�O�R�62N�k�K��HK�{�L��/P���U�IE]�v)g�O�s��  �  ��<��;���:>O�T�˻���1=���E�'�1�n��|;��$uI8�/v;��;+��;���;�G;����̻��'��T��Gg�BW]���:��6��V��g�I�Eg7;� �;!p<͘6<KX<�0s<�J�<�k�<��<�߃<��t<P;Y<}�6<��<|�;�{0;s�������9�L�W0{�����ø����r��<��(ﻣbH��'�9��;��$;��.:�W2��%��8���q��:�������_���\��f#��ʻ�����x:/_};o�;��<I1!<k2<��9<�6<Ζ(<R�<��;#6�;�5�:X��,}���"���h�����＼��ܼ0��_\������u��2�Ҽ�>���ė�����M|�+����e��J*Ǽ�����_��F$��%��� �j'�����w��4�ؼ�ؿ�����@O���1������ʹs��o��-v��i�������E��Ef��Cϼ��gW��[���$�0c6�JMG�l�U�,_��/b��d^��WT�F�O�6��)�J�!��w!�|c)��d8��K�	�`��Vs��n������Dt������t��Qg���Y��L�>�A��t8��1��'+���&��$���$��'�(�+�J�2�F?;��[E�ТP��]���j��@z��L��惍�����V�������"O��yX��ol���ŉ�f��:�s�~Wk���j�Npr��)��߈�j����昽RO��+9������)f���M���q��RO���p��Ad�]FY���O�X�G�łA�;N=�U|;��+<��X?��D��]L�z�U��`�5:l��z��Ƅ�(���*���S���s��+����>��w������|��8X����~�n^y��3|�{O��CE��Lp�����A����>���-��dԣ�����ݷ������������j�u�|k� �b�ʈ[�� V�7�R�"R���S�X�/j^�f�f�\sp��{��  �  ���;:�;8��:Z���+���R`�����yk��̗���;bݮ;�<�%<�-<�<�Q�;�t;\��8��S������h��'ﻞ�ջ�[��QP�;M���|:�+K;M��;���;4� <ްA<�2[<z�i<��j<4�^<�F<B$<#L�;MϨ;�^1; t�9ޤ�����)ӻ�r�*&���%�:�'/��J���e�����:�b�;��;���;^�;��;��������!���v�4W+���&�8�Ya�=[��t�W�����P:�9;���;��;1�</�<<�<�u�;~�w;�0P:�_�����& �eA�xEp�HŎ�����f]���{����ż�����ǲ��杼"J����a��VE���>�(R��u}�i��܇�����;!���4�J�!�
����u� �=�6Q�`Bռ�Ƽ���������4��WL��:���Uύ��ᖼDs���'���	ӼL	�,N��'j��`$���.��^8���?�E�D���D��@�338��,��0!�Sf����b�N���%���5��CG�D0W��c�W0k�g�m��fl�
�g���a��D[�'tT�ۨM��F���?��99�Ռ3���/���.���0�h:6��g>� �H� �S�'T_�:Kj���t��~��&��t����y��a�������������Ʉ�T�{�S�m��2b���[��X[��Da��8l��z��,���J���w��$D���Ǐ��y�������څ�~~��>z��q��g��R^�m6U�^ZM�#�G�<E�f�E�`J�fQ��Z��#d�cn�gx�q���慽K����������t���nY���\���	�������Pw�W�m���i��Fl��t�Y���U���,��� ����ƙ�ј��:��z���Ȕ���X���	��/���8)z���p�Wph�*ta���\��[�Q�]�W.c�%k�y�t��$�`����  �  	;tI:��X�0���Ӥ$�ק����8w�:	o7;[��;���;=^'<�"K<F�a<��f<��X<�A:<��<%�;��F;�':ĵ��.��L��(d��i���Y��a/��]ĺ@5�9�u+;bq�;�� <1#<}7<J�9<"�)<?	<f��;�):;���8�v���x��ȟ�3���\=���2��|��������R�����a�:���;cm�;b�<o� <y!<_�<���;G�;���:;P��MY��͜������˻�'ѻ��λ4)ûR�������e�Q�8�2;A��;�,�;n��;Б�;��E;�F��]�i�f"���-���Z�d}��؊�������Xw���ڙ��f��a����}��[��8�s���R�_��;z�@;�y�l��������fȼ�ܼ]�뼳�����������d �{������q���߼�%μ�=������D���¥��쯼 �¼�$ܼKy�� '
�~S������&��+�Gm.�80�*[0�6%/���+�({&�������W�U���5��a��_
����N�!�6"0��>�=�I��[S��'Z�3�^�E�a�0�c��td�4�c���`�ޒ[�baT��L��D��>���;�TS=�-�C���M��bZ�ǲg��t��A~��ۂ��J��ɪ��j=��m&���X�����Q�I{���p�ze���Z�!�Q�$M��L�)LQ���Y��`d���o�v�z�����ް������������Dꇽ	��H��p\��&n|��&r��g��\�0(U��fQ�WR�'�W�@a��pl��Ex�0~���ą�cψ�����nы�2?��:���7��b��"^��}"����y��o��Ye��g^�*�[�5t]���c���m�VWy�h����އ�.����䎽����O�����%ᑽ�琽�쎽����nZ��!��Ȅy��0p���i���g�+�j�ĭq�q�{��냽�Ή�ꎽ�  �  ^j��������t�׋�H��H��:��e;F
�;n��;p$<
�H<~j<NT�<�R�<+Ӌ<T{�<�u<ΓT<Pj-<=<��;��L;�VB:jҺ}�|�	���I����$��I�ǻe���{��J;�;C��;$d <��;v.�;`�:^�F��4˻R�
�:�F��q��\�仦m���>��?���:(w;N`�;B�	<E+<D<8ZR<��R<��E<-<��<�T�;0�y;��:ܓS��H�釬����)��~-+��1�	�&��	�B����F6���^7;�4,;�{�:h�]�����`��W�9,��]��������������W���0������Ie�H�N*�|��k���q�� ����x���`˻�k���+��[�f���W����跼��μ���Q�������`����1����	����� ��Mм�bü����f~ͼk�������:#��"0�Z8�;�[X:���5�ݘ/��k(�, !�����"}
��(�̚�����҄�"����I'���7:��)��H6��2B�>�M���X��c��|m�h>u���y�.z�;�u���m��b�x�W���N�u{J�j�K�t}S�x`�'�o�o��.��:$���Ŏ�>�R���ω�>���2X����y�OGp�u�f��\��AS���J�kED���@�"�@���C���I��dR�� \���e�ǫo�R+y�(C��>ۅ��2��䍽<Z������D���3��x;��Ŝ|��Ko��e���_�-�`�b9h��0t�fS��C���?���׀��/���_�������t��dg��l%���π���x�n�o�{ef�u�]��=V�^>Q�^WO�[�P���U��9]���f�t�p��<{�ͨ������(p���)����������%��ʘ�S&���ݍ����׀��"y��4v�Χy��o�����ρ��˄�������  �  �5���/�Hf�����|��[��:6�;|�<
7<��^<�h�<FT�<�}�<x*�<^�<d��<#��<+E�<Y�f<m�><j�<�b�;�q;������»����R�#�o��Ks�})Z�w6(�Nͻ�A��0�:�Dt;��;@a;�Z�Db��Q���iY������\���z�\�X��"�Эǻ'M�a�:}}�;�i�;\�<Eh@<,�[<Zo<�/y<�sy<�o<6�\<��A<� <��;��;ʓ�:�U��ZȻ��$�9�^��y��K����H��
7}���H���	�G���{������e��~y��~I���p����Bļ0ڼ2 �Gڼ��Ǽ��������{n���<�%r��޻]s��X�s�SI;���'��=��u{�հ�t�����$��4T��I��w������s6㼚j�ٝ�(j#���-�i2��U/��&��K����L������`X�!T���eq��#,�k.?�@�M��%U��mU�t&O�dD��S6���'��G�dC��$�r���U^�.��p�ڼ�'ڼ�y޼ ��28��a��U�ß�v.)�2,8�?�H�`jZ�R�l�x�}��ㅽt����勽Z׉��Ȅ�'�{�"m��a�:�Z�˔[�wd���s��u��b:��������y���^N��ϔ���ɏ����	���?q���c�\X��FN�̡E�m�>���9��7��6�9K9�<>�.�D��sM�wW��c�Cp��2��������# ��j���������Mř������	��כ��kv�zao���p���y�Zo���s��GC��=E���G��9���\ڞ��Q��)���c��=˂�T�w�U�k��a�^X�otP�>�J�JG���E�1G�o�J���P��X��5b�O)m�B�y�����ދ�2���J���:��d���e�������si������_$���D�������͂�;ꄽv������x5������(ت��  �  ����>���ao���'�S��r��9��;��<,W<>�<*�<�<�<�Q�<���<��<���<��<�0�<Oc<e/<���;P�:DSa������l��#��b���V���e���ʊ���F�MZ�Y0�������9+Ⱥp��R�,�V����,��O�X��������ڗ�ba�h��XJC�ϔ�:��;o�<|D<�<e<>M}<+��<�|�<i��<�̆<�~<`f<�F<��<�u�;�
;��4����@`�|q���5��aʼ|�ɼ���h���'d�����_Ļ4��YU���l�Ԭi�b���4N׼�J��0�
����O���/�7|ɼ�t����q���,�����F���!2���ƺ�Rg�GVP�s �x��m�h��o���) �Cp/�dh��a��o��� �I;���%�jw:�j*I��O��DM�f_B�À1�?O����'������t�R)�;^,��D�s�Z��k�Ѩr�Y�p�8rf���U�Z�A���,�qw�	�?�����׼
rϼķ˼�f̼I@ѼMڼ���à���4����{�!��"4�fYI�.�`�۔y��~��R?�������#���z���1�.Ѐ��sr��j�ӭj���t�-k�����FB��i�U��Ū�������y��?�������!�����n���]�\�O�Q�D��p<�%@6�'2��0�60�g�1�t�5�$�;���C�b�N�`\��_m�~���1䋽�?������dl��/���h#��.@��Ο�8s��:=��HA��`~����}d��3q���E���ţ�O�H��h
���c���>�����鍽_O��M�s��Jd���W�?�N�z|G�'�B�5�?���>���?��C�?+H�K_O���X���d�� t��P����͆��Pޤ�����:����g���������<]�����^������ =������������������;���;����  �  ��ɼ�N��렢��?l����q���$�;�w"<�<f<�e�<�Y�<\x�<�ݱ<fK�<�X�<s?�<��<���<(S�<w<B<<���;�đ:����R�I�����X�Ƽ��ۜ��ڼ�U��1���s�7��˻�M��-�����O��ngx�sŭ�ST׼����L��Y伹#�������X2�D=�����:�m�;{ +<6Z<��{<��<�<�N�<�W�<%6�<Fo�<�|<��[<�.<߲�;��:JY����,��捼���̯��.��F���aE鼺�ļ����Y�*���� E��L��ԕ��μ�Y�s�S�$���%��`�Z'
�)����������,���л&R\��^��ׅ.�pl�9R$�9�8����j��������Ի����Y�_���r�¼�X������6���O��a���i�Cg��yZ�n�F�p0�y/����-����x�$���=��|Y��vr��<��`6��������{�d�f��M�P�3����������0�ڼ�̼{�ļ�'¼C�ü��ȼ�XѼ�Bݼ�(�:� �4���Y�3�}�L�Fi�`}��O����n��JC�����Bh���:���(���s��������v��Rw��C���e���4���M��D��>��Յ��^i��a����s���ґ��G��|p���[��jK��p?��6�s1��i-���+��+�.-�
�0��:6���>�)J��Y�9n��5��uѐ�ƻ��g�����O���!���������,��S��j&��y��oM�����_ٖ��?��UB��/���M��裼����뗬��ߟ�iF���D���s�F?a��)S���H���A�>�=��";�Ƌ:�j�;��6>���B�B�I��S���`�-�r�0R��C��FO��-��7��Z���YŽt|ýے���
��������`D���x���C��!��…��!��猾�Ďƽ�  �  C���6⼏���o���z'��}9�>s�;e� <I�k<|C�<��<�+�<3�<6��<�߹<�<���<���<;��<4�<�q@<C��;���9�O�Qq�O������r������;��n�ؼ?0��P�e����W��5B��P@�:C��{���a˼
���
�cF�o�7�ܼ[��2ZR�N����)�:ǭ�;]Z2<E�d<R��<���<��<+�<��<�/�<���<)�<L�f<��5<;��;��:_����=K�砣��Iܼ������g��M���⼐{��с��5<��E��a/��7q�꫼yr�l��)�o56��$7�],��_��9��f�����Lv0�w�ɻ�Q9�O/�$!:�˄:�sn:��9	��s��De��$��_8�F7S�����dȼ�5�D�"���B�Tf^�;Rr�Mu{�m�x��j�j'U���<�^R&�k�d���� �.���I�Zug��5���㊽�
������^���s�N�V��9�ϸ�::�0ּ^Ǽ`L��b��W8���ļ��̼(0ؼ��缙^���������4�}P�G�o�Vo���%���:���歽S������������7��e��͝����ԅ����������������� 쿽{X������Ы������ԕ������r�m>[���I���<���3�4?.�'�*�g)��W)���*���-��S3��;��:H�fY���o��n�������0��d[���6��MýB�½^
����O���W����������㊊�MA��_w���墳�������z0ƽQŽ!����<��5���O���)����t��``��Q�6F�J?���:�C�8�G8��69��;�g@��F�sQ��j_��r����� ������r(��*����ʽ7ν�>̽��Ľ6�� �����&���韔�c����!�� w���.����ƽEϽ�  �  t󤽭ɟ��搽b�u�3�A�ʸ��p��.�G�����f;���;�<�a/<��<<��><��5<6� <%��;�J�;�*��\�6y��s�޼��"��=Y������⛽eW���������_���#��BQ�o�*� �����W����@��Pm�����R����}��XK�����9ǔ�k�y�lqD�����\��7"e�r�ӻ�jw���=;}L�;���;��;�2�;��;��;��T;� ߹c!��3\U����VE
���>�q5t�`�������ʯ�󱯽ۀ���p��Z�z�V�O�mi/��Z ��&���?�z�i�;�h��2����Ľ��ý���i��Ս���g��86�� ���мo+���3s�)�F�Le/�u(�'�-���>���Z�d��蟼�ȼI&���"���N����6,���W��M�ν;�߽{"�m�㽱׽�|ý�A��A0��ы���5���;��=�������=�˽^i⽮h������v���G��нdd���c��o���Tb���B��x+�X�����u������k5��P��)��v9�m�O���m�]����%��}���tn׽1���8=��p��r
�U�ޯ��6ܽ\Pʽ�ӿ�����OȽ�-ڽ]�h��������i��J��[��)���3�޽��ĽjŬ�[䘽�R����{���k��+a���Z�<�W��W�~+Z�V�_���i��y�F�������1 ���h��|�۽Ш��4��u��*���Ծ� v�L#����Ὠ�нO�ǽ�ɽ�eԽ�罹���[�
��h�h��������#��C���ڽ����e���K���~��k�����s��k��g�G�e���f��#k��r���~��R��Yݔ���������]ӽ�]���3��k�����	�<V�$-	�R��1Y��׽`Mҽ�0׽߄彡���>	�M��fP��  �  *��������U�� n�X<�)��^x��ҧE�`	�� E�:dN�;-E<�=)<="7<�%9<@�/<�<b��;J~;~{q����҃��(ڼ���G%S����,���$��G\���^��`����w��J�[�$����G�	�����p:�g�e�k��������/����������@t����r�Dl?�2��p���d���ڻ��c�#;�;ߡ�;1��;���;�;)��;ɯ:;��J��aû�^U�����Y�T�9��m�jq�����녪��d��z��.����s��I�]%*����g0!�z:��;c����ס�&�����������Ma���
��;����lc�j�3� 5
��vѼ�Y���Ky�2pM���5�!�-�jA3�J&D�:�`�χ�����# ˼M' �"z"�`�L���}��i��c���yʽ��ڽ��Ὀ�޽�:ҽN6������G6������ф����8ٙ�l����ǽ�ݽ:9�ހ�c｡��7ͽt���/���bw����a��C���,�J���|�����+�Zv����h��[�*���:�l�P��n�s���vo��RYԽ(�^����.�
���E� �_���ؽ7wǽ
P��������Ž�׽5��T|��F�E�zO�1�z���9���rܽ��½�	��(Ә�Z����}�KOm���b�;T\��7Y�W Y�d�[�c�a�ˀk���z�m������,Z����qHٽ�K�ʇ�(�� ��oZ�;�K8��S����޽�ͽ|QŽ+�ƽ-�ѽA:�!����_����]�U�������ģ���׽m_���詽i����*\��x�u��$m�K�h�*g��dh��l�)bt��3������s/��e������	�ѽ��뽻��@��p���6��h����-����4^��$ս��Ͻb�Խ���x����wo�����  �  ����V���;�4QY���,��r������kC�����D$:���; l�;��< �$<P'<Ջ<�<9^�;z�.;B���%�����ͩμ�����B��Lo�@��"���kR��Pԑ�8r��F+`�9a7�����X��������
���(�~�P�y3z�����A��-������r����_�9�1�x�����_�f�D����}�:^�w;)��;(��;��;n��;.s�;�>�:�'����޻�(Y�@��������,�i%[�S���U��������y��/b��d����]���7��"����Wm�s+���P��}�W锽f@���ү�A	��I���▽�.���W���-��~��Լ�������DQb�J�I��q@��D�V���s�R��������Ӽ7���,"�E^H�qt�� ���z�����s̽r�ҽ��Ͻ�uĽ!���~������ض��<�{�����֜��:����軽})н-�޽h��K%�4ս��½���������(��Va�)�E�j1�g�"���l�����-��&���#�Ę/���?�K�T�$�o�6È�Z���-᳽� ̽�㽼0���O��3��� �@
��'��*Ͻ_���(��ƚ��5���0ν����v���=���
�����=��� �;�콜�ս�����n��%���Q��x݀��xr�*�g�Ua���]�{]�[`�B�f�w�p�0G�������z��� =����ҽH��N��������|#�u������H�սAƽ�a������u�ɽ��ڽU�ｩ��M�	����I����ߙ��3齹ҽ
:��( ���2��5댽�у���z�*r��,m�ȅk���l��xq��y�MÂ��-��艖��O��x���ͽ=K�8Z�����^��Ʒ�U�[
���"���ڽ�ͽɽ�lͽ�Fڽ)�����
�|U��  �  �Nu��1o���Z�xq<�%u���,2��fL��һ�ͺ��;!�;n��;��<�<�.�;h��;�Jl;^��9����;��Q��~�ür#��R,���P�qgn��p��sT��0�x���_��!>����n����Լ�hμ^�_�1�H4U���s�/\��^b���\��f��E��� ����ꬴ�c�v��F�t���
����c�:�gW;kc�;�;�`;ST�:� T��΋�����j�ƭ�>��%��]B��\d�Ν~�:�������0{��{_�`�=�#*������{������)5�Z�\�qɁ��/�������ݚ���D:���Sm���I�~Y'��	�'�߼�����b��� n��b��e��|v��#���,��?7��Zz弼q	�R�$�	 E�<}i��>���j��y���ݷ��ͼ�����$���3��~Q�����m��xg�Нq��C��o喽�o���@���ɽ��ν��̽ý�g��9뢽~�=��S�c�/1L�\�9��u,�	#��x�,��-��10#�"M,���8�� I�	]�H?u�i$��y��X�������G�ӽJ��h�T�.���]ེ�н*����9��|f�����x�������{ ӽ������ë���� ��r��dG��߽�ͽ�~��5������@��p���A|��$q��i�8�e��e���h���o��sz��d��q���E�������1��©ʽ��ݽǵ������O��� ��`�����jٽ�0Ƚj˺��򳽈���꽽��̽��޽�_�a��K��XX�'������Foݽ��ʽ�	���0��{ݛ�e��w���5��m1{��u�2�s��#u�N>z�<|�����=������v���u��e�ǽ<�ڽb_�{���������"������^]޽�,ν&�½i�����½Z�ͽ�4޽i�𽢜 �����  �  �*C��@�4v3����&��N�ּ���;�o�+v�[����b���:\�m;y��;8ݫ;��;�H*;��0��+q�������L��ґ��y¼Fc��'��x0��E�8Q��9R��CG�"�1�����}��������d�������d�ݼ����)�MuC�a:T��jY���R�`B�c+��V��,񼼙�����R�<
��G�����'8��:t�:�\9ծ�c�������J����^᷼���6���)�	A���R�1�[�q�X�u�J��3���[����QӼ¼��˼)��Y�r�5���V�H|q�^뀽�����D~��lm���V�:<>�I&���_����2׼j躼L��ƅ��l֊�7 �������ɿ��߼���+��-��G��Gb���~����������Ҡ�kƣ�ؠ��m����s�|���c��_S���N���W�;m��e���ܕ�����j>��<䵽�j��N{�����c�������� ��X�l��Y���I���<�2��+�(��)���/���9��H���X��=l��Ѐ������������{����rýA�νD{ս׽l�ҽTɽ8¼�����k����~��V���������dX���н��ݽ!c�,G��%��ݽh{ҽe^Ž���>����_���g������������v��@r���q��v��d~�$��$������@垽s���=]��֤ýK�нv�ܽ��� 꽈�轵�b�Խ�]ƽ�"������n��"a���ï��$���˽��ٽM]彰��j�콚��E1޽Sҽ�Ž�A��D}�����YΘ�'ʐ�� �����D������׀��냽�������[×� ����q��a4���&Ľ~�ѽ�߽kc��|���!#����ڽ�X̽����.����@��B����徽>�̽�۽C������  �  �t����-[�2��>���8ؼ����&��qV|��F<�����+��m1��N�=:���://�8�$�w۷�#X�ASb�`O���T��fZԼ��󼖻�!��h���
$�� ����e����ټ+��#���X���P�~	s�.`���]ʼ1�����g"���)��)�I�"�2���
�������ؼ���ׂ����p���/�5��H	���vD��C?�Ǔ��m=໣)�ߞi�����Vf��/�ռ2���������"���*���,��z'�m��W�)��Xs���4����2��i���伨�`z)�1�@��P�oyX�JEX�U�Q��G�L;�3.��� �����T���RѼA���q���
d��=����˼�3꼐m�s���e.�WA�H�R�4�c��Nt�Ӝ������\D��/����⇽O����/m��W��~D�8��'5�5�<��lN�'�f�/߀�����⒗�T�����������̙�����Wf��U����I��q�]�b��kT���G��>��89�:���@��UM��]���p��2���Ӌ�����흽�����������»��Ǿ�A��ع��������ޝ�2�������YZ���Ֆ�=�����p�(KŽ�mͽ�}ѽ^�ѽ�-ν=�Ƚ�����E��n���,���:i��X��������[�����#����p�� /�����f����ј�Q7��Zq���e��M%��b�����ǽU�ͽ$�ѽ��ҽ�Ͻ��Ƚ�����̲��~���Ğ�3X��X"�����᪽9ݶ�#�½U�̽�8ӽ4�ս�oԽOJн^Sʽ�pý�-��@����
��N������H��x���+5���[���v���j������{����#����������7��Ž��̽
�ӽ�hٽ`�ܽlܽ;ؽ<н\~Ž�ǹ�z;���姽�D���짽�f��;K���ƽ)$ҽ۽�  �  I�ҼR.伜�����i������~�u�ټ1
¼ r��p�{�*12�����ї�Is���%���	�voP�����ᵼ<7ּ����(
��6�n[��W�v�������jԼ)����T��W�S�=��v��ݻ%���>��e������\�ϼ�p��t�$�	�����?�������`������5޼�����s����a���'����?#���"�6�Z�5R��������ڼ�X����8��o&�:$�GH�-G��_�����G�޼BM��ڥ��#�x�J7M���=��0O��c��{�����ҼY� �L����&�ń3��<�4>A���C��}D��{B�F7=��
4���&���4S��N�4�ۼ�~ּZa�؇�������&��<�/.P��_�%�j���q���u�I�w��Zw�zt�OIn�`2d��ZV�;�E�JG5��"'�(Z����z�#���1��SE�Tn[��q�����YV��{������u���JE���쓽�@��]ߎ�J����_���5t���c��sV���N���N�v�V�a1f�pz��_������J��[\���J���r���J��g���魽Oa��b���룽������a��&Z��{D���넽�p��_?��/��Yȥ�Ϧ���Ƿ�ӵ��i�����ý�ZĽ�
Ľ�½~���=�������.Ǫ�y���ٗ�^����X�����ˏ��ɖ��ٟ�n����j��u���sϾ�.½��ýXTĽ��ýY½�9���&��'���>���Ơ�.����S�����/���`/��tӚ�VJ�����(���q���ý�!ƽ�ǽUȽD�ǽ�7ƽ��½j����G���i�����i���o����WV�����4����W��.$��;Ͻ�]�Ľ�NɽD2̽@�ͽC ν��ͽ~�˽sȽ}½⺽�ᱽf����|�������i���堽"f��:��b��TŽ�  �  @y������Dּ���|��h��}��U�J��� ����ʼ����f���1���#�λ?��v���~���޼���߈����o� �� �G�����A!�.�ͼ�k�����Be_�T�Cʻ��^�r|꺘Fκ�7��̭�����{Q�R芼*}��f�̼W켼z������ �jD)�,��a'������r6߼����WЊ�Kmj��h�����m髼	ڼ�������&��O,��_*�Pb"�1�����P>��n�ּj�� Ϛ��7y��@����ua�I!ֻse���w$���a��;���޾���缏��Q\�q_,�Ք=��kM�ǗZ�F5c�pLe��_�wDR��*?�ԩ)�v��;�����	�����P1��@L��Bf�xp{�2���{F���0���F��?@y�'Bl�}�^���P���B�� 4���%�hp���hG������=Y�%6)���;��HO���b���t�AH��Ë��֓�i���Р���o���V������K�������r�3h�b�f�&�p������@��CЛ��9�������H��>ø�ʶ��h�������d����d��_����䋽B��/�~��Xv���r�_t���{�'��T5���4���^��u;������𴷽.q��J�ƽC�̽�ѽaҽ��ϽlMɽ�`��ꆳ��§�O<���Ƙ�Ut��T���n������꽽xȽ�Ͻ�
ҽ�1ѽSMͽ�lǽ�����'��ܛ���٩�]С����"����ˊ��Ʌ��`���烽vT���8��)Д�&=��Vϥ��*��I?��t ����Ž
�̽�ҽ+lֽ��ֽ�@ӽV�˽�a��맵�ƻ��>����4��Z�������4��oQ��oʽ�ӽn�ٽ�`۽��ٽ�$ս�Ͻ�Ƚr����c������2���Ұ��?%���瓽)я�z���������i'���3���ѫ��j���  �  m�c�����B-ּ6d��� ��D6�r"D��4G�mK>�!�*�|��c���-���̅��;��j��5l�������5�^H��O�#FK�ـ<�&���漍���i���iA����������}�SW�:i�;cd&;"�:N�Ĺ ,T�KA߻��3��р�����u�ݼ/[	�)?$���<�zP��AZ�T�X���K��4�м�����Yż���P����A���!�d����1���I�{]X�$[�6QR�>@��T(����b�vָ��펼��U��q���̻���2�{�&���f�_m��2��m�P��f�������`��B�b�(���E�.,b��{���������܈��c��3Ik���O�?i6��?$�՜��e$�`�7��T��^u��C���T��� ������Vq������D��Vm��U�9?���+�)O�js�e\�h1�������<w���F�'���$���6�c�K�G�b��Q|�f܋�?����t��!���~��{��1�����jJ��ƒ������d���C��*݅�AY�������.���⿽A]ʽ
Ͻ�ͽ�Fǽ�#���1������ߐ���s��t���~���r��=i��4c��a��Cc�!�i�r�s��ŀ�刽����A��O������}V��=�ν۽�佫k齐��|�Ὅ)ֽ��ǽ~۸�)ܬ���������¼��a9����Ž�qԽ[���罋f�A�-)ܽ Bн^ý��B���q,�������T��#:������|dy�k�u���v��|�󳂽����ᐽٙ�M�������<��;�ɽ�׽���B뽹��,�����V׽��ȽC������8���^���˶�W�ý�ӽ8k�eb����������սǵȽ���9���Z���b�����N��~��z�����^���ъ��6���1��2t��$䨽�  �  =�A�3۟�������>��=^���r��oy��Gp�w1Y�̬8��6�o���¼�z���B̼aZ��� �$-E��Be�t�z��ɀ���x���b���B��2����}���i����%Vp��=	�
�/;�ȓ;R�;���;�8�;z?L;V:v,:��q�ovQ��V��5��ޕ�n�;���^���z�zQ��L�����|�!�a� �>��������(�ܼ��ڼ����.���:�9^���z�}��� ��)�}�$Nc� �@�Ʃ���;v���p����h��MG#�����9���9���)>"�����m����]�]y��AӼH�	���.���U��Z}�]4���0������D7�����@P��� u�5�U�?�%k6���=��T�ƛv�H͎�_,��L����� ��Ǭ�2˞�C���lw�[�T�n87�_��a���{��k�>tټ�sԼ��ּ׏�#e�����(��O'�|�>�@�Z�ڛ{��M���٣�h�����ƽ��ѽx6ս"1ѽnQƽ�ض�r���h��76��"���꒽�n��$���4.ƽ�l׽�H����Nc佀ڽ�	˽'���+�����\z���-���n�@]b��Z��tU��cT�ܽV��i\��ie�ƹq������[���/���k��Y���iǽ�\ڽ<�������� �C� �tn��Ԥ�$۽�_ɽ�亽ȗ����n���mnǽ��ؽ
������L� ��� �@�����\ܽ��ɽX���$J��Oi����4��W�|�֨r��Fl���i��Lj�ån�a�v�����̈�V����֞�����X⾽'�ѽn��]b��<� �������������A۽܇ʽ�(��˪���2��OŽ#
ս�J罸x��F�����=��98 ���R(�c�ͽ���@����۟����z��s_������������z��能F������Ç���/���  �  ?:�M���o���v�.��I\��n���U��7����������֞[���2����� ��?����X��E?�Oi����O#��M����Ր�#ۂ��3^��1�V��������\��ػ+��;�L�;���;�t�;S�;L��;�+�;��A;� �t���=�x=��ۅ�q�$��5S���~�F���o���������������`�T7��;��U��R�7e�q=3�:�[��
��S^���z��,���:������@�Y�A�+�c����	��b�^�}���e�M��O9�E��:7�;H�;	z�:Y�6�H��wٻ��9��+���s̼�!��8��h�Q������r���j���-���8�������A����o�݃U�zK�+/S��l������ݟ��ô��iĽ��˽ʽ@[���֭��k�����$Z���5�I��\��d�1�Ҽ�ǼxļpǼRм��߼������
�'���u8�A�X�s���p��<N���uŽSٽ�d�J.�8��4?ڽ�HȽ2���Ȱ��Y阽u���ҝ����;���ؽ��뽣���Rn��X������ؽC�½B(���e���݈�
�w�#1e��iX��}P���L�L��}N���S�
$\���g��w� 0�������\��yb����ν@/潾������(y������M���'���@׽��ƽ���R���?Ž
ս�7齀���~���������4�N�������ѽ�x��������� ��m��t�r��ri�/�c��ha��#b��e�DBm�qnx�!���厽L��������ý%�ڽ���ZJ�\�
���B��MH�F�����|�׽8_ɽV
ý�Žjsѽ�}�Rv��#��[�����D�&�	��| �뽫-Խа���
��Wߜ��0������P���$7}�v�x�e�w�6�y�T�~��΃�Q4��(��� ���  �  �=��o��z�	�a>��Yq��B��躜������h���
��%s�%rF��8�q�oi��'�
�Iy)���S��Ԁ��ڔ�=�������#���B:��sr�Gm?�y��1���F�\��2»����{�l;]!�;���;lP<�<�<���;�f�;�t8:
э�Z7�Q��ɨ���s0�ѳd�����H���j������E ��t���JCv���I�
�%�6V��<��"��oE�,]q�ӎ�H���}��a���7��������k�9R8�����8��>�Z���ۻ��\*�:�p6;q�c;��W;�f;��-:����������'��S��`�˼a����@�d�u�RǕ�����{��hȽx$ǽ�?��l)��ǔ�	����nd���X��Wa��|�pE���Z��B½w�ҽK�ڽ`�ؽC\̽ʞ��!����W���_�� 7�J��h����ݼc�ȼ�������N���bǼ�uּp�켄�����d?6�2�Y� ������f%��3н��������5��Kt�� ��~Խ����૽�������������o�˽�R������%��S�R������^ʽb����S��B҈�u�]�`�_2S��LK���G�~hG�T�I�bO��W��b�#�r�vN���ے��\��5���"�Խ���E���<�)��/l�����c������ཽoν�ĽS�ý`�̽�!޽�!��&*�c�������w����ؽ+	���٨�N���_���|�ļm�pd�I_���\��]�P<a��.h��Es��Ӂ��\���Ҝ�j����ǽ�ὃ����Z	�������E�����c��xYཚ�н��ɽ�ͽ�ٽ�)���������%���������+� �ٽ3n��䠬��ۛ��)�������>Px��Qt�<^s�Y7u�z�o;���������ٝ��  �  Uw?��������g'D�n�x��ݒ�aޡ���������Ғ�Ys{��eM�J%�c|
����&�[~/��[�("�������@��l ��(���AYy�X�D�������]�첼���@��(�;&�;�<�<H�<�j<f��;�`�;fk�:d�����6��m��� �w�4��k�i׎��뢽��������Ǝ�� ~��lP�G[+�|?�O��.(�N�K�y��X������ү�����������e�r�==��a	�����]�Z���Ի�ںh�:��N;j=z;�|m;�%0;�:�ĺ�@��|"��ֆ�U^̼0B���C��{�2N�����|Ľ��ͽ�r̽�5��d����z��5ă�ǩi� �]�	Pf�>������j����ƽpؽ�C��ݽ�	ѽ��������a����a���7��`�����^ڼm�ż����w!�������ļ�oӼgT����Q���5�	cZ����#l��\���ӽ?�꽱������ӧ��O�V'ؽ����?�������=蟽����������Ͻ2\�D/��rk������vI��:+�*�̽�B���/��-����`t��P_��Q�
�I��"F���E��}H�ۏM�DzU���`�-0q�qʃ��Ò��᥽a���A׽�򽅨�J��r�I�@������������-ѽ�ƽ��ŽK}ϽmT�����rl�2�������u�7��2���fڽ�s��u��I����懽�z��l��b���]�Ä[��6\��_�W�f���q��%��0����뜽0��HWɽ�j�����i�+������������k�tӽ�Z̽҂Ͻ�bܽ����z>�O��x��h�D��J*����۽}�½� ������𖎽�T���T~���v��r���q���s���x��k��7冽y`�������  �  �=��o��z�	�a>��Yq��B��躜������h���
��%s�%rF��8�q�oi��'�
�Iy)���S��Ԁ��ڔ�=�������#���B:��sr�Gm?�y��1���F�\��2»����{�l;]!�;���;lP<�<�<���;�f�;�t8:э�Z7� Q��ʨ���s0�ҳd�����H���j������F ��v���NCv���I��%�?V��<�&�"��oE�G]q�-ӎ�`���%}��0a���7��&���&�k��R8�9��t9����Z���ۻTr�[�:P�6;j�c;g/X;4�;	�/:hn���V���'�p7����˼/��Tq@�}�u�ƽ������r���_Ƚ�ǽ�8���#�������<kd���X��Ya���|�I���_��i½��ҽn�ڽ7�ؽ�e̽^�������a����_�7�������,ݼ��ȼ��� ��qO��7^Ǽ�kּ�u켻���u�!16��Y�B����v�����^�Ͻ�彔���t-���l������ӽ����ޫ�I�����A�������˽���X��}��N*�wX�J����⽃ʽ>���]���ڈ�� u�h�`��>S�WK�v�G��oG�5�I�
O��W���b�"�r�*O��Vܒ��\��b���;�Խ���J���<�,��2l�����c�������ཿoν�ĽT�ýa�̽�!޽�!��'*�c�������x����ؽ+	���٨�N���_���|�ļm�pd�I_���\��]�P<a��.h��Es��Ӂ��\���Ҝ�j����ǽ�ὃ����Z	�������E�����c��xYཚ�н��ɽ�ͽ�ٽ�)���������%���������+� �ٽ3n��䠬��ۛ��)�������>Px��Qt�<^s�Y7u�z�o;���������ٝ��  �  ?:�M���o���v�.��I\��n���U��7����������֞[���2����� ��?����X��E?�Oi����O#��M����Ր�#ۂ��3^��1�W��������\��ػ+��;�L�;���;�t�;S�;K��;�+�;��A; �t���=�y=��݅�r�$��5S���~�G���q���������������`�T7��;��U��R�Ve��=3�o�[��
���^���z��y���������d�Y�y�+�����U��[�^�	�����M�d^6���:�8;�.;C�:����G���ػ� 9��􍼮6̼� �]�7��g������o��Ta��SZ������+�������9����o�Q}U�K��2S��l�����$矽�ϴ��wĽ� ̽%%ʽ?m��魽!~�����;0Z���5�,��I��6�-Ӽ��Ǽ4ļUǼ!Iм��߼'|���
�����Y8���X�����^��^;���bŽ�ٽ�R��뽀�潈2ڽ1>Ƚ[��������昽�����ԝ����|����ؽ#������T������$�뽋�ؽ�ýT;���w����x�bLe���X�?�P��L�7L�4�N���S�+\��g���w�{1��p���w]���b����ν_/�������/y����#��T���-���@׽��ƽ���S���AŽ
ս�7齁���~���������4�N�������ѽ�x��������� ��m��t�r��ri�/�c��ha��#b��e�DBm�qnx�!���厽L��������ý%�ڽ���ZJ�\�
���B��MH�F�����|�׽8_ɽV
ý�Žjsѽ�}�Rv��#��[�����D�&�	��| �뽫-Խа���
��Wߜ��0������P���$7}�v�x�e�w�6�y�T�~��΃�Q4��(��� ���  �  =�A�3۟�������>��=^���r��oy��Gp�w1Y�̬8��6�o���¼�z���B̼aZ��� �$-E��Be�t�z��ɀ���x���b���B��2����}���i����&Vp��=	�	�/;�ȓ;Q�;���;�8�;w?L;�U:|,:��q�qvQ��V��7�����p�;���^���z�|Q��O�����|�*�a��>����߄��\�ܼ��ڼL���g���:�r9^��z��}��#��;�}�yOc���@�p����~x����p����V���#�rN�
��9,��9����� �0٫��5��0]��*����Ҽ�	��O.��U��&}����H���w���"��t��=A��o	u�ƝU��?�*i6�L�=���T���v��ڎ�=���#���$��8���ଽN垽g���dCw��*U��d7�
��r������%A�h�ټ1�Լ�ּ��QJ񼩘���T.'�$~>�Z�0k{��3��J�������w�ƽ�lѽZսoѽ�?ƽʶ�f����a���2��^�����v��İ��i=ƽN׽^����*}佦9ڽ�%˽޸��-0���+��F���QY�Y�n�b��2Z�C�U��wT��V�]v\��se�8�q�Q����]���0���l������iǽ]ڽ^�������� �L� ��n��ߤ콇$۽�_ɽ�亽̗����p���nnǽ��ؽ������M� ��� �A�����\ܽ��ɽY���$J��Oi����4��W�|�֨r��Fl���i��Lj�ån�a�v�����̈�V����֞�����X⾽'�ѽn��]b��<� �������������A۽܇ʽ�(��˪���2��OŽ#
ս�J罸x��F�����=��98 ���R(�c�ͽ���@����۟����z��s_������������z��能F������Ç���/���  �  m�c�����B-ּ6d��� ��D6�r"D��4G�mK>�!�*�|��c���-���̅��;��j��5l�������5�^H��O�#FK�ـ<�&���漍���i���iA���������
�}�PW�:g�;`d&;�!�:o�Ĺ,T�OA߻��3��р�����x�ݼ1[	�,?$���<�}P��AZ�Z�X���K��4�޼�����Yż�������B��"����L�1�i�I�D^X�' [��RR��?@��V(����f�5ٸ����U��f�n�̻ق�bf1�>�%��ze�ʣ��!&��TP�x��X\�������"�(���E���a��z��z��<���OÈ��M���$k�u�O�0U6�X4$�j��Pl$���7�F�T�9u�+X���l�����ة��V����5���d����m��BU��:?���+�;y����v��U�����n�eg��6� ����#���6�ߛK���b��|������ܙ��S������S��������8��T������&`���C��#ⅽ�b��� �[A�����bwʽ58Ͻ��ͽ�gǽ�E���S�����t���A���J݆���~�w�r��ai��Rc��8a��Wc��i���s�Iʀ�f舽#��vC��E���o���V��~�ν6۽���k齧�轍�὚)ֽ��ǽ�۸�.ܬ���������ļ��c9����Ž�qԽ\���罌f�A�-)ܽ Bн^ý��C���q,�������T��#:������|dy�k�u���v��|�󳂽����ᐽٙ�M�������<��;�ɽ�׽���B뽹��,�����V׽��ȽC������8���^���˶�W�ý�ӽ8k�eb����������սǵȽ���9���Z���b�����N��~��z�����^���ъ��6���1��2t��$䨽�  �  @y������Dּ���|��h��}��U�J��� ����ʼ����f���1���#�λ?��v���~���޼���߈����o� �� �G�����A!�.�ͼ�k�����Be_�T�Cʻ��^�v|꺝Fκ�7��̭�����{Q�S芼,}��h�̼
W켾z������ �nD)�
,��a'�������6߼田��Њ��mj�kh����	꫼�	ڼ��B���&�Q,�)a*�d"�)��̪�8B��h�ּ���M͚��+y�l@�&a�4��v�ջް��%$��a�镼%��.K缌T�~�,�eN=��$M�DRZ���b��e�b_��R�]?�F�)�B��{.�٪�G�	����`k1�eL��of�@�{� ���g��qS��uj����y�ۇl���^���P���B�?04���%�B��L0�"R�i����{F��)�4�;�fO�Pb�b�t��&������(�������%����ѣ�9{��(:��h��B8������:�r���g�	�f�+�p�3����P���䛽�R���ֱ��h��A渽������Ԭ�������������Ғ������Y����~��zv�k�r��ut���{��-��d:��i8��sa�� =�����������q����ƽ}�̽�ѽ5aҽ��Ͻ�Mɽ�`�������§�V<���Ƙ�Xt��T���n������꽽yȽ�Ͻ�
ҽ�1ѽSMͽ�lǽ�����'��ܛ���٩�]С����"����ˊ��Ʌ��`���烽vT���8��)Д�&=��Vϥ��*��I?��t ����Ž
�̽�ҽ+lֽ��ֽ�@ӽV�˽�a��맵�ƻ��>����4��Z�������4��oQ��oʽ�ӽn�ٽ�`۽��ٽ�$ս�Ͻ�Ƚr����c������2���Ұ��?%���瓽)я�z���������i'���3���ѫ��j���  �  I�ҼR.伜�����i������~�u�ټ1
¼ r��p�{�*12�����ї�Is���%���	�voP�����ᵼ<7ּ����(
��6�n[��W�v�������jԼ)����T��W�S�=��x��ݻ%���>��e������]�ϼ�p��t�%�	�����?�������`�����6޼Ϥ��	t����a�n�'�!���#���"�w�Z�S������ �ڼUZ��<�����&(�-&�TJ�I�8a����k�޼1G��K���a�x�M��j=���N�Y(�����ˣҼgm ��t���&�tA3���;�C�@�Y�C��5D�E7B���<�0�3���&�6���2�a!２�ۼ�yּ2p�ߪ������&���<�tdP�|�_�8�j��r�0v��w��w��t��n��kd�I�V�� F��f5�V8'�pe�����#�ִ1�<6E��F[��p��ၽm6��PX�������g������Ǔ� ��=����j��5G���t���c��_V���N�Z�N���V�&Gf�&�z��t��#4��Uh���}���n��蘫��q���E��S��	����A��5��4���)��?v���k��S�������y��iF��=4��̥�e���Lɷ�󶽽%����ý�ZĽ-Ľ"�½����[�������>Ǫ�����ٗ�d����X�����ˏ��ɖ��ٟ�o����j��v���tϾ�/½��ýXTĽ��ýY½�9���&��'���>���Ơ�.����S�����/���`/��tӚ�VJ�����(���q���ý�!ƽ�ǽUȽD�ǽ�7ƽ��½j����G���i�����i���o����WV�����4����W��.$��;Ͻ�]�Ľ�NɽD2̽@�ͽC ν��ͽ~�˽sȽ}½⺽�ᱽf����|�������i���堽"f��:��b��TŽ�  �  �t����-[�2��>���8ؼ����&��qV|��F<�����+��m1��N�=:���://�8�$�w۷�#X�ASb�`O���T��fZԼ��󼖻�!��h���
$�� ����e����ټ+��#���X���P�	s�.`���]ʼ2�����g"���)��)�K�"�4���
�������ؼ*���ꂙ�(�p�3�/�ن�
���xD�yF?������?�3)��i����h��S�ռ���-�������"�q�*�"�,�n{'�+l��T���⼄a�����Eˎ���4/��j�伴���I)�F@�v�P�+8X�� X�ȦQ�L\G��;��-�aP ��k�$%����_Ѽ�
s���^���K���˼�g����%��.�QFA��S��8d���t������Ǉ��e��+�������d����Wm���W���D�'8��(5��<�wYN��f��ˀ��x��Bw��T�������h���{ѓ��B���s�����p�Mob�9ET���G��>��/9��:�KA�GjM���]���p�jK��T����.�����˩��mݮ�n7���绽3뾽ub���������&��'󝽇�������e���ޖ����������MŽIoͽѽ�ѽ;.ν��Ƚ���-F������K���Qi��i��������[�����(����p��/�����h����ј�R7��[q���e��M%��c�����ǽU�ͽ$�ѽ��ҽ�Ͻ��Ƚ�����̲��~���Ğ�3X��X"�����᪽9ݶ�#�½U�̽�8ӽ4�ս�oԽOJн^Sʽ�pý�-��@����
��N������H��x���+5���[���v���j������{����#����������7��Ž��̽
�ӽ�hٽ`�ܽlܽ;ؽ<н\~Ž�ǹ�z;���姽�D���짽�f��;K���ƽ)$ҽ۽�  �  �*C��@�4v3����&��N�ּ���;�o�+v�[����b���:\�m;y��;8ݫ;��;�H*;��0��+q�������L��ґ��y¼Fc��'��x0��E�8Q��9R��CG�"�1�����}��������e�������e�ݼ�����)�MuC�b:T��jY���R�	`B�c+��V��,񼼦����R�g
�&H��&����8�:`�:|\9i���e������J�.��>㷼��輗��"!)��
A�!�R�O�[���X���J�]�3���2���P:Ӽ(����˼���:���5�ޝV��Jq�Ѐ��؂��~�%-m� �V�$�=�(�%����P����ּ����̣�n_�������ꊼ���g�������4�/��UZ��1.�fRG�S�b���~���nؘ���Z⣽$񠽹���	,���|���c��iS���N�D�W���l�hX��˕�mꤽy%��Hȵ��L��d[��Nv���k���،��‽GLl� �Y���I��p<�b�1���*��(�{�)��/�7:��"H��Y�}il� ꀽ����ƙ��ç�a����ý��νa�ս, ׽�ҽ�lɽ�׼�*���¤�x��������������\��%#н�ݽ�d�2H齅&潎�ݽ�{ҽ�^Ž ��g����_���g��"������	��"�v��@r���q��v��d~� $��%������A垽s���=]��פýK�нv�ܽ��� 꽈�轵�b�Խ�]ƽ�"������n��"a���ï��$���˽��ٽM]彰��j�콚��E1޽Sҽ�Ž�A��D}�����YΘ�'ʐ�� �����D������׀��냽�������[×� ����q��a4���&Ľ~�ѽ�߽kc��|���!#����ڽ�X̽����.����@��B����徽>�̽�۽C������  �  �Nu��1o���Z�xq<�%u���,2��fL��һ�ͺ��;!�;n��;��<�<�.�;h��;�Jl;]��9����;��Q��~�ür#��R,���P�qgn��p��sT��0�x���_��!>����n����Լ�hμ_�_�1�H4U���s�/\��^b���\���f��E��� �	���򬴼w�v�	G�����y����a�:�fW;�b�;�;n�`;[M�:�2T��ы����n�j��ǭ���;���B��]d���~��:�������/{��y_�"�=�o#�������X��'���5�I�\�r������*噽�Ś�����U ���m��pI�N)'�*��bo߼'η��晼*���+�m���a�- e�̐v��;��7R���i��¹�N�	��$�/E�`�i��X�����A/��V����伽v���6��mB���\�����:�m��yg�	�q��<���ږ��a���.��Oɽ�ν�o̽��½M���Т��ؐ��$���yc��	L���9�KZ,�E�"�-k�x������7#��[,��9�]=I�X,]��hu��;���.��1������.�ӽ�e�T���l�޵�5rཕѽ~���yF��q��b&�� �������>$ӽp��`���	���[� �]s���G�5�߽�ͽ�~��Y������S��}���(A|��$q�%�i�@�e���e���h���o��sz��d��q���E�������1��©ʽ��ݽȵ������O��� ��`�����jٽ�0Ƚj˺��򳽈���꽽��̽��޽�_�a��K��XX�'������Foݽ��ʽ�	���0��{ݛ�e��w���5��m1{��u�2�s��#u�N>z�<|�����=������v���u��e�ǽ<�ڽb_�{���������"������^]޽�,ν&�½i�����½Z�ͽ�4޽i�𽢜 �����  �  ����V���;�4QY���,��r������kC�����D$:���; l�;��< �$<P'<Ջ<�<9^�;z�.;B���%�����ͩμ�����B��Lo�@��"���kR��Pԑ�8r��F+`�9a7�����X��������
���(��P�y3z�����A��.������r����_�:�1�{�����m�f�k��S��|�:��w;���;���;X��;|��;�q�;�8�:0����޻�*Y�K���[���o�,�>&[�¹������Ѽ���y���a��Dc����]��7��}��Ea�J�*��P��}��ܔ��1���¯�+���]
���Ж����C�W��m-�y_��Լ!ꦼ�s��1b��qI�\Y@���D�9V�0�s����������Ӽ����J"�kH�p�t�/������ ���̽��ҽ��Ͻ��Ľ�+������[ƍ�������{�Q���͗�������޻��н��޽�佩Ὥ
ս��½묽D�������6a�I~E���0��"�c�����њ������"�#��/���?��T�"�o��ӈ�8��%���S̽g!�.D��/Y�}<�ɔ �����%⽺5Ͻ;h��0��Ϡ�����<4ν��⽽x���>�9�
����+>��� �v��ʸս����n��8���Q���݀��xr�4�g�]a���]� {]�[`�D�f�x�p�1G�������z��� =����ҽH��N��������|#�u������H�սAƽ�a������u�ɽ��ڽU�ｩ��M�	����I����ߙ��3齹ҽ
:��( ���2��5댽�у���z�*r��,m�ȅk���l��xq��y�MÂ��-��艖��O��x���ͽ=K�8Z�����^��Ʒ�U�[
���"���ڽ�ͽɽ�lͽ�Fڽ)�����
�|U��  �  *��������U�� n�X<�)��^x��ҧE�`	�� E�:dN�;-E<�=)<="7<�%9<@�/<�<b��;J~;~{q����҃��(ڼ���G%S����,���$��G\���^��`����w��J�[�$����G�	�����p:�g�e�l��������/����������@t����r�El?�3��"p���d���ڻf� �#;�~�;���;��;:��;E��;���;&�:;i�J��bû�_U�E��AZ���9��m��q��6�������d��Q�������s�c�I��!*�ڑ�%*!�-r:�62c�����tС�����M���̔��X��p������4Zc�֫3��$
��YѼ�@���"y�6PM��5���-��>3��-D���`�]���^	��˼�4 ���"���L��}�/s�������ʽ��ڽ��(�޽iAҽ�;��%��� 9�����6ф�Ƿ���֙�t�����ǽd�ݽ�1�hx�lZ���gͽ��������}n��n�a��C�I�,�[��pu����C)��v�c�����E�*�$�:�/Q�� n�䒉������x��ycԽe�h��Ť���
�A��� �����ؽ�{ǽ�S��Ŗ��)�Ž�׽����|��F�UE��O�61�����9��sܽ��½�	��2Ә�a����}�SOm���b�?T\��7Y�Y Y�e�[�d�a�ˀk���z�m������,Z����qHٽ�K�ʇ�(�� ��oZ�;�K8��S����޽�ͽ|QŽ+�ƽ-�ѽA:�!����_����]�U�������ģ���׽m_���詽i����*\��x�u��$m�K�h�*g��dh��l�)bt��3������s/��e������	�ѽ��뽻��@��p���6��h����-����4^��$ս��Ͻb�Խ���x����wo�����  �  ��!��4�������nн/ӣ��av���1�J���dk����Q�5��������`�u:K��^����Ȼc����z�2I��f����G�Lg��������߽���xn�1�"�i%��0��\����d�ֽ@���0��N�������'Ƚ��e
���,	%�t�&���������PF˽:����Jq��0��W��*x��ory�.E3��E��+��a�� �d�+�{�m�!�����D;)�(h��@���Žl?�,�����F&���%�k���:��{��d�Ͻ����S)���ک�`n���Q�������~(�R�0��0�=�&��'�^p���ֽ�6���#��{4X��[,�PL����w�ټ�ϼ��μIټ�)�L����=��.h��6���=���wܽp��A<���.���<���B�ݗ?��[4��]#��>������F潲޽�B罰% ��X�_�&�;w9��F�ĮK�I�G��X;�,�(��]�����޽ҽ�㰽%@��>���%�i�ՉX���N�"]K�DM�ެS�}_��Pq�m��A���Ʈ�-3ͽ�y���K�%�#�;���M��zY���\�n3W�NJ�=b8��%�P�
�����?���!���4���H���Y�@�c�:�e�:^�0O���:��$�-��3'��\�ս���T2���՛�
쒽q��g���ф���Ќ� ԑ�|-��Zڦ�*����ѽ�3���s�!��8��L� �\��	e���d���[�~�K��8��%��(�ִ����*�-!*�ѕ=��P�,e_�G�f�NPe�.[�.J��5�3��3�	�Op�н�湽�^��������������� ������`⛽.٥�~��A�Ƚ>�*��z���-�}D���W�?Pe�U	k���g�<?\�Q�J�c7�v�%�P�լ����+�$�|%6�R�I�P
\���h��  �  A�x��^���T��-M˽�����s���0��c��#^���[�.d�V���t�����s�|Ֆ�n�ݻ#^*��Y����¼�T�EeF��h���*��ͨڽ�3�{k�EE��� ���m������Gѽ7���J-���������	ý�N罶�����Z� �
"�f��g����ǽx�����n�l0�}����ᵼ�⁼��=����=u��C���)S�M6�Cx��������j5)���e�Ɨ�6m��M��!
��X�{�!��>!�����|	�&*�ʽ�l���M��_�)���r�ڽ�^�N���5$��O,���+��"���������0ӽ^��vW����X�	.�������e+߼|#Լ��Ӽ�޼�H������T ?��#i�q֏�N���(mٽcs�m��+��j8��>��#;�U@0�e��OB�.��F ⽸=ڽW/�7��� s��N#��r5��>B�3.G��UC�o{7���%�-��Ͼ���ѽ0u����������2al��,[���Q��M��O�,V��	b�r�s�����Y��� ���t̽�p�����"��)8�U�I��U��6X���R�d)F��4� #�+��&���	���P@�k�1��2E�m�U��~_�-a�x Z�A�K��8��z"�Y�����Nyս;Ƽ�EL������=�����������ȋ�����%��z�����������ѽ��z�
���,5�kI�2^X���`��/`�CiW��H�T5�h#������������We'�F:���L�q[��Eb�U�`��W�ŹF��^2����X����н����6����T��g���⓽C[��}S��Xז��4��@�������pɽj��+f�]��{~+���@�A�S�� a�X�f��Rc��&X��VG�g4��:#�;������l,"��93�6uF���W�
=d��  �  �g����P�����_���r��z.k���/�g{��"g��,�|�1�/��0��ǒû�Ʒ�G8ֻ5��ؕL�������ϼ~t�+D�����y�Ъ̽h��E����O)�����R���㽭n��-���c��������������C�ս�����
����k���F:�n��Y���-A��;i�
f1� ���ż�ᒼɫ_���2�Rg����L�.��X�5��5E��;��o�*�Hja�+��������ܽg% ���� ���������kJܽ�ӻ�X(��AM���˚��J��2�˽g0�
	
� ����\Q��P��?	����ɽ⥽�冽eW[�~f4�U��r'���8伽g�x��6��I���'��F�}vm��������ѽ�n�����Xd �DZ,�Zb1��.�I�$�a��<��q/�dOֽq=Ͻ��׽��0<�mu��*���5�r�:��<7�K�,�0���
�\��
7ͽ�	��[������4�t�u�c�"�Y��U�(W���]�w%j�8|�������Uv��;9˽͋��F������.�U�>���H��uK���F��;��c+����_�'>�T���
�����(�4�:��I���R�kwT�I8N�eSA�� 0�E����	�1?��սsd��6��q^��tw��HŒ�1⏽5�����-[��'���`૽4}��xNҽ���x�P��c-��?��L��S�Z�S��yK��q=�U,�~������(��	��v�i����0��A���N��U��pT�O�K��7=�=+���������+ҽ�۽���������9��~ݗ�+;��>���욽Bv���P���#���˽<�㽰� ��!��K%��k8�(I���T���Y���V�h�L��?=���+��B��L�+3�����X��*� �<��L�B�W��  �  9���*e���1�}u˽�V������6�d�Lz3�6�
��Ӽ	���Jo���8�/d��8��g#��xL������߲��=�c���E�Q�y�Z���N����ؽ��� ����03������ǽ ԩ�Lܐ�W���;�}�]-��Pʞ�(����ٽn)�q}����s����)�˽���nɎ��f�(�7��9�H1�u��.��I�l��BS���Q�Qh����
ǭ���ܼj��L&2���_��ኽ*񨽬�ǽ	e你:������-�z����޽�����ॽY�I������\H���Ŵ��Խ��a��3��g��:������۽�w��Ŭ���R��~Wd��VB���'��d��8�X) ��u��m}������ ���7��T���x�p⑽�b��D�Ƚ�轥��N_�q�����5I����������bֽy�ĽZ���8ƽO�ٽ�����
�fe��#�j(���%����,�����Mʽ����Q/��1y���p��Ԁs��_h�Uc�1rd�G�k��x� ��5t��
��%����˽���k�������!�i�.���6���8�\4���*��-�&��w�T"�����������T��RH+�kN8�Gh@�"B�:Q=�;�2��%����(A�*���0ٽ]�Ž�ܵ�l���RF�����𻖽<��*P������ާ�ڻ����½�ս��U��>��"�8!1�c<��A�^A�%�9���-����d���q�_���� ������#���1��=��C��sB�4�;���/��\!�3���6�Ns콷�ֽ�Ľr�������ڣ�w�����'��&L��Cb��Ys������Ndѽ��� ����� 1���,�7.:�#�C�.[G��D���;� S.�8c�X��2d�1�� ��	"������-���;�Q�E��  �   �ѽ�SϽ�Ľnj��'t��Nڇ�g�f���A�Z� �`��<8Լ@驼�����Zm���c���x��խ��Q�͗�k�.�-�Q�E�x�Nӑ��	�� ��@νP&ؽ��ؽx�Ͻ[����I��x⍽��r��Y�.UU�of������������P�ʽףؽ��ܽ�׽�.ɽ��sO��Y���bcm��FI�9)���輷⿼����Y꒼�B⟼�\���"��
	���$�r�D�5h��ʇ��5��-�����ƽ�սC�ܽ�ڽ��ͽ�9��x���؋�ډu���e�i�k�"���k����e��ޤν����=�v��z7�<Kܽ��Ƚdг��f��(Ȍ�%�x�Z�[�V�B�"F.�����0���0�-0&�3�9��-R�p�n�����	m��Z����½"%ٽ�?�X(�1��8�	�s1����d��V�ҽ�����L��Mʪ�@/��w���9*ٽ<��#������(�\�z	��v�9b���,߽7&˽�$���H��Zy������A�����x���x��T��󇽑������'���HB����ѽC��-��ȅ	��_�!E�ں"��#����Ek�Oz�s�yJｗJ��~�O�v ��`�2�S$�7+�g-�1�*�ǫ#����o�[:� *��P�ὦ�ѽ�ýi����v���������Ġ��B��,�������n#Ͻ�߽���Z��O��A"�k�)�\1-��+���%��s��B��k�Ӗ��YK��콮���ed�ֶ�3��%o(���-�>.���)���!��������?�񽲘ཛTѽ��ý𖸽��������?��K�������vԵ�3����ͽ��ܽ���D ��
����\� �x*��`0��g2��t/�O�'�B������p�Ul��I������J����]��o=(��0��  �  "���ܪ�,���5p��"Г��8����x�`�7`F�.�+�i(���Aɼ{%��d����ȶ���ռ�Q�и���7��7S�|�m�8������M���䦽u����}���ۯ�7����X��u��ZBb�&B��i.�`	+�1�8�ëT�2z����ȥ��z,��2��᬴�Wɮ�Z�����,��j�F�j�P��4�g��4���߼P˼�ʼ�6ܼ���<��+1�NML�5�f�����>���3��e����s���������Q۰�
���!t��(�����a���G��<�w�A�~X��{������2��Iǽɗ̽=f˽T0Ž/ỽb��fѥ��@���F���ہ���j�^KS���?�,3��X/���5��.E��t\�˘x�Ig��{z��������_�ýH�н�Eܽ;���r뽑n�}��-ؽ�ǽ�t��B���������DF������*�����нS��<�������Y9 �����������ȣ߽Խ�RȽ'����l4�������6��p>����������\�������G½6ѽvu߽[�Y<���w�p7	�������\�E�w$�Z����4�q�ֽ�jν�'ν�3ֽ�_�w��������t�,���e��t�h�� ��m���c��z~�� 2׽Ŭɽ�����P���"��fˮ��T�����u�ǽ*ս9��(4�a�����9�
������>�����n ��[����c�����Sݽֽ4׽���Ƒ����j���7��$�2��\[�(P����ǧ��!��?w�_?彨�׽
˽��7t��1���ض��6���hǽ�Խ��A�� S��!�*f���6�����x��C�#������)W��-�彩��T�佭��5,��6�������  �  :-����������ȓ�{��۾���F���ψ��}�'zc�<&E�£&�����B��,D�Y# ��Q�d�0���P���o��儽ѡ���3k��6晽 ᙽ�:��`E���1�������i��6K��-�F�Z�Q���P��"�9@�+`��>~�����c����C���:���N���杽bƛ�50��6^������k�EL�7.��g�z��z-�r(�L�*��UH��g��?��:܍�"��ᚽC<���ޝ��������!���қ���>����h�pK��0�n��-��}���+��NH���j��T��{���y�����?೽1����������0j������Gx�����8F���́�|�i�_8X��R��Y�D}l�&���yЕ��������v½?ʽ;Ͻ��ѽ��ҽ�ҽ�PϽZ�ɽ���h��3䦽u�����j�����-���t&���6���j���O½�н�6ܽ���U�ޕ꽡6��A꽍*�{*���׽m˽Y'���*������/���Ӡ�!S��D󻽭Mͽ��ݽ�2�h���!��&1��I�����2�K� ��R��E����b�׽�_ʽ���!����߹�*f���a̽��۽��9[�����<E	��*����6(����c���M
� G�T� �ߛ򽫽⽽�ӽ��ǽ�����Y���Wƽ��ѽ%��6R����R�E}	����J����yX�n�O�	��i�M��j����ལgҽ�jǽ����N�½.ʽ�gֽ\�����S���\����E�'���8���y(����� ������սF˽R�ƽ��Ƚѽ�޽%��M���e��RK�=��/�<�y{����is�*~����|� 
�����*ٽ��Ͻۤ̽��Ͻ�ٽ���԰��1���	��  �  (?]��v�5����'���J��$��s�������ɢ�T�������J]�+�;���%�����*���D��Ui��ň����ű�������Z��������ڗ��#�����jlg�azM�M�2���������ټoü 㿼��ϼXT�4��Y*��F��Ta�.p{�1I������vP����������*_���u��䧽W����L���b��(C�֜1�M�0��K@�N�]��ၽZd�����w:���ֵ����,3��h/��g�������"6�M_f���L���2��}������u伊�f��}��19��EX� �w���C�������*���z��a�ʽumѽl�ҽQͽ%���U+�������������z����\'���m��ܱ���@ɽX�ٽ�T�:���W�p޽&Խ�ɽZ|��p�����������"}������:o�
�c��a�-Di��?z��7��퀗�#��������ý�lѽ�޽U����`����3�S������/�ޟܽy+ʽ�t��S���W���Qɵ��8ĽW�׽0R�r �C��?�����5�
�D����@+�����ὒ�ս��ɽF)���������������6������'��`�ý7�ѽ�/�B����&��K
��#��;����I��v��Mk�|;
�r �|���ݽpս7�Խ�eܽV8뽕;�����DL�����`����N<�:K�ӓ
�8��K����8��⽄lսKXȽ�輽ʄ���`����������;��ˇ̽,-ڽ-�v���rC�P��j��Wp��E��I�������<a�g�	�����M����&�ڽ�Wݽ�������o�Q�����������Q��r�wE�ۅ����y�x:����轧�۽zϽ
�Ľ0���=��)���A�Ľ�Ͻu�ܽ�w꽙\���  �  C�?�1f��&��t_���ӳ�q�Ž:ѽ�ӽ�̽r�������{:����m�2�Q�h�I���W��x�`��������½|(ҽؽ�Խ�|ǽF���ğ��8��`l���G��'��f
�������ӛ�����F�����<���>ռ�{�![�(�=��ma�y��7������sĽ�`Խ��ܽ�۽��н�m���I��- ����r��v\��2[�1o��_���P�������νU�ڽ�ܽ�Wս�!ƽ  ��FN�������f��D���%�c���Q�ɼ�e���Э�����U�ϼ��������0�XQ��{u�󖎽�9��(����ѽG�彤^������v������d�ս%������]�����ൖ�����cH����ֽ���m�[��������M��k߽<$ʽ�͵�
f���#��������q�@�]��O��F��E�<�L�d�Z�,�n�������� ���+��0ɽZ�޽�k�������!��	�-��-�
��=����ZӽY�ƽA�ý��˽N�ݽ�@��~Z�#�f����5[�k�e��ok������éѽ �½������c�����_@�����䌞��X���氽�����<̽��ܽ���98��������!�#�(��-�#o,�s�&��������ֺ�����n��#��GR��R����Q�%�O�+�d�,�I0)���!�������.&�ٗ��޽�:Ͻj��ӗ�����w���	`������`T������6h���ƽ��Խ�+�<�����T�h���%���,�Rv/��T-�=h&�@��1����?K�������T �/�
��}��`#�3f,�U1��0�d�+��D#�����"����������]�Խ��ǽ��܀�����KR���O���괽���]�Ƚ�_ֽ����  �  )�1���d�y��eƮ��[ͽ�S�3���_��������b��ƽ�����ۤ{�c�q�XK��Z���V��"�Ͻ+���Y��^� �zR���e�=�̽��O����g��7��
�-����,���;�]�+�A�E>�J�R�T)�My��6�ϼ#g��[*�\`W��J���;��I�ý���g!��Ϸ�_�3���b�⽊�Ž����=������m߁���������½��߽W���������#����㽛�ƽS���hĉ�'\^�6�1��t��8⼲ķ�����m≼�셼�̎��K����ż�n󼒠�.&:���d�̋�}਽�Ƚ܅�܍�L�n&��� 	����P�ܽ2���A*��p%���_���#���YؽD���!�
�q+�����h��	���8��]ҽO⵽E�������@p�]�V�MD�8���1�_�1��7��D��
V�R�m��녽4N��.r����Ƚ�7����Fg����?L(��#+��{'�+�����1��W��T۽��׽A@ὦ�����	������'��W1���4��]1��X(�P\�i��oi���ཕ�ɽR��c���T���}�������*��������Y���٣��6��f���c�ҽ�s�,�L��� �tH/���:�JaA�p�A�Pc;���/��!��F��I�U������L'�x���1��-��:��@�(SA�Pg;��O0���!��y��~��:�H�սQ�½��2���k��ߡ��O��?���f6������u8��$ָ���Ƚ��ܽr����Q����hJ'��@5�Ԃ?�!>D��zB��w:�8�-����j���������*���@(��6�O:A��&F���D���<�X�0�;�!�3H����h��GٽȽ�����6���䨽 �����1Ǥ�xo����[���rmɽ��ڽ�  �  ��.�{�k�󝙽�7�� �����p�o'������bb��A.��LN��+���Z<��hg��йʽ[��@_�N���^�a����Q���罽�=���.l�&�2��T�N���������Q��
#���
������j�A���櫯���n�!��=W�=񋽗ð�Ci׽j����X�u��ۜ���u�Ὄ����^��>���l����⠽�]��tݽ1��rd����z��*��+�۽����6��ʈ_�~&*�� ��7ü�񗼺�x�{\���V��ch����[����Ӽ���5.�"(_�<���@ְ�Ǯ׽�������/��$��3#��j�1�f���`0׽�^��4ж�8�����н���/
�K[�'(��.�l,���"����|�@ݽ$��T���o�a���F�}L4�
)���#�}]$��**�rX5�#EF���]�9c}��"���嬽�9̽,o�O������.��9���=�ĥ9���.�),��W��z��X��z'轱�� �����(���8�ʑC�y�F�d|B��7���&�\����z�⽄�ƽ���N�������}���0�������Ȉ�Af��@���4����+���Ѹ�Yν&X�����V�i�*�϶<��K��kS�k(T�.)M�_�?���.�c��%������z���)��ڬ,�(�=�V�K��dS�LS���K��>��V,�4%������콘�ѽ�[��/���o��Ye���w��/L��^ȑ�j9䚽��������½��ٽ5_���=�@2�#t2��C�4�P� �V���T�\�K��	=�u�+����J��PL
�
����Y%�Ά6��G��FS�N�X��KV�E�L��:=�b�*�n��W���E�UԽ����=z���-��`\��p���T���Ν�~����	��;��� ½�ս�  �  E�/��t�_��1jͽ����B���2(�%���8�֓����ѽ+���6�X���H.���|����۽������v ��Z�} ������	ʽ⮟���r��q2��P�����Ny���/�4w��
׻٠ѻH���m ���_�����qj㼲��u�Z��q���ƺ��1�^}�I��>!��O"�w��%R�Q���Tν� ���鞽���k��jbʽj;�bL
�cd�E�!��!���{s	���꽭����<����c�Fu(�����0⳼BJ���X���<�b�8��<J��p�喼xü$3 �'Q)��^�����Wٷ�;Y㽀��*m��*�D1���/��3&��|����彔~̽�����Ƚb޽ ����&&�
j4�8�:��e8���-����cV�3�:���O㜽�ꁽ�I[�@�>���+��� �h����g"��;-�`�=��U�j�v��F��9���TgнW����Q��'�p�9�&F�eJ��F��:���(�����w�=����O���'�����;�2�ZD��P���S��fN�X�A�@;/��d�����彠�ƽ����t����Ԑ�//���������.ׄ��X���Z��_V���!������ "ͽo�N���U��2�[SF�Q}V��_���`��BY�q�J��8�n`%��9�4��k�����O#�>�5��|H�v�W��`�7	`�dW���G���3�j���	����y�н�y���A���*���1��Vu��@j�� ⍽�ᐽ淪��֟�[���8���Yٽ�;�������$��:��N��\\��?c��|a��W��dG�X�4���"�K��K��T�ε��
-�9*@��>R�}�_�ele�/�b�]�W��bF�|�1�t;��B�Q<�"�ҽҟ��l_���棽�8��n����u���ޙ��ٝ�bĤ�L_������o�ӽ�  �  ��0�,�w��V���Rҽ�\������p�ٯ"�`���=�o�����׽s��E��ʒ���_��Yq��P��a�����!�m�$����������	�νߘ��.�u�T3�����㮼oo�p[%�*�{�»�f��L�߻;��YuU������+༛?��g\�u������a�뽹�
���-�%���&�b��+�#9��n�ӽ�����ߢ�V⡽[ӱ��Ͻ���6�����D&��#&��4�;�z����ý:�����e��o(����i���6��7�M���2��%/��h@��f�����O���&���(�E _�}ّ�3���Ƕ��
�V&�\S.�K�5�qO4��`*�J)�t$���пн��Ž�̽:�����u/��s*�R�8�pN?���<�-�1�g( ���
���ۚ��Z���靁��zY�R1<�V1)��A�����:������*��=;��9S���t�>㐽���z)ҽ�/��j���*�{�=�:zJ��N�*lJ��
>�r,�Gb����_J�������{��#���!��l6�XsH�otT�MX�3�R��KE��N2�[�����i�+ǽ^&��������ه�����n��ᎃ�����������'괽��̽Z�뽯���;��4���I�'�Z�tUd��]e���]���N��b;�m(�Pw������h���%���8��FL��[�_�d���d���[�K�8�6��h ���
�q�ｸ�н?������Cݚ������+��b&������2����U������E�������ٽa������,'�ϝ=���Q���`���g��e�R�[��K�2�7��P%�@������X�
�4�/�K�C��5V���c���i�:�f���[�l�I�U84�e��8	����OWҽ����X&��w����雽aD���2��l�������Pr��`!�����(1ӽ�  �  E�/��t�_��1jͽ����B���2(�%���8�֓����ѽ+���6�X���H.���|����۽������v ��Z�} ������	ʽ⮟���r��q2��P�����Ny���/�4w��
׻ڠѻI���m ���_�����rj㼳��v�Z��q���ƺ��1�^}�J��>!��O"�x��%R�T���Tν� ���鞽��l��vbʽz;�mL
�qd�W�!��!���s	�>�����6=��
�c�eu(����b೼�F����W�8�<�r�8��"J�Q�p�і�b ü% �A)���^��}���η�CN����g�U*�1?1���/��/&��y��u�彡|̽�����Ƚ޽' ������&�>n4���:��j8�j�-����[��=�f����윽���W[���>�q�+��� ���F���d"�	6-��=���U���v��>���]нc���'L�#�'���9��F�`J�HF�:�x�(�?��u��;�������Ӱ���|�2�^D�^
P�ޙS�lN�+�A�0A/��j�ŭ���彍�ƽ����c��qې�	5���������gڄ�Z[���\���W���"�������"ͽ��g���U��2�`SF�U}V��_���`��BY�s�J��8�o`%��9�5��k�����O#�>�5��|H�v�W��`�7	`�dW���G���3�j���	����y�н�y���A���*���1��Vu��@j�� ⍽�ᐽ淪��֟�[���8���Yٽ�;�������$��:��N��\\��?c��|a��W��dG�X�4���"�K��K��T�ε��
-�9*@��>R�}�_�ele�/�b�]�W��bF�|�1�t;��B�Q<�"�ҽҟ��l_���棽�8��n����u���ޙ��ٝ�bĤ�L_������o�ӽ�  �  ��.�{�k�󝙽�7�� �����p�o'������bb��A.��LN��+���Z<��hg��йʽ[��@_�N���^�a����Q���罽�=���.l�&�2��T�N���������Q��
#���
������k�A���端���n�!��=W�=񋽗ð�Ci׽k����X�v��ܜ���u�ὒ����^��H���y����⠽�]���ݽ*1���d�/�$�Zz�>+��ڃ۽?��&7����_��&*�t� �}4üd뗼ҡx���[�6�V�j1h��凼4���lӼ:m��.�._�$���������׽������%�p�$�%+#�6c��Ֆ���)׽�Z��f϶�b����н��}5
�%b�/(�!.�`),�>�"����}���Tݽ�/�� ��I����b���F�v]4��)���#��]$��%*��M5��4F�C�]�pH}����Ӭ��%̽�Y�R�������.���9�&�=�3�9���.�+&�nS��t��l�콪'��8��Ɗ�%�(�W�8���C�dG��B��7�9�&�wg�� �N���ǽY%��� ��%��S����9��Y����Έ�.k��������.��	Ӹ�Zν�X����V�w�*�ض<��K��kS�p(T�2)M�b�?���.�e��&������z���*��ڬ,�)�=�W�K��dS�LS���K��>��V,�4%������콙�ѽ�[��/���o��Ye���w��/L��^ȑ�j9䚽��������½��ٽ5_���=�@2�#t2��C�4�P� �V���T�\�K��	=�u�+����J��PL
�
����Y%�Ά6��G��FS�N�X��KV�E�L��:=�b�*�n��W���E�UԽ����=z���-��`\��p���T���Ν�~����	��;��� ½�ս�  �  )�1���d�y��eƮ��[ͽ�S�3���_��������b��ƽ�����ۤ{�c�q�XK��Z���V��"�Ͻ+���Y��^� �zR���e�=�̽��O����g��7��
�-����,���<�]�+�A�E>�K�R�U)�My��7�ϼ$g��[*�]`W��J���;��J�ý���i!��з�`�6���g�⽑�Ž����=�������߁��������½߽����ы�1������̀㽋�ƽL���Jŉ�j]^���1��s��3⼫���kr��+Ή�!х�Ũ������ż},�y���9��d������è��xȽ�g��~������	�{n����ܽɠ���$��N$���b��+��,eؽ�����
��6�����v�o������{ҽ8����/��5����gp�W�NeD��8�z�1��1���7��D���U���m��؅��7���X���qȽ�P���W�Ax��=(�D+��o'����,���+�xO��P۽��׽�Dέ�����	�]��t�'�d1��4��l1��h(�zl�~����������ɽ���x���g���������������������7_���ݣ�z9��x���Ƥҽ�t�n�r�� ��H/���:�SaA�x�A�Vc;���/��!��F��I�X������M'�x���1��-��:��@�(SA�Pg;��O0���!��y��~��:�I�սQ�½��2���k��ߡ��O��?���f6������u8��$ָ���Ƚ��ܽr����Q����hJ'��@5�Ԃ?�!>D��zB��w:�8�-����j���������*���@(��6�O:A��&F���D���<�X�0�;�!�3H����h��GٽȽ�����6���䨽 �����1Ǥ�xo����[���rmɽ��ڽ�  �  C�?�1f��&��t_���ӳ�q�Ž:ѽ�ӽ�̽r�������{:����m�2�Q�h�I���W��x�`��������½|(ҽؽ�Խ�|ǽF���ğ��8��`l���G��'��f
�������ӛ�����F�����=���>ռ�{�![�(�=��ma�y��8������sĽ�`Խ��ܽ�۽��н�m���I��7 ����r�
w\��2[�H1o�`���P��T���X�νͦڽ��ܽ}Xս�"ƽ:!��lO��������f�xD���%�`�����rɼ�L������kӶ��dϼm���j��p0�D!Q��>u��u��'������ũѽ���;��9q��K���:��jyս��H	��W��/������t���5V��V�ֽ���z��������z��9�߽vHʽ�ﵽ����@�����¶q�6�]�0O���F���E�N�L���Z���n����💽U���)����Ƚ��޽�E�����H��b������|���
�O)������OӽZ~ƽ��ýn̽K�ݽ�P��!e�0�Bu����m����#���!C��h��t�ѽ��½1ĵ��̪�c��J��
N���������(_���밽����l?̽^�ܽ	�8��������!�3�(��-�-o,�{�&��������ۺ�����q��%��GR��R����R�%�P�+�d�,�I0)���!�������.&�ڗ��޽�:Ͻj��ӗ�����w���	`������`T������6h���ƽ��Խ�+�<�����T�h���%���,�Rv/��T-�=h&�@��1����?K�������T �/�
��}��`#�3f,�U1��0�d�+��D#�����"����������]�Խ��ǽ��܀�����KR���O���괽���]�Ƚ�_ֽ����  �  (?]��v�5����'���J��$��s�������ɢ�T�������J]�+�;���%�����*���D��Ui��ň����ű�������Z��������ڗ��#�����jlg�azM�M�2���������ټoü 㿼��ϼYT�4��Y*��F��Ta�/p{�2I������wP����������-_���u��䧽^����L���b��(C���1���0��K@���]��ၽ�d�����:��J׵�u��44���0������º���7��_f���L�f�2��w���$���O�������ޒ��9��X�sdw�p̊�|��Ц�����Q���ʽ�Fѽ�{ҽ�0ͽ4���3������b������z���1��7}��|ƴ�PZɽ��ٽfw�����C޽�OԽ6*ɽ�����۱�$������G���� ���Qo�)�c�&�a�:i��*z��'��vk������9s����ýFѽ�V޽	�꽰g���q����:��̟��'�o�ܽ�ʽ�i��Ӱ�������ϵ��DĽ3�׽�i�t� �����������
�<����V���6����ֽbʽ�C��/����Ϋ�굧�C��Q�������ý/�ѽr2��C���W'�7L
��#��;����Z�����Vk��;
�#r �����ݽtս;�Խ�eܽX8뽗;�����DL�����`����N<�:K�ӓ
�8��L����8��⽄lսKXȽ�輽ʄ���`����������;��ˇ̽,-ڽ-�v���rC�P��j��Wp��E��I�������<a�g�	�����M����&�ڽ�Wݽ�������o�Q�����������Q��r�wE�ۅ����y�x:����轧�۽zϽ
�Ľ0���=��)���A�Ľ�Ͻu�ܽ�w꽙\���  �  :-����������ȓ�{��۾���F���ψ��}�'zc�<&E�£&�����B��,D�Y# ��Q�d�0���P���o��儽ѡ���3k��6晽 ᙽ�:��`E���1�������i��6K��-�F�Z�Q���P��"�9@�+`��>~�����c����C�� ;���N���杽dƛ�80��:^������k�(EL�,7.��g�����-��(���*�OVH���g�@���܍�����ᚽJ=���ߝ����ץ�����/���>����h�)K�0���Nq�y���+��&H��j�s8��Ed���p���ɭ�;������|��NZ��wB���t��7W������.��]�����i��)X�oR�Y��l��τ��啽����<���&½�eʽ`dϽB�ѽv�ҽ�-ҽ�xϽ>�ɽ������n���Ά��������"��݊��N���%��&T��	4½[�н�ܽЬ�\+�j��
�D�!�U���׽�P˽q��aݮ����0��0��ڠ�x_��~���eͽ�޽U�����J��?G��`�i��:I��� �;z��8"���/ ؽKwʽ׫��E���l칽@p��Ei̽Z�۽+��^�����E	�9+�Ш�a(����{���M
�G�_� ��򽷽�Ɠӽ��ǽ�����Y���Wƽ��ѽ'��7R����R�E}	����J����yX�n�O�	��i�M��j����ལgҽ�jǽ����N�½.ʽ�gֽ\�����S���\����E�'���8���y(����� ������սF˽R�ƽ��Ƚѽ�޽%��M���e��RK�=��/�<�y{����is�*~����|� 
�����*ٽ��Ͻۤ̽��Ͻ�ٽ���԰��1���	��  �  "���ܪ�,���5p��"Г��8����x�`�7`F�.�+�i(���Aɼ{%��d����ȶ���ռ�Q�и���7��7S�|�m�8������M���䦽u����}���ۯ�7����X��u��ZBb�&B��i.�`	+�1�8�ëT�2z����ɥ��{,��2��⬴�Xɮ�Z�����,��m�N�j��P��4�x��4�2�߼OP˼ʼ87ܼ�������+1�NL�3�f�R��O?��u4��y����t�����ʝ���۰������r��$���H�a�o�G�g�;��A�\�W���{�|g��쨽����7&ǽr̽t>˽dŽ���=�2������'��6���l�j�b(S�9�?�j3�V/���5��AE�>�\���x�q���R�������ȶ�+�ý��н*oܽ��彳��~�뽧��Hؽ�#ǽZ���*������ᕽA������y����н��R��������% �}���\�����꽮z߽1�ӽ/Ƚ�����w�����Mꗽ�+��9������)���z��������,���c½�Vѽa�߽�6��f����xM	�-��>���"���4��
��L���ֽHzνa4ν�=ֽPg�����������t�����e� u����!�����"d���~��2׽Ѭɽ�����P���"��iˮ��T�����w�ǽ+ս:��(4�b�����9�
������>�����n ��[����c�����Sݽֽ4׽���Ƒ����j���7��$�2��\[�(P����ǧ��!��?w�_?彨�׽
˽��7t��1���ض��6���hǽ�Խ��A�� S��!�*f���6�����x��C�#������)W��-�彩��T�佭��5,��6�������  �   �ѽ�SϽ�Ľnj��'t��Nڇ�g�f���A�Z� �`��<8Լ@驼�����Zm���c���x��խ��Q�͗�k�.�-�Q�E�x�Nӑ��	�� ��@νP&ؽ��ؽx�Ͻ[����I��x⍽��r��Y�.UU�of������������Q�ʽأؽ��ܽ�׽�.ɽ��tO��[���gcm��FI�B)���<��⿼*����꒼�⟼p]���#�O	�|�$�R�D�Sh�vˇ��6�������ƽҒս��ܽڽ\�ͽ08�������Ӌ�}u���e�x�k���������P���ν(��|�pr��j&ܽ˲Ƚn����D�������Ux��v[�Y�B�*'.�t���������7��@&�o�9��QR�o�0���F����8��\�½Jٽeｱ:����u�	�@�"�����(�ҽj���3R���ʪ��*������0ٽ=�������k�qJ�����c�D<��߽�˽8���,���a�������2��\�~��x�E�x��Y��t���젒�?������k_��x�ѽ1<�T��y�	��s��X�{�"�v�#�j��my�������[��X�Q���W�� �;c��3�� $��7+��g-���*��#������u:�)*��o�ὼ�ѽýu����v��������Ġ��B��,�������o#Ͻ�߽���Z��O��A"�k�)�\1-��+���%��s��B��k�Ӗ��YK��콮���ed�ֶ�3��%o(���-�>.���)���!��������?�񽲘ཛTѽ��ý𖸽��������?��K�������vԵ�3����ͽ��ܽ���D ��
����\� �x*��`0��g2��t/�O�'�B������p�Ul��I������J����]��o=(��0��  �  9���*e���1�}u˽�V������6�d�Lz3�6�
��Ӽ	���Jo���8�/d��8��g#��xL������߲��=�c���E�Q�y�Z���N����ؽ��� ����03������ǽ ԩ�Lܐ�W���;�}�]-��Pʞ�(����ٽo)�r}����s����*�˽���oɎ��f�.�7��9�\1�(u��O����l�CS��Q�h����ǭ���ܼ����&2���_�A⊽��g�ǽ�e�W;������-��y��r�޽����5ݥ�������o���k<�����W�Խ���fU��&��Y��+�u���u�۽�Z�������8���)d�b/B�t�'��K�>'�� ��q����U���!��8��U�v�x������}��P�Ƚ�=����Zn���2��3U���������kֽ&�Ľ°��Vƽ&�ٽG�����
�;[�&�#�(� �%�tw���������ɽ3ܱ�����e��Ha��Ris��Oh��Mc��rd���k��y�i������4���,��O̽����������!�`�.�)�6�K�8�q�4�=�*��7��.��.������/��p�Z���I+�gO8��h@��"B��Q=�n�2��%����?A�M��
1ٽp�Ž�ܵ�u���YF���������>��,P������ާ�ۻ����½�ս��U��>��"�8!1�c<��A�^A�%�9���-����d���q�_���� ������#���1��=��C��sB�4�;���/��\!�3���6�Ns콷�ֽ�Ľr�������ڣ�w�����'��&L��Cb��Ys������Ndѽ��� ����� 1���,�7.:�#�C�.[G��D���;� S.�8c�X��2d�1�� ��	"������-���;�Q�E��  �  �g����P�����_���r��z.k���/�g{��"g��,�|�1�/��0��ǒû�Ʒ�G8ֻ5��ؕL�������ϼ~t�+D�����y�Ъ̽h��E����O)�����R���㽭n��-���c��������������C�ս�����
����k���F:�o��Z���.A��>i�f1�%���ż�ᒼ��_���2��g�b��ԁ.�kX��5���E�������*��ja��������� ݽ�% �Ǽ�6 �����"����Hܽdѻ��$��&H��Ś�B����˽�#�
���|��pG�5F�>5	�v�FlɽfΥ��ӆ�R7[��J4��������z���d�t��?��X��'�2F���m�`���6/���ѽ���΍�o �}d,��k1���.���$�q������5뽶Rֽ�=ϽÎ׽E���7��o��*�t�5��|:�]27�v�,�!����
�+��*#ͽ����i�����M�t���c�6�Y���U��W��]�31j�nI|������+��톰�L˽o���Q� ��M�.���>�f�H��K��F�F;�2k+����d�SB�cW�.�
������(�;�:�ĴI�-�R��wT�8N��SA� 0�[����	�L?��ս�d��@��x^��yw��LŒ�3⏽7�����.[��(���a૽4}��xNҽ����x�P��c-��?��L��S�Z�S��yK��q=�U,�~������(��	��v�i����0��A���N��U��pT�O�K��7=�=+���������+ҽ�۽���������9��~ݗ�+;��>���욽Bv���P���#���˽<�㽰� ��!��K%��k8�(I���T���Y���V�h�L��?=���+��B��L�+3�����X��*� �<��L�B�W��  �  A�x��^���T��-M˽�����s���0��c��#^���[�.d�V���t�����s�|Ֆ�n�ݻ#^*��Y����¼�T�EeF��h���*��ͨڽ�3�{k�EE��� ���m������Gѽ7���J-���������	ý�N罶�����Z� �
"�g��g����ǽy�����n�l0������ᵼ�⁼�=����u������oS�pM6��Cx����,��5)�
�e�IƗ�pm�����C
��X���!��>!�����|	�K)�7�ʽ�j��GK��������ڽ�[�����1$��J,�׭+���"�"�������%ӽ;��)N��	�X��.��������߼iԼ�Ӽ޼�R���}��e?�43i�Zߏ�.����wٽ�x��9+�Cp8�~>�*(;�,D0�����D�x���!��=ڽ�-�4����p��K#��n5��:B�C)G�NPC��u7�9�%�}��ٳ��|ѽ�k��ū�������Ul�$[��}Q�b�M��O�</V��b�f�s�l����������e~̽G{�@����"��/8�6�I�3U�E<X�i�R��-F���4�O#����Q���	���VA�,�1�{3E�ˇU��~_�Wa�� Z�U�K�8��z"�Y�����XyսCƼ�JL������=�����������ȋ�����%��z�����������ѽ��z�
���,5�kI�2^X���`��/`�CiW��H�T5�h#������������We'�F:���L�q[��Eb�U�`��W�ŹF��^2����X����н����6����T��g���⓽C[��}S��Xז��4��@�������pɽj��+f�]��{~+���@�A�S�� a�X�f��Rc��&X��VG�g4��:#�;������l,"��93�6uF���W�
=d��  �  N���d�����}�Ht^��:�������	��GU��FI�)��8�����ͼ�4���8��J	���ټ�H�!:(� �[�y���ҁ���C��p ��/E�b7i�����|���Y������nH|���\��I<��� �������,�V�/���N�R�o��셾r���Fˏ�w��dxy���W�-�2�����d޽&y��vN��$UI�wj�;J�~���Ҽz�Ѽ�\༴# ����{B��G{��\���ֽV
�'�-���R��(u��臾B����������Gs���R�r�3���(�Ա�M#���>��`���������ޔ���������?{�EX���3��?��罝���*���w���U���@�q6��4�k:��>H��}_������f��澺�����:�o0��8U��Fz��{��L�����L9��[x��%肾�Oe��H���3��z,���3�.H�6
f������������΢��D���m���΄�Bje�ZA�= �)��6޽u@�����M������ጽS;��!�������`���˺�(�ս����Q?���2�B�U�{�����Pݞ�����l'��c$��&���逋��Vw���\�-�L�stJ��JV��=n��;���,����a������a��Ƞ�������;r��CN�f{.�^��# ��a�R5ͽ]���0��Yױ����]1���;����ʽ��޽�G��� �y*���I��"m��'���h��ȧ���������I٦�Q_��2���r��:Z�=�M�hhO�_��y�%��6&������^������<������ ��fg��kD�f�&����[��N߽��̽���$5�����������i��lȽt(ؽJ/ｙ��v1�	�8�y�Y�S-~������١��n���<���\��.x�������F��'�n��Z�c/R�N�X�Z�l�U'���/ä�Ty���  �  ����5���Tw��Y��6������Y��J��!cL��x�������ռ�R���C���0ƼY��cp��	,���^�����[������(���@�Ԁc��-���Q��}��H��ǭu��GW���7�X8������	� ���q+�$�I��i��c���������ۅ�y7s��R�2/�+���ZܽfE���X����L��y#�Ez��.�v�ڼC�ټ���S�]��F�>�}��T����Խ�G�LV*���M��
o��Y��N@���ꊾ%t���m���M�m�/�Ƌ�}����$����:�A=[��{{��k������=��~F���ju�(�S�9�0��{�h>�Jϸ�9p���e{�$�Y�#�D��!:��8�~>��WL���c����������!/�L��t�-��RQ���t��8��m������q�������e`�D��x0��k)�xh0�b<D�,Ea�j	�����ǚ�ɞ��S���!��q���fa�Dr>�	��m6���޽�ѿ��ꩽ�c��w���~䎽47��s�����`i�������K׽������=Q1���R�o�v��Ռ��o��eϤ��G���q���m��篈�p�r�H#Y���I�|WG���R��j�+\���|��4.��ِ��|ګ��ť�-���W3��S�n�L�v-��C�p� ��佪<Ͻ ��/?���۳�ه��;?��XS����̽�u�3l��g���)���G�ͺi�����X���7���"��4ɪ��E���:��ys��aVn���V�ܖJ�@L��i[�O4u��\��晾���q��;䪾����Q���*�����c�U�B���%�R���������l�νýU@������,���{���ʽ�%ڽr��������b7�zW��Lz�uꎾ����	����_������������:҃�(�j�
�V��O�.U�6�h�&�������\��\����  �  ��}��ew�Qe��8J��0+���(a߽�|���-���mW���+��}�`�lټw�Ӽl�߼,R�����{�8���h�!c��^����=e�5���S�,um���}����H�w��c��zG�\�*�c�������Y�
����).;��:X��p�H���7���w��b�y0E� �%���m�׽�5v����X���0����1����T�� %����e2,�KSR�91���{���$ѽ��R!�>�@�F<^���t�Ȕ���4����r�``[���>�<�#�>��-Z�X���{��
.���K��Ji��5���G���Hf}��he��G��e(�@����޺��a�����[Yg��*R���F�{_D���J��GY�q�򂉽㚠��ﾽ�����
��t'���F�Ȏf��>���.��#R��ی�P���o�8�R��8��'�� ��%'��F9���S�^�q������O�����t������su���V���7�]}�}����XŽ3z��"�� D�����XO���Ι��������½�Nܽ�O����P@-��J�C�j�= ��U���L��v��J��$�����@�e��N�}@��z>��I��8^�T.z��ǋ��<���ߟ����5ś��吾:q���0e�wF��6+���j��@꽹�ս}�ǽ�����k���ꪽ��ƽ�\ӽ,�潠h ����Ԧ'��TB�)�`��5���X��s�����*9��La���~�xCb�G�L���A��BC��Q�M�h�����������:T��TR����������DP{���[��;>�9�$�]������D� �ս��ɽ�½XϿ��D��qǽ�Fѽ���.���$�	����u4�B�P�S�o�v���룕�P���=������T���_��\�y�W�_�UFM��[F��.L��]�X�w�a��P̗��8���  �  "�^���Y��\K�O�5���������ٽ�.������ػn�?E���%�.�����6A���/�V;�e�/�AKR��D�f˛�Dj�����>��or%��5>�Y�R���_�Mb�ȴY���G�,00�������]콫��N���s�ǽ%�ת>���S�w�`���c��C[�m�I���2��c��� ��8ս*ܯ�.?���Dq��J���-�f�c��B���Eg*�K�E�:k��`�����Ͻ�����f8/�B�F���X�J|b�UXa��U��xA��5)�e������ct���j7�t�s75��N���b��lm�>(m��Hb�20O�W7��>����B�������K��⽐�*����tj��d]��Y�gr`�+�p�5����>��[��T�ǽ��������\A9���R�
Ci��#y��z���z��8l��dV���=�x(�p������B���(���?���Y�9Hq�����x���R��Dmv��$a�?bH��q/�����*�n�t�нaD��y���h��g��� ���ޤ�Vz������{Ͻ�D罱F����5)��dA��A[�}Ot������<���Ό�����/r��j��iR�w�>��2��)1�P:��L�<�d���}�����Y��«�������܄�\~r���X��@���)�����MU�����V1Խ�?ʽ��ĽɜĽ!ɽ�Xҽn8཮���}��y���&���<��'U��n�*1��\Q������}��Պ���a��,h��QP���=��r4���5�=�A��U�2kn�U���̌�c����(���d��@�����j���Q���9�c�$�:]�l6����e}⽟�ս_�ͽz�ʽ�I̽��ҽ�ݽ��p/��H��{�)2�"I�Tb�)�{�����������#���~��>e���N��?��39�7>��:M��mc�A�|�<ʉ�K푾�  �  �x;��>9�H�/�2� ����������ڽAD��^���勽�@o��lM���3�>$$��  �.�'�� ;�
�W��r|�����$$����ǽ|�jW��Z���'���5�Y$>���>�T27�Z(����� �cP�Q�˽��ǽ��ս��"���� ��s2��=�"�@��<�LU0��P ����*���ڽ�v���������#t��CT��!=��~0�C�/�(�:��P�#7o�B���Ù��&|����ս�����9����-��L:�"4@��>�S�3�Lp#����ό��(�ܽd�ν�ҽ�轇��L���/���@��5J�f~K�=�D�=�7��t'�/���;�YB�(�ѽ	;��`楽�甽�函�g��Fz�g���
���x����D����ٽK�����	������,�k�>��,N�L�X��u\���W�R~K���9�a�%��,�	�\��^�����!Z(�~�=��Q��]_�z�e�Ad�
�Z�e>L��;���)��D�t�
�����Z��<ҽ�z½����ǒ��%��m���������н1N�r���U
�����`(�@�9��L�s�]�h*l���t�7Av�2To��Ja��N�9�;���+�CK"��,!���(���7�ƁK��:`�=�q��g}��]���{�yp���_��N��<��M,�m��,����7���/p�F�۽ Yս��Խ�uڽ�e彠���D���ަ�h�)�d�9�)K��]�T�m���y����K�}�\^s�Y�b���N�g;��',��$���%�J:/� �?���S�ɘg�yTw��	��0G��2y���k��[�?I�P@8�[�(�#:�x!�{�:��������޽��ڽ��ܽ���8|�G�T���B��w$��U3���C�T�U�ϓg�fw�OԀ�݉��C��t�s��`a�7%M���:��+.�~h)���-�@�9��K��W`�=Bs��y���  �  ���x ��?��&��Q�$�����mսx���ޫ�!���͂���e��zQ� �K��V�XTn�����������1:ɽ��ݽ&�񽜞��=���c��h��:���b������ӽ�z��q������)o����ǽ/�?9�9y�E��C6 ��v��S��d��-	��=����뽝ؽ�%ý7w��[)���$���8m�#�\���[��Sj��킽i��ri��������Խ�������[k��������n�����
����kc�J��q\ν�X�� ��}���v½�;޽`  ����P	��U(���+��C*�(�$�rv��l�*.
�p� �N��ڽ��Ž����ߡ�L�������������+���}ɽz��v������P��h�8T%�;�.��|6��;��;�>�5�M+�����[�Y�����v��v���Ai��F!��&1�r=�<�D�&�E��}B���;���2��)��P ����}�������|޽�Ͻ�ǽ��Ž/U̽��ٽ��٩�YS�`��w�#���-���7�v�A��K��6R��U�.LT��nM�f�A��;3��e$�4����e�cw�XQ"�+�1��gB���P�N0[���_��=_�nZ��R��H�T?��95�	!+� ������
�(8����e��뽣9� �P	����{���K)�!V3�>=�m�F��P��UX��]��h_�e�[�$R�|jD���4��T%�ܲ�m����E&��(�,�8�>�H�g�U�^^�=�`��^�'eX���O���F�y=�c3�()����	>�H�	�,=�3��<��dS�>=�����+����Hy&���0��;���D�J�N�X�W�Kq_�a�c��c�~^�	+S���D���4�>Z&��B����c�%��3���C��+S���^��  �  �@���L�i��E�=e�Lq����.���S��{�ؽs���a��Г��h$���c������b㗽�t��}�ǽ���kP���4����^	�VT
�]E
�V	�D�� �pL�"Oڽdh����b2���.�����C���g�������0ѽ�=�����z���	�i���{�7/�`�
��8�[#�lI��iٽC������`K��F���-���C��;ؼ��ֽ�/�Ţ���$���	�l����/B�q	�_��aj�����-սü��w���%��=̎�fꑽ�E��gЎϽ�&뽀����������������AY������4�o�����ؽj)ý5;��	z����������׽9G�|��8�B�+I!���$�XQ&�X�&��&���#�ӕ��g����l��j��?ٽ��˽p�ǽ��ͽ��ݽd���*��z���P ���(��].�[l1���2�<3��:2���/���*��R#�a��E�}��bｩF��ཿ�轲`���5	�ͯ���#���.�Q�6���;�ݠ>�|�?��/@�}[?���<���7��0���%� E�=��d���� ��x �B��m�v����'��4��>�&1E��rI���K�!L�_�K��J�(vF�?:@��7���+������6	����BX���b.���ɰ)��Y5�B�>�#E���H�֬J�n-K�)�J��H�fE�6�>��&5�_w)���/��_����D���K
���xP ��-��8�szA�m�G��K�ҟL��
M��vL��xJ��NF��Y?�9�5���)�S!�.��R�	�p)����@����[%���1���<��qE��K��4N��O�	�O��"O�b�L��HH���@���6���*�/��B����3	�6���������X*���6�l�A��  �  �rԽ@h�*����F�������_��)��{����`!ӽ�Ƿ����۠������h��p�۽8;��Q�������f�� >���9��/����p�?�׽�Uý��J���W���Nl�0>Z��+W���c��}�c���#�����euѽ����o���h����Rm�l��:� ����I������qѽ�s���F���q������ͽ�콏$������AB �;������F����2���V�4�ӽ����	�������Є���q��[g�Ym��&��0>���ç��n���G׽� ���IA�#o�z$ �p(���-���.�"P*��� �����`�Xo�v,ֽ��ͽyuӽ��K���O"�<]/�+d7� �9��7���0�A(� �����/��A��<�۽jȽ�۸�r����P���������Vн�/�j��)
�	�6]�Ej)�sG3��z<�V�C�r�G���F���@��F5��&��P��8
����� �V��C�����0��@�v�K���Q�nR��`N��7G���>��z5�d,�2(#�
��?��r��=������_(��/�(�콊#���*���_b��I(�H�2�zp<��F���O�5�W���]�_`�7�\��9T�P�F�	7�8['�W�����=<����D�%���4�Y�D�ueR���[��8_�3�]���W�ɖO�uCF��<��3�)�ō���LI	�) ����C�1S��������3�G ��!�r�,�|�6�b@��J�isS�}t[�#�`�B>a�
x\��UR�!D��24��w%����������f� ��.�K">�=�M��*Z��a��c�1�`�^�Y��KQ�n�G�`q>���4���*�L+ �v��d�������������������>��z�Bv ��]+��  �  M���+۽%����_�4�!���0�_U:��h<�/*6�g(����h���߽��Ƚ½0ͽ��(���6��y-��:��>��;�fy0�9!�C������Wq۽Pp��ɺ����It���S��[;�R`-�N+�x�4�h�I���g�C���9o��S6���ѽr�e{	��p��L,�@�9�ڮ@�L�?���6�o�&���sZ��zI޽1
̽��ʽ9O۽�������"�$��5���>���@��(:��k-�k��@�
�ZC�m�ӽ')��Ο�"���Pq��fU�yC�x�;�^RA�"�R���n��牽֟����#(ԽH���8
��_�^�.���>�=�J���O��L�z�A��l0����e
�YB���ｐ���*������-���A� #Q��Y��X��{P���B�!�1�� �ބ�O� �<#置,н�J���֫�K���W ��)~��O����,���I��!bǽ]�ݽ�����E	����$�)�`<�ܵM��\��Tf�c�h�ћb��0U�O�B��/��=/�������@�$��F8��|M�Mj`���m�}�r���o�{e��qV��@E��4��S$��_�Z*
����P�콗.޽��ӽ�yν�ν�6ս"�����>���"�51(���7�X'I�G
[���k�^�x�0��x�~���u�P�e���Q���=�ȵ-�ً$�% $��),���;��#O�k1c���s���}��t�N6y���l��\�@J���8�:)�v<�������'���o��LL۽ )ֽ�׽j�ݽe�齭*��D	��}��h���-��@>���O�M�a��q�?o}�7��q�~�.s���a�a|M�v�:�8�,�Ћ&��()�c#4��vE���Y�1Im��|�����O���!z�l���Z��6I��y8��i)�l��9�����*����콵��S�ཇ��c�콵8�����|��u��  �  i��ݍڽ̷�#/�2S7�{�L�0/[���_���X���H�d�1�p���&�3��C���5�!�~�*8�;\N�� ]���a�3[��(K���4�&��W��zcؽ���M����ar�RJ�B},�����h��
�W���$�&�>�G�b�����Х�<uɽ����:�.�+�D��rW�!�b�o<c���X���E��y-�>�^�E����[���k�lw*�g�B���V��8b���b�)�X���E��.����xb��!vͽ{���U���X�k�<�H�0��5!� &�?=!�FS0���H���j�9��s@��&ǽk��K���'��A�0	Y��cj�H�r���o�7�b�W�M�s�5����:s��^��3�]�aP/�`�H��]a���s�.H|���y��m�2�X��L@�s.'�S��L���zֽ���>���ɗ��9��h���n��j��c/��Y��������gɽ��������A0���I�� c���x�B���!䅾���ZOu��^��lF��Y1�Գ#��2 �V�'��8�=pP�=j�V���@���Ê�qŇ�~���j�0GQ���8��"�����D���׽6sʽ ����ɽ�3|��"�ýY�ͽ�Nܽ�J����a�EW$���9���Q��ck������c��e吾�#�����G��*-l�Z�S���?���4���3��>���P�"i�Kʀ�͊������Ր��ԋ�f����Om���S��x;���%���i%����wc���ҽ�ʽ)�Žܟƽ<6̽�uֽL^� 0���.	����!�+��<B��3[���t�=텾Zw���k���5����_Yf��&O�\>�Uc6���9�G�HQ\��Fu�����U��8a��SOg��O��ݘi��SP���8���$�g��'�ڜ��R��Eڽ�ӽ��нD'ӽ�jڽ^M�s���LD�y���  �  iѯ�/��dE��,�gL���f�L�x���~��xw��Zd�q�I�8�,��i�H�����������D�3�AQ��j��{��T���x��d��0H�{�(�{�	�5�ܽV3��d��,qZ�t�0�mn�[m ���켪���������%�6�I�<|��F����ɽ<���4��8�<�0�Z���r�?����:��t�v�ie`�iD��'������������$��@�0-]�Xkt��������t�G/]��~?�������ν�ң�7o����R��o/�� ���
����I��%���}0�܇Q��~�'ל�x�½#�����Y4�mT��vq�]���<Ј�
�����Q[g��J��Y0����G��^��9)�s�B��h`�ӹ|��툾���Eڋ�����3	n�H�O��\0�g�� ����νH�����������K����x��gw���~�Hi��V���Oڥ�@���?�ݽP������8�8�X�I�w�]���p��x�������E���1�v��?Z���A���1�D-���5��I��	e��|������P����;��Z7���l��~d}�Ow^��@�m�$�H(�����޽��ʽ�ɽ�������{}��Ot�������_Ͻy�⽎x���#t$��}>�Dd\�|��	��l����.����֚�,���Eb���?f��:O��B�\TA�M�[c��)�x卾4���5��L'������-$��2�~�`_���@�M�&�������F���ӽ�ƽ\���*��������ʽ�ؽ@	�(d���=e-���H���g���������ɜ�C桾�l��!���<:����{�5�`��L�Q�C��HG���V�y�o�Wf���8��y��%��h砾$���XƋ�o�x���Y��<�
�#�=���y ����XWٽCIν��ǽ��Ž�
Ƚ-�ν��ٽ{�� �_���  �  ������}T�D�7�w
[�a;y�Wˆ��4���4��Yw�z�Y��:��P������g��m$���A���a�m~�*���j���9��6�u��[V�73� 2��⽳E������I�N��y#��� ����Ӽ�,Ѽ w޼���y��,9=�Ŏr�Oz��s�̽Cr�z %���H���j������h��-�����r�*cS��"4�e��6��6��ȟ���0���O��o��P���t���`������m�@^L���(�\���Xҽb���� |�r�F��/"���
�0���}���������M#�@gD��r�����jb½�������a>��3b��r�� �������c/���͉�Ңx�;JY�S<���&�HQ�{�!�0�3���O��Qp�`���K������>K��o���s}��[���7��f����i0̽�v������X���tu��l��+k�]r��瀽H���`������Ǧڽ���@�]�?���c�rp�����ZМ��O���n�����}����g��nL�ɵ:���5�v<?���T���r��剾6t��'��7����Y��D��������h�S2F���'��+�����8ؽĽ����d��gP���7������ۺ���Ƚ�Hܽߣ���)���%��C���d��9��T'��[����������f
��b���2
��ѿr�WwY��	K��4J�fW�2No����Җ�R���Dת�XЪ�a���mu���Å� �g���E�N(�{=��j��4���̽��8���Ӵ�u���#���Eý�ѽ<�dh�$N���/�x�N�-xq�h���?˚�٦�����A������ؔ���+l�BV��^L��kP���a�[�|��a��˔���ܨ�ϭ��\��S��#~��Y5��a��h@�x�$�Ә�j����h��ҽY�ǽ@���z��������ǽ��ҽ��X���oE��  �  �̱�B�꽩�r�;���`���z�������~��_���>�)"��N�%�	�#��Os(���F���g�����_������䉾	@|�5�[���6�O��)u�t���X܄�o�K��x�Ƽ��޼�˼ ɼ�Gּ�b���f���9���o�oF��;νL��L(��}M���p�����ۏ��9����x�U�X�ڍ8�t����v���(��5�u�T��_u��釾�K���4��������s�Q���+���Խ������y��KC�*�����������Ɲ����3�Dn@�H�o�y��F�½K����˼A��Ag�[����F��/r�����RS��d�~�6a^�A'@��*�he ��+%���7�QT���u����y���(`��9��Ł��G���AY_���:�-������Ե˽����-�� H��Sq�yh��/g��Vn���}�+6���p������ڽ���g� ��B���g�_/���镾�����,�� )��o���_���\l�0CP���=�Z9�p�B� �X���w��⌾�蛾4쥾�Ш�����z��7Z��`l�7�H��(��g�`3��Տֽ�½�ش�(M��7D���-��1쯽
����sƽjڽ1W������&�~�D���g�������N=�����^�������㛾 ����*w�*]�c.N��RM�"�Z�Ԟs�һ������A��㭮���������|���"���*k���G��&)��7��9��lH޽�ʽ/׽�I+��.в��o������-����Ͻ�f�'�� s�%�0�o�P�Bu�� ����py�����N䮾����痾�~��Ip�&�Y�CtO�5�S�*ke�"���p6���蠾����l������f��IP��X����c���A��6%��Y��E���|�3{нE�Ž����Ъ�������Ž��нl�὾��,���  �  ������}T�D�7�w
[�a;y�Wˆ��4���4��Yw�z�Y��:��P������g��m$���A���a�m~�*���j���9��6�u��[V�73� 2��⽳E������I�N��y#��� ����Ӽ�,Ѽ w޼���y��,9=�Ŏr�Pz��s�̽Cr�z %���H���j������i��-�����r�+cS��"4�g��9��:��͟���0�əO�o��P���t��
a�����F�m�u^L��(�����Xҽs���r |�~�F��-"���
�W���Ԫ���q������B#�ZD�v�r��UX½�������$>�J-b��o����������,���ˉ�0�x�kGY�\<���&�Q��!���3��O��Tp�g���hM��o���6N��� ��.z}�-[���7�ul������9̽�~����m]��E{u�l��+k�8Zr��䀽C���Z��	�����ڽ���;�"�?�
�c�&m��ې��B͜��L���k��}��@{���g��lL��:���5�p=?���T���r�_牾{v���)��,���]��wG���ą�d�h��8F�Ɉ'��1����JAؽ�ĽD���Vi���T��(;��X��)ݺ�H�Ƚ�Iܽ�����)���%��C���d��9��V'��]���	�������g
��c���3
��ҿr�WwY��	K��4J�fW�2No����Җ�R���Dת�XЪ�a���mu���Å� �g���E�N(�{=��j��4���̽��8���Ӵ�u���#���Eý�ѽ<�dh�$N���/�x�N�-xq�h���?˚�٦�����A������ؔ���+l�BV��^L��kP���a�[�|��a��˔���ܨ�ϭ��\��S��#~��Y5��a��h@�x�$�Ә�j����h��ҽY�ǽ@���z��������ǽ��ҽ��X���oE��  �  iѯ�/��dE��,�gL���f�L�x���~��xw��Zd�q�I�8�,��i�H�����������D�3�AQ��j��{��T���x��d��0H�{�(�{�	�5�ܽV3��d��,qZ�t�0�mn�[m ���켫���������%�7�I�<|��F����ɽ<���4��8�<�1�Z���r�?����:��v�v�ke`�kD��'����$�������ǒ$���@�G-]�wkt�1���6���;�t��/]�b?�g������ν�ң��n����R�Dl/������
�e��������_h0�FnQ��j~��Ŝ��½���=���M4��`T�jq������ʈ�*z��^��VTg���J�	V0����ԋ�����;)��B��n`���|�=�F����ߋ��ǃ��n���O��h0����E.����ν}���锚��!���Q��5�x�!hw��~�mc��g���TΥ�P���ݽ.��߸���8��|X���w��V���j���{�������d�v��:Z�R�A��1�6D-�x�5�ÙI�e����Ď�d���UA��=��%s���q}�D�^�S@�(�$�3�"���޽{�ʽ�ս�c��x���-����y�������bϽ���#z����|t$�&~>�`d\�|��	��o����0����֚�.���Fb���?f��:O��B�]TA�M�[c��)�x卾4���5��L'������-$��2�~�`_���@�M�&�������F���ӽ�ƽ\���*��������ʽ�ؽ@	�(d���=e-���H���g���������ɜ�C桾�l��!���<:����{�5�`��L�Q�C��HG���V�y�o�Wf���8��y��%��h砾$���XƋ�o�x���Y��<�
�#�=���y ����XWٽCIν��ǽ��Ž�
Ƚ-�ν��ٽ{�� �_���  �  i��ݍڽ̷�#/�2S7�{�L�0/[���_���X���H�d�1�p���&�3��C���5�!�~�*8�;\N�� ]���a�3[��(K���4�&��W��zcؽ���M����ar�RJ�B},�����h��
�W���$�'�>�G�b�����Х�<uɽ����:�/�+�D��rW�"�b�q<c���X���E��y-�C�^�$E����w���k��w*���B��V��8b���b���X�&�E�.�%��oc���vͽ����栌���k�s�H��0��*!�m� *!��:0�Q�H�*�j��#���'��I
ǽ�{:���'�ːA�'�X��Sj��r��o�a�b���M��5�|��Bp�/^��5�a��V/�I��ha���s��V|���y��(m���X�)^@�??'������s�ֽI	���P��'ח��B���l��3o��f��'���}��{u��MRɽ��彃�����00��I��c�&�x�瑃�m܅�2����Cu���^��eF��T1���#��2 ���'�/�8��wP��Fj�p���.G���ˊ�·����R(j�|YQ�O�8���"�:.���~7���׽݄ʽ�����ս�������ý�ͽ�Rܽ�M�)���b��W$�Ȭ9���Q��ck������c��i吾�#�����G��--l�]�S���?���4���3��>���P�"i�Kʀ�͊������Ր��ԋ�f����Om���S��x;���%���i%����wc���ҽ�ʽ)�Žܟƽ<6̽�uֽL^� 0���.	����!�+��<B��3[���t�=텾Zw���k���5����_Yf��&O�\>�Uc6���9�G�HQ\��Fu�����U��8a��SOg��O��ݘi��SP���8���$�g��'�ڜ��R��Eڽ�ӽ��нD'ӽ�jڽ^M�s���LD�y���  �  M���+۽%����_�4�!���0�_U:��h<�/*6�g(����h���߽��Ƚ½0ͽ��(���6��y-��:��>��;�fy0�9!�C������Wq۽Pp��ɺ����It���S��[;�R`-�N+�x�4�h�I���g�C���:o��S6���ѽ	r�f{	��p��L,�B�9�ܮ@�M�?���6�s�&���Z���I޽E
̽��ʽ[O۽)���ݐ�I�$��5��>���@�):�-l-�����
��D�G�ӽt)���͟�����:Jq�`]U�.C�V�;��:A��R�P�n� щ����������Խ҉��$
��J�P�.�$�>�c�J���O�y�L�)rA� a0�����_
�/;��Qｵ�����Ֆ�,�-���A��2Q��,Y�b�X�B�P��B�X�1�)/ �H��� ��B�~Gн�`���竽����>&���~��b�g"��&:���Lǽ�ݽs����3	�>��C�)���;��M���\��@f���h�9�b��"U���B�/�J�s,�݃����f�$��O8���M�y`�ˢm���r���o��e�M�V�$WE��04�1h$��r�];
��%��+��qD޽��ӽ��ν��ν�?ս2��(���?�h�� ��1(�K�7��'I�c
[���k�l�x�<����~���u�V�e��Q���=�ʵ-�ۋ$�& $��),���;��#O�l1c���s���}��t�N6y���l��\�@J���8�:)�v<�������'���o��LL۽ )ֽ�׽j�ݽe�齭*��D	��}��h���-��@>���O�M�a��q�?o}�7��q�~�.s���a�a|M�v�:�8�,�Ћ&��()�c#4��vE���Y�1Im��|�����O���!z�l���Z��6I��y8��i)�l��9�����*����콵��S�ཇ��c�콵8�����|��u��  �  �rԽ@h�*����F�������_��)��{����`!ӽ�Ƿ����۠������h��p�۽8;��Q�������f�� >���9��/����p�?�׽�Uý��J���W���Nl�0>Z��+W���c��}�c���#�����euѽ����o���h����Sm�n��<� ����I�
�����qѽ�s���F���q��!��7�ͽ"�콺$�Ө�i���B ����K���G����~���W罔�ӽ_�������d˄��|q�eGg���l����!)��8����P���%׽p�����*��W� �Y(���-�r�.��=*��~ ����V�Wa꽚$ֽ7�ͽzӽ�潗S����]"�sn/��w7���9�p7�%�0��0(������)$�;S�[1��۽�|Ƚ�踽#���iQ������V���Dн��RL��r
���GG��R)�S/3�Ub<���C��G��F�m�@�h75��&�lG�F2
�x��' ���JJ�|����0�� @�j�K�?�Q�@�R�AyN��PG���>�+�5�{,�v=#�;��-�������n��9�==彂��p+���-����c��J(���2��p<��F���O�M�W�
�]�n`�C�\��9T�W�F�	7�;['�Z�����?<����E�%���4�Y�D�veR��[��8_�3�]���W�ɖO�uCF��<��3�)�ō���LI	�) ����C�1S��������3�G ��!�r�,�|�6�b@��J�isS�}t[�#�`�B>a�
x\��UR�!D��24��w%����������f� ��.�K">�=�M��*Z��a��c�1�`�^�Y��KQ�n�G�`q>���4���*�L+ �v��d�������������������>��z�Bv ��]+��  �  �@���L�i��E�=e�Lq����.���S��{�ؽs���a��Г��h$���c������b㗽�t��}�ǽ���kP���4����^	�VT
�]E
�V	�D�� �pL�"Oڽdh����c2���.�����C���g�������0ѽ�=�����z���	�i���{�8/�b�
��8�]#�rI��iٽM������vK��c���B-���C��~ؼ�ֽ_0�`���2%�/�	��l�Y���B��q	����j��
��N+ս����|r��$������cܑ��3��Rش�,tϽn뽃��������������\���A���<����a���h�lؽ*ý83��Wx��#!�������׽�^�̊�pJ�V�>_!��$��i&���&��7&�p$�����z����i��8��Lٽ��˽�ǽ�ͽA�ݽ����������^> ��(�G.�T1�߱2�:�2��"2�߯/���*�@#��	�9�qs�/V�u@㽂����dn���?	�4��0�#�ݭ.�#�6�a�;��>�]@�{I@��t?���<��7��/0�Y�%�{T�6�#��?� �� �fG��q�{����'�_4��>��1E�SsI�ށK�A!L�{�K��J�:vF�M:@��7���+������9	����DX���c.���ʰ)��Y5�C�>�#E���H�֬J�n-K�)�J��H�fE�6�>��&5�_w)���/��_����D���K
���xP ��-��8�szA�m�G��K�ҟL��
M��vL��xJ��NF��Y?�9�5���)�S!�.��R�	�p)����@����[%���1���<��qE��K��4N��O�	�O��"O�b�L��HH���@���6���*�/��B����3	�6���������X*���6�l�A��  �  ���x ��?��&��Q�$�����mսx���ޫ�!���͂���e��zQ� �K��V�XTn�����������1:ɽ��ݽ&�񽜞��=���c��h��:���b������ӽ�z��q������)o����ǽ/�?9�9y�F��C6 ��v��S��d��-	��=����뽡ؽ�%ý>w��e)���$���8m�N�\�%�[��Sj��킽Ti���i��1����ԽA�������k�X��g��lo�6���
�����b���KWνcQ������eo��ce½�%޽����������2B(�o�+�N-*��s$�_�V��
��� ��*�l�ٽ�nŽn	��Iҡ�� ����L������N�ɽ�������&��De�C��k%���.��6�4;�c0;�u�5��+�]���e�Xf������潰��� `�5:!��1�`=��qD���E�hfB���;���2���)��: �������z��K �Uj޽��Ͻ�ǽ#�Ž�[̽�ڽ8"���c����R�#���-�8�tB��,K�lOR�z�U��aT�Y�M���A��J3��r$��>���l��|�LU"��1��iB�%�P�51[�&�_��=_��Z�&R�0�H�l?��95�!+�̈ ������
�-8����j��
뽥9� �P	����{���K)�!V3�>=�m�F��P��UX��]��h_�e�[�$R�|jD���4��T%�ܲ�m����E&��(�,�8�>�H�g�U�^^�=�`��^�'eX���O���F�y=�c3�()����	>�H�	�,=�3��<��dS�>=�����+����Hy&���0��;���D�J�N�X�W�Kq_�a�c��c�~^�	+S���D���4�>Z&��B����c�%��3���C��+S���^��  �  �x;��>9�H�/�2� ����������ڽAD��^���勽�@o��lM���3�>$$��  �.�'�� ;�
�W��r|�����$$����ǽ|�jW��Z���'���5�Y$>���>�T27�Z(����� �cP�Q�˽��ǽ��ս��#���� ��s2��=�#�@��<�MU0��P ����*�� ڽ�v���������#t��CT�"=��~0�u�/�i�:�9�P��7o�����&����|��(�ս���i���1�-�XM:��4@�,>�"�3��o#�9��0���_�ܽ�ν��ҽ轶��r���/�s@�$J�kK�ձD�D�7��_'����h(��콛ѽ���%Х�}֔��ه�tZ�!Dz�K������������(���ǧٽT����	������,���>��AN�P�X�:�\�s�W���K�(�9�B�%��2�>����������Q(�9=��
Q�'M_���e�d�ŹZ��(L� �:��~)�]1���
�a����i彑&ҽ�j½�ﶽ����~��U��������н�d�;;���e
�;��8u(���9�A1L��]��@l�
u��Tv� fo��Za���N�и;�v�+� S"�3!�|�(�K�7�]�K��<`�z�q��h}��]��m�{��p���_��N��<��M,�{��6����A���7p�L�۽Yս��Խ�uڽ�e彡���D���ަ�i�)�d�9�)K��]�T�m���y����K�}�\^s�Y�b���N�g;��',��$���%�J:/� �?���S�ɘg�yTw��	��0G��2y���k��[�?I�P@8�[�(�#:�x!�{�:��������޽��ڽ��ܽ���8|�G�T���B��w$��U3���C�T�U�ϓg�fw�OԀ�݉��C��t�s��`a�7%M���:��+.�~h)���-�@�9��K��W`�=Bs��y���  �  "�^���Y��\K�O�5���������ٽ�.������ػn�?E���%�.�����6A���/�V;�e�/�AKR��D�f˛�Dj�����>��or%��5>�Y�R���_�Mb�ȴY���G�,00�������]콫��N���s�ǽ%�ת>���S�w�`���c��C[�m�I���2��c��� ��8ս-ܯ�2?���Dq��J���-�~����j� ��g*���E��k�a��n��:�Ͻ����|���8/���F�#�X��|b�zXa�ĒU�>xA��4)�������l�N���0��k��-5�d�N�v�b��]m�Vm�'8b��O��E7��-�Ջ�|��c����5���Ru���aj��Y]���Y��x`��p�����N��3o��\�ǽb;�I��\���R9�	�R�ETi�*4y�B����z�aDl��nV�W>�z(���ܜ��@�3�(���?�_�Y��<q����p��EJ���[v��a��PH��`/����m��T���н3��t�������:����x㤽����Ѵ���Ͻ[��S���zF)��vA�LT[�
bt�����KE��׌������x��^*j��sR�`�>�x�2��.1��S:��L�\�d�<�}����[Y����������܄�~r���X��@���)�����ZU�����]1Խ�?ʽ��Ľ˜Ľ !ɽ�Xҽo8཯���}��y���&���<��'U��n�*1��\Q������}��Պ���a��,h��QP���=��r4���5�=�A��U�2kn�U���̌�c����(���d��@�����j���Q���9�c�$�:]�l6����e}⽟�ս_�ͽz�ʽ�I̽��ҽ�ݽ��p/��H��{�)2�"I�Tb�)�{�����������#���~��>e���N��?��39�7>��:M��mc�A�|�<ʉ�K푾�  �  ��}��ew�Qe��8J��0+���(a߽�|���-���mW���+��}�`�lټw�Ӽl�߼,R�����{�8���h�!c��^����=e�5���S�,um���}����H�w��c��zG�\�*�c�������Y�
����).;��:X��p�H���7���w��b�y0E�!�%���n�׽�8v�� �X���0����B��󼍕�F%�ӿ��2,��SR�p1��|�� %ѽ��CR!���@��<^���t�䔀�5����r��_[���>���#�B��qW�����v��.���K��Bi�1���B��E���\Z}��\e���G��Y(�*�����̺��R��W���Eg�2R�>�F��]D��J��QY��q�'������� ��]����g�'��F�1�f��D���4���W���ߌ�5T���o�y�R���8��'�� �'$'��C9���S���q������J��F����������fu�s�V��7� r�O��@���HŽ	n�����>������O���љ���������ýP^ܽ�b������K-��K�Hk��������:R���{������ ��ŀ��e���N���@��~>��I��:^��/z�ȋ��<�������Oś��吾Gq���0e�!wF��6+���q��I���ս��ǽ�����l���쪽��ƽ�\ӽ,�潡h ����Ԧ'��TB�*�`��5���X��s�����*9��La���~�xCb�G�L���A��BC��Q�M�h�����������:T��TR����������DP{���[��;>�9�$�]������D� �ս��ɽ�½XϿ��D��qǽ�Fѽ���.���$�	����u4�B�P�S�o�v���룕�P���=������T���_��\�y�W�_�UFM��[F��.L��]�X�w�a��P̗��8���  �  ����5���Tw��Y��6������Y��J��!cL��x�������ռ�R���C���0ƼY��cp��	,���^�����[������(���@�Ԁc��-���Q��}��H��ǭu��GW���7�X8������	� ���q+�%�I��i��c���������ۅ�z7s��R�2/�+���ZܽgE���X����L��y#�Lz��.켍�ڼ`�ټ>��T�~��HF�w�}�U�� �Խ�G�nV*���M��
o��Y��\@���ꊾt���m��M���/�������������:��9[��w{�"i��@���:��eC��=du���S�|0�/v��3�Ƹ�Mh���X{�&�Y�0�D��:��8��>�U]L��c�����M��\���'9����|�-��XQ�!u�<��&p���"��;t��>����ih`��D��y0��k)��g0��:D��Ba�������'Ś�5ƞ��P�����'��p`a�l>�:��,1���޽ʿ�x䩽�^��]����⎽N7��)���c��Un������S׽u��p��FW1��R�/�v�Vٌ�5s���Ҥ�K��|t���o����� �r�7&Y��I�WYG�A�R��j��\���|��e.�������ګ��ť�6���^3��^�n�L�v-��C�t� ��佭<Ͻ��1?���۳�ڇ��<?��YS����̽�u�4l��g���)���G�ͺi�����X���7���"��4ɪ��E���:��ys��aVn���V�ܖJ�@L��i[�O4u��\��晾���q��;䪾����Q���*�����c�U�B���%�R���������l�νýU@������,���{���ʽ�%ڽr��������b7�zW��Lz�uꎾ����	����_������������:҃�(�j�
�V��O�.U�6�h�&�������\��\����  �  5�꾦�ƣѾ��������5�u��D@��L�E�ȱ������Wk�>L�;<��	8���?��lT��x��3������M��>=��M�"}���蠾���Oؾ���X\�/ 㾱�ξ���|������~g�ZJb�a�t�����ԧ���þX�۾le꾙�쾒����˾���V鐾�g�0/5��b��jڽ�쬽���?o���T�N�G���F�i�Q��Vj��]������6Iӽ���8/��`�3񌾷���waȾ�߾]U�K��Aݾ�>ƾ����{u����x�^�d�~�h��4S���C���о0�L�����Uf�39ɾ�ƫ��v���?c�&@4�+'����ꩿ����Q��-i�������������`��a����(彿����-��EY����뤾��þv߾����� ���/徱/̾����헾2�e����^����i���2�˾9?����P����u��(�q�̾)[��ۊ��Pl��G@��s� �������ѽ0�ý���0����\½]ν������[��t�/�]�T�����|r������J!ھt�����$��Z��}�뾬SѾUf�����5���`������鄭�v�Ǿ�㾶����U��r�� ��8��Ͼ�����Г�t�t���K�L�,����������L轶��K�_��,󽓶�����(��G���n��$���쬾Җ˾����G��~���w�ڀ��#l���ʾMR�����|���(��<���_���\Ѿ+�쾐� �9j�M�-���~P�4�ž;B��MP��dg�x�A���%�g��+���n����� ��������  �Z���^�� 6�hW�JI��Q����^��k�׾�m�̔����Z(�=<��3ྗ:ľ%Z��������J���LG��ک��W�ݾt|������  �  ��شݾI�˾Ud��rG��)q��=���A彘$������q��R��(B� >�>F�Q�Z��m~�� ��;������^D���J�����D�����8uҾp⾇�従�ܾNɾ�J���Ĕ�t}���b�7z]��@o��_��Ǚ�����h�վ�㾱��;�۾éƾ�\��*��d�Q3��+�.�۽񒯽 ���u���Z���M���L��7X���p�΅���x��B�ԽF����-� ]�����w��!-þ��ؾ��f侉(׾����1n���	��Mss�@"`�:�c�h�}�躔�(�����ʾ��߾���Z�w۾�Dľ���芾�U`� 3�9U����a�½)F��߆��8��z�������������ý���zf��5-�<+W�����f������
|پ�v�f����ﾮQ߾5Ǿ%���񾔾(W��:�|��Ѓ�듾�ԫ�5&Ǿ�Ą�4��l󾔄��Ⱦ( ��_��׽i���?������ڤ��Խ�ƽ;��a���!fŽ��ѽ���*� ������/�`�S��L��� ��[R���Gվ�������� ������徻�̾������%���*(��|(��X�þ�޾����I�e!�����T�澴�˾e	��] ��`Ls�X�K��i-���U7������l���佝N佀��O��?J�v\�O�)���F��Nm��r������ǾkT�w)��~�}+��e��#ᾔwƾ�ᬾ%N���M���������p����̾��<�����E�����_Y޾+���ѱ���؉��?f��%B���&�n*��g�ܡ���G����뽆	������o�m����6��V�?�� ����#��ˇӾ���i ��Y����D`�$۾�5��$+�������5��Fe���,��Ӿ��v�ؾ@�񾵵��  �  �Ѿ̾�p��F㥾H7��j�e��t8�������o�����4����f�0U��P�?7Y�%�n�a����ࣽ�OȽ�5��qo�&8D�=Es�sn��HାX¾$о�3Ӿr˾/s��:���I���l�2VT���O���_��ꀾĶ������w�ľg�Ѿ.�Ӿ�jʾ6��m����	��1�Z�w�/��u���4���mU�����D�n���`�Q�_���k�Ě���Ȗ�伳��۽|A�Lk*��{T�ᖂ�{{��A鴾�ȾKmҾ��Ѿy"ƾ2��mK��Oc����c�ҀR��U��Zm�������,]����ξ��ؾ�D׾�˾���͝�b#��xY�-�0�H��RT��1̽񛲽婡�$���e���0������~̴���ͽ"���\�,��,R�A�@���W����8ʾ��ھ��ᾲ�ݾ��ξ�?���;��������y�	o�� y�9/���ؠ�{���#gоn��:���o�� ҾT�����������<d��>��9!���
�Ɯ��o߽��нҁɽ��Ƚ��νLz۽Y+�q��g�'k1��Q���y�ː��x��&	Ⱦ,�ݾo����a�?־�����!��c���|􈾺���q������*���lо���|��l��h��oIؾ '�����AW���so��L��o0����YQ�����;���1�����B ��j
�U����,�ӧG�3�i�9��&��������վ>J�������X�|SҾ�I��9.��
y��ok��ߠ��_唾�9����ٴ׾�H꾧��s��pl���о����i蝾+����c�	�C�8�*����W�
�Ia����zD�V��f���^���x�'�"�r 9�ifV���{�~/�� v���eǾ^�޾^Sﾺ5��D����.";�崾-��~��Sh��p��nf��]����˾>�ᾡ��  �  ��������������=����W��\3��g��T��Uν.i��-U��/Z��`�v���q�/Z{������ל���ٽx����U=��Ac��K����������n���򼸾��������f ���u���S�9#?�2G;��I���e�FH��К��d���V���c��fN��ڼ��/�����w���O��-�������4%˽�ѭ�ϗ��Ո�����x��EL���D���B���ƽ����C���(���J���q�񞍾���7X��/f���t��ֈ���������mJj�'�L�>�A�JU�,Qw�4z���!��w|���0��ݘ��t!��G���4w�];Q��0�q���^ ��Z߽�ƽ���0N���ॽ�穽-D����ǽw"�p� ��z���.�
�M�Ger�E����V��괾.¾�}ǾH�þ +���㤾������|�@�c�.�Z��uc��{|�d����������~�ƾb\̾�wȾ�N���q��,��}Ɂ�a-_��p@���'�X���y*�Ϛ⽉Dڽ>PٽJ�߽���#���.� ���6�}�Q���r�����|P���Ƶ��Ǿ�Ҿ�Ծ^�;�~��Ea�� ���4��ޑ|��y�b�.���p5���庾�̾>�׾��پ-�ҾH�þA����ߛ�������l���O�r�7���$�[�L�
��c�1���4I�����?�	�&��\"�G�4��K�.h��?��a☾�����<��φо��ؾ��׾��;ż�/q��y۔��υ�(6|�%I~������,���]��ea���Ѿ�Fپw:ؾjξ����G����Y���B���c�}H���2��!�F?�>�
�im�p�� ����F��2���+�]�?��X��Nw�Gɍ�����϶��[ɾ|�־z�۾Z�׾�A˾3ɸ��H���ܑ�L��T5��k:��f��̀��S��',ʾk�׾�  �  ������������4���j���M�J�3������t���ν�|��A �����Ot���N��z���ώ���b׽b��$��~�#�R�;���V��Ws����-v��[����C����Q߈��1r��Q��6�v�%�c�"���-�UE��%d� ����ʐ�J���Hr��� ��/L������be�ړI�l0�]F�3���I�JyͽE���h���֙��9��䞡��7����ɽ���/-�n;���,�:�E��a�]�}��P������ԯ�����M������u�g��H�'Y1�V�%�,K(���8�fkT��v�N����+���Ġ�2`���a���o���̂��,i�pN�7�6���!� ���������fн."ý-o���½@н�g�*z �����1#�7�7�k9O��xi���xu��A��+��R8��h��f/��^���g�z���]��I��uB�N�I���]�R�{�Fӎ�C�������7��*-���'�����֊��~y�	�_�e�H���4��#�[�������� `󽙳�y3��ܣ��[����
0��/C�3�X�q�V ��L���wߢ�B���_�����wD��Ō���E��܇��p�r�8c�=�`���l��3�������������4��$���yc��+����=���Œ�Ǆ�B5p��Y��;F�i�4���%�����������^����*�#��z2�)fC�F�V��ul�멂��z���랾}j���ɶ��ܻ��9��Sϱ�����Ǔ�v��~�o���c�|?e�/�t�3����ʗ��㧾�����Ȼ�v���V���q��補��N���Հ�)�i��T���A���1�R�#����KY�&4�	���r��3�|1,�0�;���M���a�j�x�/\��3�������������������Ū���J��hh������2����o��h�O�n�-��ȡ���0��l�������  �   M|�6Z}�~�v�'�j�S\��fM�d�>���/�� �����W��a�߽��ƽ������O����̽��罊������b%��5�1D�NLS��zb���p��|��ƀ�p�~���r���^��EF��.-�bR�8��)	�����#�L�;��7U�}�k���{��r������|-x�Vk��>\��<M�[V>��/��#�ws�����Ru޽�Ƚ|���Q�����Ž<۽����^����ا,���;�̕J��wY��Fh��u�W'�����.|�sm�ӱW���>���&�e��F���������0�BK���e���{�愾�O��Km���c���>s���d���U��QG�jK8���(��b�9 	�����{��߽$��M������+��)���:��dK�[�Zcj���y�+U���������PÎ�t�������l�:�S��=�0].�)���.� �>���U�#Dp�V����5��!���L?��Q��"��*����)y�=}j���[�yL��}<��l,�Χ�����
��Y	�����	��S&� $7�ջH��Y�bj��y��y��3���~��IO���D���1��������:��>\h�yT�\�H�$G� OP���b��7{�����|���)��񳡾�Š�|M������42������~�޵n��^���M�.=�~C.�z�"�����D���!�v,���:��0K�j�[�Ql�Q{��"��ͩ��G%���暾����� ���2��<Ė��ċ�h!~���e�W\S���I��)K�?W��ok�j>��jَ��F��l֟�Zա�����8[��^m�����������<z���j�f�Z�UJ�N):�b�,�v#������ ��9(��{4���C���T��ie�Q^u�Q���ۉ�Xw���ޘ�H.��#���'��Ở�o����:��h{��Kd�^T���N�_�S���b�7%y�fi��=���ڞ��  �  =O�^�V�o�Z�h)\��F\� �Z��>W���O���C���2�����0�M����W�
Bܽ~}�:H��o=�F3%�r8��mH���S�S�Z�a^�m8_�9_��w]�9-Y�r�P���C�ٮ2����������R���⽊��������:�*��=���L���W��]��r`��Sa�b�`��^�E�Y���P���B�L�0�N��5
�9�������,������l[.�z|@�Y�N��BX��]��_�n6`��v_�.�\��^W�ŏM��$?��-�I����H5��Ӷ�ݚ�{B �ë��$�;:��M�Ϸ[���e�Pk���m��sn�U�m�Vk��re�s([��KL�:���&�]��T�	�����������#���7��|L��i^�\�k��t��By�`<{� �{��z���w���p�"�e�M0V�_�C��p0�$��(���-����}�!��p3�h�G��4\��um��"z�������K惾� �� d�������{���o�f�_���L�M�9��=*��L �G��:�#��1�wnC��$X�l�P�|��L���Hǉ����O����������4���&|��k�FY��F�::8�Z�/�*�.���5���C��V���j�z�}�7��������
��m���ΐ�J����f��Sӌ��*��%��P<p��<\��<I��B:�S�1�s@1���8���F�9�Y�=nm�A��U��kߋ�w���{Ə�����ŏ������ċ��Ԇ���K�l��X���F��8�Þ1��2��;���J���]���q�ځ�����L:���������>���˘��!3��P"��ֆ��l~�ݳk���W��4F�mc9�i�3��6��<@�^cP���c�O�w�ԁ��f ���%���U���<��me���⑾�E������0���s~��`k�y�W���F���:�l�6��S:���E���V��Yj���}��L���  �  ]|/�ѯ>���M�<]�e�k�v�w�iE~��}���r�]�_���G�cr.�Ξ�0L
��&����S����4�ڔN�_*f�~w�������w�-^k���\���M��?�( 0�C ����+����w���Ƚ�ݺ��a��������ս���M7	����_*���9�s�H�{�W�sg�~�t�f[�
����#�n�q�N�\��XC�߇*����Q��
�g���'��"@��pY��o�Me}��S��A��Iu�W�g���X���I�|�:��l+����(�ΰ���z۽"Ƚ�k��^�½ 0ҽ����	��x)��u:��J��3Z���i�y�9<��˶��]�������sz�/d�<*K�C4��#����{� ���.�o&E�HZ_�<�x�������:��5���<	���~�@7o�P`���Q���B�)�2��"�/a����t���s���  �ZM	�����w'��9�)7J�Z� 	j�6\y�K[��X�������K��]��������X����t��2\���F�QP9���5��n=���N�)�f�����Ȍ�=ĕ�Y���_����������i��K����u�Zog�OfX���H�K9�x+�47 ���@��32���)��d8�II��4Z�K�j�3Jz������)��4����������ڞ��Y�������獾z;����i���U��8J���I�d�S��f����?�����Y�����o����������sG���ʄ���z�Hhk�3T[�ϦJ��h:�T>,�Y�!����s��$���/�<�>�2O���_��	p�t[��3���Ɏ�:B��"Ӝ��0��"���qR���;��iՊ�1|���d�R|S��K�4�N�ˈ\���q������ �����Wۡ����*R��밚�|����*�������z��6k���Z�OYJ���:�Ʃ-���$���!���$�
-���9���I�ۗZ�D:k��  �  p���d4���N�шk��	���P��*T��j2�����>Ӊ���t��(T�˾7��%���� {(�9�=�,\��T}�p���Q����c���-��>+���d��T5h��)L�R�2���I�G���YϽ�2��Ė������#���M�����c�Ľ�a��U�j8�r�)�qB��Y]��8z��芾����@	��*���-��1'��en�p�M��4��L%��s$���1�>ZJ�S�i��<��;���C���y�y��Bԋ��d|�L|_��D�ie+���N��T�\gɽ�a��9����|������C᭽3P½�~ݽ�����i�5	&��;=��KW�b�s�䈈��ו�ˠ��6ѣ��3������y߉�_ms��pU�Ý?�*6���:��SM���i�ƅ�%ꕾD��6���/ħ�����-����	����q�KW�	�?��+�s��6R
�l����1�W4۽y�׽��ݽ͂�=a�j���3 �b�2�kH� �_�$�z�쥋����A��1Q��DD��xR��P3������f���S�3O���X���n�񆾂㗾=��͝����������Ω�m4�����%@��#fi�?mS��V@��/�eh!�F���e����q��F������!��r0��hA�1�T�Bj��=��1َ�r:�����鵾j廾Q���ܳ�~Ħ������q����r�2d��Sc���p�n���~z��T¤�E��V]��A���aC��4��� ��R��� ���`k�f�U�J�B���1�ؓ#����Y�����F��������5'�Z6���G��{[���q����C����2���_���
��A��@U���찾Ø��o/���邾Ieo�^Ke��li�a{�-s���⛾����%�������ǳ���p�����#����i��,����h��5T��B��%2��$�z<�+���'�JV����d;$�"�1�T�A�$�S��  �  ����4���Y�\S���镾�ʧ��س�������)D��+��$wy��V���>��8���B�V�]������C��.���v쑸��������D咾7�|��bT�*�0���������ͽ�o���}��ќ�������|�Y���}��k���u��_��p��$��E�Fl��̊��ƞ������p���	���v���q��a\��s�p�|P��:>��0=��M�,Sl�3䉾A ��໮�4��t���� ��	[��̝����o�#�H�7�&���
�����UŽ�b��s���;݊�h4���$������>P��A��86޽9����p:�1^^�(g���c��Z���Q����������C~��p���1�����u�U�Z���N�jYT���j�/ �������믾�𾾨�ž�þ9��������H��W�}��tX�j�8�����:
��i��nBܽ�i˽�����~��,�Ľ�"ѽX�佼-������%��@�_`�P����:���ث�������ɾ��;�?Ⱦ����m§�a����"��o�m��yg�Ls��8��Q\���]��R¾1�ξF�Ҿ�Q;���˦��M0��	T���kg�7�I��I2�r��aX����g���Ț�����, �ij���7 �22�ȫH��ld��/7���窾@ξ���ξJؾe�ؾ�$о���M髾ԗ�ȵ��}}�J|��5��ڜ��7^�����qLξ*�׾jIؾ��Ͼ�2������-ȗ�0K����f��J���3���!������	� ���8��� �K�?�BV�nP&�
p9�-qQ�^
o��0��f/��� ��Rž}nӾ"ھZ�׾`̾����(+������*����}��m���Y�����/$��
�ž�lԾ�۾4�ؾ�t;�8����t��pĀ���a�YrG���2��"��a�O�(��~�����0���!���1�n�F��  �  ���:��h�1���8V��S���"�̾�	ҾX�˾@�� 夾e���q�o�	nT�nvL��DY���x�p��+Ѫ������ξ��Ҿ�˾j���B3���[��ǩ`��4������g���c���ʆ����m��3^��[�9f�R~�&H����WHԽ�����$�A�M�7�}��Θ�gѱ�13ƾ�?ҾxuӾ3�ɾ񔶾_՞�*1��L�h�LS���Q��e������⳾��ǾݒҾs�Ҿ��Ǿ��8��o?����Q�=(�J���1ٽ���c-��q���G�s�D�k��q��L��+��⪽�̽)K��� �w�=�*�i�4���+���@��5hҾ�6۾%�ؾt�˾����= ��Ȉ��?q��c�Ԟi�(������c8��/�ƾFeؾYX�K�ܾ4Ͼdu����x���5�^�w�7��#����&��ɽ�L���ְ����ݳ�&;���ѽG��H������>���e��ቾ����1H��ԷӾ� �_�m����Ѿc{��뒣�y���E����{�C���0��������þm�پ��Q��'��'վ�轾�B���p���0k��SG�>h+�	��$��Rp�����罊 轥���5���L����*�@�C�fe�����
��績o�Ѿ�!��h6��-��/־�a��O���U���x����`������+��	l���dӾ^羍0�FD��Z�u�Ӿ����-���눾&h��@F��,�p�6/
�uK �k>�������c������G��z�ND2�aBN��r��Ў�޷�������پ�뾼`��U��a���Ͼ�d����󀐾�����P阾�K��isž��ܾ���������l�㾣1ξFǴ��0��)����`�	�A���)�La����9�A���T<��Mi����~����5>)���@��  �  Ƿ�"�?���s��ؖ�o��]q;�޾���ژݾQ�˾Ig��/���6�����b��Z�4h��j��>䝾t鸾@ѾR�xa�@�ܾ�ɾ%���ב��k��*9��^�������!ۑ�Uyv��Y�%IK�YI���R�=�i�/�������-,ͽ��rR'�[wU��܅�%9������U�־�k�v���ھ�žYt��zF��ߴx�
a���_�Y�t��~��G��J�¾ݭؾ{��h��=]ؾ¾������=NZ�GU+������ҽ>y������=u�u�`���Y��_��Jq�����5ܠ��<ý�����E�A�cs�W���³��Ͼݤ㾆���A�ܾ'bž,Ī��"���;���p�&�w�f��`H��'f��Vy־��j����޾0�ƾɿ���ό�Je��9��P����K\׽޽��I��O���Υ��e��M���[ǽ��x��`��`�?��mk�aď��Ŭ���ɾ�i�n�������.����ᾒ�Ⱦkt��E����Ȉ�������樝�:y���ѾV����U���1���^�ɾ��������7�o���G���(�,�Ep���i��1޽��޽� 彏��g����l�&�ªB��g�抾���Pþ�߾���� ��������wi���ʾ2ư�?ћ�{����I���晾��`�Ǿ�W�;���I�E��������ž���'���#k�oiE�6�(���Q�xe��g��EE��潑!����n��H���[/�u)N�&v����;ү�N;�s������f�^�#P��o�ݾ�"þ)D������!9��`�� 鷾�ҾC`쾫���-���[��?۾�k��Jm���1���b�W�?�>&�*y�E��.d��������;��+���U�����+%��u>��  �  ur��BB��Dx�hH��Q���&Ӿ)/�9�- ��<Ѿ�7��Z���8�����g���^��wm�b���|����O�־<�羅
��D�G"Ͼ���������n�q%;�����[� ��Ǝ��p��S��7E�C���L�}^c�H̄������?˽�e��(�ЂX�~�������ľ2�ܾ����)��>˾v�2ڔ��k~���e�5�d�;�z��������,Ⱦ��޾r��7w��q޾
4Ǿ��+_���]��,������н���>���9�n��iZ���S��+Y��"k��~���ɝ�����~(�>�[sC�^#w��!��e���pԾ���'T����2�⾰�ʾ��rr��cꂾ�~u���|� b���
������ܾ�f�W}���L�����JG˾�R��f/���g��{:�3��+v���lԽ����d���B���Ӣ�]���%���(Ľ
߽���2H�;�@�O�m�#���4��Ğξk龀0��� ��4��g����;KQ������R���
��ᣎ��ݠ�n���k�־8𾶙 ����|��C�龵4ξ㯾���q��H�+(������ ���콭m཯۽&�۽���ͷ�9��i�x�%���B���h�#k��Q����'Ǿ9��:����h��$�^^ ����}Ͼ�Y��o���>j�����������l��+"̾���`��������/����b�ɾ I��(����l�BnE���'��`�9w�6/��g�bB�q�����������X��.�UrN���w�n����ٲ���Ѿ���e��F��(L��L���㾞OǾ���Oʚ��Y��һ��$^��쭻��^׾����8a�S*�������t���	̣��~��icc���?�/�$�4������4����ａ����������w��$��>��  �  Ƿ�"�?���s��ؖ�o��]q;�޾���ژݾQ�˾Ig��/���6�����b��Z�4h��j��>䝾t鸾@ѾR�xa�@�ܾ�ɾ%���ב��k��*9��^�������!ۑ�Uyv��Y�%IK�YI���R�=�i�/�������-,ͽ��rR'�[wU��܅�%9������U�־�k�v���ھ�žZt��{F���x�a���_�^�t��~��G��Q�¾�ؾ���y��S]ؾ-¾���8���kNZ�fU+������ҽ�x������:u�a~`�Y�t_��Aq�줈�+ՠ�[4ýE�����.�A��\s����1���
Ͼw��\��4�ܾ͂"`ž�ª��!�� ;����p���w��f���I���g���{־��y�����޾ʃƾXé�Vӌ�uPe���9��U�����-c׽þ��L���P��%ϥ�]d���I���Vǽ�I��a����?��gk�����I¬� �ɾf�����V���Q��S�ᾚ�Ⱦ�r��J���Ȉ�
���v��󩝾�z���Ѿ�X����\X���5����,�ɾw���E�����o���G��(��0�Ot�q���㽶޽��޽�#彼��8�H��ك&��B��g�$抾���	Pþ�߾���� �������xi���ʾ3ư�?ћ�{����I���晾��`�Ǿ�W�;���I�E��������ž���'���#k�oiE�6�(���Q�xe��g��EE��潑!����n��H���[/�u)N�&v����;ү�N;�s������f�^�#P��o�ݾ�"þ)D������!9��`�� 鷾�ҾC`쾫���-���[��?۾�k��Jm���1���b�W�?�>&�*y�E��.d��������;��+���U�����+%��u>��  �  ���:��h�1���8V��S���"�̾�	ҾX�˾@�� 夾e���q�o�	nT�nvL��DY���x�p��+Ѫ������ξ��Ҿ�˾j���B3���[��ǩ`��4������g���c���ʆ����m��3^��[�9f�R~�&H����WHԽ�����$�A�M�8�}��Θ�gѱ�23ƾ�?ҾxuӾ4�ɾ򔶾a՞�,1��Q�h�RS���Q��e������⳾��Ǿ��Ҿ��ҾșǾ+ﳾ�8���?��3�Q�W=(�]���1ٽ,����+������c�s��k��q��C��춒�>ժ���˽\8������u=�t�i���@$���9���aҾ�0۾��ؾ��˾���@���kƈ��=q�}c�.�i����������;����ƾnjؾ6^ྵ�ܾ�ϾQ|���#�������^��8�|-�-��:4�ɽ�S��Dڰ�f���ڳ��4��F�ѽO��)��e����>�'�e��ډ��{��A��ѰӾ7��3����2�Ѿ�w�������[���5�{�L���3������u�þJ�پͯ辴����`վE�J���w���=k��_G��r+�3�����{}��٧��罇'���:��/N����*���C��e�����
��績r�Ѿ�!��j6��-� 0־�a��O���V���y����`������+��	l���dӾ^美0�FD��Z�u�Ӿ����-���눾&h��@F��,�p�6/
�uK �k>�������c������G��z�ND2�aBN��r��Ў�޷�������پ�뾼`��U��a���Ͼ�d����󀐾�����P阾�K��isž��ܾ���������l�㾣1ξFǴ��0��)����`�	�A���)�La����9�A���T<��Mi����~����5>)���@��  �  ����4���Y�\S���镾�ʧ��س�������)D��+��$wy��V���>��8���B�V�]������C��.���v쑸��������D咾7�|��bT�*�0���������ͽ�o���}��ќ�������|�Y���}��k���u��_��p��$��E�Gl��̊��ƞ������p���	���v���q��c\��x�p�|P��:>��0=�(�M�@Sl�A䉾S ������54������� ��M[�����4�o���H���&��
�"��kTŽ/`���򖽣׊��,�����؍��5@�����!޽�+����_:�2L^��]��BZ��֚��.��A��������w��	������u��Z��N�L[T��j��#������������ž�þ����u���QR����}�`�X�>�8�z��zF
�}���Pܽhs˽�������Ľ�ѽ���:�������%��@���_�ݡ���0���Ϋ�Ƶ��{�ɾZ�;8Ⱦ����*���m���\ ���m�!zg�-s��;��{`��Jc��!¾#�ξ3�Ҿ�[;�����y:���]��0~g��
J��X2�����c�'��ߝ��L�������/ �cm�N��9 �;32���H�md��C7���窾Eξ���ξJؾh�ؾ�$о���O髾ԗ�ȵ��~}�K|��5��ڜ��7^�����qLξ*�׾jIؾ��Ͼ�2������-ȗ�0K����f��J���3���!������	� ���8��� �K�?�BV�nP&�
p9�-qQ�^
o��0��f/��� ��Rž}nӾ"ھZ�׾`̾����(+������*����}��m���Y�����/$��
�ž�lԾ�۾4�ؾ�t;�8����t��pĀ���a�YrG���2��"��a�O�(��~�����0���!���1�n�F��  �  p���d4���N�шk��	���P��*T��j2�����>Ӊ���t��(T�˾7��%���� {(�9�=�,\��T}�p���Q����c���-��>+���d��T5h��)L�R�2���I�G���YϽ�2��Ė������#���M�����c�Ľ�a��U�j8�r�)�rB��Y]��8z��芾����@	��+���-��3'��in�v�M��4��L%��s$���1�VZJ�s�i��<��X���j�����y���ԋ�De|� }_�)D��e+�5����R�Xdɽ0]��T���Xs�����Tѭ�\<½�fݽ�����X���%�5'=��5W�O�s�-}���˕������ƣ�c*�����؉�[cs��iU�ޙ?�.)6��:�/YM�\�i��˅�o��L�����ϧ�&����������q��`W��@�Q�+���^
�c���>署:۽�׽f�ݽ�w콲X����% �O�2���G�`�_��jz�ݙ���百�5���E���9��?I��y+��a���ꀾ�f�}�S�G3O�
�X�{�n���� ꗾg��`���m�������Tک��@��1"��&L���|i��S�wi@�3�/�Dv!�����o��������J����>�!��t0�&jA��T��j��=��Iَ�~:�����鵾o廾Q���ܳ��Ħ������q����r�2d��Sc���p�o���~z��T¤�E��V]��A���aC��4��� ��R��� ���`k�f�U�J�B���1�ؓ#����Y�����F��������5'�Z6���G��{[���q����C����2���_���
��A��@U���찾Ø��o/���邾Ieo�^Ke��li�a{�-s���⛾����%�������ǳ���p�����#����i��,����h��5T��B��%2��$�z<�+���'�JV����d;$�"�1�T�A�$�S��  �  ]|/�ѯ>���M�<]�e�k�v�w�iE~��}���r�]�_���G�cr.�Ξ�0L
��&����S����4�ڔN�_*f�~w�������w�-^k���\���M��?�( 0�C ����+����w���Ƚ�ݺ��a��������ս���M7	����_*���9�s�H�|�W�tg��t�g[�����#�q�q�R�\��XC��*����	R��
�{��3�'� #@��pY� o��e}��S���A�|Ju��g�{�X�f�I� �:��l+�����'�u����u۽EȽ�`��S�½ҽ�i�j����be)��`:��uJ�Z��i�u�x�m/������������fbz��d�KK�r;4���#����� ���.��/E��f_�-�x�>����͌�F��󟋾b��G&~��Po�p�`���Q���B���2���"�`k������� �� �G	�����j'�M�8��#J�iZ���i�ABy��M��դ��Ǯ�����񇔾�{��/P����t��(\���F�M9��5�rr=��N��f�F����ь��Ε��d���l������횐�gw���,��`�u���g�<{X�J�H� .9��+�
B �W%�.���7��)��g8�wI�w6Z�I�j��Jz�ک���)��C��� �����������Y�������獾};����i���U��8J���I�e�S��f����?�����Y�����o����������sG���ʄ���z�Hhk�3T[�ϦJ��h:�T>,�Y�!����s��$���/�<�>�2O���_��	p�t[��3���Ɏ�:B��"Ӝ��0��"���qR���;��iՊ�1|���d�R|S��K�4�N�ˈ\���q������ �����Wۡ����*R��밚�|����*�������z��6k���Z�OYJ���:�Ʃ-���$���!���$�
-���9���I�ۗZ�D:k��  �  =O�^�V�o�Z�h)\��F\� �Z��>W���O���C���2�����0�M����W�
Bܽ~}�:H��o=�F3%�r8��mH���S�S�Z�a^�m8_�9_��w]�9-Y�r�P���C�ٮ2����������R���⽊��������:�*��=���L���W� �]��r`��Sa�c�`��^�G�Y���P���B�P�0�S��5
�K������&��V��)�����[.��|@���N�^CX���]�Ƽ_�-7`��w_���\��_W��M�I$?��-����V��8-�����*��9 ������$�A:���L���[��oe���j�	�m��Xn� �m�=k��[e��[�V:L���9���&�����	����w������#��8�)�L�4}^��l��t��\y��W{�h�{���z�٪w��q���e��AV���C��{0�o�����.�W��̼!�ff3���G��#\��am��z����t��]؃���uV��E���\�{��o��_���L���9��6*�HI ����	�#�71��yC�T3X�,(l���|��X�����IՉ�o����������L��7A���<|�p�k��$Y���F��E8���/�j�.�j�5���C�-�V��j���}����������
��6m���ΐ�V����f��[ӌ��*��"%��W<p��<\��<I��B:�U�1�u@1���8���F�9�Y�=nm�A��U��kߋ�w���{Ə�����ŏ������ċ��Ԇ���K�l��X���F��8�Þ1��2��;���J���]���q�ځ�����L:���������>���˘��!3��P"��ֆ��l~�ݳk���W��4F�mc9�i�3��6��<@�^cP���c�O�w�ԁ��f ���%���U���<��me���⑾�E������0���s~��`k�y�W���F���:�l�6��S:���E���V��Yj���}��L���  �   M|�6Z}�~�v�'�j�S\��fM�d�>���/�� �����W��a�߽��ƽ������O����̽��罊������b%��5�1D�NLS��zb���p��|��ƀ�p�~���r���^��EF��.-�bR�8��)	�����#�L�;��7U�~�k���{��r������}-x�Wk��>\��<M�]V>��/��#�{s�����`u޽�Ƚ����p�����Žq۽����� ��*�,��;�P�J��xY�\Gh�Ǩu�(�D���E.|��rm� �W��>�D�&�|���A��~�[x�E�0��3K���e�w�{�4ۄ��C���`���V���$s�\{d���U��;G��78��x(�1U�������s�4�߽��位���h��R�]�)�# ;��yK�z"[�||j���y�ab����������Ύ�+~��2遾�l�ڷS�;�=��`.�^)���.���>���U��6p�㒄��+���}���2��,�������񃾤y��dj���[��eL�>m<�C_,�������
��Y	�4����e^&��17� �H�b�Y�gj�M�y�N���A�������\���Q���=��𨕾F$��>B���ih�L�T�Y�H�8G�sTP��b��:{�����1��*��9����Š��M��Ю��A2������~��n��^���M�3=��C.�}�"� ���D���!�v,���:��0K�j�[�Rl�Q{��"��ͩ��G%���暾����� ���2��<Ė��ċ�h!~���e�W\S���I��)K�?W��ok�j>��jَ��F��l֟�Zա�����8[��^m�����������<z���j�f�Z�UJ�N):�b�,�v#������ ��9(��{4���C���T��ie�Q^u�Q���ۉ�Xw���ޘ�H.��#���'��Ở�o����:��h{��Kd�^T���N�_�S���b�7%y�fi��=���ڞ��  �  ������������4���j���M�J�3������t���ν�|��A �����Ot���N��z���ώ���b׽b��$��~�#�R�;���V��Ws����-v��[����C����Q߈��1r��Q��6�v�%�c�"���-�UE��%d� ����ʐ�J���Hr��� ��/L������be�ۓI�l0�_F�6���I�SyͽQ���h���֙��9������7��Źɽ+��f-��;�0�,���E�ua���}��P������������7���2���g���H��U1�s�%��D(�o�8��`T�)v�����#������xU��XV��%d��E����i��ZN���6���!�a��������
Zн�ý�m��B�½�Iн�w�� �O���A#���7�;NO��i����]����L��@6���B��@q��D7��ņ��#�z�L�]�d�I�vB�p�I���]��{�͎����������!������显�ʊ�Lgy�Z�_���H���4�|�#��}�4�r����Z�����9����e���0��AC���X��$q�],��ʶ��좾�̮�,���"��[N��w���6M�������r�d"c���`���l��5��Y�����������?5��c����c��D����=���Œ�Ǆ�S5p��Y�<F�p�4���%�����������_����+�#��z2�*fC�F�V��ul�멂��z���랾}j���ɶ��ܻ��9��Sϱ�����Ǔ�w��~�o���c�|?e�/�t�3����ʗ��㧾�����Ȼ�v���V���q��補��N���Հ�)�i��T���A���1�R�#����KY�&4�	���r��3�|1,�0�;���M���a�j�x�/\��3�������������������Ū���J��hh������2����o��h�O�n�-��ȡ���0��l�������  �  ��������������=����W��\3��g��T��Uν.i��-U��/Z��`�v���q�/Z{������ל���ٽx����U=��Ac��K����������n���򼸾��������f ���u���S�9#?�2G;��I���e�FH��К��d���V���c��fN��ڼ��/�����w���O��-�������9%˽�ѭ�ϗ��Ո�.����x��bL���D��C��)�ƽ���(D�D�(���J�O�q�.������tX��`f���t��Ĉ��s�������|Hj�G�L�>��A�CU�vHw��t�����1u���(��������裾|���!w�*Q�C~0�{���R �UG߽��Ž:��fH��uߥ�멽+L��)�ǽ�3�^� �ׇ��.���M��wr�ܖ���`����G7¾�Ǿ�þ�1��餾����T�|�!�c�n�Z�1sc��v|�����ҧ������ƾ�S̾dnȾE���g��P���	����_��`@��t'�����u�j򽉑�@ڽ�Pٽh�߽����*���g� �9�6�R���r�q����Z��ѵ��ǾSҾ�Ծ��;���ug��菱�9����|��y�e��������6��q溾��̾��׾ëپN�Ҿ]�þP����ߛ�������l���O�z�7���$�`�O�
��c�4���6I�����@�	�&��\"�G�4��K�.h��?��a☾�����<��φо��ؾ��׾��;ż�/q��y۔��υ�(6|�%I~������,���]��ea���Ѿ�Fپw:ؾjξ����G����Y���B���c�}H���2��!�F?�>�
�im�p�� ����F��2���+�]�?��X��Nw�Gɍ�����϶��[ɾ|�־z�۾Z�׾�A˾3ɸ��H���ܑ�L��T5��k:��f��̀��S��',ʾk�׾�  �  �Ѿ̾�p��F㥾H7��j�e��t8�������o�����4����f�0U��P�?7Y�%�n�a����ࣽ�OȽ�5��qo�&8D�=Es�sn��HାX¾$о�3Ӿr˾/s��:���I���l�2VT���O���_��ꀾĶ������w�ľg�Ѿ.�Ӿ�jʾ6��n����	��2�Z�x�/��u���8���rU�����V�n���`�p�_���k�ߚ���Ȗ�����۽�A�k*�;|T�����{��m鴾ȾlmҾ�Ѿk"ƾ�1�� K���b����c��}R�C�U��Um�����'	���X����ξՌؾp>׾�˾E���HƝ����=�X��0�y���C�"$̽}�����������d��?3������Xմ���ͽw!�G���,��8R�	N���H���g?ʾ�ھ	��(�ݾ��ξpC��s>���Ë���y�7o�y�j-��0֠�Ȇ���bо����i���Ѿ<����f����0d�ׯ>�0!�_�
������߽'�н�~ɽ��Ƚ9�νD�۽�5�W���o�Ru1���Q���y���������Ⱦr�ݾh�뾕ﾺg�4D־���c%��i����������js������﬷��о�侷���󾀰�~Iؾ+'�����HW���so��L��o0����\Q�����;���1� ����B ��j
�U����,�ӧG�3�i�9��&��������վ>J�������X�|SҾ�I��9.��
y��ok��ߠ��_唾�9����ٴ׾�H꾧��s��pl���о����i蝾+����c�	�C�8�*����W�
�Ia����zD�V��f���^���x�'�"�r 9�ifV���{�~/�� v���eǾ^�޾^Sﾺ5��D����.";�崾-��~��Sh��p��nf��]����˾>�ᾡ��  �  ��شݾI�˾Ud��rG��)q��=���A彘$������q��R��(B� >�>F�Q�Z��m~�� ��;������^D���J�����D�����8uҾp⾇�従�ܾNɾ�J���Ĕ�t}���b�7z]��@o��_��Ǚ�����h�վ�㾱��;�۾éƾ�\��*��d�R3��+�0�۽󒯽 ���u���Z���M���L��7X���p������x��b�Խ[����-�& ]�����w��8-þ��ؾ(��n侂(׾�����m��R	��=rs�� `�=�c�Ԋ}�I���-���c�ʾ��߾��꾹V龠s۾PAľ�����劾eO`�X3�*P�*��\�½�@��$���$}��
���Ï�f�������&�ý��;k�j;-�c1W�'����V���پ+z�=i��[��T߾7Ǿ���������W��R�|��Ѓ�*꓾qӫ�G$Ǿ�|����j1������Ⱦ����
\��n�i���?���������Խ��ƽ���}����gŽ��ѽ�佷� �a����/�b�S��O��0�� V���KվW��Q���w� ��	������̾񪲾.��f��	����(��
)����þM�޾$���X�n!�����\�澺�˾i	��a ��fLs�]�K��i-���V7������l���佝N佀��O��?J�v\�O�)���F��Nm��r������ǾkT�w)��~�}+��e��#ᾔwƾ�ᬾ%N���M���������p����̾��<�����E�����_Y޾+���ѱ���؉��?f��%B���&�n*��g�ܡ���G����뽆	������o�m����6��V�?�� ����#��ˇӾ���i ��Y����D`�$۾�5��$+�������5��Fe���,��Ӿ��v�ؾ@�񾵵��  �  ��<�B67��9'�q��0v�~˽�م��h�b��.�� 	��Aݽ���S좽�Ӗ��ȓ��S��d,�������� ���:���r��a��Muɾ�,��)��	Z,�$c:�r�=��{5���#�@����0�ž�خ����s����پ,���?��.��;�ĥ=��'4�}t!�Yi	��(�W5��.���%VT�U=%��V��׽�^����������#��2�������~ҽ/��� �<UM����6�����پ�&�c�P�1�t�<�?<��I0�b������ݾVI��ҭ���P���þ��I��ds#�ET6� @�r>��1�����!�_f־���u􄾩Q�J%'�f�	�Լ�ҙҽ[�Ľ����^-Ž��ҽ9V��U�U�!��(G�B3z�;����:Ⱦ��������,�.�=��E��@�*�1��Z����?i�N?ľ�ٹ�?�¾��ݾ�i��-���1���A���G�"�A��2��[�����Ӿ�a��,l��*<[���5����!�
��2 ��������<!���e��-���(���F�T0p��%��g^�����*�VV$��:��7H�S�K��C�Hj2�G��a��\�侈:ξ�WʾZ�پ*��������*��.?�OL���M��xD��1����]D ��xѾ-���w4��e��C�P`+������(�[�����q��C�(��?�D�_�Ȗ��.
��h�˾R���U���.�BB���L�ZXL���@���,��*�����ugܾ�w˾��;;��ڧ�1��y�1�GQD���M��K�H�>�\�)���\E���þ秞����	�Y���;��e'�w�3]�Ta�?�����
v!���2��|L�i9q�nᑾ�)��6�ܾ�~�3���,7��-H�NJO���J�*�;� M&������n׾��̾Cuվ�8�.e�<�#��,:�UJ��  �  #-7�o�1��Z"���t��5,��)�����a�e�/���
�����E������?��# ��dʝ��׬��ƽ
��Kf��5;��p�)!��hžu������K'��4���7�
0��q	���l�����^妾�V���'Ծ�9��J��&�)���5�-�7���.������^5۾93��D����S�"D&��>��Eܽn��d���� ������㺧�����] ׽N��Y-!��M������ᨾ�&վM���	�M�,�p�6��D6��+�{���V��ؾ� ��Z�������c��O㾸����C�0��V:���8���,����6� �&#ҾO��6���2Q��(����p��K׽�Xɽ�Ž"�ɽ/4׽�	��	�u�#���G��8y�М���ľ� ����0(�pw8��K?�;���,��,�ؓ��Z۾%7���4��#⾾�پ; �C�ˡ,��<�\�A��^<��'-�&x�C���P�Ͼ<|��#Ն�1�[�/�7���.����mf�����
G ����Z��i�*�PH��mp��H�����!{�z��4 �d�4�z�B��E�G>���-�;�������߾Q_ʾ�ƾ3eվ�r��mX��)&�|�9��UF�/1H��?��+-���c����vξ0@��󉾩!f���D�y�-����*��W����"�*���*�/A���`�p���ģ�nɾ�f������E*�x�<��.G���F��Z;�I8(�8���a��&ؾR�Ǿ��ɾq-޾,� ����$-���>���G�}F���9�Ŀ%�����뾴���������~>[���=�Ž)�}j�Z������������#��5�?N���q�g���l��hMپR�����f2�˫B��xI�&3E��6�  "��j�����eӾ�ɾ�Ѿ�N��3	����<5���D��  �  &'��]"�A���Ӛپ���������_�՘2�����3�BPͽ������_���-���>���}�ս����R=���m�������΁�jT��q�o)%���'�e� �k������=�Ծ�����)���w���r��ž���ʰ	�H��8&���'� ��f�j�����;|p��Oτ���S�'y*����&�%̽�oЭ�j'���뵽W�Ƚ��D�:�%�֓M�ှ������ȾL��!��F$�X'��l&�[t��|�W��Ⱦ�髾=��������Ӿ�=��]��:"�yc*�G)�ׄ�i"�X��%�ƾ4-���끾X�R�X�-����Ѐ����Y^׽��ҽ�I׽R�彂������|�)�\IK���w�+����໾��例����^V)��E/���+�,��%����#;�Ѵ��߫�����.<˾y������C�,�O�1�-����>���a�-�ƾkآ��܅��^��v=��_%�����	����G�B4�����m�1��pM�w|r�|���	t����վ]���F��N#'� �2���5�� /�|d ������Ҿ�t���(���uɾ^很�����+�8�6�(C8��X0�� ��~��Y�ƾ ���P퉾�Uj�]vK�u5��m%��K�/�T���:���#�]o2���G��ce�ٴ��=栾��� �辏�	����i.�zR7���6�;�,�Q��՘����i�˾gC���.��?hѾ��@K��+ ���/�F8�r6�ү+��-��R���ྶ�<���Xꂾk`���D�gB1���#�f��UZ�.�� ��U+�>]<�1hT�Xju��^=��gfо������OW%���3��u9��5�!�(��|�8�r��-�Ǿ����4Lƾ�zݾ�B ������'�>5��  �  #����ی�羜�že��8�����a�{�;�R���S�e>��6н����[Ž�
�Ľ�ֽ\��c*��#%��E��`m�g����U���}ξ���6�,`��M��d������Qݾc������{���錾�ؗ������ξCY���r��A��4x�	[���޾�ڼ��k���a��
vX� 5��\����Xl罎|ѽƽCXŽJϽ��㽈K���+�0�yS��(~�J|��>j����پ�)����	�M���
�E���E��Ѿ:��c������%������3����ܾ�������!���$��
�l�����پ���������N��N�Y�ش9�b� �����l �D^������%h��r���
��6���T�$�z�֔��#���xѾ�C�	�d5�.���s�������վ<E��?ꣾ�t���$��K����Ծ����mc�����A����d������^۾�񺾕n���ӆ���g��[J���3�P�"����O�K<����+�\�+� �?��Y��&z��t��I����_Ⱦ�����/��m/��J����#j������@ھ�`���6��񄬾�ɷ��EϾ���Fq���?@ �	�!�����u���\:ݾ����톢�lC����t��	Y��^C� 3��(��O"���!���&��21�L�@�^�U�1�p�v�����u���إؾ�F���L��'��!��V ����I�	��8�=Ҿ��%����;�������پ���E��g��ky!��z �e�0M
����cҾ�R��"���p���Yl���R�m?��-1�!(�e$�g&�"�,�L79��J���a�e�C2�����a�ž}�循��F�xp�1�"���7���m���˾@��*M��ꩵ��'ɾ�~�&����\3��  �  ���t쾎8޾��ɾ�沾F���2j����m�0�O��@5�9���
� l�����Ὄ꽓;��Ͷ��6$��G<�b�W�@w�(͍���w��-Lоӳ㾰��4B��<��hӾ/ع�0���a����y���t�!������*Q����Ⱦ9�߾���:�����xھx�ľ٬��A◾�����g�0�J�9^1��V��C	��d���K�wi�M����3����R.�>�F��cc�-��)픾�c��~`��H[׾y���U����U�˾m谾����Q���Fw���z��'������d��վ1�꾼���;����T�q�پ�þoƬ�����o���E�k���P�7�8�U�$��A��M5�U
����p�"�u�6��jN�bi������|��󏩾�񿾂 ׾k 쾇���3 ��L���龝�Ѿ�U��d�������4 ��̌���a���趾��Ѿ뾒z�����Z� �q�󾙦߾��Ⱦ�c���S������{���a��wK���8���*���"��!�{#&���1��B���W�=�p��]���W���������ܒԾ�뾧�����)����:P��P׾�Ž�ҭ������왾���˥���ξ5a��F �����	�k�����u>律ξ0$��U���zoR���	q�<�Z�N�H�P�;�ej4���3��(:���F�X�וm�UN��������7	��|�ʾ������t���������� ���?.Ѿ���nФ����QQ�������y���o׾�n��)�� ��+M����Bnݾ��ƾj���1E��{i��Ę��Sk��\V���E��;�eR6��S8��@��@O�ugb�Wy��ԉ��ܘ�0��`&��>zԾ��뾜Q �����k
�nP�`������	˾�k��g���뜾e ��7x���ȾB4�}�����  �  )�¾f�¾��x���s��Yԛ�����Lo��Ԣs�x$[�GB�	#+�a�tt�	��������0���H� b�7�z��򈾬8��w����}��, ��|g���Jž�þY������j#���m���:f�v?R�Z�N���[�V�w�с��Ȫ��,�������n#ƾsľMx�������󥾂g���1��^܃��o�-�V� A>��(��2�����5���u�%�";���S�"bl�����^���z���棾1���3����¾edž�%��Y���0V���}��Ѕ{�*_��Q�GT���g�-Q��H���#��p����Ⱦ
�˾�Ⱦnn���O��宨��f��z]������mv���]�0�F�ڿ2��%�~��"��,/�kB��NZ�_$t��׆��Bw��3�Զ��ԁ����˾��ҾMӾ�̾���s�����it��[�v��<n���v�
w��KU��_խ��G��+оuؾ �ؾ�Ҿ3�Ⱦ[Q��H�������hr�������샾\�o��X���F�A�;��.9���?��qN�H�c��[|�&������������D���ˑƾ%1Ҿ�۾���t߾��־-vǾF��*X��Q����������1���"֛��Ȯ�oþ� վ��ᾠ�����ݾ/,ҾQƾ����T��u⣾����.R��l�}���g���V�|M�sL���T� �d��z�Ȃ������\���|\��#����ľX�ϾN�ھ�
��徱�ᾤ־~�ľ٥��	����-���������>��mء��s���Fɾ��پR�㾏w�DX�qپ�.ξIv¾���j���̇��'x�������w�.uc��U���N�3OQ��\��o�������[	���ާ��5��V���Hʾ־�l������ᾜLӾj���쨬��ݚ�*����܉�:����v��R�����'Ҿ����  �  �t��1ӣ��V��L2���@���z������	���u���ˈ�L�s��U���<�h,�\�'�5o/��^B�:F]��{���������.���楾������L���/���4���_��������χ��~q�iT�C
<�ve-�c�*��o4���H���d�⦁�� ��7~��y<��|���D��F�������dA��nۤ��1��G�������m���P���9���,�%#,�e�7�_qM���i�B�����;���ֺ��'[�����c���t���+󦾢��ћ��ڐ�������g�e&L�C�7��z-���/���>�`IW�>�u��ϊ�����У��ê�.f��⯾"I��[ﯾ9��� ��9K���薾�̈�$�s��6Y�3F�@>���B�p�R�`l�9���	��S����v��t�����������𶾿[���B��y��)���#��"�����{��+b���P�׭J��,Q��9c���}�:t��>�����l ������9)����A%���b��5���������&�������恾\Gk�:�[���W��3`���s�7ׇ�������]���ԧ��/���g�¾m�þ��þ�¾�M��$���<�����7���R҇�v�x��k�#4i��s�i��3���%��N������þ{Ⱦ�ɾ�4ʾ��ɾ�Ⱦt�ľ6��7����奾����
��[&y��(l��^k�9�v��\��&����գ��ı�������þ�nǾ\�Ⱦ�>ɾ��Ⱦ[Ǿ�~þ�;���3���)��'퓾	؅��`v�c�k�o�l��z�*���'���~ݦ�nr�����0Ež��Ⱦ)�ɾiʾ-�ɾ��Ǿc�þ���������C�������&v��Mm�.�p�b7������{�������·�Hs���dǾ=Lʾ{Z˾s�˾��ʾ��Ⱦ��þy��W��<���Q����z����v��p�P�u�����u������G����.���  �  ����ِ��>��	������#���tþ��¾����9��u ��25���<h���Q�<XK�2�U��o����)��߶��NA��`�ľ�þv�������7����a���/������7sr���Y���@�Z*�T��i�������$"�S'7��O��h��q���M-������xv��ﺹ���¾�]ƾ�Yþ3⸾�C��%f��6�F�b��FQ�0AP���_�l�}��ꑾZ٥��궾1¾��ž��¾�+����*�������r�����`j���Q��9��$��������$�=�.��]F�{`���z�����ރ��P������x︾��þ�Q˾27;��Ǿg������֕������<m���a���g��T}�JǏ����>�����Ǿ�Ѿ�Ҿ��;�oľ|	���`��������]���U���f��O���<�R0�,3,��-1�+�>���R�.+k������/���&��
��������W�ɾӎӾ�hپ��ؾ,$Ѿ��¾��������R��.z���&{�
9���x��;��������ʾ#mؾ�%߾>x޾��׾�;�¾���Ǵ��FȠ��l������H{�.�e���T��HK�BJ�z!R���a��iw����vʔ�2 ��X�����;,þ��ξھ�⾀|澎[�F�ؾ�Ⱦ�%�� �������B��`�������rr��o�����ž�־��^��I���Rھ"AϾ�zþ���pӬ��p���s��g���ȍy�N3d�r�T��L�P�M�%�W�� i��p��)��&�������`����@��Y�ƾٸҾZuݾ������9�ˈԾ-�¾�s����c����������������9���%����;�0ݾ��}��<���پ+�;����ڮ��\������i����j���:w�ˏc�$\V��zQ��U��Pb�2�u�磆��;��?����  �  ��n�%�����1���)˾�l߾s��Kc�B�l�վ�輾����mۋ��z�z}q��S���������YþPe۾���{��U����ܾf�Ǿ����p����jk���M�J�3�=z���
�����'��A�>���s�5O�td*���B���^��)��)���\��Y����ԾZ;�K��0�LH�6о;���@��Q����:x���v�ׅ�Jy��|Ѳ�:;@��p��
��-=�x־�2�����?���/р�)a��E�ێ,�^����3���+���j��F����τ#�<;�d�U��$t��[��o(��[��ٯ̾qf���������������ϾpX���0��񰋾7��g����ҕ�TV��Ǿ������ʥ������`��ݾ2[ƾM���d;���h��t�bsY�<TB�S�.�� ��������#c"�Pv2��G��G_��z�����g枾wd��fʾ�ᾖ]���v�7�o��X6쾈�Ӿdh��[��ڋ��Ȑ���՗��.������ܾH��l������:��m��%�⾠�˾-����?��N}�����m!m���W�m�E�x&9�e.2�g�1���7�TD�0mU���j�b聾^���$������i�Ǿ��޾m)������ӗ�5��y��k�վ�𻾽\��6���.���s�����x{Ҿ����\�_����\#������i�bɾ
���%���ݐ�\����l��EW�qF�:��74��5�X<�C�I�(S\���r��-��	۔����t@��z<Ͼ�k����1�Ф	�*��p����e辺�;u������'���$ޞ������¾�6ݾ.���]�H�	�(��!������ھ1Zľ9ϯ�7띾Pq������ Ij�SJV�?�F�K�<��69�aY<�p�E�f4U�i�I�������  �  cc�V���5����]ǾR 龌c����O���/�� ����	��A�����]#���Г��;��+�ǾA���lO��H�to�v���8p��=y��ǭ����]���8���h�����/jҽ��ŽX]ý��˽�߽�����L�H,��rM� 8w��T��v���(&վ
�����?���A�H
��v���Fؾ���]���]���1��}2��3���DԾU������0�������	�����@5ؾ֚���Ɨ�\"{��P�e�.�ܢ�� �.�)�ѽ.8ʽg�ͽ��۽���(�A<#�#�@��ce������;��b(žZ羿n����V�c�8
�����v=վ�s���8��~u���ʚ�����v�Ⱦ�����V@�	������h����s�ھ�幾a����(��g	a�9-B�qQ*�JQ����29��2�����C��,��;/���G�^g��1��Mw������Qݾ_����]�H������F�l���3���־�e������ᢾ6⫾Х��B���f�h���B��d�\���a�X����{ܾ-����#��-����$q��,U���?���/��5%�������\�$�N�.��C>�L�R��m��6���%���ݵ�$6Ծ�����-�x���� �=@!�i�բ����5׾�-��S���9���Rκ���Ӿ+��g�
������ �)� ����r�2f����־���ڝ�P���uo��T�
@���0�>�&�8"�K�"�P�(��A4�)�D�>�Z�V�v��k��*磾MH���޾ib �76�#D���!����b��ʼ�ʼ��ξ�+�������p�þ��߾� ���������"��> ���^�j�ȅξ2�������鄾Țj��CR�ڬ?��M2��%*��Q'�)�)�:�1���>��Q�Di�����  �  ��a��i��w�����۾�2�2�s#��c'���!����� �8�پ�P����E����夾�c��.����� �2l$�J�'�Kk!���������Ծa������5Z�o
/�R�����(ν����i%���B���˲��$Ľ�(ཛX�Ԋ �T�F�"y�yX��Oy¾e��J �Kb�y�&�M�'�q<�6'�c��X%Ͼ�&���͞��՝��b��7˾b��@��E��3'��'�U��e��F��[Qƾ�����5~�Z�J�:�#���^��hɽ{ظ��p������F�½��ٽ!������>6�;a��W�������־�� �d���H$�q�+�Z�)�ik�g��w$�H9̾B�������x��N��1�ᾑ9����w�'�Ƃ.�Ss+��q��/��E���ƾ���������X��5��/��B
�����o��Pr����d4��=�!��+;��s^������D��E�Ⱦ��5.�j	!��.��k2��-��G�M�l��oξix���I���Ἶ�־����K�&�$�jP1���4��.�J5 �O����ƾ����Ո�o3g�y�G��e1�"�!��)�l�Dd�����_!�)�/���D�g@a��ك�����ݼ���⾗���G��{,���6���7��-/�������~�Ͼ�j��	p����̾���j�����Iw-�d�6��7���-�G��r����ݿ�H[��ύ��H�c��F���1��S#��B�c$������8�&�{6�V1M���l��L������+�Ⱦ���/��}�!�D�0�'j8��66�7�*���H���k�b�ɾ����_¾v!׾����k]���#�_�2�=9���5�j�)�����w�op۾-���)}��߀�'^�8D�H�1�(%���4K�C��w�$���0�L�B�vN\����  �  ��c��M���i���o������#��k2�|k7��T1���!��9�US�E�ľ�-��E���Nk���̾d���s���/&��
4���7�s0�<���c	�9�&]���	���-[��e+�c���A�����.���e��B���-���a]��#ѽ�������jE���}�C����ξ�3������*�;r6���7��.���R���P߾ü�t�� a������B�ھ���}�LF,�F�6�B�6��,��dz�p�Ҿ펦�7ʁ���I�5���< ��Fֽqú��ꪽx	���>������]˽�j����G2���a����xĶ��b侃�
�A�!��&3�L�;�uk9���,���?.�۾>l���[���뵾�X;
��D'��=&��7�%�>���:��)-��F�q< ��1ѾX|���y����V��'0���п��A����޽���\����v��H`5�۬[�H����+��~[ҾU� �&��R�.�]j=��sB��m<�g�,������ܾs�þ����XȾ|徔�n�L�2���@�A�D�]�=��-����[4��^�Ͼv���M����c��A���)��`�8��x�J��������.h(�y�=�/\�(���K���Bþ���M�*'���:�p|F���G��>���+�$v������fܾ�ɾ�ǾaLپ(Z��k���V)��&<���F���F�	<��)��������ƾ��K%���_�g�?��Q*�����/�lS�q��Q����)/�L�F� h��x��()����о�&���f�xH.���?��^H�$�E�+%9�u%��b�A�oZվȾ�M;�h侄���P�]51�v�A�U"I��mE� �7�Ǣ"�P�
�v���������d���X�A�<�;*�]�����z�����P��I)�'�;�3zV�>8|��  �  �9e�wK���#���4�Q���p(�d8��==���6�P�&�@�j����ɾ���'����~��P�Ѿ,��j���A+���9�ԕ=�/�5�M�$�
���羞�������\���*�����۽Kc������4 ���M���:��@���v̽����/��lE����<G���}ҾX�}&�`�/�p+<��=��{3��� ��Q	�s�<��\6��������%T�����R�1�߷<� �<�DY1��i����86׾�G������/J���������ѽc��|w�������X��'`ƽ���f��_U1�;@b��`���๾�t�55�--&�T�8�ޓA��?�N�1�0!�l��]ྱ���T���ƹ��Ҿ���H�+�(�<�@TD���@�[,2��X��=�$վd����C��;DV�;�.�����f ����qݽ�ڽ
h�HQ�g�����3�o)[��U���(��\־}���� l3��C�\EH���A���1�Q���;���ྩvǾVA���g̾�'꾦]
��="���7���F��J�rC�o�1�5���?���ҾL�� �����b�Ǹ?�6�'�������q?
�bO
������&��;�1�Z��'��pX����ž���֊��L+���?�Q5L��}M�flC��0�g/�a����/�̾r�˾�ݾ����Sd�t�-�xtA�ߠL�A�L��WA��s-����#m���ɾ�7��?��#�]�_�=���'����3���%����q�������,�7�D�g�g��ǋ�ܨ��p�Ӿ���� �C�2�;E��+N�̢K��K>��p)����h���e�پD�˾ *Ѿx����z=��6��IG�3�N�BK��<���&�>�����!?���ǚ��
��W���:���'��l�����T��b�����&�Y~9���T�,�{��  �  ��c��M���i���o������#��k2�|k7��T1���!��9�US�E�ľ�-��E���Nk���̾d���s���/&��
4���7�s0�<���c	�9�&]���	���-[��e+�c���A�����.���e��B���-���a]��#ѽ��������jE���}�C����ξ�3������*�;r6���7��.���S���P߾ü�t��"a������F�ھ���}�QF,�L�6�L�6�
,��sz���Ҿ���Gʁ���I� ���< ��Eֽº��誽����:��ޓ��e˽lc�A|��B2��a��܏������^侕�
�S�!��$3���;��i9�^�,����h-��۾�k���[��O쵾�Y;v��=(�:?&�S7�Ӆ>���:�o+-��H�`> ��5Ѿ����|���V�D,0������wE��#�޽V�����������[5���[�7���6(���WҾ\� �!��Q.�rh=��qB�[l<��,������ܾ��þ%����YȾ��k�����2�H�@��D�X�=��-����h8��6�Ͼ�y���P��E�c��A�/�)�nd���^z���-����� i(��=�y/\�+(���K���Bþ���	M�*'���:�p|F���G��>���+�$v������fܾ�ɾ�ǾaLپ(Z��k���V)��&<���F���F�	<��)��������ƾ��K%���_�g�?��Q*�����/�lS�q��Q����)/�L�F� h��x��()����о�&���f�xH.���?��^H�$�E�+%9�u%��b�A�oZվȾ�M;�h侄���P�]51�v�A�U"I��mE� �7�Ǣ"�P�
�v���������d���X�A�<�;*�]�����z�����P��I)�'�;�3zV�>8|��  �  ��a��i��w�����۾�2�2�s#��c'���!����� �8�پ�P����E����夾�c��.����� �2l$�J�'�Kk!���������Ծa������5Z�o
/�R�����(ν����i%���B���˲��$Ľ�(ཛX�Ԋ �T�F�"y�zX��Oy¾e��J �Kb�y�&�M�'�q<�7'�c��Z%Ͼ�&���͞��՝��b��?˾l��G��O��@'��'�l��������QƾҚ��+6~�n�J��#������fɽ�Ը�qk��c����½S�ٽ���U���46��/a��Q��>�����־�� �����D$��+�`�)��h�O��A!�7̾�������1�������m;�A��G�'���.��v+�pu��3�KM���ƾj!������%�X���5��6�-H
����'�｟r�ۗ�1��8�>!�c#;��i^��}�� >���Ⱦ���S*��!�.�9h2��-�oE�K�^��mξow���I���⼾C�־>����M���$��S1�k�4�ѡ.�=9 �K����w�ƾ����Xۈ��>g��G�$n1���!�P/��p��g�����a!���/���D�:Aa��ك�����ݼ��⾛���G��{,���6���7��-/��������Ͼ�j��	p����̾���j�����Iw-�d�6��7���-�G��r����ݿ�H[��ύ��H�c��F���1��S#��B�c$������8�&�{6�V1M���l��L������+�Ⱦ���/��}�!�D�0�'j8��66�7�*���H���k�b�ɾ����_¾v!׾����k]���#�_�2�=9���5�j�)�����w�op۾-���)}��߀�'^�8D�H�1�(%���4K�C��w�$���0�L�B�vN\����  �  cc�V���5����]ǾR 龌c����O���/�� ����	��A�����]#���Г��;��+�ǾA���lO��H�to�v���8p��=y��ǭ����]���8���h�����/jҽ��ŽX]ý��˽�߽�����L�H,��rM� 8w��T��v���(&վ
�����?���A�H
��v���Fؾ���`���b���7���2��>���DԾi������B�������	������5ؾ$���#Ǘ��"{�+�P�,�.�1��̟ �$*但�ѽn0ʽ#�ͽ{�۽������,0#�~@��Se����$2��3ž�羑i���^R��^��
�״�� 9վqp��7��!u���˚�霬�<ɾ��Y��@D��������m�K����ھ�ﹾ�����0��1a��9B�|[*��X�����;��2�z��?��%�2/�{�G��g��)���m��b{��hFݾ{���5X�*��?���B�����-����־�b������ᢾ�㫾Ϩ������i����F��i����Yg������ܾ����T-�����h4q��:U���?���/��=%������G�$�L�.��E>���R��m�;7���%���ݵ�86Ծ�����-�y���� �>@!�j�֢����5׾�-��T���:���Rκ���Ӿ+��g�
������ �)� ����r�2f����־���ڝ�P���uo��T�
@���0�>�&�8"�K�"�P�(��A4�)�D�>�Z�V�v��k��*磾MH���޾ib �76�#D���!����b��ʼ�ʼ��ξ�+�������p�þ��߾� ���������"��> ���^�j�ȅξ2�������鄾Țj��CR�ڬ?��M2��%*��Q'�)�)�:�1���>��Q�Di�����  �  ��n�%�����1���)˾�l߾s��Kc�B�l�վ�輾����mۋ��z�z}q��S���������YþPe۾���{��U����ܾf�Ǿ����p����jk���M�J�3�=z���
�����'��A�>���s�5O�td*���B���^��)��)���\��Y����Ծ[;�L��0�NH�8о=���@��U����:x���v�'ׅ�Wy���Ѳ�Q;`�⾛��C��v=��x־�2��7������iр�E)a�oE��,�ܪ�o�C������'^�>����Gx#�E�:���U�t��P������N��)�̾�Y��������%�������ϾS���,��⮋���������Օ��Z��PǾ� �m��������������$ݾ�gƾ�ʯ��F��	s��p,t�݂Y��`B���.�' �`������G]"�Um2��G�o8_�Բz���ڞ��W��U�ɾNᾝP���p�i1�	e���-��{ӾUc����>���㐐�kח�;2��o���5�ܾ������ �+A�M{��Ð��˾����K��O���l��n2m�2�W�yF�Q09�L62���1���7� D��oU���j�遾����$�������Ǿ��޾s)������ԗ�6��{��l�վ�𻾾\��6���.���s�����x{Ҿ����\�_����\#������i�bɾ
���%���ݐ�\����l��EW�qF�:��74��5�X<�C�I�(S\���r��-��	۔����t@��z<Ͼ�k����1�Ф	�*��p����e辺�;u������'���$ޞ������¾�6ݾ.���]�H�	�(��!������ھ1Zľ9ϯ�7띾Pq������ Ij�SJV�?�F�K�<��69�aY<�p�E�f4U�i�I�������  �  ����ِ��>��	������#���tþ��¾����9��u ��25���<h���Q�<XK�2�U��o����)��߶��NA��`�ľ�þv�������7����a���/������7sr���Y���@�Z*�T��i�������$"�S'7��O��h��q���M-������yv��𺹾��¾�]ƾ�Yþ5⸾�C��(f��:�O�b��FQ�AAP���_���}��ꑾt٥��궾a¾!�ž��¾�+��{��s*������s������_j���Q�ӹ9�a�$�������������.��OF�j`��z�~���{w�� ���ꬾdḾ%�þeD˾+;��Ǿ�]��z����Е�����08m���a�X�g��Z}�1̏�� �������Ǿ�Ѿ�Ҿ��;
~ľ����n���+���������f��f���O���<��U0�~3,�p*1���>�y�R�ik��}���%������������	⽾��ɾ��ӾT[پ��ؾOѾ�¾9�����5O��px���&{�;���|��������)�ʾoxؾ�2߾7�޾��׾ �;�$¾ ���e«��Ԡ��w��đ��Y{���e� �T��QK�
IJ��&R���a��lw����7˔�� ���������S,þ��ξھ�⾅|澒[�I�ؾ�Ⱦ�%��!�������B��`�������sr��o�����ž�־��_��I���Rھ"AϾ�zþ���pӬ��p���s��g���ȍy�N3d�r�T��L�P�M�%�W�� i��p��)��&�������`����@��Y�ƾٸҾZuݾ������9�ˈԾ-�¾�s����c����������������9���%����;�0ݾ��}��<���پ+�;����ڮ��\������i����j���:w�ˏc�$\V��zQ��U��Pb�2�u�磆��;��?����  �  �t��1ӣ��V��L2���@���z������	���u���ˈ�L�s��U���<�h,�\�'�5o/��^B�:F]��{���������.���楾������L���/���4���_��������χ��~q�iT�C
<�ve-�c�*��o4���H���d�⦁�� ��7~��z<��|���D��F�������eA��oۤ��1��I�������m���P���9���,�6#,�|�7�|qM��i�]��8���j������t[��^�������݋��������ћ��ڐ�����g��#L�5�7�:u-�t�/��>�1=W�J�u��Ɗ���ţ�����JX���ӯ��:��"᯾�+��t���>@��Mߖ�2ň�o�s��.Y��.F�M>�=�B���R� jl�������������������3���M϶�r���'j��hP��s���!%���,�������{�-3b���P�.�J�l)Q��2c��}��l�����Ψ����B}��������&��BT��p๾6�������J�����2ၾ@k���[��W��7`���s�݇�F����������Ӵ��r����þ�þ#�þ=þ�[��A����G��D�������ه�2�x�k�~;i���s�-k����@��������^�þ�Ⱦ.�ɾ�4ʾ��ɾ�Ⱦ{�ľ6��;����奾����
��]&y��(l��^k�:�v��\��&����գ��ı�������þ�nǾ\�Ⱦ�>ɾ��Ⱦ[Ǿ�~þ�;���3���)��'퓾	؅��`v�c�k�o�l��z�*���'���~ݦ�nr�����0Ež��Ⱦ)�ɾiʾ-�ɾ��Ǿc�þ���������C�������&v��Mm�.�p�b7������{�������·�Hs���dǾ=Lʾ{Z˾s�˾��ʾ��Ⱦ��þy��W��<���Q����z����v��p�P�u�����u������G����.���  �  )�¾f�¾��x���s��Yԛ�����Lo��Ԣs�x$[�GB�	#+�a�tt�	��������0���H� b�7�z��򈾬8��w����}��, ��|g���Jž�þY������j#���m���:f�v?R�Z�N���[�V�w�с��Ȫ��,�������n#ƾtľNx�������󥾂g���1��`܃��o�1�V�A>��(��2�����5�����%�E";�ʌS�ebl���6_��F{��E磾��������i�¾�dž�%��B����U��*}��'�{�&_�ZQ��T��g�/K��ꎘ�R��-��^�ȾO�˾Ⱦm`���A��=���Z���Q��f	��\v�X�]�!�F�2�2�P
%�:}��#��2/�`tB��[Z��4t��ᆾ?���ك�������ĵ�&�����˾K�ҾEYӾ¼̾&���¬�����6x��Q�v�E=n�?�v��s���O��%έ��>��� о5ؾ��ؾ��Ҿ��Ⱦ�B��=���dz���f��-䃾]so���X���F���;��.9�U�?�yN�P�c��j|�8/���×�R���w��α��ڠƾI@Ҿ��۾����߾T�־D�Ǿه��F_�����d��G���񣍾0؛�cʮ�{þ>!վ�����;��ݾ=,ҾQƾ����T��{⣾����1R��q�}���g� �V�~M�sL���T� �d��z�Ȃ������\���|\��$����ľX�ϾN�ھ�
��徱�ᾤ־~�ľ٥��	����-���������>��mء��s���Fɾ��پR�㾏w�DX�qپ�.ξIv¾���j���̇��'x�������w�.uc��U���N�3OQ��\��o�������[	���ާ��5��V���Hʾ־�l������ᾜLӾj���쨬��ݚ�*����܉�:����v��R�����'Ҿ����  �  ���t쾎8޾��ɾ�沾F���2j����m�0�O��@5�9���
� l�����Ὄ꽓;��Ͷ��6$��G<�b�W�@w�(͍���w��-Lоӳ㾰��4B��<��hӾ/ع�0���a����y���t�!������*Q����Ⱦ9�߾���:�����xھx�ľ٬��A◾ ���	�g�3�J�<^1��V��C	��d���K꽔i�s����3����.�z�F�dc�`��h픾d���`���[׾̞�V�����Uι˾�簾��������Aw�,�z�<#������^��վ̅�"w������GH���پt{þ;���>՗������k���P���8���$�;�S��4��
�!����"���6�ByN�Xsi����ć���������l-׾%-쾬���9 ��V��[��{�Ѿ�Z�����g���\ ��H���e^���㶾S�Ѿ�뾳p����:� ����g�߾��Ⱦ�V��H��jꌾ��{�[�a�nkK�c�8���*��"�	!��&&�{�1���B���W�N�p�1g���b��'�������c�Ծ�����Y����d���Y��X׾̽����5����~�������j�ξb�G �'���	�|������>徕ξ8$��\����tR���	q�A�Z�Q�H�R�;�fj4���3��(:���F�X�ؕm�UN��������7	��|�ʾ������t���������� ���?.Ѿ���nФ����QQ�������y���o׾�n��)�� ��+M����Bnݾ��ƾj���1E��{i��Ę��Sk��\V���E��;�eR6��S8��@��@O�ugb�Wy��ԉ��ܘ�0��`&��>zԾ��뾜Q �����k
�nP�`������	˾�k��g���뜾e ��7x���ȾB4�}�����  �  #����ی�羜�že��8�����a�{�;�R���S�e>��6н����[Ž�
�Ľ�ֽ\��c*��#%��E��`m�g����U���}ξ���6�,`��M��d������Qݾc������{���錾�ؗ������ξCY���r��A��4x�	[���޾�ڼ��k���a��vX� 5��\����bl罜|ѽ$ƽ[XŽ!JϽ��㽣K��[�0��S� )~�||��xj����پ�)����	�h���
�>��JE��ѾD���	�����#������.��;�ܾ������������
���V�پ����Y���F��y�Y�B�9�(� ����Kg �;X𽝞�s��p������x�6���T�M�z�(ߔ��-��%�Ѿ=N��	�n:�����w�������:־,H���룾u���#�������Ծ����_����=�����^����T۾~纾!e��Tˆ�.�g��OJ�Ō3��"�.���M�t<����$1�&,�`�?��Y��5z��}�����mjȾ��龧������4�uO�i��n�����0FھYe��b:�������˷�GϾ��q���f@ � �!�����u���e:ݾ����󆢾qC����t��	Y��^C�#3��(��O"���!���&��21�L�@�^�U�1�p�v�����u���إؾ�F���L��'��!��V ����I�	��8�=Ҿ��%����;�������پ���E��g��ky!��z �e�0M
����cҾ�R��"���p���Yl���R�m?��-1�!(�e$�g&�"�,�L79��J���a�e�C2�����a�ž}�循��F�xp�1�"���7���m���˾@��*M��ꩵ��'ɾ�~�&����\3��  �  &'��]"�A���Ӛپ���������_�՘2�����3�BPͽ������_���-���>���}�ս����R=���m�������΁�jT��q�o)%���'�e� �k������=�Ծ�����)���w���r��ž���ʰ	�H��8&���'� ��f�j�����;|p��Pτ���S�)y*����&�,̽﷽{Э�z'���뵽t�Ƚ��5D�\�%��M�,ှ����ڑȾy��9��]$�j'��l&�Vt��|�����Ⱦ�諾̕���񟾊�����Ҿ�9�����l�!�O`*��)�3�������ƾ�&��恾�R���-�̾��u��B�"Z׽��ҽmL׽)�����1����)�"SK���w������绾��T��{!��Y)��H/���+����6��
��%;�Ҵ��߫�����=:˾����?��M�,���1�r-����`���Y��xƾ�Ѣ��օ���^��m=��X%������	�;��G� 6����t����1�zM�F�r������z��]�վ=���K��H''���2��5��#/�Dg �o!�k����Ҿiw���*��wɾ_���R��D�+�T�6�9C8��X0�� ��~��Y�ƾ���T퉾�Uj�avK�x5��m%��K�/�T���:���#�]o2���G��ce�ٴ��=栾��� �辏�	����i.�zR7���6�;�,�Q��՘����i�˾gC���.��?hѾ��@K��+ ���/�F8�r6�ү+��-��R���ྶ�<���Xꂾk`���D�gB1���#�f��UZ�.�� ��U+�>]<�1hT�Xju��^=��gfо������OW%���3��u9��5�!�(��|�8�r��-�Ǿ����4Lƾ�zݾ�B ������'�>5��  �  #-7�o�1��Z"���t��5,��)�����a�e�/���
�����E������?��# ��dʝ��׬��ƽ
��Kf��5;��p�)!��hžu������K'��4���7�
0��q	���l�����^妾�V���'Ծ�9��J��&�)���5�-�7���.������^5۾93��D����S�#D&��>��Eܽr��i���� ��ƀ���˱��q ׽[��j-!��M������ᨾ�&վY���	�Y�,�z�6��D6��+�n��vV�fؾ1 ��� ������Hb��fM㾫�x����0�7U:�Ľ8��,����N� ��Ҿ�K��%����Q���(�R��Rk�H׽^VɽHŽf�ɽ.7׽_�S�	���#���G��>y�cӜ��ľ�$����2(�Ty8�IM?��;��,��-�����[۾�7���4���ι�پP: �7�|�,�!<���A��\<��%-�"v�S�����Ͼ�x��҆���[��7�<������d������G ����'��%�*��H�<sp�L��j��྆��6 �x 5�y�B���E��H>�1�-�w�������߾�`ʾ�ƾ�eվZs���X��)&���9��UF�71H��?��+-� �f����vξ3@��󉾬!f���D�z�-����*��W����"�*���*�0A���`�p���ģ�nɾ�f������E*�x�<��.G���F��Z;�I8(�8���a��&ؾR�Ǿ��ɾq-޾,� ����$-���>���G�}F���9�Ŀ%�����뾴���������~>[���=�Ž)�}j�Z������������#��5�?N���q�g���l��hMپR�����f2�˫B��xI�&3E��6�  "��j�����eӾ�ɾ�Ѿ�N��3	����<5���D��  �  
ꕿ�Ő������f^�o,4�����a׾�����9z�"KC��\���Pv轲l׽�ӽ˲ڽWｅ�	��%��OO�G{��ܮ���k��1>��dh��ᆿ;���$���֎���~�4W�w(0�K��#������D��!�xE��m��ሿ@@�����l����z�֋Q���'��'�;�ƾ\�����i��9�t��X���S��=۽�gڽ��彏�����<�3���b�j���Y�������"�DGL��u��Ƌ�o3��Ԡ���9��#�q�A`I��F$��������0�����-�(T��Z|�ۜ��h2������\T��H~p���F��������64�������e�Dt;�u�#��1�������������!5�g�Z�8"������a2�@��n7��a�����;������������9l�S=D���!���
�[2��W	�J��	A��%i��ㇿ�����:���%���#���Di�?����+:�j���_6����o�;�J�C2�}#�ab�6"����}5*�E&=�^Z��(��(F��c�ɾp� �UX#�B�K��v�r���])���/���������0Nf���?�K� �]?��
��:�R|1�U�U�P^~�A'������=��#ѕ��x���a��8��i��&��η�y���y�N�W�_A�,�3�8-�n�,��t2�Q�>�b�S�g�s�PO������S�/!��3�ޘ\�� �������q��㜿~��j����Y���4��8��w��=�Q�n<��b��p��8���J��Q���쐿�}���S���*�W�/־�[��ˁ��J�m�5�P�K>�xK3��/���0���8��.H��`�������^¾���r����A���k��܉�����F�����p獿2+v�N�S�+��R���ج��x(�/J�+�q��2��(6���  �  _����؋���|���W�n/���	��8Ծ<|����z���E��j ��f����ݽٽ���������(�cGQ�~����a���H�sb��9��Ia�Ws��6��@������tv�0�P��M+�E�#�����%��m����?�cf��X��q0���Ր��Ԉ��r� �K��#�qW���bľ���Q9k���;������ï�h]὘�པ콌��<G�G�6��
d�6����\?�����dxF�f�m�X��������o�����i�zC�������������/%��h(�f�M�UYt��މ�K��l���;х�i.i��5A��=����'���ő���g��S>�W"��h�pS����������-��78�8�\�R���7����JݾU����2�O1[�K���Î�)Ô�c�������'e���>���D������X�7t���;�8Kb������������:���ヿ�b�zR:���(��n������q4r���M��\5��:&�=w�)��"��p-�vf@���\��!��iP��B_Ⱦdh��8�� �F���n�RO���#������5��������_�*�:�����V�a1�"���;-�z:P�M�v�X����u��������N���f�[��3����O���B������F�{�E�Z���D���6��G0�&�/���5�K=B�_W�hv�*
���=��C.޾����/���V��E~�:S���R���ʗ��፿M�z���S��P0�q�����jd
����g�7�X�\�hm���萿�蘿�A���h���=v��5N��6'�T�MZԾ�E��ni����p��T�ncA�Rm6�02��3�� <�IzK�äc�Ã�늝�Rz��o��3��b=��je�F�������nݙ���x����o�޳H�+�'�A�u�����ϟ$���D��k��釿?H���  �  ������|�4�e���E�͹"�d���{̾i�����~�W�M�ڔ*�.��O�����(��g���*�����2��X������Z����ؾ��	�'+��N�r�l�]���$낿;�y���_�"�>�4���$�%j�9x��>�������/���Q���o��^���ӂ�L�w�c]�AB;�b��\��8Ӿ�┖���p���D�1;%�zY�[K�<v��d��
��������!���?�j/j��#��i���\�'c�9�6�o�X��t�;$�������q���T�, 3�C������x����E`��d��k<��S^���y�Z���˂�Xs��\U���2�j��$�澆趾7l����n��H���,�%��n��h�OR���c�)�qB��^e������P���H־�`�ݾ&�׷I��j�=�������3b��Rq�ХQ���/�I�����&�ﾁ���)���w-�r\O�ƻo�����?����׃��p���P�>�-���lY�����q��\lz���W�%�?��U0�l(�"�&�,�+��7��J�(�f�-؆�W����Sžx��&!�L�8��[���z��x���򉿡��(�n�`�M�F*-����#��] ���
�[!�oU@�]\b��0���������T/��}m���K�y�(���	��4߾ ն�y���kg��(e�VO���@�k�9��Z9���?���L��{a� �����!B���Jپ�����$�j G�sNi������`��㉿�@��tre�l�C�L$����� ��[�i��ç*�2KK���l�\胿.኿|��q#���jb�L�?�H���@ �@�о���-򐾟�z�?�^�q�K�b6@�͖;� �=��1F�G�U�0�m�����Ɵ�d����y����0���S���t�â���ȋ��v���{�-�[���9�u� ���2�B6�4���m6�� X��Lx�Cχ��  �  f^�MX��QF��X-������T�ľ"t������`���>���%����ʞ	���������]�+�`�F�H1j�Y�������Ͼ/ ��>��D	4�E�K�5�[��^��U�5/@��S%�>Q
�����Tξ/hɾ��ھ����9*���4��!M�Tp\�_�͌T���?�2�%��i
�a��m��ږ�����|X��|9���"��4�A*�'�
�ڱ�t. �;�5�BpS�[�y��ɕ�?�����ݾ�X�!�iy<��R�@�]���\���N�pL7����r�"�ݾRfʾ�c;2�4��I�#�\?���U�oSa���_��Q�h�:�ϕ�e�	�۾�V���>��d��\���@��-�O�!�+/�[ �5+��3=���V�L�w��u���鬾��ϾZ�����<2�o�K�q�^�"|f���`�-kO��	6�Ԕ�����侙�ؾ���0����4���N�-�a��i���b��2Q��A8����Y���ھ�j��⿛�G_���	l��S�b�B�|19�N7�� =�`7J�D�^�*�z�i���*Ц���ľ�,꾿��r&�2�A���Y�j`i���l��\c���N��M4�+��Z������N���$�h�)��XE�v�]���l�ғo��	e�%;P�r�5�������ھ�ֹ�`������]y��nb�8�R���J��:J�GQ���_���u�H��������浾��վZ��F��=2��L�_|b�Zn��Cm�D_�-�G�J2,��X������p���쾄�������2���M���c�^�n�{m�i�^�p�G��,���k���%Ͼs찾�f��)8����r���^�ǶQ��cL�&�N��hX�֛i�����`����������h�0���.!��}<�V���h�иp��+k�b�Y�@��n$�PN�?�������~��</
�Y�!�V==�"UW�1j��  �  �5�l�1�:�%�����r⾒�þ_!���+���$���Ba���E�	{0� �#������%�5��L�Ui�\߅���������o˾A(�_z�c��P�)��4��5���-����J	����x�ƾ���~A��a����Xؾ�v��'��J�'�us3��96�x�/�B�!�4������ھ�������t�����z�#M[��uA���.�	�$� �#�$�,���>�ǆW�W@v�R���2���2r���վ5������{�b�-��W5�y�3�N�(��������۾E�� D�������-ž��澳B�w�L�.��8���7��.�%d��?������~־�@��h@�� �����~���a��;K��;<�,N6��	:��,G�"�\�D�x��+���b���b���о|?x����R,�Ԗ8�D=�u8���*�*��8��p"�)�ƾ�����ž6@޾�~�1��&�*���9���?�-^<��0�� �ܞ��O��U�پ;��bI��Fy��+>���zs�%_�PS�rPP��@W��Rg��3�z���w8���K��me˾�}�A'�{��{'�@�7���A�b�C���;�9,�1����H��:�ѾrBξ�ܾ=����#�Ah%��8�(�C�+�F�|&@�6R2��� �|/������yݾ��ľ�Ư��k��3��������]n��.d��c��zl�]4~�֞�����F������d�پ����������/��?>���E��D�] 9�D$'�j�aO��xK޾ϾѾ"��]a���*�+��<���E�!*E��;�*n,�k;�{=�&\�>
վ`罾��������
ԉ��,|�_Yl�ӊe�~]h�`�t�3����8��혢��z��f8˾Z��jg�X���5%�_6�N�B��G���B�l5���!��d����fھԉо�Wؾ�X�7Y
��y�Om3�p�A��  �  �(��|�
��g�pk�D��Y о�̿�7����(���	��It���X�aOG��IB�B�J���^��E|�G����衾�����mľ6�Ծt�徲���(����+I�qQ�GP	�$<���۾�k��~h��:��
e���`��&���yWξ���߮�s=��������X	��� �y��GIݾ��̾}���?��� ���!��V�m��?U�QG���F��R��Zj��鄾����
ƨ�@��6Zʾ�ھ���N��������g�fg����'-ѾK&���O���u��?q������漾��۾�Z����
�	�����{�#�	��� �Uﾱf޾CξAܽ�������du��ѝu�e8a���X�$d]�j�n��<��vs�����%r����̾�Yݾ)������B	� ��v��q�������i-���a־�O���Ө�����G��cr���վ� ��~�	�"����������Y��'����?����վOž�}��p����������v��r��{�d������y��;)���>ξ�B߾���pn �ܐ	����ʨ���<Q�Y��q��ɍ��ϱ۾�Eþ?���=��ޗ���Ҿ�ﾚ:��+�c��Ip"�!M �k�����Ư�����=��ܾ�^˾)%��s��qؖ�bq���������N:��R����ä�՝����Ⱦ`ھ>������ �U�F=�����!�D����4g�>��{Ծ5U����� ���|�¾��ھU ��,����SK ��!��7�������/���<�����x׾,�žbʳ�DF���B��z���[����兾�$�������U��ތ��\�оf��C�Z�C
�L��Y��!�v�"���6�E����ּξf컾ش�����yp̾�:��(����a;��  �  ��#�'��/��$�����զ澀Pپ�gƾ��������u���m��jy��Ɗ��ើ}���ͺ˾��ݾ��)?𾑯�:?�9��H�O��uD���׾&9ľv�������;���u9u�,q����K��WУ�S����9оx<�sS���y��>��g��s��w{����վM:���^������2����s�]�r������A��a���l\���!Ӿ������l �A�f��1���O��LwѾ�����إ����g��^zs���v�3��%��^����CƾH1۾���|�������l��.���?w�����y��֨��־Ia��7᪾mƖ��h��6��H���/���	���Ϻ��Ѿ���P<������o' �� �X� ��{ �������������پ=ľθ��;W���.���z��,��K�����Mž��۾��V������p�,�����
��������zq��ܾ��ƾ+�������.�����`*��䨣�*2��{{Ͼ+�徐"���D�����5�^>� ���%����N��P%��˾����i4���ә�jD��Mܟ��k���sľ��۾�&�s�$���n	��]
��
�%]
���	�Tl�?��6���+=�!LʾI����f���ř�Q3���š�����bǾ/D޾��ڒ�����	�$�	�3�	���	�����o��@�i-�,%ݾ$Dƾ�$��t9��K"��T7��hL�����0�˾x}������������	�F:
��S
��(
�?(	�/E�� �;�ﾥuھʥþE2��Hu��;ޙ�V���{���m����о�r���������w
�2�
�<���
���	�3B�j �� ؾ�v������u?���+��#a��i0��L���*־H��7U���  �  �1��^�о�Y��^�K����-�V0��.
��x��y�߾����9���堕�ɫ��똘�"��e Ⱦ�A����w�n2�' ��!
�Š�c���6߾��ξ�y���w�������t��p�q�#�W� /H�SE�ҡO��e�� ���ԓ�}��a����>ȾŒؾ۵�r�����i�;�����������EC׾�@�������7���t���`�����/~Ӿq�}�e�7��	��o�����x�꾂`پ5ɾ����E��(?��^���˸h��}R�y�G��wJ�PZ�I�t��[������ܰ���¾BxӾ"K侴���]��!���@j�<�����8�� վ4򸾱Ĥ�)�����S���Oʾ�|�k�I��,�l��u����э���R�}.Ҿ����}"��|8��J���u~���k��ie�Gl�1���L��#ܟ�v���ѻľA�վ�c�@H��ɨ�l�����#�'0��@���	�B_��\�׾w罾B9��a���P�	�ľ�(�Tj �u���ς�*m�����0��������U�Ydھ��ɾ�U��զ�\▾�h���$��q0�������������񑴾��ƾ%�ؾ�1�F}���F�-a�Aa�u���"�z �$���h/���پ.[������:��'���վ�T�N+	�Pz����!�F��_��������c���龟Eپ�Ǿ𺵾����S[������ ���䃾�������w���-���P̾�ݾ]��|��{	��M���W] �\:"��=�mp�Zl�N��ySѾμ�I���K���9Ǿ%������A��f��2�!��`"�V����w�����������H־@jľB�����%���]��X��{^��P��������ڰ��#þվ�  �  Q��"žF�=��� ���&�}$2��C5�C�.��������lʾ����b���	��pѾIG�����s2$��}1�H�5���0�W$�q��Zc ��v޾���������6���4�B�^�mCD�^a0�7�$��"��i*���:��S��q�3#��U���ĵ��pѾ��V�(:�[w,�{W5�E5�`�+����(�����ґ¾����j��� ����a޾�>�A���)�(a4��x5��p-�o��3������~�Ӿɥ���������A�s�r�U�b�=�.-���%��'�H�3�t/H�U�c��p��w��2+���Uľ��ᾤ�C��)&�̶3���9���6��x*�!��3��CH߾�þ����/���7�Ҿ����B���$���4��W<�}r:���/����B�����jGؾ|ɽ�r_��s���g���j��,U���G��*C��tH��W��m�Hb��=���)��P���4۾���D���!��1�=�"E@���9��+�:2�WY�^W�j�ʾ�Aľ'BϾy��!�P���1��>��#C��.>�I1�-Q ���������Sܾf�þ�{��X���Ì�O��m$m���b��a��	j��C{��􉾰6�����9��+�־7U�]	�fk���-�k�<�]�E�j`E���;�U�*�����F��`�8aо�[Ͼ|t߾�,��&)��2(�
�9�hD��E���=�_�.�H��}�
�lp���Kؾ�~������?��^���@N}��	l�b�c���d�yno��S���s���a��Ұ��ƾz�޾������o!�=3���@��F�JfC��7�rE$��������۾�lϾzVԾB���?�'��/�_P?�T�F��D�,W:��1*�Y��W����R^Ҿ׻��^���q��p ��@�{���m��[h���l�'�z�(��MN�����m���  �  2���#�ƾeQ���%�.���G���X�"�^���V��C�I)�������Ͼ�`Ǿ�վ$����O�/���H��#Z�_�\�V��AC���)�R[��e�%ڿ�"���9��y�\���<���$�Y`�@�-�	��������1��HN�;bs����b���7׾B5�U����8���O�Pq]�Y�^�=�R�"L<�/� �Pr�Dg�^S̾�
˾��߾o�����89��MP���]���]�JYQ��@;�d| ����۾�[��`ᓾ��v�CQ�}4�ݪ��V�Х�ܦ��Q�z�)�%B��fb�J���s���bI¾�K�L��[*���D���X���b��_�N�O��m7�_��? ��n��Ҿdپ�Z��\G���,�ۤG�PF\�6�e��a���Q���9��g��E��<۾�q��ꐙ��6��%d��^J��#8�bY-��"*��.�Om:���M��Uh�*���~曾�x��\�ܾ)��]���9�r�R�Y�c� �i�<�a��N���4�`��l��{�m*߾� �q���n �S<��U�O%g�Y2l��c���P�77����5��Xf۾�����D�����31w�j``���P���H��9H��O�C]���r� ����s��ր���EѾ���̜��?.��#I�'�_���m�_�n���b�)KL���0�_��������~��P����-�G)I��G`��m���m��ya�oK�Y�0�/�� ���9�Ӿp���ܛ�׈�]�t�P_���P�0YJ�pFK�9�S���c��z��
��ZF���X��5�ܾ3�U�'=7�ZaQ���e�v�o�Il�#h\��C�_/(��#�un��؁����G4����~�7�/�R�b g��Cp�|+l��\���C�ͺ(����@�ﾛ˾	��������M�q���^�FNS�0AO���R���]�=p�]	��\�� ���  �  �3��m�ξ���L�$���G���g���}�Ă��|��2d���C�rQ"��C�ǯ�]J޾4�����X�)���K�\�j�6��邿!�z���a���@�����d����ž����[5x���I�^�(��]�j=��l��o���'��s+
����p:�b�b�k��ei�����\d�}1�RT��q����������v��[�]f9�J�������0b⾑X��ٮ��z5�WAW�+�s����`��5�s��SW�W�4���辒W������u�f��=�Bv ������ ����������zK���-�_O�zs}�f읾�9Ǿ*������@�;b��|�r΄�	񂿠]r�T��O2���������龄���	�y%�ezF���g�대�8J����� 9r�|(S�J0����a���������P�t�P��s6�!�%�y�^i�[[��(��9��6T�?y��ڕ�����;�����<�/��R��r��z��:F��M����eo�F%O�i�-���� ����2^���X6�N1X�;�w��}���w�������o��N��K+�	X��P�撷��K��k�����b���L��>�/�7��>7��V=�.J��j^���{����*��FӾ���-����A�cd�|ဿщ�j����M�� k��ZI���(�Z�����b���A�%��cE�>1g�xみ����"��4����g��+E�Y�"�<U���־�}���ٓ�~�3``�L�OI?�9��O:�+�A�xGP��f��t����ǫ��H��z�[�*�gjM��o����<$���;����~��z`�j�>� �a\
��� ���H3�d0�D�Q�o�r�dl����ƈ�Ι|��]��:�pC��)��^V˾�q��橎�qx�Z�]�DL�.�A�tz>���A��ZK��j\���u�Q��c���  �  0b��׾����1���Y�b�~�{u���ې�}u��i}{���V�ԃ0�����p��A��� ��2���8�Zk_�F���ǯ������遊�_�w�^�Q�i�)����Hi̾�圾ps�A��=�v���g�=��޽���m����E���0�+�[�(y��W��h�����@@�o5h�"&��	���
���G2��e�p���J�`�%�Z�	�w���)���""�KF�i�l�E������r��烆�?l�cQD�B��Y��u��Ə�ݘ`�T=4���X��9��F��轌i�����>�#��|F�[+x�%���(;|���(��$Q��x�+K���ڒ�غ��X����nh���A�,���S�ZO����U�� �2�ɡX��i~�nʍ�^\���$������f���=����n�}�����m�F�U�+�n[��`��������9w/�T%J�?q�����0����ܪ���<���d��턿�X^������X����a�L�;��t�o�����P#�P&E�^�k�R߇�� ��l�����������8_�
 7��o����,����䕾IVz�nX��B�H}4���-���-��n3��?�W�S���q�ѥ���F���0׾�+��k)���P�Fx��B���������G7��/i���Z���5��y���	����C���2�V�́|�M��������P����.|�o�T���,�L
��w۾�A�������t���U���A��k5���/���0���7�Z�E��O\���}�mF��U���~�ǣ���5�&�]�i�����W,��� ��������t�
.N��+�dO�
�����6{��!>� �c�ڳ���.��ʩ���`��79���rp�c3H�-�!�
�vξ�	��ӊ�x"n�MYS�ZB��D8�v�4���7�!3A�m�Q���k������L���  �  ,����Qھs��t6���`�����h��B���\��j���)L]���5����b���=��5��<��P>�Ĕf���1���l$��pX�����qX��.����k,Ͼ���|r���>�,�Д����V۽��ؽ�@�V&�����-�%.Z�����$��'��A���E�_�o�W�������.ϕ��錿�x�ʼP��*���ʊ������u
�I�&�8L��Pt�G���)��;��(&����s�pJ��� �5����������_���1�2��f������>C߽��⽱�̲�� ���C��w��>����Ͼ0��5-�wHW�Q��u�����AǕ�L����o��G�8�#�ނ
�����}�������7�)3_��Z�����ʅ���#��Pk���m�
�B�������޺�+v���k�� C���(�r��F����ף�1���/,�p G���n�1ߓ��]��AB�u��^tA�[�k��:�� 斿�����蕿����3�h��A��= ��f�`s�$+�6W'��J�B
s��F��&����������Ȇ�בe���;��+��꾚���j����w�fIU�v�>�CB1���*��*�C0�=x<�ϋP�w�n��ƍ�\m��,�ؾ�A	��-��V�����Б�����۝��r`����`�m:�������{���V�J}6��\�����B���*���&��R4���灿�;Z�v�0�gL��~ݾx����᏾��q�8�R��Y>�D2���,�>�-���4�3�B��$Y�	g{�>���2���� ��4��:��d�-m��<l���R������<���|��S���/�~�)E�l��`&#��C��ij��ڈ�R���Ӟ�K`��ǜ��@rw�nBM��%����|sϾ�릾�͉��*k�RP��>�{(5���1���4�h�=�E�N�Ͽh�=懾a���  �  0b��׾����1���Y�b�~�{u���ې�}u��i}{���V�ԃ0�����p��A��� ��2���8�Zk_�F���ǯ������遊�_�w�^�Q�i�)����Hi̾�圾ps�A��=�v���g�=��޽���m����E���0�+�[�(y��W��h�����@@�o5h�"&��	������G2��e�p���J�a�%�[�	�y���)���""�NF�l�l�G������w��탆�Nl�rQD�P��q����Ə�ɘ`�=4�w��~��7�3D�i���d�������#��xF�)&x�)����$;����(��"Q��
x�-J���ْ���������mh��A����`S�5O�������޺2�ϢX�&k~�7ˍ�D]���%������f���=�Ն�"r�Հ��ʕ���m��F��+�I]��a����"��Y���t/��!J��q�����-���������<���d��섿��f]����HX��s�a�v�;�ct��n�"��R�{Q#�2'E���k�����!��g����������.;_�*"7��q����|����畾J[z�=rX�wB� �4�8�-���-�p3��?�#�S��q�����F���0׾�+��k)���P�Gx��B���������G7��/i���Z���5��y���	����C���2�V�́|�M��������P����.|�o�T���,�L
��w۾�A�������t���U���A��k5���/���0���7�Z�E��O\���}�mF��U���~�ǣ���5�&�]�i�����W,��� ��������t�
.N��+�dO�
�����6{��!>� �c�ڳ���.��ʩ���`��79���rp�c3H�-�!�
�vξ�	��ӊ�x"n�MYS�ZB��D8�v�4���7�!3A�m�Q���k������L���  �  �3��m�ξ���L�$���G���g���}�Ă��|��2d���C�rQ"��C�ǯ�]J޾4�����X�)���K�\�j�6��邿!�z���a���@�����d����ž����[5x���I�^�(��]�j=��l��o���'��s+
����p:�b�b�k��ei�����\d�}1�RT��q����������v��[�]f9�K�������4b⾗X��ݮ��z5�_AW�6�s����j��M�s��SW�t�4����農W������O�f���=�iu ������ �\��t���P���E�p�-�|VO�ei}��松q3Ǿ���F��,�@�7b�B�|��̄�u�Zr��T�%N2��������q��C���	��%�X|F��g�i����K��􍃿�<r�z,S�N0�I��;��6ƶ����<�t�4P��x6���%�Y��i��Y�3(���9��/T�zy�KՕ�p���T��5��=�/���R��{r��x��mD�������bo�!#O���-� ��l �����^���6��3X�	�w�W��by�������o�N��O+��[��W�R����Q��H����b�S�L���>���7�fB7��Y=�0J�Bl^��{�^��p�$GӾ���4����A�cd�|ဿщ�j����M�� k��ZI���(�Z�����b���B�%��cE�?1g�xみ����"��4����g��+E�Y�"�<U���־�}���ٓ�~�3``�L�OI?�9��O:�+�A�xGP��f��t����ǫ��H��z�[�*�gjM��o����<$���;����~��z`�j�>� �a\
��� ���H3�d0�D�Q�o�r�dl����ƈ�Ι|��]��:�pC��)��^V˾�q��橎�qx�Z�]�DL�.�A�tz>���A��ZK��j\���u�Q��c���  �  2���#�ƾeQ���%�.���G���X�"�^���V��C�I)�������Ͼ�`Ǿ�վ$����O�/���H��#Z�_�\�V��AC���)�R[��e�%ڿ�"���9��y�\���<���$�Z`�@�.�	��������1��HN�;bs����b���7׾B5�U����8���O�Pq]�Y�^�=�R�#L<�0� �Rr�Gg�cS̾�
˾¹߾t�����89�NP��]���]�jYQ��@;��| ����۾�[��pᓾs�v��Q��{4����8T���͡�UK�8y)��B��Zb����5���+@¾�A���$V*�H�D���X���b���_���O�{j7�������l⾺�Ҿeپ=]��QI�p�,�I�G�oJ\��e�L�a��Q���9�m�'K��F۾Uz������5=��X/d��fJ��(8�\-��"*���.��h:�e�M��Kh�懅��ޛ��o����ܾՠ����U�9�řR���c��i���a�.�N���4��]��k� z羅*߾�"�����p �*V<�^�U��)g��7l���c�^�P�7�������{p۾Ϟ���L���
���<w� j`���P���H��>H�TO��E]���r�龇�It��6���
FѾ��֜��?.�$I�'�_���m�`�n���b�*KL���0�_��������~��P����-�G)I��G`��m���m��ya�oK�Y�0�/�� ���9�Ӿp���ܛ�׈�]�t�P_���P�0YJ�pFK�9�S���c��z��
��ZF���X��5�ܾ3�U�'=7�ZaQ���e�v�o�Il�#h\��C�_/(��#�un��؁����G4����~�7�/�R�b g��Cp�|+l��\���C�ͺ(����@�ﾛ˾	��������M�q���^�FNS�0AO���R���]�=p�]	��\�� ���  �  Q��"žF�=��� ���&�}$2��C5�C�.��������lʾ����b���	��pѾIG�����s2$��}1�H�5���0�W$�q��Zc ��v޾���������6���4�B�^�mCD�^a0�7�$��"��i*���:��S��q�3#��U���ĵ��pѾ��W�(:�\w,�{W5�E5�a�+����)�����֑¾ ���r���+����a޾�>�A���)�?a4��x5�q-����c��K�����Ӿ�������􃋾{�s���U��=��-�P�%���'�-�3�7%H���c�?i��4n�� !��\Jľ���%����"&�|�3���9�Y�6��t*����s��yD߾�þ����h���!�ҾZ���w�ҽ$���4�P]<��x:��0�����������gSؾLԽ��h��a���m����j�\3U���G��*C��qH�� W�Ѣm�\��r����������ھ����k���!�B�1�=�1?@���9�!+��.��V��S�ŞʾBľDϾ&꾰$����1���>��)C��5>�R�1�SX ���C���w`ܾ��þ󅮾�`���ʌ�`��7.m�g�b�#�a��j�^G{������7����\:��s�־aU��]	�kk���-�l�<�^�E�l`E���;�V�*�����F��`�9aо�[Ͼ}t߾�,��&)��2(�
�9�hD��E���=�_�.�H��}�
�lp���Kؾ�~������?��^���@N}��	l�b�c���d�yno��S���s���a��Ұ��ƾz�޾������o!�=3���@��F�JfC��7�rE$��������۾�lϾzVԾB���?�'��/�_P?�T�F��D�,W:��1*�Y��W����R^Ҿ׻��^���q��p ��@�{���m��[h���l�'�z�(��MN�����m���  �  �1��^�о�Y��^�K����-�V0��.
��x��y�߾����9���堕�ɫ��똘�"��e Ⱦ�A����w�n2�' ��!
�Š�c���6߾��ξ�y���w�������t��q�q�#�W� /H�SE�ҡO��e�� ���ԓ�}��a����>Ⱦƒؾ۵�r�����i�;�����������HC׾�@�������7��u���`�����C~Ӿ+q��}��X��2����������`پyɾ�����D���>������7�h�-zR�6�G��pJ�(Z���t��T�����Ұ���¾okӾK=�6��zV���y��c��{� ��k���Ծk¤���Z ��!W���Tʾ~����`N��2�3�������F��k'�_⾽:ҾF����+���?���O��#}~�]�k�je��Cl�m��}G��՟��y��.�ľ �վ�U澜9��*�����;
����)�;��	��W����׾�㽾{7�����W��ľ�.�On �m�����|t�t���8���ӧ���c�1qھ��ɾ�_��Xݦ�6閾jn��)���3��kÇ�������������ƾ��ؾ2�o}���F�2a�Ca�w���"�| �%���i/���پ.[������:��'���վ�T�N+	�Pz����!�F��_��������c���龟Eپ�Ǿ𺵾����S[������ ���䃾�������w���-���P̾�ݾ]��|��{	��M���W] �\:"��=�mp�Zl�N��ySѾμ�I���K���9Ǿ%������A��f��2�!��`"�V����w�����������H־@jľB�����%���]��X��{^��P��������ڰ��#þվ�  �  ��#�'��/��$�����զ澀Pپ�gƾ��������u���m��jy��Ɗ��ើ}���ͺ˾��ݾ��)?𾑯�:?�9��H�O��uD���׾&9ľv�������;���u9u�,q����K��WУ�S����9оx<�sS���y��>��h��t��x{����վO:���^������7���+�s�o�r�����B��v����\���!Ӿ��>�U��� �B�����1�>�p��1wѾ����ץ�����e���ts�&�v�d���
��Ю���:ƾ�&۾��꾔n��W����]������fh���w�����x��`�־sY��=۪�N�pf���5��sI��3������ֺ���Ѿ��徭H��^����. ��� �� �� ���������뾠�پ� ľ����$[���0���z��{��}G��`����ž5�۾T���I�����4i�F�����a{�������fﾌ�ܾ�ƾ����<���,�����j,��ᬣ�%8��y�Ͼ$��j.���K�R����-=��F����:-�g#��Z���/��#˾Т��B:��tؙ�H��ߟ��m��;uľɒ۾D'��H���n	��]
� �
�(]
���	�Vl�A��9���.=�#LʾJ����f���ř�R3���š�����bǾ/D޾��ڒ�����	�$�	�3�	���	�����o��@�i-�,%ݾ$Dƾ�$��t9��K"��T7��hL�����0�˾x}������������	�F:
��S
��(
�?(	�/E�� �;�ﾥuھʥþE2��Hu��;ޙ�V���{���m����о�r���������w
�2�
�<���
���	�3B�j �� ؾ�v������u?���+��#a��i0��L���*־H��7U���  �  �(��|�
��g�pk�D��Y о�̿�7����(���	��It���X�aOG��IB�B�J���^��E|�G����衾�����mľ6�Ծt�徲���(����+I�qQ�GP	�$<���۾�k��~h��:��
e���`��&���yWξ���߮�s=��������X	��� �y��HIݾ��̾ }���?��� ���!��^�m��?U�]G�ϬF�2�R��Zj� ꄾ���.ƨ�p��sZʾN�ھ��뾰�������+g�xg��p�`,Ѿ%���M���r���m�����༾V�۾�Q��=�
�����f�ѳ	�,� ��F�LY޾�6ξ�ѽ����������o���u�4a���X��f]�f�n�A��z�����<|��i�̾�fݾO+�� �J	�}��}�5x�f��q��5��ag־tS���ը�����E���n��h�վ(��͋	�������������SR� �q����得�վ�ž�t��H������=�����v�B�r���{��g����������2���Iξ`O߾"��v ���	�������F#��W�V�����������۾EKþɢ���@�������Ҿ�;�M,����hp"�2M �t�����ɯ�����=��ܾ�^˾+%��u��rؖ�cq���������N:��R����ä�՝����Ⱦaھ>������ �U�F=�����!�D����4g�>��{Ծ5U����� ���|�¾��ھU ��,����SK ��!��7�������/���<�����x׾,�žbʳ�DF���B��z���[����兾�$�������U��ތ��\�оf��C�Z�C
�L��Y��!�v�"���6�E����ּξf컾ش�����yp̾�:��(����a;��  �  �5�l�1�:�%�����r⾒�þ_!���+���$���Ba���E�	{0� �#������%�5��L�Ui�\߅���������o˾A(�_z�c��P�)��4��5���-����J	����x�ƾ���~A��a����Xؾ�v��'��J�'�us3��96�x�/�B�!�4������ھ�����u�����z�(M[�vA���.��$��#�8�,��>��W��@v�q���[���gr��U�վ����9���{���-��W5���3�H�(�Y�������۾����A��F���k)ž2��C?��r�m�.�-�7���7���.��]�.9������r־�5���6��|����~���a��4K�.8<�bM6��:�B2G��\���x��2��zk���l���оL�S�S��,�9�8��I=��z8��*������	&��ƾ;��� �ž�<޾|������*�ҫ9���?��W<��0�������B��9�پ]���?��eq���7��[qs��_�\	S��PP��CW�-Yg��=�����@���U���p˾R��	.����'�O�7�c�A���C�<�;�#,�7��:�����]�Ѿ�Eξ�ܾ���7$��h%�18�U�C�E�F��&@�=R2��� �/������yݾ��ľ�Ư��k��5��������]n��.d��c��zl�^4~�֞�����F������d�پ����������/��?>���E��D�] 9�D$'�j�aO��xK޾ϾѾ"��]a���*�+��<���E�!*E��;�*n,�k;�{=�&\�>
վ`罾��������
ԉ��,|�_Yl�ӊe�~]h�`�t�3����8��혢��z��f8˾Z��jg�X���5%�_6�N�B��G���B�l5���!��d����fھԉо�Wؾ�X�7Y
��y�Om3�p�A��  �  f^�MX��QF��X-������T�ľ"t������`���>���%����ʞ	���������]�+�`�F�H1j�Y�������Ͼ/ ��>��D	4�E�K�5�[��^��U�5/@��S%�>Q
�����Tξ/hɾ��ھ����9*���4��!M�Tp\�_�͌T���?�2�%��i
�a��m��ۖ�����X��|9��"��4�K*�3�
����. �X�5�hpS���y��ɕ�i���Ŀݾ+�z�!��y<��R�\�]���\���N�PL7��������ݾWdʾ�`;x.���j�#��X?��U��Na���_���Q��:�e��4�a۾�M��_7�������[��@���-�E�!��.�G] �n+��:=���V�x��|��G���Ͼ���~��MB2���K�ư^��f�a��nO��6������T�侼�ؾy���������4�
�N���a��i���b�8-Q��;8�a��cT���ھ(b��J����X����k�x�S�z�B�/9�4N7�9=��<J�-�^���z����ئ���ľ 7�G�^x&�!�A���Y�fi��m��ac���N��P4������P��D���%��)�)YE���]���l��o��	e�+;P�v�5������ھ�ֹ�d������]y��nb�:�R���J��:J�GQ���_���u�H��������浾��վZ��F��=2��L�_|b�Zn��Cm�D_�-�G�J2,��X������p���쾄�������2���M���c�^�n�{m�i�^�p�G��,���k���%Ͼs찾�f��)8����r���^�ǶQ��cL�&�N��hX�֛i�����`����������h�0���.!��}<�V���h�иp��+k�b�Y�@��n$�PN�?�������~��</
�Y�!�V==�"UW�1j��  �  ������|�4�e���E�͹"�d���{̾i�����~�W�M�ڔ*�.��O�����(��g���*�����2��X������Z����ؾ��	�'+��N�r�l�]���$낿;�y���_�"�>�4���$�%j�9x��>�������/���Q���o��^���ӂ�L�w�d]�AB;�b��\��8Ӿ�┖���p���D�4;%�~Y�`K�Iv��u��!��������!���?��/j��#������\�<c�Q�6���X�.�t�F$�����~�q�o�T��3������Zw�����^��b��i<�8Q^���y��	���ɂ�s��XU�̻2����V��fⶾ�f���n�sH�@�,�T��O�;h��S�	���)��wB��fe��Ɗ��V��uO־Rd���&�ջI��j�)���d����c��q���Q�P�/�b����?�ﾎ���(��'v-�XZO�!�o����v����Ճ�p�p���P�B�-�C���R�򀶾yl���cz���W���?�.R0��(�?�&��+���7���J���f��܆�䈡��Yž���%�p�8��[���z�{����O���n���M�C,-�����$��^ �n�
��[!��U@��\b��0���������W/��}m���K�{�(���	��4߾ն�{���mg��+e�WO���@�l�9��Z9���?���L��{a� �����!B���Jپ�����$�j G�sNi������`��㉿�@��tre�l�C�L$����� ��[�i��ç*�2KK���l�\胿.኿|��q#���jb�L�?�H���@ �@�о���-򐾟�z�?�^�q�K�b6@�͖;� �=��1F�G�U�0�m�����Ɵ�d����y����0���S���t�â���ȋ��v���{�-�[���9�u� ���2�B6�4���m6�� X��Lx�Cχ��  �  _����؋���|���W�n/���	��8Ծ<|����z���E��j ��f����ݽٽ���������(�cGQ�~����a���H�sb��9��Ia�Ws��6��@������tv�0�P��M+�E�#�����%��m����?�cf��X��q0���Ր��Ԉ��r� �K��#�qW���bľ���R9k���;������ȯ�o]ὡ�འ코��GG�U�6��
d�B����n?�����qxF�s�m�_����� ���o�����i��yC�b��B���������$��g(�Q�M�Xt��݉�j��w���9Ѕ�^,i��3A�<����������c�g��O>�,T"��f�YR�������h��J0�;8�v�\�獈�<��� Nݾ6����2�d3[�V���Ď�Ĕ�8���Á���(e���>�����������X��s���;�Jb�����������9���⃿ėb�hP:�����꾸k������/r�Y�M�EZ5�69&�ev�)��"��r-�Ki@���\��#��ES���bȾl��@��(�F���n�mP���$������6��b����_�4�:�� �aW��1�~���;-��:P�m�v�b����u��������O���h�[��3����Q���B������H�{�F�Z���D���6��G0�&�/���5�K=B�_W�hv�*
���=��C.޾����/���V��E~�:S���R���ʗ��፿M�z���S��P0�q�����jd
����g�7�X�\�hm���萿�蘿�A���h���=v��5N��6'�T�MZԾ�E��ni����p��T�ncA�Rm6�02��3�� <�IzK�äc�Ã�늝�Rz��o��3��b=��je�F�������nݙ���x����o�޳H�+�'�A�u�����ϟ$���D��k��釿?H���  �  ��꿕�ῘUɿ�̧������J�M�r%������4��LR���/��N�e��^�����7��R�6�I#]��G���K���<���!�	�W����p��"Aп��%���޿�¿����68���WM���/��*�=H=���g��𑿣P��k�ӿ���0�꿄�ۿ�d��f���d.t�&�8�
��ξ�X��~�v���H���*����D����2���'��D���o�J���Ǿ-*�kx2��pl��B���Y����ؿ_�{Y�{
ֿ���6N����l��`@��*��-��I��}z�r����0��:�ܿn��~�迫տ����`R���Lb��	+��� �
þ�����t�EM�[�4���&��%"�.�%�KO1�c�F�4�h��㍾�T���龶����K��ń�Χ�9�ɿ������v����п�R��vi��~d��>�Q1�CO<�j_��[��o&���tο翣F�rH�+�οG?�������T�@�!�P���ҿ�܂���U�
�]��!I�b�>��<�<�B�bzQ���j��ۈ�Y񥾵@о�2�
�/��ue��n���ܶ��׿���A�iX��mʿ����-���k]�;�?�&�:�g�M�B=x�$P��걼�6�ۿ������1俾�ǿ�ˤ��P���.I��Q���/����~��cy����j���X��P�QoO�`W���g�����ᗾ�z������a�u�B�E�|��z����ÿn���f��8f޿������P�}���P�+;�v�=�*Y���:Q��ߌǿ���W�򿯕￳�ۿa7���֘�So��8����ܾ�@��Le�����e��+W�plQ���S���^��s�����-���IȾE���� $���U��ቿ�묿�Ͽ��X�����+�տH���N���m�XTH���:��E�ʠh��᏿�����ҿ�R��  �  ��+;ٿ����F��㤀�x9E�$���M߾�������])V�=4�~����X�����#��S;�^a�w����+��K���9OR��D��mꩿ��ȿTݿ���Щտ�㻿>����x�[�G�nC+���%�3q8�4�`�}<������ɣ˿W�޿��xӿ�����j��xZm�O�4�t��;f��z���L��R/��#�$;�Ҭ�m�!J,��IH�# s��,����ƾk�#�.���e��W��]���L�пYZ�yd߿Xο�,��xn��u�e��g;��&�k)���C�h	s�r}���N��!wԿ���W�߿AͿ�_��-̍�s}\���'��8��n�¾X�����w�^Q��8��+�8;&��)�y�5��K� �l��l��g���ip�ȃ�D�F����lI����¿yJۿ8��]%߿{HɿvW���
����]�4/:�5-���7�1|Y��)��t^���ǿ�z޿�,翜�޿�[ǿ܉�����!P�8r�!9��7��m��������b�:nM���B�d�@���F��U��o��Ɋ�%/��о���Ā,���_����_����`ϿI�����~�ܿ�Xÿ4@���1��e�W�z�;��u6��I�S�q�ؚ��ZX��WԿw�������ۿ!���*�����}��)E�rb��f��3��Ӗ���`o��]�<T�ۈS��M[��9l��)��ŧ���\��C羗��?�Sv����뼿��ؿ��ֻ�P]ֿۈ��nȘ�o�v���K�m�6���9���S��R��Y��ɧ���ۿԖ�]�濂�ӿ3鵿�O�� �i�:�4�3���ܾ�c��}I��C���3j��\[�&�U���W�u�b�djw����r����Ⱦ�'���!�7Q���vh���ǿAl���꿸9�OοN��)�r�g�h�C�M�6�O3A�w�b�ɭ���ȫ��[˿����  �  E.ɿ����&𭿧����=l�w�8�C�d�۾(M���&��n�c��GB��4,����O��L&"���0���I��_n��~���n��q��iX�^�C�ly�x�������q%ſaKɿ�̾�d���^����.c�Sn8��G�ԛ��*�HkN�*Q�������4��k�ƿ��ȿ���` ��c����G[��t*�V��si̾��������
[��`=��{*�v!��j �|�(�?H:��lV����)���7ƾ���� %���T�o0������������ǿ�ǿ/2���`��}����R�:�-��"�@��n5�r^�/���������3ʿ�ǿ�ͷ�{m�����5M�ߛ�� ���eþh��	}���_��F��48�!�2�'~6��C��9Y��z�O��j}����"���;���m�f~���"���+Ŀ�%Ϳ%qǿ5���N��N|�J�L��`-�-�!��b+�I��8w�*���1貿ǿ+�οD?ǿ�b��I7���(w�DpC��/����Ua¾�u��d����=p��[���O�]JM��S�c�,*}�bo��"���[Ѿ�]�7�$��Q�����BV��Z}��f̿�Zп�ƿ-��;b��z�r�WkH���/��+��{;�5_�����������=�οrVѿ�Uſ�L��������k���:�W�����¾�O��힍��m}��mj���`�F`�6�h�7z��:���[Y��p�澤���i5�4e�Fh���꪿��¿'Eп?tϿڊ��ѹ��Je���ic��>��+���-�E�D���m������୿�ſ�ѿؖο�d�����>:���:Z���,�~	�(@ݾ���8ٛ��ˈ�,�w�>xh�5b�8�d� \p��Ȃ����0q��
z˾�w���,TE��.x�M���~F���Oɿ�Eҿ�̿���������gV�L�6��K+��4�*+R��������'1���<˿�  �  R���s6��v��.�|���P�	)�����3ܾ󿴾s������gG]��E�K�6��3��9�+8J���d��n���w������=��2�`A[���������Ӥ�,ا������!���'p��D��="�����	��@�[4��e\����Ԙ�⤥�#���ڵ���9���Lo��/D�3U�ca����Ͼ�櫾(_��4�v���W���B��7��7��@��iT��"r�2F��Yާ�a�ʾs����;?���i�욊�3���e㦿H���R���ˆ���`���7�F_�xj
�
�����z<A�Csl�@����)��dܨ��I��z ���ԇ��c��:��������Өɾ����C.��{��g`��O��gI��cM�7�[��s�d(��z꡾d���65澑_���,��T��������I�H���I��^���[��45Z�x&4�^��7V��.� U1���V�	����9��������Y���/���$ჿ�[�9�3�����"���ʾo��+l��}���1�s��f�o�c��$k���|�4���&��X��,\ؾQS����Ƨ?�E�h��{��Ig�������䮿����}���xX��WT��!2�
���K�C�'�ðD��m����L2���������	��ׅ�������T���.����n�26̾ɐ�������䋾�P��w�w���v�EF���+�����8\���Ⱦ�	뾄��qX*�fsO��.z��ڒ����1��,c����������Nq��H���)�x�����@h/��P��n{������3����������`����\��?�p�`G���#�s^�e��͝¾І�������Ȉ�����x�h�{�"����.��
꠾E����Ծ/���ȫ���6�,T^����������(Ѱ�m5���j��uX��Ed�q�=��G$�3���u"��q:���_�R���{���<���  �  ���Oⁿ�6p�T�T���7�A1�z�����)ɾv���tΗ�⪄��!l��'Z�JU��d]�uSr�A���*��!����tоX��F���q#�o�>�S'\�Iv�E����1��ת}�� d�GvC��#��		�����$� �j��;�4��+V�L�s�t�����T��I�h��rL�{�/�@Q�H��Q߾����骨��㒾z���5h�$-Z��TY���e��8~�Y��皥�<h���۾A��A��5,���H��?e���|��ބ�������u�� Y���7�<&�T�@��l�R�p� ��0A���b���}�[I���Ӆ��)|� �b���E�*�`��u����۾�C��Z}���b������vt��ik�1:p����8���7����ЇԾ.A����0"��<�|�Y�S\u�����!���a����t�=V��5��z��6�k9��e*�q����2�� T��s�+����u��rT���({���_�}�B��(�������{?߾��ľ�i��q���4n��V���t˂�gm��6_�����J��V}Ͼ�K����Qi�Z1�}�L�R�i�v��Q����:�������r���R��2����+}	�n���"��'�vE���f��B���ϋ��؍��1��H�y�u�\�?@�Ұ&��c����EL⾮�Ⱦ����������������͒���`[��u�ž��޾�c������#�K�<�=�X���u�����L*������<��S�i�1yH��)�z���"���W���0�}	P�v�p�JㅿJ������v�����o���R��7�
��4������پ%���HZ�����#��/b���Q��6×�0量Y¸��cϾЖ龆��A��v,���F�p�c�-��R:��`G���~����`���>��/"������>f�'��G�;�(�\��W|��щ��  �  �CN�M��0D���6�b�(�G5��=�>��;���־?T���c����
������!� ��ݪ�o�þ�fݾ�[�����b�s��gd,���:��G��O�r5N��C�N1��������y��ɾN�ž|Ծ ��՟�;S'���<��K��0P�L�JA��H3��%��<�)��v���龽eоXﶾH�������	c��]���ꕝ�I޳��;������e�
�h��#��1��+?��J�ewO��`K���=�mL)����)���N�־.�ƾZVɾ�޾\�������0�ځD�qfP��R�L��?�~�1�r�#�"��y�Г �ڷ��OϾض������e��6��AS���`���¯���Ǿ5�K���S
����Ƈ!�e�.�� =���J��kT�F�V��nO��N?�U)�)������c߾�Aվ�)޾w�������n(�24?�<�P� Y��
X��'O���A��~3�%&��-������M�d�ӾY���H���S���3���f��#��onľ�ݾ.���6��f�>���P,��:�u{H��CU��\�CA\��R���?���(�WG�%������D��.���z
�<7 ���7��9M�I�[�+�`���\���Q�v�C���5�ƛ(�N���L��#�S��׾���嘮�*㤾mN���쬾U����Ӿ�"�b�O���2�&��e3�zA���O�[�d`���[��uN�d�9�B9"��0��[�����t��������̤'�!	?��lR���]�)�_�EY���L���>���0�@�$���x�$$�-�辯�Ͼ����j����社B���u*���ƾZ�ݾ�����z��m�N���+�~9��mG��U���^�K�`�٭Y��tI�)Z3�A���:��z� �0��<q��c1�l�G�߸X��  �  H`!��#&���'��'�r�'�i�'��)&��>!������	��>��hҾ+趾c9��S���J��������پ�N�������5#�6O'�w(���(�)�(�#Y(�kU&��� �r���&��Ĩξ����@����ӡ�'��4¾��ྈ	�F������$�d,(�<)���(�
)��(��&�������T����龷6ʾ�u��n����ڢ��0���ƾl��'�����X�1/%�q�'��(��f(��a(�p�'�H�$�t�B���[�\���ľ� ��/Ǣ�r֤�����C�;���%t����D�"�x#)�/�+�5,,�?5,�PC,�xe+�:�'�3��n��� ����jmɾ�s��[�����ӄ��
�۾�����2������'��c-��^/�؟/��/���/�c.��)*��!�,~�ȃ�w!辻�˾����(���'�����ʾ']��s�?�5�"�S=,��1�ǣ2��2�V�2�>�2��1��8,��"��)����/^�P;ξe＾�6�������վ_K󾡖
����(��0���4��6��*6��@6��6�5.4���.�B�$�����a���ӾGcľ������̾���� ����7d!���-��_5�Y�8�6�9�-�9��{9�@�8��a6���/���$�a����:�kѾ�þ��¾�Ͼ��F��r��J�"��z.�a5�bB8��8���8���8��28��$5���-��7"�������K��4ξ|�¾�ľҕҾ��Q����1p%��B0�ip6�<�8�;99�89� B9��_8���4���,��` �#��/�������̾�þ��ƾ�a׾� � c	�����7(��G2��7�i�9���9�X�9���9�E�8��{4���+�����������'߾?�˾Fľ�Gʾ��ܾJ������_W�@�*��  �  T;������iI)���7���D�\�M�PN��kE�g�3�tG�'��|�.2˾8�þ��Ͼ0�쾱'�R�"���8�0�H��wO���L�'�B��65���&�=��'�ۣ�rl�Ծ6���a�����N���_���+׊��X������Rɾ���x��U	�5���]!�8D/���=��I���O��M�YvA���-�gK�>U����۾[@ȾE$Ǿ��ؾ�����|��+��O?��GL���O�%AJ���>��J0�%:"����k�	�����\���ʾ���v3���V��٧��zH���������j����վ���wR�������)�Q7�|LE�a�O���S��N��>?�X�)�/|�)���hkܾ�2Ͼ�Ծ���!�	�:!��}8�K�U.U�w�U���M�3A��2�c%�E�������"'뾧�Ѿ�9���kB��n���5������󹾶�Ҿ����,�Q������&��F4�ŬB�X�O� �X��JY��zP�3 ?���(��f�v������2�۾��羱��^��{�/���E�y�U���\�3ZZ��P���B�
�4���'�������:����nؾQX�����F������.������о�(����b�����|%�K�1���?�bN��Z��@`��]�4�Q�"�=��U&���������,辐����?��{#��;�GbO��g\���_���Z��N�Y�@���2��&��u�8���������Ҿ\���R���.���C��Pm��bC��\ؾ<��������L��)��6��OD�[ER���\���`���Z���K�:�6������	�I������bM�	��G��D,��QC�g�U��_��`��3X�L]K�=��q/��H#�����2��������b;����_L��34���l��uc���N˾_��^c���K��  �  <i�g���w��w9�y�V�<�q�
Y���$������Ah��`H�+�'���=����꾱��Q���.�RP�`�n����4r��E����l���P���3������������ž�������;���j���Z�{X���b�Qay�K�����4m���־A���_���K(�QD��Sa��Zz�����qۄ��z��-_�G&>��m����e�+��ܦ��#��E:��p[���w��6��r䄿V*|���c���F�ا*��������%�ؾX���ͣ��莾H[|��6e��mZ��]��m�����L�������.Ⱦ�Y��g���}4��TQ���m�|��iY���턿�/v�]ZX��47����-o��_�����*���\*�".K�7�k����������ˆ�v�{�Иa�{D��()����>R���ݾ��¾���9	��������~��Mx�J�P���	��t�E�ľq�߾�;��#���x)��vD���a�՞|�g҇���������rs�öS�;3�I��Z�]l�$�	����QP;���\���{��������S����Rz�wt^��A���'���������B⾒�ȾB-���O��e&��ܻ���ˋ��v��,=��� ���þ�۾����
}��� ���8���T���q�[��wҌ������Q���Bo��/N�7n.����N(��d�����+��CJ��vk�F���F��9���&4��=4t��]W��;�RI"��������0ݾ߀ľc�� Z��6d��L����P���������|���ʾע��� ��H���'�J�A��L^�ͦz�����ō�_N��3i����d�"�C���%�^w�����
�/�I�5��HV���v��뇿�䍿�����%��C�k���N��3��*����3��׾��ϫ��a���c��Q����̑��E���L��|Ͻ�g	վ
���  �  �6޾il	�s�*�PS�zL�+3��]䢿pɧ�P��X&��sw���J�w&��e�y���A�P�-�؆T�p��������飿Q�T���L��23v���J��#�����B־}����ԓ��{�>[���D��68��6�@#>��nP���l����T����ľM���
���8��c�lt������uO��+j���Y���ˊ�M�h��x>�k������+��$:�վc�gL��������zͦ�W�������_g�b�<�_�4M���Ⱦ���������o�4!S��@�u�8���:�Q�G�ެ^����Y֕�k��I�׾���P#�X�I�%u�����2������{���̙�����8^�L�6�̹�������)�ЇL�nvx��N��v���G���������p�-�_�<7�9��&y�DJʾb�� Z��I���##j�v"[�hV�H\���k��ꂾ�񔾐���x�˾����i���5��P^�1#�����t^���H���ڦ�����1���hV�a2��/����T���9�F�`�e������>r��t��� X������ⁿKGX��n1����.2�n�̾��O��'����‾agv�P9u��?~�N������ ���trľ�澄	�Ƣ%���I�K�s�檏�k���fr��Ń��+k��֒�>�x��xN���-�'��
��+�;J�ӻs��N��s���<���+㮿/��i���J�w�_9M���(���4��#uƾ-���8������{��%�v�7x��ρ�蠌�vy���ͱ��;yy�	R�9g0���V�����Xz��s������wd��E�������j�M�B���&�h�R=�B�4���W��Ё�<Ǘ�"Ө�u����﬿K4��d��FAj��^A�����F�޾�i���q��Ya��yw��������{��!��	����"�������'��E�۾�  �  :l޾)�;��Lo��_���X���¿�IɿF#��ϐ��J*����j���=��q!��F�8'&�\�F�,�v�ۥ���#��jbĿ`Xɿ�����N��9�c�d1�A��M8Ծh-��C↾�`�܌@��&,�ZU!�bx�u&���6��*Q�MEx��������:�����}�L�����Wl������ǿ9�ȿ�󻿱\��%���H[�+3��1�`����/�D�U�H�9��0�����ǿ2�ǿ,����?������6�Q�٥"������ þVԚ��R|�DT�,W9�&)�B="��n$���/�IoD� d�R��� ���דԾ{V���/��wa�W���
.��gÿ��˿��ǿ�򶿖'�����~P�O".��$�?+%���?�<nk�2�������¿�̿��ǿ;ε��m��M[}��OH��]�T�����¾5���������g���P�)�C���?�^�D��R�$�j�����Q��y�þ�J���(�1F�QOz�Sݙ�vӴ��.ȿ5�οȯƿ�-��ږ� v��pI�Z7-�~*%�^+2���R�آ��\ꝿ'���4�ʿ~�ϿxOƿvװ�h��(iq��0?���\!�zþ���W���G|��i�qP_��y^��_f�.\w�v>��!	�����:#���A,/�$T]����������I0Ͽ,�п�Ŀ�f��F)��EHk�?C��&-���+���?�?�e�v쌿�;��S���9�Ͽ��Ͽ����d���͌�%Qb�(3������㾷�������$d��5.y��h�@`��Pa��Nk���~�Ք������&�þ�e�$��`=��on��p��*���)ƿkѿu!οs2��KV�������\�!":�]+��0��7K�i�v��Ζ�`���0Fȿ�ҿ:Ϳ����ٗ��j؃�רR���&����l׾�N���������Z�w���i�I	e�gi�[;v�#����嗾һ���Ӿ�  �  �O�m��|,H��m������ˏÿ�;ڿ���rؿǁ��འ��ـ��N�
�-�u�$�I!3��&X�5���$8����ƿ�1ܿx��8�ֿ1a��?Ҝ��Vw���<��L�a�־V1��C��>)R�Bk2���W�R���O�)�(���B�jFk��v��3���m��''�\�\����n����Ϳ�;߿�1�Rҿy涿�?��s�o�߻A���(���'��=��yi�R����G���Ͽl,࿉� �Ͽf���J���P�b�R�+�0��aþF���1�o��9F��+�5��f����m"�}6��7V�Cǂ�F)���,־�,���:��
t�h���_����jֿڢ���߿e4̿�>������J�b��{;��v*�M@1��;O�����B��:�����ٿ�[��߿�wʿ��������:FV�T�#�֤���[��ܙ��}�z�Y�0/C���6�\S3��8�;dE�Ѩ\��R������<����0��ɻ!�m2S�j�w���
ɿ�߿�r���ݿm ƿHo�����éY�H�9�jj0��?��Bd�׍��s���LͿ��Z���>ݿAĿ����_w��$�J����k��x���̝��V��n��p[�DZR�|�Q��Y��^i�t��������9�߾�L���7��m��L���ط�g3տ>]�J�}bڿ��C�������Q���8��z7���M��py�L����I����׿P9迣2�-�׿w"������M�r�M<�����'�<\��R���O���9k���Z�'�S���T�S�]�ҳp�ޑ�������p�����`���G����h��n_¿��ܿ���C&��mҿ�g��������n��xG��Z6�o=���Z��_���㥿:ƿ�J߿�꿄��r�Ͽɼ�� $����`��-��%���վ}4��5꒾ʣ��r�i�C�\�[X�+\���h�b�~�!��'^��ڠѾ�  �  kM��d� 3M�dz���ɩ��˿K�⿪뿼	�X�ǿhp��C���%�S�x52�	�(��7��p^�P'���I��@�ο~��.��߿�ĿC<����~�TlA������׾���X�~��N�e.��h��_�����_m$��>� �g�c�����xb��e}*�o~b�<���|
��Bտ/,�0:�Q�ڿ����~e���v�f�F�-�e�+���B���p�:���繿�׿:)鿼鿈�׿����?W����h�Z�/�-��1ľ�ĕ��!l���A��1'����������7��%2�qR����ʀ���U׾�5�?�>��{�C0����¿��޿ķ�-���Կ����G��D-i��A@�~.���5��T������å�~�ǿ^_��r�*q迬!ҿ͔��6��A�[�Nu&������c��䎘���y�'iU��>��2�C@/��3�NA��JX�z�|�폙�uZ��.���d$��8X������G��X�п�k��𿥗�]uͿC"�����&_���=��j4� �C�A�j�mG�������Կ;k뿴�񿣼忦;˿����?%���O�oT�������H4���@����i�7!W�x0N���M���T���d�K�����;i���%ྚ��1;�Ss�0욿�?���,ݿ�M�R򿩟�'�ſvi���t��*�V���<�g�;�j�R�%@�� ���/�����߿�5�1�U�߿ƺ��K����Gy�3�?��A�5��i������*����f�+�V�pmO��hP�ΪY�bQl�ww��&���^ƿ�D �i���K�����럦��Wɿ-忭�}�F>ڿ&���U_���Au�y=L��a:��WA��`�uW���f���;Ϳ��������nP׿����a��2�e�r�0�.L���վ款I�&�|�6�e�ѠX�BET��X�(Hd�ܚz�}������wѾ�  �  �O�m��|,H��m������ˏÿ�;ڿ���rؿǁ��འ��ـ��N�
�-�u�$�I!3��&X�5���$8����ƿ�1ܿx��8�ֿ1a��?Ҝ��Vw���<��L�a�־V1��C��>)R�Bk2���W�R���O�)�(���B�jFk��v��3���m��''�\�\����n����Ϳ�;߿�1�Rҿy涿�?��s�o�߻A���(���'��=��yi�T����G���Ͽp,࿎�&�Ͽm���R���^�b�]�+�&0��aþ=�����o�9F�M�+�C����Y���j"��z6�4V�ł��&���)־+�ܷ:��t�_���S����iֿ���߿�3̿=>��1�����b�t{;��v*�@1�<O�ᣀ��B�����|�ٿ�\��߿�xʿ�������*HV��#�����d^��]ޙ���}�+�Y��0C���6�pS3��8��bE�A�\�.Q����������o-���!�v0S�]�v���	ɿ�߿r���ݿ�ƿ�n������7�Y��9�oj0�	?�xCd�z׍��t��IMͿ��]���?ݿ`Ŀ����rx��'�J�p�	o��{���Ν��X��ln�s[�p\R�0�Q�:Y��_i����������[�߾�L���7��m��L���ط�g3տ>]�J�}bڿ��C�������Q���8��z7���M��py�L����I����׿P9迣2�-�׿w"������M�r�M<�����'�<\��R���O���9k���Z�'�S���T�S�]�ҳp�ޑ�������p�����`���G����h��n_¿��ܿ���C&��mҿ�g��������n��xG��Z6�o=���Z��_���㥿:ƿ�J߿�꿄��r�Ͽɼ�� $����`��-��%���վ}4��5꒾ʣ��r�i�C�\�[X�+\���h�b�~�!��'^��ڠѾ�  �  :l޾)�;��Lo��_���X���¿�IɿF#��ϐ��J*����j���=��q!��F�8'&�\�F�,�v�ۥ���#��jbĿ`Xɿ�����N��9�c�d1�A��M8Ծh-��C↾�`�܌@��&,�ZU!�bx�u&���6��*Q�MEx��������;�����}�L�����Wl������ǿ9�ȿ�󻿱\��%���H[�,3��1�b���/�H�U�K�9��5�����ǿ<�ǿ8���@������Q�Q��"������ þFԚ�R|�DCT��U9�R)��:"�k$�!�/��iD�1d�#�������ԾBS�p�/�ta�\���,��w����˿R�ǿS�z&���񀿞}P��!.�w$��+%���?��ok�3��A��;�¿ѿ̿��ǿ>е��o��A_}�fSH�Aa�l�����¾����x�����g�#�P���C���?���D���R�%�j�r��PM��@�þ�D��&%�hF�GKz�<ۙ�_Ѵ��,ȿ\�ο&�ƿw,���ؖ��}v��oI��6-��*%��+2���R������띿������ʿi�Ͽ�Qƿ�ٰ����Hmq��4?�����'�þܫ��[��|N|�i��T_�}^�9bf�^w�.?���	��E	��z#���N,/�*T]����������I0Ͽ,�п�Ŀ�f��F)��EHk�@C��&-���+���?�?�e�v쌿�;��S���9�Ͽ��Ͽ����d���͌�%Qb�(3������㾷�������$d��5.y��h�@`��Pa��Nk���~�Ք������&�þ�e�$��`=��on��p��*���)ƿkѿu!οs2��KV�������\�!":�]+��0��7K�i�v��Ζ�`���0Fȿ�ҿ:Ϳ����ٗ��j؃�רR���&����l׾�N���������Z�w���i�I	e�gi�[;v�#����嗾һ���Ӿ�  �  �6޾il	�s�*�PS�zL�+3��]䢿pɧ�P��X&��sw���J�w&��e�y���A�P�-�؆T�p��������飿Q�T���L��23v���J��#�����B־}����ԓ��{�>[���D��68��6�@#>��nP���l����T����ľM���
���8��c�lt������uO��+j���Y���ˊ�O�h��x>�l������0��$:�ݾc�lL���������ͦ�h�������_g���<���bM���Ⱦ���K����o�pS���@�ݐ8�	�:��G��^����`Е��c��%�׾-��K#� �I��u�����/�����E
��˙�T~��}6^���6���m��p��.)�ÉL�"yx�DP��3x��7J������J��D�����_��7���ԁ��Qʾ���_�����.(j�%[�QhV�
\�K�k�炾�씾d����˾���e���5�PK^�H ��1����[��iF���ئ�2���0���fV��2��.�����T�T�9���`�� �����t������Z������偿MX�qt1����;;�]�̾����GU��ח���怾bmv� >u�TC~�������������rľ4澠	�ע%���I�N�s�窏�k���fr��Ń��+k��֒�>�x��xN���-�'��
��+�;J�Իs��N��s���<���+㮿/��i���K�w�_9M���(���4��#uƾ-���8������{��%�v�7x��ρ�蠌�vy���ͱ��;yy�	R�9g0���V�����Xz��s������wd��E�������j�M�B���&�h�R=�B�4���W��Ё�<Ǘ�"Ө�u����﬿K4��d��FAj��^A�����F�޾�i���q��Ya��yw��������{��!��	����"�������'��E�۾�  �  <i�g���w��w9�y�V�<�q�
Y���$������Ah��`H�+�'���=����꾱��Q���.�RP�`�n����4r��E����l���P���3������������ž�������;���j���Z�{X���b�Qay�K�����4m���־A���_���K(�QD��Sa� [z�����qۄ��z��-_�I&>��m����	e�3�����#��E:��p[�ȯw�7���䄿|*|��c� G��*���֔��;�ؾ�W��:ͣ�莾 Y|��3e��iZ��]��m��{���E��W����%Ⱦ�O�p�@��Cw4�LNQ��m�K��vV��넿:+v��VX��17��~�%n�U_�������<_*�T1K�N�k�1���y����Ά�#�{���a�сD�/)�����\��@�ݾX�¾M����������,�~��Mx�NG�i������b쬾��ľ+�߾�0���Mr)��oD��a��|�χ�������<ns�A�S��3����BY�kl��	����S;���\�m�{�_�������Ç��Yz��{^�.�A�W�'���������L��ȾY4���U��+�������΋�)y���>���!���þ��۾����+}��� ���8���T���q�[��wҌ������Q���Bo��/N�8n.����N(��d�����+��CJ��vk�F���F��9���&4��=4t��]W��;�RI"��������0ݾ߀ľc�� Z��6d��L����P���������|���ʾע��� ��H���'�J�A��L^�ͦz�����ō�_N��3i����d�"�C���%�^w�����
�/�I�5��HV���v��뇿�䍿�����%��C�k���N��3��*����3��׾��ϫ��a���c��Q����̑��E���L��|Ͻ�g	վ
���  �  T;������iI)���7���D�\�M�PN��kE�g�3�tG�'��|�.2˾8�þ��Ͼ0�쾱'�R�"���8�0�H��wO���L�'�B��65���&�=��'�ۣ�rl�Ծ6���a�����N���_���+׊��X������Rɾ���x��U	�5���]!�8D/���=��I���O��M�ZvA���-�iK�AU����۾b@ȾN$Ǿ��ؾ�����|��+�P?��GL���O�NAJ�ؑ>�,K0�Y:"������	�����B�侥�ʾ� ��C2���T��^���"E���������c���վ����L���������(��I7�3EE�p�O�`�S�F N�(:?�z�)�@y�"���.iܾ&2ϾS�Ծ��쾛�	��=!�]�8��K�{4U�J�U���M��A���2��"%���Ӓ�q��0�ͼѾK���Җ��ID�������3��Ŗ���ǗҾ+�쾦'�6����=�&�?4�	�B���O�ބX�mDY��tP�u?�ĕ(�*d�����'��P�۾��羥��P��p�/���E�`�U�w�\��aZ�L�P���B��4��'���������'�&ؾ�^��o���w��T���e1���	��g�о�)�)��b����}%�T�1���?�cN��Z��@`��]�5�Q�#�=��U&���������,辐����?��{#��;�GbO��g\���_���Z��N�Y�@���2��&��u�8���������Ҿ\���R���.���C��Pm��bC��\ؾ<��������L��)��6��OD�[ER���\���`���Z���K�:�6������	�I������bM�	��G��D,��QC�g�U��_��`��3X�L]K�=��q/��H#�����2��������b;����_L��34���l��uc���N˾_��^c���K��  �  H`!��#&���'��'�r�'�i�'��)&��>!������	��>��hҾ+趾c9��S���J��������پ�N�������5#�6O'�w(���(�)�(�#Y(�kU&��� �r���&��Ĩξ����@����ӡ�'��4¾��ྈ	�F������$�d,(�<)���(�
)��(��&�������U����龻6ʾ�u��u����ڢ��0���ƾ���5������X�R/%���'��(��f(�b(���'�l�$�t�8��{[�W[㾜�ľ�����Ģ��Ҥ�_�_�;��o����7�"��)��+��$,��-,��;,�p^+���'�������
��
��aiɾaq���Z��m�������۾����A7�ӥ���'��j-�)f/���/��/��/�;j.�H0*���!������.'辐�˾����R������ �ʾ�W�p������"��6,�z1��2�,�2�d�2���2�c1� 2,���"�@%����X龭7ξ���6�������վCQ󾕚
�����(���0�P�4��6��26��H6��6��54�V�.�:�$����7f� ��Ӿ�gľS����̾�
�y� ����d!��-��_5�i�8�=�9�0�9��{9�@�8��a6���/���$�b����:꾀kѾ�þ��¾�Ͼ��F��r��J�"��z.�a5�bB8��8���8���8��28��$5���-��7"�������K��4ξ|�¾�ľҕҾ��Q����1p%��B0�ip6�<�8�;99�89� B9��_8���4���,��` �#��/�������̾�þ��ƾ�a׾� � c	�����7(��G2��7�i�9���9�X�9���9�E�8��{4���+�����������'߾?�˾Fľ�Gʾ��ܾJ������_W�@�*��  �  �CN�M��0D���6�b�(�G5��=�>��;���־?T���c����
������!� ��ݪ�o�þ�fݾ�[�����b�s��gd,���:��G��O�r5N��C�N1��������y��ɾN�ž|Ծ ��՟�;S'���<��K��0P�L�JA��H3��%��<�)��w�����eо[ﶾL�������c��i�������^޳�;��������
�:h��#��1�,?��J��wO�aK���=�BL)�F��������־��ƾ�Rɾ��޾t��,����0��|D�o`P�m�R��L���?�"�1�R�#�r~�h�~� �ݮ辯HϾҶ�!�wc���5��|T���c��Uǯ�F�Ǿs�L���%
���܎!���.�(=�J�J��rT���V�9tO��S?��X)�������e߾'Bվ(޾����@���j(��/?��P��Y��X��O��A��v3��&��&����X��D�X�Ӿ�S��E��<R���3���h���&���sľQ�ݾw���Ô�jl�T  �PX,��:�o�H�TKU���\��G\��R���?���(��J�����?�龓�b1���{
��7 ���7��9M�y�[�E�`���\���Q�x�C���5�Ǜ(�O���L��#�U��׾���昮�+㤾nN���쬾U����Ӿ�"�b�O���2�&��e3�zA���O�[�d`���[��uN�d�9�B9"��0��[�����t��������̤'�!	?��lR���]�)�_�EY���L���>���0�@�$���x�$$�-�辯�Ͼ����j����社B���u*���ƾZ�ݾ�����z��m�N���+�~9��mG��U���^�K�`�٭Y��tI�)Z3�A���:��z� �0��<q��c1�l�G�߸X��  �  ���Oⁿ�6p�T�T���7�A1�z�����)ɾv���tΗ�⪄��!l��'Z�JU��d]�uSr�A���*��!����tоX��F���q#�o�>�S'\�Iv�E����1��ת}�� d�GvC��#��		�����$� �j��;�4��+V�L�s�t�����T��I�h��rL�{�/�@Q�H��Q߾����모��㒾}���5h�/-Z��TY�ľe��8~�%Y������\h���۾w��$A�6,�̒H�@e���|��ބ�������u�� Y���7��%�CS�����h�P��� �--A���b��}��F���Ѕ�#|�R�b�S�E��*�q�Ek��d�۾ <���v���]��4�����s�6ik�Z<p�e��O�������@����ԾpK�P��7"���<�T�Y�cu�����$��'d���t��V�75��|��7��9���)�Е�C�2�V�S�#�s������r��.Q���!{���_���B��(��}�:���%6߾�ľ�c��✛�8k���ބ��˂�o��mb��۳���P��x�Ͼ|U�a���o�&1���L���i�������>�����Z�r���R��2�Z��"	�����#�y'��vE�6�f��B���ϋ��؍��1��L�y�w�\�?@�Ӱ&��c����HL⾰�Ⱦ����������������͒���`[��u�ž��޾�c������#�K�<�=�X���u�����L*������<��S�i�1yH��)�z���"���W���0�}	P�v�p�JㅿJ������v�����o���R��7�
��4������پ%���HZ�����#��/b���Q��6×�0量Y¸��cϾЖ龆��A��v,���F�p�c�-��R:��`G���~����`���>��/"������>f�'��G�;�(�\��W|��щ��  �  R���s6��v��.�|���P�	)�����3ܾ󿴾s������gG]��E�K�6��3��9�+8J���d��n���w������=��2�`A[���������Ӥ�,ا������!���'p��D��="�����	��@�[4��e\����Ԙ�⤥�#���ڵ���9���Lo��/D�3U�da����Ͼ�櫾)_��9�v���W���B�&�7��7�(�@��iT��"r�FF��sާ���ʾ����6�Z?���i�����D���t㦿Q���R���ˆ�O�`�+�7��^��i
�Ó����>:A�ppl������'��ڨ�NG������ч���c��:���E���K�ɾK���*)��P{�Ab`��O�gI��eM�U�[���s��,��G�u���|=�Ad���,�mT�\���������̰������_��n]��t7Z��'4�%��HV�.��S1�h�V�����8�����������O���=ރ�q�[���3������V�ʾ3 ��;g��֘��i�s���f���c�E'k��|��7���+���	��dؾ�W����S�?�$�h� ��Dj���ī�,箿9Ħ�~����[�BZT��#2�����L�,�'�k�D�m����d2���������	��م�������T���.����n�56̾ː�������䋾�P��x�w���v�EF���+�����8\���Ⱦ�	뾄��qX*�fsO��.z��ڒ����1��,c����������Nq��H���)�x�����@h/��P��n{������3����������`����\��?�p�`G���#�s^�e��͝¾І�������Ȉ�����x�h�{�"����.��
꠾E����Ծ/���ȫ���6�,T^����������(Ѱ�m5���j��uX��Ed�q�=��G$�3���u"��q:���_�R���{���<���  �  E.ɿ����&𭿧����=l�w�8�C�d�۾(M���&��n�c��GB��4,����O��L&"���0���I��_n��~���n��q��iX�^�C�ly�x�������q%ſaKɿ�̾�d���^����.c�Sn8��G�ԛ��*�HkN�*Q�������4��k�ƿ��ȿ���` ��c����G[��t*�V��si̾ �������
[��`=��{*�|!��j ���(�OH:��lV�(��
*���7ƾ:���� %���T�{0��ɩ��������ǿ�ǿ/2���`��h��L�R�Ȃ-�K"�V��35��p^�.��R���1�2ʿ:�ǿ�˷�~k������2M�y�����u`þ�c��yy����_�U�F��28���2�^6��C�{>Y�A�z�]#��]������o��7;�p�m�m����$���-ĿY'Ϳ�rǿ����g���|�b�L�Fa-�:�!�9b+� I�#7w�����沿uǿU�οF=ǿ�`��55���$w�|lC�(,����\¾uq��򉈾�8p�t�Z��O�zJM���S���c��/}�s���#��<aѾ�`���$��Q����kX�����y̿�\пr	ƿ���qc��k�r��lH�͇/��+��|;��_�=���������G�οwVѿ�Uſ�L��������k���:�X�����¾�O����m}��mj���`�F`�7�h�7z��:���[Y��p�澤���i5�4e�Fh���꪿��¿'Eп?tϿڊ��ѹ��Je���ic��>��+���-�E�D���m������୿�ſ�ѿؖο�d�����>:���:Z���,�~	�(@ݾ���8ٛ��ˈ�,�w�>xh�5b�8�d� \p��Ȃ����0q��
z˾�w���,TE��.x�M���~F���Oɿ�Eҿ�̿���������gV�L�6��K+��4�*+R��������'1���<˿�  �  ��+;ٿ����F��㤀�x9E�$���M߾�������])V�=4�~����X�����#��S;�^a�w����+��K���9OR��D��mꩿ��ȿTݿ���Щտ�㻿>����x�[�G�nC+���%�3q8�4�`�}<������ɣ˿W�޿��xӿ�����j��xZm�O�4�t��;g��z���L��R/��#�(;�֬�m�)J,��IH�1 s��,����ƾk�-�.���e��W��d���S�п^Z�|d߿Xο�,��nn��P�e�Gg;�ǉ&��j)� �C��s��|��BN��XvԿִ�[�߿9Ϳ�^��*ˍ��{\��'��5����¾���	�w�L[Q���8��+� ;&���)��5� K�`�l�o������gs�}��'�F� ��|J����¿�Kۿ0��9&߿5IɿX��)����]��/:�;-���7��{Y��)���]��.ǿ�y޿�+翏�޿mZǿƈ�����P�pp��5�����0��������b��lM�ܹB�s�@���F���U��o��ˊ�}1��� о�����,���_���������aϿa�����e�ܿ�Yÿ�@��&2��1�W��;�v6�5I���q�횕�hX��_Կ|�������ۿ"���*�����}��)E�rb��f��3��Ӗ���`o��]�<T�ۈS��M[��9l��)��Ƨ���\��C羗��?�Sv����뼿��ؿ��ֻ�P]ֿۈ��nȘ�o�v���K�m�6���9���S��R��Y��ɧ���ۿԖ�]�濂�ӿ3鵿�O�� �i�:�4�3���ܾ�c��}I��C���3j��\[�&�U���W�u�b�djw����r����Ⱦ�'���!�7Q���vh���ǿAl���꿸9�OοN��)�r�g�h�C�M�6�O3A�w�b�ɭ���ȫ��[˿����  �  �2�tC+�	������ ���x���1L���J$ܾ���H���]�I�A��3�1/��5�MaG���f��[��؄��ñ�I��=�[�����\�ʿ��<��Fd.�s�2���'�����﫵�
ތ�o9k���b��B������Dhҿ�l��1�ƭ/�e12�&�����;�^���}�Ϝ8�j4�kʾf����}�X6V���>���3��3�v�<��aR���v�(���þ V�1�1���t������sݿ�j���#��O1��w0�c\!��M�
ؿ��9����c�w�g�,Q��򇰿�;�}��Ew&�}�2��[0�9��*�5�ҿ����y�g��b)�Ap���
��*�����}���]�$�K��sE�c�I��UX��s�eۏ�8~�����K!���L�Z����m{���3� �+���4�O�.����� �mUʿ�����~�VQi�T~z�����ſ�6��%����-�)d5���-�G���r���tÿV둿W�C��#/�<;��;㛾Rǅ��p��b��`���g��Tz��X��
Ȧ��S;�f�>�-�{�i������xѿև��	 ��1��$6� �+��W����ֺ������{���s�/�����;�ڿ��	��n#�f�3��h6�|;*�m���쿢:��s6��� I���l��	������D���)���s�7"s��|�wI��ޠ���c�� 
�%��zB��y��5��������'���5���4���%����࿇f��3���Ct�t�x�7z��@���������*��<6���3��C#��p	�;ٿ������t��u6�I�
���پ�	��f򗾱���c@|�#�t���w��Ђ�G��������ƾe����y!���V�٣�����A������F$.�K87��e1��W�n��2Ͽfe�������r�+�R��U�ɿ�T ������/��  �  �8+�D$�������f�������;H��/�IDܾ=Ʃ��ᇾ�0c�^_G�wf8�Zn4�`;���L��Vl�W؎�����E�[��A/W�k���x�ÿ� ��G2��'��+��!�ӽ�T��������?e�!�\��ly�����ʿ`; �����Z(�}�*�)�R��Z�ۿs���w���5��U�V=˾ើ�7����[�~fD�H�8��H8�M?B���W�,o|��j���ľ|��</��n��š�eտo������)��)������2п�����~�D�]�[b��\�������ܿ@J	�%���S+�%)�$o��� ��M˿�U��B�b��4'�B����m��q���d����7c�7Q�аJ�C�N���]��Sy�e}��4o���?�@���I��燿ӵ��g뿅6�u�$�s(-��'�����+��~`ÿ�ᗿQ�w�S�c��t��3��\��a��.t���&��-���&�����
�u
��"��?#S��!�3P����|��@���d=v��;h��He���l����2!���A��_�ξ�/�c�+���d��\��Phʿ8} �m��'�*���.��$�J���&�f���]𐿔�u�p�m��+�������Zӿ�y������,���.��\#�+&��)�m��������E�0����뾥9��,u�����0M��+y�dx��/�����d^�������f��hO?�4�� ���ݿ�
�Y!��.��L-����H.���ؿ�	���q��Eun���r����+���a�俦�9#���.�m`,�F��<� �ѿ|�����o�7G4��^
��;۾ u�����LK���π�fz��%}�1����ђ��.��9�Ⱦ�2���6 �WS�1���񺿝��G��v'�ʸ/�W4*�O�+��3?ȿ�������Zm�j}�Ҙ��¿W;����Z�(��  �  �������g ��jԿ�����+}��q>�TA�P�޾�԰��̐��u��X���H���D���K�4�^�?�~�8����b��~T쾂��xoK�����ΰ�!߿���Hc����/3�k���olʿӞ���z��T���L�X�e�cg��sN��KB�-�_}�������
d�HsſQ���?lg�%r.�����Ͼ*˦��[��5	n���U��_I��H�EUS�tj�g��ŏ����ɾ�� �٥(�"�_�_��9���
���������A��Tֺ��葿{�i���M�#[Q���t������ſ������,$���������-����U��R"�����VǾ�{���Պ�%"u�Fb�9�Z��I_�5o��х�Lz��mɺ��q����0@��}����x(ӿ  �,j�����$�����ݿ�e��#�be��S��!b��Ї��/���2ٿ6���v�s����Q#�u�ٿP��^
��.[I��3�����1Ǿ`g���ɑ�'䃾�x���u�$�}�M͈�sT���籾*վ6��Ac'�#Y����g���M�忮a�����`�B��
���3ҿ*Ѧ��u����d���]���v��ޖ��ɾ�Ƚ��R���s����������Ϳ�>����w�s�>�=_�!�m#Ǿ���-��e抾d����]��k����%��X���{�¾�꾂���8��p�DP���3ȿ�i��������VK�q��N�`Eÿ~S��v}z�/9^�M�a�S���	����tͿR��[��Y��%��!�Z���1��F�����b��d/�P}
��#ᾩ�������?���>���-���Ԇ�G��!���I1���оei������xJ�1����ͪ��Lؿ'������f�����2�4���G��i�����n��2]�Luk��i��	���;�ݿ��w���  �  ����A���ԿhK�������d�1`4������}f���������by���f���a�( j�����_��'����ʾ�%��=��f�>���q�����5u���ۿ���ϣ��*3鿫�̿�Č���Z��B;���5�z{I�~Au�����R���N4޿ �G��'W��ʿk+��B���AXT�_(������ܾ�K��D���jH��xu�ӳf�	�e�{r�j'��O����J��Z�׾�y�oi#��?N��͂��죿A�ƿ�L俽
���������6��?m����z�v�L�96�P69��U�cs��F0��ʿ��翑h��ƕ��^~�b��Y*���|�jG�v,��T�ڊ־�����휾�S���R��-�w���|�����\��cí�+�˾@#�M��Eg7��{f�� ���N���Bտ�j�	���97��Cۿ<f��$��g[q���J�g�<�2DH���l�� ��*$����ؿ�v���x��;ڿ�Ƹ��7��Ӫo��J?�������`�׾\���2���x��{L���7���MT���@���ľ;��k��1%��ML�ғ�>f���N¿��⿔}�������v�ltԿ(V��`y��Oj�ҹK��6F��FZ�3��9k���/ƿ ��ft��T���E���%ӿ���܎���d��y8�K�7n����ؾ�⼾Qp��P����i�������L���>���ʹ���Ծo�������3���^�/���1��.ϿԤ쿶j���>��p3�F�ɿ"ե�����UN]��F�`�I���e��F���ɭ�jѿ����F���H��/��ǿA���k���C�T�R>,�yV�MU��	Ͼ���^ ��5���沓�����zU���˃þ���I�αA�v�p�i#��]u���mڿ����}����S��,P࿶_���
��M{�nPT��F��Q�V�u�9z�������ݿ/����  �  �^��w츿b����R����y��Q�wt1�c���������Kþ�ǩ��X��s_�������z��^��ei��:Aʾ��mn�bb�[�8�4�Z����9���`��������Y��o���I��0
����\���5����]��w�)�A�I���w�r������r���g���y3��p����Q��o�l��lG��I)�C������پ���<T�����̉��>������ʡ�A���վ�E���z�T�%��)C�\�g��q��F���n��W��� ���W���ؗ��n|��M���+�%.�����2�-�X�Iф�5���rʳ�/B�����4U��u��8`��<�b���?���#������@E־�\���*��m��"���+��rݠ�*����;�A����Ñ���5�ӱU�&�|�t����������� f¿����ց��1b��Pt�� I��,��"���*�@�E���o��T������{����ÿd���{��9И��\����\��_<�ٕ"�����$����پ���������9��UK��(K��~���H6ɾ�便W�M���+�\NF�U�h�������������
�¿=iſ4���P���Q���Έl�:�E�;O/��A+�P:�{�Z��9��8板���*
Ŀ8�ƿ*���?��t����y}��W�ۭ9�0�!�l��pp���Kܾ`{ľO7��n۩��J��U���=���w�ؾZT��L���d)6���S�g3x�`����H��tq��q
ƿ�Ŀ����;��ꕆ�T�^�O{<�S�+���-��B�/$h�U��/ϥ��պ�!ƿj�Ŀ6췿!���~錿��o���L��1����M�� ��qԾ�Ҿ�U5���ܩ�Kj��o���#oʾSz�P� �"W�N�&�l6@�j�_�%����ܙ��᯿������ǿ:���&����`��.�}���R�~6��y+��4��N���x������O�������  �  ?������o)��WJw���a�-N�i~=��.�����Y����־6x�����Υ�������kZݾ�!��Y7��&"�f�1�M�A���R���f�T�|�(����Ǝ�����\r���O��1.���r�������t
�j"!�Z�@���c�d���Ij��O�B��)v�� q���[�^�I�te9�f�)����i�?N��ξ,M��%0���m�����ʾ�0龌��iK��'�i37�`G�+Y���m��쁿����t���Ō� Â�+�f�_�C�h�#���9W ��!� D��+���M���p�	�������ܐ�hB���y��o�l���X�5&G�h�7���'�/P�[��@1�%�;ߐ�����=��
>ž�|߾�0 � �{x#���3�U\C���S��g��|���	�d0���������'c��@���"������7��6� �e3>��`��f���F���i��6��'����#���l�&Y��iH�a�8��)������;��Ҿ�w¾���+Jƾ-$ھ
�����1��Y�/���?�'GO�	�`���t�4W��u|��ߕ��ѕ��L������G&_��=�C�"����V�+���1��wQ�F�t�o��tڔ��]��ԧ��_Ӌ�;���F|l�f�Y�/�I��1:��)�E?�����5d־�>ɾ�xȾO*Ծ)��۩�����s'���7�}G�SoW��i�<z~�98���h��pΗ�)#��!���tw�{~T�R4�~������P� �h;��f\�g�������������ؑ�����	z��e�<T���D�%�4��,$�q��ٜ��'���Ѿ��Ⱦ�Y̾�ܾ�����!�b���.�(>�<�M��4^�"Qq��|��G3��#��U]���,��w���-m�,pJ���,��i���������)���F�J�i�z���\���  �  vY��X_���`�`��#`���`�Z[_�J4Y�0L���8��f!��"
�����ԾW�;8پ@q��DQ�6'��=� P�|�[��`�-8a���`��`�Za��t_�C<X��J�Y�5����5���3�Ӿ:�Ͼ	�ݾ����!��H�+���A��S��c]�g\a���a��0a��a�%�a��_�عV�WG��(2��`�6���5徎�Ѿ��о�⾷��v��]Q/�8�D���T�I^�%a���`��`��`��`�R]���S�ETC�x�-�x��9  �P6�udо
Ӿi��H	���65�o�J�%�Y��*b���d�P�d��\d���d���d�<T`���U�ZZD�a.����Ů�I��پ�޾�"����ab%�Y+=�?�Q�*�_��f��Zh���g���g��[h�9�g��ob�{�V�|<D��v-������,߾�����c����,�ND�4�W�%]d�8Tj��k��k�:k���k��Fj��(d��9W���C�y�,�֣��z�V�� ��ٮ��@�J��4��K��]��0i��.n���n��vn���n�Yo��Tm��Lf�\^X�wUD��-����������o#�����}$�a_<��R�m�c��7n��$r�
\r���q�r�Q,r��xo��g���W��RB�g}*�����������������'��k?�U��-e�AKn�kq�.aq�q�vkq��_q���m�m~d��T��'>�8Y&���Uc ����V��qk�H%�M�+�e�C��tX��{g��~o�y�q���q��oq�q�q�ѕq��\m�2�b�n-Q��:��#�������A�����=���K�a0�x�G�w\���i���p��r��Er��/r��r���q�S�l�R�`��lN�.�7�������#�����y,����	�F��P%5��fL�C�_��  �  �.�\0>��O�תb�)�x�j���ꍿw�������V�v�G2U���2�GI�A�X����+�M��d:��J]��~��Њ�n�������脿�Rt���^�o�K���;�}#,�l����
�0p��eҾ�9��tD��?���kH��D[ƾ�㾡���� g%�E5�~�D�d}V�~k�a����7��G���81��\Q���1m�WfJ�XK)�5�����P� �/{�2�%�&SF��5i�EÃ�z^��򕏿ъ��j����l�U�W�i�E�$6��r&����Ms�y�澥�Ⱦ	���x_��Ra��h˸���ѾT#�L�
���kV-��=��tM��$`�[�u������B��r���濍�r���%�e�l�B���#�#!�ϒ���f��̎5���W��Vz�n��S���*��x����e��9�l��X�'�G��Z8���(�����\����}о�߽�!\��Sx���|Ͼ���U�y.�?x)�R�9��/I��Z�F�m�R��3���_��Es�����(��Ê`��[>���!������
��i��u(��G��1j�p���3|��3_���ړ�𾋿����l�2�Y��vI��.:��H*��O�$����Kjؾʾ��Ǿ�Ҿ�n�؞�:���{%��86���E��U�)3g���{�h͈��s��!̗�~W��n��[}�e�Z�C]9�������������H�5��bV��Ny��Ջ��x����W���A����A}��wh�ʅV���F�7���&������v]�	DӾ�8Ⱦ�ɾ�o׾ѷﾾ��3!��*���:�*eJ�i�Z�r;m��H���+��YȔ�� ��P3������Ar��PO��60��2�av��I�q0%���@��b�ȕ��GB��i����V������ʋ���*w��Pc�,BR��B���2�"��l��h�������оe�ɾ��Ͼ�@�g������n �(�1��  �  ��g�2���S��#|������"��G����n��N����У�
����c���:�*� ��q�=8%���B���n�z䐿�⨿$�������7B��� ���⏿Ses���L��p-�a��M6 ��ݾ��/k��a��|�����Q|�����^����aо���Z��"�7O>��a�_	��C����̰��#��켽��ֱ�el��4Ⴟ~�U��1�����1�-���P����c�������CѼ�O����a��ݞ��6���qe�p'A�9$$������`�Ҿ.����`��jܐ�ㆉ��"��z����槾.�����޾E� �����-��SL�1Tr�D/��i�������as��E׼��]��i���y��1L���,��E�[�$�� =���d�jc��-�����������������x���g����_�K>�dM#���$;��#)ؾd���쩾D�� ��������}��~�ؾo:��q<���#�Y�=���^����������k����ÿ���k��&���Gho�hzF���,�it%��c1�<@O��I{��H��$e��#5���iſ�	��Ҭ�E���W����}Z�N;�Ӕ"�v�7����ݾ�ž����������8��������վ���h5	�$�,�2��O��pr��Y��b������Tſ{�ſ�򹿃����̼e��A�{-���+���=�W�`�����J���������Ŀ4�ſ팺�P���s����u���Q�u�4�L��eW
�����׾u�����Z ���)��a�����ž�ݾ�������F�"��:�QzY��f�S���v��T)��*�ƿ�AÿR����H���WdX�[�8�!++�>�0���H�VFp�����}��,ֽ��ǿ��ÿ|@��m+��b���l5j�:|H��-�������L��Ѿ�Y��6���*���5��ǻ���ϾB���T��K��  �  sZ�x�6���g������C��}ֿ�����H��ҿ�K��=����`��>��4���C���k�����_u���ٿn_��������f�Ͽ<˭�����x�\�<:.��v��{㾃��S1�����x�(�g���d��To�؜��%�������Ѿ����$����F�T!|��~��q���}࿎��f�����忖{ǿJǣ�����~~S��8�`27��<O�D�~�㽟�;�ÿe���������D�Ŀ���-���_K��!�`����Ծ����������&�q��f�_�i��z�N׋�QP��*���侌5�G-��4Z��艿����H@οH꿋X�����޿�Ľ�U-��,�v�w^L�:��VA���a�3���~���ѿ���)��<$����ݿ�	���4��_�u��MC����s� �	(׾.���#=��P���6�������0���M���������-�׾�� �0O���A�*�r�^��x���>�ۿ��G=��y��$�׿b ���I����l�m�I�g
@���O��x�Q,��ɽ� �߿����qs���p�ظֿ2��������Dj��<�y�{���5ھ󽽾慨�̚�F2���D������a��(2��A�о���6�.���W��h���ͦ�R�ɿ�����0������>�Ͽ�ԫ���� �c�D�H��5G��@_��J���ħ���˿��꿆��������B�&"ͿB���U����[���1�p8�G���M�Ҿq���l��JԘ�ڒ�3���2���R������5ھ&~������]:��Vg��n��;=��-�Կ��������y�����"�ÿ�Q��p��zcX�~�E��M��[m�%�������P׿���m��`V�����1¿�_�����p�M�RT'��
���뾈�˾��N��R�������%��|F��.eɾ\R辋���  �  �.��IA�܈�����׿����|����=�$����ѿ�9��Ȣ��>�W�
:K���^�󉈿����2Hܿ��>���������L��r�̿z���_2r�a6���
��W׾/���ލ���r��X�ZJ��G�`�P���e���������3�¾����dz!�M�U�G���㜸���������7L�H�����/�¿y}���<r�G�P���N��l��L������z��^�	�r������	�[��h���ґ�g\���%���� �ƾ�H���܅��qh�%S��J���L��Z��Au�;��Ԭ��&׾��	��4��'n��ݜ���ɿ�z���K�s��c��A�[����� Ŏ�23h�HQ��PZ�.d��p����Ͽ�Q��1��
��?��Ϡ�M�ڱ�|���dkO�ͯ������7Ǿ�u���S��`r~��[m�h�19n����YW��d����Ǿr���F%��OL�\��v�����ܿ�G��8����x�/"�;�׿��������zc��(W�\�j�����gി��⿑�[��4��8�� �S�ӿ=�������8D�������ȾU��S��y���J��&���𓈾�o��F����྾>�g��	92�Ǝf�.��m����C￫/����A^�������4�ʿ�����"���`���^���|��P��,�ſc����B����	��+��.�ſc���l�*c6��I�)��S��fd���h��U��wF��Q�Mc��O���Rȫ���Ⱦq���zOA�tD{�n`���(п���f��������/
����"��!є��1t�`/]� f��:��}��8zտ�k��=�j@��&�j6��;����ʼ��$�Y��)��9�~�۾^���k ����������w���,�� ���|�������׾n���  �  k���K��抿op����=���$��C+��m#�K����e���ɍ�
\i�2$[��q�����¿s3��)���s&��3+�t�!�]����x���#��D�>�R����ӾY���҄�2`�k�F���9��V7��?�۔S�@�u�8������`�����&��+c�zG����̿����k�(��w*�33�w��X�ٿ�.��p惿�Ua�cE_��؀�7U��=�ӿ���?�ʪ)���)�����|��jҿ���8yj���+�k����b�����2uy��V��HB���9��S<�b�I��)c�`������Ӿ�5���;�m�~�-ū�C�࿽;�� !���+���(�}��n���{4ʿ����S�{��Ga���k��	��$ʹ��#�ϛ��{#�f�,�x+(���S����'Ŀ2�����Z�ߎ"�{e��ϳ��u������Z�l���\�w�W�ؠ]�-zn��%��?�������;����b ��V��k����$�������'�Q.�o6&�d}�5��Nܼ�򨓿D1u��g���}�5Λ��1ȿ�l����l�)�p~.��*%�k����WJ��7 ���L�y��m0�B^���;��������w���v����pc��,����d���O޾��ys7��s������տ
�����W�,���.�~@"����,�῝6���ꋿ9Zq�/Ho��ڈ��X����ۿѢ�V �S�-�!�-�� �r��%�ڿ�_��{��]<�d��iN�)Ӹ�W1�� `���р�E:x��{y�d�gڎ���������m�d����H����EE����t�5$��/�	�+���t��IпF���7ȃ�]/m�mgw��䒿ꓺ����|a�Z0&�t�/�!�*�6H�x����Sɿ�͘�e�?�,�/��Cվ�ڰ�m显�É��L����|�0ۀ��ψ�[E��-@��Ѿh��  �  t �ЯO��⎿>��0;��Xp��,�x�2���*�����G��ƒ���1����o�r�`��Jx�o����*ɿ.� ��:�/�-�0�2���(������ck��䢅�jFB���RӾ5���(���Z�i6A��L4��2�YS:�q�M�
p�֒�W�������d)�%nh����&DԿ���Dp �E80���1�i�$�~'�K��4魿�ˇ��Fg�Ae�2����Ш�W�ۿ.
��"��1��
1��"���	�Oڿ�/���$p��i.�����H���Ε�o�s���P���<���4��7��=D���]��c�� ����XҾP-���>�Ă�ek��鿞����'�^3��0����S����ѿ����pH����f�Y�q��A��5����Q|��v*��c4�sl/���,C��˿�ۗ��(_��_$�4������D5��xO���/g��SW��R��QX��h�Y����������������!�ѵZ��g��_�ƿV����,���.��5�}I-�6��I���cÿ���{�{��l�E"��W���^GϿ���d��0��5��-,��S��s���<��N��P���Ʊ��Y�����rE��d^~�%�r�-yq���z�*����蘾����^ ݾh�)�9��$y��d���ܿt���$�O4�V�5��)��0���'�Џ�iKw�� u�왌�԰����p��&�M5�[5�޺&�D���0o���U��"�>�"p�80ᾐ����p��z����;|���r��5t�w��H��e����������4
L�>P���귿���7� !+�ފ6�J43��"����ح׿N����D����r��}�f���������C�/,-�?
7�]2�O��E��:п7����i���.�ޣ��}Ӿ�V���������B}���w�nd|����$w��ǭ��vMϾ�h��  �  k���K��抿op����=���$��C+��m#�K����e���ɍ�
\i�2$[��q�����¿s3��)���s&��3+�t�!�]����x���#��D�>�R����ӾY���҄�2`�k�F���9��V7��?�۔S�@�u�8������`�����&��+c�zG����̿����k�(��w*�33�x��X�ٿ�.��q惿�Ua�dE_��؀�8U��?�ӿ���@�̪)���)�����|��jҿ���Cyj���+�q����b������ty���V�HB�O�9�UR<�H�I�'c����{��TӾ�4��;���~�9ī�B��:;�f !�>�+���(�"��ݖ��4ʿ�����{�}Ga�Ôk��	��ʹ�g$�#���{#���,��+(�i��\����(Ŀ ���F�Z�^�"�h�����'���%���l���\���W��]��xn��$��������������a �R�V��j����#�����'��.�6&�
}�����ۼ�����1u��g��}�}Λ�g2ȿRm��U�ݯ)��~.�E+%��k�̎�`K��-��ԥL���3�`���=��K��)��w�L�v�T���c������e��P޾���s7��s������տ
�����W�,���.�~@"����,�῝6���ꋿ9Zq�/Ho��ڈ��X����ۿѢ�V �S�-�!�-�� �r��%�ڿ�_��{��]<�d��iN�)Ӹ�W1�� `���р�E:x��{y�d�gڎ���������m�d����H����EE����t�5$��/�	�+���t��IпF���7ȃ�]/m�mgw��䒿ꓺ����|a�Z0&�t�/�!�*�6H�x����Sɿ�͘�e�?�,�/��Cվ�ڰ�m显�É��L����|�0ۀ��ψ�[E��-@��Ѿh��  �  �.��IA�܈�����׿����|����=�$����ѿ�9��Ȣ��>�W�
:K���^�󉈿����2Hܿ��>���������L��r�̿z���_2r�a6���
��W׾/���ލ���r��X�ZJ��G�`�P���e���������3�¾����dz!�M�U�G���㜸���������7L�H�����0�¿y}���<r�H�P���N��l��L������~��a�	�u������	�h��$h���ґ�|\���%�����ƾfH��]܅�zph�g#S�K
J���L�ִZ��<u���1Ь�"׾A�	��4�Y$n��ۜ��ɿ
y���J���������I������Ď��2h��GQ��PZ��d������Ͽ�R�������1��ˡ�G��۱�G����nO���������;Ǿ�x��
V���u~�~]m�:h��7n�Z�� U���`���Ǿ����`"�6LL����������ܿ�F��7�������!�0�׿������:zc��(W���j����6ᴿ���C�0��5��9�� �e�ӿ:���f��-<D�����j�Ⱦ�X��V��춊��K���������}p������ι�侃��92�Ўf�0��n����C￫/����A^�������4�ʿ�����"���`���^���|��P��,�ſc����B����	��+��.�ſc���l�*c6��I�)��S��fd���h��U��wF��Q�Mc��O���Rȫ���Ⱦq���zOA�tD{�n`���(п���f��������/
����"��!є��1t�`/]� f��:��}��8zտ�k��=�j@��&�j6��;����ʼ��$�Y��)��9�~�۾^���k ����������w���,�� ���|�������׾n���  �  sZ�x�6���g������C��}ֿ�����H��ҿ�K��=����`��>��4���C���k�����_u���ٿn_��������f�Ͽ<˭�����x�\�<:.��v��{㾃��S1�����x�(�g���d��To�؜��%�������Ѿ����$����F�T!|��~��q���}࿎��g�����志{ǿJǣ������~S��8�c27��<O�J�~�罟�A�ÿl��!���#��� �W�Ŀ���?���_K��!�i����Ծ���
��������q�7�f��i��z��Ӌ��K������㾳1��-�0Z�承�����=οsE� V������޿^ý�<,����v��]L��:�FWA�˽a� �������ѿ����+���&��n�ݿ����7��l�u�@RC���� ��-׾簷��@������p�؀��(���K��B�����Y�׾� �K�یA�
�r��������n�ۿR
���:��N��U�׿�����H����l���I�s
@�w�O�"x�l-���ʽ��߿&���v��fs񿺻ֿ���|����Ij��<�N}������ھFý�n�К�5���F��(��c��3����о�� �N�.���W��h���ͦ�R�ɿ�����0������>�Ͽ�ԫ����!�c�D�H��5G��@_��J���ħ���˿��꿆��������B�&"ͿB���U����[���1�p8�G���M�Ҿq���l��JԘ�ڒ�3���2���R������5ھ&~������]:��Vg��n��;=��-�Կ��������y�����"�ÿ�Q��p��zcX�~�E��M��[m�%�������P׿���m��`V�����1¿�_�����p�M�RT'��
���뾈�˾��N��R�������%��|F��.eɾ\R辋���  �  ��g�2���S��#|������"��G����n��N����У�
����c���:�*� ��q�=8%���B���n�z䐿�⨿$�������7B��� ���⏿Ses���L��p-�a��M6 ��ݾ��/k��a��|�����Q|�����^����aо���Z��"�7O>��a�_	��C����̰��#�����ֱ�el��5Ⴟ��U��1�����7�-��P����j������OѼ�_����a��,ݞ��6���qe��'A�T$$�������Ҿ�����_���ڐ��������珕�F⧾y�����޾%� �(�Y�-�NL��Mr�,��6��������p���Լ��[�����-�x��/L���,��E���$�
=���d��d��"���⁸�D�������1�����k����_�  >��R#�U���B��/ؾ����奄���@������S���y����ؾ+3��8�o�#���=�C�^�����R��ŕ��<���ÿ���ti��z����eo��xF�)�,�vt%��d1��AO�]L{�gJ��[g���7���lſ���|լ���������E�Z��S;�$�"��z�'�����ݾo�ž?��f��2���9	��{�����վd��5	�;$�H�2��O��pr��Y��b������Tſ{�ſ�򹿃����ͼe��A�{-���+���=�W�`�����J���������Ŀ4�ſ팺�P���s����u���Q�u�4�L��eW
�����׾u�����Z ���)��a�����ž�ݾ�������F�"��:�QzY��f�S���v��T)��*�ƿ�AÿR����H���WdX�[�8�!++�>�0���H�VFp�����}��,ֽ��ǿ��ÿ|@��m+��b���l5j�:|H��-�������L��Ѿ�Y��6���*���5��ǻ���ϾB���T��K��  �  �.�\0>��O�תb�)�x�j���ꍿw�������V�v�G2U���2�GI�A�X����+�M��d:��J]��~��Њ�n�������脿�Rt���^�o�K���;�}#,�l����
�0p��eҾ�9��tD��?���kH��D[ƾ�㾡���� g%�E5�~�D�e}V�~k�a����7��G���81��]Q���1m�YfJ�ZK)�7�����T� �5{�:�%�0SF��5i�NÃ��^�����&ъ��j����l���W���E�E6��r&����$s�ҝ澔�Ⱦr�9]��D^��bǸ���Ѿ��Y�
�[��Q-��=��mM��`�Gzu�����?��d���4���+���{�e���B���#� �������۰�"�5���W��Zz����V���-������i��h�l���X���G�j`8���(����7`�����"о�὾F\���v���yϾ뾡R�R*�;s)���9�)I��Z��m�����)0��H\��)p��9�����0�`�MY>�%�!�-����
��j�rw(��G��5j�͕����nb��Oޓ��������l�i�Y�N}I��4:�$N*�ZT��'����1oؾ�ʾu�Ǿ�ҾLp�r�����1|%��86���E�-�U�/3g���{�g͈��s��!̗�~W��n��[}�e�Z�D]9�������������H�5��bV��Ny��Ջ��x����W���A����A}��wh�ʅV���F�7���&������v]�	DӾ�8Ⱦ�ɾ�o׾ѷﾾ��3!��*���:�*eJ�i�Z�r;m��H���+��YȔ�� ��P3������Ar��PO��60��2�av��I�q0%���@��b�ȕ��GB��i����V������ʋ���*w��Pc�,BR��B���2�"��l��h�������оe�ɾ��Ͼ�@�g������n �(�1��  �  vY��X_���`�`��#`���`�Z[_�J4Y�0L���8��f!��"
�����ԾW�;8پ@q��DQ�6'��=� P�|�[��`�-8a���`��`�Za��t_�C<X��J�Y�5����5���3�Ӿ:�Ͼ	�ݾ����!��H�+���A��S��c]�h\a���a��0a��a�&�a��_�ٹV�WG��(2��`�8���5徕�Ѿ��о�⾿�����kQ/�K�D���T�j^�La��`�!�`�O�`��`�9R]���S�>TC�P�-�$��� ��4�"bо�Ӿ1�羏�"��15�s�J�g�Y�0$b���d��d��Ud���d��|d�N`�Q�U��UD��.�-����1�徖پV�޾�%��R��e%��/=�P�Q��_���f��ah�ch��g��bh��g�vb�߱V� AD��z-�������-߾J��7����6�,��D�كW��Vd�ZMj���k�k��k�M�k��?j�U"d�-4W�7�C��,�7��(y�����徺��B��C4�BK���]�Q7i�
6n�y�n�e~n���n��%o��[m�dSf�dX�JZD��!-�ޜ�*�����&��������}$��_<�7�R���c��7n��$r�\r���q�r�Q,r��xo��g���W��RB�h}*�����������������'��k?�U��-e�AKn�kq�.aq�q�vkq��_q���m�m~d��T��'>�8Y&���Uc ����V��qk�H%�M�+�e�C��tX��{g��~o�y�q���q��oq�q�q�ѕq��\m�2�b�n-Q��:��#�������A�����=���K�a0�x�G�w\���i���p��r��Er��/r��r���q�S�l�R�`��lN�.�7�������#�����y,����	�F��P%5��fL�C�_��  �  ?������o)��WJw���a�-N�i~=��.�����Y����־6x�����Υ�������kZݾ�!��Y7��&"�f�1�M�A���R���f�T�|�(����Ǝ�����\r���O��1.���r�������t
�j"!�Z�@���c�d���Ij��O� B��)v�� q���[�^�I�te9�g�)����j�BN��ξ1M��+0���m��)��-�ʾ1龙��{K�-�'��37��G�VY���m��쁿����t���Ō�Â��f��C���#��V �Z ��A�k�+�:�M�k�p����ɳ���ِ� ?��@v��e�l�֙X��G��|7���'��K����,꾗�;玹�5��e���@ž�߾�3 ���:}#�=�3��bC���S��g�F�|����j���z3�����`���i+c���@�p�"�������p���� ��0>���`�]d���C���f��������� ��.xl�Y�GcH���8��)�M�^��S�쾄�Ҿ1v¾����Kƾ�'ھ4��!�������/���?��MO�P�`�.�t�[��1����╿�ԕ��O��푀�E*_��=���"���MX�G���1�xQ���t�����ڔ��]��ا��`Ӌ�;���E|l�e�Y�/�I��1:��)�E?�����5d־�>ɾ�xȾP*Ծ*��۩�����s'���7�}G�SoW��i�<z~�98���h��pΗ�)#��!���tw�{~T�R4�~������P� �h;��f\�g�������������ؑ�����	z��e�<T���D�%�4��,$�q��ٜ��'���Ѿ��Ⱦ�Y̾�ܾ�����!�b���.�(>�<�M��4^�"Qq��|��G3��#��U]���,��w���-m�,pJ���,��i���������)���F�J�i�z���\���  �  �^��w츿b����R����y��Q�wt1�c���������Kþ�ǩ��X��s_�������z��^��ei��:Aʾ��mn�bb�[�8�4�Z����9���`��������Y��o���I��0
����\���5����]��w�)�A�I���w�r������r���g���z3��p����Q��o�l��lG��I)�C������پ���?T�����#̉��>�����ˡ�S���,վ�E��{�n�%�*C���g��q��\������h��� ���W���ؗ��n|���M��+�$-������2���X��τ�D���"ȳ��?�����R��?��
]��&�b�H�?���#����}��E?־$X���'�������!���,���ߠ��-��	�;\H�������J�5�ݷU���|��������������h¿��������c���t�W"I��,��"��*���E�I�o��R�����#y����ÿ�`���x���̘�rY��b�\��Y<���"���q����پw�������S8��mK���L�������:ɾ.�侗[�����+�ZTF�׎h�X����$���P�¿=lſڬ������,���ǋl���E�Q/��B+�Q:�1�Z��9��b板���9
Ŀ?�ƿ-���?��s����y}��W�ۭ9�0�!�m��qp���Kܾa{ľP7��n۩��J��U���=���w�ؾZT��L���d)6���S�g3x�`����H��tq��q
ƿ�Ŀ����;��ꕆ�T�^�O{<�S�+���-��B�/$h�U��/ϥ��պ�!ƿj�Ŀ6췿!���~錿��o���L��1����M�� ��qԾ�Ҿ�U5���ܩ�Kj��o���#oʾSz�P� �"W�N�&�l6@�j�_�%����ܙ��᯿������ǿ:���&����`��.�}���R�~6��y+��4��N���x������O�������  �  ����A���ԿhK�������d�1`4������}f���������by���f���a�( j�����_��'����ʾ�%��=��f�>���q�����5u���ۿ���ϣ��*3鿫�̿�Č���Z��B;���5�z{I�~Au�����R���N4޿ �G��'W��ʿk+��C���AXT�`(������ܾ�K��F���mH��u�ݳf��e�${r�u'��^����J��t�׾�y��i#��?N��͂��죿S�ƿ�L��
���������6��&m��%�z��L�g6�*59�~�U�[r���.��^ʿ��Nf��H����{࿵���'���|�{eG�[(�fQ��־+���ꜾTQ��!Q����w�K�|�����#_���ǭ���˾�)�;���k7�f�����Q���EտPm�|���b9�Eۿ�g��%%���\q���J�w�<��CH�b�l������"����ؿ�t�	�����8ڿ�ø��4����o�!F?�������~�׾�����}��:��gK��	8��J򍾸V���D���ľe��"�B6%��RL�%��i���Q¿���[������-y�VvԿ�W���z���Pj�K�K��7F��GZ�|��kk���/ƿ��qt��Y���F���%ӿ���܎���d��y8�K�8n����ؾ�⼾Rp��P����i�������L���>���ʹ���Ծo�������3���^�/���1��.ϿԤ쿶j���>��p3�F�ɿ"ե�����UN]��F�`�I���e��F���ɭ�jѿ����F���H��/��ǿA���k���C�T�R>,�yV�MU��	Ͼ���^ ��5���沓�����zU���˃þ���I�αA�v�p�i#��]u���mڿ����}����S��,P࿶_���
��M{�nPT��F��Q�V�u�9z�������ݿ/����  �  �������g ��jԿ�����+}��q>�TA�P�޾�԰��̐��u��X���H���D���K�4�^�?�~�8����b��~T쾂��xoK�����ΰ�!߿���Hc����/3�k���olʿӞ���z��T���L�X�e�cg��sN��KB�-�_}�������
d�HsſQ���?lg�&r.�����Ͼ+˦��[��9	n���U��_I��H�QUS��j�g��ӏ��îɾ�� ��(�4�_�i��E���
���������;��Cֺ��葿�i��M�QZQ���t�N�����ſ�������C#�����(���,��H�U��O"�����RǾ0x��[ӊ��u�Yb���Z��J_��7o��Ӆ�F}��@ͺ�cv�΄�4@�r}�����p*ӿ �$k����h%������ݿ�f���Ice�%�S�6!b��Ї�4/���1ٿ���v������M"�p�ٿ_������WI�1�����Ǿ"d��1Ǒ��⃾��x���u�ݫ}��Έ��V��^뱾\.վϷ�Jf'�q&Y���m���g�忼b�����a���q����4ҿҦ��v����d���]���v�ߖ��ɾ�޽��R���t����������Ϳ�>����w�s�>�>_�!�m#Ǿ ���-��e抾d����]��k����%��X���{�¾�꾂���8��p�DP���3ȿ�i��������VK�q��N�`Eÿ~S��v}z�/9^�M�a�S���	����tͿR��[��Y��%��!�Z���1��F�����b��d/�P}
��#ᾩ�������?���>���-���Ԇ�G��!���I1���оei������xJ�1����ͪ��Lؿ'������f�����2�4���G��i�����n��2]�Luk��i��	���;�ݿ��w���  �  �8+�D$�������f�������;H��/�IDܾ=Ʃ��ᇾ�0c�^_G�wf8�Zn4�`;���L��Vl�W؎�����E�[��A/W�k���x�ÿ� ��G2��'��+��!�ӽ�T��������?e�!�\��ly�����ʿ`; �����Z(�}�*�)�R��Z�ۿs���w���5��U�V=˾ើ�7����[��fD�L�8��H8�S?B���W�6o|��j���ľ���D/��n��š�eտr��"���)��)������2п옠��~���]��b��\������=�ܿ�I	�â�S+��)��n�I� ��L˿�T����b�\3'������k��������5c�6Q���J���N�_�]��Uy��~��+q��*B侬��^I��臿Ե��h�7���$��(-��'���,���`ÿ◿��w�Y�c��t�x3���[������s�9�&���-��&�+���	�q	��1���!S�Z ��M�g���z������;v��:h��He���l�y���"���C����ξ1���+�g�d��]��^iʿ�} ������*��.���$�����'�ߘ���� �u���m�,�����[ӿ�y������,���.��\#�+&��)�l��������E�0����뾦9��-u�����0M��+y�dx��/�����d^�������f��hO?�4�� ���ݿ�
�Y!��.��L-����H.���ؿ�	���q��Eun���r����+���a�俦�9#���.�m`,�F��<� �ѿ|�����o�7G4��^
��;۾ u�����LK���π�fz��%}�1����ђ��.��9�Ⱦ�2���6 �WS�1���񺿝��G��v'�ʸ/�W4*�O�+��3?ȿ�������Zm�j}�Ҙ��¿W;����Z�(��  �  }?��<yu��eW�.�)��:�������S<�(���;���f���fh�Z2V��bQ��VY�ro�;��^Z��t۾���CpK�@����u˿�~�.�7���_���y�,���np���N�û$��2��*W��鉗��;��xd���ٿ����<��\c��{�͏�>�m�!�J�����=�l0��im�o�)������������Z���c�h*V�yVU�da��|�3Ҕ�w ������Y#�P�c�i{��o�@����E��'j�X~��}���f��"A�MM��f�����ؑ����ܴ��!� ���J���m����Ԅ|�z-d���=����տNB����V���:��U��*떾�ꂾԬo��g�!Yl��Q~������_����վ��t=�z��h���� �/)+�*U���t�M1����y��|]��5�|�
��п����.5��s䠿�
ʿ�����0���Y��x�r���/x� Z�1�0���-���_$���@G�-������-���e���������.��"���a�����N�ľu����y ��*Y�����7Zҿ���\Z;��
c��{}�d���$t�9�R�Q�(�: �+�¿]��qә����U�;?��A�3�g�m��8���q���N�{�#�L����x����}��':����+߾S踾i����0��A���ӊ�!ݐ�u8������Yپ9��ƥ3��Xt�ʵ������`J��[n��H������H�j�ofE�ɒ���迈���]Z��r���0��>I���	$�3�N���q��́�����}g���@�[d���ۿٝ��&d�i)����=�о&���������M`��&ԕ��'�����8*����YG�����! ����	�-��W�{�w�yy��U|���_��7�?���Կf���Z옿K���:�ο	����2�;�[��*z��  �  Hhu�o�j��2N�s�&�qb��gi�����:�5��3�Ͼˤ�ވ��/o�~�\�C�W�0�_���u�%w��l����ܾPl��H��>����Ŀ���H0��V��/o�i u�$f��JF�e��}^��{N���O��+`���%ҿ�E���4�r�Y�_q���t�
Uc��"B�j_���㿶u��:�h�%l(�ho���Z���盾�Ѓ���j���\��[��h��y��#6��\ǻ���[A"�	�_�C��3�ۿ����=�~`�pWs��/r���\�]9�g�(zؿy西|㍿����u-��Hr翢���[B���c�u�m�q�skZ�Ͱ5��z�y
οu}���S�mJ�H��iQ���[���Z���Ev�+n��r�����Zu�����D@ؾ���E;��ɀ�Џ�������D$��*L�uj�lKw��$o�3/T�R�-�$���=ɿ*S���V��h���~ÿǧ�-r)���P�a�m��x�b�m��P�I�)��� ��ۻ��4���E������dd��(ޟ����O��9b������*���5�����Ǿ���J ��KV�"��׼˿p�
�A�3�uY�Ҭr���x�Y�i�2%J��"��N���ż�<қ��㕿������ڿr��/59���]�?Gu�T�x���g�'YF���l7�*���py�~�8����G�ᾃC��;��6���}{��F��M1��p���Zy��� ܾI	��2�FTp��P�����A����A�jEd�A�w��lv�Pa�l_=����/�%o���`��}d��j{���￢���%F�Ojg��x��u� �]�r�8����A�Կ����`�ra(�$����Ӿ"������jg��/��������4�����CTľ�����rE��셿^�������c�&�7�N��	m���y�N�q���V�[+0����οJ��*��T���"ȿ��� �+�:�R�֟o��  �  �&W���M�{S5����/�⿅M����t�Ƌ5�V�	�e�ؾt꯾�S���x��R(q���k�֗t�� ��:���<����;���/B��{��B������m��~<�`�Q�L�V�$J�ߝ.�j!��;ֿ����ɑ���e��w����������.��WU?��mS�=hV��G�H
+��R�s�Ϳ�M��?H^��/&�i����,˾�N���"��{����p�i�o��*}�����s���q�žs����� ��pV��֑�8�ƿ};��'���D�OZU�shT�2B�)C#��\ ���¿���6₿֐��q���H�Ͽk��N+�hH��W�I T���?�=� ����룻�)���!eL�k������ľbݥ�cy������U�������N���۞��ٹ�CV�a�=X7��[t�[x���1߿����3���M��
Y��R���:�G�����l���x��[���+���㒱��0�,���7�2�P��Y��P��8�Ά�#���������>z@�
��k��#�ƾ�S���왾���]���J��P���� ����Ҿ�v���N ���O��^���w�����|8�+�?�U@U�"�Z��M��q2����f޿�T��z�������ƿp'���#��C���W��Z� �K��@/�����5ֿN���E�n�\�6������0�Ǿ�g���+��$����������$מּ(�þ?�+7�1���f�����Ͽd�N+���H���Y���X��BF���'���aa˿
��JT��f�ϧ���׿.S�/�P�K�)�Z��]W��GC��#��� �48¿����)�Y��(��R��޾<��3=���Н�IØ�˚�� ����a�Ͼp�����q�A��~�U����T促f�}r6��P�}�[���T�T=�[:�}��[6���6��vF��%����/��˹�9c��:���R��  �  ��-�պ&����W���M���蔿0�e�a)4�w���w�Ǿ���\������^ڇ�,��[��������9Ͼ\\�����xJ>���s��8���̿�� �8��)� �-�N�#�7�+�,�������m��`e�����X꠿G�Ͽڪ�~3���*�>-���!�p,�:�]������jT�W	(�f�&T�4d��ʤ�z���,���S	��D����)�������Wܾ�����#�2N�K���#���M�ݿ�(	���(b,���+��;�vb��Կ���vJ��Xf�Vmj�6���V1��i��8��z'"���-�^�+��C�Jj�3Կ����j]~�� G��~����E�۾���|r������~���T�M���崾��оd������7�\�f�y���˿����A�$'�ƣ/�D&*���+����ǿ]E���2���l���|�����3�¿.�������J)��l0��v)�ʦ�ŕ����ƿ"]��ǖp�?�T�������ݾf����-��?��pI��l���5����ʾذ�0�	�ߐ%�KL���� ���ӿ��k���&-��(1�#0'�����q$���O��'Q~��Tv�=���8z���ؿ����z�3/��~1��&�3c��e쿣V���?����d��k8�,d�� ��޾ež�³������0��*"��o\¾f�ھ����q��y�3�`�^����*۴���`V���#���0���/�-y!�A�	�gRݿ�{��Һ����v�Z�z�\ё�&���<�:|��%�H1���.�f�������ڿ�M��JŅ�MIT�ѕ,�m���i���վ�3��dа�T����-�����
 ˾��S��}vA�Fq������ĿpD�������)��92�C�,����� ���̿y����P~u� 򂿧.���vǿ������\+��  �  �$�T����A��zĿ(=��N����r`�U�=�ϣ"�s������Ͼ[��XЧ��w���s�������־1D�������(�/fE���i��͌����	q̿ ��� �M�<m���]ٿ볿_Ph��G�D�A���V�P��wZ���/ɿЭ�g� �U�����sۿ����¡���(~��U��D5��������8aȾ�u������r륾3q���1že�⾣l�����1�]�P�kx����6����f׿����t��u��k�<�̿��)����Y�_IB���E��gc�â��e@��`=ֿr���aa�WM�[����ѿ������Ur���L��t/�Bx�A
�'��"cȾ1<������[�������پ�������0'��B��c�ɻ��թ���Ŀ������n!�� �O�ndĿ��P����W���H�0U�+{�
ϛ����!��m� ����m��3��V�ɿ(���4���Yk���H�	�-�b����������ξ����ܻ�jXþ�վ����	�^��D6��S��w���������FOӿ���G�<��������࿄���(痿�ex��PX��R��g��Ԋ�_嫿��ѿu9��"B��P�L �g��\¿���>]��ۄe�&�E��+��)����פ�g�Ҿ��ƾ�ƾ6�о\c�e�ŗ�?�(��B���`��n��=K���⽿��߿����������m���zWտ\t��
���S�j���R���U��ys�Pz��&ܷ���ݿ������ݦ��u����ؿ�����8��׃���Y���<�^n$���B�����.ξyiƾI�ɾR�׾���f���6���1�y~L��n�aߌ�[Ш���ɿ���Fc�X��ބ�6`�*`ɿk��儿�#a��7R�=^�����?���Fſ��鿀���  �  ���R��v���GԠ��� k��N�p��\\��G��H1��2�'��澃�оiFʾ�VԾp��c	������6���L��Oa�m�u���������\िF��8H��"���CԳ��ǟ��-��5�^�A9���"�ѭ��-�gL���x�^/��=��V��k����ܹ��F��$�����������j��V��`A�D�*���_D���;߾E-ξ�3;�jܾ��������'� �>���S�
h���|��Ԋ��ș���T2��V����w����{��t+}�/P��G/���?q!�6�r�Z�[�����*��j��6p���o��Nu��(0��z�����{�7Hg�iS�"[=��y&�JR��������:�վҟھG�ﾊ��L_�δ5��}L�іa���u�����2��~墿V���V��{Jÿ�1���ܪ�[C��Fhu��K��?0�{&��.��H�^�q��X������d����Ŀv����>���T���m���߈�2k{�JKg�\�R�	o<���%�*������y辒�⾏%�p�pI�{�,��D��`Z�8o�;��f��ȍ��=���*���;ſ�ſ���9���֎��en��I�M73� R/�k�=�4V]�Ǆ�����_x����ÿUzȿ�S¿����~W��0��zT��YF{��g�߭Q�A�:�Z�#��C��n��hV�LY������L!�S�7�L�N��:d�Pfx�W���?�����Hq��|����ǿ0aĿ����蟿(�����`�.�?�*�/�R�1���E��j�����\��W3���?ƿw ǿ�	����*��U��}���ot�3 `��KJ��=3�n��d�	�(��NP�2��1�	�R)��n@�?W���k�l��2���Y������2���Ŀ�|ȿ1Y���󯿊E���@�g�U�7�9�Ow/�`�7���Q�nPz����u���r���  �  mߌ�N�� l������D���Q����P������6���m�h�M���-����K����t�����4�A+U��lt������"��ܐ�����+�,�����{\�� �x���i���H�k�)�4�8I�����!	������:��.[�ʲy������&��7����!��Y����>���"���犿����X,d���C��F%�������[ ����"��?��Y`��}�^ʉ�l��������G������A��А��"�������{�q�]��=�r& �]�
���������i�A�'��F���g��V��U����������X�������]��SĒ�C���ϭ���{��+]�B�<�>� �!��	3��������1�U�P�mq��b��뱏�^퓿{r������-��2?���_��w������^z��![��7;�) ���)=�����m�u=9��YY�,dy�T承8W���ϕ���&���,��>���*Õ�$������'�x�i�X�}9�V���9�J�
��o�+�%��A��;b�7݀�1b��R���(���[����Ӗ����ߗ��O��I ��!���N�w�e�W�#P9�*� �����o���.�a�K��*l��Z��+��΢�� ����-��0����ژ�����^��/�������ft�S�S�Pg5��
��(�4n�$���32���O��p���-����*-������	������.��ц��x��NV��7�n�==N�ܿ0����$��������6�@�U�av�S��od��C]��(R��$���MD��j󘿨Z������3���N����i��I�"-�d��������"�VC<�3�[�D�{�����政���閙�kϘ�L����r����������:莿�I���/e��E���)��f�����-['���A�N�a��Հ�)��  �  �8]�:~q�����Ñ��á�U���ּ����Q���=����� oe�6�=���$��n�	�(���E��o���?��E1�� ���eD��f����s���ݎ��Ɓ�h�m�<�Y�ƹD��.�a���[0㾖�Ͼ~̾��ؾ�F��y���$�1;�2�P�[-e�R�y�h숿����ӧ�h����J���ͽ�X/��'����#���W��M4�F� �����61���R��H��H,��Z ������k��&���]K���瘿����x{�ԍf��WR��<�G�%�M�^@��g�ھ�̾�CϾj�ᾬ&�7D�f�-�2�D�ZZ�Żn�3,�����:k��d���f�������u��@���^�����y���N�Qi0�,=#��(��@���f�h���(��)񷿰K¿�d�����i|��DZ��!Y��l�{��jg���R�(=�S&��>��\��q�<�۾$�������s��r%�M�<��XS�z-h��|�ُ���C���<���
��<H¿�Ŀ!���lר�S���U q��jI�Ғ0�L�)��5��R��|��9��Zڮ��迿�ƿC ¿���U��[���f�����{���g�rS���<��"&�,v�Y�|�ﾩ��z�����
�/W���4�L���a�[v��`���V���៿�'����ǿ��ſ�T������9�� �g��eD��1�y�/�BIA�qc��W��H@�����Ŀ�ǿ�쿿���z2��UW��&��IMw��c�J�M�В6������X��$����_ �k:�~�$���;�h�R���g�}|��ƈ���������\J����¿�5ȿ�¿Q��~���6���Z�\~<�Z%/�,^4�y�K�Hr�*������@��[�ǿ�ƿ[(�����ކ������>����q�~U]��:G��!0�%�O���v���p�����X�;��-��E�pg[��  �  �i?�]ub�t	�������eƿ������+�#���y�޿��=,���:o���J��8@�ƲP���z����͓¿�E��'��0D�����࿆&��@n���܂���Z��9��D�5		����8z̾������t��=�F4��^`ݾeb ��4�	�-��bK��q�B����e���Jҿo����_���w�I�ӿ��������a���D��nC���\�
2���s���PϿ{Q���Y��_�#�տ����a��F�u�mUN�5�/��������߾xJþ�h����`֧���9̾Q�����]7�n9���Y��ၿfӜ�u)����޿�p���	��x����fɿ�m����fY�	.F���M�Q�o�����V�]޿������� �O�dο�n��qݎ�v�n���J��.�:F��W�Q=��e˾Nݺ�E�������˾z���J��K�S�.��aJ��|m�Ӎ���y����˿�j쿾���K& ��j�ƨ������� {�ϘV�WGL���\�둃�S��<�ȿ���������� �`�\ƿ�O��!É���h���G�:�-���s���	�b\Ծ�tǾ�ža�ξ�p�1���=��&�<�>��M\��;�����'ĸ�e�ڿ&�����a���k�ۿ�ε������3q��	U��S���l�=��+���d׿nk�����n�����c�ݿh��K���O/��4_���@��'����� �k侽�Ͼ��ž�Ǿ�Ӿ��龑_��#��-�:�F��4g�9{���d��,�ÿ~a��~ �SL�5��Q=�jXϿ����/��@se�2R�	�Y��u{��7���d��� ��v�n��2�G:ӿC�������>y��@U�K�8��!�@n����,�޾P�;`�Ǿ��̾r�ܾ.������}�,�6��  �  @?6���h�����Ŀ��5�^�'�j�-�J�%�R&��ￆ����#����q��c�Bz�R%����ƿA
���l�6�(�S�-��{$��%���쿧���~ݎ�C�\�u.��g��羃þ������(A��h���������>���n־� �����F��~�Y����տJ�*���c+�#�,�ó ��
�g7޿q���s1��$�i���g�	��ŧ��0ؿX���:&,��#,���������ڿ���佂�z!K��(!�7���xپ̀�������Z��A\��:�����u���Kþz�羡����,��-Z��w��5"����迾[���#�DW.�p5+�[���0�g�οy���|
���i�t�Od���Z�������&�5k/��*����.� ��wͿ!x���Ww��	C���3g��ܾ4$���I�����܂��j֝�����{���ݾ?J����9A�%�s�ƒ��d�ɿ������U=*���0�S�(�2��͋���n����¾}���o�����F��q�̿50�¨��@,�U1���'�q���v�ry����b�j�#<�L��{[�$��kƾu����檾����t��������׾��������.�VmW�Eه�L���O�ݿ;@	�� ���/�K1���$�z�)L�ᵴ�=����y�Y�w��'���ϯ��>�����"��60��80���"����1��^�������[���1�5������{bپ�G��g~��	���1����l��lƾ�8�������B:�q~g���������5����&�"�1�ri.��!�M���Կ�����×u�����:�������������(��2�[-�^1�%~���ҿ����6ဿpM�!�'���������Ҿ�������N���꯾(���о���Tv
��$��  �  8;8�i y�t+���%�|���7�� O�Z1W��1M���3�W��D࿑���F`���R�������޴��^�и�q�:��Q�jW�� K��Q0�<��ؿ&,��dli�b�-�2��[ҾG૾j��~���3�q�t�n���y�Arg��ꩿ�����e�L�Ἂ��D���I��ܬ!�V�@���S�<V�gF��1)��_�5�̿꽝�(%���Ճ��ә�SXƿ}��_%���C�
U���T�-mC�6O%�%Q��hÿ&=���R������þ����_���Jr|���p���s������ؒ��N����Ѿ����i+���d�mu����ҿ��Ů-���I�\�W�r�S���>� ���1��I�bF��!{����-ɨ��;ܿ{�1�1���L���X��R��6<����vs����΄�~GF�������_�žƘ����������>����G��5��o&��%�ž�ﾐ��#7C������p�����9��Q��Y��O��6�r���������V���P��%���[�Ԇ������=��LT�dZ�`N�L�3�����޿P���Lw���;�� ����|ɾ�P��)��Tl�� u��=���^ા���O+��>�E�*�c]�F)��G�ſ���e�%���D�RX�4Z��xJ�T?-�3j
�i�ԿUɥ�8.���݋��ܡ��bο���h)�E�G�*,Y�yY���G��m)�t�Z�˿����	Ic�|�.�Ȕ
�侢m¾�����5���Ø�����M[��ɾ�������8�Z3r�b
��1mٿYW��0���L���Z�b�V���A�P�!��G����¿gC��p��;���4��R���4�zO�Dp[��BU���>�T.�W���xC�����]�P�,>"����$�پKm������������S���ǧ��C����־2 �=���  �  ==��$���͹�9X �d;)�E.P�5l��pu�O�i�8FL���$�����g$���������r���)ȿ�����-� T��@n��Iu�_^g�dSH�8- �b��¬��u�\"1�g����Ⱦ����8����m�#�]���Z�@
e�]�}��蓾F)�����̋��eT�:���G@п����+7��h[�c�q�`!t�f�a�F�?�}c�D��B��~|��t���$����}ܿ���a�;�ԭ^���r��r� �^�u;��R�9�׿4��&�[�/�����ϸ�!D���h���g��]��_���o�ڕ�����-Ⱦ���r.� 4p�/�����'}��E�^�e���u�&q���X���3�}7�:#ѿ�ڢ��W��S䖿o�������!�"�I��i�w�v���o�0�U�P�/�ƪ�7�Ŀ�/��z1L��^��辶Һ����⯊�����*6{�����N��6���[亾
y�R{��9H�詉�2T������+���R�!�n��1x���l��O���'��A ��¿�������o���")ο��i1�^KW��}q�^�x���j�
�K�%�#�`���f���F쁿�(?��&�U��W$���פ�٧���/���Y��0������L��Z�־D���e+�>Be�b���ؿ"��S;�ӊ_���u��7x���e��D��m�P�뿌��o���q ��������w��j�?��b�a
w�Q�v�+�b��?�]u���߿X_��k>l���/��z���پ������������卾a������9���������H�;�;��}}�*������GVH���h�7�x�IMt� \�_�6�	>�$׿�Ԩ��L���Ӝ��i��ko��=�$�ŠL�+�k�(�y���r�O|X��V2�1B	�X�ɿ�d����V�y�!��/��� Ͼ����񧓾�������ܜ�Jʮ�R�˾9����|��  �  Z�?��5���п�SZ��~0��zY���v�SC��$Lt�xFU���+��2�ϋ¿#	������\g���(Ͽ�
�o5�y�]�F�x�,/��%�q�77Q���&�>������{�f�2�%���Cƾ�K���2����f�VW��YT��m^� �v�U{���9���}��J��W�����~׿���V)?�(Ae���|�/ ��k�qVH�K��PT쿒���쑔����^ݭ�������r�C�ܘh�]�}���}���h���C�WT��C߿�J��Tj_��* �-�� ��㒾*�y�sa���V��`Y��:i�.%������[xžo3�?�/���t�������� #���M�"�o�m��9�{�u�b�%k;����U�ؿǧ�?���-������p���y�(�%�R�(cs����G�z�Fc_��C7�����/˿����2�N�������ݷ��?���5F���z���t�X�{��釾<��a����[� ����J���� Wſ��A=3��6\��ky�����w� X���.��#�#{ȿo�������(f��y0տ�	�|�8�+�`�/|��ԁ��&u���T��W*�E����帿�|����@����:�"պ�xY���B��Wꊾt��£���-�������Ӿ��e#,�9�h��	���߿>���QC�Bci�B`��J���
p��cL�b�!�Nc��в��Қ�����嵿$�쿟��l�G�٤l�����������l���G��v����)���Fp�Y�0����|�־�����J��|^�������l��X�������1g����ᾒ��`�<�C���������?&��Q��(s����[���e��x>����؆޿�����3�������ſLb�2_+�7lU��v�A[��Q}���a�[�9�<���bп�����HY��"��B����˾:y��l���a��茾�Ϗ��u���R��{bȾ�������  �  ==��$���͹�9X �d;)�E.P�5l��pu�O�i�8FL���$�����g$���������r���)ȿ�����-� T��@n��Iu�_^g�dSH�8- �b��¬��u�\"1�g����Ⱦ����8����m�#�]���Z�@
e�]�}��蓾F)�����̋��eT�:���G@п����+7��h[�c�q�`!t�f�a�F�?�}c�D��C��|��t���%����}ܿ���b�;�֭^���r��r��^�u;��R�?�׿9��-�[�"/�����ϸ��C��vh��@�g��]���_���o�������[	Ⱦ���/.��2p�b��̇鿱|�E��e�v�u��%q��X�\�3�L7��"ѿ�ڢ��W��g䖿����j���L�!�o�I� 	i���v�'�o���U���/�;���Ŀ�0���2L��_����>Ժ�����������:6{����DN������⺾%w�*z�I8H�!���US���+�+�|�R���n�r1x�9�l��O�b�'�pA �k¿�����������c)ο3���1��KW�P~q�חx�+�j���K���#�S���G���큿*?�)(�g��&��٤������0��ZZ������䥟������־W���e+�FBe�d���ؿ"��S;�ӊ_���u��7x���e��D��m�P�뿌��o���q ��������w��j�?��b�a
w�Q�v�+�b��?�]u���߿X_��k>l���/��z���پ������������卾a������9���������H�;�;��}}�*������GVH���h�7�x�IMt� \�_�6�	>�$׿�Ԩ��L���Ӝ��i��ko��=�$�ŠL�+�k�(�y���r�O|X��V2�1B	�X�ɿ�d����V�y�!��/��� Ͼ����񧓾�������ܜ�Jʮ�R�˾9����|��  �  8;8�i y�t+���%�|���7�� O�Z1W��1M���3�W��D࿑���F`���R�������޴��^�и�q�:��Q�jW�� K��Q0�<��ؿ&,��dli�b�-�2��[ҾG૾j��~���3�q�t�n���y�Arg��ꩿ�����e�L�Ἂ��D���I��ܬ!�V�@���S�<V�gF��1)��_�6�̿뽝�)%���Ճ��ә�UXƿ}��_%� �C�U���T�2mC�<O%�+Q��hÿ0=����R�!�����þ���������p|���p���s�%���t֒�	L���Ѿ���[g+�(�d��s����ҿ��߭-��I���W���S���>�����0����F��{��5���ɨ�|<ܿt{���1�n�L���X���R��7<�l��6u�Y��YЄ�JF�������Z�ž ��� �������M����F���3��O$��?�žR��R���4C����v������~���9���Q�?�Y�W�O�V�6����?��O����U���P��c����󺿐�������=��MT��dZ�aN�D�3������޿���Ow�k�;�9#��	�-�ɾpS��Z���n��Vv��A���!᪾�����+�?�]�*�c]�J)��I�ſ���e�%���D�RX�4Z��xJ�T?-�3j
�i�ԿUɥ�8.���݋��ܡ��bο���h)�E�G�*,Y�yY���G��m)�t�Z�˿����	Ic�|�.�Ȕ
�侢m¾�����5���Ø�����M[��ɾ�������8�Z3r�b
��1mٿYW��0���L���Z�b�V���A�P�!��G����¿gC��p��;���4��R���4�zO�Dp[��BU���>�T.�W���xC�����]�P�,>"����$�پKm������������S���ǧ��C����־2 �=���  �  @?6���h�����Ŀ��5�^�'�j�-�J�%�R&��ￆ����#����q��c�Bz�R%����ƿA
���l�6�(�S�-��{$��%���쿧���~ݎ�C�\�u.��g��羃þ������(A��h���������>���n־� �����F��~�Y����տJ�*���c+�#�,�ó ��
�g7޿r���t1��&�i���g���"ŧ��0ؿ[���?&,��#,���������ڿ���򽂿�!K��(!�0��bxپa���ܸ���Y���Z��CK
���r���Gþr�羢��5�,��)Z�qu����� �迃Z�z�#�'V.�s4+����0�k�ο����
���i��t��d��}[��J�쿥��&�Il/�O�*�̞�o� �AzͿmz��/\w�XC�:���i�c�ܾd'���K��4���򂙾{՝�艪�
x��[�ܾ�G�����5A���s�p����ɿ ������<*���0�T�(�_�������m��x
��/�}���o�	���G��q�̿�0�����A,��1���'�ő�<y��{��ŕ���j��&<����Y^�����nƾ����K骾����㽰�����׾h��ʩ��.�jmW�Jه�O���P�ݿ:@	�� ���/�K1���$�z�)L�ᵴ�=����y�Y�w��'���ϯ��>�����"��60��80���"����1��^�������[���1�5������{bپ�G��g~��	���1����l��lƾ�8�������B:�q~g���������5����&�"�1�ri.��!�M���Կ�����×u�����:�������������(��2�[-�^1�%~���ҿ����6ဿpM�!�'���������Ҿ�������N���꯾(���о���Tv
��$��  �  �i?�]ub�t	�������eƿ������+�#���y�޿��=,���:o���J��8@�ƲP���z����͓¿�E��'��0D�����࿆&��@n���܂���Z��9��D�5		����8z̾������t��=�F4��^`ݾeb ��4�	�-��bK��q�C����e���Jҿo����_���w�J�ӿ��������a���D��nC���\�2���s���PϿ�Q���Y��_�6�տ����%a��i�u��UN�A�/��������߾�Iþ�g����ӧ��%̾6�뾣���3��i9��Y�߁��М��&����޿�m�����w�����ɿll���񂿡eY��-F�*�M���o������︿�_޿������y!�B�eο�q��@�����n�h�J��.��I��Z�JA徦h˾�޺�a��x���˾���<H��H�Y�.�$]J�Rwm������v����˿�g�I����#% ��h�C���{�����z�!�V�cGL���\������T����ȿ����V��M� �0c翆	ƿ�R��Ɖ�W�h���G�k�-�w��j��s�:`Ծ�wǾ7�ž �ξ	r� ���U=�2&�a�>��M\��;�����'ĸ�e�ڿ%�����a���k�ۿ�ε������3q��	U��S���l�=��+���d׿nk�����n�����c�ݿh��K���O/��4_���@��'����� �k侽�Ͼ��ž�Ǿ�Ӿ��龑_��#��-�:�F��4g�9{���d��,�ÿ~a��~ �SL�5��Q=�jXϿ����/��@se�2R�	�Y��u{��7���d��� ��v�n��2�G:ӿC�������>y��@U�K�8��!�@n����,�޾P�;`�Ǿ��̾r�ܾ.������}�,�6��  �  �8]�:~q�����Ñ��á�U���ּ����Q���=����� oe�6�=���$��n�	�(���E��o���?��E1�� ���eD��f����s���ݎ��Ɓ�h�m�<�Y�ƹD��.�a���[0㾖�Ͼ~̾��ؾ�F��y���$�1;�2�P�[-e�R�y�i숿����ӧ�h����J���ͽ�X/��(����#���W��M4�I� �����61���R��H��O,��c ������k��9���sK���瘿����x{��f��WR��<�'�%��L�v?���ھ�̾�@Ͼ���`$�TA�ۢ-���D�,UZ�K�n�7)�����h��7���`�������s��1�������Z�y��N�bh0��<#�y�(�-@�ճf�߄��*��w�^N¿�g���������]��E\��D�{�-pg�aS��=�]&��@�`���r�]�۾ҝ�%���`q��o%���<�TS�5(h��}|�����P@��e9��F��E¿@}Ŀ����aը�������p�kiI��0�Y�)��5�aR���|�9;��~ܮ�D뿿؍ƿ}#¿����\Y���Õ�����Ź{�2�g�9S��<�F&&��x�7[����<��h�����
��W��4�ZL�$�a�pv��`���V���៿�'����ǿ��ſ�T������9�� �g��eD��1�y�/�BIA�qc��W��H@�����Ŀ�ǿ�쿿���z2��UW��&��IMw��c�J�M�В6������X��$����_ �k:�~�$���;�h�R���g�}|��ƈ���������\J����¿�5ȿ�¿Q��~���6���Z�\~<�Z%/�,^4�y�K�Hr�*������@��[�ǿ�ƿ[(�����ކ������>����q�~U]��:G��!0�%�O���v���p�����X�;��-��E�pg[��  �  mߌ�N�� l������D���Q����P������6���m�h�M���-����K����t�����4�A+U��lt������"��ܐ�����+�,�����{\�� �x���i���H�k�)�4�8I�����!	������:��.[�ʲy������&��7����!��Y����>���"���犿����Y,d���C��F%������ \ ����"�!�?��Y`�.�}�jʉ�|��������G������A��А��"�������{�S�]���=��% ���
�����F���g�؞'�ӳF��g��T������4���l��� ��4����Z��H���}���a���̲{�d(]���<��� �0���2�p�����1�A�P�0q�.e������\𓿵u��ޫ������|B���b���y�������bz�)%[�6:;�� ����:=�7��l�&;9��VY�(`y��㉿jT���̕��앿S#��y)������	���0!��1����x�4�X��z9�͕��8�W�
�Xp�ӭ%���A�J?b�X߀��d��@���e���Џ���ז�����◿�R��1��������w��X�S9�o� �C��c�l����.��K�J+l��Z��<��ע��$����-��/����ژ�����^��/�������ft�S�S�Pg5��
��(�4n�%���32���O��p���-����*-������	������.��ц��x��NV��7�n�==N�ܿ0����$��������6�@�U�av�S��od��C]��(R��$���MD��j󘿨Z������3���N����i��I�"-�d��������"�VC<�3�[�D�{�����政���閙�kϘ�L����r����������:莿�I���/e��E���)��f�����-['���A�N�a��Հ�)��  �  ���R��v���GԠ��� k��N�p��\\��G��H1��2�'��澃�оiFʾ�VԾp��c	������6���L��Oa�m�u���������\िF��8H��"���CԳ��ǟ��-��5�^�A9���"�ѭ��-�gL���x�^/��=��V��k����ܹ��F��$�����������j��V� aA�E�*���cD���;߾L-ξ�3;�jܾ�������#�'�2�>���S�6
h���|�Պ��ș�.��j2���V�����x����{��6+}��P�,G/����o!�@6��Z����@���(���g��Tm���l��r���,��e�����{� Cg��S�MW=�}v&��O�m������݅վݠھ��ﾄ��
b�S�5�E�L�՛a���u���5���袿���Y��IMÿ4��ߪ��D���ju���K��@0��&�]�.���H��q��V��~������/�Ŀ[���f;��1Q��\j���܈�Ie{� Fg�ʥR�>k<���%��'������x辫��%'�q��K���,�zD��eZ��o�LŁ��i��;����ë�v-���>ſ�ſ"��>;���؎��hn��!I� 93�gS/�\�=��V]�ZǄ�����xx����ÿ[zȿ�S¿����|W��.��yT��XF{��g�߭Q�A�:�Z�#��C��n��hV�LY������L!�S�7�L�N��:d�Pfx�W���?�����Hq��|����ǿ0aĿ����蟿(�����`�.�?�*�/�R�1���E��j�����\��W3���?ƿw ǿ�	����*��U��}���ot�3 `��KJ��=3�n��d�	�(��NP�2��1�	�R)��n@�?W���k�l��2���Y������2���Ŀ�|ȿ1Y���󯿊E���@�g�U�7�9�Ow/�`�7���Q�nPz����u���r���  �  �$�T����A��zĿ(=��N����r`�U�=�ϣ"�s������Ͼ[��XЧ��w���s�������־1D�������(�/fE���i��͌����	q̿ ��� �M�<m���]ٿ볿_Ph��G�D�A���V�P��wZ���/ɿЭ�g� �U�����sۿ����¡���(~��U��D5��������<aȾ�u��Ĝ��z륾=q���1žw�⾯l� ����1�v�P�!kx���J����f׿����t��u��k�3�̿� ���(��@�Y��HB���E�fc����� ?���;ֿ[���+`��K������ѿ��S����Pr�^�L��p/��t�����U`Ⱦ�:��ˢ���\�����-�پ���̈��4'�"B��c����������Ŀ��Ҕ���"�G� �Q��eĿ'����u�W���H�� U��){��͛�����;��G� �������'��A�ɿ%���[��FTk�J�H��-�������zξY���5ܻ��Yþ��վ7���	��a��H6�� S���w�u�������vRӿ��sI����������*���w藿�gx�RX�B�R��g�!Պ��嫿ݼѿ�9��'B��P�L �f��Z¿���=]��ڄe�&�E��+��)����פ�g�Ҿ��ƾ�ƾ6�о\c�e�ŗ�?�(��B���`��n��=K���⽿��߿����������m���zWտ\t��
���S�j���R���U��ys�Pz��&ܷ���ݿ������ݦ��u����ؿ�����8��׃���Y���<�^n$���B�����.ξyiƾI�ɾR�׾���f���6���1�y~L��n�aߌ�[Ш���ɿ���Fc�X��ބ�6`�*`ɿk��儿�#a��7R�=^�����?���Fſ��鿀���  �  ��-�պ&����W���M���蔿0�e�a)4�w���w�Ǿ���\������^ڇ�,��[��������9Ͼ\\�����xJ>���s��8���̿�� �8��)� �-�N�#�7�+�,�������m��`e�����X꠿G�Ͽڪ�~3���*�>-���!�p,�:�]������jT�X	(�g�(T�6d��ʤ�}���1���Z	��M����)�������Wܾ�����#�2N�W���2���]�ݿ�(	���0b,��+��;�sb�
�Կ���;J���f�[lj�����o0��<��{���&"���-�9�+��B�i��0Կr���@Y~�G��{�>����۾����=p��{���=���𕾷O���贾��оX������_7�k�f��{��Tο�&�C�] '��/�B'*�c�z����ǿ F��3���l��|�j���H�¿�������I)�dk0��u)����2����ƿ�Z����p�S?������w�ݾM����+��G���I������7��їʾC����	�;�%�4L�M���m����ӿ�����(-�*1�*1'���I�%��cP��iR~��Uv�����tz��ؿ����z�6/��~1��&�2c��e쿡V���?����d��k8�,d�� ��޾ež�³������0��*"��o\¾f�ھ����r��y�3�`�^����*۴���`V���#���0���/�-y!�A�	�gRݿ�{��Һ����v�Z�z�\ё�&���<�:|��%�H1���.�f�������ڿ�M��JŅ�MIT�ѕ,�m���i���վ�3��dа�T����-�����
 ˾��S��}vA�Fq������ĿpD�������)��92�C�,����� ���̿y����P~u� 򂿧.���vǿ������\+��  �  �&W���M�{S5����/�⿅M����t�Ƌ5�V�	�e�ؾt꯾�S���x��R(q���k�֗t�� ��:���<����;���/B��{��B������m��~<�`�Q�L�V�$J�ߝ.�j!��;ֿ����ɑ���e��w����������.��WU?��mS�=hV��G�H
+��R�s�Ϳ�M��?H^��/&�j����,˾�N���"�������p�r�o��*}�����}����ž������ ��pV��֑�B�ƿ�;��'���D�TZU�whT�4B�'C#��\ ���¿틗��Ⴟ}���������Ͽ�j�N+��H��
W�q�S��?�Z� ���N�����bL�*�����ľۥ��w��ˊ��'������O���ݞ�xܹ��Y�%c��Z7��^t��y���3߿p���3���M��Y��R�P�:�������im���x��`�������w����/进+��7�v�P�A�Y��P��8����[��L�������w@�������4�ƾpQ��Z뙾o���]��`K��ֈ������Ҿ�z��FQ �B�O��`��gy�����t9�%�?�GAU��Z���M��r2�e��g޿mU���������ƿ}'���#���C���W��Z���K��@/�����5ֿM���D�n�\�6������0�Ǿ�g���+��$����������$מּ(�þ?�+7�1���f�����Ͽd�N+���H���Y���X��BF���'���aa˿
��JT��f�ϧ���׿.S�/�P�K�)�Z��]W��GC��#��� �48¿����)�Y��(��R��޾<��3=���Н�IØ�˚�� ����a�Ͼp�����q�A��~�U����T促f�}r6��P�}�[���T�T=�[:�}��[6���6��vF��%����/��˹�9c��:���R��  �  Hhu�o�j��2N�s�&�qb��gi�����:�5��3�Ͼˤ�ވ��/o�~�\�C�W�0�_���u�%w��l����ܾPl��H��>����Ŀ���H0��V��/o�i u�$f��JF�e��}^��{N���O��+`���%ҿ�E���4�r�Y�_q���t�
Uc��"B�j_���㿶u��:�h�%l(�ho���Z���盾�Ѓ���j���\��[��h��y��(6��cǻ���aA"��_�G��8�ۿ����=��`�sWs��/r���\�]9�
g�zؿe西\㍿����5-���q�i��`[B�k�c��u���q��jZ�U�5�&z��	ο�|����S�CI�W���O���Z��Z���Dv��n���r�'���Zv��x���Bؾ����;��ʀ���������GE$�+L��uj��Kw�M%o��/T���-�T��)>ɿJS���V���g���~ÿ����q)�T�P���m�x��m���P�˦)�C� ��ڻ�54��yE�������b��ݟ�[���O��?b��$���󄔾c���Z�Ǿ���� ��LV��"����˿�
�ø3��uY�T�r�1�x���i��%J�-"�O��/Ƽ�xқ��㕿�����ڿy��359���]�@Gu�T�x���g�&YF���k7�*���py�~�8����G�ᾃC��;��6���~{��F��M1��p���Zy��� ܾI	��2�FTp��P�����A����A�jEd�A�w��lv�Pa�l_=����/�%o���`��}d��j{���￢���%F�Ojg��x��u� �]�r�8����A�Կ����`�ra(�$����Ӿ"������jg��/��������4�����CTľ�����rE��셿^�������c�&�7�N��	m���y�N�q���V�[+0����οJ��*��T���"ȿ��� �+�:�R�֟o��  �  AH��,������lf��/+�du��⤿F0d�!�"���ǟ��s晾s}��̃u� �o��'y��c��|���qƾ�� �S$/���w�]���t��E8��\s�3^��&�����̑��U-��( Y�r� ��j�%����챿��п����'?�ަy��֖��$��y���ʪ��,X���qR��4�n�ԿX���
L�Nd��i޾�c��3���ԋ���t���s�����ϐ�d���r�׾, ���C�&ዿ	�˿�/�.�K�p)��2m���ը�i��w��1��V<E�#`��3ֿ�ֲ�0L������5��R��I��f̝�!���y��FG��	�z��m?�B��Z!��<����9�`����Ӿ}߬����/؇����}����.�����e�ľ���2$���b�8������m�&��da����jM��e4��4���Y���R�n�(�4��/���ʿ����+ƿ�����.�gLh����?�����5T��I����h���-������R���o��-����7Ҿ�谾5���뿒�+u��U���%��E����ྐ0�j�<�R����������;�a�v�X����%׫��s��:&���]��"%�.
���pÿ����ٿ;���C���}�����K������,̟��v��ΧV�ed��ݿQ��a|\�)�#�	���f�о:糾ע�����3��0M��T��IV̾b��yg�MT�����ӿ�V�`�O�C��ǉ��.����"��:����q�I������޿�v��῿)�w_���V��9��s���m����,��S����}��B�29���ÿ�_��#�F�l��v��0ƾ�٭��*���̚��Mߦ��4���Vھ�����.�t<m�������@)���c�v`��ܗ��x|��Ħ�?ؓ��q�7�.�� AϿ�3���ʿa1�>1�B�j��'���N���  �  ��h�������H\�He$��S迲Π��a��S"����n��M���~��7+}�`w�np��7o������ɾ���p.�Ȫs�5ɮ����m�0���h�����������\���CW���O����Q� +���Ӭ�*ʿu�d7��o�Gc��5����G���Ԗ�����O�I��a�,ο����J�������[_��~���}��Pu|�a{{�����I甾_����ھ���:^B���7�ſ$��'C�g{�w���?����Ġ�������t�*=���
�`1ϿC���^걿�ۿ�>��I�����n��F���>�����|�o�e�7�_��z᷿p���4�8���	��d׾4���1������Ȇ�!��� )���#��b�ȾP���5$�O7`��9����⿺v ��W����M���أ��m��/c��3�d�z-�����`Ŀ"{��s;������e�'�̬^�w����?���C��-C��q��3_�'�#���>���l�
S-�5���־�������
����6�������������T�98�#<�����t���2~�4��jl�I���/���$������GN��BT��������۽�M���4�ҿ��
�|�;� ss�L�������k��
���_�����M����}ֿ�<��g�Z��($�����Ծk��2Ȧ��{������8���0��\о�I�����L�R��O��2�Ϳ!��7TG��8�˖�j���<������,y�^wA� @��׿�I��Sy���q�d���M�q������{S��K��yg��Gs���:��O�s����"��'�E����� ��Dʾ�鱾���|�������r۪��Q���6޾#�ۮ.��j��]����9#��Z��O�����O!��@�������~g�r�/����jɿ�-���Ŀwr���(*�Z�`����M���  �  ڼ�������o���A�G[��+ӿi���C�Z��#�i���u�̾����d������Sv������$����M��˔־X/��M.�0�j�⎢�������4�L�X�x�Y�����������f�X`7�7�	��0Ϳ/֥�E���B���ͭ�@9"�"BR�cX}��3���,���'���a��2��� +��؂����F�ɣ��*�����b������o����v���H��]���a��\���?��q��	۵�tH����,�@e\��D������������8W�s&'��E�������j�������ƿ���72�#�a�逄����qm���}�<S���"�4<�ʊ����v�|�7�6��	����G��"��[����~��8�����վ۾�Z�%��Z�4���>ϿiQ��>�:m�(���������E�v��vI�����W� e�� ���6寿ln޿�7��]D��r����m��k��ۃr��D�J���ؿ2���ve�q�.�i
��I�+�¾߭�-���u���5���W"��\m̾�0� ����;�Eqx��z�����;7 �RP�QI|�Ќ�k]��ȇ��j�xl;�5����տ�v���f��uu���b���&���V�Հ�}Z���P��[I����e�M6��.��|ſ�Ǐ�M!W���&���Hk��vž�^���^��eө�Y�����¾�޾Ҧ�WK"��1P��������"K���0�[�`�a�����"��������[��q+��n ��Ŀ{���ی��AYϿ�	�$6�e�e�nS���A����O����RV��*&�����o,������D�<��X���l�׾���}Y��uZ������������˾?��f��w0�2e�J'���aԿ3���A���o�t��h��B��(y���K��`�"꿨���E��������;�F��t�&���  �  9e�<�[���A�����3��.X���܋�F�W��K+�L��ٞ�bdƾ'���ѡ������l���J���;w\�0��Q4���d�������ſP���J'��	I�B�_�Fe�d�W�7g:�Ѝ�^�a��� ��2��������ɿ�1��v*�[4L���a�ױd�HU��77����࿔��ro��m?H�� �����ݾ
��h��T����
��L���=W`پ�� ����ߥB���x��w����ٿ*���3��R�ڔc���b��O�vH.�`��o�Ͽ�3����������Ʃ��lݿ�����6�	�U�yUe�= b�3M��0,�����ο^k��9�n���<�c�"���ھ�W��𝮾�ާ��J��7Ǹ��&о���u���.���Y������b�������Y@�է[�T]g�T�_�~HG�I$�����h¿7�������:ޘ��̼��U���( �:1D�o�^��4h�%�^�)�D�ܴ!�#���	˾��M����b�.K6����;:��;iݾ�	ƾ]���9;������̾��zw�͟�1�A�M`r�����̿�c�<�*��|L�HNc�5�h��K[�V?>���g���������6��&�����ҿN�	���.�q�P���e���h��TY��t;��9�>C鿗Z��f����X���0��B��<��e߾T�ʾc쿾/G��l�Ⱦ�6ܾ¸��q7�>�,�D�R�W���{���k������Q7��LV��g���f�RS��2��:��'ؿ��������z_�����j���y���:�<Y���h�D~e��gP��|/��
�¯Կ#���|���I��l&�����]�I*ؾ��ƾo���ސ¾c�Ͼ�d�X��vU�%9���c��������0����h���B�tC^�D�i���b���I��x&����-�ƿ�>��Zl��Z����c�������["��SF�ӧ`��  �  +���$�
������:�˿�/��5���N�c���A�n�%�	������}վ��¾鮽�e"ƾ��۾)B������+��I���l�ύ��M���ֿ�p����'��*�r� ��3���俆h������=p��&h��xޠ�J�Ϳ�����(�O�*�� ����E��.���0A��H�X���8�D����s,꾃�Ͼ3&���Q��1;~V���?��G5��+T���z�~9���Ź�]忪
�]|��)�u�(������-ӿZͤ��%��g�h�~
m�#]��X���3m߿��	�B���+�sc)�?��@����ܿ�&�����u��mP���2�B������V込.Ҿ0�Ⱦ�B;k߾\���a��)�3�E���f�Aǈ�QR��$˿����k�t%�;-�f'�w����a�ƿ���kO���n�n�~�I���'¿�������?�&�=�-�C�'�R��_q���gѿ����*��>�n���L�Z�0�/�	a�%��+�ھ_"־K߾!���!��R ��_9�%�V��z�����9��X�ܿ���� �n+�4n.�r�$������I���"ꕿ5u�� 2y�;��� }����ֿ8W�@�:b,��/���$����*���ƿ@��)�����h�1I���.����^C����~e�#��nU��N��=��v+�^�E���d�h����z���¿	x�M���"��7.��-�q����\�ۿFL��0���x�y��}�����������N���%#���.��,�����9	�`n�9ƹ��H���&����]���?�L�&��h�^� ��}�����T���	���@�4�� P�Sq�Rw���8п#�����o(���/���)�ZX��
���˿M������Ox�b�����KwƿhU�����>�(��  �  р�N￳a޿a�ǿI��$����m��/q��GU��[8��b�F��t,��OS�����X�2A#��?�V\���w��m��y%������	��EyͿ�@�9����t�Kɿ�	��\&����^�	�A�n<��O�~x��_��[线G�ٿ�|�;O���0뿾�׿\��� 4�����H<���Ɓ�i�!�L���/�JE�V��#��n�ﾩ;����5�,��
I�~�e�h ������J���Tȩ���q�Կ���{�h�(ܿ"������W}�[�Q���<���?�8�Z�JK���㤿ƠƿI��n��,���翮�ѿ�'��7����n�������6~��0c���F��*��+����/�������P��!�b�;��Y�ru��Ǉ��Q��.C���ĳ�/Lɿ��߿6��k����x�d׿Z��
����t��P�V�C��N�i�p��9���$��U�Կ������ʑ����㿜xͿ����x���`��2⊿�0|�\n`�ѰC�$�(��v���U]�^��r��:30�f:L� si����+Q�����I ����2]Կ�&������������r�п�ǯ�����o�0gR��GM�>!`�����F����ÿW�3���������KG�?dɿ���������
����yy��\�i@��q&���������=Z�Ǽ#��<�	AY�]�u��K��Ɣ���G���jƿ�?ݿ;^� ��� �����\�ƿR�� ���?�b�}xM�	.P�k�j�o���v��h�Ϳ/�J�����h���\ؿ�����Z��`���A��𯅿�3p�yWS�$V7�?��q������
�5C��:,�K�F�Z�c����4����x��%h��S�}ο�'�=�������m��ܿ���u�ء~�M^Z�<M��W��y������m��ٿ���  �  ɂ��*J��|���
������ñ�R���=��U��r��[�z�c�Q�"#0��������l�6�5tZ�I#�����������Cò������C�����c���f��1E���/��j���t�e�K�zR,�9���*H"���<�U�a�����cڙ�騿�����t����i���'���β��+���뫿����ϋ�tUm�N(F��\(���D�ۼ%��!B��wh�uY��s���J������ʘ���������v����{��3��,��� X���ڇ���e��?�$��y����#�)�s�H���p��č�a���!��������6��"�����v>��Ì��_b��*䩿y��������c�\'?���%�w���U�� 3�îS�\l|�?Q���L��������ε��!���ӳ��O��\I���4�������:���؄��J`��e=�*4&�F����$��;��U]�Qi��bA��E^�������η�V#������畵��4�� �������ר�'���7�F#]���;�'��$!���*��eC��Pg������1��La��YӶ�Ӯ�������-��O���rK���\���V��\j�����w���A�[�/i<�~*�q�&�#3�	�M�%�r�����m��*z������Ƅ������ո������ ��/p���#���ڦ���:�}�\TV���8�~%(�;'���5��CR���x�t��G�����������\غ�RD���R���]���亿+���T#��ͣ��L���Xv�WcP�B�4���&���(���9��7X����� �����]���i���ֺ�.��?���๿i0����qu�����%���p�g|K���1�%�&��+��>�9�^�������������O�����}�1J����-���4����m�������V��t߉�)j�MG��/�+'�'.�i�C�0f�����b��Ig���  �  D�����������%7���Cɿ��߿Y�￳n�i���οlV��7Ì���d�J]D��;���I��Go�^�������ԿC��-.���W��7ۿςĿ�*��{靿�&��)����`m�i%Q��N4�����y�����B�w��P��>(�AoD�FMa�dd|�I���֪���+���Ժ���ѿ���w*�5��q��JĿ����!����yX��O?�u�=�(wT�cb��p����R����ݿiZ�~�0运�ӿܼ�ߵ��BĘ�y���TT~���c���F�{�*�Y��.' ����0��V��t���2���O���l�����R���ꝿ�����ÿ��ڿُ�����^�dڿ����~�����y��R���@�|�G��<f�k����׬��ο7��R���m����忲�Ͽf��N����� U���]}�D�a��,E�8�)��?�oV�������� �"y(���C��'a�@1}�ez�����5~��������οq��2��p���%� �ӿ`������g�p��VP��%G��V�I�{�N������yۿ*z����@���$�wm˿����Ӥ����J�����{���_��pC�N�)��^�y�	��������� ��:9�_~U�er�󽆿I��Q+��b���?ÿ��ٿ���Un���������\=̿���Ֆ���h��mO��N�z�d�0s���զ��lȿ��A���l���%o��ۿ-0ſ���*�����	����bt��W�[C;��"���������w��Q�'�x�A��L^�Y�z����(��+����\���Xʿ�.�z1��g��������v�M���ݟ������$^�0�L��S���q�%;���e��u�ӿ�/�����2�����P�Կu���Z嫿�.������ރ��/l�-BO�j�3���#���<��������1�R\L�7^i�l����  �  �e�����	���Rο���,�\�%�+�,>#����2�X��������4t�"[f�j.|�N���hſu��� ��4&��"+�,�"��s�b�(5ſ2������^��a=��""���
�WH�l�ҾLk¾9g���ʾ�~�}��r����0���N�8At�V���򵳿=�ݿy�C���&)��2*�n$�^&�N1ܿ�9���ꈿ7^l�Zj�`7~��YYֿ(C�7��])���)�t�����Ő�����s���!x���Q�93��k�|��F��=�˾���]I¾�Ҿ�3
��!���<�]�n�!��'W¿.���'/"���+�<f(�T��� �YIͿ��b��xwl�ǌv��A���U�����^#���,���(�`5�C��L׿T׮�Xߏ���q�՛N���1�މ�u�^�꾆i־�LϾ�վ��龥��p�bs1�@�M��p�;���������ӿI� ���[(��-��&�������n���Ey�����ur��5��j�����˿�y��j���)�(�.�Z&�����J���̿�릿�6l�,�K��0�������Q�ʉ�M྿8�������(��B�u`�j���,���*���?濫�
�J��H-�'N.�V:"��7�eL�;O�� ����{|��uz���������lm޿�O	�a �er-�J�-��!�����r翿_֝��w�� �b��D�l%*�-#��v�F�3྾����l�!��E�/��J�Țj�=�������v�ȿ0|��C0�2}%�&/�L�+�t�����jxӿT��X
��cx��+�����c]���+�����
&��U/�Z+����v�!Jܿ���Y���=|���X�.<�x�#� �K���j��ᾪ辿k���1��o!��9���U��  �  }�Z��荿F��Q����!��C���\�U�e���Z���?�����y����%��<z��o������cA���$��G��_�ee�P�X��<���Fp���������O�i�%����"|㾛þh۬�>����X���H���+��cԾ������{�;���n��I��N�Ͽ���n-��M�f#b��`d���S���4��b��ڿbҧ�/��� ������Qӿ�8�N�0�1�P��Oc��4c��P�=81����ֿ�Ϡ�gu���?�dO�;���/�־$!��B����.������ꬾ^�¾8�⾓H�e�$�DwM�ӻ��{3����1��A�9�I+W��e���a���K��k)��H��ɿ���é��Z���u|�����{�o�=�gZ��#g��`�4I��'����uJƿ�=���h��n9�W	��w��ξ۾��¾����Og���x���¾<�۾�����g��7���e�1n��p���w����#��F���_�?Gh���]�÷B�^��w������%��Q���?̞�?�ƿ�=��E'��TJ�9Tb�?�h��!\�V/@�Rt�-U�Q��� ���^��A4��v�~� �2��(̾�o��ʾ�s6ǾY~پ�����S���(� �L�N��Ť�VCؿ2)���1��R�zDf��{h�(�W���8��o��!�i㯿�����-�����bۿ�B���4���T��cg��Mg��T��[5�����p޿/��t肿W�P��
+�N��������ھ-�ǾK��|.���u˾��k����q�7�2�U[��i���ѳ�^��)�:2=�ptZ�X i�(�d�-�N���,��X��Ͽ����g���Ύ���Y��qg�����@��]��i�BEc�ǲK�R�)��Z���˿w��s�E�C�}K"�&�	���־�ƾ������ž,)Ծ�쾦�����?��  �  �^�^��I׿�����D�Xr��;��|��������m�KK?��}��ֿ�ԩ��[�������俹h�� J���v�!���j���Ã��y�h��:���]�ǿ玿#pP�	����J�Ǿʳ�����ъ�,��<�����������J߾[�D7�d�w��2��d��$�J�T�s�:�������|q��?@_��e/�����yĿ�w������d��� ���*�-Z�A���SV��+=���e����Y���)������\�����#g<�b��b��<���Ǡ��ݐ��󉾉���!���}쨾�5Ǿ����%�˓L�vd��r?¿*$�(�5�8�d��g��(Ҏ�y1���D|�2�P�� ���U෿����1����ҿ�6�r;���j��x�������^���kx��K�����5�'��d�m���2����p��.���Y���B��.&��m��mJ��k�����%�
�-�0�5i�<䞿��ܿ����hG�y�t�����!���u����p�V6B� t��ܿ֯�aa���������{�*BM�<z��B���P��6��~Rl��}=�$����ο�ڕ��^�gQ+��[	�OM��Ǿ�/��Ѓ���F���Y��/&��@ھ� ��L��>H��j����������(��Y�J����������|��	Qc��r3���Ί̿H������;ǿ:��n.�S^�����`��XI��Ut���^��.���&����Z��c#M��D ��K�1ܾ�c��
��/���w���u���S�ƾf!�"'�	�(��Z����G�ȿ�m
���8�:h�����o��oɍ�Ff�1�S���#�
���ٽ�	�������ؿ�!��O>�M^m�RԈ�6ؐ������ {��N�j��~l迣U���=x��Q=��)�����e�Ծ�{���?�������v��Gٻ���Ѿ���^�;�8��  �  �5e�D�� ��]'��n_�f�����5��4��!h���2Y�w�"��P�`繿�J��T¿���O.�ɻe�L����$��Т��������S���~�ڿm���B\U������꾢��k#���`����}��hz�<��ܸ���ܪ���Ҿ�k�B�8��u����������9�lDr�����k��c���ߕ�}~�l�F�O��)ٿ�6��~���ҿc���|@�]x�{����E��Q:��x����x�K
@���
��z���A��A�>���UC׾7���؈�������v|��t�{��h�������ĳ辥��րP��F��E�ӿ���Q�M��e���6������[������."m�'�5�P���ɿǶ��%-��-x�g���wT�Bw��c��d�������x����g��U/�˜��=ͮ�</v���2�NA�Y�־��������/���c��	X���\��q��k�վW���/��5p�܍��Z��*�)-b�Hl��2	���Q������B؈�="\���%�WP���꿿�M���Wȿ ��[1���h��A��ğ�y���:��+r���mV�_9����)���.jc�h=)�����׾�t���X��r��v_���磾�в�rJ̾�y���V��}I��B�¿�
��0>��qv�����@{����� �������J�����%�E���)����ڿ4��U�D�[+|�Õ�rO��QF�����@|��1D�	�\�ɿ5���7:O�Z���g��:�ξn��䘤�/ŝ�����[����ɒ־jo�{Z&��^�n�݄ڿ?�q�P�Y��cՙ�����w��B��.p��8�YL���Ͽҫ���!���g��!�[W��߆����������F��܎�r2j�W�1��������}N���=�ł�f����ƾjn������埾l]��Y殾�,ľv��#�G�7��  �  o�h�GJ�� i��zR.�Z\i��O��0ţ��J���+���p��5�b�r)�	������!S����ȿ�S���5��o�����?���*�����������J\��"��N�G7����W������羽2�����_g��\v��r�_�~������˦�{UϾ��9�9��Ӄ�K�����
�w�A�� }�� ��Ȭ���Q�� �������qAO�>�����t����U����ٿ�?�׷H������W��䇨�K����^������SH�yO��bǿ 房��?�al���Ӿ���z��8�����t�E�w�:.���q���ʵ���YC�ۚR����d�ڿ��<�V��C��e��QP�����[��
�w�^$=�5`
�.п�ȳ��о�c��4%�V�]�a]��|E��)��]!�����d�q�Ȟ6�����q���y��P3�)��Ҿ>ܮ�(����=�����������Y��X����.Ҿ���@	0�	�s��Э�����|1�Zl������#��X���'���z��?�e��m,��
��v�ſ/U����οbV�ߥ8���r�����Vݦ��ѫ��/���p����_�V�%��3��)��l�e��)��i���ӾpQ���W��a���m������������2Ⱦ������%�J��N���ȿ���$F���X4��޼���^������᷆�}NS����G�迠����b��N�ΌG�S�L�����V_��u���9���|m��1���{L�tz��Ͽ�B���P������zʾ{���ů�����ݚ��g�������Ҿ� ��	&�!`�_-��M]��: �$�Y�U������_��|�������-�z��#@��Z�grֿ齹��Ŀ������'��`��ƌ�����V���o���;��=qt��89��d�V����-��*�=��i�b-羯�¾*e���8���"������)⪾?��%�⾙���8��  �  �5e�D�� ��]'��n_�f�����5��4��!h���2Y�w�"��P�`繿�J��T¿���O.�ɻe�L����$��Т��������S���~�ڿm���B\U������꾢��k#���`����}��hz�<��ܸ���ܪ���Ҿ�k�B�8��u����������9�lDr�����k��c���ߕ�}~�l�F�O��*ٿ�6��~���ҿc���|@�^x�|����E��R:��y����x�N
@���
��z���A��D�>���DC׾�������a����u|��s����\���U���-�辳���P�"F����ӿ0���M��e���6��~���/�������!m���5��O���ɿ����6-��Wx鿉���wT�dw��8c����������������g�*V/������ͮ�k0v���2�&B���־������������c���W���[��{���վ����/�d4p�0������2*��,b�l�����OQ��͛��؈�"\�p�%�%P��o꿿�M���Wȿ��6[1���h��A��4ğ�=y���:��er��<nV��9����ڛ��hkc�x>)����D�׾
v���Y���r��`��b裾	Ѳ��J̾�y���V��}I�"�C�¿�
��0>��qv�����@{����� �������J�����%�E���)����ڿ4��U�D�[+|�Õ�rO��QF�����@|��1D�	�\�ɿ5���7:O�Z���g��:�ξn��䘤�/ŝ�����[����ɒ־jo�{Z&��^�n�݄ڿ?�q�P�Y��cՙ�����w��B��.p��8�YL���Ͽҫ���!���g��!�[W��߆����������F��܎�r2j�W�1��������}N���=�ł�f����ƾjn������埾l]��Y殾�,ľv��#�G�7��  �  �^�^��I׿�����D�Xr��;��|��������m�KK?��}��ֿ�ԩ��[�������俹h�� J���v�!���j���Ã��y�h��:���]�ǿ玿#pP�	����J�Ǿʳ�����ъ�,��<�����������J߾[�D7�d�w��2��d��$�J�T�s�:�������|q��?@_��e/�����yĿ�w������f��� ���*�/Z�C���TV��-=���e���Y���)�����]����)g<�_���a㾌<��7Ǡ�-ݐ���T�������v꨾3Ǿ����#���L�Bc��>¿q#�d�5�p�d�>g���ю�'1��wD|�ǩP��� ���෿����R���e�ҿ�6�fr;�p�j�y��ꅏ�0_��Plx���K����	7�q����m���2�]����!������NC��<&���l��7I������㾈�
�8�0��i��➿8�ܿן��gG���t�����L!���u��4�p��5B��s�*ܿ�կ�da��&����5|��BM��z�&C��Q��o6��WSl��~=���+�ο5ܕ�|�^�wS+��]	�;P�3Ǿ�1��P����G���Z���&���ھA� ��L��>H��j����������(��Y�I����������|��	Qc��r3���Ί̿H������;ǿ:��n.�S^�����`��XI��Ut���^��.���&����Z��c#M��D ��K�1ܾ�c��
��/���w���u���S�ƾf!�"'�	�(��Z����G�ȿ�m
���8�:h�����o��oɍ�Ff�1�S���#�
���ٽ�	�������ؿ�!��O>�M^m�RԈ�6ؐ������ {��N�j��~l迣U���=x��Q=��)�����e�Ծ�{���?�������v��Gٻ���Ѿ���^�;�8��  �  }�Z��荿F��Q����!��C���\�U�e���Z���?�����y����%��<z��o������cA���$��G��_�ee�P�X��<���Fp���������O�i�%����"|㾛þh۬�>����X���H���+��cԾ������{�;���n��I��N�Ͽ���n-��M�f#b��`d���S���4��b��ڿcҧ�0��� ������Qӿ�8�P�0�5�P��Oc��4c���P�D81�����ֿ�Ϡ�{u���?�aO����ֿ־� ��a���O-��F��笾��¾���cF�˲$�@tM�����1����#��0�9�?*W��e���a���K��j)��H�lɿʙ�����������|��F�����=��gZ�q$g��`�J I��'����sLƿm?��E�h�zq9���?{����۾ݨ¾����bg���w��8�¾��۾����He�F�7�l�e�Zl��j����t��m�#�~F�p�_�AFh��]��B�ҍ����������$��V����̞���ƿ>�^F'�JUJ�Ub�G�h��"\�|0@�wu�aW�b�����U^��D4�@y��� �����̾�q���˾��7Ǿ@پa���4T��(��L�]��Ť�WCؿ2)���1��R�zDf��{h�(�W���8��o��!�h㯿�����-�����bۿ�B���4���T��cg��Mg��T��[5�����p޿/��t肿W�P��
+�N��������ھ-�ǾK��|.���u˾��k����q�7�2�U[��i���ѳ�^��)�:2=�ptZ�X i�(�d�-�N���,��X��Ͽ����g���Ύ���Y��qg�����@��]��i�BEc�ǲK�R�)��Z���˿w��s�E�C�}K"�&�	���־�ƾ������ž,)Ծ�쾦�����?��  �  �e�����	���Rο���,�\�%�+�,>#����2�X��������4t�"[f�j.|�N���hſu��� ��4&��"+�,�"��s�b�(5ſ2������^��a=��""���
�WH�l�ҾLk¾9g���ʾ�~�}��r����0���N�9At�V���򵳿=�ݿy�C���&)��2*�o$�_&�N1ܿ�9���ꈿ:^l�Zj�b;~��^Yֿ+C�;��])���)�|�����ؐ�#����s���!x���Q�}93��k�G�����/�˾��LG¾�	ҾC1
�]~!�ê<�\]�V삿]���T¿���Q���-"���+�@e(����l� �\HͿ/���Pwl�5�v�E�����꿠�x_#�¸,���(��6�����׿�ٮ��᏿��q�N�N���1�.��0���꾹j־�LϾ�վ������/��p1���M��{p�����@����ӿ������Z(���-��&������}����x�����vr��5�������˿J{���j���)�Y�.�c[&�+��rM��p̿jZ�&;l�μK�(�0�����T�`��G�9:�~��p��Ҁ(�B��`�q���",���*���?濫�
�J��H-�'N.�V:"��7�eL�;O�� ����{|��uz���������lm޿�O	�a �er-�J�-��!�����r翿_֝��w�� �b��D�l%*�-#��v�F�3྾����l�!��E�/��J�Țj�=�������v�ȿ0|��C0�2}%�&/�L�+�t�����jxӿT��X
��cx��+�����c]���+�����
&��U/�Z+����v�!Jܿ���Y���=|���X�.<�x�#� �K���j��ᾪ辿k���1��o!��9���U��  �  D�����������%7���Cɿ��߿Y�￳n�i���οlV��7Ì���d�J]D��;���I��Go�^�������ԿC��-.���W��7ۿςĿ�*��{靿�&��)����`m�i%Q��N4�����y�����B�w��Q��>(�BoD�FMa�dd|�I���֪���+���Ժ���ѿ���x*�5��q��KĿ����"����yX��O?�z�=�.wT�gb��v����R����ݿtZ�~�0迣�ӿ,ܼ�󵨿UĘ�����eT~���c���F�E�*�����& ������U��r�1�2���O�N�l�����P��0蝿񾮿!�ÿ��ڿ?��Q����\￠ڿx�m���1�y�R���@���G�>f�R���٬�, ο3�迡���������忈�Ͽ�h�����y���fW���a}���a�o/E�/�)�6A�W�9�����V�Aw(�3�C��$a�R-}�x��6��s{��������ο��50�������^�ӿ�
�������p��UP��%G�LV���{�a��z���u{ۿ_|�w���B���'�vp˿���֤�����Ê���{��_��sC���)�r`��	�������q� �e;9��~U�?er����I��T+��b���~?ÿ��ٿ���Tn���������\=̿���Ֆ���h��mO��N�z�d�0s���զ��lȿ��A���l���%o��ۿ-0ſ���*�����	����bt��W�[C;��"���������w��Q�'�x�A��L^�Y�z����(��+����\���Xʿ�.�z1��g��������v�M���ݟ������$^�0�L��S���q�%;���e��u�ӿ�/�����2�����P�Կu���Z嫿�.������ރ��/l�-BO�j�3���#���<��������1�R\L�7^i�l����  �  ɂ��*J��|���
������ñ�R���=��U��r��[�z�c�Q�"#0��������l�6�5tZ�I#�����������Cò������C�����c���f��1E���/��j���t�e�K�zR,�9���*H"���<�U�a�����cڙ�騿�����t����i���'���β��+���뫿����ϋ�uUm�P(F��\(���H��%��!B��wh�{Y��|���V������ۘ��������������{��C��6���"X���ڇ�_�e���?��$��x������)�g�H��p�'Í�u���箭�+���E4��R����𱿯;��%����_��⩿����P���ބc��%?���%�L��[V��!3���S��n|��R���N��=�������е��$��oֳ��R��L��S7������V<��#ڄ��L`�g=��4&�V���$�L;��S]��g���?��-\��{���7̷�t ������꒵��1��m���P���cը�g�������=!]�v�;��'�%!�P�*��fC�Sg�n����3��c���ն���������1��`���hN��q_��Y���l��󂖿������[�k<��*���&��#3���M���r�4����m��6z������Ƅ������ո������ ��.p���#���ڦ���:�}�\TV���8�~%(�;'���5��CR���x�t��H�����������\غ�RD���R���]���亿+���T#��ͣ��L���Xv�WcP�B�4���&���(���9��7X����� �����]���i���ֺ�.��?���๿i0����qu�����%���p�g|K���1�%�&��+��>�9�^�������������O�����}�1J����-���4����m�������V��t߉�)j�MG��/�+'�'.�i�C�0f�����b��Ig���  �  р�N￳a޿a�ǿI��$����m��/q��GU��[8��b�F��t,��OS�����X�2A#��?�V\���w��m��y%������	��EyͿ�@�9����t�Kɿ�	��\&����^�	�A�n<��O�~x��_��[线G�ٿ�|�;O���0뿾�׿\��� 4�����H<���Ɓ�i�"�L���/�LE�X��*��w�ﾯ;����?�,��
I���e�s ������Z���gȩ�)����Կ/���{�h�(ܿ������}���Q��<���?���Z�KJ���⤿/�ƿ_㿙l�c*�����ѿ-%������jl��^���	3~�F-c���F��*�E*�$��ߝ������c���	!���;��Y��uu��ɇ�T���E���ǳ�Oɿ��߿ܠ�ֻ���z�(	׿������M�t���P�e�C�w�N�#�p��8���#����Կ�����������㿲uͿ��������y]���ߊ��,|�k`�8�C�9�(��u���`]������B50�"=L��vi� ����S��`��#������2`Կ�)꿿���������J�пɯ����io��hR��HM�"`�����t����ÿ(W�<���������HG�<dɿ���������	����yy� �\�i@��q&���������=Z�Ǽ#��<�	AY�]�u��K��Ɣ���G���jƿ�?ݿ;^� ��� �����\�ƿR�� ���?�b�}xM�	.P�k�j�o���v��h�Ϳ/�J�����h���\ؿ�����Z��`���A��𯅿�3p�yWS�$V7�?��q������
�5C��:,�K�F�Z�c����4����x��%h��S�}ο�'�=�������m��ܿ���u�ء~�M^Z�<M��W��y������m��ٿ���  �  +���$�
������:�˿�/��5���N�c���A�n�%�	������}վ��¾鮽�e"ƾ��۾)B������+��I���l�ύ��M���ֿ�p����'��*�r� ��3���俆h������=p��&h��xޠ�J�Ϳ�����(�O�*�� ����E��/���1A��H�X���8�D����v,꾈�Ͼ9&���Q��<;�V���?��G5�,T���z��9���Ź�o忴
�g|�!�)�|�(������ӿ8ͤ��%����h��	m�w\��r���l߿��	�^��|+�Kb)������0�ܿ�$��ѣ��#
u�BjP���2�������cT�c-Ҿ��Ⱦ�C;P߾b���x���)�x�E���f�kɈ��T���˿�����l�Tu%�^-�g'�K��^��Y�ƿ�����O�� �n���~�����<¿�������B�&��-��'����n��2eѿ�����'��5�n�E�L�x�0���Z_�����ھs"־�߾����#�U ��b9�ŸV�3�z�h���<��	�ܿ����+�`o.�x�$�c �J��`����ꕿ�u���2y�����[}��ޘֿCW�F�<b,��/���$����*���ƿ@��'�����h�1I���.����^C����~e�#��nU��N��=��v+�^�E���d�h����z���¿	x�M���"��7.��-�q����\�ۿFL��0���x�y��}�����������N���%#���.��,�����9	�`n�9ƹ��H���&����]���?�L�&��h�^� ��}�����T���	���@�4�� P�Sq�Rw���8п#�����o(���/���)�ZX��
���˿M������Ox�b�����KwƿhU�����>�(��  �  9e�<�[���A�����3��.X���܋�F�W��K+�L��ٞ�bdƾ'���ѡ������l���J���;w\�0��Q4���d�������ſP���J'��	I�B�_�Fe�d�W�7g:�Ѝ�^�a��� ��2��������ɿ�1��v*�[4L���a�ױd�HU��77����࿔��so��m?H�	� �����ݾ
��h��Y����
��U���If`پ�� �Ą��B���x��w���ٿ1���3��R��c���b��O�vH.�[��V�Ͽ�3��O��H���jƩ�lݿ+��Y�6�F�U��Te�?b�'M��/,�|���ο�i���n��<��`�^���(ھ�U��ڜ��{ާ�eK���ȸ�F)о��񾞬���.���Y�����}d��3��1���Z@��[�P^g�0�_�5IG��$�i����¿~������� ޘ�v̼�$U��[( ��0D���^��3h��^�
�D���!�����ɾ��K��c�b�aH6�I���6���fݾ�ƾ����I;����s�̾��gy�;��B��cr�i⛿+�̿�d�d�*��}L�dOc�8�h�sL[�@>����N�쿤3���7��h���քҿ\�	���.�u�P���e���h��TY��t;��9�<C鿕Z��e����X���0��B��<��e߾T�ʾc쿾/G��l�Ⱦ�6ܾ¸��q7�>�,�D�R�W���{���k������Q7��LV��g���f�RS��2��:��'ؿ��������z_�����j���y���:�<Y���h�D~e��gP��|/��
�¯Կ#���|���I��l&�����]�I*ؾ��ƾo���ސ¾c�Ͼ�d�X��vU�%9���c��������0����h���B�tC^�D�i���b���I��x&����-�ƿ�>��Zl��Z����c�������["��SF�ӧ`��  �  ڼ�������o���A�G[��+ӿi���C�Z��#�i���u�̾����d������Sv������$����M��˔־X/��M.�0�j�⎢�������4�L�X�x�Y�����������f�X`7�7�	��0Ϳ/֥�E���B���ͭ�@9"�"BR�cX}��3���,���'���a��2��� +��؂����F�ʣ��*�����d������t����v���H��g���n��e���?��q��۵�}H����,�Fe\��D��	����������8W�p&'��E�������j��:��-�ƿw���2���a���������m��R�}�vS��"��:���Y�v���7����e�����E��_��3���!��J𠾽�����վ^��3�%�M�Z�r��X@Ͽ)R��>�	m�l(��m�������͝v�KwI�����W�3e�����寿n޿�7�)]D�r�5�������r�?�D���7�ؿ���Wte�z�.��	
�CG�F�¾�ݭ���������嶥��#��_o̾N3񾳴���;��sx�|��M��	8 ��RP�,J|��Ќ��]��Yȇ���j��l;����
�տw���f���u��c����&�ƗV� Հ�}Z���P��ZI����e�M6��.��|ſ�Ǐ�L!W���&���Gk��vž�^���^��eө�Y�����¾�޾Ҧ�WK"��1P��������"K���0�[�`�a�����"��������[��q+��n ��Ŀ{���ی��AYϿ�	�$6�e�e�nS���A����O����RV��*&�����o,������D�<��X���l�׾���}Y��uZ������������˾?��f��w0�2e�J'���aԿ3���A���o�t��h��B��(y���K��`�"꿨���E��������;�F��t�&���  �  ��h�������H\�He$��S迲Π��a��S"����n��M���~��7+}�`w�np��7o������ɾ���p.�Ȫs�5ɮ����m�0���h�����������\���CW���O����Q� +���Ӭ�*ʿu�d7��o�Gc��5����G���Ԗ�����O�I��a�,ο ����J�������[_�����}��Tu|�f{{�����M甾d����ھ���?^B���;�ſ&��'C�j{�y���@����Ġ�������t�*=���
�Q1Ͽ+���:걿��ۿp>���I�~���G������=��Ѽ���o��7����෿ڃ��1�8��	�Uc׾-�|��0���
Ȇ�]����)���$����Ⱦ���� 6$�o8`�6:��B��w �|�W���9M���أ��m��Tc��l�d�<z-�����)`Ŀ${��];������>�'���^�S����?��C���B��9���_��'�c��9>���l�R-�_��Y־�����������6��\���O������	V�9�2 <�<���(����~�{4�kl�����h���Y���J���lN��{T�������ܽ�o���K�ҿ��
���;�"ss�M�������k��
���_�����M�
���}ֿ�<��g�Z��($�����Ծk��2Ȧ��{������8���0��\о�I�����L�R��O��2�Ϳ!��7TG��8�˖�j���<������,y�^wA� @��׿�I��Sy���q�d���M�q������{S��K��yg��Gs���:��O�s����"��'�E����� ��Dʾ�鱾���|�������r۪��Q���6޾#�ۮ.��j��]����9#��Z��O�����O!��@�������~g�r�/����jɿ�-���Ŀwr���(*�Z�`����M���  �  �3���P��s���Ȍ�4�P�����7¿>���-v8�r:���оl_���C���+�������2������:ѱ��ܾ���UG��f��@�Կ����`����9�����������Z"��<ԧ�Ô��u)C��c�rmڿYϿB���}I(�(i�ñ��X~���X��Z�������m������-�9����^�����i��k&�����<�þ�ꢾ����T���4��R��;ڟ�����P���J ��#`�������zt2�U�x�r���� ���n���k���A��ep��Y�p��V.�K����[п�ֿ�m�b�;�����8<��3���1�����������O��4�i��E%�l�߿q����R��u�d7�Ҕ���v��5�������������*���)پg
��9����8����Z��J�����ox���H�����+���&������5t[�YP�u��cKѿ:������S�hÍ�}�������������H���$���GS�	G�a�ǿB���rC�9Y��g羙c���ª��0������HS��_P���̾�i��w0��U�S���ۿM"!��d�\����H��0���
�������ש�r���}|G����,K� ؿ����ʳ,��qm�A���������������a����Â�b,>��;����oDz���6�I��\7�cWþ����즾�`��\���3���"߾*��+�0�H�p��W��	��k�6��}�˪��?����������g��L���|u�Ǯ2�7:��ٿ�޿����,@�Α��{5������`��2b��K�������L�l�0�(�Ԩ�
���`��&�����׾�Z���鬾pᦾ�D���p���Lʾ������G�C��/���¿���{QM�!��� í�B���c���k��S_������]�9� ��K��տʧ�=��CV������������  �  �@������SY��m���bH�sb����ޟ��8�[��.վ��8ɗ��x���4�������3��Nu�����i���XF�ی��aο����CW�����#���#������sѺ�����~��U;�S��ӿ��ȿ)|��!��j_�^>��ۦ��ћ���m���~��R��5_v�z�2���������Hg���&�i��T5Ⱦq����(���܊�aQ��w��\{���Gþ�_���� �^�B���U���x+�kWn�m������8���e����I��Qѕ�+�f�t�'�?���ʿ�qϿ��y4��Lv��J��K�����������E�������8�_��	�%Fٿ󔔿o�Q�j�1�n4þ����꘾GJ��\J���8���ø���ݾK����8�#J���۸�Z����B��ԃ��
������0'������g������ҋR�8l�_��,˿���7(��hK�\ه�?������ߖ��r������}����J�d��o¿���C�m����뾹ƾ�H���|���Ġ�a����ൾ�о���NN��T�,Ǔ��Uտ{A�_�Z�aD��fl�����l�������뷢�r��z�?�����nܿJ�ѿV��M4&�-�c��m��~Ӳ��������������r����z���6����[	����w��/7��S�]����Ǿჴ��,�������Ʋ���ľ����p
�=/1��qn� ʧ��=󿼢/���r�Ĺ��:��@�������<o������ k�f�+�����ҿoؿ���W�8�kez�7A�������|��В��Ǫ���c��c�~`"���߿�<���^��'�=��"�ܾ����~G��d�������︾.�ξ�A�K�uC�Qx�����
��+E����>V��&���o������Cά�ǩ���T�������Ͽ�P���Z�M�$������ ���  �  ����J��d���|�l�=1�Ͻ������ƫz�F9��]��.�/���a����gw���S��m	��]ƾm�e���E�%�������Z��C>�*Az�k6���$���s��B�����	�_�F�%���!���C����׿���
E��}���	�����������4����X�6���߿�*����b���)����׾XӶ�Mc���A��𩗾����������Ҿ�� �6s$�X�Z�� ����ֿ*���Q�һ��Oe��F"���m���R�������GK����$ݿ����$H��R�J ���X�|)�����xM�������)���р��E���/ȿ.捿P����څ����Ҿ���yΦ�����ͣ����f+Ⱦ��f���:��cy��	��������,��h�wɐ��c��������]���G�u��0:�]�Hѿ�J���̿���54�D1o�����������y��o��I�o���3��� �qg��Iɂ�)D�}�=����վ�ཾ��*���m����ľ�5�5�KK$��yS�/��ſI����A��}�d��>���B��K̥�7��a�c�f7*�^���۔ɿ{����w࿵|�vmI������6������U��Kӣ����&]��I#�\E迁u��]s��3:�U���-��k?׾�¾̑��-���������Ӿ6�:>�A�4���j��<���߿,��/V�׈�����9C�����x�����0�O��I�#��pS��'�ſ����F$���\�,���������	k���՜��{��:�H����%�ο����H]�^,�v��$(�<�Ͼ�*��pa������gǾ{b޾>��W��2E������/��M���c}/���j��������ܰ��+��>��-x�ܐ<���
�W�տ�����/ѿ�;��e6��oq�75��/����  �  �c��f��w�l�}�@�E��ݗڿ�����v���A�&��c!�Qݾ�����������Ʈ���5Ǿ�"�+��jm$��SL�_ۂ�W&���H꿗��tFK�cu�l҈�N<��vփ��wc��N5�5����̿�p���{��𷿯��A� ���O�>�y����+׋��%���*_���1�c"��ƿ:蓿{�c�E5�,��Ȑ���gԾ�޼�������������оI����0o0��-]�j#��K'��Њ�r,��Z��Q��,��9����%}�w`T��s%�\���7��^(��������ƿ�!��/0���^�ky���1���'���4z��,Q�TV#����E������(mU�6),����'򾗍Ӿ�k������\}����˾�^�d�ω ��YD�fw�l����%׿`����=��$j�����L���Ȉ�2s�wG�ܦ�8��/ʳ��d��1c���ݿY�B�^o��݇�����Ň��no�ΝC��g����p��"�����L�_(��o�J��[پ�ɾ�ƾ�;=�ྣH��� ��1��Z��ǉ�q��u;�� �#�N��x�\����������\g�i[9����ViտV��r4��1���H��t%��S���}��������KJ���lc���5��U
��_οQ3��1<t�"{E�^N$��
�����8ݾ0�оA>о�۾�:�|	�V� �Ѿ@��m�_���nǿ���(�0�O^��o���L���������T�X�f�)�@���קĿŷ��6���,Ͽ�9��&4�*�b��J�����d؋���}��}T�Z�&�Ѿ��[���;����b��@9������m�<�ؾǀоH�Ӿ�������F��5+���N�>���᥿�Kܿ�{�E@���l��V��\���"����u��sI����K鿺}�����k��}p⿄J�PED��7q�Q���  �  �:P�%cH�,�2����/�3}��?������ \�:�;����#���x�	پ��Ҿ�ܾ�q������%�\�B�ǥd��k��Y���a�ʿi��������8���K�E�O�!�C���)�G	���ӿ`f��w�������3˕�q����^��Ҏ�0p9���L�~�O��B���)�\
�*࿳���j��;�v�A�Q�h�2��w�F��L�Q�־'�վ&���� �����K/���M���q�!я����J2ڿ����g&�U4@���N��kM���;�����������{������ ���h=���Ϳ���F�&��A��P���M��2<�q� �_��saѿ���D싿��l��J�+-�N��xT�'�0޾B+�̑�����~�#�[D?�~}_��G������@����RY��1��H�:&R�t>K�wA5��ZW뿄��e���އ�|�����V%�e���2��J�`�R�%K��5����ӧ���ſŭ���t��g���F��#+�A���8�}�y����~����/3�]6P�!^r��W������}ѿ�j�� ��!<��4O�A�S��CG��y-�l��ܿ%ʬ��	���:��`w��|6ſ���#���=���P��	T�z	G��.�EE�a�迧����h��n����b�=C�=�(��B����������i�j�i�%�_�?�}�]�	��j���f��J��S��K�*��oD� S���Q��5@�5-#�>�&ʿ���������mv����տ��	��M*��_E��S�`!Q�q�?�y&$��P�v
ؿ����ŕ��'�y��2W�h�9�~?!�f���� ����W���k2���B�.�\�I�2 j�+x��0ߡ���ĿF8������S4�%K���T���M�g�7�o���1�պ�[ʘ������_�����Қ鿡����4��&L��  �  ���8���뿄�Ͽ�����|���̙�T���X�t�L>R��V2�������-�3|����,;9��Z��f|�1i��E���<���F��D�տq��tN�������������ƿ�N���t��*\��U��cl�3X������,�ݿ����v��l����-}��Fȿ{𳿥��[m���ⅿ"j�[	H���)�����������§&�:,D�Q�e��܃�����B����Uſ��޿@��{����B�����\�������s��y�o�55V�׸Y��Az�����*���Z��������	����U�ڿ�S¿.ů����z������7#b��6A�a%��&���	��o�����{5�8/U�U�w�����=꛿.����E����п44�����\;�l��V���M�׿r������Q�l���\���i��̉������Կ$���i���%�����C�Iտ&���Gꭿ?���:��g����]�]�=���$�D��{h������*��6F�@Vg���:C��P1���1���:ſ��ܿ�t����
��:��F�	y�7��*�Ϳ�Z������a�l���f���}�N���[��^E�q�X���ô��$������пUI���Q��{���H��eVz��JX���9��=#�������1!���6�P_T� v����2���]T��|�+�ͿD��@��@�]5����	���=꿬;���Vc����f�/0j�k4�������ɿ�l��`��W��u�����+���L�6�ȿes��sU��2���𕈿	 o�=�M���1��N�k��� �(�K�@�L&`�6��ݑ�����ï��k��pֿ�i�D�M��D���2�ƅ�l�ܿ芳�\X��\Kv�f�K!s��L��?a���Kؿ#� ���  �  ^Ϳ6ѿ5gϿ��̿DͿL�ϿEѿڳ̿ꬿ�͚��0-����p��@H��/�q�'��63��4P�F{�<�����,�ÿR�ο1_ѿ�JϿ4Ϳ��Ϳbkп�4ѿǂ˿H���fᦿ2����i�W�C�|%-���(��7��#W��������@��;Mƿs�ϿV{ѿ�Ͽ2Ϳ�Qοѿ��п��ɿ�蹿0٢�����b���>�=<+��'*���;��]�����ݟ�^n���LȿeSп{�п`8ο�̿�Hο��п�Ͽ�Jǿ4쵿����U��t�Z�3�9��Y)��+�ɏ@���e���������	����˿�ҿ�Yҿ��Ͽ��ο��пDӿѿǿ[��� !��w����DY�C�:�l�-���2��J�v�q�u����^��K���nϿQ�Կ��ӿ ѿ�п	�ҿ��ԿL�ѿ�Vƿ~��E���DT���V�.�:�dx0�	9�T{S�]�|���������ſمҿ�ֿ4�Կ�oҿ��ҿ�տt|ֿr&ҿ�.ſ�2��-ߖ��'|��T��;���3�Ӡ?���\���䮝������dʿ�տhTؿ�@ֿVԿ �Կ
V׿x,ؿf�ҿ�?Ŀ�X��M䔿l|y�P�S�l�=���9�O�H��Ch������U�������ο[qؿ�ڿ��׿��տ��ֿ�\ٿgIٿ ҿ�¿n��O(����r�j�N��b;�:L:�\�K�#�m�0������є���|п{�ؿ�+ٿ{�ֿ�տ!�ֿ�Eٿ�Uؿ�Ͽk������ˌ�E�k��TJ���9�{�;��rP�@u�瀒��M���ÿS�ҿ`<ٿ��ؿMMֿ�[տ]׿��ٿ,�׿B�Ϳ4
�������숿c�e���F��u9�'�>��"V�\}����ð��ƿ��Կ��ٿ{�ؿqIֿ��տ�2ؿ&+ڿ	׿l�˿����i����A��*`� &D�v�9�(B��g\�O���ԛ��-����ɿ�  �  z��H@��׎��8ѿ!B�<����}���
�����k�̿%��]����r_��T���e������¬��Kֿ�)��Y��u� �����	̿\����P�����<m���{o�RM��3.�������3��p�V�"��?��b`��F���;�����0��=¿��ڿX����k	�H��.�����鿮$��膘���w��"Y��xW���r�2����j���i���W0����k�
����VYݿ4Ŀ����M���k��ݤ���Sc���A�Ĳ$�
����o$���� ,��"K���m�<܇�����9��a��1˿����j�ɶ�N�z[�M��,ݿ\���qˏ�|�n�@Z�=jb����Z��TH˿;����,�����$��[��l����׿P����㮿�
��4����q�_���?�"�$�RU����ȁ��e#���=�7 ^��W���ߐ�y����Ʈ������ֿ¶򿗲��5�]�����g��svҿ�񩿹����wk��A`�mWr��>���&��g�ܿ�j�������W������}�ҿT���/I��Ȟ�-����H~���\���=�&��,�)��D��~3��P�O�q�x߉��ә�p���z���)�ʿ�"㿏 ����R����i�
��F�Dǿ����V����Hi���g�䆁��Ü�6�¿@������G�!����sq�J��[i̿5�������⚿��6t�ՖR��a5�iE ����a%��,$�+d;�~�Y��|�hڎ�S��������ѿ�7�_��������I����_����{���e�.n�����Ǩ���п,\����	9������
�͕���/ݿ!�ſ�"��$G��,f��%���j��pI�1�.�����>����C,�TRF��f�q���┿�  �  �#��,ߝ��¿U7���t��A4��FI��>P�t�F��y.��v�%ݿ�����&��	�������X���꿞����4��6J�_>P���E�$m.�i��4��g���S����]}�f�V�zL7�`M�"��5��Aؾ��Ծ�������z�*�}H�Q�k�Vȋ��|����ҿ���þ!�*�<�F�M�^O�x@�!�$�f����ʿG|���3������Rƚ��Ŀd���]� ��w=��N�N�C?�E�$�m���g׿����x(��-�n��-K��4-���������⾨kվ��׾~�龎��9��-6���U���{�j	���8���}俼q�6-,��D��P�'�L�|�8��������i�������d댿���^�ٿ+^�2�,�"EF��Q���L��
9�?���J��ʐ˿kO��m�����i�[uH�w&,�l�/����R��E-��|�7��|J+� �G�W�h�����ce��TȿE����.�G�6��K�M�R��SI��N1��Z�Y����,�� ���:���������%��-8���M��S��?I�t�1�wd�Ѓ�X���՚��{���nZe�BF��a+�[���n����������6�����"��<�:�Y�~�|��V��C����ڿ���%���@���Q��;S��7D���(����ҿ�����F�� ���آ�t�̿��3�$�s�A��3R�3�R��;C�{�(����߿�`������&��S	\��>��$������`���gw��kl�1��)�svD���c�%��������޽���j��1�/��G�T�e�O��<�o���&���%¿n���$����Ӓ�C��{߿�.�3�/��H�-uT��PO��;��S����v�пK���"鎿�Ht�úR�6B6�-W����t����)��XG��/O
��6��3�U�O���p��  �  u�y�����<I޿~�>qC���n�o���h�����OSj��=��V���տ�U���&��!\�����D���G�Bs��h���K��Pl��If�:X9�����п�͚���l�q;���t,���پ-���4���_1��n7����̾r쾷q�ι*�x�T����*������%%���R��i{��?��b���[n��:\�y�-�	�n\Ŀ%��0c��g�������F(��%W�g7�
�����u�~�V�W��)����ݻ��ˌ�%�Y��-������ξ�������౾-f���Oؾ�����w���9��ni�������ʿ�	�95��Mb��W��|t�����w�x���M��:����C���t��16���uҿ�/��S9��Rg�a��Q0���&�� u��|J�1������⭿�����Q�*���, ��g־�ž�5���ľ�־}�Q|��(���N�ii����������],F�`�q�=h���Ǎ�"Q���.m��?��N�I�ۿ^^��L6��Ks��3꿎#��J���v���u���%����i���<�cH��׿�š��{�A�I�}('�������߾�Ѿ��Ͼ�Uپi!��t�y�;��f�{��������4��mO)�v!W�����Q��C���fz��jM`���1���bq̿{7���t��L#ǿB���R,�E4[�����I������������[��.�G��XDĿ�6��Ϣj��>��[��d����!ھ��Ͼ�>ѾZ޾c=��2�B�%�UdG�w��M��x|ѿ�n�Dd8�Ӟe�����X��\����{�ZQ��H"�F��f���j���$��pYؿ��".<�gj�����M���Qr���w�mM��n���P ���ŉ�ql[��Y4��)�~����=ؾ��Ѿ�־���������2!1�/�V��  �  �~��_��g\ �Hh4�) p���� ��R���p����v��5yi�M�.������ſ_��)ϿՐ��?;���v�B��Ѩ��q�������o��Y�b�T(�>��P��{]n�=[1�R�	�� ޾����*¤���R
���x��x対�̾�>�����BP�������ʿ���;H����	��
��������n���y�U��p�������z7���࿪��Q�N��Q����������/ά��Q���/����N�>��vҿ#���uV���!����о�㱾�ʟ�Z痾�����󤾿����ݾS<���.��i�K������4�"�A]������ ���s���D����~���B�v��q.׿�����ĿPz��`2*�7Ed�	V�������m���S��
×���x�z�<�dw�킾�)����I��&�����"Ծ�g���ݫ�@'���꫾�h��X�Ӿ����Ϧ���F����v渿��F)7�h�r��s��_J��<������K��yll��1���̿�%��6տ���R>��z�����JN��L7���J���&��RUf���+��n��G��1s|�۪?��������پ��þt�`z���i��;AѾ���S��s�.�Ra���.ӿ3��<sL��+��(��� ���ͯ��������ҞY�G}!����A�Ŀ�H¿�
鿈�� �R��X��m��������ۮ��a���B����R��I���ڿ�i���Bg�)d2����񾂣Ҿ���_���gƸ��oþ�}ؾ����c��}<��v��J����_#&�!Y`�C���g���EA��z��G՛�R���E�̻��#ݿ<�����ʿ2j��3#-��(g�D�����������'���n���J{�G_?��
�d�ÿ�c���FT�zm&�_+�� 辒�;"۾������G�˾d�侳���"���N��  �  S#���
��W���K�������Ҡ���B��۽�����)���ؕE��b�^�ٿEǿ��e�7T��{��`"���k��X��2л�w������G2=����D���@�t��F/�O��ξt����Y��$������|���k㠾i���뾣{��?R����рܿR�!�2�b��:�����#)�����5V��It��3�r�sc1�t� �ۀοp�˿�r��p�*���j�ɗ�,���8��(��E����ԗ��wj�(����y��|Y�E���D�ΐ���ޢ�
ّ�����M��bǖ�K���t�;N����+��en���������6�.{�{������)���l��x��������\��
 ���1�ʿ�ؿ��
�S@�
���9$��j���b����8��Q��=|���4U�e�DͿx���5J�f���Y��ľ����!��-虾xI��<ƫ��Tľ��뾇���E�'���0�ƿJ�*�N�����U������ĥ���E��*���<��ڙH��j���߿yͿ��2�0!W�]������ ������,����+��@����@��_�����f{���=����l��ʾ�r��QX����`]��s&¾<߾�u��{*��Ic���������%�zg�iS��!���:��\.���a���}��p�v��o5�����ֿt�ӿ5� �6�.�x�n�%Й��Ķ��B��q5��V��������n��:,�6��y��ZCj�Č.����h�ᾮ�þ��h\��Z��	&���.ɾ���(��a�9��{��g������1:�Y~����F�������}��dC���l����_��#��v󿹗пN ޿ ��p�B��������
��'I�����9T��[Ɏ���W�i��ҿ�В�crT��<!��� �usؾ���V��pi��TM���M���dվ_���q:��M��  �  v?���|ƿ˰�d{T�@ю�ɜ��TG��5���Q��2��y�����M�������)'Ϳ�X���K,]�����ų������K��Щ�����s%E�3�����x��C/�����hʾ�ޑ�OU��F����&��'I��:͸�6,������S�4&��(|��'���l�����������0����|���S��!}�C�8��z��տ]3ҿ[4���1�-�t��}��uļ�������ռ�J���8�t���.�i^�wt���_[�'���I��H���z�����}���[���馾�Rɾ� �x�+��q��ٯ�����v>�b�������x�����9#������G���Gf�2c&����N�п"�޿���H�RD�� T��=��o�������hд�oΓ��W^���!nӿ������J����72龚￾T���͙�b���J����>�����������H�F�8���j̿8u�k>W�w1������Ϧ����������؃��s����P���}翢0ӿ\�"�#3`��5���X��U���{������U��� u��E�H����������=��H��&��Tžb	���ϥ�r�都�_ھ�Û)���d��������q;,��q�,���-������������]��������<�̈́	��ݿVDڿ=��5��y����-;����.�����
à���x�3����5٧��$l� �-�p����ܾ�澾����� �� ��E���ľk;�U<���9���~�\�������A�����FN����3���>����	���ɘ��Ai�HY)�������ֿ����2�J�2���k����h��%7���@���������`�(����ؿ96��pFU�w
 �do����Ӿ߃��~ɬ��1�������ĸ���о�\������~N��  �  S#���
��W���K�������Ҡ���B��۽�����)���ؕE��b�^�ٿEǿ��e�7T��{��`"���k��X��2л�w������G2=����D���@�t��F/�O��ξt����Y��$������|���k㠾i���뾣{��?R����рܿR�!�2�b��:�����#)�����5V��It��3�r�sc1�t� �ۀοp�˿�r��p�*���j�ɗ�-���8��(��F����ԗ��wj�	(����|��|Y�D���D𾱐��pޢ��ؑ�����M���Ɩ�b���R�;���$�+��dn�e��������6��{��z��f���)��ml��Z��������\��
 ����+�ʿؿ��
�o@����S$����������9��~��j|���4U�je��Ϳ����J� ��[���ľ����M"��3虾6I���ū��Sľ�������E�������ƿ���N����RU��v��������E���)���<����H��j���߿zͿ��G�Q!W�t������F������\����+��o���g�@�`�����{��˓=�������0ʾ�s���X������]���&¾q߾�u��{*��Ic���������%�zg�iS��!���:��\.���a���}��p�v��o5�����ֿt�ӿ5� �6�.�x�n�%Й��Ķ��B��q5��V��������n��:,�6��y��ZCj�Č.����h�ᾮ�þ��h\��Z��	&���.ɾ���(��a�9��{��g������1:�Y~����F�������}��dC���l����_��#��v󿹗пN ޿ ��p�B��������
��'I�����9T��[Ɏ���W�i��ҿ�В�crT��<!��� �usؾ���V��pi��TM���M���dվ_���q:��M��  �  �~��_��g\ �Hh4�) p���� ��R���p����v��5yi�M�.������ſ_��)ϿՐ��?;���v�B��Ѩ��q�������o��Y�b�T(�>��P��{]n�=[1�R�	�� ޾����*¤���R
���x��x対�̾�>�����BP�������ʿ���;H����	��
��������n���y�U��p�������{7���࿫��R�N��Q����������1ά��Q���/����N�B��vҿ)���uV���!�� ��uоF㱾Fʟ��旾�����������ݾ ;�"�.��i�F�����忙�"��]�N�����v����s��YD����~���B�L��C.׿�����Ŀ�z���2*��Ed�:V�������m��T��_×���x��<��w����*��[�I�Z(�!��>$Ծ�h��Dޫ�K'��R꫾�g����Ӿ����l��ڜF�!���\帿>��(7���r�`s��
J�����r�����&ll���1����̿�%��?6տ��MR>�%z����N���7���J���&��Vf�K�+��o��(H��7u|���?��l���&�پ|�þ��`{���j���AѾ��u����.� Ra�󅗿�.ӿ3��<sL��+��(��� ���ͯ��������ҞY�G}!����A�Ŀ�H¿�
鿈�� �R��X��m��������ۮ��a���B����R��I���ڿ�i���Bg�)d2����񾂣Ҿ���_���gƸ��oþ�}ؾ����c��}<��v��J����_#&�!Y`�C���g���EA��z��G՛�R���E�̻��#ݿ<�����ʿ2j��3#-��(g�D�����������'���n���J{�G_?��
�d�ÿ�c���FT�zm&�_+�� 辒�;"۾������G�˾d�侳���"���N��  �  u�y�����<I޿~�>qC���n�o���h�����OSj��=��V���տ�U���&��!\�����D���G�Bs��h���K��Pl��If�:X9�����п�͚���l�q;���t,���پ-���4���_1��n7����̾�r쾷q�ι*�x�T����*������%%���R��i{��?��b���[n��:\�z�-�	�o\Ŀ%��1c��i�������F(��%W�k7�
�����{�~�\�W��)����'ݻ��ˌ�/�Y��-����ώﾕ�ξޣ��w𯾄߱�?d��Mؾ�����u�v�9�li����>�ʿ	�Y5��Lb�RW��t��i���x�8�M��:������t��V6��vҿ�/�aT9�pSg�ha���0��'��u��}J���o�鿇䭿���P
Q�*�:��"�hi־�ž�5��P�ľf־�z��z�%�(�C�N�h��q����+��n+F�r�q��g��iǍ��P��9.m���?�AN���ۿ+^��O6���s�����#���J�=�v�f�������%��y�i��<�OI�~׿ǡ��{���I��*'�|�����p߾��ѾT�Ͼ�Vپ,��!��t���;��f����������4��mO)�v!W�����Q��C���fz��jM`���1���bq̿{7���t��L#ǿB���R,�E4[�����I������������[��.�G��XDĿ�6��Ϣj��>��[��d����!ھ��Ͼ�>ѾZ޾c=��2�B�%�UdG�w��M��x|ѿ�n�Dd8�Ӟe�����X��\����{�ZQ��H"�F��f���j���$��pYؿ��".<�gj�����M���Qr���w�mM��n���P ���ŉ�ql[��Y4��)�~����=ؾ��Ѿ�־���������2!1�/�V��  �  �#��,ߝ��¿U7���t��A4��FI��>P�t�F��y.��v�%ݿ�����&��	�������X���꿞����4��6J�_>P���E�$m.�i��4��g���S����]}�f�V�zL7�`M�"��5��Aؾ��Ծ�������z�*�}H�Q�k�Vȋ��|����ҿ���þ!�*�<�F�M�^O�x@�!�$�g����ʿI|���3������Uƚ��Ŀi���`� ��w=��N�!N�I?�M�$�u���g׿�����(��;�n��-K��4-����r������ajվ�׾(����7��+6��U�s�{�����6��y{俰p�+,,��D�%�P�X�L���8����?������������댿����ٿ�^���,��EF���Q���L��9�S���L��Ӓ˿NQ�������i��wH�r(,��m�/ ����g��e,�|�ʝ��H+���G�g�h�ѡ��|c���Qȿ����-�.�6���K�[�R��RI�N1�Z��㿐����+�����Q:��A������%�7.8�y�M��S��@I���1��e�
��v���ʜ��=����]e��F��c+�#��`p����a���a7����H�"�	<�\�Y���|��V��E����ڿ���%���@���Q��;S��7D���(����ҿ�����F�� ���آ�t�̿��3�$�s�A��3R�3�R��;C�{�(����߿�`������&��S	\��>��$������`���gw��kl�1��)�svD���c�%��������޽���j��1�/��G�T�e�O��<�o���&���%¿n���$����Ӓ�C��{߿�.�3�/��H�-uT��PO��;��S����v�пK���"鎿�Ht�úR�6B6�-W����t����)��XG��/O
��6��3�U�O���p��  �  z��H@��׎��8ѿ!B�<����}���
�����k�̿%��]����r_��T���e������¬��Kֿ�)��Y��u� �����	̿\����P�����<m���{o�RM��3.�������3��p�V�"��?��b`��F���;�����0��=¿��ڿX����k	�H��.�����鿯$��醘���w��"Y��xW���r�6����j���i���\0����r�
�)���hYݿFĿ����[���k��ं��Sc�`�A�x�$����1��z#����,�� K��m��ڇ��}���7���^���˿����i�����M��Z����+ݿy����ʏ���n�Z��jb�������`I˿�����-�����%��\�Ko����׿�����宿����5������_�b�?�B�$��U����J���d#� �=�	^�IV��5ސ������Į�H��(�ֿT��g��~4�Z����^f��Muҿ��,���wk��A`�Xr�?���'����ܿek�q����
Y������ҿ����`K��ʞ�饏��K~��\���=��&�0.����D�u3�P���q��߉��ә�t���{���'�ʿ�"㿎 ����Q����i�
��F�Dǿ����V����Hi���g�䆁��Ü�6�¿@������G�!����sq�J��[i̿5�������⚿��6t�ՖR��a5�iE ����a%��,$�+d;�~�Y��|�hڎ�S��������ѿ�7�_��������I����_����{���e�.n�����Ǩ���п,\����	9������
�͕���/ݿ!�ſ�"��$G��,f��%���j��pI�1�.�����>����C,�TRF��f�q���┿�  �  ^Ϳ6ѿ5gϿ��̿DͿL�ϿEѿڳ̿ꬿ�͚��0-����p��@H��/�q�'��63��4P�F{�<�����,�ÿR�ο1_ѿ�JϿ4Ϳ��Ϳbkп�4ѿǂ˿H���fᦿ2����i�W�C�|%-���(��7��#W��������@��;Mƿs�ϿV{ѿ�Ͽ2Ϳ�Qοѿ��п��ɿ�蹿1٢�����b���>�A<+��'*���;��]�����ݟ�fn���LȿrSп��пq8ο.�̿�Hο��п�Ͽ�Jǿ9쵿���|U��+�Z���9�/Y)��+�{�@��e��������#��ʻ˿�ҿIWҿi�Ͽ$�οH�пӿѿZǿℴ���������CY���:�G�-�G�2�ߠJ���q������_���L��ppϿy�Կ��ӿ�!ѿ��пf�ҿ��ԿP�ѿ�Xƿ���r���%U���V�ʪ:�qx0��9�=zS���|�~�������ſ҃ҿЅֿ��Կ�mҿ(ҿ4	տ3zֿi$ҿ�,ſK1��ޖ��%|�iT�;��3�q�?�-�\�������8���gfʿ�տ�VؿCֿ�	Կ��Կ�X׿�.ؿ{�ҿ�AĿLZ���唿v~y���S���=���9���H�ADh�˜���U��&�����ο]qؿ�ڿ��׿��տ��ֿ�\ٿfIٿ~ ҿ�¿m��O(����r�j�N��b;�:L:�\�K�#�m�0������є���|п{�ؿ�+ٿ{�ֿ�տ!�ֿ�Eٿ�Uؿ�Ͽk������ˌ�E�k��TJ���9�{�;��rP�@u�瀒��M���ÿS�ҿ`<ٿ��ؿMMֿ�[տ]׿��ٿ,�׿B�Ϳ4
�������숿c�e���F��u9�'�>��"V�\}����ð��ƿ��Կ��ٿ{�ؿqIֿ��տ�2ؿ&+ڿ	׿l�˿����i����A��*`� &D�v�9�(B��g\�O���ԛ��-����ɿ�  �  ���8���뿄�Ͽ�����|���̙�T���X�t�L>R��V2�������-�3|����,;9��Z��f|�1i��E���<���F��D�տq��tN�������������ƿ�N���t��*\��U��cl�3X������,�ݿ����v��l����-}��Fȿ{𳿥��[m���ⅿ#j�]	H���)�����������ʧ&�D,D�^�e��܃��������Q���Vſ��޿T�������H�����Y��混��s���o��4V��Y��@z�ڟ������K�������~	�Ί���ڿ~Q¿ï�!����������� b��4A��_%��%���	�&p����}5�>1U��w�C���웿;����G����п�6�6����]<�M������w�׿P���������l�	�\��i�Ỉ�����jԿ������
���������FGտ����"譿-=��H9�����f�]���=���$�����h�����*��8F��Xg�Y��D��O3���3��`=ſw�ܿew����
��;�H��y��8��f�Ϳ�[��������l���f�!�}�����6[��rE�q�X�������$������пRI���Q��z���G��eVz��JX���9��=#�������1!���6�P_T� v����2���]T��|�,�ͿD��@��@�]5����	���=꿬;���Vc����f�/0j�k4�������ɿ�l��`��W��u�����+���L�6�ȿes��sU��2���𕈿	 o�=�M���1��N�k��� �(�K�@�L&`�6��ݑ�����ï��k��pֿ�i�D�M��D���2�ƅ�l�ܿ芳�\X��\Kv�f�K!s��L��?a���Kؿ#� ���  �  �:P�%cH�,�2����/�3}��?������ \�:�;����#���x�	پ��Ҿ�ܾ�q������%�\�B�ǥd��k��Y���a�ʿi��������8���K�E�O�!�C���)�G	���ӿ`f��w�������3˕�q����^��Ҏ�0p9���L�~�O��B���)�\
�*࿳���j��;�v�B�Q�i�2��w�H��L�W�־/�վ0���� �����K/���M���q�,я����Y2ڿ����g&�^4@���N��kM���;������������P���r�������<��e�Ϳ����&�N�A��P���M�|1<�f� �U��v_ѿ	���ꋿҐl�J�,-�ɓ�lS�����/޾�+�o���9��I�#��F?�E�_�fI������=���"�gZ�(�1�	�H�)'R�E?K�%B5���&X�������އ�B�����$���X�2��J�o�R��#K�g�5�k������m�ſݫ���r�� g�!�F��!+��?�*��O�}뾆�����o���13��8P�4ar��Y��󋪿%ѿl� ��"<��5O�7�S��DG��z-����ܿ�ʬ�
��;;���w���6ſ���*���=���P��	T�w	G��.�CE�]�迥����h��m����b�<C�=�(��B����������i�j�i�%�_�?�}�]�	��j���f��J��S��K�*��oD� S���Q��5@�5-#�>�&ʿ���������mv����տ��	��M*��_E��S�`!Q�q�?�y&$��P�v
ؿ����ŕ��'�y��2W�h�9�~?!�f���� ����W���k2���B�.�\�I�2 j�+x��0ߡ���ĿF8������S4�%K���T���M�g�7�o���1�պ�[ʘ������_�����Қ鿡����4��&L��  �  �c��f��w�l�}�@�E��ݗڿ�����v���A�&��c!�Qݾ�����������Ʈ���5Ǿ�"�+��jm$��SL�_ۂ�W&���H꿗��tFK�cu�l҈�N<��vփ��wc��N5�5����̿�p���{��𷿯��A� ���O�>�y����+׋��%���*_���1�c"��ƿ:蓿|�c�F5�,��ʐ���gԾ�޼������������оW����<o0��-]�s#��V'��֊� r,��Z��Q��,��<����%}�y`T��s%�K�����*(��Q���X�ƿ�!�4/0�s�^�y��>1��K'���3z�,Q�xU#����­�������jU�6',�����$��Ӿ�j��z����}���˾�`�ue��� ��[D�"w�軠�1'׿?����=�n%j����M���Ȉ��s��G�0�����iʳ��d��c����ݿ��B��o�Q݇�����CŇ��mo���C�g�8�jo������d�L�a(�n����}YپN�ɾ�ƾ��;���K��z�(�1�DZ��ȉ���7=�� ��N��x�ђ����볅��\g��[9�����iտ����4��b���/H��}%��S���}��������JJ���lc���5��U
��_οP3��/<t�!{E�]N$��
�����8ݾ/�оA>о�۾�:�|	�V� �Ѿ@��m�_���nǿ���(�0�O^��o���L���������T�X�f�)�@���קĿŷ��6���,Ͽ�9��&4�*�b��J�����d؋���}��}T�Z�&�Ѿ��[���;����b��@9������m�<�ؾǀоH�Ӿ�������F��5+���N�>���᥿�Kܿ�{�E@���l��V��\���"����u��sI����K鿺}�����k��}p⿄J�PED��7q�Q���  �  ����J��d���|�l�=1�Ͻ������ƫz�F9��]��.�/���a����gw���S��m	��]ƾm�e���E�%�������Z��C>�*Az�k6���$���s��B�����	�_�F�%���!���C����׿���
E��}���	�����������4����X�6���߿�*����b���)����׾ZӶ�Oc���A����������æ����Ҿ�� �?s$�b�Z�� ����ֿ.���Q�ջ��Re��I"���m���R�������GK����$ݿm����G��� �=�X�N)�����3M��U���o)��bр�R�E�Q��.ȿ8卿�P����������Ҿ`���ͦ�����jͣ�����,Ⱦ��쾴����:��ey��
�����(�,�6h��ɐ�.d��^���.��������u�1:�3]�qѿ�J����̿z���4��0o��������\���y������o���3�� �Wf��OȂ�zD��{����n�վ�߽����4��mn���ľp7�`��L$�a{S�3�:�ſ���Q�A�̹}�������?C���̥�m����c��7*����� �ɿ�����w࿿|�|mI������6������T��Iӣ����&]��I#�ZE�u��\s��3:�U���-��k?׾�¾̑��-���������Ӿ6�:>�A�4���j��<���߿,��/V�׈�����9C�����x�����0�O��I�#��pS��'�ſ����F$���\�,���������	k���՜��{��:�H����%�ο����H]�^,�v��$(�<�Ͼ�*��pa������gǾ{b޾>��W��2E������/��M���c}/���j��������ܰ��+��>��-x�ܐ<���
�W�տ�����/ѿ�;��e6��oq�75��/����  �  �@������SY��m���bH�sb����ޟ��8�[��.վ��8ɗ��x���4�������3��Nu�����i���XF�ی��aο����CW�����#���#������sѺ�����~��U;�S��ӿ��ȿ)|��!��j_�^>��ۦ��ћ���m���~��R��5_v�z�2���������Hg���&�j��U5Ⱦr����(���܊�cQ��w��`{���Gþ�_���� �^�F���Y���x+�nWn�n������:���f����I��Rѕ�*�f�r�'�4���ʿ�qϿ����x4��Lv��J��,�������d������������_�<	��Eٿs�����Q�[i��/ﾉ3þ;���꘾6J���J��89��gĸ���ݾ�����8��J��Hܸ�����B��ԃ���	���Z'��ϑ����������R�Ml�t��,˿��$(��hK�Gه�"����������D��k���O��i�J��o¿����C����]���ƾH���|���Ġ�����"ᵾիо���O�uT��Ǔ��Vտ�A���Z��D���l��N�������ʹ����������?�����nܿb�ѿV��Q4&�/�c��m��~Ӳ��������������r����z���6����Z	����w��/7��S�]����Ǿჴ��,�������Ʋ���ľ����p
�=/1��qn� ʧ��=󿼢/���r�Ĺ��:��@�������<o������ k�f�+�����ҿoؿ���W�8�kez�7A�������|��В��Ǫ���c��c�~`"���߿�<���^��'�=��"�ܾ����~G��d�������︾.�ξ�A�K�uC�Qx�����
��+E����>V��&���o������Cά�ǩ���T�������Ͽ�P���Z�M�$������ ���  �  `��������U�����6k��"�+׿E��� NG�Q��b�޾���f)��e)��a����S��uנ�K��K�뾜E�}�W����s��1�Il}�p��<�������o���
��K������s�[�ڙ��������s�<�`���@������p�������t������9���iQ�������
=~��73�l���Pо㬾�6���p��|ߍ��m������S�ʾ_� �|,�uys��w���d��H��x���/��dm��2���9����,��M|��������C�����������JS�b���5��z��3��Ǿ�������������@�9�����p�66d�Ə$�ח���ʾ|Ѭ�+����і�F{��ꍾ�L��{�S4G��w���?ѿ����Qd�eQ��#u��;��[�����������D��w�`1�"B��|忡���;�*�nn��ɟ�rO����=&��?"��a���K���m�G�$�!~ܿ1���HR�@��L��|̾p���J2���T���z��{���uW׾�+���(�Y�e����7�7�4�iw���ީ��������I��l���dW��س����_�K!�Z�������c�U7A�����s��o:��z���g���s���ܧ���W��>�U�+�^_Ŀ`���C��=�W��Y;*���kʮ�w5���ƶ���ɾeh뾍����<�����϶��F���M�����L������:�������_S������u��<H��W�'����6�f�W�2���6��E`�����E{��m@������)a��J�<�r���ӛ��Xzq�D�1��;
�ҋ���ž ��W���54��!3����Ծ�Q���!��Q�q����eֿ�x�Y�f���|���.�����������"���r���]y�(Q3�ߓ�)��J���,���p�Y���l��f���  �  ޵�����Qͼ�����ra�k
��ѿjq���F��{��X�e������Ɠ��C�������å�¾� �p���V����s��M=*���r��ݠ�h��������\������5O��xM��٬R�i���鿜�ܿ�&��Y5���{�����<���������������������H����~���L{���3���w.վ�䱾��������k��z-�����)�Ͼ�� -�6q��U��i����@��|��\��v'��h������8����������;�����ݿ08俆Z���J����1k��AB����������������FN|�m2���%�����b�x�%������Ͼ�ı��m��4X������O��-�þ�R�����F��u����˿�K���Z�I�������������$.��m��)g���l�D*�����n�޿t����'$���d��!��*���Cq��1���k���)���u���)d�L��:pֿp㒿;�Q����6���� Ѿމ���ϫ��٨�R#���x���Wܾ�_�:*�CXd������뿺�-�Gv�����������_4��J���$X���l��<W��=������������9� !���3���k������[����4�����$��a+M��,��̿��煿��C�:�����ZҾ8b��dY������\�����ξS�����a=�U������������D����kx���F��y��������^���5��[;��xV@�TW�����ױ�XO�P����h��l%����������@��Y5������5�q���\G����o��2�Q^�I�辘�ʾ�й�%-��6̵��	¾$�پ� �A��(xQ�ۤ����пD��k�]������a��5*�������n��P���z���Do���,��7�X:��8��Y�&��g��F����������  �  <	��ۀ�����`����UG��c�����c����G�l��?�� �ʾ�����h��Ą��7Ӥ��µ���Ҿ_���]�!��U��D����ҿ�j��1V��-�� ����������{���E���|�$I:������ӿE-ɿ�?�@!���]�a������}���9.���`��«��Ջt��2�����UQ����u�ͥ6�����得^¾�P���f���à�_�������ཱྀ�	���0���l�7Y���N�ǌ+���l�w	���г�aH������h���#����	e���&�n���{Oʿ��Ͽ:Z� �3��xt�$�������������C���_I��]�^�;|�H9ݿ>ǚ�ٙ`�b*��*�A�߾����`��7�����c⺾b5Ծ������H�l4��1�Э�rB�.����@��C�������ݐ�����Xx��)6Q������忰~˿��۱��/J��ǆ�Z��"���a��_޽����V��J���&BǿDՍ���R��#� ����EȾ�p��������� sϾA#��B�YX/��]c��5����ٿ�����Y�����y������M���Jٺ�BF���$����>��^���ܿ�ҿ� ����%�bKb�4���$������WW��t���Ν� �x���6��� ��������G��1��8���⾱�̾���{����ʾX߾D� �b9�pA��}��������t�/�-�p��%��6��tj��t������¯���^i��+�n_���ӿMؿ���=�7���x�8ݝ�Ἰ�U���T��N���I�����a�b�"���㿅u����m�<�7�_��[����ھP�Ⱦ�r���Wľ�Ѿ�n꾣��A&��#S��c��]ÿ�@���D���g����޼��4������(6��o���l�S��6�#��*п�S�c��}L��������*���  �  
s��2���=u���Y�TD%��;�u������0�P��q(�pE�
��Suξ�E��z��S/��n=Ծڰ��mG���0�q�\�/8�������r�0�1�d��a���`��E���Ҕ��S��L�u���a�v�f譿%*ʿ�7�W4���i��ٌ������˝�Rђ�ֈ{���G������ڿ�d���lv��B�#���I�Ik�A�Ⱦ񵻾
򺾈�ƾ��޾ŕ������=�m+o�	����ҿ"d���A���u������s������o�Q�9�i�	���ο���β��Uۿ�x�F��i{�>���-���ԛ����Ek��7����pƿ~e���'f��8��v�����J̾��þҮǾ�+ؾ���tO�m�+�zS�����{������!�= U����c��VW���H���
���_���*��*����Ŀ �������`V���}%��IZ�����*6���Ο�-��ֆ���[�f�'�����'㶿�/��u�[���3�%��������LվYѾ�Hپv���p�����:>�$Jj�)���ſ̙�L	4��_h�����!��K��ϲ��uJ��bP�O����i���g�ҿq�	�\�8�1_n�R���ޝ�����T�������K�������W���;x��#FS��.�a��ip��N��ܾ�F۾`��Q����Y7+��N�f���G��/�ڿ�����E�z�����.��D��� 	����s��1>�����׿�R���Z����ę�J�z?�,�����-���������n��l:�}�
��#Ϳ_��Kns���E�oe%����u����g�Hs۾l�޾������X3�)r6�A�]� ӊ��������W_$��W�$2��,i������ ���VJ��Jnb��?-�� ��qɿcP��qſ�����'���\�Oԇ��>���  �  G�j�O�a�Q�H�H�'�|��\�ӿ�l������	n��CJ���+�������q��$��Ύ� G����2�pR�]`w��������B'߿H+�gj/��O�re��bj�7Z\���>�8d�F �X������c鏿����oп����.���P�|f��j�'[�4�>�H?�T���#�Ŀ��������bb�ʉ@���#��P�����Z��8��p���	��� ��<���]��ׂ��i���ɿ�+�K7�R�:��BX���h���g���S�s2�җ���տ�Ϧ�k��iR������?�㿫W�8%;��9Z�cgj�Ŭg�%�S�;4���l��Ң���՗�ܰ���Y��9���

����>)�S����{���/�5�M�7q�\���w��v7ҿR�e�%��YG��a�7�l���d���K��(�����ȿ�������Y����¿�;���#$���H�&rc��nm�*kd�5�K��B*�k��@ٿ�ٯ�?���y�fU�x67�E%�A�Ԣ���{���M����%�_�?�ݝ_�(���G���K����濣��e�2�yS�_�h���m��`��B�^e�]D�&μ�7��ۗ��KM����ؿQ+�A�2�L%U�W�j�`n��r_��B��| �15 �K@Ϳ�c��G܍���r�R�P��4�,��V�������2%
�����0��M�.@n����j���ȿ�����h�0�>�&�\�m>m�T�k���W���6����v|޿j^���똿�����ͷ��	�pA���>��]���m�sk�9�V� i7�e�qj�V������n|����f���F��+��y��/�#�r��L���!��u:�]X�u�{�?��	���D_׿1���.(�u�I��%d�6o��eg��IN�l|*��'���̿b���ݸ������]ǿaY��P&���J��|e��  �  ѕ#�y�� ;�s�e���:˿1!���觿�D��"����c�~@�m9$�/���r�
����)�'H�}�l��Z���P��f���PD����п��|u�~����!�O #�����GYۿ�ۭ�����n�̹f�c2���Ŝ�uTƿ�f��<W� ���#����:"�/9����ۿH�Ŀ�!��C��ؑ�^7~��uX�L�6������U�u���w3��0T��y����,����T¿�ؿ�����&��O#��� ��&��*����ʿY���5��Tg��@k����(���C}ֿ�l����=#��J#�\4��7	����;�Կ�����>��0��d���u�isP�^�1�S�"����'� HC�alf�=^�����۩�}����̿�`�^{�zf�/� �s�%��^����I�e�����0��Z�m���|�Lޕ�!��������2���S&�r�"�Y���3��/�h�п􌽿�Y���Ü���Ao�]L��0�������!�R�6��U���y����t0������>ÿ��׿���y�	��@�kR%���&����#\	�b4㿇����O����~��w�4Ո��s���Ͽ���ů�jh$��0(�!��f��Y��a�X6Ϳwp���I�����+G��m�h�,$G���-�\E ��~�d�+���C�id����Ǘ�m&���D����ʿ������$=�`c��'�E%�m�F�� �ӿݨ�ܬ���x��{��!��,~���(޿6�P[��&�-�&����<�����Üۿ��ƿ0�%�����O����]� >�k}(����"�513��N�eq�����56��p��9����ѿ]��f�-��i#��O(���!�Y/��E��.�Ŀ؝�ק����v��܂��^��e��<���N� ��  �  ��⿢��`�u6��W῕�����pK� �ӿ�껿O��c��X��e<��H4��A�ȅa�����ǥ�:¿�ؿVZ�����係O�⿫�忐 �.�࿜�п�������%~��ES��=:���5���E��9i�፿����r�ƿ#ۿM�� 翊���a���
R���Z!߿�-ͿK���ϕ�v���M��8�J�6�FhJ��p�0��ʰ��"fʿ"cݿ�#��H�o��s��u��{@�����Hܿ�ȿ��������bm�4H���5��8�(�O�#Ly���h��fpϿ��T�Ә�\�}�⿔e�������ۿ4�ƿ"/���S��kk���H��:��,@��Z��<��� ��IQ��2տf��d��G��;x�H��T��_��(����ڿ4TĿd
�����$�g��iH�=�`�F��d�E:��򱥿�¿ڿ�)迳@쿦��=�������8쿓�翛Bٿ����wˤ�RĈ��td��mH���@��M�0n�(r���a���ȿ1�޿�K뿬��G뿸C���Ё쿋���	�I�׿�#���D��������c���J�F���V�joz�ǅ��꠳��2Ͽm��TD���F쿜��\9뿷�ￅb�$cտc9��g�&$��*^��BH�GG���Z��i��ʚ��Mҷ�a�ҿŕ�#a��[�EH�vK�U�'�����=ѿ�6������D~���X��F�|�H�O�_�ul���x�������~ֿ?���￞@��A�鿡쿡E� ��v�bͿљ������pw��U�vF��K��f�:∿æ��j���vgڿ� 꿊�ￚ	���g���$�￭��9�߿.rɿ���o��G<q���Q� OF�U�O� m�����,奔�ƿ޿�  �  ���������f̿oV�<i�s��f �m�#��G��	���ӊ��{�����q�ce�g=y�����xm�������0���#�av�P��<���bO�iȿh���'���ĭ�� )���[^��;��!�Ml�߂�8��2�.�`vN�>�s�u���<h��.�������'�Կ�.�&n	�D>�<�"��N"��d����tqӿc=�������j�Z�h�ヿ�ܢ��	ο�9��bZ�nf!��?#�����!��Q��L"׿��� 诿濟�I����v���Q�Q1��%�k����wN�a9��[�A���瓿.��Hh��fǿ��޿��������^�$��S �'!����_�ſ]����Z��k��tt��4��A첿�࿙Z�3z��	%��,#�Ժ�{B�����ҿ�ξ��c��������:r�~>N���0�'J��9��R�{�.�;L�]�o��/��@����+�����^�ѿ9�뿽"����!#��@&��
�������e��fy����}�s8q��͂�����%�Ŀ����1<��!��a'���!��@�>F��>�)�ο�������盿������m�R�K��21��!�3�[�)���?���_�\`��%]��T���;���ȿ�Vݿ1���^��Dl�*'��n&�O�����ۿ�Y��������z���x���������$ֿ@-��n�\%�9^'�����K�Ѱ���߿�ɿ�`��?<��Ŗ�Bヿmb�B��*�:'�E� �4/��H���j�3;���隿^��� ���οu����."��y!�m(��#��`�����?̿���Sf��� w��������������W��"�/�'���%��L�t�	���Nؿ�Ŀ�����6���1���P|��"X�g:���&�~���f%��7�G�T�Whx��H��X����  �  �S��EE���Uֿ����s)���J��b�K�j��_�wLD�M������̐��[����Ǝ�G;��b�ƿ����$(��K���c�O�j���^���C�d�!��� ��%̿�.��"T��INh���E�&�'�e���F��z��m���0�H��L����7�^X���~�ᗿ�W���D�����@5�oIT���g�sli�hX���8�I!�ڄ�g���ݒ��q��}H����ٿ���4��dU�!Nh���h��V���8��V���W������N]���][��:�o���j�M�Ob����p����l�J�&��D�=�f�^#���.����ȿ����_���A�+#]�� k��f��
P�{-�
��U9Ͽ�$��_�������\���T���H0B�'1_�^Il�_[f���O��?/����߿�(���$��,e|���W� �8�M��z�
�����Ӓ�1�����	�����7�plV�\�z�
ԓ��˱���ۿ%Y
��,,��FM��`e�Drm�(�b�]#G�}"���������ٞ���ݔ� `��!�̿L���_+���N�LJg�en�P b�sVG��_%��V��ӿ�(���d����v�kGT��7�� ������6��x�������-��#I�(�i�a��v��9���1��r	�nu9��vX�<�k�Y�m��\���<�Q2�Ϡ�����񚿥��� ]��G��f��3�8�zxY��fl�V�l��[��<�:��G]����ſ���Ӊ��Dl��XK�sj/�]�6v	�2�����3T����pS5�mfR��t�����i橿6nϿɱ��:"�&xD�C}`��un�3�i�_CS���0���
��Nտ�(������e6���������D���a�r�n�<�h�:XR���1�˶���Ai��c���f���a�
�B���(�BO��P�S���o�+��:4&���?�P�^�e���  �  ���\���|��� (�T�[������a��Mx���.�� ;����T�
s ���Z~��uk��ě¿���Ö+���`�dI������ S���f��ϵ���oP��]�濺:��Xb����I��#�:�����
̾^⼾0&��p�þ��پ1����j��~7� f�G*��`ȿA	�Z99���m��ɍ�����-�������jx� C�C�܅ؿm ��Z��Whҿo)�[=���r����c��Ü�aΏ�7s���>����;�ο^h��sk�=;��������"Uܾ�bžyٺ�J伾'w˾�g�k�s:"��|G�Sq|��a��T�߿��9kK�5�~�����m��]����.���h�<�2��"��ɿЯ�鹿%n���VjP�Zi��Eu��F<��袚�+��W�c��/����r������`� 6����A��S㾫�оs#ʾ�>о��q� ���Ͳ4��<^�����⹿i��F�*��^�s��H���|ן�7���������W�ro#����ԍ��<��K�ȿ���X�.�$d�K��槛�(	���!��.r����S�`� ��84���p���;X�dD2�����#�K��N
ݾ��ھZ$�����:�u|'�J�H��4w�ﺝ���п���#t=���q�b�����紟��&��o|��(G�!�2��5��-���|ڿ�4�u$A���v�n��b����ў��ߑ��:w���B�-�#]׿-ء�S|��K�G�)����T��j��M�ھ�Xܾ�9�W4�5��~v0��aU���]��`}濏I��N��'���ƕ�V���=���ō��,k���5�k%�E�ϿCƵ�ڿ�V�:��GS�a΃��ϗ��������o_���Xf�h2��8��ÿ�甿uZk�Cf@�ƥ!��/�Z������\�ܾ�L�P���U	�����<�:f��  �  Zъ���ſ�A�{�J�u��v��0k��������0��W����eD���/�ٿ�Rǿ�o��m�]�R�-T��ꃪ��g������7���>��������<��/��¶�p���?��>���i�ƾ�箾T������t躾�Uھ�.��x)�]9a�F>���S��!�u�a�rÒ����!���9���������O�p�,y0�%� �´ο�̿S���*��i�|x��H�����q���8���=I����h�;7(��P�=����0h���-����G�ݾ����w��;�����㮾�Xƾly�����;�\�|�#(��[���6�ey�<ǝ�$�������Y�����	����Q[��^�T�.�ʿz$ؿ��
�t�>���������ƺ�4���2 ��}��
.���:T�� �|�ѿ8��ObY�=�&������B	ž�Q���4��0K��_�ľWH�kN�L%�<zU�dR���B˿?�¶M��ӈ��u���Ⱦ�Ko��(U����80���jG������߿�cͿ�~꿟w��U����������͌��]��7p��媁�t@@����޺���|���VM���!�fk�@~徕2ξaG¾���9*ɾy`ܾT ���1���:��Ur��ˤ�����0&���e�;ݔ���������
������� ����t�܆4����?�ֿ# Կ)� �).��"m�J�������%������[���1]���m��h,�W��c��~y���>���2�����ݾ+�ɾ����0���Rr;j+�zF�k��8�I����ݷ�� ���9��n|��n��ْ��i�������u���u7���S^�oY"�yF���п޿���D�A�%��L��F%�����RN���g���z��k�V�ݿ��&׿TR���c��@1�w;�����|ؾ`OȾͷ¾ RǾik־�[�̠��;-�5v]��  �  �K��j�տnp��e��I��֝�����h���'�����@ʕ��l^����@B�mڿB���^B+���n����*��� ��������9M��֘��U�oJ���ÿ�O��h�<�j���hܾG��oa���ғ��ӑ�r������.�ɾ�����$�3�c�E������Yv5�K���H��J���32��Pk�������a�����DG��5�&�H�߿��
���?��_��A��/����g���S������}X���J��n�<�����d��I�k���)�+c ���̾�Ѭ�3s��c����g��-����쵾��ھ�
�O�8�y��q������y�M�����9��[��������P�����Yp��F�x�+3��h��2޿���ܸ���W�h%�����F����_��f���Q��*���I/p�Ed(��W㿚s����Y��l!�uG���о���׊��O������A���ϾRt��U&��U�͕�n.ۿ5"�2sh�?�������z���������i��!K��3xa�"��Z���|��i��E.�s r������������0��0������O����X�����ʿ&[���EK�.��:����ԾE���8����?������̾97�����5���t�R��������9� ��Kb��`����D���z��?���l��Bˊ�.RK��@��+뿚迣����C�0f���H������'s���a������@l���`��bA����γ���|�gy:�����;����w��]��������Ӿ����x���F��D��ۨÿL�Q��D�������j���#�����2������[�{��6��^��&�M�󿠸���Z�ם���_��������8���]�����)�r��+���迕���Hd��+��D����ˍȾ����4x�������ƾ��ྛ��XG'�[	]��  �  ����G�ۿ��%��o�G:��b;��@������ܥ��S/���Z����g��>%��u���_ῐ���(2��Dy�:z��������������Y^���������-^�w���#ɿ-���=�B�
�?�׾�A������d=��CL��!g��e¥�;�ľ����� $�Քe����)����<�����Ӯ�[����,��En�������������	�O�/��t�꿟3�n��|�G��!���Ȳ������\��[�������P*��a�D�&H��Q��7*n��
)����CȾ�ߧ����v9�������ܚ�Q�I־���~�8�7������~���lV�-������'?��K����#��^������ ����k:���4志���� �c�`��R��7��Gt��߾������/���}�z�
�.��;�Z>����Z�F, �[���b˾�1���䡾�r������8��%�ʾ����\��K�U�C��v�ῄc(��or�T���~���?��.8�����(���ݝ���j��N(�����vn�����)5��I|�����O���z���J������H��ԙ�\�a��*��пJ8���WK��z�4p���Ͼ>������#����M��xǾ�6��f��5�P�v��������A�g����_���V?���}��&����"��:�����S����Ę��F�S��j�K�E(��iд�^���>h��-i������'���@���H��{�9�����~���9���y��Ⱦ^ ����V����C��w�ξq�����F�V݉��vȿ�-�ҸY�u�����������+<��%���Pf��@���5��j^=���e(�¬����#�#�c�����q��mv���������#��x��;;}���1��|�+{��jOe��t*����޾�þ�ാ�򯾪��������۾L?�=�%�ȸ]��  �  �K��j�տnp��e��I��֝�����h���'�����@ʕ��l^����@B�mڿB���^B+���n����*��� ��������9M��֘��U�oJ���ÿ�O��h�<�j���hܾG��oa���ғ��ӑ�r������.�ɾ�����$�3�c�E������Yv5�K���H��J���32��Pk�������a�����DG��5�'�I�߿��
���?��_��A��0����g���S������~X���J��p�<�����d��L�k���)�%c ���̾�Ѭ��r�����5g������쵾��ھF�
���8��x������P��4�M�t�����7���υ��jP�����Hp��-�x�+3��h��2޿�������W�w%�����`����_������w��O����/p��d(�:X�
t����Y��m!�~H���о'�����T���Ҡ�����A�ϾOs���%�1U��̕��-ۿ�4"��rh���������z����������h��K��xa�"��Z���|��i��E.�� r����+�������0��V������O����X�\��&�ʿ�[���FK��.��;����Ծ
���ӧ��g@�����̾g7�&����5���t�S��������9� ��Kb��`����D���z��?���l��Bˊ�.RK��@��+뿚迣����C�0f���H������'s���a������@l���`��bA����γ���|�gy:�����;����w��]��������Ӿ����x���F��D��ۨÿL�Q��D�������j���#�����2������[�{��6��^��&�M�󿠸���Z�ם���_��������8���]�����)�r��+���迕���Hd��+��D����ˍȾ����4x�������ƾ��ྛ��XG'�[	]��  �  Zъ���ſ�A�{�J�u��v��0k��������0��W����eD���/�ٿ�Rǿ�o��m�]�R�-T��ꃪ��g������7���>��������<��/��¶�p���?��>���i�ƾ�箾T������t躾�Uھ�.��x)�]9a�F>���S��!�u�a�rÒ����!���9���������P�p�-y0�&� �ôο�̿U���*��i�}x��I�����r���:���?I����h�?7(��P�C����0h���-�����ݾB��w���젾���a⮾RWƾ{w���0�;�ȟ|�A'��(Z��c�6��y��Ɲ����r���~Y��}��诏��Q[�n^��S�&�ʿ�$ؿ�
���>�.���!����ƺ�n���t �����P.��C;T�"!�m�ѿ���cY�{�&�����F
ž{R���4���J��m�ľ�F�qM�%��xU��Q���A˿��6�M��ӈ�ku���Ⱦ�o���T��Ȥ��0��UjG������߿�cͿ��w�K�U����$��$�����J]���p��/���A@�D��ػ���}��xXM�6�!��l���4ξ�H¾Ǩ���*ɾ�`ܾ� ���1���:��Ur��ˤ�����0&���e�;ݔ���������
������� ����t�܆4����?�ֿ# Կ)� �).��"m�J�������%������[���1]���m��h,�W��c��~y���>���2�����ݾ+�ɾ����0���Rr;j+�zF�k��8�I����ݷ�� ���9��n|��n��ْ��i�������u���u7���S^�oY"�yF���п޿���D�A�%��L��F%�����RN���g���z��k�V�ݿ��&׿TR���c��@1�w;�����|ؾ`OȾͷ¾ RǾik־�[�̠��;-�5v]��  �  ���\���|��� (�T�[������a��Mx���.�� ;����T�
s ���Z~��uk��ě¿���Ö+���`�dI������ S���f��ϵ���oP��]�濺:��Xb����I��#�:�����
̾^⼾0&��p�þ��پ1����j��~7� f�H*��`ȿA	�Z99���m��ɍ�����-�������jx� C�C�݅ؿn ��[��Yhҿq)�]=���r����e��Ü�cΏ�<s���>����F�οgh��sk�>;����`����Tܾ�až�غ��⼾pu˾ce�
��8"��zG�o|�t`����߿U��}jK�z�~�����m������.��+h���2�e"���ɿsЯ�<鹿on�!���jP��i���u���<��A�������c���/�F��fs��M���0�`��6�[��-B��T�j�о�#ʾ->о���j� �����4��:^����Sṿ� ����*�F�^���꼙�(ן��K���`�W�.o#���򿪍��?��{�ȿř���.�t$d����2����	�� "���r��T�S�(� ���5���q��>X�FF2�5���$�\���ݾ��ھE%徯����:��|'�c�H��4w�󺝿��п���"t=���q�a�����洟��&��n|��(G�!�2��5��-���|ڿ�4�u$A���v�n��b����ў��ߑ��:w���B�-�#]׿-ء�S|��K�G�)����T��j��M�ھ�Xܾ�9�W4�5��~v0��aU���]��`}濏I��N��'���ƕ�V���=���ō��,k���5�k%�E�ϿCƵ�ڿ�V�:��GS�a΃��ϗ��������o_���Xf�h2��8��ÿ�甿uZk�Cf@�ƥ!��/�Z������\�ܾ�L�P���U	�����<�:f��  �  �S��EE���Uֿ����s)���J��b�K�j��_�wLD�M������̐��[����Ǝ�G;��b�ƿ����$(��K���c�O�j���^���C�d�!��� ��%̿�.��"T��INh���E�&�'�e���F��z��m���0�H��L����7�^X���~�ᗿ�W���D�����@5�oIT���g�sli�hX���8�I!�ۄ�i���ݒ��q���H����ٿ���4��dU�%Nh���h�$�V��8��V�&��W������U]���][��:�M���j���0a�H��a����k���&��D�ޞf�"���,��B�ȿ���~���A�V"]� k�q�f�h
P��z-�����8ϿK$��Q������\��#U�{���0B��1_�Jl�2\f���O��@/���e�߿S*��V&���g|���W�ݡ8����\�
�������i�����	�m��H~7�MjV���z��ғ�Fʱ� �ۿ9X
��+,��EM�`e�|qm�{�b��"G��|"�	���S��������ݔ�;`����̿���`+�@�N�Kg�4 n�4!b�dWG��`%��W��ӿ�*��f��\�v��IT��7�M"���������?���-�$I�C�i�h��v��:���0��q	�mu9��vX�<�k�Y�m��\���<�Q2�Ϡ�����񚿥��� ]��G��f��3�8�zxY��fl�V�l��[��<�:��G]����ſ���Ӊ��Dl��XK�sj/�]�6v	�2�����3T����pS5�mfR��t�����i橿6nϿɱ��:"�&xD�C}`��un�3�i�_CS���0���
��Nտ�(������e6���������D���a�r�n�<�h�:XR���1�˶���Ai��c���f���a�
�B���(�BO��P�S���o�+��:4&���?�P�^�e���  �  ���������f̿oV�<i�s��f �m�#��G��	���ӊ��{�����q�ce�g=y�����xm�������0���#�av�P��<���bO�iȿh���'���ĭ�� )���[^��;��!�Ml�߂�8��2�.�`vN�>�s�u���<h��.�������'�Կ�.�&n	�D>�<�"��N"��d����uqӿd=��¦���j�_�h�ヿ�ܢ��	ο�9��fZ�sf!�@#�����!��Q��]"׿���诿𿟿I����v�m�Q��P1��%����H��YM��_9�>�[�$���擿�,���f��Gdǿ��޿	���������$��R �� ������ſ����AZ���k�Aut��4���첿���*[��z��
%��-#�˻�zC�����ҿ�о�$e��8��
���;r��?N���0��J��9��R���.��L�w�o��.��Ҁ��*��K���g�ѿ/�뿶!����0#��?&�
�������Md���x���}�|8q�΂�>�����Ŀ�����<�˚!��b'���!��A�KG��@�+�ο𪼿Ч��Z雿䕉�ϡm��K��31�%�!��3��)�D�?���_�r`��1]��Z���;���ȿ�Vݿ/���]��Cl�)'��n&�O�����ۿ�Y��������z���x���������$ֿ@-��n�\%�9^'�����K�Ѱ���߿�ɿ�`��?<��Ŗ�Bヿmb�B��*�:'�E� �4/��H���j�3;���隿^��� ���οu����."��y!�m(��#��`�����?̿���Sf��� w��������������W��"�/�'���%��L�t�	���Nؿ�Ŀ�����6���1���P|��"X�g:���&�~���f%��7�G�T�Whx��H��X����  �  ��⿢��`�u6��W῕�����pK� �ӿ�껿O��c��X��e<��H4��A�ȅa�����ǥ�:¿�ؿVZ�����係O�⿫�忐 �.�࿜�п�������%~��ES��=:���5���E��9i�፿����r�ƿ#ۿM�� 翊���a���
R���Z!߿�-ͿL���ϕ�
v���M��8�O�6�LhJ���p�5��Ѱ��*fʿ,cݿ�#��H��⿄�࿇�⿌@�	���Hܿ�ȿ��������bm��3H��5��8�
�O��Jy��헿�g��	oϿ�	�%S���b�~�⿠c�!��Y�濘�ۿ��ƿ.��S��Yk�B�H�m:��,@��Z�e=���!��tR���տ
��9��?��Gz�W��U��B��ބ�d�ڿxUĿg��΃��*�g�ujH�%=��F��d��9������ԉ¿�ڿ�'��>쿜�� �������$6�غ�Aٿr���wʤ��È�td�;mH���@�{�M�1n��r���b��i�ȿ��޿�M뿥��`��E��	��������׿
%��F�������c���J��F�0�V��oz�慖������2Ͽp��SD���F쿙��X9뿵�ￄb�#cտc9��g�&$��*^��BH�GG���Z��i��ʚ��Mҷ�a�ҿŕ�#a��[�EH�vK�V�'�����=ѿ�6������D~���X��F�|�H�O�_�ul���x�������~ֿ?���￞@��A�鿡쿡E� ��v�bͿљ������pw��U�vF��K��f�:∿æ��j���vgڿ� 꿊�ￚ	���g���$�￭��9�߿.rɿ���o��G<q���Q� OF�U�O� m�����,奔�ƿ޿�  �  ѕ#�y�� ;�s�e���:˿1!���觿�D��"����c�~@�m9$�/���r�
����)�'H�}�l��Z���P��f���PD����п��|u�~����!�O #�����GYۿ�ۭ�����n�̹f�c2���Ŝ�uTƿ�f��<W� ���#����:"�/9����ۿH�Ŀ�!��C��ؑ�_7~��uX�N�6������U�{���w3� 1T��y����6����T¿�ؿ��� ��&��O#��� ��&��*����ʿ�X��k5��Sg�"@k�a��y���b|ֿ0l�-��R<#��I#�o3��6	����[�Կ����<���
���b���u��qP�V�1�{R��!�L�߻'�HIC�$nf�]_���kݩ�>��ܲ̿�b�^|�tg�� �K�%�M_�����J�"��!�����e�m�N�|��ݕ�m������w��v��S&���"�Y���2��-�q�п���X��W������?o��L��0����#���!�U�6�mU���y�����1��5����@ÿ��׿����	��A�`S%���&�B���\	�l5�Z���}P����~���w�sՈ��s���Ͽ���ȯ�jh$��0(�!��f��Y��a�U6Ϳup���I�����+G��m�h�,$G���-�\E ��~�d�+���C�id����Ǘ�m&���D����ʿ������$=�`c��'�E%�m�F�� �ӿݨ�ܬ���x��{��!��,~���(޿6�P[��&�-�&����<�����Üۿ��ƿ0�%�����O����]� >�k}(����"�513��N�eq�����56��p��9����ѿ]��f�-��i#��O(���!�Y/��E��.�Ŀ؝�ק����v��܂��^��e��<���N� ��  �  G�j�O�a�Q�H�H�'�|��\�ӿ�l������	n��CJ���+�������q��$��Ύ� G����2�pR�]`w��������B'߿H+�gj/��O�re��bj�7Z\���>�8d�F �X������c鏿����oп����.���P�|f��j�'[�4�>�H?�T���#�Ŀ��������bb�ˉ@���#��P�����`��@��z���	�� �%�<���]��ׂ��i���ɿ�+�R7�Z�:��BX���h���g���S�s2�ϗ���տ�Ϧ��j��R��K������HW��$;�9Z��fj���g�M�S�[4�&�����=���ԗ�S����Y�U�9�d�	
����	)���Y�������/�6�M��q�����y��)9ҿ�R�N�%��ZG��a���l�m�d�i�K�G(���\ȿ�������Y��s�¿�:��D#$�-�H�zqc�nm�Njd�K�K�B*���|ٿد��}��%y��cU��47��#�-@�����{���M���O%�-�?��_�}������������ 濕��Z�2�hS�@�h���m�|`���B��e�E�μ����&���~M����ؿZ+�E�2�M%U�U�j�`n��r_��B��| �/5 �H@Ϳ�c��E܍���r�Q�P��4�+��V�������2%
�����0��M�.@n����j���ȿ�����h�0�>�&�\�m>m�T�k���W���6����v|޿j^���똿�����ͷ��	�pA���>��]���m�sk�9�V� i7�e�qj�V������n|����f���F��+��y��/�#�r��L���!��u:�]X�u�{�?��	���D_׿1���.(�u�I��%d�6o��eg��IN�l|*��'���̿b���ݸ������]ǿaY��P&���J��|e��  �  
s��2���=u���Y�TD%��;�u������0�P��q(�pE�
��Suξ�E��z��S/��n=Ծڰ��mG���0�q�\�/8�������r�0�1�d��a���`��E���Ҕ��S��L�u���a�v�f譿%*ʿ�7�W4���i��ٌ������˝�Rђ�ֈ{���G������ڿ�d���lv��B�$���I�Lk�E�Ⱦ����򺾑�ƾ��޾̕������=�z+o�	����ҿ(d���A���u������ s������o�P�9�d�	�p�ο쵮��Ͳ�iUۿhx��F�1i{��=���-���ԛ�����~k��7�O��WoƿQd���%f�!�8�ku�� ����t̾s�þS�Ǿ)-ؾ�����P��+�sS�2���}�����!�� U�,������W��I��/��f�_���*�2+����Ŀ�������V��o}%�`IZ������5��\Ο�����Ն���[���'�#����ᶿ�.��]�[�֏3���������-LվfѾRIپ���r����<>�PLj�Z*��Yſ���
4��`h�c��]"���������J���P������>���������ҿ|�	�b�8�2_n�R���ޝ�����R�������K�������U���9x��"FS��.�`��ip��N��ܾ�F۾`��Q����Y7+��N�f���G��/�ڿ�����E�z�����.��D��� 	����s��1>�����׿�R���Z����ę�J�z?�,�����-���������n��l:�}�
��#Ϳ_��Kns���E�oe%����u����g�Hs۾l�޾������X3�)r6�A�]� ӊ��������W_$��W�$2��,i������ ���VJ��Jnb��?-�� ��qɿcP��qſ�����'���\�Oԇ��>���  �  <	��ۀ�����`����UG��c�����c����G�l��?�� �ʾ�����h��Ą��7Ӥ��µ���Ҿ_���]�!��U��D����ҿ�j��1V��-�� ����������{���E���|�$I:������ӿE-ɿ�?�@!���]�a������}���9.���`��«��Ջt��2�����UQ����u�Υ6�����徙^¾�P���f�� Ġ�#_�������྇�	���0���l�=Y��O�ˌ+��l�z	���г�dH������k���$����	e���&�`���aOʿg�ϿZ���3��xt������y���e��� ���I���^��{�\8ݿiƚ�c�`��`*��)���߾���`�����f��:㺾�6Ծ������i�H�;5���P���B�t���8A������3������@���yx��Z6Q������忳~˿Ԧ࿽���/J��ǆ�0������a��޽������xJ��2Aǿjԍ�;�R�ƽ#�����'DȾp��������tϾ�$��C��Y/�(_c�f6��~�ٿ��L�Y�:���y���������~ٺ�kF���$����>�_�,�ܿҿ� ����%�eKb�4���$������UW��r���Ν��x���6��� � �������G��1��8���⾱�̾���{����ʾX߾D� �b9�pA��}��������t�/�-�p��%��6��tj��t������¯���^i��+�n_���ӿMؿ���=�7���x�8ݝ�Ἰ�U���T��N���I�����a�b�"���㿅u����m�<�7�_��[����ھP�Ⱦ�r���Wľ�Ѿ�n꾣��A&��#S��c��]ÿ�@���D���g����޼��4������(6��o���l�S��6�#��*п�S�c��}L��������*���  �  ޵�����Qͼ�����ra�k
��ѿjq���F��{��X�e������Ɠ��C�������å�¾� �p���V����s��M=*���r��ݠ�h��������\������5O��xM��٬R�i���鿜�ܿ�&��Y5���{�����<���������������������H����~���L{���3���x.վ�䱾��������k��~-�� ���.�Ͼ��-�;q��U��k����@��|��\��w'��i������8����������;�����ݿ8�xZ���J����k��*B�����{���ˍ��^��� N|��l2�񿶘���b�Ԋ%�����Ͼ�ñ��m��$X��L���JP��ݒþ�S뾓���F�Xv���˿�K�%�Z�o������:������@.��)m��:g��5�l�!D*�����p�޿f����'$���d��!�����'q����ok���)���u��C)d����oֿ�Ⓙw�Q���1����Ѿ^���Cϫ��٨��#���y��fXܾI`��*�Yd�"�����-��Gv�@�������
����4��e���9X��m��UW��=����������9�!!���3���k������Z����4��줳��$��`+M��,��̿��煿��C�:�����ZҾ8b��dY������\�����ξS�����a=�U������������D����kx���F��y��������^���5��[;��xV@�TW�����ױ�XO�P����h��l%����������@��Y5������5�q���\G����o��2�Q^�I�辘�ʾ�й�%-��6̵��	¾$�پ� �A��(xQ�ۤ����пD��k�]������a��5*�������n��P���z���Do���,��7�X:��8��Y�&��g��F����������  